`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s5OZXFKbuPYKrhGgnqQLHKB4lBh2zCg8BpJB+l9H/WYqfhno/lOFAzQY61HHzPZS
ljp27H20Hj9FPhKnt8SsA8zw+3J7qYdfWkoPkVH2U2GdtpE7uklODSfcLlmtIdf4
v4Xkl+CPJzf7qdvhnLjbdsvdR+pXk16jR909sS9wFBpaf4jFH75Rop7UtxdJSCCV
s8J0TzOUCaHDMKT3H7Im2G+YuggUrfbr74wBRbTuzG+rxTZNck5ZFF7FUHzXoejW
eLK0yfn6ygUZEMi04Niri60yjWVMeRKkscLHD2WhNAu2tnxpk8R9yrkpmGbhmvbz
16GmNsRN0l2rehGigXs0yV7DVpxaXkvbBtk4UkGvHmnw7YazM/Cbyv7NL4YJbf1J
KLr3W4nLi1cwFSWPAG9477xJXZgnMJNyk3DmhN9OLx3zmiBhXIGPWIV/eQSyUWKR
RjkRR5Nj+V19ntCKWCgd3xaKThVg5asTIPy8xu/R/fQcydCsfVMOfVWZm53l8/Qr
pTHPnqYMuLPpBhdxFaQGcAq23NC8QZr8S9dZ6xsCQPCWseEuQENwRj3GsJQKZ1a4
01xkVujtRNl8ss4iL7GfWl7fM3Hj1jJ7B98yPJq7M0WMfX9ARS51BPnnKwk2Y4Ey
Gckr/OZbmuF77mZYHm1X8XKGHvBONp6keJskatSHEFywiAGqL5C/C/dDdYoUFpVE
YgSIUy5xo1etKM6vmHD2wl765sXeniin/TcUCvt89bijqenJp2DDdUfGtdqCqq6M
Dj1rScaYpBzGzQg4e73iea2f6HIOfNsEg5GZP0YwC8eLDc0juO9jChyrBvjA2mf3
cNk/fx4fP8L5MevvgqGJh/FJvk7w1OO9ZOjunYCe0rjktnll0P/wwzARx7TKt1NM
FORnXuIVjJXbO8Fco8TQwcgB7wS6titXZRjJVETAhyA4ylvTJYv0HsXFiM0DM3tg
OtGUc5HxxFDAY/XMkerz/5D+ATX7E6qgrGGR1+dgxWIbVFyVIyb9KvJF19h8fEG1
MSlnoGoEBATQue8+V0QxUTklv+cct6CSKUEc1ds8WvxE6Ej9SnDIPtP24HDFO57X
18m2b23wGcUk5Xrkk4DzRAim6WkcgCUxCh9UwpB7VkOrA/jvjFwh/es3cmGz/4uz
uJsGku6sGIx+ncwX1ATN0IY2Ah1fnq89bt1EM+V7PAebA+jsjlYpvXCwX+0CRDHD
iKEqv5AALLWfosKUUffTQY9nuC+sIa1DG83a2DTYYA/zk+bbWB99GfM9uzn4i7Os
`protect END_PROTECTED
