`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K8n1PrW0Rrtb6+n2vfKXAMEb0F3Q818l5zcTMVzJRdUPB3vrMtPn0EPwpH53O1CB
54ArP2RpL4gK30fTQhuBsqVUGbywH3DEmDMC+EruvN2vNkD/1jKiRHL0oePkBhHA
ALnEbHBM2aRU2Y3hIpRAw2x4nMaQrHHDf+l2Efi8dJqj55tRFtzNtWak5XYGpU8k
6zsiP9BjseCO2Rtcj7HICXYVzgrhWh3gJlfIAaAFIiKlCpOSgizKvB2G+6yVEjwO
w1Mt4kaCkKdE3uRbA+UDuwM/FxwkrW+rZY94q6SQ10zQeuKBK9CQRpdoh/VIS8B7
o/UjmiQCBUgMETu/6thBPB9xomYVE/jbl3jLucpYU/XiYuip0H4W0eK1q/WoMG4k
/rJGQSAMG7suJwZciq3m6Nmg4TnzFCBh7vCTSiMv9YFbufvKr7QNr81ARBm7iYow
3hyTd6yIW3L50Op0znTho8Dz8akLExebcDhblowedmDiPZ8HiPgiaBY9mg/qfEJw
ToSn1JLZhxQe59asvKTWr0Zjd7chFrLv/IjxmJKJ/AohF71ljpr114QFW8SRIuAH
yeyqVKwlp4glObFzUv0jkisx7qWL27JPS5Ca2VWw3hoDmlgDdvL9BdANFqbEajpL
9GHUTnK9gIjpqB88LBEm9rr698kmOCu+FXIK3amMFhjKr64vv9JyHbt64TxxHwaQ
i1Z0/pE5ecDWnzR5lt4jpk+GYF3DwU1Kj+xdCr9U8Vf1PjdQPyy2Xn4YA0btfVY+
HdPiRdUlkocaezlCD/bVGFZOZGySyZQwI3Aw/n8mOQeDqoHZMPCG+/pV3jKqSkL1
JqcN4Z1RhIAwyo0wkiRiBj/LXW1A6MALOjk8slW/d+qwzlJ7CcH7G15Gwjnmaz2E
LIc6lzhPAQtxsAAbg1mbODD+AmcQwpbTxlkSETaP94HvXb8tWd8ZVIlOSvKW7KvB
68meW/5fU/WL55WDQCshGCINCTrsBK+O3BG9d1PNqvQNDmt+/n7pfcuxAcYx5GfH
HFK+oh+OZV15i0YS5d8ZCBc0Ca+OoDELTRIhyb2wP2G7idS1aWYrEc6R8X75Ng8z
P55y2iFKC6QLUApX+OfT0/AGGJJcS1u6l7fhSilDCotohrewGZXjc8GiMwsxu20l
GSTDR0Te2ZkzyDX3WPi/ElSq/fduiwwbXArNv685KL0MKAn1f9RhfzjOM0Gr9uNi
whLQsPxr7p6lLKeEP2Ld6TQxhSEHMfIbFrZtXQR86fSqNFOfNuoA2KP0hq1ATeX0
`protect END_PROTECTED
