`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EpasUl5roE7pUoVUU7OJNIGebbLdblfDXGWtm544LDu5jF+UdqBoL0Jyu0Ab3Nu7
ZRFyx/sFUT1QekfSEuydvPqUEpVYe/zJqBEPckGM9cD3YcIE6m4M8fwbuaNRYHdr
2i2sCVRrffrCEFQtNJqjGJeqBqL/y1lCrsf7P0LmSjsORtqWqvj08oV7ykbZ0HLm
NU7H+9MPXJyi3S/UraUYzQLe33xG8yor9oje3hURHdySuGqiq6+rg2LzdBNX//Hw
1f+vom69d6DfQjVrIZTymfQLB+FaZRik+chnaFmckGHon4XgxgxCObKam9LtaQTF
m51iaECVnnIsqh1DIPP5Cli/IUh2U62dth7SlVgt+lzS+2llwATQkudku9qF4oWS
YvSq3RLt5QDK73b1eHSUmw09S9RfDs6MI0eWcHw3Sj2X02TbORzpfOw/Y6oJwkqA
6qcwM2LyPBxhgT1uGkI7yQJZUB97MufrdrE49oFNBgCTRE1IZSRD6GlwEQQt0VtN
yIAGUySA4kcuNW5p1LL+WlxKmXbXWhaLCclc9ds/LQuwAWww3LBF3gwNvqj+r26x
dojLf4LTeT0xLJBGnCWanH9JY5MkRz16b0P04bJJe3BAf+KlXMIcfu4fpoytlWi6
yvrPYaOQKu34baC4RZ1NfMs/LNVXa0dptbtYTo8iMcL00DsRrSCfUVCz7w5DPu82
JssVaAi3G0eJbrQvouroRKBPELZ6XjRLbATsx4tRfggSyN17fR1pt4xF+GdAi3sj
2yU2MzOaFQ0ddd5yLJvJwBbAtuggvfntwj1sNCwJO8IWJcmRX19NvfXDUETw5kNz
ruIwArMWEdcdd0eWJ9uvEaXJ4NyZUwdIsJAtRpPDscwe9xqPS3ysEn8YNHhzlMOe
bQsnvPt3q+PW2Ao3D2VxCnqlrtCcBPNATzWWOqVVsVVMZ7xXopBRZ1GfgqpmgTT2
yMBL7mYSxBz805wCmhis6sb1RzfspMrCnI2fHyOlJ+zBJuKbZv0udU/GDUayNZfq
AXKmQ2MxCy7cOSpTAjz2cYSEMGQp4VKsQqSkZj06yL+oZQMfEeiQnsWzFPO/ADnN
J7FNLfI04wSYTXpfQYwfTGtG1KvKYeMzlwPbpOYLpz3STCCP6iImG65ASrMfmR4p
wealntChZFBfE1rsHa5wC7QUusz1vhMXsDOQJflBYfpF08XQNX+TeVVpEkUWR7wU
1hQh8fLyOdMzngWe5qUo+k5bKWw0P5NSjb1qw7RB116CnqNP8nCMqb5XMNgyoMnR
XkdHfVjbJbanYicsu06bkC1BF8Q+5gWh6SgSgisJH5uySef77k6b4VbsMtR4o0Lj
+8kb3D5xdlsR6pDppbFDfTZo48cbLAx7nC01cZP5nlKI8uRQzHpHlIyAhfLhcAn5
c2qdB/3BFkdCrH24hzX0mR+uI8SwpP8CRm+F/uTSh0pYLwOHIU1ZQxjbydyg0kbq
A5Eacud7bUmqrxOH8UPHdJatFSTq0WnXlKz7sFoHzV3kmQToBDaPaXuQ87MWxpFk
oNm2miK2lJtR7rzpwdYmjT05BpmNLVHMjbyjDX87X+VpfnNi84CySdt53YcVYc9l
`protect END_PROTECTED
