`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GpIP0JO2Q/g5IS1s73cjBfu/lsIaD6IIbSQpw0f0w/60IZwuRZzAjMfyTeP+7q4d
2nWroyVAWH0RahWjRLwwhCbtQdGzVKW3TnGg/Ws/dkd6oJjN1ok46K87sCHjpJiL
T4oD1sdf1IvGxgdiqUjN0BV9rDBnndE+oMgixUVWMzH8XfT4q0I3GW68IVH6dRbZ
zk5Kef/eV3xKDceuwtyNwqsDkMl0LEB6oA9AE8vfT8X8rrIWaRYZJOXtzaM8uQ1K
CrmQGPpmqBbuDqifv80TMmMKDZaQHfk0Cyz9aSiK6XjfkVRhlXnoDIghLM/pMBO7
ev7f5gD66AIRVfmS6XT8ErlSP/bM0eoZcRfGedqpmI3STNVOjGnFzYRtOFfpqPz7
kT8QSX698qL75wy3q898mAtVjEs+0XJsB1N38/EJ3iOM/OGCQ90U5SAyejKtCvWD
mxNw9hTUrvlQ6VPGbeVKqM2A5quacfxmENY6vX95Mqxz3OA2U/JtDOZ7QAvy50BN
8Rf44u6YT5L2y62BImjDNHO0xYBEr+Nsrxk6hacaCIqaZm2QaAkbJaBy+oEqoPHL
g8E09uvcrjVc7tAflSSSVGKuQiPPgm6L6m2MJYFAFLW5FLF1NO0O/SHdS0n5pBvK
AFqxMn+evX+wnfXR3PA+b3T5m8j6TtkpIf3AZKFiu2se6wQP2s7wJfW6ZdulPOmB
UCaZULJKg6Q57V7T1DvTGzxVWhAtVasqPvlfx/WoNDT6eoMtwc6fLyN3tQiWCFNe
R0Mm7NU4opzYSarxtO3RBqLXkn5n63+fpZEhLFavFcHXf8XRSDAfuVOK1szT3ETK
LMsVPPuvZTXA05T9aZvjXgBhd5sX2NZ2NG5/+wl1ff4fCj8LPOqVMWlToCm/ReDe
WGrq978Fcnc/yX4xlTlSU9LtByNRTATM+r5pNcVenS2X7QYGREZhUDDzqd25/sJ/
YupobwZ8VHEANwREEnh7RQqDagCqzSPgWPhYrofAgfL40nWyxmTn8vjNhtqhiA8v
Phqs0x+eXeD8YtBZRUmzCSX9nRi4Vnwh52EwECfgCYS+sgVT4cgMibe+HlIfkro1
Z2MSFw9voqkSuzRbfek/2cofK8xNrD4tIrJzb+IP+oa1rq662kbgvfxQV4sE35t5
9vz1WLKqWTC0XTWAJdpnRVIJPz9+vH0Pa8J1Xfse8XUEEWPPPMT8jD5vhqgEaGUI
KB/VusH5BGdOvM24rotiegAUq80BNGkgHfEiW6UaUcaHiCsTGC9+Ntnzg22KW/pa
pzZp7aByKmWPh8MlUlhp8YiV2fD5w4mE1VrlfRvU9PA2wRLaTHiHajqSQUnIhSsg
0T224+bi1m/2AehDfsCXXk2V6FjjwOLoRGXjFyMeacJrz1M9E6i7qO2kczbf71p8
NAcfUNICDP353STqdXAZX4oRzNKrHJ6jjZwY/4Z/fpOr0NDj3Z3+D7WeIMitm7Rq
2BwTr2VI9gMF73NYW1gaeWXjENNIWnLNjbFr8J4td1xCcjNfuVSiIUP7g9On87Nd
Lhy+xCt8CyAu36Y5ocqejuTYXIJ2an5ZdnLSLwWWAdnNW7vHlyhhZ2hf73q89v4v
FVMVtGln76wm/z+57FN3RclN8v+/ildqhNrL3Ek2+1fw9juLKiF9hFIEModmcNiS
m034IMOo84L/T0Qh3waWQtweTnwWggg67stuqTGSnXGd9JT1AFRuFk978z4slGJP
ihsz8MNUlMIrUymC8VZDGFSrQEQjPHAzCoyeQ6NXnTiWXKT/z/YFtgFL9nnv/Ql9
JnDqiRcunIKT9rNuNHNw/ZrOcCUY7LGYUdbQvTZeor9ppmpYHIlAZzU88vXprgEi
40LHGTC+0J+EkpOU+u2h6DsAz8oEoBafSPeAQF9jabPkhmtgSsNoAV3gz9uQ7WI0
AtEuIuJRllxVsAcaHi2p+HCJis/AUgAF30gKDWSTX02mwBIFRgRgXLEtlYXsEkUJ
f0mKK1d3GxrwBl1t7IbpfbHJKCP1xX/ILyHV9EQz4DtqCxJVbVYDQQzJo1ZKuSNv
dejVE4CpRSwRNmzF9XDqrHJVmNkVEWosLnoePoscztL/Ee6uIWXc46q7PqwV8Fyr
aT3McJUikCLH90MM3TNINGyWxWF1EcgLY53gBtbTWZ6Qt7ssuL3SMDNcCiBXSBSD
MD5rKHk+Sp4UCExU3c5q2m+5+P3979Znom/xRJjgr4DDRhxoNVNtYFr/BTus6Q00
qfII+fWVhdLvkjJTOUu80uaQ0rPZsIUjggWTyyhVrapykMZo4FJbi6qshcqDoUou
9Nl5LS8cmPpUA+YsRbmkow1RJh7WQvSwt1IWcPfbmIDv2HUbu1J4i4Ut1xXSraRk
CoBdq0mecMg3lsi70JqKVyoZV2+n+ZELypvNou4HbR+MG3a+mTWNmFn+c0/6nz6G
sfoDoB8QqpPcc35Ro3zuyw==
`protect END_PROTECTED
