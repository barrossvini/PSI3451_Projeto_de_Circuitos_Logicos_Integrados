`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ABywJ5d4Zz/S6jKQoXVqvhidHyBnV07ZJV4dTQBBxndYRdONvpSpyh2Y8p8dySsW
xXgRNsmWgqLrejNwPjTwG7hZ+EXAEXUl8helkYYQ8Y/q34Xr59WRZCBGJuvQ0B9B
EUaCVhyzEhETSSTyS71HWwZahbH9PshJvUggbsajH/Jmty35rcL0hjD0acx/rBH1
TTJXBPDGNuuYXOZSHt2Y4xzGXWjFXfqo4LLhp13a5Hj69b0sIDHFSSLPlT9jlc4Z
e+K/BDzJ0qcPs0mMo1F59BwCwNi6RhLSYyru0oRvukdak4wp9yHgubkDEnGQ81x7
AxaxgWcOOPCDvmPgA0fbi0iLFJWl3UfnXUeqNmUDZoVFfJOin0Ksy3D2wDzAqTDh
k6xxoqlcVUo5vcuSGF/FB1D7YPRql0c8JmLIVvQBXHE8bpdeSjQcKeNEhFWt4wk8
rgb/tfmhQAzYelYjM2551O7NCd4apwoUHzR/OmveXKcdrEOhJXZe20xYOS8uFfVI
suhlyLW7SPfNLeKgcJ51pbb/Od7XtQCp0R/OR1l1VOjTXiiKEZtUNJacrQS1fTGZ
OnYXCHWXEbjr9zA5XKxvD/X++DywxPWT8phGNRm3EymhzLwGZyzk8aL35cYrcMlw
zw+OacrtF8TlpLcvfVwmglrQDTnVvTX1altTYOmiNTmKlZgNjqEpEaK4nH7Da2YN
gdzh7p6fIsyMTcyIYuY7PHPBvDZHJHcJUtfsZDSs1niGYLcJzvPrcIlueChOu0qI
eC90iWDC7tSh0+t1m99HTJ+8amXwBYxSEu0Ft6bWrnEZ0hw+4QGb0FzrZ3ZypZET
fz/d6Gsiam4niTwOqzsVfHWH678zkzbvrYvO/7wJHI89Iys9jHl8ROlg7rEqI2Sb
sbdvCThomcvCva86pizt5bBs+BmM4GT0K1yK3kHhlqA=
`protect END_PROTECTED
