`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tVF3Vg6WTnBThkoSUJvugjH/K6qD1kuBcrP1JBXx3Cqi+c836icz+YATbH7rqvCY
V5SrQBh4v7nUQrgackGUEXyL4E9ZnusyNGrIQu2edqe2KjpDVw0Rc+FTWeH57KLf
rJ5UdS9mpn163JTjpbov8IsmKppDGOVBdJVTQ+PIgVnBjIyUfNK8bgyTkO+p2bsY
rJCgctnpYLg3+CihKLp0CIc3vu2Rki/hgt2hMvLtR3VSmxhE4KVExZdiijCMK2BD
nZ7G7jI7mHfeawWRCYdkTDeEQgMZb4p22RbezIs1vHUdB1lPFpiU5PzS7vG2w7m3
8VDBjPLUPlm1lRUKWfzzK1WrxeCriAvOGSs2gsSdcUlk1OXx1eILi4qTXGmLTZ7b
3s0Hsjn46n0zidFm5PouXtSOa8nReudcxwdndYTTkJLV8lTT5sqznH1mI1eHtUtg
O462CvileCxldv7c+UuLM2O4EY6US/gLOKtUZ4fsN+9pMfIUbOtC1i8kJgX7QeN3
LqgruYpjiMlOX2LxeleTwyIC7Ymod/TpbbT88e7O2AqjVJKXF0N+P42twixuxU8P
HADEf7B0QFAU7CzdaTPkFFpKdhBmqxr/wz0OZczI/VU4GB+KkHRoJZhzqIFEKAL9
ZE0CnV4GhTnBFoLbJdYddwSUT0lAH4wORT06fykM5WCIKyyB7tBh2kEiDf5/gh+H
yukkpPpXMtBj8ajcElfoQdhiV6en11YQZA63NUziVmDHqgYwIEsGBB/W3+D8re02
ogpjxDVR04Xs3AoNwXf6OQFjtDF7rvNrRrAY52BwnsPZEysowLIMGB1pnwDd8gR9
8BeQCA4ZoxWvYgCxia6J/e+4uSbynvBlB5wCtf/bBkyzJ7zKDM03MQgLlC8Kp3nZ
T+B6wTeZZ9fjz2FY7yaAZGUJuIz+LmY/zqzbaoltNZAT93qg6WQvSviCCAFVwe5o
ozhHe8y7bJ7gSf1sUldHwBaEeWZ/0mAbrgu1PO990LyqWod9mukUaoLk1ESD5ytH
OalfcFOBUWSMzGYJykFNyLwOitcTsfQp5NA6ZOI5HwqaMBKWXcVpDXxpqRCQg6Rz
S2Vc/Ad/YuMMsaPV9xDlWSkjcvSOo5Eu1sUR5u0g0Iri8yq8uqgizmGd50ilKWlr
kNofpy/FY1N5lWvDQkg2YBZgJvy0MP2cEHB7wiF895yipIwOWEISU6LyUMP0+If3
J1aoHk/LCYAkx3/lC91DA7BSjRwUefHI1/BE/oCkoJ8jvSMwUmXxJ/SpCCwpNCfO
sjYjy9WS77f1GfDAPXEGGYdnSc6DAjHr8aNavgW7hK5EGFgnnTGLqLqT6ld24pmL
TMswp9CeFHJbWD+BE1YO9QcGZyPG3PcZgBPZtSUDJjiq1M5AfCHCnpAtONl99HxG
lMy2yPFBlnrHoHpa0XLIKK5B3b941vR+9NEpguv6PRQbysG4jK3PpAQRyffH59Lm
a4DpvLp79TO8yUwBBvHG2b2mpCnlrkl7/pqbHD8CJg0fASM0a23/I28uXsBB/ZgC
`protect END_PROTECTED
