`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ytFneAUbcAVyNXirDheBb5dqXHUkFeCQmfglPLKAWa153mO3bXjsTfv77OtW//Cr
nNnihZ2CO7AlHR3imTIt59sjvZ5jZGg1jOMcoHcNxU3/Tu+41S3U3UybyyHr3HEg
HWOnCB7JvdnWyUy5Y4b0xPi1TZBX4kbEWq1UdE9WCten1/00xXiT4IcriZHw1cf3
3NIK8vx20dHW2WHR0xJLYKl9NnM8gXWYQUcde1eTbHCINQ3QkoyaNOoYeank60t4
L09W+wKVtS3svrpnXSJn0jhD+D7Xwvcrr4O8TSe5ddQVIEVtTfrj+Pyc5Q3EAppi
8VBQCg3axGMd6RHwuTWKQw9ZQAHXzBxATz1HcZcrdJ4NB23tx2pV13hYoUzKgNp6
h1qjv0P+ii5+Wxd/etwbk5JvjNEDV6Y2NOGLs9K5PKukyap1rUgyKoBlqJxwlIsT
8e3naO2PkkRovOiExpd0sk2wWzJgWftOoMX/eeD4w9ZPPGAkZcHoa0QLgE/VjFGV
LARzT/cK01NDAqyUpaxKYB52ZzKtCF8Wgc3vYRJrxLcBJe0oUbYs5ottWV3XfHZ/
2S8L+aSllUyOVQF1cYzqlpfHthJWlY3GpXmyQOo1vrCkcamFgR+Mlr/pGnnRM4Ev
gVjAu/PjEUnykERLtMKR0I0hVNY70q0X2bCEEve++ihSytpPwfVqqaKNNeQGuyxk
8Ei603GMritEsjiUYW/hBhvjmmgd16aDKbVg4c3mRwI0XATNDpsEpjlzzeqaSNmH
KpM75RHve5JP+3zkLj2IhXxEbj/l2PnHRVOkB/a6Hwx8JEtjNoTxrXdlppQQjW6L
iUnZ6wgO+QKKmKpBORnUWPeqUXO/4FMNpmI9i/UnYI+qlzXbvPuSOx5wf7RSUQQX
4WHnonO1280o4tE32E1/WtoDBzgZZ5eLpOsJ3/v+tp/Qz1nOsMK0Jfo+x94MDOO9
eCiEjYAD4XI2Vxcx4vJA69oXxEuN63ynAgMuLgUb9X0Og+yy+ILYu1H2yGm6K4uf
CKaJTiMlax9R5vCJY3pseALCL4t5I0Pf+fxzIKYCteg5vfPrUb9pPoEstgStoCdt
EjvuwxEt6VdD3aEstE8a91sMJL1iGjd3D6oYgPBSFpqayymMVlhW38n3ROC07cDI
rMLTcRHPXJbdqdOeyRWVSj9/EMhopy1UyhftMUNd/T1us0xyGGpZTyLCRsTsPLS6
sLa1Iujz/rkBm3j9c/5ea7tUiGAUMvhfvk9XM4YR6Gb6ijUZax7AgcuE/bUSXUU9
0KVu+uu7e7MWN9lfoRoyc8x7RnbA+10K8UdrY5hdBB6JWL4tb7I/pYgc2UnNfalr
LE+g7h2FfdVloSINJyX3EAfYa9VsLwtFfBjqMaLRHLnUvR9lnt3ehno/H24KiCfJ
pPvWdW/F4icGTuBd+cMDwxhJxe5XOp0QFzjbA8EwLEWwRAeTqhIg7QKr/L7PicZJ
vAOsOVXTimQBcDDr8wK5LWc7e9CgwjTbrcRMkNkOsMQOaOk9eNc5O1fwF0dNTE1Q
TqCvaj//gQyCOegvRPNAriWargJgWc4by/RnN0M0Bq5Bl15O7MPjhERAwrb7MKoe
WUNLEgUaiMTPjLrYgOf5WvE44JwQr/F9DdnDvSRrtpnc4BMrBtdvuXJWMcKbV2ZY
5dFW9zI6Xvu6aZzIsKl1SI8Hdw44MxCVjfw4zYLODM9GG3gb7H0GVGCfHuitGriu
Faq/Ql1/ZA6Acf2j26rIGJvqxy2WlfL7vrFvQuLLXOGfAh8ExsKPSwTLhbU7f27v
qGvVN5jzY3why95PSm9PgWeTLOEdWj+cUmwDa3T/cgpuf2CgsiXnyAOyYJKNRIIH
kyDKeqdF1wDbh3twYK7b5bPp+CnHYXl2kwlwb7sNYa5qGBdU+6yxfA3QYp3LrR5U
k0jifSIyNCiuBiermYqbRQ==
`protect END_PROTECTED
