`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LiTWXG/6X9VsYg9sEuvcOcg7ogKCYlGHISyD/xq+ZbXTq3RZi7eqQFzOElNg2/Bn
wzA69ythU6EUOguK4C/Gdk65saONYSnTqgL5Gy/603FR66uLbTAs9Ae2q4g6tOoi
32JWdjPCxDGV4/I8gltNHiY6qcJw7sBNtxdqm9xhjnyCe0rOvBbKsgBFSQ0QMcYC
x7Q6jfFW8pAbkKF5S3bSuN1s6VvU6ewClBOJrO06bzunKR+yOSBaUuYw3s21IhOT
n94qxAqEqRDQTLMK/80U/oTAkd45OHWABEVFBkunsG9VOXBsOFBV5OnW/CZTtk+b
/gTVpQRzW9BkUcAflG72c0APqSuoVwvjVsfDujXf+9wyJFODq8yA3gtA5aCM0jS2
kRO07UywfDG5YXoEfGNECm5IjY5DNc9PaeO+/DLpKA56gF5IahQ/l8Ul1cTMJtwD
`protect END_PROTECTED
