`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S9BBEF3F3bVTO/h18IyjDl8NfESX2q6rhkApUAooMOr0Vntiu+CjvU6PYYiWOXWZ
LgScbqXJN1XXAeVgwjD0DJfpTuexy7N0fjWYkpNnQ+/ugoTpYHgA1h7QDBufCMqA
LQT3y/WZSzqWmhHgH1a48zDenZVe0LKHJqoCMOMWvH3ZgoMiP9DX5qPcPpUY2NUg
f3yRIQ9Fxia8gmTogUOxZ0GI28AWHCjyuaetFaknDXP8nths6cxNlZSfonzdGq4s
E0CprDRz6+4wintPiRLIhVcON+XajJWMZANLm9mg4FeHDZM9CEExea3/PiU2gVwv
fvT2LF1Sh0L6x+3wGy6Zwm73aO7ELl0YPpX/pH6kHkgYOgpf2xIzADEvJ7GPA984
MC0xrpCpn3BrUOe6XmsX8Ha7LfJ5dmT5fZyqp5RcSVtIe64/ukMad4kzHZnraJ3u
1TPF4wzQaOeKIWK+JG303gtvV2MPVq6fooZrwRt9YcNReAT1cCQkIAxCji/zZfYC
qI3v/YGBU3iWb5Pb7gKKVlac6tYHA7fQKCYtS+XQ04shSO4AxA1f72XvuUp1OoKY
omL7TnFpFYHbwuTKeo6E0I8AuO2Jxb5RekYUTvXS/M3isOsjifcYHFXStqTuLUaY
Sp1G9x1cjEzFkAb+DPZ51wIubigPDcPY4ALKEByiOD19dciLaCRqBN9Z71xx+KpX
Z9AiwemNS+Dl3fIRZhDVfmOraDwNE7TUh544EsGZjdc=
`protect END_PROTECTED
