`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOdH9NDXyOTiyF2lP5rFhJUe/5QrZZN3U0UDgi/3mX4FdBiJersaAWVMU6gVvccg
mg1X/cayZyVXMhqHJcRo/6InmJoMo6un8bhzfLpPgHWzohXM444WAUClXHSWmCMP
0824oz0HWyZ8wgywRba3w3vXsxZUDafuQPhBomopdagnLtZ6mvl4tfqtihhYSigR
/eckg1zozpomMCPwpmv6m+XNitKlM2veq6BYBc+Uu01NLbMFyUe4EYC4RIBEKPOK
YEgv0aTE5N2oBjqDKdjhIbJ1MRSgHLpvFKjFBp9LqAmr4mWY8EYWTHg9ZHaLD8oD
2Z4CaSR5vMtl2n21S9e4MQ6V24ZeVS7uuZ7V6WdgTIYLI9MrgKmN5svQdV277BGk
n+zHZzqezDO0VFRwY/s+5q5MOIO2RBuG1YHT5wt8VnBsqKVbwBC0LO01vX/oJhD6
zxRM6GJphlKtWVKXD6v5UPkhsIZfC2nGPrVQ30OiHWvPXXdHGUjTJmoccwP8yqjl
gg5PBHKPIhSselBD6fL+rFnWsrhucRT9p5qVMzIl94jglCC1AWuVEa4XOR/GCc+Y
xv49mYupY14Ox9TRO+srSaoX4hhy8HDyhrG7MVl2HjSIbCdbhsOSDf8MvqsFQbOR
dBFz7j6sySAjNNhtpRzFluX448EFNuuQkKGMgAve6QG2BZhTvElSQdKW3GmtZGYN
jQ188bLkCLUwLOZAGAawZRpiWKlDuFg3pcTXGL54T6h6vDcUXtdnNtk6EP0DHTQO
tjtYtKy5IHKOwRyfT2PFd9aYNyMWjvHQPtB/AHzwOQPaba2u1cSf40MyG6U/1L41
s3KM4PuAimNDa4FDoZvqtpPK/Uv8+l1CiOAM+kpi7YrXmretnkTyl0Rd/M90R+0R
fgN2ZvpSgR6gyWSwUI/fnj/0EqnUQWupy9WWo79tVDagowHYZUbkwmYJVUVO31dr
WY7eCvaUls6Jb+hFIYjo6vvbSHS4Hie1NotRGfOKKD6iwSH3di2D55hmMSsYgtYl
QhPunzYs2zQcVbdVAOQRAtsF8kC3/NFOQUisIZb8l0d1hwhXGR5xPxg51KAdcDiN
uOBDu4fXSYFRn4KPSKlJQGdB+GN2My/ISF5BLXehz13GEzNXG6vGxYLjknCyueOZ
B9JKkszhbJMta0PfzwS9W6qn5+zJJk2maGusYl/LrvbwR+tILFkbiKy+Ff4iV2iZ
dLwHkHqxirZPws/imp6aXjVVBSjnLsflPvC2qxK8cUTctzxSy66z4XKUvd9dQ4MW
axPGX6kBD+aY8CH04BjWTu//56/Pn1QYRkqvb+T1DABfjS3Kny45UC3mGORWH8cn
ZipuAkxgbnuoC6sFgJIZXnpc5r0V993JjFJByHmK0deJBR7fB5ZW90xq6ub07tXb
/yC4Y8TwvyDAspB8ewjeduFLiULtlLQUGSOYxNNvW15Ml1atiDdQQuOY/Zlebuo/
INgD2PJRH8aA5c/j6bTgHm5a9N4NK/2nQ+pjMbxtg2okzUQLFB3OKFCytJt6m2vl
1IUkVUMEpqtHcO9k3hkhWI2+Zj84cvnPbn2Op2qqLrn7FR8+db6ssKSzYwRxMYe0
xmdIu3VsUqk2enf3o5gOtvsSAuVBHacEpcdTBbAGdU3qtGKunQseohuOou/slYV+
zg6KM4Erq6PNWGDMEYuLBguMtLb/uS1GqV+q0/vionyae+ntgFj0yPPp25CFrY4c
DHqu/sBiQtC3IHooSgAPjnu7n7ArrsrAtKzJcmU7OK0+aW1/tm+f5eiAtID3Yq1B
V8bScbrFuFN927gmrn2B3G+Zkl40K45C35dnMGlDdoEMvwWLh6Tk2K96tP6BkSG+
06tqd82rHLbSVJR4PDC9q2fLpX7hLY40KmpkfcM66POsslc2mPrFmHqKPC4SK00z
HXX+jLuZYDdpVqRbkvzLVRanbVWmscRwaRfKcwAjNsPZ0WWdeXJX95KIF1d1NTIr
WO7CSgtArcUhrj6ctsXUUcyjkqR3+BrG7esBWC3cv/4Q48XfZ/u49HFn2rdSZG07
STYfqo/LGPG589QGAICdiY45ycUgOFTj4yfeFQ3l6/FHRtrcEiO0Wff6C8RaGNGx
QKpg35AXC0jutJnXUzAwq6hHoZLL2tE+oWAUsLRVQDGh8jFX3XWIo/Zavr/b1642
MznAUWite/J+T/tuUIS863pxDrYnVmx94YrDoLtarxkTWxFG/BGMOhGfYlg83btE
NfQcm2aBLM4kYu0wEltCc1ymrbHRyAsuR7oSkJNcBjixIZR5S6T9IwGqpoK4U+Wc
RLI/ACJnJ+cVp06oXIIUj6zI9xz7K783aww7P94Iu3CWk5ZoNKxGDBXtGGjJxvba
tjD4zdNzh5qTlK6Ekz5xpJQoXbDcrwAEy1+3iXIsOKp0vJnHnW6M3wyt5lgV8EAw
SWs69W5T1lB7YOCF+zznpnf4rl1KcLf3OgIKjOQnn6ebCM8GgltaKmDlzgFj7e9E
xuUTLRkyEc/RIw0CJlRWh1Y5onqxA/F1EYQdmcPK1czAyuBX/xm/fIZGoalAwL0x
XpXYkkxVWDZikKzTqAY/+H2fl+j0WuK2GPmXTvQIgc23COX84xhc0vcILCnJGrzq
W3muNVShAdQjwLOWknVXQ06KjJamtR6B26WdYOutOSbkRnBtfCABq9y+E62XK8op
TRMwcKwvwsReNBhKOAg1LTi/bOjt+GcWeCX8WFdK7DiGl65pZpuIWFwN5tIWj/eF
cKQurcvlCiIMDb6KQU2vksYKrZFnQ0bN77Qn+4K4A5A/7leioMYKPShoeJDtV1/u
p7iPCpvagSFogV/ieoynt/2YeIT0tfAF7LLgibL3N9R848VmAx+XisEcrmQzlJIw
z4qxA/1fWy1RCbyouZ2EU/4A4Yiemq17dCpEABMm+bm4hz6uykxeAUn/ARK6R5Q9
8BbxvLYehuJClvMlxGMyWTbSMYfDTQuhzH5GrHYSnjgBSMKp8h8QEiOSeLvtHc1h
PfqJPZhqmo4hTWR5YMAXsd2fP84h4oEha3+BPxIQ/mKxtocxCjjg4c+XmXSbLqFr
d1AShABZmbl8TJ1NG+v54t2yYl111lol/2tp1ppdZ3d7gUJrWvYqjjSQT/8mRUag
RnsRud7PkuvyYLdD2XIGfFj4qq+fEzVkT4oEY7Ind+es0Zig+d5w/Y00W5jgMpg1
EUTcEIcU3cy3o3RZ2OhsGcmoqjWfwvidijKLjmR3+RpyJyU7oppg4Gp+87K1dW3N
9AS1YX4sNy2dm2wmSkRcMfd/M5V4mBUDak1E0CklnM51UDK0uIUVXzL2JaG4AT3L
sjklSOCrz4Cqpv/h1wwhNGO+KdhqevAT9W0DUPDFjrZOUZihdQ7riCC+KgntjPa9
VD4/kXkLXj6uZTq6Zq5M9pr1ZgNyLx1eAwkUCzchw7HURU70G2EZU8cepsUPm7EU
JDqvtpKaHma2JhrVJbuTbxOM0LMebh8zxwGbOtbFhs8uJk5LOh8a2l4ogJ33HRb9
5jT0v4VPa6BZz/ic7JPq6/kjSa5S2DbWRSiKu41imgUigYoSrMFQoBWMadaSS/8a
i4BWtiUpJSGgtUQxtTh1NLPwqvgaom9woQIqbu3rail/HfJYxfitA1wCRN+nVfnI
6z8SZaDOP6ILE6e6VGuz/ucfMvSHDCrld5THWlMVx2YwFgKPGCRssSapnuHEL4Ob
x/cjqat0mqu++z7onKSf+BvlFoSKrIahNgK6ScUpOx/elC/dzICw0WAm8dOmM6yw
KfG1pRm163KEZwSq1g7zqj2mBWzckfyO3SdCUvmY/fbypI3RXU+hVRvdW4AHmBzY
jq+5uG55+akF5WQmaycLpmbnL0kohh01zXRwmLGR3LdGAachP/BWHH/NO0XWoZcG
eMNgmSvG7WBB1Y7un17x9pvxYzMF2NRaQh97M8HrGcKIOkw6X0YvnWMUnsXSbpAa
zJTUQr5HGG8ZLPesDOd07c3Ma+/P5yv7X4v3t9ZeQ+lTj1r0O6nbi/dN0Cy7PKUv
cNDpHDCxTpMMub+wgFBK9bh6hc+/G6AN+iobK3nXwgS8RUvIDdu533iwQDY8DOMD
2tbVTkHddE/MVd7pyLYICWIUnWQQh/cjQ4IbVfWbdYbjs/qNh4pdxEku0LCd/xuc
g8e3tIigrcB3B9R2ZbVUI1b4msISEZW+lEO8J+V96a2zFHTgixXr5tg0SdXbierO
AavLR060jB2Tro5DEoYG+0qwjoQBJRMKHJoGcoyrqsdjwQOv3Xy8ehpw3vTgdXx7
25HBDtXbjtTUcXFmnXz3l7v6ejmSi4cR0auCDA4Z1BWwoEYhhXa0Fb5eU+0iZcMl
nRy3FlvuWCQ4f9m3GZvw7TNxlLVxTQmmhemKXt80xRb0K2YkH666qZ5mt2P9lwlF
JhByPyI2x/jwLcBlbInb0DJov+Pmc2MicXCjRG1/j90SSd/cAQcGk8OxhtSby4zj
3ndkffgQW1UW0+k9bgQuwtRGWd86W4emug4lcd3rwZe8R7Nk2QyJUDpCX0zB52tF
elZY7Dcr4776H/cxigpwevILOswSu7rYDXnKeSFHt2nD2vp2qqDrpsT7X4BI7kup
4fJRhv4hkxoNdHWAYolIFOm3Bg9+6Rc3XeTA56wg2W3pgLjTkJ8OF1ysBSoYn6PQ
twTdX2Ibtrv5Xa06LAJWLXAHWIXfQCeYmlZ1qfTVSl7DX1jl4omhdg6hzVNFK9Uo
eLaAWP774OFTN+n3wFM21862w4j9ipen4Nccd3T5/bbacCq/OXFb2GGAhcX5MUns
zRQ1XHZFqXqRKWeXM+2UFGxGrZ52JwP7vCwgdLDl2BZhXCi8KaUvPHZT/ZKsCWRj
o5Pt5hS9eeRroaIlCIUU8s/Gneqkx7SuR8WDVjjS4CGxnZfT+prSgLHE2FfuRigY
VtF/Op0p6AbvMkKPDKp9WoC4xfBcCX6SL4jBxe2MMeVAOXMZd3K7wnaYSrmFMmgY
DOgElc893UyEuHjJ+T08jihc0PimvPnAWYKNUhKAcZW4l7m6wJveAT85OB1DdQKn
iXqDo9lLCvirHIVUgqd6JHRCFdCHrS1R+P+xVVx5I9lA6uxVg1ku/HF77Rh/Enp4
1ZiaagxLJVzJOYSmizIi7xPKj5rvALSnbMoJWE/hglrAtrzJTczzKuVrICAQ+kwq
NoDzaV/lN0I7ntQzd9/f8f2zzoqFp9A/p5OUDKPATedf4DfkqcQ4CHzsX8JPIcqV
FUNI1z3CbsYIdBCSMQy0x0zuohUJJOFA90U1MQJgCjjFpqyDjWOPNxvynkEbc29y
T8tA8nq4Nn5PRXR/ZjmbQvTbr+ByGmbn29lHm5SVgvuHh6FGU+QUYUf/3o2+BJIl
25scUW0BreJEFnOQr4poeQkKxuiAvVs/XNEF7a7bfL3WyKPMC2xFCGuNvn+mXHjm
xGLah0xuYum5RmADYxNTHdaLkPq0CW3un6FdJ1xJ3bQgR5dWf0eP8QGpkeqx5WMV
vQmwJoAYUqQP49K60aZrf+u80GH/3FAsaRCXhw0JQXfH5r8+ISHxz8bnzblcZcJY
iLZQpkAbJOs2tg+8NumIaWaR6NpUM1octnBO+E6LCdLfNVeG08uFkuJ4ISHaWiLG
6iAbnq4/gtV7cGD3L6U98pVfBTXYOUzjQU6m5F3w/HM6imwTyCJWD9P2XAhSle2M
78u/YwrKgchD0PSdnwPmn4HZRo3AA6dxHtl3TUD/xvSndlsCRzVOcinAZkl+5cLn
iIwYEK05OT5g4JZvZx9Lis8hxXdonGTNGVN063HNLKNvnHxlO64pxQkrm7E4tQsm
XVfBCLQpjxHx9THwWMCTPhEi/Zylz8L8Hu+Tsh0O15xEGjv9iM4jnxVf0TwPdDPC
5z34laI8JGHj23uCd1PsMxxag82s53ePoVG0hsXut5VRzmPuFm8Z0Hta8PHAivM7
UB2Oo9yRPCXuOeDTYuWl00T5kWOJRP2H2d3ORaVfS13BVnt1S60egyTSH2KnNxQ6
5lfDizoqSgaNtdX61YcPW9wwHcMdbniYTeJDFLTR7tvg/d+2MGOXYBarQPDdj12s
oFNZhUjYsbB0+ydwxEbrMm29NiHH3Nw74NZdYaFz9S0hzIIwy0q1k8qFFlSWPWQu
wKQlIFElz7tZUGFmqb+tAQzAGuShGJ4jrNTF+yugLhtg+t0bblSGGniQVkstRoDj
Nmxq7DErJZaW7XaicVW202zNOQSEsag97/cpsQzygibYgY7uUl+1AsNvgWyGnYkU
PkEpGlC9eMt9lJAPy+Y0xmy/4U9isWGLxJq5/wKgTE/4oK/pPBOFbguzjqUbfJH8
1LpMHL1uXCtO1IMzN+fjJ9nXWGQMu7Vvi3Jt0GClis9xylh9OwBlMBE8EVbdacIx
Zpsm8fkqXuhTGE5nPGBb2nf2A8FGS52a2CekfWRaKi0hyH0vlknIETkFExKplgYL
y09xMDlRavjHP/7cnwC2DerMPlI3diXU0eJBX7UGLj0+wXf8yerzBm7slLfMuWeO
sOzV/sNx9bLk9okE0UD+1+Mw279uzr/tvXu0eS5LjfFW3tgMoIgNk0FIbcymGDpe
RVHGlA3J2mgeRd6PMPl/mNJTLZCwHrufCB72L5YrzSbHFX9/2olYk1aeT9bwZkEC
eql8UwxhmaZuv1Shu9bSs23yyo1IXUrGwxTaO5YUjosQ88Fpx3K8RmYlfsgrn6MT
EVG1sbx8kyzMjsjblFW6upRppwzdYTtiYdiSx7GRk/pca6sJTvMHWcJKpv5QGBxU
13YnIhsw4eM2JRw1UnxAMPdjHncRn3uyj28w0qZMJd+ZgrbwkBFhm56DkE9BJwHf
wvWuAsPxt7qL0sMajgsHPKh+ejFEP7AJQKwSRvPJaykt1hqdpg0tikvpzMDZrL3q
VpFmumajJ11OCBdsmoBSfX2PXqxSFzo3dJXB2lwSzjJBS67QS9HsemYQO+5E/uC6
LHmhGkl68m/LiYiDyjUn/DgQWs12LYDpO1LkpzdTuvf80QSfPQmI/RD9OoGXUD9I
narqMFlMra8fsml8yb8O5T4qsgN/RuJ3Is5pnJZRhG1aGJmoPl4rxYggBvd0drb7
ee5NyXMYMr2/IrPC8W6imOHu8f4k28I1vPXC0xIt7G4KqcVWLbqEct6WPqWFGJ8x
0Al1Nonq/Ryu91pI5nXk+gIW1AHdjxUclLUzMG88wlRTywK+YS4LOamOlNG5Evwb
60Wr1a2Q3gHiWtkIyCQEBGqv0mMC3QjTWIfj0+xnNMQZfkITShdYxnFuYtiZCMbd
bS4g3cfcRJGcwKm2nwFi5RoHJJ8yjWgSL56Iqdp6ddb/Ciq3qmR4+4fand4ssRJ8
WtBVegPvuNeCj7j15oBfgkyj3LS4mYlhWKm9x5GDnHFKjKmUZDFfylWDJ+MpmKp1
ge9/Uu0tTFnek1AqbTt+g47iakZ9g7ueQht68kaDNQNWZJTg9Y2iUF+7Jzh/JTOV
G3toxf8BsbK4loMsniYCv4b6abMPQURD3PfO04IgUlWPLvWicYJD1lVSm1PgFuvt
vZ3zM+qYLWtP2L4CaaJqf5nYdcHmSMEvbwslHBLkAGbb8eDTyNTmVPkArfkLp7bn
scSZInX7s1AECzcjM3dZLGGjN9RLStXI8thjhHUr7I6gPp1ZfXJOR+5lMzB/3PWR
JuKqo1QBSXkB1CVlIsDzd/yThFxHcc94QNlUOKuPd97U9ZcMgGS1KtZLN+OmJ0tb
rlii2AaQbc6eFok+nE4GaOJ9AXkhSyjYmnbf5TrCevoQJ+zW3lHQ3PYDKW/fTe3B
TLFKO5+zM5/nJvLE79jJ3tXkomnpLdUMm2L5SEJz+qcLMG9uU9ybSHoFzTkZrnSh
Yqh11S1mcSN/P+iOJwOZ+v9qEehf0qki6QQA9FoXr3Z88Iuxqr82vhFozZ+z//fN
Ar+dTWWkyJr1PoWQKXmIQDExJTU3lIIqENundHVmjqmN9qohmLcFDkmgNg8XHw55
CovR0LinEGDqkXRK5Mg5NCYZ/7gxc4WGKmOwI8PkmnFcqmvL5X2feBeS/bmlliKw
/4aE7sBb41Jk0Fog3szgYdnQ9Z8ENtroBYce0wt0R7NYl5DrmA7PdjAfh8ziUQiN
597PkcDrvKx9QpzXnoqD/Tb/u3pkU84QjKc66igsXMWGqfRXliILLgUIKBarowiN
f4nmtyFe8maZYQpYeYbP4Bj2Cb/X0NWCkZlkEPT4TZ0pxv31+zfA+iCQXOlPPM3K
2SdVeaD0zEFdE1qBLpmiDAunfG6C7JoBipdz/hcgyTj3dIgRZ33RVRSQMKMytjNP
ArSlweRm1Q5kNVpegJmQRWTDAdCBxw3MlbshZDX2x+vyDlgNjRc6lDlN/kwM6rxT
GsmZ9TT3sTQXW7bCcbqfHZuJJh0aO8Sp5AdOM04Ac5skuz8/pELE3veKV4QszLLt
0lMjRxMl7k2j96OdBps5R4Gve6z3nc2cB5VajKGQ4LN7xV93WDgzxGmNQERjg2Na
Za9fswjfATTkvI4EtVjeBD+xxcB9l6F9goAOcFSUvINB9PpctkrUOug7HTMki82g
n3ILAfSiMbngI/DxKCGH9MXRVjQHkBeV+yCcVdgvEPN6U/mpGrSd7iRiDBnJqPcD
akbxUUhkY4bM2z/RO4NfkvA2viURZt4Y5eXDxaRlGQGnuPAI7nQ5WoWG2r+qRi1z
pLi95dEUkGwzibOvFQKTWFgDrEwG9plyx7Jr7k05rObMds2NZxzvrGxSm8gW/fvr
xSnZFUGGv1pgVB2eA4GoEoVEMUTxIoWYD5bQXdG2byEEzZ4HcO1MV8B/+aKsGX9n
tDKthcIt8+KHxxx6I2ityG7qoqzABeg4A28psXLzdNiV0Ba/FzcwrZyRwbN9zUPe
wwZHbANZFSpHy4vLD9TIsb/AWScHG3xUzjDwrq0Qn/3ubvFbVox6ETNuwPyJrL8t
K5dDKjY2muiFywZ9I2aE6hXHkaufrCPfBTH1l8cn/WPhOp5SiHSIuhd2p9/bfycf
r2W245dzg71OHjcolC1ykZxlUn5TysFIDszU/fTxCA9ZOd3AoOsSzovaB8BvKT3e
Lt5ixj3obuM1TCdNyHzJfAmPDvONGKSiWnaCfEVLXvt67paA5Fl6KSOaKh4PhdQk
SI/JHhZN/z7vZ2T2oVrw+m9Oh5+cUqdGZJodgxC9W6EIt/JG9G8Fi2iFdbZTpxxz
KYNuawMboUZ7a/clT+uxPFmroJXHSRzfJAqFJmz4pSP9Tf9qHDwAf5gWy17SYjNZ
zDSFkAnmA35c9BE/b/IBwPdSbiPSOWJY8I97AFQsSMIBgF98xXn8WVxzgq805mKR
Zp398yxCAV9D+WgLxWMmmfNgKT2oXUqohhLQNHuByPAib7ZKrY74ockAvDF3n+EW
57eDRrnue/Fe/qSkfnwgWJsyh213GewNQKepZVmuaJW/MhUPclNM3CP6ngnV25kR
vCSn9lVipdUCLE0qwNh1qcbTHPGSsb18fwjTWxvtFG/GuBf7fJItw06bIQXRtUoV
RmF8Xfwsp5Ml7Zvpa40YXY8VHRMVARrVbLfFgnLJtNJp9P0MHOIhw+NuiynDbRDG
EYWc9bVZKknLYYf090VF6pDdxfpsKzT7qAN06VMZ6NlGF+CuHqc5IZTpj+3HSGvI
6ISqeviHwsBbiOHblcj97zEXnYDUW3SLSZRRHLwNrLskT0Eg+LQEzY+zBpmJqnkg
/h4/W4MHELpKy0jFXEPUBIyS41Lqkp5kjkdRXCoINdzWCT3DLtKcwi+qfheR254l
PmaYSacft5cOkt4Bgudd6YPenYHpcLphb8r/9R2Ljejf1netGbRnmmWI+gJRo4qo
njptKgZIAWU3FwYwfCTH4gBBgXnk123luKcjAC/MuCjcMrcVAIbkAhDMLZRv2qcg
xbcSycDxeGL8zHOpwL8VTGGxz8/8IYb1DEzY0MeD3zFoTN2rLnloIKZCCNVE2+wq
g3lobkst3/d78hHdawO9xs9/4MV7j/zcbRq+kc6jyMaTFQhFG//ZODz6ME/R3led
zN3ww4e6X1sMTSImjpQ3DsB2Wz4QlHpqrzDBpPRaFy/CgknkkRZ+Nf8BHTdPJp4Y
5svB0FikwHgLiv5CT4l5Ds6oHZbyWP4Q9Z4guq8Ha+69y100qZz1HWm42nTc2oFK
Prurzyj/9RjyzyYdzzgaoOLmx+oP+67+I9gZtaKNFvBZSwKNWXOb+SUEcJ6IQfCW
vDlh4HvbdYrPNyPXMKBj9c6E5mAlxYbq8eW6FkwkXu2IxG6EKfSgDa272xdZ16Sq
ae8Ejso3uvnXZ5HL5UOESKzpadcx47FdQOywX0SjamoNyTf4HjCEmKhmc4C3V1rm
leCfAx+GY4LDJDDXoYEm+fQ9VdKCQDwL5feaSxpQlczybB1E9zQhmZXUGKYQr0Gq
+k0SDbu0nlasfTVU66bXjBWbhGkE01wOldGbhGmVf+UNUWfu5BWVAMAR2NwvkDWR
eBtfAtA27dwWbJbrVlk/FTlKUnQ2ida4U3MDQb271NmFXEREqza9mtz5Id4nuoOO
cZ42pwDwwin8I0E3dIaoOeBrHJBYTzVBQfXUvIduFTdGi5+ptKK+Co3Dp6n23qUV
SF8Q+A9DPfxzUgktfqqUilP5bBuIHDbVjFFiFT2S/TSDoLGq6Yg1JsNrVZ6MP8Mv
eQ7bKUumRBZ2fR7CmWp0MiErcQzbhGfB5vPcBOJEWXCYSU2o461VuIi7dj0N2l42
eydjS4LFkh9Vc2D94ebL0A0RLsCVw6Aw6zjRnKgvovPqeELtpNlNihCX4xLCYltH
b99CU0zbDKKo9IINyL5rLn5wSsJod1LcNpj/62t9cwa6iuTCo+ZmrLOyY2MM4UPP
NJGN24dTGnSKu8m5j92dMAgmwgFq5SuJP7gVU/lSabI6VT77YxLg3B8Wy3Bujs4D
b+SSeqASjTYGA9+nfSzT2mNmOmPvQMmciV8JxNzl/LIBNSVSxZf9rmasuZdJV7w3
6igR10AGmbKZpQrAVSDmzXBl1Vy8Ytghr7UEYhfL+E6XSxRLEY9QuETULXQRecAE
rJD2kvkDEhTTE00MfyMrUWezr9OVXzv/N0gKY9PsI/h3BMfZHCkC2JZHus2dPyrc
HTBWHk7uVwdMOkXUwMw2xcBYk46wDBMOveUq8wZ7ihvmPIbIMYHZAN4b/MEXfy9M
LAh4SDTQrK4W4BdArL+A5q+Dbe9ESfAUB97XnD/G+j+YU4W2WWjdAFfzOB4gvb/N
m2uf4cPyUqtRBuYY69q+CPHdKNHR3y62GlddMveDeOAzBct2Q7Q3Rg6hmJnXsJTq
v85F9GAg3CAtR1q4A7naPVesmrJlq5JKw0LvEuVIU2ZyhJn/jQAuTHeOcfOUSOnp
CJQJVUDGqu70Q3Ze2pX6OMkeC4CJ6VMnXMXgN0cMo0dxtWdMeqn7Ma+Tw2tru5rS
eV6kvrUq8QY7Pjm9UYbUPXqBdn9XH6SWI+wqmDoBycRZVNuzaR1jrDGXiQFN5g2x
G1cGvZNrX5BbjTRs7TL1/GQaTC+WOX58ClUl3Aea7j+79cn5nVIcm6HCUYQ3+grO
xtFMe+3aKRPm8ZlUC2/Nn3rSmCDhrFXV94TKKW+Cb4yn32lLP67pl5ppoYpg6taW
Xj3hDbGU7wMfdalfoTe/g5t9Hj5HeD6QSHZhwcv0nSeg/EeNkcBwJZ9pxwgItTkx
zjDHgAmn4gDdkhkXxonNRuYt9gqkXb/U4o2GxhKvQysBQ0mBMLFjE+8iNb2evj/T
YEOOAspGxY+LmxoAwz6kgUYJ4JtzV9yqjk+0oO4sz2aYbKp5Coybw43BMSBbgyQE
DrpIQgf4SCZdenFFDurUxIbEiMW9YE5/Ttx3SfETNIDnkWWbITp1G7oFMP6KVxmq
PLm4xdTAapP8tKDieMb5BqsxJLx9kqKUmjd7DgBuU/QRwmr2QV+gLCLMKuoDboYN
I3bqTaAYikoabKfHC4zdIPhHne9wBisARnoskh/9lvWq0zasjUouJQ1USn0w/5MP
C4Azu1v9uOzM/NNmUTys+Mv3RhyrKNKLg2WYRXBPF74q7D0N0GAvZZAtizNpd0/B
mm3tOmZx82M+Tzdg1C33gTCClWQYnL/tefZX4ueEDuFW1zCFJ/7WLaTNxRkSr4Ns
oEQEZEBWHG/xp/9OOQkMRESm0AN/8Dej95VBbWkF4T0iZfnljPzWaps3Hw96fJKd
2bJViYEQbV7dxA0tpKwPQQ9SLnJdFG7JYWJ+BP1d52vxEJ9vSFERDPy4tpPwK1yS
F0cB4pt6lPfcdJrTi6srJzg8JM5VbiKJB3z+3RgvXADHi6XWfAOYE3l5OfEB1khM
Fc+0ah1rXky9wC5eZpQm9xDw2pCRQFtWsP0fgpSevt6FuaEKahDL9RZXtnnRlBC2
XkZd5YM2706YTtK4KsazIJshqNA6M/+BQWUcOhGY5ZNQHpOlZVMkThHi3aFRc+vj
Rqng+lEsTR5nEslM52WPMgTiFIB76Ad8ugf2M+vZvMxkvWp9l5r3RHdOdURkAush
i7S572j3olwv+mkNZ2OKydndFIGz89RuUjxhL0EoCT3211qnFAkkFvhaVxQzuqjq
nWLzAyTFNfX5uMC9gVdLsYquTjHF7OtYv/Xk9vIGSWi6Bg8Wzfkovkrk+FhSKeXE
G6sz2U7Vx9zmGcC/pv78ZU1LtjexHayqY+vUry2hBe3l4CQPLARFG0YfCm83SzJ9
phEJUes2at5idsgGWBCrDoKHHpIcq2ywNeJzKFjOFX9d2wlVxtm1CiTDJ5kbuSoE
goLuUc7Ar7CXrsfVRrTBDaObcqM5c+i+Nt/HGgP2mJpco5nR9NSqVggaML8+yfKB
Q6lo3teo7o7WDVltZsbv18WD71l+k7BHEN9xlWQk4BfdBf/1EIup/cktB/3k1Mnm
mPXBjWaJ4JikeY1yQAsraN5+v168e7kKX5V11FVjgk2lUoWFgPSqZvYXf4Lw1jXh
wxCS0GIb5h2T3ApiK/IB0vUj7wp4CFT4xbW2CS2Hxnthrc2RE0o3BwLr6ZeNaSnz
rj6FPUDY5G0Y67tclHy038HTQ/30gp4CGSP1xcnkO9V3ykmSb+Zn0R50hKWEO9Z9
xLQBRSxgH3jh0OtWPH5Zv3RRu0X9lTJPDpiGOs51X3JUI4acfPQzkwt5+FqRIeiy
8N4Pwc4GYr+S5S/qgRMlHVEF0GbxZiZ76fEyJmn00dFH36pu9NF6Z2EIfNsR5UNQ
+dBdzxtRbXVDcmDclQ2oQFreRMhsIsUILx4SHOHShvUdtHhPI7GuJrbIFUNmjlCF
mD+h4lQfu/yHeK5RHeZ4JxD/OsVAXkOQKMH4iIqLNPkNj6CFB0yrymzY2JyE+Fa8
nGWPMcEzHn1YRT8f1uCHG/2x1sh0aJb5POi9t+QBX3pjG5ooOMFZHGRxj2bZJoax
czWYAZ500QxFeCLefN4koo9vgCZ6kTSdpqDq2eXBRen79O+eHkkvT54D2E/wU07R
xLkFF7P4rnirVRfF6bbe1sEs6lMlfeex+8Hh0RTQHiQPZphOzuJhtIMRPGQENb2t
hAP/7avdiZUufScFHZi7cSxxrzUJAGwid3Bo/lABJQ9d09AsYDOfdTF3Az6K7Iru
gagVb0+DVcfwbQauPRd+IEaijzK1IjLOH4LbjZbmcJG6yR2a6K0CI0BySE09H5iA
9KdeZOdfi0XYHUg33IAO4EOdFTCX6wtEL5o/E13rKzk0AHapOEdPot4a+pHZYEDK
g7OA4kg4r0eYw0/GbUydWyYUiDwnrfFGOgsY/c+N+NXiF17TQlI4pUlS7XlTQ5g3
hTmKZJ+AdkyEQUypAO0s8UuTT3bsRjptiTv3CQDX/pyXWi1R26nLYq0lzm8JEowL
IxziiE1Mk6t8DTBLshY3jNMqU6bRJ0GtjsUB/nPTxlBRIjAh1Cc8mAVwvA1yXV8W
puIcXnIFucEC/7YfEo+XpakoVKaIcN+cgw0uZprkX/q4iXW49K1Z1x5EhWSkwryd
XX2JEHMQ1uPrZbUNVrC9uv+duyXQaBCVN4p4ozGY7uzuW2gpZFKeAtvclIVRTY+R
78CkOSZkTpXZZiHnV2do4hZWCeaGM0lJscpKsjxL5WGMasKI1NcUShaSJ4WvEgg/
pBkxBiy4bpBO57WtzOyTuS1+vvNYPZFQRvVLlbwLy1Zq2Lajd/2LlbCMU6Mleq5e
HHbc9ezZZ5yfAzhb7hNtYDsFAIFIYDuzLP9iV7oPlPXDXfS0sQVKnvJXpBOhJ589
FOyPQIdrUML2+xxQGO+zuusVSQ87Eov5L29wC0gFAsxtehZFHo/P/K7Kx1SDKUFv
kaG6SZlIdHJge6t0awH3WIx9gbOoVEVgn37jYx8uTc2WgNG0mzteBvFURnP4cN1q
S0wW8rAV6sVzuBJgHTJEIv//g6y6Hd7aplAfC5LssUX+sy2FsOzeGGKH2VKkhLOt
HrdSlEIL9NDZIirx+5NQ119zJF1h0ZnCAVXabg2a37PEbEWJwGr46BKaevVgcWuA
On8PAUT6Spz+5peZOQZ97cFSUI0uHDPwl6Hrze0wlVATg2rSsvT3pRZfPcX2p8sd
XLo7QwaFg6zR1GUw+mbZbHCvpOrVLRwP+qi5Z93l4zZeL5uue/2w1U4j3DKL/wRP
qRm3eU3TTXul2NDPn0J8htiNfn+Ou97xRxImiBNxh9wVDAGkF62xCmRFdNVpROtI
O+7uI0JeSnI+ePNFaWzvVfy6i0gYi8eOKDYaoFZ7R+mhB1LhrRwulS7DGpgTKBtg
lrrhACR6Q1QPPnziO+nEQEBD7MvSqck22rXqgFXGCZ6UGdCqbqm8HIhhrt7fNagO
wIRt4oQFPBCZ4Y5fCkS+DdkZuEWorUMTXTbEePfzLyhHa1iRwJV1bpBwCkLzT0j8
IXOSIUifbiVaWmGTdULYchgXuKgW1+mrrJCNIbPIjurLCK3I1NV0UJt6tz2V9jFH
jaYyimeNr9rswwEGen4Qv48llfqzv+DIbZa1lGG2mVOhriP/ZRnUhJ38D3bKBmgt
aez0fkcU2lXgaKNKq+bJlGT0E8otY/67/nN2lxmTiTA/Sk3qmXiP1Nv19eJ7fYlo
U/e+gZaLr/PJDNnrkwUFFiQTnRnbPZdkiCn7dYJPBuTh68ZKMWL8deKaHiEEsOpg
1i8TBjrk78Ld4nV86CU1Ko/MjHVRg3f9u7eGsNJJoJqDtGQQ7C8zB48RtaFCpWWz
hiyaGPjLBZoaQsR757hhGrO081wiulqbAa1aDnwZbgHYJkkyRAb/IYCdVKRp4YJC
WokJ+nsIfeVWd2BXOAJ87e94R03bz73AQ/+uJ8aLFV2D917xnX6HCHW9/rd5ZZc9
LhiQmnwOaefWuECSBGnnhwt4clF+J1ZLcnkZPgpNXwmGH8ZFGDL5nR03sxx+uXqk
F9Jtm8qDM3oJ5aX1azYuAw+42YNPEkRd3GUHUIy74tpla7uf4M7XBV7SQSutW6pu
A3G9lOZYpKAvVG9/2MUTEnlT9k5a9Q7dgHzEjDAH5rWLE0nQCYkuoALNTSzDZhap
AOkqA5nAUx9y9QjIbcHYm222MhiIcKZvwkCaXzDbAdLN1buTyo7VDTxisKA5H7vL
Mvj/ihz3SplNN8hvgdLRsktPI4z+XU3yCDMSWlh5ggtnoyCblwNFK5RwLtwmlwWk
rZSB3HLYBX/9vKxkEP7YBItlig7TTNFX24D6WpEUKLfo0Pz5rg6oUzweKJ8UCSUW
Uuz1oYE7WuFgvSfe+D2jYrxebJbVI6xHxPoXNd9o1PZdv1BRaMzdbCchnK4lkNoh
Hg0G37o64IDrACBcHQjXxyzAKcAO2chicqyz8gECGF1cCMQ99UoAbfsVJ0pv8U9j
yDOvl0lMugBw70sOrsojTQW9Sxpw+lH2UsKWq4B8u6aaopvsh4bDaEquRE1v8gpc
GFwElzR4LtPkFzbPq7lWAj3oyoVcE00cwWuE2E9/TkK3L3l/+uKI3SV+TMcPzSdi
0kqku8OOb2UDoNDsEoEcJaMfDfmUUK1WvGZpPlhY43ZANcHR2SDzW4hadNU0eceA
uMIzXXzxFJ20Y0HaGgStVzBygKqk7SLCir7MEcBMZCaY1O/uupYUm2rjl2sMvAqs
XE4fI73c/dMl5VUg9DyLNhwZFG4mjceffXvTCoZUAqyBT1CyGLQigoEhsfXUoPow
VNQRUnEgQ6ObYLByQIDskPTp1xHl4g3fXqP1HNiJqm9Gf9LjaUpT1u9w7HBO/zyc
962QiFLWKZcGhUBBkfvhIe8PK71vkg6tiswipc4eteWjlDvHSCEY+tDU4UbhC23k
j5F2xIJD2RscjK2oyQkhDK1NT3YRgl2YUR/vjlCEDLwMaA2vcPgLSiXAR9b+oEZR
tx1bX1bjSpBT+sCZYgtVr2N5zvgL17HBF4GbYskuFx6xV3tgq2fSNbdyLonT0pMH
eK242NVR1QI7XeaUFbprngfZduLjwtxAGPk0/FA398pGyOz1TNSdOHPmBbLqzEJt
AGW5vsiHPu418URyh9nP2i//q9NAVcxCpd7ZC9PfcB8sDGE80134oCGACLKSGOTk
LQDusF719WJlQNPAnmUMtNDHGv90L5drgrAtcwgib5Akt3Sfp4ISB8IRx9UskHzX
mwW+4hz7/h2vIgNdLEH8R4ifxSHKABpxZ9JzJ4QiXpxhf1tKVyQad1MtR5VgUVWI
F/RCsPiwn7b91M0/YXgyEw0o3BnxBdnTt90QLGuSkx00GyYlSHD2iwQsBg+3kD1K
YyVCtwQd8zRE7kl+57ZxBUAtnvJXnEdyza2CxPc1SPEGT+6NQBFEMkRc59Dqo7y7
aU/9+3vV49WZ8hnQ1ln0z05PifZiuKk/uYwn1AIjkfy/KOubFksmVKlkalpuhSp5
qZvrp9lpsjFnxCJ0+SYj5zcHsZfYRa6ux84e+pRv4bNxG+9SAQp9iMkJrX1Kt9FY
RN4UxW0N68snpfGHSYJJA0niX5hTHOEaCVRnIZEdk9JyTNAELlEbGGXCLbClnUxK
8bukaKeyGV1YORENgWnzR8IWHhiyw6dase+ye7gOmuUVnUKPrA0sru8ck24gBV6S
0J8Nj971rydopQkgbGGG7GyhiJgtHYCQhxXVNMeFCZRWSC/G0gB/CFsPzX9kjYN+
DtuDEXABOdAsk87hM4IR0DkV0cMK5yrf3IiSnKY1FjowPUiD2az4YGDO0GfwRooa
CQyclUrYGnXZXvGm/i3dZ65X64Q5DxMtq+JB4I3KNoFsb1o2NgS17bbsgtPW+E2e
0HsJPgN5EQ5Ca+o9O2OI2xHabLm43Z1KDaZntLFOYYHieaYtyUVuk9UB2tw6omY1
7Co0iWCyDro5IK2avdBg4t+vFZNYLlNaN+JgnmvoZTeQ6CgoLnzzsDun3AjAe4EF
UjjqHEpl5987Vt6a2Q9FMcamgUFDtzdGUp/WLcktXczLx/qVIWw3+2NQVLjmzzhR
S+ZOn177vov85lEUKBjRMmb3lknqzmd+1ONpM06r4a3ztIECDt1hwJ7MBMapKOxO
+sMBktjONeTjLFbNzrG9R0OxjjRrvwI+52Yi88qJOxB+dJ6/f5xHHogYamFcZRp2
PKJzVTV8JrKCejKVAOT0VFEJmfjiD94i7Ufwoz8EBMfDb+e2JXC+YNjkOm4RBqEH
BU4cNUe5F9fp1Tce5AWO1c0SmL47L1Fg/2R22IBHRfhCNqi17aP/Cxluw24IaVGN
NmIi32pPjVQIlue6dhiO4aQhUiXOxDfQ0GaHRIuVBjLZHtEGTEmkQzLni1AX4sge
cnITqyM10cehSXgWiVHCPd6AkuCh2gwkyGdcWRyZ29ABT9xqb7ugQBxH8TV33unC
tHYS64Ds79Utl0ix7fTeKMlqvTrjMvGNrcwY8Oxalyt8gtI1mYuTmoJhBUY1GX0w
LBqZy92NM0+cu0tnfS15SjzKaKFOOPqrKwQrwMUDUqb9DFgv7WJ53GG4Yw7vbvtz
U+lMQBu8XTG0uxTUGlH7bimJHjidkCqwAd3eigqA/N6DeJlvvm7UXYgYC1niWiFr
VFBT3K8kOkyeA9Xgk2sUTB36e6Ms9I3+6Yb+8NV17HIl8DZ85uNIDLm6d8vEwGim
dvGLHRMPt9ZQPsmIh72uUmB88hxzmeq75YfouXImv1cMZcBn1usQGXPE6qNsRIhn
yTxLjGkbOFsxh4U2tpjj1hNYLO98hxftOUepb6sDmnFWDvRbZ2b1r1dxVXDgMSek
VSDsaUVgfqhKwIFRIaArLmQ/uf2n5SKiIClzBJWuat0kF0MQUPpDzUSC7Ng9tTyN
nKijVUIgET83eTXHXzjeJx9WKqieZ0REIoVpDMMelRN9aHx4TDhM/b8AGjSV+BLE
xlNYwT1+/VSAsef3auGz9eQS3BU7gdkch+vDI1PYJikpNfaXkPByAFaz7tH9irNc
80ksxy2mwT/5FTNcNW68nQKS9ZLGaJZsAAwTWlBSovPlRJipS+aDS9BO0EZaf2ls
Jf07a5zc6FmD/MppJXbefmvvBMC6/G+YUknPqHbU90N//RXeUK9N3G/sHvHdLpiL
L1ZUtt62YSK/X0+iKCz+kMNade48ovKDhrYOCBnTV/wSehlEDGxps3UT0uIKsgry
wkqHRYOp6sfShEIbBHp9fbBgxxMbGsIPr2FgXqclQlmm8g1DbLhc5EX9WGQToZhj
AV6UoFXcPQiAhJriH05C5Lf78YzMCaIcz3IurEdngDd8O2Uk3KmgIVJGG+8+GfTC
1az4N+wU06nzFytbPlef8T+SiX8V8VWfCzA4w/dGbBdg8Fkq17ke06NZENZI2IqD
5QHoFiyw/9R0Zxb7zY+Q4m1n0WTuCXmmaEIAuMm3wqG3nkob1J/H4bT/XB3uFmTE
dSgwJ5FZr8ADNcuAbYnNhBeprdkXwk2Yop2mSrGETnQOqn/y4cF4KYQN+JDHLq7L
J4Uc8w4Js4gpDfWP5Q44F0Zp+PuvljLjtg3yMrVmVXFh35SivdI798hwAYaObet/
D4T4CfuvbOs9geU074t4vdmQwLr/HhIFnGxHWKhFwf91OQJdlZtHE2TmxgoYsBQx
XV8yF7IVeOxpRPXgXTquSXMjePH5QsdnifB4XUOECzQ7BUV0a421lOGZHIU6XvMW
XiIfgLrP3lmI+T4m6hMpa/b7dl2LuzJ8RaO4EnJuYDcg8SnWxxfSTm8Z49eyRsxz
EacTsBurBnY6nNrjH1bEt9X4enNyUE6SK0oW1HjsOnAbKjwQRSMZ96k5igC2YlZ8
339R/cgLCOA6fRCEoPtmtGWEx4I9DtdHTGurlWsDBdh+7/x04b9pBfx0rgIJmHNR
p5RhSCIMZ1EqOmBmlBm9V+80vyZbe95iH41tsJUEdAMfFrZ2m8fpfxcmCiKI4tZb
KaEfnckEovLZBHhaKZMoNzwbkKWo8rwf+i0CMGb3QhOO5X3KiqB15+/2xFL+5mlr
p24fjqz050hAfAHsJTn+Iwu2OI5n6DJIRb0Fqi90FbSQUcW5PhPLweySdsx7IsV/
PkyUyHXVVccqBGVnKEMl0+LRfQteUsn3077HAmVpZdkLFNlaTmh5p2f/aR+vQAub
n1Gec+xs18uWUtVDd15iR9TVzAkqC+mXQv7MNN6PGjCmWVyKL0uzKYBfjE9jSN0D
5gIHJpcox6YBKPS5EAO8LMxzZAVEJVvuJQrfF+AJjymUncBmMRIqDKQpHr8Y7u66
gIQ7bf3uadxjFugUah8mzzte3YF2sz63nwDlftPS5oX+vYxeNfijJoego4GxP3Rw
+AV96eZERFuRc9nYn28EUNI2cEau0VzMn6cyn56fyMCWZ2uQjLcpi6YyGV7dZj7a
zc8EWJ/O619revXEdsowdNK1kjKX9bZ4sERKpkXREJyJUlO9a3P1z2OGdwbX8MJP
vzmVMZZS5jMwUjG3nHhUphxNAMFJfMFZE+IxaxyDH84hBhmtjFJU7n23BjM/Wxxp
b5QMo3mMEoIy5SqnKnCrq629FWj4TcvU/OPmKSfQnL6EPrcU3fgKh88uXP5M2B3f
/x1VIKmYz+Gtsl3TrKlbz7yPR4KCeaKZ1vRwYF+nGF3b+Ug1Ize3cYYwGpNFLcO6
hHBQjT+IeDDi55AHkhoTDwWVu5QRqh1iN1CorgGlNpbvEH5PruuC5QdSbqACeytz
CNbB4OljllqixCEsGIB3w+kPRXgarDULq2Hizn26Xj2tufk/ss2/tLmII5DsiLbQ
fT6oA43kQuN9dbMRpD2WqNiHfLtovMizTtNxT3+MvUDBJt46VKlluGY7aGL+/zAx
+idwbJHL9v5GNOJxsoLtQFNOb6KkpqYqPUDE7W0xx1eXEMHDmE3uSO1msQ99BOPc
VTdMDwopygLU+lrbyJHC9hTIw0ynxt/JMwBvVQSjeV8G49poACexencrdYFQc7ok
UkIA/JTvHbIywQF3ATRYJO0tQN2ghvNMhQglvSt9rQWfGdOSwmkwd3hF3kbmN1Dn
GzMBkOGD/KbRTiCWXP36xYAgPs6dMsJRDKohlPY+ebQoaikwfbUiSu6YVQx1ZL1n
JDnXTmf8BepIf6PKE98xudmlol9KAQwLNs2miHUudxR/Akxmll9jUL5Abhdup3CH
GD3qP1y84SAFGgk1/fq/c1vdMOxBzhgI2aZrrwc+x/OXFHQaxmCWctvjIPtVhxXW
zZrv65gEBuhdO9VEikHrTxLY0iusp28u9oza0DB26mHl7vCAevZ1pku0m7T/2I/b
g+0o1mOb42lHbZmX0PJojXQ5L8N8+V5s4WOkP5ZlVG9nGkCIriTfgrRbQIo4XlTg
CslC6U95nhH5VogLHF4kBZ3bFG0Pd5wX72Qktycpwu2OR/g9MEmevZEVkT2wDS/I
C1Jw3d1RmluQNNBGNRxgPogeHoo8MqIcMmjwf0egKF9o1kko/r09eiT+sBMChtVa
tggWwYAr68NSBInOoXktZ5tf/KxC99JGysJcUGVVVK7cz8LMtdiLgpxEGHkfBkH8
hcEbCaibQQYZx2C9KKKAk/MqhXquZ3Cnh913zzoZjhr878Ogd/bh9Q479khKBNt7
1k6ubKHLyDBY3GOCK+QbJZAko/LK7yYYtopjYy71id/zcrtUiYSF/MT1rE+3t7v0
hZT9UluNOclGQF9nc0daon75OwSrRgCL9VBbfm3cwUy5n7xYBqP+whniSKwEhR+u
bkGNVJcwGEdOu210StZ+c0v3y9y0SreT+QmIHq3hc5+rNXx3MJChx/UFObk8KuVi
DB6EECqFQcD4Vd9vpbrQghaNWMmckx4RaR0kV/FFy6K9CsrCOmjbiIAnqEGzLkHM
3duC9fNeWOn3r8H7GcOrQwf0Qik57s+63iQbCNanCHc5pTqGOzVSn+lIrRpjpmmb
M1bsl7NNjLQWdeI/UWes9h8u2zHDwQgfQEKSsCpTxpHtUleDc7dCBh+xg2o/A9k+
GQXgM4USvBrriQCXjo+Dt7fseVt8RHrKnA8Rqj0St0XXhFbLLol1Ac5Jam33EC6q
ecQqi25nlwBpXJS01WvODeh9NDxhk/XnLrEknotQ/Qjh6cUB0LbuxWBmDtUKSMrZ
ynnCnrcyj3sGlKRxiJWX69tJewzzQeBA6gUUmwlb9sjYBDwSW5lDX6yNwyrjB3OK
q6C7EOvcTlqf+w3yccYr26eoHk7ED9PMT3EYT7ZO+DQMArt5iDj+Y+Sbb1CdBY7t
4Icb2qF6c8HlKW7MBl151pa0j2/FaTa/0jaJIE/IHW4x+BcyPBL8hLj0d/Fwf1aB
QWTFSGZtiDLT2Dtk8UZlOTtxAZveTSeOtplygBptHD5a9+yGXlX9LGEek14OwtZv
YbqojYr0qlmrTLyEJmOXFmxO5GyygJ1cxNQ5O16zbNifRbarz5A0QH9Oos+acBYj
71WJ8t1LiVfYBJDlPkbJDjdYIvKZNq8xoHMpUDkIEAU7AoCHz4nPXC/T4U1NgQmp
G/PyO62+KCfl0oUQcaCgLcuZbQWm4mXS588mIRD5Bl2Su7brwHRw679VAErn0IZA
oxfPv3/iDbXGV3pwvmd/Mia6BheToflcuQmlupF7xdWERRzM7u+YawXf9xhk3utR
GMtTIy2yNHw9s7oPfAEV/AC+r5BJt9zAgjcN86rf+DhNaXdVdEIMkTLWbcbarpAa
U18kIbUQGHZrPjUDHCGJt3hWfh1mps3h5X4G+M8f4hy7g7qIPV1Zvn1Rhw0tKkN3
qQ7i35zpz9A02cMj/PelCIMKGb3OnYYiKwNJCiOJLmIbRD2AIv2UjnHGcw/n27Q6
2fXKPutNpc7ZHo7l+4Bkd5riQqzoKUtIJmZYiK9ckTxZ3rufZNqmbnAah/Qmitc7
OoBdBFeL2CrhzyNQGvZ/4Po0LW2hZ3DMF6Ti79R7mg6DaWTGuq+9Fmi1iW0o5ESz
BIesdGN8B3T3UKIfntUgaoryivtRgx1JMqNi+qizKKQi3lxRlyHuN1hWYQcK83mk
UBJ1rzYLb5klswGME5C3g1KKp49+onn4cAckXwA6yIQohOFu7cZnqZNp6Cig7Wwn
kOmVYDygdQvy2CFTJzqNwubhkhTOXLfqG6M2ItgdaXnixJWj/9hLxKQ0t52ByDVh
TuXVgkZn3NRkJRIBg8auzRRMRB+2MLgn0sAVlkMGElH7c9CGk3y8pEpbKTEt+AOP
O4bytOYHd4lT8dMF01AqGyzeYmkG4EXCwBZK1aDew7AACUFWx6y6vMKoW3+ln+gF
Xjosufy11LsvLbrnKjq0uDd83nyaGI0p/zG5NQSuF4LRfe07bMHMc89FY1lhPjnz
/PLUjiowaQ0pCAzoxWaN3RMvlYGFL0lmNvs5lnyWiw9cG5YkK3uqeXoVxAsKsdPx
012ma1dlZ3cQFopmKqhA3UKW5H21iEd2Le5XU3yrVv+9UPYBKN9sfG3DQ49ZyehV
t1skVt1cXdOUzlTYvYn5cF36RGEHjOf2Qi4oIjD/smd/ryR3kE9SYMdV132zH2YK
MoSY0bJG/hQp6sczWN8VDl2tZTJcm0NiE4Ue+UNQZ41basaF+PQSQAnkDuekO51v
xtDAfSidpqwDrSuEyUfVPAyq6seqL8VT+LLmCeCqOYsbkw5nrx5bRvsePjtQ4y8K
Izloim6eJaUcsiNAMYUspuSsk38Uuqpf43+MaoRR5RPsQm+UkqBg7bJanpqGudsa
k1hfEx0k08o0kp+UBLCt8iaDK0JcKKIXWCagRNkNgzTjAio/xleK+RjGvqRT9CYw
kXo3ztD10o0YN6cXbLsf0SQZgkBCT0JaR4wNUQE7ZdLHa4myJY15zNR79Kp5pWYG
A2Ztgt2eNaCSrXWVS4fw4Idx7Aq2pAaxbhA6R3XPxzS/UMq3TZoHkt1KvaDof+u8
zl7ScOO4MdmqJ59pKIqqSC4VzlSCfdY8tXUrFYNR+05Z65TKqufBCeTCaBQF38ug
eWkuYJ/q2m75FLWqf4GYLmDa4pK5S0va1msi4VglZOwmiVaFaP3ZXTDzxdzPPxOa
Qafzpp1lJ5EDDKPMdtGO9HSYtvDLSTgO9NrrWzR8k0BwpEZ67QsG3ni4KplaQZtj
GyjT7G+P8ZM+N5SaY98ivMe/+dxhPPTtbuKwyN5pAU9V7kIEjaYg6FLSCSmT187C
i64h/JS3tdFPVxLDOM28cT7utBsXbrx6ALJ+wOFPqlsVGR//+nSmtYt8U2pv/Oom
78QywhdJsiNbfBzsy2fUjOWziqEVY12HPW64HXlpA1iD86L+UJAnSMC+xD27BDH0
3ppoSMjokFatmDVs+LD1Foo4KVBQ9j1pQOm25ToSeaAer2SOuYj0125C19FzTijq
rhzrrsrAtXlOPPWn18zGi9zXuYjz5KTi7qojJzpJBNhbcmD6ezCl/TTyvaKeJS6y
+F79Nz/3zBt4MhQMRvG1YRwZhx/0XwDKDcrkSUO5ALhu6BIcVUOxlmHVS/hsI55H
x4gPDJmNXVifDTSjGmcCLcvL51gT29TkLN8CSZsBe2tOnce8xit+bFabofEYEWfV
NIZIX4mq4R/eCzqV4am2hMdPe+nV6xaXU2CoAHHiHxSk4kOks4phZYzCLl87p64D
P6O18ea5kMa6YN0kMgSNyWJFWcS2fgcsQZiAX+iMSRsEvx6XxVOpkhFW1kojRaaA
BKAd32/qybsNA+4bCJtTUsPyNKXcqAj5A1pVi6yXP2jkFzMqBWcwEZ+kxPqva+Se
nSLEKAhRTLvkQCd0kah2y34JPHyF01wsIGImoCzsjvo6f/7SGL/SQgDvEEYVPkos
Ut/f5TdbZtj1TJfYVPEvsp4h2nXBu3sAXDVjZEoEKshwlMqDKTD45CL5NzJRyRsn
OSRn84ztQtiKuC4IH709578Z2ymMD6tLBTcsOV3Tqf3bg2fFoDYzOi3XiwiEjquW
Iv2+ibs06NAtiEKeOpX99suGyiHYEQvErUqERd9mcTefS2rNRIUrdXPAhFLHUArO
gzI9wRwdaRE2AffPmFljDs7Y/3Vx8oHkS76B6CAB1dXASZUJqCZ9GkmJNqbAedVw
aJrsveKFJ+gHV9QKQ5bqRHJ8yXT0yOFsrKuoGHn9WORnJq7+IkjJLGb+OZwYPRVf
O0srYrAAXbUj4dDWcn3UUMTNWb0RPCJ0oQuI81gU5wksQhnfbD+OCXEZY9ISK3cb
OTbJ6jtADv8MN47kCwii72jVMlW8IceFJHwpdIz723N3HByYlCKUkortZvZ1fN/y
7XWEfagSBH0XquzAjcBm8DaFgH6IeGeWdtWJqp1HpuDnh5fuLPysa+CyLDBj8r6U
B1PCUm+zRGrfwfQzXlI8mJe3S6suEFVK3mfrPHTfm87A5PLLFrax3dKHCW743m/w
kDAT0OaJP+kLzMbl6XcxvxG+OFrTdSIYHYXCStjDMhRiH7RLVwXj2VtFBoWKbRG5
yuzYgVvJ57Oz5IDxfb/78DxwIf3ZKmo/S6mmPOADEGgFqHi659MBYo1/uSLzPOjQ
70tpWCpBZ/w6U0S0IS+wNXUkPWpoeWVBAAHCVjJpwa5rlkwlbqZZKeLoHQS6rKPd
obrzCPEUdNMuuayrIg74yp9kdlTOu+SA9VGfVQoOAc+pYCAoFLwGFxeq5BgDpjb9
5k/pz3LYfOz/NpSHSSSI7UAs5c6YDOQJETX6iMXM6j5cqYAppQ/0gSl23S6fnfom
+dj6Un1kSefoyDXCT5rGMKLzB+Qw2LcxHdGx90qhhfKuJkOW1bpQdpzuouaqCe88
CLuBqFyQ+NV1aPhcksS1ozcp71REBxVIlqgg3cK9W1Qh7ABWGEbIBVvG80ZpyRbY
5CthvdQKFoa41T88y9w4Dh9RO8FiY6jAUaNK+CXXHuvMuUJ0SlBqnTK87o6ZQ5eG
i0s42u+656N3/fdRvBHW9IZGzoq0+nFnn78b2oSkBUQYv1ATvegcT/kJUiYP7gJN
YORUY96Vof/ED+GoHnnjqSSipui9HLPm7wZYbjuFAe+ntcaxqN6pA8WR+Wmy7jjz
SOnMCAiqWmHTC0YUBFH27JbVNl/JnHl8uuEWx3Kjw9jp1IH4Aji281mI/WnNClxX
OXNwCf/a/JZLEqzyf2U/5Se6STAbvkQioqXPdzRnZimvrQvF6QAMWOMBE/2MI4TX
VDULX7FSB6xadF2rXwYB5UnKpiDVUOiW63D5HLwM7ZYlx4c7xVv3Y+y50tOAjkVu
7bqFisxs0yhwFqJfWGE45Yi+d2Jwbv6WRFq/H8nTyCfPB/t6iypD4awkUapJRe5P
yPLKXkzodWEBVYYGsvq27HaloSxSti6BeMezJEwAZwVPlDNTt0kJX3K6URYuBznt
Rsp/4jAJdmUHEruhz3rf59TONRge+f1NFRLYbYPh+KlvLRcY9wkrBErAdodnvaMo
m4FktsCODEG3+oTNOfi+qbsJU9M/njwnpoHBmkijYuV+MxljhFxPwQo4vmpW9uSG
5nu6xSP/SaV/37t/fcoHBEeEz4WdKcKpe5GihA4gMt4DOI6IoBlRRCOGthxT6wzz
fRPz+ohumvNOoqY4Aen5iwIMqI1z1bmG7Pup8KTua0U0KDT9m5pw9S0cvwWyWc8G
4bcPZDu4TVX/dfNGd/fb4/hKygUYMGCGTCepUnD6SRtpw/8AKuPykzeP8my/TeUM
88yffahQXFG8OY3QYzsT9/uAt6i1GZs9T8PMJiSR1YUI8ODMuJvMKfiRF/sfEhp+
2nEyvX96DHt46aEfmhRX039NVsbQNzonLShv5PxaPldP2A4Rs1wIMwZQNrey+agS
P7oZC6DhbKwZKV9gAGX49/zziRUcwpBJb6BRbYJgUEAtXVlmH7hrZNRin9wmsfxm
guMu1KltomUaGMtksgdBtkeod69+M198R6p+MNs9O57OyIaYMhS7bJF4d+bNW3F7
Xb5p0zHcwLvUVSYUeY1y5NDgKXj1jyOCOEIBbIAzMKpHbI7gn3aa3qVcrNJHgsuL
tfgn5OPRJ5hTOu7LLiqKAUEVRhesAO0BrlogH1Iw3MoZOZujqGr+r7ReNHsGkPmF
i2scFp2rv5+hHWvgFfNDRSofjRGMZIx0p2Q6dOgJQX3IrGePvbXfcfkGcptwEB68
LU/KYGcBxPPxQh7IA5Hb5WJl7xNdfFXXi8jLEuTOr+GG9gFMLZYVdmSJW5lSNirS
VdTnQCmcdGY+8Vlo41JJ2b7x4HkVStXd7TE9ABugPgUsFnPWIH4VVLgQF3+bcax9
JLzXDGzZhzDBtP0odkGZP2z4RqzcaPi9bE67WU112Yiz3nj0J9OJZ3XV2LsMs6+N
fbQym0R6teget6Pb1YEtOzpfe27bblvv8GimQmxyujX4vxrMeFt52nk0HCZC3Ajs
iRIZMnUOR3FJIFeiX5E97IEkbtBxVTnsbdK4eH801iVOUiawOpedV4TX1KoOnHIM
RjRvpVyybW6hacXipNpO5ykWNfYurP572nxeOt6KPt18jRoZIx42Kn8ek3kP7pgh
Hq86Q6UFqYnrvubkOd1Q3Zuu7vuxMM8HPx4zDU5+M68NyxcOhHrzn1DEppWS1vb4
Iy5xq6YNG9sJ4wqR9kdTsuPiptCYsKctILiu8Law85FTzS+7lhig8ijNtVX/2k7K
PP0oUMLF8Hm06RPdMaWmTFx5MbEePCTmmyAzZ8SXYR/drJQ+AVonvEMDctR4toJT
ZiKcpxbX5LOHTlov7OfjwTRibkfJWLZ5j36xqDMzh8G/Ne/KeLQgG29PYrmsqgBR
sjexBxhs1R+O7jles/XoKHlsV0FTJwDxUo+ya90u53Aos8Ntti7+QJ6nPkE8E2IV
pge0s8iw/zdrQRMXKDWGCaEwVejwr+4QLA7vRweFPQHM54np+CTONQmHeF0oBjMV
r+18jCLU4vlyTw5JEehhqBubFumGQpfj6A40ueCSOHdb/SoejCioqqy0a6sUnGCQ
E3FnmlK/HOY3Xy6IPr97/0sfU5bzY11bq5m/Xe7qrocMW5beJlVZ+4YzQxTeISXZ
Kj/7k4flvOPrRl/hdyR8b/L0RWYldCZQZsvPGhmFu1pqIdccB2XCiT+01b7xjPK+
seyVyUY8CGX0S2iUcSZcTtufTcbpvK3hr/VjGDFP73gfFb70HPLOph/JW1nnXC02
EWZ+yF+bbHE3lazNi+FIFyc4/ac9F2DSzQ9ZoUCLjRIX0hRk0AvgQZq86ICE74UM
OzGqGkLvsM/NtHl7BfExWz3QNxzWuOWGnK4OBsiSjI42H2aFwDnCFSdoMRYaqcLX
5XU0JGPFlPhE1lQRk6ILpF6/LVnAYWx+4jqNcz5yV0Fgc8/N+Nfw3/c2hZHFubMV
XF7uK6kPcZoV9ce/MP7Pq21qTvohak+BYqxYLRiLzQnj2O7AAkS5cel6NM/j59Xl
G9QyuODuHCaghV/YW8YvakLRshmTvrG9PpWsb8HAPZIqoH773rN2Rv7sj3S3yr/0
4MbHoxLYeJtLZ16rUNhnsr8APS0M+i2gcbew4j8WISoEnXfeIGyvLO+GMefKH549
eaefc58dKrjpEFoYlKZOAQ6WBnMeaI/vDuoE/x0VgB74KZCVnycfIptPjOdtzfgS
R+tDC4PveaOa0FxFdOij8WKtbmd5JAqpBL1J9aLux6aTX24muSvoiLD53WAGZhrY
PllhEoTMBoIQWLLkCbK1vdEys659t0KQdRQm+oHiUnWllNM9yj/v98+BqNDppCaF
/gcKHH4D91qUTwdFS9IivGhtYfO7ZloXeQnuZAtHnEACUz/FNKQi8z5wkxRW6v2H
5SLe6THQPcncP9Yi2mX0BrCOk65d0fJIRzUc+O86cZ89jkfj/Ma8U61oZg7zM4BU
4ewxwuWmKht4ZQdQzQvCtf0evL9+cObBjRFdSZXyN6a+ad+YJNcZCWTiAeBj7bBs
vCfz3JM+2qYVXFOxoYAezUglAg8/5WcPi56lEyGnBm+hjazHJ5fQCqOVEuheJ525
og4+0WdhWxgoRQFvmnsuhBm6EtIkfufVni3CBQHTidPJtAPJJtRG8LqQiOc3v2Va
m0H8I6p9mYwY1HN8UPBcBnqYUKW9yWp3I/i/AFDLZtqqmz3s73Ofz66096+SqFvd
ERwDcO1n9isYPg2e9KKdGZmhzWSOZR5NKvJqGpB8hLeVm7NHXm9IV6sZpDKLLJhM
NRrOGKGjh/reb93hfkAVzBQoetPv9S4rIb1hDQ07VgnRphFNxnrYoyCEqXRGOcm4
jU9dqdLD4k4s/QGV9tLlPNxlBb4A+KGUpwO0Ii/SI3KuCgIMdtrP8lGRNKf5HD2I
JEdHuu1JU7P+o3MZuKBqnFcADas1/E/YgHzzfd2saTmhGHWovx5wxGUG/ottya06
EOGdJqOX40GO6LjdXoNPxuoKUCxY9uKmLrXgL5G9LvvSPEtruRR6MhiiYE7FpB7V
PRTKJ64XNU94L54zGCBOtK/A2ucx+KqGdpD1Sza+IshAmMaQtaogYLZHmAxuQ1x4
8qkRff8lFnOTjhRMUlBrEvKD6K15Ap1lo3QgGDY/7ytoxWLEnA7HEeHG+FmQ+YSO
jlstRn28pM66t8CSZYRDD482w1D/rvnA5AVfwIUP9Q5E0DzcZokzOWtTMPz5wa+c
9XjT3blb/EUPylwcg9Llrx6d3jMpgv4wqlvPZWA1bpEHlFCMKG3KakJ3TO1i9E+n
i/Q1ZMhOnolWGiKvrMlE+jUXHLtqrMzdbRoTkG2W09BSs1t9X5BEv4toUU3PTUy6
RqBFa9K1RCXQSFZbZwo19R0nlzRKmWjwpNkbbHKqaXstFtLfv+JoH0fNHCltiTvN
96DXJf/lZLKfe0j4xLpiTgQADdjhTZkzNl7BN9tE45gCZAN2dqchvWFzLL1tnSmc
Qyh/q1GjTFFwnOn7SRxTQJ1OLdowgMaus9Qfn1XoYCNxVvvkzfPuW91+jDYHBn7F
OklY0ZbKMwWGKAnbYWz28rppP+v4QNTRuQtrchCrwYh6THjvHp2oGYnyqQJWugJB
YUEiEMdULK7t9CtWRzTgY8JHvxOOc6yDcZ9KMlZHDOMHAjaAmLSLTF0mzcTK1qxL
GxcWwgvxzL+XKHbMdzr9wNCE19zQ1wIz6SQn9wEnL7Wfv02OwdoIgZIsk0/zBY04
bg7Oqv0KedH5EbQnytbyk9kqMQqZW0v9oVqxe0W9IuEbP4HKyf+Ieh6WGWcgLbH8
lMp8OJEQOzbdCZnUFkd84d3d+FWV7e7eXKib34FMA9Q3i0jO8bx/BOLg5KjOBPER
xlrXY9nD+cwE3lzd5gq5SEqH4CjrKKN7md3B6RR14ohdv6x5up6N+KkFZA4yPR/d
7qvti0bQkITPEZIeEoIM51HFnFqLfNeuzmdIeDnbB1rgM6dG41S93bcLPbnd5Umy
Lt92+sE3lswhyIq2rKD2HNc3p5WXUHSpI18uDHYKU5+IqEbwHqWGcyB7CAFmhGv7
15xVbhm+lz+T/TCIkBq+gRNSbCq7hHj670gvQU1Rs2GtOcYa9YpkaSsWohD4ZUa1
aeMWkK0uADS10ZwgDhP9Fcp/OP7e7nLN+YJ770TTMA8A/CZyGjxcPoiPkHCZxmNo
6Fg48RQ115HRkYAmDH4i3imQnuADFGzzuqhfHl+cX+Djcpmo1GGJu807j2qMUTDM
jnUXrOtSpH+2uWo9Y4Zh0sUhwlmXawoVPLTfxGJPlxRy9QckULU8LcT6hrEwrLQ/
B30d5ptVrwluEZKN0ga0AeXB/9bAv5yEouxlhEFXipMf9a9HzjnazKMCzrDgZrmW
qbWP6VdtceEJ4nzTYp5eQX3IUksEnmMdGIJbhNzj/lhDYbfQEefcLr2ye8SsBM4i
sZoPZDWg3g0XCSOGpwWsp1Xx0aJVHQBYh5/yH8BKWaX/6fUR1ydSkKZnKETK31Ve
D2fzsy8URKh7Mo5IL5xsqG3jtXbHUdnlR4tI+xAhLTMTLFModz8DGxPUIp/D/8OC
R+wRqt3pXXfhdyp9YR31EgdOd1uyM90AV1tCxTUAyXSEg1SGFBwe5YGffOvetsET
wB4Djnlm7qlX9DpyJqnqi646I4f5/m0TSE16VcGFFFLLjDZbUatPOGMRXIu2/VkA
cRvGFWsRP12vi31sNYmaUxFhR3oMi6pUjT+Ha1hYFwwQAKhyiAYKEzZrgSCQgrmc
ZdJCZKTib7oovhjnEnRRyO6fPvcLfIBSBMstD+79n3ekmnuyfaV0ZxUqt32FAVQK
wCDT5ssS+thCr9l2Q1SljHvqbR+M6w1pYmIcUrxKYhxTdW/vaRFHE/HJDVt/c/eu
ga9ls1U6lmpxNfsRDm9EzFczaKwm95PlI2/4LFW8er+4KdFySZRqQ1Gkyj2Skdpq
4eGeFlr9/Zwii/eIGLoN/qUo9wAeUf8vBA3rxxTjTKNvVk+tLLubf6b8styykikc
/MRUmSZVAmJSqZzV7i2/ys1+z8IZHcxPuUsvja2EAgKgTKtFJdw+2OsIv6FL+Tk2
BBFhNXu1WouLKGLlPzSNgyeyF1vvR86CWtHIaXc0FQnOVc/1zSDiidus4RYH3i1y
FJdZ2hCYVP68PNFtRW92yU79wLltAEglvdu/WDXm5R9LkHRa13NEC5nUDq6gZTNd
21cNH5IP8iWrUX5SK322GAJJFT90lU4XbOTS/rFb/zbHbhulO0d6ScSTaf+ng6qE
tRMkRRSmH+5R+z+hsbzmIMxZ3nJE9GKQv8/wsHUW5tC3Al6pPES/S2Yqf3K5i/ms
8CyFV7vVvjn5vTCdmT5xr5T21rND0BbLAbMWAmY1fPQFTJvL+i5XwjersRVxNrwf
RbQSNU9QsNO2f0XJ4LC8xPv5754A6HhIPZa0FAFc3zSF7Pogr9Xy+8U6QQNWde8C
xSrmTMqJW4xN/Cj+ijhj3VliM38VlBo7+89AJfvt1uMUsnbc84/daBuGdTJgMjD5
Wzr79/LE/cCYAIeZmHkSZJ7CxYEvDF/K9tlNMj8xdzNMuDpH9bJaxsgpUXSjNo3y
lj6+j+P148rMuUnq3u7nAMsJFeBlJOPZCZ7DdozAnxdbASu2zScM0vkIx5qLMJBE
9qnxGM7VOsCmujusL/R+pXE9OCezT6lkhjoFyuS2AYfDTx81tr31B2RBxb3LD2L0
qPU6sMLNFKjwoWQcQe0i5CB0onVip4L+RIKUjn9kRbAMDj5CsDAM2KQlLtePkKHY
FHQehXEiX3q/wlsyBI336Nt5gxrMoCF1OHJ/327lPsnARkqYodM0MAeOoKBUzXME
7ErjiIaTUjzeQdcM6WXPUlOv/X61egL5+P4K4Nq9bdMdj2OXNcvDhhHwUj/KBPgj
hqdkCsBlhpbt83A7j8FEfxz/njyhKeuvwE0LY2/A6De3NhaH2MnbnmPBM8+0+QJZ
kBZkQDIqEzsoUxDZlS3nWlgyhc3E/IFeKaZgf7tHp/n/OBdbKN852v8udIEOnF+c
IUDI0cnFwJ91btMBGGsGT2GBxOcl06lD/AX0KGhx3W2trCVUm4HJL25D/jtc6nVV
oz2yYURDYvTmmIFB1jx9PcnSP2e589G9smdHWSvNUDc16z6EpJwRHbRnpmnDDmUI
Www2Wx8IAKrY22YslQx5HRy90XwtKYQIoPqJRJTaN8RL4vhpAYdLWD5SH4np7w1c
NWjQBtAUkQE94HDn+Kzzlr3duuLPChzMU7fT7LkI9sex/Ka1dHBwKPZg1WgMZdk8
drPlNKX1bFpHatbMxSkX7T1XD5psUw33KauvPKfKSKNIrh2pcX10mCAZ7iQZVgK6
s9weQ7r8NCMKePjZXr5hLo/zCLDFmnqo6NkxqG67scu7OfcfM+p/KBLlNOJbJDQC
tp2yiF24MXjCmSC3q2IEEaJXXQ7Dt6VOvLHpO32KSjzk+5mIMRgZ9fwX/5oYdCuD
nqAW5gLpCbpBh4yI1jnedPXsDKSlqJmq60lbK/mcNoHwZk8N0YvOcG9MFhxxJvgc
jOvy1C9ov3yncr+/Zv/3ywUbF9O95KK6L9sb1kuaOHQsWqIcxyqU7nPVALhbTqXJ
vhR0GwndTuZHbCNnJikF9KlUU2W7sr/c8mIVou5GWRcItfAXjr/uxe6S+Fl0IopX
I78dWDJdrpdQu3epD8NRXyWqMs24s64FOOZoB8ljPrw48mwvFp8yTzOIl34LQKX4
bln+oHNXXAo4Wn6d22HKubeBVx4sFACxQ1BPBwoIBgR3gBYiPdvLIjxasjLK+Fvn
etxUYqLFacXxAxgXCSQNehjyL45w/ieZzPxuyXigLQgoR18SRjbc2zukilAHNQ5W
zyCVPKoXZ5oPDVZpQrOH2rHwfMIcMzrT8qeNny5A0W6QRWScTImic9i+I9983dSQ
VrZ49jP5zGVN9Ys3xc5DpKtnrQ2Fgk8ezk8t9xwpMXqa3xR9SgfHoCJN1Dq+FnA+
y9q1+u7yzPzfurBBYEFjzXSRcW1d4pm5pFZamMo9P3S+CeRpmTiU2n3cBY251/yT
+xO0UCSpZYAUueSMPBKzhJeyq5NITPHDaq9dI0Ap31lNjLOag6RWfDMqzMLN/XMu
HKh+HiIoSZNLydtg4K2A8B/n7seYKzoIZkWJnJDzBJMCG4jGCwneH/t9iPBUx86o
zjCvat5ZuZzLqblJvjpqck+rjsPo78QAJ5q/HiEAfVW2gPyNgzej8FV5jz+xLjsr
fouOufQ/LT1fszkfpugssT9kMK3eGLbtGiZWEi5hT1egkflEU2qRzy+WI5k/GbYE
81nDllv8x2VR+HH30T0RCzDUBBmYwmhBreM9XB1PwgNCrw8RpGxYWgv89VjOCufp
YK8aoNl5B5pGvB8rUK/6J0qFI+OQOk8Dh1YoPQwYEE3nc6mmouN6kvUQ4mOEXYTk
eJJhlVReV0Nuiuxw0RNTyg+jHwPM4euhd7ZrtkXiyqXmiQd8bp1VvDj7YqVTbcIt
tQ+9+zDKIqfUJx2a87Hpt/JKUcewzk9CbUw4KoUvtXrdl++sBkS+N3a1PWI6to3X
BdA6QRhX9NrHz9xgYZKdMY9e0/6hrbOIxwkVnc0v8MCc/9yI9aJmh5fachRE5jfG
AkdEWPLaSAHS9sw1KTwyPGJlpJQYOaSlYkUjGGi+NcWb2GTeLs41TujGxQ5bsf3X
+srFTu9lT0ACib4NhdwUf7LYJo3y/AuZc7LTeTtk3k80QDBiCeiYcn5gm9dTIsxH
W+3phAMQmwjFm8q/oO7DyBYoMnqAap69Kaxj/7RAevJDEraOGg3b33kELLUotSH2
w0WpnSoNfooHuYBVDL38iMPKpy/FnbQlDjce2r+t8WIJqDHK8upICHRlf9bkfbVN
27ReZIZXC2P/mbp9+vN7lMynzxZ7jJOVaMQ9ZKDvUVRdvCaQar9C1ub25Gotgb1H
Ix4OD8SVD65CfKUFG/SLYAEDCUVQljwSEnDdGmD3yi4UHnhckGiaDOiiz2iKI3sd
smGYF3ML2/w3tnYyi298vGqOzpDIR865hH8lO94xa2au4mHI3GjEPAXKtEC2py+Z
iMt924mSzC5jcEBdW63zO5ImBwmv9YboP0mJGKExDKJGbDRyqrpI95WJxzn8DQYf
E2Yb+RI8JRe2CqSptiZ5eLl2oWVbsjKuqAaA9PO4WXxaWwQTShVETW5kgrHFRp3w
VUGY5/+UXrJ/GubS550VdIO80srPtLEHrfvlv/bKLd+Het1gz3mA85o1dYBCjelH
BfJm2A9GnsY3uBR4DUGXA5NMoj0PKZqZzAhp29wbb6E/QmNLiGl888XTpTPqr3y4
RL+fKkyDPLU/NGfulvJMZk1BWgIv90E7WtXPEPezO59xxQWm1+0Yp/tuKVVtfiME
YTJegHXm/WSabdqzB8Oh9KuDxyGaTk4N+IQ63HpvxX3WDCrJdslAeRhfKBSauqmX
X6t2RM5MUIPe4wNFHbz8+lsfgbZYI/ipxa1y+yUWWY8ARt9SQslThGJMBonGNXjv
21PNf6/HQXOIUoof87f77GW9l/ZK2+xI/lLWDUpMALFPD5x+sXtJjVUoWgSUfbeu
9/yajE1W35wzcrhQESycKGTX+c6HDUHWTI8bSJVUEpM5gtytSFz1jX4VJ7qsiwhM
OGJPvO5mqynDxaUGxZO5TnB8CE1JSAl13sVdvMDrCbT8IrbG8b3s0wiq7MYtQb3q
BGBjCLxyzOvQ4UQmz7+M6gA3fG02p6dGpLGGIOMupkzQ/rOVsAWrsunM8WgnF70h
NaW51wJkbscoDpj4ocYjZ1bOhbBNpBCgtbXR1b++0MVBwo3WdNEj2t2Y07uVnE/b
ZuXZDBfzbpKmc8ppZTVsPjVhpfKir+KCDwvwrPqw5tCkMHAS+HreRrR9NdSOH9Wn
JMq6s/o1YqqW+rr2iWGWK7w+xFna0gWHfpQz7TDjZAXS2V9nvvNXshHpc6VDp8wN
Y9GGCdl+1gEasUJ1p9FAnB5StG/2P7nbQ+sMfC8nGoihvIYVM7upBMHEVvZWNs6s
JuMA2e1Fdh/KRaJ+vBPwo1mVMBJYbczisrxHpmNZwgQbWynsq5o/eU0qtoLWFIAl
dOsTW92Hh2F9uezLC2n0+JgJYrqTMdrlWcwJWqc0DPGCQMx8m2gru+2jIgi5HYcM
yMCom7eAjboM/FDO8c8wOcKsVcAXT5xku+LpH97FRnzgV7/Kh+lTKwkqlSKUVfQG
0rlRXsIDj8929aJa3FQYyv1cpEmVUS065MBSNu/FlYU0SAmq7UBytWNvgLoZ6dbF
jqom6W97PKedBD9WFt9xYxavqIkTzcWs6oY0HD8CVYzbhlj0WjNn2aVUi6hz5TTr
IRFgPcpSjNMu949p2Lk81r4VlRv66qPRfUdrGkyLunHmrr0WUCZXCIyQ/42h/tgr
Jz9deQkXCexJmqWG5tO3GHy3ArtgxnvYiuPLP9h8dkKU3OUIfLOiENh02ZzgGL3l
9h3RfOdE3dWSTouk9wg8YOnSU/cEluHQ2B19Iz/frPt5QOtpNQy60FpZxmke6/tZ
2warfVOulP3+IVX66L64xiBfWzW9HCOsbxcgxhmsBy4kZMvDd1awxCoo6E31WsRV
8EGKVX+FD6wbymTJ56m94BdbVh3bwqFKXkKxDm8LtWf/UgTGzpGgoVm4MeiJpvH8
DooQsim1Q5G9SHYq7mkV4WKwN2cjZKwzDU+TB5LILLRrom0WpDN4NeCpITM6HUXp
kT9m/QnI9EzHviOAnWCjQZCLqUe5B1l1t2o47pSMHDsykKgwP+V0wmqrf16DZwbA
zfaBVssTrh66OXL+eLxhE67hpv7uaQNd5DIQj/I2n+Eg5t7wDNEd+9xg5nGu7Uj6
z2rg69q4WGHgS1dMHHQ9mPb73IMyzQqiCc5vzhXeNHH5NTsJ7y3zpCHNMsNqHiQ5
O4ou5agX/OlPUMANDEzqmxOGN0aUFGqd6u+uKgFfCHl4iKc+13VOpy54KMUoMAGq
NKQVEg5BnD5R+UM+rn5ZGgQDOr1o3Cbvp1C+oBhW+NrmVv8fI6Kau3ffr1Smaqcy
c3il3msWuwLGCZdFg7SfrdIDSnMTSsPjje3nqDPdjeNEYv/7i5lTDA6YtH5/0U+0
lewDZQL0VqSgBfzyLci2vjc66WWdUIoUxH8UQzVH31Ot+zC71tilexBrqYa2Bs3w
wIE6QU0yhlMj0Xur02DbtlJL3Xm84Sp6//t9QzfhljMiBIRCfXr36rPvMlc8dI5n
NQ6L+e8gZO0wtiEhrpRJtpWAGjtFZsgrJ4Pt03JkKTfBfxI/9apjDAEG7cfSoVHb
RqdS5QwzNnZJ9hP+tMfebo+vOuJuwVayekAYXh6+LkknR6T3iiGlwxI+PbtpMKBl
Yw+3m3hI8lbJ2VgXPuZNN42/nZHVzZlw3gdW1yJlkuma1A+EfekKitV7dBEBpdXt
AX/DLNpELGcYJrti8vfr9pWmfKstmVuDizqCp5OCBG47M55/SI5v95mP/wltuhzR
vnAMIZTZcUR0o7aTtucYFnWt/JnHu4wyPklPMFaDDdGUSWfCH2+0XRckNzquQwlZ
kLgYKtSFnmhz5Rm4gCbE/TzGcPS0TTMrmCv8gsTZWVWBDrf3J12KqUNaXUtSalq/
hWLHzmX0ZLz0dW9IIJvxqis/P5ys2hfQjTOgwywQK8mzwRFHzRBlUqxj2e8G7ny4
KroZJW+F0/Xq6aOTtO4u5H4Avc22AqTRc1XzCOrY335UV53znxae/nHNB5Ft3Imf
Z2iwYIsu23EJ0M0y66EN/+iBxqhmSycPkfcDqt7323MiZEaeSUesdBuPRYUOWcnN
5tbOp0S//95q6joeAlaUch2SvmeYoYgltjk3kdGWeuE0db+cCM2MTgCQVeD8z5Vw
+WKK4vb9MZvFiD21cnyeHK8OoOyW9TZvqnhMN0jEETf7oiCeHVdTfMcJ9SQcOYIa
SDbPZQb6WYzC4DlKB2ebhsKLImUmc+n+Z21lkwCdASuoD5idR7kHnk2usfc7VQoV
WeUX2iOBL6YQokRvfxhU5Et3xfkmvItLerrSNriJ81dizt3fL25YewlZ2FnAuB/Z
Gngyg6pubRWnnmASIRSgVb4c1xp+AtaR6snYgpazod2M7QA94LZZEoNt9vf9bSg1
NMpcJwlui8OL+f+Y83muQB+vprhFGzjJZcUqOnRA58hRxn604LfCiTOiFzYKDTBG
jaELH5zXA9sF+9dma9ihE/a4zydAh7avE0ZiQSlz5pTNq4RPA1KoNAsWwAsG6Ada
SKK8UunbrJmeApblIq2GZtJVal3kRZrldYSlhN1fsLbOVuwgtCVpcROa6hF0Rct2
nTg4Ft/12fEXFh1OLZHN4S/qD0XBF2wL0yXwBiIBctiBqIiozktJQKthSX+n4qZQ
7bMmqx9EXAD4aSclKlirLMf6b6pipi1C+Qd1Uhouu16jwU5UqHSbNG91hwcHPuBt
1r+NfN7MNa75kcG0j+Tl9h1rMUuyOkzaTcWZk2EXtnhaO0B3Nc0yKrcAL/gF1jTX
d+F58XpbhpJrSbz9MIF09hFecidvbxbJ63tOM5NNTp8AcHQv3A4DvcmBAku0FJjG
B4zt2Y0CzXJn9npEjkY9P9L0CcQRRTSxorKH2YlMxhqk7xNtSVyFKPKWFAGB7NYK
KYKEKyttNTQHb5E3KHgwS5brCKFOAO9M56lLUq4KFjrS8PKg2os/Qha09PsCufDJ
MLxqpS3+tDBxeP5gtkJQASeISt7R4MWYwxzxS+nBAi75bwZjCSsFFm1EiAwGP5Zs
ipQ4/lL/9LHIWUB5gbPQ5yGh3Y7Qw3iPgETRBhiS2VZNwGqnfnh2LrMg7TsbJy30
iV0Y8DcmCDp6FuySVr/nulRQzY0B/O2ch9kyVI9DO6hj9nQx91zHfUDiod+/VqJ0
T4QWBDJVKXjEdAi2jJHTPmOPynv88LyhHNlAilQnNH28yfE22mWJiD0PmtqFFI99
2zkiFfXZGCd6opehPjo94vTXubtMAV2qiQjpC6Kcr3PKBVOzK4aHMc+n0sWZqJRq
0EfnWdygcUuEj0pioZwAeNxU334TC0flYmsVRa5YmErgv+FjpFo1jF/j974a4rgb
MI7rcoiM+4xFESUJPp8QmrAdsxBwWVLAWcMuH9OQiyjJD5VTL7xHI5KIn30O8FZS
wg+B35DQrEyQ4f92zRAXYr90rIdKXTs2CWvx+220r8Uk9T/Zj+1RWKPqP336ACFm
ermyPhUxGrY/BdzSeFpKjHSY5AtqzghWnHM7/lP11nXODOk8q/M00bnUkfkEidVu
MlzQyz/hEIIgmGGcmWYG7YeV/yDzXxmfRzMhN8z1nq/QnkQ7MFmyxtVKljD7MbHL
Ua2XJo2eGrmmVhQMZk01+sZb9YBP+IJboo3cWXMjmdbseCBcKiy5Un8LJGgWLr+m
3+1wZrgfxDTC2yAzJIw+qTWoSWHL7szDuK3Vrwn/RgunEMDGTcWOBIlFGL3G8mRs
ru4szx+cUjo0KOMjU4nMnThsUDN3rJUGzPYwJUVqGU5S3sZpvjCWAQL4+v09FS7A
6RJ9FDRv+jk/iv9Y6BGQ8rXx36J29cDZYrRqXVgCXh70B2Fo4ndSMgsntEgOn17X
kBoQz7Bap10dwV/bgmi2PelRakgh4XKkh86/nPDlQlWXrxfpZs/5xXrammE6tIaI
4U8unJ0KQ4w30x7+N35yuxkYc1QtX44XwA+zBlwgO9Zb0MBvWAvDngAeV0nPhKKf
gTacN9nV4UYHqviGNr1tXg4R85bt81I4nJGhVy/A1VPXHSFLZjYDpcZp2SmioR7J
3QftBKpzAxEMWJItyVrZwMjCaWncx+8l6CdpyIHNjev4qwWBSWe2WymvBLL+Y7Kv
YXcg+D2bLGAiFYVv7WEUFmYWZXsjYiSQrJNJaJXdeNhXEGW5X+Jue1VmD+4OZMN9
Gj/sLKhpMI6Q51PW/7bZPuSJMW7Ap0Zhj+LbNiumN17mYJvN4NIMRSJJyEoC+RjC
iy3+OWD7EUgSVkSUqf8ZM5cbRox20PmJyEI6vfUMIsl8+cDk8FPjmX0sBGSmtkF1
y9FlOGlwUH0scFT+aYFjJM9vdkgBKAoDBzWGWpWHhuazVQ2MLxEDW3ODcfhJxwvh
Gf2HI5w90Pn+G6Zp4X32gKmEHrA3XAEyby/eQdh7WYE5HqMndliRm22S8MJ6saq4
5s9k+exSVM3gFED8uy8pJew/vjbbo9xWCHZeplth/rMElkIFsperAe3e1O/noFr6
PLu0UFAk6VKrseqNZICzbhRf0/A5/JCmXVrOMXddR/iWJW6VRdterMLu0F+DhSxo
GZtLBS5WsR4kf3tCFFjBbjEAwFBu8WTvcAg5egQet0BLUzDSEpkmafOcTYz6JV33
yXMihmG7H5f4pIFSQoA0b5bsjUL6EFaDxFvRT71aOUYJB1Q6fpipbFgD1+g9cln5
sItu3+EF6yQdo41qGMfAlwDPX7L4pRbx+yqKyjPBHcOZ/C2XoZQ1kt+V7ltADwKs
eQUN6nmAHHmTMxTKk36nyRoX9ybwQXyBQVHcPHxWjODevzvxzKJx7zcWVEGLiLfH
cPLEmXi6Doom6UzI+dxuRdPVQAWyMemJfoDN5uKsJSze4QlFDXI/6cHwblB5qHMk
Y9LdEBwKYKwuczdYwRCIPLhufRPFAVtvgOI1UID7DOhqku6Msb21oAG8Z8XhCD1Z
vc8rMg4SUbf8AfxPUblw2ejY3vxnHkyYG0UqKzHwXhIRk1K0sRtT7O3eWi1uoa+w
cQZNRPZ6GOee14M7k7eLlTfhjCcRWR3nHi31hWLHWjLj4GQbr/vV8qgbix1zbVR/
N9/maCmIt5NB30OJu7aAdCR77cMAb5xRsVHfhcQEvPDYzAwDL0MMjN0nCUMDZ6FY
aYoNmk30VtjcnDmZi104w+4VyJNZ2FsuMKGxbNjj7knhHPvLoDlM3PbeSIy9F1e9
y0wM5vnhIdQgm7k0D/mK7zvfhrELTuvHmCTXtoIATcMbu0lfg40MfBrZfG+MdrIJ
6E2WQyg/HsLZMmK7YgK3fbWKWbswM32DUw+lbwDCJgoizMfmFiX3Furf/VeSh48Q
QKG7PNS5Na4M5f0h0uifE2pF+JFo/4e/3aiZZFzSjTf+0eZ7QxspQFx0GWWfG+wH
kXYDukqSk6+Q2Ulmc70La+b6TAXCnEQ+2UpaR/pGRP9SLlZWl5wBw0sKUN9uuloI
R/1r9vWSOITsicmrmN6Lq3qkyVjowObG196qVW0zxJKs/r9z1WE6uFfF5VaMhNFd
70g8cAoIQV2J4YeDay6+tfWn3jXE8wxb51vvj7TkezEp3QxGIcAsnc4VQi3ympid
m88WPChz3kSaOkU5VITAcehJf55Chsx2om1doIZfQCYGMzgMKhZOS8N7zLTQ9IP/
NqxPqGz0s4mXTK0GKxOd/EEOVswfuuD03Z5xbFgz6e0Qb5yGS0mEx/9yHnUlAi9n
wsUVH27p3Tv0p/7gYVhx3zdMxkBbCc5z4rrw6Hj6VrNmxFLqjrHTqBJ8RDNURTl+
D4Nylqd6P0ayVyU8O7+hQO1CrbE1UWB2aW6G9ULanr2fNU/QIyqTVbeDqi6YfrKA
cHAW1FfIwdS0g/mkHNV/0W88qQsZYwEeuhTn4lIQlcidSrWv+ZfnlRAfs8yKwEDW
4Rdlrhp8C632SmjWVZd42XSDRzR9bzSw7qsRvzKJ3ayG4d7z9rGmQgCT57cbvQ0P
xB7E2DxQoZd2dWyFuLNp/3EMGYTZyw1OoSZX9n/g6SVMg4G1M6rPkmOSu8IboNWz
20JDgVJ5lN7Mry1Q72WOzWjGmAtN8g8f4LF7QSEieXzfNeJ2Nxxb+SWZXoPSRWmf
K6v86z5yg/h3nsciJ8URMPcdQdsXoRj7MqsipTh03uei81YQexsAU+ImS2Q6DNXN
3QHrrO1fOKO1nOLOsiS2GGKSD02BPtTh4ksMiE1XLaNatqqZU2BGYCp7291LlraU
WIF8qNZegneAsPBWgePW4OWWAFT62gZzBxCECwtA10q4hL8GxfTj3AUcmYN1XdR8
uEb8nOl26mCGft3piVacPTZAaUZZeH59QZiXwtW924OWAwcL0cKxCpCbmtXk3e0s
PdV4jqWwIkgYzBoQbqnxQWjLJNpO6XiHxbLlFK2AY5+vkSOLORcMaGgkYk5896pb
u8SIzlJZTji5KZRcA+Ju9D4BBP4kxee3+Z03+w13PdGEpe7K5wOb8wiKq+azu/7J
VV0Ca4WvM+YFBwwSPY+Ea9eTHSWS88xI+OPZ1PJWIkwvepCbR62nWkTxzV9gaPOC
sYHgme3SG3ecy7ixV9QMyRe3G6cRPKcjfgzBY/3tU6sm8Z1gXuPYfgTvW9tCpYXI
fEIHlR8G7NdFMTeZR3gEkHDrbuYqXHWKVhSw2yJ2KgprNUFfN9oHaviBlj6Yhqgs
prwqJmjqn1+XEGmQyZN46QM9/qhNSSJ2BJBLL4p55R6kWZO14RBWxNPtAdgfUOx7
rgNLJuN+9WP3D3YVf0OM+B9UIYYyyN+uAsiBzmm4cIDDsDiahF/ByegAugxW8LYJ
E3FmliVuKpoDA24iESq4rlYZdUZfn+FaVjDhUyQRLTRbbZYaTcByZeDQ1WhfuiN9
Kz7OI2a2/gy2nU9p00YCh2KMQSDuRMp+o78C81aGtuFkvYHewlmk6qR7hVV8F1tI
HyqtyOhEnhZK7zsCLpHpQ/vb1yJVO6oaHgkDbU6EKFGYECYZh4JxpU3i9pZsIKiH
I3ovrqNA3gnbAfUWDCtXJDkMw23DIh0l9HMSNR2ZDrjhZo9ZbXEzqXRrQPb+O9e9
XJ3TZtdQu5FHX8W8HWoiACnw97t4PzWHpWmVFrdKqe+3x6jF2unalrwo4WivxNhr
GOGiKsuKe6XYAb/SKjSQZOnlJlccDMy1yjU9ZCGYASY6ZiyXqtpXx35XNCFGlC3G
vrONDiAat0Ppl+2eeHO6omcHhRh3og2uUN44sOG8zw13ZgFR6YM7QgRZvZ23N8Cz
LsMY0EF5XFT5FznTtZFrs4UKRJhVZLANgE/47VIzJGYh7UVrHkBzVBQ+2dRslo2U
J2UyYKqIHStCAT8D9g2AdztRIRTCeyjs2VOVRn9r/l/OBZuEbRv8zLPHaDcO0W5B
2W3kDzNOUzFKgPFcA7FGHb7i3NuKCPjb0faOhctD57KnwTquSMNAAGR2Ds8CMpiJ
uCZHaevn6Fo91ypzvYBW5w8MsyTHgJ7qSJPtDCyiQIIWzEjivY/up9C+GTYfhFRp
WJz1jp3XpAXEfy69kJvFAXDwl2HSb93igx/79qjdf0u1PunNOVelZB2gzUPtgXIW
pFINKR5wYhX+z/dA+L7oZ5XAafQEcalxgC8E4I2xxqiS96Xlyk2RZSt+DEkbpmou
tWShrOJ4hAEVfjzz7rNupwmGviZR2i2++KMnM2CGAgqR1xckqVWQMK9qqBv9YUGo
I3ex7rLP6jtspD1QBcJAUU5smjYcw4U62smfr0qZWcsQnNhtK12UtPer5bkiD+iG
r0YwsMQ7sD2u5ED9hFv/UCBT8L9sCTpgzqYflaO7l1UvH/ymJuZe+7Qf94ayDYIe
9JnIUHv9FuyyZrvuyzKUhHQzVGVR8NrF6mN1EdXPbgf6B/PxAA4GrKPJLQ7yFGWu
5saeLE8wAJVDsMC2eO4k7sOKyWZlvSNiaWnv0zbidw1iXXOy1H+PPIlpDPZszZDX
xBAqCWld4PUd4ghtNtIQJ/PSCDoPKRFUCnv1JlHL1MSglEEzDycAxV64ihcDGbY6
kf+gWnQDXouOfd66ABoZcR5ohvQjousomKFSDQm1DDfLVaPH0cj874rVvAkURzoC
ZyMu+SfADUQWeoRwxC4euqLo5774JjotT2oCAJt0VaaPAS/w1AJrAWul8izTo6WA
bLIO4txllZWwHbZp0rFF1WT1g0j0hC3ZR8RClrPUFbw1kPg8ErkLzywfBYoL8kUa
YDxFrG4l2vrc02vJIrZ8e2OLWyfUi7jBzuVvuKwrOAROUg4z2/rzOI4F/kE0r9/1
scaoi7GsgyVtsrh4cepvczdDqjEH8XyicTKOy+f9Wk2Xwu1vWRt5VqqypgPhf41i
UGa4VWpE/GeGHGHcjHAx9jO9b4vaTcVsAz/eOWNgRYJOcKDKg4KCxX+tydMiHorp
Kun/Csd9/+W2H5JTG8PJ2RyihfeK38Q8rmI/fRGs9iI2xTWhzO1H5mNd5nCUEVpd
pSBp+rzQnZZ/0/um7aJbR7CTJbKEuZosSOKvISlFRiDMBr2MbTVDF3/IMCiSY335
dPRLhauEEqW4guwO8O9HKxfX6rE1WjAB69NHz539cCPqHqeMXGDcKdRTYthVuiT0
0uLsebmC85O6TCEkPvBHIqwN1/+VfhvU08iOQI/SMEAj6QkC9KypvNBrZ4usnzMP
qopKiULPe1T47cFvuYH1/+z4Yt/Mt6KTR+KmxQZRyacUZVVDrO+/yXSkD1udJ4EY
RlyTnk8S0aX3x1LuBgekfDQ0L/J8BcI4rxRk01YjuDp1cjWlrCK29w2nnunnOzSD
LeRtGd9qgNp6ot57WyrmbyuNy+CF70IRgcnTiosS+qQcv5SSYSfjOHT/EQzcg+kM
8qCUGfopkmzXZfHVM8BIN2JecrFnAYL5OTt+h++Z5isRCQEpu4vwVsV3JLWj4uYY
2u5fLLotXwxPkghpGBGobE1eqQjTmT+p6KIXjDI3PLonhSj202iXphPbcJyFqtEi
kW3e98uNHptkPRQ0xgNY2e6fja9NqMuy4jjWVxdzcnAc8QsT9XxHOKHaiEEYFQWK
/u6EMoC7tIkSYwqIvMUoK51GsXn8PECL653Dgo73pMmY2rEVKsYw3pxsWi3ze1AY
8adMPdTsOI4X2fKazAAOY3vuWxcSyvtvgoKM7lv6qnGIm8wPMIJBnR76YkLywCOp
dMNloV0P0bAy9rks2ZB2uE8NerR8bCnJJrhYVHKjYcaZTd/2Hsw4wBqTJxg/qzqi
qPVcOV43bwdsgE1TdDpQvVfbIfhnbqSYcod1WpsmPZUFzsG/8cNRS+t5hjuaDg9B
EunrwGMNDWF4aIJ7I3fy5/pXUlEknGIGzDWoPmOZhAWyClUecxZX64I3a+Zsuawo
ofVRnB+pLO5ghEuOsTLZYpva9M3WzYvdAZrON20Ilr8Iw2abSZE2lA0JMC9IWbLE
KuGBqygZep+ESxT1ffGXvJlqPzUJmstmKMLh1kHDw3YTXed5ZduSI9+CWDfhh5x3
FAuMJ7MCj7FAFwLY1tdlLiJC1tczvS/2HkObZVDQiLHSgOl0Uo4cuuylgOCgg67M
DobDpqJsXCghTjcBPogD9OedcdeAN/YymaXpGBL1LQcOLj6NXglQpaqG4M/r+NRm
068WeUjEZ05M95fc4l3vciV8BO/1posfbnD0nj41KEsbGDBw1WHOuWapAofFuA8L
8uZUhVxkAAKBlWCbj1EtZ9Z8JQsRLyHKEnX2DgG4KuS125WSPQ6OUqZAv2Vp1wu0
5mr+Ruaw7mhCn03aKjxDNYJtm1b9sbdVWGzYX2U2Ii61vh5LCI0Ww/Bsl2G8bKoX
oeqN3TSE0Ote+yd6ebEEnEOZmuup3P6fFZnpoTu9uaSnKMGj5l44nakjVWzBWJGI
CW5BwK3+tMlTxiJGMSr9BaBqWkOSL7pseNo865y1YuuaA3CBsArjL4OPE/0yRn8p
lzB5HxdsJZHEoMNEuaQ6hO4GRnmv6e1iDMCT5t1hLuYigC0tSfXIxNtNle89GlYP
RDXOtx7U4NMJBw26Iw11ehNFg/VzfYLXCItYmgpaUcJbYOCbUvIOUkSJXFkS+/Ib
BEUGiBf9GcsnBHLtM5fKdkh6xNr6ovhNr5b5FV9A83BuKAtDlFRgMiJLngy6dsbH
qUbqXMn1msWvhHGokyxQrGOY1ymJzKocJ9nLQx3CApH2+SYsc27d0gcT1SXCIz0s
aRiGv1OpAPS4McNGs1velwsEmeiEGsfQaLZquvkzQexJhCY4To+neAMUpWlnBimi
RiJ96MjK/nbuog1tgd4x4VfCGoqsYDIOR+KDKgi0722q6o9KnmGAe9TGdc0/yxHR
FMD1pgzLAZSjotgoINoxLq+KaqqQfooEPHjI6OmkRrfG731qAK5awc5d4DJDm3XM
oVx+7qDKRHYA5CrqcSiakl68dfkkmerSsu9kQhZEZi4BcAr7vTDY1UopYfqN44Kg
KDeywUeQZ49fm27p6E0Gbm6cJdkzVcAWZlqrFZgygsSEVlQ/TFw649g1+JdSq/p/
X2sI/TdUBu/a/tyxiJG/b4cbGdIM/zXpIOd8bAiMuM7JoIZLF7bnJ2+hhNijIhUb
aFNuM9vNXhBdK9T9X1lR2MrHr44qPsp8m1BOQ1qyU9JVJe/7HYC7xnwqo65YKbgh
eWR/NC5MwGrRy9rBnBdK7HRiqggjCLNxb2h4Bxi82WHrjFd1eABHaqoUEDIOlSgH
PbGPdtMCjfbZJ/3uG+3bX1r0kNKs8pHGD2F2v4fUW17ZU0PRm4l+f6VjhJfz8u5/
OdP1AlHuZBn8POczF6wcWNDinY3AlDaL9k3i6b2I2E4PSX5RJsUMg6a4foGZvWc/
eqqLuN7oqAvCECcWY4pyE9USBJ5A/nMenc+klPMSqSYiK9Nrd4A1J4ZKnCumbQAS
PCKYo1stoI1Q2cL646e9dZZwcgN913mbq1eE17VfxAGPlaNtS0iKBwrSgiPpi/gk
kCT/P2isGy2NtCTZh8BxNoQWpjPEol5GuH9016Lub6IPnsTnKL63te0NMtZ4TWBv
T8LhIvttUDKPjnCakU3ucToOV7nqixB3i+2aceey1Bz1NdJ6p38B+CsFMFZCPwyx
pOLijBFnQlo4H3lbFiXaOwETaOTCNUyM56rbCauUuip4d3f7D+3B7VU7sC+Czygp
lqzA8ueVvm+lj5Ax3OUh6XAok14Z3uJraP7koswcEjb+Hm5BqtT4pob/f4OFQrUt
xxDy4vmIvXYY0+kmmgU6x1BkQbIZdfd3aazF0E6VSymcXUY5ikBEkxu+fKu81Epa
bHD14TY7pWv1IXYBlRIJgmlqWtC/zDhobIS4cI1QJN9g61UKbsPmcwjVyQp4gBK9
PUO9QIMVXimBNYQokvIfLI9dUnVQ2IFgfQmMGEPh71USLKpTvOot8xRzgx7mrLxm
tEuBDkSVhPw6022rz3y1qBpJym2dp4la6lbGufNAAAOoVbN67TgrRv9iVVOu4sH1
t3zfQKBWkIhm4zEtknrN52XXJ8JalSni4WhWZLtJYS+32Kqt115mavR9CDRx/Kf7
ZJpuw+Uk6ETKAWCBpzk2CqO2/ltnHY4MTiaBOssMbOj8Fpr+wOjMblnyZcanfR8O
O44+RwGk8f0/MFhwdJZd9//HciKuwx1/LFTBgTr4X2R89I8tNtZnEoLaBfNHYRVc
jAAh8KGHJpXUWzUhKzZP3HyfsjyY/yTPNonhUlarTBNYE4x4+k3RuG/NXfZOilph
f8qAa0Ijpuy735EL4/QiE0+cdUuSGIFBW1cC4jTFvK3QjLnOKgceXAVE5bCT2NPr
QsKokRoJ1x1zbdWkIQrQUEbo/NHO64pA4GZ2EIXwv/dq4+XPrv3ppuns3tg0Vq5l
UJblBEOq1VvpH2HhDAWOrGET1W56AtbS+chw6ciG3WE5mGYGTLNYkXZsnlP1HdFJ
FFKclo23HBxIiRjeJvcYn25TJmmjH+zdohPebAHkZAXy1TKrgMilmAdq1X897ZT/
lT/e8JmjEIg5A/d9rRfpkOpGnqFkLByooHFcOkJc13f7tCsj5dI57hAyRNrL9iCE
VJ1Kld0Ib56U9u0WIA/TuHrgSX2g4TJ+SYmonZteO/l1yyFG0SVYWLcXdLjPuI1g
sEZdIRPf1kixjFz0CYxfusbvDyTW53I6yNPGoo9TjD5D8Q947wQ7Dk+7qVdWNsJk
C1hfyZ+exr5yTP5Me6UMiSjkHZzJAvJf/0Zv2Y7UdVloibtXSqurcRpmHVDUrZdB
HwVGRRmCJyLRogsn8ixd3oqrMKSi2mUFmFzsXahMbht40biEsPVnOTABPMjwNPzW
87S+mWEykPsS1uAaIs1NcFnI+MgHPLwmzNausq6hbrzj16V4l3MIL3prPXpLfEaa
7OR3DLiQmwSoPRomqNmK/5BbPeEafFsXlNfCRQc7c2+tcbf16bt1W3gw2Jd/SBO1
h15ECRSXBRUdcKYo3gaQnHu86wf+9Xxf6U8B0ePNRUlk/nmpuUFl5hlihLn7juUK
ggGgEXzTetjzsqhRtenJQAL0GeC7/TOsiT/ho/ynSgcvo4x7T4oXVCDw3ewpd6E+
sHEYhQ7L3b/KftBCAspOPrnY9O4SFIv0Q8zEKV+12luqTUPsRf8qeBM4dOiWEyKg
XZfBV0K7hLl9Iyo0wKMNH95JQE9ctlFlCIYM7lxI71enwftCYrnQCHWctyPBmlTT
LIq1WDULCxkgOSiLVeT+vSRScdAEZh36MwC7H7xiuINU/D2Eb2vIaDNR5FwFrLUK
vTf11DoYZKrGJX1ZuOv9RcUAZ/ipMSmdsSCc+80Eaat37V9FUD/z8oKH/tko9G/k
mMrrWDBFePZDd6oMAzpgitRo26/ExTohp0V43gk90B1kIG2c8T/BwJaR09EyciQs
E84bHx9YsA0HEkLUXbM+rCPf/0fdVimPtX530NOxsUNbfdow7qVgGGWDtKJhDbNs
FDM7hw+iI2hYQ4uW+8LlsCNfMFU7u5zIBcy5lkOwPqc2D3E0wnjfFukaRjAaSWNF
Sqvyr2iVdni7qK+eOJa04dhZeH66KxILdYtVdidoH43pauLvocdjoA5AsfnKUtL4
AA4o1jMgRWnyFmQV5yVzW7lW/fqdYNuyRpHcUlNmCTnsah6vNRhGuNey3c8styQe
KWG0nzFk8YJtdtjQ9U2gTxQvNeVu9wBHf1hpPEk8u4pJ/6jDuTQqZlTtkIuEZDfv
qQt6xiPmKX5oJU0CDU3dd6J/Vgj8CJ+qbDfUfqZRViXseGK5HTEdtBPCS325K95w
Iyh7vfb9ANgTjPMUiWTGIUosXl9T6h0WcMJb2E0VAQW3Qwsff2XIUUO5aop3hkGP
7L8WhJg+pVv1aEmBNatFF2VogEQN7BPOo2c3Abv0tA/8FM7qAqxQMo2j9KcdYNFW
l7UIUPuE0IMiZoV6dOB7pqjfR+yNilCsjHduof20BYKNouuRW8MgZD+TOtraDdM6
TnnWutDNiZuhFmpegEE24o9fYq4LZnNxucAM9FZ4+1dH6HEYc1L7VK18HKGrt650
LmGizYAKn1W8f5/vuAH6rwLtkGttbuqC5dRWF3iUoeMlpqRRaA0yLPu04tLxrtv0
0Y8FIFBuHbAcxfjlDWbKEi6UsjaKdQ6s9NbrpxBgOJprxNdi3X/k0jl3ZNiZg3Lu
WpA4I03VmHXn3rDOwfcnlkDCcH2851e4ij/Ckbrdkdgpl2jUAyosH0w285AA0z7w
XLqxMOD+iaZxtcDsrbPef1cnn0cP8JGu3QLENFwoSQT4BPLthAF/+zLbCzqOQYMq
6vE/Xy4PwnpcIOS0cGup2Np7kLhXAqCuAVmxtY2eGiZHrQ8TEBRsSIEYJXqfpF4V
j4Dbp8fNpYIdmZqaeG7a5Jz5kiwogk8kC1jMuy/0yGq0dHus+MWeLby+xtoiHUq1
Sp1p8eJtZMiqyXGb0bITc/SFXzpQLM4vxAtH6P4is9+eMcdDLu2bI2UmHoU1bC6Z
n8a4aDdc8DG0o0oX/hpeGLVJf/kTSTZwRHwFTpDa+8BuMoR0AFxuDksA0p7NgXfr
K3qOMTnrwVHS6Bsq/+neXoeqrv4zeTOCs4u8N8AMfdhjGZaOBhWaCCWGBxEsySz6
StUKraDNR2/LJliBP5v1ZaG277DDY19prISUQTsKqqnMrDnOA1XfNcrj5pr4bw25
wJFdpHhHTp7SrqfBZo41nIbB8Y/cls3n0df225bFv+pHayqo3GKMqx0/doKAev2D
s88rC+fPe3TSB0TeZzJrvjATl/HCt8fF5U8lmxNZfjDKZk4iNQAFD7rpz+aEKNgH
i145KZS3BlzQk61urflkPhL8IYCz40jVDovah6rdiUurhj5wL/wVq/8vL6SMGC4A
Uv/Vk5OTMjYYA8sA7pbSw381A8TEC2d7e+qqEGe17F7sq5VxeIzZh1B7jbUR8aYV
chbntC6remFqr//oCdn8nhQ3+eHBmyy7bmDPhtPUG0p//IxwaIOhj3REDBahU7jO
0I8yO6L+OYUT5B7Z3A5zA/TOEJSuLAIv6IB6aAuvDYK37jhqy/BETp79ZnuIDrbu
hjGcrTCFSRyYqH67mpbDfQhSrjUVDLEjd/cWX1FTg4+qG9tfrrvqx7E6BgRQ7O+B
Hl9H9Wgf2UVjew5KxuR/K+rX6EG9f+zF12SOCsSoej33Ei66FXj4y0tP/ZI2mPZA
cuMtgNVQUZmkvdM0EHd9TLFRAHnakRU7dnjRDroQvaxp8b7/eJtNTuMKO/92/jOX
RxJSTSnclHTPN+WnLoxIxTHOYT2DQwKWFi7Hvu7yePnfzMuuvbb1L3KARTZLHwa+
hfjHs9i08qXnK+NBSn4U3USdx2wPDtHFTTG1i11gsjhtNa/ChJjTzCkidJsMwg70
9LFM6xn3BAgfHGmUlY6LwdF+o4VRv4WCYN8CNgkP+1R3n3a037xSYhyFAXW90rZ1
yb5cdvqZfzIpk4V/KTlYvcvM1xjKpOQPL/TsQapmCbxidUP7c0g2hXpqZE6CNxdd
fxKFSyqDfeoKYWgXvt9UN7mWM5d2SAvE3+JY/xeW7RO5S7u/b8eHH0+aUbmpRbtf
JisgFxMYqQ3EwpVD0SJq84wFaWn9ZBodfbg/toO9Xbg3nbVjCaXW9NJwqLNtoc/d
ru55svLPhhYsDDFRg1iMXMDUQlKRwVsuAcEkWntu53p/zw7wgxRxdBGD1bTaDzpb
Hh+SIy0i0rK3XbuDQCDPVEY7+AmyV+jdSsRtXt1xnXwFAHlmFoRczZMzEHSGH6Q5
FlUcp9VaeLeqIVqI/2QUZzNcBqOzko+KkR1a6htF+SFrBbI8ZLlEWh8ULpaMS0Db
3LAkxH9CSuhCGCY/8O//0gFoW2l70j5yv7LSa/ms7gvKNWI16UENJVb4O1uR3/hW
Vq2gnDcSZkQsY0Eq5DbsuQU0KPLEqxoyo+O2HH3P8Ktlfpk0w5dNmofcmehdwqA3
4L3x9gsVudIdZvkfDwbrtMMUwc4HFSCBc1FcFOqjv/jOntoO1WZwuRfQ8L9RerX5
Oy84VfGJ5yHOBKug40XHjVT69ysjVURNJW+7U0tyfG+sH43NyMOWWxASOMSgyG5N
bypdvVIdfzQN0q19RfBPAnDNSAx9L/vhLh7BjNkw84xzNUoi7kp1WKJbiGsxQBWt
J+tPx5BCVv/rWFPt/thMhL0kbuYs5XHcXuJBvRmtqtGjbLwPmg+6Wfsvns/2ygcx
LaZxezJZaEL1EQyq+oH7TkMtLiLXdXjRpgW0EVr4eKh3n9fx0oYWbmlVDriTEcZD
+e+J96DunLWYUhY1r96D7lKWdWnX19jCdBep83pmSBaul3StJ+pyo8Oz+xCUYJ5a
vOqwCulhNUanOyT/0NvdFGXCxbOEH/cIKn73nqmQ6TxlG62tGpR4iUs5F258mQ68
XTOgBfCmmD+4CVL2kzgoj8FId2V0hdkFvB8opJzeDnW3EfvhAbiz7cWZuMCALpA8
6/Ar1l7jgbADucCA2uHpHR3C8/MvjsVblUBUNAlPgTNJ03GszqhwavR56CWqGPqy
6mgANyyjeJSX6WLP4f2wiLAmkPM3B6ba93vLGmC64JTqPnqgQInOzNOvFG0ao4n9
BGXzunzpopG3cJ7CflL6VsmOfSO9njOfer1/O8slJcnscARO18ofvRb+qMsmzKsB
0PeayEuM88QUy5hyT5xpSlIuoP1LEA9L1P+2mdEEnfV9DNmB6JA9tWYqJygLEsg+
h+R/XXiooYx0Gb44H0hRZKPgZ2QiMAmPiITW9sqqzl9P1PqYaw1mon9CA5GKYSIc
g8Q7SjKHyvtwilnugT/tMMLwd/J8v1UHXMoeFgdJMSxaDM3EXnMEwUFINvLdbulr
uU2GesKfLOspy7kZl1/97htRc801zt0ij56X/eRyJ2WuBJBv0nWOFOH6oOwLmME4
FcfsCSbLCLqdsy5OdaPvOTqvQtQa2eF0uvVutVnq4I/Cdg1O2jJ1zASjH1SdjpC1
dThWFY3rKSMOxu2hHqAPAzak4U2mDIqKPzWylIzaGOwJM7Wvpz7RMwIirZ6e/plq
fynVWuLkuhrnNYKS296HRElu9XnSuf3LS/9FRsh/VrMuTM476DBalEEpHst42WaT
RGPvkfVZjRzPdWU1hr1XQxMiDAiSCNyY8JD//0nOhHn3k7LL750pN9VfRxC9qjch
W10O07l1C/6JFZbsJfT3r7Y+zy6EDgz51JuXlNLrc23so4+jQtNJOPDJrvRQ6IpJ
iYJTpnDnXbWKxToaDoTsScmKQXJtVVCm6DZien21AJS/Sbd2HcQO05QAbDkuhIqx
BkwAKDx7yJZl45HBVDn87q/pRrgy8W5q0MrPPIwiUVogKj+Ce1Rd7lpFlbnUawzR
LuoSESfrFCaFQdE5XFXEmuX3YY4Q+AMFRh45NuUVQM7u5Ksn2TabQEIKz81vP3cA
qsezEnTpHP0aeGytjxVpJLO8xMD7H+BkJhE5ZJV/cWeeVDoKBQ2uVMXObcE7p8+T
DzSYTCJPx3t/keP4GRRBgFeDB1Eff8GHTuW/p1FMue5KA3nRmYn3/g1JrDsynakU
4UlJvpA4IPVISTLgClZL5ufkhAZWqE2/TRDfeDtqG7maYUm4EyQBCVqNC9jKLxqy
VoIDtoDQ0gZJUs5RAYe0JxgrJ4Krxn02K7Sq7YPFeppY2tuf8yOV8klOEJr+urSG
f+z6U5wNYv2+dKue0hNumMbVT7KS6D6WDz67tjXlwH80ROXNV74AkyfrJBrUwIYU
j5Me7/6evnzLxwJpkBcxe/gPTdsFXf4J3Pc0+DsvLPFFUCE0q7T5p/N+1M9zOPyp
enKr7SUf2QbZtVDz7MCkwkckavSCUeOGVIMZLSdhZRAnBmm748CzyVdkh/69hHrA
YIoSD9zoKieXmZX3Z8fD8hRJS1IJAS4cZG8PWv3rBnJqRKtWg3e9JaAi2uZv+deZ
ryEasrmXUF9M64jDb1BtsOkn2+NVWkJsb5EvL0IxrtGRBLGBWA/hOpkjwxAFBTSM
gC+YmuTGXYPAjWvdpxIfE8m7cuZ1lpMn/YrOhdj7ppuVraILauKgaI504x07sLDp
IXRUQ1Vn3WtB3N8WWeMc61s9/qWKI6mDutDxGy33LMPBOt3qydIr0lhExXDexKRc
c+kpa6yWi3XaZ4MnLvHd4hOnbq6LVAKJMhBLj75+gaJwepR9lXsQDo+jPhm//MEy
x4AqF+hF8jnM6xWJAS1C4XCMZs3/kTxHzwu5YEGHsUFGx1A0T4rv478ck4XtNh+V
7EW27Vn3fu0673KcAkjSZJogMN34zovVAljcvygoxxZxZrPUntUKzWwe/QzVFksS
m64QT39qTpRvV0u4zactXqLNlBhVNMSKjj5YEWlHCLrvUa3XpjOeMiX9w5fJ92uc
rXpbYnphiI1zAaxZ0X9ntXqjogWzI3VCcPxNLXpruYOdj5nhtD34flbCX2Fq/eaG
WXUfGRtSsEz4lAaHyLeI4Ok16yf+O5zSQ/oN+IbKjtybBTd4TXBs97gTAhOwz8CY
qHa3ols75khlEGgWTVemvDucTMSXLFi2pLtt2sznjfA93GArWVpFT9KepwvV/BCn
GcvsQi7IFNJ6fEpZindaz8BqoIbiMuqIdbJxbZqXSaWTlF+ILCz5bHXRriJRE0T3
9WeZqG8P7w3hG47QHeNDViVJm5OSY9ddkjSwQLqEcxS9hsU4vCa6PLWOCnoeu3bL
wzM9Ljw4zWmB3/IwNE1FMT3O/5QMQYzP9+Z912fDBddV0EZj1YS2xNGCUZGWPUEb
zsx0AofCX8oOQDo76v/W0B0ikK85qSLHAADpbfovXFGTjHY3ALyZs2wVnzGomGWV
ce4u6iiyHGLnkkFEJrgaWal9CLSnEKZrOPMS63h6etMex3+LmBYymXJ62+OYLA6z
BGuvk4DksgwZrcNU2GhRnQUcbbTrT/YszcogY7uZuTtKr0IkSeBQYnaLAkwvFR80
J3ltkxqjd/U6EoJLptr4VPaZ4O+5GzWq2eLKN3lzRLsFjvf8LkzWyNYv9SIapKGv
cJCFNos0Mxx9pg7b67OLkyiSUWGAw7FbJttAD/aXG03STvO/+9H/egAfsP4BdUoh
k2ybTxroBoFcd2lWSzVYH+VSJzue/yN/ZuQZUplzukpj+tH6x/2qMQXm29wBETdY
Ow1TzeCEXWmc+8QDNuJBW1EVhaoYkpImkSC+9136i0Z/+wWUUcYemx293/E8escY
uEwLLWFMsom6NqylRWWTHvce88ECgHXogbS1AxyEKNgjPM37YUqQbj/Q8nGak/TV
m5P5qP79RmVdaLnBaPn6nPBSk4d+3ZfpcqU1gTvdlpj7L44lxVxWlI+zyX20ifIg
MMGiTu5TFCJOBlJcomB4oeN8PFghmxvLwSWqR28eex2fdsZOuI5V8Op2fO9YCaKo
3FA4W2GlCHIxuF7R3bCbVNST9Ov1h70xQq2WP++QxKOWEgz42XgUWx2wFjEAjktK
OnnGRfuOwq28HNuoPRwD00bVYOG5Rx+rxFFZjnjmzs3wOO5iBdvgk8b1B3crmgbU
UglmN4GBCai8QBW7C4POFqTbK3dXEOqt5s4FQTgPOJqQsENpvh8Sl8vS94knvUng
a7NdMbPwmX3Ej2QnAS1hgZbPHgv+Oif6H2HVcHfcjGs1fcT5BvdMG95MByx6zvUc
BaUaHRiU1GjJJArAW3MpxXG0ZzZw/5VXD0fsWUadl6zK1LbPt76uTWp5eyg2FLbM
X6QiHS/DUPtmINrzooVo9ETloCUhw3HXBs4QmB2ybUIyMK2t5IiAYNnjFNr4wypk
b+YEGKxaYv9iZtQQhIcU1J6nJafH/sJRd+tf/Qq9+24SksVI61MR8Mxg4NmfdM6k
H0VXpbF1DRw1jpBL86kwoYH5xlUzjekTVKL2TeWUK+n9n9PwvEI6oJRmBb0e+7Jd
qiZBpX9xWTdEgIWBejCBTwcOQqXfu81su0OncNOm1KvPnHNPQtDeesg3sb9JxOr2
UFppS90keT36kEndh+0VroS+J+ENHO62p+99V2NjQVMXl2LMXrZtXt12/1B5jKrh
5gRSyU+oOks1fO104xa4FQr4B+CeEJaB8JNCNpY5zPotmeRFj8Oj7iX8q46Ry4V5
SL/Iqyj34cMXb2BdAooc40PzdMVnjEhlhcIB7cA+C0A0vr9UBW2k+ShQJuPrPsqR
6SX3DOwxpbD6ATRnEb07hS6q/EOQC0EY9GE1l24GJkgfIwDvR5L4kwsGgnr/SwBO
nEZbcHWPwPGLMddl8VfG9D/Ptv/BGwy73iXF4Y4pqYsuwNEGkZcoBBAIA/1yLpnf
uBl2Cf2S1TqxI5MkhdoCca37umJqmBQc6m5g7HLAhd4SeMGJipUyUr/o24GHNX4d
dFeI7UO0dR72M6Br67rhcN9Ump9qMo7ULrRcEyJcmKTi4krKlhyTCLZeQkdesCG1
1QZhpSxLaCWv9e/9pga49/XQpGvN2QfHpizZuG6UUY4A8nV+gVSPVFq+ZLs01yuT
FH1GvocPi0BI11UOH4HUNA0cMgTzC0DdvaW0USBhKxwGI9ERPkYVawfwVd3xQjAQ
5u6qZqnV859slXxDTTdNd4NUOOm0WgbzfyM6bH4n958Ij/clHjSaXa1pnR5rT/j7
1iVjki9Dst7i+y0PokmdJIVSwBfktrdL5spJ6MepSPgDMJqJ/1jXe4zGFt1Cg7gE
MxCdWDrWWMQ1CTdrZK5Txd3Zftf1aDkXes5JTvfeBdBVH1IZfw1GnRTPhLkJ0rv6
coIoZ47qhyExAN7v01clGKXYWsOWlPHuCb2+F9BXpUBNI0SnQrOcj2KHldfQ9E06
yGdQ+rAGx0sBx2ncPvf3m2XV2vXhr+7YSZbtIDvYNQ/IiitpU7eZKh6WjTLqSiTz
Cn1BpsZ4zblRmdzTXHo92NLDZ+pk6H38CWcTm6uQypYHdY2oddnIaStCEhIn0JHR
eT+qtfjA5Q/fJHGNB41Y6VcpKt2x+eonZ4WCZjeYCd65wQp4It48ERZQZBPN7O70
lSbbGRt9hwGKgM14Jj50aNBM19NvtBI9sNGtC00HjoefLkhtOOv5SkNiTSXkbb8K
RjZOTCEdW/6vujoI3GevTi35ceghFoTQed4rFgNIoEVM6bAqpEagffY2XAPahtwv
8O1DJvWuaOXXQ0Hl0nqA8mL0ueXhTcGbLcBB+DdrzZkzWDdQxolZUrt97tWimMvd
oMkXal7srfrQxRRVOVQfZsuVdDi1Bxz5ZdSX4zBvqajZojvNCihCdVoV1E5GUz6p
eOz2ZkQAOThlhHKFZneXelWG8Asc99+B16l5+/XQyA5+Awc+aAz/mt3ZO9hptspH
ixAaOHk5Pco+j2MjBwl57qbEDkkLKA8SqEWxq3veEpDL12ScEJSXUVSnnuGooTaB
+m+xkh+mYmocVRLc1cVCYMahRkFzk1wpsuDQqcccCEppgdQ7VeluVozz5+ikuBcD
x3NajFqLG/5KpMX5Q6OjhNNMmJOKMYAXpPRrWypss38WwLYLsOZdradX0Uqj8pcU
BKcLyFF0aJrtb0q8kbsD//IFTM6yLbsGpe3blBo8BtBBkhj9eYOFl/BE9Y1GG3FY
PHU//re2REaks7MqyYxRypNl6r69Xa2GPXv+DO1McVPaphpn1wB6D00EAs9EXnCq
ody6vyPRfYwoszdxm8owg8AGTfAOGR28V5TyvLSQIYkIM2EVlkkVSl8L2udGelTC
1HPwHuTHZ6f4QQZWDr/siQixEDrFivBN5qlKngzK8SawIZtfvTx0rBbDa01SFvBW
pn4AtJQGiehNnBa1pmYcj/nReSWccc54K/SGcIScWZIM6yk1h+BQpZco+N4FSFYg
BU5eag9st0Q+PvXLX9YoKc44vjJMcKilqn39NHSbe0msF4vnpellD2j67tXdNXug
uiVAV0TosfFkdzFgQhhhiz0qHdPzWCM2OaJ5Jk4H10ESslhw3R+vOxv9u2D++FhB
eeBs460veHjIkDB00ezjOzX+eycIEL0eFFLq1OVxrxQoIjpI1m+/xnhLuDFIO7Rg
JHEPZpyOO8SuyZIyVDJgUx2qF/lJINEV7rxxF83WiJ2B7PPB1XmYe4jEXP2ohLNz
4vfQ6qmAQMXjPzbd5fCu67vsRmwyRVMbGfXeN1hfpPu5+KWKO8ceBpBOW+vooIRm
8ui2jRa7JvEd4SCzovkwwbeMZSMhgvk/R5BvayoWgPnS7MAa2fwv6+A6k9Jtzdrq
GyzMj3yR0nFld+qLctO5dDbAO3kT5Sln83v7nO0ZmspLUd0ywcHj0clFy0lNZ5Kh
kc2vn1uDmPKBeFGG3DIE7ocA+WtpHdbZZ+ymht3SV7CTsDAxABcGNJ5pRfsrkF17
HMCsT44bhE10od97AX+Wp16zHlWUyq8GVs0EDDQuAWgimmi8GImqCFgN/sAhMW4H
b+UbY7eeGdcvf7vjlOu0SQ8QdYHGSjgmHWIp/qPYPj2wcGm6h7kAJmgfq/8Q6Y0P
kDmgqDqn9Nete1cHSKpqY3ZpVtis0M0AxLQNDKFAJ0Ri07OZc6UATdSZY3bUGqXe
G4CD09rI590HAvEEGH6pcgO+J0aM5NTGKCoLBeItws+LgSWV8VHATB0i4gW2YGf5
rY2ceCNeBlJpUCFYpUJNIqxhHCJv0A5HdIAKtFtyMINLjHfZs7nKCp1EJPKQI4hu
2hWdtQkD2S+wjyigrSwxzkV6JVi2xrS3f0Rv+KYgIiBtPXZ8DITbcpkOhZC8P//t
AHYCDyiMAYO9AvwM62XeXtH/oggm5a7KHjjt1SAJhfnGkmjpGXZ3Z9SpOv1Sl7My
dm1M2KmK25NnUFPGFsnU3c5vyq8EeRSiHuRLfdZQ3WGahVa4q7szuR3Xjf1EmSye
va9ic9RuFJIBVhKTIRDG18NJR+dkCWTK4d/elYyvaNUlmgJpcGTRVU/3k9/qrOon
XZFwQQN5ti/lMy0pbj0eAtNgnwWSWFsf0cT1gEUbr1HafxgkT+PTHdl05nHKMS0w
KFcm31Z49U9XNDHtXbA8ObRD+y9LozES5uPAbfpI5tKeWaLpzPSG1vmP/9gCsazK
bpsm6SFeIy5zpwFey1vZsc/oV2XuFle9EPcFBI/Dnos4o6H43ybFlBnLH/FnP1uo
hvSRl6dT0MYtHJZWs6Qf9rmVo1rqQQuCJXDSOdIZY+3DFsCEWJMXpsiFflhm9XGw
jdKK0SQuKbSZ+yKTUXPSN/X1V6MiXSeiIdV02S+U29IhI3IFcVdFcgT75QcBvX+C
mVA2eh+uCFymhoUFMJ+rNTPFEltT4UGm9Kj2RiiW9HvLpR4iuUZsnPCda91FYDA8
KMr6Mv44wv8zsNEZAmAy1WtO7lB8SWd8uTkVMmPzJnNuDVSVh5zYRVzZy/BWo4lX
68OCmR8mKstIJZTsH4YvNBWoMCcbYAu2TNoAjrZvlBqUK1wCTX6jEf26c+Pn9G5w
MgOFiPIJuNjmBfxlngTiyMO3G41CQNMuSW5EjQVHnREI9mJ9yGKu7LQpbf2Dw9OT
zUAJUkwsFxMKHgAN4OAVvjchbgq7C7+za4XABWcP2LYDgRsFhYkJiWKF2FLobu08
bwkcH9TEhzxyMZHr1g0S+ANwHEjUCOEEV38mCmcgtGhAn/pHcyeSHNp1+WntG+dT
z6M0XzWh/PJa5jDzh/8yh//SpVci1zuJG7cflVXhTKUlACZNf5LbmpSHYY2SPFpQ
iwphMFYS7xjJdVarRqAS24jNv5uAofixm7nngUB/OnNg4fLj/OggvFjvCugffMCx
Lppw+nrNtmwpLxSawTNP16+GSEXET4WGD0qUFOT8TfXvuM0TVHW33HuNUs6pm2ej
TIbPWb20Ngg/5udslLhvnKpNv67IlqlkwmRkr4XAHJhpdH78CEum6bL+DFd9XSnP
PjrnzPdBCzZEPIddq/nLNUA3spJJBF/Qg67hUDOuPIZYogXwKoKOqzqgkWEl53GN
JPHsP2/z9hqTBiHTZQ1CwcUg4K9wUtWFq4LuUL2WZvZFiElWGF8ANUsVtX0uGgbd
GEP1awqvGbj+CAcX8BHUGKM733vWPO4S+8vshrZZuGrHpDVUORpWplCYPGap9AS/
+WPRRY/bYkqj0tzbtTRxEqKdE4uTpexKpyeneb1/AAKx8fWDbUHDbVcw847MpDUt
oH/Jtp/a5p1M+SStTdNkr3WxFD2gAEElCA7bBYSmjPgxD6rcXsBzsMPxNn2pjcWY
jXs0iQFZIpNrJOmBBXJpE1AeyFsL2RLI57z3Z7mmCEBYLIByzetg449A3IUDi0CR
v/j8Y9qXggCuNzrEOwWV/8ia8GBUlpdK4tGf1JklbdQ/n7C/2c8uz3Nn6gdi4r/J
sfsZd/O7sJ3Vyy/Xs40+A0zAIPGAR6TYuBEUMZgGUP1Bs6TJZCr819fYL3qaL+jF
qlL+LGSytkwEbU6tI/+r7+pPQA0VAir749mAiAW/AN2xHimxaZ+1hyM+hxP4ZsCN
RtV2ux1s1luUcW01U/eU28RKfU7Gi/zVkZqDyRdMR2D1qIudVFke16SK+GOq30xP
B9rgzt1DrqLAqkFvGaF0wWl46kT4RYhXHx3p1NfEYWvfRofuFAM4TB+KhX8TARb1
meMChSAHZnZhacvoyNL3g7KqWxEOT2cqcP+wX0YQKgg0gc7WMVTdb89J/Q3v6kiH
kPpEnRYDp5t6cy2eCQWK+haoqd17e3tAZQ2tQ+iMadDYouEplwytdWbla7EvZ+JE
XAYwZdl6F1uTGig5Szjq+dXyvNinRM9E39amjRZpX7UN9JjMmulnxB3X2LP6mcBZ
IPHPzlN/HnWvCUqiNPiOOpw3CovCf+wx3lbekN+hSX3PA/wHhWZviFUXawfveGwt
3IuiJRTJvvIgDkL1pjnjZer00FEjiwUBc3CPDvX3Cca2v26VPteQIVhpcZWrhLQF
MtT6SLIN2OMuTeBGAllYjXhsApJ2rfNw84gXEE1rjAWcnQXgoO0Nbwhu4rT/oNDh
gkCS6HLsAWeqVJVa177jLhqLJyCKFUGErrTEMn4xXekHAN+J7KjTM5sj7Sl9QHjX
yj3PtMf5CTyKbcFzAFss84kB000SmEPlQQtkI20XtNxOKxORQcwcHQT66ZXBDPcK
o6I1pavO7jyCPTw6AS9AVNdMeqwPsAiw6eAij+Htvv92O3tfOaP7ZqBcvwq8An4k
RZOi3XW5Rp3wax35PFrDQKTBcWzRVFnEQKEDYHW+20+OfpKZXIWCzG4BhYaK0cda
FPnUCY7ZGlNlEJw3kW1QvVv1S0m0gTcWqVRWMIKVwNbldFasZ+cxdcnHiITladEn
3mlOFaeVbVdfb51jvh4/d3B9F5iBAs181p+N0DGbHbl067+kCwkvR9PvE6e0WQx8
7vBO+fPjUbMH9urmlfBYOkvWfRDr2yqA4tMWCjydWIoAN7pcU9kH61aNDe8/Wdvh
Hx4cN0Oo2Evew4+RiEIx77+F7ytvMNCKC2taIbJuIGeL6xzVtCsvz2G5aTB/hO3h
YHgV7gQ2QIVyprxW/O7ErEll8qxeKaj4jTF4fQMDuRJsrQuVi0eri4fvjSmnRquZ
S3SBuCihictTRXMdwFChAf2OD8A10W9GivqooDseEgE0sIMX8UH/tl4/YfetLaWF
1TKiyInSvdKXvoGXB9Nkum1ZgXGP19dpNczClthaDSsbABYq16/uPss2cKyFEKTa
QHs3ygxA5aHE0Tke3GYY1MYYx05waUK81vRprzKmADWRYpArCmMYdoSd9n2B/yeV
Wzm7Uq0eiF3snoV+ZZKvMePrruZ5fYZa9nlI6uESAH10vMEmuaUrgqG2scWlP8d7
v80Il0LRDNHDP2j2AeZUR75l4VCCSppLUBhfhHufwDLohfaKjCI9J8sRqFFurxqI
0ykjzW/Cptw8uzeT2XuSTXzjWtO7NDMHUvUy2M4SgxpsVldRq456aFuQ+vWopjKd
SGaa7uia4Dii4FXAPWjlpnJHMulu6g41MRHBwYxdpxqRtiRcPRXEH+3TWj3gtTVa
JzmNFQP0Vpmrfu/1uj1peVSksYujJC2BBn7UqqIdXzib/Oj36Hur8LZkOhjfPOPM
lSYEJ4EJvtA9GWpifwCCruNQ8nlJeYs8ekTtpWOHburGUuu4Zk11udrqLIAs3Cpp
IGkLdJs9kIbkLhXhqrUBxDHHZuN7o1fp9fVF2SZUK9PVFG6vCF4ZisYjvBTspj25
vZCnF2zX7jQ8fPMqhJ6p0BSwmgJ/uFGjICeq7wxqYzxEkOf7TdNQ+BSOivphf+sf
qg9B7mFxMPC2A7VrfdPbYTnSf0C3BoHkBPNqi00KARx7U2fgNL7WkZwpHFi3Wg+3
0YnH0IgCdX3m3LzfdxESHRjSPJcy8h+ZxGTNSrjANumyGqPBvOGa7voew/a5Qo4Q
kqAEUDfUQ6jg0BtR3lT+ZqIByDkXgJRJQpv4wOo5U+5JU/Xh/OArwFmss+4LcAFG
nMY9ug0eYBdSa3Sb3NKVUuKUgKgaPzud3FXLkG/itqLfvPlu4lcf63etCzz9kLnF
Dt1TsyoSjKJXdAg7vsCJ79/rHPOENZI7MUJEIgLg5ekn1PHo8iLZETWBbCrMbNPF
Db0j1UkOw2CwHWvoVOInQD0DUSfdEKjA37EE8WXafrdaUfgMnjUs2WD83cwWhrTZ
HeA4xys1JeblWnvv4nl3PtlFSYLVTc5FUoZnPhUtZbe8C4+bSkH9T8y8XwBO+uf4
uxFbBY+f2HVHkzZH0PzhNylnuFZwpVLHXXdPupi7wm4/l/5XbY7eSeyGpnNHd1U0
TGrbf7hxxvhDZ+5OC5UAleolHm7ESCcZJnTvKQA/I2eiz8cGas4ymPrRA+sQzt8Y
LPW8fMVjUTs/kpfcbDD3BIpJxOMcFqjfJuXSWZUVbEsn2LGxIq4MtSRVaiP5dYz0
V8FBBjJM3+aVSA2dh8wNhJ13/gmeSuhok5+gCBHTSpvxUPAzpesF0fAj6qoJFQmt
5M7WhDkelYopF/YbEm+A39VvShbTfQuY4wLz60H/hmMtjQI8sIi3nxibpeucSPDh
2NsOInZMaHthO7EtpGucOmQIIXvtDYcSnO4ETNfg/rsQcK/YBE4ZSSzOF4hOHfms
5YgCbP7rEqjuBVqNTYzXBN+xPisbHN7jrwgZjjenmxpKIQEPh6ntrQOnBIa3AL8M
bqF9UOIy4WlXibFsMpp4ucDrP4jj2mP0HGIzsRXxrpJswYZUYj3ipK1u4kOGuA/u
nT5nsvqd5Cg2joxND78QsnjwQT4YccRyDMXW6nmy3FodgJltUObfCtpZtoGh7iv/
Es6aN/9B9OC4u6cotKHFd2ZAL8Dfvk8im84INPUU/VzNvqQuvmo/A+GwqRpHEQ7C
9fh/3J6d/p3sWFzcAzcOCH1RiNApC88MFlvrAuhZbsN+V04qDTcAs3q9+usjOnms
uWoPCRjx2enBAVKthPrna8rQo9SmQklD13VArzmPNQiWvepMBTPxrhJEv570WTqa
wRFmQHtg99f1jE26QPVYsF3VZzsI5dKH66w/TAtL8reqNEAQzwRo1STZiDPscTCL
z/4AfmAVML1/6md8yZB+LzCrdxR47YMtaHDc/ReAIFZWtkkTfP8ndCFAvJvqdzs8
IyTtMs0YyJt8WVJf/FSVQLmOTEVb8uEQljcC+7nga3JVcESejYC26x+4xkVOor5X
XsEPjSy10jJyXRX05L/QtgK5cWoR4IoRRq+fFWij12ZxMwCxvXE9ig2gEB9FkjMu
w9lluQTaOD2QLL1hblqgMfxoC5bLjHhVfD2C9SzJaHx7emZ96Mnyr1U8ZsLH+zBU
6MNMQ3EwLEkOyQ83jHb2MItXF+R06D533nmSwEAOozDpmpFpQgSipOci3YY/rRqY
ZTVlQ7pnnsEsU8kqONcD+xDmelhmsWW89mfWkV+QqxbuD1dCLxUpkg5fLADWlWxU
y7oOyMseTED+BrMdl/EA+sRMhc1MsfN23K9YrJysnQhU6inWRNPHm9MIaVb6sG5i
rbng/P/i2EZ0vHnrv8sDl0zXVeV24gV0MSdT2owTQsF0BO2BjXZ8VBETknwMYWnf
TCh1l87gxE/0rS1kKTeM1bYDwiGDhlDByeMbdgE1lSYLe7NLiQ9Rv7ebK59iSmem
86ndbieLDcL7CoWQ1oKFygM6EhBo1X0tyhxxIDr3HtnqE6MRy/bCm/beSgtdo7Za
CjuIEod+wSk2TGQU2eOyQ7ioq54O0NGkZOqgw62L/v14WgJQth17RHqvmQz9KuVp
lnLe1zn8ESXueX/+LGnCq11yZ7LvSjO3S3Ie1mpdITk99SPTI5Xjuy5OxT1AedfZ
OMiyG0bhUxJslNaVR4VmNMQUg+JPh/DzsF7OvJzfHbeGNuh56vqqAXBJ1jKcpWTc
eJlVQ7A588apuMR8T4pjzpr2ALb/SaEyY2itvpSTuEAKzJ5vtOiD/yYn639lmGpF
QJ9RKspdmma044XjpwZFBLUe3vRpRAIOXb0FO3gJbCCzf3dmXWBok7o91vqjjumY
64TwKbCdbXOT9LWUc9cks+QHEZ5aIS30TTJ+1BabzgGxAiEfOjvLv3ZMQzm2hgGR
bUTCmU264JbRrWH+k+eVN9cgutK533ekw9fK1mNdaSrBhx8fVDqxWDtwW3HpMitu
4TpJUyJFFf/8KROyjCwyFJrcJI3OxwgpLbqodehY/jkV+4Yegk5RgCkCF2jxq+bY
tGLBjJZ4zRcINKneNFtkBPeHpwV0IBLsFJUseDcFXJxVu+VdoIaYLXkejH1rt1La
YqO+GJhI7FFp+ZEwZ54wobVzzUWAlwEiOj9s84LvotHI+rBVAzYcI6B4NDDMPimE
PfgyY2wxn1pfPgH7wVvWQrrYbVZacUbqMrdKJuZuwqidE9cJx7Wr5wlGotzwxire
zcj6rqfW0hGYalrYlTM6lQMaOj9Y4ZZNdaxdFnI79N4YBuSViU5Rfs2nLjABrVG4
XU7kDpo7QuMnJwjR8jBNrk63yNPVbJMnFqTmfVJCPPOWnKKjCC05rgxqed2tRWrX
BD+TQf62J4SbLblLkN4K7FHFz/AKMsy3+j+9WMI45KBmDk8xdB6EBFS56VKRBTTw
glSseTilttRfmlgBlatDA99Ws2u/TPkaqDgCpmvY15Ezr+NvLDvTGsdWWdX+tRXN
5m7rxVlzqL/fy4PPpk5kI0vJLN1ZgBjeHiIkDVAvKhAL+nVNP8zp5yawwgl8A/CC
s9dQ5mRlYdO3cFto6RCtMaeC38w3rWiWrTS+/ttkncUiKhHc3E5kKrEkjF3R7U5Q
GfZ1aWCu4tHiN1DVJdgXqZQe5H0/tVRPIm/yXvOIhOdlXpE7bTUCw2OKaA/641xp
L+zglkhYCofLqLVP998ykAClNs0wSzaum51h2EYWQgurcZmG34746KtjgZcXtzbk
POBpWJuNWb2KEUjK2cACrheZUJsdZdRwJzJGpOSi2ae47e8NyVVE+Iu/kH59vQ5+
WvE5eJJYlwKgLDzVqKIEFBxvPOIqll32Ie6uAVPjPTKqUZWP6Y6cpSlDIjvvVni6
mYqMbg054+Ueeh0j1Lh+9n1BkIlVUbkjcRWTqS1i7xeeLTT74TZpE+leKOe0D5+D
UcXcy8sF261DHmZVXnSL4bmCWUBIEIHy73ib9pN5nC0FT3x93SWUA8a9lfac4geK
Ccrlmfg2caM7dQaiAn5jb415HaWlgxJJ2/zIqAvZj75ijQW2Hk4JKW184l3XGbrQ
iBejRL0vjKXeVty6xk17p2K+Lvz3QXOKRRT4czrQlySXWPQFp5MX6+oOlcE+YgSu
ISBb68OO+sE1s5bMEdMm51+NfwJJzW9X1mg9ks/REAiY2wPGhwOSiPpgLkuiahLj
EX42j+y4SqKHWzYDfEVs7AGrTP5EHFC6wVaIJZ0i6s19A3UwwPakecNo14Ffh7an
cxzjjoA+oRWcu33E7VSzTDm13DB53jfYD5llVCa17s+X1YFwBRvKFJAr5WBmDbem
I2ec++1bCGSIRZnikV2R84Jdt99x/vqGv3Q3THDS4h7oNNM63kDOCxQ/X/oC8bO7
sh9KYZD056jgxUshPLevJE14YRYoQsO6bT61rHEBu+A1tARjgnLldb7Tca5hRJQX
Ubx4Bscsor9rR0v1rq4oltjhgJJBsv3FXsjryJYhYwjtfn5jn5rLdbcV+sux2dzr
rSTmG/feUntwqfjUQh9zB/dQlNCDoBRkk+Hfw4mjUMFtEtmJtu/pRDHsBi6IR55t
O1Rm+SsPjMGyWqpuOyoE9DSMu6XfpssnjzMnLxodr50daeeYJu7O8lOurPE705IH
eSLwc2JXiaLJH/e5u2kAC46OGHR/RP/gFxRO78++JoxCFT1b7Q4OgY/u0EXGKxl0
e7H+R+wA2Jyr7LGMJu+izigvC202S5ZS6d/JufVVd4eSpQOePRR58vC/PH8v/zVF
M0ygbXDH0gubOAt9f6xnK8DoQQ/1z6LyGMz1JxHmk1dFOfVfoFgvbYgVPxgEEgEH
DQH6gE/uZ5vYOc4kMTF/28js8+mu4FrPhsfA9c+rouiAimdrnGIoQdXpGNWjwwEf
02jOJJaPTQMvtU/qGIqikAmUTowx5+JB/8QbpT9+etbZVk3/FoayanX8Li6470OM
FZwoLtkxeH/VlmLwpWn200Kyj4eUYwtsvz3Rlz7oiX902y0N2aI4i8LLDDu51YtE
kMdFTihJDzo02cqykgcRlJC7Z+KfQb3595VO/ltR1wLH4wWJ9wvf2GzXdb/b2o6I
ebDEGNSVJ7RU+0BCtS3LN7ukxSpCkR9NrYnJHXVTSreqvsRxnSqzwR9SMF3IaN3X
gpPzPgMeCkaKCPmCS63Dt7sLkkU0YYwvoWFpLt8MzTIU9H49KrgglA5Cj7RWew4/
USsPf1C+amJevEMheI1msKZSjWTVM48QiBOo3PzNiOg13vxxvtP2zu01mtfDjENY
pi6BiVG33oWJ7cRJ2doP+4gNNzNBgcbdDfGJe7DfQySaGGWGUcCcJYyvHb2yiFZg
CMjgKsaIlJdpzArHaWRE4A5YH8618sDY6UCX7C9lDhCe/9Lu8J4l3HP5+vZ69AOC
+oOi0UXvQbVeYOycMwgOC68UWPeN57Kofsb+sd2NGa6L0Sh41gg0Vzr4Vb2DGnup
qTl7QQIQzTAFlkCp3eo5LYAI0wzFMJpw7IzzkM/GEETwGY/1nNCaiiVdkB42U/fl
RftiHRKQHyLZBAQt60/lfIKQ4fhLoj546rX8RsxaHuiewBcjn5zDso/ZzXxcOO/a
Lbl/gtbIDzykhqIpBjCdr1B1MgdbVK5eLojf4uMRXp2wG/75W6UZGP1+RMJCW0uj
NDL3w4TEiJh1nUvDd58aXidBX+HDIomRlWeQtZT5jS7Ad5iUOqFYH3JC1Dn4y7W3
9np6n4Tl70c3Vh3yeV68q5vqhCR2vrKsZl0fL5j4P3Yz/KxEmdYArIVRbgRKVUpP
uYTfwq7jGrEQ7tPsJ/txb8Le9nEdLXjVlwpbCKfy7vL8yrwE5Mbhv50UVg11oUmT
8Y3C3apLXmNtdWD+wsHxwCl2mEMru8y1ezS+oyr2K1+1o+0QZlOB4TpFFEKmOjhP
OWBmA4XZBoVVpQFiZD1YSPuc2jlEf+8K6Z3p/EIWtlA2Bij3/WgrmoI99iUouIGT
YddtqrAY6bYzlNYAKAL1AZtEau6Q8Z3a0PQIU+rlt1vpiyy3JO4NIaTTXbaq2ySi
hogVxwb3DSBvcKz2ChS9aQY6J0zS8pamOVxqEpJunQ1QYki0MIjgRLiAp30Ps9g4
9adL5nVpbinN44Zhh354H30N8xOKyQzZvRs62Pnw7OIVvvsE6+Z82QgKrmUy3qvd
WEB4rGozKaqkAhEgRyftFFAMInzvSQv9Tum20+J/KxLpTJFRSpETJDUH4cbwG7Ye
XaUpwte/PZrmrBC/ET1ehKe5jhm75DMZ1hlNQvwpT4pL5NVCxLkRanjdcJP4YE/q
m78bQLpGC3FuzSclF7IUlbH0G0UsFSAuiwnb7B0+qaY28OtnNILA5Z02wZUReshV
0ZLRRx8sdJfgf548T7RKsPXzLAAjAZRCYGtlSitZ1USCc9XUtPoF5+NeMcyFPFJM
y1bMU0+JILhaLt3xpA1XVhq9C0hfWrNiP18rh0EQ1L/OGPpCZ92LrQUesMeSuaMo
ey4NudbYvmELFPbBEl7LKq1wLsRBLlegw7W3ap5YuiW+q26KRUiHG7ABy3N4K2yS
mf7xigFaPjnJ2Tsg6YMjP8UVXVy2AiYWB7fYIyVJDWPEVmpSzJ5LRXTkB40xPpR+
ot8GspB4aGduWj3g9So9ku9r+2QICVkzb7F0Iq2KHUjK2St9rwR4hnoyELIB8CkU
YYgEUhOwkY59o96vrmogBNae2ObDs81kEYq5OvwmEHiLuxPc4K4MrWorEIpk+y+9
EkfI0CgnyU1uRC2fe25XbIvWhNyZOYmhrM0vcpReStdLylst07n3i8bvah+H06/F
Lvdnh6rs08LngHDlgEKgb0nsvoW5f3jvab88koUNfXxVAYAtNtN3Ffall9stg8RD
tehhvulbMyTAiieqyYl36Y0eV4m3/cdtKbFCWNPRVGwykjw184miEv5buSI+ejr6
AngO/HVjlOpDWEMzILuieuIaxFWYLyE12X47w66tR3bpxkrEYtmApDGHnJUTNBzG
0Bzb5ld/1TNUNXlnGJ5p9d/qWZoU1ekv5b4nbvPCWC/xrCTEbA2wDvhdDXXVHreq
C+Qb8pmeQhX1U1ivnPhB81y5cXozkVCVrmGg/VLTa1BIE3BZw0L8x7NQtb09+S/e
OORJT3l+wRarOtUgMCkQq9sa78Lm7FGTSxiUfjqoPXFvWCmBpSN6L6qMICxYIIQ0
rSa5hYs2Rxhk8fWTIe2kX8zklE/gfxTd3lFym6rM9EOrSB2cijf8qru+xHT6HX4X
kaFowHHJ53wJey25IEBwXptlB5K/yAyLA2edDCBAaIqCTX7BZ+40K5fC2vegGYGj
xksuLFFTG0wOFZafH7aBg+SsaWNRvWCBRccrENHBwcBbcnY41CA6zeg3aYijht1C
0ZMHadFjWA7x213DaAXTxH67u7GGrNRjLqWU4sBqRpwUlqfHhiaq1reokzcraVzu
31WNrpRKpuDBQF2sPDvuUhmdhThfhZlmc9EKue2DGcAtwzkSWeFCehtHcbLPXjVS
yiXp6k+Qh639hkGKkTv2yiDgF3kJR+NXCXT5oNwJggA16BkipNO2Y4lQchIYeblc
ZzD0//HTkT/cVCE1EZzFvaZ0mFZAccBbZIMF0EASO8wOvvHDimENbRbgBlRF56Ky
zqJKCH4cNCw+FKH8yaRQ8n4yaCikfDdATVFzDbuWyjv6Ja6DILqKaX3QVGmiURs1
J1Vva6gOtpVtVAhzjFr8lQIGN/nEH7OuBciSQ9XqGwf4Q0BAET2NfD/e/SXhRo+o
rMFMpdiOvQGZE8XQ9HoCZhBeNfNxiXQ0ICoXCaXZS+RQP5w1lz9y39hQBNB6+psn
u54XE7ik/I47b+lxHLp5icQJMGe9GIZLuPbhZyE1mpS618lU2NR+XpyqOfkVZEFC
tJBCWT9QOqnCm4yNDddr9MRFUG6ciXHJsoenEs1SZYpLXf/zAOAg5gL2wxAMLCN3
Pk7hY/oKGz65FF8uWzOXGagwqrws9nrlV/C83AiCutFnZJ7hc5uhGQ9TcyvUVD0Z
q/o5zoLI7ClOHC9fVBTxvEyg+DaBN5PRmsVs6v0KY1EDrXmZan6PS8SY8P/uVP7V
4Slok53SprjUf1XaWGSFPoZUO5I9qviawnVLaIEczaqci3KpVsBpVr9fL+EJ+kwE
XL2J/yJDD6eiF4WWu63o0V+Ihw6HT4qjZvL0iHpC5XJE7l6XYc1jc9zsJ5SLPLvJ
+ev421FkbU1JqPsuN7oavr32haISI9iFU3Cyd97FCyyW1+fYjP5D5IjnrlHN3Cqs
Uxq1PeWe2jUKBpR6hfSIWRlWxiDSgwa4hFqOg8f6vE0W6m4qbGC9d0+M0vVrIi5n
BwW1w/erYL/6M+J1sOK5gyjSSxZVe2JZXK8b7820O3NnTP6yBXVnqjHQG6+TZYeN
GQUvUecGINBiYvpUSzmsZ55JknGEJwelq7qayWKzyt9SUNZDJeZkdl2nj4eeNWqJ
euC8cYCWbWMQVfeSgBJcuifzTPp5fYDoC06B55PN6JRhQJd7X1YsrgHrewXik9nI
C2MbvCugSLaK7zJkMEP1Ryr1gYUm4MWakZKMrBTJJS2l/uVrsO82EUHMNbbhepqq
aH6dQ6Gl3tRgV0EliarU+329gxerhgvdy77gDS2iLgfCp8XhSxWKJy3X8Aa83hwy
ycQX+vmFfsUj48DeGH4/2c2D+8j7wnjxFjTYdk6TQVSHAo+K28KvX+uMcOCHEWn/
E2NdIg/U3W0mPfJYUHJNR9qIZU44RgTEWuPXa8wTApg53KDEFtcd0qKJJBIx2ZL4
XoIvHqDg8KLoF3Ao/81dB5jG7H9tUlvZwLIxVJy1q++G45oOJ3TSsbG5FLst9Acj
uwLpfJzuFZf9fny8gmK/GF7m9CDUDHUjRWsZtfPqwGi3HyUFBEPklRJHwhjnS4cj
MRz7ApJ51R0g9TL84UA42rioQ27PD4JYbz+i+PhaOc9lw6HV2oPGqXsR55ZOu4MQ
uPc8PqNQl/LDSsAuWSUNug6xR7PelGmOTDAuu03TLDmiutoJTtA6VkuKT2zJgeGE
2nSP6y+eeQIvdMrEdIsdnPfHy8gpRWoRBMjo91ksKcTncMWIyxwm5JQS7k/5yND5
RJfqDv+eA+52nLhvmWBp8NvgE1dCqXm44xQ8E9zdrhhMDR6xMRFRmu4dnF00zH4c
V2RHrNRaGlWHKr6kWkNv3BMYOSixQlOjpRpSJdX/4jYUjm6NEl3c5up5rZ3b0hkX
VAx3ft0nYA8TvTcO2m/rPafw1IBcmqaKS6xvJtr22H2/f42rUWa0/d2JxTjr6xTO
IqqQUnoc4UI18lz2pfdwpiqu2FvVwim/yVyrS6poxo0aWsijyWaEK92MMh4VyG1+
2gCjia4j0bNINUhfOa4g+1D8Cv/n9sC+JT7jMYTovzZYDIfpXAketGykJviqZ6bf
40wcHt0X2R3JhsC9VKiiBKOHv6Ot2LGJI+qyORb4STHZ7KZIF+RYF7stwd1EkS0o
QdI/bdNoP2ScUJ2rjoGpbba+f2/bLbvqySWuI6l93/aP6wOV45R16aEk9ieU4/uf
2KHomZFFMyV43/6dmamilnAURX/UfDcbHqKBq+yqszK2IROOkVT2nlm2plrXRhHv
h0tdywwU5bRYiLjJLaxS9LkRNot8uBK/Op/WAWi9iTwyaoQirhG7b8Wq9R+o6PQz
zc3edymkCqB7D58jtEtM6OKu0igtaFQ7uQkBnd+1luQ/JQJobRYpbjEAhjWv0rA2
odu0BPfvMdEl+R9fcstCkewktWHBZOYQuJhSWzx1zJDlurrMrQnj4e4NWq047JZv
sO59rLEqxqom1UY7Si7Q2y0VjmxbVoFGUorT/9150sBxP0SOgbM876oLPAocn0vD
oH4ouoWuZ5YWlY9IHIh7zr+eVoeAZsC9YrtqZiDEAqXRrB0tg7bk5a+qKGkdtojB
Vpyw36wd8lN21nnFmTgolVJYmCy6k3yxsuT5eAs4zWa8jDWoxy2xNXBJzdfJ6Nep
fJ0XmP25mphXLmSVPh/87fVRVuI6j4Zvq3FezM0BQJTAlyIIB01YXV5jiT6o8T9C
KvGj0HyqfkviFPAmXdqb+uJzjS2t7UB1S0dr5gltX3qQcVaR9LhUjyvJb/HFTJm3
XLutgY7Xdhn1ja4tQMrZfbGsA/nyqb1x2FwS/sF8OiInXVMs4xsV4FP6l9kc9mQG
Qvuj12254Gq+ZHq829XPrWm4+ShBKLYPodM7BTwMQlH2YoorerQa+AAbN/eglaK/
Ct55knJvLanfxBZg6Lksgk5yeBu3lBGzGglJ8qUNR4C5Q5Xxk7URRpUVstX/JxRx
yqPT+tX52cc7jpfh2hbLkB1PA+a7U+zFIHCVOkTdalm/8dEYzXFk4qESsxZrt8OY
14GkyfGCZiI2+eGKZHKNAzOaZFBfObu6QCxkvvQfLfWrx6WbHzTdNNG256Kz1fDa
Ou5Add3cNJ0BoJv6KLRtHwyEOVL0NEi7Zygq+NNpXHsz0l4KcJlaFlvWgY6xci9f
X/PsSYgV/XYaahCdHXyEed2RHC1aEjilsLLTMJga25WEkDmdd8r1jhEp3OurSxj7
OTdVCkRrvFZ7OCg8wj/utMhdearc+inrirC2kI9ItKQQN1Bq5myvSLhmNukuXzHE
cGdYKkuBRfs6qawTCQdwjXxjoBtFxcQrvzyuUqq/YSRzCfvto1Wq27+W2lsscptu
+dw8OXvHOWPidIQ7vIq2y0JF3LdhyxnXct2ztLuTdKpD+8TO4oaS0uwBLBJ831/g
d4mix4drV6raiIfv+jqLOlK3Rz4NkBGEr5SNsv2O6AM/EWk55nYmj2maM/eQqfmn
+uCLzjNOR65C1cJfYK+5BeQGacfptnkOZkQ6XHAp4c/nrQCNocW4r9NdvRwWBxNO
ghWjxSbobAeP0cMIka+wC49UeRtcZVm5i4RxqGtdw7P4MuZW6QRd/QSfcDSParvE
P2d69jDsIb0V46cvFqtbuyEwJIWtWlElDEb7AOR8Ew0vRtxKopqZEmQuavLWP2tg
IMIMil5zSqernfGGX9IsyMLhjb2BbVSNdqSCzCYK61ub7dr3ctOAZv4QzzA7gdoo
70HnXH9kXBNTzr1yLJdJBncHRvw3bl77jrRwL40XYGlZtvMGiGckgxXe+EAzHVnS
viTzFR0O47vjnNURUccNzwpXSCbydqObvlMbNodINmVNsUvADbMX3++mtAPaMUwf
oRUujszxhwzMoL8+fSPyBZO88OZKq8NwbxLaOk12AVcLn5jpZkCcUXihoOMSlKqw
sGCPlD5GslAg6RnyfdfNuiviCV+pYHlVEZRokZicORL8Fw+eMjoD0vEj6rKDsdwI
J5hj6EAH0OPd4X6uA6piMsB6K8hL1B3tzfzKELRSXgw7SM/YKh3GGMJcDAqrDNlm
zWgN5PFjbAS4Tcv1ECQgl1Spnz70AC5sR9YFAzI89ZiO6M7MvTZvpfE1qa3P0LGX
r/V86yVhUaBt9d2RN4BAFW4eyxa4p2ljoeWC/IOWZOgKdV1sU8t+LX+iR28q2pS+
WDm/24qmuKQX3P8YB5ZnSuWeDxGFRdqDpwIaF8yEv8akzrceNbNtveW+vBqZdRGN
a5YUWaVSGmGCftHbDc9Yq0tl4nlQ10EHvxJffmiGa7NXDpv7H8Jp4I5p89S9Zq3u
CCelS6b2OFViFRGemCVpJMnvSPdmoJtD3+03JDnOFYcNbYpitdNUd51QF2/tuuf4
ePpXO8kz0sktuXZQNGgIIsXaXdoqBUAQB/Zg2Q+JnUhrLKth2XllltTn9wrru0rB
GsoPzJuaHm2kPubac220WV9l5iLts3k4HP19Ff01H2bpZWgse5e0y38pefqkYhFs
hCUriMLKxm75EJ6nlwNc2uAEOJXQ5zp6vSZJUE+8Cbe+O/8DEfxiQMY1SDOzaSm/
cJekPyncV6joa6MXjBs1aRKiCmqESvGgaukJ0jYCK3W9ZBjIYvGKYEIwx9/BwjZw
WQ8a1vAsuKYYyJ2MgTdMG7tItZLbPTljvMfxrRHtL84O6Th7S7gaPb7MpNny/egW
GmyMve5S6fvkDrhg0geHik1zU/8aGBtkP+9j9kyimuHWcohyP5kxZX8ti4IG9m5W
iq+9qOAyfUYPnRE4909HMI4iUDWxCCmucDW6k02d1G+Llf4J2frrZZaixU2hnrsW
UjKeIY7PE2AYF556JGqfaeSFo4A4ol3yZkVk0RjfMxKy5mKzcV7C4xBLDnrnieO3
xP+mMZ4vsLZl3eJXZOjedTLNZd+FarvijY6R1PAjNJcnc3jVExIbzt0w934eS/rt
ZuwA+5vSqtrlm8Ftvqe10FpSQyNq4XOR8+5iktLftA6iR3w3tc6rh3ITzQyFSWaV
OeqpnRJGMhXM/Ld6Kr9ZJ3iVmC/iq7AhdgwiVcJqsEnW1ngLe1bSkKWgb8PAbP9S
2j6Xa6TQlI/CLS/aIhqHi6f2y3dh2vFz7Nq1fMlRus9q6oIrMJ0IWi1ipm+FMzkT
VzBXXxHrcknKMMZ4HyAwPX0zuVTMmrVuQTDcIxkNtq8JAQO+MMDIpATRYIq91OZg
dBGBFQcB6w0PUIcus2waXcPRkvOw9unJ68z0OoYDtM2lAU/JTbcqMH4sxiI78oRu
k4BXtqLSlHqhoy7DYe9XVB+Qecd0io20bW9xaQEcTLcw/Jc9P0+hgOia4R7+c6Bj
j7+5k0NLHrIPqFnxKrIwLDWaq6d7x9sui+59JbW2m9Qf3SWjGPW3K1/gzVbpnppn
RCukAfOaYpGVtWjDvgAAqS38MIywvbsXB9wtPj9mbFBi9KPSzkvUPE3YqBrRfB6i
CekKWAfXRwmEBe0Jj632p88DaZpm++YuF+RlU/aQoagfniLYyZ3YAY7T1Qn1TfgS
uBFEwpJ11T9pTpGIykG5JOYVIc+TWxpmCYo9Q4XfyQ/tHbFNra1gKJ12HaII8BPn
8t9ax8eLBUmP1YfgpJHe3myAWuNbbjKz+Bav1S7H9BPFCT15qq3ZpkD/qAEBjrgf
R8RQWYB0Ectf80j3ofwzxux3rp5jGCk7GC2sashozY6Y/u7D0DKCeL+DuD70YFO7
Kw0oO646bvSDEHikIZnyw769H83O3/jFSOzVtOq8+R9uKN8zrSmq+sJoyB93P+yy
zYXF02eguA+5DEwcVMH0Rcj5jhXv7/uLb6jm2gxbZR3CLXE4M5Z5SHl2lI9RgWy8
26nF08o4hSMd+KLrQuChmfu0amxvrprMO+yqnveAKvfcBmLznuqApYR0Ne7mpJlt
EDQoLJAFnMPsjJW0afjaEHypoy9W/aNbUi2T/lOC/yUEisYR0znk5QImhZCtm9Ib
cjX7DMm7cp9OLm3Tdm4SgjOmgXj8FzdWK5YPrHCLrQVo0JX4tWAIWzrn3pdraIJP
ibx/qgTIqDJOWnbQsnUmtuMVwNhMc1vMOl7On9FmRse4Tv9EPHg52m4kuAvCU9Nm
KSGAqn670iDno1ZPeD9ooKnwPf1rXzeDIz9Lk0qE6/FfcjV4Mxnm3pE/7Na3WFYI
WjWDSS64S5FRICNqWfZQQLo7/UeImTPpjjmFzXx3tZpWjvCCGMB8e2mefTbZZDEp
hdXX6ziP8eTOYZDYOWZ8tjpE07uamIIdLhSzzgULaQGYOced1s6w/Q4vrYWjENOq
D3ROkNJgp5+O60VUuiqyUwVnolD4UqYTf510OzbLWVeGq7vyWUIe8qhRAMbcsbk0
RoCIZ3nr5AY8YxLg61Lo5TJZz29hATzvD7xKCIzu19I=
`protect END_PROTECTED
