`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bWoY0ZsOXK1jeDUVaAMUhnWdsJM5ZN2AQUrVSyBbok6+3ydjEaiECL88DQfxe63B
mAYZkaJzYgsJW+Lz34ffkRVn6rozpB8zDPdOeO4uJQ4jBP0X8dAgSQCdAkodkUO2
gTE5quqrY+cVBlMRylm7FPWQsN5AWRht27CYh9fi2+76RNFWEJW99uKWyvrieEHt
FrqhTgq8aBh0X/6yO+5vrunulfyETdJEosMCASMKxBcqYmhyPBlhJkPE51CIlZNR
h24rH8RQv0KA8ITJtECoXANo9Lrfzzguqd2xAnyhlM+Gg6sMmdZ1Q0SsEBWqhXQI
PD5gUiVkhLxyRQkk96k1NaAQESUQFj2t7LI5e69q/n8oTMOQFDZSnTqdLrMK+RHo
QAgyqmnC2GBhcP0lS6V+XB51UtGuui76+SpefhxQ3JYSiK37ojSrbXgQDDOC+QFG
y03exWGHWcEaAylLOCDcU4wkuNSIeAEcsCe2ZMF/EZ34wc1Hfcic6A1a3ejbGPlr
n8u2ESTYTjGbluzG3JkaEUi3ywc/mZ8NK0KFoYplg6NvOvjLY+KqeLmUippTsvH9
r612Yph9iVpj9dtSPtAJGFz4OP1U3uZteTs0dFiiyVY=
`protect END_PROTECTED
