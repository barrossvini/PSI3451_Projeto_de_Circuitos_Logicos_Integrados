`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOjNmQnE9fBUgNXD1bxIkCHSdvb/NPM9T5tQugU6YOTOLYLH527gjunio+u8Lqsn
sqgEym2cNHDQOGY1GuvHHuoCQjKi9KedF6Xu0546JxU8dvGPFGgwaKe25sQBR2vc
y6s10yKby7OW++HWIXhrJs/AGv0G3hQtUMa8eYRBB9ioE2wnjddQPgaKYDDBbKc6
hkFUGblQuZw0qmA2/IRQYUdK+1ax6l1frsYOExH1oV96y+PjlTxR8Lc80v5F3+Tl
bO734t1H8aGVIpgocbMxW3+IHIAFc6iiZ8hHkYnu1COdFW2tv2rGImJGB27FFfqn
1OQzJgBUg3h94eb6p31LcZcCT859yOUEE7uwU/GrMumNwhBgWc4lhrJaTvatkmOu
YoMympMdRkg8C9WFLuR2bedD3zagQb+dnwwT6yvI/id86czSdfby1D1eBheY21f7
HPns1hpQE6tYG3/ZLzFKnkzABHqXto59rziWh+jArMQ=
`protect END_PROTECTED
