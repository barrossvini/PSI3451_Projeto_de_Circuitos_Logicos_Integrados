`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ueCfEGwsl5eeh5rj9osQ0kwTxVJP2XNA0q7PCkE57FWybNo9HOcjD0h1KJvW34jn
FDmZ5lZbW6a9TjrC9lurN8kM6LBXicUskbUkxONiQejPVPD+Kv1bQC49DQmwc9Y0
PWEdKAhAo+/pwVGF/AT+zZO8EjznPr0TFwabq6KzPqhRDn1/idyP43jHYwUH5G1S
5Wddu6A1OX+pKSITq5Jg3DqKCXPBgqFyOqwDfOPdH7rdmcH4yFoe08CuwuIuLRlv
TIAQ/v0aYIxY62YHUVQIyjk3fTsvni7xEIzCFtr2pBuwJIRIcTqhjc98snCHLVql
LUlKVVOyJrlMmV3+AR04rH6cQQ3jRk70FQaq3DYn/TJAOnehk4tXWppuZGUjtR/X
UEUhYth+yz7+Fd1bwDihIIPKJjm8sg4t4CF4Jphk3Oqp5bIXQXz/RBvfNTXU7JMY
KWoOfL8r/K6tmmn6iJFuBszpu6H4S7p618Z0Hn/oPEWIV4X5JVkViqkZnCrPwwpJ
4TTxRKGPFIDNyXOlW1nhUCHvmfTFHDP94sQLm1bZcb1M7IHuVhr/YumDyxQ2fH8I
V1f4wFDRpOglDFlTdoS+VEYtAhQg7tzNvtAB/v1wapuuFqCnqVBBmaERM+pF7MQW
T9n4EkTpF9WGlr4cesc1p8jPxjgFL9hJFXl+hTwMy/aGFOWojN+mGx/YBc4idin3
oNbJofpZz46iGGjSpuGh+PTdC0f8Eq+wtbBqjcz0Jh4te+PQ4LzRO9zYOOl5d0uf
nCQ4LsfpCOiaDtLcdQuQhw==
`protect END_PROTECTED
