`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hWbjdQDdHMC7OYgLxhhpt6E3H4QfO+sgdf580NzFX8AsAQRjKRhZcjQLzN2B7v8s
MSq/0B2s1bPOYkbzDKn3KcI4+Hcg0KBzYr/K91oXQjZysxGbVA4DDhuJOGe5hwk4
iPzAdA/CMlkkHuG2FNGm2K87YAOL4ngbizfYDtdJztNC9UaUOCY09koKWFhMqtPy
mOT5pHGMxy5WCHgaGE8x7ykqvlpxSpHnxiFxyay9uk4lGw5yfmlU/43xcq+0L2q1
3Af9RYZ+E1/arJpiLdLdizAJ20wpn/8AfE+rULybOkkzMUl9r86iGFM6bw3AEoh0
6wzdK17RS0VjIaF8dWUtlugZIOUVEgPYKFWcHgHnQkQqCQGnERYgrsRayHJeP9oa
RLUT9Bk2BJz8BUJTYZEni/m08SGg//HZvdGLrwum8wXGciMfH1NqRbOwOwas2N1S
4baTc2hXoM+YIKE1XynswO7e/N1JGpjMRgL+v+wh1lGqyhquteo19RVVfmuIeXdF
F6EW/XNqpp0EFRKPBXa1qpMjyj6u4Plu4JmR4cqRzlCjPGW2nSslYWGdxwNE+Mjh
DxyBr5i9Ht2ScljyTikoTzp19LmDhfcLnKgAfN5D5gppip/rTezgifrGXXawX6/z
OF1VSAgOTM/MGWHAvYuwNNNEtdtlUeE3VXlbfQ4mKRIJ54i9sq1gAYXk1HCQhNBO
5/ycdmGNECHqYz0wpjJUvpZe8Y1YXViFl4j346KrxsLMDfPaD/IjRlkKLiErfOhm
tNpz/SH7I58FvYvjJJ1zh0JaXjnKjrXAAgcChmvG3jy0ZUSXhG5pO6xdXn6le+dM
eoow7xrO5Se7grNiAmTZXyM59xJstlA19yEGKq3Jw1ih7/hIvWm9KBhvGjwFg9ye
XDMWoVQ7uY12YGndspjK4Sv78iAmUYKnK+mVi9he2n+71OPGltvoMRI9ibZ8m/77
r9ulGvaAXEaj9uUbKNuFZ0CvsLcT4POWXZgSxBBXSSY/OaC8eqkcR7E06OtAvicC
qwOCgWxPWlHfHIXGOTSWFDi64fZUyEds1aNuP0i1DzJGSblX5rV0SY79lglHTfyq
Fqd9zCtNzjPYkk0IiDVBTCn4Rjp1rFe839m3LNrHbtQ8ZUyrjO3ay0ZDiDi7Xbh+
/lHka4Ks+aMPQdwsiFhsTfz8v2qEzEy10uNvrZ8f4GqggtYQMHv6vKroTMAQD+6p
A5ywB0lozST/Q3QbEtKWkDfVHIZspm9c82sFGonRcm8pW/EzJMn8jWvJH2bh34qW
AoScA8KmnSKHF08kMJH5iEUdRluYo/gx0XP8tXeg14G5DJLeHyxxmDOqc0LCaSy3
CVaZFQ/EhyaNDQcKURsEDbBxootLeXLPqrqE6yNHJ6gxchFZHNFmrnOb7ZFE+I8f
s45teY+iNCID6xArGMRiVxnNf6zRCiqaoWrTHL6NCoLhp0ctGSDaQVuK1hF5EVBD
BdWypu4kvwQlJUz/14a2rIw1HjnWG7d8x9YeUFea4Q4zjmRf5F37L6slqCDyZk3b
ja2bVaqIJ25qxSIqmxoXxdM0BL13kF8W797C539Ws3GART3f791aS+7k958dWxOx
U0o1QSGmC326nMHzMrlyWZ9qa2Wl6IwYLl00eNE1+9hTp2bxSbVRjAEJ4W7lYOrO
duhyo/1fiDNw9UTaSRZDZ+xcld82SiFPb4FcEwpSVh9rsMYDA+4wqb9+oqybqvrP
vr/figmpe+xM0cu1SCiOqpC8nxQRSFDzH5NcnF1nqLSw5E4MZbE9mqBjwe0BKdk+
ts2CKvapL0w9ubhoU77ABJyn2NNsXi26qLHyRQPbkNPIvDrogKqfi+G5TDtGwTer
DS2JmNXTdzjKWv3LnHrGKrtvMxALuwECWVZ8pizHU7GjFWy2Lf5jK0pmP9DSfMbP
R1OuJSJ0eNaZm8WWdWvc0F63N8nD9vCchEp66oDAKblrCyIpZD6StHNryrcTBAgG
h0n5dBNaf8o7R7kRFp1TskaDkVaThjBwHsUhT89ctBGytQT7tq91SQ4rarmvbTiq
GWIovLD1KX5Fvg0R6wee8HECiFOtrL33SHn5BNFsR/yx0A3rvmFRYLXiiFRy/Z0q
DWhvYnHAhessWjXQvAcm7zdCMO8/VW1F0cAV9avWwa0yCj6GM3gD+IHHgG6KOqXj
z7jcitXLedJA0BkvcT+QzybW9fIIfHzQn9JTSXijGWZ5GnLUsEz8QUOO0SUG/tvD
bJIreHfX5aNS14jLnIjcUAZQ21UASoVSH8yv8GMBOnzZbHx8qKX1ugbapeiwiZAp
jLUlUMcP+upGNoVEAnM9cYn1dQo7pibafZTA2/jCiet06/0zRbyqptad6heBWPJK
FAtRHrYUQET4i6j9AM9V2Av7dXFEjIJvHKQ5epOGxMBn37Li98YajWbsLEL4legE
dDp9rEu3PEIINBqzMSwZggRr5D8ehlMaBv3MNItEzAj2GkiCPEY0f7Us6FLp0TXC
Ir25iTzlEgqS5DAVn2R9wBtbqdKAalYjME7R+sZa5Fw/MffNI1doaCkDzqvdpx3g
fSJ5DK4BahW2BBMuTOrn3TnEMqql9u9ZklsiuP7p5+++fXuJLBOT+ENNXpZgrAC4
aW66zru4FBI16p6YbTavisdLnAmE20O5WQu3cvfk9j18+DdVVClQ0QpCedbGDbB/
3ShawyvnTI9MK52SAsiuVjFKsqAakImNgu+A/uF6mrNyB56ZpHXKv+NF2lscXIlV
`protect END_PROTECTED
