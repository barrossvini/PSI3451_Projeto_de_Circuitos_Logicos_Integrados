`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JaEnFwPxknrfYp0p/4eHsTZ0/O88wjHOIRH8/dwoOMmnKK3pHUJ1IwbThEHPMeFD
yJtXJV5DYjaf322UspV010qjhCTq6PbFHsJEIZCsbE1NiFEFv9yG/QmmcZblSAOc
mlpJHaXepw6YtONR5VosngkyLD3q6eNtFhvD+UhApl3lJzsBRKEGzSaTYnzjdClH
y7rGripBF+M4uirTSVXeWAVwpeJa1a3TdCIbV6HmFEa3ziFDKZXvpBnVfuHcq7PZ
G3rLgknb51CV4H6UmILC2gGJ+OuYq2nOXvW6wFNFXCE+IStsQYXGRnP9qxdBFia6
iyQXR+IdFSHCm7j4LKx6CkVXNSm4tNvH9/epvu0y0SALKcA5upNyyJngOauN9N/A
RMSKM1XkXgs4bWtFHVs0cAJTViUI4639nlCJHr20RRWvyGq3TLGtePIQkFmfqtTO
DHOy1D1/M9Zh7Aw+XTLvCltOM0eduZqsi337WM3JoY+cQ8d9pSGK6pI6JBOIuriR
3Bh+FMV8d8pgd5scAeptuttvYOjsAVEFcGhSXvDCMhSyjKKXIWGiFdYmt+7u8O15
LAB5wk1csDjvcRt1FaKWg6EoqHVf8/ERUjeHX+MUBl6ujowa7lturTgYgmxZiAUo
EfZUxqH1EE70jDJ6vDdvCZHc4NQGZB4kZofmDXAeR0JQ0KehvyUH5r/MAMMe/5Za
mT6JHitbw9+RapLR8lF6yh5c0w5PNxuQ5y/dAJrjdcJiKAACT59XeSxUPFn/c0h5
D/29NCJ4Z0VhHZdfgojtz5U2Hl51ciFfC8gZAnhXMBwq4aLnpjqdA6gejPySqNZW
dYVy+RryQOhHzK+HID7wDtg+ZFO09690T/a7dh8gKGEW/L+a80bYYr8j/dK/sjE2
9XgRr6mYVFhwQZuTnDiknKb54yPheBVGeEUBNRRBXBXU25uScv139vwOz/HRWbRy
`protect END_PROTECTED
