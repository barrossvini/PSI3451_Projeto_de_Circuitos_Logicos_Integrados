`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QRTVH9c7flhNQZsBNYFfJyoCC+qjCM3+OMXZxR5pl4fxN6mJzNvT59n1TsDtVznC
mNUDIY1tL1GUwy8rQzw8Y6jkWwpoy/FJp2us4YfApjE+Doyr5T67jIJSMXd4Rp1X
U+igRDtqNfVStGtijB9EESzorHLavK7Lv5unaa0FI47VIEgfAEYHPOlMv7fP4eSM
4e4wmzeHZGNJe/+I1KglBK7kLjMAjjQQotJtZktePSl8DJoN0hK2a94n/UedBjXm
A2kX8dxKritn5pGfn3KvETUAtkuY200v8fxN4k1rdhDzeGBe2GcUm9ihRZLsU8xw
VLOCNfbH7ZYCE/XvimzuUnT8rKEhG1HZcw7vhe5EFDGRnFUZm6Jwn2xMpOk9/5+Q
BcRrJ8mOQcMiQ8L+l3WTtk2PzE01gVcnO1LTBFdmwDWbFBe8WO87HyAwQbiNAoXg
mM3pu2owhMK99TMVfxfIp0UPPYnUYyyFtA31MbUwbC4u0bKJC3lF/JvhZ3R0txXC
okeoKZWCNQevRb/3wKsGL+r9SePXfDzmWtEK1Ai48tvmxh7RgSadFOj0cel7WLe/
2ewYQjMINM6Ja0UcOqskNIsvI5UbyZ6epiqF50HdSI30KXoB5fxkEekjZXLYDNi/
`protect END_PROTECTED
