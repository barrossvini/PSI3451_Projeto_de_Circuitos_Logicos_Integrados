`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1hQmyeiGcOVYOxMC4pw3dXZZTjTT+H440VuYqSvfC85p8WiCewebDsA/kaGeaZR
/8RhMFvOhR4qJJkJNs6LiDto9AWXJUFE1WHxsSlbc8zRDZhrrbek5GDTpGjsmghr
efqqdjbJC3EkXmI7yXDzOZlyZDMeps9l36T1UMIN/02BvG5XX+pHUFrevbBxBAhZ
hc3z0vVoF29mliwXnd1kHg94hh0r8AcWXQvqkKaEG0tizdpr0IlzR59GYEirRq3F
WGxDIwqlPUtIHMpNj3Q9GDSpaqmnGZORqRmRUsDONA6qBER0RkwNRtxF66JbOOOf
2u9M1kdQ0/WlqRHWqYPsQmO/9X7rj54yRkWi5uhulvbR2XhlVhUirRP0gqOMHOmy
qGEXE9pmu4m3T6FklHoMEyz3Jr/VuVxx/6S4wwSYcAcvUlEtHK93MGP7G3c4M5y8
7k1qlh6qFc7M1BtzGsELqx8eowqeJ5GO7ly5Gu5wVSc=
`protect END_PROTECTED
