`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fb68npzQXemTOshcNHC6VVj7pLEaCegiQf58vEr2tkm/h0sG73R9qPQznVAE9iK
QH0A2jYIfC7tIZ/y8dIP2XCqhWu6SKlKivtBSqNppAmfCRIZN5N95Ll3wjNWLk1v
i30/Kz6OfNkDFdF7LjlrzU49PBSWztKAzHKUsP9QL+s5izvWOyfx73SlkD6ZbN/W
hSzrN9dE84GrAWiAlvaDq1vQqVQyD/2+zFSaf9tfrZhZf4rHm4SXAFnDrQw9+vMI
kv8vxk2CunkoMWKbSM8Q+PMYEsbEkQ6oonIFPz6fMAPBZJRUkdjRYlmfqKyCEWaU
y7iWQeqwW+VBT2t0yXtk87LPysu1UiTqvVkA1mRRmIsNSGLh2S9dgPl2OyMpJpdZ
hGj3Z8bqPQ8HhWo6mWa1af69KkTY24cuS8u1nE+ZFMdmJZ9oOtm2ODqtddr8Mbqt
KKxvuzzugLZpsP4oZs6VhcHRtn59e9e9JzuVGjSuCCT44Hwkk57AoUa1QXJMLZaK
nbRjEwv+eWI3CL5/oUw7Jfe98zsYIpQGiDdM23VT33wjn80+fm19pNDgfHS+EPAd
TIJS6dSkOuJxtwNAzWdmPHzCMggAGACgQZdepPYlm1FQwOkqs0qRdF6V5N85DOe9
wRoUvnb9a9cFSGjD0UZN8dDHKQ4Aflx9pc59X27XHG1xFIjb2FBjpFu4VNigoYo3
n060+RnzYdM4hwhE7w5zIensztvZQpmWDTNSeyE3nVV4eT+fK5MvQG49kiqG3js5
UKuhWJH8lsWJndp+J5JIMJn+p2mEENk98tAwrxHMHKGOl0T5EbhYqcA5osrUmtmg
RO3fGSiXJWi1kwLxbsq91GXkbcSqJIU/ReCeKwCmZR8utvfk0y8ECoTXriypOSHD
SBCEEerfVegmbFCoiP7e2daEwhNicxfF8qKi7AwE4QEWXdFBeIAG3s/OR223OQ0N
ihS2jYIYVcsFvr1z3RpVJ8hspE4zU+QFHrIUw9eCg/7OJzruub8vhhwghTGxXyZk
C5eS7f4KLTFCzS3TFP3SoY1FeMjJg5o/qV3+uRPj9lL69C/5+e2deZm8BNAXi/i9
cZ7QXQ7Lh49pcwkRh93huQK6a5aJzgBQr2L72/EqZGtL6MK+p9BNKKggJihxJzry
eFonIIa1c+VO+/xb9z60K80rOOwyUb3tHLWiyC2SkdzBJQv6CJ1QhvxrR5qqK5Rh
vigQW4D3nNVRJNduH6dLCbv0eWvL1GV6uKy6aBrEJ9tGG2wB4d52VNeIaYGnMtg0
r9YQrb/HqCNs0/tg3e1AcifPRmScxUTQOQsJWOGOkyn9ijDuIhBs8is8GyH9kAKW
Rd1nmX/OKxLqPdhinlQAu6aM/iAWTNKlxjPIIdxWltXZ14nafKiLAgAr8si1Z7KF
QWxpIzXnv5t/XSdKBQExyp2G+YsONmqSP+Z81wQAF52qP7pYZBm/NsAlEFC7snwr
0K2LnAQnsw0AjiFbP9i7XkQqd+rk/MPvJSvlExWTri6AkqErueP7knUv6haNDCFj
KMlNOlP/xuYsgdYdIdrv/w==
`protect END_PROTECTED
