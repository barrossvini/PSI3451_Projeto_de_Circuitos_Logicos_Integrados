`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
59GpvxjJSrCELYsSRG07th8xE4euWTPKxKdTtiWa43QZf1U7YP0ajFqQGIiy7uq1
C+9YQbD1d9hT9Z/C0mSaQQEsx3Q4F/LDDWxPaMuiJYFHlqGZMTmyEbr9x3fX2Cme
FlW9d9xbyFe/z+3Je3Kp07IeoVOxe2G0ldH6cFzNH3AuGELv6nOpzlCsu+IyA8fZ
nozbgpEcm60Vy9hlC7FQ2Wqc8LOhhjQpdMN58QX9vl/DADgYCnrLcQJTofvglost
SfIyF6YcGxnvikDZZQVg3Fy7vbXCQl7uyzJRRk00njOYDSvfBy88eE9naBtYXGO5
MC8/z3arR5CS295Fa/m20JkAqKwQOkiC7qLh/oYe2mj7kpKfWKXAHaxMJSciwMsp
KR7/0z7hT32Tl3iFEqOuf5AH6J0xCDFOP4EVk9kVkrKyTPqtUroPn4eroEz1o6YX
iKmDOgSjU4TrHFsnGD+XpnGd5UfAgzFV8QFhBsf+19QhnPyoSA9dPES6iYR4K/PI
NLXFWudB+MjhoQcDDxyU52EIshxaVjLXyUsInaCF3IO44B7PRiwf9NoAcPvStoDt
8VA+TXkP2FP/2/HLEifh4NeHb5N8fG9U2AfAWH96X6Gj8gKSGoaHXWT6WDFg9AIL
+HAW1899eYo3jwmpTfz9t6ZCJ5Scm43tx3Elphjel8kvo8iv7rUu/QpjTuK4euew
xWDkuMSBK/4HpHKJA3FidKaURtRycU0GMBySMrjha+LOK8T5Ub+M93T9WRoFBU08
CT3QkeLpUl6WmQpUXNmS6Y4rpQ2zQTOdvmI7xmmD5rg6neiW5Sa4Y81yBBJ5tYCA
RAkOLkgijzEgmI6FS7FFxoyMBRjpUEc/Gtvo0wF1A31Ws2arALo9F9qOizXlhhdD
IjgXbd9E1b920r3kcbOFORCobpE1QlU+CV9Slo0tvsytxGv9B46iG+bfPhbvhKyr
wREe74Q9Cp3F30Sgib7SkKPkDhCrkw85t8U2vIMbT5vtqI94YuerbP0LyuIJzW3b
fDJTvTZIYobzOsV2ICPytpOMmRaEJwl/ithRBDuq67rK8+j7oRZYwgdTRknvwp26
uwUUPgJHzrCU5yQGgOIoz+XK4LJMi58LMx1eV0Hm99nX13zhtqq7DWmpRCrE0JBC
BkCg+jd+Jj237sZtpQe3Z1sdqaT68YBHo2pRw07nfpejuLayic6GmDaIaPK6Aw4X
SlyXpZXlMHq3Jp7Av9dk3tWaYcLEZnA4zQm9HkmXuaAuIEenYVc0lFwb2hZp5FHt
qyIwhN8zAHBsc/ReeSyvw/uvkkrj0S7t21/1cmYOFnzQPoi30Nb9eWWJsqXVq/zD
WyttBiH3X5IXRV1QWRlXkBWUlh6upnrZPNll/jfB7MsvfpTC2WdVzd6+O6EZZaol
kpbcgpnN3zYfXVKWD0JTrac2Ma+VBsrqm1cHdaXyffLX9RDrJpaPN+yFqRuPNrrn
/al2bsjK/UW9ywBqATvSyoqjmRRnVsigcccl1TSsF65XiG3vYCuzFiUlVOCrlzaq
LyNFPGjE34K3QaHOfUhuETNoKYbwGCVKu6o5J0oI8+ZGe+mqhOysn5nHhfdfBZwD
NWV62g2uP/QR38nEpvCseAXK8JFm5ehXcARhabf3kQFLfSDjtB+5gtuccr94mG9+
wB9xAk9AxgYC6w6hCXzNPwwmmO9GcmzSmn8mYdI496BTxFNoUKNz5oZxfUlue1eJ
8Afk+PzsAzdbd3clVmwoonPV21X1NxVxt3OmZ/z/s5GvRzS0+ZdC+QrjwWuVo26d
hNGCKMkjGJHeAw+8x6zohz0scLa398KEDdRa8OVKyMKdPHIsw6T5nSItARFbxtTH
XbseqyHino9YOVUiHci0oGOvk7gDLljC9khPyK1KoJdYSZQ6yS4LVwoY3dbAYV5Q
ByDZdlJGYyVZWINCahBvHGlf3n/KMX/+nBRW/VAAuCqykFF1SoV5ytg6A/3jjkg/
8Cz4aVWJoTkQVeqj0237BmBDKrqvna2Bd85wrQrqAcIoCU5DlH8eS/yDolt/5ugZ
VPMp3nsrs+HcURvtyu4YEu2SJUd3Lwp+7r0ccqgOKddpzFCzL7gEYsqujmifZkPr
qm2cPbl9NpLQdXFdx0/+mwiy7/nIJZgBx5a6qQ6KcsG2rBpzIX+B5FERvQsMBqLy
qx9g2PGh6TREII+J7CWnRWszzh21zRzzcSEfXkrxOVv92nqS8unzqBvGXfuKJhg3
kHYT9I8LwSLVgz78ctrqQGGGfkGlt8yDaVycJBGCigBfaoMtA4/4AeHX0GhZA3yz
lo8tM1Vlxvkb2Xen/HyTS8uoyAdsA9IlZpfvE1i3/xnVmkOpfv7CJpYgiMA8yU9S
/8i476SAGhPWFdvGD/2DDN8ijIFVFepjiIYPjtTfY2d+HEFEQunWnqlzNRvVkSxA
/OZmYEyggi+MEtdRR+qeCIExCvvudIz3Z69mOErM3xA79Xf+W2J8JqpdNvkE1CEa
hhs4Hq2CZ/uH+Lin7FfuMA==
`protect END_PROTECTED
