`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H9tXuQgMr+XP7Ryfc5H4gTiRBBKW+1wdzBRD6Kqnyr+2idbiI0rnCIOR87mSuYir
LbANXf6ZEZKhfMcAM2nezDqxsKQ0A0xR6edBVv96vk1RLnXHSoekUW2+CUM5Bqrl
zVZDSsPUd6JDW34jqdJY+qRqgIJ9+R1GEjVXpIo5yeROrGpKUVDYLVjbZfOo9JZ2
I6Y99MHZve8N9Nh10FI2mlBZwIz3DemTca5vl/7+82n99RG4METxoA0chGp5QTwe
srbaACUzdLDEcqREQsqqZbdbcRUNqJ8JIRe7Hs4ETfDmusgzMFdyGDg5BGZt9gkm
DHNoa94oR3YZ0UfmQ5lHdAB7QEts/P9AEbVAV2jA9FNXWGZKkx3H4fY8BDPCNa4n
xu8rSa1a5WYFbMrzOIomHW/X1nfg9lgFnzXTadnQvad+HE4FauTGEriORZMnRfk4
KFrBtMGxCoZkHldbiSlN1FgHJuVqF/fx1J6TFpj/o5XUfSQesop0IzTU4GHNjK1y
TinJ9YMIXRAcbBVmmSmdKPOKpqFb0qbby5UaOjXzQv4YEpOSLynSJcdqIxWnMLGx
dh+Dcwg67j1Q9nxZlqe4Su/hEftSqGE7z1YYWyt+qzTre2ASReFzjyAQUa6nlsDp
bI1qxqa+giRIGA4XML49wcAS/SZUar6DstqlUP9L6xTgWw36kS6SoXA1jPUykWiB
Y/+7+KENTBuu35KG+Xn/vZKgwsTASvos5Tto3O/Fh+vNZ4ujipK6WrGSeNj1vT2a
AoKaJuVVvgLJKDF1lwnOQV1j6dDX9QTA4oeX46WYVCF2I+OIRVqpOqhHPupvjRC7
wEDdO98Y8oFfCY7HpKuzC4tLQ6QXIa7C7ukgmsdTODd6hOhPbsFUg8M2QkqBZKII
zPe4BgqdLUGL6EohpzBiLJVdYIxp4aXydIMFJDKl9hCeXky/qu2mET9HcPBIuYq8
heSCx1shzPJpUAxL25ZOv9I6KBuSuH2mkfnleb0eysCD+RE9i2/0oCDEzAgXdaND
Rvzd47KrOO0vFYarZN+t9u1cBoQxuT8TQGdFwactKlHtjDp8bhXSSSfCpyrW0Qwk
ObJxnMhUz53mfwDGseAlA7eTZH9wx1RqgIGdNzMZP7WdU0xc70MlKHL4P/Ice7vn
D5atfdbuQAe6YH6QaofNA0dcLxYTR4AhxDmftGwsdE7Tu6S1JTg8jaJhcla0dpCp
aWMYfB2UeSBGUrdMa1EFRAdTmRO1dBKOUn33FX//KaG1cSq/QMTMUZWGfMpYgtxE
`protect END_PROTECTED
