`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i7wZHxYxhv8bV4ChalkZ/vvVLbWlDDFA+O+q2ehUKAt9DZ1JB/wgckpE6Dgz3gfZ
Isx4/6AeDc3m4OFT2gwElfH2uknksz7s4LNyPPkAB/LWsnhXj0zH5SwFqA9+HEka
cbbNnzA7M9z6M8znWoiMJCUgrX07MszkZrFACd2zvdxdJEjOjYLk44zUJyyAk7Di
aEX81dZl2+vG8NQd5oYiZ0pXr0v8tsmvqNnFl4CBBzwFlfAFbYI8b7HEvxBb9xw5
TQzAmrnHEMg7e+4JAuwP9iyRRbrUXbci8YNyebeemG7OYZU/jcGMRKnjokfPaCZs
Ynk0o4Y5A1TnNo6ZnjCxkATYWebWeRkxU4BFAWHem2HFY9p31ylV5LYsuTlxtbGd
+p6UQqIzSDPTGdORTgrKgg==
`protect END_PROTECTED
