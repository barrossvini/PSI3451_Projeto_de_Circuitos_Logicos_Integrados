`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XML0wZLbe7vv3D8ZJJ60gMolMI5Fi0mkMV9h0kiY6jNALjrMaj8r/28mapQ8Ytzo
I7AbtH5rTmjqpS+gURTgqJmtx+dSmGsJdCYS7NSEAhwnnUzhmI0IqBr1rJV5gCgy
hEdFlNwx40RBf70Mc+czxkJS21tMCRzL1jQtUfOdEsAAYurycADYog3jeISeyQxv
wspgI9OtvndhNR2aXTZldOCD1TC4/LcZBj31qrwbmHAwuMj5SMHw7r9GdtmAXdma
Hl6PptLPjb/1+idvqopcwne+b/4/E0TKlZEHRLDgvz4696tBReLDIP+uq0UvBz+I
2wxjaNYtM5uQtN4yvAtkZF/F+y/FURfLV5x/TG+51OPxKOZHRcRDNnXP27essycZ
8r/bI34QeHPxpsjjFORvqc0raYJ+rFqEuEmBjcsYbNhY7CY0hDk6G8gtF4s74E9f
389zJZmcoUufkbzm/aGaFIun00OsPypmsTimm1GoUbBmMcsIqwNbxCrmE2jsYgil
9t5rwh8RWLk4vcQr++FE68loEJmyz6GG1er1S7cGPSkXgRjI77LP7LNeyzo7dICn
aaQSomek8yh1IiTJZOwd5i+U4cyzuKZ7vQOIrBKTukk=
`protect END_PROTECTED
