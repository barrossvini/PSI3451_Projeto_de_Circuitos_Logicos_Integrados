`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nF8oZFJ0NIpEMBWoCAnfPv8KoITDMZ/GPBlMBEcOigm182A7XQkWA02mXgFjVfab
1d4IiovNv0WqdUgQgU0nsT1Q0brVzMvqt3/axKHPjOoFIJqPPCwroOVVD7PCBnch
f/sLp8m3kPDZj4uGufuyo7AiWZSxnxHdUU3I7u9SHXyw4m6aDaL3J7dKjKQbazvj
0ZbNA4zKL/de9shHtTZSACGHJdDcrBZBMA/GIr7PnQ90dFd3elLdkyKvcfbEN/Wh
YU+wTUAPtRE8ppZJge92ti3SItKplJFeOsKmf9NehVh2vngn605PwWQDgrHHzkSd
Sa5Qft49yl1dQu20qMtGjijkmE6++EVz3mzrG1mTNnlD/IOY2NkAvsL/HZ0r6XGm
gTNZJKbPpjab+QBhvtTl5v74MyndL4vNR6256gb/HZO1MEgv/xlyr8iWV4j8MKbM
QQ2oyBZWsF/7GbYBHs+Ux7CiTx1NlLJzjlXwDekBAH6zMpMfEZwKaAexfkK1QzvE
YwTk8xxK22z8jy8CASQke9KxJK8WedgmzGHJgUCY5eDSWuipghIoZkCGiNdyHKZZ
9jq6g1xMVPBBj+oP21dRUGWEmz82+mQ8MatdNMLItmiOEFpIt9BWdK+sJYFx5v2H
W/ymWGPVFvFTVOhcUUqaJxJG+htEvH5HUHE/TdHvDpvHGsmAj0iNDyUSLxnN4AH7
aDmVpuCqDhlKzZqpse1TwTtMwjWactZk3LNsJn5sYEKnALMhMASCjcJee75wDdvP
UQKLpoEaY4Vz7Mqes9VavU3/VYIGZ0FCKFNgUbiwA7sqUmXsT1W8IUptLtF2Uy/o
e7mVHheeNwBhr0jSD2Wgp0A/gM2XnQssGeY/V/HvjBWqiaMbLZ2f7fm1QRs+g0eX
Lxcy9jXlVUX6PLGmyxrhq/ChlhkUqF55DX4GnrgkB07quEDt02Tj4cOkzy4ZS5pl
5BrjWAJOEzP3DBsAu+qnPNI+nm1rM+Tuq53k8WL5a4uMes7j3NFFHMzB8UzRmmcQ
/gLbN9JmftcW/ZXsGTSZc+8LAq10nyzurWC/6yVdDS251wLZZf61LgCYcjgU6NDC
wrEB55lTlcDMhMgJfwu1wnImcsz+tbsmOJGXk2qEi+0pdwsxHs50e7GLJFYwYDzw
gQEdOud+iJemQUxvzNRUL7NTLhbdwDS8ErhnDuabdzKoqj+XuQgmuoaRhFbK8eCj
rfKhLPmxs/Lmg1u7AD7wI7XvSWYdhH7dBY+OJaECkB5XQxmY77XuHQCiZ5ZpW8hN
+/Bhik7yd6ouyy8fxmhh8tpADBQqDu57Rklst2gbUuMl6MbKXlre/CfXgGYRwhzP
Gp80fPEWcdZ95AOb3b0zebFX9UqNP11E6qZYZ5/gE2dtYsk6iEI97vQbqTpXUDVo
5M7+KGWZdlaZK2x1ftF7jKTEdBEW2XQQCjcyZ1KYF0IqCSjIrxn/TaSjTr8hrKvg
f0DcAcfrnr72dQRyaUIT2rjn8qyFKPwQXpKVOCZIK7KVlk2ezKK9e0cizw+ZOX4P
a4gj5qFKEZwiYBsoVarlBBeMPvm8yJF9JxwttDhYhIwUQdqMLqS6Ci8ehkGvgIJW
oD+05NyYQ0mSHa2Bh5Bt6gSuLXhGFPFHYb0JJkRNfI7iVdMlG0lAYLaomjxCS7+A
6iy4msv/Y8b/OxKoP7QVSm/eh8O2wk95ACUjFrARSKd5vLKe6NGQirtV10mW4sCy
1oqESRZU9ZfR5wD2Qgp62dHm2dQ+MhAZNZIGAyPh+igBaMzwqGEUv4Uvvp/06k4+
wNEFcIYpG+nq8j7Ua18AMLmqwpsrI5UaBKgeqvb1rCCM51EQhKBbyfdLMwHYgA5a
7foV2/YezFS8Byxj+e+vhLmhFr+WylzpuL8n1lqStliDSCd0GXJbE4vJV1yzTl75
fwW6yzs0Dgk0bm9X9Hu/H3rPoZ0CzNEe7Hjt44/UeWJPBfgDUO4zHX7cQnEXeiCF
uvQJk59rFWuYBD8MKhI90BAYI39PLUWtvH+tdMLy0I3t2ml0hhg/etjMakVuFM/3
lfTIWhvZ4a3F4lIaQxjQVbxGBEg3pvQZRtTR0dFnc9iBToTVBocrj4xS7/0EnjWL
Rcx+7kcl8NLkbPFMfJezTIbINFqgxbutWL+m4tZZj91llbEkUOCafM28Mx1paH4s
fIF0XCmKNEts/NyKOkwVHFQhkLOrbSoVv2pMqjxM9fYVQ+qImwNmhVydzJlYTfqo
ZcOAQv4usL8FssP6Li5VzONliGg14raUwKK4p69s8QfKUthWZ9yyuIBOSEQlIogU
Xp5MZhVL5DMcRyhmlIotbyw991YZLez4oHMaBRPvGJdgvhUHo0s5pIMJdl5u6bw0
INn2bAQfaR6tpv7vH+NdD1f/EzgzEAOm50boOhAZkHjNJP+/paGj+abhCwMCHhm4
LNH5Vzf/ErcxHJhGPZhoWmp6uctvEHzXsCdkjvyWSGMImUlWqvw7HETfyfetmsU3
HDy8RzyomKiqTZMFQGKCn5yK/PU8nfBrQwlp8npWvRIYREysvFULw8IDE1q+uCMo
H3doHAdO3GMhxj5VUPUeyKtaYj9J23tH0LgAymthGL2t6VCx7c1uTdujUm/5Q/Jt
DMjHA571IYi8y+dn3t3yTKCH2DSNoFGu09A2zDkgros6Gzk7Pz0n36MpPkAwUfpH
IbKlIdTV52F/jHp/WJ32PhIWKUGca794UFopUi8puuHq0mSQtxjn24Z5+Wdpp/Ed
xhf/AgfyfyylgW13bTgWtdCUol4b17IaBnmhs/RenXkXvme2Dxgjt2HzZY9FwWdS
ci4n1fSMUOvBDiT040eUJaXFT4Jc4FmiiInEQf+opQqKug9u5rnIi3QTE/vajz3e
BwYUrHq2LjiFpQgC95n/kAHmsrJks1ICGDdRhkpJSWnsDToGNXgbN7rs5ZUz3uTy
4uI8nLWGSBmLUdiJG++n7Y5wz+uTxPnV01pQk6/MHDMvF5aG+yql0kWdcPQGTqgi
uBuPkWNWB4X8RSmup+Q/ugkN//sMDamiP/tUxrlK1uY+rNwWmdezI1e/lKoGP69h
WyYwbvQ8/PKAC6LFTSgwKfSe+vJ0yWJ9e3HoO60vR+1mCJ/Nn86mDu32ttKVpSjn
FAZ1A1e9k37/Ld6Wqmn+knsWuM16eHlNjLEWJlKQGTK8rjx0f/+zXeebBhTHc+DV
9aZduhFkg2+Ve0WjIilzlYxGzh1DL8mKxBB/m+8XzRoFECNnVk2ncMqXxLCIWYrp
y4hgiEPPU7z/efBR71BisZkt88sn9YrqRmGCjyPF6pJjJdP6evDLNGvQ3P/6q4Yz
D0UGrc2U/yKrD5WbOnENSzBLgGJPTSL2VXgcdR1nK55nTNJHi1Hcxm7NKNQ1DqdU
eba3e2DvoAsRjX8aW60JSaFEIOW4gpP09joMIybC3HRFxywZBhdhFC+2YjP3mOAQ
3V14Zco6AgsK1403438Y9xk/umFKxvuawBsUU+xK8sauYpv53jV7pG7tExX2CjzM
4eDhz/gHL71lM54CWj6E/+bMdiQCfm0LNEPQp6c9uJcVz/e3pGhYBcRlpK+99Bux
xDobCt3ZlgWVsNNVWv9/tLIF/3zZQwx6tligfEn8JNdMQTxgHHbUpk2XCE+hS9jb
TQ/Fc0S0t56tYoPf/QvYrLYpUrHuzjT38wa3Z6BLdYymk2HkpwxX4SgM0pJeyzhc
iDjYRfwOJYIXPL0Xdy7ELJ4lSVM7ctEjeXoCpOUpLJBfVkpaEKEjzQOvPLcm9T5F
OAknUAFsyKugp94Aa2aUrkj2mtSCYa0V1dGnH6ygbVFhRAIkUlkeq6Jq3jCSsgR6
AWhTYsC3a1MMk+gqnbbX4kfYqLeNaUq8YFI1suZBmw1mEKkKXxaDDSjI+eGChYh5
IEC436yQ7eGbIJwu3CvQzFKuTwLpIJrqLSAw4grMNWseLBW4tjExs/06wVISE+DG
7fLczLLmRGoVBgnqHytgIQmz52Bg2NI+nwciqiIXxRn9/FwKsF+lmG4eBl5OUqbe
uC7DgUhqL4hqf8bLvALHFHsVq7TQ09Akj32csWyd5szNQJykVc53aesj78Q/xHLe
ifioSo1GY0x8r6GpF5qoE+O/B2w84F/5QVZG5shm+dYrMcs3MpThGEO1PK0hqQVU
YxC8s7T+xZWh+5MgyXAIfpCUI4iiCP6hnosq5U5fH6KjQMcqEUG7suf1hgEukBCH
l/BpbKsr30FEPrnoicfvWwNeChl6RY2wPkDP1VQz/2nP3j3w8Z6az3NEuQTr60vV
1THzPjN84hcORKteUqyLL48IhvuIFLzqzyev0PLxT56SH3o4BCsPvUIGOhCGA+L8
XY1uZS7EUPthe81/DFeixgYl38MiUzTt/C1knartTxz/gif5w60i3QzjQMmYqWo8
Q8cnyiCxz26U6jDDo4mNiPNkLntEPWGpKoSrziA6rv8ojbh21Mvy5fFN7qm7tgAz
WBsIMZVsI0IkpulKONY7cldODFKh0M4Mj5CQr3MCR46yEIMRJucqJFDJdDirRImN
Zl6Hdi3Vz3I73zvgscu0Tj04K1IzRs+c7o4Ydwz32MsVPT09jdwsSi3qwOvJuliy
YsB17JbMPWOmvrfN2Oo05ydzKCa6LIYv+Uv/jE1/yfr99fo1THDR1I35+XVgrv7A
TtzhTsHKksL7UdIi0cI9M4OIOYwYGmo6UlIQgzB10jI2XTXgpYwN0ipFLlOtR7CT
6wVa+VB9gOjZWkybxxbVfezRsb58ObBUAzGQxYD37aXTExnacGiKR2zRADVKtQks
jIrTQL3jpaqW3nx3S/yT8133ab8cSwGZaQHLHCPBKDXnc6jbZ7RYBtZoQygK7ggn
FopIums5t8pRA1n/ww+cqUpe3ODQIknxbDegLRJtBJcBrk/RCFbLzFHZPDGljxlC
ESK05+36wu/8TQAC0dE4UCYlTCe+nGPnHCXVH4aVY4g4pKD0Sc4bORwnD/9wVFvb
wNCzBjZjqnYpRYppplmML12VgFGaw/FzF9L6VShTm2Cen4J/oRRoAUJl0PrFEGSa
jy2S0Wrqsl3UyZXjOw1cFIgHRHJ+Ep3kyO0Y4vbxaVWOTLAZBElADqkCbagrt28m
Y9GO5Jkq0PqhKop+dDt3oPyjrvcdMkBU29zUf8pH/c8Fu5vuZQ0TMYJUdqb24P+E
iBETeVGQIY4BoO0T4n22Wt3A78Tqe/vB9eneE3LDScxuuXZto+T/e6uZkrWEX1kB
U4em9bpEFlSsJbqFXRs4C7yvKJaoCs8PVZ76I8SBLo3kPmEsRMzEWN9kLvrwcgwY
9NQ8BJUpwgmYX1s1rb8gcJc+bIc4HLctL77tpEgQYmo84g0wR/587W3q/vKDY3BU
Xfj6X/bJwcBsI8mhots+CDLTlC9wORUlO/flQJ0lFyVNfMk13OYqMTrNUAHHvsP4
/k59uSWv24NctaKcoSvCGpzf/9llBlH13Y74jgwJ6q50IVIiNRA6ArU7XWjNA4Hy
6w8zt6GtWmKj5wlq7ODTNFyUh3p9YWf4Y9qcKA4h6tX0QJXHuV/7OF2M+ttUBuCK
jxqaBIaMuVMN6jDkquY8TWiXajKPV9v9GC9lCqwWRUJKcTbZAyQwZEWzXlnopCZK
0evB8JfnTh3t8NjbOs2LnDDfswfom4NH8I5rHXVl8AG/LtdY9VflcsDoeAcFkjS3
mZjnN0BdIpF0U5hfNdERNwtqgCwdGWSVK4+YXvFqnCNFVtG3oqTAhwxzL2uIoPjw
5z3uL/gFNqpELYMqTLBuN0denAbEIB63by1S4ZHuutCDIAdtQNXliSXsVgvvlN0X
Vpl8pQeGq36AVrGHBjrLZ2rMD+qLoo+OPsHtD1/peMdg1b2SSVVOQ1VzvcIIg/ZU
bmvN3Z1GGfRBdHdq9c6b3PzeRQwXyYlZy8UB4g30dXBzb31kbsaVMvwbwbBgxIZZ
6hN0PAMsEBW94nVvey+MQIy5MzXqWPP9X0FvYm+k1DDLS78lyBeV//tG6eVhtSlU
oAqJ4Od57H5xaS2J8asPSGEdJ4vshiWOdlbxxnWvuhvAPpqc9fcrsQHY0EgITjVd
NgZOnMJjYLMaLg9KMPC32mZM0hGVuNcdjG7DHMKxwQR5pgJg9Y4HpyAEbTQKRepn
YtYevjVwff3rh1ZWDFEgkBGMq74c7V2kEcC7rJDm6y4FpywrQv0Iig33A/SI1mF/
/oAdMXOu03QEzhOKTx/w1IEt8623qbZhikZl7FWW6tu9gSdxlUb25O8sRzwi0SB9
u+zdC6a8xyk2l34mSZlEcUEOqUiIGfwo+h0ut6aeNuS1DwCvdHKtfnD8xGjfJSk2
n+lUXy7O49qvZGB6c2nRFVnej9VpBy1jybsJ898ixetAOS4oYwmZ6aTDXZfL75ld
20yu04k+ChrFA+aot3cyHPdai1b1C/s3pfuUg7XgiOit8RY/vjwnqvxvZfLM3xoa
M15R+VjdWVbAbe0VrUFBJIL6/v/79oFcQlIPR6aIBV/XmfRxQ6ec39QGg4pAD9ox
a5iT860KyUS/O1/NiiEM2diS98u8N9HhNGTMEccIpviipDzR14cTwart0hGxvD2a
nE0C0zFzQlgrcJqKUiTZpohkpMSxc331tHxoAQlVwbrYRcAlYWLcaxsXapChbf20
k5szNxpujP0fGncWz1DmjRtSnFVDVauldUzN4H12i0SFw9FLgF4akCc5NfOkex0m
wS7vBfSUax66xMuEMcNT41Cez7ly+aawTNODL+2WsfXvePn5IefCSPOEWXZpC8eZ
MyZaRlVTEqagLzS9o2Aa2UCXaNDG8j/QCVOb8m4lCUTpUR/6RH1xrx1Q4qvpg/M7
h3T9S3nFSV3HFpHwXO6FFgLyV6nen2H9oKRzYGsLJhlYzKEOKJmJRtXH4dcKmUYB
FDBQR77IQ75NJlfuAK2LeGinqM6Zj8m80mVFOjJH2DtESNXP4eWhE4EhphFipiRC
PzhlpATMl7P3VOH6kl4pLgorCwSDfGgnikcefhCY6tfHbYiy7rjzg9VSRheSEAkT
+ld1oI/B0yR3pxe23964A61zMnvkqs04yf0GVRMBL03B/RWQ/lRYAIOAPHfycngG
hGGNIjPCRfN5FcMSkT2njGzblceewZqYPthqWDwVs96l/b8XlwXiNJZzpoypB9W9
uVcxinWwhiqWwx7ZXN4qfX1ilf94lAlBQyvCFzgvBm21CErdtbz7Skv2i6R6vAuK
0yTzSGDW4BOeEc0u8LSy2LRBT6QANve9+qTi3NcAWz/tegER3gyi/7UfTG2sLBt9
AZrnqffM6+UQce0/m89W+ooEK05pWhyeEVE+y3LafQ8yzXG5diXPI3bDix4OWvms
QZVSUcK9YAI5VKN10IXI9VwUkdKqrUFM9q/CBoxG2YXEHBLsFBNUX5jrMInWP0ha
UpnQOoTtsERET36gQw6E7ZpML3vvaMRDAk5OcWel4ROOA1dR7h6mR6PqzjxKuNTf
OILsDhgfSjCnqEAFIlBT2k13o7qjQuJPIlbvr5wyJF53mff0C3Uxk+isitwNXf+z
sN7tl+5ojLVPEVify8JraJHvyp1H0Ir35dJZLhMpK8PhbAcMc5mUaFOth9P1wf7J
Yif00KJV/tCvjYJTcGe21jBEqddWV3E0QnivgnTPxGk929voyqZGFo0mYulVihHx
kt6ajmYGGBCSmp8/G/53G15JW+Im5TqUHcE+YNmhzI+DWesiaz7PqnmnvAC12L3t
NvcdqfR7k+oznUDEg/MBcFqcC0bQRnyymprGy/xI55K+w5z1Kt/ZuhnyFrFkIPJm
eTpDCSnXMTnKK3gtvwspo4Oa0L+Q3ENC2cfTZSC4ACZgEO7pNHP8DOQr0htdBYPO
BqsHwY2X0PmxvtyM5PzU5GRfszi7fi75EbmEha/cZgAFAevfYxZ5v4rECCtu5efO
JWG6HxhZ3/kY2WgVSnVniCGTUgvSxBFf/PlpsxQY+fVt7QsHKpCOvFfDv4TNqmKp
MMiFoVICyVgyarOT7TRvDXFr9rpAovrg0g9Scjq7kcOQ5t3pGMsUg7OEQQmOOBw+
p4ntgnzPlOef5F90ga/i0TH5Jn011yjRAGqf8FaN6c+cxvDynYs6+Cmf04zfvQ0d
pf4DSQ/sAK2bn0tU7jal4bQdRy6BUUFbF2U84pOA0ilMTH0AbwY/RRUHvu30pxlk
nkJqt4TBSbkVOhC/5lg3eF2jmXSslmn4sVwtNwh9p2UgNNZxrt+J5vtPBoZMO7b4
JaHMnPznkKbu1EsNv3SZu11i2Bg6X7SihEbf2RCXntMYU0q6SrXCfibdLKi1Kgne
SfYTCXq+ZKuElJrvclQIkmUjgbKJ/r6Y843aDgePWa2lqQmUCkG8GbeoyrPFFXt/
mCDLfS/GeQEQx/+eqYQC0Uc/B5uG+eaTAmRapmJC9x3DDQ/sIotp80rfr5G9YuvJ
cfa4z1PxQWlgMh6cu6fzxMLZr7z7Yp8uCnr4SUXLt1zQI4fhIpXVlGbVO8KH1DDY
thCA0FP0N8M5RPTyQd3h96t8mKpRhrPkoZNOuDbUKSrmkwUKZ8Cdrs+W5gMVUQcr
r6BwRTUrQjdkvsY8hJ1MOAM8Uhhf7JZi5Q+qGKkPI3YtrYsGyeAcJcxFCqJiMcyl
3zFy3LpFRWsSV5kLXeL3otzHM/WPCEwRd9MGqCEP53d0Mgw/IBpl29LdoEfgW3zc
CA3OpcMOsb1NnTBAbQDcVja8TNtDi2U3wu3FJ2qJZU2ObBfrHIQ8mLWdlbSq7uHg
mEIijA0/q9nuq/FL231+aNsQ8iT4miGBGU7YrRBZ/HGuMqSGFtaYHT6XMEqhhG+Z
/JWUBGYkwnQaf8tlpMe5+AORG7nLymVW0y3mizr9CKSOlWjQG3mFf2tKBxLoVzYy
gX3EOGA4uO+dyi6GeLGk2tWocrU0rQBhaVvFCIRqq+V2SPDt9GpKrHWG3YsaIxUp
bJ74ImhOLY9JKGIZxf/vbcTxMcSAaiEbEi2hFse/o+rKDBvFr9uqSVbbRHb3fG0l
9fx20Uh+vhRGafHMw2EoRv8GVw7FnhteGvTD7W3KHqgH3V6NNE99R+vrIZ16tTk2
c5tYETf0GCo6nqSAM1A2iZmdfe9o+ykmbl83k3xi5Y+qYIC3qYUH+FdEaGDg6pWc
Hb3O0ttkPbzxyGzbo+Am6h/nwfCzd1IOsn1RFJpERJM+LwqE+fNMaDbiSI0/Cpi3
rF9AbcWjRWutV+YEUjXQfjkV1LkRn9hHEhwm6Sn55lxpESOxQBuEgK6NACrxqeys
6zWondI5huAIbL2AHjImxVHq/DF3WADbwLYb1NoVb+tT553gqfQi1JWes/6JZeEX
cvK4y2TehNepa4vTxp9/AV0ddjk16tgtIuvXpi2L5PAUYLtNYcB/DbWnn99nVHgC
jcyv47jB9wMqK4yfUOqo3CXQp7S52UIFPQCPTs1LsNmOTuR2Q96yXnjmodt/ywdJ
G6VNYl60ib/Qq84nyo2d6aI3oy1hfblKJlL1vCNvuXjB1f7SlCWDX6LNh0xjexk5
8YeYYo2mDi9S1gD6a+rpRC6eXFwgCgzzTZsw1/NYNBieqCFKuI9F1rBphFZHnFJC
AzHSXfbtNq2YwFgBTwSsTGzMylNLu1c3WTn9rpXuGUvC8cxcysnbMFLGuLOQON/O
FYkN3PyAb9fuJghlwRHlzCMsiiYDVYXTgt8dmyafVvJoA0DEDzh9DTdOEObuVE+H
ebyGLBMMnJweg8aH4Sl6ybAE4oR1FBlfgyka7nEukGy5V9nLBlWQhwt4Ebeviu1a
/teItjnoL3xFuf8eC4f+LNE71zUPgHWUwQ6l+B4eM03qM65H+SCTFrXLDkc2/mhv
BfAAv/jeTtApFdcrEMh/AZmuhvJhpVCQDTIAcKHl72/1iz5K6B3Qw8qRtqsz6TrW
FE+aOsj7uGOZ05v2Q52/dhdcC/NY4qTHrNRm3IHNrNre747C7SXpNxu7nc2bM7OX
5517zCJXSA5QXdXLgeHzRpJjcGqSCaWJKRYYc1OL3uRcjchvtqzRN/joIUs3AkUh
cHVt49/NcawhRSAvSoH7k0XebCTxjDBtQ5r/L0K5B2LyvuqLFPWoXIfR5aFU4Sy2
iW6bq/fpFGXDG2OPU4dCGk2TfbOMHeI8TlE+WPbWDZ1YXqypIUxbkEWLWealLbnG
6ogf2tgNXP6Y78TSLyOxDWs20RjQxaCCJM/+QawVNzdJq4zncaLDxqIDZr0/U8F8
N9JvSdAxVHmZqqIoHvVXvyKUn3L7BIZyEeD+RqXFG5K2ipJW0d46ViBc4QSKNIy2
hNv8jpheqz82siH/mdPzoToYIrckuc/ErMkZ+5HThCsrSy996f+X3VAQq7mpd7FO
CtSDiBJBWqKkvhYpGrSjb3+RvcJzYk7/jEaUmk3SPE1kfwHn54HYgzEAo0V6imWi
MlpsCK5Qf2ySzQ0vUD2U3QESVbWEgtP9vcmXcUfYh3NafL4SfS+Yq00lUf0MJmci
+IEQ3iQeULAYUiVlUBWtQy+jQG1WSAiVLVl3IcEZa8h0k7tHb7f4zUEbBjfidVWm
/D4MMTnY+BJ2EBhP3EN09E7FeD04nu86u/8Q8xfrXOjaSUptS9MAdG9HFAFPnyrB
v1l8AATcyVsMKo4NZ9/py03z5BKU/UZnVU/hm9dnzCwGCQQVaU6UJQrMHo/BLpSM
c6n9PI8SiHrIOq4ch9VAyPSsdQSYLifIHpK4KChytewaDiGSzLVxmyCB+EmvfODa
dqohnnl4Hvkt9Vk3TsB7bsGZmKe0QBKGtYMvs/PZNaEYYlsJ6eXPz+xS6QmsX7/w
I4aEz3i4z74Qpohd5M7ewq9drVeEzHiUs8TklPYdlrN+OYlfghECCIPriN1GIDez
f+Z9+6yXSI8Qhq1pZbYxUWAu+03Vc/Ywn14UZvWV7lr/A0ADUQaj+ZsJQRYuZBUh
+qpwYgz78Xc4NGvSQXTeCkV3mtb6rDSYHlN0L9Zab3I94/DImf0N7b477pKAsztb
tSCb/GhIn7Wc/MnkGNOiQnAu2hcu3b8rtUCYHFzmf1hJP2GOD3P33L/KCM8Se3sk
MmmdeJAVyzyAe2WgYSF38QcSFS7WeeFh3kt1go2tC21YWMn1LMykiwYWlNtZPH7j
1MxvPTAp91gIEC2VFKEgrymwK5FRRyKDBOfp1KTgXYlxbRpm3rLoAVZr5LkeSaMb
u0pS05MeW/YRlD4dlcuSPzEBQ36FBXsQmcEbyaLoo4prmhBz9EIOaZIerYtTHPrN
dBqUrrK6hn9iGTVtEKrDgo4kPrEXP9YoXEhLgc4rLYnVXm1aeqRfnFHDqio6+HgB
3t1OfHHZ+7aHXiHDzgrIFng+6u1eX4fdce7B1Wtlq10Z4juiJ8DJOPxzu5dBn9Nu
408LkTdJytlEvHgbmrBTa48bpYPubsV07LZxcPV0k9JdVWF3BVMBUzM9pbP9YF6g
qu0co02d50t/zELJlxCQBeYM/ybkJnZuNFKlnHTgDx+zFFSLLadkOv/+M7S+yrR+
/Lgs+B01CocYrYPWbKT7NmZ6limMzRypZhDmTEo3ZDr9DSeX94oQMxeojZfxHfsD
QUphepT70pNiZ1vXgmpJY1STeAEqFIPUzqOt4s3BHnvXLL/LMO8HhOVcs8sTkT8x
09awwOTQteA6tN47YZJH5bHCR3/qQrPdqTwczTUnuHa/jsLsBUld0oBr2ndWpvQz
2qlgPu8u34MIstifWbV87Qgi/f87K0SXVDIVtOF7MUgYC3wnLJcU3C6kA2ZPZ92D
mgj+KZ5t65VXe0QYe2xWNzu2YWB9nn65gEwIEXKrhu//3m4kWZxJSr+Ff3fGtBWn
MBfjLm+rkOuzyQNWVymUU2J+j4F0ccdlSTVSvriQjqgpalsMIb0/RL0MXvMOakx6
3puokpPIfSe2HFER/RFqZfERl46plL2x35YjLSwY/ZVegAzsB9hkoheiCOFhS6SC
eewPAApgz/3HLLgoQCHl6tExT4+qkhI4rBOmZBmUHRnR2IerqtguKDaAS9Vr1iAd
Wyf8LolXuEs8UQtKq39TUnL+fe3K1hhLZI0ydMZMLT0totYomCv+TvZ+NzjYD9Di
Z1AWv1f7Y2Q3owOK72lEi4d4itPPan9TKRGuIrpKiEiyn9pmV1J655fsN6t47mHr
uxyVaN3cY2FfJ/7iixpFYUyQT4aUCoI0hMIiW90G1i7DjhQGZtHKLKzzxv8eJt8m
ZsmEIf9CltqtQfP9z45p1Ei2FdKpHwe8tSkYCEvcGOdHSifwA37zS2c/qIgvvv/T
0eG1t3ZMcagiSGy7VhnX62+5Ax8HL8heDuiSMsB1E3D29uan/Chh8iLts9XTF53A
yyMEBuulRt1DHR7h/jqHgdWFHrFlBNNmTKecWMZTwDc0DxTd9CvZ+rXuNK6yQawN
BIGL1w4cTKmpHYjKBeS7qME9AWCBHvjuHU4IfBgemoZE+OdooBlhCRzShn2qBE4q
r1JbGVlMu+zEUHjlrlPrEYbEOmzEEghKCnMUzYcZLQEm2J1AYTR7zC90F+fklUQT
a3I7V637YaVBK599GTfEJQ5jl8WaZhrEYK8joc83PoW/v5t47ReMh10kUPUmCCWj
Y9z98dmIWLh6V2mHHGmN4RhTD1imgfqwuVSWNeHFZMyhOZY2eR7vrj1VIoGPAslF
LGwILSO8c4IBinaClFeIzjslGrMm1PnEesbun5DIp44EZ1kXhFGaucdIZxgniAZe
479xlvAIR9CE3IO86b2ImGnkogKl8cO7T8EZK2UBztATic4IycjUJfuheFC/OQOv
P+BfFkZxaxWynKkYoc4WpSspn1I00RoroQVJTMHzIanUz8x4BxzcafmFOZkpLnMS
6fDjh4sjeQw2YQsUG8EzmT1N0bH81gHOFMxWCDGp+hCRK4KsshyUa9LuL/NCm6aM
M2jHzPuWy/YwI4daV8sb1EqZqOJEcB7eDNoMbmbw1b0jEa1lZPh1SwjeN26G77lP
M8mQiSYTHqDbd+hE2HOmE7tPCRBvizS+Cu0qqLz/QF7AJLvdthQ3gG4FHL//aVBc
2qNsVkWZAFhQ62ykYzlHKUycDuiP9ymOiQ41ZpeQyJu4gsaIhtc7o7Tfyvdm+7vY
qQwKDeZbazLxZGmiJN5gRHGn/JEi31WeUeVniGMa7wAq/m3RWJnE9p/gwDFI2g4f
jr3tx8A20tlGkLuNbfbfFzjDNT6y6LU4/EamhzSeAVzZWDmBksm1crIBXXWzNJru
`protect END_PROTECTED
