`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VlwbtVY/nc0rqEIR73QdBerrzgBL3dRWKbqzZURf4Gv01mRc95BmSxaci5GtbOCJ
YY6wm39tUKmkHeFmXMPSqXBFFMCRHuTtZFtBdDTsjlKLfj4ycGjJ6KSXZg/D+VGk
CsnROJHf3tuIsV6Z58cwBYtWaieAonXO9BZAS0huvDP/DHbk96hlANGAs2fFkCaz
uLnkthFEcQGkfuspQHg/FZRkgEol8oAEVv5QO3PrTBeONQKXaS/FtSXg2mV6X+vR
yVRPj2ERbFOPDuRsxZcLmmUJDCsgKIymC1ofznMCJr6lQaFh/Y+sep/isuokcFX+
iSRAeHcqfZaKD9ZU/YPDxPpz6F9fsfC4bZtbmyAKcUw38rkrI/tKoB/rqYmn6xrp
pqmWu2FQusrQ3XeQIVq/LHq2EARCUgOOd5G0uCKEpe7AFB6ggFRic9uJZdUeCvWO
/VeZ6GSaVIhv66Y6VhmBDndCRwLwSinqBx6+atRxaFPUVktkratOMCjAma/KIHwT
DEeHRsHfEgPskulba3PyVZvflRPOSmGOpQgKApNG0RMu/eLTKNoGEDM4wdwbAUPJ
ElIYKMRS6TXeY3dopT6Ixgc5ntAXsnrlC+QbZA4qxxSh+RNQC0egamgJXRzc37Th
o08ZtQOMp3kHORSHerimUSDdBGwC4ouPAKlzQrX0U6XZqS4c9Q/vx1ksc3PUlnYM
0YFKe7cZwzIsiZd0ESM12XMVqf6azbAaeHSdiKDpA5L3m+znv5YVM+xnFeVb87lK
vIkY81ylxZ57bjyal7gvSPXvKz4/KR5WxbfdAaMCFCkEMgvtQW6pr+qC4kxrqNGf
/WfrKFxYKy1nH2Hirs3z4zwgy+DZpSOF+vkfIIKCWKSlws5xjglfmZgnocwxPsWz
atyiTJOO1MEyf8PQkHLrV7BaS+JCIvBB5nlsHsaJlhMSTAmojPlgIk7Zbds7mZYd
cjV8cljxuGritraFL4k4ixfSs0ZDIToKlSiGjrscfFgFFZU9k0zTx47I2cmW0lxJ
fDW9EFACFxfKM5xFvSHvFPxZKS7B+70JHgtbZkx686/527eMDFMeg+UkWjMXbhxK
F2vuJAgEsTUVzvCyX6ZAhA4Mf4j7Fl0o6ym0HnL6scbQgXA9chcUXazUH1tI9EJ0
/Bm/yg3GpR1r/kqrYmbzcOu5DDULR1FQzjpxn2HsGvfjdS1bpjDTRoOirkp5VDW/
zRh/WytDesv774qoo8S6vl0BUzM3yS5FX0NIb7HCzFMuu5s/m/iFBh/lnBi3l7+C
rJR+QpJle2ZmtqpCgAbxdVkQgquMFBo5G8s+sXRLFMbfbsdqVpY+5pblbkXxizdJ
AegvaGs+q9fo3o84WuCz326SVuEasypwSnPbp4V51i8muxxeFhqa6XFe9HgAwSzI
VBAjRD+iSOBa6nwaQHD76sJTF6G1gj381z0+NAVXTca4AJmwNlgTbU3w+Lkkd0XM
HhRPAm2LzTq6EjT3rM191VslsskqRbfemM32J+H6ghiZ+PDaTG6HHzhxOEtfBTNx
FF3NGfNXn5qbrJrY48qDeuryEShoE3V+LlHnsieglrFwpTVQ9+HsBuUKzHSwdbe/
ECAHeg3JrBzw7CVHaDF5XqTZuShOiC4jvSOkI0uo7FtypRD2A0BrEIpfiYjwVSzN
CqtWYAsDnTJ9qQdKy6zkqmndUU8dzA4WyluK/Vss9miN88MfeKTlBsOafFhVxMQp
D3xBQOW3l39ZJ7Mxm+snTJPHmRA5L+aUWse+SlVAFcn9vgbwiNmIbTWG1kCL9Str
T7BLkYrNJi+vxOWnuACBzhxKQ55plp8y5DyD5gPyAqGmqLU/FLttOF58V2aocdJW
V2BqPmTAsxbNLnUG6zU+LlrqFISub7rX10FSmT57sFuZfAOD4w6+SepafLZ6a3rT
lCSqDbFBPBt8hyYkRG9GU3Fz7+Z4VJS1I5XrCAzrzRd1+1V4RfLU35Raz5GIuwkW
5MMsJwqQjg+qL+YQLQdmefZB/PytCtnO2Te6KTYWar9krqY1C4CJI06P0Vyw0Zly
QLQ+PPiGsOL2VewHZyFNVxK3FbONH9dVDX1A2F6620d0E/Yoa+uMDFSy9DYtLJWI
41GOYS9gqyzk9JXTqEI1xzedldmpYZWs9cCU+mI61Wo+v3cBBwW8TuI7Gaw3otuA
cK3AyKyxdj4vy7dthPQJhQyd5ebZvpJyfGnaPPXYocanPcYQjuzjak0cunFHlW44
VEZxPPxdN5cBnC/Nx0VwTu3zBAvpbVEMLPTuHkGlwi8ZwEgTWHi2dYsGJrgzeXrA
U70DaMJGDHk4NHruovvf9as/x7Ecips0znNmNtz+kyvsZ0KjRU/yqtInMeErnJRe
pBwpWz6+Qppo8qvkoBf8ZBjSn9DWkJM8GCep5QkU+QiD5GUNCssnoVaKTIVVyPm6
MQfFjDY9tAHNi2UOANwpSegrJUb3JN6CwqQ0gElY5N94j88RBQ7q2eWUqxYP2eo4
WpGPrLUGQoQIIJZENTAGhoxERcr9HRVuBXmqvRA2d4iSiJUPfLcNppO7ZxsKwA+L
JOsqviTfzR0fdcWBybajg0hGjn/y6u3j6vlh1rDaQ8NjeahTAjJ6RyusNDKSlgqe
FhHdoyZnci9KTPEguH8J8XgkH1hP0ekKcLKE5IpyqRkbAWov5dxgaxAxDwQDoq0M
FNFHljdn/yQoIwhHLlRsbdKgYDZ/kSzf8Uw5YPNcZc5YM8uDfNogtsuiJHX3x6+E
kuF2scEg0dmclpCTEZYzbrzuXzh63EeVQ/Nvzn6N/xNoaN9HCkHZX6rnmrX9SRJq
JBPC4WqOmjSPHIRbGtNliwX/YKHgBc0J2eGB1KRsYRqDfPPF/t6lW/T9Exr9pNk/
yx0MBdUmNJz/u7aVSMHFXdand5HhTBB5kZ7bCV+LdJyqM9JDqJZz61YOgMXpo9eb
Mq1YKfWcIrKGtyBNLvtMfvBLelUDUwEbjq7mAy4TAQQIoqfzPM114YSw+PbnlVbq
8VRrlLgs7jkUhiq7dplRlwl5PeVQeO62WMMoBCeM4P2WUmbwSQw1hqNE3srTZkbZ
W7RfDzi4ssPSbxfoQN2EKoIGW+piERYU4j0bogLUOjxcDXAOX5bA2nv+59GRTXDH
zbmoB3XOPoLpAD+ta/YaN6Hh/z81d21k0xhK/RPw7XfYOdBaowu85v0CAb5JZ0cn
kztqKYmdmhBi4nV3IUD8fM1O62wz8U7Uu0B76FchgzukvrUzjfLtVhiG/dcRtl47
ni0Bupc6hJijcwmr2wlpS+ZYn1Hf5cucmtr7KgFOwaJlkYE4sCZmrqfQ78zU8/l5
gVdVV9JTCgjpFQhpWolFwEeMWk78NwSYzL2CZ/CgBSxqLAJ7hlz2Wbq/en6H7F4g
3B4gPtPSjlgmwE+x6p3NLdzddfe/WfEeqk6GfKAYX+ytzC/LQbAn2W+o1gho9q2k
Mm2KV8rZeHPJNqm/CQa25Yjq/WnsoNzSJt2zDoKg9Beban6xOQM5T5P0sKqnGbFo
+9u3H/wQMfg/y6P0thTbWlH+W9QXh+XMBOu50+pOriLm30H5e5JD6qnA68OYmWfZ
AItzAr01/+fypcC5Li9nXtx5+Dvs0usrwyHDv0IA76TnsRlwQ5R1KrUPEpfyJNjD
zXtsnDOOBxKImFf9hXKnqrg6lXJdbaUj2BKneSZVC1nXiTBAO9rlnoz3OskhJYyt
r7R+FsLGKoJBdmpUn9ybvT4TgC0s/7CkPaUYDU99ubSuhHj7y7rNknwDcftbFbGe
m5IoXi0T88+vXbDsMIhHbqST4ugCYRWRH/q8xDoK2EvTwkwar9Ij7eeYVtWNgr6C
sWFCq7rYLorrSA60ZiQQ+HVRC/47wP4hdMXmqmPCdHoraklNTdKDtkKyxj9vceWB
svUeewOMm6U/EPndfo53EGYqlL2hB8sjHM0lirAjOOi3AzrgJuWy57JDUbi8QNhw
nKP2thtWOBubmEMdlvL6kGF78FH2n+QmupVO0as8NvC9sIyu3044gS733xf29eyT
g1C4ra10O8LGJGDTgFDvYTKqSBmWEjipI3ZNLbXOkbuke2J6z+aJ/xhJGtAGv8Aw
/HlRq/JHO0QXM4Q/W7vKw2McKx1jYEA9I+MxWg3GUlI/pCjEbnjyEpxN6og1tNwr
oRA0ltZrpteSIdKbG8SjWHJSGNh9bQk8JK6EDKrUtrEm2CGHrkVM1RurUdbYiVf6
tORoYVbGqSL48r6FjRuNGtnijXcBCmn/WiP4wMZVYlnuTFQnTur1F/55D+jCbVhK
HN74BWADzdA7qlo/oL3ui4YZifu7h4/osq+F99LyGHAHxByKSpir3tvW5fkub/kY
n5vU3+En99QNLXzURYcCARDD/+V5VQxzxWwQkZnIbUPnVc4VGxq3FV192DT9kWG6
6z+DbPtjJaHqao1eSpeakmR+RsewPC29gCqHh9ueMeKvYqRBO15Wa+0ykjvP6YiM
66iZbp1o0tdDVahiricisjZGkuhV8lxjpEiJb55OyIpZ5S9hDbtb3yurBbQ3Skqd
cXrLS6gK9NbY/dutuhhLKDGaKs/MPf+HoofiiXX96jIU+wB2+LM5RDC7YSneDv6F
mTP5y5biC/qPITnmqcshdi3h7t0hNzQ63RM6nwSygCR7mu6hzrvLwFcSozm71V4u
TSgIHl+Ds+l4TqQj3Ku4+hL2xOMMtJNp3PyMT0MkPCXPLdnFKq8qs+xKotLBZPGq
SdAv13lKajo8JEV+Bq3X26XMQr8AP6UDef+lAFW7BbN7Pk2CoCETyMdK2t7fYUx/
566muoReViPoYCxNmj8xdkmAIJs7R/+6n/8UYC6yQeP2JZ9jdIlkDuK4trEpEhUi
+QvhJpBuofw3ycNeqtRRC0yjYMQ4HWr3wJ6hbXYp6PGF+4fKwxyHIP56dWGA6mk4
10yC3PAHaU3mnf4KX96bGK27mOQqGXZVowox+23HVi7or2eOtkcq8hRVHm5SPLZ7
F5i9evta8Pg1x47+CuiwhI9DBKeHDDiUeLjo3XB1LxE/9xRDFswqNaTmtnrzc8in
KvPDh0pz+jFYFOoIzPwX0J2akLfnzSGRXG8lUGwnPMDQTFvz9OT57fN7Ekj2u8S6
K1x4DQfw2UvJjWUdc5xgPr+3sfQn1aNRu1MQQgv+qOnoI6WQdeKXPTjYni9PcPEk
/QMMCh9gD0gKeJWOj10Iyf5RjFNAEp5HFogbXhdCID59eyGCTfTU2mZrvD5eJJHV
Bd07rRYuXYXwPH1MxL9EZmwV1y8v4ufvIvVku1A+GudVSNdoxPDzOg2qJWHz0Tf1
jF0J21F1ROPgDTkaZFV41SKQd8M9Br/2ETl1WXEd5/arogXtLlA5GeZ2lbgLtqIs
egQeyX8FDk3IRh/QJUFPdbIsTE/6DYttfFjP02ZAZoVlulT3sCqZ7+OvgC0TiUy6
2nK4MJtrg1zTW21V9NWuYWLU+HDEu1RljWHDuiELz6s5m2fRfGYF6gxK0m5JJ+Vp
NGLtKmP1MzV0pMHX5fwJf6HqkRufC8mVf/OStj2yLhDceuQuhKj2JwiLBwoxSVih
0hMFQyfMRotfKW03mNi2rOWGN2ZHiLjibJWdiFT8/r/qGL5Nco6PCugGYbFnYs+3
ocOJAXbDeWa15Jg+Q1v/8J3ndiuhooo4uBd6cau4XTJuyJsjUbMCZmq/Y8vI3cCx
K6knf9sBp4dcQ/WN7lVwonpmSdOmRCYVU9kJA/g1X6zFdk8rE2Qn7ec+GTJQoUxd
nq/DsRWF7ROuK1+3WZHAiKdCtjBWCWxX107/0jfuiVQQr9R2OX4ZZb5z2pzqS4o1
JOeP+bAwX65/1Mq7pZvW8IX3OO3Nh5hwjOIRfe5OjXZ5ukK1BLsbws3at+KxDXJX
8JFrqWlW2n52Q1yGB33fI3Zngt89vtgCRAK0e6uAEIcSP20T3gjJffX5HXY6WTGL
lfvhS5Go9ZUDVYIpnewiR3eKeB6IZoOyVSWd0YqPYaVJp5yR1lGmARsyPr+NSrPX
k/VatCmPzpJuQS1zHCYPIa/LWUqv17L8xFZ55b2ujw/AQMjhXj4zKeB4sPZIy24X
t9qFjelVk4GT+nXAIy5ThiGGDWxHUmHW5Zfi/9r00NVSI1pOiWIAyFLVU6z5lVAD
r9iUDRRaYcJSJCpxora9OMmLgp7VHUjBMEX0uu87F5u4YREXNjNIoOtZimcnjcsk
aspvv5xw8WaKGhsI1iUJtb32BlFz2Oi6edR3UXeSEASUZdwv2iVjnMZloA6RFDCf
fvG9lkK9DHtP6RxaFHZusJ7ikKeYzh/GyLTdDT7/znCLr8BQ1B/ksHkjsTj5aRlp
pqxMPerfaKKgZM4neFXRyfrPmLc7rgLx6xU+tNTWRk64V2/zHPCvDO1yhG49Q4n4
xe32NrXZFssowvXXbB7ZWBVxEOHtrPGvCjFxqeMz1aqZXr2DjEuiGsXgRwdliqML
qFZbBu4DByr6mKsA6FFnVpJLqAOLX0QPB9cqh6YhH58x+EO2leZP1g9VZjGuyGL1
Of+uMlipSvQbYVoy2r/cIW0z1BdhawBfkHNWk34vE5MWLxCqewidPyDzcwR4Z1sm
av8lKh/EEC5aCxhFQ76IRm9KWjp66VC6SzXk5xXoCSa3+uM+ufRD6e0qT+USXXtJ
ea4RcSBSWMdxe2aFuAUzazJPYPjt11zfSO+B4yfbSnM3CVA+85CYL+IDGm8hsyEj
wOeE4R8/2VZJfXHGlvgoEQnBfmIzHHbVXiw4F4dEtc8gGxArV9t26SQW9TS1RbJ3
phjqS/UdYHDZcwK/fhh0vMADBeZFAbQRLpLlgBaLM6a5W589+rm7KFXncgOm2XAc
i7WjJpHD0nP6lE3T9NSUfYN4WO9hxZK7bHN+gjUqp5mAerMKYH7OdAsFRy4Fb6iu
sDhQeq64ZbUHp0haqWfO42oLhUw8TRCeCE2nYllUuLz7nVfwfth6btfwag+b++aC
kPnmx3fGk8ldQwddBPrU1yNlBn57dHx6IUH/1a7SsjXgkIRMQG9nVUEcqUbWYe1a
R1B8G8IeQh5pwGHX0SrQ0eorHOrbCAgb1pgF93xDCsNoRo870gz1QfSyHlII0d4o
l0Q+8cpwYAwbhLZpWsNBvJTxlAgOebWdovXUv7iR94F8GmMWvI8VyYALdo3oSt15
Oxfeohbf+cXVmysuFHeur8qw/KfCNqEnLmcsuHDKxNKTgtgITQpq/YwlKvOpzkCK
nl6NXMQ99mNQTeadGi8tqKpKDc3GCtBPdNTV5QsdrizO45L9cmpbtrNClYwL78x2
B7P0vG2pBUHEHwKEivPyG4cCETsF89GhnO2dnBighroY9iy1pslE/Jd2IT+lOmaA
6tlj4CM5RnEsBKNEblTSaaLTpjgQnW5UcF1OYN/zCjYUm+mOncfaoz7eDmiR2a9Q
R5kLI5AES28vkXRtRtYydaG1AnCNL6wISr9oaG8bSdW/SUSzUbn4CyfJNwxrI1Au
s+vmivhs+TtHdZ3px8RLGk9obGrlG1VgJKUju7jyJ0ZCHCymPtgGytBCCz03ucTR
x82IYOfKu8pw/5y9ulk29CzTYvOKNYfvE4vAZ14wwZyuDZ70cq1W8tQsNDIihN61
lVDEDttYc9/kF2eEx42U6FKeSzYFqDqbW5saAQZM2ErHbsrucN6Gug2cI1cthlx+
1cUZEz1NExwJD86IKdiaf39d7IFTv9IJQPYDokOpHDKt1O3ZBkvN3slh9W7OHmv2
+KcGxFa1c2tO5kgRsQU2LRdDgwLbyAeAvtuH0BVgU5j1MxoabK4cB06W8xKpu+Re
b4MKL4smmSxfMULD16/5VXhEgNxYbsOgUvP525XbVPyKPYyHHYrPfqh+XyoI2gOP
sYYmncfQjpUHlcZkBbSDZWd28pALujfRssEvEZk2PoFCtwwYs6xoRLgS50nQ8Cki
LA1OIH+we61einb+qWb9Fs9rB9FfuYOPZOgQBQ0toE36IjeZ2QnHYDtXop0zs5K4
l9UaqaDVW3DiW0aaIeSPhRSjmGy/2VSitwjxMXWEs6BfbvtxI4NYWG1jZi8CyKhy
og+TNr71tewrSKY/H0T4UlFvDxNAk6ZCJzfTkhRqw+Se9+p1/EIdK22F01s2bkdb
jFqNtyTyOfUtfs2/z0lmEnRFFG6Z00LTjHnb0c1TWS3JjX5nOBtj/UC5Cgg7aO7n
6XBkTK566V628LjSKHClTtqLaZShJySiyp96Y+o2lpttJTdLuOaW7Gk+qxcOL8VN
ZaJt8KasoJmXa29+1MJICX77gcIHP3bPusVRhmfMpQtqRB0X1/PoDZYnpSfUSuyX
TRixiKaqrpNZZDatEvGvUcJ8FlSefnNBhwpaCnv3SILKZMbpMMPfKUrqgQSRRniq
RQEp+ZzGFm/JGg87PQHw8JQrdQKXhQmUOH1Nrz4Pn2Xum2LIZaZISOPXgOnPKoaD
pmqXGuDl7cJOOi3bVC5lRcsLe1/cN/1Hhzj3m+QPToFD3ZqcisPENSQxeKL4UqlA
0w9YKnXEi9KljY6XZM+IryVKwSkT+oTYAtMSdmNkLu7Q17n6EIUagF1oEUNUz5P8
T6SdpoWRK15jWAvFQVQYthsYOZz3AIu8QCAIcFh6g2LKlNudFZKNeU4QF0wURmL8
jx6mj6edSb43e0m4Y6L+yphsquB+b5ev8N75wUeVpQKYuPW6yvYaeywRuZ+7BpaH
LutZDPwe+0gI57/gSzvVYsdDDOy9xV4lkxGJf/HTqA770Lwkom3qLvChsRDbHHbi
KEZxzMPEbQ9t5Jbils8CMwF1gJkFfIRFfu5wgNm9cT08JNcj37M2hC26xU1MWXtl
vM2wL6nKnMOrKcgskEsKuFEVRf7oRCFZFRv206f95JYl6SLuwT2cgpFuI/tmDluX
BCJZsY7SpSiTEDNxuC70dLsmBbXJvLxyZ2icOoqHDC0EBj/VWZG4Zc+Og89Zno3s
eB0VE+7eQ8VH6Y7dFDA59op9e7dfo57iAvCZn/Z7p4gPZBqCTVrk5FAcdYWHB7T3
v0O3oFBoL+rAdvKbT3/66/F5jUdorJjBanrty58ORCrjn673DbiHG2unBZvENkjy
xeIYuLMY4IT4CptgNdVL9e260zeUpRqdH0wUQOlMCtIP3s+CwaYMOd6dguzSz5k2
nvtfhDwQLGvDNSTg39a2Z27SEG5l2XVxUwCmTTJIwVSLOiQmJM5hMYDcw6rZE2uv
3+OqDgBb4NcFvKOUSSlQ4jwI/fP49F9w1F/CbzEDABh+w0vARXjV5ypp7zsb7P3U
QKxYoBD1urVfAcEJLK8AEFsoYG91xTDXBY4x0xlRjtHXnXsuoN404uCl3Il27IxG
IEZZPivU5oXG+SY483d2oo6h1uOb8AVpFlWg2Gsd8O9qXoEjVe69BKHU55jtJfoH
hUOJn3NEQQoLg6inPOLRfFR+7/8aCQEspz/PDtbguB1P5W9gpryMiGYfcBro6Klm
QHnJq5Y7BMe03dxZueq0UrlIbaXZSGcTJm8A5w/1o2gscihbEdUx0Qfhb9M5F8tb
kUpf99lMJcEWU28ePQiEh5F/ZtuomNxM04TziABc0Wm4PGC9+vfGvycYi5ClPaAU
1EsFTPqVcNQt2qKu5FAWW+5KVjdEJnKBs25Hal9XRqDzFL6EHKwa1r7Uwlkv63qC
gEn9DFJvTUKDoQjKTBK9i7E6Ki4aOkNHsxFYT91P8XQ7zDcrsa/2APS9RCjeZMAQ
pWhB0IsynjQciNPWSR1xiMPkxnoa43DHVKAPDlX8katV40v8WCf4CkEmxQ/obCZ+
VhYzcB8xPIckk+3q7u9J4aiQ73gMnW4odavV6OKYvOUTw+RhnG6JtHYxLRZ3MCs3
08lhAHpKPkI3VoltFjy0MSwVh/jZ/pUNYZJFyRIh871v932rKiUbP9T3MREPSOVt
ymqiRk0i2StBvuzCTjstTne7h9ASlpR6HzOW+GjPPlU+kxlcXe06n0sqvlB3woZY
XQNQqbL9BmdG6GYa7NoMNhyZhd9GCrgR1aV7W4ASjLeaZYOO9qkEyl1HiDjHeY5M
gzZshwZnHc/rRI52WbSsX/4SOE0fCaSkxa36BbH+2A5PpL7w6m0IVoVfPE82siLe
OIQ+/IxWMx0vZGjvI++2RZIOTL0lhRs0u6lTNSqxeCubNPdTN7cAyH0csD1IAuoJ
SySoqyRMsW1X/qzwPnPLp9DLoAtuByrVZRMRaciuQYbv1LhlIm9mqGotkrlPYm51
JoHCat3ULb1JI01OGBltRE4wmXP5GJJxBMC2PYhuDH+dB3fXLEmkA5TeK7+YLoFY
87G8BddFdj9i5Qeq+JGgr59OFj+V6/8W1cBSPnn2thNgiJ2jfrq8RuGHdd5DGlAG
49t9UYkQw8o3FxPg9QUGUrSE2t93qHAr4sfXvT1l8aJQ2yFAgRlo8u+Hg2OiQX5z
baFcqdBPkwLEvtD69gGocGtgErJMNzlUC6ukTDqouoyATma1PHLTjVUmmeCxy1Ck
DG/8oYFD+ze8guIeixzedKHlj0QZM/Qz+ngz56wUmmtQsoTdYlVd0uLAp6XaJR29
22DvGclUDwhAKieogLMUaiBdeJKkTPpjo6Xf2xMlm13YKBCMo+UtPD67DfYdyDfU
B5GM9oiGaBKJXojF3ydr76j7PRfuzd82FCPDpuqSFow7xw+jKxzdtbQ90bFH09Yt
U1/Snwzi1l1yS2Owg8dVVXO+bSBkhgegTi2gZ5fGdoYNTj3BN7g7fksXTmn3VZRY
XZNXgwb07UFKM1ZJ0YfzbZGhC3AyJge5RLDGvwsa3a9oLj44wOCIFqxBb/gL79Y3
6Iv+xmXIS2FWYKBKRew7Gxt/3YRRe20hV54kEgXd3/p/sJ7au/sKaZo45mWnB+sV
LEAL4t73AGPQ8saIJbSdXsVSzEYusldI9Q1VVl4WrHe1mK5eBYBwwG/jje5KYdWv
PMUk5MbMDk29KRGYGrJE/LX4DKVMyIWIDr2b3/DJtEHjTaJpBl3XjY8XIuRfhwp2
hdngPHhkw+VLB2FDqH+ai5x/H3+9cJOirSbiCFxpVVu2wAjbl73PWmXB72hKjM1B
stsiW1Ur5NzKdveKCeEviqnJ7ITrI1gLa8jQlCISDc5yUIi3fE8NXm06nxQPQV6f
uc7do5P7wleV3xGtuMnbx/E2AFxuTKQ0r3raL0gKmRDzuLFq0aRzWA6VAOv9Q/O6
kOfV9SAXbNOQKgc+YlBWGlDazBvlDK9mH3eEvrz2FRtiPZldEcTs4MxN8Ei9zztV
13JsJ+t5kInRqL6UIfhsBw72RzQt+JehanyjXdDEoGU4AEFmchVweQ70//4d0q31
NxoJQEmY/U4+1TzT3kAtiqfvooD4WHvbJNV8PdCBsQ3vVcf7heB9mY68TpafZaEe
hN/e4Spf1Yx1hrocS+SKk4o+EI7zCA+xkjx6s9iMXdfjPyTbbAwYWJ3Z87l31Xbk
s43GT1mAYTOZgNzG8+R003g3M2ZQeI0Kq1D1jY9LQNTd9Ui8qJSU3nUnZCieOVGe
Q2kdCqwagOF1EHy+hcvK7P4ZWQpQg/q7ve119244D8bfCnWFeZ2T+SH64MJj2XmJ
SsnvYxqw/RSI9iZFp/8y+EPNqYCP3oPZfraKw6B/sav5c7B0SCghnzyTuyE8xMa7
2+sfsEauB2EqJInOvZcx8J5fgEuqUbOIKI3/b4eiPLeq1UTuo1OfD2X4X3CMAzYh
eiqFTnLJaQqOQbHfF1dxI46F03LEfrvpJpzbf/bqzmoTMuhnp1K44YwKyD/vTTyU
pg3h8+ZL3TyH/0qwX7Q1Bzi2uUxYWdiaTpk5yp9vp053FO9flhfmjY5+a9j4R1is
Kq2UjQvgT/vwjEV6aarrMLx62GcuSzMORCCAWP7fkBsBSE191vWLCJtycBzs9abv
1PZlSt0kPpZYRw7NcvYR9vWMOk5tQKsV5c49/m49c52McDs5vLTFKGvCOegigAKl
8sJcvHkGulSDtfwKNi3opzlu32/39jez5NA/9RLiZs2Rx3KyZkDZ+wL5ZTXIKHGA
8PUjWvNytoYxWpxZY4ShMnQnHLLmchqz9wycK9zmAeVWMAenGHNnKeVQ8x6gJj2/
KhvxA2PENk8LNDo8tdWuqPHAtgcujXMTx6z89HFPRetXxqjLURKVucZ+SgPSe33e
atm5x1KgfxYTd3q9lu5ijQ67wqOfHeVy+BePLutz3UqRMil84OsyS2AGj8ULdez1
mw3TuqDbWJ6lCrI75JZJOi4grHVhu/5Ioeo3DrsaNrFmmWp1wcxwkUgVmZgNsMPA
zJh0+kKeVmrSsVO6UAIKfceRbY+YrJ6jxBnD5ifUTunsZ0CagrlDiXo0egn/AKkK
JRNjV3qkWO9jwe5DW7IQegdby7Fk6Q0bs3huqhvTLtglat0rqVcAoMYDDZ7M7GRp
KHCrKKjO6x5IHSkTL5lQOcID5RLSPrqRUTIXepfezBLOtxecN983ir7E210D9Ngu
z8SzXU0SPUepjlV41CLkSdZc7P5wguL18ZnZqa9HvOP8IU5ak6IXNtDxwyqei9E2
wAef+7BanZLoihNxmWhA+4Uc5Gvh7WX+S1iKx0uOvwRaFuHzK/PMqdRr5N9FL93m
DOr7AlQoG5euLnfxgBqNN8iBIYtCGtRp3/DRjbL+17ZZnduMsIRps5t95Q1mRfZQ
3d0dPmSB/jAJB+Jttnd2jdmP0R94Dke5/v0swX9njDE2RerwuDRb58pLQtlUOMlR
GVhMIsTXvPLYbKAXHCXQ7z0ftydh1aPgZ+pp3InEGCVnjuY9DXqIaZOJjkGL3x9G
Ynng9dnf0PTS+bbgDnOMFwgJ62gAijjqmRTCGjcHnsvR8clpzTGfd0adCURFtQm4
9rQQ45Pc9rH7YTBdqGbX42DIAJ8MnnrzFP1imY/KxHgobvIne83f+xJvGbW7L9p0
o54wAsnh6MENjyMVW6jEky7x2No6E/IuyvHnmXEMCa0/4UvHPBFesjtYkLljKCMl
FNc65yckH0SvmIPrP3bxVM+35QHQQ88NV73fgHlyo41I++ek0Cx7eV4TryGEAYA+
lCOWv48VhriC/j3bpqhDud6tPUfWPXnYZGCmMl5pjpSY0b84HTgpOGUVzNL9xjIR
mL+yMLfCpKDKn6CIPkimrQ6NYSJqfuy5QWpO7p6c9I3nveVDTeNCTNXrM8NjMmOQ
e+XVVjRj+xuYgIC5OUt3vmq4sHLaNFUjC7OOUHzcaWhLz1TT5G8rAm0+0Y5vUlak
VBneA9bDWD2KEy0TUPiF92E5g2+vkRWgYB9jEYwhIc/e44dKE9yvxLAq8tWUH4lk
26eDSWU+R9zC/k0THWoPBEJXoVvuWNxqTnWeRtr4R7Ir+2AHSV34TFbwj9Lk8izy
xqt+XwhxtRO/sYispwwSn1YYfU2ccNhDp0pAeZkaakPZ47fzwXmNdyLnmHePafd/
DjE+BqEavM/YyFgGpxQ5ixCUWyh0HPDfbB6KhfiHv1myLCcBRRqBZspW01Wd9vTc
0xRbEE93OlYMsIWHjbEcVetToWuSCKvkpIJnGzgsHEf2tuLtE2l142pdqyDWPpz/
m7xdULbakshipa41GrlWtzLkcD+cNM76flyfTrP1P3LiVEKsD5NWJCw0IeO6yWRx
UUzY7b6rOmjJMHDDFFbstQ/AW7A3c1MX7luycighG7kg9CrErtPsINBHFvfAKHCu
Z0QIsDoU0qYQJ/gryNnnyWL5P8Y+iwt24Zh3LgdcuVDbtYsU1I87/RsfmUIVMaIc
iZIZR5cVbalb+Jx+v+Rbn4qocUsnFqg+TaQ0IixRKe1vopNMQlqFBzg2hWO2CA7k
5SwAYO9PqhrU1BUdVQPFYEay3Du6Ry5ybFNFSoN6APuyVMubZSk8r+6ukNyFuyA+
YY5qCJurboOe+kpyWh/6Qovw1GcwBr28GIk2ISuAaqY8ohESosKB+ptlurKCyDEa
OI0KvYulww5kZI7/02dl/cZaBLIqG75oi8qiQ27wAT4LtrndW2mO5Osgkt5gKZwM
+RX3kqX8zXABcrsYLKgHP+7J9raWzeLlGFo8CaQN1Eu/kvEJW//T+L8UW+bfjIWM
N6YZbXQYaK0f7/FJA/eqkJRSi9xrHLYU4Crf3WTcwUBJXQxRshW2oUwaLbSsuSgP
XdAC2S1+1iB6Btw52upjySTJi8HRtGX86a20yiyI/fcaJHx1blxNrGbR/10RU0LP
3YZOm5IZZ9TDRU4jPz5f6vxd1vG+kNpZbfdRuoArsEXN6YYkR/lQm2P12vkFXfPK
8HwWM1vKjgr5H89iLzC+FpknRhpGYI8vXxxm+Ef1hwVtTCg47KisO6qTI1L2cMgJ
RPa4xcPIG9LuWfpJUQiifJHkRbmyKG6EZNyuT+vy9/SzHYgTsx8tTzSba968OZAA
bVmDwPLzRGqFTf893N9AjfU73CLOOhoPLTz48iyTaN1mz6Z6S1hSXbjDlCn5z9Pg
AThEJ2sSyvDKcN6Vu95beN0A3M4b5YJdPJ+YZo2SUwf2jbIbgbYAne8F9yS2IQmt
P006MmnjEo7CPsj/vpieRNo83CvFd61Dg/zjvqblxYXcX9WFhSzUwAiMaQVH0z6p
M3mlrVy6b84PTZR/v1Tis2pY6sCyVyzQczL1kUywP/mq0uOnkC1/M7EvVDkLnEaI
v/gKffd/a6Vd3L6oUuX7Q3nd/ZGtaK3812PfZRxUbgzUjssvyVGwvvCaU9YwcTYc
FQJaWejM4FX4+Mdp7EUkbPXHD6eZWQ7DbySF30GzdBvTWT8Dk9QRGoNrHxNyx1H/
4MwKfox6aBsw/H1ff4hYkX/5tzWnbHv/mvLMDOWm+vnPenHcfui7ak1rs3oyYX2o
nO9j4bJR2FPpAwl17sdUi1cCPBeOxa+mqY6xgWO7/3buw0cYfq3lOlO/7yPMX1ea
xqrMfSTh/PJcO8uWiJ1CahLXHseJgUTzKdwnKh80i19A+iWZTaj1AmxHIP1nFQbL
jsQwH3CowkFuFSPDtom5YyXBTjWcy2CBdvUvBN3nU0RkCVQRV/CKPBUmbA0eqPpw
fxKlyDcyZw6B0GZRxPFKQSYxcjnd8W921n+Bwzq5hSaJCcXCX5YbzMiAw6lAU5e1
XPrpyx2cQluUnPICGqGGD+cR3We7KAYSHg0pKlwYM094OUT2+JgxFTNbHRCEZKWU
Y1GXhq9qVXxfrucFAkiSbKZJlDOhxjbx/sKSv/Igt+/rUMroUser/JwWXpJ+0FhN
Hs792Wg9ug20V+g/R56Rdk9KB49tZyj+lHQaaCYTX+DUu+fnx3VjsPHZtdG6cM+I
lVCN66IebLDXic5bwdhqeW2QL9J9LGYiVaLtePz01zTHMa1MWpzn0xOBJlsIZBAM
Vj6Upde5WY3scOujzXuAuAc0UmwJ7IL2tC7YFdAizaT61l1WNs5T/xn+kJC6C7rR
oE+9/0VDqEjft7geKp+3kvpUBFtsq/ACq1UrxwwapkVZMnZtjN9B3MB7f0XRkpzI
AtVeiSYryFP7QoJe9GvAIfFMWMehLXFJdqN77TmYQUFuC/kPWV7+Xguw5F8pe/+C
NrmPzX5G1x5dZRuiQ09DN5TL4/2yIyaFvyYoZq/ZzG+oy93IH/gpyG/V38g3RQIu
Jt77SLYNLiSqMoWbxYxFp99Z+fN1Itw9w+RM/y0XzEqQDTHa4kDnwjrCw5D0y3qD
bnZj4F6aFffCKB3X+rHmunK3hWqGSIwnPuH8ANCtrVrr/rQviC7dCih4Dlu3LnHs
NSmKr/DAsaGeT4P33PXqqOjhbFZxNe0J6sAXFi5yg8jMgFF+BiEdkarPb3AAj9Nl
KcvHyTXtmOi2VGvNsQ/GkzY4kk48AL7ZtiJgnbZCIxxosaYcc3ZQbGPHG4EO+Stp
xtwrtg0Kk2UzHATluEOaTj73az+j2YBeqprRYG9wk5faroGqyi4ruLC9oyupRMqV
8lnxArVWAJrDjaxNvZdJbVKS6OHPmSWbUqrlRO46cWC1PPvVnS+6gv1Nk93jhx7R
EbEA73Nq1JLSa0Cl8j9p6PtjxVoo/sUwPgIPkBVbqgYGqdcXbABQRYArMuLrGDjv
PXHlfmpLqvey/xmduYkI5s1TAQMyLoF52yN5liqRAlXQdcrfw0/39JVbAlP15Fjh
3JwFAHeIKtYKs1bZCJPlIGDrH2vo0OuO92JLY+3uP3zVNhHsAkzBr3yufb5jsKus
0fhmj1K51EAyHCnMquDdMUwCKirxYULDC5+/XKwV8qTnkHyXhW4GustNFjoe9yx8
zDA9U2uejE3I8poLajAgPOUonPfTxMu/Xz01HW6Yj9A8wFAb37ydz/j1mOSuVenr
nTe2PbZQHcMaxQ9ZWKc1YJ8T8Z6QoCoMfqq40zXocnxmQrfoHEu/B4Y8YEaSTV//
TtVL6aEIEY+72c5diJ6IEzw5PkoLXtnjVGSx864mnn6YrSeeANPz48IV6qSb/hNk
9MrFKLko4FFqxpDD3beFeMM9UPXwTQK5W1D89eqUteO8LhAYwbLM7WAURcuSI4mj
ZwqRObDVedKTWnjo7zxAUR8IEPHvyXIWtGu0Q+04FZziYGqxetu6lnNih/6XVYf5
nnYYFE1k23QCd0qp1Gx/ymDotSIkRTMOGBRnvuRbFxfJ4Tn/xnnMKx+F+diSnwJs
JR3l8ADBVk6+XQ3DAGCxVA2bYXcfGVc/FlxplY1eLPAlk0L/T4NOcjQAx8ZinNo3
Qo1c09CurG3dymet3XYOU/i/n341lgURtdNOKuhHgJV37fwUrfYZR1FG7XbIkwja
okizU7Rs5ydmPMk1NNp/5K0kWP+tB5brd3FoemNPlozmH1wpAX2TBiJVK5GXt+XB
JZhrpkqT8zF4st4l7yrl05dPce3lrAcBdQ6+4emQAe38v0WfxPnQcqkz7BcgEbdr
SRkcgZg8lLqLf1Q8joOEXmYcWHtqw+aMQfmWd7Qt4cQsw1QNtiy2vo2H8KhYXkKn
Qg5Jx6N/dEDtc2g1qyTIFukGITPY33cFFdlMfILKiMzjrMVccnBl+4I5N8rC6Z+Q
6UX3qQXBuUZ+EzLSTnKzdjxkojgFrxrYL+YU6hWqIwb8qZSyUdJKl/Hes4ppTA5Y
hCNe5mGdGDdYrG9xSQGmnW+kXw0Fvmz6cAQOcOl92132GaVlFTdYDkasL11B17Qt
SbJCbz9AcW7GuzJkLTv4L6m4HRHaU8iMZp1BzbAL2dgVtsgqnQt2hhOuFNHKYkwZ
9H2c/EftJAAUja3E9BO7ph0+XtfxLkOIzk3XKsHqrL0u4rz3Hrb+itN2LBHtzCqH
FGpx+db3A9lEWWAMatzaWwrwNehzd0AAeNu5ZLLUmyW27Q6DT+kd4KMbr1WUAwYv
qJ225RHkw9W+1Zc5lrUAYsQHIjoQTy11CxwSm66bJKROfFJy16+hL15YQAj9o3Xh
CHl+ljtVEpq9uRG8+GSShRM3TMEC9JxVZ9TirPaN80KOyjtc5SnUevQXvigqdK1v
viuG6GKZ5VJw+nzn845m48xyZnJAr6UEnabfegO3SiOwA+KCH8YcHxoPYiYvc5bk
YJM+IUiBkMLVIriB4kkke4VszsOtwUrX4ZRTeGkdDKr+xPjBpPWoxmLDBx/vlF6k
EQpGJie+cyidK8tA/g2NXvbTNw3IvdegAFBtUBlBS+YwTO3VpgdBtjZ68Ekd7vtR
2BMAd6NTJx3BnI8oD+A4OSZuIna4/oZe1ZIGz5gat5+zWwBLhszInddfvBNCgxAR
b0dWY7yqzSOoSvQ4ThNhGoVF4jEo73dpTAb+f0vIUrjpDd1Hk8kVR2o/8b8wecjS
IRJ6+TC5sHTyDRPl/sud9cn3t35qSv60jASUW6nL/6tCw4U7bMXHMzFVXWc0gDcg
rvYn3j7LAjMgTAqYfqw1ZVKIXFNIDst4q/Ve9aUokJ2FApoZmOO5Y4RU1P8sEmWV
wp73yBIlUuRxRAITwR0GDJ3HyvgLEWxJdnft6lR2kFUtoIHbBMBbaB0R5ihz1PnS
xMTKwcn08P8XQsbh55Ue9wOMT9YNewa7VAchdU2kPsoRO47HF9BGRk3WJhYKbGl8
5nCXaXeym1MB2UKF0PUR6rLqpAyDBoHRpSK0on9J2YfqPAcHIDzKLrOhkGd/ccE7
3KwliaoPnJ9cmACcPS0iYI1MaVcMN84aJM4iCtkkfmbJl9OfiNdNUmopbPOnZSKc
ICx57EQJJfkbtF5IBXLf+eDYMiU1ZvM3b7hv6Ody6M0CkY4nBxh5/UEUjAFPfK9D
N+HHvoNliJYuLVb+vPFukiRasYhelrpRTxGoH7HBJviLdjsImWgtF5mDwqoroBTP
74Qaec42ZSdNBxp3mhQRob/b/n8bcP008YY1UankRnZUaLG8fKt/TwKhnwvgcU8P
+dlrMJirL424ApvS5rTEry0VyKNp5afc9yCq86C4wMl/T4Nm6SfHY2TiHAYUak+m
RgPIJra0r+r4rReocLu9x+GvgSMs1aKHiQ73v84/4rXukX+OfcAvNr3mp+7pfPvl
b1uIuNsfcuiFvT0CKrngwWVlNRk34wva6IYg9fV/KpylP+KslJKoTheBabK90pnU
6CRCLWWsAg3aHBF1052jCf45w4APnPzVSOeGy3NuRH29pQvzV9KveRakvynbs6pI
c3cclZYo8cxDvg4UKYjXi5RDtmcuc6QOlj8xmJ5ZOKJlRgjMDsMBJTaO72BeaXzW
v2FKPnjWLFrZJxQBIN2Kr5r/Wgun5hMXvF+iofz+t2WS/9A5JzlaYTY9bDIav8qZ
flF13iztJHBoRa9ntAMdWTVmrpxFPSWFXSPgO39wo9gZ1iJo+wqIWIAmDspD8HC5
Y2NIXSHMIkuK3Tyo6Z3GZtb0d0RlsuRqHQgOopIYHdYMtjZPxK8kSiPtPs+F+gNM
9lHCN6ouoUJBAX9SGwyJUDjOo+BMX1K2VSXTBxDoSQraoCuPNvTDhPOglQaQKlqF
4ajJUkCkhaj7M9yhF7C3Tt2nvaOYFCOBRSIbjoT98K1KBDy8+YSjfsCAbj7tOCFg
qxbRTmY6+ZOYfPHaNeLkK1EoRrP+rQaWf7hH1XbmSpXCAHUiYfVS047aAx4DRtY2
sWThdC4AZECrPX+qqkvaQgNzu4bGb9CWMmEjw4GxQRZ3TmYFslQKwwYUk2QJgA0J
A4EbZ0wxKqRTfE36LvwknriVYGyTW07BhzSCkZ/v6u794Aoo9A3AqB/g+oLeSUxa
EYRKi6NUczYnKIsf7DRk9z/juxRCdDZ9HFOozv6xEC5KY2LLAROZbut4UKDK8UHE
6dpmwu6pxDTSu93dPzNTMD0wDovaZpSABomW0HXR8fy2U4KCf8ZvCkHU42swX9B9
GfUZpWmRzUuVeT3G1FUrQcO4HuImaErPdObfUuL9sRsHlpHp8pfLCMnS/BXanpKl
RYzIlit6DLZc4QgdZQxen2+uczwXevJ/aeIvnjYhU5zrS/o7Gkataq3sy3IgO/kd
xIcPaJNoO2jkcdywQ2WFFKZDyBziLR72FUznHw4b02tmzK7lHr25en6hAoXyC2zW
4pYdP+otA57UHYi5qxm8cxfpE8uNb9G4VVnhtEiqp0Ga49cCcUISe6ZWH7s/vWRK
jRKaWD2hgcf3M23bXDC1FnmUvRLPIkI9M+2/X+KvM2dR4G0Ydm5MxFe5oO+LTqIj
484yug6e1C4PybqFU2iNgM+eEG5j6svivdQXYyFeWbByCowmC1NukS2F9WCcn3z/
cUoE7pOClb/jZUbM3cNoeHcNnbSl5+QVtbwLp5doBR2MY3byMUpovrw+P3hMOms1
2FPp8XZY0ZDrgD0+hO7aq3+tJFloGFs32U6Mvy3zPaP7edQwAUeHCSDJCjuwLzGr
Kmx9CSrySuNH0wxpIWxffksCWlFjgSbS2j2qlKfWukl/5Z3RnvrfRrjR6w+PF0cO
s0vB3gP8z4+YxU0BgSBnUngiTA5yeFaClVF+85qBJZx9ICDRl6x1aNC+OXYVSqjC
n3feuknP7WNof5SvrZaK9kJLqU8vaK8R6nfbsg7ixqWoOwrtEuUcHZYe/+2YmDyA
URSL2hE4t87V9kcBpIigZoOmD+1WAkCnshc2eCxxF/2ZwKlVuaMvvJ41eeNGQ7Ut
oVn9DINcbZbYeteQcqnIUcEHRg9lgu1KBXLnRt9nOozkXD7kmL94lLXooKtiicIs
kwnH0c8gAWttrhL7PvySz44ITNAeP+xfH1Vgv+SwMyKQIgmUt2zYoMbJMevTj6n5
lpB+GgWNAqdI5HoggCpqWw9yfCj8nrZlrODQY1Nktx5mJDPRec5TqFyaYmDI5k1G
FyyZ99jEKiAzOmVYfsXK2A1y3mVBQmv9VMIEXLx+pNflax972ElA//lv7s2JC559
3RS7pSNIMAZpYBNaCxVSAE5GOtDsjD2H1PW2uUuQECs6sEF83x78hKw2vyeRPNOZ
p4OsoQEsVSk5qvDVHiTFcyTzBDb1WMmRzSw28QFpT8ZLUziOp0ruLYoKgfB4Qh5q
XafoM3aiVI80gS/vVWqSI0jsFRQBS8YY+Gi7Fq5r6LqyMAqzs6Giagrr3p2Nm7ys
VtwBGAFQfUdwPoxxcTiO0ivrGul0pyoZbn7AguUDw6RGHNyfkiyt/99/ugfT9Mli
19wQNETKPAMwYTohoe7DKRwlOVRsdh/6MLPnYGq5eTQIIFhFlNNkzcYNuZJPxVIZ
cSP/caBm0SwN3jLxdRt5GEEr3WVBttDh99mS+XE1jtfk511OAHQTfRUkeLrMJfK7
4LV2MOg9yhDZEHN7s3zdZmCmxMzAgbUxUmICDz6IBm/IFLMvZZV3wSsADCwxAxHL
PwxPC/gPIGJFhgWHO598pHNcIP5CmkWTV2t+himhWDUs9cwy0jExPnD7+wxNKdF+
NwKy25FGl9faTI4NOIwFvl03fJEOg/gTXXtSVuI/1YeLYErjocNDhAfk6KkWU1NT
VALWUEp4kUldNgvHU3AycQLACkreJwHaFvukarFy0YADz59RVUrS7NEu4VMfbp4T
BjVgEzovbpXpCp3YdCISVJT7iT8IZVhzYO/i/4ZfaJFjT9cyfZdyyGhVOrCCHsFc
3xf8daaqQU1Z33IeecMk+xEf9Q6iC55PsjSw8LsINC3FS1P3MyXizsB6ybI/omH/
RG/tf6Pyon5YyKGJineHvQAzz8u3Tc/xk5nXCronZFjqToK23CNne3eG9gOERAN4
fkp/d6RrLBx3DlgruSsmqKUpulSS3lKMbozVKlonyVTHm4sUpDeBsAs6zOXVKSDW
r0lXGFeABySbEWEE1SDIrCaobqG8ZoXkMs4u3u7ZzKJYduhBpcVreuLZYI0Qk/+r
uDJj6+BnmWMC+s3vfGs04GcMFOj1F5wk39/SoQn82qECTrxrGkx3Q5O/ldiq4acL
7qLNyEXXxMgVo3IoSmITJCveyUXhOD7eR31K571J6zCZe4WaErQNosMVJtkQBjMJ
8HV+89SFmJTWPWzQRpLeqvUP7McFBMf3qPelpUhhLPACWi2VJuxDCcOi3wm/f10J
A2foJICr7lAFGtzkvy7+ktZ7D1q/d02JDRIlD3oyqmyMr/+xyf0bQk+tEe4ZWWrS
nWxqnwQ+S9yp9of1bVdwjqG1qqqJAghLvuprmApdCLmO2MPBpQIRIzpCHLhH43t6
UlorCvHb4Hx6V62H8Kytc9e1CwRGXtSeuOfGYA9sEJ0oyluhM7ZgojhRauIMiAeG
SMAMcuDnmpmBq5bcQD3ppUhR9eP9eFXt9p/iMUzbj7FN5N3+ikm+siQF9JQxt8QQ
v2McH4yb7ubXGDrI1yXpPiyYe3XuGhcZn0/ICSDYG+loLqDnIXdMsVtliT66f9He
Y3fwpqGbbyO+Ls91ZzMaGlTKErSE0MsXcq8G12JZW+RSTCJ3aUHqubq8M5gRgUAv
aGjIQjuNZlb6rEYY/hERUvb6TP5zjxXtyeDIKTDsghKJKULdamZlffS3eGPq7FVI
stUvJkDj2mSDLMCLg/idxYdYPwQzuWpZ3Cnm82dCPt7ZZYyoe3Tt9kTPZUrOeq0s
d/ONKlA7pZNKlWoHWbsGwV2ECLOgE3osG6NpoVuA8PszZJDY+DrHkbOTvU6VFM5w
RTFs+zzSdYh/IC5ANWG9VwlJKT+BeG+T3bUjNgqLXu4PEYTPeBYZEMnWHrRS+GCb
MQpvMIu83fpvujUtjaXygvZ7Wvj5NB8AQmcvpCRe8cyDapQi2VOb6th7RKnuO2Py
zgdCaMM0F+CACx6eHLYdafaA45QL76qlzeUzkMZkoMjNsXmTe99GuluZK00Xt7uA
+nn0IKDxJ2eatAXa51uFeIDKbz5SBBvyDpMLZvl9A4I6TuUVUhIQXDSsEEikWmBs
9nc+E78qETPImc2sAMC/3z2MFUmOw5w2RJ14drbRz7inqp1Q0eba+dx+lY1dUN+Q
8O96tWoPE/oIMFH5gDbB8T/qAL4Mut2TPAMyJHFKTe3XzxYS649RSkXBeRFddj0j
IE3MD6MW5fEVJQAdWc4fVDnDIHTKP7uN+n2a4d18JYAkocw+A+cndWm+hUGeoBmO
5yr+RkDQInJrg4tsfSABcQtq8HzeUdvItTr1vLXNKjUYdbHyYgYSOuheSpPHlZl2
BsTIMoyFxaJL+U0CxgvQ1+vJEF9qtN6io44XIuqCNfnguy0wfNcb3D0pJRKHIExz
WVqfr0qny3CHyxpIbdKoLVgsvxR3E3L4yXKvgjv2gwNVx+v8jwpS39OKkgZ/dqMa
nLeEkXJs1C+1by+IWzD0izIViAirgvz0fO7l1Z2S0Mmfs5L+6Ijbr7oOq4U61uUR
11MCW2yeEtpBiR3HM6ypHbvYl3w2PvpvSpdIsYCPkGic4CP4ebeIqsO53fgClNou
gqKRJ08kVEE6Naurn8IxNAwc0VRowhQspubo4+qC46k+vRO9n5dtT7J7u7StZGI5
lPEu0bId72Jps/3z9Wx0WiDGW+DqZqBRZ6sunHjyTzPPi0NyGsqL1OpS+LzbIloT
jHN9HYNjAysA2EHelil6LOWzNN6bt0g7rMcARPBHNZssYsnpkIcjn0E6cOaeb1lU
cOnWMXz5Oc0v+UGr8lisUOK4b/Pqbucv3yMmjBZyL5OEsDmMO7Nt1Qkt8KsE+v+P
n/oAZZLe6AZju7W1qAorLG5BzixNNJ7AQ29wEIi0cfui8sOrETigX/qiZw/BZMIA
UHsBgKgFURaz35xFMeyvTdPj1Tzr+a6X7liZXGQNY/zES3q6XIfXHDFqLZa3EnVo
u5HzWfdw4vQq1M/9/HNzmRxMur703HmyZNxmQ3/+2vaVo64eun17hXxrioij+O9I
sYbExJwZgXvtjujs34i3qyIwfUyKTCFuK2tS3t3SzYvzHX2iTir+HDl8meMVuCwy
WWbvcpzTHjkwyNE7SIFcdu9xZt7io0mlKv3mpbVux6s6XmSxHH4fX6YW6RRsyRIh
3ZUtdXTPFyt2iizZaqrteYmnZCmZDZAbfkqaKabzmeFY6YBWYVp4VRKSTwEf/qwd
eyN5HUvPiIVFGrWco9jbd6n0Lv7h1gHS9x37ZyzFnNZYb0a+jZhNFMNRym9tQojn
gWHEN5jMZ7gKXNzTbO3GF1FzaXMT9iJsOuvLuAPaaL62R/39qZyeXxvGN5O6HgW0
1Ah10+N4Si7oSW5TLKMPkWehOUvbF7+VSdUuxgOlIkBUcDVwkpD8d01dNw4wi8k+
R2uTmKgly8yFmZbParkNOjz+FT61orqnj/BZNvnxgJhS57MJ1WkIDsZbFSfwBLfj
WXYtvyanP/L2BUSej60VFhkq70pHq+YTEPMeeO/3rMh5HytBZUtyimbmFHp+QC0y
+7tz9eqzmTn8ghwF6uiGFxkHBujHKzNG52IwkdvuLTrKIW6NpGsKqr8KVHH+mCyJ
6S8fp48vl+JObscFyAT0G79HkOLPtiORXjnULz2tG4584j3HVaFOTijg0TQ80aVV
7gVd8frDmM8yJxf28CefI+jcoE/cfCn5ZM3CN3+UD2wirrUBgsAAJ0wiqEhytHQO
6f1T5cnD3V6etPK9619A0TWJxyt4mWrTA0jSaI8hjwzfiSmJ8R4XDuzQvdUhGRY6
KB/Wb89xGNG4E2LatwPzPFpYVjbwfLDhVglIAHFDwbh2cYIl2j0NPCq3snDnWgM4
SLHSekFCvoMM0OS2mtVJPCfIxG/AfSHuMpTFg+hiPtTz+y93PVWfxmx0P3FUC26Q
Cp5y2FbMLlig5XQuRkH/XMHtez3ujkPGpYzMLPMydSGi6FjWcFFNgdB6TZcokCqB
/68dkE2SAuAaTPp+ZnxIoSiaar8pHOpTRO4mXqrlWuR4RGsuf0u2zL5y/FkmwQS5
+6b7d8C4MhZVr1/3wp6A34UWyk3TOlk8HbRrBibeFy+uUKynlsJ3/WidjmI3Vk2Z
GJET87bpk95DrVW80O+E/tvc5p6Kkgd4iSUGMtdmHu6ORH7IITe3tDQIjSobG5bA
HURfUTzSmY02B4sF7t4/YkV7gaxmH6RbeNmAyxQ+RqbbCm+TMicUJ4MW4BU3gNRP
yBCEaHyZ/jLnBmHSzR1FSlpDtLQWodbYd6CF6DYtbN/SVLvzzSYpRGuveQR/3Xvg
0iZrZ60+r+iTwPmo5ggJZ8G2LJ/M8SMcAAPYS+iEWqfzhFZnin0zU4MyGT6X0cJ6
PBnQE64nL2/mfGfn3H9jRUObH15PCut2vldcSVhOtuVPRqan1fPTHK49/4qo7BUK
eMp8cZuMW2LP/+2llWUnNp3Kbrp8xpfvUDWg5amxdZKMH/YFNPsueeJm1fBfD2uE
OM3flOqmf6KRarolWSP0vAKkEQac6U8mzELmX0WEbj+jM8xfS1s/2UCD4GE0NNh2
vSL6cOcXJLJ6tjcVOVeOSnkMTRO6iav+innwMzScqiPvb/RoOGic0/4xlFtz+o5K
8Iwua4CazezAd/Sa/eJRAdURwH+wcBWpmMk1bioh/caWco7zVn6iRdPHZmomaPlf
lT+wm/fWo3J+CcMTIvXniCBuqeBMsiBfxEUxf/RxgiFU4iwlSgr3Dj4gU3Ar93Yy
r7tfsCj7Mt32Hnnp+yPnFT8rs4y+3/B2GXNQWlfiN7ebdozRBRmuO4llIG+ck5sT
1d/guU5KlzTzGyJOjCnBKCq/Xv5IUaWtwyJND0P5d8ZJxvSczMxtl9oZ6y1Z2t3e
Gcug9YgrtJHiY9Uo8Umlqr5y0yCK4mdjLTXea+whledQcnOYBl237JheL8w1TbyV
Vl6Ao7S8eM9LGGoJ3G9S4l1mSy+OmfkgvOGgbIsnlaDyTOT92JQdAoNWFtJzFmTH
en8QB/VIZ65krAhvYBQqRDMPhDuVKT5+R6SrDGQ9lWucVI4bArEQwOpPFPfr6E9g
CbsLr1FmXhEzDqZ7Tnpl3EBiysKuVlxMzYb19YKm9bXVPQjYkRGzoVQs8xZIiHV8
UdyIQRJE1lC85TD/b7BOl03ct4cR/PRA8TwFjcIPmdOZNP1hnLuy9LW6i8C2Qm0f
boQrHtIseymp+2JhiOtqPX1ir2dUJxJjrHkYqUfAlUAtHXix89gGdiSr2upkiZBc
zjcf6nE9Sfz6fMg1fbUR7RLGyN8JwJjARNuX4z72v64QNjPTQfUXvUeyqpGlsGtG
w9jEita5hax8P2I/ec/WxdbOZhnL08qZ6aUparTuGQom4uOKcS7K9cdg00GOVAd4
Km/ayG5eE8j2nkCBmbRUsTNSbY2nLVYyUfKlIvlDMkryMkXQVDU4b+CnSeI6IxBu
pm9Owz1eVLxEHWd7WyVvH1DV9m3fh4xY5TGOtSgIAwpoItPE9mG2VRBu66821r7P
PWYwk9b2EdMeE9zPqpkPjk+Xl3bEy+15hJV3oXJoYrGo8NnCrZBuhgZq51BseMrp
MLiBGjBmqIqMEmE2wrNg+2/LF9gkirVKjzre4KACFXWHOy9LqeTpet73KArrnWvO
uyRAJENshdnhCVZjMU6DwpdxLRYaKUqNcOZbxhPx63FQ1bFGaU/H5rckI12/OIN7
/P0POx68CU/yFN79nC9FZvSmTz7oukF1nfSYDft2Rr+ggntyYBs75Zw11kem00ln
yh8rc3C1LyMDAL8QEb9yT6xprbfjyCfLFJ2EalzMTwqo/KXwB/IbtrovxIrLYNgp
E9oSs2Gv9RgN35WSr1EWI5eWYfuiuxEhmrLJHVeiHJMzGWgVcQt8Yt9HiLYJ/ZIc
Kodpivau14VBvHzRByO6Qj0Tf1DTfm3kKiSg4Q2iPrJ+cVNwbApWRtvezlF7gxoR
jt6syzzgcuswotmh3obEzCyFhihgdMM+XV+XzF3saHcUs5UcGKtRGt66AGKZ2Z32
H9NMf7HlG8qCyHoGuW4V2jB4Y9oNdDPRqS5yHt4nDmJPZmQxv6ebf5oRHpiSkPna
wR/zGNbzgvSSEVrsFWWJHK/F0eznpzSi0LxBQU0C09sJWS50rk4Gpia9UYQnq35Y
2hsbxbACFIEd8G0DAPdMszBmbxB3A19ONQwt0+S63ad9lgnK5kKMc68Kj6a0aujL
smwK3xHGclhsV1yGYH8mvd+wQci1lXXo7av1y65w26mzK7Dt0pD7tfK1//tomlha
PYQEwz0NOObjB9BEbYFZTHkRagcm0TY3xoj4eHDDDoUdMEIUbzt/6att5YdFoX19
9+Q2YKriJP/ZCnt5kTMU/fmy82iOIwRS1hMLEjPblYZYXoprnFehRklApie7TFgm
y22E0zPWh15f4/ncxU2DoVDGA8ZJGn97NHw8w5zoFaaI7GsB0tOE66wyi7/Tsbb7
h3H+P9LirvwDxy/W0aQ+Tm+ddku8x7sCDCh0Jo57jdx2GPoS51cnHh8r1mjWZRJg
ItWWY944Nv7QrwHgwWHOHA7dKkebMtwwLZs9rmYArHlc9EziriAaBBsoUNl2a9lv
ukgLT66ZgqWgNrvdA4Mnz17BOZpcIO5SjETeIJkRzeI3SYgFSK9X3blplSLs2nzW
6BKaGnd4plUdSwFD+QkbYVX1E4DScbNdj/n8xfnErmmF2Kc/W3R0iVqkyyOmtLqq
2bfOKvOcUCR1zsQlKe1Xshtsp93Ooz5MnZ89IJSurRNysFX3ocjWaavJPJt1019s
M9QtyhFcgiCB9nuBSQxUOuExrDj/hYvMlO7qxcvMFOJDFyfAckOzbDSSMVmbVXq/
kn4lMHBDHU7K/OPkttjFgVI2Jy2ksvwJsmY1wQ8ILd8vm2hqYfyITxGzUvUagpFk
el6SvbXPma+GfVFCKjTZog6cgXHM/GUVQ00zUmKeUGNFq/BRJautzJ8dWRvmbK0N
hUalGn0XqctGuojkWX+sO6ohPc2LOdVenxXNzMcqSwGhzIaGtQV0436w1h3Dlq1H
Aa+OSRiFssRovW59MO229JlSZb9KyoFRtBlIeE25fxApWolIlvdI/nNJtHWj9npK
0DhkaapE7lKM8ycxPN42uO1NCScB+mrtap1ZhKOrOBKb6KKXBjvWZ4T3sE6NJjya
2llLSTjHEnswM1a5/GAIxeIsvJ/LA9C35xkDzWqb7dwhbTueuyMdYk3chmbaw40o
Lb64Damyb2TwkdDB5boQjjNWQdTtql0JN3E+Lz/WjirWYcR7Q5wuAj0wzH5hbbu+
fv6bC42fcKH/yVSk1x1tOx74dAaXSDebjfA0N/4vWJShR5a1N/+/3c8Let87pjCJ
o0gsCEOVbdl0kQ3O/uKFfQqlaTbaAKQ2xxgywVfQ3BLix1OBpcr144vLrPGuAK5F
0ZTAbjy0c1xchg8gBkIvT9gmRWJnj/NHR9JfmldNOPya8dTRL0LyUPD5/BSW0xpc
3ieRnIt0MzPrg+u+ppDDyfsBOB6+YbZdItMgezRYhnUzTwWPcxRXcOtHGpqS2m+t
KoY5Co+uKCtDrRGZfTpuMG5UsWOL9SggOrsSNJU/i7c9+ol7c9R3syJcsqQDiiZK
HDRSYBEhx8cjz9mkT1vXgXIlty1bUTlClHAc160FtOgRf6lP77L13qcWnOwkAai1
fN6VnLhj73T1Um4qYxluEBxOeicp02SDKE+Nb8T5w5GJTKKp/SbiyFxVN1wrQchS
lQ5fTU8RLMNZzWarvdfp2zFVk5MwYAd2z2zxeEmCLSkPQrewqcLdR5WYycubMbUs
5fQej5vOPWj1yA5bx0HpDkhKc12s/aLtkjCAZfF7o/Pi88Xl2V2k8rMRYOyRXokE
7JEGthv7oyxFJhEJwDgHmY1PaMNx3evS8abDY2qd++JA0dsVVMSXi/eUGBqrcGMM
0zCf4WHq85luq84iI/5RtY1tKRX7XsLZ4zobdBzPn0k+0HvoI+ja7lxokxLj909J
gE0lQ3ZGJcOx6hv9Am3AhkRxRuraifqS5kO3letu6j9mbrjZnX3s05kywuC2cg0T
oOtWN6RZvRb1J0hhdhdJJ+FqSw/QxE6klVRfhw9LR1tkUc3IGN9TpRsVPNguaHZ8
ZdC4k/1BIc4kCyTBEYbsPBTP/A7YABartme5e3udup6PeOpqS7s1Q0Sjh5V+/zNz
JhS5A/UEf5RddncRVHTRsPVZdAxRG+ftvKMGrN2tAwN5uxtQ9UTZns0U6fM6p7Nd
jw9fsTdkGFsZ6STw2HvazNrZU5Q+b87OTcYodxZkpOUEMpRHvYSyTchddJ65a2QG
jdlf/JuZ4j8pb8zB1BmRbyUreP2rE2gn5TsIpNopUsw9otoxljKtLePCPrWF2pfw
0CyvnRvtMP2LiPwnmuBcGMNbzTNH2ENm2GX8v3VVpuJ4MKV9RBeTb7pACDZ48dGb
datqIL/0B/U8V/emsQwQ9q4b9bJkoP8W4DkrO1jfa9F4s8bldc5eGRcSRRi/eNyN
/GmO8ijM/yPNxcYYmtBAcdvpI9rRk/gUxq+xuDVEXis4Q+SZ9XK1HSeThUuTLFWM
uNVBtIyaoqI6FkpJHE5UnNiwFmrHSKDnFh8Fdz4e9jxmDVfzjDo30mkH64b2LuDe
X0PDVS8ftYHuI/YvORV8G4SHW0ZfSN2gk+3weCvdrv0DL94fg8VbXDHLXH6Ba6RC
sjLiUTya+ve2sw+fI+oGLSofhnK9K8FUq1uoWP9ugM3INPQKxFBxnBnYR3PcmFsT
gs9JX4SIl+qDjjTs08lh7XIhRRDsxcMUcpveqGvCqmgkKZKfNeFGexRdQZGTxNTN
JyYldnnSYN6fUz8xEeP6/k437R5rztsohjBfkYNjIEe9PKswT4bgQfvv59FhvdSs
vhpol5b1diwOTLonpPXznlkDpfmlb8o21Z6uML+7LgWDKSYpYolCIiqU8RK6MDNS
eepyaO3l/L1akfCzY12r4SatANOSz5ufPlayY3YZD5gv+1ZM/oKLjqj+P3VHY9SI
ZMRsWd63fHRM91MGCRG83PPFKXy77OqsLoBsJtvzuxND1z7mJSQxrMVk6mW1Acrl
V4YmOnPhQcKYqyYVbVZpAY/NxtngE+A/LlOvcoBgAFVKXRxe4rxZJazvLcGxHf9n
DbXkGhtPGvPxHvlXiIK7nS8Abe5tv1LVt11tSt+LEtID7Q2Yt1CxIfCbHanqWoHO
g4BKv4EGYt/KEVc1fif+vyyv+HMHoiE5fD0qoW2YaQ+JYnTPmzzSK0Zkdg9B68+A
gZaxi0Z2qYcxmfFHDBhVhOpauiYTjsxFmHFEGF10D/X9uFTipHCE3Fi6l6U/oLZ6
zZb+Yv7fJQK+KqoDTqk7VjP7rpavAatmx4uNjtjFGCYwGvMH989Pls125zLIBBKO
2Yf9zEQTER+xn6x0UBU8zp1vIgtGMIHQ8fpft+oAsNJzYRNUHXwCQk0vTEAy28dC
NHCIQPQxlQEColCaC/iC8k4I73LWKMNxPsFjmDxGW5gDuVxAChRAc9yo9e5LuXbF
AESofRkBAqwwOtiSyIWjIfBsHqpH1o9uG9EO0GnSlehjGA59iy/UgHEVqX+YQrBW
k5QxG5sjhFlEycm0MmACrDe/3rnpg97T0m38OFRRGd2dznpkb+wDYIETzuvZIhre
TpBQtNxtRn3QmXFGpK9fB1nmDRap1ZS9W2laHPSlU0SZNVcderXr6xlCz8OWKzjl
vQaX8TpMWA3+Zj247GlYca2Y29QsX8MekjLfvBV0KH7kCTFKGBsiVND5CcBgVfKa
2LbDaHzLbNzJjHQqf+BNObKCqje9reWtkDm37++3rLjzJ1yvBE3iMrxAmwXMFM84
zpz+06oZDVMVM+O+7NfxfWLZmO3fE5OfJe0UHA+qkSTy1JChRe9HasXLJ4axmMXC
7xMfgB12OGGybmuoRsWekOfhy1Xd5H3HT5z0J8X8DXhlJqkyl1Au587gprfXD+f3
PWRR+KMPHmyDaAdsJx4LvOWH1dWrZrNInVNZm+VgiB37UzKdjUYXcNF+cLtecdyg
Cgg2UWACky5YyNx9dSr9HxFAyUu6xIj+C/0x/VY+JXRlfo4JA0O9P7mcKWXgS8sZ
/RtW3YVD+kmuuZd1j6DSFcL5oRg8ULVkhcTuLs9rc2vg7bm/0a7kQblcJ8VXsT0Z
4BrqIlePQaAL1mQsKlSI3Z3ehRnmrK9sCISSJEusza0ocCVG7gHJBZF/T1DztFJo
cs2M1pd7jYW9IAU5fBWmcO6Ww3QF310bHLtMUXgNichL1sMzAbe+GiQtkzwTRxAG
8QrjCkpxqQBG5XsZylgcFMZg9PQ15TZmJzzsTiyzG0wLSPbi15IbrQyz0fV2HQyl
xT9JqqhsiRnAR0Q0n6tr1FqdMRIsRvxuE2r2XmFo3/nDRTucQ2z61B7ROeceOTEo
lwdELFSFO2vTveBxkouraBUYDkfgKNwbzXVyrI/qch7CfEON6XoZvdEuC0kedhMF
5uDKWLD3Stv+9ndgK+fg+LLwCk68qV0fSmzWr/r0cNZIgs0fgKYQnyEyB6r4Oatf
KD9O77q0dEQZEnffb+INiJt8znv/qhtAm1vMaor1v+hbKdzS1vtea+cYMthigjX6
YzxKj/P9KlaGamKrMw+w71Jg6BmWS/AAw35jPfHVdIGWNWiVYGTZGqd5uKVoMs5U
t4GSURxU3DKtAznTgCcOapBLVmMkTsiqNt94C2AA/PDlOmfcd7QBFG1lh/04KXx5
14W4t2L93o+JLZzpRSXaxamlhEpz3NkcAOxXtEmciNfr6+f4fDQJOlRurTRHbc5k
i6GglvcjXp2pW18A4VfPguDquL88xIh4nikMdVO42ssNO5/kgzP7lHF3ilSo64ak
bEadAKq7QhunZ6ZoV0P2ap/Pyi48idBLmcBkj9PMsFRH4BSDGTkSew9/FIdQblUv
vdSYfiirKTDOqXiX64I/5DkBYWJNcJmIMTT2nVgYVPacWamRgk+MsmuVzHtlU5Dz
HL6KhwZXBXvBhfrviYkEFeuNgXZ3seyvvJ21h6g+g04SF+VdDqJ0UEYrgIDHJbYV
e8MfqORBk5NqIXo9On7IM75iK4BoiWcwZfKuJouwHhKxkeiEqdTJaQ2ATYWehhiJ
G1fpuSFOlaEwhM8snUPKIVrfYZv5POAeKO9EmHtz9GZZPZaxoRAgPzxbJdAM+FRQ
1TkaLemm3U/QttS1nwoK9PKMA0gm6OeNkaQhbEef/4TBJCAKlJKyer5Cb+UR5xgB
9lIqq1Ku2i5LCdchW9DuGHspScC3yXFghxNmfgF4bMVRo5LvafMlh7KaEdeqX0b1
0F7GdU1Wb7lX9Peu/tbB99ScE49HAjrqOXge4fzkq+JRoJUUYu2/drFHliTHOYvc
qifgLyjh/w/yaz3y0MlejbYB4rXIWfylweQpnN234zgsBUnEsI65wLCWNPVP94/w
GtVWrOJ3EO14J0+Uno94dB/pC3ZI/RKeSqW7wxzAcis7WdA+qI5Awc4qFs8sZCrL
gJl8B2u/ezuumvDsG+oHwkxs+1OJ1HNFzSCmuh+5tj+vAOSJ1rJts4m+Oo1FNRyN
vMg0jB8s/zCkpLCzUkJ0thZaPCngMD4daPMXJ/ix2HzKySQSdAyDNEu+mdqjMf39
R5HRGoYucIRIzLzf7XsO3J4BbBcSGjFr1cAU5K3hmNsZNLdoH0oS3vYRwrUPIwuZ
R+NkCicotGBUfsxlk7F33es+odzx+YUIshSv3TzwQ+3Ao7aluv3Km9GNe9KC9dy3
gyjgxEFSMMMWxMBUt9xsbxbfqVKOz5urlLDm3N41xxR5V00Luxy61YgtgEN5/YLW
hMALJL0s5Uy/W1JpPydBSB7g6Hf1jyeIglvzN6gUaat0nkxoeH9Keq63BBjyq/C8
Tb0rjHc44cp5o9+rMs46GKeUpiN0LMLchn8evwrLPb86w3tIiS9TvewmSLJbaFq+
A1xbngQiH+1u9CFkhZRbhgZFVCpLTfr8rTjNXB/Cnlq8rG93YRFOQbTtTCwHn+Iw
sziagByk6xP6BnCU7KwTSGxlHeRgMq0MdlEHJiXlxv6I18vmFkhGG31EnqJbVvRc
zMfEnLniMwV0k8AyzAJz6vXvz8NJW0kD2RMWkkJXCl+AX2eDhIKFnGQO/WRTLptL
YlMay/AK3VUcFDeohavMvKTvD2MeNEiSa4gpz7PbEFzKNkzDrapguXgkJxgAF1A/
aWMchNOzn9Hnr3vMpOo/6xk8ZQ8CUJP+MnOJWTaCqHD3+X1eGvLBZLIjtDdGIPhl
sOQsTlhbtj1IA65AVWMTkpmDlwN9iWO746A1sUYc40FXtJfF6lfCNMW4FgBJS6M0
ZfLg1/1nCsYiMo6eHK/WOtQbH1HRzBQAi518XpEq1KtvtVecYyG+QfR8Wcs5D8MY
hAFDfcQoS3UyhJ6s7bVLYfiLgfPXvIoG8exr6IEjPUQN06tXws0Z9uwfwWkYak9s
uENGLKSY+7ouvNBg+OX6kCDM8vAt8QMDG3zhDiSV1p2I1GHRJ4zVF3+iceQrQCx7
Y7UkSIb/rSlsyM2UuT/RtQ+Lz9M5tteCD5RUzKYqhoD6EdupKhfbAlIUmFO+/I0f
ZTPgC487+3Bq8aR22M6kTnaoNfTd6D+lVJr6i3Abfz7/6YkMLpHQrA0JJn221has
5oHRa9U3zQ5J+RRsTm43o4BMVKVJBkwg8lxLNBQruRMbC8xOS8gcXqL/JZTvsxIR
4ri3wbmVbZnTlFjEM9SXVnr0TgOC8ogltqfNf1CqCbGvwm510DHA9ubfPJKDJZ0L
NxE5w4sItz7meLNFwif6tRY6YRFLzzNY8Bo5pLietrB/KxGGW5bV/sTzbiq1hexp
V2TRychWCv/SUP+DMHIzBOy+KqcVho6DXmjUWkh+JtTbvIMIWZsRE/gfsJkYQooU
MleH8IPARWMKQttAW1Ba0UwFzu3yl5vGg0036CLJKPyW4M7qYSXdeFm2Ff/r+gD8
j1QXW9iniOqAS8pfbvbzcYkR+dXoqb8tmBRlOGIsvrFCqfdoTNLlkKmaF3AM39gN
4LSd5Uxi6GOGMJW01pmlt9PXp4UUi6uC86uVfdgWEMNQTn+2VqGztrT/ymgImvPk
eLcVbGav8lXS3P1tk+nSUuN22P1+6VhuQVpdvFui4gUPiW9c/w0vFuDYXpEolU1l
2oR7kEOf2lCe+sZbtt5014T5+9NFrOiz2DWpU0M4I26JkwjjqxY6USIIMdSNh4gc
JuG8hkAdwSj0Z3jzJ9NFhefAxjtwv8aJxTZSiayxpMlWMV9hMe52XdtN77OG6XZS
G19yQq13nrPsSFcLDzpnLUrZI2d8HMibjd+16TsWJzaRom4fmUf9bVndeb5tWQ6X
BaZTLVq/P5LukuIGvJxg6Sw/2ao2ipcufl2P59/XPk9OJj1BBTVG3DqnXjN50/bY
Ih+b7J8EIVbudl7njXsTsFs7K/tieYbRKHBmPDEO4llJCaNMjeW6DBaFh7TYqj1h
N0K3pcyvl9adzJV8EBlo4mwfzu+zCkZVjY0SxzFLARG4hWXyIygOIHElUOGTnfLU
uQWVkj+AD2e5vq1L5Ha28Q+itmYZC+wAokyemayU2kPo6uxOiyb0Tu/+SAYdI58M
vAUgVvf8PlPBRCFSsoJ2zQsX8QGO1/lgAKKi5oM5SJOc1lVVpXRh9OkYyDTZsfpq
07eaLQxaKaSnhmlYlnyKO8Ko72R/FBvhGClP/DCSwz7zRkUR3FbVLUETDcV47S24
WC7Shn6+X6EuuZ7+RvSXPtxGL/E3ugKMQDiS/TLXbj1spnjGsZKmJk8spPg+yyOF
phlrWDIzngKMj9thnPzdUSDLJVlyaKuZ0+HEIMmj6BvoSWBo4+xDFbZo0gbXmzj1
9WHER4k7gAswRHRHf7GHr8WXT3znDlzjGs3s1VBFxlve+TLY5OpEMZ2AE0H5XVy6
sJRzPGCnzKeC0Tqm89ZfataMEDImihme6qcgKuyL7fUoh6OLRuUegBtaX9/C76RM
+JE5Te4ndqZJLtauwcaYgED0RrfogJ5EDVi5aLkK+8fH2cErN3lo7zaiXUDalOvI
CyKcHHVcDG/QC148ZFZTCbowGaDpB0ZbxKBBHY/+HJkedmqSR35FTpLqP7IuGJvB
2oZiagf/aU0ysCFTLfFKpIQ0GhuaBSbDg8mQZW/RliAVo/Y9pL2lw2Sp1YRJntXc
Fdg9b+TUviSraQjUfhVDoOndh/A5iHcMUnietQPh3hEbrcjtEhlI/JMAVBdiYjJE
A+1/V+a0HGOEjlgCzHJI5Ug4cCn6g0HEaXaBQ+wd5D30quuSquR62+otR+IyKgN4
il+ExO3DKulM5pCoLe/EG4uRlm4jgqRmHdz0b2eP7zGm1gRNsWcpOBQh0QKI1kg7
yigm2Rk8BimpbF08jOO3JTM8rI3KG4WGA5vqqcLB65EGPdgpuhOycil9O3UBo+1g
QDjyKo54RA1r2ISzmhZz/yD7tu64N2c0/oQzV2lqTWcioc2bKa6XMQ31k55/UPCy
pzHJF8Go7MKOtghY4Rz/1lCyo8DekUcwFZMBJmMOAXuG0hQhVp667garjR+1RFGL
Pqf+TADcHNjq7Oklo1kaZVSAA8TZlInA/BGxgsJRJvDVXQdgMw0nkqm5ZLkIwfIn
nDYeXcl/F1E3xCGCFsa9S8/3qYHO7a6xxYvBDXLVIiqCSx85UNVGDx0z7eA3xd0f
mo1yMGgz1Eqeuss7c+i3I1TnWMORKI9eUPM9I7GFAAuxxJgDFAjWRqxldTxz5WBy
2m859v1CPqdCvfsOgu45KQr7JEomQ96KN7c+/I7LyA06yYct/dbUg8WzcHoAFurC
g8TNl7UGsPjvnFzSahjYxhB4kZA/lmPm8Sre0DZloTbmI2OrQeLxfTu2u5EMjq7l
GxutZorixDHdLs8qCepAqqDUdXxoB0TCdXQumCXIwjz8Uxy4gGUGW5u6DnOaL5iq
ya+38EX7AuL1RhiTTgtdtDWDEG8RBBiznvL5aI3hB8nyw3aSJ0xGNJimyGZl8Mvj
WYxBRzkbVlfXK84cMzeFn250pk8t6BoJEvnfw20flkwn+6xVjc6sCjhR4zc/MJjz
1kM91+a7QZ9uZwFxPZplDQldBwFHI8c69V+34M+r1hCCOEykOlZKd1NqeoC9JwMV
R1jo9PQwxReqjwLnba1CHON1LKjppNA0Od/IuMYb2IUHpRu6a2sSiAdQ4nEfUzYC
cnGL8IMEHHn0WHhzMhPUKgLVYOoNzKYeLCAuRsJ6Tzi7kC+KtATR5ypmuhhkpXsu
ZWnJy1DzBcNVJRuYLr8L24nhDoYTsVuvm5wUs9ZLEIlJ3o/NVhjqyPJewtsH00qT
WYdTCSkpGvLlU/aaK9FWK4VPMe3gL5Tvw/OYgncu7eiRvAbAjh9vX/sMzaQi3qah
Q6l3HGXz184Qs77ELQPFl4BnsMdgMh5YTrNIECB3xN9gZ+Y7tFk/1PdXAThP5cqw
/rqfYlK6vuu9qvu77bjyf1UcporCt9vR6zFS+ZCYJqsGaBzeGa6L/zxy6WjAzilv
CTu3ymYaTuIoh1HJq+YX9U53ANlaCftsq2Z298Zu19p5tFtCl7rvDt279zt+d9sb
LzBU82hiPNce2tUccmhNvwlV30PHptsl+6S2C9fUL+9l+NiVtYPJdzYBKjIj5XKA
xABmPL7VohE8/vgkt3gnwycul3McWZfYV6GiTDIaWaQrjKebPv685i5f4SNcBQxV
cublu9aAv/QKzCyLiRwGEYmmlstbeS7oMh0dMF4o8gUss0tPucHN8BZ9a/J4Lcpa
/h2nIS5bnsjx/+jU11axP2lVkV7dCPYT1iuSwNZpscqzL9zLWIQAs2xxei4+cR1i
4MaXrbhryDpqI89RPOqwHXV2jXvasVYz6DyLp4sg6G0zMa04NILYe8j0SV2vC73K
bIj2LSUgLYtyVr6fi0n7v0/0NjfF+eoqSh+pq/bDsfXDqfH632wy8mYc8BmgCu47
0KPxA4wFXuGeqcCxXkxGsI4SfR+40eGlOHNmYUwCSAONWvN9Ap0P+cxxJbmEWbGU
drjVZLnx/TaSe3Zehuq4k19ODCj+JKscfLAiASdNtuOqbT2ob6sCv8QsreBFEUO0
XCAZhCA69ru8Ia6VD7reNiFsQcS/hgnew52iFbkcn1iTmpcsnITD36AbsaBAfAMd
Ez0JW/lrJvl2Sjay0gQsGCZkQ88V2YpY/rs70btWzbv4bMX0GTDBaQmGwSKwodxk
huSCE/0FZtzYp+8HdTz/9VUawvoW+dYNuUdJ4JIFAh5jS9YOChmDjYWZQkJWVyqN
wfo222p5lg1fcJ2WxErBTXGFiOeP2x1y6k0kpF19/sAxAGoSChCKmHnquCP4wAHI
1JTspHN8ZKBg1hZjYTQZqu6pHnvLFRO55TXN0mB6OXFh3vpgan+1NMWo6uKApddk
VyzRUKjzp3H1YdOccvVcc9AuGGR42roKiRgwfASqJZPidmruMZV/mlYc1JRhp1zr
BQdKF0lzj4yXT7GbWn9PpTiCXBkgZ0yHEOr3dZ0vMP7IrS/KlRzSniOxDbhF0NAI
l1sOiLK3z3oD2YHzROOypUPbT0MjUqS6eiT/+Q0kGk47Ww8W5Ly0A4Ypc3KIcdJ3
q01rCACOrRMdJPUbqu9MbY4yysU4s83d/RGp5EC+rIpGVE1ZsgdAb+CCSfTlzpFN
874TSnssbX4D3GckDw3T3DripRlpIsatCxMMiuqdYI10Z84IA965w+oqquL4Zs1Y
/1+dLP37CVcrSn6QUM/V3Tqk4xMUhrjBtt2JuDhd4Fe4m8mriUrwNwkTIsOaLo1G
PFMx6F0h3WDoAs+vorymqvNYBS3kO93cToos42TVhzw4WmhdGXdZYBD+TOGCFpOS
yMfPLwwoX7Qsyjd+ZSHpMv4YdAk6rDJIO3tyjXui11NiqzzyJs1ajbA/OYe6Ov8t
fE1xXDvRL38CBakJDbDzjulJTgYHXhVW8q/bi7NwMeC8qUjmQek3r1XP8wqu4/pZ
BzetfLUBmPJVUaQM9QudYbZoJei/LAZwuRbIux8e4VzZM9/UGzFVV7k2N85atyq9
ePXhDtj13O/jNxWvd0Fn3Uq/BjpceS9m22iXuKbpSlwAJ9nuIXDzaWS+5qnlOYUw
3RQ0E+z3zj74REEQ8KvZS3PqhiyO/bp80bPnXsZeLrzfBZdSyHbxMYyOfFvkxkse
u6ZNKxJOFRF0BesruY9llCvMadeq05xfMymiywFpyDo85mVaHlXNHong1MZZkjYg
W1KfcT7myYoA1BganQRk5ZgEJEI0lNGDJqvsyKmmhXOU+S5JKI5LRky3JL5T7pJW
ealnKKCcmiqt3AgKeWrOVgfEBV6snx5pSB2PmJ/db9XpwcmwaxZbeZekneR+GeS7
KTIrdjiQGm7iU2VzMfHjYJp6yd6LPg5xqBV4rQluxqmtvR6F+0j2xvHGASurHlS9
xxtle0+tbsh+E/YVdBXOI49r2LYCLyiJ0XtWoQwKlTc1E194nmmo9Y/X/SA6msjz
QfYC8+V+pbNP7Nfi2Ze3dxi9BivTLHWE1Q3A6/8Q/ZcOlERs2kezllaOzmYwiyDP
LTDmk9IaL/gDayMtfD9H00mWjMKDiXhA+EyAAxC1jgxAQGxj2BHgA5Y5PrFOoMbX
G6GtQEKyfqfJbSbpzyMYk6xFDcQ6nWJ2xOgz2Ymi86RSy+LDhejpcEFjxivJITPl
EqdGhXQnQNaTzFrgexA61f/8kV2pncF4HG0qM7dbgtxc8EXaMHW6Q70rMXL16ptT
oQMX12qt0PeaxzqWeuymiadDlTl0bDbc7yKZQuyDBbjLPS47X0lXId/IIECy0InE
vWnCfLabKvAhmyU/vO2DKsE/WnS/fNlzYxMA2/BdfuZHqf+PzAKHZ2YkLExVjEmw
dvfUC84oIB0y/QwjzBIsgVCUdyPA7iTalHkloWSM/CnPzmitUFs+22As2Vu4ebsU
m2gLnqIzpLC6PRylZL3NAyRbX/qd3vj/Yu9iTG0XhjpD67p4XjQZNZtpSAJPI5LW
R/zFzkBXvs4yOLgMHwGwXFCVs8yDHPEhITyoo1g8WH5fIueU5/zm6LU7m1aQjGjF
EFFvjxVYF1g0fmJ7tLkILSnyL6wLsGy4ZI6VU/Kw8OtJH677Lgb8wKN3tIA6rIbb
c/pog5tJc9Hz9kkq2Hrj8GQS0Inkl9Pj4TNkkNUkX+ZmygcNVegD69S1bVb9mV/Q
UugAMk38ga9sKBgJkndW1GR9nQ7vFtzJPq1ORVwzZi3XqgUFSMNABSALnY5wKjCV
pdOiE2H3ja8r1cLvOifXG52C4jLYzI9XBRI+MaQxJhT0Q/D8WVBTs9xk/bTcdU1Z
oYdg6YwKU5qOLeOqfvQbVT3wmLXre2EY/kAAQihrJ3/Z4GhHf793EaKYlbze1Nch
I+XL/LBUanlsj/R8+u2I7MBsBd91fif8LkhhCe48Iz5TqWiL848urZ8pdPLwf0v8
eS2ZQKgGBZ7RD/LQGghXXfB9TKMKzGsL3SQ/wMCxVmI0Zb/fBvKS5LMnibs6Kh0d
Pt242qKuZCEFAxFLI2H/SX0fo7QLyT+yE5nwnhkOpm/3hR1aRV73TvBvrSPuPNpp
x/R7ZavANkjpze8RBJHkYyfR18XbCUSFjcDWsnnyqAQ0gqwPMnRI3poCMzKsDcl1
E3v22G2QcI5Ed/wT/i8IRMSQ1azuAqBqqt4NRChsSRtfGrhXPVg6tZayVf+xdPyq
btGdFzewKwg1cVinRXSkVFVlrorXgmy/yxSBaBKNX4neCov78xrqQMO9pHmlhm6e
b/CmDCQphl+VY3Wc0HqhPE2hvrGjzu5S2ZmTKuc8A+KIswra+O/06BhTGhkjx53a
+binr8HCdjH35+bVu8HZYDoKCgszgLcqB81/CT8p6btNEhsf+LVXA5AWEK3qfbNB
uojb4y7E0vydEG/Kzhr2mRu08tFIJP491n+n2M8FjHP1hARAPQQeaG/DCh5UPA4e
3+hTssj351R6IrEmOLAlDXj+xrf/YPpN5fmgCEkoP/CFIDQ72k0gM6Ue97hjmyTI
JjfkdEgDWq2uZCLeGgAyrx6+xcgASPFEnHOGK2LbIGpuppjIbs1AYMXJk/FUHMxt
H8BiVoI/RC3/RDf3BvEW7A3GzwbyJ+GDe2SyaMLuA9v8at4xcCFVUiRqph6FLMjj
4iNnjy9UXpo9RmczUQmv0jG9bLjtv4LSuYDf4yjdhfCez4EiFoC1AyHQ/9/Htpb0
peKsN/ez7Vdxtwn96bikzXJXNJzl9HMP+6QhtHwMwN1fwfqslF3xFVcEIDOoY26Z
l/WbCSXYH1q/vB+XctXgmBsyNAnnCWoN58EKEUP7DJe/CgHT+AccHu8/UrjkIX5p
QRKaXDvOILUv2sO9VpKRkysUidcinbYMXt1XB7SW9R0ouj7TfJ2rrOdgTYUx6WCz
LikoASgyLR0wfqJC6aLZVylo2T2L0vSKRb2MIzuQilgQx4K/9jFqjSHoZ/Vdr+bj
iXAF9pYYIYf/LHzjBLhr8S4G7Z8m86MrE4+7fq64NrQz//LioL4B4zrjCk0DvTwm
nG8Hzqzf5P2OkZuaXBQrcrN1CCZZ2Eqx0Njs/tjIKNxW68N0cHCcKVih/tsy9btG
Vl4QxaEfy4fy6PQ5kD7j4iCx8x7qWYs4QrXqJGPj9ueatK/XH2Rwb/ZEBk/juZNO
0rSF8FGVzHL2FA9PBw6f/zPEx6WLe+rZ2Om8YryE5Skcs+LdiqmAC2B5ITa0ySYI
xWjCZ3BNvw9WVTFg6WYmsrytFgWsxz3brbPV/t3AXqc1IU5A3Qe2TmARncA4/WH8
U/xZodN6r9TMV66lnQfWaMN8rvrAO0Q0oGa77AFxns4Q0OaymUg3tHup8C3B5dYE
hn+A8OEQcrPRMuNU5PhDOpb98FCqzPewGRlMNZ2OM6l6DnN+r0Ki6WaKZN7KJISp
apmZOSolPey6f9SCcpfQYiZog8C84a1a962sFlOwZScm680c/x0cdJlK5X+Dttem
ZKgZgvvVfPXYP/BC1o1HRg9uueEsiW62QoqyreFshw8dG7rgOObN5OVBBc+P+8gc
Ivi4ewfS5y8zOQMQizyVzwf7Hjb4f3JXIzJd+EEqGNM54bNJ010xuP1ERPaJcX8P
imjf2skIw2NoKwfq2rXH9hXM7NAN9Y5RjDOI7T3oQQMRfhw6MjfTqURouK6roCfg
cubJ/SsT+9TlyeYet2/fSdFq6ZOl6IT7QBUnrKKuPhJINjAz41OvB+lvE7CdyRT8
a6sxkvEZS8eb+h1QbCBrEZS1e+LJ97duL6K4zq3jn14DAs9R8J2619fVAB0PTxDK
W0e+aGSE0AzXdAioukiIFxrq9JRjzTLnzLpmTcc4sC6OxneOzYWyMnejqj2A/WxX
7stjk0k2lPnbLKUfCtWSkt6WbFTqWdrlyG0TNnSUDNit2US+wPQi+nDVZEPXEc6J
p01OtZPqLnCeTPqpy/WjTKbRr87epgDDi3r2zEs0bU0aXyDhKsaQJ2JZSoQTnAa6
zvsH9vSEIWti9XtIm6A8WL6v8ruiImgTViU4aaWjKVRBBUecFdszCTmZNEDZkORB
g1+WGKRQF3OlwGqNi2RDVclY9G7W8vWQUvYk+Vk7xxdch4HEtwk8kBSlUKTSQ5HT
b9fP0F8n/QxkNgOAwcd7FZprXP4GMtt8q0KGcm8dNAYwIb1lz7saUGRMc2lfRLjX
3zinxfE6+06WVbWTIaAGAlBAewMj7D/yEzTdPqUN4QLKYZy+syty5hoRzyASwfxH
JP6vimosK0JDlEyCZBslpQ4d/WMViCTYscb8C8dYUCapbtuR9DwaYL9yFDcvgRxb
wmHhBZdNCHtPZT/R1vtQDMRUt1d/8M0e8wNOhC5BIUgNZUmidA2W5wuI5zbsgwm1
QziZYYAExJUNxWnjfO6jU2Bo9nH/aKahJZRskUx+j0+vM/kgcNnSI6OjRrUk4aTZ
VdcsN1JrtgauHXlVQLQ2fnA6QA7oR3FDL1X+9BirnjsFSctjy6P+CkdcWgpUwWja
RHettyHX8FAZujadC0a+v7YxCu4EWvs8gkAiPJH5d74KoYOXGaSN+9CHgt5G4FEU
ZL1ueXehKSnO6tMbDip0nPbbg8//IyhBxeWeDOYOjkoyBS+MDuJHLBE7yIr3N/5F
CycIMS70nnCorOdqOf597eLDJMqbLlXQjRFwQVp+8Chfj8KTBF4EhS8L3Zxb8jpU
r9FdSNkS4y7E3Ny83ba+355J0BPYfl2Sqw6htr2q6F7UgBvuCFEUmYQLUem2lfEe
NpnQJWOgzPvy6n3aZDVkVx0u+BaNdKgrIGYnKbbZUhHikdXJ/3GYdA5MXKFtApqc
wEkQeAqMzkOlER4AKsyoLFI8DZVBW4LFtOgxlF8ktRsBZX2vc9jojUrY0ZU+Ep64
JLV+JuOGwaa8MwtVdQFb9woIm6aSacJiaKwgWTpvxWK3D2NQTAqCaesXwCD7m9l6
V5vm/yHgQcQBRb+nRTAcD5RifqHOX/+7Xgx2UGrUUY0p9vZMbY/1esvaNO/XNoh0
cjG/p5CUoQGc04rfU8W4daC0GZRESmDSTism6AXIZ5cx3exHBynCBWQX66xB1epz
kZ9Qo3Kh44bJ4WSgkXiAJ+K6/7eaaE9DQaKvFAMnlaL0qjF1s+XxVrgEZaQD9eDR
HuzEdd9tb8XuvhfTONJPYGFjW7xNmxsGCFvpSfyVPmqJcKE3Lh/5EmTWO7Q8OLCz
m8gPZPCokJOr1cyXdE2wDuS9WCphK7dthlgk3FWSw6mVzVcLjNYVOG92T35Jx8uh
SSiLkwhVfVFreJoDyB0+9mTDWZzc0nn0G8WIejSXiVOYukHNXIvSNXYuaz+T+kvD
uYyL9QtxhrGmoN5Vti0ne0bX0rVj1QVVyDEcIXTByH4yfN3jDJcCSAyivctj1sds
xoycXXpvZ3PW/PUDrC/WWmUZBI58bs/SrJ25285LYx/MhwiOlTu4047GNKEAUke9
5TE9oBnE7NPrHlpgPjdqAdXmzpPM0AuCKmkDgsTMi5xEriMGHWeCxcQWDRi39EY3
hj8z/CgFHTkXhkkW5jkq0hwF2eHu7m619pUOCIXczEvH90BRq9Nya/0/boxPGrzk
GdjW/XnE34Le0aocpw6JxX9Evo3MBZurYzWon3EXPY/94kjgTvYArIuwzdtRzVZm
Pa5Kv6OJvD6nE1j2f47immyBYG9fQFNkvH5LzH2W+tfUzZzeDmNmt9crB3CJnusy
QiY1GQhlIwZDqOgoF5W/rGj2CO5/uRHI+URMbltFp5RtJTxEBa97j1htWjervZiL
yQruh5Yp4vmbfTZ30G0Xi2ycSM0SpzmSGnN8UFk8YVMinOmqlib+H7mcfyhKAjYi
vMwXDUn42bJcmBChZYPIhu/mb0RbXhFgsCj8RusnxWtm/Hc0Eh42+HY7s67hHwaX
WEk0zL4ZC1yBEmzXlfacsJypiHKf3mM/IQUUJZeI4kKT2Eqxd4hcVKx51Y1iLmHu
0a+HmDZuNlXdkzA/9qctbJtIZiWvA2pR9USLY4Dx5dgOv++ENpq5ylTixKclESXI
OazDudR8s/Titwqal5UHPQ5mB/K18D8QTV/P2rSlNQIwFCM7HOR47PjNHF87bBDs
uMDiuHBY/klSdAcjNtgbuReB/CZzKDrag2uTyfS3r1taoJJAiaaNHWOTJ6Y+EJJ/
5vbS+MSgAlhESJibYYwR0TH0lEppCWlBYwkb57yUp4CJ/IuUFUhk9Nj6jMry9ugc
jagRAdOVkMd/QoZNKDLiD0RYN+HmY6PZox9gskN4M9gGm/FyVbBYNWNS6bsOhXFG
a2qLFg9XY76llivPUdbBQhciNw1futjbgcl4NoL+5YZUS+jERxy7KS30/gnkJPyA
pBCf38imRNwx/FRZQez4uOd4dt6vdzTSzAmqlvFQZNFjgxy8Htzxa6QdZe+wYsMC
JFCflNlddisVpcKImiBqXoIOM53RITXQB6Sb3Mi1AsgEJ0n32C0dmq+cenjABZti
Yen6NA5/DhKApBjEMHGcTzmcF6ytaz2J0fVciz0KhyLyuwPC4hLIBeByDpuyY+x7
edaKAE1l07a2TjmZEqHBhd+BsfI4kcInGLpn2qyHEoTB4kuCcbHalsMLu4AJfbiB
Uu0c7WyMsaCuNeTEGTDZ4HR+kMEPDwi6VzxJzo+pgistIJhcG7cxz0C6UUmD0F4L
QEwwFRIXx9MGFmYff9chBrPmAFQhSShTxN4189zoCa/vrNu0aSAA2edF1NyCDZpe
MDD/BVSZcpOluKNHHfAvbvMW7WvdBkGw54aDCQe+Eec55a5v4PVrJl965mwvASAW
cmk6osUD6w3o7Qa0dEvMTFNFeUtCsidl3xfm5lFA3lgfdXGVsNv+A7zxQ6oLCbh/
0hn0/wmXW19mV1Ayp4IX8YXzgILRQAi29WzOTJ40cx4seg0rWOxSOt62l3mUTBCM
8G8XpT3iuxyWoQOB0NEgJTGDMXUBhHHWxNCA3ClOButKgBnjEGkqYRW1M/OzzMrX
P5aOH83+LOVTB4hnk7nI6tlWN3FklvlexZ3DosVciVnmPHBeQeg92sCgLMA614M7
1U5ygpKPWvqbkHR1lEEbnySSDcKl4r3P/pQeUNFNSUsNMEGz3z9bwbc1hwJvVOc0
flEKXECRTyUPpKWUfLfJjsRr5I8sm//lyPxo6kUvcKbSWwCUAFmy/7LN1pK3Wq2M
+hfkGZ9YofMMEEW8fJ11E8A5WSr1d4yn0rj/rHAj08Ckyj2Z2lwKZyaLnkvplMGC
KMfaKtJeoWThRgzwNyhDYcWF2NI8sQmwDFv245rIg17bbh877hrzRvImuX3c0sGX
1Id81vxygT6jyQJfW2Tf5EPwvcaNQY8NaFRJToAKWq1BjAFNeEtj+qDUTPWov9Y2
rC+l1FNEATHIC3PTFRoagqB3XOZsRZsfOH//4Pg2W8/7YVi6AlGU52QHPvi1E3jJ
NmPePqRzVKA3ZEfo5oDfz1dSrrnwIKpf4D/qMMki2htd1kVuL012zA/JvBfCzFlW
jRR1LgsWPKWrPEpB+f+aDsu33jR0PbgfoY9GFmw3iCpd5Khusm2WsHHFLwKV3RXo
/yovvOWaWm9o4+8DNYDAKudwPesXRyx2tBokV12IBPoYx520XEIyoeIjydk6zLrJ
bHOFffBFGXA0cRqsf0RVkF50qyQKbFbOCw1PHbDiFPRAUzwlxBNoKkEB+mMG6YXQ
ha4g/oO2uW42YBEsGe0ZOpVzynm5Z03iWReUueg64vb3n4BjZsv7mCeN7OyISuQ9
kaB3/yoatjH18X6saSwjQ6+PxjZs5wm/uS26ZJZlNZV533x1yUHQh2fF6Xiw/jyG
wXwIuyrj6VsJfvXGH8nyQyaaDn0//gCYiTY0cugGer8XzZy6Yt/bTnqPI60JNP+0
vBvVE3RQScACXVT1Cpso6TfIcPesq6InrQAoW2cp+iLTo4YPK3ZvIytO0MeZW5LJ
RixDdh1Q02a13gQA4JB3rPQfa6BnIRK7uQiK/pHrI9Rtw41nnKXNeoj3XX3f79PF
iNcCLM+PKZpw4Q6BQAj1maF63mda7T8G85dTzg2MPu7YhrcpwYICzQ82vxCZhr5Z
HCByxEz5jdwCJzvtyL08fAZS38Z/s/R5LamSayYYdHQZWSKtB9Roykkogv0WgSaQ
X0Cv/tNdCtRGJtu1eA3oRYpARJDpphqAVC8kQwQ079hbOCd6p/T6sl6kjLUjgxN0
OBJvUYr+DDHUVhQaVeKaU81iP7CFkkVvDbibvZZRfp8FvZ+LiUHjiFFapGQly4J3
kmwO2TFdjEhVn3siA11L2/uvhdwXqeH4PpPSE2f5pg11JtmnI7l2aulPUsyZTwkV
hQOyuS0NrHu+wWrrgljgM+diQk8vZJzROU50ygNSmzU3vU/W4l18A9O6BdjDroSN
5mbr1+mrsheEXzTF82i7NzTI7ZKgOx54mL9q50ipT9BzA7V/K3i1yaG/FBcHQkUd
mbzzPvl8PFUcyHEfEZgfMylg7TsKcQft8q+B5piXxp0DdHyKRxXXAoO1rVyOF0hT
rW8ZrBzMiRZC4xZSYcLKI3t2O4aD1I++bRp6uUsDdM1kIPrjYWATQm9WPK7H9hEi
DTWUHDNzEBEioMDdM/x+BLfp7JMgYkH3nJVEhzrVoAcNgwOXCldRJrhJlgh5KSWX
2Q/YmRUewALL58e/YgO4IesZNI/rlzFXkQA0PPAhALbAYzQF1bl8g7UZf8hKQSAu
XssviUi5U1MwikbYL438BGcWnew6CIXd1p42SexeU8zpP87U1++roqBKDjDLChDJ
K3R81ISAN37HgVotoVs4iUDVm/mREsDFoMKHGjdG8xp47HiHFb1o4MZgbdqoL5Vo
Ta524ExpNuLEqTeQaVjlOefjcLQ5whJggqkiqeAOeHzVhfgOn+z3BgYKBWqSCYLB
EsNLUfBGvbupTbtR7nybSel1Q9d9q+2i71kmQFRUy28HhrCQc7iG4G59IhzE1rve
3f86Hh0ZrR14gDbu8uFus3W9jtNDS0MsDg/jGXCDSwnzvqY70jaSsKzqd4gvwuvX
ZteaVD9CThNoGKMektvjD9M07C+fdLzi6+KlBGgjrkn9M0v62bOLDoYS0GEknf2b
UI8TIL1cdHb3JzjBgcU60MYdL0Imea2xqaJ7qEeplXWtChHkg2ylMoDZmnDdhxr+
F7NrLcJm65NdN57VrjTjklkYxvXHrU7s8OLFrcGMlvDffsiRKTavVHbsq+0+gCNw
9jKdRO/lRmJVZ8Xx+8j3PGY+PBd1f92va1FtjURm6Wf75dA9hUzWvDlEH47xH7V1
EdEqes86D2+/hI5wB5PnXPEEBNRHEoK3pgty6g0NFMSVo1oO9MY/SqZHeIOSLaum
sbKexXA4PNxpce5rKMBr2m/KfBcK0cOtWPfxPMtZOaOyEU0/8veae3iQS/Bv7lVA
GRKUqGJ7eYzDarl0/pljsRb3D+i+0uTMNn9KmZqpdEx2gIEX9xKuMJyFxfkD09oV
DOvU1YYzn73vag+Sgb32MSS1XMGU83zx7Sm5LaXBpye6WrJpS9IANAqi/kdMx8IP
Z6HfTFvY6f0VlIDpflP2wFSkJ6RfoL2bZBSZl97wDJOo2vs8jvi4cMOBDXSOZ0SF
8VmJ1ToDhlK2PIzjx8xv99jcCUU2mafA1CDXS5BNpvp2V3n0DvSje1qtSBqpyb5m
O1xizuh3pAxI49KPEBI+a9RKBNDTY/GElsHeg4fSFskJUg6Rv1N5jxgIMMVAqFxg
zGgvfrSa/it5sTa4ulbxo0paA7LC1FFkFKt2IWOm2R74/9tCfNhYo+96JVKqectK
nnVPT2NdSYUu6F60m/2n7w5hy3GrwcGOtsRK4OCGM2Pgbxixe73sPHDe1dHj1nYf
0KspLfRhoD96j0wQizgIjf9WNVr0Io952JX5TDqACCbGurXKiywWExS6PXF8jl2A
5qaK2J7iPxFUA429ip060Gys7qgp4SrB9Ii3Uv8uwHuUEfkcMGltMlvloIPm8YTn
m/GOHPuK9HbOuGGFg5yVXFHYv40wfgsPnIZlqxrAvRmOrO/nYKtSoFuI4RgWNi+y
b6CVOVC7GrvsZ9PzqsbfFXm+GW6VANJhRnIyHgDxxQv0dxWLNGKmIBkwTEzikgNQ
X6ATbBRcyJRvOORQzDPigkyOvqJOwZykEITPp5EK50cY/h8HN7DJUCRJUfAvKiln
iXd08g7+80t/MhjZyj2d3qm5j293qdLV/cCEvLwxMDgA+r7JF87Nmoo599PG2xwO
VZQsGkIdoZwDVdW5ZgT6vdM4oJk55OnlM5XCUxAVZ66wLRpEaHoJ8mOKvSNmstQi
D97hALaAXAYew/n9TXU/+2e4yDMUMqBaIrPA+k+hmsQ6HRlPx+G876LMORvS93Uh
XSobxrzTX8gavks4tRzYg69XD5n1lxBeUBYf65AgOnpWGz6siXU4pqsRDnlITnG8
xTsmJ2cmnfmBWAOF7zCAqN16/p2DJ4IlG/TXY8jgSpfVQqpE/QPhfdZemrTbW77z
vHzaq14jilBirzKWWHQAYQLWmA3JvZwUIjUwlweHMpm055s6jCGbrKbwmw+zO0/h
kNakNJPYqU2jkvq4CxxEA+5IXCRWxUHFS7dCU2V52wXcdecVsknkVhEoMJYWSgLx
5CTOAYSoOARsPW2ITCvTqRnioH39r0OrVY0vMZey8m+uaBxST4wwzCd4OehidatT
bVKS37xfbksoNlGrbpafPAnOYnEy1nL7Tz8odQgTsAJ/mVamKonqfcinOKqOnjAK
/txB9nsVBBkxJafoo4nDkHosvrPIzUoP5Rqc6gLX4dLHB1xpqX9GuQZnOtXGh/yS
Blf6PdRvua1FoTwvMd+r9mJMv4v8gJ/9PYojWz5JxrAnRo61e0XNQW6Epl6d6HWM
c/p6AFWoaD/0vLJQjlAb7DNY82xwh5DtRB/wYRP9jibxNpEX7ojoPPkpms/PmlLD
grS4pT7QEx7XEANjNA22bAtPPHwCpXx7YGxIvwfUqkcPCwhjjmQgV5ZUmIq0/sO9
MOo7Fmh03J5LE+24Xnm6VumNGY3qQ6aoS5t+ZPm02fYyA+g1i8kqCbW0jUmccrSU
7I22/0jwTHntMk5NloueC584reBvCXMRXCrVlVBaF0j97MQiU1A2MaJovBnZAezh
auJgVfc+B1KY2xspN4VpbXTt9+hZ5rBNWwvk2x3eNqS0JIjJ13VyrlxND+ciU0wr
6u9eDjKzPkqCIOMSXTZ27yROH79vM0RmIR/VLsrLfijmPRtRiUmCI20A5SVE2VOo
MuwLgjrByVKvr2ejyEDbJt82trHjJ9o1eu4rePayguoju9c+bI7csPWwLtCo3/oG
Q/ohqn4uG1wnWxHo2cX0A8cIC0SYzMQKRgakXj8QfD7XoDui0H1wX7O3pnYVgYWz
/ESkfXy93nMAofmSmCrW2LbzBW9SrkkQJSnPPxZYEgFNHuS575n4VVzd4AfF6p8N
GUUY+fwU+NY/KTDmWu0aL9UH/seCrxp5gUTCjMrRFae7ioRX41lyhNob9nlD6Mfz
EWmwbUOlgl9plkDyv5rixd/mLhHC4wv+GKMUUGP6cxlv9qU6cIzZlWco94NADmbi
/FP5MGHV6gvcW0+fQzSCeY3Rg79MkjtQDdN70cru+3Avt4LkAKTCmXyXLgwc+HBt
5A65Qdvn59rF0aH6frA8Psjux14amOf9dSXmpHjEYLDNuoebD9wiUBygGIMnu8P7
bJodQdHqsYvArLLkD8Uu+ZJ4T+qEZr3+tSfPEzs6e/QW4/2fRSsirfHGzkNUxZot
AGuJ1Tb4Vr3hNPVnq2GOUGx4SbQ1AyIM6R6U5rcXq7CD+WSveZosrf8Qwd+Vu1Ic
Vq4Zg8bHHRMARYaGTCh76ZF2SJvsaOEQZ9Gm/ruktitJlE2bEHBsnkPsjqxztQpI
6LejWZSIBu8LC2JF6EueXZcuzkAVXYuPxdQEkJuzbiAX9bHw0kvazLutgTDRcQFn
uI9HlVe0PsSub2wP9RJTCfnl+/YWrm6uSESLWaW+/Bn07x7GfmFSKSXc/k4gWG7H
q0OWkSIWul2gZUAavvUumkIJgiN0r6T3Ds6AhWnp/op6UZG0fdlyIkZP9WRqb+qC
2lABpy11UH5rremf/jgJjQ+bz+Vr7zXlBkYO4Rbm0aVmBVrKYajYEf6yToweDKDb
dzjK0yaA5sAKmPeqa44PnLRttLS9Vg4tbkc2m7UicksSw8nHue3Ba6W8G8Ye8RmW
813BkzvCNQBNV+R3FSFG7nO/SHPGk93XKDjVKMnq5eKJ8WXnYd5W6k2jTKKqGfji
g4h93WYZnoBKGuEMaL4L1BZG0PTBBs8hTiKTYdzfstbRwdD0fnBDtjtocqHr+3j/
nQU3yDnt3K3ArxaDlRFe/z2vOlzEVQsiQM7O5YkhuY2ghfBhnx9odl8bVsQ3Pqpv
dijY27qc+SHpNaPuNLeQtTVg6rSTN85dYTlGRtAMBrZoLkFWEWDqJR55+CSVkilB
RYu7BQRXPRVxBj6f8TX7pzM6V2ZXgnrPPi2zBScnUqm9iVFRPFxfEiCsSdlbKnRo
cwANLih+VbtnLRGK0FKhiEFIddooY7B3vVYrizuM2zpVzTwOe8kaEIPR14HDuQZA
IVZ5RgZFyJL0nZfjWl9gbDNXglfiQ3CK4glHqp46gxZQIV3SigpHxD3tnQ5DYwWv
slkA9yHwe7M2OIEr6BBZCUB3O98jBeP9PEfd43pEzLJx1pL645w8eOm1+WJDYUPy
QE2UG4+NE7sKwuC1T9UPyDXwi2M86QcBa1CsZGwhwhSucwvhksLf60K0YyzK+Feu
wpnZVtagN80Xr2qvBSnlA516hGtHZDYaZXTWxL7TMQl4yl382gSR2w492ywZPPnD
O/HwSfglrx+2oWlme3gKwy9qlD69Rw/f5amop1gPpH9X3OJ2FH5TrOHnyQdKEP5T
oBah0/LmhuA9gEh15lLox3xT7zH/MMsFGl6Nd0gRJqhOkpvBFRnjnP0G9rrocbfO
5ztuO14sn/mWPFewyPla5S+xYR32hDogA9bEeNkXgzdTXOGdsqMh0LuTXX6tXbj1
YxvqhVfW8JeaARpl70gNa/tl/AukygmC4xYuWS7VRZ+s6WF6YpSmslBSyOB8205C
dmkkmgWLqdsWz/wmJNXGLXRLq9P7FIdSqE9u8r6661bHapc6xaBM8qgrjR6WJ9gz
hOOKOuiMTp7+Q58URn+PIiuPq5t2+NNG+MDLPB25k1F+3JmMgehxZrv+sP+vJ1Bm
tMOhLjeWyrKfQCZkXf1ckDZfV41ZR1rLU6I+nf4QDWh2VaRna1vdrU8BtKozhb7F
4Vvu7wDZzsl9N9JHebYyTdt5B9K7shN4UDLrS6RHaeAUxLb+4sU7cGWL8exUnZfd
eGIhQb1v7EM3sOwVma+/kHDNEgiit1KrOqizyparCe0HdNRILhmWnIYoDf7rZmpW
T84DMfJRezb9lbIjy+i/+drRsmjZKorbkN1NfqxXPChFsvxLUEaOySWfXpaW4pWM
BCMETVLfo2VCD1a73jE9bho7bnUL1Z2tpCedkaKkoUjGjfflgmrbcE9cCR+GS34g
BNj+SmVz+FuklqiTCSYB/CxaIvXWPF89DcluogR/lNB3r8vpwoEBUMwqek9zIjd4
GC8RkKk4b9hZuDOEOA5zXL6HiUOwViVYc7s2YDgzVnJ244IIz+v8d2/mLxDq8v3+
m1YPJH/oVgtVkJwxnzmEd4kTyy94O3JS87hvYSDLSv1Z18POmpoFTa/errXPcT/K
Rw6D8uU13qXXkh4DXEYEtlllFV5keyATBq8q1+MLGRNcZM9fQiAS1HYqW/0OUVfP
DVjVBVL5dh5jlfzHQgTxGjKcIIj03s+kboUt56v1Ql2FQckvUjmpsrKjZZIx8/ON
O6Kdd1P8MfEJhXbTzP/W3s2svnICMTUWbZHPVNf2GcrwHV23aAgWfWNHsQD35jik
0ZfborFL5wu9Xcce8WdTTMXhzHB6A7WcFSa3WvwQA8EXWjV10nhrRj9N0OAyLGHn
umkVwoBqG9r3GMb1Y5NzNpXde9zqX/lkEosezNse4XEmD+epWAsJCu6oAX/7Ji/C
66uE9CXaEobGyuRv6RKRM2W5QIbviM/vPGpvUHay3Pruo9wYSahLHHX8lRcrHtRp
NLOe7rYMZw/tXywPSUjv/5Z1SSPQWLeXT0EbHSExxvunLL/Ew5uWassQ/kQjYBfV
lf2wzLamxwKbBeIYMgD5rUu1L1KQoXvGWG78H1gw24zvVDCI6IShIQH6Iog5Fos5
I5ayVJLIfQvbtac5EUt8TertQL2hc0lj8EAgFYpRfcNlzP9jVfYNOi2w/cTsAgpd
eFilIS7OOSKEv7UwlrXTFvvtiRx2ZHLjVbI/nksxUBrbUCappj4FmYsEUZLkzGAL
CLMm5XI0QB4O8khR7c6OjbeYCBWFxRjkBXGMXRoaV53SIoGGvN+8fnZAh/z0qfJO
vI7THYq1UtyOwcepbKOvhtx1FjgYfViOJs27c8N5wxAFpBP1fZqjD8VNP0ZecSDI
FdHR3mYXC9UDYeeOvAEp0nXRBU6xNW+pu00Z/H6SPhwtnqAegEXg9RXS8Yrlm92I
hcceEygGXcWug4sBzwBmuyBhs720qdQfDA7AAHVdMWvwcHzPg/qPqJnDGxll23eC
9A0e4AiMJ6wK28nL7sj1KQfQJg+sELG+1ayFMBbjzd1rJmr/OLG1JFL24AhM0L1P
e/BJEgk8/iBuqoH30dfy1yCrNM+MqEV69uj/fDoUCaY6zMWVrLdcSaKBa+zeQz44
AvOALg+XyXQ0+1lIsRHnIEZO2Av2e4cSoK6je8HO8I89NMoAhtY7bAQaXV/lQ0aP
p94eC0aT5SgwB0HByn+DAR4Fu3+57yRawfhnbDb38iW6X7wsuFBfEj3BljricTmL
hB6oPGkB+aSYRREwFLUfID/HNaipYQZjr8Imp/213e/muHHFm4D+IiY/wYLT8q7G
I7rEyot+90DCLxNrX+jS/wHWz4Tz/juwjtygbvJnrHgj869SE0FPasIPA7gmthUH
8swNKr+E1ueGWNfcjrJ236HIJMSc3+4Dzph5jxVYqJcCOoDfR5wQCz8rTYVuhnYb
b+g4BT4cQXX8EVwUePg/UOYOnwUq99f9AP3YArWwzzsijZVoCZxh4C0IPSQ4E4G5
sLAySRTzKzEdBYV2HAcz9A0hV9u0dKP73tI7o+tY9tKyoyvrxxpUFbv4isoUoIML
5oYVewyEXgEny41IMf85hIZ5W6lhqh6mkf29F/Yzi9YIukqGPTx4lLWfYz7eHvBW
RKlE1Onjl0USXt+K36XXW9mSG4ZFfZz44wyIhyWB6mAdFUq9+j4cYlLEH8PhmSvI
iU3VyKI41F1T5K0FZxD5D99QPijvPNBQvkny+ip6Eb/Sdxz58zg74JY89CDyAiBW
Tm50JZMmcvAn467ri9sL12xAFF3//Tlfad2cgC1RV7onu3xr1ZbANLHQRskw9jSH
LzRvEIVRUMTb0oN9T9xagabHH5kEXso2ILV5Ns3Gj6hnCSStsddpOz7jlKq5y+0d
LZ1LsTS/udmq6UOyMnoyUcIByvaKNNs7VUW/fM4azOSj3SRLjUai6TqqPdpi5Gip
pAa8i0glqH4p3XDPH0UbDGZYYWQo5DniL0kqIoYoW0cK4xX5svdpFZZP7pJNirmE
uoSer19FLEd+7zDFqrx/IRablZvTBPJlvZAhTvZBEFO8GYjJIjHoxmL1/lqE9M6O
0RLUH+RfVLOm9W7ICenPnwDf8dQ9Lv4HCIykUwtNOvg7tFcOWD8WI0B9hyaSppFc
aGFZNb9eQfu6Wm//3+He/AU1TXobBQpzHxxGa3KZsXXYaRvvs/o8hGtDfBFFPFoE
ZGwXX4UmynovXx8H9+eoH/wvTbDKygxkCbekdnh26eftf/yLRjPpg1UBmaBBEsKx
6PWE7VWQ6ffjLaGXn8xwb6Sg2M8bYfR+tXJ8p/jpHqc0EtV49PKVgLvdrDmba88P
aZlKi0+kJv3xYSvUvok9qwD9gH9aQtsOG2l7y8EDyyzmmYIWYJBvno4/5J806C0L
0uC3U/EjuGu2gVWPn1VZDJIMg9EAbBA9SVtu0kvAN/k5KXFfi1uvr7xHmx+kADI1
3u3SlMRRyuaBHEtBVeAhu0v+01v8EOY7rHZy5EdNgGBEylR5FC/tiUPS5jamfjJB
zdNeQ+AV9pjKY+0NFX6y1X/xHPXAserJPm4a/H5q5zpCG0xOunq6h0T/LQQAzjkB
pUNhHga7v2J70TtQRxCAmhw1AO6qPEDgagKwEszKHs1EvGS5SDdr6UJqvI9BLBXQ
OyD60hinD30qxMa9L6Lgkvtt2/XsIpuXjB8e1mhT5azH6mJdY9u89xZUYqtHcvbp
g1f4sIl9kODf0kMMhgToSXsF1aMAjKNOmcy3TYDavQykYiF28TQ2P6j2SfP5B5V+
FtVPJhu4UeLEf93pTLhECg23dHtAZgdqahg6tV4Sl4t+HOJDjSz0zx0RLt2CeBpB
myn9BPkFkg5IloYvKFEv7MTgBUfN6ZMxwFEVX7M2OfhAolFeIzz5IDt822fqHcc7
APkxXTKBEuCfAlm035G66APvxnFmcdbOP5ZUJPJNvmuOYt5NrmJuxWTqPFtBHGX+
FbdSRgqcSRj22eD712fhs8Ir5Y5vAQ45EoyRc/YCbtpVGcxPqmub5nUc/L68+Zri
byto26Mf/wSACyNasyS0r4oqEHxZ4f3Al3Y48346nS6/ml7fVmESSNqIBaTrYDxf
br8fqkK61o7bgybD2noWubz8tVumWMu5pBB8i0KMvfRbChDzzWFgtHWZM6jf/jfa
mtowxHx//UIaELez8TaHjQIqm4FS6yw79G7xaoeGuKq2gVCGFVk33sKNIcRFP1o7
3aYrEBZ6XXpnXmRQsaU/SYrmvrVAOV7RlvIIRGsz7JU1DcDQFZ/ZW46SeYZcO4q1
R3CqCsWqZSXhhBZ3SlRu/OJR0ddzJXfZnhuO7nftsbY1sqCDJLYZkpvjqkMqtIcl
T2YNYeOiPD3BWrVghDjvqw3oPzEvnWKQPFUcxtgQ1Gzx/DjOFtbdXy5PuZV7gbBJ
YEo7tVrcqsmohSps7Z0zfys3BEOyI898m//isXRfTdcczsdfUyhl3IzWt9jrrwXB
2VijJDCUmwehll1JQodU8rXcOCUHLiAU4VmJjNFwBBmKl8Gb+etlulYr93OSsGgR
ZEhRrcrM4gZ1OibMMOtuianZSIsPaSYKcNdpVEUAh2gddOcY1Y+wkt1voBnbTDUi
xic9WdYGlKY2Q+lO8cVwSgl81z+C1RoAd81d5SGKAdwrdmWf/1AhutDTNEBo8euF
4TkVlEJpbyY5aRokQKEnDqUbvptCmzHp9Md1nzMsA4uE5Z6vudY1EU5R0WvRpIK8
cNQFZP/Xp9biZzGt1tD3l6bk2B+Kdt+4sC74dSbA44Ew8088cZoWBCs0rwtOu6DY
tg+oljsXYtbrm2sKhi0qLotVnl59ljj/655mgRt1ZKSmH+Ao0jzYEPNYn98USIMj
PjwQhXeosoYeLhF6UuTt5t8oAa017gcwiJLTbcpQbRcYFKt3ZhpgW36mJkPwVvJP
/wdgc4D+eTDjy5W7/dV36sKjb6gpYEIKOJZK8yco+YzNhCuew2pMcMSTVva3Owod
PG2VIDGt+51rRQbkxLgdr6IBmX9iyp9P55PmESUJhqOalZQYK5H+n7yAlJckmRdS
W4vZvdFJ5CcpIo4HuYSCJ2BddGpSrWA6d7Q1w+EaZJxvcUyTHcUDKkaZVfDXWpA/
ghPF8CobpGvAg8MN59Yu9lqyWZl2BD6SWjyE591ZoY3gzOFtRPG03jpjDB9Yc7mu
SZxnNal46WPelScjksxOCgD0YPq/xNQhDcCSKc833C+h2irFjcIXzAAzYWLGqueY
WpdFwGG16RcsdF0coCEIvuAInmCWlT5VtYxutgvVFGQxAV8hwyKc9KLLio9qUCJl
aPzDNuD2pJ4aja7+jLfCmvq1ssXazLQmtsfLs7obcE3IxMYhN5CbssULDpl3Q2tU
+K8wY+q+9e9/zR1sPGYtRawn32BLh7YAOq0XerUobw47kleUZgKkpuP+mC/pwBfL
vjA2vLaz80ZppZz/ARST2JPKYbru/bSeFEJ6Q10HwFVcTIpcgFSeBUWNyg+OYbAR
1jQkgwSyXGOuN53aMaIfynSKE9ww/HYB9OwSnWsxOBvUL2bIsZuR+GEoda4pqllz
yDgreA1KtvOYxkrxGCR1gGOhlmQMIUxrum1N1JibCMR6EhtdnkULbTFN6iyBsVfw
zhINUkJ62VDLQ9Vuk3cYMebX0/kkitNUv8Bj2gtkNTaI8UW9YggoIWSBThHDxRhW
gVJ1k8M16Jd8yJvS3C8eNXjK1Fhcb9vvHGTGQD/No4dMmSSKdIL1bIWPdozUSmXT
aPtrKI84xbs2R/zM6VFwYficqa0DCwaVs5F86k8BoknhcGgKm0sGgogloriQtagf
lBMDdQUoQOn91jd/bdI6d7E0RBGPigwyVFSAmicTI3t6v6Itzo2eU2FmVGZnJh2U
zL5J9jYpfSQP62zgiq0d0t1kbUYxKJyrpaRznxrSvmlBf/7Sf9wN8h+96dkTtTX5
uWSudDXsnB4oVtRwi5yWiFBT+26Q+NR2q27x0h2T6zL3A9wlTStC0mlAHzajYq6U
I4lEkeFcbsW5cfvHxkChCkvvE9GGUoX/dCF+bHiEn9g5Re16j6eLIzO/0cz59Kia
4NOMB6EZsknxzF+4tNWteSN9/4lWkF6i2qbNN6mZYF4hNZ+F9MUpYH4sBovyfjlm
k6aXVB2l5yLCp0M9TA8DJ+WTeczArVMSDYkOyrhkSdtSKsiqSs1KrGJsMiDaf6bV
cW+UQedgjeAftjmQ6gdweX0If0SgVxSXkC9BZuVPaubQaH5Kfvvh/O1u+oTDdyz1
H6NVKQTHcrzuBvDbPOCyMqWgEirqLkZ1T0S7ssbBlDhV877fQEIyQmFTD6Z7Qqiq
+iO95wnt8tjb1S1qrsi9i4LbwDSIzX2Txxw3Q0kcdTumQsIiM39NNAHqtJpGmnBZ
cIvkIJQT9k5aFm9Yzl5BWLm8YEW0ujiaWpEgBL4KbEmQzfhaJBto0VKxgRdVw6W7
1SOj5+LK6Im3yjPl/wWHOHBp4y4hTWsKoEdoDPn6zJzFLfUva371b82Wq3EG7TMX
aNj/n0K38PgAx29gQfZ+jg9uPDeG4VjAiQlBeKLPP0LfJrDA61BULIZ7A1wm0Nwn
eCmwHWopsYOZBkY2mY4nR4c31d3BQN+gOaOXBTjQ56EdamddIPIPTWszZkRQZh7V
awlylmg7JhPKZcKJ02KGfk4ZAwf0NS1o4MMcRm77WOTJqfttFg6duTBhBi9NfH7r
Bp3PfWwvOD8pvsn9eYTy73rZ5Im+v60niDID8DNoJlLSAgPbNnsccl3iVDxH064v
3pXcyhAzMNPqN/hQ6cpoUwUSw8ixo135jZDZeRkVZ5K+Pa9NlGExYEEc99HGJjU5
1cGRzrlC66rDUzEOeKX07xECWgaEBbZZ8z8mIGql206k2jgAHTZK9S47wPV1zaLk
IXAm9d36l/bs39o70Wdd8GtEynSZFmJbj9CFXhqcwvAPXTGkN8yGy9oivTpLtEsB
+vI3nLWbCxnz4taGnQtXIU+B6uF94MtsKqZ3Ra4Y6B6d37HKXkDz4pPdHpAfUQKZ
vqUbzw/9QedDncGS+Q95ZuXaIF/KM0yAYWY7UWzz6PQE/3bzDBOFf4Q1QfVu6FI0
NQwrjECegwzLnuC+eUWwW4oa6Dc8/kpRfzJ1XeygGmJMW5F19ikQ9CCXxaizcXEN
E2ovxR3F+rUg7aEZ1yYkzJ/IQuHOow/wrwwwGw8WG34qdgs84b38umgkTLMVD0Ay
ItPqFktOHk3I75RyJ6OyjbeiZj2B01CA0q7s+V9gmsUXL4DWVQov5dVoP541e1td
lSvuaBfswGoZHH56vOKaX+ffL2xhhLoEyFYJl/uvlBJyirjjly1gxzz9FaBKxz3R
XQVEWw37ESaFGx6MHBNTH+obm1yJlIPvAmGGGCOEBpgM3W6EQx8j5Dmwuq7r0arF
CCSsMq6VhGETx72mpMK45FvBCYQB6Hedm/nZFvp0nFToTISScsqzv3ugY/oaXoWK
ARA8cKl0I0euq4/XHt0QWt/cDzz9z4HPgKLNX5RYBodte4ZWXG41Or09pGF6fvM+
58RrTITZEMCggekWSDlwiwwgBLFB/WArsbR13IgeoKi8RWe7dQGsXZh8bMpI9Z4r
+MLVOkck4lUWGRBLSATMNBJmRE6paRLDEvKKs80eakecn7kEPnhVg61kNhfqg84F
d3NPSQHXYbPhSVkQo09C3csnkzodj53FmSnIMIP1ioI9W2fTC7jT3AS2A92PzCKa
21jzHg1rincmGBN/YPVQOdwn+Lz1rCfOQ1V6Zb1TSDp0UBsJDTVicqiC0g8FVmt7
dCI9m29Eborxk1Ez5XJA0OZYSPqpR80ixoMkFZxIUo3BEzK7TdvjKWHaytVxYtVu
HF9Ftf+b4BFEQ3fGxzY8ncfz4iigUVtIj2QTK0+GH6S4lx9iWtAZnl4cRXHBma+A
ity7GgVpgHRQSUjqssLORX0m0lghqbbAmE/i/+jlJOiDhmTUVu1vVhu3DhcusHpK
MEncsZX7miml5qNrN0L5CRRrrfD+roPZeCTBzqUd/j9KlQvF1/087HCkz9UhWpDg
W92GZoLen9c972m49da1dJd5/2XxryLQPUKkIYG/1syF4N6Wdbfpzp4uorWKT3Jv
4iAul6vz7rWEd+6Vms37rBkO1xOOYvfMoe2R51P+EFBBnzpaHpwhV98wOctTHPzF
xr1ZInp68Vy+hedanUmpIlpQmxeU3I0rlXScL7LP0QkW9o8+BJ5BndykHv5Zn/OZ
rsDp1UosTA2naguYmdgm30qpK3K+t44RXT5x1Ps1NJb+FWxlBKs53hS6/8EqDKxv
7kbJxs2Qrtl0D8XHc9JcgzmZvgBTExYtdQowGQzLwr6Mt0s9ZtFiO+aZyoJ3uebK
KX5wCNrFtDYIMe4oJUObR+zEs8wj3J71GSJhBo0H0EPCJUPg/LRDPrQ+juMxM8dE
7R36g+T0lUSW+8VbtY6Ou/K72FYXCJPRytKe512HUOQaUjgGbN3SQiyRf36vZw2V
NJjXka5z2dR1d6w/5h7W1w/+EJvIz/toakjo04WqeEFxqtgwwqehFRmvfPypWWG6
G11vyRzbL56WgqOMm8Iw7Z3Wm782VEyEhK768fd4z1TSHdXzaUik+MAT8UsbtQkq
HWqh9R/nBCoJdX7GjGZLu+Cy3UYXv1CK8/6NgFY2p+Mfk1KY1n6ljPOM8znf3VU2
s6SzBFOW1nrKMipxkVvxkZGYInr5Gobhj6s+xzBmU+V2oSrFyLHdQ2BSzSCkVMda
qKspvujq+0ReCbIltf4DDipthzw6vHVPfvAoDDZJKIdSRHXMonaViIZCdLkkdlUQ
8ELgPoOEX6nY/lgNKkPyssugTwqOBnZTJ9OMfCQ0pSORx9oouTSCs5LiRC0b+ogW
5Sbfuc0eOBRk0RokmTpK96mGVktLQUGGbeykZZ2PWuR0xpoeW3LSKqDDZ+Oehj7n
IFpt6TT033NKTP7ek4vxXkSkO7nfe3diIAmkyR+qfEMkaFO3NcJREapV7zyETxNa
3EPx55dZN9URt9+05x08/GTJwHL/Tdr07Ip9c54weaEq0exbs5lL5yd8HZXc0Vtq
4STq4Z1WmJ0yiexDY2RFAKs71qzDHuRiqBZAl9Bqh8+zpYwCQNY/xcc7IZHhkyDG
k3exWeqDI3w3J2dMs9ufyUzzzbo0o0XOgxF6RHUT+UEiCGc+p8HT0b7aClLRyuBw
9riKg9U7dBoVDmpkXqIuHyqIb/nU0jz88PRenSFALmvu0OWskgfAubBoGEQXfFBz
tV3c/d2AxPrKbeligedmZS3Vq2joTz63zkPY7FjiDX6R4jYb1QFD4QHsYgJYUrSM
Hz0zD4Um/CSkKR0FjBZASc4wTUXO/4CMa6SwNqVhgApsbCeUsAoSApxXik2IY/fT
TqterzV+ohKiV9HCfbpjeZ8U0Q26oywj3Dt21PSex8VgZU9OnDZKKvd0SjPOCFer
xsSW8di05HM+zTwNt7yWom4VrlskSALsbWuQcBdBMh6b97mA1XhYjqw9alZNr2vv
DJlcn6PsEYu1FppyVrlxbNghH9u6nDenLgdrmVniVROxkAbZ4LwfYcY1CkyYL3hg
dtYgmI0nntVA2QbSiS6svS89ljSzF+YOw2jp1JZbDQw7JCJW3/GTaLTwRxR1cr20
KA2QLRxX+Ten0ImN2CXrAZQ7e3sKSe3INETDuZRyWLBQTYmTkuefY8qkE4B8ojeF
5hOoZ9nkvT9Mv9P+tMlKBvF2x0IH3pcQVz0mInoQNPJGyEuA1uRhGAG3E78yb1DO
ouk9LfjEJFgGl4YcwuMq8hfFMOQHytRZ1hyfgRIjbcZCK8PoMPa5EbAVb2ZzY5/5
ufIglbMXXss4nq31zfEpIAVX0MUkIRufMjLN9Igbl8kGPSrYY2J2q4OEtdzMBLMs
8Th0ONUOAeDsjHl8uuWIQz7keS0yemGkJzuSSonM0HbZdxb6aSZipqs+FPwm40xG
LAeLfnJ/Jrv5CFCxyHvvfCLpReObdmAp+DmDet7oMk8Af4Vl1mVpfc49sOtGu9Y4
Z604oVe17suhlG1nMqIgSU7Mj73M2FvRMz/b0LmRHQ5xVQ0/V8kE/kU2ZdfetmjW
0VZ5kJ3sBey79ymMZmYigIv/KWkn4HTr3sxdQQ4BA00TfEjSMPMpHrXyHoPjnlAw
iaJXII3HjDFTqk3DgAx82JKNgFuOrYBRuh2Bh/cCMF+txgAv4mX3ZWbP0H+t15Hj
mRRRYYittA52nSEqmcAALGAlN0XzCC7Ass0NcDUS6JQ+jUhy3did+dUwlP9/w6Cq
0I8tNg2QhvrFzON+LfhUUcY843QEp/M296efjnrsIS7PEVKTeT5HcutJRjchygTq
PaLOelLOqImRI0Lf9I30HzOOoJPLEfuQn7YfIRYAbvDMekexOKICF+x6I+pe5s1S
O1pnpZ4nCzb/Xo7VqjbetaMgJE4P9+aSdOvAhNy699M/FkfU2D43nIyzI1fU6Rzo
FBm8aSVqxJKMBpNxRZS+phTTeGiIo16RhyitrJohGUeoZb/d1L6vs00yLQ5khpgu
kGXpq6xgtwrfWB01on20+l+J1p2Wub254r7EyisK2ydEACFZCzZpqxeANQk1Lx11
5Fk+AbUXjtVi6LuomT/JicchLnELzh/O/2WXgj4ccY+rESMpUYWj3jF4qe0Ms2y/
CbSs4xXpy3JLKW31ZgnW5pPgHAbtu34j2tAJAhau6cibCMaIp+g1bXplhDrOr8dy
UN5G4TKpqc42iaUS26+h/Dc9516xlDuiK4KYSsjXl/Tm74FiwzDQi8kfaFs7KCVX
gLNPokx2dT0CRjyBeoByQLTZG1/BFCTq+r5oafjYCjgFBJhfXAs7/qeVbTsZatyY
1Z23+aFUktoeCvHEcVsJ8NkoDYiHx7PF3ambu7YE3ky9a2rIxH1cjDtxv5CkBsh5
Fhe7sQfPdGa2jSf5GtTmEPqgrp8/sv0FebZYzZPmToRodY+sHNpaqcyb95LNEaYd
NOasoooPvost1SO2dPmEQPtT7Pd98nZC8MyB4H0cJ1gbUmUqMYqZHeDhQ0pRoFZo
LF66Io+3aSLB+JU58GJCGm9oKKEUvFEH7MdaGZHaF01zPgKd1ePbGW7RgWpqECVD
vJrxAdKlmgz4BI4AYcD+wKj0cjqFfmlK9tdoTuurWtoBL3Fj9jU4k+zIpmorBKAe
pYneuuPAZtLh3jg/5NcQtlCBbg7zGL+K2WlO6fqS8munujt9q9EgcHBK+s6Ma2mq
ix6WCT+1+/kSpOupfErmUfr2LvC8fJrppgWWKgxVCMrN6CYpRchiAb1osFxfP+7X
wW81VFhQG/w2KNSX6VzitXMHET35ghhbinNUjLhX3djVOWqbeNVltzrKyQw8GlRa
YN4cS5kZ+w9dU4jZvP7kQ6LQCLGkQ2q4zrBuSy/gy2VHqDJ06w/zOGBSXaYEjgPv
bxjNqnWwWj3Q2/vIm9JjJyc98q1m3U/1iw3J+T9rQdJQkBIyLiXfk/FLICdxR5Yi
e53Egofn7KUKe8Y1OLWBvq0WnKHrw2sHLLKOKvvS++Mvz7yQca+OHdPpjZA8+zeb
BpRkY3OCl0qdPqrsi1vCvQGaPWA9YseT5GFiy+GQ2PiKNgdaDXHgVtVBY4EnAmQG
juOk2RltY0523AhcLLrMKZ9x8nE6XX7kTYkMJs2qGyWbH5yqB+tN3uOS0gGgse2u
dZ1RRhf4ys2ql89UhzifHqOjRKDrkOswCmtG+xdoR5mj6Sug66MdbdhGWFdnPuqP
/zWYWKbP42Mj1VmtGnR2woC+BnLxghqUpTE94lGXdzkVrJgJihWRDxk32uGMWzqQ
kMqVAfz+nxRJLCdKH78eH2KvUTAHRodLhBoKKbEHifgosVLsUIs9FF+vf0YqOVkZ
uVirLxOhsQCzLGCBlLmIkzLyCd5FLa5RQk6RBAh2/hr7fmUE6P/JJjtJjHe2rp2o
q5iUXnBvh+262/FF0Owt/gH7kK1n9eQ2qW8uefQjXsBEFQTdDhME3I3H5hpq7Vd6
0ajfccvgyeU1lkLh1Ua3+qFKM/8WEz6O2XEj1oQcF7D7kfhr0kwZF9pqJ/Sz/ri7
fVstlGC8aE8hq9k2B8EMCq/huAl9yT7Q7RmIS7n8WM17adVxSkFv7TlQsq+qUd8F
7Kz/8Pweo7hpHsHwD+WIcLi1r+mEISZQ3SF3Fak9XNnb2S3SM//LmMR4k5piIEb5
vWHR7KFK88Vb7/aYEfLyLgiG/ecawVgUY2cKkZNnd2NLGtlpZLMnzuJscQWVyr5F
RuWYXx7wjWNtQW56JN3VANPDhKITLvbZu86hjh0ETI+ALNnUtF90+UYe6sRChgRL
/lpuzg95PdtzbsW8/wagMKZo0lNI8poteyE1txK37mHGrrtM+NHSaykHtytJ8rvV
hEBbm0JxUa9aSw6N4L6eDab6JxgmOxdAaIQxXuDkZx1sfT7KBhqYQ8y8jQAWn0g8
hLK5W97EewL0Xd5y10RhczfcpklrK5QNZmPYCpC/bNlt0T21KAtnKmJYB324etid
IyDodbUJMlgepQRDTV30fOz1wWnq0d5lSWX2ihosWIhi8su7gO9+ogvqTNZ+Qrll
fmhtwcp9I5PqJ62ZIX1RcjCR8cVhHG8L4k1Q7pkVo+AWuY6naFmzEDRCo7EfkGea
9WmzqQo3Hkh2JSTp9sGxJLRHiEJklexeHIsSfi+wryxiodbF8s9ZFpzjJCWyzPjy
r2YDmMeolZ0M4KVmRWITM6hBU8cmOMoY/QbOGQJPLCcYa03bvdUyd4SDIx64i8+C
3rkp2RDSi7GOBabyiPQeaT8cT2P2T7EzHHvCkmskRiG+cJEHKIgJ8aknVrOrlRXz
3VELIKkPqp4TCRdraEvLqRfMI1ymAL2WBJieuCNEeosyIz0Qq0a3J2Uv/rD70jIL
iZ0B0oYNh8IpYuEeOCgM0ge9SNapqnyiYPqPe1s/VYakwFD+f4tgrhclO0hJ2IMU
108ytJhyRXLSyw0pvCOaruMadSoJPm2uIznrGkkl+Ly60nGcP1p/uPUc6z+pTqOO
SKiw4q7LwrrbEbtw5TJmIr4ni/hC3jeinpIGHSIIBLuiwiH6vY5X4IdKhvJfUFyI
f8UwlFE4gGsdh89OjNnNmmTBoxTLYno6ngHdWS7C7lh5K4xkNTm1EArLB4YfCy3Y
9QrLIHrbUwx+npCND9Fr5TG8yTpQfKZ/1Qk1woNhezrfjLLoPZyVHmhbU9cVxF/i
7iGblYi0HVnF9TQ1zbUvJgQTKzkinWlL8Cx+6OwzClZni+UFfBeKyPwerBX5AYcd
J58aiySf6ARqsmOnNz6fSa4AZvrrJjsiEE8J1mTSIXDfDG6nTmgP1Ny5r7BUJM6Q
qA+n4bH+aMp5xXE9A6rrjYKp9oDrP3Tp02OvCi3HZDPe2uz9OIX2GIyQxk7r6Wsi
tXrcaRk5NmFGiXEXtAwhngvCv2Gmse6ZmXJH2mA6ldcc999SALt36dUDOSX3Gkki
y1fZ4c32coKUYr8ZNCnFfklrp4AFU9ufSoESHiXgQ0V5jaiwWZXL16yOr2wSnlJy
UpwhmnqBC2A0dkQm5O6KfBrt1uwk30QSfhBfuZtJJt+XET4hQ0AHMDwSPDaKRv1c
qZ8wmulhKn84RdaBI6RK7KcCOJwfKqTQV+27WdbfAnSq8ZvdZAhPnt3nfkVZrbVO
csRNBALUbDreXOMeUnJPQorgLloN6cT6xkP22bYzeBDaq98mZadosfTqm29lI8A1
E/t5MZK8SQY3mAiim3AR9CYECX2J5+3XE8URZEH4Ta2c/FU2rG3eAN7K7+T1cqZ/
UyJKvwuyOLC8+YKMVxND0avCCYDv2ID1OsxGgx9FngWoednichly5pWPinuTxnMG
HL/IkOlPulLA9p027+SFj3af/db5upqbdL2qAHU3dH3zhYdAUmNCVK6c9WYXRTEr
CLOy2jlCW5+6GrnMW8zCEdVplDR6mu/aYxo17Kiqd60LKIUAIu7zDNOyy6/Obm4c
HKBDwYaz4IC5MX88yVaY/njF6FUWqaFZy2ws30+m6x+TKuo7jfxsWfA54DpLqCjX
NzoeX7F7O0lR1DOwAUU+a7MXBCKThqQKSdEggbTicNGo/51NU19NnbyLpBg6kga2
o4tp37jhKhKPfJW3pZczutmtzzKVL8OApWkYM4aYjJzlvG7C89jfON2ljA93n03N
yLHqsokfkeKKQ79cyW7AhI6fjz8R92UjaFyVUd5c4/UJWPX0CPEKFDaNx2ojsaSH
8220aFFVUbieaXXGezbHesmx20Lld6w+iMfjhodFk3S2CJoPieZiw5xNX1WsRsm4
tsA7X9DUNsxeV0kkfB2AdAUuqoXgARbTpfK3yLkBW9GeH8/xYrCCCiB9SREGAQzI
QI34XbLrp6IE/uq3HTPLfQRTg5ChXAuNuncR5HTIlZQPK83s+exzAcPqilOaqRWY
ITHeqUiuCoLIm6H62Xarw2iER4wxN+0cIK2JVPbghAOlznrdrBYC9xNH5Wok9Gga
UIuSUl2s1Sb8QD59xbsMA9R8LX5sWg8p5vObq4wVnbtxF1VEj/fBrK8bsmyrxgiy
rl9CuZjkgagnBaFq4IaWRWR10j+bnpYfNX3kwZEnS1DBropPbQ1JJBYEhU1TTuCn
oXljWRGvirhR1SnezCNwSnwM84CifkUiwKLywL17cmH0ynlGVFEQtix4HvgvizGz
bl+rVHye/QIzzrC9pk4ULQz1JL2E1TX+Vm9knIoJE/k0RW9wOFALPkocSeZGSfp6
oEumDD71/fxZmi3d1igtszffrUgexJvUsRFNhX5elS1wF1og2skIbnBtGJZdjj5Z
TOhO071Y6PcdebrkuuRwkPcw1ATJTrXWzfbDt49Cr+JHQNeHG2JR41bLrP2uYJvk
EPv+onLy0ew4sgrILZzgQ4K58NJD3PLvGMy3I1vCBsWX5fljzROyAvg84Ps8nBu/
sIk1NXplFb85wingpRCawdNANpWwK320V5HtrO3jzQ/CqHMpwJFC7gUdn2aXkl3m
XNWxDKUgV9swHVHoN7GOA+loJZivCDzQaY69TyfyDOHIsXrcCLkIGYjMv1KDJI7L
Dvwlg4D2otc+TyP0iF+TYTE2x4poOVTUPY9C1vq2GGeqYPPWa3n2lCqOhEOGMRCy
+Yz93vAHREzZ4sT5qAwmazRNADAiWCJvOK5YULULNwxiShiUVmai5OE87iC2yckk
98lmmGwUaY7mO5pgGvcajhgWSI+GUf6JmZH9Zt828avWsMl8AidhSNPVjboKmgmO
ekFk9c7xCnYmFuZHvQ/bRaJHb0TeZPCbqgatVDIAec4+0xQb/5HYCnlZUso4lkK7
BwqWdSkDgSbvKlcvaVlAlpremDixzZV115eo92QmK3wSUllEuXEtNccli+vkDuIr
kh7g0T+OQxhwn1l91xGvMwLNGKuOu/FZZDoE9r/dNMDI1YU39hEriyTJ9WdA1O15
vr1Q2Dnsp+/d7gr+bvjlwihB9ao3GmjmhigjTipSKOfbZ+KYGJjGO0TzLXX92y7P
yy9LViw6/YiIlvQrtY5U61ZrD4LAxi537JvP6Wl7ZE8EaUm9clUWHmO7yM/vQt0Y
HASkk4DfAFsIVj31xe7zuocHVIfbajOJETgYBydTlq28QfK0YmhNXcXh77sC8ByN
hAPQxADyT9J9gF7zxDOZGMmSjYvdGkePbhJZ+GttsC721QROEb+/KIkP3x44uCIq
LjSXckQiEL73jML2bJwIOfvhFbcGMDBFCNJC6x7WqpOvamJ8YfHvUbG6F24W0Nhv
8CURiLWcSTAWQ1MusgaCSPQ77DvMtEkqWiMdHqrYFsKHz9HHbvQ90m6U9ymYPrcd
kLWK5xOnTIFU39evHxhHuYgDCDAOOs4ay3cL++Qf4NVlI2/Rvk7ipYSzsH/yd8QM
GWjDxA+Zgvjpaa+C8JXtBNNroztnzCKahyWAdBHSLpzV/D5FRVKxF8B7CEkK3bvL
RBmffAziM4zeoUj4aDkoLMIRbhlX4GX4eaNM1hY8Ymf6CvJwRBmu5lMgURBuoF+3
2+F9fVzOC9uZWfSlH3+K4Zbtlxf2igxVfMu/Dj3Si0umshhBcf5cSNjiwE2tKPWL
4oxqHcb56xv4WAI/OHuC9Ws5q9XnDjZxAWF5c9RuyfpKQVI2efgSR8YTu/8KdueS
Zf6p8n6PImtTI1bw07qnGnIYc6ainaOeMFW5+jGeYpQQMdgPL6PMlGkIlCyEt++T
peVxLm+kCcPrreJys0vQ2n9EhAc8cegflAp0dzOLXuN8JHSFVzqN2o5LpNLJkJBY
xg4kua+MDf2LN7j2gpaBL6OOm+ElCPzLEYPwv15KQLbgFtN4aFS0w2l0pcSvSUhp
bDBPjmvM6ytBm0pqYW0gi5iYLc4NlPFa+NZtIGcag+gYZpcnUKRZf0ydPnGPlooU
ufbFbjPE0fJ5ZPOeGZsHrMU+nqj44zJmKxfdcYsizC3NHqf4PXgmLcU5yE19lJK9
K31N4iHy3n6K0iNwqkPYLYRyC58TUIn/9Bam1/Igi7i1McT4ySwAAffNaw2aV4Sl
5W4vPNUeLfAO3LzTcvLi/EIUiq7SrHPbZ8ElvV4eE2X4eKL0yR09SgRUyFaMCpVi
/f5BGYfBDVXbL6nFlaIDXU+KsS+JG/ffRJ6PuFaUDd/XNfJTN5hxQA0FGra65VH4
cEpa+HBye0nt6NTranpdkhtzHTz7SK8nr1iKI1et9vCG5CLzq2Jzif3EfBxtZGns
fmBTNO8K3XvJTZBEBJSg0LQLVIccoxnqE3oBzhYnugAqGskTpVRVh9+Ae7K0Ldui
6cMEmeRapRmb+ogxuOBhlzFS5/ErTF1bJePDP95qvJfB4i7wP4gH0gp9kyVzRlq3
dagh7kmXhmFIt6K49+ZwUjBtelC/OzDp0FWbVAaxODSLByYu3ap1bfDN4gDn+wli
qC8kMLd3cPwA/n7v/kwj3bvq22VVpfUwfsPna2+MUI9ybRa6Ehl0C8fWu/QDwox1
i5WobxfHBbDeZApDP0N8VCR0wK53fk9VeSUeAiePwINr54ZIGCcchw0ZaOulNwTU
pFMzk58u2cIH5XAFpE19/WRN+6BCtmSyZq+p4U89oEM1KQXbvD345tf7yKGxdxdB
zCqAlGsgQ5eDXB5B4HAd170jSvxQ0nlpqOzABT3EuWS5/ZBQY2e3XkgxplvtSh6J
mJP+JBbn0I/7h5G4nbHmQGvi8GgAYy9bZ0AOnmf1z0upZRsdlzK4xkBrz/ZAiOL/
aaAAhojpVqMSnkLILSn57p4yWHcAAYK+y0Qr0arrBfitjVogafPZbD5PgNnySx1K
KqtNAETYoiGOUwB1hEL4OVu2AsgahOTICgOBqIgZZ6bq3IKlE1ZAYS3k6jmHjLCn
CIp5e/GAXodr8xkOdyIPNMHJJc0Tt4AHyueGfjGENtppGEidVNOPk+Sq98SiH1Ho
uxjXcOsEhqW7uqFphqxx43hkOx7H5xNahV9TjtmojLCK0Wq3HQ1qRAQO8A+RXIZl
eIcB0FXH7plXLy97Z/9JKFuW6o7SO2jla8qv+OKU2anro7bc02W2cya/sLjRsyxX
OCRX5CE1oOovhcTK8vtGHkTd+2Ug+or4gk+P/kt7wP4ACNQT4qdvu/WJ+ue1TmX5
G2u9EuxF0YMzl4y7lNT1b1gkJ2nUInTALoHT6n0kdvstCx4V530nI7SMgx1d1Hgl
D7HdwYSTAyXMeDCDYUr+jc62QKG3GxPoFzVnQwAz8XoF0KrXBrbwI6CIqsQwooVZ
9Ayz/LVLSE4s40eDwH6ybaPPJ0TEePNNnLyIVyQ+OMOQr95yFamh9hxaflpt8qVo
6RYToHiV/MfAvs7g6mqzd6DBCYNlvgfKQSfw1FhBDh2FNem0zaJjvyYdycF0ujsj
+42pMyyaEqAmlEfBWt3Po/bt4pcbSBGUIwdnKU5P+PcYabhhhR/Kc7Bk31ep8aCi
odpRNUe+/FnQN2aYm+E1tnlqfgfU+/zzq7gzbvY7E1iv8jVgekBrCUJfKfkpxSS8
xInC2dsGHHOQof7laPy+nQm3s6DdBRBAESk8KaAnpt89r9m3SwbaSWrFniOhympJ
IomLvCS3VWvOP50GJJhn5RGjR33K/TAYKpzm1U3IL5BQ3c21H1eF+ZvdBHToNKM6
NR/B6cmOJzOfauUjss5Ycq0imYIPwRByLvIdYLDlu9JRyv8s6C+HcqnM1y7S7PQv
IRHpaCsUJd38z5Q1aYhwV4fdCKsVMdbvb2DsvzheypViqLvHivG2o1mgboQudYAo
/2IHeeVB9w+DvboIGIEsH7JG1DfEq8AP0QOyUtWz2/g+H4tYZsQKR2BZVFR6A29H
5/q9bU988NP6TnsgMczIQ/c0xueW/GbXV4MXrWIgk1rodDsI/JN82CGn/BRrjgYB
QZfdiV1uYfr1+zbaTImbfvJX1aL91pd3zGLBZO1bArDbhL9ggCTYfG4fEN6Ae5ex
RIqvRAWOu/lzcodJNNvi8wu8l1U2ZHMIr2LQFV9LCyf4CmCKBlKx32ZXooUUd+u8
xGSTwsy4gqSFNZKeV9NC1Rw1xQGU/EM4ScMXu+MUmFDuKUrghkkbTqmM/BEeRYeD
cYhDFepU8YNu0uAUdF0Z0heeNOEK5OWlqpilUYDWuqDC/3H4NBu7WQLHGHj7KRol
aw/Dxqiw4J7iiW5GkfswLQuS/vuGTdkiAJVvf0NIVgVUOIjV534sIXX/2KFJ7x9U
AHU80WwIdDqEzqJlsUw/q1SGfMIBUI7ZD9aRZLhdEbMYMzKAibuinwg6QWZdC54u
5bD3/OJQ4UcudURUT69OmLpIPzdn+oZym5/EJT36Nwer6PY0ipBj+eL/5hPkEgtf
AxtnRN/QD7O2UTWjFdT6SPq6ZsfYYiEQQ3tCGM7JQ5U0W+954YFcsMCxM66XXjLC
YBbXp5qWAwTrwqmvmAenX1kTClX9LkzwI/kmwwiWbV8nnqazKjY5uxpiisGwX5F5
iFfJ8as5/GOu4JqDMAtFAqNnA6pWmJgU+wgAYERf17+aiFXvoROoPMFHNSu6UuxS
UjEHtCZ/80wpIOVwomxw17rgzz4RaQDqgCxhPUXGhzwd9cxbQ0ZjVfFA0yj12eVX
NY2q+YfzchFg3YHqd7Wj1p/7QCFjKBiDe6ftx6Zj9GzNYHb5fXYYPUnaEI23CjLp
P4Mq5F1gqvnuzd2Av22FkBAeeICWO07UWDt3MThs2d37Y8jBUgMZf2ULG2zdLsNf
fKUm/r2FSRhm81xbPZ03WnyYj7pt73OI/M/hzixV1uvcUTtBObgspYB5dfEUHMrt
LhXxepZVBhqEpWdIlU+LhPVwxCSFG1FEQDMrXX786aJHsoo7fdTeE4anSlRq7w+B
fe5tRCMgdAMznLzAaxePBEObcEJUzNmvo0z81nhLotGLAKIK20UjiI5a/koIeUet
LrPhkJRfGzgY+ydoX6PsfZqT+NSOyx7mULBFYqsVzXBx8GdNmn77Q6kG/hAsMXZk
6PudrwClz3TBdawMwkzMsThPL6QU24s5k4jHXRN4w8YkBAufUYE2dnHa0YjjtsWf
1lNn8xMsUjGneuaphnhQvmaILV/0f9/bwSt0uUywzlLx2UOy6fp+hzq7BypSccZZ
cSituC2F0K5podZanCPV6Axcixxw+7YHRP9sJ7GsBBUS7fnEL5l6KWWRIfiwRch9
KiSDMq3plDXRM91vGY31z8jxIE+KutOR/FLKDlVBPL1+Q+PGngfVGB0nQLyV19Vf
gbMzYJVC9uteiO12RiEQ//DUbo5VDLRKVDmWI3PzaAPl+WN2HtURigFvtoF6F0rB
ynCPNawjWvKvtFACsVWLtVuuzFmCLVEqg/AmmF10jA3XBhSlBD8osvSKL6CTafIf
GqOq7J4PKL0eg3b/1jaqIvnEu+9cccUti1F74+NP7QzyhbS9CjM4Ljgk6s+v/yYA
MSJN2VQ/iA3OR1oDkcy0HY5SXjWYmd/DQ9BTbLeZMHoKMFfmlGoPdxG3LMqvdzJV
mgVf4ABnZZgi+1IkTjZAmpFBJKeK78KqpjcjylJ6NWWIsvTCH7oTwEGjGNs3E1cV
dZC5c/HYMyh4KFD8zr4AouypRV0jPeuYrnsWdoTzuj685PWPtjeLqzpuzcidceZS
9lq0OgPCVr1bmOzD3xKMU8yWNyjrm/XbGA0z5K/HewDihghdWt/nlQSZQ9MaG0Iy
86zJJKV/mj1lQmwxnIB720G15INDb61OQqrr4+sn5Slz8c7yTm57a+jqqlV9GTAl
HfhlqVhS84bYPbEIG3kzCUzPShsV6mr088vM10YQao9OhwMvW2P2Eyg6rCChtGI3
CuLanhor7zHy5TVwar6mX8KNBKjnaqMd1XG1DNggxFb+TbxIAdXz7ymuVzZFyXly
9FwQ1+0NKiehwEQIH5ERCVGJnzgHX0UoxRvmSWecv8G0q4NQS5ESodiuYPm3FbaH
sZkokWTplBvmPAkv3L9GVLfOTwQUh2SycMJdpBI95qTTnkY/Gve35n6fnJf+j49R
mXUL1SnqnzEHybtyOKSBoP/U+JFn8P5cOcKhyC9Fyw8h7OkokdPEULTcmGFmfs/x
2zZDEIen1EzJgx6sYMZWWmXZ0FX2sN04TIXs8caQcvuiu9yV/umMQMF8E9lXbJGR
vLbVq20pc1cWlQiI80GD2+716ks7qozaqCOuVLiLzsnhoGC4LGDzbdjqTDYXBrKT
NOXaqjXXFaBwCslVSBQ8WZlTi7EJd7YgxTaIYEs+gIuile9etVxzQ92Vgkd+Nm2W
lj7krIlDwY3e80EuevJ9/18xf4sdS+hAS330nzJx+6/EbtepGUuj9Hp70XIM10Rj
xeb4bMzj2e2/xtSLe4XSwvB+GpDVvRgWKxlWddGvl87Oj5Lstu0YwkFq0e1bPNJE
y2J2DFdSr3MZGHv2vXAO9KCCKigamlZPSYTFYIZjrdsCMKXrktwQeQjSCMRFj4fc
ib0ibVmB3EHlV2IMSsle+PHUZazOGjFLFl5fQKw/1as9bAsnY0bPw931t+c3HYje
Dk9Zh8mvvf+rhqGC0l0QSOwQyC7lt5J+Lt8pFqdEN5iDS22JkT2g4Y0/u9yGF0Hu
LLldV+geHfSu3SwMk9ZAqH4kep6KqOfbKhJHaHnNPhfXJPOE9SQm+rHHGtROqSZi
I/BSi78p1KX1V5KqzXHZDeW7XWgmfjH6ePLZWEpPlEgDnHUSML38fAB6acqTA4vN
/nAIcv5o5f+TAksJl4ABI4zi+Kou12FvWpWCf1E8NUgb3tzaaKI5cdCvNChHn3Av
DVkzZJR7vuUhHZd2ulAutHAAO5yzt71i7/Wra4Jo0V0uuvfIfTx9HQrkYxI8+Cnq
8QaN6kxMhJ8irPvvEV4JE8Aou53wM4iuIzonREi9KmzP9jpp/Aa5XNNR+t9dymfB
/cxjI18ZCzBlzq02imWXGHiiDhCKorzEqLZdx5U6RDoGQ1JhgoXHELtiJrDb+jBs
6gBmUZ2GaoQnx/rH6Okl6K2nyvCH7FM8AvDB9ZTni3ALZlYvtlvVMS0ZHvIDCEFZ
8Xi84HjB14XzJb4V6TyklQq6YXo9HS0EPsyIqp9FZe5/6AYiREKi359d9wT3jbpp
xON3yZTCTwJdEtu5fBuqy1dovHcBqWIOK3eOeDTdzhlr/3oQW2ThKYbeSPkj6TSr
iTuaQXCB8pyvzR3ACQUNEvUPYJDS/EnPCIAcxOOk5CUuVdsTwO4I/s5lt6AbAZgl
eb9JqMwegIPSNdoW1FIwOOxggQxW9b0UzxlDY2tzCN1rZHtD6CgOCvtnZGfBvIjQ
DAPJ6SDblt9RfSMgB8lmwgw7m96J/w1h3yOjL3f+HJ6PJR3eLoNg4akyFOd1fVM6
i7AgbZQtAFCGQBvm0UOUAVaCoUPDrqeXDmN5ECyemY1kIo8MdqsqNWvSYaqUeSWn
8yCA16kQRWpV2hcjd6sIvJq+vSDtDeU4ICS8bhryHV4L2jWvAZgnjZ13bH0Vfy32
K8zJdAfjaniFo+oLqfo++psvQykKBpoT5okhZOiFi0iRwg2OIjh+fRsNYv1n9Qo9
KxeNjOcU+uCpGRHPf9hK0JCgfsU7wovs0GNgaAaC7Fv+nXFQOQXEksXzXkQmODeU
2vyaPV1MA8OSOvwgtnalYmGRwswp2YpMsd5FO3bmr2WqH+k8wk6N0URJwqMoDFYm
0niI1CEtRCkHXhRerAQIqQlprF4KE3NWbfRJ8COqKk87xdrf8uKMLYIfrb9Ae3kE
PllZ25B0Ie6CEqJTM+ZHmM0hTngFlfM+zPQx8b6zpetBZCEsKNey306puzwoX+B8
X9oHqGxIsoF6DIRdFKjr1GXlW8iJH6rQfmeXe4o7bBM5DLh2Te9YCxP//yXvW5I0
ML3da9P+Z79RljWbVqhdyeL++PIZv/KVhKZhCB7y1WVHEHnTGQtxncXktIbT7JlB
RmlGDIvBpGJXd9Hj5LruJ/HCTNzd55ICbNZIj924ANIxieaGT18rr7ch3XX/FY19
Vh61F0LEXbA4K1VO2TBh/XCgaHIursYdkcb46OyX3jvBXdvtGU892OM3t2CL/PCr
E48gVCTKOqoTr7YbIhyZ/fowZnLIJIMrgfrBK55NHC0BBztZX/kRXSyX9nu5Kki+
ev9Nc07XLPvSFkkwbFCc1BE72C87mk03j3rERyLDggLVt4AWLMWrrHYqYru75p6R
0yaZIlg5npiyCMwMufIgTGvsPKVAw+QYQJ/GDTy80IJnKUHXCSb0Y+QMqWjIt+S7
0fW7AEu1uqQpSrSf26eR1u8KFhglD95a1hMXr+EVSn6y81rY3v4XFNsBYokOX8kh
JHImDvytiI9jnSYJj9Lut8YTfhkSdh6SPWwB++fAHevO/7t3fdBjkzUq3/A/Oki6
JrOrqmu2nzrEtaE8ODiKxNK2nPDt3SppBskEowkTCHzw5u0xbn3vrzEspbZI/+zG
5CB8vK2t4rJ/i88uC75pjVEKBu41eEkCMAMwpWUpEiQFZgN/P6XxW17h/7VNIQes
kXposLBASrao9nXnJL95o3vSGP2/ZPi1B/yX8l5qwiW4Bj8gv+K765TBBN90lP8t
m0Qopeh8i7x6lYmZAfRL+kXMlK617QhGNBpkltgjRocbW+VWaKeYwBDjYRWyDTlM
7n+T+ec4QDLRxes9fimo5besmpx7mblRDOyQ8+PcrxIySg+Sxb1fGq0Lje5/xCLO
Bg1nhe8k5bvD8u1c3rgK/vwthPpiZI9xbQNMru4UfxGFsSdn6jmQYk8Qyyx6wuut
/sYPuIj/Y2qRTv4YtPqjRFj0DDkn7VMCg4jc+SnQEPJhz47n6O4EE+i+VYcHOTri
/KSNDna68YA8saZG3LGHrBy6/u5iUhfEbs/QM0roWfQ8/eqCoAZpZgNAgLigcn2V
npFPtnlckaaqF9s/oKGIegGNU/+r1ONDA7l5MPelgfE0RULuCEmXvVgGIhXA4nrO
sSzExqxBZz6klrOv/MtKx2fDSrIqSlXGpVrlWwFXvXQPeUBzi1ggstDultF74xqn
Q8K/9bPqEU4iMzuZyFqwbdW4plffdgiNLm2PAeyeMZSIuJDPtYBfWIsVceY/myor
XXn2oYVzVCNQi652RrTyUF7kkIWRb6aHWkDpO8Yv+veOJbAm0cxcHDiOJCHVUEUr
aIvoDd16tXHZmDwtLJ84UA5/rT4mpCzi+4UUu2dozRYwXfF9SCKvpvqlVvTtKAly
3BY1pu9E2GlsbHLIAUHpoVgIEMLaobwu5x7Hw388YfDxWQ1DVO+JfA0jTtml/3BE
XMVNlZqKvALOjCaDLAtlMrQ4s/xkpVmyQ4SfVX+19WqwdN0Mvrfb/x1RQAyPWRUV
wdjpHq3PUeM8GPZqWR5rCpiUWcFLud3yb1L+GaB3IRaaTkwE2Z6SlxTDD0fFCNAa
gCnCRx51wewhcrkNzUAGuR90BE6ONaBVGxyxX8ZnW48WF6bsXyLqQeOqaruDEBXW
BvGwSBKRJFkresDBGDAbvuZa6/YuxIIGo2DzxofRTUUAN4bxNJLlMVgSA52Pjd7H
3PfZoTHY2T4Fx5jyEWEl5X1innhVQUgRibduU34APU3FwjkwOaVQSkbQwMe6Zd/U
38v0HOlBZwr1x5Q6NUy0mrvjIWbJO7/8QFIb7TP8PF4SOmA2a987rv44SIhidq18
/f1fhZffILa5GceCz6C0BjCXsJGXyIyqRr4Sj/Ah8G8okqFytCS9HW2dAKbVwm+e
3PhEwNt0GQQGemNESvcNfXV4yNnBTZAhTOZ46mW/NBm49tQ9cwdvzrrEl7xkKKqX
cWocwlroZdaHtlu+fYv60UYSrkTE7B7/s03zmrsFQ5UDH0HZR5XCHDCzIzQLmKh5
aJIXDSmAaZmH1uYWg1JJHLXRlxatqFvCyk2/FGnOV4yZZAoYGH0zZxVg9evCrZN2
xGDl0DtuwUinJCUkIJSz6Vbf0hYA+uTktv2A7lj7eg1YgwtIV8B7C5WUJHdYh9Ub
Zc9AndhUv26ekrQkim9RSAtoktxdkpJ49UiYS2FAPhlvVg1zKixZ1VSMLsSRKTWN
zIjb0zcDky+P3we3d6FiUarhEwr8ZIXaAc+KIyp4WSha3sbS9wLPB31/b9fDuDc0
BIGt8O24RP5FCxwiM/v1MsIiVXfcVArd7pYV3WdtL9uPfbLiImm4UKyS4/RI99TS
J80dHt46nFzukDPk0dap7gOL4ZRh99/2BH03KfTTI1N7go0MucplaVqJXoFqRY5/
yBhdWktOUPffeY4MgSln6IbM5rzIdpDRVcZZi+6cWkM+acC1qPeHWnLcBRjQv/yP
PWIZu2j7WldqmeJWA00/U0pk6PP5ydlXEZ+pm8BZmK0WhHjlkncWtzCZNE/mi8Jq
rCDjejOam+btMxryGPzL8bhojY7I18WKPihtNHYk7wm3Y059LPjtFH4hCohw/616
dwAyryrdU+8DU5s0dzoNuMe3B1MXGIEiR+IInENohOzyyMnfaYbo+GTFgI8Xy1T2
e8iGO6KxWwWX1ZbOWis3peQ4WJsvcOKOjRpXWAPtg4LaMolIMFaqW6WhTCdxz3qX
4InmgFziPgGf7Ke8SMsP7rvXvbB1J0caAhEzULPyfWJLxsh4RmSGSUz9ZTJ3waa5
IiOPmP9in5/4rg1DqOhqSwPnmqxjiV00TkYtamHscvHUdfYBTO0zFGkcxUarcMac
3Og660YFszTtVugOICkGLUkhHKJo9fki3urYzG0rH9Twj0YEj/fALsSiiStEGXWc
kXCZu85VBaBtfKCIVljLLmpobK5ngXvjfFqor9ODZ5aQA+MbTF3L+/V7PyIFnScu
KI+pfOjh/uIpfeztxzBG0TmqibOMr25sWPZ/DZIxPgukV7Qsvy3IjhFtokAcE0IR
FH4m8GE1j0OEpAG7wemmcgJ3Q7sS6tBDQjbJ9CcE9v4q8xukvUHdW51chWGLJSAQ
UmQX981Pnh1jMQfEIWnd36iYIa2qObmCmEZ433/yhiNpQCt7lnHb9i6J3uxArR+a
DisgerLxmOCfVGbh2CrBkv9M0yt2ssJF4Z4Nj0bD8Z7XsQrh+uK6ctdzfXwBgZxw
aVUGtHgDcd6HVjVFDxnAkB/tOq2n1VhDAFGn+4E90FehpIP/KEM3Xm9/M9QCT6vt
+CJb8OsfMYiktUsSGqkku/Sq9Uu6rhkDdpxjN68KRWrIc6HmXjjsvorHcoVRrcZz
Vsg0oB/1tcAuelpltz0VHocVK3pM8eAx6ibmvjylFoGOo6ZYZn3prnMVeEuzJU8S
CjfblgTgsQcONkwUTGuEyjUgQLLGegOo9+ah7IYG+ItuyZtsJP6PWnh+Ja/02TiD
K5VdS8eRGAguQUyfG0Hyqznj6HYvAr3VUxv8oxn8NIcZI8Aq2zgPxvSnmMztm570
H6Cb/x1mdv+8f2VJVi75oyU+jQux6BOmDjT8DRzn2dwF4E8WZWYjekj0x0opblir
JUj2JzIOr5Ro/sE4QyzUwW2a5G7qxWlJe8b8eq4uNp255WmmceQl3bhfvccO/NLB
bXm3MCtWXqapmvtEXMi9AX1i91AegwK2KKHY63lwaMcDOabc3VYd9tcNXu2OLTkQ
1KQXLiZc4QfBspO4DoSGexSNzYmUulcKbhi9vHvkLQ5HGse/WBIymYiAEZ8zMgL3
cl111Bf4L6Jnrdf4tGH5Y+RIPsTrnhCGTl1f6soIR0p9KD3BNJfyLd1X8C+eW0vs
jvaduSH1TnQhRgF2m0+zYRjrVIzATCaZ2KpHBPzMaKOfT49gT58KZMhAxRs5g2IX
tHJn6QFZKYRj+UFsSmWz0ygXLcpODJ+4ikiYD4y4p8uEY0NMSyavBFa/3/kZqwsW
Om5wz4qMER2M2s34xdeEk9HpR00/CXB1tqS7QGHu2v8NmDIJinhegvn6EnN0Hn83
zIxF+uKvgfdv/MxmhggSV+C1L+eijRPRcTSk/qUGMIw6SJHcGeQWpcgeQ3T5Kzqk
JTg7Bxh68ZVjhKMqr4+THzFnuoXEOobKxtIRlIARsKyjxaiqremEez442XUx2D9/
+3avNSbHoOMEwOxU6iHpxqfnhWMcXzIzNceF9uB2BoibBve5sxeUCM3fItTa6n1q
X0WjDX9OQR1H+z1PA88Y14yIjV8X0VzZg1v9xtytMPrLBWQVq+yuuMBdFvhNFlmJ
MI8r7zFYqvPTjPVwP7FGz2IhPRj6W1Xo7G0xkzea0UoMPefApOzKvwp8zuhifP89
3iOz5mGPqN0h6E/FVY835cCgxpX4IJkeXzZjYhXowzVj9er/6hr+bEGq7eLpF4HX
HtZAd+mIoby+Y8JuzAOP6kg67BJcnsvGoLDye4qEkZFXGc8q2p4TEpC/qlNXkoMo
VL0GJbNMTEqPRvUzZxxBbOne8oNKFbGCTvOb4kAi947JofXQXPAlbNtPIl1IlBMb
zJy1In9pula/HVx3ESZXyo78deDjgPqpcQEc/1FJjF/aLyjJS9KEDpXajma2MDj2
399nzrMHcvuV51K25veN/3GBsz1mLbLY06Wpd23FK2IH9PsyrlKrpG3R/Ll4raQe
3iSVhxYFet8pzWPjAoQtj9FQobW1OccbfcTW2DqKGW1PIUN9eXz6N8VGiTWmRK1B
oyaf2wPQRz4Vxk5KYgIFjivvewmBrnTbHeJAoR9zVuLTDReGBKqsCoZ8Hp3v3hoc
BcKeTi5nhFa20s/9glkTZ8XdOAIjxRPJY60gG68kcPV2gmxOBydEC9dGKh+P0XP1
4PIy70ZbZtcxWRvckNzYFkfm9Gn+IPd/JoyrqLTVsKoJ/CnDHBIEJHu+Ps2pK7rx
lCdGRgwyL3XhsRvUstI5FHae2BgmXFeYHLVYJCKO3/SsIUc2gRlhGnFSFg0jh/kr
JBTvAwbjxdvlSQH5kUq7yYROgqkOzBoCEwyQnVwAf8vMh4eybS1dPkWqUN84Y+zy
tFXpHskCK5iBJNlspPjF62WvehwWROEZdPJsye4NxjnEexdyXCdwCpzvALO7wAG0
VpFLk2E+U+cFtFOVHWHb4FlzRG9kd55V/7cPn9TfE4Cph+omGG2iLmJD7BUV7oLM
ijXDA6IgHbQk7y/8qz6Pq1z144rGEMcP3J8+FR/0fTBkWNDSh7b+2FV8EtvH9X+j
lQReJHRV17JwQoNrkCZT8SV2Yf3sZkzRlCAOSjPobuY209nRV0uUFbwxUSRA4HO2
xC15ube+R7hA75dFISUz1Fnb0Rd2DdsnDGtD9wGLAov/JOVTnAESdjnICc6yUwzP
B5M1n0pqKUtOvx27M/Wbcw1mezVNU3euvP3fqjyR3zuMIHWrEK+yHzpKbNgiDl2/
V+HlIqmmf0b0Ibla3JQHPYCszv8uuNQIDcVxK7z2Pbme1oSNQ2dJ3FocVzb+6vX1
4qurcLrEN+ilwlVMXBBOFZhZwuT9L6KXcDqnliNRtlZiwNcVefXGfR0LODe82IO3
QN8GCLa04C38+ocY0+COqPCB/kaNfzJptfeDMyTKeLKNyMSzdG3ze7I+M52lcivg
FoyrJLhUAueRbrAu+/xEEgY6sxDHDoSOSskyC+KaglGedlXWUPxESeRDTQwk56BZ
TMyw3v4ZhbkFN+IxRM+bRWA7H9FOMY1+UganfpJ9nIDPysdechXe4pHsPPm/Pevj
/FyYs35Iqa8nkbzNb66Aj59UVAePD2NoitNRu+9Qospl7wR/7V82zxnj4HashfIH
O5E9wG4l0DdzsNEiVP5QRR4bGyNLbmA69keJFxnLS/4E1bU+0qWVoGixFQ4hBT8a
d6zLvKfWqFQeJUF4WjphYEk3RN3h6TGntEb6G+BzpNGJ9eSHvbfgsAOO0q++4bEg
UULy2c0d5mjEkB0naZFVQLyGFempBr7+rTm9oR6A6Q1Sb5b6nIhUXWPj4PKk/rdl
07ShossI6K5alSaiY+c1oOTjC6BfuLiS6Z5fxY4yPHdjSqLbHN793PQhqgfq5u38
Qzvagqj6Egt4AozpWkJdDtd84HGcGsBXPNrSTqOgxPe5RpS9mC3t1WhGb1ck/jXH
DJ+HgqTtNh5oeeKrYP5DmeqsiIIGUk8rOtZtRStSPnhStBzedG63cLTVJvRNcdlV
Rx0xb9SeyCPUmifwf+4w1fwR0whHU1bdkJ1hRIFixRr3ogU2S5ApmCTL2BknWQMO
HIL/KDFLQVWvO8DkdxCGnvq5Idu8gpZpbZ1i4fa2JZfn5DE1Ive6uVZn47Ss6osM
+I+2zXI/1z98c7okpd3Tu+o5mGzxlHbROTHEjYApmHkonLhCb7cxRlVP5y6nfrzE
lbewQSasi5B5rxBsmYURcwmTfTjrJE170SkQCsRDZ4W5jtYqYZVNXmFP27nmTweY
Im3JMhvsv0Rp0VN/DcUCqggFZArz/pnahkMpEShDTg1upcRiImZJVtpTgf6oN5Jh
/k0fm0cZU6PAPyE9gyfheof2zVswJpWZNiowRxkSgjNlB9Ow3cqeYCL966Dk0UEF
qJG7PQviHaX49xAANPaqj8AL69fBJe/vi4fPolVEQK9YYxE+ZNVgHPAC0rT5uvd5
ej/2J8on4xoTw3R1+rUm9vydr58bRglTg38LRJ0wvFGcJTFY2FPOGbiaawI0SwZd
yFMSMFL6sHoJkA2wazOZrKeu67utZKxJxssc4aa+PdYd1R2g9dJOAytU7G8d/K71
q3cj+mk/v6wgVD5sJ3NOSjvdiE7yW143L9OZ6C/DPrueyc9MFRlai1tAreZhV+v0
jXTfG11EOcHBLQCoayA0KlrKwPn/dT4sq2oofJEwBFWTg5wS1xEyZe5GviTDQbvy
67F0Xh02k8aG2n20Y+gDrRR3wtzkMtWSN+e1wGeKRLD2IIDZRuiVMVNJKp8ZVIlk
gNppguI1an2WFZ5+bMb9TcnaVYd8seTtuf+XNTp5JUOUcrPwuLaabR3Jwrzc9ThZ
rm8aNwo3xkiQHGJNemjk397iEB8rs65baEDm1csiXt7nta/IwIqWJBYlbI5oJ0Cf
z48iVSlu4GXDmwKq7ePuD3MGmXUqSNNsLvmgmXA/khgIxNoXipBzlBQoCpMk5Vko
oDPl7b/wbvX+ogfvcr3pHCzProUFzdQlTUvfXpZ2XCySpd/LsEX2KCEFsrT7C6k1
37Tm29OnzWHJKca0NavseK/qpCWjYGGzrFy2f2l6p5kOe7jVzjKqK+H76IH3Jxxi
5AsS/+1CZKIlk5zPLvaq+5hWZRYk2WO4luuo/XjCih1r8BGXiB+Bw9xFul275RKo
CfinmODFOXDX2hc1NpH0kBJ0hDKxL3vgRmbp2tpfPRDs4LOb05VK7Xkoh+gGCK82
Lkk+yhDYSif4JgZbg76ZaabNl6g7WbCnkqUcWCjeVTV2XWDlFAVel3BZjXZbkxp9
SvfHg26PG/FkXPIG5zFbCehBHcC40KWyOiAyckNbBBws+eM5l9/SlTXQgO/d4j7X
Uu4wOYYoRTAIYLg//sOH1CuYV053zRA4eyE6a4coAwxqzbzsZGqG7pdzE8pXm18P
MNKqsWOaLyAjLT1o9XhIUtaD7jl4al0MQWZn4DMPSBVUUF1F60bTHN7l7UBRtZow
WUI9RZlqqzXvDaTpUbke4K+J4Hymb7kq4jJ8J0zv1/MX1cosjx2YaBc4hHzlT8MG
E4Ywe6ZhX19aaDRzFNy9ryPSph9j4C2dEepHv3NCpdeUIr8ME345d9FIYitovVmM
R9prSEzpzgw5sZCK4gTSrQQqi+CXKwXcdDRPbDmDamkNEn/U4oZTRX6hvH+RCtwk
1jwMNnmZl2twtEtNd49Qf5HQ3KX+wYnMXblvOIdRgzR6Ql8ZIBh8++tJBoe5oXoK
gN72+uWgcy9mSV/A5luWlnn6rPgDkpNE1eNOfHRzq0at+npROSEnaiNYoeT3JTYQ
Njt3saLq90c9R7/ti9ivpbULBAvn4DJcY+x4fpR8PQa41fuoNUJUxmqpQJCcQYPX
PR7/qssF1tvqRZoX46UxDMmBsKbq9OwTJoofgiPTB+xl1gWknmVPR7GlJVY43qNC
4QyaeDYxeNl2BPkhH+Wa/8UDv+/PLMRzXkz127QKzLLqBewFZriq7tuHOiXX7roR
qkCr24w5RKVMGmWcWUU/Jy3n0QUoTVflkXGpv24MX57QURG8b4cifpSeeYP2zyoh
07DVlda8HgsyRau5yFSLD5gvDAnrYBBZ+36vLyOSee78fEAVrsrUvGtjLeK5x2CE
qZAXyCvHZ1lbKRj9nsHpNJdkCOIBmJeIluN5KaAq/LEnRrSyKF5Ba0F/qTGfGyKa
Qz8cTB8crhPLkDaXmJq3pk7Cf6YnkOG9dACmZoqPRr8eD5b5+TATHqgSipqKSVDa
CdEzSRKebCK2hk+9uClsiGZYwPe3JRm375ku3YzJcBvY/UNdmE5NnSanBgsqLVPm
3FCxd+CVvi89OchLLA/8IqKg8M/WMl5tlvM7VxzFJo74xWo5ap2gEJW4jsjYW26+
VJW7wffNNhzFWvqwysyKQIOcZxmGtQ8ISzE9Z1xh4R2TWDCO4AhthXkXAa3KFN0h
w8uCd+srYvTFR1Fe/J17338fsZ89ZMQ2G6+E2WSIMHN55T9KMKce6vsg+1Qq5S0R
fA098Vq3f9tIOCFd/mJAyRWlAP5l18CYjf/0bt0VtA3BfRZJIauyP9ZmxpUpzHCf
yPvBqd0seHMoJCC53OCe7XsfJDBjRXkDiTzy//lZEuWINlmgN06iK3mTeSYtDKW2
2o7aEH1TvKXVcnyboY20MMlUFBYGJjTShSbCTLYrg51q0LxtdcCAsC5XlKLRDxPX
fhmiHA1n3jssOuWbffLcvTkg3TsEDyBdk4fmrlBlM2RDFWkz5+5Xygtfbg91zo6M
del2LUvjf0kLfG6C9+sHcxL8KeTSjTwvK6K0JDhqPdsI/HcV1zMwWDtdLqU8o9gZ
B0bA6dp98h1rEoyXWE+tHc7onh3zfZAVh8kOnfQKugV2KdDVYD8QSY2bwLOjrfak
ioGVyf3yIAG8+6kaIRsAFlsPZQa5Qo4gFMJSHq5heciiXqWGqnmJKC30gcJaIuf0
vzgwJEaMDHPCxWhauvaYCaCFea7TiFC6bT/zGRXJNK6TIWg8qvZbH5eLgDCKWn7E
afI1Q6jYN0FU8oEfWl0cMTpPzAInWkv68Ljkc3uvbIpLvYnPwg+xJ+XB9JPFLwk1
JxVUR4WsV1/FpSH2EOU/psbnj2CTWnB4xM4/ChS6C+tEeJi7xK5qzCnVbER4nhKu
hFO6GTOdx+0St6UQsFzoVFZeD5v9A18BTDR/XPWhG+zlQD8nndxIjrxGashz/u3J
FEXfXEvqpfW3cCGm0UG4lbJdzNxObnpe2WoVsw8pbEYO2jR58UyctidED1NLazT6
l1CayDuMAY1J6TIplS2KYIW5oZnJVAohw5UucGskE/IIPSjSwKqT/jviF6xGmGx8
JsAEYPjMD7dkChtsNnl+vXEubJ1O3oNELqc37beuQwh1CiuBpWPztw9MIdGVngxI
zz3Wv9aVfupJ5+Yf36FAdNB8wIVol8NBawUBkmQe7mUA8OaJj+qyU5OSdLnCJGga
NTnYrqN2AmvztYGRw1Kf/CWbUdLqgS6z7k35si48KOUHGqFAj0C1bBxMQd9rWwmZ
0augDeU4+DlDZNX2vthvCHs8E4QvVjdkyj2aHDptiDE722tedRI7j5g/ci/rgQLW
A6Dlm5pQsWPlKlS6VuuiD75bLIloXpkBWdISqqvgdVCN2cKL0UTHxcH5+hJygCKZ
JHiOEM3PZX8nIWJE5a7cbws10zaSceyfmORKgiq7vGbvNolzmB/ZhiotmBXcZceA
ZJQTqiTJa301PpQjY8AFDZSCc0pYSF6eVUgS2BKWvGwYIW1d8gqxVsuDfCm89/8Q
SB1AKz5lTWYaZrv7GAV8//9ZGMMs77aPC2yMUNHUd38c6fg/k0ER4iTUb5VkJrUa
20Xt9vAQutedHfXdImhYEojpIRI5MELBC/7nOsdL0NU6qtjJ/aOYDBMmIuR181y1
yduvMsFf4peQRJ96vLdUeDsYoIJyeJXV1uWSr/YLUquAEMMi1BtRyfxu9ihObYn7
ywIxlfLhDBPQPLXNJGxJ2+q6woAkeaJckqc04hci6NZp8B5A1p/RL/rBaP7afH12
FtGrgOdUuCPn35m9uyzCshe2PpAOsQzgw5r6Kpo9Q3v2XHNv2wf7PO6qdwrLkpxn
Fx3URIAjRv0gxgQSb97rGzqDe5Ys74KFXcbsWFYRjPcMvlnT6rr1/tER1Xx37/6h
K0Ak4WoMB/rzlM5IdtbGZloj5E1naYRh/ZLEFFy6blsTw27UCNvkv4Bpq7zj7irW
YP4vVZDGuEW77/9i8B4lpA7hzBjVbpb3ok2Mlk4XgqlyYukEvLeWsQnChXkIFjFR
YeQMBVPBo0xJfLvDQ6kCR6wD4MFsSNahplDArbWbRdDpZSkJMzGa2b64XxidXmCF
KKbIb3DpIhNZtiDJsu81ev8/r9ipreWtMhx0zi2TDRol5re7Rv8jHklOYLF7f1cz
WKT/yEhZcHyrlPCTLNeE17f1yMdU4wRgo3V66n3LE4n4JbY1ISxkalBTFO2ehNWW
nFxq8/gV9Hm9jmVLAp9ffAl7o6AQv5WXmk8ksJefoYjAS5zkMxjCO+gwRJcpnRpN
0alFLsFGvC8rHoaO37xHLqprDnMTzLPLZUmNHLz1Uz0os+6+Gv7FXqE1Kb+5ZmXD
vpiPzEwaORC6SwARFMfpFR1mugriO/CfyfetlFj9LNyuR20Fed9PQJauI6jjL76Q
b0ZYPlXzSa6ZMuq/CWi1Jh6eWIxkoRw5jA/X9byZpRlTXqfz4d4e9yCYuZP2vHGm
z8qQHQYXkI3OjMs2feyJVblNmrIVUi/JWFcet3YpVy3UE9Fv9LPrLDRahyma1UGq
rmJDT4EQsMp6s/IOxtIVXeg9o/4RvYbmdfQsPoQ1gG/8dwIds3SZXpTU7ne3xr9h
RmxiLNJKmJ4wgH0+BfbL2DkQ1o/qHU0baMbhE7pEFe8HbaG0UkavEt4ACOYVW/nz
lOvI4IHWwU6vGiAj8XyFpcPBHqug/hPKJNycFFI0p4rASIvsj7GVlIPqD15nuXKQ
xSxHbm6ImfFZ9rjvrck10gtSPhZiZR/WpjN61CcyD1aqvy8x7ySmwHaREsYNo5X6
1bGKY1FWbCQteg5vJUXM/7f9BXUmCq7yHBEDxLGkMiVP+SFvJm16TZKV1dlEoiAn
fm3qgDYEX4NevWShpsU/GjRAwfKFeC+OhT4DKKj5uOAr8CY/A/mmUI4stdo2kfK3
Qcj7IumNHSIaoi/80s7yXx2yPNtXrtQBxGuKJ4PMx6QlsC8bIdg91qumHJxtEhLY
dp68a2ibXPULntLi100NG3AaIL4Z5U+59jZm9G4Q30ZaLE/eNt1tpn0wo2+ZBbMq
XJkbFnb92KM4x6RyxZthiN3P4oq2MOezMPZedGmtqfVX0OrqO2Z+YfTbIP5XBOSL
R9224KkvTc8Co7gqtGqgXsOGQJBv26aonMatGax7+VTYke1kX1+hMvf8EzLXB1Lf
bF2Sm8q29G9PRK80iS3pgqSLQTfwVGwQtq7kedWUqXICFIFGJkG3EBb23xtBozRg
YUuzC5xNlWkE5aioLUk79VO5RSw08enf3Zs3SuTK63FByZG6hVGBZhNL1+Bhjce2
evb/ilcKQHSdkFxPBlefdfDwrdR6ky3U1FcuF5ioyK8hTw0+isTxv/bcQ7eGvjs4
hf90zMQQHUfgP9trznO10LawPbPhojuzLfxt2TsWMWfjqqWO9mI2U5FB/rE914cZ
Ttj6hsZX+hrrxNKuw2lGvnwL3qU5DBhilBbtCI0meQDfVHf3Wc80F7kNsQhHF3Uv
PzQv5KiZJxsxkwwJcWLz26jiVkywENsT2mHeVoXXbWaFwEbwGRRqEyWzyU/r9LjH
NDG1muuqm8u9dmVF7KABHhGSFCY6W1ai+BWQs3jYb1OFrbpx97tsrmY0/lnCIUDL
IVsZ+04/L+eL3dCLW/kxIMQD7B4/L0RINZc/yW9Iv7bv+r0NPJV9lRlErhzMYgCc
HyfptQhsEmynbTsem0fOPxSpcz8oNf1xqcbDgLrkc2GqGd749/V0BAT1eOstMY6M
2T//nu+D2ugWDsz/DbcU9QJH5qU6BrzX2+8fCCj0XbznNxwQw81ZUm1QGNYmv/hL
KHumOxaIMbgPp4sLqJvmg/2rlHITgBzsNQREbNbLFajyr1LV+x68X+nZI2Z1jrwx
OcRjWWqotf6hcHWmSFcnbU6G9dHGHLzgAI5c9L7BRaOcmqeBYya6BZ5qahGtrmUk
lWSzFXPdd6vm34LvtHp9HszQYE1VJ4urVnqgVMXhsSWPG6hqPsOD3ArhcCDrhXIB
rbFMzN+Hd79KaO5C9wvd7+9ppeHZ4CabxoIrezb5xy9k8Zo17ccZnmfqTa19Dcgu
39NgrFH5GAljEfbF5/jspMocQhz7oJeFM4ul3GQqceY9YYJJc2oH3ST6fWy7CJp/
N6znsd8/y/6CVqOqkok763p1F10Slqjl1Gt98marCm/Tp423IEb0Q8Tx8w4kHQkk
9PlvvOinD+8KNqDQHJXwG2CxHAdRTKePef6RYrEOhjCDVjDvZFKAViMtI0fb6brv
RhJ/8GOQcWjlOxSD2HgZlfz4mr5VpuEoHVcCBTAg9KYDBGXLgs0yIyCvc425eXFB
unSOjAw965QPIoJF2aJ0dLsR7/IX/2SJwp1WYOkJV3Hlunhax4L+POL0NVi2MTYV
n9zVFVwZWBk31pWJ8LXszrYNLddtonJHZGvBaPFMEyH/F61f9rLR6cV/h17YW/as
iKzaDPBhCzBGLQDYVqTEfU0z+4JixgBcxy0ICLyxOFwyIqPmKTogesikCZynSZcj
xkQNRus35TaQv3OzVBgtNty6vyV7O4oOniNVjRWD7F6PN1KezSV5GU+cX/VMQmlv
NXcWIamDmk//j3ME/e88SkVRyA9cfhqHCJUFHPzkBstO8vEQ1R9A8dlbNwGI7p2L
Q8H2sMakglIjs7a6OiwA1iBAR5WStCpBoJ9JoTMo6Se7pa/gflpQ+U018FHHDen6
n+tDIi4r3PvhgV1mUqthIvUwoQ85ZtxoOUtJWcGWq74RXhmlBaH7uHNxBQg3UaHq
psW3VBoHP4N24Ye78JeKNt7u+o/zawbLHPCRjOFptsQ05pM3Gx9smMKBI/bXBDdi
7ACAo+xnHRwUZ+kmiPQIwyZOI+w9S5cIBQMp+OjP/HWNbBls3ayXthYYew8wyQHw
XLBMGJRsk7KPF8tEC4+0YBZq1BOWPlx61ki8/VInso5W4/JNUeHIeSq5edKEm+3G
X6G5Yka8MwVpTxcLEWQXTD0XGjMNOCKCSmty71dWWGX/jE3mvNbOFZDrpIXC6/Ya
nvtbrF3QpItG0v8cTn19hBYjBYsSoPa7AYz+ahW5Ak0Y7Y8pCkOEKBp9tRASk9SR
VTAgBHQnPr1JBhaPFVYeWKO1tJCViNvDPCM0leqlBOCJuLoTDPTvwyrYFXNVcmrw
KqN/f4ddROe86r1opmhKH7dX4VKjkSKtJA0ua3cWPNQ/cFI1/Wyx+wrZ6sKtQQ97
BbdtOgwFXPkLAMd/t43Uc5RQTTue4VNi017xuHnctOqeM8O+Khnm9TUBjgVz8Azs
Gc423y50GFIBNlhoYz0Fezed4x27AZThsDfDtBF1i1CRoVXtByybono05wHu98X7
4g6r5BinOpxEVi9TEfS9khEbM44Dwui5oe5veNzgVUldTfnBu2CwQMwgIFGsmGu1
Wcbn4HDAA2z1JnWgrG3+WZzYDimlIAvYtZh+Fwunejaj6jHwmtYcQPtNT0PJnDer
ZI7jDGc4DEIMm94uz1tY1WIRPVFaQ5BuN8kPINxfaBN2WDP7PjHhqqcbOMbOW4vi
Kr71EflDqxUTF9kdhRiDu4gSsaCONJYmJaLPa5e+lAb048nZw6XLcBiE0SDBEmgd
NiucCITizc7CTPTa086esJahNTYDhdxr6HrBpvLWzks2yFsQsaS8AR8IUacPMR+f
6ogGsiFlzsNvu4ECJtuTC9DchkykqnqJqOQhBZ5XAO3MG7VWQmhHPrSGqMZPN8cc
OoXSIzPVNJNEQ/2NBWZGR760W0x83vFcPtJZQGfDxDfbBBjdWnu92ZlowrKMxdBl
mtn+aUf3vrmYYNAICLhQlB75EWsKBegQ5s0ioM387hl8bKOnhtiw0EIiNNr+9r8r
ky7taZdeUVqVS/0vMwfXk0k127gsXEI1+7mMRX3QPHtDUxZcUS+yTxTWT1no113a
mwcl/aMyvVDtFhkALG4mxjyN/Z1448m2eobHRSOGRqSpqOiK1+x9VwtlK17iP3vN
IsOnjj2VY1ajGLngXwZMrlYrOiJdPxCcC21aQXf9yKiXqqCjooJfi3JaoBgqJBEr
BxcCZ3U/0rkYzmXNFjGFCgZD38+4psrz5SHzg7Ox1Pv31yJt5jN5b6xZb1Q/oFAf
a9EwgPputYoPkUOt9OKgyT2s4ouHqNC/vi6WAI8xwy3zK1EGqd9Rczua2iB8L5d2
8gl8AVP9QGwRm8evst8Vo8s0avXbAGQN8XnDMUwQTMkqfLyqJvlo2zc0NlQZao4s
6LfkhJMfHM0axAsEqRNuSYhyAdUCKcOpBxMqUYbqaGE61lAgSpwC+K9P3J8++PDa
iGvTX9sy43EXElabf7Ioum51309fyD3V3gTAGa92ptBetSPU7rnQhaVt+i4IKdgp
asByvQHQX1RxPAt5laajh0TsLOeqNUfy4awnaypM5r1ig5/AE97Lr4CLLssXq+ck
jU0K+EkJJtD6peXcPRPKIqKgfl1t5xQGdp66S5totLjPm0VDtguEUUDAsIneeCgh
cJMecvCLCJj4bgCCbJMI1RKFPM+yELqkaTVzSnmbvlc8aIzFwqfexnLGuxXPu9HY
29tLmfeCxXvEit4J9+1F2z9Ke0nrNQAdqXHYs35fmh8ZHpaf3fmw2icdR8F/Q5UF
XK/1zZCMYpJKAHaeiyKyFnq+2z/RaXBtc9Oc5BiVFWUmX9lH0A9wUHtV7Mq0BMMb
kzgwDAHwn0tjawHekSLNFxUrDXgJwfIcIafcJOwUABjqucpxrvdFLjWUdsrrn5bx
aVrb/7UUrbLKsXyFVQrIOxLo6EKIepSoYMTnWN30m5YmNUyCIJVDEGJCE80XMH+Q
yuH/S/TPd1E2VYh/Vpgafo0wUTWSmXyZUFBLeTFPDVeW9+d4/icXl7FU1sE4N+WQ
W/9l2hkMOvBAJdfE521uVQOwpNEm4prcNeKp80s5EQaV7Mm1ZjnXTs388jiSc70/
FeryJi+GROLbzXH7bq66lYoRPWE8tAwcV8vDqPQ+o6Q64lJjK44n32ehrldRgIVJ
x6cN1goeeoY89myNcUpulbbeDW15FzkECB3L5AENdY9Ro0M/dWHVEVgTc0pYjIJx
Y7f3QQA3IFDLj5KyJbjXSdkJ21rkRRRPluqhturksNTqyPiFUG6LPY1R1uD3yGB9
PvX0B3SDkrzAlavw/BsBdwTb9YoNPEKqIoMfeLz1J/0XydcLen8UcVy88XuBWuAQ
St0GLH2yUuT/VnC4y8UDgtuuFxm9e0BkpNK2u3Q7YPFSbgzuBH2CJzxfCzs8eKjv
7bcdFiY6AY8eXuQN1bdoeAQj9nI9sTiQSeyxA4yPPPfq0A1W3ZCs35hYFM4l98+a
qAGyr0sV6l5YCOMErius2Zfy53Cx/vKQ8KgaXfd2xyVIcIbhvG6Azzg9b63+0drw
TBM1uC5fHflOu3TUUNP+dmbd+Eo+I5sU6Ff8m4KVw97nrX1fOQhkyzwTpQEAlZPz
BiS/ycZ/8DD8E0T92PwgeuSqCRrB+EpLKc7dcqjEgJopeDAe/hhWJU6ROFZR5BaF
1SgPZCGnjaGNqBAPUlUTKRpkhlHsXArlW+Q49rN3S+IleipGh4ZKdPNIJ6fvrjQM
+0xOaZypzvDzJP2Et/wXBl5Zy36616FWN9ylzF9Wj7aaH95Se6cZXU2Dy6yD4+WC
FEfu20kNHGxh6FMWgYvr3u5vHWE5GS5TI00DmNjmj581f03R1ads9Z7mDi0Z19NK
VODD0ljAQ0POkLk77AVDFQ9N3SnCVL/KlficeF+hBCc19/2hfl6/q/vyhIzp/3r8
7ofNTr1tVd8cyAPZtcFHWvjlqKiCeo4qmdpk6aAGK08rDt3hUYR7Z2TlqHkA2lam
i0fryOR1uNg80POlWviNS++Az+eK6DKtUoYGV3gIqwV6gl9NM9hKF6/7HbKuQuou
JnJIUhcPFIRnd0sHzyqHHKR8GHolj0UpObo9C+5fhzXzZcVNa1/olJ3Qm7M4RsAf
VaRw3/kpNcN7mtHuTzT4cbacNR1DTo2XxZBWi0DJRotjCqNZRxJbmqzFeaWWxyhk
QfEmHn29Btr7IFxM5KOEhrskONSus6ZidhZkTigOhiwZLx4pIiSsCOkfA4B5vHWL
pVwc6mG1cQ/HOLBeHjMwTrtbyBAwnGXauDYdSipzJdq6Zi4C5sfT9uxGiF6j5bAD
BxlkXVb/SEbFbNmI15hZ1yvn/ByfzIDkFz2HJ8/cy60GG4V+puYCRpZkkJ50v7uJ
yrvZoF+TEmJlV/fFnNv7jnvhPwYPoVDw/bnDoUv5H2QGgDzxQ/cQ/3MV0DnLtPJq
vr6Ki7033CEOzvH1lA0+ZaIuq/ErlipF5OfmaGQWLfFF1p3N5IUYNkpuJbGVnj9x
qtgbWVqm2jmuL6/HOjZyf4Fwxq61gETrb5rvgbqL+0JY2fAcW5BCUl8ub5ZcGKXs
UsXC5/lVj1f8gJikJMeUVZqWqzW/pkvpTB7fE6S+1ANKsy33CLLC5y6jXjqXd47k
1j4V9JPw9s3JMmQNiMEJ8Z/n1Gdqa6sOp5WlznVtocnA8WuMZfJzjB7jkz1aM314
6mfB+OJySWbTR6CL6I0oS+cLUutBZh5gFVg8BVoMGI3a3fRuyJ/o7hKPTnedGHeo
9b4Nk1l85PrrFeN3dledogOVDFS1X8SUJFMX0diYLgEgEfACcUD76K1mA7UlOJNp
QdRUy7km2Ex7Tkl83maU0/6vt0h+rrXS22+cYieR5/rrdlLgT4zCJCUWRE1a8AA4
uGTLZwPTBlqXfQ3bvsigTPQNHsC63wphDCH5sy4X3Omb0S1wa/bS4Gm68akzODj2
bhwrjXf55uMzx04IM+VzO4ZIIe1f0yrkRyDhcWSCBQTdR0WsRt3cyeLvrqWh6t3L
LiO1rV/UM+U93B379WlnLbnPubvFCEVz6GFvrSDZi1OYmxA+emDOIrJAemCbihWv
LNj9AR6TwyhsAsLkO3/UacZhrqTMajbw1ZEvqttg3nt5AgDPAm8m8n3f1Htg/6GC
SWnn5E50EyWgIst+cZrXXp4tfEO5Au7/eqpodTWs0Akn1tByLou0ldOkvaVO7iXd
VzLvOR0sZE5W7lpy9SzVndRAre4zGQz7eUfaQytiB7cztqkWElMBNW8pXbhNbWtj
GMebT+nAVuJ3+8DSFPFMEi2JQ8a/YgvfyuoH7hgG+tuqU+iVqo1XLoEfBKZcggbh
btuz4ffHSjCRNqz1zm39q76JsH5v4qpU/7Idu28n8SeyyIZviZ54hUx5xE+jEMa8
Tns2N0AALG+L5QaO60qdban11AEDEiTc/PWSu+x/Xzae1hCcJ6GTJNiPz2i33LEH
izFfffJDPJzUsC9l3uhMZo9eCyHMw937p5/3FQqFsiDUDOCL7G1pimD1vBCoKm2z
3+dM9iTtzO4NWr/UzENK+fNmCvFUzsxE0sYPyeczYgj8zeMZmovEh4PRaYw7dlQT
D3S7No2nHuUpb5Idw0fD+iYwa2KbZxqVXzVXOOoqfvvNIeYvfz6PP8qyk4N2C51+
jaAOPTW2GIVl/y+UToRwHo+mV4DfR68ox0RTpeS0FuQu4J5IvqtO++q4/wqLmg1B
muZoEmBIUWrLonkeXTodOG33JwcDqLF1jvlaBpfXUboR/ARi1FF7ca3KV/0kX8l3
fUlWPl+QJa0DsCmBOPtQp6DzFtxxoB3uBpBTDJ+N3715m7POrJWqZhBka9BjCLBu
ygIVidBLMaYdSqvbpGZKoFj9JY/bW0ElLQ/fUN0zR90/TID3PapL9io7/oInvHjv
CwHsZz7DDo8rdVoEw7PKOPAJ+w81KSaf8GXM3xd2+PgBqYdzQWoWJ+vo3yzaeL2w
TbSsDQ+IuAS1362nUn56wOWMz27dv/1/9mHfa7mLLCYC6W5WEvOIazg+/ZqY3dkC
cF3THsTZ1Cm19DtC9o4ITRcHYrgehp7V//29Iom55V4iMG7sAqNt0x34VxWqx4wU
9ev8/jmmKFB1ZkBYRAN9CVvs/EkFwR897kTdvf22MT3543K+luvZt3yjLllzCH4L
NwYivCspXCkdZmD27GfOWuZnKEPVjKo9385KYz4EjRfBKrtlPM5jJHGCM3TR4qse
qhEVQQN7QXzAiCWxC6zY4D+JiVlvIkK24TcJ3o9ODcZ2h8ESQkJtJfIdDCsH3iUW
jlBpAEfsuI2AvmXgYsq00kM6YC79s127MA7lRDLGTPWnEodawjflTHvTdkrYo76o
hYVgOQ8hamOG9KEkSvu521ilXunWlMmCot73BAej2t+PpMa0mTl+4Q5X114ZgPAG
T+9WRtIrqNk9oyZYCT5Y8KDUCq9Qg7uEcLupaKT1n24dMAXygJgoTzZADKdaHGXW
/mcPF7XGrYLtD+a3NgbuQjnsSNyCTuAUl5hMzzRaa5+6CzIxAgDXm7uDaxwsJI5S
mym6Ay8F0bzAMoW6ejQAGJxfO0rSsoKxsKKNtb3gINA4s+TsnobJrL0VPWAFJdEA
BAkGaKUfHnK67EvPxEz/KYZ30HPvsHBg2pJIL5PZCqJUI3pPyboxlAWapZxm4FjX
DH7SFeq0md0XkBhEjyj660TgHYYyKojhFUamha+zAjk6b7helbCujMI9x6PNh+N/
U9+oAH8JD6gAKZfqFRAGSqRwWtgTOv38rnWFP6LJhnb+Q1wGUKIo9+bArAdGCxCB
l1B1jB6kfGUKi1jqK9ujc3r72vSt+K1o22MjwLSXeK94tbWExCHEo0mxFAZ8AF/n
XtnnwC+/CE/WzbE607MCUJmsU+pGj61kkRcMBH0zruPYbvfbo1U0007dUUwSbOQ4
D2/+Is9hZpdnn1cmnMq3laHqJoc2jPHona8S7IiVj/NdbiSXu8THpHHO8Dac7LWP
/6/N1WNIFUEabLMSK0lhDQSv6CuV7P6L9NyI7zCbhVKVgn53yxjHkPQVcqWXkjY/
5/yP0A/modt/8sPf77sHKGSjDn0HbWZ2vBAfPcU3/NEbZNvtGW+lU7Ke/pfWLXPy
Nd7Timp8W7HbxgxM1J4DF10vprXKL64EtqS566IpCkYf4kKb29+G3GKcZ4zu9/7p
h0KHEJSrYR712bwyjnZhbhBsn76JaQchup/+dWkyKDjRZLY2HpJIrFSB1wNQkMNP
uNqvCfZzHxBXOfYZpaWx+WxW98YdXPk13RxdY3vT4GLMGGdGKUXhA1sWMYHstOGe
o6lu56VUZEJ1vDwVF2R2ww8bvkSPSl5c2USw84VAISGfAdQjK60bjpC0bPQ5cTHt
CVdpy/vDVqEvVwG29csCl+qXL+/Egc8Y9BGNGd1GAZSVC3o2aF20Hgxzercp6bP5
47w5hSodrDphUWc1J9USpaJfMz7Gcn9c1agUnfPOXx2zfonA7TYLeMbp1laD2UfJ
EQXe4+Ccm+ILZIIkWOzrMT/bNSIq6sdmm06AZvYpixj22egOpYfIsMC7UeCJML65
ZZ0QVIk+ldP46m77chbUEA8PgB4YXUZg4UfZJiPQsvumYJyRXRR0kK5m8p06S4H1
Mp/aPuQ+HCx1WLiD+Exm3geavRxkHbsX+pxVC92ikcxjCjm1FDqEoXCT3xJ1fTQO
S/wbBNX0/1HV9sjYPo+6lfx50LVWCvynd6iHF3G2XxGohkchHbf27HflKfSlKQ8h
l7VJCsbUbX+WRt/NYldk9jItr4yTcPYcixP+9ZF1tUjM1NFZY7fD3RVFNcZG0FYX
o+uxipNMDoQ+kv8Z3F83SxnyKZ2H4jR/uXwuHNsVsdxXrXWTOPJZ7/V4vqnJ6Q91
HAbnTXdJJMaBCDD5Z+eMBENzxLSvrXb73/fjtYkjJDV+kRvSwE8hfOBScLW8RZNE
amc47WBMMTM7e/ckGXexvzwoslMkfuZT2QduM2HkeGS5lD5SmZMHUnTbHhZLfFOY
vhWtPewFM2z7+2gbJmYLgBwu40vCQpHWP5BCwkQGj4eBknZPFcz6OSvTMSNwwsO+
H4sV6TnrKWgNFDTRC8iw9W8HV2QC+V9yQ3eUXkVqQiccF9mTm9czLTmMtf6z8X43
kf99MZae/HghywCRiIZRHCLaOjSo5mOqgwT+2Tdu71mKd1RVmrlmJ0FMQzSnItDS
JiYbb+IhkyJeu+6Fvr6G+fH24vXlyMy7dvPZRf059z2t7iOHK4px3EMrc30ruE0c
1E4zwIS/d3/dsijMVqAo0+l2UPyjUNoBOHPpOsP9ltyaNrblXko7d8Lh/fY3KS+Y
DYbWujBc3Ey+jAVrfdCTye3nfs9GOsEJs6jT9DqcfeGksCKJhFTgF3I+lwwuhYnV
qZk0ize1Sz4chvpKTm8lfgl10xhRDBOupky1lqmpTWZl2zHmAJ9K3Rwot8tSdT5L
UVSQueuATNOzeK7O3ug8Eclhnig3eOWppcVS4kX/fu4bRqvtHQB+8DdYnLJnuFV+
nZp2U1g2PlsCsNZkgTw0mMFdKy8f78O1m1V7G3tT4t1WNRFvnkUEGnRMsMA7dj9b
ialX9kYQkgoWwB4yKYzjnYmb/n3u0vNEYuxS0SK48Jzh0z7mToqPOS5DW93REnyN
8OLHO6HBUkJTg5huopokTnZ7pGqteOSr78YjPUzaGosn5l3hEWL2If0OKReUP20i
mQ81G7q1mQJYJ4AP/XO1tGITWeJsQM7E1RWgCXO3j7ej4GQrAfAZkB3vwpJ/63Si
5SBzSOoYmqPFbx1l+yFjfLcE2eAwnbm00gZDw2kABar7xQoQnsC6LqManlVqrhtK
pZxPiLOjaW5u0zuFzCeDNmWP7tDGhTunjWTY+ZZ0fuDJS0k90ciQieTID+jZ7Ixb
YyFGWh/tmSGYutwdLuPZS0Z43kFbG8HVGofmcblSRTQJh38r0Mx+tJvGDv3WJCbu
19ohEpTp/NGilraE09UMoH7/WsZ2J3rvlHfhXKu/XQKxuL/FL9SJua7XtWsiVCso
YgZChvlJea0P/bUvhbAl6BOo8V+EBq5m0BpWyzGeFU1HYyISe0UxlzJvkCsAV8AZ
5wzVw3EcWbqj6ilOgJFziPCNAdEI/HZapXtbp7wWwDhx+Ca6K7Hi7+jP07x0wyR0
87CtPK4VzMO2p9d8LTNZZJ6d2SQXcGDLYitO0say2I5LhLZUf/teQYoZWSCMb0Gt
L79IKRXHa4a+MU5gbs3JRaLFVN9+uvqmGv2RrQYLO7nPjOjkSEtyPwFYb1r+dqHc
YajlrwfMXMiLFbGkUx/Iz8o8GPNyA/9UejkqNiXhye8g9TZ1v7IVo0B5JZIsJwwM
Gdc3Nfnx3IHOQOpUyZrfy0hBMrPTtuc1u1BhRSC0Us2px6mOUtT+8tF8P6cWb0Xh
HNpcbIFQHypnd9dXPBmqKsexXoq1ji9OmMjN3DQkfRlj9vwtuP44qfczqg8di8JV
as3M1woE2Cxk51sPYckKlYIWAPfwozzruiYDDHrTTFNV+xERJS7iu+5BFHCRMtNI
I+0ULQCI4FGoyhsVNP17VuKUtCNDptryJim04yk+5oNF3PUXfhevmV3jJ0S2idkQ
jtKzhRtSbpu7Ip8gbAc9eQE5+mU7+R3bJKWCDWP4MzD5jAx8ujmu2l4CMVzXs2zJ
dpOygpzLXXHxLspSnul4yBqWRwS0Wu8s5RK18M3tD7aOGkn7SaGG3a/XxDPZCp08
FN9IXApAsC9twBvly1a5z69XRlAd2puQJREbzrbKMA8MBoM4y85F3wXrT9jGXs9Z
Em14vLyaGBKTPh7Ko1uxjp6BfDebjQHp9q2x+v5qBvgedRjdz8Dofqe/6SsPGq7N
kTlK1KZlJ8V1gmt14sLEYn3HXTp10lF3IvuKMNnucYU/Rkc11p1WXHnUgDEZPKYh
k03WIy/WIe/3aHPUuxEgxu4TQCeWowD4Bbuua7HGnnOfvmNRZYt98EkAduwu80i6
Oa5zRYl/i7yGZuJAQszO6nRxQzcjl+ysvOLAIWfWcgy9W3sFv/tg4+s74dEyoIaM
ujUxaxa83xGPD5VaxRuXzFn08lu1hylf90muAmVYW0XUkMcDbB49FjMcbuuPMQ8P
l02tBIvaoVKPz1L/QKcca4j/tvDnRc/ZRbwRarx3GJB3TT/5uvLl6XjvrLMd2KAU
9B1dwDHAIf2qzr+FViK4LTiemfoPf9sEtTlYiOvlGkjb55xZU0KpJxSp9c7nTMq9
uyRSJKX/lEEtdA+205G02ryBCOvkNkHNq4Y7bbK+lceU4SdZitdrJ+kQLK0fbvDU
hpB0ru4xJ/VvPe/AesjxmQW4fiPJMxsH+tsm96cDpZ6KIpleZB3l00BxaIeqUsGS
FA3YV1oZHINV7uPxVDn8tEwQPtkskQ9OzrzWD5Du2UH5f+lvEw657MmQF3/V+VfP
6GzBTm46OmZbBISvFuxzNz0aJwghDZX2RDs3TB+JGy829NGjbC4s3mIsN+DtUMt4
3Nq2xYF2zlUFjjK5aNAqwa3Pz0Y91Q3oRLDLBczwfNr/6vNjjox3YhDcOibJ7dqV
nI3huqT3LIzQMQYUHo9CJtMb+65irvRzNaeg3qAZA8w2ddHMnlbly28OWsk3s1Je
gHy0sMGrlcTv9LC4LDv8YsmGOUt1H69CkuEIMvGsarS3qkUzLPAlfLbSSZZqw+fH
KGIeqRrezFcSgLjpG5GVIuzhTRzHpoJUif9eu7Savl1Q6I/zNnXshFHtjFUSsLPT
gTvQp5avYS7c6qYefxg2Fq1KkkbfMiEg+XpSyXKIZMDrVTFppJl4x+yy4RFLydGu
QD4dbMz/54d4To1ykj8QyrAO9JhuxbWAEVgoSq6SMLj9/xB2qq2fva3wwnyULoMT
WZYpHXT6oyGH4mdgfHX59l5JDGRELLersIe+MSX1ohtfwhEUNKLnVJvxGgFcOhRK
QoWA14SZq7vT/h1HwAi9QyejPv/e20Hw4C85pOLShjir23CDGtc2KAfFT6mZqH4d
jh31vDY3nT0FhqrYp2l2Pm00WBfFhUyql/Rah8VPkV1wJSkwCTe1kRSskubgVWmK
/4L7DyXS6vs67/q12GT22WxigprO5dJa9oOBgIXfVzVlz8OorRV5y0YfLPvn5Eol
mrqDBtESY5JVqw4zucj8UjMbIqLRfzlTA0dsiMJowQtqZR2pw4FQHbTehYB/lWp0
7zus5Hv39MlkAB/huVX7yqnZF3j3YkvHfFoxEch5Zo/eHEkKzgdIoq5EvybJoV7C
w3cupimrARIFXRxkeBdoA8ckfuqW7g9qk/naLUcQ3B8MOdfj2TCuB65S+MA7jjdm
OCdTRxPlfk3FDTmG4y4OExMNsc72vwgOSO2lF5/5K0yBvkG7nzkWMF+HikqCkfG7
T2I4n8Q6IxtpYspYqh1c5brofM9kAgQMw2IuHmjJJJUH9iAxe/GwBJQJ1vxaz+HP
ul1NHQRW/6WI7F/+UhLseEU/X71J8iD+FokMrGpBjH2A3anp7Jui4NDJWJK+YCqN
N3iXEx2/IG74wrh+pCftMTT91wcXEM+UkckyTL/XYT1JPlwRUk1UtV20sBK+k6k+
/RO1TD915lvhKNtBMp6JvEu9EBOIGBiTxLwf94mtMFlQ0JaJGB0yLkyzgJTZI6Su
88/+OC9tEaWosBQ19c/0sgAgzMHYQoPAkKamYAK3eeJ8rMBqOg0aLOOSmMT0vqZ6
TBZsKKgS95A/yFePI6xA+c0q/WQTnJfUuioNR54ykZ5FRp0AGQ7i5DM+UqIro8zb
P0h1mPP1O/0ysZzKFcM3XhLil89k5BRRRdfnf9/b7jgvk3zI27AbukJkL+L0tK/U
WkyODTwKKP2znIEQ/6DstJ87hEtmkE3ohMMJKYN+wrdCgZXaz0X4FaEHIPV0q1Bv
BOc3CWQ3AFAUaKs9IAWxkSPmgz3PyW/F20rXx7MzVp+8VR3PxCnbfKQXcIZc6ZBg
UhfwoO0l79yQNXIBmlZsZfqBliu88bLnfpgAoTVcJ0KbHA9vi+Hp1Fn3i5euVRx/
9TVlBitYN00YRW3YC9Hrh1xenHEPu/ChUbu72IteBCH9P4dRBin/ZI6PFURw4lDr
JbX4R0Z8hXOuCA8XytxZf8MASm+r98OWBAnMU1VFGTMHI6mah+NqFfiK+IvopCUN
k5g9v9i8T3i2WBnSPfgoUv7Sde5QzhaXPOJMKOZj1EfD/gglXuyDcj12PXjFac+h
58jfNfTXw51WIQrg2b03zX6hQueUShiVWXXyo+u5eRaSxrGTgILQwSEy5TgDetHX
m2HJUjD+PBecTScu5W53I8an0qecsl9XHL/0h3q1rpZv2n+jUc9PFXqqhRQT/kor
8Qzvf9y1ia3Ijudgve7bXnhOF5vW6Wd9y5Fk40U3LblocgiXHMH1Tdx/Ia7W+CDP
d/k7628UYK1+GwoLOFKjXO3caMNS0eA+6/2mUl9SnPxYPH2w8WYFs5GL/l/umNye
Dk/yPbCjzjjL+sDfyxq+GpI1O+/opabPHO9grPnuS2s0j7NIzmmZs9WmrWixE9Zj
te8MduPcUeOkMzpJi2/nj2S7ZddsT+t3W7njJ3AGUcLTv61FUAd5fknwwfApVLfb
w12skRhpmrVV3NWkGwgMq35c+3EN4xR8HLXZa2D9VWaKn2gnv7JKZIzb5JdqQbAm
IUm4IvCXGAf+JeWKzjge70sIUJEcSOAW1Xp64T/o1dzPfR/8awZVQqvNI3j12xAc
S3NP1demt71GjJW4yhMnkSp9HoRNZ85XMjQEsogm1ycI9QHkXHXIO1FO0qFCFW01
DSgILl0r9zAbtoRPrfiYs6Mb6nEhAYVTcMIG+fBwXUGJT3r7rnrnxv7tfx8EzUp/
H8sP/CEbZ2A6zkWJgb6tU6eui9ONr8XXwq51B52S32/zw7KPsgB9DOL/yFXf3Jcu
FtzBJL+gNlPjZceXoI6hp+omjF5GjWEHzYHrprDQEkKIPY/FCN2z6G8LH3Pnlw7V
iDm7ojuusYuvR7FsxW8AC55tHLowbkgea7xnhSxF+C0luBYrcDSG3DW+4oXT1Xw5
wZ05gy9wLrbunHtBpl1R2a+zyaYf/nS2frvVjV9OULjhaUjt0cUwbCZxPkhe1ul7
CR6vydEbAI+iRXPrNkAReT8C1YRD7UZaEE+hZv2MKttNmdBRq+Duapf+iADF0TI5
z0PinW98p7Tm7FI1i2/70e9kpwkN3h1Ztt2VUI+F3qfFKSeMDfywb/CS0Q5nEtnj
KHnFa1gW1kBkEcERbpb+DOyoYIGcbHCHyXlIrZJP4Cw3caeOdXF1EeZfBWv4faXm
AaUQuhAMQXmKYoQV6fjQVeKUkEjiWTXRVGceSkvaLB2RUOsqxNSIPPzvDl7HHy12
y/3VSmiseutqD4atcOFHku80ZKrb8geRU40pRyGwFhXcTgeSQhmaoMK6sgdaTKdy
ntcmwmCJWLpSJQpPzioToSxE1ZFoHqtjyuLq2HE42jhxKi3cL9TYgAj8Pq07BRa8
OJCBJCAJQLuUYRW2W/1J/2Ovuwq05FVcT3RWmJwsXYpCLCvtx5YzNKR/Hlig3fwQ
dBGsW64qF0eR+oJcascrNqzPJ1/TkxjLWKXWMWYVJdvR8AO8+U8ykT42Vlbp1u03
37VB5N6ErryNF1p6bVqifkBPV5ddU01F0VcQTu6sZsnwBvacgP39KtWKuDg7i4Za
H99iJfOHEpxoW1xqZNCgL8UxR1p74vBj+x4CwH5hYTF+XgqbZfu9jLnb77zqs65P
tsPdnymkFjR2RKF6Ux8VSfPFZ/R7LP/sOK/sss8+0yMDwrt63X0lon81XwL5dki7
MQ5lrhqb1f+9VLU1Q9CuTbbgiIGuJu9iuQqWDb5YGXWDCz2T++zN4WdmS2UVdXFu
k3q0ZNoolynDLdJRTX3Oy1Jj6SqZI36Rz2MoDbUTu3CtMzqAyeBpFNLqLsuJtY7D
yTVlekdH5OBPt3IcGdhCVNZMQuruH/4R9WbtK6LHXYl+vciABliubx8vQ4fmZOwr
mdm2isMRpq8muR6/MrR2c+vF/tvnCBUTVUq6C6yziN2TtbXl6i9mOB7yjuaa/XaO
zYxmpYpscfCoRSZ28CMFM4aDUUXXBb/EB7KtLJKqOEscChPb0BgTISylXriYxTJA
boffQyvHmyD27ao5kAGkhb91hY6MdItFmLwfdt0ERTmFEi6wzF7dSGtJCtKTOeJH
z988deyjdchP09eBWax+YdEm+kpuC1L9WHL0MLyDlwpq+xPwVUjI5CVSD2EYd21R
daOkL+0izXiflyFtJgWdQIltvot7UDEWiwBhBvUNzeF2t3bRtHt68YUbHGQS9h5c
P7TS+/4djP7kSTczNPxwBaSLcVUivaRKydzVZgrQFUM2gId1mAv8PWSP4Nv1MCZx
1RcfQ+NwYwkPKlyaFhSl/A/DOxkOCc/3GNiOXu32kJhO59OG6VKS3VJsYDsaRvju
111Dikojva8A7PlkgeJh8eQcYdmR27Qe8yQusNiaQonfjgJXHMPNWIklzObw61/7
jfHjsbEw4broyO9fvQdosQPcdFk5DlfyPjbikGLqy26wTuKo5cDZy+EFxW0+K21T
18Oh05UxMgwkZhCaSVcdOg2Zi3DM9XTIAryGlUAM+jj6d2COLwsFgETkxdDN4I+K
YzCgUVSAHuqDDDhoDHD3ZDc3DzaMvFSwaa5oV/7he2LbfLuufMDIXKueBnCOdmMR
7HkbwRVsAqEX8jhxdAccDlcgFa1/haCBq5D1GrfpeT4EbzHWowzToSxqzKTeVuyr
dQWl8nLamQfTv8sx1R76pw9KYeyHcvegYYwgy9x1vEk7KFprp3E9yksVm9HFXkvB
wlQ2ZVb0DVtUzADGerit94EXxk/aVkmP5NyoIpYad9dXIMBbAz2eaNEvYOOJLx0l
L6JNi802tknrXhaDb93enMdZHwg5DT4VT/A7ZhnPBlagtKICzfN2E6oGN+9/9B5/
US4hyCpSfDrnx0tAZosap5ls+W2ZlsZ1YpkNTMw5pAXd6sh1tPJUgeajDsvIqMjt
wdYv7GVevsgerlGSD/6q/pvbpYq7EN/BKegWBCjn3zE/nitO2XYLAdZabawBbIMb
D9X950n+Zh6BdtTcz/Qo/XcbDTdx7Orf7P1rhJ4vCDPShwOti6T1P27sJzkDAxOi
ocZVNcRDxaeuw2z6adWXOvGKFQzRARAhXMWkIjfmhuBvJSo4EfHBcXwd0CSGrJ3E
3mNptXwT+vCLv9rZhHf8popSHxXpA+q/dUBVN4OeE9SD4ozdnzpp7D96KY8H2J7b
zXdbGhSbkBHAkbgqmEGawPvwwZxJbOyvVBIZb12KcGR5Pk1hJeFugKI8CkWcjkbo
lJQYLTK8nqbEAHZgRFqKZgDIsHJVoxqpPvoog7ZKR65bu58MM9ZrPy/k0O47XcJ1
qBVP2Gu8R4Ad3DqGMNwVkqD7ldknmnzW4LW98TcCZtZnvpnBT0eGIqxxMfFzl/m8
WY/4c/UlOh9LtfitReI5oKyCP7+3ifNznkJEpJXdemjKoKf3Xl/CUWLBQ539nRN9
BZS/3cUGG7vBmHu0i4e2oNkMbMqFvOTuba3MFn6Iij6Ra/dcxX0Uz1MZVTu36Ue6
PRzwV3CVhJQfjJlhcCmKDdPafaydKf9hLbPIXaqBRrChCHyLCKkDYnP1zYrv/1Bk
KapelSwFszH92zLlBD9aD6RbSi50WwVd6XRkYnmFlo0k9K8TYjYn++4EXcWegCWG
9zq1MbHD2KPATJ8dyjej/ITrJnMF4RlQ3qBFPrrzv51SKNZT876D3s/zmv4zMcdd
IDfv70dflV06l/TaYXNnuPR0ZVOZoVZMw7Mur2fo8E/6CufZw0hYtAlF88dDcXl+
4HD8g6snfzxkUDKtEOh215QdamWf3aTpyv1vl2p1kplrF2Ip33NJadenXQXfLC6O
0YpG3pVb6J/2RUBDDW5r7n9ONRgk7Rc/RoNbz+AHAtHw1O7ZgbgdNDefi8Kj8qI5
TuGNlhbX2KgEhtDNYk9+9D8mrm2qwyZJeO8BfOZap3wLjC8ETWqyrnjByrEDfM/+
GDgnH3usrTmSlo3XUygcUSjxkRosJIQnkLlPt9uSy1wZ4Bs98d2sC4nhA8U3HBfT
bZ5dQx2WP8hWhx6R99ymXncUvOin8ejpL2wQ/peo/X1l/MBGlrEi3jkbuWv8mrY6
zHOex4+2uS9skFUw8uGbvCK9I4dxe+WBsj2PxHjo0PIOCd3bFcEzHpZYjHLEcxWr
ZTtgbMdFm/5vytbqanM8EfNuqho8sbPx0MrCPXKgMLCYqYvCWDgrYoVaTYjQr09n
lHfYFyZg9UD+62f6N3jxpIdrJpFfZdpIyBMHvu34Niu+liZltAK4g7fCrlierroG
FTAgabN/K5OaWAGPaoun+Mh7hMP+F/CPuO45o07Dv0Kn9LHn9SSEpb5znCYppB8a
hN8L7z3ULtw7LmykBv32Z8ugpAlyC4fJ+GXdv8iAcmt4mkHDJz5LQk0JgfMQvdyt
ST8Rj+Bk2W6p8AnTz7KT0nlhhfjlMLdcndygKsv3Jqb4ZWHts5rX31WEosEz5uQ+
S39W0lxjqDXB0jgXAzeWgecw8qSvTiT/Xzscw8J2trfdS4kGkXofYctEvOVOj96Z
EP2TgPUieQmhZyDQLN59hh9rZEHMyITDX0PIb90ik9otudwNUNhnEWRTyBuJV7N4
oBisKOkrySMu7a8uwuW+2I7tYSPLOlPOpSVFmvkCf2MGz7RvdDexL7u1N8/OWn9K
+q5MWmEUl58mosfZqys7JMLpsmL2LYxhlQBPfiK+dg91OUffKcH3TxcVfMUNzcgl
KmH43i73HAPSTSe0sWeV5zGW5d4nsbZoq+Eh9H2R5XSG9sOMrnpo/7bGQ5Q3Jmj5
F1vTxrHVoPTF8cccQSu8r0ZXqUMI+7y9hrh2ABIj4O5czG5vx4aI5BMMP1O6FeGT
uDBAS6NSnjVinw06X6Byen4Moy9E7k0RdpX9dUtavihERcNAEAv8RoNWodE9vXfW
TwZLOAtXwlU07DIUZQqal2rxknxBYnWlswZvjRqOXg7NsJHtxcuqPCew/7HLRgIG
fVnMCP/DHSw2F589f605MnAhQzxC9ux2zlGqjl+4xmfx/uny8/NOTG35tsfjpugN
IcXiG9FoGLwy76xnVLKDUS6mU1v4uxruZxcQsKvKmOn3wvkkHwitr8/br3qtgWqs
/w1nkbxC1WLd0xv1+HQkLMjXT/h8HhxXcL5iG/2Wd9CRh6bkZxjifOHuVXXT7Qpt
eHVZd3TK143YEGJi8BdYuLxITeGE2UcLR8C0YgihC9H9GBeJTiLYqBmiDk6ABLcq
I/oC3JOfwUvr0X2VyTFGyyPFkl70F5IAMKybYJHyad2QSky2tFHrgKVACSG0nVgV
ERDIgqiRt7mPqISAp2ENdSlivhVndWq6rB8QdJTFIfzndhk0EzehOZczcO9cLxTF
RPlJi9UFmzV9tLTbitbDa0A4LYKIpLdsh3Oc+C2gwN0Yj9KxA2MEjoXJa4BfMN+5
d2NYN/ZrF5axMT4mGnaNF1UlIYqkjy12XSNJtf4s2CHeynZEO8zggfoppw9Jpi2T
FvtAZCHnrDHduSeQPLEhfn8cw2E2fdS8Oia4W9kqfaonJWkBk7KYWMl76C5vUzG/
rhSMZU449t4u0KKSqH3Qwi902Xy+yLTqOM8d5Dy1LmDseUVUOi8dqKOH+O3xBJED
hSfi9QSuVdVDX8kFnHc31/184WjRISvJ67UF+icNHtoPlkaEPUB5Qr6s1neVQWM2
1NAyNlz5a4H5H3+tTRPKlbqF8jO67NrrUW4wohNMJXFM9GywIpebCq9Uux8AbFWB
wwE7W2nE5rGZHBoolOGLLRMTOaE5b52KOx++x5tw4J1w49aQR0LpMe6PmNqPX7/1
GgmE40NIQ7Q/V27RhG9AUcSZgHlBEyIaMQz2yCwKKh2W2TchGPk5f0NQ7vL83yCz
l89tpba8rFWdT4jdinzLZbofa9az52xHWskpE8t9QybF5Qnl1ynAnoYvVoL1HG88
+I9J21mGUFDUvKBh3Va5MtUVet406rB7JuLyeQJP4ehyidtYsGmKrLHPQ+7KqXP3
N4JCZ19JD3dMhzg29dTo6s195tVE5oUgnH/XCNfQhjx+AcrhdQnRq8qxjtigt2sH
BJP2frEt9scNbt6LOv+VlbwQPQYtiLk+BEtUuAqvRi0noRHWGMfX48yevO30ZtXK
XoEoBvUfYpwatodeKLTa1QrO0f5KmpV1nj81nhqg8JuZMYp6uSi/IqqNbbOSYpAU
hKKMVstriTFspX4ginthcRLTkM/hInlyCT/hjH7E3v+jleaBvoTp8NTID0woI9kz
ZzfQL5jCwgxJXj1JzSQW4pXA6cm4zEO61oVhSiRjgwa3AoIzWWj3clljeVIkiPFw
g5CHztLYWldpGwrmR58oCZvfaMhON5Qw6iohmxda831oO11BpZXmixlEZLbV2GpY
t6cRBsxbZwM49p7S7dRdCgyF/OWUmMPTLoMDJz3Zeo1j/HA6Qt+IyVATN9ZBRm+k
oU4XEneEYl/PW2LM0iICAMKK+Gnyp0xB98O9vyYrrMvzZ0WSPAswpQm3+2A5DlaW
9pDApNK4QB1GKA2PvLDgX5Y3/6dHRaNnnyMIxc0+JErTW8qW1+Os6EZ+wzj8Bf9n
ynDzKGKNC2SvM013+7KRgqekA7ptbP+r+VQtW0ieh1p5Yynwz510GHS51iuj3ON0
LvCHEFXFBGZ21XggdfjQvnBD32iUnI7VnkKftYJ42OeldDx491gI8b9nCaHZQWfx
guWjKSn7nbYjCuve/rnKrnzdZv8EfYlksGbv7fJwS1MY8omw38nfnhurylNokGdU
5yt26opqMyM6GoY0Of8oibzY8I2Offui4GoKnl3GJsd4eLHqi63Kc8l7xI/25AN3
Blls+2P5lbYyVDT2NkUiYEgHaGCiR6d1maRde2b4aRhNB6aK+IEgsWHulU7K1ASM
wuhKbwDPbOvIJlUgndjRu4GdQvvipoeL/c0KFhxT/Xs+f1oS7AX/FIUx1/+n4yBN
jalMnKdLhB1OknMk0dBwF3VfcXmXjeVu9f8iXCvMP5MI1El3GhdoL4+dSZNE1aX8
EMmzXQq9719UcWN2ACpDKXwnuTz8gngny+eybUQtewZ37Rp4aVLjdiz9xsR8iesq
OXdeeDyBY7/jThQAZWB40W7GggTHi8cvfcpgBLE+PhacLm2hn6HaGW+EoxKJQAfk
fBdRDy+wTX/cx2i6XDi+kkmxw/h4s2Vu7Pj1Tmq+hGFkHG5OUg7n0On16PLQstWP
+rWEgo9wEynSEOoh8lgiQmPzDXV4rfUO4fkmBfio0czMJEZftNsc2tWC+uZ2/n4D
4KZOMADI92h5k7HcTIq6wn8FqGdBpooMDNyMERI26fRqr7MWZk/3vDxbrhRfBT17
RAN42LBUYF2l6i5I5InPwUwmyo5oN4X0ioezyZD+hbxH51JEjcYOfE91XKD03m3h
o2mk7/iIlwaJdRdqi5xz5WMPnAkxDq618TmbyMR6uCDufPdewwPz1oHfPPSlZfWQ
u1p6TCyCTMEGl0yaundtdmriabnabSB18ibq58r+cOh4OmMgeBxrORWbmrnuZe+y
ZHd4SoVtTNDKe4cWuiKW8VCw6LGJkhBZEqjV1jz3tic9BbQ8SdoLkKt6yyMGz/cH
jbhlcrhkWYwuX1tFi1w0lnLmkK7/eXcNYaNTn2BCA41in2vEiKd1eRMmiNQQ9G05
w31hTTsLQttmwybcmpTWkstyamjp4OJJpoO/IKOYbYpukYlYIsi/Kd1yaPP6pkkF
futdx3MdA1t3fRvMaxinK/osJo9+P4m54vLVLHs8Nc+84fjxx0G5yPolVx0Q0LKh
h6EyQdAjz+OH7MjtDTTsfTIlvH8zfXpfPSKRVcjxUJhLT/gNYhsjJIeRbN39Thx8
yBoqTEXoWLaM4dhI+wjwLZf71aJNk1tPWGP2yrquZZkaJ1qx1caLXxvYfcKB4H8M
d9OF3ajypSl91NmaiTF7vYOosQGzcNBVlhG1jDSyqUw1xEr0wCGWxNT4wy+xO16o
3a9xarSAezCsg/QW629s0t7OYG1bcxKLLIXv/iC0BIh8Uoc8USg1Y5C/GJ3ogGRY
9ftE3eFyPw1bGTLOujYrcSH38W25XSREtd/3GG4fRoVpZ/qJNqzkgsDioeRywQkD
yd7k6kahwiWUKfAupJ686T8njAiysHqJAWG4LxBMkuw+xskVeYD4AHfXXQC8wAAR
9SgOcvyp5G7Pt3qIYDn/hID2ohoSqkRLxSybQF8WPN3rNYqBbnr26+tbQXNOg0Ip
pMKb0tGdOb4fjigwlAhB7J4KMMmiB50tfOt+tQVZhVImxjPycRWvV4/w+7x21Ta/
Pgjnx11cd1xsnzoAX+hwUYQYw4LWkD4xhsk49VtnbI2eAolU/0n72mEtA32qptyf
S9T7OqzJDsAcvZ6GVd4Z2zkA1stKotmtkGh+ULe1+advYh5ZFNo9nlwMPaB9+/72
GX7Mpqvl8GThl+eBRvS0mzpwBFBThI99OjtmbFKJeHNewnj1SSnC9SZysIvZhg7u
CCqncTmxYePbduRJ20frpSgt7fEcEGC5KQsXPz2BEteSGm5+B2VhFe/I4A/XOlxv
c2SZZBYd1tRR7nFq5aaxHYTBzr46IYP7qL1G2waL17IB7rED+ze+lHGskWxtZL02
alVMELJEGGKRqxl5UnuuASEd0ZD0gA5yYh8gnGvAxuVeE+L2BflLmv3aIY64dWVV
4iNkg7S6kn4QAvG+ogThiyUOD7JrIepPakNezHvGSN70/6N5IJXvTAQK/QXtJfJ3
7pA/JNWdsDl7GviChGhOiNTyoiCnL2jFXTcLJikXtk2bKtatrT6CfpTzEylkWafn
Gx2+Gg5ytYckxBZv6z1cHAfruyBrtJ1iO+PsCXkw9Tb/rdP3oMwtgBtERXYpvpHh
kVsZAnLyGOrcsKuW0h4yj+4Ml6ZtNkUNHCJvjDH0fYtYDg1Gsa/GMi0vk07Ep0Ak
ZAGi16BSlCK4Qd8IwgK8lyfEZqbOTaSZCf1znNkUdKrU6PV6XQ3aEhmpnDHApx0O
DPQ5W10SmE5MwR1sUeXwFEMxXvTfiWq5GBUgs8JNL+OL0jpCs3y2K/emiNPconAB
bWW8j0FVJLo63VQxAwio+wEHAnDIFlgyMrs9HnuWbsVryBw9NvCJDmYg3JjOaEAQ
rVIaB43FkYeAZf0g58qIPZI5LCg5QLD4agEh7ZMbAAoVQxOyKAF39zxMD/vmyuqz
xy6eLLAhLt1ywgGGwJHkMRwPZR8YC7loDxrvct7RgdbKr8OSVfQ5hU1a3nFzBRBH
es2XN9SxK2wILcgAztqDstE9oY8WE4P5WWV80YDmN7OvoFDmvqdk2o5iQeyGSWpB
zuX4SuCfQ6ch3hNlaG0kfbIDvI/3siyrdSpwmlAIMbsvCCOwmXeFLcyEFiqz4Ay9
e5gnVJ4XWg6nePm4pM/BbiI47aj0zBPArpkBgHtpQpzEO+4+3ifUp0/l48oVZIVh
dVLnE8f/2r82djoDMYgrqXpeK5kUPCF/tlqlMsJGBHa/a6xNYUuXZ6IEASN7Ylah
j9C41BeVBoaAlJ/kImBwLZnFVLSR0eQDSHFIurfyDkYQHr1NnlgCTmXjxDBVMSU2
31wr8dyIB8i2hu9czuW0cQpuGxd8GqDXt61SyKF9jxrneJyzDzQhuThWkvji887f
OISt4H98LSKkK84ZD/Qm68HN4MjgJTBL/VaxZJYRG1tkeFrsFQIcEQ9QNNI/tIcO
1W3Ani6o2kcNBV7h29ACbiFD4bov+kbOVDAXkeRzuDgpPgFng2Ec0JMOl3+Di5bB
KEZDh75FHAv+3Ak9rignAzh6+Dc/04/rLD4i91oV5AT5PO4dU8bYfZjiSdxY5+9i
9c44sKocoxuC25kL2VghnvE8zGmFXu+Awposx+hXU+bAv+Vxx/xPq1d43dJTUSHn
Xt6virdV7tIsURprL2ou9jCyQ4rp+QzWQBjrudmix6Mf3BM4cJdxXXDaFbxspXII
XUQ9Fhm5Kkt81cCChD3ThLPaR8JYfckPXm/hgvFnIb10lO6jKzCcqg6eIcAeyc6V
rrMKYkkrq/Rdym8jbJRVKr9yuewn8MP0IA9URTwnEy94MdfFJNx7UBhaf08xhSRP
3YA3/9Yk7fn6rHJxpNjKoGFtZ6r6XYNALGoX8uyFZVsYvqogss8HnTbUnaeazBa/
W1bEBNjZ8JexKLQ/ueSbM3l2S5N82okL0pM1h0mutYT5s6sjJfYCRCHn3O0jPhjP
HQnNiggVBVmmV3nLMFxKS6+1PfjCZ+JC7bEzo8X8FWmGNvCaOK+YvKrLvbOp4Wzq
nG5SnILlvmbiNki/+tyFy8ZUSs5V5Nr6HihH/7wAkobOO3TA7aCbUWOc8e9h/PBe
mAkyyHgCmju+Rd89RpQvzzmjlj9eQFprL1NGVBS+jzLlabPW93yN46vtjoOObJB8
zhM0/ulh3avuTTk4kKByoPClD2a1lmeD1YPhGpcXjwsosT0PJPjYk27JN/8mJ+ta
MZtE4SSjtACCqVgcBtgYilQe/+IjRiUxQO1IcweSH6hM8L2ddDuKVZ7gOjkSac2z
dRlImuH5IhYH6E2jFdav6bbHjECU11a2rpr3so17RstvscU/J9lQtq1pA14c9tVK
PiNaOe37cJf3t+5HJ35cKh6rNVDR/ITyDOubewnL/CYJc95Rn3v+1z0tdK12anIV
dw9hN30wOaifd8pOwiPrX+GYx0Ee+YYw2dgP+gZ+ucT9ZWR6KslDFmOg7MiIE7rj
dLh6pLKRGwhYMCCSZiIJ6/NNvOSqmo9LIFb90GTZMZ2eg5pTcO0KQNtkXzOUUREI
n4QKkxHxmm2ti8VYvoLWIlFQRgximd/7iR+zysjTVX+xvFu9LG4LGZ/e93SLAD7a
03AyjbgWdhlbmRcRZvJK61BuvTo9x57gok/zBRqwE7yQQ05Jzs3U/LtXTScHpKi2
hWfqbZ+dPq9ttAJR7piHfZIxXxFdePPZMFYJjHUdubpWtk/4tYTv/zru4Dy6NCv/
6APlNzGQbby27zr9FhWYWkG10OIb7eb5BUI/9508UjOyy16TfNpDXx/SRF0RpN6Y
nvmoXGighufzGhkzmTXmczHRRynfbfA0u++4MMq6AaYIaWvU+DOm/Yk2aMC/6X6y
pYLbdvWcfAh4YhJWlmNqmQY3eaUHye9FYlDZlMXYwGkbsCc3qD5WQ+U45ICZAFld
KGAPqSJtaY3wrRGox8oPRwqjg/MGHPeezHWEtOJefDXvVeHpyMI+b8N7Sv0JBqDt
zr6+mH4i2JKuU6I8Fc4TCXEif2l/OB+iDFsuCU3MZ+x8M0/4hvA4HBZD+Z56UoYj
6pHgze+2wcOAZ0mjEXcTzIhv8UpC9MuQUnHOMmgJFZTe6BbYUGd/CWxUf29eXgA0
fdtewbMTAAx2Fz5GzRbXNn0fuUP1Hbv2XVq/JJOI9L5pFpjxEQQ/QjH+94gJ+Kuj
zFe24iOEkZ921MBKZDZub8Rx3yMeBtyyJ9DEPDS/xu2pyj6TmwEo+ki44PAAX+Ix
zKGI2ZDHIpebOkVudZB9n0CXCl5NUxd8XcZiPyQD3vv0Esqh+tSlDOd79Cs95u72
bVSvXRJzRQU+NhEOmyb8XP1fBFnr1PpG2SASglqByeCjigPpIF2oCNfGJK3o46bW
CMfl4VSGU7EURcs5oS/K1O7yDYct4IS7/b2BY/cHPoP0jXBgD3pIbQxcaEDXY9ds
yEpbnOG1IpGEJH7w/J8zL27mnF03UXpGZBOri+Q2gZ3GLrV+XHgR3UI5NhyOeJ3n
TsZ/pvuRunY6CqE3BNlc+0ScbNvDZpHhgrLf/p9CmL2mnEuibCf0sJzjP3/CxaSC
mdTku0Kvja0cg7JxHGYv+81A+wQ7AKllE6g44PM3GmR+YtztT3eJrna9sby9ViWh
hLwUE9qGBjyD5LGqkYguVOz6jsn9Stqkwk1yUWgKjFUQ7Fh4WWISs00btQtccf1i
CaGT5t7EMkeinDbLLAYSUlW8QmJwhpzh4qgDdCQgcm2iQSuJWNY4EV49zhTJ7AEA
SVf98a3/Nq/xjaggf1g+7Cn9PItQ+pdi/ulQSkHAmu5MCN11XIhFRLwHxNkcYVu5
Hda0QIdZSN9w//49Fp2+W9ARV6IVOfxWCrPDiy2ClwPJw28mb6CvbZ1Vyk6R/kY6
fJeykdR3OxWYMbG0xcrP/lYjcxAZaG/PKERJxlS/jh6T1m/Cc7s1hQrWkZF3zz+K
iNfEMz9PF4DdGA2bxx0MZPVNnAguf/6IWjBlvZ+ucupAk0KZVMnDjT0nt/g+WbVo
tzZU7IVhT1XdcizJ2Nw5Ti6s+qXjGtrLCTgN4YsyBNf5GMj6NVSv9sQifDgKfBQN
NrjLlUq+QZ5aZGN8OjXJy5hDHC/rjKlBKlUgJS1nzkJ0r7NEYoey/EXWDP8mk99q
WIz//bwiCjyJ+xtUxCVHFLp7XWLYAv+qbFlpHeMKTqcNq8JiZKeGdM5XAGei6Sh+
4YpuoMiJP+gj4wVA+30+QRhaAIDCibJhGSk4KkBKC9uGTmDtMXn65RffcEKhiVHi
z2IwPIU7Q+WsR78a/NNA5oH6z65zwc/Um76NV4iFB5q2uaqq5KMYg8P5sL6ZHAS5
trDLHSaX+hsG9K4woWO+/bJowc+peKA39NKHrF54vcr0IqjXQYiQN/17J4Gi29i7
X5IfuXoCVY55Rc3O5iQY88fwrT2L0UfJgrd9POPhgIcPVF/lyYZeK8wKn0OGjQaD
ygyuTB3IfFfd2VBTrxmGwTgQsyaWbbuWSCsZXqCIxLP2Z4smh3ES54BVQnzZCRVO
++SQ43vms+3ixo3WsRCrk2aRE7Hc74F5Ga9hqwElvC+2IjXCDxM0WbD8KpCz3FaT
wDKAuE5IUrBXKF2ikoLEGvWvC8VVgDQ2ROzcX3CJSHOk71YetXl5sq4zNOqY6NIH
7vguBcOEwDHsKC9qlP+W2nya03aehiNkJUn6bLbL9rAOcl3o6D8ZxXeIsvmge7cw
kfzkueF5ImzfdIcU4QPzdWPdIxDJJZGuLXY9yj6ZcsFJLjwRdJKxzrXUWTFid9LP
RhWTko5jrCvyRXJmM1Y1ELvPExIVUWe3mKWH+pQgxyuPq2zzWLHpYKdGN3yUVzKH
SWKzsawb4CtK3fBdzR89gdsOory0OA8AAXvPB2XveuDji7nqUVSQtDRNZCxDYBxV
A923KhSGoCThifekRQQmMe04iO5rpx6UZN/sVoD8e58vX4OAFSNaPz28iKB2bvtQ
qObpjzaiHqqvvhv1ZPW41NoZtF/zFX34xpVDDJp/3PYG21vXvsZoXM5KOMZxmjQg
iXe6SoeGaPc4p3RNmTcKz7sBFksPixAZbXxfCwVhyL22f8J9LJysHh30KChLSDGP
lKrY2vdcoJ+q7FhPl5KMRkYy178Qh74GVkfbEOgmsu3kosEumXDaMg4YeXE/FeUX
8kRIQonUblco1x6cSLw3Swxol/h4TD9WzwL1XzyHOlFb+GHKGLXuVgNa6O3OaDdw
t1OunyRi77I2R1WrZpimLGQytat2mMpfHYF6BXGjBTOpfZjWl7Hc2BcOVx6J7Dho
DvLkjNH3AQE3AJY814BSSwGfLnWBXng587VU0MhvVRfK2FuFG3BdQRMilQqoZfos
UEo+a2MNB4DmdYmOQCebMHHm87RiPU4x5hBGnMWQACOzZbOKGPl89IP6Rkto26/y
Pi6ri58959oYJKO54Ivts3X0oWeX8TwRDrvaSBP7vYpLH+6sIYu9F/X3mMgOT8Zd
CBoq+NGtbS06FQ3izzXI8clyDGd3nt67dH65B+NEwFifSI6hAnvdv2iH1rgBKxgy
bDh53C633gBqEigL+xqpG+222cSr3EEH31sLx6ygRRjCJ+sgC+mwhMNqfoh7/WJC
nwklwOEeKbfiaoKTwArG7WE56P+LJ3TSYSbthPeYaQ1+xeX+XWfCEmKx/AROe7cN
n1+lzzVDAfK97rzaB/3RdNgtZEeQcxGzWTLvqce3Y0FBWh0WK2cbIajEtXmc+wGP
LZlOq7OdPYThIQpKCCXn+eiaHWzrNj6roxRoj7FfEPLmbhipOOxJggR3sllk6PyW
l/3TBDIgREnGC6jC4eu+fKsWMrRWDNI9LPJL/p4qTj1lGyuaqPBTsWwn7qDJDhzU
t+N6xFVOCPWPm4Zy34o7melpwmjlEVxv4FopeZuQFKbbreHxVrgR+VuBdaZyXbXE
vffwtXr273y+Msb99lIatcHGF7kk6mCcsY6w0QH9ckr+dCepBmAVkC+L3xFj3YiT
rWJWWzYc+oZ6P4LeQcWlptldvszLghCWkXsEFYkJ3NwU4qF/1OwTL5262KjR9K42
tpLG0vQA0lRG10/w5m5CCTUvgpJPNWuBfFDUzOU8WOzBUhzmz1mU9j4OBcAYPORD
zP1+rdZyy278ViA0BaqCIvXwc5hgGMlwGIgrmDxFuwv1g4rOl0JZVYK+metT6qwU
A4tBv3j7VZPNeznCsMtRiLsEmIbXhmjgSmTv2+zUHDr+PzAS055tfWjpehWcHbJb
GTpXbNKb93+c3eRj+cCAjgRJmE7BYYasm+6NJ7cvM0ppZ5czT/ngLKZqiLwxgZaK
I6zTCvg2EJMKOkTJjICJyLzhPL8YqHlwWHJ7v7CeV7Ap5AbdkgF0onSyhjDltoc9
U+jBjemVOhGJ7qjb3usGN87g/1ulAPPjLG2urG9FQA6NDOrqMy21nxammc1VFb0A
+z83oLUQNRJX3btE/J1fDXJ3yDxoA9Zt+oOMcjz9/wCWiOfHEhTgCu26D0Uaetad
df8LQpMYEHK6Sa6LbYDnMK9YDiiMXhHvlCq0At7CkkVVuVEM4ZARDEgD9Ry1TPC/
YoJxJDVQLY4wsVBMNoKTF9xLwRvpe4/Mcyaydy/h/LPiIrhMMuD+nFDW3JW3+sFV
RpCCbzHIHDMsVXUFu3T3pgkCfL7o8wdh2xvYncoX1iXNg2smojxpIVVdZJHzUSOh
ndmPyehOV/r8SIkpHJwLpxQz04wQjIfil5chF2hjfkRZrMg8AJT9DTAwIeLywb7F
QxqjoObokE4LzMhKZpbVfZRmq7G+/xhh1/2rnGJCbEjF9BeU0sfNw2tAc/4m7BQk
WRNZRIDLNSgqphOE2IEDBBt1RWXU2QowmCZ5whaa/UtUA5t0wjxyMUKYR8u8J/nQ
odr3cJHZu2eGgFTK8iffmzuvtPnaJavQ6q36r4KoRlHEOHZnteKXqb0YMeY6DHeq
NjZaPxWmPlMrOT6i7JtVyPwWS04PG3PhYDQyM2ekBHXZYIUUD0ZMuPn2CZ03Q4sp
NZyT0d20f7iIP5aslCQLoehlrQP2ES4r+3UX/DiwhV6Y/gqs5CeEE+YpmWHoffmp
lSHJ9xxrPy+odqZGRDoCDfM0DDvGOcbOJ0PbGU1zj1ooxO6C90nhAjz6Jz7n2/qF
QsLcYW8VLKEPJii1tDayg3Yv0tbYsNLNKb9yKSMuO4NT1O2qpmrGgpizoTuSS2JS
AeZdDBbKy3x9N0F0eGS3doCtPI/Zaoq0XTZWCxwDm8wXWtNFYyjAxm3xCEBAV7iq
jKX/WGhO9ToiZ08uuHQXo+iNAy9PAVyYJU6jD1Wv3Wibrr/WEw2XV7VSHSaSLOiG
XtV4/SuElCYMrdBrTh8y53UMVjMU0VQjedJ704FQsb44RwspqjhG8LNa7YrU2zbR
hFJSMrzIrUNELDzr6ji+sL/fPRnb+xsy4myFRFMYBGUny28mx8EacQ2VxqktyYFS
9iEZmaf2eJb6iYoQk1Q/kvaRs7WE2S/O/qGuyvVN0dl+HcCm2E6WvYKS/Fsx70CB
Qei7J+n5ENwVXq62Dj6F53YjbJYWfERpGMWKFpnXoEv7P1KPkGJcHQtpI/whNbd3
ZANXNsGLD/QT0xYQ/fQWJ4odWJP+TUxGSCAyfn2VaJNKv3luOj2z0NZdHMB/Z9ai
m8zq1aq6xW2Pv8XdEbPG+hcgpLdMlcQzprIUuMgDtUemg11Xil0uoHC+RtNKQ8Rv
NJj0n7uZ7fDJTJIHrWxAR1poSk50vLNPgVS1mhoP+PSRJf2PcWbsjGp5Il/vEfLd
JtoUdp/EQK+yyyBexyKDhwnT29dqZzYNbGL0eKCcdBb8Jxxcyv1U24E5YiOTYS0B
prABDrAIqR9rdAhkHStz9aqYsi6L9Hlp8JUOWR51Qmi9LisZ+XqpN/Kw0R0L4DI6
zI41cuXxtz/UwDOk18Qunjl59+UHl6hQbkt/33shOCx4J8oGhsAEoFfW2eZXrd6O
VpwvBv4F7l2Xk74H0EBhn9zxYB6V0vYrhgjSJ7GltJLuaLujObD1undjzrb7MknE
fC1M62h56KMwpk/902/dToisP8xsm9ezFVmdMn+DR7NFUKAALqCDeVbp3Lpjw9Dc
gTAOljgKnOID7wsgG4qhRrYzl06LQX1FVnzXH5bHIddQ6lWayjAJXVYPezQJks9n
4ZIVi458q7aqEJiTrZW8BQmw+kEx3DPQP8tnY8lM3ZSN/tpBqdB/6dzqAxWomI7y
txbuUu62PL/5DmrkSb8PShH3ZzTuqP2U7WoMPlSoj0kYH7DYQ04VhG3MX3Qizb71
6eN+sbp9rXfwpIufwizHtIvzOehaQZ1g2zj3gwCiMWtOVElZfpDnwcR679uj6vP3
IJWQoO6PCHnCNLJ3KMd60o84JCc30XdY1TUN+aT0ncKZP26W/l92fLrx5rzhYGgL
mQGS23ft0c/GXcXwUD+IDrEixWopWcgsQeJkX2GBSNn4FdFBKthqzJambAQI/Exu
hQYtqM9SW+NDCrYFoDuiE6foOdALWJgN6c+t1KSFbXYxviFr/88ERUUV2DqERPQa
ITChIYUDHzBXK+NO9ngls8joPUZ+elqdInw+X8vTyPtv9bgaRKOnIclkhkf6lxXG
pFlKaVo//UXtJyD26jYmbcKEa0p1VGrDpsFek0lmp9KzeGxggvqzreWgX/v48bnZ
hPhzEpuMpuB45Kb3xshH0GO9ujYUoE+ajY5Wx0mwX3jak80xfYh12nmll/4lvm2u
pBtQYaFbxrMTqYqBW+pcCGlbN4m3aBYapIz7uktMAD8YNBoMWTLoXibmfw3FtYDa
jJMUiyFRgEzEeLwU8WKTJLOQFtNGsuk2o0VSHGNQpTPFVZqS2qTWBHieQnpUfQTR
m/O+HySqFYv9Sy0cAQt/JmQxpdGYZt4ChER3LxVN6m/pOcEA2qk5RnVofDaEDjqa
i8X5pZoZYnbL5oNlhaLk0WpduvNnLgy+B0A+eqqfFrjpuraKf4LHcRTg/1avpnoS
heINXrfgl5mE0hyUaF0/E/AZhC3qJ6BSEI67/UbnOmWhjh0NEVvrIJMX+BR4yQQs
USBSOiagDflfZmMsJiRBv9ejZ3brneakP5hisAnRCZfV3DwWDBN9zfn+ZR0v2VXW
YgMcplsxLBgp4Db4Jpzi3RX6CUWtdx/FDGfwlM19vccloY6dY5dna7k0MfdNI62Y
BJt2ejiSLbz3jL9+C7g7T4qsn4FQw4Ex8MVzPbQVYndJghrxuG/4/+N93sQ/if9M
9y4AjgYIPQkBjp2knZ7XBqX/A30zyqeS0d/yHqfQULdG8BAg3vXhHRnIhnO7AY1i
/9a5xWvVShj2pn7LCSMzcZIDxBkq7ZFhtfb678Dk3L01QFYuyDmc9B9d4E+A+/Ni
5cVdCrc3ahlALEAKNm6rz8mzhfP9zcWP0iGBFh617H88egs8okk4dzJyxoSlpECg
phxEBozAvIfx5VzAZuOumDccmHbZQTSz/leHa8pZgefE2Y1ZQMqA70EkHY5nHlmt
YMAN6tUOH+Q2w8tXAr0VEv/4Ug/JRaBN5c8AMMUf19vFz8p9ICikSLantUZ5zSBk
EVppqYTUaMka3rv0RBbAMzrVCQgcZy1qD8OwC9xsaqjrMP5sj9LIsL5Yw/757HLf
ET+CHaQG1hm7ssQ+w9VH2GVqNswAHjM52EXk5TB+7e/1sq7TqSKMld8yWHqOzE0V
Gfp9t9honmPPBPgsoWL1f29sMnfQPGBxsQsvQ/meDpC82MgPy3T9qul+H681C0sX
hw9VYEe+/PzBoF2ov4nQ9SjbpX2H/YKpAQigP4U6CELFKPuqyV7bl/77kjrYuCHv
ZT1trNYp6K13s5kklbKv1UFZikDAeghG8e/Q4S/tbtm6wUntIb+MlnoWPWSEJcNC
OA+/bIqy2I1nbaMHp5idcHZZ/0jgIFVnqjL838SAwFWJ+DdqHKevuFioustfbRU1
jNUqX3Dndw6rRh8xdpDCI1KAw+1mJSsSA6xRK0WXSosrAxLZ2roWhcqZmAWYjhrI
h+idiFMMjrcO1b9SxS7f7GpKSg5k3EnbmyI1UETcSm2hAGDoFuFVNiqkxu3iqMpB
nb5at5AYSL42zIc4a8xp2S0pT0O4FQIZKHbnsMklytGP8tfXQnzdIESRC7NFyvwV
F2YZqKfZClpkauqSEuOXfpPYsJB8SLV6sLr6oZFVcZ4L7X2t5jCtOvZkCcbBYaSf
zYZ/EAH77opUQiogUJJUOHNbUkN0U33IUpUCY5zrsTG4YuxTG0YX5vhpNb/f+53D
oljv5XTca+pULoxXcsG+Q2JYiNbqVN8wiXDCa4mP6yjTuPa4lbzcJolYY1CNJDLe
xoXWsNRhKK/y20pcP3JbzCIDo/Wh5f/QEGyxR/CVA3ItpmDHE9K4V1yoIseyFk+X
oS9CJKmcwc2zYhCs+cmJxrRh+JQ4Blci+UbCBuyf0hbG0KtkaY5zIXnpvjHVaIaH
9ZUyZvIapRGN3vYXE/2X+wMdJxqhhbsTaVXo44CaL9rKcC3eCY3c7nMW2Noqc+/I
QIukuhPAobvpmsPtE9kHf/cAszueA17ZrpDep8ftW7ujPbYn24FEFap1PwcDsgWO
88zyRqOU5iAe/Dq53S4uoZkdu85OYg8FnClCvvqg2dnk1DqGPeGwZ4NSgnSObPXY
R+rhwyAZeGyBwWgpUA485KA5QjUYsUAdxH66u4e1KUyIXZvqUuhVXTIAfhNWP5QL
+WIR4l89PPGnNd8GAcCMjE9LDooUYWVBG6Fu9oYrlZ0vudatv8Qo8jWCntQlqHQW
qOBNWpMGIZPvv2cu56PHxG16VtmYtOJXRA9scuSNGjO3gvtCrXhtjXYE9YOA5brO
KS7OAClJ9Z07NuLcphHvUQZ8zxpo4u07/HNH4KMjqlFQOnGCsn0f5nFnccNmuRid
Xr6yYuGGmZ9IEhlx8iKY0yxFA8e25liAqRhQuv+Qhsv2NaqTbpuVlJvKpS9p64MR
wm1SzjAI9JAXaF2+KINjCaMkmYuyh1BoVCniLz0HJTl5znZ4vn75ZFIgwbAlIUBa
4OkqTfU53S1wqhAHtujLDqjIZiQp3FLm6vMcIBO7Q6T+R/JQs54lYVFQxvBuEU9E
aRaQamf1IenjisiB1etufgLlD40NSP6EpFPbv19vUIHiig7mBUXAWUOBAzdpg3IV
UsVTKjf/txHyeaLqy9ytDR1pH8DuowxaAT0pkT8se/3O7tEKTkjcSZGN10YAcdTX
1xR7slXoQCcF2rrU8Npxzg1tA5N+Dsaa64iYkNZ7ZZMJ1idLlT6P2Ur5wh+lZS5b
2ybTbIzeUwQghvKBH6URMNExkftZR7CqsJpjMC3fcuIiS/iRSoNkyGuFD7XOctVZ
3YwmsYMZf2m3pKPUIDinCafav94F1CQF5eLghce84SuSLtuWrgxVDSqGmjW96i+y
OBwE3M8qr09CQ0Jvq6VTuInQva4LlaHDpwm6VN8uNMJe0R1ZFl9b4LMwYCgZHe7q
1b+q85zhBQmUy1cNGFWHiOOoIRx7Cv0+0r5Wm7Bld90xKipwnzdlbY73DpvZ1C/U
aM/mHZWkAorfZHLw6sgubKF4b+tj3WSYJ/y54dLo6a4znMBSKpOfs4d8l0x47DJV
Te0cIZKSPpL+ihH5zm7rWSWPYP2iUQAxtjnW3E4eo6ke1X0yYbNECNmnIqBomoxg
PirZ6P4umBMOtY0p+TVzLdysDXgGc/IO/NY7XmSBMo7uSxpqUk/DPm017GCmyotM
xHOHtrHuZtttEwpqCijuHPkFc3r+Ihgn+IQAJAy0CDpEW6q0rO1x0Wn8XA8KisHJ
AFPnHfgjcBlDAQ7xndoAlg6/Uhv6pGoU8BN3NpOptbdq8pF5HY+R7zRzJ8x1yctC
a/racEuIX5QTW0Uy5RatrDs76Elasf532er238Z9C/rN9vIqlQHFaJJOoylu/1Pc
IOEXYxK3vzT81njVMjtYKzfL9GNWLGv0w2Z7Esr4NonroNhClrZhbnhCdq9eUwZI
a2Kyu9lDs47I5d5VGIwnzNXW4IGr5pR0kz+sknQgmV85dzwdQmPY0UjyFP9YIkII
LmruGaHlZtWFFDWTQtAbSZDSSykVJiyHuYaI9a6pvNwnV5V16bg3Suvks8f6O2oB
gG60mZh/fte424KtSwhntlFgF8yTosgCb7ExiijQDVlZG1rsS2pIAKBkE4suhjUW
j6yVh8qHA4KJ+8i59aZ+FtHF16tY5E3ChdcP0QtfASWBreiRQwAiQsjE2vuAovKJ
OTFiGXhxr/JFvN/4qB3p2tugEz8goOqQQ6pdh05c/TPo5iOrl1O9pzf12fWGs/RH
C+zGVVffvTnZ3vI4zYriFEPNPkllsoznIAq3lndPeml+qR9VBlzbhvfjH/dbzIFs
RxDNgrKJETIpUfAAeGGgr7x7LVGkqjzxnGBDJWuBLukTNZAYe+TsjqZbUhe/gVyw
/GYLBqP6ljf3ucIVxlMt0vtgMk62gFZ3zPOADiItzPAu4MUmac6piJwkelpz2lqu
IRfu1xXNQv2LJZbfUiuKRgCY3KvBlnK9xjFZW13IPMLsEfgCaxplVvOjMMx/NDzC
va+4T+CT3EmUsqztHnt6UCpcKpmffV8Xjy0Ib3ShwfRQDXXFPnaNPcXcTEu91PnR
Shhm0xVzu4Bq/CDOEghdENRjrkx1vG9r1TtIHSRzOZyVWk3hAnRR3bp4MYxpXRHc
rW92xRyxBbzV3WZelQ5f3faJveUYW8BIZS3vn6WmfW7n4kNzWR2hTIYDAjVLTcCA
JnYdFAOeN3Nu5a2RueByBGjD+TPTZQClpz7t8YogGrMJi4qBabSAy1WpkO4zajUO
E0At82Kktxry8Som/8jSnLuS3ltjz93i46oUmvbPnawHJWe86cFhH+OBEuUMI6kC
cq4e0FIZP+kfjsP9th6tpu1bP7uu864M9PSmn62TlhDSNQRrtLkQXVNpminryUmM
dTNsMSmDQWLzrxF1R9JLOsWvKr1zT9GotkUU9VH62r1QcQ4G1KRb1YyOD3R3qPFY
8wnsU61ioWeQj2cb4QpUQyls82f5+kUaDBrf/1q9F7k8lsT510cbl9ryp5G53MrA
M2EVFnrTsPZDZTi/iq4FBhSeeq0UONK0qbFIK5fgf7PMD29lYaVVT9jocWOKXPO4
ACE3JX7t0dBmHwjKYYmrbpxNjrdFn65POMqjGuuMZAo1rQtG2u6rkaPktgJ81j2B
GemV5cAzpx+bLVHOXef2br/fdYwt7lKwquYHeulNMutss10JbKFpKcYSW7/KR27S
XXl1qLbXb+2z5C2MzOP7FQtwjM4triTBO6QlkNB4pUyHN+fCRByEBBsQzGQZQHbF
XLN0CTxLrjIt31kcktsVVVK3KfEryOb8NTOwSYjXJuJsg1Jo6gXvdzJOfxCSjOZG
s5Yr2rhvTEZihSCxuQPv5ZRgUawfaa0u5RWcVznsR6dvR++9Pm5qikgxgBBrUsgq
vtiZ9/zZ/6vCbwTUawVEfpTo2fQaZXKqZnyvbES4o8os+HoWYkTkH9gcn9AsY5Dw
4TQy9VmbdCLoGStIASUX9srf2Z8zQCle+wmxAyEPJTmyzPEOp3+P7fFR011R0h7i
5BGD5UUCC9OKtBH8waHv0BTOoJTfnok5ceu8UusRWW+8f57/KcgscvmeP8Mtlm4j
X4yWXLIhWA6JbadOIW/RY41I3zJpmkD4VNjm3hBTmPCvxVEpV6jn3mYJdD0PupbY
mSuSu5jBfOcIEalZKfBcF6ZmdyZ0iwONn0yeZ8hDXvn553A6C+toDAL7E4n29vgz
iW/pvT/dAVIWfyOaf9SHpmbJ4kTa8vjJb674vuQk8J/w9Q6w2suDitynaPJ6GixX
AJwdnDUB2R58CSVd+8am/ckMxQBHCeEdSFV9Dwzz7evI1oC8h9tDrj6mk4+xgUsn
vDDn1lL6FrVyp9elpYm2gBau+FB91elgLBHH/8sz7zj+axS1Sx9F7ulc664bKdbi
yk0FngjvI/mWWavPL5Jd2eWNyglc0i2Qn0795iLxQUQo7Bg6SrwzBKguAdFaBn/b
Yfy7Djne4GSO3bq4GyXfSqbi1Umhld9xvGlyZJBV9ST56dw1AK669PH1Z1vrA/qb
Cm16ThE635zQWGVFpPJhLkXslVu8P1FlYloQOEjkk7vM05iTAOObxCjqWPSmr81B
We/rQe/q1fMNtmItksYEY7/4SO1Q3pE2es6YaR0lil5vKx9dhsPJXlgBOBrI2U//
mWGEyqXRTijPqSv+KRf3gF/pvG6J3UasYfCfhr2JnVUJTaJ2N067Gsz1e2dIsgsu
fPRJDYI/PU3LNT5CKOlQs/zZ+d3WuFE62Psy9aYkr10yDEiD7JguPhcL8J2ALszs
msq6LwVGmv/uPY2F10Gr/cNqcpiYcCUzcOXMUPwpSPJashpyFvAEBTIlVKojgXez
sZcWf9UKBTloHagX62rYBG3uOUGOnLV6tD1jYk510SJgg5EPKicFXEk1XiHZruYi
fYXWOuITz83TY+BKjfMlmHVwbI5F9J9VQ+MeKjq3Xyct2+J2BK3NBRmna+Wm3Dx1
g69tnjavIcfkU8UVDTbqN6k4gW1xCEhp2nz+eg470SZopLx91JDBJtt35dHyKgLP
s49JjnuXyJr18EW/G8O6HynkANUrbMCTKTQS2/p+BQa5wFs1FU4AXr0N5fqxrHby
4gtbEaADC3lORl3vy+3oAhVwDDM1x4cRXM29shDWLwfJr8D69qghwtgvBBj1BISb
mXKg0GJ7soUnHmBi4mxyGZZVzVGcn6GMir2zmy2RF2C6ATHutKa98IEZsSJY1BKL
Jy6wqkJ82zamu5uWC1LZ2GnazgIQ/52WZ5EFMpVJqTdLKfyowo6wEFXJ5RvF6LF2
3QvLQnUlVXkzaXi0GP57/GzCeVxjSzcgiLDG3uPluCnZxA584nUNWqpcl1m9o4Xj
fKGAcStT7Cu15J9niaDUKmJurL+gZTYpKc//nd7XbAay3ZdGoDxKUPvSL5Mkq+MI
XylK4K4hm991tp/HJmf1FHkcD6YxOuyyrDrkT7kJN7xDty6o/2ja/TPMjOqL+kat
gmbgPBWGyO8qRofkGGvMmdMKmHz8XI4h+6GqLV/Lua/EF4fiG6oQbnmFHqDUHSoU
UaLOR9baK1ArUbzYZQChV2vjwsDjNKZcTtq96Q6ThmpQx7wCzdDrWAEWVAejna3X
/kUGiE2wD9Yueyj6si893rBHuxNVpNQ0SjZVy9jyijhmD4y//GWD/sm+qPeVeYP2
S+FkWVeyj+3CGSIj9c9ahMSfy31m2Q32EBt/7vu+N7VYhyTj1iKVlzy+CQGUjNXO
74EydXVuJ1C4vdsSasBpWyUrgCcDlxqCCSbhKx0+ZfCuK7K/BOAHlR6fYs3l+ogG
9hI7q3Gbj1Kv97V6DS1dlXubaP9Lw3DS9tcbupoDEYtgWI6qzW+TsrNJoI3YEb6r
yROv8+7mwlGbQYAvKSRpx9LRUlGufNbJRJr8mc2sRJEzKh3Hmnj3M3MA76aoPdNJ
QwN9AWmDP1F5QtsLWE51FwUsujw8HoMoPe7s/QFIGbP2cHukpbxQBRSNZ2GJk43v
IRdU6GzmsStrhpwQMuFSxBVlSdtvVFznaOW8doKPbMI6Z5KfmunpjnU2skLxGbxP
6QTPx72BkJ7r9YgWs8JhtWNJmnViyU8yOo2B2Q66FPqqmWFOvX7JDyp3LSHS2VAk
b8zJcaFU2wASJav0a5vdvdw9CoBe2L7Wed26259AHTj2hTPWbZMV7CPBhpmrJ7/A
hJ/Gk0V/Lpr/1ALkZn6Ho0GZzdd74vBw8rdcFielL2t8bjtSCCAVWDQlCg7DlyHF
113RnXU824tC9XS9Bjf1GoPG38eqagAFK2qOFCFykAalepMIPPtH2v+lI772kxoo
C3soMVCCRAIwZ5svxqXUCDwyIcrmf4wzvb3xtVXqWBK33xsJD1lz0DUH6aJJggH9
tQNsql+O/bF+Bx3bzaZiVnU8FYPyHyxFlGy2NHR+3WWMHdY4tP11bwTRTvxDm68D
US1jBhEeCxMOASrpCvfijqMOmPu3pnX+H/Rma1dVzoY8+N/xHdxCPS5EzAQIpmzl
3NwDcQ6lFEpOvIsBE8nxDlHCDb4HgX60Mgq1q3f7rCICLVZZK+YECgRfLDM6W8ip
r87M9cPnek1idurH0wlgyvn3apJqFtRg3X9V1rgNMCZc3CQx7VzR7cioXbll0U11
tjOp0j07xZZ9y6NJ3Kf7i9rSSWMX3lgElFVkeOG0lzfjW3U7+Sn3EMRH73/6nROd
ch3kIxh9/+xKoh2QSOfJV160HWlXYNlCmFK6dWIGCstz/ieO5Im97DT8Akzvsw5v
Fj/WGgB24GUy74LEGDtEBKXavRTxD50wDHUdk7GmdJTObhM5tiXE3AHzjq8VdDMw
lhLkmS13a+9cz6i33/0BlU3SzwEnAO378Ee0lDBFzJlDkLHtG6mLq15qz5Il/dov
Nxg6Ly5aI45lnUQSOXpziAmUZnDmEc2nloeJ1NHu96Nr/YUjZ/TY1G7mkzHzs3XI
o18ugF3ygYa/XuxB3SFKVv9RKmwGjIlByUIOywr33gHt6XpteaHThzwoAK4J5V60
8f+ZyMnQLjC7HDjNsmGjLSb9LJuNSVYfZ1hfLUw3HGXmuJz1yZgUhiYHVayT56hT
lkbSN987IWAVCz6pkErBbXwDE0tHCdnHTnFD7a1Poaf+JJIqCVrnQrMakV438Bx6
HW2L4NwWgpvO2rQIa480Ia1+CINVlGrrwZUkQphV/AQhzrmKH8vwq2TB/3ubetcX
O9j8p0J4IN1RTAksMp7mKZtqNlnhN93GSIqptveAMX7Hu/Fd9MrgUs0pg7HuOgf3
2elBFO4PAjFBPRKiyyArRhVVGQQsPLxrh1ZIqu/aGZCuZEOI6YSzxuMsqq6oAJHq
ISWZa6SWoRyKcpruUKkantBSEh0M2P4AENFVOfcvTRVGCoWsqiJlbohI3csHMUyg
g9aHsvFMdejJquNzeWNQz98RuqAYXFxTjt9cp3mE99Ji9nTlpNSD2d/27kNhezY1
7llTC1Q5AwJcWyxlNPEqehXE0Ch1zbEkbiSWUEU54rcgrmlFnd+Azz/u7G+8FEST
tsQq9E9cpleK4mjEM0nuCP0/8uzasuyjcdIcdlqj8MqS3FptHmIRIjIL2pYT6ll1
rk7N8RZjDZMWN59mJ0Yzcqz/WRtUks8jSPkN9ItlA31r+xSbI49UXcRlrAysMJAm
MBFa5hyav6DJCusJq9hMcgQc26H5HSx36/owqjLPAW7Aa6JCEM2ZVJXf1ek93Abh
2ZQgxNchgGibpKuPRJeq+yxudrSn7FX5AKvMQqVLIXQRHx3nEvXjB995C6yU00Wp
rnB2FYMmaqhV7knhEXVSXIab8NQ2+EAArAb61QC0SNgCZ1alnMIg89Mf8ZLO7qcy
SO4FqXV7i4iWR8DGpj537xfi8PsGnLLW9dD9rkGb982/ZckUjvC7Rf0RSrqgFJEY
uYvs3HTfjYcK+kS1NUoUl0afKGSbaiKbBX1ADozpXDxWKj3Gj9gowNFjUbmsxDRq
MFGlT1LLvJg/IxrCv+n2wxwR0flBJZ0F3ivTmo6GYenXnwkn5EUhkKS04uWkxnu/
LcCnBTRZ7aLTH4RNLtH3dk2YRqfKlDV1z/GG4bor2CNF9BbvFETbnaesdfbnuSYZ
B6YkFFLMOQk40piHyzJ8m1fn3LL6XtX+Y0PZzl8t4PIwSoq+nDz7gh63xfrxQLV3
a1WwRgfwenodhbDSDyDBIf29h8bBSbUBacPMpcStzH1mVWB5cNZtYVwaIgEohsc8
3KAGgvMzNJP3s0Mrm06iyJo4Pot8UVTp6ycmWYwg6mM6C2txK6wKZLNI7G1kW7hy
fXxDj3XrnE1eVjL7WIorYvkWrkzuZEyroV4wpKKqmGGl2TGGtYWeLQd7rK8Ie/J4
IbXisyHhBkLPBZACj17e/1G07N2XPiC0oprlUDQDBA25mkxr6hPMQFmNfBZsV9zc
yzR3MpueYYxF/vtGTrSrN3FuDHfX8e22BQGw7nltX+4jvjj0GigJWdIVHzYm9ohv
ryhLbrWHk8/fH6zYROueGPQhR74djtQAvYdk08zXNgyY5nmidCUBUEkAE+/nuSv6
uwpAxxznDx41HIKL6rWdtkRcKgbFrCPmZ96rxa1BJuLvDehBu2K2rgUkk8oHTofj
tTYNJwH/9tBEHzl8niVJQbril7G6VO1GbaRnKMR7Haa2otMNMeQ1YWGrMoquCI3i
E4McrhAxYSY8Dgs+wXdgGQTsBXzIdUn4+z8cgddRVIN9Ooeqdk5ROs4CI5FKB8/E
rCphdk3wuDbWzBBq5ZnLVL0vLuQ+mmjRIhZyHMaeqYWsR8lScRb30pdJVkHJqgrE
68CCFTaevG60cxnbDIMjhmiea8o68fegXBEu5zpHIjSimgrGeZOfHYtBsiKgIbQZ
gtCP1BF99VjU6PxxWznMn2KCATkh9X/tgZyX8vY1xT1wk45YeQjbsYm1W6UhR8ve
2IVAwRry0NahKwyEPXcchKFKuTFSWGFV8guhuKe6fRpec8Pz9qbUpFRx00jZTgW8
RHSQM7qPsjj4o0KpclvjuUAxgyPlT35kMa7GoOW1n23T70ttN20aBtBo+fUSnWVC
O62VwgeI//7MxCyVTZd/WyW3dxR/PU0BvgRQOKAOOhvGSJOFACiDtgOyKUkqHpi1
r9i+ASHVx4sCOtWmwVrVVTxM/ViXiuKoWH6/m3BO/1LtyWqcQ7ylKm9m8cXZ5ZU6
7mYKmRfn/kBgvsUiZAn7CzGMxyyRzgZtu9wXmJvPgyer7smCneTwswz/8n0oyDty
jO6j2nLQVACL4cjYlaz4Li3c401hr+GvbEuM+1Vf7BCqfMSD1oc3Ey4aDGRB++Ir
EHOnLVmU81HnWkTt3341snS42vFwB6RFBMGrH9yxQD9vpjpev4h/3RqVpaJ5ngyP
pjhoKE4pXkXB8T4OJntYWzZkRfREvj5l0pMiQYJhPVXeYmme+FqjHmIIAcToAXOQ
/j9qj8fLQHHLkiNz9GCMXC/fJqJSFcDFG49h0RoyjqNREgnCpO5YG2gqIlpoXj5w
TyEEPBeMUsByPqlTytWLjEG/6V20ChyT8zV4QFfbr9eTBbr5Asm4uMzUfm9slI0e
Xvr1mM4yeLHsRVl/q/6DJBgFcYnBPDeDhm7UmMcvCG3uPLUhmJ9Mp0l1ZruXc0hs
Q4snB/Q1pZYlabrBUCTupnNcvHMGy8UdfA1RwZOb8ycVklZeOv/AoXXAM1FcLjsF
SiL4wcCVvnG21WrCkxouzv3P+/CgEnRY7nOLO2GMAu0/anVYm9FcCDZ8qROGK5vs
LmkR9DL51zt7pW75mdIxqagw/ikphWdBYQLWyPZZEmsdSFXBpnrzBwW5hXA/O5kQ
IDdp1Wrh3Vdu6pSmcigJaChWS4Wkq3yCoiysfIRr/hqQaxdeBH5D8eeeDKKf9JlA
PKz1XHufNLIQrxha1jFWQny8uYDxW4yDK/4/1ZlLW7975JU9Ux43lPl7Qkhwyssp
wO2LogSwDwZ39adwNQ4+P/d86ehXq39GaJ0wFyVDz4HRBHgEa0+fyd7KIsGvZLVo
1iJNdIHlQVBz3qyXabpmYcD2sd5Pz/yrECLN7MyjVjFUIswUVsimcOLURvQnmiJ5
WVpYM6bJxFhdSalOCr2QwAcWh8REpQHZLYn+pU3LnX8fFl5DYGM7+6Som9JW6YTm
LG80M2mWmSstIVoxUhw61L7PXS4p7cDAvwN70F6szB8f3qs/JXzBYeyeIYaS8XDp
k/JRj9Vp5EDirdMuAoaLK5Qo7zP+A0lhsQ1g8TUhDM6Po7wwcoFv6u9p6eotfWoL
JlwdbgLZksy3zcF4NfEd+GqzRgsZm4ElRoL9IEqYdsskwQXnnZ6KLD+AtObnY+RD
LaqOythuaURUage8bIGll0wLyGpnYu/QzRNuFnWzy850KzjkLfkoyCO36b6QXIFN
qU90v7aQA5oOnfo9ZaBZ6oOi3/6FzsWLYJLleLUc/arxbY311P74ugncKAEf/pQs
U99ICqBWEToTeQxHduJtcPVxgKMpb2eajCRfXdGSCnEvHFQBFRNkTnG/NypSlfrF
jh9QSPYa8Dyh2c0B4LBt97kRveFW9VeDUdBSgVGP05834AzugoPgrjBwyXgLWaZb
s+xb3oAEP6m5w4Y55d+0Ar6mpkjRc8V4NjKUxCxDXuvvn9Mls3s947vBdLO3l4MI
USVt16Mu6TrCjWdnW1Vildm0H7LNT3QmhkNlDRFG6kyqSEMUMGMGLQMwrH7AxF+h
o2oC+V+0EnszyShK15FGeAepRConJREFwz5f74AQb4spgwhnJHh/Fv5HvFTHTR6M
ZelSjlW2Yh+vy/MdJ4iNt5COULow2L83p4B8xz7N6Bctk8HzBH1/hSeIJ76MzWYr
ucjGLxfms4MUvlO3SwSOjphclhGgbkVLxfxuP7/HXzytlmjajbUMpRfQ1M2yUbtp
9pciIHwDfiQW7Y07/J4DXBP6EYXMlyEqlco5TYvcLRO61twk2bu7x1ibXssmyQTJ
eOVC1Z99qgnjIkc1D1o9ojEIBlIWuUbpq6F+embSYszwGSdtkn+uNJx8AkMmbjMF
uhhMtAPBJX9lIOc0RX7iZuOvg/rDB1UleM0FGoeSrRd4XNneMvh4QoiVFKsRImIs
LQhbDQMpKxb+hy/0ZdlhgLXm/e8LtpI0vQWiw4n9wOLvCCn5FDogRMMp9GG/SOnI
jVrd6urGqxi1RZf+I7gTca5BTLH7jDwQBnZ/r8O0fXbyeByHzpVXimsA77NjCIeJ
u8P1+k9/gZvE+sFGBTGEnhYtxTZGSnjd/XQDfse9Zt0NA0TMlGbDJhLVxM8n9gFF
4QgBdP0j52T8l17Kue9OZAnXZoNxaUS+YpSkTE7z6MgvjxCgL+GfLfeRyiwwjvKN
XX/8FINBq+Hn7T3lAuWDh+0BpABjnKW64MLhFTG3UlSMMlxPIzPyvM5Hq1h1cuxL
LmdAIojWBd73gsyfAjt0e2zEYkZPkHxVikinb291I8TbVmzFXt3q1DWLHfkaJCTM
l2M0hhSG+yQM/tOBOdFmA+WhsTYyftYe7gf1SmOK5iVRDrbyKCn9W02zH8lqWodD
04GAXRR4Lp++xFkF9z0k2E1I7jYjUuncSa1vx76CROoSof9+9ddAm3XXiwdNmAmM
SAkIqgu+rSS9gelNTvI90PSm+bQu3jnYTBJtToosHcatOgGeMmI4IavIXXAuWhik
pVlWlF2EwNmYv0xBvJQ4smVzuCthfQCPfpE45qzWUas2ABCLe3qaGhzTz+A01BuW
uLwplbj1e4HAEjT6Bq8GYs3eoYqBmjpGNecLWgcvVWLhv+i+PcFAecBAewb3VO16
GFC+hH47hKe8HuHFHzQKVxn3so4IOpCLwgQOonGEcrLUTX0GuV49aFOATrfcly1q
cPmrSjIqZ8g3gn7unmnvD5POSekmAY8IO3Lgkno0ZN+JnLk8TZnK4rH9Hg4swkAz
ksOAWKf2e+eHAHeGjm46kSebsoaEUa605hQIqZDgqCavRj0irWadOdr1b0SZCY+/
alILO5a208KJqjn7YGLdNozMS69QN+LRRHBZbxhMZStSAQ3prYj/3V7whCgDi/ER
E4kxFa9k0ynvS93P19gm2UwYXkejPxCfX2kpSyhqj9Fyg6r78gzTMvF9SfeT4YMY
J06yY4moXIW+o7L9ivKM2R6iB5gsKHaW6vsKkMiXijJpAOtfXuttenKZq6A8hK3d
dx5+tghgerKSR5yVuMbYry39CATCLYItRqI3lctsFMnUD1J8ahvC4/a5ijWirFsB
U0Qj0VqntIdIJUrYQ9445cY9qGIlM7prXNkQJYLJoMx4Wf6MRH6fH/KRcfZcSYvm
aWU+GPrHX3zkXmnDHDhLnje7e02bLG2aLTtmRdZxGpE3aB7qMyBn3hz7xegKbky2
q/iMrBkWnkfDHL22/dHRZX2h3gl0vdYWe4uwAoaol1FodryQ+kSCCMZDuOZ1TK+c
nFTo16iaiGqhqx/EFsCch7qMeJwarg6IPT7tGSsZJxGX9NY0t6PhEJsJDF4UL0bF
ZZFyaW/xt6y6nwseiV08W5oYKDumPJERQue2k1PhVKe+LUXS/GkeTSa1T6lIKtzO
FC3Uv+mFJdEAyBXWTw2T6oAEQuv/oG+Rw0/Vmy7akIeXvzHWZJbGKYkC8YY7og4m
7oHK0IF9nxiCGLtvSNdEn8+xbqav7Q7cYLSo2+Zf7cFDOvzFVTVIfQLVXFmybP8u
0277AXPLxLCo3wxhxuxhNilL8JZQUSoV8DKAGpTbocaQ4TMGJWnEgZA/69Z3lCZp
Esr1bwAj+LR6SCqaQjQaKgfaO2eqDeCMTtm801mr6WfKxUou62xEBX2+w0OfMaRB
GdH/qiEEyi42lRN7PbS1dnjC7NvLuckEactJ4dYDtenm2xQIYRPSZFDBxEv/t7ds
9363j4vqZepV55btNg70xphd3L1gmlxw5vlULTqXKb1X1mI+JMH3SzAIXyKrRa9e
M3DD/lGelzWXsC6Z21oJQRvV1Umg2wPDvPuYIq1fOMmTBJqbOGvHWtj3/tDG0t0z
rRSTcPr6/2lNDPD48uXpOuOlWZJnkmKtnfO7Vs51QXoJeFeVpCjSTDWhImypmlLA
LUjM9QfBibTTlLqB3UzJImb1oN3yaW8aTqWfU2NFSLa/4Lyl9XlZM+w7ibj++TiV
rxL3P2rYdSWkh2/lm96NeZVPH86u4jr2b2Sk4kF9IftiSykbaeZalBFB4Vm4UkdK
4RuCgztq+zhpUVweRSBxrPSnDrcJPoKqGXfxYhmzMRKBsXJ1FeLLRAxI2+xyuZqI
r2ZyPc6Rl6BJuxnDKVoyHcTtATfTU+00eeooIen06rlH+KJ+aklErK0hvvPPf7xZ
24iIXl2i3j3Tz22E5A88oybQXbvJMCTJZyMvdyTtW1r8TGCOwcLIBgG9sLxQuzFk
58rktaAlo+PC1c1vmkXYg+zeltULXjt1s5ar98FEc0Ni2JonhGlQp/u5MqNUEnZA
WLLnrlQtCc1mWqX/0oamdGdRrZJVUhxJMdB3+eX20lB+Nd/4H8rElPOj0cdQAOJ/
WoeqpieriIBbbyaXR8Con/MSJf97cQY96Wbydyv2Lzt4qxUXG5wsT3i40G2BHvT6
goAYmUVIs4sLBVyWg3anhqGGzSq8Y5HMkYvcZ9k4Dp8jE2TPy6TzV8x9Zwh6CGmB
skwHP5nhZuLBSjNcn4LzklZ8afzZUY6/lUnyurfOjwmt6efhu5tyZPzvtUUJcZZj
5UI/Vk2SqNL1EAanuQ7ifipfuDmRjVjdG/bb+TT2/Nes1avdkH0jCImnN8FMa8x6
fAtuP9+vWpQaRcFSTT7rpja/+pSkFIcAKMKQzN6vJ32APqOS2Z0n1EkiGjAzf714
sY7DSH7FisrJeBlTmyv1keUt1HBziE0T5z9qIjHUNfMM9cNoBmDpnu2GXYmJI87G
3Z9ljEGbcECXOvEqDfReuASKsJXgHpbokBZs+Ln0aVt9GgfDhLiaIIUXGtQrnccG
buQgLjylfXEPJc82tcQXj82luhaF4g/txYba1wiwXTeKXM9TvZVMwF3OuIq49fdN
dy6in1Dw+KFIScRdHQYsoBleNyv/zQ780wTpVf/y7M99ShFkyMoI1CTvkwd6UbRt
cqLo9PJhI5iR7MdgpLZ6LgvPRgv9T9/iBXUtkxg5Q+NyFQAx3s8dCNSa41DyiFv9
ckmNvTbAgs3UKhSC8dsnnDU2h4B2UnGz7qmT1F5TxWqYDjBYaFkoEWll0huivNhd
+n/1SnIHlDGjW9KPZhnKAvXsyvvzGCuto/ye33oiKFXqoXmBkwj70HwGSj8Hc3gs
py48pTaGERTspJg32pZoNkWThQpcb1ialWByHAlm/fWQ1hk1fjWkFRBAdumxVskc
QqxtJb8F6qybQTE9eKkNbs4QLgtmnVMYw1aFhjR8rUIj4h91Vo8o+0p2C6+5IeW9
pD53aB1CFUUfT+yMP8nTsFiT9uV6QDTiG/8gwWEfLvTaq3v/s99xuPR/yr7eDn4q
cCOGhGJo9cHxVXkghPwr2OihHWeZJKIfFMxJzgfh10TV+/S+Sf3PYH/Wt6yn4GU1
3WKpyrjDoV4wtsAEXvVR7cgHuxWwW3hDxq/ECDlBHV46D4ZPJizainBMzYwoXAz6
6rwPaOSMkneGOLn9bLWEM4d7gc9kv9+iyWSYyahMifYRDIsI7dqgvxz4lILhgC/U
HKkZbsYavgG1O+5pFESDAneAZdIuUv7wrDUiKufGQgQaGmq3plNGjKnN599l4u4o
+kicj657vU3tLMv/kTCPfsOAHalE7GOgmTpx0A06oMZOLmwd08K6lV6d4d7aVlOm
eDFTrd6/xz3J4VZKPkdatFbnT4rtut9DIhCoom0TONbD5TO/tyKzgZ5thw16Hjg+
/VA/3CsmIwJA/0y/TbXweZbSdXfw86Qe5KKUDbztjBqrsKW4XANOFwtT6x1/UwQO
DhAsU+36WZAedyjjYoWqMfLo+rnAY+9hwDademm7ThXvcLLxziDtfhp0no2Sd3bK
uxA7h0HR29avKufLRO32VVd5fZeyvTYtWsMYUPUHCtyoOBSXOl8tvRKGRNouW6QZ
6vx5yLVMzR3/n2T4TFiTEvcmVQ154XQO9s7rTuxBJdbg+OjZytt9ZURqmhiyUUXh
xF1uK7DPh4YENqqmmzATLb/WTzPCPolxD9gcIOZoHUZZAf19Ic8/fHYxsdAVhGqB
NcxWjYiGEoaFtA8BkixDboltGBv8w4p3D9RfvN7hCqDcjq0rYuL951rWnrUx7yhC
C6zo/VufR80Qbu5aUv/gfBbsutgVaCQdwKQkgt/3LZfVSzXuZyPl2aiTUY+lSYXZ
MbHeavo+jjzQ0wzAXMv42P2U8p7sKaQNLMu3jcpfVOS4eTj/34jX39IESSSR9xqP
pHdzhPWRZwiqjUqGZvZy3C4IaytXLjxfPvrKUUaBr50mECDKLO7YNvbq5vI3nhSN
HSTIb1wUuu2kd2pPSBK2JBnML1N5LuDuWNRCH+3YXqYfQd5kFWdmFXYx2kk2emYY
rkhm3zgRsVmMoZpqA0MIoiw0mYBEru41IsLLhLzrXndcAhfwGH+KMrxBMnj95EX+
Uf0eQLJ5zFp4kbpenIZYdKKmJOHBbP+4ZZRbOGxu8kJjIfENxqz/XpzsWYjWpZBf
Ice/0nl5qRAAqudl9MqWl8c4nkfr9xZQyjMKQPti9AR0tgGDE9/39w2tICaJtTHb
6BDmJN3A7UXC4VVTXNjVOGtdEDWbtStGVPfE8jOyTeblU17pH/yuX2ZZNwRSrxcC
AoCgElbCVsSiitAY8B6wEo+/Al/PY3LDh7uNFtSFP/1VFYQXQXwgBtkAOudSvARK
rFpsOo8BA5UdXYen7sh0qUYoYZI/FH/6PtTXhiza+zTmdsWpMUagZHGeepLKxYhB
xz0jYGvmme/UUpjPFxp1DpMQiPXppRLIu4Pa4CNr3dY6LhkjYXoK5BjsLuG5SEep
8vO2ab72iIdLwoZcxMPD5LZFy0cSUpYIc4OCN41AObKA8zkHtOM6qmXaPOSK8l9e
g2J8dJBpDcCRoxamiRk/ONeyaTPx42NJDR7mMsZ9tCtMI4Ij8aB6nvP67vkGGSVw
zkp8AwMxzgQklkN4zR95tz8fHLKKuBjz/s89yZx5fs3z6vVB1K7o2hy/l7RGxAEU
cyO27khqAtouh2m2jKEd+qV4u+XPVZGlpPhvu1fdz7ZT8UX0nK2hiAx1mzP7DaL8
YAkBWu71ZQuMRRDitisWIwuFc9uREEkyP3aeOPWLs8IjZA40+oNYNq9MEUKwrZ/n
ICb0SCFDoF7+jCp/EPEHsrt14DLHKJ+H5P1OxVFj3Sess+1C2/SKjnoS1k2lATbs
yEXJpybuOyRYYbj/rZ8BMAowiHtyPrXNUrbA/pxOnPlToID2hH1VMGDNUmIEuIiS
g6WM3YEBxzQqJ5ii6ee0CiG3CDaG8PcHhZuHESqJW0QujldnU/L7vNr3qcDsO4HK
iumLMev9U3KFvHddlT5+X/rULJTG8CyohmJ8U9z9bKdrQdetvZ15psKflynC8Q35
hXLZtIp1ou3wlWxFc7/j4l72+4jsZICwz13GezIYbrepsYCc0c4ID2vxYi/+3HhY
L0CeqriQhbHBnNVK1fKf33kq/2y0blkxtbUhNRAhiCy9RVevAjVMt8waOgzfeDsB
M0t1VI0a04A4r2mrJbkVRbDSWT7JVo+MgrNPJKNrOONKCrWhHZmrB3wPa0QkxJnE
otnS8OXQ7brXF5Ia7x359N2opyEizbjWArup8hPbVoUydppAm2UPl4ySLnJ6TJ7z
Zy/ojfpAFoyAfPBMcgobwWSwsr9TrJWfA1orZeFQMIMoYMVoVhd7HWH2pzUcrXzp
ECZFLKHMG0m3XQDZdvklevwI287GxLE7EMKr26yk1AbjMfPPT4ts9e4Fexa8gLtI
10C5qrjkqUon8PShkA8EB9XzbXaIuIALKpEuQDyW0l4xI88cHZ8yyThcQatyiBSg
HabffJu3btSpKwkNhDRAWgSW4d5rJSH8x7+FDg4zIX+YCn05BWwdtbuiYX0KZ6Uo
L2Ecub3VHt3FECxQScDeVuUYXAs/AK58Gx+tVLdfP0FPiES7wWqnqy89WkGB43GU
s1+iH4Tfrcq+tvA8LKItNspbh5XWXVhWzGpdeUUlBC50Ic+Hwn9YKW8g34MvmqSO
8hTQ3qXBxmVvrZUzNUn8Qrk4Zk3LVdg91i7WS1pkkIC/rcauJR/adFv4nKnxH8Ui
WKSb5ZNdv/yJL8Xx63+jGAqi/u5vOVjnnwvsNGQmSFbjuTCyEIE0fTa6aPs1hag3
0iHe/njtRaUDJhkJuT7IeGqwJ4TA791XN4j3gHkY7yqqrb5pmtsOPCZ6KxKVf49p
kn8GI132J07Y5Ld3YeL+OgaBWwYrvUE5igUqwrfcfd7bHYpdKfK5jpValcZhkhtx
cWKnH5O8sFmu1ffQrGX5wwqQLW8e/NAfLpKX0IoA3MKR0MKrrriigg9b2dmgoZYJ
FoCUUId4Znv7V/5iYI1UPzaS5c9cyj0xwz0Nx+9vLyIHYOg1196TjYGEIUbo6FHL
kSutReUG4RGDgU7bFOxalPmmtk1pL6YJ2neI3zt6L+54HVTH3R+QcnUCZn8bKcyJ
VZr/nCFfwMuVMQafg3JH+VqYpYNYxuSpX5Jig0g7g2xNYIR3yihfbF3eu3nxZ5wV
4hZ8VG4dsZjame1Uo6SSJCQmTs/aAtHiG9Qj+NCjEsSSp5fMZJCMByTowo31Ih4/
4gXEtymaALlmokN+tjodqsmiXDCQdPkAMtNPy0cYUsfgD+lCrjCRp/188pYJDLfz
RLw+QyFQw31nSKUYa9LAVgs5KpsPf5CNwnfxjb4G1LhvGRudxfJPqTdnG1omnMtO
/p5L+3dzBsW1sdcUT8QT09WhF7pvgTr8sCOROkRWveCbCe5i0VfmqXTB5Z1LP62x
K3qC2bfiUhR+yiP6nIa68ynopRDm7bhW7GAjFgVw9I/6ear/ynY95QMyPwg3zSTQ
KDUFEN9g4xeoByyPPRoyNaiMfVFCFZfc7RCJ2YFy3BwRVHIs5yxaGXd3wiowHlvE
g3nelpYyPemYLwwCXDRjNiieee3NoWNQfZcsxLNRD1vx0nx2TeO99CPd8ukPaJbk
o5U8MJ85U43RWWWgYqk7PiBCx0pKDJswBJTdJZe18FC4YrWccZ03SkVl7K4tTqjx
xGOYrDzHNvp309DRE+ZygwIZeCcr5DFqjYxeuxbb6X4smv5yfpnRmMuILy7zYytB
g1Tcurg06ITmodyPQaVNubeRQHweD3pHYlKcvaNPNunHoiqpMOPtXIedBDGgq1Dn
busZobCZ/Fnx7P8lZHeH9PSvgVGlVNRqCSg25tiHgvAE9nAOjNoWGCov6br1WI0x
7rXdzPq0B8Syytf1/wByef4LOb+F/7bzWzfiQ4uHQB5p+K6VovLK2pzX6uV50qgR
qLkkHKJngrLrGyR2MKQV/PU95N6/QL02nhc/Sdm1BdHzb5yQYVxLFuErFOfDkR/O
zHPswKe2J+fcgwG68opXAlNRUd8yh8wCdEHvMUEisM0Lm0Z5+tQDzgS9eQmSTH6B
bbrPu2CvyMiGpifRa/JnbNIeyqVMvMuaFKU3Zuy+6mCDbjEZrjsgogaQvuSoOmca
zTtGC06WFE4gHePDTouio07nooSclsx1AwJxsstBPqVuGh6f4S+BIjdsZsSPoM04
QuVGTqJ7p3MbEcybWLu+YGCFrk3MXrvwYpX+3bWojao3cyWRS8kRN3591ib0EY1i
GpmGM0nlL9durkvwiXnV+DpeOT8AwRV0H23n8mFHfViAWdGzAr+GpkSoJVHtRpMi
Xi52asOekjiUAb4i8aZRASgkQ8ObVnAaI2g4TUA1jVDtl7lw81hKzLl23Kuozgsv
s4yyvPPoRqgum61vBjGwg6KFpL9beMBxG4d3qBi8l2YYVGPzobmFpNCPpXmXPnTV
YZUCSV18fVJbMt8qdgm6ufQCW0XBdgQALpWINj2MiqhGkuAJPxoZhhhqopvsfOCD
cCFZg4uzoJ0WuMGrD4YIOljI8UkWmt8kA6wvNp1uGpWm+T1ITnT4C3Tn8uLRpgcK
arSjcJOkDEa3G5Z6JFO1ADQPCOTdwJehpPhL2E2p8LFpQ0rIlTYu0vXb6WN3WpUd
kxc61TreVFiQT1f8eY1rqYb/gGt1jaN5LY3ZHdO4KCt6PlJ2XvHlhZI7HA/p6E5v
MS0e60590un/90DR002+O/e6lkOBv7iPq2Skflit8hmJ3wDPCyfHvCAomYSrPhrb
KLN69NKYrYKL5uvJZFbtVuvD5Wh3NwRgHjMmzfBs1r2Hc2MSlARWh4wTkrL8k8Io
qg8kDJqQkf7hSnCgLNLUfvvDa8bu5RmrkUHhLFsWJKogmHFbFxmU5+Wjh2xIMjWI
uaH71NLQpoILOnmG4r5n/Nju892vHa7juTpYjlOxhsOzPC8/kuH9nyhQTpoGkgNa
5PvvLDDvuA96Q9dqgJ4pwRgYB4u+Mmbsgecf2rnoyT0hC+5rdPnitLkiDwMbSKwl
Od7pyHJUSXX8nye5KZ7fObKrQ6yD9+rfRUqlGtAnQlUptDdYBNbZdxWDoV5yBAhr
ZCWIDvgEgYTBBtER6vMJVB4rEZnCODZr03FXso2C4sApkMwwJbU88XBbmcDBpOQR
MYlFq8No3paBe36pGI7F/aYRJ4FQVYPKfMAsH3pwLFWWGpxiBZCJKiUIAqQ1x3dN
NsG7wY0RvylTwaPbqzFP0BL2I48t5Cy+ShVE/iBwww4Qi6CMa3R02cC/Eu3t6s3p
BvwsSBoFzYwIv+YeC/m3w+avbP8eViXNkA41XxinGKDSX5aPmJrvAe6xL4/EIfTB
NVaI7ZTcesDRsMQx2QSlWQ1DVBuOUCiOS5MbdIrevdLZdPxYMpjqfkHTmn/8bHZs
5ZmgQk0/aBOBRgNNLxhz0yHHO6xSNP8Op2AEDxfSrJ+8z52XM6SxEQetPLg4wpBL
Z5wvaXjxSMkf0eVSPQZQvj3Nyye9dfx+hc6q0HEGVlntFkm8E+F4sVKtUYpNOw8U
Bd/FvJkgwenvba23XassQD9iKB5IzgJy03a5DEDO7g9zePohLEpt6dO0XLZNxjCx
aJ40EJL8Ghzdsbja4wmtKopTzIUA2jaAqEY3g+J2Hg2B72y21q8LO3c9f3q9rIQo
FjDACsY8n/2Qd0IG2ILj/UwLaCw+Z43K+3Oo6wO8p8JxoB3dfYRDoRyGePEj+39t
v8Q7n14F+hO95gngo5ivR8ubJtEUb6O0lKHmZkqfoeLJ8NrQ8ZhM1MG7Amzt0plC
llYoYqK7/rL03JTqW8DeVaZkJKIRxCRdkUkbamubEXJJgnvmHS84TNl1+P1t27Ty
vGXyHTiGmM0RQI6zkz+9W9P6Gs1yuSgqdKk0jsgYBcNcQNMKJIXaHna1SDzhQFO0
/bqD4mmUwPj1HqRpKrcDc0+HeEp/9+yjvBBMqVIIOcDZvJyi1UIvlx6QK/5S3+qs
usWvPbboV3xlJENR+KJl6KYYLJHxxny3S0uJzhvo4OMQ6c5cTr2L/RGvUVZhPfZB
0tuSxCNNUC1/rVt0jDtJDy85LHHI44Ri3bUnLEAxDHURiCc5LMWQIxipou0TTfFE
NatHMqg5bASG+X2c0xj+he7UShH84Tj53nPGQdz7sipuFmIgbGc/nP7pB4f0Jktz
7QZWmTu3U7FUNtNDZt+PjBEAPt+UMnkf49vrG+gNydoX7sbiTK2Ik/tlIuUkfFxN
219mnVwhMXDJgnVbQIhsHjFNZcKfGvlX7WCBWUFGlQRzWimdNDbvMl0ULM5mqmmy
6xGRsF3wCdqwNX/CH100QM9gqdpHNOsmDnK6dK4LbHDl3KFQlDI2iSSRBxo8dN7T
5+vQ6LQ9xO1JPc4owDjLFk/y9lIlbD//PvhWp9aaquRhP2xDZGOQwrQSf9S1HkBr
9FwItXaa3n0+KjlmH/DllzcMQF1Wu682oEtiYbl9soK5nY4S5oNjJBP8PN00BvQO
UEBaoJiZ+XfvqKvht/4839z2+qqv+Q/Yhew6arGrvUL59VSXLRTA4Xhz9I7Qu8FC
8Xjv0iRLmF7KoZ5mng27d4BEyDCPmtQDJHdUjm+vAp6LarS9Ud5AsRIqce95K9Wn
ZmkKirTYn2NciyDcvx91SYLWcy61eC9L9JOuAF341mj7qnvjtuO+X5BSI3cvoAi1
9Cvqs77MPfbs5nAITJbxAJx0dNckQYuYGAtk+zUvLMOpO8dfdmZWcCfrmbaUT2Xp
1o6R1ArdM73So4uKHqnVHwX/BFQaZOEEEGSw4Ge4hdxzJ9ubCzbFeuwo2gb0w/rt
n1CJp39AJMzFdX2xFjk/K2Qm0dF6xAptZt3eSg42fqM8VWFKm9bMi7uJPvqi0JLv
F3jXLhEmDzpAYxkRYwU9S0VS/QmhWRPQquHXmAFm+Oqg53HYLep+BqlnDqclf84S
YMmfhfIWXhEiB7NZ4OnNptmVLLXiXtXhuJE40Wt+CFJlY2kQ3XtQLPfl5RNHr/yQ
NMsRfDc2+8DGH+WPnnEP6IFF/MxGEAAdepZeKpy090C7ZVTqQKUrdJi1QIcoSU4P
cN/VaI56VWup+jHUJMHQDO+3dN+XsBblsN8PI0DHfIpecpGZzdBqm0yIYR8Ld9ej
h8JsuUXD1Xfov77sJ3jRkgdtbGp2dwx0P4ekvJPUEfqBTNfqftgGBwfx6rHfV5n0
4ttoGI04A8dcujsZwOurG55Hdm/V8cCrUQIb6+u1IyBjPWnyt9MH1avsLsA2S18+
Trd0/zAMx63UhA+38myTXTXmCHL8opIP7EqSSvvg7YXNpsWuKg9N1MXSWrttFxNs
eyhuIeY1L94dfdWGfEW9L19q42kiBI8m31YmSLqoLf2lixdBjagvLkGqx8AEq8Ln
XUo2cT3xlgg1uhjSJ38BBhObEs1btTZEUyxX6LUPQWKe5Q7n3HX8S10a7kZBEqTU
X7fQXMQeTsdCPobWUj0JxXyfiIAc0BbQwwyGvaXkVHopqSZfiCul4oumVjsQHQ7m
GTRZCIUYQsT7gh5RJq4mtvE4uTyIe8kdiPBn7bzJfxLFbAqrXL41Kc2jcQWJ/aY0
61AtWhKLzUJoVTuKisvrtS93jZntarYprY9yzJ7NySBGZqmFv8JAZTTm6k1dUp5v
Lz7Sh3xHQbP7m8BlLDf8XH4yH2bFe9KTxqwfiiiWRgccCFuBH315eoVRRhmyc01a
rVX/1RvxWOudc9GzhhAeSgbD1vuzp8gAd8a7WlF15J4DlqaNzb9iDsSV/Seo7iKP
9SBphyfGowwCuCPf0VTmuiWW/U5joEy9MYwAgVuBEJxfRc4URiovavZTiMZo/wQi
ZPb2SFcpFhGP2Nef5xjt1mLfAVbN9lmJA8zYA+6pq1UXxvrp1f2XTyRTjPQgSB74
95+JZ/MiNn5HO+gT9kSHDkjKw2y0w0k7IWV8De7lS9bsHSR2Gaxp0EBtjDX6sjvg
B3+o1ClYm8asiIsiRL9LEzapUb3SQQkcTviZz1YFnDa3ejXHUnWp356j5gnYvmg0
C0tsVVmfp0iLePY277gywGgvVfqUOfSuzai6Oud4dIdVvI38NZ9TBfaDsmZc4zQq
oU++rn6WkzlFAekkQbpwE97BRRkMdS1f4arHy98q5HHPXvgnbxrQnjsqe40lFd8z
+iP+hSqBlkKbBHIQdT89kMdR1qGMb+tXJkalzE/DUqDAT0+EroHX70hbpy0u4tXh
jrDuzLDTqO4f5Fofd8ScwngbcXxRCCwQxbeW0ZEzwnFdeLJ2XjhYFvXPpVCDA8x7
pNnjnL6h3rqCtfRYAllkdgBLzqlX+68qt+kGyeO+cFN3FIPvEo7vo//rLpTO2Z2u
VqMjC2Kl2mCPg/ornBWImCYivRfgPPYXXsku/kGIjFLTduJ3qDuhsLDiEt1R1lXl
wo96ZR6ZLCoWZA5J17luXxWLa2dGw+akCvh6ItKivHI+jRbzJ7VXNTiujTglLYGK
GG6nNPuLEh2oFOqzFMH969i8u0oN0Unj/12bEejhnpgVA71kbC7husdRydlmy/qK
LTDjm7C8X0c8H2zqZZ9NG3ej6ch0EKVwUc2Q5FxD/g7E/Yss8Df2QtjvsJ5zzJE8
tpBFQyh6j2a2IqMPgR2hpnrW9c9XqsGTIukYUH2dAyvi9fS3NRedRhIAlE++HRSw
CwFUW1+IL+x7exKVFJYqZh4/ePqHItLXWqPhmyZ/1IuPTQk0MePKo2ydfjCBTc4r
2TWa7U/DNHjpSkPzUJO9tE6Da4qoG92At/bmqcWVao1+9rjiAMKuor3mkOIbFAVU
eARKC7MTjc9k1yhdF38l8cTm9An5Cz9xudISiCf6OJzNU7BUV711++6D2wq6ONc5
a+btjSFwhyjjanh0NES8/ImJBmLEFj/mwZ/ZVxsDn50Q8w9eEn/umKxyMsDJfEnA
9W7fQuSpmopbVN8Mw07fF72YXj9CMcBar5kcJebGFv2KIVQ5Bo+gXAq8tnPHk1lZ
ZfV3zKzC80+aE0AFg8ebLrOYt5QyTYQO3aUI/E6EmWIEKTKUFJtrKyQiQRx4S7xX
/uf6DexEavNT/ghL8JZolVYnnWqdd8zL5TdKXFBGxYCFb2HScB7HirqndOlRsTN1
SC4Y+WrpT7VGBjQSpIxWKkLx6Nsc+Mrha1mR6hXLXQbmW56ZOm6OrjwmZI0OhLBa
NcSkhZ9vUiQVEJBN6Ehhv0Plpm9kZm/b6PsABad3gV/GIKxl575oExaDUq6KGVZi
W/RGN+7pVya8ms/8J+9R8AXMetmkDcmRxgBbesCHSagxtbdrdlJAHR29By4lk3aY
+twhnHXXgrEPhbHmEogQXV/hnBWTYfCuy4cZZfrrpm8C2kJZEasSHT1Ssfa+K00M
4hydPB+AhgkE2yX7O7vKbQA0UXmSreT0daW0AiXZ6Z5puX0A7TKkrWPeOyiONdx6
F2LTtzGZ4uLL2oqBXdkcGRTicheuArQtsjiMxr1gADjIar6VPXAuDjwUUaOTqq4S
PY3ZYtGjlQhECZ8F0TYHz1cjsk2S5ot+f6sE8ywwNDh6c3mKnZd3W+pybQOz2bA+
5YqHeRsehB1a5OReXI2kmczmQWYVJ29yr7AYIRXHpVViV5k9WCFMjPjQkqTDc8Aw
BTXxnBlmSSZ69XHp5ovlgJxVOVOWQXChYmHPp3wia3g3ho3GpwdIuEgrTboftHBq
sGc0CRhk2MyDYQBFAW7vIRK2qUv8P1hDniOp0dEaMYtkVl9VgQDhPrPTbN0SDRtq
TV5Q2CdeQ3y3T8YyDZHcwxHgh+fp875gcZymZo2vW8PG9snkMKFYhbl+1/96GSJN
gjlV8yp/hszj27JSguZVyJg2xeBsWtkMfZQJsXaUTbNz+knh/Y9Q+Ndl/H5bZmKL
Ry+vEnQB8/ZL155CGJdGFU8A+zR/ZMrpIAxw14cwuqidsHUBk6E5CH5molaB3Qon
zGldiajJMAwCkdK9tXAfLQXxqUbh1Yycc67/DW5DrzWVKFeV4hvsN4dIe3J+l+Tq
IuU+tloaG1CZqPmq2dYhn99/jVR+CxBGKFCgR+IuND4piI8Ylde4eKzD4ysGJqYj
XMVjFkui4saGs0u4MnvJiYDw1ppSfGORl9EoRx7L+AYMMrvnOXkOtHlBIQ8qvzfm
378gNFBWkzjM+4tKatoOgBnLY25Hz81q5YXzIddIpqr8zA5wW8LgLJRDgCSQbYFb
OaoO2twexYTLZrAaobaA46VLDJ3RUICkjYuunXJpfZcvsE06sgpUvsOnob3KBLgz
j3AGEe01Q9/v6/cf48TaxVKTLsLq4TQYKi65Sx67tpbOJWhrRf+xAxaJlIB8iW7U
tA06ZqiCqkkEIr1aWrEgjGKh3c8OPVysnNa//lf3iaw0RN8sWKuq5i9S5IRd+yll
PVBn3i476j4BqLCC1onZHWctk70pv/AzQbP9/WDDsLvME73TLmzzBhXG1l3GQFKD
eSy6d4Vnk69+9M0piIqYKLcnH5PRy6evG0Km9VwraUf4I/muhPh0yHYOfJGqnoSe
ekEaeQuak3VgbobNtFJUNEST+RN6w08DzgiMSe3PMlvaXn9CQcia1dLtcsWS95rY
hj9/XmoLdgozWT79iUGxGVCOe1H0Ph7fqzjSrYpxeNQbnnv3yBuWHJggUXezdQ+I
l6JpDjCXZu60EQQakiMnWKDB78R9Vgif9ho6An8Stnq7SIZnKy5ulGNHdWe3EPr7
Dy5Pqd6KD6g/aNT7BkP6rfilN2xJKpjywAl/2mK7x5IFXgLlrxUbaHFy3R2kzkVs
nvWc9/WRxXfIDv3pxrK/Z1z/f8dgS2c7gfVPXpqo/vxnO+pB8Q3GIcjM47XrJ29B
xg/AEt/sX8ilieg/TQlyKeKl5Fm5+ckPBTfxhJ/3XXW12QV90T9035vSaDDVA0/f
1toA4xHNMBTNXB4MfeNHcuRme1GDpVl/TcUArxmkSBYJ5YbtVAeUYbzdQac6eA48
5/bEedETDJgnx8SdZ89Eof3gJ8WCUT4W3sBdr93BjtPtftdbldebeUscSQKA7PLf
AKM6YrHhuwDRVwYrPlr8BHKY3G6VZ121Yb2Le55JYNoZqilD/SPoHrugGpyRNG0u
zd1JOUJORufrrLByahWSh6VkJcv0lS0BKECLkB7gxGAhO4HDSWVKVUu/hz2EzoUx
zmjLdMloIxfMi/6GoSsiSJd1VgUv5lZsQF50o1jmP3F/ARYygbFEdsl9K2GmL64r
u2tU/cs0xYWL6dvVp/bBTz4Bf3Z0fuXVYLtYEJ/BT4QMfOK9/LTeDfpQN3G9BUKf
0aIHwTmXeWntJN06pA/cttFvqoL9AM+CEAe9Ud8/GKQuG/8nMIOOcSS3VXZoIw0I
yELeJajCv7a//SsntjPJqq1KQSSrAgldnDLdcyvjTdrLVE2gGLcfBgJF3Pjn1MoG
flIa2RHM3BuOfCilHwFuST+pVSyab2TUFnVvjNMKTyf+4G1ykJc3zMO2T4vDLkXI
l8FdnI45JRVQa0i6JLSPNt2g1dNsyUEYek93wMhdWZcnUN1rZAvkrxzOFsTyJ6Gk
Twe55ECiB/KajUI0E7BI28Zch9nGma5A4areMoyDZnsjXz9BY6rr1j/05xJEtdnh
z0NZSMfckl5go8uxPc89fmRRNjRmCfx9LZ0ro6IJb4/tPUo2Ds8veT10CeLUm8HB
uLaIGYsDf/zAwSdOimF5AeU4ayqSIjhSbQhXpqa6nvcaDhBSd4JGKbYWHum30zQ2
ESr+oQ2RSHI9e/Yg7ifbgsjU1EwLnzEEnhDOBn2MZL7mrm54x6GLOUGJ0q79qA8Q
y4l9w17eZv37xzkO9B01V7uA5N1/FZplahS0l9X27cj9sVPSFdW8DgGoAxPPUbcM
18tZKhVFiygfsE/dYQ3pM8+g927sCwhOcVYrp28iXWAIcgxdMDvIQZD8HtnsJi5b
vFyy/2OMgr6gdQBsD2+I6+k5nqE8REFNyDiwEYpJItMtMCkf7W+marhKAjftMZZV
3sEZNL9IWuCJAMErpQbl4TEY0MUCagXZ6Kyqx3lxEt7D8GJS5ZVj7Ng9kVfk8hLw
cwvwhec/Uf1cZGonGsVjnap6MH83biSMIJYo6+CxvZT/j+/WOzN71EX+w6MkBMhZ
FMx1wq1HYQkTweQq2Nf74s4Vxlt8rIQObsJHIjfH1W7O/Rbrcy1PiRdxyBAAkNxx
+7CvRFY2yq6SzVuTCeYyVlUhIVOxdBJCJkYXhy940W8p4czpFLWsVWgBlzDqYlAX
T+UdUUk0IvPtq/IhiH3hoCk5uO5NMx9ItilNSuSIlKgB0wnF9e3R/gtgeGtxfRcj
po751Z4I8xnQhWY8kIyQVKRP7+rih/c7RBIYPhGxa+DUJ0bzyLqaK/G4V/NnRGpL
4TDU3tZE+xQX/9b9GzDI2L+qmc/oVrgP6junzS4EDyBmoNLS+QTK9DejJubHMUh+
tvzCnzOOkQIef9HD1zyur911gV2SZqbmsX2La0WnQgySgYtkjXuUzsEP1Z0F6HYN
QTB68dMVHFO4BHQajNx1ZJ4g7QHQQtlOVbsklkDiNNAN5yWXs3AB5WgMbotP2kUe
ie4g/NapymKqcvC99GprJVtCYmCym3pq5LET6thNaABjNqMbWeUsvf4rGHwGOjds
CEOPVTOWjz5XXhwRUQz787de3R2RX8bps0rTWeuAH/Ftt5IVaxDkSZb+t1ga1Pl+
fJHnx1Fzn/4caY0sQnSg8c07IUBSN4mfXDpj/34E4+JBXwkX6D3x+LGptaKNHrEg
cTk/tk0bs/irya3xHz2AYw8g2xQFVWxHdR7/36OBkiba4aJ27wT6Czv79c7AUBIY
2BozZUTLv8OZ85Yv60Uj+3/A67OLMtVdjKUxs3+VBAFzYSdVODzklQjqIbjk6uYf
1BXJnMY3LrZ8l1t/+pdDxuw1/jNYIyk1tv7wIX1RTKA9I9vIiEoR36tkHVIn25tq
9mqMU0U/XzjTf6mLyki9ZufMtyUBilmNQnpMZsA+kKsGTf7ywwMEEBaVcAne3Q7/
ja+zL9rt7FtuXM/v5gPSEwTFMKvL3gh6T+/BqIeswDScp9n8Q4Kmdocu0ZZLqCrH
/jjLzFc59vgYQ/SMrfHF9fMaZsuXhhKDu1efF6qpG7QB6C76cQmjQCzJUFx+fWLi
rRaCAqBDhQqszhTDbrXQtMULjOCHagJML6l8uTL8I17u1G6fiu2TpXkHvXpPTiQO
Do3M6rAEoUzOiP7371izArFmw2SGtnpgbTAz+vnUOzvV+/8ExS3U60WR0gVnt5kH
u18ZKnOh/A7shKfSygN3cU/uMqLrAy+7XrotDn4vx92Ejg1pE0DkzX+Ln3iJYSlH
skoXuw0/L45qBYhZ1UXzV0tBISWpmG8x/DM5tDxpE6TX1HKt+EBYfi8IwNQD/WDC
OWq6+YWYtfuVXmhvkcZzBUz/DGWA8lPkJL8VW6GE3QXUBmsKzfo7sj5yGFlcpKuZ
k3mE+MqwJPNT4+a4FMp2iRZUvabLa5MeNVMzcB1T9m0SwqGKsYrSgWu7fqsJ+DSb
2qOPJBOV8w4DZIbPC+4b8XEMl1SXc/dy3r80aZVrY4IdenBJSensSVE9C2rBdgnV
JcGBGyLI+OZmJxLYsrdpj1TUJpqVovW/Jtx2WfkDypdDhZOXhWt2IUkB2a2k+BC8
LJNM1/vM9qg2UfydHrcLDII6g07tL0ZLz9RQTDiQSA2sRc+r8x1kPirdUPXuyUNp
XLxNMw/k9IDga3cyPv26eRf89ehsE650BsQfPt8r/VMfGCuscrsZSZRnR4gpWv+f
pPTARyeZfScS6BtQ50rtAbD6H+GzTBqefpVaoskCShms2nhrsJu8k1Gl52GV6wA9
ZPJvClePQ8kGzAQBdIZi8Q9iEdxt7IRHb21cZTvlqRI3kkG8Rnq2SdybLy8FWv3b
1fewLmUX/PHG3zZdyYoMFbXlzSNphQISS5VoXDqvo1ZABhaxNMKKwtk4lUNQuVjD
MACgJqbZDJNVwZmtG37M4YetAob3yYoxmOqQ/cyCJ5oZ00a7GTfd83va9oJF/R4O
OXw5j83Rckntz61XLSCmZTFpuiF5fFVVjTrthsDrwYarK+144F3Eaw7j/N7ZYQRt
umewIy8XifT7JwZzm8N1j/hnOFNvp4nl53Vz0KSOEbxwYGU1D8E8zf6SW6aWoPZU
2KjSgFsGGnU6E6DOi0we5AOspjCys44VkhD3oH1vNtOjy33griIIbd4EJ3aNKhyY
kJUaFMtx9hBMopyX0U9KRmeUDfcUwiGVqN/Np6cVAVuaPxf8EgFadoTi7IjfGpBd
ieas6QhmEo78gPzUO99G8V/T4dck5SIcaEs4JgEhFzda8Bg9kdw/u6x08mZBnvPG
DFY1UDbTPj2Nxl1mXBfri7yvHaoePnwnHbt+BsYA96JaDF9etBIAAVdqtdgonAn6
wknNFdpw12FmhlXlLLuo794VBD+agluRsfq7HmEf/rjdLa8qnnPKKzR/HSUanwCx
eOvEcLlcIs0WmHAdj/ZqUjs3OIvTlXZouJDPFssfCJbxxgnWdtqw1Vm0MfLJMA+D
nRe4OAfOQkARb1+kU+ledQ6cn8lGiME5UUKv6+tyLjMnLzln+fWpwA3jgg7EImm3
+FdAWtWT19nFGsREFB+Zh686t189NuSFBm9v1EfoZ4tVEZgGNTVJGTZoX5yzNbrH
pep2Y0mdjydVS0WtMokAKIpaZ3c/biNz6AdrmXDacKjmYCyuVOcdxAQIBfQSQTAj
Spuc4yYw/jD6BvI+GayVsiEX1IXpmxST5jvKnhq8exRZaxqvgFWc/mc05ZRUvsgi
htrOmRGtqdvewLz7wP3o8rBu3Hmy5wgoAJGsas26CXmwFzO0go2bf+SxyXp2YP12
FZnPDmrS5nglkywkKqUiy4M9jy9LxTZhaeDvjDndUfNMccNsxjIOAM27sKbqkcLp
O12ZH4WyEFORT4TqaalMWm5sH3kAXhvfFrvsR16kdFl1HqxeNUI9CtfUWP41FEfE
h37+dyeFncy+en8WvidIBZqbgIoaJauWLLhkS8Aafoab1LLYnNnTmLJoR9MKQ8ER
CCOnMlWKLgsZ8nEUg4T2JvPYVOE5R7Z1v9OG2UcBv0vdbVu/swnW4/nR+TB6GBRy
Oyo/TUU6GIj5CLfiYCMMLOLLvLPrQQej7Jlf+3Mml3Oo8M398dlsJkuWegHemcnd
5zfcYx+CZHn/03H3Jf5h3hAMEJb8xzEbXcvmGkxJZgtuq3c0ZedejTJmOsq1oFZh
P6JkK1c1FLwwiInpj+TUEXyhBUtEGG2lJxTKu1C8bENaLOn/Q59Ec6Ta/79xhym0
fH3b3NkiqgYND5okPoaJnAsN9oEUvIBBDGe/t96+ZOLMnSZUp/NsWFcb74FVC3mO
pJgldbmpH4yyndFTGR+3u4KfVyoChdcYU4uQN6N8OEmPJgowJdXUACP31XqYTMO1
jcHF9JIjP8Uc2guhs16y1L3EsRi9I9jCiW6YVkawQsx4LMqmk3xKPQVUsUs8gI82
jouKiH8aS3m8ulf7jfFTQT1BkJ0tO0iKfz7uplF8XtNGClhzAck5XlZ1kxEDNChg
kwk33ZeNySpiNRuvgPDGH/zXpnnb4ePQZ/R5b+08xsuOJ8fsxDsknvNdtJyFE2D3
dn+p48ujUD4a9v3fqmiRY17SNFDGNreyACqqzgo1Vte2UcQP+XSOig56MK2of84b
/JGhfR1NV+sMhwcZLg0Z/RgbxFYdzxyZOiejnsD7SmPcbOaLe4cedPOqiue5uskw
6ocyhbE6bRA8BHM0Wygzqt8TK2IaM4RicvvXa/Jp0hBsKRZwOBBc+uLm8zdxJJ+l
jOMOmCnAwsCFv0RFDa4otrDXiYXnd1c9HtsuMK4o/f9ahvkDiOQID2jv+hWFOyWJ
G37J50ydHfmJ6s7H2Va7x/JKp4TdGOv4SUx5MK7lI8fOjBMF1oyDadUTHPw47IpV
xHnYeSBkAiRnOhdI69UmXV4QMel9J1PXQi/1rqh4aYHBsHQKnJziyt6WSjuwqLCL
scQf0PaMwKT9Em7ojxnyYmoj8Jurf0nCjE6aDg7HfPlH3hVD/lGLZ9/vlEjaJ33F
4iutiq5kjJQHnlWjIsg4wEh4ES7c6CX2ZmHZjmDIkY83XfI2cCPqqmRMbVbOC+UR
ugJZlL+An+jlgS4ocBEeHO/FnNPusu515r86UVldO6N8/evUlWL0ud+r52TC+L/K
cI18OPfJDP94qSu+BhwG6+Qd5DFTtsxmGUpg+umK8z4ekflJ5K3PE48gdyAL0O69
4JVsj4MjFfoZafei7uJQA6mrzz6lrGdut+rPWU+dCy9LDAnZRi/l/qd1AT+6oC4K
Jvm+ZWwuSoyilwFdfjWZ5d3sGbS8DrtgZZAdx8Ar2UnmRmzdeiPFI1NnvwjxN/m0
mPsC7mlH+qRVFcvOoNJdTwkaw89uMcCI72gIdi6I6GHc4cX7PfIywnrRzQe0Xx7y
8faZe0LjMq3s8iZZWhFPRyAkyTSpkX3gn2zswwjOPZ9eT2pMYH0tMAyT2zs33sd+
bzaa8l2tjA1ymIpqFyeOr516wd8U5yS33sBtod3uVNEutaQD2lL/+QuoqiU/RLrT
1cs7CPFrL1oPIxLfDFkuHkZ0+8s6XCNyRPTp+Nhpm94lu+R0xPR5t6RuDXH6CtRy
rlHHrtRVSqUGaF8KTAPIEMvrL4+Bd46lFDLGoftLH5N0Y1m7fDOpnwEnBxDvsKeG
eQzJFffOPzAz5ObgsbLNu1Sb5qUDyZ+leU8sd/xCEHHPo48yu4Z6MOnbloOrJUnK
HrClsHpMc5pjYR3J/x3vPyB0lyEJonyniJqiZuiwS9js/FaOHfEH1/rb2vbvvRi5
GPf1/bsV3YvyLGYd80BlFqLQJIIfXwhsV8dTIlth2iU/n724EyabQUGDjJ4yS/79
O+xOepPk/IPgXFsvotuGRN31iP2JHOGUb8j5BJvHZXo8CvsiKb1/LKcwnuDSMdXv
7L21YqWUURJJB+3teN5AtEWl4vl2E8SsmJo676dNT/BL8osMJ6MJCaxAHkTfuWhG
pShbWCG+ZWinga1Pd3G8lT033nZXwh4FTILYht8L7HSIGEkKHJKIonoerXJdPPeI
a5FZhj8ZxLYadoDOf0D84GZaUmDpCpvdKc+btJ11loifLtVWkihDb+Gv6/UCTtmX
Imk8d6onmpFjd1szPMP6PVWztCFCrBKmRP7PDp6cCKp7Nt6bxb3bteyOBQxO1+HP
tq1stzlLb0LJdgB9jhSUM+xU/fiOsAJh38RFiNVfJR2/I4e7BWG6mb7PBe1AF65C
UIi8vWAPWTqdgotGp10BfOKpcO8ZO+VA/Pn7MiCPhqK4X7dOcYUq8+QXHm1STuV9
VZOfKVegg+7o2/rBgSbTHaiyEuT9MqFcsaqbyp0u9LI0HXtIZc5XmDG874liZSWl
qojbNYdkKXedms4L3b3YwY/jNwEMvSqfKCcIgbXsb9vi5fKFQM6dmFCVkFhXf9Tw
JsrXTC8aqzHZCdpFQ145dDKuTAUo/2/X1roWU8hFWcZEdrnfYG4biE+W8zIlhJrr
G+osL3+Ficvrf6+ij/DPTeqH70HhRKavdx2xqRDu4l3iWw9pr2QTygkGqhqbAiOd
JPwRLsV2K6X3HTBQCEwu+PoGegV+otU28ohjoOlSUkhPH4YEUiGNH0chUNksc0ui
iGCNBPKcdaHIbKXCGO3Dd2LGdOBnsB4NXA2cFg9gqCa2OBm62WX2gaRMf29kWtnt
xtChhjtkBQGwBy9WXQrA3GUslzR7B6t1wy+2ln1UdFkrCqa4Nx6Ab5WJX7zb0zhc
5M2ZqZZ7gNsTvFCy1efGTt1B1G6cFDITIqapW5SsvOF4AM+g3Z1jutfBIEVqWkuD
BCr2A4ebOCpmxN3g6nXGXriRVUYtSqtSeH5asSXtGORrmHNhH0lLVQSEOImyF2oc
tggtRuPSLazL5Ownh3bLLvNQz66zPruzIl/4cVO1Da31rUWMqWU0RxRg4NEnjxap
j4i6cl6PqFnJzcgXmdd47q4+quHm3v4pRFI0fkRT8DEdGgFFCT8HZeBsC/OqslmK
D70+UhHgBOI2i8qik+gWNlv0A00bdYTgiuqb8V2ILYevrUXZq8dW/BjChKSnciM7
vZ0oZ4DOgwOSapMfkuw27IMp350LKKWqG56lWcMZ58LpyCTwnLmGwshW2AjLbyBU
OA1Gga1X5CGK3aqoMUa5sZWxLDwwsWqsw6WxIK9gBOi2qLKZnGnMZuvKpIrQfdbo
IVViepDWDN/+sTKXoM48S22FvEoEoCUAyE6Ucyb/UroptmgF8zShCDNYSkCWrRA/
HbCQ4QnI3QXlUuhYqZADn+ky0F5Vj3fqWmPORzpzybJyuRgXZKef5Jo3JOgQvgdb
/K74Xw8bltHZ2IA/6s/hD3QtvH/pPsG2uNw01pbWgNObwwKoykPg3r7TB9IUNP/y
Z8M1vPRcHYr6IffWCNqD9tNVmZc3xwgnholCMbBe4t6UFAR0CklJbASHh3p+bDnC
UC3YlNigoVo2AgPYRs+EerkurREiokbRQadGpdxq22Y7r5bIrL8UYZy+hWAXd6rF
aDJKqa17yJ0VVam7Jy96cpYYV8wgKVsJ01uVeADqILPhFZPw1w3Qoxm7bMAhNNKU
xIqibkCgRreQA8tDqlebmDGbnPK+FWABpZ7zke/LGuecskMTgFvpiN5RC1VcxREf
ixv8lTDO5g/RnZjyzQRhbgc7KOhNl/ivqsB6ZkvcsLIudClsoi6sQTNyVyVfR192
S9vdYhdLOemDZVM0ge7X1gHU8sZN0Ml6m9LsMAHMVXkvH95WILt6Cmjwzry8qTL8
Y6bZxN1YmMGaugYsuca3igszXnhDbG+98QKnvY+u4wp61BnrLCqxVvKfRFFIxoKn
rmxruN9b4CZjYcbGjfVT48gDmAkDati1vz7hEPKRDDuprCNphBfoZ1xREzYRQfVa
b/Kxn+8s/PccHeZe67vuSfZrEZzP3xgyKPMykBe3MBiNOvyFAuwKRpea277KyaH8
y8GsQxXhzgz7qCYP+U4MQpJ0zJx7PkpCGb8pxln/Ec0osZbcYuiTUECDs3NAmjpx
s/ClxUygK79QGv5IIT5Jt8yWbhkxmfcivsWyBn8qO0USfmoX4zu+C61Kgt/OeoK/
98JywZ1814eQrHfEf7ekCtu7yRaj9I6QS7BbnPDJcrM3bp9/dK8HyzOUczmWb156
XmFeZKW14ThgvwCGf0R+NjhG/luSCLbnKeZ9poEQ4hC8vQDHSY+wErtih+JL2WWv
Wx/WgHGxrs4DW6kUMIuTeXXm3Hnme3sEYr7rSw9P0rFXOwbhoLkaityiDWiCkpDG
PwOR6hNCKYxBo2kxKIQQmbSB0xsPAaerSH2yPe0B55KAS/h3RVVyx65tDwEkb1Pi
Mnovt1n0BUlBT1zJX2fmtFYMLtYZNkXC1BX3jiGlLuZdrAoVDIVj+azrbNeZjOpd
Hp/sKmoYvTTkwWF2o4CJRB1owyE+1aJfU7zihFXdPZxqwcB0ffFItkplDztV8hA3
di8n/HQo824vOVLKRnUefWKgbHAGKeaGfaBUzL5ddY79bv3J6skVgbDs4cBmaC77
DVihKXd5KJIEBZP4eYskuPHNUcV3PwDrQ9N8kOY6TgmF7LVNoD70h+gt4hm1b0Cp
vpIgpqNiO7aMWQFERviRUggLxBre/o5aK0dRUzi4keywSeELr8wY5updeS/cndIf
irqhQRJHw99+1KmFRk0rPev8J15IIGlMgHMFd/ExHdmnOTNPBjhL20r/BVnsLg8c
1DME69T2RRxt0ZErHkYNnTArO6aJn9ylsCXjskHsp04VAhHJWQZG0yChm16o+61Y
H12vWetkNDFhU6hXoZN6F11YXvJyQNJwPUQW+NtqdF38EYc5wc68N3zP73HvOcQ9
v926SKyVGnKyBk051nPPxpH5Xgu6XPvHnGozNF8+gYRVmSHhVgQdhomg3DDSWWrN
8TsMhvID3tW7tfOfRSgZI9GcpVNUvF0dj2lt4ZIc0/mjBZAcCACTouivEMJvbuyv
PoRcwVl9RmlWKOCQt0LHhJ7rYUJqtJuNlPs61aLnMnamgTnxcT7vCMzvZ3LJESj2
+s5+N3o6gDcq0Dvg15PGb1vTIreE5MCuzPGi8LosEzK6nzn7arN0Y3nXcjyaCyON
Ncu9l1f1HFmrcMKpdqqJ6qZtsxFh22qvtUAyVzCUo+Uxtjg/tBn0sK/pbBsHp4J6
LSxsgyBS74QABwOKPqIyZO64MEMAb4i3rzD+XjHfqjWlzq0hjic7sMp+h1Xb3We3
wHUMpKyrS/XKLMPcKtVSHgPeUDHuEkpJUNk984yffRZYiTBS4wH7w7jQ0KEzfLmJ
sO/Mq1tAQ25l2vZ1Xg5CdlT23hoVcN5jKPXcYYqucG82BFprOdLDOSk/qXX3UBYh
Wv6aj4GmeWq6XJvhsVhlERZRtFtxcJWVojrqM0FS0WVJ51mfzZCn8skrjyGYnnGm
dSXYtPcoC7kTTftb2IT2ev847i0nciQx89ocdV7GogCmxN2qzrDwVjXZaxGmWZU6
zOcpjfV5ySGolKOkXYeI85iHLOh2+5ixq5Aah1mGqb06i9lbMI8wRE9aE9GVbiIW
+Dhqf8IxLI0P8Jixq4ZEEhOgO0FnBmZWIbKTkg6pypbBDMsIyKUmieCoW7MQKR3R
HxtkiT8/jiDqQAwfOhtrdAM5Vw1qCbh4Lzxaf/utFpFmV0F6kxYNGglqivCnd6Wn
YE2+Crbynh82m8yHrPbNkFJuR3mPCilt4wvihj/qZ2NP7kc9cJsW2jJI4idXfitB
6SV93sXCKHg/h8Lojws9dEXcemOQWkBqV78uH3uXfM5GDgUyiuVcfLw9UQ6E3jq9
QqmvOXneuAIzRMjRE3fdaj47KljJB1WS1+8Ppivy/0B+eOJHX6f+v3uL5EMIldbq
tdfQm4RA5hMXbUwPW1hVngdkCbmEmHHwmttK+8x76/dgOEGVhEp6eUguH8+vS350
v8mKjbu7QIto3m0TtnYxi1ykGv/a+aHjVKqmSUNvuG+QGxpJRH5t85UYi4hMXCcd
GEMJTFhwO3t5LhJRmRRByJ+wI8uGKXt+HcxofdDDNfg4hkOYFfUjF6/hkMCBAC1x
pReujHSZciujUexGE+gVs34n79k7C3dRHtwo41JOMBMgE49HG7vy/Jk4qYt0rLCM
wbx+FsE2ThXxrN8LMsbGPLON3Axe2/ig24gbQa+CPzVHtKlP84Qz3JBAN803xEZb
shZfPwz9nC845M5iK2LsX/5T3p+hKdI+myqhdib9zkIcMOUYGzTa1o2vlsmH716h
EihySgH2otKeFlcefyLMINc2iPLH6W9eC0tR9OGKIGmJ3h+S8ogjw5KY39WJ9Gua
uv/HIl7qZF6+CYi0Jeu0t3fKmSWIi6GyxCc1vdhcni+YkmyHUK9aMhorysPLu93C
xsejqQ7d86J3q0BMUxviaZvr5YlOLCTd25zlR6FVcT+9u2u7vqwHikgiaAamCZ+K
8MqbN0050+j+TImQUXts3olMeIJD5PJc9TyB26y/5O059yWpF2xPBfCP1p0CFEo5
3oxzfLYkRAOD3nYKjm/bpSCyt3S0XbRcExE741H3GjBwFzdO7kX1sMOfUjXWxhGj
mJMlrk0MNnlqvXxvC5xSKz3ohwD2r4gHkfG86TIOwQ64XYDpW1js8aFYuCJxDMMi
5f3fj2pdO4kGBKyNoQ8KJxASlMHlEe3PA6Uq3o4VcLIuhpg1tiaW8dbPzBO4Q9jj
qPFjcY/+TelDhbdUNJOwz4Wg1wGOYsQqNwL+phrPL7VvCPgbEG99VJs64b/dNT+d
qkIp+eqYzqDqJC/Mm003CMZBdxwzL5ywk8BUSJ7fLBFWCtfY5MPQV1Bf8mpVGUz+
Qwml0f7ZPbpk6TEP/61fuxUtVdI3n/LqKbk+CTT9cOCkj9t9jCZYeOhBQF9DINf1
8baSL7bzq7o9ydsUyQ5nrpnUTufmVr40eeKGE3zPYHqRyWA9THuOg+z6oB6xhzWs
ogBeERkR00qAxp0AtGFlVO8VI/iBQ7lYH4zZ6+gKDj1tD+csFZB+qc9oOZR8uE/P
/oa+EvVzmbp7ls/mrnpLSqAkXq3OENzTNGAqtjHa+84Vn1/sygBMCKP4UCOdPE0n
BgoiUTba0+qGjiMkFdmRZjxG/vCQLqkeVNudhpGR/LR+eD4MG7TpmJxplxDgG8Q6
wB9LXQuTKpAtCZIW7BY7oknCkqHMpe13zWMq2Yf4GBE7oY5aIRdW0giDMv18d270
BjBRB7YhRsfaBdMQ3My0jcgO3dPv4h2IEqnCNBLSNMUoMCnNpo96h6He/GQvnVnk
lsNQHEETyKPSiN7bzIWw1ZIeP/XALkKHsl+pCoruZ7SSocQZNxIxjlzH4U/NmWaF
IGAofYFL0d6/8IQgk1MjpXFDNHarInTC2KY96nQlMMC7fMly+f4IVFX8j78TegkI
82rKTmNEbiTa7SKBzBRcrmdn5AMFOhHclasbE5NmCAu5HOc7qPHrEL3i+Dcwizva
51kM6syHWIL0n6ClzMzMFiDfcRPDlQ6XAMOKYt9z6Eqv7XrfSwqxYQpkjydptd1C
6xLcSIhPkBRRazEGN1449G3daYh5r8K4KczgiKfhTOdZq6bkKC1zYfSr/O9QuCfq
jTVURNx1NNYUJ2VtfZg955AD90DEi8+jA/0D2ChMrEr7ObOCVlhId0SdJojMIrSt
MtC60c/u8ZPqLWt8yEq99h0fnrH+tTGG53wEJONvL08BxHRoP5FCrwOlG4PTBnCy
sthjHfSOpBlD1iY1S6JaJtk2/ftFwYkgM8ZrUozhpWWSZEnmxrqKv2zOQB3HntvZ
fuy7QyO16K5dmWE9cTg9Hx0XycDpBN5652yko1NRJHkqv2cXVfJkTX5XeMs5r2Oc
VButD6gH2UKmFwOwAm83IJn6yFUPjDrrKA/kxXabC1oxiWA8Q6yWZfqAvxBQjngA
/ZOw93MGf62kFxbLzwep6XcFlvLS7cmGLH6SLtr3pZnkle/DQoviC1HjZ8WdCcpk
3BKmQlruGXp1ctC5FRpAT8HZzqA1LWCFve68skLMU60KLFx/mphC+cB7eMoldMVq
s+2H3qrsj0nheaSqNDKjUYdB3corpmaKsJwWSUzJ2v/7Mz2KBiVL5nrmDFj1zy6h
PWVfIV6QWsDVWm/uAmgqsh8nUmurCo/KJSNnnO8NNaaDve0THfLVSG2Yz9PmGUjr
VnxE0H/eCG7RdkJhUDwsCOipgh2TG/VS176hMyrWkjpQlp8kNsG2mkaBbe9+QiYp
Idbv46uur6fuv7+N4NIJ742uGtCjWMHIawHMe5I+cvQkSHRcpzLNuUrRAB/gPVR0
QXqeku0Hw6ueKnLCP6az8WxZqi1UI6Xl5fvcgnPII9mqZ/kt16VX44evkG7Fe32D
HfI+QDA0ovqJjSjZZvPodWYtF+AP5Cm8NPy/Zp7nrl0DVC9DTiKbvc1HExmCSV4Q
Snk0BC9A/+LQs7SCyKtdz8pz7UAjCd+aPCCGaS1R/IHIKQYT82kACTqFD7bWoEH8
P7X9DiEm0OoAr95QcsdCKxqIkejc33FRaU7edMS7xWMukEF9p0jOm99Qv8u83mRv
MQ5AE6Tf4Y/3ERPp4S3pp0PN+fm6W52/KcHo+NxwoCLRCdHpD6wUg8gWBw/EKdau
6Kyirs3C17W7S6MxNXl1ewi17Jpm2lg/JHn7oSVKsE/az2xTJ9+M5En5A6Gz+qNj
w7KpyWEq2L4XSlPHB151Xbf0DDUihvAeunsT0oFStryIHSwUoflKqXR50m+hBe8Z
aRaR+ByaOzeIRJlNlTK/JkVDa8adjjY+4c/OqmNttIhYHNiSP7yS+GtnO2fFF1WF
0mMVAPqkuHahkkSbHfKRO+nZ4GUqj0Z5RGZO7E/yOMGjfAKEXXr+DzO/wmxiogl9
KsRY855iXiT73jQMuO37R81WzvHkbCzvWTx26nDD4PcUiNY8nz/QnF3k4YoOljW+
4y175t3PxpNR8mLaIYESzFp9SE4IHHxA2bkKwwcZK2TtYgQd5rT9KjA1pWDAxdbS
gdkw6qU2PAEmOOrmq4nYUxnVlnit07wkdZPcFg9mZGcG8NvLVRpLuO/afvo0Z4Ve
jRxG7NgY1rGi9lwvQo/GURIo5tOaCwVOOLMoqJSVRBhcN8fq9MSHJ6FPV1d6gnfP
q2Dg9WvDhnwZE8FKA/cOx7xJP9dIGHFmu8aa2IWB7pW+w+D5AFvLsFyFyIcKL3XD
yGg9eJvHJm/IYO/QgPmLsQhamJHbD9linOoBcooeU61kromlecdChdAVTff2ZHFw
3ZpI/orgSPIb2ZOb1dnovSjuHbUrZl4f+gH5X1++OlUVPCLdmOaKssnVPNkGTYj2
MRtL4V6LPkVWsz1HeKjNor2CY1tMukrT9Dz5YAwQ997Exrj+2obcCZVB1iTHpw1A
Nu/31Vrl3eEZQRpANDcKeTcMFirP3zUFY3bzI8M531x5QAm+1oxtvCzTuRtH84vN
0jC8h0Z0LsMICbYSlsVFxn7lWc73TUo+RPx1vvvPJ3Y/TuPL3gTqD6LoYZSFVyA5
bUcq5M17yriEMbhTLrWueRSyP3uTr0pq3ZK406IBbBG0TQPHajQgFFAKFYv4z0xs
lmfKUAYF8fgHqWslw3lc7XJ7dvWnVzkq2mNFa822a8BWpmErDu8xk2XOKti2wwY8
sAJ17vPRehdzkuVk5LgVmW0mXznoF1RXloF64TTlOwqRpj6AeU1x663q3r1kHFLH
eux4jrSU27ewXs4aR8dDKTAasYXp16iyaTZWITOpkdGh0W6PmqcbavWbnXCGxpMt
3uIIfm5AoiVELEFGPREKdCVq2IMbdNoHl6GXZ2I8/6z02X0w+p3r7PBsh9QddrQZ
b9BO0nDzg3qVCsTDA/PiWZ63nPMmetwukYXyRyZHllqYZIUPdOngro+5vtgtqADU
yTMaPhzxp6zgk7sDjiVyuiprAwkHPDylrsR2cTLaW9eFqBEwaO28EAzZHphzFpbm
XRnDf5ZYnzcO7L7KfKvPJn5N2RRqfwwIeCFDYRmU44G9fZRiDErwY+rMbrq7RCtZ
hKoxisSwYBAAoeWRAUjuyEDuDPO4ZLXl4ni2JknuTqRhsOjcIxv6cokpJH+HuwyQ
YoKzfaAMBAJHFilckh9Nn+sspbB6e9vuZALcEUJCyx6Uf+dbuOj7h/r0u2rpg0k7
FpR50AqRSbOYpGy3NISqFSWjAd2mVe5oQVTNlcL7e2RsacuWN+gmgVfx2poJ0Bt4
Z0VQ+ELgwZM+aCmxk9CCZUPTzldQDVFLEeRxkfaeQicScD4JM4P1Scr780WM705i
DDDcEMCGkJXF9MOGhDs3Vu6TJJgF03SmSeFs9sFIDlvr1J2Ih/etnPv4DmlacSCH
ZijH3D4O4tkBnNmM+Bf5kvIAbG4vwiEmyZRlWRLeap7fOZQelYG0e5G+edLciADy
LdCN1h+4PqJcJvXkwVBW3HBGLKXWhAkyRi8F5TgL8a1ToRWEFzMmoUYXnqESHCES
vReNDOGrLa1l9eCOB/nXKVheDOpgBqYUGdUuNHTV/KYZqA0IVrjlRBkpkm3W7sLk
zVbTLRVYdydibT3fKPYN7vRZIqhErbYSZNoJTOPdi2cMvUdYh0DJhSxftgmweYLx
imDnoP8Ejh6Y0kIvjhO5OMhkq9ua6Xt2Kiv+vp8HYUgFtgtqV9tcJ0gXrIu5dnaH
jD+JS9DaE93aCDpDU3ZarqU0wgZG64KnNAFtnKVQziWOHPF1gZWvtJIr37WOkyYw
kZsx4pacA4p6K9pTCPQqsIDf9vD5kIDsVFRgafPs7Q9rWEon1SHQFlhK197uw37m
UMmBzTdfi+D7gu0oln0v8Vy3clnYz6h1fleLRFo99epFw9kI86UzzP/T72DimBWE
lhYsYLAtwX6REoQNEpzrQGdNQjow9BL7L2Y76QGjZWW0+9msHXiiqos3Ba86dBZ0
Zp3yh2ZpDMmd4iVRzIavEGZzLXHdxncYkxXUilVUvyrW5DZqyFpZgHsm/fBIu/dF
nPY6GTbSAQvx1e86IEfNcfj5WoFiN2kLuGo7/bD+y+f9lNDX99reUdTiV3EFrHDc
lbpyJzlzn6kXkm+XhOARaXgCJjC+LUPf5OfqjX/QH3p8CAlFJfjJg6r9sZ0nNorK
tb6VZTP5VqjiHUZb8Ojf4LvJJpokNlwmTm3R9bpMNL3i4gLRQlEjnIp11bUcRjME
tV6OlFN3xsGBvMHrgPOtduTC3m9LDxhcBCMt7fI1YoJi6lM7qu2EpFaoazNIo3+6
H7sP54xnXEH2C5BeKWi6cHFOFX7ejfTqAPCgGpnacxzmATxIdLyAtMrMWQjODqog
9WQDAKAaA/VIgBONK++bTFLQWZN1g/PrHo85U/Ahs/XszEv+bVQq7aMbR5RCi6BR
2nQQzJTMr7OeMxLgdDSfy19ByXZSgWBc+9CSF/xTFiHVyE44yaKuFb0Pgpy9vlDv
3rJjgZJvRVmupYu2KGcJb0E48CKM0Fn8a4DBBY3S2CK2zrC+XAy79vq7FmtP79SA
NlC6JY/arq9NxikOzuWEOKnVucOagn7FZU4Pq9Fw4mkZWyzqOszUU5q84q0c3VSj
DMe5/9R0GGVnW/eTygn+79qKb/nb3tK3Iu0ev99ohxXjra118A7wPZtIOUBRNzCk
2vSatvyJUNL7WfluiZw/cs7GcLBbXW2yG6YwTgLm8txsxFn0Ooj09AbvmH40pLra
E3BH/L9rG2hVwJRbmKiK+QvXPv1cr111Gc4uBBG8/759YzLS5JL4bB3G6owxoykb
83Jg8uj4B4DdkvbyhN+cpP15COV3xGtjc6hDusvn1yYrRdbXMZBvbJS4ABUEQcSG
+WEVuj0531Nl09gan4SEB4dLVLHM15TtQTDExZq3QUwOa/VsHC3zgP5yJsGAiQcs
PRpSgDq7UtVIhYTD6BUCIpf1lYv9Z3bstr2oNAjjDjny20BO9FRA5iWYvy3elowk
tJuHJG2JYXQ6C5N/IowftfAEgp00/scNBsLxzp8400uGOnvsIposcu6ZGfZBuZZy
+2EF/zLE3L+ZqgB7hsohN/X+Yja4a08kWhLnzyZ7RHueuYRnu78K3xD8aL45gQqQ
gcP7dFSVY6LWEv4Sj6q+8kwm3fhO3BM3MUjVLiyAHK3lQDFwwkT1vuZEFTIokaJU
xPIUrowNDuhCs9mladWtzhkH3WBTFg6LKQtoNLpw0rhU1BzMZGtm72FEikYoRkNZ
Hh8H6heNm4wmhTpLkA1UHWCQhn6NXYw9KqJwx69OHcKMYhptIax0VWhFR2tYDyQb
/yPR89u7Rcpg6oiJrGekwDXcRlA5fY/je6JLa6/KXHtIu9K0HEehgzhYFc7s0m+J
nmVo0KY6nZj0As6WnZVUNveZTpUxMujzrTL9tYnRV+wdcVeaNXk9qENTp3eKyQCI
KDZVEAhC+E/ATa0xjDn0L6LgwIxVMccr+30HkxoLG5iSpTxG+g/z32+QuX5hJYIy
z8F3Z7gZqkn+1dM2j8o7wNpCuvFB2ytg0gU/PlzTvwvqpnHQQveuSixW0Vzlh23i
TScypgFvxmETc2nz8t8y1O26aYks4EP4ugaDOSKzYC0/URV4UvjKI5NTUDnoHiN5
Zk7sW1CO7V/mtDO+lXk/fbsVfB7orniqtGaRDnfrB8rLhhSJR6pCJMgEhBeHUgLv
8XGo17DCW4LCi6icjJ0u+XnB0RFS4v6Vc/RoHOlwNG4vpHsSc4vYqudsfFYU/FZ1
iApXv+LaUOpJ8RDaYV4sWqUT0hPelnePE2kRGo/2cXx7sRN3jyxaMixe5JYwZcm4
Nk4cTZ3ADlbdW0cNGHjg+pY6GME3ijwlCOLCvJxl2jhoaqGCZAFx8VT0IsAiUTtM
CPqHzvX9ksrD78VtobvllAkLTEAzGuStd2xAM1KJn4AzrVH5SXTe/1+yf/sJZ1Wd
mL420bYxG3wsMzthIOuDXaxl2kh0QoKnBpByuOmqNQYcPKM1uEGHBl25BqSLemVw
4xLpmVP3vFQ9jdjM9bGyWeDhkCRzc36eNKJMIg44O0q5u6qu4sivT6NJu/ZvqPHd
Qz1MtqejPIRMn3Ip/f3LVOQfSlD2SIAhfdQyXquzP8FU5inZcP/bdQDB1Q3ARWE0
Co5khcKe0dalau1ufjnnPDJMoXOlJNJdV6qW7gTEkqDGwcwzO0j8IXN/qiobXCyt
Al35waOpH8ou0hqL+xbU7ZmJAgHpUd+AOlbigmhZeB1PvXskubSp0FcGmSMUd1aO
S/EFjOTHe7bnwa6DgziAsiCviOnUzZktL7E4b59ClY7O1mEK4Z5SsZxijLodA4rz
jEiz44FYx30U4uLnqubwrZiYJG0fkNRzGW2dEJk/tWk415p03yQwcYJ0jBnR+YWU
8AnZ3LGbYSiDBPTM1CaK0eyIpgxmMxab9a7GijtXA2hq60be1g5SE7Foc2CQLeaX
Psc3kNF8kl5RERBTaRT8eWlDABkyktet815vVP4O2Ty6Nf6APBUQbEYqoJsHkhTQ
oLUq7daWvAMNcR+E1YACIt1SzTbzqRmGnSzQXfUZCrzCSrxhtosaPVsvKbajQBkd
wy1DpczAzjknz1PhAL43meR9HiFb367tkGvNlrp691e/Tjhro3o+AyS4dgcyyAqu
0ZGrsyA9MB0H4/COa1mM279/f6sEf9e/NYcBnkv2BXPAe56h7OFfon6QUct2KhNs
XvdAIk1G5L10T63dplLp8+lYECqwvFQu+ed/Cph7ENNdPIQrlWXd1bULPVJPUcUz
pAKEDo3tsFhxgNQz3SfdLwger97nPcyVP4k6sy1E1D9ZTqBIRrS9h1aHvh/NQ5f0
if0+yCMhlVj+5c3GSJ9CT6eS72b+n/V7gtEwalqvsS8CvgXSozozvyxkOLd6X4Ln
0MdUhesTAiALjF1DZUEJAP9O+HlsWFnn+fJ65f09zpk2x4kSQ+nBJ6nI0T5clO8a
3SpWOuV+mVETlTMhvjrOicpCEmlarGkwPeuws3FS7GwyEeg/2vu5WtOb4pWGs5oI
vsnBwmbFROap43Xyr+U5cD9wIAxQl1J643niaHWhx5BYdFaqgJRw4C7Xji3+wags
Hf2iUxIJRUQqCqLc4OeBYlNVOejVaIAdNHek9VJKYmfMvc/gKSfubUflHWKFrstk
zLGgTcLGG3uXqTIkfHU4hq+0joYqxzhQVrlFIY/Ha8Iz8hTSDeP3PMfzr3pAML6L
5LqNBi1iZ4vEXxdCcy1KAJBs5r9BedkQqH6vF1h/28kConeraZtIL/iQopWn9bKC
Bp30cQqZCxL5v1e4YikXJNPc7M6hrTDMem/h6Ary2aZ5qqOQ2Ymp269ZEETa29SB
z5R5PMlf6t1N79NBUifD2gvmqt+J6aqY/O5FwK/e5BQ87sMwFVs7H0xK1TEAt+nT
Wtgc323iYk5Ol1vk3IkFlOgQvUg2Cnbj3SCUkC7QBzVpAZQMNIOHznebMa6Le/B2
loXuQ5AD4odJAWjFbcZP6CKIbLiomu4vx1YIjZgmyrvVNnxs2ukmImQ6qC9Uk2bf
UaxTEVj50MpMaFLcqj7uENkU6rCO/1oE9F2Ir0kRTEu0MZO2zyYDAyB/HG+g1nao
TfQeF4BQ21f5ikVBFQR2RT+1hpZJU4FRg+yu+Uuc5uoCOoueYqJijWGvrfdr2a0s
fc4afzt2f+epNwfJZ06DukBfMiHxfnpYYdcUxjg4wmlT/Tx4zaFvKdtGsJpT4r7a
1wM5GleUwBrtxXWGfxXkuIQKS6dgNvPjegFK4bL+95U5OLJKxf+qo2MFUKSQsAK8
7VcEse2M751fEnmf7xBCZrbti9xBLSCwAgGYZMPp3D7kzmEymB0TFQvE14/V+/cq
Xm2r449198K6HY6+0IPrNrNfQp1oFnQKe9UnxpgaNVJlaz4HJWuhyKOSZBLfKgB6
1orMpFapRVj2T3EtV8LFG0ZtkVsnxQVSGe5OJDd9lm3aVwfXOEhiZ1evkN7p11A/
TTsfbKZCbEFU+O7/UeZ5lcuufyv4xYhdK/sODgVPd0oCtwORYX8aOT8VFcwxaHqq
ijUEXr3dwnP9lblHfZVgjV5/b7r/m0QCtLXL+k0oPuML8aIEPFCPqIcjeS5T0d0d
gcUDX+N27nz/cErVOZ7OAuZ6AkZsdRV04MmzP1B4XbCRVxKdzNT8/qkLgPlmUJ3p
0nNwpXNxApQGAOSaEYTo7aPlucbwQb3suCZDePhg22fuwrrs7Ehl4vfR5M0j5wNk
jh3awlGi9Frx1ReGzyh1pJIDtvqi+7IZhTadVg55hnVbuaGHZ2BnJsxfrkTpsRVq
eNUpXUnnHxwloGg6tPsDTukT8QXbuLzAPtOCjqK2q/5Qh0gO5JXKnlKm1SdQ2wXD
tk6GSr9ts9lYRqQyc+dWt+bqc5ILSa7F471xFp6hnOsO/y8wFLs6krs1KJdV9ELY
nlcIrlJyjBNUE6IBfER5RxLFSTMwsV5slmKfJkkB5aDxN6thEkjI4DVqSknbSrx2
ec40b1LP2n8jtvUNzfz4xx9TODW5qYmXlX+cugqkEywLaunsFsh1CK8Qp+zhhPh6
j+8iQi0sT6uH9+Keq5EeOomzqFKMJQik5SNvnslPXsAWBH+OfcbrSMlrbpDf/t2E
EsF8c7gnZ6+U2prbhHkXWICReRR/PimsG7FGK0/B6Pwf+1OhK+Bst3iE3+1Bp5mX
+ZBCUwGOa5OCn45GimBWxcFlCNglexz0+4xm+7zwGystrpM/aljNjioxecVJbi9v
puJizsMUeAA7YrCJcAx0MQ+G6OIwvUJgwbpjaEp9/zDkghSyeD+3wsv5F5Z2qrmn
yak4QcMpT9PJnL1MoppODXAkn3GSCG7dY1f/MNH+8JxeXNYYXJ79TGOlL6FCdiaD
D45U5vABxvZap46k+vhxmj21qMtUNgpwoAP3v1fChW9zuPxq79aUJeG22k92KAOH
+vQRpfbjzxlK+cY7l4M1PMqdHQyuzeTU/ngbL8FBe/l9hskZx4u/v23aJGh+GR6i
6p+nk+OmZhbEakdMZcyxU4qmoxPf3/qUTsR21JW6eI6k8OcZ2D/Lo7Ph7vrG29oE
czzplf60D5loBeHCZDHm//WSf+7qt3Ad1Q909MoVhh+svcThWM5aUzQY/ZKFPFLY
cwKHupXzbbhiptz11C3DdnhDWY2HGOAf2B0BxfOzfIxZAgCV2p/JZXflNE76L7m5
zWS7QLWFLazlKSAcjiI4PzV79vK1YHodTBHB+dpx5vLtV6E72/hvRxPrcLEIPDdm
ofA2vkIfCOSWLahm6JQQMMtVtAJOGXcv5nqa4GLGAtF4N13n87Q9zasBzgY3e47m
65NWgxvRa5dcI62sJ5poBOYQl/6ngckmfxVF5YHjHqIR0phFuwMTfNo3EIeDJ32x
XJcG4bH7i/3niNBU0uUKDnCGjSPJ77uF1oruAu6Df+AJS9PRIIHaApqH7XebR09+
9ybYLpVohjdhBjhduWsatttIdgG+YpO+vtdABdNU3XW1lRNw9cmbdoiu6yvWqdr1
EVb85CMd6HXam4bEyXpjjcvZ0N1kpQsKJfzkkv+vV3KL3EmWIdrT2s8nsaZa6nGP
dKCdH6g6B5W/JNyUGe1voVCNAe3TYbGxhZKD51aGxQaYYKv18MWBwvGL+X2W0EUh
SEMoRPeYXLoNzAtcb+TDKX32V/7uwgfzbRbcG/W77HkZDSaoKgzIxzo2Wokxqrr/
amtmh/vt8bnvFIEahsLZxav1Vfj/dqX31Ew6iX7UL/EfrXZhUOZla3Cb1ZCO1Ml/
3GO5G4CLAQsWfnCTVWyHD6B6G4Jz8/IfEZ8O7kbxHmV+W3W7esKOellosT724g6J
eMAP4KgVpFT7jPHNSXH5oQQAvmyODuLiMwRxY3n+Ci73fh4UnjaTrShQ06x7+wi1
6OGDsTIxX4kL8BcyTLTpaP2tf8F1lrhMuyDI1F/xIxA93KCP40zHk95CxTwsUUTt
Tdnfxuz6E/gjc0GGlbPaZEM4jrL5f3eeKO6eonpNikr7nXCiPe0QizAokH9UsxLh
QE04IDZ1hrbYzThBEMVJSfG21R86oFHTrroCwG/X3zD0HWIo+UUN7Hc4bXyjLFBx
9DzVrnSJSjCDxXvufjeIT4GyIJRyhN70npe7RQimaMz7FiH86LYCCVCgCVy0kvKx
jluRzMzpuXjtSH6pA4lF7Wr2Q0udu30jVFHQeUyLm3Vv4Lq5HrZJYgrBucW7DMwY
f8EHqro49gSwnjlIRoVmaE8jRklWDLpYtw3XJcxQlGZI+HhmZUWQLtPkacjX/oiQ
bg0jwPDCVc4TpcYJKpjiqR/Kjh7lV/O8/F7Xca32v5qJsX9O2z2gUrnGKKZ+UR4S
jIMhOv0MTpAaWKGz5WOJPJ6OoeFL0wvOuz/wm0We0oFGrdqnPhCjlR+p+h0y0bWw
FkOjYvhyLKQy2a8JB5nxJ1L6K2NvU+E8hi1BcGo2Pv4Y0L3nHDak+jtd7JDacrjg
+TCR85qnqqcD21+J0Z+PJkAj6ryr96gzhIrbULsdWVSjPHXzp15dPHJtRga/k5Tw
YHXL77IPBrI6l9f4Lsn0iQwL9Qa9VJZNXUzDQiS9uxz+Clu0eCEN+0tH8AZcWt6a
1PBFyzRq+QQRzaE17osIshxmAgTftsVZ7RkJ9XXLYyAnTm9R6EobxuSy4Lgdl7Jj
6TvJqBKpwkwU7POZC0thco7rzRfJUQnjGgPVGxgVeXUcKwoFA6ImGylSSewm1tfs
8l7glXQq1Bo0UtC1yOOMUryldnmFrdKy2LQ9azlMyu/CjJh7MjLuIqRntGDREuqH
VCcRojOAVyWum11Fb4cPVLD+sZ7XXA2KAvaYiZg3RgfeVCspqY0IVyDenzwU5ael
J9XV5fgFK9p7tZ2Z79sIBsot61iNxT08mrx7uYuJZ/e87ozce52don/sT6UZoxoP
WEfzWV8Oi7s28o+QQ/rddbFN9nu7DzYuMnNXy6sNj7dNcjAZaWPJI7NlwPhJM5uj
n/uUoh4XLR1MOZO7OU9K9aSB/CV+qmJFNRNOy4NEP9z7pGrtaLCGC7at6VTSDlH2
TdMQQ5AIiz4VhmJX2kMI3k/OG8AT/gpZyeG1X0bHUEAre4wLm0qk3IDJuHgYASXB
+fjz0XPeVKV+WfYPpbTjzm7lSh5K/dTWThaJoDCURPkU7mbVxCHhzQhuY3jDM17I
pvlWOQo6pup/GQQJvJQjDWtqA56cEN+wmijI62kRN386QRyV28yTZjDxz1uyedpo
feBCgXxr+Qz2UDtO4pdj6nSu8DZSkDCpSo9n+UsdXRj4CZI2WUmZkVeybrcrxSVX
gkXmj1Bbc/HVaItoWEQCtaSxTPJR1gLMIV9tWipYe6WtuCHhx0ojFM1YZJCdIsnP
YPIHcdNvwfTSqIqNSHc7YhavWKPy+qFqo46rcMvXKF9tbegelpK4EpwpGtZAonoj
2BNGrA+dj5Sf1gmMTWIchLyB6QiWg++HIC50EvyTJKR5lIGMo48AMFYHW4K7L60/
C/XAX6ImTnboDVdwc8sZITSNW3aJTIzsy/x3Ip9AL8JdI9y/1D+fDftl4mk1WZhm
SiDO5vQ5hnV+/fR7slrCUpCiqnPu6KrtzecHYmwVtVNtqu6+FCVuRQcR87EgUxVI
Zm54QeXVj38owNifGWLZ5GuwPmdFEUFujCmJHxDoaWa936e5tE2Q9lZ/FxsTkjzn
xdDd90Hr8g+SSLPbWHCJepWYOgU1Ese0EvyQ2vGkz8tkt5SGHXjODOW87ZH+qfsa
Fkt3d9tNMp6XxLQdmxZ/Om8vY9o2jetjtb69vT7NeNcxoV6GW2q527+lj51+TfyP
PK/AmvQ2XhVWBQ/aBndaiyhSp8ngzMxGVuclO0353puBi9OaW/SD/kO5kzKp/1At
ve2deViXFBLBsr7YBydIVG+uu2PData4GIvOrzWQQHrX+ene3cpRj9xWdTzUVOle
lpJGIrsiAfUWVddprwCyq7i8puJlRgA2EY7kL8ernjSOrWDINKzfTlNKby70WsFI
j+7AGlNUzuQh3opvtQAT8nEgCMISed9bUgftu67kBbKjj3NZWwlK48BHivHPK/wJ
MhfQ3qoY16ZXeXCRj3sDcylqT1D7JOjyYftw0sxt5jdsTx3zF5H/GhvGZ9/T4V3E
SVZN0ZOZkP1OUhR4p+gVAJUz7Jqec0Ci4Fgsm5/SzeUvP9PTWiYdylY1tMr9V5d0
hQ21qJn4xFn1cxQjgjKz3PDPPpcsppWz+ndiSNcjlVpxym3S6lTWWkKuix1julW9
2ZOVjVhoX84CIXUBiRwvUytxI73OvDac5B9XpatlwO/iYT1GJk1PBlvY2evKRmSR
r2rYnQX/NnshwXqhDcuYoGbtzGOTzGzg7qPrtn180obcQ5Rb5iFUJiSmhKDMKD8i
OAi8Q+LhcD/e26cxRypb2C1fvX8yvlYe8tanHC6l5gzekpEkjGD33E8wTAkQYJg+
WYlxrsyLo9T4tOhuwfIlGZ5zJN2oqMYxW4CsXzJYJOsJcA1mLyli0mz4zpQbvtE5
yT2mJDpigMxstkmRiB6gJhAvhGIzF0SLJ/kOU1r/tQ4AL+F4eiWvLS2lQcA2zdei
9y4XPknE9wyd7+fXfxMlUppuFHRIRpcUajZrg57r3F5GFly14cum2tEUcuoD54FH
e3QilGO5+/pUDgS/uoqlxYX6vlwRKs38Ft8F93HZAK7KRVlUQr258IEfkowXAXDA
yyjuRDKgiOgp2NZyoC0b2ruYUcoQkSrIZEbyWycahZh5D0uIW0iQ2+76pFHAlIEE
ZxjSkpd1/qsuozQ0PF1sM2KmeU6VZVGV+KA8S19vJ9iaGKx513eEKYOiH5SS9GJF
n4zesc9W2ypLE8jV11YmLNREZEZgOraPzwlHUxZxfQOutjtbysr7hw3MroQh2AP9
WCDwZe0J9XWTVoTFz7sX+bgjBogZZiUbRYUaNzmB+yyJV++Jh8E/ubTUERfdtBjI
z7awEOnTEoIZKrb9LmV0cvz5jDnlXrkW6Npjuh+Hdp9rvwTV25pdnaVLgLqMPROt
KaG2ueLb3BAdyatI07LCUM3m2XRciqq9kJCsoP1QSh67Rd7354vOYsb7bxl6ANB5
ctb9gMyBLPQNgRvBveMv1ZsNn8GkOBdHdqFw+cTVNgjTetTJoJhdP5c9XBBSigHK
ggJL3aKvhlzLgHX17h0DNMadDrz9Uz4kpDr7oqpqe/RuPp5n5wz1WQpSWiexvtWz
tBv5emW61MgRrQ239spdZS2wZsD8wlxk0FDBj522Gx3okJUPZYQivujs1gSSmySe
Kk31CmLFe5X7zZl79snZMiUHcEL8ww11BXmEWkuqtDdk5AqnxiOwXDw8Dk3/KdtY
eJfOW+t4cHYJVIzAkh3gw/i8TY2PzpHlRjTwebJEpKG3heCtEjGgLcEMD9kq/ZEM
svNPmf2XBJLvXVJefvQ3PNDHrpio38RXh2wUzPvKnNPXikgj92kUEBckIolhrUI5
Jk2gati9fck1SCC6KLaNHIR6QJRUiIg/OXKrTO07/KOFX7tBlfaPVrdYts1/Qz1t
8IIw+WqY15LUz0pWkSjITY2ZjZXqUvCltQ11i12XkQlk8ydR/D/F5Fp2hwuvtUVn
7zig59xCVbtGtXTEsQiiSaTAVr9ymcps608HVfvewg+IOp+SHmxdc1iU8jiGhdbM
48Lw5lZfRavKjAvZL/s7bBhh8yBEk3nHvl4sCKHqTjSOUjo4ysTkjzIe88c9oxwA
8+DGp3/Jj7MaYTbuab+2uqpFfLFKk5uSA7JT4oStKNUCU2hPFq96Z7/RFdqjH59P
0qc9npJbS+FTcKBQwnpgHJCeLE4epBsNOWTxJOPM0DlA6xS0WNM90btxaxHOrLe3
JRgDr4kS6rLs6xEhYQSlwhmMFSQ3BcGbQE+7sIId0/X5zw2WFmP4dGPy+KfuupJl
Z0p3Jt+9itmuz/EiIMi2julHuAXgykTn9KgrnxjZ/Rh0ZerO3cj3pgWKHrd6XczL
8CEvZ/Eho4fujviwOX2UimXsG3wf2TgyblllperxDdl+E61iue/gACIJ0PeDvU6V
9WlHIeorO7odlbo2LpmLaGaRumSF/6tli0jH6ftnsbS8Bo0uRhIUDi5lgf4gh4rm
przeJQS6djUv45KeV6Fj31ajwNBzVunyVGpJwSfGWni1Qcyxq3CHrt9Jc06uaTF/
tZbWK6XfNna99btTTtRgAdDfczX301CQuCJC/QAmg0MFAba2dNSbHpr83IQ2lHRe
RFdRKt56adXjBM8TkwK5U+dEuqACYDBquyjpS78gfOAGHnFARkVNW/64EhVfn8Y3
FoDZp+anbniae20uzjTthSPoeHAcPIq1jlaaNwVNuzpssuAF/KGLd9YbmMVZMMsH
ALur84JHrM559H7OON1UNOVDum/Nhjm1+u5cgR1E6WpxmrQMRGG3SX09e1aGrEG+
0huKnhq2ChXsYD44UvxGw2cRiAb3uM3MXJzkVwbc3vZ7JBWMHOYuUpD9mHwG365A
07fU4oMjEOTzU7Ai3EqWvedtCQstaqG/tJdhxsmrbSZv4nW2lJ1bdLO7BO/OFaBe
EPBLZkMEdQ+isPi0oX/YGna1Wt55jtQC5vDckgaibZyfW65+zt9j5/xfuTLPHZ3i
A1YflYNM0rKAbkmi0sLQCXC5ekLHZvKcBSr2y29PmkFfsUbCypwxD+S2EDJXuURZ
XW+Swdkh56Z++q388r1s5nZ3MJZSt0UzLWnmRPqHFSCJzM5g2tkHDu+kBn/1qjxr
EwfM7OA3VrHVE/8rGaZ1UXJwBNkYY2Uw0+Dk5Jsilq0oZnOS1zDb9tvpKuljasL2
lXTdbAsi30Ni5dxwJYQqwTwKC51ZsQaRwBKW6d9AAkRWDNVvRAMPULhf4esw1hac
6n/XfJ/UiORZHGjsVJVZtIoEi6UVq9wra9gAl9gfg27YhZUEVgn1N3Xrx/GBhrNy
+FgwUNF/yXmguK6SQiSaJe/MKGvn6Jbofgqpje2+5cgN7pRnVMdD8IY2NVfcZTnl
IHDcFj33sPBPvldOt/KGbNtxe6Lm73Q3C+LDEYywlIUPaQi05K/u0QHST7W7A+d7
2gS0DUnXCXNnxhILQveTzm3+JQ6S4PwSqfjaQmCti9jYVdymMazns9HukpNVxH+g
nvdf13XDkvAtT3B0szXdhjxuwjZwIdfn15nIsayHDui58Dff7R6WzVT76DW0wXLa
/0u7K7mplP7SlqUPS5xayAmkVkFUJzAKUGESBgEzRsrJK7Cob2OUjanbbz0Ba0TA
/8Wrdtz0HJP1AGxbF2IxVtVJAwMS2O89yIUsZhUgXoppVjNwgH1bbWo4m+0bxDU8
6nPA2pT4mU0FADzd2FNOQCmpFz1QBsublTnDUKtKd2MMqxzKZw9450btfq3pzRAL
rqy26I9mHQWfw/bJIT6Ujg4WvzHCPUlxINb7SHOmy+r0z1pMy8/0+WXhEiagfdax
mg1KZh7fikxIUH05uL0kCOaBalgdnvjVBvpcZWuvLnkJVggCh6VkDnEvoKiY+AoZ
QhrvliQLCXJdY9JOXdvdd8DUpANghBa3ig12kG8fpEs6qJRDD6TF1DZfxc2poIM1
4oG0ZJ6h1xVhrLBDRJZtxd2CpjWDjs8cve6quVZIoK+vVLINaUT5M1jJPifYQavX
gdPt2sg4iOjez2ti8mXmyFqWg3idxoizcxP+PYuJ68vL/QWHH30u0gAVwzzhbdHF
IKeLYZVdCAuTRK649Bu4/LBv0b1yxc2zLmoVlEOtLFw8ZDhgc/sVrvCzHLQQdtBG
P50EbGCRLRCUuF3mAn9MVX1hmW1U3b9RjrK4bJ4WVIQWgObgs+UnGpJBuvxi/y5d
VzcuqyBAuDrWOiIuxZoYkkHKXIgelUo6QJfNgw4rxdxxyBsnraj8IV2nS9mxXeuB
k4+Td5zjtvEqIKCXxlFYftTqeWGHyZ0QpzjwKr2CLvYDdVCHsFkqybwkoruKaUXA
ZEVqHNIydOpAfCtA0OrvzpSQNPh75B81fEggWw0GVVTCP2zVpqqapZXDobU2lcoy
oNmyt65p48LFPltp0gdTwhIzmmNe+ZnN2xDFCsx0RLlE8fSVYdt/rsf83a16PwUC
cAkL5l3yloD4+98z+uY2cKtb1w8oLLgLjFynU7brZm/ExTdodVA7GxvtCzV2Fw7U
+GtEfPCq7kCURdMUiCG0nj16Jo1QVB2Oo+pTlJFiWPKIGBggnN2xjlMpEKnaQYKB
CE/Ix5YfTAICqVRWNG/6um1uU34NHbhLe0fy0c63kY5og7PiQIw6l3zCyQw7tycF
hRyYWtpXDzG6bSkXWIVaUpyHrTumL0MzsTCiEj+faWpVgvtcCiedlzowetSI5evx
CCcnPJ14DIeZ/W5bOE7OmgmGFAl/sdYdzH3uNwfeNnkYj+nceBUdSWplnJ3U6ISF
0Ot1J8c4kgOZ34qgc1GCVINSCLery4o5PDgCJoCw5Gerl6iw8HvL4XSSSWG0aSMb
O/zm0NT1yAIrIMEqC3r2clekNoiFVFpcFo0cnW9hJLKduhODIhn8mT8qzvO/nxCh
uCFOXuNFYKWXDs99WKtCqVmPioT+KRuKp0704aLedWAhDd/ThOSQbzKvUjrUbBUl
5Tfr7NVDi3ik4Snsvk9C/qW0ic9i71608y4s3Fuiv2VHJne4RoC+e6QhjKqg+Un/
Jm+2Ir0eyfdjeJ/r8j/1dLU86liqbLbTBzAytRiD4lYlhbKros0B6oYdMSWb2EmM
Agrg4RR5jBAyiDUZls/xJutq1Yce3T3AK6h+Pe7d5IMww/acWFjhEAQs/PxU21Pk
+Pg16quQgXsCWEPbbPGKNExEjCfQWcc7LZdrHk1klQk6d3Pv8qzKhZYe7+qqfyCB
+Q3nhbw8MwOQT+weZctNrJsfmQfCFjZ+bX0gLoVpBw7K36npJoBtAy28GoZEd22n
Ied35J4lLZYPMnf1csQGDKN/f42JWO9ZHznySbULoEtYnsnkvt2mMksXHTTJATC/
xavxZ+wu90+blwXRKdNfbBbnG4lGwKs5DaYImcfeHE5ytz5efX1E8IU+hV18SCiS
4Aku7tdzNMshWIoaTKCXN7or4+HQrO31LDepTZdJn5e6Wt5FIiclp/QyJqIgIUuK
ZxfYlf02/37/7g1Lkwuod+q54A72Rd/flDMG5CItpZW5bXqTwpjPZ+1Lg6IkO30X
CbH1oWmLJN/wGUrEsIM6f9CZI8QVoZtL5rh+x8VHKCkXkW/opOqkupo0Rsp6emSn
ATwZz9xb4iaHLU1Dozxba3Evb8q/L4iDMBSVVurE35A7V79VtlOxNYkjQctU2y+a
k4GlhRN3UZ+6OOez8RzJIcezv1yH+3rxpoUJeklDUJlutWHIgp8aM3sAB1whavGk
L/ngqJTVnMJXScjend6sQ6B/Epa8GFoMWac3v2GIa40GVlYglRt6j786Hz/YF83Z
8a3q5DhUtp5bGnSXsqsLCJDoRRFfjfRCGW0R2YS8crGYN0OxhIqu9FSuG0bsp4/2
kTWJkMy/EoHTp2GSCzvXGJrrm1DejerxMVGSImXa7n/VjGBMoGPOP8cPWZ6TvNTH
idko5vsFulR1Wi9itzNGJ0ShS/uu6CcuiU+mx3zFtiE580bSB0/SG2K9UIz5N+xK
u+s/IpZtuDj1IG9Wr0TXYGVuc/S+SGfazzWMFazsTs80dlAyPO4wpttLDTw+bsUa
YS1JGu4GYa6CQBwW+lRTgI8k7b4DqlFHqQAKP4SJNM7IJQKXYA8YA7xAYurZOsgT
rwf7DzrIhy99HknoZ1p3ye7yMp5u5ZMPRFdvBNbiasEWR/pgnZmZXrC9iI86YgVM
5mohaoxSzRLnItaNAIJGR9P7wUjhwMAQR2R+qfT+rqCYM5ECSy5/g3Zxt++H3WSQ
qYA4LbBp4eII1McLrZRClKvVAuvjRQpH8p8axXRxMcvYmSsDSrCV1lEKGpIWOrzv
v6q6OwrcOAXI5GW1SvbpgiCr0Rz97j48Q3v03QoSqlUe4z3EapSZX/tWiyeDpQ3P
0e9MrLeXjjHlCfJU2CqYnzbgtKsPQ+9+c+swH/V0tEoz7BOB0Xd/xwQkJNR6RuJt
LxnQGv75OtyJIDbi2Cd9InjgNsygq6t/dtJ1vIBOzduxPQJEIxylhS0aUYcyH4DO
f5kQH4CE5qJxhLGhsUFQ6jMMGPnocDz5I6cfw+JOxFHcBjFUPcypWhU1q5pEtH1G
VeVeOwz0stwQsNwj4BPglUI5PJt50855wv9txongES14uJcMqXpEYasSrudnX055
GYec6fLj3PGl5zTgiPa8WHxb/WCFSg71DYipjq+PgzMhGGqqBTijGKUxUe6+ZmJD
351E9zqM8oNsuGzadIm1OxLQEBNY6p3QyM13Jg80gNzKyMbg6zUvJTGHJAXY8MTN
nMzInVSa5btpoIw7sxyb4lBqPej9QJ3ZIFc5LmoATz8XhOCt36wPVqhN//YmwvLO
qSHRYUC++xJaqI0SNmlKMtQSyxB1KE7G7mmx16IpKqIMjEpNDeW92h9xW+kuKKD5
AN8IT8txmHyMuDwFN4qDif9qBNqBUy5cdP+MjlYt7heF1HF89yyHKDg0+lKAtWys
2QYqBkG6vvmMtOUgz2exEtKN00mbchrEfPazB9x7uq8dGHJdG/fJCiNiYw3TUkzU
Q7rzHMzNRkQM5z1PNQ1x+0nzGynJ6Ce4CI8NmDAkXVDWFTr1/CXyrE0tGIuWO/Bg
aUalLUBpK5s0GGkC9jpG/KUPFXuQs4oYIlunECvJdAqe/39CTlkS3SA02XlGB7N6
lDt4z3jMKA9QdX52aXispFiqta5/6UYLBkYut55qFr+723myb9AuAMU3PNknjCuh
mIjz7bTDSpASexr2T8VisgdSsI1/5N+QAqgAOuSl7ug4JUkDOPsYrldgZBWjSexX
WXlRSF3rpCmSL5rn4Kbr55igKLQXNFvhscKDQJyjL2qcq7A9NdcvUq3pRifPikKj
nh1tua3BZcKC2wK49pZpFp14EgE8JB43qV0iY7uQPSM5i0wsiOGjL6KNDnT4XI/u
JwzDS33HqV6fIBgsXjE0uT9tRTUrNB93q+eOsclDqHmV5Oo5NxoCKsEe2paxXyNx
LRy5esgsPszr3CAJCRzZ0emu6OwnkDo9e2bAdd2nd8SgsrjqW49O0fKa1hB1O6bs
VFd0HSCkr15l4Z1gjINoZkzl0mUYJe1J5snoKZlPpAEOgdbFZ1rcz/HJ3CRTMB//
pqcCbfycfbUCdxzzVHhxGa4inEt7nxbMTp8J83LMwMGgpfCuc4yTP+uMGQeBxM4a
iGht/hFe2Z1+IzpvFaOXU5VkqPWAcmMLRvzc600eTrKm5fxSZMtVwmT6qxmICE3B
9rEYie/jU9+Qh/5Q687qX1xtstazKSXQsC1So4q7BLz77vmSfyANa6PUYO98zelS
gMglR0lF0pGoWDA/U2JpE3TUyFdQH9/+ZAjcTYC35fYLxfB6V2C2AfAf1YwsXrBe
y3xRcI6ZsstWJ/OW1zLOY5c5Ga3/IJTFSsD+EC0N1EDASTMDELbeis3F1RwViATG
Qc85pIloGsxaD+3xfJuOhRYq8jas2F/zx9HJEXfQ6vmC+ps+u9UIFngtx6pjpzdo
L3oPARDDQ+0Gw+4o8kvnqN5g0kNKr7oM3rxpEAzUywVMcTNWw+evBHiEt1+X0Nkj
MPtyYI/ox3nub5n1xAYdFnI8V6Wt3RTxiSrgv0qaCv7cwGSleUBVwnDLs7RZi70p
7zMw6OhUjqbX4/SBQnNIqwUx1HjlerkaXY7zkgQ0KziDktOgAEBabO4xMhr64p/m
Fjq3CBeBZEMTG+RrAESsBXQ/O45PStwQ0j0m8xtH4pjQB411VkzNbClrh//73Oob
MUrcYsefnBUO46rR2iX5+Ff4MYOGSeFgLTJVDWf4Av6k2K6XEo/wr5B8hNHsmnvn
E4bo/FPgUUKY16zZ/38IAbXNnnebmNQ4bCWSXYXIDbc7WHItvBKGQQrCj6Kv7F6o
yOPJR0z56ccK82dKRlC8OW7aaYsi1m0dDAF0SJgELUkpZMiasiyOnf1nV93LldF9
AwFAxEV1gV9RS8/IEp+J3QnxkfDUfo36LCccoc77tNhBTA04frxnBhQScLmwqnzL
0TI6JJbZ5ZGHyYjlqRfE6fwqVl1uTPSZz2gcIkgN/sfg0S3DTXkiDdBXYe+KzUws
ZOyuY1+vWJOoTVAUwtf9SPxOVFKT8VXv1LK6y4UmCYHE1dNn/p9dfpFStrYWLgXK
CvnjacjRD0VNslcFqxBJG2Lly02Kc/MfwTDac/TMBd2shKQmiv7bSpA1gUEkm6SI
JfH6JnxZMrYfm49MiYaxzZ+FUkzt25hPpiHPxkKLzYRK00FJ8TK5U0HwHlQWSfIx
FnzEgMcY1LCYYVIEAbznPuwf8dUSEC0qC6giW6MreyADWwH/zFtWR3nQydIRp9ew
/HHeBG0y5u1ljox4OlUtguRsJCYxNCzxpd8Ur9R3s45alCvGQJgl0pvf/mh2JE4e
Sgei1yK/i3a9aOn/l7gEGtSJgfHVGGMmrFakJ4R+m/F4GWTiYLcbsRirxgNt9dLe
IuVuWSf/42SJ00MiznB5K8Wu7pMWB3jtp7+8nlGkEBrM7Lu+XRoYjGI0XjrwWijA
8/6MwCkYGzq6DG+W2Q0D6zNFQiUXVT870ZNooBmswaJEoukCPQRw3MRMQRQORg6Y
KHZuTFzVWqPznH8AJnsl6kWM6Wh3A/+9YniSB4lIrpq+fz0GnwQwbCOP5y+5ynMC
xnbNzi3aiYIpAspPkYGsA17M73m/dhqpoKxF407qGlakV2YfkxyYm/WkplO7u5GF
S7iXlop4Qd7uTq9e9S1TmSmZIu3VX0n71VW/dqyWpI7KpZUfx/tVamD/vrIa0+w1
QorljWc3NrKHT9V3p6eq0/3FT8tv0UEXoHsEiQmW/2vT6wqUMZq91HDU0wn64Iaj
4UeVuv5/lpR9nEXZs2BJR83xkHhYsB1LiSbTCR9mkb7ifTtG1z0FQRaQ/dkxVKWM
ihKy5whmkGWrNYfF2sN8GGCB1VGlSXHEG6b6wH4JXdad48vVxzI69VAjMekCkFbY
bA9HLJMrnoNIWwrZu7lr37k13F+BZ+kOgFCFZTyoFI1BE7N6k0qiX07EXRjIZWTI
RoG7/JNeosPP2cs6Fxww5ZM7HAh10TLbbZzNppPAa1Sm26qCQvXRjGMHD2aubkiu
iDDKbWjQKivg+J8tIZ49D7/KlKI8f7yehssWa5uX+vJaxEE1F8Z12F9hTrhu0Z9X
jN5NE4nMszyF3dasfnM9ni+nu1JXzMrBWB/Mh61dLXAmTqU3kaKOyefl84pDtHWB
6hKWMHRCALT4kj/X+V7gSohIX3b7IRZqInCu7sgLbKJU305w0hpcYdd5BxCNrEFF
QOfykcc1lZGJY6z4wc1TPKdj93kw4PW/WRBenIh/mX+QLoXfce0rZNcs22288TYh
nroW78fDjFqowYj4rWE8gNObfNizOA7/WRY0g+Sy3zr36IRv/iKbsw2FSsw/B7yQ
k+sydlVbFOcfD4u3wU5brtjpr0kuGXyWdArY2vT6akvO8bMUIc/ZlfNRksDwd7Y4
v04i0ERkts5b45T5CaazOxYdIOyt2cuabfB9oaXUZ/j5KGExWrH7WPKd+SfiwT77
CwJvWllnwMD/2QnqJU588iYZRlv+fpIyvG33n/22VV5hCSoQrhzb/VNWsM1llDv6
sWfPJJfBLJu3PvaKmVAfmwMXRDarZQH7B3gSm43JfW1AZrqxlpxoHwPOa34wO87M
BidfxpBccwNTGLLoMlRpw6JunbZlUJ7Pabv9H2/3mpGcZPkeg9rS47aOHXPN4aV1
flg4UpbkM+IdXSGna50k/KpNw74Frw7NY8jZgHcE29GWBQB8cG0NIPhtuCbjaqSE
wOxBBUr4w+tCSyQyUHKbehcTWqL3irWp/Adaet2PrylVT0Hy8YfD7D3STILeFzuw
KFLmK/U0Fu02GkUrn4cUHiWrk/tJXTUzGpis76aRKT3s1EVVqXKM/Hf3f4UGR5C4
ANo0dypNM3yV8ax52PFd6uxRG/aIGVxhhm9Ls9f+XiLd3pMGSAuX9A+9XLEKC9+Z
1bGdeorLNv2PBPYHOed87o+hRngwOq53xNGk9Yi4HJhtjncy5Ti06HzA1ve+xPZS
OXW9woXOj5yfoNoIy2GPXUAi0PoN5vj3UL1hN0fZB7thwwlo88emV62SirA3hgPs
SOOtBWEaZztuxmVa03EKzdAMr0pOY6Sp6ZsqU7rRnPdRUTulR9DBuBkR0Lh9SShh
wUV/IkNKJ65aTF4RR6rfjnM9T+O82ureKv5Ro5WwFa4Yz4NkVHF/57HXuVsba0oA
adcPfpM9/7/vOiH0Yejhm2TKGLZVzc4eXm0rZnDwcRgIW0athGpdQKYWXkW+IZ7K
iSbRKVfSxMrmwZgMBBescaPlxd7ongpvmCkTWlmK3dgm4oBv2TSIDmtnxlg4g+71
IQoSgc5GMBWYw4kxC5iZcSCqZvLSYCUH794QTgzT7URd8LozKZFeax/5S36YPXtP
FFV1FOyRbY4OhXLJ166DZ1d2fSKPXeg2peJRsVflm6J1OdnXqyG+69v/qWWU4vc/
jJR99mSMaKwEmEn9SuigqFZw+NMg4+17jZ5fkXRqUcH6YOaQSnb2kPa3b/2d1NZj
W3V5b9rCalR5BVIbvBNzKX0R8YfBdJTKgcH2t9ODKfzJNZpPY4TH99PIhaW+rEvm
YLtJb7y1RsfGmCaq95KrnUWKAjZD6e7LwqKJhlvTQEoKENg30DyDQ0R4AzTc+zyF
Bhm3o3wKfV/9sjP4oZXkuNG5gnEkk1zo1O02MfLH6YiC09AWc5HU+t8PHcXmJFv5
zckB3OpRqNknKzYXPNkQQ6JbvcWiLiTR7fHlEmv6P4uRcq8rpGYLwyX5iLuB3Cpw
uqUk32i+zF5LkCMeuous/eBQJ2NhqEBsu39i8CMYdfAW/X65HGoKr03D1kvjvPjY
LkxH4jD1UOpdM2JuCHAmKTlOMzcU5/3vhOZa1CdlZqsIB4T91h7oOfa5Z1nFoKLH
qPS9+uyzcFtXh/TYlvEmtgZEV31Hqm9aGpNKCoe52CPWVITP24e0AuPfD3AH2G/1
ANW48dNx8fU7c7fB6T+ZQnDcitneo2OfFbt+D8YWRhYTuk6+1XJ7ENurFheK5aZc
lpat489VLVt4ET3QUrmufgk4+DIPSSfrmQLkOckMulH6evhPAAcJxtSHQzu96e2X
XWeeYVZWYgljL3d1VeNGLlQQjCte8xajrfGxCSxhlHLoXMdMOMhbElePCrsiHziA
VKpwJYLOLXR6d3gzXqr6uF4lMJgmPXi4QmTXpsmyjKRAxcE6KPe2aPU08Is2ARo0
qN+T7bJp6p/SvU5mZqutrcAQ1iKYcRbn+F3qATGvbDuDWb1ejlaFOpWTWoGOM44R
dbG126I9xWorUQ7gL2kV6Ky8IyO2WJYSOfd4TXcpD5W5HRGbcFUrMCjyk+wSpAh2
mEBGr9OmUpKM/RG9tjc5dLSQPyMiEQP3c+7jSTwglMZd7e5Cl37WX+i5SiQsu0g3
9mWaYvZSsmYdFc44LZzzczGz06T8FWD3txuYYTH87u9py8ms/pkwmq/NQ1uTpML4
Vu0JGoQJegWx9a+5oBShO1rJjXuOtbmJeoN2lt4pQ3gUmyPkvWs3j7AbW03rmSKw
SKjCIyB70miyjFb5A7utS/BiSTZgyNMtRo2CvUV/4g2zczCBEL3qVM/aF49i/IEU
SlJIk6S0xQ/EV+vidrAmtSU3n9RRIYS1gGdj0aJX0LF/KqeUmbPTWaG83dAPnei8
v1a771WqBl5RxTaMrXcx9mO46STk+snEJVYG4Caiv5nO88m+hUbgvr+d0BLZFcBt
3xqhk3YgTGUrt49N55k/QQtkJO+QBuc4I7FlgFvX+HujINtnhY1vOpYDUMPF4kBs
NtM4b9snqC3u6A4X/yDgNx7niwXc7nw6e+ALKj6cH9R5tHLG5wNc2joM2AZmd4bl
U3/Muvz69hqbKxX/Hmu2Wp4CNw8YGNnrx819/u/bPU13M6wygE00xZr7GrjMlOuq
dspgTXqIVUYThW6hPbzqZNtpAelRq8sXA9pIBaAfX0WY/FcvkDOGm+5BpIUM1EHm
oGsTS5vnoxA2SljuamPpZLq9EB51CkwwtlV7aUtEPV2yFYQDrMwl6MlLMvt7Gksn
RR3ME+AoP573D2TTAAYBjwi4fSPmj650AcqHV98FInWdJTp0P3YHtqaCaI19EUyU
Wbc01jmalzAu6kyRbMWWu34xSWAhq25SG67TpP3rDoIyIEiCBmYOxB4qEz3rFVjp
QkI7jSmhb4B2uoXU4/vSsjS2pWErUtjyccLp7BYryYjRccEnXPkvkisG1qoDM9BF
l52HesB/WQuYLbU0tZzxH4ka3MNWsezTubK1Qn9USuNACgH/o1iexbN4kVtu6vPs
F6Vcx32CziHW7HT8a5Tfi20RMlTH/ia2Uhkof5ERG2T92V7I0hRuTpHH7WOcKnwb
zr3kmrZhazotAFfXsPtlKknxnmrIGsx8orBFhTUBbEWTX8zmFuJ5hbvCqnHTgLXE
DbeN5SyzzkpCkbAjS7wNtv2ebZ7Q+QCinTWbJOYxBXPj3qTwEN2eceETOEmuAyQn
fB7dxTZjsKDs0RbZeH+Zf6WOcqIa8XxvVxE7s02s0Y4/3jYndhDr1yEm8AdnQily
s+SHx0mAqPwZ5Q4XP7rjUan99AlW5ohhe+lfU6HqK6kVukDJEY/XJbIYahvyXHYb
oZlPQJkKC9D7dZ/rgtJdAX37r30ejgfmrgg8XGNC1sUYdOHx3+o/rXQgNzuQ2Tif
/A3xYtvYckbGP7u5dS6xRP48q1gQOR120zqZt0HLCti19inXrnh3sGp7WbtQrBNh
vmU/jzy2ulQdCpnaj/iCnTTiSKTaK5H4WV+phd7R+7bMIAHl76D8wmIIVugy7KLV
IfWAgNt1xFsc/PgfWNpP37NriOX2UDaiifBaN7ryaWvmX8SV6XJinhbV6Idtoty3
VFC2TOsBOUYlTnDvFhTEq/kF0MAJjlgALLL0dZ+AS2A1GbLMrOce6UY/aDXWnSAh
Iaa1aOGcLnQFPUFP0nAqkjK21MXhUg8XdFPoDm8FUWisLscOUcCzNstY95On5tNt
7t0FD8ZWKrhv/pyFZgTMMP8gyBKHC6zuEEr31IgDB806Bsn4pYrIrLKStQQRsqJx
AZtUuE6qI4JL+ZRXrCQ2AeOHS+Z4h+TB9UOtF/TvWfTJEZELp4TWJxMN7U363r99
eSrkovBHcQTO5Ejs6d+2yjebVfCF31ycjeCV9STQXMMiwiD/6TlxlYwkQK4imSv+
G4q2d2ohMTDHFJ2PipEfSxeE0kmjJJZuPZYIr/AaEHeTHTy+7ZRHBr2lEE3zP74I
mTek43ryIs/YVfcT9Ld1OCh/hBXXEOwg0jbAAii/vueS7rr9DhQIsROdzU425xCZ
KPvX7+O1Rrdl2v4huI79MNFJ4NC8GcSPX+Adn1/rPUOvTPl/4HWfbqlrpngyBIDP
5BVLGh3LbEyx3BTivn1ZSuRpbYJC0yDVlrog5NBCDK76/rg3/JpRWx+RyrrsrEwy
7TgYTmIhoAS311qfOpqkem4tTffkm9mC9tiuLQZ3sRXY0CggiIapFN4+BXKfTMZq
yBbfkU2kQW2q9Zmh7RzB/0aoKD7M8BevbJFaRa7UJcmXuTtu1PcTebkUsawLt13k
/foxW7Dvzr9a4V9lyrciik9PHDpGV72y58Z4sCsnXiPpabXZo50eZWnFcdZcbNgJ
EpYbD+l1HcCLVwjGjx7qBjWGLLcAQ6AyCOA+79KG2ibo1Bh+iYLqcDB712xdKcYs
NDoMosdbIkY+fAY40FiCbeWiN5p5yLJklsvrf2L6Us0pD+L9w+K8N0gE9frQwkw8
pZgNP81LoKbRmM1ArnWUcCwXcBua6JPHeBjNHdqZVRHbMvvJj9WwAdlCZ2wueASP
8/Ptrq8Alv3DsOW5Kn23L5CjG1Cu4fly2+DgkCbpGGf11NgrquTmgeHt6AakOsdy
GRd6JKUQywUMksiJ0gnQPF9vcvFIQ7XVEXaVIOc5W6F4jME40nIv1Z50T+Vyp2M3
wc8/gDPvAub+DbYrrXNaFd9rt6376X45IJBPqerdW+9NlV8pxusXN5gr2NuZOQqk
d0/+zqmrEzzkSvAScBX4YmpdmpLpr5X7M1cNYJc8Pyfgwxf2Ios0BahMszSGfmbj
K4XETVmbmfCxm+/Gky6ci46bwqUYhO48yYkf5nnSSjNEV3a9D3hG0Z+eQk0sAY0r
nlYM1cvJH5se70oNtyf0CS1guDF1IPsZBWW8Lw+3MYAtLdgi1Qxa81qLvDT8h7LC
y91XXhfQJr3Vs3DmfiXy2Ij12lHW5yzrh/sNUUqLvWSIabDgEwJk7ys5yztoJ2Xg
lrS/Sdgd8K33Ae0nS+jNgZ7YnN0XQ/SAIhqiXkXZeYRPnKWO1CZSyV5cbiRUp6bt
8OVB+3AfTWagH0pDsQP+OsoexeGD+kj7EtTD39l0XLffBPOzTUlFMb543nFkLwIM
xyCySMdl94AxJwaibrxE++aW3BiCLSMkkJyEUblNMGuWfwcXfchKf3P7YJojgwbZ
np83T+JBMdjsjk7mkInRE9Fm2UvoBITuukWpM9G/4F2Dv7YKpdx+QpCTAdDh4CaT
C7W4xOuOeF6y4iMgH8Sdvn/pyo9g7gBJHCaUN2599TnR0OCTkUzOmSuIjrsVP1VQ
nY59inj1KKiTOHuwPT7fRaOMMvc6D9HSGtb2KzC62atPzcuJa3iO0W9EXm3TGwV5
q8kUREgF2x+CgHb/WN+fgD8MKzDrkXCk3efzKp0iwkx4f8YDBGubpUDilkaFg6To
5u9M8iwldOd65MmedB85bBU38US0fl8QW4ZA7fQks5SJ9wbkXA6lA9m3GT+3TJX2
AREBW3PO5g724rPjo1oRq5fVdEWdv1s/epsJS83IpYT55iOGlCsvpe0cPs3cq0V0
rFz4HIVvg/p3zaVaZRjZR6P8i8L+2akE728hfT60zeM6kUZvWeMnPsSnq1OyXYXq
rG74ZENK4zX0YZV58tcvn+dAgNhYtVKsJsj3mgBjAubFetPDujXnl/wwUjxnPsFO
ntfkEqF2id9uueh6mathrphbVfzjb0CrRoZpi+meyZ4EWredAQhxhC8kXV1Pj+U+
2Z1xDNabq6Yl+e2/fpK/XZ5T4EBFSdtgrnAlUF5gbrBhWOTPAuNhZ1r1z1FrUUjd
bPeCr5m7m/dT5O6r/aMDkKPJnI+eN3d+/F41Sw1xBBVYgxk1N0zi8O7qqUOdQDEV
LKKq05oqxAi298whBDPGvOrflW7apEGZ/54a4nM5QbQCaUqQDS9CTrW4uU/rXOVh
FRvYtuQ2iM5G9Vks8Jw39YvDyu9trCwoQNTOQ2WxrBb7lmTLqOVIrsyfNI6TJuTE
/52frnAXvMPdKNBHn30r3Ogf7+DexCg2bInmpv7TRR7WoA38E6SkTMTw3rSxqeba
SKLzCdhScV8XtmKmcEd9t4aw0H06itRI5jURgxrF+CPL6QVegOBFiTLTFtqYYCxK
GiAAO65t0VS2GvWGXqWo7nzYKaCEaD4gygWms6FspZGP9u9EWmX/gnSgWbpT3j6Y
zqgIUxQpEWheVu8zkcULQZK7Smh22j8Xmd2eXDAORQ70+ni+TXDoGfnVi0PCIQJ0
BFP6oSWefmkvDcD4uhiYUIRSSN2IWDGv3d+XQOqqdo+4jXbMze6EM6Aytzx03PwT
ZG3/A0MY60eaeduhIOYXhQX1rAjqE3PNcFWfcLE8jZ4asKY6QVl0RWIX41oK5XoX
jEyItG8mlw7n4tVUgOTO++waIG+9pSNn69Ru+2SErHveq58joB+gIphIQT1t4orj
m2I07y+tdMgLsUZSbyyujkdqHRJ9LIkLc3QLYtUSGw1VmlsiRJ7XQ5uuoOgK9q9Q
U2SAX78Dn852kwJj3znPpO3O4O0ccPhZB8MasIgOf1f/3eH6zikX63LTxVwpVZD/
04jEzJ/xznXLH2iSnWFro89ko/fpQ5xlMwjmqPp38rT7kZNcUKA23ljIRGqdJcVD
SxxXv5VbFsJAqE8w2DnceZTQRGaITeCLTCIMDYKR7FU3VFHwi2SjLGxcy0Xf5Ej/
DiVRl/11Nu4IUoo5U5JFJYXl7+a71F4GJ+/UL14rMqRIHDhP8tEupI4YM68cmIAx
UAPtSCprfeCTKeYaXl76xE4Be719dAsXKrpsqKdhJJF9RD75dPdXlw3D7DyMTHOR
L+ftc8m5wJkVukaq4rhlY162N14RQBfEHpeJMmno2l5+UPZC2zHwzY/DqmV6b2HE
CsQclz1YipCdd6oGqcHw0WADtv1ljNliLAy7vl2QBdge5jxACltX1x+htGZYM0WB
RqX4sX2dI0HCCcD9mZNSLodPpTp4QK9XtylF/0nsouLWNtsqGnqEv8menKNFU0q6
RErCpSJNHvpToMtTQPnpcmn6Xxa5UG/nClpwHGXCestDiQgg/cU4DXESyuccLvx2
UC7wuZjqJXAxGQE/iRBi+pC2/WE7OXnKg1NmbfPPT5HSjnsgL6L8YJfxnpl4PnOZ
Vo5PHKpEnrGKml1vBHbTIYYXAV7qAav0x5mW1YeRmLVGE4ktCKUlZxwNY+B/OSMU
Lijb3hQNg+yKwKRN19lk0F/XRhYfvtqNNVkL+PlX/UddCIwHCIGWfYQLb9pqySTW
VgHftjhkk3MclEeqZweoY4O/ckYtJjF29u3ubypEZA3pp0fCELJXTeA+AfrBgAeX
ZBuwSGye7gqXoraNJ9RQkdCKnWTaVLAc16dxIxnoW11snAHX6OyhMkBlg22BzUwp
MO1v4T0ipYE008b0mjZMHWZN/Euxy85qGj0zoU46UzpgMVdxInim/1dKBr2LMOSu
8F3ht+GJhRnHRXiLX2Q+cuP1tsSc5hqOdVffwIQERVzl2J/iQWptm13MGXIbUlSx
H/yfI9UfRwvHOosN++hWiq454eDyAdjFX95tLvniNzTldhQRC8sbqc8NGYhCT5FU
yYdguGiWeqmu3go+a01mfP4k6R2oLDdoWBwnjwrwxUf1ubQfWgKytYC2xaihx2ct
LB4rgAHPvZ/redzslWNmLHco9ad4ytZzKnN+6HkBU2/xnsMK0hfAgiXmq6v5CT6r
0lA/xfYR7fvNxjoPr67n3ufrOgjeGPeMbd/0vfr5kRPMFTCwclZ5FfPlOp2/dWdC
RWjtVDR2QqguvrW23B7ikH6DoNB3/TQbx8575ZAjFd29voPi1q8a+X3Mv3hWPNkM
58Jqqz+nqZDVcVlGnOW4kC4X3B0XrqUZobaBpaxKDS577QqQI1Vey02WuWVROinb
MnFfGb6s9P1kqioOkA6z151oc8i8iffITdsfMJULGmQognamHcVU1NPANrduU9Xk
NLOcBI9tUF6Rs8uiseQyVfGfh7G957CmuzJodAXX54gBHjuC6tGE+MVyaEEQ2+qt
TgQuBqnc5leO/Z2CnmjJPyaTuFMZDKhu2zPzSxx0CZs7+SEcmCkO0gy4VoDQPNFq
uF0sDNWD7E2c5FyyZ3+5x7liW+KL+TTrWbyFovGx1VG0a/cEAR8l8QYLMkkq3Ye2
p1+s+3k5gwV5l4FLOr0bk99LxZz+OUttyME+jSHzBQ/thsnU0fxkK1iwaEbzWDtS
zELfKdfQUZmK1bAuJPmqKj9ZeOO1xC69fNnWOj4wObx8L+uaxzAGTxBtMvVJu2Ye
HuTrk0hQ6+KZXoiP/d9tYAmJnjYXzaTdeQhrY2blIQaKhjDZs61xO2PBMEZLIhTu
QHbsio0ttC8pDPi9u+az1mOfRBjiYCGvjG2R5fn70ot2dkxoLGq9bvClF9xbpnBB
G04fChdWhKZhWMEdXzAwYHoLBIFtWBEQP1R1dIikqlGUIhfqhfTRttEEqjQkDWWf
Xy/mPbuPkj67nypcSm0YqWJ8AI6DkTUVLCvVCMqiXiOv8Knx1up2U43N4WjuuesK
OhMGy1q4FBbBVg1pIfWCWAFnFjruCWc5MVlZB5Dwsoq6QjFEeLUspPjALifFE10G
ee51XvLv/LC805049t5+/T6rQhRkoAqzhLjveEtvBNsVRuDxs4AOTVF0/wuiTA+X
R3VQtDST91moq/hYnunjqvbpZx/XUmOkAgNCFFyyqtIJJl8t6ttuRBfMJgAQGe0B
jQzcPSeSF7L8Cp469tMccE/9fJQnsjuprl5Hsg+C8FwyJFRMLzbYkNp5oBQNLaTt
5bEH3acaknptFZKARXOmDANoC3ZOL0z7vb5oGCazeNWOubZh4jbohsUHSG+hQfPy
kOs5dq2VkI6XQuKnA3q83R5hGb3fsoI6fHIid5MN/kqcZ/aZI1eNwWZ90QNIbo64
xo9xfKTckzeqHa8vgPQfqQCa4ZO9f1VqcXV7tqIgxARBMG2drc+C94ZHU0patxNp
XMoGoWYpt89y/CyCM7UexUauMhkdZcJl3wLivhJ3muk90TPlpcHpsJxmJR7+xJ/N
i+S3EutBl0HnMFIN6wi0D/pmi3tAyP4DeTzbUE0dArISi+Fk5/LursDpxIv35nMz
bXfdMK8Nzl7ftN7uG1C6STUyB8moONjbuCnG0dGEam2dUqHeKoJNtROucSoHBzK/
GFkriSrq7Q6zAOkaFgPOUq/wuutTIt+AkNnAUoEPcl+cRsmrau/b6++jgMwgmfpQ
MUtx5ZjrY/VA0ArfvYkDcNxdg959XctZmqhKfy8J1JXDdsV0IyPsiGA5dNIhMFge
fZqfcV8CcdNNFykcai0gkDYhoyINT47tLhICoG4BTf3gw+uvHXAEixt5jNQmuSYW
am3+N7f53cdbZmrrBu3IIUFjMxLmFXRbh9rZpnxMC11n9MJp6stEIr1NF5Sw+XTv
2AC71slsi7Itkj61YpWHN7GvkMkQiE6ioZrdFYgmx8lvKldZai8FZiHMDwY6GF0H
7B9YfNSOSvipVhJd0RQgf1k0OrORz4bbhxWTF77D0aXAaHeP1iDHwSdPYo9r3EQY
9WF9H+xUD+Ji3gijCpe9pr8Nml91BOrjH6nlB93LUHb800TlvI8STdCVmW8nN4BY
H6aERuPd8moiqZq8opkd0i9TnLuueQsYZT3IxF7zsYemAAmKHNr56tiNffguTkqM
TI3hhxC6W1u7tx6/y5tq73+cjm9/ZViDCKRvmYwt78lA7il70y2HtqcQpjb1iRz+
Vc3i/CChr1vlfM4z1MLD9lyfm13EhoNJt6sQRGLzgPh+0XFpt3TQqnb5KeKqZCxn
3phr5/QZDIjmsNkSw8mag5rNBCZYt+O7RlaKAa9ms5Q+AIaNpbsn9QROHJjkrQs2
VV3QjxI2W+lUkHE370hyPb+k8evDCJa2HjUDr9N2i4ijD8PzdFWna9lNVFcjAz8l
AZWEB7GSk6fIVs+N9YwdBPeX6aTwk9iNDJgsBf7aajuQHhGCCcq455H+jd2+YN4k
6iY40LcP+tHto8yqbdmCU0YnhemU9DYw7VxzJ4bqujiO9hRQZzaFvxpPTxOnAOd6
0/SYRKbYS2jQfLhyrP/SbLuf8nE3fVzrhxaH/PHLL/tCAg1ZQeRMlnIYE10f81jq
Tio0w8ExdlPaxdYByr7COuhrxaO87y4JdHZ/AMHTy1uUO2nuAd0N7uD5MeObnXTM
zYxRg1lg8ogpOZAc+QQaHFhoca6XymgvATTY2XkAcKyquAGNiv1jPHBf1XV/3Soh
fOSwh2dgtGd6sVxJCavJKTe2BPO6PoK3D8JsS0rbsXxT3lH4rQi128W0TWhHAkXV
7mm6j8o7CS8cA1XNeKbuuJ5y7dP/ZTvtCjm69GuSJ1r3kDEz/0i5Z5f+0nAUmynY
wvpB+E9yb05Tv5IwTWQ3ou41mSbYQtI9kLvslz04B7TSXH2APku8/TSB6ibuya8h
y2Xr/Sxmd3K5St004/zOys5ahNGVf7n+2nRrcN1VTfWbPcJO0+LVZC4XLyqPrxB6
tYLQyog2Q4Tuaht4TV6h26JQlc07MpvnkiRB1W7HQFzX3wzt9n+xqN0ues9dhB+/
tHOvW8QQH3DyhAM1p3+jApXGeyRc7bwIp3WpdR9JZIwjLZtlR5p574b5MVJUrEyq
K5eajTwairYeYk0Xw2HImnKFM7JIhFxiOAL3ST5nEr+5AU9US3lfTMH6iFVe4OjZ
3FSD1B0MyqFh43c/Bmws2u6MX3rozNEejQXc5hprOR1vbhTJ1d81YVx2NJqkwqJA
GctKmc7KKAJgRtXjfY0Za/EJOnDsQHRt1QeBTaB2dLAedKrS8v/5vovGv1+z0zNY
6+2K16qMLS1NPSuEjJcUpImTNPUzNVqZBLyO5QQiL6t0tbh6IkXWAn43GK+i6001
00o6Xrs2m1cTA37nyftjP3iVkPG3a+qJiTx9GMfQAeVz9gllnP1H1j7zn7rGznI7
YteS2PijJXpeaMEA70i/B14a/wf8ZwCe+AKa+pkLd2dwxbzjciGL4+zdIrFdyM/r
zmtMuljhfyPIbJPxGtVOJBhNJ2k3q+Qoed4bRP7XmmG4sE26qiWPnHAmO0Jg217x
p+Uyr8C58XmUfMKFx/bJqDLbLen99jgq++eKorAhNfOoEU1lKBB1TMkwicVJuBda
V787V3lIGUzUu/U8jeYMfN5z/Hq4avcUvbAusmeNfgX+1uOZeh0J6A74czhNUCzo
sFxPnNkvAN+kTMFnFp2fE8n7MPNi/8bX7AA/0xKCOOSqeQWS27mvGMJFmk5AUMpL
WSh+/EbKx+MXy1UDujPOlxohOrCX7/ijegZToX2QdS9QwlafTqc2aLkBkIlZuNIQ
+87NdeTLjmUc/Qhq5uKmt71AJXnRWzfM9DUkWgDk66VH2beNIrQ5j6ey+W47Wrid
n8JJqSWWkstMGNQBIAijx5hJuo8nZmH1r+Z13b8B9R/KPuCBg/XgG8vn+CAjsAx9
9mofr4OJnA0DmlXUcbV0cU2olqZuJotiINQKFKlNFAcG5+akA2TNk+G/hJ7xb/Xw
NosFkko1b0vmwJrwVveuZFSaBoQVFh85hgX5flPI8cwgBumMqgnjVABCyy0h86Tq
nJlp0VJ2AAyjMYZ1tDzD7yJ7ma7566ruY9AmwNBS/numudcpR1jGr2MCzz6H/yEc
kPxMlBFPkJlu85E/KziyS3mc+auPmYQz2L4Tc8ICzv4QbDDmfkuyIIIX4jCfvrbB
BJmGm+/jJrUQXjVFngPXFvsxd7wSTE1KegyT3nlN1iSvdtzBx/Kp9PDrrFuQyw4m
o/oi9hn2lroJFmcL/RVZQO8Ot2D4FMuA2aGCogoSDZmN9k+Z3uBEBT+LB5Y+jW8y
4Df6YWEK8oi3pbiO8ZyyZmDl0y91Yfh2kMoViwkVfpby83YLWlmIPGF3mrtwy+uN
CTTuliV9mZoG8v4MQyxPmyUIWYo8b4REblLjOSKnEqIG1yIdSdO0NSpRXK/4Y1RV
LA7llhKSKqzCKJTUvyrMEwtWvc7KY4VgKzpQO9paYZNSx1hlswR2rn7a7V6GA3DP
Sk/RhSMyulEkd0HX2yqgewL5n0AQDxUUh4ipHRUkWIcLDz7lJfMjaV3djTwiVKcV
Na4XvBlMLvSlTFblKfHdzY52peghx1CB848QpI4HzzdK/edL6xoSDez7KGythNcA
Pffe+gOeNUh//ZxG9PUBbPfyophtYfsRrLFYPiR8fuaCCxm1vPKD9u0+bv73dInD
GVz7+Edk/0kFkDVaNutXN8c/HkdSTzcQgQtltzQ/ZqcA42JpfkAnCBgK0vJUmCct
RutqZtltSQTNJQicCGdqvtYWV7bhjbDcJsfhjeYj6PF936xGNV9Fi9mxBqBn9oQp
I16o+EIcl0VdnrN5pGflaTL/JdWiko2PQOuz8lv42N9zWAjEwpyJ+kS+5n4i2PLc
3SngUq/eXJ3eM2UBINm3gOnMm0S+X09WGPftMCO9jiFBr39JNP6hOKVNOnYqzUkm
xHaYG8toSFupUZKGLA7PettV1VnvQPICWv7AFEIJsKrLx3Dvb1JrraWxXBWiHV3q
KVE1AIVz17gBye6O0kok89/gJk6wQXt9Ozl8X6Ht9I/mNpJOMtBNGM7meH0o0vfx
/xPe44XxIFZ/D0LifjjT871rbINtIcEX4lBlrIVi+/WcLzHzw7zlplTzmtxh0KqY
sCWLITQPHi0PMUhTz/IPUPcGubej4CerpHP0ZFgPS8gR947D1J4Il9IE5XHPvTkC
tVmCJJa5ybB0aTZJbG0IqZHIFabFBTtd7UdEvah/xL3mWyRZHX9iFQrY4ZcYoE4C
oIKRHf3mUBuKe2ZnCs8XdHQ8HUUP03Yn62BE0y6eJO4s/Vt57lHuj28i4SIcAEIQ
i+vPm5cu62EI+2XjHEAip5yUljDD3qpN+eSDjo+FeTF1IzJGIArIX6NKHKoX3l/L
YsCMsowDjlvwymzomzeRCon+m7Z5VW9uQnFTFQ6D1P4XeW0vEF+PoAEeINcIYBIV
1JYhGX6/zuNOdJGgucMfgyxcfdWP1hUfVHJX4mIBb4XXmMoITZpCuzv4D6H3vJ0h
Z+7zh0ckO/8Pd5PnYgxvqUB1Mjgk9DUU4nP9c+ECU0yXterHiGEwlsPlsAYdeIVI
gKkvS2EWNS2H+vW8ILouxvnugH6nv1pp7AiNyH5wEW14AQMw8CyQqneObPyBdYPP
AregmIXkItHruZS/yY+GdDso4HE9Hj8khkj6LUvkO2MYBCTPsFPOUzKcf+kNfAiZ
7UumH+S60epmUdm6Wi8wPQM8ey+ED9ej3gc495EFLgvhf+4iWOudDfMNxenIm+XC
jNalA554RO0ccE9FPZpFlDH5bL43gIudVTsCjO25koRIl4PSRZZYKmfz5+tJMI5F
9yhH9VTXkOzSjF6G4nSe19dOFPlpI4Rmu6NsXkqrrb2Pf0GhmADg/+LU9o2gXSQG
PsZzAO+3HDXXC6UYas2qAOspqBJYXYb1ItpCBqIWAMV1qWZQW/Fz6V9xY8/834ej
jfRDHFdVeqBYMGGmEbYLBRDcLvei+qoenVtwHH8itbvQRRiyvIYhYO5ESI5hgoZS
GwsbZ8ebq+BlBwMttqsABZNVoMqqtsQlu2CozzFlGwTd/KSubBVm/dkK/CuFR8Fj
OUpfj55oSo+X+zij8FRHyn/ZMl2ITLo1St0y8fPGGmjcT7IXRCqmd5SYvdOIer9N
SoeJiyg7H8nY563ZKoiaKt64e+W7q/TqMIMUWiLSPjHpJi6KgYjP+316xqy1UkIj
iOY1twRU+mqzxGkHEVN7/oGiz0p8v1eQHslf8iHhgwZOffwvX1doolkx7HLSQuUp
36NymcMX03AqH+unBimoIz4aqjfawCgXem8+Dan1SAiOE4MeldA6R4sX4qiCL1FR
/IWfQs/62UE91rMvx1CrC46AVKF8n+sTATZfG11eVrk=
`protect END_PROTECTED
