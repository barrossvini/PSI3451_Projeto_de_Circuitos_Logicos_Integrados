`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v5Tj3HSIAYZor7miIxhg3HTdNyVKZ9prBH3S0Z1DHfE2grqdWcatxte5+T9JuGZ2
k6RfjZH0c+MxODf0mhdbKiKnnBrluQJJfZ8c0m40mrE3SawJPGF8V9bva/fGStK9
c5anfdvNQijyZHix734SOluWV3GJ3uELcK9N7Ro825e1qADlVRHDApkmy/jKJdnU
Apt/lqjeZXZAb6rZUdymjGRvbXUj5QCbfHAPi+GleiexBIYdT6US3Ua3QX1LiHq0
MX9i3RPVPhF1CHPk45aNyXgbalaC5zZG2aNjMDLMa0bjtXVZew7zZG0VSHNKT6gE
OkW57YegAtJ2DV6rdeb6j2VktB57ZdcYE1WvGpXjkqkRGTo5MEqlXT7KirlyEqEw
jbhKsi4C8S2l0itVy5kYI395zEXQj5/xkDegLRRSuN0RMwmCeolUvI0O3mwyqGZh
GfRq/MFhHbir047aMrR1Sca2/nMKhE06PL/v/XNuKgvAZH+XG48be0k9tPVRH0OW
8E19BgoF0pKS1xXhcXx3wjrYTvp0tN3XtmPLopK5F2Asjq8QmZwnL9ONY1Ymb3od
u0A/xHLKcsIL3jeRNnUeBuTg/sm7A6XGVO6wdd7BOiOCiFNZpjP8HZlsPnCtBcBr
HqUTuSZn9y0z8O91st1r7Y9QjPGVkCvMhDnaLLV5ZcMD+hD8E4fxQ11mml8tuQcP
`protect END_PROTECTED
