`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bcHqePcLVkxfNdNu0NVbeGHDhMc15FEDBwnndUCHywQngY6c55Z4L1tNvKhWGdam
+IVPFLsD1roKXVWnl8XmsBPDxxbJghW25I7DSW1dswsc7+JtLl/dzDBz6p/5K/k+
tf4tjxeszBbgwkvZRlb/+oesDHSsgnN9Fv9jfIZ0J4XTNRndyhAMgrBODuyJa8hn
yLM6BYNd4/7b1xn1OYEbQVb6B1YlOeNRPpwD57+ulPXKpYaN9lb8eTUA6T6Mh0/m
OYuT9pSp8el9wMs8luRtwTXQmeA80B9hf7EFwLnkXIGO+ucsySFYU/QLfiKo9SUO
0B9VO+TvBvXFzpGj6WLPqHPCvxXpsKcAin2yh6HQxPSnXp1pFTnojKSk7VI9sgX9
d0tZW2ekgta8ntFBo1fhfyYZm/W2EdDAx/6rKOMOjBMy2o1erG9xLXx/PNJBCAEv
TdM/OBxq0byuN+5U+l8Jk0R+iIr/UihlFsJRshnstX7zsaw1JYopZTFON3vOLIZx
Avayb5q4T2Urm5C2H4fVrU9D+xJPzXiFZcNp9in/+/Zo06iHQNdIQKcXsXMcwJGr
KW/PxIqYdUjAOdbHOa2UocZ4Xl8i53bgRrSHev353biopIqD0OWppGfXwlc3r4P3
VskkYh3BZuXiKzxtvRGVUBOu5Z4hZwiVHKjfTCywkuXqA0/fFEVDwXvOCN/jVGaz
1vmISP9PU0ntGN1mByviQ9Hp9G5x5jJBh1Eaveeyf/gVj8o2MJKGFhCQsxiNabKa
brwB4lAq6jzfWrFtQKCkyO8MNOC39ddaeJRoIq69y0OB2/j8uWVtmXEIyP0Eg4Vq
Oy2Uq6QRGuY6HmGJlfQFxcBp/8wdJwd/vZEfIUPUAbxaC7e2UyUkFEM/oWlwGVUs
dFa7vzciwPSDZVWS4aDh4d7vZYw36VMERyCnTVMy/TomDhpa5d7+WBv4aBldfEgi
TsuKFAYHTITRFBvf1XW51Sfo4YFsN5Z2rgq8J/Fd4KLi8T8jkg6XAMnzplsgpsSd
4Pea+0o0CFTCM52jvUrH2/gtKEXrFbomHq4KZjIY4r+TjAOd/jZYSUOlIElFfgLh
u5H+S1cks/DAItsXI6jadS4Kj81DKBEquJfHAeEi/hIIkAwww+bu2cukag2WbLSe
Egv1sFkFmM1YlsRCNGj1UdLNyii4wY5b6LehR2PlmRDF/aNhMpAz59QLdsRuZMpx
5iDiUp5gMkK3QXzuSHK38PmYiESBVMDs+3eqcc2K/rq5AHa9hSo7T+rKamLiFTPg
cw8Ki/ipTw4tl5tSGoIb0q4mRMsejMPosXx9LGXeFi6kI5TRCvZ8+nsDD5Vs9ugi
fk7A6P7uG85XnF6xXEF8I+2xegTF85MFADS5AUwzdRCaRf2tYe5Srp+KtM+7P245
BJhaQ+xy6aHps5ayi3dpOMQh7JldbFW5srQ6zkg4ciBAcFJgLlcic74rgBjBvSJk
UH66SX9UqLmkvbxV0JNMUZjBhoab1J3TzHEaJG3Va+WSlymCWaXl7sVAx4Cil4BA
XLqiZGP7ULNxBQ2kf+CScqUUQ/YBrehadoP6JLbR+iAwfkqXIJ4EB3ETRCKFNcpl
FMOjLIY0edi4dqAQ04BEx0FmHtjetnf+0IiaPznzuGfjt4i3D/mXbXeFC3ZFFlW9
E6P0zIKQerNCdRVD9FuIgq/KoOk1pfzJ0ru0sPUbv7IfqXIeEpohrQ5N2Dw7KLNJ
iD9es0PI2gLdGfX/j5ungke5DF06OMUe/3pvYWOsdU8V60Vcc+aeyOE/HCoaELG3
+Fug/zKTa7AoxLxGU9XYRPz4dCla9jWmekKGdtIZC2QJgurn5W1iXstkU/rCoUz0
a9HEkXGCSGPIzwdAWdFgeiZMILm7xStFh0Y+0mNBmLuUB4zKs8t673nYKMFbW6GE
VNvVBVKyfPBGy3ac90ZVdRKARlSe4zidN8m13GK3FbTF4OMzM9ZUs0fFC5+shIWv
WropoWb8gYlf3nIloQUtfu2DBEROH/kf3EdhnNfCMj4QnWbJyNfjEsU4rSS1ukiG
m5UhBWHcNBv79YwJoloMWPr0U0wIAkeWWMWs2VigLylxGWwM7MQW2KnPKuzykRfm
Qo5ZB1Rnc2p6UbyC9Zq/M+Dtqp5ow90QLTxkoSyl9R/ipkEBSLuhk6fNzAuoqjzD
F1E/ouyVrDHcgGtDXoMiW/qIely1n5NPg83sWDLdMqF7KgiMMpfMPgABPrzsXdQh
DyrH5VdVP9iQQ8i3DPIsOSFrbSdYwvW/BMvHLgPwAu1HG/XDGj3jkdiOW1wrMjzC
eDQJTqf4WTAAB83zkd+Oao/mM91dIpXD94O4JbW7LF7DS05Ck0be04RhGfCCUNsS
1631482VsYaXdw1gjl3RohzDqwxcdb/94dAiML3Pyo3DtVmIVhTnuAg8PlUG6/Xp
1/qgnAFkEHdHlSIE3S3gBWnPozjh0Jo7x3CZBovQnB5cyUS/1bbL2IWICzU52E8E
svideMUDbtnhMYrnNIsPGebIqjwIJgfqMrLdrv9AznUUCAJegRLVWw9VMQaLeXPc
6uqI/0VfQK7he59QIBys1auY2pFlBUYt/d/f6Pcf9T8SF5iv8qN1Jc7nGMH4NzEO
7CLS/cEhN2UWnKC2nq3eUwDAsNTFJ7cxtQdwKDwksx7G4PcjMFjXUtYOGkyrVEKj
OtGon+weTUY/RnBv0jKtZUFqPV1l6CkHy4Bywb7JLQm4TmXJrwNGT8ak+J2JkXDY
bTchyZ9U239q3hHrN32TOhrDmTYuWrUWjTRWhizaM7Pk5gwD1Jvoa1wboBqK+HC3
6W2zRvCXo8Y1cHm58A1lQSHRYfP23x1eNF678oyhHT4CmdBV/9BrwJioGSlnr4zQ
F3ddWYtUxFFBkXC2p24JKrRRf6Zz4/KY7tsCVwaJuTvhj78kfKV8Vd1NA588h1CK
DGx0QvoAQRsfHQW43EYKHAHTvjQLdTVTCJASbkjPzNq7hrw56U239a3dVNJpxGWy
9AaiNQ3sdTW8HA66NAVypgYvIimtNBrKBXdkWx6QdpKy9lZ5lo1tLuxLnrEfjFvE
AbOVYOj8UGU9sVC+bqKevPXxOuY7p7eJjI7nrXL+EUYu2Vq4dPSe1qK7aWVpPMnU
cvqqoy2lY1tZ9Kcn3yuXCOywnS4w4eSyL40YHf83p89UJ1E2nZXaYKQvEGs+HUlQ
8uqxypQKm3+EDLgAnIXaHvepAAZyoJsB3saUEAOdnLLqcucsTsgpGpWgc9V15tvS
7kW6vxlG+CtKnV45HVI55MsUG3VLaURljPXIHytApqtnnZv6SKjXskREYkq30W4v
+Yz124rhuhTC8yW1GslGQ/Dn67YlMmqIeVdJZi5sxkOtC85aob7yyFeKolMIHuan
rMUHmnBjUL7lz26cJNGeADU8Uiyydth4CGERN31R3IAXXS7IV+urkgsoW65R+kvl
KLXb3HqFq3mD1OUQJrwGyS8SDjMxlArOcBTQvqfQu5qVSQVvPmRPh6fvnHZAIKhC
2yanwYRXySoYMAXrfzNSBnhy74YUOsoazkjNUG0lg9PbCBPECsGCK2Qmm5FmC4kQ
EaIia1XeHJeoew3Cy3a6sd3+G6um7YMG2k3lTtitem2KPP/3tsTCvrC0eBbZosnk
AEwRQ9/L7BhJCnjOjT69GiF2qn4bCSsD9r80W8w0OgSLspv7tJCdz+SwKS1ARnsF
s6MmoyIwOYwc4xGzEvstTqltocwcwZQtrrZNT+wn83cQrQC+gRqoUB2FVPm3FQIT
+798Akot9F6zBM10hE42PrBCL/d6libTmxMGmyS/4CW06hy+4RiZe+ATVCKtp8kG
K7rqz3rAl6Ulxufnvxh/NCcEKawLAZLlCMX689+PMys1ARvaZnKbCOFAZadU1seC
y4A3PBRodCEhMDLC1cEAvA9uq55iM6+Nrte4cjWh6BgJEw/iCAsJs3aBld9cWAz1
B9Kudg6IzfuFrafspE5xeupAe7voGWF2s2xWcl0l54kZPgApa/V5GrN4j6tmjjG5
Iq0tVcXcpoaBTUCg2VVyX1WfzBDKmzvHTTD0Noy0EwEPXKsptgzB8JWsjsFNgN5U
LCGHiVpgn5V/eGiKG9c/i5Z5TatIxoGXI3Z2S2hmb1ebwRw9PmtIbkWsh/Ew6vjf
bQ0212bg09lMzcqmfvpbDqOPdKH5qeMkD8jlRslp0iXeRiePh3oyPzIvrybMZ+jw
ufDDQO7dv73C4h9hFFsp6+/cUkUQVkK8aBsJnMy2/Gk4mVlLAczDVcVAjj1N6+kc
5WK1p6Hs78VmRx4ZGx8LhCViO+2nQ6C/ZeyTSepFPWmdZhF3B3nntzya8p39rLGS
CLNgrU/wg6U8I4BuaEj/XTS9nFGNoOaFLovy+lR9hEYmu3JCWvz5KwiyG1IiNVfL
yjSFlGDL+hAN6xdqQqmftx6/va1hVoae3AzQg6TgOS6x0pQi/wZK2kDaCwaE6mEW
alyJZhBCzAgPXRyvqaVURScbvMmnPky7SYb+QtwhUBdZivupxeaIYbKaJNaKffgC
xi8tauJ87fML93zZgmON7YZRjzNQ5JBrefSN+xFkYY5hxo6HYB/kMUr+22vN2UIz
iC80Cpdv1K8+HkitQX9KPKu3DTMLXFyOSgAhtvGmkyRiJiY5bzfwsUEp+YSQMI4x
nkEmCaJVnuKjIytXmSAePt6HQRT2V/dpJyXpnRuVsNsKmdlsuiDBZzFL9Uqzk14S
2a9YZ6o+F43CjbMRYtP0bCoyQxjrb/NHLwY36I3z5GvV54N9RMCx1iClXEshE2W1
MYIw5O5IrTTfu3EFWVQYu5uA7spEqPJz3nHOI77K5a+lX9PaA4+gydcP6GJ9Nctn
oPtNKXcv1jmjmizO/d0OogFvjZdEOQJbJoAgjlZMCDhA3bU+xq19rjKbYkHxRYd4
9ehFRBY1KKZE7z98360FinONExOu+Jtm2145hhYlDiClBgc2wqcuXnKseVfFypnR
NFKRFTbzMydYMkhtRPZaMS2lj7p3OdhP9wIo4RWibwEU3CAvY5uHvPNciqRbfjLy
AbDVAvEmg4ENSey2S3NfPdOmB9z66g/mN4WpguhrRrjvEaZEcZRo67Ji+RsKqAqG
7ZaXnYcZmjWk2r5rWcGHanHdn2V7AAmKu9of0coPy+3t/q3XPGy9PjuqLfKxb5vm
9ca6SCRv89jm4le64ng0+QS1I/rDZibsWWTWphxCuaX4HZdPY6J5fWQyQEyk2A7b
djn+3ii6povSZ21ybBvL35kfWtBbtZfR0HIK0xevHGhVMzOaYxrxo5EHkETXJqrj
k2QSwR03/tHeOndFSE3CjFbNvWswg8wnonUIT7KUz2zCbcT0gE8hjxdqLg4E3IPs
+IkvuwgAaaB5SF0iBB81j+AL4+7xDuPuNEFtNm6nJAu/OIX7I6yHM76RMaZY8iSU
MTaGfDt2otfGuIUTuk2/847TOnhGhRd3GR5y+35Zo7g4zWckY+ETCDGBJcatiuNB
TTR4i1Gcw/lNCdK3JbODn3RTYPATOnLlld6tDO0pcMG1upuDUX5El5Tbi5RUddY2
EPGjkLRPN6WBg5zk69yZuCSJY1JbFCMtzOW98LfPMZmP7H0VEx37P3gZqHui2oEl
GM8KqjiLJ0MUyHEfpWNk0haHOpnPtjYBWYEXj5B6zQBxTlyZF7g7ZmPFBaEFjivX
oNtaiaZdzUj0MTfBAvndJ/X5hc+W9U//6AK2nw4ksiOlYixuCmdeky6vlKW2dLNe
Tmogan3syxQgzWbYs0cbd70JSI/UaL9408Fwf8pFR3+6zyGdJgO9hEq+9vZBSMxE
MA/8qsxTSYY1yTCYQIKglmnfB+0VlF9dOAEBDI3zoHNgluogyZ0OrxMQDNBokm+p
vB0XN0jxSDIrFD0T96a326gGa+8Y/9J211Ig2vS4VHsxHTn5c593nI0bLgs1Vhqn
mtO1pIqkz1QmW6T7OFlii0mYBso0HL9La/vjImFaTwDxouOLjegQpNRGLhuK/eg3
+4Loi4M36xz6UdO7C6gvVLOq9kkn+CBGqs4GvXLqdY+R0SYSOnlD/GLdIkfGULjy
UYAWeuc8i8Ub4hAsLRpZ8icjqksTOhFC7TWzbpjZ1B6IjDbZYDvLz8RnmMh/X7Mh
V01FZkktk6c4dQGricIAMhhFrBokzV6vcbBmsL1QBvro17tBRKO1N9r0Jz3289mZ
jM8xvgHHrGtK6lTZcevskfzMEmntjb0oTcTIqjbhlAMk1ryMaSl3lLVNY8qnpEhu
geKL1ouJl//92Xe9ce5jbXXJ05fg3sWF4mcMTezYJ5z2q5xXBubfB7dZoL7YXhSj
Qn3qxklpk5e2XntWTqUqElZLUzjet9fJaqmFQ9UlCbaZpwi3sjXyc6fyTpZunmeO
cer7g6RIizvMuBWj4SLV34TEjKzJU02mz5O+FayGqx6dtE+1WRJ9xWgUJuP9gYjz
kloIYoQDxI0MnhDaiW7YJ1x1MKHAT4zvfGEQfqxeULiqd6HQLpQE8nrof2nuBpwS
rkcTHqozoNgQUidvXQvOJ1o5XPM2WEMwOJ/7mAonQWjgjDzpNzIuq8s5FFw8/NgE
9q5dIZFTcez0cyOhPMl+9lhkgBP4VEPuqrEbfz+CAQoBE5o+QA2fS6RpK/Fg7eAK
AwWTWTIj/HzSp7451e1/F3QPumo8Cx+s1N4Bbt1aGlNPXLX4G/DPSyvgGEXTlQLh
8bKI17ihasq/dp855rccxecSik9iU8LF9a4hawvM32dAqXQqG7Jt5dZsdv+2HDNe
EhmTfiexDNUHXZoqXTAPNJcNirJV4IGpzva791E8+GblYakvyZmP86xa3iut8Hqu
7yOBlDtDiIeYZEg0dOmtdFk7dG/wQp5e/QKRH+xLNorezAJBJzYdnSozPs4ZBiHi
9XfCKzVhLkShyP8Fc0h71bsB6JWWvkG4JO0B8iGoIMUXGHgBoZAFqRdFlD36T2hC
wMPyWL0u66VnuJ31iOWsscC66auvHqZ3IB41ygfU8LCn2zb9rjOKN3eQwIgd2MP+
W4leP8dmBsst7DLsQp6z/E5wttWGAlywXZYksBYtWfm5S7XlwZtAK+BvkA1uuT5g
jTKqqXTCCO62C/KhFm4A1fP7MzByJLTqIzYYT0H+bzZU+syCt3JQS6OQkc659FPc
2+V2RWItjXryYkKyXqjF7RpwRo7JR78KOl3SURtz6Kp/CAkhwl1T3u949/SLLiZu
ucXCn3ccg0LmEH3CQ8yCUtQdFqM2RTybo7Lf0uSnv0jjX4/F1/gTbUeEVp3el9CX
h4oDfxa+pNlD9t6e7jMvDUWqsiYuJ/w6Uk2+7PYCITRGe2R2Za7Xc6xojqhiv7aT
FOgRF6ASa5YJA4cAHx13/pDjtEpFeVgTUk/DST4BjfLq1dY3r4Jr3JXusH5KXNaR
3hCaX1iS+Mo2zJ44MT8rQBuJ58uKkDn9aE3LjRxYegJ5/Z04YbzH2oIuv5zKN0JD
xhWHrYpveEMuytsvtVYlOd1i7RIkPQlrsZUPVj7ey9Vr2rcRk+a1wq+PlcycVHIv
sQ1elGhiaZoghwbOFALkNAOaA5TvJV/ZblaKz7a9i2HSrIj5zkJYz5PomlrR6NPr
pAHliW4atr14VuYWVj0q/nRmQpfkZPA7U6K1p9l8mt23/vA3acIxBAHyVmKng+1n
NQVyJhnd+e3ABTYHNbOTNJ4a3+LL1VlWxEh14/IPnQZ0yFHZRsMlbfWJ6Ws/YEB3
53MB0GhGi1FbF6E5w3d/Daxgmu0MgY0xuxpCPmJcxywIY2Gzkxa18lUKqIA1y7ua
+XYFfdyEmXdgTfQMdBgV8FENFgSX87acpZPTRDiVu6dID6/DQfBs8hFDRbEs28yI
BIMMjpaOs9ATK7Iz4nXmEK0VqspjDjr1v5fzKQwCAwUVg1hb92WRjMBIzSIO7chr
NtC3yEvZahsdUrmoRLRFZ11Wvtc72lgiD6uDMSPS7x+otJWLAI+scLZG/YheAsnh
Wj8wC5VC9m6xDCX0+Tfu9rGRJEOrA77DnFf5XoZYaX/OeEMZwZyjOPUura8I6asC
opnsCxfXxFu9KT+na9oeLfunUlEGAgd79fTf3RRn7QVP655FDHHApHApJ6D/FM0L
xzeTdVOh0tMXPSaIJIH27l5aKL2r8TQ56kh0NWNb8Aen59Opcmeg7eneHh1qmsmp
Mx+OSj0bci/Sp/Njwjw/ICYLVnD3ZAXeCF+76isDuOMf2ZhgqKoI44keQPYEsIgC
nfOrr7tsQG9Rqh8PpxaUkKWrxIrBT9pS1oAjAn6SRbHxC1Y9qmCyKMNiMwVFBDX8
ehmUDkM2US56OlStgaLLvSi1pRCM0IPGZdAFT2tX+FKreBfU6Jkjv19M+oY2gJkH
nOiRj3hpA7seq2BRO6FyzZytrsd2DSshEizTRuTeFyR5KbGuiY0SUejpe+TAmKDw
vsj0QdIyGz2rvIaHXV12xeFTLVTSVgP+hW1pBCvwW+ZTzPEfw8VURvRB+uDZu6Wr
QVpDO6Q7Q2hEcj5A8bznb1UsV5RsL/eXX87OfR78ymYQoJhxi/Rg8Oa1xKybSAul
OIemFBLmkPceM/K7wAn6nSliusVBVbSVUzyi87oRT8eUke5PCoOpqmozBj3sit3t
lzYJOu+w/WuKptMMwhkfcE4OvA6eAe869cfMV6+n7pRP+9KJ94tNvm0sE0Qe3mEI
6QCXjugdt/sDKkSHgg+QO9tx09DiD+s5jUbhuYNCAhHHgHJoa4ATbjY6ZecC1Zmb
uukgSbi1llypFkBkbvV4KArPbP5ZZxcJbJMVH3rhbrOKcAM0f/2w4W73wP7BqkT7
pF00m2pM5ggY1b8mgz7shFVXeLAjsDZUThZQHftkay1MZ35HjsWt+k7ZAWeq/FPm
4htRlDqxkEi53HYCYUrXe87/xeUsGANb4vgey8OnRmtm8xmniABYJGIlKzgmgW7H
LjO9GIiioacAxbIFI2kjhfCwGtPglzcJ61dVpDuMsf2Cu4Jdi4wQEhL5jp+T1MvS
ZhSibKhiuWY22xAA0XUF18J6QFuW3lSfBL/R7C8IfLKuAmX7GYohQ2aL/CNWWLuY
qomwfHtfv/gSjeuOylOOIGwVFLM2vvI2ebDYlTwZt5vOa7H2XyLEdirYsEsuull8
iOrUYZHhOyBYGhvBHiwh+wKEns+YxRwHaUzv0tb7F2rXszZKP2ujQazHQWX06O4I
9nObz0aq7ICrUGkcgUc8lOPTt9j58YDpr1O7JZyEpNnHBAOSuU1awvISTy9F5fg2
RxbvnIdCEAzRp1MqqspRF5Xyoq8J1v9wcRkO/jJSgVT15t+kqHYKvdIC2yEq0PCx
OWj4hmBQk0xYoyZEz7w99GZxI5B6T1cneqI3xMo7eaFliWH5kXIAHDlSKoeOk9xE
h4iKL1TDrwd5XaB/Asq2cYXFNrgVT3Wq2dqYkSFcjZSwnCkLNtFVieH9u1+OtgXR
ymDxQV0I4eUxFxI1mZvPTmGXh3+F2Y/Z93TJiqEOQntjY+qAmorPz5qu4EKRVxr0
Nc9+8+f688Lnf7wtEosCnCdkzM/QBlfa9xudZlpS0OWqKlfl8AANeqkMO/L1ID7M
J89xqFDszA78r2z7vjnXGlUaRZJhz4H83UjpSzcFQwMvzjEf7NMv04orguQHfkh0
XyX61WfjvDeM9ArDsVsN8fXtNMaiFC70/EyLo4A27XcUo7PR3V0aZ+uZaewkwrff
3YRrYy2DJrzGE3tmDMA643kwrOTKzITpXGt/4zCHrzdxeYdFFep7QSH4mWWFHAVi
1bfi7ALr06f1kMLc04xqYF2IXnqsdek3gQlmcT6QvChQbLaucg1SCgU+Avl9coKg
SXIbUe4/QqIvvbTAbuqpABuBG97jCt9ZB2iFuZIFsZed4Lkf1SURLnvMgmFGjgBg
U0kVT/bvl2tV0D1DhHcrH0PfkiMVOIrR0xqefG8V/R2dmF3zehk5KZOAzNHctGuu
OPVwB0To7qFAvEM098C4HIbbAJE2h8bb1Wofo63rawsYKnHdcRhauxq5EYwByPom
8Q28A5un+in+DNcO++A6ytlKH/TS4UBoAZPY8lB6SvXXauzIZeKp0d8Mmtk0CxLD
QA2CWmiCQlxFNvGjtjkcDkRQrFkBmDXW7fEc8CpgqOlz2H2yaoH8E6tjUQmZDYTe
zouKSLC0cvCHzkUFDvSjDoXKQmzY/VHXkFZ14cBnQ0cyORHcXYnwb7+QJ6aCK/XK
aIlPiOkwUnsoKBE8KTbWlyvUzLwEVB1o5ET6JyMoVsFy8phtg58AdW69RQG4FZk9
Adi/5XzQNPFd3fuxoUTH83TKyoUB07RrHp+a7Q5CAteWt3KPiQVF6H5SOh8vYfmY
RBLSfkcd1hhAgDXoVTxvs40xQpRYP5iBVtl2FiGdDo+s8NnSdkgPf8M8RU8cYCE4
4YGqu35aRRg4N7V0vluvyORPYYr4BftixH1SEWMmqnx+9FhSZpbhMAe6FOK94Byc
QGWrcSw3HiHiUvTwrRyntW9INCgyrzXgeNWG/4JQM9mS6PUliV7iX4AzI9pUsyHR
/bY0NE7H0bBkSeThwqKaMfJq6nai1hVMKlWmeLGn3XekjlBAE1gTFdVlruG3qwzY
vwIAX0KW+1N6bhD0MOsB5BW+5ZfLk9DcwP9v6iKJPXBVS3d69gzG+5wl8Hg0DmmR
wbv4h/mZIEO+/eo8qtlRlVqQHTi54pNdnuOkMVQEGJW8AUWJFcHHfM7rnyoxnkBp
3v47GIZy0hxUpzwpbaTvXHVJGdod1zjmGQRctHkIv3lPUB2Oc5fvg9SHa+/xqbgK
TAujtCttLapXds0A8TL8GvyUWUKZEn3b23hQionBN4mY2yZs7K3BS16FKH9gzmGG
X/h+8P8WgVu9E5KdLpFYQ8Axpo+HUcOsAjZXz91uWPRDX8x/UwDjfK2Nc1U1yGaJ
mNRX9ZA7t05mKD1ARaCl8Bf+h+p/SNQab9sJgU/xW8d1HSnKLonz10BJlRvx3IIS
puzME7jYUwZ1RKFpVzS6phqC7b5D7z54/t7l38uEfY0afAMLcvxuORXHAph1ej04
OzvT6Cc8l+ur8jY6D/Dr3/r9ADpKK5XTo+xw+0e6tbT426MiqPHBQB6Dr0NqulVJ
QEjOAq6NQn/7lH2D9rY77bEn/JwN+YUmo8hgqP1QGkvGzdvGSfbjgrZ6PcaopwHJ
DROA4e5BPMXEwn3wSJKc240WjluxL7vYIGSuRvFsZxF0wvLuPUKpZyB2Nf/0O5kS
cyYr67VgGwpvgFxzhVcOwxiv0XQ0vphfaHREDZMlUf/QrqWhyXphs3RAgbD8p8pf
NG+RMizVkdCOdYqw4owlAUAw2mRRmukF4VrZNjmjPWhR0FH96wMO7v0VHr7MN+DP
1ozslF8q3NUWUhm1KW45oiQu3kwZKos04mXWOzLcv/LwgDwSmytzfQevr38nUVU4
i68v3gYo5s9xSRBWoIJGQhdo73d1j0iXn06o039Dv+DOfGWbDhzjlAEau9l36Obg
uShjl9dK82QqMa7J+GBiXjG3b+R7RmpkOFDFHpFsPTlsfa6cw8Iy9uSt36e6SUos
4oOu4KfpMcd/qJQvU0C/M3hxyQcsZsfnwVCWIM1dQcsLhJ4JsZiWFbp5Schc2UBY
vla+H5FdoW36hURaPznPXOS0d/wD6zgT5RwADp2+NfVjUGM774gDrtZDMS7N0Org
fG+2C7nAYORwcSObCt7NIPPly9ERjgcNoD80QuGayxBiRP2ryFtxm3J5DMjL2PSj
0nlp+glp21K1I6plFi0SZF2yEtuVuix+8bP8p35ISpvuGTcyV9/mmyKlt1y3SkCS
we9SaInYBeOSrxFucCNAt1aj5CWQBk9JCwTpPO0yo34eIZ46MW/84+BsALkeIsxE
SWv1uGTGChZ0ZQBTBOhZVeXB8+WSeH9Td3ayILioNgMGk66iIdYEjVj+GCSABP+v
FOKOTb0NGtGG5MFzFAZhDz6m/dyw/L8HQGDh6kMz0+rdYaXMUSwH3NHMi2F3Q+FP
Y6nELe2/cBUCbq1ELoVMqi9WU5HDf9JI3x/UClMKkGTCtVllY/5xI4pPapckin+P
6ShEO8u34UNGatpnu24l3TjHck/9HncvIX1OpJbeS3jcF4C+xbHVI+yyUmgqKX+f
0+5gnNYEMxSMQ90+sRTnSbkXlxrQ/Ri/nM53+hYH85CUKkyjcXQfy8dckCLk2OqP
VQc4i9P86lcF2r4iyd+su0n0leLvKjWE0F7UOBcJEknic1trQq4VDBzPF/PKbrwA
B5qZ0Kwz5oaQPqkN83k3NQGC3zuTX1Lf5n2qa/dOV2mD8Q0cjH1s+3y9aQ+RSx9n
jXQOScPqhrZ1Wz6VqETorJucg8zDzpGcYyuYeLLw9c6gfUD0jKnt+Itzv7bds3kL
KHddBGelaJmMBLxk/TGx0U3ymn3JLTgmxtig6AXDp1L1JTl9Mjj0MB1RZFk5mdDA
qzuLGvqOMfrH3ZVazG4POeJrZlLnJJNr/G3hswCrD0p+/S0lTAA5a/vfsa6em2Ec
0oa2JaD4tXhcDE0LfE8Ju27gCXEJSZpxHm/I7zNOPRa0sFMeqEIoylYc587in3uf
BNI1M2hrEaZc7jhEnvFkjKzggfrJREWdIYJvRfBsWB9sQvD6W9tUdl1EjFCVd/F+
RGmwKS4hQmZAbMo9Z/54PxprCojCSypIXLl5KmlD+AALVGkTY0iE7BeVDrhtZi23
DJ7SMaFDkLJVe6V1bGohhnTqwM4yfy2BPSJi/VxiGuiVggu1P6dnx9Wf9zq1bL9A
27sDuY89XY9z6bY3icrjpNOkfRE0kdMlhjLYyV1qC1DN9ebWkSBKMTkXIp1lhEIE
/6rOONnAHsr1/hOyHF/P9DpHwAl7sX7ymZC0nctZCxZAAWkrSAk5+omtBkNSQvwZ
H4GYRjLImR1TfDV/O5ZNhhExAtjJlh/XItVtqP1OPVFchNtNxtHmF8fotCE5dCx2
Zm6/CsyMIrZEtvQPuFG0On/ea6tLBiEt8StH6aAxaQhwwW6VpiIKC9DVvNMpKrFk
G/vf+QpDUYHw+vLLLjqilYYdF/ChUWLBzt17ncs5zgJlGdnu5FQpwNrkc4hhcOus
XF3o/6UY2Yr/HMgDeXFOuHFti5s1EEI8edG3uusrUP/XcJhIcGBU14BiKT/ydYU8
dcXOuqnWPbsI73HiM9tiEeNC9bVAup/KRxqHTdxXcjqq9t+Xi942Au0zfuw8rmTO
`protect END_PROTECTED
