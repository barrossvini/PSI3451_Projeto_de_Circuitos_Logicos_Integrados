`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ET0cUaEOW9+FTptHNdoN7yKF5wDokxQVjIR/2xA8YrjGWVBlA0ArTVL0iJn25wxB
vHGcM2Hs61fyewxnKpHAFwMKKN0zhr37Sk7qhbMt3UMVhZvWGor+EwR8KgZzPb3y
y2hLMXNHoTg5CMn0daYTvvJ+mXK+sjX8yfVAv1cADee++Jui2GLgBgNcL7SQ/C0U
LBeeGaXeqyRUQEwXZCTdI1IUnmL+O4TG+lTsdJY8QNiSn3sbd4oRXr+FqrICsC+H
PwswdcNwBPbHsE79bVtuDo5nmtVCMniMpT7jSmdbP+Ldj5EsjICzLtGWtUS0B6P0
38sfMw5G+B2EG1gFv+1zPyFQ4B1RBmF1trPtqP/Pdk1kHXjXAk+IIMXR1/aCYBEF
2Hmd9YZBt443d5Q76Z0MPQ5wXnBProVMEgdOA8NL4y35Km9lgdV2h5Zg6j+LDK5u
P49K3wXfV5XDx/OS3SmkKD1Kb0/BTSJ4RQrKm9NkT8aiZzgg9uTF3iPWJrtd+bAd
QvdqRYTYO/udYHf9cWcxSbSpB09xN7PDP1tOGTMOd5J1ui55pY+GQLxTGmcginn1
ocrjP30Bg8wYWn0dDn864F7DemsTS7BAb1A9xaPrf0RMmbAnw7jzWtu38oUKSfHk
2wOv7Z9Wa1MGMDKuT6Ox4h1g1xAwy6XXzdV9mmbmQBDjTQqU+MZlPJWWOn5sJC+W
YbvEnJXOXHVFSVi8aJO00vZ4C9eyMVkJgEC0vuszY4DsuenvQ+Jb7Puwk4HEDKaR
8aCPGojS0mmXrODgADwsa2PEsIruVGKE58vfP/2hmwtpmpsfWhx+Gc6k21285jTv
uLj72W6h0wO4/Lm+345ea00THYNzv5odXah7fl/OuGY1h8+ThPNVSNx2rzLXiNOc
MhUb+7NRoX7+vCuZZNVPAkS018FP8ov9CxDfci12Pg/fce3VZ7kakoOZqmAZEpYP
lVPtE2eDXZ1/nR4TqcB2Xrm8xJH9EuCnBpmF9stR38YUI7rm+bFWn2H4QsZz9YBG
xMBtwu1tteM56CMTETE8zcNGHiFyQkdU18aEy/ZgqfY5wI81S96f1W25TrS4b8p5
B1iJQjkNUVqc3ORFXuC8oJqmalSZuxGmAn6aHK2HteR97bOpEqQKGzk0ZQzLw/wv
0IcvkjX05FlS/DDzUF+JaP7AMBZmNKcedx42KS1mqNUmS2NfUX58BkUvUlASdZ2o
ySfWlla+33OgsDVXdLijtpw2XpzJVOzG98UaBW34fp0Ooxp2ZHPnPba1zhdyJN9Y
sYlOLTd4JEv5Ds+p9pmi5p/JmyOStapLfEk1ulZcaot8P70dxjU899riA4LJRkS9
q3wGxToYPJ/EeZpB/C43zaLKYqXvXYJAsuTUCKqXJYUTYnsqsnV3GbDels78ay2z
c/VsxUBJZ26jUNYelVcOCDmrzUT/8GxJhV373NNDvtsvDKAGTT+JMKRfxBLfi24C
f/6yXwKQ+OaSL5MhR4rP5srTIKad+n+RbKYwPEcPozHVyUBYcE8yvryX1kWsBq22
CLlGTEjoIylUa3zfLzYxHT73SjEHjvX7lQtx6hE/Pj5KZ0Nwm0cwa3/DhJDgdLEY
wOyzn39KKGBmeZPXWscObotD/yE0tyBjSAMeVyeaAw6qTEkw8HzimjKQ4JaxnqSk
LwsCW2EP/s94INdpGxTSerKY+iSouGf5/WRniZgqnmsDf9kXmbqnYafkwb+Eq16F
bcqt8R2/B/LUOPnquYtwyKfQkoPKwUTWa5l6r1eNLyVz+aW22tnKD+gF4EakCQNN
pxL1aP9sIpfkSYwFIMTrR10/fqEQ7Y2jLbEBO/duj19+UfyQ+TjaXukq0EUN3ngf
Win2/h8j5XFLQY5EFWxQFXbysIHD7R6iayZ2w5usSxvCMhl0z+9TEqfGoWDecaNU
XDtUdaza6eECV7JB2e+PBNevSvTVVyYvnfYSro29Qi+qAIs2DU0PcNfuDxQX5H6+
E9mVrGwVKAGzIaho/Mpg5zmN068k1QAtaiw7+MNvGx8K5PiN9nfj6mhGgG85p05f
vMyVW/QyVpGO2/hXlVvisMKIMWGlmxOmAtA2tKhce58E0MxHyda/XPJAz06Bd9XH
Xw1yOfcViTF2CXRu1hXvFqP/yZaeIYoU/w8/w6GMLOiav2gsLU4vj3ljlJrzCoNh
/5qtuKzm8kjZZYsw9QBXpmSbaofm0ZDULRmlHWrtZMkRT1CMbfPb0Xe/f7QCbNRj
RO2UKcbmPv3Hf4Ny7KdDu9DDV7rA6MQIxDnreUGnyHv/r9/NkuD3RmG1HCI8mKMv
WHLTc9os0XVOwuGlUSvNteG6ZH0ySWNMcRcquZv+SrNxcHFN+FJgjlIIHMToNMAP
6TO5LJmfAlKm4naMV8MNeWoTlqbVf+nfyTHHZWFZz6kD6NeP34Qpr6cvtGwaVasA
GfcY4s/HL1Se7i070JuwJVpNBWkv+92XmtTXKHv+eApdfvU07UUyFHHdMTms/Hff
OoyTW/8PfCgKT5h3ENNgQE96HGzCDT9V36jQ9wgrg6thXYb+6NcWB31/nzFSUV/V
mdJ5Kjg/TCD7cwt/MfDssTJf3sSCdgAi15QDa0+9Ahd5elme7fcjCK/qkTt9HpGX
3qkhvllJy2N7OhYsCh/C+lquaod5QHznqnkD/Y2q0rIi3r9azPr9II0J+RXsmdyV
CRrhaL80UvIHrUBA8PBLX28DTGJvTauWxBQZrYd7ltv3PvmMce9jucVEENb5Y0aA
n9Dz6ikzEFRHb2zCo524yYT47hZjFI2VSFzCfV5JhzxJIqN7Z57TjtGWm1cM0Hs0
rtDFa5uGbW+RN0S8KTgPml3gt+Sd+4p+QH43ClkEMTT8QRMFaoyUI3ysF3tSprhk
2EujJl73KZPkU1S2JhIzMxbfKHE5N4/02x31mYqKiN6ODwTIU3Iv27JU9KTjSUrG
b431u8+hOQlj5NL17ianCAQxOxBNQpz7yXc2Fl9T9YI50z5mBaa9icOZ0gSMsc8o
ml8NYmGwIqCTj2H7hunU3gvoN3ONCBPMG0qgkl7O7MREI7CSAIiorobEb21EYzDZ
S2gE5rEavfo/xakTX1rimujrwn85bWEbQZwHoMa5tnbzRZkNBc0WmqPBJrm8Av2F
UQNdViKxkcZiRBy3tJyYMqoZ7kPtgBcqiTYaqWF35WiXcGGJ0IvHJZTHKGpybE8x
mG/jy2ikfDGQySg+cZmxCHRvIRjqlrdvE/QW5ShaR11XSnJOZoObTIVDvS9lobzP
lcf/YeU6uD9QAzBpLQE7mjnLFE94RelFTHHIrx/2RNCgukgmDUyNv9JpQbgv8USR
U1gLJP74D+/9M2P8z7LqFjFqUIbCNsNDaKWfXXQmdkBoJWoXM5T44/lt2nNkB2yX
gSpoB+nA2EKERupzb3wTDcL06ebvE9RUmWoiXKVSCZWXZyRVcy4B/MY/9QOYUgTm
1MHaZJoY++W/QKWfLZkGqFhOveFgrKrtZR6aHXI0Flm9byxsi9ClJxzOGa7QcwkI
GQSb7ZrrLN9r2JGLkDG+GjkBZFrqzq4Bv6gnrDnUJGBi8ua33O8sg3gZvfpDtuRk
pRMDXA9C9Qx7CllnzcNFbIuQE4uIPzTobqPqc28qM3oX/Bjr0QhlwaAujl1i1Mq4
RSvMFtbyAfNJe5oAaEL1F/Kcib89OAobqPrGtEDl0eQakc4MhB4h6IwD6bhlg5Kw
dEX/R2iUj4hovenHM7ui/uH6jNxHq+CN2wbRudzoAxz9mPxxjQMybiu0h+5E2I8W
tLH3gJ1jYqT1aJsJkCG7B08I54Optu9bA0kbg7Goh77hWOW+yhrBwGqOooe8V36t
oVJ0KH/9jRB+FDOuQHM9Z0HQK7rneghVzpOOcEJ06Uz/vo5mzvVxiMqmup5SeN6d
pG+Zu+AIcox0HEB8SjkR6ygDyWjPubuiH8bVub8MtU3afm35cbgGbCInSEbdZI3V
AINr41LvxeGYhPGoXYcozAmrfTcrxsYyMKshBHrtC+82IvTZTqT566w1DkgDVrCg
jnpmdtPkzX6FnGD/dRy9QXunyiMdg6EXx/bJmyTx3soPOV/Z5zb2Cu3XbmIZ2+Ff
7ntDcUc7vvs4/XbmLPqFkMv+Rc/GfUHdgY+UuOCYU948thHwlfwSo8jTf3z1n9mt
RDYPcZ91nJYu7oWwgoyssDgZRPKZ7LenX+JqpXYbctY/YLMDeKK8gJAu9vV6qzhX
kYZ/HRnlBnIIewTSENvpwPUhzJib1cSxz1d3hEln7DsTnevEMA3+uOqFDtlP1QHP
c2/yUVVYiq2uNLh0bP7kFRZByCqrUW/xmz8nhUfT1y5GHZFzYvv+KTlCzkL2EWem
qLSfqC8i1//B25wiCboxiBpOUQUZ75VxoODYNdAphag3Mhn/N7Q9WuEWv5crZQsf
JEJrVd8P7UcWOjenkPO9udD0eRyP944CCdyAjXuDqoQpBjNX1U47TM4K3X8rNOYV
MQffPmO90/TV3JB7BUxTNk2LmY80JucCxW2v6jGliBEvr8y0nxJyq2JEmQl8tT3A
JU6r/sAybTRu88/qXbxkppqqJ9ZfheHOegttfz8haMCpcd5F3zN4EZZlesdxjHua
AfSxwQBzZ/rfBcV6g3g42e58MZYQjrKBQwG3PRKRFwKYgE95TYwV6KaM3+jczdGa
o+oyHXDh3Xq8LyZ62c/zJgh9RZAvQTS1AWPnaF74Rm4aurYxer618qneeWR7Vo2x
0vlEmHw6jkO5zWqGGuO1J9Zi74quO4sJCWcEED4JGf/VlwJcewjxok2hQ6lbFF5e
CmgPeiSdW+DvPgjDh56dugN3ShSjMDSnG7lw/YwGS90+fFOxw7eaSth44HeGfVEh
RBgKanIMOrJml7ZQ7Lg7YTv/SZmohmkzpvu8+5bU3lmQYjfZ69tpx9Cuxx8AwkZc
8E88Vn8RSkV8wOY5CP+m0d/mpBwzIZ3KinFzimCC0To7Uxn2KwXKOj/6t//7Ez9r
1W13go60HkAKNmcrQn+pqcVnmRUCvnqhBbyY2WP9IacwuB4OAxCfJgq3rlmBmnh2
j093fBFSg2OzCcFo9pDe4b0x3KlAhUZ2ZgpgsycmQFACjdeFU8AXmF2X/8sELSQM
17i4FqdzptV49Yy5FHF8mnMkn+qUzDAziEumepyhOieH/xuI9+hH+pgS6XRk1Aw+
4RD0RG1W72XiTgfHa5hAsBZfW24DEUbREJlyIY0d7wWWN3co8lWEjsi43MCb8tZL
Y0QseJR2/gdgx/MHCX/KGuZeu9xEDrNFkV5+iRlzT/3FMYIykETVfjBsF7Eh0XmA
WqgUGdAntu4RLfcJbM4sTM96YpeyDTTjA9yOzbGviTPr2tM8ymy4wby4b7I7ncT2
EP1fMOwFNayvwfzXEQNUbLjgFKG4gCUuwuOfmQhIyQuC/JPJ/f5dEsK9ItHYcxO/
6ic554Olp56TowWt7EzsYSTNoTFq//r3yW/Cm/CPBmhx2K+lgy3sg+EGAV7na0Sc
0Tp5jcebMjOEH+FQfu0wOOsoWrQBhl1YY8e1hrQAc0CXj0MjpnBimDCiMPIiog3c
6tFQjvTdF/sv9MEImMREWVOxJgoWjxRmibuINq4XuN9sV632phVtgWXbbSaL+Zii
/ZHMRO+EpPXGg2A4KLD8c8Gs2orKXRuUR00QtJMxibLdClhNJ91b1kSnWXexOZIr
FqKEDiKdYB50oDSfOYQSVPbCC9SVb4gmUm8BD+weBv7RBJdtOSH3V4edNjU93XTY
OS35Jij1RRRwnNG/dmu+QSyNOVrmoFzuVKevLfmvUavkrUtxM4YZDW0xg+ZW9HUR
LOXLgfG6UJPIayKx6LFHkCMW708e9+8wDdGwnBIgpyKqd1eC7fEskPh7HSKqYR+d
nqyguODFLgcpkFHIuFKDfiZArGyV2KRxFjeV+ZZiO9s4ZjcdH783m0M9+/fLA1R9
9DZAnKuvss5Iamy94N1fB/1+cZvmiXjo82hUvzinUoGt8lCvMuuQAVcSX2iD4uXp
cm+bSfohUrNqIIIjDBOTZ+JQ/vES1P7F6cLLS9IxNtqB7mAaqVXTnUPUNuV8ZZvh
71V2B/ba97+GHcBBhNCJNo4+Rpz0FcBpZthBJhpH1NTouNhQ9F4Gwx1Ik3hRKg0o
spT1T1of8PPhncnANkWceoy/coo2pR0C17RT6QZO+KkX8uWZWjvZHXQOhjimwOmh
o2eD3YkS+NkNcHw0hJgNfFFNhiIA6ElWp5a13NfXydN2XACaIuKMRxqxIKAdWtym
AjEYquTodfkKL3xeCvw/cdxsHHo61mB9tNdSn9xP3L2lslua4PvJ6gKMadP0QLiT
73IgndAqvCd79V7szyBd9n77E5yxzXXh9YezUafGBG84XGTdP0sxJk9H0+23qSUi
VFuHGA7g6qsdGezBE9bVAMxdi1uaf7Rp4E6JGdNqmhvYpRQK7u5x91R1Ao/aXfWp
h9NhhUb0URtz5YDkJFTXSHzbkquXY9+b4e8EkXmrENVX25t6sR4XEHZewCdQMLS4
nvabSxMBNDbpEHhwMi9dPyNRsHveDrQ891LbkixeGwJQ3UWu92k7ks0p+PZ4tl/j
x+nyvYD3bHNi0OaSVBgcJ8UBMbCkIku7R75i8S+AU2IO/zFfZuP9h1PqdN9VwQUO
5eZzUqMMyRSF29AeGeI2p+SVI1wr9VXis8f4FgIED6jkWpz8+IxcWvvqgtoBAlnG
Jt4N5RywMfROz6EwVxNL1bfppSoBhwnwjxDVzdeem2zNda/slO9+LfKBXtsxwBBn
+K9+CrVgObTrhmFXb3zMrWJh1PO+/Qbizsf4aCjphHUbaO9rSjjo5t9K4LPvjBWN
v6T6IO2LH+c1/WRte2FrWsxkYWRjZZmoEi64LO36ld5Qh1IaQ2KTUTwzyQ+9zSfq
XBS8Oc8LlppQsPdoYRYMnhIOFX5MYIaCNNaYEnsTPK/vBgpib9Yd3d94OaUDkE3v
ju56QMCUNUipaVGhu+phqGR+GRBwdqm8kmwBGFi24Hf7dkvPmtGNccKb8O5nKnf4
pnjnpyDgnip5PMTpoAZN2VUPbx0l+USBOpem6iycOPQQFUJmjBWa+hPrhv+1+EZN
qJFf2+sVMiHDgaUtouotAJmhi2zNd7N4NWCdg+C/0VengzNPIqldjF2gJzBVisAD
z91eyoOidDX2OGVVzr13B1IUCdY0TVXajCMZ8c6ZObXFV5mt+qlpWc0jzt3CHPjb
CkSnSyTIDkD0CLaExD2E57nT5KvuLPjLsoSrmG8dTQ8=
`protect END_PROTECTED
