`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6q8upRSE133Yb/nG6rshj3XahPx2Jr2t58aytJ0I+sQg5nfzSAkPVbOZNC7Bi+no
kIdgN1wg2mu251EobLTdfUwQpkApKZWEF3o7zMNQw39Iv8mdv7/KiJzbgnOPhrPv
Mw6mYltn2MGGDJncVVqGpeybYEk/CDJhDVIDQbLAAsrTdQ1g4E02FcMAkzeUoL9M
0wx38PlXAm9ch73Onk8jkC7LbJMIrXPNR8prM0XhhxLURLQQMzdAaChS6xfUKYTX
9ra7pijCfan2DitIwxoyH4UfKc6d88BAL4PWX868hMg918jVuSVvd5SdLWLIOMXi
/Av56RodqI0urfy1cI9iBGJD2HuTxSyI1hMTrhu1+HImMDfKpFFYRASFvGdhvDlV
PLoYpA7zqohYR5soZNFgMyRTeNOGnukovcw9gdTQFHfjEp7Cv0zd2hvE8BiJP7GB
losyJU8iWFwsQC2S4LvZZcD439PpGiBW8sZ7XF4X6yJi4rnZchXp+y2Qwpr4SL/A
/PYe+4pOZBTSedJTdHTlADwItzSg9t5kUJKPwH8rMnhLeq+YN8KWs+7nAMeF2bNK
qWi19g+8D8DaWHWbWQB4hCB+e2G7tR9xQDo3Ns2HOCfWsuDdshuMfBMLozTBLwiG
YzNlDsJQnu1I4EfF9WEraPrSg80xVttwh0T3LEJFNvp4i7D5v6GcQwAlh/n3PLP2
Qw9NHGtHy1i5IfMHHaFbYrmurlvMHP5i3OYmvfr3kAJTvjMUI6k9ef/VCbOdWuph
ZDUBnbE82lB7tOMnJAh5wV73EIvAUQurpBgZkYBzWuCL7y5SnDZNcopwAYnQqAhr
tMk4RdkruMO2LKA3G9V4q3bgEmfQAlkDA1Mkv3h6QhpycBpVhnbmalC6uYDQV4rW
KyIhvIXf7E8dCll2rTYQ/qyvwH2aCiYE8njSHrH9P738QzdvAyzxD3EOWFvLtMbI
Ob2VgvDfNu2KAVkVJOYlEkEfoec1CMpwOIRpNUEUau1nm36nDWja6beGGO5bvQO1
9X2uLZn5bzwMsqzeLKBhdkB0NBNkwZsXj1SDHjz5CXG41AXP2whodJ64TpbBPKpu
JTLQmpmnSYBBGHwv5+248Rep4G/GvWF5WdxBt9OXkSz0pT7rkva4bRbn2PCe+bOl
qZrkcN1FsixRlySIAYLkSqy7GUhjYcIIkxhDQFdEkchk324RDiUmLV/kRhq4tu9q
O/bMVU1AWUjJDiT+gvJVtNgB5RGUulZUBG4ZyeI88yB+0ZS/GUKYVKZGZaSqjlmN
3rlv4vSw2ERnjPvHwCC28fTJm+oARube2HXI1YKYF/zLzK2XVa96CqoKjE004Amn
WO/aURJka5PDfchwjdd3Xga5f1u63noqpGkwUTuSVzY7gN5jKTArhOZlXUBhJyPN
XD0s8hOLtI6YcVU2EhZ06QtoFxyJa8HSTlEi2O0fGTolpoh37ZfgNIPzSqJ5jfLr
C+ky8ZQiyMLqjcBU2c2PhMvxcEZN3/eyxjxD4WrhAHKBNBJfFA1HpOEOuBikLZ18
ijKe7XWOqQ4uVsKhrj+/7aIpd4qiE3jRteeyF61/myvISnvKd9MnstjaT3pqu4pv
+lYvM/lNqXgpZVD+CcNMPZC5W/lialhHU0VyCoKWVBFx9Wp6wrsgd/nHEqEqljVk
Bg/uLy8j3eyAc9Mnfc6wlyen3GsNF9sflQXHXuezR/KP4AuFLeUwkVLHiXGSqjxI
X9F49n1uHPOTVBdfz3fcBTYECeoM90F++LJJkY5JhJQr7kDGEMzA+X6vmWaksoKI
7OrIJshFmUnqJoRfZxYxnMpW17YZdA6Z6JQfUlVw+y6nbhqtw6jrhXxUsv1jJgmS
q4Rv4cHDtjsIEiRGhp2x5RmX3s+wXiYITWbE9WOvtdaFEndXJJgzv8jfJBDxmLCU
7J9uq01gurGHx0z2vCWC6nlgzv/U3sh102TLLYWAJD0=
`protect END_PROTECTED
