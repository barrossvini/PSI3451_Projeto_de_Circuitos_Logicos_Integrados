`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hw5hmi4iTDsc+Mc6O/0asEtn+Mwm2pXxQOYnGGZJwsRLX5iZ1jWeNjdSS6tnjzbK
VBgeghf40gjg6EJ1C3b8s189GL2/xDt3g8saGghg/C87wKkCHJNaSfeyM9omj44s
ZgI1uf5/ufxavgoi8kVC1hoGXryjqqsPJarfp8KLIKveUdt/ZVLuahbYv+ptnXFr
f+DXzOfMZDQw7wL+Zy/FGTEWw0MIUpGA4qzHQbzgAzGWiXXDT7cY8n1pQ1H4ccnz
oG7/cbZ0tm95CZDojRLcC+AUoUnhZjI2w77gbbv60jTuoObkeVBtwgVpBzSGyPe9
Mb70DRJrwhCqKuxo7jy++vwX7YUhUUNQ/MNpawtyULDfeM7BzFLboLH5N8nPVjrK
0HBQgOIO10xqCKWXQJufk1uPID+wEdpQdGjn5gZawf6u5bmvgtxwpyPlHI1sulVe
/xhcVY1hHoPjioZqzL5QEv2Nbt3avJP24U9cStu8eMmUvga9AlelwjUYH9+A6k/4
Q+zjxKUXUGmYDTj3Bkf0uKYcuzPBajb0wc9NhxglLPaGuZkeP9kQcna1E/kUVqoA
CSQJRxAeEwWRQS57xJS6mV5lDbeMEDaMlSEd1tbvSPRW/IYxh6RNguWBBZizVVb9
9F4HekQqg8HwDCwFYamMweQaF6EKAYtrBkX6t0hxIjtgK2X34EovXXChPu5hGWMN
PJwaCUKEYU5YeCl/UQknA7FUgyUZwisOYi4Pe9Ubb3r86ZZw0fAFnbk51wXwEqJo
q2omNOhQ09+U0TIWKjM+TO4L8yUVUaQLq1gLPAbllqpBvosu0EytFFeaaNMSC8TV
Gj60lWlsjUCasQv5TxOE36AFSZ456CI+/GPcm1IXQPQjjX8qeH47oN/iob+CTqe4
vVRo2XhqH7eYiQKDekvTbIIncLsDCTqCWAcGHcBBYydI7D5UBK1h4ZkaA4TNjG0v
ZGziExCHY7LDO9+0G+4HiTr32sVLdefz6RcIyV6WMP/nejwOdX3G0g71x39Rb6oJ
RPk8NKI5VoVw4EsNLM4gpTFVu1lOqMhxt3ZDCpOtMNcC8CG2GzFLepg7A+mZ2p3s
1Zeq73OTDYqYLKSxMrNZX/6llrqI7X45xZ7IqY5yNYYoY9HPniMf/Khyxywu4i69
Ap7GdXg43EQOMfZ/3UGOScmzOVKDG+3j8sN59PA5kG2IOiQdeqc2hWQ5dbeJmx/4
P+ZeCU2OflHC7SP36oPghkV4O/WcJEUKYHeOjF71hRy4/kKSSgJc5GVm0bQvN3aY
BHK8DlBEPcmb1eUfSLPiGyQruIUhA3PMuI6hkWltu9Ot5AIsePxJRSHbB8s7hyZY
p4LLJIcXVDsuaPd0lgjquK1RDbA/EJgUCs+I0uZeJ38O7P4F4W/vl9haJYsJBIj+
dUegTniwzCuUw1USI7p6zXsp0y1qTxjbHr3e/Y9bnROrUZz0oJrItpaM3T+tHTAU
zzUYe1lFGYlsBWc9NVwM++2McEkVoze7O7CsYWPJYjS7e1TamHBCm5lFE5SSCKrl
hyJTCDLbsh3n8iWLTTXp+kZBhLsnlBFFYk0hLTQqzJlqfrXAB6QBCY/y20nftBqI
QKTEdz5mMPAxH6hHWq2KjOiwkd58da/m8KZ1cJ00rb16CY9++t+O2TjdlHxw6qWj
`protect END_PROTECTED
