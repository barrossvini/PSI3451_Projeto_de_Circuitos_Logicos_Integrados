`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TzycDxyrKvovsW8CWev8NIL9v8ZQTj/jr9uznjEA2J8FKk2cBBzcjgXawOULM1eK
6tA6o/lxNaW8NsW/bhw/tFj7tuDi1QxSl/CbNS7OzGB9Fwu793Fs664ugPWOyRpR
4J3Su8bgPFy9OID/6LMKRZUp/X0s0WtNCnZWSr3W+tkO76njCbgY/MzbO81pl5Eq
p4zDHbcJ60TAInNaAWc9MOS6pg4xhEczTHGZQZQdEPtRPlxMz78Wh+fldT4KpoCn
nKqIykSNMzk5EFJMRIimY9XrFlNCoINR5gt+JS4BMOPMfNC/u51Nj0KE7ixZ8Q1I
o1fXVtLjaho9jXWyTuhBCPaUKfH0c5sMy96jmTv8RvF9FxbkAxVKiLiUyILtrRrz
p518iiJbQm4apIQRhbz7q2d4mF2BpxafvgkI4P0difgxVRml0FQBg+A7ZCkiMZ2h
`protect END_PROTECTED
