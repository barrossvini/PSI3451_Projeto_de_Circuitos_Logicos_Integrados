`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L203ht8ncaELxnMZbAnpj8KaPvhjlvDx1jux86DHjGzjxn3ps+6kS2KHrKBQmtMy
MmOa3KMfQM0H6ZTOgDcIj2bP0Y2KTKGrPkbtxiYTqYd9eO52GU2s15etZHHeckvs
rFNpE7/79QQdgElr6/QCNjWFN6x9pEn2EqrZcDFyqwT3q9V8HselvZcXhuDseEq3
4bcICra/zVYo/hyQYEBBDOZlpUfRC5ZKySRUZxKxSXC7K+bW49rPg3LNTEkXoQbg
nxd8aMZNiUVp0eRHiZqWA/t+cSrwZat1LXn0MGalEhcyMa5PaI2NyFu3d77zW0bd
I0fBNjxePG6y8baoAtVNaNOfXnbfECP6vzWNONGiK6HRZme9aXthG9l9Y6AN777D
ZOHmyAIRAiC2eIUac8IRJXeAMXClZWTnG8uK4wZNlaZa5ySPZr2iDU0jhYhUzQaz
bzifRXYr5wxCR1O9rSEjaMMMhHWF52EwOXguVN2vLWj6kFrUnzgG0dQjIhyUF/r/
6Gx6CJFGY5FyxutByCkj9cFT1hhAt/kq9D3Aahh/tnT2/7lOaYXEsL8yyiCAe2/A
gKPtWxiVEppjIIgwCBkMjYJRYqJrpK4oN4aas0eCJBAbpdFKIMWfEBVUN16gfCFV
35d79JYBXOw3pVKpjarNqckKAvoWBSvm+M/vU+komazG8iPPemQWQEtek96hgzHy
HnbpyqOSyZ21qw4VOGQjQQqv0LJ/P5jEU2exE1qdaAWEiZ3ioUeFjSkZLKpsM+CG
vV9PlHhhcnn1MSQ2Qb3IszYSO5YfdLXODCrdMevLh9ZcVLzIf7dsLf5d8a5ZKMLX
aZlWc/J/2DafxOQscqzeTJYHXSmGv2jmCUGQwBwbwg6BfGKI/mqCtyY7VGruI1YI
aoQv6oDaG83/SUjQPBJZk/gYN3ge2Tujh/RQpm8I89emwv32yFOIBS0OjZA5ADwJ
nmYlsL9e0H/fn2TCnbR23saM/HeqqDSU35UCqqbffTdQlgLWrxJjiJ/hR88rvi9V
reijbS1dtxjgW3iQN29pR4aSKDz/XhdjyioVIy/5ZmrPldKAsuQgYf8fXgQcHRv9
vzkyImBDzf1r84Bdme9E34JSNw6Am53CTnUjVwc2NaLjgWy43Pvk1Kum+NTJHWPw
Vv4Pey7yIeJqly+sRDr5QdngTAsTcSkx5UiJtifpm8IZfuprkJngY2/L+XZLO6Tj
Ebh3fsWRoweteNKIUR5iR1s9F+8+Hd/jaiGhwFOnKo/w0FHiYNLXNCKv6rxtqa54
p3p7EouWH5GgwFqnSNOatwXyjS5CnLfOzA/zoWzzQFS09vt0XCqx/n6Xc3IlrTzq
KAbLp48apevLvT2LTBrLWn6ATRBlYxOadTxa85upGru3xUtiUEwidI2NGCCeO0wj
G8ZSoB6JIUMldQ/RYnx0zw==
`protect END_PROTECTED
