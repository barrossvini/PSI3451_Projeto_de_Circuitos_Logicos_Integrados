`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZA3xp/gtPFQytgoeuI6n3ddRp80gWb4H7auabrJBOxGls6Q8LIRG3ZLAh72iDRgd
dYSWJTloNpCXVgIAX43Z1Po6DBmscDM36AyYtq3pUPQm6gGPVCLq43peAbOeZ2uW
Y30SHBHmOnxIFx7t/5SYkpHUYYxxbxTBHrUUC5oO0/D1GDKjcAkPhsyrg4wImt1x
gwlgPesRcThmFgaSqoKxUl7nJiIgq3EpFO7SfI7Z24GB/kxQR2LDOmdS0S/IAipO
uX0zmkY6TMsDofXm8h65oQ==
`protect END_PROTECTED
