`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QDkN8ciJjXpypVs1Gz+VzpZfpgn5jx8TdyHD3z/l9H4WHAZ2FF0l2r05aOExPt7C
QdOZfscYb3Nx/tkd+clblGZkI8aPB0/Q4jSzk83dWLK/FNxOfnaj97m5cEmS7VvK
8ke6+vlQf8mzxri2fo/oFcOVp02+REJTfiopCWZcNlEpye9g0j8aFU3DxnefzBoA
qM9akbfAKJfYoeqMxPbOu8ANxHHcBAqRT/qh6qOchizUhmBxOPZ+Wix2i6sTWXF1
J/JKt7cSLWavILEMqZ712IwICYkeXuJTrWg5tnhsghznGXjItGtUeTBTJm/S5NH1
9ahHCPpPiV77xsf+U0kdldVupO+cLh2rW5O0bfwNFbE/fVEbGbheMcGV0wvCmDhD
h2eYaNg3kJWWGOkUvs1iHw3GINaqP+AyTNbNReTZ1/bauyePbu234F3ARpEocGku
iAXs6vqZMmO8WEAV3aBMa6BP+Vy8oShlR8UenFUx1BLLN00D69y8O94cxK/kAIdk
cpqKGMN/lDbbl9pa2FKEuNWzYnMzFrcEbEWY8PBqwQv49W0vmJ7rSMv1ZyQ3sYaX
HQUhCfVYMOis1JETUrn31OZxByC34lXAck0wPP1e0GsmaoCNyqrhI4Sqmgz/E2+w
BPVK1sqDAMV8bsoYhKdJkNMQBMBuLPjvI+jNwfGDmARJx2Q2gcNGxBKU75hTTabH
2j3uwkUk0VfEdUVg78jDDXyLXNx1LHhC7qSEaysHUCdb2/0WUit8wkPKDGeXAixb
4dsjAh+930PYSmtB6ra088YQOu9xsePt+OLSNS8V6/qlSN2MUD2bAh8f3aysBBJs
lTOFRxCecyDUUOps3gmQ8QirSAmZD6ayS1QUxo00OHuqhW/xho1fD/X7Upe63ofx
ULyW9W1qQsCMcTK3Bf7QE6DPfQxm6K9L0U5aNaOwLQ1tsBp6sFE8SXASkMZCOlcd
tEHNAfsJsDd17O3yBEoJ2P+x8w75JzSUmj67lSbN/u1soNsKeRjRw1Vnh3d4UlKz
R3bk5JLvUm9X+p3IwkUqTHOeI85k+3bODWt6AMBN5P6S/XE1zcDDNWXM7YkyD1ko
OwPxGHSL/z0UU1tysz7wDMEYEtyRnPeMKXXHPZuPcdc48iQ+IrW2uZhhvay4VrVp
AxX+PElsnS41PIG6Q56L5uC9fvnbmPyUfpwQElS3trPdtAkrmQjfxKLGoT+LL1dp
MKsG7Awu2PYO/HUQQiFp6i7qsiLXQ87WfsRcxctkx6oeiflijc/mZcFbigSx2baL
MSd71KaQESnVXKfJRV3YT90S2MQAT3M9jivKppN3D4XSwoQkSp0B4s7P0lFSE51y
KMS+uw88qjV6bJn5hj4/ZCIMjDNdQtACFk92VhXbA8w2Ap6PtHR2C0/SBV9DzXz5
mZKI2BkIyI+GcTtResyn2CYI90uYy0zTIRJX+z+LR7jtstZHaocuovCkkWTuKIPu
uaGsFXkzEl2zEr0cP0V+fpCwV0LsZLAvcsTKIl+RvZyATPGZ9S4LFJI9H8V1sXf0
qsV8ZtaZcct8QUlbIymCJQ==
`protect END_PROTECTED
