`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ELSTshfwdjv+LYzsDxudGPYt9/QD76n8yzo3begVY74PCQob7pnRokYZnpOvUwAx
wFRs/g5redhhXkcNerWVbaIuHBqEoDuPVolgrPVRZOziGjldKdGbZd9yQm3MOdyK
a6pIb48oP5y3Qjz6cI2s0j73Kaq5aG6Prm5Z86P/A4P9fnu0usgVLRoi/12QsQm8
Kux8gzDdt0CXFN5wsgQiMuMp0ewagEiCpWXEBau+DUMsrlBYn3rbNotooxeNBRbo
yBhSYlRwbNVw7QyPM959k0O1xvLcFqB3OVKiaWjTK9zbNA97LbG+KPX8ywgOtp0G
zomi4YUoYOPxGHaL2BcbfRXnNaSis5kmMNPeRQONREVffBBQYTHTgQBhTadlhPL1
r/iK1PxOb9dSDt3v5F+NU9U9kadolpWcyA7WsI5hzFs9aBFFc1/OR679WDFsERHT
Aasd1unNcIwEed2B+6MnmZNzc0rW96GztcPK227gxV05Ig+h3OnMbn97miHGFiH2
I+jsPpy8NkOmn7Mn76Q21fdoArYTBDcz9AYnYuBBibctiW8kixP+c2wjFue83Ozu
ovvsi2ZCiYr9lrlASNLm+leYnhSv2NlFOPK9WSka0YOUhRoZBuWa8MgUw4/VGu7a
O6zrzX4I6UZXwQ2MIpV0qqXe4s+gT/VPzwXi30pLhXKdVCInE8VIyplcJCoXUnbF
xBDqO2HFYDQNwgXKzdjYG54SeR7GcIn5KtyFSaLK8JW8SgjwYeqOnQBEzDj3bKBS
gvX7YwwypsD7e6Y5PUCrwkJ5em8Rn2ha69SiXRVK3Ny0QyPqUYA/yugvJjEV801R
9aoNluOG91Yf5Y0wqsX0cwQLyDKWmq6hwtrt1Nqsdq0maFHpUw0Go4Bl+fryj2oq
tzu1dubo4qzaiLeWaRA/Qi/ZYD+0C3kk4QGmbYyhCbXLQ5X6CpN3H7hz3DYdJzX0
tw4Wt4WbMjKfcoczaQFuYsjOtaCXvfnB3XGzHAD7caWBGdOKnzP6RGzL8hz+Cpmt
iY57UIIrE8gAx2tD97MLAFHL7IFBtZJp6MePPqSUTEPoz75i4MQAE/+6o5Zejw5M
6u6fm/5vbr7AKQ8+FH+LVCCojFxOUGwzMPr9SFh2NA91nxgg3HTPhB3QFovo9fkT
qb6b6V3PLYI16UreMbWW1TAQdyUip7BS2TyVJ1VAcAXEa52ptjVbVDuWWK2oI/qW
Clw5bgD/Uq09SUVFjohKHLCB9Yrf2Iwi7yJ2kD+Y81JbxjFlsejAVkNcS/naGeEF
PQy4fJ83+loJ2lEVBC3HBFB3i6FeytllwouQS8TZ6/sv4gTBjvPZLlN7nuBqxl/R
M+0yGIpNl+2LrDLRj6x9rrG7YMxIrz769KIO70sxi3JqnVWGBvtu/VJw1V2egxBh
tg+fQIM+TndsJ4Ej8aoP8lYSNX2fbSQkt20im/1kGBm6FIB6lzLsLIwLKJjPmyXQ
O5lnQAbFz7S9qEjXg8l3Ch0ntGwyoK1E7VOlxTIfVo5pxEQb7e+k0mYgxbC/PrtB
eygWhqwNx05jbxBJ84kOwwIctrp1orcTocp5u4RRDejKY5Jnwj4oWBm5SDiOiqWt
EeOfu57tAUZBKd0LtZ4kU/fpJLN03iYoHWcRaanTvXudxY64ZcvqpinNp+9aX5sd
apUZRj56aYeXC13dio3M52nvGrWNIsD7/3aum+uHfx4S03mn5L4aYPBNpwHhW40H
ax5i1yrwnzN3/Jq3VGCNZ55fzS3+Q/KViUsz4Fudqr8FFAleCfM+sOYdvtY43rtO
K3hj1vVqVWvgMdydrw3Ib7PYIoQYIQkURPFLJ+aDKc8m/laqS5w+whUXzzEASC1Y
TMaKr2YfY7/Z0OuVL2Us2pJgxl9QGvNWTsJ0J7XsIzB2fixfZ0Sh4H949q8/aCmH
sc3P+oxmzxzZVHhrnpYuIT4Ozhh+62bjKE1uQadvQDq5jh0IyIt2AH+bTA56LVI8
C7c5ttzqrx5F9EYWobVzQBbTf5/fgi6I04rVBNyVj2JKol95KtIxNtiSvfVJc+kW
4nKVvaRXQsYEXzsOfou7NtZ6sBl60y8YSX2bQ52NBUSdh63e+iFklH8XUhwvm3lB
Pj3oWyQhuy5jpVauD7QPuiI+xOHkHpS4CjCqW8oxNrLKRHr96Cm4Qo91fjgUGkdJ
OUMNSW8UUXy9ul3tu3k3yF4TRM47jd3Zarq2VMrVH3EUx8hE0a52b+5HJqEQwBBX
noMvuB2leXHj5btYbktV1o2ssmrdeZXl1nHexwmoH0TW+dfGe0eNUVlwVdkDfkjr
4C3yoKRKIV74DBTqaL7ErSm1G9vph5Py5oKpW+mWC4c1XCe4ybsiFzFIsZLtCF7p
ZSgztoG8SkMbdVk2h0BqCFZm8w/Op2QeDNHQ+CxLgtsIAxnwlcJdPJTsElglzgrp
obntL8lG82lRk3degZFgwlxyNjoH7QGOrCu0NBoNU9JO2lgzB4tuoqeqkQEDKYmT
1/13mTxtmRlHPptPIIwDTtYs4n6Ez1KciVdr5zLmiB+OyNKD6ZcLuyDU8WBxEUY6
e1+euRG5B9u+52mOaJBAydjt66fK2jedaDSTLNDba4l9fqof+/P8GDNNk75Bmi89
vxSFOMNH5onf31KxeF2BE8hvqEZDsNhcKMAPQYRvxE2S9+8NFIZV6dU1hv4QS+ap
xyJ/JwlbMKOy/56VXxDTScA3LODoAZMHfcPipaL45fpSvp0Qog1TFmcF+eof0p0u
fvXz9gatxfmHNtjL0/U3RygkfqlFxOOoexuIWMWRMKhF+ThklwTzPsLyT1DS5w8z
FZ5J/Vul+kLUpG9cgh87ybfdYKPw/S9o5YLgQLVj292zXuD4eUeAQ44CqAvAwix1
eT3qymm2RA4cofYmYhIbxY5s7ZEnhnuGPSaw6f6v1IEpEKAdfxm0c8nD2wk4r1LP
VfXGQ+q5nYmHPkAwEljMjRwspJKwUucSAAfj52O5C3REEfD5M23AJvxscHLYKKax
NhuWK/9LHaVoqNAkeBtM9ItoahMF2dLvlHgtF8/qZ+z0T+/Soxarow3T0WZfRtHK
aXjhVYHpXkoq6CWFyGcMgzTWdHUhEouxeSOtVMaE4jA0xO0MTAhVeD1AdYSKditg
s97NssQQZNel8M/KBKvsVcFU0pCyH4ULUaum5j3AtlXbhY6Y2KScDzVst73JviSL
Q/Fk4SSoqZyEPeiHcbhEesMMjC2u4j2YpRgRe/e3Els3txsc60Rz66YEqBbgA0mO
OV8jPlvfsdV2al3ptJVLwXqUc7R7JQsYWDv7mOhmJiNlnCbckVeb0JGsWHAibvZH
+PENoT45IFSZnwzonsLnGJb+jgLSsm+HXIVX+l9I0slIU9JRpmqpjb8c1dUq040I
lBFb5iNWyPlbxZhQLo5gNxu80uAf7OvirGqIkx3eL5rAModlMQhwGYVT7NCU4IJf
kD/wSNB7s2a/NoiBtV6VYiTvWXfqV58G+pJYUOUSGFP/R6VjNqZCLuw+quMwbuag
iajWXLvIXVIO6XX1jCk7imeNJ0UP6YnO323BYvugUTNzIvdwwlYaiLbEdHbm4azR
Kx2Zby7/7aMMUWhdPg4LcpRN45qkvl0wAkpJs6jAu5jObclEHbG8giLBcqNcWDjx
aZeTRwU2PeXbOVRHbB48IDD00rF2GkAKfT0jQ0WGNEvOIcTsL6iHmb1GBHt4BAe9
raPgPfqgQnX+5am1Q6VfjNt0rZpwODEsm1W4zbgYjMIVDA/zIve7xPDNbS3fIHWZ
8i7KCj7vG2xml8iMQCw+OSQ+uUV/ZCbJ/bKnnR3eBy5p3ZZtG73CEEKVSvd0sGHE
NftHVc4x8Khil4NfRR4A8UJkhTc0EHP7bwc3wbnl/6UsJBCKsvXyTJKxmFgW9UUh
y2aQMJXkFTzujKokJmW/CiRZzyOWGvt755dLuLRP0moEyIG7yoPfbD3OstYBI5Fk
tNdTKST926bBmo1yuhz011IreWzmom6+vdcWiTvY58T/Nr41Fc12Kw4KviM19hfP
t1rSWrLtpnAZTucciiUuxOavuKnWFGWBWOh63sSHIfVhgkjevvZv+5PUmFPaWKh9
FUfE7ek0D+bJpck3mlbEDkYqUP4/iPmAwni/nwfSo0wwaKQAILcel8SD1Ng91GAs
AOQaeve+xBDHfdoQP7TOC/Q6EEKhtdfUozJSG37aofZz1a3zCMj4Kozzbx158DD5
OTRUdCHB/lrOVyMpVgkHwUAvNVprbgr1dkLWWqcGsjvRquQz2t0hX9suxBX9Ax6W
v2IsNaj8J47CtHGtNFcFAHOE8kKMh04CwOjANpjPAqZm5lxnitJSefiNvOvmoY9C
kcvBoIHAQMmqGH7rWI/ytI/fnsHnDJHDYWiYIBhDVY9z7BYiiys+Mfb0yuOSgYfc
kPsfyQ6Hjh8NZLSuu71wMsqvnin31Di2nRdzE8Uy1YDgTF9c0EzHCyFXCXcc2Hcz
y2i1cVMdkIW2vhxwV+qYiVjfknRu5x/7SvbB5Lm04CzRzeIDu5LiesGIEZDDnY+f
pMZPqu8erulDvVeGI1AIK9NinfrzmBtPzpxCUuGgPNlot9xnEBMuoNCP/8pEIoga
Odxtd70XXfPV6DzBq4Du/0TG5bCvAAPS8fNuBsAs9E5ne9VVUlaFrIb53cmRmbQH
bMuZbxpcK2s4RMzY4Nm67hxRPO0RFsBVCqbeejiof1XnRt3b859GmqqyoSrkpOGf
vIQhjFRRd7sQsUZeTxrXeWRLM2L+aUeuh8lHgUMnzBDFfgVqKKvi6hiuFqwDpR0I
FTaa4EH/srGDAqNPR3LgAWjzGukuc090ihJqUqBzLWPXOj47g5e8OXYiWP8zTdOO
78wOcT/hJ+gpdzuhKFV+CDsKlWkv2wur1YXX2w3BoxJ1oXXz8uT9k/sjztF0+M04
XQrljYHMMvl2jp/cj1CXq3+4+xRTKOP5Ect5uNKb+6cWkFkJggVKR3gBKrOCB0Wl
/7ABUlviQSJuwC4Ac/Ym6nZefLXPFkKydeNbC6giTsQQujaR3gr0sBRRImN67fRV
9g26FbVKOfxXbijugZJkSxa5vrFdVuGrJ+K2zmqAAkaHCt0fo7n3yUdtl//wxD2f
k3vo5vQDYfXIoQJF29mY3oe1U83gzwFdn/S66+jfpPs5PBZ4kKDckY9Ipsgq/uYp
5T1WpHNOdfTak08aaZvJd+kfYhYFDP8vMb38nXnCDZ19sU8ICvvPx4R7Ueapi/z6
W3AzrNRsPh07zWCsHD2m4ZX8XqEpkIwCrQCctNg70b+S548Vv97ODSUB7ZQcuUmR
Sddob/DNcdz4I3SrCgvg31QVxS20Rc8h9A2lrmjO/4Jjhk495U1frCy3IAV5m/9P
mMjitBwIfV5lEJhORNBawdKKEQLIxo8xaHbGHgUotVgsZTQcLmV5GmIx3W5uPIe5
P6wyy6kGfQ1bTkfpv6YAvuriKKxsNjyUavFRYPkHaf9QJb/XJILo2rNhkeLeD/1w
4z8bFb/vKXrf+eYHC/0O49ZlzIca6Umw+Wmo/8Y6ecNqEHTLzSKdYKBVSuz3vtQB
Kzj+gdz8Bm/gWy3+Yk8QPyO/bxJmrZRUrHL19Wft8txqdJDZilmgeLagDSY/kLns
BepcCLn8txhaK7jLKDaWmb3tdTJWJWS+z/OGZuLHAQ0j0nc7sQSC15Z7heZw2yc/
w50cOSickOpJL1Lr+xjfjzHYAisT+b5FNMyJ5fqNMqm3MbqeN0FYzTBqKZ1c05Am
/oEwQBcoT1B3WlBXfzjiyfNvDQAXFhKAXOg50oUIoEY1XylqU2aX+bf0nX2sFBH3
CUNuQYlrRVHOuAMrDqSrvHCpXzpAFiKn68msHPm06QQHQtEdfikx1i+eywwKeyPN
kDnWrCITaQ5oLMp/r9eB5m05KevzrAlNQK1ZbnmpTwLfDIa7N543RUX5oXGJIG2R
WHOQF0awrkVP949ot9JogEdsStBER01VeJYZVdtVerGq5cLjPo4pdpcd8ehkBszU
Cgx/9O4RIdRqnb0EwD2qcTfYt+Z7gUA3ZYeZ3W2Awy6v5sGvzOyuO2hRpyxVR76Z
s/8nPWkfuwk156RzrpI44cQ3urJWQ1itdlh6MgMPvscIG0sGlZVD9MxRBVMN80hk
fanccn80Sc/HnIvIC3ZxqTXHpNKoMivUk7vYwdjMFlnJ5CJPBQai0K81ZANpqa+a
M9GGZ592GVdqiKSszSo5UK3vilDfLJgmlNIW0xVSlQ5UciJrIBjiLmYc3oUqLwLb
NUXZfxOsnaaCkOpFFd2p7uHOxt6D85Hft8/HppPNU/Ou1HH//yOrixuITDofmaER
5/c+A7b8TeG7+HHvg9N3lnWQINeBQdw7aGqiSEJo7nuj3Tt2ypByi1JetSGPXIm4
B+87VVUhE/kb5jUvwSCUIN/I7ZwSdQxwZO1Q76KGDVQ06qZvjN3BGt+LaVq+KgPC
9PhomFsbmFG0yVOtjA4PU5baa0uKzCtraegUix+BeuTEGRbhXgZylN3iJNmvad/J
A8eYmVLy9f1SQYuGjdZKcbLl0NPqWWP2MEdIpg1oVRI6YPr00EUqQPlh+pEtbP4v
mLhXDiatWha0rxcnkuU5LF71mcf8Na499zYDv1n6Jw8feMCddrJ6ne4gdbnsDi1G
iUAKk6KV3l3EcyR+fGWB/7o+mI2gonvfFlF18Q5j/Dbks3eZaVIfMKa/kRmqYYi/
f7Aij5w5zoGDPmb+IaBI10J781dqPsQ8KpZm5GbiIaLtzIuNzrb9xHFBwibtldeD
9lNAERrzi9yB2U3QRM3VbRV2Ehae/4uLIiUbq5yxf87KmdxHzHDaPa+SjpVggqQD
JkADTo4HzjCj3hNRU2nUckEgMc4gQej5wxbcpkKPP6ruq4XnIUJL3mOZ/x/mMWL4
w5s4cYwhvn03tuQdrdZgVN5zmy/EBrpJ4qDcikNH4m9HZiocvkAwWoqxmlizb3S6
hNsplftQv+uUqVz7zM8sShnK/SoCDXEGYjEsphiBJOu0yYXv/G6OwOQO+EHf0W9O
SGNbZ07zRMYVltwceJ1Jz9BUDF4CQQwh2ms7xMldW7B0FsLEGEp8EJBAwFlxApYz
ouaDGTz53FriUZdjJYnxnobJQ8PWgMokFB4CH5uYlpaPIvTW1od9YE/Bttwlep4b
74jPjBjxa4oRPDJziy6+xsyXHgo9GjCe831txL8bMkzIqpMLu/u+zXjeuo4cBpxl
kaqPFRZ6CVDZEMyZq+eO+PhTDKCMr7m3zfDVxrwXtvXXXVKyGTa3VqHBXDF4EoD0
iC05bS0hlHt8zkhIChOEl3R44jO3wCqNFsNh6iUEdvSq+Ft/e6WRFr704gw7AZbh
UyQD+N/6vaO0P4RUvq0y+PDGqYbhDBFZk17afgjp4nbgTPnfgmJ70Z6epT9lbS7y
PnJ57xKCe0zoVBU7wAQNLCJqsqPfh9gC4Rz+BogHXfiPZlj/W5YI17O51ONetze7
yyhEuGEZFTFjgQ73nCxcBnlDvu18Hcupe5Xu/Aq+7BiMnTwgSyahNG+6NIt0CrY4
/asBWtlSTopDQTCI1ptALZFftxRD6TpCn33QRfW1uffomy4SruaMBCSBsvtUP2Fy
IgTD5fBYlBUVW+OaV8YD7++9nn6sq0fvje0b+fC6O7ZFbTmGowYprWiL+VKvg93l
iKb3zrFvwzHF6u563Hsp6qMtJn7nSKMhNFuFkKiNNndQNE/d4kiLMnJDx2zdO0rt
CmfB2g0u1sxLYuzorraNobvrBA92qtRCNP3vffRKqL8VEyxBil2AmT5vPzQc2c7a
jdgmrelSOqKtSvg2avV0xjMxsvPQXY6cb/aV5m7NZb4Y2DGjUZ5Gv9JpIhYSg33s
JIddFdfzj5u6raHjcucXhAxYPPVCU8d4nhQpYaNtkBiGzV/Xoq+C3MjmIeWhb54/
jAHB/htJWTGnHBDgYGZ6WeZtm1nQpr3ci8dYdiimXszwpzz5rkb1AJO/Al8D80oZ
rKZsQ2pn3fKUh2vCwPhhEdxGBJDTkoJtv6AWKlgIzz+sz6xP14z4pL+VwxE1p+oI
ESVyUHgpiR5Eg3j2R4yGEl+ZkXsnl32/3rEqXiSPB5b8X6lcZdAiK9YxDoMWsyYK
GsWy1hSscy1ngrKf4hJvDdzsvT4jqDKNKiPBj36K56VpuqyP09LAJpMTRqssJ49V
0mL4GckGUJgGBK7yVvXnqLJE61EqrYwQjf93hZoeagxrAvxUvXw/L6m9MB/OOx8K
091iQ0KoB+BoryRkVDWs2fYmJ+JxuJ/4//N6RE2XJGqJP42YZUHvJFKifiXRDPAY
+C/VhYIFu526+l0WFzyp2eZlOYVIY6LNTeSA9QO2UByoD5Cv1xC2ceS7EZzaKFXh
8s2+W/899Ym1OiHEJZEgY25Bi8NeW1tlRId/NoVdg2BS/6GkrkBOBtUs9DCqYp/7
oPhXNEfaxujWo/lA7lKOaQOb7zRrsTbI3tGIRQr3qyxnaGNjnn/XheUaXxRTwZTs
6rgl8Q5/G17rbBdYWuMwd2pB+d1bpsh0BXXWAJsNbKVcqu5Rxb3tzW0z5prln1Lj
k+5vUCNNYwQjzcoPyw16snMQgMw+19xwLKHcJrCnnobHIpH75xzhujacThK9ixmC
WbvIQF2R/1oKwzBUzG0KqoXAuU4qoRKRAk2shB+jImxyc7sgLuNkHjkqgAomXb5X
VBxJV/3LUKPE14yy8FNw7u8geSOuD1SKaVRU6aXayp01q+qDoxLQmTHjLZY5yvWV
rToPtrsaOtII16Rx4jOsErUaEoycnj/pgGx9VYZEch00NOp5+q1uks9YfBooaO4D
D15cmLmmkqG7joPgQUswievAFcsC8XZvZ5nn/tnxXC84hL+StOhzOF6yIN/b4RW8
/6CyWFmY4bgDDBFOXotPjshEXM3cw16Q4bP2o/ypvFau03fgeVmgfREfWtvgnhIa
7d5ems39OVbdBY3znRL6RbuVubw5dmTaM2j385w3akFql7f4gVDd6Qa6Axus6bvo
DpLDIbxNgdDaERLoCoRvxWvIbjCExQc78U0+z4Rs3bp7eP6Ak944f/dIkdPAB1pk
bQyJoFxQVQHV53a4aQ6SVue0sM6Z7TAHC8Z9hOWjVwcjtYYXW1vv+xzgqeucCEPs
EWv2R1ZmZPGKcwH3187D2E6R+WRk2I9O4i/nZY8W5l0/3rZ99baMCUuRMP54dk+t
HK11l1P2ySH4QpgXxctBg4MdU6VYDZ/nqVzH5jBsAMt/tLmZntrjkkVJwvr9qj6n
EVKuddlOew+Y6Ie2xJVQJEVY2RmLuZF37SDrfXjnSFqqs/wjIoTOeXF/EHCdTboW
H/eyiHrMN+uPMhqL655AH7hjCo0BmdOFz5oxLmQU5E8i9PU6KRWOe8a8Ti0JDQZT
qYppcYk96aEud/MhD7Da/cM6L8BV2Tkg3Ldf+2JUmVIfq5i6SnixTH0vXRUF3Qp8
+NlPRbggWqY7MCjldMdR9Vhv7HGaMMfXo2R9AMLfyfpDXRGm/RHKy4nnhw9zozqz
Q3gsP9iEpLGLXF2yOl3y3kXCZYtpgqbPj3tIADMeO9Jfn2tf6iiHaWrqPY+mHdhK
BbjtHyT2MmNzRoBEk0a+eddDPNQvaC9apBA122OUO6hlqdZk7LnxEqlZPHGNU31P
I1y0ng94UgYb5J9z+7YtLl9BbN+uVau/8JHtfvbGtOFnyoQQABnJrLvlivt7j23q
UUL/cG2nFAuS4l5TtJ/NkXbOTAoUcmtF2AvtklaFEyYC+dAmpritTOVNW9Rpy675
laFMTdmKQ4jBP5E9mTHWFoGrRcyHs+SWdju94/4H4pFJ4uVbL/mlJEDzRiiOX1Eg
LsClnl52NmOHXs0LgJETJQkPVyw9uFNiQkW1DAwCIU/RXODO06deLbl1Bq6FCH76
QT0AMhNZ+nsEKU8QIwfXNvuZFjlqZ3Y+ai9Jkr3QImNBZnWD0RehEth1l5ile6jw
Ao9iCBXLNqvWZ5R9ngh6sHRsPX2PlHt7cNCbVF99Qp1VNbDYXqtXpq7kye4no7wT
M3WVHkdAzJso/Fnw1YXaEMVvTzFAxnFlk/m5lXfC6INDNwTQPCRcF0LKJVddlP57
MQuWjaIKfKXzgEXQ4LZNFQp/t/+ZdEjNY+9zL371Cb2OEWWTHw852EIyCS6WLPbJ
yyP3YTguYOu6Q7mR+cOmLunfCaUdTAG6x/93O++DesMDiLmY6MZa/2PXGuLNqSU2
p99Pec04apTqG1y1qX4ZbdDy9vz0fzvQGGY5Jq97PMFOrPSHgaGRBR7XcC9w7Aki
phTYKADmPKbMsbQS+TsDDvcTbZdLhM+snqc+GdZPvCjD/VGdw+rxl/EfZi9xi73x
00Y23xrVhX1WgsAb259RLKUQGksPEmhMUUoKZ9rsdkx4JsUgYCnO4WxEJOrl8NFE
PErH8xcsjGeoHxhk/kIZKalQUxhbp6fR5/Lp2uAJhmznQnyIMS7Xsegl4IEq+EsJ
zX8Kswl1jN+pidtV0mZEA7S/S+5I1ieLZbUmJWpj3HAPscbGbadMYvc1x6EpnAys
XwSQgztD0re8avQfZj1qi6SxaB8QSK8wb4tD0xjOjDHEhdlofuGSn1CMJpmyEJmL
xK99WOcnE9XzqWrQMS65CBolxVOipF5BTEEsLeF2ht+irQIURwwyzfUNoKu8+Jl5
1FTmSkBPtWgIdzmUtCRf9VgV93yhaPi5d2MQ4ZjMpAGAwr9tgS6AgE0c3mnbWD6f
niudivrITlie8FTKN9ATGdFVrsLlR2fLqPL2QKgl8mrlWXr99SNrSUXQ/V5fNSjr
Pva8LtGgO0kFX3YhKG0/FM8sJXKcBK0W7zND+QhTAQyS4F/KGiVVSt+Zg49nIivc
o8JHa9BtfP9ERGSGdVZSlmyrgUuQMgCOTiWKHRO4QcNbLYuzZT9wCnESalC7skQK
coRjZn+MJ6SMB5xrxVMrzlDMDisrcL8GJJzwuR4JqqmWOTpIs9+ynvbLx0V/X35g
LwCWYwDEHgMtSQxM+O0wzY8kovB85l0ycoYp/j9fAlb/mbxt8ia8djXmJfvnt2fU
VJDJCvLXvdYmY9WcEZTXFvWOSdCU75lQysDJyI0DIgI4NzGz//OhHBkqoktLnalW
YbrZf2nwN/9pFZOqf3j+h26eZHLlhtJqZG+pPAJnFPUNzlzVRGYeXXOZOjUR1llq
v3PU3FR6/gYxmQn3s7CFXj80pvb2QxARFH3hy71qqc4O0neqoWuEHHJavZqt6TNu
tzXvfeKmoF/XkPV0DRAM3JcJLTnG/VDr5yqaBd/MKxc7BP7dyU9Gx6FTogC+Ez98
Vnk0MQjpQGLyml/zsMzFoKHHboXbG/zif14re0mPlu0pn1HIt5A0qxgDmFchAXRr
6aJBQO3fLiIbliawNJrvB08kZF6QaHL7DHDnDuSOi+wVqLZmABV5bnDuVVDQbTTi
ksTJVMpi0I03PIwJKBHrokT33O+mPUiLQWQ9UzodLURZZzajbG/47dd3ewlkPN6m
FR6NoqOVfUcGQrkuvbrc4ur9bBqri7yjVfb8RR2UdoxbjagHMOMqA8ZOtxFwEjWA
ThYpvuzX5bKnrllfyXth66rX4zOEym3UWfp1wgZQwgfDfU0VOGBJp0s5JR195/TK
/WoMMPdnlcwADIdpqyJ5hzkyZKoQRMGDJxAjQyXVWkLgt/JLcVplbkl7OmTI9ocm
aDob9L42XAdop2yho23Z34e7XrkEUogwVVb0IiMdesM498/YmfUnGx8wJ156xYqf
LVpaw8Gk3rd9GMZ1Aryc2ioeUBinE9zFOLYpX7m7m7EYsOKSQurvMmAx7c6sHh5z
buWUmTMPSiwYCSmRVm71szQRmnfDSYWCCGV8k//wZmDzBAWMkLI0hI1AdLZOYGfi
nhaQ3AdxpXJFVq9KN8YBPVdrglJdthYhYflkFtzH8Z1AvfsNp07JI758Ta+dYYgL
PR11BTd+wfMJLE4ySPfk7B9nkc07OAmFepTNWKWapi4MOP3Rui6fl7gIl0I0MzmF
ghpsK6LMF7kzAMUDBczmCW6iajWXIVZGtI7y49DwDdIIxHGpcnOSS2QMLDTkgHPp
6QlQc5mJP5+PP1mh5j7rlFuV1yEq6u1NwHZplZLh7+84a/a5agYw4adjG/HA0Gic
eN0IqIkDVC30RNjcAcAjlDH1rUUMJ5kAoYt8Rln2NaZJ6pkzH8w6Bhe0Z/zQ+YHd
jA3u9c3R0lSFvSqHns8d3djesQsdGS/DdcSiJ6DeQOjDfaiW72qIOPwBUd5fncaX
8WBmMhJ/mEbHjf5A2wybUE+zxATBU10VDSfxThy88LuRvs66ElRbOVSexc/gYEDL
1yuY7f4MspTKUV2Ni0ndBkpt9NH25JajUJCjD9mNhqRWTyqxJZ0feD/f+dD/JvdV
aJpneJbWj3Y5RZccmcHvNmMFHbNmYnI5QJZ9PMIhvPCGXu4xuNqGp1E2cDDCfhEu
UNDr126OuHjmxjypVmi41In2edqjBJj9BUQeoPqLNX7R+AMEF5Fk1/14ORaVNQuI
kcku65sCpHb2YzlcYghqSl70bIKnKU9L26I+SI7VQLgK2AvFrC2sOsfZ2sVbH4Sk
mG6amy4jwGRpEeURQcs4rq1KHsWB5kUtL4a0lSLjAK01sDcY1tjplA6Hab7MOTLf
ERtz24owFTLO3yLLHBieO8J7dWpSF1Rl5ymuTaR4znd8VmfbZ+/LJCC80Pp1RD0G
IIjyj3KjbTd3N0ik8WdwAdz5EACRPh0Tt+Xo/97CYAyXZnyLKAqaM5CssRRpK06K
nO/YoenDs/WsI6mtO74sr1bKwuchYXnVxm0ob0F7kHh0bvLmStJGUvD0GnCTEdJG
NQ4hADxu/tWI13T0LaxhnagkzOFPaz1HRIkai0qoJi0inPCwezpFTeb5YDsmyEbn
IiaBDWSBTZ8RoYk3ANyPhvQY5d6EhQKKLq4G5nfRt/7l0BfG/HxKWIJOGaOSjfhv
Y72XGibBahZKbDmmPhFtw3E7/YOvbEip3R4fwfsWS5QR/rIXHb41DWqXB80SK74f
LoidNzsj91CZboOYVTVSTz6BVX86+/8gKl6d0WrOtVzCGQXEQna+oL1yatd9cJ8u
jHwsTJSzfeHUMWRX81vrieICYS7HknNJhKaPXUb+Zs7EEGxVnuzyvTqr3CPozfiE
Z87/vW4ZmkKJYjeLswhF694/SpF/h4jlIT3V3rC6nKA91z//tVVcLgOQwtmx6qDx
jfOKYLeyT+0Hnc2arTLGg4jDjN2WPtPQwSuNOZ8HeQf7CdojV/Sme8KmgJA79Afy
ZmIR8308p3XU23pEhehQqhM/A8JeaM6lTxQr7Yd8zjigtPQ3xNLDnUUaqcf1Dij0
XKqQ7XmqjHTBjkT1g+pVwFWtR3lnU9jFjaNfKgmPkf35zt7UFNLMEipfg3Uzfy5b
ysNAar5n6dXtLiZCHVDfZTWoEH8x/nJqOtsJPXUiWb+NLhKF/Cy2PHuKIWhzCxvb
zU0KsywweDdk0+szl4pshPJI9ot6/uQicm8JArO1VXKDkIYSC1ftGY2mBhfT7U5Z
oFoWrCoit20Sy6jKfNlj7uaIIa9znhoequ2vXA/eeRBg1Demq0uR6KSNg+V/V2la
wPe2+VDjWPSEqq3DQhB/q3xBRRxg90pjaOcaMBgspDjGNFQUQC6AH2PRSAE3fYwh
l+tkZPH/EXPkbUq3Afi4IzO9M3irL0oKOo1IWXXqorheKlu4dP5F6f44CGxFo3C/
iKRB7s10i+8h53NNF4XC3GCAEmtA9AqicuSkWlRIzULDMh7AOliA2FZDMxXeYXPO
9PS+ObeUsnKkOQAEONarxDjs5FBsxnT8p2M0i3Mk8tEn+Egf7+IxAhuIsHq1qDR6
23/67vFQWZrQVgwR3zAvoD6eJUbp+H9a+bZLbBb07OtAHe8i4Qlv0Bka9edLuOcx
+Diq2wVi3JVzHgyqNX/8W8EOx4xMttBaQPNy+ZLTMAHGComUHHxAXMJX2dr1iXAW
2qzZCCoK5r5RrQ3vyJfo/LksA144V6Pvn5yj1D/ramo7UYAcKIjj7q9oVRgi4qBF
kVLYO+TtIn/PCw1Rmo8GzezbxlzlN++d2wPpCp2enSyeJmoBkPfUBdae5zCinj17
C5KGxz87wDabE15UghS5ssU4HIF/p/eNrIssH5sYacynNoRfWKb424OKZdYWUZq0
8PE8P0/GWQh9ZqEJ5PTZe1GBpALDulTISZyRTAIQ3xkgUSpAFEuQaYrFs07hO4Pd
JSEJAAa6h9BdfznW6W95qCf4CURpU3P2UdQTMRETpPxKv48lyrwCcT0kgU2FdcxS
oNL+cHwYTFdamt2mGLogFr97OVNRWmg72B2HJ0moE/OP2DQ9FFujrJ2A1+1dpBOC
5NUNpoHYpbBZ9Cfzwb0AJZrr+G/iVyNU9sI8cdKwu6QM2xl3QGOATz+VW99dNV9i
UMG5gaE/nePRXNFtXcy1LGqw4Y0qxLi0ZamUtKPMZIb175QcijhAwk6uvqIwWX12
C5NkAzxiku0R8Cx59Tqj9smZqVT6HS4zQAgxxFqYc+7XXiseoGhh7gmdTXgBKTk4
j4MNVFk7J+YgNmg+wR+G4AGdj9YAPNewSDjk4tgnOUlxPc5HT5tu3V+t90pcRgi0
086FgioaMTWZ0sBzjpXFc4nVzzzOTXukbPl74UtzSGOSQ5aqn0N0bRQ4+EJl8nLx
HKxmbxGI2DkIYVDgRsbBPYFuA3jXMUB1At0T74dtgwspjYfz9t7hDNjAXlANUkk+
WbjRru6i9ww733UDhvFd2czumEkXMIGGbgEj/NjZPPE8tA0IdwRdRWp8x90qnbnV
cIYM0vsBhjV5g+aXAEDlBs26ActvKNQWyg/3fURSx4Fme4yZ0Asaltnvdz0tmSP8
YYLYR8Tt8KU147dkQsC1ujWMM0r5e4OKjgISrPu9DsSQ4OfxnX7jI4cP8qJTYAHz
HSN6zOZddex2o4bOM+2aZcnElZ+v8qE4x9EUwXMjLycFEGX2H/M5o7otmzCWZV7n
zgncildZs4VPWf84j1u+T/kfHU0nqccuqA5OQhkkKCSKkEnH+BCTw+g4fMYoC8Qj
XGY0CACTJy0+xKdxFa8Y/ZFRCNesDB2qE7bDyZQY/IyIjZnk3R3jC6SBQ0varWhJ
asGYTKyJmZiIWDaaMGXClgDDeR+DDR8XY+z1cYKLUz7JyL4wuGbrMJJDqzJ1uJDp
7MVG66GtwXwIPw+S3NMfyZuzPwYJ3GaE+GS3H86xZpWaRnPuKTngvmUpfuQ2uztV
XVJm5pXwpX1ARGdfKtiyqUc6caT7QsQTSGiaoQUp87Enp2MxfhYR+IaqVrlF6KOw
oKImHCHOJ9j3906hvda4Icya3rWBdkEeRVB/gxY/1mGRB4ofu1/Tv2cYVex9iARZ
IChnnNN8XrcFYpXtF4x88mQoNFQhFHYCzf8VWKbiM6XxTgufriGlrpWDAnGS+8pR
CgENQqrzM0MmNpvvkzadQ77WyozXSY7tceWSl6YQX3y8+1kljAngaKwhrHxuTeMK
8o99Jk9Di7DlDTEyzHnlqooN7reBTX/0bGxTpMyI8iw6gy8jgX3tbvGI8Up3lw7x
p1ag9cP+96oSEy7bFC1YMj5+akRpwcYuAXxOM+PZgKga3FR+pnC2vlxzA5+r2GbU
IraSVg6VpoVEiP43G7SZb65b2eG18wvwlBwrvz2TVNoLgmHPS3YwhQGfA+/H4iL5
Qa380f17vOq9wmAFa/nIEIgALKuM3Ti+0Im+691gahRI/ARj3tGFAHRvpwpjP4hC
QsuwymSVk3iFXq8pC7Y6gQuWLwcZykUGO2Z58BTptRCobDBvdWs4BeBR0GFUXH9j
8uK7lmoCiWRcbgfqXgmjJIMjk3lJ+cvJp/JejgSgBlPoxiToFwa1oHIG7bQunMv0
REH5T7001foSIRjCAIbR1fqhYjF4ReyZrPncmPMa6TkjSUl8sSxq+rZFanNxR61R
1VQUo1e9sear9Q1OB9+NCSOyURzOCOZDqJUWivLurAZdUI6N03L9+Z3zkO6yxGJJ
8x1QAvIUdNWoAo0yqvSRWTZdQNnpqdjrH5MgH2Jy8jdCvJ+Ao1/xwXJPEn4BB9HR
kxbVyMJgQB4jm9loEZlaKsFTX0RXa/E3sBNNgD0++h+T+zyWQKA5c9/lO+RisAZg
ZPirZEZDCIwggk3OxrRfG9ZRZAXrp3rBzXGoZIjEcm50xwd3O0hQQm1meZmKiZS0
e9WFM04zFp4cVqZadU/dMaksJUPhQmqwheZ425WIhm7BEF8Lv0pLVi5RuJLe0tf6
XqG0zU7SgwSCR4rRUurytWrcWKRX1z/MjVPbtXBs2mcIBaBlwQega82jxozGBeCk
tx+btx5bL+RS9BxavoFcgfO+2l2nRFnLwYkGgt4fUmCy5B7CmBe1aI/d+nvIWsA6
QdayJbSPiB9uu82bxACN5HT2mxQp+tprpluwX8VCJpAeQnLRBMxdP11NKLiWQuZC
EVLYJuD6AZQbF0nZjebhknKdodofzJmHj6Cq/M0+TetV6ZVt+cd8uKNSDCib6K8b
3YsF2NiknetpuuQB2jSq8XvrS7DYi4Mz2ALM3J/fgIKLkboNa77eI86qZnsrLN+f
iKFou60AiyTcoOJk87pSmF6KLIhUknPRuslk4Jadlo+S2UCDKP3Ob2KhWHWHxdsi
jhbMM0ajdHIm7MBoKxtKyPxdTvB/KadniGXeX+D+CyqXYfftg8TKKR9N8o2K/R5Z
kXxJEukX+8lkjiprw5gpePPtsow1rpL35CuCmZIW/lfYyF1N6+B5Qz/0ZXrX4Mbs
CMYznYNOm7w/JMT7zyUhAPZjL+XPpiWgp+7thzJ1ssIb3lfkxIO55PK9KnQ9q7m5
wmjiuv6tkVDXIlfg8gFVeRcLFss76eMU5/NNA+vg5YjMCnK7GKnfGZ92g1iYXyGn
y2mNbgIjmZNebyxuQF7D12Bjuka0a4QzDe38jWmZERWJ6krKFMBgMhMxNC991yDJ
g17YyHxcPvjhguTD+k0jZxQs9paVkaGruiKzw2OdCcumzC6BlSfwfv+a2AtUpUVa
ZzIPm5Kn9GMGddNG8/dDp6+h3So1+CImeuEgnxjNw4Lg6LE9z/a/trAICY4sWaC+
kVP53/mOlNgyRSABgw4KKYxyCOxXFr3gtlh9FKOGW4SqQ1UVei4hDiUcu8PCyWMF
dcFVZ+/D9BHVkkb8Ng9s3JhA3S1iE5rJEYup+OUUQfCO+OOVe5N0p8S60QOGhqTv
8sncCbmps+R+lDW9koOBcQyUmjEchdSa8pbrz0ly6z7K4Ppr82I3r3eYFqAQ5xNg
ELNslW4+OeoyoEaMv6JB1GFa2WSIjBnQSqDS/8i94eIWZmK3v+nOPeVzxqxWH/kP
2VVRPV2VPSf05w5exOjRQ4IoxX0GcKgnZjhOoJ2kv1vSsMeKcqnignRKCVzSE4RB
j2ff6zwXluSxFUfOiB5Dbxa2uwMJn9vHLIFmz5dyYjZ+EWYshioYXsjI3PJe/i/J
GIaF4aqApH8BFne5KnoLrD0qaxyt5YweaEzkM0Dxkfw+7bUvix6eVQSnMN9SU+Ll
8+6EOgZ8oSeO1n+co7lmmYY9nToYMD3x8n0dpsENI+rxatujC6A2yFnHIb/rZoWa
fCChfcoUexgvF0qWZfizuJAf4wFO513cx4HC8ZZbEUC0srO/cx2apaYIlwvZ3bXB
n3cVNZwyPR2Mb5+Bp5eNbEzOgfdZRDern8FbypkxF/v6Q9zWTj6QtZURFl4emKHd
DbLe8ejgdPMPFPUt1JbqdMiEz8qaFoA8sLWgvMNgZwaj65h2klwnd8xD97cD4Yts
9syV87AEmPmuIo23verJzBApfEWGAPtGkMlEK+YNGhcFGUDcDCKc7GQSayPriiBI
X3ZGR4K/pWeFIN0KiR0enbR7na0BtRcgUHzEFBeEBjmRRknjXRuDsWqr8ngwD3YN
HfDL0Dfghbbyp+hDXuwoI32dnRIfFCvSo2MxEUbo+XGbYu6UKSRSLOT+28yskDTc
VivqiJFNb9pwPiCbiuqHfB5uKG6QkMI9qb83mUoVYeNCJz0NPb1W4lB6WG/rumkr
qYTwDE+bZ0KVmNGHKgfnDavW4FwTVHlkSqUDEN+97eTWLorOagWgqHpKA5Qnz8oR
DIJ+TChnYhIk0ykHf4egqWQ5rN6M3D8yzhJKqGEfaH6P3rNUObUX2coqN983+34O
4iogphpwilbG88SuJtmkPpm0dz9lUsN4iLg3DdHsMjjUrGsYHcwP3MfrTnUTvZGL
kn2cYaEEOQzxait0G2caROE52pQa6whhFPED6xuFbPU9eNXYw+ElUOQJ8d9pl+oc
oa9bjPxkF5NCpEfp/H+0+8JrYWasvX00hYi5UTswFtjznhX0ZFiOfLJ4XTTXBMAw
zHiCiZifhZVsHWjkEHZL1cj1SJjOz3ygPusiw3aa8a/JDwNhyvxJCC4CO4RlEg+D
erNCZF2ZMwT6srmIPIpDrgU3qjE1uTDqY38zemFs8sCXWoWhomd2UpHZeiQ79uMW
9Y3KNE3BA2phThbrSgqSnYDRPJSa/5L/TT9PAPopX4jp+6TiFEP/GSvz5o3Mk5ZR
dv/bGlNQEaZoRl3tYckMrUlN+rH9HkFDnmzAqDU6GiHig+gGXeprX5sasgHGOy/g
uNNW6QqVkg17b4BZpu89TvQZ/b56CYgZQmmitmN/MsOpr5f/I7J6N/t4d1/9aB8j
+x9UwvWWExzH3+dgI6PO3robbS0t7PSosfyljp8Hoxd1CJhSpbR6SJEWznXfCWwA
g/3z0+A9CcAyh4wq9LXOtrz/hEWJohGiAxZ0z7km4ypDF0EcckWsoaUBx6UMTFUB
fOO3Jrp8EIdwDAxCNMKdXVSQTeJ1AvJWJju6mWO7XQraMgrwLKDktYRsdNJS+WuL
CFO4SL8KoBWuGD2opDrTyfokID7Z5QjV2LoThgoJ3NB+6xvVKii1VlNXjYuOZQS9
OrmVSHHjxuFxNcqJexb95WGaenIhw+Lh+bGJ++9BzZ2k0Upw9otgzF2L8veeHx4O
vU+cheVm6RNAWpzWztIHJOSaRPte3wr27ho3ylP1XLHk/i0y9NOXIyF8l4otLLnD
rOyVHoTOtrapj/Mx2b/O3gZtYfOubeerOwcFeVDtxfJQ6SNyY5+WX6FZM7ATFUe6
dKq9WrLwOvqcprBcyEai4Da635LlzO0nGDnOdQG5YoSQqiOcPdL35KzEB6Udfzz9
zyphXX3oAV07jlDjItZVN9zEjtovs6u16jYb/pA4LTQ8bDDoSS9WvGcF6cgPzgD9
MGE4XukrirQzMlA9o8v9f6IAsDw4Y7aN+mdrfvWLs53nKQrJwyO5UjdGNaH1h3ET
XP2Uce9/0dC53vHk57wlYb47AS+hv8A2T5TFuTYOcNmGhdUt23btHMSODoDy+xpD
vZIOgKazwq24OYjpECKvhOMIPlt602GmR0qUgNF9iNPIJ+/FoTuM3UxquOs9gPtZ
2avORBfcjEm/U/IdKgfVISNGZk8Cpv1mX7KeZwqg2cYqaFMm2jTu8g9PleNcTzD7
f3Bf6Cx0XxbtgE5oqUASfAxuZYpqLrgHWFBlBuA2mR952BX2BkyLs0SvMup29jxS
JS6PVZyRXcnRW4De0P+5lH8N7AIjLl6k9H7SEoq9vwO//A+OjAQs7rHrWuzVpOFR
/JHmLuil69wenp5X6UukDhAZxd9Jv/z2qlKqUNPs1MuqNw4LlG8x2iSlJefaQ1il
F4ltEJp2W5ySkX3xd4Ii+UexM2ovT8UTaUVpjL8469R/oXRfINTpji+YANZTFJyG
zoBItko58qPteVWUERshV+dZKK1vgyZuULFAiJ4O+nqVhE8kuQ2Cr9m+Tzl2jjow
BntH/u/YaMyrddpj005tsf1yMjrE0Gu5MZgqykaf9HA7OK1LHJ95rUrWhpQ9M02c
+KElBZgKQ6tTlCjucDzPDMdmI5SXKjduRw72W9Q1V8CeOL5aLkwtuPa3zcPJMPMq
HB1/ym1IgGTNa7kVlp4fzhpkkz81gzIDcopEh1IZHSqaiFmgbGEpqxbu1mc6QId3
06JL2SQR6WJfK2PIzYPnTndA4mjww+hW19RCknHcJexqd0QEgrjYTsD4IA/UfDF7
bBfFiOzkThBBgMf0v2U6QvRW/bBH5IBYlvsaBFXLX+Jji2sKCOtLMwKr6RnnnWh4
P2Z61/3Arat5IKJyjjlAU/X5wJ77JJ79s8x35wcf1HC9IDV6QALLvzzh/UG2Pyoi
ZQzXUTzon4CvL4a6g5MwHi4Riydo7GH91e0ekW26H6QaerImzXQLsRLmWDcA6nM2
diyAgRZyNxkgst57NCguvf5ShDaavRpzt+c8ZXw++qmL2E4m2nbHiULzGJkuZxFg
LvuCQUwbqt1xhIIntAm8dE0dIqHv21cWSuIwKSNWZG7HTIE5K8HwYKga4A2mdJ5Q
fQNdy7SKS5o3D6+26Z9AFSWvgu/cT2idjUXBDOEwgDOoDfNSB/HRYtZ12dhp4i3a
34eosZP8SAxAgZs/Pe29qcb5t2YRJ/EQNvkDbLfZY7P0fLII0MVQ+AAsv3mNC1Dv
XYPA1Ghf7J0JRyloTAv6vEE8J5AYOZ949sNPoXkF/1xK4QJsPHf5mVAoBfUfq8Ye
Z5CNj/xs/6ySNvfq7SJDb74WlxEfkEg0PoXYaDkFgMIHr60IE+UZ9qMMTIu8ail6
WS3MCGN83bMjkb8o6nuZG5fALRAQDtZWeNhkRT+/meUOOlaleIyJdZ2tWv6XNepV
rQh9LFkQZyS7kruhuxerUJajRoHvQiszB4omCbgg/djipjAK7R5fAJdIA1toWUwj
JLU/WIGcuFADkUReGjrwSt5tq5V9+AjyoAB+nS93KJ3zLxRzfufdB/cHiTqJC36V
6eHGJma03+h4JfZ07ZUvsJ1LqZTXUEfNgqskgfykBWx+9F++cUXuF4q3BBes/GWY
cwVb8D9Cua/hWZHWzcSgt03gGb00/WpynjmLBYLwEUfmS0IVx2kPndrwREYByhBI
R+JhK8GgOI18MALlxnM942ErvWoIs0xLJ5ylit7+w8+S9bN93YE5YQvoebqejSrO
9wB7ps12I05svwaq+z+46Oi7b14W7ISNwQSQu9J/mFIEbv9epsSX6jC2BPitUJ6w
NI7lOV/C9iKlUh78A4FzSQx1I/P//UR4OYQGDcl7z5YcDVjLAq7UMhu2QXubpZvx
wnXHrZfRI/W1DkmhIQO2eCtUAuu8WM/xZWwasPGQa0ZZIu5tYJWYYzgxQRTo1nAg
QmyXwYAzFbGbsg+JjnlpmUcGAew0NzPwGP+HBshhwKm43dyz9SD+2NxZ4Gq46LJV
yAuFjwFPxtAdqgXRvXJGBXhZu8u86jGSiDiP56SGl+ggvAMn3rCIce4Q6vU/ECfd
IlZVlESAUiakn8MoYHaXVzL96A5Yy8/B7GqUlZqt+5iUVKJxJYkKOVBPbP7Rlr6U
Gg5/1jTSRCn6FNSexB5Ptefh2j8KkN1kLuNiattmNzESES7O2Ie/gLMltbHZTuw+
bIBCFTIOcqMgb0bMJTHrd7ZX2nfTfdbXNUZDiGRwBVG4yDr+t0nfA607RFoDoKIx
EW6eGpg0McnbvXPtmcB+L0fBad8wv4kDK9bi++ejlOG+kM8qtV0c0c3L/62YVCsb
YbU4HiM1t5m8YMBT22nkeDANKzx+O1+IudDYnagmuzRhnulXU5H6Us2TPx2yld+i
D668sGUtEXxYx8WDREXgAtaNy9OBymuMIP9OtlJDjAYwIeKSDkk7hOhKeeb/46lB
znPgikyf1KxI0bfKp5CQugIZlWL6iVrcr6FEmBFHFaRBECZl5o1+0RmuAc2R9pcY
yEA4WOKYsRFvNmKrWTZ+xC6hYIolYKbP9Y2zJVc2camteAFoXTU7bVlgt8doBqra
Km2omFKH4cv41H9wp7FhfUlGVi7QKBp4kk/faE6s37tMZ3TpNnCa4T+qok5IUaAj
cXMEnFnmwH3RSsM/hljKaQ8CXaUrs8sJFmOdnjMGuLbMEW5EiEN7E5emFOuKESE8
AAXDr9leZOiw01DW0FrXjPQTBhdM6oYRMr6otYW1cHZOEOIJChM2Mz7RYmdtQBoD
sluSvLCDQ/vpD5v933W/FuqMtRAIRQ3RDZ33Mg5n7ZPSArrrrTS5Gu2qc4FY4FU3
cbsuCNdkKmB+N+kH3Ys7wom9e0/37+AonIPvSM9SP/8ME68VbBicCcHu61aLTGgq
uijndRjRg/k4ic0vM81OUmDnU8m451X4U1r+8X1qYGwZ1vj485/6LHySpVmfXs0g
4V5nhQRzSyKE45QlYnbWcs7FdCRciIlMg2ZeKaxj0Su4eDnWxQIDKQbmKHZC/sud
clFc92XX64p6iwUql0lM8w9ykQvcZEpSrSOginmcGPxO+wTkw5CWIGbPh4Er8kMc
+JHtI2izWhgF84A9h+kijWkv1HtNLGkYV8ikDkW2iM401eRgyUcclI2+Lyby3ymD
fgUTr/kalEEeh2yC5I62u1O7DtK6oooPF77AVuiXGPQkrDZUKXqNReQ5s05gI285
yHc+0Pw/qho9eY2VZPV93ORcVGuJ4i+jA2xRfrYgyv1Kh7w59MBrVIoR4JntRSGX
tPmChmSjqi+q1EJ0B3XB/kHXRhMQu6Qk8CfZlbsLDHt3/reJ4BuTDnMaeWS5yVk8
BgzppVo9fX2LgTVKQKbZTvWUCV88n0SQRR8xwQPKyj4dU9qgYJluhD6xmLW7jlZZ
ArwlrQFz4G1bsD6ifqv7ZhyvuFqDou+qEchgs6Q8IyHWclUeJLX2Fj0WMTqudNt+
l9m+nyhTrBzYYphfLE3uxtCRugX0ww/94tOnyrPBmfbErFGUaeZm39zWz6L1k0DF
N6GLacEmuTxgez2GVLI/7lAAh4EhEJXOClqd0d42fKALemKGNQEe/H33XdxBc1mO
VXSeVvN1UMbllizMKG46amsEtUg9FuCswnfQGuEonH1w0Vl7S0MBHNJuU/lNZf91
SI2IghJ0JSSd4V58ZUUST2gDtAvvw1wz6rRzBnCHiqTX60kDuNtG6ejeciC0vMqR
hOM8tOFg2kgOUV8ntG5V29o9QQ4kXeWw0WwKT7qI9rvmjeniNgwxKBy96zKic2x7
7EGSjA5KI9GYQ2NVAc8CfLDBFWn27ulpPGL6/phQk4nmWq/yl7cPjQzc9WeSeLYg
Vrd961GvgJ5VGeux5ZXype7NYfrkN74rAgN/SKDXz58qAzHpBA5fcSxTri/RFbci
ra5oC3OzIMVhucLaw/wthkP7Fo7ydFeDidEbsXECeg2QGANDvblUjPIfZ0TqBwi7
LGqID88T87MkpPPokmBtXmGyi2j+nsBtSs6n3EuBaFGTX/F0+JknoVVPdUIzBork
tRQIDP23cMKMx2O/mU+coX4jlRj9un1O6Hx5MBj2N0sKtGMY21AjjzffpavNTYW7
OnPBWKntzGp7Gz3gQfHJNTT+8nmLMzMvtzutZPqwDooB8AxZSgCdv2rRmdu52DRe
ahwtRqgMt/UadDjxQBGflB6DvlxIZ0VMJfSs+whY21jjjAQoyVIF/DgOgaAi3eBy
4D2hC3mqfjDQWgje4lXzu47BP8AspaA94i7Z8CkQrjMcYYQPAQyMTAzn2guXm9Dz
L1JrcSU/bF980pisE1ATzGtTm0gJyDkpvJ1KfM0spePY3WuPUBL0cT03ZCImW+R7
/hOlTGrwF3DOgOK/cMCyG1GGNUCX5DxLd/RD145aSckP7fIGzM7/rlq1/pA1Xj6H
fdRks39C026bgPmU45cBiGzKsFYErWkvsGdjDNvXGuD94IW70GCWOOZ7U+XEUTMN
C3jMj2coVe1IhIaQmJwLFo2csxeE+2Ny711HIG3n8hyGzFMV3mIehjiQ3gnoONyP
zU7T7DPFyOrHi8Zs2a5QSFrMlpCPPTSkrgDlhz26ZwdA4mrWuuwYpjEWVP6AnBHc
Y+WxyVYtcuR8IIaXrpaVPfRPDK9Aq/lM8CHal8fZpRTlQaFb0g1kgrSiRZouMVZ2
BD+P+yN9dxJ8S7bdQDUEe6tfa1A3OVu/KIYVwv3uDiOlfeKMqQywB+koZYMfjlUJ
rZsAMVamFRbfPtvnMq8ANzoNKY4aK8Cl4C6rr/cF2HP2L+RAXU7nvVHSsvFSBI+p
s44Ezb2WSzvY/dweZKxbl1cPO1sIf0pdF/a83lFA1IBjilJdZ+YsGRbwI5j8TSgO
WbkXqSvxQXALL0BSn1gJ9YVtzexLfzHt1Jjs9AWHKgB+Ps3eRob+qrAbO3/LYdKd
bmj4w1VhwsOVOfE/V0bzSWAISOVO898dmmOOAZILfBCV7vZR1byczOhKgLCigT+G
3yyMQlhJC0//yg2hkkrjP43p2C1rcprUFOwSLgO8uCtSS2jXJv/x7WDylBLSevoy
Ck4e8jSewozY9NnYp6NU+mzyukKvwcq3Fsh9z6p7tzn92KS2Z3no84jJnRdd24PX
Qpk3AzJSDvRHI5v6kSP/htF6MANiRXw6L+n5fa9u8KizqcdIQoo+QpkMOuXd0dLA
6UUrUI8k6/iIfPG5bzKf09RoxHQFns0mO1MtCShrBPJY0edQYl+EYGeV1LCqHrZ3
mRpgHYkZhZ7RF7Hk448iXw3eBxywLVmZN6xNYNcHHzCs+ZC+i6XQJD/tWTKJIS7l
d0jtvR3XW8BKGowQaxS4U+o2eefMCtzKPdpCvjiap0IhcvxS7zrYPTgfYuUq321/
xQaqfQwuh8xum5u7CydPOTAKB5QR/P++FRibGzXR3EAK4kEjmBSLMBphnRaGgnAI
jCvMISO6HUoQeodAG3Z48oLSCp1OKYhxXdjvME7H/LpF+SAG7MnuVcikr/Ov4Rhv
O/DgEU7Oy6UM9EOiCvGphV3I07kG5069pW+rGL3H7YdaWp89cS16CTW2TngoQowt
gY1Qq/7sEvepxco+gSNEewmPnvV5fjZdkFq6BGxiasKuN7jpffoE3gi1G4W22u0K
k1lz+8ujyYPPJEZZRUNJS4aa9X+KqaJy7Aw987dFaLTVunM3Zke5wQpmLLFAa6lv
TZxKxvRFh0gwwVB8WzRPaiRzw/ibqeUpYy6atlpGN7rJPtJcLmq9NjBaWho1dmXH
H/O1XA5uXOeisYa2YzExQ5qgGV6/D+J6/vw8LqcBZBMSkCl/do1UA5OvAcPLgu70
rtoiQnrYnt64xuJ2iYxhmewylYeSj8UxomsVY7aisUcpSqde4EcQnu2OPQ8OFmxV
ORVWWM65nowGvIIX7668Y2uWHxjwUVsB8Ab0lvrz1+X5BgEaIGdGWIIl/l6HIfky
dcNYpah7PUdgUCmHro6AtvwyG+MhqAWQpZLcg7LHzLI56dU0/Ff6lVNXA/aNpGuM
rkPdiuDDuSWdbbH6WEjDNGOZX1lO2zFbzMq/C6NjH5EYQokObVCRK1uK5HrdIUs8
iOXj0nefBJ7Gk+Rf2q4RJBMDGxzFnQBMJARPqGRUi/iLG0qv9UL428AKa5UI9HHU
m9rI+KeLnkSlxC1HYRY2kdAqq1BIJymjfutn8RSuFTMA1AL7NM9HGjNjDQWiWFXZ
otTOwt7MmDHLmkSfn8OuOCKVPjk4kW2uyAB9vnbeOoLOKUXrbnNfOVDlXbPMfYFK
scLdPGDm6AqpiI4UD7QdgR3ZX8ub36LiVW90McdfQ5orGHeBNmki3JTtK5JxTy0d
5JHPYBb4YFL7Bp39laATT6t/c3t2dpPsCPwkUhQEjTxZQ725QUksyjvFHcqgKvKa
a6mFvzQBfd2E+efb26xeE0EgRSXTtp0ci51OKWc0hfNM67vP15A6A5op0RILWJdg
1hAiCHaY/fDpDt0gggKDmU/vofF7ZLuexhbVnBUz+lPXUhf3EMn31kZifOg1wtQg
ogdw0oMn3yMMIgvUlRAu/Dg6deEd/+rnts8awDA75ZOsQGZ5ovutGgPTM1qCA7rr
obB/jfaPQ5I9i8ujFDtjCoJbC6ZPt0/vQMwBs8AggrnaaJ2LUEAQdQ+LGdUP+nZR
zeCBxFE6fzSIO4NFx5uDE+d0lpB4Oene8FAOhCiyvoz4DGcoM6G0t80NTZ+6qQ+5
sARBE3CeBP7poAdRc1zGb+v2ecN2ZCQquiiIlQ30Opj6rqj/uTV7kzcXV/ExtYL0
u2q5uh3JYhER97wK2WSRYd4vuWxSIJH7tmUMe8mUBMtxWvnN6TB1ARQXfCc9vnSv
KBzSJU/TWnDnCDlxlQnnZV9Qhvi3yV9Cypr2mpNnAdn3kuo7okqmkzZ2VM75x95F
qR3mCw1sm83/snl96JNfOm9awDgdtdsPWeip3j29FFsLW5RJVGmEc3zniEAUaflN
9ex9Go6Tk6SteW4k9ImtGhOsU1A2GtGP0I2WjGe4H9Gk+9DI1mHTsM+W0BW3SrPo
v3zJar38MkC8Ay8kaauE9XMj6xjt4vcHtR3drgdCuYG7EeGGoWXEHQBEnNbnb+NV
YYlr1SGgp5Zky+QnbnXSNi5hJqPZqStaGtNWiXlUsc2CrUSA+vIwODMvFaH8XqRB
YqiOpqCHIZASiEpWwKcYAfvaid6pJVleSTsuOwkT5aaaIMZ4ipMO5Sy6fsZmOVog
vBVBbG7+s+Xl9p1Tl2Gh393Yj8YBbpqDsXPUhEdcz34Cr3UYwf69vPxl/VNDPnWV
90jZGm3aPn3Bn2nzmLaoMwp5uxw67D6cMKkxnTvN5SgvFK1qTyEg228lqrtZm+Im
PkYIaQBTbpNygejsvTbrVEIfMLYvFj7/KEG0z3FFsTieqzIbM7+RM+V03y+Y7mJL
vvAm12mrY3YrbS/iLfjwcAw/IQ6JnuAK1KnMfcfjeLZ2xkPouC3tY3FjKOi09+fd
l7ac9/vpuO0tRK8hmvdt7knIhLOJ62quMNPUi44viOvIw2LvNwY/EtHKttncFXQg
y/XeJK/ExaBPd720Xem91mCDrG9cUWhfGpuybuDUz8nRo5AQvK9pGaYCf59Gnwwb
ht43NPma7P2+6YVb16WsfGqhTXzI7mr6FLwUtyCEgxPOLkvBjKm+mDp/yHLRjfDz
B8LweMnpbcNYSVkPIWjB2fSLBzUSa+wUHn5zAxLpxksY5W/yfW+M/Mho45WRJL5l
iuDP6tB6hL9AEqyLRMVC5gVexBnfRsnER6MG5yv/baCfUoBFh3UI3n8oy7/cPYuI
fz1miwgzDWJfAjSOtWwEz4RQRmILBhFBPdhSGyA7ruA6PIAV9GGragSfyhDsnTZe
jpLK5gblHn7vAODjsKf0yuHdWro59nSZlBsnlF4i236m6xDyEZTDy5VFWsdrb/tb
ubsfAEl12EMgtqUddXlOgi6TihZC+fY8p7gG36Zwh58pRr6BiBeHKEL8fzcIwDqI
yQTcQxf3VQyfXV8rp9C8XCZWPt9PJ7IzziSOryzSn+R43WoTpduZknXO2iPivd+O
uwH5FJ4OYa9t06FsKhgFj+Uc7NmVz0qURcZewcusx1ZrKWlzakVel4pT1gWWa1sx
fd9ZzFfqTTudsgPQxhr7LnwxfpIA8rs8dIDS5dTTb1VezVA/DOQ2cgxn7JD+8SvT
0L0rVDuB4qPJmo/BDt24ESSJHA7VNT4v8uFAR1Fl+My+7TSwGOJq45m6trOEsRPl
QKps76jZbrce1riFKo5kNwZySDMWOthQH1oepwmfGEN0oEreDGpeciOxZ89jKphe
94iVCAyvVVSD1VNWgM5Mj1ulmtrk+JgmBybEBedx9zw81A62RjeX71pkUBgcktup
V3Aomo41hw09mvryO1M3dcrsEA1eUTkABGmU6C5ewlHcdJDe+MlA0fqtWgVbNUtX
Bf6/lqB8r1SDam/b/vEAYOVQBzCoqS1YPWH021mhoAHTWS/3xTs1sh/JYpYcasU2
ScxRbEnCoOnA3NEywLbjHJok7uzScHec1FnxdvQEuUrjMu4Vb3RRRiZUy5+qJLPX
Obji54I4ehZaJoUePvG2FCn8NrDNtUVPPhVEom9CiWsQdQSPCMYJNkUaidK80GsM
oF2Ctt8vf9oeS5fdqwLtzNRbE7SqDzSEyJopsyD0tRfropIQ16hEFiumz1xvGIhj
9+UM1lvBPNB6hjv3I1yASgzw0lRAhnA1iwyHE/cL71CQkKQymlLZ4vUFIEgWP0yi
pye4XOTw0YkOkUFG/399nXIuC/0XewiwINYw7Q8MAVnPVQcqpRyRV/hGGxWi+DUB
KEy6zKtGgEj4xb1XgQFUh+oUPLHBqUo+afYQtjWz3lqNgBAQxzEptkZ5Z6lnmGs7
1oMNHaAoT9VZvrLg/l0IaZvTIZFC1NdbyOb1NREyglF/i96TxbGoNh4aJTpAiRkN
tWuLZ90QkHRTcTw1J9DAS2Btx8RWMh156W4pi8XHVjzjvNMYBkekzO3KtBEMNAJm
qtwDdg44/DgzHEOueGQj9LPVAPBJjt2qg08RoqF40Af5A5AKzBLjO4X6mhvVU/uc
GKHEDfUc4sCzq72OKhy1KV726BhdkVtWV4QX7pnbyukiSA/vdWwzmHNOGqz4/x9d
CxQFc4c9/Yi/Tjhor9QnjjoGHBANS2FzGWqWV91iwxy+RJyAgCI43WDYpuMJmIjT
7obbk6tPFyFPcOsFKU2G0HOmnqIZrHA+eq6zoQPbvV/xeEDANnHNPdp4KnPWkaIw
t84f25ohoycNDIxj5Fq3NfpQHy6iliRhNiIlYDQB2mp+1qknCjzf6gFmDVsj8e1D
2B2JBAECSl7JZ1IGzIsL9EJoQ2a8Lx7sPB5BSvHqfERqmmlOwxkw5ArlGVLhrE86
KVDtbTvGJouO3BZvs81XssLenFuJG6q5K//yhGCX7rrUZtxtpEpkCVAAFc6Ag1ik
OLx8WZ4GOPZfizF08yTL4oHUFVlYhcv9p3cc5B8qOfYrxdC3Cq8M5zJyrlkMhqTO
UTs+txmDxzCYVxuiinC0tVSQZ095uOk3QnOMo4y3flrJfsvlQ2njLGC1siSXZtXg
ijPd8vVDw2qUrvYQgLNX9ClDW5YA9kr0evIAqXjK0Xp1Bu8ZAq+9EFGUaj1pQNeS
i8CLc0lxUC2ulxiGWbBigoUPCpmV4oG89AoYfEela7UarPO9EVlIZBpQsvbMBioN
qazEAa+WcEHXDBEVm18D5iXguJSRJeGDwi9uFqGwIVZu8qjEQJp/2kqlN6HF/NIk
Ohpf49iuWqGASrOEnblcowQ9Jz3Gha+WHd5wrNsJZz42F84mDojci9Ob+gk2erV7
7qgWRcom7IC1aDmitFE0flJK1x3z225DT6a0Ywq45pRmKWlTC/jHYXylCmkQ5Cns
Yy/e5fV1mMMfsobyTW8KAby8QnEnxPenlmUVQoPWXs3O31W++0pTohfEDtyNMLYg
7n2I54CSYWNjxE4ex7a/2VJCT6nKcNz7xljE26EwU0BGiIhsz98AY2IhPAgkO4d4
cOBje+VjWT7b+IwZCbpnNNqDTRcua7HH1iDl204LTgLCsiTiPTJBU/pxzOjYttG7
0pKlDnn3tyjA+rsKZ+qhUY2ztYJKMH9LoPFAvIP4G/9FyQjYmjVKtSyzcg6NXoX0
MCjRYIW9m3yiccqE7qJr/v3YsYk/Cf3bWuyc6t90TPegiqcTsHiuCdNMEOJL0Rwj
7OYFoGl+GCsJPvr/B/w6iYUyS1ArgmstcEB+im2y7pTyJec5GuhSgf3UHAl8A/GB
VK74xeRHfILWRNni7JgZhYioHTin/sXOUqKuZrFjqNvlxGbCld9+vq4YWwr6EQj9
a16cPq+sv6t0hU/5ziJnCED3mmg8i6qgPAMLXX0COXA0m549+HKbjQTvdB71yc7y
0vbxQNYEk0ngp8r6Qxxtw0Y8sQxNapBku4QUAfbfNqONQh3LFvN/a6KDlwDUXUgJ
u2edovBl/U7L/PqJ8/r//hCxIHUcqXMlTmU+4rKTNU2i3mzhfnJvm9AqhHiaL2Y2
DDmvLc/HclUndvhDP2+A3omY2fEt7gfRXwFuCfYEUOCvbF8644WuYWHtfaNR0ecW
z+Jmn2VxT8SAd1ss3YJl2HCbHHaMTykjIu23rtt7YQvtKdbTQjSXdtdc4DRBGvdM
3aCMfGC87pB8xzItnTbECgXL3G9CQjgZdToQhcPCLGfZuSWegQ73CoKRgo3yPwXq
NCBpRzTJbTylI5S6mkCnHogNoUOVPGblHqNxYF946zi/MSgSA5tMMnQYo0xenHjb
gq0h/iEOCzSEGord6h8ImErnBBTO4ngmmrgtBvv06xeq1ENXDX7hi+AuDMTSQRYW
7+DfudULNGe8CmVT6WkHfQEppGqBSXr+qeBCmphVpHBRDhc9P8vYK9LFKMm1ZKDN
eN8agqsbtxr7UJkh9bX2DcnVK+guHy/wJt+Nc7Pj2zgmVpcufwBp+f3GE021WDYY
TNTwuuEh/fPENTc2n3EVEqu61Bn0U+OEu7LUznQc2/2UscnB1JjZ8NP2/E9k4UN+
9ajiFfKMm9gGiVrRqYkeyROWu7LXWbc1yfqzbcZXqboKGN0cgCHYwWx8UDOnC8iD
GTAXoece9+HfyfmaXn86B11KVJziYVf3IuDOQi7upytDFI4T9JxCw5VGx+Eo4mZT
wbaG6HAcqubv2YBRTk4v8J/oDzSxGQ8s7zcqug6lzWlqejDpZkJIZuAxsrz3tD1B
/6RuV7ppJ+uH366x6hrQpjUEnj/PBQVX+VtRaoDINjc22gKLaRPcHrohmziAyU2x
6fVKvVi5T0txBKKd0iR/tiAoYuMIcvg+1NHARYJXcwehanpR3RpL1DL2GruB5IMV
hjYCCRBCkJrurpjn/1kORJ/xk2HdDPeVNwDpOVJHbmc4ZIJLkPS+zQ2Xjj3q95BK
Wj8RgRAvvcHDwLRwquNNojORjZMWES64fB5X0qZurBjwW278Kt7qgs8uc+d38+d6
BQ+Z3Z1g/ZaDUD+uVyM7H+x6JY55P+kEFPteGAZOkKLgzfLCEK9p8NUS8Y0j+Lme
1bFzWryEEukWRwfO43PnJmS5mh1lcONvLxT0qtOlKFCFc5fVwpSyp0pwxxXVsQMi
JhYdJGAZXty/3O9SgAelwGxmNyGzvk3xR2MEa/zh9GZEP2g5Oy5XX548hCQMwK90
cqO/h8ZKPA1EaYotRfUJ4kG7kx7Pux9sMYzHvWd2U3nEzl/fu3pEqWPLaA1xV3Il
ibp4vWa7mZ153Zp0xPhvsZ9Et2HQQz3AeBLh1ZWYr3ra9Fpdoi/DQaC8uItbFrLZ
eo8Y9e0vqN9DPunKNjfc3AeleYveNbSOvn2QJ8TXns6oEv9k03mZWewmQdqcqeP3
nmGvutAiPy2SlGEU6zzfasVHvTKKumMQMAAWmHrB7JkiG+Rt+9EVcsUSsbwo2l85
c57+JnWlXT/wP805GoECk+L6PX0mac/4j+owI2VA3aUYmyLK43iu+hzfNy5xWlx7
8fAJIX/3/wSjLs89dDdIZiyR5LDVyh6bvVuzDKGL/zKUaZhbXAndpd4+jcBA36Zz
m6gD9oO7tBaRh2vSkos0Ez/+OG+1uZNvGt23vCznRojQc2rr46K6gA7OCcDEiqtc
xHl18iWkG6d/X/wRXxU1JTwmTtXcXsUvIxQv1ce/rmoOjFAGcdOs4d5TW+cs+e/t
gVLfTPOVwgldsD1rtSQPJpf3kM8nqbicC3WtN2wX5iJKiXNq/3xyCbdDmX8QHqSs
t0tVDBBYafdpsBAZf0T4AGnLfZpzqPILjxP9DgdMCHSVX4KAUFrENqJtD17cP66J
LvyHp46jGUfbLp4UGXTvvuTUzlgma4NW6YRa5K+lLmkGWyZePNPHxvdV+9t7Ho5b
uDWG0T60fqM8tn7sRZEBPL9Gc2sOOvfJPdYCwcPbFe8KL4VfACkKPsnZY8flEPvt
uVE0hyRw8KRc1EkAlj1XM+F5zrGY7K63hupVfOOwtyKxoGEM9C0bbVRmTh4QAe8b
3TekMge8FTg5f9qakk1ZrPDdlxF6Jd+V3TclPsDK/YgsOXRHGB4y5lGsw5JKF3jG
IDWGufNVMAY3kUt4w3J+6C4izs0QR56LDqcMTkeCXNl8D1D+/cSprUrRDXgYIz0e
iu9LKP8PvNR+qJ5r0W5tgBtD22WjJbF7D5SS4AbZx3bLkc2NFhvAlp91Y+v3mHfx
mFsFkMG9vtyKNtkBEgPVQm0Ca3fhTzPgQQJTCM3pX5ZaXrxsK1+/YM2qvyhj7465
KC8XvaTqgDHUiwGW2IQ6M2dgrkmGaPdCmnJatKZKv6lIDaossHoXTc3N2WXOQqHV
hCrK71touxg6DHAzjcIR7SrlHEYCoZ8jIGl4UuV2kLLoopr9eO6V95Pwb8zk6woe
BYnaO6c4jNSs7Ergzo9/PHAGCE6qvZv4Mp2i3/TOQGHRO9GvB1vjkzTtsEda69T0
wJGCcyDucUu0Bc5ge64HeSH9vhATqQnhVkhBBlHCol6DMLDun/lne2vM7kHYR+x0
3dIvTueOtfoegU5x14gjj+Zodft3j/RTsmRJbp6J8VUJo8w9iP0xXlyMaXgc/XOB
3uskvfyAE7u1hD9t4itEamy9Z7eRs1gkeUmOqkZDTQFuMQ1ek8OYyu5bFJ4Vy1ts
cHiId14lKZRqIikiE0NlrgBj+LgdW8CJAe7l9gTj7akhy+MfXyvw4NWBRGcVlm13
Wtz9w2W89kn561w4qG9ae2QCjCZoRCFiaRl1p5RlBVDrJZN8cSGgVCkD/4HiGsHq
ozAGwx0NT2SSfvdr7ylKnTaSGtsJ1tMs/FqyvTRIy4MIhEVm7IKssDu2xGvKzDx7
LWpZOpiW37JMQLUtzKWIuBHa1Ubdaw00qWaIxUwv8vOUmh4dG6tOp/G0vEODkrcd
txWnPY4F5e8rVnu0RxgBBvMu6lP/COKD8WTCyAVpN31OYc8XjX8UjdLDuLGGc+oz
jBQRvbsZ5Md13dPh5wu41l7AkZ8VrsIe+zvSkk/OjH7SGln9kxYUndpmPagzX6VK
2WwC+d7CwRyx4QJt0ec/v146R/JsBSLuCdfeMqyJE7KWzOFYc8YdzfpYaj3EFMH4
9ZQCeLWizS1H8Gz+t65eXMCX+ODzkxjTjwEVU5jdzC8ixJpnndA0Fv+YeRgcStYj
w7Z/xHtZo9kLLM8TRpQI2ZBZE0FhTPbth69Ak1q1ai4BUzv0KwcWvYgkIZQ9BuOJ
x4JST8dIMcsJKAIbMkPyZU5yZ/+KGe//Zzo6wd/eOHfnPnBP1uqePDwCmPgc9Zyd
iYQWKGTTxtSh5n7L11sBat5zy8FDDs2IbAKognp0DfTwSCea1hH/SOfTw4GkU15s
Ruy51jzM3YIT42TBHn3CEylgY/k8mNw8xq/4xU33REtBjhVccCtQyJDHfsRqWbrj
J7UWBWy1cbfk6JGF+lSjXq1xRnCgPqW8e+GcDEGAk/EXmJdvP/vk1Cu1kD0HJshD
GUkZas0rHiXT3+oMdWVVJCFQ6rVqFuql4nUjLVW+fi9CT0Nw/m7B4H60itfg6Q9b
VTxxhiJ4XryEyaWtA36KNiXwFasfVTosfh+PKSTc3JhIpMSGISwvRh80bpOP7YGR
yhpxYIC2jHlhJvMgA84Rl8CCBk+gilGG80r6fMBYB4EALfahr3f0OXtRTlUZZcd2
ufiDOy+iUmdkqlYDrzYtyDNW89KlnocDUx/+etMTC0WN6QKz8WXETPDxVcTl/P/8
PYPp5xGGaqHxt5HEepZej7inBfWhtemTL0Ouak5RwVpw1EDQjU7+FlbnHnaxAi3x
X1BldHrv9M+wx7oM0nNmpG79owtXwWiCVZKOMdVMD2NscxcHXz1EkM1UPPWcny8e
2WqibKHLCgyRvDMYfqo4Kug7bomR5RdWNdg/ahCLoQTPkc4FPIkJsuq1d4WvZXP7
FgH3S1/EMTT35VADvZmwKp9oYqrAPgL7ZSyImQmuUOZQedX2Fi1DpQmX2NmEF2Zi
zG81NIq7JUF6f1zwcro7MFDWbfi85/9BTZPVq0BuAwOpaPv+JPZSHuRFR7vf4KWE
avFFxoU6AjSCITLBj4Snz+hmqQJzSfRs/e1p+YgPIC/f+OqnZDb65Q/AG9RmCkI/
dmDqA+sAU6mFJITUb04PX71iavt+V2tWjZBe1JJD/74J27vDcyKUlTPYY67xNeWc
PhT1l29CZ+MFIl9AwH0WDqxP5SYaRFehWF64tdyhazidTRABNTgxn817edywYbWw
L+CnUErylny6uqV02Yf+8JSKgcTdwzXHHoURozhXphnBU56r942qooRWqk0aBOeL
WbaU7I8HCEc74mEIhM539Imy+k/zYS8WgIVCPY7gGYAY31B//qkXt5IA4iwtrEzw
AlZ+Tv9xK1hQY3g9NN5sSn02dEvORTdkQwjT6zduhW4xHRAxEtdOIEkvID+AG/g6
ZxfMma4z9NUhc2HRL/hpDgh3Oo+jglg0PHAQ5rt5BFHALR388SbTmNJhntqqpjei
MxkHVxdo4WBMbqEnViiG4KiTnkjtvBIt+y99fuNqEDPFnijeik90UDyhwO2nLBdY
xrrSWLoBjJQ1kdj5XxQcYYkJyAjMYKaNqC1mOpB5/LrDTDVY0lRVn41zY19LWn/j
heQg+D1WA46Tdhoqc+xo1J/p+BkCTK6P7htVHuK6hjVJRvMkZZgLnBaz7WfL0Q+q
jkcSKJsncfvO3RiK/qT4LWsu3U6JKYHIo+CDo9k8eAdpqqnBjDH9o8XR9TCXOY9d
n3z/K1TSCK4GoaypYafPbV9tWMwOdUAhjTNXZ/2a9xkRt0SRg3hzFsSxqh2kmbqX
YL3DadLMAGInjJvR/55L5caNBnT/cx/pU+xurZRVW97K8a9u8OBTLoy98tbL/Fg3
2nvzUHIgfCT0VUcC6o1nDqZT+K927GjP6Ev3EX9xdNwMTdwu0TxZI1TWlCRYi52S
My3vrNuexSIjUaBmut8ow3AoZtVOxJFB+cwiUBfQlSgBCZctCihc5f/DWuDvHmPw
DM1e39rV85dPXwSVsmDW/Aj9R0L4JuBTIoQIr/R1igSkNUbVQcwX+Z5t2EKuiNbt
dKOpY8QQjVW81oJg215WPai08cE0yfo6hTBP8ExJErY2dHIcmz/9jVJadHIwhoH+
zYfkhMUKkfD20nhEcA/+Twk36ov2yYfIzdM0cwur3aifeCnZyUEE5DWffL9YBzcj
mFJyoLcAxJ5lQkjv8i1w3XQy7oKzETc2SFM+BrdK1vAjv+TYoptWLk4HNzXZzg1x
Mlk87Itx0o9JgK1wHH/FbJqK65FKwjSJDFGr2Hor+dkzhomM4chpMQj/a3sgAuHy
H792SriJUFsEuNeAgVdtQojJCCrE2stIQIFydz2RBvWHabrX6pJne/J0m5VVh71P
JoVdmvVjoCAXuhXTrUAqE1INkEgRn8Hd3JZpkpCgKnadXytC8xvN6KQ+WZZdLQRl
cMbu7lv+vRoKufXJTsr1WBeGH/hAHdPCyvn6I34nDMn2Aqjysrp3AaEUcLMWnAeH
xirHs+J3ms7ZpZQc4xlPEq7W0kNDqvyIqlGb7sGzj7SJ+MOAV/28TiRZypt+x092
AoJBZFKx2z3+J0RGas84FX5BAyowaySaajs0P4C+HuBMoRxcG9q4owNUWwUPIamY
MgB2xqEYfDt8Rx8wt6t0pba6ip9ltgzdCElWnzbEEVmT2iqQHp1+PutiyoVdl/l7
ec08N6G9MIwZvUxk8/rHGSU8+qc/kMdBafsES+/TQIgQPQksCMUDCQ50cr9HJskb
IGanOeSSFzJcPIxTKZYURW4f8KfpHTqrMCKJow51SXVFZ8cAeePXYDEewqG3KfSt
iNjusMwlkMBZImblKn+zsZ9LwICQJOdGklu+bY4EAxHbjxx1m0giw0lHagJt3f1d
0XjgRo2xmpkdyNjLauH0gQHMuk/Fz8EkRmGQOIBIAuDUfpPWBT7+sbBBsLQ595lU
3WPCs5NgzY1rCmYrxAxBJFvGXbSk8h2/ASnBpI1vDvQ5fWDYXSKK9WRs7E1mE0Xr
7C68A+LN0YMEPu6laKQBznVkSI0PTmiCiTQDaib8yjwpI3EBYuc4GVGvj3A/pI4a
ugOfnTrgNoFbaIGkF6obVb6kRUFj29DGRwARBQRBDLR0lBJocc6yV6M0wGPBhMh3
8tmJfUg6HBJ4fqJ7Xep1gOrKEhya0pkhlFqL1MW/6rngsV8VFNIijn7NXq/ybc4Q
EKHOPE4acuyctMYtOQDFuYbmNhtitj7PjxQhyWnNy509gdHhgUn70Vr2hv6WtoT/
nV0/3eKRSZNajUFNr8ZqYSMscsZ9aYp4sealveXIkknfA7sYFfGd13W7oVVqH8af
lME3/ckpuQu39TC38QtK/KuYc6g+pfJQQh9nxTfVxonRbQgupJr5Fo9q7xCd1iiS
PVeoxEo+kjUkQvh2eCDBGqPHxPqbahZwnoknaLAHpMnx96qEkvoU6B2uOEL39sPf
mKo3xcuMtUIHLsz75G+4kE9VpUKOwq25aDo9QywYy9CvILFzxM0Q9E5E8kIINxq2
B4Aigv3USFJvdR3DvMAG3bHMhEzOJ6z4kDysDIZSyz6xDoYynAiBDIgq3UAlIyMl
I/EeoKVFZ0Yvp9AERx1751eibGuDk91fJJZwVI8RGz5w6GxjwlEZvQws64AbFt7D
jUCSZkQNCf7Un/D/AxEXC8r4Y0+iS36q9kF+aCm9LZxBu4133Dm8FWRONCi24/GP
pLyROlLoja9Bq8VRAIQ4RaOFfloElXcpoaxkYmDlG3EyUKQy6a0HlSoREfa5l+CX
FIO7LIGooc7RjJr+pLK6t/TZl5MEFqTDQn76MKGUbzSfPRErUeTSvGsfUJAAnKSn
E7XfjI9XbsDNAm7GStxVYGFO/8GY0Fj1IAVfJ2NIQe6yrTHHPOdeu0bjeopfBq4j
3GEJW3qql6WTnnFoYPOJAU7e47b5dExdPJgszfQBERqMIdNbr1afKJuEkt/nkB2X
fVlPVFraKvfKlUAS/rtQ9WRSCbSfylE9I4GFXyZtv0d9BMx4X6a7I31dIHIRlSLc
DFuTZokvEDJzpdU8O8o2CTSpWqTNY7BBQJtzs3xCHmxFCfNdM/rCCD1RGMrf5GQR
V8RsQ/YJ/6EIZX3vAVnz/wO1e5PNAAxfu+HENdEhI0D7qpXiUxwnxa4BhYKTrWEy
N/OF18wGQ2Ikw585oTzl3bxa9wQulQ47B1g9knObg1dect9KuD8TcK4OdGBqsmxS
3x5d7EmrRmgdSsaVHIN0v2Crs9irJ0kAymUwimdUkPeG9e57ggaQi3pBC+K+i289
iWva27gu4akdsjQI4lyu1iFEDelV3bZogmahNkBr9WB6+Kquh674W00BNXShR2PE
eJktORSsZac3MK9zWpfPREl543Ki5fF2+PtHOtmJZkXPSMSW1y2vIhAdMyFuin9M
qmp/VxIkIgip5dyU0Om7n/xzTH0vD7A7duvWbtse1UH0n49XRxWithU07eRzh9sA
ADsgGmfhV+XypJoiyFZ6KGLkoseLrt9C9VGxBUq79XXPsj7McMuPMGTc51BEqeu6
RvcnZHmRgH5b+jlq8rbVIXI+1NbMAhlnPF+lF3vWt88VFa+6lsT7wT0jnBswm0Dg
bNsTgqv49IJ+Ve9t24um0cCec3GkTsxc/Twt9gY5jeF4vFStbTO14idTgxNyLvwt
UA1R/d/jWcCk7+dQTz1z5fqBZVeV1em+eUmR8sLsQlRnRNJiIz3iVYPzH7IpW9Pj
TKjJhj94WmhEF9Xsjtz4OdfmY4MyxH32poy/zIpIgMZgavwqccUZcwEzvfJTbEqm
1j4yvHOIlLernPJXdyii0TyOMx48p6sBAdtA8F9NgUDjICRFz9csjU2YAbPvF5Y/
tGnRB8KJsMVjir2bGVH/H5lE0t8L6EvDnaKa716tS+2AuCEEFTMO3jM3VegsToVG
dEKP1istEr2uz6UriZKbgzpeUMhbRkKc49BEVncEuWPwFG+z+fDxflbiSaCpuo/G
xub5vbzkpk3dcr/kK9MBF9UcNruY+HolF/ueZM86Vr4mJuTwwHtExjIJ+jmoTCn7
Qwcze4zBIxFoVzANx8NkbXMNhJnNKfLDb7WcbaMJC8Xgk2p1bm5vM2Kc++8Sq0BM
k438isK1AyOUVBMALKE39qr48Jc4QtXiUgZ0FRyu+kig3FIDBzqY9L+3U3l3Ntnv
b98yrCpa9oTzKXxf/3AJzx9YaHvHUyAx+iaT5Lj5vpK6oMx3HAg3eRw+ZVEkBFt2
sWnEdY47JpAwiw/nBEF+ZLJealyf2Ut/kChUZg0lb6piaShGcHXoHlxOsC/qAD8b
VezDfDhJRwzZK1tQZGbqoH2TRTL7g8ozYSNr0jrH57snyhni4uanZCuDy2g4i1p3
OEEZiHdZdoOeLEO7tWGmDhdxEaBLtWDkKJLYJQ6UWws8IZNmcq3fat//LYV2HIK2
fobAzS6wp0FzCVb1xhRsi1fne0wD+s0gO42mfigqOT52vgx1EllrWOTDQMqn34jj
6rG0/b0oG+kQgnPlDBbEwhd0H5z/KEyfSWXcC6C1ks45EVPd1j4WYyZl9VrNrOjT
0K6TljVU8ATjo+1BpqiujQzzOOLfsCHMEfDbmybhuPgteOv/gnfm3DhRMl572t/r
eMUF3fKnROsWZckZgFNCLatd+ZwJT2WGFgzqb7AYkFQXqkXqOUPVb7JDqyhI8197
je7jO9yRoRoFEw1MDBF2deSdbfvje2+y1Jsi9aBcSVLekZYDkx9S7AN8bkAtJAx6
SVFcYwVAt9UKu+tVKN0xyxVC8I7U1E/Fm3pGZRYXVAbcxfNyeSjbstY3tq72IkN+
SZEIcj7WvcznKlmYrR2hTTG2735asTwqmcaNNi/PLLW6+DRbUNNLZ3hLTd7kDMvM
Tl6ZpCC1zaTXKK6VXsXSzytvUkNuNAC/uGOu70AvKLemYfy4C7DKBukKdUS9Q7bk
R3qdgnA9H2jYo4hpfEBCwv/ntB9hcrPLZfZdKNuubDyVvyzXMGG7iuZC2ppRGhYo
GJyCXjmXSNZVVN0/3U8koqDzgQrzO9iuezVhPiZr05GfYMLju89Yf+Dc6LmnEX56
V6lVFfbDc6yZcFlqog7/2ECNWMhWtJJLfVYVYwhgICAKl3EV0DgNtFvcTUs3xPUd
emlgJU7JsWyog8TER0QHxRfbeZsxkN5uPEcw38WRbWb1nqO5cFQCKaoxv/vh2qi8
KwJB1RvXVtfitKUKnIJALERDK54Z/82VxBptrfN66UkEuTbKHQoRsv3FHWFLzABu
tNX6vPExIaBljQOwVqLJJ3Viu6ha/lIEBPQwsxAaAdcZ6E1jjLc5UpIlgjJvxEbD
DxAqDdezwimmJshy1Gv8hKBO0GFelcK0yXU1WFGOPGQPf+/D54K4FLjnWJfN4z6t
tlxo1qexxKoNyRMxYOx9iBZ2i/8P0B4PycEx1V/a29SLWvV/bGh0YygfJi6ACPgO
2oT9HU7lIUpnLiHIcZ+yYofECN+mN0SQj/hA175H2zRyRVtPYhnOqWILJWeRbqJp
vboZliM8b/kqmecbFUdkwR2ipN4gs+1ImR1LXfCh7+P0kL46qD1XbceP4ML4fv33
Kl1fyso5FmsTBz2FN5eSVI9tSpuUpKQTrkJCP7dGYBfwtf00QP2X8EKfbhaO1SyE
WKbSpskvT2mpnBHAY0FYrSsUJvYLVqQLoQW7mMZ9izJZDrloJbaKkCLLL/lnYy/U
Z14opTgYhF1UsHChP4PxNc6bVYu+Xe6+Uo/esNarsgWxBVbjuaRs7S05ccKjVYYc
aL6otGcUFlzjerdOIQDGrsEDdSdNpi2NtdT+m9l8R5P3n7yEHpJLFHnGVUa5aXTO
haxiAiKckjqGhMzIQhBgo/ur1JPt4CE4i8Cb+ClMOPPdiE3zutRqDcyGqxgRWzKA
THbT/IBZ2wSRprL+MwHH9L0CzAQNTa52q/XpMh6YPAvcuUIT8L+W247NlH35W4h9
t/a9jHSczQ5jJcoolupTBkAIwqD6wNqgDTUGdl8/ORFCQ9od2WibQhk1n5wq3X2V
SiGyztfAv1I5MUetY+bzOFccRSFTzlt2tEUAbpM/IRUR99KwLKQmixvJ6nMYZWNI
YTceFphHrh59aCy6lixX9ecrjcYvxupGQbJPi8MJR9l+ei20V0MdCQ7ETiqd4xB9
v9X+jEaLfQs1brq78ZdBMJdArZoOx0sMln8gaxur5t4D++XbNdCNUnF8UiWdEYVK
EWEZK9NkUqIr1ZIJZOtAF+SPD3pW3N5GZu3FCBe390f5UeBYiaQZ+7lXBV01naKV
5Ngmb8wLolASeS12S8124eMdk3CH+Va319iNla9yBNbuPPPIof4P1fDNDSjM3qgJ
s01EHpkzNYA5uYyex4SkRwd2c+ZHM36yWvNQzhO41gYGSVdy1i/Sd4yA4IKItj3c
sWukE9zIMpl3fbrU49ZOiwgUZQoCCH6Ag4XOsk69FitV2J/m3elM0Uq801LLd9Vb
R6QkSouyax25yRzWbwbqDZzl4notNkLtwA8COmzPs/Hamthu3OVUF7bM5h/LIt41
2wu4Fsk+NA5flxjQBBymE8cj019mqkgq1jDigJilJ9x4QXBTgi7RT4UwCg8G1Zsx
XlkNSQeSHmsgZhfp4yCssHprINGTJ4491G5krRUiNY4K/1+KcwSMWQjPKFR6JoSm
/OrsYAdHr2DCRbcwDBnx0QGaJ09vywRhR1Uq6EHozdT16vfvKL69oJKDkX63TsMU
yz5sIzQgViBLAbrUyWUIbQPIyB/uOkuComKw3usjp39iNpNwcIvi0wdFrHO/MtoU
YBFqhYZYkafelyxB22cTjwy/W3MrnuY9XAiFV+eo4fl//AZ60NbNotZnRIEo8A0C
hyg+tExdpQJxGvVrgaFnLCy+GyMSxZx2F8CvPbPXZYRFZHEAc4vFoq224a7yfHq1
7clg6hGxGlqqJX6z15BTSPD9XSI4iqDINkYmriMpTkunhRAzCxup0aqGEfALHZlI
M8Y4e7Qe5TMra9U10gIU2dB37xCOz1YfJ90g9EwCVlvUhjkCyqxyFEf1LC9xaHv6
3snuhnD5B43Z5sFtVogPC8Dufdu9GjsXEzHXinpDgqh8ldHTJUq7Wqf/SRQSlmIk
l1WMjkpvFXpmofgr2YFcgFMtmNXHKesl66RFcRbHaoLR9cQ1ltAZ8KBxwpOq04SJ
+yy492Swd2LLtgF0hiSDXEvOai4TTfBCdKZo0/RXHmQctSGJqXbFVmXgY6jtI9XP
F5Axa3Ct3EJjEY6gt4YOab5qCF8P1iOf1eNu59hY3HZiLJkFwlaOaNYrOh4eQvTc
3MlWUnW5i5ayiqM+xwU2AJDPMeo0ftAi5Kd16vYfEBjmSBDSkrKuJyd+NkaCkxOk
abU2+wU8MgBGsH6ESUxRGkVsVfFVlDxbJ3TcUkO3cmJOPLPHvNpo+Xx3W4SBPbbL
xkLA2hzbYTixS/IKc1Us0i4xk8d675kUstRtVHoahkCNnzGCoN5JsPxr50+GR/R4
wLbAIj7MVNXrzMTOtTRaLZzupVwRfsnZz0l0yne9q/8nx8HMLvTi375u5UW2zAz7
7F8VqIDpWgM+8zKMm4Z59vQTbRZe3ka6BVEQoTydf+x/zZiYIjLcw4JtpmutQ9e5
Vxda1m443UvX+fXBTN+48hZSAWi52Ts1IbqWZtmLuHGmvQkik/UqpmYL5j3r0Yvx
VNCWpWGPZLWl8xcSQwGl8v0ItpFd8pQ4OlaEU2SisXEkNmsi5wXy2BcLVgPIZIz3
MPgJjHaC4WUtukh5KNHSUeMg3zctDxvFBb6IzbiHRJj589PhoRbJluEhrbIZcMAA
eG5zorCVG0QBsbyR2PFl8KnSUs84NKDrj+E7FupSXt8u6jtZYPVG9sGpn6yodPNW
niKvdXluCREG8bM819bA4pWQIMjWzFEEy8JjPOJfQ3vwBfaGgMRVDYbb0HqEVuVi
pRtfdxEVA7NAV1++NbmoRre7Fsb37veLMoNl/HbKsQ/376l8QIz7zHJl5Vcbw9Eo
jT54+14NcGPzIlLOGgYwWHpXcreMqtX6T/gepcr5Z18i3WT2zYODmeRGWx4sRTSL
KobXj8BKInYlV7apChB9aPExCxQkcpMkHAtZJiE1Y/9DQKlBGPQGY41ZzclrIQ8G
jgjsWfsiIH0RTsbG0uBhhUhVzzO05JXx+UfHi/T++PEALG5hV8dr/p1hfe5ERIyS
jxvQ+MS936LcqF3PD3Pip8D/UTooIZaAYJY5j5Y1Vppx+zhNz4rJB5S386lBk220
xEnULfvmX83Q0XnW58SYIwODAefurPBK6bV3m7++NPNCYlncD9jHxg+v7ipMhhjW
tAhaUpjOy2M3i7JmyfUaywvuIuSKOiwBXpcBSX1TdXU2nIwaF1/yhawsOfQbf2s/
YdtjcXFLB4jDNs6yGQGpdNByMKt3Csp1OHFex3wvQt14d68OWfTYAKJGErChIlWw
u4MuSh2qRb5fB0jXf3OI1D09m10qQBcrsFlvq+F4Qbi0h/82cG2VyFfgNHzZe0LK
cMuRNYjwNCZxMJwHzYErbYWVjK8m/hyk8cHbnG5ko/p+CPed8PQeCbM5grUpOO+d
cUC1yUc9rlSQuVd1nfj2KcqWQnC5QVKzDDTPt2bU1fMgHPZf6bth/TDEAZ6nQgzr
PKAaYIXfkzOe2pp2JypWfHR7P4FX0YW5HP1yFYbSfB00ilKhpIY80qVWPPQcxmPh
R66IH2EESgy5RxWbcqjqAdgc3+P5V/qrjVr4C8rzLdItU5v2WfF4vRuBn0gis4PZ
VfiJv56xj1tm0w74EAgK+M9GMvM/R+nvhjmqfeHhMxPwNcnaaU1tOqCxfGyDjjHW
wmrFsxzYy0XatjTHkYr6Nro42h8ulVuaI5kVV3rPV5gF36Twm9glAjXuKvm0gmQU
YNvjGzarEvTuQXAUAUA+NIImMBbD4JRXidYy76kat8tIcwGeoZZ3l2J3Ss1n8v9s
WA23aC5+qzQ388LS1DVChNwxdAXL5ILDeeN6M9jIqxi1war4WwfnHcqpATMcVioJ
KIpzHZS1pfb+Z77Brg85WijbZ0AkJ8IaDMDCLuhni6UGGCRa0RfTT82Gph2IGGYg
WuLV8BCDGkTzQDNeoIaaW9FUuSmIUTcp4qJ1SYFgP9v8FLvi1anlZ0sF79ChMHvh
qAzzpkq8q1Y3v/eHBaeWv2KeFJPMEIjcWGtMnrgJya8N+UZe47c6VL57zcGgw1Pn
wJzdBQX2mfu0oknYawARWRZZvDs/h1Qa9oUWkZwwziLMpBTwnlAPWvvkVH6GzvQy
l4bUXFXRGdakDy4e7oU8K5mFUkbSsFTFMasrg3OzH8Ky3gVM/CJ94u/gvAd7RWLe
qdKlxAbFbPJSipQdBUPnzG58fLsVKNaDp5pdezi4T2Fwf430CIoQDytdpX6jKs/e
f2EqyERpLSFEyR2r7tSHEJL1NQgEZCXY2eI3dLBA0pNnhqmpRVxnZMQdrLB+S0Tv
w89ZHSTrazBAm3scV4/1vE5yyqsiiXONLrA2jJGv5PhVy9QCJiH/RXD/uLPfpqAD
k1yEdo8f12M6JxNN+WLn3C7BnT1ZqwqBoNKfVeCG/OAktWF8Of73ERRWP2cor30g
01GzqI4Xal0jGkM2TdICx2YATG2Fgy9VcNN4OvcZsV2VwANLwXaovUoAvfnzB1Nb
zoLbd1i8CMxPwM77R1PByzXngym0MwVkP6EjSZOqWqU4yKGIR6Rt+GMtIgPb7qA+
vbqvDYt7hqdbsB5pCnsapv4yYJfcRYIamxE3U9uM1NseDJVWPrBKw/QQJNc6B7/3
ZS5pc0Ad7+Na8lvyU4tfG4w59Z8dkQ3atg3ShPIa7CfKIKc43BAdqv5KsyqABosk
IdDwBUP+Jm17NSaOZkrGvStrnzSi+tpEeWkLTvETk2BOLtEgQzOcfy9xNU14k08x
269c7XQD8lj1UUlCnwf9yXU3DLK+Vk1SkvKRm+uErXBUNpXdoA36pk3VUn3TzgT+
1zoTs36AU/jOwr/xQkQLEd5tusXztk0fPGRNy5+LZAK+wPmE0/rvNbtUQZOnyo48
WqFhALKfySZawbpdwMX87Akz3xiAJ6I5SUQ4SvjoEQ6qU9UZ5MBOcD5xiJ1ky6Ra
a5qpaZj6CsnpoWL5GcarT0jbv9cBj3t5Gufk/rR8/jrndV47hLCdvb6eCQLldg90
NqYnxkUpIcqrZBJS2kFKOJ8xruEonw/sbvzpygZ4DwBBK50cjRFXE1Q4NVbRGtas
Ws0g8kJ8qgSAQxk8Rqpnk/yUcAY1LaObcaYGEZegG4s8HILnLf4X5s6ufHF6TULx
WCT3dKbZZgQcQqnwoIzAs4UVFQvgbmtNgZ0hlAmdD6srLfwRlV9ehhLHLy7BCaQ1
8IKtGiv4iF3GASw+1yREB6ig6kadqFX1ipmV9ZlbkTdcb3ktX6J2UMJa17lFn5eF
pLK01sxeqGEVMUF7SSMN0pdH3/FGf+6/ES9KvUcuiJ9ddwZhqzPKAGl5XMfYKVhT
I7/q7RDCja6/UOAridtuiVkNyL9dJ6LWX/0y7i8RZWoNVWD4jx5Pflqe0byc/V4f
llOJpBRMY0Zvj69avo/WaKkjpl0P37dTpJn7AE7wgKwFhTPU6e9safk679+rqa1W
FJ5nwsXboj8q/rZDo4xm8js0IKHJexkwj9WWkRtJCA66Rt9YpDy7///MhxC2FCYi
Bb7qL9QZxxMlS3QU3ZF0oRfv505HbrvlJJf82DkumY0lLrbjoGzmp6E39lCiTu/f
98+ibyZNDtebuqrUS6qt4oxDFrGtUf/Yx/7TVPb3erMtY+7E8Ut7wWh9QWPRx3gi
R2A5XogFRfcUvao6tqyVBazrc4H0BfK9Lo2JEBxEQJtd15XmhqnoniIV+kKssYp1
AtywRBBreN3jYI2qKnuqJDI4k55HWE+w8BNXPl3Z6pl3pRN5orxAHIBOTDGHk4YT
LsUiU7EnE+sShcbP4lzq4mnD50AbwBKAGDYKPAHYoHF30tD0tnwYHh++VbU3DL+a
EmW3yXwnmGJ+VEZlxJAT3umzE9bsCNpLW31wkpX25Jbr8oXOaPJwqnnD11Neyzjw
xw6+GuLToA+ofWajuids1bI6owAa9vYy5dsptj/50EvRF9rOJqpF+5m16SC8doVz
mxumDDjcRalawxZFN2eWIApzsj7m3esmhwPyoj970bupbP5wVkOz2JSYxsVTBfhD
wekM/FSEvAlZ0WY2LTAAqfXa76/kkh5brWvbt1c6PfCVRhiENJWmNXiBJhZHEWMp
IXi+mZkC5QOUfwPJikIxXrfB7QJkLFfMUdMVzfhvA9jdCrsoNBFGGrc5FGbfYtrP
H7yDvB1AKHN1Nv5g7YEZe+t1TxdZkYh08/v4a+KUEPsJF09907mQhQndy5OgntBC
uLWmW+GTvtTFSJo1FNtEAgs/tzEIU4pPtVhyq5l6mi2s4OU7Gu39sOSLUUG1OQhS
K5bSHXrdhUan9AxQtRWOgTO7BJ+Ii+xyhwFnw27gjNcByQy4lvEpLlQip9XmKkUi
K9pDdW3eWqL3nFzkNwXpASNXGQMOrBzWgH9KgyLNrsfG3PQ/AMd+7wE1mgkfKQsf
DlqcJCv+Qa0yw6N/D1TpEwkGg4cMINWLE9z8Vkg1tr/YqcEXNjlhR/+kMWmAysaf
VPWaUjyAC8DhMq9n/P/z0LKI2/mwRSG+i2ILouKWrmo8ie+lxf2jYedcn/r4OqvF
k+6J9URaJU/kCel4jCKLhejL2UlrtSb5hHpkNO7WExBHGGOOPQ8pOxIp8730qwG0
PnidxdEpf1vP8eSBHfE0XfpPQUxuFe6wEjR/tMi2O+qYQlozTbqMPqh2h3APs1li
osAJHOGGG1bf9I6cUMlE8miarmDN5oprajtkD+FGJpHJXwB9M8eyObgfevHTQAtA
ZtCLAKFloXNNAVKM7z4gMixk1lYyFE0w0cALgjA9txn4rIe5DOSh7Tz/HQzcBExg
uy4O0lD14tI60xA/ZRBosMiA40cAe7O7CWc498g020oEQf9o7dozm6O+byOv7kkd
3B0jybfUKaVKf1FfMS2jH9Db6546JNX0jxPP2WNEkiqJaMTnBMPMSRgwRnvTNHzg
iKHqM03iPZF5ACAbsV6jF1rzNnrqNKQC7sMLwwA51ljmYKIMiRH2y+YtqfTULObz
NHsBAcxkPTtfTj5dCmecqG8JrGV6d5CH7H89pmihK7EpFlTXbr0jz+iK+wNm7wzi
l+/2t2GmritgbEqEOwDkhUUt8VaETZw/E9aB0DLY0/gb8ljwJ+KMFwgV3dtI+WBG
049ceRRRvyL5K4fFRm5JvYhTNLSog6/R3NsjU5jNidRZQYUn8R1nxRFzbjnrsbCg
VfPTBsXJ3pnJJJDXwR7a7U1z6YyQqxYEDun5xsmtYssyg/ekzaqsojIYdYwpKaoC
Z6h36nSSIWA+CuMwb9lk0/vX0Ne1J9lOas0TJNBoBJ4Dt+HA9Iv4B6I+kLYzazPr
mrGxvlxc/IbCZ6roKcvbrKd5HAvMZKeKamv9Bjb5U8AGq7+YZid+NJYZPcopNJlT
NmhUJB9cnv36xmu3b5bFJoGH4ogA8OCpxskuGOAZZhkaOIWBBvGt6CsheUymIgS6
Z0oNBEbUZCtTsI83KV98wDMlmNQ0VUrqqb0dmNApmR1iyql+lodifZpQs/JsG5Af
4AeKOJeFkXOZIn3dIxzp+cvpyQXs3RvGw6dzaS/P6A2XFWnobJM064QVIIx8HFnD
dfLobfWUy/vvwEzTmbNvQ2lqg8H1eGDItbgazmwHEFAY0FvHtWD1Arpg1x4XuKcf
eupwHNUj8uGzVNL926RK/59qvIaDFKp05Ql/FDSzSy/b3m1uo7sDI3YKLwSk7wQ8
0A2GZiW6UZZIuzCsg9++5KQQ4A0t/FXk+P8cJk8uhCeb9G36pUzcQgYdnAcvOZZX
6ev2ptv+fpsyGIzLg36ndGkoGw0ltgS/ivTeb0XNLuUHeNKkQdyYu+YfIJDdwHit
hQ3SnrqDnX5V0qHmfrut4HTCL7vWrCdt5SinZcTml8x+Lgjh6+SjTX+N1R6Lo4cH
K2H3TXggLH8AdDnZXDerJl81Lky+u4NLLtOELZk4Ci/sqMhOEIVNQRypJKTud0m2
5ujrgWBI8lO5Jo3R4WG4lgd7yMm2cClpkfnkOB9Qfcpizblruq//2PhhX3ThD3B4
2TEa5FFk9/bRKCaYBeLScKjZZO/GuQS/allURo8TlzPnHxHqIRBQS0+b3SciWEo6
zgmtG4WVLSRYEEHzPpeUDcDzJ8I620JGp+Ly7Fynu9oea5+K0iEzYWTb0YCfodRw
gAoaZuPdxOesXlCftU1bAphXDksDn8Z33xSKisPGQAvdNtfQ2G/P/rE43PIRaB+3
DLQNM4hUQRm2D5T6S5h3HlFtuwFTsf4okaMLY47PO6xCmUcdomlNtmIbSlEbj1r7
1X46/lIE+tSZWMsDNnCcWwrIfoV4dGa4+k+d+0v2PVuo6gdCYsnbkILhT6B0bRHA
Y9obCSqxHrlBwbx5jQ3QM32j5z3OOX0350D7l9Fyp+YEz03uP0sKLBtgZYBUP3mt
oSnaISwLVDaRDUMgWTxy1qWhiguUUQVZoSRQ4EqAe2f5w8b/VL542qOQ1Kgy8jH0
J5kQqs2+ve9sgD/R+Y/eEzsyeH5M2l6kC3R4o2lJ7zn28VZAivsVXOKRBMDnWfBC
O0K6TwYtJrb4IJKH9KoSsBFXLMZj62SjRVqqffYBwD2NfARrj02tlirEDZjHQnYD
gzXTSe1S9QAZw4DueyvbVF6NedLaZh9PbYOHAqr+RsHt3QDBOR8mO4TKQ3NQ/c+j
PKuMpbVlXfoMzQaFXWJkOnW8oEVqtmhXKHb22NM/RW+vQ++iUO6Xk77e2aQrBs0Z
aWSFLC2HymmV/sTkeDwEfWTG/wvQPJEWi8FhAJv2ii9cbZtsb/8r9k8gYIQRbMeU
DznL+U5xiH8oxPuib+UWizsui/bG5qKVSDYZ1sg58dGA2PcgCys4WhO7EMFAaUIg
/f+p3iJ2eS+BaM/HBT39a56O+QD+gHaJE4vPk89yg+H0W88VFv+ckjWQWmJyXTgS
Eaj3cNrwAn+HE5/oUZs7iffWXLTf0CdgFCYNPR2x5C3orED3ntBrs5KaW6XBk43U
JPzVEAwSBdbpXOD5UyVkzD+NU69qwcA1WlwjKQvQRhy0lswngfzWcKWCvUr+4Sn+
wuKpY04LPpvrkswdbgegr4/ZY27Gz067DwTBBiVuKx6B2+IDpERiBO7olaA+O1vl
kIwV/geLka6c1StWg+jLJd21MrfH5lQUM5Zp9aN/w3xWVsjvkJxZIYtgFRtlFS3L
aDZxs4vnoi4IxKkHOW4O1kZTbQFd/p7pwNfOnCh2m9DqCNxeSuZgNlKhwS8Dpuw+
UNzw5+HEm8hOIxTTWT9yuAzQK6JMWQup+/asqwbxe8WEE3YFTT8wsIVXvcUAK6QJ
dSUuX6SKK5dmhkhp2Zqax+h1NhKmduIgA+QRCBjtSu260NfSfh7KXxQ840OVNZmn
cYpdVtL9eVhvAK9ttHJ3q14VHylUDtyBpC0MZvBYlfMMw7qw280cIdgqdSbt3W76
JNjokYVeAaplGbClycOMydiW/aRlZGAdh3+c9UiJKFHgsrWPI3CPfTTlDrrPN4jc
Z8srl2kTkChmF/f1bjR9Cpju/PNUka+nSZL36lvGiTycCffGTJqthmtVhKfH8x8y
01EUI5yr6lydgV5yvHEQ5O1nMFV+wZ01skakRZGr5UgZM6yv1FZoFpbL9IQawzpi
6I47FZzdMQnWqUo02/Hgi5xAmtMwjYzaLZYKZL7AJ4fuMIIREvCQY30KztK6BsnZ
bYB74jbR3DQSiCyELWOQBbEYdkTbBliugCJzu/MYgJ9whE8/vYywSb3K26NgaJKT
uG12RJ9DXPBGj8PxdUytnetttK8M3LD1K2vWB/ejMXy1ldmTnlPs3u0ovXFasJQx
N68S7DtOkSIP77gpq0+rH/Uc9Mk9iq1POg8PVWWfZgE2qkh4YuHUTzanfS0q3qEO
adeEbjMVZs5f+oxULBdbyExJWpl5xQQNYot6uxYvomwwKyzqgXX/6pGTuXSiwRkt
fm9N5Nv5tbIhoqywz0R8qlKm96CPdtk85GBAqmZehcdf0za/NAG1/LAXoLD2iakC
oipQsFfLJa3lqFpJBX83L/7nlf4/iDuOH1gQ7kHGWr/5xF6YOlrVQ9GXseHxXfok
5ZrIUEvCLu88t4ZT7JUWZCVEWxkqF+iVkyRtUDKggc8TbWldWM4xMHtdV+BYAixN
FHeMW2LKOKGRCZ+iI6An18CEE8enAnhphfnBLxo2r7VodDV7iyLTu6zNeKI8tZeI
qvpSP0PEa7BGi1SsE0h980z1A+np2X1iBvFPyWreBkCltb2R23z7P97AUK2IJFY8
DO/QvOQ9JSnwkc+1Oi7/l7JnT+xM4Y3k3gLiBbm6m+hhFXHjFMk0M9BR6MB4V/J7
Sdbp5eAC+VngKa3h7VJMFNFvmZMrVjzKNpSCRqSECgOuLZuLs8yVd5ICCFFWudpm
dwYIKeX4bztBr5hcE2Bq8CXvu6FdsHpX0eTuKCrIcqX14LSadHXHqedUo+0ObGeq
5T8rxw/7mDghm20ntPPiov1iYTJ7TBORKjvTMeQAVM7hYkgpCaxQjXuw1KuL4c5K
9URS+SlRc+LcrMVUa9GXkxIiwJ9Ys0XMxLsJK7ZaynSVYeZwVakwGC8IJv4fsfoc
7ISxRx2e+nI+QrQ49tM572F28qnBkP/raeiusKX7gp8Dq19OhPc6j+0Sdepz8JgA
9Ldgpt99BZTzhNsDsHREEoB+PQjitNB4W7lF4YpE6snNXNayjuoYkQG+W4OE9cZb
6rCz3ccA77awSbTZwdWd69l71/5h+KxU/OY+M57820ebA02Wi6LMxSXBazKuoiyN
TgqgCiEP66i2kxREaeqaQf/kaVrtBhlQCQ/7qmm8xDYgvBarsbAdwtLMdMrjCD1K
ur/ZI01kY8/BQgVwm7AbxaRtJrWu+GjZQQMS7u8ihwJqkk9cRT3pjyVZMaa9p2r5
m6UWNqKwBqx5tZgBOzxr1Uam1WBnMdKjnyea836a8FXgBTNpJwxSPl06c0HyuULm
mUh59cEXxVd1s/iUm//9edwmxvckQJKesekEG2mV04n6/jRtV4wn8GyOFnzDsLEQ
AmYjWcByh3n9ndKuFMYoEhvHKJvHFBDup5aWASDfCou+drShaBS+hDfOBDci2xqA
a0N/Rl401H+mtCyCS4tBgOnXfJiAYnWFleHAYDx7L66qdRl18L6PJIZ8LcfDv4Js
RqyXexnBc2PRRV7sa2isLCN7IA0MRKa63LPPNboVmka5jHSpbyG8E/tgA7dZmYZ9
hNfOjsgzb2XpFI+8V56RcH0kRHcr2gxh33slz2C9cVe1IKGENH23y6QqFSzET5lx
4Jx10VlgVB4wiTelyPaLeiC8qjEsVDaDzE/lIrsGKZVJaPLGJvxvBnu2xIkLFRjF
xugRKdUbqeqDaCuctCWXA3OqHhy2VFDbpSehKm8WSJHWmzGWEucEisI1GnuUI9Wd
97E6UFAPzLPwV23sEKHD0DHRFD8aVQqgVTr4C8etLP3aXcY+mCq4ErbN/QBuCYrB
OX2Q9+LbPr6B3nq/uU3i5uBqGsbmRReOL0KVjSoF44eimsQWD4yer6WgoR4/Z6Gr
xw7bt3pa9U9dxoVgr7wY9JjH0Sr4PCMOuTAAN3N+NwoausMidq5GOR3TkFv4GSFN
4B/yme7mP1umjOfdUrdfge4++yg3+DUA9MAFlLh6L/qXGkiYcsMz9o0j8ZFaHsxG
B6/fchDfT+hqv/EMismPZjM+a0EZPLG7O2gJObBZYbN2Wtd6Hc7HdfDX1EEfF2dM
cH9Rb91ui0sMCiLznkihVsZkUscolt/oaAUFbmOwgVpfO9BDLdSN0Z6i2OPMc/aS
6i14/SdNswU6n5VYcNAXOTKMgtUpV+qgySnXXJMjfzxiti1bFlyvVP4fjilkVBwK
Enjt1UByiAI1HDh7ZSm52BlDUquGyB/hntZGGfImPffHuOHkZhplRk2LKUgkmPy0
0MalInWf34BFtqU2qfjJU0/UFLlfeK7CwLZUnQ3r8gCS3lv3DIAT2QQLJcm/ZAy/
SLVaP3v8hQ1IeVL6e3S5srV4q6hvI5PxlesDcJmSeUvXDSPX74Lqo94Ap3QFFJfa
pYkTo3cD2jfoa4ertVwYQMZy0akoHuSw7VLtobsAeg6s6rRJEf/SoFuxBjkpCUgr
thq3fcfCzBxcjM1U1ddsBfWom3yf7zgNmCMy8/3bt+ioDOJ7+eyQMZJtm225NgZk
70CcEPoEJplNr0EsNtvkj2BOVLYbSqnFZoKliLgJaX7GnIjXqk9Nxtj4kJvw0dfu
leI1JEyqSWiKfSrIMxxEJUgv4tLgTd8LLOgOII+8i+TLpAR/y3ATuR7mPU3Cqwaa
y1Hz7S4+3cRRIdOmbjrayKxJXDLlOyZuFgJytjZ13diL1IT8Ju3k9xjou5pNFUg6
TTOBxLk0EegUU3OYv6t8TmQRk4BByzrXwlDZSHbkN8g+IOy6ZEPJU9XyBWLye6E4
/EtKfpcH82XNxvYKeFMeZl/WTtnIcQ1bmu6A8U6UQcnfaZB1+UlYSusIFNW0sc1I
GcxOq+dKdwzjpHjHEsfmG63kOOyfAJNwlErqk7FruFhTNub5wJ/tsYGad2J2AjYl
ZEsAR5Dj+gJ/lkt1mrRmplaUdqQnS48gRtwmML+dzNq0FF2kVh9kzhC/PN5ojdDo
20t8OUw9QZvjGzCUJ5UqbKaehd1QkgzBSzE7CEsyRDT6PujTGZduZt+TzsBix+/2
gl12FHIwb86KntjK4pkW+90NDq7aaJmn9rx4Q0tsKZ1PvkMNlcVoyGaw/O2wCyvu
CD1Eife/A9aurshXn9uI4d33LHMm4sz5d8LGuwrY7ZWXeR/vEoGK0I5hc9/4yiSE
PJNsUQ74V3TWr8x5c8w+9RQhR94+xhUBoVz47/aUI8xgDgJbiR2TgUpfkOE+rrNc
TNM/x/MeH+xN7f2f759UCfLYq+SSGSz5kG05fOYV7Xn54uliWGa5GZP3yUwdYc6M
dekGdjXmw/qcUr13xH/cUcVqUw2XM0g+TrQqZT4YEiWoHs+3keAYxc5uVPq52Keq
9pus+s7p2rpaxqDviUylsX4jLi5bzS/90OnvzsESa7tc3q1WZ6SthCYwKvWv65Ts
7cMBF5G3QbfFtDGGdC5tfaPIFCiQRtsd2OcoK8rlt5YbiyU79AQbbqsPxrRfj8jQ
XDB+IDmyO8D7kxyuNH2M8xXOEAxkyak26ENztT8UbccRASfhTX4Fp2V8WrbNGGGt
3WT8tGHbuoqu0cgTf6D6QVijszFi4sTRD5aqi3Cvpjl2oP55Tz4XsTwvTiNwDpf1
QdcZwnbW6ZXVbbAsy0DgCXSNEVCIK9xiiAE/ggGXCJaN2irUNIKr7FdBqFdjvVd8
NeecUpKgv6jfolRXxtQQ3685rYLF6F7qopCRGl0qtW//LgJnvoT5DvmwcwwaTFg6
PL0jfcG9Hf3g7kN5OYPuPeDj4h04jUgcJ+J6jjwsxzWJjjxzncuiDiKer2Yvr3lv
vg7UzbqMuSBcP63vfNzakctsnNvpqNE0FoEwku85C7+eokmzJaagtl1awl4XqK9h
RkfiFKqW+E1V9yqINaRLCfP0hBHaIhKIt24Cn38OoAum+nKUs4C79hypLyx/pZAP
//58f4sQ5WokpTQf+UWoqod/bgsS6ZKdzmdJrTPBOL6S9goFtbTUW3/SGLTGnYAi
h5XhoUvhz0DW9qliEQAQKV7PxEz440o70n1udonsP0SUHLLeWAOW71hQuZ+gdp5B
PYgb0UqRn4wSijzLyMDQvUmUYkGHC1Jt7A2e6fbXQAzA8+LqTB09WZefKZH8GklW
HguLropb04uUtcr0huwxjkHUEf+CLu7azgLPO4X0DVmCYQBKu53YkO2YadLWkIAK
8kA01GP4YVeaPpHruCY1lZBKKt4hAjNNFOk5e315CRqv5W0d9BN5nVofmZHcetPb
HYsTQ53z81xfOQpKhzFhliPRVAilWQ7TupTLEhYPJ9MxRHpi0In1AwgCPISfZIwc
Gk88a4z/DahCTjFiXmF8arQPEtJvGbpM1j2NH/2eIexs8GlosdPXJA++o2XwNyQa
PKCCqEMABXmWiQ8ZPeZZuoEb6oC+V73pActBr1pvsAXVaRUUiDOoGhUQhBmh2P6Q
wB689cy4r0n/4bI+KzGQNs0FhYKDhsP1B/rWQFg0aXrdq5uph0jK9uvQEE2FMsSv
+iWG+UMoS5iBqd9xVBdsAnx3Q8jo1WfwiRZsaBgF2wfa+qdKZAHzBYbVAK6FP3WT
i5IoZpAr3tCfqYZfzkrpFJVk03jpaxM7pK2qCPd0T94dsYlZuVSMuR9+Eb+XcB6g
TDdOJ2xPDXGXCp4cx7W1y5WH8fh6E3tYqMl7T0fyfEAa/+BK+tqo6YGnu6vpJODC
H5aJ85z30l5dGue1+ZriCeGHVfWXbrB7bFvp8QkvrUEuOEt/XWMLYoMCc/CQuPts
uX0JRR/2ISQxeJyhhHZTaSQ4bvEcRHL/2X0bI50CZrAESanHXCnMnbSKZl9HdAub
B1lOpMupb9KY/Q8WEh7meWRpFPfzFqPKxixochIMCEx6bzOMwY80tHbzI0LHdTXl
c9kfb1vFYljB4yqSu0RgGLJTs7ZpW+sWhdESZ9mHIDEYN2SB1qiXQrvizpfS69Uv
QjcTVRZZvrae6y2trRsnHrI0TKiG5ABL2K1kjLU7OaH4oylzzHSXquoqbZ1R6W2G
p0VvGqqeXyai7UP31lu3/H1SQr51OL2svt8KkpGBbj3oWk7Mi7AbMq+HmVo55A+S
n0PONuq2TRmRujw/X12Vf2g+0JOcTWL4cWAMUwBCAIsw09RDeXaum1ElK4yur3VV
K4S8jZTWmrzsr+LUEgpgs5QpLkZAkGu66OgJPQeeDiEmpurPCEcNm7WNPRZYIXKn
Nu8GA4jzHBeCRi+LDpAToJvhDlaE4+yfAKWlGQO8LnPWLSXj34aXB6/eP8d2crl+
TsEdru9zNlIsb7+P4lMsvOBcCpZu7z8aaOOLji7NroLURTjSz7b6eZYrj9e86nri
L2sL0CHL7OcWa+hXrXwAaHfktAaE44m8S1aXGUx9ml/X0jYNyTB59WoB6zunVtnR
to64Y6MtW4N42lL9Jm68F5DF2EqTY9VuL3i6ZOfQxyBOyY3kp5FvubJ7RUVXOAXW
7qm3PL305B6xiTnqfPKHSGJnE99/rnoBt5wqL1uxQeDtntPvPZ/YXVOrjeGjzR2t
4rYUi1eHV5x3RxTgDSinCsYCBVzZfZc3fxVPPlCT6lyEpn443R55sYRiKP4bratP
Vc7cGUG8YgpkQZ3xtG+7V79geBht6Ham4coBFwYt5Sypfiw1d6cxTlAn49DPZ+b9
Y17V/tkrT/NX/gA+T4HpCwJMkInIfc/zpVmQ2Sm/oVp6/07Wiaa6jnEMUJNU5N3H
w0Jgox3Bk6fMy/+0A+trbuvtMbAS6QUo0Jgwb67/uOZKQhWzkpTMcFDktTviitwJ
x6LxEfrkF1hzO5hz94qiKszmMOtauIJNRa/31nummWf/uJCBB7MdhTcZxw0lC7lR
sOUgL/1SCJsjlQSmjndVNpeQKOJsyRdWay65+sAsDv9BVoaQLJQ7qR4zsIcZyJEf
Lm/MIdXofCsUKb6viVuZFvTBSiFKG5Ekx1BoPFvrImZrkJ7lqkA4dZTQnIkHwvB9
ehVTL2OoxzHrE/OfhNqqK/ZQR4AmfV/gXAr4Bd24iawgqjKsBzhuMqOkPdoP8qC1
fM3OvC9rGFrue09qWgE8hQm0V6Hh2IrA7gLem3HwA1yyrH1oKQCv1ghU60KUSnfP
8qFseGwjZsfKDsTsLFzxZKmyRTo8mt3yHc/2gFhraa4l58F7/c+2OCh0S68EWtLE
5XasUUGBbUl2O9VXt+iRNTMuJ2l/qTBF+rVb/cUdLcxQcS8TYGDA4pQVkRn5u+kC
WknST8ew565NOt1V5cnkcGr7OFskmh9Jf99Ch9AxpykzofwWUztKcg3ZT1B70H42
R5pfix3Gjf6qkhVUu1K5WXN6HcMJL1EeQaUrYEexOV9GvYq7OYfwytre2D6461nW
82YFXKGsaKBtsiys8+qyiDr4N3nKeiqBh84GXYjuOiYGhmIxEdZxN9jnf724jOnG
vlktunUZEj68ZmJFGnnx8XXspIxPUOGdSyP0G+58qlYmVjN2dNTMAjCKQ1TVR1bc
/ff8uxIeuyjMp5zqzjNNsrP8xSr6EMWk9553FQfmMqs1QsHwnMbZn96VCE5SWgK+
pnv92Y4YdBaTNuYuTiG+0iK3RiPKNiLSy4D8YkvIeVLCynT3KhKfJ6r0sPwMxZOI
SjzjDxa3zdR9J7WkVgPSx3iu1sePWp6oeRyCOPmfS/D8YVRbA/hmg5DCkeL+cgmt
tIskdn9y4PhP9uZ/edy6D6GE0vYL8Krn6IhdH9wA7HRqHdcmrZ8e4Y9y4EWxBrzZ
ldD8qY94jswIuk9n4t2XbuwkMefdFg0EsyVEi5XzWv76ANV8e8n/Xw02vnpvQbh7
8u3PTouIaC2xMw65+IT1DK5ZvAJKQKlPz0EuylYaYosJiTm0RmPA3u6OSVTjC451
0i7AmdztT3Q+Q0mbGZ4nNdxL8tFjurzMS2uxUQ0bOnPNTsaYLpCkyuQtMzXfm7p3
PUtGsKSIrnEnk0XmzX1rC8UiB7motnwWPE0j7met9sZX7vIP0EMiIlYnFJX/xcKJ
k+ah7MKCL/ms8mrVE8oDANQ1nAHLI09E1nTsRqam+fwdExN3HZcCFw6dMXv7MGV9
GCmSTDeLJhsRxDjrMtDG46/jReaSumrlZ3a8xgqjM2cIDjKUm2mcF1esWJfd9U+L
KxK5OnNdPah9WD4TPZ+3hIwS4b1RjdCDAJb0U6bHqIAaMvrPst7xj/iN1iNEQ2WT
8BFF6unprAafr2MoF1LiT357/MThv0/DFTg0wuhpPVEwYGvHndNQ4Hsml1KoHX3m
ca9po2kuHERb8LYCi+v4e+UkmcmeTps1REoIEZuGE0Se6h+JoAk0FATvJqW65GDq
C5+FDG9T7rAVMZoTCROD3fSNZVJjfStgS+5U1wtgElI25x1WJH5CceWGFHDia0yf
gljKIcLskOnYrj/jQSdUe6tCORs3SbfOEMxktKUFgnqxNw9HjdYD2yVIWqDgyDlN
zctDqxav4OTbaJTW1BFj8NvIayLEENr9oNWqLBWqWjJ937Z4t7F7QvzpHJDvekPu
hLYf8GQ0vuVoX/CzBwP/3/rkGRiw72jQozN24oqk8ikqkpJFg7zqFjiVqoN9UWPK
mFQcaxBiwLLtaatyxxCMzcML2QLAJA44i+MOJImBeI+4BIPY5mVd4Sj0g5DbgaeZ
pZ6C5m8qti0V5sxCCS1fN4idhMgDQFZE0y9ssOn5I2nNKKNDzpJmICl25olQeL/I
U/vgtTBejBAg1jIZAsX09zc8sYnIcY6nQ/DQJ0efefwkDGssy0lrBs9qeScWUqmh
/o7Xqg/hi+CGlBREP3V0lC8h/5F/mTTw93bv2GdlO1VTloUG6MQB1KbEGfaGlKOP
4nZmn8vbhtFPdpcDF70nUBZXhieyaxG1SqiS6Sinm30aBbQmdJcdZ78cyuwrpKLo
Ogf1gv0ZeQD0qt3YWg74hX2aXWChfj/bVKA4XQxwvXuoEzZu47sgOdTRjsN07CIF
nfXV/3upqDqZ4JFdgZK13h5D2crjDmWMCObIBg8cZlc06/X8HEAKl6sHbPlXeSCZ
oek/yE/qH4tD051lKx03d8mtq3WOvCvNhlED8TSVm6z4VOrjSD3tLhhYRYT2vpp9
zOB4bm4fKhCAm0/z1kueTFSFuLZFohdknByjXscCIvUY4XkzZ7ktBzS/C2jUYbF7
s1kg6bCP3ArlAyRyHnXBfVGI416zkOqXlYJbIW1xSki/N4QcX7s3+dAFyFhdTuVF
AZQJ2C9d41xK3lVtXX/6JjPAyN26VLIC7YhlphD78ItYFlIrxweojlws7bti8SjV
WZwUM12nbxrYPtvZ/J84NLtOOaWbqVGDGsSpxcN7k5gVlOUiwkQKg5cHJ1Ok/60T
stT7WV/tmsY60ilZsxQs/El7uWhzVernPJZjTRP9b36Oxen5GVhuBLdoJsjdEOwu
+ru+bgTy6+ZarW8YuVizU57+8Gpi6YOPl+xWOJDrfC3jWJGkcOADg/rJmfO+kF0k
4O2SlwCbKtOjH3ORcJFzUKlJ9BtIoB+NUJdCVLOSu5dETDjb20q5BNHj/cOOnWq7
96KvEQzm1OPdxFJ22VbVFQPPvuCTQUsslInn5cTR98w6SYh7swcNo1gjtrNGbLQH
nV61EMxGYQoSiP7W2+CFF1w9GZ8lTe79wjRnTIhbbpAVoAAqOYHky6+64U91EdrM
KmJFSA8sQUaaWOoxLU0gMtBZ8fb7zyyB4fsalgkrvknRegA2eY55/SA4oA5qyf3O
F4+S8zxY+v+2o48rH8551ca8eprn1iTmm4isKgqzY54QY/FshA6Rmm3ZlG+H+bWt
BjlYajYoEdpEn4tjwKqRzRIEvx+/OF4cQaDUi9M/crrcsPfvDIp4wv2Fvh7uJeDF
8Ns+OeVtbQTxzD7fo/wwSo5/NYolNcj49i35SOZudS01gjqX0SIsz1zYPbt5c6df
91g2dqX8aw8smzFCr4EoUhICrWEG/cZqtEVPvAWB32ChHD1iNKJlVK8Ga/leBTXO
Vw69AHjPXZ6caFClOYFdjv52hW/hZh9gi5g+FOln97IK3MRKX7ODja/WnjFPpRy6
syVgh+ebm76gdsLO6VY+24xdJQZV9W8L7J6ljqjxTWuQK1jYlJI7I/7krrRX8y3Y
lk1H4kGkhKmELWR+gYdICv7HtrMNjNm6Adv+Hw9hnxgyebbAsuI5vRLyOk2IQZuq
JFak2MZ6pW1fxFEoVq63xSLYdOXniFoFpJvFGuGvk9hQASE4N3JEsi8rxaBNurhc
d2EBJColxrRjfsHuHVp96yx5qZaGtqgGK5oq9dwauwP4otBqLXnSqd/FPazSgpT8
FpmwReBMXW8wQTnmlZUeyBAV9g77vzZao8pj/ABk7roIPbNjDhHvV221RZFoFRfK
wk7N/f6JPoIEGBXKNatZxOxWeFM29Xm28HR7b0iWvFMO8r36xPZpUOdhWi9CQ2rl
93X1gJeAE/hWQsrqvHEXQ496QR4ViT1TJ0p4kt5fS9tSujjEbigyWUx8hMqgD743
Pw21eZmxBktNUaZ6qGQQ9hhii4Ks+HJVnfwKOjEXbk6tKyNogQn35VCRHrgXX1Mm
7/EXgyPHjGamBftPYKKz9OnxZ6gLTwLGEB2mSMNQGT0AJm9NXHmXjEZFNQgdC9Bx
MEckD1oBgm4HDf6wJUFn3GZQ0qLauTdQ9ixZz1FPm2/OQsmeAVWMOs9lhjM2GQXC
GDfI1wznq/pGADPLjIMBCqOv6kbejAF4/2BGFD+6gkGtAOApb1QN7lzf20NvjtYl
T6BrCrijBakfHRUWI07lnVQisMXd+oqvUNK5nWeiBfjbKUx8nW6C32u5PCiuIgFX
+m6GVe+hdVly5LxdyzMMjRX/A9QtvMLT/KvgXxOKHreHrN6YY9NFxC9v8bEla7NO
frbRq6lo5I4DBBQrEru4Zl7cKZZWbQTXTskmkj3dqsnrlgeQJJulkn9ilD9VXu7x
gPrKDj1XIfTPrCJDS+QzqdpXwUGGB25Il9CopeEuDRLaKJr3i6YZxoA49L0B97tm
eldhDm+GNN+o3gcV8NeLN6ge1GvJqTroztj+FpFbf38n4Jn0boiVm5+4ehrSmAFr
vy8LINI44AOV02yEqmQJRJj7QJx0qw/caozKNrL/i5rPgyJ+fzH0/fegokQlW6q3
c6eqftcM4puR/M2Km1kbih1S2pLDp2aTytleJk2yFgQKxHFnEjCS0J8qddi6ZJHh
pbYoA4jt5Dshj5b2pf/3IPcQTP8ye+T+reZTYB1xsICkxt/NMlhbIJB2Zhy9Sct2
H6ftgQ+y8duA+/HSBWsuTaCYln0+AxBx+/38A99TtwN2MSthx4unPC3OCLpv6C7t
NKzmkmNW1HXfProjnBLs93NuX1QwWvRlH6eNyqtqEdC8jQp6pm/jNuA01+MbLejD
jtVG3v8LyB+cyr5diqSNRg7+a+Klqb6qTHyM2XCsh1yi4j/qPqvLHQNh6DtcL9Ev
SpW8lmLfHfmoKV1YcGqXIHzzQHg09dsVLhrteg1eU3PnN8PKEs83ctUtHMQQW6k9
bW8GAizvHwDzcefmc7c9jL4pm5v9FK7Ha7oh1Tulcv0s3O9hl6H5SoIP3qS7do8k
MBuHyb/C+O/Y0xsezzdvA8EGEL8VX/fI4RFt5FtlimgGm/Vht2mMi0Wv4gLLr7qe
Sn5jdMmcY4y+OIpDf2Lq+pWyy7uXyhJTl808GmBSDGImAZUEVu91wsyArn+RZzKo
LrL0+mKE1TU0HEBV/H6+yZ43V3fsikFrJ3ov97fzWESEK+RLtzBQe8HjAy/zj/dB
fBzroGfeIHdvTY1GRBUNWKHaz7p+DHQf50qK0mz5EjhkS/DMJ4XirGofAxSlhryr
BdjV1/p1whoqo7HZ5rYEVL6xfxr+Tm+5JIg9ZE/0Kd8onj4en+pVRANUSfcVz7B2
EYbZeOBnz9UfDumuLmS4VumxEU/YzzwzAAnmbAWr9aCTBe6YC36eqoAjjCF+/j3z
4X/YfmK2esCZ8b15RcXJJOk8OAEsVcQ8z1fZjRi7rrwsVnu7Ggkqtdc5nWYwSNkG
j2Fj46Lpr6tYi9KMbwyZ/heRWWVQMvwg3l6jLsR7VbZMkpNm68sNZ8+UgTXKmfzx
TYc/4pU/OQlEi1cNJ5ZVomS41QhLPo8zU7ybLMcFSPxwrl+sa6sRki+F8uG9SCzu
GPehIGTUCClihnU5ELX346gEjkPV7kM6SJ/boneg6n6iGy2QLm8jfAPUcTFTgdxS
gQ/24QWijFtXNOp5KRHYESK79p4LodhtR1YxXH26GnlsTrcSWWpqqu5botfZ+Xaa
I9Dm0y04NyyIdLPf6PMX5FszHDrYH/QC2KmVid5QIH9SjBYwuYfJt12hJqlklKaq
HS9kk+OcjEWEVWNYRwp6Fo0/OsIpyBFvg/ZafW2Y/xN0QL7inVfOQy575yfyq2OS
yIiaAz2IQcEeEXBwz+xrzgVFWXySSg125hhgZAHICg9P37sc78S2WnA5iNVrsIQN
WrKLUPs1CYddo01Hz6xUR6ragEN0Ncn/KN+jpB0ippSW4SC8/UzaUMXa7hl3ZeCY
8l8LNxLr0aOJyo9WHt/liUlN/fLqoqueynBDelekoYmKBf3p/DYH5XCqNmbp5UVp
ANIbP6LPzYDVHcTKfornr9ggxNxCTluHv+YssEp+SPoBfbbfKxsbO+yh114XC9xp
hfflDdY7ts+eFs4mgS0jB+LuIlfIzJhth68uwDUHeY8JWCKhaYEdgATqw40C0y5U
3IHwrphzu6K58e+SMvzVmG9mjOKAxn41NBQtyqYOOah8JJlPCi7nWtrdMGpD4sQA
rQB9SCmZ+DdYI4eqArHnOz4A74Ghyi04LopWUDIR+cvLLWpVaoceBtcRizjUhvhq
9L5nqQC4McBTgiqeyCf4SYwkQSx5IowOVVF+tT8fhlAtEMYSS3L5gxUdVWajkXks
4uleridmY3DPhAmZjJl/z3EFPjBrfun0/eaz7FL518TQTZ30FjBvtdEX+tpjz+3F
s9fpKaUL16XgLSQn6xp3BTGZnogiwhE7KnBwsCTA5e/Yj1npTT4NeFJUY6gk+S4d
34ngcoyUYX57aTardBTMbeohBSUhE8MpaCpm7xQ7b4w+/uPdbQ8aex/Zn4tAyYQC
aQMeqvYRAUY37quFTBZGSREMbAYkMkYhII6duW3Gcvpz/fI5qfYIwKDWEQxOV5QY
RESGOgMphAV0WFlaBiL6YYl+pi/CBJkIvc0mAyhuagRpIpenLqZAnaByC6Kvdp9Q
gDENgLmt/yyDaKIWtVPLTqi7pRcyPN56kSw41lxlyLcOc29k38ns/Xh0xfatRlRv
Fj9uJIr0QURSDF2nkYPfYGMET22F0DNLULKOl8PnSWj31kjakZMgH8eoNRMuPqNB
o2GNuFuseO0fZPAMRX3frkUmdCiFAghuWklzKCnQRC4m0pkDqm9/OYUMzoS1DQtB
Z4zxiP+HCf3rNcjKNWzNLLbkUgcCPLpH3K9HjUKuHAJUDbB9UZM8YIJGLeAw+qyN
OgqdvPRsvojujFKSZL+dPIZxb1/MXRozQNqM7sD3WLGVGKZJB/UTrYbLAYFBdrmD
QBTCapN0+rhS6U7ATNYVwD8czmlF/Ne37rcpHN7MNzBxfLvA2I9V/5nycyS3VBKD
X5Uk2DlWRFBykwAlmT0qEKUCWTHUdCT6Cj9Ut65KYv4bG21p+cJF4OEP6GQvANXS
+CKdPBIRkcFVCadGzLIIu4HxGaRK8HXtHjps41/uDcEU6Ojn3acf5qADaSNRBwz3
p4c07sSVLJRO/n5pLUCfczKWz+CdQYL9Z8E/cRnDiYt9Xkw2/wM9d1hjoRwpxkvl
QJxc38wBt950MzK7lofJ3CDHozJnUSIOSPpOkjjCCSF5PMN4kSwb1+qlF+eMpu7i
nba7+AWTrgAZ8OqF6HR4oHDqnAJpfQdHjGoDRn6HcJ3Xw1haFsfuSaJseSrxcXWd
CUFzek4o0nD56ahTlVim6Y80A8tDbBz/JKauTG4EqCaQshdWBUxQznsiVe3QmIyC
qZa+ocQSPApwaZ8ZN2rIAWUbHBdEXvMxr+zRAEyC/WSCQuyk6oo3lRK2uPO1A+Nw
do39Dovk3N0oWpLQFY5Evsz/Gg3dUXCOxmLx4AsRfENavxTxgc9aUHEs87N9Jd1B
rVWc0DxV2fPuFP20Y0ssjdkC2TaGggMqwNVFWpcfV2F7RFaXY7PPxGoDXURqSYe1
vtP8kXwNkL2ro04OnxgOxGUnEPU72WGoR8P1nvaentlgwday5znBUy3ku7psnBpY
fKQxYkOjUZ1qTJvL7pHcnkWijGk0S6Fl7CoAyv3/H7ifTkbP+QvHdGlmhyzJ/hrN
QXtMRKcju2aWOv9Nx8CAKvVewW6gU1Ju7K17gvOk3RZEuRTsa+blf5upG3OsoPak
h2894e1rpKKDz3Pd4c2aH3DwIOceJr+xTidWskyrk//ehAH+dQJ1Qy3D5gbQaH+b
XdC+X+rJI/ftk2XU7Nt+pY28gRMUUU78XIbs6e8iJAxNT/TYIPZJIkZMuwJ6lCqn
DZs0OmpbrEaoYdc9Ar6EG8PFBW9KxUevmj1DnmfwGSZ/Lf1GOlYVQTVU9fYq/bmJ
XsadpGW+EBqTYiFk+Lqt7vlAS1jLdGyt3v2MsF4u8Z7JTpCxR87Jpr/2OBZRacnv
PluTr3rXzM5UpVJXOMeLhlUSpDnXe7cOzoWi5AeQ/5QoNkEgyNiqwUJ8o0NnPGUS
cB4ZMQKwtJ//m392ClEvqkVIFiznJBG7NSUoq/YGNWM2wL/UoLNCbERkm+o4LAKv
gq2ELZDlPl2TlV6FoZjZVfJVMFbt4dWQupL76zZkXTiR2OXYAoLbZFMs+tLaly+j
m+Ww4llqMBBeKNgoukR86kFhyfJXOiT5pgJvyrljdUL2pH4Jt9gMZu01nr/WuT4h
qxoKudX8h9zC2Ew2lhJp+xDkQpnQUgbL07hoykPpHVWL5pf3p9gUMNggl8FbD6HE
8yv50tzIkNnfzTpD3XoBabaacV3ilm7zOu3KhOGwji6cWF3v8S2fp32j4Jf/VZXO
7kEop41nFHdL//u555OR1crR7imkIXtGNvqMysHIz6rXT5fbzH2DIbEt2F3A65BS
LBc2IUozPeUoX7WtM6Lc6xF5ronIjPRlYkGaPmtOIdpbceCVGCp825vTH9OTJptn
pRVN/usKDQ2F3zwLWLEp8cURdlDZLGuUYd67pzW9TTuyoV+ApAPzx2EQ7suEUSRQ
xXZKxuaMzFHD5IkaccvPz2Ozny2NJyKSCiwTPTuXZzgemRtmR5Qi3MEtyaR0C/qS
SuRBkH7C1u/uT2/r4xNdSm7iYS6/hPK+4t5XnoxUwDmTQelA1aiB15AXJCgio4cZ
78GpRe3gr6IKSGH578F0DIjtrqyqfYzWqonPVSGVEybQGHSoRz72nQs9BEb5m6xS
9ujOgrI8e8h0BtAtBYMMYKzxrmAim7x4p8BIe7m/WJysg/T54VRycQl9Q/WnFQ6M
FiDNEfvMixgT2zYGhoYmNgv/Oc3myEQVucO8XmoNuvkzCN9Dg9Q8sz8MZOZpfsZR
6FOOIxnSQJzKBRRunYqTgnqQGxcCcJDRPWXNbW3GZbJbk3qZAV/oVLqftx3zdBiy
XwNXX38TS0YmCELtHv8CBZdtOgpM2mNcJjCeBkRvoCJ0H2S0SnCeX28ugupH6XST
vphp3Jstx7m7MjgfvFpY4XV3BZd/6mTa0hDrveCAqTNvfKYUa4NqzJ4ZZ9jJTZAm
iTRDHkYmtI0fw7Y8gtSn5HK+idP+pKlL/r+Jqn9SbLij10PJWXc//bume6e7dGi9
bYtqofYgLOrahn7S1VyVUHGu3Tj+s7cWq/lKo1DBuV0iDoFQS8mr6c/PLR3S7v8E
hXISyeqyioCJ8mUhF6wBD2m3WBnBWFp5TKmeU4gm+AmiqvvJ2gbx9bZsQgFA2eI0
TNZk9osyCJxaRoErcDbW9HndGNE+hyVJQH5gVUxVVTkT5phbAp4GomS2lSe21ppk
sy6qZcNht/XBAExjiXF6AYKAXoqJC2hAsytk0vfEcms5ZK8vf4Jj6athpnXI0rBP
NYMF0S5c7m+5dANgQ8+LDgZULOLFhWBHpr4NK7ptHUus/zxyyJ9Ql6foax51lo8D
jvmry+0vT8WSkFurPrJuaPP5h5AQ7Bqy1fXa79By9rLXxM7o/mgDw8hkjGUzHqjE
cC1+upyn03V7hpjZjyWAoIM5OyMhhXj7QhvAUZU1I0ay9F7D7lFGHNbaNZ0FUNSe
0Pd8Hazx0mlpxhiOwdNlILImtqmgLACX8DcFiT4es7p1LhXXweUWwUqWVFYttwxN
Vei/5wpZqRthj5yIDnz3ylWjEC6Spw2p/MH5m/TzLfhBWR2JrD3eKE21822CbqMA
XbdMvO7bCakd+SSMvq01DWwMj/nuO36B/RnUrseOcQStrBvSBDxb732YI7QxbxXL
tL73B+yIlwl4Q4BS8oHLYmofi/jdSig7GX6eNTRdKCVPdstIcR8JPJgVC8tgmaUy
AG5jhKp2nU0TYzmnFc0KliuXi8ETj9sublvhrWtMhMWZZ4vu19snFJgN1emP5hr3
4MzXLoVe+WpYH3hXSBngv5UW3Pqm86bZDBwWamYkNd4Ds12E6ZrIVckjvWY3HrwQ
ZM6b2cPyirRX3Iy34aKIrugoLkfY5e+3+EGrgWq9m0fLT6bWX1T+3GUk68oYe56A
orZEWmDq7mFuGeq+PPQXDbCQwybhHOJYWHEEv4wc0Oz2Dq5T9w2Z7gXp7oLjuKEs
tyes41nPMF7H9GIOGy/69hdxudZ+2DK1tGlO7ovRRFdAbsCHTriw2sLdI9Qfd8oU
UqZIwusGeG7QLlNRUnJxZLgcWkGDTCBQFISdQv1LMp8CR1GFU3oG5WSlJfGeJMGE
ZXIZ46e86eEsa5mKDLbHSzP9+LLJuKwEogzanOOgLPuGiWZG6Mg5GA98WRaz/W82
zI1X5DZeEk2Z+BpUiAjbVW0G/TRjBWhHFzfIMM0KGbCbDaqe1eaNLzptyJ98s2Zn
vMbcd8umAwex3owbnEraXMz0RiCi5IBrK1c979GKh/kKRqdMtWChvxYmC/59PyD9
HR83GDrnVrZYPQUg5T3IMcptnltUr1wYcc7WOu2l4qliWNNXqJJyNKnRIytf6v5Y
tvUP0DAyvoGZB92iMmv2dAgkDTr/n6mEjGnNxdnH1F/SHiPz6V/hLJvy8VracMay
UKG5kDafASxOy16apA721mJ6Tq6ilVl6Hcf3HvzooGCSD6H7JBxiPLe/gqcz/oU/
p8OKjoVyzws2z64pP/iB9uFDy1SgODzu4afhALonTXevYk7X8EOV1jnxZH8TVIQU
0T+62W0i0615uYTfYQkMGHrVxGnhigWYuQwdenVcyfJG6WlxSjYX1Mg42yfaqdvQ
Gafw0+c8MJ8N3NJ5bxqDAHi+tuSBEiy8ohc9XUvKtc7E3MHq7hDMBUYUbaOEyZPz
r5n1UWI4FDXQ31JVT2VbFU5T5WZDOhadgrzsvPifWxXC9plsatrCD+ExvyYft5ac
QSAk4OQomdHXNkXqxOBXZQGzpUYI9yKSik+YS126GhrHhDUjd0Xke7O90IkhvbSE
7u1xhcSBtuF+frVBKvveQSKAf8eesIuYc11M4xgrrxGNlFERCTfVPQE3NGawiw0x
VY1x830Awp8WwTjni8bE5GVprG4nl5sOlpYhVm6FxHRMLu7ikyVzSY8kAE6z1k7A
L+mX5i5u/zEZpZWzwXm8DE0MkRfbmBtbjIzyLhkGPhvAFYriUL9pXhLyXQOd8qYt
hUtJvaL2BWiOnUFfWkQJSOdVFDZF01JdQJOLgrBxFpGeGnxV9D3QG4GXb7h7QlKf
1Q00TgGvr3WtNvJ+a8cdfLzIF2OSFSEj5K9ipp5H48pzArXzsUj+70qPIcpn4gxp
euk05kaU4/bXKrHQ1zj7C4NObtljx4YIAVl9Pz/9pp9UTXJo1AEdNYz0tetcqNiF
54p9fPnXbcfsKZTn5P3y3YG5kKPrlKHFJPmvMOuWspxTOn+4fjkxKggIq2humthq
gGR9CynvPaSVQAd12B32Fr1eRT30h6tP7pOY/WgLIHhd3/t3mMr6Q9guvJ2yNJp1
F6MGD2RyMMX0YcbdnCvK7yfZFYqXF/SZ0JbuxUlRrWiBg+Gt4IuqAed8Lq1GdSJk
u7HapWQzQ58gzE0LQVaNFtPxWMsxk7yvWWL/Wzbs/8FT9+TAaJMKKrcow7HrgDov
03c7AVXpfy4S8pvP627jtAbV/ROlHt1QBDg89P1f3X6p8a9dK9GJMstVJQ8ZPdMv
vlQoZCtWFNggJgU0/tzlHFKchK0nfgKieHKM5RyX9Tsh1QqiZsVBTsq+VpTVACeq
gKJqvfxYRC7jdAV64Ru7E/T8E6pVRqXNlT3rmBHb/6rNiBulpmleWMmzv7o8cy1Y
oFfh/Y6TifJDXKjLi4qRg8G4V2q0sm6h8pD5ghrRZbQUJ64v07RexR9d6gAoCeX2
mz5E8dfbz52T3tg6kNTm5LoJ/g6sEpq55jTjL99IETLN11R7ZA92ai+tYiujtJxD
tT14kR77bCDQcxGBAxOF+ezRVIXjoJ0aMob4z9KDujn8LH3K6pbE0dBM9xa5RPdW
O+i1IWemuj4EvgaGezufW9e5yO//rR5uwDVP7SQW2H7Av5BAZADNTXw9H0zUuVoa
I7EI/IIJfyLeFvXSrIsrY5i+ZvszKoppus4nQCjkAl5WBxADeMheGfeq1LBD0E9o
ZF4N/wdciEEKoYv/FrblcrVa7jFRshWZuvjcQBcLgYqMH15EwOIaA2Fk4R7rNCQ1
FQA+sY+6qX3OF4PI5Pey4Mq0WEkmcwjedbotXqgK+a7/mDwTLeNzcIj7WLzgv4JK
XklASTqAjznY2rQ9cRLUBnGH47WLGx1XH62HHaLSMla6LaHlO3d7kI1x/HrpPd3O
J65DYxbZtKTFlpAQUoiTthVJM20Q1kPwP9WJx4syYHtK0Nj+J4Hwvi6+yJNPPXeq
zqEWuEnJu0PyhNK6W1c0YvqrdnYYG8DyN7CngKbStMHrA5nR8cjyWRVO+AHp9aIx
aw4hNs6ZEWQXYDSlySVzLSpR/U8Cj/3KhGJpBVidlvChLHUnOJbe/jEbgJoo2xVW
FhPHEPqj/91LsbD/+6gZO2IhSFlzkQ+odLz9JibVm75N2yEU1JNI81LVQ3F4wKB7
i2ItqwLIcRJN2qr97DwLxWWNQHTFLHInTQY8y5iFZ0fwBGwIzecb6tlg+7sgqp0B
Vhw8yxrTXLMZGjzCnGxKPz2zURSRwhQsIsH9DoW4tCibyHnqgA07ApFonLPnOYfS
TwF5baXZHoT5v6jeGurNEr56egggutN34HVvaxdgkq+otUjwoYhiCfxkuII0PLqM
Sln9yvr06cd+Aspknott2D+BEqmFwJKaC7tE44GSR9lOn4Qoqdl6mrOy9wtHDPQu
c339qmjDSGLF4CjdilmqXPNI/cifZ+WRIW6W7JnC4aW3itd/YIjSiVB8VoOCEZ7L
YUbFnWVCcpysL2CYXJd7TehaEYxMC9NNwiLXbNREJyKZaarw+KvwthHJpMnmhU5U
HwLzcP3RMK7fL7wWNzjn3PKbyAe7hRS4abJoycrzIViT484ByckP8s1LeYtpmVAi
TKKC+YhYvi47yBOfByMAhe+mncDenRaQLreJQODN1zyu8caBjJdHVle45BdxYpQC
X4DivRmJru/SL1QZDMK8z8UaAWMF9wU09v53GJZxxC+evVGbxB4BUn/etBN/SD72
NZZhcRywdtGoPQlCm9c7i3sibG9/HimUNh9bvFXQZGKh7+W1ixhGwZ1wanEEPmrh
zKw10oRPjrUMqr6KIXA0UMRR2JTfWOlCJdPmZcDSFelJTYkUbSjGVe0nDq/0tVJa
UbfGOWOz864jMEFHWrSCjQT30dl/zHUdCTtGhAMjC0W6JY//dc9SUeJ+9BSPE9LU
XSoIpP6fWTENydesm9uW9Qs54175QCTm9bclZuT61TuQH++famGwRjC6ZT+wZTtl
vpDOkE0Ur6NC+Z7JKvxZRozWRJH0KS4Cx5Hri6A3W/yGhe7ZB0fRpZ+WxD8LIdOy
VtNV2NHWod1XTnKGlkRmeUzjMJRnBRqFOxj62gesWv+1Dl+m0fo9y6McFfEORLmc
Fq6bHOlsQL3vARjcCDO68vaUBW5/Wwt+uZQPy2xd1iIbRTf297lSKPre32H6UTRB
VWIJqUtlMZLu94QvO3JB33tQG7sW3W94twD6h1Ea5f7rZZbSVKN2IxSIs/GbfENi
xsgxukncXuGeNf+LII7TYtMfSGipnD/SnCPo7wER+7obf715Txg0f+hvkgPt31/+
HaI41zpFho8v6rvgeIJr3jXZEUZTfY6b7tNPwpMgJG9vGB6YZd1aO558Enxgh44k
falJQOMdug+mzpqXG7rN7xOzmTumXdwfBcFZb2gv3FKPpG/SlqtWy8MObv9c7KBN
r8Z61Ng8te9WkkQMdkdRmmbPjTwB7j6xotOnK6ZnW9nsg9wjrUGFrTjevlzv9U2S
XOCLoRXsAP616AzD+59sh4uy7qBlzFiNyfzq+EdXNZMXtmX4oq6FOBVRyKA9r3Hk
+uNthMC2pGNg1B+tuknB0TrmeIIcU+QJY5K8fPv2IYdZuDuIzYcQbIT+MHF+Qpt7
vFEkwZzi/0faGBlAheXCavm97nN+Ktk1ic7148BPieyCV9op1O436oMx/HXpNIvP
kZYkPNb2z1S3I1warl5IpOG53qh4X+LicvI3LcB9cNTYeDNbbF0nKvXeSEb0HyVi
e0BZkqF9Zgk023dYSiOM8c2J7ub6nRZKHw/PNF67W+Rf9N1SspLVMfJn65xRfT8v
pmxnhZjTWzDMRCdUFU18LQE0WsLWFjB5QAQbmjFAcZ5xBlG8HWW5BMNSGIFlRCnu
g764WPAIF4+1n1brNZqLP4gjhxhCIS0HCHrpn/uyIlLoIPEKvARPuCx4iOYX4QYe
qO82WZuYaluWrlUPBNCeiz9YZru/wa/s0LjP7DwIH0NnI2eSxMbBvGftK9LZ06Pw
b4BZxAJRfr/GyaIE+aSeHhGtQEXwIWFbUZTYsjV26gh/1/hoohmBaRP7oPNxHJK6
xowkAt+xzX9QwBFPCpGG3g+A7EskF+Vi6VTmetHCTyE88i8KGfh24dCFVP4WZHCG
VA9twdsm+WZ3T7lYOCI20JoLVwKX/3VNCAII56Z0jpag5xsUm3QBlF81TlnXX/0O
yGoj57ovmYCNF2NiZMYB2SDyZqlegBdz2NjuGHBH72FWgi91tBEmnQmJmM5wd2wL
mCOpGHN+Equ2EWTujCs0DGcPYieLFMOqvW71kl9Kqn/wrZjHoxiyXjR9AWK5VDe3
8ngz5JQWTe+3Bv14Hwm8BnYAU7mxAk3eP1r+fTghba2TQerZ0HJM7YccQjwsnqpp
QLvygPPcG+gMJOqW9VlUbra6NOyrKnHgSWCIUWZCB3/+t1luQCiIQ+8g7RUZOmxN
eXpFwCygC6kDFDZlxqE8v0eaREsCzkeO2+ys5g69eCg61TwjwPV/t9YN5hdghYXh
eCOTglkN5oSS2j2UzSxs/Ia67Cd57I1RmUI2HhbZ74C/Ayuk1ToaYumE+lubq27Q
B4R7UcWZzhOZCDzjJGaCFFP+WwDUVhJ9Oxq6wxrijo2hCHII/iOy28+S6Iy6XJUb
uUQ13V+N421xPyQhmJgAKhDgvXGUpIwi0hMEZN4Bppakk9ymjXJf1YnNllQ+hC3d
2lwVQGyrcgc2e+8Y+UY1mNju6TDgMkzh6utWc/dzgyvzJNhjBdYP96uTe7W7tZ1i
d6svjL7MX2bx93Yk7oUpKBnzjBZlCBHm3FlTNMPMKSqwJritVqP9aK3vV7cjmCrd
ReiA9WQyEKPFpQ6F7AYpcQCi40wu4PJ9FDCCHqLJt9Lm55r1As5DdOTBS896R3Du
WplZ3JNAS8udBrWVNDeEWQTB/AAVFjlYOE31jeLTmI7VqYEqrEkwLULVb7zJE3bf
5geXsktjqy7h05qoCVE1zh33PplHOjRKb0TBPyTj3vWwZ0OZC40HX/00r39wxRn7
RzAIiiwI6RIBStUjaS9900hv3/djHtXHl+ED9Qkg02Ap/UiXl+/Kjkc0yiuu1JqW
8ZAsPBP5Ok1Vwfz6pLxv4Do5jWyrfe8JyD4Kq8dT3CiX79ZbMarlZi+eWSzxNY8T
E0uAW2S309RI10LVekOHh3d+wIpne0wQHmFVK8ek0d+2rT19rSk9x4d84GbCMkTg
1XLaLxWdKQr371CNZN7kz3ixmWjRcW+L07ejARFHYqfqyI7IEwQDFbKafTd+obvf
MzyUVPQ9V++ZubfqQ0aBlKJz3sWiN9MQIyai+XL2buASVHLlvOj2cM3MC2opKmVt
ucEs9EhtWRM4Ib4yS9ilIiMWl6u/BOMArECOKUklmS5KVfzCa+BSz8WtXeYHtKRu
f/RsdaqF9Z42udjXfNhTT9arwnP+NWejdG3eUgZNd/1uz11MaplcBpsI0xX99Xv5
iTKXPRe0QunJ1DO3/W46KPjRT3sq+ZwfiwMbMpmJLRs9/AxUVpt82UYiWbiGlvmj
GDHoowMCMYP3F7gcOpIgF0pMgEyv3um7u8nvBd05ay8l8Dxy/qMmw526Q34QyoXI
vcA7qY4vPiptyIvANkLH+nZhpiC4POKAHAk5w3UBCzBwRyfD7nfujR2bWZPBbrEI
Hprka67vP8loyTbUowRaf7UCoxwAH1PAgzup7vCPdqBE+dPzR2eAy0Ijky1++4I6
QqBHotrwqdndyAMhGjQPl9ZPZ+OOgcSYqBEX02Knn1s8cvIbd42mnqjw9zdm5Ma1
kTFnc7oagEgi/+6ydKnI1zjaJfpCEnmRXHfnAy6iiVwLFnLoBE+zo1rMSYplAJsQ
UJdjd8YFjuHUK8ERgaDXTZVEgWzGu9JS3OeKyrMBSFRwx/1KvNJrH37/euHdik0x
/U4JpF2Aim5jIUCTNHKFQ4CDEK0+MsgA2KLBuMatWYa1o8JxELOU3LhBt+aN0hpl
AHM807KAjk+ein1MbE3/ejv6OV0Y+HX3cWBUs1mtglA71AJfwAWa2Latm+H7V+xJ
08ZzgcjAg7AZqFc+Q0QAnbapR1G0Fm7pS5ohvxBiXBpjrhZc9ldKuZh5hZS5GZE0
9tYMxktZWx6GFP18pGltoOq5PUmTQpjpth/qIjr72wREpAOcuN2DkKPPFPVg6mtG
gqVjnEdTlsnKY7IGdFwI4/x01Ob2MCl+Jr3QQJL1Mp1ovvnKWPRXy4g0TPGGcI+2
Fs7pyC2JiiHYFyxv8sWgLWDevy6368/dskN4RUpE8Xh/D4clMpUWSx6AmpTGTJZl
otNvdzPYDqcORAN6j9R1ckWePfghLkDX3EmSzXjDAzmyTIOkiMl589DV5SQdT0LJ
KhvIpl0+lnTOmJIa8JyLktGjhV7ase0tWKZ+TXck6UUBVbebuZqEnDJhdb/BbR/N
3HXdVgjWdL8i6DmKM2rm/pyTmK0GmQIEvtK/+3C7EKxCW8ueeI+IG+svacOF82gv
jUUsH1f0BC5iiSemtIPnrfiuGNF0dLTFK4xlJeuWVQZHv4Eao0YHlr1IwwlMAoBp
rgLprbbwRvL10R62NxZ5ceCSNbPglbgBPoZN7x2iCDgLOPv/HW8RB7PKrZt6+hKs
VYnCck2EclJ4wt/vH4i+UYfA1QxLLJcYbN7IvsCBkN2E0qneQfzy9YZC/+R93N6s
04HlgWeP6PKuPkV9JmDPPK5087+Bv5G2FW8SNEI15Gax4NDnUoJh812XnxGCaQKj
WJsTQHMfcf2AXGOnNH6LppYm6bAfUCB14Puum2N81ueZiZY7yCiL4rNB0qypBzlb
pG9XBDJsrlPOESB+gUm98JNeatLo+xBlYiLHBM8Z8FC4E0rwxceH9Wc+ZYe5GYWm
kO0/xfeVkvCxZbZgH+hR/d6NnlLDfhuWF2WhTcjdpv1Chavy6jGqoAYppqxxlGsh
B/F2RDJVowD3c6UF40AddovWaQ+/6SM6ve/4BguvgDCPZl/3izuBG/XbTVvvjvWx
W88dF1TC9XnvkLDRUpomRuo+g1RZCD6R6d+bpHocn9rPmPjurLHbHZAJfppSONzd
lIPbU41PUwUhu+gLLsdZYHJqDG6iruZIU6EjZFnE3AnTvN1A9m0pUM3OsRCFUKd/
63pzLeVoTfSXCyKbY7WfMIK1Dvikpo1/+sVEf26/7GHqUAZZf7O3n9xdbRBPok74
qaZ4913NMLZ8pJxTD8ZyHpl6HpSpRqtjYCmHfH9YKXClSAay+nmqQ6TOGoep4qdi
0OoOhwgQYYb2rRKtXxdfB+XpPLqz4HUMynyHTO1hfyv5GEaL0OKnFJ/nyZ1GxkCo
NZ3rsrGfMacR9qoYjtSgAkKfP2qRUt+DM0WVtgPdkLctIQFgveExyIsFLjjFTTPq
5f4G/3Nf5AISjrFtp3C+ciri8eCK92AC2yHn1xsDd3rwTsKXE6d17vivOgoMEZbY
UG+v+SOs3tGI2GKtfJ0pS+pFU9rLB5ZLMOd9V2jyuYpbwS4nF8CjA+4iaN0b7sr6
5n151Ntb4xOXwe9DZt4rCI0RNHMhtuwQ8xppvnGPpgApr0E7IU3gHR2WVHPrDD6J
BQ6WknfbyaY6fUccLiAR9YeQQ3YUoDINLgzkXCeERBDFcsygxJdPeXZ3+WcPvrUQ
lq5+L0N+WBE4UQXkJIt9RqIAgNzYVHjQABHDUVfndK7oYMWRtxFzOvapG2YdtvRL
14A2TR/LLaQIw/8sLmFA5PkTGEMXMvgtTgZAEgJQSWFqDcwzqT294J2HV8XsytYM
KFNVCwnCRhdvXGdI36p5PTnI+flTmQtNrcPIU6gJlaFSJqMO/ANmythkUlJfdw9L
2TVfBmcyxMaVOmlcRbteLoRAABn0Cig6J4qmUCKJ2UUOdVpCvSU2tbnUMYHtDTyN
88tjE+mrL3vSbqmTorZYe9f0BIR4y9ZRtZ/Rmhd5ge6hu8Vy9eJmU6Rsa8JWYMzL
OAP7dDbw5TBbHXzsMCEiF/xQ0KPkoVva4HMhyqdYcavGapdzMJSJ5Y15W9P+uUU6
bC/TsmHcPKbZnIXP3ZOMWlkO8CPrJamHUdQ+DiMcfkEAxWac2NnfPnRiLApDcuaj
47g/VgL90NipkPL66jekniYZm2Ehr1tvGSuuUZCpCLaipiXUEbas6XdSnO3pbSNf
cTyhPfMW0Z+9dhltUPOKum7iFlE3P4Pz9w64kQIqhAVus85BwwLdIN+zsnEFU5MB
mGgjfXm7+uZgXml+p/cqIPTtjgrEEd44T2J+DtUmEsosPoOuE7ajpwnwhAig1b2S
SvJHUYNqrDq0qsC+xkLwErptRuBrgHxBhuszZ1Fi3TA6THTZ5YXoANqinj1riwlX
1eko/3wCZJ0R/ty12wN+EudMpzKYDsEhzf741uuKarsLRBfXHSAl6IAZ/Hh7blW6
3yNs4B3N3WP+oPisqTmHmBUk/iFD5+F7ISkApGPA+roDqToS3Tp2yxjSWJ45pD9T
b5Uh/TTTImhu/l0FT/NZ8ZhiUSCM7itg3AKlY3wzt2sjcOdauBIfbfCUUkqYnmcr
oSQWUOnX0OOhVIQMquY/cy74chQTC95Vzq4MwFu29W76wDMjwmv0aPsKvbP/sllD
3gjXyehyPFyghUnmyr9uPDk5aCIqQSdIXXyswHYpztwBgchKrUl2G+LwzSQ2isuI
6XYRBO7aYcjAyy7JwX8Dih7izjOiBTiQXBCsEJswsd3L9ZZjCJGr7/3Y09rZnqzf
WXMZUdXio6d8xXISqnFksmKnp81b2UWpqY9qYrKpv45ohQL7HQ/n0jNrBAxBwr7f
oIzf+CF73ZktfpKjBfLrIHkNGbYkBGxWciiT7OvF+AfbNUuR24ddZr1KvC1A7NAb
tyiQp9GbcNBgfoxUtLxt9uEUE2+InIXOJ34NLI9c16YXbkr5OkpFclXX5TyvryHH
plYWkDfno1yeeUDs/FYTqexGYhpKg44A+jhb8m2WRHLpydW4MYfDixlgCM6VGm7M
pv7HMdS2k6VeoTlf6jLQr5Y3SxAEqP9rjnMSHr1RbODwkrhJ8ve4uWrYASWdUEGn
PpiAR0MXI3oDcHVTyIHDux2U74biwloj43pl6xppqDdE7XEwch07tJkAi7ZB9zA5
81X1dtKFmk+wmaNBPAdPJdyYa6OnAOZMXds/ycb0MpHk+Q+4KyrENCri9xVta+mr
z1xWqMYCR0bJABE1kYBDKHsHm6oDx+eBvqWf8JxFETimQay16wRAKHLQ/nP+DdZX
k3JMB/K+65Aai5H3UJ9z7kr1xN7EAhpyoxi2sD54S7FD4oGD/Ecpegj1KVBcaxt2
+9qbjnKrBGfFiPQbRa/y9mUowvunjDYjiBnXM6bMQX53NeoDzh6OcKQDP9UnZDJE
gZuHNz58qd4ptbZjIQChr/fYgSoUk+MSXAgfhIi/B4hgxPVp/C29p8ZHGT+WWUPH
hmqKcO4j0uekz0eXTTCuxvHkmcxsDW6xu/rSBI0awzlT2dW/goqtCC729nX+YNr7
97m1quyB/7pkg3bnqqEtjRhLGXGBJvEpHz2FoYw3bLxIpNdYCma8Ypws4GDGtzG+
dpTQ2DB3b2FSJk7A8r31PAiHEIEmLog3/YoiG874U/Rj0S8tLspxmr+5U+dKMuCj
3RLg7gALoItj6rG3uAqG81kC04/H9Ovh/R6VFlwp/eIeCTusnHwjOXtJzEoHN4kI
nm56rYTIpokWrXtbFyGqznXrwnfzclq2nCNXuN+bKtFcB0fJtNrV5fxPXD7vwa+w
u8/x5+60iTQtEwkXOfoWRoYIBNdXAYTA/QWBeKytplrNt9CPJTaMzF1/qyrlvSxR
IbUZESIIgfeMXbKYyb3+gwHf7EU9FsBFu4aBmaNRDQC5ypojcKAy50Q3oODukfg3
EaEPLb2bXflyTX6vjmFZyJLbLItL/GiwaijA/KehUUTYfLhvMpSkFcuNJeAjsVnV
AgDUsNscSClW6vIMXBFtPNP26kgCF1BLj25GEvjMrvWUvPgZrS4JPxaHRcpft8tv
1po2cy3O1bqcJQ69qH3xf4Mwld8rvsvD+M31p1aeJ1bzsDi6x4pmZL+rcg6WzPVb
y0WKec5fIq3VBgDefd1GbI9yXAcwJDVEWru0eR1JCMFVfX0Hl7m0SjpxhuDLP1K/
OPGzToEblGJ+fWDKB9fCoaQJkgTwGaSLJ6XVdJCGF6iVqdL1QvnB2FBVNGIeb4rk
eG6GRLwfXrOmvdgrsHPIrrTpvyZqUZF/v6eIxHapne6GZ0C452j08y9ulmBHJWA2
ijMaaaHGOeamgdrE87fuZComd5sK5oUpHjixVYAuazfYXTeSmWH4YTikqwHLTPZN
yQIMoFfbAHPogQWAhwRqLUOD9WnfRlmzE2t4LYCXb7Qv7WePUYRnZ4ueRveIeWzJ
riCPU2P0u15AX4KmXQkzSGKJ0iaDKy2ZWY0kUInSyndqnHpN7tgcL7BP+s849eu0
aHqC7QMXuYJ69r4iVTB2vythGRosi8C2pzbslfpje+U6kH/0sEdGWmjLj30y7fOi
MrBUhTQG4yXGpTxQVdkciR/Sk3CFcI0BspEtacXHfI3eTTcNb2zPr14ewnloOG7s
PG1fli3VaLZYUNkTzfvZCuOH8NtMRu6hJtRik/BepFF9WiwAAdSnvM3SDisurl/8
1/vNsHgdTRTv6CSW3/SptpC9iC/BaQzdyBCAl9Sub4VxsNSJscVsYJERZkPKzVi4
mTSxzm3NugBh48sr7lJK0PFb2DX0Tjh8epvMu8h9gfJQUV/qxrET3O9e3NlPyGVY
TQTpZL1oHHMKHs6Z2iyItcqcHTiaOwUHzbhQs2YzLTGqqndXfN1lGEUyuuFK69QY
DYgXHB/dC0XrTC6Z12HhbVXPy06NGsYJ/Wex64RDoSYUhTCEGSFnp2eKg5CJ+xjD
TveZD5HCXAOviYd49zaeFFt4+rg8anHTLhQ7618Y8T6+GRQ281NwzlFf87zoXFfK
lZv4tVTnBXv1g9LHjaUsSXjwTEwDw9z490iPrVZTkh+W9oDRbGZxbyFwwkMJjRBj
jWmdhIs3a/jAkwev3BF86nnP3O6RkyiI3yU1OhQbLly7gN9fUbgF3TZTOY5Rz6ob
vMiJI8O1uxdiQWsR6VM1t67kf7h3moQaUu7zScNGJ3x1PxucVjNGTjyuVb2fo81v
9N7U45VhGWnQlJE6c9OQOPRLsbojApVHqhckKXTg3c0WPns41vR8KbbJzFvFRAAI
QEjzcLR8p0F2B+g6UwLPar3E8fI4AE2L/+de3faiIpFOFJwfbWQvVhBXzJiOKPuz
8LwDOOEqiYpwpyw601rgXOFnc/dpWg6ZDgOMZO59yOo6Atc+DZVvzWVrO0LEaWvi
7JyWKQ5wir0iiojfJu5pmXPhAvg77QQPU1+q7lOEbZvwGahKhJpF/hzxjSQ0gBCV
C0deUdS/X8J6Sazfj14L0MD/ashbplMsUixo9ll9MnuDmFaaPuKHYHoMf7+tyXfl
TOSUySJQCoWZS73I7cmRNRMaNtRqjLmO0PfdmsTVN2RVirITrk6UOsidRxA7CNjk
i9leCyBUKzWrl3rwwVNDTSCHi7BTOlWRQCanQN3v840=
`protect END_PROTECTED
