`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmOvjpdfU6FTM+0MQetBiYhQsxHTFpmTjZTEDDXaGzvJA3Fe39yYH8mOTLSpihsw
PlekMJwu+vUexeRmt5yiuQRRFk1nTifCXC0ARQLmMGki5AV+IxHnKwHya24gbvUj
JmQOdeWQtE62VjjD84YuSU992vLNmpIG0J7nhuplM+2knCrA6tgtHpBog0qO8u+j
5tqMPyqmghz5CBsN3Xrd9Z3AAUpclQRN3bLp/UIgQoeLmltsi31GnD80tpAyvLEm
OjaGXnoiajRnZtDYvPTpPlQVm8Md4k+HXtokwpN/RkNnLkzGv+SwwsC69LYQLxLs
A2SHEh6o14nGBfBE54Il3yhXqiQdvX34ShrAIaRQ9xCWmG3g4z11LR/kDhydXcCx
sd7dvr/F7Qvk4Ri7uO8n2Mz3nUbluDxCV/B2kY9ruJzrWuM1GAZhOj043vliPfIo
LlTSB7nvgdkmgFEw31iD4jG+N2FdDZTApQofLXKoH3VyK2I7Dh6B5sLfo9R4oc5A
EeG/9CvLe0Z4NM+khwXYhwh/Yfo1WpP0waTJ9U0lUidg7QeFnFEzdf72bpBo6NFZ
PNUFbS7GEfnInWUX8QaClAm8qkWiP8M+YkBJyRenBhyEO7HDdWNR5mtXqEgXRG3k
kVoq1eHMJzPKPWDcXj0XwJUZKGsz5TCQTB5nTxcGNsvhYV3xYDK+t+benHr1uGyF
Ql1sVONfYZavW7foc5mZwJWQmDjPQVFKOLPZAz+NGrdy+yC+2CZNtcYHXpWee1cL
B604Qwl+iCbiAHL5QZqLwBI8H/b030LpG+0PDc3+9Hwi5m4YF1Z1DKQZLOjrQyHO
gDkeDAI5Fk6QORqLUkEkpGqpgqRbhZZmo/KHUZ5kiEdw/BqCEb6ECaJuyP+qaarj
E0ILD/lnqYHLPL4Fh1IN2NpNXzLCSE3eij1gIVEaneyHRb0mN7qI9uEMOB0n+MNd
EKmCCzemrfMUfBE4jueZxGmmar7svnbol3R5HOdUrVYC0yIETs28IBgcU8wBPECL
97qZwFU8mZlbnrhwkv+v0AiZx0cgWqJFYX3ELaEx5LDBKQgM2IomY/0lSUTv+Z/Y
gGbnwth55cwwAVVomr8rIhU80auqPsZZatfeM6ZAMSBVVe/QnkFR0AKiHWjjMqi/
CCBTtbghoe98ZLLJq8f0tEv75kn9SrlxP5ESBSyNQwKDV+ZbNiKFdV+QFGKuD+9F
WzKEVjBl/7OWkMzjMFMzoALsmQSUfi/Xdg+vFaV8M3OWpeYjB+q9VS4MlWBJPrIH
QCZ0IjTYRGAx8WESGtcYcwhmXIvZPrFvn1df23CqQQzz/1nzczY1dI4T/rTI92sv
lF9u50dX/oEF1YmKjl+44X4GAKRUasouSQjHPnx3c3OkLIkX4u8/IhUnUxhEjj2/
etTz0j2hQgnFmAITmKMRLQ==
`protect END_PROTECTED
