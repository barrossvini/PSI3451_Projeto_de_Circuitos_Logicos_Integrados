`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FcMC8DB2Ij5VRzBvDogWDtBQag8dwmgJC9QWv7YAoEy6rDvB0mldE+gySpE5K65L
BrYeZ6ZxP0/9UvS45ns7QaXI1qJFiJvde8AeF3NeoIrF0hs6j2UCS6oS/12U5Gjf
unY5ytHTX3ZoIFkrK+PTZCoIFFu8aYbq6vht7eWcGX6hzaqDUvccevOavxgEy9yf
TW1k3uk+TaA/PP0hXuu1dSHm3IEIVODQP3uALbHw5+zgIiSt9PgSqasI8906fJPQ
J9jVqw/hXjf5jG3DNVSceTrytYFA7AhqJBWq21wy3z6eyKwLrVKMloPDE5DGHIIM
Gj6bitawMgOvbWHlMCSelJeQ8FZHlDQtK7LsFLtMBlM9qCfHHrtuoWbryJD+3AAX
8xa+2G5XQ5GBSnYzy0dL1xqzy/IT+4iZwDgblPwjIyiQsIJHrh5y8HI8mmmB1myZ
8rjSYSJGa08yWVgVLSmulFoG7ZCr8imZQ+tH9JsrpmlTp7KF1jOzOrhYP0B/jfca
m0Xdh1BI0pYXgn4/AW5PD5Cysb+EHFOtbsMzY8wHy1vTP4HjAPQ/kl+ObYFbIBXD
tIRAVAzde3NgVppUo7N5egDO+yPxuTw7qATumjFzwPyv4NjGU74rEsMAU67lb5h+
MZW6LCMpZnW84FGGIwY0h8ibxqQG6BIoHDdv4dIzfcN8ZKbihX8rvmeSVhJSsimf
2O+DLiqc901STAgJQcZUN4FDBbjN4FzCvy9y2OQFfy6WAN3w3dJBthDqgLxob8PN
ZjEdnGtzMCl0/XQo7CszyqCmkHPZf2RRtrLERYGNS9KtEfA7xn7oMUYIbdmMwFaE
`protect END_PROTECTED
