`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cQdROoEzQBXXwnT7Me/Xd+gjNLJpI+DvI+U1PxHhNOYSuvoFkAjHgbwGSv8Qi/sJ
hPUBwIOAlOv1LbHrdZmhxo68co9ImujxIgek/MVXeFGPatyUfUOTwgRJZdfkA2Vb
7CGeqQm2vkECJ586+quTJFGOYPdiijCUt8jOMArPghJkbnnE2qLJWyoKOche9jCX
aceb5mxJqUCXqOf4BT6QUYnDADPxEDr3FDpfLshfRLnQyoCJfD9J84r5g1Lr7UqQ
HQHOqdX5AsIXpQ6YHB8sBGS4GIthq7uWKic7/nSe8bEL6ofda2EvPow226cHCr8A
CHVXDB0ewKSbrrtF8SYKNwnOiiiR/CavHpXdnCI8N0XqFONm9z/G+oddgfsK+6bI
T8LYP8feKfkxT7+ryMALJqFYu7SUSCPjYs56ULr74HI6Nj/BxPvF0bKepZEbaDcK
6Uztkv+0NufYzzC4zmHlkZ5Fnc7jZvJmqoSqjRvRQrWR1ofLA/MP9pgFq7X9T/cx
B9JHPcpEQPRtTTNVfvUR3+6xVmJCLt9I3YfC2NYT7ObA43Twmwky4LMk/9ChLP0T
jUpBps9Je2+ARocNMRMXymDp0VOF+qmd9gM4bLvjCHwKlb6RUsq9DWscGluTcVvb
u/5YXH0UKjTueYmCxbG/gthWcKltj6HbYTi9Zuf4xvW1N7U3/NCC35IuWjGcqC9m
+b+qyaUX/E6mSH0kfVNkKRSvadfVzF6dtjc6ci2uZvc=
`protect END_PROTECTED
