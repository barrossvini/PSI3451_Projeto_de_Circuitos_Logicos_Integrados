`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I07mdjz+EXDc528pDhPhx54q6vClfv0nfa6mmtsTXA4zQlDR0jmBKRTLKYQ3z8GM
/J9D7KCrlbkEZnUTzS1/U9/rAaJeWqSwqscbxrW+7U5WsrScSPIxJpqqA7+1hf3/
oaH6595i+Knwutnf7crXCWdp909LJyE0BoLh5YToKAE7sGazhttfwJWWAd9xIHZE
iNqi76Li3+4dkijOTYHrJnTFybVglBxn31FjJIdEWrFygsRoOdDlYynACLk66iCk
idt8cKodyJ72QCqZrbocwYb4VTNQbviNDp+Dr+wm7QL+2+1q5cekNiB2gwAG83+b
xDOozF7lGF6uoGcdOp7lZ+WZBCx4F1ZMF2kE7n9eh2YClFJU9zSPcd6ECAr1plo4
v9ST930ciKZGfQRobBXAvgk/7kQ/5CabwCXkVmIOuoaseVxGm5kr8+6sViWuYLkS
vFGmmUqEHS78B/bDt3cdseFkkb5ufwM7+K/GAOC2Ih3hBoEdIOy88ogJ883ez17z
fjlsgdygmw9EFS9stDNXlAN307Ik0/DLGOjHUNoMCqAHx9nCNY7vUCMST0AxqPRi
vzCIuottVcGmiS1aiCr6aj2EW2UKxiw650TNGS3fFhNcIkQkwlGS5aWVMZEQt3u2
`protect END_PROTECTED
