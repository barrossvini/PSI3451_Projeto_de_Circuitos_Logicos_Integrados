`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
faY+G1YvOA7TJ5KCVndDkZoN1+ehGWXFw0Vebnry44cYG5Q2cV3lOpGuJtyGsyFz
Nv2Lq2TMpUc83i1GOORsPS1zNFiIgZmS6nyU6soySpFgrmlPS+5Pxpt0gdYERqaN
Z9dVz3RLUbPcFDroroFCeDf06TVnEz5oY6YlFtyGK4gA8YsLQ8lmyH7eyA8k7niQ
YOjtOPorXWm7/9opeUG8UNOK/kAm2WdSppOeo67lrMr7JNOyutsquTvoCs2NAqN7
TpdssF0D3y9DdNKySHiGvnY/gQ3uRE5jWw74ldh08JdXhWn2x3aDRxm/f0wj6JKA
uLI2HD69JHQJM8XtBNjEhH9yUaChB4lKQJpTYGFcCNL5dZElvmRaXtw5TWnI+bqv
9hAOdnOgI6HgIWOfg2+5Uz1Oz4oaBxGOgCSwZBOSnCYX4pO2XH2L8MR90DClMbLW
v98c0h65GjBVU8ynueevm4fV7hn6wl9bvoi+/oCRdOjbkGB2KndtNPOylkqkLoBb
pXo+0LCPJD9BL0GOv71t3PedPMBe8xbKcHqH3umBZahjenZMy6a6y1RyWl8gsw51
ubGt6DUqQN0A7VsDc5qar3FL3BowPj8435dljro5QulgW8qenJPlrLWiAQPVYm4v
E1M9IGPoS93lx1JpH+jbjCcW055ORBiYovr2qRJn99i2JJlQ2ZjjYUnneJHMW/0K
6SPCmg2AplQrw/qbqsV+e4m6ApX/0AxRK1WPzmpX2Jo5tF3AwjQ3GMmQEiAmcCJD
FzpsFLK6O6eB/cmVSsVHBsqDVY9LWmmK7bSm2z+CCjTlk51w8NqYokzBukpuFnuo
1R3j2bSaNOATAvgVCflKtQAFK56JU/lAva1p1eR76oO42VkvYNOe3EXAdgMLf3yg
18om4N1R3/EgezsriwJtrIec6bys6boc1/l4w3N8V/38I8abeNHcfuZQDKQCI1Qd
xuvK7kWo5RRQ0/eoUpi/tmJD+8A4i9X8F8M5Rj/QLcuSmwE6h0ZF06r0RibCt14B
XZy/AV/tRfta2H6w4wzdl+xCPAVGLWo8tN+ufDGfdJm4bN9+sLHhaZCZNEbvnbFd
7pavy6Hb/mJD0vkBf9827IdFVgtQb7y0IaLtTaZeEFJOrFMyJsaq9cphq6NA6O/l
Fo78qUpsJ1JoyiAHk6ybcs2QrUOf7ZPSf02TPMiR2iLvBG0Hnp4hCtqFWQEu25cm
XjEKdUqxxnHodW0vmtwdXhgXMRsG+2KdEjkjIndQ0MPcu6pe8NTUeUumA8pf8z5z
iqqiCXLIE3ApNMECmra6MYK+y8JstpmcSxIID0K6hl+MGPkO3CTJtEJsE4xjl+MZ
W4YVGqkfe5w45SL1diN8rZmrng1CKqzX2PqecvKDTwL03sKb92Mj7HSejQsxnEg4
pUHNj5hdoMSfgWG/fIcgyczZAASWeximqAR1DPDbcqemEDjD1JYX/YzS8I4TMNSA
Jd5W4IjZMo9mAXa/sFYXtEoZt9m+eu9KaO7XaWXWSPAmXz8e50uHCn3Yyg/XuKBx
GmvZLKmAYippHDuIR0AfXysrsWukelRrtdsCVYn8dCaVxaB3i1gylF3TGWVq0PKs
CDAVMFW1YG1A7dJfszBNalR2T+dlDH1aln7HzssLlRY4j1PKzrqyZ/hAyZLUIpBb
xNePpioqpR1pk1YbQgEZwyilttFd0ewKeJhIv9oGla2A9cVx53DyS8uCw67pT9h4
QYnaOtabYyiIaKE8fmj/4lk7r+m5lznD6BmNUuDMWwF01SDZLs9+SOxeVmp23+hT
cgGEjvxJpke+1V0WKQDoray9hdozs3YxwApJ7sDoiRa4OPAq6AKiE9JT4fbj64BT
aSrcE/rJnVcysxt6M8YKgcpbN4z7+RlHZKt0xpB5ikAwV4sufjT24HtTL6jZJh6h
QfaL3iDjrp89PTNJp/zcBonLpgaohi1sUipZVJDznbXTwv/u1JohcHuYzyo8c6n3
mW4r23W/te5Uk5AIDug0buDqf6H00euO/SqC0EJeK900IAigeANJjcInpPH0K2L0
96LafEMLki0rh089cInJnpuLGrSwVHcctv4UrC2icGPS6puwbH8jSpnwjNbz9dGh
+y7hQlMvnZaK25DE+B+5PG9GVUZrkVCa0yUQTuyDWXC1nkYy/CpfFsu3hWp53cAZ
OSYlvFOVQDayBfRd1OiXxK7s7m2eUFRsTd8La946vh/foS7aydpdYXEpMFoirdHE
EHuBGzpaiJxqLlMRsWinC7QmngsVhDehQkxva1jFbUIgnaVI96Z7xvFkSkeRpWQb
a+1j47UcL4zHoTG2gr7Uu+kuR2RPs7RjoJFidEtGmobypqktR+d7CACQUoBQJdHc
PG7jZ309B5L0I+iEpbnfJ1ECgkXE4wz2h0GU3f5UK5JY0JPe88a2t+keXx4BPpw1
xCRbpn99LkIsre1CWcomdw==
`protect END_PROTECTED
