`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vV/Iwr9XG+Zol2U6nBs+qeMamDw8TaOKaw6nepsh8fpZN4FqzCtL3jwemllP2lA/
QzUah22gMh9WrsHtkbQ1Q9Efa7CPzkVcUiOpUfuywlJ4r+rN1WZca9Mc/wO1kjZA
fhSIzoMBqp8/p7rVYlsGVyrRnVNK9LXkkw/V4HIbS/SPlzSHG8oiVoBM3dBdT5Af
GGkMw8muyN26ZPdR1lmzRAv0LlZqiqWxHzBaaYkxIL6D8lbwPp90lBfH2mQtwnqm
uHz+Kkg4RaLMFQ2Ewfa2pn6ZDqNQTaA/UVVR9FRixU99GoYxtXiXE6b/HJBAlcFg
7WLlv8db9E7575qX/NdDgFi+bSvopLOXiu+nPUOycJaj9GD8H1acQtxfpNiIfKW/
FX3NY0pRC5Yq8Vzd4FkvSTpacfgDo5PF48rgESZ46QS66r6Ijp9JXphMwl0fpFOQ
MIa7RW1R5hSjJHrJxoadR7oEIm28OmVft7MRE3m7hKxelbffpdflPT8JkNhbwrt/
rdyM0qB5rf4gKYW7rDTjeJYr8Hb9vGXHRFMCN/6xSxULxKxLdIxfwWcRq3nfPd9B
TeOB9gPKVV7O197GIridk24mtuXQ3VYSrMtSN83Rj+glujh6/hA5Aap/ounTGs/p
TkVNvrACpPoNg3ALxcHE6bl3pdIEb+EEHOjyPS5BMEFfoD85+KtRufXGOFL8aJSe
8NNMOiqV3/7PDLbVKvvIcTGAtIJr9ZhPdkD0nh4VP9+r3awyGWc3ttAtFgsPUXU+
1W3pw5CQsuQB2z+qoQwR5xudVhBNj/uFAJItTilvAIuK3dp115uwcIkqB/hA/raD
hXTfn6m15sQrfK4rNCbA9/E3+9NTpQwg3axEU8h1FCCQtwnGz7NJTw5wdJguftyh
8eIX3UnttNVrvWZvEEBhU1hIwwH1GwGp4xov40AYbjrIblAn5LY7p1Z7gX2+UD4F
B5Yk3GO+I8Cf6hZt0dp9aEXYYj1w+B4CaLz4oaFkLEoO6/M/GHYn9NOn88ojMpX8
joslxT6tgxhFq4kAewTY874h2K/KyCJpyD8ASiwHanpt5tbd6F3gMT751feWy7KK
LoZiaEPvBXAwKUPDoUadfF9dL+Zc6JRGjf8SpqReHHOYoTxQlKp41yeeGGP5uSG+
PVgNfLFuuxHC+rFvy7eSMWSfLc6m8kuxrO4TYtP2UBBKVxPuiKrmL+oMOUbrw/QZ
vIvmY9gnvZiQ1PXHDttG6c96yBuNSogTt3LsTZwZhYXjNYMasAnmGyI30+noVDoV
fSiYQCf4x+ikjRgRVLSGZmDpsGC2a0jKvkK1hvLmkder7MA174fQAd8lixdgnbGt
ft9YdkX50n0VZbom1D82c6OUt29UH4DziZzo7bZLQZ2xxe+bU3fJmfBBQSIFL/9Y
vZ+cmGrYrkwR093AHgUudg8+kykRBPvvL1pWHuY+QptvnpxW6JiXhT4v8Xv4Q4i4
N9xIwcq6mohcqrubcyy3hsVavuAvS52To4cicgy1n/bayVoLW0rbwprOs01umPWc
guDogZdgOdyZnjNJurU/FteET95ZHdkK0xaBf8IB7iDA3xFHi3nIIpgU5mSBVpnQ
5FAGuCE06xRazedTC+q9YMOUN06dwHiA4yoHndZA7r6EG7NviJxR7LsBdHTB2p5G
ViOgFhG1NvlrC/nA9Alb0hisVVcwFHfGIqYstwiduqxEVGWBK78TNH8isP4y0ykt
3oJQHVJuclkgU6QJXgSzLH/MwaGdW7nzki9oaJiygCPPvX4TTopb6JsRgAb7UwBY
neQRKN7IO5XLd3BvR4HLPjEGCZEWfeRVsKuIPs4rs1mmfMzWO8+3jtfxOLdQcnAh
grd/RSkJkITU65343uMMeLb8Y+UNJeyolBPGjllh55epU6P9HBiPkUutzj3nREA6
wtXoYiD14uUCxG4thYxoUKEgSNN98V2txF1uyKHayh0wHtlcfL61duA+r8tTDO21
Ac67Jn76rHjTg6D/puU4IDFkEpXNopXOGKPdI52N4DgN21ccOZH5ymnhLbwF/yRs
2lKa21aNdDYP+FsEqS7ZzwwuSXyycuPnzzFMF3aLo9ZrZwtAJZXASsk5G+dHtced
sg1h+RA6f7RKvwj5rTHDsDZ3odiWAFdq9cNb/jzxrRehCsg2nRtuIQxdLdYp0Lv1
3SJ2/jb1HHIDcWnlia1fmF1ZTij11z74GhX9LHciKydRvZpJ0HACTya403YOTXmm
iDMAflikJvSea3QaQQNG7ZsCf78bj2mOZCJR7Aw+4FNoHLcI6cenhWhoEab9vN80
EiIN8B5+xIeQDhr9Y7fdWbZGpyAfKcnCe0HI4waNXAEr62PqtvWA56ue50zns44M
yJ0bsLPc3JT/oyLGL5+xWt/4+9k6UN0jMUBrjOZ/DKAsbvckcFP2TDRpAnAPNrh0
s3MC/3wI4J6IItZMjqSE0NkWiQ0KDxge2LPwId6pO3XluU01+j/9dEcamRtWBJlZ
/s1OIfPFMgOUT1nZ/IIgJ6BHB6+hgjZQw2jcwIKLhI9KNvF63L4Hy20mBqRMQdJM
k8cN6jcKgP2AE74x+skh2cUXNYfl8G92LmqGgRyf1ek7iB6OxMwnpy5AM93dP/Ba
bwE9Hp9u6s3pXj/0wiZ4Aw50Z/J3j97NP2448tpSZUTKEBV5v+qiX6X31+Kx3umc
uRW8oI2EAeYfCqBGJTfYTcX3UadqtFEFozo6Oqe0A4pJ/oV1gMC8/Au6UepTtDMH
+8OutDlOB+EVPPD7LrSTueNXhjqyGduXDgZPUqJTzmUgtmlZFYo2AVAJY5ykjC6i
VEj5gEGe+sQsWc9ZxSDs/elDL8rK3M0v9hTTzAjnBusUD7OFqqC14eYQUmhBOJnp
STddemNclJMWKF/BFmvXrQZYpj7ym4h+UZF365DEVHw4KNWpw227IfduR/IQmOdf
ufVJ1C10iMJ+blvO8+Xc80xOjGyFNljyq5yTupA8m+PmwJ/xCdf03Ij+fiAHgTm8
wLrnkg0noG7nNqlQh1lYx6EeaAFmJuHbvbzqe42xNxM0sYh6NE73t6rGYLvxui6d
1bDnWtwR88iaCu8blu0TKr7WQiZ+7HL4YnZpCEZ/lIz6ukO4wfwU0C4JscKCXA+F
ONAff4CMdQs94yn5YhaQK8AYXyYG3XUfWd90KqGFvF5foyxTyPHXgLf04FUbItYO
1wlhGcedP0I5zD1bO6/nz/afVIChN8dz6xXozd0WrzhHArHYpBNYEZaRT++lLKkc
oka61/pXPmqV6nZqDOQaXYCcBvjsi6af61YKaslTgiSxvTB/aVmFAfcIsujmiq4n
tfxRrvgc+mO4Ji15HYCt06ubP6iyTXNlr4on5A4wJy0FqTJqCnO119//wSToJ9f0
4lsu9KJUjqeGQoKxe5fQ5PVZoqQl194ZH6A/et2LVtsixBTP2wZW0ujL8TWKz7yI
J5dsXxtgR1XL0YDyFTlbv99F6MpfLl+iz0kBOQg4bgTCvAXgeK+eT3M1zHTRr6xB
kFeiqRIMHINmIsmoIiuH5rtq35H1u2+DEUxdyl7pRJiRr5HQ22tCQXt8c2/BWMrO
ez9sGFn8nOjARAZZ3FhDjzSuQ9l1T82vO6qnmktI0zR0OTOV9ROKWqdfffvrphmz
sLWt9pgpNUyezfuH36e0fihJsKb1l0sHkqar6rrDdCfzkdax+epkLvvuGnwP3AoC
Q9yqSzb/Mdbjx0UYEy5SSCYfXmtmnr7MqSOTJGzvF2EPLj66XdQNsxsaNiAjXda5
GHJzna51ejlHSyCej5mNsBZeRyMOj7l13aOPGKcH4Ur7HsSCE1kAAO3Y+WP2yzkF
D6dZDON1BXrALMForTjh2oojv7E7X8Rpa+ZRnvYCATOTOFUbPAMghFCMdZ6jMcvg
BLJg6N91NDF4bj85sJbGF+AfskrmCWPPiWywWSkHKvgLRgTjzifqSKd9O7hbIPAZ
88r0vkKICJbQNhnWiNZIjUugnknCdj5cmUwGweINskQgIhb7EpkXlsCXqIJksPrg
/d++UsnFQ7VYHnfkpoaB+Z4cdBrRVg3Go9pxf/1MSO9WVdC9fdfpE06X2JlDqPH4
PkNaEfp0T9qrVF7qCg7Cdw0IHtoJsgHbS8wgoViTWINvn0XnZZgJgD7inOA41BXu
y4RU9UaUPdhFEGHMT4nkQlt7B45tbRmWfbPfg1iUmJbN99K7G+L88hDGWropu/12
l67d9QvdAf0DiiDEodt/zlhdJ4gQbQMFMfvqaZX3vgSIO3HVgMW+dfSYR3ZTusfS
9YAQlglHetZEYMaZR1Is/eDAyPCDfJn2MjyWoszYpmz+m2AN7eH5R/AXFN/AcQSU
KVtGSDeyGacxrt/7d1yJnbIWcfXP88zdpII/Kj01OsuNRiDa+fomtpcy3FcPEg5E
wfKnrLQDq4myLG+4U8nHT/SercXNKZTWgNCpmyFbMm00MiolxU8bAA7lg1ZS6Qoh
mKiezGLGuFVyXb+5UaprpY2WLndxWM74L62/Gg13D/PBthZqPGMlLcNnDbmSLFJE
d+vq3Zm9HqmWKMCRoSc+FRj6bpbkUcleBSf7Md7KSx/f+gaQjNsJGHY3yNKfNrKg
sH6TIlQpq7/nJ5BVugOJA6OigXIhm50OlX5qmZA6N8UBoO7pauT0z/1O7YxEmQ0z
mLmgUO7xIlBtObqbfCyLEOAFa9AGhFeCiN23XiUHgg1dPr6j7b/6IlkTWqj6bOrm
qbtqFk7OkYWVU+5O0mwLknPOl/3JNx5AiOtrD5Tax7OcfBNxAXbSy/uZTBvRCm3p
a9zL4STV8eO5zV+GmCa/QWZk8lhyRqhU5G3Vtwkvg5Mp+qdaEepjGy4j6aL2fRWg
/jfBS/mhUqWL2bvoxciFg/xNgF2gwPUXULVDMNBuoweOXs4gPv5KZijB55XMPqF4
aEMckvRqiwQ6cojU+yRrns0g9yNNESZSafkAanK1MGVZ7I+wcKpTFPBL2uAAg2Fm
+6tIXDEG1pTcJDnJ4reyyn0siQn4WTY1+uUh3ycq7InUNDkH3xEmiFiJAiGKeqyk
QpAmyVRV7VyAT/XOQoM7P2I+n8UYBO3mnNpZ+VmcKDLj0eFX50o7w1dcC3GLzK5M
kiYieM91so/Iwr1JX3ec9zoIZyoo+nBT5+VY2/koCVPh0WQh3T5NM9ZhR5Im2uaX
u0AGqf6nROWemB0+NG8hVgafPJFT9Zh7YXoLPrYJI/xPVaSdf0/gyX6WZL1BL1tR
2Up6DT4gNsqDjbPLvrGPEtpXB0jryfG3BZVNh0SyYlkcGmyTK3kI+O942eNkxE4z
9NoSPe+acZok9x/XWvkOWtzGhf+ekQepp2uWjXKXGQYqNxdqhDfT53TCILvOJjmS
raMXeJQM8OIuc/6I63m9SBiIoGn698WaM1JweKUpM8SwRrKE5J5iVfYgcuVSgeXJ
uxX6nCUtBAgtTFzsSe0Faz/W3iB7vIu0oWenGlOecEC2Ak9zbLMswk7OWYMvCiwy
GGaVWadzQ9DqN/yVT8keHJEoqWHHYU5dQqlTATjbjwXYC3DHlmBxvx0rXBX/9OAs
WdPK1RGUNIqrPQAmZHQb39Rvq+88hQuIJ3mFrKXalZyAIv0YQuLL2Ew6RpEcG3lf
Vfmg5fnbCEGS2G9Pr/RERgaPnjLCQdqvt2p+VAVNOMfGMDTZKrAV5hp5XLgE8LJD
PqrMxuBEMNSV537p4uiMG74euRtAbL6uVvqc4VrY9WDgyN6m+UMnQRyWAH86wxzw
C87JYKEr2mOa1Lv1VkTAye5GikJs9pOmMbO0ptA7KtXROPEXAStfeIss5khahp6U
u2f2qOqJRYfkAW4IxugeE7f9XIBuPRfXKM890Wqpbypw4FtA0fp9WPGo/rCvYfSN
igFgcPsP3MWhCFjPZk59dlal6SBiQ/lpRJno390lFWP62pF+JlwUco+yaY7iJJV+
yT21qM2qGAnfVY+nbond+7aBkvciEhyekSvf3/W/iNrQe0n9OfOxNs/Fe2hAs8JA
M3xTfBf7IGOmSjR9D0Pqu2m1sWGXvGz7qpeUeJddG+KBYA8th/9SsJce0aPrNypI
vY83jZRZO3T56gPKdMuT4kPAjKuMSQgU1+2qdJfcaqZLvLpZpYBfM4jvoTHiAdwc
g7WPG5lbEXi1jowXRWuCZGBwWj3XmFw30KE0E/ZnxupoOdeJJH2/J6MJ2niS+aVq
+oCORxj4bDZPTeHJ78sGwh2zLDFJeSHrqw0J4PvS4Tk2iGbo+SLn4NXX5Tx7cmQg
vTY0XhY3s2yRdbedu3B/Q4o7jj81HAkMLYECjnN9nGMU7qsljd9K8/1JTa81tO7C
YIvNPRyjKTJxhKmDBeBr3MqMR6gIeA/7gyB+htN8ntbx9cu23f7aJKYym1nXjf3n
dLHCsWmfsIaW5z6YLNHTD67Z55RF96WoKkqgLqWoElRDKi8Ln+Dphw7DMzMrLDGw
8x1YT4BovUmNPJG5TybygVXtubfUwnAlc+Z5s4ERt5RGaLlOYMd/rM1lce9G7ByX
hiZOmKcylZF+7VThpy/g9iGdTO3KsGJaBOeThNVowlZ46Wn9IaUfV23H8oXQet1R
puUqrS9qRhV+m9/gyk30FBFmPVnntQCctnPNJ+DT+5wSsueDCsPIOjTCOO8VHTuV
7KqFxQGAtDev59r+eqaAU5b//SUJQytbzSR40SF5UrsmjkXQOqme9Uw4iOESBQGl
B9qYw8pUK+ToJTYQSGDvATiZJV2PF1AFGuwOHycGL14GyeaeVY+CfXvDoaBqn9Kw
nKkjB/dVQVUTbLyLRm6EBbN28aWpDM7BDYPoqGx6ZvcCaTDqBvvwOqqvYxM1KxDZ
QgTt2rSnk1lnIU2DTXbw4670aro/Yv7n1j4kzC7JVOTLUETewxdafSyBd93PmrTT
YmOc1m6Aytd/75sRUa1SJwVHZg2wKPH+R+xZuwwNqRUdjB8Zhqz+RH2jecoHQ9Bh
x4rjFyYEQGZLN54HPOVltilUbUP2Hlw1FFyXJDRQAgYOCXxFyX9o1ZvlqKkgAJmw
huI8cnbPKW2VhkXaFax9zl9ANEiO07R/5rsyaYnq6VgqpwW+563yYCw5FBdmghor
/4ZE5glScVdAfLtuFPOTXPeyUqJQDGUdqKVXEkhiyYShKMq4wfdLyda4c6dvrbOv
IPTun4uhkb5YZ2C8qYtFZ6mJgvkofCbWylnAIPxWtmpkSiatd74cbzKupHseYbIP
nlmQxA0Ygw/VYcdKH+fThVMxMETg9uRbUx5mIihgh7+iklgjE6kHV8rZB6ueU6uT
JSEvP+zn6eoz4R2oHIn1P8TTzhEgql95m9Xb64GeEojbYzFyj8KrDgn/9oEDVFDP
6rd8qyN12SHg25vRrJIE7DsXmfofQRPidFTzPEaiLmQXbj0nhINvxCXH72pbPTK0
O6HB+wAaw/KEFHA4WA/Fqk3/dQlj3pUilXQ5ib6feHmQ9s5Bze04mh1fcG3q60jF
NreJ03wSiUbJdnyOJR+wMajh3TwKzGMiolZi/92XLkA3nBoveNBqz0UFpbf1Zyyb
JAbT51cVgcN+2I2dg7HJK9383gWQ3SmniyCj3XCNt+D9eVMZvW+P3iekls+zOqtn
MtRb2fjALUf+pumF7KbzRA6okpksrdGIPFOxWw2TLMNCzNYVYaE+yX5GT6PcgqD2
9eNf93iAXdziVLOQLe5ryJgsJFePQUycBSYrXn5QU0FikMBE6jLOumjPoUdjmdbf
Xo846lJcNnkcOP4I+DvGsPxplFGvfBjUZP+hnmqBfstGBT7LVH00yLQwkS/FnOaU
+AtzdyXf8lOaSNZqRZel069CGaGsoMNAJvpPBowCnH2mkr5ptq9UoWWzu14TInko
OQcV9p8rIuGETn1nyIho+G491HbaChUfQiV0wsHC4r6s1AOB+KOYUaGuJJLHVS0s
vocaTCYclH3Vx6hI6zev8c4S7iVQMe51sAmyqqo3N7dy+YCl/2q5ojEPtRnIJ+SS
Qy6L8iZcSzhZawc4taeev9aTQOIO7Y3PqeVA9lCFCQ6UDLB95jePRLhdMfrpncTQ
pD0kiEeCq0nnv6UJOuFFuiH3a8eGmti44BB569n4hD9ZeJg9yRGWa6qZGnT5PyjJ
VsSNjiA/A1GKmNAcr/5lzNoK8u58A5CAe3yCULNWBCED0+QiVQVc/9GPkjthAfQw
u2EykNwjChLrjdswr2roTI5KHWE6G6RzQCKcwxjxOp4gCj2s9wEOx/QHdWCUunyt
+/ZrESWYLBNSP/5L0Trk3U7xaAaW+JvnHkIoP74Rnoa4XJUj7ASF2RJgDEll0vvF
FDDHdOvuFNDm+9FbtZbHeCObYEWz34Y+VTipW+VPSzvGjXhJbmd5mGezvlbuCqUt
s7zA03L9T6gMOQYJBCd2NT+Hr0gJzy3bHMWmLhlYpyGMxOXsS7ZwSxQybxf6g3Ox
LWYqDsfWi9yC73iqBcCjpeKa9LZ6zno+o7HVojVcBREOa1az9yz0OoLlwpsuOhLY
hFSUoPqtqThGHrxGllZDqCeoxIIe4BHPpQM7ahU58pBg3W5GADwYitep1hP/HfHz
j4pDs2K0p/W5q+D+Z0BOP1wAaomrcbHZDIqCcNt+BQUCAbVQorrGUWc0VfCHMAn/
8YIrKe9MCBHpSefnivw1vRl1q5laO0w90WpSrOlt/CPHzFzEJ4vUScxWEhgJG3qq
QmQRVMxlBgd4BakDKd0bv47iLRC/9hkNO8tS6jZ/SoQzR7qZHr/UZXsV6LKl0FXF
qj+Vj19u5IJLpMoOh5dq1q8jXbRebMkk9EBzi0NGIAZAZ/a1e0NwPvvjVP3ORet6
Atu7nG2lIQMcqxLWCWuvUoodURth7hPcgLms9ImRMK6Rd8j2KRWA8wTCCvJkRg+8
VLjU+9JOLzlOdT9YzF/KEU/hxfHt2mG9g6QmKXhWf+GlnebPH+EwhYQargFmnQa4
j8vWDnlYeR0NubFNtBnGWjudW/p6z4Vz7fw46ceRvUbKkZz8ntX7EJMXQm3cV14N
jzJY+/ktBsC8vz2k7OUwAeThkmWlUpdJXSHQgn4+h87MoFAnlQ9izYTuTaykM7Q9
RlC2gbrXg6KaqcHN80FR+biUpGntKTxZFSYB/0tSd4BXzEZJ0POqzxCdo/t479dL
U77BAR0xcPBi/eqpSA6mE+DFOmlyFXxOnMb/M3ZwOeL0azh9Dk76VquCfTDRDVBJ
ScIS1teyavO5DKsBAZff0WQxOpRpeUR7Q9Jk1A6agRa/4UkDo+i9CxjB0nq/a5j2
0a3RGugHfoaLtVZ2EVESOsIAVF325QvpDPdfU94DLRUlS7HlSj7zjYyfPFiTrSBc
BifqE/JWzrtCcyqrUtZG2CktQyTi6WX9F0WZQu3CqG8LLE/lXIeJYD1cmE1e/5m3
SsyP+Dd/wXm8ddWvrkBU4JSefSsYOd92n9GjnCcfPzbztrm5Ov0UwIex0Ux2MZyB
I1X1BNkLF29iUod92a9VK/9MiUKWWoSWKEKZAmx7U5LCJPk5/eXnFWpmsmve0e6r
35jmifQNE+520BaWOKgjdG4u6cdhQEaUZiC6rK5cApY646bujRol3XCmTHNNX8/N
IH18+RniQOYIeEvwh78g5RN/ER5Cagr+hq0gvTh7cXjWSLzaQAQ7gsKgu2Gl8FvN
6bO8S39OxcMCNBwU89R28jV09m/S78CXjAMDYdqhpUMn/AHVQRehzq0Nedbc09XX
eeewLVaIMDb8OS87caTmdkxAKFl467PAIH9rMj1fQEjevOVxG/jsxPWELCZ15vLX
e45hUwtMRSw8/EvH17g+Hfb8LcDdBgf1fxYGAyVGgwtW51Xjp4LUZBp96i3yCxk/
s1TupdHfQ6Zav+PTUIoipUAYtXcS8SCcWvsSIrF7FaeFV7iiYbPfTuVUdhZjhxIf
oFdJXH63H/M+gPXll9BOkHJqu9BYj1fl8dwOvcdB9ny2ghwFmWkqT/WeHLYOBFSd
zHFqhxATYzH2UmaYfLzGVt9b5dGpWlK+4/SHypKUGt3SGVSu6Omzu1sFWKyM2rbF
AwZ9HHwMO+PNgeRyHFvT7CEZgOKGkjN/MC530IWmqdBr6H9MZYINBA+KaJjZ/85i
HE5Sn4qOWyasY/RDH9Vostqbb/P6vAyaH3FTHR5xG1jpwCX/oc/8y2K4vbd+T1FT
A9/azAkzFvG7CeHdDPKII5kXouHs5MXb0G1FkiLKafSmaEf3/Okl0lUZ60Q2cIxg
Bj8G/YUm+7U3ZSKd1qNFP4V8eYfeVhUm52bDG3XDcWHjdJwVpA5uS/0SJOJhx7Er
iw6812wyyePRUyeyH4Y9MyxguyE6L+5flh9onMuHDhGdw0U8h6CZS5kIDa/nT+A4
T8gBFmM6RksSyxQm0ZCuJp4QztDPcf/8/+fS+kq/U0Ziqc5nXRFhQF+tuTSJqAn+
ybr/zpxMmH7yxRVQ14aMBwiOBDTeNiWfgGIfF+52xUEbVV59Oh118MNcoCbcSE+5
0ULheiIazI1/VOE5Y7nongJhXeX2FiwJJjFpRFyQ/pFl/rGt/lFsEb2uAoQ8Rf2v
Z9S+8uXmeFbh/ytZs7mqoETcf9bfS1Ns7DnlC3hNBCzJqggvtu711k/NiP1whiBQ
wgkezanxWlIUvvKOXRvXfXHc1Y854VhAnaemEFcGeLC7Mj5Kh6DwWg86ITXLiLOc
UMfEhBMloFrYTPNPx+iVW5oyp5OiwI2Bg+fvM56wvmEMAafu6qT09z3V0OuXPz4z
SwVlLVyQQspTOXOyQt8UzMzbeVByCGTBL5cfRZJUH+vUmOfz/YZLQFpkTGW0Tl3c
FvYVO0Lbx8MS4pLS8aMC4WUaZqXonN7ECiOUrNqnR3r8U13HWGY9bljBrJNH6GoT
uPdWTp3TvA1ur7QmWRtzXwgqiXxPKElGHaFAhaw5uQQ0Egd8ff5ve2YHcblU1jYt
QKkTkVzrK87//pIjKpkvwb2RyiOp1mCb9bKTjxprZvtlMT50p9lxCx0WL+WVWxP7
ZZm40Msr+mP1wj27hkxTS1kOjuzSUQNEOhJXpBFtJT3bD/3s8p/o8aMvidi/4WOt
eZvBBi45w1MqluvKLfgAak30cVxEisEAe7s3hcBXS6rgJY+Mz2YDwDs0BdjyuwnG
VfNgwHMR3lCzpwSuxRIEvGMcZDuEmLpVA1yKkxcg76vJrLTE6W2ztnqcTKHiHVIb
7W3x/6puUf+cfM44QThz40jRa3qGCdk69SPTXU0lNkxcR4hR3TQHqqRw98YNQRr9
qsz2hyKLZslPEG+G5SaSRxAmzL6pVySn4g+GD6pn94gTT1wgMwCeMjihKps2WJkq
z7YGv6b6AqFpGeaw+AsM+8ROxcDUigKoikec9bLarSWNzKEokxWytKn4IHWGRzJw
j7Apgyp5zos73JMDqJ9OSQ04zTNgodYRINxNtJHj6/wqoSsqAwgGUQU1brFB88bt
UWEgwhSU2F3DQXyCknzBsBeuGfeEO1ZhSKa3V2d+EC5fHHZqUI9VUMoAkXUymFU9
NiJ6VSCol2acVkHbpR6b9Idw0rNvdCe2A88VuHx+IPnZUbZOJ9lNwAPPr1gAZqQ1
rdwqyJ49pOuhK6txLznqt0GT9rNbHzWDxCxIwLRLaC3l35Hu0yJNXbgb1F3DEy9G
Hp1+kRuPVuBEajkGTagO8wDOOtHRALUSPStJr/YeuGwTNfSZcie8MzTd2bkPxoEh
Fvvjr7xsYLZoKcdGBYOpA8xyLVmCRDM12Zmbr5f+MHSvkwxRwGGACGBMSmxjPPq4
aUzLfBDnabuXkjL3sa1cYMWLfKcti8jfe6MKOxBDd+hY1JO/2qr8NOqBMwjdNJ3B
Pf+JDdv2jvdPI6TJf1boYu5fzeagrjga/mpT1FfCM6U3ZqYS9X2OmQdUfQut5WBU
v0HsHUiy/EDgZLvb9m45qrWYNfkxX5AKQB+4vG/DfjoXIDYJA/EtfWaozbEOxO8F
6GXyT3epVn+CWOeTxeWqdwzi3OJaGslt57uowe1lh6zTXfNhuHHZUGLuBSZ6zGmq
l1wOC9VUe1NXabbtu8hoNaa+8aymkCkvA5+jQQAWJ/OGVJ0J7JIa/dAWlh9ZcTHa
oe/c0rtDDkaPl+PNOI6eBkeKGXJIK7BVbPuF8QsMfLfn2H/e6dUn6rhOoatxFTzX
DJ5Ty+r9Z0s+gvzMg8o41v9WHvsswSL9JjjGEOKoYIxqvQKRUbSYBhxKuL7tc9+O
giR6MaR6ry8TXcjcK5VJs2Y6bahKYNeH0JmBIpJKzVorWyU5LMzIrGfNlhQUg1tP
JhSJ33a0jdnRjTVkfSyKwk7n9nR/I/0wk31to3Mz/RbgPRXP+6qZdXMqkzSVTvca
5dX95Uo3st/W8VR4+Ogk8s9eD4qGm5Di5S+OH7Ps+mKvBfqvRvRh75vSo4K3n3Pe
nXygP3hlR1xcJ6lpuB2aPJMrMzd38qE+pnZygWSRLi6qLm1OmgUg6rt0KJyiwTRb
fRyoG0xI+0LWPq+zBw9mYBe9+QaGZBD1E8MBjD9wjiYlVfISl2RrET5qPiJdONF1
GlQv7zv2ogvj7hLQ5JzWEBtrhho5bxI2AFWkY4CBfX8l3SBHnt6A97cpTd8LDdun
PS93ZxSch8Dpk9Nze8FfwUTN+K2r+uO5ZPFw34z/57SFZUMLHHnxkB5L2oZDmD7l
oBiwkFbFjVGMxzgN5C8o2G9bEGUJw+Z1i3nGIE47ebuEmA55ORGHfXUb9JdQrRXw
/l9w7Mpn21P1xrGTvD16fryn4ASonDuNgRVLH0DAe93OCmZmmBk8Tcq8SEmKbVGx
BzTdHEjjuDkDNXBQLN7u3X58WcH9VGqeH7+dSGuZtUxy17E3B7nJPr4ATRw8dfmF
XwY150JupzRO9eh6/18hy2OvK7bTKCdm16S4AbgUaSIBmJqvYlpBNysfr/BpcW/V
jCt9QlwNECq6lM+MyJFsnI3WeRRTsCxBCjU1UoTKPAyJDZ/Vqe7NriNg+iUsnaWU
gRHNocjL5eidt+xdPnN4WNDqwCxxgz0uAgLe6g0pvYf13QImga1MdnnYu7rkqrHA
4nPdBEcXs/JpVKMn9UPl5OjsNcelb/UBzOXzetij61OH1e3H5CrU7CsrlFGhL1RC
uhXy8cRx2+tsoxgltC5bUb431KdOMiEFp7i0+w+oY+xHobBWMe2WMMzNz2SHNejp
XX144i7xRVtnsxUiyFyAXMZNqpg0tfBNtbyIlr31xKRDQK9rhJhRAC/NqeOwnhx7
QdNTssxJ+vqnHrKs+v/wvjaIsWbqsuRHu42b0CYEiQo3jCOm3V3zeq3kc8rY4DlT
krhbJgXns3a8EfB6khk06FGBLRE4eCk+mhAfUO9lDjNd6i4CAfsHbeu4xmkd+2Tm
CjsCbO1dIgG19guDzSCUfwu+yiiiEMghazZEZlNhjH4Sb0V9BYJRrO0Gz6pBoC3j
HQx0+rIEKnU2IapBz7+ZFRpjl740M8TNLY6ba7W6l8SXdsTnC+esp0rNpM5Bfw41
6QeAD8gj61O+KD2zqBtKNcUE12UK6XCvYG/jzmhwFioENlaonyjnxmf6DnKQ7ccU
cXBouERHU6NjAjorRHJY1H2bVtmcak+1tRi6OIXMta8m/3Y4KUgQZRqZH7P14pCr
bPoXdDsjG8XsP4N62kklARP2PEnq9W3Vnv7a1ZvuXeQC0y1zlJ7EW/5nGvNscOOH
r6Onqg416sEEU+Ae9T/6VnnmI95Dn60ZfO8ELrqB8pKTS9zVH2qIjBpZBp6kncp8
BAxBRT0pS9032/e4ZPaxS/+gV9VxSJ5QUxUq3qFkb6ZFLQuUCsBw3Z6wPDkdi6x/
ZjtAGhtFsuzuR1FKFsMEo1XF/7wh/Ix1+jJM4Zo2LiYs7OgBvZOhw/JjldQkTKBw
82qmSktnekq/JplDI57+j/iBoLYKk+gN/Sa375LdZp2dLiBB4FvzokJEBV85Q/3h
pZjOYf81L7Jpf4WnL+0m3FVGR9XpwiPVJjAmjCKqWtw0BYq0VBTk31YBN6NO3rDY
H9rmCA6bAQboLYMBw6m0xxA5eyoUe1+3NalJpDa6pGlQKAcl9WEc0Lae3PWHu85B
LqVe6Ogt5KGP0jcDoDzKlQeYKqD/vBNR8ZOCTe/f/XzewEbzy7HVZYU5O1rNdB/c
edFcsgicE06QU95ZMLVZKvH218V5wF3R/N1VvQzMlwThJTGZN/7J6/7Nu81bbb4N
qtjr11uE5zyisAr049D6zAs0gyjrXeIF2d4nDGo4xfYngo/xlba4AYQyT9Vx5bAo
8mfctFLl3ykoMSYEFSvQL01PLJpK0wb+qWp1Zma7IeqaKoILchXJkZaXeMkohGQR
i2Q2cRcazRj5dtklGEobrEd1/0DQB+gxQgfp4pz1n4agV3ZqgeP8XCVuGYAI93tK
bbIpIvaLUbD0Y1+wlD2OaaLje5SJlSbamdP0VGCmkivu2U0GWNodqWrqhxgtswmd
8mYyPc1sp6mgLeGCycjbWMJKbtNZsPwTtQK6Ke1bJ+HbuKVBh65BhHW0z/15jNn5
peKzuLjjbDoAVXYf2SfYyq+OXEd00zytB+U2L2zQz4FLfLYEFfAbEqj0W1KqrmBV
IiK9X/6t0S8awCAq/lAnY1X0Oc3QWpVuOijJdm62VUW2Qgg00WZ2Xkh9Wf7UGkr6
5AJf+z4wfFib6Cq+V+Rnywdx9qLxZIhPWquh2wVQVvz1zOL+o7RnIo0MvtVeTYUd
jPSKsE84XUW/GhGHdJLyVpQ6Ujum6bRvzLZ8HjeH6mRUQAdVvt961OluiO/PDO3L
kUFQnCX0WHUa8F6JdjAb8wqGD6Bu6Q+1KjlNfnhJblxDRZNlwQBuWJIWJ8urQVAv
f8FdBFXnzIe3WhlZcFffV83+LfYRXXYUWc9c7CZOiDedRpQYwtbFMZA8e9vJ3j4g
JSOxN8zwqQTetzngAPXTPoLCP80K8awD4KAlrjbkovidctDRP19T6rqpoH8VCLPT
+4v4LaujMklutiFn9N/WWjPWtTfhzJvDTcoDCURJALvxxDxZV7/QkcqJMcde7XwX
+rqjypezGLVNZkp3VwB3Ty2kVGWInVszkF+GOlVcIkB97qsbLA8jcLN2Y6nJ86VL
/ehDVVdMUP25z/d7GN+ZPe31OsdTqecmaNf9j0FrQC39YkWv4X+D9lbFijbka4S4
GT9RRlVvqQsVYmGyZaDFa4OY6M+kC1Anty/ic73yu63ouefVC9rjdwvQ9n0sJsIo
LB4cuf8gnYECC2V+p3SEd3wZ9/P9y0ZJPLSZdTmFUYPG7OXHNkFAalipKCGzAv4l
jCRqFtuHYjRyEl+kif9VPi7gHm01ZPfeTIm6llPqQEsKhEYxsBNw545oS/ax2QOO
h1swAXdBVZY4oASItBZRyfX87xWm68S+m3kRX/F4Vn0ZGn7O0bXC4Dc1hGkOXnFA
yT1knkdXJHeLy0rOfeMUQRY6idOhF9bGcN9dAOKE571fT/yBQqHW+99fx6KS4rZo
RLfr3825fngrsgo7yFTSW/uCTqMzkcFFr3e5YHwetLstoc4abn/cD6wyFEBR1iVe
N5AbsdJiuAH1L+OC25wNvpFyUyLCRatLkmHihyohHAuQp19lwsJKf7amVCFvuzAx
+a8QqkCdJj4A/LUOfvPNg87PqNruc5G1+gRPU0DZ3SFab8cPviZDF00NGZNaoWhn
7muV5/XCfHK21GdDabYOVCZE06CJMyzew6Kgay3cHu5U7bBRO787EFq4Pv8w1B+4
sussimcOYz4wn6qIE5JGE80xYI1FDSVSYXZIRuPIAYFUA/VDxq8n1wJibzOiVbxv
rmukRCY7I6c6BnJjEkkyGwXajeFfWVaGFbBW1cL5MSIyjzw2yVBADYXJ0gHfbE8J
nxAGoOZNZr94Jlnm3SC3uKl7XB1AvrTUBuSytt/ZbHYY5JIsuB4dlK7wN0xieAMi
UbV8kJJfOYOvQNkuLfKs0G1giPuS/nJzWfgtiU2aYuLK6LjJr5F/BDZr51dK3Cn+
A+tXMxhVxZhbAIF3t1ua4t+V4x2ATXbnlx/o2IXfjQUgY/j7bRtWJpVwmtYhp3Be
yXv0Ksrooy4NOF95UpGv7QFIXSOHfB220g5Sq3oNWpcGbBVYvLp0S0HAZME2UURW
B3DFWXidcaGUWQ6/GyvgI8lGDm2Uh7UlFnKcVa61mDvDLRvTdIWNdHY6wkA/hu1z
BVl2qEOXPYRihidnz8CQdyVsDWPoefLq5J35DwOMVMmpGahrrXH+E9UyT2DMZ5fd
Y2MZAx1LeuLZFrdq1kM4CwuU2jwK9XQ0P7RDeDuFeY44BEv96gYy5QHyGvKbeV7s
Msmh44B6/X+CHxZC5yFoQoPB7NUE2zMq2clZnhhcGemgI8415XNSPXXvwGIayjuO
3MmGpEjqzlulyCOe7dEJ0mVTRen8rJHeeBCTLj65HthqF6PXHtcKJBjLyfAYksYr
eDH9haHbzs6yj42/CfF6p7otvby6eMYgfpJk0fJq+kVhDR8kseaio1upP1Rb/Qp4
0Z4zvA2bc8uhDwXV3dQWP+BDAEZFiGcizB2nPFbHqz/az7oP8UqXjMzmqiDO2Sdd
N37IVllgmyI1UUj5nCB2IwSDftVvZ4Zyjub1tpQbYaXbKuilCk8ElqzHf6XBS2bN
sG8TLab61TS3TMbc17f33MNn0+yZ6YEPkSkJYo+2Ulk5QWjEqEqq5qOMrIFFyStb
9Y4j08lFU67dUtI8IgZQ8LMuPrHmTdEQrBO422SpRGII89fZzUWfqr7IAqvjdC8x
Lh/h8q0wQBTvcdbU5E97MnBceLbmsUgjMOa3d8szWdBg8AKViH9ZJiMZHvm6l1tB
ylp8jJU8HYzazprMZsGw+7l0PYOtqqEbRnfzFK++JIs7iwD9LKXVNY/oPBCY0TpA
sC72htY/iyBOmjZ5IBrW4/ZRNSgL8SckTzs1ccffXbhlmzKJyxxqcBxSQUL4F691
TAcjwS19Xe6jkcE/AeGA8MlCeBs+s4j7k+G5KiEfGazxiOxIgzTOZR4OfTgVTdYE
/SVxwNxJibzKJFdgqc4XJ/V+9xUMjloaKprWMiMb+ddpUDqX/pymyjAX9Jx+CZky
V1CM30Id7PN/SRYUfrgXwL/qU7mOCCsWU9fppROfK/n3KOKb1VFobjg721Lsj9CI
YDa9H4S1/FxDGaoroM4JeN6DI63a+Yb8677vqX7+exLuVfkiAIV4tiS+zHVW7IVI
Pky66XAJi1cetSf2yo4rmB1NrSBpvOn//IaLwKhtH0smhKxC+eTX4wFQKQcQ43YP
JEVXr+M4orzxZQDeWN82IvqsXPDV3rTLHD9IRw1+olNqUytn5zqPW3LdE820flvn
hGUK4agHL0KqWhh9cFkFNVcBqls4OU25/jjRCSR4VKM7qPNp6ecIJUoIDjeSNEix
i2dNyTDQA6cniWdIkMGrj9C+clPHTI0MXYlrHID2MzCSi36qY2uUln/wramUY2WG
ald6niHiA/rZvLFW7wCJLaKsDd1REkYYvfJcdq0R4DsL0v9IztUrgMvUvo0Cq9mr
byPZcHrZB4PLsuUrIqKTe9gHMjEjgguT0YPqzPvS8NvnP52QAXHeuT9SYv11LCDc
vc6yhCRu967yNz9b42jkL7kwhMoUQL8RS3akoF6xkv8zbeQl8pk/sg1uLRZRZIQx
K1Go+9N646LlhVSUgDItwUrR16qnaHztdwL51qzeh+B6Tibk8o4qGU4VjWXaHc5A
ehlDs/QWR1OXDMkiV6IuLLgJC/SXWKutAfOqaNj10orubrx6hGJ789XZGrl5Y0Do
BuScwcWcAIuNBDtj2Uu/JX7HODagvH6QAAqZFDHvR5+aqpRIYBecr7MAI5krnay2
4OcCNd7gp8aD6SEwgYLmBmwzcaDguEPRR8PRaqqXfaMt7jR1fpWJZr3LhNWmH6/P
lJ1hg1/xM/SN/syOqi3sa0ala9pNHjMpAsrhvqcR3U3Jy+XlNUBh/cG0ANbacfAU
wVzmCySUnhh4Z60+Pn+tNFgP2L7Tfchkm84V4fxn+n1r5eEjvSJ9ijjq6+LHZKJP
Y4l75EPtUML/quadTrbWRK09ZEt5DtfVGS9H3A42V775m47UvJdxt0Sz92ZSnG1F
hWrMkWZT2sfzmQq0T7821/KBUtf/EGVsrXiFH8Tf73KVPvbPkrQhQtvVNlY+DfXE
hbqdgs8XEIQMIjk0WQQvF6R9ClBwInCIa5sVqAq97t5Eo64N0Qu2a8aZOrL7NXXF
BMHIrFF662zG+wtwddBnMw3LOSfRzqpd+JwzyxE3csX9bszdYPShvah4HUIhA8O9
0a/jfn5hEXClpAK5Jz8bPlG7FzjuLLBJ0/WoGeO/D+f93tFRt5JELo2IocJZWR7Z
yD3Ex9+iV/9UW9Fpl/OnsBVLm99COzIF3l15RkmA5WQv2nAY99sLHCbM0wHM/IGs
05AbpNHPFpNderb2pbkFuW304CIoo/phAWAdLV5uhl6mzyLqmF2hl0iiCR/OC7V6
BIJfi+cWHHFeqN70Ir7GHaLT3NLpxLWaT66sulScaW5aumsXON/wZl1JfAdvxAUG
Kpr7eBWUM6DVZXKa1xV1oKd3xyjefvY4tg9bH/0F3QWlWBDujcPWuywi9EAaP6G4
ptHCF7kaoSe92uN7+42rxmCTnGshmPQBs8nBLLKQUwc0UO+mFsUEJ35iOvF6udU+
ulHRJz0VKLL4KQjrt5ZpCtQF91Ae2pwSKqnEWCODI84k4NoQvXO9DgRRTqipS/AB
hAQnQbvJr6kqNSI4KzNdhjcJQyWDtJfZDHVv2RjzCqhiHxlEgvEw/+C75STAYzab
c/Ss3rgrREZtWFinhw9b6gceqTdGQm/+8eNmFSV1ENVBndpiuCe18x98kpap4Bxj
YaXhHYcHF9jRboM1jFiyK2BB9jF9E16uFVac77bbUjFmui787fCvV324n+eT/Qe8
ehw40DXJK8VY265NnU8NMZFrs5Lm64jycpHmDxzWn/qIMMq9B7VQ2aMwaJZcc+n2
qufUJ2OY8DPXUBSYlvSnlUEmdkpEC3quSlADdYOuui0UJ/EchyHn7D/WPEgF0R2c
fERMRdPa6QpN6CQQEKRec3WtaGsCn98CH9YMlVZE7z4XbyRMGdLPooyXp7RODhsm
iWFOTaL7DJBTYVeNXQOwfCdKIIy/QAq566pAiqYE+9ERZWTHe/epSyyV7zWFBjwa
pFkcIPYOzdOopA7MWgxGhQpgaHP+4Q4dUc1YAlkVqH21G66JaSDbAi/zn7meWCxX
m6dByRNXprarHDOx7SyIFe0kQ86PV/5tmqcExg9Yvu5iQMin52OCUXUVWNAwdkHx
lBjj71JvQH28iXdnY33MQRYttdYa7viD+ftSYxdxIJpQ6AH9bnA2s+LuccvJ8hxN
MGUqX9JU4CbVTNL6KTmWZWpomKxj04jYCen21fwaqi2tbqNyjOKX8+u7CumMW2dp
yz9AFepg8d4wG3aCP6f8AchAXBUOHZQvi9FZKdQcYeA2ktc8sljT8AmNi7HQn4ex
cUXMopJhUkoX3PAVbtk/Q60iKH3jePIhU22DCW5dSugS11rCR+Xysl9N/ELKINGn
QChd8FUb5qpIZa/sIMD3WtYV5tF2lw1xstJRJggoYJR3wx3wrGTNE52Olm8gwKIP
x2ih0LZrTPMqDfKuMFjRxslD0y5auRaQ0M8TT8GEUjnVyq6GhoJ1gseiWi8zCEV8
0q42ZfxAMQaeVZcnA9HSP9YUZAUFej+2ayacOpuRkFaxhNY/u1gloPBmdeNRmP3y
Akg6QG0keJVKYYc/LeXP5GEkCLxT2O3mpwoNb/fINhcckFSJXbswanez+kDzfhOp
KFZQ/N8eDC/eW0+GdmrErggBR145hGgDKUFxDj7sXvkp6MNF3XcYSOGJsqPhOSCD
qK4V257QOw4Ia/sj4ng90OH9U5aixCTsTO2I2sId9ubqJe1zpS37G1/VNnGOmdAv
Vh+ahdFLp0f7jTfw/a9ZqJJ94UO1gj7V3uFVxfrKLcvqSZ/6wzjwm5kkg5+EsjFf
pzNbXQ24VA/auke9cTX1aIxh53R2v88DJjCeNVPig8/OLg1BMo+K+FXy7xK8IQTW
1j3/fWYQ/ER2Ip0ihj/xDSUTgWv0xXn2gc0A2DN+dp7dRwIaPlyb3M+3+vI9mBPt
Pdh7VapfDQUg3ilG6nZC3r67U0pVoaxefr26WMha7+QutmIEYU1tBPDzBB2GfhHs
J+DNTNZ5cM66IXWUZMjoEjFP6l1iOFV6VGSH7+pyPTYUmFL+uTDI+2tMESJ5tdGC
O/EgCKQBnwtDz6MSD7VdilodTBN3CA5PlAbMh84PgtIF3tgTN4vq+sqddXQjryao
nX1tuC6I6TlRLJ3ANuSse84Cquu8cK+zJxPiIxdQ/fB01YGL04+gbxOkVbWlWGb2
0VxohU1nlvBfdx2ytMrYvJIzrTdTVX6Df4KkW1yKRwWatVVbXcTABGhrvDNHCds1
1Cw1QPj1Sf+L4T3emDVtOgQg/0BWDsy6kg92wmu0RaeYy9ywErfqpoJgdFdPQ4KR
CReW3DV2DVePm7fDSq1W6vaGS9Tof70aI4ccV84PxMTVYNRoTTIqh0wLfWt7vFH4
Vz2ljVRfVlkv46rvzQl6+DsrQaBd9hFzQTShVlaOFYagOHHeM6IK4aOnpCDA4iJD
+k9TQjXORBrmE4aowL5YpSfhFi7rjeEXIMYquGrpZjeaSXu38/N5tESh8TrRcWLA
nB0Hi1a+nUn5EkoYKDhSDP0qw9/yPspO+CHxgX5/VfKO/lZjdIoLFOJrjlmdmJ/x
dFXnSN0U7wxcFXuEdtJ7RzPTYvkcAO5bEtAza8d+cqkA8/YLew8lVu07jMpfhl4T
uFjEWgvZNHwRqmXCWzCrLbMeF2w+twVY/3OThvrpOs+wcsy/7lloc3rPcKzbm0eu
NNExP6EATizUvOJ14yuPDmTTs2KdlJvviNn0PvzD3ofZnrrfBOhYzmXGQVTGlaT+
S+BKyj0zQy/K2VqDlNRruilsgIAh/uyHy/lCPSL6YeQAfTuPH8Gq2ON9uKPtzG5k
V2UgS0bKukYPOInWWOoWuhRPh9Nr+t2m2ZNrDwvmlhxHFRKKWk40HN8lZLsmSDFr
tlpbDftYmCfzWK1bjcSVAbAGGpSQsxx7cBLgg4eTh6diORXGyguU4+6WVwHLPkBm
sio1p9Ww63MKNIn1fWdEwK2g00NOKD6LIDZJe1cXLbqhWHUvWIjqn+5xvXY6bq5k
uYssRARQL4PuNiyOh6VH4Hrjp/4bnx9qc/KI9xBhIjIf6Yy00CJpRA85fSgfVd6u
cLdkcj+smM8SXd2TdIVIcm1ToObQtFhkv8+tNPPLttTjIEsxVmusgd2+vEByD0gu
8pOaPg1YRQJ38kL6MieMK+6d2T/21Wfp83Un4lAVjC+pA/AhQrhOOIXaee9KIBG2
Wln/xtOyzUEfXShu/wGVHQV1ygbf5p93m549apNyf9X9byZeuEbaQJl68V7v7aTM
L+VnCNI18QTd1O0juzLsIZts0D5UhmRlBdMUKBfb0cOEM65UUHqV4Ia0WVV+tkWE
LT2PScUT7FS1cksismWLWYW8Xk0//JrfYj37Cm8BtIqV1QoRP2io5OYrZ9E45dry
Bj+1rgqRjDQn/kVbRghe+oJcTcCbgtfVAEGzPbjqcnJYoqpc3LGjy5k9JFQZYNY0
8hXgZCMVSQ2eztVRSx671vuq223QfGXatCPKUs6kM9DOa1R0bEW+QuiGPWlUfGvb
Zldn4SGXovIM0Wpwf5CTBJXsvZGToMUkWTIZzGD2ox1WKSeem3ga89vlUUEM5qDM
Vy3gKcZHFuY+KrDay6od0xMCli0L5YBdsdagPcD9m1BvVQQ1LwmrqrzjA0LryJgO
h1MudaNPjYYBzAVoN7Qjwx1qZ591ZkS8oKrzc9LPZb+vIUQIC2W+xUJcGnyMUGZd
33xRZnml3KwJHNZBIMC4aXGSjMoKi/e5HOnGVtaK5ildF3aevMIklh1RHKPytU/K
zV8+p9guV++dLHaG9Fdf7DXD6mqGdrvT+HpxJlIGTrfB95DXzuST/FB1BwBvk6Ql
JHUou9KoD1fZql+zqR6z3/xSBoBN1CfDefGXOFmeTKjiMpBGR6ZTCx1jfbK/sybm
UFOZSF66VR6bpH7kgylGG/0/hRLi1MefS+GH4jIJpCOTNTU3zvza9B8k20IJJGUB
CXPheFSryQwT1LfH/RO42qfxr8ItFMQP4m9F2GyNrmUPBWW+WSAwPBzKD+3WzucV
CC+fN/7L0nI9S7rOXvCo1XYFsslBMidXqivlN9DOQAUw8GLEHk6Oa84H0ORKdN2k
C//eCfexTqvAaySZrvC6MMohVf3pwJUHkPmohUtf04OWDeSkWS8o/iaxqrJBRR6w
H3ciPcfGn0asBzTqs0RkOksrAVCFkGU8bZUxgFu5O0Y937kokw2kCkfd2o37TSi8
OT4EgRBLbkoe2l+fCWiMKU+0p7udRExeBpTEj3fuKkbvF6DOXQrnVYZjvdKt1ZV2
YaJmuQFVPTEvqL9Q8s9qZE53iAFxx+4gkjNN+91ZJSGs/K1L+Jux+XMUHpzufpKh
j1bbICVCWtys61gVJo4p/gjscOg3Iq+EDkT7JvctwTeH0gHk5Ds5Mvgwstb5H5o2
wBnpqkP/Mo/EOW1aMIgba0rtCQ5yYFkKukvLZrWNrPx0vWQZf5WQHZe3Fb64S2A8
xc6ff9wHJLFLL1UELOYJo8Kv5IF9xPqIHd7UMCeu/oOVozmH1WA8XbWzv2dp4/P5
1Po6YLr1Tyz7oQix5PLhujkh+q9k8zr8/DuCHzbubHAr/1bKn7Pg8c40CPIxY6Ze
SDZXz1r6D/IFH1C2cwgtlsDFDszyfTzl06PTQYFD96ppzEEcVINQaJ1j+0K58QJd
skx9sfOWdZj479S2UTPvIyw3inoiHnBI6yRphEblKu8+oe5LjXs/lT0y57vR8RqF
LWH+z7MCo4wK7scFN/KM7zr2G7vT3C4jkd0xkCHvEHSgUMikX8BJieJ4nZcojSzP
pgTYy84tW6gEOvXHizOEXV85r5dDq7wvxFMa3mlnS+uDffcgDALYVxnbjqXfrrUQ
uGOY0t8wThTCtoh4L90g78NWJtP0Qm40mrDrF8TELUyH4V6Om50VzeCO62pO4Z+p
JlqUG4GT13oWR0dvhExzV0EuS+PS0JKjVkDKcgAuQ6+8VKYHgZTUVtvF24yc2B7G
KmO6Lx+dR/7CM2NsEQVtnnNFDHl7J7lNgwqao1RJGfsoKOOR8SPgVAOR7eadrFir
VNIoed/4/qDnfWrQYjlPSFICUTGDmqLElf0H49TzrafrEvb61DPsN9nLYPQK2uEH
6GH7z4XkcNgJueDQozTf3rNgSIEK/o3rI2uXm7YiZya/FdRly2A7XzpnGr0q5mgU
1Dt/p1/KhDbueP0BA09LNT2q+b7Unc8R1NSyWq0v0Kj0uOC9D0ipDdJKnoJoCmva
43R7G0gMJeX+6y2s3E6Bs7bZ/ToqReRD0OJYfMrT3yZJq+EhN6OuOD27lDxW1rLY
ZxEIXk6armUYqDzAHF2XjnbQf0slYY4JtieqVI9k46lRKco/4PH3SRT82VHZmn1b
fRYqV8IR6YQ/3OxZa0PZQnWCkveJaDMDmT1PR5ZsOpAMAZ1Y9J+SUo3RZ+GPnc0F
x+7gx7u7MMeMHUddKGvqQfx3ePGgmtFu8Mv/RnWd7EU2eORoV55sSoGkM7+PQtBC
i9GmGmC0atyuIHpFt9sKeCh1RGJ9Q6JOB5R3fh3o/ypZzPOEMgLv9ssZRdXM7cCG
sUYS+PJ1NYZ4OZ6N2gb0W3sZs8Qq+CZC8OxO7cMTfUOVHa4Zell2lN1JQpip7+7U
bGct+EDBl7KfLQ3lsYWNEe21doT4X81czO8pb9Qm+0N3uGmsjRNMbTbDkGzJCszz
IpsSjAdpxOpWGYLWqo+3c9QJOgGbKYogBQyCSVHVa3YlLdjdoO2HJv0W/xhIcvPC
HyfWs+kczQyflNwSoo2cVEXizNcCssc5gVs141Yo1q/nZpZHIUvvW70rvlN2llVE
tczWJDQbn823tp9L3/eFPqsSdSZ/U8/qPm0PvXyNthofD+xsxCgzefxZEdQ3zevd
G2KdZG9PUO7M8loAVsMk+RWg0AG2nSvgAuwEjKi9a7Sz8m2pIBt4q4r/1doHsUw9
CtKWFRMvepmA1CNZMVutKG6pgBdWP8K6Hn7qcSXnfHGxJF6182IWPA0YoAyeNk2X
B2S8GtrJJ6o1SYrTgo6OHo4vUnx0csJBEkeJiCRAB5fTywYASYhAlTXvm12rTdgJ
VynAY7P+jBqxiH3lJ5n2IVZBJXtCOG2lAKYOjXtxGUoXqitK/30usLiIPfkCR9Q6
l6oboOX/lZ4L1Q3V8e0+pIsXCmfPpD+7v4if7DLmbtzcucpxE/dDpKvXFPo/XlxZ
05X4ytZEyKaBl2JEKxiE8N/KqnpUC6V8ceG4p1G0GB+FqQxAXe/lNzuHYkdjSaOe
SRqjYoudqq2O2LjhtsTRKnPllca9KoLnnYMDO4aRNDV+S07TVHGY8uckfCRpRB8k
wlYiYDvTWDlnwBDIiiI/MmQLRpahmUoZT3i8cYiWw/YzjADxLm3Jkpt/Xob8nY+Q
fyBc05EAKlcjsLMBoFjdST09UtMqu2sGnwaBoH2KvZj5JKUO/EbdZxRauUY0F+Y5
Swn53Hfv/0+TZz2bt1vufmKx1GHyZDhPRcF/7uPPgETiGnJf1Joa6Gy1aBGdgPrH
vdyqvwGYTJ0MTYajkQco5anDrtbSQBJ41tM82qPGoEhxcsZeXExmUWff46RKPPBp
5lMQcpm+bEbdGKR2S9EPp5zRVgtpIsFoKgMAWpvJVOdqwwLgFNoFE0sGQ6yqMgEJ
/9kKDKlqZRrN7wyu57Y/pRjVf3YS02ECXtK+ywoGIvrWjBA07ptK6PCNOcTRXuQ5
Sm2sbit+i73kjfXGLdmrRbljd7OA3/P8e3fc2e+7UH0P7qFNmEOfzwI9lqRS3dtC
RajMunnMVSqqvLgkjJh8kH6QWyPVrlgxZMHPtGVkOzyqI3Q72dHbdlY4wNMKGmsc
lS9ZXJ08pELWkL9v2GGzBySP2NQLs7arhui5P9T5DSQ98MogEcB8m1/0fAuw2FWd
kpWWcxXdxv8vwrLizycge+zZnbtP5bywHT44JWZBn4AJklDghjjyy0n82zzdtfe7
bgu4Jb8o+UcwTTVtHzxedqi2QVgrMuvYQilsgQq00JSP/WaLmZ4xRFQcVRZqOl9E
hIHbP4RjvEKeAQoxfQ2Vcz7zSSoY9fZEfqkrkutbBt/9VMunaHxd63U2oV2OmyKp
82TD3eoF8vf6FrEPo12m9eZ08S+0nEJxJYdl9NzFGDrngzn9PfMAk3XVdMWxWFf0
UcNt71GrNA8SMpq98lJF4OrEFNn31h7x5LgD+aAy0lWCtTE6lDPNNcKxiXlDgnuD
W6xi7ZYcFI5E62XJ+kNfdV/TwX7WYCqkEqZ2AsnUuPLKoec/llGAaGGwBTZPMXdb
vuYbZU0loDQZiN5+eMJ9xxHw6GNzusjCioH/8Ryy1yLv6KIlEAN9vQ7QL7Akm/0o
pMV25pSRMC5Ipkz6fr88h53YOsVyhEGyo8iA5rCj1mS0v4+vkY/sAFyEy2JkDAfe
eAkMKzkMnTC4/vRURYmYP9sPPkoIsuP4O7VOw0JC1FjeXET55zjPMjniPq8zmoJ0
9QzpHn7hD69DnYauh+vM8A7IH/uVt7JIs5b2xM3jpXMh+g4tcpIzvPYFm6gAhxE6
K6lWsex4eJLG8TkxbQiLJnX55oZ+HnEsloqOWAd8TZWTZq0JBtI7Kwx1QSiHz8pn
FhMEeMHYcU8VtqMfxDH9VirV8/Tl7yn9Z0UL1fsemUFugkqUF1xV5bcZQpFzoaTG
0ClUdAy2dDg68bXNWsdPs+AUxoKDciiIEN8kWzh8WaG0JzkYDRP1Mj7+2NXDzYXA
TerMVtDkZLKObh9COkC3NIBoVD3NDUPc9rM1nkTMrlGGxlUeZHgB0hpdbKLnHUJJ
35gFipa9NyV3EsCBQG4L0VMZiLqKYah8DXLBpgVdLAMJuseEKw4qyqqjXLlMUIKy
l85+yJ4NM+jlDH14Obj2JfJ+utEAc2SbFLXouPliGoqYcXADmCDGV/VfX3CI4ufQ
RlNb6FXkTZAtLHV/m4V3LRFlKzGUi4Hw1WrVSD8sI0KaOOo15FhEsJwnAX98nQwQ
e3/7n1JUnd93QZlny+BUlboki+AN+9wrc7HPqHWtxbmBfBHGXibQBThZh7L1owO4
Cg/KZo/QRqYr8FB6u6n/nqux08lR2417dVOAulKnvmitLSVHqyEtyq9WKYjKH9l/
m7iw+8VwQaOB02GPTXinD4HffZH729lEDunqr3ZZ/3J4rQ70/G9ufPyC+RR2HJKH
+AfIaNCzwI9JsFE4VKYgqL9/k3YEUGZxH3IeiK16ejIaPs6Yr7I0HqGmyvSZnfOr
0gqKukLEw+jyWC3AMZ2hrKPDDZKXGAXJKAj+2fVS3bJBOJcHLOMxMipHo+GI6lGs
bbVZ0hY2J5OAxr61QErdj29oQx5KAlLd/t8EFe6f+pWa2vpHjIsh2OZOFq0r4gFj
HTwhNNAnQmbzMWmkUF9YYDY2+Jwa4qg8wWKlqtJo3fmHFGqOnpm7/uQx6KSMwSbu
tBBS4wdvX+YaeMZ48S6VhcgQJnaXifO4OXcUx+y8OLp/RDlxYVVpPdPJNDlTyCY2
MnVNzAdTuVusXLc7NkjN3EuRjc9GlnJShV0MlzZ412A/BCFAnCc5IlANWaFu3voC
bb7p9jowovKwFWa/wALybIWt0JmWEQxgcg97WGYHJjTtfJQt2AOtBXRF89PjKY94
p/eEFxdppIcfEzmoERHnjthLVEsWWzEbeO+zei+mkGX3N5e+IfjNF8xPqJpjZP57
/qFp2qAamWKrNExCU1Ci+Eb9TS+doHW+uhPwG6+iL/xlEX6GWDZD8q6ojvCHva59
kRLW9tTW6uEO6oqLX+dB8bWxTabOUgpmX1zSAtTI4C1GW23lzrbrExCzaDxgUIwF
CRLM0/JRheCZhxSMe56X/mAlXYVvkXPLxuvYhX6bKq8eD9We9KdzchNNKGmFUzBk
BBtSifKHKmsDPhA0SCHzyp/k1YtUaZHzZOV237QOC3KodhwG0tBvuD5+Qu5DTgZG
vOCnxpDTP/xXsx97PbFEXKwwUo/VK8I53Z9EwUukjBomr5uzfc7iAW/+ZMN5SHkX
VktKJNtt9RUJr65nsL9dqe3TEYzmVB1Oxp86SofARNYurTOFQ85qvhW0xxv+7dnz
ADl8io5S7HgbE4h8bi4Iv61WaJrpSTfH4ewsLDCOghtYLGs9XWlu+if96WSO9+lp
BnOeMx/NkZiM3SMER/S0t677Q3cktdqSmtZXASPA3ev2MDMtVW3lkLc2mQ03ziA5
gy7z7lEojdrNEh2qMcnK8Z2F/Q1gqjnlbaNrvrdksy5pCy+xoISGTxv4zKRMcfHS
nrzbdvmsrJTsTGCph/IT+nXydaV3zVI+AlcyPSaC/+9Vpkf3awoTlAdNjDkepoyU
WVpomBY+xt5Zjg0vzQ/rs1CFXssrkw7RXgN5SGnP2bXIrsMQas0Z9xO7jUiZrm2h
T8g+q4ORChCbkd1xNerxlXOb61kTFOqUoyilqxS+nTbFsnKbR1b9xL8C3xATgEHc
O9doX+kh14y5Qf+o0hoC6DiNUrdJrVgaZAr/eWlKjyryYgvvNrWgpfgyFoVlWDqI
kVqM5b4DurU1FbusloaJFPGL+81XSa5NpUlvDWhXTKqzqNKuDMJUgfULVcId0w9W
QEtvXe32IY/yEemF9Iko+7cTkY3aos+mL1HHVeGEHOfOp3oOq72lNWMxwRzpc50X
sqMdtt090H1jJ8HQNNpDDymqxELqGjOeZz73mGhW1fd15/JlKXtzWdasctGkYOlr
vCUPcRn0WJA/zTyCh5lxkQ+haGYlm6NrvA+mE1k1e67bn8926dWJZZFLW9QwKNIQ
KZRGSr/cI3zvZDoRA1WZo3Oi95m5UuSNnjn6+vZS38C15S6ZZwWLF+pGpznjsYvS
+TkUvfR/A3L07k4Shr22jxGbqVF+ou6o0M9Iz11GGvnKAt7J9E7lwy1fQ8ATAw9V
o9boPeYWmvgNSsYF7dr4/Jnyp08bLBVRDK723ta4gF9E6J/hqTpKLeJ//u2ZtIHx
dR41cMq7FS3Rh6YaEbiUOLVyOofhiQbU7N09kRZQkCB0W1n4Sb66vbdFPbeHf/y3
vOtxmdoEN6u2ZxIoXasB6bOBe3/06NPu5NPjbrzFLExXThWKxXECWj9EOrpjroAI
I7H9eyDguYiPe6N2DY069NWG5fBWVtfwnUbFBMGeFBIjuBXT7SW3BZftO6VrUpEV
hdArpR2e4jfMbAyvH7z1wsI16oh5J5aOA6UzMnCNu3pD03gndiQGR4UJ6DqTz/I7
b/tXAvfwudoP6Qe8LJtSM5FAynMycRchMLs1JHTLk+cvtsrcbCfGzTYOhwdawv6K
V6slAVof6Fg/ZjSdolHsd/44nUj2HQH8Hmc3QWv1+zkEJBNhhdRUs3lAm3CASFIo
1NFa9GRHPlplUIc/PzLHO2w8SksW64WNArf1cp3VGaL2O8rhGSxVQMfZ70XC0LQw
f2bEEO7rsAJ3jAJjW4SFSyjhiOwho/rflEsgEkX0mDzWBvxTZ9QlsYiRrilgMuek
AQ+PiMhjAFlJ1R9Qr7DfJkdQRAz/R9a8ujy3iQiUuFyN3o/EHKBfwicu8ZO1H5re
fVUkrFSIW0KafBFJAUnSknhoezKCmws8UiHPS4m+s7VSNE2IZmFbiYE24lleQK9Z
9PNMtrl49ePnzuEMm5aSngE01zVPIFYlFdJSjGY2nUi00zhU3wBqaeifGm+CLSx4
H7pPoKKZDb863T80TsBWHtI9ia1ApPRyngtkgnHHvkm71eTRevreA97y2w3MuyIN
/dLzaomXWHNOZZ5krmhS+Z6VAIIoGygLredKLNVOqJGW4Y1zwcHuIIp3RO0JrPBm
2uBPxtiPfuGVj8Lkhi5iv9t2p+O3d4wRzjSOfix1ZMSvO+NGl31NEAGaXy7lw8r6
taP6dCYoBEeHzHOGd49Dwt9G0hM7Nm/0Bqyd9gpi8Tce67GVDhiHImSVdg4lD7Y4
b5/KbZrBNMXsdDBk2UvSfdRi49R5D9iXSOweb1M6Pp52UrItv6KK7zU8NXaG2sLD
2jRy684fsDVfT/EXpc+Lz3YFPK+LNeF46RBmKRy4trBEuSzFpWJX15HquvUIwx0S
T+af9iVK9Z09DDY9uxz+xpi5LN2eirmOxF1wnOgWzlhMTwtVXPPNXg8oULSm+YU3
Wr0MXVhnSM1Gz3bJDcZ5kRkpJY7GKBaTBcPXj7WNlhnrArfqcyzJHm31+udjisPy
0xfl7VsayVD7G+vjpwJLkALtmxY37UWt2r9MJzquP03DBmMxL1gHzJe0F2n7zhKq
f3yNzLQpnUrp0qlVl8kAWRRUVV7i4hJJvCsdt2F0VG3+AQ6uSi2miDqWR6O+gti2
WNarwWcn7rdAJHyp+w1+R3qjSXMziDDFDrVxc3LPxBSJIQw8Eey3HLgklwutfuhp
rzRceNVgZ2YLXPnnwpM8u8Bbw4ly0UV/Xez5ushGYoNvu7wYOJcmRpa7CG4LZFqy
S8ko3PxVizWtfmUuYp8TPPtdzADTYXD2+S5pK04a5i1RZJ8Bp8vFIFhbOZuOLzTP
3gWGGghmrLnTUWLRbZurBD/iuvcmQqpKS8Aq6P4izeLpLyKyb6D9mXjXQQi6jmOp
6iSIpYwhs6HZK7KEwv3eHMGqzb6FAUrX2L3s91bBQnm33+GsCsqAhNnn3vN6+gvI
9+0Gbv0O78FFPA12hjfiMyMmoj42VjTyrcE5ksB01v7h+hcoLc1oaQ0RrekNE3Ev
vVud7BFKJ9xSPeyLQ4gfB3/ydTMxkbH1NgEMKhu2+A59NflSolgXNCKOGGrUDjt1
VRJ7k0SGoONa6J3qUpsbdvmpSv1kaAiw1jCiVTzLHgzg6TuBdW62hvcLPIYYe5Iy
UMUruAkt9fe1R5DdZ/DBafFFuOpIBBMFn6b2snaOFxLa+Y0NhcP1lxjJMokeS6Gp
/QAZ6gn6GPnxH6gRtlLt7QhpLBLaAJ77G3tvk+US9u3XQgLHf2f621F+9GVx4+XM
0Y1XIQymmhO6N71WNFQUcDlRqvOV7PZ/tigKegtz/NGMPmwbXkGLoIXpzwZ7azms
/jG0lYA7SHZraNOBS2Ut/xQk6pvxM6+lQrF62ADXfK00IP5oq6hQ/4Eu5UoCwv4+
lbfQ69hRcgXtwoXC930V6n5v03K/VujBNqbeaP9drZWgTWe4kvA9yIJQ6hjgtIZn
Uz5+o8Vi4652wrcSmxnlfuepUNprm2GTkweMmFlNO5pldSYgUjupZscb+o1os3wZ
lqkEFGSG7eIlKNKGD6iaDLDAl/aOHSzLMn9AUVvwDrQNiVrUomSlsfinwkqy4ixf
6qKHM+J8+BvYTwzxCyg+vv/CYZotBHoabuk8WpulNdBvjz57Vf9BHB16yEvu0HtK
fTKuEUvG/Vjk1FwCr3agtMuFE8wS3rAuSUtG2MFj2SRzZN8+1gRlEIP+R4zUY8BC
eurBORsJ+4lXYMUWSvuIITQhndyUZhPDVBTArhbZnR9HDokGa8Kh70E1+q3od5N2
v2givhXeSYUlKMJDJuNF/9xoDotLidwLo4B/Vc1+CdfyPH76AszcPBBqLFNtx1Fx
mqc7wkxUzBEY2SlS9Aj/Y+JNKaE4jRbPedrVMGBeRVCNcl4E29x66ZQV6mGarCrj
n5FRrJKpsBrcU+Lq+/sz6M4c5XSiS9DEwG5f+Q98fXLGbU6htCA84q5HbwZbRAoh
TG3tUA/d8aznvh2QFzPtHqijr9WQ5+gTcoTwMRpGfWYUHLjcNv6AHEI5h4swX/TM
iezOaUUfwomwZp9LscFy0SiGHie+lGwvGVTPCOPbxKk34QCJqpYtxDEvq4lQQdsC
tgy841V6Rn5Piu89BkZaZYm0bDHcgCDWloU7h4xVqK28CYtyhMcHRXh4aiPxmhp7
Ih6Y1DWVcQ/QwUj4PvwoOIBTBBo9H0BMt/a/9TQdmKXxH0xdQKav0kvn8TItfHvi
EtyrtMYlVWO3DXHTaiLnMoccKLkYsdcD4Kskq3zaDxhp/MkM2K6NMihl9BUfDUT7
B7pS4C6oKhPAMXebKWBfXH/cQg0sj294ENPmzd23w7J1j4LKz52SLuL9Zdg9gxfv
7fZSL44leSl4IBTD3vGhaavu+mz809aKG9RMZu9QK2KDf0tXPyNV9VH6QcL4Dije
otGb33Z0nB/T8F7hyRX8M2Ss8zxEjspowdAo/pyEYRcbpkqZ2wrN5gLKpZtQ5WNF
xcAy4xvIo3Q+lho/ylxEKLsV9w9WQDSJTN+j2EG8nw/TqVoZbmlvVbh4F2/SyZEL
z8+HtoVzw89IglDrXKP8r1qxQWUD2L/xx4iuhTluufm3Qr/GV7ptBgFZorZmF+C1
jF7ugqMcNNETtFUXsROCzrVDj+lsyo0Xg6HnjhkGGTKUjfkWA1yYJ0QUsF3D6N2N
BbyoL6XJrFCan/KWcQcT8TcS2ixiGdPLy28RDw/5LKq0WvnoSBJN4P6ZqnR1Kc57
bHBFQ+5Wvh3dQj8906yXNv6DXYvr0CwZUYiLU7A2XU6fRQTX3/nV9+/wrFotMArO
nOvJ7rwooxNB18Ki619Yw0nyBTbsEzsmGEPGhEwTk8cF+TEiOvPqb2Qak21asHoT
DjI0eUTIpxgzQM2GWM85yB1760bIWMCjgUvEvIzQSHLZCqAcKcwhrlM1JBH7ah8j
NpNdPr7BuChS3vJPfojQmJJTe/yYwt732fTV8ffJnFCbaDlGB6E+fzYXPu6PdxGD
89wrzM9JsDAl8csXN1CD8aakUr2GvvBxUx1rBlDDcOxFN+zTayNKt2CMsq1zX3kX
muocK8CxDbM7dRA1drStcksZ8T5aE18POJJ+lbk+yUwIXfFdq/wS4vveDFkhm3UN
FVYRKQK1vr+FHSvIahcQNwgXmXrPUeZQnFCLD+Uyb+qM22JvTe2FqRT61CdmZN3u
AwVHJqSTmBQ+ydZ4uMfwhe/WIATpY/FE0T53CqAEPq4BxsfpZpkdgBZaC7rjaiir
80LOD3KoMClVBWD/TUP0MNJ6uSTkET/0UmyLN0H66CZ/BC4x2Tj1tJR+bcEWmCN3
HtMtVyUXYmy8qxXC8MY7ljDMURoxxiPgSFguH5Wg0vbXfUXdvE6pngADM1Tw0RzR
xoIW76JWIloNUVA4yzEZYOt1giIbaOl8zpkmF2ZHogdYaK2qeHpW2NcG1kN7BpaR
bk/EY8hfn/nj6/99+an0bMgLmG5KTqKLR0LXZkfp+YfHY1/io8bVVRTtNlmXTdZH
XecZGdtcqVcR+7aYy6GGPaEsqyZ7n5/0PiM/MU3xDCT5/JGVMEbIYSAVfFzNO9yP
0avbKeNLErvA07KFMrPVCO0gv0uWuN86QHTJl7CZnUU+g1ftn1MZvmoN1hF6CLxl
1owj+Rz/QBa5YY+F/ph+fyF16s/8DSncft9lf5flyN8J88Qb6oO74KAxNXOn+U1S
CiZnvDg/ZCpuwDl1xMLR71szDY9AVZ+QGorZuGD7u1DReZ+FIswVrVle/YGEqSvF
XZgGdLodnHqFnoyWgLGL1r+aEtApukrZchlABYuRi+/iuLMveDu0u7fb+eJMQczp
mMq/rudX0yL5Z5VoT3IbG9PQ5jveEVw0JA6T07rUfm7jYA7pWgmJowO+d5S99Yiu
Ubx6CWBtZoHVyl8n1SELERXHXxRlXFTR4hoybv1cZSBbCV6i6BEKB9GlZcm478P0
MkzMPtFD4FUaZifqb75D6Q8zwoDJPswNvpZIrLhKlccoVUQwB8xblMXMkrmoAT4K
6+3kkMrLWKyn6QlicuIHmYAHIUvJ56mbuAve+oswJyo9Hf9j64ORmu8DFFX7JSzS
KBMi+I+DRHg29ED+kitm25l6POimvsjS0Z4zmfqYPEEA+rC8OO59NS7nulqzwPbn
N0IBJ87OQ8z70mOu8Qx2byQowxaxi9GXDAYeor5Ou2+7BbnLB/ETA2hWXJp5sl4G
JGqLtbr2evyoOptdbD+YX2i6HAHerzn/pA3xAC4DRbJ8a3iUSxFQyhRDFRRPKhqM
DNaQlRWP78QeFo5R+tgNG95bNLlIzWBYt49vFuRv/aH1nayn2QTa+oPiDdx0zBwA
o6596ikhczrT3BpVJpaJjrCwQvv7/JOJ0kSvLbgEeAVTR/aZHPzPD2c1qjv2/Bpa
wWuXae5KaZgU5DZDV6XjjyoRk62jYBPs5EUnLfJp9VzjVPb2Gk9ljEqvhgKCoK0o
bkmb8GTY0Q6+b0M1IU/mAf3gjI0LTR5repcQFCD6KUS3els0l7xwe4ipgwck3e/v
msTlT56aLRqwLcVk1P/5clpmihXTXXGDXAI/K1ycMLrXQupfDKA+QiXfSqqnIj7d
dGWQCyHLNO0N5BncBX/OzCRIDKGnUPqv0CT2gbHMvXtt8ZLAJ1B/B2DL7ehTRqB4
d+kXjZ+YgfJmCsOdgyOjrLg0Z71ilDh8okuKiSPG3HJJsSBHgajbfTHEyt5gg1mU
ZQo7AsC/co118MILmd8djz+BxIkp2j6k3ShWFVvqr9rZL8A+zGydwTZzMQ7fZ08K
l00amauUS9VPHByPiO5JuWbIhbAEy0dLykkphqG5a0echq/ntFeBD294c5GKh2vD
ZytjJ+BhQFhQCuIxQy2SCaYmE9uqyTxTUsCTPymfgcvj1bCXooz1rSw2/lEs2VXk
msYESZRMYlvNtN/rSf60VR3/1JZ//aqUKXAoRIXviZfTu1teMfRL0g4ufogl2I8A
QbJ33yap6nVv3ppm/vyUfEFkwX7npne+OvvL0KOxBvcJZ6vSdmKHbOFJjefL4/Nm
mNLanIHWbqWK3h6E6uQN6mIX9ro2ExA4oDr6KFSpuFeuyXPZXNgC+4PNQ+9Jry7n
mfRdydCp2mjY1kElG5CkGAAFMYaJgmeXkGuP5pZBMVNZhL7/vNwfnF/gXD1LgwaV
yZ8XSV0+6Sdjp2gEujKseMJhZ3kxxj+NwIYX392x8NOkroPbTbQvhbMgijOjSV0o
6xaK86mtv4AwhsrmDL9wJV9oNJqwEfMYRaKpkv/rJXDTgTDUjJePj5a4Mja8GPxA
hcunPx6JcAe/RdF2zn8tYXjoq7CPxus5s307aEcrtNBRtJ7dlJrhdmE/Ad6mERsG
Ix7ZnXBQLDQ5Wjhl7G1A9FiQ1+mASMlWxIRITbXcaGPV6i8mtBAxASfzI5o3pebL
UPoCOYI8KsN2U5zQ7KWvwub3gPHIgw9WTW1KEFORbOXROU9SUM+hqIZ3ljHyJHhG
wH7BCotgeDCGfyZFh3jL9nqMyYMK9eFOpmJmFSARB0LElvQqOf2RLv8LQDmzQPXg
3RhpGKRjcV76/IEfKs9lX1LXVJHeC4TZBFc1wnnBVN34F7FM6QH5nYdqnECOgLit
lRKVwuf42v1TFm9XkByzrxmZ6a1l5D8FR5vy83x/+vqHQACphaVlAns+bFLiZzOh
+KbjDywpBYxJAwkwnrZuMowaDI0s7S0+uJbEdeT+jAmKvIEfgHN7E6Wxky3RSloD
uiEvdRPMCekKU8GDMyoruWUX+S71nlAZUiZkLALgoI9Q756rtIfkbUDFq9EnXLIU
hnKJ1ehY/B4szaNZlVl8x4xTAvACNsc62zp8dQAsWMzY891OC5ct22sByrsxWqlN
WB3y1vam8NIqx8YIx+pUCctCWBEqh7gQtEompqFXN7Wo5ASvqqQvIvXr5eYJhbJy
NDsohSndirI9dPxRPo3Qtz9twnIf93sTIFLFy1Ag8IFYwC87+jM9dbIXT5+SkZ1e
/GKP5O7myftA07MY7+ncf0ZcxrsOxQhQl2TP5XftEZsOYNFlFHYWqqf9+sZxL4zT
5efFUZuGZu5XLwPrROSJvynYxNi3mcxoh1JaPl09mWQKx5RlV+IhysDQpoBY96CT
q2MFPCzGqjgrul5eLqTYXekHonWcTtntJmeDH4wGYU328p+el34OvMh0OzmlL2I9
86bqbVcw2+jqmSwewoSxdTf00kJ2EGkDqHyKjN3dGmMlJszYuOh/kwTOw7Q9asw7
ldv9oaGCWjBShIb81foRYBbeAqJKoBekqVKx/oZg+d+p8U3a8EeoN6aGuEAYjkVd
7GMNaZxOq3VXTFdXI1Mr57R/jklwZ8VPOvdGhdorfc2f2/sXCCpy8U2kAWZo9PZx
a/tqyM5D0egSYTfNSc3tlHeqVx4Eb7dr8res1WpbGUatMQSB5vwZQbYSqVuXQA0P
CVKRd05KQLIzIObFCOYMWdAsVy7+Wrm3M6Pz1NSVp8aF2XaX6u4R3m5ZYciZA3Wb
boNOzQt8rJ9lkEhmTJgtDg8GFl039bEF4k1wcF0B3E2IIOT/hvHH27mh+0S1SBMB
s00QB0EL3dpFVDPay9+KxRSul1JuhbNFjbTEGpbrK/HnmUBk9kORiwopWPo7luJs
xoNgTnjKE+XHsvRqYnZPDJIG/oUxFuhSCd7UKJZZ7FltctAv0nuXOOu6jKwwAPBn
HqoNTahC5BPOuGv8xLafrGhsoQL4hUNIePAJ0j2f+55CiV3iqyOwHg+ZYSO1VGFq
PbkgvbkQtnm02BSMYjh6+cQXfk4eTKWy/FFtR1udxNiBoNmS/iIiGF/5F/kryjdB
LRdfwoJ7bc39rBQFF3Gv/Wgzgdc5ZEg7crNnA0z5rjypslwNTvpb23L0pADQX7Ma
lxdKM3sS9cYvFDrvLRYtRbtWxShmX+uh8SwOVpyI0T9ovXFGQyhYdDpuJiB6HVW2
pvVM1DmajjxRf9bqSCq5fO7Dh//0WCXEpQ/yQ6F55tMSzKYDwgCbIjCxDBENEs9k
aMlV4ceriRrlk5/YZ4OJh4DvEQcWpFV2cmD/e1mkKLzouzu9kwwxJozVmaLz6R3R
ogeu0s8X4LoxdG5+r05rd0k3aR94X+lSXXTMTL0QReWxXMiyQcxsW+ilZVktn0Oz
VO3OOQElPrJkWTG7YHIlRVhMkEFxIMlL1En5BANJcY1OyQX4IW7RB5gbjwJtsO7b
s7gOwsr14IPnbLcJIfKF4Ua7apkRlMhmLI9RmLts34PLFnbJ9uH+Tyyg4a6Mj4DJ
See0UCm4nri2g22L1qvv6JTKWibEIDLIsMWVZTtPViFqjg9SLvqt7NLWtslZysdg
LQUmhuGhXaiakloVLj9a0IBE2DCnAFEDU0dlgvxVVRqWb03eMBSMG/pqktlzRaJm
sN/lsndi6u8fjvU5cuuzAge1ZI4IERxbUvrfn0vNjoBg5qREsK7cg+6LNjACpsi7
a+462JP+upyX6gDU91++fLis114W9jQnTr696VRuLX47/JS4zFncB5pCFfYSMP0R
fqMlfHOIG27tqgtQ0aV/dJbD6/tYftTWmASSTNb8AOlSKE3yr1hTXbpLtRhpmDAm
90v0orMdT2Zczd9uh7NUZtTqbUxHdTJQ/bciC2wNdml2aL1vGZIpid82m8aBF+93
u76kDVODMkIT5OompfNcXx21RYJp9zRqKvCITPeXJolFZHCse5WEzMDB06WCKGOm
komk2MS1RD3tXAzNKvKgShLPyb2EhytKWwZ003RclMJFJJ6F+HbrMZvJ3Bvy28Ov
aZ2vNMM3UIVvQBUFaKEpsT2GlNrRvk7EiIGluYu4a1lkgdLNnvjjDRWsDLu32O68
c7rHbA59tHYFFNegsmOmRlPtzun3Gm5KjOV98GZbNau8M1MQTtNBjJ+Boc+OnE8S
7uhH9MpmErsosTFxb/1DSvUw7xm4F4ZRgAN/GDfR/ou04oOSNF+cZS4pstYh970s
XuMX8/q0sDX1hPWd8TfCqcyktxIRiInpVnI5iCwWJbGkMDNLGG1Qyf+B8kUeWFfr
O2JetpD6POnv/WNHa0TJAH92CazCJZ+EIaqfvf87lQwpHonwWaSOiu10dNsnJhwJ
K5CmCnASThZut3nJVeuSjXdR82F/ivjYoj5EChiFhkiom8q5B1dOCoMHbaLVBjHc
fgRXzQUUNmjNtCgfp4TgnZVycODmygVs5LPBfhB1kA3Vw6H1TWRB4mAD11TBrZ0P
ElwMEkCFmStdUL0hF7C2kv3N2PIYNY7pxZrzLFDgfRyirYXaYcXauG3O/q6ZgB8S
LlBqon0Y7NWWT2E/hIuOgScQCbjfgBfFdnO2sqF6gk17kmFclpMWqbDZBYRa1X+5
nBh3VUZExgf4vxrphZAHRsKQ7P5JX6/OjCLGoyR17a+5mVedCkar0CUKtVRSTM1H
60dJ+OAnVyTMThimxccZllF3DU0JV4f7PTGy4ngKMtqoapJMyK2DnI5t4Ohz1C0F
I98ePbr9XTX2jePoMwzHqnPB2u9p+jafTPw7y2Pntrbi4wSwxefGY85VzlpeoM00
LNWyT+Qr0/3LZJITZITW1uOl28IWrziI9wXIS/RHJE21H2Fvd7oBj+iVok1+FVD7
3UlpDRMfiewNwoELhZ7TbJqIzRt6u2MGrihbhY6HbOQdQ24G06LdpesM0a3xXet8
v1agpKSCvc0m6zfbE0QMJjgpyrEYfeqi5fb1h42hQnaTLnZZc4nkaYb82p99Uh/F
YkndP4vuDcrJo9Dx8tbnW/0dHcF0i8JZPh4aAvtx/1SQ6MCA9zCNvkrI3Qx+ILhH
eu1nDGceRDE668URkGamxvRmvkGWyxcW4SCx63r1PYppOMMYjVgQOOjOQKh3HkCK
3bPDYqdeQotjlsCmnSdGETi6JGmp1x3hDpOuH21taaLyPSHLzzbUfnDaIzAw3T8a
s/I563K2xuHqpl8Mw8mzf7OpMkobXa9J4mKjn1kiLK0EfJKGlHAPch29tS4hn1yd
FbttKsYiKG3nj/YOFpvGjN+lZBAK8b3+kWHyOfnApZxze7/SvzmkP/eO+e95u0ta
Bs/7AAGI+lhB9xNdu1igjQvDiZUUcOE7hwWy4o/TBMMet+bLDop9OCdS7LoepMbD
+Ocs4I0sDmTH5uzkbNHUuFBtUyH+Dukrdqq+ZZkKY+tIT2eMVgbJRhyeiu8ifBuZ
8z7UoBqsz4R1L/XYckmyPyqyw4sHpthYQ54e1NAHyGyM7471NK7ny9R6tX9Uqork
BBQ6hgt+qeF5Ow7zvWG3axzy8j6qJR3zgJ8NHrPNol+DUK8cVIM101mVCUdCbX+q
yDN95adCVFMW/8+kXBtlr3FMTxtGLGBpixh06vwA+db+Mnj24y6iFYa071Y/OBzh
vmcRcOHcx5vGp7sfLccEsUZK2XrAlHxtY30Nvk5QdUx6bFC8LNPu6W9r7W6e1eBY
3/Hv0nGAKC/k91yEa5Enqyx0dltOAyzmkT4KZpOE7+CuCUOiYbyPAzFLoR6OjSN8
MMigpBreGFqL16KUx3/i8ZVn782AZORJ0ZuQmULfxINkM91iIeVh90xdLK+w0hMl
1NUh7jRgLXLY0orbLVNqq5lAzNJZ1ScH+Bd/BY+tBR7h4PkwbiYhuxtXw91htQQk
xCZ0sZfxJtrcQ/3N63jrEuhwc1n3xvpzEdJXu0V+rSSeAJAZCzcNLU9gZoBR7P0e
z+Ww/TZMVWuR3MJENysVLLRruKTdi0WZfcPNd9/GOQmCrBUymOGB1x5//AdVTHIi
jjQwUt9kfZ4Pvs8IDVs6oah7gDW03g99p6/0h1d4NO5XCGJICaRfgSJ4yHJLgOWa
8Vx2OMP/pz/XCITAEq7kYCg2NmCJ7yHwwlTG4FAWfIK/OYWoOIT1JMgoiX9s6nKZ
QbCtgeby5Du+FU18LXP+G8h1IOVmkVruh8xw2uCabNjEFcO0G4M4QSIGyTAz9fMR
AU+yuAfJ7PlbBs9qe5Qw5Ig/nINPyi0jYjPshnqe5twpkWsFU5wtIjhstsygpVX0
rYNSfY/f4N3NAzyoesC/tXo/LRQggCubT4rE103Ei544zLAfVbmO4SZ6EpR6+PcT
by0GrLIlLhuSxYOZToo29GfUyuAyXSgMi3hkJ9JpjwTfAIr9xiqQqn7SmTsX/IS3
xDt5MrvMceIiWfEiPx8eW7e4yegYh8cKbbfKYOtgclhBZFffiU4LdHhA4c69ejJj
uiysayj7W0kYcQDXMmKPP8Zi15AFY6PWfBtDKpkoLheZEXsAtRUfFHfbI21WLU/x
iGihmv3OtvAlqGpLxKnegkjkWmCk2Tgyk+Fdq5xv6UHtuEmoEY9LvHFywElr3m0q
tRPXN6/CWSOz32xXcA0jlf2yWG91ulYZu9ZQV3tFZN8vq/a5SKo+RNFrmEwF+pBj
/D5+D0aTWegGcXIpPunV04TLGRrA1cvjyxhRVJpirUnN/EJL0MQddFuQMc8py1LA
NQRkdNZzvn/POmMtJX6FgaMSkzrL/f1Yl1e8aVziiK8VY9V0jAPMmf2y/yXCyV0I
sYCsmt3VfPtNDAqZyjYFbPBqBUK7+4EQDY2kLX9wjJX1QHAXPn7FZxQjHCbPvmpH
8KGZ+GjUp100yQzhA2wfwf7f8p5Qc+zYHqqM1Eop8ISt+5/I4BcGRHBaNbYLHl71
vENx6GJeDITvmpBD6gHwgY/571CDJWJOQ8BpnfhrnPvo56bgYcUKLg+sYEphWk4Q
ix5YpsyeXelx2AMrX/c4dmkc0HOeaBcPYxcN6T/YjESxQZb0HZnZw1ynAlRWggsB
wjTOBjok8ey9MIzH0yT8sxfB8/8umklio6r5esrj2VAYUJ6Cn7+w8jocNNbDdMG+
GKVbh4lzY2giaT0r4zyJu23n8Y/YmXdRVcFsaUBDAOqRwXCZRqlPVpVhRwyiyO9F
TeFJc8TP0w8iMRE4t5tiNcjH5/tmz2jFfEd3xyli3NCZQkRHLhFwLoMBFU2uT606
fUMElCjIlOnuPVfftL9pym7tAO2wNEgj/HRugGaL0FLvaqTpfHNw7kgRGXB8bEEl
le8uNm+9DmV+M6Nx0xDls1lsuCY+PLAGm79H5UjBP+JNgcP0IrOPQRacZ11nX+n4
LVFioah3hjy6syEDTHHnaE/CVxUsYt3PTObRCceR7nEZWhkgW4TFaa9XUxmyhP72
YEyy9q93Ur6k+iZdn0cR5HBeZxcQFJnT9WXKmnyUbmjtxkSw0ZXulkUi1WJ3iR4l
LwgzqmA4G+p8U9vF/EhOi7HAXRZi0MlpUfbIFy10wBgNYV13gG1n/1PzQIcuPmeN
Uz54Q/7GzhSiCaicjrNNbEJqfO0pYi+wF1OraFoLE4xoFdOx5rZD6EIDKCyLE8jl
RB8r/hlSu9w3d2i4lLalCqC4bE/SiEPdtsFxeQ+sAa6rAB4/xhry4WhAcfRMFpoQ
7WPmI9P0LfGtF7OkaXNFv4xOiyLRG1QX9tJNHFZOc6IG3VR2xbzc2xFlpYDfz7f5
Xe1g8DLSSkILP2G+cPdQU3O4thIM8ijbTlPTUIUB5KIsdRWX6MX1KQ2fDp5aeyXt
rVvfQsROjQvii8yupbRmBjSabtgxuCF14ObRrzsMm2RNLOOBRWhWoZDfRuOcApSO
LFt+2lnKPXk5xyqYP6W9Jz1YjXQEWVucsv9xaYX1kwF/IJHa2DD+8ZBrhnTAtkWn
CcE+Hic9HRT6Fm/Inooqwh9YF/U7g7ImTRI6itPlY/vRzXFlUwbRv4pqtm1hgUJc
UQLJclwKP7TthCx3Dxp81ZWPhkQXxPQf+mdCaWP4TjMkwpIkBuQ8xic8axzhLW4S
Ox+gIbdAeclnIZuW/0ufc93f8tj21J+Gf+1Hd5bxiQscZ1YohOlfx3Q1LS2laLT7
D5CXHdiwYUNfJc1gdm1qPvUTJBzx7YKsaHqEU/OcY39vqzHe9mjAzxRyluFqPJwP
L3RLHP6YSeIMclfXlmwN9EhIxS9L/6jhgH6Rg8VQ35a2vx6EJeOMODd7rbq+nVtR
lFQHjP0zJxiZg2ElKIoBiz0mzhimRSPZB6DT9z1FlfDNc//8skTyM/hjPK8Cv4qI
EOhmNejD78vmZMN0qK+3n/8DQfbVJ35ac3VLY1IvpZ1K83oEXTW6WNFi548G/Kh2
Ttb+vZShPUJuCUNILT5iiavQJZ+9GgZuQxGFKVYiiQ1bJsTp/LuktXwZDH9aThZw
d1S+rxJcyOoUNPzeA+AyofNgiIaVbN1tn9390CMQ38N23szs98zExegSsB9GW646
/X2K/TKe165lHANNrRmcwqMw4W23PCGOzstHSnNqNS5Zpqjjd8FCOSF0+7e3Uue+
fGl7Z2wc7pc9LkHFX9BRATn/rPNDLOiK8YqtbeJj+TnDDLSC+jYnNAGlBMKbjeQI
omJ6wX8xVS/Siz5Zc2mB1E6t/7NrUhrMP3SNISBoA53bbHGokhA0ifSuFTYxJlQO
TN4sxBoKwQa7Ge4YuE8tOK5bmjQJf7+vZkZbuGD6IOiDGKrn6RGI+0Eh0JV28SmN
DaKxMQ0y9e8+AeOkjWwqiHD5z/ktJxYNmcTZSQXgd1K6+dY7YtMdYSy/vfcT2csB
3DpFe1wPrn2rr2F6vl75mMUD8iovGrZ8ckbbIa461Z9+f6LsZLVnKw0lRh4gSczw
ebP7SZUyyyxYdtU0AEMXZOe4ApCbRAG9+67oiK30txQFEczJxschgnr5np9JGBqC
/7XjamUquieIErx2wxMH7b0L9Pb+beDY3jUzQBLrDO+U/0BxLNWs9Hd3xUNCY28S
WM3VHO8N7PeJAlleKDHimln5xzBC+ayq5yZWVWndnshjNqXHE0/jghPEp58Mxkmy
zcyaOFkSp7aMp+NeVf8q4Y2glA8VryFBMCDMBklZcVIfqdVuM8vpHxrdFmWYCv05
YJMeM3Hb6JteoCauDvbWGQgQ7HDwLR5ucm6MjmikZurRy0X/npBPGu9rdy1EWfLt
401syT7/dDScktIWxHQkuEsOrfGUQFXfm1IATb9+CKa0pwuExG2QKFjid5LnHXR1
SqR6MdhvtDQ9o9L+WiNIyuTujQXVQLmPeQpvyNItdhrQRs2JXYpOhODwhUBifEYj
fNrlp7x8draIcb20h4/C6HUTrxRaAdSNEFC7/RngP8ms2XMicfBZioFV1+j/s1H2
DCrQaktaJpnj6c4rZyxYpK1+RQTCTRq9fNw4xIQo/L1sU4uDn9XtLjI5ALF0HyMd
mrHja+AbJurR1iK1IRawis+Yk79XLzmwfEo4c6eOXFq+lKDkbStx+InpVfOV8M5n
fvLhHkm52P7VbhaMM4T+EM4+L8GYA+Z7MMop6RCkcIGhbwQ5br53h6EpycN7Aysx
Dl3e2fuGGuLlgSvWvouJUOFTKRq6UF4JmXakGKH3CsLrTwhMbuBTdNWOTR3DSDFW
4F8PjR+3vaQmkMbjn3yvuQX+LbjusliktTfQ9dib7rSlrjRuWDJKqltMkdk8y6lf
T4OFChHiLD4pqBzRz1Ovihk4dQgkxc4wvylKoxgT67/RAPZZ0siZbY788agSLz5O
F8o00G6EBxSfvaN1Dy5Ho7zQ0pyY14LJJz8bTevFci7EfLDZ6ISnAoyM+4GvFH0g
UfiZfiHyEP71YwKjvJ08K3TTggo4o0UmQ51qFstF6dGKhhjFGhkG+hF+joRu4qRb
974/vlfmWx/p5pmCmAiKNSz+J2eT0PReB6RUYGQcYb8boB+r3fOhjSN28Knsgcez
HcKNV4OpNppVvU7Epm0Qlsn3c6BW6VWOaWdZV8Yrh48KbZTbEskimA+i2zz2kgIl
4ykiBjFjQzH6SdDgBkRH0dqcv8NF1r6Hllcbv9cy09gkWR6pnLFud4fA+M6hgzbv
Zxxl1eWuo8uZ/Nn8A4URDfWEeh0mqB3DdIDibX1pEKCIvsgZ6/1tS/AggGG0WpBT
ej+trqG6nzsKn/OkAlBggDMNar0Tp28XP5lbvSMsUgaMUwjwqzHvDZdxzyAuBTti
beWt92gbmqWqkQGFjmNSAIzIb9TqdM5yn1TNmz+Hio1zaodq62x6EEWC26z2xDlI
q2jShW+NWKwJiNd3DDyiodD4agA5nk2VLSM6/IwyRY0sRJPsIvg5U4LdubS/a2nc
IMI+H9yXQeK6DwS1ZiObzvY4WEiD4T2ynDnVlWtBLFPvHFtG3MinGWxNYTW98oOn
h5TC6tsFsdLnxLcpkkrM3cOqy+1K+Cj5ebWmlXOV1BUjQlP/YKakcuTEkZgnPbyk
MxBiKMFYYe338Ancxc+Xd7Vx+mcah8/s5Z/VRXYG3nfl1d2eHrtOVkX+v8+kEGVb
lkWXhm8BfzcT5Hvf+KvlNv9SYqWJKWd0stnk2BFujoBNcBJxo+hYLo1miBj9zg1I
YHZkaDCGlwrC9WSRMEkACj8y1C0GxMX7pwbWitoOB73yIGalcEkxuIiDoy6bHSsF
3wg/ZWh+LHFDOtYna02r7DLbUMTHxjedYkizk84heMidMRKfJ3X2OnH0CGfc5mMI
9Qdwnhkh0AKe/guJQHDxitFNXfosLorPms7An3cOVJfz8CzxkCkcz3Xm7a3xb6if
K76FgctmyzcZkzL3BV865PEGQ1DCKodbt0RzOlinpmgmWts+wP+YjMSEDt1C3qdi
AOezzqBcF8QXmdQlqGPycGwxdwghEyufGkqSblcjNxRWl/mDyT/gI3+4GH/KqOx8
5lYJABDqhbhS44jsoPKUJDMLZb2Anm7N2QfP4haD6CGk1yN0loajlI2wIYicTwxg
n4x419EY/C+bhvOB/v+EiTakVARNKfX2ijgPyQ+Eajb9Q5Eekh9EfaDKOehvMv/v
EKed7TqWxu/ZGfrLPpDJ9GcWRII8xX3Yxko1JCJluYcmO4CwqkQMgM57nAtYBXxi
nv0sbFGfBnNi730EqR+LAeBa0eiHkeG7ZH7V2ZR+lrP0GflRTTnpORT3suTFic6G
H5TcwGhB92+jOG8uhzo4NqoGITI7EvyROJxJee47cq0fA9yGptZd29xJ2YwbDYfX
9WsQSb5s8AL0sbUNqFrjp7rptdVLzoDuuL9VIi8XZ5H1miqqqY50lTw6YxtTE4DO
1vAfSDDu6cbirN2fNb6g5RQ3YrjiMSzpvuhmOefsDKRHT+ludZnI0g/iPkJ7WucF
crRlkspnzui5TZlNNSMDeSOfIh+XTOyLhA0qyez8AAwe5DhGbvEi1p85f2BsY/7y
U6YDALcYE7uYB+Vddzea7ixvlTHk0IQy/rPqiPVXsLTUsy/glg5Z3kFT4Rlj6L1l
oUp3a4CH/uTRtvqoe4OjeW7h2oj2YnUee2wTetLcqEnJjI/YL1ktdUJD6hAO82x8
abmeM5aONzIgluvcHCc31+f2ployzR7wzokpJjN1FSGxTyzg8PMaZ+bABrnRgDIb
1LHSjDBhalU7inqiWyVlJ1QzltF/vykOjxirki26B1KdStIcS5xdPYb0H7xCe3Rw
VWZDWqqZfZdp/e6r0un0bDfBVd0rv9MjSobxJ62gxs9NlBjetslS7rRjfj5fCEhc
8NrYH31nxOduVtZcPcaGNnCiK1WJdBnwDxs6+jlajunWEX0w8MypTQyV8qm2nP38
UZ2BKvrRKbto+bVB5JdbpvyMu3cnfLIMt+Sn+6OpcnZd2E/WczqpRrpPY2l5T8D4
VDOE7Nakjy6fOwU0qqU0fF1JQHUrLpriG/KqS+fFJdz5kylWEO0jZ213m4vwzHzg
oYxSslhOt6o5+yMPYU7ylIRj2T7DfekoBQPXl7xeVZCkfRsuahbk978EswcxOQQs
SC66qfgEVHXw/58qR/3xthehgRUDv1QwOSCIu4XVMZy/17hDPdLD5SSOOrK3cHZu
sT2VLL6jLwxSeSZv6anPAmzzYAbRBhtge4UCS0iTR/s21f6SAXL99545glyGvH0/
gCvq7riEoUpLp93M2bGuoI6/e9O/o1DRpExH9jun5zu81pMhmTB4KBZDBgQ6Ws5W
ubjYrJU4hzQd53R74pU+frdInECw07XEo34resQo/lZs78h1V22Ov+MKcrIHOZvW
WZckjJ5v+zVNjycVQFGmiUUCMeWiVR8Z9/kxqGvcV2Qot+euu4ufn0xCrYwJ00eN
KjueJcNNuBww8IXPxkhkMc4lp1NrgdJhdpPWFhineyP75yl9jf0AwMRfqwNo+xN8
IgJsSOtE23blKFrs3G6MyTxdV14Hre6bBUFLphnFvymqJC/Fuk1rcO7KZow35csv
zRHeM7UAuWhlzQcJLAh5WRmDsZ7pOP/wdvzRAOzucxPj8s8LPxOYaxIyifRZX7Qy
PA1c3lTGuC17XK0kE/5jsGJ32hI9osAWF3U28w5uapmb9+sUeGceP2oedSH+voQl
M/bZXpW2eTttytPuQl0Nr3VQG5dm5UPxpwYGZTFWj6JarSwKKY+swl1ddReDp1Ev
IjvuXeMNGnNv36dXsm9blGgYNuCaJcOIBIMlknxDFie+ePs5e/BWaafz2xZt47Zt
LZ/bAIWGDTlQgVJXVvxaOJTpYi12WJ1SQPAmVUzdp8LN9agwL2EoUaU5kOv5cvnf
iRTIHsg/NgHisckhlK1HdLkjRRPozXEbMzfVekgzE1JBVwl3gzsdJAl3pKiwQjg3
BDkjpVBmeMoZ8RIiWVuU7K5B+QkQOVG9fqDwxRFoeCB93fZu9FrO6PiuyC/FCH+b
0bzte2npyFyeng0VvMeycQmnsZVGtHYhNwFZ38iSo8+l0JRjlB08FJ5J9gc42mA5
W/6sAfKWbzQrddxVy5oBm3dS8qXBXOG+TytU/CoB6XxoUUce0iGdwVi7a3IUXXLb
g0A1DP1pvwplc+CVkPWUdpGAH6Dlts+o/MN5q0aiS3RyFqayOuPzaa8HSrlfhZOa
+cCpp37xkRep6Lnd5I8uVYRBDp6p8LJHBDwG4dNn/AKSVWlbQm+c5XpKg1TBV7tV
xWp7xTX2lYNj6cnuR7stYWSlliwxzty0oWAWnHdESzhZjG/KmAD0Zd8s3P322LZE
Es43teDX2MJUN6IEhl7yuAuYiMLVypfWGjEaagKdqXoj4GBDvKVM2zOAd9OBjFgi
Dq38XmfTBI8I3fhqRQwCnNQRKLg+Tcu7DOujUlISUvIXm205iqSMYGSMH20rOMhZ
r1irgeGTXAd34Au4epv1uweAKF+vYkE6OxsLe7LeEsBuewQefbqtJPhxWL0rMxvX
lyMxYmnXstfDZv6hin1jMDF8SF/17XKENezHOJIpD0asqDPeIbuoYMKHF/yoQewz
bh0ROyTz24LYAR87L9u8/L8FeZk0CXOk85dfoFRVO3yCDlM5rfiOpo0mB1ffw+ti
RRxLXUJnGRC60Nds83fcz0r0+HfUD0GiZiGZNzKqml09HWj35FsNSzbImbscS/d5
45JRo2NGpsy4vm/CXH1Z6d5ehDleHiUgQB6voG3RXkNiMoDHXuXaBytyLViHDV77
lO9/QxmCi8Vv0eJdyu0OIaPaQvrz87+HVlI6FddvK2EaswYX3F/r9el09h9iGgDL
xCgNGbgKMKVkPOfRgcbebOkuabMnbHsuXgX1vj2URI2gMvOzh6nCybHTn+JuSwDj
alYL8GoFyM2DCKwu/T8gJjQNH5yjQRKceMjSKvNP6TyteWvySanjTiSUrbpfpom8
lL9f/mQBap0Vc9O+7NUiYSIuJbkJ4eG9kUqXJJjnAEi1zz794ccZ3U1KkOs2GbOo
yUmEx9auNbqBTKtWlhndLhzQDlEiAmkr+Wun7Cq7+v7FwW3kLCbpeTigeem9+a8e
1XhpRbcE+PJFg6a+hUwDeXSmP3GhwRRrpxujZznKjnGZJeRSwhrEryN8jF6wvlgE
y+L1xxGPI8Zn+Fmj29PvqAC8YExvC2CEyb0uj28gSASmIrIgh0iP2XQ414eg9d5j
i4d37wisj4wBoeWxwgZyMwV0xx0Qs8o04W+Ndczqf4xR/vpLUQzlTky1wuQtmBSw
BVsAhrdndY4tJb/aQ+czledGN55QF+Eytwf8oKrfiP8tKVyeXb8zlbhpOuCsmyo7
DIZLsw8FGFxarrrKRp0SFpJcdZEB7EcHWakGt8daCgDHGbnJcfUg76r7qKMjsv0U
FCOyDOx3FEXe9i1U2DGKMaX8ENoiwCSAOTljT4l39VgO8CFuwMo6T7AhKmPqti9p
DtKCcLXLpg2RCCiPF+CN/Nju2dfmp7heDMeQ0XE39RPqMXZi/NQzY+E8W+XtKoSJ
9K5SbON72h1/AX7fQjuOWyM3Z8AP8nmYKCZ2MUIZ7hCKl2DoPiab5i/GyvL3CHwl
22IC/NTTYA4KkVwD8z0/j3cl7fLaS/zOj8LYmI0Q58UmC3TRuxUqVHbga0X2L5A+
NEAstEZkoRsRce5nx4e7xkVZARd+Wdu0cBjItxI7xhpt3f3APX6yDFXhcjuC3gEE
Sk8U2oKveN2UtFpvn4A+TQeTnAf+7oGA/cU0+AWg8TQRU0wSJt1hrcA1tw5XBQFD
lMxn6qHN+EKm9R59O3BbxiS6OLqcxV10p6HVC/SoOb7NeqHh9HFaxVConsJ3alel
960S16gQ+JxiO2eutW2hVT1FoRRjjGLeJ6pTOyaUjYD9fImMmyqxZ6ZP7BA0lq8V
7XzlqevQ+sLfKKCC3Bu5lBv2dvM41JDnc2pEVCG48pYhHCNe25T8VnD6DxaFYfgs
Vc5kh3bHmtYFreipLvlSNPgBobt6knMdxE1WR9FtmP16RaElQI2g9E2KhCaQDJ82
ms7tkqiGStlaYvPLKvAsWbc4iOgZJ4n7KVrhZTvsk0YfGCg14JdsflIIb9QI8Dn9
9h1okPog0OFUq4Z9IQVlr6K8Qqx7SBudL0N2S809RDEpslvynnAuJ7dUOfULqH3e
na/r+Cwb1nGUzKrU/Kw8to9YafJysZ+ELZ7bJYhY7rqA38sCUNai/xGlLHcrDq+b
+MtdR479eQzq6+sAiYq3TB+SEvn5E7ahUkmJoNpSlBFgFVJT8gId0mJhfHtE1u8w
7DaJ/VJunrZ02eCNT8MhSSvU8blh8JwFQ16/UeBSqwqnSwkyFc/+RM1yw+ETR96a
kBzpYvsJpP+aI5kIfhQGCa0ks0Cj3Z1/zc2VBnlkBSldw7FXG76pM9sIf43bYv5e
XZcWv3bkN5Zz6evMS6ln6UC8kRIfwESgduHo3HTviffKfV3Qu8TY+DhGYCFFsbRh
hJvv6vB8qskhuFVETr/LdMZNhxeH/E5nlF5Ox9KwC5mkoORX2zJqVfel9ZpahVI9
d5B080EUmbir4a7z2n1GwFRu39YOLiFP+OYOcsl4yEEawFPdaYfAcsm+gb3lMlaA
8q05A2NAugxulqS093FsdknlKHfrixH0zvUh7QRJRHSNjuJpjDDJGCCub0FoTO8T
o34gQe/O/NNpmELqtosRcULLRXI1EtqZY5RgATubKbknJWZ10sBqmDqNoVYfSV6o
QdUMSWOuX90hDayw8oRL3PMoOuBqob0HbfOLQAXpgH6L1+ovBeiVcUhzUYMj4OIg
Qr1TmrJFBxe0/BpzPND80PU6cZhnb6BgByDr38xhGE+YN7Klc9ua1Jp12qw+RoC7
RWALQgVH8hNmTPqiWceaY/Xs6tyY1gzgMepKD9QfdrvY24Gh6wgcpy8V6q/g6kNK
D7ra/B9qxH4I18r+mcdiO8ryG9/Ct7qZWWNQL//aQEaJlhyl5R1fRipkgtVPfZgD
zF0Wc43DDhbv6z5lJs+qDLrkD2UDwn5xQUYgVK7hzt1VlWQVHn3+WEoPSRNEig+C
6OPs1DVqAmNKR0g0wPGvYOiWpVx8Ki525mbOZ4VnyRbDxTnW6SlUSsaeQN5m9FSc
xdvMfALGSnmg3xFylOv+C2KWacd6L+/ibJvcn8IhSyEqNOAmZz4rH0+8pKCgRQr0
6cB8oRLgksIf+bCzVu5cFMdr63zgXdSJZf+1Gc5r1QlscdY2ux6AjqFMIjffx0AF
eTqKIbqZ+lE3nEgGxdkiHevQqF8tdvZtSpoi+TTm+CfaYrusGIiHNjCiFo48jKU9
Mlb6zY8lfrJP6MoY+6qVvserCjda8bmXgVaL74muYev9aKS5P7cy8j83OLs+1vX2
12w0jtPAXbDvZ1YVuvkXSTNrWjXz2wapO+UBiOuu9X0LBD3UqeE2940NERl9ajSC
iIRXP6htoU50WK3+Irsy8RJtscWKu6ArOzliAI+OriK2NSItZzYxbFr9nd7JllHx
R3tTIKWwLoBooJnvotgyt5W7RufG2GavjNMb4KJRFS9YARK7xqS1J+a6a7Prm53A
J69vommpWAiqxwJEVZT0FNhT29eQCgIilHHyTIwT8noXUDR1XLePZJunDxPCIO7W
xX2KRlTeoHDL2t2Qux8CWMVB2L484+WHX05pY0LzDE3pz5cNbbSVQVQOGGNszFXv
lr6M6MTfptPPESk4OSzQPE2TcFOYYRMbCVNCNdXQ8EWQFzEEMHTu05UlFlAclELR
XB+kgH1hVFJe8l2m2EpNZJlJaYB1C8qwMhVXrxLmmXfKusfAGiOB7ZsLRb13XX+h
x0DokHdASgoa9nRv6zjZ4IlRQqTKmTADuHTPWqJVOrTaTAfdugGOwIMBCewsM+dz
6NhAZR9UnpGNekjs5e0QvJryjdI3Z8Nk9YxL5JAo7ybbPChfDt++kC17b0vsQi7L
ultBTGZosG/86UxW8fay6VIiogAVoyH2vbg2gczS7NTRXqpUrkHkcg/yXyDBRQE/
iBsZ9pvIVP5Ndm64sWt+Mk1HfuRSxj6LmhWiRLIk8UAORUmMU4sAEyiNiandN2Y3
RV6XMIMUNnhb0SP3ZXV2leH0yzOxhjRmKkMwBOl/rgS+Ya6R8QFLP2VkmNbJbpSv
kM2szdst8N8N4FQvJ2Tps1rf9tPxK+AtSweBITBMs+YYow73E4b+tVJ8PSN/VbNN
WBDcN9BPw6Abcrp8ePFLECxr2zXw1cu5yYOIeOeKe7HbAafyTCAP2yIn2nBxfj6p
hTBHJ76KGJksvTgo3+/yQOxnbk6f2Rqrc169xY+ej+5iuNV5uR9th0N1dzS/2Fxo
DZXIIV5y4Zlbu1ZGN0yWi+m+xo/+9kmE3YFEN5fEq/k6Mkpqt869YQrJ1TVxxxgs
RjotjtbP8+xb/QXCN23+Q19eaC+JsidLt9J4gI6gJDG/1P/bstVNcswpJp0LWmB4
sN8DpNDjb9ktazpLB6iNuuCSrdBLhabnbdWnri3ZDhuBr1rDzcStRSJTvEwxmGfi
ZD2fGMDvpwO2YybpN0i4lpGb7sNWQN/DqgB15VS+9JImIgEMUX+Y21KzUO7i8YuH
Yoxyh6uettnLI41DX1ttgqinAgtiP/K/+tzZibU9hJuuDeelObH/99/BdsB7eeNx
YLNg+5rUwLN4nWXvAP8niMMpywWI1F6kla6SdqrczFg9Yvv/8m6j8Ijd5JApBnJL
alUkKTXz2ogRQD6YXdbRef8bjgXH2iS8DDHEwoIH0I6fQKsLe013ZP2t71ig2goX
RDeNeNuoNQGIIm2UzQKjPzDGlGJoZLiNqo3qA6mlTdkSgXyHxc+RI6iM/ifU/2VD
/t9BK3mBqoipHhWnQh94X/EhPHA/ZK/raI+skN25CsufXQhAJGpwHkpU1UgVdYi3
QRfikb572/4uORUka43TWxokv/Phn0wQy2bgTJxyy5erEqOyhM3DHTe1YsWyeYUH
W+TPirlV6SaWuHXPPNIAbYOA/ec8L63dBnFMiQFWRTarBRet/M+x052Y/+S+8ZYK
uG12l4/O44uiopZDDJ4aHKyJDnjDlztEx7IvzZsOjJsUepWlZ7tfQNHawQ8HCsmp
k7oMK7VdVGelBT1XfmQEvVQ8CHpS4ARZEm1DCsmhkfCPyx7WB+vmRbk3v5OeCbwb
7EZuPG2yfSeuHT/q/lmjDCR6ah6s4a3mQ9xFFH33nJcJ+eDXOt7wRzy6Snj7O/kN
Qt8kGz9i39PyClgLOjLwDlntHBlbRH5zQUwdwRuslwcDrnegDosppLGRpwqLU3yb
lWbXrYaIAgPHLUbSxMbFgyjWRU/PS6UQghU+UgtpZxmW/pOUVIYPEdwo3yFJnLb3
zF6tAo7Bf9NlFUNtdB7hDNnhOOhSxLnM+Cs1xjHWkav697XVJWOXx80z4cC4DKwX
8jKaXdHEX7HbW2AJ8RC9bbWP+igCQ4z74E3YZmOvQfL7iNd6RLuxuwgcRfn9n6iA
TBy0JEU+aHYxXIFZQsWO1vC68n/Vk07opW6SqdayTTsdTlV3sGaIGvMCQZQqn4Gp
RcreJfXlHIUayKujjS5Lzi4PjIkBHHhyg8QYc4P7Co2PV6DuQX2M70MlVkfqfX7h
XDCNeKzGCk6BlO02E33FuXtcdbl4FupDtWZS6vbJrCd+Vkg/Tc3IVLVAinqxPTHH
thVvgtLJGUTqKszD11yPKu2gbE1wfCG3GUezVT9qSH5+BoD5weHIlLfzXaRCOEPB
ZsiQjGYKwswSaZ9WKuSTgpVbelUiVLlG7g6lSsEyN4HqsaRMcFKMIlzp3N9660Ow
jmxkGXbmLDvSDp600NPVtBR+SQ1+OoQrVL68wqIqKpWEFS6+Ehxjj48bf2x8y2Cp
TFn6bfdqrLwPyVEWWl1iKXSJEuHNe8foSkxwsEfq4mo9GB4f/zE+miy5Ad2WLrf2
9AsdZubiWfaLl0XcgS/oThPd4O52a6QkjclhkHv3hpLjxk3aswUq9+PYyXrfHvYP
mniAVuPyhf/iGgKdWgcL0YAOedEgtSqh93kDoHNGiM9AAHwSyLvTG1J2chZslDNO
gueImNzwLEYjIK5CXt5CROn7tr2wy5YnVfLdYfl3gURo+c6bs5P41bPSlmWj98SU
ias2MH1BAZaoHOOpdfl1/CxcuAcZVVgv49O5N7IUUjIn9N0Ttw+SRs9Jb2XS8X+m
18QXzUQQFP6vKGl+yZeuJ0et8vPGzgKjamFC2NzqkIeRRzNT8jYf+f+20YPZAz82
TCLYWEFZ65eRgURiVjGn4dibJpyEuSsiysgAdJ3db66+Rjqei0TgyXEIgw0V0Be8
+s+OUEmIKlAq1tn28I3pNrUeZ9G1QkKWZH028CAe3Lcp5ng7hRGe6n9JwYQ9omL0
uGCweAUX/L0+R6qCJykfKLW7mnWrfv6tdmFEFzDNDkxjL2RdSH9IWOk0IwTXixuI
2h+dmZvWuV2zhyvJDoXDkWgNLrhroKrV67Dp8wEvW7ChyFXz53ypsNtubIk46LvA
U0KKopuZmaaXvB6eFHmscU0JnIf1Z3F3G4+OfMbIImxJdVlgJuZuztzspgSGUqe6
D3532NgyFe5cu0mg78gBoxNRNVPuQiuGzB//6Vdcd/LgrWRt5Yrp4TjWxAl6/Q6p
+sKza6T12t1SMAJrIjgtDwK3RgbNxLwXE8agVgtp3cKxksCqrWMlILzCChcxh3/Z
fPCzbdaR+q2+v8JawYfOSZrSMQmGYLrNWIt8xsCv5GzqUyiSoBw0libdGKHF3sYs
EEeh9Zoih3a20cjQ+46V//9mOpM6iatm246sidZyUCwmCUVSUB3U3EAjQflZk9aK
Ultwk/W60TzsdmUIbkAxlTl7NVXIDXdBmxbjLDyUw/FM6zihYgcVJrnKtZGIC46x
LbzDgvV/WQ/ppRdRFdlgxJNsVrtJFhFI7YyB2poIAjYZPM1g7r7J1GZaTHaFBlpu
G9yPoHpXvBhk11itGVj/6rPgEPmri7sXWDO82RV7uWUCIDCIPdMHcFEzBGwbzEEF
yRJuuEo4eC3Zg4CZ4yDMfUZaW74yl4UWYzxN+E1GdGtc8T03Z58CrG7ONcuwZAQr
IgORXqaHqQ4Pk7w2b4oOkG6a6d6KOnw/+SqDp2UDdTAWhEStMvuALObWx7ZNCGRa
yQNRRHoaEVnqSEux44ER1IYRQ8m6kj6ZrGrCDufPsv8LkFiXyVi2DqX/O/XVanFg
vfdByWvc9hLTDRBA6wwe2K/H4pjJ/ieULgM4motP8G8FFcrqc91861EJimfz4pDv
sJwGlteagt9452I7EZHfUkpMEF2cvklixT35yElGs27kwuTGImXpau5Ru4vCDw+D
Sy/l3HRtLVBANmoH/lHV/fDyaq2kSxR6kBl7njc2yKDh59/NRxONpkSropWTzL+m
NdW90+W4r1+TcyphxyJfgrPNBN3NFwd7ejpAAnVA3zXODX0Nx0J/DeJBjXo+os+F
e1IASIQBOo7Bmu4dMy1PLaKezxeH7HFF3y4QRtepF/dDB1AbEyoLwmOg6KpeA9a9
dHadZeWHqmBFhN5yXG7d1vIPCnhhns7sFUmBKOQNUO8wqRNkPygLXgUJ/SndFkTM
fFKKP9jQP3uX06AMuHYCLUL3bKvo0323JhQmu5wuqvz2yzRHs5ZCU6vV4WLpOXOU
UJj+AK1lS2JfY/Va4I03QrsY2/VcC+S96O1mPYQq8K0h/PI06OzO2nX0CcGx5lZp
01NUItIoy6aqOZa9yFLCp9wVnFi2ISapZ2KxGyonIfxgf1aN2wFwAmoemQoTgtI5
XJVT8suLLFvWW8X0lxAaS6+W19ZJMHF+yksldfpHfI6nLG0UoGDVxw6Y9l7I2fZO
Td9ydLWLDLj/ECyhQviuB7ylzboOhQzTWNSg/sFZUvV7x47nz5y/mbWeGGj4wIwl
aifkdi9UF2G1c4dE34n01XfKXtSyaqTK5AARs26C/9QJmv3yqyj+xOMUYstYrFNg
nas4F5BFueAQkIleRtTXclAuR1hMtkS+LcxAkkxpmChzujH/8fS22Bk9xi0d1OMh
WB7Ns+sh127PPltYgR5Xf7a1V/oAYPLes8Jw32mIsSbKw40N2Fc3Lno2PMPvLImz
ttYcAi/XyShXnyd4gme5Z2D3WHFyPHtngNeMsRwjjF5SQGjLrVHm4FL8WNN9kyh6
wn9RYXdVvy+926OGDwGw78wSOy24yZems2EJ8AwAa5krAW5cKdZjcQGaeAy//VZq
AfxxadqLaSswOeEZ/vzp9LBsc4FrYigkn/uk9Rlc6sGQEY0Drhf0cFD5HbCS1G5Z
HRuzoz1OvwtUlk77yblP9V811Om0t02GRE0FDhJkp4CyRbaoa18qIfNOGwDGOHne
4nREXLIeqD2rCh+HvV2RzOjBc+gVvAYWpziTWN2Bf/IkbdTsq47H53C+EiNpGl74
q8kAudoSKrMqfa25lB/k6DdiSmO64E2ywDMcxUlhw/0dPO94AZPwrZLRlf4xxKnC
B4vRPNLPsdB0luT3DRaYqLtKMnxKjZudPVv2MG7DL4TjGjhYyuTJGElaPoOSR7oB
8AmxD5340IT243PPthGB2Wc+84uFXTin1AvYV+cxShJG/odSxV60Ly4EIJLS2gDA
wtQzlHQRqfrYlcfZ2QPKs8Z67+Nc1AyBUIFvuuqpbKdjCH/Ke2ndYjDDlosNIeU9
j/yTECRjF/wo8Uc277dZIV46CnUyGFaS8Gu8rFpKYI60yhJJCs+bNgm1VIkVNCMC
66tDBQzxc6Utzf8NsTDxXaX7u7sQu5OHxrtcY1FKE2Ml54WIad0fnozxDGoeFVh+
3r9ei97d5UL8tcOMveebUXctW9ubJ77ShrOyWcUBdn5YDE10rM3DTM1Um/IuFg5h
UgeQnqZnpCp57klDV15ysWRdDfXFEJjQDuL1fgEFL8OX6lac2VzWZ8YU62ZV95Dp
DINW6yN2du+K517oIkdS1wWS+lbHmLzOmUNkBtr8KPNxVWiRz0F/6uStU2oaHd+d
qXW1qGC3oMaNNtAPdTI/yacooy/meRkSRt9WENzuFFh3DoPAsP74vbYpPzVXloWO
u8FFN2OZMCvXvbUhpzVB0FzAJgZIbhqQ+mQJsI9Osat9WqbREyCoXbafIYC1iJwk
dpHNkoudZO7I7Cq3ABO1qkxDBJ4/zMfHn6zqVgxUa56m5jZGGe2mkX4hG0yzuCWK
KMX1VT360clsJD8Qno7lDqj6Z0DP8dlUTLRl8hmdQMhZWAVlj5lLAAStaMtMpDD/
dwsHYqERLAu9xrxlPpwTVqz5wd3tDWPX1jf3eg9lv4T3//fzzKtyE2FyPfvUp/T7
Gz6LbwQFwLPQKpS0qFiSTOn2EtdJYs4LS2lp/KCc3E2ZaSkfPYKoK/AArRpPVlbL
fVTweGtcnHCosD/JiLkERn+m95ln/RfLWffV3dRDE8S5tsubSEIi3Lc9vzt4erI5
R+Y2ZVOwTscIhJKwordKFtIEiT8T6/Bu2m33hofkkd3p9iZwychLkiFyBvfRNmy2
yl3mPr6zSEPE2YL1qFhvfdxp0TyAcSBM8G1eU76vJufyQNO1ni+QahJ/UVCg0pUN
J3o+x2DSb5mQa4uWB0TNqhWUUiUphrYqW4po3W1+gwR+vABhXTkdVDoSx5y9k6fm
Bc+/1ro6kW5vHmvRUlHlPIZyxe9HPSP6giuurPB2hgwN40k/nkEZXnxANssr0iIf
9X9KkxTdENy7r2XQFMSKdBZMQozVC4sqcZY5l1pDfAm8yUD3X1cz5OxuJXLg/mOw
SwVd90v5nKtx0GrRQ/PxBU4EnkESM8gwIdBna3b9iXOkxEkNp7ej+j8nHDe8am3Z
DAAWkAekxFR12T/bz1LldTmnK/ak5KbJc8M3bNV5E2KZ69ctdUKZEFzTA9N5a64g
RxqaSsD1als8/9ZRMCXK4hftIIs8FzHwHO/Uzp+F3dzsDuKMo1mLL9l1q4K0nmUh
ZvKzRfmur7vouwXEu/0ZefJ4GsB+uirtC+JB2HDanMdZVLtt+KIDQjTpHQvLGAKM
tkuB2PzD9NmUIyTPQSFKcNmOkNwCQ0P/wf6/FzLt2Ln0nHpnzLXEB98RyjOvJdjr
wZnPnxVScomTSSCEan6e3g7+1xO7VY1Z8qAInb9tlhTlXdl4eBLPG+JPiwvl3sik
z6NNTkFAvecSoQnS9hWnbF2bg7ooFIaor4lzFP+ldTf0pijvI9kVZ9my9FWQXKcI
DKtdzJ06CHQEIpS6K3lZjwaq2P+zrh5rEQVd5s3EuzSgS5LsmEpGvuIO1feONHoi
yPEd93D4UPSEC0vhdxYggQaua2FXN8nXMUjYsGfCFGDqL6J3WErAMg1X6kEsCBRB
hJEIaa3MZd8FkvGi/1YHtkAK/1lWbpHxTP6BnO4a+Md7KJI8ht/AoXvjiq/md1cU
4V9ibvoMugyfbqg+aDoXbmrdyd4rBct3ckPxp1yEBDyR7PrlAqN92OoEqjG+HSF/
GawaTmUA4R/zO7k2n1ASUgC4XYsw71FxD4lrV2nctyUQfbSOVSBbuP3QCDxbCZ+C
rwcA+siv/scoXh7AyNiZy/uPX2IhJjah1/kC2/qlvLXMeuh5ivY6ayteI6YxZNPj
YchCbzQPYiEvvl4Bc3GBC/GVzeJDksj4STADynItvmcrb/zGUw3UN5FKANrRShtR
ax64Ap6PLrfHeLXQKd5mjZERu4tzzAGaNKgI5aaiKbmsR+VAL/FryycSySXNfIv2
GI3JITBVN+TBNctqvsJI24feMVWLHqDMd40TRyyA7T72KHkFBUfZA6H+A4aW7fIm
ZBD9CCAThJQrl6pBD+aM3P3+8HVrEUkTdAIUTLxzhECT4rOjkB5kJ+bhQICdqYQW
fJpZj+vp1v+KtjPWQM8cUhJolWxGSWrSVI3b/bEN/zN1pTvcI5DZ855r/WcmQHs+
efBJOyFdNxjVYMHjCSkhIEuAmmm4iNTuAas79EkfrHpASJniZeFJXyFMfE3CaBX3
PWn8PAI9cpJNFbtIyz4K/kOEUeY/eb3l6whJT9F6xUNOO5BkB9Tga17S2wgG0HNh
c0lVzjjcn4NjOCufNmEgynD//jzSs/k9BpeNN6Lma+tdl+4r0DG1YLb1335dTMtj
o94LlzwklXBeGzW+yTFW8+AYodPLJw243afeCp9Qer0/hiaYsFSqglmUlqWuDyv4
Um3nivP9Yu9qhaNhelk/HcPNnr+dD6trXKKgQUh43LcIkspLNSbmGpwGfi01rATO
dOI8p71IKtMVjKN8JZ+GRUfPm08CQBWPwVt38TELUc2Pbwc0z8aSUzCBEdcv4pZl
OL39s+GaSTcnYu1paACLM6rxzE6cDkReBta6Vy25Xn5BcuS3gqqWEIyHcHsUE8/L
PhRjrEhNefIw++4ah49ThaGJKOClZfY6eBEt0a1DdMpBJqepxNfXpEbH6RjxZ7/E
EVs0VR3lm2bJ47LIjjmIFaZsdwS7otbtstlEXO/tzjZ3IdfB9FxkN4J57KD3qIqs
EWb7g8NUKUGgajSpDmw+j52bQfC6mi49de3RzgjBRCU+Bv/Nm7FRN6d1GLoQXOgY
k+CkcYbfeRW1kdd8q/nvbjuVTtvB7PdEfHC+UeXl7M8scTTgJASqE8z7cURBNzjn
7YOq7z4/Usmpz2wowUNFTJsrA55I7KqvWmsY5Z6OJoXzezXnn420I76xRVRdH9ba
9Hj/knGiptFoxKd/mKPntVhBYwiSKueNtPAAMgzPpdXGFZ+W39rV0v2wrCTYts3i
jy1g07BEvlAGRLJQsyWNiaDp/H8Hk8RZJ4/zOdJs+ypO5t8peT1rhcMq6lZTZ2LT
6stldi0lvBVww4LSU2w2AeX8jxf476OiKyLuVCuWtIdxM6SMQAFHJ8C4mSEdtUA9
DE82JBPqx25qMORQrxjEZbNpFMUmg6DwJ5e8LHDIkRo5GTPJZwreUBGVDgi0Z/BF
XviNg+7JWhQYIKrODwBMApRnos40/PT4pd2UkHu6iADMmAMreMUed1qYJqNXCC03
KpcIlTfrba/B0W6+fkNHF701X+/DCwJq9HPFrSFWodWo07S/A987tw7iV+eUbE47
LyekYcelvU+9kmoYG/r8ClMkJ4e0UD1uZIhe2oQpHmc8wc1msXkBr9BHTozstNw8
WyP39kxHFK/Q89Zr+enFCMhZowwCIcTEqHs+hwAPrzboFN4Qb8gjvBAnMHwvUTjC
8aThV0GFYznGaZB3Plk/xB66CB1brqXPmPtgMruuM0Uf8JGnQTzYOtofQ6/M704e
KteK0JXgKJ5tN94IGfpLBgDUav+HC1/wgstIF5EJBm6wucJM39QJNIddKzwaodSR
lLtLme9KE5RHVGRN6Fs60foGoMYGciFU2P1Ay2CEzGOQbaukLud9CEc7tY5z5Lsw
7cgkfWfUZ+ZzbJN+O1Elsaz7NZRSd7X7tO+YAc2ewQqIg5QCa19OYW6M+9HE5LDX
letgAA/CTNK5Y8VjLt28Vf57PuTP2q+TINuO4I2X0anX6hBK40i7Z6tkU9vgEil1
RbFfb4adzQ7jh7Vudh3sorkH1cyk6nBpsIrg7oBtzvPZBCWvpoV1ACYwESbw40b8
KQpR3jb94hsSlb3uLcRABvvqMxTOt/7TOwJpdomRp8ZVIP+lWF/NritKEBtgBhm2
JBMwLEDgHtZUrDjirDBfoz7G4l7XLtNbgx6IXuj6qBynWtQ2EMBc7KPtB9zPiqv0
jBHoitUG53vXAuRYL8WyqJyn8S2PfOjrW6K4v/NK7LtL9VUswX/Kshsk5an3u9m+
qJIDpsEmMnm91WoBc1M4xLXdeoo7HXn2tC19DgIjY3nDwq7UZlqcUt0ZCnZJ7/M5
V8dvASsm/cumB/c/uLWtvUHk2c4P+B6Sak0qAIgXVOspu5KKEIWalsjag5xe5mBZ
5h7/Tpu+Vf3Nmt2gMnQ8yMnuormhtMmZDKOENiDa1yPbcdE+/ruAYSuID3W/+qSL
PlO7kb7dEJ1Bkr+LoXOeIIZLdH+RevWSqj6Nfs9FR1NJR4oXTLaX7tun3vKuXwGz
zpmeQ+iMmIuwuj4RAkOj+pMkTYB+nT89FKvqD9Y/4BqBxrxbAHuLS2Vjcf5B9P4o
28c9Tg/u0pxF2+0Ati89CqS+oMz5mVOYbOfssVx8MT4v+UCh9HMZWGmtcQ7/+Ido
VmMoCdisIILQOcYTDj26Sqj73Nfk9yh1SZFYhp8AEenoy+VqlfLbTdbvAVcLNujP
gQsM6JaXSe387GYI2iHIR5OexjVJ7yjyjzmqU3An6Ez096xv3VSLULc13Y1E8to9
cMcnuSj31JINDEB2RuS6zGgeMjbOT3vLq7aHQxVD6sAtWJqP6EkwS5nPvsNIXbkS
gZqL82r+U6NnQ9py0xWzMd7Faz33dLoNY3PL7xjBYBZTMnrIC5HA24fhJ82504Ar
PnutZoSb/YTXsAC/SshIqUTeHqqKTknQZaSmydZMYGZxBIHRBAVl5qtAZBBMhtMr
f6yupdCioJxezVAhHkG11sd+5TvwD7CgcKwz7ae64VIhHb+E2D5MeSbxmrJxZ5NN
k6SXtoIYmqUsICInxevFFgwazIvTw4f+AUvSnrvqu+yQ+GP1DPajcmQ4gKjdPoZj
t7tzWvPi1hkVrB5RT4lRZHAevwPFld+W4r2iRRlekTz13szfw4H9fnRGIDknN3VM
wLegjpU1ZatZXrEr4URwwNhDxbohzRdlIzQQCLzlnObxr8DHdnjgUb2oUptG/enH
67dxlSeIQufbVsl0nEq3T5c4Bhzr/qldrz0xKkKLcMU9so8LkLph5/k7W3xdXhhP
ZFxWzp2vtTN6drXUPxKp9O8iLPwFPKcf9i3Uiw2MNopPUTBB2WU4nYDBHvYBehSJ
A2HkUnkCWYorN6z6ZvWsK0TP6Aq11x5+TydvepOAPuhkq8M+2BWMf6rRlrXX2+yv
hJH+FRSxyvVP+12iFb3GKj6djUF5RRAADMuocK2Rpq4mNWptzIwABYt9Bxe1by6q
d6Rt+Q3LTfarcEl2VA4WTobEpwF+jLC1pimggfQlCLbm2iYnU6+0Aml5yiTfytEt
qhCIiAaj2hMZOG1WEZ8DFwFD6xz9HeJQQNrjEro4DNBzGtS6LHBoED31JRqUWmpt
vU1alR2fXKnOgQ6fsiN6tHkr1RSraKxZcAo7/7P0EEN7psQq6CCBVSV7+L2uQEJq
tGtmnG4REjpLffujz4dc8uNjk05qTPfe/nanJsdZ7VXImY6FmAmFXLzzGhV2szFi
z1ELVRk6vXlehLYFdqDR7wLYBA9OH/DZS3nWV6bXGMMSinun0UArN3ISS+BjUW4E
ScOo1YGPC/vr0TgIZzeoiJzVNQfX1lVDlpZFgVXVkWvU5aZFPwespxkqQ0/C9IR5
dF/79c96R0ya8B7jIAbIIKsVbI2sPYzEWvyJtzaRZ5nBXUDUV5R7GeGtn5uUt4kd
bU3nwXu/cqGqO/NtcPrM4lldkzBrhE1znk5PtZQGhk/wWJAHxe0/ZroyFIbby07P
qA6Ou1zYq7wKmwuFp5Ajw0OL/1mwFZSiE4LCSZc4sVmWalsUFdoWdeJOGUCtPi07
esFsVuA/7ZpE0swF6kOpKgrOaJt5dNOVVd2odInqBJTs2Nx2RIqpMWZDoExbZ2FY
QnPmv3rw/GCYG8WzO62n93LU0QPXh5Jv0KJrstorADXHnpbenuBnocS+eFASq5mn
dOIL2zp5NFMBfsDo8sKAdTOaIuaM8O9Ogm8FMbK7mFApY5pm0XfUW+TWaFMlaUge
xVekIPJ1U4XMfgDW5ORTK8f+JnsUYcvubSFetcdV3HD0K4MUQodO+2hUafvARuzE
woEBSPk0hDoz5clE6ckKpnGdFQiOzq4z5hvdqDU/pdq80/zZwGSYMbSofRX0FiTr
dq0v04XRzxUKpdLLOic1b/XQYHeczHS6yxxvZPh82C9UMAG7XTFMuIXMDM7oFfOy
oVvVhIr5R1i0nOn7P97N0Q+/DnO10CRBIN222e7Z51pqiFlV3+5+5N3FI+q1hPf0
26hwCnDs6pR0CaqmZFIkYWb1XHrUlQm5pwnypPjqZUZxP2xPpEiMfg1KB64675Cw
Xj/Y1m9ZVoaC1zcvIFQVp571aJnEv6pChvwo+oBx7kWeVKufGXJlbgWkCYPtwNai
biVGbu8VfwhaCDlzNUs4XUd+Z2V8QcJZEs4wFRaHXtH4efxzm4ZijC2oKC4UWMVt
R2ysQ+Vo00QR2y8vwkwTff4os93xcUyyvyDOL4Goyjs+3O71mGVxCWb2xzy92dKB
VjGUsHUPSTDaKaKHdMy6vQ5IM6yMCzRxUERwtP/56XQMEu+sLMzIiOtwtvSrl2G2
1IZNXXQFlSWUVuAuYGZn1dCFcVuwX6mFQx3kON8rJ5zLq/GfzxPeXzK93k2o6wZb
aO8uA2vTj/6kbB2KlHDkLeyiqWypw2XrKbB5YwvRqjBza30dlRVU00QBpQE2IJ6f
pAPLJiH5x2a5+J5sh9xoJyo0RNgek88f1O51j+IuCDNsHYHj+HFN5yPKq83RA3r6
Oi40wwqA4Om6jtS1QRCh3QrbM8MOgLsDmdxXgq6QYGuXeZCGj6PYAdGnBJclcR+O
qIM8wmS4BhLLTJpMT8eq2/k+T/xWUK4c3fYK+HeeVOYfDuTuMv9qJlBPthsscuOJ
yfrjhIzHt2H7rS6qi15kCZseGo8+ARhz80I6t8+4nEBC23P0U22yfZiZSFLfj+ra
GyhXY/60HQsPIG1b/1DkcBGf5GGEqOiABUjI17PSf3zebLt9aoUus5p6uTsmaEnz
zkXHyOnJmB1XBxsePmW1ENjJGPz/tCISKSpIGq7jqCZkpEOFtnLbcztVfjf8lbcf
RyElvhmeWfy6WbEfUou6wKCpZqJwF5/Fp8VjyFSKDq4gmMw+ygIPpA4yvNesU9eU
+JmMjBB+lN0kO8f9wRSQK4KVlnDuehIIeCgO9MAVPHbgw8FsAgNgF4kxDnI4MMZj
uhSkZuzzlE7IYv7wJaVIiyzC2+kb8K0k00MnxOl/n/cJWYq+uS9GjfjiOqM8OV2Y
l/XuQlGQlyco8fWm5oBteRWH5pWVt4PFxjvlqYeXI1qdhiSoOlH/9AFWQE/LDAnD
lVswgQCiNnFCHSz2bMPvyDsYuPKYESCZX73yQstJT2T/gsFqEaTgZWdY6UWJ0yQf
Br8m1LA9EPkQTmDPvukBSJ6ewDAkieN943O8a/cOigvW1LHNPDGp4Pi0Zja17UTc
7NsQwQQD+0hGpMMAsQFV3ZD2393YyujMVmiHZshNp7KJwzVu4sSgREXHjI7frWGh
5GPoxFJmCcaerMAcMHtfeIrhf9+9nwj1m7WQKBzBpobCKKjWpV0GGhPSs/V9rWcB
mn4rzg1zIWPNgmHEdHM2fLjNVgJiZstAFKEZmjYM4/sUaEXK/NgmMiX/ISavfRAi
rbDF+qmb+G0R+e7/HuHKtRUKHw6DtTT//LRgAkrWPZU0NnPWdm19/il5QoGzfJh1
DFATunlh7cib0Fubd69+eejDsXyY0dBwcSCITzdxVkXfkidEHnqcSoUKX1MMwv7b
Jnt38BT3g2DlNyXlQP9UvaRfuRKRiOkOPczjSNfE4347t7CZtljyCyQTxsejr9nx
vn5hfXrsWcIwuvDVlv6aarK5JTscIYiejOXpRx1I4RvwajiWRtYjJGLapk0HbFIY
0/q/8V2Xn5wdwrLx0wwzKrpaRRLK5LGrzZxer0B+Bxk24fRuWEaxYY5kjMais+VU
CgM6mI7AeheHAsNEuQ3iYwDTwvcfRFz+goBlN2o7H+mILDds4HkMlVynC06BpbDZ
7W3SJDwEHaG5GYKLOBhZOfv6olq8q2cLS4y753h+/TBc1d4W0dTmvPfeOQ2hWUaT
z8yU+6IKE8sXPOFmFHf4fojru9mmJe3aJzzvy0D00FXaTDcEzZQWxiQU+MMUoLJI
1NKKeiqHu0plkRErkBsoTHY9VGtrDvjyoirw8szOZ3nfCbTzZBVtNlvd/4IihRD1
KYVIouOyZpNR4zlfMeusZUcQ1MZsDRKctwgxRMY6z3vXf5GlM3bViAYiMzYszbrn
y9WlPmCbk9DonOrjPqTPqYtWUAkioJOCm6Jn2qTdLERYnXFF8FmFRGN8lfHYgO0N
3msdrJUixdGDHtNu2BAepIkROP5wgDbzKUecDAuEXsw+vWumUyRMv27+LBSq5D8u
nFIB5aVdTrA1RexFX2bKf3XO1K48Gt3Rdrhi2h0jd3Y087OfgmFosiaE2P4hU7id
EwfAKNrbGDncH/5EjcLDu7YirCE0ekrlAZDyu7uO2JnbnNRA7Mdk0uwdHxdGbRiu
YIgtZ3d1oXosC828jHuTFWlFuP/LXrN3zOwuGriT24vD0A5lKKNb6E1PAD3kVn8x
Qs2i1ygCfpj7GwZRg3ZL+tEheVAKa6vqWnwui+XMeeISIMYYJ4ZOzjYNxzo5BdrV
ccDYbIdszTUVTMrRH+A9shNK9bZERa4Sol4e+f0X6CNnZkS0V0F5B8Rfew4xOkSG
pcPjnysrUfV5Rv6c7U5KUuiHKOB0pFEodQcTjlZnxxpy2jhVx+re3I+0ul4/ShBI
4NgQg5ZLhrnxiZFqGPPpgZ9pK53ypWjtaCfIV0jweYPdVjvuABZyNV8lm95MGkJm
i/6PPyO52h4zS19hZHckl5RNAqtQG5xXIsBvRp+DBFjaT3Gtyed0lGy7E5Wes7Gf
xs2cpK4S+I8b+zDR5dO6+OOdVvtx4jmXFg6kQrHK4Qh/yNPrVycvZLIaQCMRHdk5
QGEPnRBLHi5cKVpxX8QiptUZjOF6uLEProhBKe3cvGzvGJVU3FEi7Gp9nzyGiafk
sxgJSwjnHKgAAcZkBmfnjjypR8dugZmYrzY3zt6S+bdLVDkLjHnibKgnRFA9oq1y
Ec5mpvrnXeGA6LLCWOQJkpzURrB1cHquO1FJTDXi1aioMnxUK+NOAWq9Kh+gjhOM
rnC8D50NIHx07++EHnE+OHKLxkMiHJfm2t2KqVWMI0SnHl2AmXWHgQp5mxI5mt8Z
fkXCP4Mmhnabgxtf3GMtX1maUq6JVPsxS7MOcxrX6K9L1LLB4wBNRM8Q8WIJrDmJ
RUVTzitLN4aYKeWGa3ORwB4gAtZTiJ1uw0h0aiqiZauMtrHWrpz7nbb/bT3JPPgn
kbCF88see26QYdJDKxBiiLn7ViYgOo5wGfowNvcnOFuWYn1BZcmGOU+ZKkcfK1sb
AO2V/+YXo1UjJ/WQmHtdbL4E68sHYRE/bfFB4m5qRrmlFXvwwB7MJoIFpXJnmxWa
NHC1iELL2TIVU8VPshuQDzjPh81HYX5F9YFr661rSyURP3lPF2A93vGUK3WBAcm/
PJQqYhq8WH8xdiJrnRWIpWQDP/a0bQ8Y7YzxWoXlDeDLA3PvxUbiglUJVrzjWeDp
lImiATF+zN0Jgk56RGNQMYU9mkxiC0X0c9c1wk3D2IAFzEzVhh+2eri+M4Qt8SA0
xYW6488RoOWITRWbr3f0bqt+N7lE6+xfVtCsZKrgwnIWRJEsbvyAw6oIUF/QP1f2
gZ82JHrP/OAoTJJUTiL6Lp0nY3OZ2d0uSwRfwba47FOCcDp8TANyEDRL4lALT7UX
It4uRug9YSr5tUyObdwqBQgdBXCpHxeefcy4Y0SpVRXnMDY3XerHxGQ305EfmDry
3b4zjQH0JHhc7DgOrBZg3IgM2w6Ej3Mm8fZ/H+hEWVCl5x/VB/wycEPBoY9mht47
N8yTbRyF8Vnl0OXWAYMj9e/1e9vg+Fk0DSSwlmOYcMGbNE4U0M+vCJGYkuC/5gcb
HCazgQzzupvvKfBCWDZYWtllkOipGe/Sks81Kio+470dgB4LtLOZ9xbf0cCvMsp1
IKOEMjBHGc09w3QKfVbUa67FcMQyZ9HHlIXm7yDZcD9MHfWI1ChmEKnqlN7ctWMr
w/y+Hcip7h6mmBZ4bDNQ/xdr+2NyKGJSQql2nVI0zlP+1TGiU6hEU6SJmF6pqOi4
dp04vZW9nqsQZLiiv/St3Eko68Os2GrFpiIIanzTIYPjGlO5nevZZERT2Lo4siIL
UA7UbYDn6S/7VEPqDvfvXDd0hZE26wfCZtHrcg34N7/ap8yC1yh5gtp3anNBKV6S
APs9d/Yfuc5C57CpeWVhCFMOsmOViBhN9IY0gO+Uh2faBcLn9AV3WELljVxwAnb2
HwKrcseLtjmfPrmhFZ+AROw8oPEmEvHIYxhx61YZNO45vqCwE6iWdC9CYHoO0KuH
pdXjE2mp3uF2zfVFWDITESsqJsfbHBnPxzEcUU3zNT5NVwRGzTmskbzvoLSJ4ZyM
B0KMiGQaTPUpLhXLielR/5tc4z2pBMNhQWdGKwVynT1eL7AEWhij9lRF7YsrWppa
s/WKaXn/v9SlYwZBzOUD1V61Ahj6oSvqHkE0o5tbxYkhG9L+wQ4gSHgJLOO074Pl
tct3KEJU1OYAchE/pToXfDEDIJ9H5ttKniftIuFWCD4YJ+BkymKlmCS1vC9c0FCt
9cPkSP58pZL6jIdmW7WWPUtOUmA3811hCedSGqh6eQeUKJO0to0DLaK2OpMYymaB
dR3XY+Za7tLavzq7uI5DnyrvajlKcY39fGgZ2ZqXZpVlP+xb7WgrmZ2IzoPEHHf0
jKOSHuiEpQzdgxKcK32A/ixb94DsYZMEyqMUHu4bNbUonRrGjeSHX7aZ1QRMq35e
HaGVa/Oa9sDJTlx+1sg4nrN2FAcK78ex2HkeQ9k8ZKT2+C9CQgLsTAhtXzmAOQ/Z
Xbw7DRVB8HUwR8JL8RaVqkTaOsVGSZ15y1fbyGnq4jWPT4cWLkqRz+s8s6g0vVW9
C5vlAo7igPsDvb+2VOwgBrVGAX3Q/d01LOcTvTlh7Tx58LCxgQd1by6FsDzoVMim
/qvn4x6Ny46rUTV+ymnrFRdsP7ndke2icpNFiV7km3PIeb+XsMrs/d5Vz0Epf7PC
wWT8dd7o3S9RcKywJlzJPMfLqbktGTufETqwor1Ow0YtIl2AflpHvaWzahOqFaJe
+xjtVq35CD9W08Q/LYTSJLWnjBbVChObuhNvj+de2W7aH+5US+Dey4c+uLXI5v0F
ARMk6WYrRDAaRfLKTP35Gvi159G9uxtsZLakellrwzyGQ2vFNHI3GCOoYhoDYSMo
RE67BGs8dkLbQEolVocwX1x+evj6s5hT+8O7wpbx5scGkjlO3L0ccKhUkLaQ4jo3
LBYNd1XQlMx5G8KgUvmadPUIWSPApmzXVYnfQCZZ0BxbbxbaQp7G+xKGOSNcRc8/
X2ZzmUQEGTrjdqQ5k5ED41HE1xLRoIhlkwbzLqOwi3luVawk5Sx0Qacbw982ZivB
fZ/UIvQqCrt0BEgXmfd79TU/CczYQjfBmSllIAhmEFAQwFGhgmfStx9mnye09X27
OFcwbwmuMtHezkyR54Y7dZ8fNOKAjrBIKJoxWjoEfzoSF3A/Tp6yWQoF+EBgfCBw
A0CXlTstr3laW2NgKTuGOxl+CadEg8TdZHcm2ApDM+srz9Z+mcUm679sD4jUot35
8v5c5fenCtaZs0M++yMJZ9OoGFKTHLHv7DY7lUgVwF43Dmk6qVd8iDnkmysIvARV
ubSc6mPuiHAlHfEEVMRIT2R8Prh8QhTksVujYVnmhsm0QWzA/HlXrQiVgtoGvqqE
MRiWKxo76SZ8alrn6Mvx7zcI2i4K8hPRuDhXh2DkYOb0K3b0Epl5yuqsoqZ2J7mR
SVH2Z2l9vtzuvddy79iADGdqQENIp9T2j/iNnx75CX6btlNdDVLn+BgTWyAfPFHY
ZcE3E3ld7tm1yHx9O8czFCpH5hPbn/3Emn+qAquaLB8Op62on5uwlZ1wg3IzdyBV
93Fq9bgBeXgpGum+JQOfQsCJCXzgy1+95cIMj3QOJXKqRzMaMOrmBMulthJBJKEI
xsznJRz/vV+v1AldMPuIlC3QIoLrcat0eDHuFyxwYrFs3h1XaZCtkR3GuGodg3QD
moj0T5M1nj9qgpuhE5DRBR/METRsJVsDdr02kQDJBQavr6u/8D41UrQVkXAcc/uQ
UaUZN6VNG691cXMq8RRLiivxBM2FWcBgua8ri8WqssRwpfHIlrEkeoT0eXHQnHCc
RbSfrqWnJvwzMvRFfEHZFn2g/Cuq30soRZjwRfMPe9dXfg97S2wY5gUKfeJzarMD
dJst3/M7Fphbsd5G/fMWjTMttTGd0AALRB7vzKZ6LsrkEcyIPjlCgtbdQkp4Gd1A
LtitmAPpDO9TwRtcMgzMbPmatMHasJMyka5mDTY2OYn6KY+ywexSivh4hQ3cOIFd
aM1Ic0BmD53MkkKJHekTsu2ta1evH6+qJ9wLryH4WElFUg275EA2m2rd5Pv349PW
mwZuY0E/ybLstvotYRR8DfnW4bNC+EAtV3/ULsmNin5VcYt3vvKoJKNqKIwp3/dR
ZW27r1hbjnP0CUU14ZVm35eRxudrxmW1MeD7gN2oLjWc1qpKGctkwJFfy+7tFMej
XyEH/1WpeZXXrLhLEYOwKHQDEOPbeyw00eJEibZ/kq0ezqS0oH76fqNBD0ZQJZw9
emZHLyUH1zHLfLy72EWS2iFYRlG53PFNiPmrS21HIkl8IAc72+N+cxIAXAqEpfuO
zQ6yarKM5HKfJ7WhRu3lechnRfx13qej+qYLR7po9o5BSEfaueXp+ijaWM3O/A6S
JVSyd83ztpED2vcKKMBBd9wpSKvFY5nU8q/G0ilNYYWOTXMhcbsYV1ayD1FrG9+j
RM1VBVVHa8U0qZ3CQvLn6/pLPo38/Tb/G0roLkrJ91SM8fxDaJ+SJEn1X4ATcfse
d0EWKD/etmcMd5zl3TMCkc561jeUy/g20x80ds04lObi14CKPWe16yhN0wxVn6Uj
vS7wQgVKPsV3BERaWe89rcU/+lx4Awb32E1qFI3n/D0eGgE9MnXabtcUBvyKl+jj
lOWE9O4LPvb9IczqRTSnERXuPymNThDTIghbH4Ekg2lbIKNbvJaMQXFbt7YcrKOe
ztR6FRc7Zfg6HUvp7VIRiDV01zibClLveJfJ1R4gyAXtZNpbp6BsduQol8z8C0JH
EEI1WOvT9H/1txOO5Ck9/0FJ/yvxxkKR30v63CbuJehJ59IaiDgR6u7EhyiWKHps
gDjxT3lmNxD6p8VJzu1Nl4SAdeIOv+Ejws1wVVpUdJ1Z3srgbyxxW3zsL+9+O2IB
dUY5/GaNtditV6SqMVp9WQ6bxrnlbmAyljfubDNg4NMivAldV9XuDiv0c0bmIruO
yBpleW/uom2145WhUiwmbeMVxWCdMhaixJOvREhpSrW97xumobgJmErhdxeNVQJ9
QiM3xW3BZbF1jXSK0Vv0dfINiUxqytd//L1Q0bJw4RE7z2AD+EwMOmNfx2fIJtyv
d94RyQPuy91mgYSFqeMljN+OQrO1zwHJh9pWjwEeOp9qC5WZS9Dq9VlTIF4uqzLX
2GEXJCl4A7jdbiUlVwNn6Q0cMf/Cx6a78EAF5UaKMY/uRNz4N8U2HreBntF4k/uu
t7gmhmn3ACmNrZzCZpJw131ECY8IDBSPhpJEXId1ALbPnm9VreoMY927dijJItCI
4A6DeAQ89y0tlJa18LpLbcl9IajuNXyONEmLj8vMDA+rTNdg3U6LmBer0TBVEiSP
E07TlC9hva61x9x2T+uSp0l5kZhHfBK7x7oWyITXASyvAPd02zEFL9WdAuIYD1yX
VDmyetxkWA2O4tOvlVeErzIS5yaePn28npbvZtdjTM0dYk0hSYkQU7kS75e3iRiO
1KteyZ56wN70We5+zPvbgIzUBYy9vgvEovthmuUCz7EHY/wqk74PJZ5Hyu2BzjPX
oQl9WgKutkV3jDbkL9bqQghoXlf6EzohV89MYbwUWSp7JhBGwheySeKouqpiXL69
7nPdb3g+xpP4hmlzP1ruxuITa57EOS+0bzCBOFU7dqfN069sbpKGDtalgPyHwYKN
1oQXpoGMYDO32PLyV08UmVv6tUv2lHS4UrKD3IuFvyi6cDNBbsvfoahlj/aTFEYm
qO3HLSqQXxEaqWPT5XZUPJIhbxbZYmRTkU8wSiVWyEnhPuUZzFsDMYvZ/LYvTNzW
xhlzJrWq0jmXtwMlGaURsImRR7rNo8Q2VErsG/X+dJ+9lYA6JqtLpLlrZ5V9ibp9
5vN1u3W76axE9bVRYfGRsWCVlXUNenD3T27UASsx2mqJ3zWElzo4FrL9QXmo9Rms
Dy0WjR4SUdgc1geWA4Hz4kaYwgBwTxeGW5DtcZZjci6Q3n0pfuYrSRrgJ3kLf7AW
1j5xPMROGxNbcQcivYq+7G77NlXShFrVnYtJfGIKgEgzh5fSlG/QvaERCArD3ZU8
T4CHEWH3Lmms05hzFkpAAU8coyydOGooTBi+Nc4C7v+Cj+A7/Sdcbk+9uYCr9+iA
LPtjjjAhM4/LuA/jVi656bvknYJyRXT67Bl44xeoX8un6s8kEEsYbOxAT5PKKm8+
9L9o+wmav6RulRnlvuS3EK/OkyV6LXBEyxc97ayWEqWEtIh/7QoW5QQ76Mb02cQH
JWorhz/bIJdUH6u7UUZ6GDj0L58wnXPFENHfNU7V4h8yKDjE4trAc1lWv0eYKaSp
GZbhKrWTq2kvPkST+ntPm0GRTpS618jiJEdFRmDv3f/qNpnUFg58CQ+02SMyWmqN
U9fuHH1IfFywvJ7PccJFhcQL7RRI8Y+nWuBofm9kNJJQNLp9EjGlLOSaKuGR6fMK
Zv1Ki71z5GQjNbXCSGoXmkv0U6J64U0/CKCp/996tM0sLaGam/cVkGBiILkdSBB1
0KoiXq2m5GyIONOtoS02kYGoWQxkKTjqCcjmg9KK+1Gwz9axxN7M62gkGHLjcsQD
jehdX1r8SspxIcOtFFAD/rRvTETcjY8MkjanFPe90fLadhHD5kP1PqrA9XdsaLww
uRFn9st8G1Mifp+ldyTIF4wAqdPrtHAu/fd3eZVdAd6vfsN5hxFaB3HdQu4x8CBD
Z+vUKVhHhTfIrPmhQjo/egs2nt4Iq9TfTZo9oKDwWzKmGq9nIuXb+iOvNwojV3c5
ADMV1AxfR4nKHHLB5KoxzlphxnEuwNplKie7PVOV82hnyyOdOUUIXPnMyFlBL9sb
8UXRf6GFMfq4VRYsQYhgHGRyzQJObe+Vok+XIh9fcs+103WexxzT6pt7qo0ke/IQ
KI9VQGO4nFU8Zs/LDD9ROnXh8VJT8s8aMy0w2wKWhUzG0xxGqlbI1bEdjA3oc5u6
3XOGQ/RN9QqMRfVEnFLNlKIcrndFOs/u9rHi82ZaiZLtF5awk+RJglU9/DeODVw7
YuR3vtTWZjbixXSa2+IHkpuwSgOMIrjLwceoajZBMcYK+cg70f/TYQ/CTioH7VtO
V5q4KbhEABqCNMUPYKE5pj6YeCkGODpBDCr7PZjomgjcnahUWklCqfNx3wB3jVPZ
pA+xecZmt54QAT0bMD1s2R+hmDAnNIN6fkkhDt+KReBtys+ElYarOKLQbTg4x21X
7omIpRyNOYa7pcT380QBlEjZuv6vF/nCAKQ2UkM888KsXwgdnLyV2vkhhIbPKf3i
SWPJa9LlLGocbinvZjoWqbUVWOlUU01UavdCPfUIcW1AYtG3jL6MXeUe4m6++F7d
4tj1fjGjE0Mb6hTbNNJheEWhqJkp9qC/fZ70LtemW7ycNMACC/fTK1uoNVfXkhYW
y9WmkvdVlTQ3SgDKv4JUTv4N/Q4kafwvZ5FDcidRPy1EgPYCR+GO/WHznd5rcUFk
WVqEci4AOirJG80aFJYjExOzhEc+d368FsIgOnJJznbal77tMxfGmCnMiwGUQiEv
oNo/rrp3Kar2AHgU/qjCZFdzJcSt+kgHjLkTYwx52BfLcjmH4RKy7OBq+APyUdMK
pKFnql2/hLQ6JIbMgbGSDXs4bIO4XbolVB6PikbrUA1vZnzrk2OIVET6LW1mwOgE
ndaLUAKvsKF1YCWRCvfrEoqcYALU7fFolUGeBJHl+rde+7YUik+hVnO0iyJH4PAM
wxedHx/Q5d2garWo6r5EoTSx6FOi396/ZQSwj5okfyn/voyktZq4nGQG6nHioQE3
xVpd+y+2/NTggC4EWzfXhre8wccE/OrFQSlLqm1eX/WR5l19fsnXb5uufAnp+cZv
Pt4AuXmF2SxjZtyXvVgQ/hCSzRBjPWS94Yzx0pVBKI5dKXVJCCjfKdHbrJn9mzds
MWJdAnH8B5GCbwaFM0SgEzlHSsFVxL84RoPqSv5cP1VyBCKhNfVqoHz5752q6Uwm
yQj+KisyKR7fIw++dmuVAwBhnWTaWjJ/JD8CEjrJcch8OlzHGHeqBYf84S1hIfdt
JwETHJDhE0RmBng+itOgmHVfowzyeiTBmVSwF2l40e4kN5Q/bECX92jI3UlC7rsQ
SM9mqg03PZBcaxfhpDYpJK3B9QxoqrpZx13pWlFX+CP4Qm9NsbOYr2F/feiThtDD
L3MX095XFZlAiWbXSR1J1GH4XOkrfucDIjN4QISWe/NXl8OucsluRPxyXqri2uLe
r+Ma52bQVf4Y7EtOWuf9W0SITk404/DI6bzhFjcBWiLL13n7XlAuZi/SYPIw4EAG
Sj4lT426+8l5bHv8xfz/frlJSNEF6MafQV7u37Fno2+T56BqN+SCqv6dB8IjWkx1
LLq76vQkTgt+Y6xB/XV4Nl08OJOUOPEicf/zKzsSWmz5mKOhPsLcp5OXHKLDX8u0
lqoCKj+lKNbVGISB1RGWu8+r6P/dW4eKnLujfeb8fbp4ngr0ftdEgjkXLqEaMWuy
z5w/YxjAe00R1dONjZSq5BB6pcJeUfGpnsZgVPMAJykBruUx4X0iAioo7yUxSfk5
1ofCCxDfkYLAIRZfsbCTwvAHOYzxsrsbBOQP0Hn9gJBPrj2Q5Ppvw3X/oVpZeXqz
/C1JvsA3eQ9FW7ANvaGB2uJeGLjCoQwVkU/2iZ2SsljU6nYYAREeXQlVfDcXeMTs
B8/LmhIODM15+oh5DoMvb4uUZTFP/yXRM3kq/ad1u/l2mGVHOnKQAqyxFLh9ihf+
sEY9LKBA74+gs25w7xLVQQRzNdlR+8g0inQyIqvXqki30Rme/NGTrBsxxVQSWCEU
TuRVJwzIXT376rT5pbJI2vZUdbwEbI2Tz/Hw1Eso22ZYReED6/5U65QJl6K8VZUu
nviV48J3KVaGNsPiw6QmC+OKYICLd1bl21S0mSTLDbkUv0EQVQkalgDbzhoK/h09
WGjjkWr4QquMQAEhlMQCfMUVw9iAIbJEDno2+pPoJHFEemIqiizTvKmm6QuVXC25
zhjtEi9WNy7+7KwOUJr3wSH88l82+uNwXgw4wELlUE3tu/l4dWuFPB403D2sIbJn
v9i6T/liw9eZ7obKpPP+GSfmGPBrGgDmJE9VxpUe/Ok3kYslq3UQ5aW+xNO41nHs
fM9IcuH7pr//9YAoTuKzdIFgo+cfsb4NE+oO0givzUW3W9SV5I9ytUokfkARcYEe
V5taahiupR4GlXUElsjviZ+HVR3ha8ZwEGl1UetCd3SCwpmgKNQVhdJhbsF4popn
WuSpcDDRDsfXUwYIi9569CwZRbXH2rCgCLlkRmuc82yGGaIiP8MzqUjKstHq4Az1
E1xLC8LB0b8MCk/E45dYF/7tzG1oBdZkKU9v93WTJn3jkxjR356JHCbPnD/uwPd5
esX4jOqKb2QAhqW+jeqU4aSXqZ2TSc43bko6GwZQeXMbCRMcQBH9w5FpPgC0xqE6
KbQOrzRga7HVirtq5K9JTT6aYT7YhDB3sOLiYbDfdipBX5yhNlnPeZMQHQ9Rvy8w
ccQbKIlsiWZR8Ixe1JCNT6DToPQIHNxAzkLogWUpSc2MmNuv9/FDAiw3qJFcY/zE
TneQZX3zNSn/wzBBIeALVKpez8dviR3EAhQSF0CyldTEPVD1MS8RE2SYjotoEd63
R5VOUJ67bRDUvGwdtYX99mu2IHAEdnR9JHADKiynd6nPfPIZ8MQTdXGN2iLQDLd2
XVGaU+BIas+a12PTg7pBuQaHFUjkPC+0csHF0T/ngpB0BgiYBJqNMtHyQRVQJ8Ep
y8qbjRiFwffLupcD7MoBRpcjIc6KzZIuZj9Dv4AIcwdSjSkYTbXEE9BI3PNSTYMx
qj8zrb/ulhpDimPOXCEpKUViXoWhhPopv26N2W8xbkXQruOoOMisXMtEzdJHa8Jr
Ajk8dS1zANo4UOTZhLIY4//9OpnnY9AHe3dpvVkyQfzCaT5mWcvMfBtV4THH5jr4
izZvUcLTVoEFqw2I5r6SXsYlQey0XGJ034wfhR4KS/yyNq3g+eud4CKInddQDf6o
7caJtH1y6iO1CRJhqysjSQ06e8CjFfOSxKOEd+lQmEU1Va87aiSBKpnPf3aGDtQi
4FD3vXhLzBpBCSDNHh6Bj6Hsk/xLvzsKqND44sN7vTDLG39DpVy/U+WI19DUPIcB
JYnHAOjiayvwvWWvSvy7e/KKlcOgIAcQTrpuvc+IE+jCmAJc2MN/fluzEbWEiHbG
EqVNzxDUMJDa22N4IvzeV7/OSBOXsE3DzHFeGHt2ZemEE0fl+qpcGyGPBTF0ZB5L
LNosv9SffRUlq4rJ0ys/hhPV4c0FKtyQOb4YuzEkdl9QiZWdQ7MW2ZOHcHewnqE3
CKOe23VMgfxo5T9k+Upofm0MihEbUBjB/6f/bbo3yyoWh5jz+oHPekkl00nanpUM
nV1DZhQElHYlJiUycMRojTza2AeLH9oWx7zrN1z4NT0E7zwQbyqCm/W8HD46Eadh
y45ZD0aAl0qbdl3MYaXgfMOK18oFmTOS3obzZphCuSRZblwr/JF7ieLc5WJOYpJq
1GmAcw3sC+TuwEl4bpkTzpBVU/Ho+zTTeGA+cnk/tRiEvxuv331oeB9J5kPN3xzw
PUGbXX3BgYQUHU+UB7Ikv5W16jNDFLc1Y17flgi4ZuAulwSRCLnIeZ/zByEXfFFn
w4v1llCKWlWZ/DaIpnWwNFmTMlyGpCvU4mm03mhgnAb9bSDaFb32r72VYRdf5bOw
jfZ5HWgHUjDkYMzBQzm4FFGpV5DWjlCF7g4uudnR8C3Tedoih0oYMn81oj8Lr08T
/KjcGtCW2BPBJZ9zFzyT3iRGGiCrRyP5Z3f+ELUK2LBtAjvyfbmEINdPSy4OBaX/
tgcwpjhZhb/OAf2oM6qx+7h+Fz+Mc2AgiUqKnAvch4h6l/zDBcJlM9K330gO82ln
Sk7fPYVFSdGd74ipBQjyFogB2lGE5lcXyS14+4Kp4wh5sIhngtI3RjhiFDbM4n/S
//nko4AOuEB3t2d52P1EsQHSadFAvVpieF3YW+M/d/zCrUpcijV6Iv87O4VnTQIB
nwiAK7wMoz2cSY/ZT7hKuejQZe0sTxpRW0MDVtX2RBw5gAuWlkJp1wW7oAwvii6z
ZNvW5wbaXJqhZDeEaAhalAwKHrWm3vPC+WQaaGlBjSQZpU03GGi0Y7VcHsyOlesa
tb0119hxWs4Qs4wrSLVAC0dCXmHGj4DpwlSQcPy5TfyBf7sTSZbB2d6CMU59Sw/Q
6217U19k1lvMk6uTcF0qfpGqSii8+DkzVD0kO7rcyyvdn9ZcOVPqNMbAJT6AiRcp
gr5juqYYjx1eMFoeNvltjELoMeK8M1Q4sWGF7EFkATQ8oJM2lYliKsJz6h4zb6Wr
iZkUvUiwDYI0VdHPCGrIpipqpJUoS7V+kJH8KtoC4tJOw2ivx/dR43ByX/c9XOJX
fM7KB20dfhGXam1+kTtC2fiW4e/NooWwh6ZimFZ+bOGP34CVAbh/sOtjrroyQsIp
kpFpUDbL2Huv/iBaaYu4VH5ideTOKC1KrzeniW/ExdY62cYAMstOh3igTbLL0D4m
nZvEjSpKF4P39HhwLBC4V0AHcjoO+5fbvpaiCGrGmHX7mwITXcQeA1EoUP5/bVD3
Yi3Ap025NOoHdUgNJbITxCq4dBt4KhCqBKYYFUqm55S5h9zdej0N+N2oCQliM3Z9
XeleWr8t+Mqsyt9wZtYqe5xRHMUFWo16G+zhTY3KW4Agpt9c/oSm6KVP880Z5tRv
zTuoVusSxfneX8S0VQJsIkahK1iJlO6Zy1/6M80k499YtJ45bnEcn+viNzgFbMVn
PVaZIZVPB+xEAojMgBS0wZBixr4Mem0qv2K/5m8uyc5dGOW3VDtgTAbaSSS6QC3z
y2DoOrmns+Qf9uuw3BHCN14k0p24+OYmf9YalZSPD2SNKfvmJ6yMHjqrobJoeB2v
8wsT1AXjgZUv3JQYOjXD7qZeMeFD0inB3BMjF6Sup5Y/CaDwP7+rEXRgtWfmT7sO
k/ASEATRO/+EDwJdlrGHK/VmUryX0/FbYWVTz2nbOtnw099TZd1lQ9NUxetRlHS5
52EIv5C1NQbkj3h8jxeAD4DJPbSDNrsnODjuOz3PgNd/KODblyt+nCNlnJ0kvJCs
Jrr6jZVGuQOSA/qjV/1qUrZlsYACkwVnQ2xbJ//I+F3HEkl3ulOBM9LZbKgpZIgz
YO1Ia97Ra6XiyjKhAiY6katl1SmKGFsuNoWTkj9xNO2FitlJxpNlRRAcjoEOSdf9
+njT7kU9YXbYx5uJB8J69Ebrc5obxhzmrGcni4SfT/BCogy3nv7uZUBykxZl5+Eq
RZQDVVB0tqRHcuE3yLd+vF1FZB61oilnpFWqRmV0726sKX3MvuxGTP5SIRu+pp05
r451TRCYm1XBWMnLbPgYQj5REy3JAsoZXtX819G24MQ0BjgxmouTl+51G9FTaTa6
E2bVwNjRhVjy5a7rfYqlezkHmDqTFs9sij4OZueamruJJhVrSMS4sTnc6tVN2DGx
97XIxGqzN+3R5ExGtqCG9aJrUiuupRgrhkRJT2GV9O+Ob1ehW+uJGn/3Lpl1xizq
R2hWStgWvv++KGdIlKsrPaXJjr1qazn1y2502NioHdYTApa23UXMC7sCsg8OJPR3
4LDP46dXuQh8mUg+V2eM5JvqkcgWPKH12O3XU7YAH0c2/TCNbDdIePLOAZjF37rR
h3IxCpQODUXkt5Dq17jORRTkznmNvO2oIxQxPEivEshXGiJmEZEN8o8dWVHl72gy
JWKIkChYzbJm1p7DMnlRkK6oT0ZgtXV7yPLmBnKoa+URj+lyaFW2xs5JinezouaE
tucKjz1z10poQ56itcweXduXv1f4WXm7hCZmu7CO3EqvLm0blTEHlfqqZkVTgQG5
Xoi0UFa1ee9XskFMIbyhXMWH4pFk5u7g1By7ZbedQ6FAZnf44gyhHTOzh9oYlpNg
RJv3nsttIaO6x6RovNh2l6evdXy0KqfQUVnHNr1Vy/bF2oCIy1tFamqOj+SZxQK1
w2LOm81cC05I5zi6utpW3blgvAqOl0+tlk3cpj4p38V9IJb2L1Qu/cBEHDUfX5kr
5vkTnY6q0V7zEKM6IIT1Amz9aa0/VNq+G1h6P7mjrEu8JhksZOw3i4WxTilEDzQ8
8jZdsGUy90fW3/G89GdY5rIioydAnOYvSlW/hmiKjKc6lWc+TXlsEh7hosFV9Vw2
RikRVPl8wrt1xopvu3GzryiZOn5yyqX6Bmcp1ApdwmASLnKcj1M4FhBurVQO44O+
AMDZwEFiTLdiEYyeoAk2z3eghToIyDlBOZJ1RaskVOJcxqR1zHaTh9MiVaXrq2xf
mqwpBQvlBx7Wmv8ewKDg3nLLQkvL76dFb7dSNSGJzI9bP7rfYATD7k+aSGoUVRx9
p4LRHTFaBjXlYVWmPuVBuW5nSd0aIeuBq8xlLpA9yhf1C1Yf3934dVNO51ZrZH/V
UBVJBZVOk5evGT+V7hzKQKhItR2TrCDR3zYtkgNTiAjzJ7T7ZdGBXEj40+lQahNc
xwKCnqNDwY1qxbdP3AdN6LuRryOTcOcvJkSURCfydhRhIzU5Vkla46sLQFuQelpD
HFLtJp5c4i5/ZGGKzQ1BhGYeiRw/HwDkedliXEJV4U9sOCOwJ2X7+GsmbppC4liB
F8JDmHLOZXcqkkyFbqulQNB2D++Er8VSjHYxMcdC8hRhklCRzYgW1nMikKlq9BK7
Eei4FlTmkJJSmuMzT4pEiQH9iKo8vA4rgoiRKh6Gj8x4zk4mVcWQg4spk05w/gDd
ASSCbPcaNQv7cRJHrAHPLBSMqZacIbGApY5gagGPlEUnR+T8md1by+5c7BQykC37
YM3HI1dXUbIkkIM16EHniI/b8eyEBsrsRZCLlJWaqZpr6KASrGVxwbp6JupUcwpU
cZTvgRsbSyS3CTxiTzTHeknC2tUvGn1OB7DfYC7G3Li42vxuQqDyUDSWu4YUb9cE
Mn74h/ZtV48Jv18hYZAN+7KeiFjheocTMV0qv1LyVtUUXSSGsvpKTeRfIor+AiM3
mlj+hitdqvEn1PoKmzdP15vHGoRjuZDrFdphbC1sj5V/yaRQEWo5wyMdVizBMJUh
zaDXFQnwVWNuC3mOcIlz15KBvq9BHCTxH1VcTeSAGQ9lXYy7nbxVbLhQBeXVr8yg
LG8Wd6LajDgx6Svwp4duAuzOWqpSamT9dQyuI142co1KoyBuQOqYKsDv0Vt3X75I
F5Mcn6kI9Oe8qVSF9nBYJrAd3IlVKaF95j7zYPJsV9siDCtF7HtZXUzX8snJkLqb
iFVtgawZdBpnM4qiEpL3OBq4ID69F2ezfbhldi1pKwCBr5qOqlFGlu8wX0oVMAvm
Uv8y+DnQ26nM9czQzew00l0diCR7K7Tustrrw6+VBelIyRrt1PxWOBg31FDnID8f
MUxKgIfqVMfzmY0zJ/V93BFwwwSTp+HDYlKlYbIQquVDzoquBpYhBI6ncFCARAMF
g0r2FZO593A2KTy6VqrO10wan8iK10OQb9g5lgkqeuj9XU75vhdMxTQ/vGui/SwN
k6DIVtZ3hSGbHL3frhB6pULwd9NqG7GzN+slrCarcVvCz44NuRY2oXqnhg0qAIkl
yFPjZfJETUAGAlPcUUP/8KKZDd9iPz+3yXsD1Iv0SX+7MR50JMT92RBEJZASAS1h
BopTbIJTWqQ6W0ajM9gq5zkqKY3vSwxD/eyAqh4rEeTqnu28I3PtUntU/BIID79S
IRSCh986lTTqvdo6ityaZl0alhellcH2DIE12hXpEkFGd9D2ibzK3n4vfllcGO2O
ur4ELATRisuv6BCWX0yobtce200ke64oqiNP5gI4q0qfHXC5D1F3JBFzNonozAki
e4yAahYylzYyOb95rTxQP2FrUSeSPnG5ih6HCH6As4migdA7FhJ0KD/87daxtcL6
mS+V9rwWB+xH5xMexqhC4+m63tDeT8ByzBJywQm5PR95jgIsKeDv96GfPJQquWvh
2Q2c+UrvTYjmECzoy8qBDMuwMvmcBxapj9oHHyfieA8TxTUqVB4AWeBgdb6Ms4Zn
4EKHzDBJlnTjokpawhKDE+FuaM0y1wrUgZbfbWsXN/P0jQOkvRq+sScp8O2265Nt
VceURvu3SxFnPeTY/4ir3ROIouOJOqFLZYRgG6ZQkxhhg93ZVV7LyYPaKUioUYPI
JywUFM9btXSgVw9dcZi/jhLR1dvcu6DP2zYXf11S2r+ZQ/1vqZJZ4IAKFfbfPozO
mLMYMHtk5o6awfehotpOf93ISDEiwqQPtwwnpiFLRpAK9/UUqBtSq15BU6h1MK4F
E7q0n7wOlnpdX7u1uW3Shqm/c15iGlhE4yOOrA/wFBFTaGZkppmpJPBf6GVch6Tc
NqDcmeGzP9sF/VmJ/LvC5z1HJrXa75VSbzz4A2dGdWn4iiNmCfBsgqk0V20AAq5z
7zsTmkYPwmnb6f3YoyL44kk4/wkH7HRTEGxnEC93UOcgTV45uU/R0LVUye7UviSU
cO+c/G017X3rMGZhzeYTv2Kh7qrdkbZti6i6GNQTiNivGdfKdhNFg90ivBo1wPtM
sGPTlwh6rBMEU7UTQLZiUtkUFagK5n6wDIbknzADy4Q6a2LHlJFiys7dWqdXRm7b
c3K2nzeAzwCwenp2FE45TMIWdqrSudb4H9zaJ6E5ebczMq+cot+0GfX0ZAz/m8wP
+M5fPNDdD6ogonD5WKNnImapa749K8jYNct/uSdJ7A7dqv///xNPmtFdg2MhBI79
+359VIy3sORBacq7PGyAfsyuqyTo3dNJnrgdG4/qYwDNBpxmPiUvZ1iDgWU+AJnx
0tFyGcDHJK8Y39bXj5zbUCZjh0/A3tp4E7YxhTUCG+XU2kolEybVvbhcV814pXIT
tZruRMyj46ADADkVmQH2ewSWu00tC3C0kfCv10cW3pq637KpNy2HiT30XJrPvGja
0baWzhDLnIPkF6fcFNeH17PWpPSRPALIPgp694GeXNR85TlP0TLAK1206HF8CG6W
owMtBvCn/zqqKj7OvEXaTRmQSitpNa6jGqBRg43fQ+e3jkMlFhMcK34Q+cgOiP1b
KN+INGRPwa70hgFGhz2MAaIJD8pw0wQ517wp2qkUriGcF6QOg2H8F+/tt4YRSr5x
wBjkwZPfbBHVUNzLouvnCy3UTp3zxd0GlS7Z+OD8GSAFv8ADjX5qsFFyKjm0gHwJ
MLdl0pdUyvwrDGkPYUl7kmbTic9+cgU2Kmm7ST8A5ZAVD80RiVm+bHxJctxLCwap
uXdaN4QC5b6d/HOtmNYMmxxoJjRbSigU0Py6O/qCCWUW8uz4hUm6n2bsJYnnu6hX
mq70jT7lYTDhs3I6HGbUEDaXI9viqnI1jX8627yW9nSB8vB4jtKY0ybMVN0ZJTX7
R75eJZl6N6BPwAaea2hOdtWTEu/cArfIPtzHk6tWrTUoTEidLVEEr/nRdoGEKESM
8urm7UFEYhwOnee6It6PH5wemwpDL1l/Y07I5mHHkKyk3qFyLBGJGSdTxuVWGV9T
uGaL/GnLr1LYFLQJhb6sRqKpx8LK/mupAbC2XhfgI8cSxtDaklwfAbKURDNTE/wT
T7peV7P/7xjFqtovkyhqK8EQr2lMvWBoHFC5dP94//wY8vvrwc1jQztfEN5Mx+/g
Fsb1Vh1z/R7kJLufoJD1Ne2E3BG/hkJmV6TPBvMb7FB4zE7TL0RwWVTEEX5a51Mz
Xrm9KqN7S8MLzQDuelEv18QP3npvP3PftAaUn/cg3aJbYtamvhF+NpoUOhPMxdP9
7haARnmgmd8ENCcDDVaIdKixPe/Efy33t/O3Z6dfBA6r+vihbEy9dnAEWPKuPZ9m
bmNh0aX6tcYZK1lTTa8U8DQkV4mMn22OnnjaFeJFFj+KPaD9YiOhZtubg8DaY8kk
qvU2RlNBPRnBiK7en6JgJT/579nlBhfCmWQSHS2RZIPVNxTTrpQicJf7NhIl893i
Yw7VKy6d9EopY9/U5sgiu5dmKgwsYHYxejLMuDy+G0T58kWPD44Tz5v27673tliu
qac8+ex/jPibaq9sd6lVEoMj9HdvVSE/Jwql/W6rDB9j4y4uQHy0J5VUBgpJFHdx
9cG9xrDF3mRL0+BZdP3kQX4aoaNaVrnzH6HN6ngWfGTc/NGmHoX3DgWeTqLFD7tP
vRv1+dR1iMMXaOns6e8WOG6ZKYeFcwhBhNcUdP1WvI5FjBN6an54/UEW+24Lgs99
lb3xfZ+GAvojRSWu0aNbEUcayrlTEiWVpQYloMDVAhMBVQKvtXxc7O+BczViRM8I
2HmDUF1A3vaP7eKKtmFOEL/X0P1ln6Ic27elNwMm/JnoFzUYcP1TUy8zHcj5EfnA
0L54H3T3uEKr80GmM8XPdNWhEWKhjG6gOe7kV2FJbDjAO8VC0W2WxUSx/mbioots
RJfg0Ikl5I3YzbVt09NwT7wannGWATtoF3F9ancby0mWCr2DwDGcsaBPeQqTLZbo
BPEUhgvPc0uCj27hUhnoMmWPu9ND6n224zcX6Av17tsxGoKHaxGh8H4tmuKwZdCv
YdZmFY5ErtRN48NbT25MydEsMmXOe+VoII1NSeNdXhilwUyt0awFXdgiwV61/L0D
/inPHf0EQAmNanv0p7JiB2rmXyvRO0VYrjlitRKS2edC/bfJmgQFGsBYfuoRN5iA
VfMakU2kElYW8uGOtLWS+ZrqIKzoHekB0ZDUeRwXXSJ4lx3uCNIogLuiPWIY4M55
qMU2wF5URJWdbDo5WrXAcy7BoGPqQBaz3dCyC7raSP4SZVD3UU8dZ2SyZU6lrfDr
TwbOiWs/POo4145lOW+qiLKR7DYZ9iN4OIwgwoKIFY6taiAObAgVNLTs9wBOpXyH
XH8bvMSQNqX6J3X9ARUFbnmkaEucPUStaJH+MDC84TlrlJDterwDHP0qpJkJUypO
kt2t6YmGOgvoxxKO2zuOunUjVOqcyyQETJsFYQg7Am8BKohXUwnb7KRQrz2aeEri
QZBdczfmZvzsJa7+wo+iIdUwpSHYKTV5VtQsyE2I2Zx9nfZM9cLX0Py0EOBAMmhz
e3jv64VHUyq5kWZOH0wj6847WGmaZC+ku+uckGuLPqaEYzwqgEt7458lauRVDmk8
NSgy7tlGOWTrr4Ev0/EFDZCy2HG84V8s+elP0dagVkoYxuoLDxaSLckKdI590xwK
GLxwEAoC6/eDIbmraBHu94Aq/ZXQ0M6ACRrikc7Sfl9i3dDQswZvBn2vsjfXxPwu
4tDtAB/I4bqY+awwpFfzzzZie9l36ut+jNuwB86ygE/ne/cF5CMCsJPNiTaNI7rU
XGjii9M0TfwA1Xf/31MIQg2AezaAtrbdBnvGUsTBCHUQz5/5ujiIInWkmU4yRazh
P+EWUM+/UMjV+rxlDFjmrHHDbI0Ko4kylvTWLkm9WqAfM4lq2Zufg3BfiTslUPWc
Esk3WuhDRTsT+LJiy9NoVpgpxNeLrkA6bRlnc/6S/T/h4SBkmyDwQlg6Ii476GyC
li1qaLCPxT7B5c/jO44N18/AGCyGdsaaFxT/Q0JXm+Atp4NQVPEixnmNOQBHO/7O
QpQOb2XQf+5yiHagl8mE0MUBxfo7ReU+lK0PGAEIwUOmgjwgksW0LL3xTWxAzoJb
sr2zu9YFyiBB+C3+zkem5j/If06KWTPFs/pio5aP2cDUaLQo8ItSczUApqirwesS
xBMEyqEyRhH6x706GboGavJ//2bf87Q1JmCm4vyO36jvRfVLUpUXdqeMJfy5p0yv
uXnrzYBuKebFxHgjct3iNPZMZYWaZB9CyCN/DESEEoiD589PLOL8nhW94bV6wJXd
d2M+Y1lU/XDP89YG0EW5g7O87mtiqVfRr6hAqBg6dgrCNGx2eZBy+OxowAN1rv/7
nxzq6z3IjVuLZBf3nq21wSPHOuRl5Z2BlFBpyA9sl9YgxlJ7N4SAklDwPaF6ooSn
3O8ELfE2hizTR115Z8qk/1+KKxrhMah7CXvVf/tY9PQc6Gxtg1ctdZnmdNV2RaCm
8H8nhfre3VKvLM4T7AygMMxJ6YRQyPad43tek6QT663TNgGeNC693uiK/t8LKczo
PIIQ5zUdmfBj33tiqEvMwmg6QuexevCwdiucAvJ9KKIXXFftUaZfBPsq4JHSj1/c
kBtnOSEcfDJWSG9AsKhVkZAacuPqhwCMY2F4b1rbe9pdFxH9BY0B+Grl52aINvJc
yXmpDQ3HO+kAkqMn/yL/yKBXOwuMHPusQjamZxs6suTOWKt3DIUTrpeLl9rCgdRk
gCQ3tFeZUItKfixBMbpBT2JezGp63hZT28O4Oh/Wlnas3Y71ZJgGawtxYyPR2x0G
BARPtSwpGNZbtIhy1VUD6J1WvCYCk+vtSis+V6QRu0xAGOcxX6Pc+gXR9w4K0Pe8
nW9qPIBoACVGUSIPux3gy5Cr0skF8K1vLaiXE3J2ah8VYzvh7Qf+wO9Rfvp0Y/fI
b0ehUwBBSK6EUzW3BWl9XjEVnF3FwSiDjbqBoGtZ9qrOymVQnvpeeKJgi0HJ6UgQ
Asi+ii8wxxkQ7eLqIolcVQoTWC+tVKn1DWRhHBh+RsHol6ctCg3+jCTwgh9duHif
0RXW7YjuaF+WHFq8usbVhvbgMVVJGBp8x8DKd1cZGQdc6WpXNFM4TDxVPytPYBF/
IQP6urncfO5akCShJFpKG6diSsR/dOHsUZi+5CPmK7qUFdQxCWmeXOELbBqRyayN
YEb3rI41JH7r7Pz1NpDLGhahf3wES9gBZme4ApoQnlCIrchs4BFJHoR3Ct0TqmgR
jSIFU36CC5Hik118oB6IkOsomP1S4+rGgkg92BruCWWoK6vebKRaQScNvaNcrpH+
E9kbHhoYsJn1wJegqkv7KXJRjkBpJFy1YSSogl6nWdF+bboQUWdWm+6QYYMDF0RN
pnFP92i0dacDekv9OswmjdBbPtzqSOWQnSaQc2xBJXfIRr8z8bLzP4X0zvL0j6XX
ZQ2wGulPwp9WOiwFsMEbHagyUfXvjAmyJkK80XTDb8za41eg1JiqvzOSuZqJic8d
+0lTLescg8NAdhCHZmqXki88nqRoeCgD4jDx7zXTF29vOwm8pfKwJB/FtoGOW97l
ZiXUDUggIzPCYK40EyGqcL+7b2fa35RDtt2OU0RZNFNZ7Tagtf5zjkjcKXMPNg5G
93UpscSxji0oxISCuWmStWwDJM/sCMBaBY3Bzc07WhrtvZspkKHveSYp7PlT4010
vM5VWasCAlir1dRkoZJac6lz1Bjf9pOpaYgdtLXi9ie8QmCdCEZh2u/wz6WtDZPt
/GFgb5CWHfp2QI5lBd8IbNZpXXV99QYPgPig5BW2qV6phez6NPlok9FP/jPR//fP
ZyfUQd71+4NPmjHRRfZJwhrfun/9zKQ+gCnmw1tYCBuNy7zH2mVjOBnThX1ZvM4R
NVWPZ5TSHe3wnWHPNsCZn2jzfgWN4kD5MTehSq6IOKEeOMzOJU8Ns+ZrjTZAaipX
KBI12I91CeANJPrIgkMdJnH7Aj5rurBzIOeg7FAqznFMo11/4hj750U9jo0p1rHI
47luW+zBmfe1pMTO4zLD0RyI96zNLxWbe1tc9zoMKMkEKwacwlFCXdJZ8KFqJDfM
gxnMJz1Rc+TZG/UXESi/yIR6wkKTOGpCozjQH3fI4losb3j8gnC7loG91oTpJTi7
NqNSiZPfUJT3H4mPyWPKLQV4C/oXJ37VAYsUMUrJEOALJzBguS5GtUW0BWx94GzY
BnV7vtVmgkmH7j5NG032EBO3QwFEhMKD5rUWrhLHC5y2o7KEiI3qihDWNp3+4Jos
MEmseU2yXMbzskfxETtNmhCqI1JmGpAt1mqJH8/80PiODsYGFY+eXhekTWPZsQCs
pD1faqeRYWSpsC0RRAYUXuUfFr2pie6y9ATj6lC5F5ta58s5ug2gv+DnGcgqlb9h
C65CByrh3oasmlqsVnW/yYiVjoT42RP/4UUlyEmQ7CZ4XSrknan2fRWFePD1IvvO
JioiVJc0MKeIIE33fRIlOeYpPaSGyARJ0Qp2VlH7lj8vWdYGkbYxfanMcRpPzyu3
Bgo26Y/GD3RSaNrzMVGwSec9SHdCcmQC93XHp8AbFzNbbNS6kuBFznmgMLoyNMM3
FsUJOjsACz4zLxcbBZ7kOD2hBwNTT2LGt+t1bgyy5kklojjEjsV+soEEqp6fJvvZ
Wu6CyiIafgaF1FnrFM+VDiQ9h+ScRT8655hhHSNmpkwA6q5Ivu720v63JsrXQI1/
6EyTiBLlVdAymjMNo1s6K4Y186pYvHnITC3P+Y/mJ5pFjw7lH5/d8IL9JJzQsCN+
lHzZ0+Tvd1OfcpdonLVPPRcyBOad28pSKp0mtfCu4rC+/B8aOmNpm4yt25d6ln1e
Ggv6ia5zu0hLN1Z+HeZ+UKzMJOe1hloYhl0McCCCVPVH5L9leFL43CrVkByYyv0m
sJs8pBGzpvzRjIw0JLpQebgxqGoPUTNdo5bgvYDPQWEno4OyP2wrccWQsb4UqU2z
Wrc9oL4QFZyZGL2vq/J3ba9tZFPNAJYF/o1QbeKPX3W6piABCzdE0LbfQWmNagRG
1J4QVxAz86+0IufnX/VdxDyDpq/mnf5oKm8eV2d2q7+2dgwk6o31of/fiE6RZZOP
aNNHTWMUtw1X4HBe9ZpyPzzYc25v/dMGxr/U21m2pFg+X3D5Ghu60uF/8qC6mlle
9CRGJ1yanWQ5WV9KiuH6Oh2ULa6hB8bwZc9tD0IHI9hMAdMZwGkaDF+vhKBeCjT6
kxzWMPGS0oJVtBq5dknFLfd+JRanBfLDgvWB4mpnMmEiKSxQ0/b7flwORH/MM4vS
zt7I5QJ6OtQN2xprdDEG6DlpyQGesWlpNJvyY6hDtXbsOn+bEkPz739G8lqkIAfQ
MoKMLa7OXxeq3SezF7nj4XboVJsMOMur86x6mm6XcK6QU8BxfUfUQKyevMrqnZRW
EeJtd5euII253RcMtpC1yObV3c4uuWFypvffTnZ2jqjgnHwzt8EKB3qHPA8bG15Y
zRAF/OxxVMZpZkfCOzabTDGLzhnvN2zQV2TEMgsDVI1/hGKYMCnL8FOnFXOv36r5
s+g33Uf0bIlAxIhLnnxPZgqMc52k3KYPHuJLMAjYBMAjUIuLgQgVR0QBpzpTBSlm
M7rmaaRZyv2ZN5k9ztsdCil+l1tdw8Yesm6C02ATJMjJ5tr715+7XyWocQXJ//ZL
41duz9rWH2rEfol4i/0HbLFEiKiKoAwl6taT0TA+tcRAFZijonADuHLMsFdiwTbp
/lxfgU2Z1igp0Q05ASQKmGip4v/L+nr1jFEHrh0pGb/z2pdCEs5XjgKDNySJHeNU
F/CD+UDUnCbelzXYA7usa2LB3fvQWcC7mg0lkOiB9ZCL3UeK0iNadVAr9Z2sYGMh
hMaKcZctN6G2eEnHwIYR8BcUU8JMTMFBEiWKDOvEEauZx153aFzvHVlSkZMtJFz2
d/iGdF/ecyvF84ZhX4aCb/tk0jTk+Q/1IpkooD3zOthMO9Y6/iV1FVDzYOQWoT+8
9IkCUHvUtdEJB46ZoHrYlLrtouftRN9ytqKrHcz/G6DkGokw/g6C+f/lyRGRC79M
/p6v22dAIhpQrNiLNKcNo3iOgLkJWqpjR34nxqsONJqqhbp+kph8OmuvT8glYJwg
bFF4H3TuSfxDQ7PNV+jP80AOSJu/aFLcP451jgRO4WnVURA/cSL2uDtMWXVaL6l3
7Un6CBBJutWhyItcn3kKqYuzGYMnmtaNuRx16dNJdC5p1hMLYHvh3x6kdp9KLNmt
0cvne4MaRxtlzw8LMqLB+KNDb5+Rer+s+IlaUmbHoe7tTO+5Gh3TkplU5sXRQzBb
fwPuvz3vDbM6DlJ83LIKiRe++mWtpADTYRJQIQHN3m5wEdL9PiG7KZrYP4SEg1ua
Gxm02+E3jXXfre9l6VyQq5lb24/RGz46DJO11NySpBjUgttI82pfscT2Ww/7xX74
s4+S0vCtCPXEotwF2QUOmd9BJRZRcrTBNcAMIagDdoSx7Ujovjf7r4Hbh0NMNfJy
2O30ew7yp+VpbCqKgJH3cL7Hq7P8hY8H3/wB6ZvG823LglJ75jnpf75ylw5jonTH
XUzyUHjVKc1FMH/Wl6v+YABmlS6Grr6gFxXO9rWDdZHuqrChHc9ytJcj2/1hoCnQ
YLrpgFclRavU8514XuKhmBpkj/I3oMZJGFLuuJY3m79IimyaGfGqTjJpmrn8UDT1
BqqqJ4GZOAT5Ppp2xxLpB1riJKaQ4kXP199jjTcNBFeVViJ9LpX78vPuYY92UvQj
PAX/kgrUPuIt4qFdNV86rbVAL5mZuGgGVusr78GTV2eoZPFg9A8fkUh4AfU09XhV
XCVxje7piB/tuTyieq9sbE5DyYM8yUFAt19MfClnmO+5ncmXkjHphMSsPHOwGFzU
I4kcDOtpRuQHYzQXzPvVSmuXg3cDbDN4+QSs/g+kY1ht49//sDiG2DPRTNAsosvt
w66BKnWlioiwfeklunHJqCspm09tolIiAKeOfjwTUoOoq9o7XaTub0vA7W1gdn1P
5R/nZOAj5gF3w5vK+9qs6v4lgS6CWXxTFgoDd6b2hHVTr/hxktg5/3fwg7zYgz0/
MieCZBxMuU+lqh2LV01eiUsueagCgHj72zYC9lKRDiChaCH5gpmS9MfUvGXP32Sj
aYqTZkZ7B5ldOg166sS/PWuQ/KchvzPWm26lS6FItctXEJ8ffM1zAQQQf1hh8eXa
gO7bUlMORdDZko8eCPxsyWA62idrO3JMv7nwGyjPcDnuPbErRDBjm6uvv9IGLV91
sPbZV5hRP7fp+TXhWl6/If5ZuQn1VDZ5yC7xErgiz5hCLabuGJD3PV9+5yIcjLPx
ex1ybUdrfUHzOqPeek3ZEJhF4T9o7raSLMXig5hJKuS/dst8qG35WvNdCTndWjic
/ou+WiGUfFhRVa7kMyyzVb3K3H877KaRl8JqEp+yAIIoh0FE++Wo8UmVWiTmLvWV
LnYJyrEtFZBwm2x1BZqZWUrOHate+yU+3C8Fm+KMALCk6Vi26Yt/iSUGWrNGRlO2
sWPlLzN11pb5KvLJX1Cjg92hBmfLwJPzdfol8Mkzj2pCKB8Z7C7x/tOnIPMdNTRD
KGQFYhfvZ1xeReOn9zfw0fSKWjfrUczbQlTc0We1WELvwgKiJAIGiTmOCbcjiSL5
VE8gmiUYmFBBE9jpPhoP6NaZpCL2hsuEEGaeRdJxPWLKyQY9yEqyDDTnC9wdlRa6
eNyE6XZxz1GYEExMcHYsPwdw7cEZCpB9nfhFcRuQ63BuN3QeTQn8aJE5Pu/eB6lv
WNsB4I/nhk6GraWPsrspQ2uu1BVjzAPJNLVgWHm1Qqb87Xrssfhu0Ez2K1/3zda7
p11mEr1TDs+CNjfMZwq37Xt9gKJ+b6A0BbbcySF6w+tlHkpc9ypddbackqGpikA7
B1Pne8AGzI8p6VVeWu+MqEYEf4kqAliYE416LzY9yq29QwLK9Rwy65429N/8prQO
1ETLfw5hGwhwrN3mZpFYmyvBKaHlkjnwgVaFIZxkSHF/2W4hP347LTVt/3iJag4/
fJqB8lbu+rdylqHxesg+YECdmUOcfscgf/IrZUSilcknYB3i70ze+e97Gn2FhP6m
h2o+kck2vo21P3oFJEQTq6H3l5mItWiO+G1mg9U8a3QYl1c5Zm7FfXnbIZ5toRXG
I0kVquL2Mg7WUgfqDDpo6fiqmEJnkVGMelGccpysDy/ulaBFSyXHYvbtqBO8N9dG
snTk5fTYhScpo8Oyra8RBNubJfN8jAH7Ck8Cf65gNWIpPiXp2iU56Fd1TRFxDR8l
FPfEIxXHp0LdCKcXnWBw6BpCqjOiPenFJ2Fd9hJOj154C+xlSvmGpS09RaA12JUe
4jbNvKpS6lJqb1FDXa5bJmtCX0lNToNRSmiIba2O9o0p4pDJkvPeL+9Mcg9vjmhi
67jQlmtlb1IfeVG/hGdjXrOBH4qGhYPIwwug5p9ww8ABUtJMqBPs7k63dzulW3H6
l+knD9uO4fsiAYTPqH7ATR+uR8cwKz4t0IXcKXtZ1RNPF3/Hsjclyw1L0rEfsMuZ
/66ccZb3OLKM4VeYVLZCjjItyV3tvEERLEF9Zw2a6eLD0TFABjIgI5dAI8sESzx9
hKaFURYp9K66Tdcpzu0kwe+Wq3DEr45hPp74xzfUSBDA6qRbD9YKg1K8gIbZqa8X
M+smkNkotS31OlusS+aCbAJ4/TabQgHlcA6QmANrggMWyUkmokMLAD+X7vjo1TLH
yr+vCiDNq7pd00wBn+jVrZOQB2e6nVj2Xk3dx94BAhJhfryr6RfzOKm/7Nhe/8Ni
IfJNxeDrshg2a82mGm+5StQCfws52HhRNP+D69wu/caruwRVrD/TvLv6tNIck7lP
5HK4HMNSFIWESqgoCH1o9RD6jBESpPgE75A4y6io/42VzgEUP4h+4CbHlbFYocdO
rMA0WNE4A8iVV+3VX8s8mHERVYl/zA17h9Uz4BkLMJ+2oQHHhT55tAZtBlwv8js7
eXfphBpAYcxUCKGI/+THOzqk4DCuAVeN2WW+XDmZwygS2LiYxbgHxm6oeGZvYlQ2
K7CP6fxxuoyaegcetABE1BBqG2nQANCHIXbnqwm4F5y7+gv2Jr9WDCJU58jTGOVa
/lP0TebWyzo+6sjs9fotXaHHtYqWrUs3Dp2gfyNAM1RpabF6AexF7kKeEO5S6z+U
T8CC2Uy0TevBbqbfhibwMaDVRv9S35FNHiEP/vHx0iOXNNK/xctLs//HSDnU4IWY
RoBrnZoYI08KHLUHlQtmhQ+2LTJm51mdQ1H7WrLiYPSGjlZqR7BtlObgdBFc+16o
aCIohqkOIOjsF3pZJj7cjYquoXjbyuNFvSfhcmDa7qGFf3OoOj41S5XE3JrZKjRw
C9N5/1lqMjbBqcTRRnOZO5BxfiCbB+CEzavf2JDgdoRa4ovAC4h6mJK34YdbZhUT
xvCVl9BzWC2O07EOHAteMnHS5Ty43t9pWXZTriiczE+lC2sebYgUkpSAfpm6RIhF
Mu+nATWVLbpg23oScgLCkt+juoCNEXObNeCsrjB2LsMMstAppCqZzpiBI2zDdZkw
Z2cy/MBKKxQct8zXFEoP6ULmA0W8YUoref4qGOxWRQ8oMYwB7Bg7o46Gh+PEJayY
8ZLPNtVlZ4O8hpFpKd36ll3L2XC/3BHJGWbc5Jy4rQy/858M+9Y0Af9uuFt3Zs+4
ZpkgyXBSGWil+rURYAmyXBQX049+Dfqr1IbJL8NUTVVsJhfXysNzzpGC/ojcC20c
fHtJp0pDD8okySNstWw2KpUX3oLQ/dFPWXR2/rrxGfaAEMUez/rKnAtDbI8akpyJ
TChesomcsl2WpklwKZAvAIX9Vtt2XwutGy/oI4FRfDo/U+fnjS4Abq32ft2BD5Xk
ID2H+8lXnvp02c5TYDJzMUjASfiilcTEYg1RRua6r0oBi1AQwHktW8tHX2FC9/qd
eICNNscFxFdevoIPx763IrBOlCJ/K5A5k2soJ5iemFq4VZWJWdZuf9wXmOVoLYI2
2hZI/9E9H/3IrtUKoRHvHQgLqak8pRhFXd2IL9W/MJuBbvR7PFjAhihr4yuQzl5g
NVteeaNeIfBvx8Z5W+aKJOuM0ba4+z5iYKrXstnrbXcZeUVzA1XNiEOBtjz/Y+Fd
EOHC/EcO6kZ8jvots0lAd6JkIy6V51StsJebPv09e5i56X2qRcIsIGZOgHvBMGKo
3mGN2tI+UfW5EI6vNx0rHFQSBVX+BfxHVzSYPkT0QTOfLQIk+S9/LfgbjTmQgdob
T5f1FQbJHWhEBgjv4fxxnI8fDQTg2IdKMRJNg0MEMIy4sCJXnZvgO2zVOjVFOERX
svqf/5TNOsz3rzvRLZIxdvWwbIU5WoKLMRtOVvA+Uz9QpLehFMfRJB2XtRpzWZ/t
p4gaya8yfSPNzHypKNsIc+wKLNMcvXaTyloV5kCyWHdw2ovgJADUWaEB7Rc3UQ0w
7ON3iMDsMXdnMPOKXpLlwvVxyHP/hG3xarUye7rxeRrC4KG+bs4r28+tFt5krwSC
kf+jN/u3cQJpEIOHVrvMNo4yyss/Qi1tP1WsLWvr5QagXQXr+m0JIMCE1gQRLzt1
XIX+7q8Ztx0Qf6HC8jV1c8joq5ocMVmJvO7VkCi7Web1iTnLK7VlKGLS1mz9Tn1a
djHEbRdg74awj9jaFUZC3DJZ4arjlLXB0exA4A0QAci28Uqhpy5jITROE7EhpAsY
dMFWL49aLI684sSDHzYGXkrn3xxKsiwiWQUhKjon1LFMNPZt1FNkWK25XezJkM+t
EQZ6eKEwcOhLLEoDc/GjpmoCmyxPnx0IyGWPVC/AUlF9PjhM+fo9uRwtjQO4VMFO
qkrZeSFb6Q1nGCJXaWtXHPCBrFT2qVFpll3T/yc03GSW+hBl0y+5fnFXx2X7J+0O
ylxDu8WTOppqx2s/EMTQAEzTBhlJNIMiJFpcVvcmAnRRzqMtsI2S+xK8J8ZIOMno
FbSBg8Mqa5ImYgNCIkqRVWbmY7Q/ZOjjj2mzIQ8l0v+kM/b18h/wDVTe2Uq0Q0JV
hBUq4pjwRI+TyW2/shg9RiuLsNed9tapj1LiAfxfkDOLSw/cM3vK5g+uZS03xe7D
6LZAZp7HcIx+EsP6eWl7weE48XQRofwbJ8Z/OzTW7tMLG+xy98Hr1MGLWoXcXE/D
Le0hdQynXXoSHGgGP9EDluBZT2LIi8NH9rvp7Xoj/J8Zu4Y4K+4NlG8zhyC3t4Vo
gQ/Z0cc7rasfgzrthuF5dbWR4e6LZTXpR0RF6RwWJavifkm8okEwOEVJ84dnz/UB
+wrbf2m0Ggmd3umIKtBCcPAQcwUEVstykDnWRd6qssjcH8AFBPYroGi4FaJ41JLN
+dHyBrg38HMzmktIJygyQdB4AJy9DM98zm4bT/215ZRClR5IYnXbMac358UCfgHa
nDy1ni1NhIjbfEpSD1BTz044GaMX7rJjV2msqsb45+AxQieCZmkTWVu/Nb8ZExZU
II3oCjDYQfVoyrGacYa4O5GHlTpAVHuNMJisFcdpYF/NYd+/KzoyQ96B8Ca58YcU
zaBwS7lfZ1W5tTgUyOEfJZi5vp2pp7f6PUqS9VB9bUXwmuzqKcAqCW1HibsR4W1P
9rolKjt1bD6xJzvMpS/BMFEAVuA+AXBOUxN5P4Rgpq1OqoWrgQC7eCc/yi0eJTBm
O6NBLKvF+gx8VUmfhun+ntsM1j6KAbUM490ABe3Bo1m8+xAs3ZKyTaviT59MHkbm
GNj0szEyNs0GFYwNli7GKsM6CHxnuyU8P0PBYO2I0SgNEA9AaaBChYTNLi14KTpU
Go2jztowMz8Msv5wGzxM5f/GTsChxikIe8OYjeHgilpfn1AiynpLqkgLem9LBO/o
0gzZSFMFiJRu6Rq86egnamdMUlHETlX9zBiiYymd+fORUkjqwvtgkU9ZE6GH/JTm
fEQQWnSC2gV05c0zjiFbDZtokuSMiKFvFgjVr2jg5KBZTescFnHRCcFiNnNMNS1S
tTqSdm5dUCz9p4SRtOPwyCkPdXzJghcCtusfJbmYJmuoqfou3SE/mxwBIcD0SpLw
ean6LjavlMMG5e/HD5kqhTEA0coCl2ulxK57cOh5Qmby+Kl1jtlDD0nQ5I6Kbzv+
H38WyJ5YQBIaQg055H/uEybU+YmmCoo7dTACY99QyIz544iSUgl0u/A3gSCj9A1M
10FvzO32EbcsD/COQy2mEM8wwd9cvzOqRFLcQgVcvkhlGEbukk6bAm4QODu/C/Le
K/UkoBffcB4WEVG6MyRtgls/dYGm1VGqBZ89YAfqijjlTQ/B0xEok4CZQeVv/s0P
wjxR3v1wwgWXqib6QLM7FOCfw83sXZLu7qxCv/tv8V2+FHVqmQdD14F3icb0kcHz
52Gt5x9P4QGdk2NKVz562BKo8hQg2iD1+yH3mruE478SOtNYl9Y5hwlTVi/jERsf
hu/+7KzNfRVMPWNVF/tXUh19RIzK7Yz/gCqPcYZYMdbDIUYYzEe+jrFnLIStmGSz
9vRXInM+ke/jLnqquiNbL+PpnL4kvdYc9kPBhdrjjVwV6c19pHpsxNDn5vMSg6Ml
I6rm8yWl2AJkpC9byu7icpKpvnDtB152SVPLjbjYvRifIqv1khnaiLNyS7i2zSdU
g/EzrUwwWeoO4IbY6gzz4zLl1vA+4J6pZ9sE35feLXS92ieuLL7FuLKPh3cD+gUU
LXqhJf4po8GhCnK5VaHoaqQwnBYCHGTA0DiT+mgJHohqG+CRLPhYiZJaRDyY8VkV
VxXNBQvEnGLJepfuP43XGv7kuqBKpMr1I4yLoAEK4oRcrjNjJV2FwEn0AC4qTjIr
p67qc+mVfD8EFdPGPxeX+Yx5ApTRGkF+6ZUkU5BZNVcEAAHdOJ3ihj53Ja4LZA5q
uptaUq1oVQ+WXwNAn+A7x7LiqHL5MOQ5V6CuYl95NxfOSfU5bWq4tvnaxJUSZpJJ
FaLakiHER2T0S/fxGll82Q0NmjAaMo60LBS5gpPD1gFHpxhkV4HYeZzjCpytUh0W
ju2OP201gfSZba1xhouq3tAb5fp9jK+zCe5NifBmBxjYsJOj1nJKlsc4OZ16prEL
e3OR0dNLdYQsh4331wHbCFwsllHJhCmGnfbgqZb4odbgl9sQPsiUPpBsX0PmqyWf
PzA/NzRlqkp0iGkz0+MZB0a65wXrFb0EbKXctRGX12a8QnurDs+YbKCEmqT2mQ8z
tU0E6dVw6LTzYLsLmWil8nnwAcD8ajywTDK8olNStR4JC0KRFJGopu8QEpCWNcUp
u+D1nIJymobpG6xBC/+2dxNbz0UCRN0vB1GsQqF93m/g9gm0DQ46yZVwJpQpmAtq
w+6Jrc9ij+5UUqy1LoSKu7dLNU2iza9biH7DreVbKwcOC3vh11raj5ZTMROiZo3P
UmGwR71MJyDqI+dw93qjWJW83ZC3XsfNDevh1f/7Y+uB1p3ZsJygIquqFulPubr8
ymIgIYlsoac777NGYDJQlUsxi6NeIfSiq5LAITLIAG85cHwq1kQB+Wh++bOS8Ius
5x9KygE278qVG1+4r8ctatkefSrItHCwNdcx6JLlAyrKL06Bp8adjgsCjQTfpr9f
qZyx+IqoVgF8nbvsPWXD0kfXPSfHRZzIfbh9NiHBlxpvemUSrZXRgjBpqY4Y89dz
XrtSwhRnSeGd3q0Ycs53M2ZLAAUv/rzzqw13U9LGio/1Yj6/6PtaRxZuu5lQUCkB
hRXPIa9EONHjIavcfwtYoVH2eHzpBxvSAKtobBerIGzwQJIK3phYpynHd6nvxHwt
7arPw85xxwvr4MwpTZk8yyxr1lqxAnef7QBhU7QOS3PWOOASR3gCRJ+7CvAHibqY
qXLewfxBqahZL5RDzZ6c2P4tNrI1q0SyowMgKYbrSrkedOCOuwwJiugHLwfrnNcX
z8jDJM4acut+sFlUVHuinaRQGF6k1Ly0FSCV/4hSUF1GQMMMaabG+HmUA/YLLPst
zN0NaBKK++TfWMN23DSuuC/rJ2msSiSqrVlVJ/CBjAZMd2bU8OGfpokmapVBtiJM
8gGIqMVcoYFgKWE1SsoF+U1yLUJTHsCY5EZxvk1RcGoSG/xNiqn4MX6p6Yoqaxja
xy4bVLF1OIFg74Mjwnz8jQH+jhzr5HyL/g7kInZytNzx0pEejNK8w2EavVpkhDWq
7Glp0Qvc0dNipVDZqrbUxNo7mWNslXE/2dNL9qkZCXH1BojH8UeQmKaMfKKK/qJI
`protect END_PROTECTED
