`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cyk6q7w9i2sKsYIp8Bq6jTGerJJDF4SBx7B/5TsvJGJalAwt/b71j4SJuB16mJDU
iq7KuFeETQhogbQJg0VIXZMQBopUfqrpSQwMLc9xCjBDYcmdMSL2H31YxctYZm7a
WeeYPWvHGoSvtn25B4Eb9dTy97Yw+1qv8dPjeYYmEwGN8qIUKvdcyRE+RnzG36aa
ql82a1ceN1T8dzLxTVrdiQasZgoObPOxwKSjd7+CqUXO1+ctJHPA7asQ6/kTFwVk
iO8/VvgxsSXrjNmFcbYyKFJ4IgbI4zJF1M4gGpt5j894IrRpPh98mAIakvqEITyk
cCvcM730AaapfmAyW+kD0FumRFXqR3kYpFiw2VOodV/Q/jeCWpFzHlWeF8rSrt8Z
P28+iBsdIchIQdqBd0pK83uOLVfwBVe8Bi+ADW/B6OEAcSVDBzJdq4t1x0TOrqMj
v2Mt7hB6ThSQaDo4qwsrB/ZPpYozYm/Y7YlrE68UL7XNgD3sTIPk/lxUhXcUhOWJ
orh5w0HfNywBORQEtTydLP1dy8a7GqfNoZkWny7KNMOthInELXOjt2IfB5HJtPhT
gi0GzH95kzf1WvbvyJuBvrGs6d/F2tlf/Tl4IN6aqQ3BivKeqo9k1VJEpebymWZs
A6Z9BCh36iaurFVyMESsIE1ivVccUv9+8UIbZLvlE5BoWb2lqpFoj33X/GM/RUh6
RXVJLARDQUXNY2d1AiSjTMIxN/4OygsoTQ/uC6qNlq+fa/5IwZrWxly8u0MB+bHn
0ooZ6G5bO6N3gTQUc9TiVAGQWbY8j+HgztculNv8md0lAv48wYhhSOLjGibIR2ou
enP3q+Ar8ddJn05asehz+qWv11pqcn2a9fQiG6CjvGnYBH6rEApRmhbKzihuh0YX
EQmvSlEClnfxoZETnvRog4z/jw0N++cRbOdy3vnBrCjTgxS5ARef7+D381N/Zqh4
CWk0dT2uJJLbWodRTuE+q5Uyu6s09dQ+SvbN/JHv2XPR15/LBJeTtVxQl/vWvpQC
O5DoBnyRHOKh2UXVN7nmPD6HQJYFh1M1QQFK+gABH0numKXYFQuiXETf+r1H1Vyy
`protect END_PROTECTED
