`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mf4Ru+18p8q6D+DIO0FB0b6J781YLS99XC4YBrtvL2j1YubtF2V3isj5nRDNTUTY
Vm4aYJny2eIhLEZBeBEpHJz7YSbA5Ti9SW5/EomqZc4RHyDTge1Q2QOU/mszORpV
uJipniidJUxJFUvocrkRgAsSKbQuec6YG42sLg7aQSQwmYEZHNv04Z/p+HRuxakA
SyQeBhCAe4ZsU7olZNBZbgnJ+YCbye7l2/B8P0amKvV3t5mOHj7lJXe9ObuDsTxR
dll9BkKOs9nukMrjDSwau/cym2n3RBjsT3NAaE7UAlhEDT2S7f0xOt35pkDCjbZ4
582yYiSs5Jx9fUHOSAwJrip50kaLDg9sVnce51I/yNX7NBrFTkY3wImk/siBVJHW
Wx57a2vHACJep0R7DdvEZHP+entqUohzfVAAbZB9F3ZYDRI4jaep7jlHxoj1kNJD
rcbBfhzJiDVIVmlpL9NPJ37hzSvKDzqDI42mVlwpN0+19AZC6ua2YAfaR1q+4wXT
Wm4QiUDPk08EeugEZjXtMPBJvx28B9RawWnyFZGyn3xOeCowCLGnm92/4I4QJ9cC
wjhFAD3N1xJ+jFwgzgWjo6LBk/Psgqb61/VB1FfamvMeXyYTgbj0EYxH7DT5m5ux
v1ccTNUn0zHY2P/VYWmWVe7WL+FoEPruuu1QlDutiMspJfKX54yGHnOjIedrfVLc
x0U2qR82XvWZ2fcFaIveDmV8dumj5vHWxel6zTLpA34xU6XabsrAA6JKwUGmQNE0
YU+b/UFMICWhmIUJZdT5s20617PceEEby7vg5FiCOML7e3FIfofMSECwF9599wiq
zLcqqMR8zvcttsf0DnLrDSMQevBCd2icx9oFAEcR6JzLfowWEDvpMHTMKT74PmGo
LQAwgMDBeBhDoNKdfwPtOwaHYiWDnw6hil1hiWms/rbagYaezBToJ8doD3YuDP+i
4H+vCCl2EZBEakgtij34vozbDEiPFYy5zuF0bbgnUne1B+/XWWc4atiMXEvM8P+7
OgSClGchQyVcTUPEVjMt0ZtIkpPpGLsD1FAh7BIxSpu2T4KXIGOKxnbmq3TqF7PU
0aU/1Fc5KU+ZjNfp3weolNyQ2KB0of62WbUJebwcusqwkFgeVPxiLqzPFJ696EWM
cHJGZDdt5H7+X53BRoT44oIcANrT20HfeDDl4Eqy6XVNsgnakf0qmOlpy9ZzPZfN
P4nyL3Xyjt8V4EjeH5bObXmtVszwnbA70uIHvu8MBH0kU37PdI1DVhWRwhi14AUb
JZCc4H715G4E76wxKkMs/j/sX+dy4IxoxZjmde2cUx/H82Lt4Uk8YXk1NBJ2uiWv
yTV7XxTQqAVebEvTTJQ+Uxh9uWcR8oAMwZmeaQQgqt8clVdKw7B+6NEx0AGX9YOm
pW8U0idrdUWky0u2MdrS2Hf4olg0nKXzmTElKkwPs1abp1kBW+FsXLCF3EiHL6Xp
mW4r7oTCZ2v4D4mwUE93QjL48nFVlxSGQDiDTZeJa90Um8JPcIJEE6tYtZz1TUGL
dMGHAQkof21UtXOnTvX5yv7g0VkZqRLpS+N21uxenN3tYNYHOm9CRSBA1Q2xpGeD
FSNJmM5t0mGjZAZOUTEUmhHToXUigeBL+pnN/Xgk9Tw30Y02dxTWHAsJ50DHiFvg
UrgD3xlmRZ24lJ51MQZr5CCGw6B9jxCkdSl7LQmj6VRDVjazW+TM9/pjztI0FhEv
tAxCCHgdFi8hi+qrDHascR2tiFsWW1to3mS4xoLklCOqzBGwxGCowtFB0z9jWAqR
`protect END_PROTECTED
