`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ivyu8yKq3Cdu1HNz0TwgBlUlYp6YKYgWwjF6R2AdDzZds/jYdK4l15txs4bKZAbE
DhCeXbAlWqQZox+YfOxkNCLDkbriznss7jC7yhNwpzUc7uCYPM0okXqtxI8iYYVN
sHtG5Mt1sRZcFv9KQafvvdwG5gFQHaAgBZID0IYatIXIMNAGQICS3W/bxHhBfMTR
SSwy5vpYuZ07NSpZYLDUCJ81Xe+80TjIJ1VvsWxtIwLBn/Is3i8hmJa60VkSImOD
qAetwsaiH3pNbvUemzo9DIy17juoH0d0ftXG6Os+aOe9y57PYaxvPC9yLhEzeUN3
XH5QFt0ZhmvydnDyYBk/8kSvVMm4c7lBulL8vDAzThEOsWGPUTREDvif6D/NsVst
y+GAo8uBS7xknm3X5wMlMhq6/5bs9KwTuUf4YH3ilVJrZMIkNYRfmZeJS0AOQ1IS
BeDKr4CRMxarRJZ/3W3837F+DwNNFuQM+UeMlrT9yTOcfgfNcDtrOwwOF6umYZrS
wpGTvlO/vED6hOc2gT5WfyVHp/0brJsBo2uWk5W6l4X8WZs1uK8Qkn35cTjxoryK
gyQI5SxQmZCZ/LAecV1b4UBKD9HwsPI9Z/y+t7xn9dEpGXzZyiicdps/fdC3ueYS
RcSSKH+JphzIcD6so8ZAgwtaiS0L9eGh0xTbs76Xp5MVzLuAN9bARmQP3b3LFHY4
Tv5QLuKLlsRLnQkIbztxsZB+2YKUo0KUn27IqikOXhtDbtGLnNDA+1B/1EcLdfjU
uB+l/M9rlFcYL4cFJBZrfPYyfMifQK14KirjhoIwMbn0TN8rrAvHPgiH0sVl8RjZ
DxkF77eDve8CLHyqDsyoMEThSsAq324R8iWqwSFaV4NPvt8Qo4LyGlS3F8nxRSeP
pR+uI8FNDQI2bGkJyXSBaYLZ8Jywo4T1Mu6YZ6/vG98EKmfGVX2RChPl/QbL1Muy
+1wlVc4T/TfnNKEUxlVx6l/6jKg+4fQYuPrqV3KVIRlffFTAC0H+eN0q/OE0zWxz
vbEFDi6DTJaUZfLF/XEmQY1qOHIyBhD9s0XEgKSbfBs+eKixDmrcovn7C8rZ0QeK
n1zrhrfUGZ3EGF3glC3iWPsd84PIAYS+Z8zegsIDveK5r9aAjtYwvULvqAMAJM9X
z8da2oy5aqFFl5IyfDuXGmnzLC1wpKT/djstzBI7d4S+9QwRqWCIGqpfz27mhF/4
t4LTzZHgfB7cfZzWPO2WenFcrkeEeW+t2KoPcnC2KSJnV55NnqN6h4gFjdzDOWTh
QGX9Iw6ND+m3T5OUvZRLq3pNOz0ovv+iJFWi/gZcVSq7K4Kb39LZzU0JHsnMZgiD
0ZQmSjGB+eZ3e8SU8Je0a2tS2SXKeo+XCVFlDzOc4hqCdSZwrLVgectjYj/XZ8D9
e0OawMkPUmuWay38vCLNeJacixfELoH9dHLx3hSuC3jwzNqVAO/rIEBo8rBO7flr
W7yHgh1HNjbYQOkHeMZTWg0LrpQsKqRtKBfPXPrE0f7Tt+I23PRpeIbfPc9yyzzG
tgMY/73dDN1zAAIAayxJ/vK/BM72TS0M3Uh7ZDUa+lbIXCxBNQ3hOcvzbbveBPoC
FEFTpTZMJHpaTB5jkOuJ2CpEWPYbNvLYlge0TFWtWoxq4eGIvdpYl1YjgyPvj6df
gI3RvaEngPne8hbCTM0I0Fej2hS1T0WJtFG6adqItJsQZvo6fk4PfHzEUhzQhkk8
dc6Grxrzutx83Zg/hx6p7R9FNz/SeaGEEDbqw08QayE8dGS92PDpr6LeQgT9QdWe
MvO9/haNX6wMBjaTMgO42uW/MQT4cOpKlOVvMV5jnoUDq14cuWn3pJUMdgoXwsMi
8ZITJXv4GOmkvEnv3LThLUbdb0w2ryt5wl9VrUdHEpbvpJfRFWnW4zVoXRxzjlNh
ZCn5Z4Y1QCFmYe6lQUJ6zmBMtFFdYEHK9T0eKa1INh6c8gwteVLb2E4Q84QbFyhz
euim6ekRStUmVknpGCmXXX302ndPDlsbFpbsNgDsYUz3y6XX/VjcjwMZ9iXr02df
UHAHRSrXOzjjjcAQL/nRm8pQqWoZHXspIWQ3gf1hqSxUyc46gHD1pR/+rYJuk9hf
ch2zcJaWr4grgwFPFFsh1FdNJQW6oKIH9EXti+ifqSkMcppyc4rqBhSnG5o5mHm1
wG49ORC9vkQZB6FhEwuLYjMWU9d2yEH0Aot4gonzp6ZN2fHvgrU80WKVn6UPRFZd
rxqmtg1prX/omkUukwjQglFcpSemDY6Xo++OMfF2syX8ASKOVcpElvdaVcNXdyhH
Y3CoH9GwULAnO+mg8Rxsj0KEl+Sj7LwP+HsbaOOqjmYzfbdSHchwsYdyayVVU6eW
soAamwonNQ7J/OqvQPvN3czaYENE7+xTG7Qzj8hl/jJ83BSbU6mMDeeWefadCB78
uFd7hcfKFJKVnR36rL1Yei9nt+u/jwDOc5zE7JG9fJqo2TcKm2NykB9v2mT58z+l
9KbcQ23r2A5aQdIraWPJbFBYmfs83Kwgdqtbd67n8GhjYtAFjc6+NHgcYCOpmAaO
`protect END_PROTECTED
