`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y2rlw9LqMrB2o+dSyfBHS4SOPfbG/dTQ2VnRSn+ilZK66UiAvbPn2e8Klop1b5pT
SCOxj0LTBhPztSUGW7t/jJRK3iP9FR0eK93N1hndtMB8vlY6ZnUT+XutoHEYG0GS
cHBNsInbROBlN3XrfOyfGMMapKpMZpBxjNOCrib9UWnqmz8RL4OYS/IbQjxI+Tr3
q7h2uXf+34sQCwzkdy+Rx5UXMnAJss3GHI3AHVewbezILmDnoLiTMMoMHaPUUkYz
n5jpD5lnPAWnu5QL341DyLWvPYhz9FXIa+Qelm9ztMRNe4Ue7F2ydHS54G5JpecO
ppbmhqKIgIXF1sS43CnK0+sIFpObC42EkxLYqsQtc2Os0Jqovm8z+8um2nbsjwuB
UtvIjU465tsCmm8wle0ptW818UdV6uFTyIE6xoCmG7au8AhtuHtAjrLHLkSC2HVl
nX0y3BxVBNB1p7quI7ygvH8xgzICAERL810cuBy/Bph0q0oCIjulnWgAEoV+9psv
aICZNw19NNsrcYg8TfXrsuAFUHazSCtn4ojlQEnlXVZRJIe2Fvrs6eiqxAhcY5X8
GXU2j7xl6b9rlhzXtdV8NwCJ2eaht8T8q4aDhmeIu6J0ORF6Id0tdmxcEDTifzMh
ifurcn/RiV6zUHdRQPy0tw==
`protect END_PROTECTED
