`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xIKzgF69pZKoFmoLno4s4MuoJF86woYykAZ444dMTVny0wlH4mIHWSn4kPbzGBRs
Neu4fL4yOPSZP7dALroy6Zqxe/YPrcxta9d/6cpt423xRSuqXduMoSQCdnL0QEym
QtReLfRFHQJVmyMC7lIVjKoFj67HmXeH1HwL0h+Sx64YlCTBrGHNuqBMmokt2E9m
WPSCyCwwP77SUtPdM5Q8qHiopGs2h+zEK+sxAB45P3GFyQ+m5LyFaD5JN5zhm7Nh
+Wbbfzh8FE6jN6DQs3UpH0KkrjSfRImQmzqZYWWKC1AAkoDvc5dcNvCl2/FC925t
+YZCUcIZrezd/p35a38eVOBeetesG/E7QRQMo9IiQRh2/WJ54GdaeAbJBZwUVKRg
tGdDK5eeeZ4hYDn4SCh+QZXlQpK+Ds/drrC7YDN98QByp9hASN7j3UFuGg1gpb9o
U7hfJUujZTk9gCm5Xf7vXM8kKw7M/khFHYb62siZv0iPRVW22GUCfr7kOXagUFXN
s00KJnsjQK260qExcjw14ASIXTQMLQn1krPvC2UhFlebsmGYDXDpRhJm0VV4On1h
xMifJ5XmZv6gR7Wk2LBbnFinAujkaCYPJu2SKJbhFIASv78tpCHGC/moW7c7qSb/
RJUX0SLlE94l1pY7Z6+veNRRLV7dN/Fe+4qT7vYICoihHDcEyHYL7npxl5rE69sU
oNS/OcxwBuXf8qzB1jd6vboGiI1bfWUQdFN0T2wYSBSiQGWCTVk3j+08qpz5wpCJ
`protect END_PROTECTED
