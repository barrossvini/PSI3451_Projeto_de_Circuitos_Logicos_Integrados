`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ZV0lyB1c/vcpCXUoriEFpBdlBkObPeCiqMBwB6OpOTPiBz+hh27xZFIp2EbEEyU
hyLaIWcps1gW1ZHtK/27ijTZEW52ohu1lsZ7BxYV7Z1GiRcIzpqHDAJE18qN0Euw
BDmnkmGmqQsOENsKl/1rtWXZ1JNuN4gHQdLuhd3JqmH4B6VrDY3UWHpbpaAhlLE8
qgthF+7FJ46joEwvqh6aiGBHkWDZ2DCnpVhC45DKLpr6tUb1Grl4S+xozYLgVOIp
QYOlTjs2Gd06vfXKGvepfTs4c6tGirWSDILQMsYcjI1v9qWLWE964hUQ/iCUMh1c
ni6DULoErHhw440sTBDMjnPAO/SRSatHZ6nrDqnYc41nfVHHCmq2B19E5Q3sA55X
+ERYcraxRK2Ky3CNrPz7IefIm6IqW5XsnR7Rd/CEbsjt2BEc/abqdqYAgyS7yW2S
89Y08y6j4+i3iUoZ46+QpM79ttNxbatzZsU5eIvl76kmt1C07ffhJIYreNpZcy+a
SZ4yJk9+jiXUb7C/cfYeMdBrIWrSIKTK3XnisiwzbFxmabMnwcY3FspWxSnIBvb6
AOtl50OR5sm/ndwWgm6Uhi1SeUOzl93B4bXmWGNxz2+iU/Vq+IM3zSRyut78FJRE
qFIw/MsnfbFbJ2eLj9FMPz0BpUqnqZU0twIyl8FS6p6V7pEescI/lzhdSZZPtYNq
PnZmET7HkSAlpiJxdnWWHxH50GhCqdLU4DwMzpiOJpwLbEEYr7ALYAANuIJNiPKA
yp496X8wxz6Z6yw0p2GLffvHpwjoOVgn1wWpRNsAn4VNAVbTeRd/KhN3BpXraHGw
OMaesH4PdfVH7WM10yK3ylESIUTlFjIShWOSoUIZxVdbZAu4+qhto7BtS6tNIW/x
wm4yJHAcj66hOsrtFOxSE29Vw8YBGC7Wzm1x/ipDTzjl8XGMoJyqwl6srRO2ca7Z
4T56DmOV3TvZXGKtg+tugwKoP+pv4vr2g6rAFTGdnw72XSRSZzmTfBNnbaXJDGuM
T7EoaPVqGgpiNHX7JjjkfEGgmDVu42ucyz8oQQ468nU=
`protect END_PROTECTED
