`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MeEQnsgRmqTiOSxQBb81IaO14m8ggNAWmmGU7DLYus+Ad8Q2cQXSrALOl6ZkE531
MJAP3f1jdvKD1UWnaY/vErErlkNU8SwdAGVFwoKTC0aAS3LmKMv92ShtOZraJkVB
6p8R02QVjx9wB9j5E8fowXnrCjt236/o5aW/s2rkn25SQhazJeC1UqDAaiDXDYss
egVs6Itqtrt4/QJl1zfxa7lfG0V7bVQPfUFTiRgg9ymwb3AKvJrH8Efkr+PVTuFG
NLGt7MIpqJ6f7FrQIQS8BOnBaIRwu7Ni7ME2gau+vyZjhqF5w4qOvdd4/iU71y9C
1fZ2d5Z7kaY0q6Nm211ZdM0VQFnDFnGor+qQwUfzThwMSFEnhtL3DPjtSGVvrOmd
gWKueHzHFevpE26M0sfQlNaET2+UhwbHwsQMRWs55apQbD7Mm4ooocUfEi8aJUk6
QMGncadwzdltlcy7pGhn06irosaXdLomC4zWTps23rpaFu64GO1Wy9+bReJ3jf3N
rz0g99CRJJCWIUA4WbkjWGaZ9eMrFdI2GjDFnEAXxxZvr5DEZc+5PmL3CigP1WQM
pEyKu+Zedh5MjVuaadtXvfF4cvzCslEcrcP8CML2p/MA8fvQA7Wdp24gPN8MW+Ll
LJsWjKPTgtR7TazgXs1B90g+5m9V2wnmISYpBro+zXiCDq/OfcfyWWhLw4OMjnnG
qOaDZHgvcsUN02LPxnXu+Uslg0ec6Fez8MKhtxc1aTmyybfGccya8Fmy6x2t8csZ
ImHpBTyKZoT8EM6jX6Cn8ZDNKqWW/Fq50Eor40upX52S+1nID/GylMu4DSyq3qWe
PUf3cUlLwJsQt70lNgHGfKq+U2nIQKCvixczJfDzzrA=
`protect END_PROTECTED
