`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5QFIOMXHutJkw1WZlf20ZLMTEPChy095foFkGUGEjtaJxWLrY4akCUDPPw+HPozb
917trfAzHVee1H6Ni327f8gvFEWjDRiwhydwQ0jduVjFMMN/QzMnSRzxwFwEJgpE
jllwtzPUfvGb4DMoyZMbL6e4AbuSFGvQmVJXHd8xReAe1dJobiITMHSZMmqgl01u
Dr7vb8aMutKjJw4q6sFF+fv6piu8sDEcjxkHo9Jh+hvUVsWgUoes6KDrwnvot6OL
cOklAiFIQc3B0nzz/FvoBw6McIwW3uwNDq6p5ZLaVIhi+tu82zcZVQxiscC76+//
6PeJGx246Y+kG4i0t1Mqm980Mfr66fEulE4wS7arYfexca7uLOSsknSEJkuhmYfc
EglrZC9BbhICPSjwr2570L2joLkkf0w97YSzCYdY4BoBxYwLc9XtVsJ1Cbd00m7/
8te44WvSxFx8LZpPxGQ6an6R65a9qucwCwL2CgX5ddlQP8/ffN2kTguhP8lftbsk
dLXIE/SwnhpANtIA+MrXSABgivxcQfhOVZQwy+JDeBq1lvtWOOlwGO4ay+w+mCw5
kvVWcEMR0nivS8SJchrKURIq8icYgSNlHAoOZquPmDSaet/BwuJYvJMY5l/UpCzQ
S7pk1ZUlZsvJ0duRNt1yTkW2olIDDnhUlcJ5Ba1icfB4b+U2pPWIu9Q+X5cHmhHf
cx2xxE9aHTgZ//Dq7puagllffO71ixbcVJiIVkv75O3/im/gX2cBYSKGEqo+rKCB
YECllWB/tz8x9TjPSHjCm2a29oGYxhoIBS5h6CX2yAH29v44UU9yV0lm0SAXoDfN
MA9+HTwOvNF7zMkxd05BDGOja7kzpBX40ooem8tUF0Ov9wu5H1OM4msMxajeenkr
G05m4XPYttT7Iyc3R63rHrUVl32DF6A3cujOeA9Ifeid0GQliUPjOk7jQHfm4SII
tUHT2SsvewZH5wy0A/J0/zlOcc1jgQ+gTAWUXDrDZ5t44HR19gOVM2vDyZWZea+O
78vxd1r+n+kI2j63t2D9oTklIILPTL6qj4bGqgLz/ZPjuCQdkKIsA5OY7NlLJ4y6
XF8oSGGQTRjAEqzTgyilcHDg6ZJ4lksBy/pYgLH9IkSZ/n/hJcV0ncqoHpEq4KT0
aAH/uqCHTMBmLt6eysI6HpBODj1wRNep/q/3I4SaMyZIAqgxNNHbaJqHDQjKa2U2
LG+SIILub+ogVOxTQcHVdYxs9j3mu13vBDTySKHW03OMa0Uesxu8LabCK9+eKaPk
3DkSOvgS2HJ8HKzGSlbpEvLIQHLFUEVY5rciIica5p6dvR5ops6CaFthepSQVwO5
bNNI6veVxp5IvsJsabnUFKHVULfgXLwJdBCXKel4M0FlLC2/KJaVnijQ1vJQdI6x
cqrggISz34o7SknFhkLfgGQPwC7OO8v8oi1wL5AQqz5Zn8gN0zG9OVDVtRB17k1J
ExelXqoGpzWjOkjzLibh8daERsJKMPtlqYNrncHMd4MkyjsD6okJH2h0mR4BrIc5
pBlF8jv+rk/rJIkNpGzyvYGI3fUo9hVs11ON1R/Zi3orG0LQ0ArXbq6hWjy4ZjIe
gr76PGFJbuMhNRSXrV/iE5o4FyKMKtzJHcVKKq384gKunrm108dHlEurV/4esOtR
fyGvAikZIwHYF+dPGEySfHr+UUwfeVXNun8rCw080XNc4riAxgR2J3XrnyOqVPJv
jkpSPyihgCO2R/AZLTpjlS0MW83TpzBTnv9TZRa9eIB2fToypWmBe4YI6FHqSkeF
9ebIFLAn2vRkjcasfa4MWw0gG1gRnma6lmeJ30u2LKc/lU9Wg6oJ883cM7fsmtGC
foA7O6uHNUZeZEzNN211NGw4goDc7UmSaK1PcD9LzPiwe+zIualEGEnIwz3iOVP1
9SHJkpGKfqxWqoucjywoYFFAXlSm54DOSvfnStuTU1hSkLu5uYjFXhHsDSlEJ+hs
a03Rad7hnANDpwKuI7kXhtnm7Le/oJHLOAWz71z/ZDVvcw0oe/wFNdPxIml+WWhO
j/Xq7hJlonmnew4PMvkltlSN179Yc1nhtpEVUASefNI+h6aehQWXsVFzkZl5ur9C
pSfxRBbtIzAimTfUNkQF++ctNOSoVZRCuR4qpeVgVnDxuAdsAuX0lDx8zizjs1m4
IjrTtz/4hhPgOvfOkaPNkHLHxxeZoayD5YdG5zi2zYyL1bRVUwskAIOe5Qwfhtsx
DHAPIx7UdMp2Mv9qMbyHTWFk8qTXdlO2dcaMH0DxSZ+TJspH2CmFZ2YUqUgImUuY
TxquVp7U9lpXs0xKPKH/cGCpQX+EOYEnh3qDgs0USE5yGCUCmR1/SHVd/qCRJQF4
BmWx6NRhFfSf7vMWuAxZX7kIYSJM5AE7h8bpC2UPhhcBl6YyGykUqiye2Utr+WHt
G0Y90tyxvaoJq++X8Yyja4AY/Th9VHGFKB7Dk0oeIf6+BqJwlUp7eoDZMkLhkUcO
giYIlEVRXs0iUScA6mlNvgAbzB90KE5WNDzaJKOCCrZycGqihDYuBxgkgSFrNOyQ
6dl4dyb98QOtwtZBsi4mU1PqVH8D9rjdkD89KdjjveAOce/hRmq2uYl2m2BUUlyp
oEffuXIzela24nTt1C2UaFq//RwwBMEaECSh3NwNffctUedgKk7BwgQFGCEIihnB
0oWecRRrcSHiGH8P0D2+Wc0O62Yl+vAUTR8mmewbsygcJCZjrsGARHcuiNPqLnJa
AZi44NwpQ8SVEoElTofHeozuz/WoP7Pu/a5Wk/ki0M2/0ZopZM28UIklslp//3ld
EroG3imAM+B/kDz4AknzesWKKFJVBgZ1B6op+AGfKaIJkrymEnDAQuQIoDqFkLie
Stu/91GYAyiXHK5lPG4LkLx+bjexdVMe8w/SfFyRQ5HHg6GzG3Yt4bVEgjmVdrGR
VUBxgtxFgqUFtnvxOMDTHCpLPlRyLU9fT8reNGkorMLPRJMI5YSnFAYAYOQqqgmg
IApYFoEY/stRxHmdj8B8j8w8orRFAbXdGJcx1irqucjkfDzNwG4u0WVAtn/eRbn8
E8jgrXvr1JprTKlyYnySDF4P+qU2kZZnjT/SHmWNklIybKNadQxHwTSLcM6reAa1
fEDxL2fgKDcnCJW/JhVUKATkKgxEbwxl9EIxDXR2iV/A5XSiQ7wznchmyYbYga1l
1fKVTTzjP7dZ2gguNVoteq6WxyKt10VU/3MPDJklsPmgqSYXd/vAiXzUlj75H0l7
bKxAa4izBwgGApt9KO+oXEP7h+j8eGouQhIcKJkCM/ds9oP7Thmu8RP3fmzscH2a
L/ViV9g9nwoPJYZbp1QPbi58amGGt7Z4mP7PDwKi+7iU9FC0xwncTopBgmwVkz5P
55rzqF5o7CTw2/cFcvZNYdlVhaLxVwLbnBCaR9+xztM+E4zCaIZ8+veXpw4XsQUb
3Q5HReX51IAF++lCzgGpYri4spYPlcGwU02XKUdyqwZ2AQpZu37ydz7uPq+lmISC
YFNu9UK3WND623bFwj6q62f8pj2Xj7iQgUPKYp/mHRgcH8oqnWYiH7Hf4onIIJLc
JIWxawCG0rdYwYorL5/TkjhYy/DWTqN5PiCZyFsf+c4j4Ec8UU9K+3BsGMdwJRIf
hDdED60chkxAXDjuOM43MLvWfKsE0nYPstL0mgDpMQzoeAT4nFq2bey2/Ob/Ly2N
N0OpPlRV5uNZBjV5PaRsNlYOU57n2xM5SvvrVqVuWc28v+9vpK3S89QEckvJLR2x
AjhEbOMDINMAUDlE7/z5LPx+j0u+C2rXM8hko3AvNRakasEKccTcqk5nqELMJ61N
mHwH/cMDKCbXWJ7EUpMCSlx04ohcuFtp0ME4lvbQa9wAFepGraCmgch4OEiHlM9Q
/i7QoxgxJPjU57cbZMgwBvfX4jJN0n80lNVx94VPDuryk4jqjlL9dPs8eegRqpgo
J24WZVIk8AhNd8mLyuBOXdbh0JjkQuM3c8mgcn8rVyR4TKeSvN9jST+DRp7aS1lB
aP+4ryBwr99+bclF0QbJr4WazLChEh0BUr7bM0gHf4M2Oql0fF03SncY1nbHSics
eNje2Hjl1D2/rBMBhExeITgVQgGmGVj5aRMiAp/ZZFG35nfgxJ9f26M9fEtyvi7V
q8IhwcSODTiSXBBKH46CBHlwVBhbyS38Xszt4jqmUlFFRipEc8AFfxUPa7QBtSJ5
yXclSYZErfyzFp2gSLz+8dUUbzZL9BwzrZP7Z04U0G5i+A6hcXwHCB160T33TwXe
DwCjvcBmjliokaZudgRDSsdB5G1mFcgcjJFANXTlm0rlM/o17AE9UYaopmZEnE6S
0IQSfDDW5hCJZ2zFwsOVA9VPn0sEgbxB1AIxyHu8/y63kHRqGCyqzdexY7SRUhvw
ajKSSYmQ3eGSrhXuU+N14rTHcLY5Kr1rCHUdWskWHXjqr/+87YWmN2VT8DHteVxj
6216yVnyl6pbtSRr3Avzoml72aGewULiHFno3T2bEtHFsU6570tNjJpYyb66H6LR
tMrCxwvv5/siPsQQltvfyUNfhMvrmRsppzN2uoYs9kDKbQuOTk74FuQqL25TpLp1
8R0qDprvZQFv6FICRxC9+hg+uXjpJPWhIf7R7N9JnnOgXcLOO2ki9tlV6B3UlmPS
CVsV4PW4W46JklSvCiORCIv0JaWgqOj36t9Xh68m5kF4YyvEWAq3xG6WVE97vI2i
ny1Mf1xLewUq8ltQEmo3+nBkS9LQxCHxJKy6d3Jh92xAdQyWebebvrjOX3cMoi8O
VFEoNvPsxMoyARm4zxsCOa6ZNXA23gdA4D3iJs9sShsH/UkNlTeNXAKsnLlwSAuA
c8KmdnezHMS7bR/MZWSfUUI7rhXvG0a8qHYZCSqcrwKp5tcg/xpQS5RpvKX4PVwz
wvRTKStVUhXyro0SzlS0REOfo6E/BLDkFHrNJR/jf8K4VMoy3Cg3UnlUHZ+QsSi3
vqxsoMCvwCvBQ1FTcSDOzEUKWHM8UStEGEEjHnFBpuNk6VA3IIuLpDRbFUlLiw1/
FnZRGmumINxI5f38PF8Gw4xi4apYhoVmSkFDgOhl9qM+6zfVlCkZHSE/I6Fo1n4z
81gYZrYTKQ94RhhJDxRYYDk8Bj645F9UduQFHGtpVoJON9yxY7fH5XLPOOwuxs8w
kgAU5gcozQyPLg2xW8aQ7VX+6s5fnfQCj7oepO4+gqixRQHPKKToCQxwAW4qZthL
6bLzNNJVMOSfg0B/+3SCd/5awJFXLTLJdZqnCqz4PdWURQ1z1/BZUGMTq0CrkU46
luK5D3UNLimeyp0qgkT6RnXVAMLGb6BLa5jo6ZTpH3BrQ6KTajZnWRjkx2Ysa3AU
TUo7ZSblG0GHPiaEWI2l8C4DddAWmuml4T03Dh/okVgJtGQQzTvxOrpqISk4kUve
I7FoY70gVtyrF2K3nR1yCYm3q+aybaLOZ7jF2gr+ZrYjnhTEBZQbN+1z+ysDqfsJ
orL8LBYKsmdGXeglHvZ7ezkgSZ+eZbs+7HkS961bdRHz7fmRgapbybTO1k9IY/aI
vGSrxeyxqmpH6w5qNnMjmfI0hLH6PKgVOKYK9hXwLNwWzF/BCsaBenwhK0WbTm5R
jeOXzsKnqzLhkKJVwjrUiLQbRStUQz+yjtX42iCy95QWzD6aikZ1/kSpShwInIX9
vHT854WKMd1kX8G66/VMD1ylia3TFEwedv5XaYTeNwmdi/gT/sEwlahlA6XphmMk
u2Z4ucHxeqEUX+gUNCIzWdICHH6ImM6O2bcaZpl3Md0NmoMnsMz9Ro7oXdlVExjd
ABvTdxjhXgQ9b4vSYHMLPANzQH5a27b+bNG3iFnUxOWoqxoImc8ZSidFzgDBEwne
ikFBBlsgrAWBMm9cyHdAf5qUTP1kbeNGDFPP3S2oqJ6R/+dnuQagq/+WFVpdzmfD
pJGHXX8hALJz1lNVQiop13Yx06EwcNGb9zaqzSJf4DyNspRV2eoOFVnxWDDm578v
kc8zxB3yzl9JY6PwINCVGUhOrtvS43A272pbJoQ2yq5PzozMjFEQzM8XZDHIk2e+
00q20at/fcT6trMudyOw3pLKFDoI8KaZbpzpHHgwlMEWjlODw+4+Uz5nbXXzQNJn
Tgub4QyhVXhkTo/dhnatDiXpuR39JBvqw2z0rGEA9r50s3LWbu7kl0UJUhkxKSJh
VodgYHrHxxAnr3uknJL0ihbQt9+OZRfO/TiQ/3HBmfa2SJ7HP6BH9KZx1Q5YEOPX
A/WIGftkQwKFfHt7+wBv5x4XYShN1oKp9CpbwzZe2qPWGNtEiyg7Zlm9ghIC1X5i
tA9hqcUq/GCsdSyw3JTWUD7e9+wFV7B3NysemW0w8zbykQXSWtzbz1x938zqq7kI
VLDr2HB2PVqv1v2izJaL1ozoaVvx/ZJK/PuZ2rIkf2z2xjzM31m6H2L9ta7ry3CE
QqKfqsOYfZ95I5kzAdpJhhD2Q5jvUpX6RtF4QInStGk6M4WV9A1Rqo25nWSfsqDA
vtrhgSPxWsk/qy9Wy6LUjvHlaBEHHN8tRUrk0mWYYIRpnQtnmrMwfCq9AoI4ivnj
e90JefcUx1PlTPkBwwppv+n5oCA7pjUKOmh2toG8mF7hOyFYardQbIWQP0lGozbI
7jxeGyDdEoLxGX3/HxhuPofcQ/+08tsxzTtUAazxvecShgQEDkuLTDpmXXzITlgO
PrpzkJ4f0wqY22cott/qnH04Sw/G4JGWYJFzhxwL0NoLolYwi5CHP+KsDjgG970d
RZsBA8anvgDDRR+HOl7ovHGcoaOAeo0M4FcX1LA9uZDiFWgAanAnvDoyfljZp4xe
`protect END_PROTECTED
