`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vwUet9W+B1m6nBxb4QrkGkoCEyRgZke6Eo4TPmFjfRBZk++S5utgVjTRnV+nJSql
AgQZda+W/1vtTkcqdfu+Mq+0cW2i4MHo7rM5oEl6z9WFNx3M6s3vjkZo+72mc+/7
QS7/Kkzprd9NnOlWug/RwAEYL2YsS6AcEbSu57hITuN3QZczKPnAi4ELfYubk5Jc
POLKh6Hr3OvgHZaXmEFBznh5gqVTIufhI+ufl9gBFs7vyDredOuugUm+5iFFmgSq
I05cPoKvEqa7dYZaVQNlQzMhqNFHlAx7zi7TtdfO3yC2HaOfpoEZ2XRRjiMkO2pm
mO12iVvNkcHTgqD9bY0jQKa80ba3BIf2ez8oEd6nS6u/9p/BNzxHeQ6J8KCTMtyr
AY2JWF+71lyi/krkj6cB6eM4oTt13x4vqbIpqULJeZSxX0pr8i1ae+3iaz+mH0pf
bTh1q/LPRYRBcNzFkh0I3jcM/yFs3qSGnxG+jz7W4SyP/35ooyLdNBgnjlbV2xqL
RMZSCR5+9JXtThYOcqIriH5+yb55or5TaKZwFFtMmYmfnspvQC+y8ZlRVwSTzNcL
iuKsgm0bCv9ZLyqD9qxzX5lZw8dqxvf87rZAj9b/nEf3RtJeLKGxhV01u1UOkmU2
LHOV6wYt1AEhY5xXl7lBvb67DmWkrOAwiRDfHOeVCRAtivRDo540Nt16R12JonOD
6bMAn3k105imwp3M7614YbZZc2NFwHMmaBw3nFmU3NXXcAe5UU0lP6W9x6ANejEu
SJRRKe41xSqX6kmKtvZdzIjUbUcRH248NV5Ixt7kIk7x6tBxTtWCnZYq9TwUW1x8
QAgluhDxtx5KV1dcTa1k9F9F2ezre5o5LJVAM99QOn9gusHr87HHCqwIH4S06pje
nPzVMOJ+AjXkGGLyBJbtv6/tzVw98Ffvfh4u3TxkyGCfYTU5zxwSUV48q69Uj8Gy
+iykvY3iPYtZIr55aJhi55c1jO06+Z44eKZXdm/8WUx0kc11nE17AaGb3gsZcbcM
OBD2YHKY6lZcsPH69Lok99Ac1xmTwAn0DJK5pJKDl00HwMh+wxbBIjnol7oUUbum
TkhKn+ituOGsz5s5xOv9B+ZkKSmjwvTZ5A5Xyovtt1uZoCCXRtnNHbOntbxjEZic
26+z9AZe8G4T49qOFxyzuOil5DejonZxCusApTlgfw2puEaLeW25D6A3jnv9FQl2
hqU32FTjXDMXfBQmlADGVQp/Y7A6wAH4m9WTCnOtDLxKTlrDawSwhC6EDc4XZLQp
vGJGGf7RF2MoGryMUrjEAr37PsL0LaGxGBXIMCDgDyAEbC8hESMM130Yvk7X6RFx
xr1hwV+afjKuJQ/rOu1JmFMX1bX3UJD2Rp6i/+ZbrvOm2r+CxkNUcr2mEBEVhbP8
XbingLKn5MjpjfKaRbxnzXlB/WyrtkvNchxz91eKPVM/CzxthPxUkuivfyFR7inz
VY5OE8BuT1njvie2NcFKSCSfjv2oR28BXhEmCcqXKVqMwavUNhF9uFAWqGm4cJek
eZ7fTxDKU6yPhCiaGmrQTWVkXNE4ya8mJpR7kVytuKU=
`protect END_PROTECTED
