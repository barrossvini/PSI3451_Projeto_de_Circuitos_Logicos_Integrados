`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bG/Wm6uwLtQmDakO787zcP01gg96S6vVC00C4kgN+Pq5lRhuC6yYWnuEV6FOKbOW
dLlCL/APHqxuppoDon/yjfGYZ3QM2QVKLbFM5+mexddPjJJdqOgGd5e7dmvgTs7C
f8294O5BXyE3ehjzd3/b7HBHWysR0NJ5dkra9fQSW1YYnAw5pGGegagQBgEYCpgp
KxWsmcXmBjL9JwoPbC8dWQP/6BPh6Aa8efqNizGFTh+D4IIFfxAtVTRaN8BcOc2+
rbwS0DaPeLD3YZXj39E/y5HgvhwRUhvRouNRpZgE29VdF+8++MWjKpHwKLeo51lB
VRA0IO5k8csCN+YOOKsYoC7Ncs9VKOZvu+oby81wugYiTmE7uSIsK9dt90kHwqjB
dHpHpSrFBBAYfPRKJpTAlundp/MPgthHEAPQsm/nyTSCgDHBWfwM1xRDoc/3H1aE
ZhnuL7IPReirz6tTDefl/zxc5nJYKrlTJ5bPDh0KCNzWsvrQe0x8/P5KTBPyUsfq
x75DoBiznX6pcnQU3ZwXCAxZGBu2tQvWyozXWMr36z1anLCOWx97Vys13wzMrVUF
JP3iP9uqzWv1l1s1/hwAA+Q2SRhZGLhat7rbT+u/FD9MjlztDo6j9gzo9PofZlzG
thRtQgkP9TmDxkS4cwNBhMHXGMIAVv9svDEcvjvDSxcTmryRJBksaQV4kwmzsUWl
ISB/hv0/1eFgwrCf9TaF7NBYOMe0jd0HMz3f+nTlI3JaA6VDK6zrx85RYC+jwfn6
SyBGQsit7/Hts7+V8N79HWMOdkp/WtJpSs6DUqthFSQ/6/b7Y0vUe2Y+f/iuF8VZ
CPWUC0TOArBcohbOsz9nu6odNJxp93NWue+VJ6uFpqaZv4GGlvytQf4079z6WKPy
cl4afwRNGIDWyAfkLrI7SCNuSh8bAs3IUtv4J0LrQdAHG0Hg9KPbAR1jQX4YJ6tq
Io2rVwqGWcLgtw5Xomya+8tVM/gPn5+gmulaKLiS2jKDQVNjGZAUPB6saO1qpQfm
vH4CjStNNDUL+XyUukqRk7ohD6FWHzio7wwcKnJbQ61RMDlA0xLRoDK1C3FC7Ala
woT+9xXl5gDQEhTn9SmlI2JdJwS9zXvlfpmegczBuj0n4oI8pWQl/P7m8fdv6CyF
uKX8K2cyJshmxkohmX7DGqW1ipvAt6AgQPpzSOh3VZZnJj+/uAkwnftwpoYhAZpk
c4S8kZ9Acsx/yb7d0M3KpRL8QA3b+wIM/5fE/l31OSgO6YZzUeIZRQPu2Qs+0C3H
ny/JBzTPMzfOIQ7vb6kHWG4/3Pt+0CrmsyQ6M+kkkaez7Ky+NHAd8tJkNkQPE2Ql
YwXM8/TiHCMmTrDhNXC15J5yYVoAryi0QEo0xcRYSiyir3g0xdWB3jKY+oygCjdM
jge+Y5gZBN1h2EtD7UwbIP56Z3JvAhPsMWAx87CG4VqqBlHF7L6+/3zWJRZBDu6A
9+xA9QEFzSYS84xbOyRbKxw6DLsQ0Zq7gmuwhWs7Itqsie4aD7vo4ZqxHPnz1D2A
mmuCh1/FjRyTKWO4fi9Za6/YuoIRGNBlKr90Ng4vTf7rpGd500xyOM5FR878Lbw8
DTujVblrjewY0gKZPpNan7Gyyrm5YGHtNiPpXO4JIG6j43O6fwW+DX9gtgbk76po
CS8eLscQacP3gh7acMApMua25gmvapTtF8uFX5TxCiWNNEc3ShS8NCGCsA+gVKla
fvLgWAhQzj0UeGNg6IaMI4R6DfLkInZy+g1iuORmWXoA2h8cQkogIx7Jr0503qnj
CrdkTraM4lqUw6VMtNY4+nuuIbfREIRrBKYbt03/8i+yDIPrsR4426HWEVdPOORF
csWEDfWgMh1vmEuj/tLwwnrJBWGM1qE0d9iu2FyKK9IgYmt6yMdY7L5XthWD6eXV
jgXvlG6cWoBK5swFDUjQGDdISpSw7+lw57MUmh+hINYyfJnxcvcC8/zBsMgSTrM+
yH7K2T0RYWM9uWkHuc2qBAtWLdMOONqU+njCMTOalxYxeGVJqvSn5TpDmRxeRjJC
jtmXgRjq6H6CIO2HpETgGLZzgVIQttF0fnCeCwzScUljEZy8+Y3sPQCYx00s1Caf
Rgx8+Bkbse2yVbudgY6xElUK/3IC/rkEIV+MeaEueOM4sJbccjVUXZHUAT3tNrBM
ShKtc4NFeBKQdVBqWyCmR5x3D9S7n28fPLOy3VBECWMoBlJHsAozRarGmE5Ah80w
jRyzPnfxEw0VaOYyD7Pm3NV8mu9Eu0DVNHIbfsR2qLy9ZjKKGXkNsvdeSopcPY5I
B8lVXKyG4uA3Z3Y+7FeeXqjGSqZfZjfpt2zuNz6gcBjC5Dartw3EWNdiFU4nKeQj
lcwKMNrWdGFAvT1Y0ikAzNk43/nF6BFkuLtAl1suPlQbxV4UizfzSKp7ZH3m2z1D
FKHMl/2KFVgpIa6bH0seTXTZHCq/9Njr6a6oOtdRlgG+pf9ASi25hvr/4drlOhA7
t6U1NtzKL2yXnOednUEeDaov9znew6Jle+JhvoSbGnBVOxwPZjpkvPUaaOipTNt+
nhnBGMLQMsFr0yZ3jwR/9KLFw77WpMWDxjhrEvCKwWwT8irTjDO4jsq6HZasU3a/
2+87jPwCHIupxK1X5MZL1nB+RKJ81uEmzHGhqUFXcnzUt3feZ4wnC6Efgs7PObo8
h3EjWZt3qJjljd2LxDtrDRE4nwDpgGaBN3FPZlb0wOZTvJeZ7f/4GXSEUfLVd5cl
kCtUt08hjKvwA1bQFsL8ksuUuFy2bsfiRnGmbdpFyjUOhVGVXEQHgfi0bDZz/bCx
oHl7XVJ2UBStSJk0Cd+zn3z4YnlZTGVObaTNc3aqL3a2XB3t0d/B4zw3R/KCK2tO
77WzDzH4UMNPpQumtS1Ry23Q4PSoaljgYFMYrON63JBvHhdWAuQLT3GYa3OdYBNm
QW2vpyp7vatEDQ5KkbjUG7CNhcqdjLO7jpH82IKswKLQhDdNWqDJxJbuhHoBoWzP
+fV2GBJiXMR4BiuveYAxv16Z9W0rIbo7TgWIsDNukoRLHYzJW1Lo/ER5SxZyaIVI
+P7J4tMpqQFFxTNP3gF2y+f6Dt7PWuikdYjHb6S6s13eThle3PYexQFesFp4SIty
KuBlCT3B0CadQ8HaTIUnFYNK+P+pSbYlGB70Ad9ioNk+1JofYazGnyJ8/5t2T/dq
XNXtOrF6+CwfZiwohjRV4ziz4ak7Sii7YsLL2mXPVwmFtfzSFr4XimvSD3Hq7Jnp
xMyHCKJP+gwndEgbMF2ky1Y2hr8Rt7fM4TVee+wxncjInUO31HpKmuSVqGcty/e+
AyOQdJQuf/5HALGtdNzAqPlbtcaIejcb27mp30fzW+V50/lSo6qSths1K+PNxQ2c
e6ueujvZSHwk3JJibwU7LDBNhd9wcED9OW560tKYaF/jljXADBdTgxIMYwpMzR5b
4DqS6qx/o1+ePASoBpJJTin05pShs8vXDg7QvQ6GWkJw240DhyVmW/4Mj7ZUV0Lm
NjkqicvNnJRj8OKT3W9oj5BXPoiKOMdcVSgHGse3ka6YHdR/KYnx7dLa6v9T0Pal
QH85wKy4taVseJ8PbIMhHB5bnoe8dC2/PHfJMMQZ11GlETwHBiD0xmwTqC804xk6
87NmdemeYr2AaCeNP2MDDj2QChDALesx6OQCauKeAnYfaFtSvWNv+IE18pwvE3yC
u5bvSpjAcIA4m/eAhL424I4fU6bcnl45VrkVik66kKCCBHr/+SnDKGtLTohTlvvA
ElMJ91F3jneXAZSMNgjl+0nl4+7TQWgyIGId1w9Bdlry05xDljvnIJlDGP80LWLN
t19OStU5VKEBSkoNyTt8kRaoR7LyQpud0ea082lbsiW6ERlh/dEBE1/MpIIWHXqU
Ijt/9RZlmHqZ5uQ5+3hPFljHtOuwVgM2QChwGvmsD6m/RfRbn5MwlpS7X0Zym1jG
ZzdKOz8VSr7PSxFq9YYDKrayeo+PUbt6dhmLmqSCGe40m7ApYYXAgK/1Zz64Kyvv
naeqNb1p9OlGtwtVPghrZSV3+l7H+PEToaqNPCLp+bWotoOAXcMdLWnOJch3eqlu
yR1VQlRU/06ElXhi5b2/VHPhAD32ud9To3qCm4mp0YLJm0wHywqPnbfAzmJWl98l
Yx7xNszTv8PaVVaM2BEdzhZTCKWlIsRvEgkgp9ldrjoSvu+4qWU8ZQJChi1yphWo
Y8Q6k8aFNZ/6//LMOLCj5NygH0UMMfB8lLWK0WInx33zls+dots8PxVSwajVJb0d
/A603y+ZMzRez/jtVi3j2TcHbLvfjhGscntjZ/829l/RlF6wQhHkGbU/Da+ac75F
pxqKH3uVzIDlTCiUMzctIRmkczVyIRTCjZWc4jIWmCrQSpA1GwsZH8UCG3B2kbI5
sZiDAdnQ6WMj+esxaUnrXmV+jeoPJevQ3LcgEeEmes7kK2EoIjW20DONIKucvlJr
RTkE2qFMb+t95+ZlvyYLGOsj6kK6SDib1oiO6JwzLq0v/C6dOj8kzMwn/dizKt0G
BZ7tPcYhdEVPPtsLu38Gg+lcjnGuta/+cGXfggcjJAJu8ZvZuKAtrVz14dnt73YN
LRq+AH4ZDCqZoMwqhn3NHPL66PGNdJy2JJLtVPD100KUEcpN43jwj+tAxeL/1Y3a
zRo5yMavWAKkof40BJiBy76PajVrplunxnaC5UgfdBfYFqd4BJbxm2m/5sUC4+Vz
4CoH7rv+GLzShGdN/Vd6pfDeQjbmQMhNQmvnBWySM3jYR909w1eKQYP+bcEBCWCZ
5NXJ8KMo/9ySoPcYMRjhNpE0N6AzhyB9RRkKt2LK9yjloNcbG/m9nVuespEcJKOS
Kcwun5XYLpCzZrlDwGgX6txjDy/PhuATHmq0FQXZeW1nLqmebp0CKOe5x14mHmCH
RT8qpj1I96ytw+oDjQce965od1YRSukp4XV32x7DilWYH0V0oAwmk2zok01YSBvk
H3Gyi4SpUKHZE3LailRAtIQysjFnJiltFMlPQjarX9DTbswNt94VIBQeYqVStUjU
7GAoM2fn1AgjqgezwBkyEruQCUppGkvgdEB2sKMg0bjVnHD+Zal5+01s+9INUABT
LWqTmXWQ7b0JDdoGkDQh/mt5RLdKMHrB+JnkMcDsV9WhaJ6JI37BohTDGrDgdtTR
tW1ZkU8OaF0pruX3a13u5hBwhy3QUoYDxxp4idUZ5KXjaqvSi4SlEyDgjCof+MQ5
K6sn9E++0RVs/ovs/Nka+b1i8wwdOOGK8cbcytxE4H1Mq0UlL35JagHXl1usgczs
AWGF8Y+Gz4uxE6x0BITdlcqlzgHqz4PgzQdBjeLxpS5+VjL+H+A8MkSlW7uQXkrc
39/lrNjVpx/8Rzo+sAgiWxHYrP19+6N3yu6JdIZF8M8c1vmUwOFA+Y9sjeG/LXJf
vzk6Y9Xwsmd7TlMbYu3aCZVXlvjGA1YfWJEPBQlyZt+dvAAW/zBCEFBrKRw2HXix
9Tytn+FJ4RYbl9LCcC6rTwIoLfKZgct5IGh2LQN2B7S8TT0e8XOPaadtUpxDue74
Y8V4FS+P7YcmzzZT5WVQ0WIAwvyTEb2zMHD7mIaerD6bUfxxiLwbpN04NHTFRrwa
xT5d6UK0iQoAyS4scmNlwqSRNdq/3mQXIM4youbbIv0e44vdFo73rWi8G2dYZTYZ
JF6u0P0/40fVe6Da3dmrf33Yk3WsoiXeoYdH4cmscC5+ECJgv0GosMnvq35AoQ3l
nzrYFQKhbq1epVHnDEG7VrjQYlNPJ76zzqjvjwjttB+bQqn1sbMADwLh7aE5llY9
tvkBHgfv1MM3LXTfn96Af12RvNUoXfWG28ud1D1kQYLIOfP9johCkNQd+8siR+Bx
L3JsrVQ4pRtHfSiog5E+AlYNdf4FY7sZFfJwBNrIVcPu05eyMEdHDh53quGcisZB
PY7Hi1z3NpCmDHb145c9HpCKZKSd15BSdRWxMQ9IVR/yhktP/9Md7CbwhMm5LrTh
vYHZNUD0Ej9ZI2zvoDWSktLH/6oTRipkrYmhsnTLroGuP8avkuIj//I3gc1b+H/C
m/dR7ipRrFZCUjpEbak7e6Jo1yjqWaLp5JBka8wV0ERbE+xRavQ3k7auGcjacw+c
FYI1kGLz+ESrht2jBssub00ZeUIfSFgfQ+KEGN/zNVfOo4IHdA+ExONyOwoU0qiq
/PZs2kHw1FQfbmiTEMEC7/bhbPy5IstF/k5M8eGw57CobHtOoa+ypAe6T6GUMDVH
5gauemvn/FmF/VHbWuPMvLSXgOM/Y3LT0Q4dWURdtKlaL1YH0VIiyflPYsuf8YMV
Mc7CvnsXQGz1Jueij0Pw9QBdTLmQvrrwxjSieIuAt+vftWZmVyiRXnDlMcR+5wvH
afUZS1a2fb7LMNVc2vu5lCf45sOn1VBr4A89v1XsMTW7gOKu+r601RHFFZcTXdPN
NWgWZdwXRaRsa3KL0dULncYqLC8/Pwnip0oHFpBG7v7qZtsxvZ59Albn+MBcLddv
LowF+AQZkkMGb2H0QEAnxdvYd91+vyOGSrmLa2CKnB9wb44sW5fPunzSZ2alGcAL
Ss1skQMcQbYnMnoZx7bDkwSU0Zfk1OkwTYzS8JYfkvnfBe38R6UYrWvgM3Nde5Cz
U/odYvDAKnqbGGfA5LlveCjpANkbLJvd9mRPv5X2jIeMGnsTGLKmygOWzNlkCq9c
auq79MNDrWaSzDZn2iAS0i3X5SNuzquPTeQubbLijj8=
`protect END_PROTECTED
