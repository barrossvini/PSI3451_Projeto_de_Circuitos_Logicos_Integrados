`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GVHXCsYuDbprwBWwRvIfjyvl0yiclPHiUBS6lsZtJQ6tNZ4lUgy7WRMBho3gi1Hr
Tx1By5UTT7rQhXMn+jaTBl7L+MbQgFDN+sHnjT9jsPS97w3PKcHug9YpUL75/CTE
IKGuR9g5XhFFU2TxtAI9xXBryb0Bb+GmJifWuovmu2FFeMFAp5BiSp4G/XL7FwZi
welfoAeTTXwar7shugFsQIQyRcplI7AAnv+BMfdWhvz7KVj10B2e9xj/bGgeeOo3
afspgyDYkUFC3TrZE0y8f4ns7DJk2tdDqQsQKHeAPCzoEyDVQWDzX+A0mFoccDVF
VwsG7YGzwBGq8zwuKCht+ThH4etU+O3PpipIX/LJ/XYHbTerAaVPnqCYE93201pv
TM7/Fn2EbRQ05bRP7mlhM9+BpwRnIFggPvuNPyEVc17dCx/2oscHmx+AQ8ZtmFKB
1f93AZMPbcb//zz1IgEyhGpo4rLUHpna99SycaWmyNU3Y0jDyCf4qx7RxYdRdraC
ls0rhtFPaq2O9HcRtaMRA/NYefqYLaPyG5ovnloX/dXuxxzBrSMeBl4wU1Q7uiSC
t5vvKn7OXA4VWFgQ2US+wBjUMFU1RZWoRAkTh4hwyQR6WC4ZUJVlyLuWpFjwjmF+
irlWijA8Kz42SvsFbuww8ToWlRhlYLKo8IOw2UIwHuq5RMET9bMAP0ePQSUzrcA6
5Cr0hGJ+UvCfY8lodKc3UmxYdmC99BKz6jdmQfkFmaSqVQIsSf00etecAiqDtOR5
Zvc/r/n8afBNws5FMnwD1q8JbnxU8IqbiBLhD3Jjkidj7M3bwdKQswdB8ozTEsbT
fNnydTk10ysPJSIi+XCxOPXT/olIhNznM1laYBqskj9FPnSxB+PdT4tfziYiK3cF
T7DfCyMuJj0/hH4vVdNC60lMNnbuItt3dr3cTa9zGPUxwn60FE+yUh4KnwsbpYP5
koV/56MpdjE31pBn5/dXmk7HGjX7unNbgvvB8MnH5Ivu5HwNm7xQ/Jkaz8N5Yltk
Ot8p5bTdkQvqi1EoCqNiSYfgKVXEfpVOyr/qZOrmifvZe9DSt2ZJ42TpiEVYErMO
lKvoR+ij+Y6GuVjahhdcEk0ZJVKgYcrf8BEEVRGnw38=
`protect END_PROTECTED
