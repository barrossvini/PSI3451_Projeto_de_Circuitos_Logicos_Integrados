`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lj+TO2eZYS9iPWLY8CzC/QtUFLfmK5XYgdsPN/37rjj0/qpL2sKAgfeg5ZyoqKmT
T8D2ibaJm3hefs0z2hEb0VrCI/5Dm6Bcujcaw/RGLPRaqD0E7upilcp2WNzYQb30
JXt2yfM1AzqpZf7qgHb3gyxsKzLmt01Y3iisQO2Y60jdipqHwCKHaiVGnZoNpfbj
Wrh3kgJHdqj+Et8y2PQcO3pB3RCeRdlITxOfD+gHiYx9b4eytE9IO/oqyKefVtMM
xPkJoUGRMVJM/NTs6o7PeWub+DeFANW9RU/KLxO1t+Vnu18ouxTXP2UkOd+7OV5v
aGgZCuTEPDxVQwPGPC2y9K7Rz44c2bNOwIM9wnOZvWvY3VIz2TQETYeRnPILGjXP
qGjpDNh/ck3ye5rp92nbEqjZQ/jvIBDLlHK6Znn3WvuJuzsVIA7IlH+1CBeQ3OEv
QlGfQ4ji4kIsdVj1FAhz5Y/Nf1AXt6kt3OwvOFP7yV9FAMO0ztkSu9HM3jyyVWNJ
RQwcZU+RVYog7BtAcOVeMBbH4SCNg4dgITYFY9haZt6x33oCkf0ulipMyKJC9YIf
5/cX3cPP5nmMKHGNWUpHlcn0jCnfjO7yXE6TAKp8yx4GvkHb8ekuJnxgEpLv8KRZ
NQnW8ytzNloyuiBFiCk6em4Nsoze6sL+YeoP6w4iczaEnmJcXZ5BdX9QC7BNkntC
fLjY0FCimDoVrvEJADK8IM4lZQqWQ/kqsyG2s3p/6wShJwVnjTKH73oloYkS1qvg
/yc6sNji/apYV33FWZ7gPAMLOBgVPKywUZVLC2M5O7kUNO+lbJo01vNYHLH/2gQj
VvxX4a/G9paX1hWEigvpTk131+FKdY1BN9m57G3ZdZ8gS4j3DnLCCJbkhR8bxjrL
QWNOoT2wipMKw1cvmRSSGApP1jCuvZ+v34Q2LJeewBtQF/6NyCwcTkxzPXLKZgdA
Cvr1zw1FCrYJzzV7t3NCNOzd0ig5Xs1X6IRXCBYHU7IAmhycSsWUo08SgpMpfLQ0
y4cLByPu2iHWgZvjzFvboFPWBrjou50lENoO0cjoOJa0RK2EDTjQMVLfnGS6q4aT
eulCYqoOMaYyBsDZ6F0Izst//mGbD0mpVuLYJCm6Ip/Ft8MGzEHG8StUCiaFe1GT
VKsXSiMYdXI7HhZZNxZErRfcFcJ0pN0Cm7Iohll17GAJ9ZItTnrychnD4ldTgq2K
p/kJ9Cf8wI2AQo4r5QX+roiv5l57nhhq9OLZYmBhRwTjzPlyhciavtO+pRX31WqI
lK5vcoRYf47Gkl/CNDiqhQ6IyvD1TRqaND8MeWGfGA2b15FqZC6te1749IZar92q
VF4FaEBkZ3u1Be3fpwT7TGoOjPHsny1iEPPxZm5bWU0jNHdE5L8JEKe23j40xvS+
H5gBjXpnnZ3K5ev+jPqqLIwDQzSWNsubVpqa5sevsA1MxOyQG6xTmzUmoixbZ4F9
hiQYo2J1zyw0lAV+xx2jr2Wkh/mpkvcZkqkBIcoESbwweX1XGpPIGL6zyy8DXTJa
Yv7SPzfbUX8/Fxl6yUw/AjbOHii0uCTjDrJ8/rv/ku2VFeWrjtOcGrgjl1FjvMnn
BmmftHf/sxwEh96i9FhW101ihMYq7XlK08keoGL+fd4oi5zzEmmcSjxFwnQR2mm5
k2lGkE9Hua+sb2d6yN7ppIBG7ZXZF38v5knbr6u8YWNAc390ilNpHmk1ZdlXPkqD
2eOTvXRCPFOd3tu5d4SWNQXGMHzyEpc5+6jAvEduzyhvpgJBXlSnLcpp2hyKDM38
8s+/vwOptNeD7HQJXusUDZdZtseiK3TT7iu4lv/VELzwNDOobGi1rR3+4pEiZ+UH
ByZK+GTgBIx6XStLg1XXjVLMWmCdXREtQGMddmJhDkySFIItrd9e/rT9cgVliDk+
TTBd2y1i09RgZFC4kyRnXB2tF/MnJI742uMbZf+whDiROX/SJdMNa12g6VZZtWTN
dpRdBoqoJigzrtsVb/cYvXqzWLGt2aSPHDjPznLj8dRj3Au64HrYIXgf4zj4fFQt
MRuBbutRX5t0FDMHN3MkHOVbTzGU/rH95ZbxqQvOgMN+9z/bHvCmblY0PC50EwDD
M883jHbxD6OSQaw8HqgRA04fGYkCQt3VmtTrfpmvpsXfHIUcGLeVEtdF/nRatx17
niyZixO0dMV+mkKLa0KToJwIIyuoGCcPnxPZlJh3h7VmqhluK//ldpFDsSP6jaNI
E2jeF7R2shC1yxnkBnWSV/XsV4TcMWmoiuBliHC/Aun29YqJhUElYmalYWM9k0P8
kHCLC5s4sfpLubUnljngylWHrzu49MWlcEqAqqoBboLeixZ7C7Vs6kFm3Ko45ZzY
KM+HAzcBhVqh/4+CTHF5v6Sv/5rRfeyLF/LktHig8QOn1ZdiGb5A2eedGHwR+bVL
MGqTp+dj1ydXcoqGI1KphrKjUt9NRLiRlDYmiR+w/Xy6fFi5XcaIcj1TSUxlVIVw
DeqJtbdDVMUPbR1i0fF6wFz1voCX/I5KpibUNBCja67phD4BKmcOD2r+dxS9yIcV
32exraQZYDQyU87N0CJS2nO4wlcgIe9KfXY+WOeWKXb0+bzZmoP0gSanM8JovUou
C+db4JVSfPnSlvdc/66DzJJXnkoV/CuVG7zQ9+z5biNQG5d7sBON6zeKcpxdrjBE
pJSF5rS/6z4PuJHNGXt9Pd8dPjhNGrmvPL3vX8oFecbk+oiKMfEguvQ0BtMzQeR+
44lBgjlUEj+G1MM00N6qTHKs1OOcpewBigJyfxD/Gwq81eq0GsjjlCmuoskzLGO4
WWEsDnHdTUWLO0xDaWq4qk7q6nkPYu8a9NMkWP0TrxJjhhGRMIi+37ZzK6h0Z0Ey
EBoH8hy2S+Em9H2ki0NCV2HOjwCfPsXdFe77c3K47SutykZkGYpsJoum5+nhn6KP
u43K8M7kgou64Y4SCizgg7B3fKcIMhb0r9DtD6KVH9IKrXFyLliqX06ZIp3/W0K8
47rG2of+S5ycHoqrHev1oyRiGlxcfCVnUL0IjV4Y9SVLJk3V92Jfi9fBnFzSsAS4
af6nAQHe0FjSkXBGlH8Uu8YrNtpkuc7F6SCAAaE//tvDmjutRctGFvbzhhiPyrUK
8A9uWCyW9BUoyY3C2tfqXd9av5h9j9pLSc+I0cSe96hCuRnyv84A9JNRYKbpf9LX
C47knYDU/mlTdVsYl5QX43H6T3plBje6XMPxcC+uosSfjW3orS+javmAsUbJFKA6
BlgzRHImdgBzjJJmGovexurz7GTyQ0FP2E/x+bFg7QqGMu7g2hUL4zrL2QKfFCRf
enihezeOb3ds4UAtQ5X2bpFzKnWJPb2cLX2G1oTaM5Bqhg5vb2yLZEEm+mTxaUIq
w5BWWw5DV2rLgCkgZSOxGUiMOqc+bnWaJhV45t28kvvE2aLKC4emjFIVhP9+9txi
k8TpJTT5QUvvcpxnDxzMO7TVKdaIdtsoulzzu/ILIbhRXkuW8SH+HWTjxJxdXoyp
l0s9kz6X0vj0o1JjQgTtrTEO2JTj08rFvt5AHMIMmIgopuXy7g7eJA/qRzwAUMhP
s8kvqwwi1pBt/11HxcnWkal0q2hsE4Az3XAxOBs4wJubTnZmIZSv+uzQccBK34mB
TTVkt5VzWebRpDAFCPS+gvxoUAdYNPfkbz7TglMYrxeOhUdilUaAFzb9FIa1GevE
30yJEII+JLuXhVe5dRjODzAR5pEkA1gvmYnXULDIsBrUebAE+eMpe975nMYXgT4U
Bmy3ya64pXKW0vkkCkGpcoqlnUZGPN06fi0KWOvFuqnCui+u0v4mH5I2rVOFFOc+
6mwdlQlzBAFLBM6FS9LuFnZncTGpOQAxOx2G48+cGIUWefg5CYYfARFSU3cULlIe
SWOWbZ74Tr0qr5bTcq59/67UclHTCiJrM6Uc9iO6383eZC4JkVThOjCQi2+QbwP3
gE6LruNc/ijHmGeIwqBYauUgPDh5dcrgYsk7ik28xWTpLE0M9ZPr8HVS9MxQL0QX
eSBTCR5phDHCIUdMFPswX05wafQx29v7vHgmf0SSOUrY4sXYNXe7QN1GfveTUJew
82jWdVSRiFuoTli+maQN4mAu7qoUjn58sI79ZdZjPwWCK0sTK7HIYbpJvw8qiTra
VEqzOKSlAMYAwCVYKCiBEtQNkBSTbr+THXvRYtpQk/r1uDhYNUEjyn3yy6ZvWhgW
0HOapGf1Zg2EBxiXOGjk9qHNdgz3F50hP/BtOuN1/OnIFdGQ+TC/r2TmJ3Auf8Ep
nmwRJYOPj/ItFVNC4FU5ctBwxEOUjkHFJGDxdgbR16awCDiWgAKjwBAufuixtdz/
oLTE2uxhsHAAzqwqEp2ipIdF+sPFGGQO/45aJqPw7HlOOiy3i9UOR+PwKvYBvqld
K7xMfMChqJBbVGeQ7RqdgPv7bO0e0gHjd5NMk2B/1f2lLmgsjudCKdQepcRWUgBf
aUaVFRVR/piKVaW4A+eWrs2SkxswtF1RlQ+6AWaz90YIms+jOnCy08gQQSvkqzhb
MbDYWk2aRTfQRC/a90C3BXcN8J+EAs5CvFSEeOvJeQLRyEkKR3vvLnA2zeIxAhCV
DH5EWkmrhs2H9ZSHJP+efeupFpkEz8m+hYia/P1eJwtIGrfq1xzVrgj+v7YOoXWY
tAvOdtwgOXartrliQLWRQ/Lsrqa4pLKf5ANpWQr9albZoS+Xv1XiUuaZceoIUj6T
hDwyUdElTI3XwiJtVSBwa1lZmkn4tthrpzPA4EGQn5NKrKEqYOl6VBFu7FoWMIfa
pX1OuYxMBm9wUL2w2niBKnlkvlaK0BBWSiaMcpRBG5gGn2baC0HJmue0MrdVMB1H
RjXjO5ckzOOI8jCtDk1fTvhDM4/HCypq1KpKndsZd8mjmDjLE6zrKNuig2C8/hbT
UhdNmCwUlEr8FIgRsSETite6K7oE0WitJdDDiBo3udjWZ6Lj+fUUohYwHWhRF8Pj
5LgKECC2Ocs8VjE07JjhOqUhoEHt1WmMsgmKMPuCZ50jBQgG0ejVabBMLJ2Bfmf6
op91qQ5Q8lG1CL1+lLYLoryA97GEj14OvLiq8zR6ABUlFb05gD/rshtRJilbpFhS
/ocTdSZ1YQ35bAlWowIVs8ghde/RxDmtIEnytXUJ96SBzLO7r//c7lfmUIUEoT1J
zyMLP1bp6Yi0k2zRgUsI1sL4zfjsss2DgJNKl5+0QyORweSyKkjr59YsdlKk/Q0V
c66TgZLU7En0NGVfBIheNPxEDiRTFWXe1Kf7ewnplCEgNrXNy7eANUGCjLmDjBjV
uAOks7fVIjFMrHQyy0Px1B28x+eRRdy0ghE/EF8UQat8KKWL2RpQbPBRjallGlOV
WLSYeuc+Iq3nvJGCDFVraWWIDKSEIjMO1OWZGS3J27k3tBLPO78BmmXBhkx8WRAv
qvOKHWw/X0hnR1RbORiZzextjy1k4+5KSeUXxzRn1bK8nkVpKPOsDn9wHM4dSwWn
R2Co2tGUMaUnHQytP1oGR0/3w+n93lVkP395WpW6CdBQEhOMKYrOdlvVHujbZ5xr
5kUTO2mRSvbreGhaXwNG7BKLAvIh0EStFNYTBXkank064Dg9aLV3m/PrebdJJEkn
WIoj1vV9SUXSJEBrL/ab7tMzIsDy28K/SZj1MAbeHE1NzkDm5dwm4POTTqs0sCXn
0vucXZzxnoBlO2gm5egnHZ3HDAQmTXDk2UcD/8SxA/D3Toq+SvcaxvtCHnNdFh5R
DRJOyyDV3pH4BT+Mmb0J4j/Td+XvIJgdkUEd6ymhYXfNG9xmQtzbFc3ZWMe4MhAr
IZzGrUTPOO+XxPc1oO1aQf/9kLJ84QdIX+pMrivWgoBNSte1k6MTdrHzikLhc/5b
L7nHDeaI8wb/JUpEAZ4GYNKLNfIG3Hlv87V1wGACJ52DTUqVrhChB/lHb4O0uzWE
FEQ9VwHWb5qmmTGNomGC2ulTj9zCBuatTgi760+km4vif8J+3eUBlZ5sxvE9MWyo
+9U0fmQshZhvmt+g2b34eWsJZ20EUbzqi3xMvBJMFdMaa4xHiBk2BRlqqNKFGI4H
XtPxuGasuAEhU9rjWzSzVboDbHJLmPVMygmEYxEx69CC7qmvNpXgoEfxELl31Ny3
DK4vlOYXK4zsD/XAnHTexLyRj6vsCoEkro9j9qnnP/ibnfVsGpdQpbRcy1JgwUD6
/3snghd6fZFOfl03a6Bp+BoEqqXvu2dcHiJHZqZ9RCbaJJ3cYLGRfyLTHgEj1pBt
O/tgx3MYGWepeZAa63AD2Bsw9Ql5BlW4HTicbXyeKmUKoctmmg8FxJ7G0yjn9WQe
SxHbiZuJBpuzaoUhH9p9KyXmeARqWBCnCU9KaZ6OltOAUJjvEdC4jDzgtEbHSVdU
XhaKKw4NeORjTMLdmq/4HY9kA02aTIfYJ+38/Xz5aiGLOCXEXLvWlpgGHlwjxErA
m5cwQukpzMsQM0Iar1JMJ6rPb7WjWy8fxGT/K87V7VS9HfEiXzRmpZUPty4FEgTk
tT6z1UD24ZIJprLdO27Ph/sfPMsW1tv9J2rP6TDXzo3RxN7gATUerhnv3OjgydM6
H+OSRVAqdL0yr8tdRKbaq2Y54R0ssiOv5BDr146xsWKZzlQd5NmStb6fWJGCzXQ9
EWyMFa5KuS8UOk0lkdBA5AUNFKvsXvidXNu1XorZDzQaNOBmVKL/InPgFLE3PJaf
Ba4SPZZh5Tena7Tqgt9z7yDNfFFqma7OfQmftm/Pjq6Irw8KBZUPKuTjyPlQurA7
NS3Dc74/DZueTYBYskn9A00Apu9lnCw0HRuJr92beVfkc3RBo/KCS2aCkch9d5dM
`protect END_PROTECTED
