`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AuvBF8UTevUXSWW0yx1dh3HYTBN4AWdibXwGDc8Gm8Aaqwm8/FnZawbJq2oVSkWO
1Jaz7+vGLvP3pVNNdNPLZxmTUv5b810Sf86Kmdes2SMbTAXjJEEU3exN7J5XhAHn
4Z87AuvxZ+qZqTFO04id0lBtQyRZhzLSsPSsOG8SD6YS3GHJjl6rj8hiCyjT2gFa
5d1hJFxDpZaUv2sLLhu5AvLcb3X1kzGR2a3EPfTfLwGnxeYobil9O7gqYVUxcz0f
maM6G43HqXDu6SFHJ9i/wDtMKia5ues/KrbeGgns1k7YDfrWKdzVMWWj0mHiQzrU
WOWZ9fdn4GJB70SuoAebyt1DR9etf3HQnbQw2zbiRceHWK4oqiMQZ67u+aKnjtEz
lwWzWwdkA0+udsJfyJBcd4XGP50gooU+tWn9iDBnWpLfcukUXWsfTJFruiZlZIvi
updZSB5xjc6srQbet1jTSZimQwF33ZXfwsN9BfxcIrntmaVHekaTVVxRg4/rOSYb
PbIcoOcXFJw2NEtNG+8g89mEugVxlwd5bZ29ykRuTA59Np8bNXqQ+UqXI2aa+u7K
o7FrBhsyzJj2f4VJ0EQIgo/JnbI+jyKerd+WiJZ7MRTdJMgikDWtIPEu38PGQFdm
BZpctdpAdIXYu3YRgihs5MzpgBVOd8SMPRhey8RJ9pCxY7ymyAzzqqQv1A9rjDLK
IIQuE0SMyDYJry/FeEljBrgfoq/rmwtzgn3fNj93eEx1671twyuwKMwBP1xUydVe
ZkunxerpcjXQ/FjpuoA+sM+5cLk23YTdA+MkdGfkkNlos4WKOMjIWUdhrSco5KAu
Winf5OoX92Jd2Jdb4Olv5ZqqhOPkhLNG+YxQK7ezftFHJkfVEDL9c8TKLXS8nSwF
Qj0UXHr1XMdHUI5ufDQJft0SCYxLqgiRtdd3CzY08Nx3Y+4aU4MLVOe+eU8NZoIJ
WWh3K0DInO5RCDYkLOr1gELcZkHqn/da5wH7Imbf7mLMfrwsxK2I66ryEqC2LeBb
CzCeDqcfjIQP1DJ1fSJLow==
`protect END_PROTECTED
