`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yea3xaxH7+HzDxX40FoZYHNXJ3FXSMVfu4tU9aub3UQCxSC6pZjZFt4ShWnebTa0
uTe5KEdQC1SKgxqax/ASdoEl6dVFg+oAuv+qfbbzSEqEf/R+94ZixjjVydQmPvWK
0CVJMOQ25aKCdj5jZ7wDR7KRl6d4GYVYjco+y+pINbzGAZpPu5tliRS4tRwzqfi1
9816gprOS9shvo5tGS0QPNfc2GJBlX6scCZKaPc+KdIxsb0V8Ke8KwHz457RFzyw
Tl+dPSjTOuf7ECfJ1Tayc3syS7FA0FC0I7n84IgOAPpU+b/R4IGAw4RdXGtT0dNR
x5ew/krRrSzOqFei1hVRY9ckjtDAN09xFMrgITdXlzF2dc7L0qnbojod3PFBvKpL
Gaar2KdoSi5j8kUqsm5AKzKAcy7BWqRnafrxzJNUM5NiN0d6uYt2BJ0/Hbn3LJ71
PXTch3U5oISBIu9B6x3gOfx7e/KBNVD9jTmWOlVSaTNNlUVMKE4EDu68DRHdnD6v
UsBY4WbIJqsIndjMsgcP0o1RGwqzTWz2e/roHY7BP7NuzZ9nyennqOa1+/F+rt9n
Bq1qpn+ixZleBxRs5u2SQm8xLRdlzFPLvybLDIyx5f8GDt+2LaRIA8U+UwpxAJ78
0n6larCEMLuSXQpnJ8hb/BGOc7eyqaei85p21Rw/YVibbqemcXcbZgaQW6mDPyyB
y95subsPDfW83fFSA6vj7svqzDUjRtHerBEzKn+oHdLrrPoA80x5tCgTg2XBUZSM
FxbuAD/QjcE8tS7A4azEfKoFS00hYkNajVUgWr2RN56IUfnKenlqYcqqXbLZhuKU
ygVdCgtcBdu0T3wcM4lRNnEdAb+b8i9LKy4SmpbQLTusTZjwuCtkI6DN6v5D9G9f
j7msfYiiFOv9atVkqjQX1FVYFf3X1HOwXzLYDKKtczZ3UW9oZZdi0GG7cM94X0u9
PEXXYw1oH8LKPR4T1WtvMI4cP/JG90d80F3E+/VX9nvUpHAHPSk7Y9sgTftwMsRs
6fd3OzL9Wj/pxywS7CCeum+sApT0Y+vFCqHuLyc8mHSyFih/Z9MEfL6wD+YZtF88
Z8VNfDNaAkBlJvjjlpE49yBF/ri5M7HTZZpTsZbJhU7UZ+px66KilUEs0CWlNUaA
OEi0e+vIwXBoh1PgwmgyngBnICrnMB/h6VE8czV7g6UGyE3A43X+eA1NFKtQW6UD
OPngZpr2vOru0thGC/21v+xKCvz3KjDBt65VU1Bdkq4+yKXVnGwBicHfuBQqE13N
Y0KR3QGTlwwSZt3PTc5Dk66ivDM4NHOyHnCl7vBs3BDf00l+uRtS+CQnGbb09nOF
lWFESGFV4pLqcZ+AdFieEZa/9vv6DGmUq3dK9ektNpFZI35WUaHZVlO0yHd2eC+W
DgtEiX0v2QST19A2ZIc+0m0BSQxE3AtEojz4Wra5EyPud+aCUK+WB2BgiC7zLKj8
`protect END_PROTECTED
