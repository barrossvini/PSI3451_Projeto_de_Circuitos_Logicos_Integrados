`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mnO5MqiqYzpf2hCn0Wn6T6Os6/2OOth9M2XEVkOEko9OEnHSDBkJ1zZlbdjtWegH
BL9zJOzMq/pF30ju2UA68+lKGwqWi8cIYAXzLszXKL6TckosMTq4/6/M3eDQOMNr
ue36boRG3tnL7JQcybs2LvXZY5A27/dw5zBErv5nera7ofl7hZ1ak8RHayxGPyhL
Dfx6/DRlcGsyGg3UKhQ5Bvbos8OvYQZKL3B0ESJE5IfUaEpgGQvpFo6yGIfjc7Zs
Dx++0M75M6529RbxPWJDY2VVRq0EYDXKnafMO+S7DmaoQbhiE2uNJuqGj46dYLyz
DxAsRmzyUQZPXCnrJKp2aVcNLUpTSsJmOD226OCqpUZk0sqm/uGV9ZYBR5BCatqa
7iPUwAWgjjdCU81q6yHbSznDvXP+G2WNApSzpVRCCTHH1z/wYHNt/A5AdZaM0NTX
tmeAajxAj4dT5uDEf7vZUta4ngx6vbczdyhEGW4Q/uUhqj8+sy+aBgZrHZ3ZgEVR
g3GS59mPgP6j5mFMJrYo8ZD4LusyylUZ1NSV+4c/gqb2ojTyJwQj/3MX2GeRsTvo
WmCgA7/wLL9wTQ9WQ/Zt/ptzT0C0u7bj0fn/0Xb7Df0Wyq4DxNlKxfxyQxFIbXry
suE60e8zxbxDQqlz23Er7whDHPHtMoHHWUDriC+eT5HTgJ3+HmzHPhwCHSbgRdor
Bcbnmt7UIUY/6agk4lydZmScENRtTRjcG8ASyn5rVGlUmldcAr3MbesLzG9vOalq
gr4hc0qc595bUt7PvyN5tgUa4bGTjKvAopjCRmzymMgOjvZlNJXLDogSMGpfTSQ/
`protect END_PROTECTED
