`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D96ajrv8Rqx+dyqVqPc4cOIADnnJu5qyKVdbX5JbiY1sGjcuCzr057id2Ztgy/1e
B1LEXtmnFyYgDUDAZfilY3J278Q8YVSfpL9tBz1RTovtPnF2WBOw+74v8pfIHF2B
N/1DwYGXO0xmVp51WTCwRjSJTpyaNMLnK3HFehtxUL0=
`protect END_PROTECTED
