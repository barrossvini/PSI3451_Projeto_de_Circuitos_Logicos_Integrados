`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b1QXYxcJ0ZrIm/IsTp/bpNiNs3yP7+jn3UnWmpRRfh7IGP/W/C1fcvRiF3h96HSo
QIXMPh8QdVs8yb2arEMp/YXEyxLJ0ABLu9itD/t29h4wx097luAILLmLEcGU9Bcr
HyHLhg67BWQLymdJhgOTw2v4Z/+Xp76f9qM5YcRCnT/uFNgukx3MTBgEUcDttCCZ
ZblfWsHtvDxvv0mvb+iYpHNXw26659gSioapbRzOz+K7XFHgbeDOFcPuyJ6NPTOa
ZdwUjUJIFdw8aphMEIDkWmoP0Z5iQ7VBMDL6FgFFBM7B0ut7BO4A/OdILrli8YG5
CxsoWTncQcOFkQ9vHyO50f/pefKBqM3CtpSSzyES9XAAkvFsvkoT2Sf0Rot+lVmJ
4XaZhmiCzuE2+y83uZrea9K/ahOa3wbH/9zB2BsKFadtLt6USInhhHPaZ/YHUDcL
mh62c5JOgcLyAJuWt/JzCRsNrFhcAonxvw3e211GOszVbOi8RYvQ+zHDu2IaGzNF
P1KerzdMM+7W5y3ky96LWk2gd5Qk2gnCPN3IWlhnSNPrOvX26TyV73dhx70LqPaG
yGrlONUemqv6Hl5pQWVU5Jen7QNOb2HNr3B5R5pOipJn35GQTmd4TEAr0Ek0DB/m
xCnqEI7BTpJ9jNxjf6DSHWL2fNkpA5k0Od1PNs4nOvKL1L5RH4K/Civ/oilAEWXd
7ivyCA7p0R9inr35ZtXmwQ1Z90SsLEOWaO8djM2I5KzETvm5TowMRgtxDzaJdpjK
oPzJo3s4Tag/Psj7a3EVA+DuvQQ9YB9WsDy0vu13LtY09Opzk9o6axlkX4dKgaFL
97Oep6xqJi5SoFADrOnv4rDqADthj6qoliUzAyVmvSqQLh0p3+hQfB3T474St3u4
SpXw5OGiEvOftHxkkvr/SYjuDwZh6viMc5HdYMfB1E5i0gl7w48UsvpAPjwfLA6y
jnWAAa8qDf/Uy479JgVZUHuz9wL6/0JkxfR9KhRIjg2irGEmcowX16irbHlFy68u
shHxagdVKlOFHfEnAFp8SGoN5CmibGfzYnBBCXp8mwmds9M+OCRt413pjNDvda8N
Cl0WRKKcis8A8n5LJ5deLdB1V6pjYKE48uum7FnLM/iduPmQwGuKRYJrkKCWZj1L
uuoOhThmaQ+kpNvjL/5dPQdxkVXGoSNpdkU/gj0mzThMgRqxS3uI9W8iUxcyBbzQ
GqbIeZ2VBiirImSm+p1SHePlmLeO01JmiXRXOHXa6wo1iW8kSk/CxXhszi+14bth
xfKjgaSeLwVj4NQE/sfMtyKluWLvLGJyl6hZuBIKB6Rki4TtowjIWmqcDxU2yi6n
s8rPZHn/qZAjNX9iSCZEUWVarEl3ipoD5yud2xYPaIixHE/0nauhjJpwKhFj4Pj3
`protect END_PROTECTED
