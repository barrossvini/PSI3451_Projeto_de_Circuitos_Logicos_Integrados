`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pH7qmry5IOdPCu7RpL4AQvzvJlnnWtTkz62HYuY4v1KqFXvwErVoKuJ19FgrAvWV
C3HFyzgGsBgxmNFeSgMRCr1/W/2bOchzI7u8WW+wbqeCa0RchKVOjxgBmQS7wD8C
lmfmYGJz46oUw5iEhsrOgqeIiKOA5f9Wpm8dQ8jefc8MmcReZHy9l6flCKc0Idqb
B0DBwxAXaILooVcM3S9LHtaC478UKfj1n3iYYyFxBaOte2lh1HBN0C4vBSvsvN5Q
xMc5f799gKL/dt+CteOQRPY25ura/i/wAEPjOUimFzMxZSS6zM0eOKfggx8OmOdj
Ao2bXlS8PZ8dUn0AyOngP44Fv5lYdrntgbF6+Q+Ug5oGaiKdtucW6wvbsOZD2Pu0
MBxHgaiY5JqnU/uDQL2h+vnVFUjYUCGOYn/UK5BuhcPJVHIkR3Tqn3gecBZ0PhjI
m52Wik+M6m1bCq1JwhNQUgAFuj3b/h4ZiKnUK1rg3mQpfOtNnTbLaK2sAyryvSlX
BbYWW6iBkYSiPVpjwhfvUHNVZbuueTYl8/5amTgpM+o8xs326K9o7cHC/kr6mfx7
zjUkWFOh3VaNE5QcYhsdCvMCsMnns+xZEAWAxSTUBzRk3Fw9/g6CdioKUK+tfZ8+
p38PrROWMPnb1kgAwBmaYr/x9/7rJPJBr7Ul59H218hsSjoEEU0nOGSat6p2toIk
u9Rp63dXHO/VbWzVnP/Wt73zVQfqX+C9sXTu5UqxkISa2HVEXDY+PDgNlcN4ZIa8
dfxLVRtLndhDwBkyoRKT7ntdlgvf/g4y298CdSBRMm9ytlNgiEjQQ/4SwWpOQPuB
g3kmGZ9rzNtE8wMUfb82/Q==
`protect END_PROTECTED
