`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLHzCSxLYKQXNBW7yOxRa1YXpKFbLWHUWEQyAY5Y0xkxr2PfjCAK6SVHZwA3FxSC
bEQ/oKZ/h666w5DBzB9ZQVe/tMyHF7Ce5FCkL9at5B900c+h+xuXPlWk5Mbe0xIX
/xJPn7ML+ySAdQig3VLyCrx9XE0S+guicjDdzZSDiRwi7kMPFseSutgsaBkfd8l4
m4QIMoDQRo0qq4YOfcueAB8Q1MIATfcojLrijat9mnzlH0OSBryHHm+HQz0XhFWE
KUGKGPPaEKz+nxKlDH6rE8+SDBPfUQmfSUMO+v8tV0QDlK/NntN4SJvYhxHZS2tB
IGDPxJPFWD1Zv3AnW0UXid+AN3XT5VGVUJhELNzlD1GRWbHsjzuz/3Yvl1h7OfTe
vble/VGvW4K9IcWk2C0vmNuA/CLjwGnhY/u30gk7uCGD5bEdvlg7FeMeOwEpZe4r
3d12YGRBjxNE7vRkrpbE2q2zj+gOKDBg+kfxySKjOBAXzHhOEfokIWMjRB4W/rBL
1WKGyS2WRJivLbcjUh5dvbkRsBJfiErYBJBap73N6B24A7pq2YFzzoAADLliKIjO
f4RdIMQY0cEgQ9yerze2CqW5z/Wr29fn4dCogBNfiIiUvfAOYMMyAZpppvI1ybFA
4QK8QMdiJFdG6ibRoYeeS8m6LQnzrVhxAjIFz5c+E5cIJxYod7Y+UwPE8dsfGh41
6YdW3M7Aq+XAiMzL0vrCbKO3KYTl3UIQAHst7h64cyVC+HpcagIpfOEmyq+u2yYi
2yyiWhYJdC4xJLy/9BURopr92mfyVCBTbBlMip4u4rhprdok2EcDERq533Mdhnlf
MasbbFkWKzq38OAhfoA7h/3hQVhOC8U4pcTnHXf8x+Rz8lOTzlaf3cxuXKXCavV5
FQbNy9tZREWEoIpuqB5vnNLOrPbVb3XJMNihFv8KkT4JHl63tdmbkvmwD17LFKwk
LTR53tg/f7PYn2iab9fggt6dDBSLe2D0wJcfd4aS2NXc9aTxkPYh9FKMZ8fCGf+1
mRxr8TsADvhgnUMua8aLHv+Q06pLdFrBVn000DaUikYI+AYEDHgulVxL3+DcKiWy
+src9ykI2ZckQdMaoTwG39PtGF0biRTLhlazwho3w3kkZxf0rK+S8RTHsdpl8qKk
fWWOCT+pqAXUIMEv6zLs20W+WPYoMWeWJuDbmbZ+XAsRwqhDF1tnslmIoEnDLzwx
Fac19K+LgPo0xQICeCs0SqRp95sIoWNFBlWdC8h7bdg4JKzLG4o1XQXPAKS0L4kM
Na5urByUkNf9ssvzwoxrYuPb80PuNb59LJ8a9ltA6GsHKAiXe6NdmzG88cplFMqg
LLkwBqD3PDdyx4YKAfOBBGeGEh1QMOp/8+UAFNumkFHg/Bcn2uJvhfCHTNYf/2Cx
m8OJ/PRa9TOjjYVPED+N9szRAU/Qq1JKODtAXJFohzWgTVh2nLgiKVuwfL+e2SWy
W2tG+g9YUUAcPcFGq2/VC0SwA/nzvyi6vncYsRvRpfdkS6erS452HElTRKUrb5bq
1UBtyAGhR4BV7pOpE9Ykg/spRsx39OVkuf6sB2guNhRs8as4nh59rZ2yQ7WlkA5A
v6MGNq/gpLLE15t2pRhBKkld0Pln4yfnMXuHHcVNAq0lwJp7KeaENDQYAziDnpZw
VRNEV01HbYauqnFcrKVgPV9EJjphY6aizDlPAj3Jm2GCNiqQ2CwddPEzkWeVCfh4
6jIjwslscGjFmyQy1zKiWoEcfXmqMioTh0uPNAJU33wGr8yRXwo771LD3eM7wA1Y
r7KfUevI4RZDKPVEQBSg0rqAgp4xf9NNsc3gtvfiI6I6I6L7EO9pK3mmZUnAnIy9
0qliJXlOnU4vxKrGpneSxQalbg730ebd2W0ogHhoM0IkeipxlUNk0AWJaa4PnapG
90O47MmZ5tk0OkqVPyvdH0WuTaCQtMu0hS7zKyxWKVYCtkqZ746lfvPL7xroGRIK
uF8LF9rYXgat4+o5sJWO13wwemU+/1Ay7q1lGYXKGZ+3OqzBnDiyPZ1MiTp401uM
YIVdTOy9+oetVWAUFdoXx83t2s9Wt95uSdAdRzbojKWB4Bi7V/5lvIlkUgCBji6p
aa6TWWFucWg0Lwy6vi1yt7NJVX1M1YZcKkMa+zpCkkFtpBn8nmWetM0SpgD1FfyD
+FmDkeSW4MbCscGHEljuR/C7Yt4AWbMIE0YnjnRBiF0VWrHsB6eoCShANxHfMDud
Z39ayNx7hYO+Jiq1kOtgoPLSXMsHvdb1ptnmFyjmsroBet/gWkMLX3F4dYH1Evds
rOfybTNgSFAigZD1/HgXebaVuE14ZJcm8jWHb1aWAyscNTmAzda8xyeZTr5/NJQs
J7it0jUPfUkGxoIqWfANEzSrn2oNkHXsG70TMq2KYzFYNFk3I2774zrcIQFB627W
GxEWWRotozk0rVdYFpx3lMKAMjNOKAusLwbD/jdkV2bA+4p6dIIDU+N6eUmwf8pw
s88pbX4cFKWa6gKiCVlIvmFMe2Caiq66oM0mc1CC2TqMQoR7ZjnC/jG1mzM7GCWk
5kOG2JRslOIGBk/oSbFqZSwQZfpQ/sqYUKKfpChxGapLnpPhjWuk3okg81+TN7f4
dyBmEvjT22ASw0zkJcNTvVdGiddIt2kUhj1Q4yjiljt35ZC69KbJaEcRBvWykI2x
XEVRuzEdplGTsCcJuRU7hfXF4Xy8n0S3NoZu6+uGbBc0PldTMZUNi/cJ/xckEPF4
PMrbzUJ6rwMpUu5aa+fJmAtgC5yJAfWR2m9pZqa8pqeOkp5sp3ckS4htthyv/3Hp
QpK75VXAnFBE8htg9zTpJGxC389+/id2TW7BeG9eENJVDfGb6HCTiiaLgXdkeZoo
rx6w9lpH046WC11lMhmTxrcENg+mxQ8TGFuUc0s2tGyVQcQXhVJHzadO5NbDwRnm
s9ut79mTFL60tn3OxDWl1xLjhqocntwTJOalKeIjYWp+1hS89In/muYvTTckjhsZ
TuNOS0wurCikV4jocyLBeQRNYtnezLLcmGN6e6cuyHbPe0jaVHQMTeyQvoCCu9eG
F9Ir0nuqla37PaxiL10QXi+czf5s50AXYoXChvwdzSqq+0RNOmOuKvBdsoYJ++Ir
1D8Y3aenSGSKcxz10mvvW1kn0io0BiKogQRQMsdGxc2/d5OypVxvzraieLayVpMI
IToSBVlt9S7zbCX1GXj44WRCop2z4kJdRDYJpYUhL7IjDYG7Hoe7JuqxoXHPWYNS
p/zkJjawoJN4bG2wq0A/KmLgyqBQ6u1pexBrvOGCNnjggpja+nx/0vHdvzM42RYq
/VPqXeSA9fT7NsqOfd9yOmevTkKADn9DV4cMc5/nPCBRt4FGtTc6+8+95jb9wxZM
8EMNRnOdT3JLu5BKnat8QIYSpH+A6QXAsFhnxLvFXVkHCmWqVaYwEUzvLcxGBrU5
lqknck7H5Y0G1ueG6OO7XuIvMbTHPXbBM3P562HN0u4cXzK+gA97kPEagCleJPv/
fwJlNo9lAkex6wGpBF/qXMA2nDXDZeD5zbJ3oogXoe1KixbhDY/Gt10BEnGlBEfc
63wvLnsd36z2laAUxKTtF/dObfUnI4BlbEcd2Dl4JcEgCn0n/j4s1SGkmIm9RIeU
SqPvHM/FffTwx6uCXHpEEftDeu9w33XA7MbVA20V8R/jPFjy8lWrFNoT+/ZPfQR5
GIagSrKw5CH4BedrJ8UH/wWtFUe58BiysrzE3qLIzkwiSkeb85lkAYUgvSA1VbPK
vE0Dmk5SSVDHtCBGI8muZDqSGc3qmzj5WfNsMSNlWif4kdSi6x1BClEBHQ/yiC+2
4MhajripwzYo3C4dFphHjT1ChkQHwpqdVcIvz4NrZ6jz02vJ6WLBuKhiM/uvzSnG
oRsbldEP+E20xTkgON1Ts7Mfe64OuciCaBApcYgHxEDSvwZbkaGPqbNunFdo/5I9
agA8+Jp8JXJpzkhOTVBfCJxmLJg4yuaMHgIINYski9zX9KHeNRNzghSNxRska7VM
L4VYgJk0xwirHUck/MO3CwViYn3KN3MBkgbKnx5o7NtWIC/0vjirB+r6Gn5mX4yR
O57ZMrmTrUtztTgYGsg5gQ1YFY1zNp7kVJc4eaB00GcuCw3FEOvgaaEUgiRUcs2q
bV5Od7SIhPoCEDzXVAiC6hJt7fw9IUi1t3mfGeTDoEZbBJO18R5Vg4LqOPIeoOBK
h0w7w8k4eFK2x1+p1SOKs74YZ+x3DcanCtNgPGWIIyrxhE4XZpPZTgIVLHQIBuxa
N2/cKXNQQT9sSocsXeT+zt1JYBWRkwmuCwigKaEJf/cmJRZw3IhHwVUTb4aUwOZf
gZMq7kWBlrQe3LsDWCuk9C34oCb0K7vY6oCs0gCAMsmqOzEmdlaNJ5QpjFP9xsxS
b1kYhF+6e/SaADzHWhP5lz0xd3K924IRAl2BOPDxHqnaSoobIIDYkefss7on3ZGC
j8+z70oByoxHeOr6sRd1snfcczC9FfVPbB7d7QsCIer/8YVP+Hj8vFWtcWqzRns8
8o7587CMul6QtgbBOf1xWRXRUqbp/OUy9S5M8qaNienXUm1109MlD1XPvqcf84o+
t0ENJubMn7Hlrqoe6kqSluvxNuzpjRPt3/hPQAyi9vvA/hHpAmHPJgTV9b6sJn24
F54zbMRe+c6PNRHHqFnWGruI/TOPTZGMkVXvVj5V00C4V1A7Rh7nrf+wiovsO6Yg
c3IxAoX3h3CLe1FLeRc8ot8y7rxCocQfRM27lLywAZu6kZxmTEWwVzAP1BR7tV/W
tGh3ZV42Oj5p7jq7cM5KPZvciPGDonh212RzLEv9ZHscnZhCPi2kXQO6yNrp0F0p
Kd+PQK0RbOhv1/W2gtiIpjKimXNn/JfRzGm0rd6kQXGJQO7w9ipfhCD2u7VowSiV
6cAOUcVHplwzOStFwKN1zA3Vo7TgX6V2u83+Ac90EUL6GechgCCAUU5evsCegPtJ
iQFmO3HoVO+nB+q6fqxWs4GzWTDlKC60tOqiIQs26kQdCwnXEFW9CBEmLLShv5Se
XPlywOH/cdo8RayRUVjwuOp7avddGE2oCPMmUu7N5g2pmYH8Yev21eIItYQerb+D
M1eOyyBot0uCTlBqm20Lkv8fUaKfJB0Jjcvj7AVc8ipKXVBZbc36q6/Q+dWiAR+w
4/eNug8WNKuyFbifptRalwilDYytCQoTN2AWNQonzqXwKxydiPtyqImxsM8wdOiN
rkvgB3ezxrFe/oExwJRQl1v5eE1w9SFU/CHwe4C5fdgOqj9UE1dZC+GWbp8pg9HQ
0mfiNSioH4ZgSHUUG42aQpzHpyM1HaX0/WmCvJL0fckj0XgQVkb+MNIQPCr27Fnu
6JpL43xp5Zrui+4YHqBWpak1XQZFVlBI7ihXFiJLSuxZAc1SyGc4sNsah5Ot0QQL
F3yyko9+9+g70okvTjuVeByU96z+iREu/klQwb6467esOK0KUnJryGklDxInCNk9
2qJLATdNqdNnGbCf3SzMNARmq79rGecDqbGVudnFtaGGA6VGgsJni0And/dUZJXa
Bb3ePuPM5qdeY2dYZ2uIcb2+T8mdeSFm177ctOX/YM0N5TNkJzNjnnMRy6VUJEVy
kvcQX90aqTVJf7UULIkvtBYRK/q4nkyFxxjHI6fi4EZddH40R2OUkDMnz+lURJl3
TzMJW/mofhpK4RvzG3nal+vnoePuhQQ7eEgtXZAxbWkLsT8/7cTtCBJu5hWmqvaQ
AhzrLOZ32l3B6LXi0k/yj45nTxbDj8wuBMH9Pbhgxtljy3guapPTYYrMi+UQsDAi
fNMsNjEBwLCaZ+xDSmqwzxVo+BQNDkCehgwxoK9sZFDIuUdRiJMja2MrVA7E1zMi
8zSaR437+J5X9EwTdxoMiYNbcFeGWIX5kNwHZMQyAzAP27bvwFf1GFdFzInI7BeQ
rv5ACaqkh7JV2R76neBFAlGXHGgw2WdHEc+OKbu54qDb5h5b/HhEvM7uXZgVDT0+
hxVxtCmtr9OE2RnXdpPcd4bPm2EvkBb9D/xrOf6iWyQnp8aqd+5no3XpQChzaPGe
EkTFi8e+LYe9mwWHXiEmet/I35OmKtrZvEgD8rUR0DudyXggQV3rTYHBGMOWzinM
vewHea5C+HjDmr+1nyITeqiVZ2xjZHVb7PH0weQTzmUrdkXDap0YpBfxnrWbk72o
ntUmq8E+HjOWC8f2OR9czIPpm1ubZd+fVFR0mnmcVf0IwLjtANEAr7TojuFvco2k
YDmSvRfg+o7nfxw8Rs0P/2QprAMK2CiZLgqvoFKkOWju127v5tR4AAw8pmvJsjmy
6IqxgTUPXt3aWawbqn/Z3KecAKv3pzUrTCzBx8FXuSvCQn8n5ejOmqmqBimhUmYg
t9lD7+aKSJL0XSe270XdVYqvizxNsElOehAQWcl6wbgBI53Y5Yn80bLZHAGJPams
weYof8sTnYSd7/JWx8HikPFuiLq/XztPt4HTbmpJG5R5+pjaFRQuYyrrSp6j2Ouc
5eLpZJcWcFnh4Qv/F+LX9DdtfkzDOFfqDzp391eYN/wLiwjDFcTJ02dPUjcg8bJK
XeTE2sDgUgNCQ7U2iWsLFniccxL8zew/ywIjUtNKU3109wClydJBmrKSljyUp5+Q
fy8nn4Fb/jxgfb2cTfCcyA9mmFw2m0nTFt3AQUfFx6CyYw4/S26dxrNYdQq39pkD
miUclkR8UbJDcO9FgJtFo7NvpLgf8/s26ssHwDJEvK/QTbtpQ+pAzFbUltfoq0j3
QwuJkk3OKItvWEcxpdgm0pSGbxlT2SDSZEAFtuZmXUvq0qcBfZGa/e74iZH5XlF9
TbZb2JHXxcxYensKHtCNCywJfWfahHf+yod+kgdqbRRhnKGoqdEgbbvNq7Z3D01z
SVFBGMJlM59qeIlroaMzYhKqFJajEIL1RW5ynOuZr1opg3ZWAweVjQ6LIC50D3Iw
jTngJU5x/cChiyAtvpmDo8Z1A/W6VmslRReic/YRpNr2CtDyFp3X1LdeXA4w82LK
rKWde59jXg1rXeknX+fTxBihPf1n8Ibqgd5V+jO87zJWwfgZ6IrOhXnMXnMz61X6
k/3V+6To12TfR2EYyopDa5HSX9ZHhIVeMRsItAL69YrDSb27pDBSATpxON3Cgblp
DTaREmPZI8d/v4LRuznUZoIH+TtrFhxwZObtw9rll0t/07+Qv4EqZBFXTrr01UU9
nZe1bm62mt20elQ510HoT78S+fiAMcsYrfCsTO3X7wDyxBBSGTOH1BauLIFgHv8N
nt3XGjLRdlfGNoeJM76nnxu1yOv56kiqS3pWpWMsmefHYWuAKcPnrNJwkGmLo/8y
lnb2jGLwprojftbfxa61GgBTveD//WxPwGWA/Xq4dV6fsqueSZw/LeMW/CS7mqfQ
FgddcuewaYP//29edLAbu70usga0okg3S8vjiQbsuPxD1YtPzqzQFJvoE5Kot7aP
SYYH5qmtvsShtNPpuv5dq2frBplHPsEwZ64JsiYA/puzSok2BZIvzUDFuYcvFX8P
Py89/PXIA7nkgqvdp02a/tXwrnzBF1QcW6s+8cmZ0cf/tAu9GiF74NQt25MCHnrQ
eAgmspMNxbjgccBZA1IOHfvj1tutEtKz2l+hDoFGSIU+6A6slsGM1W2Q0eKLOuoD
8ZvCcEHrpJ711UNRBp9Do4cEqwl/GHabj0SSidHzOzFauLvojFj9zcyUVDZ4CCcP
kdwICQF8g8p2BcUT79W9OwjOlxui545jH+qMQlYk5DlygamkIDzm/3G5NuHoyCEp
NnV2sT3KgL4IBpuLc16IQZPTNJbeJsnZTg+l9m1wnrY0A2gW1QkT5UyzW6k5U9oq
oCoYjSf85zP0tUY2HXq6Hx/Hs45FgdtCDJdCk0x/WMGIc3NVqQUSYs26uG7HVURJ
z3VT7W7OO+WmUbejK/aubcM5ltbfL3pb5GU2V1YFF/VZIiabH9+02iw8z+8h4XJQ
FWl/4L/Qp7e7WZWUe0C/LBXRi6Y/tRKoZBgZ1K8DH+kgqgXmWSwNV6wwcFUQH/pC
Yi4ZCkWNzVU0AzdF/X8zT7EB2Fo05elRpczzBHPUCxJLq6SVVe4LiGy8cp3uGy3t
WQN7pMVtaWEWLz4iMi92eV3bouL6vBeOxi719qRZAQ2PEapCZ49w3/+NBRRdPstC
KihA4/GQmlFWsPmMzVNzby+5oJiDIKIU5KJJAwOpPrqcjL408redxbR7xuHKpFtE
6IV/v/DhHHRZIAOvcMWcbnXhQvfVOZiLNRUkGCyy9uZQmej8tFZyAb+NmJ31EnsU
KZ9BsVu1o86qEpMHnbJNeqBSzQ+TTcH41j3FqIhbORT/dpMXXHbjcU9eWoeX3Wax
jegd0/3weD3421XTRfJiJ7ijaDedD4b+FRLwrIgCQum8C07eKwY1bKgh8POS9K+o
WcECXWROUWawbp1i+QaXnZ5CbHYcknS9FWNJDcOhesBiqP05PINnVxZ2ndFbdY+y
mTqvuGSswCzGrRE/LpsZAHBABrqVoy+QeQ+ZkxUyp7BQkiffg3GSdsSGyE9+AuHp
m8QsXTcZRV6mSaCT1esJaez/zGQ1yRAO6VZwK8hg317YerM0slLUpPIKkB1EhpNA
lr5Odgxr6GNdueIe3Uw4JrihD+hBfyAWEA7wXJ842nSjP1OYnHO+mt/Hu+28lnwn
j5NX0AuEN6CdZ+hLbnInR0/18GzG3jKFAnXh5nPoqB7d88XMIA7RwD80sX0VAqmZ
/3UchKxxpIjL4uJhzZ603R1d8Wl/Y1R16NtZD3PQJl/z+h7VF2iD+IwB3I4FbCwq
riX1a9XSRkQT8w7LcHkWQOkCOw6iMI9hhMIP8PidcnJhY+2gaM0TC6WD7RxsDn2P
l+lltFvv3thSmY3oROttiQAc0pBQ9r7hpvQi0k7sDU/VwFBauFSkciWe9WnrwR5+
DZbNFIetEgau+t60F8sDyYWO3/IVSa/8Hv4MuKGYcD0mucx1Px3UPWHRs4rmsF+X
wQpZVgAbmvsWTRtSieC2e+7W6fSMgDO21aw3nBrsUMBugu3bXq+X/fTV0yFIH0xp
w5z68ZarVGkjQd9P8L9xYEb+mbTIoGu/HVKqHE1kl9oM75GM88dcO4pPRaW6A3Pf
scw98cnXBS3SmXpBVfi8fs4PxRR9yBieHvXzOWnqX96yZaAVvnted3V4Lva40OvY
ySap3r37lJc11ilP6L0Iv1/P2O8mCU0PU/XE68XnQbLArz8mYvh2q+0gn7W0Haat
nlaISMseGShgLnYlnvwSXwF0fFqSpPEvpuRsxjef+WkO1GMbPx7rGFcyo8Ic/C0m
SueJ++X9Z+VnOTdnUq1DXglWhHwVtn9JvNWpJnUvjluPT3xHgDZApxwW9UT8dpqq
LKU7yK489HW2DF1QW+k8nrtjYSjBrHJHP0d0TcZ1xNgEtnoRPGyFg1HsAA9IBX5c
c1QkIZ9sy0sjcd2fQwhK75jiNahPwNKD18WmSarMsgkfF2F/7ld8CfHAsgUaeCYI
qKn8uT2dfI1hIU/zbtQJIeHxHbOfsUgR/Ywpds0xcar5fOw5MaWI5Wc6yDY4MvJl
Fyz2BRMUQ/4vCqavEurTZQglp6dm6MJHsodFqkkRMQoxxmY+0JcEsZWoULQc9H89
e0mn+ATMtYV8uzChroi+vKfZCNfpkLR1+Crqf3V7t2tmQcbAhKG1Y/LVZucSKOK/
fj4MJMizrm+im+sBqj4kuMLb5l/+tPy8XV8jT/k/F35XlwJXqBNBmU0GOCDZ24h3
lypCVf8TK5KRAmw2mo4Ukmaab3U1lDKrmGBAyLukwhmg+BV1XDDHlMnWiLf5y0HR
56Pyi3786BrakYsnLh6bOR1rlZP8jwWG+0yTF3VBYt2xrE/CudGW+hIgQhdANuOR
6TdjggN3m1EVz0DRN86EEVmETwPBiUy4i2R2ePJ3LuNB8T1nLTHOVipUZMZlh3wC
ct70+/5D8jmt1GsYB5maZhhvOBH+XoKkdO7S1+V0hdntf7+pD7LzEhyuvyzMRT37
XGYoO4li4B7VssBbKEXaEpVkmv4oaQJIkNCuSxcADWFd9Bm9wBtHuo5Z8yAsZgGs
4KaSRCmOZ6daXGBWFW8PQ6gTfbicL8KdbX3PvBQiaBh2i/oL2KbK/EXsFq6QUbad
Bk/O42IXXxQMlHMUjINLcmq42AwS93Cz8SDbfktL7Vdx8Co4ks1GwtcI4UuIReIW
zlifCIt7+yoV6HgkxPBnKX9hPrLIJominc9hzt0gaXbdcCHcec+EMvIx0CfEAvtE
iE4/XtphCj+wppbdNxjny4fNUti/HFAiLnMAl/hJqjlYZh0cd6VJNt9dD3J7i+q9
cpZM5L7egMTPC2xkZ4NVHw0dizoIjh8izWVkhA0ovADmQsLXeAVzd0rwus2g09pi
3dToNBYJZUBIcp7LJf1ipytDBRYDe+7+CHbvczjWRYGMRNEIxJnZJfa5QhugnVMa
5fbLmRzf7LpjnNs3OsFRV3LTKEItyuz3TgA6lH3v/u69GT4NqknrxwRDZo+Q9+cD
MoeUeJc5zMByWkQ9tA7Wk0BMqGTnNK8Nbh+AwKx54OXtjTEoRAjbiEB09QjJ61N4
kEB89Tuqm9/lJsoaLDgJDT9lRg8ih2N3rWlJrJkzf9D9ZKuHHchSqh+T5YTTSoJ1
QcaUvbQmKMRG8LOq4YJCDsYXnSqyQdsy/SApzFcMjS0HYEUtcfoz4GeEOx2ih7gG
s+We413uDdtYzijjvO8vSg2imYTccWvRG1hVaizLeaF77DDMp5a9tGzfcen4PmUn
i5MmHBr0297PBUKlNolkY/rU5svEmJfwqHo6VV+iQoGNiXIJ3XF5wZ6GlmIiEyTW
0HHJxTBlewNhbrQeT4kPeoi+Ttr/H046u7LDtgWI6xF+jtB9UFV7BWVvJNkx8D6V
K5rjsCWbFHewvOC9D1HkJbyGZons0rz7KXE8GMqRNgJxailS3z4RNt0DZCypxNgi
aYr7LVq2t3slywjNEzt0zt+TJtNY1QMbtQ7JBQr3bR12qgK35QMWp5a1V5Md7xO5
gKFnEPIN/shXM17k+V7O6zuxXNNK5jMYXD/GqiIHmaFnFp+u5yi0nrCJc3mtB/K3
DMfrtJkWcJSiLQMI7/ExUbStHn95aY3u40u3dEWL3FMAzxvaTJ65r3vUF+1sCI2y
RWNMvwVunh+r6u+mKg9zsd23slHcgV8ZqqWa4wPU8OI0u+D2T/eKXbi6LQ3HyDOq
I03Qz3sS6t3YV6VIjbcWJOujIx/rPBT+kDZpoiXJDbIlBOQkKJvvO38pGMCFIXOY
TJLdCabuNkma1CT2Acadn0RQyw1xhPYzRhj/XXZaJtdYwKV1DnPvXEXO6EV7Oaid
QCRJoJlIb2JNnRXYtpL+4lp84QMukMsyyH1ifGpYtfA+eUWecEONiSsdJUgXSu6j
HWzmbYK9QUWQYnPKolqAFKvzqCJdwl69QXm1lNnDBsHN5Zo3S2ThVy4QenZRm9IZ
sVnfXr8c1nlUb/rTob3b9e6M1QTeKBwQIb83xovfWIpGGCzVJ+qUQvGMyTYBInWo
CRQPafhSE+AwzkpXdYdCqArROdWOcfFQYs8vpktQ+XnE9DpUjDP9bSJg5Vs/q5wc
4YPBIUVvbLEvn5VzaoNL5A9c/0QQktA/lVd51o/k5jsWnmFM9K9TYBko416L8ygm
HhbP3Te/tSZBg5fKKyKHe2c2oeN+rvfy1Mp7PDyOhtX3wTNrhLvIkD6D9wH6tWxc
0ZKpuY1TfnemD3iHygnu+lue1tz5rmRifMA7n5gcl+leHGg2n8AgMPbMdLyKDTlm
6NVuPfQ6vCJIduqlwlJIDjjobSu5FEAsuinRkVAgH489SJ8DBLrUGRuFqwWwaxpA
n0XAXfgFbmrSY0duurx3R7Ltv0WifWiJTpfAo8GKNJIsdy23zPDTq6iGS2PnNhnZ
wsD0x4bCr9EjN5wfp2T6vyOrO6++l28O0kYRm6LazQ4rApuMKPCV0uYhcj0dAnkY
p0+qed7E42plTCmZrQIymdFk6KKTaRL8QF7dZrzHLL1h7ngF+epZclUByKU6BpsN
vSgAApcfOWiFh38ciL9qxV2MNyRTAtI3T37BTtzpSr0UljfDEYe2WYCw2Y7jIkSr
2/jQUFz8FYDnV7ZdYhHLQy6GmGrkcpnIJob0X3iX1NU0ikES7J8wzzrmsTeTAPjj
+e9LyyoaIUI5rn5fKcF2z1hB87Zf8lPH6GNYc6PTcLE3L0lIWw4/O0ePahlOV+zh
JlxSYLBRiUiyU9KMCy8YWpAavBBpy7td9Dbx/vDbCIV5H9fUxGeVQ/dmFeQ3YnJn
1Nz75pBPlmzq1AaWqRNxPCfbl0rqKnd2nNbR6Hs3bGgHExXkEfcHuAtqd9Y4n8/Y
rj6hKqif/Hsc28MS+Q8ivVxf6toDPF/s+iLrsw76MpMdj0G+D38enLiJK4cEFe2I
5JcxG2NlzcfyXAGkQumBtzRZs7u6nQXVe+Dztg/s4CNMXt0lVHT4EOuIdxDvMxge
wUUQL1n2waqQZ4bkQVUdvUGOu8UVo5bsnmtsw9yiJKKKksrtB6U3yZ1fNNRB3zdb
MO5rhLv+DMNBFL9rHtlJcdRt0vKKU7S47MNSYpcP0BK4WMhQeSUlF/NnXpe03An4
G11d1IIpL9K/MiJS4+jXkbYXkPgcxZWBNQhUqYgzTDmn6HnYoNK5bSKWyMFrb4X1
XK9oY8Zp/Tu0lNhGiNkWHicFjM9o1fn0yEW9obuvOkHcQTc+Gz8jt/UfoI2JvyMD
XnvM3FhXLfKH5BYrl+FRXD0Nv4A9d7e+WNF00U6aN9pmVW2Pt6vxNyarPrl9miKk
N6k4ET+cdbunzZXJostfluwWYAUIRVcn0lXnjKCbZLpITDK4/0T0D3UTMi/OEG99
t7u6UOT/FVePGW+f7Pug4n0IsTOqvfCpx/J9HOBMZ4BmTnczUsHT0FDeFVkHN21r
seDvjZ+VXWUbNJFQljjgU9tvGxj63/xibEN5cPdIrykWrjkMTO8pmSAbU3yZDQqx
j7Xmu7IMZ6CK16YYAoFS25iEsCyRp4vz9mjVqvzr+rtTD1+/S6fy+JTrC//d6hMm
oDPc3IGmsjdGJw8u52EhHXBkOWsuSplX1IVrOCurdTKeTjUpzm/lR8uHxOTMR07P
uXIpDrVTpgVU5a4GHml8Fwl+GgIDlIl2RJlYSKpMLzE=
`protect END_PROTECTED
