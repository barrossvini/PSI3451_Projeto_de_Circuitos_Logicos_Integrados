`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+6EkDgBcUnEbODNjYsm8Ib5tG6cZ3+VHV2O3FAtsaPon1u2ghnIs/CoWF9xSh53
Yb3+gZ5AqU2VJnesWQ0G7n1TFjE8iG8+90P4I8bc4B5FFli/rOOUzRkyFxP5r/oT
rJtgogmJI34Gv/DkP9MxAIJbPKx9lVUp3+MUK+XpPXbfK34zwh9B067GDJY0cWBL
seYbAia3nY6idLfM5Sa6YqxrNlaWVT6H4YdgdFL6mSuDhgwZArU1MBJ0oL0uoL7P
+egDU0GkLRud0oAX3VKdXe56Pjf6PfnFcydJpwTB8hp0LjbzzkVqZ7nU0/GYjuJZ
NIhfTtBdahfsctzkq18aT2ZhOOWQ6hf+6l9iHf6fPv3bP+PJd9WU3cdawfV5xNGN
ZHBIMLgODgcGoxLzF3rwrfUpjm+cDbuE4cHRUpk909wbm8S/AYj7Mli/wBVlKcXM
hhJ9+g8Z3aCtJvGVy9KgBBecC/oaA89FEY0H18BVrAjJTt26F5c/+bItQLsYxLjw
gwFOqnBF88z6I5QkEqP5FBCusiPpX4lMglv+G7661XFrXJbhV9aUjgVoQIMHarrB
BnCTG90CmBZIKlgtU67gEGd4MOp05+zcAe3WvbuG4yn1Y688Rq0j9THh5ikghMUT
6bbufCL9JkpjiCPOyC2ivxcpyWv0wNRgAuwK+pXsOS6rp4tM9iyvUYVNQ7NZHd8F
2Wpg8b+Ontqw++HOrugr2pQyz1MJzGzMWnSVIppf4PdIbGuV9SLe/ss2iIHUzu1e
rKX9KBl49ZB9qKfLaaV4oL+zJk6z6eXrlQvTg4W0On26moQ+rJIMBJnoeA18uchd
zrOwPqAaZxw4q46j8Ux2jPLXWhCRV2qUrrM0Hs6f2bs0TBtszi46e1hkP/od+Z2x
qefo98PIVMA1ZtoW3azmCSPlrifCrLmrzjlD6OZunrSH3HNpCDVpRcWGmiHb5miq
Fd243zcJGakWbANR0vnozYMoogL6SmabXNL76ab1c1k+VNW4eD8QrDsGhQmw9CPC
/EsA787BHQMw8NTCTG0nHdF1+ixLc/XRM4bdXrOpHCLH7dJaWVOp87ai7Q+Q57FE
PFRjz1GKYMRRrNWjf9zZ17Tn38ADdbB31lZpBvWBV1N/dhCTmaD6QF2NvWNcwSlI
ymkEAS19JC6NE4Ekx+S0vaVC2Jm+SvqMw9DKnS+i2jMDhMQahmsc0FjjafUVkNTx
ONp+77sOZj/ANEpO5qVeiz8y9nwDdwjGvtQflnjICt/LGj3Fcs9XkUxoA4Juakxw
GK+XxTMlva7FNZS/fysBZ4Gy9oYIYwuEPdk0VLBAMnRL4HY9nrTh3GfJ94/A+M05
FstJWeve61udxUwVV75vF5ubr7akJesyt9b4Nz+dD4EZGUzD5zV2SpizPgrzwcev
iDyHk4wXREO1zv6S8HtYXM6j4/XLDFUAQ04hEN0ISFm91b5ll3TjZffZBYpXFa7V
+ETswiKvwuP1IhqHgyeX3ewGivcQGg0SPK1jKnKIpv89WO93KXX6cMXplH3bxPZs
OpQrhCzZCzW6S1GUAyz1t9HgC6LgUn7vp6kchOG0LJzCpZ7isk7wGZDO1iBqIgng
lylH//AiSfAPl9WwP6iPrnmiZ3QN3PDpfwS42ygCZuahPjHbCvR+sRf3Ggrsk/RF
u8Y5EJdjBZrwYr0GH5OufyjyHkvZs0PNEaKo+sTubV2gvLoXHpkVKfGNS2DwdPMq
TcKXK/+R6ci7fv81+ny3DJcJCrV5O3BjMV5yDzrRqaVr3KsZZTs1FPbu3IKJ76JD
I4YhxZAvHE1i3BqBU3NAS2jbV9pSHY9b1rCFp179I0grV4g8jgOqAfL63ZlRHKzW
iNevgW/C1jQN/XM21xsv/OXZX3LOmrgKCoux8Ujnwokr4hANYNBOd28ulP2mLKqC
kY1TuzofRALAuHv3fFntRfcHMrXaMIVtqJ/83WGiEmg/E9FLuOc5+opLbps3zMxA
VDRl3s1epWndT01fRWouLKJB2Bg2qgPUytuYvk6chxybJxtoUSa/bbMknOyg9C2N
+UPb5MAztoZLeonznmTWMdQmgKaIyyKOOlpr+m2xZSJHKBv5xyQ6M4IhQZViIc1Q
BTO6OcxPXGJcIvlZd4j/D0n4cy2g6wmjS/9EO8JgT9dOrEjbP2cyh/rKg8OrL5VN
3z34/6K7+x2S5swcbqJ8m702xdPF1loGU/205CfXfmPEJHbq6NakV0SZHIC1RMvB
M7bkqqCIbd7UGbYyPc+yeOhwnYslM25vW/eR6u9gOLqUyq34SZp961RcgFD3aEQl
XB7gqwwQJPYnai6YJdeYgXpz/cwScT5TgUq3p8qe2xnl3YcNqeUNd+KipN+zUGDJ
AOABAURZarTeqt++mcrCWF0R6q+20vyLCJqLbxbx+ZuoxpGpzk/SpjFxq10fYmG7
6Olfmsz0/fnjFLMlZQU77241lbgK0iFrXgeB+/qdMJDqIgz5bpjF38+UL4ENlpei
ufHbT4iOoON92Mc69q4vmTSZ8Mc9N+q6t+LxOt0VlpJeotvp+ZMcgcmmO+jX6rda
BCyi0ixJNqF7LkGqvMbWpLpKoAAmYc/oi3FBoEnZeUdpGhhpD0NkLJPv7IYfhB2a
28wTXVdE7SMLJBjsIp/9ulLpcuzGZG4Aiw1MN1PPZrAbqLfcZ2KWQ0zEABd7rEBX
WGfjtggiNozxhL+Cj2Q2LGWAAai0loCNY3X5iRqcHwnyJCsg/K7meNb8Haij+gp1
I6qcmAYWTYvomhjrAtH5hg==
`protect END_PROTECTED
