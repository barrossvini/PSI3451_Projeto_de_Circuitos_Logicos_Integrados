`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dO+Nc5jNZzzOxBK6trVJN00iS4O+rVZ1kBCTdBj+H/DeA1b8wZCuXj7UDkDguYOf
AHHLkCUp/WxppWiNXNfk4PUeNG7/eGAwCP+9jSVjk1/c33lH7Cp4SI1Z46I/ehzT
OSR0GlJAE5n+N/OgU0bPIkqnOzrPM3+DZKHvhXjke/8/vExqegnXtE6/V8yGef/+
0iWS9hK94mfh4kzenpWIKMjHSAtGMqzzemTurJDnyzEoHvHjF3ft58wB2TzBIVfe
94/49JXaSflq9HSm3Ddk/LmRlgasTU3ecaimZo050b3q5GgAZ2fg10O6mGiFgxai
o+O0kRMcROrh2t8x1sbubV7LzgM1OefmcuLwnN45xPZBSjV4AxEFyyxmdx1wkH4m
wbngDSM4lSFJ9bmb8Fjqmf9U4+kmE9oBh5VM52WrfRZC+dHAuw7sowfRaUfUpmOg
zq3DgPu7n7DFn/+IOy7BvTHPxWMdd5xbIbtboBSHN66cGB7Z1+Dskm2yHLlVAptf
hIAMeY/YIJi5UcLrYH1+iYmnEznE+NKnky1qMj1qUotB/H/Kke3eljtJSDEkusDc
QXt5F/KohW4G9n9b62CyDQMUSsGpFb5z+gwde1Bh8TDj1xEXVNU26I4zVhiL+qFJ
bkgxIjYDB8FjHMqulVY86ITWt6xk9MWNcLAtjMqNsi/OOvZx04z3JVqo/Py10mm6
C7AJHpshFp6YgwZkZ5BxPtfqMQNx/MrVgEkxKon1KvfPA4tC9huKVYFgUQUlHmWI
L/fFk8XapB5rr8584n660+qdGndHGUHUFETMswhWzahRdETgHgcVmdA8LN6JWyUK
IjWbc5AAKH85iTkVcYCAJX3/m/YhK7WaG31mcKwDyRGuVw6eIfQdLrXL2utea47s
QuIgNEKdl93Xn1T/4DrhnG4r+8/UvyFKF9XBpUb6EjJUL8/lSPbVV4N7qZF6dIYJ
wNKe/A+egjZzakKMRz0szdUF/phwbpgNxXImoJQe6IA4/Iz4Er8xOULp2otbkMZp
Okr1k115A2zpPTsgxMB8sQ8hAIf48kEgRS6FTcG4mmJgViPPCg9SccuVoTnxUaVz
rDUcSIIniXPCZIuKNuZ3xA==
`protect END_PROTECTED
