`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j/GKHYfnekWcC5d2Vzxlsluo8gkaNQQTVvOEoVcNzYm2qKwDr6rlhY9lJTaabcdd
i64BY/jY4bKcIEcECUOQ/yZnTckNlWcrGp8pY8a9Gn+ccteycYTZFKa8V0hZF6yt
/HsJ+cKqMINx0az59YD5iIkbee1gQEQum0ee3M1EBjUdu410K14AprhVNitbsrKw
UK2ld/50lQhU0DYaSo4GHtTuHl6pacpWX4tBBYQnKcGxsjS60U0hrRa9g+L2dKgj
yhMsMx894KAwyz9i3PatPG2RIjYuHJbE6NLPhUVg8z1snNrEfTZA19U/IdQuT1UZ
YBCzRYOz1TuslYlUxed6tmgwMRS96RTEwfE2JKhEjc6ze/U11zFnsTiVI6NiDree
g0tbUfh1Wv6Cor5OaBmAvBKvK6Dp2WNLEOc6KPqT8dhfzx5iz5LKOHKgsV7RyLdB
mQR31Wf1nJd9iM82hfhu4+XZAjS2SGIo4znuvudqY1Oe1s9R6GPNl/mphdw5cQYr
bl0voGmPF8Hmv22ht7v9NoYinjqW2tA5dC2WjgkcrrepgS/vnJFg9qeL8Ck5hSYi
2tkLOhanoCVk7wRQHLOdZYD+163603kTcuBUSFnNbsJ97fmYtQa2pd/KBYTfGlRH
uYKuKrZfyJ7cSUUB/M5B5VTU2KXwRaYRQB0YoBtHOjT5PDo+RjO0psiForwLCjIk
xTsaLRl+2ai5fBJuh6Bls+bZBLK5T0YNyKqo2cUeDrpNfI6qzJCEWn7dqw1IeWxp
XMMrMZroyetXEz5gN3dzvdBWCknWzYoX5K3X3C80+zFPDeXirp91YDOJ/bZ08Lov
1ZoHzK6Q1a4+i/0cOPT3kfvROAdieb+h4SBCn9JRVwlDOgxnhDQfz0doGf/5K2YN
Vbff4JhivQBEc1JG9xav78mbGyx2J5DwAJd6G5DChiqV3vwuK9cf8irlUj3PL4ui
cKzZJ73hVz1yfLufbkpZtrEiuZHoscAjHhh5UPu/khTD8UKRYTs478i2d1w8HWce
3bSPtYyRbHoSXpmcxbZlghr+pm5xLC2bH/n92Qn2losC7rMyUOxQm8lGSDbKl9Qe
n14yVbM0o/WSpk6CtEc/N6pkXosGEoI//PApNv3nNK9p5TTAqdwbYnypJEowq9pR
xPXfQMOCfXD4SIyf8/A4WGbRU1XbQbgseO9sjh4ZbHU2QqfjL2ILFFg/RRNEM8MW
whm0zSmk1oCFhhxF1sfWqpDSaQWqagRMuNrTptwjnWa1qQetEuR42oBFQt2+rZNF
cNRHap1TuZOrQAIp8NBPnf6EhtWIHnsy+QWrZJWiWEEKYkGgD+V3LlzslmHrJxeW
+5Ec8wZ90iIBIEDDhUc3Ie8Ig/tthCKUhORigZHiacJGUGP1vkFHefnKY3jMSas/
PupztBtHRYUQXKEi0qBxYjzLUlYWuJVg19vShK+PpbY5WBZFQNBiL60d6Apjexm+
wlj45VGD9k6JMeCgVoWXUzZMGt/M1hBiRAvF8ZdSIMiCww2PhqfYT5tgMyafT09T
KG5A2jq7HxmmzKKUsh6kx430r7+het61EjU1Lz8XsFC7/83Ot1KiyS5k3ZqlauDE
GMVXMi9ykUUTay/bU42GoLgfOVAFDxyoFtChuGXDJ0jpexuDiILloimMFI9XYzKr
cMXxVpzuu7ER+S5Ft7hWtSxEEAsW4tVgqp5bAJC1qXLeEjvv4oREg3N8w/07RlOj
JY9kjOy/inzV0EnDWAHFgkXmvDprgrLwWzaEiYOQdnILBpiK8h8Ik8jrfQ4h4CKC
LcKfaEZEieUpp6laIxfWT6q6VND/EH7aTkGagn/ppjaRCG90Lth3uxdfj2CkwkIJ
+eZYKbKNWzsF3IbW85v/8NbYz4t780FkeihO2yWNiyM4pML59T7eFphmJxn2iJQm
FXvQfC8hGI9PoRdvCD1aojeNdIs2BCvS3wRCCu0cScYv19vsDl0M1JBVWCJNpDzw
hF2r/+l3QqMXHJHhnUkI+nDYgB7aEsV7rPCH3EDRpct5aYiFIuar7xu67k6ztf5Q
67nRJZk/Lx9mAxv0dD5Mxn0yADUSpRktsM2efVG7v0mqI/St4atEipvAHl7trTGd
XRFF0UCESsoqSz9ATNLvSBEilDbDjFCQX80LCWVc/QM0R4iT6zWuuPqzcbEajwvT
cPlNj1uJ36Fb5BFIIdnKe1/2mJ1LVDGLpuFXheX7+Lu9d1Nx8xoufcf+0onXTMOY
Vsy/Hf6eJpY4A13jME4sFKRDGVqUdKGiI0NshpuVpuuke0mrZS4UVqGXlG9+vIIK
bNUPb8gS9RHQxdM974vA+gfEfmuJqsOwGQsWlRALrq74JuEN+R2MEprcjAkZEqK4
hztlD887w9fJjSqxKYFfRoSdZgHuuVCs1NmPIUjeemLK5Cgn6r6PJwWVvn2/96e+
Xys168O615EvWLXN6qSb/8ypslBqFMUhPmatepCa4VEqTd/Am6PQLGZvix/7cKiM
tK7fSx16K77xShdD7OzD7xY6SrO0r5DRrKr/iNkPvh6G0eKp645BCZytaOjgB79r
LCzBn1eFgAX93FiEJLREnsnuRkLX28Va+t9F35pMDvW6S5XJRUOyLd74FfN3KejR
USQfFNmBzJRLIYb76qB0HFU5JAca2L9gFCgDiQs8i6tSfus4O+KhKGqH78rFU7US
KbEqVMwsy9QrcW6Q5VSyus/MA7ea+219CkxTyE5qfurMDArmWSioak8pvMoVuIUI
WAXsSDN19sE3iwQulFJsM537ryCga7XnrNv0k08GhY57AUoAYmkHvZYp79kqRqvr
GwbR9SOu7I1I00kJVVdPaQR8wv8lJO9XxuT53gOAxs4sSalRWMcdDpLM+SQTHxto
cL132kaaRQx15pbufequKXOl+JwqtopaIAlWvAU0nmzAdRdC5LAfvGD4L/t6+Y5C
+dWK00pJRlXx32T+VNYUuvi67A6FzNDiZ5bT4oewj9TFTFlL93QhfTfQYe4FKvq6
VTWtP/4KhWMQkjE6SwAFB1TNuS6xLRbxgGZve2jl4ibJA7ko546f1juC5YVjJ1K5
LDLArB+17ofwRecjchp2i2RU8VZmDXykQ3LFhBaJrYEG7BNeAdzE/uycOAq4fw2y
PTMkaFM8ZlIx7q22kzfAkQU4ScUPXMYbdQEPwyKL0kLDeJwVsjttlE1wQYWPqSoS
ep0RWOCfrFJ3omullOwBHvImNSM0/9SN2wY68V+L9Ld2/X+/aFEzWaqGe7Fmww0S
vjwZE/ZoUDMs+/YSNlqXiUuAtGPJm4lrx9GqFLUGQTFwpbyenXQ66fR3wFNGQum4
JlxPDIzxiQtBNjevXdEU0MTNzBbBR+L+9FnGANn0BtNInsI87cetenVTIXODTWrp
6h0uGgNfPVAOpzhRxaNlTbjyiZh95nwkgOjVoUar9oYOA+rygcsENiT4njRD7qgz
29m1/EbY4O/RMxlA2/U1SJCY+3UvcbcF5mLGNKhEbTeA8q2tnmH8ceoISVsP9Xar
YFJkjEJAM37FOYz9aDd3J/iE1aNb0LWlVIQ6UZSZPuZNb6sqLtVChqO9+5/9YeNB
5oEZ0qPbKPb7dyJSFnKY9L0rQsaDb6lTneEU+03rJ8RG1IOiVIaatnbHxzPLuUuY
D0NNKtz1EZV7BCoa8lwIs6XMyHFVvvtD5kiVCl83LY0NgEYuN+O2jvaCmkKYNPT/
sMSDTatwktm66YEilAwjK7fDqADANYk0mDrctfcWEC/zW6JdtpXlddZRdskEo/+Z
qrYUdjLnQy3ID+vg5PdLf0SKFCo2OO6GALDr5hP7k4WCC8OrE3pz/ibSkZXzwmjB
uv4T8rvmxuauz+Uje62RyukGLNhPKo6X+gZ1rn6PQ0joPVJPqjmiqwCUEzMMeTLD
BBopzNuLAcIgk0/TtAm6IhnRgSmYb4bFbOnzLq5/tzMFU+a1vUhQtFvAtDcT25dm
eMMfY1+gUqIdUQZOEPS/vNFdlhTm94t7cUS4PnLC1khxIL88wEiMRrM7txCWI29T
JQ/h21ixh78gMZbGU/TXBzjTC5Iedbwku3KPErhgwiVbdRx/lVGK980RTMnxSgoG
Pp7XoA7bCAt6q+p0Vbdu2tbJWdf7Qiw2RwjahwLB5EYd/GMO2Qfs8uouxEpCDFY0
LRmHFtFP6+CoE7dFxpDKd5ByvvAczE/aDfHRYKlT1v7OqTVkkPfOe/n0gArwegTF
Ud2S77xzpdmec6k7CSOscj7dIUMS1/YJfHwTOgcRQETice5e6J1637htCyNBkSmh
V6htGwPA+Uq9CkHCB+leL29wnbaPPprP/ZFR6n4WvLWtms3zpBnR7WiFnKY5pHjC
/qBTcN3EFS7KGkxMD9ARD1GL0DgvhntsTvY7BxXAaUjwT7OfpB1NvJKVP/eR/dE8
eCiH4ZEbIzMPTFXHONMV+14ic3tMBY50tWCoQ6wGjOzAPcOW9T+4jSRs6XrZxQW/
z36zfroBs6FShWlLIbIDfmIM3p3/zclfC7DUNs1fEF6WsftEvpfNtZXK+Y3vSvVk
5Y0Qm1nIcwBigtPfqW9Cd9+AqJXpONpmG8BIwUdg0jbE5XkcUPcu9om88JY8NVrs
fPFdzSG6I4TXF4tiTWnRG2pV9emqrhqqER3lI1f0YiYHWPZAud255ecnlf85OECc
Xy3v1HvY2uU3y2r4b0a+I5vX4jt9my878mn2vhWEN0s+EIN618DwacrDuCS/ryeF
Bm5hqJFMu0IFGgDz3dmdQSOurYWCFdG8z8rb/Gxqy6CvIA0hOyFt5LVZI2LdOYDe
ko9vexkylx0lSg0BM++/ExC9HBOZKB3f65bg9kSC79u+mu/6VJaZ5Crbsc4ifpjf
dgIj/lYNDOvFhx5Mu+QfI10EarbrRJjvCNxRSgpb4mWre1P0t5zNxY3dxgWaNMWn
C/iCiyl3daJ0gk9JWaUZr0+rSR2luvO1O2mHQOwTAFrFK7UzJU9s4TdJOtfxMMYK
nnIaMMOEn7V0CFAqu7qAMRS4WuEoktyO9QTnAMgsWxakmkL+BZjCSuNiQtCQbnCR
l2yHecAKvps+YEqV1Uf2FSWGYRfTAPmMCgMEO+MxX+3Edmcti15JErHCTMMpilFh
2uOgWLY4YFpe5WeCxTGN49vBP8Er52+p/v2LM2nCtyIX3TAdDI4XhhubZiuSmIty
W8SV4uW7qu3mAkg1FdL1h3ia88RLzElfInUEDW5cpsmSJykRnXoCCSj58RnEK7/p
xPgLWA4DOov2ZAU+jqmre/LwY9UA3nCwmZGN9aaywqbPCNp/989yruicJ9xr90sW
j/p01al3D6kp5BYoyppLexUvBqcJqGTo/a+3chlm+ynF8ygyC/1xS4XBkZruw6c6
bAxZPIPNpGE2kfboV5FpJmcqwkmqXZFl0k3kHlq2zvvOQYD9J4TsnFsxeE+aKKeH
YE6bMJafRP/eOZUWShvzld4wVk/cIUeSL55exDenlkBofpLBeOTRPHaaGeGXUUfY
3V0yEu3LEKhQ09Xu63SA+3cP+M4EWPWfT3DUHxbvbOpFeMEbz9/bhCUylwbxIpv4
OA0BSqkihkCybDrWaSNm5ghZ6F6ORbiEW3BqUk6UjuUE088YGJz4V/x4KhrSXC6L
ksG5pxR+jtV04gABMUCJN+jJpdDZBk+5k9lBUBC/FebUaoqWTfqTvZxAfaGXy59N
MSnMzHT9yYhuHw9mgjUKj9zZUQIPR1KqKrmc+bU/hcpJyGVM1QLpMD7FN1w6zxwm
kYj/HFb8eDwk8wTzi/69zzh7nyJau/UVz9ZQ566BjE76fjP5dBirQRdloa1lz80q
dnQDbf9z3VEjT1d6+ytHOtzuzOkPI2wxNZ1oo2GotmQ=
`protect END_PROTECTED
