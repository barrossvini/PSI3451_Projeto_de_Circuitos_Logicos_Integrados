`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CaJEmICcDFRun5S4K3jqE16eRAdbjV2B/5FH/zvIJD6dj6pE05LgSjDO7nYgNrYP
MN6wY/JCmD1PYZWaG5bD678elpWJXXhXBMTg1dMDQQlGs/QtSuMBPYLaOjFbXgqF
1TDTLnQx0/khvXxDiF4DTiVzwxVNy4FF4LV1ay1TW90NwiRgxbDvxNVgjmQdz52D
qATby/yJDr4W+vaUQ4tkLYay7jSkHkWeLX49r60lCqwJAVFX+HPvN6iP+pz4cesw
cuIVcqLNUwWdvi0V4AprvihvU2e1AL5meqTnFEA4pX8Ytb1O2DIptxycrVnnKJm7
SGEw/rHGgdDBHQIhILTcENHh3Fjty19AE9ta0tUi9UL3+7kjZK3CDb+ogujGK3Ks
BZBMI6lGm/RfcjaU31tE6iz1tBCKuguhrwZuqtYpWyJ+Sr5p5ymG6Nv43dFfj6JE
Mal3iZBv0pF0Ewyqxzo+stuNz01R8qCnpPMt7BqBpmHbzCgW2If5IwpRJ8zITNrK
dUDQq4KeKZMePSSSfmVI42afy/9D8wGz9DLGh6VTIjqTn+F/6E2zB0UaNtrsfX6I
TjKWsRyLLHlD8h79wQXM0I26TGGp59kNls0gw3jZZ48VO6jULgi5XoHcPutY7dpq
6aODtwc0yq+PvpvUAdY7c1xfW8D54t3ycg7a8QXJEjFkskl15i0ZFHJhXBk2hGi+
8nuUu8iCDCtLsjWXdjz+KwP84zTZatXxbXLpQmi/CxqhjwsTp66XWBEAhq7t0vI0
RIVKTXci7CSnhsVvl1r78fPWX+ISqujN5bLD9PNy9/pPiKQJUK2UFhF8Dfi00YqB
HDnO9zLxgwG79IbPq1FUGd0U+2yrBtTUtaMWCw0XWm15hB7XLA02+ChSZLM6c/zA
qyW3Cx2UqlBjCzf4JZEICqVz9jw6Y9VuH3KheAe5iTj0ddC53egpoKrIui9R6J6l
70YTbr+osAuLTFsxFIyjYWaTVOwKTwgpCJGmw9KNDaL2DttT6rfPvIFXlMi+LB6F
V1O0oyPMq6qyBVKkUZjDhSZu12kZ6cbwbnqj8u9RyxLYvKqQWqJHYHYVnNS34ijk
iTvqBQ6UPwlI0SDl7Ttt88d0uBKtfHMPeSRg3j0GvuIf0GFCHGSJUKdYT7YUVFth
KkK7kWtEYsX5pKjVMCZX8tuBi/822iskvj4xBn7zvtF03SnLlpaU+m9K7oqs4PLa
kseT1JGjUdMrUBbP19t0EbyGiq2VOy92EaXl7Gz761rXSfmrjgHbDg91zL7z0M2r
LvhYLj+t00wjFW4WYxTeX+YT7OJcOs8xtvjxi5vMtpW3M4poOhXyVNTtOlbG2EvT
D2sAiqRlG3pDZWp/GtjPvNEptQmZWRyEKUBPyq76tam1MDilNYpiLBK5VZEFM8kN
x8Q50ADzHr/7N1ojEl3rotdO45KsWPStjzX+SyBmxzJD2tO26rzxH2+Px4F5TQE6
acPqNQYZolJzIDF4XEcvi5hW1fAWibivgQ8lC2sP186ZoJ7sei8wSHS+BYgRWiCs
FLbK+H0AlZAfdDMNJyaHOQswas68i7rJxT9R9LJx53MfLNWkg2TMXq+xE8B8tBs6
exzYU+3pv0SbCECR2CH4K+ollEv6gtrjyanGnipmHilfkHmo0GOShhUxYfqKa+Vt
M21+z74maJg7IWRK7+r+9LIBodtPU392sC3HsstJD4bkNNGjHsrL5BKHkBJQaVBO
CZRCm+j7FHg6RmuMFfJaUZC+2TRxhQYuqt//flHp0cHimqngdESxqvZSliJvMGWH
60ZUHBQxB+YbqAlYp5C9Ev2Cl3g9Qph+Y+7lqj5mieAzU4Ijg/mrsrtNI2DExQe6
KTn1JX9TlNzbw7/p8jJQ3VGZibyr8uLgFAkK7f/PFXgJ8BBkYWnIUoq7yH6+Emeu
WKJQS/AsBvUneKVv0ENdupC9LzW4FteHCwW8K+64SoO7eKlolbdm85z80dRx4mkp
1NOGC77KCB7LrPwyH2eVaS9DOA2cIn/hFmGcNmT/F8T/b5GJ7t1i0dgqT7EwhDjZ
TwarHGuzVsEUuNj9govJhJihmVsGDcP9CRtRF7K34mhFvy/1w3lAHiDPv5mkoJMd
VsRL2m3iABSpjRm5J4ROa+/M+S9LOntkf22VZg5tC+ua4bY3Y0+4Wt+a3pVCmCf2
LF1y6kHHOpJuau9uYQWCsMWUPcNEiXV4/J5hzpWMZme0Z/wmxJQh7vv14zl/9GZ0
izVPRFZd6MoFnThA72Gc5sBcbSY8DB5YpP8nUMyI1JoNRtWwzD50gxKxzyW8cdux
t+R6jW0NuPHhz3f16UCsN329tf4RxqU30Oq1ey+StoFheduYoHixyVfTMS7TZn0e
NKG3OE4G1/5h78MjbDvNjhMjTiCeysPBzgIIqISKpe5soVy3Fj8etT65aLpIJ2c5
K98X78jwmalx8aQS4uyufDqgLdxNMZrMIKW2pXYZBk+4o7MHB7Wwakq/onAA+5f6
cFzB5PxATiXQ14Ww292S9bqdEA8R85cC9vUJH+Arkpvs4UCFIoPkJSK6xo+sfq2T
PymVyuMmtBkDLKiGCDYLnYuMJwvZV/Jjo7wCJem7yeI26Fl01LcqbA/Dik8Io89o
K+b/HLlwOgl5tgmhVRGjH80OgwcTFlqt2WGufkyqL9s+a8H0VIKWhTrgHFywBGL/
GVGDBDUfkQVXfmrpdrzEbB1vCKBr8aZh0NRlUWJOWOpr5e6b6q8Li6gclakzulFu
U/pesnXOL7zMnC6Wv0QxCEtGkZwfEdpliEsJueNsMvMJ1yVg+2c5sVQlmNJGy+nS
mnVgjUt9p4fg4sTT6vlwySb3IP2gXXh9ekTiqrMCI2U=
`protect END_PROTECTED
