`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NzYgMpmpPDxam2hHuFzSGgjA/AUjVMatKkjtiWqKKMtBoPVeB7aPHZutPfdV3Gnb
b4BBp0+SS90JOSjj4zyNGWn702igSIAFCMHRT8TuwpGBRLE/rwggI+kQH7Cf6xr2
TbuUkaZMyrXkyMq5ziLIcEb0btuJD8yMvvHGBZIIBbXGpC/Bzao2THZFz6ZPGxZR
OjamWNLMLWou2iTKrIUy+08UAoEso8oK0bR2fV0aKrsRbxUf7od7x97Jk6aJCuZ2
zPYXkC2ckRb0gLTrDnHqeULslEL+WXLGtBHuSPUCJm5VU5g/eJSlWR42wguASXXQ
5lqNrS9UBGKS+Xd9rQQdJw1//CNI+5fYtrt59ZN7i1v9pYi+Q8mt1sDtBwJZsnPl
SPLPwulUD0KyvQSFj8YuzeVnPK9P/JqxacznDROLCp3wIH9yhenvWgFRNxC6JaJE
gpSSHraR3TQIE/InlK0x7xoPVriqdpGYURqiuVVeNWDNDI6MewKPhlVMWfwNooXy
YYMx4e76YnfKGY+takrIkqSzWH9tKljOc0XSpF8zp7vnNMrlBz/tiwGgRLPrNflD
yhIt9emUg8cctRV10rG7BQ==
`protect END_PROTECTED
