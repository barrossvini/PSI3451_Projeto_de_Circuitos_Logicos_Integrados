`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rhjn0qJ3UWhTH47yshkN1LJjEMQEENlHPwQTaSAVLu7C9/Aeuho2whfFm70Hn+Z8
GaRNxUXv3ZRmnJOXtolQ40rixCxu5BvZSHEsMQLbrVBpduCA40z2PZatVxvLW2VD
4daqFMlVEnPbc6SD1xR9rokCgFdfHiEvxOAFcjpiin+NE7/vSYBJeLpp7NZ4X3p8
7Eiyxd4gj9sdazVdRlarACOKOlVEbY9H+3VXDlIKj8wLJGSziv1a8Ih3/oedexu8
mY4/va27OAGR7MLF4imwhd8tDZzJIEwbDRaRSA/71j3PGqs6GZJFfjrhN7S7GNN9
hqSWkruA5xl6S/uV+r9Ud9I3I0ghnvdPZ8loLOSx3N3PAqZwmga5Xo1Sk2HTEvZI
i3BTv2fJxTfo8RTHyWtBS9B+25NcS+uznLK2xu64R2unBVf0aO9qbkU1encJiom6
0XQtZAK8Oh/N+omsvKz93QAFmCcjJxJffE6zGh+n4fHC/p+5gUku2C/NZi2RZ41e
JgiQ4pHeG8Cp+ueNsp2V2r5mNadT0lQ7njhL0c4ATulfPGs3Im/rhH+udDexfEYs
0T3lCG+HzZxpao4vV+9p1fbIt1AhGe8EGG/F1tP3xHeE9VD4FUOd6/iCNVsXmOo9
JFEW3vn5ShW2ij4dPPRHw/a3DVESdQt9LWrw1F0zNb9AxoBgNJr9Z1qatrYiTQrE
jZZ41qXN1w253/I2uJru4NWobBs6mSW+gobHb8d0Xzd9lQe+Q/aB7L7fpt9/JlUx
fbKoPENgQqTN2xL2Gq02URkYaITgWDy0B6Ul3PZH/gCRZfUeh894ImGhZuYAhJt+
MXkQl8fFzIJg24qKgOXBwbCkzAG2WX8eMaqJW0op2IAZNTs8/fuQbcSa1UySMmVB
Dsh6omCRufFkk55PeD0MZHTZQ7OtdNiObXd90wifuFpooZuEhGIzfdY7NHmnMHo0
6GaHFOQpFF2qmb/peTcqWAFKSwm9204HeeBiBQmEKl1AYBzL9Nre8IOYTXJERYLV
MIUomPwLOnQ9vvIWqMa229Ynscxr+QxCyc9fmglkXPMNQ1kvkopHx99sNYr8R4i5
y/M7ea6X+pZOhUyTzY/mYfYTgDPLAWrK1qc5oTENscu1uGgc2BoeGn1KbmnBk8u3
y7hAUUg9P6fTIBV1POo774bqXYt4GGWZN6Aax0hU5zPplmA0Voa75HKR0NDZO5xP
wCvDODVsULKmTyEDUMgT8Ki+Zc+EJ3RgZhrgbtB/e8W8KnoxDJnRLtSKZL5VJde6
6/1GTZz3kj4MpKQEAKPLpdFnl9ajyyNOpEhVCjL1FkzmnictTx8nzpyMCvJh2IDD
CrEf7qqcJxpQ//hITiLKCeSk2S26BR8WjiyEQxqkgJLYCWirjjycKAvkgbu/GPiK
bsKO/OSk5V0x4JiTtQc2X8UgERTp9mylVDljkPqW3y3HdL7ltahb80zI4Zn64QNr
hs3c/o7bFKdF1bjqzKs7qxiQVmtcNc1C6IMyvlDobTE0lv9r+DLcnEJQDmMBj9sC
RHXPEH74gnM9gDIynqyUK8RtRHd2FK/rxl0PaW1imQ55K+lv0H3c0HYqvzP336bj
saOr579m1voSVDsVgS1TYDZfmHmhTljco2RaIOCJe5UwxNUnqOnvJeszxYzV0K1q
oa2Vu/CVCnmMjeIrbR1NtL/szt0YzornVptP8vVGe2aLhIR43WHEB9RHQNI3Kawn
6HEsP00F/20nk1cv3Gkeng/5yYQqJAsCH5d/haCbb8altydJ4SxTLXifUsxNsYXd
hWTw4sAttl+AOtvmGJGiNjhLCwaiD6BnUczqwyOuVFGJVDBYwHftbc9/4D8qED8v
3nKhrHpZDgFhPZDrRm0M/VyrOnls+a9fbbqTPPPy3g9stMsVs+PmllNZN00mNXG7
l75P45BGDCe7Y4sN1c/jmvCFkQSggrhSre7k52XilK5BWiWw3Klg9Z+pCcza6EQb
XBY69b+VLUu/WdBrjuVXFYXg0zuLz2H+VPRbxaTiVIBj2rI8GiGLcnUWhb2s+rAy
tvFDB1u0LtQvCm615X/g8MQB579RaNEFoqC1jgPu2AUxjiMAOzV3RHdNTSsLplCG
J2GCRmLCH+hdY6H4RABXszqm2BhCQ8sSnuMpt60q/6ihX16xONHUEFy1sXc20rDn
TGMx/Z+P7urq4QcRhJO3rXoberx5gEIOnmN6HDgbUFtda2zzRwxt6+JRhDJBrVsC
bG927mnItlXk2GdAM/3RvsyT0hVda6dTWpHo8PYE2YcQzvgWL89ClIk4nij0abjG
LOSUXl9qiMrL1n0TI/TnWGOYVKtkNyZj2Y8czmNr+DVWwRmgj4jGEG6CR2/Bh2ja
wZHzdk8J3Ky4pCLffspfbULEiK8hb2QdlpS+Pq11Foj63iJ35Q5Y2U4Esvtg8wpD
rFAfDKw9YIpQJ8bPP8L1AjZuugIpivV9YlfvShH7DUdwEih0sBI3HcxYm8+yBnyw
4E4s4iAH6/xVLqaUd7Z3OAuEI/b9NRKv0iVyuftf3CzHdQC3zHStoXplaeeQYRIv
BFotBRYEUbjfmm3VhlHWp0lCkVhvJ/8y96TgMFI24CDwv7fc2EoGZqnG5QYVSRNX
e76uvhMw+Ul+lWkGcPgUBUxJRNLpH0wXXX6x0mwe2XBqeXT1JAgY8tTnpBYR6YHf
eAFAhS5iD3NspIiPBkr1OIGKF9Jmb+1ZHde8fylPkXmLszhLLKpAzoIhMfu7DShb
Bo35szLOh5RNfDYfl+8mHPQAHzGOboyrChjOcCWltVsmWIv/IWaAulT5T1TgtjyP
z6B6AsvHILtxdtHAtciVvZRtCyYhp78eBClMwU+f3zEUqcCJ9+vrU2XgyrWGKb//
F/l+vKNlfycjVMDUJp1W8TJzpB2O+qEWm9Pvrqm7XcejW4o8j1beoCkZTD9uJi1G
dlPM1uh732NuuHS2ylWxj0eQr0A/FbJh3lseTrIthWxoAhTGi58kwGLdAZ07bexe
AJbniryYx14KAineCRwf8sFQESe5NbkbqHG97WxoxEf+9qC6K+eCYLEjRdUbE6op
9MtXEcYn3ghabqqgUxVQDc853aDfs5p6Jo+ROBIuiTTAXtZRVx4jEcui/r1NwKTZ
MW1p0OIq1i8zOfvsyQ6+4+NBhFHejxgJNOFiDh6Ojm6R2J+7f747kKealFKqLgoL
HEcHzzBbW95scSDYRkemG2d3vn63la34VmsEbDdrRs6/0O6nUPBxZW/msYwN0FKh
lNr4zjsJX9XJe9ACg9jpTnkxA0LR4UtZc3TBViuUidzt/O4gUmYISDdZMF7lNuGu
mZ2H9m8XV76ea6c8WksGMewD3AaC/v6g1LsR1PUPM5kUbq18sMAdy0KInZvn87HQ
SeVxJznQhzMNdaQgfkBnJnQPm22/buyy5RspCPZwI99Rzv+ANRR0jg9mMDs7qdri
DA5gqXVnzT0KaAp8VdEPuPTG5uuwvaOjVDjLJTc79A78TjxPgY76FNcH/KCyue7u
6Eez1sl0PjNAQY51WiG6KEpgyBiCkG7DQtE7ZXR++Fp8E8jH5IwtZtHqe+Nli9Q9
kitm/ARaHfyfOIlC4UPwbRFpzMNT71I942edWfhaTUD2/Av3EBk+hAtos5tnvhyt
nFPXlEdQWL7L1zPkljcYKHz53OS0nyFTHlAmGegE34qChh9d8t3paZ6o4zNI4Oiw
ov9xFdeSYR3xlz8Jno/cjQrr7f5WoX7Ae9+8arxRYXJ4UA28xJxOfd1R7iaJGeqM
jgqTZrvVpxXfrFC51Pt/PfGE8PzoxRTnJ9H+jeGumg1ygXRvQOgEvyC7kENQJqZE
4sGSHH9Izt4iByzeuzNxNmtwq6T8JFTkvX7Bq9Tp0ERUa5TQpR3/gKimSaac58iW
x33nW+pdgk8pi+lEc/4WjrxUWaXAlgVN75Dql6OrRAypaH1TQ3EhVIWA9ClSeoKv
acE6eHmhMb7K/dKVi8wJGpiNDnZAvx4PqNzvwujkqPz1V7BL4KQdQtDR/dNbiZWU
h5DZImyIIQ+UicG6Z1hDHbx32DRwBNpOLOR+CQHTnV116G6Sa/7TnqHiGPTKv+Qg
u9jsJZBuBruXS1Bz/5UjbIhNQUmZ9LdHZP/3QYpqcOgJRRd0IlUMeuA/btgrPACq
8F+pMvP3VSTMzgyXhFbR3SzjfsIDCy6dimFDG+uYZx34w+gzBsDLHnLRPLGIAi6t
7I33CW1vIsJXX3m6+bnX7+uP1sAkLZANIOD9amjcdDOLKLSpNZZNmby4TBV/IEGI
lkYLcKo0rDv3mpYA3/aRBrAFfZdr30VMH73REVc4Cng8QMRxAb881LIhi5qh71B4
tr+KnD0MC3hJl3/dXdNPZnANCJv2hv3D21d+5g4yJv047oGI+fkfgn/mWhP8IZlQ
1xA01Ymw7vOCkNhSeajP2miZhdf2OBuOY4fJrD84eBpURRM/my1UcpwMOYwjvg1J
nGfBpPr+AOPtoUxnDNsTRVD+If18PPCXVipmup41v3NNSZZRtO1KxDVTf1UbEY8t
jO3vay+NpOQXJcoiItL0sK0NEK10a2vJVkf5/bujefiye018bpOQ/SYomHQbpGVk
7/W7t86EfmiYAqSwsha1XxU6Eyxl7OG7iVbrQ7mSZRr/4pYpvOhKBFWw/Wgprilf
HqYSGJLpaLMPqbVMhnRIUb4C8hzXLENyHdwoyo/2mPbjQXqoOfBORqpChuBU+kFj
vVFLtU3HdcgXSDgdAECq121RglAQwYXpueWnp9n+FTlWc8Zb0i2WnUXFrdCcnqMz
LTDWXxf8Yho/G6xRkXFkfBRehI0OPoQRZSnK28RHjEC7WQst/VrFtmO3XGhof7YF
GbFyGimhg0fQ8EzAX0VUwfap22MfimXgwMNoTnw+Vgsk9n9lx6H1cp+dvW6Kjs0U
PXABFnByBufcgYsJLYiM6B+FUwANhRWeGzyDPXqS7DVjSwXQa2zQpS7BY8gxevAF
4ydnPBgF9REJp0BYaEywi778OgowIy+41RUHUlT1Dzn1NjbRUwMtNMXzHMJ3UzCE
o5Xn7TrMBeNecLT6jSd7sgrmuj3AKBqxw2FbUJEWMRnJCr/BIOen7c2NTKqeoIEe
oK7/GZVrzzBfJAYjrWad//TbjAGHxBs2a9Om01hBqm4Q+WuzED0Iww/IVIMpxT5B
zZe70p4134viCvTQOMlA+oxnL48RsqSAfMGDhZnH2kF+h0bkq2NsPkRrC1NcfWVk
YLG2znOHivINDc2iWuB4tNiiLYDgbrjuPmvZK8GCGp5axNOb/tZwmpZIXEWsw4i0
FnSnTpOvb/OcIqFEG3S9gsxb5HgUZJ/Ye5PrK2e1qbz0eEkU2LKjJmf6HjCppm0X
BG+oo985RH/n3M5w3H9DPUPMdiukR9z/G5bFFEhb/yZwKEHp89B4+GG3sgBTvNkA
ZVIyS6V5CsyKxb8seRTdC1ylYg2ChbbfqJGzYk09NtD2A8NltlKJlQHe1BYCS0SY
6/Z9OQCxDiNzF/V1pMBleBQ32fUTRNlg3B/VdiWKJMcKrhWqWxuHzSCXnjzZiiGt
06sbGTx0FxIZz+Hu3VO6IZYypqB+iwBC8GIBrnZ90xheTGWTI2o0qqhojqmbZPGb
+2Hrtw7leRXmwFic94Ippo8B9O+UjWrBYEnGBio7rsx5kRUcB/Qk2oI0FiI2dLvd
1Rt8SROgLEyci5Gz84ZawGAEnAbmaAr9wiKOz89SxmzUdfVGQ+4YLUlnsq1mzgiE
NPt+pMibkDFnPpxS1ka4Vsv5FBWKNzqQ1613uoqWbinCFau9Hy3OtAhEXH2Ae+bH
ZuBAxptIZeVTBMp1UcxdVaUB1Zt7pU8cHuqk5hlu7lkSeUbxqezkgXBeRfAeSJDR
gNdg9nL+xxjnzRQGrt5tHA88XXa/KcdBdktfBoEZMu0etT6/QsZVWRgzfgOGUUyk
VHfddQkDt2dHljt0pOq6bCCdu0ORaoM9DeVaR6oIouuKW9O4xj3WDuIQHdmIvOfd
n3U0qSkJUaSE03RmUOLyg5lhMm7RERDj0xv/qGQhsHYOx545jTnQHI7V9AnCWjek
b3QJddj3g9tWRvSjJNBlZ4TsXLoAx/sP8QE3hio5UT6TL+Lr7ngfvMoKQQYcTQyV
nFVzQ+oiKjqxbqfATsjDtOuxFuJ4IETEIZ/4pwVqpHxdhtrFk9FEUUVB9gxceiA1
CjoVJ0XbZVhZZ6ZlO/fP4E56O360oe3shn43bCX9K4XvOKBoxeoboYn/Y9Avp794
C5pC9NxDCLSGbLThowHCqKR/OnaRqz8HIF4X7FGO8n8ZH148LbfbFX93vcfbP17Z
vlvuYjDpw9tgy6FpT8ZMvpvNh6TMELnx0i5P9vJ0R6QVB8Pzu0hwc4Zs469HUMis
zAHnYVY/RDICjZOLUqN+jKms7mR49kjZzOuWRv3GIuRDD9R4+3E9ehakhk22EIi6
3/ZFxsoHR3JJ+1jN+LJ09cNAvA2QQV5Nmlc3cZbuYlTsRodOkjgNCVWKvaoY1+yP
ZOIA60fybVZTvFRSpwmQwi9nGVBDt64fs95B4KfgIBydeMB4K+FyVkFLCdy40hD2
Jzwgw+PU2Zgyzpp9E0+BAv14S5nQbnln4BbhqjkhFeUHlAHrbUZVuw/grQvMPGer
psI+qrzzm8lbfFkWp2ofnQaMsMJRRg5rohDxirU1/kDvf5TeX+z7xM29W/JSk3HZ
vGIYkoLlL/o70wyLZ432cbjJ01HWuaFLoLDDaB5gh8JJzINLqWX6XszCj3NsNtc7
u+4ySunCg395N8hcDk8c+wE5IonOWEYw7KpBPMmgZKeGupejgDBuyzC3cSVGTz+y
3aawDLqu4vT4yJz/HD87EiwPEGk6OUEUpKolMbDN+XCY3psnN+lJjPlQ7Aj3jKMN
Z1umMv99mtkeExBD8jZS/8JN0moLS6957I6cv9htCM86a5XYYMPk65HnjjxCEFbr
HiHpV1Fz7/c1vrLVgNPTwTMR92C2RHHHr0vIC8lyUhaMC+pPmXxd+oEGHpy/7P6F
FdABuWGXCCzh26kvev3rzUV0ve4NyYmjUiX1llL6yqioLCB/cgDSvNPfHtXVsqOW
DkatCQ46FLOxQZT+BGE89eKs9hQedHSNfnGAcqWpQv4Og4rarLJD/PQWPupDo+47
IlZf8Qoy1vmfOc2McUX+xI89nJWXixhYuyv5Gv7deZAkdtVjw671WHryEBFwlleD
RqXBlvwf+w7RZ+1OIcyCHtuVGwatmAFWNQpb6dwFd224nFEwWx6nRrjzxToqwgO0
95OPPqotG1QCryCq9W6BfA==
`protect END_PROTECTED
