`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ufAT0kjzxmyNp8mXxm2ymkKeoNKS2CRgUrXHHZ3LLpAJQlVqCYQlIUrBeLGZrxi
pHt/tOp4bEEmrR5sl2N+JQC4GOIEJMz+JsEyW90LLpABjmJ5NGvxJE8NoKiGNAVW
RkdendgjjT6Bceu4EC4+47Lzbe+M0dfaKrShbVHkO1hEmBwF65B/d5NeJH/g8IEG
sK+FQ9st5nQ4TbmjpmK2kcRDVWus8lJQ3dViq7nFqOiFLYDpgDbr589n/w8rCfO2
qF86qc5xquaQMYApXzM0Ea763wC63VuIrXrqsHliP0zYmeqcFcfsAjpnGis37wyi
+8jTLjoTU0x09AiBXL0+0D/ZYsy2v2TChCfGFOVVhJKrfZi0MglIthbRGgApsIb/
Vjj4G9y3r0rV8R8YULgLRwrulQu6FekR26bPPTRNAt/pkASlvjKJNLRSekVZXbtC
PTBxfbNyktWuQ4gFNbGJB02FNOyYAAbg1yW1vWT7QdgIMyy91zb03adKP9+s0Y60
`protect END_PROTECTED
