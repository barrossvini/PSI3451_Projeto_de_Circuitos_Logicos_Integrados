`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hDbiXpVowcvGQCJAEpTlqLSmOpqS76mlzFB9dy2L3DhOANf5IqiZa9vKEQ+upohL
SldgpVK3NfeyDjWUef7cPfiT8vx3qXHDvOqSdFFKm95cdWtnUieb6EQN3G8ETjxV
zrpgXLOCOHadIxbyZ1tnH2fNQNKYAkF2OCGOcwEeXkskGAPpAVIR08rOoLYIQrGM
DEIp3wV50CvvJOfh8a7wOgh7GTFS8tmDtahB5FxsL9+3VFUchl7JC/B1TPwn/dSG
1IHusBbpdtKJeJpVDLUkzKzs1EGWrsDE6DD/5yn8Rpw9UnVFBV+oMqDzUKYivWUs
wqjxVqlYgt8i/jKYaLo1aIXez8N8ddxkeEwE1oSunxLqgYnb3Xmk0Ph1McLhtIxO
VKyraLE/ka9RuicvCymsmnY22UC6Kg3rY196k4HzoD/S+6fOER0Vi5wvMR490/IN
r5tgNYr63u7A1HTwLiVth9k1KsZ7jDSghGbYt/jiqwgBaXxv5qM6HFn4s5img2Lp
aPfhwKJNvztHh7/8jY7rHeEDEA9qd1SMa6DE7ttaoNtqQAEJp2qr6e7L/uNm4lZU
QccDOIw2TXif11F+39YKpcPtuuGl+JGgcrzO8Vqcn2sERO7PxctCO/x852LCl6Qj
tu/n8d97UfcAY47StTbVw5syOUjfrRrnIvofv8kGd6t5CuRhheNnC6z51Usq1aQf
gIaR5SFF4G/qmtPOo2tVvsimbn1u3Xcon9ZE0FYsZXlXmAvsC4ZlvYcklhA2C7ob
NZIBOaH0mBl5gCJ49V7j3km5wcZkQ40pEw8f+Q/bVrpinVXxHy9bIfHVjkmhpcUe
u7ZnWWZVcvyztOuEbe3pwElgwvfqrMst4+D0aRoydAqyVfvmakWKQ2PwT2fnDNDB
1bKvEEpYn2wGdJVOBzr5IrY4DF67cKokKiyC3CVOo1snWDbD86ZBXgGiSqgme7Uk
S70afVZcJgZoSrkRHLftzVcDBogbGYgcNXhO6sWFnbco7qm8ifpouSHoSfnDntR6
eqcrHXt++m6+dhROXFaKe3SxqmEVOTDbIK33tW9oC8930kuuiOjcdj9KR7LM9fff
/9GZIVzB6tj2oQWt/3y3+xDFYOQnLvAR0n9etrpvrAY=
`protect END_PROTECTED
