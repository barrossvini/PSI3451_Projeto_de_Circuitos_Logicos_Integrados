`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uBmM4ICmc+qpYs3IUSx+ugdzCF3OUF7AzRG/UyeYCW0AVgbVJy7cbf3y9JiLI5K8
PsRYA6wKRgyUU8Fat0G2irltXEtJIJziOgXqu4XhpZv8UVxBD9ZM4+s5T/fgQ6tc
ct6/gd097YJvaoEB8REa6FDIUunjyiG9s3ciiVGYsC1BIIYnyz01vwBu7QTtuGY+
f3S4lnVt6wvh50LNvXUG8UZOHS9aXcswfjuQh3SxcssC+WK/eJ2w/AOD5M1a6S4Q
fcHfdNeRdU04xOzvyV4dNSgZyKtDsY7z+iqC+qMdZFCI0pfT4aluJUGUuStXlNkx
obE2gtQeVFCGa5yTZiBtj78n3bXJdHvxhNnHseb32ep8DLqcsrIxrTBsSJWyT1qi
752/EPhrbDcFyta5/Y9Y7NFzwuL7NdZjVb68BncMuVdezZBJjFrjGSx8RUZXIYe8
P7oaFCWA54BEUJx3/xVfQq+2ktHRD4P5codI8aRnkSWRVoTkDH6oMNGcs6O2WcwJ
K4MGqnODI3a/Cq+JO/HUsVZCrstt+bOuC2wrRvyIHYRxVTXRjd0AKCd3X44E6pHw
saOosl8U5sHYEXUFdG3E78INGkORI2rG8yBRcU+4IuKwHikcbd3hzb4XKGZl9Ncu
1Z8DnRZUIrQBwBojfD9OjQ+LOPSAxnQeEBcK1AenYRmWPeO7Eq/ixiKzW3n2UQM1
HUexMhP3bGmIABIis+ZZ9Lay6v70bTnXXfMIzuo3MB5eAEDvwjeH57GMM3n+FVAp
in4VeMiJtpkna2DbB0wz7uiwHHrrLfRO5yAJJZxtIuC/khNdPzTvIGaJjKrhRlsg
moVEelPH+r0g4QJb/MfkJkkklKi41VWOiHRh6PPuFKaoAZCUTU/VpeArS+7aL27U
24LPMET5ZGz+elq6KkJFdTH6JltnoksKa/kRWhuD96JhFDxV0bj7GxZzVLe1FkYS
arA/sramJJ87tloWZcfnXysyJ4SuhQA60Bfncc7pjjM2oHjsRY8CohNLx5K7DUTr
xAj/Va5XMVg0tPslkMILILSkhcrvS1WrakI7Rm56VM0Hx/CrDey2qgRxbTHMfIga
381y7v/Z5060sXymVLJAMDdabkKfEzzdGke+2LMSAY41XN//jwDHxCXJk7f1tZTE
dBW+oNge+YYfb2QAcuY+QMdXR6Khl3mLUcc1/T4OMNOMBTpE1GnbR4D43E1VUsO+
nlWcCbxMFdFDUKgVWWQ1jGkN7NL6mlVvXhszYiHG7IA41XVxW9IoOs3XTBb1UIvH
kre13Kql1lL5l/JP6Bx2EAtMsWj232ORgdz358vX5TmAlaLeU6gJcVznqPMp2ZOY
fuNzccAtsmXCwYXJEGFdTS2dNYXyzJJ0oNx0+dxPrmaUJs8JgJkdKmMz7s9gNLmt
3HidG7WnlW4TVD8bGg3BNWlz56DUZP0vNLUVm1dQgo9yBRr45BXEs/FZF/Myo46k
VHrJpDuoCFhGgJ2VVhgiKeJAaUrbtDKaHn4Ug34/g1Gc8f/5nXZPnYHE1+eq6uIa
V5GShdlbk5lkiFhI9YjleOdlisWJz3f2FTi6yajUQZsoIUhZEz3+cyO57QQFtnPC
RHZ9bnPL2ZTMakTA81S5zRYDzKVjYepUyCBm0mOtT250OLfL6rL5m4ptcwgzAaiy
82K5Iv9ntlc2P+zvFCfokkH6nU/X359D0zI+2qH5vXAcnwAtgF/gnM/KqcQoLbmq
DE0l8Pqcetj4tMrq3XlkjUoaYxudKd9BErquAJp0BXjmjMErSvGgiZ18FGLZjqLA
ptuhMylEg3qYADOsKJ4RvdlnaKHOydn+wiFJPb8436IbTWz/sOW0u1AgH3+ZbOGh
g3s8S8ugmR+SgfF/xg7GRSVw7SZzd5ACMJh0VnTt0OcnoyGWFbElpA9EarTzzGGC
`protect END_PROTECTED
