`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QRpd+dUSqQSE5KL6+BK32Y4LPFRQXo5tjIBqBaxwYGzXKirYzTOSqLCkDFHuWqP6
wU6BAj7szOA/1fdcnD44rIDsAyKEx110s1qySdhEveVp0KBqXpnnTp0HcPyOrM8X
dbjL2Cmfij9oNkq36SkaMS7R/bsO479YuAq+vS9pQrnTy+vmGaQdq9mH5XHs2jFL
2fMFD/beVDTgPgHN98razs7BH8wRhpKZcp8GgsIQYoT0oVDrxI20eGQ8f/g/BwQa
St7Qizubbc04lRfGlLmlolS0PXfBMYNXpysS2xYV8qvCgNF8KsdI4QqxZ4rvLlN3
1a3ddrg8Ve8J0cvGAqTG4j2o9BMsZywMHpuQrHIWMbJD9LWzY8I9IzZPk/70yj4g
ReDKDItXUQu39qbxREBfghB7xflyVKrWgRjzBMCW9XJz0CIViGiLElrJdbdHVXSI
Py1rilFJtkfAmgBFhN7bESPUuYqWiIjz9CurrQ2Imr/A4lGHCHhObzg2+0Zc+aA9
`protect END_PROTECTED
