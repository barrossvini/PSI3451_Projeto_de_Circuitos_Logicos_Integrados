`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDEVcSvc8APlsonWlycBGSVtJNmIrFkZ/7kEwcceKa8vDVZ//u7ki+OZ70mdhPb0
QUz52pLsf7H6ZaA3nIk3MQat0Xy29sSGYSqKx53tzQ4axWiMSiNl29W2uukAQ9W9
qW9tvUnXVGSOekX6i8ZqEb+RYeh+mIteRZ045AVHQ3pdPk5mFR6Zj9xXVD0lZpzG
ex+U8jwpjakL0K33farsaD8UTE5vLT5fh5dHFc+woTQK0z5tkXS123NbJmilEb4A
9uKKuUF0SdLSIfMf66xAJhv6XyMVlQKxR8l4JzNc6AZQiII3unVor4Qra7/IEaB9
XYQUGM2c2zJiVqKPV/gugrKTYtn7VKWUEINkFqi7A3sv4Ztr3WDZjUK0X5C2D1wc
jhp/ZvDh1z54jaZKpu7pBXmB0chGzB37wL7A1ZV9EPhCD9V3V/I9JORtxNeQsxt7
EXBt9f0e+RT3nLIYBuFowxSQuwWYSpjud5/XVDRrOlitCH9a/AQpwn+1xERZVAqJ
euFqoA4u3KsPGKJzIQTUMdP9fixpUzxpTgHJhgyZikC70t5O5JP8z7dMBZlv9KR2
oyspmmTuFroC4SiEbpFICEZfXbTQH2r5W2ujDf5lOGgjYP36KO7oQWPy5qWyZhbM
R7O6d9nislmlHZxdhUroun5nJGp6E3UdNN6O7AwfEJYwJTXSlfyStATxklezCcpR
P5iMW8O5LPygZ+bqD668b2lygLIIzbrSTygxtycwK7pmUXET0Uj3D/apdDyjkzCk
ExvRllCmBEAW994vnpFvD1FVRccfIcYmE7axOx/HENkynEw8mlmd/FnlQ0BME9KR
SniAOvhtDqJ+vyW2IF5CLFFRkqUMN6VTLxqOKOw+lVglrb8QvzmysCFdVLAs7Enj
hXZEuBIyM97Ja86uU4gcmRUIh6sHtIaTNUQ87zSK+7wcYe86bIpPVtODj6aKj/83
ahysdfiV+k5NXxCFpicjHJVe4B1BL2C56Hf+vw3A66RXtwvzu6fFuwa950hTf/nm
MwThib8XtkkezzW2UIWD1NNrwJI76aC9jckOyYwB8CPQ/ds/CVMXNone+D6ll80F
1paDDAibKdnuJcr9eqU7Mf+X2lOhonjzfpwR+6ITXtj7Wt+7u3CXAztRyY7gNgq/
rq+oMaIg3B67L8Gbr1IoI8QCFHTHdm7ywxvtadagGLNv5KMz7MOMNTVOcpuwIl9S
Zi7KJhM4b4in3J094NrSWp5gvtPn2FOsrnBXfCgsJcl2vBqY2mz1dFmEhsLCFHyJ
`protect END_PROTECTED
