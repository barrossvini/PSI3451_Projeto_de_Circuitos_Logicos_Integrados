`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kxm+8mxARM+aMAA8vs9JErtNjR3+zhvgxzQZAUfZCSkQuUkQdnKeYqlz7G2ByVKo
rY/8Zt0nmUEYfmwTuXL2nkSrcO1UcoBas/e6LHOA+jGTLQl9cpsxVPqep5IdEGRC
M2CFzu7EvniqLkZ0RTe2yrAnZTGcc9ioQ4JH44wX1+pFGQ9wTFifa0m9ktG8/4k0
EuyrpEnMn6o8tOmtBd8HBWrtZoQOB8FLXhVhfByCgdwZuSxBm/hXqrUis3Tok6EI
ridv9Er0ifBzW2fIB/idRLIkye6LUYdXRqll8pzEiymBHRGuC0WumU+kpeOAjJpI
UMvZo4pu+bDqfvYOVBtZ8Q1eKgrdUBPNwoPjnUTSt8fTmb2xX6++Z6pX6Z2rzfEG
q+BfHRDNJCZqDAF/qtzEYdPBG0SGVE64ddZqenqiDW6QmWaWiTeMHjOKIkMaBnci
HG0p1hj6PVXhgdq42cu6FVgUgDzEIEUzjNWGQeVAzNFVGiTQ5sicY7HOMTz2Eehr
nNJ9JLFn/hQ1Vd1oiG78ezlHHcva9kENPDUV82Dk62XAj1LD7XltGfvwwD6fhOHz
X8BVTxIjT+wYAOmecs44x/AhZRTbg6KXD5wSXC4eXGMIByoN+jKyEtfa8rlU4ukM
d6wkdOTQdfIqPi3f97swCfmXJnR/DVRy9ec8YOaI4Zaj5JUS0Ds9zr0/JLfcbhO5
9vH292B3MOoPwrVQAE23PtSs+QlMo72myq18hrloRvNperWKqvdl4mLTb7ZvdT7y
/sZknGeGqkMW8V7vtRxX1rqsYaCkefHQeYZztsSvmYTWzl3S+bEHHgUvI5JGQs4R
5GsBekJOwqIlUK0brqhzh7RpEyS+lVueR3/WDfjzvu9NUtmBIC5YBz7XNH4KPezC
fh1DcL/eHlxB/gWWAukWkFNF76PB+spiXm6VgZhtByJmvDPNRB64/Et+wvBUGsCC
8BKD0Hhi4B+nwfpqeNYWdHmwyl80N+Dqe4/UgvidAHiH4DrcCRR46+bXwhQKGQcw
iiWCehjBr///F7JFMRjhvnYPFKAjDo4h8YXcwpUTjSH7lRpczSYO2UbfEHSrIH0e
Zz7n8QEjEgBE7nH/QZ70Ph08FW7zGn5sQWc8wLp0nQI0+ANirrF5ytz0tisr5n+s
5n2Ggo1XBhTQ4ewqG8pcCw11rRmaFca8oWtx/3QLr2IE1E0eh57p5kvzECA0UdsY
oHdkgTYqjypKCxI+MeJUiyXgMX9sbApRZalrqTwH5y6teF4TcheH6Yb6jmBntk6H
ZBjIDSt2EM9vJHEn1cnfIbFLqkwPUURnC7Lq0XMQK+eCUtd7G0Vb4W9YXmFRHLPE
6D6k7U6RadS4vemBpeEdmA0gmI1G3NyvXhGa2pq1zHUYV6HcyRteCxy8Aj+Fa+6s
zJ7R9985vpMsQz30C2+KtsQUH72UO9Htn1tqIH9T7Dp/2xllKUdXCUE8BpQUpO4x
zg5ompXq7NZCxmKycrHWFVVIPdHFp9ZMm4/aHtPNlsyLZu1LvdRBIzwZJpi8yd14
7K5967QICUYsB9jwRIkfgX62q9jFdomI0DgnKW15MHY4xnbY/EgrrA3EUoU0wLKe
gS05ZVdnt+VxY6CfcZdBhS6c9JD6yTZYocmXdemxqKdqldnzaiYlrPmdG4bLT9l1
0uwJcAJsYDBQbNmlAjr+W5OWsUqxRafC5wXBfBz0tOiMQVC5qR9fw36+uZ5ondu8
FWPKg67aEsYOu3YLPr6lFKpW0GUGgrdE8DQrxS332z9pZOE2ShX6ree0cY92akBB
`protect END_PROTECTED
