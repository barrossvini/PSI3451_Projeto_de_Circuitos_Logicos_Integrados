`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OSESdSwrxAInV0zL4bU8yt1UH6JzU7PM0LMiDnLpzQ9alzwqilMCYZ0JxOaxSgjW
+ZNpSDFhna3UBRbBe54Cs1TFKWF8Rz7M1N+ChMSAW6dXaAFNXdGRDubtTjxhsxmf
1gtp13gFgNox8Cl1+avWJf8lt5v+yImReh1s/vGSFHB6U3xCxB8UxHmqBkP8mYy0
50ahZBaYQPgVpzYpM9rNXL6uwEEuaRAYyoNCKnDwXR8mqaKRSszIOlF4QXQBR1wN
mo15h+XWmjfGvuhYQ8uVbEMyseGjl0hi2brGqkwURDKbv/xUaY1M1kbo8WobjWEn
HKXebbXqM1PlOgbf4nrLD0sydKR4Vnp7TFZyIqkBPNn2BiINfCiu9YkV15MVIb4w
arigrRTQDs2hKXFmCeCutsTNGkGQXZkVs12gMttKwLVv96yP9T/4t8P0j0GYwIWT
pBmtXEJDM/vzrSViwfbLVxh6skOaQuF4HzzhFuR7HOdZlVjWEZ2MXq2DvuOvH00Q
iCvwBc74V2Q6Db6YNarJObmZGt42t28fs1nzWPMM+GYZfVqDIWjv1tTY/SKaSeZZ
DLg0tOvtD1Datb8HK3gQSXtj6esG0CygJxc4we98a7I=
`protect END_PROTECTED
