`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FxOGrlOxztTqVOIi8P+cxR7BmiYwnoxvyZNyOx9UYf/8iv4+En87QrwLYL3pjB1a
iG5xOqZivm71ljZypPsvtTiDg1aWUPT6Z57ulJ72PobTQNIJFQvQ1FF6tFMVRbbx
JgvELZVsQS4BZBtMaxNC7Yx5CKg1Lh4D3BiADdFkBcVQFz0aQdqyuNpgXiqpaUaU
gllmZHx+TfCVyWn0eQx4WBP2jgk7MIZk1Ysbzgu58UBiaq8m75h4TBxz+OXbyJbR
pHDXMuC2+tpADnlMG5ubKSPphDNf1oJoGuh24EYtT/YRrt2yq/FkU3CXcwRWW4bX
d95ALVOZ4SpYnXWzalGTPhWbB2U/50mt48j78LHelWynaeGB4a53OPhLSFhikpo7
BQBZSF72GX/MQhI5E3TMsFDZzONOVp/z4+O1zpJHawI7O7B/XSLvp8KBh9Y0Ytmv
FgsfHnTxJjeL2Jq54bDxt6Ojh3eApvA/tVnwGAgu3Fo19Mw1ZM+TVgIf/2WK3PUe
pTSQoqzr7pSFDCrqpoMsAtwsqG0DWh39iVeiVUONTR2mYMYmqaBHArm24oXQEWIz
RHnqKgqnbz/TStOm9Y9L1O1ByLU7O7csWe7t4etWvsP3brlceUvRJMcoMCPBwx/B
UHCu3Z6Ra8QyD4Xq63NgItixEekoQT8gt0BS01qp9K4s23MZrSX3tEV+4Mfa0TIJ
ySiywjFVZ5E7qIzD12hQMpsGFs1RnIH+38PPXSVL1dhhmnRAmmFmcT574aDxWEHm
QIOretNx2fWJ21jIWW2y5sHo3LVw5F0SJg1Sep+62ks6baCILKWbawlYZv5aYJC+
mBIu7GUtzS6X1X7fKCSuXU+Z9krvWnVpo34NzFHtf3Vlihs9I/nnJNg2psb/AMah
F3kVZJ+ohRep+p/z0QWIBpCk1CQmyC1ju0GsrNusFjDKNGSSBQbYuUegqxec2pQp
g+1tLbNurlff3eY078UuBqGZAOip8UzS8vG0c5D5JbR0+rEgfCLw8QU1eHftiBJ3
aXysXo5239MtjBotgEWe1diuQCTw+w//wfZzVSHhb98+gTzB8avyvWWzGJ+HoZed
ev6KcOmJrm4B+QHYNnimaoBtnRmo+C6f0+l8fYIG0uDG6i0tn22ItW6NrEGElrkW
etpaTYtFfeR7E+DvomABJG3KpZi0uvw/rCCJAeItgd1oZthxI1uTnC4q1gShn9EY
GpkM4Ow96gVjAgOjTsCvYj3rpQsADGyxUQB0dd6hNiSd5zwLt6yAnFPgBig2EXln
x7sg9TZ2R7uQSz/Vk1RZvLLFHoqw0LSfSe7unM5bhCAWYjUIzzr1Tv7F3mV13RIZ
P8KApCNXzH0nmJ6nLu+raUgDymCy+CRyvEvqPJYcYwVC2TTpehwy/vAZpiyxlQ2O
BQBT3d+fCTEQbvPleNaThpWmVqPKUUB5eobouY7nvQyNSsCVwy9plOMDaCOOR/d5
SvR2vUOCEDDEmbONMZP/fUrKKfffU6hflkkdqrq8JwhjQvnhk2BeTyg4Y5zL+31L
H4jXHkZE9U/upX7vNzh1Ig==
`protect END_PROTECTED
