`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CZUn4ARRFLgS96OuZQ3kXOAj07ATX7HEhRl/Evg8JOrRe8pAcx7y+zL4x5ebsxKP
u8UDP7l0L27QUv4wP56wLZQ995Yl5xfDsFRVR50/JYWePqEZ2XOhNhoIrOqnWmmk
9nUd/pj3hHQb3egGc0ke/uZvEnJ/NBu/7r/rCgBbMSJbEl0zZ41TVwWP6T4zS3tI
KHm1VJ7WjoYZVgXAeD75H9+SvTiw/DZydtFtx5sJv95GAgz5ldk6FhuN1EcrYlGe
1w5o8FkYzOiO9VnkXYFhpe+tm+95doOd3xR6oGxvc2oXENxboSC4ccQWsHeos2ZZ
4E015e/7eP2iOM/efk1aHsf4QsFYoDRxh7IwI1Tu8cqfTwSWXMrRwTMUp81i6Oas
pR4X/Ix3yaY0C+FwA6aDGqETCWeJ+g2qHQxXhlHUIW3thepHw7r1eCR1oBncnNQv
wvkWYHNBxM6Vf3Kd2OBxFYGuGxW9IESLYJl5Sei7ujBXuVigPda2Acs1sB29Xp1C
0XZtUTqphPdLM+ClV5yHZ8735/RAw5zoFAT038w1JvbK3g103aVFckZZ7vfWfFq3
2zQX301th+39Q77czOnDbFhsDNDugvsTOgVf+OzlmnIAfNc7YZpkT8xdKmgAMdyf
qi37tFux7QJvGMEwNL0d/Su5zeItV/ccGByBvxr2wiHW2nzU3UpIIlyd8pOTobU8
Dq+s/6EFusFctT2mfY/cxndelMTbAS9V5Q0d1ZX4AXlOB8JwKkYQhMVmC7MUc+lv
WUpBaOk2yOXmlAeZAO12uQ==
`protect END_PROTECTED
