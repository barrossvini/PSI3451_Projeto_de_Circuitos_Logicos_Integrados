`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3SpYMYzEIjBv++AlMWaZwxB0kMPtJcxgJFqV8C/iZDU+iRczA526yhDuw+nYfeXO
uzt3dnSWRIGqrMjVXl7lOUW6gNTDC31DNIkwxpluXgr486d7KR06mb0XlS444BY5
O1q6jA1efIfTvZia7A4zN2FM+ouq/EQsdmuNvs5MLrQyStE5xjNtcatSLLirsypI
/DRCIC5/74r3fJVjKIJTOHQBKKRLOKPDzhxOW6ewY+OI3jQunUKSNlleKtJtaClB
egZAhhyzBuYeEzulx9uyynBFcQTC5b+hm5iiYy+/anau0yIMva1SvnTb9vaGuyKh
pBWIp9gVXMq5RN3xqOvF12yhIloxgksh7gxRnqM7iBQsbyw7vuywBtRinPI0ZmmI
xS2yVaWrAW6RgWU/ObptZa8yX32VbJL87LwJq4vnWMiN6zIyFY2/91lkxqCKX6dh
HNOXlplH81fdiWTe4SR2hM/GppXNpCSAZv59rt7Jf0KqQFM1QwPogJYmupCng+2m
fkBnCAqU+myzvNj4e+j6LmW00sMfa3QefiFMrE/V9EquZgXtl1cU2qnncrmpTXfo
4MG6ksobt17mi6F8IocKu4lrU7FM8KcXLQQ8e5HHUg30VlTjFN4JY/xUROO7pSOF
vQfYZ0wengF1ZakeyNfsmgQrb2dN6iFuEO7zy+bs6TOp88lxgCtHstEoci7Z8mKC
euxaHEYb0YhgNfXwNOdxsPdrkOeRkjrjvoznwifq+GJQs+UobptpjXo2MVshzkRB
YO1DN4lsyZKX1PoZSjrGBNiRGSESXxWLZlz+BxlPItCy6xieAD6MM1boQ8uCRTkW
2fZZoBgavO94AEQE0r+KXCElVQBe7V5O7W1g1EWOQ5fxcTMbzPf/hutf5kpidL8D
Vk9p3f49bn4e9FU4/3rIH8NS0fARdugu9zq3bfTuJ/Oqi24/7SrEh2zx9EhtakRt
Pcamz9t2d7puTg5z5aB++6pkpf4P/NMnOsjKThb0+0NBNzMS0WEf+cYBKRlJQxzO
TWyHwkSmYfg0gzA6KWve0V5EDLTYP0g12Cf7cQmHFrB8K6CDPgmehBASlhtgESRV
l/UxJcyvmsLgVOvT846LW3oEmddUuZIOWMmBKB97czOJc10B2jQXTUE7zQodInyL
IJLvdPEOthTgxpPfsTlM56GI0fB/htJC6P9Wsve56SeoubtWvH8gpANcjlXwppjW
xYurTPGzPJXf9BP2ClnluYA/KKdeOZDRV9vVsKP2BUithaJfgpBoMz844ZVZ8ctS
X2y4F9mSFFnty2Esn9q4esd4roWLeSt1YPJ+9VsVrlwQqafzjoEUpY3uO0f02QCw
xn9LufI85f5XfUqiHhiJf8EUWOp0jRwei5hBXhEYpY5Bz5oq4uLBoHzereTSjVw1
/FvcM8Y6CpuO4SoxnD9BV9WvYLX2+jV++OaUoHLLWVFlM94pJbyTBW6UCKa+qY2G
vKeGcbBHvXYi0FW3LQ6u8BBcW9sc3nfnjNP+cL34n7VwIy353VMs5OMQdTANdsz6
cCzpZgCiLCzC8VGF94O7fN16iyAYavMuqxhwOQr8qJ0Q/t0iYQZdWEBFLgGx2x5h
Tp8Kxn/gj/OyHoWIOcDz36GNSgc2UbUHmcK9C+6w4/jcZC2g77lZEhn+5X9tPLx4
3Gg3NRWhBwB4aZQapSfXNsfoMLS9c6RsHNaUF31rH9Su+HbAGaSFDWf6lXmz+hU4
dM2TNFa6C34pqp3bnD6zkZPy0O3clTUxFD+v6uW63OCuzc8+qPrc5wbVvUhEaIQx
KsYSErujTiWbh36xVoM0OAaWXk8IRm8qESsVKmsj6w/fdP24T1h9Iik5doERg8YV
l+66wIWdrRW7eVtWMh2zGtOGk8SJCU00UzT/+PCdHKWdUxovNS5i8YjIKhPlmjd4
NsHvTUvj/xWoLkPsqAmvlaSm54pVz5KQh8VGaZlWos6S1QFta1GExKZKnywchumX
/iOz3CAM9An+6QU04rUSVz7orp3HtMG6PLNI40EHSuDcScQnb+nya6DtRecG+93v
WP2S0llcBA4QGGqE2iwleajxgA/k3w3xCUMKLCbjEncUP2CUN86fayX6g7SwTTh6
F7fZ3j4V4xbco96y6ACqzzJCqqlmXsh3je+jYan6mxvkQzG1npDWHemwl/3IYZob
QsRearx/gR9gzfVtl6MblPLieQsmzA6eaxAOjvXFxzBXrbVJOtSu0Nw0OqZmFQhl
FWMCGwULp4/Xxy75lvtdYSHHdy0ziD3mWA6iqxqZGQ/9R8mVbF6bIRm74k1k42Wa
SVA/biIrazCz1vh//HcVTqpJR8xqw8xluohNojb75MxaO1DhWQPsuPEnPlTFfpYq
u1cMS3hDrmgxpUlxX9vSDf0tHNzW9hsdJOa1KglqLykmGE227K764r5w2T7Sqtpl
U7xJCgguqzEoPqwzZ8IEZGUGaPSpJtyFNPyuLqUuMzaKZd1LHpBcGaSReysSQGAP
/nf1ds2uGBVAIO3sIfV76uWMabuGVFNG1XVCc+ZrbQj4uP4o+tpf5gEsKeVciE/5
YFuqbcVBli8ArostUdu6FXKVKpbddAdNmU1lQJKvxYpKyr+TDXb4FGoPhVXDjYww
F4qKuQq0GFQkO7mN/ouWgi8Pp8hgr9MDIdD9PpaRV683rIaUj4PBZJQQJxNfI6Mb
QYiLsIsd3x3AYXS9bHSk+wnZNs6051XoR1LTi8vQg/wvVcO/MAcf0IYSunpuTwp4
KQqW2vLUi50/MQIEgF9OiXP/ODtIusOKxqaJApyWRRGOpZL77+86MaXfS0ajKykk
GNc6EQ9/x+rnI8BpIpd7Gg75GC4j9k2ZuQxMIzcBx1hSZJ00y1aiKF3aUsbiyaSs
e5dSnR8tX2Uk6HbHyH/tCrSgg6VdmPKguvdYdsNHMTcBArPUctcRdctbn4tZEEIt
tgSYNasJEDTcPPbQcu1MgPu/QN4qu9KKUxY8bRciuvh86a7u2bA3wiY+0aDXKoNQ
YD2GTruQJQY9ix+5CZx6+gRAe/4KpG50P3wVu+oYuN6+LlxPr0e7Qy+YpWBLzupl
jq2vhDxQ559w77ClaY0TDS/d8nu0UsN3OOabXrKdPyhw3HaNGKycLB5PpSi5/jJl
akRBpfd+AWYU5yatjSU93mPW/ntE5Mq1E8W4nt0SZWJJveqtE4zHoD6q/Y+JQfPe
cpV/O9KXvA4K+O25iPo+MGRj7qpaZ8l/PyZ/7boW9JTtQMBiqUTxhPOJ7rT0S425
cR9+opLl/S6WIhxXcrp2NO2ZUPWWUHF0WaubW4ZKfTV45g8WSiHDoIQbz3DKwBp7
LBRcZzPMKJPPZEVjAq6opFPHXXLwiCm1h542lI7IklcvlwaHOq9yBhTqg5bUroO3
R67ud+LBmy3CINfTUTQ/sUIQ9u72jeomqe3jgG/KZbo8uQ8yUV2G3hhBVvT3QKy2
X/7hA8zY4hofI2HghFn5R+Kftba7+EJ5/iK6hxYuWwBVbiZRZw6YsWvYQiM104zW
nn2kmxwijgwtregGBWP37ggi2qk3y3lRN/+tAgh+xyLPjkDC0JVkzybIFdzuWdxp
t/rB2mJrMyP/J+0NZ+79shxugeeTe8JVEJ4hiBD/XtiFEo2NxHfodMskD04QChpo
xD/Z+35T8BvRLn0U9HcwKQ6n3dLTIYdu+3UakKVHTjOJCWAY7Okky3hbCLM+ySNF
kmo5d6e8hv9jWJ+q7fVGMg==
`protect END_PROTECTED
