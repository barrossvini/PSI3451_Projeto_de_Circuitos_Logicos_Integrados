`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GTJMWXgvSOlZTWFRl5lpSSPfL6kK8GseSwu+/UjXndNDOjmSu5sT/4qjh+PIFQLY
QHn0t7vuiZvuxtMeqj9lyxdK95Qc7uCEoW1ecHycn0Xg+ibvACHotHqhA/6RQfi8
IdqK4bwMLW07T7fWym+nr54C6IwvCrK4mTqL78C2DUaDuoLjxA/oHN8ShRiVrxKF
FTjQoA9HNKQCNo85Kl3LF9pPwflxTMdA5eTbS8tIooIvbRO+wF/rL/7X5fvyPbmE
Ef86s0azjnfBl2P72ixSCHHhguuZf7uy/92wniHfOQWTVmXoKclI3E1HmJB/lHKh
bw0+H+Gwx88xbeAce64giW+r4UwJyBAfDRZs+6zHqwfGxuYOCTE1CH0Fo2Eby9Lm
UeMN7SsXNrAGNrGo209TNlHCpbYJ1JIW7hCpC9mp3/zPcvEFC/i/XqSwmx4oW1Ww
ZuytMCJKQu7d9S+3ufyLNYtJ5cmFzbOHoropyP9s3z8t/6ZEwc3MnQ5NIZNRphCw
/U6eLmsp0HwE/VZJmX2E+FeP6DKzu/tIoLLF2xXLLhpFU0ihOVeu271OoGAR3L6h
ec+D8lK5cCi6qW25My64l/WHrbu2UxfuKx8mcpknpfmB47jyp/J9fjXQdPZBKArA
EylfOHPdA/aIcFDNAoUTqX5IdmTfvKY02egTGeO8FfVpPzJmiK7+j1/Ss0cfIOSu
4pcbIGpbz8atFA/4f38WCAR15mmPY4xnADm9NbRKtNwVxAeweuT3SYGqFjXh17Jt
moWa8KJtgcrvu3LGu7YFAQk4VxFQBY3MAZTGJhbPaWOc/MFZOECy95pqaaF55+tt
2JH+T0CV9/K8jHJ0WInoeKHtl35QxtdpYxTRvb6yGX04PExoCyIBFB2nLjA//+PM
49ieAdvWicAIvPFJ+a7QtjrftIMpwioWSLUkk0GBcMNxqkwPUch8UPHXtb2GWc2g
aAfPU36RLYEe8UwBM2LDgdOnBQOb8nVU7+741NrC6pOrMklMrMaNxfiwppzrrE6V
eavbh6uW3qHz/GtIJpkH9dPEMjo1FhWmAepYNamTGfGjAjHcAVy3NA0m4tm/+ICv
EcN6/V3BeYrvDqDBhZ3vPYZKJXAlhIRqHTJI34Vhh71K16UPxfI6Q34R3+D7Vwpb
z/y2tAf+dyNIhgzvVYIsat8XnZ4wiA/MbnbXo+8fwOs2jGJxpi42M5XdyhZB2gX+
yc5RueQYGrO2Re49litEkw==
`protect END_PROTECTED
