`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+V7fV1HxBs/+346wRPnHg+3haNOslfS1A4dT/YuD7XrhT7bSZPvFWhNuYerNNrqQ
4DnAUksP1/cwpUHFWcgW5cMEvRof5WEhP+dfgiUqQt51zuILuYlc4/Cv+lRoUnGj
97oXm4UOq83fTLgvq43JfRuPIatGSy3jd/11n0huUsARRnoVfPfy4XWQ2pCJawzm
vKYHEpYdZhCK9x1gudZ9fwi485K0P1lXX5Dubu3b25UWr/xF5BO8SZBYpU8t2RcV
eTVEEhkikoYDq+uMoUunzndc06iX9wvqev0NxQbWd1AjvImz6/mDyfMjazX7Ywjv
BvcEgllxet4MHf6kGuNN/XKnTUh4e9T9d0iS1gzyHCLI+AUXjcglNmRupSN4kPiO
E7hkLGAaEFDy43QVKdHlM+9U+A3TWaZU5DFbqTJLigHMfKq26ywdnj1FG2XgYp3I
MEjsDXI7GE51ixl+i/rrSwWv7dRMsth4jc5eQUgjpmhIkL+SafkB1sdChZRbETn8
PVCqhs9pRgmYRIwK29qCMpvB1H7T4ibiAOcNavX83EPMm2AODoP9S20c8wQW41KJ
sIMOcGPJF/BDSLvsBNpOmHWTqCXlqP8f/QPRTX0CgUTlDyNJfR0EVDcjPk9ovJYn
MvjH+wS6NabqE+1FHd6BkZzw9V6zGX7BaIXuHRocFoSkCr6FFpHuOIbTr8p81SYo
Ov3v0BYaOXHeyLEpyI6N/SBnYJI8PdqBgyH1iY9oAkZMb1HOS7b4PwW8eykI8cmh
dHiztBRVutpI6Rv1GGscC3JcT9K6TqbF3LEnRiPJkMszYTL1G8sseG6/qhGyOWo1
cTmtyUMJx0zXHHJ/KbGXk8RUvNKMR/nEacdAVHp+y31Nndrk4b74JDXpTT/I7h/H
8R51K9DwKlgQdf+zk3yfQOM6RMMSVV4/sRCZNc4A5AndPv6ljzepCxTuU/S6dy6S
0fzXtYAgFyQSeLknbPtNl1cBY6Gmx7TF0cP4qwJT6zfMXMt+Epn8Z+rAYhzNT7xZ
PwycoiRgidbGPZ2NpYl8eUU81fXhLYBiKjTp44Bso5byUejRWvrUL5SdjoBvRGMz
vNm5Ye13icEgYCibK0MhTtzOP9r5S85z3CPi/QSp0V8YgrdXuUtRDgVptF811fDc
oNQ+S4KEIftdupDKLfuxI8J/+rGdlM4TRiPJY7Y/Ccm0X19fE/NABzKjYcL41gij
hOkCEn52WCGItyaee4K08ufJpwQieW8J7fHe6CNodEo44aAiZJIC/XK9W05VuLw6
iTLIlfrN0K3VHICpEDcMVIIf3NLzVL8DXXLRhOymrBp/0mgAt0EwDfZ0Ao/Vak1y
2C792DQBnBYzbG/L+fkl5bPXlnzLo03vMWNsZs0xp4EDO2HvOdkIyo4GwHSVt9tt
wwud8q0BnJdCo1k1CIvO6mnU2dB6BSALNxcRxWQr1oiKbLqBjsbgxi9gUWgJ/Ihj
HK/v8MUMuC51MTytxHNP/iIDkxoK34FonbVeXUm+NZvwceLT62/M+VIDDBxuv+nn
qMs4qU7j0Ef1snDEqBIf+BQKZJQJIX2TCtkj01rL0pgKVB4NquBf5u7UcS2vV+0F
fH7XyvwAz5W8OKhORLRrm62ZCtbwg7r2K3qB7EjsiNLrirx0sTiytPyDusoNIOSe
jqgrEMyI1FLi1LNyIM7WJIM3wzQhtCIR/iq8RBM6gfY6qFrRoAhdCWfUH3G+lhdt
hShnjZq7yeoIvzyv3dfwvI2IwAHr4Q8nHMZyGlZGVaGzuzDYc68tNZyHer3B9hRZ
URBfp318Sxul2irTFrgZLw==
`protect END_PROTECTED
