`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QhHmUp+GLYO0QCwpIlR7b9yHBYVmqEfQCUMFxotqxUrDcfk2A+5ot8HcfMQYUYKv
rkq9fOFnOQ6PRDt+gJv/NdoxzBkJ+6IHgTxsaEJRt8b2Cqe+N5wVXLqOLgJELivG
J6+OQruldZEssOpjkpogrHJoI5qChzhHpCNwf3jtE8UmYbWzzI/urSMmm9U3mIQN
kKUN7OnRZqDcfD7u3iQiczB+smr3GJlAf41sPwOr04/P145K4hzs9+tAnZyeOAP+
iNqKy0WjvjCIeBd7Q/1gL9vOaeeJp5AWovgsdB8yBLEw9ghMp0OzJzuxiNx1jBjG
cd3ECRtjZXRkMabc5Cvf0fv8MHZHY+qCHPtkUh5L5HJyb4vhTwOGPAyTjAzX/TtS
awZGeBdP0jDo8TJWZE/2TGZCcbquaN2hPwrs9v2ziRDi8YrWEVTGn3zv2fg6OkN7
gNSUzfIeudmEuws3qW1A02+3jqYx49KqUrWnNywATb9uis35ylWaf7v8AEy18Q08
hsT4d3jPGulnWV3HSUQu4jTYxtJoTU4yQOpLbqgJj+/9sXSzDVcFX1FsCmyFxG9O
IpyrQ2I/ElLvbYTZDAdCB1YNof39MejABlflFdZPOe48mdGJhWKFlRZlWlfdLFD0
3ZCzM5f+Z8ct+ejbP3qWtwjuA+X6K60YybI1MClLDp2S95fg/CJ1oHtOClMLrz98
6lJTJgYe+1lGnidBLdEiVkTzOCnLI0MkEOYAi2Sdblc7BawHNXySlz3wu0FvVChv
ELdGIFPGFvifq/eLijPQstuOzYOfUssm20b+HR7T64WAupWRsVFiGxLCstaes/RH
9sTMsRSqmYASbEWKsuV+8nAPQ1VNIUMRHf24n2g1jo5B588Fj0fiZk1tkPpXCxDP
SBWKT5hbIjUSQBnZmHi9iliRGTATzKKigrq7g9shFaJgiHIPutNhxg97Az+kaCxi
O2cHcFP4wNr3bRjyaJSU14sFntWDoBq99I1IxeCXEe5IpxV16CSd1tW9jkS95LZV
NiJSL6Ny0n7QoYCBYIzasIj+APjCcs/TqA0YvKztl//dODjO9cU55YyCGDEqereJ
jc8Qt/AXCuQ6yxu1ZIo5aoAiGmhp8jpiF9nc5Gzg1K1rsEntXU3hySIN///ImScu
`protect END_PROTECTED
