`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZzCTz3Z6yvmJHzl8ulI+L48fjIN5nqM4qDlQxx9lCUqV4cjvXqfZv8IO7SVxNyeI
ujNCtK99YZTjyLunRf07DY4yJk0jOCJlmsps1qDEtAzirfmmTeTVk5EJIHtLozyr
k/1uNSxuyJnE3a+jPkfmVW6SZlE9YZDqSaplN4rxsnhMNHpjwYsq2CfV7vPxhCcM
Emq7xddwcoaDrUvleW7Nf/IhXK1RlJK7qeDpLedY+8vMl1DCnX1PsgzsC7MzxpqP
z77LJKqIJBB6agq/DOpPkjlosQDFw9sXZYwYcep8X4qQFQjpCME+KujVOulNn5Zn
mMzbSswEXijdWRMYoPHiLGgqtYavjRM5ticUzQ2M3gqSuDCAOpQdSi7yjHGp9m+L
4KThd7MhDz6TmXmfJfwK/L9ptQ9xRs0okCaaqA5sZ8gvymhXAAccgFUZpJw+lwDb
XCFBWno+a4/C/3lihJnyzzOH50fJpdyUFGXnCW0lO4Z0k0fiPG2bRXQHM59eg+75
ippm0wHHar34M+k9jiroLTzan6FT03gpJIl9qac0Pum3pS3Vk5Ajbzc1YES7yRSC
/SgEa4AVDvlKDVnfXXMcRu1NuNjD/oSrdK3uT6YUi5g/4pdC5f68AdqqLTXQgAI6
vPsD9ehIz+rBuefH2j0J+Wcx0uX2+fKFBn/3pSRkMG6+iREOhN8XaUR8V+Fcydih
`protect END_PROTECTED
