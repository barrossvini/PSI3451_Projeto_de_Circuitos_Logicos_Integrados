`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26qRlimDxTUsdXgsDP20OyE4h04yZIBOrsIahK6SSYnZZRau3xZ7R01c9YSUuKri
oS/XT3TJYiPEk7Kp+IhpUHz7Ls/a9bC2smit0lmwnyBxwzZBQg/dFVmemYF1unfq
fkgiU0UlGtAxTNz637hZiJdu3OTT2c4hklhfZwt5G0c0GA6IZAS47Y0SVqauoM4g
cLuNI4+agmrnlUMT28JPEDbhKb+beH56lIqiR0dhGo6M9sI5rjCNmLiCozRHF/8d
m5cq2IvzQhiVHYPQlhG7qNb1r4odPWVNQqUSYizCSzui92QZMWHUE5UYq4MkRmPB
06xsnvF/7WQIzTZEaOYLF/ShyktdNvXQjPojVkAokmMIfqxek6ir4bXJhIhLTTPh
uYmYBAXoRUKSy1vZa9nBGvnsWjnMKgfpRCzKQq8wxGj/nyxBel35yTRD/igDr4CH
o8W6aUsAE4xhipM5OTw83WH1QlspwhbIaszqfuZooR9Wi+NkemfsqgJkdiOUBUqz
Bqqf8UeViFhrU+3elo27sieaMIncC2BT24MOycdtELPvsLUSL+naspVfE5OccS0a
/rOnrJ4BLMOfeOlXWf3M8mG9UAnrw4BUmFShVAT2mof9UD9/lk4ynVF2ZumwCd/V
ICNz4JuE/+3Zl6UtNc7LsXbbNxWKy5R0DYlDvRho98xvl4jlQ2XzmXCCrEUEiU0H
LCApSwZPaWFBhI2fdFquo79lIgX0ICcdy0SywciFAts+g5UzG65e8o3DtmcwGCpz
0+FlJFfjtqNg970fZpRvYkXxSInInHs9vbuNunr7XHGXKXBSfzpThcViXR7GwgIA
HnwaAoSTp8AQqzQa+btDRu6KFaZGpe4Vm6MNu5XgAdYnn/gaLoLW8Pp8F64Wznhs
1F+suHCVyiCy7plEwKTr9oGzHnIt+ddSwfOhonoTE/Q46EyDAahicyjQDax5FS40
X12qFoVicGE/J93lkPyQwdU8ZaNbyvTrIrc/xrefv9KwHZG7oCmvZPp38VqBcV95
4mfdwv9Yqj57iEMNjvs5ymMJJzO1JbTUbEDwLzh6vNdPr4MHZZ5Y83s/2h5I9npF
nNz8Bq+GsD6/tK2QDaddTZrWlBP/dcFpHiCBQn2En2o9wnfEHJ5cwriNxHVoan2I
9/50XXJ+7psFDuffiE6OhXsstIaSfOzcSvn9zQewCgNE56Q+QkJx3rVU8dbPbDt4
MkDZTxb1pu/urabaXnjKB24WhGt4BS3f1fFXJf506e6hL8g6PexjKnoNk/xJw8sz
+gsK8ML7wqmPW9/neVf6ldlvEN7yMCFCw3P/dkiZVAYfQGgQBlepTj4QpbxyOfbG
Ly1eix7ZKCXUwJdWsqamCM0Rw6Z3jq9MJ5CFBUUV12DRXsc4/0sRZCFVGzmgJ6a+
CcAIkYqjrYTmn8En1aKVoTcdGl0f+MRASVJb/nK0dfbTz9m52olngRUTMnlXYUl4
ibpMBAszOcxAF3cTlFRxrnpsHHuWyQfUBjCawmGG5K8tJQf1mz6JAdXtogVpgYoW
hRp1am96pF+mhGdzpgBcQ1T3H6O+8vUBfs67wDBBMtClSZOtzPUdv1ZQuz1NmMcG
I+aPKh9J4qIHK/fGYpnFoOIhYSQ3HghnSh9AP/XIVxEhxOcw6GUab3CO5ViKGUrs
rMQADAB4POh5RyV1iSxlzUCs+J/irJn60R38olbTF7SKIPCGkzw6v2wTUq69skGD
NhBOpr71igTDCKCQ9eRJwAMxVyaLT0SE55eOC7nQjAvH8wq05NpU2Ls1Ka+liJSU
vuQkMAPFw6GH13HWtby6ZbWo+MdEraFIhZCAGa5gVEXI9XSKszKe568jeub14AtU
XzTB0wOhJ4UBNV5DVTmZ76/sZBrx7VvRgk7g7GI6Y5/zGD6zD+IHU22qOxWc7KJu
G3zXNcEjtF2iviQJo5RggIhYcyNaLBxyvGg0hKYMyn7LZpq513/AfpfSYI91XLrg
M8U9732QkV0RKdJg3N8MfaMhAR1sMlhHwFo4V71o90O2E/b8RILRj6NlHWr7y5Vt
9XhDXK/Fg1WlAjgDezc+2qzwBfR6znkPcm6lA/OFUrTf9HmBqDfblcB9Jg6EDaXV
5RYsx/S+awiUq2W0a/Egtr0SsdR5HcmLD1zkNGftx/ZibRtU/3HzjxfILtB1cVzU
uL+6oNcAyIwjup0kH0I0VzFTkGZav9lLer44gQZ+Nsy5WsFws19KUD2T/WfAaxQM
A9DDjhsX76T79vID+88D1GZJziNj+M8GdmPPmNbacQSAs/w49/l/Svf6qOUBIbBY
mP5+I68nGK71zox0O1+gYaLccKsgN2gbXezHQsEqIRUdMHf/xKtxG1WM0TW3IvSo
cPyIt92oPuQwXpwNZOxMLB19hnbbfLuElOrJZblaffx07KmjbPXg+VxIVwinZhel
nxc5q49xyDfQwim1CzfpZspflbD+JtilrdqP8aF2Zh5JixjKOF48RIQklyAiOROL
VAkz1k8XBhhLJZzd2gEEF/lmijZjRhCykaudV8qRQb5QP9OZ6Iv4uCRH+of/bBhZ
0J//9rlP4FGlPivk6xg3bilt3AKx8zSLVjH83ukIwa8fbNUSl7HJG6T7bVNBNgN/
EFPizA4pWLc3Ark1EY+TQx0F2vip3m/7Fdm7tJZGz4qmjjU5zCWYipo7va4z0m/d
GNsYFue5elvIjkTTk/bLY9RSyKnjHDqQdQd1OyFJMTrfIhA5r+FWHprVlTsjMZRr
7n2l3yNsZizDgB1u8H0vELr909+wGxcyPGUpujPq06J5uJXml7NpSHczic4letui
6JHDQegJ9OEo539WxinXZIBenqAOefUVLQQ/0G7wW++Tz8dmDbfTlVCBmYtR140x
ianwdCs6r8bzruicuQ1JsmW58GK03bj9fFQbpgfMmt1umLI5AemvZPGV4IrPeQQW
+WE4u/8He+4YZ8XW0Ogt1txA742+lvImgkZRWOMA/H/vK8ewNz3Wb7/vbQdrbAhP
fus6kvMkOAU+gdvxKJJq224wRfpmVcb+Bz0iPI+BEFOUojiJGyV98AK7NQLrkYLg
0I/MYGwIoadT5R2LZhfh5kIUeMW1j7756aRfdl8fiEKtGBcgyyl16lWHpx84huJG
CQzo9ReqGHRgJzZ5OcvQo07rPoBcjCaFR+aNmMoYpSgm+BDSMnX3b2JB6dJ3dAsj
tMK6cCCsJe0OvXBfklQm8AYZSm4qYoHwJ84zWO9QXl13crh5cIqq2vXkLkmiHYPy
yjvVkJGLaksGkudGscQtd4PBjO0o98RDPaHwzSJwESJNRaOpIRapapTHV8yeYGdE
6f+NkLVYKES6I8uRDle380a51/mSZMvHBkdYAiejn6qifPV08s5vMG4y7gRHBZ5Q
IUu+21m+FP6AUvqjv4r3Wjs+5rIYnh0qLLu4V79my7Lbgocd404xNPBboPSR455j
XxTMeSGUykFZ807WGTAIeL4+cpXIe02vdwaraYgXjL/LL4sOjyvfy0XnbtkspuJX
/Q4C9wlF166vhwk14oLcfs4iCMJnF6IF1j+L8QsEKVJyorTgtHg8dt3V+NlPL8TH
eD2jVbD8GPH8Wc5Ia36HttO/RjP+XXJ0YSY600slXumKt1uUmuJd/E8EBopCXPId
m7UpKDTiQH+NYbF6uzH4/MgyKdN0cGFjYA7WmsHXPQV7x/5Qm3K77xgT7xsQmgpw
dz3nqno/6dZRuMj4MiHrqdT9N3LT+B8xh9s1etvPxuS0295j/G48Yx1Wxj8PNBcn
fQf2RNJr4dhP9TmiC4C6TCbc/gegflueYzpZQ4N6pojdCMhtj0WkIO0UmtHWr+64
Il1sixhfZAzctj8bisvLpoermXFX+NNhEt1eMCMuO0LLbQf//OJursFvwp6LceEd
5zUAkO093DkCXzVY8fnbIjuNuE/LvCvBr3YhpNBhF1oVUPEh9wXWfftOhEsoK/VO
r2nU8do/OX3TomCm3tB0/4Reh+/UN8LProWxz/rUBlnDy5cjM63/oUn+2F6j1dYO
DXUbICWEHGEiGqVRVSuUpJaYCfki8A3t2sNe1EUZwyk8uf7bWpJvrNeU2AKhKiYd
ky1OZ+ailm+5wetnK4NxC/Cu1cXgE8xwmu4cu0rQoG3SneRA3++X5RSa7pQOgCzm
roPm10W9Ot3K0QI818zjtptsJvjMlw7N7FMI1CLE/GNdpkWpglxFJHv6yAfikALA
2NbDMuobxmHqqm1FP7ePioZj3+XfC6Bkxr1PwJnwUlH+AAE0oecuLi8v60MV3R1S
nwrQjNXtAaQqAUims6pFPbuMw6RWVMTDFnVaZNvlnamiXdGk2SnA+WE5n+NVr7Un
gexRqGiAi6ZzOklDhd+SRxIIUZQh4l84ANC4b9lv3/S2BVR0FPJCxeV36UFSVMGE
Kme4g7cxCtK8bzPMVHQcOVS/vdSovVVDFMQxQhdICMnV3KYIpQO/7sC/oWKn85Bd
/cSSCyrmyhYEEvohefvZml8MQJgu8EByEp1AFTZ4/ZWFD+hhK9mOAZDU2hk0eh1l
rXHvdJuuQvC6p6ZjC+faWA==
`protect END_PROTECTED
