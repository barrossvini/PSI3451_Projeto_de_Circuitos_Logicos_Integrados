`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3LNZPdC3IOBB9huyogGNuMhE7NJ8AkbH1REimbrpBH9jhE6p7anCZ9qu5YQcJxT6
Puw+/63Ys366+ft9MEeE5kUuECfzh/iVzXm6YxGXSr4DNvD5hSxgrFz+7KzuonTU
cBFYxHUI5lgCcdJPRSCx3UHsOWRXhiIqOA7kcRb0Zfnr2nR947XlsaUl3yMEISB3
MR5iD3J9hAnNoJh98TbXgNu7nosqD8OVUkLBAumg2Lv/pJ8mQzCiuBQNzrRbU+0U
tDguNV1ge1qy8gep1/wgytjLJOkGdVt7vP387qVxDE2r8qxX0bRpP6g54adNUlyf
vSo/WHV3RRKttHEEovZShoFpx8AKX6I9ZPlFTh0Y1JDXNd30M4ACNPVfcEVtlM6i
xe3MrwW+V35QPEpKn2pc6rT86wkKi4LOi/dankdHwf6zuDZvhcr9dn32vZ69+g/3
zkVPM00Gzm6NnXb6QEqoFIvKYXd0GCXZc4FVGWB2fL2Y/k0JXN7PegcpFl5OcPgk
zeppDV5RV8UVYILjGGkZEa6ebW44LGRCivxvyVnqY3ioChxWPj6MRCktPCVdLDBU
oalV/YMW3XjqL4OXr8VwUvJ/Oc1PDAfLcx3sNGMPcxowUmGk7IIMTh6rf2kvZdGA
LMTyBS1QgB/gvNXI5gE3mHM8EnC21VXrDpqKq4z2kfxaeQVbSOFVoLaHHnIlo5bI
0npgjQQ5HzMqYkkQnR1lroFmHdr8Xh8AGSRYX35aeUgAaT08f1vz156neI2SDW1j
qkl5jfhNQlEFrDs7Ceo4Irxd4o3rTV/CvLNy1NQl/03t2myztAN4PhA0fYlf36uL
XSsGHdi4d8YZJhmcTWW1jEmA4je93zT9flIxk5JcWbC3yBXYC54HipCYJna3IsMi
47j8gqv7cixYJdSxmdg5OJCa3trvqeKVLuW3NkxaE7cduwPqEcaUhPc0A/aQW5Md
Y2ThQ3YdkwB2VduxBAczAy4fTV8c2JHCsR4PQ7ywCJpq+qdglh+XpQdKpXE6jlRR
L3zKMFRR8cLTTzrtRf7p847zuXoNbOAY6kFl6nZmyyyUJ+GlOgvqX6pfaVfgXrJd
P6TCsyZY0jjtKJGY5CvUkRdrWOZeKjBzYC8r30uupZ6ENTU44Bdmqit+IkzdzNgt
w0KKoPYqhyFptZzYBEh7/PE2RYVXTHZWjWNwx+0J4i0THVrW00bgHgPTLXDlURdX
DslUWwqEzfWhAYFLr7KMJSAiP/Htf7dBgnqw/Av2jO47BMKIymfhGvnfBs4HroO/
PpF4DWieS1i3qWNr4YJBusYIAkz8Uv0NPvbzZSKeZdY+zF/4U5OHg8lfcDW4vuGq
jw5cHht5ZqBgQ+W/mjTdHwAjUPwR9z9niR8EekaJb+92uhB3Svrnzl9abDHV1xyL
IMgTIx2uNSFIHh6DwZC5+ZrlHR4/tOS8ffYCctFJN6B5buudVFJvQkCck525XvOZ
58UCa/H4WiA9JHCYmAaw7bAPpQ/bNmTTu3WQDraaejGy4qp3vUB5r5rkK8zow7GE
EYmQm4eip7ZySw/gOJylOoVReKFWedsPWZpLByrY6kQibsyXqyGMvxM9oauv+Hw4
rWGQXqCL2jabWQDMu46TmoMfxlX0RqPD1dB40vYKRJWraMBN8rXvlBNKnuuUmNm4
8EmpWCR0qSJBTqDtarQsI8pJWNLf8UIbXOjOL8FjM3uyi2DU2xOB7pR+rrIA07nb
QVF9/8Cu816S7Z5q8wphOPjWRrLsx2ajOnZF21dZv8M0xolr9za6UFu6wusUVnVc
0yum9DUih4/GB3p8yIuQgyikDmpc4yOHKHQ1uDQkdn6rpeOkLIl+6Kz0UgKmSwhA
wFDlGjPTJOgTKlgeCSRu76lTj2ay2stS/AR8/f8mqcfrf3KR1fRcqMRGhbbiK524
LPDwDEFADtOeSUHqfK1yfOabVfIBMlS6Qd9g9KV1EMmMPj1OF/77l3eylxKXrU1I
+gkQrIOBC4Lwy7C97QIa/kII4TypPIJUf5d7NLRD2bioGZVF5msfHZzTLEX7VjyU
BMdPscMQ5Cmu3waMYSeDw1w/S6SqyvFcsrtT4gJUwpS8T1MgqsD0yXxtONbmszwF
pODxTKaFmlhLSVH1K4x+ukd7NT0E5pM57yW4DA5rrVU+tpJZqp+CwNjfIWEvrNy2
yLb5b8NSpRkwr200aWkjE/f+ZIDEEggawSMBoE4QVKktrqWRQiTta1Akx9NpI9tO
hhHWtgAAAKI2Hvzda168q6zaMM6AKJ1JB/00JUq5bMPi77H6UmsGovILhEEnEvJB
lYQllywBhNbQEa6Ze4FIa0h/k0cItHMXmi/pFFWMnTJldlUcaEg2hg91wV+xOluS
50sgLN8xI97lGZ4H0t31CQV6/KLVIPdfSGRJz4O+70lyi5N0GV5H81cdhbUM6463
1etLlpLUL54oPusTS67X5iTCJicdyq/mc1ZMllrZ+OsQW6KfdVi2PNbBd65dPe2+
CqxACY67BrQSP8ZuWPLdIjQzjAdykh/4FAAMuX4tNfURnfKe1V+VVwtFzRgNNaOi
kyepdjixqIq1LtIVPgBkboHlLS9lhtmy1niSxV6UJdsRWlEGsL/4y2ivZmXh60ev
6aRH+nhd4e9AELTLn5ZE6JsZxCyXJPziMi1Q9jpnEx8JdZ6DKNJDF3q0jt+z+QM8
vk59N5RfbAbnjLMcwZaHfTPxlBgze2Y/F0sOaRXBRgc87bI9pqI5bEw59115vIvn
dshp2jLiFbTXiUmUQJyAO6fmA/81AtUPvqYAD0rNqTlJQX9oAbw5MTIMbS86EqL4
yJzBG9uZHHSRjjK7OcGb/JPgNjKfPC26X0UMTZN8MqS6q7Kpev22mf8AHXyPVqKI
dbbz3AXsSlnBX+V1O+PPqBOWewfj2wLQ4ZN3CgIG8xUrT1HiS9G7HRB5rsRAe6UL
/fMMF9Ot28ZX1ngPNC4HuPMBMRQU8mZs8AYwn81v9qRkN/+oEsXwvh/Gsl57aJUm
kfx9QaFxHHL3/l3rbf2YyuSwltEtaudTCQKtSwv2EihwDu7QELOBGyhw95WzSiyB
sdZXKd+E3sn7WSTrLlRQC0c26deoQJDxv1gubk/EDIAAKIcqOIjfUUFAc2UUmxCh
DachUwVeWWjMG0OfxNrbq4fstpMGkydg5A6AmoMnaLJ0LdqKUgKFM4idb9Pfa3Dl
zucDWp/0DRfQGGN6BBaq0VV7/PWjOhWxzlKu1AYUpCg6JmT8cYeRnnsmwShIKktg
TIi5sX/hfk5Ai4KonTqBURpTT8A6Nr9nPMfsehhn713mbMEjUbC0jgYdFZixmNPh
Ad2OT9KtCms11bEz9YImethRPjQCuQjbCfp56U3k7PYwG2af8OffDxNfcGUMatNo
smFi1DK4LmsTuLgALj9myYD4rCzipm9EzpkYu62Qk4L6gKaqhys+a9nCJRT2jGDR
3HprDL5k6Smqh0rsZqnxV3lQ5U2FOKohUHQKgjIoxFApuTOd+Z+X+lNSu2xrt5T5
qeI3cXxCCvIJ/M56E64KfjIq4Az0b+RM2++Lh8jA6Udz6a2vH1wgrm1Qg14j6HvO
k0n+fms34CtEcOddTDBa/mEZ/UQ1r/TREBG++/fJpI976HbUzy2IP73Rd1FSnVEk
SsZMLGTG7HxvkwnJ2DTyw768tQDUrE/YK/dpFiLHCqF9c+D5r6Nds1Tju0qazj2U
TdmVF8aJKFYsHbmDmv5/mIxmobKJDP6Y73OPmKV7jaxmJeznt3nDGNDvzPW2bRf8
MBTpW1qSKcflDZiYH8ntmGTfBDs1/sZeUt3YeRT+nsW5LXQ4ADs1T1ySZuHuCX6F
aBGZxQM/MUlSpZo1kun+IN1kfmP6bbrqaPDpcgjyRowIYBNr170804A0+YWL2R4r
AuLbH3rAeUg3zCCLLbNdF83fyPbqJzamljMAoiKc5vJcnknIbYpgrHk/iad3Xz/o
OZ5tAYvwgns/PkzptTPPDlSzAMSGB5ofFP7T564yaWTnBp1/NupRb3AQAaWLwMsq
v6UtwUiDR4DRnUvcKSmEYTpGDA/Ye9zd2CN+V5FwEiIbMOShwF+R43K6efbHEFcO
uNbdnWcKITNyY2jDBorAk8lOLOl6cZxK/EyYyhkeBrIFSJcUffOHrJ6pkuke4mJF
OGifWIJO2QlTfPfl0Tarf9NqpwXqJQpJ8KoCBNizqJYROm6Y7KrlDFMbSza1zUhR
fe4C95ZA1D/841R0Lr1xYBcdqBFaG4qThNXFEBiH/CVGhwTI/ouPjweazFPfE4Pe
uH6b7OitnNqtecnaT+jH+r9QEiE63AJcgIkJmB4WccrRmfJsbPYyJZfh/VCqQBZi
3ksG+1sAu1rm5W68aePNz6fDj9yEOot/ilfwdWN/tRYUAVeAxL2FSTH3f3+2Q8HQ
6M43s2KpUoHIvpVjhoJMyz3stPHIfmtm6/j+tV2tttMmMlpZg6nSW19L+Vp5JbkK
L0WneETCqqNP3xqBoHnVwGcQ+elSQyIg7u1GF+ew0jM32nHvQRgBr7FY60d1lZp3
Caobw3GKhqWSMMFD+0UCzGU9mt54pZhb5yEjw2oBFzzjQ+Fa3EVVOwHgdjsoxAX4
tqRD0kjkHfdHV0CRrp6Ug6oXJhY48Q42tVxkt1VaZMPkczxk51h1F0CXqIO2AjIC
wbsoGuzjZarHnsPTCz9t00NKW7oR/ILiWIlrquLUivnzlvfzwrPYU2w+KlPlhplb
Z7LxVOJ55L7jyUceK11PbescQsLtlWcuVYBaTYWsVsnusPdBV0hQHtXjcPjb2jEx
5ebagUTz6EWk0JxT73WwxU3zhN8scr5Vj4/E/xfW81LLUqJKBfVt4a6gdP45UQSh
gHgXL24EzixWy+kk7kKg58TFn/NvJrESYP1S3TxaNXxaE9iXeGmnpWeO+V9qeGsr
sAHotuNZEtleRdfQUokkGn/1LiWqpU7stpEatz+QPKManvHx1bFYpLCqO5av1rx6
0DEyz3gMRMUytAxIxc9R6x+WgDPW/XJZ9BUczf0I3dP7usJ/G0Q28/+O46bz5INf
0ottMJx0bm+TdDlMCdqRaGe+j0QrTNbRu223ojpEncCVmtfAKlFD+OWJMg6WFcEI
MQnKqTKh01SntS3lyXAJGbiUt3XyEm+rGJ+ypnZtwCqtTiGgoiO0wWvvle3kEvf7
SM1UjVd+Wm0Ct55abEyRMdA6BbZlx2kWcD50JynNyI+/WsBp6Xl/jn1IsY+vANd4
dSU8Xo1mFPXvXF6Ftv5WS8U+CnBKF5xl34kAtsZ0dAsAtrsgBKpZQh9QlcoZZ5KT
MwIHwFMyMYWsceUNmxtN66s+hoazQ4TZsVCkYM6nsuEIjbilYV3FJBBdQJ3qjCaA
3YyVkTOEwWBWYjgXiyXOmsDYpXlCPel8vgKYsNszy/4QBGO2Io8SRyuK6EyyuKiZ
MJ/DbjQrmPyFdcJzD9nuEy3JqiNpUJW4nmT8tenMIMgRenpdzQ297jGV/kbtH4Iu
pLuxGj9d25sg5fbFtFFaGGrj7socKFFNSrNv4pPK4rbBBmaYRK6zBLseNHCsicfH
GS6Ey6xM9K1c6nIqQxDrxVVmIm9z52kQbc7u+Rsw04Wu2Fm+3+70PXiZtjMIh39U
TqkuF1SQw+PCqQ94XQJY//xxNaU2RjWuckQBMpdH36x4GsNO3GAsY0ttZmcq7HRT
cQM5JNSXEaTLOW+19ER319qv20kyqgT/F35fcFtMe9qSG4EQ3MkrovL/75CjSw3B
L01uxF3K2500uzWCkbT5MgVnCXssgrzHLnXVvMQDB40XJqznQr92etTPgjIuJRC5
fzAe5YSa737TVQNa4b0tBawISZLyCBw+2O1J+OoQlGE=
`protect END_PROTECTED
