`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cdsROmctGiVb9kbdtmDwXWILxcifgJ2SKfUGlJqW31P9aQK3eNrWJMXwMFHR2ymB
yG31Yw457oJOoTGsDQCT85uNMaJY/qUCuuGU7zqoJ60SSAVCmcMGpMiVNrf12Yb1
6XZ3G+gNsvgys2L/EJeKYEsEq87VsJ8rDoL5Cw/V8oCB/ZC0L0kh/vAdpqitjSrf
an/Rcr+H4RYkTZV9kLM/XuV1eyK42+nU9onCXD9fjTePXVkC+k1eZHfMBWlv1egk
Bgwml1xUH2D4I5HVv3XmQe0KkCl7ggBKNUD0A9RcMwB/Lf+68ODneFVtBm5QzfMb
gLn8zhUExFv46SB0xYktioN9cPAGhB/cROCtt6AX1RgDeyZniCb9bqRIDRc78RSz
H5/5s26QckwZSQVxE1NL1hiPL61Tmdqmttele6yATAZQmmjxgb0Pbu16737SwrdY
Z7AHjjPIpPks2kF2g5QTmEysphlXEDJr5eZCB/G7uGX+tzEwEKBSoNOnjRJ1D4r4
x9esXPxgL1c64h7/pJLq+rIIX9nzPQojdiSJipRZD5r9YaqT520mvxIkzRaAI6Kz
nB3p/YiSSg8AriWqX8l+lxYw5MeVcsNT9Au1IqbsreICPPCRmlaHNqhf7r8m2uNC
70aC7Pm1Jsv+ZP0fn10mG4g1IdfDIXfG+MQTPaBuabYDl6G6UPjWoKqSi15tLuDv
dqJ/7IiKIiOM0lxxoH4RXM33yEDpyAi3if8q/EhIR1xQuqj9EEmh+4qsNah8Pj/D
9HlusDicLyO5W6qiIPGgTWXpH6fyQNhYYi+/vo2Z8Sf6UydxjD28B3wg3GsSb3xr
lELSjmbNORgO71wWutPQju5IvDXrEYhMkRNAmAbjSr4YRgzio3J+ngADglPmSEfh
l6pQsPhZuXF2lwT2SjOj54Oq18sqm5AeFpxFJH1ZuGK76gDHrs3QZDXJ1GUh1TsS
ovwlRYhcv2so82HidRg+M/RYvgh4clvo9IxWTQLgGBPNkb4h+L5e8kWwXVUUtpRQ
l3d8pcVwTRxFKGO1DBjVeXByf+GIuvnKJL/1eA9XhlyEMghTUpuZS6SFfhW9OI/r
Pe4+Y6STLGuCHA2YgDPgeUMTLXkotiHCnkz7a1+eaRtz98MICD/L2qD36VXBMoHp
oxDBY3WzrR9NbI9MQQN7p6cWXtRzto0t8RP+bfPDtfcNSFwfuasjbaCMYl3Z6rTQ
7RfOkYMWKj/OYrxLZeLXZDBMPfp8jOfqxyPkC7bzx2AqxXy6HZLu5yEMLssQk+cK
+VkvOQBnEGpgI8dDlXrvPhafjmoziNjGeaGkPVdBtCz4CjXXN2mE8ad1O/bAqhro
cHGvy4Dw8FSHa+QRIbY/44QNPFlNod7STI6eil8/rltU+dLy7c29n1swrMm+aLcx
MDNHIm+Z9vQOxXdWSsbKd0aAy3yuvSK1QcB32iSpcT5Am8a/5b4EQrSd1sPd5V+U
3fRFvEiwwF84wsjFigL5t5gFmS1NGJaB/WlAEdmlYE3bPgmmsGw8hb2rHI56UwBK
whFqDEksoujHaWTLtL1AhIaHAC/jcml3fpzEG+fTxYmUAJA36mieOznmxH7PdCIK
GcQyVchRPrZxWRemfNdri2c+GBYCO9B8Dvp8EFVL4r52Nm3+rOBMdcsKpBpPqOmV
/wxZ/XEALgrRVQeQhtJMv2lSObRdeEI8LcdNXlcJa+U2N4e4NLPFwP4/m1i9j7ol
Gpzyl3vhLLWonKe0SGmeqTut0chpO0mgPB2CsS2ew7zm6ZiGZB6bXJeiUvghn6w/
ZJDpHTEqX9HXmGl20+Eh1zWojuR0DOwABhhSd9bQj8Pq54D23jZbkIfmIW3bvmmG
/nHlylU1jdE6b562+gbJXBlAQGPouAJ9F0OkjckHcrYnCHgCWl6w9JAY328mwf5x
4r4w01ZvtbSAjhVoUH5wVh83RWgWmrknA8rBtIpDdoaPLYkCEIXJVCrRgaOURtO1
AA+4PpqX0baLIrGU2z6WOqTlCE00zcalDDUE/MFUPGUYmIpzZvwjUtO5q/xvndty
SYTWDeQjsIQxCHs9lai0HSYSLbE7vT81z9lpeVL0FavcHUNkHWzknfKHseFuRC2X
vJXeoOYGvCVvlHcncwM/V7CWmA09FDbGsncC5oUY0HWoYvYUk14UGaBD6X9xmXW8
WdZqO13hO3vCGKHH/D8F0p4wJoFprzlDQviOkPEjSaDLy7ql06anhLlM1rV1a96U
ljkip4aanmMyAod6KqyBAb+NzEioOMRnXuDT76D4C1dArkEurO6Gc17QOPt+JWWY
0wXomuSy8nd+KX3QRXULlRxnEdjgVprrsBM2IjI+OTuCbQ02Mao+roGGgECjfsA8
V4NBmKhXRBAyPN9oLQ90cN3oOAud7FavpRsHaUJ0vPIUuV/hID8arb5MzPpxKcgW
nRBR0LOaQrDSoZnEc+Sjm37TH08pBsr/1oh1zIdKb3SKaWTYKTrMr/Ual0PBngF2
nOh53rAxzVC9PKWPUyWMeoQeWx2HOy2/RrKf2vXr4turs9kpBuBxpSoDzjJ6gLlz
FPwdR/9olvF1tzOV/ESHAMeU65Dzg6zXlEldhj6hPxjJ/KT9ZSzpG0Crq2m7cHRu
0U6K/iLJAlXbemBbvOMhZgB/uvL8+zcylmX+k5kKkmoYsq2Xwef7Dd9u9DhMD2eQ
OME+RnwecXu03essWKamV/ZcvCaQCr0+4xJUyQhK7nzReBp0Hci1jSP08sv1rvqk
yaNt6yhMoL2QV6g0vGOkwn5dmdXZ1hI+/Vq+qqEllLTzgzqHBIFqWjJVeg5aR6sT
SgpNwQKx1WLyrY8j6R5sHSVUHvE5R2kicyY/wphulXoR1g7b8+M60ow5nDWikBs3
OlSjGHiUPaxOOdrHPLpCG4alYOcRAhwpBAm52jVriu3S4rQ2wvj3zT9w1jNJ7Qo6
renJYPj40uwDcwrUnT3GzXecRDcR0PFdZ4v8//KUv5xIRnPser7po3J8IxII7C64
/frCv86bSyKKbAXqZr/nlN83xNuwnQvKYRM5KmU76O07RmiH9ZN4ljDkpwwX4FdO
MxG0gamBCRiHlR9sX4LvfJK6tN8MZjZMXz0u/QDuoCqlIUo3Ex540OjbLgdSkueR
u5GCkCpCyvFgYP2XjqEKLJF6/nynCL0GPUWOFCbS/3g17xJHdSph9HV4ER3Ft4o+
90KdrrtBWYOHP/T4XWK0/tlRacB8LHOycnztLaLd6htxOkJXAVNQXF6fuEagdaMH
n7dSHAUIPSW7AbIWJd3Es75YbvjfQovTKFDmH5d+U60SAodw0O06IYqgRU6JKBCD
HHsownLe0topBLb4WtUHGWXQCNuFmQSvNCRNKR07DAj6C9HhL6k1pPFMi0MgGsjR
oQWculzbYBdX/Q/EhFrdABmJmMXRm8Vv/HqOzSHWrvegxtx4yUfhJ3Es98S1UuCJ
dQ45KKbZXc34PaIHD6EIXtTIdY802gnTI3fOVL9qfoJFXvi4MnFeJanApVrKxBYb
j0pSR35F2/iJokn5eQuxCK3BRrHvRshV+qczDsGfyVgr4r2sDJpwYaSBtvLgZCRv
pLxisUZnCHP2dG2ZZnhYPDebLLpqLKaiRzfqP6nVN6HQkIfBzhnsPR5Uz33DZtz7
G+2bULNO/EqYvWj/bLikBNvkYUM+AL21o/J7OcWJZE0cWCPMnH3We9aR8hscSkXf
ZCI55GVXVR9ty6CYq3KnQJwb1Z6unxTZ4utpWNjAEJrfJMfVL+mHx2s9fMsGn25H
+sUpTPqEX48k5ejp3IDrdG2hfPEp1feo0tI0cUwRj8TQRTxZddPQGRYanWf7K8qc
fwvpKNtizFPxBN6UveQnjIOJqHxFCkzeEUENFjgnE2YDOwGIsow6FjMLBRDd6zjJ
DfxmNDr0g1VOfRDvo53mxEBCQItKMgS0m76RtyyYFWoIIUqtIgZ+X3eClQb/ctMY
e80Eh+Af0//FEn7Dgi+tCU8LGh4IcGGQNftpW8PTVK7FJx064YnDA+QVWicrSxkV
o9nPeCYEE2401Pbj7wctPdLMT/kDVeCfaGa9nbR8vXAFAMUzzoPdK30okqePxMoH
rZzJQRkFwypQHeTvTI7bML7D3YqlFY5AvhTOP18ebP3jP86l0MI1F92Nh/ZL3fLa
+R2BQVq0nqvgBIY8DvPAvh85HgX6SYs95F5ho7BnH0DYi/5JmezFjmf/0niZ6+Xf
OY2RNwxb6UW0JdcVWZeF7s+j8zbC8GjVL9voJUWnbinHrmPEJmX+z09CYwiE6zhp
pWZ54yFqw17ovL02qtPLcj17M/dfW4tqdbXvvt4Ae0Zub3L7AJZQhoZXkIpMiIWn
c6VjFnpkCxsIv0tdFruVSDkXXoRAJ7/nawULHE8r98wCnlyBc5dY6RKQToBrDvsq
VVdXsWQwUG0tBzDddFj2+blBge/utKhWxXmY7EiaZuOcXIuf3LFRF1yPQtPDrxFg
sU3LOE2UhAYAQUzyujWQkU+8yXbFHGN2RRZM1vVUeo/TBLU6lEuVg4c19p9EUaBa
ZOQlZ+pDzS7Edau791vJu76pmiHUC0fY4mp7l0FiM4iJoDGLlGN0uiMxSx0NzzGd
nmJeyrtaW3v1pNI2l2f8VK0itjWlbJpPlqQQ2Vx5D2hohVaKm0IxLkm1apyDvwAY
CA47+EW+bCYjxSOK0aGQAIlI3ObdBAiI8K574r30gNj8MzpWzsHJqCVkfPayJTAC
XBPDSo0B4Jkjm6SFyiEtr7UUO3u8gpCg//RBpkobu2VUncdvPvEVEGcQygLorEZx
VpjsTd83lr4tS/RodcqjzzYmMTzo2bzPKXLsVVvFND/dIeEwwtsjlAqLQaJyiGrE
deT6cGTp1IEwqqIoNvNTFfqo3B9bMNLb+UPPSn1KRPrysgryuD9Tlys0mBKo/3OZ
DFH3FiYTJhwQjsBkKuBQF/R8JfrFK+6imZo1k9IPnlk=
`protect END_PROTECTED
