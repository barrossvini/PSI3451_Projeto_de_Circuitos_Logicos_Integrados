`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4eHm7Av5vMOmwTZ0YMaZCikGLQjGJPsNCBURse/xtnmmzCZYhRWxV/JP2X77WR/N
7BB1fbcLv1O5O8EUuT6dfqiHEZnp+fCgc9auENO/RZ4vgC3/qg+gm8GFJWC1/Dx3
dhXvVUX3ELW5CLWCX7hnx1J6NZOgWW5jhhLcGdiPI9WjkoYRBa8p/rIOD79ueaZg
3TxAaK0+kfJoCfiaM4CmG6Ui7WVWBpfP7V6xYHQIE5/HO234+pwR4cSlWg5jDh68
jPIZUZCwJzIEtR6F/Uphyd3lFwq8McnKcxLK1l+2LEUgO3sU0xkJPR3oLG1y4TTE
5z6NM2qBsJoNe9B4GdFG2SE5/7Z6+as3TbN/6J/kiahyJnWy5Z+qILyCyg8B8A1U
Ky1dQCPjyifUHwiEjAy9jS8dSF+MWMRJ6VarDDXNJilzTKoEJ5ecVzQyr4hJ/WRl
X0ivstN9iLsaAoMLYMWADZJQWBJKQ0vJojT0Au8PT+8xFyYjrCQU6ZbhLqaf4OQ9
wVmdMywmK16Ng4f7mteLS/Xe9Dbc7kHIEC0l941jHcnW0bMgn3JTkIDy6xg9wTfT
lhYOJhOrLvgh2Wehj2O0yUgY22jvfqGJ8Hcja2Y3Nfk5HFq/3ZYUXrn9hSQD/GUr
RoGkVV8MZPhz/zNvuVun0zogMpCp7nhdK8P+HpVNuF1Ng1hhUyHDmjyHk6cB0Aip
8z2DUD3LzMmA8qDEOLBpdmWCnS7CEHiqpvRQu7k9jfTwUD/hkWne9mYpQJswjL0u
CkNiViWh3qO852eoDpNjCR63+EAVmj59bVVqOEknxYjBLNxquNBS6oCEGwK6ljaR
gP/Kg0DiaQowodvdW/zAhZQDlRbiVjlYqRFUZhzI339ai8BJVcIzUFrLj2s0k/pD
iMUCvGopqwfKIp1bZ1nQuogr0ToOGTmPLhQ8LmmbptLjc9q8kpU7DuCa3nrOjfAF
Fluy0yRh/ZdbgF4hM4BL+nNetYY6UERYfiLq2CfbFJ+vGyAwQRdGWJD8dqrhEhfy
ThHoMt+uKr0XXQI55n0Ndv2DdtRwCoLXsR4pQ9g5P2/vmjnR3u63PBqdeeLad4A/
cCKy/9ukOPjHnywE9WndFhmadg5o056lKiXTru/T/wfNmxoCHMmiDVLkEvQMETGP
+w6/9iJnjqJJbjwS3CKKTOfzF4YoBw7Y5C8lR77HmrZgQJreASvN5D5V8gtcX9fH
s0yp130W8o735vi03V+Ur3pw0Kl/t/flYRZpDPQ17we54gA/ZQyQoYU1urclSGur
nZs9yICaUUtvGOfY4X5qsGnZGMmJI9i25K7LSwYp0Mlp0vwr856YYRC+niKeX7E+
arxCIiB76gkiGx6WCA0+xTZnNTWXwTLu+lzIvbrYkr2NCojnbMJIwm13m/E/DdH1
PW+82w4FjLeXLWrrWyw9+vdjkYJeWs/DonkrmRjKP3gcxcybXNnL9Q/fdN5+kVES
Nq/rD+JQ0AW5aeIVKnY75w==
`protect END_PROTECTED
