`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LYwxe+X311MOKaGE+HqKt47ao+/rX5bCijXJ75sVe9hxi9RiS1Z/LoJ4srWLUNfK
60k8f4SGR9C2RW10ye2B4bOyU9WIfIKoCXGYoDBTQtJHmTmkJPul0G9hGzUaYDVH
z8SyUtEJX6vhvJhmiSC3XtmAJ3knmPd/v5T/RK6XTsJrM57etT5oRhFrAcgeJCtW
rjFV1cwyzSdQEfZMyc0byoFnXPFeTvsU7HF/Z+1fLvLW0GkbS+xA0TsYKtUe9KWI
288bHbrzcgjdfkb44++z0o7f1O6KX3bdCwgy9L3a1yny6pulEeKfSWDao53xZiLC
tcw/wPFuUmuoSEE17IT1uhcQBtsw4HzznNL9xIdab+BQxLNVl+gJ+QDQ8X9Ywrsv
sgOvDmH+ay4bFKu8wz4yoF6hcp4Hq4BmwQbDRuGEfHaa7GLjAVqShEgRMo9M9FVP
KOU9auSvKyRxTwvXTnr4yIUXgneg6ZROlp2/uMnG6qt8xWI0kTPiXVvsopsT18j0
9hcqQ8Ui58SuCHxLoz1ADLwSOBJWFcLFiJTzEEchd9/PoZHQDudedoRvMe2qAF6V
dYSROYI3wgqiIE8eVwmgYGzO6sJ5pWqnw/Z00BPiU/kMx7oXpbFqVoPTVPc37/ul
asRQ4riFATBoZkZwV+viavLsoZhvDrbSb0jX2KT7rssHX8+S6R2jUMFReqShGI1a
gD0VI07ufy5yFRm+F9pg2a0y0uTuTuZ0o5f975Hk5Yj2qqJPTq6r//k/K38Kq1cG
zNEJaHC7qUk6rLCbEYnnxuSXtySnhVARXndZJGGH9pt6OOnW2AyHQ2kEo46XR5uq
rMiiATVqTaYxhCzOtGl3fQr70J1wfwmzNDY1s/4YV8xyeAyq5GqTH6+iiGrypAgD
awMvEq00Pe/7FjyAdwoOSrwRGsjFXHZQ+88sjHxygP7Mg+q6PKkvEvooH4zApJ1I
ABcz8EvuY59swYp8eE294HT4uS2OUYCy53iwBQAbBfqcNxyB87LJ5CvPOyxZ7wJI
Nn3BIx7Y3wUC0+yemCvrCMNjBMJ79JAn/i5e6e9CdGpLF6ddwzbqCbJYyw/I6yXW
wfPhT6KgDEUlvyYYV+Q9Jc3/Wuykh/vTi3GDjsM5syXr7Kljwc5YL12fzrhplGdz
D5jcKRdhLDluZ4m9i+eZFGRsHw0+A+USKnyhz2a0hjqDGJOxP0YKV27wz8mdhLqi
q1v1C158tYTlWntA/9c7Zdbt70A4IZdsUaDUcVFAy5iYYYPENfNfvh5TmZg2moXo
L++TCKJK8dTKOjcnBAWs9hS74YVQFpZPlooTL9AJqPe8c1NS7Xd0hR2BkLvyCCVb
08bo+M5TVLBnA/ndzGhjqR4+TcHGzdNvtYAatZ8SvKGMcIejiSbxbvhLK6QCpOca
1yRuBVGkYpXNeFsF7SdmnFBnv+v6kCZfTHn2mGR9EexaPkK+aKgmDY67+k++IXxG
gq6leBSDwxKAb3n4tgmtGD78bSL4e4Ny9i7hm2+BF8p8Q+4dsYIC9h59u4l8kjiU
VoT/8Of2E2wieCydJIUEr9QWvqmgCNOG0p+Lhtug1ObC7Tl/Qs956gAG8Rb68wl5
eoLCRn9SJ0jVn40SjFhsv8EjmntcbPv+B1jpri31Ty7a/6rzm5RiJkZ61J+oyF4T
k0tG6spyaL83OjeARtZLkOhTZdkDdBVzcBBf+hSiHEuZQ43CpmmL3d5nuT4W+WAh
tgqiGKh7fSl286OAonUYCXcFuYGA/IggH1LbsgyaEVZ5r07YYYIIoTM2rIPdFBGA
CUW2e0hVWhsKw4aFnENpEvCmlAn3mKyfjqaKuAFtkD2b6ufe6/UQqViOV6T2IcpN
axCY+2+7l5NPnYgaHe/oFORiM8wU7bVWBpbCf4wJ6kA79/iYKybyPXqbE/icL203
`protect END_PROTECTED
