`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FAPgOXbPRDh6dqJ/97RT2xa3Hd3NANBsD4ylElYvDdzet/D+Qk85hyS5R36drOU0
Jd/26i4DIAyv00karojtjKFrvuhZYOzJ/NNZzXUOz/dKTtQqU7A5jGQtuYso7v4B
06bm29NjLHsBh3TIhWb4SVrzIUM2YXvkkwRUuLW5JUWNYFSQlKAmKFeREZPV3iQA
0JOJwZPYRfaVey57cE1uXD6NoTa5kh2x1mN89vg2IzPx7oF9XRBFP0cwnl2IkBSy
2jMwYj9hvnlJj8jedqcO8X3mgXIm1c8BowcwKshhxwocIS4jz65ODNTW4cqjEnkR
aQX7OWtQRhBfhnaT5yBCgHfaVjXHM/wNTHZpRkPrp4NuzjpYk/60g+kf2eDq21Fk
5lrt4YcaqhE1cxAE2XGFgYitxfqAojWIAdkmAxbYrgxUszTafHRyfYvO3V+BgoId
sb2pW5dwhAmoyFL8CQYhUtCX/1JbAkvdbB65Ye19upp6Vgalpis2m5sNDKAv7KUT
9vfgC0MgGQSx9yWknzHOtNXNKZX3h9IZvDH6KY5c50dyLQGrhJPNdbZzEm1h64ho
TIE96+QTKToLCEBGY9Fk8BEb4omwta/YeHAPX0oxCqqMKSOuNc89fv4mvp6ALm9i
U0K5/gONwBcQ9iad0CqBbPtss8RIM1a1H3wh6rcUW88V7993iNrX4Wjwy8JXr7QC
oXgXzNlMhuuAonH8UAxKkEpCmLGnL3jzrnb5ITQMET7nvXdnPeYUylid1huWj1aS
2DJ0WoK8MikNDyfS+dLixc1Nimb9pOo7zkJdDzgDJ6uoi4WWlMiUKl3plRB6AkfV
NwI8mciO3ZXwsVCLqtbkyS56ZhKza0mIk/CjDkgXSrNBLOH59IFQa1Xh7x3AzKe+
3G2LgUvQfq0xGlLtUxM2z8sAqFLRSq5Ak3PxD5wJeg0mWLe5/u2hYwTttZiEQTbh
p98SvUleEYcSPI+HZ9/D+JWhy+7NT51LEDkKiWa1wD0Gw2hi04d0lBWifHEIYEI0
9hzNIKiewq+WaGzbC93jbyFT5MPOIa9IhO94eNdHiu5+Yy3AuQgJfXD0zT+lQ4cW
`protect END_PROTECTED
