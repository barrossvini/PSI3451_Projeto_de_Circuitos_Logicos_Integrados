`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQRnyAzI4oaJIM4Jw1zKp0NgH7ZBbrQDC6o7puYlhLuS+G90LHEY+alQAEGxXw0T
nbSqSwtS6syjUHhp02vQ070DCCMqQjcihCZOAljC7p9WqXhualoqlW4ai+vd7MoQ
jyv+F1XhVH+74tzmGDaow/g/s/+O9C6u0xnvGz09MxfkPlEt3j9kV1GSCc3zDgO8
k2cKO38BOnKgaODvbdFz7h6YM6GLrzllooLyxZBy7lAO+Nq+B6t+PoViNLKPxMLy
E+qV3L8+r+p7589cujMuooPlCEpHHLg0/cLdjIf3x1/N78ZtVsvVJk7IXStpeIMR
rc/9qwWUTeOMFFHxlCX61XLbrgZ4Lr4oE6H0MvmUN9fGdcaJM9XYLaha8ytFUEdI
W1bR0sfYnM2KbzFOVIavqec0UqzU7YzvYtvSWX9V5r2TxQtq0DqE8JYbM97Fj/b4
`protect END_PROTECTED
