`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lLiGsAoF+cXTxHXUrDS82SRHY2wVuxFrv8sAq8w6MLlE1VJ0oybiOjzXUw2kzQJC
XZNgaOMlIRl7wUeF+ZQ7UHOLWSH6ujRMKMBX7290h0L56vbK2fQpdyhb71UPbxON
qqB1P2Bb6Ys0ZsQMc3D2hrSCXTH6ZmU8AcB98nq/u3M6Lo1msyFnuT2pAQL7rFu9
3kNqWxxbzvTA6sQDGmo2NrUc3lGoFJyt1imsPyDtX6HjGi/U93UiUXNHa4q/54FD
uXncybRGOH+AyAYvg6VP2VJ2fQPnocK3SaulJuwDtn2il59QP3S9nmLCLld9ZwcY
XzYqoAX1VapaQBWiag02WUUPlFE6UaLWsJxxu3YjtWzTyoYlm+jjk/idbUzFcjCR
P3RsHiMN+oIrZ8mgy9Ke3JISd0OcX9EWutx5uMAr++CULU1AyH1j/qbMQSNC6+tf
ZUpGrb/IMoYzgZMrZ1QAZOUKVfl+dnaBdKXSMOlOSItjW39wJjtGiCDVfKJ9+1Sb
iDhp5qF2X/pcgRVQHwXhxsiP09jnmUpS02h9UpESjZ3Jno/T3YJPtC+0SsawwKyq
sAIBdpOVB8PmgemSgSS0uEiwAzbepVbYhLnttZxQWnC+36uSJhFUX6G8eZmAdY5L
OSNVBxEqX2LkxeE3EoUseu7Lwo9k++/zePknP9n0h74Ot2G4TXzaKyuM5SDzCcjD
+Nyll+DXPwhwhkNzkHrVBMIQBl1V5Nr/UFyC89tNoizso2XTatiN4Mi2Izd3yg2w
j5im1LNnRbAdiPKX1O/M5hoUQLorN/aH5MEBrLxvfYIGMN2eSlwNF0sDhk67FPBM
7rgBMPuf2mXO1ppY7H9D7T9Rys14G5epk0jmmoaet2o5+H5WeabzJoKk6gvn4KHd
t1YVye+M2FNsY9OxizkN4wrQwK/cebUOEyNXp2UthPeOsLI9ejgABuT+8NMuBXTR
OouSzN/3CwzziaizijLuQR5HjEEsd5s+Ab0AcYkuPz3Pfzx0iTwVEYgkyPwNFgRY
pvsxpE4+U4hoCkDNH+prvDAkQhoLKEJSZt6kobdmbDMtoIGYcUyWWFQ7fGloE0CQ
FTblsM2jeetFx3oNhdvNW1fhRow31cY3drwww5wN/iAS6k4Qn85ocl9JOAoKsQbr
aZmIACMIYSWLhrEu7o2KFKlL+3Z2xW1idXm2e44svNSeGUP88pLKoWx/BFyTuo1w
5PWL8Q2rqkvzAUBR4qKDrajqmj4Wkd7vgACNgYV0nqxAps+v1XCct8iexrgx1BQo
fxUFjAnG5rDRveIBWTRN9yLVeymb52s5toaleLRJNsgn0PiEpzx7TVZt9MenajdR
gC3RMhs9ojc7q2YhPwCFKjo44sWVl1FCC9WUc73LeulRiR3hyYlScXgdJyxt7T73
e/tPN5EezeG7rDCw4m+n7sInnTR9hY3AK7tYlQF5wZZVyaNylGWXRMWadnMvA2gn
CQ2VLWE4YlvGjTg8tXuAa3tB2C8N3ZzaWlDlvra5dMb8dl6YftckpLw+PmWce5Ue
oUKQZcUWmT8RW/nBBBN6P7PhvJ6TDTRrb6EciUzNxMEI0nK9J/HxaQCnT6z+3q+x
U9KvJYbSjeXUI5/FNHGC9544JWENEGrQVEsrXzeEKl75H/AM1GyqZRSd/cuqbB0+
91RGpBZKKJxrgZg2ur/jy/38htTJnyxavp9upnfmX9IWSBoSzpYurhMoGN1V4IFt
JsmjZzOeMnQ6Ubv/10n/6arnscWOrSiluB04slteP0bfE94TeySifQN8Cfk7LLFJ
lFCDMGf9E6eYVrOGzSxJUuuOr5VbByecRHds1/dLxQIjyepUcRyElAn2ReCCrEAI
oKPOgsTbcED5KUqXZa0+eMLJDQLKZGwKUJiQUoiT6n3I/vbmHQIKBqOqdoRhV/Uc
Cl1s1Xtgw6YzlkM4R3Bf6fdPy2rXxc47NzTMRVbYvKJzCMOVDab4xyqL/UCEOjZw
kzWhqTLEF+OO0f8hTfLQwRy2NX5AeKuWzytqOlJeb8/Z/dQRjLuFitn7TBezwCIP
u9Yk+WUDyh4yfAUsIcbYOX9pE3tQdVf9GPRTTLOzzKwotwBrDhFhQy729N6xO27B
AwIBH6YPfdc+x4WYs0ofbCr/S/tThUy6rDatrOV+7I2FuPiCK4mr3ZtngbEjBa4i
33wIFWJVcI0Ztvf/C8EyC0SWloNTEstOZp2ozyLwpLrRJt6KMtd+1BM/chR9Cih4
eCrV8MZynVf00JxIbau4Xr+ejvqR7+IlDtP+vaxzfJefPgcwhOQReoM8AfDHJB+c
VIO1kSYOk1x0Rn2VSOZLbTiHECZ5kMibbxUuSVSjo34Qhdp4sbzMtjWdrppmka+Z
Ne3vh38RdJ+Y4rlD6qsoUnJb0kKcOC5N/sDq3QpEazrTQ7tnVIbGQFVKUq8GM3uQ
xHMfsPrlqr5jRbw2fmYnng==
`protect END_PROTECTED
