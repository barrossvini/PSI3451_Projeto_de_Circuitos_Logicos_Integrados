`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lFqxTJx8kuALuQNjv2TZ1xkFb/OGhHqV7LXmYLr2WRDMdzC4jC2W8hPxS99frG7/
jHquQ09YYQzIYd8eEVK48T3a+h3yV55vhBog0zaHhWUFYXtDsCDydAfKyX6tJ/O2
2BGA9GYL6u1umf08ddgNUOvIjFUAepxO0nlsy+Yhdi1BYpK7QzylrtunDZe9Y4Sg
GDFKa2sZPIBRVaOy6Mu/huJhTnL4G7a+Jl4tvpTHWl2XgqFKtfLbsJ3dt+vgVuez
owHFBSeIcRThD/o4/YGyNtwwigrlVo1xwckR4ShBgRyYd5tnGrQzX8ne/OimnduN
OhVOO34rOZUEEXLc7ebGJE+qFAqrM3lz+y5ymYEmZtczG9maMQO2TYueGlt/d62I
/ndRD/wK850qSBqyR+epx5k9yJ0+HxNc91/gSTX5mqnCot8A8VrbJl0khQsMFzSl
2jCDd7IBjx8aeiigLGXa/CHjCHwHEjazHHJe0BaYPFi49HQycyX1NvBiqm7z2l3s
TPy8oLmUPspd21C1Fvcxk35iqdT8QxtcjYpWP6xM/BhPzaFFdkNvf5xS6mp4oUy6
HMntiq/lmAyhX0D9xYyFfxnQKLk/823FDct8CDJRF4P3uVXqq8bNC1c7HUa8kUR1
Bh8ngwjyxB+e2gXGb6rMnHZ5dLLT8qkI2QNR7/rM8dSwZ6Qt3E2km0S1EUq6WxaT
c+oOb1UMxAdhgRuiQT4yog5avl3gpl3sGMev5o/uCji/mId5qPfl0Yppgw5poMqw
wS3sCfM76nLl2CuKNmywwyYMPUkq4YNXNdVVuQp111r+RNCs+tXDyJISUb4YeW6v
8bHjpPblTu32sViiJzfLxwUVYQyz57bILSNpAh3qLuDNrmUCpvhMOdpujy/XZNkT
OTpHI3xIXZ/n/eL1gILmuKoqXQzzGR9MFhiqpHrMYfyuNZDYCPraoboDyf0g+1Fp
hyQQfMEQZcywHlq6eCU/zXHLajqlGZwVAt2IaSl+hm6VEKPWsXKLExX2hlvbNPra
54MW5C5m0tNuMDeMnmG2o2FYTWwdlAuFt34ol4fka7E2s5978xjDqnELd2LXAhXd
a8IhW+AfFKmoeLbD+w9tIv437E33ppBMTvRG8r6g0+3zcaOndl2wZHqYWUO86nrI
Riu9yhC3ahgfoivHLqeZMMNiYKWP8XrscVgHtrMMouQm9KZXTcZjsOptB8ElWEYO
KTLoKHnsRydd45MgNv2N+Cxq5NwM0Oqvna0/pVcMy9G1DmRMM55QYiFRPJBAiFEy
3gkclaTw5WPqh051RHcKmnRLUIv9/ygzOHOWDC0S9RHWb9BDopDfylDh1vYv9rDz
BlqIJhICPgMJfJ7bxVFaQahoxEYUNSeBVcV5luUwpBO6FL3+NguOVrmwPRrODSfK
y5E76NubjP7ISczkuz9n0BXtE908szd2n6Y6H3Ox9Js1laXyf1LEvY89QmhCLjqD
`protect END_PROTECTED
