`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DiQHyDo6S7Yhozp3RmIA6Tf/wVKwL16tydh4njJSy9fJAW6DQCNfQul1n7dj7VPk
HXk+aWCGeMSyEe8lVkA02hembyqkdIj5FUk0b//sti5N1oWWEl5fYYTFwJsgzHxY
+Vjjp+vbvMqquzsXqgBLGe5capnmGN3+tCS+mO0J8D+5qsWL0PxQP5BPwIGKqHUz
vXyJ9QoztY3Tl3y0YaRg3nFrJrNIFNLmvPAqOYrfLOuQvW45IeJBQTJS8eRpZwlz
a0dy8Nhd80XRgHz6G5QjGw8dYXOLqrM9zhy6VhrZfFRT8UNSz1KGqCv4g65gyYpy
GzNLDzFkBmM663dPt7GcWmmm4o8C3Kd3Vy9i+1ogAMbak1nCaENUD81MMWfSmhZv
/hSIWqGXFmv+dEiuVDZ+jSIPrCgHbRh23nLU38jllU0jayGqocSbl1X+U0zzdDwK
IgLxCEO+hk8Y97hjVdyNfEzkYdDess2ycscqFpsJfhnlF/SPW/IKg0T9++jI8w8d
xNNVkR8orB8iN3ccEjQXg1PIaRsX2WeKSc55lPRQ804V2v+Bee+Ylh/9ybiCN0dk
sxFMJEJ8VY3lNeYZ59fgQYUd33fNkBAocU34g/DXOOxI4rg80+lOQw618qVS+JX5
oDEbeAzsNr4IcvHdqLsdg8p08Vl9bliX0BfPe8vr/Y5yhq4hftpR2GDmZzTEjDH0
vCzou88AnD/iKeDi35/+qfbfV0XYQDPMtBL31jn+B9Trv15m2TobzgyFsmgWTBfd
a/o1fli0GOojYiQmETU2794c/VbtphmBuM8IEcmtD7iBpD9cWaba945YasgRPUe+
uz/rwF4diblvxk4g8OTAUWzjkfSKSD9OMFpROr4bi/fGIa5ERijDsAMtD4NcDhCB
5sAGI6LBDtKQ4P1RSk9DwHZFwnCCZyIQLWIin0vxWK0CWHMNZwrgjihlH/H+Mxef
5Y6avrl+y0SCaj40Q1P9iJmE2LqRKvcfmab5RtRsJzv1lTO4xGi+g9EZ6LZLJkKh
+h0ssmOrWdDQjo1czQIsWgNsWCfgikzKngB0NnMFu9EIKzPAph2PY8pONrwbgOWJ
7F41qF8aIWoUPQ28VkRivGRBGZMjyOU4wwaqnZlaOmrnK9p6CPlT/43wsJZEVTU2
+/iETL3N0IbssO9YueWtzi1W9OELMq714AmFOx+lab7BIAwfd5r98XDyKJ+A8KmK
eOtMuxJu7lAAPtVdBm3DGsacAGHzlAdkyUdRx7WSbEkjsT3j5Ovp08d3phVuk6Ge
Vu5FdodIabs/+lA+e9U+OJ2vQ1pbVhIL+xoD6S6xrgSYcoLsg1l5qr/GvPYA28Pt
dy3CJkYw/zj1PDafbbkBQjRp4ZZrvkkKi7wyjWk9FqJ7Xii6lKK37bVhstyxdxSy
7CjWgDKfRWhRZY3FsOXqYdWdTTOH0QS50huuCcjLoQflCp14O4hpSCwlsCqcL3Mc
J8jiBf4Igioi0e70jdV9OqCL1IGZRX7gH0LUYfPsv1QHQC0IveOs3yKrKpJ2pRAe
3nwUxCb3PVya3cs1BZkgYL1qfQy+F+dW5mMZTrWQwxKO8zKfH8FUDTRiTi5Z6Mla
TFOKmB/QbFgsGPQBxmb+N+9Gtb7DtpIs+hOCZp3FWifRQ93t1NBok0fiN5vOTCds
ujEkIAjKenPeFeZbTEB5Y5v6Mp8FjBAzBdoGJO4ubQfpivlOVLQ4ITHS3JnMcKTM
8Ufxl/2Nio5wJh6yR77HvjSxSn3pd0NHYzN8duo3/kc=
`protect END_PROTECTED
