`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+34+ut37BHWFRjkKgKGiIWgl7gsSvWn7PG+tfLcItMoS+23ARCwSEnKjG1HehqUO
g/AtQYHGISiiMAqdM0rKgsT8cCtHJfiMwQtupqCKEgcTVM/N+BfZDIFn28UCsUwa
Mp0LkeWI1cFm9d6HwvDBe03midcWLMFSBVmI8vVfvRpn0JrcBa8Jl+lsivTunWBB
cs4Y6JQAkil+3Tb0jXHiqZqmK+uKpHPhIQ0iBvEeV6xqzisYSfxVFOLlrcL+jK7x
9jx7HHqiHiXeJ+ZYJr4XmQwYy86+7TLgdtYhm7PnZxvWCJ48oTdjBy2VgQVlhiHn
AJvqv+m3Im1O+y5gE4AreVNnfWo4UkvP79oADnoYmIBrrWUz3Pmm1WXJF8UUiBO3
FhKF8bl6N6HTQAB2LdzMenTjfnODypKbThXvExNeBb1xrIIJyp3YU+qHuAsJ1leD
3z8zo/+tfHgRmNe86XoQtlQgZQmKvm3q3Na4+k7zoZvwmxsnjyzry44oNQz2b546
5tuoXL2x8L+ZN3OobsrR6QjVRoNIfssyCojzJZ/um+T6o7sULN/IN+JQXUxGeCzd
CwODYaEn6pOPru4AURgaYs6dciRrX+EcA7hzcJ2oIgNFEKgGaezsakCA0YENl+8N
HA62QMmpTircRsiqD2t6ZdJRu64BNoRNugrDXqhG+ibSGLd6ZhL8v4ljAkI5IXzv
8gmMzpW8tS3bWCL7z8X20lznFk0khp0/2bSGFjc1eA3d24JlYNmhXohiSNoGGE0P
XOt4rFIuOjemCZMOepjGl/ZA/1IkG9blj7P3aYnm+/J85woCRxVdebZU0qTseak3
oSDl9hwltnUp5DHWHAFXdIVJq5AvL4dyViWWop/OPRN2Wi5oPA2bDbrNjvFEeDvJ
fy1fYQh5JCJXywqzBgO494AWy7Md3M7MgWYbXyaUMXVJv5WOTQg50QMgcWti1q7A
rGewGgjuG/bOUlT26ETha29mqe3AAheVqA0Pg9DP7UNEZZfjhMNLY/K/LWtvsSmF
frCshBiP9sGunIa966tADhxhc+pg71vB43SIOaj9PiNZOCVzyn+wZvP3+HRHPigC
sgQFGCz9YqkxvQMGdCGGrJf5qQ0vOzL8hVHP95K0LPmp3IL6eU8+wE/1lRK1e8WX
IS9hEUy9Eev8c6w8Pbq2Lg==
`protect END_PROTECTED
