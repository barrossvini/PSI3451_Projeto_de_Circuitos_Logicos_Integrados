`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eorqLgPuDqmJKy0G37hpCRByII5rxYDKYdSU4jGPFiiAioRo4D3ylFNvjNh4QdD2
A8IqLMqvuxRnNX5VHdpZBDqaPdpTpWXCLa9XLfn6EkFfyU97HS6MoTWKi5IEciNT
NkwfJSBOkH67T2jKT9iVSKHK6atkHHcWrdv43OfUdu3W8Da/wwJHpoUs3RtkWA52
Sn/8RXk8PV9YsLfziBAUz/lDKuiQ+BxW8VR8Y18a9Aj9Wc+LQvIuVSMnpSokoBHM
pZHo51IJ0hImWwK2MMid1ogLJJbIA/lPQVQEH6D9q3iaw8w1VXzm7coSI/IXWLfT
bzhmusS0FGp0MyA/VuV2XEhiA02mLoD8VnqvVnT3wsootT5DDLnz39WMZ1pw8PoP
S0PNfLTt1Kir1GwWiOtu2x7jGsScKKzv0fEEfAuMKo9//dkcwBmGmP2GbDjnM9IV
d5AzLsWRJh/gtvjLi14e+YdoCIyboumRXgH2FHLtKT222KlomezqkBHjYZzHvGPM
gJRRwqS9hHEWmyEx69iLXoPX82hG5saYrOxVfqrAC0DyedCqMBTSibma5s6T9Abh
Sqm0g9nvYDBHNQM32FIv1cZfuKbiF4rwncbr8lKY/8xs7WNpn8SuaQwCZCjiglRb
Y1RvQ0Tk0mv7hfsTXhwYoJZQGF81hhpqSY8KDJncA9HUiFTfbkJe5gLbPflchEqN
LeqxibRPSFpjV0+TFAQMM6UvJmYbry2ZHXfqlaal8jKQS8rQ+gZ1AvMHVz7O22CM
aEvizVqmLMeE0AkSvVs82D2UhkPyZ8o5LxW4WYFtFBnZvVV9SaAFHjbjYjuhh0ha
P3Dgb/H4q6PQknvlFX2YIYvRtEknSxHMftI54S9c3fXpAfXu21zrE0eeF3DCluYm
Z0uTePT5JfBcRyQa3ipXx50WghUoHLpBfBpcMafgR+MKAF4cA5AfKy456vtHCNJB
ruonHRMju/yX2rwkrj6sJR0z/uQQJN3jvi72BKeEWFrb2GzEzVQ3KBCcIl1gYazC
ktVhIyUg6u+j4M6wH9BBVLbhZt5aoBxw3E39W5QvB0OA/bhqjzmIXX3v4/af6C97
8sfP5TueEjt/6ggIixP+mJgrhQ8bOqD3hIPy7j0uMJvi8NA4ykNwHQJ8PKf7LlaH
YOBEQZ/EMrvhyFMwoLpoPdiUPWqLVi0pWaUIFCReevmsBj6VQKeuFUUHuSoYfXu0
qMcaetZDSLmHGA/iD2X8161TcI+s1ZmfPb/O6s7/5IAGrIV8TM/LR1iOsCkqSx3v
faJ4v229wnjLE7lzwnMCtIBw89VML/pqaXvsVWkJOvz7xSN/GaVybH7Q/9tkG1pH
vasFgt9cWZe2Iahlhv4txz3HdbXR3f4mQ79RxQdeRl9lmgEIECtFgmga1KfN2RWX
JJ4KLQCuUh/Z8a45yb0rWxHPAwxzAPI0ajnT5IKGrxgdy3z5O+/bHlcdpV7/kHH3
I53hikQ7TKGMe/qrGD+7TPN3JXRYrF/l/Alnl7G79zIiYOw8tV5C+hqnxZh4SRVe
DCJifJtiuwGa9MYGo8FKCCSv+Dt3OUY96BHdju8B4xsz021iJ4OphwHzDoAnKR3j
61YnMLkrdpoopW4dgd0B7DhcNkkQLmFQULWxpd1I44qYZfk8SrLU7P74LijKAb/H
M+Dw4ryxX04f4TF9sBaadugttmOOt4xzn0SIM13FL9y2AH2NKMv5oKfyCZmwybxo
/aK/ZNEAmZ/hbn5xV0IJBAcRXgGpB/NjsFRzkJ60MyoqXqEkCmDCOcX3dzaWJPB2
Mrl7n/R087d5DVNiLWGXkFcbR3t/fesXB71dgHZD1dkLuEzMBBY/curJJ0Sm7+9I
u5JjphgeeUBJVgg2mE6gDqdvMvzTHrJ4pVQ3EN8EqBAgmuflFkBj1somVyTBc5WB
QPOVqLHcd5Doq+K1XFhEnK7J4ES7XGURUTcnNGKstWbD2Vlw9SDjpSBrC09/QGN8
zGCVXGF8fBYCUmtzWyFYnSxaOmDXonvMdFzrc1Xm1Yuh6L+4hvsRFmB8tNrj0Wci
S1ajDNv/9PXXVRToZdxgi96sQWo/RduLvinbFD7slHkv1beO1k1G0uCPkkML5EZ4
7YTM4t85vmi/tFs5cxCELTdeoZI87W3SQmj9Il86jP5Q6gpqOxn60dUfsS9HxgeD
JVYCH2K7esMmqpmURZJUFp0uwsxrt3hrXeKqFulSzMoWlfCPPb5z44bL/lfM86dl
nJbSfe+dnj5bexN+dFiAAUhei0hEZmDBWZSvtCxqDP6LVWZkbDxLXOSLFQAzTKGv
njgXTmvPOGm2OvzxNGMz6noSpX+aIHdTJCfcxdJ9+C/BdkCgGOnj20v+Q9FdImHj
OatoUI7UueDxYySDUFV9W5nX3YaKCYre6y3t43uqxdWFuhqejX+1qSjbABT38+bh
pvt/NEYu9Ug6782SpeWlUgEIkU+75IIDubLzGOxoqEFSVe1aiVJnjDUmcHRqUptW
udO//3ehwPEoSIW1yenwxYR7BxSw2jRVJchp3UVaaIbhxIBf+2sI20ViF4CWcdLO
w8obMmcy73YOGFTHKgHZhnN9kzMTTmZiB3ALvJQ6B2BkpXRifSs5XLC9ubK08Hao
b/4VQFzrwf9F1co7i8O9dhzzrfIsUmBwW2WOszjSXyl7gl5kZKQsblC3Z6//1j/b
U+iJpLKL5e84jOYjpGB5dZi9Gme0pKKJj9JcFFaP8tloDxdWiKhFJRGndNFu4Syy
DJgIFUkJ1zVrjzTa4LXNiF1Kqv+Fo2mNTXBEs53vzktEoKG7IxXXJnqOLDncrrOe
QlIyiGCRmzNjqtCvL4b5dRpwCPgCf5y0sWUSObGrWmG52SJmDfUEBmJG0ykCXIlK
0sV9E4/rPe3vI9hRfFmrOyipYpQP8IK2peQpxbHqTUnBgjfWWvtEGSC7nbriMnCs
nsqiRL20InDLFoGkfBM5F2wU5Pq7maz6L+dLQgaOLQK64jTLdMjju1b2HJN6CMlx
hdM8itXkWnSzVOfV/kWFIoHI45uCYknJsu1GG083HdsimMmjI7XqcsBGSzhXi33h
pghFeE/urFh5XqiEWhp8uXTuTLIXmBeYy0vl4wVSNPSLWU3hcFjfsOm5220DrYDG
9oYthPkML6P1c6n3hV0+/cFvwEZaRvZberx6F7pODp/I28FJaPYNgvshVk5crKlq
jHBrx1nFIYOyVVXeVRK4mZI3LSCKt+mNDHaNXd76njlvFoZiEfTCP9OJ6V6otr5s
75Mw68T4q7nlrK6AMiyGI4EGdexAkMfB91PO5P7nLBpaynyoW/9p/+ZtLYfmYOEj
kDA1Ykh4yPoTJoh8NQC0XrQh9GT9zqIslwc8bbaFp7q8UDWhUgXX7qYKQpYlqZE1
MdZXBk7uU/ByWHACAgHkGXqneD1qb24YW0JO04lvmEAEeWIWsiOKhwXmtixbIooz
MLm/FyXjjsOsB2ih0tx3RVKyllG5svqaov5KoEGaAR+BCAf7us42tZ9k2nOXK8L5
oCCzJWHjl51RgbUJeyC22KNvitVj4vT3b6XxMI7mHccal8Jlj3vRVAtoeIYnFBXb
dsoz5SP3MtdfVR59NswbOvnXjZ4g4lRdvos0r/6Zgb4NooZczAUcS/CfDZUths2H
7hlMEFFmmjVa8VD7d25gnYu91JyrbgqA9IAtLF2ZnLqO2fGcVgmLbMGCG4OubWLo
uH/Wrjnv0oy/2rN4R7X+gBP0ooDss0zeswr33ivYYRKtR6yb7cV/flTllExfJwzT
NU46hvCiOdBewNyCMOpnPjktDRL9iyBhscRZWODuwLIy0HvC0Fsyk4dFGmb2KKL6
GczoQ7TGWnWhdwK+z0jhxmejUHRkjQpBQ6v5w23KJxdhTm+isbMZL80VBEhmqnxJ
qf2uDAExbuJPGku+217nlOZFJNHE3ikBtPRX069lSH33Nb/XDnMl0WGHuTn87t8r
4sf/NxjNOgThP5p4px2PzIt3LoZGzhHGYWdaf1HxT6zvGNvGvibjQlCRGwuqFKek
n2C6H1hdS2/ynp6AOsot5RWZ9wpN1hECKLqD3q815Ijdi8tgwyFnJODYZ4NjijSd
h4IIsJH8PydjBmMRbWwniCgFGjJ4mTVhcoKCe4eCCNW0SXeLAJlBamEb6f63NqEd
BEQk71W8xh6zrIoSsMRTv1fkudZenCCY2x5q5pl0pxURt26gE6+VxGHWJaXUWb7q
pxGzYbGWUXH0TnQxpADuweYof0i8rhVmoYMWhopVh86WHSsDmcAswmpDRoTHX1wA
GZHRdDIGP9LqC1p2M46welBUukEXSV0dijrkhdRvY5+P9KS+UOAsYXU3smScoWSc
mRvmw/o4epRlII5YzBkNx3iYkBOEwcvp/Hd/PC64Qk2l4NLh4jykUV8Pecqr0Jfo
StnjHvJPqFrWlQMi8WsNbKXclQ8iRrPk3NRBzn1XKgakpRBwAh7ZD9Cl63Z+a3IF
c8WJSRSP9EUyHACO8l22IVe4Xrqmw8jmCE2HgbBt2ssiMoWElcMSN7kDg9opunFO
E5Zdtb1193knAgfo8oEz6a8SwioDARKcciOCP6l9LuQN1ltqu5kHdch0OREE04jB
7J/ydZS7HNTit9r/lxnzmuSV29sROtxw6LtY68n8+uSCr4d2ronoKYrsoMlGUVme
lYHahSQMqkoQiTWOJn3W5lwCljPTfr8NMnOMRUR/S0o5k1YZBEZqnzZIvH0b5pak
zaVV0sjGjylOPkvOKOfYaIBCFf9JJLpACtb+FlywvfJRHXFBrowXHX7IQQvKGWvS
vfgd09gu50/bOaH6D0xf37pRYw3KmYo8ummgpIVbTf+ymIHGG49a2MI3C5/1MG94
MENArqg+yqM5aLF+qw1OB4Qhnesn3vyPQSRUYEDJ79zegq062KIfASKrnCStd12r
u/MpNU0357rFfd8RF7x5XjBW1zGksYs6QNhhyqvYLalBQNf9rpxUbmMIjqFpOd4X
oib8tzMlSYYfvo2BBO7aljEvMY0do0gA0B/bsTrqMZQ74Tpf01Hx/4p0sHB4qdp7
j6bskkE6Fyc4+SRiiruyhHeRtPYFKcJu+MRnhlnp7UszfCETWbb168VeBk/Fgflh
mmSroUcyXz2JRQmQ+zWgavojva41UXu3vX/6iQsjuzFL81j1LcIZNYvqD9hMFEdJ
BiWdEfwfHiWNyycueX34kqx5R6EI/6v9V4Pg5L8LQVoM6NtopKX3bG4k35UKHWpU
nIspYepwKW9mMoLlf3ODF+7hIUs16LMtAhNYW6vkTi/Ox2yDVGO7bYFuAM/4ZHPI
cXp9W994EcQb2MUCk9xjVwpGYl+e2ndllrx26Ofvf6z+Y7Q/NtAxI8O34CHjndmK
LXq78kqdO16yg/Xj7SCGcJgcw5m5r+9bQE1pDU9gfyyVFSSEvSuAWloLL99ImXbF
VATfxfkXgCeLrQ135VBVwk2bpNpftFJvm2xGo6am/dnK9z/A4R4rFgLZhqLnRih9
hPUlRmyTu+Fqzi8YQTfiE/4mcukzwLUcAqERirGxcbGRBrvOhPffM3Bbem5QDpBi
cmYqSrQvM9rqNvsA5TRLwr7MBI2wOpSu1t0q5e5AQRUTXZ7f88i5OcCraMTLescu
xyIAADMnDKOfPHmBNCNyWAk3SKrgcExbZGB1L6fNalSbH97kDUBVggRWGo7UXxFm
o+3fpifZeDcl1jgX9RDatBWTQNxVh66iLNwtCd053vHWdDCtZa9XAzemH6sxtqOS
UvO9Mvj+y1AkgGByFGYxLrIquC3Lyeec7xorU+ePH9A179xARaJnNoQL44K60KQ2
7Edgb3a/e179tYzjPPP+Sb3X4Luh2QMjAokyMFwQEdm2fnSg2Cj6P9JBcVLYNuvV
z33iFVNSAgyNVtqMDs8TAxXFpRsJfkkYYjtpC3coyOIPonw+Ec5Kp5u+yyoP3CGi
jh59q0iEJ0+gV6SVxGWOUNv8z0jbVKx1Fzx0/hqSTWco/bx/C4YctEwoVANq+2mC
mMuUbkqLPwULh3AkeqsqEbhyRAAJAtR++IAJa4whd2lO2NJVrMgYvnfu29J+88cn
HZPShVDZmsDjP3OLF+TkiAIXEHArNQJW5uAGmVt/XcRLbjmUW8xqjQjBA25xwdX/
Y4mYiMpWD8IWHp2EipswB0wcBzZ6LPYJADb+J89iW3F/sHvn7sxDM9vx4qN3O2kM
UxxcD5uFpT5b1uQrrYyZ+r1A6MnWny4Z7xNawBNt9OMGMY269AL04BEEdP1WhDJL
WvR6xbrlx2fFNu2Lhr7330mFua9Oc4TMEdpofz90nXWIG7g1QfcHdqvfG3DI+mGA
ljHCg3uLUE8fRZczNGOK5TE1V1TRlggY92uD1GzBfKjFzelaFI24p+Tms8HSHPhT
fOC00qE0SpRyNix5Vr0HS7K8ZBWbKbyIMZFp+BLfQDQZ4dRQYqh8KcSKV5Xk0TZx
gfW0QNNdXU5HfcISjx5YjnsPJ5Lhvuw4EUUem72f9oODmVSf4F+eDJEHxMI4lSrG
ednNNlqYxouw0E5LcYOXPs50TRXfv/YoFb17zeAZvZPXNS1slsqpHZlNzFAir9u+
5oVOfbrBGDIBm2vgsTCmiawRnweR6v1t8ZhJ6EfrXIVK6l+wlUGtiIgEUUesd6uu
OUzzDpddEzXp5hUqhFPNQLEoZsUkBW6Bl4mkTJIhy8yvqx8oesYuzH+ONRqBCawT
/s8Lu62CjbdKsoBwlBPB2ZJnPyKDmXas5X8T7lewd9NXbOAKugm8lRe9oCDxmaNx
wnQFpOfC9Sof0TWtGcgrnmk0Uxao+DY5JHoA/KOC1yahiUGl9+gvaKyooVtq6sSv
ZxYtIKn1OyQK+SyfM2+LU9wsV1NQ3CDZBZmbKejE9OqFiG7FOeC3hbI7iEt2fOcS
BFGdrmdCSJZ7JdGfE5JOiWAzfCvOiFArbKw51jaScplDoborV/bEWPwqdc92ej6B
9ndoTxorj8v3ekLWiwJPfK21SioUoDYV9Jq4n15N0YVzuTCLUv3Zgg9YRMQViAqq
9svjQvrFbKR1Dda5nz1w1pOZTkBO25rMpqvJ3xX6nO/G2kCPco3WgfbK4PPU4fz+
zPNq1yHGxnpF2czXIK9sYsfiLhNuaPGDr9RnlHoA8U0Vu6MahC1eZuuNJyCNn0J2
duxSs/5uiAR7rS02PQ6CqSbYw1+xZJ08Sbp+PlyOiFCpzz//+1wE05cnJ/WfZC5L
42rERVlQPpMPXKl/E3uAkzCM7ZBZ89NC1TCXM5G0opQzcxJ4zx9oJiOTPZX9MeZI
CQikFJ2BRzKi12Vsxe+Qy9gHPgsddSArLME74krC0RQFHk9SteXpeoAGDxZxMRP5
adOjlnboitmnwhsEssIZ5RE9rdEzA4VDI7q3C/OtUX3iJ94ZiyynZcWnVUgtfo+y
pvAEIcI+MCl1eZ1yO8ISMbSFLvdHDRRQmRkKqS9Uytb2KKt7mjf6zk4DbkW2txn7
BYrgDkl2wJPM4ADnNx7wl93Ew/HcFoTbyRMS1cgVTquUQEyurCbaKVudRCMnWkQo
gztGturuIswoYpQUuxdKj43v2qDukVrWQ8v+e311ch5fhcHFv9dBaad96f3AS/sF
5Qx5y/MLiqp3QguexC1d52YTzmNJF0scpB5hxG8KdIOdVixYaLw+NAp/+ypws/cf
K7CjpH0HaY224/W5BbqS+q8kmU1vzrNZ8C3DdTj6506eWNNfepzyofwwklxIjnfd
a1SjWDverF4Bv1p+2ed3vxVtSDpkVOf4zsx79ewU56RkDnQndHKUXllVL+AnBxlL
4zeeN7NvvP0flM2fLl3RF7ZEohLpP0THN5AGKEgYmJOuYQMEwO1PEMmJS1euowvx
G5EKLpJ8eo/9JU3uz9v7LfO4cghIwqNUH7ehyS8LeiEul93uXmxg5jAUg45jJHB/
EIl2lt6b/A3nD3QU++mCK6AlorHb1u8shm8rKnsfAjKP0g6PggsLsywVL6tTyX3f
eH2D8BNVFLSEE1UBcNSx/yrYlbygMYUE1QFIgQJ1pHTjFPjLiBqRSVh9i+N1T628
jZVxO2b7Yz8S7C5K/A6uyVhJ9VwFi9OCB82DW/OyV853RNx8i21mbVwBTlykqUnd
T6Gh9wzSY7/IY2sU1FlZIgKROa5E9/BB7MJPIR7ep3yNphTuiXLLvw63P6L+QhqV
lEaG6mgMMO5dRGfgg/XIqJafBaRqH+WjfYcDYuzNMw19BOenvVNPtr07XzTriYSs
ZISv+s3til2Bw2OYVJ9x938bAtFAYRy1nELfuSvsrdnBw9Pmzb7vbBBDwk6k9KNf
LrPnftVGW6SWtHuqvKDvUGnZskvtM583xpwsQwYxlH9ZqK+K+/6RhXg9o6J/mpNz
UdgmxR0iooFXu+pzEcec4SGd9Lmtzb1QIXPLbOehxp5ZpgKKNHNNJm49WrymUUQG
+WkszzsYMi5AMcQ5w19uXm/02+ie6mGhm11C7PqT3A67QhudMC9KKycF1IZG4tXA
Ryuq2R5uih9fQH7+HW+jd8z16ASg5btvEOslUW2qdZcvH4reCcfav6vl5H/G/u9N
obBMEBCMYRK+blZ8ajRjed3zqmu8kDclXrQIu7Rb4A5iBn0WTV9pP2Zv+lJeJ5Ob
F7z9n1VcOHHh5wyhZ+PVIS0IBbWLbRKFxKH4DMoOdvgAt+tH3VD/Epr+aD1vZhpQ
2gbLflq+ObydWhlZ0Z+KsNBnRfmZxu4kDMNDzI0/kBhgX6WADh/IqhSVw6ucCknS
rcZQOv6eb03Wt9AxP+tw1HJ1J830/oFioLZYw9ZHbdSgL/1g9noUjSPH6SkGukaV
78Zmq6TcBHUy3egxITwt/0xjmmxYZ+2XMNyazmcsjZj2VriGXvAdYvJvOykeMubz
zPFvCSGn6E8TSqrTYLgeE/aER6OZSRlyvYwaMggnIBo+qnpxLIjvq92+T1TEQe+J
AgIt6jqEKUbHowy26K4rZs28pR4HVM7rBa5iJqSxTccy+AY9M30kkGaDblJWB5dk
H1RfF5L6Mna5tV/6n2H+WPYxAsK3fNQhrGlnZBHrpI1iiu9p58Vsz+uD9iUbYZc/
Zlv6ABiuTzLwoHXh1kZGM8Z+Wk2zWAzGoC32VrBOsy+FsDYESfiFv/hV5IDrjRFN
AwyTYc0kX+z1fotzsKO0llLGfqbXlne1MOuvVDSvUanAsQrpa7JESlGAoTuLfGWp
u5Hw57Ws47M+dnyu+aUc51Go5/93+D3Q0VlbokEdvTws+GWK7AHB0QqyR+A9Mu9u
spk04Px+9ix+UfjPQpV3/AKgOdU6cRUceI8UT+rqTLZnSj1hqhpD+iE79FWGhVhj
fz+Uneu0UB9gVIczMKTkdt6SU5yaHe6090mgamDbuXrKpupGylrH0FPwMCyL3D64
f61/yYOV4nT06yI9GgqsTJwFQyJ1D2qkowN8xLRP/WP0rpO/1LO+dOsTzurPRKmp
zQdQJuM/q/jXhd7OCcQUtvYPTWAhNJfR/EsZuGJritI2tmNnd66i4oWic8+42dUB
YfS4LYsLbCMeOKxHAGOq3wQpNUOnGIte2e3TScaid5QNnhzw1p9gbI+TWZASfoY/
g8DXZSM8HDQ4as+S8NBo7tnJM3ceXALhYNRb1nYWlYhsdHXg0u7rpGdjwM7O0ufH
9P6EvzFlmZGMqTukLDme2sRA4zo4xaw9ZN7zONmWwLpqcth/SJ4p2sM0y5Y4IANM
P/cNo7+4FWEvHVud0+nT2OsQuBNzuMPGLzkYTqbg2FLgR/UB3qTNp8XbCn+nj0uC
/5oAimmhanC8SSEDn4mYBy41XkKDmXluRSKo5VkltENHR+ukBlIkEXQlVxiokizq
fUMSdus7jBeqt4Ro05FK/D2SLrPAUqBVWwhiT7jl93QphMLwCYxtJaM2wshqoA9n
6XZOEPu0vameC5I5SPuLSETn73JnrAiZCDd7X5No1WLe6t63BMlCRLpL0U/9+yyP
hZUp3V7vlNrS9Gno3IIvV0sW6embzzvmCZIhit3HIZ0dGGH+g2UYEsfBsYw54hxk
/rmDaYiT3jZ2QKTGGedWtzEZlDkXOCGKM78NN5lIV/a/jM1JoARNHKqNH2Jvl0tu
FwqeiJGFktXMry3g12i4YzXAyA4OOOIaT79ZbJH+khdOQ8E62U54XTRw+9u2PX40
8CerSq5RsG3eGfZq2QuUk+gulFub/Y93vvhtrLGHf9/FSQEOK3xo3yJRG8W/vk63
7fJ03SX2ws82ijiA3YSeMlLAD9+1+90M6nUqXol/bhZNNRSU2gI2Jw13r3yWo+To
p4Gnj235qqKT+qOptKW7TsLjgStaR2PWgY92Dc+tOTlbHH+2whIbDVPy83/2jFOF
S9yqXQn8m4dU2YqCKAymFt2V88JW1uxAORPx1M0r7RFxkx3fdQKhRAcElhCwuz53
blN2e/hTvv8Fv45QwtWKVaZCHeEynosukKiCuzoQjsO2q7gcKi+SfrxejQ/6i+ep
wAqXkDIXuBnUSz8hFsDP6Fndxi/3LulB6l7jJ6BAMEWMyjQnhekY8eZHtLwRJa3K
xl3p5s0phgf4vUgPK4YkYPAFvjTWtqKqsBX2AkfYrUz+3Ddd97DdeJv0G2aK3sbx
9+kM144L6VFcg4h8SFjVeeeo+SXpKiY54g+rI/F/iCs42hyOPxwvPFmcGlDRhLda
I6elNQa689UAKIpXUu7B98NUIQDJkRnrFOH497+VFa3A+KQ6ty6Ma6vrWbPnUjnp
RUZAZLC5vKcSEBq3VkYjNWQGukqB5jETYDBR2Kk5LZ40uVJobBzcyp27U8i7nGZ9
C9edQUoXwo97rEa/mwWEeh/hJrHgzZ6ynQjaiMwNlvoG58cvqk/d+lxIPKnojZzz
+Rrv1rb8oWn1HDbOAQ4HnwQpBp95W2YipA4ck2cCEiO+BbfG80B2niTa1nz5ByZU
ZU/qHP7YVc0zFVTgDsyIvnfA2r12gYdKJcBi9h5SfA5mLtpMVOf+tRZNKRbtQ/Eg
lNvsFEPMRRxqT75CMGn39SZTt9E1bE9N2IlSdNEjFR6mPiccjaBzk5JIabcHeIC4
b1E6stV+0vq4nWHrbPIxv7Yhb7giMVQboVC6bSY1EwAPaXxd2aE9xnvFxWdV5b1c
L1zLJBe4pnZc6GPHhSaBO0v9lqD2mSBbZd5vlRFzbt6uR+yMoomg6L7neMNFsKas
Gis0nlG2QgBErAjx17sIg+94D9mPEyjgJcjuX4ctL/UIpEQXou+wVEY9D0/LhWB0
KJfq2E+maJsKQwOVjFKI4TbMyHUOzTiDf/IvjE924Jfj7tRvQY7fIKRQ3R5Bd6hw
8UbwyeTCvqmhwZpIoB7sUbcKv9DRPYmqWjsHk5qDVb7z21kM5tbDInv7ikt/POft
edG0qUT7ZSfUfYQknrsqVuZfaUIj61cPqRxEMGzPy1bHdndbRPMg5v0T+Vov1Z4a
8yHlSXCsjFBXmgQM5oD3L5nnwnE1nGG7El6hQ7uDgPl4V8V7bLvW1gUk4WbpL67o
FS7hgWhkbZ6DAtKuQ2uFz+kdrFpZFE62BGGSN1hUi9KWifmhQknvdibsmp8hvVAK
+ANIY26jFi+J0/E6R+QYXh5sa8YHjmugVuNXAouirHS+YLEga8s5FykzGAzIm8PS
EHjMRE0MuZ/qjWMdSsCA3I/wYsQYh9T2PK9GdYPewJ5UDFaS5r4a6KeLG9xF/S4Q
7TCzWqgdeyfO9+KzT2WLd7U6/OgfrxxSNAipql5fRMeqAhFYDqOpMBbaAZr8lwKm
AihwqfIKMjrntGyj9/3Xwo+bnaxPmZ7g/4QgyTh6stWXZNrYaaPOSoNNShWIowU6
7NhLu0edkViRYBLc4Nik1FdcbQgtxUGq9f9Ar2848KrPI0x1TeweKGFmjNP2myqj
QzLiy6k7H7HD3qguw4hyLdryGfJCkI1hc4mXs51KQmWNHH0KVX3mig7IVcuKB8G/
v58HPvmFqCmjAR0CYaEcppFlZK1LG0ONm+JFEH7hTbZN8MgIKLuKYdT5tWoear9O
SPhliG45FIaehrknWjLmOgg+of9OAyOIQgiJ3GQT4EIfKdKHdOylGt57Lby0nucu
hsiLE2EwvBdPztU1zLvOui4lScQ+fgDNtOZQaLsKrrVSTF3c6oTN+maizpELx5wT
pvNTAnxEJw1FzFX/r0fJ1S238zHPeA0Xl2wD2NpDseR0QMDTLZZN0XZyCOa9KSqC
M7eo29fnXlu0XIGZOw3qvC4ZxAdIDKnzSYF89IQp7bRufgTxXa8LVLMRlk4YTqjR
z8ytx/grCazu8QsvAK7TJ0e1c8vKUd5dEg77l9ZldCbr4SikqGg8B126v5AZclD1
x1CLjT9bppheSqdHR3SXOMVfZDfRXgE+q281EaNA3KS1u/EybhED0wr+fwhYPvnl
hcGqf+r39XX8VVQJi0ordUfPlXsy6fkLx1yv8OvUpkCVJdejSspsVfruQrxdR8MY
sGYn5ffJAmqHkQ4CzqJR35BI64W2/4M/67bS95CbN9QuCsO4i76uQT7xQMHmtgwK
EIzGgl1axPpZKK5uD0g5j9jTDk91xMWiXdgf3FT2WSZQeIszMEt1OX1jsH84Zgku
Lg6+WvkfO0tz2o6+ApAm0dJ1gG8iRzzcBDI3oZNnQ+tr9cCNg/H+KFIBDsDUqTmw
qVWGIr/eQ3IGmJtlVZJYr1i1BOYEKog3mDRlm+bcMzuSR9x4tdXUJxouUii3RUSz
1SoZ0djYBGce6nOBCW1e4CXNvWOHxLI0QGORZT/OaZ7t9PYyki608VBhGoUt2aJs
XMWaY4h/ODSbisGb9KxZrGX1sg5Bs4Kpsl9VH0mqntN3Q26rzfM7L/z5vWUJjszk
PDV3rTqvh3DIa92y4+FuHfPKbfvrGaCzv/9Odzvr1yiWfrd13dfZGbVfNMNFKHgI
Iyunu03jl18q5v+nLr0lFCNdun9pf/QQthFxhebRKxXi1lqeQsqm5/mkS9nvCzxo
r6P3xhztvvldwiKhc5QhO3pVs5M9EbWwvu9798eNPuN2chXaOPKUXiFSHMWpAqp7
hRBnBXqF7MCUzWTIg2QCBpNOom3kvjhqbGA17URuy3HiIuiL3fH6JrdI9NrpoGLB
ajUzcFwQKoPRiB4GFHN+4yfkYQOiJCPaaMFGWwn2p/sJsB1NnZ6cfbduPzVRKfTi
HpzRv2VLxCcKKLfSoYEMuRymaj7hQtxB74Ril9OOKKbT40w4AzxJN7Nx3Xu0cjgz
72v0RiHv1EBYFBi4XD/g8+wi1PVcw1xQFNyOaoIWrCNGZ3PMKrTJQMp8Z/0NzudX
7Sq1CrMqVJlc329i/3KcHIBwxzH9+vbPIQpgiNpyWmwYitfKN9dolFMbUFPZEWsi
E122Y8zjiZHjHPjyHrEf9dEclo/s1nCLAEs2fjOZcRn3e+v6KYRRZmOV7ojiXnP+
JQXbqzR6wT+Bv79+9sKIzh/ty6u6ZeJZ4csgsAn7DIhWsWdx2WPIsY8cScN0RwaH
T4g4qGqRcQe9Rzx2+trxBGG6y0ExYpZ/MV32ftExpto/AcraOEx7Ymj2skaWCOlz
Dathc9YeXq8JUH5mWxBO0UY4+Jqk2l+0TjVWwyIxNvxYcXDU1G8f+TUggvvukmvH
MT8POfqGeKUKqPUJzL5x2e0UCh9E7BEEG6JDjDfMFaIwXRCMmiPxpxrXUO6myUcu
SJHcw7Zkuyy7uyAxkuUZzV/1vn4tr4anqO0rwkpCho3fm0KOVoWfEmtfFCYhYOzE
5r62IbWyj+nw/ZoedswRD+477IBcASQYMmTri9YaLW+nkAEXOipZSym/91j0t0e3
gIx1yz/WKg2dIBb6dFSZVLcNvfhhTwZF3biEF7SDBHjZLzA/sDzCXoGhOlyXsmm1
2bv3MvWpYOBUZ74pvyc54eKKAoPia/NqVPa++cSTxEz9+jzSnosCb5KehW9gONqA
DzQR3Pw82XLtSptnAmWKMoaF+E8AHDcudKnfEvVbz+SvNrOUedjEBkQ7nlIMWbNp
B/Jct9cu9DhnEwT8tHu7y3w3nx+vysuWw0CS/T2URMIG3lrC+AkUplt8/g9ZELg4
nD9VPiPB20UWybyAE7IeNszzWfKJpxqWyCWYfNSkkQOCFUAWoNUaVET/0tHVTnoH
Ps75tqk6fy7dFM6S35SkEx5HI6mBkNNbRVWyaewDXIBUqBH109DdLDm6DONLs6a9
IXe/+CroIEdUKxJlBagilkxDzX0nDvuXsA0MaAmR2jMFmyzN+DlYKjw5jBCwl1sM
q7L1SGpsyVOWPjWGY8qbnevqj2AXyODJrgkx+bxmlcMu00fGBvekhFzdJaBIZM04
rRC3dn0ul1xuf3xGNECExCJaYViKCj2TdpumLbGzWZY3FH7rrqVTkh/KVtTLl/u+
ieHGrTA9uHzDqz8kHIR1vkqTSGyX80gPnpVFjYKPWhAFtA0mwM0X2kNMxi+VGZzy
2zUODHPRUuuTdmJFTKKbSXW28gTvk0UP9l46NEIJtiQ3RcY48K9c2Gnq4iSrXV29
0gBfqk2vm2Wq1NawzpI1C9OEPNumSgMptk2kZwuwHhIzuWb0tAvCIaTOcn7ZQ+NV
YOp3GR2zARQRa+WvjnHSSFJvxB5V58Tyj+K7iYjsijQWZKtZp8a2GaTIpx4eQOmE
uY37czAfcA4YuRTaBd0k8FSNa/4QtRxf7C4yxAjv0I/XPeyCwRTh7bffnxg6OgiV
Xt5diJ4BuQ9CVCvSMTsWOJVhCXpMgi7BYwGddNjyiYd9aOmJrwO5Ou6b2FKdjXxO
WKOehT2EWO3T8uoEN15PWa3+L6xI4aK3aWV78yd2RQOf5aIzohg8HnJORDFegdk3
P51Iw3FRJBizfsg6WyfixeozRFOUX2TszJrcDeUtjp2H7rW+wbDB533zfK4C/r54
FTrbdhnEjeX0LDZIFfJR4/OX7TMIiQaZ/J2EKTx3+l2ZM1JCVK0oCBPNhnPrDklc
Ob+XgOToXQRX7U18DhZIw28fr4UOFtX5hDdU+AIJKwvB/CMhI9JRWGhE+gHCm0MG
nAfB6LoPNb69sSHeH0R4bG7byKKUOVzkwV8s8xyL+coNTKayMNbPobcTTGP1BCB1
fBHlC2pLyAmpRNiRimbIKZ4bWxPn7Z5JpXpCtfWy/cMnFGU4EFdeXjhZ4yebptAq
C5xeAwsPqHU45yD91BoxyEb3uKw1FXLZvyXlbAuBgWmS+36n1Lp/a4+ZSue9STmq
i9vF742REjfTdngpPR8GGyy9nXyhYSWVnMTqvB6Af+Son0HdGaNqfXdC7uNyt5CR
vvi72VKjVTWDIIQUMsixNrXuVx/np2Hr8wB8JeJf/mpD6hWHajkumBg0HaK4jtyN
PMNLfM4Fhwy/aP8Spxen56DhcaOYOEhgdRlL/twQeF7n1kZ6WcwwnJEE8RFu7OnP
vIuTrYnky+AJDekhSkntiP0dPGMfzS5nnj2o54bJCoUmf6bcVJyUuQhOm7mVsFdh
XTyNDcSbryEP+tVCkp+k8zNpnXCljyuQuAf3ggMfrH56GWBioe5wLrW26nIE5c/I
9qkZHrG8mHVNvxYyUVJglTJ7qdZLhTgfuwpWkiaOnvZUrodRx6CpgiMoRancpKRG
o3yCEHQdxw/pA6GzWcOMlANi6liYVSrdMYwFxJp1yF7ypaLqrM9G7darSfIQYk1F
M+I59P12fpjeQvccL7rtoCV722SxYygffw9jLYBffnaAjKYnBM2zB/rom/OG1lZo
UIq5p8S2lkQ0Z6Tkl5TbZtosdRp44DNKyfr0BfZiEjd0bEUc8o5PUQOI2CbMn5WF
gkc4zciroq7IY7P0En6vOOMFM4GKyGkxEBqin7IUe0zW0B4MhGNQNbQi/lT0XeFF
o/bwOmf8pleVP6sdqpyGVzb9i3YCFYk/MQoQPlaDTIrqF0oKJSAZq5n65bu5fZjc
nHZfCQ/2LuIXMqQ8dbKsLolXnCtEy46WadYnymgfE4b/DvO4EakSw77g7s1nU75l
94xqwP3SZNFyDNkoXcGlb1PqBRASnv/uj2egKnFD6mmkzgXuA6uwH3ZJSM9NUJ9X
iWjuJ6cyThLV8y14AWSFmUiy1T1lDhAVyi2Xx+D4oDRde0DdnR9bxutajWHsKAEF
Da8B1uNEOrZeJO5/RvWRSUnPFf+DPSDTHQTQRR0n1F4JZmdWml0qtM7VbJdaU67W
3wTRw1VoxTrVMuZ+O7gm5WfYcy2aC+ShgtgyFbcTbgU1EohPJGhCoJPmqmgoaTUc
4o57nWeJGkP65KRw2hthajhh1oAdiIwcd7TAvgosKfvozkZAywIPlEeqkMgcKplI
7HewyV4QS22IOIVfYS2W/ZXGzFav4XZiC9uIe0Q4pbK8A96UV0G55k/uoPM5XnHv
DTvhbZP7qIbKaqI/BbLZ/N9L683h+3wPqyLd9HYQE+yTw/+mqsZR88iJMxEriIV/
2Y6Qz2+gA57rz3qkmvy6s3yGMbrCxiV/O+j5YoieQXp3Top06RE3yhfsnMxcBj1L
s1ouEIYHsnrd+cdltcLtOtV67Vs7lz8qwU3Cnm3yAeuGG5uejXrV41AqWlqxSfg5
4IHajB+2HAJYMtIoR5jpC+Jr8yuM+JXSDLg3TWlrXu0OU07qTqU5wayb/RJVIJj0
2EiZGz4EU/emqNMi2pGK5qORaC/Cy7trhs0GRdkaWUPhdQUdmZZz7R+RwKK8cqKw
0UJri4PM/vRBvheOkqgp2jMwQU/y7DXfbGkFcBTEOHRvBTPuRy6pnJE5N+7Ii99O
xVkRLjj5Na2I04DIdwzjOTKSaebskJ6jtGPWrVbGTYK6+5wFqEd3W63Z0HVKJu9S
R+Cjk6ndmnhb9gGiQha+XLfN6wZFlE4o/K7zWJP2W7YQLYX5ec/O05wCncr2uSGg
Xlva7Kh/qxr2++chdLmcWS5FRQK8C31hZbUQllB7TJD17URLkMQBmTpwe847Q4J+
rW3mZRxLlG0GUVX3csmRR/vkJMKSWDHbiHsYguPKnNX81e35mRoxIX+o9pfXo/uG
QnHoLstNBo/Mg1ixti1687tY+rwe5PeWP08v2ktd1fRXj5EIeYsKDTWHYO+ZSZQ8
9fDOf15lD5dGWpV8Eo69Sk03zL7kFuoT2E5qvYUyBlG8zOe7NetdmPxKFJQYOcJ7
ZdVTEDQ6dStsU3Vr637jsvQ5UpB4SI6DD9aSzkD4VzldhjHe8gUh7zdBIoeYZ3yR
lgFFUW8AQZsrABbWxsEq5YlCDbY4Ys+mnZa4elDnwsF/+gzbffGnE8iTFcz6uvxZ
+WjIprFbFYPOJkz6THI+2dCOjRDAi6rSm5jgmSmtUtLpkoC6Pqv/Gv39YUo32ry4
eDsr8dbFxXRcHhi0Rv2W2uKAFI9sKIg06iXmdnasQGDXg6E7m/CIaVRbdiEb4OGh
KgohLkNMUUi5PuwXESG96A/D/l75Oj8AXhZ5CKxUwtWLGqH9GoXlEaFiK5lHeNYp
XTBNglrsKUH1dXO9oeE+FeCCa4Z+Zlnhpqxo20EtB/5h/mbnG1GzoSJeW2kNZp6G
JhcJqVSj8ZQPKqKOhDTF1PAUaqEtpu1naT89whylYUTKSb/4l/0yrk+hQ/FdWXGs
TE5gVlKJjWvLuEDLdNtbxfedIJl/+QqglXy2sPlJr+Jq5QlFDBWZCVeo2XETXulE
OuW5r5qIRbxKQIm6xNjLYddXfv1/dhunb4EbnoRQVCb8s0ru87+hX7cpTULChG0j
mMHJcK5TYr3ADcBfEIRICPxyACcyh5dL08Wd8AD/zJGTC1wgIcGTkPi+iutPPCoP
JvDIZZnMPfPkmg0BqONIhJfKlIfh/foDxAZdHX4K3DHXRnDW3kAcydSdbnrSrUV/
HF9FI8zhOrMhoTOdci2cJfbs1n5o6Jx4zJ56sX3vFk07zcUbmDGhbrXai4njgf3B
/e5OeQh2bqdp8enoT/IvwF+SY03aaBrTpxw+YlpOJ7ySAaotCXGlsjaHhBmhKqMe
Ys339wyNfpQ3NHZBkdtrKYA7aWg30EA5VISgmNdXGpW6SDu70fGQHaU5oSBk5ecB
1F4w9QbIn2wlVmf4rLxb6iRQa/hDrZflURVqRnTJpuc1tiK4T0cKwPuwtkRWQgqC
WqZt+Q896VsQOCkfMX7LXLrev4MfAtzmLydgIrnz87JNn4cU3umOyaoqSXIQY0cb
JRcM9NTj1ldTnAWiA0NNDUMR52lxEkBU1QalGgsW5udX0ollaebQV+Vwmb80wLWa
Wv7GXnXgVkjttdKYzYUVUoIs2PoyH44zXNRBftqOQutM7FGqjZc8AiMkPhP7+P5r
wOoY/GC4diVumUJ8vNxYxBcMCFH2YXBVCCdd3dfIaBDWuUaI0e8Gy3zoMSej6GA6
sZzffNU9sXYF9opDPTY4UbE1z6/B2z7y0DhnUbpYdIgyBAKYSOwnNm+5zvsCjE3f
3/V/gy7whwSyJy1fBg+TekaSqKFKx2D/k3B+Nzv8mzsHrUbhHxfIKdET1CNCgey9
XzcNFX83IxJ9Eku6hb2fUtCdxUE0/sMNn+erSna/rU1wFTKuJijN4fU621Z3LVic
11gV2jR7Bh2EAW1kPSLHVNDSRKiPMvjDXIJUl7l1kvVpDkCOxpJ32BWXfVWv2nxe
lpO5i0FBNpMqJBV+cbrTxXnU3kYSn2+HfKp+3dj7Wo2fx1g6c1tu7Jef13jXyfqV
+UXACuKQue2ndwZeN1qBBY/vGAdR/r2rPlC54mj5JdfmHjp8NRHq/UOVCT5rKqb+
xjT4peUVqDE/1s6oUc4ekaQRORkAr3b14Pom/Od089Qp99Q1/8B45mvTZW53/9l4
bXzvdpT5T/pn42ztuiA9S8Ss1tmWSudOpTqzDjybGKyeh3MRbAl5gMohLhCQ/t32
MI445+O8bixs/ST8E+Z/+QsGwt6TMmfubJedt8vCpboeMqIbOt+aDkBjujIqJHEf
33qwTH+Toqvw/0FxGRhDe+IU3yJ8/+JUBMFRu/g2SXhV/X0ze4j8lbPat2p39Jc4
11dTpS1bVLynD2sZS9J2ZJA9X4UB8LXfxCr+tAYnlp+95mtSFSKgs0yks09/rcRq
pBDQ5pqZVPGXHfB3WfxOJt5l4PC4+TcwmblXfLHHPlQ9U9u+pFfxLqdFvFCBP82G
f3CE8rnLulMHGh6RbyqkEgqLaUZuwQqdWc5pI6Mt1fAoauPl+jpCSmi+n/bgXwqY
Bw0ckqa77MTHxrExYuPSBR3BA8yHfnybb3QLzmwoviMqKANC69voPFynjDdOC26e
T92xulxQ/ZLUdlqP2ZRMgwXnjC50s9JFjpyoQFIvel68vqxBC8qQl6gH5Wcg6VaX
2E5SfaZjkkFI6B9cynZRef9fV4HdV2m0QD050cBGr3US5Nutv29ffsNQOx6vCcfk
tLA0CEItR4hf0ERQ7Tdrv3v/cSByNGQIxEt/NYzsxMceCShTf8w+faKOxw5/pEKh
CKU/QE0Ceb69D3X1IILzxrPik5CkEt5Dgr2LVDQywW+uC928RXIPN63TRTfLbjgl
x9gUrRfrIcHgPRM7rMr6BtBCByCNDJRsLTUNsghKkEmnCWUzRU7taqEjqfnzvj4o
FbMjWrkKq8eQeVHu5SJ1In8rHittXGN+xX5sRU1n8cEWE7K6HJwXE+YlQjfPyiOm
MGL2v8F6SH+/5/+MESwT7lk4Uo/I3cgg7kDbHVIwokb1fBYFEhnBxciDaJDzxvlA
71JIP2QZmjJJWiCisYRIwdng7dqlirMQAMscZBBbwdoiF35tYA61Nl37atKnkQnL
culaHZc8gFo2jLt76vGPyU/+M6/cZ58M5DRQOAtUdDLENX9GH0xnHc3GCoRw7f26
OPg2DE6YN+tWIi8S/D4fSGqSfmpkeLiIVr8HS4NwwWVd14o9ONY3le9Xo7RJy5h5
nxhhtG+p3iQDfS2hW3Lgv9GZEvX8BFViGtsH096GJaJpUBEI3PeuhRfsLXvb7GXa
gp7qZZ6obTxxuwVjt92SfXnrVqJ55/7NrgEoBAucAMFjKXWdwRzEk1+39ZYMUkAR
W65wrnjG6czrgHJ6pHBm3iVaJVD4g/ePob85cngCdYeVCXgIJii64Aha9/WAu9oA
BkXpFZRmUEZGBEHQO4bHBsWaSF5+oMu6dNWFzECJKhHJydD2vlEoLjTXC+/TVj9h
bsg1KGmg7k5KC1Z4lnwGQCMXQPI6QzM3bgdID/dphZ88ONqBJ6Lsi+hlUqEWj4es
pajvRjFIWlIK5t4vwJXGDUdhipNkQajZxVMPcGV/IARuqQ474NX5aCKzlx4BdbPE
54TXAXQECctSJx815cLpCW6UzABAlQRSls+NyxELBsuT+juJUrg6Kx5bbvg3MUfW
FkfP2Rzp8SdOoBe5VCU7cIWctryrI9nUvB4JDg81aaEAymcfp3AMCaKuZQzWV+XZ
zyRhZJKwRbuqK7OEz1Q69bDP9XoRWNX+JcVqIY71eeqwR2/5Vnct0zaGFUv7GmRh
qUaq9LpCMwM1x8nuVgBg0WBNd+xbnTOtiaRo45bf6hsena97SvZvGQnH6vqRttRI
aM0Y3589I1+A878T+LcDqi1nhti3aHPhyraM24YpfffuJI4S7yE26TDra8J9oQX1
aY9PE9Qmliv9l9p1iBjFif+e+EVxFh7CYmc4ve1fDhJAqEATDURkWZB9+5++P0Df
68I6gFSIVLQh1MKVTt+26r8vYViQvNmiJbvkRG8gakf69yp1kkH9GH4h53iXz12g
i1KttEqrEZietpkd2DruaDHfF3zEeazsZWDkFxk3moXZwXNOtGor5QMWMBEXDVaV
mDjIy/MCy5QlFHvxz9I/88APZrdwJpofmaJ2FYPmo4qnePHtuQV/m2niX1WTiTck
V+Xc/4YAe18Ry8m2SKbyhpeK5ECHugqNcoQI/j6QE+i4vb3DJoGIPd3l8ytNKhOM
7QNStONTFtz/1dAizTDCezHuLpm2PDHu4Xky2uKRQfnw0dXrkTli2pEIvTilgNjF
99POEF75As3qZKsd8bxHbQuyzc3EzO0kqSxILEaLk0S7E4F0a30XBgg9VQrXIK8Q
VJm+SJFqOTZLJE69/7tVc1t3EB1uz3wxquGT2BD/8RANUoMrMFnaFC1050UqNBuU
RK/1Pd4WFQsWmafgWsofsU/P2LTThYnAePK1/Rmxj9s4ckbgomUICMflc6qGnuRL
fkEfD7ELR/xq0srtdfZjn5tSjzBg1boK8D6K0n4y3bA1ui6gc2Tj9dWRhS2kcw+3
OIt8Kdft5qOYQyCmkT6J49vcfSmYkGCs4r5nESHP88dYKdD/eldahQv3cjQ6s3d8
YdwOPhmmoPmdutflJP2A0RoAsKsYJGcqrOEfDEWNUmO9fH2xhxVZfzqLHKwLDkG2
WPnQa18Fst/v8Q6VT8RYIkqEsxN478I8OYmDfOhatvG0DaoDVPJmOiv7UI6W8LcD
2mCo0RU4vkz0C6jnvK/7sh3QzhUdqFs76PjTeJoYwQRAxdOPBubxngjE8MtKXFBJ
eaLKTtCZWKCaAkwjOb3c2MkMmFzAmMGquvAykx9wee3XjptUS+hngGx+Wr4Y7v+3
uzXlYCcFvS1ced8eGBZ7L/l6UrlyiZCeCBnBu3BZaRaPXqCwDvMYmagtHTUXOpgH
DwyBvCkXlPG9iTr6QEVcsqYPN6wP7+tXjM+S/akQhGgY+jV+wPapQrfzR2zK0QdH
2JxeExa8yJQLjW0zgt4aNsrhr6BqsgZUpvo2a5oa5i6ZQJxwDlLLJQ2vzmT1YbWe
BjtskO2ZCSndRJptaixu6G16YjtCX841Tui1PrK2EPEJVNRRT5gN+FwlyQx6Xw+0
PCSyVVbM2tvrqAPs8gJtbV/iV6+8S8B3cDYfo4PpJpOXTqgRTrS32vEbzlLPDZ5I
b6XsyEYCfb5cpvBb66UQtBX9xAD1bjdSF3OG1bta5AE9Rz3WBBlmYfxidnB2q6Rj
uCdjkvL29mk7wbWSuoOlfWgYb7yKKDEwDGkcSG+6WoCgrDpR5jCfbNwfhzVd0krd
mCAfhzaQ8gzdfTjjS/8RVN7NBnIzVPTG8+9tEWowZ9cKwWl9/QN0ebEjXF6VbSjS
dSmVjn3BQI3QO7uUtibWG+X4QHiwlY+fBpnh7l2bKU/49ipHYmsxBuwE5MmEi7t+
IVyQUvz3qqHIy4nBbOPNxhmeBgIkiBKlvGa1qE/itZbUrdwWP/IEFiAiYUR2qumz
GR3LILseFWZZus3Oyl6ofkUMBP3gb5KpwIFp9ped3Ll92CnHmFAIGYvUuy99JdyT
fd+SNmVUrTmckeqaQ+C7W+G2t/bqn3ZzOHgmf6FHj+uoBfnaKVip6R/qut4454Kl
4pZ380vWKDTy8ENm8KXLhdaA81OpQCFUuQ14K93LeeGFvIM95D8LrZUq/vV6vfGk
SF3jfXNcxvYrDiSApjqKM8uQEXqt1fKqZPYAbmunwPj/jK+uPr7QnrdPPAee52hB
mC5EfvMTYmmKxhrRcNCP/KzRbw+ZB2RitBECI4knFT2ns/bg2yM4Zn5tEZReCA9s
SePqE/49PjDBxXjqituxAQNE5E8tlUQ+/gl3h1JyiIubqM6iq6cIgzX135gXqg5P
1DwGoDGXOTATaZ1tkHDHo162iEkkJun8o0lqJEMhbN6Mf9cAZWepMZeAWqziJzTj
ZLUk8BtGQ42vfUHbogq9RWPhdADocMRPyuWPEW7ZRhHll5vZvHr/CtlPmATF4LUx
m00t01Ml3vot0CTzaHBGnCGuFEMkE0sv8S4sXmBNoeVvghtm/lXDsCC7jafBhr1a
1cfya/p090+7+S6v5QGJ9QjJxf6ONLx4xjPRaxc5pQejl8nyayV1flyDnk8yWaaL
ZaXSOeT6RgEfq8Z1m5ZBYxOKJky0wsdOeCNS5m5hl8Zdp9BDFFfZ022nQWTHlLeT
ucoJRzPFiP4zaf7dLjfVWX6Q6nTKYhNZBrgescTtT8ol4Mx+546mYuAlUFhLAUtG
ckZe50K9pT7ZAuoRHQDJuQKDOM3B5OGAdyx5Q2qEV8yFIYJMUzsyMQ0+r2F9qj76
GORHPf7JLqKrm6du8NmwP3yZWlDiwTU63BPlUKmFUCIXuiKfX2srD/1mhizLQvXz
vpBy+MeAMw48J3PZKHdHq/ZZads/ypqAEhVA6e6SE4W+Egd6rbf8L1dxcX0hokYw
PjHn8hIbizZ5xjYw18lJMG6V/GHJafDi4QgVVwqu6PNQ4DCN8wU0YiP6NHXu4oxr
+mjuufhXxQ2uhmQ00zLLd4w2X9veCV344MEO0xGFPBEgFcd4MCx7L2+sEGQQMDnV
YqfjxdZ+wQpZLRInubuRrn2HuFAhTnDFgBDOZPa3ij9sbUw7775+RQNlp/HudQVD
YT6u7A3rGUDTzSjijctm4ifS1u1Rs3pd4vkvyVfv4C5/5CAL22XsrA629kUC83HV
nWJHCwz0TXJxYk3xKmcK4r6PJdvzU7tRb8i3scZQIaxEbBXT3r6ij5ZkrAr3cR1a
Un+slz2gjLUFQF2cYra6VFBuh4Z/+wTkUNgZSz95KRPdtcWOTe6kNytvJ0CiHwHr
gGHT+OW2XWHT/CZAyqCiT05GfQNtAuTXNJ3YPmCzvGAtZXCGXeLCU5ccg+cZ54xe
4qjYO8/Uy8qOHEdW8UKMNDYoEBR87fzsCFb4ME5FEylxOefGwhlc9UklOAK+2DA5
4SiWu9z5nPXdYftCh23XWO/zlOf4ZvL+oxj8Fu0Z4rRR8l7AFgLbmxi/IWbrEblT
OaVGZvmRvd0fBhdzcPsBBvvc0tMsKD3s8UupuVKlRHfCbl4nxRfsEieASgZoG/ky
YxBn7dGcVtSEeUmxCF3cfLAbdk2rbtBrG6eDKNf4ZD3T3SoF1sVZL9gMai3XesTy
e40AHzdFAuPJP58Ii/MNpMBq9gaqwJzpRU9a/ItVqtWr4vnCqe7SLuuf+uzgRCO4
JuVRIN9WMb3zSjn5xGKWiVe/YxW6NV9lGzqQY24EGz7JHXIZyaNvAgAGLFScCVfl
eKC+x6vHTEYBHiABFpJVUVqlK+3n5l/Ij4x/COAaFWPTjB7g0BpjTJRCj+53aqfY
n53SKY7QI/h+6TNEHvOL27Xd2ECGt/y7/CMDzZ8QX4KQYLnHX3S8yNXYEq4WGWtF
zyCdgVPCNwC03NlAYOrPu/trhcr61j+KCNap7MG4N/VZb+OIAbJiGESMwCU2X61/
gUCkQcc+TbJdBj+eamBQYf6JyfST67bbkNOELyZB2ERYCW3rRF4OS3m/UQGvYOxJ
RWcdZdpJF57AU5j/B47HnHqaT5BzTK8MSSvGoaTz5taknKPgZ3lPa1mt9w77HF9m
JB+oGCYRjpcI9E7C924rWYMYX/pwy43UIdvrOWElCMqhTxY0SAJm6To0mGJa7DQt
ZGIKRVcT6d5bDH0IzuVffVmcUUMpivSJPsaY5U9FQqEDIgyzyeGCHJTtnytSmYCB
5+3JnvqpR8QXVFFYTavPH+HovotBcQhArWExrGbb3YgGyx2c1tGJ8fHz8fEai8U4
nlYI2Kz6FsN6O5jWlNHVw6gd8m/jXjIF3ss6d6Xl9U9yV8N6YDA/C3qbOoSsgMYs
77Y5mkvWkgXyBWyg9lY5iTFPf/W0QZEX0pDWFZKi9+zee7HKVs9B0c61KknbATXh
X7g1w35yCFiJ7do3qyMy+PQEt2P6xBNrcAneH6mJmu44dqW1dQEOHShCxZCW7x8p
RkOIh8bX0hYl7YGRzRQAOH+ca2oR8do5HYb7re6yr8MnhopDVk9fuQkonaeNTj7g
mJ0bxPHRxwru9paekEjqJRLh1SerqIa0ehek8QDNAmK22chybx9C2Tpa2bTP1RF9
GZgs0HGFL+Ov4Swqz81t12pJtEsaKh53RnX4oBBdYPN3+PoYXFKaydjYO+6r/nIL
QueTUxkUyPsi6pC0Dc4RBfeyCvuTt0kZBDuvWHokLwSkw5+dT0f2m/eeeCG1uXxz
sjOlCgE/o1/IDKhjvJAYbATFpv98ogGlBs/HpN3ex359YLXvRcAwLeSyl/2ZDQfM
Lk2tG4iytrij4HbNfUMIZ1h4clohzKvnD7Pc/TXmts82c20SqdahmGW9/f3mX0w0
yMfOA41puSIsEAcWlc5JDoswCVS+Dr3yzthaWibAz3bf5RA0/koEU8ZHxgYaeZO9
/abCXbJnPhsxXSq3Hyl1dqDxZ2SfRVrLxUHTV6gH72BGDb+rp7ZFS8LGTgOe1AWQ
pKgPvA7uLwlo+Ao+LjlU6keMQtram1fx+zsRhdN9btSNeRkvVYaSjMC+hqCpJ3q1
QSGo3NfUXZNNZOJC9OC0+ayoCLYzjXV/aSjtinwjbtUaD30yp0aVvfUBB5NWBGUz
RkxVmx6kFMDu9kIdE5X32UBUlENNRueNZFTAabrHPQKIQ6j+4b2LCEZsnPjRAtra
1/ehooPh+wmS1j/a6lpGvs3avmteMsn6E4O4IXO5wPo7GsFIexqnGJi4sQWc7wBZ
bhBFiv9N/G63sOXdTczKRxZuT/RuMuKwFMvn76n6dEMCDURSRa6fJAlBLKoB0icV
JbDuLUgPzeMCTRfeRTg5R+OJacBXXOcsXaUFmdwAmUe5uHuWpXfil+zJERFmb0Bb
9Rq14EBluRgKkU9tzQdkID3P2/SU3beFXT/xZ8Vb5GXN4iC6xz31H3nTYipnsXV5
DurASwI/+tw74f5StS/c8EVs6nuL/vbShIvWP9DgTZWlNbGvRpsR63JOlcGFWWCf
ZVQfCD1tEoFoEGiPKWQRKw5Becd4K8ymWRWDaManRKIQfRMdoQsLugknCdySm74h
ZOXJa6pCdlKh3kpE3AYOKRktZsfc6xmlP+AmEva5Q5hMVpp8TN368lVhNHQqObr1
41bM8zi4G1HXTQ6F1zpENHlfQ9cOcnY8YWe+IBKfBSoFsvZ6oQxrxZeQzM84J2/Z
RfWXIjeKD316YTJqrNGCvHTeDDFpZirNx8q1neqr6XTyXm2jTqUFCHJzFpMMTBsk
AbmLJn55iZ7GVcDKinA4ZUVMCccoxRGC2JvJxQRsMCJ/OIK8YROYm7pXFTrqA7s+
V/tZ06vUDMeDzpNsLzFcLakVkph1rvGWidsyskErAI+/B0UzvaZWpoa6FNmN/7yp
hJTTeP+btuM9lfcfrNYLvDR/2dfgX5jjPA7rP46EWfSnMj3PdbOYe9DqB74IavGs
hnqOpMxsglIIt2RDXWAaWrvezqfPqYdg5MEp9HvX3ci+ibuoG1adeXtENGzizqDd
EwU/IBfK79qp6umzsEc7hbSnNPxIBB0YXZL172gQPToYAaspUaxMQrrT/6C3tpkq
wMiJ9OXMmbeKJOF5PyiePYKea5AaCbFHkWuL2XwiHPTMBlT0axUmwb9updb2aR9b
/HvJDIFUOoj1anR79nJCj3Mm1/R1IWls6kmDV/WlGIhq7AZGVCGrB1rECepPPeQQ
zwuGoKb4LxY7kgiU6b07QJwsk7NVeqrIjgBxtlZPwaNYvXlglPyzvh9WYCP3yyTT
aKsyGdpKxCd0vT71mqRip1twrhVvkaSNAT/7mx2OENCc5Fw/JBzVUekHPN7lgqKt
q4wPnCYacCntGT0TaYGmV7COk+g72O6xcOtEyjhPJSqljdT0MWCiID5D8l7BMB+u
tQKGnP0nyczEfnq+eP1v6PF/j1yODjjllAbgB5VEm8cyYU56sauEoSDMcV2oye0s
YY6VsE5+UraWyNFn+kXgFbYLid+wFtxT/sNqnI4yGlqZ+MifqV3QjHU+43FWcTkP
HSYaPVtL4uC9RME5ZQmGKafhr/V5W4eh68UJ+vRIwJkUgLEXn3nVXWOvDyn/pCFd
KfOhd+yBYoFfokWtuMilRSo9K5uM+VrvC99+Ij5Y4ZGE6dDqwNTlemenzzkoPNub
Zn32FSOn3KTIbwBwfTN5dse/Jr1vx8PQSfGko4Prgf+f8lRhH3Y+fUpoYB+OVo1W
2VGRp7kgJq37XEQ5bw4J7ecE5fH3WwZTyqOfz/BZNlikncmqobu4MIN/gpXCi0ua
a+vmxGPWMBVSxSXcwn6MmJ6sEXGgJgBFHyVHsdL5pOjuckrCjAqppkFejMs4wbeR
xds/w30Yh7wCsrdESNa3K8Jz5HesilHX8anHh/pNX+svBKO6OhO82yeMrN6XbQUn
snuLWQN1ItWlFypVzwM1I9dSGKeb8RxsNBtmaoUtl/MU1+2xMtM5mNDXB0j27i6X
TDcj+d2g+qqgfcka3+TpW2BDBEqC5VROfUkA4+MlEZbQdZF7VaMbW1xTOq+UJ5rZ
N7MtuMSSsmjnCS+/72VeOpjOfQXd/8/3lU5icMP3yfJXclbSFm3Tiicc9zg8LabK
enZLBzcIPvCnK7A24qq891X1euLGLOK7OFjTOsOAkt6Aud2VogGirKrg+9r3YyKk
w026Y4ttHsLbflVUm+do0zBN7l3dAy7aMGDZiSDIHtn4p9Gfo81YqCEE532xRMac
gaW5YmCMuGhOBduvGoCxbmvMUU6yTlmo0sEZksJisKlccwu1FRDhJsLRg6sq0wdu
LSsF2mBJmqnu7y3NNt2NNiVymSpBe01viuGGcuTXQflgtxLcFslfMDApMRcUWef0
n7CqMUotCT3whik/WfCynEhsGYk1Xei+SkYYaoygFruE9uPZfe90gSCwwmN9tWvH
OQzRMayeuYpoKKSGUDf1CIMOKEUSAyX0WBK01zx0zXKcsWfDtn45UQk8SQvR4Ype
0nTQDpYXPBI0LMK4R0rYo4I5Zij+TDfOSnwE1CCuad4HJ4XXMOnEOBVh3BbnQrIu
vQ6xSkbtV7ZxGzX86MK8wOMqT3k2f3PrevtGYMkuTAKzYY11dqtQ6FO1HCdekiUK
XX0/wr3PdcrUFakKb0e6khcaLq4e5x18XRRPAU8R1qLVaEUCysQR3ZQU85WFtvND
4AXggVyt/OTkiDKFEN/MwhgaPKM1nvOgGo62c4cqvkxfdVNfffPH+D0305L9pInX
unsnplCbn3a0loWrXQzlbI2DZ2/qobEZW7sbhORXCCmM5pQEP9zNS7ndoX6sTP76
s0VjoBnfU6ddlGwIJZ10f040SD0aRSrKubXc1xG8iAS+SIVSfL30KRGtARPX4E0F
SKF7M+38/7aRmFXN5Bv7ymm4lxEwwWaPhRVbrfBcnZpv8uPMrXfHpD5tOjDvL4+N
/oFHqft9kCexrGLmfRGOHl4ZsUGAxdpZr8h3WBe440fyqM9CVkYz9ZbejmUFkgwn
GJ+cHQxiYQeZ2clEZSBuG5ORrap2/n1FoBpoKjXFyqGxFHd9MNT/QraeYAZEpGIV
jpsJXJ7ZclYOSqrImMdnDJ4frC4Uwnp0KjujA9RZ1N8ANjsgas8ICQ0NmM2lwO5t
MBqaTvzO7FWAlvommip4Scyx0SvU+C7LOAxH2nlJmk43ylq3nfnIAooevceaH/vf
M+c1fJa+qdGKCY/nCtsch9nbxsuE25naNmjdzZvxmyQABGw2yUUA5d1dqCAAlovC
q7lCDf1YlfnXdUn+UBvPKe0V71CeGA6nkPkFyi6cA7wzqHeOltMpqXy0xXQb9b2P
kl9m9sBjff7zNHkSEIRfENNMl94bhila7hZWQjoq6NuyiKhO+W7PiSgWyW4ozRXy
bh+r4ZzGNUGwv8+bLIYaOsln9ha90bK4jw0QeLQQBXpLdjq00EdvtBOvMQDoX9mc
U72glGXXlEYONgLj/WyXijueKHjY6jXxdsXIiDHluCmSHLJ698hYUErn8XAMcgIj
yQ/azOsfxNIXdaaEhxvFUs0LsrDLjV6yNwjSuDkXFBW6U9D10PYwROFwlBhf9sgj
I6QsM9HyXZVZCUKVzqE6YxjNrJMNZfJbSBLm3DAqTyE5QmfRzJ7D7r4qtAeuP94x
cZSRzsMgiJzuuAb2q+RoxgHScP//q/XdKg8kv+TgQ68VvpOGbbMMeq6YrdnvkWGr
L/96pITCp/YG4Rlx5e/uPVE0njWHyeGHnkteU261oWuGvQyzhSAvZI5Fsc1xWS+5
AYdvVNIlkhhSzgrtwacd2/v6BHVPi5bpVHAx41Zxg4Fpj4tOEP2Il/Sg/moyB8US
PTuGCG1FnfWPy8SgwO/sC0Xue6FtTrGy5yeJj4Q+Vri5nSkOXlv/IBh5i+K1d0o1
BsMtHY07OpWyB67KTq4zN4WzGVSbzN2bzB8pcGpEmm+7KjygajJSm63UxACm+yqo
j0qCc5nOewTTKXRaA+fLHfW4GsZJafIEAsNconJdjjpMy1fIVZvpO5mAKFXiKCsd
55vEeGt7tXqwIeHgGBbQ9lDOCpxjcLDftIHNgYai7O89GvKSMAgbxGhEAm5atj7i
V0Cgg40XntH5MhgS66opyUGOGBvi8oncDzRMnsb6ThAf3N3I48sdjFw2cs5dtAIt
1e9hyH++3jy/CYGwSdly9T0/jZg7wUKZKdP1hoOX3l60QRu1QO1uDNSXrlEiOios
UFdbmyuJq+xtFseaJI5iabJG+HV00sV4UB3zI8TNjg4Ji53kQopnxxneoUJtlX3F
Eo/KSFJ9yWVsY5rRdqakcnxYC2ct550fg37lpAq5p9mPxLZMGDVy4MZsYUXaOi2U
YYpNRNOwKRvirn/e7Y6eK18Hwm93Iv9ngi4wam1IvHoXn871WIXySh4Tp9mqNwJW
xar+hvO/LjMqUEeYahv8cTMHq4JHrpYoh0eZa8VEJ0m83XvDJk71mdpIiCu1cYv7
uvyLjwhifZcjtw75M8t15Ozm8M2mkccwRoYkUv1epBl4AeJ2qAo7BmckQuAudo7D
Giu/sVCMxizFEelq5ho0UCihZpdQH8TXcj3ws43vtexeqxkSId6A6vKxdfYJBG3a
IrqQ+fcFJx4mBZETy8OIRI/CXzouFWVAGc5+JqdAdeiqwhmtjh3wNScQiSUb/I7C
V8griYc4o0B1HLLsupcr8P6g51kgSxvlQ2wHdPHRaiaUFKPe4p/QiQz1dlGKUzmY
F4OOLRc0u3SF//t9UXJxPmAP+setlhsjCr0rQvsD7p6EXa9D/enHqTRYZa0nCvYT
BZlqVg2PgUOkDfCCp5YPVUfNZy2HNbBWVAkoSs2rNuXUT25taArAPXTX/S9q2mWl
PxkAJnk4yh55+m6FVwG8t0uabXqjdZDg9KOWjzJ3MaTJMC9/2IkffKe7srvuOpek
ENd/fzSdWvHPK8zUsSAy0GeanQdkK07fC6A20C+vvXdz4MAYGHasU4atz15U4X6y
HvBgXoeINcU/hj5sjLJTgnS75hTnE2JOas0cGGLNp9h1zeKf7sQSZoem1XAiB91F
mLhrVGA0pKqlJkPeOF/haodhMpdfvQEiZi6vH6gl6oBr20UrIQuKTdUf+xmoWmpG
xAmRO34lmVgVgtGkqLt9yZaa3zzgrgVyvFgPNI+Nyv875IPSICjsWa/mIPY+naLS
25nn8JFb+BCMN1lAa02RSA+mzY69oKwxOFkeHoRlKuGoU4xbGcnp+mpechuKGcNm
Leu816eh4TvrdQtm0a726xTLq8CWM3ld1fjyIz2t7pVH7EnkQsWGZ9SO1xftcS8J
Ynw2p2K2dQczKstWEeuGPJu9LzFKrwDBfM+xltaLnOHLYq1eSB4ongZylPrTFRQW
Rlqrxpthw3g0R634owKZTSmXFG/yDFv4pcorzn8j0luUBBlJ5tKWjprvSJcKROfS
GIiEKrVn0zGm8z/nATUAOlRwDnQj9FdwQ73Wei9oIWgwDBa9Jjxg6LiVldRWBdkJ
yw2ke8tobw/tSsLVqnx0sWYx2owooSQSn+DtLvtpo0HvbjiDDUyEi7ftvVuRu1kf
E1pjv5ddiDJBfAD8PtBg9Mt1b1eEfakasoquTX0Um1ai+EW7SXi9WROMwcxAlwjC
kYMn1OR/zQ5jqO71SQkH/DFoNJ4NdwLNhWD4T/wdvU4aAGkf1paokaFco9bnOB//
pUEUjqQyPeb6r2JsIB7FtXg9fIXegAdatYvo1Qu5sbblu0FAffbIbaKzBYtatfCR
cmk2A/3yKPq9ANCK4Rj72cTZGq0EjkAbzk9ULixAVMEDNs9YtLXYt53wnHpzJLyb
T3imLaBt1UE2LUseaTi4HC+U9vp4in3+qKXhVlF0r9/wzOf6w3cMiZ1Nfcxkc/Ye
QFeoiAmv49YGB0ceBLrojWoOGX5gExPpwdWMmkWHqOnheRFOCDtGyyL11MyevH36
Hd1v+R1pjWT1mqN6euv7PSYNjAVoK1LgWvPF14Q/f7KnNJ8mpdg9eO17JoQbNzcU
vQke3kqDFNDuMQGxbQWFRABAafW9LPdYeD4VHwk1YUV11uj4xSV8YpRsmUzP4l5J
p1wJjCQbaKBYmc2oFfp1aBQnwtiTW5fsSuuSUmgn6UMidtWbE9ALdUYChMK9u3jg
U1+KKwjPhkEU7aLqND91JULsS+9owwP0Kp01JobEOe3dWmsnPBpi0dgri64mCaJc
9LI+7C3Dr53VwHiKyv203p5YJwvGJo6dDYj5uXoaWiFE7qD/mK997IWoi6W+0+9M
pvCPjx93GyN1W5aNLM8xeGGSpP0BxBmxfLAhToPC+95oa/c2oYnCwVGE5dA2NgD4
91EyAkiNAbCS+RrLe6TCYjnQPDHBKYyxWFg1wV/T+Jr5d+HUuJX+6b0U/BrGHZrX
/VQq04o045eFLVMPXfpQK/nbHDjEmPmMhWlt7HMCtKq1yxp/4vbSO0/jD84HXD01
VSDPwcOMQrzIVxEB+sFfqSeqZo2cNmdVdGveNvBAXmKdCZt7RZZkrQmiDXGJEdcP
0OdywmSAFs0IWxPfgg11JGCDV+T3l22aXBawxAfcABNasycl/CUUmYLWFqJyqXdq
LD3Aieq6sFw9bCKJQVsT56XugPHETHUxF2siIv7AEFYOnyJbWcsWUjx5nsZfzvBf
rrQcZzWqiAX8hQPaftgshdk74VzEiMvBRPun0JMi4RPqawxuzwSp56L1buY549GS
veIxzS49P162RwZOYWeJ9KdovJOVnOj7pCfyQwdlJM5Gg0zJvF9hXCvZj/JjN/XJ
puBUY6VzNqVNMRcSnTRtXRS/NBBTU6gvut73xJK4Bkai1g4tiMKinwOUgTg3Nn1Z
4xi3aH0KK31Uw/3um3LTiPdmEh5KAluRtr+GFKeocgGJpcI8CDWHgAnEhE0/3d+L
ayqWBagszeAO4ONGB2aQ24j+sNJLCZlIy133YOlXUAATROy5oC4VAeffQYiRZt1F
YtJpS6ghgXl3OUBNAamCywvGaUCLqiUtrR92VInAMiFNx9c4JLlIy48jHa9Meha0
pLUN69+UmYXahnjcGlrKcEMZQTIprEu42QBjmT6Mn7VJWU/NKWctmB5C/J3uR4Mu
ACwwL8PwVi7iB6VgkEePWndCKmn8xoJlRKeNUz3ECk2JCcSC2+ML8N/wXxqTulO5
GZT3QiyZEGISkc4/El+P+Z+hJFvB+U3CiaJdKRD/aygM++kzI+vTshsHVjC55qWn
FdUpRXttcTcssINKYEUlfu6IAoVoKu+mCmdJDKMdIE3653QgXVf4RmbxEsRlcJbD
og4LvNgWuW0qqZqKvPFdfJ/O9h9e++TcDvBRPDBfjkCqFL8nGNbCK4omssBVIAVo
8kN7vIfQyz9HzJZBqO4MzK4SlqPAb2RjXjx/xUodMvNrut6vntqiu6/h5OpY4sMt
1/wDBlj69zyfLXAsL8kcaVgp81cdC73z0KAwo/hDtg/NdqtiUDiHUEfu3TaUZJxg
vKZlGLw0KEIo9mfx5L0RLQmFVzLNBUytyH5SKkTBYndvuLQq8BIlmQ694Qk2eXcr
qlhZOjM2g03B8kUulSZ2VVvD8chh4k+DtE3uOOyVhw1BokTKw2ZX0S8CN0upKaI/
C557dStndTbkOQtLdsMD239UC8CII7JHuLCkQAa2aHeNA2tF/FO+KP5sVdavBEy7
66sM06S8OSn4kVMO3nsNua+dRu36Zjsbb537CB5zWSb2WvmSnRbtCuqEX0Dix+fU
yZIwqhAyW6QIeoZ5D7m2xGaYEvC4y88O7AocclNAU3vYQuv+5UeWgwhYijvsLk+y
VWq6aomE1ghw0oSXVapiYZwD1fsM2oTbqlT47yhCaLyrSb+MbkJqTfVxoaH3/Uek
E6qmvNTuSQp5j0V6A/mE4IMlaBTjaV3tzwFjgtsGpzcr90pbYWhBTXQPBskbC2CA
37BUIWie8cRtv/bYotEXP0t7bz8DF4BBMt6uRrGSrBe9NcXwDimbMI8vMbrBDiqc
FTOXGRsGSO+3m6OUXbQqJAVZE9uTvodsumXe90CEqg2wZF/a5YCVLaa2PgR9/ORB
OBCtuzV6h7eYDn4PLpJxdQM3T2gCaUE1catc1jl79G7djABQMpX0h37AQvlDohIB
DHzmMYCt7bxYUjLBm0kgUp+qEL/sWjbO8yUDGWuzQfnvO0WsuQ91LDkLMIy4Qs+3
FCTnTiIbbGJw7w5ytyZzbTtq+JcamRtK3EVRHRbfSq1lOXnUyGhNcfL3DRckQwzT
me9MHFW6bgbqxF8nVUJmN4qBppUhCIVD+jnxxAuNU+svO5e91QOhX+NrehJ9s/Oe
8zN82Leffmu8EUc3RVr8z5dsYMVEyZ8TBTFZIJQ/lv+ZvtrEU8SNwX2/klGjNihF
vpD6l1QnFcGNrFWA3wqwTteI/fpsLOfA5EzL0e1R1F9GcYDLh4Bpt5d1AV1Zp5tA
qqfwvK8rqHGoddI4lN29WNaTXEDJnSbAtq1vnuz7P4qUVpzfO2IV2drt3krncfZs
3Gm/fI3MsIoz2y86SqwV0nLZgfzDcbiEMNk7GRHm0WiKjHPgW9y7+1w0R2OPTa19
rm973cajDyG959dwNYQ1AOT4V73xACoKqOjRUeN526BPdZdahn41bhTAiTVTFd1u
ubq8tUDXYGsgQ+p1OqBfdYxnxd67Oz6L4NNCIyhMLTgwDr42w0KvTyE4EvjVMIfX
7nwRvMO6p6/PcU2eTAAzkDI7xxpuywvFOWbEibL6HY79qvLURecoKhvKxbG/qN26
oWrKJDSwckb/c9L6cno/u9RNrJI1erJZ94uFy2UK+S+MJXpkjvVgnyzcZ89n1AEz
qjcBKLrxMf1O1L9yqvYo+hwK/F+BVfLBSIUaKcAe7EQXN9NdERy7i384NVSCL7zv
p5FLdk20Teudt2vpJkFlA+RaaeAt6oxDNheSOZBVpNMT3lA1BO/EYS5+qjWv79MV
HGgPz3FW6kVsCma9rTF3Odx/NP8L7RKZkdsmsHVpf0Vok3ARDvhCVRJTREE70kwB
T0VH0tDl8X+ExmHAprGNCjXgrvGuMocwJlYZIuQ6AcSD36VD/K2VFR5yKrAzyfqa
WPrA7f/xWnLBddYchf5snsShiwEp7CNd5P9HJFhvp+lyxxgj8U/7QGQm3op051Kf
JJILmZWYaK9U9qcv1X72/nqTQrMDVg9+QxN7hMtjZP9WVcq8l7qhhGFwO3ThumEq
ZIEjrvIT7GIhB79BZ4hiBGdwBmSPkLWtriIcwkcHs+Uab4YDnGOxZPQ4ZefzPB7M
pAbzRd4BsjmxNNom5drAjZIqTECdvUgoJkrXj1CDFUhEIwIRtefkdAl+bokikBBD
SbBdsRnPl/I1YJJD5Uz3R2XoEuxUuKROoqy0iClZU6Dbaj+cDF1dNyoS2H/zhyTa
BEe3y5y8NxAwDWg3Wz8xpMkuzmyeDe9VfAy6HwjhTITRyQ2Wr3QmqShiUCVzMiaM
HuVsKtKVJf6VxUP7c1HfLp6dYLQXE8pNXyftbOSNQHpiHPmOc9iotNc3XsTIT2E8
8Yv1K711LYXbcUmFNdYOKYO1Ad2MVqg1HDO9FNBIH2Iqhxo/82N51AqXKIOE2WOR
0QDPDNODaKZhsCeseyf/3bx7BC9bzASKcbnahfZzEILmVH3OkQokrYXY63sd7S7S
Yj/ovWCLuwfgpIhUjCyiZY9mSUygka4kfR5MJg8Tu2nEiJzokprXHwCk5x31aOZv
09mqtWCyLPy21wr/yh28b4UC0riyMWBz9ZZMbOGwXYCi0yjSpTIQcR5VaYvR1YtJ
Co2ShCP4GKm/fJ0p/rdBzNEuoEl+nOwHMQB5d5rJ8CwK5LuS+b8jxOn2meeFYLXz
g1f+x11JIzOuqA1zdVwVSVNWHdEfZ5G2lJB7D8YiVWo6HElDs5lYWslaRYj1Vynz
VoYOgWZvNBRPZRbdwlOgHB10e5dBIbQCnadB+27CH9uL7cHujFL0oMX/yztJEJ/E
4Ed8cSEMm6/zfo444pHjt/ak4EkrldsGirL/wVDjvhScwC9ig+KXdA41g7R7QAvo
01IA9rMXvXkd+KElfpZPW9xsNYlZ0Ie0osJnhIUVeCobqA24lXUqa7vjOHhADIeD
XADdoQAo5A7bwXbQs54u4d+YHJ5QCtb12QQX2bq/svVqKlcgiVptWA2UrJ2o7aaA
VaLQ0wUTw7+W5nQtqFWAgYDaX+LeKK0U205wON/AwWm6clnH7R4cLXZbkETskSFx
kK2NmQeh5IQJfR/mnYjG49c7n0ghHIDLnJgInBzgsTOBSCYn02GRbDVCsoc8rUq0
D37c9maOnWWo2fBkc3X1NsDmkkmUEj5v1Fq7rRXwrZi6LjEpAlaNKXwCsuE2eGb+
6ZjnFQegX7Xag/FkTk1YH/3jMO2+wzV24cgvC/aALFtkPR+UOgANl5VruQvAFHjl
ls6ouICmDnKBz9pcqth7lbP12XViqhJXaIEJlA9qHpsyqIrDavfNnFTfqBFniTAW
G6aIBJ6MG2VB+z9m7AtheoOyrBic5mgJ9GtUTgU3dUAOEvwrnZZjY+uTtB8pRxfZ
H6jWWdOaPDy+OEQP/eUFhXCWkB5aW5zBBz02GFnK1Q08OhzndG2SUEndPDZmd1Iq
/u6SWqplhellnK8vFxezpI8Z1L3mV2E9bVa+AMl5JLr7FEkrrJbbiZuBbS81AEdY
kv4ENyS+LZqUXvoOizPo3ACc7BNCoJpWFqVpID6OorEekP7sK9KK2TqJ20ySi594
M0ddw+CNNG1oaarmB888dM4BNf1n7Bmkxd0rQMpgiJjWJXsNBHJo4E0fQJV9R569
4p5ssYL4UHmpRUr0iS3GBV5goWXEnlZNRCiG+C8yl2uXNgFJgl961Ogu+3hm7FTu
8VfcsUGIPnHgVp8kq6gp2lN9zVa3awYMn4m7vHSkSbJcfYXF4JjkPdN7V3nNY3uj
3B9Wnp5wQlnJXNm6qJ4L+ylke3Q7PH05FcEM6IjWMKevWNRaIGOtLTvhOOeCMTTM
0j8ACUKLxZwHMBOEOiFRYAYBcaRdejkDj9sC6bai3ir7MbumOMiqn94d77/8QtV+
NocrcrOysrohsi4Lgb4IDngMcwRO0Km5OhqTftBLQCAopUEYuthmR61G15M+avFa
2dPnwlDtxcyEToraZMHocJh88slil6wAMZWwe2gE13iQfIQr7OPS+zLwtGQdZggF
Zk+ecF9XVzsVe/k8wH0OH7cQ/K0AfFTJ7Iz7fzmWUbiqlpYbCew37iMtuKTb/MbQ
h2Z8L3D2+n2IcOcx1MXYvNjgEUY3V1giF4yKiEBt/QokZ6+gz3HlLd1EACB0ih1K
+hPqGIzAZqTt8eUdT0U0MsLHIy4+dmAPNml6hWsIqvOpeYilcidQUIJ8lVX3sEmj
X6/mLjFFWh5LKiIESMS0IAXNRqLMQzgo2IGpTqEls2YaQXTPtakUPxHXdyyKReJM
ldCX28F+v2a1y2u/WRCH5onVhlQWSCd/SJyDb6v3ViK9Cax9SAJvJiJ76pO1epvT
Y7PIy/uLAah9onaINLGXkjYAAHCxbQFGMx81Om+rc9zVIU0kdRPvzxaXGtvDHIJq
x0QvNenhOHKePBJDzOvCe/zOITNA6+XJSiB0cFJOW0H2KJA5jH46T87+8c/3lfKt
mOj7Biv8TW1rLbskpxyz9mldhayqIELf/QqNOXrzqBnkFGbIdrg3BmGHlU7VcpsM
W7bZWp+UIJPCCAvGkP6m3cIvuRy14A6eZk5CnmGq4nbTu+8USBfs0o+yG3tKDbGh
iDWZ5ba/Gt7DYhGSUgMGcR95U39H3bFsOJvDwmcV8gWEnlo1aRl3RwaF3uF5agy/
RT008bw9SjlXIQh7kd4CJWLxR5hu43zKkF0MLtwyvFmMvcYg8gRt1hasAAZMU6p4
TSo0ARWeXbqX5IPEQOrgkZkEwXDvbXDVviJJlmmbEkUmLR6MP21aEqeR3XQLwbE9
AQ4zxXgtjL0gOY1v2V0x9NAdVHtgxrRUhHfgUa4oBQoHaQFuQKB6dQobPf/PZnfB
UHm9J+KzI6MYpMYtDj0e1vqkxCuUNQYHSRfpGUDddZzU6b0sud4U7LuBW/oOImmL
YNjq80N4wOTI4iN2GK+1FC7hHwTkism72QhNEC7zNhHMeOlnk+X8Cvs78KxudhhV
9qKqlL5cE+yPKYepobqZH9UcuUjAQO9gJVd4MuHB3w82lMewWR6VQD66s4kJN5XX
cYl9P+GjiUInt+Mbto9yjyeN6OLCw7jf7CxRNAFbTAS/3F6RT7jx7VXtz2LhhW4N
M78LBGYee1BS5nMjHcQvhdk5obv4zE8UX0T7PmIozt+zhwZ2nu469uNSbBgGdVfw
Iigc25fDKLugJBbjhIgdTSb7DaVvok6r5tT4HIlbJDDJvOspU2HutKXnerhvXpQY
V0qUlMng7slol5r56wkw8fash4h8EHpviTScsYzHrRGYrt6IBNIZ37wfn1/AmyGy
rYY8NJ5uak8v1OwsvZ6aByVD/DfwhZVhdvbSzdXjCtBawT4QNDfUX0nj8nfoyr9L
T8WO6MBkIcsyJLYhLggdnEp5ZRkXALWWqq70veDjr4SP1uTHSuPhNDy2mGtYwpl1
l76YU1BkPWk+ZW9YnkO7EPjyKWlzV0TnVZsqxk7MnCnQfAs2/XqfuXMTw4GvH3Gu
1HyivKOSV6KZjJNqviBg/4dQOmf8gzugFcsIjrRxkUbzetz4AfswwIMnRDbRSz/D
t6VP2ArwFsG7OIzStTGb9FJBGIPfmiRIe0C0erLXUf8DJfV/B/6jVkhWCi/5ghsD
0gXb5svwnVbE7i1Nji9VwAQdCf9bN1vqi2RKCNOBfA520PzAhu3HmA6g27NhLhdT
zQLeaVdCYkSdj1mY1EUG0udiw/Pd3JdkzGS6oEHrdYk6Q1x4apiStKxzjv28b4Pe
ItiNRubuD2PKD5oYoDUATw8CdIAH6os38SR73cDw1Xt3znumieZYJIVI5BX/CTUO
3RM1UhTu3XRhwaq+EB7TgRAFRR8YuXfu9EWfZrZ0qC+hWkyNF6873IJRphWcLIJz
hsm7GyWtDJ/MawhmuVPVBgqjWzTv8cthirp0a2/gRTFnRpc6QDg/jyUVrIAYt7bM
BpvE2zBab3FVkXL/uTRkQdhwRaQfA3eEMAnIPU8J0QFwmSva/7PYbygk2W1osGMQ
HVGHuqzhoenZe95yoH40NwXlUvZmMaDZ2cNLx9BuYCNugej7kKKDRNjcFn4X9434
GjcXN1nYxaMVVJGgFgwWoI7Iv195gfvizM18KZv6qJ/j0tWzVPET7fcJaVFUaqSq
+IIdPY4qXTYwF+NmrWpm8mEgwtg+y/gtIuQC8MmMNPTn+W/OzPD7C/p8DjcGihV9
hD73At4se4PYDCGvoFh8o8CetVC/mB6r3Q5vI8o4Cmyj65FvzzIP8KRnGq2eIEzR
+Fzv+XvYcdpVGP16x44up7Dgu353IBULMy8kj13ca3VMA7TCjDICImu8Q1LFgn/b
SMMPRcDm3YAulnlRqlaP+SQDvnitM+AmH6Lbyqyswcc2TFJihk0Bm9XAXEFaeQOZ
sXKeuPNorjGjycHVzVn5KheJtveC214ZGuSoODtgHDhQIlWyDD12NrPwgB7pHDR1
4BR+JCUPB6GeIQHSV/gyuIoGOPT2WKRbMQR0xqQL3Xrw6gL8gfZ9nungGbYAyPjp
nC/QitPavtIA6QCtOIdKYY+8e8UIA/0yfyNxxsZxIdzDeNhHmYN76O1u00eDQlWS
4e4feXb8mdV0foNaHWAR7dLdwyU3/KgoK8qNYYht/55NspRE9eLziRYJm3qftllZ
pWeXBgjxEQdhan6yf/scYY3o2xtzK6K1MWoSPSFYY2saJr+2a9ImZjHwqi2NR8ue
LbSqQe9izLlYYAdQJDp6+zZ7HPRzJmUnyeXjQ5qE6jPulkj7/isc40rwKYnI3RLr
tjd1EKcRJVn7xEX3jRwgQot3U2Jbspm9+urRsOxPiBGddaS1Oq65z7VG4BNyDMZu
kQH2dXedVv47W9lNLAddL553zhiwPBI3cUQN5Met1AweA0tAoZTv9VHbrzJXtvGx
Blv0ta6mfTrf1FwHPOErpdDM5uS/g9YrDXXthhKsR+bknKf6vpxPEkpV4kIY9jb6
28sK1Rd0U+AVdfERRnd25gegp4j+KzyJLqiq056WxScW3MBOoOWeaPH2imzXS+rT
znuXpL0T/FgbkAejlYYMUlRuLV6AksVMLTLnq2skU4GfVghsaGH6Hv6LwdsZKaG0
M6nHj9aNjNURvGzpB29Ub83KxQekIMUx2s10iEX7pRKazrEUWgKpzPiGDyyivOOP
FTBUro7+s4JvrpzVZYzRKgEYCIsmSj8HPRLRPfYnXOD+k8E7TOg/SMWZ7NrTqKxR
I9c+z5IPOyevNBBJ+v12BPXgUXE1Wne8XsvpKAfZgV3WxdRtj4oP+/cZBY6oEal8
hLNxv7ni8fbHlxoEmv8ef1Bck3YG8sRAK0bfH+hxH6+SaRFc1/jst2pQJn7zHIJg
ePSjt5yAYrum6hnQoX4nPSVmhpS5ebm/jiN9BdUVcKocEBX3b2+TINMpAEu4ioqh
jvT0gaYNpKnDGyPdj+D9qhhrn20vZx6ji4o627fx37elfEyXvfzJN3PdO9J5cRtX
Ao4I60KnRU2Xs01x8pU5tjjg2VQNg5hUWB+Uek0wE7TgJVOXBJqCyqXyuKKHYtfR
alvwjKoGQjf69N9C7mMuXAwtNmsOQ+92IzsyTHHc3+4HFCTPMQ99t8rIaWYp4UBk
xtcmTu/3ir83WUX1z5qa8Ie+kjKJoi8vUm0ALtwBa8AVEw57iud2S+bi9lTkxXJV
KFbu6ELNlNuP1f1I6XFoEnoosr1+AippCaT37KToAKStPQ3P9hNudnMgqoBqmZh2
YyW6P3+fzaUJKGeFuszEKZUnPoX44nov/HWOXkWdTvC83wQPBE6dyBHg7cme0bNC
6hIRt9X1jzZPm8rmUVzu/+7Ho+qbUTIY0yMey6H95DKwFXRT1EdvmsUaL9Hb9qBX
plj8E2UwJvd6fLy1+gi+FP7PKvXn8pqb94ccLlK5RBeiOqIsA0pzr1E+N7THrZxq
mndhmKSL5/ov1fIPv4g2v0bqHaGvNOsHZfFfqMU7CdXK4t4WxzqO5lDTa1WpXpWX
ZsS1Y/rZyg6grrra43Y9LCICsK1+Y5+17beU7HLRfXLQe0ds8+qnVh0miwfDaJ2D
1uGDTHKxAH7efDxVRAUafdmVLxGM33zpmJ4rU0ZFAa1UhZjfZWytLrRZ9mPnOwC+
7Sq/yzFCxyRc6lcQvtAXf0bHmc9jrAp9b4BNi0t9RIdnpIKbdiYL9GOpqgiR+IYA
mggkzLIKoudyninbDbGDfBjiABaslo2YkG3ES6O9wNO7pj/3UaFM8MgcrXsAbhqB
Kicv/f1ygSx7EZXTa5IC3i7VCvA/OhJ+OOcJdg2IQekKewrpD3tu2/TGaasDOX4K
hr8iyDwsqst8PWj6mueFVdN1c55flaZw9NmQGnSjOKBzrp1OmySlwdFBeOZnYMAE
zDk33Jq/theFJit0MIua3aJWAPhm6SMPBgWairfWVz3WO+nlKeiwmPfRZNCfYFdd
HMvSbl00OYYS1+9sN0v7r/tW4pKs8hrQ3FrVfv+KUrx3zpO0feANyBzUgJPmkN+f
oQYFE9YCHUv87u/VYF4A2PgZKyREHeN/emDvC+Ios4+BqiqazhS9/7B30QnajuOA
fVi1v7ivwcrGTW+24PigG8Yk41ASdkCiJRFf2vOff2whq5+7E/QF1MFhecTaX6Y7
5hBXYT7C9jIhnHNRdizPOc7nbdBQmO2v+Sra1qmJYdAui1Lf5JNMGC/HKJ1GY7Yg
uzvs80rplfnKOaCpPTe1NIM63zi47sR4rl+fERa/xvU7oZugi04lD1YgjWdVCWhd
lAMKfs4hs/eFLZkwSPoesV0X2iqSo72s4eKNIR8NBuE/Iaer+ZJyAP4Qf/pXA/JW
EsXZbOptZYDwDQgz6grYPy+kLazSr/NnPOv+0zyl6TB6LOQQXlsDlctwa6mJuHpj
eegdOqDijEuaODwhaZLzytLpfQ9h8Ft4RLl+qm5i5zjahGQbGp0eE0JnJM4r5+YJ
CJLojnz8j2qR41qNQ5DH51TGEGXJ//1CMQinvXjJgIhlyZ+3pUAD0hxcj4QxHC7L
OWFp04YtaM8/Nm5Koj9CmY/RfPpR9U//8VAha5q0hRtEJ3fVKnx151nenQyLYMh7
bJAwIGegZEdgtEXDHy+n8dvlgT9Y+n6K4m9mQoEWEzFesmoq6e+IJ2k0fG2FTioE
C/b9NEy+ofm81lwOEaWRGsmjbvFXzqr2XjOPvC43L/0Z9v+g2ZWgyuNSLk17jdpT
FYeJgOPvNhMgt9wf5VIKWvcJ7RR9AVw63awv9RXN9krotqEIjMQAPKwN9Y3wNiAp
eL7qp+y5NTyMkkfBTifLWbJlFBhKC03ZoXP0b8p44e/K+H7/0m9MNwutwFzvXwvN
fk/v2jWdH6rDUszzdgDP7ijXH/nPQPKAAUtIwvw5FRny5n8Q3av+JhiBy815XmeI
OW0+KDVyrNyCGCQ3bfbxJ/MTd54cTN/7VxxKygZEsIKa/mAqUkifsaeCFrKvNW8I
pc8ifWokY6ALRPLpiBzWNo0ziH0cOSmOiDBefv2aZ3hcxGf4/UuSckyqLETJzRJ/
YtPpd4j6GCRBR2SifFa+oyXc8wU6BnmxLXqhKs3xH1HqOTVV9TQwnztfuaz/+plI
L8Z5SsforR8SRvotvw6jF/NB8FoWgEFiz297wIKzzJKQOeUCvo6UvOOnBJGBv81X
tBfn9hs1fWfH7r1fj/oQn6G0j92YLDInEa27GzDFU7m8uYk847TtVjB30L3o3VBk
83AIsxeSTona0MHarKiuAWelVjBfjFswbvXJhgilWAnDVGJl5f5ZQRIxOaCEcoqg
vI79c7ifa6xW6l+VfHnG84QQXSrGRZotfyM6XS2GXD4o1pygt7vZVsBE70BgbOam
rCD/TfFnTZVp0Uar/vlJHFgXZ8dFJEz4dRXBXeYeCdQGY3AiLwF33I9oxhOaCjLQ
OEri/xCdiZ8Rku2gh6A68aTe8PNTCFiO+3AlnB2v+0tAgudj2VNYnFlca1JfJaXU
W4RB/lHrj/FPjhGkAHWADEy3AKUhZ47Px2f9Bxbv3+SUKOtt6z1o2F6NTkfHGAqD
lBacBmu50TKuWdn6i72Ixd6eIV2iVJNE38cavD3Nr9F1M9DN5q+e6hKFHTqNDT6Z
bXEhYVe5CEmL1/d5OnFOsj+cuO2gt6KsIEctLeXibAaKQCoaszKn4PVScFzySnNn
sXjb7BmdoMgoFU/ghxNpnEWlE/ki2SLQ+1MW2s1Lvp0Fq/sQ9vunOcU//UKQDR+/
7YscNRdbmC2Y9BKThQX+9vBFToQc7KjEmh5Ntddm5Py7Lbt0Wv6LW7uJ87VO7Sbb
XF3shjNigfRv5pd2FUS9pjVJ+5/Jkoo7ATe1m7MU3Zd6eyZsrPqTqEf4PDCMJ5yD
pR45DOC5/kHyDmJCv9RFif1V4aYOm3e5t5uwVU0sie89LnXtdcSVeRpWceKk5f+S
bNd+oXsrU9Iu0Rl3Ae8B+rzBCxDYn3otxTpPCCkm2XZVwK15zoUXIb0YP3Zv43nt
Y4dRASwxOyPRRhY9iiirN7NsBRQNBhbubSyQ+zi+Tyaqk2ORrU5OrgvV0NA+0YpW
kXDATYNOUZVxClQGDaZ26SNkhl882zLDMtKOSW3hRmLIgKZ9SrxaFnlaBWNSYedL
2sciTU0oaVeguA0xMdC0ToR85U2JHQNKIyHIaSc8GIP4x4gv1TqppTtMTR0IyKMW
Tw7jzoThzvMC6Bu1l6Ke9t1TdnVx61b8FHNl3YdC25ZEz8Vhm1gnxz4+knbu6cjn
MUntT2E2TXOCivxGX0W8HiZ0vBRL7aVMuq4e4upDp91JoPBAxHDkQqvTbYv3D3V1
1msLZydJPktc1ygMfd9JFLkT3v1A9yzFGc4k8C1ZdWvFQLb/6ixjCTgjAysuaG/J
63wSzenDYi7MQ8ko2CnpcHrY257aVoeRYlF3SgdGrg9fcYXSvPkgeP011Xd0nqlO
F1JN5kbNuYhYPux8etiAGQGigfRpzY+OtVw98fypa4nMxd+l377Q/HxsTgr2IMcG
pFgEaZuIFLVQD9ElnW+mMQ6ZIcAGvjf9EZBAEsLG6VFDdLRoUfp6Cm9z41W6dpl6
kmm+83ei6uj2YsLL6l7qBRWsNRkiGZhf7K9/i9uh8RuTl5t0XEfEcp5mioglaLU3
NfuCE7IARaSqU8tCBte9jZIL8/sg+g7LwwBeOWK6VhrZ7tuGVTWqY8ICQDqvRrQE
WiK5ESQIpo7p7Buuz6dHYPZqew5JuIL6W/x5GzAJdqRWYgOdOWQOT1T6K6GiSO5M
kE8c1kskrHyyh1ln+0aLP1zqs3jmwXZiVu14xOKnDKirgLxy/yzBkjFdhyHgmkSZ
MEr+MS4Fv5ispFRjSCGYQ8upM5P/7Tedog4LnLK6vNBOusKPKLEoKfbnj1Xpy7Ie
APSqQ1zIoBC1oyHkW/u+2cfW0LtyIMjZVlNTSbu8UaBfujsYu23/tGGPBQqEs75h
aqnBGIA3VSmwhiu24Qce/fXa3Io2NaVeiFAA77PsL+bJ9WY1WXQLtTl+bACgUBm+
P5sj4eAr01DsJ7GkicN9yT8b7zfYr95tYwWHvGtNJWASv11GP9lGPJUr/NyV9771
0T/H4e8WigrfvoZAKQCONGX3kP6+EbUzP27FJrJ8ECoUtwlcksf7qc3Bua7aWKDb
EGIdzC5r1AE65T4VPQ7DzZvF1nvJhYNLz7FYke3iM/gIn9ghO9bm+ms3aki5NlrN
btqXnacuQ+LDJJ6Q7fb2e5q+e32QuBHSUn2+g4XprGPhjx0SV1lh+ITia3SDTlk6
mRc/oy+27n3xIAo2gk0eOLxcbs6fmsgAa+87WFKJbdaxKQDLL1R52B4IfhztkhIw
9ubm/tD392aP5oiCO5Yg9nlb8NE5nQPvZF0Z+jOk4VxpL5Lr8e4/luCbOODRv5bI
jXnl1h2LNppAR96lH4Y8CRlMYMjArw5Ct2w8/Is6L1oH0ZDDrx/hFv8kf9Gf9BtQ
QjrvxQZ6cWraZGc4k6SteMZNIsrSv7OnH4RYFLNuadsSTYWcgUNNxgEUunTEp76J
Lsl2b3h4nJDCmbFZdPdTUC57LzDzwrOizyHUxiK7PEqt9EviO4z5DE7jv4X5tQ3y
ZK2fm4flemG8HNdoHBX3qKS85bm42dyqDIwBDNxMzvf/MO/uNVbnEueBDkF4rc5e
vyX94xcUzbbbjMy1R4JK7tjD3M+uEYIqBpsD3TLaG2pRKcCGzl1ezJoYv/9jgig2
UAQoZvvo66tpgx86IBBh+eHQ7fdlpCneBWz3maX3BFbIUp+Ibqlfs9A6z2YUNLYY
+mmJuC86oCnK23MI3o3vBNUuliDbZX4dtiuYqnGUQmlOKRzjL43KYL0ykLvixoC4
sGrZOzBGNgIbBRDlDuUTsSE1mT99Mf9LWvPXQWu+TjDB93EV7v7uQsMF8LsXDGHJ
bXRxUKGT8Uhx8/yDiQ2FBKc4IF96rKFqWByyoRoNZURjzF7XHuwI4YUUnEEn/FVi
b9hYmTpO0sRwMwVPddyNU+KBENem/8JYXhqy8e/rnakbEbStR//ZAN4Q4LfGr5gL
q6Bc+YZazzJCovgP97Mshnz6mHDaLxv3LYAXnx98flOKHyeRTP9zcVOF+Teolpaw
79RyB15bcfAGTnvcf57Ys/YX6P5DjOKf1Nm81EKpHYgQo/PdDmS7eFA4TRNGJWAU
bI/yjbz8Xz293d/SXrxjyAYVu5QMPA/8vFUXDwXezS91FZppyLC5AX24aj64iu/w
qxF7N7W6XrRFjdCA64JNcJXACZDCVqn3YiHSpNjNAdu8r1zO5CR19aeswcwmKvYu
cUiAms0qDbWZOgICMoLZY5PPXznXjY8ebq/777cYRbXzZlikx9nOWVpEt1Ed4czb
VgMAW6ingFOXoOo9S5p8kX6hJegx08T2fgqVEhY5tMg8j+5UugFbdSMhuEUVomqQ
7D0yTiStCkNl1UheRWRqZ6Mo/coL89IAoL044Y2o7YzaHPhLhGo4RM7wkgDSc/to
A5L8dgluZapxDWJJHEK7A1yfQXm5GB1JYPuc/0TrkrOyI+1iSmMDAb0USjV6HuLZ
J2k40hMQCXoijOUH6fyc5/oC+FLZKkvIBQQvVtmG6kzo5fTfk6qjkXoZzxsGTboi
zAW8ojUuxKCOii9NnH2uFa/4KB+6tOQhMv7KXlpv3fvvAdBjqlAk/CcP+J4HLuWX
Mop1kuk+hdJm1tSpUTitmRM762HZRH8eJIMj0oWRJt/OsvHEqqlcbbeehtoxJ6JX
kEtqm5ZohJkaffZIN7HvkkXXK9RNB9j6doFjld+3UqKBC6xsxc/QJHArEilSamQ5
OHnp6YR9jGRlEvLB20LtyUVuc5yxgkGJ0s4P5C+ZDZBeb6G4syKDjpGcSq9PzYW/
cy8D5zV/HdD810Hzp2vpV8XXYqFcsm08bCXyc2rsCh6Cfcw54iYaVx0F4JNrR+as
5CyN51JTIkqOZWi8UBDXhkdZNY5QV28g5U3YwkWClbfo7JT7DFtcnolNGw1hw8Uf
Y8GsBAbW4V8ua8PfSU4y6BlxM37gBEWxWZxtGP5+yGwYgHayViJ91GiOCiyD0Vig
SKo99/5hc27260UoAmvrZCIOKOSNzHcP0Zk3LQe92fwpFiLbOObLVHiSY2Dm5n90
8EHCB02BLPfoM1BqduRaot+3PO4+0vGFLMO7rB5t7+WlHxA/sb36I7N0Xs+EVOur
96u5L1SmmgwvwLf8prq63x7ZAzdrl/CrR5Oth0eQuH7+LiNjs0L+xhzsJDH6ZKxt
S01dNupHFHWHg1ZA6uHpt/jbSZIpMOoIFEs1MhBAuV+j+DeYFSGQEjjJKNQusoqa
fiyehX0Jsqmx6VlrkRhifsQoOhiv8DMiOz4FutqBqYTF+XokhQ1Q80vUjAF056GI
TQCeNrG3Bv+KSS8cUHbFgpZpOd79s9KoaSymciiPAdarTDKa23uMJAARibN8zKY5
ur3TwTySgSH5K/7v2vpoNb3niLJN1eSKQjsjhFEQ3C/cezzfXWHPVaqn09KRHR05
9ofMcfvk4sZkaLw1PBYk0O6RXPttAmKKhfHBYeMsSP/VyzCgBvcSQ2HELurT/CIi
xpO6vzuPKET/3tXg8W0yk//TkSR3xHoqpwqP0q7dJPHYtw790xYBqRr7qYFryjsO
9xEXuVR6KvApy4mg67p90CDBQoK2EqKBeCl90b5jR4nsfZ1Zt47Jn5Z38uCIVeAK
9qa8ZVNQMT/vu68hGqU4VVA4J5mbdornMJTCvXQI0bvTApCIGHy/nnvOpCbtCBeD
1gnAeQWpz2i0+s40hgsXj3JIc+d8ac+GLFODfwXFlmh0ji9Zw3dtj6AaLHwL485Y
6jDdMf2h1IYuyXP4mDPj9t5k90FrodsjfvyfNi2l6zpYU56ErdQ18QvRLqoDmVLx
D5nvnimjY9gAfscFW88LtYeB51UdF5kk3Rp/KjEOQWJU3Z4TbLOXwS9L8Dwf87OS
U23ZOniW2+Non7uJSnKTTIcJxq4qexoJZU1jJeF45oeOeIxS4sTaMgKURAAnV3F0
I3H0ETDTxRdNi4UL/ol5kC7XshQDqh7XRIkCC7M733B6MRl/mtd27aKiZYS7CQZg
/QjznMuRwi9hGc5Ue0digRthReJUuq1JNHut/75WIonFlJLdkIMNqHC3Sp8vHG7q
Ns3ZGZwA4/8ghWUUTCZ7FITGxEV83VJxE8t5kfDRAvg6ZDGA+kI43QfWWFT1vK2x
6RlwK7fmwaf0NB/2D8StSJR+rssjr01jNX66LVQwHflJYFUE4ok2P4az00W9yCYf
/doRfTsnnjhUPpVDHMsxOfJ5qgT7ywefspal9OjMBfW104zEUrC/z429Vg3acc6M
U5SNfTV/q4GZkgkecKk43ExHm2XhFw1JDOkkFVpAZ7yGNzSnsnmrrcdEa4zvoG7P
y4VPdmVzu73nkPHboumVTZLISSbYnbxvN9IeE8NhBm7lN5sfnqvbU+5sUfJvl99/
8BX1E/NNZ0iYnBMgxIg/ot5ugQJLkhh3EHOpx6URReK4L3R6Kh724xbZp92B4g4J
eKAjWlUwQNFDm1DNn0sJUFTboX/XYsXmxhJta6ol+c4Sngj2PUtL02KwqLUclMQQ
fM55NBvqeb84A+9woxfKPYQHXu+lEv2AmKfW2ocsLkRtSnvUx1AY2UJ8GY6fH1C8
V5C2gz9fJBPQDuS4RuUknmRS02aGOJ1UufEcX+MFSbq8Ok5FtvEmExCeR+7xKkz1
3RxQB8bYwfaNKTYFpqqBS9e1udOBHCGVbgB3eTIvhi6XofubpWTYcvI7OUh8cIKW
mMN6NfQbF/BPQtpTZQw4jNuTzMJBcsS9/twM5lkMVauUQnB0uH19IYqQB8lYZBMa
mNAO7XbltFZaTbfJq8iwCcSHGYi0Fq6YWccve96L9aB4g+c0mTZZvBrhiGQr77y+
TUviSkdDPzLChCsLeJBuxvk+MCsLeGVohIYZ6oaUQGNJzfjx97A0/yI/m8pqGNSs
a0Ahm0hMJHPqqbUCOKU/A5xTxH0nbxJx5/3P3hXnaGc5QbWn0wrC54ETCs8Ymnhq
dCeerrc05SiM41UPk9sqmGWi8OmFKfcSng9DIdcCbPhSQKYvqPpXRF6KjVgPvWta
KXqdzMx8LyxrA/xcjn5kIODoOJlWr0QT5sgh+y5RPXQA9ILtQCZY4LPh4J5uyqzs
s1k1niPjoL1KxHQn19cfsEEjbIGsgHZOg1kuhLyV/7Fs71DHql8t9HU8TMY8bruP
ffKQGtbvvdHP5l8W2QWew74it5pBoS4cx8UGkcv5OgWJtbsUqmx0ls7j5YE8oQrw
iwEz+sLv/QngbVGIcEbasHw/az3p5ycsxQjIVmY+ItF1R1A/8PkbggloEi4Oq2C+
UKuDfNupypBI7N62PFGWQHthDlbisV7Lz0eBxC9R3zJWxxHE/mciyB4yWWi5lu+Z
zerYSNLqnGl7/88Dx2i7PcBI1hFezANAlICXd1ncoogWKvxm+2q0EKsdERIj6R3J
DZKm+R1jTXgZfBrABsPB2oorOWCwdWthioSae/EZKGgnV4fEpkgvQqGKr4cExqhB
GucoccvIFoqdVRNnvLwHl7MQVov5l/ERVXNkJe2YxyaT72TRF7EcLxXru2EXigOf
jQJJheVjfaMc8L1Xuy3wdMlnZgo7cINsxIhFxRtLduGL4Jq2Vjkzq/j+0NUnICNq
DAWia2Ms5TtGTcZH+3QrXM+zYkY/r/Nv5JLfuPcIW+MpQb7395Qk8txXUITTSY9I
W0nX4OwAZpLuP5V4JxZrAInCKz4BgJjnnpErH5Ykin5Y3i3jm5SFZmyHAU2RqnOs
eWb8u2CFHHsO42OIBLBeATbP+UCFHGJY60U56hrFse7Sqd5wjh2y/F/SS58t9ZB4
TjS6pqZpWvEO3Bxu5EGscSqTyflkiHmpJD0uxKDEfnBn+Vb1vOYqY01Ie4/vx+lL
9a+olQZXoATL6ppHHzXQWGqWRlimNw58+rFJ7gGKwzcz5uoM8lLRmwiiMvk5Zkn3
2Z7LxfiJZ7nELXBXksGxP8hRJBBHzqgqzcklHCDQuPwG70DGFne5upxo3OXoEVXz
lOes12EngsUlVxoG8QIAP0RY2S1MPeYWUrdkWfHJkc1kLnnlf+L+L2jqKNVHZNvb
b+YxGFzSL6N7ga1AA99G1RfxSxRlto2TXlsYaVyYr/lWplEcF/D0F2CjxezJP+pO
xeXnO0FU3WiOP4FENkl3IDx8IJUZ2a2i1s+jJBXYrQI8RuW4g6HqLJxeTRhgsPtf
fld5627iZHrua8Pe2mlKoiG65d4QIgCRV0CG3zYoDvOtxfRzeWeDIzNukQ8j3vTa
YmHbYMG8qrCcj3KlUFmHSQwpQS4XRyNL3XxHQ0aRdedllHxKdFPNouNfUVaq3SsY
UgxoeExbpjKzaKqiFcFrpl1nnVuOBa9jEMJ0J7lAUdbFxDPk4TjGEFhU0vvPBKCM
vpN3QzFP1FOpFgTJ15iiz1AbqRVZ4vuTpI1MpigKDaSN2214eZ2NICziYC09duwc
XgghJXGYpQgMUDkHy30Hv7R7cG3zUTsEuqWob8aOrTf7rZH2Rtd6nxeCJWhM+OfM
Dxqq6j5J3lJDG99mWzlNE7sg2WK88HfYNDxWgcGRQWdHJqfchji2rbG6KLgtughC
z73/8Qy4hWmaaf7QfEjYGyop7y0BU9F1AgMfVZ5DFYMj1qp1uSen/ZpnTw91WmWI
daa7bkMdgOjFbB55gY/MZyqS62NGg8AARQAjC8GnUH8YDCpTHfyg/49CyvCZvpJs
2J52N5ieQkKd6EKhLckV5XekAsbMmmJlKQQdXP3+t4wQXdQEdrlb4mLLts5gBRyG
CfB8yj3IU2dQigHavOBrcEVprKc08pkfUpc2HAZt6w3Xgq7Du5Bbe5veZ2OzeroL
L7rC/41brsxU/HhiBN8WwfBLxQoiOETHSyaPYg4CKlkIEb2JVKp4/7NrsrYCFcb2
9QYGKm5rlcSdLA3iXmuOeuPu/+bCm8Zcoy/mD7zDuUXr3iQNXAdlk27S9LbUez9d
M3BTqhIT+sEL8qsrYhp4r+GlVMnzkLVnG+YI+kHASYrZlhsdxBnYQodfCLMXRibn
RyaofQ4ipvuTs5n0iUJj63qtanrHaBggMnHU9IuMcQ7+KlZwNo9r25xFqcMgEDoc
g/FjVWSORgP6ClnUJyKxH8WV0zOFpSqXid+c5yS2zY5VHzZ7HnSy6BGHS7cKMV32
phNzc4bTBFGV2HnzHWiKwnqSW5mwDqcPj+dMOew+Te6LdHBhRrNZq+HuD0/nMAdR
837GKlVvH4vvjIgO0L4hxlajc0hi9pGvds78VpmvuCo4x6xTvg+4HcxJB+OON+mp
GPzMfD50rsQH7sT/87BfLmtkah55GXB2LULOoFeXFNCMRHQ2TRW823m9MlDe9JI6
KKJ4ep6vDwkeLXt6N13Axoim8SrpHhIru3ms8pwx2YBarkfyzFwQkym9dQWWbfBo
OcMUKvchaBdAcWV+ykXt4tAsF3a1QTYWDnZ7RG0BGSlIpcLmEvJVnVn/5yjj1N17
qSzfqzJfex7FY4aPixBgq/PWi+LKB3J9Idqp7YQiQGWQDavhflZLQJqOYaTZcgRC
93g0nsP1OmGjkuy/Y5rp5Y8B0y+NVXgbqtE9IJzBOAUqyyXPrPOuSlJklHP5vAyU
/1dJSzqgzPtTqWLQUIqKWYX3vCnTqwqwrsMiCvX8FUy3+7BS6+RYXUBVl+eNPkqC
qObrR1wzEDeLV2BL0gOIvq3dOwkTC0vQ/kPuggeOOd/hynRWKfbspW7gEHA+VuI2
21/cNGOBVXWsTxFJt3comV0+Awo/tbGYJduEGRJ/Pd975Kml/GOE4+CvaAk4iWLz
ZoOToTNwEFnEayScIJLLtE5PBZQ3iLtSDJXMfDGFMJc3d2VEbtFL7PuAKsbgSHFk
NFn7vb6+f0HIDY6ZcdgYOu05yGYRoxf8jgHxh00dCJXZ0K5Owpqs67+P4HroQM9k
JLgLEhAKlVcM9T+DN+7OB2qkFNf+/YTCNiiAkbwIA4MQje6cX3DQJWjjyVeVhlD1
HDEA54aTwEuajy0Oi46ibBQqClf0hLITl2jFMmwdqjBHlC9r+W6n4gToltFIF/ME
20PSEKbSFUONjdV5H56S80byqLEizXigmEdNc1mh6UpFSfwvayYnlPf+MqyUGmVL
hwMWl+YRWqPbND1e8C9bo62p57Yap8E0QWx69U58cZdrKphSuUY/PDtQ/hXEmhAd
j5/iHzfDzIFRSa6nzMPC4GtH+zn7yBGvhZRo0H6tgQPFLQsKOR2hltyJTWMT1Qps
6wmM6SMWy3D1Tdk8c4xuQ1a5+ROqMn4oL0amyGL18U17YdxX7C02A6jfdm8iCMZK
/CNA/7ImyfGRpAzZoCBiPCoioTbqxL3akDDkwNlPdihLpHQ3v6oGlufR8JzCBqh3
94mca234Tdii0qeXzLVEAzveGz51aortSyrTmm3n0BAhgIKJ4IkHuUs6Ju0tgI5H
2GekN5me367C62Mbb0y0uPsqnMaDeUZ3/JQ3Bzmi8nrAdjCqhcEhRDCRdTui01US
Bag9lQqQdQfDSInFh6WfNLIBr0675/CVnKtbu6CC165RxUPc10GdUPfd1ijcbJ05
jmAjNiYADkxn3Gep+9fif1UEFuVmHDm50wC8702v8PAlcSwKbWZcvzpwfZm92ba0
ukBHtEM6J9V1g9rXFOt06EsPaJq6BpVx0iOCoP4BJRcBWM7aczhlK8dncDJnlD9p
wUQReiLjJ+CwAFQtaZIRjFyQ8hGrmF4RcSjzJ6bcOZ+Bvysx4I78fkSXeJYeiR8p
dIRDZ3Ct0GAdXmRIOGyf8ejrVFxkEh5oshcPmBoui7ovRMxGGjii8abihxp7Cox6
hFx/d07qhW+YAz0deHKXLonoM/lx+wS+s6k/umRKc21iw0Vhf4r732Im1SXo2+Db
QbkJNvPrJLb5g9TK50CEUDO4T5/IvSARZ0zJHw0sNXmuuw1Z3wPFJx5/o+10AlBU
8DRtuHDkV2CpYTR+85za7lB0hm8x2L3uJmBGQAbpwRWfCXfrZOvhASFE11Ttb/pk
QL/25yY0S/i59xFORXlubVBf+QgWGSYAHuYj4MIiYd6GkOwGhR4nWhm0oRGc4MdL
vKAjc1KH7Yhd0MhysL2po+It6zPrUfO8g8wY2znGuJWSIy6YupTxlULwQXhQtYDJ
5ZiGvW/lZ4XtCg38ExQYcse92Z2X4jGD/x/IdeBIBmqzZBKCeJ9Uz15hVz8bVSRi
p7U1PGfqzZof0FE5qzqHPiqo/ZbmhO0WTx1H90j+kVoyCC79rwbom09WWGNrRALQ
KAruOO9sKY7VPaPeYeAd6xz2R7lejpDJVwKAmC7eJLiicpnqRHZ24VjZkpAm+09H
Ohl1LluMw5Q0TCHEv8IgSj/rGeVcAl4bi69YP4TO2LsjKQ/bCg0EecTbAG78f71l
MA/buL5lCzQrVBB2aLl/pKDNmJid3txXtOY38KXB3DijioAvcM5kXYknDHWRRAN+
f8dpha2iz1FmlluQDawqayKXGdSFXOSz2eXw65KDn9fPko3tR3d2z6osWzr9VZtI
sI1H6UIRAX6dx3tj5b9Lhc0qN1xleDP3OTEriVuMu5rWYtOn/Nq8T5J7d6K01c26
jObfvjkCQjc9hqwyntaExgf10f8X+2Yt6gskyCKaENFrs13k5tQq2c1UcYxgmzcD
tzaUPmv0vPifsUDm6Lh9qVT+RZwasU58mGfBx9WGiqSqnqfXQ92l3qOPAxXdTbDI
XZ2EAZh/pDETb8QSJAjDWEboUp7kRZiiHUe0M/UIBOPsdfPUpnEE2Czd/6djeXj4
S+xMynUYj02JwOCsE8I9vfxGnCYdDcylR/gepapzD4flpukL9T+KbxSEQ1Nt7li2
08CQGQbYT8BPLhYQnLrMe5DjVMFEvR+1ewYL0w4tj3uS2bk89LaOHmjdZ1Fkv3iH
jGyOjhYOoP7nLHr/4TeCGZQ4VMWxkiWNmSOGV9u/fmtjQ0mUrJD1aZrzIwgVtj02
m1kACOsl71NZS1PZdBcyJSJ7vN/ocQ7BGrncELadttolbmdUcKc0M07NfRbGZy5V
o/PMkKODaRVaZRxYtO18XYXJSMihER0OWsD5G1KAoGzG8ZBikVQ6cltFCtV2N16v
1Bx+Tv22QvZV8fgWjts/9PYZ+cAA5UR1KgbnpKFBPiX0nmhpzm/JPXyhdTfzzOcb
FpJLVTlhu5V9jmdg+scnN/qDn8NdxuqwPewt6XSxCUWXAp/TxLl8W6aYfgc7yQB5
mEwF/NEwNEyG2cEe81Ldt9AsGncoc2UqvAkr78GgoNW2NA1c6n08ku40xgwxyt46
DVVhjpoME5rJ06gbaqQydPVeA5d+4TkYcyxSVhNWBW2MWgmuNyzGbHHVB/44AOwc
RXZ6ZhnX7szN2YNpC530VvLceKiAt7ARz46OyL5BmPfZ/Tgq/GJQu6iNjuHRM8Y1
B5neTEUQz4268QUiox+aL09YTJP8JubaS8lNd28IDqJTJP/6hJZWRtjjrt8a2JYq
5f5ytKhXtN0yYyK7rwZ7GFDhJ3utdx3qO1N3daaa3qNGGYHKVbEK67pHqZZ4sIi8
G7KOtTD9ZRIPXfoZuLdXXzy0iJJVZ3zdhDUCZBiGCclBzzqlfH5PboiaGBZ+Wclu
5fa2uTxKKLVrqA/rN7Fv9RckK03yyiGLK20/Pd611ucNyg0OpgRa2MFml1AaAu3m
IpJBXzkxzUnOr6fvR0Ua60kxiO+YtujqkguDwLhw1iZ3blhg3e69n9UHeQDR51YP
fPnPmQhydVgcCswfQ7Jelx7VFH7+t/RsOfuNLo12XYc429HxeOLgnQPBBluU4PCl
c3vMhNUKMfaGsFsGGOpuNU4hwggayg8qgbjZ/vbvQ2J7P+kGIQjOrf2Zr9oldL/a
0c4thbluuEV3SRLdFVmdpwcALHJqaJoTVv+ALuosHBNqG3madFLK/BeHqBksg3UJ
VDwYZoNG3OC430L0IN1f7XNiOpfl1tDD79ShVwiTqn1aqO74Hoq58QPfD1nOUBXB
9TGu8jrYpGDOPefbGI0sqlAIb/pNot2iP8r+bHbefoStvjjFcRisqNuMvmPsVX3p
4r7MMmNBPwv4RTn/u0MqQqaspG+AOgo8rxKZKz2+EyrN5U22VM3pDjMUU93jbjdU
HTaHdjTPI8BCUz+ttEpVyuUXFV7eouDp35axAFLtihVT0GPugyDSJTsj8XeYyoNL
6mg2Zw986KnxIZZ3gQHoFz+JeFsLW2+dm6WWOmr7jgEbO/m9Mf5Zus56XH4+nDKQ
gpdAGdt3+c7Yi6hAtlAVWm8KmaDzO6GkhIULBAWpMRyT/sDkhk+/ZdQDfiyFBX5K
NdfUmKlNyiJQGKmzjI6310ha8bruVMbAyTQmoM3v85X+vW/UGrjEx/spnDiJ9Zxy
D5LHBg/X4U0D/pqEdTtUekESEqxC8Mxi8xyZWBoG8nr5o3M2He9KGPFKxzOqNhWI
/eTTF88TKIU1R1W8Ie69Vzh53s31kKhoCZcHDBBnYNY0S6TopfkKI+CNMAVijtpm
vWRnGJWqMFoYDzo7EisW1YpWZauhgxPTzuqwnhHip3TNt4xFyj9Z24CLG/5VDZt+
ACXZwLkgrryLEe7PHJMIweLiY7t6nRk2AyXoMmyHm7hm230hcimwnmbpU4SETx0M
mmBMZgeSMUNiyvH/fL6OprQBKbnGxz79dm150kbVkxQoHoJiPb/XU2Wm8bCJWOgB
y0GLX5ZGJroQJ6ZJPNenA/Ao+1SQA0ZciwPFpEeDDI5yBtdkT+Z+yUmeNP8RPVzB
mFfYg7QAj7qEa7YdRsXhonS4xWqPz3oslz8QJAxM0YHj1QQrVVecCMitP9bemeoK
XWl2G46AiRmW1Z2KqrEhKaTMbpeJLQnymixYs4cU38wFEgbxFdRyhtvxLZ50eSW1
thOLVrWzc7OWovZ21jZh3Ac9y0hVeuRQX9etCLeER0aFdW1kwT21vl5U3m5jDKjw
x9GoRteHV3tbzvjYNIIiNMFVDamf0gtMe+LJwRKjeAZ20yldmGb/NvwYA7+RL0EY
qMDp7OiYQNeAi5XocCwQUeSoxTuT+DyextpWkMFPuzophSZuQabvpnDvv9XD7i+u
w0YGvvtXt7cNmE3BOKlpVqK//n6nRy4C2BN2ITbxwo8xyV0ceL3WDC7a4d1ew8Py
65EEQNMdW5WBFGy69rSvaUivxzdDaDIiuVq04Sgf1WK5WSq2bMsIxeWd0xieJiLD
HPFyVakK6nEixauy2SceHjciaDDnPtB2N/1Hkb6XNJ555uMCQI2KmrA9tTdgXkC9
KzPQ4m6IMevQ1nOzP0UW4/WkBkwL0gkBnUUy4PhPp7z1d1KOY0vzpdu2tACyfFeR
r76fOQ89R7WgySgsxD+1mQCjJSD7bbQf+81/YUHtJJsXv6HlOKK4fivhKoz1RX0Y
mMrekHvw8FZ/hPUYvgwhWPnJ0h2UWNQi7+FlUtM79PMTZnMbCwJ6Hnzjr33RpgL+
1awEvhqU6Jb7/33zYQ51ijVaDrup/TK7HQbS++LuOOhhshjrGYpQi8Wf7ddxDBWp
UaN0tfk2YENYcCcdeclfOQ2SjyINbDJWj5+q6KV7gim2uT++XQk4KR6u8mFurZnl
Ik1PzgCHE2mvSaoI/J5OE2B3//T5Im5EjoXHVObNz0dhgj2ptHcpJfwM+QTJQCQK
hYI6775svd+k/PKo3yZ7kY+pTfYcFQ1HvZWIu1nwfVdDjbdopUfU1n8kD5c1GnVV
WMBUYN0k5wwEVaxInSf1KZ0iDU4lUY1+Qn2QKM2PjRNTzjz+Cgt70p6sALOgStWX
J3RlkruGg7OGzJxQA56u2PvUlCvuraFMnlANKhWHXpbibUWCfGQj71pU7DAlc4BU
od+5GzXcFQvYDjg5WobfEP7Cuxjb6jNRjhOQE2XYvjAurRCz+y0QY4bMkfB2ffF6
qZFxNs/oXc6SEaZJLycptJL0Otg5svMiNsYhee/atCKts/jwrE1DmU5EyHxr3NeO
8RBUv1Qhj0S5G2gkXWn3hV90vyvIW64kmu2bvqURyi7A+nWxbRFTbRcuvRqDI3bO
FognwIwdQU1SRwotKJZYWOUCZo9vDle+TbaVf/ihMyJGRJg0nJLb/i8hZ/l7B+zR
QRWCKGu/ZZ0k8IKzmxO6u6IQwRP4/tv3/KaubD6ZOuRojJqWtG5wXvigx+4fOSOx
0Tp9TJKV33dOlO6TdWxXiMYbhhmQmBXKo3XS3j9yrPmbqzItwfYcowDMtjyCL2bR
eOLdoEFQ4a6szoBNZ43sPJPNu05NrnYUGu2zRfWLdoW9OGkt339BzHVdfT/xHtJt
cAaZDvOf20jAHF1BRrsyfi0a7x47lTR/jh8NKdu2+sIgOFv9/h9THVNVZTocev7Q
W0UHrLQoXkbK+c3sJJ5k6zMMnCJP1TQaC/to4UTl6U3XAhlu/wfsQkN9K3mdbBFy
0pdInlQ7Rw8ptnwrLioXAU0/X2sgo/AD5YASNRPIn8nXUS9LHe8O5y+eiR/gnEpJ
FN5OraI8Tzqg3w/NkIruHAfiBNi2biZMQrgDnd+vzUc/FsJepHFJlSsv/bTc/iZs
+AbDBczgvqgwW+m/KvPpSM4D9p2dPzikvAibZ2IXatdkQiF7KB8JtT0gntkY3VK+
ZeY/7Rz+Xfg2e1NkkhHfiGiGhmXrq2y8mzDTkVL3uQES7fD6nelYo1Rf4aJ0Y9yD
ZKSmeDFPuBBLS7524r+dbYPJBxW/AsZIc3aoPZBW4cPwlGfoTkGl1fgdLEAPTCtv
BsPx1t7Vzs+KfIYTUJZguHST1QLe3toqpH+gG4+dPSAT7UtNnmX3d9aS159zLs5P
hIj+ocoNG+o4Bt/D9i55wBciLUTHlKbkkfVXJcA3m21XbeCKyZWnzMJuN/iFrkv0
PXqZ9gtLt2+EdpK5N6nNgfviGNTihOCuGwGNrb/x8hjngiumwA5WSMx3jid9XQqx
pn+qkTj2CeeprkknLmDTSTwK3ouOAWccc6ykYHNfJ7wpgvHgZ9KhALBxu6czqjK8
kP9CHCXVWVETpg5TxyL4Nhp1pZ9gFn4K0zEO6cle5ZZibp6IrDV2gorqCbYBTbxO
p94SlFibA2ecIYF+5ysWwwzFtYDJOoPwuAng9952032Jyt9qyLhw4pQo0mbsi79y
r4UHnT6qRnsZ2Kl579oon4ZIkSRaZHvz/fas80APXQohwaq2FDbADc0uhXg1yv/D
W347pj94BPrPZD/+/kRMoZsCdfjIXvo9hnxZleKxgPBjl6JIRMznkNRkPUOzDMz1
SyzHtz1o48P1y/bIPPK9Z/D1EBxUyafCHxd2zEE8trhZiHz7OW8Bj9iYGjKvkAbO
Vc1n+ses1vihFajlkQN5RHcPR3Fpq6HJ9Sg/jrdFSASGxhIVApK/zGrARvHOhaf+
sdd7YC01dSDvrxg49j8c0tN37b+/2SLRPoP2bWMcFsJEw6gXJ88aQjBlWPD84ow1
wATu+zFajR0ex+vEVicsENL6/cNbrGsS2aofEI0Hs1WLVQu6Vingi7TkhE5fs4/b
kBvDK8QwjGtuFERxjqMKFvlHabio0NMzYcbhv8M0IEsfeO7q2RCOwv+hN9XK04q0
qF0jMkojS/BhohRxrA7MnyYcqOKhcCMRJPzDGTqNxIS+CwtbdNS+t1B3WrGT+xsH
XLI0xYmyS1GDNmnjHuPCqwlpbuxsYqzFx0I+1dl4zhLgC/FLmI2plQQUI2l6WIOi
2NcdyH1YderQoXGV8wF+e+SbomzXvT3isS1mpWPXZNwQrgUk6fwNRu2czkNLAWl5
aM9HBftTbZhkW0UHqySE1NaGnP/l0deUIqOMH+dpixc62+hWm1Pr+R5gD909lrHi
JtyA6MDzrD959XacUPpuYhnHNT6GVNB+vjhX9ciybIlFCLH1ty//jeIhz9pWFWwt
MIxDytsTJLW5EMcR7V+L+5f2ajXjhPy4RhN+AqxUqHkiysj2jnbUpF+oYGz1fjRt
Bf89HPxqDi9ll8BiCJQ45k9zCHOPJY4kLr1e455V9gTIeiZKa+CLzhiVwno+Em/0
+t2OobSxmLvlABPRUis1Yc7d7jnpEiqT9qOA1VU05YkDrnlScwxsesPCJfP4CpaZ
4/NrgJdXogIHjae+nkzsNAdo81XDch846CnfLSVHEc0ioHB+deegcAJ7jVofj1ZC
ZaApbmxYlrLk7IN7OYqa2uzLL3CtjWkoU5zjV4IfCjSFb51o+KgAUpdY8FzIz5IF
WkrNNQTTo2umCW8qdt90Br6iKBvi9favJpbmB3fe3TpgrVAmhgiJhEajw6fScF9l
bub0IgN7dD7652dPV4lzFGbx9Vs83fnPaLGptAc/OE1B0jmrlPqiTCc4nJy8/wIM
CPPefw4mFUPqAIDxAdbES7wLCTc9HSofJ4D+HHkJ4BdgTDxyHJsn9vBJBmYjnZO9
7RFnSqHj5ODF8Yj73bHZDVmo2KRRZiNkT6/VmDOjJfJRQF9LyCdOEFo2kQeDxmGh
MgZ8nUJywNav/WJfTTWV50pxYPXMF3pOAj6KK+iRY2nx9NLrNvtQlMd9peDWv85t
r8/a82NWLwR6gF2MRe0nGoiww6JOpR3qcU7jmrgKPRZSVz9k2h1cYc2cg7WwwnTd
LNKAeg+bPR9bsF44do7nigULd5UmbshW6iBbuMAZgUHksXJiMjOYgv3EMYzh1eDq
CDw3OlPQjgxYG/OepN6EMO79CXne6WhZoHIHSCVoiCzn8iOizRHpuQiD6W8LVSAo
F0QF14arSejUwjMar+VYFEJnPcAgQGmMwNXzbuBPqiLqJ9hcKZAZb9kyVXyo4EV6
4myDpXCd7/o0RyhZm8XXIAC2OGN9mz/g/VEGD5cTEusFVEa+lNgfI+pkpsqlZGS+
clxFtJfSHx8slHW7PsYsDuxCi5uiO7Wy6vkdMqdygcr6M6lgSag0FzMWGhLGwneY
Za5hJrr0d3cJXoLIN8jXnnA3w8evxQyGrM5pqCswCqQ6wXzyIBOV1PdbDBMVLLWM
1b0a8LUBfEDdDU0rbnJsSLrQNbX/U77CIei9l4d1v5NejIakYchoKBgHm718nykw
Ec+xjW+A9bIRlJC0EoYu+ksASgBf0g6fk11Gp2xOGxmU29fOlBxtTi+dLogSMVpX
EaWH8mzMBVZOXI1KpKH04ko3krTtm6zNcyK6Vb3kuNp3EffgEYR7lBbSJ+VVO9mr
SA0dyPDZXYI8DiSBSZL30cr8+ljkMJ0SNihn6TGZEpMjrlFuBzYWXJJNF8YOUuVo
jGzgjtbv/jOp4+z860M3UykzwoXTusK0rKLu8/IWueuXgxYusTRtWq3gXJB/6GLD
gFkJ4mYGF3MCXmxhMAMc92VmwPZuMzbhKFIgI6IAH/oHZIFfGykHNbglsmcAgOJv
x3mOs2JpHj7x2EPL3oVuGqL+etzyzcOGTUR1NpJ46hTQZ6BsuG8T5i7ywDFOxnBR
E5x01kbhWp0j4wwIboAYaNgp5ho1EVYzIeGaEgdlTtcopU6BzUXm/0ik6k7KZGka
pNgchngn9Cy8CueaM3oA4QpbunG3c4R7UDtuQ2HzUuVnYu6OCiAuCxcUNb6gcqrk
8k6Xu35G+9kn+cdfwUcNFJbqEoaTfknmyBtqfNqQ7lYbhh+jpSyzlavWaX9RMGm+
Q7K+uz4c288l9pQQshDqXicfTH7y9EKck0Pq8UEZLSZccx8SU7TXjRy2z29SjPLr
n7vOj1juZrCSEW6my3MDf+KdagD5W1ERlZ0pSwE4VgQjJH6jMT0RLfE0qk7/46yA
tU8K8Ll70iL6ASv2vX7pdV6QLGIjXNotwHHcT5tljnHIrpq/1jPz/5HI8EY4GATV
RnrmsrR7EvTZ2R1xd8mUVTQqHgJj4OlertqSitcL1JkGGTxczxQv3NHbxruGAPuB
fdRBJyicB6SHm4u2vTU3hLsHJae96iKIU7pFTbZtAAt4l6VA9ODDPz9SYdCAGJ9k
8AH4cljn38M2AlVXtBepYqnpu6d7jDGj552OaF8VAPGeSVgCviWFUMsP2WQBYzFn
KMkIOQz+HRhegsbuOVbumQycxZL9gCbKvagapESLNuaZT1shEzrW+E23vH2FrhAh
n5vGd3Nk5ggJXjXLEL8MFLfrVbZCGbW1LvsUeiD7ZrcqlZv0Jd9pGhEKckMb0sn6
nfzvSZgbgLqox1fJBmnygrFr9GmZIJ68DC4GRYnv+aoa5gMO2EOXWQNct38Veyrk
lES7CBJQkhmLBDvvAKm+/QMHpUtt9/iiD/Qgnv4lALrO2iFHhiMwE1GGx+yYzxNp
kp35kVXmQDbXkiJwBvHcH1GIIfRy6QpuldWuYmwFSG9g0+4fLFtOiM2CD0RPlpl/
cHGx8BfdL85LXpwojOtA6KTI1JWVZANqqBPaMWL9g9j5o61ySAjJW3/TqcUzQPMx
Aask3Uu31v5RlDXOoOcJ7Jf/O6SbtutYSZz4jSjVOJYy12E5xBWNK9gO0nrOrSx0
IVtjc7pH3tR84HcUoaDffA1RDMnJHH/C9rUwcWGZ/ZkKw1Fpt97LV1UBIl5MP4WP
kxe10Lct+NVP26hKi+ND0pWLCnU9QK6g260uL1OK2U3Dmvwe9+d3ujPh1FCL4sMS
2SnDnehQdCjgX7YM0+9ibd76u2r7MpJW9q4GH7NUEoxqoO0X61XcqCeA9SbgLU3+
7wkoXBQfsuAriRWK8oUaOkC51LUGcuaFD9duwmq1SSSHNqUcMKDhScxLJpYQsRe4
G+le7jegI1tMaeFQRIUOQkEVALSCc9W7Whbxcnw56hgPhDOMDoiHW6mePI1n/1Vj
fTggQjRThXZ7RhUlWBm69WKUiSeADrBal9nz6f4A0Dcd3gSCbLOcw1dZ0xNAS07Y
hJoQJX35M0deTWhDLdXEtQpWDgjMznSyQUPjdlOin7ajttCHDtIqIwCW3G7fSS1U
iWL+pZ4K26yhIzYV2ppf+eURwB3TP/GO4qT8tF5foOrUXzkRr2GGLx4q5NwoIODw
v4gyVMQHWztMkZRYz5DfQqKKJh4If+OxJu00XPcHVTOWZp2ulzaa7s5cC0z63FAa
quxPBRoRGtCk8ntNvbtrrGR206ZkphVNFmnShX6AWjXeByug6nT22HL8Fak3ezOO
eYQbik+a4oEB+LMVMNHsNu28IxpR3gzJCAwgPm8cjou6aWRa0FL1CyObz0uInD99
w40islYeW8j8N6lMJVIRYYgY4eAWRCFOafOTQwy01Tyz9zem0GIQbim3HqnhSa9C
vVf5g0/kohkxapR19roAUl4Kn/CFnzyAP+OZI8VHjNAa8c5h2ya0lLWyXF7nVsW4
+2OqKNOZwRKelB40oy8covsLscJhgIkiwvx70U9cI96dIesieYV82bcwqXEieNFP
a1jZkQe2Efh7E8uacR5gJxAWgImAqwQO5u/R1pRp4g8ybY7jwpdKya3qFhK3YhlA
fiYRCkdnzHyuUvpEUKn1gHSOgwHecjJrUG38XshnN5A61R5j5SU39z2oEuP1QKC9
gF5WlYcfb5EIIsfJyeNx+W9Uhv+Up+xaS5WKUL2n+hKB0czT9f8WXS5R9uPfqaKF
rsNKyjVnuZ0cmYhR0wC0+2WAPo1BcmphEAVclncuIF/Uvhi0iu5LM5EzvBEBWkyw
NCV6kRGMceCrSD5u51hAmwHiFDbJ3lKkkpdykAXf+V3r3tCykCGgA8o7hzRafqAM
C/mdSQXvIR7ZrCg38xC5EdiA0N1916sW+3TGQIKMtGLFwjNjOVLEu88aeaL9S/sY
3N9BIRbKQi80lANQKjxYD870ZCFYbYiy8pdRg+wQ2CMrHidY/jPrwfJV8fvcuEgK
Ppg0Kwe89YiQ5hAAnh2SlyzCaV9//g/0aDCP5X4aOLC7wh+R8wzWWgUumwhuYGp3
LT6LFxiTuU2logobgYDDHQjtBYean8bc8WoWUXhcFd9AEDpDtguyTbstSr8J2OIw
xsCv60VZk8NQEyRsU6Hhga9bkVH8ZdQOhi1oyM5tWBCinr8GWpH+v+Oix0wGWBMB
5vliuwcBLSXXSsvhXUJzFsjcdGYGjCvF5JzBCb3iL5+FtXldvnfi+OYPQBccjDDX
56Yk7o7wuF305P1+oBVPdGfJmAWkrhB491IYhBzqtADqqBNl4Fn1NGsqJcMhjlkd
P0Eh7LdbHqqxbIVl4QI7o0EQnJmIkR89BaYhi6zoUGt6fTq0wRx2u9el31J0a7hL
8LWEmOnUDLwulBxEC7yrE9M+FWkmSpv+zxvjk/lE7SlOcCdyM3DYM7KK21VAaghc
vucRtGD4Zkxh2iww0sI5igP0FTgfBFbgAl6NKg4ZCX7TKlG/cTGloJx+ZrUOvgbN
3nWctrgFy464vi6nVXwfdrSe4VVpUyDGdFiqdC6oAlXIuTmzBhzDNoeIZRIEtCyP
1lJ30VgxzmBoV7E9tlOz3KSHrfZz8SieiYVIaf2ThLuqjEUYRW3ilhMoV4KqpQ/P
R7xoHN6XRBFkfPyNpXOhM2c67ycuaxHdU21UXK7UROcuhYuE152LbYI+Ah8MISPw
+yLPTzgCrlQSArUhLwvDSAG1YR6GzM61rDykT4bSc8+t4RgvzRdBsbTu/G4JUuLd
RyqbWLGq+4RZT+mEzvAby9jehVI4ZpdcoMNx3/lzDbbFTYIFBgueGXfSqIpRVgSh
n71WK+ZeM9VKc3oJ+9yr11bBMqd73NwZL5TxFG/Z7xMjkfDPxxGmb+StZveQf/S1
w6+qZYCNXOLbELwlnRXyvHRShJFXO82n6ARhUkeB0ikMluGRi1Zt5evjClsRVoBS
xTThRhxrRoxof+xXI6bq0HyYIhyXs36IzsxrDAa8NsXnAfKxtUMGzTnX7o081m6u
iwp6319lxScR+S5S9uevQnyAHCun66yd43ijzWgm0VHzL19DvSJ0uQV0+9W/ZYuk
eyCcCoHW49uPFoiQIfA/kj9IKKuM4QZ9z43XC4fLGLPUaw1QZr9FcdLbfD5zFWu1
0sgCFSBgVc2Z17zjO4inhZRXPhceJX7RWigOEkzbqhS66qxd9wGsSsSPPMmVOzxG
fnlsIaEV/ymAeK3zIaMAMXphMsr/M67FWAEbhcj6UDxrS2QF9VMBw0c16YVEcctg
2YUrMmHwJa/V8O3ESy5qYySVfV2pj5+umnKIJuvcUexPdLsheY6c8YzgeP1FT55p
elBlzHB24V7oWnxSkhGcPfVfG7xDpo/pBSwBaaSrvutBlZCkJgkhBTx2OcnAtOMd
Pmp1qo2RW2XSKc2AnPe3TdXOKORA7xUx5ZAPK1Aa4KicxFpoJ7xpm8efLSDExXzh
gZc+Ge3MVdOBfrgeXnyAKZI2VdDiXGaxeVkJhRW4QoLnsYOBerOUR7qi2fAsNSdq
5VxlWqX77N2ghXMjduAyI+iEJVu0m5PisT0Rqd1U7solLUHS48z+WcjUtTPnqk/i
v2dbBZ/LmFCekqO8rq/LyYHe0akIo1yivpZ9DK7iEWVV5c7PYYHoErahSH+/CY5N
n8WFqY19pN345t3MCTUYAuS69yo8AMWJKyIvc2y4R7hm1IxLjVSmGiMnXiEy2kxw
IrsQSf6WsjgqI8q1DEF21MZk/mEqHteCBdNZ5b5SbvVAK68EFcGD1wXobbhXCvwl
6sar19m0nrZ2lIiMrWSiX6adYDZPcnkhJJX+xK54bjTXEDsa4yBxBQ6a3GyVirmd
CfSOjzCUEkKSmCpBOlIqP/ggQ3+evsuwZzPyFPTDY9/hMN3PMCzVLrN3PGnjftLP
xaWiaOPCgFTaI8hm5WXFS4V85BdH175VQWz92CL6NPw3RATvMTp9TSs0JE4mOQSh
N9ct86WRUIU2+dAvc7yp7OtAR2XgiL6bBAHJ5AuT5yQwhTjKQ3uT6V6wgkUl8lsn
bSxdLYApmhQAFcmnfXiqC2+zQ+Ei87Xz1DLPlxm761F0WdZVXIesi6Rw+p3DuBmr
IR/lxrhpEXOPytOzTaWjXwWq8pB+ovOXlltnyCzHBwNV8YnH8QlG1hUNG+MYT8Vb
yEWLL9yt9sOyXTkc+10WRqmVEM2zR9xFaP3OKlFMiKKBBRa0dhGLszKf7jn+r0C2
74tJYGKrh/HlS3nRUsemoCmkf+6FlRRb89vAIyPlRIYp1xNSVjb6lcolMPCibglL
w+4NaYofbtN6M7KgM5TFWNWwU7A428VkRap3ZIMySFdyYTl7WJgl24PHh8VgjBr/
R4WK6Esj7hhiHPpFgOJGe1Glo9qftdcGLxm4m3EGyP7EJuzrKOUGETelqcUNPPON
ZQBJDDOfKl4ubwB66lnvEAaPO41f9RwnOB4U+3zvn3/h55MdoOuv3a1fpOYKiuKX
XqIt8uMMgc/PjNNluewIn34k1xmCrQVymp8deHsL5Oi+GSMkYWLD0gt3baSX19SR
aMHCi+Di+neEsivYRhkwT7tlUxxIqEbmxJnjG2WppTiITGrxnIaUuU9NHVFNFCFz
tn1dboabR5RQKZpF+x3xLl6RnYgaQ87/Zg38xF3Rp6rEJ+bQMEcd55An8kLCnZqr
ByiIk3u8A5DVrINcNJt/f+4FUfQKXF1ZEYJa2dFkHMTxMQKpPgx0DHE8Lsdq2yDJ
XJdvbpT8N2Dd0PRMyMEiJ/0hcIqUMeXecuuJWaKoDy/FNZvxaFVDHM6YkCX920Kf
xH/LNf72EtO2oXB18T0nj9Yu/BqXJ7zvvySDLrvsvL2F0y0cfeqeUA18SHH9ksbZ
wTFC20GQPqBTzjhVkZSEmaTvn0F9UCxu2VtFazIhYdWQoln1BZexlGP7IECj4hqd
u9rNIs5+gp0fzdpEzL2Ru5Y4QHOhzZu4K0lVEF2GTxN1QU4MPJYGnVtR8u8QHfaS
ihmmsqWyf4hVRX7W8+wXLmKeNdzXW6O6j9MpNZc3lPOzD8p3iI6VwGRNe1EnzIeJ
KUSxJXqODszkxS/FLBCButYn39F2m7L3Yq18eIty/Ngzi3CSX/Hx3YBE88dMzuRv
CJ5wVvi5FB7Yf/gU2VroTGEY5RGiLGCN92BsfJ7WntcjNTwG/JjYkN3MfiFiO77w
9pbjaO6OblM7Dt8CuCIU6oE87v713zh4JLj0LvumVWytsSaXyIcgzw5X/uyFt6KV
2dtFSO0XsAoptvXYH9Yozvbd8q4N5Dt/lxgFyNOL9DkjY4wj6jMmpn1sLk7vHevq
ycibxmUa+6voRqswN1ouIaiVMvVBibeHZde/7Ki2uOvs0gNgZlSi1babpnfluaLm
xhDwWhHsbjX/d8L7LE/CHBmZbilQ+BpdGhEpHKYSFcvl73LWTDdQnqGROGgJz47m
mTOYIJjF14FzqXblWZBB3tR4mIy+5o81AuTL64zY/UWiA65VriKMLC/i7q6G+8ru
Zxp0NrPlIU4iBNk+WlYwPunD7oMrtVHaEKp9NwuzlfP32mjn7GU/CJq3I6G8KOFm
agY6LtJtW7lh3/moZq/uNociPBeuWh0BG7lMJ0fxQ83fkmlxRJ99uBtG3RWSjcDd
xUBfSKY39kJr3GBTmC+oZPchU+Deu4XuBlzJCLitzuDdcM6XXErjgSGJgEliJ2rF
IGlOjv9TrpCwWZNM/PJIWcQyL0V4ZduAlpa8a5aUuqrPpxlStdUm9yR+y8iKXr1H
B4x8Pi2GT9KGABcB3ydoB158dI6fxBVuZ2kUPctlKffFU5liG+mEUwUjwR8yPk3f
oLl3X0ojLgdj91xrJ4bCz22ZvlpbLOlU+Be/fM/osTBmbejFcXXbjQSPCkM6Q7Au
p7KyXJQ+M4eu/HmFtzIm/2ZdZ/xGc8uQ+YtEm+BYdK2KR3W4X4q8i7HTBMwoI0jJ
etBvBe9VFMzUoHdOfyZLi6MqVm6EOavWuj9+q5LmXI0KNxpJAc3mqt8xfDHt8u/O
/jBbynxwXFyKA6tPX8UvlC/WNGNx23cpKlStzKsk+SMuSFouHfzxB8zNEojYRupM
ojp8gSPrLP3f3frypm7UD7lh8mGx8jFqURhecMqTtSru79aK3C1LmP0M3TQDXFL5
12F2KM/+/9OG402ihwcuf2SvqcQLKJOvCutgaEquhxfmjMjy3Ycdrzl9BeToKuNN
yzCa89rhl9OHw8dX7xe/O1kJQ/z9fp6UepUp1n4wx0VFK3zqhasXJyYRHsdGl6Az
RitPT874GZjRuT6tK+t3S8DGzYqvKPPU8u4w3B78JixiuE5s5Yd4oGxrf8F4yTwf
wrkMSIVWZ+lOWjTlfAqJx6MN667NZmuOw+aDZEZ3i2PYWV+KCrlRYtie+9o8MK9f
HwI3AvjRJwQhZovRoCwqFvPUtwdb6v2ft0V9/t91vz82tGW5feW8g9fqyayWPGiD
wH+UHQBPAM8Q4X8+U8fe2jsM44q805IzzFSEqTWnci2RqlPUFEmri1KJw5kkbhlh
Y29/bfPM9LmsKa3phwzRLDWweMvCT5BJjhyzoqXAhIww9sNnFzgAhaytHMALKJ0p
xq+Ldjl9sKTiLxv7LEq7bKooCHldwOpSoNPFeJV5SnUb09lSm7octTnYBvySdLab
2CE87cj8BIDgmxo39mcwNyrI5J/kxqr6cB+SQDDrdxBM8MVbUgsn8OHzQiYCEXWA
QfLZgI461mizL9KATZmUyo37sMFt2gtjT2tayDHzHHJIDJ9dHridKhDL28v+vczB
5RLVvtkR0stkDBvPkdeVjKQuxqtMIg26XR1IAx7XzvFgiZUWXSdIgLA+Gd4cpYfF
KmCH+L6aM3a1AuPoUhzIPuKBAeNAPtSF7Bmktwi2ziBxTapQjN3XpVVd6vzpjp83
DvqgnG4f1zKb6K5aSXLMlmjRWpPLxuNQaFYTMoUesj1qYQBsjuI+IIC1mQCTu5pI
pq3K5GBYGhu0ZSoq66vV+oxAVJ567Q7eBZGrenGmR12aLah8NJBez3kEMPh6XDip
mVSg+ykWlAd1GGM4jEjxYrr7kaugr0uTrHaFahQxC4F86qDqZIMkBLgNslIRicTs
WGvkOOKLbKCabwAcNovY17hFz3tcblAldGHodBOtV28AAhyvcHNTKFFLS2miO3G/
TxeRCpuXDENzaXRHbT+vUDyKKB9J87jOZCZHuxq950ZTFZ3nnTmU+mMXzsUU6AYv
PsW/kBSjxwLr7m5rgTCZrhwGLUH6foSrSH+VEB1pFboUCcba60L8HsQRyrIVF5jE
2jJ2d3YQdXenfT08jg41YJOnXweNBfYR/E6TSZImLGufgWmbI0BSjYJHhqsT7Ngw
IbK5aDzolTYys0W0VkQ+RIEFFcm7/C6wxdurxDL6RagxnSn/D+HQ1JCwO2tka6pa
xMlKiUu4FPz4O2J/69fr9pSVMLALy9Ymb1iUy34HH64zXynNiupxrJKZiYpokCyk
GJWixLjQrA9DFUQWB0X+6HpUT6YlGEGtgdfjd3r3tifCTJhINI207gjsU+kA7QTz
GgZiasofPf1HICS6oTqHhjH5BzVWqCYlJq550Z59OT+TZDndu/bo8PYYI/zWHwbE
3Z7bj96mwwB/k9fqLZWY+7557C77vu0KCRMEqMRXrtspAYzhCt8ou0AS9PJJM4Eo
5NI5MMOOcO0NHanD2l/dJUmpfrfxdYVEa8FWQQn4HAPWkaLH6M5SllBWOInYHBs4
wYwjAun9WV2peWdH22xAq18SexzSOMUrkKAWYRbLmVRcl2rZ3Zykde+yCHjlIzzo
Fynb32upCkBuXIwwCB4QazNACsfcC4lRa6z9oUAJNeGpkqsLYnzd3k/kCG6k0VcA
2oAdc/llvRZLE+2Kd4qJhyfO+xdBw6Zl4wLZMcywWN6UajdfzUW2pjNLVDcBQF5f
9oW7kumETEtrBs882/D+/ZG/m5l0V5zd5wmoQcOZLhVx3BnequRahwMANWuJo3WN
3GPP7I8NT5FjibOjaJS/MteflxMSFWlt3LdaZRuRBRs4VqlQwo4pv2cwk/4uGgQg
5cN7BjD0Yandnk4Xxrh/EThCcp7B0a/fuSHlmSoJk9R8iUlG3CFRheSRt5ZhZv1N
gYix5xI/k9Rn4AHrgjm9tDfP/XVHp3VF6j9IHIdTJTkRYvE/HEmjZrILzynvxDzB
Urn6WxROpKC5snRJq/gwUwAM6TjCw2ncndhCRRnJ7JT6j7+tDpTx/H6g+qx6RLJa
N7x4a47NZNLhi2iF0hTgl4NM09n37ociHpFbC/gRsP9s6JkUBpdOwIhqiErKoc4W
tmj5wjc3JjLuP96a0Epxq7/fNkpB0EZcQk27KxFLBUM7twI789kUHLy3TIMm9knk
gaq4LQxIADGnfgDC1WwmaQ2RGhYaSbh485Uj3xpdENsc8SL25dOkLU21vHi0sNfd
2W+aXVuay2JBkaOn84q2lkwP1Ik1v7H/S3hyPCzIKDDPhqUj/Jx8MMkr+tFgSGR5
P/mZhlcUUhtp348cuEnmzfRgKhjELIM1aYMVQa8EkZmlzPpwuegzAvSRi/tfQqR8
LnJgCdDxGRWJU5ctDZAaxLAm7tImyewv+mYb2b4a8fpFwRqj6yt9cby5huT+2uRW
XNtRMzzAomOlcr9lZ1UULK8Le/DpQph/dxtAZZZdRs/5niTPvTERDtGFpUo3DgzY
l8G1ectc1zGDzXRj7MEPRwbVMgQTiu5qwxJ+4q0bVRDhZ6GMu0LAhmuNyMVzWtDw
9CqIfgHMWTxkFjzQ7O+RsbMq2EnMHa77WRwQwooZHcGDd0JQo10VLeNwOND8Cq+W
6QEY01/rp/VvfXtlcpuBpry15tB61e+6wv/EdLsJccMIObb5AZsfWUNR976Yscgj
ibXvfGyxW5oeDNhtxPmJJF1ru26Lr9FCpNavKADygUDInwUayTlTzmjsVZOxWbvt
F9M567saeyj2JolXVxI3YgWMuyK3algmaPNxcChaEtnKwk9hLvmDAErjCzk9LOHO
o0wozwlEjwWm0kaFPxIq4aQMsxLiEUBE+o/ywZSElYZkpdqxkTCIKVAZ9Uotpw8d
ASFimI3SjTCM9hoEMM+Z6lkFnAKUo8Kiqb1N/csRv/ikAy3Lvo1ELbJGhY7SqXYA
ulxBWS8NsCdfIUngGXH26W3TQBTtajYldM+O7HHVB4wrGaCr90dJM5/3EZbXGoQr
u53D6r9SBIMPiqi19klkBBiHQkoew4TduvQfkDsk/dgPrfOZVMXZft8wKLOtoTsm
Dg/EMNIgK5f/FO7p7AQLkHSy/w2GtgrMhISma6BgsmWIddBu0cS+pUmVNNNJGJwI
Uk3E3cxuEh8zn86b7799kRyfGevkCli4GsgSIYbwJGifnFvmojSke+lV66U/eh++
yQSBZNH//1F6zgwyzm/V6ys6BMmj9zva93+0wN7Hb7Yqx5UmZ8wsUtktZ3L2zA+6
QEdA+hL/pPwjkMPNlGlIEGtxiDMVeFmgSEAXAi64WlxPsKBx6yVMKqgpjC1bJgnn
/0i/LNhg4hVfZInYrW+4dkDMTv9zgRXPJWF8SpAb/Z5wsEkXME/wmHV6FbB92pX5
5WPWC8+Uyypk7AgIQL++ySArY+81voRSOuPBvJV6JqAo/SyVL6Gsoek0IgsKCmOg
r92lRAsXQ1Wxyfozi0nLY9pWhQK7PddT3SOB5wF+0uPZaZDjDgsPlCHh/8UllJyS
+wfZvs9CoKFPtcp1gHmhJ6q0xbLJWPhiaUY/LXa4ALAKuRRTgE4+4XOe1tTgtwdR
zreaIeRuwSJcmrW2XGmaeYcU21OenD2QDqbmb/IyOrFTll4OztwyOzu0PNURKPIo
NkU14F77CCY/7IDbJ8l5SISlz6+Hm1JJERRr5rStWyAmZrdQWxR/JDcOcXB2WRWE
ZFOui4thoXXHBhlI464DF72VDYZAM6HAW04uMN+qHBWlTeHKIeMiS906RT2CYi9G
n1GyuIcU7KMj8//fzQXMBOkIcaW7szMzot4B+a9zyQhZUUM0EnH+cB67pUZD6xcC
VNmU++8Z7Bwxj4KZ9ionOS2OPxGY+7tkuypbXqbDJfaPyZGEl4IG0THq47Uz1qO3
lnnbNe7x3QXd15MB84pAhb2fHPT3TbQoT8Bubir9LsFuBtF9+QuC1JfDmHt6LpA6
iDPGPhTKPA7gdOipzLwGVQXdOxJIhxXlSc5TY+FTKo1ePNRRUsbN4Q2z5xJL0cve
S7ygT7VSZS5Pf8qQy7DVl1/eXWu2NMOZdNLHySAomIi9l+cp6daVP0XevwPCEsCO
WVrGdNH4jJzLxMGz7srxtr6PH71UjJuAwkVyg7fH/+qWMpt+NAg6mgpTmLhGq3fI
3jtCMRu2S1uDgwDMdGkTHIEe3/nX3NhD9xJjH/c04Yyagb9IwrDoAxp7hiS5/zgi
t0AmWJ+53S/qL1LwbIdUmOIm6oK1w0a3mJoH70pAFhiiJIW9ED7HcxtKLydkn3Cy
WwhuO/BUn5wnSRSWtyaFIxXULZXC4UiiZGD8iHWvfSPqeSXaD7KrHK/Mi31DWMdY
m559PmuYrSDiTxBx1mmVtC96LKKy/tiuNemmpUWre6PRKBWqboxOQ4v/qFwODyq+
lHJEE0N2Pch6p/hWjeguRUlRcqEhePHaklwG75Xr+iQeyB1DECQzALVsx6bYS0S/
x6rXJHgump18Fx9PpjeAbOgLm0sJ2PoMswmvLhJoo2KqelJwf2rfjk27It7diHyi
LAqCYTR4z9+OIs02Md+5U2fKeKPgxp32a9Qo55WirdxeCrpP6VSm2QzIpWy/gNpt
+i95vOLtExgA3eZASSITaPCs0qYE6id5AAtn3guVJoL9bLNhQAIQnyvgpDVRlOBv
uHNcQ3MazkCNjXPeZHqAj5+SCvaWKGY7CMyG7WjBoX4IyWzSYcy7JawIdSBF6Y/P
J0sYJ0yfqcqbarNZ8i5jPpoUxTP8GQRsqJwg/ZG19jjXmD0sdIUFcDqSB4rJlbS0
EDcMi5Sw2JBPAYljRmgA/2k10FFXavBMMe2z0LjVfw+mNfrEP4jxH9PEgeouNOkX
Ziq9NfnWGY2DWE+hvkROrm5u74ZAu5ImQqDfOj3FaGpAEj+2nkvgl818X/yb/qD2
d6vrAlXiGANP8onOKvLIBPXASQH9eesUX8S4kL/Z6MHpnsz6APNqglI5hvdv5I0g
ugIoJM45yGv+pVXRBSa+9umyZcDjOtiOy9pb3fZh4Y+qzHpFkS8cInxoeF0IXwUu
XwQSOp5zzX5CSGjxF4tsn1+CVm3SrDOTKgBUAHWrIBbeIrLayiB0cejkodiP/zGS
PV4lc91DgsIO9Qx4XzMzNAq7LkjOUW9Q1erb8DbMYtnaCHCX4n4uldPs+N/hpAw4
N34H4jyWskHgGRxwC3ZcBdWPlYlr6u76UyGR3tlSGFflqiA743AFc3nMmWy8i4Qv
M7S/p06h9PX5i7phaBtEQ/w44efJpy/7yqMNrsDPVL7QMHnBJCTOknzusal8efXE
QUSq+zpZ1w1ZM9ID3NO6N7ITbIt5yphr/GBX4aREgwipDaXnq8CoY+OTAgrkoLPF
5yBVCBwomMpuQJH7GQrAD7IjiB5Tr8A8KSfC/VHLOacqDy7uB0ixUJVFN7tFQG1t
vMtYSCowr+MgYl0+84qbQFKc4eQ8a+qZLtddlWcXfxe65jFwmNracPt8+4xpxMgh
WLgA5kmbGizbuGVU5BcjKwhmhI0W8pZZK0u3QERLnMPKBlwby8u3ATgwo+rXG3RE
nRq0Tq1AkCGIcfJCSpNIdUeTXYbyprt+1ejnq42TgCQ30y3QVJNaSIbec4Zb0Iox
fAvmivGQ5JO6v2qu/shibg117X8MUwdo/DYvXci1bCRpyBJ3FouB5bbHyaJOcXqT
6IkyYSjZSkdobQnoGvB9SsT7TX3hSDJlrM5QJa97ZgR6Wqu6WQjP+GVmSzQ9IMB0
pfzuU4I3oiog/wXGaDgQ5I0mWLRCPsxhkLAr6l0cygVvPBDc8K2miDdKagQPAy5F
L99LhUMvzV/j5uK/phnUIAjRKGYfU/2+ZfDn6frROz6DC1Y5DDKhMJi/JbHTeo2K
WS74AnS087Y8hsBcd0HU5yCvTUixwRpyOpJfR6/hrqzwdow6Q7gWnHKBkOQ/Nsle
Y2uOXRvJLbb9tm27tHMV8tdWepcZh0AVtd5vyufOMTmIydi0PpLNm4YCtiV8Wxjd
zkrp2kFvmrHXJ9mTH4wDOp2X/MFvaMHE38M4beSMKGgUbw4Cxa8a9YegsZ9a0XT1
CBpmgH8IWELnwTZLCgklwDyx/K5sx85ulyNJ93g1TnJg5gC6kMr2o+QTXSGjIL27
0uN/61l/3Y1oy+qgiqJa34yndG5UBLzhtNt9mLyssmNrAqthQXjQC5NUynIC4Sa0
dyB4bZraKEQJIb62N5d+44kGCyezLNnwDH6is58g/M3UG9tEPumgTPO3bndSciZh
yZtPQUGpMXcf41J+sMXwsGrxUPyzcwZKqPsOESirjj0Fh/lXwTMCYCs4lXt18rUO
64iucShyv/s7t77OsIebCg/0PX25G5vnTpXyLNsPGZpxczqK1yS81c2HSweGFhDN
z24pS1nvCVgdSvNrwQpzMvUd5rfmD2f6EjDtN75NBO4BLJFVswUYjaV1dSU+V8Bo
yxZ62DzXvbtM7x4B9BLKwM0OUnLkkuMfqQXOjxgSSBzpDg2Bb0qw5+TNDnVXCuzW
AM7WlBVB65IIZfOFGRaDZ9ruO6T5LvS2E8qp6GHCD9EkRygsupicPF1GtP/D5sRN
4UYAgdIb2bnoWxLSz6C15hSdGOMES7aN5iPaQThGD4rpYHdhdUglkv2ZVeMBFnkc
vb5ydLUqT9Tj+TZYhlcgeWykuhXxvcX15xZ6JGR8Q6xmVZ1jHECBz8YBBmKjqubs
OCzI97/KqlyrUf8VB7oSlPW/2L2UpBnQQUq3Ki6UftO6bzQkdJspvJePBqEBu/kV
I5ydRsBtrOAA5F1h3h8PW9XfXyzH/WZxtxdz9D/vgvBT7t3EB1ZW1bv46Z7c/8E9
eLGXDcX4jN1gDhBGwFFlv4j0AdoilFEcdQBF+4wMg5+u4aqc6XoAlU5lD2HvTlQQ
lO2zGz8vJACWW+RI6fMRtNNORCkNN7nes3xf5XUJHPLlVkgw9/xHab7Xw0f/NvIl
d91+9HH599P/74kW6AjiPzvWeP1xjlwnlQT8LKHgWbvutD7WZId79NQr/wY/1xci
hJ7ZuSc1d9rBhefE1g5R8apGFQGtisB89CBH5FCjq0Q95Sg7GTF+se/h1DigvTgs
OBuOAP6zRPP74itnxHvqvOm5NbJtdpc0VCMVsHZ8spXGv1AwwrFBlx1aE3Coe+qJ
+t8u1Rd+Bl/iwF46kzuNwRreZELTqY+BsiP3NrW89B3lzoJnJ//aX9ThSXKLMAbm
Dnk/TQaBc1y/9oVDYWHZn3lVx6OL12D7ZGyvw7sJ6Ivpf2db+VxIjVsl9NR7KzgV
+IfzD878/Y7BtOlJFc0O3NaNvI6wxeFvTy/Z/3WQLuspUSVU+fsZR8ylJP0JXBUT
CEy+eXYLzZ3lvOSZV1LvCXZTuZSveR1Pgq/GPzUMjnWjbl8tuZFzkIn6CVj0PCd4
Ior4SZlZ/KA71GBGXqvOmC0Ml+ZeeO1mNVh4Hw7obNDxqNZBrhqRV4fnk4jv1BXM
gjCwJ+wkLeNAG8qPzKO6JB4ygLuxEP8J7EDiVESMess=
`protect END_PROTECTED
