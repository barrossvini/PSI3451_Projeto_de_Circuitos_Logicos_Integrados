`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p6Ut36q7+VCIlV48bE2iY1r5YR25ghrwha7WbSDdgDtJPwvhxvoVefg0TL5C1CYs
gEY5En8KWopdZPwzO9+/rG07aIqWnN5jX6erwJ3BaPVqjnCiczeXRR4mLeqbcuY5
8gHf2bhCe/oHRZOY0ZAhy44rrcBsSGtm3na7dhq7B4eLuLXEAXa6F3DCxdArw2uB
uwC+vR5+GX0o1RRjiKUMnvCpehEXqmKHjeFYKQHoVLLhvc3Iy+plH1Tn5FHzRo/j
W2rC5hx4hDJE0/nzQ1jYKWV1xJ9NBI85CtPq+yfnzqfYlSZrGv6Rm2h4lxcqxzHX
B9GrO8EGjvAAk2ifWcO9ufQCJuXdfRX56FDcZP8eo7FLhd7+2Vl8smqt6BVzo9q1
UDauG1bl+6/9zPgA9GOMrHo1TNcqN1w661qGAPOhzj7vLNBIvKVmT/2gGSWV8kJQ
lLwUUkqdUBCM4V7BXrDCRdoxWkgrYuTPkvHkoXE6m3U=
`protect END_PROTECTED
