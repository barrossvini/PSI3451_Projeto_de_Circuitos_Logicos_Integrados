`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1hlPAZFm1mf2M5g9bOoaawLtnXThhNs0vxAi9NIyeWpQxqoPv1v3GpVLmMZAZNiZ
fHn9xR4nfPBkmxBZCF1h/YGZSJtB75swUhOgEBFP2Gsrj+lM6AdjJG9TPxcdsC0L
UibEdMJbvA4ej8VnNaa6+BNM9xULEnI5CPp2uZwajlOBxe+6ueKiPx1dbf8EEcU8
asodSFOkvubzsDPMFjiaBxSrnPsyJW8gzAyuSvWXYkAyPPbHYT2Qy2g7HuGVFQbL
Tyryf1xmeXsdh8rszvwzq3L9UP7ckt700DSTTPnfHaGEEIRfiorMYggW8PM+SAF0
cuetsSSTR9GTb2a2rY4CJzCoem3zEh/H4fG5Mcu9zezOi4vJ3quXWhUprCZeC7/2
yspAxl4CMPgz1bRCkWedSDlIRbrMWx9s4vyiSGzgc0+CFmJ+BUPDnq1XvgNCaIz3
5mluSz4Y45/DPx0jggjgmcjphBVaVqcqJhPMHuSQhz6VzZa7LRkJtSHowU+6oSGV
IhC7qDk7Y6wwq+GGFZW7FRK2EXKSjVzD+yZjn9+DfXEfF7IT2ekdnjkVfYr9oS8V
+94sVgwlhZHS9PcriEzTTUI47ikHT7tniZXNWKcK5NmuJE+ZNIHz62VDDBy1QVUb
76SHxzch0I8MxLwbcCQC6x6fcXUlLgwZjYvsbv/aXx93wjTy0Y4RevIFJVmC87fv
kRisPlxla1BswNqTZjiULwNzNXkS1a/r1rgQaHFBRQqAZmi3FDAZWE2isZ4ccTCt
ZECcS38307vmjaQcXJ9JqT4NOw/ZM7LccWWicBb0AaBPvIoDOwgZgDpgZPBKJS30
m31bcTI0Vt0VYXYVkK8HoR5oNA2Be3Ya/29lbQRw5lVFsXi/3PS7N8srWByZ1ylo
zEJVzEhbzEQauYpuS/q6X7pO4UuOt7dcReUXVzjp81YiWGGq6HffZ+ZG9DO9zRCZ
`protect END_PROTECTED
