`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+pW531g+YshbJG7bZSHYl4Adp2P0KszpZA5mp0VJjD3P4PDkQ6CiLjozcOpAW4S
RvGXKfD9VUu1vc8fgVQ1X/7aMTkCzrXFl8gWQ0wGcxItFErdTE9Fg7d3vvdGz0lp
IoJr6rxwr7qC/nxNHTu/La4PUd1S1gWRhr9fAA6ZYC3yBkQ/u8zZOH2clmReuANl
dTx8bhg0EiTtCxm+3iZVQXt9V6lpfhR/cOptcbMbhKkUwG3xjrBqPRJzyLaa/S1j
T64CNupB+TUJs9f4BRtcdFldA+GPWx1T1N+o6T372fZy0yQxUVZtmV7EyH8h2pXX
WSn5OwZn9zTQ3ZdkQeLIArB8J9w3eg3dCoDbi4KDpJjiv4LucDJPybk9w6PzQs2/
xjOJXQQeJplSQROyrMVRBbARifPOifC2JxtLnM5RCCZYceQM0qdnMyblsKKukTFk
+kZXkgnJGbRgMtc5PZHBg95XVw9mUAf2C/twnhMjlCJitmP5MibmuSOXD+rSWWSB
94cwrP0PdXvRGL+qiOBROTBtjBQBYhxw1EbrFMZX3jPu2V3NRUn17krYF7em69zD
2Vw7vZPDODYNkV9npR19oqJtu9Qkeh4Q+KUyzuUkNC+jrA1aYHRLT0rvtl9G/+H0
WKnG+8zDzJdmBQOoJ3XlhR0bX09tIdt8749eBKjM0NNi+oENxQrLjlixoCxFBAib
6gJFl7fGJd/VwMwbAqfFkZUewq72+SszLq5UyUk6UD30LYqQmkQZV/TVnJKYAFHr
QhJut6+rGWfEAT8j2+1AYBPV1Ecrs6FdFtR4VN6S+baLi8vttc7BhInK6JCMsTGF
bnvXiTQRswpTtMAbatMnQn+Clrs9iflcoqlOQRKyCY1xeeroovHYINNHN9lh1w/6
y/Q27uXz8W5bGRjJTBsO8jGij5kwpAptLGotIVGLQe/JTtnjg+T8attVoi9qAXwm
HZ7pUMbsTfqO8L05NOn5NF0TUmOVxjlKlenGX4N+waJ/fLAujkp77619wllMuZxr
q8kOT+Or7WXigdICvQoG+2lrlm+KkKayNheo2R57gVDeaJ3ElmhQ2apfTWd+Gmdy
tnxDh6QKv/SOnVVDMwb4ukeLDq6EAFPyx209Ul1YYTJ5i8nNa5yS7M6LOQvcl+H9
7kFSnJZUhAcgOMUCcKHDs5ZJLnN+g/rhbaysvOm8R6hnPLNzLtoPd/A5o6K3f6g/
1Mq7uJ/kGh3N0pL+KaMFcqc7JyjA7xwQUAdWpXnVfh8x6mz7itKENnwNamggMc4f
josn+i501V7duYHfKElt3rOx3LvksyAJ67T6RI0rL5mIkSdmP1t4Q3wNDfgx42Vy
/IaH0qEFr/vsKQfk8iFSi2DdnvSFW47V8iD1kdubQhsHBNKpliDCujHyWKvvQdNH
/UmB/kYcETx7WWdHwVhS3XdB5Uxfh1hC4CXihvYUZhM=
`protect END_PROTECTED
