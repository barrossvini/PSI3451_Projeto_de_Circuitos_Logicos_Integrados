`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4sinFuEBMQaicbohMYxO8o9iwASkHdNdFkUtE61LvdJw30J7r/XutXNokYalwgbE
l+7kcMOv7WhxnGL1S8hd80Lf+JXFwQhXl5UBeiV71olzeCwmzGZlDQpQLMUjzgAC
cCFfIkzxI0o8GIDmh/gO+uNPzTwn91FRd5/Db50J/Uwj5vUk7ZSNCGDEUWozYHyD
k+lAQlTYicaHGQtrK1mOtthywelFHucAORNQxPnLUKKvudtaiufLihzH4csbhlSo
pHLzwFCPl+wtyY8bxsT+5b0DSQsqvzyEQ63ZEXlC7xiDZw+71ZYI7QM6QSsLGXr4
4svphaupaM63f72vA6loNSYWLOO46HtA2kNd5hWOnD113TNfNqKZzT4z7ModHIo7
ZfZ/LXOSHxN+9E8oozLiulR5jUfkxbO2tFZFyo+TwDwxi2Yfd373FmlRoz/KQddG
SWAoa3qlzQCynRY8qtG70vesF2Otszu78ztBMR1uk0DjV3dux+2GpTTPDB//lNwd
tK0ZMxQgNzpfsRwjMLsTNLMN4UEVCgAMrYApZ4gFZjphvZo/hjWv+XqA0/Wk+l2U
td4nwtzEPQ0kOhcHW1xPZvL22w0pyd+Vc3AiQlzfxWq5/3G1EoEcJw6hXObNk4us
Zif4C2QJ98tESPbcuVojwr9JDFnTouly4v6fIUXzt2m7xCM8zVkloZSupvqgmxXG
PHSuBWRlptWMF4lrI9GQ8NStk/BA91mKkpKDx/RF8HH0bppCQMOXEQGGPerHuEVW
yfBvpG+TJvko7pRgRSi5VVrlXyiVadKqGFRRu7Kx9u1KLeFpuYV/+Mv0EiZHpBbS
wcedEhPKfhovXoM8C7rXbJnUs+Mn2gD2WvcB18UIc72qjifs/BHEtlOTI70byxKO
tgnSrrf01oVPe7rPhBGx17FcjmBPvrXMec1uIphTEDhBA2w3UURo0HMyQIxTCVfz
XsRnJ3NG4wq8EC35oVV7Q9GEtv8IBZ0e0v1VN8S+VUPC7oezYY5n8NjD3x+8Hski
UsM8d8Pqf3uwtg0oAuuinQAWv2emvegZwdMf2dPiiSol7/lI47Nu2/a7Pqi0e8hY
cw3mZb1Ca02gCUHbabcetja86octiabHP/P73X0l37xS9g+AZH7sbn/xFLqynwE3
sk/5iMBy/xhvTe9wfoL85PWZtorynUkMxEzPyOnVx7EWUvpwonNsuEXZz4dUtAxY
MEA1FZ7ZlKh5x83qDXCsvz868wm0zs6F/5feTpgdNS9x3bMOe0YuOR5VchR4C+E2
zg7gEBdb+pUG6ekuYixi4K4aQzolbNXH0BLxp0hLSHgnSaGhnTra4jo2d/rxIvgG
khxwNWoGeCJsc5xvotdZzDUDPfrit93Ny/uprXLhMWyBQucL00vbDddLAvsIx69q
wrwrBEwo1RCX8qeaeI95J6QzSeTxolm96OXNf+TFfbTniMD5HSY9UomeEZ44DzFV
984yjSuFRncBxv2v06nyRKYl0l6kG+ECYoB/+rSwzeGZO8LRFf/8ITR/aaerHIEs
m7ns+TPXmk4H+VvFDrACTurtH+Ncf+gL1mP3VQTH2Kl57sf5wHjLYWlJDxR0rqWG
4swu290HJYyMt28/HxExpxxdFOVLCy8VS/Qq32ulr/lz1UObtbR4K7q0+EBiSeEa
kqEo0dTIp7APrDLD4QuVa8f5cfNhzIm0hRy/1HTXIw/fFZmaKtgX8MueMcHWMvk/
+iJt9bcm0TS9KCHTMDQ8tlh5BpcNyhbb4VgFp9skLLBm8rmUNnbViOjkr21Q8tWN
qqn/bFfzVAOZDo9y19sLCZ9ynOSBxcdO2BG0DltVWEdaYFTXLdilz85p30fLTrPI
tnDPxj6QA4dzW+QJqWDgRcwrHE5rovj4RMwf6R97+IKmIvhkzq0pvHbsb+EfCD/r
2c2zN+L/CDn2CIZHnBKl+BHYg4LMdrhg0yOPLXBFWI0eLUlQJZO0hZByQksG9wTz
cPI3LXpcqKWrAXv4gbNOc2UJItNj+/5vLtC16/Cz+T86SB4zE7aXNX8x8Rf3F4u5
lj6+iMX8zO/wZokjnCwi21ZHgLG4kMZzfMV6WUWo+YQ6Zhbua+tN6qMmGn+5phgW
J+1s2rSbTnZZSzqt5sA8NhmVPM4O2QbNgS5PqCqApqSRvWpjmpe7xAECbn9kD9N+
lh+//MhClP3+WtsLwZcrem5igtJixVSm4Ox1oFsJzzXR6P45KREWz7oE0S8rhfqs
YspUbr150z4WU167Qz/TboujrYSz7T4bAPb0vjm6QklmwU/C5tQgiNvzHYkWBPjt
j7PSOLWEwpOO8E4epiK0YPsAi6N/6HHQe8MnuwQKY8FSYcwHXVVsOPI1k5zZpnDz
5/sklaU61kONPnSQVxazsjEOWU3x5fO2Edw5Zhr4Z7qS8wz4aKtkWArb0Ax/qhRW
cx/OB60a+jG7VSlVoI/NZx7y5dn3zXgtDfmztZM2b/ZET9KKYyFUwOAr5t7LOCDu
dJmRre1VKaKZSWx0+6yXzKSBEtZ2eBDgAKoHpuPYDBvaRZ4Ga4g85U0UTgXF8ZWD
GppXqy8v5oyMPHWznyg7gvYcY8YMUrxRHkJLOMbWUGYs0UFE5j5ypPkJaXj8HYev
IFb4ArpRMqhjVImQKvPj0+cGcM6vOUqykvYt184tUxZ0O8khRUU9P/ohqfJACZlK
T+9bk3WnkAbYHeTs33s01cjQipZqp+8Op91U12CeFiDygNpc8kJJQMhnr3tP7i8v
YlGsstJ23L/LeQTosd+jswIFgC+WsB+iM/5Ds5nkU6uGCy4OO9qg3uWkC89lSqZA
+Ag88/b0ABWNgprhUeRpnbKWtVIVfg5S8uKpAh/wOxEe6Fug4Qg7cgZiWYca1+MQ
SSa8f2dq+zILjBRTbJqaNYw/QBZ24Z4f2QW9yaiSzBXGxqSQmzBu4/62VNw0dYI7
dRBoP5llnxvQ2NHjttCoCf7ia8P8FS9q63CBO0HoL3DBohElMGYKH3ScuHEJ2eGw
Ih2WESCugTh7tVPSAQlm0/sSQzvUghCAOlS49UENE4stfVIoQUVC3vwyVVuEGxyd
9jDigoTTDuZHg3ylUWrNiuQuhwSptcmE6vhsToDy+BXh00DDNF+ZycbHsScex6x5
jLUzTpBkyeuv4H6YcwQLV8PlDOAspY3ebV0kr2nfNMu9zXrfu/Dl3EiB58QNYjqk
Ad54qeQR51ij3fv8PB+mDa8HWTuFXi6OeKvVdJqyrXuTwLqo2BfG0p8AFEoeIs++
CxTEoQfPx85YDbCkaxJWHnxeXdlmUVjNArGHn4qC4W35SPh3vENQsFPNOg87vxta
X8/komhUZTqdjN4xoWHQBTvUmQQX4uUDawG0csgPocF76h7qxFlw544IUYDC5Qh+
DrFxV5XIPOCkWjo9AGry5bLwbmN+aL8JNMo3d4ez2QffZq7Wsrlu1P8lHYV2W8FQ
g9/ONKvVGk+dtuh/CbSuMEwv6ATr8+8oJNAVDxcnEghEcMXs430hQDayLKkGc6vj
wGlIfx0Z0Sz8N6fsWI0KrzuNF1RtaiPIaoHgUn4WXI9svPlU/kHT22X8Fu/6hbRm
vs9Upz/VAqh2R6mYpLLDP6AszuLRmQGy3jvGivGhQevq1R0ujWx0qcRrs93NqYz9
eY2GYzj5G0NiaBPSu6ZjL3myE70q5cWUF/AoMTqTHtaKCWoKNlB/PjUe+yJ9mXPw
ShMT7LFzTsTF5oYkk/duXFLTP9qb4brpU3lkfvJeyySv8/Z4FNQsVxAAsNQ/hU32
PY2KERpwiSVoPXG4zlqLu1YOIlMNTMKfH/IOZxjJ7ytdEG3HCA331CaD1hDS4Ecu
peS/5QDUlBSfOxTxBkMK1J1RRca1tELUDAxkWbMy3G9wBeeZmAwv25R1DXO+rkOh
t31ZjgfNEz+yvaOmEak1FDZSluiA0AKeXRT9MgwnLcKmf4ItQXg3yvItQdx23cxH
haMa4jOBvgLb6hL73qzB5hYuJyfklFdkM1xLBTvyxYZ+4fL6rYWii14NOhRWP7Ic
GjbrmBw03uPDkCiIzyRyEsHoabLCq4cvu0dBkRer9cqw009PIkmG/xGX4s93rVz5
yxSmEQVRPAk2ZMdQZJtkagKbMNgKyI8h0du3aRqc1CHSzyGaWJHF2eoiB7XVXksG
Xczr2cVgZTqU/34I4+UNZYGqXY1X3z1mJ/sNteHrhgHAD8fBT216szY70CWIfRRv
nTjPqbrW1Z5Ve1/gWyR40uKQK4t9gwBkr0nuWkTt5t9Hdl8QHHhONYHQJ7fDavAV
seqM5hBzxjSnFwaz0BOapXcF7h1h/70xHSnFkiZVbs5ycSo89uM7jHBzegU33U3u
lWhfaU+ZfnzD2oGvBdRCVTl8GkUjn7tegU3VDEvpX5R/IQk5v7443l5P2MRiuvxh
vxlsemjkPA5AUgTUvdM+I9477WtrtZRUw98RmK57x7jhF2fqyEFbdcL1qZXhP979
meIFj1CVD5YQXVviDAiuOpmxL0jz5ck2T4msC/C+GPZRvEOC4z591JDI5KhII7Vy
jhNjpnUgF8sSsESczXv5NqxVF0DnHjon+0zBo3WqlXRmvPZmoeIM5SsufHM3gt4v
`protect END_PROTECTED
