`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ltbyVun1/suSkWQP0ySlk/mf7oRSiUPUCMSqnYAjb7kO1YAmU5Ms20jL9680k0l+
/9VC71PbMJbqNWbXVvMG3JGDf4SpkzHFrFOiB8+Jd/IF158bjAG346UV5ERPX9ap
QaU865jcQ0w2eXiQjZRdtQ0qMqmCwyRilyjd4oU3+IzIUwMDfji6tdcejuG9CDcF
h8vL7oOepzMOvTf96pDjwQH0U1J3sGJL5nLmSvPoaIjdQRMet20lpGNHfTO+s2e1
YNuexxjtdMEedpmyCuRZiIE04M9hPpTsN//yBnxYfwzhidErG0igBmjbY2XOY1AD
c+Ie+rMHTzuNJECdqmRexH+7b7mtVNyeNu20Mlwc+R2HnyYnXknzMro87ixuppht
rlrW6zJLs69Ww5EVPMdyUiqAde7E447bv3Zh9QqhQUhfJHngFG/Dex+ggbpsjuH9
OxSp+p3ear3f5kR7FFKT/ZrBQSsfnMmLsvqFtZUyRUrJMBzg2fHqcl42xnWsSLw+
KfA7OXqmy0nuLqagvbbC1ZH0UgFeRHSJ5VY7PWi5moE43otQwb3c8nkCFlMGbEgy
PCr2oVzLYxgXRvsz9E38EnEvm0ODMD0NviOMRFAj/N8GMR6BOteIEfrFygMzu5U9
pKmxCtBPjVtKtwPoNtMKIWihwRFA2UVL5JdVKd5nbrAXPx+qYlIg6oaQPcT3jhD+
X/Ra0YTqcIkSwKHcQ4tXkyz53wSgtRb7PwJK7v3MayhVAZlIvSCB9ZnaLmDobTN3
g5csLyu8tU/c25i1upkQ7i87l9aBetLmb5hzDGoLDqy/i5brrhZFHBekb+3jiWyj
rwu5f4vIYNelJ4v9GfdZ4culdZw7+ZfOTi93boBxDUB/c/PFHQicI41xWzq7RxIq
Nx74Z60puNMQnLa67vpytSqMcBlFzwMA3WRFdrXz/B21Amkp6ivwADXlwNayY7zJ
YA+dRUviMyZkslu36zweWEBm4Tr+uq9eROgLfhTf0PxsttWouIiY6JULzogw4wZU
JLRTkBtlXgtVt4bnLwLhuaSq8ho+Bejel3Y16LNlfnmrjdHBG82+ZhY7PArLKjFW
TV3sTNGfQ26rn9akMW80mzQga5XW1C45Iu+sao4PM7g+fL1bKsY15BVWEt9FBflF
5BNx/4QEQZLJneozdbF3q+ju+GngcchDoLtdCu9M734WwBuE/M9Prkh2To9Lzu42
zVLCOcEEaqjktkGFz+tMCFX4F9XQlHOJyyKV0eb44ytFbA/h3jFeJLvdcjQlv3ou
J1Ch9fxAZjM6om22Kd+4s38KyDv1J78KSFWpPAmBsxLFT70yShg541CpghqCd/6g
FD/XerSa5tma8sqpdDnPR48AXic1JY/f+IUuUNSir0Wqb9dH8TJkJQVFVLr5nn3A
o9wQ7qGiOK9aKaeyinvrxYNwwtnKnoRAWa/WQlILnxUHOaz8yjMaSY7Km0/Q/LS+
zZ5UmAsoWGKIWAgcT/pcU5Tw4IUj9NkTNSNuQ28VxxlhBcqwT/tMo21GxSxtDzOm
QfUXIfrEfn2/JKV3arxURdqSslGWyDuAwGKSdhtroBo95N1XzLuw0LsB0Onoq/5J
dKXvY9muDURyeyk8zD2nle/0WX9o45RZXnTozS3c8QV4KRQlkUqGQ8q4lojV8wl1
La1xs8Ek32Gmhgk77evMM9dyTy+pW+XA5PckekHOi4ywopHPyOVsNwQNK1tYdMtC
EWye789atKzbCQAxKWHoSJ27P3fH5IizZjviZ2etw986fqMGo3CSE4UdqvVYBYMp
IGF8TiGlRR8S8CNgeh45UaBtWzSyygjSm/9E00EZ6ser/LR2TZAfR9CCAkoI+uaL
Rww6cDTwVlSj8eCfUDorn/XB3mDQGGqVGCxh/BjUZaFBgkIfHeL3lrPnb4NVzRS5
ZqUyo3t+Th7cYt49BtnocPo904wQwWKVqAI+/+E2FA/ebPkjgaJ9iuW9QK0P9aIT
cd4nIF6qy31E0+UipxLsumgZzNlGgPjcOWHt6uHvvyIeZkOd7BLc9L7zQWf2r8LD
quoVwSJCJtQr3kOg9xaS6LgMpwiPaNemOBgsuPuorZ571uzbnv4HnnSfMngf4HW5
IcznqQhx2WEjE+Ur9G4BLSPx2i1BxIFjnudsaKTTV0mVXxC5+4vUgzs7QaE0su29
0JAPZbUeVrkGWsMk7CNlipsiDB5535DZUTPmgzdFs6+Up/0f5mIoUpzVDxdPHj4g
dNSAK1+N/RWERg/XsojbfDjOpuzkffmyQXEkkhj2Ayh16JrLRxdZy+UAjeGEpjRv
UW63BkD8y/OgQgkyg/GvMGVv64PA7WdWtyyQY+TGivANd+Ti0+b+4rSaP8lA+FAr
zvQNHCE49VPrC4zxSyyWqAhEjwOW+OSLUWEzaphGmBBvzmlff1oWKh1OhBzOiQlv
onX6fSmSwanb3IBpu4QfMKsX740tW1zlw16lKhu/uLvBHcwEZXl6cgJnpSMHBbSh
L1VhXNnkSD7Y9iCxYHU5DNfM/mwbzRCEWKie//HHauVwpeD5Rsik6993nm41K6Bn
r5zCicjVT1BZ2mnHXg7JOIAPw4ECHm2uwt3UtQEtshkF5MNNBdxv5lHyvCdAe81u
A+AJvoTi2hdDr5FP7agWIYA1XdfPXe2N8AclldzBD1AZfE13ej7yVQFa2DiaCztu
czqMqAxIMNItZQYQqRIY67CLOi1EXEG1VQo72bRmrvtXkZwFmXcH5jYTZ/xrgPlo
wwua8CyevSNjpm3+7tMW1cOsbYHzXk+5aiXTn7Ixi5sm8vGqN1vSPBuksoCtT9w1
cfGAFD16C6hT+VIp27ksM2iYYX7d7cFawz854jqdp3HLdQmkkvgjMzsIi+b5WsrP
0TcnSezk10wmTO0cO0qWfTn0LY+NKTF3dszhLSKMJMPdlh2zy4mmmgdxobb/T/ID
xRqR+vdQ1hzJXeS5C8N2LyLOGTVE7lZ9W3ESw0+d1F0SEEMfCt7KMlGFkCAbLBAu
6HpcXFIG5CE8JU421aAh6UrdmFbd/93s4hi1tpt1EgN3zw7zSPF1GQlgfcZw7X5v
9N2sLzRGUvK+9hWbQ9lkhD+BcZzCHLmPxfqwgJuwMTeLmSSuLePoNqxUcpWPy5Op
VDZlk1K49lx2OmtS6OmOUo38bU5QGL+zWWZ0W1IT8taL1vUVC130mlS0XgOKG00u
QDmtnYEEY24Ui/W8obaCWs4wsKe6K5XBc9dLD09UD6Vi5YTGJv7FP46a8EBV8gWA
avO6iqLiZgw5fNRG9Pyecxy996Lnlhq/efyxs9SrLe1Hn8OaObeCOkFaq3UE4Xjm
MWIp0LerxPJWhAkcdC0oZPbSwotF/cqzozbYin8VFFL0K/gdKIImM79O1njwtWez
faRmPd2sC6LoQykh38zMMmjEGrb3l02Ziir0r6ddYd/gJI2LGRMimNwhjAOOFNZX
//lrB3PL9NIARCPVietXoYswYDIc0Zw7E+NQtuOQvEC8fjJJd/Ld7GhkV5bL2C+H
pcYwdXEi1f++KLcmxV8bXV9WSkXFPvd3iDo9GGyCt5ceMw8x6EW8bgROIDBF4vPM
PX3C5UpcZjcJAaQJSCJlIM5ZZEE1hD6/P86XKzb0V7LuZk0rjd+SBh6S91vydl4f
EXmaLCh+OmHmOpVGGJ2FxEyEWeY7OtqJ4l2r0s70ssPBW9Kmk7/g8/h2fMJrnr6K
3STrooAKB1RJFus+BBIwdcRvGcpAJEAgC19A3mmHY6gSOzBrkHyqlkCOX90odj5k
O/csjGU+vq1ZsNCUeov2uuFisXkkHcwlPdOSqT5tMKlgHHhGDMTImYwGLQPL/Xtu
at2AjsRkOl3YcmC5wmwEYP5+UdtLorqAoQz6O84PYPOON8x164ivXjyBjVwGlf0B
Go2TSy1nitbqblccLVgGz7owJtOcwj+iMvul8fEfgru8K9YCNdwX6sI3gPtDGKGK
lAodqEXc4vm0h/+js09hkqwLm2h6U57NoVJbMLNGFANWQoaJFCPltIAOExAH0Jal
osFfrBGg14RWDtP8zPWQlc4fJZHnrEJBqjZxyzXxzNa2jR4UIXXA0a5H9ZQAGZUw
kY+mm3ccVI9HKy/hrlToxlW1d98NCYktlo81du+2ZCruXHEtMyAnywKMt1ky8T85
/HHs6LOc8jqWE+cDcyGC/yt7SJgF96uPI/pzc9oUXZ5pI9WZ2n9WjUJXQoAZPCs4
ARLSjg/TUwn4B0LE9JXGrGmuPUcrZYWjxdhGO2xFxiOE7QxrSR67MVxkpQYbzPG7
7gwtBuDiiGJJ84Jl2NKpeVHGSJuDuJpok5GpbNvusy/qm3WXwMvKNuExJ0iPN8PP
7oArYQaRF3wZtL57KNzml0+KSipX2PzPUyFw8jIfNe7yeLXo5n1JczfDJ+GAxwYg
PxUx3ybJ8/TSj+U6iYjb0uthVkShaI7NTDVb115KeMsYwZiDHTxjNqABxIo49gtx
p75J17G2ppEq9UCZYTSUDawtr2U4kqffa2WQzMXHosfvmQQ3DvNhPFrXA9nP3JGL
3N1cBan5/yedcA3Bhl3qIudWMPNxcyWBFtZIPJHvfGBhoZU//9LUNQlNi5SAG0cX
TtCFmS0WsNsCrYkhCq5o3sPmRHniP6/1Xy1efVxeavTkBwlC+XL0IaWMbM3nI/0T
8gxmkxhNNtCJMAeUWl7YFcj7hYBUXyJct9eN41bVkbxE5uNsNzWDs4G2fuwLHjzt
MyPw4CrBi6VlF93SK8i8WFwo7IXPOuGMAOR3u+XLoSCrPRtc3BMSSQuGPLsXn2GG
7Wf/0I9BD9L0Ydhp05BoDfx8gbfP2Zf1/G5fuoIXUKEFdAzKbCLW+15nd1MQggyX
JSlw0XsoI8CGBPo9AcNFDHwtQZRNMIZ/VfMAHF/E8An0CsjuqnS7yUGdlKn9yhv0
3+TLh3pU+Nohzvb+BemEOBz/X/LW8W0YpDBDMVJPnsaYIKSqgLmiXyAxf/rzhZRb
4RqvK9jastMmuf2n4nw+qKVkiwjmvtmy4EwGTqENUWR684fAc1WcUftnyFbCzmeN
q0ne7e2hKUUU+CfWmcwMYg/YEtpGU91hjlRzPc6s8uPkSciG8jof/5pNiSsht8cu
j2PUdQGWLVfUE4rktPbx7VKQVac4cBefrr0UBElkLY5sFilQbI6ED5BE3K590QQJ
Y8FD8sVc2qJYqiskHlLEax4cTlalj9MhaXi8WhjHyW1Wt0BgAO9tYJdBSgh1fOgF
AVNK2bl4FpF9Qx21OFnIBA==
`protect END_PROTECTED
