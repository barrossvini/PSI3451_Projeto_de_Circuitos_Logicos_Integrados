`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
clhKLejB+i5gZXoeJt94ZCM3WBVOyo+ZA8+QZSYyTBB0RITSzAE79lCoBMyKXMLn
KwRMG6Uy8RZXDGRBsOQBOzlAHPwPKwAEncyBerLTvNvsFhE0GroFEJR7/BC3SXEe
2SKdZ4O21dSPbKuil9wm5NGmolUezfzYqFszVVB5BR1ASYzdU3UrMu0k2OKgTlg2
+89sraWU+gzI64GWUrX0XOmJ9UXys6uiShpAvSBvG9wi5njt9I5cVvFGejdQ9we6
o9bVe6VH9dpB+WB/2aHs6hA/sbUa5nV6oeMTU4nXI8vMD3scbB3LY5L+eWxskG5C
Rk3ZceN4Zj1FPi5qjBN7LPtT07AX3a2/4hEUXEW3/wTdfup8UHohIi/aGbXX+YkI
QwG/H2zt8pgHHY4rBpaT2c0WkVygRwXu87xmfelqykSMRmtCIo6b8gJ8rlrY66xx
vni90JtoaS8BUizBigpcAAsH69rOL+UFCVOcD9EN42Mtma4t+e/Gd56MEgFjvpog
SxvImtkFZ0zSrGzYHQQH+uZhcldQDHw1AIPzjjemneOjN26LRCOZSNWsf0JzlY/5
bU8pC8mmULJLMerzjqJMsPaJSeCQ4XKUEyw6am4gowPxTKiO9qZX97dFvGo78uIo
abSpflmDgn77UsTgNot8/WtOEV++FYezDJLQVAdIslIHQjrh2zqL3mwbYKVonQmP
bdxrtOWfpaJuyNKMSU9WDEnH2MA4Y+YkPA+ZM4UjJgBPJTecZNzkp4hijz06puO2
iropvY+S+uYqObHcx6hogfpCzK5Sx8etNEN9akTrr/4nvTXhvIAT/Azs7TymeY79
bRWytvpGFbvPOo4wJE7sLlqDkxlbGqpAfYybEJm9e8tmiF2RYTQtEP8UEa14v7jN
pNLlXcJMwk2hV+/2G1LL8zBnX4PE1wvXR7daiGI7+eI4s1A77KIvUXmiz5e/3igR
Rni9AcD0d29g3gX8nZdTkusPSYvXweiwdQ33HFEtA2+upL4hVZY+75TmDuPZe454
cnNS8eUpEhbyYz/+1gkapQL/kdpfZpROGpj0UqyxbLm3gxfn+soLHyALWc4VH20+
xjNgxKVpdP32M0pMldW7wWrBeFQc0uVhw8UynFMSBnqYb+0bI9l/3U0VA1uZk3+u
42Qan/BWxHYhEmYsrDfIz3oJtE8RdciG0d24SAYlnXHLQRCLfKShV13FnNNEaQas
DYY4rdDMTlH5/ewVhLw91z2RC3ouRylRL25P5g7ZhwzVqpP9l8cHTHKoHlTs09S4
vFc9ZUwh7KBsjkGwUpqt1sQVVO7Di37K3AFzs46eE+hNmbQkeyD9RkdZYygsKhRe
nacLasIFwJuYn9buKPknR0IbA6bceOIelPTPllJns5TybfPMgRpMOo6Mgfe8lU/F
mhZYogLNOwr12lNfqyOB2aJNQT3ud/Hh0EbmQPHRDhpKUEjBHo18auK2jJ60Bson
psypvBdboj1UYxT2zJ7qiQCRN8Z/iIarq+ZjaNdLmzRxJ/1O2q3agQXjepR6a1qz
wPd+SjdHrlfuMUkHxwACG8SpXX2ni9tlYxnytOAqWNNHynB76/ymLz3IiyUmw5AC
74ntC8l5562o5h6rvt/z0uegFPohUcW/FNAeJuMuDg0KL2bhuwx/JImHrd7cbPG2
93LVfqvuE6LxFDET9Y8zPdNZZijQtM/S7C4/zT2PT8UfQJ0BHDoW0gtG0jd+ErBi
dJrcFnuuELGqnLihfISUbji4Iziy2yJMmCu/bn2yT7Gyu4N7jO+NxYXqgPT7l+rO
ZBJWQm2rKCAdoS+NNRtHEqRSppXtqVQn5SeqzZy01X4cwaTU8hs5FozcJ1BU0R5j
+7NWI3IKagRJJ7+9iaKraY3VSP3kCux+5q+Vzg4lqML9qsVOGrYQ770jYmE/uGiw
rST0sA7sBK+Q5v/DLV9lg+m+SkTFHqSSc1O3fsKTNLwqv+Nb6b7piInMfFeKbuKC
FHcKwrVZUWYjtykUEKjxBOlNCawT1suTRfh13tk2srJpQXvZaGncTd7iqtGOtpGu
7rVY/BsoEhG6G/fijabu9pF3P9J3m53bz4ptK1OOd6T9/n8fm88RrJ2mWE6EE3FW
PZC4cm1vNa5WEnHTD9JthMUU0C3mIksgO7DtTam5K7lTtJkbLlOryPrD1z6O/2XC
qZTcpeCKR7BkUGqkYuNH8YZ9Ase+13mNiO9YcH1ZVUN5v+o+fXxWssm6VTFs7wEU
vzeJL4CoNrmW1G3Vm4EGvZKHVgilcz7tlo4H2p3Kb7hmq8KLRburs66oH2ZJJdLX
9mcmXodQDOp2rXbV3Se+Q+YFrilxEn7HK22ArldePCNZ/rO3oTYJup2PXXGyEtYb
z4Qr4XQTcvynND0B6SizBi3MTiI+rYyBRPU5wOPz1Dc6o06Ft/zYwAhmjaQGS+X4
YiRZZE7OH/H0/BbmajslsH6QjxaYcef+JhNL47KMqIRzBwo6WDiZig1uS3e0eQ7v
gyl1t9FjvIv7id2vb/xet+vgSfvyrf1NSNPy+26A6kEtsIWj2T/DJY8z7Enrq5ej
1eYLMxw4apJktxf7qjWGXIk+C6cE/it0YD8zaCD3y+NiZ+Xh11XghLwnAZw64OL1
Uh8Gd90xow+w5am5W8OmTFZXi+Zv9w1/ojLY1RDfchlEeiR/4uEcN8tMw65jMLga
WM9F+Pt0mmvW8TMdemsRiZAJYsHEo/r0SOWZVHHsm46RNNy4j3KQ9MISudcsIwhJ
Q0IoXDKGoUi2h6Gm9vycjyvrSqpzhb0/CpMTHR53y7C+Eey1NRLXQdYt7pIStwYV
9SgwpKhRDUF3NEmi6pgrHnWp1aHghmvWX+3gohzk1UGhC3MsMHWKdjXmE4hyKCUg
ET3ouzEdDNf+d9MppSNNrJGDqZjeZFe3F5HWbl0TMrEigqADxvIBfgBYF1YJDctT
NNGpStbVI3WDrmJ4NiSTjr44u0qBJi4eF6K1eE2EmRkJWYO8NVsCVuBaEGnt6bwq
/lpvRAgI/gBv7EJgfkPavLncpQt4iv9FrEnSZHjK+8jfJeOJerBOgz+dfHqkBPzZ
w3ez2xQeyRQ32OvGpSvJOFhaiuhoL+m5a797FKk66jLqgz9uWWL7gy/fmUPThN01
4Er3gWtEHK6fm4wluXn503FzHCABAPwhTwmsMZl5sYAQ0MjRlN4pC/n1ptK7n6nj
bY8JhcvGnlwgj/tIOrA4UbGa/k8BNMNVvqoyuYimKh4h0Y3AHiKdPmKQSmDLOUT2
bpL18Ae1PgCEjV1bdHn6BQ3TYbAbovHobTqg/I5px/nJjfY5ufbFM0YQOO1EIMnq
69zkEMX4PIwF91UKS+c/SxHrBg/oCXn0qIGJFfIfET0yrCSA5wKFm+tme9ICd816
JeWzp9EAY1OHy4OtWlYX4XjTZEp4DKsaZqnaBK2Z3ctGd/cxELzW4+1C4JpPwpNr
qzWeL5kB5OwCddym5ay0zud2A3xpasXME0XCTCKdYtCA6YN8N7+2sUriPkd/51Bl
K2iGIH962BC9W06ROuPOGnO162Ox/7E0yu3DHt9XQHwVHrKOIqiqTJKIcdMUHUnH
tkPetzPu0TZLz4LHPQ20oLoLB3o8S1ylh3rRzDGPWU4kNgL549g0vivRFNbYdM8x
gO12VTvl7RviZRFraoQzLJhEDThA2yQ24AWr5r7/PexjG080CXWzQhhoAcc1xLkN
SW02gpTQ99nrWesOibZFvsuSrlVAzzziuMtfIqqYQ+h5PZ59HMxMB1trBk8zplGU
KR0lrVrU0nv7TYytbWi8F18KW8eVnqwk1gDY1pC81+DC7z4tuSB7JKEgXd4TFCDh
6dpKCa0kbZVbFXGtBXkJqhEWCGiOjSuA01SKPr6Mk28yBgmxJxa2fYIvApni+LBa
Dz4v2nkZhnXaxC1xUO2Z2tVfAincHgQUWlwxpKNeZAevW/Aupv15S79S0N5cD70a
F8S7E3JpWW2xmJWGegf0M3USy4VM+iUL2PEE6fag1BaTgMEjiE/4pZQio5MDVFYX
qR9Sx8u+ICaPQXyOqstiuOz/YOg/V/OgSfhTnB6XSMqV/2Tjgh/5SFtIUDEVrai0
sNaIQQtku+U83/RZ5QJGr0ZN4GuJ2OMF/McSu7mVtfw/LRfHeA9wcumlpH6VLGLT
V6aT6VL8M3W/+eUN/wvP/yTjRpHp0rUOhF4zgVWavvczKamFOo/V8UMWOkn2rLzq
AJUVyOtfU+BTN5gRAqMJmxt2C8Jc8cCyCA6HMyxQgXaaQ3Uar54q/m/MFWNduplM
3USI0MCWyGQMzhd7scSwgHsT4RKuAl+BOry88TCxXrGAk9LCKORVtGnY+p1HuSIV
MhWvRGNRUkIX37Z2PY5S7Y/ZSBdx8MOGinBdcLYsxSPnmtbVzpauUKdgxeKcLKfb
55Xr8DuLLMicrDvzWzA6eTIqUzvFoihEjqUU7SsagW0uU/ZMiHAu8SoP4mN2IdIA
utaPq6ndR96gUVzXicgKT1f0WHUuE8UzL4wtsIwi0e4uTwTG1d1VcShJIbsxmnLN
l0xHfIXQ4tQUxfRTO9mR7noRS5E7QAFahTPlVa1WiWA9U5X/ycSW7IK8lrfuOhnV
LXa9dx16+9fpX4N1GTGGWLEaYWJplMoMrAD7Ob5M8Zr0x9ub8HYbvYh6JhczD5Vs
PfKuvXAXvdOKZ9boQG2egWjCbhBWHNyNutCw8p1MCsv9z6Oa7NiIW273jd3QChuS
8M/dzP5We6e3N+I/uCvV6stQSpbtbJmDr2Gq/c0AAW8PvOueOudHk6Ru0bwnZiWH
3pfhFGvYbL99oTpHZ4+3C5+PkwDoZsxewl/Q8Ad2pjkKPU+mH1GqFBa6Hn8yR5yN
MmNBkWvjXKoMqIsE8UmGz3X5ATEJ/ft4Kbtd97Zik/JwAK70O77vsroD7cxERrLq
J+vD+9NvNAjTrvqkgQ2Vhc/qEB5r0VMcTS2B5mKSLJN1Wg65gQRcGN9t8HwFbR2U
+9JeEIMN1af74Y97H7e9zHZdESKygXRzkfvyBGMxMKKwFZX2sDJLa37tBdHLt7ro
DUxKq9SXnQfxtP2GExvWWGoWWW1Strxbr0Rdv4SGS1+mOscf5IlI/XMt7T3ChDSH
N0xwfFmZVzjyByTvvAeGfMApAOCEHo4RKC3W3obB6Uqty45AUFjrkdXgp9CKku4I
0FxHefnUOt83CPa4dqeorzhvzjxldM9+pqWA0l9ol0Tkxq5+RWvpv4mEqxU6qDyt
PIV85GiiLOlocVl0hvUnm3PGGLo0SR5mPh0l3540Kue366LG1QtdjRovSnxQP5EX
/w5jZFt9O/ScPUDRfMji+b2HLEiuNciHnpunNBpdC0j6xsktWWUZInUwkEGg0bbU
CuLycgcmvKdGegvotyzmy/P6JzFVTXFwZE2KP90twu+BR5+gCcW3B6U6tB87ZLfr
OVYu/H6phhGFWDJv1zBdiVqpHvZzDbzEbDplNLLiaAsInIA2It+3QXPzXev7y30H
vFF3LXkeIJdB2BNuyeCfIBIHOhqAow7wIsZwG+dP7BT/c2ztSA42cU4VEGRgg98A
9iArkICX0lrDXlSYBhUmiKi8vW35RZl3CSURRCWgi3009lMbEGgIzAC7+v5IwgFw
amQBwMgKi8jELJMtCxQ1PgS/xE5NF5wa62XKdLOxfZNV24SO6V2CmXzzQ2iQWYUx
TxhJLI6t8aTkg8oqhNVTDRw/k171Eb7+rfUFH3UgWo+1wEl03xpdcJrhpEvxFgJT
LdPwJYG0vS5xpR0f7SI65kAj2Wblpmf3GmzeKyIO+2dsfgr3iEk1MkGFqz1TldYT
j70Oo9yYzsbfY07dlIdRsb89GcScwrqUikWl3TsuykeqKJGh6Y3NIGyRLr49M49m
59pKADua3Ru0vNrmynIk68xfHgz7UA+/DcHl2ZVO8c3qE5vG8OqpNFaObCECZ77o
mYWUs4ju5D0T7uDbWToY2STaD6KR3ZneFJP07sAG+kPLmiQbZZqOdbOeo/uSqidL
6Dq2FQaqkGVM63WWBwQMgvSBHkd0b0ehVp7paKo5816PVsi2365PfOkNadBFR5LG
jqrdvyrQp/K0m3Q6zpYu6/pMk2UmKDnC7F8jkm6oWfZotmDpsYnUPtq+ffEayu7Q
t4ipPRv+mXPzvlMcjcD4O1bp26KS3JG5Ax7UzSjGkICcsZZ9bwid0pbveHOwLqou
gZdASuByyBKlztMN4kI2Tj+1n1BtJ1OZS2zuxvhu704HRjNuEbZ8+C1QoHuhfyjB
ral0uNYCke0NvDTAOBIudeonyElbZsffykuzm0vwr5eVQUHB94tnctzbMzry8JW8
lPd+srySESAPJKlhapz5G3wxIyJAbCsdBZN4466R+EZg7TTVz6CEkW+PRntjIXT6
p9pTq7Fbnkhdz/roUgQroQkVnumRkxWQ3FhN5GQ9cQnQB93ddSM20fbn64saxxgT
lmUzM2GgakRxOJ7vwOySMi6vM2FFAseEQsZPFXiVoVS8y0hIB2VIveo+9ROa6VTG
w14VUWdd6FRSfXuKDEMdSKVThrRjPSW/j+U1KPlL5sxGgk6JJVVQW2uBtn4Klwxg
hxZu2+yGt1tFeMHWrVGzu5ccNddJimJNdShijXTSyXx3jhti59Syl9G91MPC4fB2
A4q1P7dIWuchIbbN2Fd5ow0qtAKAJvmSaEPQiCLDFPFtGj+iMkWS+EePKzmhddpR
Xe7/owcSANtnjt9xGhkTe7IPaGdmnAzhKbi0owSbG3OcPRUv7mcxtMkFrYN6t83u
OQTYildN2gm1qCkmSiaepL5ALoFnm5v1dtWkXCyjHd7fUrRpabcwLdIsJFOc8nCN
4q+meGXFl26eWICJw2kQmE2PkYzrwMr45ZL5Va8UDpd8ubGiA1Gsksp5jIxiL7PF
VCIMrVYyODStrNBC8f0qz/rC0L4/ax3wKgS72e+nuAkfo7FMfo+6ACoOgCF2Syhi
ZEn1L2RqMGu0wo9GFIfdlKs6Dbc+2LeGRASODRc5fahVeAGHWR+2zenPhy8t3iaT
AnmgDs3kt+z8W89CH3lWddMhFJbywFp08biNhL9MFSvZpnqvlsA365iM4FWdyxtm
njbBqRtJI2IkiPrXjIrdupjP9x5RQ7xRSN9jwQRwh7mWVuXjHb0DCuaBuRr5iYYx
mit2oHvn2WACKmImyb0o+X9SfHWXo4LYlvWjy6j1Ub9vZBuhT/rGupe6FWow32fN
Fblb7fbtONJpjcOKboYc+KESWe4BF2YYW1WnUeIkSUU4bSsFVMahPXw9DqJ26iQn
OV7aCHC1T32rZH9wkxOw2fLOBRmzTjldCMh4GAjzmzM4dzx270b9mM5xQ/wyeOC5
DP1silivJEgpN2UxfYCEgtJ7gVjxxjBoq2bvoXmoNfnTlWmM3aaE5S8/Zpjf+lcH
Uzu9HHDzHuCuML6dvx87ijXxWiIc9C/el6VCB9i1yDPreWSLNyyLk84Xp5seX5lG
n3teAyYKYA/xEdG8IFZFAstg+vvGzTpmM1DAaZpVyBYcKYFKSLAkTmLZwoegK6cI
/nHX7nfzRhgU7i18qXIcFysgpj6zhAl51sn7nwdmVdZFVy7e3q1vDAAfslZrGSmx
iH0AesBgslyZCxMHWzaq3Clf5Rsgk+AW8IO78YEplvdlNPgwJ9iNIJptaKNVT1UQ
woY2X35I/CAJTmeMDmO5U5m0N58UYRxE8HtmX0AqiYhJGVJleh4L6EAaR2lBQ3tC
3TelbD1TaGGHxi5jX+4o/aHdgWz/suWBuzIpOS6lJO4FQGgDvCeYR5FuI0X3ywiM
S/uC4sKgEF9/HkxFKfyx4Ok10JyTcfwUHplLI5sK+xC1Kw4RROc9OqhSHIlEQ22Y
r4HFO5BoEr2uGvnDBoglmvFwwbtmBAKqE8i3jUs+za/UMRYKGQP7yTOxQFnTN8pW
KJ8z3NBX28+BVMgtl+SSkRUKcWcZsRJYcqb9+UhMeJYqQthukaLF9pF2TQugyn/G
ME0A+IWDS02rY6kDwBPLsMK0mxX5+N9ka5vPaQu5+E5GWGTTIVpZ59UOFmn3j+Yk
YqyeYuAterZNacyDfNGPJbigXSxa3s5q9idoNPIhPRS44A1lJDeyxUaPXeD8Sr91
rW2dk6ufldlRzS/hvfR6qz0IL8w1cfg5BEAkNXke88PQOL2IkVGNhyQ6mDzcl0xk
pJp3nNRJ2PlahA1LlIaM7BYxa3ZBQt6ieQnYOcRr2E5exDHc+ayEgyUMld1K2b/e
J4zMmSNIWThyVJMByjy32ZzQMdzPa5zHR24nELE2Ev7Hr5LT2Y+RgLRQ0CmGpoIp
K8p9VlJUcabJiD4tk85avfW1olfWQ6Fg4GdQBPHTFifIAvX2S+dorxNklhs+11OW
Z/3Fm4XA/UVf3iKpgrMlXn1qJMYLjPyj2EB8sTO8NgrUAOd7Z+1GYbkBFwaAeohB
7i8N92ivbsB7nZX8EDIiTbyU5zR0mpTepFEvpAZLthMP5FixDlbJ1JpqmqXZd1ST
gEvjhDbmlWy6HimwjIc+iiJQdnw2BbB2XzefpGzXg5qrRMtKrIFiGvjH/uPNY4/O
VZ/G/N130tPvjRutantiaM5E8BJFMSp6wk/Yr8T6xgfkZrqL8xz/P5ICCuWxxa6d
bJ7eej2T40H8d35vNNsxy2vdMShvoy9IbKt6Fpq8GeNEblecib8FSQA8CVJJa8yw
5r8pkrLjtDuNwVA6B9+SrOPGxjlaBca+uhnybg7BTYa1/1SlPFZD+bras5cGfH46
RfiUXNwlLN1Bev1E4PAOyImUA0edAgDi+Og/Uml70al+V4wJtkwUIo4JziAssi23
tlUXVEcimwLVLtxas2hAROyJHpS3e7Rzychg2VEkhHw9FGjVK1EAnHAHsPmr5dv8
Tpj8L5Ok4eEsHX17H2Q1MD8y7TRL4aFuYB899u0eR5UeShUUyVAhYlzpq6q8S2U8
GohwazqHeQ315Bwd2dWRyrsPKI1ViMXlDuA9vCNgbQ7/+7ILBz/wjAez8wc9boaD
uhhHbSuvk7Daob022zQ2//jKJh6uMVdh5lUcCnVAa7MHSHq98kkJ9mDxKhbrlaJI
UA5bi7sxBAVsN6PEYp26kIlefqJx0BdO2ronD3tPHC4nUni5mfO0/yPk+yzpCbXn
sdCsTSWh3423YH1jKZbMNZlXUpIxIL5folFSyXHnvv70qT1RJPZPzwzuqgNkK4gx
kubaq5o1Sj//Trslk6jdXwvc99lMdlt+OTSDnpdWfrAtDlqyLhmdJl/Zvg7nS1qg
/vUPWSwdXZdVq82plUlruEzPCT3RzQPD01n16TlWTZaxw8lchKSsN6tlY3IAnh0a
Q4mCD2oJAFPqV6gYI0jrVd4LLpgAmZqyo1Zc6x5sZb48FjNtPTNaFJ60pO0G96Ux
LnOfbh3LBMjA+ZKthEhf/jVCgfmfSZJ9FsK546oyXyX8MkxWHsLWde1GArBQMhbI
pYbkRShBm75h4oNfqS6KE5lG3fUpUHtFhNuUrS92TB10QBhFf1BDL6LrrRqxbUM5
oDsWpUupHgDU3g5MOcV1cRapHESJcsaDFZi5vnl/nn5Wc3gDNSG1RE625cJ9kGT2
SJvEMG4KqfPFpEZ1oQPtI/4p8OF1Lh9E2vbb7sL+gRFLY1/R9fJRKNQ6e6XiXnMA
LjpGuWXhVidLF8MCoDCikefnYC491DC7QyQcSojLxr1rB6hfJpZa3g8+d253v+os
t8IWTiDgN9hNfnHeB+pYhOi17nE0HRZOE3JbrFFIeJSmgSoRiQfAT6ZuB2j+4N56
62teT8SJZ/xNvPNqlcnJzt6hAiRQIOlSbZs7piwnZWa9dDVJ0nZBRysthTP1wEI/
z4PLPcxRzicBcwwW6ayGN9eMcuEh2omf5V+tENmy7YIAjv8ZAtt8umcDIAeoUHBX
jkT2rGE69V9+s8yDqMqAHUsNHqUUQxSYK/NCAlgEFq5vQoOiNaN86doKpEgJd6d+
pns+On7uiokRMKdOtguU1QBOGYgwBl9VeRBacJr4HVLKo/Cu1Nyjisd//1hBCTHz
jw2o5QCANSy0Nj91aF4OkqsRDZ8UA3eNVO17+h4izov1yVQ7FgIR4QiDl5TVpzBY
5Qm7kN3BH2sB+9dJnziNKzznPCDhX3ZfKxMTY3P8pE9FRqUrvVucLA7QS56V5bu5
sIcVoQ4Ln1rV9Z8KV+y1nFluHB1FqKK44K24sSgOSKQhjWmpJlK/3ykC+ujtoAjL
w26PvlE8UFRD5Md99ZquWnP89FGSR5XhmZY+X0lrz6Uw+zzYThC4t1Jm+YClqwYh
85KW0w6VuLF/7leKN2EVMSNJCnSr+H/TgqrPXm/Tgw4ur8jdj00sc/RaUNEmT3T/
FBt54m04FnmJgr6kKodbeYVlaT+xFKVM/QdoaWC/+2cx6m2+8P3KNBo8rFfKC/nc
XvcEuDb5bjT7sShf6XEfIm3ZCm/ZKj9j7HMrrSd/EDBBXdx3GEzcPbxi3oZYvRys
3+cGSzX6P8K1TNkPQbqHLd38HsaRqbBxC9r0wv25+8rHj72a5M5lDqTl085oZEWo
6jdr5Rttr4xXf8K3EW3fFgYNDQwB4IH6+6CjVxNkwR0ypbNaPB6U6VGBGGBT/+4B
IVnMnTYyaX4dpF4koeDT3Z+P9zGk0p2f//Kp2AhC2vYa6HvqZmRXtjk1jhYlCIM2
Ip8PIzb7bwaMQIzZDFEFKPwQxKN+OQmdl6wdV7kTO5dX0lf+769dhSRpi/Mw2GWE
Xf9WKFl2of9U8Vh5fwOdX2XqZRPuS5rf7TCGipXlZZvptLn61DR6FZMFPvDtawhY
i0u/Mvk7EXPLK8UtIg5MNbRBgxwreJan7y71r+mWLswNlf+wCe/DrQxogRhXm22l
5sl5AoAhip5g0GWiT97hhyikcXkOu+HPyiOD3H/eSWcu2NjLgw0uEaqlpvDN4ljK
zWX0TMeebZmGINUtodJLM2/39aMOeHERNq/KK+o/wQ8tsepTcKmIiuj24i3DLrQB
4DU6QZCXTcESpaL4mNE7l/m5fbyVDeMK74R64DphGW+OmyK0Hwa3PV9Bzn0sSD/H
+6hO8y5+tPz9Mwh2wJIomwrydC1tATQj9115CuZY9XUpAZDMD1kfffhcq7leVQbl
ZsRyUaYNV5UeVT49iurNGmBXKkRPqKc1dPdm5oSGQzQ1srzBshDN146Z30OwCE9q
+PEPlqF+Tcim7fDEnNkJ0nKjeJa7xAyI/8HF1iJnOrKYDSruUghfM3QgBeIE+Qsj
sLC/aL5cbqkAhVulr3Eu14F5lG5v6UI608D0YGxCfV+85E2dHqlT00LE8fI8luBj
tcgn0+I9I/xflNrA6G23HRAuUhNtVWKlGapqjcPrejS3helvv9A6yTpZTFdfp0Y4
r0c+PpQ6SMhwVh1QrRckIq3DVwaFROguTZhvGMLwqtHTbqW75DfVjXp4UxlRM5rx
BAExqoNmfyPmuFb6H22bPy+eDNz5z1Tn55JTFu1/RfgoVPnXvh/NwhuzYo84AqXI
LWtRBNlL8VkdyjFzg9GJ4qbS/kyczkGyj/FY2G6ebHHOKJ2Hk8b99RsaY2aPn2VC
24ow4wF/8mS0/u5rxMF8FRb5P1mckq8pr3a0zQ+NLTy9XdZsK/eAzEHSHbFH0cR4
dcD1uv06nNiz8pdOuUuZA4qJK6I2fh8S0LjwkKieQqs7ht0ogIhqV4McxCoF93Ju
pVa9EgeLquCktc1MvDD1/2Izbfb6ZxNS+v0VjvxKfXhzWr2MnBbFn78b5gqLRYo2
Ab5D5POJclqXVOk11gbgYhcqC4asX4rKM0Zxh1gM/klrlJVBlMBKgnEZWkQ9V3nD
9637rhSTUMx1IcyLRBDOY20THM8qb7toHM21bUJGic94kfUb5Q3UXoDx4jASwCjq
BIoW/lmJF7Vbg8Jh27bdAxHZDMkU+6RTbAzAX8Hqh+Y/Mu/MCrf6hq5ReCmD2dTP
hNsGueku6kyM3RUG+EMouCtbJpmL5Q7mjAtL6AyCZg8WJfl8F5M1o3VU/xY13EjS
0BH5+thnjWM0baWaYreV7FZAQOc3uknHh8A0uzcIHGz+/S7coifWMCjR1e1/YJAv
MPxzymwD55SaAynsmnTIco1T0EDcE9dLJjssJmEUj05Nha/V4cy1jczXic216tsD
4zHmOLOrI3S1+xnvechG6Os7kSr1UjJ5mmIIh+vc3bo0q4wjRW9htSWp7inLUvmE
rtCbWQ627HaYz/QQxv/UQFfEKV3Hdk4KDU1DZMly9rbuM+YIF4A4PDKsSlg3iS4t
KyJxuWBvthLtuAEtmcr5N0y6OYlgvxq6OugWCF26VdlHdFEwWwgaPH+cg+ZMU6M3
7Ag4n6C04zyxx1Rx2B4hD4Cdc347ZZQXQIi1/BPKxfkh4vHVZhbbmZhKQacm2izi
KMKQTk6WWdhKKP/gcgZx2r4P6Rl8ITDQX+tLA37SHKkL5czT5BDD8xXbDf9gI9ic
Ht1SC7DBGc9w6uRno0Aj94xNkxyganIjIXQc2MNEEQHAnYlr6p/pBZubQlQO4Vjf
c43Rh/igFWZtMslyKz1rUUTriLolXc9MV6lDXTNMgzOKr/rZX+HAGti/NbjYoVNA
dGSicwo7GAxvTT2DQl23s34i2v9L5SWGeR9koxqCCm1qLHbUwsA144PAWXz2Ur3C
yZCz4+QdDS7hfCFHeiAB5HONTNVOyIzyTBMY/j9EKxh4sFRrrDN1qskih7MK37Sr
BYOT+vnEMZ1hLnDljgYPJDWqnSWaGjaj5gNx64dmHZoEmXklsvnu2QuqUUe13Jxk
zFQ+PtWhJnB/E7iwsQa8mTmN+t2z0UN+4vSulCzBXgEh1wlYwNVPR7tfpR4rr60P
u1lVf3Qp8d8zOonHoUu6aH5A3dyod/a/hcHpfzMTogiZcYaLsKmrxnN8vujX64YO
jtWsoMXracCGH3EKTXD4bDzueuDz/CWgJVYekqaaSDLlOM58SuJGpmvWrq27pgMQ
ske3x+aq/w2keS7+2beYTwwQP1txSdbL+f6z6fsHz2/zPmYnuXituywJof/DVc+M
CePyA9PBbX3jGC2lgbhSxzldI32iVZtzZXUbfESN7jAzxWO5Bna0hrMV6cKN3Y7b
UKy+xqObYvgPXhz/JIsGlx2LzgyZPyjS6fbrn6XZbvhikw1dEx8FgWikJfFtrDRU
Um4/Mlfq7ZHwLfbLIAhnFhUdDt1HHeoTWezqDCGbKvZHZRPFjkNZTa1N0UwKbXYb
3A4vDBT5yUcOK74rxAQOf8Yn+fdCU4YfaEzNT3kQB/u+XuRCS1vnFn/tSyTMxb7n
0B/qZ2CNGQlPu974O8Z3XVt77sgYveqtU8QcrfmRzNxPCJ5H1kvbr58ZvMa/dmc+
sTg6z/TpeYcvhhL7GTNcUW0//o6jX5TKd4EFFK6GqNCC1IDFZ+lM17kM7Y4Ir313
T/xLBZa+4JQGAm2bR7gZgoe6B4fdzTjE/g4xLQ7UGA2EvDE/Mldzn/1qZl7A9Dxl
pIKbHixcKuDq+vKjFgKNPdsJMGvAxJ2+Et0xifmJgn6eZikBRHJeQIzGvUyJPJs+
myd7gaa2p49vuYek5XxQdEFY+E0XSJF2wLIi0oycmeTheQhHCMZy8MyqaNzkf/41
O8e+ibjsvYDatA7nzW7ynQ9S0INz8W1iLXZ4yzg8lixqk21GohDQyUk8Y9vGRq6m
Aq+08RmglRaPluUg48zmII0GS0wQcdXRf4QuGg8TSZrUFM3cfot1lA7C2NzRRO67
S3Iq1+krxlc3uTjzYODjwiSH4vovzFr9qna80HLvrlsgWLBRZT+s27Zq5qv4HQAS
MisONxvPnCUls8TnGKB4gYvHRe+/uj06zqjpJ34hACxx9qYDj9CTnfE1Th3C1eph
m+1vebETEzxtzvDzMQ/CFvDnEMtc5AIwZ3ehjdZQ2iLKd+xrbNxMnUj12s2jd0c9
xgWPHiJ44HFA1Yn8Q+xZM/EcZS53J8sVSsL8IW5tsIGSw+kJhs5CLYyyNhxAENUn
qvXZzLWW4tzxrgLha1YZg51IBYNWLStpprTVKw7cRmjt6J1xQOPT34NeYL7q7KrD
PM1eeNRIL0Kx/NSRCdYugHD7hXS623Otj0MHtmGWtuk27S2IwYcH/lSYe5IlE8FH
aqg8jnQlsb2fpkMy8RRbBGKi7Afz4G6KIu/UU2+2hZpjry6AN44zpYpHzVMZkuTw
gmD4O60dGNROD9G7bkE6VmIVVauir6O/d70pE+vuMf2rxO0SlKQ1ilQ21UwTa+7I
rGFOuAiybJh/n6oMNamWmsC1UCHfEHqDitAgVE9Oc04wDutWYB5vphuh7FUEsfbh
Y+ZDLpnpagyAqD+Wr53E815CL9V5qZdaH5+p1KBonrr0VXOFEcipSnr122LCN/zx
mpxsAb2fSRzzAOphqDc8lpMTzKJIBX80uuqaRTD40OMw7/5XG2JH0iVTMweOyhIx
QWdYjSjEnibU9jxxVFO4Fg+zRkPhrmbBe/+yZ1XnZIPWFSF6hPmc/2iWUfj5UXZb
HJhLinMfpJdQjEWpIduOviEyVBiPgt3PSxFCsyjC4Imaesp4U5dPFE9F8ji3ryCD
WQgiLGfCW0UQMniu96qtNErGPNf/d9Ok4Y7o5NkeOBL9H8/IFIarr2QvXQ1xWVCd
kf1bBxUPOrzKXJjezGoaRt1y+b/M/zTaX5oSLuhGkhaV4mJk/uhPxYuxZgB8oeUT
ZVz3ikoybEeSqgCBI0nBoYyPajsKvUSSThbnY5+ivKxrEeXklExLjhoIValpGSZS
PxPwbPOBdSRW4Uf2d2sVhx84Sil55EXZYDYww0Uk258XaeyLjOJ+7keL5/2zqoTL
98pvq4KvQLTnLB1plD8ljJekBcVFpvGPNDxGTdd51VBTidnDjHYqTm8c3FNydJ3S
aMWa1vSNeKMdAGKCxtzsEnibUQICv7MYCNlztgu6w6lDkbC/b1XTSimFmCBrKdhQ
4iJkO96AkF8FR8AVcv4Wqsel5cQVQCQzTSa2V/YW/YYcLiJQoAAc4s6d0LRX9tz2
xO+5MT2cOrmuDFdGF6aHksSeW8mJXgBPUKkau0rOM78x96K2bjcY5/E43CNLzvQ9
TqVE7v1rlzTtldQI+8rZSORABA8IonJafn+GqsXKhQimahKWMtEK4P2gKbSGLQfB
nfouqZono9GsRGm4JIrJ2c3PrKVYmcqawjHNDbigO3T1cyAO3AlZ9oHBNmGULoHM
/U9lPAfU0jL0PpdyqCV3oh1gU3Uey1rkHpoikrruIzyCWYAH+46KlosYDKGMW5xy
/PtRyGFaXVk9tLL7poyaWW3i9tyoKVs6aDARKMpX92t3OVd2cFBqDAqQzRYEjtCG
dW6FGlt5jZONo0U97ZNIvxdQQGMPYKJgR3W+EFm/rdEchT/udIdt0ERvV/x79UnV
ke1rHzV6hAWVp5whUB4+5xtwFOQORPVPtHEbTdp7eOLid1gi3NMQkW+F6hE+wcrt
GcjeX8cE1H/isRfX9HZV9OvKZ9bVR6SN2I3FG+0ffgAsBTzteZHWN0BCdVRbwqYF
29hUq+70F1yhrnSHAto0d9CnTg3o0627i95/Ynql+N2K2lorH4LHghQ4cogO2WTk
a0jbKJCFh6589Z5yBuM9ex1fBU5vwpHMvoatyQg9eboTgCmzYN7PLFr3GbYaC8lE
dpeV851rIWBxn7zkPQ6UT/kkqy0jN0f+ylHHecXhSw+i7w9gIyZ1eJf6eNReqegE
97lnJxwydpQsiKkgjPDFKFzShDGgNSqp/wVub8TKbt3m4e9HnBl8WzIczyZ6iN4r
o5KG9jqeQ4q4MU0eohKougkloyrdpQiON9jxOf+jJLyqzOAIdRD1PzQV+Icj+078
e+4isTbd9SCzD4MGk9uOZboCAHVAz+QSQei4sYcSWVMcsshEcxqqcTKTEvNB7Dmq
Ojxp2kIQkTVMSwCsKBYi69AifFOUMv6bPatpIojrYxEbuI3zy77gxxFznxN77qTL
FsXQnlSuh6exgotXV0yCOdMErBOtNx3L2o4esPPXAdthNPuvpClPWUmJOSkdMGim
Tu5qTl9o0QAOjOSI7MiPUI0Y1sbJqmYiVveOrc9ZwaFEVYQT+TcxbDvy4bsrA4or
lGuhb5pUexZgl40xxY6grBn6pEdYpV7/T7r/UJYWGMvaaBIjVBPyoGzzEJLNgWw5
W8malVzrOD5ZN/8paqr9rye7mo6NXJsCgWOle1a1V8JQ6oa1aylTjdwgm3m4fx6F
kxkB8NEkEXyJEzhTMmGHn/5dCkRoP+y10GvVa1QIIo+bYkksVq91SUUFcU3aon+p
47G/DxqsLCoiX9DPKAU787PZcb3dqMaeXceRN3Mg38CBHgqVDsaySy5+RNLzkZt4
50OnzoK2g4/NLkCs1ngXGJf5pCGvAUn5Wlgoh/99ea/MenYmWTYORugj4Ob+rSxW
l0Q0CDREmOwC7SkdZkugKAeHyGX5xVv5HOe6bT66FWxfOBJ49G5mtvMiQvSzU0Om
C9/seehqyxP7oeqs7XAGqDyVukoA9Tt0DRCksDMCmEyNXG98NiBTE+UUhZIAPr+A
rCt7LJ/4R/LpNGJbdkrLflH947ceIghGRfEBpVkxljLmJsmM08zOKZUWToHyGYL4
0zJkcCndiwMTksjw6f9BvxgoNb+lyl1Jw/Q5lkGU9OB0H5nJWA19j+HlgOk1aNpZ
gr6VO+wL6mXfzhNpdh68NeUI6kvVPMgFDMlq9ikEIJ/+I1AfBg+d+Kk4PkPcmJr0
C2OZ35+q3uGHA9B6vuzwBbxInUm1ge79Z2mnGnyhAQ6pXhn9J9vTuzot1s66CJL6
EUFF+FYktuhWu8Nd/utm4Ttp1RdDKX0SQJ3ukH3QB1rJXfduw8+C78oJFcqnHBUE
WbaRozygOTS2yTIaLbVt7+IZPUankRSNIcniHzuTT0NHW1xzzL+lTUkLwW/0XMo3
amsKuDib/hvNdNOJDzEC8fOlh56HOJtjSkKApRrTrsv1JtH82B/fBXvHHHeGL42X
RoDTGd8famnx8PtAZx1/2fqOBAy9iNsXaNPSLJIzSD6GDq2NOrzRoyQhEDIMxDAA
5dVMopgylOx1prTF3+Tk3tqxNIZjQ4KpFRlkFivJuj0Tt+nd/UjpR3tIrVr3GQT4
LZEqGhTZm3U9PCxk5QZK4HIZkQ78SdbCfCNmIw4OeT18W/ulj9h3jM3bz6NWPRKo
IlGUBUC7d0/eARErz6ncNUQw2q8vb8NEJCHXczOCQKW0Ht8cmbDND8fe7SZ/2+y8
2vbMGH3LbHd30dJG/4kkRMr+azbASruyd9lOa/StJvvXf5iBgGn23bpMe4kLIXtf
tn9Twvha/SVSOAZf0O4MD1P9GccJzkzEquGvxMpUq/OAvfDPta5qPpXiBWXQHDCt
U0AzQwwSn3cKyN3dyn/i+oAN5mnS0268eOY3Q32WyMc2lpJakHJ6v9UMmWzooNnO
mr1K0+5Ci26ToAm2460833cEiPfLFSiyt5H7tOV32vFfKBA326K1jTps7vrRzKEW
oqEsxmwzHvha2HK6MKr2kphtr+PH+xtrqeBx7Vy78VSTWu/tu20SitHB1vNRW2cm
4Xgj2flkdxeb6E0OGx43MkItdpQP4K/4zy4R5qd8j4nlRkyfZhaj2S4H0HO1/oG5
yqXfU2puSfTkOlBomPJL/O/o9tV/70FidslkELo38VN0IlOuCHa+noKH10SE94nP
ElnwYhBkIFwVrkuALfuK67yMIlOpjas8OS5qj8MdDz/8yhvZYCubpu9Yx1hg3Vv5
Mc6++jZ9R3P9DgYBXS6mtRfpv69kZULsFmJvw5LyLRBozO3G80uGDR3d0u+zjEIN
wl/FT4FPAxHlim9W87vRwjenbaqvxny8NTSVpIL7y+BbzXBlQPq2X1DtkAdMamO3
xlmN47t4CiNvo9p3otuygycGQHwsW3uE1gmQEAcv8dTayRtfbKpVwNaZanqwmP+G
knJJVOYWsJTU7ENheDDTpgsLGugf0aP7wsfxGSHAqoVXH/Aj92TQHnk26d82RaX1
PoCs1iG1BCF4TQrwgm6DilW6v47XN+AkLsSdY7Amx4NU7ACAQVQ7Bt8HJQoPgST7
J6UBnQq4lpSQLBN+vfnW206Tzl1I1sSP9bXgdOgVNa59wn5YcqZolT333HM6iayR
NkqhigED2Yb98fHJF/JfJd1OGhOxxDUX2Nw5VF2DsryLAB4ssXWmKmRRjHFV+OdX
WDhGptIaaIbUoMqbK4FZxyFspdqr+MFBqWRC09YCU6/Iz7gCrXWZ/MJjMbvFTv5L
uYTutAlCdcePgFVtqwh6TT0NgQTDx+Vmq/6sXLucystLN796VnCdm7I8xRqkS8ir
9hx4FypvgC55RQH1S+R4bkwsdmZofVrV57+JBz2BsfctH3F6SuBszlFkOmy3E6QG
kquVWVhijG9AtgUCMCvnUav0cDkfWyIBiseU3ykhLcqLqjcczhXkLz4YTW6dq228
8Oz8sjMCXH3zt2MgidjcddBDRTt8vvue1oqetLXgm2j2C9jN2OSCImed/pAgy//S
dBYiUu1n6l4b0bJCB/1LeTwhroL3peTNCt/dxQLloqrdfAEsG1asTVKd9TLAYUoh
dSrSeVW4r/EP7pa5l18IwOHg0jf/OVBPBodhXXzKycvA72ex85tOxb7Y8qYJa3CL
9HaaGizyPBPtWxZdCibdOmJDOgPKUXFDyLkqMOrutGKamY/+V7/4l4hgOjH1gB3b
yWfqEAYDuHSUECsn7ZUp6GQOhXfRgx3CsX+eFQv9dwYjHrk8Rax/ODCbbwbcSqvV
aGDslk4cpyUhG2SIX4CrR2dLdCJKrjpu9GaMzUk9SvMPTY+Av2xpQRw0F3cRVUQc
zXTaMTLpa0Td9RCVE3cxbhVQMl7j33A35Luw2mNABcdrNQoi4LG+UnOFxeS5RwEC
wPJDoOiK5Yzgumsdr868qMmR06qKljp/tEitRevUcJWYGmShpHdMcZK8KEhtyqV7
8p9JnzQc3fmbKBaf3BnEhH4uv4II+Sb2QEh13FC7o6bpBejY0Ir+JMkEtoP7s7YL
QBer0r7iyIEpHmcdQeHOnNgPW/QMouNyNAkEkwb4LMqWKb5rpggJHxWuhh5+wkTW
VHinIUL+tUD0r6nuY72PjVOos9JTxXyGQv1oVNFqgqKOqpVkfaJIWmywAcxqxt8l
WhwhEaehBA7LwuYoydzoC4PYcx5XctWs2r++aEx+Ku96nmz/vEhQRn/QwvTwU1w0
TI3+OweCbOhtB/oCPtUPRzYwFzoSADWWUwVJw7pAyk/YXn811VX/1iLhBhqjhF9n
KdKD70v4oUPlsQuLb/6NdOFLEXMTO78KWSYcaHhGfOy922HPBPGLGyxdTa70u82t
SMiRXrz6glksAQb1LBVoHZjiOeN4r6rBC+RGwTh6pqKQEPATxK8+SGfIBcrF1Ipe
cLm4Np40Jbp2aZVCVZcMQMljCxMR+5CACux88Z4Bu1Lq+09T2SWnS7KqbhO61+NF
GwOYOyIB4z9Ppw9tokAVtDUFnysdl2AWilFuk8FeiHpietv4gPvjPt4D9bCFRPqw
gS1hAqdKEFQQaXx73xnq7JbIhVDpy3ueF06uIgSjVqvrJzsuY/v6kLVIIxS544kG
8gxpI+dyf+PWDZl/tRld+ha7HONlcawGRWuOv38fBxP+JbetyFzt2XuDojyHj1TH
vKDPVfns0sQWdWakhGqURx1+ILDv/ehHe3RogadXJqNPPNjA3wVC37b1TOu/XcnA
+OB90y83yduG8X047WApDCy/Z3sRTRl5qaQQXiFC1sUzf/+/uRoHgGLLwz+RMYyh
7luKghtn4UFo8HGoKlNinIE/ifs+fh+KCXx4BKrQM945eTBuyNlEhZoNigWkKr0G
HvGj1tl/iUkalG8Ak9AWx/LBrUKT9r7RPwA6edFXyWmMyiaf/xkBra3YJSYTpRW0
LHdfWqxcvn/sNe7UYXMZtB1QLcPu8vb0oHgsrjaCrBU/H+POlt3IPlbLqyWQlE4y
HyQG8rZuTTBkVZjANGK7vgwrcUVFd2671uJH0rt0vtjfAyZvVrgpLeE4CllpxP29
C9+1gLd4+9aVKfVUZrgek6KJSu7jAqWfjMGzSUYS679/8Ea7WOQv2vIhVGHCchRM
mNvMM4qGZ3fDJc5naXbmRfxp2IyYcVSVg9/pIR0+zdrSitbG5959ElY95BNxit6m
ie7PxW4Ka4LmWG9Qjwa36hSCKkX9qaSw4NXKdktUGavA4EFA3BStcb7VT80zn3sa
MKaJQ1jFiCB1PYWHjHUygmEufez6lzYDv+Svj4613V0zqu2pWAI5nM8F3rCNo5le
slU5i4Q0TQNLLAi07KIsCslUXQdCwAOveuIbUnn5I5JbFt7FVk2IPAhOVB6GSAHG
Xk97xfTva+OHMMFHcno5D9XGBzeylr7NjBM/PLoQlKcV4LpBumGc77pbvjIwr2+o
1bUxReATldWHxFbvLUUca1R2G2bzBS5GqjjMl0hOU5WhGxg6WDlYeCFQZNciMS78
A52PutgSoCTWrFj+xppRio3zgL5VhJ/0ceDsor6r+20bOKvH7Ln67O79QoCAkU6G
Swt8LEeSeLh585B5ZXA5ddImkdXusIwSwuBoLaetXxfpgpX6ZbXwClZvZlEK5u5a
gk7m6RtVb7j/jPuu8exOMyju8g21OmbesJcf87XctzpszfJdbbSxyWeEY5Xro+bi
Lu8fB60iyJ9VkgqLotp0YtB0XJgPpYuwOwnpQCH0mM2day3pGeF5dfYOl2OnyAv1
Ii1CgoIM6YsRmfXRa8Z+SsVR4TVGLLkkrYKzAAHJcQq2Kg2apX/+5Z0DOHGwkxFu
O7r408DhWILuLN3iSj9soMqGDMgjMODeRGfnr00EdZUtP1mEcShFYc351tyQDKL6
19dV9H+O4KiR9JwTGk9Sj3cnVtzCVkJoQgsDtx6dVzs1nqccP/HB1/bFIcLLOq/v
0cEvC/1irkVkk7HwolQYiKteHrCuCo/akMNHvgFVQzhIIrUqvsY482tW0ay8EVDZ
mb2lQ9kI4QWOiQLazZLDwYLavJTYv0PvjmVw/Udi9OxRL536t262HRLPwn8OOQlr
xA5XDEoSNl9yWmNy3095NtJIILPOnxikKj1WDeXazz87fATuky4hYDz8bndbpCvp
07SOj1BsCKRq/ez+2XDD8cUcC1OQbuT/1U6/T39Alf2ReG0D7RH7PkY9cuPbyfvc
9jyx0aRrwgBxZZaycoGftkach6a6CSF627ASwJ1TPfFE7M7ve8kp3Ki7SasUYB0y
uDlpC1PCT9vnCkLro8udJLmoDka173uOXUVAQEGWhskdlgjHYvbzwAwN8rrzuwVj
/Ic9qBklyJmzc/0giPj0TsAK6dOz8sPmSVSy9Xcs10BO2ViTS+1jMpHZupQLaxN7
pk+LGFcg3wF3N2nFIFsbaU2QUJBKhniD98qGIfnKID5TpXGX7WDn739mQHJI34n+
gJ5FMuM3I4t5eTuUrij7HSmMxk44Kd60XrJkKlVwHZ4Y7KqMlkoqAx7dXiy8oBd6
WsIURZ7wixnYDmfbW6NytEWQl4rs2NF/exricz6hBGC/OuXz3Fn/lnhK2kmVzc7v
dlnZEB+jkkWOYOMtFwtdY6q9SQripHikaYjQPd6Y2X1dXUbu1BI8GduE+D3JXC2c
Sp5k7nsrmnhN8TYzHtE8lIagV1YCACRMeB+RXIcVaS9a6uzllmPglCDnNksUAfi1
fNd9MK6lSQqrrQMjGwif7BE5tgOPViCh4SzXHSXoCD9yr3hWl2luRictHHzY7456
EJmatsUxZEYx24n69Xe8GJfZ6d52EaBl11s5Glpt/s14IuwQ0Ng1NXY3HJqxsLs/
aSRuVZ3X62Uc+CSNd3lezw9Yh3PRcUHveIONGEpYky3yu8X2zs1JYkGQWyXI14gP
OWravvqE6DFO55cngbzaY89hpx1MeTnb1af4+htA9ya6IL+G0CJBzpDMDiW0tPdZ
Vacg7Z1VzIlK7tKFOeZR2oTpAjNqt0RroYcaOpTWIqFOi7HG2+ZFFuSemC7tLNKe
u5Fb7gkurknIizfsbhMmMyLDMI2vN6926u2Rrk91XmXf48DTKUshUjP60dCXNs2n
D8DYjxy5cULRwy2u+C2KueHesIjcnZ0CMqNT52iTskiE1BVNhcr4rWPb735zWsit
jVjntiNsNCVmNSWsdCClQ4kNZW1GAPWSNQBsLinxbBS4Y/6U2/kcHKq6aRcdzBlw
FxuMUnOTYSvj/qTYA7+yCJafEgbWzInjZwh1PAKtvod8bJ+sNjzY6jSV8U+iCgkB
gq1PPNVksI37SpD5svdvcNsmznxUV7BucEUqR4h8jXObKP0gnd/b7W2AB3LljaCE
0hpQGzsUr3iwuXFb4xBFfINKk6+OUaJ5gFqjA2h/s0vzxEbSW6+SptkOPOO0/ePX
yMAhfO/kjheaAr0EzpARRSjk7MDTfD9I+jtSv1xNnbhgfqSiIJTO+UhrjZbivVdA
hbIvxRwcoQUlcPeeUa6HWl6N4+jVNxWe8ZN3itLOhV5oBL6y62gsvNKL9MEjuqQB
Pm952f7FcfhhTUz1tJE3hEsELBgu2VZLca2/kl+r0bPpGPE/n+506ObxFyN0CuXy
fZf9/umnBlpHTSwXXwb46ZLRxpznE9GHvUZ1Sew6Q2yTI7+yJ/J+sul5qXHJC5ua
79IqJq55vnYVXgFJ+MR1lzG0xBnESPPG/89E/sIR88ad3RFkBh4uSdPP5qfYh/1j
q+40Ti7UycA0w29f1ag/okvRou2csKC9AdsabCcGAWKhJvmHYOtmEj8Cuz7Yym+o
1G1v+MOOtoh1twv4A9B3NpNEEBXTEhbVn0vlQtwj75kypunIArMzG8c5GTqUfShT
MvABAKHZT/tQG8T6eBHNGilG1sQVmA7A3eq42WsL1NPd4ORT1lIf41til7loAhVl
EYrMAmteoYscq/jK0rT3+FWHdncGCCzTX4URYe2Gi/+D7SawcYG+dnpg5oHgmvsc
jruRguite9Oe5v6qhBCDxqXM7PY914uaQh6IlExrl9F7FJssc3CkSUSBpvzRFvk2
GuPG8bi9Lk6+2ADO52eGxAihUUZBcAUmFBM/AX081pMmoe3sYNsg7gSn4bKTU6gh
Wsj9brRyRnCj8iZxaYQAmBtRZ7c9wajcfxisTnl+Cg/mvmnwiyYUmpZ5FOVxCpOp
W+2sCs0D7HhTkUqSPJHCqaI/y+1dN/0JfFgAuQtB2FmIjilrBGSEOD2SepZFsAeN
2L4/V2TK+K5UoUCCz7js7W89peHF3IBSRVD/ivB0hPWCsrv/MSgc+dhdk6Bc5I+0
ysgz51Xt8lSsHvheuI7w9wb69lm4C5JnApzwIUmouJqtXWCWwZIJvOiRIQIrAVuq
9yQ4Q/y/+1kUCpyGNPafkvOK10VIrD8DsMStpFf3dNDQeUdcoo1euqrOXVSNYPip
xFa7QVPTZw83YMdAX8PpA9uF9kOcThJf1P1MddysOr1D0N5ap5S89HSq74w4wdm0
9GZBPZcTz2O8k/fXx9FHgofQUmG94tkEoH5coCZyW6aUcHksyOApM9PNGUHeiZ4E
EvaOo2oLICEaXSQBzOpxwbe+O+kP+/3ZM17vui0Y7pTui1akV3PLMoAWw2NUkIb9
MxxHSRb1zK7OVAcYMyJNeEEW+bDDnMAWdR+iHbeYW2ol7ikSVFtnwzfun2xBVX/a
Jt5PkJJFtpTpl39jOrj5CzO2ZDM3G5Kr1SOlCbuThp/PgKOFh5yJcvGdGjCiP/sM
pmHvZIDvu5+XtaJR1PsvBIlygd3iqMjQDB2O09+3TybkJ3vmLIyFlBznOaDrI58+
tmhcxBkl1Bkxi90fCdun0WsV5BIQVkikkLoQfObpYgPe54plFGE0BZQX9t7vZskh
rDlHowHBAxxFYYNv4i3xt7MT8pxHGqnsTRvSrgSoykomW0wKq7gEVImaEUVdlyO9
X5+XdhvztESc+VdFGdgArWMhGLfkVhPrR+gjInY3pobiHMrJ3QW9f3pnxBw+ILqo
byxB8ef6yZR+KjLRYN2o+/a6Nc2Tgt4xW2X6vCUsW9FqClY5u36Agb10EdeQ7I4L
T87KIE/XyO4AaJL5aJRH9c7zSqzIeQcO/lg7C0olTjXGX7e9aL7Xe+OvSz2MQo/o
vlCGPo+JSEbXIBf54/SkQ4m6yT5gtyYvv28n7mB8zxgjDb5NpkVxmtsMmewv3FMd
jLGgpDNwKpBXLz0bIHgZdcJ6C+AYs2Gn9b6tzAZxk8cJsrdURm214mm04o32myen
wPcNVy37Lficim4yly5s3kvmA0aQr8s8Q1X+HRcjeD0lsfALNLc9hJWgmeNESpKQ
fwPLZ/Ns8iuDd0bf76dSDduMb3dcIMZ4mP7xrQWJ1xZErqgrSLpu8uByn3EXwYC7
latQF4fRdkYF4dsFWZRuAr4W/6bRLqcI+/AZi/mRU6wO8gPREsLOQsSdbhXFmwBy
l0ButlNDyAyUFCtrsCTUAeulCn8yd3B//1lgwpAeZiP8xZfHbS3SIbaBVVdpZoKp
NrYMftOtf0cmXxLJuwzSjFbTsGsbxV60rAK9KELGPFxCZ0r1NznZYdddU5Im3VOi
iQ+fTgG6MoTpgBDsep2b45C/+3I2RpRF0CI1dgL2loVdiMkvbwI17wlNM23QkLB1
/gPR8AsUdXzHQz8pebOUORgAfpZHGlOIdMmzV6+zzPZnk7aK751nVgKtx2nCfmJd
RaRWvzcj9RST5xybPxk8zpV5aoJa2dDd5QWc3AqTqJU2jVjl6U90dOTmh8t8i/AA
/CCNSaAAIYXwQbxPhReZS5IqXZx8Yx1avp8StiP+sHJVUf7yyqTpMcN1XDTgzmD5
zFF/WXwT3J5JsuSLCqBMrodqhqj0Xe/As+e/s1sWcV6wFdGpm5oyEB3aUFUZjdxw
OdnLhQzOyAI/QQQAhcoHfq7GmpxEiFtn5esD5t8wdgm4W5kdmln7vZdfA3vdUIQx
SjdgcyeosDc7OJ6B6qQPsQMa40DMzouMDuVPLF6x3YyGtCEkDIzqV+hQxej0iVe2
5SEbgFHWI3Rc9bAQcPDTVJ3kWp6eMb/wNkvjqJ4j3HI7uqdrqF3CRyzRe94MfKe8
SobbB2+UO9w+URPiiRUWfQou7xH2bxwbYDZHulyoYc6Y1WVafTiWyZTbN+5+97qA
ZYJaOjIEC3APIDuoH3dM71Zi+KyxqxyGHPQ7MAQ/NlwjjPTdUA12QXsfVkofV1Sd
Wkp7UbF2ITB24FRfzK3DSc+GXNUmSqXavLxZU3pMPi4uPkrzmW7kFtmiOBW/b6Bf
6y5wnfBzZunE/PkT2dpBTb7WwhQmFLzgrfQFFsQJc5fDortyl8nib7s+WGvtJFp5
bSHGXPmsy0dd1tZCjxY3qQl1ZQyvoWwmOGpMiYWc91N/RS+80ZDd+ZkdbBA2lpq/
UJ4720xkUo1V+RPVVL18LcPPa7Xy1+TY6YkhdWL7YuZMnbTrSQcX5/Wjt2m9dLbn
BTsusQtO0vxKpy99QRHqT4ULB6QsxD1KdQVcmbS4lYC5oSYVyH+wZBrUQ2KKoWPz
tiXT9mKoNbXy+QKmV98zl1hzhKRjp6AYisWqrfurFgz1blh6dpGIHT2DefotspOZ
ZJ0LoHaeu+ZWni0oFWH6du50S9dC4DhCruA/olYVRlJ74TL+KlPeu6TLr3Uv0EUG
doXdhZrSV2sjuoCzkH0GdvCWvW2k30oivKEQSLu7+dnKevw03auNmJEGZV+48JnK
STIX5YaD/kJWplidzbpXJrIvXR1pMMofSw2YvAr3HKqvW4qbSHSzCAz+5NgCbo5o
yCMmJASIMtXN1SUDHU2OzcXiUyP+GYS49y+HngKJboBqAIYo4vYEDpLqeL4S2WfR
ieRwwYU2REYXvSeI8iQOqdsJ8P1hhqFOr3R41FqjiHNrx6yC6oJiIMfjTDqu4e5m
OvQl9gDDQkNSaxwoGr8j6ohsp3nlUTH8P6nkfkaymVwbP1u1xoHZmvG7igdFCRGp
aaoE10TKGA4Vj9Ao3cJyyEluYaeMeAwFnVUen87K3hSb6jL1aHF9F05hVHepFfmL
mydlqkgRNKq+uvyl2LpJMiVmrG4WSyvotuznT73RLJUoReZqJViXimxMCzOsOCbS
ed+/z8Jf287mN755hmoXjN3J1KO9DfTdjZHBb0UsmWjzjlgKRhI5tVjF7J2DopmC
UzmOEpuxzoYcCyfhwLGSKxE21MLXwrMAM+cS1G+DX/qcBNHcppZnivjXw8Kw4i01
DzzvUXWJCYqZaXGcljiPPiSYE2Kk2Oa3eBp2qCtqqH5tczT3ngyh/TTIa7ATKQUC
d6Tp+MR2X00ACSLSThS2UK1TuKbdH56LGrK/Huvu/PxS/vDf07QMpcSw4B9PopQR
V7lxGq6zbnwUMVFfIBsGJ8o5Oeg9yaSrlfBH1/eySkmyFWSIquhAakjyrotlABNY
DQvYIyOK0MqMm5GXXRzN730emJAZeEUp9mYpqSYULvYwHCV/QmPYA57rTCcJLrHm
OJaB7hvUAeXa1v1s5rmots3Azen1dGXcqCY3iXVxZRx9ie2QCbDLCmV11BuBg69f
S09rqVl/MxWrOhBrUgGyTENDEaoNEks2n7qFOxG/o8OvVEd5TGpx8yODeaM7F+Iz
aqi4+XZmCTNvSevHGeSwRkTa4nKr2VXssBbNIzVb60k/cPZamA6xNhR1eEbx0Bx/
xkRViv2gl54bmZzYijy4ErATj4w8iZtrj9l0+JAeTFrjTS+usfHbEJ5Ht5b9DI8R
1jAYxAeSGPcsVDu46sdtTUjjmAjMDAzcf9NTdLkJzRzXs0uA4D9Baeo/qc77ArWL
FjRBbK/RdhY+8sCPRAP7ynZdlAQh6+Koj9iOydL/Q3JMDbQg8+bg3oLPE9iaJC2h
8P3dNKMPZJznqSc9aPldY7jGghr7Vq5N438l8EFeAKba1UgSwso1jiUfRhd463hl
Egu7acPlhmkfHUPb3DHZvYE57q8RyD5sixV5jSeQs4eSu7S5bL22Qx3k/15oyHjZ
THXqFW+2pdf2tPfdbY4c5R4JziOMJOBgaO9TRAQdJitZWt6C3v/nV/n93nGHSaxo
jv8M4JGL+0l2cVfFAC7sjSlKZmnXfCfABWyemqbW9w0pxzIFckZVpGH8Z9koQCSP
ekOTiwcFZtrR3mh6Pn6u0zDNw/0tmJr3H5DeDXjwCZp2/GcEHLq/Y9LdHOcv2sIU
YxsjKK70dwGyZARNl2v/ieiXBdKVss8RONOIOrWwUqRsd3EfwpKOerE/0OTZ6pmK
zG1q3fVAvAhmlTTdOBtkQ6wBdvFQ+WWNEsm5JDSegn7lLaAP/2y0+cZHKL72mLZl
TP4r10f+6LZJFMTE/cK0119Qx6BJXJZqbi87ux3qOB6uBkDkkkyqn3hgz7OOFG7z
w8oQ4jUbL/MylddnjKrxQIs0xFRusWXuOkWQwfiBo1PZA9cZn9luumh2qQT/6BSa
k/cKQgRbj7Y7d91JC/o27dJ+4XtBmuVhno5uJD0SGZE6Xo8YMhiKKAoce8AqC9g9
RVAhoIqurkgQTJs9rELUPp37Rvg40OuCxxyD5hHqm0q+YQjCFJ1zpFZOu/v78QKm
sDNF5ClssnP62j83TeDOZR+ITcOgO62jYo1onN+EErEIc4YXHAsGsLANB5WNnOWQ
guuS3VSJfUlOhEvTblW3mW6Mi88AxFP0+qAopG8x9M/WFFrbO1KZcS/XffclaecI
jO7ASIpvYLxQNvTirrJvHFQ1i86/ugyuE9lrS659JRE2qnOmzX9xowAiL1pWkSFS
MP5+ETnb5sxgw49C8CJdQZIWm25YHMLWjYiBTQLWgDatodQEJHlJaSc5qmZKNYqZ
FcThCgokGhWczwY009XAwLAlamJhvG/a0UZaSqvdEuCmXZQu1YIk/agG1bULcmbA
uWh6Ll+FUgt+1atgUsLuninXB4i8pa20HTcTFbiLacrKURpxlYrzaTrPKzHhWj2l
fnKuikwvk+sLExwA1+hz1HvXAmYViH+D92kx9+tl/qMhb8rct6vHdH5J3g7JEHw+
tMKhb74645gTu2YZrSYqUhU1CDSDu1YxHOLdvnPRdG75OyHsp1z7Qk+lUY6wnxvY
OJKAS/GNFTDteFEFq0JwfaluJbp5rVyyyFTQeHAlD4jUVN04cIXRctuvMt0Xr2TY
UG1RlBA5thLsGmmVyW4AdXw9+9JL08kiyMO0BNF/XUZsElb7sArQCBxhxC0F90Rn
DeY2NMGpru5nQaKo3RL9SGXDrXRVzaIUeugQgBUViK2OKflwxS23TLAcJJIELkVY
Tp7YtPWKFZFS7j31+g5necwA3C83btB8nN4X2/Hokkr34Kj5u6owfIgoobPxnMCw
2pMz93/72oDOjrRiRB2ZgHxwWeCrpLWfrT3kh+S4enC9CMTqv7c4dt/VHZidH5bR
5FusThXHh3MAEJK9G+CMyku2kGIQQ0Oj8nO8VR2sDFBbLQk/Cno3A4OFYgoI/egE
ipV4BJo1BBZxI4pBk1jJljRmQ1bfGIMvm25da0P6tLB6R6jLshZMxkNsi2xcsxzZ
VOFIk6HSi27yjQI0XM7xYdmSHj4hK9eqFH3j2NuZB5J+v12y58TxUBwZ+27ONKGk
BTldzA3fnIECLj9TAFgg172XP2mBvCI3PXGcPb61elIH1ibn+tDWp3tHk87Nm2ph
oMVOSRqe8cQXQw6c5UdxMXQgu1ueGLRhbvHMzIIVw8pz6QmnohXZnWh2APCm7NC0
qKBiCnTgABVoY8n9h14+7NgW28/a6AZYu8capFdJJ5UeNdQOsX635hp2JqSeR++X
lPgKgV6qZDhE7fIexUh5XcN8wFZC7ZFIpamVTODTK0Oe3r0PRrWApNhFx0RiCLNS
RqbaA99teTHmJWOwErHuXl/XbJr8BF/4FUFfwR+m8+K4JXJzRQNKcY0wr3mCCJb0
cVJiWyhZPFPTfZ9yN+2Rutmzz4/eAYqddr/prYWamNVBxS0lnOq9Ci7AxZt++bXC
X9ycAPvCh3B/SuPDDJHivcAFrP6BICR4I4SGlzNkW8k8qs/HdEfz1uAM60v2vuYb
aQ9+pnhGlr1IvfZBqjbADyeOpH5vO7KPU1hPmFTYsW8CjdfzPWSS59F1E4QS1m0o
/sM9OMf5fmzfJ6wvNkmt6c2yE4Lx01pzRZg1xgfLo39V2Owwt1fe+laaLrJPnZfR
LZrRa6aRYl7JmMzWuY1awIapArSQAhkc40uOxmvxLwCidEXmE63vzW0y+uxLTkZD
QmtsgT9WcCNBpNoR4wu+q8OzVB4J5SdTtQuWb2ehAkzlQAffme/fUslDX2o8IC5+
Vkb536OqhpzSxtemmIOZG0U8U7yehvyghhIFcxj13XV/vQWGDrViFqEKAwAlwMkm
6wTn5VcIRGHS1PgCkjECOQg0BkZeWgV4Zdn9KL3B2mcMJMoKfUk4HGfqTEMjd8P0
Z6dzHD0vuJYNFuQ0bikyVoFpC89hW2aliixx1AFzdubHziE0PLX+gRAXguViiBLc
D6LLN1CMD0z7+uPXRnCp1xUoSI4YeXTDyoa9jciu2zJHiTgarrer51Q/paKm/Yb+
cnaNILGw5Ya/DjTG8PP4IT9xfO3Uj00UPS++9e6/oBpF8MHHsY8Fd6EkHTVPrPuW
LOUNjw0TLRY6DewgzfeckSfEGXYAstn3d7WcVu4+YRuxx2Gpl0ZLCgaF4hIAxe0g
Hvt7MyT4bieUbV1iTE67MbjmwNEWBZkOGY7nW0bc5piWwX5wehIeOdfANPwH1AFH
fvqH7pI7+qoUqo7u54hTpfQVGZIEbzUPZYLoMT4x/qz8guNBX82QrClG2Dicq3Cy
FPnkHkxR7hnfOSFdrGzZ4NsbrLCzkEQPt13wu/XhFdFd7K1gnkPYiIVGpbpeIfFe
M9/trWDzdDcFXIMuvLYBEOfXAoigM6rZz3rF7MMed+FTQN81O5Ttzx3RSMKEZoS5
UdHA7a3MWa4v6e/sh1NwCcxWNUMm4stCQ2vGtZaptCPR6QAznha0XEiN3OONY4BL
P0R1qKL/VpBwot7+37Q7Lugi3CiRVa1PFrc9GZag78KEfwGG7AkqeHKN4Y28oeWo
9wIlkeNYG05vgxDPyJzH+j0m409v8K6L/yFaAJytC0Nx2jOqfOnRTez/9spEdBvV
qD72lPx3ZKT7mWRhgRqzPNV6NTVBQuRAgRNUqdSjouyms01rQ68g/ZCAN/oweQHx
aGn2tslJiGnesPfq8FA7w9SrikkIeGX13SYrkYVdjaH19INqkAxYnOH467be09DW
yW8+wA6TO8GGtPlFougWsaSa+w8a5kC8wL3TO2H/RcybIptoiCTnqxC2qDVnwDkt
aGLEpZSIU/FfaUU+/rGjNztuEwiybQzVq88UgfvhJDgP5neS9EmlkH6S4CW6MvpN
6HhzJyPRhgxmaiunRe1kBj9+W8SSJCN1b8IWxUtmkLjlAmAoxWouGwqEL5TqZI+4
SAAlAVaaqLDMGratfGIMZcCXvglvql1qFy03Cs43VGXywDv4OwOE87ORFRXjGRh+
ckFYCyMht3GPoO6zDkYpSgewR51eoXuyrd7o57903ShZbrmwyQMPeoefO80mSGHC
RW62wFpT2G8ojBVyMHgpCEeGXQqh+dS3LYZJ0QP/GYln1lcL6WPZQujSUJSCHnNu
l+hpCaqEj8J4wOj6xuhWK+rCq7sRleywBFmHXypxoCbl4r/wTemwXmpipUfxHIFh
T8KBbz42U5hmrYS3rPS9tUvTnM3wTCORuzX2tQWx4My+SmKkTO8ndyBHHv6wpqdW
BXSv7y1A2CdXm5yqAK4AVmualdClLGZtyY51CLGJTIvhQm34cWN5uLJgYtukllbE
9yqANp1Q5+ySckVLzxns8tsfSbWQkpEirP/HT6JI/1G2PuRx4XbRxSQ8pE8BjKTK
iNKGDuZjc2isIHL8QZm+H6phwI3ALTQugZ6LszFKkeXIoMfC7uX3HEahxoP2NNYP
NgvLNnJGYN0bHP7xX6TTnyY7MWcR5pYdfDCSO7YwuCWHNtkKepknle0fNm+cnt5t
PlFBhpwrgnA8WMNpksEg04FsrEPdMHLgEYqfxfQCnxCXodIyd1nmwz0Aqhc0zCxY
jZHR5Cpl7U/KGd8c/I0p8q4bXWiNflREjVBO11SoDy8Lgkbp4H8pVpjM9bE8E4Mt
Va1dhh//9Bx5ExKVNNFtOJi9z5DTmviuTE3snXrWcKbTW1dZdBMrICDXJ5FDt7yZ
7TcUmrJT6jf3I0trEYEydfdjnYhCFW/kdOOefzetxecuRH5y5T0KQWmSD/aDcrc4
4Z6AL4191/DBR6TmvNL7B2p1Pf1zmFzaQBQIqxV4yfCZrzmUCLToR0EQjQwI5JBX
WxBjyfOqD3FvnJWAosqCEmpqidrU+MLZGcwO6f9PZSjZ3axDQjenoEZEwdok7cXS
d4SommNP1DIwLZPCUfjmoel8bWg+YVXYAddx6NAytTnPLqItUZivuvb5RWQjCAMD
Va/v6tuByhzhE+eOg4bsl3osjCISGhI3f8DOJ3ADRIVvw5jc4oNTkD6TPkTggnoi
25SA7k8qwF4EfEqmwfwRqfLwGHUZjm/6sxLmpeFumh63eNWJVBwDBboFF1Oj9yAl
erjVpzcuIb2cOcLpuE9FLJAKV/Qlbn9674VcqhNfUktHuZpZLyC9jnTHclmKZY0F
txJcNhOxOgnlzfeAiEUhbxUBOK2hVEQy+QfcQaHxweW57FU9A94qVmHieeSAQlio
MZA/+6nUsym9TO28hu6D13YLXgQBkJzx1Ujy8EStIRilqsyOW4UkEL3sBRxxAWIv
lg1cLzkEBUsdFUZWaazgemXdTmpX3tVdeK4eJUU2j882U790qg5wMIcwFeHPD+Mv
DPMh5JT/dEQLTNwOh4iAwNRDJZTwoo8nn6aUlDH91UQRiQ176TVz3nhAHGogtJ/q
tvqnbU2c8akax3oki2SUBXz8fDs8RzwBhfaV/MuDplL9xHTsjJzvQnfF/dKpcrYz
AZX7+W8yxZVXjFsJ7UDlHQ9lSTsNqpqrx3hxwU78oFWil81S8knblPr7Qj9jxYz3
h+i4gURJWzRmVDKgWr5l3gXJN0vUaks2Ymgo3tspm7GTfairafB57ITKOmACKydl
dKalnfDfX4R1ogLvtvv7Ggfx3h3u1oDxxFYSBBrY6op3YrCwUis83fbkpbKK/o0c
OpRhtg4/T0F6XW5hSNoOX2gleq8XbAEEm84X91HtUxiIwlKGJfHXv5UnoQPg+FTP
mjSHaHcXIJy80hi4O5WLtu9n39WlXvJScML4SNK8gWEjAaFzsoZTu+fg+wRfy4iT
uSj6qEV2Ui3NecDM0ivyQU6tJOtvMmbiPTayzUvZZS0vilUre+Zr+IsAe+RsyXKb
0KlLiFME5j39kx+rwdloF+mREOYPE7s69Vhgx6bnD8QZP3Kr+XJZIOo2CyVDxQoV
ZQMU4BjQq4jZeqf0VVWAIjxdWm3IUsA0bR9JTbOq1IfuMNMVnACIB/mdqAsbcd7Z
GEte7J9R5+O+lJKVsJMFK3NhCZMi4nfOG7y3fw3yCJ57kjTjE6oMuODobiS5iZT9
dfA5glO0nDdKlIwEq8gpL5JzZfk0W5wh8b8pgq+qYVfT4SAoPoznqpq00cYRkD61
4VAQh2bRJogtKfMZTN8sQdAcHIPZv7+ZWoV6lUE2d+Q+uQMCYNZ9IYmgBzQev+FC
QcPGxEsDDnMnzpw3FroMspazs5CHKV0LKgN5Lbgs663MmXp5ODQB4ZY/6/PQyaum
bMevGvOTBIkgD3OqWdm6llbUQ9hbpsg4JoOWvrqoUmpBv2QddWuBykSzl2FDje5S
qTfk2pHvsoEPc/hg7xfEHzEaQugBlFd8QPHW7DJAnP++6OTdwGihhhQFJcgl/v7g
6SRd/dlfi3H9YZsFSrLFLTtIwzCm6gHg/KZ8Uv6JdJzJZGl6UVtS6XCaNpbQKFu5
FC2cE1CYybuwlm/aJTJ+hm1EwWvughEACNVnsM9+hfmBKEiYw81rzQAEzqoauyg9
41f4lMRAweWRomC2mG5FKo0ZFS0S7xYogKKYpf49Xv/Z27BInHHybcoRVEnjtUMi
YVNd+t+ZJqO8HxOASHLL+FlHn4iNkakI/c2eJ31DchSZa/Z5K+c/t0UsroWgf7Le
I6F+OAEMwLMYcFN07PYwS2l2d+sfyTVOBxd3XjnOfT6wkTb+SUFAdFoWvbMdzL2/
MPLqN0BQmHXJmXZiWxfUummvaKtXl3B36qeUWyHraFRnS2FqF6UjD+fJh7ygTOLE
FG1Ck4MJQVmyJK0hvmyuOBMZFW1v6kNERbBwaP8sNr5s4m/z5s9MuRapgoeBj19g
tiB3hhSH3onS+MwTB6EnufIgBrsvZocoHBUDixSqPGD+4bma16Oa0nbgrmMRxJGd
/JXA3U1Js8ocXt6qdQqtND2e2GNHnG3zton6uNKXUbdlFynfiiBM1min2eBOQbpL
qfZ0s5cGu2aPqj012H97dW5FNLwdV30MFyiaBDU8U35CI2mCdwADvSD220y2UtYa
PYdYQXTXF1n2QmzZO+UgjmOWN2LHpbNdqRURJm8Huc1ARJhZjtu6FMVEEFZVqvZm
MkoS3jwx3+IadsWqM/BT36qAf9naaUWSqNa+62Mj2Mn2Xk9MQtCci5F+0Rofm3SA
EN/io9NrhRYEjs0Y7YKi7z8+7ZFrckdKJgo56t+eQVgnBK1X5viFSrjiezcxvLbL
zpUWgy7fDN1czZ6FlyXUDvhJ593sHvxm/yS0Cpt1I/hhwWEhy+EkqTrOB4nEXkgI
nhaIF4MKOy4musYZwhKFYrHNT+F4OZ0r1bgb7iBxi+D2Dx5twQjryW9j39wpB4gS
xEMjHpwpGFSaXW6nkaR/9e9Ly2iJDeZzQ9zV0pSdRBBaV0Uhk8wlGgONhNzYJaUb
XFWO8z5xM7oykR97pDBuQWXlP3NLPqJzac4Q4XDA0K50kyXCtbYtKBqiFvNsoCq9
TOPBA+nfNlo9ZF5J2Ob/xZ/EtXozFraFzTyFzzrLESz0vEMQ2FNe0zqSwiXVCOum
DUzNzsF4az7VGwiO2umyH7zdmKz658n98Utxovz8rDN9bH6AgFK2jyiTvvuH05VU
IT4JFBqOdGOAPxLpNY0yXi0BejX0S78cwPN8hajZO7gM/WsTlo/I+lCgTxOynkZ9
jvBzZD7tJW9f10XX3x2Rda0slbL+ErYw3bJPe5DmpTN5IISA+oVspdps7VzND0+R
7KGm/ebx5oQvBpBoe77jaMUFlYk8YEMnUJy0wNNxIhxhCeq1Pbz6VyquFy2iqdNc
L7ANOldZThH4U7Rx/DQvKxZAibpVQaHys24lwk1Ue8H3A1W+eBl8Ancw2nd+DI1G
zxICg3WX7Os1BvTVCl+RH+ijV4Qa9Ccwta+cvRFvdcVtDg3K9Q1nq8u/HAZcKm2w
lWp/zdWSZT9ATeSmHGvZXDb2jD5+9RS5V+tDI8qbDReS3VJqPazwVgQcGpe8S/My
MkAdu7nvpWf2NU8NaWKi7vvyC4om5zZ0aNzKg/iJs86qSF24cdKC6dM7lugz0ZWy
dffzFupwiNAPvIjLXOQTYKGtjrYtBZ1EClZnR659P/iEB+cD8YDdbaGboMuaDisI
YFvsFg3DFfrQPnvcAK7XSdAPKNxM4OPMXMUFNBoHA0g9LqjuzG6OmbHbN90Bx9Pj
AQwdM/Thg2CX6vT2mRqA+etyc7niKqjfct4D/YDNk2nSFVV1iXzHgDiE2e1CD9nD
nbXZVjTzrKr0UmKk2lBDMaJqM14JNQFB+5XJc78JqbYyJXlHoL2eUAt8zksIVsM3
wDsP6A4Sb6x5kEyPVOEk5NtykFMgaU09q5JcTUm2QoDjPxdTypeuBM2/+/ydLB0r
QPnny4WHs7aW0QXl962XIKGkjVk52NpHaSXOrA4aftkrU0feWMXsDdgarBtvsDSX
iQjspIBDqQmYukokQ7/VsIQCOlmW5bdUQ8AUL241By3YKw2N2JITAabp+lz1cpGk
NXvKwzRr+4IBKn9vX+68tP3/p8IK+5aQiC8T+BNs0SUVvShmr1w78BNQEEcEEI5+
wzi261cPViJYNDezAJ7rBsZQcIQWRXuENB6g2F2Y5UqpSBUp8Jc/a2VLc+kDQEpc
j50vqhMnYOzxLlStVuR/INxy+8xNrynNvXRgNB5WN1n6m32Uot0oVz4Yutc6+hlf
91XKbLIVeKS4ogZqXc3ebFKaxPpb/L5lvon0TOdqVCzXXyB8vz1mY1N4xHP17rc/
7UrWw5ODmBVPlCym6QIqERrbe7vNRughoDf+eRXsxr0MhUCrLhgjGhvfUt5oMbNw
3XBM2f9fyTUU4ePcJDeuNPPLLtQgMnLb66bVBAQUKYZ0ylLw+9DvvgOQj4ypu9oD
fIIahNv/ZuJpMb5zxZNSUgtEiYZQhyKMnT/ipvpZ5LOhhjPIyOSGfwjtVhW3M6Yj
j57US2Wt/U4Mh5OlBrtFp0RQXF2p0X3T5DNuJZSa2mSxTEwIiNMyXYQ74ZLZRnpN
3FTUaXIP5WFScKvs+TGDNqsMD0xPvyFtizW6BRx/spTq5pxwXUiqdYcmdakG5Qz7
tMM/oGtf1Dyq0nf0Y7/8lashJJ2xSWxZb8FXu0Ry563zHLhe6/UAdeOhoLVlG0/Q
2hLbOH6lsPZ+ufnMyURD+Lyo9P+/7PUyABCi3GD7aPt/4N8rY2iZwBpma/UGjUiS
2sjE/6N2EavU8w9hJryT7fixJT/BiFCT99pf/0ckfAhG0G0Uxl2DVZyYIN4LvvIe
diGPt6IFJs7p65lezdBbnTE9G96ocw+hfBOYgWetKK+A83f8zuf8mYooxiMusHBC
vNP5uOU/rIyICnSwDZ75z07EjzP2UMnj6W70PHCWMdy1Wajg/Gh0jhUvFTRqurvC
kVxR8uI1wU8i1JJDPK6a4WrJ6XKa1Ob28ElXoSJaA7OgQcgiMKiyhaG5v/yInp8P
VshGY3YZWrEhywb0dyF1s61IxisWide6t+B+/GeBjKc3bsVWNNoURodqFLUlOSf2
ptRXh5+5vZl9dkflvTTEZQ3Xr5N3B5dYMuisL8n2s/UyCtNOZtjj11jJT9gWJZbJ
AEelAtnidw8l5R6OKtmBuf4P44wIff5rG/mWRi9iTdC8CyCfA7mamQ3NAAnCoP2o
q/Q0U057BiU4+gXK2qu5dsYXus6pF5JxEmoq1Yb0ig/mX03mMpu/gPHuJHCWUim8
vn2ZtuJ/4Ewxdlont5Qz7kvac7/HIen3MwZCxKGrmvsFbwGRPnsjwMrkqctCQ6oz
Q5OsdQWBQtnFGO/GpfHjFZZFyoGEEUotbbqk/4pAp/Qy8Udm/JBEOQsi7yXahNrm
yPRLc82JISdOqAslGekPQbhvu7qDcWisjT45OKN/Cw2bnTKFC+USMnUs4WAulwEn
uTFYWEDvAAd/6Pvv9siWsfMccsDiKafbit+fF8Azn3oQ8ni/7ySTtMsw+rNNkQfV
VCq7FDaL4IWNQBDm9F5jIqyrJGZgF1DFQSwiu16s3GZXpvU3dYvmX+yWsyg/vENL
p9xxdJ6b9xcTLvXcNaxR2pFsJn/usFs+gQGEbU+v4v4LFiZjuRiEDcwEIkFLECWC
mJa/nwvPBGQDebbReQ3i8lCX6deIfeDw2YBoq3EZ/w5f6DouHylruvKivHkj3+UI
C6vJhPwd7jxlLMfhWQ+ciw9fbXAubYWAIWK1Fhl51UdOw3P1op3MBVuPh1XcHc34
M2lKAs+pMMkVTh+0ygzGj3kuMw53T7jZZUPHVdiEFsOYas93FpDnPYruhf27KhWx
JN45JvYwO6e4LCxzfagzJjl4gcsk5T0jLtQBwlICFQgI0+U/1bNElGO08+8UtE9x
9WmTqMqRPlTY0QbkAZOHaA5rId2pwFahgAAI0yAlT2iB/B9tIcnDsmXpojoRWuy3
l5jPeBjHK7lJo3T9UZ2YTLAMeGihLeY1dCaT51QsMBgh3tnSbBvdgAC7ITSgSCMz
x1bzxrLzDoKLD6fY+EtvP7Ij0JXmFsnjfzvFWMW+6zbzNlR7V2GqIfROVCbNrG3G
m3KhSqrROg7mh50lWsS/G/zsyOWSwzMWj8ePy/TWppotqWkpREwgeoEnk4S+TVbN
f2h+/Je0/AdLqoUqAYyiI7khdpfNJ1sLi3PSfpqL535tX0JhTz6MWNJoAH61EVqb
JhCDMLWH7juQ7/TxheK+lmIh3YI/BQvHU3hnMISQC+n+ZdkyUww9LELrpm3j+yE/
E3lrbArFG9lncoCLmuZ/E/LCgL6ynmTVgxmia4QgU9FccQz+1LjXRwQTgud/FyKZ
cgcxQdzoR7q5twp3kdi1TSq/Z/gIbcC0qDC/f+3tXJ0VcOR32shNFGeu+iIYXnsS
Y41FmFsdEG5EeOvt4parmhdu1pk4H+LrSbNZo/Mz/iN9g8zUrUAaNGKhjGY/gQ9B
0NsMMv1qOCe34IVX3p4pjUNmRiha8Dyv9CcOlTGcQ/zjCw40J/WQL+RULXZD47wq
m8KZ2GGNf/poYbLXX9L54ZsmWoCQKXtjK5dLuJ8TiY2/Eu5EhkTNGg/O1Q7yOEE6
8kDAxvvpq8Fr13ClBefWSMtw9hQG+WlzS/ZuD3CdvxqJUWIarGt6OqoJW9AKicsW
mPbqAC62r6Gp/JmY9FJHaLUX04EG1NKsh3wllJNtLgicjTrgNCSqQqw2oDhiL65D
RcVrjO1Wa8/cbPuHbyWXaWo5WE9hIf199geml9ugqnmU0PE5V+mUaXHGIJ8/YzWO
wZs+CIlYAWBRa17JngEKfPJSJuTPWUTF11m8EMhZc+XX1RyI6lWarRG/XSWbz1Nc
VYlvHAz0t5F1p6BhSbzLTT5X2tM794j5icU+VDACBKdgtmWj5sVlQMz2TtuarFPL
Q0VAZWICy1vdGNw7MAI4+4KSxbb2itXaLf0WLhEia9AKYBx1XWktD8i+cvLnIDJ0
CF+5UQavWgG/KCNREqmJ89Muj3+WGHfxmWxOiMoHU5dUlF/xwC/WUun1aEYCVKmy
tQvbITZuHFKfBYch5NTrdyF8Tg4ZhKkANvcMvhUc4BWHrNDYfMO5Se7aT33XR7pb
PgOT8H085GLC8Y7Zi+dDSlf1iwJCe1glJ2R8SBiowq56JQYDRm/GzhTQ+9t+3yFG
38q34T+nLUYXfgZE6lU/108MP+AL2JKQEn9Zqc+AT5cyGy1neum6lPl2N7Ugv5uX
l/92gRBktdJEpGDMX4tLoWMio6BBqbDnQ5pkRrEjoYdKPLI5DHV4168j7kqoqJg/
HJPeaaF5cQIufl9PYm9fRDTH4/sg6Q+q023xEL8pFajHQMQzwL31Ph8A0rlAhRqR
en3/ZIAlTfLzpNK7wxt1/DqKTP2GsrY2/3+lZ9bQZPCewwW0RrjufJC2T6pqtImw
2hVE3c8+uPKzui9bkKLBj/ZoCpaggM8+3WU8YY64hTDX9ya13ufBaNO5BL8VNfuS
wM+gnpqmZ4l9YO0vVY8Euu8epiVbU7eCkPUQZNKU+Yo2spLIMuLPJVomPUueAxa4
9M+1pvq3iyuoEJ/a3OpJh8wYuktLMtDwrlPZHlB/4SE9VNyo7pcwS2Y1eJn974Ju
ecjhGiirr0VWFDY12XHiloy7EDGVAz/h8/fN5q2C412y4Gl3f3p5cAeLVEDKuFVU
karfRInUfYlV8TQKj8LCjvp35DAYmsXPT5WpJ9z+4AnsYrOek4KeOclCIlMK6zYq
MEGkY6bNpjpQfVrZ2R2nQnSBPa252qWtEcrkmqpz3aBoHk2gpSOVB1bL7WvqZ7sR
1S90/yHQbIEUAaKISkQ9a/czgygUJn0sqA2oeItoKz/lOL9dkzX5Y4MhshI6Upqy
I2lR4FRDvgl8E6mvtyLP47CrYucf/04sPuhZB+pWrotDU0bG43R1mmOya83zVL7z
KZhwWFfWp26YGmJjxtJ6KABWM+aAGSLXGVEuu191Rx94SfFO6sAGSBvH32vA/aQk
YUpUC7nYDpB+gOBVDUlgiB4Z+3sna4DJl/B1SqyXI5P88VmjoHRIXt/8DH/iEaF9
y47g+Kej7XEmR0muAbqcpxoXhJse+SOJX6vPg3Nj2Xs+J5BA5XMOrfw2QSK2Um/Q
Xi44zua8UEDq9OKrjv3gVpUsK8itt51IAufCxPInmu3Kyn2IoG7LaA4IZshCLOHv
Z0PVhVbTFYgpFNYP1aSzcCi3lnB3APJpttAh7qMM88UTgWiHGbCl+aObbVeI9qkK
BbuhZOBES3vVry05ZCUr5Wh5/681+uTwV4Aq7fXZMJ/M0O46q/3hrN7RoEMMBMW4
q9+iWMXbMllAF1gh5YTzvrD32CwfXRqMmB5+nbdNs9FspWpfuyDb6+WdfBLzCnnr
ELouMm/2Z8DwdxHHtqy4a5GdzPFCnh5KEn9rDeYEFQ1HLIkpE9ZEecIYo+wbbImo
vDYNGHlwmKJ5vXDPkUTEGgReI4fLL1uf4bTJCGKDURQJ+De7HtKGu+6rMU7btGo7
ECfvIlRj3S9cBsW3q7kWS34vPEA1rUx+VwmF6Y3zUyDZM4QDRxnhQ32HsZrNZY2d
Y8EmtEZa0AVb/0UIMPm2mVztzMDT/UHPlSkvCcz7gsbSqTBDuFcBt6RISgX0LHmA
cP/i6a7fobdiucHtwKLSHpRwN4RPuTMA8U9XnYCPL133to35081HQ4+F/aGAqQCr
RXV2eF8nayKIZ/mBhITHZAz7DaTBti0GvUCmHFNTdKi3L04UDDC2MGUTbfFfOpi3
Vu6uV0GvqUswuJKXXw6Jz+hkr+g9d6qRna4zuZxbjlSHKvrIJA3m38clMo5udv/A
ZBiU6glKQCm2WZzzyV/0x/DX6QmWWJZ3HBLAdUjF+AMpMjvUg5/O1ofJCpiIryop
5poe9M3AmYRbE3Bdq/mxdH5EyrYPCTJ+MBSjfUE44VhsuV35ryqN37gRTyzFs0R4
J2qkAFESMPFhtyz+12j3QQYVvxgApktcFodr0iDoiYZx0zUg98qvJQESOgpObkRi
QHSo4XGztYkKv7PSnNheThuGlVuxqLWzzRi58zZyueffcVdSAefM6gtXFFCWxDM3
99DU8TzA1yLZM5EXrs3qNQ43pVQpPw1l4iKIR3LQDc84hIpVJXbAckllYhi5A283
2nPzOLdvyKkkbou33IxrQTR3cdTc9biggGzbS92UNfOM3vKT070LC0GdNZZhA5XR
jDjQ475EprjGIJ09XWKJxscsERdx2TvaBuJ8PkDf71lsn81yr2rPqqEKxufftiHL
/znvN0TA4fvrnIoyfWVA8YFPmjEt7/5KnkV8RX9PxtD4RuRhT1p3daAqtN2CNw/U
s5lsr98hgp88ya6nU0ioptZJBRQGUjVEjKMmLNFeG+K/1XJPo8IdgPHrXsrl0cgG
dgY+9Eo2sjgXMmMOE5FVI9eiNm8zCa+9FSDVYBcBNYeqfonbX5EFYSnQJz8IqC1t
Z89o5o23U7EWvT6pCntkTQUFx6tcGgaju39pnNcghPiT16m0Jrnw6dxKcIMQUIai
MhLeLbI2SDkMqexemHEzmJSWdzrF0ebA7N9Z+WZcb/7oF4PQx4adausZgHJp0JnQ
fTDWhWgm248jew/dBiBo1KQD2b21O9e0jWdB6hMQXbcAHivy++8l7cVxODBdB5zh
mXM6BUnIt+LFDuxjx2Y2CLNumEdabWuglTmBa05I0jmT41qPpz36zE088rl9EPwe
+JQ/QYbMTFE4HjXrToUvjd/CqQ/LYvgJHYo27roGOy5bEqLATkyqgofDiEP9cZdM
mXed64wcW/tl89nx+T1q8f40V7rdPDOuHckUvBeITTCLBFYn922/bcdrhRG0fxau
n9hzuVznFl899JLOdAKwAfuUUq3Mhy+me4pIuEJ8VBNi++HPCpcE/xMpQ/GOxnpq
j1tUYYJKnTEPsbl21zaqHhlEMkLVPRDADtG+cxeiXN27ryvbeMyY+qlA/8rcdrDV
u4Ps4TSvKQVaw14wB7DD8BNI9Be7XahZydkyO46ECLdXNaVK18FFsMNgw8DyncA6
60RTEyrWUGi0sMt+YJj2Q8z2NuRU+XjpIzk+F6d7o2icvS+jKKWQXsSEkn3itwG4
y+see6VaaLXSq6s7Kng+5HAEKzICuQtiEdyk/m1OA/3U8sOG+FbaUiheZqVWEOtQ
qWewh8UW3hr9qxHZgcQAXIzMLy8uK+77WD2AjKw6vbzMq+J1C4Mlx8kB3QCte+wQ
ZP14AuZFVz5vKAqZQ0d/x7bchhoDLCJi25eO3GoKIWcmvBH+S1ZVM0j5SANgQ971
eRjGd83SUkmr7fcKLrcNhzA0XqnrFcZg0OkMmToVrTLIGQvP/wFgGLsOSfUNNDAi
m/iJpvkenmm9v93bWY2NaPBL0qnUhoBOzSkITjTjE36xpv0TsDq5YdYQK0CdHar4
Do92/4M17KxnLPDUWJIIJhE+wzi61YU4/qwwOrbVTgeLZL7aVZ7GB9OYCNq4JbND
eNQYZZzzIoXiAzsyo6Tpc9s85PwlvzNttf3IwJXjksMu/Mw5zhUH76d0rEMcSwAp
/faIc6hdj7jtX6glucfpoz+wsyXamnbjrjbVQe2TMYh5vAaJyrNRDBBy4m4rd+wN
OTJrwpDesyXTkoh+PBSMVeCHnz/GDgXawzldwHmqbNcJb9vsbkYtgcHBobS5qj/V
YUZG7SSviQ2S/KAPD6WxzKta9a0COgRN1ZsLhH1nCdMK6jee2HpyIy7ujWrkxkao
4qPAtXrtzA4I5pYlEoczwZYzBjHSdVsjYx1yWl7r9IU5HmaMHlzSuVHvSa16jWG8
9W9FpphiAvk1CO6g0yUJqGA/CGxitg1FhbqW3p5ZqC4c+a0xZie5SZklL6a7mlNx
J+E6m+7Sjg0lAioqWVJDQM5M29gVp480MSTH/MmrmHQMm14GA1ZoyaA5toxZkNcz
rYjajjUgqXO+JUecGixTADSQgIMqV2rJx/rQXT7UpbVSKXxeSMbaM02mZ4QqSXZv
tmYL0eFKcFcnm6EcYDpScHzzsegP0iUZoVqSWraKxRiAepojHiQUkFPs7Jt3vD9u
u0CVAgsl2DezaoWqh4k1AqMRpVT4rMXMeNbQc71FiLiN7SA95iGh0OSgkNX5UFU1
blmudE1C90MMGopryiBOoeXwDbsaS9dScmPWMSoVCquLGqYuzvh4ukxf46RBAfTb
7HR1SZKRzAFUDd0RnoflmdySxUdzjIgMJeP5D/CUj/2oFcrVXiHRHz+jFHp20dBB
1pfqSD1Qz8IYE7wX9oIK64AP7odpVw9AdC03yP29Fw3qhQPSDOyX1PPMZsVZydpD
R6XIPWtcm1XgYvKBqeS+FK+qSVhuQh67/G9LoNfrgh8uh+7pfVfCS7oartUQhk2N
NO8G7omKrpIVUkn1yEhLtxXjZIL2lKsy4XcsUHWvT5DRROdfB20BNiQJlNo81KDr
0rNzs+O+KlsiRAaZUPeznqcfS5uQiiFYMMFmd7eGApn2Mqe9ZdCsNI1lPwoSdN2i
/v6TRPEj5jUqZGlUS/dICwqQQF1NVj0Rnp4QZU89i/7bKM53lmwYftvlXlk3xiMR
86rNyCBfWVao4XIahIXuG4yti7y0OFTrWYIX/IlkU4VOwO3jVHlVWXL/mOLihVPK
4SHNA74wuznhOGH1Kf8DSMSaYHtGO02n1lCLNASk6h7lVjI0RSLlfIgeqmYDAGQg
KkYp8y8m4RFOCtSIxh82caS2dmv9qTO/ehfCNI7xmtf8bCWxGF5DyN8Hibxbi0ud
zwaA+zqrrWGIMog1KHM5Vy9HtcCq/QUYBKy/C/6s85kZZsl7Vidt009OC6ym+3PV
+Kl28n7wHNhMkqGPUlvD/0/M2hWiypyA8Dd6w19d24XcipO4pmE9HvZgIudqh+pw
2NUH+7ihOulb26qDa7l6F8QmCaw421SFLjXE0bkwM9E89nfXgXNlV5msEje1sfiW
O5cnMdRzU7rJhbZ8z/bp7BOq6fPbbBAlaoDlDjXw7W9K6JSpcUXDwKMSM9dXLf7r
dzFO6dmvQwIqombdiE1vXMy3r1nK8AG4oKhUNgo7nRC9LT6Ye7VHM+w4bCqRVvL9
iQ4aOVTzeXrAea4WaV9D7N6IgqcRocelT5bbuGWR7Kvx6mgjRVAFjOizUYyW2Fgy
jL9qYf7gD4TB6kCVADDTHkivTfcKJGhx7HhsYt4CHYiwpoxLQAfARC9Pie49Zupf
21X4BJjklZMLhGGmF5An4XNd7rBWl8fRet8VExsVvKl+YJFCv/8JvCUFl5oB1Aa2
Z7KUTWqMtGzGC8RKivoXREGAwxtYb2He3IS8nPMAm7T17qR5Fmhx2zh0wyPwSxEN
zoD1iK17TqNrqWsssOvGDzLM2COYquhH0ZoZ/R1rpPdn4eqOFSDkGLwAKK6AI2et
EIo4GTS9BipMzTkJUFj4+ILCSle+sa35bZfKAzgVI1iBGfqV+EHfOTP7FqIS5NfB
NqeHGqlwONbxN4z4EFiHKH8SGRN6WYx60O9G5cAazungiDooQFBolr/BuGkv0Wlk
SHIZdXf8EAlfZLTVFdjUu10UMbv2DTmxffIxIDDrQKEhFOOzyuedsrB0OxXpcdje
ViTTwO9K4M/b+eRMQzpgCcOwAiN8fAVfuAjoj0sQqRCvDbeel223khSVIK2F+MSf
TkOFezKkx7t3Nh1JgS+nDJ+xjgdfBdY+y6D/ArwUiC9MGYRczAr8legrTMZ9aKPF
GfjKCZtQnfOC6QRV7jFZJfg65kooayrIVvX9vG+jJWsAMrwEpycP7+fPUJiuY43V
8Bj2XA5BNY1nuJE53/02/UIjPCzD6zvWdvNqzvmYbSey8qCYn166xHMcLUl35HgL
xkiEwW5UHxabQ99+JdQrbN6lVqfzNradZzepaLGx9Bc/SfcgDlm8ABAsJ13CAR/J
Sq5K8Av/uN4IUuLx1LS3ztIYcggjPGNVNnpy6T1cFJGjfECKmhJ9Gbm5wnpR30+/
k9qHLAliU7Ncr4Tb1vnR0ucUohoJ3ORGtBRCuGj+/QHykpHyg//mZr+uHyLxVHwJ
he0Xpl84w0G8hxolWUnyh0/pyyaQ7cynPE26JeoTUZE6IbpMAgFbBr4rbOAMcl0r
h16N1dg6nK0sA8x3kJaUCjCgdVTd3hWTm+9VXcKLj0QC4r3BZKH6ML+KfyRl9Gbo
aQrw+Fwy+nESko8NbDfu5s8aGoQV6I7BWZQTejHLaWl+h0/jIrwDZm3FuoA+HYmG
MdU5IenR4fvuhiOt9HSEto7UKiYNF14HpEJIj0LoiIJNHiAr5ur4yot3soTtkLMz
EJjlrVjEE52XgXSLG6leYKUFkzT6P8bjAsD4GCfZOVDHEtP4xSA2qqw3t8CLtxRk
c7FRl/nqvpfNhczcMGlYgvOWX2z9mmqzOZbizoZI6qQjhLHEdCASeVCVuGhCYMPg
yrxz91T8n90JPISVnY9AsoYn3+Gd6StyELcR/dbqq2h5u2a0iq+OQEAIxsTTr6DR
ELA5scf6ntiVQBKnFLlNMbLZvQVkmRu0oFZKBUlWVM6FrqhuFxXpN8w99JMtrsUi
UMSH7VZ0JmSAf5qt8auAPgZVlqEPKm86M9qUKH6H/IKDpb+SpDroSeLQb5sw6sn5
NWsnE/FbvslM2um5aMyz3VdQhzCQ04qlLjP4DbOkLOR1wpEg4aBr8jxA+3eC4whc
K5fxJpiNk6RjWgqCzjollX+OMenkMlCsH2noC7n0uXiPrEMp7GFyIovw/xlQd+UH
CnNAEFTBuG3HhHNLesaC0p5agkS1OWUk95/H4C4S32i4RuAR8EI//J+jeXJljQTK
nKKxVHqQZ2eyhTmR46LyIfVXmQJ4I7AXzVDYtjX9tCC9vUbt2xAiA6+l7DOIrfEh
MRMGDcwCdf1jRWp9GeTxjbLcNU17cl1P1DhAO4f/VC8OwMsm+JMbauasIXNMwSiH
Qz1C3k0rC+rxxRod14lZPM1+FDfka+L3/uiprhVKnUV9bQAImhve5/LEYkbQgD2R
vE1Uyw+MWzDgobXcyOLbU4VrIRMzz0XOzoBIHGsvWUYpaAEpu/wbEp41wktIFPG6
o+WfwCPnWZAPY1j82I2EehbiVXC59kYNKALy0fqXilQncq6LjNfi18oUQ9NmR8Ps
2KGT072ts6AHYLnJdbNyN46w/FoiDVWBYssZBnlHV5K7LuUwMB/Wjgr4Nh5vsDiN
V+Qdu2+QRSA2sgFVFbvBWsVo+QyVDkHTxUAE4WvgY/ilt/0gMUiVH6p/DrQbRDMU
PYX9OkapAZcFDDq2BtasfzQl3AkmQp6UT4svZhcLugZMX7ULzW8wK/ODPywsibE4
kdZGWU9iT3s6tE3OoSQcGezJ1egM+sABcSe1FQ9PGopcMCHS1Zi2fnNSyEPurToT
20zpe+7qu/AeeI8UxolAckWB7nJ2wRCKWAXS6sTzshffVA1SoHquH316bHRum8qg
yGKr1CmpCluUqy0u6yWURIj5ecDSfJLsSIbkP5f3bEbpPte0zuYdXpJHk/Wskmvl
RhVlxnG16L/CYlHU30MQ3OVEm32bT2qjZMkbExnRkaWFz+QCJn6wsAM5BD0fZFXC
5TRT7kPYmhDO2qKfaPtp+31/th0I/F6RNScdF88FUoExmYDlhvk2NtRHTkfn2CHP
r5m33SvHOO2MXcvAAgAR7b/4ONgK7Cct6DiNgxXF8dSSX5r/FFViWMQAFK9penHL
IM86p/yNnjKFrFHChuAdYBZtyOaT6njBBMEYYE6PjQH9CXj4bhQd/YyvzHff5xGk
V3eB7w5ub+8QCzuN1OXdKOV7AldJWt+50RnsXa9qDYCa2dgcPTyGqVER+875k+vK
wC8fDzmapz2ycMucO8JlWaO058cO40RB25B9w0hp3tZs78LgZnxa/o5ISuWg7TOj
qLfuWeIZzoVg1FaR7IeJthv3bJ6AHiS5Bgyhvv3+ZWHLLnJ1F5MTPwyUxxOauFna
QHNBO1pczzWbArgh9tmzQKE45GpaulMNG3noQLnv8eBi6xOg+x4zA44COUo3nksP
1sjz1O2z2AYngFKY1aKCFwpOvOekagBxsRPugI3lL1eGjWABcur4FxhrqQ0afY8q
4hHfKX4lZCXIAAMDchn6yFmghWcXNuNrQav9NNfQvhx2HYBh2ddyT6+SGi9d3fR6
762MpsCIsBxzEW9QgpH6dUJo9gdxI9aTtL0by4XDx+y0aZJbDyx3kcYFnkiCUxlI
DcyzRWBWdo+j9bDjDj1p2pEoZ4WWcHIm5/rvDwVYz8K1CXSiucc8C38gjUN94HPJ
iFuedf1MiB4sfVGb3E4FNyOHfD8OzzCB6pT1zFFezcFHxN/FPp5iInwpQ85aXQEu
okxvT+fF1OP5QHlXVN0K4RNtvsgnEwIkN88ryosVttrGm1I/X81VgMXmAcPfNvNN
J1/EjzBTRQM2J1bv1g78bg+reXnxpG1mcLoH4yENJVGAGLAMLtQ/CxaFJhsL6GMP
rrmhiIk4kMBjygM5W1K3P6hMT8L9rKnvnZMnhJMt/UuLNZKUiYI032TiMoThdQ8p
vK2ntPsnS2qhzsDuamV66iZVnFOKJntVGO/b+z6cxWJ02bgHD3KA0kbPETTHigXN
D9V6wbrnEFyaXVaDRNo8i0VXDMJyAipqjg562McjHbkYL/I7is/rk+XBEHy9haBC
fNzvdEXq32xp4ofJOAfZ2kvtiEM4bCSkG0wBvXOSHBltfCWq2hU5O3X6PaIB0iPj
2AcnCc81UXWah6tHsn8MM/9xHDfIapJF0a9pIHfOKGwStkg/3+9SFNWcninVAsoY
R1krGTpkZELQlzxdig9zlS3GN7zmAnJ/pk1SqH6Xp85ofu9so0oTP2W6jkStgoVb
VxVrOF2u5ugifxd1Xk4U6tTyKxGXqzDUCYX25p8g4erD8ERogFzFMp3XilW6uPJd
hF/6+z+qKehrsky3Qj8y4BxGANTlkC7rAxpWrOL65V8EXfcfHBhbiM09j/IgdMJ2
CXn2h2MPbdx1ngp4QHy9UIwTx5kERuNPUTmKVlY9NUMfQlR0w9mO1PU5yynqqNWh
DuE99ujGkR5mVtqRT2e75YnZ/tL6WZKa2obgUIXxpkXWFIl5xlhxXyDX5L9Ugnns
TKYL7wq3y2rwxMr9mn2Il0lPqhpcfFDglY8x/cCG5394PP07IYBGHy1iarYX8vyi
GfKpOyps7dimtrpwE2SukhNpv/vBf4bq6BJrIsXqxOG+l3/RdAjwsnt52L5OB0z5
VlWMF7r4ANoP8wrMBigRihEFZpxQ9Ih9Akn4TdyAW2VK2Oho+ZGT4dhFsLhe2mJG
RVAzwbuPJlzIuT50dtbpuHjWlQOwVnV8Te5t+oqhBtkd+NsccZfiPVnSLtigi8hA
74wuEYuLZTnvj7PCbkl75nB4XVa/0BbqWY3QrtYKA+5fs4w9QX4aohwEIv09lBxW
cbGvE/XRAvTS3VMebA4OuEj64POFqMXZqM4fpW+Vrhe58YNUq41Ph6n/yu3w3+9k
uTq+kAWZc7vp0HvGNcs0G9HGELbxNonP8C0JUbvKe5zVD8xSZhO0AnQ1rb54XiZb
Uhdr1ccFbpGgK/4leWkDOpKTU0S+bB+ssddjYDDq5fa5CF2ESEZrVxAEna7jZaof
GY4H9UCMIbpeEpIMLagRJvmD9qlhC7CjgKht5XmXR0HxwZ+725eHIzBebI2Bd1bq
uPDzW+i2io1toNfkUvH3S4sjs/mlSl5/WfhdrEI1Cwlc2G5MXkYDv2cZVVMvKfge
yHZv1vkhRo0qmJ3LvsWK8czGqQVd07JoIOqoRggKve0ePY2wjB7b8TbAut5+QNxZ
O0P84hxCTIfjeMJ1bhgsXzdtQUq9P6DDd7xb4VOeqxsN0ZzcyjfVjsQ+ZG8OLOIp
X2F1ClTHB0oj7Zq8Jt6uoSFWn7ZOJ3joAP7XJJcWlWF2iNIE5NiHVD0E5nuTG6P1
DLQnPUbdbxBcozKb99dj033AIOAq7PyeMv41gjLOW9Diw9tnH/3YB81/Z7GW1jBG
nBeQlkwxT14VxNzXI3EHCeCehdkOwD54JhTnOagKyLAl3unLhEShPZx9oRFJmumB
4UEEMuifK3zhdg2BUxUTAFS7WW1GurCG86Lq3JmpzEhgZXfZGGa0wqeX1/o9GTSp
3Ag1wP6Tt37NywSkBoK/MBubdCafhf3etlvrOdfl6PvxBZd3eFS9d64gY6/uQVcK
tF868GzmGr59tGXdzGti9d5WANt/1AXhuFJGwTcymWa3TwK+mC80JrpBSZ/D3K/I
BCfk3zcz7Pvja7OK+VRnAczZ94tLQL5UXYPZSe02EHU9FzfHWqaDS+2J1V37yqQ7
Nw/EsXwtw9GxBpA3WMed1ndf8Csdb82UCBYrk+nv7tSUH1nqS1MwpGXnPWoo60lH
tTjgA+xyOZ+7/+ytClRTe4ZyKH2sZ4f7QUMDa+5R7fePRiIjQsbCXyASNoUTk6ly
AER0tAc9jzECLcCdcfdjwGVoOTXapwikJXLdcPdphvY/3QAt0afQnAcZZs/6Svnm
y1wJjTSw/kH8RG2PVVRvImW8LJPUIgPMvzx8OvmT1PJdjT3XAD8aK2gkoHV6odvj
6LaHdHP0GLoYeg9gza1uqudbWwMagYaa22xQmtmKjF/89a1KOAfu/lleh4agi+0u
EMQ74SCFZ6z/uyqgeDBGZxKRE6Ffg8BxKlspGsfQA/f9+L9xCgZRs4bShOPEEFNl
Nzd3bAxcAeyp6ODhbzzlJFSUVDQOD9kK35+oV/1rI9y29jhUmZ0B6mKo7ggVznrC
9PjZ4YDz+ZhbgBNiYyYaaWi1F40PFhHOxWys2Z59VNOUz4q9tLm/YflmNZIqkWQG
lyqMoQXQm9fEKDvt+BhwVcpWXSqL9gkSyB7mw1cwBVWaeSWA7TsecJChFA1OOdt/
lMjR5Wtq57VNmeYcFz2parL1vu/Anorj7gbE4S0ntsy1iQg/B2UGQCKDowuO8VQO
yAMSCsuDP+snRzLaQwE3L1KAdD8R9zgXBTJJVl2fAhw0ZIGMoSaNWCutossZRSzu
7YS44LTRQB7XlLtJ6itxf+FkoTYG04o/5UaRrv3maCmlSO1TWH3T3xhKsLeqH9c6
9jsWTqQ3cO0CpbLHQIFAm21OECwGFH7XJ/QsFe3Ji8NsWUmFSO9dUYLltTocXxrt
/PEaaE4iioppWwx65dAliOct8ns2WPmrbhMfyxpyxafeqB+d4vYD4aIk4pRMu7jF
qFPpqv+vM5mSEGYbUMcPuDnDJfvuBhzZUtSjq7ZutejIgKxm0AhY2QolWZ4O/FdS
0Cvh3qHqKL6SoFRbQHcqV6/hebqJNIm7bFHhX8x4jdS7RSiVyfyHxgoWKpTaSxwP
kiV3xBa6BNOz/tIbV2xB5hGxdAzAROUO8Hgyr2i+Hq8VUHnSXQfJLT3BE1b/zjar
wBguo8ENHP7fkAo2vpnm16XA1+Y3D43qUdU3Co7UOpeTeY0bGzbk/CwXtpVYt4Rc
MxJNdLxlJaaJBPFG1j2VssU26Rx8cpX3GjwvN+PW/PGrR47+Fkoktgk1iXhWzcH9
lFxv69Njn0xUlnn711HAAeSO+BYBoRPZTQ7+KH/tTfdqlDYO3EEqwCBJJ/QVtQrL
p36vakxNIR46vOqTFKrOp5/CVNx1eSraWQVxwOkd+V0AJeZacBtKZhCOTdNV58P5
9NIC8Trq8DmMvuIB0FS6BW/i+Lez0KWV0r5TAEOKegp8fd+JX5XF6Mf81oVXe2PG
1DpGcOQj0fG9aQFrYs/NUQojcabpvn4Ub5M5nPZZX5zlNPCbsSA+a5Inl6zBc8L0
vToinM5NHXLWkjDeg0itaGkfZrPinNZoflgSiwyDNSS2Xu2RVOYpJA307FXq9f+z
93kBldVNLJVvy6hSaJ9iREoiboc4noF4pgYHnkGroQJup4GQfzQ4Qe9Yh0l9c4nu
xsAJkEXu9nZ8trcOw9M0jFUp2vy7h4qmC6agLKfVxd435PGjFrIuVNUib1Ybh5Bh
7VWq+mU/XH1ELvZCilapkTqWDJNt7ewPrrY4xTIbm1hZJR+tHkPL0ChG5VKtA85S
4iPsGZ79v3NM+mX0BighMKbWc09GeRkWlqlY4e8GwcO/WfzF/EGEcfsBCkh3BEjz
ctFrCXwH05dJjLgilsKyanJasxCcTOd/u67RcX7nYLNrCt1Y0LXMAAA9wXoRJLps
RMAAyTx5vny9AKJ/V6t/BljRmE1cgcid0BoxBl7xOIY+hwhnFOvLj+o3tsSqdgA0
nxUEwFL38cteuqw+SsxF+m1bGRr5/aE9tXdaSV+Sy/okerWQweJGZj23H+SHl7V/
rCFK1ReNU7Uald88k3fkhGy/aAt47N1VpFruNvJlTHlAh+BYRNRO2Viakxvzb/YW
Zq9wffIzFsi/mwsECs1qEqhcc+HzoaYeaR27M2PS5osK1KREMGHKdLrPgYYfvrn4
tsu9JlN1CgJfLlNg970sX9vxOjiRXeo3zrE9xJuIoKMxG0yxHDhrl5E4rqxY/sBN
gCgdryARO4UXGXM8fCvW29/o1gRswjsuBz5FfopMshWH+wQ7D2yAQZul/1mr7nq4
A5zWOdL39pkdmJM8ovzv2Z2Z3g90RnoUUOk7kVdZ1tohz/P7R22a26Piw/H2uJeV
lTiAzNBPQ+zPbqqFrTUEwDerV8Kr3nVr+cxiQnYbh48pXlCcJYPoxj1FyDtPyj9J
5rKeYu50AR9VvZR3IRXWOdQbD+w+yAFJc5m54sBVPnHO2enaugTp7JQddXsRrTWB
NBAqK0+igwDq6MhQ8o0BG0EEwgrSlI5c5QiJmLabP7hS8vn/qnwQR7MS1NUtf84N
gq8I9ME+aDvLICAF5qhkil2Ak+pnSqAB0GzTL8NCvxcyf52iWMZcBgsNHyWpdzQT
Ph8uezXutitB7abejFsD+MZVCko7qPza+XfDEOZD/geu40HoGF+ZeafvYGcUWjrV
iJlMB6CSKLUB+6wFBCloFB7FU8xrXZJOqWj8aWa1VqKXGcya4akNw0Tc8YPALpf6
b+qWFRXCTnSuWzVnebIzomzu/FbZ25ZcBiBnu7jRXTBXowhB1iY4PcDZZEH/SUi3
pPtoyDjKKzZvpKP1uimDahXIWx2xMZhlnK1yyVYZkpyzRTBv3QwCqDZk3IboXGj/
egiozJhuihuovpiBRAF/+AtgseibQv+GZtwyKXagUkgxDtU9Vkkn/j9igFvy2DLB
76817ps8YNP6nMB7SlLo3kpQcfCKZDbue7ZjpqEoAJolLJsHNBYjfnqTGF4nQkVW
/fvQ+Ydix+vrmkIe7ayDXObN4VrfNqTaBTA/KjqnRDkKAqD+f0r3L9rMDGHNBi2P
nf/VnuvnWP7gf18iAy1oFGdNZ0U4y57aVqXq2yrwNboJ0ubjuHz/VxR2h9ACuXNg
lmnM4S7QQTEvKTbGSp/jpkvQH59ZpcxK0N9R72ZdYFfq2bIw2w8TUlq3koZScMen
2MZhX4vDs8+3caGFfgQmodbc8cfPpJk6OzXleGrhVG8qN/UBRoQWP8/WV8Z6SnAc
HKviK/01WgyLHH/bgOnkyWr/pRwrYU2j+EsBwrBZlOO8tYFKwDM7vlOqSEx0TSdD
HYTzHu+LgEyAm44vzuePH/3624ltcQ3rvRozQ/sKfN/T3xWFA1XYrdUeUTovrJMQ
llaZY40ZRDOQc1wui/6BgJ4afeA/WxfPo0RwuooXEqvthbhX6PGM7xHkF+UXcvnB
EdTiYVTaWxafi0S8fvfYvKwYNV5eJtdP8WqxWJmjG7kzuHUWgCYFujpUXHH3FC7X
dujUMhdnXy8SxdRLWOaX5irTwk/EqQlcLSblmN3iPMjLwiXMJDd0vGCFzWCjVeVn
zcnRxEgMKhMCmrhEog3LpDb5eCV0rtJU+lu7YF9rDq/4DhdLOTJCKROqq2hxuP75
0v7D6wM4ymK8nlroFAtQ72R60I5nOt2f8+t6uRLVppqzNOH2FlmhHJ2GbONNJB6n
3bjj4dlqWc3OvogsWcp8V0/v8lkrDnzDzVQSfjWUVjod1jTzimOX9iqgQLvHWtua
zVsuYjym8MfnB8aruPXWGoxT+OiYffWNfy06vBw9cQifUHJiLaQ35q9tmBKAAq2g
hW6HMZeCmGr4bFdy0LDF2fuWgSOE50qHF9wsCuRkyw1dRc2lwqihlZLMskCNSjqg
cACLry67WSREWvIC5OpuYBGjtRFAXMSa68cagT43NZsniWX9pYWZFQM5KxBsOZ1L
QeBpsmWQl1J/k71337HXZNH8/86ETv+U45UOAq5dwzJqphQM6XG9ulsqG6XO/8pp
McCFVs0k6INO2VUAIbwUsRKj9J9SPiofHxAnyyZ7tiTfa6GFupDZw1GY/R8rNjgy
ganseUY4hI8tjAxf1wHtaG46h08USm2dyLcl8VVF1No4lA6zWj5XqsDlbXkgYGXM
B6Jdqrhiw3DT81Yx0U2vv2Jic1jFKyc0edkq54lv21g/ap96Xw4jQEpK66ftsEBe
ZwgWPb/zd6fBpfLxqZHTKS1mG2EdDmWoALOSPujY9gP5dmFk9YRqmx8CsdS9p87X
cYkHXfyO0ESZNtxhC98jhz+DF8iqz554hnYHxm/cI+BPPCm4hpd8GJSbNNnWB5dg
78rXO34cy/ymUqGThKhBT6v8ectXwwBM3a8zFANquWQ6Zp0dWyBT3B0MuUqvMbRx
J/IhiIMUm2S7NO6TguNZIL7QYhOv9pkREug7f0FwNN8pOsaxVrhzidZQM0Xn4vG4
FM/nJpyNsyj4E9PgPqg1EL2m0QIdMRuGs2lVdn2tZyYmJoY45sesUeOd2V7iIMQ3
55jqZd5lLAkVYlPozJ6LZBZMjFKpX98S8d2qEn6sWeVjhRu3Eqvi8uod5tTXMljq
6gkg21DJzCsRktatP6J8vcOGaNh0N/Zkahm3qM9JZjScEawPAmFHkeIYlbkMtv3P
nKPSdfrTeb0nUwh8Nt/CzbLH8L0ONEDN5aGPuzyrhnr5yOTV/Cs4zmwRhh+82Kkc
hNSxsM7wAocSrc9TefQrF2hXHR1js/Xo8da2QOsjV7T6HUmpqhjEmCGaJHefbKf/
xu7W90nOSPrWgOv0A52t3WJ/+46o57KXkY3BqyaOfsD8aS7IAVeaWYlG1DRO1qMO
Zwjvgg8vdOGsKrNmA2gSjBWqQlW6i9mVYkS9X+Abp/4Bnrd+L0jKNN+C0doWRabS
QoCSOJpCAC8cVkq05/p1WLDouRSqy4AMkQTGh8s2s7XF6f3YAnHgcAsBy1dqde/+
uLCOMd2xAHxuT0aUpyH5xXdwSzDT1R8L4W4wEJTPV4Ncysm96rrPvPip9Jvg67ty
Dg23XCN4EF8cob5yavBJTIcrEaR/Q5LiBShGSyXbQEc1RhVsmnpBDK1bpPnIOe1Q
U6o2iOiMGmqM84uAG46RMB2OBnArKszQigj4p8zxnSeNOGfptDn5FSLnsHkZnMW+
KwZdtEz3JmPRBORj3P6FHqznLd0vfTm6QG4w4LjajVh6K84mTPzx+q49bqp86xwK
dBL+KXOE7y+Hfpq0wrFMc/piwel6oW/V7+5uuvIXXOWj1/TUpBAsbZLo2y9QS5sA
SpEi4F0EL4a3r2a5sT8V/E+rkZrlrQJ0GffA9k5b73MuyEyVK1vYb62ND1xGkEEy
YZW+ueUFuVIDftvlg4QNO9Kt8Kc+qm5OlwhIidz7qbap+qTfQ8oYMMCDEE0leqZs
kqjfJZjH9t4KgqKFJisLyquTrfN4nfVHMrfITRnNd0d9KEZH6gt6t+A/YK8M+eov
W4Iln4eF/DEX4/X5hdfs/9b9QrmvGow0mGCrj5LhsTr7wyGF0cmvJoMshki7lqdW
rz0685lQptsiEMR0fxNBE3LLJfUC17/PfezKV4xHXgNzNpKkQfQCFmQnEjjagKl0
Ar/oQHpPyDzwGvPebtWo7QLZyDOXviOXGMeYHdCEN+y4pQVanZid8aP+bJgJ2aub
tUtuPSDkxXdU9/Ps3tgLJg15qvXcXJw23rziNnaAKu2WH32ewuBJWZK91opmPInI
7HMVam2kmKBRLoKVAWMLP7lfl5dafgMIhwYl/eqtWOMdzA+PNC8SH4oYsZy8VQJd
5D/4YvwX0IIYBfOCmtGaZSJz32vCpohJhOaxUt2xCMwTCQRAVOWuQsS84+fPDZFF
hzk9VEyNrraXLB5UdRpK3udnyQTRHX2/uIMfUHQs4I7laM/B8GkLdP9g3jIZ+APq
dmwi30dAcmsUm9uINs+6+IX+x5Xve9vuQw0MplgDu2TW4k7ouxFiCt+ysFgj2KzT
o4uRl+jvG9L2nXUVbAoit4Ki82g6n9X5+uChKS7YwLVGi8UT7EZKw52gC4fHm0uT
/iSlhgxMIlfK2oHlj7/vrFGdlOvDMfokT6ZnADoqsgbclpVQ5TFa3IZm3SGsNCCz
+Keq12c8kIFI/8HmnfqNhKXzmFiBtUdseFa2FhpP1Yk7B3935MFxXcHTXoAVPeMX
QhWm1k/b3D7rSaNfprWR6BVZctvHhYfoJKt+jui6yLgW5HHia0wXgWfW+NXOHZVX
1XwFjliN3cojHkmQnpPWP+3uZD7Ocm58j8JsoLhMZSZDjoLPderIgwMLN1fmN3nc
glwyWT0Mwx5saS1ptAnWqDd0Ckz4JCD4AliFmkOoyYIqHNy6a6Mv6BKs3Tv1kHVv
0tif5cVJdmu9Hysu+uxh92rJqIOt8a6kDS7bF6DRsocV3+D0XFaukPPg0Fc3J2SE
7zaHXEj1UPQ1U9r6Q7AU/pbfxzpnRwrrt7CDVly3qqAZcbxyiLUEnjMmx4fw5XH9
4Bnx7JBmHi5IAjIXRBRBFGu0S6EspiVnDxLd+orkC6Wj1D9knz3cfp7vxBY6qEpB
owaWonhnU38KGuOB6QH7p4yVbHhj2omSBEhBS09S2w3GVvtSOsi6X/O0L9p8beDQ
xxRxSmKKXhhfJlr9VJR/jaOWJ3bl0AhlDLsShS3Fjg6gPESxLmVPh4ZjNWOZExIu
7QX4kEbaQs1058/K5Q7dCWwmpZT80kXMaUOZQZzClQvkfb+K6KvCq6m/C9VkFNjO
yJFVOoDweZy+TUp8DCA4FvsEySMA27M3/7ctnGJ7Jzt34zFmfra1RgQ3jE4ep1rm
Hi6rmhTvqyZDixvPE1FD1oZYRAeXyDx8jZRzXIpRJhfNApbDxTVaUNmNe4CSIKAe
5ECO1Sf8Vz5GjIPTD8WhT8odV/gHt+2dueovhDzHWVb6waRf0fE1GcPMJUDxsmyp
o8do82DvTYCXTdZKX3NKSPo8myvQExTjfONm+JmPKfKrKs1EO/7Vm115QTQZjRij
Mzto+NeSrteKb1A9K5sl47dR0seSvAaIwsXIXcrPSgPdvZhKkWHUIKjASJUz1w9d
LcL/znnv+F1h/Jt2oq+DbXadhQlEI01GRBPes86F4fEoFuFTEEBTUihEjJOY5JKL
BLVo6HRxuCbIohbliz2RxdED1MxaSz7fZ7J1g0SUc5Hz4Wt5k7MZoe85fsfmqKJL
K8cwPiymb+8AbUw33lgNyeXKXj35Sj5FFWBxKK3YrmhGCboWMCzvDeGQuhh93smw
/LoQx3DhIHmKK5eZBrU7tWT1r7I6lIJ0ZYYYgP0zISAmCrembi6Cc5jxvkWrw5jp
RQrREkJG8wAmPfZqE5CYLdbaNL1OUC6LZPpP9Q6u8uiwSbfcZUAhbxY1PGq1QPrk
pH/7iSPUMbtFawHu1EoHiBwd42QM+g7stznKfazztYpUWTX+BFRAhc+hQbS/WeIa
BnL0AqUWwbizz9IiaQ8hEj/V7VKzA/eAJBh7kal5xba5DDINo/YRS+vV2tQ2gk5f
CncvJ3Nngk1BDZ1adhC7MoLM5aFtT7yAOUWVNgwxiZWY0R7oJEQOWybs6JkGsZmE
wQmeC7y3NGKcKnF4rGrAeqLYYbvuGIf5p1gO19tw4gFtZyNFPG8x0cCfvxahLv9a
00VK8+c2aegoo8MBsIbXAgLEC9XCI3b6jOrYtGInz0/wak5l0jheghH/fLKrvFAY
3KfcrupCtnO06royBQQUvU/ar1K3dDMlAaPvLNOVteWeeRR5A4xiKHXzA8hYUcqw
vIYOHUdy+C6LBVNM/FV3nlIxhXz3zhEFI+Qh5r+sS7IbujW2w9f+UfN7EIzo759c
Q+v709+N/UxxqVtV51fbfqRQFiCTCUH1qNeXTLL3EelXQAhSMRweQZVN4UWYEA7M
No4+Vd2E2bxOOPBDSfIjhPnjHLDAE1Zmvq9qhN943cRvVmwJedAEwwcbZxJoxO8j
FoekXaZcakxZdiO6kWJw4qa7s4GYnYTMLP2xJULtrBlGXxQtISJexPkPHnzmxDc6
pNvcoUMnK59xeCZN80/7fnfE+z4zCkUvrBu7R26TJsB8torktYXHCA83CWCJ9D0c
bHjaGlvv4bUQg8vWD7a77VzowB+tjF/Aj1TgdA9HyBy3LsCj+Tgxj8cXCQik4ALC
d5CaQYdDjwDUaGrPgm5gIaSiRTcCfL9cV0L8DdyntpuNjiq01tcO1DmC8HCBjs4g
zsbTAV+WP0ofP5+MWnvRocK2L1dOj3Q7iijzGi0RR+YgQdXLDSU+/nQvjG2p/24c
TfY+siXMJNNWVuL0bFf3HHiZOU0tOiB/WulZ/3en/Ld3KFQhwZ2w1URNrvD6I7q4
zsl2aKXs323hHTHDIuiTqoXkD/DRfchvZ2ch9Q03Aqg0wnf+q7z8N4bvkm7j6OLb
utCofqTlCXGfC4IArvanlr5Pdcgdn5Gq/kKYLg/VU9g2wWuesz7/2mdS5FE8kKJZ
hsdiZNVpA8/2Uc9WxdSdqn8Th8Cn7CSnQH/wC4W44/z24wOivmrEsVZVs1BCs6G9
1aRN4QgqzAADGQErhsA+vxBg8cLVZTkJGXtR2g4gtBRh1xIn+BcpBp9KjTDJ79/O
rPG2WlS23MWT0+GHIyi4x/EVQMfQ6wwp0qm16teeo1UI9TO2B5mursCT0CPDs7gk
nq7aQ6bjlP6ih5mbgqhqsaiXkONchhcbcwqk0GFUVrx21zXWgRzB1JHrJkWlo6ro
TmjA3qSUYzpCnqGfuqJdXlPi3nAVF/ZFJbNcszhgOb3x/3xLt0dEePU7SlTHx7qF
6mQvnEaIE0XGS3t0CUcebZ8dk7OIIHB8L7LLmrRxFjfW69Dal28aUHJf88IH97aa
44yaaNTcDtdHAXz/9eEydYlMfbDyvntBnu3OrSCuskmA25cKpPTUxY9aEHZc9hat
fM7BkmJBhDaaf7Ch4PROoN0OwF88oZD9ReOkGYZ10C5vknXyDJRkogvW0uV4tdCg
4tAvROTMhN13Fm5UBTkTtoHxdCN1yBiEcPlUeQu/eqSUSI9Mo7ZYREYnVBPA3r+T
VADOpaCaGqH6dHl6cEGWkh0ysW8p9HNyz3lC/fivQ0yYezAB7UMhLJPlj1XjMuKD
kPdGW0dcIC2yVF3t7aPWcifpL0bxXMlyUOKhSoPQ4X9H7PIKCI8mLMvskIzlF32x
Gl9VLpbndfy3CONNn26vsUq81i1eH/owmSXLTIqd503eEyspbFj9xQXDtGY2wV1V
eYeinLWbh+WTgLDkoacaqD8Z2SyW63HRmVP40371curT/tOCZ4391pcwtUoSYXtS
nhhjnNVglXTFbLzU8b2foK1knkc98bQ3W83s+7sIBEVYDfwYBo+U5loN8RHz6Vf9
vwgQmDBpNhlFy5lPbyeZtAiR8p/cr82lZl608pm2OgVir8cGr3BxEtHQeYXMYPGi
gKPzcUSq2vqMaMX/ZxQcqn+tH/dpOkGNIkbxiI80jyYmIg3Xfbiz5ATAZRGEzegd
gOysz/hG9Y9vFfTUazeOkXB8HpEhDgcN16TT43jVgRxR0zyJ1rKzpT3ujav0gnho
ESSwYahe5LtGH5DdB5I/WpF+Eg1KwJh3vbzQ94POnBoP1HlVagiZTaDi/Aljpx2j
1atW66/83dv12aqr9nSaZh/p8Ixz60+TG0I5ZhRaddF65VsPn7v/6zQpQT2jnaM4
CgxQ5W93SEvLdSMBICmRR6ORRKggwrVySrKztiXJ4GaIqY5lGpRlvAMEDnkGsH7o
8ToAJFarrmyNvRV7p0igCxVjt7UDb66NwT5lUNH3CVt7mqtlbs+Sg6Jfp8BCcUue
tGyDbCpUnyz+TGxF4rvcSt3ZQ8umzpcR4US/3/iReRj5poDJVHpa1W7dF3wAoHAf
PpBBC+T2iOsLcV0UMSwNhHSTflUlOD3GoLIy8Rl6Y8wWdHN9/s7bJkZd+tEJpwbS
FMYeCytEou5my9oIL5x7wCKE2p66n7wwXm/UQzINetOgUWP6Q2UBl2muI82QgDrO
D1TU4f+ltr01tZAa/kcvOdVQrCGV7Yu8Mq9qS94tGwW51GBlsVtZit8sCZdkhhu+
R3JHPiq1JR10ve14Yd+DHKP91IrpOx4xy0zk7409bmw8IdWIU+3UnoU6AUGA0gzb
g6FGZAFKzUvHn1cCPa42WaGJNcyk+RADAQymms/ZwWTSY7p2Gk4VdA51bSP9fE6I
5O5WqGoxZbB7JKWy1F5A+NQWIauFYmjz6BBL+oTenOo5lclQ+GVEc1XizcbE6XVA
EtFOAfd/oBc6bbPKsS1uyLZYGto803MYpwPy4lCUfUphfvS4dEHvaqkPvw7Vihru
lsJzAeOxO+RsaFgnAjuM2Rr+Yxu+DY5G5RIAlOCieZ8T9zc+h4m21QBqoE+2mBlW
N8h+pPF/pocsOeqWZMebEDkRP6oxK2Ws3jbXZ8XzseYo5H7XZKFRi35HARU9MW63
+8a61VaDzGzsfH4kcci58qvYTdpLdXwitZdxYDdlTcU6Wsr9oyuZ495mNkL2ELij
xRNEq3r53Ull1NhMbrtzZOHRpnhIDKVSLUxNgNOTiOfTXoHoEJ0CCmUvswMEvpPi
/Djyou8tWPHhTKR0SFf7cQISUsMAyg+mflFyspyk3F24oKddXhHowPkE9vrUBv2w
iq+wdqNz2yK5lXt0DaEpQKS580xfd7q4GtG4yuetDkX0EBWQtRM3IQQEF7diH6Qe
Oz6K75+Deb1mz03O0whLzXf8aaJvY5bCY1yNPEiipPEXGcWwfU9SlT16Vl1JzB/g
MLm/YKZDQ4LHYnDjnrHBGct6vEG+ZsVrpZ+9enhLsXdawNXTnJqNOMGRADadSlil
+VHYoDJyRDbaxPjzMKhEDRINLFS4dyyQ+zoR3OXcwKqxwNsLjYivpZOrD1Ron0B4
DFoKpJ+k12FkAOzmx4YVhV8GHLpWqEMBNwZnqWykbvk3z6WjNv8OvByXBm05KhzB
aIqUnoHl3AH/DbvRb89qHA/oRqE7ToULDIk2ppgH3agGEyVLIokLLnoLQoHf7Kud
y+7q6lx5If394d6EsLabWL/9DQac+xNL7byFJO1cqxd2ZZo2HkweUGfoeacEJ5OU
XD5za/go6ajVqYslP9bIn9XzJRxTLDGW2TP8HwXeB5rfxQ8bJdCC8gNIwtPl1wHw
ELJxQk5vl6pWJQAl47vnRR1TPEXo1etd+dyioL27IBGQdhXEzDXaLJY7tEpd7ASi
VeAVjEoVSrrG3Par2MgE1jBJncDfODpCt5TCFjRunibihgtmxW8yPv1nPdiX6vcV
DZUjz3ai4JsdSXvzU8n4/RAUwhwjUSFGABfX7Azntaz0MBPFxiyUSuh1X9/mKPmo
RuggiFPyoqDfVttDJUG2JXTY/pSDIWUtOgCh2FSBM+6xjCuXHg/RzXlHA+pQUjTI
UsnhQ3UsBPkOkc6sbtPgXUfxBbKMeNiZ2ckSb7oecWekNVl7z7YtGDq+4BtRA6bg
WCFopF79LiKPVi9FCqTkMXYeSiPhmKNgwIi1BNzP7wsLJuJEnsMZdeiyLKEIEoxi
Kx3kjpX+53G5lopx/ue/tKnj0kZl+Q0u33cEBdu0sMauv6qSKOM0VoaWdkHSbBl2
hl3pOdMnBrODJBIyr7q5u8yPmta/gHsGmCxq4BrF330qDRj1qouIHQjh2mq16L0u
pCd5c4TxCZM7ihFt3/ClhnGTii5p+f8Mw7UPTKUN8nCRe5UG5thjJTxC3xtJdSLl
RAUzV3Iy7ZX8G17Frdbkkf2p1LLBxYjvsDJRYv0iiBpQZ+KIRnOuubiZAJfhejuy
SxQTa6BpBOEw2YnLSVDWjCyYakClT4QcPiBC7s9pr7Cd2oVdO5U0hKiF1rtN2K6E
YMaXY3UmwlZcUarVwPCoVrG/CbAnsdwjdQOedxx4d/0wQun2cZnEKwr3TIXyAKMn
UXa33sM80YGuFI+0WiXgY0xyT4ihlqgr4E3gqXsFwN+gtzZe2fnhCdf5uEiV1WlP
QnlQBR5wmZZJmObPdEt0+/vq0eZDMA8fs1YH/1JRSppHq4/0++YIzZI88hSo/Bas
F7RTn9N82+r/JJGaf4HbHnJHsFVIU89WmCft8D9ZY1qVKTBZactaungvMIb10IDX
LmeZYKlPIHV62446SGK0ViIICTlaBQXoLuR9q8uFnrB1OwFPvCSBNsBEiS2Tpq2Z
SigMKUUgxhejwLnIaJqHwK8MYqsQpbKh9YR0iFvgF01Uq8OyHQmsGRVbA+xLyMQe
WLFTZayx8x4BhmTvN9FIPzqQ7a4rm6mfNXHW3FPA+NSxEeNcr9r12TIuOcDlOLbP
0bVcNIJCK/aB/7vQjW4FSQj8RDyGDs/wmdRnRz9QcEn4iX/HNXF/t9JsX8WXPy6E
qTOnC2+2fRg+8weXMi/Zb/mnspvIiPjdUd17nLhqQ6mRBDR1DvqDF9fhmKRckeqQ
FnmRnBqaEgsMDCPEm/1cN7Y/li1N579qB5cZLqAONU+zDAboSrn2DGR6PietqBkE
Xj1u6AfNlzTOjlqG7zw0NOf8l/dCy/4hhpPwKv5+oE/XORNeqO/tRKlV1vsHlhNq
fujVsDgxRrqtl8j8sqasnwZn1kPaFP26svWlgo6YJybQTLscD3UkgqzPVcRp54NC
EQATGRzqHKEd0vqAcxfluKEwcJ67PVa/IMYUYMCO+m1KvUJqvlGvMTWBqh/ZVP2P
Tzbwygv4r2HhBo0mlgM5S3nNsmdTIY/Imiyc4HDjNPDyhH/Dyjr0y9qpS08BjIY5
jEI7pEN4e0B4YJGRkcDV8qE9VdsZLEyDpYC/0PR8wW30KqlzOWkpITJSd3nK52VP
JiEZUP8AvantwoYqGdTwXnTGNa43CfiWlwajdMtAIUozhhJQzp/O0ZNZtI6K/+gv
U1o0o5K+XGIDmsmuatlisA+tkFXDiJhlhr29rmYJhao43bEsQjxPzNJ/GgCN0f13
SJssoIjZ9HDOnN6jLoHmFNNMJsRIMNVzQMRoUPl6/+il7cJwCh9Ut/IRF6ZcdcVI
9jBLn+QaxBD4RnvU5cdaFpq4+u8Qh0fLVAYNA69o3aIcwb2MxR4YVqzYGkkg4/14
oCw5Ug7BSymVtXnLP/tDilR+0cyHPczq9G1XSeQQBd7pYkHB6Sk10C0uD8dXOuSX
IRS3DnBV+5lsVn6Y+88o6jxHsdSIJ3oQmLIlKUOTzHiuXpOGznVQuqcZ2dV+az5T
iCXvD0xBQR1ZggrRw0+kL69p20n4CY84y18ynXKJSCT2qMNYRv35cQz+N9Idu2BA
/vVOBKqhxn9KdmjQ6r4jYgA8ZOy+0pS0ULS+cR5Qq3+CBJHvsD1W2MygHtYs8LrP
lWDd1/wPFVMOWKB2wheI+n95NiHSxMq4HfG5mK9v27ngoIeUoiTcLrtYtDHpneBY
7cRFkYEughtCgThi/KKRk4jyQsNYHD64LmQepPC3UbTCbDkyWQ7sxRDp/IX+2pTF
9bESBYigQYUmdbYqoukEflx7Efcow8oxwdT2KmqMyO60i2PUjj/o/1/yLAsDmY+7
WtnLTrK8n2dOXoH7Fx/I4F1HGf1lCsNgG2HU5C4hrfAUasG3qIyPMXg0tUWIB1s2
mSn2XPUI8iBCFHP0HYWRPajQWdAnKJDJ1+XP1WA4OOZXFkQr2Rock5U07Vw/an9A
FqLBsVwrObHItuEZ5N+KGdQIfLqIywqurfF5MAorElYBwuvn3SpJXKCH9zHny/O5
qXHX6dp34QrrqLvMT5wCADJcr7K6QlC4nlUmt4Mcx8FTQHhQT7ZM6MfM19MQ0py3
UZ3GXX9rG3g5lY7xkd3aMDSUwz9fv4xg3mHVWg23ts6A2CNRY7MqDZmz7AIUhBaF
1IeY+BbM7SF9m1O2FrG4/tVrntLMqguGA/tZXd66mQ4IwzsXLqSgYVf71Zb0H0fz
b88BcdBmU+mZKgX9Nfs+ILpzL7hFihFgNjL+ndIjBpj+ls6/bcl8dyFmcnojRZt2
MTSW2TguP0iXAW1/tyoWk8q0/jyzIgXniAgDQBtxuzfmHBEZ4tSjOi75yNzXRCpn
kks/ZBAXmAQU3d846pHmr5MAJgVnF76oxXISQChlGwY9CqdOE5juSlTwYrsgjd5E
LEcRc4/6G05fvvPxLjOQ6TzhO4dOf+MHptjXfzZ7TjEG6QJm4VSNvhHpXciVRGlX
ZLNNUOSoXFL8SGELLELSvmSfKvlhQZ/EJ4mo4J9+GVnO0q6ubdjkND9Jhn6H3AEF
igzA7sTuuwdGXD6VyNzIil53N08Bc5uemIu/ynyHYd6Ep8VnGRIR9iUTNdMkhMvn
RWCIP/jGFXBD2L8r5n+RWMPC2SVxSUaKFPRFR/XuT+4pH4N3NJ4qoXE5GnlqNu4l
or73Au5ZVtJ/wBpgaxepwSLGmmiSq/3D/kHPiMfCDMn7z68W4rag4u5JZR4Ptxoy
JKF+I8EwAeSRPBN7ECUT0p7iM/Aic55cZUj2mRMmO6D9UhzeMWuvnLMnNggEID9G
Zv98czjUHC5ZjPpM1Jzbw7bftRAn693ow8WV48dDej2nz17AiOL/fSwe2gZm0XUh
CK5kFGAuNmsrF4V7y8fY/PxQMocQi91SvVANDYG8u9XgAs6J8TV90Sw6PmW1EV+h
n2C1y5DUL7AT4AxXPqZg3rph1eUPoE7UnjnGZMY3kLjZzCX57mLrW7YASwDAE+/6
cLNpUXEpwaVO6XlkHtE/iu6VOVbR0KM9XItSepNqxXDwMOvGbDyXWk8VozDCKoA+
cnWfuEFjDuUz/1OMIT5LAnqWiFCXhlem4JzMnqjpJYj6M/UG9+jUiyHzD9oIMzkG
I3q+5jNxumjJLqvjQ6EjWVa4+Jry8gfo3ZwgpKr/d5Cg2BEs5IpKEWmNrZKKVbZr
I+k6/5JKftJhRuco6gNl1kD/H6s7aRvNVMKd/DvkorD3cZ044U1P0msHv2No8lcj
jEVU6aPUx8SQLokP20dqIrUIi9+x6OwC/OLzD4plX640qXwWyoTYgA8x9wiUi0gt
cxLqI0n2sq2+lIybwB74Y3IX00Ssmg0RHOkUCX7ZsBE4Cap4tXMRuRGMK9P/akuD
AUIzX9M+bYDo4XhjFs9x/LrEPAH9w6sWy/l/fjJO4dgi2dBEAnl89jOslwUlc2de
vbb2mDzSaEM/h2oZ3dzQVXgIUU/ifkvg8nSJ0I5Agj9SWgW703PQSX7xJQd8d7SS
7eDZukDNdjjEbO7Q7qqNoC3k9URCq41/IubBpIVaQlx+B46pYLS9J9zwinXg50sU
Z9X3PdH3wu9oSn8AMNo+b9ZUd+Ypxkl6vwsm0A9KWwT9illluEz4SPNJM6Kt7cD1
+U/QUlnfEyuQk2jrAhFRtBYxNZcillzw6DGIqEPCit9yfukcIaW/AKETxW/tU/bG
N+a6Gzom79f+Z8mM4x3hAgtQjuOzLmtIDIiXLuCFV1G6qJw0YWpHvwCyHst1iIl+
cptfmtAgPYVDmJ26/Q+/IJaVgt9vKsoK18WMIcSg7I0fg4UwxhUGRFPcjmYNV58W
jkR98JeTKrOiJj/8py/8yJCwoL4NTE+ikXdQ7nxvkHSYRveUZIfZoLdUQ1pPCI8g
/u7INRi86CHZi6n/l18dW1H7Ezc6C+C/Qv7rmdTAFlIYYf6wLTU8FS7BiPGG0YQw
eybIoo5xIDUX6va4U6qIJIPl94scBLOF7NnJe80+Bq2aBoAb6QEaplMNi2QfllX1
zSwHrwvUkOaeGNQjzEf3xlNBP8TwmZpEi590ECxwju98/rggwh9qz0+HgDCaKOQV
cNghGWOtMgctgiIeNC4eEMUbrvbBVrQih2EgaFPQ9M3+5cziADYIBR1UHyKEdkVf
y8HL+0hotBO7lp8aMBUoiupYQ/dSAPhZD0I+kR05doyspISzVLvqaeG+fp8a4YwJ
zdMrdZiOVvDQJNZyPKNHBBszZJavuST1pY1OOl5g/bMGp6PH1vL/b8W51RyulT/O
OlEVkMFr7il2nqkEhu8t43BHoIOf5J/I9GrOFO7kjIEa2t7pH1OAxOR+HJLLzXUz
sKtjoQOYR54Sgrcl1OpSmmNa37YrUy/LbC5Xnv5xfrNRtMpa3x6H8y4qWhLDAvQv
ZLbBUmqVh1ALhQI4nj/+ZY83dL9h92UNZyicfk+CDVyG9UebPEhI73VsgCf6I5x5
o8I2fpWVZOI2X9y2IwoZ99TLw6ebSB13JcuHhUO3VIcrxA1aDpy6KLcJSHQVr/AR
nu8P4JYTlRxY9DhJIFwWyuKrfWM1rDqAfqQzx+hhFysbNhDl91Kv8K2R57+Hb29n
+ddu/yP5uonb5cViI7jfhy/K/XAsp4yzngqzzUPGd1/Iq9NEWWnHG2BNpOJt0gj0
8ZTwFX1ngX6PuDuFiU1KDl5x34qWLkISWj08+5dIZEif09JPvjDOnbIna6elB3kP
EEB5xEoteDHmBi/qc2p/HIFksDiJPcDGVAbr51DPZlSJ8PIcgb6wUmMBDXcvBzau
7LmE1479+9WKmbQcKgPETtzk6FKzhXJJDJcKL37DOs/HBgzxK2dGAGAyaoI+seEh
3q+/vjPEEOpS/P8uszqeGrKwr0/O8BKAtEmHfYIHDbSnrK9wBOG8DtynoQWjhjBv
ETWzHvwmZ1xENH8GX0Ene1dO21OQVI/27gFiZ9vK0tYA6ux3Fwj3RcjEtoF5mQX2
bGG+wkZv5leD28/Gt0sm8dXX9fUutf+oejejSxJJ93Cl36sXdlx04kRzZt/+5LXR
xJBu7YLEmDCa1dY0voanHVVUJ+96dsMVaySIjbn8Uor8ntuemiJAqvtDOHjjXj3m
km314jAfFmVc4HFIf1fykVrCXZlkau3JC7cSEzQa1gOIw9ypyXRUiH2mrzJQo5A6
qkVSrfMrZlJftBHh0O5pzljotf1gRit6HgfGvKuTTQhK2ADBewfiAmUVdlFSLxla
aUy0hheKIoDVFsnrUZDiZQnsozEiQK6rOEuiN73d4vfW0Misf4b1jvAuqCNcFMkW
wYQu10d75gQLgsDbHhIUZm6ilYHFRxRubUr6SbpVCgR/lCBQY1GoJhqarCDEAPUI
PH7HOClf8zpGiTfXZrG+Wz0/2FcLkMxaNdxAJXJ5aliHAb+FU6hpRFuSHW+3Nm1N
rjtSqeHtxd0lIuIeRUDF2SWqABHUZRfcjM5eVkBmcLiMaI49l9Pi5GqKicqfyo6+
rGDO/NP56ji+SvF8v46+kCpP/+XgN4+IINwZk2QnduDC4LMizfceI06BhUGko7oC
7KPuWpYLF8ictA0l3TTl2r6XRbb0TmL2a3uD/QulNkNQSUEKNtykeQcuSKdPu1M0
nR1hMs0eEHa9NR67huTjw7aICBEHgu98RQ7KQpSGiMFGceTQewwVrJBrjFqXkyJg
o0Hp+X0eFWXlEiVTE9p/voTGxGgEj0f+l62zBG96Zwckbk9HgID/w1olJHyQhrGZ
PMwGuWYnt7bH/sigtIc5ycATqLAux7v3vb05X8pxMHxGSh2WkMN1NQGGI0O7S3nR
zXV9tIzgElWUfdwtYqcURGSxEkgaslRu4YIMAkq9EzOY72Ykfusgf9DYCZxVKajW
TZl9fUs4VIjWxIt/4beZAyK5BhmOeoskNHzRvuzapN5PjNhnQKf8Ho1UuzXdSf52
G2jhq28QqX4rMicvh6zbqAR0zvNoP+D/kAldGot8+4ponoBpTOHiXjI/sE09G/Io
iHxROoZLO2G/e/sutxxyqyWc3fp9ZHpnF+1Z5tYfc7GSMb/LG+ogpOJTbX1xlcnf
jkEdkTzWoxIzpzzNfGWJlow/JX6LE74lFSBM0R5ruy+519ETo5cHOa5DOMlCl7pw
lw/609lSa43tmlNtiIBHa5UZjbDkJhIz7yEmQuSEdLpSh/BpzTZB+SktkjNzX3XP
Szgr64egwCCV9yeXiGOXL13h9ok6bKSSKCjBSBKLxCk1MqVhLdugTMm6bEmF8g7Y
foqZMI3N93cwKYNcn71/Xz+/gCCz/U/uVpfeeamOrBGODIVP3BwskFagXFBbOvE2
DTN7Vkv7Yx4aqsu9AaeoyvpQX4Qy7BKNfoqLse0xfHsxKtGYsnP+c8AYvKFne4+G
rGOJgKr9JTT6U4H8MX3eInHqi2F/XHbhbVTuSspkAahX2316shJ5Ny2xd8P56rx9
SRhiiMkaWiJ9fQn1mTq+AZiyAn254AR4TkwoWGaeRfHRZaDQ5RD1D9PFXeb/yGV4
BMKybTtnAMMdnkWVRVFj2xkKwKY9hMmcRcWzRaqPjaXffFZfh6BMR3V4/9ox87Ah
IAVQ46zBY8a+tWBdGMngEqfowhVcD/pC5MOU0av2Iq0f/GUMVZ/yo++ieDhOBzmw
/Ry2FB6CRqiHw/MbpryrCws6fAzMlXTCD7lVi9QMLqDJvUY3PzTYjzFunXoxkFt0
4QNkOcA2jO02/8/wt9wOjmV43GY2mt4GSyrpF3Be466Zl1GzKy73dPIPVvs5m0FH
eDg6phug8Pfh1Sd2uqzTUkV0Y41aFXHHwpzJmY3fp3jHk+phBhqoXGpf1tuGxXtN
skSmH56jC56qfUQIsUf+2Ylcrep+XLMfU/2fFM7kelQNZl917PysN0Ve2qpEyqAs
xCt1ycOqbbqWKrNoDK6aC7sOziSIl5XkEe5UsSPYdECK2W1zUutn4hvQ8oTYunRy
qQMCL7PyCN9CRSq2uYxSuIVUqUCY7C+xQhAyj7sSBy/BAnpDK6WN49W7jc24AeEv
jtEZvlaRankj+yTnyILv1O5P2M5gjn+asrqBJvtvA1xbIp981RPwpnRTQlx2f4jB
fk2TM0/JcVAQK4MrgK3n5Zj+QMxDBSIU/FGlE4OFs9WNN5IvszLjo56u9Lc4EVVm
7kDXroj1uKuRP6QPIrXn5zrvWxIbL2Fpmwap3xf91ja+krhX9b8AZVG78tc5De2f
8oqVzCf3N8gaKTnBYdLcshgxGFUmAs15ZvK3h+cDku1gJQ6wZ+EaoLufSgLMBwkG
4FfHHF3TASEBGlbPT4phbTfdWexn8yR48OiVxfMkbYHhjtJhvtLAgZHDXaFuTYef
/Hg2ovLglSp1jQ28cdeexq1K7me2BHshQ8e1CW0VQlbFCRoNlmOLDOEFrXhqlFvF
oUxkrHdjq111yXU+752eYwkn4/GFnZXnxBVirC2w+rpAfdFmGgnkB6rbjcHsJ7ZT
WgXqw6n6InPdcm4WjyDy+d0VrMXvSEiW/ZlZzw61pihltbystqgl4FVUsuQgkf/1
KjJUvc5aSShOQDIbRuEDQZSckpvZ8nXxJFObOLvep5/kHbKVNoVonaTLcLak2Wod
7y7pJjEg0343LOarFkeGOVBt5zq4xd0JNwSM6t1akK4CsD92XGZpnj1tQnntZp0B
pJAWlAATYsG33okYlWJtcmTjmgAOzbV/BVljINi3lchYl6/L9haEgYE6MImXDfES
v2Uigyt1LZ5RxNuTeDAdwEkKyk6WDdW1FuM6PfXmLG25Q4C53bDf1UeCus2WqbU+
ZAkuOwK8WzZeR2RvH3SpfRPKeY9lUazc5P5xxCSUEtQI7HEy3l2vO0tpCiYBK6Xt
KrICfE9s0lL0k3iNzKv+PI7kzggzlqHWqikOJ4lYOAlDT1OJpRg3crTniDle+Su0
jgoK8UMvh9/vlcVklXODkEfBaMB5dpdgenIZzYq9gQX2y0qjLNhlsPhIsLZ4wfFf
sDkJaPCyvYF4IiSRQeO3aDEOu3qi/4CXbWOgfg7DoMVQynK8m/DAXkkBuhlnwxx/
1sB03uSJG8qRKOnpJR8/GDWLgEeVlntmOQB/0Y/OCZoUDiMqNt1drAbOHKPR3fII
5Q8qZSJsgvRbTeWvoHT3hWk5Q/heALCGglmLu5AY9AR6PJ+Y6qw9dfxWghYS3ow7
XufOT2rEDzg374Kf3U63Aw69BHE37Am6h2IPwBin2q9zr2OLjv1JdLQw2l1AK0kZ
/4KetqjytmMtfnEYJA5ZDC2QlMiuMVAcK5J7NUerZG+C7FQEAfQ1qI2WskZGzQ+W
sePcRKFoF6ELgp/qb4TXlWg6cvgy9sWpzqtfFBCMmO8otPFmjiIq8lUVF72MKEBq
ORdYgRleCnuDJFQq+pYp3DaXdhQMtWAc41DAUvihdRPWcz9KtKAmdClBe35fn/7Q
WhiG6LvXLylnNXtfGtumWdUaFWbbdgPo93HTwf6UVJvMEZF5+H2dJxEzO4QCwYF6
LXjbJhqBY4oN+mM82etkKy1oTJLk21Y/7aDppOSNb42sGONiUEHDH/sGOYFq5sCl
/MlzIboCC0aHICW+nDWnFw3GurUqanKmxWg1GKHAQds4h0chvuhvJAdTiDAzJosb
xUGY5//864OLs/KeXZT8KvW2l47m29yzV4luOQpNilX9b2O8PiuSwWeAM/gDF7Ie
KeUxv5ebGM3LYU1jLdxdJYGHr5jVEB318voYpEsoxwJtInh+gxL15TcpqezupzI8
bzBg1m6xWL+b6NvQ1f6NvIab0orBrfLUqelVtfMbtis7FIXcc52oF5dliqY/zE+8
rYRoT960dXdEopUUgtZpJshPHZGJ2imQ17Ad2DXQ3YIcY5SoD+PHh/8wJC7/kgtd
LK0rKfh8Uf1V5gAp162sgc+uPBKB2MvjuJdWveBDfuJd+Vypy9R2Pp/+BsZBnht0
H5UATx/EstRG6lT1hlitQi0kvwMu6rGfJSjxm/Ab93GEs5HsaatYu6f0IKJeIhJU
8L/MElVrMzbCQSp2fT0nf/5kFZbr4zpG9c9Br8dkEOwtN75S5t6Wqg7bV+C07cEt
gBV1Qlz9FU95DBWPdTnZBAIt6dYZ6cY8K9uwbYXKXbw5NOVwMQfH1Qzea1fYwhqB
J3X0kt5tGesEDN5oNEF1YjVUUJ+KjVo4iUP7Ab/XaMI3ex43CedtumfRlis4F4Tq
eUJas7VrxgDxMMr/vX2ea4TYnwu1W9PAHKTM3F0MyqRzqYoTtbvPrsgmZKJP15+n
z0HP3MlycQZ3wSiqnP1I5hWx9YmSyl1MbzjOTVOmtBKU/57CI0SGcaFhXjK5dHFM
odT1vUJOOgUui1+tHqcAk0bn3sZyuqTnsquwsJc1MLRFjTxTc148Ay8mIdO/8l0M
XRQC4J94OKc60OdsQLtliii1NtzMT2P/IFuIeueZg3ZubfC0/cv1CyECqyqjCi2M
5NKHPXch4a/C6CnEkzO/ZQvmX4B4VtXTt7+5NjIoAO1yWIk+eP2xj2+bk1cNyJ8V
NguBXNCkqeLVmVrUoo/1ge95kQ6p0mBbOL9k5j1+CxB5FWkxxPtmf7VAtdEdbcd2
P5e0kQpI/6GVp/D16mEG4ZsHR5httnoYbfrHDdLIv/DQex8kFtOOxMqbixHUvC/E
+NIsCdZy7zJ1LT6mjKDFdL97DNdC+vdgOSGmcAWHhqcTzfrrBIcAPlA0QFeeOuMu
u9u7jVkbyiMgjiUiAfdGIAdZvwtqnKJhn5DqBEY2s8xoDDabRtscAo13JC89DMyH
hgaOauy8/V++NM4AD4OaI2RTDZR2WYArV07lFEgGUy3T1n2rw4NQdwdLLlKn64rE
7yjwIHJgvTVqXTt0b2v5vrn2Nwq60pCbwssDxbm0Li8V9pHiCH7k+k++jM55A2tg
HVp2PpjdZMFxVyszlvMaBoFjnKBDtZsy6ef2Jmlo1K1PxVgziwRhOONKNTUfabMx
xrIuzzZehhbXbjGa7+jyW38XcjGVdrzSVskNCRzsFIRkWtKL+iC6i4ZqYL2RA81M
9S3zPtN67Q558pj5dMBp+V5FU9qHg4Yk2xFaXHq8URE+4dd899EMwvXqMJ35IR9O
yKGH6pgffNg4D072vJr5nbdGoTOKQtecOlvBx5lExSyrI/gHqmg/awAUnrm9tUY+
pUD5m6/Bkz3TM0SA0sS155UXOU72446f908zPhFMFqt5avgEiHpZ4NejA9pIBJYw
gJRcvqd7245uPVkUD+wgpeLP8xJkmxcEYhNoE2af/N7nOhMVmFcJhWioRDQWmxkC
sjH1VsY54/5xH26oO77uBMm/fc9q41j7FCtFp8FBaay4aH9nS5+X+Y/4h30LBhTH
pReNeV3nMA6i50VLCSr0Zzb2qIk8Sar1gVb+0v5IQigoLFWeAI7kkNDvmPjLAUd1
KsvTLkqCM2SaGt6T2V/IGqG9g+JPm8Jqp1INrAjUFGTdhDD/wSeB7hjjbbdxYHJa
wqQx5KvN4VDdg+gxkY1WCYBM8YD6y0AEwTHQRTI+m3HIKDgpd3pATSBh0LFlvlMy
qMkf8O3zPVEAU7h1OVlTWRry6dbi9+0UziM/OlC+Yj/VHD/tpQ1OTlLUi1038V/z
lfFClIz7wJ78D2JEQKl9wT6f+k3ZCfbP8mcIy9mq+/XEThdGRq6NwVSE7+rnuo2H
Qb9n3DveurDPAhRAxBrKg0rMR5s4Ltb0einhMBPM3M+OqFsQsuB0y9Ya2KnTVGLH
WnVTDRWchufC866J4V0W+296shUALDQ1W9A0ZCbxTA1byEh0jFTpzU1M2zw8hg2D
f9fxT02W3NAHSTmMYIh+FjxXeln/lWSJI+yvhTce0GIVImKgWXcUM0CtRyJj+xU3
Ewff13ZDH383p6ALvEADeRTADEDXsGTr7f1lXDRl9mtA00MgoqssUnQGSDT2UOgQ
9sKOWBF7MNcGAf2jNV+z0OUbzcNp/TZJX5vPkzjfdsCy5FQqQVN1f2UHPXBLOprR
K3+BnTJGY3Dh7iw0n+N9NkDDcJraSgRKEVQOasQf743JzOqO666UNqZIOZdv0hOb
aLEmnqN15/VsbC3lQtk81HoaNgHJAUHj7M69lR7Jduly5DlgB+X0k8IcxlrABsZd
ElIie5WrxBQcGQ0V8JZLUYbmxEGYrWn5VCeiVC1P4rFQlF/gt+Fz6SNH6MPhwF92
Sal5xmsV1U/6YqqQ/p0PKKbhJpjoQvJCELNh8AstXKDsILIG+QYOM6OAyItasorL
VgDtE1vaZUzdhrED4OzCuOAFk8FMCNPeOEbE0SfY1Vc7wJPGAzONkNI4bkSwvZNh
auu5IezAhIYozEfFxK9fssqZp9EpS8RJHaBZ5LmJnlN7BKCUof+cSoa6LgtvfEFj
AyRYVfa5TVaaQc+ofpI92ogt2Jz6iEU4Ilnbqw35RLGlk7NCNsGaDqE9gUCKMBkK
DXeoarcnEnl6tX2O01VHVs2cc9NgZBjHc5JbvumWXnNfUF7nf5d/BWvFQT5KsJ2U
WeCMyXNOyDWLdgG1mvYTJxhhq2I6c7qYxU+CJEuZ/k2yVw5qycqeaOBMV69S2Oge
mx5ZAFqykXzQ5FrHQ7S77ADf1yldgE7Rv7WEzOeqN5xjmHlr/n1nBtlHNtt7lxos
r/7cUWMeEGZI1bN1wUniQXkE5JYG6lVwcefh05WSrfT6Z4RONPTDKJggS2Tdsje+
NSJ5i3lrnoD9tKpTmD6VmRF6JtyBFkgFMezHbRHg8+Ws4hxXSAq0f8+AJwtUo7Jw
x7nVBa2fIatKXoqvVE4AbnR3Jyezwml8tmtyoyGZliLWz2TgCSgBFb3IjZmkw9Or
ZvcIswQrm58tJA4Jq4shyZihtx/NPOO1fKrmRp9tlE/Ra91lI0IxiZhSNvXq6Mv2
X2P0qcxcH2at+RnKrxL/oR07Y1XNDbbwZho6razv1YOvoQpGZ1A+zcaOnNGxZrJb
i6Fb+aWTRAanHucg2tMU0g1lLOzjVGD73w8+qm+nj5f/kg+ih/f5+bwou5GP68kx
BxVF5iXOAWy6mvgujF+3zk+tNqdtRJqhYa9P2cJGXAQQW1l3iUgrHhqOKqoi/xeC
6ksdsGPQ7PJyDQNXpnqKlnz8Me8cW1fauy25+Sfhv9xddg0uX+FP4vVFvCjOWKlS
oBX/wz8n4m88AvJnAQO5OVgMN39P01e3njTULVZ5mQ0AX7nDMIyGUPz9oc7FMPZ/
2D2tkKEw9K7+Kwo3/2GaW+uxuloXT2a+auaVq2PNC+c62NOdK816Xtv+vI+amb9h
UqcY3wpy1/hSxQRo+gCfKFYOPyYO1IXXk4s5S5uitOHs2sdi17eNReBS6HXTMALP
rsSbb/D2e5rpIWsnjrYHRM35Ue5Hdl6QZW68JPRFYyKSlyLuxyb4Si7cAaEA3BzQ
KfUS8xKwsbaoqf36h9csn3eI1j258oXCFiqPl+7NEPh6o/g0024/k+DZHfKMJtS0
nFS5PFFdV4PocJqo07AWpbNGUUGVlt6RydZ0vH+uR3R3dbaSFJi8gphdEJrX33SL
CNqeSLgrygYcRzWbXw8rN9nm5cScfYeWNtjDnnQhFA357+VkktDwWoKy/p9F5ENy
Crz3ND7Rp6RR3fIgXEhgvWrTgbYPWMZSQESAwcUlFJ3Adzt4MPVS9BhC1ySN8CMO
Y66BFyBytwpAQB1cIHUBjSM4Pnbon6NhB7/1Z2XKEfwF6UXqKpTBq4PrcCb24DZO
47OCVd0b+7mekHMzLgDi3jgIyC+67WbbNUJc1Cn+bX0erEkf1gEF6IbHJ9ilMTJR
mebKx6xComnW7cEL1AcAO/z50rTh7Q7tOja/oTu7PFGhKNJ1oG9iOF13IrDiiG+x
NPvA8DigObX24cMSqJ0jv8U9ymle6xCWPysFtMd59vbK1YINa1iNRJ6ls5yiaejf
nL5Fjkc9G4AlqN1Xm1Febj8OEsPN9xzgRr7bAJZ97Kf9CnRNkUAC151PDxHIEibZ
wiEyvH+RqX0cG+Sy8bN9HEEH4zNS/5IHZYw2tDUxyBh62Odw8AtNx23Yn1T/UgPr
IlNH8FZ6RZDISuaYYOIJ3qfC4MTBb+UHlF2hKhDIAPGeJAzNp0s7jmdSeyY6pJGO
6YkQlDLhIB4rpxNFuK9z6cwf05M02XeNPf+GBo6YUZ3eZ/VrgMB8AvkZ3PjTOFBg
9BU+wDRscKTiGlNvC4qARw35CcIGde0f5aqJ6+wK7LSMPrRbnvaNJ5r1WVwJ7SQb
WiOdybJ7G2qeunCm7OCkObTPzd4SIgHgXG+hblHsl9FVwjhhx/EqOXzlSsH2Ia8h
OrSDKfXsd/UhiX64eHGybKZ5nAefKNUp64aoMxCv1g8HjGQIR0EfnSdJZxPSlU9l
nE5KUEfD9qKt8XvFcUgICmyXraGIj1UGTO8DMqmRnLvqhtjBn140Pome9zTmyjQ0
gRQYU3C9ObcQ1qMXPT/Af0+4dVEGFpxQjjoGLn66k9utBRLgF/8N8E6A3Rc/TzWu
HVFBsxwyju6k3K8bCP0JDRNlQgvu8i5GMuS8pXrwcG7vDhYRYKrzvDlMt6EkZ+5B
3n8niKPDTT8lEmSnGYPM083PcZlTVQFYjU/RsGCTyCaXqdtmZ724oo7iyYQzBffS
39KjH8ptJ/964BUyIFGMIYjeaDhduL/DfGk9bmtUU6XgRBJF8S45CRgsaxJprZLz
XSBf4257PXdxFcdSfrzZUV+r4iJTmGU5cmWFXeS6gOgUTlMHU+7HnYhkhJUjfBCP
hJuZerLQ2E4YobrCzPUm/1XAo2gLJgJzUHGMgXFkus6aJWaU0/go0x6qq7Yb6OWV
+sDKWUazvTNTZo9iBQlIG7EkG/BkeICwsELKn+/fYCgDaXVlecgpRwdwmmVD6WSI
tScgZmMKV6OrmUGYHqGejp67mg5j8AT7lIjeyoFRrkAtuuUsS0HnfGUtiO4wMqMM
mAYbr9SP2EK4T4MoLYtrRfytxS4D8C9wpriVYbS67Gg9hln5+mHUJcE/Z24+JCQH
y2syQpZkBMAFwmxBBeAt9cKj2nQ7/JMeJOR+7DDXSkyPKS+m60ZWFD9PTFsKVJpg
gyzQpZSQCJv4II8ELntp2Wu5MalkdCjTIGxlxIZp5pDXxKxq4K46u60Gz9Kj3sP1
XJ5LUSrVMZ7Xli/gWvjRa4avW7fCTt73kKEtUfKucloF2Zz/WqhO6Rx/2xlRXfLH
inlBOs1w3HqaVSrNqyTlIIxkSUIEQGscsFpGolkayD6anTTY7UuZib6pxIhfcAuf
pgutwIgEIi3fWo6TDHQL+Aa8PkbrOUG7H5Ynhya6A4v6pfSLUw7nzIBxLQ/iEQsf
+nM6nV4HgOLchl9a/fUWn1ZQL/DW7nvm3+0nzHG1gMoMChFJK5L+HC8CO2L8Rauy
HU9/PeULP8fM6aA9rGoE9Kr4kE5qS5eKp14cLTiZJWOVYSfgoqPI1MZ4ZbpVn+WK
IfwLMGLQbw284swNAMkEOiFYaLkbt3yvxaxYqCuvm8mC6uhP0JO0asFK+rT3chxR
XgTC6BZCIzKpOH5HVbILbra41PwR5N1H478ULVZXcCE44gjrewgoarOYtMb2KAxq
jWgx1TXbuK8jy2Sz60BAS1H6w6jSBX6KP5JGiKzuli8dIdFEJnHE+jAUDuau2Grt
zFNhGFHYB/+c9VT/+8t1YRuJsSzxu8YQ7HUfzLDQBXv0RXqtF3XwFo+7yOtE/XsI
va85gcW9bSOc/g98mO29uFk9UTu8/Arf/Xqx5fqKvFHWpGrCR8QFYq3FuGSrMfTP
BtX2ikIzSvO2VOn1/YF3EydCeqpWPwo9LOF3nFiRbiq/Cbd8pjTmJ8iIDn+9XCRR
d5/H8x0zQ/kY1HmwqRC5DvVuuFzuo3P7AtLuGgrsnja2AZdf2tCr3qg0m5gOkrzj
36xWr6ybZTTaAvpQ7Mxch5pLK9MIMtATJmZgH+GTKdDM9orEOB1z4Myis2OhzF1n
VHENvdhPiXkQ5pPTrZrIaeV5dQSRT2HUTo0x2gQ6DcSAFy2TAopg8VreUHJxdEXf
odxO7z8GYS7XoPVa97+BY6ulRrBBRlSqNgR4uqQN0l6yjFfI19750We7jmajlqIt
1NQ5pjSPLpPfESfPKLI08qi73BW+lWXmESA1gmwkLoruxecYPah8vCx9IOaRMa9r
NOVk+8/CnYGJdad2GuaEFH4MVG+Igfu+6CW2dCs0zLTFNqOgJekRRa83Goj0fY4O
XOVZhXvHdfZAeg9u07pj4r4DFyAXk5nsmf6JJzhqiZOMJ7eyKcphPFuvAfzSl/5h
vAE/7Zw1CQs4D0PH/5vMVk/9+J8AGxHElMzIeDYD1rRiSUGiCF/ivHPvdbnSt+Zt
dqBOOS1hMInBXsfm8kcdCgqQaO3dXfSc//FQSqrxIfZeXDweFOIHYBgDrNgX+QTn
yXZy6iJCVaYu3kKM+iHn7bX6kt6sBOs2xkjn6c7uOGVGxah2Lo8J40dHmj7IvYle
vAvE51/eo4Rp/GjJKE1x+V5oGMG9tkpbQAKo/exQ8CmVvxHD0S7LnBR7Ma3W67MN
p6vE9NSMvCLiQGBqZkKPyhRdb5kH1v0V4PwN/F9ym0VhiouW94dFlMCsXVY5iKBG
bXLCNylNP7LaOpNpGuOaUyHMVxLBI7vT8vZcWWuv+zrRO7On3+Vwh++Xc7GFjFY5
Whuyt6P3sNYORv3P4XUqY/0D72hZuNEify/KAGtlhFQ3N3jXg1fZB0VhTq8jDLWp
GtHgkeKqANm+lYiEKCPWa4JQT6y1vb/Mw16Uw0Y+I4gHS4hT/me6D+VP9put3XZC
VLR7TbfRjFa3FAsOoIZ2QYUjCZtHa5BI4+eL0BiaiDGWFxjbp8Wgzabp9pFZTsEk
cwtTTaSKY9KlXwIzE/8bSxO0yUSk0c/jHnReH60DT9YifWLWwk8tWxSe+jNfq3UA
MDQ/uCAJ14HqBMwFGUoZWwTeIugPOXFMNLjixwk+woO4vZ3SRNmK0vrI4GJjjY5I
nl8J22GjSXEb/Swh/hFUGxBbtrXe7F4tDzHTuEPoSJhYs/bwaTmItLpoL1sGYpwN
GQC6LdxEd1Crb3EDEoPkZHeke/7bdyG2OOXOKdUMQxTP6gf8mPoPxstVf4aRPlYB
v0dOORL+JLycyiAyFvYrdZrxv9pwVBLCsHftAyEwy5DqeGeyalU+6XLlZpCfBv11
x/7JA3ICiy8tHDUzQAk3EThlsFniFXdtCEYsrE0As1u6HY8f+FcQUlzkT06rczwJ
7B6kQzA6KGVcEAbqEXbhjeWGtzv5JWycJ3DJ8128wY6KLJ3oL1EX1wquAtw2B2oX
ussjEJyu502RxN/KEkA6VEZlfAWvy7yFo65/WeHhNov/pYv5xydLQhfmjxpOxVUf
1EwJxTivDKJ8d4+p/oOURii8BQ5GnPrbX0uTds19nV64U8AItnLWTR0XoqCm4FJR
eKSwN0D7eKKPzmkxIUdPe3rxcyQm/+wsGzyAlsdSnpxtP5P+IWj+gnxvm9Me0f4O
nZHvKTLM2ey7WxWRncbs9v8DbgCu5L0gFwORsbGG/9/2go6NeIdX5DTt2DVS0/6G
2bYXdkXZPi3b+Ng+/7XjZq3lPfcYjpDGQ6AmDOLbIN+YNWcwRdlM62/9ZVoYIV2C
w8sNWS/pYh8+8J0+yEpk65tuJ1MFb0g+0Xf4X/bW8KuT2C+pu6AHVeDKjuLS8OW8
qYpo3VkOvDd2MyE1gd3jCCXDH7dupp5tJDmO45aiy6zN8+T1cw0Xmhz7LZgq4Yyr
pNyeUtKWD6+Ek3ytoFdsIic6Rug5f8STozmMxLKQqhoilYZ5mYF3HDEGjLQBbf0b
R5reDEzc12itWI2Mga2VkBjs/8EWuYlio3r5IPlYtk40+LZMA5mUu/DUPXl4iLLS
QyZX8NgcS+dprIPxgapuypk3B5YQGoXr4w/v+zE+Ijr+Notc/fXHT/ZjKX9DQl8F
Qo4nG56mDrO7XfhOMZu7iHz2XIS+5FVUwWIr1GUA7VYIetEYeERXMmlvtOeemtNP
KAZWYiNdOqm4B0NoQUAs01wU5o9VSZhTnwn8PdbdzKC0t2FQf7DuHUp3Fi6iyGeq
GlE8XmV57TWrOpSTRWoJcw/8lpYzI/a6OQe2mJIkKofNXIra0/t9n11D7xwQNldi
V5o0sHA5qQRXnH3nLoobZnjf5l1RrUkVOrFd1QvifZgmD5Wv0EXzQH6G+WSrE682
mBPkj8PQuvSI4vjrCvASpPcACmcUd6CDxvDLyo1YeadyQxzIiOS4HBKPWB5dPcKd
xjb9Q5oMOWWcis4DUT/FF+KQXQsTL5cGlYk2NHLflXsRrKudqvftb4C8GvBdJpVI
I/lmypmf07nz3RwvTnav7BZl6bxQrRqS6xKGZ0Nauzd7nHwqaYF2GFSfbMHFmZON
n8/uEUQ9Kh8S2K1Ou5AjkZivREokbcSmhliW5tFlQMsnPZgQQ3MvhERdswNBV47/
WjZKgCnPpFQa7zG7eNBOVs2k/HdvQgyIK9zsrUkeU3ne3in+Fa8jrf46T7KpdxIl
uiV87NHhqcRDw8bg9hrQhZ58yPhk0L76jhpiB1/qdNRFCkX2gDjFwEXu/9s2FpJN
Hbh0rqcrS7Q7GU2ZoRK923Z9V7Owz1qeGWhi7vjzGO/z0/AXA9hlIrTnbIZWzUEV
eEP74KIMKv1BHTZaJZHCUMcdzgASLOYw4j6dxXGj938iN+VkiFwN0iXW/BGUw2xq
VlMD7418pYjXoe4XeNcaZmdmmSoDKtXbX+V4JWQSSTLB3v4ez0onck/bvucNhpz+
LF4znK+wgX4l6KQmPvNRQHJjGLB5IRcfYhawwd1JjoYrhBBWbxbH9zIs+L8WWuaZ
9Nd0FmAo4Ezao3e6grs/Rla9PCcDP1f/BI5BZ8pFOZ+uxStesKssbcxU6Gfi18BY
VZ+ROf2vHuftRWJFNiKWxc3/9f7iSX3UKmZt9MOfl3pd58VJyFXhitquGW8L+SC8
R+paMLMuOyLEakSzJh8ZD+vNeFVMFzhDRY5bqgvVnO7JeBGda/GrIep4nkSdTAKp
RJgYdtrUwRwY0tpqeCBL/0ImUtGAjOog6/M6zt6sOjVzCBpylz39txyjfTLVOxP8
NrU5j+eXPBkWu8Wg9F2cR1GBmsoQ3uhNFC7pHOOPtfEMrDh7HSqpEWcNf213ztgw
DX1P3PfhJYOGJudBs5tl4y9xmO0QmxMOz090w0HH8Z9jbGBm1cMdBbBbJ7NRwSny
x5cDW2wK3mTkzbzT7IPTYGQ0Xc48cH+peUUjRYkepOSDFmHT70HFe6WNDkcdA1/9
Daor6A3T4PAjTCiy9vDUZJ3XyUejIsfEnHZ9tE+ED7xU5lCcwu2q9v7iBNieOXWN
zZOPiXPqRzKzEElD1ZKnS84dDK/d3/QbaW2WhN48/T+3XwHRSTQG4raMIVWJi7I6
KzmgT5kku5uePUwczlhNCgQ9dpfpq8J0xqsEEgQlsO5710lwpV4Z8sKHz/Ps4rNM
vbbth6cR/mo7ipe/e5Z8pLcZhS3Pl/l3JP8RXovrG7BTzCSUu6RMA8P5cVei1dZZ
zp5ySITqXOiaTNwJFmI80VEbawHwzmk4utCiJukMHmBy7UGTm27SCyVymYrdwxEo
QnrGuLh0jJEb7e0lfnOH+HCC22H8ouv02wpis2lUl4z3Bf0ib4qm/p9f5RMTKsVw
ZNsx68Z87ElEX1rj9SkETDHvwmbmyvX9fxdFj+78eXiKVBOAg+o1lmVXwExP88mb
rq+LS7RjaZxVNKnOO8P24QEpoK+Fg3CHvBltfmTf4mBTMWxU0jl/d5Nsrh65SLjX
0dUmbpT4kIjrQd3jK3VZUsEtFz0RlHZHyKWAJI9I1C4r/hn8VTuRC52TIS7snCc9
RjDnoK3p0zKaIKOqV8W3g8p6Td67YJaTbLxolky473PH3VD2heV7OMuA53V1YnVN
etHLuLioY3F2twQcvnh/C0Mbdf3PsQLxzia/kkfb9NedSdh+nB9dK3RnZIc+jvzq
Zh7FBwN52n4qalos3+gyCch6PzwC5HNRa5wTXdTOYzSGuBsvxIwijlqb2ZPtSnng
0nop212oyQ1ZyOlGwj3+vFO2wpQ5x1keY8aubfbwZXGQ4FLUA8v5ie6IeutO+652
pDAL5jp9TpU16i+blJ9kVmLQIUFIkqH0IJHPz1vQ45OjuFDLIdTP0GF62HI8mThv
2VNOOAT0L32rq8WuvIwgwdYX439PAiS3PeZnklB7L8vXvB/nQTnIFp4xBzRP+0CO
qs05mxxLUAQxpNjvm04CRqAj1sAy7RWWUshhLUkbG8BVGLnL6yx7pi51FW15lxg6
W47AfeqsKsdLki/PhbTCKp91rwqTq3O/p/02Omtt5SR0HPyphQQ3srvNjQTRMI0Z
hLjKc88N7skwCom2FM1fWrECyBjvmjMmNQodpN2GEKazxY7FVjEiv96pzUmYIEML
IZzH8jo/Cfys587wm0xybRjo78m2N+StTvjT0ksrSsDCTosEniExr/2p4sEwNBuf
8QzFatZMiff9ughQxtc8VnPmOG3T/Rp4I3YPLQq5uaFPiN3lxvdD6NYk5BwdYXAQ
NxOmGGFMhgogBy/n4msvqC9UlYlI9o5kgSOAWAPDP8DFLc0u65IjQYMhHENJ/f4Y
PXKOebsmEouPYvmcx0NCo7qJVfTdCOewD7NBALF88bPo9Do1JNea6M/TPEHLRNaS
R0hPOprF7eFEn9NcX1T+wtAkL30Nzj4O11r47XaiVXn+8AFKol61CuVxF2u+nn0H
JKPkO15c4mJg+/fRBwvwafL522hs+4Jl/fGxWJWGp5Ue6DimkGTHY7Ts0jEXN5Po
MoaBldArSDHi9OuupVQKDqVas8oY4HUAH4s0k3yzKBOfj6sm4FBr361GejyRf/tU
lzhMkAJhP8IkP/Fi7d3sHdU20JjVhEUWimHTniarIvMKGM0xfSDiI/9Ns7UXsaI4
BPUHHZq/R0WaJHd/NJJTlzFasZlZvOLuVdsvqX+nMFeCX2MhDNfnd6lv9hiC3s8W
Vp3nRZagbp32BKJk5jhah7AXiGIYpZoff/c3ko4hUEOikWpspiIV6/BHvSgNCvTl
WVgmsNONRrTl4Rs2db27SQl/n4vPSxC69iPHpyJKyLMvQD0DApYuV1l2RUQFSVVj
DyqzRK7Dh/6f15+wEr2CVPvvv0v2Mtf9sTs+vVQI2ZhfDVIRpyVpovKDh3iXrFT5
zUeRwTZa8WGv+/U8Nw7+2rFRbc4AbUlrYD8lkk6Zx9pWz7VNCoXA3Niuvj2w2i4b
Iwk6zdKcvB3I3Z9kduH5NHLYvEc3MBZz5idsD1sOV2yICceThxYLzJ9b6lZMDp3V
M8kR1t3sfsU0sDJvHH6Z1+FIkigSeYyw/UiyRxaF3FgUna8yiUPWcRFEjRhbw/RS
cyGuxtdyNf8EziQ0LFEowCBCwq/6ZPHCu907/sdW57Vyq1rHJQMjC4cQWGW4nwFM
zAdgJgxHYFZ3EMFKogW2/1etW9x2Gpz81SyTW2XhdqBmvSQPWlY1PRle7P2im4pU
kqmf8r5njruakXSeCwFAB8loOQ+2SEftE1DddqlxftwYy7ZOE6epGNYsILjUivG3
oHxEkJ2DSFQJr/2q5Jv+3Po9qYFKkvg8IEi/YlwTDtq/52bGCaMUY9A7inyivvEv
vINwrkU8QTx2tldWjiOYTOs5Y4OjMTpYkW1SAr60gofMJ5dOsnXU+WtdEzynkday
eP1If6Z9SjnA3q4WiRwPbYnY7ryiN7K8MwPh8XEQ/51KvzIFuyVcklpIegjrTKpU
7FLhklLwKyHofPh9UGqQWMkVdp0ROzrMCABYeegt0zsVb8mngNyyvoOZomNufO5g
SQWIzwGcsyuRFkmBvzpBWgmv8P0AwFp7cpj1m8QcVIoGEbxUh4cS9WubzVBk02Ls
DKj1zyMDZBj6YkDOQ2VvUm+Lb38sSkt6QkXxR9aPtXcySRAOFWoGhXht6MNWoCwZ
D7Wb450X1xxecp2ex5zOtEt/w1g0330Ye+fEMZbzGG/J/21KY01W4X6+O/PlKMEE
zsbCnTgmabVBG8125boS4acXp6h2la15OX1eBM33OcV6l5gETK8nQhemF/QyNkzo
nw7/eSLSVeGFu4d0JGr5BaEBKpMj6z5IdK/3AhIcTHz6qChsMo3MceJAD81W091/
v8qZJTKDAmzHAzKb4zvpV8UeUvk4uL/tjU90HKCQbS3uNnZgGDAJ3FI4eyFctMXV
gflo/9gxiAj7bVyMWsnHi3sm9anjS77AhEAQ80ry6epj+EgFOQ/Kz7bhHzbwCssw
KVukRlA5BRbaah4YYJk8+17AcaADk18I2lw2dxMPzbxWIY32tO+drU+UXOUuKUGg
Qtm3I6co2iRD6hXw2rP2H8k9uciBiZFBrIjuCqIWjIBDS8OefB30GTdqbfKSbE+B
qGdUAwxkECZxupLkml8snRMHSqWhsTv87+jazC2ud7AvNuOw2tp3EvryspakWfVh
M6ouHPDH4nPkQWaQDE5K49pIOHxVElkTttt3suSazNL7GEBzlZZxoMsC9KN81Hp7
T3pxIcfKYHuWe14TEhJRPnZauM9yR5jXBi3MBYqnTgEOCvWoCi1YwuiK8I7eLtXp
qIPoeCCPFQHGLJGnAHwuwFUEHCfFSYueKC07WYZ1VzdWwoEojajhg+/9vgoWJgVn
chySE4zi8mLEYZZEbRCG60W43qvNCqsIC3bD68BYntMkAXDpzDHBHWUHU6TqoAyI
n9+C1x4b3o9z0OGdlErEujPhiUnRKlMs9iCv7CBoVsUlCmEsKc6aU17blTBv/blf
dnF6vp8VKTsxR8tUJrf4WITMWDhJM58G/b6bUOoxXK7L33HKc01tofKdXPvuJ3OO
GNyd/gywWOHn1MqsXOqaULpALcC4Zg8Q31TZjyRsQfchh7WxKM7qYqCkJSI9LMh5
nv8BPpbxnJl8nx5KEyZZTPFekAI7DSRRJE5Vi039M1ryUWIaSEfXJsLt8fAXlTwQ
vt1CSJHOFhgrumJe3CstXY4f/2YTt/0OBhBE5GT6QL+mN6uT4PNO8Kl+ZOGoyswI
AVaj5r5kDh3+qpt8K77sPtlPswoliBO/6fs4vq6VCZeXoE0ASLlReLqSmbdSk4v2
qKtJBIrPGkrEH556VCbUrNO4RZWQkocCeVrB74SV8QPJi55+B6+7oMqZLOacviRf
S+qtBDQM5Fxwc94eNSy4v1V3LhaUhnN/mvKCKQsYT8jYw0MQr753kOiKZKSUtcY5
TEXM2RN7MKq6fzWPcmPdk161Bo0RKLZy7HqLdS/XITqzD4vXc21FgfapbnQsEbVN
MUCRgMGCt3GXbzdfC7smLWMoFA5dLhgRmj3HDPOahM3dhnr+kltZjOC350iN4hlg
LirQE+zt47C67kJVdEwVld2rlW4K+xwD2v9KF7NxyMAn5oB3Xj0MCo03PlmV2APS
bqllEIkWY6CzV7rMyc8jB1WaJyNfBMh5QpJSXUBCuw+xzNs5F83oBfTkI3B3wHXn
skj0yC5ppd/eOpM9A1aWe3YgkEOj/+H5HrQwRb2Al9PX/qDdQXX4VZAZwNOb/n3D
QpHjxycUyqEt3Pkem6dGkkuqJfgFOflYM4Eq0iODK22xvCA/KYRoj3APLThWbX0H
7mZqhkcKaIMeOLSF7cOWN7wTaPbu2nnfVDQngFsXSX6Xw6ckxkXgXihljHA+D0/O
qNcTkxwfxMi1ZCN27x3LtdO1nQkaf0fGDG4dlc4FYWxd9/bLk4jI4yVK7xpLG7Jk
DQ+qf4EgsRzaUFDbtn6OwcC0zE62ceB3DGLPnln4Ujtv1J1dNHpq/QqPNAaubMQE
tpQxAG9DjrHGTbhPEOfq1wVbU4MyZkcC4d07vScxV3IdRUIEUSpEp7rPaBBhRYnt
HrhiAbdbTcU0t7T3AssDF2EXxD7bjUtTL7RKp4zD5OJ07uvvbiwc9ffNE9Qv8kKQ
Ikge/2cxTKJu529LE26P1W1Zyt0UnDDG0TU0DH71SjTauupyiu0Dk0w0vBo9qZLJ
dsFryqbaLOCqg4ArvkcffgHU50MKOwtFXJcF9odbJf/RDidVcxwuEd5I9SDue+Um
vL5as9JJi8/3wBdjVdrK9uDQEFko8LhcSxzm3JG6YDb+TcyOl2w9e1JRsORescW7
Aaz6bTK75iu1z3KSISIVi8aAk+YMjEDSeLOIb+QJaRNvHKpd7KXye28RYAGNJTi5
llotHlgxNfNchF+HeUz2/8KHcRLNoc+ydctDGXSomuRtk+aK1pFMTn5UrfmFFI2y
QJvorqY+1jVQKHBXotYoMVY1sZWoG4MN2Weh3P8BEw9UMTiEtci3CyYS9SUSO31j
S/a+fR4v9PwZcuSZ5gZDWtGHSYkbIMMDlHd8Lz9a6Y01IQZyrsrDLyijPXl0dFwz
D+QFjTu440Khqs4boSNxeAvtKsKe6tG/apgAaSSNE/yQZ15YeGsSb7EnevdKXNRq
u3siRWe42LGKK8/t5DbhAw6tyYa8oWawcg9mN6mRUnvstV0QJ0eyZZ4VujzpgSZL
/EqM40k140Nk8Kh1AeDf2NeE3Flfn+16eFlwCmB9Vx98ezl2nph9iAJU1HravchB
F8o6cfrNf9oMwUnbKdsBIIgBef/NYOD6EUcbZ8Rp84tRO3CHgb93enW4dKjS+krR
ludKaMxedY9RkCEH+CpUXpNF7gxJ4b+LdrPk6ttyr9XZ2ZtQbHYsxcj9RZY1Cyl+
tX6wOhU647GOtuCV4SQfnDGM7lsAXusVhwYrWS4bWjD4TsC/EJvl1Eo8zuTCnVx4
GKVpvhDAWaoRHXOeOT43OK5L+5kdr8kgzvHLVxMln7YV6T6DjgpmcbDiUqkZpehG
hblBcqQ0VaPPRqTIlAp63akVcb4k2fveRd4kr1FdkX34cTPNb99WEv5SasGGkir4
Lp/9XbUfRly6phJdzeLsJHCbj8PlLjJGb/7s3X5jP26PPW1zbfxMjBU6jg5+JUw9
b/3RqoORl5lOMoMIPkCFZNkGejq/zHKNCohDMNvRJB5lORpog3C8OhVQJEuUsrzF
pL1N46+f73a+matA3QBcAfp2fsuPH5OB7xo+S0Xe5PR3WmVuw6Lv9gZea89hciHV
+fVv+TRUpULNMkEVeZfp+ZKqFOb6GwOUcREBOdHNl6gSNI4Etdc/vZMQcs2isfnJ
EQE3KGQOXCc1VG75JPYzDvGXKeQJxN38yvkthexXXp1AhTmbB1pWfxJzUNuLGR49
+EsHSrT4aBRMI//MXGlNCYDfjsexlcDrFFiLgx55AUXWu9r186Q1Ar6kNPyBXdcX
cVbAxTfdYJ8NvtJwZUoseJsJIjIYErZDfRcFckJ48T2nTV5Y8igvyvLJ41pxv4n1
Inb9Q0j02N/RxPbgV7zvXxrVYJ633u7m7dsA/AC3MWaUJX/NYz1Te6IZEL80r3aT
woTINeFDV6oU49YOoWF/A9bj8w4GXbVyY9wSEIWtQ3Evi4yOfRdcV4h0fseiLYt/
EkNf0LuhRD68Eg358zCotsdb4cgdjRaBJK7NNAMjtpy3UOeJ8dZ5fafTxtmYUgB8
8f9IiZjQNaksniqgKo3WzGMy9Crt1KitFXouxdDv6ico+62o9rerr+wfb4hPl6wG
GIjQIGm86Cne/fq+quT1n35ZwWaiCZ5BCfcUJK+PK5Q14AXGzKVfqr6ocHhsQ7N3
yNkYc7D4LkKm89d8dTuGZPC+0J9NI2iHIto2Yo9u+LfIvM2bJt4yIOBgkqoyuKXP
xzmKtwJ7lo4tjVhTSHFsaJ5Cg3VKi84JgiYCjDZbUk1KiwaJNhJ3Boz8XaxOgm7H
nOS8N3W6u8lVeN0oYJuBgCuIm5/fNEegAYWi/rTABEDHcqZyEvs6N1m3tiFLaVpK
3Wre35tCkzD0JhQUQiSZVFQz8C9dAUDj8fKd+y8HUNzV8792VsTr9IV/QhOXh3c6
3FblHlieCEViGou+VUd4CNw+R0aI4vH+XHJSxkVaG/X/mpKvL/cFdEljCLCaYXwi
ZILsuoVA20zsRK6Byme/4UlxoQ49Jxx1v6FxINOstP7cL5g+IGboZEDZ8692PSrq
0PZhMILzrlLpL+SICxWzvIctfEWU8GJnJxXKW9M22VhgBeFC4U5XpUuI3ASwgBIA
n4I7OGjdK5oXHgvAJGksMMFs+yggmV+a5Ht3VgXfTBklUq7rmdB7q8cKuCHs7iu5
VscVhx7DyOX4jVZ3SzufGHhAPkmO8az10xJoFR2lJnUK4+Y4COBGv+nKOO9ZzFNZ
ach4KRXrXET0/O22lUzTnSoiXin8FymAmfPpxTRWKxMjzGZBahGYGYN/ireNhmWU
MzeoPAApYdwEorYubN58kcy69mRq86hJsaF/epxAkGTxBRmK4J3V+GxXY9XBfzNy
K7GrdgcrYxf2x5eI/4mtGaI3Kmc5xHFJUkKkmNawaW2sQFO0ye7QT6rAUJOnYnjY
2r32mBGBfF9SrTVrOL0jD12SB/j7nY3rqCPLvIoiZBmxbOslcp8/MHZ3Ht/E8PsN
GMQ+q3N41xBj4B2DV21Cx4JQ7phJAZiymBT/ldv5oF6Ymfsj4Ocuclwzyw0/Hu+T
dSWKHvxPw3oIz9L2T9fFHDWAArUoS4sOxxwHpupFyXYLOCj9xLkTFJnGkM8nhNcY
iyHw0wR0DqAe6+kn/Dyo0BXyAfpIslL5SfYqA44RxsbxoBo0kJur/PYFtY1EjauZ
z7muqeSEISdZqDza2hXvslKfPD0yrDuR/SS9oG3lTHW2Y2BJsqhRycPKo2JRE0YD
YoiLApBpt0CJRlE+A/Kla7NJcoEr4rlNvHfzNwRhRP9qPs4nBDFQdGmuKgtlSYYm
WbgrKWXSPG7/BTeuG+XGN+/OUbVcjeeZxCrOiBQZBGoLMft6qT6apbI2PFdPJXZT
9HqFLMXbUWGXKNIs5vhCkWuoIq8B8jOccu5bE/xiouBgB6vNTocgYIdvwicI5jR+
MrFxBONzgBhczGhDO2mSF4tTFHiKIgki1BbBh02R34kfjyl7D7o+ST9PZI/BS+jm
Nj6l1+2ik8dx58AoO8OI/OTtWXMKJr9tucYe1M9uUtqLMepfPLeCd3Wu1IzEmK6C
BOW1V4R+AO7x+tgoV00yly453waWApWjuFC2B/4/Kp+2R7b1N/D0C/ewdEQjQRvg
CupG3H3cpMn92RTVqmhRPd+JPTS0wMCOWuomvUhAvJYfOkmSdPX4Ycq41YypfiV/
smBSw64rq/GHnto3OSmR6seGwBGgamyPR9a9qn2z9QfDY2bzCQM80chsNsUDbf+Z
PIRn2mWi9YrWQ9SevAvc6CILOH8aI7LHJkJgJtboDJB85xXqlgKJtV+yqtoPR3p/
nwBO7l4DJ9VioJpFWLy2KfRofKlOyV6CwbXTxa9XbCbzc8wlxPQIShOx3YQvapFD
UnFtfwsKOQIujDAT/2Yrp3+YJD1n+iMp5OLNKuOC4pbwtz9nlW21r7VIf7JS2M9d
iXkwNLTb6GTFvSZBDQzbuqag/CXsLf8+g4cNBejAlrcVjU35pYeWWTrp9ZzMKaEf
VI9bSAqGkaSDWeYgDRHDzHqitWaz4pUppEWrxHrm5jqrvii4AFMbZe8wwcVzqg3M
PtmUuQUE1EYhOZdT+XZpZMqujaUbbEYk0UaEaWY4ac1YxbvFWawOrR4axqOu/C4I
A3qzrr6doEc0YBoxTTY6zztXXxYa1opRUdZHsZu4f4wT6zD2s0WgFuSp4ugWbHWS
x3V9A2XFIdiAdXXB5ox3qcvhiIX2O5QVvxiBNkWhzjBrMTJRSekTDOAwu5aNZRA6
JjUczmWMnf3z0093Aj0VhW8vT4Wd+H1OqYyrZElUM0N5I/EqMW2Y+ze+/PfmYdfc
fRR60561+V+cuyMz90m1Nc/jZZrtU8NJklYFHa4vY5wtDyTFNAH+8e+fD2e8kX12
qBeQnkc7PBDdusScbVoLahTfDToOie0Cti/xUUd/hBstyMW+3We3/8PhMRg9wHIZ
Dbeay0q0o/K7hCjXZwn9YwXtvxN4/0zclBIvDze/lsX2tKUfbW2z+GVrYkZbZWCo
SbDSA2YMQlnznvQqt6CM8OW0tD6IU0Jtir9Eno/Vu1KCCdheKrp/HkSCrEafUpqn
vvOmXWNYU1zB2+MzI5NqKpEgdkjD+S3ERKd8FDS8/neHGNi/aEnPvOuc5mSdf5q7
g52q9aFzPiZW+lOpOCApgnR39QKIJwK3UQ5uwHbqzEmFb8w7S/ss5DFk/UYo34A5
i5qS2iVZ/c9LuhalLe21bNYOEuZmHsyWMrhBWEJPIQW248iZe+2vlfWd7fz7EvH9
qo1XMlzxyi4cQBOhNG0sI/rskJPGFyObBxldl/+UqkxDGZuYfGEXjlJoZC4Zrpxl
hbp+iMlyjJ/QBRTGHXXZkkmnPygkQazopU6250kFvoJHO5xtuvvxoRIIoCSsUFTp
XVQlug2s9enXnNaG5p7VyMuN1VwMIRo+f/GbB30pXqS3Pg6bIBt7QbdsT2DXESWI
E1rF7iUTmm8IRPHCMtG95KgO8/XissiGSHO2TBnDmQ0L91vPbnaZYmXjxR69JkG0
ilVs1EqmfnQNm0L3kMVwc18Y2RYzjiH25n6UGEbP1Fqtzl2phTCQ+LE7B9WChcNY
u432DZ3K5ec264CjD9lsdum20ya2GsvtMrPPrIxSl8M1fUu52jox7LejxniReXpv
IgBmaugPc80TySWmVxhGEaIjqABTYB8IoKdLCD74phVEVDjkdt9bDChWtzjsR67F
1GhSvAKUXSrOfYWj3rUfSuu5Rum1Xyw4Glg3n78iR9OYTiRVULjpXE7hm5WXPCTF
KtW5IQ0OCNcid9vN5aRbl+tNhWrsXJNwcKXZIkskRrz9GtKkgF8a9DTxQLmP3wJW
8Ds2xEjpI6tCJypx5RGxAAB0970Kp0ofzPDZ9j0tIadmiQW9sMj9peigMaRjlqEs
R2PA7spLOSA2v7K8t5vGrG+NzrFff9uhQ4mqZ/uU8NOKSZOB0ewiPU+FJG3O3sYz
hoNBr0YRCN77CrfQUQp88zRywFmCp+GO7zFulYHT3kl04nwHK+OhEddNE7CQURBm
P7HjTPchcgOTeiHqB+90Ex4wql4MHOO6iV0nAqmRNGAlslPOdR21k/Y29UJY9M90
ugRne6+LdDwTGwCLPl+fWVZZ2XCbZNIyCm8h/RCDsv6vIv05VqyrcIaMb/NABbNm
/JLPnTponj5qg/XSFWTC8LaW4+2PHgky98PMgmMbrlx6NkOAhiq2oodyMywXYaha
zBjlGb6E4opOAgyCoUJ3ACzGexDJ8XUy6GpMS22hnWp409ZTu+GLCsjb6lvYOpyt
x8hpsS8T7FSrkVaaX4yxwBIIjbHNiOxiT+XHuvGJGjbQLcei8Y8CLubpte7T0FtA
jvymgN3AvgM5NRFepjyAh0WKkbrs4VsdnB9tfV4z2KoegPPpCNQCCPJU/WZpIv8V
wze3BmRUEH8K84l0mVhw7/WDsEZL/vwE3ktPyyq2FyMXwmp/9wzycMg1cfOD1z8I
D6GkXP9GjGxebhPhbDrCrupqwa5UT2BxFDm2sushbvqWtIvpwjPYERBxZjj1H3Xl
ON8N5iD70mDbQ43zH8z0e7woCDezHrY688QSwh36F48TGJws84S+sO0NUv8EY5pE
JAEUSqDkjjpRt+NVzOQ8kM096kx1ZVKlqkgJ6ndpSdvMSOzrDU9IWWFqlB7BotB+
bCwH2chnVjCQrvF+Npg514q8qgw4ssmGuLbmWt9MKajNa3BbI3lK2j0UoLaxLz2H
CLlIfRcLFPLP0cB+RfKnV5VmFP7aulkQeCGKH4lhNjgINMYeSeG3EtiGSUSBbwnI
g8r/Tdh8mkGZLy7/jU/LJg+60IU6NlGzub9OBVenmKdHNs+62hkYgLWWBec1IQbd
Mu51Wkqnp01iijF8vJVqry3QaFJBnucPk7wwNxFCyzK8Oo38nnpih71A5Lda9COi
T7r8SyoMatCtL7tQdWLY+66JJFMdUfbf2WpeLcSdXl4ksxXOE4m6Dp+BmrsMpoSc
+6hU7VOd7/Ouztnj+uOj7vBMnZCGv7h6GsFu22ydnyZ85NcEvPpjm339d1SwgxCa
XgT/E9psARCe6pSkRXYOCleZpBGY2HM6huP/FPGWbm6sFlIP1T7ZHYTAUndjGoqR
7js+Cb3GqS30D+k721mL2KY5Rn/o9T+6FzDkwpaR4wp2NoC64/inhXmmxZreBd2r
5IfdMSIQNtrMlmMh4P/V66mjwevBM8Cz4D0qnD6FwL5L6+NzMKGPsZCfkB4FrRoz
AnsqR9YKB68B0J1StStyOpUYkxi5ObrNIe+5dikb2RDuQ/EuHBlQfsN8h8fIVhXN
wF8oAY/S5NxwjXeQNmvjxGA5MxTwHat8ottISFOQpoeGejuikgZQRZoBnQx5Pwbl
EiqWV2VUiWxx2rv3jwVG03eEA2dQd3rE2PB6+Sdvz4iJqPsZ4pIzF3xY5CHRl2bx
z0H16wRkM8jMlTm6tsP0Bjg4eI1VKDNeOYSqLP9PdgTdQ4YmCGV+FuahDVDSxw5V
MGWsCreVGB7lSCvlmYaQ+hpvYSYXHiV+ffV/m6FVQYyMDTuddfWeOMp6T6JbLVsD
7akmZl/5ZhzM/Yk6xRWzvfdclfG996s0pUP/7F3ZGIYDThhKIS1D6sjpp6cBQCRw
QCx/m+xPmPJZuWW2YrFYBUGy+HjvM7qp51/L9iMRhQNyY69lhCccBaQhUSgaMCRR
4az3rKbOPvGxQ9BIuDTlKILuh+m1dJLRdvGpQrRt1oUQC8sYt7pcE3CDgjTkVSQh
hkJZday3IH+ipaXbM3qxVL7FRElR1Ve7yST5eYeWCj1dgqA4iKO2scULpWFrEjmc
b0OCPLTFGZ2xGm2iHe9CUfjVG3CcIecjWfCfFIXQiDZTK1UK2uRaJnosnU6+O5Ei
4VhqgUMiU/9oGluRr5OS+tqiJNeK594SuTWrdqSJx9RuqCGmQhU3MatK9wX7OEOS
G+0QnF2O/TwRoyTcSo5FIBQoNuzYjNWa1onUq45D6hgDuXtWHvMZqYF+xVELafAG
17x8k1RqYofu6VbbP2ROtmXKm4Wv/Jss+9sue7xys/eetrQXvddwEN8LIQ/ISWvS
t8qWoJMdSUeO4nZkmsDWBHoOLNt/IubW3Fn2EQXh0Dt7giEHtGXoCA7pr0gEgIrl
DKvKAEJ91yZtcibmpGWWUu6maN2dJC2WLSoZy24n9L8+5H98fBp3Yd16seqlYbkw
qlgNbhheVuQLp/h3e2eTL4TgyxNJug/7c22Kodb4dw3U7YWIikPKu1+zXJr+MuAR
PXgG8w1kRTroSAP9J2zoO6lzid8OdL3m4IvIzknIIie0ranyBkhnRwAk7SPIcpmU
mqHtUhUBGSCxsbg6nmja2lP/qwhZUug7tPfY3550QU70GK3yjQBSBNeXEcJV1Pdc
+rXz1zoADoT55XC+shueOSiJsRP6zTx4GSqdB10NiyaL1RIUFHbSkbuAB4uTG90x
1NJucPz4HzBcytknccqsnkFbdk5/z9Oav/DZ2qIPZfPF8mFGjTYWEbbZhuAugCdP
ECq7ReqNmzwJM/TrpkETEQTl3WCPRLDpSuwjK1E/93cPhWaHq/QUGTVN0woZ6wQX
Eo8sDKGsHifatiAowf6dZHUr7Bkq5CuhdmQ2+PLG8bwWsb4s2aPFVx4v0nvtKTmg
JcLzKshD1SNn4p5DWi5seFF8hDPpWfG6ky+dL/L7hag02xSwkkJOLtNMo7o8m5vm
P69cHlsxH2csHUQsy8rjeWrDiB/goe2upsaFKZo6pfYkPjtmgRaqYMeQEi/qtpIr
SAph0cRNhdZgNs62rtiO9s1pcEDorCaXacQBjW3QXGxF801Nz6fEJ+MzKaDf3/bQ
3Z1HWvlfdm//1O+ZMHw3qrBmCLpwMYWCQclUAuayIRj3Vp08+Dp4/QDwHYgZEgu6
NI5+ord/r3iy36go1qyuJYF0cQCVyCX10kKllgiRreQUuKEcUji+v/XUnDkAPMLQ
nEUEdQYoQsUU+yv+r/CIb/u22QmeL1u66afkay6LaiuEsd1Ou70mqSDmySH0AOwY
lUQ+50ohYdoO3F2Xad4sbZkVTN9ayU2WWt//VedBo+4xqmmaCBuE8WhEcQpn5fFk
KMuh/CxyWCcg33ha9yVAcqJ8g5r5wzdu4OtxZSY8e0wMYDxHlPnt8zWyq7akCHrF
eP7nS1SvZkiXTKzIM2hO7Hu5tj/jpBMnDpBNNTFHbv1MreXLWH5c+6zfgc2T97eq
rSoW1H/U9ze7cOcawpBHEcP5C5T4EAwiJGPXbxj/34OvLgOWsl+eCHjUqvINogYe
s87mWW0rhAzMm1L25sR0JpgEAI3nK+JZP0KYt7QV76WqsVKk3lvVea2j89raxEcp
p4x9O1tSvID7+sB37iPtUuvh5gL9lHED92kQU7ayT7QiFWrQ6xduoDq88v+ND3DZ
p7oG9e5iygP49gKjrbGp2cUy8m0LGKWESsXIMCMbH4LGyk5DUwFAu7x+YnPW118L
wA9vzxwUsYVobINUwTvveMy3gzNrb98Qgs2XuBv9eHt0kQeeJcPWRxJFf9MK+x41
xD/4IpWKD7a9YWgtQ+fSuv4BpxxKdVYurV6MGSv517yh1hkwqi73st4XSpBOWAG2
XG2WJOJ+JSBjdVbkz+5yoUepnTqYtzUw/U9RuRS5bSuW4zxvHC3KaPQpikROOXPs
a3VrB4TJZbSe8MIHdmOH/0irmewfCFYdryMCQw2LBnKSwYkW5TE8P6LkRCeBjNHI
6hIZkbIr+BaklbH94O2WyfWK2icCRXYZoo/ad+HrY+kKDYV3jhdunmyodsh0ade+
kpIAlhUfpOeufLfPRcuPwcBYEcDXHtzg1lLmhWfx1mZbqHizwUG38bQHp9c6qWs6
kr9U86xFRXaJkAz57kMkAYg52SSwTtJE/EVgBoQvIEX2mkUouc+XTvtotz92pi2I
qPzjMJ2o1FrkPFlfwK4zHqXs+i2ld1A6krWWAQR8rqyEodRGmDwRwA88nUiZ2SVC
q0dT3YkwJ5u46jLaDy7hDiG1gjYPqYyZJP/iuOOPR6QvSQYnnplxm/jzIba3Q1Ib
3Rp7C4DW+u/G4A1jcthLHFMsshM67f4aU8qu9SWESXsXFSl7SEejA64j+DR+9Uwd
iSbfYbO+2QoRlaLe7DjX4sLjguKIwLmlLdTH2513IKn3TVL4LzNfoliisWL2qRzg
3UJkofx3v8yKfylbluSa7rzofA0CMt264pvxPGBTu9uqTB6DUKDg5qzGlYT+iWjb
70gLq5c++X0sMTvw4E9+K+z2shr6JC57uAlmz4Uu+8Wmt6uXIUyCskqQ7kv7kcYh
yQZFSk74FzTHko37Bhh4QdB6BPNL/BZ0ssbYZPFWzgBVreiBuWfCGUQhnWFHa/kl
5LeAAywybdNQ4It61gVAEPR7XGawdhDbnhXOoeK0BtrZ+yFbTD66TOpm2gDsVzH+
dS8Ad54JEOZ1+eQry2Y6kdMJwKQ4Yt6WLoPRbEQ7XSBeC6ZDVPZYcCLJWrrpS329
3Q15GHPH3IMySfGSFcbM3nHsA+VF24enalIIMn6P51HkJqmQrDC15+PWNkC6l8bO
5zPP6a/lIZa6wA1OZu3TufCtqRhSOLkNgkg2XrfXieELwwiO5BkIP0ps0OdZTeHZ
1lMHEkhHdtEXSrOS+USJZb6taBV9AiAx316nL1HM22BDqh7GVXhIn3h6I9S9G6Ih
aIzap+Th8GDxam1DdcxfSuqGT4TD5wmcxvbApV0HwR7AUQTGEE13yf9hxFj/znKA
bj4TteVPcaqZWuBDWM82VzTApePxxEiQw0/hGSlDcgMPAuRMv8gVLbKBsgJD78Sa
uhhj4t4CCO2c7VLVup8gCT32Y9XsT6cwtw3XcaVGbJG9iwitrweEvZTj4aGD9qZ+
Mn/W6q3UrqmevEc2g4GMKbADhtXxlDyJ0Fc0e8YoFexYRD3JR73IhhnJ3ahKyM6x
SiYx/RMyAr5k3PiEme1+2YLHgMOCbTpCQkrqNVSapTt8WMQDPZ3vBzw4Xg73C6l+
w8d+vorvgogWYw4cJoEPs0VnpvQWcpxP1a8suuAskjcN4gWuWZwSgIRBLb+jOxUR
J92hjnbNNh15hbz+5dv5FlNOBVqib47xLLvEAjTbbxwABuUKcfR8Omuh01zfS4p6
XRBozhP740Co+oJMulM7BNFjv81Irrc3xrMvdJx4wl0qYrfuLR6VvfF1IIjMCL5a
UGMiv8ABf30HQX4DrK4ztTIRlBmd5ttiZUJZMQphJHRp0wk8y/YXozGnt0KLaQmH
G69uRs93HwJkWqup1y9LvYxjJU/oOOBB46EbH09W33pmm/gz03WEWIorqX9ejb2M
AOMZ0IOHav9DZ0619nIdWmIlB1Z6CRvsd/gUyXiNw2kU8+6/Ax6KodUlvloF/aMp
47+WVubb7/gORv2haB/pHi10tXQpJOWkKZ7r/eAMaWBa353ZjiTgVh/tCEh70Be0
VHjnY7DzQCtwX2EBodt9dpiDp0b++ZI4hJXmWsvI/XWB7KD/mAzKJoa3VcfJs9tL
ItNq6A4ej4MCLjo8+HWob2uky1dqu/EDi8B2ZayeRfak+54YgIny8uRvuJx1kisY
Mf01jWOCgHh1eRWdufPDbcnUQyHybnBhgLG1ZExKIRnP5n94SWm805maZx6FVRa+
`protect END_PROTECTED
