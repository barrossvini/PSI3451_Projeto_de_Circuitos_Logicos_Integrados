`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5a2scul/uAwMVTTOaDzH/etDZdcyZZqC/KNG+qUvNAi6V9lKII2c6OkZz+nFs4qx
WCXWMEUuqWT5oPiR7gzVtVs/gQz51YPUHuYGLLUhmOC6BXO3ERm5PqyWwDa4j2Yc
Itjv3yi3N6hpqIO/xpeGn6jlTaT7Q/I0mCdRdu5Ut3mKzrFwaEcK1Q89eZbQTuuA
enTigIqRCpnv+c9iDZO6CVv0xVEtnf8zqmyiU3GW9wyvr+YTFW4ARKyrIejSdGOl
Emiadc3AUtSgdj6KsGzoqOtKRTZbIG5xAbAB/MH6UhdL9LXUD3GBWz0D4cPE7flY
/JcHsNEAdywApUUV5+6DSsJBqO9gADZLFale6jVTli6xTm5muEJvPMews6BlbeMf
vuqDaYAQxSgshGFieUp0s+cQix9TYO+dIo1UVE6g/F/ne4kNtkxugscxN2BGvxC5
14FWKZZcW2lO4jQVwooYZlAGaT4cHRPXHbw7VxxwhZ2r+pyiOjiXnKGO5URIQxrd
mAO+chSzShg/jb8rquwEZEkec++AKwHDlmetuduiWBs1wD+qmfIT6UF+USwG0861
Xk7OyuPCWMuC05TQhd8XGwZbET4B8W34Cahr0hYu3vIpGHRdvKT85hUHn5P7fqOB
r3ZJxA2tJzvuucr7jnSB4PrSvTtN58SUcXCAexzDGWBBseDEZzqyGr2sI3+Uic2M
d+PpGDeyY5yyZoK35lc8MwtcHZHBhbA5Oruv7j+e2e/jR9h6N8e8DSWJnNmRn+Z5
/KEEiqWY6hxi1nRz/cg+eAOVm+jYoHCBV6ZKMc3+KT8kHkFpPLt8duhilkxOTpXF
Bo+yA1weVfyCrz5Ris1gvofxpQZqcnL5zbOl6mT20Vye28M4o9TEx1a89f0JBT2I
R92EPj3p8A4oIRCE+TSFeCRgP+8GIKrWVlTLtttmzOkmz6qoKlNAD+NHELfBRl8y
TB5+q0leX5zcDKLMHI16ZkTJc+h6wGHPCWn2hUEKiEWvtVKwjvGjflmQ+hLVIcUO
mHNqcvQ8+xudhfRT8BPVzrFl4H6K+55ofLjdILKHlTAUPvo9q3apNAyJ7XCFDz4T
KEYLnHfB+tM2V1bAuA/UrSR7m6cx8QlzzfNZpZvU6pD/exq5kg4/kAQwBYfNN5O7
1f77/SzUMh2hKg/OrhPwNwNHdS8yGcs7ZtsqIbo6anCbHNW+YGnh9uAOOGeTPHHk
is4FSJMVGcKsPhEkdSHVYRyOZJlvFcC7glFKbJPObAhw2fGw7Wsl313PB1rBQ23c
DKv5TI3lw+sHMlcnim+L1UrmMqOjGHIGSMpgQLF2nUewWnJDyXHMkauHVVbjOrvP
ftV+U+zEtn8FojPsUo7E1xDsFYcEya84q4HKe1oyrlPFBebMaJBmElI2iRzAnCit
BjiaJPAk1MYjBNImVNym9c2ZmLx/aeUI6EY/0VI4CSS6kGJHUV/x56YAXkDUL1Rn
8hmpn6tJULFwXkh9JTZGnAl0ugx+DpoHdc5s/1icgJfFkce6psp+nnW+lCoS81kP
0KF2kNr0otfnUBpskCrYarlq2vWqBcsqbUTiJW9KW7Fdibwc9X84icm1h5ipvBTH
gKnJeHy8OzmJ4nIv0byVDXwdjSce9cKB/VOZSsKhWFAQ9PWmR5jDE9rM4strz15+
l3NP7hOVqmoX0pFM07cl8dvxbZHoGpETk6L2DZIX/mjgOFW8hREsev8kHd85oava
whCyAtztv5KfRiKGvN7K8UM6cb5W9wci65I0eyLdWyPf4I4rbesZiarZu/2XuNAI
LFn9nWbndpqX5kHXa3KgToyos4iKhL7PK/J/ClpmdrzTX9BqfWBGikYGJdRIiZmB
kstAEle5dmwiXBNhTguIkTl+mBPTGwE5BURJC4urFze0MpJzKE2DUj4M5lB6G9Rb
sxjJzIyfjMiCiFJHpIYgQa4jdYtHvuqhbOTIGn4uqoBoBetOAcvVHwYdYqpvgB1A
hQ/+6FHKsRvzwBTGNXwNVZmD6RcmsXWfICAbpmztjgk2IzD8Svug5CyoX/1E08+G
UoXuwvSeQJnNXIMZ6sNt3bkVDKKM7DkGSNYC3Ha8DxlrAjEUSL6OpuVT0n/NRYmy
5A7xEnlugzGm3VXz0Ope/7y9MpY0iHAEZcfIPrvYPYZkuYSSZ55oYbnDw9nb0r9t
pIEV/BYVZZIYYaQY365RL6HAfT33gJMV95ACBxEnkT9V7FCOQfIHVKHKDNcqzq5Z
FpVQcZKL4FQD6ivfDc6x5zxvDol2DM4G9LGTswPPQfXlyUdipfFUc517IVlLhzFC
POXjV1Ezy/zMxLRTR3h/CblmR1wEA9SuY6foytuouAM1APh4iAPhdfPOLjGOb5il
/Um5T3qg7qKGPxdI9s/TVrU70qCoLBZmWBN3UNeLk+ulwMQD7fxG0f8MUp0XTnwQ
Qk662F5x17YjonBk/jNuJVhsUONzqPzzYOL1/EGwW0m1QXQ2qIgmX2hWpDCDQzdA
Q+w6QSbPqEAhw5PlU5Hp7zlxcagpAJ5TTUmIy9+7qa12GXOuc/xUVg4P3Fr6zv+A
0xd5uw6WlETD7OaZOnDa/K9RIJz9xYjp19LX7gcXB/w+VDOb6OS0s9FUt9f2ktku
PaQyeSfR1EarUgzh9AvfySJnfMwGYa3rm/RHrm5Tf/o0f0Y345Ld+lRaCmzZ9f5Z
+OSFtoY4/nfnCsv0eYEFloFxs0I3YM5am+41ERQCK28ImWsbhvTgV9y3pcLRzLsB
AkI9IqZCg5KbrX9nFM0kgNSOCpyf1ACpRHq/1H5v9Xigw5rlbLTBRVKKYz/ylYsx
hgow0Vdap9vLbGopPU0ZBof+I+MZjIwC421uJ08ekAFMqY/eQDX95hrmqlJMlzZS
zwZoBl7cG3IKhll/4DygmY+BmZVdQzvnFl6oS8RAEc+keII2Ica2ffHATELFh9gF
MbFQxvthxv8UJ5hNwSL9HnxHD20bW3TvgqODpuKPwBDuQkbfYnXw8Le7/2okV8J0
YvWZFUQ1U79JgOu7rLqXADU4o0N42jYYCUCVpxMV2tZAZVdeUQE7SVEuc9Vka1rN
mRqzCR17Ozbs3XDSye21ETntRzjU7ylV12YML+OkPBWEUcmXzQDedY3MAf6VncU0
Agib+pjnegfzIja+1l1zCXmn7QXRGzqIiiSm6X3ETWVuN+6fM7HvdjZnjCIS07Zv
wJMdPa23ZuHaV7Hr2wgbKcAOzhSYNL9SshfIA+YvzyvqDCnk3MISW1NEQBl1iRBh
AitvN1b3X0IO9WxQ+4SzpD6VIAQqOxSEv2s3TM/2D7uLK4uc/AELPL9Dpoi534xX
A5fvPABQ7ui4ylQ1HOFVV/Cny3UQwDCtxLzNeLozy4PGChfMZxF6MvAgxpcS8DGA
tFywwc+K3j7blGJMZbTdboXP26fDo3b8eCa1+ec4WK5b+uNCh2JkblzNx1LbrCLj
VUbTF2oempMgtGmKDE6PZQxuqND53F7Elr+i68+rpi3AHh0m9PTXT/U+IbNOhusi
ZkKk84+XvnQZGLtmf9/G89NBBVZnM9nybI+wxxcOFc0OChw8Up5zDtZFMIztDVPE
ZE9KvSpvtfail+jhLksM3mZ0xbngjUeVfGZ17+gAp0elk9TglXnd1Q1owIYJbQkl
T8kfpU8Dlr+LexGexwdPe0v+rKVYKbC/0j5iYI39LgEd1wZDZKfoSU37wRy8Ivln
TrzlnelW44wHJXGjHzYBRsj0xd5xSA320B9Vo4AM2vXQ571q1XHJvmu0VmNBidMO
VatLiCrnbOAGAO3+DNbEyZuPirvzgLiwa2iC+riPqGdrZFu41Z79P/N1y/dqHSNQ
JqVgAYVgBTh6V8LGRrHCStLRJWxxqNqRtT9ypFwcwevY9MlMtLS7VyGQfhMbrD1l
K5GTvJoxq/maDl5UxAAZkYR23GJDGkW9BGeGYNOjxJesUPlI9vOKU3SRBeJWVzoq
gHOJfKjWPMTUp7ybQHmInG7wRN+T9EmObkUut4BhlNeKnYGh1P48UXrK3yFK95v5
KlZ1+oBTBecyEk3Zlwla6TkVIctKivRZ0nJaOd1gqKQJ0JVRgNRPkSZX87HjzSxK
Nm3Qy3ABKr7DYJRoI+Fjg9vlmNfe5rQ/2u5Xafb2Mc+vzi8RmByewG/DPuU19vq8
wdjvtdR5v9gooeW7f8vnYQhTEJfM3X8BVan3T69EZ1PPDBcwRRZ67vaHXJqXgVt5
si9D+I2dwiuVIsYNS4/C/dtcOQlWyKJbE4kHBBuN/xZWGOWB5zua/TP77BVK/ycS
2xGxlbuOwd5WUJw0yVjpG/DaHUswfo6DxyIPhD4cgDWYJ2wS9YPvrznv463xXxPy
N6Ozgr3gIIRd0GdQEeJlp9Os7xMPlABsFwyBLEy4lqWyV7VEJF8H4sxkwzs+htXn
olAJlJQSLhnlr8JByI0jhJO6L9JA2IRsDxpcOx2cQQsLQtj10BbDzyVAK7hvxOq3
ithYO7g1mYUPKtyBKh0CXV8IHF+B7r0E+NUlmfFyBZYp9eAwgSlEfTPAoWmsWopn
/BmKyry+7KjUkrjCZJZHklKgAFekI/VhXN9HJurV18JufUMlTFXFvldvq9gYHpaM
`protect END_PROTECTED
