`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6l6Yxb6duQMWUSB+Lhe12p0AP0/sKEeUFwQI7GU1PLhWogTPzUuoTL1P/NBKuvzj
zww0Pa5NYn2py1XgC0nxKjxg8hr0u9O91nYkzEYYhG0rK0WL6Qjt1pCyvnUhjN0E
Mxzl2Yg3WoYC01sp04cGkdR0ha1nrJZupclw2uMlIMqYGwGBWlfTwFzU31SMXuKx
KClz6yLV1YTYrTRo6qYmu80WhtEGmnnN5/I/QLgAhSLcSkSkEQH/FuhrAQrCDcL/
hautRK/85BP1gG8gFMc/gyzLkoDxPjI3eTxMJVXUVUzCxm1CuRb2ekcrdsAOqOj/
W+U4BbcirLUWt/nOWVvQM7EQK8d+wtM1OKw8pgEnIkwyc4CcPlXk8XN3DQKgQ40G
DnKpdzMtypac4IXrpLIsyXELDY79uom9k1xhdUEZjojNfp+avCx2NTtR15aOysnt
93BvbDAXawDOs9TpzTeaVfpFVFfAaksyXcrWJfvv9ZTrc43ktnGVXaDZdwPxuFzp
KqvxCJh2WotdN3yhydBayy7hCzJx1z8qulhlocZhzAAbl0XohF70XBmQ+izZSejM
qvxy0r41hlvVAc0Z8pxenGq7Qu+FfNij/zNY5/DNACXfcR5UEhn6AzBdfE+XuUJF
Vo3DufMZh/jkJxIPAHbtw+ZKU+ItFVOPnXhboZRqTWVymXIVvZjOakM6fG+ZnKxM
/md/Gwo2X2lnuRgqbS9os6qLSDvGbkfZwEgVRzv6Yh8NVO6bEO4ah+YEm7sieh5s
aM694xCQ0IBDH4Su69wnaX6Hfv+ADXrl5HDud6v7H4HaKpVrOgurr97/ckyRYPC+
5vFMN3WQk0Wi7eHtyyP4p9+gOpfjKBBYid/XuHOghdyzp1jgYIwtclTqJWclyyhx
9Ogm6IcrFtv9OlSxMySg0DrIfq8oVkrDf9raKeN02n4XtYjZkC6ljwn60DQRVbgJ
mYKH6Aykf0fMmCLhyJ8U2iuhvYYo5GCs9JdAZUL002Z/5+Ss1FmAU5kvewFUkB+Q
5cDvSYLJO4EC1ve1l4Rk1QLc3dmzmmBGG64aKbKHo14=
`protect END_PROTECTED
