`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
euUaHBVd2+hJ+lmqN/rVWlKkmw9HSpoSpEPPoVx3Q6IzwSe4v/n/vgBGzadHZNz1
qRZTyZYO9jPUgYDv00pGRpXZiMXXVxR/FBCbY+zRWQvtmOfTDPiwK5IqrCvdq7T4
Fpr6w+Kk7nhXFG/4tbAawH7AcONZ3QZm5t/+mVrsXjxgUYXb4rzTby1O4WYmYUfG
qS/WGngOV+WXD18bsrqSp0ajI/FXTcwlrAkDTZNi/Q6P0OPRvV+at52EhxtkHn5t
QmxhJr4o2IzHoWiQxn8sjDK3vF1Di4xV+pNTczPiWp4qY9twH7J3arRI0ZdnndzG
qSco5+hZ2Ztgs71VlXX2qiHYIQIG63mHKBiApcRRA1ca31/9eqV5iUTVZKfWs3tr
m+KLblzhx0bKMNXr5OeY+YcU/ATXoeMBNyoCfxf4pgtxPs/cKdb3xr0rLYRP66Ij
IN9U0MbA2JEVc5gJxzw0+xgtJC+slYX7ZZQzuaToIqlvCfSVT6aY+3IjUjYaIne0
v72MaQFx8pUtzNZt5wixZzBaAEdo2rtLc+cPxdYNWvMA7eQwEqZI/q0rLm70RmX9
ncmeU/JxhXt1Dx733aQxtNig+q3Ir+r8K5gbtEn6Lyn0zPu9+M+mLGteIR9yxwvk
QPYhXyeIa23wndEcG5B33L3XEyyTIqv5QDq4XJzoW+xbVQqDsHwpDfErZz0Cteph
lclgcnKwtS+a4lR485eobzwv/MZNRRl5dhxDHghPx8yhfJ2pJIW7km9DStT2OMcd
6LrkghclsU7mJmOD2ez1OQBxLx309yKU9y7Rpra8vYDAcnZQ/9HbGKhzKcXh6cXg
67UsXzkj4jLErgKwA64sfzpYm0SWeZxHLnuYHLKTWhTDczumUAN3Jx1JRidopvVT
NglSjBsAjVNRQUYeIV5y3TnIRE6gMNS8q/i5vhKXCuZ+7IWFi7/oA/ch9SpO8bYJ
BecLYHObEu8mOYCwMs8+DVfNmoeqmQtm8p2J4XuFBSMWsXXZfQgMP/Hp5nXbbseK
xM39ALdU7GBfZVxrFAkj1fZ0YI3u69ucgETkmD8KFv5q23RBK/gNtHfvNNBBT8wO
7rrbPbMDZUq8CE9fqwt9i5UvpAHUfky8F8EJWKl/0dLwtNTp8qoRyCf5Ld0mbwoG
BirCMQwTHbSYu7MmeOrjJmJx01+Qd7kMpfM+UbnOToMQdc8+bZIN+qQf/q03vIL9
XNmmJ4t2noRPZc7ikrLQtM03ro+thVRsipKKiR1auNHo3DGXz/t7ttfFGJfVj077
kPBi3aRf1kq/OXIETTvB1dfqoQ83fU9SAbrdW3Z9Nbdh9xO6Hw2AaGMByKZ/U7Hg
5rHwG8BrT0f8L89rOUr2wYL53qdGcbGtNait6Q6NGu51IMFfvkj4b+gPj0+2pzPk
p7WZWmDnxV1gsv6f7QIgvVfD6JDmn/KiL33yRQHsIFccZpFDaiAd9IqL1oWc4NOw
FqcmezJtApjVqn+W2FcoJpCf5DK16JHgh7zcJkX6KtSnmuWGLZYWg3zEthbr+xCf
hQZ4quxTbC8DuTk5iBMp44Q5X592AOpCiaYqIHGymBltXKeOss7H79YLOjTH1QC4
tgimd3024UkmooHo1VJn6HjYXxe3REJ5bs/vAi7422ABc5dWsW/70xDj3GTzxnWq
ol0gxYwKiUv1vI+dVhNKJszZHDGh/Igu4vILoegkmlHSFW8uyWYZyhU3v6jsvQBk
hIxsHyU6CMDT5Y7d6VInp9Pt1HzM0uNUIZSAWxE9lA66oLUJKGhJKzpt3axQklCy
`protect END_PROTECTED
