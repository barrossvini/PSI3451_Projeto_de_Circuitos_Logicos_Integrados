`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wjcbr2JTJAbGq636xSXE8cqJSWtp5dw233L7pa8zxHKQ7mVm0Lx1jLT/Egl48Jat
js5P1BJ5XNXDRyhgPgKDNEMfPhqWIx/aDnpHqih5vEdQiyQF6zVMRyqy8UT7Qiw4
r07yyrKlk6+f2p5GinIygYxShOzSmKbhYHw08ioDhPagFSwyTGD4QrpIz0R8mvCB
`protect END_PROTECTED
