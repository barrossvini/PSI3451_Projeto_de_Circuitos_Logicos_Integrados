`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WO3SS6GDlWXH0cpgItH7vkrXCP+RDQ/V+S2x92Bx1HXwDcSwewEx93v+MaGJXyVk
/7yAMy9lrK3ysHgvxEJQcVSsdfIUb1bEfLHMXziOs43zoi6UJQ0Ks+FpOI6LX2Re
3a7p8jsePb4elRjEzewY1oz/cEo/Wg1nYw4S+E0p5tu21hY9SQJ1HLpQOTIKmgul
C+fgk2Db+8RMlhwuxYh5HxYjrp6JjA+3ySdAFnOZFGeFPlArGreMcnaogdYyEqWw
epRIOfgUcfvi5oaVAWI216orzAbsWIlgNs5fssLQFIIaUivDTMljHgmgdZroqxqY
PfViLAOk45nH7PArvzjmpgUPV+Ng6Fk0nwUi4pdGc7CKlee4FKTG2U77HzIEuwmo
fh9XWeGsUm0eJg7AE+smAOdA2xc4Sr4YS6rvy/E1DS8qT5XuuI/0e2UICdU4Z911
`protect END_PROTECTED
