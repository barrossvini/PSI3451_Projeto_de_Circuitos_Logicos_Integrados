`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BgoQsRQqwaHVdRSEliWB5BBDEaNcSDY3ofBr8/ln8dFOxtAQI71J89YXhvwFcJTC
GHrECIVmkqIAcw/FhfdmksFXhB22qM/uvnFT7Q0jSx4bZRyMgYJJW3N4EqNtfAdx
RrMO2obLBRRiGehVSdAkBumcPYkTOMRVGUtk+F0lJzPI+gs+LQkZkJhMU+4Q4AE7
QaZWeWrNSGEKgEIWI1g2YjTacKMBgmZ/bbpBNsKl+xpBOd0T09b6UduYhAH6wWLd
4N6GJa8s9nXPjyHtKifVUeOXt5vDT2bIK6LucfyFFqnAawG2zLLs1aJTy1lsPCpG
6a0GA/agkZXBIam1ocuUR3VshDmwSQaJYGLfWrY+SY4CUXuhR0cNpT3Zl2odFHGu
/Mi+ExHAbsMyM6FbAAVVisoZhzGEDTFrd/sxpKZs2Eh8OSOjG2Dg15obPr7m9sho
VHnKtm0eC8Cn4n6eUIt+mG8h+os6HKo2HZlZl7bMDNp3jeaoj/4dau6U5Nbk3JOy
VNv10cSbs+SaUjY52FvUG2ZjnFbWZZkVK1RUp8iGUbtr/2k/ZhdL0KqXvZXjxLAA
2VbmuzzuwA65zP6b/rDB6GwYK976v0x5ZWPlI0Kvcd5318xfTf6DXfPl//+7D4ON
3oFUVM49TdabL+g8LZJXDYZHjeSgQHt9R8bh3fjJfUS2SkAu7P8yle0q6Jy7ZbE+
SjtDWAWHlVnot8fxvgFS66GCkFj0K+l+QuZNB/fTI7QA841Qr8dteo1EQHdFF0Yp
75z7nt50pBsKTOgrPUoqdKGBRGjl4zlLGbqGqZZc8f+RLwQifaG0d+RswxlPycdP
YcdMeTtIbJ1zluKpFhFyJAcZVRic2phu93na1LWD75TWpc56k3VglTHG0flXbwaR
MJLgYe1wCuMkn8VZmLcM3jaDfdWt2P79e7eM9f6/Gy68IWJHWLVcVYOHLZxI64Ww
NxCm7/zaaxaYovDjpIdZvKwKm7sI7JjK5tZdYZaq1OkzIFpz7l6n2TupVGCCdo+H
gxvuyA9YC/I7R82fiAq7dpkOaAEgFj7eljcOMe2Md4g2OfaPNXYxCNYfeqRlVq4n
E9Zhub7MhLD2TPsev9pW/I7X2A11N/qmzAB7qy6pocEH93FHK0iQ4ezbg1zCuBmy
8dUrIsGTBk9es15qRy2ptOWvH8gXCgIx22p7nuCv0J9XEbVrr7kFiWZ9pmV5sNT6
0xVHif6zLMCvab+HANqLusQF0/Zc3KQN5WwZ4yjUt4ywttjTOV1yPbdQuziaQFhM
iNwldQ/ey2hR4OuJXgVWmecxbMjPz+ZOa95oC5idgZWXcZ6OM2Qumw2zSI7bw8mx
AcJAtzLVourfe8T6cL+lnIRThr0O/cVwlFavy2bIFa/evJESKCTg4JbWFXuSE6NW
7vjG/2zUpmBzsDzwM8aMojJFiLusg8QtLNFO2bxwcWYASefyXQR/4FQhTzoOJ5g3
mKpYbBoR5uOdbZ6ZH0YDTp9e/EQf53u8xB+w3cqJkj+fPp80lL4mo8wAqdFfsmgY
SMc07v4wBI3Hpx8Dk3ir+ZtADdtA+iRHlNB/mYAy7Gs=
`protect END_PROTECTED
