`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J2EYt/sOfe9vFfVc1WIOAbT0ec3skORi2Yqfp6zcUjABQ9TwrB1EC7+sXIV7Kbgb
9rX8stuRWJenWb7UTLmW1GuFjA1/+PPAOMTiIpQVaKR4whtORr5Ta8x3A/WWpD5C
NgOzI1Ndo+FFr0AZnA6wiXj4MBeO3eudhquEyOIk3bZ92tIzXY8LuyTYg35fH5xs
qEXfE/PZSLzbYbeQi0t4gowBZuDOUtZI8n9nNPG871V3e+UoRS0ZqSZIZsLiTFLQ
5tCie4B2/rqLZG6NvmYq5ZICaouLcnNjFbixmWYcxgxetisWTbh8Yz4d7XZCO/xI
++uDf825FyDH6V9LfNjb3SW6ciLM6ocPet7lBTSAc2KQnxYYKUnvaL5Vqx528AfH
KkOrpujjg+058WndYFkEQAD/MJzIFETyPbDhtWFrPKHbO3seb1PMxksUIgHnBwTm
zcPmroBBVgSmkWCl7yvzqg0WsViZREmzaQrE6SCEGpCDVoxu9ZA/qMrgFAeU5szX
kA6oy6pbz/YN2tTI9vTMlXSvoW/8+lqnUi9O6bt4MhjP2aR6oIalT1T3sQsYtmEx
vMiJl3Qhkd8jcEN+T+Ypr5fGlw09Sl2DqJlIIadLHztczGS8N1hKt+YOT9g3tFx3
yMcfpF4EwZoW/c7FlxTZHUDVMwQqAHYsgnAMeIhWRefWx64uKxlfsm4kl8zHFpAr
PJ9Dhq895paH+5znow/1IPO52J+4QhrYvOZ94xF+arJ+oU6eMKziOxAd6jwoh5hj
7DBsZlib/Gj1qhdilOPN5w==
`protect END_PROTECTED
