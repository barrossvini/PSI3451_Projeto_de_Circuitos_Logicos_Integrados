`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LvL1bN9nzaYqCyPhxQq/R9gyiSUkBJJ/25fn2563+Qo9+8LolUvuzkzDOPQcTHPF
Li9HTk8osoxRaTm4Ew45KiQP8MjtcPbirs9LRQ6OcfOB0uMtrdQqLERUug5JyL4y
QA2oT5PH8J62fxqgSFusidSYHYOSeoI+aBvUgzZC2Gpyow4UBcqvBsplnDIDgGyk
dwbKy4wwxDZJf3T9F7piTezigHHFjWeVC2pJuQ0eEJ4JhLydC3UR8vZguqAPmlfW
W7LpumeeUoocJsBelhPzsCnv+F14yCtSlf9oub10hPqM8XwDqaZBN0zAFKZtcyjG
jRpXOi5jXUYZm4aQMP932SmftKk72JLn/PxfP9q4qCaVjkCjkx3qC3+Xmg55D1Cx
MMF2s/ypwZ22TdEhHZvDLlNGPmOVzcbcvHcjhmfhQO0WPcCJBtMqlSlD5ltim075
ewTXmifjjo8ixcpPtHfJduWhcnesR7Eeq116T5kVefJPo3GPCWJ9Wh1nWi1lB/Vd
aM+7iXI8m/8sedl9lAdS8He+/Tcg1+bUdH3dJfQLNCWZPdAG5QeP0Zk3DXn+/ZP1
RD0IanbINh334wlkC3MY2vKv1exgl7SBrs5So5GuEys/3RnoiNtazFMzLptdIN/E
ocnzWfACrXnldIXQocwiLrwYxQz9kQltAR9X5oRLELQeJbvymL/lAVxTlGYS60ia
4DsFR4FBtHK/X1UijVBWAV+yFCX0a64jHvH7ZOVLGMXmiyL1v8drMUDc2eZCeCEd
183300jCZ9G8pnXlAjyQoxNA/HSi92Y0JWlroivNqsorNC2bZK/ExvzoVlwYt5oP
EkjclcfKwbBQYBQf7gz+uqyw70y1iOMMRN4f/Ov7Ndzd7Tv+s9xUKBr1pn+8iY5s
`protect END_PROTECTED
