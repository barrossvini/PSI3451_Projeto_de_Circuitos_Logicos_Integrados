`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ma8XPqdcWpRaYXtwRRKg7F6u4dzdD9KeHiZfLvFDrTiAmG2mYD+mmxAN2gFavdaR
yZP1R4TSy/D9+YASF4lyHv42LBlmwSY3bjtA28SO9mckJTbH61vzUeK01X2mN6Qb
6u1hLcorHsWX9zhHJz7vPZnXXZ0fY3hh9eslsDqCtHf/It9PA5KyvSTIsYChTeAt
1of3H59JD0Qbbni3e+5/xc7Hqs7SXr0RdkrZB9XRQjXvwjEiDW70xTNsBLQ9ZY+0
r7Oil1RDmN0CkXyCGK7sQRdXVf9RZmTztwQtFF4nK8x2UxGeb7m1Auz8eT+JxqRU
+A2xqhOOYwJh2XQJyKM40PdTf5JrX+91tAANoB/Fqp6SXzGZQ9UT1slMT/FRyaby
sqAiICQPWNB4ResX4HhxoaYUjJudltQgapW/KxJ09ze/BMZ6e6M1SyACbsVBckBo
ha1dE9SG4BckIw7MKitWofKTYC9/30vl2YuZYp/OaV5YXZLu1ED19FCpg2F6boa2
usTz5ebaZXVyfMEvmN4RNTj8kDvq12jHRxF4b6gDBrSZKTcco7bUfVNcfHrQCr51
MzYxzQ8O+ukW5JHPkWzE0IBsvJ4OUEVehFlpESNLp/gcseMvW4YvjjYoQkT0XGgs
1wEiIyD/sjxOB25s/ROD39+EocSQPEHMGRZP1Aftrhi0+3We1mOtdBpF+vaMF5D3
VXbg0CjHfWfNkH8lgc3/5oilwYwVPpVrIpd9lXbkg1/qssjnhSVGAPhlQtdCIFma
uMb3Cl1HbJy0DUK68O9npJT4mBWhxkElwLCPpbRobXVvxNRxePVbRSFzjwOrC4Jo
R3h37ZBjWYLxISCsf8NObSclf2MK8lidV3FlrJFlTnxTATMAYecQyQyIZTrtddaI
KELKygMlJ5a/hghe8ZzjxSw1j0xMAlWZ9+ZrR2QyxImA3sgme5UfO8n6ICMXFb1o
qmUsXAebOQ3MKZMQGuqbvMXZe9X1K+gZ9lAdctolXyO8EPbmLmOiqUJxO8iBSuwK
JeeM54nRz9WIpr05JwcbHOkrW4aJEaQFd/nKBlNpdXBYbC7mJyGoN3EKBfEfzU44
KE7fIOkivZCJHRPUPzKUB5w2cGTnDnGOPiZ0BWbjbakjAitJyEN7yVoXnmFqyj7f
mO/gMBs5s17KXmQOSuSQvN9bATvNWhQ0Zrm7U6Bz88JzxXoK7t6gQli1Egs7CD46
tjupZQFy5kjtG3H72duiv2dQmWap6QWBxH8dHfyqd+la55j5kbmPh5k5floEHHzz
0zywv4jcuaY1p6PGHWJInyJ4oI33WbXTuBr/bfonHLCno7RfwAj/1+vhqSEHb7Gl
AqIkHcTSpliwGgmvbFIQaufFwuJ4vrAR6zmGwNNJSQrv98XfaWpkjWHDLCnHcWhE
KfWYcav/NPF7QCNCG6g3Flj4ami0dS93AsAPM/Noy51KzfuiMc0gLSQCkwqQIqNk
rZCgFfTbNcqLt9DD/U5BzzeFLUMWhe6cOo2kNBWDG+4ho3XMiULQX3a1LjMjzf9Z
hjnglCmX3Apof66DaIGw66aOmQr8ssZ5iaW33Ykfx+GPTQgSmoBx0QJ/XsALX00J
txQm1POAHU8Us9LptARmviJ2+IXRKv2EIE9xghVg6wg=
`protect END_PROTECTED
