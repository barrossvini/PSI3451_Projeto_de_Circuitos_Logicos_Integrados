`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
txJlGSN2oSqYKYMLTeHvcaoDlemEiZoAKIBCGj66jr4RhGS1FAooGK7kaWpbD6js
5TcGE+9USFmX14JClay7qLjXpAuq4v+8bLhf8+KjheiiWvGWOehdDE21JhMWZGAk
33mN+jS+7TyRaJHxnjO5hJV0kySuiNVAgK0RZ9wX93zmTw85DjnjJyztohTBv22A
ki8yYb49kTkUnddwlW1LV2kwD3EQft/ZDrj/skhTZsrQAhmhTVtZUQgR8FjoVm6Y
dS4XTIfpY6sy0HCrfdeDsjHb3CpZNwmEw1BHCHXkqAvBaCOOzBUxxX8XURCREoGM
n1ahTMclkK65pfsgZyXA+7aiSJP82B9FYMU93i5QAHebfct0ciBoVlAMx4AE3NEa
RDAFW16Q44GniV0HHLcfRaGYdmJar3ouRIItDJdkPBdgRj7MbTIOZLSJvrpvIGM2
p4SAe/OMiszRk0ECQI2cHYYyqxJtNa6izAEN2sqmn65783A4AhvrAzFG5OZS3s1Y
YELfx1piiuXFPK2up3jZmeGGlLwewzaGkmXSAV/LEnTgJ6UjIuebRl2Y6iX2J8dI
LPBVwWsyR1CM9gr4Bghs478pMmp1UNqCEqWgu3JsmSljWvdW6y/xN3P17XqPyWSX
RH41hdg9OdlO7Tev+frWdP3zYw6o79d4SMjXrdXeNtpozak2SsU9GpxYTuORYuL2
DZi0ceuGqVFrQKs1b/+N0fTR08Lg0u9Y+GOWtOLFkezsNiVH31FuGUkgsOc8hCnm
xdMcCaFl969+8Vc/COq6wUNn5E6LCUA2KTSAJMiRpLXvfOtsuPwuxpwjZqQrbRnW
fxCBrrnApdhT90/u4HJr97Bh+qPn371At0xF72EtpiM=
`protect END_PROTECTED
