`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdwZx2WaB5y4VdqE4lXhdnFB5t9m4jFOp2kZuV47Rq/TCkD3iweC1alVRqc6G3RP
TTZx6nU7negPiP6lckWiXEIfbv2+bkk+u1Lp3GM7XPm5Xlf+itoUJMqKVacDrgbR
wbKm+F9pO1TkOg5AsLITTp8HuwTUD5w72jgn48gstWpT7BHBmcQRQhuYLLT8IRBn
CFoolZL4G4arBpXpWPwNngaSVbuMiKJmIC6BJdkL1fun3jugDHInmG3jw4dHH9Pz
n5Sxr6psdxwSekT63yqXlaFQv8iUfTD3Va9zk2wTWQYmmlC68vn65b1xY0LL07cm
jtVVyBjp4sGtsuJhkc+0RAJW5tlpi02256mUVKgPefiXVJEWOSVHNMJic7n8bDNj
AFUt86McsM/QMyxp1K9jKHdSacjEW9NqbEiS3SZb5vnzkdgJfWSKuLgtBOKfwpjU
ezzwAU+VtDfmKY1zJjoeNJ2cJH5LlGyU1AFAQMkNx/g+TMm3eSmR6riZuDiXB2xS
s/M1sm0uFBJXHb9zMu93eat1XZqxst0ERVuGjxTmjsBNDOplm0havMdJWDW9+1uz
uEjwX9jzVCR0VTVRIIRyk7AKV4yAUdNC5AMuacXpuaCpGZtZunq82B3CWVOz1w2W
En/XTsZL9HM4vcnMTpG8WtxjxA1LyBxuACC0CGV49nJm64sJ8gRw9alewaNSil8I
cqKUiJOSilQ7nPIC7vfdqS27236nGnGPUZ/mSal6poc=
`protect END_PROTECTED
