`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9XM3YYWefAJCrvZ+1HIxWTrW/EClwKhh3025bXllHl++KrbOU7NUWVIjKb9BGky
X9cTTGB4Q3mggUjFw2PXX1l/QUf5qjzPDGurri4HEbLwRv6t/P6o1Q9BLkmrDOex
gaM7PS5930iuV3Tt/yL30+KDzTN8A5irlTgjhUyNU4RrkRunMTJTdH9giJREvP7e
YUWy3j1VTKgvnqnGzv3jbBwrkGYYUGUo/svO0uuGj5GfNQUTIyN7MxJnMJ5TIRtz
X9yKqz4V7YMbdlV0Kzk2t8gMvDQYAUbShIGVumNLvHuk/Azz0moYFdKyA8WH7u66
TZlO1LauWxCbtVugyUuUJjM+wkZrkfenwmkVz8wjmiB0LnFb1V5ZqYr/mHujw2Z/
RBhevPnGh68y9AYUOlD8RzBf9cADQjMnXW0iLaizOyV5zCQ2KILWt6w8Tq82PkG1
oX/zhffxNPa4wlmRJPMSCpiPmTHdta3KTQMMg5cYzgj3+HOQFZ//l9cJixK69M6w
UBnuLJ4Bwr3o+icLPUrWhwAVWmx8ulaLtBROYJAVggowUGrnPSYPB6zl/ORkGkpT
h2kOCbpnQbmOujBTCG0UH0dKNtH0XGrKHvbcoA3zIx53+gyEQXB1bNb9oc0qDwfz
7SXtVRUZ3tOfJN4SKVCdSTR97pH3f1AvwjvfV0FokmZ7pl7PkpNwv8aydLODe7fW
sImwKjxwf6T5VA5Wt5uQs66YcWSP+5auSuzLt6g6NQjrMvhyyTTxoDJLyPtQKUSY
LVeKyb71S8fRHALgYvU/Q8BVIqZi90SgQ61oYXNodqBCrNFBAROSnOeK8nkvpglt
XZ3uKzpQGzDA1ExRQaC0dw==
`protect END_PROTECTED
