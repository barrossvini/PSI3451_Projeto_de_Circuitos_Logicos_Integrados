`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hTUkh5Fsx0hxTVpXtbAvsR/OBENHLOXbw+HHWUdlzoyGXkU80sj3xmrGTPS8kQBa
W42B98srrZPl/G/LcB0w/uK4C7A2jJqsLdJ4CZpezjEdrYGNXqyrdWH6sHhwIze1
q9WOjgp9TEQa3qFxVVEGZ8WWmcp2l7crxqAZT00TZE3uaZUG3H2Sx44noQDK61NS
PUyBsfXu8XXvjRWbuCBZRmauP+dBZvbvn7RoV2icXQoxsu3mhgXl1+l2wsk79IUS
9Dz1doakaocvwr/UUF6gzhxis78k12vRU9q8rp1cBXKqim/E9VDtrF7I5+BWcZnN
7/o23/4lGPN6s95GmWMWoYzOmbPQnlae7T221EkSmivJd/q8RCerbOZaq1TSeA39
9I7clss81bZu8geDZ0a+EGHotchKKCXZhqMXCP/GQ68Ww8eGcuKsVe8Epukq+PSM
CSnaMUnr8jble6zg1HonIRakbGhxWV/jJwsi6qHDu70yqNJH1aObOC9NMMO6FfvO
Qeou+ah5pLRJi2ckSIx7kprqHcV/nOuEzaUXHlyeOFXPJnDtycuWFFjzC+ZKUyLT
zV5PinlBFl/mknjYhF3CURq3tbD3WlZ21qF5IEBjE85TXCP5SJnXMqUz9OaJMvre
uSqnAhCiid9DcSAR988fCc34Ygm6rMlr+q6P++zeRYV9q6nANf2kl/2y3E7/ItvY
I5Lb/60Htqm3D7EXMqkstOZhS1rk6y4D8u4KWCsou4Gk5W6grbh6ggGPLZBy8dpo
aQfWJNmM0ESXq8azCehbsNznj/83wMdJN5SGy95HobezS4KzExc2CkHmJFQE+Dxe
8CrLBEQkRW+1R0/Zm1vwYrI1Gww0peh2Y4y6dB3rJ8ER0XVhq55cSqkm6Jkb4H+M
twvWAyQTKq0q5YTX7gYEl3R1/qHAUvQ2/3IC+94Xv5cTFDGUrjOFneMBK1VTn6Ui
WrTv/nZdxpB3CBvZL6uPef8+3Fq8UafnCZ/cUVAN88R+K6GXiM9SxGLvVh2ZxHmG
hVuGT55mIJY0k7aa1KRWmAVtkZ4eXnsO+vnThoBt/TtxRCDuBrCZzddVjwur2u2z
S+Zl6jV6QdVdvK9MVEpatEWXVMFrUvH1MmbPDQI65lZ7cHRVPahPj5ytc2rHV9kl
rc1sAIUZw1q7q9G5pZWFF9Ruer9J4/ROpG1xQyeDSeF27fPbRL/NadjT6QCFxxm7
fNlEsArMA0FNaSPEQp9T0L7knLu0pRGR8nVE4A6GC8oaMZmw1Tav+Ve8gi62v0Go
MJTuL8lNbmES6L4pCUCH8MqQBH5qIgqC5nEx8ges/VMfcJO7eE1O1J9CWuxj1ran
oVb3YFzQcCp8LadT1RQOpmeRJs1I3M795D6xvEdJu/S1+37tVBEUCOO9AESgU5Yt
pNTTMiaWyBkHrJbdtTwG5yXvZB/TZBbW5uxB3XkOpKmwq6csBpCK3I7KToSmDqUe
3b73tsH4mCBHLK1RAyYdwvxOviVtbsw9ifojBQxU+wjBWitCqVMZCHxpp2s+eFmt
J2SuyMyTgoa4YtNWPLiW+my1Slp5u3cU9lw0goxeMRhHYg6YE0GsIxsrozDaDkSW
UU5tUg605o40nacFIZo0KhGvZvw13/upPtKd0ztBa3RtBvsd1pdNKeyvnpCl8Dr6
QQJn5Dn4GDImbwopoYRH5nqmwkxhC2Sv9obUy2uHXCiHerJkw0Tc+gSG0++tzzQP
rqte0bSe31YTe9a0OTXqSOr1SNPK4+5SoVZWsXMdwmiTgtSKQxp31sg2UFmAZNMt
bW26450ED11wiPg2b9iJSr2Yue+ufNjKEK1vZzDN4MvFKAhIkeUmVT1+kvAXb76T
1qQ/NhLUMmEJWHSGO1huV76N7mDLbsxRyhARyaV3VAR8Za/1uTVs+55XmFW9W4br
8uRLy9R6iheI505Y8hJG82hjLFsm3htpHmBi4Qpo1mIo4ljciquU+KdF+Z4+LRHo
OS4iQrUNjNtSUFD8l4SmhYbhaUE7wLNL+F++8Ur6/ruUHv11xCgQ1xdDPxxdSx7G
mL7HpgZuc1Hf6l+U3IUPALmwaOzLNCnv7Fw0He9vCl7Wls9fGGydOXNU1EGrc44R
f5z0Sockzw96dBnhUhnsuC5CvfhGKIQNMD252yOXlmFhYSFGgxq95PQAfnfaE14m
2nofBUscjnyrRHGChU9AGDNjYlag6Iiw8kfNc6HmmJ2t87OTVFiRdeCfZyQx6w+g
rMXdAbVVI3OA3WQ94uOtL+sAw8zC0ljBfa9ISPFkdsvcL5N18+kQm55OjuG0wIMJ
/LbGmPnowFv0VSymyu1uoOINO1oc/K9mUc6OYqja4CV9cSgSmodudxOkOsHVimkb
kZ7uG2dHtYS4I+RO+7AgfMiQN/FI9GLwlxdNANvcxx/LF92uISOb1xqAJ7zTlgP6
rvDWQZNSzGvUUYTwRlZQwJchbLYvfmopSZelJEqZVIArE9ni+7aJW97YE8ugYlqE
Yhg4+ZdDpHXKnjWs7j844WF9biJTATCAaBK8qr6qWtJN/tzS9gJ2ifpzRUI4J4oy
vVyY9jDbMAAHl7/bz61eLqL+tiAQB0DtiZtg1Wu3qZWnim6PyiejIVxUxqGGB0mt
ukg1qboF9C3JYMQAeaNxCs2v6bY2TGSJmrY16wTcuKAlX1ZnbwcUHBORUDUq+mgb
STGvgyQ9uguIUuXxe28416mQi7LUhyywwnbh2D4fF9dNDr7GTQJB/uRccb3jyRXu
3XHU4DF24wzFpbOK+cCHaJKzkGTAd/wiiz5zTR4oa5kXDsfxXSCXLwHq2s8q+xHz
elJP72pELT76RLHx+ezUnPX52l+Y65ci6dQn16jeh01eryTNnpGCtwU3WlX5ldII
0h8+2s/h0DiEmzdL+u8hjCXbaYM9q6RNh9HKY2ZIX2Z7O82bG1Z6U2V+ZndIrJh4
DNhABqTf3VHtR3OUoDENQ1V0/Oacm88KKW432VH4jV76GlGHejLUCnRgeeieH+cl
zZJ9aFQOfWdKdqY3K+VGBImcycJ66f3cvBlw/gkYJV5zb4c1s7iiiPhedSqQTHBR
6DVBWhrlYioba1UXeTJlTriZH9GeF+Kb0u6WBLs90KKj7AKZMcwv4L9yBRb20c3N
dY/OoijcoxynXyPsRIHGtUtm0jgc7NcwpnqpzCx+4+ZORb3tzlK95tUHFiWkRNrx
ec3G2n2FU5KM6tV7FvVks+JT1sKJsccZcZgN6vKQ3ArZ2+2fk+/H6gmeSt5uD7Cj
iirD0SXEqY68hywFiu78yJBr34oujQuf/Lrl9S6Nv/jN9tgKvZmVpcnBrFGENWly
+pAUB7bPP8x6qMQQuJwmfctsK/prZYrvKxk+VXzXQfUL9jQXt51ONdKtHK2+MEtI
nuQn0ALl0fJ2yu4m9wmVCb5TOysOb6b8M3YSWWEbCOdqhNvfMRkq8AU67YJsJZgN
ZcWv+Bpv2ZC9MGq5MWOOG1bBgL3nIfQZAuUm597aA++k6s4aTSON4TsGYhrcLdfF
ZyctwbBuaoJ/dkt8V4DXllhGqX2BwdzFckUJHOTw1uZIq/uOatG3Rx60vrR3OS/q
jlmISVJuCwMxFHK0ZklIgzaQzE4kYHtnEZZbEnN1CYN2lAUbMqt8mvr/74CQ9crY
QZDJUn0njxktUAiKMe4PnLh6+M4uSCGEYx9eNuy/bRp+QfdiQeHF0J/nwDoGDjFx
eoWbwdOxBGA8onPmCkBd9377OPAyF6OlwCtki8OaGky+0i6tATDCx3eYYEP/5KRm
M5IRVefdPMr7JEGBqMmnkIDCX7qmpvdK7GEww86IQAqZiu5TM/yqWX3JYQ0OMF+6
MyUCAIIGi39zdvyLbpRfQu+hB41kyEsPwM2JRsnZKqc3b4RL4I5lZ92JdnrCy2c3
rVLKf0q3ktpQvLPAAGDsSs3gMNq1TKATlD3BTxtGcjVPlMA/ABpxuTaAY/sRYA14
iTxDDnnYzyJX8vsJDjW1bNapKEEvVsm2HBQCj7BKz3fWJuHimrMdWJvioRnzXtC5
4ubGfR90qChOUhv/dKfo1yx2FQukv5o1sjef6v329HZN6/NXMHFkRyFJe2ihjASr
AO2yC+ATF2YtcPRCXTefLEH7Gox5QHwXYEpTMaDretOdSmfKdbRd/X6QnE1wiJwW
74RFiy1kfFWvZHnpCQ4/9OQtiv7O0cnpWYP7mO2CJp3FnFM5efawiZP5JmxXtwr9
S1I0O1XosP1Dj23duR2Cjj3Y7PuofLu4E5NVQ9M1EBJExEBoogB3dyIN6hVKiB2z
nG8RvBbYYj9PgPw+wg2Q07tE6lm3krhFsoHGkjA+xukn//DnE/PuiP4ZhWn1xKhJ
37Gfrh6CsUeuNlJ3laKoUwuWpE2i5dr+etEoMn4nwA9zhiyAbl7Wn2doyGwitTd4
FOWmyNcLL/YBoNw4NXYKL2X2Kh9sHV9qECXsZZi07+ElyCDuIgr2fy8ID5rxBX84
6foh5GEB/gzvVo3fOllDbwzkq6SiZPFRxZI5IB/1ySi+vuwxEmL9Bd67BhzR0ofR
iy+DVscBQ38dPonju1JIAvaP4dhgibM6ZnvQ4De2DhoijV28/lna5dJRkHPWYj/a
8O6BKc2sGG30X43RpQRrVy48DZgEJ0pFG3umbtSFwNpnVF3s9r+bRmpufSc+YRSd
BXwk9LbmcDW6zOPT24UiITZJ6Y2aedTP2bOioRcpIBPM83XpsjRjaGSvQZ9mqokV
H71bCI/9bRfKCgsc8opbF+cu34b6h54nrg3685YMGJyjlCcjD3wGZ7ysO5fnu/Me
`protect END_PROTECTED
