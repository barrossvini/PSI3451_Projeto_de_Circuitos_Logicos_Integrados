`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fr89XIxup1+ySCDBbeo4I7QoiyqhKt6Ud3xMhKgH0HDcHfVp51bqd7m3pPQc31yk
BIFbTBeqs7E0zWEyGx3NJ7YzaOf1hioS70Y21YrTG2FioQfWm1bvOo5+4YLfal59
71ac5+msHksVrothPvK0PjMl9jK8VSeks3Je78UkFKWLBSUdz/FzhaHSmP05JR9C
4kdB+9DFsx7eSE0qpcMu+l7ag9g8PRjWZGApXe4Ow4lsCXDzkRqxdJnpcZpsGRKi
PmNJQ4845YHHeHndqnIt3DQpHTjdjF4N9YZ1Yxqd4aqgFNnH/i/4dIeIhh5qhbc1
oBKk7VqQvs3TEmLSIM4hKUMh26EDRX3L3jKQnSC6mRbfEO0Pxc2PjsLfCEwB3dkB
yrS3fSZh2qHlRoqbBynXmkdoW6HjuMzhx748wctmN0FrrsYVtGq1IYlFh3fH+dGD
CGL+/e+FqFs3fDQk5244ry38axIzIZIEzZLCND3lQhqlsWND3jTZbSsvlK9VuZ2v
CxeDbqrd7TSFkyWPmDu0hUoPDgaJPmvp37x+Es0oEho=
`protect END_PROTECTED
