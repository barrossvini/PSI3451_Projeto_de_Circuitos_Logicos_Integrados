`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KvUeDuaG69iQY81nulUFw0HlcquYRRd6k0iq9b0uY5C0j7X8HA7ugJYn38Dtu3SV
Iq9TovN/3q41z7rrUEh5tYKp4bj9TsHNgU/p1iRV5cG3IjtgUMTPwsQeWjcAFzsp
2o6BvxORCWe2Ic4JEtoMslftetbQVl/rd4Mu83bSDiJSUEaZdvVTp2iuM6eEuvEY
NSu+q/S9/Tz4frfmXYZRhcpirVH4gavNhCQRAckljpK8dJUCt2LwM6yw/DPHsxBU
CgdGQa4GjXPkuN18e5amI+pWu2BFFKAXsLVWDYBuLMeVxJoJ9MENT2ocNYmfTTRW
NR3ilBcq0H/OSSYKYwG+lQs91NAb/+gtbvcLq+PdWwpQ6S7Ek2cEXVRfvldLONXA
GIw0+O0SxiGk8ZA3zLHZFKH9njNCwePfkAsn2OBSfpl659WvTh9mZwOxihBIxelu
Wmyu31mwg/pBCqmXBPpck+o0BQ4+SWWaljg67teO6nPJMfzZKzEGVUXPz5zXz40L
t8iW/KL73+YUe3OiHwYmJsozqVBq2FnvxLxPn6F4MIw0RviHeQWmFytECGzVwfiM
hwHAii7Djsnl9uP+rW+8q48Qlg5xX0hFTRhHZxLEeJbTVegx5lbw5IEotvvFmWoY
Y9pXDpRpoZAGrC1cRjG6LT8bEMviRlWQ0mSOVZI/GxNhgV4I3tTrbqv0PfZSL6dM
HK9rLW6tSAQXcOt8ds2pKYvZoHtNdxJIZRPDVW5NY2kWPy3Q5pbJFHr+Onrgjg5E
MlNiJ6Y6DaFeSfH+VQDX2b94vMXMh2dhxrjMK+tFhee0/yOfNX7G5hOvLOTMYk/1
gmIQLjRSs+H5ATAw9MgdwimJEAyJ3WgyAlu3NkQfLmghFIjm1CQT9Md6/NkyJ/LE
qO+ThtoQBbLbvrsFZDEHHFsSU6EdLkZr7G1M0a1F0u9GcaAWjsw/A/FSLbPk80Hn
OfUmfej1+n9JhjIb+Z8Fd7yY6ycGbIrAcQcYmbnkNlBNL9ficPbW13xkqpyP8tsG
4hw7PCXstRWwtMUqcc3yeLw+p9/BN08c8VvT3+9hXJlo49qSZ1m4UI/uYZ7imJPX
MW1Dipo1f0RlxDP0f1rlKD/HEgwmQLOqyTJfYPvqzBCEyZlsREAFPfmgxtoVqLxw
XtPnsJcHfy37Fk2VQV1B0fXMmb84/0HaeBWsJjF58Fggw7BJaDfknHHbVe4GZE0k
x/AJDS7GmiReI3r1MyhsnLK61Ep/2vk0ba0H5gxeveXnmGFola0Da6MUnyC3ynop
We2IFTv/+/Ts+ISb3ORh9EXnksLxMerLkryrsxEZN2OSrzoVyR/9wlAjjscrkKgq
bfKvkkIHxdedDXkelF0vxFHmA4LZiixvxJOagUUEe4JhNFR4JBPCORlanSrXihBd
soXfYawF+EWzxX2AAV0Pn/1oSJy4ntD3CJl1zXE9HB8HN5NR4t25RYJ+AfmYAHRx
5WSPAek/RkggT73gkE+PY0HAO8GS7iOOXjGWL0YNDzEJTz+e3FdTZejWw/YziXNl
Cajwhz3myLLtE3a/tOM5J41lWkYoe4CORePi9E0P4pqUFHnADdC4BRjbOtkg2HKT
PhaWliYclUiuYoSwlX5EkABQllV9x9rAUjWCDfGLopnYmo43/uTY/sJ7oxhIFyYh
AqDf0yYuN1u9MqYDcVNyJbqiGcZBRmRHfYGNIdnFlYRAC033Q1E06ne1H9envbt4
fd3ngcZRnsjNL0StWsyrJG58Gc7IZmzWJNPEZJiqhX1/XwrHhxfzX3tnh1/VE5Y9
aLXjx4A9PWzm1QXk3DyAEaxA+wO73ieDLKEEtjt95051k6Fzw6LuFNTaCzEXRHWx
iXhB4o3aFz1AhYdGo7df6R6xoh6Ul2eX33HODyQRStoEPbUbNoggmRWddu8BPa0n
GCrqj1xtng7sv6KBi42LfzuM1OwJj8qdIDTk0EtZGjWzdOXBtCJ1iFI4O0LMXgTX
kPzIaeTRhERTwQ7COTxtudmzIQ+YYW3/ehmyKBqWWufZRw2/Jk+nTGvdClaNWHbc
MXZ3vmSMwgkAJDyqPbqY0QQw3gVU4OEqQ6akZTTBBtnF7WDTPJf7Qt2QgVFS3LGI
j/aHnsPAzij+VtBdSyRIz0PDQYkiVYXTPfHhCxfPxFBLg5j2rY8vcf+r9CZ5GHNx
1J3hZ1R/xYcmqwpXiGQHO1rtXVO3kbpHEOOGlMKUITzYfAhKL852ftrsJH6lw5NI
4WGx+8Wi6pkSBhCfBG4gDwLgUiGtdpoyFKFilAygdD7wo235dQHMyeq+SvaqPVWH
AMV1F6wcav5TcfQdQR453uZjG03WPrRMR2ulUjo13vmGHkNiqzulnMCdZr5M5Ger
BQ1J1my4HoEWzpO6801eeWvF+FN2xiv1x5/7/vMMTiyruzz4Qfp3VGXUgOzbgfYP
jwfDV6tacZr14GVkJ5RfeiVKdRrFgPv+TBMQt/Q/d+Hi5ARZLoFwHu41IcIit8Kp
Ka7gGCishgbFgIjOwW2h0/KLGEeqrwBksNqfCmVlBTvBv0lLqBx1m4JwBHa+Abk1
TBVj6955nP3ZDL0tYb7l9P5u2Cm1rIzlrh0ktq9wCrmZNNezstxgQffArWVxAua/
zEYHb4yua/2gKshUVORkaUO3sspcszDwfStnjpZQepv7IZ0jB9z55yTnREDC4w1K
k4kTxfCqi7KMdXSyPr/jGnwg9TTzKrxwakhDHXAX9+5qCXNPn9CHbq0P5exs8ekW
GowfBeFll8cSVLRnjpwBbE+UrU1bRS/9URu/j50LVU7JJNAbjfAtH4p/BGMMuwt+
CBs+UV6et9K4UNniotN17LM+5yc3jmnQaLwmjSR/+f4SdX1+669kMgRjmayQQgMY
JzqvNcBY9YssduncoQKXgBRyVh5FvPT6gv/pvyopIcH39dKnu7OR2/ajwP6EDOwJ
YWCQUSPw2AsYzIwns/kESvdOvRsZWizzSkUNr+HjLFtC1YPfW9V9DOhdJS0SjLuD
y6B4WTB4/3mXDKVupdgujMZcKzPgDYUzp5HyMP12cHLmL5T96fIJfn8P1EtlHja2
QtAcVhHQejpJIW3fYhXzvWTNU6Cv+amzD+X/wHKHXa5q5n1yK4GJjwmbrYAA3y/E
c/b3KNzlfHkGPoQNqaBdwAYtfxCnjycnDLkxUJQ0BX9uZ9z94XG67OArT5w0P7Ya
X06L4kNMFDoWZV+MQ2chAkELsg3vEkprqeH5I32cpCZg1oGUMyeB25f5FsA5WGel
Fv0QgCeU2KuzAj8N6L3DZd7phuGI+wbkRleIRuvkKqP7dq7siEZtn+Sx+NcNKLDC
bbbyFzOv53DCuz03ZCjj+9ZyH4facWiulDK8Be70+qiHeil7RvfxdyimDWPMqqix
qRjt/0lSL2hyi919MCNZqT7EgCIP8sNijGkXd55BAT8teJ46iEJYp0R0yUuGY235
0TAytlHtpY+1IVGRetTLhA==
`protect END_PROTECTED
