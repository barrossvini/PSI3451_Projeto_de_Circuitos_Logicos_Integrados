`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YaAXlt76+z6kCdnLR85w+QO9LctXc/Ty+t99H369vhYTVUXHnMM61B5uuRMSfvlS
jboghCFmnlRpdIcCcr3u/KNFXcubAcOaqgtvZ9wJOTJ4VUTzoSj0Ef1sCcS79S1x
J4gmA+YadxGKCIW/Ty9ck7KkWdYc0kSpwgSE8z4XGcJFMmI10TSu65xPIpCEjix0
8Vat/sSw+9eiHlDnwnLQfBzELw4AN+sVB1Db0yyyjPhjJZuhSboVZ/+vId3bg1hP
V9fEiTHB2vLhTJb3W/I+Hv8CAxWJYACvMpIQH0H3iw6G9xSwAo9Dup+7hy5iN++S
SxOVVyP9RwSWJ2jMt04vIiyrEnatzRIFdpyZ6VFKJ3NnevDUXiZGlyYpH/JLESTA
IvtNBB3ejMfs7TIoV+SM37idWgEOvgf0THNLB+gXP4O8UeaztZeXTF0J0l6R6iKg
Sw5ex75EyLIS8OjRLaIBDSQ8MRXUPh1kBFFLb+dqapB4sqD4irqbMT8P+9mdu7Hn
OTM3ZlBCG6lt0GGybBjtdD8+sMmElYLfFBebJtiXLNGvkSb9/7xe2ej0PVYHQQHw
B9myEX/DtuSGtJ2Aleeo4bAE2+FNs3RyyXSmO7J0OeieNCa3ubfFE1glnKCDf/Ry
SxIPek/29S+/PM0udS9QM4SakqPUVhWQjDuiKIwkn1UBTkiWPY9M+FBg/oNIjDCW
oEgzyzHGuMVlOqoob2SU6E9NBmkkLjriKhnEldhx1yzjjiwTjEGVsTukcTHfNsf1
C17Y3YUHMscssMmyRK8rIasU+gm7k+cHTODfnglzp5NeAQogui3/VWZwgeh3jYDA
IfovQA5c4gNcwckQyDrvrFlfl0x8FbOu0vdEgKlRCE0pJ/zbNK/I7YaWvmPKubcu
xbj29i6US9alutdcZZIBW4KtklxlTebhlhFGnkeJ7UvFdFP/vry1WVj4YiT/tZ1l
gs/V/qkk06UzXYEACyjv17skJE26gRNJPfowP+HY0ZG4veM6azQqJPDpuWb2MhQl
5S2zUipZbdpbmahIIp9P8xw16So27Si2FsuuS0QLmdSYTkcAW2w/CeQMDgMydHQC
mSNT6roMQloaIgrEE781PF2vvZw0QYknPjUJ76D4lzV2sNh5oYjmiM8pfa7znotQ
29JVaVm7tP6+9kySNnzuBOrrgEmfS5R++Z5yHrYvrfIYFVMqvlkK9f9IeRQWJsID
4scnyCxkchLNcPN8R4Fjg5B27ePstJjuBIYsfFnSGG2uSNAxJt7Hy9ej3Qjbfw6c
Igxalqe/ojLJ6H1HN8CC1CM+AD3hotUZRuCoGwnczRi6MtUnUIizPxeRE+/gx3P4
iQ62Lq4KPluMnf9E9CiqKqPQvuoUUUvpNiBfL5f9upLGeCvMAXNOvdb5W6Z/Mm2t
5AmpcVEjJXISNlG4Yyw0NL/D8KVJsmzWylc6h7B8jl/UNuk1/swLm1nrTGBLkGEW
4BJK0MUuH/K8JgqARXb//flsgnKMwnuzZAyDU7dwlP5PFkx5yv5SC6QEORzPExTD
izYbiUpTyZIrjcDOtiUepColLwNO47Scx2YtNtsPaF46Tahd71QrokS+XqW1xkDG
mGrhjeD9aNxcKuPhfp8h2f8Tl0e2IyPjta6qUOPFuVlaeCjLIqK/5dYl4SbzHh7d
kNxbhwxSOrZf4T6HyBR9MK9OCD3t95DUsvrS0NqDxtm3aIaJnAc8Wh/SguITWdZp
vQPXZjZDigIq9sKoP9DRgroXy+xoG7Uj707eSy1po2NEAQ5OZt+YiTehm6AMNOtH
6JoJfjhGz1Pzsspgmx/GVuxulVt+xsZyCDGvc88AXh7TVk/IBi5IuSFdUIcqW9gb
b3gU8KRNLI5ypDZR7glxbg==
`protect END_PROTECTED
