`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Hxzf10yMHgsmgr+tS+joXN1JiZZQz+LoMo1p1c5X4+HewXwpIECcb3H3JtLFvEI
advIWDmREGHY4AzaoUORiTxrym8lqPDTXs7aYGidx7HmAki8OzfHzDzPRXLO1mBG
4/APPcdRxI7W0lC5A0GlImNJ/pdblnY1eSHm/g3R7f+GYIFqn75WkO/+v1mwytEv
LfSyZw/76a25tEcRBgRMGln8DTioMi/gsNR/woIU6tItsq0wRGzOT7CxVE1WghBl
4SC47AKxw/cw4P5XlaLbzgKfbU/i4dwrYHji0D7BqDlYPUg7wLhcYJr8X4QBUvxM
S/HxeNZyvvA9ckTztZOxk5+fyLRf2O7jpTqXKQNp0CEBbM+QkwG+gAt4JIx1mxe3
phSxg8xt7hfTn6XsBR8M1d8wsdKsZickko0OxXxMfPnlUNOb9Llkz8PTUaowmIg9
uxJTOKMZ5X5ivWnCTtyr5M4Sn5FnQ3wEKsOeKbqMPViqK8HEfkjfAavm+/e7KzAL
iAE2x7LnldUZcN0V2rFfM44YYEeC0Ca5APtbe5+HnpuKMCLRZXw48Rzj7HmJHuXS
mzhY6i9Ipttdou/ca4UhTH0HRsQNNhKEXhgDVT2y6p4qwAwvlLucpmsyknxZYI4t
KFk4qY18eF0zPrbAFpPusEecoGxX0nPjA/ewPFc2O7Y7aZPSxGgHG1BEwJCrJ4dK
KhyNjRK8P3jclz9SdkZeGyqqj1d3VAouOWgKkzouof6zAXwFhOTcFc+WXppbGi8F
2PCZWO3nKIDFfWD7WEGVpCVREVlo5Wq1LmX9eOkRWirvT62QaeYC/eNYA/q+MFwJ
ikp+Not49PU0QaFnfPzDsvrU8Ki0LGfDYN6nMRTT1Cg=
`protect END_PROTECTED
