`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y0MnFuqR6VDAWR+YZ3aBKFQ4+A5u9QCn5KMCYNvxQpIdPt7JF2VVPSPAzPmFCDj8
mgifIBnGqTIBFdQf1I27rkS/oWH0x/F1Qi1nm+uu1CJkMJmbwf12zhRkp6YclDRb
fA3ercYvpyLvH9lWFVpwG1g2rkGFuyml/3+gGQriO59aC1HavqSYkYSvUJUy6qbY
Hw0tMqSCwpnWc2xF7TQ/wc1oAtWDEjjTaOWVdlxZJsycy6nJEw3MUKdluuv5+m2K
WR9WZv1/W72TfvOeotrCRNWBp9E8BsnNne1XwJC5sndrkM9xXsnnY17mTymaEhGW
nxMIAeqRG1M/twPpYyUvYrBcpWgErLE9MbZH9Obxj31nz6oqhVKJjnIftvtNJqFC
2DxtV3/BFAax0KbqY2npAOWKBBM0UPBdZBzbKEgW0AKCTfCFxZqWC3I6z0cBEzqT
cVfe/iaYlgnpX4utiAOOMulnOIWRkHFtRsvbre3EAt1d8zr9CnOjAcSJ4aAcQeGr
SyzSf7OI2O1sihXNNTPSsB578YwzMMhrRVUhDt8K4ZgON58ezDa0wWDuWWupVZ47
vLEbL7ikH01FY79fTbKUJcDs+BqyrTnO3lzMFJDeDvpjQjXJ7PasRHENNgv6T1UN
KFtFK2RzFJiSAXf8QqQNWPBYVDFvS9Bz1RtoQrFc3w1c5dFGFJMfhYLGypWSV3ht
KHW8UVHWjB6evPjrysYh5X42GnYtjCBL7jyFu5espDNGfMg8Yo6x5GmZJWrz8oLx
OqfS7RNW6tabGaTiNMTBugChuV7Pwpq3n/+wb00gZreA7fKHCJ2gtIjzNVcHKbeb
nhPDKhdE/z2aB+OLjYL+AWSimEv0evwKY8UcX+zWNyAY8ybeGdEUkXyn4D6eE+cQ
h/BzV8AR7NiKac6TLMs9y65iN+b/pUCuwlMktJLb/8W2EpTAXBOwJqEoFJegdnM8
bYtszTZmX85dAUMcrkiBefUvTYS6FmpAxmnd8/bUxDoxBixx81XkpTeSRfUh63HL
sRy6Nl7Cjj07IARsqw7PHR5DhMlDYVbPG/FuC6waBoxn39GT39h8zk53Dp9UwT1l
mZeWqtOdCbTh7mdCL4bcDTk0sb6chJzeU5Pjtcd+j+M/XPkXOaSM11GjPPQi27el
3o4JaVMfT8tNPInUFRo3o6fpFZliUix6dWP/+kdZVZ0lanqqJAg59vJbSd4jU7TD
xtSyMUmI40AM03vZXhK6Yw==
`protect END_PROTECTED
