`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FAhfuXOMU004e+x6vOncHhR+oWc5Hggn2PRZlD6wYyabvBE+CJxz8lPpXWytpvn/
yAixpkWzjYlPtIgJmBSMbh2m9Trg2Qr3XbFIA31w0+8dYKzBqhbrH5toeSqC7sS7
ONvCCNegjzmGS1EmcukFoMzpIStJQKkdtRh4Abw7Cup2U4B3hg8h6vpRNXVWGgRJ
5MwVrCmOYsKxbv3WxaCOHqUep1Zm+H5jI52vtzruXE+LKL/KXRO+Z7XRYYq+rp9V
CLHd7cQlkTwDtlkk+bFJccSrT+oIU0wa3N5ewdUGcz9Go/QY3O/aUeWAqLpjEHl3
bg0qGEAMx9ppoHj1+cQ4/P4OdG9Zm0utxXIqjjYtjR6YX2zW75UD8o+AAoTlMKxj
g9d/TwkP9ac6IjK8pSDc7edoqi+eZYglZsDnatdw8NqIsHcD5lDEhuqyokDzepXY
dZJBttCfonrts083fAgkRv859YCwEpE/a5NO01BKeivSozI99XAXGjzQaDtU+rtA
qgWgcqEn/BInyFn5UuU4I3QHHJbk7oQYIJ2lslR1ZeMVU2Fgph8EbQA1WDLA89Xy
U/T8yUxADa9EBWpnyI+hOUs/u5QXtcWixEbM0jGQLFtam5RskvJjn13fSYeJh+Xs
mifif6k5JSvic85i/lIavE1gylnb3oHwV4SN1v4584xgEHqDyLeUwRUX4KrKWfqu
B9MmobzQeU+Wm7GNOPHdOSp77u1GcDl74uBuqJ9RmVaLExVdT5HpDj2lkY3DMnQl
Ng3poi0CzA/1QmlOtECo72CCCuLvHic2TtvA3CZku9ZUKqQypQUXX6LRhJULl/Y2
5OOxmk5Zq6o0hEJuHEoTTx67lIm6lTwlnzQ+s7RYIUdj/yNVLnLT3Y1VBc1yOI1s
wmD1B8MgP1amPoH1yej2oZgoduD3PQDkRYe9PMyeWQhf8Z6nWBcoqe2X9Vy0nbfB
9LLjdvmnsICDnI59Cs9qwkuft+LN5q3O7KA/kMCNPkBhrUDXVNbYTUjZJBKDtc4+
kwkO/jO/fp0T/MsU7zRInizlSNG/gDXC7S07wxesBKqSht35UdoRtFap6p8LNoDr
s9kwOMH2ioUT9zzZZDqfLBTK9FDzYX/Jm+hzmCLj2H9upsrx5mNfAep4ZkkWvJu7
vNiw2IgrzIyLg9yZhRUebWxX+kbfcbRqMV47D5/iD6jOsHFrlSlbJDcpS0ES0DMJ
kQg6MOhMvFJPGhs1937YLy+zNiGYh+8u0DEkjcIKJBS/FIw/fYFIzJaOKTBGr8il
jEi1ns4FFqAz0+NmT7GT4sSJgPp59c5NCsMq4Kd0fJ+IgCCJJoBfaeKb75PWvQ3C
rOX8kLekStOKrUqrl1MOsn9sOOtKWmfcYz9f+3d3ixVdUbjC/NSdLNHZRIt8BXSb
h5op19SL53aiXWAneSJwy1FDR8CMRpyT+sAx5GEIVP7pMPupNcPnyJEKqFhfgzdg
G9ZY7wPwDTdLQjIclDSIM7B3zH6sysFKOR6yxw0sLDPTTT2Z3HeLcDztRhlxf9SZ
uG4iEyZY+i6+fnPrGgpcMm7w3TPhz+rPFnfgdgsg0hMk3s5wRcRkTCOOcIkNCkmT
0dTXJ+CtayhqGptU8O7ieYE7tl1VudtVcX69laVAyS3tAcfcWsvFxSpiPYB9S5A8
H3YokhLLR/2CfayI2h9OOv/jC66U+kkCYFpU7wkS5M3sjPhzbP44dFqgdr+HdJFh
KIA++CrllvLjFnpLd9b2XHsB6FDMa7OeT2gFyVEhxdUqRTY3uuV39je8aegf/1lh
3jl3zrcb+kd9OljZ439939x+jZH+zFo4cQeX5vy68bQew5rjGaYvAdcezr5N2TeY
HY8mBgF7u4SBD2brNsWGp55hapC07Z+Buv1aE3ywoFkj5r0egDUT6Wa/iI4O3Xln
2Q+br8gaREC6JwJTamfY5jlNZeWJ0ATZ4Qu7QYWW9tkqocnEFTnu0XwczlblRF0s
UrwclKzmaMiwWA8PH+pmtajHm8O8P7jzemIvQnSaZXPjhcG8u/+5XM9fH0iMJSAc
NojDdsqFSX3R/aTVYa+y8XVuEkG0whSP4i4Ssvqqx/hAvmlDLRR+SLkrkpoMJq2i
QKoWxoFbxIAxK4j9bZZdHl1lweOJjgpkmCGifjqOTwSzFLeq5X15/WJjmu6Brmbb
yOMf5dkYNyZctai+67QjNElhW5z0uo2wW3woNUZ/CoHVeZbyO9ThrMQxI5bH0YeW
9wvKP1ufcIIQGDbzGgqR6D+Uc0adyQRmwL7FW8iOYBfWqdS9QL+j10bK8tBwwWLP
nKYwaoiIG5EkpuiVquTmdUFrb6ZFwn944l37kV2QxwcXLdE+RfzcjGP176ggS4Hy
o/DcYHBPTKe79UwvN5FQ77F7eW6qhM8Ya66kWO3N1lmiAbtR8BE0TDdGEYihpEDM
`protect END_PROTECTED
