`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkhq/4DbhtJ11Kx6P6+1arDv5ZWCGvMRQx7pDPXsbhpU373tyG+R8CnnpOdDC7A/
elLAFWOAYF9O0bvLrfvJbZngiVTYKnd33RLoyfcR5RYPgyL+/vOt2f7gYCogQjKU
1oMCGvlpf/T5giF+xXXOoj7uVt+eHeUsxqmXmLcmONpy3RVUZrTjZZD5W6qv5BMG
Gb1zdz839TqsLWOvAKk6BH1btme78zmSBeo3fDbl06xfKM2uyy02zl1Rqqm/Hs5m
6DfFtFwQqY0ZIhOfIRfesXRTkjqAEG09UmA9AVvpxvIl+jXZEJwA9l/XsYoR8e06
scZPxKqPNXZCbxoTiUCWu9shPIeagrFzcA9H68mUGzec0eS80zEqp1+jFw3hFfsj
2tTRWYgoKR0eY7d91KpvPLC2e5zwE3k9s7K7VEwp5FM3vXDIbszYXQjg+LabimkX
vT4mRZYuTNN7KTrP3snbNSevkFSTAOaQLjfDDIFoPx1ldlAYNqQ3mnqNo9H2uLoD
eSKAnaug7NHgrxTyxbMKcbFVfXOuYGcz552S9cJHff9uI0v2k71Z5IFPvmb+9HnG
TwxOISr9PRU8q3qgxWICDvzxtxSLmgzTofLJ0KfUSHg/WNgrgRauSKIh3jZXvj+N
CA1FGGgxHjB2LmgyJHjcvT5HZ3XRtpXevWVeu2ItvN0kREKpDPOFgo9ehUyu/N/w
kpOYTLA5GuGg75GF8pF0WFJMHacyC/jc0JIE6eE5BZLAg0kn4uabiTn5MoXWv0cf
2j72F0xYsU5lAdwzsayUmY1ZmM3v455uPZpQdSIFBgYWjjT8jCBE7AbNgODeo4ig
ySwefdfO5uIuaViXXwZoOQMAzLN1yZaY8XFA+1fMtRc=
`protect END_PROTECTED
