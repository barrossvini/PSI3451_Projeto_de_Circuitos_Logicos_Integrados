`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KytyF9dQpkuT9jejWHYbL99cPw4iKuprZ40zetpA5/Lmd3ryDEMHtPTEjkIDQO8h
R46RKwVTCGXt/B+gD3hOXvcUFGgD9jxmtyEhUgwO70j0bvjtbU4dnfP7DwNsJ0BO
vCuX1J7KYnhXQ+vUE+HeUc/VpE6WYLZnNUCZud1FjS9PTDDc0snnWBv4kJYiuFJ8
xBAOLHzCV20C1hbUW3Li+elrACKDiF48PUiG+QUDQW/Gt6IIhVxOHRBqdc3mRw8N
KEvQu8fZLXd+KXYiczHDbVkooAQgdrxh8NbhwLTr27j6127Aa9mpPmnkvbZrbm23
Edu19s/CV0s6uWmy7zBPRUJyOearCbBCfi9l7Cu+bDq+arfJqdpvxVYREfiJqPyc
zbnFOgKRcfdkfns9Y6BR03/9mmtWqpPuV5/ck8dq18kWVs8hl7+ouUp6wJ90+rju
C4lB/FScCa8pJT0PPc9Ro/3YmCOvYi2ZRhBAnw5ber2SMRzf2UqhTtuPXpf4HwYy
X4jFOKQjsgeFS+kypIWWtyXCb3nsadvjzoWe7MQpHCl/ud/3blR8Vx0DIz6gUdqA
6U0/+Q0wyVGcUjwqg4p1s51Z/p+TLQe5GbNGxW6whcwW2pKF8/RR3ZK+M4QBSwtk
wRgYrPN7xhSh4lJKcwLxXhE1+4Qoqhp7o4sWuhPD+phjZBmJ6b72pmTqzbKoFPtU
2i0jsl5U1MGD8ZcIBj8yvN2i8JBPcINlj/7a56k3uMqTJs8pBUQHYgrNiZGs/hPW
NUZk4n9KZ1ZxcLArDx+WFwLE627JRwsu/fEvbF4OR8hrpOFmx0wQx+6dUMk/Axxs
LSOuKGY6BdL4fM7UU8IAWw==
`protect END_PROTECTED
