`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tzcEkW10UtRtB7dAs+kPs5N+ZT53mGdPPLTJfZit4dh7VNZE9Ers7n2OicScbnJJ
bogOfs0lqRkRsRh1I2cytc8xuJJes/4UDacQgBryBNq4bR1ZO/Z+eGezO3rji2SX
nF73jF31tJsPJmlQnrRusIC9pfFvJrhE3QDaRfinnseZYelTpwRDt8uwNyWbttVN
gcpi0zXx3/ETPQ8D0G38wUu+0LfPX/41O8sW4ieqxVd8kPRYE42LMpUTEUq1bsNX
vaZWylVnBRnm+jyFfPROUvxC7nqOATtOBUMChlqnKODTQF6c5vdFo/uQlXnf6hda
OJzymEZOQ0m32CrrgkRV6EAvkMDq0H7DptAeE9SM2Cbd/R0dn8BjCLdVCUif8CWy
fs+sEOEVwjazPASqqqUN9TtzcdY9PqmhmNhMjJikJmq2V2oryBwTx/E6hfr5hbIs
9UOZqGOJL/3Nhk+oUAr3GGel6BbWNwyN+WvuslJ5anm4MT3oELZLS1Vj4b04TBdS
6x7hAwEh4jOKkDnFGgdiB1dYPH+sCKimXzAhti6zALLiQdRL988gel/BngBgcLG6
Tep+5SVlL+DUrp2Xcyc2NLJG6IC88mj7Ktg5ok4xytHh7RUwnT3WQNYO3CiHMGVi
U2Bx6MIDH+3uoL2ZfVMrjj2nGIkG3MRogi9qQDupvD23LNSx7ydMJVuY5vKsFAj9
90kJCqFC/JG1UcfVjIOdWH7ogPkwmf6nAs1JGwUFEwLdnELoJre/bj2L1aWcr8pj
B/xUQD8vqSaHgjyz9GqFGixJW7jINFjmXEmCEPuQv/7ApvbV3KLjmYIDHjoflvEQ
WroP18ufFSN7Njj8pMrqXYI9/8wV9K49ZqaMVEUxGMdHkExUPQ9Bv4cfX/ags8Zp
7KW+qEXTPZCdJ+RY/IUl6+R888J9ci12bLxk4jhZhiC6MtuE4RoagbCZDovYcXLP
0cwKIlOOxH7yPGVoTpNfYqTUCoaYaFCKucrqXukAlNSsQ033mPDyAurjgk3t18fN
C6e1zqdml2zMXIkqsfCDwcSBhdJtpRPBj9Ks1004lZlGkEyZasn0Bn+H5XUtNEZV
EdtRK1wB+orqD1rrZ10+9GlLRuQFKr9KE/CGJkOSXMoxmlwxqMa+eMK+tdiCtVhY
d71uRJWtrsRrmyA++Lie5v/Rzjq81aSKd+pTp29QKFHR3tN/Gb35w0Ex2VYYzdE8
VoSE+ZGd7wPQtfLj8Vr2W4vjo7gaXAfQlmTOee8N2dO5JU1j3+tljS0YPeRBhmCI
rBUxr7F6nfIb5J+g6/c7/cirWNU5rDrSzfmmdZa9Erx0rOkOpkKxyGo6xEcgcglM
rwpIdtcLxTVS+CPzIC+ku5TVpGiNPdjbi0CtRBLsX109Aa6TJ1TOaxDSDSrROcRs
/8+dw2IjEznZDfcpJE9c4vmCL43r24udI3FMDcB3YzbhlLhvSRABruaZicqc0bwJ
UGkimPFA4BXwjbbblalkqieWuG+8H1cH0vqaeO1MNA0SWSu8pgeFAAPk4CU685K5
DpSiC3Rnxbn78lBhqIKK9HqDOm/5ZKJJsygfnAz8yUOmscqmi0qlW7P5y6/Pz2Ph
HWw3Zqf2wMBiVxqG+2OWUDGA5Xt+uao8D3R9t2KWFqisdPXA6iU8Cir8ezw/vqDl
SJQxRMO2uKLPxv1oTGeOUBlmqYDZe1tb7seg7qUPIxACdeJM1hL6gGA5xgQdhPWd
GgQeFvIauMjhea6q4qhFE2X9Qs55EEd9NBTtwROZmnHRPcMCrG1zQhMlM1t7tjex
MZ8M2vVQyVE2MZRu0WFXusrD60nz1gO7DgybpsUF/3mK++LXwXCtyjC1gXgQh52T
VtVamOZmHRpbexaXNhTfyA7xMrmbInDH18fII9VAc3JX/nI+A/TonFfYvt/c9l1l
v976Xv/pVlVC255E97uCy8GR/7b7Xy2IgLzIM+HyFuFRmDdPiURgTq+8+ojBE3OI
yBtFAo2rlBQPCujNZuaKBcbclVZ4ZZvukAwkSziy21nRa0i83Jr3IARz50JbijNT
U6nMqDUz/KRGCoHXOJwedstSehDprY0+ljgXpSCe/QGcr6pAn2b/MhtQI57uadUs
HNQvWclZ6iR26D6N6+I4qqcsS7ft6CF2BJ9GDduTGJB4fgnj4jKxZ2etJokDI/fh
PR3It7aoZHOwiyhmkncDINtcy3VU7jy28wITCI5zOAaLmmYvxa9nfuTqBWuhztqG
BoTK9ADRr7fLy0WgwfzlETVLsEi7Euy7/tyQQ95aDTmSL1BD4nV1qp2z3lgiHywR
8BvQv65wK6F36o32wZgEPfEKiut+KGCoJcORjTSIWRuQ147TjJ+ey9WQz0oKJ6Pg
j93/g77h6MaQez8BiOLzecvSKeSRY+kv0NeabTbkkoiIzswRvMN8CXHqCs9Q/OsI
+8XjlvOodLtMrUsmekDyhBWRNQlnJaXQIEKCUiIZs4mx+14bnohocZX0G7ZTCUWB
G/0UX/+5c073hclaq6IVaEpARVcO01QcC5HLjtPvD30xaZ/CZ8RJCFTje1yB2rSz
v1Oi7S9RkIlX3tEZYuQx9nxfRdCAPxjEXL/woK802z6nNj236s6bQOERJHHVT39L
nZEtYdGLx/dsFLn5EusGs96O1fPq5qDMVyDKGpwkGV9qMeBHiKXbh8IU7om/mIUY
FNv+rtnB/43QfkFoG/I2ifH18SxzKHPT/JyFEh0IoJI80Pviw13Q8+gG16cak2l+
PamAgctgp7jKhJD17ooADgDPfOsWPiWPWAJLoBFUqKTPehG9pTKPPWTxlZtNPOts
43BzbJk71JQbrCU4KbFp/uGhCykHY/IMfKHXDExDX05rbH1CfFioeijY/4R0oUjM
+UbeWSgOcbR3SV7grrSHXD8TrAafFYt/Wj55CqnNCRC8nutw/5OeNIYRsMp6DxD+
4VfqPcKMdNvWciKTO7yZsIdyLppZA8+uJwcfL/XNK0ctgai3dX02kUiL/ZpP1gQJ
0uVxtNkPugZGIhNa9URE/sG59sXhkr5zjzDWQQOsU+YiYwsfR+NfQXZ5Uk6PdUfF
DyIaLhFeyjfIP873rWGXT9tMea+b/i+/TqlBp3nNAs2QKPSJ7rjQ4KavkT2X4ROX
OdhUr2LsjuN2w7MhXdkcuBs9EzycbzkIk2es6RIQ3S4zHz0x98OrdN1+mypQvw5u
SYgdnCEIyWmpxjFfCoRsYCGisOy3xUO4T+YhxVgP0YxbGwIFT4MiVJRoVyK6GqMb
dh0jA8zzoAH/oaoBT9+tFRA7r3VhfKJZBdhg90rlW6wCO4DL9xqLeYaE74x2/WRY
R1LSGTN/bdht4zQmZr7zNXHO4UaC6fQ2eoabrISRcsvWB3iQNWhZvrex8ooZUgiK
M5pZPc1TojEpzAvRk+zrWyPfYJtjPqVzsxIwBIP2sLpGiqAngcfnnzWHbim/xTzR
6faAbH3ffzxAov9+OnagUwSSw0TYNEGAVk587uZiyCpnz6iizDeA5fpomPQk7Vk9
pUjZFTHSYTMSFnxUT3rUaWHijiwqrCywtiCh7KqW5bx2qwkSFpAAnc5IVDgkaowF
kKKl+Glljd6Xqh0MVTVTLqctAvQlQLGS1RcRR6NkQNHu7nSFfDxodpbR+7faWhT+
jwiKU88KGDqVHPqEu8ysieKfzltMhUAJLaJ153qsi3/Qf5CHa8EhtYIP3GAT4tEa
bqhhwamVxFN9YB30gT7GdTRK9gIIH36sSLjmh5GLKDVQdMdFmlIPfVUqxZWUQRa2
qTUInQpdd5S9djBdCtVQW+9dhBVGGMUdllG40Am6tTsQMQrisRgeTctEiyKDb8x7
wnuR2lylAYHEVtlZKSPoj80qUNt74DWFDiEM1ZVbNAbW/7tT6kXSnj8xHCHgxsiz
yT2QVVlNUyPAlZMt+Ng3HpxfIKDLp8gDfqmlSPB4nfF62kzEXJ1X5vgU8Txx3dFG
KlDcclxGiY7wNZFWaUsV0fRN0cqhaeKpjRtAr2DV1F1yQoGzcz4oIM2wgVdKIf6w
rpAz7On34wT7Od03blVTV/5yajRwAZ6HL+cdEriPpj8r5ozY6/mh1rceMye6ZQNP
OfB2KZZDSFyf7Pa8PsCa21fF9iBdHMF5j8XKRqv3co9j4lOfUJ3EeZbe6e2KYV78
Qlep8pGzFRlp9ax7rNxvgnXMi3qZZd7IFjFBYpiWz49Z23xZWmiMFtGybUstZpcB
cV8XECNCyh48FfwqAaTqOddx7O1L92SgZLzcGagSL7KjCISDUUUMblADtKBZB5aY
5k8tYmnsl+x2XdjRhVifrALeWrirtlnJcMsZho+Tc/1dIpCekqmpCEL2717T1PzE
zbU6mKENb8H1yjZcQO4LQ9YlX69Phboh4cjnsDFrI2abs7nfaxbJAr2VbmCI7d0L
XUuUkEFRV13Lndi5zI3FUttPhbAyAxD55KEGQ8Um5v/duZ5zRKQaEznF8wvpZwAL
WLcoR2dpQ4ckBtOLFiARVfSJAorMBK1k2CzkYqXq9VcoLXTNQo7QJ36EsyMXHvV5
bQOWvKDy4Z8xBsZuQ8SmA8KkjLOGiswqHCIqoEIexCZqidBtVy0UclcUfG7Tfb2t
nrgGz4dtz1OtfyyvDGbtH42+BNtxs7702UvAuLMxgri16nCX9kCD7N0ektXYXdo+
U5jHuMmq2H/sz2t/qfsrFSpGab+jP/9Jl3QrvyjXwmoi3Kh1sRnnZ8hAraTgnyX3
X+07yI/IXqdH4jg4CbmlnfZYhaqQRVAzkTdghyJK9HK+gBtYTbxysZVNnqZWkFqU
eempSrSpkJjgdJuqbQNc9QFjP/Hf7+4eG6hoG2EgHwOxo8y92QcGutFjc25Jtbef
IPorkkFvPNPYmvWrlnNvy3yDFMhgcNEX9SK5lOb7zm0XBk3kxkCdZAuJANWqYJ7P
Eie8j5/sGbrgpd73xnooP1qOCudMWJHZkSsitVbToLC2+PNM8gzdBVvpMp5v3pQ3
rpkXdhvN0jQw3Rq2EkNOayT1ZdsfSyHrbBbO4bN5uRL615lqZP51N9D0boacNDTQ
nMvJGCIf53OqR1cj5mhAW0W5JjwF75uYTSE33SWyzs5whRt6lnC+6mdIVSLViFjV
s+W/SO6xVwDGewDneLATbfyrP3Ysqo86s6pIwzFcwuaOwdjZ9T4Cdb15m/8eUFdD
kelF5HsMAcg3KYl06+42JZvqPgBPjv7AhRZM8z2lPB0fY8Hjcp8YG656HlluHqUW
Hgym2fbBq//gKiN97nUuyXKCJD+wYj9zoUvmbmcFBNXvZOmBkSh0YM/NYG/E2Gzg
PWttKgo+s9LdnaAtgUr2o0TArquCvx+ifNDQTRnbOEWPVgVu0C4OCbAFHZeQMdbn
qRR5ex4DvVa4/P68SecphqLGq0LqANfQfT5ly5Csy1YW9EggU0OuVHQ44YMCNJij
ZssVTPVnUY1CTqWkJpZCS378CyzgrR6MlPq/Q8Jn/YBGBbqVfT+Udk2F0ehzQJDk
H0W7TE6+D9KOYzZ6O4nIsXJP9P2DoeVGaOpBUY/pd2/rUI+QjrkyDhulqO+Eenio
ePPCd/t4rBywlX6suSSkmX2TQVUfEsaBjJsFLOU62N1lXrnuqse6pP0tkLU5QZ5r
18iBjuhw76YAPVgijVMdwpFTxWT+GS2iKRCxGx/3zf9aBNntdlbJI4R42DvNuO1A
w2cGJivc52TRvnTaxtHyIfYcT/euYi6+RyLnYdy+RK1LHcypiPs8tebu95cKCX2L
UtQsbpqfbAFd78NZ282vsdQUh157c4Oo0OZ8FgZL2UP5oV4qpJRCJK5nltKd98CZ
e4z+4gFK8EXXEcXL4eULRYTuUFLluyqf1Fjs8HWxvWz3cae2NZnTbh5JCgRBetOc
RwM4gMkXgQQ4oP7Ajz1/cEeO15nizPL2P1rDjgj33fUgo8ZcdRpmQhY/fW7CkYGC
+ecV+Q0zGuQ+sYQ32kfuTyQksxq1YcPTLY+vt3PX1Dc=
`protect END_PROTECTED
