`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ekk45gs18dTW5g2NanMOE2DQSgOs7u3xgmJeDka/rijX+rNhR/zwwJqFHA/GP+of
k13T/FprUXcJsupbY4uHq9gxFBKSz5kwCsIrMgn/mN4Aa38nIfGh1eEWT5B20sCP
1YVfGrY1tsyC40tPe31sgQaZEDnRdXK2yXGf95lhNizjh0VgZM/gOPCiNVaHu+gI
ehZ1y5IL4+24nEAcfyOAFOkgWpjNIEOGzqvVStmKZQEhc/Zi1ojIH7hDL06ykC7P
KKnNvnn5ktvQeuasfwMUApvDOD4EJ6FGE7vJx3dS81sC/a+225vftF/j7/cUnDYY
GEjSBlh2+oUslR2zicRJXM4HPbyywStwwgtCIr7SCXR30CiYuNNgpdlWp0CuQN3X
+yIGj0KDaDjxvhdnzidsnwuY0XfO/aMCzn2YSsGp0oYzCH4B++yoIjC4/DkUukau
ITbwgLnDw/LerRpANLWHe8SqrjnSl2m8YzR/UlRTTt/nKkoTemdYeDpvGslGfpPg
a94l1+nxEU4xgPIeJFYTZTz0r707UaNiUn3YhTcsVp/KBXjsSnVRgiBXvEJHkH4t
JghjF0ThSBfEjoDfEiBS/yWujjPd2Uuq1nU1VrVMTG5NbG+RmS6YA/0knCkt1kGA
kuTMy6bH20XD7oGieSmIVwkLdmI3Tn6hTTXa6JW71xt12BclZL+MaqgfExIiOsCg
6nzyBHaOneWvfVhufnGmJdTltG1bnBe1c1V53fny6QDIcb5qvXEsfzJU9nJmNcvx
vw3FXti7aewgENtfzoFCbJCo4ZYvNSuagIUZQcmAFA1HFnDv2lcBt1+ySm7W/Psk
ho+yBISlb03MHJlekZB2zZzyCMqtuABoQmoGbl9FDZHrhpwgyWejohfPx/Jn2/tW
uwv41Uyh+wxgHJsrfxZOO2h2S4kd3J4VlDIlnxwxGC+7GT5zGuTiT6EtmyaVCuxU
MzQA08GZhiW5hy8MIl8uU/YRbSj3WN1ChwgrsbSifGb5Gr+Psp9LthaOzJJUUrkp
utGt8k4ARxk3DKQt1Xrjk7NVcDND94TZkeo+yEg8i9oarWt4Pty6YbGtTrMR+smA
ifAYU7QOOxaKaDs8Z+aoiE2HdAr/dvuhghCr7tSsZoKhiN72hHpLVYQcvrtwVOKT
IQYG5ibgoAS+n4piLqWkAPW+75389hnQMdWObrlI3zPtZEWE6fZf8u4mgdJ4e90O
jHh1OQUxOcd4Rkw1dtsAtyYMbFol2GRH/68wB1tqFAh+dwn5SOYsUIjwEMpvKlt3
8bOAFG+jbpW+ZOI9rUzVa7x085DJ8askRc3Vk1zGGhdNAZ8B/LE5t0UR7LmSOEhE
7LFlnXETLQdGPGgSWapRwPTrZj828WYpfcXADwBmsLdvRTkgIC4eSSJwsjh0y+PL
jPpNMcuIJLLxaSlpUMT6qkTRXeUMnagGL4uASL4gx2m6AoijKkaYV5UuqF9nJsHF
fFUBHC6hC3xvnQJ+ROyFHlBVCv8KLsdrXcic+uk5mkdRoy1ThsWo+TsAzTmJptTi
3PtOWFXkU/P7h7aJFH/ioVTV5ZZlF/RebEbDMDuRx1E+VD8gdc5O3HOIhMcspvgN
R4oZtWimp7h0pe//vLJijoPNR5AvuROwFXylQkz9MOOQjp01UjBPWoyX/FuZICnp
7zBU3rlsNZ23/4SehvCYmAINmjo/86yanY12cxvNd/Bsx2vTywY5RiOzrNUSX50v
`protect END_PROTECTED
