`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GE/wJPEKxcTgTGdPbW/cvqDGiefLuGyW/oxG4MvY1we35f0WLl7gLBUkrQV+3FeC
jQJu6PVztRfS4e51H7neFZGknppa8Td36aFpxu5ns+zZzMbgKks+s+RnIoHMzVjC
aZvOAmVLkbFZJGwCt0MulucnijGVJu1VahDuW18yZFPmxVGOWpHTaPuUdH8u1ZK7
/3rNtGbUOn9zQoGMQEwT7Elg0KAx/dBSgVqG/on0Mnu68Xn/Mkg9EAbzmluM4DkJ
j1RsAPOUeKwTdoSdY5sBRDoRCGN9LzyalmTuKscVoOMuPkkZcLKUfD86TgIIgV+P
FIUNanlOFza5bUnNK2LB7KhZBEYPuVpI//CXP8iHCL4OdfcKbZFjpvywXTi3o1Al
JMjGEQflncQsZ0CRonc1fqXmoVOGLpCAXVT1fg9CDcd7bTCpNxHiuWYu+VD7GBwI
E+5bkC/ALoTk9MYnDOcs1T7+j2bhRIf4GVsKh6VY0v3IFpYWAZUlpu1EIU7Hi4oI
14qLQ3Hwed/3ml/omCa2/dvRC7OAgkHeUxPMLagEqnhrGbMwXLCLhf5w+zAvLOHT
qdq1IY/Q6L+/DWrLeMuzhgpOatLNDbhr/iFDdF5/g/J66CkJsclMnKlRj6tU7lOK
tEynR1HTVS9pNPu9onl/m4AsZ1f0pHvWigR4uLdFDiWR8PG8cdPRlySd3Iu3lsa7
PruIVl6LBy9nRYcuInheRyggsnRFux4tIV2xRebZNOx9q78TuaF3Tg5MDT59IwDT
jR0hiPZZMoO+rN1RnnZHKHME5RD64CRSP4A2amtHQ3GqVE/A3GHP/au7JAvLk0ro
bxyhO6V9l4EyuCqwTU7oS5iAJL61AcD+1AcCjoJw+/7P8zSxonymOhZNX018dMxc
MMwUU/o8FI9jH/gcJdUctIf0P+Wnq6vAOSjbvuNQytKmlbIJfaYzEleBTCWYdkn/
0HJxycpqGv7/n3UVkdfC83w8FwrcLOSKtrkfmC89cyzEqFQTSIjqDPU9CVNzIMHY
DHrnZtKSq77FcuKcjkPZx0GOo5t4d3EoHkXx0h0HPMe/Xf/ZJMIXBlj7wQzT8S2z
5RoF/YaecTgMCTTlTaDCXG3PFRIQ0p/C7rL7fjPfhOd2U59nwYi7ozyL0p/hDigY
8N4pSQd16tDRjTv5fuf1K/ljBhuKA1HoKtHdjho3ebrkxQxncYfuHLBL9XNqZRGo
JGdR1HvW5oyCi5RaXcR3s+OtAiptE7Z7i+IFaDiV7C8nhZTjanNjDvQPkh+5vtLR
2xuROWtKbKkchKbcyovQb+IGxQel6B4ZUnuLnZCcxmYcsrhACuu+XXUATnz5c8I+
gEvZBWf0UfdYnPnc2EFa4uJbhLv0szb58dgIOL2BFwhxhKCYgMlKvnhgFEdzmiBZ
gr/u+D5TkjE5IaBzVIS0UwxwIe8mgQyNpP9u94K5G4tNbN3JoHRG3PyB1wnk2fDG
QLoXNaOALQ6UdIZ0zK7Wql4yzsLFTI+Uw2eB7jJEe7tDo6J55sduH1MBxaRZQT+q
6YPTXdxKfpe7vTBLjKEgLeDoJ51IV4UWi3jRCu19RWILpa6iil8oRO0qfuwxrrOR
XPUcu0FHwA1swEx8JIUEohhLAh8w3/NRynTwxyMYa5uyqJ59k/boAr8fpIpasAJ3
SDOW4vw3TQLd+8EvDJ/RDEeiqAg9xgB7CMnRX1cYUFp6txfFZib4iizwAXA8oaKU
JfsS66DP1ow/2YO1S6pJ1jWnQNcoaj+4z0RsrQRt1LPYUOOz/Ql92R7s2ydsqoDb
JXLOzZ9OSTlfHHLp4qv9Er8+EtfxgWBaD5j4Yh3lxoEPe4c+5C0zIF+a1Nbttd8I
tPgofB6WpzFhoU27+8y1UcvVBpmIvIYmYPrwZf1JJlS4dHv687OL6vgVWxtDSf2R
Y74bw8SDnF4CXXqmqrsC6VdBYKDH2ZVotQUnLN0Owniv2Wi2eQk9EZgklsDD7Fk3
YbOnQIK/n0lHkoW3jgiBNFIKM8UBcOPmORDFYb1aZ1T7W1J0wN2IxZ8P6HtOnWBK
hqzTo/iSGXEKUBSp00AbA1RijofSb24EDZ97gkzAg6KpGqUt7JW5WGwKhRwoubq8
th2laFJMA9NMyzqK1VghRgt3+vF6OXi9WHlgZbONZmH3W+NQQpM6KcRjT6E85W+8
gom/i0DHUL5y8TfcXp5+DswRhhj21s4OkepFhTMQ3EGJ2BiJMd0OL4UIJwEluuzV
OVu1IbmyV0BjaPrv6LHVXfhiP6Uq1kXEr2fmNQ4R1Ognrm5vY3JDwtCaA72aS/c8
v1AL1Ot0HDNGA/LwOsfRow==
`protect END_PROTECTED
