`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KUIoFXLBTlYfWtruhJqv+nY6OoYtO4VZTKS1nsAIH4vZSslujz7Q2hCOJ6zHEvp8
FsiHsnZTbfF+MAvItcyp3GBTStHNIZ+nPFd1fB2TkvM8d0WE8mD+AF5nY8hyXXcM
tACyIF6LziXprHE0PWAozPkZmH9Nk8Qjk5vHJx3TJ2qGxXunflCNBh7uzj3WSbNm
PAkS/wWGpN6ldrojpb1wgc7Ldkpli8jwPtxYBWqHx96LBic4NsWrzMIzWJgwQQdm
QL8DR2dLRUqveZC3k/Dta/oRZRAJCqrilTQzhN/nuNSTeoYueECmLqY71If9FErS
29BaGNhhlyPhVgByZADi6j6nroyNE3+UaMRkhhUftYfswXCX1AvaW4zLyYFQkvqo
Rs9jG3zX7q3mZq4xaQ1sesbIVLeu7O9XmqAQDC1YkmzFOeFJZyONF6Kia+eKcmYu
weliB2ODErgurXDUHdR5r/SOWhpW5inxrhTdwSGJV5M+BSHcWgrRcD3Omi7VpS3+
BrLpWSuI0BGff/WG30eZ8Qdtp18U/1ZfwSM9lMGqMyAqGCwAvlFnxX6S84wD2CWh
BL1x9pxdg0Ck0VhuFXj4iz4GBUHZ4QjLIQAiRpph5M8V/Zrk55HAGsXTK9VdzI9S
0brKD7olYDzF4dAlz3ZGPcgX5X2ly+7pBmes9PWO+wHYoUOfk/cB6WzQ9kj+YECs
8z4XJrHoFyyivIYViSPu4qXG7xKYbYrp2NfF/9BWtepKNoD4RN7PcMINHd85tEb2
K9dgVC0QbQ+u61WpIsaChydlmvjdDUg4aFgmpH3ROfBZG+KrMlkY5x+dYZhxYxSq
`protect END_PROTECTED
