`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K6HP/1KuHRYIGb0Hxcxckrw7WJrCtDfY5tEyHrUn4BRijNPMGqjiiYF+ZI0nXO5c
HAD/H0WGotzvRg+oz0sEaV1JitJGfYykPs+MhOQl7HFTZQrg5kAM5U509seI5Z2t
7ISu6JNFbK6CjBr8lrX3BDCVERERa1WsmFOx/1sak0FlmRfS+HCo8w1BokqGUvxS
T8TLUB48Kdhghiqi21vhgKz6baQYAkCb55Zno44/yzkwljFHoYp+611Xtb4mg3K1
vesEkCnwN+s4k075k5UFlTOzweITRxisdh2h9AVgAy324bfRVKSOgt7p23vPA92F
CPSuWCk0SpNB+Id18fAbt7jfHY0OVTlOpiPcR16dtoPk28/yrqorFqay9qt1wEWT
8GbsO2nKWlooATzhOubCCA5iprB/xDafhEgBXVKIa2eAszwzJxF/foRVNMj4UaBb
VzdNiObhe2e6dfETbl11nKRII4RPMtXDfIra9HtSM/bJ7ZqbSh7Av9twlLD5Sdap
heWhfwSmj+3ERLTRIrFxJG4aF+8xFNsz9AhFMv/a8xrpvD7EOqKbIAyqkCYLrTmW
sKGbjT0uJbNzXi0neo1ZumtJAZHbZb+G6yR4WHiyTBXKaNEl9QJ7ijZ5JthCaAE3
JtEn5LIFfxIVGjiH8P542onZA3Xg6/NJQbtwr22wYv1iMj5Om0DnHe0MEJWL+DbC
m0e6dMPne6ov3M307Tq+nXJpNbBvdajvDYMoOW6JzI9XcvBPuo6gDV5G/HWPh5Jd
ZYsNsAwNt+gPH4Nx2Evh83SGL8gfbQVd2YffTouBnTJMaVne1pmZR/9dUj6RlYl5
vQlcya7rS6pWT3UoEtnSTojqeMDCBe5BLShe6Um1oMxMQY2lU0xI6+y80wkdcVWI
IEmz1Bc4FBeHCCHsZrZfa/e18g6ybpLEks+8GeDi5y0XAMuuFqkS8fJALuv2KYr/
IGXK9THgXSfvvrIxLFz4bjemB0dhPNhgdKBJOSeir3mp1W7yJeqFpAB0IT4YJsIt
7JyfVqAQRTEnM2hAC/6dleNYNByjMrlEY1KZ6io8ktTn9Upd2vwr4Mic8Zs2lWlS
nHB1ZbhjBBQctba55g7Ma9aD4lHCzamyo1Zx6cG0GQHaSdIgYK2m2nqLdPTJ+qsM
hTvsEran9eB0k6Y26XVOATLW5xpCNfmgv4oWLxayYbq5dUbVCpLoOKj6wSClBuWg
RXVsBVa9H4XmOLJ6IzCPfpuv1lHS103b4quxjU0OSQfleeHBT/EgQByFh7VsIyVo
isg/i220xnXO4ooJyDghy9TThX16/aCE2k37bJSwN1TDb+HEUb5654gIruTZyqwf
mKnf2xgvajS4RHpIhdR0sO5cAPTZ6Xa/bU/sJKVMihGyU+f3y5c/s+Yk6/F4qGVB
S0/fNcVaSuKwU/dV6tz5x7Y56DTJy6VuSHW7yEOmej9n6tJnosK/FlqnYXwGRaOZ
Pa6KVsVgFqgtHvVM2wcrKesTl7xn3anpxz6rFtjL41hW4Ukb0zVOV168fcSsEwjh
bzxM9yDBjxPYz8dnnYOI5Q==
`protect END_PROTECTED
