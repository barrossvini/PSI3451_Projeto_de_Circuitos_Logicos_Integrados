`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QbQ+dGfQiRJkrakHoZA5UA5YZdpnwzz9i/sbUruBo4PIKRXXjU8D5TwZRqeS8S4B
vzApK8FcuDrzotOAjZlQ4auCvqPvLNNJ6oYf5eC4Dvd5HniWGLHa3fFzeoMzB2pw
QRxQdxrQSXVsxmdeA4DfGdOxLYgTyj6wL5GAAV4iGkFVQWKC+uzMLv7FiEbnTc50
Dj/sI6j3vS/taauKngwHW5t0NBeckK0Dv2cBp8zNSTzf3RVOTOLPg6R4oxx5tElE
T9Pq4zWPb1qFXULhsQ9e72mzlSnRkIMAyeBniqwzY8403+pPboCHJEuL97uv0neP
hCrhgfwOIvcYPG5yFMagl085m3Fcr3mEcjhWYUAbUw7xXQz79WdKyiAr9EHdtS46
7sp3eCpVGVPcbmgm24VWHYg6SxaZGHSAII7DyGdi9xmwe2Wxxx9hOLjC0IA6k8lT
YvgE7JKTs5FNVFyvM8TFBtXzCmM2jJSK+064iz1txOFVu3/WQcc6F3wNz/varngD
8cQWxk+hrQcFVzLbyl0tMDeYGC3oYA5E7upf2SP57yGMNGdvWB8ZeF/cNiDbzSxQ
43nYEKS+tBr/Ga/JryxGJGXZ88F6RoCbaSKLQZdPBy7aQT8y/lP4oEuc8EXQ08+u
69hzSbV1ve6CLY/Mk4T998vEI5LSM3ihwKw0qIVDi0uDSr6ngW+L8QHV7xj6Qx3d
EZfwzVnOEpIthns9IGWbGMWuk9NY3pqe6nZ1Q7PZpMajYRfCaDCYT5jUcMm1awnx
LtLB/OOd7VcmZM7/AHmTVyDD+JhkFHBGeskQBOFdWXkJMYL3zkHPaYPZ9YdU0o0g
Nez61ayMj95EFIwo9w/SCkTAACnQgrcnmbgletlKjjFxlA9PceMd+3VvUKrxJ5xh
yCBh8ustBipJtMhmIEzzmhRXrpGYSy+Mjw0l4Z9PjNsdFpoHmoR2hMh18pkT89lv
c6F9cKUVmFWf8z4Z7xodwOQ1U8ECw2DxZ+Hd6YqYSOMZeEGesXUUhpnVYshZrgYp
aanCUDxHUbLdUBJr3nAHbvowdQlDhiHg614oNvkaaJ6Ls4N/SgRI5+wfSO97Gssh
nNEOjflMi5UYElvUNd5M7vLMICqeSwfBIn+5VrFZMAIa6bnKvHgAegD8c00Wjj8v
w7MbPAyTfwlLzshRgBYVcNtwiqRyFYk4PUIFyLke67lvI0oUjaSvAgOQruW0Do22
QHO2YxZIbWtS8uwlgfFf9Qwk5CIj0mH4C542Jr1dp/8VPBkpOhlnJ8X8FhPRcOoE
2HXj45JuUe8TZpq1INBI4lhpMujUsWk6uGTyxHbRNAyP810Jf7cb5vm15o5/98zc
Uy91mrMprclxOTbkKximKSoa6BjiBcY/QhFgvLeWi3JO3WKNFEiLIyRhCNGeZCap
3dKVhnSmaktF9p4RlMDirw9kSv0+YvZsTtV5ujphk1eke6748JpgXLREpox3XPsz
Tq4UmYvkHyBnu+Ng2PPGGHnGKEwjRe/6MJCGmnOBa2Sr4Su8TAJX9CV3TcW6su9/
mKDbMB0ASdKMLoHIyLbtDFn4O70JTigNqOqVFpO/JDRjMnEhUAp90rCe/9B0npvC
FnBQWe340XY5hmmXK+F3jOm1U0ZlNq/FWWMkfZqFGFC4PDPQ2oz5ezaM8C5aZwWM
LnMARxXzgDE/l8+oYrN4Uo9/f1GSXz+sucyE9hQ030SUBb9GCPBFh0ZpDtv7LoIb
R0sPNA/1H27bh7D3RyrB+A185x9oj7Hyrm67tRM4K4gEpCE36pdioMufAoF4dtgd
zUr29nhASptuZZiTuF0AhrEJgga5N17rFMvXWHYSN411wXfrVlJz4mOr1JpqFG2Y
mNGYTzXlJsRS8DqRsCY2EPHuLbs2JSXoVtt3eNd3zVLG4A1ZpigSKwAuQd0oQm6A
Qfp0HrSru16W4A/5YeYi4SkPsmrGl9RPjT1pvDEUfgCKh7/cLaAIbhWkJoB7F/jq
on9UYqWSaOJyyaCJKSsH80EM+U0YeRSA9wkViQIjaMMvk7I84UAyYNkn8xtJW8k8
UUGhLkcMffhRHe8rURJoB6a0uOmqCg684myVAIXeodfwJUTHiLqUU4qI+iSUJM0v
pDm05Z1OFxS8qHQUTsrEwO6lJjCOLJKRLIwx8p0u/9AgNvYDEybEaPi5mOyCqI4s
r69AFZ5TY/L7gNVskcG8iRp2gQ4e/8HEPHSXQOOY0m22QleG/J4/Ij/uQeDYJOj1
672qKs70uE7eaLUSnBhtHHLCSJ3wcbONwigZjG4dwbcDEFNfLZh0ncYE15Qs5bGZ
9e7E2ZtLEqLR9b8NAXHGAL7wmkLPLRr9TcnKLwMK8rzUFHWwaIOJoU/0dEw5BUgz
f90ai40Ci6lFijzPXNdEg0+NyTLT08VEQBzzUy4KvZ/JQZ/nIn0WM4cvuLVzjiQJ
sdtYsyYUh7YWKCNUel3oDQwKJ2rj5y4gtTyGiFFX4S5n3Ta/0xHQAiugv/wuSXu1
W1F0KPBqTnCKUqCf5LfdP0aun928tQZppE7OLdVBkvDN0RwQnqAurL3meGUBFQcZ
8UyuJX4VjGt8WnkL7lbJNalm8HVoBGefmR9tDOU9nLbQRX1142RYF8UWD/WSYrQB
+8rxuUv36RtKtqhk+SLXTvWzxCkfSa99sGIz0Z9XVCuHsmE3s0dO5vbHI/NgLDr4
k3WrQzJLTcM1TlrwJLW7D/P9EkqTSyJcXrXb3uTAShiGIkHvcw18SE0GpywP3HBN
SYj0o7NuTcwUqD7bQruqSzlAU7WE/DsXKFMxO4GV31+MbBXu94HLhB331pYf1Slh
YN1fOZLBYcB0xCPzkdkQJRMoKD4PK5w+Qm00Kb0DbApZ9k4dgDXGL2/neLULiQ6c
hIneP8nOJz4wwgJ9cSvpb8A9swm7973X3CLjY/zfe+M=
`protect END_PROTECTED
