`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ltS0ZXW1M9Ok/Mcui5/9wIRmpEmeYcxfAaxvCgA0PtnjzWYpUGKgYgjwtmPRhh+I
6ZnMVqVhyMgZlmdYnXbIWUHZgykvyxV9hO8QGO6S3est1tsm5cXartVM+TGNMWiI
BSRGJkRjVVq34hDDnk+TsM6ygZ/GEJ2n6kIG/ksqcL2rymVMiVg5D0TDloQ09tvS
32iYWZ0EnoLr9LN0MDzedBsFTEMoRewdfdA7IoVlA1c0A8ckfTTApvfvP3u2eyKC
D2+s/icMdjSIZiGqSALcFZvVgeeEXTpny1T9OEhnAumH7xTTJsyiVq8Rh/4OOn/t
7a3zsV5IMmqdoVTS3vjgjBCxFmDHnPY4MrlH6IVvVO3l8wAxaHsLJP92wxuKXrMW
nQ/sh8L8+2BNb8GvFlN+2EN/q5qV1YIC/IHWaI1TS2kZgYrf4G8Yv+ZNHQ6vmxDO
9qs/9CR/1qadn6x8do5G6rXX/3kiAYjwYJuv8LleBKDNFBZ0tNACKl6eEz+O17m8
bi1IIJ1Ev4hqIoPW6YYybT28IHoVuP/14D+c6XJkYPJP5ohmStUw4v4ELMEF0wdt
tc0evBKsoO5z/FfGYTD12FVIDEPLTow5ndw/3ODSbNWnGVzxLOK/I+TB9YZr4bPz
FjQbXoQJkPbwd4QFKQLRTM/PrKtEK4aotnjdFcvuo7gKUjtruaXf4L0VOP/H8lYb
1rv6TaWybVUmxsPtCaRkj/IjhuhQMh2JuWMivf30a1REpsiWqwE51NLi9Y+c/Wr2
JuTBtwzl7O4VXDv8j7JgTQQMFK9iv0p4fWF6nHHQmjVKkKTibyIEA9uJFoiYOi77
47Usk5/4N/sCNcmwYDoBzkj8X0LmdMSVze7KOTrQSSy/hzUi0edl10FWSU9Gbr/H
j4gnlcjoWVm2wLaPMf2IrI4mVPdh33LBoZqHyBgZ/6+pWU63Pkh2MXUXVtdvj8BE
tL7JbFCvkIY3wAfIESvlVHH+3eYROBKEztrRCmWpqh1+7goaHGqT+vksFVylkTXa
J6Ob9EvuwQWYpPe29+JKltUsgYKLX4WKw5HBkUZKp1OhjzjRxw3R+eGX3/Qho4Aq
ROHBsU0ozaCWHwFpxDJHdPY9CXa3zVlwjzvwWF7kPjaDcaqxKdUW+2FCJV6AnjiO
dp1hdrtkwRdvypsoUMcgAd5Xq4tIzxH7e+jkWHTAwNz6xbSRSzaauRN/gFsNP+jl
rWxHI5h/vxjEi5OhNRr9/kJeaaodCAtB6Zquq06WeUXATNJ1CVAmgr6dODkub4l0
uFBRwxagjoTP8C6AwibMQ0PQk5h9eIARKn3pxyaJ4LbsGApF9V6QTPhB1ubK0bgz
ElwvE995lCROcVSnKU1kYFXRQsgqNN+MjLeZxpiToXaelbXlpXv+x84j+GZZUA7m
wKyDbjjjsdWo49GOL5LhQMCzojze6EgbggcQsXJNnla7ls0Y4dgqeoZX7+zUTKrb
RaHx9BQOUN86CFl0llyLKNy1FdyDXQWOamij7ey7raCANweJFFHu0HANZ4+rT9Ay
YCr/yKCzpq/maZ7hb0lA+eRTGZaTWR0RRLGcJxOi1An7TDkTqYQQaX34VbzQi/6k
ZveV+tfP7PUpG2t6lnY1m0eJU24D6QUXDwX/Gn402mxY1bjOT4TqHJimKM/iUxtU
s05MkPnxKhNqc8hvVvLO9jPjAFi8sO9Cmr3gpOiUEI8=
`protect END_PROTECTED
