`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
olU0Q9QJllYJT2zma3yVMneWGC7Hy7Jgpwp3bRbbeCKnuz3ZnwajmBfvYRBcXGjv
v8l8myjMNNMytoFfWU+Jy29B6+jSLEmG2wrbTAd0bFuyV3Z8CRgAkFbgfDIpx2V9
c1xHhzeY3ZDjTVLRVgmNRXVyDZtO2Xtpb5BcZKY+pDqo3o2xR2Yu9l+khc6hDBsy
HSN2BN9WI5ZtfD8aoadjVyhzA9zOlIIEQsh9HEiUSBTAPAV91F6Z43Y7xiiVySQe
m0xJY8NNrQGpHFEp/D5yBWXCCM0eYMDL4YN2kCOOmKrTe8CbOOsubDw92h2kthMI
Me5LQ0IQ1mpuyOwgusTRow44RQUqCV6DtFym/2Jx4v3EKeJNB6a/1G6GCz2eNWwX
rHdA26zOwoKESow1Z/O535DnY01Fp+BX4zKp1x85ww3REHy0BafnJGIO4CUDntJg
hqoV48ugiruwUbxrarQJ+1xt17MPeuc6lBOTx6JPSCe2elbOYVm+JI6jwMikisJ1
HqaUjj/rBdzolPTJKF4Pf+rNch8DYn6JqOltHMG7ejszrVCqFOekDu6+/ZahMl5i
I29tNcfdvW0bJnQH4Hl0OnUVy08SaY4gVl6kX2vYqC884mjpc5Fg791IEJqpqGGa
o5k+OvAj3xq7mS2JjPNNnx6mV49Mt5kSufzeUUEw8dplUHBnkIn1wV871vvxew/A
jAgCc3Tauu99qm9ok2qcx7CDdLtPFalfCkIjhcP1Og5MQoUxVotJKR/8qxUdhDhF
PhdicEQeetOwxXqqNz9FTE0sCvkdkElnt9/PjbloaYazWfkraGWlecvC9anPTWd/
URRhihthKrnMC0ZWnm+oQUC4wA0wT+AX47Mt/YTZLpk=
`protect END_PROTECTED
