`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Arlex9UiAMNkOfriAdMEQ5+JGpSwdbLG5hATCuXkU+15UQkrRPKiobHUKmZXqrZ
0For+i0c43OSzyUe8/homSlYuHR4uwe71hEO+AHrmbPeZxw7iEK6VrqWa4tFUN5Z
xc/B0UQpD+YRFZBif6Wu2J47GjiDZMmRuY4/LWS9cTP+8nNYkgSoyuWpJ/GfF21S
E/4iiTNtfVJxeV3DLoOzTimFbtNdJy1Oq0ju7pNmn9YiNwOh43/fAOivVndDRgKm
+NcrO3ZhnqNkxEN41ZcVTUnsWeAAoXlYyDJhxvB38mrL6aTiZmC0ybKgb7yYQecN
XeP9Z7RuOKuOYtpg0pKc1m62e7VdPQ2UkbowBWuxnZ4zJ6LXozy+9S97iHvE8HBC
b6dciNBPiz7LnZTvzKxBhTV9vsz2b8eGpeS2UWPRFMthdUIdTqqWHRgu2jemkmW7
6W7ys0zqhq4iO51Ug075PArkjeMnIvuo4tIZpVbBeAGNF47+QrBP3NTHsrcmDpih
BHnAI3kH1WFzcgjWCD9dRmUKDO+rTdJ+sTT/IcOXtOhSrXy47FhX+BpHeubEAWTE
cm+okw3UnIU38Wpeu1oqSwmGdBY3HWqfiS3WyjpMZOdrVYOg+rs6eiy8ahk2WlNF
LpkEFanLcsdiSbG/9r0Z6w+zaHYL/dSkHadxLsFPpphsbgZZvENS2SGiSjS4pLjd
GH20lGyzZg18bNDGN0Cg5DPSKooT4X+m/r3vbTIVMlmxHbqLnYfcYk+m+dNC/XPA
TjALHzjho/4tjWZtEJp2s9t1jao7hGzv6AYIPRW0SBtWysrOjHfHdKMGJyevKyd6
KnoBneQUbpq1CHDEXvA5iQ==
`protect END_PROTECTED
