`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TBmXzr+zWm9LLZwSxD+VrYSOzWVtGbWSEhOuEUi0mFS/+1EVoMBLaGnqTebenYFa
CgwcEMX+R7MvZx0dBzNw0NZNmtDP4XnE1vWeXcGRVZ18GDBLzNF91KtLKcrjiZNu
OhWhZlLO+lto+7OB/cuAmCTkNzMQikFrLWXhNPyjfU5dBWaLUdhUlkzGgCxiHVEH
7cI2xgzX+bNjEGp1+ERrexv5Kh2tNs3lhPkCEPRWltnlsg5QVW0GVhXKKEWr8o8N
7F+Xep7hVuSINMp2l0M5qFg9tn3OtPq0Sy4XXHXjXKksJxfdQpxJSKBAd6+GLRkY
HmfEWAIuLw8I2VVyLaVobW9SiDUkFpS6oRkI3MVkLUaSf8zASEb0/sBNB5WYIcia
fUaSjwvDepZzBVVl4tNvgNuhK3i29NxvMGppKb6W4pHu7rwezUOhoSyL12hVK0Oz
4DJ2MhcOpKQolQT1WqlT8JwO94QGYg73/Zk9UQhrqvq1X36MXSMufN29xTOFsFUy
F1KnCHhTsmluk8lJIcJ7ez0aFWgmOPhh5H+nPOzNHYkiuBu4ibgVOyhdYBSPk2+L
MstaSxuOWBSsAlRrKcDc8gD6F9EX3AN0c0hsxiENdjes5UA/6kkiiqZEzxlpRagH
vQHo17HreQCyeLck232Ai9JCYBoJaRrLZGKBr3PQwFT1T0eHHMB913KGLDpIdJ5I
EVxUjbzFVPsV3WkUTCipdZDaeI7/WgqGKsVI50vmcIAkC1YPgcIkXSe+YtcxGxV+
aypkXorSHYkPKyqcSPVslN3t5ySEjtsFH2Do/VYxfrkZSZGV8FPHXKlPpHqFQQIj
mlpflNaoV2Z4MXnZ+a4H/oBnV9vHn2D0h/AbPmpioTl+niHr4TQBdt8ncFPVC3/R
c62Nfw7+taJnlKO4aLe4Iupf/9hAfJgrBXQnlSxYbFvXLUDcARpwPjgBUGm1R6e9
5u7PzHnRkBJf2eqImFFvPtA/2HB22fOYC78Jk+L571bTNyCOWmfGYfm8zPBX5gmw
bTZo2XwXwJfeO+ELqPTZULq3E6in+CJ9Olpulf9Phr7ofj3K2tcZLQ5cvsLCkEtS
lQtcPLIDqx/oIVRA3JsHvT0OgakOj+IEwh3AXBFgudYMwA5NTs9Sl/fcmu/Oaw4K
nq2D6E1ubx60a5gwl63OnfMUlAouay7UIF3vjCk7V1Mi4FwpNXcfM21xvFZpFuTp
bX+EzjUHvrpEUqg4pzSh0FeBr6I0CuRBQwbtDIA54pH/StZNcGLZeaPwnqWn/3rm
mGnWKDOZtu1LENs5Hn/U7yiMKq1Yhy6YcdQo6NhU7z0aI38SDdblZPbB8UFjYAoe
Xn6Amsv/n+3vlcDTPH9MgaonP7gzOSUrXEdvJLbWOb6jaE9SYri8lLrQOPBq5vMS
AuahAn69Oppzh4wF+JtcPXQaS5NCuUETUvQ8ZbhPpqF/8uMMnj9ZyQjeArMT8FwN
VJXHnVRnRIMxz4u0ImrJyeGrqpSV+qGMTpWy+baimYQjM/upf1OWKSlAJ0wEIXjn
uJgLQ1iggErs+xprxH5WZMpea/h0wT6kxtit6Tq0+H5Zo7Ruc+AWNbqwRy23GJtO
rOxrZxPTTaNrPug5yV/lDHenoLJFaCFYGmfe3afd35hZumETs2wB76OJdCRXyfoN
yLItDaWe/WzymHyoHdGHh+goZrJfe4Xp3kw/mXIElPJ/p6TJ7xaMYRjeSMQtTtAZ
H1EfV9PxIkfL8kdL5ZOl/JS/TXmyjNk1nas2wCF7WyHVHzUxsJMGqGwIB+nRgoBW
kRcDdDolcI6GL9p70MGT/saQBL2aIR3fkyz++3ouvGYOwGV7//uVJG0y6gufd2br
dytEhREw3aT2uzCGaIri7WphP62fmLF71OndFfoJR0uR/IipwQMWpCiqlQCGuPqX
TqcWaPOKV71pCwg7cmc1hm73+1gTTn+qutFNAz+3ey1LKMjvE5iP6nMNJ/39j+xL
Oigl66mkyESH3l02huBRzD6aIQ4MamXa7Lhm6zkM1eq0JrCVEiUXhgOojc187qBs
b8eKi7dKrYQTO3znTSUSV/BSmhzkbvBk13/tTn17Ms/u5RAsOr+Ak+SDJMNZw0Mi
/UIRvU/lxFUhRvNU5IfTxbxdDN/yEfAv1RbKc64WRQCqUUyoYjrMbyQXEf7YdGbd
Ppu3aztFVZXHqyWgJsljj3Xf3HRr3I5MlR7xNRkDL2imtYzwbFyAi/o3JbAYM3fX
j4Zi9j+kP6ZOagtyz0Yx4EPdVZYKn4Qy2jV0SwUbaLWdtxwKroylCUjXdi7Z6/IG
WIrnF5AiTIbm97siBjEAbk1DHg/aTq7ng5E8rDSR6sBj/x+dk/Mo/utshQ1qJzjZ
7RGS4NCtr7kAsLZEyWGv9LRsF+UVO+um2Pswz7LwzThRQ2yE1imQdnL8cO+jip8m
nK+O6uKHs9jp7UM36DHdTCz3XC1WKAXqtLr7LSyPv94FdZAE5qvNmtDP1+eKlti4
w82haqYYVp/9CgRpx09hvNdRwzCPYcJIgCcTa7XubaHhrp5yq2j5oAhn1Sq3jzZm
E5QrxtVdm4yG8Guk9c8NcZZgrtmY72Hm/DPrhiHfOdDoMjh3cpCu90FD6DH3YzJW
mLRlV4crB9FrvIm2TOBYYhxEwGWvoODpz2zwF3i8rfiNDjzQR8jB3rqwauZhY9Hd
iYs4siWVvhro1RPJ4x/D3cwrGi/Vy6gdhzyfnh6CXAzwNANtFuxlazZEhdnevC40
3HWQuYWAEAnUAu8620dSqX7bZ2uvZfaYFerMKwK+0iEDcpX3traglIX0vkUKthD1
2JhGoUIJd7EhvtpFooTsqIsuwoM7zq/4O0EXdbswp5N1fxp2pP0QWT0MBD3rWtTi
9vP2nyO4FAOX/jgtd/jhjBhMqcgaibBzwCwuXl1A2pdyKt28QK5XusZz0tvXg2/5
S1HD2FAq2YqLwVTpMeVSnPcIbPRaspY9hOxP0NaAV1FdlZ74d2IVY5JvkglqfxNs
UOZkfng1XJNdKfo8RMRL+KDsHirF1d7UlhNdaeeYBeiX4P2v+0R5zq4iwU4ylI/o
JFP2vog8tVsz1+9KwfCXjwOjAZl/+zc+iZlkUZXk+Ol/dd1Ex6qU8QdlDo62Rx1x
PTeQReoUSDN62oVDN8VwB9ajS4Kr/GiOi8HELxsx9rmiUcoFnS8+aD8IMWnWhG2u
uYF8/ffqpI1LWaD+31w+avhiEvPv74mxW6MNMjy4KWN6L+FzyhVqqNH/V5zCeqNa
mQrzApNXNIpaRGqRmJZVO+WPFe6IDFMOsB/nsrb6SgrODQpz2pe6dmRZEZgFuHId
tdNtbFnVQhzYwxQ91h3aK7SoG62txaa+tMlEbhYbseqqkircRh/9BajUSBSAesXt
AdMHx3v2HB0P74VGewzbQAhN7uaQPv1z/ZZhSc3OiDy/4M+Heg1wySXOXcUm8yg9
1SPdERQiiUqLXt54sGbBKSFuzhQcurv/KqN67KOKry8N6JqnOYGG6TXnVdq9r9cT
SBNoV2/hbxSIviNJmxbTfFzW2ULom1EIgXquxTQ82u/eKGiRdHNBptNDaHGyTqBB
tEcxJyjARsuf6JTDXGHot0e3oyVxKZ4YKs4RyEpGZ8pjF+gPGwaE+r9QYxm2qQGx
AhtZj8TWm9Dg8vCeZhoLuEpgwEa7gkZ2xQm+5CkXPytokF/T2qUCYivcB66wcHvO
KTaf3/tB/tdjdn2ceNgb2moRRTqG1hkA8buQaXMLPk5LTeIM7VTv7aMOOZZcv4N9
ibS3fmkBX3pTpGa/pfbOsQiUfvFEfbPiaW2SflOvwcpYtFkEuXgx4WCTZYxi8n/e
PlVpR8352SJYIV6HU/ghyFEsic3MLvakIElusIAzGwdVrYceez3O7d9ZMHkJngVQ
YF50SmEllWQkjQLQMIthbLnhqZO2asbalCPxbcCcm4WMWz/RPbdnxDypjL5YIi7v
7UPIfhBoAvmnH/UUKoZL5q4Mm4lcb6jlkYCtuaf5xr8eHgWVKGtsMxswonMFO+2J
wWAqWBG0RP7NWGb9m26yjV6V+9rBzs8GfmrQZ9zMZaV4oDoufNzxJFkHmKNRXBQz
6pQvbzo5QcYRRZrT8N4Hi7WE8mIkx+KjmYBY0dHTzuKdz92WrBIekV1bl9Bpfrcz
0jj9Jq5zBmeE47o/m11cGRQWuBT9a+HuCCxpRR1VkaNLoTMDhJrZ6I6OeHE93ZgA
AF10wQe1aFDRwRN9JJS/3bDMaqZ1qBubthTV/RQlI7r9bDUNYp1aRSAmaBZBhmCA
0aTsAQ+wMCTdqZJaWiH1wJ2Rj3IkSnJotUOz3gBNu0JyD97M/O0tZkKKcS9g/CYW
pg86n8y4V6GIehEr1e0tZT9CvXK1jPrAx1BNf9kTiCRWSk/Stvr2I1lUKMxLoFbm
azJFJRJ8iUfYJxZrP0srBVqsWO0QsBs53hu+GyVVypQKo7bPMeLxt2gxbxT0RW5j
7KSt0CPh0qcQYKq40/+wBre99CTxZWTBo859xaRIISYeMIgq6DOmibOgz6RUKrOa
ixjvAlRKhj2QAux2y+gqn+Z+RVNvCzdnotDX34eWMUU3xZ/3vt17+VJ+RJ8IiJeS
CZsVmwQ/NI0hJ/Sw4imAEO2vLa7lOULt21PUk9E5Ki+rzRDsf9pCQKqlmFGCI3j2
PtyIR7oC+5Hvh79vy0PHalx8dFADrdbbKGhq/GRu+TNDUVTu/ctWeI2q0DwfZM4y
ZBeq6ihJJ4La3lDOWt0aS/V6VzSs8SrUinrppbTcT8zrnqxxKeOqH8fT7UWC+Wd6
N2FtRyTX2rifMUON0ZBdAYu++VSBCwyR8wzEI4wNWfHVEzcfiKZ5OgienSQ5JlWc
EDs4COYXKWzDYzSmsuTbjKEYXdqCv6lW/M/XmI+C77QMizws6hoEiu65Sw31n/X0
OK1Lszf4wNYtYKHkvDS78yydmzYwmTUXmNANT+1VVS2ELX37oLRAie+lVGlJp9N1
R6iInjGmLLluKXFTzm6wWnDcvmk5KfCe/1Fmyg+Kq/1HvykrJslUEseKd/BJwGt7
E9ckMvI0a/VxpSRwHYDtFlUOmFUFISkm9fLHW1NldBV1fnQrO7nbE7tqx7+j8H2L
9wGoEeDUEL4VE6VwRpOVEn3nvWTZW0VfZAIMRTVUo7V26Sft2M0hQMzYu8wOlj0o
nQkpi+GNXYtomI6xqQdqwwQdlBjam3QnqRsn8KtgOxDvFUKHW3bVTqZVjz/mOOPt
+jOvN/IIn4q/09pk8nAGIkJSnWHBcGySNXzDhYA86LrpERdaC2EMEz9O6/C9sTUU
3c+n91SVu6BWMN7FONT/Wz+BJOuackWfB2C2rLNl/uzvElGnT2Djjns21aDcKe2o
sGb9BHfTwa81wMMdFLHL/yhdqR7ZppUcn0p9oEtAkCiLJ9vVX2Vd645k4MdWCPDN
zXIjCmqpt96ivp1vmd2jl4Z5IFiP/6EKqkKIGRTdOaXcFJ2EGxzLfdi90MgClEUP
WSlf/uwUqssvPmba0AqEG3+liEIuMo7kPGS2Wu0DRGtKypwCi29UYEv0PdI+GqWz
dPr4q9eCgZ39HTGIsD0kkDMAxh8TIDloHjyl5mYD6EpCj98B/DwZ6ZR442PNemqO
NyHwT3MJa9qNYJYZ1PLP8mVOsJtlsc1RIsbFp/siY/UtXdiS9UzF0EjQrwaumSCp
ANm7UICILmvLZrUk9rWeiKfv+enJAbz1hi+UxC669PvNhjZej8UeLM/vjaHldjkh
1YtvyNMg9f0aQYjghUftLlUz8r1W8hIw2WWd/+LXbNt/Nsu2FvPJEZfjbRIOUdgs
roxVOahqyhx0BLxwRR2dTrxfKIqT2LD4glMKkpnwEhLs4HPjLXZiB2ksricb/dKC
hgGcq25HBSPRa1Yu8xJPPy53jG0ZdBtCoRVv/mQGtZTP1ZZGy+uKISoVSmrxwMns
hrnkKLCVupPOhAX7Npx/LAZ09tl2AGjeGK5BT3s7HDGs8OVCUo+Xjm2Gu4HnXayt
D/UYtZK3/ID7L9IDn0EoH78QNVKGZ+SepkgKbpRJujggbOQZZGRxFaG+3qddM71s
t9kShw2x9cf52fJ5dJdC9Usl2rJwsGgu/wCo9bRfrXgZsQeCNTguhDgMcdGyQMuc
RNGYOsiMYdT+G4F2GDk0Y82GhzExpkINUXbBbH9Km3jWRFGIJiQYCLPLoXg3Q+Cf
tq0610+sypKiTr9GjGuW8q6QteWMncPs7y0P+rYWl4/LKrN+7EjHa59eBqZt7Iqd
dD2bGCgbOkxzWQDJMaUuBDbVWeRlcJjDiy599UsTaswPuJImo3C9K5cwmaorD0L7
3opz1FcTrkOVH8LiSJuI8jAS0fTohPe0qgtIgvDm1V1MBsRTaqGkmIbz/RHdQFa/
63HH/6Sv7NH+55/BQAd7IdFDvODkMpfR4woj/yoSVRdTUttP+Hvjz+7j0Ue/ysPW
rCkdaOlhW3pPLx7n0fqHGaQ3Mro95nkqUhiPBmmvowQ7ALdHY1jIbSRfh/yhCvnZ
9ZtaUxd8yBv0K//wxwZORYszAwkMrKKP05W/ajs5/q1ef06vyL9MJVts/8vPXLoW
6nZv32/3blJ4juWSWyidCJ/M3GtWJcZINdSSzeKEh/K7kgGlKx+zUEvkxHPXvd5A
juzX50Q/RGegOalNYVbQ5iTHFBTv09iwlV3ur0B0EkXiZPYrKcnF6P5ewvvsV6G1
GN+J05RgZr7+1guNaYDGiR6F6Dd2gUDVj0HWy8GmCpDs7XMMdxpBPJv2OogQ5u1A
h6YtklgiWH0S2DCrBTwGF3AO5JRQJknf90N32ptXvJ9GrmVHZXIRw+WCcQ8oNMkN
+G7GV79lgrZqIOw2srOjL/vLO0cpsg2fijXZ9dPNHKLKpdFcAg0zDN7Ju4A3/Xs3
aw/f6n3KJqQtSw0Oh9CldmA+Te3DHnNsGsEqH+OtBnaLJzGvbDayN+TITJaGB76M
YH30sFlt2liR9ZzoryUb7BQbPMk1Iyyo6IYSICNLetAjyR+TxDKsJMmdHeZAkPUN
3vHOUOKLO2MbcyHHzL4f4/5j6A/UQmbSUahMSRG6RYR35Zbl7HTSEeTQJqSC/5g+
b41tw+a1u4xZRdL0SVg7BJQNZycFgEXgzFLI13m1iPuou9E10ttltYlTQb5WmSV4
IsILXpNX6ouhkFYngUJ0pK5W1D9hYbh3uUu6CDl+ySx5O+z5L7eNFNrf+/N9abhc
WXFy+9ZddPju7rdLfOuT1wPpXsJu8BChoAI7c5mULgROhbVja1RwvpibZs/ajVOr
4p6V5niNPwWS/rGubX6LTwWjkmbsXLMqt8n9LsH45t0ovBXME9O9cUbIzj2sHM4u
AGVtPU0xa7ZRyMGwJ1dVsvZt2VL3SBKouBcICmKTgjDVspJLXBDGYdkE1V2YEzYk
tZHAoYzDZuxRH+8upZACxExrW/jVBPr8a/2rC818HsOElFi9XeNTh7HdNYOjae6M
bEHWyjIWh2o/bzNyJEfagep7qnNDJO3IrkAppXy7Vs+aK3TYHNwUUXqER1uBxwpd
XyfjsXEMVzrFGEjclXu/OzK1GDU1Av3oLomdnNy/VBbpdl3hvUI7RDelZiwhqTu9
vBtvRTVrDPvpXRNFEpaNe6mwf8n8iR8x5oaTt28j6hz4jlpRdMP8dN95Z90zqxh0
UREqrUf2S99tdHPYjkPe/DQY+o0LW5iT/QTk+D+BptbiGex0gVq8F5LCPQTWeMzs
KrnG0xorjpmDQsDdrnM5TINki/Vztg5WapCmnim3zJArpOG/DgyStL9SK0V9scot
ca6ghDIuVb4bEIfAwT08beLk0Sc9i9ZlwkFXd92dRWrrCBjRdM/eLANFpogCzq1Y
FXeOYCnA3XyCHAYI8JKhbAy/J/0apPAd7dbTxEuz0xyBNQyqr9CuIJx7g4UyyJeq
hIqz/IezFhKVACmNV7zP5apDlMfpTWPT4bWqFDDtAZ7dIMhexzrOOXxqSKNyhfDQ
LZyH7Jhb5v0futhEovogBziLVU6E5pKH6VSO/XBK8C5Ym8WasO2f0cjI3w5zNNGY
+AP5oj7MUmxtNtWcqwlum2ps8/pRs+T7J/8fKzE4vC0/vDT0A3y1aUxdHxG02tbm
JMFLL4kL9mmqx7qP5u1HC40RsA9qe0bPf3yO3tfseKmGBfEGLCEdWHC5Rm0MvYoC
2r6icvgoD9Ksn8UwblXB48tYRpQAwxyLLkIIE+3oT89rtM5Zrmx32H70N64rM0El
3dXWThmQhfpsb953XREeNdeLg5UhojDaeGtj3cYGZyltMooQU599V9M/SmjcD07U
HrXfQ4N+WZ+Q+gnPBSw+NDjrtHUFymBnwhV7UBJozDJwGR4famye9sv/0aKBgPLf
yh/R9NXDyDEZc3mCpaEQAep1pGsjo9u+6UVaMFXkN7TNycG4VPJxhtAPmyRJqkD0
O90QTYeMD3G0cREFT27/kyRZRwx1iUqDm00BSDJXnymLD10AXrBkyLauH68rAKcY
0H9ODPnKIJv27ibPEdlNMcwSNkImcuKsvz4nCdiEpJnEahOArFPEeh6JfDeI95dC
FO5E1RUj72NofSb0HnCw9r74UYNcqiMraRZIbXGMrjpKLHbxSzS4wJTWdMxq38Kx
XwOgC2T0zbI/P+zuys96fpTNorf3Ef9BZt/Ub+o2bX+fCQ3qu2z/lW7EDgvudind
Vh9E35xUnw/G3iTtg8Ud38xePf4MoxZ7ZyAvdBFFhu4vS9gEjB+UOfFMQBhj9Fsx
0e2WAmPow/or47gjgRz/OOKiSPGuZJwfq1CqFSuLaY8sxFb/D7R1eQWJ3nWOkljL
UEP7yvZFo5aGmN7dIQKXDUuhZIua3d/5C8QDLRW/Z2csHFYSv+n9MlJ+Ej+fPTGU
yr4RcQ61jyFUnBrBqzMQqOWNVRCDuenm4BqtSgEMFIGNvXqfbG51b2oCr2U0JvcK
HAsklKrBr6Li36Xg+RkfxDnWILU85b99v+7rQl4teVlKnidwSRKH4hpjHloUR9SZ
1KE83BOQQiyh85QtkQXhVCP6K1bGeiad+OVlIFb/u5JOJwtKiYUXGY/QUzhcGIfC
+DDp45zdSSGzCaAiLfAqsEqieo9cxLyyzoOJ5JLjdUeYdLB47VKLQ2LF35cKJSba
LRuAQJPtGRQhCdmYjHuRBs9Ra6f9Hg1CR3MVx0iFsptpZPXIziMkXiImCPmZhpib
6vUnIzZ/1SWwn9N+KBkWwxw6cvCgCEq8RbJNZnBpSCEV0oQISS7aNMg2uzIzttA+
vu/zvedGyjEZHYwcUEpF2xSN1b+RA7wLBguAMRY803RhB6PKIdhdcBZR63YVU1Gf
GTx3SosUYefYaARl3AhwwHYq7+URLUfv8tiqNjXpMN2sPQAitL0yJDsEBOC/pjzb
tEC+/ft1PWxK3oW6jqZCuUdUdfw1zQjtl26t0YKqWUXYojG8f0RP7zCX7LUKuwUv
UBaKYYmf0K6xul0VJrDErz5trXY3FneY+sazgLUlf2gAeAt/+HU+A7Dl0DJnaI+q
omo6u1f7JO4MRSjZHdBMna5mbAmYh0JF6v5Pn1ECPZGEYZ2mIlmTVpaNL2pygHWr
S6wdd1QJxtKiDCDGQuzGeJttsjkzdHuEKlEdqXzjHhjf6mfBTy5nwEc5Ml97IfYD
oNO+SGlYlrF5HEwzF2hAUsFo0a/rMC97ILa84q27Jd+dZBnr6teZRuQf7m1JtLkl
7Z1ApWHWgFpXK59i7CHYEym3TYHKZZlnhD2RuVS4BJ3G0+LRMN/idLb66yKLgCJM
dTKeD89/XChCVQwF60AM2oVrqxfz/XA5fDIUghCzIaE68kCT93rkPekih04u2BDt
Uyyhnn2GyWKr03T9GBN230f/t8ZvnS/iEmhjaAX+CsoyRszmr7QZHqVIQyDhk1ly
/DX6feTVTrjwIvb2bcP79drLWH7oTc5CWpGdG8gNOBOHzTuiD7CI9MdgX+W3vGH8
zhfMr2bkS6wwWZJ9xNv/tFOyR9rfrpT1f2w/TnFWpKQ+A8Tx6E+C7K4R9s67w2Xp
MNhudngzAJJ1fYfMMwUgONpXdLWYruoOlk2hRchwddaRLFBDJjF9p8hEtEg0QjHz
xqgXzME1WcxZi4F8++oX7iDvTqPi5XMx6BQ1vIer2X6g7NnM06SYE6XT2XA2ByXS
5pFVyvf1u4Qc1doSa3v0OFJh2OkrETWg2HxKi/gKmxXp60d/AC+1hSluYQiIYm85
mPhDDUTq7rpxMaYAjAJArB1load8n87WmWRIATSx51q7SPR0UWLUteriYEn8CmKn
H+IyRgBRaPLK3US0wX532kGTd/f6e8cC4kk8nyrAWr5vriiO3EBu40dMSCPF3qfy
TSSdPhtGq3mGittBqs4ROD8iiBKc5FDtTz9Wkw924N+RiODvfqRiiVmKo1QvLKFu
DGwdvpOvBv6RK5qIWkC4RfLndpcTjf+FzgOglkaV+PjgnIrbBb0TUXlVB79Rs76q
BzLYaXkSyE7ouox2MgTj6qU87QSPiQ0iXshm+0rkZDnILJ1mElzViQ5bivkRDrOe
2I6EIe3yxC/b9NuLT/0Fjs7AiqcOnwxJkRh9yYy2DsYFb/V0OtgaI8jZzTWBjnAh
0OGdofOI7KuxlGYRTkxzwdW7dEOuZVDtIrM6MAHX8ZqgyShT5l/tsBueTkPdBZew
jC5jaGLdsL1J0xbvfUa8M9nyQcodoGIL2zAIp2mH3iJ+7YQICwFCpyrdAppMUr3T
MX72VoYHrY155UHP2R1CC8UZwQhElcG0ndXNRyQg+9vas6uvpGlrHXsUnRFWvFPU
mi4AudIwT0i+orouVn+zr+sobae6zowJmZplk/M2as+r24dW/VK4GAuaP2uZOnBO
GSCgRyuKnszBuwJA7BQpzRlRW3dfiRlGr3oMbk02uJp4Fa56SJKu4dzfaTuUMtxw
S0YdIQO8wacgWziyYLtczBtvA2kErFTyiNpJkRqurmei61ERhTzqHbcVfCMGiZND
mEyLYf5yR8y5vIkykddQp94O/zEiiZ5P9qgMmeTl14Z1S/CMx7UXLvLxGDP4U5zY
4MgmEhKOGW97VyUB/xFTFRa7svq5kSpPomDEmXDyYem8hoN60KTLWA72S+3sphgN
diBmdD0CCngYWhGC0MJTm5QzcrNiiT1u3lDVrqCnDiDBPofX4I/Z9p0U1QTpDFX6
XTJHZpP56NJjy9qoK10etmMKws3rw+LGiIQljjCxngC6c2iXOcVc0XKYjgJTe5H0
dL3DPPEcT/R2DAIQoHlnEYzF/hvPGOjlO53tKKOdxSuZlVO0exsxFNmTJGIEl5t2
Wia0ZMoB+aAkdT7w5YfKMZpetTqkOqo5i9n8bXZzOdPHS4Qkla73gFy450mW2jSP
c/YhQm3AIt45Y2jL9uaT13iQzlkoQrvo11dULcfCEp9VnjrKpCA7odIURiNHn6eX
fbWukVa1x94m396t1wK7MoGMMRmB42hquANwI0y8vhMKBNHUIIjHmX3wlQfAUcTK
SL9xlvRccQIfSBj1rz6xwWsTeHbABP7q2GYwcUom0auek5wv2yvyAMJ5aZjO+kHS
+3Fqm7I0F+Zvef4ejlivJGLUAm9/5zTBNOG5MDP/ESm9NI3+RSegHRwDwwi6yEut
yWoWoHcOiwft1194urMs5jXQY5Gg5qwC47nwqonEBmnBLVvfGBR2f+Q79jrHbW0C
X5ibSCICFYTFMpCKQxcqzchmzmaoAHQXP50Pb/zyHOjfGTMbJ36M3kduK4UGRDvZ
q0QSEwwTUbJiHR9indcPunInYQGdP6kK4vc4lUZbWxpDcOxuTBUxYnVrThtvUkmP
KSYm7yF5E2uw8wEL35qQccxqutJdiW4O2BvhbNZ7AJARLrQjkfVSeNSzEvkc/gUB
A/BWEJe2Sh1CeaR/qiTblKR2Q04MK5BlUG8Xqgf3Csq/QbizLHNcGod5SZyL1V3h
sIdnC270oXeCZbs5IfPhwjDOJPRWySVvJLiCnGzzYmWIGy/Po3410mWJsPPb2fo4
JddIDYoFiAK6HGU4rMPTdEjY8B86IJDLtC0NBga3fyFZiUEhb1NHTn0dAN3s8IR8
q2zhOmjPQQuNn/9BlD1zMKULhw7+AOD0P/IQQJCtyXqIIinjJ8jmi59+sy5VLe9u
ye15e63sorWWAjxq14C+UPJfAVcpRYUVJno5l1efiC1CN/QRsxGwWUky7mSYPVHb
XgO6LJMOw936E9rs6bk1eB0p0vmuz4ICNcPk8XmsEODRRF3mLcuiXh4sjDFIh/C9
BqAtWADJgbodewWdlP+AOwe/2wKaFnI4cHOgs6alQLRaFkfu0vmGtOTPhREvKq3Y
eGncHTvFHytTiwHFZ9jxBCBEeqOXRMoeFBeiHNQI/IZSUWgEuVOcBnlGM53nu1yy
KNDDu0kfn3FxSaP9rmZKkLA5Wxs+2MkorwF5h0mcXe1JSoEJiHELP9T1fRElJ1TU
iE+Q7HbxqCHKl08ELpFEX10B/p8y1fSJFwchIvxmF8sZ/RPl7MS2ij2IowKVhyPc
4XlwCqjN6h5x2VBJ6A5KQxbP7kVuX3RhmvkFdDtUpJn9uoI3oHSxutCmwteyVEe7
63m26K21dVZEiRqQqo0Lig2vq0TcOzpDjsi2ZmLtj3++uQ6RwnDn+Sknw3tOkgnG
gYPuUsC1PX49EvLVTazhJNsuRvyUMFjKXqahUnx/X51YQVBAeBfY0zxhuxq8zXgg
ayBW+M5LwiaGICNJkHiv9J67d5QKf381oagaVZ6gKCYiynAj4ERPJ/jEuoultZMM
1F46Tfbsgl5/p+KSunIOVQbCCwQCTV+ubxb7i+69OEYzsDWWllRoxVhW/nKiWE0G
LAbHoBzc4VrAUNYFYYey4UuJA1fuBdLOHIXH7p/01VeVYjp/6gY82dnllh3NiDSd
XCY8NOxEzxVm7o6t7vXkqS2TWRWzjkmNDHV65vTgus4Mm4TOZDTYbVxseIbtfN4B
++iFGCcKcXnpMmH7bwen4wflPGKo6BvdMrkLuihsdvUx8AZ5HPm4Hi3WHueYJlpD
FAzDB7LDKuMr+9boHoyzZZ48WpUMcRMJlqD/ISODaUcxyczhKGKdqpIUOLl5utEC
OUm91QwMVMzEPZ7hs/+F1bEn53cU6MDPP28qlSYWmybltw1IdNlvZqjCqwyJ+y9v
bGoiCNp+1b1DQRytaiN768AnL6hAMlYBpvUxwRN00FsGHeMpDJDzRPvobckdVUHN
PdYlRjyA13QNk2gF9G5xDasfl9n2olBJ1g6BAM7UZ0/yLSe6onM6p/zvusNtvvkV
W4q8TjDQykHU2tf7VQOtiUxWzfTpqCZY7AP9eDby4/2IGolgaq3Ymd4pHI+aYnOF
tGDzHyvKm9O0S1Ra7pwsr278+CMen0fV+6YbBqLWVrR2FGO+yLcBLkpwvhpxL2ha
1f1MLSof2tZ3DEDgK4zTimhq+jyMsZjLfyN3pGaxeEq2Fj0QqENLi9oBYaDjztzF
/xv6FfDwVovbLnhpMtQWfyPkeQzWBnYCk9/eSUysp9MQFVvUumF9bihV/g7iHZyM
2HsJJNAOOJeXt+dnDluGFYpFQ52CrKj17Qh2uupGguRFH/1PHVXLzj6CWOqy5uAW
ZgtPdlRbdsxglzjDawAK8064hyX4CD/crjnlRv0LGKB5NQTHnb8HAVq0VUELWEY1
WaS+Gx0sVizrS/cbJYPtzyEIPD34J9VYPEh8GRhzI9itqURWNkHucZ297l7ytxeA
Ijva2HkW0o/RuQrA/h7FxQ7OpCaTthm+HH5tE4P55oN+4+4J0z55XMb9ZHuq4iEd
V457l4VKFwyTUYENgL27X1pnNDflOcYGzn2iyWIyG+9jEF6VY4SZ+aFZqcxAiTEA
DDslK33LAcOYNqRl5gAtrxqN8e65qndd8Xp4WnBvTSMVX9gN/dTdAl+g26h4MRyJ
z1oHRuCXlhg9DtbL2Te2N08zY0T0l7d3/oypDECgran/NLrlFPVW7sa0puOIyJVo
/W0+IVzLiieztSTdWpeEK0GWhKJ9Ub5uF1z3MzpDg9GtGB5sTw9XjjmBKO+osO0R
OgXnf1zZX9Sb9NAjCFYvYqGTqCJ7MJO57h9oR4EFrbKPWAawo7KrrLJdV40HFo0p
ah8pAnHnA3KeeQjuyiQLwAy1OqYrNyKi6L/zqHUY+DKl8RgtovXfPOdrTQYDnF0T
F7KMegtei85HHoh5jvNzIx+Z+aszO3g9CmsXEhuB3PHUNX6rtJ+QoWp0BVMMxPQX
1j9i7BLW4TU8EnW3awLw59XG6M7btg+eIjLgTyecgaabQu6xNTZreAiqN9AYEROH
chh2VhdZJBRKvO/CBEK5szPmGvqctpB+QWGk/6r2JbtZuUkySQmwSn1nRBev03nJ
AzCoSlzg1ENmHpNoau07dGvbPXDif60LEIK5f8KGq6lVP8EZ/bbu9BhKR3GeH/vZ
G3Z+zmpijGD/wQ1auqrEa5NakBmBtc58fjDy7WUaKeBv39ZkgqoJqOhTxbPlttia
86wEr72nBF6GGlHzvX3LyC2+w05rmeyeZiFmwJFC+rsVOrn1tjRlKELT5gl69+Lf
t/kVxIH2+DoAeGqeOC27NHffDRCtGAXqKRZi5RGcsfQgFqGrSg5J1BN1v7uJtZoJ
LX6ZoIFhG9vzWMaukiyXzXPSw+epZLVmaY9rDLhDC2GSQJg6IHJZ48zTEtlAF1wB
Gteym/vqHfPPyLlZ4ivcn+XJHU89I2YSO/UwfvCaAWYFQtlSxHrGoivfTH7XiP8Z
5X1DlKXZe6m5o4Vmb0dkW5BGW8lkw9LuYQOgn6OL9QQgqZ8LvSkEiuHNk6SDiIz1
8sLW3Bxu+ZWTnKBWR2w6jBV2bOIylW464N/h5UJgK0cD624o6O4tgeJc/IuNvtCg
YreHRrge23vWzmXzrQmxZPFRpV7CaTUQXE4rpi4lbo4lGyaV9bPXF5Nm/sBsDkwV
3qa+naAtc3aeV2ujsQL3JWqDuw1X5o9VrtRnDMCDidiVl3c0aW0Ek4RavKP/MHpW
Tt5nbHEdBnKjBURvs6zH+QvMW7Z31T48QlRbrOk2neNzP2omxFzX8uTkKQgFyrEi
qFhFWtwdQAXxxQ2FlvCks/BeXfFS/dEp9G0ZaC1FAhgG5x84hc9S3anjLWVdellY
NyQlX+9Z1gL5O3Th1NaUU2+6aakusnTEyeLmWcUWewjhdqoko170hw0RV8yxt1rz
WTWRlaZG42JAzoD/PRMtphu2xsBCJYgLhVzVH4+lIVxCI6Bj6NtxnuWkxSqzu+e1
jpHfl9Io6dd9YcfZ9qGOg4hsuuaylsywicU1RhUW6eph3RXmEIKDPtnRblcOEHhd
+6j0Qat4WHz+FDNJbCTQcCPtgiedo5bW3ujhYsf8Zxj0xfmW2lC6t7vUOckQ2BlJ
rf4Syi43y9QUeJ0AbX5xdcEqrAiLrNnE3li9p8XFX+ki7wKanl8kcvqgC8YnV8md
W1iZbn7o+rSNvnPBUDfcDu2DWadRCjcHAXY4yPwVgdjfQ0OwLhLG/qMBkfn8qju4
dVaB+YTOs40/+SD16so7eMn7sphvzFLgWxL4lEUyhPHT8CGtTVx2DwZvOII7AeI4
eMDrv/9FVrA2a2HdaADjEbo1aay21XRyIEYwdPDWLvRwcqnNryBjHszUcTs67WOM
BBdlegrI8ynrBgdEsaVCqA9590RUfY4al8BbZtoxsk0=
`protect END_PROTECTED
