`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E2iMnbAIajGo4YWUcVGQ2xqYn04D2SVaoW0ghASUwOpUfsjYWkWzcPvga6F+YkOX
GYSFgcDUzPzU+FzvnRMVtFk7dZNLQM6fYhDupJYFrmMGHmhnoU/Ul5vZBbmy/wIC
cIY57ET6ivbpTzw17YYrj/v3dfe1sVekuGaP99jLGCOmBVP2UZRfmWwf3p0ZS6r3
an+bqtyGFzuF7M3DQbAZhkLawWsD56b/21GZ4rtQrviKNy6iidvnMjRbwUwxJDdW
l7oQd0NzuWdcxXlU14WBQg==
`protect END_PROTECTED
