`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T2EBQlfgzKqVOoT88f325JwHAPkO9WKbt9Lx4jLpDRXiS4kxGJP1XNceo9yECyTN
zBqlZ8/u/mtt3XIvCoiTXoIxhRrfU753oYoFxVrqN7/7r/y/4SSjavLQ2GiHqsHN
85Wx2JlU01dBbkjgyPia6+YhAXZ355i9BIbjKcEk024PxdMl7W7k+QVaJKV4x5xF
sr26kkvv3ttuvWh8rs01di2tOrCpGSnPCkS1LRwj7Ebqgh61u1+q+Mx5Hz3q2l58
VxsOCZAORWuZ+WWqCopo1P4JOJC83fZwGNfPtkew7faOo0uewwDBzmVHXYccgrN6
3sC18cDzi7Gg4XcOXy+SShXDnbzb6hcvkp1GR547l7CP5NnqW6akBfuB+KIuZ0Mk
ccFrxjsCjX5WqjSw7s+MoR5fEhkE8Ihe4gknHZ45f/nWObiS7Iz4cJ/qA6zm0l51
l5OgXOsvJ1mBdT4+t+zUwrZIVDVaM8RCIoO769hdR3DWUSDMGDskZoPg94E2GVZE
fl88lqGrucULenD9l7l3pYQhGjhqK9JYM/YFlA/5Ix1fg3Z4sQ+vnr3AFFAOq1YA
88AQGNi49EONLxcFE35xbx85BblvtVevkZ/W+1OWZdYxOlA3vzkL4F14QvR5aOIa
g+IMvsm3E6P79o1T9yfTxYv1dOXRzH0xiSTmOlrgtgRXJ1wmFGtqqt3zt5qX0p6O
++gIG21ZEQiKMDIdcf4yi4O4wg2HIFi/OQNNXXL17SlswGOhqzrmQkdIYxEO/QnY
6cfudACMrqvRze8IRfNyeUUxH1ml0vo8pnmwK/htN/mPIB6R6tmTgjd3xYUEzmWY
QfuX3UD7OvUhb6R9cUaDTlbydNm4x1VhhFdm87Bvso++Cww/Gy0+Q44sxHj4Wseo
C+z6tvS+TL9WJq+bGa4VVODRNS1sLYGMXjuV0sQ6R+KEXPBMTGT0UA2TpevBODfp
UjDoeCmqdt4XcdS+S+ISwUskgOIH4HFVAM9yOBn5fZyCkx3SHPuuBFRygjlXSeU0
M5djmItWIqvJNbkXF6312YZfSgWNFR1SmLhoGazHqw4EonoxepUYEYegjw6HBUvd
ZHdlU12JK3Xfzga+lHzCLh2lQJ9z5xhoOiWBzC5GkY92LpHX4W9QMZ6k+J+if1tv
zerc/Zae3LfVpo1wq7gx9G0JCoAruH7i8IDYT9wmashD7iTU0gvOAFEZLWsArj5b
ZtM7NIt8cR//oTi46CHuaUnoUVh8bGTnaH/QAl2m4fZHU+HgB1gfDKaA5P/9DwFB
`protect END_PROTECTED
