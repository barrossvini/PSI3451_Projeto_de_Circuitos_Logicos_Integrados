`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kW7xvM/GpoVu6Jz0yOV2mA3P1yMRn7K1iQbU5cVrjS58rLYzG5X05iEM1/gr/USS
y6/thhKsIncmzWBvPUc0MnC2M10PCA8FEGiZhZ87HSXMSufnISNO9l6bSp9qD73R
Jgrs9pzRWLxhvHR44EmMZjQdLw4bvWStMYsUZS90XWFW60G5vExn2VsavwgXQjKH
iNmcWWsrRWhDeCVXEGqDF7rduhKKBMqYcTrM8l1cI3uueA55H2XLgx72nnxT1Lqa
4trl5ak4IyZKvbASNMo5bu99n3uC7sNnB7jL7nbt6e8Zbc1UamHHA+mR4epdiA76
OAzqnoQl5zcPYWH4TwVz8tZZCxI8QcpWJrWQ2RM8Ox1qfi67+tT4ngDjqjeY6zsN
Ns0D8Vs0RYWhiLVoGPEKgWwFqGqebni4i1hVQfFn7DfT6Qd5C3depSKsBo0ud5GD
V2/QYkCW/3AqTll9c2SAdFtseprnzQuahesuk2Jk3uYwWSpWVFVJzOz0k1MFexNZ
VN0rEgDqIfhoSdleeWQFDlMpKBf72SCjFPu70oEHqPHpa59MZm2IgWXs4tEDU4Su
f06btfvdC8oebYK03XS9FujClSiGpsxMfBQ3AlUjxokzX2/eaeRDd0f/uVE1i54D
ykpdJ4O/9EXTntRRiP8+WfKLz7FIRqKW0E4N3WIXfN+kdMCyxZVYKj5vOathZZ3A
CJOiEq3qkq/LjL9XiHaa2VwgVA9Yz5/N6A/52UIriB73titMpPWlIqhLrv9at4ag
rrqwuUPcXEthF5YRCiToxLvcEMhS4px7PlUpd+vfs1+nkSDv7eT8DNYc3cCHLa1B
zmMuw40QNCJoMos7VYlglk89ibWKRikYFlSeeaVAD8P+W4/YkeT5Ws7MxZt1jZKl
lxQa/LwqlnlWwEpEKIhb2CNvTewGIlcW82Ge0vkS47czR6p5QvJCXuOcoVxeBFIR
S/AavwIr3crejvdHb1jbvi+uW1MLEyTvZJ/IovumbMNK/t+PvFdVGlIP/PuSuiIo
cFIMvVi2891F2jY1RJL0IODYk+Ary3RGf7D9IBcZsgi5XAiH4PHjh325YMm5M2UO
y2q/Yrmp0rprNbxfgFfMlaxDjwcDdOhLzM3CsZYA+VajM/J3cVSxGpMyIa1K82Dp
k9CzM+4OhmDos0FaiJv4Va09jhuA4TMTAJrZd/d1AhME1G0f97NYW/3Kn4G+71sf
/YLM8VkMFdxcY3L0mBapvpo6vaZDl7s1PI/r2alScOddr2tLR0gYUtG1zvET1nGD
s6yjRvCJNPYm/trCPPVLSycEQ2zBWDOigdMQY2pLhE+rZWUDd2H3bYg+DJpXg35E
N+MUfyYFpSWVu3oTtoYLjQeg1MeaFpE//+Rgiln9IbPI09P/H3Z9VBwsDFCIwvwQ
PlUSs2e7YN/bmi7LEh4RnrFWr35vkWasmAQ+zm5iJoz5QYJPKOykxMuEl0skzB7u
ZdQp7cmH9WTBth1dAikbKb/lYdfhLWqeC8UstvtHFHlswkNG5ErM8k/f0bqj1ND3
597iHZKYx6gLIbT2Be91SOEDgfKAAnyMCKyqnC3SgVTkjlpAd2wAvKerv3RsKMtA
1gUTOtPwNyph3R7qj1+hPHP4kF4CFy6+4ponB9rz8A4CWXLQTEbXgEkNLTwrniid
1oeoL4JjFWyPtyeGgSmWukzeWgUonZ+31s0GjasOnMqZN07xaf4U4BWY7D5evzwj
qjP9hCRpnI/yH4Ns8J4F3No6OCtjPN9Zgvn6pHiKUdSJH+brfFBUKY2qmm38tZDI
`protect END_PROTECTED
