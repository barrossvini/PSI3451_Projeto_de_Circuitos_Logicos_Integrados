`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wNf5FiLAAeelebqjQB0Ad9m0JOrBndP15PBHqHoZgwRXqcr7cxfDAv9lxByABu+C
F9lfLrjz82YMgd8k1HzHusZ4yMD+SGQab2kbhqyYbtfE9Xrk6/FicZRN9AJIYouD
qqy6k3wiZVgWb0cIae0yvVO7WGCtcbJj90t5c3qyfRa4LBf53cfHghBq0iEv5f2F
ph6YmfFdQh/LSwysNMXuMSwNvRK/wfML69Sl6bQ9a9zmh8DVWrOXNWZ3Yr+HF4OK
L5jiDDqtNqbc583eaXsTSLWWrqFapp21rbm38AlPyGN/UVvq5Djtw4JUjJgeZXqq
/kS0rvGkzWRHCVg3bFLNyHKIgP+fxDx8xIfLLnWnCs+9qR8Fs4xdhPTWxvSDYY8D
iOleLshz45a+/iUTRDcYgb/sJ4xOgpC6f+1r2C/lMmklqs/9FMS4fRCN5ZnUgT/N
g/myCW02mP2WnqmouVwtEBXOpPweVtIWK/wCcFPX3VjWNgfnyeQQuyH//docgqmO
i8DZYpn792lnh1uHbDHwsD5183DPRJCg/BOZ9BoZU5S7qvCFehPBBj6IftZTr4ud
S+a8uKq7z6BoShOr4aBe+F0gJCdxYvvOLQTcxmNetTh3ORgeGAqyuRwxiudF0m/W
v2yo67nUJWEKxqMJXldmPqr8PJlQQOcytRjkuCIZdqWx6y5LHqB8qdqcYdiLiiOx
m1MGG4F5yMFt0ki24YdTQh0EQnXRvWq4Aj227UhOqy7Wq754tKBIX2jRIXdqDGSe
HcomW6++rqqVCCiOzpfgkH7WocH1swp+Aq9VRUephydBdzut8+edYlF6wIfGwQwS
VF47CC3nRePB7D80WrKMnA==
`protect END_PROTECTED
