`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
604kB6/gib3vs6AXQViSO6a9+/TmaekWjig2aOqYFZA+bSOCVbNCZn/sP8KSD3Z1
BTVX9gWCSmJ9TJf2MTiB+rq2TR4Z5iCLHMe8X8ZJMJUmIVZHxJuKDq6JjlAYUif6
oz6hy5VoMa42beBB2H/HAdALQVJGY2EE7sawQU3HLZDNIUVydAtD7IAL14czQSVS
TMlBWm5KVfnfi6VJ3bR9Znz4sVPEBpb7A5ijq4oEylERCIKoi1yBJT5UcgY7x5R5
RMfOI9MiDRcdUWZusXPt3deSc+T/mssfDmbZQYVoFfhv/4gsZKcnSXuG4Ejt5+1l
7IH/nVZZK8xKaHIrq1RJakCabkT9vs/UO2l+s5Vbv3BReu56IURmWoGYZLZDdMEi
4XtoarO1LLDNPEZy2jgbw6m1PZMCgiqUJdJOwtkKmmpc+ymUjQwI/2awJc+9uAiI
quu6bguWVcbsdDVOPdHWlNpFLwqKPnfd4tpXSQ1LWqGZGwHoOJDYe3og88evnvQv
sdEc0eJcjK2LeksoSECs/p527wSN8yJBxryvQNdSF2bflRPm1+9KLS/wVHPvTeO3
xhdrl/3sjPzi7mKk353bCbEQ2Cx5UZNg3p5XILm5T3fLbOXLhKyv8VyKD9/3zBMY
/kbCoHhkm50P5Gu70tM1FDVOTXBoO/pXau/O0Rcq7ZhZQwtZ+94iP6Lqg5orP4KD
Ky3lrBNR9SpyqN9sZY/C2bwyWnbX0HnA8lhC5nxpLNV21BF8izH6Bvf8pHGAB8cb
NKBLQMeaDCZV9+i/lxy/oMPcOm4xPIDxH9g44PU6WdSrIQyvtl7GBnvMo1ovU33s
+W3AHOsqg2IFmK78mGh6kS281XoZkZTIMZ67qaPC/37RVQypGJK62ytPwdmAa/I4
3cqeHmz3vZQ46YNiZm2SGZhXZvlgxDNblHUxZY8+AzCxBdGyW6nI4ethXlZytvir
1TFWugtgMVAXuYsW4UYxXN7myUXRe/wmAM5Arzt5SlBQFfjeg+zcRuK0fkumiACg
WtEZ9OGO8vxolpDfdntaWskarthTanYQu1oNEyaLt9K2CTByETyTvAH83UDlYfPQ
9wmJdKk3w2YZJJxzAHFCSkL1sMyCjkjgtl1/rf1vG9WKAgYIJwcH5S11awf1vdvc
Lgg5oSkuseMEkLsWuUIpmaWrXxAi7Q7u9ESbT8PrmHVjeBa4M+lGyN/thb6SnhE3
zDpF1mrw2UCthZtYASqihJuPARDOGB6qyujPoU3EcsYGy/u+r3P2LhfWss0Kjmww
51Ej+yHZt4WxOZ1qfJFPCmrwcTsBu8mZzaSVDZjp0OUNa/9rPiuOYaFS+EoDtIn1
SdH/hfl5SkYbKILjsxhlwhwTmft/PvIbGUcOMdcjJeAVv8PVO20ymYlu5l+iTM6h
/nKMNGknNQnE4kEk7laQo20mJ2CUj5LWHHEaYAH310CJJxbIWck/5hUOsrhrBW8Y
hWJMJEReWFYFT0/Yfpuu4TW9BgFMvQwlwNmlS3ww3aG4Ug4253BJWBeJVbWsjEcy
kdBuddwLbx0KJGWgGFUVlfstrTtIBdE7E1Mg3mSFTbEHjnNGihfBkMfEqk7yis5I
FfpLo1D+Y4tcOZi6lecOxefogbDId7Pq/n9Bs/ReooYxYqpIyNMzQlOrJxLOltnw
nhHU7k0VxPJkpS7sUFPhGR12+J7N0RbW66tk5F+v5hYQKjOoQt9PD6IHWhEZvjiA
EqhJ6/5+7z5wb1hvxRGLvTRsrqUSQNoIoFB53IhTSnxXoez8d9QFFEmDDB1RDLZV
mR1iE2WunW9Gb6Npoh4ANjAylLBjy/mqyByrQ9HGCzg8NX/5bcBDLZFPG1AVTA79
qSFiX6yseovn3Y74bWffZV+kK0+X5D8RSezG8RGBCCx3GEHBoB9N1laNNbpGOKh9
yw+yl1Lqa6eYjIm0LZeJQWiRaW2feZSWBczSj8ob9rIOh5+ESgCNuViGgsLItrjZ
6MF9uAL+VXgqZXCWdj/MFBFhV7YaE30XSIpJBpvBoq30OnXsecvAaN8NGB/rqyr6
1UjfhSUFMcM5itlZ9SHuRKz7+cS/Bqt3s7gQ5ygCcKsyIDHk827aIwahjofC8Mpv
TYPf4NRsSSUJI8G1NjCou3qdHLEYkCTwU373FUT2QrJBntma0ybt8QR0O9Eessl4
75UI3iU0CosQFCkECsGCR/qSIFNODIMYye0RSK/mQ/0BC/zx4JZyOtCHyGssiuky
EEUztItQh0BIV3AsPnSxVvFgcS6qMi9k44UmC87rrC5Mwh+TxAj6VSJ6opq4clUW
V5I2wqWCtTOJYEjDMhWoemmQVFv38ToRf/JNtp8WJD2V3hkz/LXzgAJOVQb3sAmG
afAX2bhdgFiYauGxmq59S6G5+LV5awoDanCaGDMMFeu1EcWUIL+wlAF+j/86sRna
WqJr/fbA/TEnfmi9pUpZuBoaMpnZNC6ddxyuu+n9ycKQfUl5wweP5b5V0O9g4ZYl
yEcdZrDEls8IZcvGcv/p8Q0d7W+z/KpA8ZrPpL9m+F4ZeQDh8eifKIHajB1oBGbh
nft3MlJFQ4yu5h4cgndbbg9jZzuZNaFg5A4Lf6xTiiOIqd3U7pb1QrCtNL4S9049
SrS+g5VWrKiNj5igdh23r9xh7LOqt/QUd4UQgKxOuYQZ1XflRKzFf499IZap56Uq
SKy69ATF6TIdAUgTxh/+eVN9fZkh5tFcSBIq5YCvguHDdtPzIa7g9VJc7osdrAXm
hsoxtOB48ciqWaRHrBUDnW/M3A8NRPAjzX78Hjo2e9HqoAPHfNfmS0grh8ANJeBI
cLmKt+7RndOlcsG+C0Ax6wRiu6LDNJNakMgjpHNlY7m7UIH5dO15XIfSA9E3Wxj7
wnBmYND5MEJaBSDcc3io+sWm4nJ2MFLPfaxRgYcn381cJH2M7WLuSf9l0dU1Jppk
9NsR2jt4w0lLHrzFwWwjbWfHz5+yecG8nr+glNDtGRDEHOxQvZXQSU6OyE+DEIGz
Cp3G2KXaVfAvzPIsEH0f3wEG59ADtTrtL3XgwnLF0ctk2PKHZwiZylmJKxr1irHq
vs4k1uzmTtrITAUCT1ogbW+cdbTcI9yBhKxecWLISay8hmmbWY78JNkwUYmbIVij
6mj/dZxwI93MQKce5p4zhlbetQdKUX5xiQ+Us0n3hq2AUS5LVgAkwJBS9mEGrSlQ
B0dHJHlFM56F9oGKpQapnxCXwKhduf/kB3LszHLI3ZPKAzAmB1HOpqAkNLWkFEQ6
dpman1GdeC2IiCrSjAra65pbsRBUjn7+C+3GcC8hpoYLqAXO1Y37YPjMeDtieKIZ
HDOrgc+TBM4RlNEvXvROO3HjPqcyqcz8H1hdhvnw0Lm4C6qV2eNdgZo6I84j1NMv
bQHxxbAhPBsewrLDxehtP4YoOY+pPNcxf6o5vGahcRg2Q6cy5lbtTxPOa1MEQsbV
iJZSTwNqkNTRu7tIWEJxn14+S7Vi3KCf0QlMed0N5Ca8AxceiroDrAQnliDrHCwN
4tdnMS6qTbeTcEDlnj8i3BYN9k77BmPvO0dr6+p36YrB6u2rvzE7MGCDiNNVvyZ8
BCPf5dOHkfSqkJonVDMbTcq1eT89PNngXNzopnY4zBa2sFwGNEc/AaXIavKhFO0J
VxLBDcWMeQo12iP8x4XYcJG4/OvafuQ1OgvHDF8ITE9lNg/noG495eYkTdZcl+ST
nJphgpkOrsbGxyAdKKGXkWHv2Po5LhJDd+hsc0320sq7+L6kahL+MF2K66IBYQOg
fY0RSNdbO3prcEDprKzydwDBHMApI0lHLENAoK7rixk0Dpb3nBI2r0LMlA40eOiP
8bO9V1ZBAQdoss6nN8PNW0d3ia6KJgcucaP1wgnMCbwV+7p/vN+/zZwCnzNfv+Wa
hMAqcgbdo2TGxwbxmvQ72++3QpCI4gHQ7RExSoKKt4/4Iqn98x/kkzv+XzQ/XAjF
saPclAwIU5tDhwpKEH6oOGBRfPX1LWZ+FGMREEFLGzfLSqpEb/x+cmUZsLpJ0ASB
fSnZbXru/+ghEBVCBJUwzpvKeL2f3e8Ur/0Mdi84JOhNke98hwZ8UZc5PjFSXe/y
BnouyOdzlzzMfN9kszdErPmc4niHCF0Yvuj6wAxKYXf5kWiqNsVLnd91d5IeMWnx
ZDb4CSS/VdJ4Kwtj6vm5fEHoN9W9+tbR2/8yO+oG7Darkw+wX4B0oxHohClfDRei
6oTBRh5BRPXdr5ly68lJ0zHusEV20MUYnOWviTWHlzAdoxJiFDqW/zYAyqoOPpAo
Fo6VOBRajCiGNRKIgPXaD/eJvcRvUpjG5XUwFjDuuWvFgzU/pzoNyL9/1+VrbWTW
FZGaxrRzSLUqhztT6lh/7FTLPNzjf9wV6wqJ6su9h6zJnOqXwPYNmv5Ag/wW5Q9T
ikNOCeGPumIgyZRjml5haRoU6loNECivUuNUCW0Zwg2zAOwfelkrTKBfXZHYFnWw
1ex863XtNfeoLBMHkzQlLFuPDkNX/EWQ5QFKViPPEqfQdwBhRHWhLtDG97KmCZir
o7l3rMI9InRcOW3FPQYD9psv94iOElODzMHpitBZ6U5udE58n5QUV9+UAqEyhv+I
lDnZ0pd8JlPf78Q6jFHpOWxEhpXqTvjkra8TmpNr7p7/kU/G+n+dwWRZZQCHogeo
mJQuSWF3SOprqD3IwLxz5yFtJXmAVJrNJ35EQ1O7hBD0V3WdDMqvaWMtfSqvygtl
uK8LiM0RH+QlhyK0ap2SM+c3dTSOqLZkuUYROs2Eycj4lb3V3KeZyqbJSjNAOw4/
9Luk+niwihz1Yc80GEbAmiJ9piuB4o0PJtuq+3RO0Kh7heuGdhf9G4eX/Pe4jVye
w6N/YRODEs25yJwut7v9aMVbfLC4xLI/jLOo+D1jKDKi+4S/z50zX5caX1/cHHKG
EQZ1Dv4SVG7QHr08az8UVVF2ICOMKM0LnYeSHgBKVz2U2yC3147dXEwIfqdEuizA
P+zImrYeq5Oi7W89pWeWWV/82B1VYSNQZbbhnESzYv95wWa58Vg67COs45BTrsA+
Thj0upvGYO2lo6+OTLOvhYRMe/vi8fJb1OsxTanJSYRNrkCfChySfUCdgfhjjlsb
U0yQ7sPHkxHh0ZUX4Rc3IcP8DZgAoDztFWJqUmf6A51PanUnGPeu3Sz/LXRyYE27
6zAxeGoS1uzWwbAu5qxvjh1GJXDMIAhHUK0oyDwk+CPoh770Z3OUeJ6I8nrEYGha
SN8sMVY4VXuOHRcQfGfXO0yn2NBm3DTNjI23+470KYXRL+F5Io53RMvWi2Z6HFDQ
ib4mpGPiAnW4gBZor/UHu5Kc0/KEmNuaqVyGVfzJkuTkTn/FYnyKPOvkSrHXCrZO
1mKvsdhtcJtCvqVCeQbY0zu/d35uqKhhuG5ds7ojM+7fsbC8O4V4SyZ47tRF79/e
5gWHfORhpd+25+BwrxphLfhIcMCkp3nWsgaFNl2U+SXCzyINQk5dkolPMWJKRSxA
x5ZWP58/ctat48nSY8ugUNY0MLguj5TYv1J5YhpVxsuZxesuFQaEGNbFU48p3yEy
S0OfOxJGKtdPwRhnXKFMUdt/yCyiJDqKYb8PhLFBfmP//NQR0T6EwGosidr2NCPW
PJ//NiO4qS5BG2FnncfkuAUGhr1BL8ShgtNnYiXIfS9mfPMkX/iB1ac+zoEAl9ku
0Ni8rCNxdOmMsZOdVZF8ULv4U/OO86iyNpobCmNitVtFq3E1pnX2oOggqV4MnYeE
9PmUhiCPhgu2tlhUd9NIweeo8CclW3ML7jJ/e9yeRBAB6AxPm981qYBVOl4pJsKA
GUFYb3DKtkpB7G/DQ9/CqcBYxODDAeufI7eTZGJpRF2z8BvVz6FATOeuuCxqfTlD
xkw9+smVoXnfKkt2iiuSUIxL7LsSccxyGFhsdD8v6S+f4AZCPgvgoGWMcAA4uOAR
0dJ6bCU0qWKy5S1lUvTz2FvjZpKBYMeynPA4vxdtNOz73Kes1IS1DTEJz4kqVJlb
v3qdiISuqxrbCQ8hKxroAErFuQTPoAxrIp3jVD7xqtmxbRCXUyzzkOoOqDBVPoA7
hcTVzIebi5skFGMF8Dxs4U2a04lZf2IoLwvPxLGswOPHrl66Qpii+BAvMo0Vhiyt
oMe8v5wbdIz2z3hB2//kCwNfQJqKhT/Uk3VIEQKbtDLOltE6iI01rHbuFAldGTXx
sIrXMelD9I63irILVTr5fDdItIc6C+cCpXS1AOBokTNqkZo4Hd82a6dNdle4UZyk
w8bYMeHT1IrXU7+ZVwx+qCb+Cj8fkgYQo2QEiy1mLdx9swV1BXWq0i8CP34iSm5Y
BgH68O15NPG/niUsq0YFT8+xbGvDrN/oJ0CR5WqAR4VvXxDcfPe8/cwbBbV1M4zV
Dztoft8kWQ0aREwnrMtwp4/PXvufH4jJgcLJR1I+aQrgugvOeH5fI29HvJ7lTAKo
h55DeBrtlMGDbJ5F+50mIzw330e++iru4yzPAC9hHxWurQvTfKkMwRMr4GMAP2LD
+WPfgO0+ZCId695XyiAF2xr2pvmuNMZU1YDecu20KeH87RBwhsoCjTzGqqqNdyWB
4KX0vzqmuDAxJktpevq3U5MXicbEmTi1NRcZhq7/5Y+RMCMu8JIQH2kjqZ8v+9D7
coaH+6iZZfDqTS/0eRu6upMeB865Og6gvdMk5QSYwlPJZhTNR/0yLS7e9oINwb/X
qdb0Lb5+bUIlxH76K2BMGphY9ucW4YtwR3e0KIlGRWOyYYEZ3doBAVklJhjhALVg
utxct6HTlrFHBRVnug0KFCs2wUK3oZsXo8D1AgjuK2tqrqLzoVQ5fgs0MeE9c8id
3yIppDICjAj/9XrY87maiXGmcgfZMWhiArR/fCDdj/RAWSzcL1zc6VDrTmzNOWEo
HxtWlrOkACpueKsXlxeyqV6Rm2QUEJdPtm/ovGDPWbKKqmIfXdmeqlXaPZt6ZcSH
uxMPeeol3tCQdKIqrvhvOAMqRiH54cW7pehfo9dtw1NXDQrDNUEg1ZMQko/+OZjL
l8e3XG7ffcjTp+e95c5YxigCEo/j7oeNQKWT9gaJcy6gqpv4uyyzy/IkR5S8q7EE
eKOj2ou1O6L2jtEon5qNFftUitsjL6N2ReehD8TcCEnxwpaBvIRnO2F1wc7I+IhC
Kxg7+lKD97iK6HOvprfNdQqe3CeOTqScJertmCgUg2oNLxFMHzpso6zMvCiI2VCT
mvRIAY6DsDWvr8hsEUyoGg0uRHbIFVrY1WkMKe/pMUZu7Q7W7hW/BXo0bLChbFVd
ScVrnG5feDAv2+s6qLsV0L01HroUFFUT89Fc6yeeuHJkeLKKYCrczZ5oreK7i33E
Ljgji2foLyhVVMizCn1pGwnColz/3gSfckoE2SXCsOLFNdLtobvzpJnOTUfcQ33l
/EAlGpR5GQkIQpomZwnn5FLErixdn5AFMX3lNZHp7P91S1uBEe8EFfm3eesDF7hV
Xu6RkvtnbEbOdPghfUUVDMbHOwEZ5lh/FfTMf/gJvpDwG35lhbft0E4z81584a6b
7bdK2yanMKYHgYOyORvcjgOlMKsdNB9KG/orPG4UdELrI08ibSj/BylBTRWjTcN3
iKVikrXkNnXtNMYezNWXqgPy3lQa5du7u9b0QLNFPZ2v6dhgYPgr3rFNwjNmlZYK
sP/JBsUeKQmod/9pdhZgBr2ErIMPljTbTPpNQqUNK3HagfhgaXg6RTgDNkNmcuX4
Wd4IxGv8IrpmVMZkmEtFdcrfSaEnPVo77i0Nr4XqUvMMdHlnSqj2DazCLfS3NSry
XyCxIYkUrsKJsfiGRP6t5AxjDiFbOjZ6rhCXGfQSwq2QIVOHX3jrfTzWCE8vDEmM
8kNhmiKUAkhxug5xoaz6OBCdRwkFGkrw2ylPY12FutOpNzwJS6zHE8ZLzZFNbxhs
DP25v9hKwWVnTlCYZW1VsHePKiavSTLCXXUEHcQmZuM/HlODPsj5Xh9zFtq8F4RF
Yc0IztDejubzR2XSvTIsebczKyRFC2+C7+KuzlInhDxF3nB96NhB0HimKjYv0sYm
YJlO62wsyZRfV4GdAaXvy7IqwtP9BCxhD7OFQtYL+ESfoByO80wVL2HYkj0Tf3bW
p/B6nukVD7ohP0qCHOXx6Sa89ghBZ7gWkYXc1G3y6F2sBUItF1HOcG15rUlecT4q
IhIRGxa8g43gcsXYSCZIHg7rJKVv2XeTBNiLoKKt2rGOJC5LzyJL5Uvu3JuOpDEe
asFwBeZBVn/5xO+TkUKYZLHgyk7103n5ZH91Cbzq3hCrsUtkmJAwp0ryr1JWu4YT
vg7eig14x5ZcT6Ki1jOPoiZzyC9C3YkB9OyYjzK8kI2a4E4CEoCYWLddVzNVVPq2
mDr1UZe0e/PiPuYnNCkce4CaM2bLNnKLJdE5eM1b0g35DyAwrKhZIBydJKZBd2Bj
uj+IkemlMeOqKM0TS9+deBBoFJEJypvuqRe9UkTN8Wtkd/cW3Gix9noZvYI8J/ee
9v9+G7+e+MKrpgVAvCeE4poqsbLNNKVu1DWXNvdpHJCo1PlsUiURBnWfHFSsna6C
wpnEhJu+pNp/BX1l+vKSwHyDdZokSNGPZUJy4I7rwM3qh/gkBi6UifuNYYhu/Buu
26j3JO3ntj79jUaJJrT/uRWsaiyBCKdLWNEuarJ8KJBCxW363mvXrdAxE/raHEKE
+KYIZHa/tNSphqs6A0SitYzFnzFIDONDFHj4JvZaDefIEPF5IlVDVTY+nVXOVFWM
yMKpMVm809Dp2SjjIL3/smkUZ2k1qfvB8SOf3A/qFpOMy+vKSD9IZUiKQafLdg3i
7seZbqoWPEy7GC+I6rstJ+wa1k70D4A2GNzYL/0Q17DF25nc5BUy0pNRZEzfJwLg
V5CGvYojxqbNpFI3k6M6aowQlD1Oam+7Z8ateVF5ZrnZPlUwLQyK6a9sR514zpHT
v1ZCRRJt2ovjqJfEWTV5iPU4JRU+hO9ZhSeAym2OyNCGwFN8vLfT0TH3rv/6jMgJ
Tsfr1gH6NyhZcFKihgFjfE8g4d2GKXZPEL8m6V4SYtZ4sWMXzpQzb/Y9Fw+ABWM4
0pGyWHYtj0IQqsei8UlsexnH8wTmQq87iHxbTPpz0WrA+bu5is/SXmve40ze8vzp
+6wj14ZFkJlgQcie4cy/IvLBSg9+b4X8Q320tFcGtNZmhyaqufcw6T3ClejdPIfk
3a63Wws8ZgqJpkst04Mdpe2SMAWCTeL4NdQUSKtgsf8xVgCUtjfjuNOCSTrLZurI
df5a/Z6lksPA2jjml5qoltm93P7InRtKU8D7k3gP95aSXHBpXs34AYRoRD/G7BJN
g2PSlbxbcQ8/XIt/HPLVFkzp90xjhz107yvVqJIoagn5XjTNFGtm+wvMr5ozdioY
sl39RBK7rLkbKWG8EnbNgYSePEMmr01C89cXyKC+/SKWqPaixRXIEes+QtM6bQCc
JakywkYTL9dbbdo3wBadYLs4FlxbghmbfPiIIhzu4RaNGV5VM+i8qPw1Eupppsl1
qDsAyEhfWAeh3kqu1FpfXkvL9N5AqptJPSDaX8Q2PVtUs6tXb2JXXh5iCJBxC24a
NUG4xJz4k0L3GB8dasf/jufc/RGF5wWjTws7N2lEGvYp3Rrxt16jgmzd8jarR5vk
cfeM0mkodhj+d/rvi1yPUaMIH0Vh1CXLYy1fTqX2jS9ctME2l1iJrmnSZpxKFWDU
g+OwWUHYbRCdtQjKAuWYP4LWQujIKYE4yrySQd/lIaWyL0fgO0e9QsnP6ks32/H+
+TZwlngT7yd9ALqbpD/VnZ1YfCoassBeAwXzUI2C3G9a3DSH+ncbEw1s6InTBPA3
PQpl2Q34m8mnd3wPUujFh9hIDVrcSZdlxXKnq1nf6HDKAw/KYzWaZUqDuaqtMycv
CMCJDKyMZq8dzlxTawZsmalB/Mr1psG91tCTmSA7MeRTSvVkeCbKXk9wZ1qCvprV
L72pLKBuLiCmBRsbM43tpzTGynjaqJ5UR3QEVTKoNO1N/dOk9DqdH85faTOopv7A
vjrW2YHk8D1bM8fPUnjPJCD7TUc3mBlxEwMY07Qda+XKg4OkMvxS4tI37Wj53S3+
yDpJA9OERRnCptpxX5pqA9E1EeMgAlZoXJ66GS+q3haK9fDcV929SxTSZ8mKjSaV
0bd6JXJoIIQChtZcuxoIAWYKvyiegCDjU6CSj3nHkY9PT5GF1A9NAUYYNJ8BkV7S
gLQaopIJWEus999PVAf5Ic9kZ4NMN2yLXgTiTjTt3hrUgHUUj/57TcYJWjoOtSXL
WJW9sjagnI7EGsWBaRPzS5dXkY/p2xDx5jjw0wUVqFBzqMnMcHpOxI71yb2FChnd
AE/0BvefHrGSxvw8e0/5lIC8tnPvqwCtuhuFQ+o+nicQ1wQlqYpdLEXCRYO98RGc
WtiCB4Tr5vI7BXuREhXf0Q73cmnxPUSJkmobxeVBVHSnHSg84zl7XIUNX29JcKWE
Plz3tffaNoLgnZZvD+qTa7b9VV6G+guDSk4jSUDwpP8CV9jI3OoQYXGzxXGn9JW8
d5kYFLyLdc2bZrm8+CoPyIrCdzAn/ZXt0Qb7CJY3Dm5ewUxttanQrItr8MKVWxMY
Umcmc8+4i2ixhzCw6kMceKSG4Vh+kRswSyyOK4Qht/+qA2ZYpxtp2HKSyNVjMeNs
wfvAz6QmFAS5Nhflnt/C8A3r1nTCXZqWN99VMi0Qm+o2NpT0NX5GsjA9Kotq+Ii7
PfD1znXcFJrxFGUJm8Uye3j4STOCYFkLfxuc5kQIw6MDbHYP1rR8Z8s8Pgd8Po65
bJkcATpxuN4ZsN0s2rs6fsSIIYoaCDeyDnt3/+TZGG+cW9wY7BmBTod/0sjPYOjZ
Eu3tOofb+Hoi5V0TRqceUZBeYVRdiDtmq1biVhr/LnRmbWf2cSPdGF23V0uuuwN7
jtwYh+Uf1k8SliIsSi3DNjp1ut3CxRUkZZW69XPnNnfbHPXcv2KrXxc9Q7BUazhJ
W/hpvx04hgx72FUjaw9loYZSsMazsJ7/gJ706KMPdlXMAVse7tBwSAymBaou+mTu
knTdDZn0GOJMPMfaUCasSdO5t2Q70ave+WORqKKDvCdfKSn3BXsVuoARrGjHjuFS
tzpXMvLF2j8aXHZqM4bAmjuR3DeckbdzIdGdqQYKJgCaKaSIl78IJvvUUYsF6pJW
DNnkQJV5pTtkMXDuNzjpaQJfK1928+6YptNMf/PBHC5/RdKlEmCIb5qfKQnc8sS1
h+N3lcwxPrR0sGivw7uATuEnRCmxr2mar7CVuyXNjXUf1v3LRRBIbrjWgWN1YmTr
kffOm5Cp1y7O9KjtKCdUTMcI8GgvFeuThZ42R4vbTrp8tpzczRwEWNHL4Mksk0zq
VlmUfy1MNxLi6ngZIBZV1hJk3SAnSULc+WIQzR9VNouI641IpzxBGhGhKBvTGEpy
/VMhA5OGHAk5z9JjXlpq4aqkb8ofTPyecH09feR9IdbRfZWQ7F5hsZlvtzuttifr
XExIURzv4geN5qWEg1lM4aIWJcHznzfkn2+Pgzh6DO/rlly1vIXuoB56TmCXukXb
HCuQk+YL1+fhZVXejsaoG7ol8hLe9wSXBS9E4C1V2gPiOlkJ0LJjsgKWSOjvf52E
gyPft7ss1Lq4GFEYKdpvLUSFwdnHgwsmSXUnrWAo0I7q3EE0BML1ivnR/4ePEHuu
73obgfTYBcXKzRofMKi9Ut2yiaIiPWBchJnG9z13JtIee66kWHF+7LMADWlCrROB
TR1cPE046xgvadXClZbE2Ey4s7izarJfOyTuzffzEBQgTXRNWUjjQi4TsiQAclrA
xyVzlgJtDQRIFYENxgRfqoBUcKVslo0++W1+gqtDVp4XvN8doAwafDDm39y7at6F
yA0nsISY4Wmne5ljhWzYK1h5VMwWaeLHTkItTq2AE2nLfcmzvZYXUrP8QO3K6QHN
uNLufu1Z1wbSEMZSKlWWTfTnWJwOn0MJ8EJk5hdLh3IxD/Mqk4MOTgywObnk80Wl
lEjN2djv/H9NLJ1+bqVrBPouef5xyltFJi7VfmsqBMePCk5iU89suA2jYGdf06No
MbUqP24qi53idyOc2Blo5mhIyVhX19IhBp3T4iDKjUfx+Ybg2EILam1EckYJnvhH
hbqhPRYyIcLVDVQDph1Kwhq6Z8SyzlCkvpMk6Wb18nRfuqvZ98oiPNL+NYAVGaKK
6zyPlQJ/y5RxG+dYyfYdxFKMDMHYTUccGwI1JYIhClvLKeyAEZiLAeQBmezY1pzd
uL29YMkEquvbX9wm7inBdXZ2iABizDVtCj1SzC1Kz+4+iPro3w9L5zrvxmsCCHC7
kfii8o/xHPvKOejJ02EVhRi1kYzbxhnlX7XYIUReeKSGD1gjiVje067RW5Yg15IN
k50nQsE2dQwX5oZ33n5mtt0locO6CmDZzoajlL8ND/zdqzkzVNyWDsYYmSpQwptq
VQ9onDem6TBYbkXSjf2G3dI4CYnfEO4XCPDrgNlVOWgsi91USlaA/rqDEfg2x3X2
zNN7erRBnAAHnHRHLkLoJHHWeNv6x0M5ETYUgflaQrlsfVuWx9e0HSFbY3xw2Lvw
B0m9RUJyvBL3NqiDjQXqu7ERXVtun2+T17k1qYEu+ZJX6zE8AjG9+w4Bo5G7jEI5
n3N3llGhnPRiC925X//MR8nHIZH9oYPkY8hiRExn9MokIoUaRhVkVVAPl+j4cpca
KO5k+/wp0OMN+na6um8TEs82cyH60L4cTQOcwVZGCxvmU2YV6g7JjYx9Hg40FOFF
R0h5ru8b2R3/wSZBsRsdBd3sPcnTcXzCxqokFXIA4LXbbVYGR5IpFHcJCOnCachQ
T3sBTpJZTiYU4VE9KcxnPfB5PDawySleTedMs0Q9MA6Jxml7swUwWP1Hixlu3ugz
XdlUgmfT1ZDmvTkYOTjW3zIxTCXI0nygqDUIX6cNAhtNB9A5vte2eZG197G6Fsfc
KMaDYrd773T/6MoAB4hh7+wyyXInL4rP6Y34M85TiqzZQP3Nw1WGB298rAXaFv/X
xcsP7DpUslIbCXPPxSPvPivqlmZj/aZtceGS5FPlD0PWLitdJqXMG7gdlW1XwBzE
/72juIj3HEaraWfFVSia0oeKiQBpoDV+CKHaQvNtxstwvKAzpYE4R7L6T9svsxrn
Qp22rnY8yWL10a8V4vCQxUq6C7zfwnhrh855jK9LlqSOiZJpJbkpH6+/rGgeGNqo
dM26GNdCQkpeXnRVPXmigK9eTCZTJTBMe1zB9BEt7/ZPksDeNOHwlf9pKG0pOeJG
2CguJuVeaKDJCBjVcYvabGoNou/ASwyii7GE51SSGLbFsXFhnd5mvgO5PrZza2j5
+udZlwoN4y/OZS2+OnGGqCVjJTkgc28e9s0+HElzIyd4kJBmBQgx6KfMgdjsOzeJ
9A1/AjvCKXYbjP1Q0Mvgw+H+ntkRaZpHRMqg+ldifxNnXjwIEh0ZqgIvVqugPRke
gk2vnE5B0Pp41uEjCn0y1W60vsOpL95HXMGm1JmFwsT24Y3STpOGAOS88ZKy6ri4
5wb6b86ZyNdaqQq9QSs4mhS6e8bv+T5iDlIZ4g5+xHO1N33Ddy0fFAQ535RCRiw5
vvWVWGYkaJfGFAu920fmnrkyEXeygnJUHN27FK8rpK+PbgNbZaAPb/VWVaK4nOSt
ZfP2dMTqLES159qUTygy8De4kpIazpzup7KvPTm4VwMXQkYOhZOlvL4G9SkK4jWv
Qmt+U7CeF6MGG1PUdJxXfKjpXYPQRwYJ+yFBzvlYiidqaFcxHCDcWick1X7wzo/g
ZOm1W/B50sD0ehQoC26JlbKZZ+hd4fby1CSH0KynYNlzBWwbUcdS6wsSykmRJUPU
7wTurXCbWod/AfZzTfvwU5iTz2cdndqmN9UQQMK7rdZcS4teGqAlfC12nJflTq8t
9zCt1BH2M+LcGGAuyyn8q28la8+2wL0paHBC8Efh6gsXoAOVJisUtkbWKaH3QnLA
4BLgqw3HHB4usvLRqjX4bMNET3HxbCVI79/52G+Z5h9Q3bz/EWMX4VGeCDmJT0Ic
qHqsndpCD0NE1p7U8LK8hT9pmEtGOzbynNNyG7pEKDyv4MYcDmVaf4mWWXWUjyKU
5ko5vcCHbiCURpHQLGLtBxM2E/4ucdSaydDQ3WTeL1OkdAWiOkakg5Pv2g35SEjG
TsYb7/qV6MMhrgqr2KfE7PaNKh86RDFFe/D0J+eOPOcIM67Ygn/GOiyeLEBmyYGs
vyoLAEZJruMDhcXJT1E2l2jaqgB3RJGJ+b1P3+0qVQPqYUGp3BvFPspTPXiKRl3X
6/Y03XVRjM7t4PsDjpiwAS5tXssfaZbzeTXnizFknD7URFXKa+pBjm21uMdpWidA
djr4AhCj1aNAKRc9B7TmTeCD1APL7ZeCGQdddQrpWrosAjCYv7Igvgrv62KNNyzf
whfVVhdAV8+ENdiyu+W+ivIy2MpLuzfn+MhjjRDfVuIjnSo5vENdVBgcyrnje5gB
lz3XAd4eaLDM1gJtH9F2Q8zmf3pKd7XpjzrNvSboaG7rKGw68geUcmNIBEzFp1Zf
pNlBALMDeSetV4gVkflKkPZ0gpY5bQIcxLNWpd+WdbNbMU2T8LVaK0GDqOZt0XFe
H/ipfzyZgW8K2mi/FntxmT+Eb/0HUf1+dcg1WQCj8EoMT/TKePnQQNzdpXrGXKsp
68G7c20h/m3J+C15uJ1d1QSPAS98EYxiPHdwjoWpkZwsaiWAXAOV1B+9JqPj/CZQ
XLn/rLMdqTrWZX/rIATpMz72u+k2KkfPW+68S5SoOzWZVjVmMDEKNKrNlJdbQCl2
fkonP6uKUuWDv1tRsrnOy6Ezd1yMEm2K3Enx+VLRnHXj/BcrF7+LV+UA14O1QCRH
A2PU/RYUv1lWNa6db1K/Zf6PGQXIFNlh/lNHL7vXm+c//J/sRdWeIxR1v2PZz8LH
MJOs9PybLDxrqJtnrTDUSVfZLyn7epHebyfJI1u93Av2nwTBFXP2oTvzp1TOSyVd
IQsV0KO58heBA+JvXyUWzn7ZILyQhKuYLloNIjyXrD88G9UEIVjJ2ro16CSIuKH1
X62MVRTXBUr7k1cgbJ6xv79hOXW9AdFIAOihEBTdrX5dXMUFXgCSr2xL2CEUE6l5
tOOCBuMnKEFg0LICUnuandYGwPcR0+stZKqYjrTwLBmJZCPuW2EnwWIigGAveqP3
AV3rjn2dC/kG190ZZV0qAyqawNxhANDfIoQ18JdboPLF146vHWBLLowXTG2Ciq9L
SwUfRUo0CPu9hrEgPNQqTBVkb+2gdMLovBjfHQMRS7bJzYl26KOpKq3/iwk9O7sf
eRXgV8lpA6/n7trnQNKX3MkqdQ3KHmFCs/uc5SsIoFJrx+L3Qo1m9jm7wMIqu1lt
seMm0AOBtPa+D6w0h9U2lTrrZt7b7ZvZ1gXQKDEOu5DB/+8O3edstZLqvdwyf9iA
x4oqPwDSpCQKGewlDyqROvzyjzjvA0++4y8LDh+1i6CUK91AgLgsg1yV43nLvzA7
VZjleMS4Ue4hsrYQtBoAFnQUVY6uIdzzpSwX32tvZDRAQ2jdPYaWCaQTLShxu8Bn
dIp27+IgvFdffNvE8kiix3efIClCd82LU0t04fWzm0gkiVX2MEWruUivA4xKwnLi
lT6yK0vxQ5yr7tvP4hFJ9kj/ZugctUWfOgYQOw1N8Mpjohomx4g0fPk3uzCgaaHV
mXpL/rf2NOE6wpdA3H72crsAoKibUTIMN3LCe3lZ8pdemL+9qAJQUjBpS4k20nH5
mNkw/0145DZ/JsUoj4HIqxzOvbQXbHsN2Gn7Rwv2ETQcc/pgGkLohS8aZkApYiXA
1eWVic2KGpdN+v2oLLW0IpySLYZvTl3TDbZM4gUXPp6b5UJDZgkEbFKAgGwObqMM
ayZ57ltAtgprA7BqOvwot4/J0vdV6ibg979luWqQEtowaY7ksIxyPPRFgiY9rI6h
u23I7au+HdCwVJGd8fo6NyvO16QCFJzaQbqoWC2QaeQNrOZYbE/gYd4EJ8LYVgZX
8NnqhxUIdTbIfh8ZAwpR/sGA5aiQD7wQd3XzZyXC1XaxtosINV19DQEL1fWlW2ym
r7NEJIgZUHXdBd/yULfplmThqLmmATM0wL9Hsf7epladbAYneouVzQaT6vhjLJFS
rNAUSuzZ9UyvH/JTAuIN9QTvbL0KhMqhsq0AT/NkhhLjkjN8Fv1uZFIeCajlChuF
rakvn+TyeCwQzaD5/m9m+ADjp0TBrrJmq+mHoHa15Lgh1JFCJ8pOz9iMjlRH1X01
mzoe6KwCBDOPr/j1I6tFsQpYj/M33SYHIN1lc9VBFyW5sLHvzPHQ14fHcpaSMasP
12cT3PrNhQTSFU511kTEvV9dm9o9SH/lfJpyR/utVNw3EghonVBSG79ci6s5qIXT
YlJsZJhaGQvTVcHLgT+Iu+v7YIH+4rCFKbmkvJd9dQ2yk6OunvM7TZqWhVQM1Q7y
W/Ug3FCwcnrftx8MQ823wqc+862YDlMiliYYacsKyCMYYwvOhucNN0qE7kgmklOn
utmTMbaPdsMOv1/vijZwVovQgEf+YX3eShJxU2wgGPKyXz8Qs4/EGcMD4pxyHA1z
7MQ+cYugC+bao1HTgi6jXmVAtEg9r3rSUFZCoyfs0R6cUceEP897YrQfzEDRD62t
G4nC4ltu2vvIe8Bden6bTj+xbpghftFypadEsBiaVF+m95NuMKrSGdxGyfw3xTvk
jpLwmGIu4MjO0gjZ7iChucugkLz0x00S27bT4F4CMep0hFhU+yDBPy1uBIfGr2wd
HxJCk55m0FZ9x2g1sf2wJ5oiRhNSrMzscxP5dL+91AZjH88VsV6gifmIKjUZw2Ss
dmK9H3l+Sti9kONXdHJ5mKxZ+lM/qUof4hnxlxcrDJrlxZ+bcJ4t4zJcOEJz0PVe
vKHx9fLKSj6K1zYbPcp2dk3ckG+rTxjvcESz6VlFyO5DDgUkf/cBVpMKvO+IHbzA
BbLDrSiTdf1ARbwlkcRCdTmwfSApRSbKPCTwTEs9zBA81BeuNMcknH0OO609xaxA
3UMiKur7tB4CVsSgx/qCoqn4JSqUu33yzOpMrH3JKgRjnVd4amZWgkqSd3hC8K/B
c1LsImycLMmDq0zCSjPOr7zZxQhXLb/SYEi4bFyOdBRhj+A8GMYJxFsGI0ECEYeX
lNHK6tI+sYoe/CyJRpCEeSHJZICBxAoVIB8aA5kmHzP7pUgrsRoiFXY6tGRd4S+l
RVTA6K/fmX7jnHu3HiVzvcTVZDbd2XzoYwCruMjUwa3tn1Exrwl+vkLA793IUzVe
hCHPw818jefZCZRMiVVYSf0I3fAP4HROkP6xCm5/Uwd78s1Fc13/YEmKNsGn/rH2
ybY8PJ6RTMG9IJNwRXoWGYpjjcFSZv4CHn2QEruTlSss1sNcs3mRYx9C9KI2wtHh
ghheI2Ioja1jloP8eK5l45Lz8C1fJZwg2gImi67jPPVn8CwlApCJLc/5LSPfCU8x
bLW0SrEi1jG0p/ygGHH4M1nuxV3I3FB3p4yasXxRxVg7/Nm+yI9tZXlErGiYXju5
LVOgnvgecAlm3xYoaMOiMSjUiep2BUsyoh1vn558ukKTFLjMFyAJhSm0X1CuVTyE
kPSxVTBJNsHTl61T13F3EsKyrejCAXQ1RGJxyJQygFX0oaufVFBcVlvZRsFeqgzx
8KpryTd7NJfJXSqKSBJk70hMooi7IC6j++ZxtzCAJam500lJ3ic6k4k/3nN0Z2gb
La5w5ruyyy5fKLUndHkF+mYkeoahgQMAyEAgD/s9f2nXRBVpoySQ+y2BOayz1coL
1h9K2BsYGm0hbm34Fbi8YIl9P0k1qeGzU489zvLI0JvVrq+nS6WK5DzBGDcEkAe8
SCW9jE2FnVO+WLTmaPKv9goc4IpDEy1IrBmfe7yoNdGoC3SHDZzQ0jnrEtQfDDyS
zBizCtWhieV0IDGRDk8DrHxo2TPqnLHq6voXgbrVGt3aBen0aOHfBQb46PqjOTnV
trvYyzbNEDDJAtbm3qlFZDnWqvSAVFodLXQM//LYuAcAJYl/4phOfDDkCWutUxuG
TxXY9leLk3mp/BKlXYIPHEMLaIdO+VZ1sV+K33xP2+pKH24wbG+zfuqsareInEj6
j4PgO3LiLh3TP4rVZh1K3a4VkMJHEmj9T+dBuoxlkg+ZJs+shGiuEsv6LlLnoNln
CJoHf8ZqLEEd/wuNPLP69TTDN6Nz8XfY28bDMmMzj57gAqSJQvAIzJVbvmX19pbb
9yaDemWskdFTBecDFPKOuD7pIGbmSjSDuE5gtLqnGFyNTC4Y9kROzVkTfvBqsHMa
+y/EIIZqDCj39PJuV41x+/OlcmA0/qjtcawCCSMnzc0PcjXtKhbdNkXOvtNaASfY
LnYTBG64zmK9+U6Wug4WpwTLa0vSFibz/CYYLitQpprG/SxPuFXpYuzuqyRFLc57
lS1a+WNH2lsCsn0vR5Xz8jXzjyuWgMdWgw/Jvjoh81Etdx/NB2+XgztHuQY2hUMh
SUUKyLI1ZwCHX2fo2VZqCQveuTUTU1NXO8rgRcWdhB0wn7vP0FO5yundoKdh4Xym
2W13Hizddi7tX0wQ2yO56sdYzLBVed+bOsy/KjkrQMLye/ZqY+FxYPleV3wbF1/z
echG6Xh3jub/63UgUsGWTq+xOLHvR859u9Fj+EoYZUNMWsqWkCDjm24/P1H7Wenb
lzMHkDKJr7FOBV6+eAdPJobChjIKS0BPax51N2ba1IxH2rxaKoaTW8HwytXHgUVm
8t8dA3kbJjCrDTvKYl/WXDGT5g8eYlN91BKRRyyY8p31i9i8s0hAF4sc9HS/JnbO
cFZBm354LeovsjhQZnI/QVvM7cDPjyd3nNW6xZd44pccM4cwZaMFHVSjCrW6dh3K
/s2HqT2Z0/qk5f4n2xZqHi9sokCci6LgyVT2+dkWvdP5HkkafFJ3JdIESXDYe950
AtD3t9USvf13u4x92S9XVhjVRjB5m4S+65FPr+ViHDM/3+P3skzehI47/5NdACbR
6QvXNEpWO0Kkbir9H783c55dTGzlD5xPX73X8kzEhIZUdsVHXkCtKLMpP72vN/6b
nmuILBupX/tf3MKI+dv7sIIHcX7RjCBv1IcGwEkeiuCTgeckzERMGaT3j01ER4ri
0ySGRLZcEopp969LbZBSvEZzyJWTEUNNWY3C/Ph67ws1zIdJu9thI3fjghIhDz6X
ic5+TywkH6XMC5Wai/cJIZTwTQs8a6COEUWu5xeBLHQupte8Mwv1YbQ32KGh5+a0
2uM45p0N0+kfOQ/FzqsMglBPdGjWr+iWN813XT6TRgrn1A9p1md2zdt6Tax8EQ0D
TTLszd/4hNHKUsqmsYKb16pFPK4QF9652K5DAubt+YBFCCp7YozZx0iNyIT3eHfp
wfHqy/7UiJ7nC6MgX4+8ffSd4xkQTLUjGmMh6igLGQopvi5bYp1kAASGqngU1aKL
YjxJr4sHtTtQKDOgn+Ak2nwdfLJ5ElrRKhtzWcSTcLvWJLDCCSyn+HoMckYpFlZn
AP59W1nVUwJMYXbliqLWeHXQ9Jf/zdy6Iglrj1NYpo8U6i17rHLaWLJLCBMvohgn
1Q1DsWfCIWEdsKR9diKapfS1UMXnbrw/rUBkgl6csSRzy6+Umc9sVpOPGQHGQZ6e
SRb/wo+zVVqgSPAUOfePmWDEA9ATcI6a+xSDdEm5UiQXNkVcNg2J2DvGDgnBPhE0
XyPZeZxcGAzvUkHl0BBv5UzeIBB55i+2Iazv75AT8TaO1aRFIDzfRuotk6ooQSaS
lkiRKtLGKXVu1TMCql4s9k0vvz/Yigpy0jukmbNgKJdjc8qGJrK+X2DKs4DETDMH
zPQKQP1fER83zYqwqE5k80cNH2Ajmskv8xbRTELzQ75sdtQ1+K6V3QM+d9MQ6DMx
LDpEdme4/izxBdX/AKyNmk80bJF8limdfgYM5HKLWG9QmdKMB/W9s5CLdTWJexTm
Ba5jCZtFyluPJAj6d9NcETs7lTlCL9rbQ9TZPCGSY+7lrNNdpYfUaBoCLDI5mHOy
Sd9/2cTprnpEf/Sc/rLYJp+gZ5t3vHitXI3qyzYoULW6QwTCXUA7fQtNVY05LU/7
bnCdWqXUvZQP2b/4QE38vHbQxemcSqULcndj/rtlHSBrY7i7Tv27SkXOge9y42SF
FZHuuTkLyaWB7znTPbyVxIJtRf3JwvrWWVI4d+Y1GgOwJfY0BRF8x9bYuuJf1oRq
0PmL1mTDGDIwH8BBG+Xw9KX5mwYoBySdnP8go6r2mj/6aJG8AldSKLcpuMe8c3Z7
p4c3Tn4fgquMUunCAuIYTby2Bk8BCVGu+4K9wQKjnE/YXFV19lCABwbpFxyczSMx
CiyPUpDn6u42uaio8MKRtf2+U9v76YXBW72B3sR0/jSllOKYqfBDhVqoIvR0TnQB
b9ucSlLP/p1sRR7ckJVRUOMEf8CWtU39gEUSHhrXlGE+r4L9ODdWM6aSVcKP7PHS
G95oyUH8a3D2fcnxn9op8VWFwDzBjl93TGNrUAz4aZaeABE6+4sH7CNOiL1PtKon
/vFQt5fQuDBxfgyxCRfrz6zI884TWs332euA6UxEA2BMDxMpErOtXi++6+xvEr9J
9JN++3Oj3JuPtJc1VDA61umC9TUZnDJZdM6+2sH+9cspY3xbL8EwAziIkXC0sFwg
QXTnWyUnqmguQNvxmld5tPV4tulr8/JL4cfb6Ay9qpSPyaPbRdzbsaEb2dIyOzBD
e4jCszG/EM24ESbQT5bb5/FeMxRjZT5KZCG0ox0knn5ZZHyk748sreWolaxeNKWA
Hy3cT97AcjGt31GsyVzX3x5y3XpRj1QtfU9MDsVR8YdWd8RMXYzN79KXNc/ngJWG
j23cAdKXGRpAIy5bAv2Ds5maK/PER5Cmne8wOXiLv+8BGylCJw2Vkn1cOVuVaUHL
Ev1G5sowYO9VWnJrqv6+mzGH1fJcpqTX5u6u95QtDh4s/ibI4fNSkAu3hLEni9xp
5yswKWKyMaBR08vauuZuZjtl76mRQ/vZq+LkUL1azimvxLjj5NRe29TKgKzlZVmz
wlOkFXcepTBu8vXCG+m6kN7Bt5aaaVF4B1/AON1Tb/ttC0iRS0JhDHuSCgzVKHRT
UiUndMOOExTJcrFE9lUkAL1ucbx2t5YEWZHcirDaAwoU82+mgA2CxTUSfj2IaZDF
PTEyuy7jsNll2tRLI4VVTtTnO9IbWfqZHsCrSjmdScEap6N/bUveXDCQRUlkZtMC
5OB6TzJ65Mtbq/m1cr4mzRp+iBH6hta8T44XHodi+3qRQtniiHm3nKwPNDB6xIOB
FcDNbst4BdqM6nJt/npEY5zvhrI9YLvmWZm31zkBQ+yOPXmhRzysqKPwnfN7HdyP
ww+7Ug7OqdsRQZfKltvq0s+70IwzsxAzSb9IkAuXh4eA08puYkVMZtybxx3aocpx
D122GBBxvTrvemK0mCOIY31ymxMU4ph2yU/96LTMmP1IuxclL4j/Li1fiFy+Ehjp
VMNF3CmcLgzEPWG0rrixPvdEKdBW1rNA8l31+nvvOa5Htf7avUP0GdyMNZL3isAc
XfwLAwtn7LGsWXLb0u+yseDSLmMwStRMZC7Pwj3lKUWir2AjCB6MuVXcGSNvosSQ
dgjsT2F5t4tZDdDdht+1e15xkkSq7YvpLZe33SsMz9tEnq04B2UWU6yJoebMZ2tZ
cjq6Od9gmxHs3zT9Id4aneRmRt/XTYRs4Lf7u4ldoANXPkaDhMKn/mYgZL1adJzT
h5oFdUViQcUDhOZ1Zv5sWJuFbbsx+v6K/l/x5EZx3FIfrbTL0mC85XxHWYevUQnL
qpi8VlGwRuiPYZeFhH5riHFAxDPDTMEkZNHCtFHcK/5aSI6Q4W+myzGi1DpHZ/JL
qJj5QOKeOjbbmRBB2KIqW8kpKDRFtVEbv38+iNEUoYk32sUXybKroYsdV24CmUw/
PZqvvqV7A0Cn1X0BsWYVi5h8169vtZKHda6V7obR3p/0D2TqOFoERN5zzSRhjMlh
Hq/v2Q/fiuD2tSJYeP9sbxnT6fUoZKIQJd8LjK7buOAvajmCUM46mOU3lDPa2JpT
76GFTXGYRQ1NJdQTO+1KXSyjUAdri3C9TXu5nP96fcPrCKyH2txpuLDkOmqVa4Yj
LNrLn7R0D2z6FRYU/h9FWc7J25UnlMx9vf/h8KUhVvaBID7D+9zzXL67j9VL7IZM
d9Zo4pHdtlbVGPXTj1zOfRgyaSeuwN3SufZXtgad75wzi5Wop5uJpUJ6nxThy2J2
UDuAmSf2jCHLrcGxUmIGN2GFuYYD9DOLiJNC+YQ50aP6YJZaNF1AqyT+I8+SfB3P
yIV9N19akmAu9yPu759Itj+eDAFfjHao0iacoTYjq/uHJtmyE4M168jWUMy2r2Z3
ivdzMwya0W6unL+wPDBoauNmkfPg/Md74PDt2498HhBF5sbn1h+bnWUknlndp+Hd
UwUYM9KZirw28LQCuGsxKOqolNHVmc8ce5WhYM/DdHQ+QxAJ02VWMxqtM+QjpqM2
wtFJ/m00S+w0G5OiKGHWARWmQhSiCdBAsNzXVvoMNjDi0WF7zpQfP5uJcHvHTNL8
1Nyds5mmQBaH3oE8gL0cE85rVVQaJayWMefdrkk3E2NTiR2SLJ2JklAtrbBAGmc9
qvxVgytjWZszzObTK5U3w+ArKv1u+cst64P5dez2J0afgOTbvJHW7EnWt1sTzOzZ
N3utZbkUryASgCdCdXU8ER8jxYdEvNA3jCU4obAGfr8TSsHeg/Cq589+LoMW+DI0
MqmSAhl4pSyn1GHzbfmYtNlnzBydv2UNm6/Z7h8WtTA2+Mce3CWPVfN5//IHYzja
SIrI+9ZsFdoPvVHmPRM9FDImNFOV+vw5smHqHqLqCeDyL8VkOK90kBT+sNvXV9Cx
2srOy5njJ8Rj+eLIYO2UbUQcXjPO8SDYwP+nEotXcuyBQ3RDxNu4ureblkm3/cBI
N52wUXKbsG5x1TpfSn51gXiyy0f+fn7bLBb6y2uLIsV2fmh5sBBqxNJXZwrr9Iuf
ih/V+VgYQSAiMg3EVL4oPX7/wWTmLCvEwL6x1WlfMJFlC4xf+470PxUSAdGYJa6Y
NX2og+3AjKRQGDXAdOMsb1BONFOl6W3zKyo+/Hb/oBOEJbWMSKQySbcWXE0DybVt
+AGupz2Dkyuo74iu8DogKT5ydH/qcQWWNDPAaed4Dfylhs74Lf87ufaWrRhjLttd
rgkY5c47EsF2otr82lWg/Zv48MBxMjBYWwofZbEmTy2sGrz4GjVD4m/tJve1jPjS
F4BsAWauKfq1EFlwBo1U7+ejcPUlHaPhvxibXxc5ZRZBNp3zB8Q0aHFxstpdspvh
qOhRYvywqEW++94KPabDND6X+JXdpVAIu/JEYhkH6riaGaJhfYN14hhR5k1qzquB
Y8rkwvR45BjBgAWChVpuoNhid+cPVJTjaA3BkmG0jAqZlCM07gTe87wLfLiXS546
n9goYIYkhHeh3h7EsCrefDoW3Rd+S874lzXzw/29odoyjkvqjhLfzgzSpeByjJL+
ebpVQzmgsJwBscfDeRoIKUKV9eVr/ZFtDTi+DNsU11RIhr4XNuc5DOA/3QjR/5XM
B/VbLsj65W/mupdb5NFPpKVrmisrOBrOYExnW+7WZlK0wXiXIpuZScsMzDGoILpy
p7ASggMlgXoyT1XO1TOJJM85/XvSizEcOv7XCTAdUDAT9k1fJDCOBrlsTa+ks+D3
QIKIdhr1aLlkubuHURAvxWedKTYSNFyjct2vMRFsjLm4oMnmPsZz4eAq/kzWRpHw
4Z3SrLCm2bqzLy64GEA58GB0q6YXqBqjjutuCwWZz6iARHtKxCustJg7D439JwIP
E2NBIZ3gFsuR3icxsgjBI274A9h9VYZN1nNSKPKl5XT8Iyz/V3ASb+hr2o7ad1Hb
d/uIrreXLw8hLdnZqciRZKQrj95293HZytWq/fqUWnnZSFJ6CBsBMNjVQmPE6qaw
zEwBGexGXUIzcVwqzn02LDrJQH4k2/bXxfAtfc4TbixJ5djehaGcWgxjGbD1qzN2
AeqPEszIQk1oQqrLlwQ9c0HkaRDOBzkgElZZXCysyJebXi+xQjYAIPXEBSmBFLYG
3YMCsXqazLqvA7XQN2CAwTVl80qIOek7eiQDch6V0nkQHOu6YJ4f9nOnZAxuEQWP
VgW3Ebwht468YLcRvVUCEtsB+UyI74FVnKOh5iDMEZkEK4S/YzO1SB48pNHLHNB7
MAb1Z7SnXE4e9aAhkVDs57CZdyOV6wjhYmWJnIjcV6x2HjsUNH6h9LghgBi09HUY
XKc98NcfOeKJy9osdRrGAmph6OytjaJsTi5Oh9jJBVimboNWyNpO8zsWOSiaNDj5
Ve+Q4CmFU2VIzVY2Au7+qFzKoeYPZZ0xv07yUvEHxBYm9E6Nsjw7ZsKD+kuNwECg
/gwmJ/WxJwKBgmQ8C8JW/0eNDJiY7YWbICkjpIBLbTFsv2PB5cXyrWeHxN+i17UZ
gljNOEwkAINIBWAWhfsDZJfO9KktvndFKY9E9R3guONLME1QKXWOBALFxfeQywmD
tT2c6zfdjswmB7WswWqMC+hMXZ8oxU5/NOCgY2gN5+da1i+LM9mskdrpL2oIQdbx
F63IAsYvIxa2g32PCbXl2foIy2HO3yjKsp1V+U1N19ddQn/U36TJby212eQWeJTO
hODYj0BYxCz/ni83XBbyW58QnkV2D4Ux6QRfSe6YG13d12aGKHpiumqhNSiWX7rl
/q9OsgrA+XaMbnJ5A+21gxwCUiL8pFiXINSpvKzPfg/5RsuIHXnNRmQda6isqkfr
L0YQjIzww4LnByl30fy9X7sUQXzqlrnN+yl3NY3InwXHDWaVc6HmBdXX6TY8M9T0
2S5lyDBcnzKakngO8YWirDe8Qe+riNT5hg8nNsii8OvPL2Xy2CmU+puqP8qj+d/D
YUf9ttXpsIiytZh10iS4NOLsoFx3aPmPcO/sAzPKI8qXK8z51gYN4Cqx/58oS/ka
1WMCv3FnOht4aqLYu9qBCcHuiAmncGOKrdLazJG/tNTbQqpW4FiwRY7gp5zGUccD
uZe/r/dA8kJVQqtDaT7ksHhoByvDs84ZV+kXiaNtv1RLQjTb4vJ5zoeHwFWl2hBw
fNUyMNdMtsyksS+dVAw84WLehqOMstuowfJmAjyhQn5dBAGPr2+p+W6+e/j2tErk
FVeb75W4uRShy/DnCWmaekaJcudcUO42b5bZt22kg23JH/z4B98QoyTf25oWqyfd
RjI2PafJ/R57oAzKlrQePlkrJMJIDddmLmgellzBct3fJbD3+040tmf5N0j+IriP
cKzlmZzT2oWFLy4KTYMOPa4QGrLrEb6Pcc1J5ngVERS/O2iO1IvY827ZRBPorXzt
KaTHrDiqOziEh3aFMqXO4pBDIGjVfoEjy/mmZo42W05doRX0c7j5TVeO9bP6nKGe
WmCpdMG6MYZ3yHcwdSHaBKCckl29SkNV+CaGmpbOFSUPltjx0bmo6Qob3qVue/5H
yGKE/47iIxcSXZzQ0s+E+I6BvNbLTQifDqcYYo3eA8PEZEKLYQ6nOj3Lr0ApBl+K
plqvcvG8IYk4rTBIee0cVf+Lszx09O2c39KPgOD2U2VgYeR0e9i0ocUtfKBD8gs9
DevKnmFfzEwokONNcl7Szo31215qWDaWdvCR9zaiAri6wH7x/r5zNpU4PYE2zGeF
l/RihZSRkBNTASr4aH6svXZdhiz1kq8wN+JIum5V1vwYLbz1OIj2xi9W23dh9wzZ
oNLqY1TQHNLn7n4cUu6jB2NIbdia6zesBKsfuiTK4AFQ1X1jghAp2FQdRfQ0zRJX
wqFRezGISCfrTa2hflrmtdiIblGbY6NPDY5xkNLolZnJjO8tP+YO45csmx7Mv8zy
V0J2Jie4blXnmRQ+k8A3fUzFsVMhRswXn1vlynO+qFuFpZiWx6WhLL82LxWzndhy
0+JZGhjMWA2aWJOi926WPy1eUeD5eP+XLOQwjAbYBQChLDB/DmQKJxIKf9FdIB/j
0xWncgqpL5o2tRiJ8uIvKIGW5HlEtUkOL9OsO12enugLyNcalxP7xJA/0Iy+CPI2
iftaC3YNbm4ZbuG1SvfGh8f/CfxAbd3BAM5IyrmzWUKbLeMHbAgKmsJteWQ0eplJ
aF4N2zdIrUPPtc7y2+vJxXgmOVoo0zhSkx5gR3wH0IEGEcOmc0I9LKZ4erjIGcIp
R88UklL7liVrT6uQgFYvSH8dFg2KzFceayGnyQrnqGrBQygfmSMxLntpX8vgzQaX
eKQYAQJQJj9jFGjjK4myFW7khR29+aza7KI+JLDwCD4e4q4kw8vIMd4aOyXu5oHN
QRSlY5NG1f++62s6SCAcoO8bhhD3h/P/HGaCIDDWfy6QiZ9My9jPAdUIzVS1RRD5
+103fFgDjWymNEGSDlJjLnlNVS/lqapGFsvkoN1Gyb7/k09lodv75dsotbKOFZXf
5lmJu2gWGIIMTkx04sEy7IeUmfePWpS+LethDJtNeBT+sUyPI/0n/YVa/MOQaCD1
2+3LK3b8o45Asu/K7FyDtBw/ADHDjKkIHbV4a4ReATjDG3lhPchfzYOKQJwajOvT
trH01ovFks2doGpQv/erXPG4P1EkSxeX6iEO1FS/TDdxbvJ/iBXXx63FHrG+zGq0
BLuz4Cgd7C368B2NAROG+1gwwpyaVgG0MmchlviOLFfTfI2p/NtQmrONqX7zSm/S
1IZMH9DLCRfOJKNPBMt3rchM78khNKTfht/Hli2N7ztTvA5QYqGru/7wDDQwqKg5
nJfkl/ycYRgXrY5sfywI63pbuziEM7+enBJPEmy0hGHO1FKqYivzNg39cC8CzOsQ
EyoglR9zWgLWXUOu98mD7ZOvzjLJQgAWfLj3Deg+csCULtay2mOZbZOOF2t51xeH
xlk2DRZMnoMaPdD5hSvzUouXggqOjwU6OwyZaJ7+M+LGJ2SYQuBK+Wsr0tl3fKko
nZ1wMn4HHi0poftwNkNEozIBugVc1KdSKKe717ypkflckA0IR2VwS7M8XuQ0pXRO
W3OIJrds/QWAkZg4sP0g6Rx6RXHJtiSohTXC3guipxd8VzTmBbLxxVuul8eJx2KT
uSXcNgCCeXesYD9Sa4izjFjhmcGcnAo7Fr/X2Uc+SX3YAgfcQvyKiPK+vFBcQGQg
tjHz3ckA6W1peLV2OZCLtHimYRGVVWauhaPeWq1Fay4FA2LfNpCwxiyARiw3RpK7
NAlRmrexl0QsmirI0+k4Ubh1DKElsx/Et2+3HH2ZOeQ/fKxr6rRUv2RHtgo1JLO/
0OwfI5kcXk7rLCJT3x3MvqwOKSV4wQcgtXU3KJJ6eq6OP9tC8Qa7IIpWpjjkXHj+
4U24YBg9Y/ov9/DTXKBE26MHVe+EvLaKKeW/9825+F0wBMHjv8LCmuK9FANty82s
lqsk+06GrOZtcW7tvkNU2L/o/s3POfCnKpAQCGaxjoAxJbQwPTRYgwE+2BS8uJdg
rVS02RbgAP1FoTzsE3NkweKqiB/2y8KqW+OciQEArlTUpZo906ND+jljvH/rOZkU
u9F6RPKskWcrTnd6OGYuAm1vAAseS2ZgvCj2qEa3KMSS4a0x3znfNcyPY2ToKgay
meSkK8OKxmEoz6ZHMNp5ZwlTdshyrKQh0RiZTDN+CJIE9qjAiy0fxMLZQaJ0Elzi
Gp/4NVvxug0iXVEO0m0pP5vM4CB57CYEWWI6tTCgv6Aq0RI8nooZ+LilZXnQ6WpC
lBuIds4ZmeBhL1EdjObE0i25oT4kSrfpeapI7YRi8sRkAWVr348oEkoDaG8fDC7m
FlBkpcgrUSf5cem3szBLjvfkQE4r3gdXuu0Akp0tFoquwaOANJ77BGZD/6nfoq2z
FPJQ5dznNFemZ0H0wTizPrMIwzKDCk/J1iqgiwOoNVuo9fC6H3MjxtDCS0OBuvqy
X9z9yYH04/hxMeP1iDLTr8I6N/QYNU5LsNjNAc7IJvCL5S41I7VCEmiOgKJL83oz
y+P2AWnXvM7v9jlfvSds8ybnicr0e4uyA4g54VErvoxyI1ACo4mE5iMymaWoJa+I
v//Gmpwu2g0v4M1ixHFKzyW0otypwE2iIpii1ZJzURbOxPMHzFq8wlsGdrsIq2QV
jVhUsnRe5v/u/j5BVibNOPkWQx+qH/t9FdXpt3ojU0aATpQ9qhUmwqAfcjq4sWRk
0WNYr1GcjmymB2wGluXw8EPn2cdWbvdnkkdK3zdyIQ2Lgg3DI0cejc9SzWqz+aLh
GeP9pnikj4cKX8/hJbYRftjJPzQo+zwjXPbzqseZ+HfIktbHXzkqoxEuxXufvf+C
yNvvR6/H4jKpvgwxuKua2AqOciU29AH/pWha9C0aMDLA8QeCbLDrWTCxKbxODiw4
5VVDaytQTjiGRlOlZuKYyzMlSmafhK5GFnQdXvswL5msR7T1ffDaVsz3KKmwvY91
1XYUCRQhh2pE+FGVKXjiCLHA6Om9is0FfnK3zv5ju1JrH52BT5AFTry7xxQBwIpI
wFNsBs63So4MPSBR8TiWvzjn7/so5MFZsp7smX8kXiuCf11xB+gLHudBOthywkdb
cx8d4GqcHs8RKW67rDWYPslJPWESeezGGZDxZyzfJ7aAxIPQIAuk1SGOHYWL3UHP
hffuElXvPZGwyh4wwyKVE7ZqpvRDyTBWjNI5bRPSz0x9yUCERY5TV0ddzCKa5St9
5iSyLY7NLsUGn35odgQ5Lx/tFPiGNX0sjkr6/bfS3vsw306ThKLvU3OJ+sCPnzdq
eFNrzi0TnmNWFrYgCvLtYrDp4PcYcMi2586J4vLBzZZiXa5rB/wjuqemx5OHsC1O
gtOvwEoZHC8de2Q1hDd07aj2QlnHEMevr172P5IbVToWQ1OtfHzOX6ENHUssb3pb
fff5gIGbE38iXRfZj22s3c27HAJN2qpkguZp0ba/dGyLPFnwNFbbbLQIf9vTJ0hF
Z2igiM4lx3taVNwPWhBGaUTIYLqn/0xeT7zKPH2iksKvJvbC/vXsHx1nhz/oFI+b
6B5NypiD3plHkPVHPBproT0zF/C/oE6VH0G4XjLUpK8AoqBU95wmN2ddN5nE279s
qJ6eSkDOGB9h3ZsPZ865BHs9mvQd+gOiiq6AieGc1UE6Q9KhwGanMrbe9jsG9ejB
t5xzPh1bypQ4na2F8KjXDXp4AZhRcS4oipGi8gglgcHSOpMTh9F8eULDeerU+f7A
6F++iCd56HvcG7DjLpWii2oDflaYSppS8iONIsSs/xdf34i4au9CDnpGhAEjqL8J
Eu8gtHboO3FjY1l5bO0L2whZTX2MD1KJxHNcSwPL+z1U9h9Lpx/rz1LO7mjxIBDm
qelGj5ujhP4sdvNRzo7iE917qHw7wx2hJorG77J7U5FPRW7fk1Y/FSn4CcL5H66q
EjOBj7UD2GBLbVy3SoHh6FC32yI93axFAB/JyuI1yksUru26PcGjE/G7u+kPE3SC
p4nKY6GVnOlIHBq7+YGSz6hY6D8j1KPSNeU8H5/c9xDMrD+L/UvsefDfgut6nSyz
h9OfE92hVd7/BFLeeY2xxW2kDmcTjtMZjgDd88raANK6hUHGnZyTrJSQqWaPl5M5
E62/zjVU11y5wGGRsAwc0iAz0eo4M3JyFQCu5ycYCsIJZqM4LNVe6piWQIzB+cRH
9NW9H/UjX0V3q41orPQU9aLlSzNYCHewQPsSEPVeGJPt3hJWfg1Uq9J3vCT+cGhc
M0EQ1cxQQQ4/McZjaYNOTaHM+FduHH8AUMWCS1XbZ9Jl/5u7w0RnJKzDpn6ypauz
9pTFFtXkis2jm5vXtPwl/bcpAEF9bH4OhIXLU0Ml5QbegAjXx81dNe9RlW2jPbMU
wC38iMqoMQ6EnFiU3fPu5TxjKiYcxaxcCsF+wiuLs8aPgz9872Qt734CxLegmFhU
Ydx/fqk5P0sq4v62IcJ5dTvq1/vHEOg1y/+oBmdKe0x32vgy8TRlNRnI0TZYG/ME
3azv2p/CKcvnyNF6dlUYgRrTrbP4nw6NxLtfS5PSTJauyUQpF7Pj/ygAgXvUkUrp
+ohqCLxKPyWvgpZ7jwh9LNO1ru7ripJvE6myfrYHmZSMjiKAzU2DapTCRHo56b9L
jFJ0/haoVgfO4PabgP9+X1hhTgg/P/w3a73qTBBOR0TpagJxZnCUPK/uj4Gg86xZ
LE5TWzz3wOAXUB0gFfdbf3aC8lXvdGG+8XBfYjf6t5yAA2p4febk0S0KRhUQUkad
D35btVZEsJvGK35V2CQZVLaZNQ0TiDwLJOxVL4oxG27uDF1lzmIV9TUm9jpDc5/G
qTksTiArW5Axz8IfyLy5x9UNyz1rYU1AnU5Tsq72Kr7t/voab+vajRcaJF0Wl4ny
ybFDGof7Xy+uQfeW6wxJU9xwjWscHpiJZrudRnuCkXYJ+Fr8OkJejRJsj2+HNgy9
e+rcSDe71KNyvlR2GStCnO1K2hFnXonyHwjHuAJrrs0rUGe3trGC6CNjX1Ql1kKt
p7jK02bjqtuT6g1SPMQbufIKoXQgrfsDce5D3KyEUhXlkkFHJLH4Z5rAWtaFi9ji
1Atoz1/vu0oiWovYhsZIv5eGJhEwD1YaW8DdrTIEb/OOIMFfX5GNZWC8Qk/o1lOe
IUqrtO48E+YfrSC8qHqQryhPLdJXGN/Gs1X/WY9S4Zmw0sJjcZZXzj0FbqjXqAFf
YjhAAVObyA3pnouxucy8lNP3eFxNodxIMuuM1HkC/47mQ7/l7ShcJMtFbTBH2zaI
mhbD7/i0UZPTxFEZgwNlg5qHV06CXcRzb3C9Y2UELf8oEFg6cvL4UtvWlXLDeIPB
D3pcQ/G9qlnFEu7/9N/hbd6005TDo/BOusIP3Kzc41pnrCxKGsvMoNNSQ1RqM5da
76aYAYE6D1rZSgzF7ZXxg27fF8iVYxatWWQl+EgTm+TXanSpluIJB1FGpnM7Aiie
HvjnjUXADeA5VUO1ptC5c8YEOlBeBuHdyiNQhiVaXngH6T6sByZDTnO2uksJGgr3
E2jbEmS9giCyKK6qGvcu4ZbOuIkrqDDtBzjzT6LvoynunCR6uWlPE+H21GcNCRNF
c7H4drnSZJlz32AmY9E/wXPxkH/qpLziBlysXfi1BNYUU+KG65ekJiftTKF1lbj2
8Pft0Qo6Hl8oeCYHNh4ZrAioiETJSN9tzwBpOiAg9AGHZ+YAS469sYSeDaELJM0V
LgSAZpRmTe2VUxkGvEwm1F3ynif/fWqEjikH4zc8FBPxwGA+EzsqMa/aGqcUcDul
sPiTpYme5EkDfMuq1ehqieYEEUSLoB5hgVJX4vWX1Rw4z9GuWDOsqYAOtyzF21QF
F6xYMakusuR4wU67wq07EhCg8H6glKYI/SJWuCeU23ReEt2YPoLsVdQszJF/psm/
Tu+RJJrnFn7Z04kaTDXK48XMh2y03hhk6kbyXNTcuXoc557+f76QtWrHgFpp+ixa
MPhh4B8o4tgptr4WXM5SntBA4P6w4qpkz5A8xtKeedFasz17SizGmauQGS8bX+c8
Szp471m7caA0rF9mYkdCWRLPfq4YB+iYxPz9RKPYQpjHhe0tqYIYuM0IVGHQgEd8
fPJw/g7WNgT5/OZ/k+kuRaAPvqFtYDByoDKNbEbjLR1Vi12rv5SFZO2Gljj18kyW
PT6+yRFrDGu9b1LcIUPWG/aTbTHgkZhJ3HWyuVzPQ1Fk4zJJHeuZFVcUFp4IKeDy
0Z4pFErgF89LKS1f5KGVqrsgKxgKUd+wJdXLmOX+KyGMMDgkRcos9ULtOJywMxtF
hDOh8AyTtLs/Loa1VH/TaXWWX/qG/bIb6LaRsHj+x0RmufGB7wZo+gpu3W0hwa5t
n55bUTD2J1UQaCm5Olcas2hIl4AR8XdcJ656WulBHRlzoD48+td3z0ZjobJ7QFcf
XZ+UGrAaKi9KtPPjy21ZZ3jGlMMUCvRuuiD/LiiR8nnlSJSrjWQdVPxf7q/IlFXa
aJ2IrAJLTUMHRKO7zaFE+zwza2dMzqy8C4I8ahGryZkSZe6GJcHV/FR2VGJbEbJx
xUuCqNpUlzbQ7pkKw00ytE5n/D8bifUgo8Vfnfd0ldz3/TBkhesmL/UrdWc1eruX
e6K7tTwnlwe9JkdbrTn1+wU1gjqRaAsvl2Gf6Lgve2mfh4us2c5GE3d87AlxrxS4
8qVRBCx1uoUhUjQ3oY1cK42a8hcSNwoHHjYD54EHYJgo2zU421U/EhZxDILbI4DV
pIXs4X1WbrPBDJ8mpc09PULs+qS8ptBSnl3ps9+5xjGOmZvMNEOQcJXz+DMcFYD2
3wUkTTViwFT2N9Dh/ybgD6Lnkag5LZTtcBt+koEH5QwmtAxwyUMNrMPTRGQ8JW7V
RYiGxEazESo8Y0ghOolG5+mx3Abc9szrrbIsF7QLqmfpn531KtVNeKqFbZaOS5oF
UQRP1YOyfHLy/Xa5r2k3wSpc7pVfeN5g9f7Wf36vlN5ojFNCrt1IUSLiGvN2WSST
+g2ZWAQvJRMHMDFXibGbC6yObdwOUFSlhhSsLSOQMrXvy22iVc9hl0lVacchnGBa
et5VJTplJt4Ikb4Y4R58ttVorrIz2FI+Y9WutjHv8KKBawXQrDtOyshM0FvGFrb3
XTynVoLwaEy9+RLFHvuN7hFWnBX1PL2q4s8dxyQdRB2OrZ23LA/YD5gNsEKFS+fh
xlbbFtcxbDYSfYhqQaq7g2ZZ8wrAkOz5cOvHSGnplvjY/lrGSn01Wp3CTmpzVRKv
zhi80hwbWJF4exUj1RAV+2Mmj4nwy1oFJ1nqvEU71elZb39Z8E6uH5r6X9wM9tYk
VMWaSugtBC8p1Ld5Yk9msbM6bj9IowThRuDqx2JTv10LugHhprd6lt6X9qBlRS5R
f7HRXApyLlhgFqnD8ckLmN57In+JNx+6b7IRAEl7LCrcQLzcl2lYm+scVhvPiU8m
BGsJIYLKVv/dYljZT/PoFHDIf1IQGQ11EN+8EJuuolCT9zxRty/8IS2RX8B0cmcC
Wo2k4O9L9LKA0l+cGXm/5WYUZ5OkaX1kO6pqN/M1S+0xeEWTC+AOyU90V0hN1w28
qOxDOLPr7a34kBYpbnh2ZpZPUOgvmMw+RbD+ZGz/ikE3g8VuK0Sfk0ip00G9Wsv/
cuADHoVxoGo6DXf/NkilPJT0KWZ2wNjTl8hCXM9aGhkfcUmZ+gVjtIOYEBOc/mDY
fAQgrcunlT6cNJa1Kz9U5T4YA6Qw8RGd3chFYsu+cK7kZ0zV/kWn3vJnLIow9Hx3
SgFCwb24B1IERwOnEd/B0JOA0OOfgwu+d8U6ScXP4TSJS3GIn0piKtJESECeEcD6
inFJ4Jv+bu1TNcaChBfSnnoF4hnuH3IgzsP6AyBzRW6436OsiHVdz/aJf6E/2+2m
n2hX9U5LUp7xv04usG14IGsF0NDq/5UgBcbHAK2QEzg94SVNdG2cG06c3deEXkOq
ld7VT7it9xU3iVEpDqRRu6CFzALy8k1mmEXbnSo3y1PxY+rYCNEWm2iaBkGzohPv
1jLPcA3W6OeQVma277k40jP+4zGEMm6WXqjX8PRYbDGht3ViB9AIwNZ3F6KNANmK
4pJWKaWv9t1M21SUgL6hwSu5BUCFSiAdVRXft68fbmzWRLG2L7McKm0oiOuQymVB
QmOEK+KHJynOwZf25fB/8/bNPaS5HsvG40WpzXIgPwy6/doFeh9YGbLXgx/X51rx
IU4Y8sxhCK9uEh7JMolvoXaaN1KBy/MS4cF+IvahailNqWiYLDghJs0ZTjns55de
b/CyqU8PToS07Lp5zfAMNbT5AMTlfne36xoXcJKagOPZX7V72i79IQ3XBqP4Bb4l
CX4lEgo9VLkMNpkAn7vEZmfGIwbjYJNtHlDvGD7n+miLWbWN0xxq3tOk5t2lOLI1
xUlZv6TqgYoUHttjnZqE6QRjhgj8yw+6UNHrv44X9RThgixDSJxNTvQwG6gDsWmG
DxDyHjUbh4CHBuUFapMkRqBUSfeStccVdQsEBBwTirwst0uCRjLuNhuNKvg8V2Rb
oD2CV2iJKK8wLYG3ncL2UQXmyJmzlu/8AqfAWQdFZioQWBya0rIPtlq3IT9lWdQ8
PbGkic7GkLb+ktm0aiUwZkCw4aG1KgReF5bgonFgp17+zguWBNOXx5eI2zGC4VgS
sqRI+R1s7toTlyCW7Kts1Xk2CUMnHxZwJrJltPpeifjQk/os5t6tE67PzUoboYrR
qq0OxUO70zjtQPyy+OYsgqwKD0e067D508SYT/rZWMAgrU9yCrCW60/AGnqLLyw8
I4vcVC2OHp3lDzWNjVoHK8gOLubdt51sOKKs+Eexzwkf/AQ/Qac/MUuSFIqqn5Rn
ilowdgNvlUrx42H1J2fsE63ovS1ggQ8QDoivW1X5Lm/cJafdLDG/bh2w8ndZUnNl
EI9hPaHH0nBE91iRFQ0G/l9QhOTsA2Rgh+8w52/5c4XWpBJ8qUazo4NuVFxG9tC1
4ZjiNMDRDWriuemn1py6Wd/JyLAmcCfnAE3pY09zJtBTjdsB8YrWec1kiK1D1/sY
97awk58qMMZvLzfi8aRnIgerFuSMSuQ6DpAPdTdpvt76O3H9bOJxlMr5mFuGuJI7
rOs+tjVMzKo1YpkhsBZyvWF71mphFuDOvFW7unw2nVIqYN5WxBYM/jPgdG9JHkPZ
rPmMkOPWhiGZSkrEcSm1rOvR6jgAaVc2Q+YlhelUiFFISWvBHHTkXLFtokvs4ZpL
cj3D5bwr37xAOzq6HXG8AabRaLO3yc0TWuwqPR4VKYd5IaUL1Skzt1sjuvZRT6eI
CPxgB4V32hmv6OBTJPMN9DRTY87mvRD8VmaZyLQ3m7kARXiH/yZhmM/WthdLakr1
NThnB0KDuhVlgUz4j4DwsIO+Q0/4b2WzaMSwa+fmIFSCt0RgSi0aTb62N81dpXML
VqzjdzJH/tylArnMv8EQl8VRNInyGaOaqpCKP1uFV3iJQybDj4l4AWqVJMRrHcbq
eYRjTopmuZSJNrlZ8ZdAGqicjx+uDoULy1CSdiOV/pibeSkuf4sC3rWGDL2FUuJH
ku5sbuhvXeye3dsbilNWOaUAUFyj7KIuzNlj/6mpMHSjPs9Y5t0fPV4NFk2seJXu
REd+abQV8xR0f+FOJl/AGqoEuIjS+HomeIqXfVXHST0tnL5kurr2IZr1B67XPU06
iqwOsXQ8xvUpTBy6+zpAxLcVTLI53nU/rJwQeWVMaJ96USDMfvqxZBF/wlSY/IfC
pGQzMT8+Qr/z8CX7x3xee9gcrwEg354z7Lz0Dp3CdYBNCvByerDyzQuKX8Lw7SJn
JzwH970V0pL50EBeICA67f3MD0Cko89zyNw1JK9oSIngemygdjDdR4NTMpb8l7pV
/e6Ok5Ppfymlcb6n0ueVjZb6Ug/CK1Yr1c8MXhC2c4LZGcW57OmX9Mzg34FXbl34
JziUC542a1D93eU+nqtGA3iK7loGWie4sBXCoNCnlydP3ZUO/JZhfkLFnOsAPqR7
lPaLjVGFG5UFzJYgMzxNyx91IQv/nDEX+aFeIdef3sDlvjRQ69ki6UbHz1qt7zvH
KOMkhAWdYcZADRhQekaQ6VbAS+eIBTE6/nkFDvzcTfOel/cWdNEFo4tv/K199fPe
rnck7eZTBoUgZ2ruUbulHEBfoPbaukRyzPlVjbRF5td7zwVk7/Sks0DPRrLXeI/m
Qjp8jd0ocDcm+liQzgt9O80/4JSstlumvm7S27Uvl7rLBR7KwqygYrgW12bCRuXL
Hla1gZFz1aLYqL5YBxKpoZFMELVjw7ndDhz5bShd/KaNrJ9rtamV4nn9EyxYzgGm
wM6mwIQinobdorbPuBsRm9gIgVdkqqZ5OP5DWC9nf3WYAunpE0yFnSf7aP8ZX/CF
pRTFWG/70SNft7HWcKQts8XDPKy8AAoUe4iOMN9tyGzjCBK1THvUXoIwFq8OqH9b
uUNyxdhloAZCc86D1aF58k5m2X5qq176YtSUnDs106adIO6+AIcroOTwflelO4N8
RU7F8j0UMhm3WkL5BbvywqCJ5BzouB0H12CEmUroHgfXUGPP9AxO4htZXeLHgZFn
ctWQpof3i6sH3aAP2h7Z2fR5ADM6aPMv/wTU7x3it+btzCjFQdVn/xaj6GihWbgI
9WqawIUb4lxP/zdzit8eqk4enllnkPEMjLUtXVAf7FPpJ0WuXrkdwWbgd40BRtEl
o6diJRlzg9jbm6jK5mBt3Ha8q7lsX/42Lfrb4JFoa1t1MLEBK9Jnc36+IpTjDGAB
JljtVIBu8Uny1x5H8hX3SYWlaUIttb/gAAgrUj/tfKdcsdkwwI4uYNWNN1weVCP7
Y/p3Qbejj0OCsAIpzgHoaeKc4iou/a2/nD/W37kLteFRFNSWCdhL1wP1VwbZe2p3
fVCQAj2XRykUr7dmIMOcUUCh3WnBJaA7kjNhMLBygiAoo08J4WWtTFojVadHoe/U
/uAyaEcwvMExWp9TAEJ11/LsdtSvAUsHUqQaYCNmDfg1EpUKQWRErM8Ulc2MkH60
0Qj50j+ZhmNz9vy7kaTlUa6j3BB01wdZApe5y3At3PlJz/queX3w5mT/3nfK6o2r
1iO7QMtHbpWFQlgfSg9fyRGpwxuroiKkEp2N9rCfH3DTsBxQFnb5Th+8SPCrQKU0
bekH318GW7mO2TESvv5u8TRCqBid8u3Ck66z7jYqN6XGUm/mkcI83sLdy0E/hDqT
IzLit0kPKtBfWnQlXz0LlIlWgJPAzSuevPjZzWGANt9u3DwmrKFE/G5wbUGLEH1/
/Dx9eq6lJS4As/3U6FYpiB3Pwspiv2wv4v1S1ZpH9JibbIrXrj37SQN/LomOJ1ZC
0SHIdItLSHlkQ+MVwwUm2WIwvmgSJgVh/N/msZs0kU0D+G5i3ObCFc4Wam15kM49
Yx8hrBQsgLQgDk06fGEErPFHPfxf5gM9nR7UbDxO6LROhTHDciPhxv2cmh7SHlte
X8VRZArRubTlvx2K+EH2G6D5tugM08nO2Cf6G3qNCb0YbpCMHKn8RcUEgcP4iqfg
pseSk743ZJWRCINuZRX9HQ0TRdkvKyJ4c/XmHZyas4ukC4HMOJ7k9hivLIN0gJvw
k4ZeLS+zCSD6nJiB6KC84zjDBNwpN8Rn2MXycvJahOIX851vV4bv2ayzWj30BAIG
CT5hUfN4i4VYd04p47Mj9+u4X8Y1bDRpqBWhxxka8dQi7Ps9/y4LrrX/fshruo3w
M/4Lf58VX+J0z7ce/sK3eNVI0zFfjr/DFnM2y5+AuHy3ymXBPexe/nJYn8tw2WhV
VrAQ6W2wZ4jjdztCGhUcbNsqFmkGW9Dfh/582NhL9jnAy0C1a8JW+ectad3LX2Cm
X+axj402qgHAZydeuu9askJNJwJE1gTtnTXz/8AsrMIUG9ajIbDlE61X8iYsmqJK
HHv0DRVNv2+dLgnxui6Fy8jHK7oOIXgRkisEaIeiezmYV5wNXu5aS1VaPJFgkb/G
HcSJ6Ci5+/3rnoABu4DaWF33r1MtvFYipNJV08aC1e6Ykk9co15BojdJ8JuBSfc2
EmeoVh7y302VH5p+QKWb9DxQ5e2hw+h8o6JUdhUZRo3S6e+zOVVae13lGOOX5sKB
BpWcN0S4rIyzeXb7mjztN1+KqbD932iNqzEAFK1XoKJAY/Zew7cJUIHBfjzflUax
4NBr58ZTfbJzCxrDtO0XBZrSaM/14OtESUz9GKUH0teZvA/XzR3Tp1Jn1ttVShGC
izeOTwsXgP/Wj5hSX+n+hG7OXVu/lqBOXeSJaYHn7cRVejwXOO5Q2hQcB+zxtKYO
zrM66jDgVnT2RoGa8QRxn7JNVvsF/8xivF06D0B1qYE2E47ZyzP6to5ru0O8/OBf
jziQaLn91F3IArhnI2IUAhdKgGiVZeEm+6ZQ5RkuvUgdoPDdJzVnD8wS1fGHsR5m
/FlZwZMXu4PuRL2kQhD8/Dli9LwT/itOvUulFf0AfaqkAr+Tb9lLA06zp3EJ/7Um
42KfTdiCZJOThPDlbz2dOZuER9t3K6zXQimwsOFLpBQFvgHBf0QoA0GsILV/ZPTZ
zdz/2yxBeb3UwKsTce2kV/OwFbxwxTaPy8CNSQCJWga7dB/QDi4pHJglKTgbPhTZ
WRnk3aGKKl9vhq+dYVTPBIOp1WUvlMNkTv/b1HXtHLy8LOjTcH2zv5xl3iG/xReB
w6fcP7wzVSrwV3/4bLyw8w5kcRtNNbygteHF26wQnPEjaNfM399FNIoputA9wDOd
i+unR6rMiK9jskK/YWELHyLF9nttyuUFO2wuenw0nETkeHxcRXqWMwaz8Oa3bCFc
9xbeeWP/c/WyEnvtC4UETOqnb2f++GoXoCaXlL2S7USd4uwggR388XLRRpkh4AY9
kjP3tTsPgGu77uBFAsizgAdhyhxSgmhmdxWhPt5osxW9b98qHdx7/+wrY3pEhrW8
nPj1HHikSC1xlvimeHXiWuZy/q0owY/F9oOlR8VAR7sNNVALbSCEo5t5dgG9kah1
RfdVADYHXUsZB6yQraLt2VJyOY5ghCUxOBWnZ30suMxgult7T21aJMpf6dcaCaw7
1JVH/K2vbj0zHDgRzQv4EykDi+0HTB2PqC5JOADGgLeFXFRvOn3a5sQyGsSlatID
WuPRY9FDdNijYYWaY94MEyW7keBQM2TEpQui7PUB7lTKbACsvPuhTuKjr+17K1eR
3uc7UrLBvFY7qW10zkFQRmZX8b93kyPAc7+70zW5iCyCPCZKwdrtS6153mR1s7/D
8r7i7M8ssXPX5QOPKF0A8Nldt8j6EYBbbifZxC7PXmC5bFzRFpMc4+BfL9F132Q7
GFZEMAjNKV/sZYAr4uyD0EEY2hxTa7zi37HU4uCsYuICSi81K5FWbk6LlQtJf3XU
8lhI6zm5D5kD+b8SN4X7nUPLRqe1XsDCZ3BCcD9bBiU/3ejSuhWesZdqgn5KsuGM
yzTQ49dSVuP73ErHKFwXIUNjGOwhAqrdwY/BQZuDQgm228LMTokI+mZ4RlQKXVOv
3g4hFxqYUZygHWzLbtw1wC2nADeITiezdGhdTL3eNa+0qtQBP7jMc26pAB6W7DJ4
NokvB5p7ZFwIxXh4R5PksUuFqaHHfeCm/8tovlEOu4Vnl+fRMeVDwX2OgVE8S18V
hWzaEX8xm+8SJ+VKfTXeeUUMsjszpJkTZr7xAy+z7vAcfKXnNyuQBfRHjXoG7ggn
TTX17gn8+9xJYm7VYZV/a3Huoe8bw9g+5D6buvUmy6b3reyPEEWrhKLsSbdoAZT7
smokVT8j2bXcGY/21pVQSHAT/gbuYrx7tXtKRvSpB6lH7ML9nDi9cIcpBNHmz7Nn
lACeRH1gh1wGzYyyu1+HnEAbMNQ418LOnvrvxm7ZnjU6dSBbybbZXXAI72IJcW+E
nWOtuzdJBlWbmDn7W2rUEjzkEBNF/KCNxYGnbmssudCxgguKNlXaJryFDiE4asJA
b3CFTTKoWbRYHHMCaiP4s1Rf0VTo7v4tMOBNpU9/LAL/3doF+RR/5BxdTMCAlARa
B2GC+vr7t8FxPSGUkS/PMRySW1jdj6BBiZfaGfF5z2MuZNtkuXVXQgJevyXAgFpT
On0r7x4zcBa/7+wwYX7XuhGT7BKZfQPDtlvYtO1b6lderlV+mUeSirh4H26aFWdd
CCH10pOWNo59BeeWm2avv+U3cB+YqqEIG0zo5E3LC4oI/Fl6eei4PAEgnFkeVx5F
l5gRt0LGsgAvw9mPF3/0drhB5zom5TJN9z0vOaqQbIZS4JqvsnZwqs6xU/DiVtzY
nIgLn+49ziJ+iCe/o0hvr0uuruRhEjhfnQh586Ft4gfD+BzxT8NRWMJg+4haHj8a
00wpGzY1zVncggfNqAFlvq/jNn7MSWTk3V9YxVyTexlqsv2eF7uNDGLOmG3BKHm9
Jpn37yXuUpoijqIiP+g0mU0PjZOjA/qftdvDZQCEV5vpcAMFKHe3rpVwoLpC/UHx
7R36guj/m+vQa0NW59FrCp6vQDv/ihg4LYAANzdnqBgAyQNyCCvqgbYoimCCxrYG
GdrCPBu4hsQ4fFo/Cs343RwP5DwvPtia9biJzPd3AInAgGdQxAq33acfS4EQoo71
QQ8XYdQywqQw++XVRs1rTDE2irxlwsebg9KxnbdRLh2F4U6EBad00oWc5CkSLjyd
6ODxRYXs0CEEILgmH4p7KhK1UDlr3bK5TPXhdFEpkxfBV+HweKO+T3t8+Mwq+CEU
42a+gjaVNCu9fGq5JZDODraMkDrnngf4KRgzs1BjkBz3lbB71rZeD2W55N5mWAcd
7boYhOriHoUhaT4//Y3aSkmzU8jp9v+ggb/C548YbUxTaTK3Uxpv/48a4oLEpp7B
5hmf2iTKRnbYe8025uMZAleP/IS76uDYgkAmptkZG6g0jw/aIZPXZSXF6yK5ZZm9
oxENLTrde84N820oQmGqgGTRJfTgGNXTX2LCGIjZNPKhlEgEMmzpwuHK8IUYHt5S
Axe5c6jVApO/0S3KbOAeDJ1AulzVMA2Wfg19Rn95dUioYxbsfFjL8dsB0IfDu1iZ
qr7yN1IAwPBaUHNyDo07Acvvx3c5TmU7gWQeUJHofYJGGV6Wn8goDBMpuIr3V8XE
2pi1xmrp3pr6T0+cd62kk96zjCJGmttIr+pCbPZOY0G2GzWm/W5F/3kKvNlIANng
sRpMingFD7YpTF+UYAWoSf8fjNLqNIc90tH0dv67eg61dXbyB3TQ65nD7n9TIdSs
9byhtyHXR5hm/QMXv0HoLMUHLMA769D6gd14rn0UIBZaomMfEwp7JbJo49cuSP5K
ue4QQYos5VKnaxjYSuWgaL9P8QbnsHbhDx3C29FWJwkcZX7g/qhCAii93FRIkLoz
knC1TNYO1ViyjTrUJz2zajq9igI3i75sAx0IHbsR1hL1Ro3LKJW56fqwO6OMTkAh
9EH5lEh9mhKkhlDC6PXMAib2uJjuSg4AczT31zDhbRYyIBffy5DHT2ibOLIIiPmp
j383a9ADChmkCorrURTIHOs6O7diTWHgD0AVTOaGOcibkcZrC8I9Tqx6U0l3DRQX
TLCmZVKlOU6edXskk3uVJo4W/ssxn99RFdfC8SXi8GaCyiVMxPHv9lKIqmlsc/1p
+OGnW2hfH2OejyVrPbNwDyjxvTS8jckyFApPgydAYslx5NAM6KZXMLCHiC0hJwby
JbbQMnkR0iLzOiRRqcF3ie+199CQM1P/Uf9ok4tSvsUWkS3yINzmQpVRACgEGoHC
9GDu4kS38AZRXelW7tFavwR6d+UDzjOmddKUifCbLcBWm3GfoQykLB3mwAaPZgpt
uUm9xE2NM93fUiG8nOyU0HzFZnYx+Db+mYfXFSfpJ8meHQyoMC4iOXyOOhYZCFeT
fBmwVX04SBfBeof6Jh9WYQirP/bRO9pKEdujFjm3oTOiHMoulukIXX0e9ycCs30Q
7ywOINRUwuNLKTxDvROlVyoaVobXrYHxP3kGrjeHH2wtUfx2v54nmMZ2Iiz7RDuw
D3ByOIJbaq/EImgNlw5OaR8M+OUztAj5EwDT3u+YWW544uRedaYZ22IT6KoOyRTa
dOZHS7LCT0p2Ov2FgEfQ1Gxba1kmGc4YJqi2D1gL3wSBMzFBZjHBYXr5UcD10XXL
Iqb8eIRTdzeRsG/mJLHsEriea1l/r6OlJXLfqSgAakiQixMkI1u/o782d3Y5hlxU
I6j2+kAAVIK1snjL4jnS2wVaCmNAUjcw89DZK+5GGGaViVHky7Z7K9cU0q1U7bSx
iz/9+Z0pJemqOfsHVeLZLXE74wwM18oIn7iI6HYp108AeXdYqNJtKjBQ3U+PpjFk
VjKa0vpn0/Nb53I6D3zOAXCDrKYCaCb0stlM9sxMYuxagfKpxKeOijo5LuCTYECt
oCRIJ3WQkpmIJ2ERnSL5EkzxtvzvgF+x5M1DVfz9F0JRP2siL8R1lom9445pWv5I
+Fb59F7eNmR8G8kgA1D0Jwhd9Iwry/HZZaKkK9B8ivf9CDUH72nBPz06gQGfy7pa
4JgOzrere1KATvosIH+AYnEnnBc+bppbLqRjGL9up+RuGV35k4EmzNEOri9gn9Yc
egD3J8Fjp4l1kT5LenNTwkV2nqBVVq0I0pkkXcDgq6Gx1LrBtOu1nIWsN17up9ae
oPf+EXP5NQucUE9+X24OGeG2eUhrSLfIlNamLBbuV66NUiP3TLCXTRRenN8F6tHj
ULTXDn8TJqFQFUZeBScymB3OOwqUB+jwx2403U3+vWBhfDAjOUvFPt7syZQAIgMp
8Djr13GHAj/aP36gvk7rab8ewMsKG4HUVSfVm9IbBe1SkLJI9pFcg6VQtPltxtxK
yyGZZ8qqBDT6Dit7/U5otcc2YzgtDfS4zyaL5saS5s57x76hb4DcgrPvTkV4Ai40
Ek9/qr1dnd+oiCXrlHDAsYAD57Gw2SdvLzFsVek3AFEo/Jgu7Q5pDlZM5bGQL/bS
oNqLg9+IaAz6fRu5qm7g7RihMbDNnh1N7Je0zrd2LaFivM0h2PRK8ryqBxmLvurQ
pRoNiGWpNZbvl30TZLHG04fEoM9TptKlRxZxbp4pEeaTvxK/YkvJmsPcB5khXGkx
igkct0iB4Jf5haUhl3Oi1KXxqee9k3cDogYMEMLGbjNnzBSfTt3uUi5jmI4fIGB9
Wdd554SRlWrvrOJaLs9I44NON9eCbyM2uup0liJGaLDOiwQL64ekj2aJcjAssrTS
JlCFnsFyxfSyS0b44VXljSfHDvlPLUht3w6gpjI4klW8M+enOFKc9dspOH/MV1xv
LqhDGGFVbX7BWiKzX60V+mxQ26zUDYSr+OCQNwKWc+9QpqtY1FpwAuz3hB87NCYu
xZe3RGChlnJlOksTZjs2YdSDRW6juXpowHU2MDRotLgkr3KL+aWNwkVr8JAB1Tsw
nGXUO7OS9xk8QDcmXyVoi4k5ziChLQlMc0Q6dX3Fabn1xwazOOxsZGr2mnU0bc9y
c/aNyS8nXs+p6iKEwO0xy98Tmek6kG5Usm/4I226hlCAXZNMmv8chopqwuINVkqv
uQkrTP0bekD36uFXoctXxmA5CIakJLoJEJ96uGgfPawI2OAqKgkmvm4bxQNNZLQC
CC5M1220fyVr87mHrdSPJWePFcyqH0y30bDVOQJmyMmbwcDspm6j08cTsq5fTdfI
7eSstxGUbCI2G1LCFB2K5n/uL8/36GXA7DhrYFWRb3doPN9Vi8PdfTKNMb/1LFj/
0l+P+yAlEgJulocqgVebLNcJSBngSRc+Zsf0gNWvZ78rKuES0Wv/xyHPIFmLtm2z
OV1+sUSabWSrR5QyxPJX4CxQp0+UG/tqN2pKK7PCUYZvH0RyqnkHyYsIHcEJmRw3
R7Qk19uD0PR4NbVJ1m+9TVs1kVvjaJTt55vXK8fK768GiW2t4n3d/Ni2o5eFivVS
lDvsCz5S24tBuo0aKE8hh4O3kyTXMpuFoOz+LolD20AG/QjULpnmdXmupqKifdmH
ZLwGsABwvNZwBZuqNiYyxJtvGBvq8/kiU+yRfAG4bzYyyM9TCbPfVtakoaf19XFM
9+saQAygsW+nkA3B9rJe7uw5XsEgVnGRK6s0PkQHigO26QrZkl6hrAqU/iD+ObRl
jwQY5s9aXfWpiRdSWaPFtXe5LZAJHdTJE/zKCEozxgE9Jx32TaUPX5qUSP8JKFeg
JgzEp6X0YF/3Zo+6PGYiB+9GdNFJBCfN6JjmUDEJZDeTApxuKxjZxFhkxYKOPQi8
heK5bjZkTAwgkRIGLTPJshJMbYaeu2T+/MOwm4Mn1pykbVgYqvebSzdVzbq8HtqO
cs5GsIyceMtVWCogzhAIHJt0j4eACrAhAIizzORURVM+Pie6KsqrOdtnmb9Kl6Iq
qx2HsJ82ybvZJqi5JVKEkXhQpp+RvPMEFxBhShukY7x6cpVVFJfMj/Qs+j6lkFu0
GWkPh6PIEf9TcjU/JnpgFyQ6a9UXI9YBcOAaVXczCs6z68rsL/ODo8hSlwArKWqL
BkaoelDcTfvZFUmAi2mkUxDlqMoKyhYShdLM+ymO0gOG110eizYLjH+/kM9QSQPx
yRfOpMwftFqf8lX/SgrFweTPM1kuhu1w6zFFNhmiLSTUmhibfwqHsBs75DsT51Ew
/vbTWdbm1F6EM1gJy3UM7D5AT4ZK8X1QkTz1Wq3g47l+wPJris56bkn2PqLwFagk
wMWoGzPNRrAL1tgtl30gEsdGm/facnnzTcqP5utBDMomo1naE8wzE/aPi4aU+s+Z
qKmBLv2o92I/Rs3EDflizRsLPQcDisRfApIbN7AqnwE580XqVBZ768kD5mlPG3vR
ygP53ghblfRPMacvop6CQ7HboNwRBHXiBmEDoang+vKp/C4Z4qq9QW7Kw0FvcJSW
9czdG5ETP5fyb/8fInQjudDEhYfYxCGwU6n/lL3UQPgE2BSl52JaZuGMU0OyXMjS
ouk3zQK7iODAMsnT83K5QSkoHW9mQQO+QMlcyvzPnaQIfES50lctIH4IjPI11PII
/yfGUQO38uADZPi89T8G8zrxcR4Eo6PHLoXQ3yUShSLAcWnP3MddIR/K8cFNDawT
cliQoQV3SDOfabZ5gif8XjJFPU/ST6NHAXqJnN53C0ck9gV5nVGQ9fdyQSxGu2dx
NZ6/QM3bOK656+8nFzD1rLzrIZ9vGPzbNfnOwc4pwyOm4cJp6u2cqueVAw4ik9Ms
96VyNOS4OwwD4vewthe8GFL8+vXoJe88K0mU7MkI/dX2lhnVNC6nX1uyb1we48mB
Q+m/ry4FUiUfhzqFKDe80oNsNZd22uuIjPTlMeeLfr/6G2+ljw/dWQOYY0BKiAGY
nAX2je1L0vfbgAQTnZD2mwxqzrQ51rOsncqrnr+hriPMthgiZ3kcEeTZhIBazzHr
9cl1aVni+Q2QlslfqrBXiY2UstrnQIK3WnWRTTxYjb+57g0550F9789D4mO8v8PT
Dh9ZNj01qJUlxebJBmhXju6N5hW+/MHZVpeFKhQ+pqhq9cgKK4JmeZwALXd2ZH3v
l/sCe14a4IVVNtopYtZE0v38PJsSNBLMlt+wU9yes5I+Cl2dmQqnM3IWyLfGLgaw
0r7PSnsHCDdFnmlVgR+pzNcYde3ZMyaE8jsQ/s3EOC0u4F1FZafdUZl4DwPCuA9u
anhhiDHenjPHwnbkTr2E9t5KuXr+rR6j60mu7ReQ173I1uunoMl1sYytnrKm00pC
rMpAy0VNd5AlaD6pXKBAj/AS0TsGZ9t1/QmK7logGJGTFxmV779ZTOGTPw1JyQKv
a5RCrYu5KCkZ1lrDl05MmSw+TsniHVHdIplimACsM6OS2zKnWvol8efKH67vXg1q
0Vaij3DYeLp3PVnwaqYEplmXDJvcTYx7cfTvjtceRKjVZm7FqlOowxkMH4cGfisP
uCOOsKMEvUj4vPXKdkIRo0DSFhtInV6/+izjyaYijU76zMZ5TPKDmU9+4nuN7MZ2
bYfaczOHrqvrvJFr+b6sh36CSLnOzZJjVxU0AIIgkFhtqXifcUXEu5dM36dNE+gO
scNsE3+2bCLnuB0CPr4s2T4GsEKEpvdI3Avn/b2wu8Mf5Jay/vKdE3I0ZkMEsK3i
7ysZRo32nfcGQXyxI5vCpQnWOVz7qO5I5UQcs+bJGRNXId7H0qIoTndknyXy7ogL
4eQXT6f9k3SmdtWQqU0U7MIFMEido9i4MPnce9GXvE6/kZuX4IlBNBt52NJQDQ/Q
mwzjckXDxJ703bYbb//qX56TeHiXEwNI38vjB/aMZu/L76PoGSiI8+X3hdjUo0Tl
JCe9G8oPIDx1G4gnaJfVZruObcjpJ+AlOlUDSnhCbrtjM1KGilWGTJUTkMmqQxDX
d12gL3SWFyeJqDpBiE0Q8l2BTlIdODoXvfllHqVdGcx3+CBf+zbLa/RSOWT1JT2f
p3HqjcKBopJgHmbfgbQsaTZ4kH2GFY23iE2AF6UgmDuYipviof0zvAJ3eGeCX1Os
cTjlQijxHX9JwL0pCDA5VXOdSaCPJ1/Io+cXhx4cwbh35KltHIsVHueG25zycoC2
+TH1J7bHb0F4jKy4nYJfzPNnawK54HKy60hz4U8+WjuZSjra3xxDaGvzJy1IUu9r
SgxRv3/ulJbDLgU2woDuhlYdmXmippS1B6rAbXyv0JhviJFIkZoNyW8MOgM/V3o7
V7otgjby40/uw3kRZeBGrZcJFQIJ6Mn0tMoNr8VhXvhVEb7S7egRVgPCmFTf5W70
aS8ELCn+QOE9lKmiRnjgtU6itNouFnWxq/CzhaNVqW2KO6Jrgkqj8J5OBxUxlHjf
nchLpyPXb6SUS2b7N4ZfCuuWeKNDK/gGKFk4xKOa8n6gIE81zdnzjFBmDV2dfRnJ
rTyMJiTVU8sXp6QldG2+gKauzulwxDNHKYxtlGWbZzLZFjacj312EiIsWvdkn9z9
6dI24p+151bOeotezmX/OluIuxx9mc9m6FVTe/1ZhLWJBC5BFv1O9zQvrk33veum
hYpiEJ/Etl+C8B28KYIfWOWwYuVjtkPJZRZMfUbEOtT9RTc7OIEvwfmgVEN3Ahu5
PCWk/T1uyuMten+DfN+Br7XmZkIZ3WWss6yX0K8cnZm7zupjWmeexH+XErLMNLNL
/BV6hmmMl/6BX2rquTgVQBCPiVt7bKUwdFIl2yCWgfpKV43zu+ujKMrRZ+zS5FrG
gKQHK1zvRTh3hwfC+/GDBu8S51sc/AHix7/aeQXoEdXCv9DkPqkOMwxwjVbT6Pu/
c1N1IGs2fesQ7jYyV26vsqHC7FXG8fsS2kiJwiQXUfMt9/G7M11+YiLrf/iUSaEg
jFprYU+5poCkWzLAExmK01xy7FmHukNY1zbxJ90eu/wdwfmT1ktXKrs2c2jdfTEI
o9zDfzusLsOlp6NxsMqJ8Fk887iawj1nyjOFsPd/h/8fO4vF32NS6WCD3WuDN+Pw
KWt7XZ+qUsvinYHbonXAQLb73ZO4ROgYlqQ4uFib8J1H4bRcvc3XkoS6zUYZFVt/
oLibI0DLE+qoO4TOAFQmEFb2LpHPoWP+QJHOfWEaZLlRVxlKMKnNAVLaOO3OkI/g
ob4X9dnPNLjLsv55cgUUQ7IOBAsZsw0rUlBYekf285HFCunuAGUqgljcMkEao4aN
eJKx5PtYacfxYQecO+o7mpjc4WmgAlih4OjpYymJ8uXhUmMnxjhVJQsKNTxt373O
qqHbtTYi/Z1QhGehekiAkdSJoCH7shim3etBghSLmgcZv0My5qeJ7lVleZYDcPGl
QEDw2nnBvVQajZhjymijRqIlRiadjAhNlmlti5jal0wABr6jozg7Ys3Hsc6BYrk+
bYCUi+1VTsK7tRgcCRkDwUWP93vwqoeiAc7LdU8PQ9mL+3Zf1gA4QvxKFAs6nMm9
yauigIlaV7/h54YSlPkKdLky3TtzGN/KeuUWnKbpockx8vlfpglKDP4iwJ6OAqD6
IE3nyi6TtS0bn71x2GIh7lG3INzbWNH35sv4ce5pQVD+CHIfJirWQ4vfTudvoR5U
pfZnynddEqzTG+69i5FmgnXFgH1xDAWXfdVdnpCdrUZV+4Mm9/Qq6rZEJxS/JdJt
ZhMAN7xo88ultzILCWe5Rl9+FqdXAn14k8W48i7BJpqFsCMKNzpHWmV0++fJKdtA
ZGaYSw94mx+KZZTXuFBWHieTlgSt7JoG3GrXlaLr2EwHTApTM6emw4MnnXgEUvNV
trq+xOKqEo7Q93xv+1jFADzs2jM+L7yWJn9MsQjRLCn8PPXC9z/blrP8MNJxmkX/
nEewPaeOtKOV49NqJqDh3BWSB97CcwlkIkBsYF8+W/Q66lm1YcIybQdnISEy8JkX
4ocXGiCJTQ2KMDrpK4ZZftDlxJGqe81IPwb/tAwuOMbI/lq2NFI6jMSdW43mwRTZ
nV3vVgsCBQW4pVae2MBnDf2AzCIoHfO1kBwIwbmQrNxFWrqm5JgLjRYw/53VCeaK
8hlNP5jFaLNpZNNanrq9Uk3Nx2bwj00gIePxM467WcFk9oKUmICRqWMgk7g/9Yde
4MqQXVY7ZPim0LDM6NU3g7Nv4bXJglLxttRMCRa7d8MYa8Ix/D19MeOcr+mZ0Q40
eq2J6lxXLphClOVpHhCorF1/AVXGCY4KAFkFH4m3tdhfs04b/ecEZ7Z/91rkMkug
nTmcNan/Mo7x7L/QRLbesBbXroqLIOKKMW0/xUJ2ox/q6/M/uNF8G2/xSMPl27re
W4JPkWEMoc3BkT7U84UFrRupW1jrYkMXOVrEgsG9YHHWKc6yNmij2Q7/jg1U1PTA
cBN2cdarR1qWXJS7+1DviVC7OYhKSA/Dw8iPJnXgGsphyOvrQ5wbIAL7z3IZTj9/
R+eETjaU080SSFq9wtgLSpSPcHLT29d6Cyn+n1SVyxBfCqjCk4rNUe4Inc+w4QXr
9s5lNxDqIu79gi4UhiWr3zhGEIeFQso8BJi/ubk19tzEHGtgrmWQ21JjIAZ+/FhW
KsIu5iDCzwL1BgTgS2hA06Pp+OHI3SaUnZ8q8UFR5//VWLSyIoEE4EFa6m6bURdZ
gbrPOKv/GTWDG1Vi2iItxmvP67equ29G9v02OTXOVleJ1VEIs3hoAXoJAcAPttlD
CPtbgso2b6FGQzQjwHZQ6oyeJ4gdo+CQC8VMetBjHbCxgzHIHtI8Qd7sQw6Tf/T+
ahMo1vOkH4pBDTwGcZj+Yz4jP8HKmn88NVUH0PmPbUQ3bhu39I7bOpeH3T4nVA1h
7u1CLnVllKO1/XVXPffn7g8f8xoqDII2rnsRY074bEroErmEtipuCbew07LI8gbm
5IVwkpKsb3dPyVLAI7xmhNLlzmd4GaVDKAdNke80/PM/A3bdXJPJttbn9NvQ69aP
8xXLd3T5hLtlzB+Sjm9Ly3M+/ymOE4RstEUvvFQGBOss+L7nTZ1NeEolMSpHmSnR
Io//R9REI7hy3qwSqq5xmPYVIZK6E2o8Aeu0u5ApVSpqSwXMySvJ0QlD+yLAmlHP
lfmnQNMn2ATHAfSowbH/kJkGkN3+yx/5s2E3pye+LGvJMhn9h72Pg2YIAAsuSGFQ
AyXHtEvlCvrLzSK4fiZrroWN32Deq+8RTwv7YVvoMzf4fyTAzkz6aaxh+qYPhHuR
l/y7rKcdY28OCQZoZzkG5mefgk1EUjJHHprd3acsTvHaTCiSnPwHQMrOvcLPFM/1
PtwtMC/NkKvzxhxsDcM0W42/hbUpjOGGg7/WtwFJdkvVkP4mj63kThfjcS0059yk
SzkjTUENumEMkWxtvCzTZHZsTq9gPSUVbpye92SHmz0Hcobfy4hDSVoE/fp3ScTZ
Q4aSxTikqFfQ26Co77gVTa45GfLdTG/EbxUnliDYf4ulEyTEpAnyr71hZrVJtXGF
Hbzg6iGPIr1Ci+7kRZhI85AD99xBPnJlusB4Sa4DP9OwbhnPL3AlW+CdVN6bBlht
/wLhm/9Dh4fBfNg/UqJ0b9ipGi8V5fKK3Tv/MrnOKZd/Eg6g5q0UlEU4Hq24ASa4
PNDQrori/mUNEwfXgrV78jwUhZy1vVnXcVSkxMd2mdvg+pLYL4/r/GdiTkM0SM8G
d7NGP7hasgT7VCUT7bU0yZ+r5UEdDDoZfTDCFTQnOWzu9J4EAYFhC6uRrnoh0o41
hTtmZ8EppRvXV0IS9aY49FwtlirjYgZ+4RLqGXCVVDmyOQPW1vHml8wyaRUMGFb8
9lBXBmC6JUO4WY9U1QL2MybQOu60NfpCsSASk818GFr3NvWvO9TiHEJO3bpvFPxk
fAtX9+mjjFZta5wazNriP1wMcFgxqx9Tpo0gyK7uqSxvPjEusXhM7135tZdxC1A4
2AYzLQehgpoY1YSSEW9AZAmBRIThuyj+ZBagLLlOCl/iBI3kzMgsu24q8aQqKQhX
PnmSniHZ9xGyIgPaoY3X1F0s1wvBFYu7QePUXGn9VMzY89IqXgHQD8k13sLuUEWw
X3wBhnD+un9aHGT0uC/yJ5WSdhLCexX4hFFLnWNXoAjlC9ycYN3MUf5ItW6ucnBg
D/GchZZ209+v/Zv5e2dg7Va/Oj3WrjQag4f9OFeMH8rVn/UE9Yct+C95kPPk3TKc
ssAJ7n7sYE1vGy7OAzyjtYL0WQlkThSRagzTIs8e0tA2X0RkBjUwt3xPrrlw/Oq8
UDIcAsb4t9CZHLPp4fssYasEh/mbB9wPazczFAObUwlGwB08ulsD6MPaq+2XjErK
zRM3yg+A0KXJUcD1sovwBGm71HD+nnJ+KtXz9IMFqj+Eis5xNBJHScx+dEkI23KQ
jJOssnDR5yxQnB/AHPdE6M0mJcUAkeQ7uvE0aJ7R0hb57Gqg5wrQj9aXI01eOg27
88ZH3dx8RQYM7LXoOz6N7Ak0AdhFEW5vuIiRUjr94JsUqS2/oxjMHZ/4UTjBrYkg
vl10WcoXmQnOkC/boP3Ytaqog6bLU5bTToRDMx0pM74gnZCQrkXmUnGML7I6X9RO
7LFhZSQwXrewFthJj1JvzVVvYEHmeleH2Ak0RSMYYwpGOmrTPP9vbzA/1vBN5WM3
oKY4VRKNrXjgx6uY/0+tQaqx8BPwSKWVJAKgKTZvIszLtknxzPCchN+hHytP5Kp5
XEzy8lNwtxT08A8c2tEzWaeBEwJtHiYQbYKM1LompPUz9hcYaHyiqjIi9MBivbdg
ZLYK+FICVQSVj8dI1EDSt17J9/0Piz5HfkxDB5iAmjFHJNB+xEhTd8OctLVH/pBB
Fpyoels78RN9YN4F7/znVcx6jd747mftsfqStWwAmCIlBN97GTuA2h06PJDdWnRr
C0q9bD9bLBLHnf6vKLBU63ARv3pt+kjNjEXQt7cFI8j+VREJLCtDTLVTIZbg2Dlk
g2gGI10GpoheqQzzAWzvBz0fMwpG99nbkbwBqlbaMWXQQl4se7poLavEtJqy+d5i
3TN2Vwjdh2qlNPgnzXpQH7uLLb7YL9CvU0rhsUAsTJqs1WOZeW7uZArpGTASR4lh
ObdxPM/knGe9/ALVEv1kZ3uep0pxCjlkKgCFmgahjpiUUoq2resoNHlzN8GbgQHF
w3Z/9pRqkAOYUQaGq6nd5gJ8rI6jZjDyiX/fmCgaii0m35m6MgBhXnQOPk1cYNpK
P2L00Z314MrW5EruLXAlj/wGf7UUiSuPVYyWn7eK7o6mc7V8R9o3OxAjL8Hbc18J
qFfH6hUXFgBlGlZ+EAqla/wYyTRgIWRMS9tYDJME+afvcaPOeJcg/QlY8Ke6EhRf
8+iQ172ycaWuf/IKbqpYCXn1LvQwQhteIhkn3YSxbgbHDBojHfqAmcRnqqSRu83u
wLAoUW5k5+pCqNv5a8SchbVDurgnUT5HwuNX+xRKhcNHA/k7SDygoedDE5FyFx/d
FooO5Q7GMOzmr1fXGqtXV3ehCTe1bc69FySSXWa2Mzajv/3jqlFEI7867BJPnC9+
ptGoBpbWijOP96TBpwXp5N+k7a3PULx+OkNQW+mUkVI8yvHZIG5pUJg59lQI5hQR
e6ayQo09DHO1moxaTbv/ovInYF7MqLzjhKQwMAiJ75rZ1JbD6y51SUwfNlL6ExWn
f5MLtyXTOV+ehqNoIODY6iDWNFoHzATAAJgRhbPHIo+HDDKml6d1ePmc6hNVHD4Q
Wx/N4ZxHCX7ngtNscQyPvcC1B/dW7h+0GulziIKRQmCH1J7aL1eWDgITF7chvCsL
P4K6jpCYQbFh5OZ5o15jUs+VyQyqcV2T8L54oBrqoiVcxlsauU/MhpUb3OvbUCUK
8o8cTgWXtdPX8/mKx3tT8MVp7u47ydizicltPKrx3MNj4vi2VUaD0xeCU8wQqjoY
op2qaHAdo+PtGSrc5QkmTFRmbGGrwba7yuvbBCfuU3NBYZmVjCpHv0YFfT9CN3oj
deGjBUW2/AVAmRURo+QWArIWy2nYSiYfcK0gHLgqsOgC2K66P5rjX0b+9LcFyTsm
R7EDaWVSRSZd2zbI5N4RRzeHchzBX4k6fUsGTKUECJUaVwZ6Q+R7gmD1SArnnz6u
KmVg0brIUrgfnepD8WQblKVmAyV6Q4On/DN3nI1X/3eDfGKKtyGJuxDL6xFiJfe5
kLHwawHtqXUh8HP+xSj8KUmUlBAps3fmNwccyiMqS1k5uc03gDcuPie5WYSBpB4p
FIEmF1hucD5a7mQVukFqSQGIyTjgpxDpdWMhPdtyLX13Pqbt4o4QGJ2FPCQZZsFR
349f9IapeynMR0M1SxOhNAXn+IsuLKCOs6Drd3qXeQAZb4+0qescMqFxn7dSoL3p
zH5ZtaZ4bP1l3qxn3l7FGeQcHR2SK7ySm3/nKo8hrzl0Ih/AjlwEt3GnoO86G2Np
XWSsz0k/s29E00j0b66/Ze2D3Anc3hccaWmwGNmGgJD6E6pOhjJYHnpmRPhoz+JX
7k/Y9Mf712tQAsbQ428kSb2KzBM5QDEhB3S89TC805zGrVEH1EujydYoU6U+C0N/
X80fE12HpPXIJ0WM8p4lLsNeHj/prdgGGbPp2mCOpk7L+ZejkWZnHYmF5GWbUOfd
hkbpp66SqLrs6WlXVtS28gy/3osYKl7ZEonZq3AzlLEZ4fFAZhswIb68uZ+LdO//
SxqCFryFzRtTeysdA0gxYM0MlxWEJccV69KV+HLIapuPKlZ9HP8RIYO8FuzkdZmJ
PQ8DEEul8/ghQ144aRwOyJaOZKDYhKnzmRNs5G654m4mtZHpwrt1+23FAUc37xHm
DhAKHEy7dBOMaHKJKRuwkgmS4ld5rxYd1QM+0zFpkt/onn681zdgZPPK4X4OcEu7
JX6KshLzpWTKVpbT9ewg6vCYL+BqGTFFpD+Ja7HVDIUTj2ZnhCfBIAyzALsm5Y6s
BJkUJ5ON/7+bWM725B2XsrzJnfAwE6bfW2LmBGFYxaQGk+13AH5eWCEStNi2FOyi
E6ZTBJUfxfhV6GC2RAa+9MkfPhzoQVTqg3965zR5/JG0aDoAlY0q3yKFirUeJCNI
BffeFDpc+VuX5UMhS60RlYx+RPDJgxVsWlGLgJC9AkOFXM6TPDMZXC4Xf5RLDlEt
ysrXcze2Wl2t2Ydctk1pRu3EGjlAv8Dg/Wnxx4uBczp/hXHprO9slgAuJuwRVOy7
t3hiVY6dkaxwDISIuQpV2GqsAOLMTm6qi341WFvIeY+wufW4KfDiwuNfrv0SZWr2
gK1/cYzZGam0iczfK41N0hVbAQP5h5yFiQQpWsxSSPgmWU+n7NE8QTUBOYzfc0lT
kcSfU2tOIt44au58aN7UdeynluvAlRDNUSqcIetiljebRKToGhv/Ml+jfOaM3GpW
vT3Ht/wCy1xrDPW66LZFMga03yRo9C8//KkN7xrgdUFY+U8vdEiyc9ZvXxZk0OnK
z3kdfHR1BFyYAF94+xmZ6mu+vKNOaj1dYKOB+qWdvY5xYLrSZ/br3fFvBRr88Q3l
tDmtaTktlCtNtwKPMUSdWkxxmc2W+jz71VThTXTsu3SPPdvTnXBjjSTvNZkLbWg1
NtShZFXirWthoUvSQ8YDK/mA8+j9P5+r69myiiOa+ecPVx4aBtYMBrPn8xGgYIp7
MUwySfAd4VpXR37Tt9c87yKltPrHrXEGxyHcsKPMIpau6Fu3ti/qagLY1wMgm6Kt
E6Mme7z19fmF363eWfFgku0JSxyujcweYFb/dl/0rxXDBhvEFGip+ss91Gdy7lpU
nAi8iRCLjM3KXbhCfvr+EuEBKslt3Dszyn4d3fXEsMmaZweZr1VkQJ+ZHqppkG7y
NHj7pj7bBcpT67NkhwT4WI0vpFvT163OgDjSqVVZ1r8Mf9VRXGoyjRB09NWxw/pv
wqPE4IMN2dt0XZpefk8FGW1nVmvLazeRZH4wZTit1oN9SagVARhvDdf6gEsh2dx+
zG1FuuCH+Es7hA8D+d19Ls1HPn/GvaY1iBkMnTXuKIBvaTGND8avg1eDrLY81C4p
8yk/7Vik0davaVotx8fg476HDKtxXLtUb25o7Fr3VeRXlvCX0InT37pgutzT2oGn
Q3WTJABS9DnDCgrEJnS9YDwW29cFPxYmFpcjyLd1l3GD8vR3Ew1kKYAZQV/p/ATB
47GobUZRq15yHwF6DngA5pKFYy4SaVbjU16v82p1f+cB1jdf9OSRIm+bM6L/3otD
cADKr0/5a9RS3XhzMNDkN4AOwBp3ukzVY1ESLI+w1Prv/va8WkhYlWsGHF5tadtW
RBRTROnQFfEJe36z8IF4h4uWCUxdBToKhE0pBCNEw8q/DnBIKolBnerS+YF4mgNM
s1sLo8EL0BCiZVottSBkiI4fEA3epbwXTQjvwr5MEEo/OWz76HI2GR1KVUqE1xWs
Q7MFrbWvDkYNHS+d2EXB3Uos1nVuEP5jZjVa05k4o0ax+fEdPdjIDHh64se/N7E8
96Lv/U4YcgxknkBvpVHxvn8rKMJ+kbq2n0R52/UNbGwIn9wihTzLp+8n/7G4Zb6C
AmTMvfKca+k/0v68SNEsOSaGPWMRCZTY7ME7ihJmeroeq+JLgd/XRj5xbWKySy0C
cqvNhKSgqOOImZUrQ1aGNqyDVn3+TkLI67Nq+ObEf+16nWuE4anV3XrBb4VqY/io
ttfDAIN20rYRIp8DGNkwlp84RcyHfC2a6VqAzqK9TNgM89tUkR299Llk+mhXHb9R
84/M+Ig2jFC7MNX0rddi1xJjDPM9oPB76r/hmR/zdTMgNeotK6C5UwbB1vSN9xJ4
SQq99ZhAaXeMakBm9MkDcgCSlSvsg5k2UG8Y1Rdz66TSX/0zLi/i1BBXvQvED6iM
9MxvDoYTh5X89WoIzBE7z8JUGgJ2hg+iNC3FnRS8qwCBUajpzskAGmthJjZFAaFh
RePz1UoPZ82XKvArI8C9xAEKoz0ol0Op74De2gCOyj0/LiWj0HRarpC7NLKUqQDo
+vcgOGOnuA7DcO0PihRtzkZg26F2MugwUJ5+Q6E4087lqq05Exkep2FAA4A4XDfi
9GRU1FY8Nl+RkUi4R3ukt24We4eaDDBNQI7pj6HmRwE3ACzKPeMIUT8VvEfrFoev
rrX2VoV5cbz5gYL8uNZmYNhT2xDY5SWua/q6GhPLVzPBGqmB0G4Ih5tgngJ4u1P6
RkRO133+y84pHJekHAzXRHprVp61eqxN2YrSonSWNFCZx7OqpIWC0B5im1eM4D4b
4uG14zLwLMeJUl3QtDQdRHTgg3MTzhimmJ7apPc6i1CxHuKTFDax0nDuouMrM3St
DW4isFxyAAnsbrXo1kXL/34E53K0FUWL2uHs/d14fO9LKtDD8nreW8Lwp0W8zRKH
RgatR28W/t4iPC+lY2qfLqmUs8eyUV2RKO0+eG/azPXok8dU1bgh3ScYkRdBgefB
PKBC34HEeelqn86uL3nwLcxbU1G/fGR+ZPBdfwQL52LaatztSJJ84p51VPA9DVD5
LgMxQB52ys0r1iHUdTuXfhUnohwVeZ+ORDyJHZO0F2ariLjdXF7krY7l35CzSSGz
NLaWNsHySu1QwGUzSpcBHo90wpcfAvzG4Iem+oXlwLI5J4TQrZRkYapegDluIhzP
jq5pW6RQwEltixtr9qFa2CA1bdSySuolIGhb6dDSiyvTGewP1HwIjo3x7Gzh3PSf
ir6pbvOGny/mAguLgxEGYOvtl4hGXPY4l+Ca4Bb8RF9FnhFrFug7EM9LSENBJbJz
ABBc6dNbSVwyfhExCI1cBBJU1Ym7jqeCc85VEHASXaK8no51hWVxkdEwDkVvE/1m
jAcja2wYUyLBBWch7Ya9jh8fQlN0PN5mHK66XAPmYwhjDYlQYZ3puI+LTWKNnJg6
azCPc7yDnS+vJHSVaOCs6dOaFbQ71pVvqeCFcY6sJWt3ToTqf5+5RrIKh5n2YY/a
XyM93tXi1VRoj/s8DVIRtZIihmUmUD5Gd7SuZPJb0BHT0CXPKzmn7vxlburMGMyw
y2Mg+GM54WDz2cmTH037bBEIzruJzeLzHY6d99i+aSA6C4uxyJLPE4K7GDa5Nkms
YAGesBR2LsCQhy3iGXyarMg6x/IH2/zIXpkKrugIfW9YexBqeq2ka/YbT0RYZM4Q
gQG8MEwfmqsF4vYNRgHwmcRJUod2myqkFUNNf3KwAxqil9v8PGKqpOR5bz/XssRg
mXILRO3ZlI5BMiD3x+KYlcZrFJElbXJNFoDRHRh3k7QBiR2XcxTkqpWYfWjxpI1q
zgwVakjbXiW9IqLlUISP3FGQBqDmnbzvuUn0a60gie4Tf5Q5ZbGly9uitlh2daRl
Q8SUKnreMz2vkya6+7DdRCKaS0Zcw6t+Nzl2ZDcT2h9lPNnLheJpYauQbyXpBBLH
0QqupZv8eszQQ1VRKlW3OqSVHyHVVQZlrgevFEcBJUtV4xSi4wt2QsM+kt7ArIi7
N8G8kIuIxu2zUWYY0C83lzf+gMRawWONaj1+xFbwqIBltr+4gUVoNOgmVqHmQYRc
0m/9SlzLYVMME50vwkd1QZKy0kSpBBN6Y9kWBMSKMH1iHvuuZrxBQPf9fMFHZ+8j
QoqoLXEsydtVMCJkuDQFA7nCaEF5OJFgp/hW/7DgIIaRfS3XyKycemnwubxM6o7e
hagdy5hlkXyG7f3wJVEzIhdi9gfK5Zx3GWasj8n2fnx2vNsbvJUohI6kdSereogN
tj+oEIAzm8TMmsJIl80ZoJMek/MtIMZlYRNwEYbmSm0VjbFb/iFEPy3DU2W/e/Vp
yEY80dUI1K62vTGUBy5LzZh1vZF9aGtRDpYa9Lc7feT3JrE0ZBdfTg4QMgjIJB4G
keSOUNDxL9cTaJcQmgAVtz9K6gPCTSojr4t5Ylcj39C4NNUKUpB2RGWyyHmY7Nnb
hkekEA1+9buSJY9xfyji+OSVSmQs2p3erfQ7umkA+GFtmG41ANYjyQr7ER6jJyVb
qNl0VgBJZ1YDM0P1lOT0wQRYV44zW6BVXiZgC3N7AuQHaEThTyx5W9VlFqXvN3Jr
juc14yxJEueWNVQTd0c47GYJjOB5eeao3pCHVOQx3SFX5lEBHZKCjGFj4BHahul6
gNWY1laRhqhVQcJ1r8C6oEip+uviM56h6ltE+LrII4K/2cgLg1HXtd08/sgnqoOt
DSHIjyhGUdAjSkWfHOvNNTDWCrzpnU27awwB09wJ6W0y4KHii2TiAiyd2I8ezBZt
RVTG/tch4KDcSYBTsGvmaEOfQahIYI1mnNqXhEJoSdjiHkIoNMeNNxWGY/Ww/fdw
OAYLg9dXBDMvrodNxc0dT1SXXMMAbgOAeUUOhWxIt5cM6+L0st/VxkSehJqSwbXX
Rl2I/198wNZILvhjlVZnEa9+CxMtA313JKCDpy3Jaa3UF9D/4KwV0nnJtVfQ3Pf/
uPLj+ondABvq3AxFBY1sxTuGMwGiyjRINsgppIN2LMrLDxQERMOpX/qiFzpy2naX
2b7zS+LWsPY1y0Kp28F+c9VBYqUUHtFScadanm1ltOP+UfvEBZk1VNxm5Vzt9jGB
yusWSZbc469AdyKHXDPBkS21wqmGyFfpfU/9dLyxGenhewE+5GcEgkSRsWs5ukdO
EyH46qof0eezF9uYEI+QGptxNwB9qY/r+8kTL0IhlsTvuFyqQqI2BDPZBV+5BEL/
wbpBBK0fAUjMYfJewKrDzq7G8GdpTsAe0ob5Coxlb8gX4XbI0jVsK2HutbeeuhrN
TkabrBOqAMLGng7FXJCpKhYtcOvZBxfcneuA3FenvNpgV20sH89yINYxlEC+NaIQ
WV04yG7fiJ3M42y58PSbfqUWgqutPCnKTkhPiHjw44Rd1Zj30VGG3rQDJYV0sbr8
va/mFzu9llTGwSQo2uV+8cI+cjcsrknaun2uA3MzcQoDJ1LyBQwToT5qePsEmPQg
9FUb9u8jKMPDqGznqid0TH+r5YhaYOgryF7qp/T4mGDiXmquMC4P1zobPuR/S/ho
buch0vMgKc1Et93RdaPdE53NDcvN+ZS1aWFvr6sVnaHVLIiZs557nADb9aIgaFs6
Ea1eqGBUdK64VfYb4JS4AJXz9/84rfEqyHKmNG5g/Zk8H50ndhe4WmknUyecKfgX
zIfu0gwnlC6uxC/Al4zeE6VpO5oCVMWmbsuB0eL550ni4mOf1wWvL9XoNbrBluQp
rbtG8OkDO0IBsmclo5GhDgIlFlx6wrKE5y+GJbrLLDIiOVoRCR2jw6fzQqeDsEZE
LfWpFdn3NSA1362ajYY9NPvUN3vxhVXHzpkEokYE6bfkVHy3HYhweJizA3b6wqGR
/nZZhkpScw1hJLFJsIbeaNkWv2DqVBO0yyxaFLLgxFADIXjhbBL6eNwpchza2APm
zzyDWObua0s+sf5qqR3jt9E/yTcbEvhROu11vtsGSJzXCNzx4a0xk29gpy55JRLX
7mHfpdU28ovq4L4orh7wG2utxw5MdisBsfdfoz0Pqkv8Px0gqzLAUla17K19Ffir
P0gbpQWGQgM51+TXTAAReej79x8xTt1UfBjQgMN7NdWMBT3OVDDEChTlHsAne+GI
dVPSg4BuERDDtMNH2NllhB5EuJT+DTAhXfqvaQxgbIJS4Xa0RaBW6UIZG0I2Oman
+jlgUmKN+fLM+S4GEwq3lB34SzTLiR1ToCfafc7H230MGqS1J67rLSWSEa6oIL5m
2o1sb/zLn2x77tOg8riTt5/5Kr/9HPNqk+pgJ1u6Z2uhTr2WvWqwRXm65HtDNVM9
mkjRcq3QcU9HAu63j832c2o5TNQ6ogDjOX8WXChvpHe5pwHwFQTXZCxuQcPHbWFp
0VxeKe2o8HFXLOVTkecB/3ASIMqCSfJkJCnT/yhrpcQemn8mxjPiJ/vJ6ltb3WMX
qGvZwH5dqZnPTad1Mx6OP3pJ66Pux9z2634gm11+t0N9sI9ziGJ+1AtWsG0RYJzM
MiVcgG3UhbO12fM8Btg+f2FSalcE07Gchy4DRV+D7+cfKcc8fhs5IoPSbKEvxWhd
kpzjvDYAqMtE6MZPu7u6aIpIrjwI5boDwdtuZ81ACYbKszKc/g1F2+VvQ8g2KBSA
/77TamatTP0oq/Ugpnii38hF/vObZ7AFeu21gaSXoJTe7yWXH0Bt0qnzaoXEYCRC
N9/dnD+yJiOU8jBNoYZ2f5ozo+YWThFfiQ/Qsxgxz6NovgnYFNRqwAVNQC7k0vSa
04ceFMofgeLOIq7BHQ79kZhv3rQZMTD8i5x5xCIgpEwbJAeqGdnmTFIw8meCpfHJ
qOxxpEYQYBBwYxhzEC5tBwOqq8BmSpgnGTfP8vNuoBDfxZ/URyla/NFKSEHuDqAk
T2WTkB9W8Fzcn10WpmKTHKLDnxGkzN2BZtmXz7Msf/kSnjc4k4A9mRhCFgeBWdeQ
lBdN0u2EA6cxBr9adgAWnkgaGQfABzlGcffwPkIuojSDc9UK1Nxmrjxz374mes+Y
IOckbM0FWqsprzyG/+E/Q0RsRCinYWHKriR4jNebVfLbPKVeGqDbatkozDRO6ZTS
5Ev3K3QllozZSfjfKMMQLBXzZcMhfM5jl17/y+XnH6ZC+1m9PX2gP2vk1P9aCtGW
raFfRvRsWRDsFoyPrWVr7+8kYCNtjcYZWvs/IUiuIgosmFnM5X0Yj7m2vb8dbPbs
CJr9qzJNXUA0YrBPPdLp1glzIrajQg8mitziHWIz0EjV6UVlKql0tOqd0yqx7XsL
1TrWG6IOuBSTiAlM4aKAVP7VFn57beETqNUTe163AfBSB5fGKECYyc67FcDvqkHT
bkZ4a2f/TDrQcZWrVLWW+202055vAyTu3qmF575LphOjHDS7ahBJqJjiyvRrMsUi
Kw9gXKssuXigdt66+0kzDdY91j3RfweblCpo3ynJcsPbI8RSJchaR68SW2QT5hHN
+LvUKFV82zdhkI39GM2tBc+w0gskljgkami0VQ4L72SUQPVtC6Ch72kHS3samb2d
DsOUCY9k62xdn5WDc3CDQPTQmdBD/gR835/bjp8KF4HWYB28TWm1wp+6w9FuuHwW
CEuhip+hE8rXjjt0lDeXDFBgvaem8JM6JKrXKmCBBAaN70xgRjG6Is4vYJIspCXq
glub1GwyjotR6+SLzSqGHnXCPURdMKcdKviDzy4KFbgW48geRH9+vyXiRBvi6rb8
qO4rIocJW5KA98C8nHcimdJrB5+0+CBgSbdT5UboyBlfSqYxKw4OyPSjYsbVDGpx
ObQXVbMi+8REPQN8Sj1H/NA27jIRXcvH5KwoJCLLM2XazrReknDG6xp5vfMSmyOo
uIhqMRhAK4Hr4SUplRc0OA/T/6iR+IWV446HN6f1NMhfyV3bHJvS0GxIZqycIBdi
OQkNuJq28s6/Is6N7lCiigYgNhTU87vjjoAG60kcKOX91osQNRD7iQxSfiKoq5Rk
bVE/SNDHx7UH4TX15Wu9GEAwpVgD8//clW0HTi2jDi2tT0X2UybrIAgIcN0tC/1p
c85M3XjN96ijXUCmkbgVOOkOwlcof9VgDnxPRG0jmSmILpuPJ0SmMIKsYYFpCDla
Gh1bnt/VJX1K14oDSs5jmVqRy6RHbM7LKaihe+0DNJKg3Eo4PEhg5xjcBpkysRXE
kaFD6qpPXRO2gzQhNf3E2aslLtLoDkumPammT/c9lkKqlwXJXtyYafK0HtQLx/Tx
CK/77WGmywkaegm0GrVfmwK/FkNoIElvc1oV47kxfCQSbluRoT1LMPdnH3sCQLwi
ktRujyFSUa+MhO22mO1QVni4LA74lZ2KXz8jQ7oSVTQ1n2FGaxxxWuC6k+vYHxAR
TpyqpQxJx5vkk+uT7z0TjDskXV6ntPYCMfcCOATnSbE2UMHkABmjBGenwUeLE3iJ
VyfRWRSowu5o0vOuZJFJ0Bt94Piagoa+Xwu0DN05zToGnhXQBOIL1H/G/Pitw+fa
AHGd39xP+ss4TsXkfzTsljlALCLp41Cud29dBKB3zN2iCPWO/Efmo8Y+D05XX4VX
rYHP7zcsSnGEWwaucGJOEdZmQilU01KznKlEx7Hgd/vTBSVAPLGMIPQxCRpKqF2Q
Y2Da+Vvyd62zAJ/rzrkL86/jqD0SUrtivkHDX8maqB8bhGYHYIqgvjBvG14SZxEv
VVy1q9bsmY2BYkosOz2D2jz4at5RZ09t2kcqvr5ctNXuIAm+JSfG7W6R1fCnT4bi
I1TY13V7aSkSPZL6N+Qp5ocyj5HL2hICBX2m4fQDPeeUyVkLMRONGapXZ8SshSpj
IRjx///xf5EmpJp5rBme+Pakq1wqTosRqiwEGFK+ks/XGPbj6SuYIRv/bZxp5sKw
utPb61wT4RtE7wiOlpnwaf/FKlevWGKxxGbYANmXANVgRa5woSlVDw+mtUStsnm6
m1Dg6np9C9qZHoI5wJjH3sQT1W7Jb4teXZPYVYtV5pKQhNdJUviaWHsW85NOYjBS
QF1wcpyMTMatA6YqWmbU5AJGHhVJchAWzRyqcLBcio7pNw/xyBlQOHymOThlLhXD
uKY5zUy/cPNEEvXWZxyVpGWsUeH9bh6iCH9BmM6t6gJM1fyAUJ0+JE+SuGNniIYD
+HeN9ASB+DG1Mdg6OkEH3D2HGCqUfSKYmJHGvLooGlXCa1HvXl84YmhEHFCHoZS/
acYlU4EAUz8iYR9xjTedPofADwzc7ZJtWiNmTYQazDmL1elBlEraGp1vSUEEfbmZ
/Yrp355I+gm846uS6koXGEMjU6zAtc1zjw+vMeSYkgknx3OuZSj9fnZf0uNnpghJ
8TUSmghqZxKLuaterZZGNfEkFI8wTwlIGiFNB6XGuj8xA6b6uLoc7AbeRR4i3wFK
KVXMrrLKgUBELfe/dBIxzVWHHxQ7adB+NBIlylbAW0LSXXzZeglLRW9qroAVhcbT
y3AoZn3Ly6QIDLuBjjSE2wqjd0fNC1M47Zj8KCWvcWm3RpPVg0w7+tF9x4GTTwSS
AbjanFsJXb8s/2ePIBdD9bROaMhU+sJlXWP0pFtaJ2ol7PIFi2JYTSpB5tSTOYEi
4ZJDQzG1bhLvoAjYPN304DhjWClqw5KR4RzSmIP/3afzIXjPQa4t4Q0VfpU4GfvZ
4sGxNR47BwvpicyMGrWzMwUCXcUf/9PGNHBsrfX4Pf5mDa9C1ZVqtrxsCTe7GrHt
GL9u1gqUXg1BUXi5/0fgpTL78jWik4ZFsMkaKF1oTpxHOtMHOFR7jZvkU1dg4Qyg
8R2p/zM+n5w/7nnWCPD9Mjg1Svl0aJ+VgshlntqKYHPAHLFA0xzU/2bnLNjmQkZP
o95syWfkuOKN78bZcmD6Sb3UyOpxwjC0b2J/4zxOVr4bzXeIX8v+2hkZK5UoTJHf
0nf1H7+Jh036Y4ATgmYiveAuYfcGwoN3B9ILKzIbjHNO5fJykbU99yfXeXIO2jhW
gpqoBxxOg3FrSuANpfwxgJTupF9G5QLdTiiscwBJwy8+8LQ9vCTYhWNlvzp6xAew
vt8KG82dpD9lzu8spDqAy5LXgOEuiBDyuLPlJ5Ya10KDQauKFTk1y98IJwuVYwTJ
/3BVaaVgeC5hS5pkxmEp3VHvzeWwOFIqvoFEIPtOqi9mfTKKehlvj7IiT5QjDktM
mcMcpgKIos7AUiAWZEx/bQVWFyiFQ5Qfg4N/wLzowTFuzdoLjMcG3dTQjksYpNbr
E4LKoHUOYKWXgcHF9EbYECkGBUd3nSYMPYYQ0jBUUFfkp9iIHkg9Q+NMhFVEITno
46NDpVIQSduLWn9KMBPidIbeKLUamvRR2nJTRhIF2gZwhTM3o7RvHLMJG4j/eeH/
Kqgkio2hacLXH8QmEDhg3AeMH+xwPKDZcCzEFj5QmNthZASTM/VfNAGpkSEj8UB8
SvXE7Vqgo/gcVU+N+VdGaRQEgds0TPuSXB0XCx0mX4jz0QwJPaHKHX1ZS/ij8Q+j
nNYDie+CQuJXic3LbbTU54ZK0bjqUumj5JC2A2g8aS0r4UxV0JlXcoMFClFqT1sU
ZyOLgSAqftwTxq9CWKIcU7+APX7nuolWoGbcKOZpy5BfPtcqbnWTSXQIRvPbd69l
YozK5lqq0bZz/rkkt1lgNTZ58+riDC6h+towRkCDvYkjf3l3ltmSo2OL3ZQ0GG70
ebZ4WNvk3fRgZ9fYEOS+8rydh1+3tTF4RzOmbxCGsjB+F0vv0rr/++ZgFSs9rGgN
S5AY3V2fvylUcxcwKbYbrg9B0GNNceSW9q/sxlyTfgYeDy0l49ApDMuyjQ6vvgQf
dOZJx1y9OaAdZfPVkoFHWxaQPXhFpw2571v0mWAqHXqQBi+TwfuqAEx7ue0aJyju
UBf5lafflFVgbNZUAttu04soTT1WpiUXJBKQLCffcMnQaI1ElR1KAS1rhhwlhNB8
M7Rc36fQMdievbw8yMN6Ik5OP0G6uYIffHfOTj1DqNvCx6SdrGXpku5q1lFaLX+K
VJTakN+Xojljefq8kX2o5dWEZp2m59CedcvK6geoQEzzPAX3HVVechdbVU9+eItJ
Ezc+7jvShOtin3+Normfv8UrVKfhURJE/1YPt2GAkd9fDHBtfr/e3p4w5rgcQKLJ
VKVKvb6H4d8sgFDTn7Y7joieqms9qFgRM5jhCyyR4I37wl+w9yNkulTf5FNFDChy
o4FnU2gGG0eynxOOT0jEcsTGFfIw92nWiSGhTE5enrSEy+pJn3Bh3kROF7fjk8TG
eI2Fht5qJelFgZ9ZLAvvUZlDPSw/CtUbHPkWPWz/9h46rDGVUWy3Pxl4tYb1jfyf
yca0Dal1GB9SOaVT3pRmtpXl8QdtNJUK6R3wZ36GgikFFuEmw4kHcNXLMkvH/x+x
3hTUUiqikO7L0t5gkuTVhou7I7MtNSo6prMegRnwyH7gMtJV8WoVlqTYcKLUMBTy
ncEuE4rmxmJKFF43bDvJbmd0lwx82tDBiSY0hmN1k4Jp35Hwnau8YJHRqNL8vpit
Kf5EQLcu0WMekxTLtbJ+5ya8iGXx57TvcxUAz17d7DbEEmDZscFvjd/45COGB4Hv
y/TdRUkRhnm3jG1HLU+HtHmkYxJdnhNOeN64E84ZrBTkvLsK/7sf2ejM7wHwWJ1i
GM7cQSnw5BLUFROlcoORlKhLrmwFACrwjsNDC0XdJTqEtvWKe5EQQ8winBmVRLZd
GaAoMYI6zuQjB4+p4/lTaJdN2EgaSKmcdaHTfrA8bFa2ri0MO+t+IXC3jiIHHzt0
t65TJ5i4Nr+jvSoWZx9vbwPEAfsvlWRRF37mpzE2vJP06bhPn0gfrHEsAjt21/7Z
2I6M6NcOUgzzQQ23kErr+or3kPoeM87mVM6fRN1JlXDHmko2YoFXuZSGM73xBFaK
0428hVBZRHjO/ehFqPYB8C7GWtZh+6iliUVFS8NQ8HNloGmtjg5iFc8TkGu/GwdJ
8AsISe0Tvzbulhs4GEuwdom2WeVSMYCJ1KH9XezlpnoOgnLJBaYMjeQqTGZue4zu
8FtMSZKBhrGgcmMQ7LOirmHBS5YvtgqRLQo0mmIUrks+RJb3FE9KxK684U4YujpN
6dfW0hbzvFZLgxK3jtvE6cNhL4qJLZxSt7V15K90650HeeOtL1rePBLzksOyBJQt
vp0NuN6ZV27hiTZaey9EET7JyMs3VeRmSA3wr1CW4OCEIAK9NkhQiK72YuQYB0TL
6WYkiF8y2RodF7bOUDCjokyfz1nxewLlNcNJmilUq2Dm5AsvbAOeJhbCvj26ouGe
vo5dsHdjatIS7T1kgqYrRYBNB4K6ehH1uqOB7tArP45ZkMcB9VpskIOCsXQqgT7k
O8vO/f3rCz0ysHpeyvxgzIfEY7VrwsuhRB0i3hbDkOL6IJFkUlojU5jIg7NN41tB
iGOBMw4BlwEnO7KfS2QUiDjgg41BeP7QaOclclPH7IByfNfcjW2mjALRSg5mcJSA
KV4rf0sC0aIoZFURPXmfK6/g7AxE7IHSt26x7gi3NwlqFWwmgI77vWOIfrTwziM2
LW8enZFH5lz0VyyNn4hXXsAV2hBT+W1T/q2ci174m40kbliKDcTqRINt4Hhb/WAj
3YOErlpNz7toOsCdVPuI/faa0WMgzb+tc+QXZBG6JuUYAIcK0fUfN5mwU8ni9xyw
c6K5VhiN63NGUqn8rzEwHyMwu7fvZjIH9xgjRwVIf4sHjZ7IvU0Sj2mXhj2qPGpH
Kz6H8khdFugdL+bLoQsU4Hq66B9XH8dSiyABNmrwLszZ09sUEgjEjBbwQvZ/ooEj
DWxCiaMDy1kypDi5mceiCG8EOHNESYsucQ9W0Gc1O5VInmzwgGJgIBlZWxY8PkOL
Py1FqEiI/isr3ULce+YvOp4BH0jX8tmL7ECVLF8ZN5T0NUNJzeXSqG+iWTHi9FSd
C5cukzk8uM5K+f9Tj24wtrSMIFdEJwoBwjv+TbWUgtazDOrDRgSHnWgWwDcVTs7K
gV4A0FmWaq85warjOlPnPz3mKWUbGPQX46gCQj9IjxTyWznuTlvfNoiSRhQ2LR+j
EopAzKDFrYViyu1wTzhG09krQ8bUK9W+nfZbMjv1OHt4Xbps5c6ds4ZpKj+bGyvI
UXbWWrcXiSayOo2/xWSNyNW1J8VreWLxqn0flloK8jjYw3jXd4J5k1WCvnfKWC8R
NeCUeT1BxZ4hlE+547V5v4MMn390bpAU0Z77SHciaMU082Cr4/XA8SIF3zmLOVdn
ppYSO/3ntdZGU9vyfvMud711Jvl1r14HjVrl85zlsrR7QbgkGhf9xbjaniC8EtCj
8bNkM6vLD6IWAOu9lLYoTGuacFxlU3lcUS52QZAVpdQug2nCqwrQp2pCZn/qKWMw
bAb4z28Yuh747SBgejSJiPtxoI6wyvHfwUKSm+dSNleaY6WBrRz1Cr+LAQVg1JeU
WSIA3wiBp+22Kiq2TR+keho9yQhFvIQpTRnC4tWZzkf7Hlai2lcSVzBVZwa7tc5K
Hj+tGUGaY+A0mSbCMJpDj7CBjkG3zA1xAZuzWUeeANndZo9fPJMzHcMLS/EZs/b3
Ymongzk0gFSeMNuBR6+cQJWtUSvfuQBWb3k4cBWx0hiPdOUebsFpH+ey1pMZM64h
fsccVqfAmzQ8QmBpoT16yjBefVVyTlK1Nio7Sa8LFWHfVBfkDnJz/CQPJ4EMYNDe
x2NaJZsFzdLoSjXPuXYxG6xzJRzS4aHfXx3pZQNad8dLzR6l3BBD5Mp+/xaz3SxM
DTUpJcXssKMEAzmzytpAHqCmACXPS5+C09bobCcNfdkEDrAbisyg7Xsyek4p/C/E
72epNldTSRQ0vc5qAfSwtH+j8UiDwskG/QDUeZuGdPPhJ7Rjo/KolDOd2oIjWNAv
NUSmJKP7Ccy459mXTD7tAEJ14t51ReYKStJ4AHTJ+IHPAzkAoyAOjkYDgqRPWDnX
mDDxppqOFo2WNGlFAuH7YoNyKNpkb4vmW/KTyU5RemtnWy2y/gc7bUNJWoC2pD0C
QUjvj7+9HsfGqyQuGHNeURud6TdkczCT2oNyY4Y7C74lIgDcFvbo69062gKAm/Fk
gqc1H0fXngAcRIpcqSwokMoG7cGYGnzf6VSp8YYDKmhUC1J1t+N/8j9umrxrFMaM
Wnkv2xOrHsA29WmeFGdOwAydsyaDon/md1p4dQmm+sTdgNh6HsMADoBBnZfF4mug
dw4K8PHxmYO6FkLZBnMb19S9+nxVFT2xEgbh/ATLWH/6E1DBN3ZZzO9UMQm6Hak5
sh20hTGhTqGK3eBdjSaWv1aTvguOEiMy12/TigBQLz+smNEpn6rXy80tEg6Gcvka
5S+Zh0bU8e2/RIUmIKBbtsBqqLWcPIl+SZESaqaWgZu69IZhVb1FALF0VEZzs19o
xtjiKQaCwMN7JT17PJ6EB1ge3PFVQgI/oDRlpTAcwNNNvNcG+BuA4Cokq8RHdM0o
Wk5OhD4mH+k+NBfbLrll/1+oOMin+uUQiDXnLwDja93nUldk8vV/QD725ZUWCzvj
raiKWzel/YUBqrqSU/3OS6MgPiOqbjuMmu2Gya9EtIeP4xDqWNY6i9QouJb2j8uI
ajb1SwGCpYsPCRjWhO9MnwRqWDmgnLnjOCsxRXRjPgOSaNENMCfzXoaGyg70ui7C
hxWi2LVmPe2gMOVW3K2MIiIyD/wqWhBCaaXPXONg/g8H+LLExapi1wOo7iBjFpGp
7s/tpcfwWyR0sY6BsHPhHNtEDwjx9ZqPIo7D2MLx/nZIvPE29Tis7xv/E5XX7oZS
AQ4qABcgQHherMAXjo/01JCA4DRC2C4LecBsp2/mImRsu/X3J+/kbdsI2CWOr6cd
XvFe5IqZm9OuRINnBFx9yxAOOZ8/G9mE+BFk476ARTTurVVOvw2prjB1dNGVLbcH
bBT0gbLPOm3RDIqvy7B7SViv/g4+AQKyvRN0eaglXvbwT1gUC5j2QvXq3CPVYM7Z
/J+jEvCzhW/JLsGbWCTVRp0h7fmfqeiXF8FMm9ywfffw6HggHLdypFOJ/S4sk/0j
UkSpKn3hLNo4GCAodT1pUHdezepvX/NHifLaD++cYnB+PIVw1U+PkhKkkVsEykCT
Ij+HMIfIphkxj58Hw8Ie9vqd+3VHujOaDXNyL6WndzHUwy5jm8NdAfEzSpmYK1MS
uL88y84gRfeF0zeSv4YsKcINigEVxBJKuUM1Z8eWg64DG4TB7sG7nGXCN/78YKWL
G83DgCS/PahbsSjQpg7CR+8qEVmqSyS8PDGqgvh8B0CPpse6lZh8p4ui548VNSAt
Dne41788P+OGGgV/8RCmc8HY9LRKCK0bUPSB19jQYEbvIRYWbEGKJRB1mAXW3Gm/
R9KquZa0J/F/9II+EMqujIFguUOthZQHkrevQ4xrYxVh42bKJKjBu/EWDteweDVr
hXY54UZoU6wBnxrD0zh9IvWvFzoz6QqCiP3iVG8ij/3Kl0R40t8g2FrK8H24qEfH
9BJta6NPD7LsxAigbx+5rryk3KSf8wHr3As9CXSxRkqZC3SgmZvPVrubXPMqpSN3
hkPlbQ1dKK8yDFy0/6MMhabJ+QPKMgLCkvx/JNUM67fiG4mPbBnc9cNTDgPqJAnv
3g4zR0nx/IroF2lp622oPVwaxalrlW0M+KvbFleJj3NPLH8XH//1IGjlBS8H8nhu
lvc/NVp9M/TtO5Z1YO0AGB29oZo2tdjqannzBArIYYtina+B17WgwD1j9Qp+f4Zs
0xRG2aZi9m1eN0FnA0Gi2KMzjVyD6xxxyKiNmwo3zdMfrcqWvO2Y9aOcvwwCZDZ+
lEcnWGzwbQLfX7cwxxzA9XS/D9LtS24v2xXMSuoCkR3F4rx042HXG4eA1eqrNdxn
z5lXJZqnM7gY1C033Op/ur3NwF98ty9ehJZQq2AbKQ0KiIGuSpoQYPGY0LVB2vPn
vxCiphKmOPAcD2Ke8RV8gEHihIQ1NJFNgVABwKI2N0w3ARTXjh3B/7U3Rkom9nNK
b67qJMnwj5BimnvIIwWVA7F5U8BR2W+DRM46IEYZsqVaxcu6dVIG6MoJLNWsEHHl
XyAJaQU0gF6a4nqpExZUYLu2Amao6UgOSevoH4XmjNVmdKvDh8PllWwweDuVzm18
04WzOWtuC9nAcuCkr//7eOLmEP13X0reluSJyoEqUw2U8Ch37oLSljTGx716uhaH
klKtJieL6J7Aie11gq+/6saQySAchn3CkUmZcgSNjlb7dmjbaWq+8GaeMbkgk7A0
ZFqSJZ7+OG0ka/K5e05HW8gT5xMTnXlgHhFKADscMP4cJEln1jnSK6esOTO2GqkP
fpXzt5DO3+RH0+Yij/3S+u9DOuQwJkllClw4J1E1eJ6mPwTZTDxluuX+YtqVEq1W
5b21Ta0ls+tgpX5CY4sNmZmCUCd4CWJQDlS7qM2wi2tjIa6SD++BjdZlsCDk6Pea
eaPixWB6ZHj1/vQZys52fdaZAsTdIL+alAQ6NZi2PTUVQsGLPLO8wI2wFllj5zYs
i0GBlXNetHNJQcwlPirEzeU2R+dTaZJuecT0eGxIpHiJLbz2TpFJSLnhF1h1Xp+v
A8LXjyLUZLC1t1nSt0/MV3UR9eHRH0EbDYLoRQiGiWHUIS/cgHCzw9ALSodmJfqx
fzVnckSaC17TY420rHbgQP0NVaPWmviA0QEMdkIYPT8UvsRQIXX6IX5lLu7FKx4s
xcPVKikUC0YQzUHG6jvkKfH2Y22FMrqByTxf7Sk1jvii+XnDLJH6OdNqS1bV7GBx
0MYR4RXh7OCm7RlP8ISTr2FHxbKFAedClSZwvQ/YjeqaeCneteRFE2f745Qsu657
yIMrkGRbYoOp3PeufeI48vYSrFxSWBktuNyfjxP8Q0mePqNRqhe5SAiJJVRechp3
eH8GGylu7a6eSgLxnJ7FjXK4T0/hCFCVHa3P/RWh2xwCPzRouJtyJZ1xpt0XmlVR
j/xkZAvUZSrLdaV2HuV1iYzTSNMXLCwXoDvwDTXAFsS/I6Gw3WXrrsT/MG2Q+zJs
Lkj7lXkI2IAGDmRRoViJSebSVQJjnvWc1zbSWW3ZGNw4zvku/yKg1t/kIa822fP3
CyRmqawqdgNuL8eqUdRZuHUCMc39/GRFv5ZK5mw9aZp5EyWbJEUJRCrOKMmL+OtM
KTTKfXOpquPxSscD6sLPmzo+0ymZ+rhpHm2DsaZu3t+U5T5ZbGj72XUAFpkxnIcy
NKBuj1po3w8zi3EBMA+Xbkmn0Ypo5YvM1wRFhYrmeg6T1o/9NOFeVy1cev1gVOnd
UrtVIJbaMzQH8cOJT5GluAZ1ErczcA7j85wAtbwAE4UK70xWxoGMxzVJLIZHRkpy
4yQ2T3V3mvvw0c74cOwHDMI5gSMwpjMOkNzRIZfuhPWZ4CsVZuhppBWLXyyFfF8W
D/D7i5upTZhkHl4keM2f2S+5LIcmf+Z9QxLCMFpP8fSLI3dEX4uGnAosphmO5ftH
QZnaSipLLIPAik5zK8svbCAtL+ZovUuFpJwAVYkVYUnk5j0Sy4xIStQQ2dCUGjQx
MG1/lJG4VoFN9QW0Dk2ngp9yml9FvoKjlZZGf0Hj2XK8fSBjbhJiOhEcKPMCCTih
JMRBJQrbqLCadqirkknr7vTGNTq1OKsofAomkWrzBIhKGhTnpn+aOOywbbWUzie+
2AtRwVPzVulYJlhrpQ6WJdTbkIOT8iJcF9PXOC2owog5PAzDnHBjOp2cumkXac1M
cpVRtgEU88R/rSDEYDoDDqwzqR9gA/YnzJynRodpz03PdlvQjOvI9DtPXnYVNm3B
MIb54UbNFw2wF4pKf2ntS0010AyjhicDyRtnXOMDcdl4N0S2ITkvTzLamJeJmdwD
S5mrvX23WXdNStp9cCe+gXTngJXIa+cYpgrj1B6z6SZNXTe3Kx46ih5SKAWjHc5o
M5T1DbINbqkh6TRe+1gsePLDcEpgsUW0ID8LJPW5LJUazEZtMK0pOz1tyS0VUHN1
QgC+0J4qgdWWmePhNis0AcKh6b8XC8TNEyVtpZQiu0y36UG9D2mePT3x1ADH9s90
5n6beY1wdufgUsyfM9NpSmPnYIoMxYuvnf79H/o9Msabpojnf9sSkKFwBwo/S6gj
IW2PEshNmQTACoeTs7eEOny2miyOrLwsqKh1gn8iK6169TlaxvSrKzOu7WPaQYhQ
R+0/wzM8kGqFE0zG/QpN98kHfCtdSNeQE9XtpMt36Jp2nll3bRufqvzCJJskkvo3
VViCl3TZprzwW6PXiNaY2bB0C0CWwg5gghr6I1ah6/zb4bXamJicNxuXEAvmsDqC
qTD7i8pAGXEc4oZVcJ/K1T8a4hNeR6h4Vln7CpLTqi1VjVwUeQNe0YNkNft0otMg
xyrxrvEXDctUYmqNeieg+OVL/R3GHNcnsbEMnUHkq5UFvfi7/Dy8jAqeveFIUuEa
v3XBa3a016rhTsTjSa0wC2Zmn52bB2dMEbACX76CBOS0BQ5/4i9UHH0t+R+fsHLE
cZ4jLGgVWpz3VJzJXhJ0M6aTOLZ/DycyKbcwP8CJLA5yQGPu57GBPqJGtuh6gF2o
uKabVmCBaEdFbZZcRMQLI6fxbnFnMoVs1hd2cNpraJjbcbABuyNjvX/rsRbpB7XF
GH9Iz7EpKTrteQRW4aCNPxMxAkl57YYAT2WrbN1eVuowEfx893nO3hlwzakbsG9X
lBuCyY+zAzBVfFeagfVmxvqnQSDaYo81M4SyIZfOxD4TGYulcUPjSj06iVBWm0l/
OytUVmmRTWvaGgSp0p1SeUjC1KDjc8UHE0izLnHfJw6JbL1ZU9qGp7Q5jTpf2jk9
YkuqsAmQNSBEFFgGRSHaLIo3rRw6BLhrfxW/w7e18XIwsJboDZu1uovaISJBRepo
TVuI9s8tCvoBMuIqPwKDEAFzGzvOuVHZ9QSmsb7UqYDaJqeQd6G2KhGWI4e44a9L
kV1hNOZ/FuElUooH2T8viBHe9byskuaPQnsy/E5ffENi1IxaPtZv1adrC6xoqbYm
pT/FBMU/oGl9t1aPoKpMQIxpD5Nn0VJhSrkStf7yybBG6BcJ2jJfqROTZq3jpl3y
JU+EnVo9hjm2fpmH16mwGly6alZGEYrALAs/3zJKepCUTUhZ8pG09/KUuBE6/1rY
/7aRcfn+4+YinWW6ZIAB1V2eulGFLH5fc4XLD02TWBSvSJnC2AHjeeLHqknLAcUO
uhOkwp4DuXo3Ih2RDEHTg+pyz2MOcON50Z/D7Q1yOhHmjHqm5G0feYRREVwKYJMw
OhVjZwPo9yOAq0Ktrd/TKex/W3A1Okyhc3hZFmTALs3bwkIwQkKF9AMpBoVoWNC/
wQtGBee6v5tM5qczVokUZlSXwzBY9VpX9zPi9nEC6HfC+jIuqUyReAUzmlKGUdJk
6GKJpt/Sl6eob7S8sRcxSydW8jdBtlehW6EbVR/CGaLFEcB9K4Y99+fXs69FRbaQ
pkaYAoNvsUleS1Lp3GRytDTbOV113utvwf04QeT6DjrlQQCIlQ9hLEJXQC3P6a1b
4GwK1Ah9l9zS2RwT8omn7CR5xcySAJSQD3dq6AMr2U6f4qfQico+6E3f/H5xD7M+
5wmm2jYgoMfc0W8W4O5A1dkzuC7mcJ8E3wuH8KLRaP8CsU8LSge7nxNf7qli0ilo
lHbtyovQQAR0Lc/DnOcAcm3wlsywWHf7WVXyHQhguh/dkLrxt8w+7Te/1oY3qMZV
0YUNKffkF4IQ5CKFvHuxC5cDjUWTpA1rG8Stjkqo1P7/FE14uc5du8kTyQN7kU7C
yvrVGxuZsWsyAHGDyHhQf45SUc5XcNqY6ugCn9zkYbdi7aC4AHNRORG3I2Z+F5J+
l82YPBPqBCYHy8fpeKI+EJMUVniq4ZKti0sEOcqvLJcsPWyziGpil3RPbyoWzcfy
QcVDr3mQyrHuisHMtO26mmpFAM0U0i5ziC8uLBWOEsOmgI3vh/pjKzxSvFp4/2V0
m+4+276vh8MhBNZs+bdeLhGZYNNR5Ce/Pbtw9qP11zgM+SMKuAs2CPmets5TIOGV
A9yIm6PD/XLjeAnCdT2+1sEIwvZMS6khcUIQ2Dl+8daBRxSX3+qFcxaj2ZCL/Ze8
jwe0o8CtaForfTh4JZAXXs+6fNEODVn0lCqqUyjAAvxneb9lhAqJ4xPesw5voLSr
Bcb+oh8g82YNjmnS+8Ma6pOtCUDnNj5qN7jDOZDf8hi3ECroZhtlPCQDCMcc+EBj
QYVkjI57mYzlX2mgvSsAvI1u1bsxnw3wB1E5iYt2X1bBYqgCgaC55EFurOD7v+6+
V8SdUOc0be7z5Lz2wgobgT3LbWPwo8ZC31q1T+HZTSTBo3dohseQ7rs3yeyVHSBb
kYyH5luYch7IoMLhz3cDaRdoaOvbQ/gSmjdW2Ey0sp/+4CWyoyyMe8GG2DfY1wFl
bjFOtWsIzVh67My6OcEaGUIfPHqL++poScVDLjJQx4j8UQC14g8zjjIM0EwzTnOl
BMtIripk5qDZQcNFjjKKyttIcNWJ2HqASYw/MjuRxWYlhSL9YflxFqQ1FVoFkG01
7JBHbLJA9nqbXRURGnSEudlZZOtPRaNOLz+nr2xD2RZtGbK0Jsegn6yK655qIFeK
wvq/q9sn02HBFeTbADVdU+8Maf3qbK/YA3hBBD2fytPzEvRnCFLAeDzVKGbzKtqi
1Cqq3bQQdT8uMc7fUJ7dton51eS6jUQdFcmXFeLz83vdXdu11G9NKG1YNPFdrdFO
2PYSunb8ZOX7JDekkg0CH7wynWA7W0ASQoBHVqIKN2qg2YYPkXsBjXoqA09AQGTb
DRtWMFEi7kKB8g6F1zKj25qOiuslcaYv+iqToJiJ+wls9rJQA5T7IlFd6LMucOJW
IbdBdIe6fYSS2xNxJxpx+DSGLyASH0o49qBenzYxA2CluaWZhPlWRFztkiIp/2um
AKkmiN2Dd4BtUwda6LZ+gXER+HwiSdjenfUvdgc1u+70I67mxzl7XhFJt6BVjOiN
RYetZK/bV67cQK+ios8oepXw9Xjs0JTVRyUrlLnenQ4ufkIDuh1UAaQpQTPcqyrR
qAgrAchWoxMnuY8WBapDjONC2XMfUXFYpLaULyxcCW4zU+NkgVPahqWRkVmu/Log
sdI7lRg9QVzitwF8idaIjs23Zbtbqh1WihsqyxHgoqEoCJFoVxoMmR1+K6pu/ygU
NhQHbG2eedZMgqTNC4pbJg0QABZR3ler0K7mYRywtUaWf71QUXtRdH17iObYI6Bo
7cv1J+7UJhAuRMiXPcrMG7ZOF+umyfShvEYwzSYh47Q4b9BvFUAAFHMgy33EHBy5
Lo0VuEPrAcrPJiMkYV72H5wGseiE/ccxRYpH2u06IfQ1qguc9mjgktgA3QOUEEKE
/Vw2hzhHR2rcfE0TqPkPWNvAlrJr7ZZXTfwUdkSv22uVPBpjaCTJv3AQkfmsIX5f
RGa7s8Gcr9lPzUKVLOeKs+8RLWJrQY7jNsFuunkxJmkLq/f5d+VFBBDH98YJqmCS
N+l8Z4n0fx1+Wx70hH4m1iAGPucK1Z/crzgPm3RWMjIhZUDXo6UYIZ4IeO774Srs
NwN5ZTjRjUk1eMYAaZF8Cu1emKDHcX09APw0u1Jimh5ZFkDovl0IJrSerkstaPGx
AuX0wq14xbcx4B6tgWUydKFztOnBX3BlK8ZrA7pSnUqMttkwQ+vbzd509d/DsCOW
XDs2LM/duvGbEaTV6KgT7kD/oVUW8XdolD6PEucL7K6e/X5XzIdXXovfXwaprlCj
2cQ/zEBIIF2ysHY6hkRCzsv1cSnzByNLz5vtOTKHAc9TzjWk8t7FAQjUJgx2qeZF
wnLeEJ9RxczTp5u77yJuUBx+LZ3MaypBGd9e+rEefD7u56PL7SabrndEs0BcO2BQ
pQjE1O1/zKW7u5B3PLObdXMZ50SqEVJ3sQm/mPBqukQYi7XTjFD+wRJqInJ2OMAv
4BBfVgSQELfc+nj5Iwloks1V2rjEnyBb7QfKafKmKEmA7BCcwJogJpDNTa06rBsp
C3l/oe9wWQlQaehrOh+5G3I6mjG+ULA7f4ycX1jDtYmoqouzCM5oT//v9l+PidbS
K70H88DHyHX23bPtkLiqD3SCDbnsg4rAhkVnd8OJN9acStZiV9OUepkOjPRHg1T7
NTAMx/dSMA6UGp7im88XMPCEFoYSRngW2L7R/11IoF5N0LmcxitgMTpL5JWbrE1V
zWQ8JpeOS69H0/4pRjMMJbUlfBZdIidGPD3sjRwLGS5CAU9p+iTDIvafZV3dzo4A
kT/RyEcPG1OSgxP75EvPaL3Jo7iH77jteFtb+3R73eEnjloFxcSb4Vxjz5C8ShZP
D7/26eq+OAxwSOsDI6MSQvCIO0GR04FhsaE13EhNoF12a3JrxpQeg5xaQ3au6LWL
2pUO17vUVvjE7p4f3YQTeeTPrIoxvrPgmZlW0mgTfu+afI6WpY2rfFm48Sf7quI0
U3Zby2UOduZpdZuFj8i3fEpvgctcCma+9ZMB1moTWlH7jw7iFVHc819F3T49r0Tt
Mda+k9Ni0Wj8dH1sxsIiJX7KSW6/KC3AdGeC3sJMg6FB7OPbZe6Ns3ZpwhZr9phA
46pJQbxkWNtCKINoPJ8eLAigNll1PRvRBkBRTSzBsyXmN4Vl0y4TW4d5TDGIRy2z
6gwyTxSzI6UJup/BpIIedtjmXa6rIEcr5SGAtLxm0cqihtRc5d7e+vprEietuGfl
WHcpVR+gAbk/HXDYH50d32O1Ook60JU+riekOg/bY/ZY6xXihCUuGTSyGpfj5tXY
pWAPDfTkRZ3sTosQSzeweAhTZ/Vc/hNdqkHjGuhg3bPaeqqgcOKeET2W9oAMLpcV
zUSV1ZOE3CIGVSjxQfLpV1oQ3QuoJpt3GIhYdFAVGxVOLwJVRq+ABWcAfKNVBTvD
lmIPQ2UIHwGHQPm5UNve59j05S5Noyl1nA/lMRj/BXp0itQtgsyMRjuZ2Rly1g6o
2OW1vZ6gSOd/DTWgiQCI3uyB+pJpAEvXeeRYpSiDIYzcEAHGUO8T7QRuXOzbbkO5
UJMCwYBdWo7rObS8md3TDGeJ9jj1C7wVewXKw5TZaqeBfrxUF7/FEMm4nAGKUzhi
2rUadv701iyN9mpcKsBeJR+A+xmyw/qhnR/JsLYAqYoPBrcwnfXjbTrXfEefCzIK
ZDrYmStpeSVDpMQQSJBVvbGcyMAnggIa/v5n5mK8klpXkPs+dY2Qpurb9AMk1eC7
1NSgNFp0VESsqSLLaBvc/LtiDvWryRe4OQWP2k5wotl6btBTQpAyWtukkmUk4KUp
l2S4Jnl+L/KKcXMHpILXEE9N9jNwa3VhvLvPayosOEx5l2HvmfcRuYX5O5+2oBIT
zWmH15gl4sLgZpLSLeMHqfCNwzpGy2yvn1tsj6yk/PZqWgoIqcmtPo6JCStrlJdz
91s3NRSjXdRWJ+dxVCUa7d3iL2IpjVINrDIk9Jge4J3hWZBwLnuYFzzd+yhKSp15
4QJOMGuOkg70kqqzIrcZrGzjYE6TrxMaDGIUlluaZKAwGXJwAVX1CISQHtt/9h2b
qRZ0uL4MoC4o2homn1X76CnC3d1RF23rSrS0hc5kMoP+wyD/rS5KW1SqhlNxgG8S
LJ3ISRUHki/xDnx35fs8Sy9xofF+mQtZmpmRn7NJYWE17Fxd2SS4a4piGSj2EWUX
xjDb2UAZ1WBIjKo5W7S2dxYzoqd8g5QsoOM7NatzlvDP30opqZFqZENBSby+VkVU
XtGu6qj4oRp0N4fEaM89w8+lMLN1SUmufMnGQtOliprt0PeS//wCjYf6//Nkmbr6
YgtXDeFiAkRid6pqv+AOU3e8WjyHPj/GzZdJOWSD2NcltwFYlw2YMwPNhnjbHDGL
mHFyEN0W5o4m/6xtek3zPFbISToMTbrL1oGaB+wW3J6iXkm7sLB7fkrz9vDf/1q2
57Fm10Up0QCxCgPWR5evLgZY5wUm53qzmZ6vw+fV/iFNgX9AqnI3FbiubOPGoG8/
LYzVVzG4iE1xfxEZCEqX2g2exfif0J9MxXg2tjYaZKc=
`protect END_PROTECTED
