`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a96d5ZLas0GBhE9UeeHFU6oWKHggQ5xhPbzUM4xCx0UgtMEtenliiIktFctgwLQn
PMO7t+r4/2nD5tut2u6pvU8F/GvLHrlCntKUv/0z2Eov7jmBL7+6iXgJEe9KiL+6
eRDjw/PeNI78mIR0y+HCNxhHwRIZ3D8w56BEHznAGhP3hgFG48XweqzzdinkI7TY
lJ8YWYY4rQw+DfiDoCZh4iq66lFbq54x0EluKeMA4iWhkLLFageLpqdiOjPahkgH
R+3NeupD02+OvpEY3wAbP6ZvG2G7PaZWTb+Hz8NQgl0aFmAuBnImtHOMjDb01HFv
DX56VDLEddhsgm0v22GBh4W64EjN6DaBWpvJmJWSdjjsDwKIAOVa3aNdbQoU9h7h
m/WN8mCf0AeODukblYAboEZUI/ysqhbvvyPn9SMlDeriFsr/O2g8Jd5ts9xrgcSf
PXYxD1XrFR4E7tzkQOnSFeYU4a+mZAwpz+Ho6HUgzUAvqgHn5AnQgE5xQkN8NjlA
eQ2bLaOs7DoOOygjzGJdYWQwO2zRHPY5HjNbwpwG5HC+hjQUbQPLFsJkbRAKs6Rp
bcGIYNsnqDzKPl5YG0+/JXaf48jOQBzxy9Fm5SW2jKtKRblbk3zbBMONIYqrVznz
G89RnJFpS/jfOZK+cSej3RvBIqMxbb6TxZymgvYIVwaU25ba2XxgNkgWpa/K9ZzY
qidEis2fMefzPIT7IIJZ7VFPQLcQVWRbkeZXP1Jq9ZVznvwbr8ceRxomOk28+DEb
zdOZOiY02Vw+mt2lQZaSJeWdCUuxGb+kw8sNaGdRp3nugOrKZ+fx3UiC3nS7TXZv
A6OmQacjIv3zd3F6BYHnBdwmlvG922yQeagNwGcCzs2ALKi4Ch5f81oNs3KDncx9
KRQ0X6GthySCTpj2It6OlcbYxXbGbHuqzqsIy8TLOJYLs/hyPspGz3gcsDUptTWA
I4bIw9RUzwiHEO9+J8/SLOmUNSsmFnZLQWy45GcZxEwKCDYtSiyUHymqpV0FIqxA
Lx/NNER2LZB49EMx0LM5OnviIxNBPiIB+LyANKNMqHSpd9j/SeIuIFhPJGeT/l9l
okRmlctbb3/sHWl/gzQ+oQvXzNzucMVTkoltdmGtq1XBJg0Ivdy4xDJY34/oJ1e/
ROeG1AtDdFK3fItvODDxATSSseylhz0t8gyvMwbDDB44O90R3VMxAHr8jqbZpsiU
zI2UbV/7GHTWQjWW2yBX6gcBqFVg2lk4NbFeHmmk8yU0uqSBBjPXrqqaza9spG5T
KFUwm//Igqg0vt2/we69eYHldfsX8QZLlFY/XHF355H6k+/PMh7XyJZ7MTShleO1
bssiSkY8aUNxrPXmrXJZmqPNKD9RZa0kf1Vp3cH16YcO9Fav+lczcZYaHGxT2dZO
cmaXj658QWGuC12gtNtX6rk4LM6U6bFyFZ/yG/qh7MPQI1usgTdf5XWD6B206Py5
0Zz1Rdvxv1qLxHngdgUssk8NzYMCx0u2F37ZM5GcAuirV5FamuDlPuDD7pVxrgWh
PqjJ4rbZ8zNjhgRY3Ho2IQ6sf7RvOiA/avXJHRJNU8Pl2Ayv0GTh3hyE4DJ9driB
tIks1yWePV52gBkNqQ7hhxC4FsP9y7XgWvfR7F5sBKntoax55xXiCRwnkT8nMzx2
7PX9FRixjEehI0zyiihX4kFFdqIXK5EI5tDKJWY1P8PvxFFqoPWv0v4J9A/L/5OP
odvOS3aqBj3/oqyOfBzW6ulxMmyU9+tablkO6dobMD8dqGxDrI2Ov97tjzrUkpPg
st0Y2JTtsYBB+UcCPGrdSUbQErSFrBdRuzeunRXj5x+VT3R9TjaM25DL/8o24WYD
yldjky4xdosgNm8midXfzQ==
`protect END_PROTECTED
