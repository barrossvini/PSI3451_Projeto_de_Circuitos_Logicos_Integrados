`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YrY3Lf3ncutkV8ldkdjtkaCI8GWb85JsvdihVFfyhF2chd5jSbmd+hQG1O/56LIn
wgFiVUjVNGEgMoS52xLUNNdQzckUsATFPcWW9a/QsnXH83wvdl/dERW97sXb3BEO
efmNP8jCx/Ahytm6QkSaGHpLUkkjCyshJvT0z/Mx6+2Xjx1WFHRTdZFhmjQ7AfZk
5qfVJasD64B4jgL3Nf67+Zhz3kW2aoW2UFt3IVm61cwd4zBvIJjjzQvM7ThzRGqn
Z/A2+UmzvWvmOUvDoXp1Sd66lDVHNTRkNQ2NzuhyFCcx347/aYymYxB8h7chTlkP
GoX43fYXrY/8CzGvp5vJHtf2q2ZVUNnoP4xutLyD/LCeqmts3DPO0MzbTG9nZRiD
zPSDo45jLSdJ0G94NLlISm1XKskrxP4y3DIHVbGQXEOBtdCK8PQVQe9HjxwdzbNw
LZ+2uAPtjWRXJTzYf+w4YhWVifhd/WFKgHDB3hhg2ZWC4OgNz7IL7Ao7QYX+xh/Y
H7YNpe+IzQoWwRKQADmLl6D2BJ1HzpyYJ/NwjMHKtzrgXOlSlc6LXZjM6gKvcLQK
oQz6oFVGeFj3TOs0TsBb+sse5sLMyFBhccEwFRImCTc88B6Fl+Y3xAnk1bJlSDJD
9Q8IMu5IsRtc49ykDnJSJt/o0exdXY6Qs9jF900QO84lhKwObdIOEYRvZt27pYBr
YyILWx65PsWKrUYuako0NQ7+0mVZRVEK6rIVTA9AdEHop0zPspLQu4dzKoVtREic
4ogSfA94hUP0v3pHgwpfaWO/uMdICpmZEtVm2d/xO/4xINAHDS4yLR38g6zCI6rs
l4taRzaIrTiszJ2jRNSjhSaZS5p/J/UV5dLYevBZDe+sAzxPx/8kYoZKP2cXotSc
OCtp5iH5pDiYLXC1N1vcAChgs13LTNFJ97I6FLU2Nbf/1mMtCzVrpw3ud56Nbaym
oi9zVGHbfiPyVZaSa5/9kQRlBmk3lxCYGIn621CrjVsDDXDj6n1hZkpyyTZuJnC2
48GMaSDctiLIqS4IgHY7+VeRcPvFzpymeyUM0gvLja03KNMkpMqkalB+4wC6qd7E
eaOKnK84wTy1HuLtrLnwGB7ZmCYxSRS9AQCDL2c69ZnHCUJ82ra8XRB52BiWsN3E
xgbkX2JgPFlmx8JH6ipZHAGfm/nVDRLIExlO51R5SSW218PwGh8VZFrL/nYI1t7r
vx3NWSrrGybib2QRQZrPpgk357QsJptPpD1OhBtzFZ4WmgcXRG7v1eDXn2kxsPZ0
fOR5NJqf2q0GPssyHaNz3ehp+TKHJ/8dminhJR0+N2WADjTugc6dzuWzzsxFF96y
/1Cneek8WFOz2csrcf+lVm/J/oncEolGwu8n48V3U3k3+15n+gZnEXWaqeavz4ul
gaXJ6eOrsJqpQmQCbrR+OxTXHmVYEMuQlpZROH3SAMBAEIbbT0tcBdhq7Wdmjfi6
cK+jirgBTZJ57e5w2CZQ+DJUYD6+npT6bMiSL0cNXhQ7b215ygOoyi6OM36AbUuG
E3NevcdG8CZHnKiDcx/PYOhNDvXRvQ2y/eMqQNJOOZhMcL7gazgxrkqF+FHn/2iR
o80onW4eJ38LSaQFPfsej3w6/PeSCvo7KP5s1IgS6tgevo8vVbxPK/U0JqQh6M0p
GTM7Eu6PQDKVWCxZOB5IUtBcc+vsc75OWVmpNHUZQEaHcho3i5Rl2+88G9yHoVlY
YCO5Y1NsNKqaVNMO95qqLA2OVxQTyUimZl195oIA/6Vjrcayht4Op7lk192e6OOp
8rJUqCh63Y2YBc5cC/8gWANksE18HoNP3rkv0cINkQAgWy0Qxka+qzeRk9GVFvSJ
uzjQjR1hTedUlT1iX5coC8X2aoUJe1hpkAw939IA5769vZNDWyJ088ZK+0ZdCsfx
UAHiWANr/gaBDHKUnmSD4TQunr9BFIqs/rdcJ/PKstO9nJ3RJenqgS8eMt8ObR+E
46rb4gdGScJ9GWUsTv9tpkCKLNQvYdUwYpIAC5iNw3FNK2Wq+XnO78A3xtCZALqv
AqF4UaBsmEQDqv7BPUIikaE5CncLxJU/fibrn2WynRHPeEHr1gGmEV4Vmu8SCHny
Ub1GZIwaJsH1YEBFq+WIIMBqEg9rhk49ZzVMvhVv4M6GIaEcjbgQyYyQXlHqEQ8T
6CgbRZ9lpSlKJOzcnHxUnSxSpAR1x+Guaxex+LN6/w6eVCkcqMMyI1CgRIQ2XsYW
eQ2E55wakjTYkos7sVfvBSsqU/84poEqglzkXqFf2ySMmQsHGdvhohaGIOkORIFk
24//Kk4Zjrp2W/XuuMoIkNKPRuLzGMutrI5hUXEC36zNfov/Kbnltj7OQpH7CNE3
ROg9i2PkUVG8wt7Q6/WSkTE3BSyXY95wRB5cpCGUDl1r67F+KpPir/kSvHhXSA5Y
ANePbZpukW5hDCnVmRJj8HqZmTAZLJiiN4wK5oadbAaku2Mc7rDUnF/T8XD2GrXt
gjmG+BmfeTtajJWHNxDpZG+vwbpTgfVQegwDFlCYEd88gb3SEBRJXKz/nPsLv7WD
BiJ7pjygntYQrEADEtJPLTfL19Xk0KKc3h4+8pIOPE1kBB1Pg8BieeDybEPcns/f
bmKwSCSzJTIm5h3eZEOHh+cTJpjIPkgtEh+bMhxlYjjATiJ6SZOHqziLuS+8zgVU
g68sY1Rya35AvNWS9FoBoFFAufFaCVGW97pE4wXIgFSWusjyxE3TryLnoevvHwxG
msH27HNaac2LXJLdF15L5m4SXb9jPrwBOaUun0qL4RKvBO92V/kAemp0IT6k/hA5
a0+fskjKr8txhj0zjHFfqRp36WTmtUveTI60pH7DrpG9MhSoDtpNQbIgsY9i8MpF
dt8JM3i3kGcdkTXViUOV+ZdOz7DEV+orwsfmn+7hJ8vtaY7pG88u/fjGQANiaHJu
KBrhpdSdf59NtVh53uOVKIbMPbxMt1piqVo6K6j1f1dwvZYwylbr/xddvA+na78/
MOiiq9xato1YCo1lxC+oTUm/M3JDkLy39s18QyoI/cK78hRAcTwByc9wrZ5XzoqO
nk+IUTnooIkGpUXiaSiQjzipAFkEr8/IJdQtuPaW6AnM2j8Nn779RjGQ4sJmIPrA
zn4zgy9FZKTowzVRRu0A+09Im825PMxEGfjLqYNp/NQ/yRkxuuVjpBwBoz0NgAEU
+jUZeb2GwexxHWvrNQ+yHiVigSlu2PWWlUW1qE7Q7HaKnpVrJNsdKyr8zVAOSX70
Msy1cMPYKlt67079BmLBiO3S1m1bu98w39gv2rZBCc4hcYkntdqkriIXdxttRF1e
kdSD0X5/8zmqhQ0N37vB3kToDWL9TT22+mRpY5a9YpLKH99iqR+KcTyh58MmAtUm
2kQmqHeert8/PW2tR7Q+r2t2N3WFjuOYfkfYG0+RBNgs5S6fGjgG/NRb7qQRT62P
JhdioCb9w0JktVyB8zmCFm2dTLzGyn7DE28t+OwtX9vhDPqMXAUZLsDkdCdEkBWs
yHmHmon8glCjrok0Y0M+S3KSycTh0oc61So+h/z3hgcCVGExN8DnA2eh+j63qlW4
+MfOAr7UZZwWmWmBnU0+gJJU9JEXbHbSumhZw2GIHb+ePL3dq4v2pYopdVUOcEgG
mEGwCdGYpcVzWjPMsR3Lc9Q7edpzScP1hzqSf+zVjpO7JOYsVsl6/+Va9Snmwtpk
boZiRfSXHqvoljUgEykYElHliW9djHA4JfG+UodJ4XBnLlyq+hse8IsXGsxJmtRe
v3nWWKK42EmZTPsbLQLoBfi8yiB3csLoRUhX4BUT9hku9AVV39l8gjFvcGqi1fQo
d++SHjQ/WWKN3AbQQjtXoqbG2Jd+h0fk3oT2uNWW+HNtg68iEEpTwzA/9W9W8jtb
pbZcCbiMGSemHi/5mluhzZQ/IJHunnioWg0V4OC7yZ42H0ge6iplSujLvxNfDHzC
+LSAzCFYa2eS/46y/qsuZ996RK1pHS3n2eOQmX46caO64b4GpPKm2Zg9POtPE13n
Q/qaQ9X540MQqhtXEB2WRDeV2o4sAfiDIQMYZKe1ZOaMnJUouNcu8zZzpfQqkqb4
iOvoKnnQKNmU/Uf9qgPelIx3xJqA4kNgJywlH4tmRMlY2/O8R0tVeC6G9IE9imEa
C49rp2bf4Nv8BJ1UdtjsPklYJ2+CN9C9bgsw2jUWOl/KGglApR8gSve0IGthObRJ
35MuFEDMJBMG7SFXzAvkVP4sW5GuIuRWp8ItbMk4l+h8rOPYQDylGCqHsGz6LG2v
ubdDorpBH2MRkwOcW4eK3qlYYv4ajbYavPDabrkY9gkfCUsUN900GHzTjJPz9lni
+77eCfB3Jkz1dRph7IYNNPok1NKuKiGq4iay2D4NDhSSnByJfqlnXYm30A4GieOR
Pa7pmEF0EfKF8u8rIGQaryCGRJRj32d1Eags6pJ+3z/QPFfcy+jjAHAbYZP8l/tl
8VikZ6PNAZztI5qKNViI1bKs/y0vPEl63ryqjN/XENJBs1t2919qCK3XeU8x2le8
laRbpiqm+2z0e5bLeOzdMuNU3HHh+QnxC9wYZLPLmc18lVzpWWPlAXiy7I4qBzlv
03K4jDitIORT3n2Z5pqmxv0OYHPQc9zjr9xy7UqtnfoUo/OPtNK8Mwp5iNZa9OFp
WVHfdRjiRNDMXxSzzV/KPcRSB82CkIu4VbL8+/PR3u426vBsDNthMJfgaL+o8AB1
NOXCKx3SFOP1wpFMRum5R++Mhx9Bgx6HzQVM14EAVuXRjGAA3Wv/g+mNACgAFC3P
yIqC3T5mhWwm34uU/HsNWEoXqEXvRp13Yuzk4KC+iGvzmT0M45WumufStTNLk+3e
zqgLDE4Uavaz1MhPTDqCvjSxQytVQQbYn7xt8i4TD3t3FpG3+QS36uXu4ET2L0AQ
r0BKLkLOyHCOIvQHcsiBdVQj/QzRLhYrZ07EvCrRh2ZbihDrSYp27WI3Ox/2yqQ7
HtHWlbLbLmW+TnXUr4gwnbf6itZCtc5A0KqwDuZ1E33OGBH7bWNNC7VtNQP7YtBY
TllW3aPO6qsKwSmZQ2ZngFjzDMwXMRlDrnJ5UExOKY1TrfeUVdGlmH2fCTJVpMpL
cmseo//ZVgRreQeS7qPysqp9XArxPbOMMqw24ejAxUpbrIotfPFsro278QTvvzVK
E7oFE5cLts7UsYi3LuaESP2nrXs0c1k8+oKaovPjJ1292SxzApXhZZQ0opS9HhRO
GOVyj3/JzcE+edGfjqaiQsimXZkrPVJ/WntEA3B5eje5l5T5yQ5RDPrGGiST3G4H
uytLPkp1tCC8px+kE9AeSOhthadRMwoHB5Ts+lwbOg0/Wv4n1xarJ3PxHvDRplbH
vM9Vd/JFJeozJh/11gUEy+tnTr3Tsm2SW+7oGCAEfaCZ33HrwFdsr/Hhv/Q7L0mT
6amf3CCwZCItLRpBPxb40I2LRipmK/onWuaBD73P6N3QDtT/yioZgZ77/uyeiwN6
F09knSWYHRYwXRJkFEHTwYx3NTFZw8C/LoSMRv2FnkAqoAzQvlUbcQiR0C7GqBKL
+KjdrXctOdeGIgaq+V9KvtoCIzGHF5ndtQJVio41gJYIu/1LUmdvklDADeKey5py
zMXr6u7nC9TRglz+DYaU4vb0b3hKrqMM1naEW4iGsXMrQa1GGXjBryPMxpnbxqlx
guULksn1Di6hm6VHmcoIdw/u6uF2963HG+XBk/BZc/D9DHGCZSGPhDsfBKnpKUrV
nv+h9tgaPQCA3puLw0E12h4ao5uy5srXSLaBgYA/8njDf40/rJaFKoOBjAovFgQK
ZKgc+DoYVTd3GCyivnu7ElLkP5czu+1Xuxd3g7vM853skzIjDWzUQMrEf28b11xk
vf6bUwGbeYpxz1Eu1QCq0NKoifWtrsoo36KS3h0zXGGTCOOCrHVMM23SGZWMSviW
fsdj2kYu3JYTKbpqV8rDQRe5ROcOy1Tu/IPiAPtOfzesKwUHixhz9aflvkZZEoaf
icMbZ7CrWDzU4yBlBsej+R94FU9bB7gTNothfJEipLR6KEL/497BRJGK0nfaAmv3
Mgo0rxtNYERd4RxR2heaJs+509SR8nCLfeYOmiu7hM7+BCqkOLOSMQPAsC93fQTV
vtuInTX7WONCmp99qtPLgLgRQu2m2XGHOXhIBd/jQg2NR4vLgt/4WqdK+EJeNHbh
BGcYUY/p1sqZ2lcbdM3deZnSImvQVaON1dVc3ZIrc8BX8oXAfV12/rM+5aWcPJVZ
mUeb4UXDPJ+Z8yug+b4EWBBOdwPbbjgKg3FfZZsXgUqs374wCKhoioSykz74RWlQ
a14FtSsJhJjPR3+Pl5j/WmEzqUVsoa0I8pt3hPZ4GJWjrkDcksRoFWxQDpY6RlK7
oZ7xaihL/vU4UMRJpjHiYRdHibbKVPibpgUSNxYyWyDR3wSa+3lhLARQVHZqq5DF
LPHWvbGlOloQNbCq7ZRp71WApHoiaM7/Wo67IDcpm74PoQLUgZq+TxVWYO7oPZmJ
FRudCaHjJ2PAubAexOm8SSZJPMkkfjMBwUIpYw9VM9rxR+3S2CKcoD+aspDiZkga
yafT8jccGPCTetmnUaaaPsT1kgHl2+qconZoUb2fANkM3gnnLEVx5IkiScDNITk7
ttdZvP4ZJfGper4IgV1IIeWaUGOfoRac4MtZkE5zK2SOopOTSLwj8XdJtogBGPPg
DDS3k6ljSd0kvOo1rqslzX2RAZXI1BJf9eHUZsl2Ecvsww1a3WWXVP/TPZJi+L6y
UHd134mZWDqCqKqrQB1A3YZavyEGr+SszM0jDYeKGJsuju8CpVk6DjRfHqf7sljU
FZKvHSRVip2WrMYKfuZ3AbzX7sNzpM5m5qaDDhY4DQn1Nr7lrCyQ52jNROuzSNFx
wH18vyXR/TpNL8k7/6/klHu5HZ6QU+4uXKLE1wZhvIntGuF8afe2dIDYgnREjjmW
6aik9KlGJS/Qxevs5J1xexQqY1JuY1q7zNrvyUFdbiDFwt0Gb38FAdU+wNXey0JW
FuImnz3nYYbSxDFz+nLae6PMYm3AQuIcVng7EWPazDkuk+SSLtp5bMXma7t9kIT3
W/GeOsFEL0Qmt+7SykKfpfHT4SH8yV44Y+iMVAsBqz+nYTdaG3Ncloq/f+QsTomd
tDDLTUf0+J6+VN0ynbby3KUtVlzlGsP0V2rRPXJ+F6VRj3GUTRF/5k6hIl9KDVJt
AX9T2u3e0ErIpUMnUFT+4id6dH6hCdo9928c0QKvXqoq0UmGu2X0rdHE5GepnbdK
GEhyqC8qdjaS+pfGp33ZNA==
`protect END_PROTECTED
