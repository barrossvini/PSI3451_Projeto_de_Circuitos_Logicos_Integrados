`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+JmdFSKVxlKrsAOYI30fBi900CXemPk400XSIAWuXUIPpQvV0yYjn2jzqupPrDlP
omWow/C9d1tXdXlOuiO2NbG5RoZwMDHWECaO+gHHqOOoXozctp9DEDxfHfXT7/CN
vjIpmzGehJn1sdOfx5kMBpn4way3rq0Vexw8+Ie8qzNPi8eZ2Rwi4TeHC/JdLr/6
RFZCrhYSvLE/JX/crIJwcQ9HKzE+DSBhXhn6R0A/WhvYWJ/XbJ00DIDjRqSn7un1
kWPNsD7L6KSBhyRXntoYnRoqZ2ly1b0+FQ2E1wYyXhKC8xw9WokTdN2TfeTGVseX
a4onG1GUqaqWLI2lfBSay+EJUUEPHPELYO7xjDSv74Ov6NK+D1jifq3WJlnpTtLq
5eSxbBmVdtbj2mYNKxsventYDY7DPnDeZDskneyOwus3KkvCiS3c6o7jajJJL9BM
4L2E24jLWf6l+BWBUeBjhpUCbAnLeuHYtQq1Bw5Fcnp+Y3MOusLDCLC8IN//sOO0
3t+2Ut4cQShCGXroGq9cFX7Ba55hDePDAhI7N/6r9kUASrD1eNBnWOnmYgo1tPra
sAgoVp3akFlbrzvuwA+rRcwZgOmHEB3YTADF/2fpX6uGSj4rmebuC0erg697hcl/
w9RXzhUdU4tGhAFWQ/NcRpmpaKx5tkwnn0LJ9ZbL/M+hv0+hjYQRG/Lrnf4INW50
6zJVISO+diMDoMGaV++JUZ+rs9cBiiMZE/UgZfwvafIuyezUmN9rJt++L8ChGmeF
xV6pVXEwGsr9MuGc9x62XAVsez5i8aD6ZH+6NC7ndKSln8AEi1RrlrbJjr76sP2o
PbVFcFkt2ZzKlfkPw66PWsOCX/jAlmrbB3eTDnZBbUYAKXLhGugFg2UYezqsug8b
S+vwQUQ9pDB487p5538NKwiFzGvf4gzT8a+YE54yj4VfzHJGRuK4HqHcyRKLxHO4
hnW6EtwLXU37Nabphoj3a140Ku6ztiKgmZ6dII96cA2a5SfVaSZBebitOlukYRv0
XACB75FBrD+rrdYYRxUx8oUyM4WvrNDeUxeXEAInqoq6MaUH18yiy+bNdDhj0xu9
Ri8BwTtkySMoIIqUZpgjvB4yktlXXPpeXn74Hl6IgM7076FN8qkGUfVAEGnqzI17
2iQAYQKeh2tO8OQf8KDbRbMdlOc6RvcBdt8hdCt1VZsJ8jB/m+HTG90FVbxCS0dw
LFZWujJOHrk4z4B4GVaIYeWyoWWjTfV7HiQFmoOZ8kzv4Mx1PI4oS2QcAyaqDvg8
Goc2Drqe9yh4Tm62rxeUNqwtHNn4g3sQHXLmRTnd9QC5U0VwO+MMbjbZN0jbNqlg
ZNaimAijccRKh2VwFNAllAgtwpyX7RWymNWU5MaggCP0V6HhA0+E92souzFwEyA6
XkvQlAve/WogxyEfStEaQbuVOJONDEgdXMB8LsoV1NHBzeYdosv3bWrYoBuJdPIG
OLUEGDwBUDS2mOtB2HDrNT4UK1+6WYCm0Lpg3DtnIjytK5KhANJwyNb5VUUVJ1HF
REq/tB4deJGAfTLn4C9/0zzHkM4B6//gc45RTlEA8R0sqIS7MWQ/mRGWtJ4hT9PO
eCcmszOa9XevhMCoSiYBk7BpLBB4PE+srjU3HpLB3msbCw6yuUBpedzD9mUKwUUz
nxd/GBLFzI5VUBldOJz/nylHqsqzMp4/fC4C0sr9ApuZUYlpZDUqUR6PISunj1TG
0sYh6svyTNBy/K6nS4A+JPn6G7NhZAc+t1Iloj5ga0igoZB8+um35aOKXTCD91VJ
CbMOIWHwXhQHrBI7YQ12r3G/naHOPhpIquixC0HvHW7NeSLRS5bkLbQEqwVb0B5j
n8zbYOmVtUGBngXABiju5+CXWB6N2qPhAsuYRbgJNYy/Y3eMNWZzmUfZtjHgqr6w
jaq1j/oGeNvwqSb4g+NfPDG1pL9HUtBPYmHUr0FDZ05gsyZ7PyZY4mfv6EfHWtcf
NVK1IZJI6w91Xbq9Eqf3KgtrrrV+TKhjsGHO36+CoNDDUZvraKce7EpL+X4XzFxN
8TLYbxBpJ3SCrVSX+mnpBQCkEWunc7ztW+ZcvRr6D9FwI8QIVVp2NrpWkKbPqdRJ
xaetOE8f/aed2YEtehnBfaoXpQ0PJIx86Ehp/UGT6MzvZSvriivP7HfY8mBGnJUg
jCkw8c/U7uEHSWDkzkZT1wQT7BZMgQe5wVBgaICOpwrb2Ffp6eg1SAlrbIHmGakf
Ok9VVAFfBc6z25P4f1F3rTt47lg1OcfBEcrp2CepO1WcqFqgOrmpLzs21yn91Trn
Hkcmg4WdFe31hSSs7zHvt/AG+qbp3FIYgVhN9bLLR07EtkHFIPsaJrvBvRefV9bs
E7hrcRqeZUjNCXk/lzAMxdQ9qzNyECacKxnaHEDb3nWcrafVxVANIJc7kl6zBpEK
OzNgkqhwfbIog5eeE9EfYMCjxMwO7mRul8aIGY+giXFmkdDMOM7w9EAocBy8CSVM
GG9XclMLqjpnLzkL9vMJOQ4TOm5+rY7jKPnUq/HMjzAC1DcowlXRHsYDosDepbQi
DKM5EmnJ0uc59vkSz9ye5cCFyYUalB0Pj5J07wuzS+G2GDLp6CSBoXhD4xKA9ydA
Fn1NKXAihNmzqUEbQ3dhGc5C8Icqp8PDX+ToRyPcV6id4kiCiYivDcatGqdmgqND
0YjA+VqEMZ4q1WDP7I2BzzjwsrtPnwh6L/jAO10wRMCJ2Qb6IS0V3oPy9mUUMY0W
FnktlWCn/OohKY0MpcDWX3dxIzJSzIUewvtA/4SbaAtq2SO37RF0ukIdSSISLPPk
K0qK4iIHjzdVFpjtZEW0a9ZIfqNk9NWquK9fmYuAmfyz/QoZ2iT7ClaCYoywt8oV
Y/gCC8CeZhtertZhUMh1J3fF2K+xc5uwPmWhfLnn0OQ=
`protect END_PROTECTED
