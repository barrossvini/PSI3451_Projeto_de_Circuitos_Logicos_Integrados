`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oRNtZVqaGSzZi/fgRwLhm2kKPAuM7c5qD7GsQEvTBdW3Wy+DDxmSdJ9LXbF6trWJ
9+hxymw65v/qXprHMOjtLnB1Ozc0nVyoDwxmUQnF7tJxMjJioC3Y4Rkx0RDdRq2+
0w9AAD41NBLJGmM2D5BVi3firaApNGcfgdJWex3YVNpGLSLmGt6xowEDQa/GyGAC
uI+5XVzGim1Lovvii6VzVIyq9vkBGSv9rPsU1Oj4HMZ8rSGNRHxZMTg5YuJI8Lwf
suwSNTF1eBu9trgv93Eh8hSo0z+LFPFsEaC9BuB4uO3MYGQytz9zbuThy3h5dHIX
WFhYVWbWTg82Dond7TfgiREt3pzJ559UqJp9n8ZWJjhZl5frZKkwTWPrbFux5dI1
NZUvr6ix1RS+zpfPKW/o1LD/KnyXrzVbccpBwaioBCS7VYAPXVCevelcnPvlrjIY
VIqUOu/WlYc+m/AUgvrmHwD3esibNsy0rCDb3vl3p6WaOjNBpbP/ttEuN4S0M/O7
BcTTQqpqTfpgemHGTyTsn1DTJeE121Ci1yleY4KOrM0N0q25ojt+9e5gUFGBlGXp
x1RlNB//NTrBaCd4mDPt+B9uQLeSjAS7AQFKamNDiSO/SAny6G4heotFl37Pwnvn
gt5qPRVguld29jpJDcRO9qOvemvoMB5kLa8uc7A2nVZiEFeOuyVeTe1Vne83mP2/
mQZpUxEbpehb2R979jlW/eLoivsDLeeDSHN29ot+M4K9w+yDgZzTa9dyAntXXYGX
qllboJ+SOCMT2ssYHBLgvylbYfNr68AcIXTyYjHN6gwzJd9VAEAVg0jIk/Q9P39S
rkdTPquxekvmnynpYAQWDcCF6JEDOmwOTNTiqeGbb8LbKHY1H1WGiodNDCgSTS4B
TXoTo2VUF/5umhXgB3l6KUtJjED7tewGFEu1K5QbTEWSiohH5rMWH81+8ZkQ9Fuy
FWjiAFnKjLMUnak2IcDzjuOLKDMt+M70bBixJtiuTJHmM+19TJb6AoTSnHGoEgjR
W0ze7DvF5l5/N9/WKCknuyfqQkdQLZGSTehdPrdDIy9D3OYUaHolGmUSAOihqDqb
kaeq6hAODoa+L78ClKhT/677fujEtCCei7716zM6/kUzqmJuBIeJ95+Ou1jzRIKl
vpAd7HPL8kxJ9rxlgV2V6AI5BIrf6JY3XqeyvZHkOmOJ6q2EfJiNHu+sMA8ox81B
1C42mexHQNORU5u7pT01X1MFDBmOmre57vu+ZIvMMq3+0hwjTX3QDkjMlAzQTSPf
7o4QcA1BPVhmI9jsmqd1/uL30ug+i2QiB5mWGH42iQzDi120lIwgTZiRHlrDeWii
AyE1I9SQ7CR/LxFIOpBAQ4KwROpdST8o0BCFE4Z82URPLlsPlWqgwsQbYPSGtKK3
RbXXiGUEZ37tUEhsEOwo92E6AEgw6ymDj99wP2ckaI/RVqM+fnrFLv65juBV8U0p
YvfVdJBVrjJa4kSSGRKccE+lmjVcX0tLouuHk/8PbKcb1voeG8Mc1UZ43dRljVN5
PcqWNiYK8SzVEsg9TlAsfrFZ9nKJnt95E6PttdVP57YRsc4ESaJTwntoPXmsIbcN
8F9a/QovZllQBErbCijI4fEU7989aZ7gapMUvoCa6agLDSp7fp0Tfs2fIkeCzGwZ
iB2HRx0GQBWXxoos5NftJ545sSkcv9xAbA42mC8xhc4YVXMSuQXnzpUo5Pza70yu
p1kh9DmT7R9Ke/Msj8jxgQMjb/tHvCBVthEQVfC0huzdizXMPWtlyqwgnkXfLU/J
UpRioA1SFXlewx7vOltuYFxFKMWHNBE5UVABw8LcVy3eqDoBCTgnfFxv45CVr/LP
Rz20286cnBxYR061v1KFJMRbwjjC1lxts+LewaGupInTpOC0Yyo3ZXNzcaHMbceh
yvh09ICuRmLDu38+xiylbPMw/mMnMVyryzxDONKkPiVzMuaR0f1u5PL7ipSNu7eS
pEmiSh9wZP4a3UIHlsUQxMPQKBMbWkyxF50QyhBaN4pvTlfkSM81vg8eKB2jUOiR
8mi4VjJM/0BJu5ysbTtk1+BbpCKAs8Vxa8NcETjPste8SlQoCoJUsU4HR5MqR1+Q
pVbJI1PYtYnNev+2lgZkhPYobJ/ZsAvpWFj6bWitq+fZfs8GPqfcQhHPOdteEX/z
y/PNcEKKbLXa1fQX1aTs3c1rgpMB9F8QsGdFl+45TMKTmZzFrZ6c+6vhpE6B3lHl
SlX3D1sUyYLD+fy3WxLkxsZy9mHj9saQW8ibw71WLglPM0QRlTVVkR69XQx08e/w
4+kjP2jHIHXTGfYCD6/5tWsdwAJ8f3ShrWIJ1Ndg4v4SjTqkRueQShLSWUjdBfqM
ikaUfpZJp4xscaa/9F+XM4QXG45K2Cr0NDqSRZqzs3ZyPzodB9jMcIQn26F3LwkA
0kdVA+MvbtoTyBzoMfsBElAe4zRkecfx7lC0thvUpGKmK09CX9YdbkhdKoJHOiJu
cSwKgTv/xcKxIlikXmVkLiwu8V82zEFLbeQ7AOsNHyCJ/Int3EMaxjg+jwf6bJmC
wsAGwGXBK5bRRkF8DemZQHEc6J54JzwNaCzssPRYGX+yQDrt6WrlCUpbFfet0UF3
6hsuzMdxLznahUqpsnFD6IDUoM3B7P8CCSXd93tQSaKC+zcrZVGLd1dVjnJV+xDe
71PgoAp0xdy+Y2boVQX9QxTNYVj+BMP4IDENClyClkj7H5RqV2bcS0mJa6OFkMuA
OghuM4ndJpmFWSPxvqC7+UQiEzHVhMqvy9u3g9NDVYvK815XP806/vuscg+jE9Td
USm2Zf+GeCD/dS63UuLCyL16934G6TQT70ooH7joDwkSF+mWAKzvhotLvC6YWygI
tenorIf1rs/qS7jdEiFYA+eKDOPu77vCzokxXPMpPU20+FMBrBAuACWV4eKQ+iUr
rVeI5vvYF14lSSbG+K7VxR6KFs9u9QUZfwpKoy6ef2DWNHBlTcZbeP7RlzODrHnj
VSvjcbSaGhoJYlKt2EuJhmoIeZ+uEynm5y706cL8J0LbKBdqct8g18fBBWDR69CY
Hy18+bw8juorqeCXFkmJe19jn1wfMBQ72EXITKGP82peZsllJ7BwVE4VzhPHnv9I
71eE7t58m2tg1qIcYRQPeNA+CTMOhQO0f9FUOjENpoeILcaG27XBrE5syklZ29c1
pctyH4fPX0RSm8c+v/E2h3WOjZPE2HOiXKGnsAwKuG6gnQhs5FFXzRmq4zhOOdpJ
iAIk8icpOv/K98UzGFuPxBCfZQAq3iF8+RolfeiLqisWzqTUbBUDbTnB6Z42YfGk
hdyWzYEkPFc5FlH0XN7IuFzxbsM+1HgUSkTOP94GQNdhqMHzgxwRep47d5py5MrL
6wo/albb2YrWjxJPnIGJkEp9a3sl9HCFttHiJrwUaPTqzgdDRq7zgb5VgXZ3GTMt
fTJEi4eBeNhagZ6IM187xW3m+Uizi5ym9SSvPPjSnRqwOD3QA/OqsGxZzJ5+/Oxa
/1/FAYwgbGlOEOCWrDNFedjoU6axs/z68ijQ7rfrAhzhbM4/NDV9nGKof7va3mYK
fQlqX59IfxoiXNMuh7+5VuA/KnEUrQAizDzzfPaQb7ay4PH4ryJCWlDMuTwGH4JF
9Jz54HiKux6mhBPawVs+HNUV5RDAfdixR/rX637Qr1WnaVDO7gWznZPTujHx+tAi
QlxU9bYXSasQlZoGhU1m2xrxYjKpRK4i6qdNAn4XMa7F3GV/UC+t+37MecZrzjTE
awajunL6lGj9M1flswAkv1HPXxegAB6Nb0jULJpErcRnF7bV03dc6mezIYIQjLvh
uwdSkpj2FRpEEwRaJbfZfHWv/9s4p///XV00igOda55nMuRir+09/460jbujD+pK
XYBFA6mmnCn+CYUeIrBDpWWVwn2+kFcyzoaEvvKn5UcvxqDEmyIOK5D/YacJH8De
JYKBRHhZB9JSb7QyyiwW7AWzMtNHidpsQ10Jgp5mmPI=
`protect END_PROTECTED
