`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VuJVhXHBlI9zcWgqNjU1UQA+0eOD3+6lO18VKg02uzc8TLNX5ppdtXUKqXAWbaUq
+q/UgOp3ylupHLJJlc1Yp2ucS23+AsZsb9DYgwxRVT/4zPdeLFBZcNxjLwNuCQHj
biMy322PUPvHpAXFzEd8zf92PU93fNbAVi460Mipo2O2d2aVuLNu59Xfne8t+BGO
jqwKpBhHoFMm36PJ3WZFC0YVLPJzQK99gOEyxpQEmQMygs2+PaSlEL0zYz9ZL3/+
07UaSoEh7uaWMCMrbg01wWsDdezPveUd6Zw3Lcv6+qva7kcAxJGUROX7eLWNPUuD
vj0s6FhtJFU70+RtY/Vd7JhzTiV8F8JnvF6vJJvw9FzqWDYYMneDFy5wRWgAvpua
RI0ZAHWu0OXb33rcy9xQEF4QgHC2pkBgDKl9VaJQvGOlwGVWBbUNyoaODubiIjci
tXhNvBEG5lbbByvK10SczYIGm9UsaznTtSvYAmIujvy7lcdPKP+dJkR0IRY1o6Xt
nbtHJ/NHXUIkbP94lQpO2dP7aMjG9lMiV+jfbwiJ+vAmxiZ5KBP85EUC3/ezSnwP
oq9sAZSzPrj+j/BhBy384MDgJW6q2oCmkPjV4Eebajs9j+BiamDIs3CIe2i0krRU
ZQ2X/lhSyb6iMaTAfQSlNEiHWNvF62vXtsY2M/YcDV5sfVB9Nl7N8xORYH6OkDbt
UkRU/1VBKIWoOVmyOLjzH/BpYms/eJQnOZe4WILSzM8YXFeQbf3wlwdTqN5CeLyN
glGOy1H2en9owa9FtTjLIlknSVQieomS+373U/0I6Of+fVEeNZm5zQt5P5TFGJHK
Nevgl9wtkDBp8yNjkvvfmiiuUgwaSv7eew41vrxU/KSZf22IBdRNT4n7kGeiMFMO
JLJt3crUNGLjZb+RF424LQj/ba3mVinaMi7PIybw16rHSmmlLlZUWQnVwptRe+nx
DRS0yZq9Iz1yhkCQ+YGHM9wnFA2vzy+IG3+GDn+oXaqehnM3x+5Opqbp7vLV1BBw
nsRD8Q3WW4LtEmrDiyWRTNJazdGyiSI2E9uVwBASYn/2efRnnmv9qjiQVaioQ1VO
eKZZZTSLQeJ/jOxyvjM0OiC8bzfVQMTasvyAITdiZcrt1GY3166XE+IkZUP5ON/l
LuNehKq54udIosLpHq+0Dg==
`protect END_PROTECTED
