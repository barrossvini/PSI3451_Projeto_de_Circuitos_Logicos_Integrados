`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OZqkDttqAlV6hdgjxBygo4qrEghFFQ/s6f7KYFOCUjcj0Hfrp9U4Tj7+bkdqwYQz
WTqwmUOLD7Waq+oI3zW0GPXhfFmM7qgUHFlFQ8tYzDgMC2EyuFnyuokEEnsjAYmx
5tI1YIraZvwXphHrY2aSI93Nd9dUw9jeTL8seAIX860=
`protect END_PROTECTED
