`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P3+vFr69oYAKLGbJG3lDwo8TDe0pILw/luLMEtfscAvQclIq/FsrPz/YNZzl6LDh
o59Nw5gwt7xwkCHTn/wXw9BaRraHZF/3s3Y53J6thzKnSSO++xq7S8pxiZqnptU9
qu1sD1IWYEgMnpeyZxGL8KtfoFC/ps4lYEGycgNLbJetFSWi/cLxcb1Bn7d3qUa1
E/yQQPVvVS2UZhpY5g+oWNfzpLHBlTDatwd256qXjqZw6cQn2Q4O75PyMxfLEJ3U
24vFaMsCGmotB9B4Ch4dkjvnqAggkxh5IqMnPhJG+kv2F+dE+BRpnlGckw1CHjAM
TJ7fnYB795olGkU5o7XUf1o4laLR6Z9TXKhKSo7tHUUJO7ZhxYWI7knc8uYwvl96
K6MvqL23SUpc5n0vAQvGleAYB+afYPR+rIKOpsUL4A8GEmiFiQfD2Q2qMLhXjpVi
78XOp2utVvpsCXyJ0QPvaZaLjBiViRUkSrx7kGXHu0FlECXCVK5cP8N50yQN/kri
8FHO+NSXByfPFwzSsFwzmMsGwmf9dl6DZ7V02GIAc2LhGEm42gQWXIa2gY7t4Knf
kkYis0yKge685qVRQJuTrM0LdIy0ugi1tuZ7fVt7YQSsIEN4bXMVXTLuoIMxp006
`protect END_PROTECTED
