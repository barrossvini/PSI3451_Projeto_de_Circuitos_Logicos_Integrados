`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X6xte6Y2x2POOjlp1DzXWiSxUACpj/1ypXzzqpUwgBqeUCXHmfL4M+1BKaKlR5Wm
IHgnVQ0OBhrvzHeINkXc8QQJvRQ2km+h8tLMxGmy5HGBmb8Zrj3tYYBbMETBziFG
80d28nESqtrURtyBRd77L05M8okjYGsjukGNv4YbNJ9r/hz+qw84UJjAocmbRd2A
MDGklHWSnOy33d2fqLHZGiUOpCA6TIQTBVazwNoIgChCX8CX3hrCg4hiwQSxMHlh
xQc/N8CdoEyJjissIvrLYcWP5l09kYwPSDM58YbTQPoxy97/yQVhh9KS+0Fo/a0E
7c+rFWBspAi3ivWkSUsqN5cK4ahPtyP7RCrgw7wAPXoxQfIcdI3/Xvu4tmgP3gNG
wy8HRJ9fXj8AIoIGR7evygA9LfETBtxxY31gm3qOVmDntjapRq8cZhjIw60qwJBd
RJZ08v9389g3qYW1L9MpgN/488rxXqAFs0tveYkJwgTaopwCESsLECilHM4Lpzdc
zfSWfzt26sWZFcz89ELudFStAEHEEi6X8aDxit5xCQoRun4/8fDSgyoq8o+YWg8j
+CyqdSSvtapZNkbsFNsluVHtvTww27iXFI4Pj8SeEFip0CWUjVkcirDToIIDwV8e
5g54o3HRgr4yYXnStYRkk1hLCVyWHWOBUbYlU1MXCX3Humkn4Igu+yTCfSOxTXnh
VpJsUkkeIkU+3XuBLXFlMUGVKd0Kf8I48IE3EW8Dp/vGPlPhSRXh/xYSSPVmD+Gx
gugvao6Kszh+EjaIFOFYTfMt3XMIrgzZLwc4/cqufZt2HiVUi1jmPauPJiamgphs
fNr5kpFkKmWQhoQs7hPIoQprO8gTm6oG87Vyb+m/zUImtHNVIqSlbzxTLmIk/RvF
NoHytRYpJpjs5/amX+3spxtvE1lFIR/60NpYTC4Cd9YR8jGaqMFd6bqqs2BL66IE
D/lxXFY+7/fmstYU8A+UQpct5nVSSYu6MiQSDuCVZeBRlEHJDLIEBa2d73yqDcS5
5ASradWDfdSM92WdPjniDizIKpdtIr+fER3crT2QGxwn5ac5XFVop9MaP+v4rala
WOv9DAJvgU2g1qeN1r8RuiGfCJXKjgUizpMC84ZqRWM=
`protect END_PROTECTED
