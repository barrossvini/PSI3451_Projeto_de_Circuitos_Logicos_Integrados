`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9zWAEjrVR2zZOxOZkn7a39+1NKASm6g9jH13efKX2/FcMle3L0pPiBvuuG9BasLW
RgFDjrNLIwNxPSF7GMw8wS3dI9q0hrbnTmFMtuh3wpD+m2ERC0jIql24J55PRm99
prXNhSGPqFLab0HUavfABmGU14m8EKrCKdDeZLs7If2AO+EDGj+y/NjmlhGdQ6gB
9zM5de0/TbXxSrrYOCfepkNAoe3kF1Fs1890eeNLZmU42N1jX+OAN5hJkzRHuAyI
f7nUcy0uTcW/3xPWjht47jc+A4DqI7AcseSz4Icd9sxCuyier7bYsESRm4W3e0n+
7oNv37lTEG3htpIsEgK14O5JD/0KEEIUOGzgbVwRaPyVknJ10JSUIu0ZNPdteaDq
IX4ITnfJl1W6jnHWR6XSLOtA4Y4R69lB8vOYok6+lqZo4OLjh2mE7PxZszVNqCkW
TxpyBZR2a7jwkbu5/1xGex1f3kl7Eqv0gUjhyH5VjRAtO08xsU8BCq+1YbmNTrcW
ZlYz0oLqMYIw4dbbUUb6r1kiAi3dDxsctEDKjKuiH/jgD9JmtDP2OL7JQzL+fkmY
qAPmYBZqYSn9kTN8kFmsSA==
`protect END_PROTECTED
