`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cvi6hsbjK4Y4EZiKRI25UHW7/+Yy3Gcqp2BYKcjQd6A1UCyHH6chUMQNDJ8y/dEv
PyVfk3ElOp9EKwf2fpG8/CT5K8f1m/SR7nZgAqYW/D2OcpDY7j6vu/CVxILAoHbZ
/CFbPkKK/30GRS5yVMnT4I8g0BL4/u9awOyaJif86dcDaTqWJsgopgh4EPUzEbDz
xVm18CN+VWyeyC2RH5Hv74Gw1XhCWDyatyo7qp7hDuHI4JMXk8ZJd/tOdiU9jw9E
cxAvf0IuU5a0WE5y8xBFLVniF5sKgTUInyDQYEk0ZMvCLG/EjFQnixYvmqKB2SW/
8foWGNfNdgrfThwzxIF/FGFhjFcMbsa9NP+xdIZe+GzOOUP6TkpgA6vo1KFjrUFL
Gx/oDjL/Q7gJWyKAtn1UhpZKyNODMgAS8w50Mp/J3maUCy/yWC0meZRCXwB1LbRL
+qyasQK1q8nNvKGOb3rUHAf8KF2sAjfpZzFy3f8A366XKXMRJVe/0jrwGOkgveyP
3DbQFrngbi8GyTn8zCWX5927gB1oPTweFU1QFYKeLTPersmBZCYYQ4OGUYvGMfWW
qC5b3kwfa1mVqHsg7/2XuTP4uVCucHH05TnyF6b4cUvhUJDeiaXzpi4XX3sB0ido
wJ5H7/0ZF+SMFX7mGxwKIt3GzzNH6cfY5outsY/e6Mwtj+YEPvWMEDXvnpY/ouM9
Edlof7TdZVInVIoCKd3o4gnORRxBxcexTUQRSJz4LoGrhOmMJ6XkxCDsINGt0svR
ib1LbDbyaYCjy7N+yKdkXUGeheBvqkSdQytKOO64hHSvtmcJleQtWbJY+cV0JND8
Vbm+MZ9GrfoCw41Uuj1A/tymNG7qhpxTlkBRiBv9ycbxyN7ywCFhEA2rScB1b5qg
lwz5msUAgSvC+IvTBwkoHl/rLaiL7dBTbxE6D1KsgSye7Dxz0FatqvuR6sT8aosv
DgUstZ+PTMLf8i/nw0NThtBIsOpXIJbzq1/s+qusLsCX6IITcNyO27n4jZFRKNI2
NBhozKHop1JjebQVaobIe/MyD348Qr/eToi6RmALPflkhFp4KnLAgy2fLnRfJUZk
SpzU/5cW49C69CcfzCk4/QBBdTWVvbrjKVLX36uD4355Ef3/zcIWZc/Fp1uJoofR
BWzp9LcFhKlHSZZBfM1POo2nT6mwZgqMM0g64kP8s4aW8yX8VlfbP2+EQBQaN8aO
1TL3VxfO+jFQniqcRbUdZ1dUXKDFldwrm3RACrWOHLYMVjLxNN0VvhTmZ9RjGrTO
pfJ+tNWYkRKCN2a2MFwSemu6vLdJ54Ha3l/W9jics9OlTFvXZjbRwc6LtMA6Y63p
PYWz7dmot0PxJWyBXG3eGkor55vUyHrlbY9Zdw4DecIpmtAZRSSaij7fMKDJD+U2
ynrBKV9U7MgbRhdI8OyH87b6csJV4NkK1dnJxii0CTH30BEq4ecVkDG9e9JhoSsE
XDeOWehn/A75oEhTTnp5ndSk6KmJFccgJx2IEZaAvO3gR2auvzpcKRbWq/UGRKWE
MgVMv1pPQQadFaLeANCVn81gIHmPMiiIVyYJf+jNY8leWt8M9XpWMvDlohlsU/n5
aAe1yPsXZlLNZDRLRd71vKuLSBwmwHTHqut+SBhl43W3QCLUd7GMqKPgI8bZu2j4
tnqxPt9r7DtNUEhQubaIvfS4WShsJIVXUfjRI8dq23Q=
`protect END_PROTECTED
