`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ynamb2mu2cilLVPccGAUTFHWMrG6mfJ7XYhA53Tz977jKXZQz6kxytAzF058flBA
rjunEYELf23xwjK/73Jsy7RTP7GunTel0PQatkNH9A9bbhV643Vg068IuCvgyDpg
yihcbPUYwLanU3dqoPBRG56PozuWPGt7it8+zphy5jCj3V6zUlflAf0lTk31qwYI
ykXR93u2OxrDV4E8tP5lJA6ZZmQPZiXvPDXlhH31ThMgpNhJ4MIUmuaqaE7VAnlB
tfZP6rYJ2VfvRYeWFyPU2VSZHylhE55bi3qp7LKhCT1b9U1GqRmwIoGuAIScOA9B
hyOh9EPBv8+9XVS6kbTTiPdrQMdLBDfGd5LOUwr5YtCDFWN0IlHSvnezAdYBkY9w
w8uGKnU86AMZfYY/FfwYypr2IIO0bzzFP56g+fxiJJN79FaRkSBOX9oDyeupHrfK
jocUUzGNuDfKW8ZY3c/A1ww87PMWV+1MW2ZIxGIUndC4+yjl+HJyr1Q5/M6tRQ1y
s5IstnvsFqVMK8IwjQ5SFM9xrT0KSlowDz5Gr+xxGijYoaIUT+/CWwZjLAuxmFAA
DqOBFPSqaGlEOL2R2/rNP1VNJGKTKnxjQyKoxTutqxHLwCrCRPtqiTO79yXdYJnk
mAHWzMSnZlDeW9TIJvAqXm2kAE0C9bbx6bKPVBRcoaUtt5UMrmPZgNhCHDYNKFCs
tdO9ZdSBBvCTn33X3eYoZ1SBC/EAr2NXRxqnfIPl/3ltLamLy4PpAVWx49VFtQ+M
Sahe5fsefpng5fVS33+rJZGmsAhd7Dwuwhkaas1FcWFyDS8OzvGaO04pBWWrCXL9
3yHxtagGzo8hipj+3mmp3HfyRUnTYR+4k+0gP5qlIN/+0WqZt7AZyvBdF2ISqsZS
e2L6oGJt2DmAHMLvby8/4n+jXp8AtRH2PAMrxULH7pVliipJxnJF3ogfg4gZ0Ihm
t/oUmMlZF97W4Oor+PKC0PyGXhAueAKuOt5Kg+Qjaq9vZeOl8VEPW7gjX+APkLMV
80j9oDVusRdYEF7J0d0mJaDuDLtbjJ257yh/K3qaz3xMRvRy5Km2EFNiFVusHFMU
DYVY9vqWUXZsu/U0LRdX+0/IeP5bfGa3z44Oe6UXesO3Gd68fWLFKc0+ONPhD41Z
yef/KzsoEcp1FllRE0wfb3/x9KEXGdpn6P+iMB0EW2usyihQwutPrNs2le+VwEz/
b5vE+NHx9TYu18O60uZtv+4gCzZF2O9xQnZZJ2b7YkNxQWSkLN4ozOSQa0sbN1hQ
giveUVYcEJiXBCrMp9MMrxPWQrlFO4Y1QwexO26SlJxDzcPkhHqFLC09usY6+xqK
0o5q4935XMZQ2tDHHJpgw9dT0j0W78SBbnz+f9/X8KXC4GIlbWrCEpLoXr1bCgwo
2cc8mtiU4GxM/uxbXrOATtjI/TqoTD4nxvPCYE+VNUlPP+vUQ5dpR63LeKnhIBt4
rxvpQ8D9obUkcTxoJOjta5FDg7rFLjgoYlyCQViZqUzIJNS3arNEbpXkPXMIsHd+
fe9Xb8Sgn9VoBIHQvrMjlzwSg3oP3sAxz73etatPjt9tSWsqI5iM8UHvnrF2xdVF
PFnRyTikFc8Lm9q0PZgONY33L8M4f6yRLnJ7T3iV2ePN/rBOMDTKfKUQVtwVkPYx
ETqSZ0f8C4wiBwl9qT30LE8DfNS/WoYTvUnlXLf5boaUUHMsoxtx1SCrElkVu8Si
4ZOOrrXZ9Mt25I2EtndA+lu0FlQVkEQtKM43F3O4Ip1hsxdEOeCRxUPLDVKMkM8u
bSV6jlA1gbB3ov6efIDMjGW++kcnEKuREcbWzYxJ8/xnFj3pzvbomO0TszY2LRlw
YVQTXxDQfob0wt1sLwotKJRAgX5ao/CvuPs59AegSTiO46rigowF76hJtLrPGvN6
yZEFDdcOM39/v5Aui9hawznb14PMZlAloFttDx5EDFk43oxarfOofvTiix2GSqHN
sPqDHp1ezwnVxskmVWdyw7ymqh04X/WK6orOSFxKMkiZxIAkXAQwvc9C476z+AEc
oYjY4Jke5ED9/AcMrz0TqaUEhQpA6lVWF6po0erXi2sfRLfny7+656dRh62h+0vB
ROrRFepWTBBw27KiyKn1MvbsZwQibw5/6JTVY4XPiLXR2lJCwWJWbt72m0/XA9Yx
jlsp2ULzEM4rBcrallokKv8yTBlJumx1pxhKT0wzAE0v9c/s8c53zf/leJpoFo44
OG/ggJ1OlFb32NANWy7qI+qfzfJ7sq7alpzwNBCUtzzU4bbvSEqHYu5c5PxMt9Fi
TMGUHDDWTVe5XrfAE8KZrFSFdEepTdgxl6T5EIzbROaJUa/UJxLv4nFrlqLcKyRH
dPJd29tcgdL8clMNRCWsJ23ENbFpesN5eynkbv/NyHGeKyX2af6XzEYa8oOP3dpZ
73mv8UMcn/dKiLUm8OzDLsNFwMumskSTelL1TsBEV+UKWdLlpw0OEtw+oUgdbuS2
WARb3LHa+eyTsj905tElfHuJU4Lvhrw8LZqQXsC9JRmQBU0tWf3hVg3qiNeu9Vlj
fMZFS499CqdNbVtCQ/9CKjpCcr/AkKFlRXll6u3QzIYWag0Qboi9DZhT37P4DDVo
lmYtKUEF2bOoEn2ppuy6PAwoTDYi26kqZzDo8w0Fj1crHmWcmGiU258/RObH8pkR
Av+vecwtSBcwWh7MTN8wH4LICFE5RD4nM970lqvTwK7v/jFa+ZEPJa66twDOj/C/
7FF9/l3mZ58aAjCl297Xt2FzWqDHUhFGcAr/e3PwXxcfRe6r5yFXV3KLCo2XbI9t
7F2mVCk+T01JSKuo2wrFytukH8E7edGDcKYTdly9yjdAsrxQPjU1/YWXpBOnryMO
APyEUoI45r8iwoBNIOa2YaXdlgjYhuIcj3vX19UjjLG9geF4+ztr1DJEkOvtVWns
OSvs9T3PWCTRwFLgT/euNSktxzVYvmfcLofyVmna1wPm6n0hTUAHsHTlICvQ6/QF
bJ3Bpotg4QNL0uI8ozwdAc3b2IRGC+APXmePmBH/eKFVe3BUFVkHt61CvLys4XRK
uUYLJi9il6IznRW0np+oCU7H7k9ijGxHcjxxA041BubdjK8cdGlOWSk1O3mZOWJA
PLq5MvDukncYWcXB1R8uzCwPoblFdLeoRgIsU66jKaM+mXh5ECdH9+DVl0dkV8Sz
ota5jk7O3esSVRswf2Tg+/QDluOfMBnCF8IQx18DgRmOJEhBGSlF2y3JmVgw5Qh1
Mgp49yqqqzpIPRE/IlMXd78iX3isGjWWu6Q4sRxPPjjsjO6V8PgyrvtnCX35k7fc
j3Sndjb14h1Nc7h8zOd3AZCoikkhf3APHTSxn1xdsOrV4SEy0xOJfmm3Nt1QjkyR
HTWZXc3wuyTL/EyuzG63gw0aATKIbpt2MahA94YZfaPc2EEFV8MCHOVQHl1Mc4Ve
c8s/XsOsJJJssPIxdDRsate3HMjrwiHjZRDxWT8ra1bytiQAhscbP/p45JV3rAHP
G8BfQ+Swvkd1caryr2uMhUH3NveLj+tH+z5X+61ClqROL/ijmau1/JyUFfHza1mP
J/oNARs8hLOfEhCwP3K/RfYFolEhciMKcnRQpJJGxftlECDN3eGKo7NtBBy9WON5
9HsEHfDVnWvZBnQ1DJa9ubE3tWcDiYJ3OeLALTrPF/eFQYtTNcqejUZ29Uj8BjLg
CEprCOkrwgUhneGBA39SbBseZKoinkkzNeOvmx7F+6vIwuph8qacEaFNYD0UwDaC
xtKZdOQL/5gIUEdKfX7YSeqhdzeHScDIQ7izs+gTurDwO0ZrzpP4DclW75Tq4L5G
NKqreo90H1oK7M+dhvL78T5ddQY3p2mFIuqbIi8JLjmQGGHNWVX6qV17l6NzCzUy
XjsSzuh7yccKFr/Sl38hvUDbtZhB/B0QG9kOi0eeJnJWNCex5jv2hxLn0Xh0+S25
FI7fKqNntjOmXowpEAI6vYcOy77FOVeUrOSOXM86qAzCdDI177cIamcwclu+9ZV/
AnJuRixK89dCzxtuOJsRvqkqfsn662Lyw2+IBHdqGl4PzfvsAAHwEZ+i6v98S6sD
Ce+EELGkjsU4Qa8quU6fQNCw5xMTyviVfiKBF3F6HQCnWcUqmv6dPCiIbblBSTq0
5f2UzffmBxVCBEbeYh5kSayInjaj115N2GUYrDhWxJ39jkp+iqkuD/8S3TahFMqV
F6xocfGffk3LrRncA4AgaMzkKl66vVIxn1XhM8UGfirJhBxalRWGpLWmqn8G43dk
T/3Wn5+gzTzt3HYKKuXlpbK7qjEa/vr3r8ngwbwpHurjt48kqRWtVOrtuWX2QdaI
WMEizs5zWUWwx1VnqCoi+KvkATYSWYZCr+iI59oNK93jiNIxvC3L0iUXpLQAEw31
XUjOia4H1POigfX7wAI6j3ITpqLyLLKhJUfeaCggbL4FRoMZIWwWdXqFoOSrNrI0
DFEUcEm/sHS5XRMChq5iHFKrDjecJsI6wXhi0jDpUhtS+la/knABPOpAzXIND7fM
GILkG5KNyKmeUegMWvt/Q8iAmHvp5m8anD/wCeoc+VMjBiY6au6f54/xq9q775N9
kqsht34i8+y/08KGnPB27hInmENHvyvCOEarEgtoTQ4ey0lXyaPrdaj/DosmeE1i
67++WmT7ZZZBYJTBB/bx512GjXVU+lXtfcD/KK+dEL01D7HA6KEpO27iJb2fcB5g
qCaeZSSiStaaTAQQsGzidKQNrlwDmsfJpJISEoBy35m04VEwIGone7AE5P9J6aRV
9jTDPp5xuyoxb8xd1nG4BZ8z3SWJHTRNpsuIuD/LARJA8cF0yrgJ75/tEl7xW2Px
7ZnCCsKfF27U6ZKxk6n8bvPN+tCfERxfhl9GMrTakr+YywdhoAUWntS1s9QuA4CD
/nBSaNamj9p0/CM8nm1q+ArkmrWyd7MIfYB1m0wpP813S7IGCAxvuOyhG1A78aH4
GrE1QRXv8REbfMjUS74l2DZ38Hg+HErNmiwuQQxFmtNIAS0c5zkaIjfRWp1CQmd1
3wFLuC/y5qitAcudh3zyQw6woRIF4DzLc6hgv2R/6LcA31O8lisSWw322MTZhbv6
6yX6q96Uvhxe3UOVcxYsoIlX3q0KAEW6g7u+ca7ubfE8JNkjKmJPrbpRDFmaB/TC
gsLvK+kbx0Z/3sj6qcrXyeViM5+8daY+2Fp40hOcfgfj41oNSIGjL8qpizzTGSHt
S7y5C7UoDY8HMrt+ahX7TLCcRVU3I2BZ5GKtUDYaWh5h8oHx7SAavK0Mo+005nt9
tsaxWcix3ox4m1vzDIzKqT+vIF3Hpl1wlEbIZx0FyRU7GbwD9wqdvNBfgYZpTBaW
lmDRn7+QRe48EoU0M/nryuWUGUiQPP/maRimcwcHfidL+SEoG+YpReOhFKpou13e
QRD5D7k6iXzmh6y9Szr5NXzLkTYB/u41GLTn/uDOzySzlr4GgBiyYAVuhwmHB45v
MgS9V+6LOHuB6VFzaUYxtcS93hDHK8JjlkUhJyf0AKEWSafGj7/+Nefu7Lrx9/aX
5kTdPD1L/iTJJ055iv11ozV6trmpskRGiyCLZQGt/iFm+O8b+oi6n1BEOg9cDpXc
CE6ADc0bJsg0PoBWURlk4yIdjlQVdecwZDm7bLJrcgeQI++WmBrmTN8Y5tSUsPph
iFW91aXOjJACwTsil3kou8p8S8aQLBsFu73FqozfmxrPIyaMNo/a3HvMBjyTEbOv
spxvuUudea9LPxmNJBNXjwGA4yNu3YU3B9E/FJVXEsNPw8gfdRSZRxAjkDKN11hA
P5n3c08kHtPFR6Rpztg8t7DyaGeebAdmjZve2/TUkfR5IYS885ThG0s2noCFq3lM
Dx0hmcVVZFV95GctTBXUH+vlvEmc6XcuFLc2/YlZyi02uCYu8xGAnlYqps0DKAw0
DxDCkyWveZQKymHVmuK1mRnuSB6/+phaqj724QjRn4PGcFMnAa+nUJZZxgzjaOQ7
Y6FNpLCzs19Se8zlXXoQCBGnOPuqmDyfcYtv+22DslanIUp18JY2iEACyauR0xMP
M0NJvquepHIl3Fjqo5BSBUKTgzihynBVMSCmdhyBjsUOi/5DtbPfoU8b1tDlKjD9
Gcjuk2/piTIt0s5dil09Cia8iximObpKGKq66B+/xzMei6w1IAgEgbDPQx87SwZ8
G6GOtVck9VBF4X117cWkVmQES59gemozQpKJM8BQZKLMDvvbZp5Kcx95csWT3Xgx
sl2XkaXOLRTVEQaUJkESEfYl2WYNjybD0sPxgEjiZWMLB+Tc57sC3oYjKCrAs7gp
+spgWTWf46aQO7KB+wKDNIxjP+jPJ3D6gFgpqYaUqqpkIbo2L50h48EPulibfS9z
whLFGwe3BIpf7EfCDSiFAcZ5iKNfFy6W2sBiwg+A9ZMccpwzdNst5FCPRlqIKjiW
FyXgGsc4BKNNygJWGGv70wpx53S3ecpaJXwKuqTKy7ME+2yHNGJLVVBL4t6oioq+
wDYcw/ZJkGzDcH5FS/JGHocfGNq21vjpEmW3CvqdztGIjjO7wBSsjYUjyltwCnot
OQ8a7aCRcjYzW1Rprsfw7MuJsfLO3ZVWaFsys3IrLo0co4QT+ughSwxbuZyS2shq
YDXJDsspkbpMEjV8X3lSlDOgi6Z3HmQoTfhEpY1Ppxl6Y4h8sHyhUFLYKjQXn645
f4Gle9xpRSYK4JB6NPacJ6vs+sPZETuwkly4ki174rjqobSh/dEndrDXYxwnCVMY
LuRVQMjJ8lyY55NoaRpsh/xqZPdlCvqbpCIgb52k5zamp3btjNBo8CB2g+mksat3
E+7CgHOWMa6rbdkm+HyLMhuWadreEZwfkdEpWCDeP1NpexcdagRVfqpRnLTDJnAs
JyrUjhw5ZxwnaXLqNHE2m60aDgLjBvA+X9x846F8SlY4SlM76kwnbCulPHpxnyWp
yu5Muzi+5M60Iw+LsxzcTBbiuRdx0EqWZDU0IOdeUXNO9eAt96RV/W03/5v+npVT
JvbA0tSogGDhMw2nFiXCM0rlJuQM3c0DfcCqeiqcF5F45LiSMqNFmN/mkW7XvED0
BGIYn9PnR1lr0lJuxOreSrBzuf1B9ztGtWYdgwrevk0o6PO6d8HMA9osAUOvyfNA
1t21KOahUMI5KAQHd4D66Um6iASAQyrhvKHppz7Uh6TWvLHj12Qza6S6hCKwFbgc
Nh99tvJnfFkm6S4Kf+6/N/M/gTBM5FbR894h+nGj+a6OKjg4GGpBBgbFoVnKO0Pi
/gWHh53uDqKbh4fKbxazAzESKQT+qh4urDmmnpgw7PeBkcKfjFNBBNO7dsKkmiCD
dn9O3BsEzOpJ6/N5uxVEOsLzHFejL7iw2630RiVOOWOH5SkRsEgMkoHv2UiHLecW
S+QaWdHMn+5Mb1upZc8bp3pess8Dbo9oyDN8oNpinTj7M2SGhlBUiWwLmoib4bYb
ScMvyR+74E5QJJTmZXDFaT7JmXs2By0zZ4o/sbEywgKDuq+3OVN767KISftU8wAr
/840xA5OavXO3g4SoE8deHX9ohsE/N4q1RaSOZ4eSXkSjwv9DMdlLTUTyr7U4S/Q
2cG7PU3A4Fsv29eJ9ULuvMMPGx8a3T6BPX5F2/hRRPEx4Dy9eKGe7q3IdoXx6szK
jca+Ta6qcLyehHdcwZL9SQUTg/amYdZEx3HNDv418+XTEXx00XC5vv37MxkhW1Ay
c+P/PeSbfNqdvw6R1oEVQsQOrEx1T9/pySi+cefA47sZK6pa+rosj38z6ShVz2YA
U4pwrDnsEsOgPmO7sEb48qJRw/VLYSgJi3N66EyROT9V1i8eV4LWl7GKo/Z1gvQT
y++TYC11z1Ip6n49/kWiXvQPyT91MKy6YBTTru2nAFAgLvW203xZbH97/Wda1taD
a+R3MrWBhpq6JKICCrC4pGuHcYL4fEjyJ2dkpvcf1liP1gyuEqjDa2jeZznHq1As
mojoRexcrPRBBKmo9UfMZmbsy/bjRTe0ayvU9PJPW5+2JxeSJ+XcoetfOcFfbM4g
xYPlybFNMUyqzJRkAWtkMe+IjemU9fOCQ5ByeMZWw1RE+tvNNrw71fQiS3z1o9zJ
7KcOVqUFBlhj8DHNhAwLhkYhOf8Q16+qoh6q3c4G9UL6Tx556ZlUrH6pFSL9oy8V
GdEFfNS27ZgDHsmg+aAZkNGbhdKXC+3hMx5aKzvV+Oc+pxbqUKLU1mwJmzlMcGLw
R/M+ZKBPEMrNRhI3tURdVvPm2JSuxnPdgGGiccWLCX0FLbZf5Q3Fh+kcy5JLURDO
VMVk31l5zhMMCytW8RQS6wxiYg1MGPv+C5+Y6KLvzKUdXW1c2XvtQeoykLyGiuUP
YX/MRgmhP4Wj8Yplqi+uojtL28NmZUwkIi1zVijZkyePQMBNKryKjw2BJITf3E7b
AAxPMHpLT+VS14rgNMsWV+jpQLycZsuEnhpeSCyxfDDY58ITg3X6AW8UM8Kw0bSB
/4vycHR8dY8isP5omr6K2tWfUvQ/EfEDhwEeLI0UUjWTYsZuWPkhe/bA8My3IXGQ
NN6Vkrsv3Y926Vtoco6fMP1cNtj9ugTDSVF5LACFGV0S4cIsr52H+/DDdWqCns8A
a4TF6J70X++o0fRRq7mT6bUIHKeX032psMpK8bJQMOudDJ+2tuIMLT8Badn62+80
EiIGFX3zrRzmdA2h5XEjl2vH3lkE2C1hjHEo2QttayawCUfTBjD3sYMgzvC6+c3r
59Jjz0+y642liwY+GgXzRJAQzjs+McqzBc7pXK3F6ZximBvQWezSMA2xXrrhDD8r
WZLW1z1Bzmn8rRUkmBBTQ36KdRsaBb1iuL9Ni9Ii4fSE9Em/aUsEPvKS/i//p1P3
0HY2+2nJLOOvt8k54uZXXimwPYNVx+l1Ln8jb77Xi/ojvZU5It/V8of9o2Ugh8MQ
4f4ciqHdac8lKjIcSz9OYzGQJp9jZk4DfbUZu4Zzt61IlRn8IVuBVo/dIAmCFfGw
pbOuBqCOtV7pmiLtPYa3zIBjIM7m/mjZX3WPwgv73sC5XMezGL36Dm9FMLmSWJ27
LjzmwB+4+dRtGbJjeSoMwvk/4uCKjZzUhkpNOygSnawncnHGYd1NXrWxnc43dU2u
gOWzG+U2asv2EerGHcqujzhmQNGI0y7FGMpN/ZsitWdN3f6kCGn9YMMO9waRaBis
NrhlhEP4CbhGl0aluv6uOdWJm2fIn/zI+rNry++t0+7cJDNX8QA+BVJ18dfHtxbl
UlaccsX4kX/FuO4pdTVGiCebBpzn2352JoecrzBr16BsMEiNK8pOJTfMn4U7dano
xsGCmp00SWo6jnlTBK6BF1BsPcJdPy9ot0WhUywO+La5lgnXKPs1fuYQ+iDSRWv2
7l9NZTlFLCvcrfYoYxwTMfu6L1dg50WmDpr16I9EaWnEChfsWJvlbCXde8cl56FN
cjsxTLY4vvXJW6GNN2662CZYpPJy2r+x3wOAzvbO3zJpyNmH74cn0DHrevu45GuO
mYVoVm6fPmLr6tyQsuVZMA9amOob1uELruTr0iCBUJMYfjxU+L9SUit20dUrqbZ9
1ai6HxSUA6dsdYZknWg75jDxZfLTMpd/wNIi1gKftnWtSQNAzNV3XRZdYzEGvZGd
ilVHl8yANjD6rh0pJvf/vQH/B+gTTPwjIJPuyqAojaI/aZl5XXSW/Exa0v4jJe1Q
WJFaSLmEQtENQbEKY4avE0pc8lVjzTo4wcX3qR5wtUowqZFSoai9ae/SzG/Km48t
+lBKJfVWGCNuSW2MTRFn1Li9V8g/VN/iXN/Gk0+I1HbozbUZhadugvKwgEsDt+Yd
4RiIehrcqsTGty0RukC6S5lBdj0zK6nTzEuzsm/6Ah343Na20N9AHh73hy7Yi08c
IFAq1vQx90h+YV7anzovbs/daJT0k0t93XFUQk6ZZic5c5CXdUhaNyYoKDuN/Qr1
N7gWj/Bei22LYpGoKHgblPWoWTG4mIW1zMV3DdjcQZU0+xcNPyGmLGKRLi959l3c
QGrAiRmdqj2mIvSU0Rr+UXWxVsoQmQxzwR6iJSjnOmcM++eeC8DcljBBf//Jt5Li
lR9hv0sgM5PKkLhTnE0roGlGn6Uf2CXotUITWyigmCQQ3IMtRBd2mJZvSV54ECJo
+0hMJ/fYhl4gGv99b3XT2cGUOabKe6pQHzDb2NtCQ8GSaY9UelAVhtVl6iQu4mOr
WoDZ1h9KpmyNVntTi39u91LuW7RTvfE33Wz7/5tZ6OKnKUNzreuUSo5iedKg9Mkm
V+4qFYK54DN5HRWyM0b2KAxrz2fnTIWXf6DV5+jL74BYamE2siapDQssotubqVZ+
pkuH0nV28DrL9c+22HOERE2YVctTVsIlpGnyaE9NAWWhB2pNHvENIG+lMSSiru6U
H8YVZkY+UKBKSWohpY83IPIkwqLC2RRG6M0/AXXzvrG30PXgxpBKvvwwVU+Yi2Q6
vo/fYoX6BLFm0WaY3xgSi8eMnc3ii6z+yYxTvDhebrgy5l3MktiWBaFV4x6II72k
9C5ubBXylw1Q+h0pgpZcysQOtNCfo8R+jJne6zzwKBVdhwUi1L7+VxB5ffyHNZKt
x7ybnZUeJVj0TujIAsHOvBaDnWu+6jNEoGEqxiCKaes8HEByHcwh0zXxCXOqXnht
GgqYdkezyfODBiCWo1dg8/SNB+qXkFn3t1+JCcgCy7J6KGcwhTefdMcbSmJYWkCS
Vzgaa/1RuL/bN0HgVjtIjsjWeu0+z7JhKQRhZZde6pekVT9QtWZgjxDw5oDMVYjU
ZjaAdm9ebxHPivbLS6f8Ab8MHRa62js3UwpgSqqN7k8idPjCEDMDef/u47SmKb4r
s4++Db4BizDUduvazXUfeHFZfqIKkeORf29icgZl4vS5QeNRnCRcYFalC4Ua6Yf3
+lFMy9x+ynHT1LsAotXzzre+s1caqeiKFxcAekkUchTUMnbOFXshJNigo3TKKZJL
QkwtBvhoOL1qlw5mnZJuULj5KbKmUBJMoSXl+XqjXaZrQOmyYRzySOh3rhU20MYa
WVrqCHN9VBqBFMm736/OQ08Ksna70a+nu0Cd12eXc5Y2Kuw1FQJRO0j92yhE8599
X3Ya3kYbPJgR5WYECUJLSv6CVn3cvZ+yXiuBzdx8w0nnSspsoz33WkEtLS5wCD/v
JKZ6VPb/9krdG61rTazboO3KPuocQvwu61/LQOWXjralrso5JFwCe1Ic5tqY+nIN
J2bS9Yg+0EbdM6oWRbQDnDbcVxmELUyAc03WwwUeEB2LJ6oVCEz/YTKX6TmfbF5u
Zh7WmJ03xFcy+uX+9fdfqsszZVObgcDm+qval3/TLW+Y8wxohEO1vN47yM9LIlaf
DrOOCx78AF6+B6iuuIsnfQt8MntHxHUXQh4ZOhgygDB1dgC4WJfHlMO8O8hQGS62
csQ7TkPzWLNM5Wt5E6OalgZrbLGKTGDQzwulKEu1a29l4GY2aOR8ILGhmgrsw0y9
xIgp7fT07lAnZlLfI2ACuU87PeX8dzDas0GldhT9CoaW96aAvWg3SAIJS06t5L/9
S8T1IRJG2eI8/+9mb/RSSTdniU59xvsV6aOn6zwxa55zUC0V64yyjeKpl0CYpsBg
14t2UcGfxNebDbzeZ0SDvP9t8wQoTNNCR/QXTWYbGUodaLv3x1Zi6klz/3V2kn2Z
rGwr68uzzjInvmgQSe+P1pmfEGRkoxSXBySsFgGTA6AEK2D+D2szjkM0PSo4M0Mt
kchrhzu2X1VoD4mfRE4CnbFMtjpa20XsdcGNmFiEH8hB8hYBZOeEGcdC+yCO6M0d
2r9njzI04EuW9xBd3GEaMTwRJSwQUXqfUpRtGHqRyL7usd2L6+FuAuYaiMkZ+cvq
+31zwXMtApTVMNI4Rj9VvN9YxArEg3N1TthaYLoZmTopOgzGeKQQ/ArEYWexcc2m
xeHG2Q4vEfJeL9g224Al4d1YedJ4N2V8qqbZkEO0gXB8ZY45XqO61MhKy/7CIy6v
Lmp27J112q8s00R64P1G1BniuiOpg/ynesyKhGOuwmhrLTSNfpRDL2mIBX7UViht
g5gfhOtn7msuG3Fm+4hvA4f+MVuhCb1R1v0v6/8Cn1SSNH1H4igNqwJsfZZq/Wyr
4/KNjjR4NNYP47v8MU+6hN4fxaFp0SNZihGNoAqzV/JNPLJeDZzMre7JgdUXAZNp
3uUHq8EmuBEr2r/oQq5t7WgceeeaRep+reQW7P3q+Q3Ms8bkRKN6oNuRgECmszHP
701RO1iHzI35J6c307722PyemssAZUE0ktXOnaGYSBoauQqv0bH/bqEuRn9injfx
Zxz1VvF/YAB1gBMYVHkqgQeGEVITRKiNSXDWxLWFj0SJ0aZ3ybabQb/O6Gax54/I
kAn0IS9XIrg0ef3tzLZg/JS1QOWgqjd3ApQIMAVsA6W1Tcw8Jr5szRDXJPLa/dDg
gTSQbvE7LP1tPo49ew3rV0b2O/uZ8vAlvcZuWH61IxBwONGswOMKEps0AHuAIKKD
trZ3Rp+RrwRPZGmnKluGz2fVrAniVfML8cJWWTrGw3GwLV8PrlotJyFgR4R2SFkc
ubsHkHSSoQ10i7NCajlvb6v/rY9fmwyZdeFThpq4Pq86uXuAEDgqas83qUPFj7/Y
gcON5sIl+kSnjkmozBaxJT3GUjNoZbTzVKPdNTLVOn4h/z1ZbmPM95jUmFMpPNEo
H5j2WHqAwiCPgwn6Wmw6ni2q62JBBbYXqvoYBE6jSjUrThFEqt08WTAsbQYCtnCy
UAuI857By+grveuPPL5XT5taD5QhHU0vIFsuOAmvGHm+nPLvMOpmVnzqc74JPXap
bh10uHNNaBXur4z0QRR2npITd0D3LJwJ8dD+bbLqsmeAe0SOnw3G7Z1e4f+oZxRs
ri/Skn+RYc/xPf8ZZBFKsFtLLih5CtaSn2R12tNMFerpLWb0gsMMgcFoSaOJ9mLO
qbxD+LiTCdkovvx2t99zbVYEvj49Gtr4TcvPHXYkrt5hLrbzAV8rQhlLRiWw6uEf
+XQvyDwbqvDMNmFzjgC5lccUcr3CAY3ffKTs7NwSyA5ScYH9lfeTGiZZaJUN67rP
SNo63Owz9O+kGs0cq8xPCOuVwYQfPKBbgt0+GxrYSrEDxBGQfxKviMhFJK7sBduW
Gd3wFSNelIkOCDKb3/O9i22xa6Qn3vN6h3DDHMR5+2BdzyfG2ekfmqz+YJm3dLCV
vDIBIMija5I3jZD1I2sMNByIKsJk8eyUJvg9jOSqbwjh2VfsRAmk/V6KbcRMJ9qj
tR1A9vWeCEh5TIzL5h06c2wti+9XEoZ77z4KeAiHuDBYRa5iGcccxyrJFumAlgy5
AY/pFXwvzrtHqBzky4EZIpqomEjNE+Ikfe37iSPUWciIyDwneirmV9xb22U5crq9
VZJzPpt2BwhOhWr8mqnOnHaUISKsjOrSXEPRfxiC2FlCjQP49daqHbGhuPtMwKdk
4Mm0O8YHLhAXhv/NKNQODETFV+dn6PsUuRZc1py1lFy2QKjYMnfkqxiND0Xo16KU
/yT1p3BdGktdEa69Vwy0EVMJQCmfTNqHBO7MhfalUUzCjmdSzjgndN/W4lb+he0X
MmmIIPuhsJ4t8VNTH7eteZgss/NLbk3tiNaMSgBgExq2prHMLHA1z+T+5A6hnnIS
JWgL697DBy+YuyMghcyITFAKbA3zidps5vRPRIU8pqhECiU6Ox8qWq2dI5Aka8CN
KslV/gAOuSDpM7L8wnHoDWDhTnK88+H6NqEZLpYe+6Gh9f3GjE5/zrR1l0ougJga
jKOxpFi6hbTcwflq35TVOlFvv95WPY+YVwK12o5923zu8L8kP8PXpT6MWPtzhxp3
A+3krzLm0wPH34FqIUU9S8n0NumnP9z7vnhHR8k6JVZwAkrDp2ozG4RPd8vsGKra
4yCLcC6ZGmHMIufPfiK7Htq35N8LzFFTslu+IYUJlUL8jZKRD94yBYVMuv+ab0RR
Zyh5kmHJslxpRDa8SzqM/bO7bK92SoUYYVfg1xdT9SCFOLe90HuN4tV0tRtygRGa
Nx1ImFtWk23pB7TMgNnQjlJ8hc4ddN7CCbxxi9clJoLBYy9t/b20thCYcoxo7qEV
42C2CjHdW3nWCs35vOj0CH7YJzA/8KuXiFOul79xBFUX1lzXaPfivQi/77TySSxd
aTFY4t0a+AVhss/ebO60g0OYxMkl2nAV8PhjPWaKtxx6oeqEsZbrSpHFy6qG6T4n
H/eQIQQnnhIH7W6P1nog0JTFFJbVsnENu/ooLnyQnfh8Pzg0DawE22whU9c5oxsv
0RKk3RwoPxL2tWFZgmJrnF1EbShT1I16t+LSMH7a1yCEUVqy9cyZu/3U2pniW4tq
0/GC8tNW1CynahabZRv5V2VmnLLJOfTagxnHT9zxYpnUV/dtMhQfoRpJCZbKo8Vq
1QxRjcWgK099fsca2Ge4x7q+we4gpHb6IwhpLE1mjLKg75jzN4EQqPJ6K1YsZugX
5akyhtp5DbBuiDQ2T4o8V+AV/oWMigB/upFYHEz6PMTvwtenEL6y+M5kTLGHG7jI
GT+9wnusu0mFOkjAAvV59vhA5iy/OLOXCA7RCJpgOurB+UCZTYfKWjevuRGwSHjA
Zv7Pc+PYp0fbo+h6GRgY302L4sH1CnjpcxMnU3ItVF3eZcBrSy3PNQ+fIH6kXicU
txUEfaF0fHxilA/1rCrRUkQBysrwictsxd7QYp9WdaD5ixzjEGagpsZcSJGeelRL
FzfQ44TLZJb0xE9CGOwYHDFhbKToVxjN1KkS2nUt5TSn+04Ig2MkWejDFJW9BG3B
3DiLxq+GGqOovJyanmBqQn3MDmW8ETR/D4p3Xfc+IP9m9wgUm+P0KAzLB74D4Duv
4sbTZaBA10vJH9ALt013GzkTLEtxtiGcV8AjbkM/kMmgkwQpe8ZWX4f/7/bW5uuZ
v16lFpOY3EGrxOBIJdxsW2mDG51XYHX8/tXLZM419poOxePlKjf8BrkcDWaI8vO+
Mt9FDzqwWl+4AQRZQd4WtRXjiEbBqLUXW4nesmus3G0sX0W/NWNpH4PtpX7+ri1/
EGtc6EFPJ3AAjKB48MpzNDu1oK8xexYJilKPY6yntKq/omt1LGeEH/K2J/wrxqZP
0wE70w2V+1RjE5I49dLRTmiwGrgJDhUapWKeAQ7ZRkyu47HnVHVuNF1vKhKncvhb
VWoZkPaUT3cwqSX7vw9nSz+qoFmTYhSrN9giASBZMEMfCBveMvbuH4wFKpDugZWN
vhPxIsVltAGiS403QbFLAvpWLf+OCnw6LJO+oSxlNrDpy5N+lwOjC7L4J77c+GZt
5V0cAG9NivF369mOLyJQoIXDd+m5zbaHmj2lgXWkR8d61eewVUMpmZjSS2PSX4N9
pBbWaTQRjklDrvp57XoNSVKQei9Yq9AdPQw0lVSv49v9Jx5+K7pdbstHZXETnBa1
RoNsm9OpyfM0AOiFCxGk/2Oh41yyyQegUZ5fqcFBcMmEst8/TMTsB1F3zjH1oZX4
NleWPZ6zPS5bsMwxlPXtOnkYbM/OHd9Gpgu/2P+p9/Qg4Tka8ulbuiAT4Y6pzpFN
h3ZtAduyarVKeFLHMezPYCcS6CwYTRmAhUMEiYdi58jkohhOIhtk4eb0iUGUAgxw
eTvi+9aOkpmx2jRkOHygdzr5UBlH+WTyDxydkDCRC/F+OeaarB0pgJ0QKFk+0g4R
LsertY5RbDcJUat8jqEaW9iJcaojkw2Y8m4w1zVmwVg+GCa45TAbxMHxILCkI8YY
6jCEoKfYuDEvrJ4eUBCBNe5cjrjIS04mtelHfl4+Jnwb7KJpc3NPiWz8fv1pt61C
E8Hd7R/8KUak1CY07OtMgIdIADZgrRC2VCmuT/E5WRkwclykY5CYPNGKPO/B71wF
MsLgq3NIRCTBB8pftNEQXjg1YtYtaY1Axwxnu65bLAzCrTGXiSwOeN3leNTo+J5Q
fOTilFqTwEd+wuZxqF0fqLO4fLT5fxSKMGJpbPLwTm9/PMIREoszTBZ6V2dHqsZS
tzLC/1cvXRu3dt+PpyxBaOL35aIm4/wIcgK2ClXcX6a19GGzu3gEEYHcwXK4ErTh
2zpNGnZzOU5aW+T8amKeq0O62lEcR/saqAzJywVKHJbxblbVwlxgUsTHH2t85ISM
HGr8h+gqZ6xAExYoT954YCHchrQUA+sOb4kku028e9Wq6EsuRVT7uB6h6+RNUGXX
BTGI9BDClctX2cFiGeqGY388w8I/pG35C7YcN98MyzhT6WCBs5nGriGcImEKxKCD
MnVyu6YR2jqVDrHYRCRE6C8wgWA9w1HnMKKKz2B1hbbA1mc7ONFfpdq3957j2K5f
7urd96Xh0Ajq1zjlCYH2JjhaxJOeeTbvc8mbtppxm1aRaoF64QeWT8MGh0BAFPJT
mkm1umv6DgbCqtlp5SnCZTd58xEdsmyrXqksleoIOGHh3fRA1z4bXxjPof/eBZ/n
wplb7r3oKOVKQBNufrDarpG0lxk+hOl12tFrs2Sw+PWfSAwlAfr1FnLe7EbyU01U
FrTCZGwiQ0HVE+/Dj+ptNPwRiAtdm/axoqMJIRmkGMzXMEFzah19c13vYMRjtktT
r83ufppzS/GV9bpktjuR8e534PxiLhDZ0pPl/O5zmGeyBvdLvyKZ5ao8RKK9NEQ+
ClBcGHex2wC2vfyteOs2aljTyPmxo6zpVnMrV7WthQfj4nlS7w5bPhxFNTuk2R8R
nzWcUdFjvkpUS2dgVfAld8awHl4q4QxOU1sV/nPC0hOlfzUVEU2N1V9/AixF4z/H
EUCO5NBSvvk7ycsvIAt6gIq+Ag+9JuMGSU6QDo8L7NyRTCoxEfShs7sl63zsiKLF
t3qacixReQ0H9+W00AKWHxOy7tP6GTdLDks7q9/DTijasrcYqYT0Fg34ik1VAtS+
ThfWVodskGxzD2xqM0nSLcV6+urDciqIV29g+zzO27+zeB94eOa1x69fis35W92R
Avb1VzILnV7A5m9dIckkRxOI7XoEaY4xq9AktFJb2QdRWbrNBgMM3WKMlLwlzGA9
ClWAf+qTBkub3kokhhZMsuQ8LVqdE0599fJKztqYNDvMvnIByFtNdnS2P7bpOp0H
jr8WuvtDfhO/Cz3pCt5AM3/vIsjwgXYMJ1TMpqTj9B0q0TdAL6dRj/BjHY1iSymu
lfos67Z7CTAQ/gI7oZvM/pqt3KjVl2i7jTIQuE18KOSD0mrLqH/05w0KRgQbOb5J
b1NNi/sqfcBnrm8UzAFZOYhJ687b+riVOcIfSRpNK0iJAtSywlhmVDBis3I0O59M
/eFRTQACAjYOwiB4wg6wX51AD6lBOF18t+mlP3l/0C6qAjpdooRrMo3zv8cBS1I6
VQ/PH9bBLmWL9nzF+HCIhsINniJ0J8XqFyFnj1GC3hltRKWToQjh4eIyzoa1etbP
AKo0IS6inmqfo9Zgy6zXG8wCFlm18fqwhhh3oXkiJNlhvK/cHpisUZtOzgBVE0FL
ICJ9cJzt8gKUcYpIHFAz49yYOP0KZ52IDeV/7ky+r1iH1Yi/BZmtbZjZ4lSj4NN9
o4+Qy5x+uaIlJ70g0HHZsyDrvmaZ3q2ttexh9+Le60Y170TuYDzu8PwBcalr6Jg/
j9S5Q7i3xfEPDkFhX5YZWz7y2UVxzYKgBHmiBHY1gcc4RHXgNadOLFjL+8gqtUYJ
sGdTyA3B3GfVwrzSIDc1Uory0A9XcEUJ2aJQjQrqw87ibzFZ1hNDDJY4iwhDmBBk
OnQlAOGMyNVvPwxsJD2y4DM+jCHmzH5itgxZ34pOEo95bFvmIRkKtUQq92SWBS5J
TSr1W5MGBNLvGKs0sykxKsHFCnKsOBy9hjsYZr1WX+5IPg8sOKgSTNSf2yBGwvcR
O/kH/oG0Fmi/R8DMrKiuan8jRhdOe0O9+FktiPpvo4MXtuWSYNxY1Ul9oWp0n0/r
AQhDnyDkloMyjavZYyXpOdaTExFVVVs0gja1KUz0Wfy8H0UYqlrAaQq8Q/XmUkJr
157wtaZjTXsxK1P4kWhbjDw0vuNq6vYI86i42rBghwIJLmkyYQnfGEVSooCo8XLK
ScSwq+sIPQI3DmqcGVnMWJZPG1UcUerMbx6CL2bzle7Y1FfwLSw9BPB9zTOu5C5j
OmGb5bDec/ftZt/I+es6ZBvmq1yimcUPdU8tnBehFQGjOyLtplz6K53G8IhJj/mX
gAf3CfA9ZBDkzV/qbJWIbjBVKLLFns/c1/eQ4lkuXEjZSyqTZgNX3e8DmWhrnOtg
FM3o6YA2KBLO4e1L0uE2j3dhIQB1j/3vb+i3r2HhCbYzjHKzaKVlOEe9muhB7GdG
yQWtaNzyM18ta88Lbt9KHVRlqPMliyrcZfJxwvm7Senhb4FCNhm/t+LyiUKic+8O
GXeLLpPb/DsmAJPTGVkrTS0dBqL4CFgnlw6j1aqpcdoy5Tm8btfkUQcAlKUdakfK
LpqsvF7pR7oesAL/c8LxK7iZFR1PDDY8JxxY4v7kLbzFK9ptQJy3ViFq6i7gtTlZ
vx2255mHPrOBxD7qXj8U5cGD5cytaawQEo0LXajSAP2X7KaIAxdWVyYPSrKwVrJh
oFZiOrLEF9l1L3yYM6OIBRSRUN4h0lbsZcs5H+tg36BJdYgDzca/rNwx3AB7+61D
dyyVi3t5i9XdOkxUaSGFS0/fYApRg5PvAN9SSJCe8kN6JgKilmeiauv3o8RqBCxg
x3nw0n14e0xJb/lOtzkwt6cZaiCbHJh/Edw14isJzASVhcXpoxng6GJQ77lHON7A
6pyirLV/HFwuwkyu6hB5W/8XkQDEqngFt00p6cy6MvRkSMPDoZwX2wlPuwXsbUk3
ApbrnbUg5/CflBsnQRw2WbEBQ0hCLGawd4lK7dNT8+HUc4UeWBbOQI+IZ3qov4ty
eIcwX8OGbMmUcktjjEV68xUzUbWNDxsz1iLaKLpF8oWISfnX1wfaxINRRzRp6l6n
9U0o689jIhwDM9VIgY8WcyzJ5rLzgLIsW18avGwUpDL4HCPmj6sSJW7u5BGlaAut
KDFQXvCH5feWFExbsdyydR+uvrX/LagFR9d+SPuzCyZP8RCtk+OfLTDKeYyVuxeU
A/6IMrNPjue/+pUILOfIYOKJKmmACIErO4HLNLNGVW8IfwUji6Hbz78bqFJAUtGV
FZYhhqKxnkYYe48evZs1iWbJML9c8NFe4e1iL27cWTF8Wdcmexlqctd93A2aZGbo
XXBMti10QmmrZ/oodloGa01Fqyqj1VTA5Mvr/s8y08+2DEjttZY3sqPrV8WKnMzE
FEepAjGtK9icPvbvBVgZ/Hvj4NONy2SuY0+/PeL7QzdJL1XcsZTogfHvmirSK5ST
InvYuG/X4Z/yy5Nr06CjolZ/1UdtgGEBO8o+aQWwpgXldqnsgiSYs+tvsj1oRMx/
4OjnMyf6GRrTRQQX0dZ7L7EzDWKORoTliU75LcqDPTMthmi32hkXHWbz1RocbJ5J
LaS4GOSDwt2SEIvSkP727q4BXFRTpZyo0mHPmy5SHkADzoBUObYHP4UIFaSqDCS5
hQ2IRoBIkqYl5cSm3rRj4dEZHJcqggV6mgJ1jHgtsVdArWqOK+NjzG+qm4y6UA5f
MhPXFINzR4bf/pVn4UEfky8znhBkyhGw6H8/nnvM4Ddjsum/yBr4jPCIYK3Lql1r
3Md050s38BvsTkT1SLtmSHpf0uLZs0nJl2TuPOhqDhw8wZHGRi4FEhhW0RWi0z9W
Foju2PYMX4H/0DsgsSX0YkEcq6TyHT95+0GIgJQsta6kO/Xoq7r4FMqj0TP2onB5
my8TLtUjdvkEHEw4w4RnyPg6KB9EleuMKGej/f3z+/V6Nn7Ih/7qEsqGVJpd/Vah
e8QZpirU53FEq35Cc+q29qLFgYKXS3e0RGae9iL6UAL7iF5a89O7Atc+DZ65/R0k
FrAVc+Zl9e9IpXLgN2Ue8cXuBhjCdBVbFfeR/bIyUmISBlMqs1KWsPR7iSTE4Kme
A48wQh0L0CxdxtpToi98ZTB+Aja+Nc+GWet4OK4U1kDRKMRl8GN6SSZKHcCtjHD5
3MFXmqpTKuUHE06Ot6ACmuQ1/yYPx8tUWfgqE7mzCwSkn7xfBamtoaRa9JVHzTm2
msm9nch5QL7bYaK23zYcWb9fgBFLtXAIO8KcO0cAY9vj6VBJ8BiziTebwdyUIfXJ
nBStyEAF8SfKRTZNaiREmX/+fo+xJAErRb+8YoYZIMb+8wK+I3nY3pg/Z58GPoNo
BwgZtdfAnn2rx3cmsXIkppWZvHGP4a9hn5SIEth9cqpHKjYTEpPUELeD+pDeAc77
vjsLDkDCVK2E/8XfnHFMytuAILeIs2aXgFphIiqBf+M6y2ge0h3KrZ4jk5PIIznz
8IewqYBBuauWSMiWzrO3vplpgWr6S9PoK1V2Ko3ZU//q26Yev0IXZzMwv7TBnJud
nsBouBBaKg+Fe/5Vhyd84eOrMpS5SxdteqDzRV6Oafgfrln2bFdjIGry79tp/4Fj
XwBgG1FCBnWidoonnRVY4fctA+/XzBsvM5kQ200sHlTJrXSDEn5PvEfaBIl8DteY
mPUn1ncbTEw+3b/FXYR9TzDK+/TWo6+2lJ5OEk+GeWENWx24yP+QxNWghzrEjAbn
MePEB7Qv5RQDrbVhkJvs1zaKLv+7d7UtwNApfnDzdzt9k2a7UNlKo97nHK5QiLJY
flpccbEOhnvONyJIgC3wSK0EBs7FRMSxbl+6cTu4jfGBZE3IxFe7zXtI3Mjga287
Iy3c7XYpw8qBFOC0iO9Y5P1V0CbOfp8EeBlrrsLlFNADfcmn0GPl2nxnDy7EQ8Q8
70mANwslI1lo1Y9AFw+Wpixf865opy807/YlOp7ECDKomQt/tSxJ4q6ZfH5R6EDy
hmmVZoF62g3V1fsjndw+1q6/GxdTRs0JmqWhYPmQdHP8ig2GjlgJ5TdqzkgTq7J+
2zUQpEGOfluUwnHNO+xYWBguBJlbcWus09m5Nq2E9hWtEbMUUfVAY84FiTLAY/iu
8PXPS0lA9Z3Es86O3DPU48RLI/vreapWwmkueU0KgloCmHqXB2t58MjAg63Dhnwe
Rx/5WA6LcTyYvjo0YcLvVoUz89rZ+dOpW2lycvrL8rKJa8onk/iz/JaxVuva4qdw
2NzQH9cGAF65FpgeUgT8fBRscP46tfv0yAVrcQ/++BIzbS0tQlKdNLAV4pv4KfEN
08ld64KqSp1d3TZrNcHYiIuOJEs3fAAoDu+nNFEFVFUdjdmWHYcBufs6jMcApCFq
IWT3Z5gY4MfjYrjDowEn5an0yn+nxlXGNLuSx8ZAHeOiwPU8rJWSZIyawZgF5p4+
7aTrObB7nI0rTwoiaU4Gx//2fO3NGUWBMdbaJajnyDPHOQOA/9jZsHtuYs0PnWYE
DJCEcJsx5fHms2zLf411VZgV7C2xx5A3+7ewuKh2Huss/vAmSzGndk1EVXMdVS2D
Fug2jB8nFpM+Crb3bTgDDazGV/uRixs8d8q+9ck6vdXmTtrpGhyQ6Fts7MCRRFAD
8S9PMyrkCjRAFAuUhFKZz8zj+gSXaNeazO1Csc0N0SJJHAV1ILXvZ18tZ/M+5Q96
zYuiQWHHlOqfrhHxdpXydIEDlCuw4nDgG8MIUcKOzzpbIbrgh7Of47cQq5Z008s1
H6+H6N62kD5xaeRnAjjfTnI9EhsrPZed8fQrPAR2eg9L9ebnMFeJcPl/J39YsogP
WYKrXXsUAVaka790KB3SNonBOW1M4VVs7s+/M+hy0N/715bh6Q59xxh1wRK296Cu
S9EtKOSebYcbmmfsoinY9p6J0wc0TPV3SoQlyknuanmReNjDA9Hxlp/AVFhjfiYD
2pzzv3J9M7QCVdpcesUJhKIh/gb40C7tYDOwSRMjC0/9q7hwEBQwxv+akPzpouIM
Lp3OwbghI8tqQc483SFroBGeUJWEP44qiLBCDE3rqWLvMtvY7oFKB2RHSRw49VpK
u3HkNu+OKhN6e/QctWoFl7nWzrYc0wsPdjf4XXzZw3ssivfv/aVe8waN0ua6bSkU
jxz+A/+SkfWgCvuD6H7FbDmil9srIVoNV+wFSLbph/u8Q6Uy85HXfLR/Tk16Ja75
2oPrpPI3zLsvLO7sfcy8bSfZIVYJ6+L9RRQl0Oe4vYD/st3RgoGNVhLrEoEpvJ0r
fOyNcxsCZupQEJrsVFyypXLOZJ/YmHTkNyMzpnDgOJnBkDX1F3FtH0wdfqpMkLVZ
vmYdgsDgHXYfJw8IQhnlW8sZJkDnscPvjAEFx/XKYzjlUV05QNwCCl1CN2jSil/Q
iL5+pt3SL23ZWsJrNZ3Se88P4MKkSXL8uQfMtaItfSEusvvtur0uZ+DC1unWAuFN
c/Zeu8znP3DC7jxwVXa3+gAXpf+DtEpUjT0VAnJFUcbwIQYUvbG7qbQv7kZ9N3Bl
usE7q9wsJlDFmI1p2f9lF4RRUSfU8zmlGkmmGcPau1JnKvuwOxnrmX/aP2dHivSi
G6G45gtIYOFtK38k8n0Avilb6gMmrKPVcXo/zqqr+ni/R0YYv9iI3BZumePlfpta
cpapqJRKx3z+rbbo75muAiZnbzR77hnddeaTXbVRq1MN/zevO+YCX1wlrJciNkUe
bT5l3a0FbpjNaXzi8OwTmDoPOJq2ueDCd9PVb8uKvRRuYE5beAZcoAYenPkE6K0t
nR9OoMjjuGxyCJydvGXtFblHZE4nQetlBapPHTazo6kQgi5NAtTDCrEM0yx1SjEy
v/uSmq5pY1KSB++1Wrk8GQdZDEfJ9DB44YMHPH221rKfHf1+BuXZM+vgf0dkUsd0
Jevc5jjpUirk2KG3+2wuhWYqCsZyZ6bxovjMYc/E3kgDvvuJiscVuyMQqBOfsDK8
wTmX7jZJ8PE4AhxjXA0OP6a0emRGSdQhEE9bMy712eYGVnkEyeAx1stshly0yKFd
DMdkdTdY1AbZRrW1u+6sukjid+TBofjKGzjjAe+2jwly8YhQrwAWVCuX8W3EXHnO
bk+QRAbrQ7D2PI90joydSb3de9ecPVzwqgjnbuiNPxOgOL6ungplD8Ou9ueT4+Gv
eOr9haAG9okk+iM+Ig7Xb6UHSyrmEsCbrys2v/abu0Gmq+pDvdP9iYYOR7wYQAKA
NWvfU43yKCN86zxMyDWFRxBj3nKqZ5CI2q2Js5e3+2p1OH+dEaIHe/y6zapMROsE
TMDyC8E7YQGkhWqJBahzYypJ+yyMwEMSNdaxu+ToASrBrwxGjPBI1o67tR1t/qaf
XiSqza7kyekE3fxtbWuNrrTzWgHZ6GMgX80+OK8FCMuWtf5ytx9ZpUa6GD6/Nost
FkbGu0KX8tJdbfXlOlUsMqPFnq0AUa6s1FS9nfEhpk9DDhtC4gtAxW9BF/zHfw3i
+aX6X/h2mDQ8AElHQJypoSebzisci+P8B4QRJHUlRgh6AR27RbHMocDY9zH3KTYM
7YdZ6y4/rSCnGdbZDFNdrjnGNtE2pj5EBhmu2OUwqbv5eBnb3HLwqQF+wlXEWBFP
yN9P3kfOrj8gsahZ0tOcyAjJl4aUqUQN1h+8cLHoA6vpExRtAY4o2vv14sFfy2/h
GmbVZXx7hMrjDknvN64ihwlxdt5amZwgV7azNXeLN0VrvdHZtgYdXM/4jF5FL//5
a4kSyIiubiU+A0y+CMZkyQ5B5XuLBRgx+ttYXBkGmrqOLEb6aVPU4RITcNXbWete
X59AFQn2NTHtDL0bgvMr50gwZSf/TvGfqMFZeG5Ha2j+al3NrpSVPjS4Xs/Jkt6F
Z188WcPxuqVllvA8RsMUgYN6VE3XQV1hOUL8HzT00fZ1GawSN84Kl8KKJ/xAtaL7
XC0hEvq1f5z/tYlzg1wRcboZHmR/QcoOgvxswkJCb2PFweWkMV/o4EV2ubVpvAeP
oU8OGdDoEkLj6NDzRTosg7Q6dmcW8kwsrOO0FFoxGj/pCeW5AItBhbhEAf1Inkbp
5ruYE+gfT3JPadXxavKqZEEicsnogEzGAKu2PkPCyakv+43Rf6SpAE3lfSXrs4Ix
OcyryhEWUDGgLgJjmomsdgTH3w9nXOX2Ef9vnKTQ2UtTk6ZVU9MT4LvijM0NbVQ7
3uCLg3t/5ptUaiWWv70SXAEryWSRm9BfKxinbOGhOufWRsTKiVEvhppU7LV0OVoe
PLLAJ+95s8uT/duL4VYP4Y5eV0Rs82qDwTIusD8zTzA6kNlEmUnbPsPqUvZ5liGy
bi1Uw8EQn8HAJt5My2S0DRZMJxtiD4W0+kN3Mx1Ut0Kj5qfSj4VhsTDbO32cr9on
7R4mYmSJuB39VZ3Ga6j3pcZQzAO3JLwWkaGY1S9biZCbpWbaVcq9yrBS9ZluSx5I
HN7pRv6Vh5Nbbx53cLhv4cThgEHPqnW30UlgjiERETcGDsL9m/+Kxl6ntGNQynn/
K06dB0PYyLRoYTCPdrrQvNmBvinI75My0zpYJZpQz/8KlPqTU9ZdokwZPGENXl+b
QqBmVRKgM8lx+norq9sk7p2UZ9FJGIXDtYbBh4KlNKAcpar2SkmdXYr8Px/5aC0w
GaZn69xtxbVsV/fDOBClD/20fqgUyASmEn4izZuSUYxQA2DNblW+fakyjvyO5RMa
yCrU9PIJLIpW03hhXvm/RVm09a4s8xdcwflZcz77/mAiu4RIW91rfi1LTwMFM6kG
yCfzjrYDFiK7lgRuenrlYPOYPnmEMOxHFg72C5M9In78HxQQvdj05n7e3hVYx4u1
8VEFhoBgjlvYAGeB717qpFMCTDJSZFatH577zjeyG+ecqdcZ3o/2uJUFLfkCDs8Y
GGOlucmDZUQvdcOnJZcg7Z6iLSKE/RSS6McrMRhjrwFbeQNRQ8c5mfJHY98t06+O
WcIm1Q/B56KNgT8NQWdUx3931UOvRxfy1EQVmKoEyK+1kB3+adPyT7cl8MFfD7Yp
4oBqEhFUSu08P2r8Rm8LAKxzMXlg7gZCu5RO45DqqqnFuaxGb2kipeaAI2hB5wwl
TZG05Kab5UmajJWpf05pqK089HT1ocT1O5k969OMA5X8smTbonwzoKTqiSIybjJP
ip6/X1+kyT2yWm9jzu3A/xGyWXiA1J0eM6718Y5oHRRF05cKZOYOwvdh+8KwBtl1
d2KD5ZLe8rcF1RfMkemrIYw7KOtDAErBrv0Rwp+RRJzoHOzl1P+k3BHzi6bfo5zY
qLfMLF2iXyeA1gjvwMS4gXtMxzjcJrNSAS37aMDEmQf5iCes80a+c5+3CBGFz6Qz
h0VlLvFPbaTi9ndb412+PoTiFnXEjjOobpF9UEVXPRcVvPNKUYziegRBBYEiV6UB
R4Axxx4+903U9Fs0aR8S7fFcWoAP6k4rt1Y4c7IzbAtY8kQvx4xbje5tgah7GRLC
ih4iGtNecwSBRShSHrCLD0nQ8U8lQN3RWSmSqa+sbWvMq9M+pifIhOenzS7iuhLJ
Q6SKeybvmrxDDhf9PSqDjMYYsBgCnc/q/1iTbKjVBqDiUB+zp8qFz7N2TNlhTZSj
cG5bhVHTABUEF5mdw2Z1CK3NyZ1oONt6UML1c6ICqML4+4svFtJHLJNZbD65BzP3
nGACGXj/x0fiojd3TA8+m0Hy9kBx7DskL5b5+iRtvdT1IVpyto8OpIOjSckhPeG9
bD0IudQrv+L70626xs02e7cpPQcdNGTJ5Z4AzpmqJbG7jplEjq6j/Uivaz+GoyRC
0lyxgjF9kF2Hgql4BKUGmwAN1HUfcpbesjEoKOYaDGILkYdaqTE5zM+kzc/lwVKV
3G3+zQ+6esgmomZIA4ycxJ9eOacLJMDtPhpF8bGDh/MDjdUC77ESqWoBO9/P/uJw
Jnjjto3xXQKegU2oHpIOjRUf/u+U+lxFctzYBy/NcGRGKq7wwjVB6I252FawXSbF
/p3lLSgGwo+ClpKHr2i0pe9OTszQ+Ec3/fXwzASo4ATyOsgmcF7FqUSTytCI/sp2
9CHyPsEiLnjdeZgAKi6mEkCHnQiBSRjtZQTp4d+OXtvAPDEZxR5sIH7Pw9tdcuaL
vZsKXOwKEcsK7Sc5Ir5noU5h7YfckxoP8pAlxwwu0XuvJyusHtmfyGmye8fjOIKw
JaHkcv4AMSatHLoxoubivuabRZ+z1qLChyG/tw2enXRqzTOAVreo4ULlFVZoo80F
xzOJakPzWTkpsQ3W5UbBnJfyHLIL/J/83QrDJ60BVRhlHP6qSLUHQqn7oTiyST9F
ACoWq8c3MjT2KxZ8fb1U+Av936FnrZb2jbYmGxATjCAw/faOUh9/wjg/qIFeJOfF
KaMSwx9IpD5BJ2/O7rQPCZSxvelLNE5/V2ZSlZgtA4mQDHvFbCVmp8FmsmEMkT1T
kkE9TLUnJla1uLnuVbb1K7t7344DwO96rmVQ4JqBouR189uWBO7Fv20eX5tHMNUG
15e52beElDcPK8ZcKkAa+LvWeKoWTOO26V6+/UHSENqwInwuK0IFZGJTmfEXJEMj
IhmW1A6I4n2L0HpnWGdrq2Qxatl1JVsLZjcouKfniy8yC9v4DtzZrKWzBRkM4WOC
mXD9XEMVEkTqYd2zpuboIh0z6PYLQBZdlrJp7ssZbLcZ3jWD263ecrwJ/a7j2RC4
DnCg2sRzXDXuXvExMf10gYqCq+n7AqtB+TJwnx62WsTazlwXNo2408Zf/hkkMFpn
DsT1139wXDdH99fe/lpICy0lmuIlKtydU8S7nOoENd8bp6hhFFrSQYqyh96R1P8W
6mog41TUSzlDliIGPLABKsz622mUkY7rB2x0J4FMXFh3+3meUosj30Bu+d4jatIa
UGXlnMJIbnosA8SSs6Htkhp+HqkFe55uq2OYYqnMkVSiuoAEmyuKH0Qf3A8CzAjj
cRHBcB3KhBuryWFTwVlQwmrxVvxI4eWP4uSx3MZT65rquY4pEI+jKzhTfuPBER2a
N3O5oO+vLTdyoZdso0CkhwmQXRuMRVHx7l28VWFyA7iVnf6IcM0KXfqRrws7dyD7
E6HNXR3YLk1ltTCHpiv2do0SnunWcGsgqXZOQ0fZHt37L/+UP0C5voUzFTcHlmT+
jmhk8lZIJ+ygTZEf0dgDdtbneRgXb0LJZANeYlnm6Td9x4P01ykxqKPzoACjSz1E
C6QpnnPoDhzFsQezpAZRZkEa1//RMoEn/cBYMgcokM+Nab81Sq15IVZaxadTI2qx
SSli41W1oEkV45VtOrqKtUNOL4D95qoaA36KLN6lM3VMjG+OuItpSpwAemYOUOVh
7VNrbi4WYup6N4NIPbA2U9fvsacvxufriBj+thUfWnFwcLsjno5TJoYoM3Zefe1S
TZ7fSmYmx2XGj4/+pDG7xS5ahT6i/MoWxgMzC3go0gOYF1E25zopGNNm+0c23bpu
ECXXaivhTDb1PitMvhXheBiJ1COSVy5vRMnlfdRFs7Ys7pUgfBtauL7loEvxC8NJ
edED/nmehr18/Ur7yEBlRRBm//h9fpek9JntehLr5L4hyoKFyBwX7HD6FXMZKm3/
uAUlNp4B6xwrYAnAfPTbxHlmGnho+f1p2f4nexAQNZERMCAzMVmOuf69Oe/2BipM
lRA2CrZ2NttDpNpV+tKABaqUU/+BQz3DgOI+YBKJ6yUGkyHDtP/MYGjTRA30Ksaa
LBuba9TQqdVXMTiyEePfmYrctBBIHJqC0Hje2g47EK+441j+dZF5rVW/ybpKmJEI
I8VqH8Vd8tVTXF9/hYUpErLhgOhehu21pGdfSkBs0XWv+3/J7jdqvsH4N4Qb6KX0
1R+ZZ1IpYfEa9JWA/cVe1SyOrWJOy3jOEZTHG8wF1B8omjjgdulQldndyb5svQEM
/wy5bBTZ/EDuDg26Lu42LglAfvCqFEi0VLGdv32nmLL722CogUaBmDspkKJzwT/V
AcmeKaA79U5GTS64HP3KcGB+AyCiGBJDzE9B6LLlAmnd5L2OalMyMfVcARqT1V37
/MqKYaNoE6C87nImvHeI804oxawXM1h8plc/JtHWb0ybo42m7/f3jO75HUNQOG4I
uUfeUzE1nbai8W1eJNfeOMGJai3jFYME44JderlAmCbUKMG4wWV/NEunv8cocWpt
ipRa48/eIG1pKlM3DPgtMc834KHWxBoK19m3B6I5BPLAN9ZzNllcqDxrVxHHq5UU
Tj8g91IJU9L7e8r0MtNA4ONrpsG+Q8y4gUHupbDMWIBlR1TJRLT1yicMN4LPRAJ7
p/1XzFEzEFjX/iFafl/AL5HGl62SCUuruZW/8uXui68K0lBsDuDEu8ZqlYE/xSG5
1JqXGsSjBV6HQA/deL/8KWzQOeJQ2AKdXmQjJLlas7mMtkwm8gDC6IR4aUAY3xmv
sKsct8LNYINZgiSzPOoL1sLbAOLvphnO6eDCunloxoUUkBiDOOd+NmENJgJJ9pzs
kCxJlh1oUxthfnWkw7i1a/MTga5cJNDnCVHRC1o+5uw26cbY8l9q7FaxeTT5daOz
Sln8pYfh1PdmLl/2U4JIQl5bYIBCIQMbJtrTrlCkxu1EbZIUIDeSrX3JjY+bGblN
HfHrr8ycC2tmrKlJssltnUK3n4fQDUUv2axoABiJ98hagLKB92TjcRof9t0kIh7F
rShppdYQJN/oIeyidLpnc2Npbkqm8TDCe6jGC5rJkt3jYVx0YGMSfQVj2AUc8xt4
zIGaVW2QUOPryhO2Pd3xMJdM44ZN/btWvyRTMfWBJeZXVEOo83ZTb/btpcoFE2Gu
TujHhoB9jJ1Bu6nH/dtb3ssYoVjMpQOquMTcySgmYs0dMRAwmX9znQ7LOh/lv7MX
5Kgh//ITikqOouzywbRgfllFabCzXoc2h5nH0OVm4nroQ86qoUE3jKToefwXYUJS
QeXEmtvlILU3iAvPNWUb/om+a4NZuxUww4W/JDxyru/tISN0xsgBz3PkbVj1/kAZ
KYcn3gmFCWZ39aK+Qbv5ImP+dQMi0cRmOGwR3uMIqHCbAiubEmLuPnK843plsZGn
TXhOMNtHBA7kNmJEBEd2AuN/FnSzMauVTwfCdY9M8//U0jtWMoNpV1mzb9n5l2B/
5zJpbZvJN3ga5vW1IBC6gvQiXHQxPoSjvkUWNqFYPoBmFdhMy4todzv+/6fUGS/L
O+1PdZOsIL/5HAjVoisimxk2Iyzo12xf2B8JhE92UJ0zGtfgGD0v+JBOxsyowJA5
O7wlOAWLc3ctwlGACrtlcxD17lpdMp5RlWzjTk8C2KNEsd698gnRntToav9Q/wEP
X6/vIouFmlcm3Qxa8A35BRHVnG3E7Dr8O6P2yS12kRnxJzoCwLo0e2eXbKrhkdmS
Y0OFaHPxdZS3kHj+iS/AAt2z+tJr8i7ITEIRZudLhHmZZHH/vtiAKJYwKl9QkZya
xvGebluq1qJmIRIJFEbJNiC+PUr28SAsoalIT4HqZYPtPAc7E1GOSUcaP0yKcQdQ
CW+C8xA3SDpkpfNKwvCFlHG1vNiyQUaaxve9bwKQlWFj3xvbxgde99tJqQQbl6gy
bfSnb/YRTI4iMX4B5OBpSFG0MaNifMFrhpyNpWhi0OV6bBKQCLzgIwqMLpjvcn2u
1lF6slhHM37k3Xe4RgzMm9VSjlJmMGgd2ip1Fgwez/+uP5iSJHWMydjMOv2G0TDq
jCgSYqSoK3M1EYrPU7UbYGBGgXzgwiDGzY9oEc+8f9chq39NzRnK14fzczY65516
ljhWjj25uVe6zToKdTgK3zMEu0AmGHOQyTNvdSQ9wCwqbo56heOLwQivd3C+Lo2b
LaRaTsHKY3CR9hX/btWGRYfzXbFDFf6lfxKlHWBEJXUxhTBkRyylPYG+f/mtYAkA
MiAPFVyjalX+4Cq3NkvjvJlb6EhT8PcO7wqxVWGrUxBzryWz3HVyLHG552vZcUCk
eSZUAdSFxneWY5+zQ4feETku3DsRtq7iag7ZJ/eWUnfV0u7j8ySjv2i2DDg+OGh4
qGyevgq1/RNGchFuLgmYJTKZTE2RCwHhqaxTpVM9oQf8Pf6os2g90Doha6i6xlTB
MhyzbYbRf6LGvpTK4x1udkx4pHDxiji3oH8vTUHIvX8P0xyo4juspY+J9YvHBO3E
CL4fAUsFFGa5xkK4sZl05IL7yIRQEGbKtBlQmDS191Jp5m7gfGkLqZ43CJqo3ODP
0P8ANgI5kpqhJEcMcYAgm6gJC41TQPcrFWi2pbW1du0dq+tS7BP2Gp/Jm+7UTKDq
QjfXvGHOLpMfkPQhKvW01nMPDsNetrXJ03En82VRPEYkFuc7qwlQwfu9GJ3qzHIA
YNPHxw5qQQ3YCsq4ubMP9UPrC8a6fg5FZx6iyBy9NvknlBjTVD77Zh1fCGEaJ4bC
enMW5lJicu9vjFcj1z+HxSKqJ6+HmKRlbmd9RYKaZDCx0cuqmqks4A+cheSWrGDG
5kbRVvRwgSyiuR7jorUuYov9MSAeeuKDK+Jxta0APNUHZG+iBW2KxC/uO3M7s5u2
+wNBvGzUWh30yqgo7r0OdEMg17YWrMOQZ4lB7ImSR+TXTcXt9qo644h0ykAj70t3
+/jtHXdDymAmc1GtrngO5V8sieietPEaLCgL34UVaH9xbj3g+d643FlyxumVJvPd
mKxLz9/k0XOW0huTgSEvcaDLPr4QBR5Wk9LnQNDksI4M0qFR36ZmdEhtAwQKS/FG
PlecBcY6MPpTVuEOLlJhkDe55hjHhCszL89LYlpFibNpNLhuouj1R/mWfWeFoH9/
+B6p0T7YXCL4nLBUU/h8Jl5H8FqaIruseExfPyfezGtVAneRzd2I/HXidjZ1T9I/
curEt8uCgPJl7ulgqwXK57a1yxRuhZfvfeudrPAV9QvFLRpdLh/WON7s8ulIoq6E
Lwr/Zlo34lXH3lJStH5TPfbr/0dHiUory90tHNVl6RqNTiwATGdZ8QW6t32rr0GJ
Y0mmwUT7/NC6eEFEVk6VTPp4newEowXdoDgwa8/4PaPVYV3eL8O+jhbzHunP3uSL
lsCAmESfzP9EsY/r8iuqIAGOM3o7ty6NMU8M9C5efy0qdCOf9zUq/ItNeMVSTb2q
aMwCBuxx+mbmR4qfx8u4qnYAWrxtC0M6PHwbmMtHWRoRJ6S8PtfhuFe9vH6jruLw
W+iEP04sEpVV5fYrE4ppIcbBzTOTqENJvR8UsTCuUOMe1xSg5+EPHrNeFNQxJkg7
7a/j9+32EudA8wbzNvfVplkK1fjyMOou4vxjG1xyYDkxcehMqCaFp5rL8vQOCoaX
KOh35JGCzRyZLhuk7NAKJRTyhWxOrOJfECX0D8g0BjdCxsctuB6lpUehwmTz9vld
pPgDUpNw+v7pAM3VMApsz/T9bNdcREd4jTwwGj3+gZymCavZffUKxch2Jd4QB0Up
P21vGX+BtWZYLkTtquvVcmyBveHsPxipsMQtGsNvkFDbhsi8xRKSYKqcEwmzMF1g
br9XQfzmY4jWu7ZRgBM513EdhMS85Qg1SDtmc91kQ3Qy7V9ZydM/lL+0vBhGs6Cy
Llia8p/VzAaWIgggkRvMjmgU1K62wBDgk4yFy2aOkjMr0asd0Xg/orhfPSZ9IhrI
2EzbDV/FuhlhSS1jxm1caQvTYecmtzB300dKst57GI2uWwiWkeOsVCyJ/zziGweH
574lC9t7uEeqAyfRSK5UeX8Yl4jGJYrVqnfrLBIVEb12Z6wBotKteZBDRSVf5szm
dHBZLatwrAshzmiz/vd91b+NDRpCQKpRs2DZ8Qe0ElwBmTwFvObldYvLj5amW3RB
SDlg06ob5WdSuJk0lT0P7OvoCGqSeBEqVTXiil5rWrjQe8YZf+MlEPmNxrX9z45y
OvD5+WHwfcZEAyRj9kyvjbxoI8cuv7gzCq+NgnKYgHEkG6aUmqm+tydXg/uxblH+
AYr1URHzjs7ou6+4V1pTfg7Rs/y3AeAdfZNoOeGcBiKUKXTzZTEdoenFo9ebvPVY
pK7ZWVFrFWxLms4u1NlBG4fyFCNI6NuaWBAYGjpuEtWpn2dgctMewcg7MKTwHuOH
XWDOif0E2/VNtnHVAwWcCzqTj0xPe2gzZ2Ce9Q/OD3QZCPFbaiRWuJa9fNaPywfw
72Sc7Mlxnxd5PDb+9/YXYlPjae3/a5O9SkgIjQ315eadGSvxWawxECr6GcEsKDfO
kQrsj5x/t05gDFVT0x8vOKvKtqvzaSosM87F8S+gcO1YNR0K4O/D6u6PJq01+vFh
MndNUHXT9XLXvdup8xn553Ut271X7D4T4i0KAgxsdnKnhkW565qUKsmo9StMeX47
UB5RpNiOWwsL/SZqq5v19t1I99UWpH/j5d3t/cnUTQahIQNEVBMvW+91KznmmOCh
PrXloLZb6tMI2XRrNSFBEtns3vOantt+7a8KiLWyMLPO+2f69qccV4iPbdxsa4U1
WcxB2b+whl9kpkQNM2gGzWA7LDhfcgkV7/ehK6mAaN69V6BF8j8Jk2W5skbrhcze
kh9EyI9Np1d2mOcG/C1Yp139e/GjnePpKCiIPt7Fe/nLe+v14EeT6FtiUAJzSy8a
nf0ACrgt4+c/F76MGGr+h9pxFqJt9Ue+mm+fcJlH8dplkM9hpkAYMlCHrumqeIYP
PUC/Qw0ZJWThlgjhf1+HQ5wNtgca1gxJRxP+0RFSeQJLe8uBzkSjGQwLVgjrvLEq
S/iCqU5KR1luZEho0895w9G1poXWEduxhHBsB1iTSQ718QKIIGlK9uB4rCYWAapO
qsxyZ5YUcSVfB1C3BisLGHeQS37Yr+jzjQe5etbpypjUxvp2pnoM2OWJJqCazSG0
m0XkX9DtQvyCTmcyFIu/tu5b2Ovqhtf5TykKNDx8yeWXrpWRNMHRFyVWqZGOpUyp
OKZ+kjumlqxVkiTWgkeW04x0mD9WzIszAbNQ39Uzrm8ryWjVQ3kSBzWwEQK3Kow/
SStV8rLIis457AQR4J53egU3KtIX3Vn3hYyhRrhUDa/xdqe2XqNowApDpb6+pp10
Jr2ALlBmTS3MI+kTydU5tB6mtnO6f9Qo4ZiRFMTpVLGs6ZnEFrcCDhZ4yHJA/iV0
GhAfoUHtPmveYol6bjg/PNZn0B21laAbGbPhIlcEX2FCLmsZCFZs5vCCp3tAwaPs
cVCPMH8hQwYC6t5BhV/7bidiv5eieUd5E37zguiRxb5bXHubQ+lAjQWWZDNO5Wh7
UfYhFckwVFAfJo6e33V9ygDvFPswV89XZESYdaEBSZmAhAAnvLwzZIqOEeLMWls6
Tyq02tTEYktS3uuc5XLh79C+PhmQN1Sesmn3hQHYlJ8lj2Uk5z7LPDip7lyzX144
JoRWC3brVzkdHnrhx+E29ExDGsCxSgjVxjd+qHFJfxW7uGAQ5SiLTgVdDw7GjSUW
JP7ATKzo0YxNTjtIRoVLZrbtmgV1ATQUnb9oAw0L7Cd/lMTnOLXSCTOP267Jep5t
ZuN2u97uY1w0lNOtpx0Ut1H1+wmh/ePh72sOGJZ99NWwF9V6iK2kUHXT1lrUn5Rs
SiHEAi32s+N8pIfrqjY2KpfMXsBXS77o8PFQv1kt0wk9k1bOa5gkbY1BXOQTglLS
qO/mbQHVL4WoHsD6oee4sycF43jXzCxMuAop8NEG0OI5TK5jbGAACYIaliIigAhG
2rdf7FYVXSXcodBv53ssnELSr/vqI7Sgimk6rf28CX++5m7OP9ojahv9qcMPKmy/
IQWRJ5nmfRtvayr+IA12sQrKhUYWwxYH6Q89lc+gFrKAYyP0rvkpUXHvW2lWm4Qu
cEwrhc+R6flIehiHEGN2E/zuUev/zIOSZUfOhVohIRm+bqn4BD6CcrncJg8d/9XC
tkwBKF0KhAnrnv0OrzuyPy9UjLECVcO+bzEt8a6XLW9MRGDYXzEsFb/ajX6q9OZ2
IKxHLx5hwx58VQwe9Iyh+1rHSvU2kq/1vMDhkf9geSDUubYcXXlXcJh/prBJ6fOj
/oumFTrDrUIe9rLzt8aUA+vuoKRgjzUVPqF/e1FdoFJALGb+WTQsDczG7XgmZFjg
VuZU3fesCmVO6Soij5nrEdPXvKKbfkhU3PwpUCSpnX6wLlRfNPA33x0kqOfNWoqz
lHfVCdDnCMadGt4fOEiqczzu4vzQddQV/Flq5S9iO+QoyN5deT2/bb4x03VuJEGC
rCESNIRB9i1yLVhwvIPk71iBz86u8ObWhFAkAawc4MXim7RGfElUX2FdN5Ar6OKX
ObwNRfg5vmC1QElI2jRc9nxSwXb54p0PHOOQnckK9mbn8NcVM2qD1KRE0SrKF9Sj
61rAFZwqatax47gY8N6koIM/IXEg8KP8KQBI8UbYixyOifJDH64X5CBzjBueJ9/g
nOUdDvhlLWCKQO2CWVDjB82dyevFL7zY2JkJStvgy1jY0gH4F9GVXsBPkyWFhhC/
bA7LhUjLQ8x8D/ceUb6iB6CzMc55Iivw8W1NATeDOu3/dlucU923mo/AN+qrJxSZ
oY/OEDvmQyGvtJaKNIYpEkfmZHuPyv9eYPNkxXfMtUYTs7fpDl4Git2Xn6uhHMNK
pflNXbnGzsoAcwOTX5bs8B6KnbWH9lSYf43Slmi2YqiZZHQWg/ygDKS1wnuytCbP
c2QdpyKBVxEyDmIDs08qtoLAVf5LShp1bUq51dN00HmiaMs2sjHRd6pE+InoNuKz
SXp+rsFjjwEtlEv8HkH207SavoEy1xvr3Yz0Fd3bm67FajjfTOZXQ8m8ic85JPHF
kM8SdQe8XW0CXcYaDWyPi7gFulGGecuQ9PIaobciHVpITL+N5qaChE920uIXyK+G
fAE48bS00QN5eF1pT+g3tL7CC7B+MgiqN9hA0FrC0E23DU+Z5Dyv+HUuaULFRkGs
34I5ZA8cG1CC0fjpJv+SuImUpmb7xNWMsXPMRcV7N+8Q4Nno5P489iXM3bZ/++ex
BhTm2vziZPiZzlKLEhnBLSOhOpF3q5RpUL7Tr56fMbQ8nKARywCu9sxt4ylGhHev
Z8UPoWvPu5QaD9W0zABtWXikvKoQNsnNgGRdekzXStl8DkvXwp8vQxzNr8FsxfuO
qx+bJ9MJlU913csHrqAnqHNyTjyTudp+u5DBwmMk6OYpKfzULci+dVuZZxLim4Bn
hIUOd/gKtZ1FIRPx8Su8LXnj7TNg0MztInEht46tZIihZP4IS9+Dr6STlv/uDt0p
Uu1+g0O1yYURruXLi1FvT++G91Y/JMJLfr48ES9kEhNWPSqAFYcI9osVdN82QfBt
7rZ5B08J5PhXa8+uJNGLpCE7odAseLNqkJsqovol6rCWS5+XWLRPl2V8xHiGsSQV
CfBexSpTbTMBIZtkNp/c4LQR6vFI+XWkLtp31wWojGV+d6i0kqA3PJ1QfmCaDSAy
dz1+aCI9b2sKNiGsa8BLbw0pcZBDnnGPW/N2g79OHizmvfacabQB6T1qy0grDq6R
H7DkzF+14hS4Pjqyr5C2gYv7eq4f/cVlXnDVebAGV0NkCKT+YUZ8HLYOm9NNPiw9
6sYU07h7dgbOTHshQgjN5+4Ws3c91ugMz2psqIPfNanIkn+EigQ5w54b4RcrwnLL
RcScB7As4gFtFTIKJ4QAHC7N7nYXQ0jUJKncLyhQDEVC3TEzooUz1YcYJ1GA7LGY
bo+RMPYLiuuGAUNQY2vJMQu8FQ1VitaIXNc0mTdGQzooVaHku4tnW898QA7oKniO
ICGMurH/PgKEJhdhYh/t8spQ9GUDNqT4WzKhf/JYB8B9UhPqRxtGK59WjLq/luMc
6xfNcX5J4PSB1fxcNMP0ZMGpYIbFMOPUvQ9KSAvuRuKHLYihAgPY0JDuv9uEOrrj
ZvXfR8IE96IbR29LnAwvh2EYuIneCQ7vCmNAcmm8dueKHGATcfsld4q0sSqPD9SI
yakf7f+JXu+f9cFcICg6R8Z0Qx6mKAiYnOLnrKYxCEQWb2TdAdFphrgVEOHK7lKc
/1ooVsKq4HlcgeOkVfu8zHDsxACGGVrGaMFh9kut4uLRNM2yfN+xp8YbIpsnNm0+
967094h6GgOJx+krP3akX4Gf0VsOPphScuHx0z1ozhRO9F2h3U2KNFacwyFLZCHw
Hr7szuGOQ4Kz+VbUlUHDgJL+QZlRif9HMfcMNczF9Oq+cETvkQStZEtttl+wCFx0
JvZDABDVqjPA5XMlEpnjgn1Bsp1MdrIjkRful5P5paInFDJUVLJmWigOF+caL0+q
T+8HNdM9qTpf7WINUgFAHQHv5OSUZ4fvjmmH2VaP0DIBMJJ9ximM9VL8cBI+RBbQ
VAQripXxhtK3qwAVXfEj/caCFaWBlYoiLWTvmQy8Ad/iMKBm7c3GeYB3i6pT7yLR
JylN8BM3t+t+xp0o1eqr7f1kCGGnztDwr6FhX0V6TP0m9w7h3/2l47E2863UfqVd
trMtRcCFVefBJRFZ7nfCVOXt85FYRhPlMvqntBC6Ccoi5fyKAKE7+XTL2nM7PRBa
82nrx5JuoN1hZmfwZPg2HCpv08AJkAiqagHAwZ5RezYq0pTD5hDG6Vuq1v6rXypb
yNgZj+mA7b2FWdrqoWcw4grSV15ei5V+KbVsdto6gzvfv01qeScVH2AZVz9X24R8
nwzAuou76LxOfHPDm5RUqNMdKVM0SyBq3Y45GsdMHVW0/s+jjf0dDIbMNhzKKINU
fQDmDcyq5y3DHoUf+PvJIeBzaOfCjwJZjj2e6ehl7yb89wdRM+Nh0cE5oSSaW6Pl
4Jk/83yb5u25TN0mETMkA2E/ad/kzZJJTfkP5yFUWgQrL5ex8IKyb0aP8ikFK2fr
lCUaFSDpZ9tHqRuPO08SKDTpzjTSBL2QzvCjyXtQFy+DlBMSmqMKSBVjPo/Jarcc
KPsDAqhFfwKwsR5aFnNmYRQfF4Mn4jUY5avFNbhDppacagqpHZtKIYDylXyUe+q0
cRx4+Tg10Pk4uu/KC/d1FXfwgeNIKVa3SXjDxMYk80IbK2QUIXfek/nmD4A5G6vr
x6n+CD/mRgJ9x0O/oq9R8RVfpGHlRPbZYbxRibONlwNQODvXY+/Dnmu/jXPbyWkQ
4eivNdHaYJbit8LUwud5jKJEOoFDCrqSeZ4so/qzrxGfp2Y70XT9dImkm/Ns0HiV
r5cSc6siC0j+9wBAcmKjj3hac1yFWaSVCTYPQTttuKq7Qr39NL+3c4Vrts4DMSBB
UcnZ4+ZvpMolHBdBGwgZLUd2Ylja1Sc0A6qVgYIjCvb1Z3mFNIc8W/RsC7le6uFT
1zczYtkx+jmn/XSUG8KFMahI2bkOKY0AMQc+0kWg7HwMZ9dN11jxXA4rXb1T3oQJ
xG27L0Wtg1DWd00uWV1cldvCJEiC7H/MPgAu6LCBvhZoQo4Ts33kBXKsV1SL3arD
VbAmwTpcUOO6LDJ9LRU067yMF00Jm2FrTkBA8iGyrWS6zJavckdb0K3dA9r2XtvJ
QP5DPHB2KZlUrnmAl1lgCkxjJpS8/HM2AUqAi0HSPfJFR2xP+N4YlH3hpRXe74Rl
SGAXD49Om/p7EHnjpK/0KAFUzKYLowwlr2KFAbbmdLhcZ7rmSFNP3IffghgwQtsY
ttwRvs7PB+Q5XhBAtX/bjc+KBRlSeo4eIltRsChHLIyHfyhsErKgXEqsYtclKMBk
tY1hh59Fcn4ypw19R47cbJbyZ36i4Jz3CGgjZoMSYeJ3zYlcefYHi8fXlzgTIgF0
v7I4dGcmSz/0fawgM2yd+jJpWZo/csLOmHRU1yo+cztXRgPtqUNsGWBLMlTVPVkW
YmmaouWDWtWxE+x1+Ejuz7OrKdWYKT6mCrtAFuLptkcuYX2m/ABi19aT/fygy+tJ
urlTDrdAeOhfvwP71YWM3ftes1BRA+Ldbf747LhJQQt8PamG8Kr3oYaRmGq9DhKO
MgN3/zrIjofx04dNKvEqqj53Z0nXNg9owtHVLadc5Jz9T7VkYhrRA7tnTFckRqKJ
J61XyrPyXpjWXd1fn19jgDW7OAkc9yohNgqIrZo6DtiLAURA1i97xMSDdzqYJdv+
nkL6rEGENkjH4jD2pcipx9zv0DusH1ap+kKnVpzU8i2agkfKXJtPBVkQHdCe+yeW
aCQHuvycC8UE3V9rLpXH9oFFtjyUABw+9MeYZwRGi+66oDDST5FNs6yt8k6fCeB1
5g8+GwgMEQZjTk/NHAIpzjSj5HJ8VMyArh9WeXj/yG7OdJT9huJZ9utudYxheWQg
uSYzpjsHxX6rQNRRdqp4xhGyxNgkULimRg5sc6LpiZU8JBBRhmCWRS4J5KHvexvm
64get+VQmefdyfEOj4pgaRhKwgN39l6zRj0lqTxe1cxa6deiNaOtuZkW54u7NJ8m
+lD19r7BhErTkHJZJ28zPc1O4E0NXinOqFwGcJDXv7vgyRpST2wVUOSqm1TxrLiB
ZJ5g0NFImEQv2rbmEpXjRrrDHjV1RdyPLRE4c/dURiQ1WBn20vaYEPz5ZoFEhZ3h
DbC3H4wIsSG/4qFTitTAKPwIdbhyM973OwgIIrHTL2yA5t/KMYk1bFcESylPEqcj
+TKdQI7r8oQcuGPd1vo/HZkThcFmvr16GkwcZNJaORx0uS2qJBWfSeTF2Ns0fM74
fLmwmE5HSKBp6JIoUpvPpjuh3l8CV3f0vHfgqfuH3MbzQWJn9nl73h0hY+Mdjyj2
Xkq0cR/y1fICGHqyUl6BpHKc6grdpw1wpTMly0bcsNnx2Zm2nz472grVjiWObANj
IlMoTl0HAK72kgymhOqG7g/abW78tipe6WXaWC7wZxBJxIrUM3LfaKdaejXZjDWn
L5UyhmkOEimAdrVzzUfHHqsmLO9uiURFZzF/YxowSY2za03fd0htnVXsuRHspkxA
qnCK9mtWVdvnMOAtwkXqmD0+vbMfzsHre4e825hI/4Umf1ei3YLvg/q7WlCtpO3I
/Z28fSLyYp4G9487tbWECXO/6h2gkxTraChr2RvZb6b+rVb7p/9CntiPR7KF/NKA
lg7JlawecYESAxun+bCPEzB6lqR04ejz6230qyH5Rx1prUpqi0yylrDcEilTRUz7
3PBbHdeIgmk7+833wrcVTwxOrohVKygL0RN5MzKx+mSSYvhODZrtpgTRuPwSdLrT
Xjf1ZPKnLA2g4kCf9JU040VAxJcX9/a6XECesxsCDacPm9u1YnCdJElYLYJYNr2P
IfFOTZ5f3CyUZYvhOlp+SlAbRDNfECo9Pz16Xu1dLD5hqKFFTJjd9/Pmp6pKwHF/
Odwgk6aU/GDocAX4chEbgt/hL3bUomj+9ASWT8w9/uw3tAwp3EaG75Z88YmlqZfl
3za573QcYT+jEt/GuW6ez0prVzZ9VIl1atzl7JKAI1chtO92BOYebAL7cMm5Ruk/
vMBVxCDA4wnX4JJ5djkRgtJF7AZCxRl8qcCMi+SNkR2gVp/MqIciUu9mxTGXMZab
3yR6roUNk+j90z6Q2c+WLRPrHFqKZSfesyqwULIYZzx3zofeGVOBlpZDr5lJECTf
xiqwqRHTOUBM/zj1mInaYWJPlQ6+o/blM2dd1zrDhgUOMuwM/N9oHRYbBhuNgt/W
OFjov+MoeAYNok+N8naM/884YnTKGgjHFfhi05ew6eKTKAOeT3jjYseM2pMX9lYe
UD3H+r2xIUFlwSC9QhfUf4LNZDJ+oxk2NVquC+5KOHi5E5ZzQ7t68Rg2iuKNqael
8mnU9aNTpDpTYTa33nSe5CrOoDBDpjMM3B3ByxMOcAFf7jsmxl+UqKpSc+5r7X/S
IZ1dWDnpzwc/z0c428snPAiMkiVeDF8gB6xKvf6nNKuS0OoAHqdUp4Xh7DBxmtId
00IOc+ZOihGnwq1OCDeIZkKJhizngoS7unT2+ddvUwmcSzuyZ+2JhVt6pJ0zdcmq
JEEyOCqs6vYOgMEknaMEpuI6R5M1yfHUuFpXFFsW/r30uS6/LIFio1MyxX5x734Q
nhLK1SsdVUgLgEyFz0hTtdVlzz++KCT3pTrZF7UdaOH5Lt7IproZBy2SP6kCPOxe
HqgXLOpJnIzvNqqCk1ZhSNkKyabdH24NvByYeN7Nf5yMbO9tx9D7ywLjWt0bFH/W
6ykA6vee3UHaXl8gZNCpnvcU2zDlXfE3XKAOh0dByGtGshUWNsNeATwagoK8gLR7
UbGPdg3s9iR2y5Pd9Pc1Fyg77HUktfpS7pG3FuGoQJ+ZF1ENNDbGLOkXwmWFg+/F
u4ZTZo0zCRCLA83nji1KHvg1+fJyfkwBV4ezxgE6EVbgVIADfTNssXPH071AYNPd
PTYTcE/sg2qv4A5rFUi8Xd9H9a/j58B1PHJHiQFRQasUZiHjTD1drxQ843mjA/4I
NAnxkbFvZ0B880YVOka2e2t99l8SjFvv+3L7qP4z4wiFfCeZ+IZX7dzVEevWw1sW
OJwWt48YRS7mBjpOTBWIrsMFcvcx0o9NSkpz6k4HqPQwCle1uQSogclsnQYUL1aJ
HyfAGcucA0xbf/XaBcWqp9gfym76eumoYqiExgV6/fLNIaH/FSc2P6/JrGYZbdub
4+SLbY8astMKWJ7vUV6wVwMWQyYRCE+SerlyGYPlomPNTBEA8XMhzDOcMAeZAaYu
79SbJmHldEH65CZ9kpwsbLp08weaFGUAZH3NFFSbDpgALxGCEZHBvP04FavyRDvp
wYOFNCQfAfzzxodCf0DNDXbwn0Awpz67wMJlJiCzZh3rhhqcYv9gmlrS966E4taB
a0GyItkJwcZg/6QNuZyt2XusiQvvzqFUc6nO1AAfCCYaogq7l1VkdGdftKANfcL+
HyorMfcV0baY2ANzDf/ATIeIztT+3N/UiTG63SW+YegshmVDJ7z8GQ/ypEsTnafe
7JqBVnVBl+nZVHguKaLs8oW1XIbR24os+bdu+FuR8nSb/hdxp+cI1fEqeMRNEXhk
OiKi2gXRoOn892eJmBsxjKCdp09Ws3IDiPsplLSKqqAr+A9MkNCSP1WmoIkRvk8c
hqer7x/V1RIVPlP2Y7VniLZxhKf+FbtD9qMOeBMR7TWC4vRLofaG4TMxf6ZDdTEa
/jdsaSwYR0xUD15hXZzWMCY9vpsuPp3326f2Ix3bhIZQzdcv8ne/NZVg9Z0tZhA0
0JdZTYicbcJQAzig2bGydT3b1K2UVitdLvkQkA6oOVZgj0f0mGHQgUpRY5htu2HF
kMD0dTtWaMR72SDtO4OgQSN5Dz56Up8qllFO5CTbLjzbeloJwYdP2I+iX0o5K0FM
iH5eK6IsOMpC1bdyMnrW8GBusmfZK+jkOZlzY64g1dCqL/RcJPEHiJwVh6eDQOiO
mvQljmF969MyZ1MuoQ10KUtGczQVFLpY3xLXLKBJZ0w61TkkT8HYBjaQeaFPrIG1
B1udCtCMxNy+BSRsBtSHBTMkA8PnUfrLh3hAwaabgU1uYux6JYsJvalLqLVJN3ZP
OiPoFbLsvf9aAWB9fkBWL7OV5ysSp5SvVs+dalXRhWyIAHQQ9BKYWKlsWxifWLFQ
lLIbXcH3heJ8c4VTTAzl+bZMhfjgM4eU5aHSSnC/jhdwrrtCyS1nhtJ7S+YtTc0k
jWgJixAfdmbDdNuBI3A5+1YHWqF/zH/KVXU8TRSUIuaQomYQgKfk4+bpZ6KLKNRq
33VtMYZBVmYzhXpXMY565frCIwN2tTxjKWlalnRYEFJXebtGRaLjgCZ02A+49dDo
qwgXc0uK/XcgM9PIGF3/xrHNC0+W/cGKhJzeBWY3sj0AD0P+K/JJRWY+B5qXRkWf
e1mL51p4JfZlmvSt23rmg66QmRe5KPptTcSbRVdrrzvb+9N0U7gZBuqJmxL988Tk
FHPUhjQ/6i7qglg4KfPvtp+gQxBzMd5NdoZtVDc2Y5tKSukjoOGhH8dtIN+76YEq
yXeZEph36qG0/JxTvJFU9Ng2/nyapSGGItX0vU4GQifM8RAB8DBhFO+YdSkgRblH
+gxEaLKm4NzSOCj91JWer+2G8+hvMZnjknsiqE1tNTOFiijpsgfah/ocJO5JSp9N
UlGBPEBTMnKGQ35a2zPbADcTnnV2SsMx7Sww07ud3HHYQlEhhW9R4NRVNDxefgtl
L5MdB877uf93hKsDBhQpzUYz1xSbASt1W/E/GA74KKfmlsWaXvpgoBU19gn1vq1i
Wfs2JJbOlHncoeUsWm49Nwa85IDQmjX8W5tD8zMUt09zlklp03yfMgQSY1vRMuCN
G95UFFc8cVeX/O7U0sYR5+drvA2mm+PSMdTOJBDps/yjr6tNfA2BTr+NGeA8SH35
9AHjpejvbLCkXwWnx7xZMFBlAJ6LuRIEkXHQSdBT7Vrsz+X+LYSSt/Eu4/W5/Afs
NnLZhJXqOEenVII80WwOxPC6n1OH/xrxc7KZubpcTzd9euZYy+7/QmyfMgEWCCKG
2r5Uk3k6A2GTxAPb7zstQi/y9bBtrmE10Y7E3XATMPorZm7XlEcFOm2eZGsL5Pzh
09JGM2c2uxq1YFGM36SFvFbMhw9nYMVLftRzvi80Futvr6TSwojV8iGlXhQOwzmk
4CH7u5xdMU4Qu6RrejLgqc1hncYRoPWvUKuzr+MRrJRAVB/nH58o8JIX1u8uc3qd
HhfjvjoBZUYTQXkxl1vpZyFcuIKMQGfxjDmymi3SxPMbbd47sa0XYLhTYcztKk0+
oHA+ql4FTwx3cayoHnsAxYCvN4jxlq3FxGYXKMabEnDcBySKBovM2iOB8ChQ9OcH
77VmqCBpPF5cxuAYLry96bsP1dst9ZPnmFfi9nlYupOAOhMawvIF76UAIwrUt+ED
L0Lyb6JBU466839k/wjGG3wUnkhej0W7fbQGWvaoK3meoCCXgpe4CGYd6hoteRyl
0XmlRu7W4EYpTjkouBsJucCxEAv+MUVgtan2mDebEoJmCFk6qrQ1xvkH6wrkLEZj
m/OWd0DF29aFttzD1h6Rr6TtyGlwkiJ4zHHQr/94DRvCaq4G2E/meIcTSZPSDlSx
ulxMdtEYG/9XQr/8kU2GCxUxfyalt5lzqSZjeAAIR87iY2k3hukSBh5fzs0gK3D6
lYvxpe+g7G/efR017NZN6D7sU/otEec0gHXbGBnEctfYwruUDZT20I/IM0Hg4p7n
Et6BmZD2q1Y/TA7r61xC907NGJMyEzRsKvNio/JQW6r/HNPBbz2/5b45MmJeVdkv
rXmuFwn1s17APZWONGDTSq81oJmqstweCLdIii1SUOod/HUXtIzVanXxd5SvwLv3
1CYnQJ5jmdtObZPzmCplvwFkrsm1PEZCefO+jDJk70+z3kpdaKwN2NjGMX/66POA
xGDCqcuRuXtSVZ+rd+oTBC8GzBFRle2nM9D+4zfVLqsvwrERftaMtYTCsxG4LUoo
LwC5rKMHhzFESRm1QYQFqcp9wE/kUejOtQVBnC+IQOC/P4/rnoM1k1dUWaB8X7eK
MBCgpcTTy3hpyW/9/WxmGkJcZjPzoVgHWmUqeeXOYDTwXFbdEAVhmzgzHza2I6qm
NsQ7AIqOBgVEw9apXGi/6/45rLB1zLdEQJXkoRxOVTfDm+rMqngIdVXEyK3eMPyc
hKtThzaecmOUs7dVmf0kTiCaLnbjLO7o2aMR/r3qTZCzdnSIhS3XwpFhtQlV3YPV
ShmO/L+X+IZru6bPdJn5opraqMIWgGpMTOuNJ5omVTFliU4dIFkIQAdCzaBtaS8Y
r5TUv1YJp31JWZu2Nf/oO8tMj2NgQtMBmaNql6vYqINLgYve/QRRd/pPFegCQOkX
XVudC/2LtZOWbtaMWwczLs93IMtwfijvUryyLrV1FJJb9qZZR3dlcaTjTCdg5Efz
ehp9MAO3taxvKDu5TQdNK5C1jtGAaZ6NsvaWU3ODaKKRQyIZUvvVDKS5y2V2Vh/X
DXK6WC0yZ7fqnPk+drlyQ53b0YUpddRBIB6AdCdM8yhhof81PvsHQLJVsKG1IoVn
AdeNCZ8gY0iHDZ8q/qNsxWmuf9xkcWhDGHQMzKbzHG52Y+tiW3nCXrQl5j4+Y5sw
vv544H3Iie6FpVI7iCdVhxdqwYlrQaP9jgHAdZb6Dp8zerA1QPt976KfranqCSdc
t5sR2fW7AbUbkppRcxhMld9exARF7caZqUiLJiHAQ8FiQ9Sr5ST8zlZYgH8mxB70
kkNOpvlVs1Emrsji6su/+rJJqjHZ5S0+Ax1+UWfYfDlbzjvw/GXdpuuEZnPZOEVS
Ro/NKGtlEro4Vh/kfblb+4NdENWn69WqcEJMgTD5GHE5wby0te/6EQI51ejRMz8R
89xy1X0Is9bhuihq/6aK6TL0R/v8dB2W0a7kMCbKIlSMzzXmV9QDdYwWPlKoENjW
iVFuz4HG23aI/CfBJRGPD6PBRSR09Es0DQurHFjhZgAvoXbJyv87l2mt6xFiGA2W
0HN85JPi3VUuyo5jRb6m5I1U9/STi9L+Tfl3O1uXAFG1KGd9Vt2eE32XZ4uGaZZP
/IUuLNAhQ0Rj61cOSOcch/3cj3mbeH+F409HVdxcpSbQKoP+vcnN5b3l/34VNl+q
iASXGaYELgvfErzQJIKLMVd5OR9uk0R01NuirvmjZ30JV39Z4whV19ZOHsg7100x
jLbB3+RZyLHi3AmS62nNa3Scj3HpomDsjmNx9/aUC6Bcq+AoxaXkCXxIejWs4U5z
4drS3PUXUSkiDiQ7dUy3U0y2eUQdI/N56BVBeTsHneEBY/NeFQ261p/Lfx9OTRsG
v56+AeMj7hMJrromC8y9OVRGHQ9gComw2iCGHuW1SvbVQVCxlQHfwlgh6a4yG9AH
155vnSYrtQSDWTyKP9lkpcwzIUOK8q6fXSot3GgzMWH8aYeuhRIpCo6TTxEITazZ
2QyqlbTY+Zodg+fK2AymRd+Lfh1/ZPrtkd3zf3LKzZsNv9UNaIv6G51d2QdHw44p
jlp+hpVMiPm4t4W6ESzZ/HUL6H0cgkBjXz3NNvMt6G6WkR2oaZNhnz0qE6fdfK/i
eWTucKeWZr2gVp8ZDee2uonX2sNb3E0L6DBnY28vPWoe7rLPlL4wnY2TxwtXxMrP
/TkRcd00J6V0OBdrI1qcTmp0dkHfp0FPuCtL3p/VNgLZIWeuaxurxGM8yVCgHAz8
aGixRPXoI2ekoVFLT607Ki7Gs/gmqspt2toQ3BMAYAEb0BJKMvzLl1E3wtcZ9W1+
q/NUnALe5Gb+Lsu0AmFjIw/vMhnJHTZAinrtLnmhARQlrmMK42fSx2e/oW0kDbMZ
rXzhZF1+L42D0FTBAx9cl/Thc4W3T2GAadPPcLYEMSmW0m/R7V4McSQpYvwp+0Xe
MRaTv6rVA/64MkAdhMFmswqG0KAYd27DQUM0Gd34S08pSCQXzGQ0+I/bhGj6zaWZ
y3BqUvGmLWlxehOvBN1YLrLcnApi+43YkeG9IC4UTecVYMap0BHZNLSaoTsOJDtr
IhIf6IGyAqS+GcnpLOJuvdyDk9oyNbmpRXyqH114OOGdjsm0Enj6yFqVqIK6WEbP
kORVGTaGl+fCps+sOprApcc8qT3ojvQ4k/BVWU86S6odmFCioM3r1We99q//g4V1
Jy67U3zJ99jsDjUQmVT3x6vfLw3k/OCKe6PTjizyTSrcrrqoZ+rawIJLt7Hb+p4a
XlTp+4dfkUJO5Oc/8qTmYCTJpngQXJyQM90gzjQ/PUsLm2QIDSWvUPjvuLwdfVtn
nDrmuAYE0pZDOvHs68cXmoke96JzwxDuHlNbRVCcsXxnhz00NZpnYWYjJB5vSRp5
UryEsEXPPe+tfCeHFZA7ZS1hiQUZ+bFH++9zKig5RiScCKwEdMl4/cSMA+ges7j8
JBKPBVqdfFF7cf5NoHyVOiiGnbLkVdyuNF7yY7JZGGh0s93sV7vc4BXhF3mBoEgX
DtwtAsBEiCQb3juxuRcYBRYasSyNeaavYuaQQbpKVtre8YAJP//nV04ifLkA4DLZ
HaPAN8LX7qYTB8zBU3BTYIihfDtMb5Vb4YwgkNwm6HtnwJAE2fLFbYBSf8spKA6V
RxbqnC8ndS6l+aLG0E/7gg2BzPAxlfQJT3YOkMXY3Y95K2VavbwXJkn+Rfd90aAz
K1VagmT1vD10hQPuZ5peCagy+n4CkuAY4BqnBn1MXXBVuif5eaajwmMG3s4GMRiI
VsEemLBvDom953fEzA9ezjKr4x4TrA9Ub6X5MELK3xZdycTTCqAnlzLB8IHds7xr
qTE5JGoDZiQgS7M7KxamQKcgL+lNcLc51iCg9cBWuq0sIJFJxH7RO1E8vW0oe0bH
wVzAhdadcdFJuREQyI076ZcHtOc4mXXp9kepL+gD9IWb22MU46J4RaviKfbRN7+Y
1kZGdI+j9G3z0yPXr/n5vZ19DKWZwLoBnXNrdZqGiJ51H0d1mLBcZXjDmMeKQ2gE
Nm8iMiLkiRQ5woXYMiqBh+qmkVXQLOBh+HDSb/mRyE6ILNHbcZ1ytsmD7wvg5L87
JMBwEOIjPqa0SxYy58j0pVitSWq4merBgWHjXWTLzel+/+O0q3kxVxCgGiDJKuW+
IcbJDtBSHvimYwtbMN2spujbl9hiva50WJPFyCLWvMMtxqzSf8lKvLdkH6Szoppk
Mm+ta0kGCvZzIfkj7QScBxZOeTemPdqFUlxqHXJowDxyDLyRFFF7MfzrdqIsraMZ
xHFDnGRC9oSme53XjXzVIPKq7BbA7G0hByFhbBxwukVQ5VSq4xuc3omuDbmqk3g9
4DPDuJngvye+1HYggGFf9OxYqiNYQdznlKISqW9gfx+frLXYXMo0FpJ2VBjOp1Q/
O/Lakg3qFL3uPN6894PIkfw8i+kykZtigGeoD5IaVp5rMXh7zpnaz6tRLZ8L0YQT
dh12HlC9wMHpmW0dgfWDS0cgP9iK2jdsGVPe3685+vt8YdCONk2LLF/dcKSWyzqV
eZ3zC1aFHpecgizxw9ZAXrFQ6/ozEAeIMFUVcDy4M/YJLhHpuqV2XHIeuyTmACt3
W57iQExVg+gj7NRir7Jb8at2ZtNNMQQk0UIbtilqRLwIP7EHn0mjhdvUFIGmjXQq
f1cQVHas4bnUYHvUO5sifMZaQcuFN+wgs8lUExws4bWuH82iSBBrdMad+KiU6a8g
ptamN6holXe3rTcvpMUd/8qxbKeuftX2pqTYSYXukKkUgBXlLGTHPhtiYJ2jACtr
/6gfDyqfRz2jhu2H4UFdRFVknDtfK51gtKmAThIRhCk2x0Ut5SXy4uSo/YR3oKqH
tUm3VdO60l/C6da+8WfFvZtwqgcMObcDysJrPmvrx2P4OyXmGNTYvHWkgZZqC0D/
DVQB8GnGlP7+6p6VZXiU0BdCd6xDBb3dqX0iqv3OPGzN8RUA8qco+8r49VeT1Wqz
V1hN4xKkOseQgNmDMoV5BqTrlCa2khmpPC9RmN0Tzx4XT4j4MvZknI/Lr6haA1N8
UDADcmLpKSnADDvRjk6tXFMIIg6tMdI87G+9u1IWXzNQ9L5wlps5g+bq5C02Nu6Z
IdThc7VB2e+tQQ2dDzIgUE/4Lf7rVrDjymqAEGXNO2Vk3syPo7i40Ki+Xew1FaGG
SAI4yxWylXnIMzRbwNMT5ek5GGNJpgyUqIkmxGWwYDCLonn8SvF2oemLVKMfgr4q
S+fLyMWarBCVcjSGjh0MHRI/jopmKOneCu0haxXBvOaZ0I1gk80R0LWqvBuaVbAw
0aGnIwaAcJQXUwp383QoFuj3HLHQ2aXnzGzFuir+Dhp/Mk4RskeahD3afda594yH
/9kHkQALq1F9dz8Sjp02efmdkz4q64dqGZSNPQbrfqLJa3UZ1BM6P07J+QoX6Tkc
zQiy11Ta9fHaFOHtXOYx+E60TyxrzUAho6E6iIL0RyJQ2w5m9WjyN8SS4V/66QR1
QgQGNkFKI/tJni9l0kpszzI7bFXe/JWVOAvVJTriEPhkqBbZDmIv8LKxoZPHgKUn
ubmg6NUZv24GzP7cLLxDqmJhznfNpbzMowNNq2xgizUrfBFZv9no46w19p9wTYhD
CYH8zVuyNCizYF05Gg+n2WxQO+MOFOZjNdLrE6A71m92eJlFwhxDVEdouxfpkwj/
dC9iZmJVsb6qa3kBbF+KQiX+CtkthYSiBlbqQURiPyZV01w3QYxXOpoeUhe3J+NJ
DVVxWWBagfqg9VCZ3iiPZCHW8s7BzdzlQZDJcG3PGqOlvd+jH6lfd2brM6qkKHx4
V/LgQxqkZ6KzLOT+IMoKvbmMOGw8ipSp/SFcaStI4CEkszqH2rKON1UaFwhQ7nfq
LhkM1dP/5lVa6qC8X3Tmtw1pQT3TYAwpZiocZlaZE69YAavaQj/o45hI0VNyQFJ7
pSZzbxE1DAOcIM0ean+OCpW/lXj/fq2sehJg0wsKhO2retxINZjC0qiDYVY7RYxi
igSmXqtP8qIGm9SyNjrcsXNuPPAo6TxMPXJ44dGMXzVoFNRDe8YGvyz0XY9JJ2xO
a0hm5FHidyv4hiE/8Q6tXL2il+RyQ7zzqzzpSfVShLDV65FpVG9WoHWzcmZU2qL5
p1w0CW8S3sYDyyRH6UIl05EAJMmNI1iWLMrtGfAv1iT+OHPEJLh/JZQ9Paevi4cc
UsluQ+Pk17zjZ0ed0IgTCOmNJ2cXLUJzRVtnwQM+SoDAb2AViHaru3KVNum/jx5O
F2tGBbEr/UbzqV+nVQesEW2rzJuiwvCrzW9SOZGv7tpla7JNE2dIkmpWmgZXnuAW
w0016TTA9wSO9mAbOasTcnu/X0CoPU5I92nmWuXyFBw7Zuz0f+QhuTObGmZkh8bu
yZX1lqOu36MBEjlzVzyZ2IvddW18AypEW+Gkr5jzPBha9MFLIp/mLYR1BbzXRX83
cXTfHAhK06oA8AJIUYVqZza/GmkMHasGQ39O+aetkaUk88xZ5IYGkJnY4lX8i5Hg
x7K9V0kUk9pQwbP6WWoH6TkqNnApr2j/3NR5TDdO3r/s4e5ZTi9DjtjPY3hN08y6
nhskUG14zKcuk3B+uKJwsCXSobYF+RQ4kGaKZWYm+M9F2NOnkSPUUDUsxkd9S9Lh
I4P2rq7Q+TXs4mHynuIfeUHlxjU+SfPQSnyTsHIet+0CRGlOvRDaQMcLTrLOjejH
Ec6+hcXlffK48N7jCS2qCFYNK3L4cb2WEiDXtgbQmHNOzCJZ9NBNnR7z9ov9vUoN
f46mgC3FBAN3qHgcFy7diW0KAZfoPsMgyqIbOmTIBt8INNJUSxXJ57jZ3zLQCVmU
ISzAGVIi4efJ8PxAUbRSICiEMiACfWK1Smlvr+HRdK295gntgmhQ7X6EztHuAner
o+LV9NzuncCg8NcftVbCikQs5EVCCwQ6vuXQj6WM4fi4LO0nuqHG1BCwPWjTVjgY
V9VRLtTEul7gXLIkqYTQtLt1w0mFVBGfd2JjGXf18gYFXFmLrzdaIzHNYteFSwgj
Dgw1/AwRUBS6w4CoVD3J6lNJs6FaFiOgjozRESlHkGajkOZzJ7pRMSD8u48fS9ud
LUnG/sdBvTy9BtIOP2BnBnwy4PKEo3p97TVc0cRrDig3jKpW4/Yb2Qa6OEPA/xcw
yVY8o5c9jGVQAcRlXih9P0hQB++XU0bxChkMENTKtNBu0Bav6nWQ9ureSA0/Uvbh
GWLuaoj1azfjDMftKusIyOxuP2fAXm3elNdoiri8eItiNgHCkN3rjeAVaqsmY/v3
muqyUJBhthp4/iJjAa8Q5f5hK5tQPRHTsdWuVJknIPmouJNVd4ab8OQ+jb+mV8t1
SyIQUamqjblPYTFSuygqO3H4466vBD3LrhMq0+9Za6RIpv02naEDYiGZewAHTbMk
OCYqcH52AGZSCM/V0bvZA5x+o6k0Rys1ZODMBuE19WhY5iWFdhbfyPmdK24DVAro
i/ByLfw03gqUvKCzT7gPlQ69Zk34Ilky4OjxGsunXlto1BOu+gzVlVkZzU/lz7Xe
fXBS7CAT7e7SJAmXXuW4arwjdnHhYKEWu2ApsDmrKA/Ky5fcv5TQihTiD3JDKuav
EMrBMRoUYgaNN28aeDs1Pyq5NeEO0gWc5JtTfTX9Hb2cxmx3GlxDz88SSBuc/5qH
lSOXlhmsCzIe/pe3n4g0AJVq+TknMUBDpB9zmAAbhC8+/IVJv64SxCstDZNfb0GY
8cSzuDljVujYd33L6twqcH2UJ1Qf8D/g7MWXgmS9TWHbA2okl6HybNMgD4XSo40v
0EM/SsMX7rd7d5q0WVonnOh6qpA+XRTJgXFkWdFs4+m7+sLIV+4HM9nk4efUkzc3
F/7PAdaEm5xznafveAtMn5bfCJzqKVFkqre+iCnPb6H/3MWMxxIeXSQmfE1/pCyl
LvNU+hiVCEBM5RQEYpUyuGJlPFS9QCbuW6PErx+5yIM/KQXSqs4mwovAqlVQOB8z
pakz9rl8+j1IiZk/ICtUXsUXwgkMnq2zJvhjKOCDL5nw0CWbW3d40ej39xUnvzql
`protect END_PROTECTED
