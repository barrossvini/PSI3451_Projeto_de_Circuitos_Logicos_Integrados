`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x0v1hqFy372jmixf+W2L8Xvrgxb6YrVPtgEPIaFtUN5n0lbyIE+Ae8XZsBXFjeGn
fTzo41aEYQQvqDlf5xHu3eG4ML8yq6vdQdXMy+IAkV1iQQDnViZPdCpakEr0vemn
JXzoGKnslMu0GVrMMvupGsceWK+jrpFR4hzCuTwTZBkIC69KfF6uyRDVWz2Q6QMs
9ru/s6OlGSM4eKL7z+Ixi1vgC7Z2xoUgroIQD4VeeC+EwZaY6Dm0U3Nw8TveDOUF
lM01c5x3v5JI4qMa0FwU6pnatfdbMvP1nQUBEE/W6Iu+PCjtPuXMyvRwN2SlVuzM
dTx8Ot1FTc3EKnP6XSel9kApaqv/O9xn3C2b8dPCULfzjqaI7qDhzS2QyVJDAZbb
8d9SZkP9nLEcpXyZYFnItK+C7M0DDKN27InlDfRNR+SxRfA7kWVGsFXDQh1XXHWy
pRZBTGSalIQ2HfdjvPBYVVGrK0R849PmGIlNrz0ym9DltqEtsAVBe/tgso+r0py5
0X3DfF8N2Y7sVnShJ2Vsda3JakwTU8JllMdyx4lR9mXiAuY2TlxkvL940B7K2lyT
FZoXo7ZhFttfEhBNqZQ1D7qNz/FhCvULJ/BSmVgrMElRgW9ZYlJ6vmgp9LTDyjrZ
vpkk5KoJt2cYbuS4/bq02/mSJWCsC53ibdfbOftnKoTLB32tz0ro1DaNHqOmHOgi
x0pnarNHA9XbSCqXrWdwuV1Ejka146TIci9C6mTqvuPwjoCWY3jGfZ4Cg2Atk+mx
A0wXGwAi1eiBWTlRudyXuPG3dIre8W8YeP2a7pyCJ6PFLPd4l54Af476pTqJAdFu
/NP7EaBQ4L1lndosvWz+WBs+2oQhbOZf1BMahKKGGHB9bu+LSBcadSab4itY8mEs
6rmWi6BztynI7Qwx8k/4+Z03BxTlhfmjUrC2NIujkw1tJ0B2uIT1SLyr+MpZaofG
3C4ebEVtvhSyixGZoWm4/CH4JyxeX4hz5irwdda56XQqWuZeaXQ4U62tr2GhGlYi
NedK+ltdkw//17VmiL4q5v+GQnAuef7d2yrsYgDE1eEUyhpENAl5TSHummb7JNqd
EuGScYjUdhJjq9oeOcZxBzdzDID8aBRg19E6rQ9nAHaeOsohTAER8yCus8x1J+4y
UwFHhvUkfzUlIpOxzOSlqmy1cX9D20t9PwWTfSn++P2cr7Fk5IQG9yjMUdly3Z1u
7vzwB3zgRUdQZrqI9f9e+ZZjDNpLwLNNbyHvpAA6szfvTeEPCnFl3WbS4SN+10Pm
8mngPLRuNVAyQCEGV+fIT/3LCdw0iP5lEtm+g9O+4zDhRJoCXrjyBTAbWJeFf8Cj
bMrdXs0VTTYPRvCf51w9bX/PGaUTgYA+2uiKsYGhxZxz8mA+jICLCDvbLc87/IPj
xagNaqU9NKSKw/VBFGKBX+JF1xAUTZsh2s53dJ02+tfjAGSP1xTRK1gdzVYnyW9O
mR8JxWNJmdtkI3eWPGW4szFLGkEVdeGgVUP145mCFSFI0/1DuqV7hXsuIKCeeGR3
f9XR/EeTk//B3iWfqSr2mZAQ153am7SpXtKWGCnvRYZsf2M744qRyKLvoPA9K1AJ
`protect END_PROTECTED
