`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MzP9GifSmYKO8XgSF1Li/SRANQ6HLTLMldlLjzZrSDL86QyXLpBIWCEfkeHYzY1G
DLQRQPYV4fsM0Q+XuKwfajfnLrLzSYVykqmO0/N+mnnf7N/q8iH4fHBbCqVKcqXv
GK3SbkpNagwwgQcG39C4Dhr6FtVraW6bqx0Bf9Vs1QEFN1IHVtE9vNSeSCqNaReI
5AB5y2pExs2yDn85X5u81QOt43LygcYq3Kpu89GA5Hqbx84ap/qcgG5gmg1Ca5ja
ATLbSSAl67VUVjEixxGEyTdPeFJeuddbBq8WwLCNanHbnAZlTzzAi2t4ShA1fkq7
iGiYqI64y1BKAUpBoca535tBR76CSOw22hLPJ+d8CJ58BC0B7cD3Gzq3fdhNY+yH
rj1po9iRgPCnQkZ3sRzEoWZhMNKcqXvm7yY0YbHfrHewhpi7VsGLL7x890nVq3zL
5YCaf730q1XW2ldxaqp3iABz1YwKNJJc5XFhU/+b2mfmEzYhVHNRZPcMs97ZHlbc
gpgSw0/gniJWQ41M8EsTy42Qc85Y6+0u2wKi0s0dGVIsrqb6BOVe0j7Q3eWo4Mbk
klH8cLvNlN3elwnZNFDSpImyigobEj8OgudAIZoz3q5XR1iLTuGpRfqw6eqNvqMA
xhYGXg2a8QtSFFyI1xrHiM85zfGx3R7JPspbz7AzWtnERFTq5OBPW2EELL20xBWs
45zHoma/NrdbKX9Fj1LZ7r6IinAw1vJhaM0MyGnZG1RwnRKbpetnYr094UnAcjuN
52Zf0WRVDUBLbckrQHDRxGTEoJ0zw/iRngonf/zkSBiBmcXwwSKvAu42MPWu6o2M
VrCIJfmhXijvG9/SF9yCHJ76h2nQ3Yddv6L3itwVT5ORHvuDQIvYd8GFJSMmXBDc
osymO0//N36/UFJjpR7RdwkS2xzj3iGdvyfv5UXKZL1N7bBZ3nCHzfIxM2ppqGcZ
FTo2hxRkqj6Hg6n5MCCmIliLwX6XvoYDFnxNU7EY39+N5KoT2h6hfgOh45LtPvLG
vLJvK5/JzsMoapXoT2UQ9fPnuXtSF4pZVpnyAnV7OTiWiqS4KHfOZO3p6TNb8qoj
6ZlW7eRgTwucezOH40JcDaX6KooDfSmqM2OmEORHhtb0Nbf9NvIdAScbOhytIgiP
HehsFdiw0Lyz4YLW1OE+DBZdeLjMzZj67nJOJmkmYkxNWHft8APkXv/gkcQIOj7G
vNmJOPj2K8mzljBEHNl7Zm9GaH0qnATzQETz1g8u6VJFd6lAHZLUSmhvFK/wDwFw
QgZcjFt+5jtrboT5+i3E+VMzPcd6svOkED1UmXdxsBdTT66zDQfZmJH9GKxHwOp9
fJ09grN58WBfl1xOipuWCJKzmpi9edI3b4x2xTGJONw2ieGJ9cdgIQyPGV56pdZN
QgWP/iBz7j07p+yPmuW5pQMrbIDHi/H2i7fQ9flmImJb+ROMdOY6NLJzpizdwO1k
E8/ozdoWcPyBiclR3BuOeOVIITs+kYoaFMFOjhmL6/v1wdYzwl9+rn0FjQZMniXe
RISbibJ2lfD3GETcvRKgq0enJLJ7zSQQxbHLeGz++IjmIph1T9Cv4VWi0GqXO4+t
iBJpqyWUWCps0cy7H91R2XEFw7/H9WKx1Jt9NfvxSY/bJkdIVlALw1qi/7WhB44i
qb1FClK5pzgc0SgURexnf6agX027r2uuGJere3d113KY7h+3FxE3zmkpSFvpc8u9
MVXPs6LaQxChYCDtraNV/Oh5iFttOUAL5CZBRZNRs6JWJdOhn2qKnsFX++AlSeMF
8ldv/Qekq+uqLgULo9LUrwPn0UJotnCFcGfnvtDrmr3a71aL5slgG7qEdCs7u1tF
I0YKdNfzcEXI7olbbZyY04pH6qpwFcpB3kORwRh1gLNqlugr7Gy+GiGdyf2PUvde
kVPRkUCI5f2o/QonossEG2YsuTqYpAfs0Xa8QT0ODX8OoGaspfwF2ZkE00i8FsoZ
b4ArHEVPiOr6JH0mikIESX/sBWMgqOA+1Rm8JgwtWSQ7dgO/p8a5n3YQyGWyl3Mw
iZEsjhk8q+LbWxSYHDkt76B2mK0u5EqY2iakN4RhEdBtSG2uV3MrvA19UYClEiR4
pgiANYKZnt7CXbMIHuuVXEgPv4HSkOgECqvvmADHfpXIXvoE2yjxhFGsZ0xuT+E/
RapwpXpmfXzXkgO2fuHR72oVYhTL2QWzUHqenbTokZQpbQb4+RybNC5NGlfOGKR2
wDHvfxnHxbDktZrx3vp79z8tTPAHjntFU+WGYQZTUUAz+OaB2+2+5Rg53Dv3yX40
Ugo+InUm8/ON0IFqUh/gt0jg/g3Lbzy8Np8y+K1xxvRC0VEXuzG2tcmlQMXyzm9k
ogl+k/sFTOUzY98sSl3TVyVHheobMk33TYV5MMVy1F4Al+ci3K+NrPsH7s6FgYXe
S2PKbhTdjSn8hw9wx1f6E53Ln1PFPFZRVOZUFXLFkjxrj7x5XbZ/pl+twLXFsyGM
1u4oQlf/yLCmrh8wz27/OA==
`protect END_PROTECTED
