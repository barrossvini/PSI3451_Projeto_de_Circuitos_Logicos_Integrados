`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
91gm4cDWITNwYt7YmjetGHm+KShhbk3yxKGgLxJC2Z258AKJPBOzvnYDnYM7Gvus
UAK5uCPuyitagpksSEN1B7Fxbgij9yUw3Qm2IK/MnVauDaiaUMEiyiW9j4X2TpCN
D/HA+d0sIuohwDKmjNKeAHEso1TFU80LJ+xI669v0hQdIJiR50q21qCeb4GApg4e
C615u4sW24NeqngIgkvwo8P1c68CVHuu+ZYpiuSRYie/OYZHl9kMIGI7KN6+7p6x
91AdiCENc0CAX7xYFwq10G6Mgmnz6M/DxcQ3sRZ6nenebW2RzKrRNPZ+K/zywkc5
GnVXgmJalHRSiUebR+dMHM1/eGxc4XDfir+bS+WzXGD13kHrMKaDfpcwlv3WBbQm
IhPbkrHwONd+nIebcVf6ozWXE8BgvgyHypZqsV44CLqrKLcSMkAEGohgE4hs28m6
JChljnu7tbCfmWcFY5I3NZUaSEneFr+0p1nm0lHXiRm1avTnbBcEpNeYBhNNFD7o
bJs0KkVtZCFHcMwXJy/rL9ee94/ke3Ohud3l4/nt2D1IlWjzNq8G0Ami+shgFBqF
npnAFW4QNqFOdBJiak/+Kru9muxKlXGtgEioakRyfpPb9m1hzHiMiopLw2NCE+tp
NM1DlSh1l1YlpzTZ6bYcZw7bcMDYsqlkGd2Dfv6v5byyQNtZVDlDkGQGEdeeKhrs
DeDG6SnERgr+9+/5yxjkYL0z1tXu+qBenJieNrz1bD09kv7snxjk8FK6f+zkILIw
zEX9804YiBxHAwu7lh7NeB1E1GihslclbMDW8/WGb2wY+gjIMBo9hetWex0PUX17
k9tUr7ARS3St/FocrncVXzjCHHZSLPaR/LKUuDHXkvJDuB5GtbsheUk8yuGYyIzc
53p04tpEyuuVFgB43fTCQ7dZBuzygeR/qvcdPsyYc8WTxeGMLYV+UgskJlFERrJq
sNNNnRWKj1jM996W0rKXjjCMmWQFMOFsKYDwEQTcQ6WsxtOQ/Ecg9jDxnvgUpSf4
1a5Lz5NWVoxKbWXKA/8eycxfc7xsCn2J0u1GZaQrYRU0+gAlu7oqlAPVAgYzwhXz
t10atC5qN6ae+9saC86PVyw0I+o8OWCuYPSGDOrYElpf6Ggf35kyikHTDaZZsIdV
BAkaqnD0n+eo/wxQPEDjgOTtrnzvkaWE3TXdag2N5d2dxMWjbog5ZgDZR8u7PM5o
HhhpbpffYcLeK6k1cgOb1ZH8zRNmAfxJ5LY3dn2vmNVFcnksvS07jA5fWxPIZaKj
7sFJaUUMxyxz1QBIvE02mgAZKMuaVCBMA14o7alBc4QPMFexjj446CQCea1WHEFZ
vL+anmdI/q41i6/wy7bKtIfCGxWAju/bm/LaX6EMDpmzrFc/9aoWg4CjI7OBCnmr
v5rcL9x6ljhobcYpAdYqJkn38CSDiCUT0sOVyBfNrg2VSQ0K/0cANNwD19y+HBau
8QQBpVSvt5/RJZfXFMFvftNifndmgZ1I5VHFMBg70qAt26F10L7weQtCkhGGmJnr
n0p+GUwexbkZGcxCfaQkxgSfYbx4HA41QK4jbWERSpW7XQ0FDH8IDG6uqQRfoOC5
1EaStvntw6hjLzv3ilV7Ff1BF5tV4GSM4gA2/9oZXDDVeA5l4GbFMjKGVqAhxoOO
s0HP1mK6zN7cRdydvhGu50+xcwcKaJcjXCxwGg4uVFHB0xPRr0rEoSpI1bS+nshO
q76kX6ZiQdO+hme2THB8anEBEdbuWntKGe9ubi6UBYAQqtPYhIs1KWSi7FBl1zVd
4cQR01ii1fVw95px2WxqGMAZ5EResLQxoS9BlbKR5IyWyfIgzjlgbR35JzZU7+dn
y447gdw08pPhlB+a8Phqapyz9cYhf9gZ8cwwQ84Wz7vghbg2DaZiQJKXUw0vjnoF
VqAZN/Eh1sBKzNf5pEsaCAhi8ZR5BImM7jQM51ZxCtqiS/q39w0lZbYeQyG18UiC
hCbPMf9VUDglRpZYSJ5vAkkaduYPMhdmsI3+DeT7tvv5PieEn6LOKxKOAXoO03t/
MLW3hjeHnY16kIClTzcs7mb3RaAfEbBJJYNOyZlctfsQ6hxv+SxlScBITTp4YJUC
ZncV52OXg1z6C5i9xYDzZjeEwakQpuJpVIEB+v1or8oHLTuNUgE8FAhcGTodiKZb
c8Gax8VK5RVtCZj2BhWIh1dRSf91NKwhjKL/oKZkmPH5hu9psHtjwKHi8G6c/B4Q
bTXzSDB9FUSiNN5mVb1kYB2uCkfThAxphUwE28WhSRMwOofZSTSvcQ34bxJMM1g6
u6S0LeuhLvGz0dtHtdEPFiJU7VUu/VW9VntcCN3EFkrXxG7pmoY0BTEPURWTxgJm
3Z5NDEeq5qPT/bO5FTu7wcZ7GisiLBtNGPTALNPkkiPb/ITkl360wt6PCzmqhWRf
W/eijWu53NdrQ1/76MBOUot98vr8lqzUbe+04xYC3aaZaY3CZ+s6e0VcaRoiwCLn
jDyO2wikW15fPSp7we9Oz6/P1rqWdrrjPGStoC6rCwpVLbi+ZyuYzA9UYARMUpJe
9xy/Sisl2ZAsz8XInMYQ4mg6VExbpaQ1NDk+WeFGxMIwdFV8uDF8Z1wHXkfkJQq0
N9xuPlWr4O1tZv3HnFMhvkBqoiua2rcMa3n1Z03rcihBzBBYY4slLhFZVQXeKmtM
JBVq2CMIZm+KV5nhRfy+4jP+M3IT82/sAloxjVlVXHBU/OdEyrnhAiTIQwuL7kne
ET0dJGJ/lIbRs6skWkOtOjC9YDIdVqXgdesNFmx0VoM8FVEakQSH3fl5sdM1gKel
51bYb35StoG9PmdzF1IEXKrFNhkn5+c1sj9PgTaUS1Q14JTkC+qD717hP8Kttaup
AThmlI+c4K7DpIkkx72+uT5XD1skX+OhSkFrtPThUmDc7NcAgF5FItauQkXymVmK
k14nGItDqLxgeJUh4m/CWDXNiLD3c38jsnX+OBrxLVO7wdUG73AUf84TsuU6nAso
ST2rbVp53jshtC0LPG5l/KHWLPnb0FqFhe+f04A62Jr0Cl9FTzq1aEoIeN+WiKnj
jikeRW/0ZesqDgzxQ63B+edbloejmiTsIOS2SlAgS7NPHhjQhOssRZzDt2yzkHeo
Hp9NBkUv6oY7/LxuX5dxfI8oM9TZahOGwcVkZS1K8A+p6sUNwKwGk+fDt26/BHQd
2S9Bn23b2BFt23dn7Ifjg3clUixXxmqK/X/PLI0smBK2au2LvBWdhuOGwhHNiMEJ
gASLw89jkMYOlGgtPrkm5Qex0mTJNUe2yWfN1RxzCIhng3kwbIT9cl47EqyRe1vA
CUSGgXNqGM3wNpxRGGBQgmOKCRqSwFyQ50vLFYkWllsA6k7a8PGtQId6pxQCWsMf
Uq90cNrJG0LnjyRwYFu6JNwOnRAIKtmZ4QGYe7ymTUYUA9zcqaMdBmOcMhZBFGJk
buK/nvIFH7kjILchfZOU9dWhahBrsi1e1owXFk/UKwUedx5dljdHUZJA/pKFWS0x
bug8IB5F0vhR5YbzE5oVxrMT9TOorZXJ+LcNyH9J8v7D0hbjoXS14jv+4Pt0Y2dw
WN56FxtbAcocTD165lZeisgLpWl9CF9ydxgiyZFdJzq8P+gi2EceCbo4NdCIzeQc
7eaxadZ9bTkAT8s1xo2KyDLB5lrS7UZhL88XWwUyqVRZr6wjEau8O0XoJ06tPQQE
Z6fqaJww7t3Sg96jCcCbhZGEf9y9dljZZWcUH4rz1NdCjEHdbuy3srBi0Tmp8S8t
0ewZG7cC69h2dgLhKx/nf7P/D9lAhGnjFTN+p20d3U1Rsqi0lW8hEdhFmHr02kHn
U/Y7PsQpKw1TtxvoRHEgWD+9R/eHgBRTULBerXcLadl5vZZXJRGxlSJbketfdL+N
pm3fAZecppqBRze3kv7g+sxwWQEMIXjSc6n6nKquPXKL8xYewGF+rNOkW0nWpCJ6
e+i4Bdn24S5PX9Z1fGzYUNVipjXPMC9hXSLbCbjaTJJveOimWDb0yMkLVmhUFPjz
yzrw90MzBUudy00HLzOpfPiskLkZvaKArUlizoKh+XZekarzjPKYn/7EGmQRPOB0
txJykfOknprxEfvxuctCkzUfgKEPiGuke2gPMgKtcnTuWUnvosESwxL1itHlpiAF
j71JIDdBpWcYq2quInENbKHNqXWGbXsdf/rIWXqOiw4EGS25M216wOAgxkZ7QYz2
dYbQfZsZwuGU9JHXkCBAFBNcMKrRoykesnr8qCjbAbG9AILCGWBySjCZ9w3cpgxQ
oPNJsygI9PiyHVhT3gZ3gxB+FAeKY0u5z5hdGkPQUujpnGQ+6wjdVrMTX2sFYt8c
Lenb/xvbHCMHkDPYwoPaT12lna1CLvJI8O9w0Q9r0EQO2SmUTzGD8IctkSlAcvNe
6PwaGcxRUaztoUNiP7KpmCSHSUNjozVL0uIXElQvwYB08sMAbnxRW5yobhpBVQWl
iDtdELzwAETwz7octHZSp/EcMplIxFox7G4DcNpB9ifOJ1twOds/FIYzz6C806SH
8nTjy2Z9G4RlMinNMeu+Ymi4bSM1xv1YBBGNhPPpYTCGyLPZEXx5rInktbG97Ia8
iMhMDY92WTwTNkpQhA6c4lXVV+9/CJxAGVqlRfbggOsVKEWu0tUWWIXqDw1BgmO+
rNBrwUL+tqZxAbPiWIetpBVNc/kEEL7tqeHjqffFiT3BJn4xemPAdaQgDWBFF8JP
Yt/e6AZGJV+agQLSSTbeq9bcz49zbqU+k4K1nq+xeXhvt+6RVzQozDD2DCdyHQDC
bIHD43T1HxJYR/Lz0LwX1bSP9vi5guJj5HWOrHOKkmvJ0HRkzAoW/VimtrPbiiBk
wpIiQzqCKR8hThTT7TqtkT/XbFHgQHwsLCFY8Zi8GKxPJAYYUoBjoghOveySh96M
rw4bdGb/22t8SWc7HdfBii/A7Qb6uhJFWV20wCp6U6FlffG4+y3MrLJkPav3jbmy
nRAsC4eJbzekoSzCoapXCxRbgdcn2dFEJrRzGeiQsQ1EpMXoK1IGhJkT+vrJWZye
ublcMAePIOwfSMNv+p4muU7APLJV9ItsFpaor3x1tIPQMEkl0AdmHH0b/7Yo0zFf
h5VV9ntY8B4u1g/yS7mUqm6dwN9c5NNEMT0Hm6AEZ5oPflyVYloHwdOy41b657wr
lD44ToUOqSb2/lDtD5R0FosHXtNspuVk5uLiNFQoovjnSgJZl8FiAo+lshwq1FfL
laZ/8CiAQm1dKlDh+Y7qqDP/JXpS//oIMii8elIhGb8OewSasgIP1Uhs5NTC5ksg
qO7T/IPuSqObLYzq0S4iO6380NY14r0TRhNxHe3e0ByaNBi2i7MkHLB3Ns5gttNR
pkttf3eb7l2q+clH47le7MDBwtMtWHpB66eg7wIZ1dFb2z1QkwZjtjtyXAL54YFL
UoCoOE4mNxxy3Wa45f7MRkQ3oYrkahsCH7gXyKyeugCKzT5dgRP+eGIPw25TFztS
qlIG+9n3kI1e6dYgqNE/IiLDDZL2Yig9gsyd7sGhw3hp+BKiNtfyxZ2foUOFZ4I9
krz8GbIWbo03dfz6+rmuYRYjaCX6CDVLx0gxFSj9t5aNTLr/XKskjIUkQLeH+h1h
cxdo+Afyfp/QVL2o5kI1zG5ktxFsIFJ9sH7rc8g3f+H76ykBSXBbo9Stkt920UkC
dZindC5YPDqWJTvuKBGS0ZuV4lr8Nr3eku5QcjzKhr/9qhQ6LYXD6HMK1Jn9xHkT
sVhnahIi0epS6HeObMRX81HtmM0fVeA0ne5UEP3KaVqbuVL7AneRCigG0wyE78Cy
NKhTEE7iAwDNzwbUPweHeqVL5iP4+wfRu6iFO99AUt0CVIXdXcMZ60Q0k3rWY3Tn
hcn7hUCfoHmZWult67HSx1HDYP758WKGnbdK5aXWyXMiq+trs9cF7Tw+G1STh8/x
Pi4mYd4x1EvqVw0govIKIXe+5qMh5MOv11nJTeOyNEBYttJrrU2US8S4+M1bL46p
WeVleBBApcglwJe/pmYKo8+XbKJZmKZxeeKvv6vMRFFcEunfO9wYsCPLq8euyLmf
WohPkXrA4JlaWiyBi+7XS1H02wb3+am/Jq51oX8QUpvWZ5w1J+dv8kULPRUUahEw
3MRlyzJL67igrhvK4aeFoeetioJ+221jDsabgfan+UMoxpGLLe5rTbar7Sl8OW8G
SY9xe9zJomoTKu25aBYl2En0AQj6db3nk/Wj/q96+GR/V0/78hjVaSyKzWlLdiJj
QbIqBSOrLkgJBxtyc8UX133cUnxRAkL6BpZvalW/PmW0MDTrnXPGFX9fuQIUySDA
QGg+WszViFRTCnuI0ZzSi/nAWKAjyDFXddjXn9mfBFTSMm9DclqXectOiOY6j4fI
rN8uuPCMNsU6t9cpuv7rYeQd6VXGsL/g1YGTgwXTXj7hSgBnIPD1NZUe+oaogYBc
MYmK0zrwTY14ZnYPMKi3iXBHY47aylSIoN+psapFjEv3id3hPypOiCGhYmTskEDc
xv6hzdO0QtjHZwbOtz4KmAxJNzMSbEs+7liXnqaDp3fvi3a+mlxM4rc1XIC5SMr8
r7vpDwvl6WmmZm2sVammpB8JPXGV8KZxhxsbk/DymJgO+3TT/TRqVch9KX6Hu2+D
wBJ/S4pK1GubaquJBj1bwp1GhsHavzUnnBxziPVXqsGIMkIMGkbyp1ucuykdO5Kd
jOpijxogN5JCWG7oPa2zLrdcww/5oWrKM8Pmue9IVTsblMyrd4EzglPI9LLVW74t
O1OuV4uVid8RxiIFvh6H2z/LNkpj2cGH1hB6r73E+OUZ90jpqQC0Hqc7NUcvmEzP
iXazmnpXEBSfWnwe6UH09Xx8xJ0ppy/kT6wV/gXnm8CeEXfHhnfug72AK/xbQKQA
6l7SNZVIrSZq7OPPptQk2un/LavTvKNF9bWZcOHNW2u7moqybkt//QzQvkSrxsyh
gmnkxNx0HtQ8ojnRr90DB1hFCoeVeQg4WD10Atmu9QwdgN2UoCPKDQIxRUVP32GM
5fkQ0T6hZdF9BerikdjS7l0Y1O/ZZX7oOd8he4Ipa3F5VnEABcjYAsVzV/MnWQHN
/c1pSsHPEtoH8ke5yep/afKR7gN4Yztb7/8O0uIVHSH4eDGXemoUbi8Jp9/kxjlB
HOKYDQLAT24H8z+0Eg87VqMuaaT3Rmmqv8BOOkiqzx2qCmnsRqbaHzFzedAgXUoI
kFv19oS5Lu46lwO6Oj2IioG50mcbQddSqPtoDBps3229PpEC6QRqIZln+nXucoFw
Wu4JOfgspFStGUWfvZEmijWpqdWCyO9tz0G2Dc2/1azT6QwVhdXeOXJYSxih0Irv
mK4bB5G3TUvMFJ1l67DXXbE5aJIvspPosaVMRZ60HpN2Wz0SSPWN9sJhcRS06Gvc
NUaTdRIGNpVqz+zhGdk1LE9c3CIXvqPGcjimYPcEKu1wo84INAHpKv03Mg5rLSmS
FC0Hhq2qbowqNuj6EALDP4AocfLDdQqiaIPLRG+66kqHVQdVMykDpBfFmC6zIxvk
/7Bst9pDGYh+LFT5qDqYi6Fyb3m2ej0fCPDu3TM8naV5+09hGSabIN7eaZdWo3G9
58LzbfPEoVE+jXENsdlnzWPoJt0wQ677xjzzgUZ7m9p8wDk5SrobD7T2gYK24dZ5
xFj3cDpwMj/1ZIZZ4qNzuq4eZMRAAaTntoG2Kz3iuol2cul/UgAEULt/lsAgjw8+
pTJgVGmxVwWldGTAiZsxMLmQCXgBrodkxY+5SHJF5YVeKmh0J2QKnABofxIRmpKy
6KFW8boul0q5GDLBbgSRjmY/q3NfoI6Uhs4EQkKVnrjlEGh4m53eHOV1Qlpe0PJV
0J4xvOxnyGHFPnR2AAxJJEpytJyD2UJ9TxK7MYFy9kTKhMAZumBHgnrItp2iqpfd
hSEp4g/PeCpMVKm6EJ8DbT5sdTXnt+hAoR+w4E3lHOm5l3Dy3Ehwkghr3uF+QKgU
fnouPAmtR8H/jNrIgL9e2s36aNEATYMteUo0e1fftPRrJbjJA6pMip1ZxKzXkgTT
blxT/hPHPev0zstJHVLx+QLGfQTnOPy+LTouzXxhBBLAYlSwbROGZGSrZJWkvwaL
rWZYI8WdRoNhK/Xx0uG7GXX68shGxw1v2vbADcL0ElpURYCzn6t9YDD9GSVMTTzZ
rMKYirQs77NjVOzae7MNJgmkAh6mLP0KAtP6w8kmTnAJWp/PKQ/ucam2L1zevVZ5
78YAnC5zkHfr7p/QWJkQC4MR6nXjR9xIG6wgx8LFoHq06b7lciDzQ3YN/OHcmijf
MgKBusASAouXiIWpe6SkYB7l/1SQ6MxzJ/ZyeE1F4NAX0aErEbCoswQBuV4SvBBU
Qa3Yvw0jAEqqbuDm8kfDkiNgz8lV9iIEM1IOJfRzQEC1iad0SnkVyxV3EaN8WSor
vPYPEclSan+3z43RzK/Ah8GZfzhDf4MhV3w7t7ybIaK+x2CamzdVqBeTP2/tC96Q
tgCSQKkWFr0JweWY6zlarLn/3fMHSw8GDGwD2edg2IGD/WQQxdN5JaNUpeuylXP+
Q20JBUR0dUieh3L1FZR12g6DMDmNoiQDvX0GT7LSACBkPN1fJwA6fcuddMdt93b4
bveUJBBWSFPKW6pn0Q0GivYJgKyie8DObiU9S90bHAvSfRq1lPvybazip+omlB9p
CTPRDmLCmwSgaiG6FdyY4ECCyoXfwBX5AFM++oymoP7OwTektH61NxLDIsRD/54I
/+ZHyhism+0VkjNNUypwWP+/EF9Mj4qAJo6YaLi6O7oeh8WVVT2lGf8pv9MHMrr8
vK3WKYZDfmNvUi0Dy+rjlfUoPpC58e+O4/mkmE6ECWMcu3wMw9lMuydfY1f+nV3e
/rozoLgqUniXfVoO1pdS2NC41CHdIm+Pv5vYjX+7Bh1o8NKA2keaVZlFvljhG+Ib
GsUF/8rGP1omwv+tf6xDDal7RI5ja+7nrry+tTUuOavyL4mIzjo7JwlDnHXQudsv
YT72ucSq8aZ/G/E9hkyU/YhuHbxWM2xSc8imG5Ak7lbJfqbTx26Jook/tnsRBBU0
jJ2PyKtwOcmvMFsn3yvSPe11Z9Gt96sQ+KgEjQj2+e+kd3Kj4dg02qkjUhownK8W
QZNEJsDURvV+wTJpBddjprEFzj8W0BWucbjY91aBibxEVbPcH0QBQ+FspU8AWnLc
NViNntE7dCiZjfBwXYy5FJIsBHfHaTavY7PeIEDC3CylZmTW+DxoiKGGdRF29sO+
CVrGjm1HGEuVHOkvJy7SGsGiqAQW2SHFS2vaOyDOHRMJQvoFj8Iy3mGmSTYicTK2
raybOYkMujudbF/QBYPA1dWBVrPkgT+nRq+R10P7UZ+zCrsZuYQJ5BspYKf/IX2g
eiwsWWezTW0afm2iIMMlWeoYOizRDNFLLDxUIp2O7zhgQ41GT/DILBsPvHUjSpC/
0dkbTWM0VQkvnq0UWmJ5W48GWCaZOTNeXV4NCGVsT1VP9PpFUs6JiyywtK0lMiXY
z1ZXm80YfvVTEE+35Q5MfWzqUdf6sOIqw2idVUOWk/IMX/W+/zhAoLQT6eaDv8sS
mzKCI3Lj9wzqTkqMx8f5/JOQhlFYNgEJDnWZ2ckTWSl4YgWbga3CEx0vYTt3TYw8
gR/5ph6GURYQV4L85XmW8ojhII/h4SStIqhWbQ4IhXc1Skuxz+Gfqxl7MuhwnyFk
qvmMKw4SFZa4vYlIII9d1eRRIGBJOAZfNuDyIkt5VVusaPW9WfrF6trgmlrmY7Tc
RyQPz7QXLUHZYHupuw3U6P+DFvkE1SZW3AcdKRNtmaRYFiC4QVEOUKpbDLIT1MVp
Rg1YMs1+tPESAqP/XDLHxGYUs8L1PzYW2kJqR9O3cTQsDsUAOfygbA3L4J8ObnAu
BiMQyuQbBcO0g6X6c3RluUPusiKg5sYZpX2ZpITVnwwiOXJPrGv64nl0FrhhBtyO
BLqUS5DO/i2jS/KSKfvrIFhBGW47gasw3GJ8/7ILQunLn4NKkdvibIpGEVjJQ6L/
vwpxF2I1jrtHde5PdR1MY+mx7A5CVWIwQGAH0HHZxKUxp/kEaQrLCEhMR4QSjbxc
a4kpMaPr9B1wUuxEcOpTHPCoC/i7gjYKNLW6HZ5ECsayMfCR8FSKc7yOhuj3kh7O
1cKyBPZ7vIvp6q/FEbusM1EZqE9fBLwoFprtb0eVs8bGQIADMvi/Pb7KFOk/VuvU
6UmbzUKmxMz/VUDg/9loIV68lxed4XOmFyYAz296TOZowxMc8sYsbbQ0ZoGnl5LW
OL6jjFOnVx7kvN/qT2pJCtdx9c84rSZ8sY2sF3/Uw4tK9Wz7zNmD61QSOJRVgMuK
qz3jxZM1RPfkFyQB+B7ZWjuUSOPVd6m/QsxKPwjMj6z8iVIsuHSBx12KEeaD5eRd
W1lACxpU9rWmWf/2nOkuBSp7lBXftHoH0X36vDNT+vIA0neJDjeQWk7vdzfPRVDe
b8KDy/czZoO1K23wywcSJEd/4SylL8q+mAVwB91EHHNcS1TF7/mIyBGUPxhDMnEk
L1ZMF+xU9qCjfSnaccll9fy1+1iqUIZgJuLrX8e/MLtZ1rxLrPmCkIqOgEvQt35Q
IyhvTwa2Buuz0MGRx9x0ARs2FPBt0q8a+jslWeULKWtTxNDyX1TY1//dRgfqEsiF
BwtuHTNG5c0JFrH5wqzpgkDiBxYCLqeex3eITE95ywxAs0ZVHRJKkDYPEkaJvJaR
k3Eq7iynlJnE4lXQi5wr9F3GNXAhIe6auFPXdy8IqN7CC2MCOwwWIlseNDjtgAuD
Vhvby2BF7LXtBmjeBqnJyx30i0yoRtTY1nTVBe1QY0LiuZ2Vc1aGorFvTNhjA8oG
a1Po20b3H+sFTfXzj8Wc7IBBfGG65/oKNgyC/pA5XvsaCNJPr3o71ekI/Ds6Cvcl
Ba3OMkqD0pnqY+aixEbGd7AeqxFVGKTSu4EmOp0QauEEphgRQAYHBwUgVUa2gkf4
Jgp3W0z70yt0cEAseayq07oF1O/XwrWsGQrQezIUwRdLVpnHj/bkQiJyVeXm9fH+
IkF0yAhRV+tC057kelAsNpdDwowAfp9BHiBOV8Qqxo2IEOL7lz/Fhh11XWW7EygU
TS3yZfr9jaoV8s9ETLC0ffF9H+KvkOINi5kxd2lNBfizv5f/X7nMKsb6btkE+BkC
0WhJ1dQC0OBMKzt4w2Co5+zjMkHBE2/aaukgZOrfbFr8K1jFr9eTexUsnhnq62Wm
ZmJZN5noi2Ii/fTzOo6Zaqra7ZxVKQwNRGJ/udvRdgu8IrB01K1bKz8giR/7Kw14
sVpx21k+Uoh7cbkPjsJjemgVM2rlkX6ySF3mifUW6Ei7ngGZuCgCTUviZQYdwmsP
3h4ouaRhKEeiW4txa+mkVVbmXlMeUOXhF0NQ/8d6na8wLMmctuSfIrxp2MJlRGfs
CmUdZyGVRQ0EhqsvvGXTeur3PMC4xkWa/9SVic+rPGhfkHQMHELPYl1H6KDy0oTS
RbLoi33CBZ5NW8waba2/Fgx1I7qJztIAbhmvMTJhcqfGG92po8GF/IYd8JBAeS/X
fkEDQQsQjLgbEi50RjoZKF0Dm1fvHTJeiZ04gCv3yHIIFuvRfKx0pQZwA7PlpJ8b
A88qxo2oTydhDiea2WHuqauOet0gJxQKyXYHk9W+QJHxaVMCsEUxa50lQDVx91aW
zflqzVLlRLmMi0ahPhyn1Oy87phH7K0yAFnLggdIiVBm5GI1jd6JM5zT3tc9l0zE
tl/f9BZS6gYCD2QEGGE3DSVRy6jWtr50RCp4KEnehywzpk927eECSjmj/2FZlLfR
yUlYueUgv2hIzK1OCt85Ieu0d5+a8L730xZwoL5BV1pM7L/3VhMitrzoqMBM/TT3
i4VaUYHOqucrsrffV0UR6LrQp7D9TAcQjPbfsbX3m6mn9E5PnMr+CrqwwonMJbat
RcbkKUF8m3mrV2154G73GpMaZwmlIqTnmmadGBXBEimbQ7OzKFwEFpIbXCMN2FDo
rwLzsOQOq/t/CJAWVnmW8qNs2qGhUm2S+mQI9xc9dgh8i9D3/5AdHj0qSKtzYbzs
LOb1EfQ/JVjylfkEGiUguel+SfkDAbll1wKOJWT6bzYs/g+qkOt94IqewNqluPYx
9KDacpT9+EbqWz/5SDpWx5tBjGXA1F3Iprqr9xJxYLLcdVLbkne1JYFmw8Kdm7cP
cySWXOKB9XG3+rSwX/zvPE+kskDrFLwVWPiK8xMmIm83caMGJ0VLnd01CDI1kr2o
FVlVy1KZTSJaeKpCa637YkZnGa9xPFa41pZctAU6j6Z52mRrTg/tVNmKmZQfmRM8
00ne2AT8BliLiKjGJBxMpPgvvXtKHc4N3Goy/Gloe/ADr5ud5ewyUAhifLQyE68l
ah4wcuzVox6A+67/ZCtA45DtJO0k6xh2zqzGqmgSV7q2l9ntcwJipUASUPzWgaeY
D537CQIU0sqhufLYmKLsTwm++p2qr119F62OWCS/AYTFsBiW/Nr0d65anazZvxLb
/palpny+mfykQcddry+vskacEobHEubN51HLVwVHu/4rui3V/JD+GS0Ya4uLJX8q
Uf1dRf+g+YFP/w9QetmM6GgmIyWjejwDHtEfyrtbxnSOqv7Yds9kh1/G64pRkcuk
uEDTqGm4SggdtZNP+d8Ae8RJLfbI4d9Q/mErIFD17kGa0i9RHPDvCH/hY9FLEGMm
quaeSXpvLW/kHu1SY5SynLStd729dt0M3rj3YpHWmmZagzrruuyLeCnXsjwrfsva
wD4EdWCpqzdjrh4z3TZPJ6QDAPXh8FZTBA+Llj5eCAKaJdzZ24H3c7USqgkIgmsY
gtdqfZACqdFwwDMT3Q8VqPpnQ/8kd/FojigxhA95x/8cwkKCbwertNV0Md2f06c8
Xcv0rnqVYz+7xjJIzyZm/b9KLXHc/WjPU79s31PSfwMCcIzZulTu+vwvIteVZwHk
IPvsZmub45cppkIu88VxmTyEHCop8Ck9lS9dEpht7XaToq80kWVhTQfjDgjHYyKP
OCgDwOd9DN2pB3kCr6o4nzcf8qKwb3oIKh3nYA9Se4m81WUNxPClIZZY4XQNovMn
pH8/7dvxZpO39yMKMiZsdCUjfyklf6BtPMJiJO/mXxqAXsOA0qoXKxIfBoP+NtJu
SfhEzrLsGrgxJ6hOpeVRdBrkck99Z03+zwAUjnbQmcb4hBnW6mZbluH4Tto6If37
kV7lybA+kAqvJh5S3JnpFG/smL70grIAI754psm+bEZM7CZP2UFbzXalmttmi9r1
m0gYVNaGQjRhjtr0i0bWd8rAOsBDAyvKUhf9rjv3D2XPEFHR+EaPHRYnhhXrwtdc
wAXsaeJ/SQ6SonkNCI30ix31yu193B8wOAD5Ultvp9qAx5xF3/85hpMdYVh/8dKK
Z87RWEu66ByBx7rIQlIr11VFfe4O1GrnzxXc32wn6prLyzapVK8BUSCz9iIQA3vo
ENvS7r00kNTxPr1MFSJp42svV6iizvcoddnDOXKMmsjB6h62c5FFRsLcH4bDHWNH
paaKUWMxjiBSNlO4HKZyZpHVVO16fdsIVvs4Ffp6I/DQr04N5YrnyJiuhSxbqipm
SfTsJBItaFXczZXyTDbaFJAAeJMwZJHh7GEsCefeDE0UIprD8L728dUH/zDfpN2C
c3hMwhdwYiaHFfrpPssCr5oWyv6AHWUrL6ey6O0XQsXMlCHrNpm1UW3R3DOwajiD
4dTMADcwjtVHYjufB9NF0VHKKMVc7qBH0nW0jYSqJlWyPjIp6wpdlGfoQCiQG9Hu
1ed7qxiRJrv5MZ/dRzIfSluUiq5cnDBYTFQ8j2kJga8G5ZEXCSdnPLVmhPRn9Ekl
myOUSsKw657KE5bdmt8oIRovo+c+jVXLTgsKXnswInVud60kPfr6XkXfW3Aje5PR
yHfUFdi6UttMIzQex43SRBpZMotLEsYDoO4UMS38GfCwh2vaSByUnDYRJ4GDZh+0
e81xt6C0QbfvjzynmHpU9QykGS4njTpRE9PSNlQrOb/dw9WspDMPoixkzUf1hppu
VSQzHXOfOwlfRvJfti6cZ/gt7mgtTOsBzfxGIdNLQKa7x6XDkbi44TDR3hb2CfOe
TcNHmUk2ykXi2O3Mdbv+e82bKtQdeukOGS2Jr1Wdo+b9/0x3emD4ySZQ2R38Kpph
zwLiribaBRORAxBbz5d5oxVShAZNkJyLqbQy2tNb4HvRI7Pttsjx/uElLz3MAwCt
MfZt9zAgaruiMyDapUOcFN3UbGHgOViFm/lhZaJsx/hAPgk5rjjXHaD+5eYU/IBQ
ezKyBZIF0iQm7/22fMQK+YTenowVf3O0ymSFJFhQbKIRMK0piO8irPGfHV3tlr37
hC5TdDPYsTj0Crjuepj1r4gxdzpWrm+xeCRjIW95QmjPbYzOu2rJAqjRSxuzun1N
LLMJlIuyEAKQXV9iCvt7Wh1ZGKUXwShA4UbbBPvVHZMyNlRRMMqshP9BciJbcT6r
yXBwheNIaXp1YDrleZGoVeU/erUE66+stILWcbk9vgMqF2s2r+/0UYTFTX5FKddp
aoF9InOirVadyhDUh2t6sySb3dw6/Um9wJhLtcqxJs9QjrvqFsNXyd2Mp7bp8W4a
ZJmHUzw/TJdDJxC8oHZlODYQibzfV31vVwBOlHmcBmjEZtbaL0MC6jhgR3Ptu2+9
Vq+qnYi0Mn5y+sUxY1QdGRQgsPOn4ZBkWOXauY/B6NG6WI+Ja/YA0X1Bi0KnlPWO
2avz2Yh/VkwZAjnJdEHm4W+DPQzzdf7nTyyO9rFOai38m4SVWtwtj9u1qc8K6nDJ
JU6cIsGSP5mNaC8MqkaARLNTMTu+b9PzMJFG42Osi0GzdGFfftl1lIs1VoaUZ/PL
OB0Nr6Yf6vtOMyfvhLIRZVXwCAW0qlgGSKpgxUYN/BPFKEu0S5HPVOgQ08WfiHhW
sdqHAhPK1WqgfU7ZsRFugTv8qFIGrYuQJmnZRlcQgDOAFms5qXhqg35AtT1h0QAA
mLGfGoFmFhpTy/ytOdixL6XuMfMVuz9q8rrcF7ZyDIv9qMZMdkojoeG4lOFN96lw
59UDdlo4UMyvS5UZ2+efxvXE+LKue8OW7JMu7sktAZKBJIX81AiGLT0r0ymdTXsz
4I8dVZBiw7CMnTIjAab27NMqLIRxcwy/6OFqa6Z7HIiqVSVoezowWoAlaIn5lNmg
PPuH51k1y8bYPeLz/1jSIyioweswcNDr8UaSB1sUeY6UJPLtlOzgqvKFvGEdGMC6
qycsv9G76wZLQzhlwgXN2juO6R0s5y4H568AANB8+6kfHCC19CoI/7C1nLzO0+Zq
5d92Akxf5BR1SUS3Mcr3N9xDwb7CgkgEjhNhTQySdBihCX6RS6+7ohUXMIovB6E2
CjlaP5PnWZoshW6Hp5fb56B+6DeQtP0P+4LeYB7oc5pCdXwfqKZJf6kCVonV2fuY
1K/QUqEnX258k84JiIhSeElaKWJ8kNHMdYuKT1BFffSSa2PJvnlmtYy8nLEn5DSQ
h6GcJdS4z609SZ2qC8+r6X9B1kQ3B69jRoJOEn+jnlXTaVWO1kRcFnHKETYvWNi6
S5QhCx1tOJIt5KQUtXevhvK5PASppR4dBQobxIB9qoI09Slql0kwLPLopYXqjA97
YUrkH6iQGNAMxs84FNLVU0wT73f5RJBDk0yqk+bjlaxv+xHkIQFJBkJ0LE/oGk4v
2YklTKD2wYt941adgpLO1SjVECrn+soYIa/kouxCsUC9NYUeD4vSam7rq5ZuJFm/
evVL+t3s/bqovkHT9VwcOAWl/45BEIIEiAVr0S/2NREWbn7759g33HRwbYIX8P1A
LsWGvefGjOPrveCvJZrnSo1dK9BQ2aKT3amLsyZY4cuC1RtuhFRTQvOfznVHPCgQ
4sf3x9FO/mE1n/trXwkn9KJw5n0zM49UPzxeYlLMNdUh+ucUrq/dH5RgngR3kEXL
NAO0YbPn4Sn6Q37YfWtWX8kW2Mh6ByP8N0B+4hbGs53dfMst3aGuNoOtpH7HUHVq
JNKgyc79vIlLu3+35gIF4sCKhyY7dTDahoD8aO/q55YUlY/jFGAog7CSKlPH3bhL
tW1QAkPz8OKQY8bdcPW9IelQ9bNpYs1b8wsFD1UjtGwDNPZdk3KQvzbtR+6kvSK8
w1nAmtw2WIDIZWW1/AAFz0V91PvaAzZhVSsbyOlXxlsKs1/KYaVZrA4cK4WcgxP8
mVmonSdZqYkwlPPdtQqeSHoE/0eb/dLrRxltkqNQrcc/K/mBhSbMUAn2saCfgJBT
c7NZ2wTnB0YqJM9IV67uVFS0BfIIMb25DhM/Cbgec1/5L4vGsf/J0ylYfXCtkrHN
iLKN+WF1tAVB23SytfpPRbBnX8ZTbnebKzbgSyBKGHmyc0fd34+P6zySCwgjIVs0
UnWhFnWXnDomcnhXhuuPSSCFRNosmsSeBLD7OYVGnlrqlS+R9v72Vnz/Qm+TXRTN
jetcnjpTEJecQdDvbxdXhxPeTjXT8eE0ntLyVP+u1BfprvwYamrhosKpfJjKRSWg
lqsKx9nKr04N8xC1UGIi4y8JlgeDbqNZcEz5IT4VJ68fWro2baNWHrn0kZgbXziW
LiB3drhDS8uaDDoUh4qOfgjZtaDWPwn9fPqz/jFSvdoGOzFLRAKG3vyXGgRxvJiy
v4ZGvBC4nnLzMEXZZgrToar2X5H0BDqXg5rRVcosjKZu1RSINEwXSYw6EQ61Zebz
J/UjdwU4BCv1zfoi1JN8DYFZWUMepDx4fVAnJUGBl5xnpKL74zd44lx+ZFPi0XaH
pSG97+VtOPeogj7wXh9siEaTfQwZdxpWQaYzN53bZj20IwkjrILVZzleSnhG4P51
hw1DHcr/CEeOdG4RbdnP46lpqoX3wGdfx8w4t1HqcfRwGzJ4P8gvKVg9Db2ueH2+
ZgcOm3NZXfbgo8WX4MCbMZbyYk4P9rO942jQB7R9G1yujt23t6SaqeJwwfjmDgwr
eA7hkbh/M3n3MtKAwUxNlmsynmjfcb9i47tAbJea57FomuznxpDYl3abS3HYCmkU
8+nOrBLu7Ch2z7+Wz74l6fPvQ1Vqr1HIyu9D/qNuIEN3kdn2DnIG8HVGEQ/cSfuV
lvGhU0SaeCwjhfpqZKHYDDETDx434gTK1n8dam8oqXsrKfN5x5FvlFs+GsXKu/Mc
pRDvy/xk9aQCuDaEuwc0OZqQ/h7aULd59tNWZl0huOyWaG/GMWfzaheKKuvm1jvC
ynnw0j5gOwKqeT1aEhJ1yA3FXCyFBLaQkgV+pRSWWtQnNleG6V0ft0Ovv23E238K
sv9hx2M8AySlYi628vFth8dw9cu5dxumtihzAZ1aBpR1e8gXcB9lNulMbB3nFctG
zx0NN+l+UEipSqsLSkjFxseCpf8XMJ8SOqRrvQHtu5VnBbv36o5IXmCdaajpyaDU
JAnhLlihbL7Dufq++57rzOycxUPFU+h2O197/VJsvU0GouuqkXZRDszS/lhx0wg4
yD8g5c37Z4BwqNWkx1zjel4Lg74adfCNI70Ici/48da6BrTU1rkybr4GuuyTBZz3
YT53DFCb51+a8lgxwnZnaIUEWIVcQ4dtNXMFuhe0BrHyGBuR08S3fpxX/pWpQwzt
w/qm5xTp/oxzHanQCOrssMS6oDA6FAT728pkhZstNKuBDA1tMw6mhes1REXCzZSs
2PwZ9FP1HHfdjQHB1DcVAEBHNMRqN53ZDWInQMrcLD1ihqsmpqyVjmRhNvWR5qRi
X1fCGUWQzveJbIkL71dhXzYyRjSRlYeBpnnU9LDllfQ4gKKhkaBLvAhIFKTi39Dr
Fln2kps1z77rDQn+2L9NLtDai0LZWg5zObE60+VuTeS0Nb48ClT077JXFem9mAah
7V7OBTPwp0Y4izotNVlSS007j9N2yt8p8AnfIELHwyuwa4vXibnNcXotiDhORciE
d4B0Q41/L7ohX/B9uek+PNmv/tRXGKjkod3RQRK6gW6UkRH4I6NSZb2cU4BI93qV
AsZBCEUK5voKrg/0Re355G8v8PPfMqbXZ/PiYSh49HXv6iuP7RO8bIZ4YDDGlTip
k1IN5qmQg86G8V91U4+eWW+Jx+vk+x9xLlby1sMve9KY0KZHV7za0OPCRaZut5wo
WQxYwYmJL+thdXyEj9Kjys72sHyH4uhAI1QHHXOY+y22kGzM+HXrDepYxHdMO8jf
KGfH09j+KXAS+Gm5miSgI2I54R0xhi2l9FMvK4/qpqHjoTSQ2SIJpBHfs2KeXVgN
8CbHzPJtljea3vgJwdU11W8g2hYdPvRmPcc53Adsujyxji7E0VgnbJgq8LQ3IwQP
dX0mxCuaN3IeALWM9yEU5qMBduUG4guTEKDFJXQI3EEytIcrkl9a5MAUefje7voS
ckkYI7wMoAp1tD7Ki+zKwWcfXENbVmltnpFTxvmQk9R5SzZV32P4uOnq1+JAyVIc
qQh8GpcVIxxOmTVwQz/oLF+HmETm2p4/6y/aSdqJiT5+mZ4XcO5BamfZSTFzXncS
ilI7ZNHId+v6Et/+e83FjmmRSyIUtfVYOYf1qLBBMe4OlIHjBKkGGZaj8+aX8yaJ
ACeSahQsgQ0PBgMaqXsoU39hVR4g9XE3zQYB8tLNaxRiP+CgXeClRNLWG8IpeKXj
0kav8wtVEdDNZD/eNqMsWsxp3Th2sOGeHy+abBC21bEjStHTgueHJO0rxEKM/x1C
mJ01YrV/plo8hQgXQ+jlf/lmiktPXUg6AHkIx1e5lafXRCFAcTL8ruHhDeWbHAxq
ZGADGsM1X96hmSZ3BSAi979fxUsm8I8fK1n0BOJ28pHdzCqY8oSOJHbuBJogHRFI
/FxwvTTUOSTQgjvr72CnEsNxi10OSxfNDAZzGOakVEFZnCF/OY8TfR5gyt0VLZNI
kHu55RjbYBZJNQVO9ZZlA19SVyZueO1vN1r7I4T1RhI5mkTTt9ZQHzrHRcTezj4D
shcWZeMrRf/oQP09riksm8a5vAt9PHvbiHK1suyYALxR0HKLeOTkKPQ+fOLEAhsd
MDaNytSyvXWyfB2JntWJF5EKnYnsH8EXkOk5PFMrmsK1LRA2j14Tqu9r/3pgAKao
Jync0XMlLsX2NgjGJ8vMyGjJ484ApcbRwSMS3oVWOnYpy5ja4VEsr4O2Umi3y1U1
Mx4nEKZFsd0+bXllEavtialhz/2VSTQz+YwHwsCqZKCiV1HYeW94ZoE95CZlyoM0
7r7erCYH9lGAbbC4j5kHmS/qzFKTcO4XCRvEyGuw/CUGPp3VyCHhF/QDOZl41Vrb
KIfWy9HHdSvmmSeWXutQEiJB6mzQw0oMe18cOogVupuiNb9UR45fCKDgTINv2K+n
3UOuQDIeAnzA4za5NJegcOYZ8tpYlu/+Jqdcl54Y6KSGeAE0Z8HcbhPXMeJrMOq8
WeWx/gs/0G2L9TGP/y+TGnoWbX6hARwtsjqbNxcTS10hDQdP+y1IQluXJd/QKtWA
GQKTKrGuDcEVoEVvCN8FujYZg6PPN5iG2lM0J8I+V/bH4hx7qsKrZL2gnksXVgy8
cJlVX4huYteWhgt7ic4pU7f24peCb70TaD/apwxvlVbQPNWEMbRR2Hoc/EoJAsQk
9/7QtUPJZynU+z3W39DiXNE7Fnu5/IU3CosR4BX4Sgahl0S1O8Sv7RU6z2N5CIVc
E2+GEmpEyqbws1AN8obSdDRBn/Xu7VDxoZk9hg5m3UHNSIWk9kOosF5+fe9dyL6K
/y3Py5dtLj3r0VvIFZQrvXswyMlzIm17SPQyJQdaBzwapAI3djevWDuk89H2JKTj
Z6F0pNOoAOI3GKdlLMWu7Ast2u7ZmNlamRA1Ul24jwmLtpJRoRGhstBWrVpMe3hS
W3MUKbUbmrw7zhdc66xkjHdvb5A57NBf+SPtMi2E+4bbn8W4mQsnRjLsnT+T5bGc
4OyIrVyOwdypONEF5ElGqkXrZcOl8u3y8KUjQZ08EWrwJM3itanLUdNhuYRZx0ay
5wHOHFXOGZUPBRj1jx0Yo0M5Up7C2JY7t4LXzZGJ3ttvy7dgSyyXS9qbuNiY3u3M
FuUJJLxMP9iihYDQ2wMrXLGXb69h+jzeQ++vfdV+UotlOYAkjfJ8rnAwS/5BXPj8
H8xhjrdDcPUEaigHHYQhg//PgXVc3tRg5niFsByQRHqpIkbMvSdNMgHjdWSoeqft
6IVX2Kfs49eVvdu56cBfoQ3jf1pEBbUeBJ6xLiRkbC+0BAcQIan5+GOfUE3WYV+h
P4col3ZDWfqqKiZn1vZ5yqj25Vmwbh6oL4Vsny0yhjeFi662x6k9DdUFxqz53iB1
XkzMaemKTWrIc63yU6CmYEezyMZktwrFNYX1dvJRQe3jTKEwAvRvHkbqqogjOuta
SqNVtAlwOz1lICW95Y7gSp70lK8SxAfAFpXkz0A0fiFkheiOSTcq8LrlQ4kZwd04
nys3EItoCu6S6d3uqDZRZvMDee+Pa/ra4u58Gfwyr8CXCniWfEWabdTSXRFawiEK
XUQtChEkHk6LcJucqnZeXbocBSHETt/gBCXciCHHs0OU/Qp8KRzPspSVwuuW1dW3
tP4KwdEnRgR+btjoUNvzLgzAx8inFGTQ0tDetJbH5R9zPWjv4MRM4ZnO8MaEiWte
MZqUShuDJtf0zKevOfbPxgtdAy6UMcznuuacAr3yZd53WpMIpbM6DXEYNBM83H7O
/zMrTC11eYYrclUgyejKtq5k05XMCL6uLQzhodZPoZjq+nHyz8BmaNz3/e0ZLMhM
tGz0bWQg1KaqA07JO1opW3NY/Jt/x3Gy9NFEYpqdM9ja1NexU3Dxs4h/FwHY9gZC
NOOVHVCqJdC3Zv8A3aH2BqiJAM0YMS1c+GsiQYzJEfwF41nZ7FbeBUJ1RpS5+LBL
+/NNNie+Ibw4Zntl6OjdzxkT5Y27ubztNmH9oTsQh+iNVOxjetapAx2K3yebc0FH
UAqEAXILPkxTFa73y2Lil90HWQwN4In+1mB19lt8O+1U4jEfwVqBldRG6fd1ZAof
SBwxphOimxcDfnztYaqLcodcc6SIAJtqzCfGOfh1i2X60P/fcaxpY0Urd6he7btA
bA+MVACIonDLWGB2CNmzi57Q4LhqjEBlsrO+3lif40/cWs6P20X1ONp90urWhMCb
RLRp3Ej14XW5tOeKeKIZA/Oo8M/s3Clf5LxMZHCdBINLc5yENgIFNfU5egs8G0bL
RVjPX/Fg7TyKaPTzTEpZ8fHFA8uTMoXzqU6Dr91cuZ9XRFxZ4gL/nfetW2G5YQ4k
7Fqi119XcHw9aZgTD6+41s6IuYY7BjgMPX9093rMM4WW61l7+6c54JCaCdUem4Fr
2cFYiMDMM8bHpXadhnwbFsp9wnwXJtJidHxNnd+ii/Zcbr1OJqn1Nx1btkrFNOHC
Mps0ANrIH0gUHtuQjYu8b5fhRgVXI5oKr+dsQZLHHdI0odpbzfJWsTY/CYEI2ZSO
D0OyrgZpe+8qoedsySP5rSIEs8l3DxkfBIjfElvBAN/+ImRVAffU4FZDN9Klobq2
8TNgv3+NcsBKMOOAkHtAliUhJ6nuTe7u1ybO29/mDW4I0mJdtTdSrlZHByL0jIuZ
TtP8+kdhReNjKyWnGa4nN+sV4tOulE481dLNGrnDE0tDxIGw/hNJUI7K2MgPe8c1
DYzh0s+3dJLu7HoWG3hDQ1/9Uo0DFt8ReKO1vRclGrvbBud8pyt1OCa/xIUJb2Qi
ix8PGwGrWNESP4ilxsHyycrUlFn2KIu699LBKtsgyO89SmHNNat0+kecw9BnfN+P
9ofuQQKlfKSAY9sGxCQf2rCJ7RBhWQZODs2uJLrEOFo4nU1dhxGkXBgXXpU+qns0
0JIFAWouQbRhMgDGEOt+d3CmNh9J+2l4GkWZHgiIMo4akTCD+b6o8XJPC/lt3uhu
1MeqGKgRC9XvV0Laxf/a0yCa6I0MxhruT/99R8O7JqOl2MzdjObtb3g3aqcBqj11
ek9UemCzJX2XRI4qs8PyhY43PY0KOKL0cPCbOoNVfh/yiDE+qKWkNNEVXe30fKJD
zxHPc07dOiU48bRHnIeYMy/8Z7uj4N30yrtzf4Wudfi1nWPEZMp3U76zcxvjWlpQ
VPcJ/kFYMlhsUuyd6ecTN/SX/bUVynsQbsduZ+euywTdDHeAjxh76GwURlkYaNjU
+46eyttqpOtb5fgkbhfPKxFhwii4WAvhS1fCWbGdaHfiNcSlryfHT4uZM3GERYUJ
6E6eg4+n7gW/zR1+t6pTsAd3th2IZhZIRFGa38qU04Pti9O1V5yjEsm6+ZYDNthL
f+3tCZge/oBINGXnlTaTUUOgbYkZAPHedCBAgOpFxB0YYrg8QPS8pBqyiRJjQtJb
2Dvj1MkQjlwcTeX8ohXHMTyQZZFvpXfhRC+8cVl4cpCjmm8/Yy6JlQz6NcupEdEM
qMlNy8mCPaUCTmKkE/0mk6uwIRoK+9CvQGmojs+vaXMm57skDpOaDteQkPVXTS0L
r1/MebPUoYD4zgcvXkdQnS1TQbsl55Cz756Qqdk0BU/zHjHw3JydUCfouAJHC56Y
IeWFdJyUD27FEDVXB2lYJmn8lFsmElA83zBWWX6xhQaooNrWvS+Qc6CVpAm4LjiG
zDIZq2y80cwnFLcUvpeaC8Txc12I9qgJSjb1CejRoEuXk5A3Jbwz/Undm7H/CDd8
Z6He+bSC7c4vjNTQLD+Bi5UrZMByAoOE5+pi+3mFRsktH8mkLooq2RC5DJw2sWiT
uYfqouzzie4tJO6U19oGMVhC3/d8knI7hT1Yuxy+p1I1lk5112no6AjnLF+eMa0k
UGxQ835Slaeun/EbYW52ACMG5OJDEBtj06OHL9PEoJYbbaOKNqndmTqyTRASRcwR
YfWynnvzgEc0VarBLNOAN8NRwak/YewKocudhGbYvjFWZnFzRzoOFYcmhYgCGALe
DVaOXIYRNdxZF0Sj5H084IurOff7n/ir82KOxkh3L8XAA0vf99pzOLJ6ItdJ8JWh
S+BGR5gb76wt+lIownwuF3QnIYzFmAgQO7rvaefNziCC1qH/0plQOaX71l7qyyuV
zFt87jbpi837GIQdLV6HtGf70hqGpMnOZnZ47RQCpDMSa6Z6aIbv5uSmvTIqcY++
Y9hiZOgXnB3N+e7CV+YkGQUK2jqJ4bRxoMa9fM5DuOAjC8xu7cNjqTy8+gEhuFxN
2stndJGwdv8O+ac2ubsVCO3TnX9mA7yUlt2RUHjBLPu5NajtgkckhcmUEm9agVaL
btkxDtqPBTR4Udkc1eHwy1RzV9FQ3j37kJsyKSBdKhSigJe+jA8GUPinM54Kpddq
2d/JCeF8giGTMVFTgb64OpktgpyYiNvHLD5dZfkqhm93/ivwzePX0xlvgBN3HpMn
8TbEQ3p3JNs3gFAwolAKYDE8KPqzFzplk1Lfr/+XXXI5PswEpQziqHIGH+g2apTf
wvR19q498kP7L0xsRjfBr2WH/YO2diqlX1aDIN5BiJgkdEgolxzcGYE4umy3XQW5
jvfIg5Ft4xIpGo5WnR0kBKDnULqDcXuKknGPK0cySFd1NVrnPwlEjFJ6aUB9+omd
b5ReTqFNuhlWs46i63+yu5zR7z93mTD/U+qr26dd7RUFb2/txGZhPrMAB5p2lFYY
EeHOSV37R4YzFSr7UmBQRa9tBY/VCwb9PjoyOckPhx97+hWp+Wizhm7tPcXZvrrQ
qI7niCD3grBTguQNolMjsDGyGx2KuRnnbbnc16EJJ5aRr7OVHiNqinU8ckaiyQJF
UgAGPEXt0REMfJn0Z3zlFlk/cg+xMO7lsZC6pSpQqtymXu27Uy9rHYzF8IwtLiZL
jfb4mZpjeLAgMCls/5REM4uieYTVj+Jc3aI0JvA+ddWiZPKFp+6vf4EPonmCIu6F
OIKXDyv0/jZ8qe0Jq2XTSDfW5UBuI0JV+OwWBAhDdmb7UT2q4qkgzJ2ReJF7ucz3
cPCLzfcJWsYtilqWjmc4YUyvdzbodILFzo6v5ib0bSWEQL3HFM8XNLwcSjPWZD4q
g3pBkPGQy8qL8Kb75rKzlx7AmaQuXLcg5oqwV3P1QngHqCSzEaSQqcJ2//0k1Own
CN91DxGxBb9S4EmVH0y10vAnUsG0c8Aws3BuVYtAYGJWwa7UsoQQXzYtS6+Xy6ae
RCXa98kOaPm6ARd+KIxF72oTTLJbJ4rbGBYrCtbZy1fjlluHweW7KXJwz0vhgVxV
B670kE4cYGJfQ2kIZ/ZWbClxDKGspbK+VW//S83tQYxIXhGoUjxVZrsc9PSRBKRL
YROERdeMbH35ah6yaWEPDketqqM0yK5+0MCw23yfr6v3L8iUSOXI/uSy+gVa2+xX
fMbe0JoXSB50WvmRIXPT2m4tHRCZBWTIw7Usz08uiou0ztMOlav/oQ9riIPACgNC
KuYxo/Je5PMEaCn4vlSGAt4q8A9lh6AbJpZZ5AzWP0fakfqjuJCOFuX3vzOcTGU4
DGoDd1fE79iSLsNL09TUEyghbU525TJ86dwHnlFus4ANEbSG38xVKFcVauBfivcw
zPFDpPaZzyPF8WPhDGmxk3VE/Z7MEAzhX8yH9eZGTYgDByVc0BTxgZ/4Zkt+QWHG
xhpWkBH04nmKczsRHi41Yc5twCIvWYJmwEu9ZRHLlWNa4xATD8KHjRHhJnuHVJ+k
PcFiCL+SLvGEDyPASSfAp78knmKWLLdVJdlM8vwbl8UgmhIlGRSdzSzugG/ssKIb
HTS5VRG3MuoBCCOWEa4H6oWebE3UkbjLd/YxCystv45mnyvt1NmyQ5BeTvSawzMM
VQJvzlSMqY8mCYY41mGKAuCobaHw52wlRykeLA8UomFjuoh7e8mqGchZOLit0Hdh
bDnWNILKgurjJS1NKrBq56R8Mgw66V4lzL0M8qY9SZY4PSmRE5WoBOp5knF8r/du
jOKUHCLMPPEc7qz8oZPHfg72Djy+eJDsHuAYVqpZLN3h8s5r2ZGkjz0CWJyvijNC
dFQn9PR35msrwwkiDJm1sFjpBFpLw3Gr3OscgVfbs4fX7wrhOc0bSe8qkiLEAsvY
j19yfhCqbbfCVyWSqozRGQUihpUNe55/Qtsj1yavdjsLcoH9LwgREDKA0f+fbcof
cqWq+242p/bJ9QntxZHByT1bV5h7XGGzdti6wdMEQv6cH1SWEBBOjg2ewBunUK6b
ovoYm1VeFBzTa6T1+OG7klk6fY1i+btbdkpp4zu35uZSDkH945L77hZY6zn0RHgs
OgTV1jE4Al4sAm5DZkB5GzMSf99Dc9k1mfqOSJwE8qjiQV9Be9L0UPESzvQms0rn
NOD70yCBtWVsIwfggE5e03qMyocfJvk6ufzEyislIGXrdSuYrD47+FchZPDfZKZr
gHv8Yzda7jrO6x+OXqXvy8A6tpod8pn6FNs7S+KxTKz9nCDyzvdlfF4xh1jUx24c
j3aQAXBgvkBmHZWGEigAkQAYK7vdKsR+r5+BI3ZdfQGFHbAkzy7W+uIJnN30Nybx
gey2JPqE3TRiwa45OEk/I5/0uQBmYXRMezQ5Z+kjWpmUNfT8OsWqKo699Oa5WjTD
iwlugzN0V8/FPKmbu6/AhWzSpV9UDOasK+gAwnQ+HtEKiRkCxMUMV5060zp/az/2
B86KwKK9aEdNlo+MlY4VuypFMyocadjEX3zdGXKYncGjqh9xqYPW+D9vGn0p5b8n
2ClksavqDYhcFY8zjDO9Yt3Em7It2LLGm/j9zQ3pDDbJ8Yt+AJyIaKXQ3rS5cd9q
SID838bfMWf2d9z+GON9MByyGJVPCwlnrO14e8PvFFiRZAJmE0qo2RD3wEAh5hQj
iYZDtBA1MM086A6Rou6fVmbhggdawiugUIVUZEtXC8jVNhjckkVGkUNc8Eb75D38
c/xqaH7plVvgRIsuw3DqtdLlZcWqW4HFD1K1d+xv3XqsF9FpPNUW0U+bpXsCJ6jQ
9BodSsRcvhjqymN3MBTSbdWZta2QvVBXKPZFWNgdMBpJhW4DeqIg2ilns2h2Zd30
JYmVrT3bz+uNxy0lDuDDRK52CpywCl6pObBZOsGDjcvcCin8QpZ6yV6vtZINTmvl
ugE+km+FSoT25T8tAQFuQ9yrupKducZoj2mK82snBeyXpiULEc/yymvZ2KnjmsSN
fSkFk+c+NOyGt64YF0IhPCWJH8ZTJcs3y7GOLyqNzrAftUpGDwZKlNl6+TmPIBg/
qN1vvO46glYa0kUHdEEqXZRgU9S458bm5u7Fcz3ZmRMqINdDw6EMmgALUcGaRH3M
qIgjwqU1lEargmhlE8v/OOlnV6g1E3xctuSl9JckYCGafyGbJKC36dM+eU0mxvFN
Vxxjuldxc/melT//oQNbR6ZXGNUEWy7vDYAdPYPyzeGwR9hct0UuCqCtdiTIs5Ec
afiYJnQ9te2wxKE1faZpPfzuo6eS57ZRCEYK5i9U8dbnDN5Cu/KRYXM+isFEiRVe
+0h/bOiGvqNqeExGbS0Qeg80lViO4snEdAtcXnp5pgP2jpnrJ5HoUHjwMBw3k2/y
rFXx5WFkOG+NvFGjoXWydXZUjK3TLF7L+G2FSCI/FBr9jiU9fFo41A6pDrdo+/0j
qZJMcG73GTO+oXiJPlO15LHF9IdmP+jQ0TnDx1qmKBTDVhii8n+o/pII8VbU1QPm
CJWrLfuKr149A9ZxXPeYJ1fOk3OTnG0CTvy5hoHYUFHvNZH2hMj6dc9nvHS2onsa
xtYq5IqWVqKGyD8Y98uKRjs7Noryaoeq+CQXYi9VG3xHaLPi0quVQ5qPNyMtygfc
QEjSBhadxy5p50yveynj8N3VdJe+2YCRQOvv4eAZV0zmCi6v9UcLigDc08yHlUym
2u4vDsDu69vVLdHQE+TSJ501T650Gxe8xTX5guboNwnkIIN0TzFEbYqtuqpmX6cD
p8x4t0t1bPzz1J8fqZVlNq2FTYG9+/hdu3lE8BA4cC1Xm4QJhJ90ALSd/lmoGcmn
TaUIilzhMO7UNj9E7OrPHdFde6zw1NVqwOtIa71reJkqMXGi1P/dUrPXo8d1BLtf
E0sTjcr44zOn0xu6ZHkSvl5GFE8p7TgGYZpVg9a5/7x5rosX8aXXV8i3XI0P4JBP
13dFFDwMArMQUXPqAL4EcyNpt/5DdAX9LEUU0NC4NUXqXCclmgd8cPMMsjY4Fwam
PahY0u/gUEf1xpjBRmb538yhtSjNMyi2ZV0m3vbY0z9HkNoQK9gfgnLQ3dutSujc
YLEDrrkyMC3NtWXH0TmfWWkoWNJig37hOT9lCBn3GBZmZR8fao7axI7QKgWmtbIj
TjkatGUl1KzqtKsnfcXpz/swJoEwy2gQ2HUASAOnC4VUjYzJZ+5QqSALh2sUIqWl
exz9Rlh0tbYr4OB/kCjO4NahupOfrnR6NxzwzN5rSdyVeVx+SYtiDxrBxn2HdtjF
Qwg8ZVDP5IGQfG/IDJCcxu23kZX61dxf62admwLsVeYYPOHizRyv8xajETp//13h
3GcTS7CjUWUEuH4cfpIq3TuR8XuXiDB7N0Tve3X8f64LgO1WwAidNfCMPKWq7b2/
H1SX8Jv8Bc/4ytl2HuAdTeQyHl8J6SwwRS8W8UvfVO2pFqqtVSyTyJ1TrTirdyzy
QTDcJ1Ae5NU0q9oflMso7iMgdxCvcRqtpGGsUU/cx7fXIybCvXEn4jctZsEIv71I
meVvlNPQTAzJgDZLW0UAAnQf8AeTLjY+zEJjF6Q9PZYQIM3r4wn5Jy9VSQ+QSq+i
VYfuX0Ib4GcC7LUburmJne2aW7MWDqREOU4YaUAJ/qH0tH+R5HxxkfhFjApfFi0Y
ByjCaDJLrglkSZlq7IaodSimef7R2p9suE/ub9LJOmO4R6v6yxFO8pO6Hw0isFTL
wQvuKAletp4wHY3ZU881zaPIT4vlEy5s7H+MZGQUZX/loM0CPtClU37qkEcjSjMf
XmN8ZJ/FFlx2TPpueU78SqVy88P8DA8tbLj7v7HnR65MbnFuoH5BzGPPT321Kkav
EQce4eZFcxOT7BrJybgTU0UwnfBxJt4oyvhoVbNrwIE559sL28tIcR7iGTqMV5PG
aCxVUh4UoCrAxgOiGIw0j0PdOm6PPNppq+MEj5YS0mRgJIEt2l78VQn/qKEM7kTX
oP3Z+UL1Kj3d68jOq3ieqhT79Vf8a9kuAdXpbkQ7tA4dJUYQjEDXAx3FhnniKleB
/2ZNOYvaj5HJSl+RS/EQ9ZH1ZsxD4UXEWO66X0hLDayNssV4UT9hCdtqvUiSAnNr
fRL/le9MFpRpCDOeSifLPU3alPepUp7m4lJMitVu22SqTj4fHZDOUn2Zj5jNxlN1
g/Dha9oHgpCjV/rH/UJaNx/gs/w5bMcekJwhv8OWnkKqOVpO/EcQyoOn6Ic4kXwQ
i+oo2W9CRgVY3aeS81g5IV4zLK+hZ7WaQBOcITeUvxWTXxiYQWrdwyl61PAIA516
wiC5Sxedvm6XBp1CuIUGaxF7DnfKJb6x1FCbbdYcVXJPU/KvibPynt556psteTkc
E7LT5PB9XLR9J1zW0y+byMv/scLjyoR7gOwU5bL6aF9DG8bma8e7jYz/zwgKP385
pS+dwFxO4VN8rTCl+TVXIs04jlhExWzhh2tPXw5sSebkHR3a7+lSsJRXSDIYU/H8
5FM2WPyXORjjXobI7lwxmw7ZwbPxE+8PlYnv+fukG0a3Ps9ixtNqqVPTc0DFy2RT
xNZvYDjXxRc/97Aad0e047HO2cYbuuCqFdactb/Fazd/L1hEDGINrraPnxUoxgdH
OkB8ByXtT17O19MIfTWlTyPAhgj6DTIUNxskaCCHkbRLv7dAlzDb+/BJTXqFTVzB
HYa8DoKWT74gqtLIHT7P18qj+FK5SKZVuKBrJ29bnW9xrIvNlkuKwP9VlCZtKubW
vUgSNP50dEQgUhnoOHtJlWaeN8UdF1RbEpJlZR8eRXhlBWNlWREJ2UFMwD9obNh3
9mcPqr8fjriGuHYV9SAU8Qn/fU+TEBafeTH2tGEAPG4F5lHYhz37Exk20aIffLgD
tlbb2gfoY7WXnYlzHTssqGZMJ4pjypcUyqB0jCSesN0LohRX/mr6iZ7EETA7YjLo
FndidK0HnNKxHIqEZYpwNXIsQCitcah/BS7oXZRK0g6YwSPdOKkCgKrBosbGlSXZ
3heeSlV02X9tBlJGouc7wLDnpZN9Sy6z8OBcHvYZuJKIQEfAwYap3NHd2pMY1+l/
DucvNztFTYaqdfxzm8AQrVWPelZqFJY/QWyaMhoenfEOzR6Hu/TXRB1KJgratZMg
noBr4ffUO45X/5Ou/s8awLUT5h+wi0/AZfK+gxKhc9qUMUp+jPaIDbB+7R+PX9fM
bexQwgbhaAKCdmwFa11MMzs/BePyLNZN36XpWc4OWVVbvBWP3CWG6a3fEHP31LuI
i9HIKVP7Sq/myFzYTEZ/2WfLijLjE+d9ItO5ESkqzXc0ILWBwnpfeB8XD9uK9XmE
8bmt8JdAlSXPDvJF4ZNiEINdineXXBsi2/yjMHQZMaqVUFf4C767Hf3j94DQjxW8
Rc3GPnSBcCyky398FG6GjTMIuO8SZNWeFYs9B0dR9s9wg2nwMhXNMbJeC3wWGI7Y
uoHFXk39bgnS47jmrAhofgmQt0e8EFNcCOePYslUtPgRgFfOi0FRZjR+VwgrKaVJ
zDZhTVZol4HevnqYSCbyByL1sYVZVKhQBN/kbsApJ1MXLXkknKCKaytIRXafk4vu
sL9hHh14jX6cmOEIX4vDLUGFSG9ooy9XNfJZyhxMDPbn8RZ3cM3pEKkX2rf3g8Vn
z++Zqz+BddXvyobXVNkW8bLTIN2+YGmH9yiXRY+/UDaP1hBwNlMzDaIp+FGKVDqI
J/lkO35Wsx6h85DfVHICdBTk7PhH2qCh0yF/2+PvsF39EkIq8i4oznceoZvlhIaK
1O4wRgHVuSFfOdYwBVWXCEOlVsjkbMedQlTqKMnnLdFto3dNcOMEC88E7iDG6CEj
g9SJwEA/+QPQjMUiRLoRWU4Gn7A9NfSy4J63lP0nV9B119heoDl2LReMcbarmLcZ
E0q/4IOcYDD6jC9n2FNy7AJjMXuCb7cLxa2+A//B6fTPOepZBF/+EEEvwivKGrSH
5JPiuvCX0i6det2n03GLqMsl6x0YuUij7mo3p/WB2mY+4vzGfKG+YZU2zdnFJYlQ
tvZOgf2DYIXnS8lOY8gCUxC/naQCpngbUZA62jGimtX4wDMlPnDE2haqk1oQCp85
zTeBMI+UzOJLq/DezCBnepdPAVj3m7eJhjSYrnPjvaPVwFHNV381mnR336V4lOdK
3HKoCNGYEqJbYUeyt+NgCQZ1+A1gbFwufnKSvaV5crv4LWrUpzP5djlWbS1NuS7E
yBF6HOp0H2aqjl0JZJdroCgi2gGFxk7KLdq2sQXzLC+725FjCafbR808u62toJx1
wRnwuSuDFH4W7YhO4ZKbmAimgltXNnRo5o1Tr6QmAaWGn9BnVAChZocupq73Iy1n
0qZYUvs5GCuiypT5m2oVtLoQepunhFHuTDnnJhxzalDo+gbMOw3OuEOjMbA+TLrF
ZXWuug2hnNzVXpOvFJ5b4d+cHRETEQV8J51Cs/Q1JF4NHVlX9cxZYtiFBPeJyNQ+
BnK/k7yh6MfjpJ8nT+ZGb3SeDSZ3mAD/Ts0CVef2eLZMN3hOvg8ZA4lixIla7PtL
+6dz12EvJJLagRGB704VmUQwirP8rIoGB6EIcxBEQp1urjy9Rx4jSFWulnXWYUQP
9JsTwx+fro/4IEBEAVHmqZVreGuyCKI6uQmB33yE4GhD1RvKr5UBRAhKoKO35KzU
TNDcylVoYTT3PSRdbG5kSee+0ZS1GEOeoVdgv77H/hjD5li0dpP4b4dvLziETXcE
H4Ye+6OKG8WP5Tqeg6stq12iSLy3LFJLqTJc1ZOE9GIBSHouLSw8zRueLV5uOvij
OzZfmNG08s/ZNJST17vSbkpBYdYlTFLyDzkH80kZGn77ED3MdgrVJBDCBTcPCPuf
s9iRKWYVlxZQT7WZmtV8PPm9Xrob8CBt7IkIHkJU2Sp+MGWi+kgwsD9KSz0zI6wS
gD1CmLSYSUPjCx+wRLsR6IrH4Q/mOwgXFjti+1odqBlBGovqhKrXMQcMoBIjEsDF
ctMCIju1BZMNZIezTWNLxXGLIfguMEzmw6+jkpr9Nl6KZJg+O+7q0+niVbquuNYh
qooEG3EiqoUTq4jadOMzt5lsr7aw6EQId3hDodc7p7O8IPmAvOgGp6SEUfZl6K6i
h0J2nZWdb2lWSxAP2mdH3EO18dxgvr20HKzIxYLkTC+eArRjDkVnzvbRdUG5AfgS
gfo7MLExzfIhCJTOjJBRksUdnrxX4SFTL+KCcaN808e+u/+myRkDRHaEfCULiV6a
oyzWwsNOy7of1tjTgLMc/l+H6/ujZF36uNbB4evA1liZaSpo0AGrOcGuoxwohr4t
zuaZAlkxpF4byFEujv5jlDyms3vvASoLSJe2jtsq1DY9NL63tP5x9IVz1VAqKK8i
tyy07C8y+io0EW6tc9HEzBND7ZKhEQF3Akdb/oIe2tmUFzNXUQ3nPw8yZnv+vSbd
stwbKHl/yibVzEkwoxLBCPbIK3DM0muq5cIWbi/PNZwVUijVKqo6ebFd0zB28PKu
Tj+mzDIKdzAMBJgo1n1wGIy8cKLmuv9j4SVaDbYr3W0Bbw0mAfLHsmm2tHPx3aqm
iyJXhKVpoBCzh4Jpy5XIORs9AN/fkxqXXPf+9ZopT73FXf1cSKsljo2JBKCqPmT3
Ngu+IV7C2fFpwHM9QMv5T0SHZ9hzz41vVZrky8N1/nA9LWGFaxOcwBkaK0/P+j99
OHHud2iErmj8AbDr+ubodFza5TX9qpgdP8DOeg6gpHP7HU7YfXoli+8TIoHAfR6y
WdscErGU1r10qx6xovkcn+6BHAUttOzLWXcfeSQmwyBNFX/aEwjHxuhXNgcF6W3x
0kTsn23JzlMuRHWkQpDKzPtDnM+y3KUoUtf+evv9AsFb+bZK0YPCSGNkA/xci7NF
DL3JuX2NdPrRRqMcq+iTbonQrN3LMvkCQ6X1Rt+siepp3A0ms6SJKbt2WbHkuRwZ
kFLZ9wu7eG1OkZigPPzUyVVahMwj4W4fy4iFdZYaXX/fbMdeCuD7AI+ouRSaYuMR
TiN7EWzI7ee1AdEd2d0dNsuH3aJMsqniPOT9PQkLwqN0ml5IgTW8I9vA8eKrhvCz
NHv7V03Huh/4w4k4JFwpbcWDoUmgY0XXOrFHkncjwM4VIl2M5J49h6mH86w/+/UP
KnFZemsiB0BxzHZ8/rPUwUPa5ikNs2STHp7OiublVcnWfKNPHAB2+8gWeCWdhXme
o5eAcbpI7k7h8zIy79fhBHA7PqKahFjNwmhED51BRBUuvXlQKjpQ6Iqy8vYGzyqn
X5eE8C1r+s+ZLT3Y5UdtkA8G4gNZKuLvNH8m4jhMNoBONjofukFbU8r+f89DKkbJ
BANRCgRBRH2gB79DYdIsymcUIvq7APoYIbtylsK1AbH8JfX4NyQyWEftE3DdANPb
i4BuGaOo4QnDRwBOBUOZ+hxR6IKaFjHHE3oAfgNaNo9py70mFmu75gyAKEqeoojf
6PIQgDjjY8/Bo2rMGQidVF9527vYk/SPH+3rS6mUUqmbHooiF94rYxUEjnrAjacx
tMjPMvdR3WuT3cGIF+3FRDwnIN9e7j+t1mKIjPy9wt81//UnRsDqBOkLn+FIIKcD
jgNyIK9jwaS0ebjdoL9yY1aRl0+xtmaEfCHMcFwnhqbpKZM1++IW9QWyTQ232yK7
tiwNXAfgg6IfrDZBYxzGiaG4O0K9CaYyKTHHTkgphf3POUPVvQl6+V9x9J9X1WRd
Yatqd18Eeu8mdqySDqWxcltk4YjCtXmny9Ybahur5O6kyMo1Ov9vNaIxFX+WTF4M
6C6PYf2/2eSx9xO6gtPTPVGkYb5nLO8UQJtq1Y8TBK8Ac7LAgTesJRe2TQmCoa7u
qg7Po6eKx8CXMYtwvzIxo3x6m5By94SU4X+eaZ1wsPMFYkDU0RTgg8YRo+pktZf0
MapaQk4L/cgBT2Rk35maczOC1bi2YkslsKFosGAZhaBrY1SC1utGyCVlCLzQULpa
cvQoD1qzGlmWb63nVi5bgzk0FR0hq19ht63BzSc/a6TsabgKXJ29gMx2kY9EYEC2
Z5hjzb7z4Xkvw8GFGpqG3lfrcQs2sue00kZVXHdj2Fkgdhe+3zSXUu9TjYTlUjoy
TwnChDZ+1m5+Ix0TP9HjGXC46T4UYuyxXQ1YrqXQOw6uVMjj18WQuS0ArUvb7YS/
g3HFTzAQ7SrxQV45xCe9JyzWTBH/PHwIbC7vnu6545shcFcNh7uSvRmqgHxlRF2d
eeJMqlKC58V4W4imYJPxt55BgWkfvoydvTskSZsdx8cdqeRBXzEucgDIh66Gb10y
x9E5IzKTMPUXeFHI1xqe2da2UNXJX6eN/zEev+g3jR5QvfNdWso6hEH0VUpykBPz
zYbvfhc5aYU4Hb4+tfHjWO0jdKcgjcnKztUIYe/kh1JqqvgQSFuaPOP1u9t0F5ks
EUEHk7bgZd/cotYydK0Blm+BRrwRUWvRSPU4+1fcFp82/SZRy05K2wLiCInCFjMG
Us2okvSiEMZ8RnAqBEeD9GDU7gki5/gN8NLiW2OEiB+TKNodCxmSrmp7+1Ovfmc6
lGoT6d+yQjcoWDfz4FRYdPG2e6nKukf7EIWm1Xj9iigDKdLTZxcz6n4WPYT2oxok
n1cbGf6a/gC7HO6kye92nLdm8IS57QiRa3q3eJ3REjmRljXSfYzUjguZowMTTXjC
ULGgQ6XfdQRdxwrqdJfpTC+h5oYsFtpEQbbOI36p0DRv8N1NXD4MjuLdHbb7FcVy
BSCn/ZGsssVf5lSelweikf01+Vkz0ewERsM89qytFIwIbLk8Ks3vMhv2VB4jC8V3
hTW+UvuRgTRehkHSEOspXK0DfSyy9qtQdZ+yz3GOXRlT7261VyV/AluDqRHOHfW8
qE3WD2s9HBsv7D0tp8W5oFoS8cFGDbqQNe7cETn7octEdAf3pFKQPu1QxId5hkod
FProp7CjyLlbNY1G7qJV03drKgGHi9ADaS9MF2FiKpytnt29g3iXXUBackD90O7N
5ANqKbakW0z4ldktZltT9z0CaMZnoBMLOuf3SwpMCZ/pfKtZDUKvWHkjma5GJKya
t87WqeuHIhhX7NWnpCa5tk5+wKrvwt5DfVy+MpgYF5ASSP/GLSERlywPVe+Djrjl
uYh2aWkdqH9yZqFOScrI7u7JWcCnqlDLCVDNcQ6Fxo/b1NhfpiLCX8yNpOUjkzff
PBRaxBG+FUlrK54AHvmE7lpoRQ0sgY8zFAqmqAWuirkkJB4m/3hLS+Vtk7LCTtA0
EUSuIMCkv4iu0bJRlj8+OfkNHKPh3dbdR+GQ2wvcqmjyvm2dusa9CM6U4HLaQTZb
FCL1BSpE2/IbL7PA9sLoFHGd3S6cpf7gFnR/GmwKCfJ/NyQjlgqy9a3xV6C+5sOx
dIxQpMBXe0mM6KlawyJUy8Auc2D54r1uqCTz41D/wRSRs5f/XINZsEY1uDpvyGw0
f0hxzGlNr4fitR45MgEHA0z+g2e/nzjVEFfpaZx7VpNVRwcneNq37h3LWAI4+exQ
jwrbxeMgXPLr5Y4teO++z7MjbNiddomhjeiJfqSXuOGIh31Jlx3oDXAQxxRA4KHe
yya9goqh/amS0OVjlIBWJ4ZVn/SQxp5TtHrpj8qeGlj90sAPyljIV+ABScKpSdiM
Xupz1Piys/fbLjyqeykVXFp5uiEy1w5s9F48OoJ8tj68TtkTOy1qO0VXwcYCE7nM
PEeMQzEAdphVZikvEGNazeTyipYIaLSX8NnijaVOARxRTVLMrMXWc6tiCDoIUWva
exMq/v7L0HSc8YU4M3hwA10tSuTLQEMD6Nr8RQRUVY+o/NM0mMtxGpKx/DuyFYsF
ZFFdJ9GxURI7Qn8Zw/OlAPOz7ll/5n3kFLeb7Ghw1S+iHO/5jDQUCLp/CKj0oiUb
wDBjUNXwxCrkP6AnjUXiZGlhtQXn3e3z39bUpXqE3AHHUDxwOw9xxannGujBqy80
BDvyhJgvJ60omfpQEf4enveolkXoJrQhXwTRcBX7yoHlKxBsQ8wK7XVvZRHaf/7n
CTuetc48R0q4Sy5hYpqxQR2pDd75kG+l8VJWgk9A8GfQ/2nUieCUowsubK0CySmI
jBY+mKsrUT9k0kxakzYV/cR0yHyrlfb3R9sHe6aKx1gy2gSQPsq+Q0QbqiUJLZVD
HYRi2uTWa591CnWC/hXtLgVwiIXplPd03dljoUdjkMhlQYNIgfKcz+P1aObLNZym
mb67+VAPhNF5W5Fq9YPqY2opWHUmpnArxwnaRfvd/W6Litkh6YjfWZICrBNrphY9
RBKKQrf5hOswKL9U4NwuxmDxHG6M++EqsmAYKAbw0GyVqRTuM1UQx6PuHmglF8ET
r9Wn1UI5dPF4FiwXYPFLbjbaXYK6Q2TgJYVV9zIsXtoANufBpUroXqDEm/BI+w3t
X4uI/VFvLTj26PftoFggMTkJOe8K2b+R2XH67C+aN4ECEiHGPwdR4h8mkKWg/mhX
3PBQsf9O06rguCrnCZGAZ4YycTotPMUHoEbU61ujUL7b3yPh6htu8flgyD9Kmfeg
rLMsxmgDdjqkifuTlkmPj2P4oz1M8r6fDX4d2BX4RKZJYJJe9CO0EbqD5292oIyv
O+RqmWrJvrhXESteP4i6OFTp2Ytk5RnY2FEBBfq6PxTQ95EZ+INcXS64GB9SEhF2
L0iXmWxvEnapANOwTavRWtNLPl5OOJfqSRLZwer2CDB9yoq60WCkeHdGwf1T41OH
7OtuAK+9B3w4np2cMKIE79pUl3xYJ11imIblbpJdSQOT3VphNGlWziyWBH6dy2VQ
WcXMBKSSJ7lSs4slcPXxSUe8rEaW4dm7+sWifGaTETJbUs+z2yI2U9ySiwphnL4h
/tJNlsaZRrEVcP8AdNiJ/f0jYMDhnPb0pYE4qNzGwPG9aMbZ4yB35XcwmqSW3Fx1
CgZQeXc397SxZHIsXbY6VjBD4dJFrjT0V3TInQ66aDHN6KQi4PrdgaHKs4ea7DKv
mk6hy9AHQYfalD1x9W3aa/TnLnnwIoeLXubEvolI2MYVxDbJF4eD3ZupVRc1aHkz
l/UzMUDzfc0m5LMjNbq70wJnG/xiVMqgKfbf9nzDVrDFlTsJiF28RoQHLDsWB0WF
jhJFZ9WMAGRb5BxQrSY1ZcNBdPYeZEfuPxGIvEEUkZej/JrtJCSacdb2ryRBnPT6
hG1s6a5fjLhb0lFx9W25lcFt6SRIjnq+tP+5AhSzw4wVNwS9Oj2b1AcA9E9bFGsZ
OW+dRIzfauWzU9qNsVOw1Y6WN7px54ZXXngjYP5bZlkTrlteHOzeIooTo0rU/JBK
qhxodWT25vzTo6tjo4g+epz7RI6nfRNNheWwwnnkJuBthV87Pwr031feudtF4DNu
51uKvD/K/YWo20/s9qPVO4K00rAO7uNX63jeVlukSVOxGuusKIQ/FyK8FrjkePaV
V5yWAQGiY/Gm533KORJIxx0cYnTqGIqhtmpdDJfKWHDu3OjMoZV1/J78PewM24Z1
XrJAf3aN0jnCpAolwUQnTok/5qe2QRwvOwsQHWPL8N0E15RrkxZlUIm1Be+R6VlB
bIhZhNzARkHjbktRuT9KvlMdTTFWWhoMgtjGoIEqVE5RN9mtiaRb4TFFUmJYT4y0
keXCdjDE7r9b7q69479/kWm3eVBAOemrm1ZCuFEKeKlEqYS+hrym7jJvHIB/m5C0
1MeFNPqWmfA72pwFUPwJo5nK17mgyq73X02vHed7Qo3gVcUurJVWNzUa4shJRL/Y
ZB+4wVuU4ZsfzIOtaohHQkgPRNtNikFlDUjREpxJLGa2fM05rVkjd06CcI5/9M/o
ta9GkkJXEyUmDZTHG9INYVFuDN4N8xEJMHeA/DrwSPIQQ+obyuCCQR5anQGyxxRM
H6qZsjP/03BFRboiRO/teTmmIZVREiCXOnTNSg10H8cyhzVh/W2+87YXQvZ9jXNH
yxOVe8Hh74vlpc8yF5HAETAZcDBBaxI+dfVlA1pPaHLr+2LuOINtTHpq07erCzXZ
miP3hLSAZD9/rE75pZf2fwA3u4JFzSOonw1vxx8o3Ci1LvxJN5avSPj/KB6W7TX5
xBZZjjkpxSfzKhOoJ9V4aiM5xlGXsQeEDRkTgDuSTjFdnBMuZ/QX/CwDqW2awXEq
itfuFvTNfQOYcfgYXZ8Ouu0mbA9WzzYqLsy9dYtuos0lzhm1/j5IoGW9iV45OYW4
er8vHH0RNszqDFrK5zpz2Uk2SFNEL6rSnQpk1PcR5e+SI58k5npBDnv0PHupr2IU
ttUA2hcpAqYUItix8BmN2biYhVL+TEXJ97lf8bALWBuuM+aF8YPzlWQtq6Wm9cpr
O1K7PJ2lJefHsIm2/a5mfDgAKBsJs5RSf3ZwiEJVSYIe2NGaR3yt3K+eeHtdRgK4
mF8/z0jenkgDoJGjv1IHTLkkvoGqz/itRy8mSzvOWgqljMMhYug2BItk1nWYYrUN
vxqJ2Kx70LnVmkY5LzinYnAj8vW3MFTkutDodTLJlCBHVh0mUV9197FjZ4tfj5Rm
AAPzNoUdQXnRS0o6ruk6AEAumHenahFgF/ohxJ2/XJolO3cSlLT5i6AaMaFJRVVg
elsp0f88UZq9gcAg0pkEHeoRfV9reReEGAqTUWZGJOHOAkzeg1hheZ6U4yzu3TOA
ZjDecoBCN0sHWmvocAAGz3t1lgybY8f9CCmBJk3yCBqPjI0qoi9jBSsId3QI9AT/
GTXe98HOQWCdB84yA/xFG7Ypjyl9WwhD1WmmX43fbTrC0Z0A622TekStrSHYC1tP
azE5e+cfOGfH6UcvZiyIT5hJMivWRaLUcupZlAbLcwTKSZkYOEhMhnPq7D5D/3GB
q4YeudE2MhHYlZc8UFbziQ+maEh86SM1FEgY9flzYb/yqIJDynF2e1jt72KWesRZ
X9XvZ7WVnwDyc5jMM0lrHm+eV/RbI6XPg+se/O7gr5P0doXfbbIp5JWq7vWWJ3Dz
MJrVrsnO/3PtP53IEfbE2jLBTu8DKCa4p0n31gSAph95f4Nc54z1Cvf2EAfoZil1
XjJ9AQSgCg2jqvw262K8qmQiFeRKzwc+K8tZsMg8c8tuaLxMm8dK4y5+P4Qu494v
QObqkdhtnl36lWJAjFrG3z4PwiZNz+ATVAT5puRUKibmIfuUDpGoFq+RVRGwe51b
u/7CpOLOPTTsdYNnvRQtHooGtcAZhb6PKSXTDQMRkgghpEk43g4VUqRzBnbxjwsF
ku3lo5/AB/MXiLfnDetof/dSdEGcxE3UYjcDvKF7EK+0kHI/hlULZ7l1TY6uw2Wj
B8u88B3U/i8u12VhZfCedmcJS9l/w5YvhCgiZhYBoZ9jPHb/Am90O5j4zphqR8aT
zP+rR4UbhDaXuHn8w1RY9SVd4UpgSgtOvAXPlNJJBBNAxgo3FQp/Vu0sq8t74mC8
IYLn0nIdQuqSW4T8RoBg184M2EHq3OSigAZTFt0p7eLk88fKOkjuvSQjvk6v9NNj
udiYJPdm3YImFoxxT4X/mqH61BojsjfSwY5DJ+qF13PEuqzONvnI1Qvb1oZuMNGR
7KeB5Jr9PeUGKPpYuEjpoWyzQK54UixMuG0lg4yuwg+SqVuSDh3XPvbiNRvHRKYj
9SxoYCC2TklGo0pzXWkF+mMBqYmJDiz/1Y7Fj3JpmKSHFtrC89J7Tn2+6ckFMqMl
pPfjjo0v1ajUOaqnLuaRmmzrcFrDbRMtRVDrvNXkGH0+GAHuHm1CB6R68+2RHkpE
zEIpn8GMNcdFB0nbpXa1GdNmoD4hMUc8SmoJPdxFPj+4ipEZHiKBFm28rqI0PEw1
ZL2M6143pDoCA8Xug+3Ld+OcK9acpphFQRGh3X3vAJo2qUwEP2dlCPBTlc2GLnWC
dd21GCL39UGjsCdKArtMKhzoJgq9CllXK5Q+K6XVIxeL7+/+rmkjtT3E4ffYdcNb
2qFuhCLTFh/BNWZMqUkSQ2ci1rLBwieHoUdx/TvQVSDY1mYGjHy3qw82f/1cJKVU
ei4qT5SewxPUHzp0PwtzrDQ3MVs8ErT959nfIS012s2f/1j5CpvsP7dnbjAlODC6
pmehr3rIuBTE0tjR+wpTRBHaE8A7i8YwC0JsULHd7DrPpuLK4H5vXradGYtQD8rr
S7N8ZW3pyJNORGN1XkGN66msrThDiyz3VBNXGjWj9dBuIfzNWQnvgZtjzjzT8xti
+h3gmzlpcj0jv+cI3NsePkicZB5H+Qn4fVVyg4b7Y4lHlmiGndv5mDJglTDlSRRj
RKQGz4OSzM7GFZM1e5/dugQGHfn4qmdr1kxCzCqFIRjAesryLYGjrXPWq+7Bhil2
mxP5LEbY0vYSOQqj+pYScGbT2LPLqHMlYpyOj/k7Rlg7We9nrdkRyhUDkCHnUxAc
ALXPQkxvQ69mT0I+HLDUnKQ99UIIIRhk+TwJeKDBCi1fTAjhJL1k2lpI4vUdg5f6
4/DyS2OzwI1Dtt09X2ziZa5WaWidxW305rPbeRcasso/dvja77LAxGFsYQooZzCZ
MSyILBI+QUGUij2ZO45S2LuPyJvTLrGuQe30rncMiVl2znx+eNmClGI28YFrUB6M
XgM7z21jMEfz+vISqOI83NxrGx71AUAKMp4k2bnE5lAzOWeou/P7AloekMDcVRWx
3seWJxqRbg2KgHycfUF/Fiq3IrWUPQhb1YQYXakxOMOyqMF4ZeWSd/h1jWgJ/1++
UxaFnwKO3NNKBeVI5Y6sP7vx3nzEmjXrDrsSzj34Ppj+biGE9j6MQ5Rwvc8Ytse2
muB47MgnyNLNI/5/vaIwdaDiFXoKovfB/9PbCemSFRX97WkE1owNTprNPCZSat6b
D31ADv12eOXyZ9tfL4MR3dITCk1PixEFLsAn2QZzhmK1bOS2SNqZTnb80/jgWY/v
UDK9jHcYYPzSJC70RRAL8ipozeWLhUuNWbp0YOHqncAOH1slsx6bvcWtzjjeL1kU
GQZuoMtc5mmnKPRsicDKsBsSGMuwh0tFmJgP3KkgmVjf/EDZVwGgQJ6KVT1hqBPK
ArWvvs26Vimapd6XOhTjLmyVZoX+oSefXJzXbVfrbbltcM5L9XQIt5T7XeSRFl9i
qtYel1O2gXTqp9BAtBDmIReoq6KgIP5IkDq5qw2QAor3obWKghcSETfoMp8K7eqL
iQ9gBzyoQpojR4GFGal0wkPs1IJbuskAL70wYJ60VnbakR+Z9uvVNyPu9PJYtYso
SbM8+3ZED7hx90lDeStN1NCVhkGtbR49rDGEqT5u6WAYF3my//KSj4sAclMiFYE6
58ODpuPS61TV8NwBnsMywpcZtvS5NeyzsNuBGBkftYXfEIz95Uorwxx+86DcSBi+
Uh8H+/bRlTqiNRSyGr9sXfy2obeVmO3aznsjH3+S91uBZPsi5Vy07BDSq5r1Qh0a
rGClu6dXYSsyZ0R4mB4KdL04KNAm+0cKxa/9vqCnsYTm0pQU5tdmmTYzMs57vxWJ
5IFGb1WgbcxFO2If1r89up616XMOqlw9gdh5zY8sK5AN77bYF335AtOkUKb7GT+J
+/DkuvTHrmtf+u5dnu8B5RfXTjdA4C/cWJdMZrM/POip5dFKKBqjr/2bxEVsBH1s
o6z+zqIPxdsYXrnSxLgDxJI/HRxicePhxl3Pi0wDNUge8QHJWKY6w9ntqowNTn7S
v+rDNAmJzasYLk9ZF/clRJP/59Cshzzg5WDCCEwooieFoa0Ogp6mIHTICvielTv0
NOQKxv0HKwjwTOONWzVBPMbeFNUcFvDPZ+6v7J6iRYrTwPrjZ44DZTxsULu7epxD
Kp28ogCpyk+8LXp47tlucgbdFaxFOUS06bMtMVjikEtPLtrv+xEq9zPryqiyUnrG
sm5O2JxZd366rjCcr1theY2esb0apw+yrFyG2obImuMYovmNhfJ9iJjk0N3CmsK0
OyWSHt9UCGQ7j1+RT3O+ypCt/tVZoHsLc2bFTh6fmOdgRUTZwYVkQD59sXVVZ34r
WMbrrrHQfH8wibP8dzWsNcjQjsDI+lOuCMBjkcComTYsAclyE7vUsnXwsTcR3jRH
Ti2dKiyoIEwkD7c0TRielLQnwiSAH0e0FiUE6EfwsBhBSx26NJ28Z/zK+4JX3vP1
tYgR2KIzu/b5MEr5Ux/yjnBdaByottEzvi/gn9V5Psgzfz8rymaQ/in7xMGd+tav
A+SNJlj0oFf7c5Sr39MhI95WR9VzNExCovqKFUXhAmPWxXxEDqg/0jokE8fq/6tJ
HoY7XHgKf5gBVCoHDmRHv+dtOn5bFn/Xt2oqa+/BHiF4lxTU1gcqZAmWG9ffX88G
bad7bEyvTdVeUX9fJHo3U8BN8L3xWQPX/Mb+gkMPCAy8kjBG4RlaApILQZH/SOTk
7HZpuV00PZl7wY7Rw9c+S+z+DIN7i+b/JEWFPm9GzJffA5KeY8a76Orju/5ITFsS
rnokhwkike9muFV1EPR8IOfrn6sguKg9hEuD6lwPeyPCQiK5iuiaR5kHe7qZpqPV
jsxIB+IITXgRoqpseJMf2m7kZNnYn6xbK/S8qrFLajNbfH0aDput7bXVsOw1r/HP
6Yl1aYAtD6i20vbLd3VRQsvk0FdbvtTEkV/2okS3D8k3ly3CNNEQ6F4+3xwMgEXh
awbs96d8YLvyiug67d3FMuuO6LmpaeoC0feYPMclbPN0D8PZ7uP9Vh8OoH9ED3Yx
SeqZ4INmMJVaPaaxa6Qwb5e3xq9szipfZIzILw5BEFeO6/D8HTr7FTJ8wTZ4Ezjv
BSf6OURnQU8O2zVwxB/BdSGObtsjoLA+JE9lmJKrw+bKnroxo24zURWybo7Ay5G0
jac09p6OVG3iIEXmIEYICXww+iW+kvTAxZDOd03OSvtj4dfsy80kUgT2ZOFEfsjA
SsYiry3dALfjT1B7dxo/8Ii4bq+TYRWCEfWkzP+ICRhzYC870cIk7JszH2+i+MMP
LprxxZgFhpojhguQGZjwUaFE9xmhDAS5JcEjU02OP4gzE+E1O1XcTavMC7YZyikK
GKHinVlasDmGMGFdobg6FJrDufC6Z32nolLApd8iyvkkcuelmnIe1cTVuLeceS5G
B1rJD8yOlPiJ9M9X2TXqjd8GMm73GflMq2XaC4yVwdVBC0ZuKFFclA69kpc3JZ3j
SynFzr4UmimCdxAB1JBl4aQYJgQ8AnvGurtrwQiR9Or7sdHr7fQ8nNqCt73GG4aJ
Ppe+KVyBrWsNyEx/cBQO9Ys2ixVsbaTPy2wmzuKk579SfHRFT5+jPcBR16oSt0cL
PGSh5HJESa6kLpnbMCFf8ZGLLJKXW5BCJfIupnE6kfYJmld6HyL0uMPNBxttygcA
e+VFm8kZXApjFi9Ku6bungEipsF5OsNoPyTekW8UXlHjzdrbWj9S9idVWtOqs3T6
/0Jqb/Y4+OIOcFAi+l+4lyFSFGoPrrVZ1AC9oZzWUKZ0Z8mKQE694uBHpGOWfbcq
8yDqD9rz7CQL9Ni8y/UUlO+7g59VvDVR5npvwSrAYQBsAYxm9/MgEgg0w1VZfl97
HXcRntlEQ6r/HkyimIYTzw7SAvxlmgvvsHxTrEBf6WA1g/GGbRA1pAqmffsz+3PN
vbaaLA2Wv68anxr47cVp+QPMuQhsaUcofL1IGX4RyA/N/s1Hx7JCmNzxe00sHx2g
KOE1IfnjC0Wv01zN8INiUoqMhPJkbqxQfX1hGFe/oaXQpQZGEtVsa5QA440Gq6dD
y+pwHwwtjQcRnFrv9z4xV7vdox1VXJwFafvg1GYVdzQ/xLCwwjtjLI4z/uZTRh13
cYscPbAmfbGiEDoy60O6+iE0x44Fe0st8tltylLwHK/nuws1Y2vFhmJcKnZH3YLE
9Tf0DsGJ3oxXy/XWSfCQpKuWeoDPba7s6P7SHh0mFvOlFSizCezMNQs0Cl0laY3F
PfkOz6HvNb0C4f4pD3ApNExuUpSYGjKoi9/2fy8InbOAsx2BwuEVX5Ut4CVAs8FY
BcRNwOpbWfppVUHrlyrCDJwU/xg97DWlpLPUKeY1Xw8T07O/ViEdf8FY5IvkHWH6
2teOLUQ60TgYjXYMhjSXT6rVF1R7V7T+gr87Pa+y3TalsbGLfPhVyqksM/bTJKav
PQ90bqo8Lz7+08Q8so69+ZfaYrc9pvYE1T8IB/kuhAtRSRg9oUvcclyonPOKrVc8
TVI/BRnVv9tJgTexDDgTrn2jRDX+xkXxMaXMZxyFqg+GwrhQDFlJbH1fkIVK7Xeh
Gj/eZr4aJQxJNvdXGuKBXYNxotSAstYOq3cnvoXjkFrLQOE3KVpjPEo/XhqVbBUl
/2Ac52wM8/ZTTfT6eOagvJffy5bESKObRk4YutPmXRaHQsM8klnx0Br//5nx9dtf
sSmPy4zvYQFmDW3E2XK6PamGaV9NRK2GTF7R3TOC9LORkHRzqUdO7q4+kQj/LVeT
u9g6ZF1XdXKqcj8HK7fWNcLUxcFyUxzq6+DpMjiGQPlmAqF1k8KllFEGaNCFmgXL
+5IyqKn6HWaazNCAg+OLWlCBkjo7CmbSh1sNz+P7L8PUGTNYjJ+EMScf1Vp1WT2R
yVyuHAi3sR0KBM31c10UYwFClx1cPydaSNOP4KYAzyd01ztCAsHxO0gSycbmlpM9
5wqISxQggz+pjENYgTqgwCrIyO4VUNauVBaD2oXnwdlD0KsO9BQxans826IAHLaK
Ect/xmFfXhvwJeu88UTiTmeYCUpqxaLX/ThYuun0oLSF2brARKpL5T19TlyLVt1O
v3DFJ6tQyDOWJRePXLRKO+E+VfcMQ8yJ7k3xzFboQdC5IqhGl+2kdJzK2eme+Gtw
BIqmYhp/cQfoCRyS+/5kSGaMi7lmtAGMYA3pbaNSl5Hkcw/IXTqaarriKkfBhzL/
ogq2xxWxc0Yru4RmWWdfVRJc30fMYlkVbmtwfE42BQa2EnDaYFXVOD6/5V0/QkLM
/vL7V2fL/j3ILUW7493wiD27GkjQ/GHoHRn1v0Bfev6nLuy2zFWQzuo7cxL1d5xP
0xiTRgCmeogAqUCZ4CK4CVPJt/jkRn2FsIjLXTfHtjLhkpGCGwQQcjzWXTWM/Gw1
ZkTVbNJNeP16UUeNfhiDAIJL4B2KzOZN5RkXlmsOMC6zqMmINax5PenWFEc23JZm
VS6tf+CO9ru/WclYPFtZS4AvAeAtrkkKkpTp9bH9gnkCIXPdt8LSGjUKbEMgm4WC
T1VzNx/vYT1IjgEY+AWuKpqHjGjt4pfUmR1Ks+w+pPZ3Ob1BNQhf4hh28xfAevR2
ZdJlYFA0s1nX7ws/Nb9VQ7Jy4BPkVtJQ18r+jCEpU/UGegpESvAdjDVhZft+zl+C
1WeFhexJVDn4JFR1GMEcdK6u6BzHwAdP3topC8sbGxe8X0IjRI0m+kGpCQqz4ohH
1f/scnIG8/Fb52fjgYeEKDuiSUuH/qGwfpYgxOj1EseLaGeq98t0v6TfLfT62d6h
kyzsxxfhY48BbOf5KjGb7gGbnA91qVO4PUjLkJquS39ApfBeSrf7uefneS4kYAxt
VssJ5DZ5HsBeDiRGYwD961Ki+egmhtUWpGEMFlCKusWzIjWCJxntAszlOadl/8wL
+9nJU0TiHwme6gRIWtBkCvwRnR19h7YVmFhS2M8opY2WrG1us2NydxDsc5SreTul
G4xtX/REnyDxWocbOXF8g+4OgeTnkBmqSLbSdPr7KZ6DzTOEDQMPaJM4exkVLFOD
vihzgF5xtlZouiqmlq38Aa9UpyddtYXkFEAJbtKiT/JmZ2tYpUnfM4BhL7pa56+r
QEYHdMsY1Va+Frdutp1ZXi4FqqFi9vqOMN7aGgpZnzCZF/lm3ZCll78abBPRWnxa
83brlZLsKYB6PsLrM3Mcgmn6F6rJiqT/FG7tjEr/qum1CfCce5CuypBWllw54qy6
8kxh/LryQX/vB/yKaZNa1CWrAIeTvJxU2RZuWfXLCYFPUXpjck5aOM0wg0RF27XK
jZiIbv24MfQHYeHSqgv4lnUMIXREFX8CvuUPMYud0dVvOXzyF4VgdCUi6NYw0ldU
AzfHUpCq8y0VnAAwfCvZBQnbcfm3aKNaYyS3xwjKV/SmwUYNtiK7YIqfRlibUeTM
Lgekbaa9GNz1YeuygL+HuU9WMWfubCHI2xdu2/45kfSCs/2jMo6QtlGTPF1xOyUR
dQsAZ2nKU5VY7PJuFu7rgBpjgEuuEs5OvCNl+O6JY5SZ04J9K9yMIoQegiN5dO8B
RRcJZUvM2YejGPR1VU58gNMqKZ1UI+QNg8PMRcsOrCBvn0O4q2MOobJjeNoZl7kp
VgvZuYErg1yznCN27DQU6VP6pbeE7g3czY+6nU0MBDSCVnVjFR2K67Byz7NLrT1o
8HeXjSFtepcIKN27vMMFyuS4O12dbYgMX0Wt5goGUKYZ4/7UNp+f7P0EkhqRdNHk
iz0gSu9y3+CtwxuhjZmpgUgUeYEDvVDQ7AL2LuTbSz4aXA6pi0gN8AuMP4220ymw
0qwwhj8Sr9Rus61l53Ukb6hkCdkvHo21hD6qY9D+vCGBIgB1/7txTezJhcygGDio
6idJXCn/ow4quYAT6IBUJ0e52fP5ffVvpJpqudRb+qBxn2DppLeR3U2Hl6GBKh8g
B7IuUp+pOAdoAY6UIgEAy895+dAji5WwW0B5MrR17poQQB+QC11ii5YcTBdPMdWU
5/y1NlZ6y/4JZG7gL7Iga3Beao+/u8sQBmMyQC+Q5ruzpm5uBpMwA4e0bM1a8qZ0
Hhcbdp4Q8F4IDn+Cqple4KBVYvaMIB6pwB9TZdP7OK8dGmoJnrhiHP+B69lNu5ex
CaaoUrYUtROAw6H2FoUD7a6N9XuwydmjTO/WssTRR+NKohtyeBUXAKejoxBXIV/g
hC0GEhLU+Ylx4MUD0NB9dnbT+tP05FiKnclMMTizt+OiEkL+TkNZ+W1zE/icimo5
TCoDwTR/XszeMKFd9qvFHWt0Oolwr/dDvZh1WvLCr5uT6Q85bCKrGXpDGyf38CXa
32lJ3GbeaFOSTz+lkMpm1kZz8iBewwqHqaryv7a22o1TQ32DI9UxF0pPkG0KVQWH
RaoigG4pl72qL6yc/vez/9MwzMT723kzrJNNfjAasYJkIK62oTJlZe3BgOWOYHW2
r4HX70TvURbZjQ1XREHnZiBhjHGvm/QJBXZnopjuzPL+6jWZEeuZRJNRwXESj73L
uum3zz52iTnfPP213Mxfn9IqIzbpyOP3Hox2Offx4Zz/mOs/UFf2XnrRDfjtzPP8
Eu2e9o07w7rfE91O4p8yl6yUzEnpkcTdIr2TVXIirpA+tJYMDL4Btdm2IUBojZrY
CUMQzdw8snpkuvDzYbsD0Y2qwbzTiQJs/YoOMx5Nq0f7L7BROKJ7xE3GPMInUakx
9pLV5yIvifxebFFFZbFOgTPS8JcGx6wrnRQQxbf+PTh7x8FgkMRenJKQt8y3tBPw
FZsUQmikCA6QhTpf95F7YrZMk7lHd0/bftK6NEHcWRjCXQbbaRLIH1QRaL0GSy68
aRpemsKzOX4HudWS+2usQg03YvPwa3Wx4Z12apAHaM4HhKxaYldwVARO5eamwabG
xxXxvDJ7Sj15ov78EOQ6WLd4K2fJVzWcz0pf4TNbuAOfg1r3CltgpuYXU7HtNpUc
ruvSuM7j49bowCt2tJh7SGL985ukPR167YGrdwWhfUftUoracgxqORImLaO8niMi
I+O9ofS/9DcP/1JHP8B+pNpms1R0X0lV7360Xs0/XlruB2+iMDQNPVFQB+7/avBT
JPcsgKjsHoSF5gHE1kX8qtwfkb+L6nDXVlqG6M6sc4dzWAqmcQgzv+ZBMBmAMLCH
IZ4goraKs4UDHblqBg9UsV1Cfw1cnM427Z3CX+NEIYukcRqVYOvXEACl/bjucErH
90hdUCt1wh4hBIBDLslAQVa+QJJop6exYdKpITELke7iO2SiqV9esTL59vxdz3GC
ACA/PBka0ROAeFl29iWTNT57uubmbcHFDjG/FrsExhqyRAFJahaa8n6vFrbfZEOm
Z3ATNpkSbKH53NUzcSIC8gG6yvcS+ZfHtDtn+aMT3bXT6nk+Q5q6IrVhofYtkR10
mXt9Hpy9AOQM34JFxaG5UmPF1xDhowLPpwXVmyWp3PVcImmVO0ZgWSOa7DTrQj5v
O+O5A/nQGzHTFoNiawg9nscXi7dUP5J/Js6jpUQaH9ii+cx6w0GAmmJn3S0+QJOn
gUYnv/hEYCqvR1AEhURQUxNJ+wmKtQ5BDfj3KVmZrw0zxLgOsyEtx36pUxiJyD0P
q5ZrAr7/PLXbq7GsvcDhkFs1QJ8GvCnFFksGemEt930IRUhCI1Rqa5LaBMBU1Xrx
9amCE1ohA+Ye3E7woRK+cL01g6WfIBvlxXTRvzkEbTjOJM9d51OWs06r6MmFosfM
/jbb5N6PRMceBpT584oSxWuTpOd+nxp7Z2TOEYFxqucoitBs4r++teYm9fD/fEmr
5OyaJQ8vF93b2ZgUEIRbp6WgJ00dJMbw6+BKro0r5CMgwCcdV6mwXIGO0nQL3eiA
fAfTcEJX0305m0N2ZvJyOmP2v6VRfVaPLdt+5BQFpC/iLy2AXVzNAKfFUNCOjjPk
ICmHPmijaOqdjUviSLTYabn2lwIFUiydADKJZQNyX3S+qYAJCtblrLjuCrDCBtG7
lmocykfkh0slG+6R/LTPTDE6eIFH6jZ0pHBby0x7wwr+4kpC5Z4VUyDnjXvCMpPq
rTvI/thj1zW64qWv+hPlr3G9saAyYhgm0uD5RAO45H5ZBNUaUItVaxi54agz+boQ
TP7l2Gn/6V+Nagc6HGg+FRT7jtqSZm87kzKkfeGmVkYPzQFuuN9H1/dCqmdm1ya3
RXF4DEFxHyHQ8qgzcDXW8oRJ06CSta6TLmKbR+w1E0HmhInEUuiXJ8IHANwrKbH4
kOlQ6U3pyf4l/AFYwU/6qWmBdvMhoKYPwbyf8zHJC/BYkPRXPjBq7pceckwlUhyb
MUncy+k/TBBlpTuRVW0BSj/KXL9wG/chgxX+aezQEjYSSm3LtBg+5R8YVT4Q9mOg
IO3J7KgHEOopzgozdzXG2BM+6C8o7dFieF/cui3PsHkExu03H3IJhJf+6mYU2Wx/
MYLPtfvIuXooLkQRMnDaIcyqrHHQTEtZv+O4aipDYmB8bvIQAWoSUZIA3HOTRto3
DDP9D5AEgd4wko+E/k71U4Da5rRcp+ImoW4PkWTvMbmzYwwQdO2kVdLPp4/i8VS6
bStocOHeUoj/QUchBkPIgxucUcB2Sojtll6sV2eE4BoKxNCdn8trVT2ppD+o0KrP
PE3FBum5fBycUtgk8/hMT2NeFmYekcagCvLO1NPXv1zBGs9k5YOWCugW0NHaPcGq
EYjUs42maWojhvnms4zOWrpxMsGfUFrY3IJcaQXa+q2mJZq6i1ZwpSm7RxHwoO0z
/an9VUaiikQAOf2OBrqZ/lHXyDhaADWnRruRM4Kr1lYfo9hl0emOvplz6L3Q18Up
AFmOidkg5h8/GkSnA5fl5KKOuYJuP2m/YS0JtbMkyy+xZDPmxDpelmHul24tnG4n
+YRC2rVYdZWrDqcsSkonwaZRlSyfVZNfdFxUNr06iLD9z3VKAmAhogCYkxrGaePX
+G0HsJp4WwGTMAbcXW6eaFpvYW+zgB6yaoJ/7tPeHZ7x1Bv74GaOBVNdAkOiFzSb
f5CZykxAfPWoyOfpAbk5VKIaJUUjihtVvGMu+XUeLI2FnMJIvRDmnXSAO0ShlqeS
jXe2dNN4HI7rKcJmVjT284easjLc/tCY7D3rmslpCRiVXTrXiyXKGeW2gBO4ymon
BXjFApgR9ZGSAVffl/qoE5d+CWPURwbKNMzCv1ohxnutMiUKJhP6WOyXij1+QN4P
n7645+Sm0qk9NJ2X99zhgj4nCK0uAL40SEMZczPjyzwNkIzA10VoNDiABaLq4IaX
7eFARwXcC6UAa2QBkOSysrEsQfbBgKyFxowcAbZVYdKyhY6xR/O1HWN0kzWV8mGb
mKl+wYzIYxxYTYe8c2Fq2zZ5pQZ15lKxT7CfqciJkmAuPOl9hunef7TAaxdegZy+
61wdZCTi0RLcegIQ2FzBn9pDGVFrvN0AafDF6iJ+x7siIzWLgfkb1MOQotK+boe1
MIMpFicH/FMUi+y/9hHzKSH9yY4JisTjikZDz3OH12x3nix/G9uXV0tQWDP+iL3O
dw11tNq6MDTLhtDmNQaSe5mD14P3uPrtmE2bugRfUGpCimTh3fl0TTx1uq+d0UOa
dIquY+myjG9diUKE6WPdoaK4U6kxlQvde27+Hcu0r28KB/m+F7WMBmGrMXrNY95S
GsYHsQyZXbwp1Vqao4TzyU4+XedX/32uBAl3McAlQ5B8nKfmVkpm1y37EvGFkPRS
BXchDB7vK/9nzqeLvoDzIfnJvF8wiqjX8L3h19CHK395YY5Af7VZ3XsDPNIvnWuq
RRKFik4OK9wDHZN2hXrtMxMYqTGuyKL/QC0x5nuEaDWrslv2cn/EdXv6VT5x9Q1X
Jf4IXGUw5AhDKJd9gZi5jFJQAVvGi30068BFwVPB4bk0FDLMdDYn+DArguxmsw91
ia/0kYCSX0UitYh0t4EFQ3/MBSn7gP98r35V2LxCVA2/QzD7eJrZspw1AZk7JYrO
tGYINUcMkyH6Au3Cm6CaJmf+vCjTro8KW7C3TYtOMJBM4mBER6+lErV/RNEccT/q
oXJ/QCQxbQPauvTmndsTDZM0JIDA3igYwlFlIaWff29ihJv4A4S+PfNJVUh4ib5D
fdDCExiy6vho4iglzrxpgaZ22R+X8onOLTFNdDPbEfZd0i9O4ikt6ILMX7RdtUQ2
TkvNKQapypslK+7MUbygYEw47IJ/WBZeolFwiUzUHOMuqWtkuCznGidop1ngCcu0
okqBc8/6/dUWVFJEy14FsPRh0Wsevs9ijmTqMWF9sNDTnbjndFYkhoHuMzXrZ+Ol
kz0H0hBqXbMxxWvpPnT9v2gO7pdn2VwVMxiVb8tmKHdEphy470MQKu2kJL90X671
Px0ftuEBahPpkA+bUJIvHN3EKbAbsbxADUnoQ2SC6wolXCwmaTMf42AgV+avy4/V
pGsjNaVYXa5STjSqzPTCaGmM8XGABORADOHEZjbnazA6Ehpcsob1oCibi20BxaZI
LRkR7DCmkAecVtWw2jII8H8slDlBQG9aSZcDz9j+f6CnO2qg/26iLrjQXyNBBvo/
PHT7VSN153Lsm8MD7tKxm4WKG2fQ6b217b9mGK/d1WiBbh2z/CugQqLkSZJdMYc3
6UTQwG6M9sBf1BL4ZFOw87bJp0ZhQQca4BSgnekh2mpjplhJ5O4YUIs+CAbES/wA
emGBTLRNTXmpFVelz6XGbKUlhD+kFYupEHzZUB0vdwgLgX9J6ImwCDrU/Q9zNTZw
OJFi/M4yDxEKxKrUgXSdeTSEr/9TMei4Ta4U7Xxb77TpJF4LTaIXPD3BQPdC8n3y
sposnkMQiSIuutbpML2e04+0V6v1Ts5g60UlOq9dg+icNU3dLXSqYP2v5PrP63wL
c2nHabtawXUJctgAduscLvT9KcY9XWuvSO80wIhXwtWUreArNsaKjNe30Yw5Me3a
eeywJZFW9gMAz8kCMoOoLnGHyFtLHQ5ccBrczFkofhnxywFGy2GyyvoksJOwhQlr
3NGon98gsSAILbgGkHwhdJgSUTzpAO1LAib7wBqw5VV7+F1MDSIIO2qSLn5pQgkG
D/ZJkIUYue/wpFlnm9DE8O6C6MtAY6WV55fM/5AVfO6jH2vdwmTL3PL5cPkKUtSl
/7VggDnl8YIQEpz3yE/lEOs8P6zgTfeu8AlRkXqzQZVT95MPSbkHfrxCPcEiAd36
x3t09AKPDsMcLUGEndNDWyon7apKjIaCkKcpFFIksx2PpU0+wQ/yTZ+O7pFNFHmC
irE/ycx41bEJwVTYyzVWFEknEmjpdp7fGvBEeyWjV96hRRLpw2xVfYywtAX3U2JV
zGXNNhBF65gshBxuueNXB6jHekMsAbNvPo+hF0gj7xQRz2K28xcHN8dfSBmzvwDB
DL1UKsS6j7RWZrRr4MMvpSsTnTCQRZzESqQ2v/PeYo9cD8OYt79RwodRqVT/ga4R
APi2VvGo4uLKoYhw74zwPoo/N3+yC0QphCP/MS4hFKShRYdWFRipug5EbOXuoWMY
JsG5n3wJzFIyoWW+obZUTAaJ+TTAfuol2XfW7TmScUp0tUy8Jz1xizkCC5zA793h
uE+reYsE8lcxLVpNtMNnZHlNqtsaZUGBfVwB52DlshJE2qVogsj/xP1HKCEdOgTR
8ugZzV8E1CxmuqrpOGTakOymFltfmYpopoJzzWANSeV75uW5qJvwLAEgS1Gq/yvB
/bIZalHpRCE4KuLqVw5khXFYDAoxL83SoY7DBJXl2wwqK5o6LeGlIrNTzIawmPX6
xW1loXOi06dXfSm2/ZORslGn0XjhQ1DcV386GcORUfMY2n76DdOC1Y31PDsujPtH
LcGxaZGAphWoSHOzGWqczShaa6fc7ooyrSamBZXkISeOgnGMxD85uLIsY/yndqys
AlFU9aT7PLeO08yexsRMvgm6LI2LDsn7wzVpdyiJ2LIwsjINiqim959/owoH5YVd
hOHToLxbr2ALwZibLB+Kpl1jvG45DNnjpcU2gW/LzucobrPIdVA23j/pXqkLWm+v
yiq2hGKmpIVVAhJ2dfxDoTHmBtQuMgkIQL62TBTR6NxB3jHQ3Ps1hRAYB8fm1YX6
Zr40dXtGqAjOo0mX5WFofuc0qWA8MEOKbTSEVC8++2i08buK2x/2XbhmRkzLqH3y
frC0B0p11WP5e6kOOlGkZrChCsbVdkf+RfPojPAfrP4Y2Fru39F2GS5+yCiZPVOf
WTHN2T7dwQSAkudaO1gTdx7nd9c2qpvUlQGVx1hEOu8TEdGGsg3Wrq81Ev56ng6x
xIfGPUWlF1lDquQzHvHgjLp1Lzpki71TdQX8ghqnIqNusjNm0ET67ZTavj6hRLYe
cOlFLbUa3A9WvXjm9OKdV1UQe9QZaXyTmyUW42PiVIhc2xfKEZuvmG+Gz4p6ZMZD
ViGT/K+OCexcbEsxKoB1t7OX3pKu/0O6j3g2+WL8LtEGFyLunZR4FH7Sb/3wxFJA
MpF5CqDCUqdB7ZE9HbsaRioOtFRAU5JedSldQJr/zJSiYRkvZ0knO6jCly0TrO13
xm3hGrmUrwnRuFzwaEiwl4HzgQrRgS+R/SbNPg1rb3w0IfezbYiBB4FBstSNDno9
U9PQ9PUR1e3nBYTmz7wuuQ6YBiWQpUCgZQFWCqCrM4VE0HTJRIBV+QKdDilIgBMg
+3poRbQ6+LCPczbhwWPWc08dBG3lB1zTAjEJC7DSo7vv23HXUvpGcKNdb2oihmT5
prhYGGm8dZyhsHXrFoca1+d6D+XNsG+jFa+YjQbzukkRAbltEBnNKgGb6tXO3BUi
Qx1XGJNTnw8IKG16DPB2rjxAHeFr/es8hXfNCusKeVWFo9faojiOYJd/06cSHoYF
Clh+8acGTgozGuFXSidTj/dvtESUnxsg8BJeJUUtJs6+07UNxiTvFjoBZf/HJwCA
LzJajshnEmEwOobfAPxd6OlsGebat5HTXqHaHwGHd3Zc8on3e/bWov8FLNkOs+kE
19dFIPYgGlnIiviXjSB4eB4mwrlYAUPb8FwDeshO7PIyjnU4UaLVbuth4SHNGGob
3fyr8MRx4sn6uqs76nTUm3DzaQHUX1HnRdGdGA0EzOous90/LUpQ5z9Vi8qwCiQ7
mxaLXazR0IMPvmRLvqjUHC/Qn/NXUh3KKXamTcwH52R00xr09yu3op+AN9+8iQ1+
e2k32Af8yMnO/dO+GtBK3YfQZE4ni2lGHQPRlaxPB4SIOmvnpFftEKNyfwXMFdZS
pmOz1dd0VllZqeLznDEHkcUe2lvUyLdM661rmvcTGFur2Ten92djMNyjUY/SJT+D
CmiagxOBCuN3ZJ1Eu9AUD3dOhkYxThGEeqvyysPQDttayoQJ46VA9pIBoMJ///SI
zhgwXxdqd7pTMDFhQkji+1+3cmWbvzviUfxBYnwsuq6lLCK0SqkNUVq571AJELXv
Gu1BqBMHa27srxkkX59IEhsicP1fOn3eWiY2dwFcgfj9dSe7PKgLfZKVtnE0hZDM
KyFL6VZA6CseA/NUqC/uhKWrFLSj74mS5N+0bl2OXWPtyYYYfwtpyWtCDJqYIaNu
2z/e5Q/0xakGHxGBarod79YggqjrrrmDM40XaBWcmpnvED2/3RbPUDFxfIBGNMHr
HGg/ktSbgeNVmcQCcUZpbfgEqNoqMsF4NXUUScLH4IwaHu/t7FGkFKEvjiBDR/qB
nH+xjhT6nb/aJe03OaMq6jRFeoyhpHOeTCa8eMJUh8strz5RN+s7kV+3oYdWqKjd
IMyaeuBXUlYv2kJxRFDEMAqP5TaPtOyGnAi53sjhhxC3XAaEnNk4WlhU7LUXR9no
4A1kN94eOUf0tvQ2zNUK+FCuN/oC7x/HpG7CgsmnM2ciFvblEzx5CsqKfaEXIxcQ
OmX4kilioV1KRzC+rgKiTxvzbNAtCAe/v+5gWviYODr9ExvucO/lG4GU2O/u+tOY
dlgdEpCpILf/qvuJkD/Pf18XXoZTjQSdd3fQmlovub9Hcs5FDCklBKJfzAtzqWid
zY5w3X0Cl1zP37LPI/bdamP+JuA3B0HA7QP5HXjVsjlu4ZgaavcE4hQrJfJHqHbp
EoLuYYBH4RQIW89ytd+Xi369WWUXNchSbSvBO242NVJkTHBNYEL+3zfgeNMiVrJP
y0XwR9xGKDeSGE4a0lcA21Ht/FMh1NaMi4Dj527Mu9vhhIw0A+rRhL6VPFtdRi9M
/28/5N+HAtjx1nRQdflK3zYa59TyRz1bIrSPPvmgHtgnucTT367R/e3sUNwBQUDa
/+jExRojsQ9pTZTUWKtH3e8Jj9w9tjActCkokaz5Keqg2sp4GGbHhFO5ORWyPuk1
F7TwTUvxlq0WRWDLEx+co85zvUvagJP1rKMytX9M9pa7GxQdEsxf7oR1EMVap5do
eIRIGxFqWSbOzeDPEwS1SNvOaB0VC4ibBt1QRlCaEc9BFkHvmY06AFHEc9h7DJ0e
OZcsavdFMv4HM8148kr8N1inbD0nRNVwkj0eX3FnpzJw7VFKI1i+G9ZsBPOPi3JP
DAcQ5f9p8ureVxWAMS42YZkLClTzki5+w4lq6ipbGg/ErsGp9gYsE2kBv84eoeJ2
eXH6TKW5XO+xX8LExHmrHBod1W7+eokhqq6/Ns1K4YYnJUhsyXYsxXMpJp3Xrqzc
J1U7Wv+szxPZ30PKsyyY8w0UO1tgfPXTHaUP1DAroDxwC5aBZUSdtdRXyRh8fd11
DOuLBz9Tss3HJq3u/K62HYNQ/qC2B3FkSkO0DFgQcpXgrMuWoGBwMYLj/jJMMp5v
dQVZ5LG8Ic7ni44k6Noo5u6nRmJImL7v/fxHYq/oxWHYrMhewWvb7n6GfmtR0bpl
mS3tTHElq4c9xoFa9FJhGeg/0bwg5t8n5jcFuaK9PEASDJ8XECcYiMpDrH9QpIJv
KbRHi/5a0PdUG5mFiRiOlQZUr7BpqJOT6fzav48PMkHgEfZ7+dsfcA+IdtwwFITk
tegssbP0gCxJh9EJZna7U2LML1JElkjnqKf7rTtj5sg4sqrpkipLTSEXy+q6mOLH
tgV97JkHbWJBncCbLX8LItG1ebipp8SXdbmdTRp9WosujZcMSw1TlyptcB4tOOJB
WCe7aE8Wm4Y6XwIdwFL8BPfz65wxezECXbDLIumujk1hl8fSHVpHyKHC9pTV+BOv
GRHMR9mW6M+sWTTkvlzhD2rEwjvHOSPs7z1V7YHZfQtnspjUFU49F6ZSitIl0BfI
Q16IiRXGxdRofOht0SarufUmnQc/jJ+oH05JeJZiIs/5YKP6+QVGbzexUIkXeSDH
XjGAsdxu8VtcNJR44JMh8dwcSaB7ToxPQGFMnCaDcLqCi5BQp9w+Aln4k6KhikcG
5rqHLXv2dlF5eVXQP66sYUgPdz9nURZP9wnLZ001MDQEbR+JhZHazMJeoAK4DdmI
m8Q1PdAHa8tBApd5MurYw9ivFWEdFG/H0R0PTCExadiihbnwNYX9fakJTMerrkFl
P93QEWDcTTzwZdzrfPAz6KIBnSB2SQtFeFFRuTUrV4nFS2aeJYfjtFGZRVyp2+mp
TY3IHcPz0DNDFEwZknIQ0CdC7NFaZuRQVAaoK0NnaLReDtr4WZyVFXqXpvOrmCyF
Swx2sUorrN2/hR9vAomq5zZ573+LmPUrJHYaWpTDSm3qWmBLx4t0jlNcFqAL7E7t
rQdA2I1cD8mFmHp/P9nHna9HHrPGKn/f5o6P2VMle9oH0DLXiLZ/aVbIN5Pudayq
qxUQTWoq27tuCE5R9QfCaUri29Xz34exioW9jlyU/YIp8GFGzkH2iTmZajQY5F2m
37p5T3PZNOEnDLqo4c8v556UHYlojhtCQemkRjRc99w4U7YXZ2/icxVM/qxZ5MJT
6/5zYy4/nb6K1Y7NXET1qQ/vdxLrbspFgwbfve84R1p6t+aGWaG0C4tigtAwxCHB
aTEYW8hRX/zNYJT/wH0DOn3FlVH4as5z610Sygrxda5F0rEwNg9I0yqRZekkBg9R
iQMN9sfGuUK3GoeUGqYb44YeKWIZ8ILCWJiQJPgM9VY9kSYEzXnBdewFtCeVLcS8
FOgsUEliwf4JA1MtnmT/7nkjeYIFvV71PvWAq6kKYsnTHVSTcvMN3S5O599ohkH8
vc17rS/lnLtDcmBxF1vhDBB66CCqxaknbabqyaUoUSdlID1REIxsCcg7PjtRKJ9T
usPm4tGcFOCKpsGyRDTeUN0GVIXDsstofPXRvT4aJgS2K5RIAA7FBEPGE2DxK/1w
LtUw4gHYOmua8yr8Sian1Fj5S/OTl5S9Hk5lLG9EHQbwRcuVznOzwCqyfQgnKcGO
xepLoYriNb4dbNkkX1BcExrUGZwhbsOJcLLD7DLZ26zag9UwnAUTXejoFIbpRdSv
6Xylng3O6Alyu4qybkh6h8O/ACwSNMBjwQx2bajcmodx0SmFESv4stZmDQ7V0ArA
gMujFTkbiKymfRMs7lt9QaMCvpwFED3Df3Bh+Gn+/hcZt8fTFER+DYaxBzaiCKWV
iZ4EJH3ukl1jg0OUDg1KGKJcNgnb5oA++VT7Lhego/T/9viv5OMhxuQPld+tlsIg
4HHRwVnmJLMxiI+3/xS7dT+li/GoVVk8cE/PhoBH9ZPDiBaUm8NHpZbx+NYsrqPo
+No++i5vdYLjELCBAb1ZGsBphOd7d6E6FRZfc5VmKj0IOcytcXhQPFM+XM2OKWc/
05i0NBL7fpu4fEHkY/rzSYORV3geisHuWUymHAfMvaIGBr2KUnzrSsBaS0x29mEe
4TMXP2QmWusWPMDiguFJO2nudyBzUITPY/bCx/rsv3zqUMVVGTUaKfdvk2m8CdYT
5Mu56BVGlE2It46wiCg7oeK1sWePaNs49Sj+d0bGoF+K4VvfYtHtL2tPrafvOD9v
XPJ4NUGFNgqfIE01NPxa8z0E4nrBn7VOaJhf3ZVridKguO/BvB8ENZiaah0nM79/
tp+P8vXXztRLw8V0LBzBWwnXBiAQlB7ty/6+ye6JWVf2gKHeoPu5dE9tFyL+0gig
8PLKjrCHQ7LW61HoJYIJ5bwa1qnJZEfWDFC/tHNNelUC4mmyq4pIhUL9ZagqxGjG
kAU9FlndDhdsIr2NDMUSc4b6KBl4OZoidjHse4mDZU42/KG/VqsTGWnhID8+6rtF
Y4+U1+gR7K5k3wWKfHa/NVkLc2XsY3eJJObiZVZ8iW1L/C+v4XW7ug1RdkiY0P3n
j8/L1t3F9XJwKBQHlufV7u7muEAENJZi8ca6MvoZ37YShoETDpLFT80oLClQVASQ
BgcteqedWHunW7RPCAV8wAOGCBDgD/FLbKQU+psI24qBvPyCcQ+K19/zBQHZ7nvo
ZMsQbX/CkOy70zBZhKtJx3S6FZ2ETL3aVY+B3P7tLibHIoiQIFFfHRrw9PonSJOY
HpQohsjdZ96dr61blPTwA1LiyaR1q8FpE9R9thX4jODPgnx68MFlQqytimvWmcv/
Owr7KV/atj3jzBfzC1XAjCVOS7LikhHqG4fvkLxKLf2HeQ8B1lRjRQRlvQ55kxEw
xnR4ObUR/ohMlt2Rj3FmhH+kPpZFwpTO0JMOTghJh3Z5FG9RcEKsKYAupud1OOcu
ovGl8ot3uOmgcwCzB4RMiOz9ZewlAiNbKOZ+UEC88FWjFrCP1EP0t5qBj9NxWth1
RzMNuMSQ5EPlpYATErQnqKO8YdhDJXw4+6665h0CY8f2Vf1FaV3ys6NZ6StE9nz1
K0ZkwE7VIEvFlM64fD61/IkcTJylh+Qf5IVXM647tq114ftsgHrPtWI6ESIYM+qH
uQkM156839uKbq/06bhbqwOxaJdKnZ/+6JWXzETeMAUVsLzf5ziCemcjOk0XdW+A
SvUXmJuBWXL1/wBT+XN9h8fe7PDuMRYlqlMEPpZI97FhBXGUl9kJSmouW68bZWWR
J98jX6y+8TgWsdKgIi01QOZ1UAYi8F3fdxbe/HIeNCWlSE/sR+gkf7rdLIpExlER
W5fTUrygc0iIy0vHgD9IekxD8rpLm39keKXpCPq45v/AHnzzPPInpfJ/1k6Pjs1l
2iWgdr6kkbD78oOS/KNepWNZ4qGk35ZT+2pojEeXlUMEk7I97HVmqQsHwkPKAseW
6bmcJCDrdKjFO4dxql3TzF5e97g5lFa4fS6VoL4l4tnxWNIEhs+ck/MWPUy4kBpu
ep/YDdoo1N12T8dAWSrJ92DBYNiKnSberb87N1+Ho1D1gBSj5KTWgKRT2D+Z0C/k
IL05Ws1XJD70yYBB221wLD43gWmw90PwtUkEIJCptk7bNNktoeSdhQ6CRq3kX9qw
gwUUIPig94xb8/KQ1rwfIXjyCQJeW/LWp1fW8OIPG95RadTcKik9PEVkV4tNVhk3
3LxMmJojTtBTJ2Ds0CVLa41Cy+fIhHjYeORV/wchlDq84jGGspljbdaBkO5Ua0FZ
CupIMFu8ol8ZJBKMDDbbzTy2k62RglebgAhTZirF/oDGNmC+jLRHwvfKz5Oim86c
HCeMPUHcOiPNwtsHYJ7Ls2lvtp7+E9eJ2pgD0cjrhEHMPmGZoqbuQaCQvYRwYds7
9XquqjZKvgZqfXWnGaPFtbEDdOB/yAyoAb5BxXcGrGHNDQcMsjIBxY+akiQezP5/
SSbeU2LELhOf9mlNVld8rccDfxX3kmqgVzeugbDHff4yWEOpQv79/zuGwmkvwAgQ
NktSHSuCYtKzorcdsdUdTKU4Utj2VIbeShW2nqd1I8NkJ2lVde8qlVwRtbd3pMm/
h6E0QnslCrsmHLpQ93nlU5T7Cv09Bv3+401b/lTl2TidibbjstWlQSV/MK4IhYd0
DTMKcEi5Xmt5B/5ghLjrEglwdjie1YbrMK4IotLGQ6/eZIeULvmIrIM19yK20eW5
qHdYi7peLwgItZwQn+/GtTZ26dI7y7jeAkoldX6BW+veApsZvZOwjftVYZoWzhIW
Yh074BnXjS0E0HvyJBuNyq+8Djf1sQLST2LX6JLSaGGl4fqN1irHwLRwXmmV9Kvx
3eJJaPAEblmwr0ddZLXE5zq01TNJuKT3dstIaIhhGAMn6AqsLhAnZ/HGF+jD/vn8
qIGXAqdwCmN4pg5QDqAbzNqyQiUtVHYfRgqccr16r1JOyeifW14oJGKtLai49hax
diPoN+HEiRvNbllFZTC5f1NqFYmYHnY2K7p8MCc3b4ZjabbRcpg11MnOwIFwiNaH
O1Lu5EDsqA8eNi3mhLs9Cc+7/1ahJxdZSvR1aDLxxKkQnLUcvdyAv/UcSqmFKHTr
b3rmwGJo4FMTxaX1UqWy55TcURZfi1RAHaStHbWcI22zODGiaRnGibLAeGTgNv+c
hVrheHqOFIryc4wMc58A3nvNieP2RDvMvqb1JFP5f22Ct7lCts3A78kj097dLUUZ
EUb7kYNHSUBboO1tHEyIkC8XeCmYccibHHL9jNLHSVbKZdvykXiuASfP177QJqAJ
tRXOM0WKaXeaDVpCQq63Tpnw2Dnj4Rbw2YVAOD2FC1Z6YENDnTHC6L6FBm/fezhV
P1hGJrWFan5KqDK5x7QbfIIarkfO+vZL/SSVYcXY3yq/poIb4PUORyoSZ/PHBHU5
NJ4l/LsOz8gZREYnRGA/T9Vi0q6UxUc87B/aIk8QCgID3DlCU4c0rTgXtfLdKfna
Ku3TEBg3TMIgBeLHBk/FJkGj7OYSsjp0YJNht9n9cGqKoUIaCoUBCfbJ7qsHTuuw
ziLRDEN8tRRBJSgu9LIvVK9cMYA77YupDnzvkpA4jGBgsKDkkTcpQbVnRKV4t8Uo
yKuhUozXdmQh/Nf/ly6RTYgWDj5OBsUvTqmsA/wvglLfkAYfw1gSfwCbuS1PL0ve
tvTPdrCsPajr8a5/rLmsSjap/Lhwt1lD5dhrdEmtp2brgKU85IwanSGAJecP3tZJ
lml9xNGMbqDUZxae4Z7xrxKqTb4Z85hJ6laUoNsWhTeAB46+WSP4ZUFhwEWd175F
kVOVXUZwAhaUeRG4dqvCoZmRsRoQOC7xbR4+gBJ1tC+HSSl86J2Ovx7vA2MQGbsa
8XR2Z96LByLY+GvQBg4GLRie//6OV3Y8wmzdwxg2oDsBNr4HN+y1dKvKurPOlbZG
oZ/13Vi9nzLwPQt8360/y3RFkTpgVCRZxucDPVqWIRmXZKYE9wsVrMSidUHicse8
XYabkhYif/CJ8hUb7pcHOT3LnwnGayU7Xpc6EOHJauqXYcuqLywZvNMiNj67D5uQ
8JaW+yYWmte0gbgvuGgIeUMRLS5859kupbFTRcZ+4n8htyzcwQLBftembuMPm6dO
kMhwbv+sT3EfqHdPZPz+HxMA9uUhTHrWa1CvVAyRy/s2rx+1iccppEIcJjpnomS2
TxtRXTaf0rGDAGfO9ndqi1XgoL2YDgwA1JPA4XdQSWgrxYEP1b1Cup5bvZ318p7j
XXd0nak39gXae4RMHGMLEn6prAcVbytO1qtde8VlbHhPyJeSEHr3yIDMS8IRVvEA
QkkoKk5PleMsrE1EVZycytDdIKyxEw/DEiDDyuPV+Q+HUyLdRMD27IHSbl/DCfP4
MU12oUxjOGB0Rw8uXn6M0DC5gsjgWxctVe3VFNp+qA4pqRkJjIPcCVktdLbekIT9
Bj9ZsnLsPbO6oiy0M/aycvV2WhTfMHQJt6FMWin5FGBsrhbs6oX7FV5IrnM2Dmus
xuy8zQt35m/pDSmRrjVmAOCWzBTc+AijQ6TKhOs1XThPnN4ynJqycqYpLkQQPuro
oxa8Zqjx/3GpSm4LzT+e+FEMB1nTHiX6cRR549F82vQEkqiwovxhtYpnSPb19oPQ
EQfoqk3+NZv4gslFkVqe8G6n52cB5IwTK6ZUpLbZA8AoxHAyl4zhiOSb1epbF3z7
dkNT3CSgDZ0sSfzmUAHLEZNdJUDWX4d8yAvIyBzhTm//vQzJ8r60Ifa9tVGII85g
9r1AXr39AJi8B0DjvyRYTlJAZ52y8/ztQhMha91qpnMCM4B7qavJXlBLB+VEOrTO
wcQyyOmRznfNolHYsQw+Oqun8XPWSoHLXa01H+9Ye+/+O5z1LR/IaohTJV1rbyOO
duVFsE8wEd/dizIfKCg+ce4kWy6lqTnuvWiEnktgaVYhNNJIDN4sdrRLEsXaJw7q
WGlfexoOQF5E7PfKC7meGbFJQGYHO06p6wfoMs//dM8wcLa8Rrdu9Arbv5pSiOl8
SRTa/Jndbszazy36/boVWINFxW4gT2GqeqGo0T3Age1SzJwy7ov5xVX0T3sTq4PQ
rxA6peN8GZl5VnkQ8/p4FbXJRM3zZ4R0MucOh1bAIcsgE1KIXVef+V+mv5wW938u
X1sefIgM5eSA+zNCI/kJ6l0V2LTCqbTESlfzN0fB7ArU3JLonf8ar0YTq5/847cV
62Ng1ECbsWeogwmVPStuMpYJwPMd6vX0qkRzWc7JIhxtdQGUVVD2Ymh+gs6LmX9b
nPIiOFjs3pYyd+93bLyAxVDhikFG4eQl+Ap6xMHM7u/ryiNA6YarK/WMCNQTM9qe
14uKackYlsEpp9AA8cPdn2im9mGPNNiomjNgphNSETuTHmnH1WsADeu81lQqJe1J
Xwy2IWhlcdB4QjeJHuftqafZFRQSTEirKkpu6Om817bceBEtZ1lcvyBNPNR7mdre
lHRAh75dwssvGSsPlZohzn3kqPfyTuhlTCWVimS4vCpzMfIPgzJ3wWQm4JlmzfA/
59+STn8P7JsQjGI+IS1IRLrh0iDtQZDuanF2vu4J7Pn5J1isCKljYeKliln0gINP
WUvo/e0HJCrHxNRN40gKnF1gEVh/ZLHWo9cs3oZekxCozJbFeVzbD28iKCGNZIuy
aKLH/QLQceFWCnNeGm9vjGANLZ9yVZ50aYnVdW6r4aPnQNpJvT5m1bLd7gsIXgtR
rnm5L+EMPiCwLIeOTwhnVnh/LdX0oykZsfGy+/Sul3CSZJyIjWgHMa48zBQI7NbI
SoUF+uzKlGCE4ua1TV2afHnvKTDODYmEjtotW6yYgqNLPAqm1sUEsQfClxifxBeD
wJWoSwEknGSmmF1bjuSpcJ9RHySQ4rr7yK5lbNcUrGpcwg4m7E8KO60SJTJrj2Qg
7vB9Ryq8NBwmhoGhLsWjLcYEX4t8Rh4IdYenwp5rJKUQmZfMA8iKf5xjmJNl4St3
W0C0GTbJ9g7d6h+wIXiGa1pkaP5vF+OSV3I92O21muv/AhozKN51c8jkYJHJCg5I
a5WAGCxL3YYfddr1x57Yb00+Ey4G+5Rg6BRAI4brfXM/F7ol5N7wwNlQxWaDTtzd
W/QMju3A1yiTslmnhZ2CqBtZKDHJk9a21ElIBIhze6nOt8ZylFyb61pnpmb381MN
INfw9feeaZ+I+8IaIDSRe0I3DnJebYQWJ/8fiY7B0OLmxZYSXzVATwjldVyw8zj4
Sh63vSNQFTcG9eMlGapYr0NNwvQSP4UvtWVFhV3z5tAM6+n4WjgDV3/ec3++iL6a
WuHpHB5ISOx8lFQaSL9nAINmU5YzFqepaZo4wayzKHypIGt4m7SoxhcRiNPUrkhi
X4pS/vy8BgY/LcMYpDDrQ61BxgJM3CoS338hH+BBMhO8eFCxOX4MbNTjLDwJ15kg
FbAzQBHOHTDF6ww8JE49WOc08aiWTZkPdD2BAtufphfGJfghoj72mZ4ILsVX8/RA
0TJ0Nhx3da9hIQYQLBq4bk66jOHd7mR6GHgA59xz6dqLUZf8e3eKjvPXxi9gS3/e
q46ionSm04+c7Pb7+6/Io01d0l7cGhLr/otSLW6Lpgrr6DUsygAvypJnBApKwAy2
kSdrDQp1oD3Fx8qRfDjSZLJZKTFdi/Yhb/qS8PovaxZsrgQb/RQdW6b/Pi0XBiM6
Zyq/4bdYau3DxLY1U1q1eBlviWJTcFhFu0vGCBo0iKBMh2Wsn1UIEALF8P7uYlB2
KjDVnUaplkGu3UQGCfM2+BVQ4DMnARQfukN/JjMXEMqAtgg59hE8a06wdrnedyyg
5prWMGn6q6O2Uz1UDlDq+ciREscMLzj7kjGXoj9/7bWzP6Gz+/nTQXCaIKS7giYt
R+8Co2rudtgKcXfADzmctfqI3ox2a2GHN++7BOapnS1JR6y9op5ZsUEYLeydgRjc
aZLbJxOWq0BzQc5E9T8P56zdzy4SxefxWFS3GdjoBWmpMKkHj+GxaKH8J6FS6uH2
k24he+vDuF6DzVZbkJCZ5NUsZUYYy/z0JxfeJgQe5PVmQKOAjNJhjfiSGpnPjG4b
5YZW0+VOC8F869ZbMTR2Bt3b8jt0Il/KvjRfarPSYK2GX2+xB6DZPXwQvgzCMkOk
ELuGhDNRtlVnz2sFrs95Lk+1vEry04ZiMxDG86Qa5nLiEYv9tRsBYpX4pzRVSRfe
yQ+JMKd5PLKrDRjEFd90wq3LgA4Iva853766sXzb1G1oe8NjIi0STiJxaIKA0vHP
1vC1uK3XtD4K6/+h9pRslXc6p9omjfNQdNGL68N3SoKS6dRFQ4EfTiiqj3x4NxIv
4yWB/mPDPxtsNHBCMeuO9jtuDsejgGHVJ2DaTZzks5IPYqiFkPsI0g73vtIFJerV
ISwArEH2KMvkakOYDeM0xmgf2iZGGZZddbldoi15wUCQvIelJuj0CXgYcuxidMH/
pfjKBEodEqL18xw0TSntU36sbwztM7xOnYz0yLKyfOw8yILonyzcUJ3Z+g0tKrON
3VuBTcIZvKOny1bLHBsZhEG9BYDIudTav78g9jykcOAGyvvnw1HAWo7fIUON2dNO
BPqgZu/sV83tcIJ6rsIgST6lFzNPXF8w+LzpVFyNMdF3m4n2wcNb3eymKr31xLWN
DcsRvEDVpWB0dDEA/L2AZdtZlrgwVJBo/XyFZIgWjHB2AfoksL88hSWtkXD9ruVd
BgAUXPK4iAHWtvIKJsCkrQXY8bS8YS9ASeeZ+LUwLH8Uszak93NxJPYNDNcFvpgR
RgamzulPY9V/HmElrxz9d2p6yRdoY7vkIBO5nWGxzyIFlmN+qZ/cXiJ3SiAU8ewP
w00tX0TFQiY6WfjobKoc2decL1OAzFBgF5jSebXybeOAmHRX7sAQ2yYgSTYTf8gV
BwJvpmhdpmxTVuryZoh4L/2LTSxG8RFe3urfRLKx3U2Mf63xPr9O9w8lHhRQnnOD
/tTpwzCrEfvZG9a5It2ElRC59aKH4iKz9x1jvCEP3j57q+oBW85H6uqcFtpWC5hc
s4kqOuXvKAV+bsWNiak0DUoiekfT6zrgBbH8bs7YyVXndCfhD8qLV4Wsjr61empA
GfsOa0rMh3LJxhDHErUTPAPMUpBqJZ7+kttLwg4Ljt6TkI4t9gsTl0BCubt4+Ir5
URDNh+97mXuvIC1O3blX4WYM2SCu8pdg3sV+lFkJAe1Xqxxoli+kpc6lAa7iqYOa
NZR0BnZaUXAZgX0OKhz/W7KxlDo+6JR3bVcd7povdne4TrmNf1X5IF50CjOFsGcT
RjEkJ/cKOFh9U1KB7H1nBysUqqJs4Q0Aa7JRLqsSIiNUxZXr9sQYhJzMwN88VvSJ
2gXVrPUyPWbtZqA2txCgzLzYLXmW8jmFkRS4f4xqlS4lkk2Lc9otSjTQx3/GUNFs
VdAxmpwCmhlKkmQWUByGsxRicgMAO+9RjFP4QpJ3nUaJBrrM0lgXpeB+WFCDjaib
mfWI6rBEtVjPWBqRetRhjCRmwPbOSZHwaxxpuL8L5Eucf71bF1V5xzex1dSQTcjR
GH54yF7eud8zj/iqLPhqB7SrQgRtL2qqpoPypzGvJ9CrCXjJp22N4JKXSjgTbhnK
2KqFSZET1dNjAEo5InkL1tzdNDRDURX/MP/VDd7It5hxp9guRRdE3anuJn1ksfFL
+QycLmK5OgRloTCHsMbhioTwZB9HDgIl++Of+dGY7TJP1SGR+4e6hD9uKsru0VCx
qfVLoLRxT8+nHAVF4wb5qeOPLPFi9j+l0A1rFxI763b+RXoppMXSlksHT+mvbjrV
z/iaF2QoG3mMRLHpmHNZt1uZR9ICKIjce5jQIQpUqhCCR57UgkiXLjD+CKPJOSbz
LiplYV0UrbYU01eJVJR4gIP4/guiK6sJ9pu53huLuYjH5Hlyze5ZhEoB7nax7OHi
MCcC50o9hnnddLjmjIwwgmkSWYmaEgcONBbZiB+Dp/5GgrbK1yTEBMbGZchF7PoO
keal2kOTUjlqBdYKHrv7Qt2ozxv0aF/eu3YpSrlxrsZqjq+vTHgyboj2VTRVSO3L
F3SauQYuYIPjYLbceHuoDhyJ+u6ai3wctBtB4B94yaQCjH8hOPH1yGJhC6SC3ZRN
7IEe35mUeNG2zQYtBHAeMORxLXXwqa+QJgtUVzdCnY9Z9oN6ObjDJ2samEcz6iL+
8xhIsNV9fkUFUAjyj/mGcSOtFeP0mlMYhWcn++Ne+2SMi8J/xQj2EbpLCrP7O7Kg
1zTTK0XNLWftT19tg+r2Qvt/7xq7gzEJq+gfxZ+vrYJoVl7TKLwoDV5nfTgD4mtG
ky1xTWQSSwXF+KybmwZhtf8phkybC51kedKVNPVQ/fSIMYuMpVCG3V6dh0PVzyU3
BfoNAgZ3TVMCIk2ROAdTQVmWCG42zbM0PfsBAf5OaGzCBLJIzIJM8q62bbGuiip5
nW7wasNoJJnJ7T0Er5HYAyO/S4LeW7xa5JfDbAh16n/9dpGuAHrCOmar+0XJtQX3
eY/gZTB9ubBLl9QtYuSJUSrDlxLi44r9jJwb6KQWV2EYxQVtquZ78I2rRvAZcKpZ
7FBUYLSk9sTsHmhMnUYoJZy+P/JATvlyBj60LFMCaL5n6z28xZiP53RtSaRobbcn
9LG0RXYJGkhbm7i7ZrZWempLXKx8m47V8Hpd9DG68J7dubUru67JyXmtWLRUEMd7
2w4B0y1KZi1fJd4ug7Qu6bQhLWJMgBJWuOsNI3Ukb23L4t16gVbzBptfQQrfvbrH
cDmPH2BZ6qmtpXugSSiF7e7EmtQawW0QurFX6Y3V3iMCOcMPgXIZ9aHov1S7zQSp
BxEvMT6PfDK1DQ52pfBd1yUBrjKvrENY+wvvWxy0BOoshjyrEO6iVlrf+rkyhB3i
pmwV7FAs2GH6gtlgihfRV0SXGTXT81t9PPzhLgsvSZf21YP7HjB9JuMncKMcJq7c
tthDKJnDCeWwIil1POtekYWMsRGnE/HaXnoyRIruXDctVrbrw7a6PaHsCptH+Fyt
1WDDTg701zFJSFGKBsea4ssOoZn5WV28N7NPDeJRHvvjotKxOn9bcsocl3rf3im8
LmdRAb/fRc88hRLgTac1JuF5oHjLna0tMBqq1P45umUd8+QIWvIIZq2uUDjVwqYE
5f+FwcI7XszWX4/K0aD1mEINP7id+4bY+Sl6CrR2yMRB5E6GKLDgUTao08NxTQwz
MIjQ8i4IlhswWF8h/OFwVVMLByrDo8Doj5TLY1MADckKPJoLZDRV1xakOHEvMeqR
cPkSJqkx4YxC1WjZXzyb4DgV+5sNHmowTSc6JP8A0FmjQstq3W6Dh0I+GJwRUXwY
bOoek1kBL13MeYVkOui0wWZd6r0JQ9wbLWG13fzVt0IeSSVVxh74INZMUhi2kWep
3YMCg422xlaLTCa6k9gWnMvU3y3hSNyNZZ7OkCYTWXBpqx6HuDP33gYmey4/oYus
RW4Kis5iqasUg/GwD+OPJyfCMhTAH7aINiipmZ3TQMQvn6zVq14djV8Mz1GPdfKN
Cg7D9RhaQFcTk4H5o4oEIVvhMgqh72+WF7FG8KGCMoAsOGuUDvVMjVYxNx6ywLl6
Ly8mWN7gGu1WCXc85BzbnTZqQ5maXvFSX+T1lCxFLzR86yJh7Q73LpYRh3nMgq+R
xJKmQvwqPD+9p/mO0laQjkWf1xqD3ur386s0GvdUd34OD4p7AqJbWZvzgJH4qLOt
NYUP8V1FSD/lwgP1BGCmRs8wP92pNQNnslSq+K3QA2MEPj9rHNhkFAxZJLNIEPQr
PwciR9HSJ88zXSRYouUzUunT7AUoILev7vqHOYZrfqPFmD4wc4Bh77BYDGYtM9iA
tvI03JcAFFnnCVw7LHCQ41Ckutc4BmZq1nWcEYYHogEpSRB6B/CgzPpuSpG48Mbv
1QgK4VuiwSRzdG9W7k71XUE9f/rr0p9qKSIG+2tiLjTDFdGtdohhhCY7a9J/26CA
wLbW96FL3UbsnO9dxq+p1rMke5VEBoxufhAND+mCSRLI7m09BqGDncw8RBHbvFbq
AkzkSmskqBKUYiTt3qQWpOQ5fYk1k+7oyX/dWtF+Fe2pqDe0YRSzVVJpVa471PyA
10iUS1g628O7cYGXKBCmPPPZ9+z3KL+WNuRWW9PSKpgmJlOKCS1Efzqs3/nQzM2T
DoXLBh6Vcg4rFEaiIfkuuXifjOYZfYt75WyPepijI1IAI2JEDjBdbvaqYdC+NIp/
HFvCGwM/eNlQe9zfgF1XT60/1g3dehyEK3EtXbKzej4kVhv3m73DiY1TDOIT895Y
cBwU5JchUE961tWIYZmRvwayuvlR/Hjk3SImHldPwoP/lM2FEZTRjk7GAiG/oe/b
UfBtY+RMGawE3l6MONMLbjXxBiODTam1Xxgw0SZdJkW6jvjfibgDZS9TFOc1LYjE
75JTY7Zr2Tco+E2JDBW3yxOHcYoLxz1N+b9XvJw+0PkjydeJjycftrOulEAgcLga
DAVWuK7NzezgFDdmx2gg2ox5abDMgftoTVp9tU/AyJQo2KpUvoqRb+TVN2ABX1bO
w9n77BXpLw98Ee8xKEJ1MGHHTJenwTQpQBzBcIMCq7qMI/9qm3YDqOg9HL1QYV/Z
bzbvHWm3twirfmz2lJ8qbQ+Tzj9LjFCCG+ROjgR1q+xCuGF+mAL7T4P50oik9T1X
qnHyDbj1IbifX8pNTDlZ65Mwm9HLOqwXCietrxV2bPhsStsRKj+FqvR4RHfvFl7R
zOAop3vcK5zlE2VXXrmfttcIlu8VMRXvZtD2hgbpqgnvC+BdlkH8mFMcCZZMwkrT
wkZKymZCj7bpM+yVwP3DykDxl8CVZZ+iQpRYv5XxKpYNvUt3QPbgdUymfCwVvFrh
yQ1WJP6ZYjvLLR2dnBDX+Tlm5kqZZoVf9PR+wC4NB3Rb9W13QZZ6ESnJJyJn4G7b
C0YgGM82CvfejwdGUUhVO9XXizyfWz+szOkQMpARzccXgB7QLYBxqOz5eBvKUiMQ
4ixa2NZ+p4G22h1bXxHHkKA6wcYM+g3Rl/k6ftdhjaZjR4Do62HqAVR/TSoxbR5q
3dskTx4SEJCjXDq0mYj2sg7BejvLa08JN1KL0nYWlhQi3Xia2Lyti8iMsd3Q7O1c
Drejf0IhGKLGBt0N8KMTclM4RHp2G5jYwEUxzg+4fNueIOmscv5CTk6h4/kjD1Bh
QRRD+g3u3fA3uPichOl5xeIwUeE/XyoNj3DxxQwYn8RQpsWt3LlM4Uve/s64pIc5
IqBqn4JjdzkD0Hij39BOxenEts3zVVylEeVx+s4jIZ+9pProsu5fM/PKWXgh25Jm
e95v9ca84q+Uulps4KZf+PyxYjfHIrxPsgW63TwFuE13ObK6y6nlzO5qX4haUU8P
LYPF/q2ZLgfTbWufalqbETo18SxJMYn4vAhM8Wcqp+YFd64bnJmIqbifHaSOKseJ
j98Ecc61FsFuIEim4tAfkSTHM3avFMvEnpj+AY8k0tAUHae7U8BXGZVdIJ9NunCE
WmwzzKvB5+1ndInHFdG6yDKThkJlSyxYhSQQj7rou8ygMPsoYoymCArf1BdR9RB+
Ecg1lMd9hClMksA1PGtrpktWB5d3o0AXhXDQeYojFwI6zowlFKCKZSD4JbMV9+do
hH7fNEnzto3T0T9Jq+qqEm/3t85XV6N9pl+i0dyH8cGfHsXUNwdTu8osOkUqJYFF
/exa0FFqIiTEVqGUFpVtyYneTHtCY5ekJOCElu5X7aL/XIplQm8SwmwJOhko8yXU
GQXiUwLHw9/kuvuh1b4ZBvUBqtsW0vQSRhYesEhoosSLFOxg/kQiV1o+jT+E3ont
7xJxB+JndZOtp3nEooFVjrPfPzA6qOqynNn7wDaTxAWgwiasp5qzoSqbX0Fy4vcj
C6iPnMDYA3QAubMxkECXE+quvUDMfZvxPpzaUN+fwjeQ+EYlN6Y25GZJ9HaC41PQ
C0bQv48JrY2+GmppVvXmfcHRr9ZQdwIMulTWOkHuLuf1VXplIsrWjdWy+j1sfMye
siyvjVltz4rDmpJJdM1eovEFytp+Z9H8sXitIdaqicDowo5fcGDupRPxvN8nRP2O
nD1snQqHCwX1guLY/Sx8Ap4qnET21tfZlKt5gy+UiFKyPqjBSA0X5AgHu33oxJDc
QJXB4jTcauLaJnnqtXbtKoilILgfrJ3YVYQP0Q37QwBhUxCZuNddZlm8xKu2p2Ho
ydnn/c5Y0kza70NZVajiICg4HM6HoF1GSr92qYtDSKaxxSxhKObue+YHeKLZzIiR
lle11ey4pATLFp9faYeBUQ75NPp7fixkiTnMeqGdFuxNT49nfRqh16Z6EebE1hzd
h63fuisDTBKPOiY7Rn8O/kRQe1Jkda7tH6+bylPQcAU20ta31v3u02aPrYcjZLyl
JZsr7W3UTFmJDAT6PYCOLzByEtINeDS//S6eTiuNjnm7l6Pgll4oXuyv6fHAnrsu
pJPv+1W8EIpEgBMKnOQF2RrJGJLcjQiq81eUCQ08T9J6jc9yvbMmMYRvlSuUoIC1
wq+5Pvpdv3eoUq5GqUj7UyUw5P+W7VE9/prOAJ1cxpp1bYKowoBCFicytR5QkFsh
xcUJliP+GDa/8KPd3C1LBHZfFRBGEbkkPB+vR+yv7dgdyOKSOq/jhzRok75XGC7Z
4B+GqXssfcbfJMDOypE7McoBM/eTzOq6/ooxKFRhyUWIwBl4ChMWn8Jzv67LllAh
DpWtek7Nlq0cYdlq+jkqQ8VDHMJRlIeKfpT4D9SnJwXQbyPprGh/obhkdYgXWUTE
4+z3anAAFx7g9oSYXFLI9Ih7pwuHGXmIdCRQ/HLHQmQbHWsN82y+K+TLO4YiS0IC
/ZxFCLjsA+/hnDcIAau53Xb7NhQHj3/P/TMNrKKwUPNNYg2Ld5P9jkQrm0wsCJlJ
OiWD8keu1i6S5oLDiz9VIROKmxEn25zyPbAp51OCV5L6rN01hmMc/QAeY0aBodp2
waV8J9O0dtm80FzZS3C8ioM8b6KHzVTfM2g4osngyR2oTsBabX1925Jg83HklfNB
FcjrgON3g+IZikQ7lzlnsoda2rJhdXZ1KvE1prN5vrDc3crhTODxvf7W40YHEVpK
1EUZCbNi8pZI9b/DyYxRMN46D6Bxgu5n5GwbvvDTmJipfm5ZBIp0oPNS09Xml2YO
isyqU9WkM1c0s6PatCQsviYLbvAwVQRyVKCA+U+pjrcugsbZWd/pwHUuQr/IdPQw
FNmI0clFn6OnBMS9X7IbJGviVUo0dBS9iLTploz96fcXn/te435miKg7q8LuBx+d
DMJTLkl2jRNomspXY5TvZ8WSZC1bi1MtWLi9DfnMKGPoNk/vyKz5RvEDbVzqV/gy
PrDU4vrzb4gLwuJxTmEZo2yK3qnuFAqNgVt4Lp5/ibtV+67HS3+q/uDmA4+B08h8
T7yubeMYAIwUt4ERZ6HjNhvwQ37IeEMEYstE1nZFr1z5Ooeyy896Nvdsyv1oWP9H
BS0+cL58/vahH7NYvnJ3cddZFzVy2o3MUwLdIeFI+X5t+rTELZVUvVekpEhslxi1
TP++5kbUFX986EsrANDNN1hsmNrrqKifyqLDHeYgfXzCWe+iH/jxdJxrOWLNYNbM
3xGe888mHrucOsG70n61tqfWZ7G6WcI6XSqVFER8oyumAQ6k4OwIag+fmNPhAI9p
WlRXleJOHnB1nBzVgkvqf8yxFweDDFNXlZr09g6E77iHMCj+DNMWcxKgqbstg+6Q
8loIDxaJ+2Ima0YAl8foayteuvAiYBq5hJDGG+eReW/tQ4eduqsF93BW35u3icVk
OmL+LwI57tC/Ll9bclW94t4QkHJaGPH9C2Dc6maNNrqqUMjSS9Q/ychrNSFHj20H
fDadNrA8xN/1YO4JPoKdbpk7MBP6SoXK5A96X8Xn6R/EigrAc3GZpgalzWnJTQPj
Lcek9K6earudGlaagx6dR9kBrWn+HzfhuT9TteiY+bfBp04Z0NKFo7ZS6qyAfpke
1n0Uad1IAVGwFFDjkq2iZNK+ECN+usFNhvtaC80o3sqUOiKrCerUGRbPwvsLr2eg
u2CsuLYLoypBMzYpPezw5sz4x0Di6Am8CI65pxhcLT5nzp1V94p3znFXFHY3NClc
BjeIipSgnQjvRjpru+sLC3+DW/REdA10ZXXpeCh9JiFO5i1Rwa83f17/Z/srSmD+
aGyrrFMim68I762knsCsUm7VzoVNsq1FC/DT426DWMT/xSHMbeThO2IoTDO1DygO
FxqipcIMRM5P/vMRRLx2Czdl4CbxQzXdZk6XVGoZ7iIkY1o/vgbeTbwScliZ+5ti
pZNANyj8YavXYKksUC2vyy9HLkl9Ua4c0k/eCCn3GcJX5gCivUV5bJhlPXWiQdDc
nxrbZJd6qJ4OrUlS+P0G7zEH3GO6XG/8tupEeDreQbEd1g91C7YjwFcHzGfzAZhv
Ub1GtdlnQ5W7il14v/PtZZKTCn0sp33WRIpLU8vs1Y6V/jHik0IGvUK08nCrd5P3
yno1BnySRZ1zkt/ZzuGULlCanBchOisk5tHquWcwLNry5YSp1RykFUSNzyT576Xq
5ZrYoFNwHFEjOTG7zkaQOkdE5aSuNloihNLoPPljqHorOujMELK5C+Tk+dmz17gl
ptS9yLyjiywUfE4pUMjQaaqHF3cWz35CXQnC9i4SrvvtaairYGphXvSi7b1fvXyd
QPcWlJ+YKM+p1fC+KLlpvdEifOfCh9LrYcN0iPjW6TMznWg7QsvjbFJXv1fZNB2t
2du0FfBrNDmf+xNTzz0WuHAhzAiqhJP1yre/hdTp7Mmd+CbXa+rSh6U/4Istxh2h
QhOiuIBWp6FHb6ptJzlZHy0p96pr91xxqUbylX0E7g6BiCXu7wVMSj2hP9u2fJpG
zdluWRkA23v01V5NLglXkLjsBDtVZp3orDnWR+tCNSk/a7Bczun5YJHwR3d20j9T
jPYZDvQ0LEeWuS0GW9Ap7nlY1zKrUGjus4+XKwasYjaiwCa5VOdzh4F4WE+tTGZ4
xVlEJpSIhmCAG9V0Cje7Gs+/zLVYNz49AxR5t+ebS9vJ1bJeaFd8iBCLEl7bgm50
Pkzh7i8rzDoOhe1wWEEg9EQ3PfpNXuohtwCxFm0xcAGn3VojeXY9Xe4F3Ek/ynEz
xl3TI2qNLxPkaKxLZkXPQubhcyEiSCrLB4jIIbdTYZCQ2D0OsGuPiI13l0g/dfsM
HO8CfTv4tBM9BaTv/2hPkFT87MqiPgy/AXx6jYs3sXxJECbL/A95B2w75p9av9c5
vlki0JkohQev2JrQckGYkSB+muBuKwWPkk16i2CjCrNXqKTmJAK77ObCbLnDnbCQ
W5Zf5772ZmzMMA2jxjhRhAoTlH+IQC5D+YJhWNRVr8FpYKI3kDDd79Yxw1tWtslQ
gNml2DBH5VAchYe9vBYJXnsXiQLHKdv5N4Srbnk8eu/imlmq/3lGG87+i99xKTL/
jyf8SdshoextiOyqNiSepdwL+/MWADar7SNi/YByuG9TgoeaLyvQs8iPXLiNdLdV
/NQgOjZ4NsS85GJY/FTw771zvnVs+pOw51XkCINGtvd50m+kZSxAOJWUs3QVmJSY
8ZgT7DnKKZrPrit7R7NHVBc0UKp3suKMB/JdpC5OoyH0SkSMZeYnTCkfGPr7cKOn
CkbZqLXmzsY2P51W9tQa0xDK24URXpOm5Z3DjZHI8AJ+fXd7Fe0YOMyaPHzZx94K
ngrZWcGEYyYaExc23ZsOIeSVIRfyDY5rF/BZ/dQfp9UlcDvcIqtA2wVcSPnQEBvh
/3oxNbhIHb5/uQPHg8LoKoj1RLrf27qVr4GHYg4cp2sTfWt+PNlzluMdZoombW/K
Lr69wtR6cn4xdHM5OU38OXMtxWBmxax/kbw8qyIE+EDgIS+IZXQcfWKb3XhTEd03
dtnI1EjYH45ISd4QancZPl9rCzMAjCPQwiyYao7fCZm9HCDDalHAOoWVrDIGjMQz
M1hyN7XzAqjBFPW9b9g3chYeMUgLv369oF9IDp345l+91/37oMNED3th6Ev1hl6E
h+kDT3Ar4OgV88l6wmcIZQAKTRAyFDk5vFOsXoE9WmcLMZvLK0KvB/siPi7oBzOl
iABVuYdJjuU71ErAZki0sjvg1XxQQwu8+OdrTEEDPJ+Pipe/Tt6QKBvP222VZVym
YL7X9vky8QsI9FuA1Qf/OzPgn4TpTR9EvbkI7jM1vq491FDHpotm2ambWJ1VSVwp
YyMG2bXctPoIWLacHKtG1CNiv/5LOUK5gq/46BoSr8/wTXjpYJftm+ctYcpptoQL
YdOAWEmQQ7jdsL7viFdMQdjLRa2Vu7aZLlu2XE74N4/R9JfCWGH4jHK/3aL5xwjK
L5Is96/H5PBbS6QB7+CYVdG/vhUMLFiijEkMmXIfqGIy32GTaZ4xQ4lt9sZ5i/go
9KovjKpm6N34JIVddyn9ZUqY9OkAz1QWadLlJTkvVFJXcdemx5JYoL6CTdMR7ekB
8RkVkaYliQT7Pu4rFzbf5s5+pAWIosdTvEYSsYK19IMPI1Q61IpmfgGpIT8lJUkN
joGscqn+ooA9BwNGrWMA8sT540yl4JHkHPbuft2VKjAppu8W2VwrIR4hxs9RtcmS
eD6lP5p9+2D2IvWc3txpwSL2HxFFA2jeMHLTc6vhyE/FsCQqdooFZCXmEy95zlRq
xJphkM7iq0HrrgV9nkPQDMoZVpO/Eyj63m4pAx8ijxg5irAThlOh2qONy8HmEf3y
FqH+2Xw52vubpV0fyuF9sugzQnoaPZ9FsoyXvVN12+RjtgFH9YUgMTqwr8nLZGS3
3JSPxKpAFM1URJej8jiGq1Wo0fRmZ3OGaVRjYy8clDpUDNYqH9ifJUd54lvGA11x
5oikUCPnbcrd9+RSZvS11DJ5UTkFHbKceBXz5xB2gDLtwimJSx7ZoI2mLDZaMTj2
9EQiTjztfzc72ya50NDzx4M4Nj0v0ujFv75xOXKqiQOOWSXGx8oi6M3CCinvFJMG
lV0rLJy3R8OgBs8Dmm05MkTZAoSYVUVz95A7aKyH2fuPQ3XG6qu+HzCwuh8bw/mb
XDCIK8UwyXvJOPGQ2ycVue0mkz59BNfr3H0QNWI+UnoV252M/gR6PjMwNe/3CKal
FBXmSzH6AOT6DRqX6LPicg0clyU4JYBthuF97OHwMxj7RzBTCAbWISBOk1yZSdCC
SOfuu555EEFCzcB3z8MQtyCqyJUAuH1G89a8IgnxAWwJC4fqzg4tqSqUddwSIjx6
wLek2cz1I6D/GckNGJ89APIpyXw+9k0L5jnJWvtZ1AYZHF9W8HwskKFAZXk+uPXe
SjU3UZLr3zSaVxezysNM/lXli0kdguH1iLQcCfex0S9RR591Hl+XEQs3UHC+b1r9
XGACcU6rNkJR405Mx/+QBI7m0Of0Je6nlNC6VrnYOMH2hz46u9FIMeUKaqJIUJLa
8RD9Ndc/iExGcLfID8bcGC80I+riwPovxu/CpJjHp1gksyr3SiV8hqF3RTOPvZmo
ZvApXz3UrauU5EmD56a0pFmU6wxNrStg8nuPzu091dtF5zdZwRXSAAgMz1eh0nF/
IjmXptntTR4GO98fc3a1P+1dWKsO1SV4A2BliRrMzfJki30gUHVamJ17V1owI0H8
qS98EVWHPu/LToc6354EWl61cPF88RzjIQfSKUrNc41YCpo8ZhvgG8g7QufSUvNc
GcY9/fe/I1L5ToWniw8PtsEn8BzR4iD2G754HmSM5KP+Yfx3nTpdZ+4rxnhn2IXw
ig0fm6oVJeZoSVvuajeSdH8X2hQ/Oo5v3Yq8TSxHC32oma1OpzwksW5gkbAvv3ZG
Rar5lkCbzVLCFLT6/SfYwhhIvjNTTPiXh7Nx/PuGpIX7UdE+9ZbhmORhkHtQXSI0
sP88pDmZVhD1Zxfe52KV5lQ6c7iMsc9rWrp7Sconr51H9kDikCmLNVMrEX2QspLP
Nnzg2n8YteAq88KrJZF4YvrF6HdYwIvi2SeCRGbEUZ0OG8d9NrkJzdxGjqd0lWId
64xqQJPk0N/m11iOC6FO0SlrQOKnmFLjcYckF67coGfEgO7xoKNg/8z5xNpUWkPL
d9qySm+oQ7cCJ8svI30Tkuz0XhOpXtAZUbNjhy5zLHAslDH4GBGIOsDwtD3tvmRk
VEualxPwTD9NgMChYOEHsOJSndbSXWS4RHtqdexgrdlCt92AZsTdn4GLS4PKdo42
J0CCNMF5ng6z9PEc4a+ySxVKWx2iCtu88MspcfHaT9VFCZRVwx4LUQOUSDRVFsle
qrRKFOz7k9UkbkUpAuNnXhEohTuSNrFkplvB3p9mWkZ5xmPSTkeHSZBXPZJXehiP
/VD4ZGJK81bdPifa/TDmNCFbKdZ6zhY7WRg6o0FbpOCjQELikC82mQG/OUcrBG2L
Gyq85YkIuisdbPphaWeu20PrIO3klw6wRQt10c+nO+Wu0t7c32cd8SHZKoplABGT
CHdqQeEv3VhfjEHSvxpYCIgu3nGQIhwFBehfL+MjylFCDkMyFDq5fzrXlYiQMWyE
XdJ2Wt8KEvupTnRUqA4/LfXygc+jIa1DJOcBwN5twRjKeqt7PF3eBPfvdT3e6zT+
r1H/uUCmA0zWFn7uyxPQUbp5PJqAwoaTJNMx7jh9kW3WvhMIw5zf+/HvKagmGFxC
mDbxWANGDbTyn6tee0ij7pONKvkBDaRlWyEc1CqqGY7OzLy7WYyixcpK1IRT9Eit
A1ewJbc+9h9DqQhyo1z7b2KCzF3LRjeMpmHD9gLKzXZQAdakUyakAYWwQkuo5MaY
qQNRMvukimGGgsSrcpFiDNIrPyDddhKPfuyoSO9UQlTJzVLPiU8jwLt+fr7ibsNn
49wdxLOQq7P0+L25Xj02XZjrc2jlALzAKMAEK5FZe3UNZ0XHcsI4yWYB50QpX0z+
sy5LJXKHa6mZV1zkK10ip+9/seWK5xpChQzVc/HVvsCVrWKp7ugcYEr3o+xjHHil
EhF39jPE4lPmAYboprdmJ2FPYLHH2h/YoQvlmEo7Gnl5zK7QjV2zmZtHN93hiWvD
WfiFNCr6LRREFyCGQy0LGYu8ukLWu3zQoFhcXDBfKo/G9r56IAeX+ONL0rkTidoO
8lqmK5ujBMToUPWaLymhfhPu875TkphTFHzTqciDP+Djs/+etGUwIy1PQIISuqdk
sQbFAd50X2WEYrJiZfxexqrENyjUbaNmeOSpg+ADEB5wuoQYwteF9DWJwHym51Hq
xOPsOyE111S7G5XSNeI4L3Bi0rTjcZugl5ywBmed2IzYs1NkmJrB5XfUA6A+Vgwy
qAaULtzEPjUAicCzmCryWr/p9Vj9gVrBv03YOTk3pxiOlcNonoF9X2cgNas17T35
fT2VJA+afhyBM+lm6nIuEJy8tDNBgXT9F1AVqdhHVCnQ8LpNiXODrCtXm4LVCiW7
8BKFDmXZJ5wk6mR8HLNiseucCGmZWHVW2HxzCy0+9/E=
`protect END_PROTECTED
