`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WCoDltdOEjiAJ5PV7n4Fs1KO2OrOYdYm/FSuZK+KYdkXaI6l+dQ/hvfJ7D+egzXc
LJ2M0RpQIrQxQwJvPOALovW1SkxwwGrF6Ks2ZbNTw8VidzhTIkvL+O5SuY+VGxpw
SqXvtHW79OpO2lZspMergGyHl66BSR6qUNZjkfeTcjy+/ZQj1pYFV5EWXIa+A70N
qMa3O+HTqlK572IQda5xd67dpZesHIW55vYLbuWddypnIWx2hz56sQgSM7VGw0JM
8aUOjmUg/gaYZO51tSDk2viwYBknWyBreqp1UOyTH9rZw3XqG/4ImM2t6XQRXwGG
doiZgqG9u4tMNDXFViMecY5UbPn4vHXX/FhyqdUx9upMymuPZXAFGpXiXzIiOgOH
oG7St+kR9u9yLB/J2Y7E9eNQlJS8vMnydx/92Mo5Z6SyVfI1ClNFy055nyDYv8vV
`protect END_PROTECTED
