`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FLXMHaK+B9ECEfA7fGApdI2DLqldGnlxhLkZOQmu2l0H+1Of/W/SMFMNzcx7AeLa
9szmuFjN2KbaMyvhhLh/Rv4bURma01a6dmPAkP9epyl+Gwt/vZKSi9XcPNL5ewun
G3Kkg8Xk24V4rgJcmhlblMvZGuAW6WTkaaatkW97ADYNrTAmETUdZwMrx7O8r4Wu
747d9kxXeBg8l82YCXU1lucf1a+kJB4JpRhDKPlOPQpd0u9R4RsXYU1XCqjbEGeL
WBGyNWAugHObr5BIvbdagiTHsSdG80mWp9Z+vkGaOspT1mFTHs3Vo7tJ74bqLcbl
8fzYiINHUUu8l2YaJ+nvgZDVM5cGy8Ckxpb296KlGQeYB54EW/3FzokDXW3xEOpa
ihmuIctWIR5P2iJZxAc6zYH0YiovO4UrVubCAszg/9aRhkrFyPVVmLXIocjudV1u
Ezjsqkm6Qe1jkqjxdyjjubOx+ePKkuu0qSaY9Ffv5Bfsip6L6WeuZOV+C4l0taEZ
acxxAqkzved85ZRrSrropndnT74bV0cgesXzf6JpMVptdmS4dlj2pGM/ivrvG9kB
RlHBdvkyh/zVZNXzAvAiPTlh62jI3xsU1Tfg6cDxyremLLjYDRWvIDngYU3bXrsD
vMiZbK/c5RzP45H55vVIczSyWw5T5TAiJRzQVBYkb5fzraCS7p+ojXr7r7xkhdx2
`protect END_PROTECTED
