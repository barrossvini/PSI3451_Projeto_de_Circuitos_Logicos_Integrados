`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kwO5f7ckfUHejwOeYhwQD6NYcgxAY7oVVj/BhQV4eqDh9S0VvLpYKz9fmx6RqI8B
m6juBxMflzzR8hhCIEMaHuovrOY7SRMmusRGPnf7X4JGOVvhLnfpbe3vlQYBPU3t
NGUcm2Us7wpXUJNVWLN+Fh4vXc0vy4heEpr9+G63+1TvyJs75hhdLV8Ele5XPp3u
FXbiNA+XPnwYfeZRm3Z1qiM5ehz0gjl9z6lNxXFLgOAQILV5dcWmHKw8UhZUweG2
TaKCI2UlCtIfPZhHuyPjiqyUSTcwGEWS+7dCDwrm45kRCwNtNCifN2Ig/cGw/prC
yAIYldqHjPW88C7ip/3HPUCSshiVu6vEAbBGwl5e4qhWZ8UTkZQ8ixzDetZiBBcY
Laz9sOV2IVCe9w8ATzs9qGHguiTGC4/wf14dlsOJiLXI5VoiPDGffGnjJyeZoc5T
/rvjLRa/KYXqIl9ZUYNbP8xjx/90A5OyjouWupGdaavjBwVdnWHURKsigpDiWWN5
QxbL0t6xCtke7PfhH9q+l31LM1uJGVJYTzxMEip5lRXEYJdNDtvTsH8GlaKJ8pPU
p42wBKr0GceDxMQjRVuscsXir/Fk42W0lHWLQQhdx/DEziEqqZP0YQ8+v9HvpsPQ
BT+e0iMejKMnJdNkqNxKNKyiz9oT7mwwOau0TUwTk4LCo+k7Smsdpg9zTpCqp/El
t8aFJCodp6F/pRnKicdNCOf/7+i9YmGEU/RTAjoQRwqlTjZDWCMDLR5AirMtoYm1
wTXv+Xe9qfi7EBlIjfTrJPIMjaXMBJImw9ATkLVLlaOda/YsFGyL4cNyDxtFdx2H
dV4KVkck1W5VgvgUOfaLuMJuDuaoDDaQk74SnCOLVmdaoPm13p7fyY0LfID7xPUL
10S0Q/E30GRLVSU0Z9U981IyjcfzUIRUSXuxbAedoQlImKdtj87dsftQjPfKjxM6
Si7S1cIhccMIirtk9oi9QUj9haxnlGA3TnohgCv98Rm/b4+DphX6WZN3zKAZ/2rT
b186vrOVPNYd/Ry7HNPI9Q==
`protect END_PROTECTED
