`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wLhOEpBvfNC1M1ljWutxuRRRuPPX+kHN0kyTCdMK4nECCVJy7Szf05i1p9paC/Xx
v0ku3zGAKxwKrLQBjCffgrEzKcMPC5FuWCbJD0NamdeccMHVOURh99tdq9HEQYU6
03pOX2CIzteV6E99Zjcq4sJid9+VqaVAsFXyuiltrF5bdObKCrHXLWcJw98DLdOD
6RT9vV7p4qAnEDDZOkEUkfDcASIa4kEW///XUF2jMIuh6HmWVNsMTymJMKJfBvmU
UvQw15eUGc7FZHOuOiu8vP+TI/JKs/7Xqkp7wkCRiUgFjcioDpghV1eXInk+ex4o
9gcZZeyeGvDoXSFUJH5DCVXT5/2suL5WxC9y4gEa/dKSvpaAGdO7NpholeDRzR0t
bDn5pdD+/ZleMqMDqg6eR4kFr9Jg+ZDRekeSOhXCZ2oXOvJMVFMkNiqXCdcmI8Tp
wNSPVejDDm5EiM1CencvLw+TZualemgVW9GG0Ro2Yhfmp6yi7ZLTOMf2jGnSvxLB
/Qeq90E9mSOknTUscbfI0KjtcymZgIfdwVA3YdpfHegXoJ3prZMUYGXN4MzFr2JP
apudn9r8eaDo/HAyHHq0hGp8os60OwXpDq84T4xxwfV+MAfVayX8CHaGROgBnngj
tGYlqA+rboVZ0qKU6ixpcRtqeehY2qf2S0C8pJZzTqYys3t4P/Nl6zZ+IrEK4WEM
tfN0T1xSVWm5E2L+uT0DUQEfTV+GSc3ugHauFV0JTowVyxKFzhtRrf4U+CzaNoBz
ZuVU6g3szkNnjv42PooYPcCes7qcDqdWITCLV46bzBX6cOphUKqTpf/i/ezZYju1
j3cMGSwTwhgl7888ESo9dX1bolL+HSAqbBzqBZDSOm8zYR6oHTx1z/MwPOF9iy9/
hspiibKtDVL/Onjky6sb4xpLnQmuUj8nD5j6ybwBbjcN/F6hLbubt1YyiTsmPbUO
0nUZ8WYA42sk1m/ipdLk1K2zFfHNleb/5cc8RMRUJF3VLsX56uGJGdT6Gks0WBOb
6zMqp24YEHA5UuZRWU6+8Lxc4kHr07ILvet/Eyjjf/dz87UT1D+MatSXM/xL+t6Q
vhaptMmpge07Y3p9C5aRBeLwywgzE6biB6CPR5pyao0MnKuHlc9sDTU8lR3GqmSB
kHBVJYHN/JYzkSbbQWjxJOShKpz6fbQEkhkJSuAfAkqnEON6ABfmdBIP7goE9unr
Z68HaIamttzb5wgxZiZN9rs8u1qVUFfQiJI3sRS0+rjPCd1j00ksV1Spp0kNEHIb
Jtk10nzeeSxRsVPL41f4XdFs2madWauvDslQtrrBsESNzGaYbVcLaLugKC5LFfwk
JK1bh0hNxCtl0sYyFmYEGBF2NljdthThAxEay+QHt4NQRIt/wRv3dJl9ezszXTdw
HPMGzJy5mo6jvtO752N6xqIo+FTauiCnjGyMJFu/Y7jU5zp0mseo9Dpv91IKeKPO
Pwgrmw0luldsL/vKo1WGwahYUsc7UAQrLH0+Yq7L9qFfy2IOWNLTU0XL9QnwfgIG
Xn5itPhBjbCdod9jARkrHReaLhKjKA7toDdlW5vxWZtV1R34Kmdt7H/wB9zG7mAx
pn+kMKUeK56BlaQp4bal71U9wR8aN/gMnJMVXsH99RqzTKVfWWN73wa6v+iDR1wq
q+5KXW1hJbsoT+mEqCkBmMkn1b+MU4r3i3S6qeKJtGqIAOQ4ZLk+YfYu5AeyGgvf
GpmGanQC+fLLCi0bCAUzka9EOdx/TdZwrrsi7GJH7UjnRj1rOWjC1kbrJhN+gr2D
lAAd2S9BKDvgUNB2PWm3Knav5B+G2IaJS8IuMe50ScpNvhR6VxV+ua/4VV0HLFV5
1CJXLOlXmAzK2Gvy4jK1FFOqAxhJNIVuPl2F0CRtlscxmgUkFy9AYVRs6Xkk//at
Q7rxTCoCOfFwt2IxsujVtZDVDeoNX8j814Ua3gtyNi6y3xEFLf6JYr6uoegFXSL7
s0DZExkwAT5rIFpd6lcLMKPdxFTqAiYhekC32eBAtXuvAZABrX2/Qel6ck/CBlDp
BtCCurKy/dmTF1T0QsqXy2rpmNjjNXpKHBzRVuJOXXqeURsqxuegWM1fXHeJ6e/L
Dcdhkxn7MIUjtKtJYKKr9eHhkCf2u2Wk9XXh4hlBPYROr6D9qcuDyMEFgB9119n5
FGB66R9g79hHYEFGUxa0hS4gZOHCJA7vGLUlUdZ0VrDCY1K/ZXGcKxKu784zwbjF
UIDJ+cXrypXQkzIVt7lprDzzeWErjP9Nifv9JHm+y3n0k1ZZoGWV0vFI32TOvz4j
nZhhuWnluCYd/FoFd8anLM5JPjFDEEC0b+DfZyubDDc6vSGhTxZhziiXSCVcRW5l
Q1lsLDkUzUx4aOjQ3Wc4nzPntMhfiwUDJHQbCyuZS2lt5bdY2CIxUz0lLhQAc5mr
pZ2KCFeK4Be/D4QI19KDz/cfPMOtYMiS/KXz9KH6HzMgXEh7GLRQ9Fdj7H43jdXx
FWTrOnejgB5uVkF4gsTw9UN3DWwIbxhvE/blruX9ej9wSBukWjm23zK/OvdBzyDh
oMLQqi0HSImsSx7Sv26PK6Iq5zMMTFsRLEXsHvAGlE9xRzvgHnGxthFNVx0qoVJo
ZXgdyoxcaAzKx/zfiqXqVSB0TVQJ7EqqgNRBAbkr/+EJeB9G7DxHDC6ZIm9zUIhR
hKQ/AREJlxH9DtJjA897IqPi5305NuhxZymKZgCOxeCPA+7LMouPpRxqGimRxAjg
VwG6cn5wvoHnErRSqR01ch+rEfT4UTJmDaJAMeBo7WEskAITVGiq274DbRU04INm
4lUliqgjlQLLW9SEo81JccWQBFeVL/ywoqOhksoZ4cBDM19QKzVZNXTSYZTZMKri
6ZWQsFrUhpEjONcm62d60h9e5AsbQSXd98CRwZZu2J8p2B8pGqp7t9qKWUjSK9gF
BGcy0ixTSWf9Jabvcd5aL4asnDmtUVrl1wpHLmiD7XVjr0KDrEwxTJ2blubbC5Eh
xN6tppn5Su4y9S/2VLHiixau5ranZ1AFGUInwCuObfTXgIfhljUiLc3JUv7QFN83
uGNx6zq+ZxkxWY2uQFFoO2slOKP5Sft8bHefTqzx9DPmLYiWrfnoSMjDgYkMVamG
mRhdYN1OU8yE70eftXbFKDeOUY87AE8UWQjQHiTeYlGsWI1jzkSNiPH/Mdplcn2y
cLH74JtIgTayqYem0oVpwtTWToo6Av5m6Rt92YX9ziCXXExybrGXhvItLH/En+SZ
8caYY77/letWFjpEa71ywTE8ghHEzkDSekDVFR7DUhmWu5xbIkpYJ44/srKklXM0
/9NX9OqOhJkCc0tPNLU8hFvHq3dhXK7OpqhP9jm2nlsvouRZaplVZh1vH3+mvFz8
AWcolk6oNnfSdsunnxRLXWl6EBX2PpkqszkKWZBdg4W4ikzLfcjMUAGe6TLU3wEI
35BnVJ62eSYuItiW7zrV1vw48/EgJzP/EalAG2hefUtwOThTFbrhKz6mQhx68fTT
MG2mpZ0Wc8/YJ+Mi5awAsQDNjY8AmcaenW5NF6AHOtWx7JoN0Ga1YkPjNZTr30Wu
yrOXKswc6lYlsOeUohA7fqZ95uAigg1Obgp4BRJBLXU0CYEw77BValaHzl6BF+GI
8z5Q8YxqWsIqK+/kDiGDfWpYu0K+LbEyY06iZSDWyooN3Iy9s1uK7JpPfjwF5ANj
BJtjOdb6l+tK0T4VVK6TZOhZ8zQVheOEcpSZ4qhzWkwrjatn0X00m8Max9hOduyL
YU00RL08miYWQ9ixk16KMMSAJUCTBixqBcWZBxCqCEXwwu8WxuVbi9sNblifsMnt
vkTK2p5BDLJrun1YTJCCbQsA6rjZniFUg8pflYg6GRqXtBYRD1aQ+ZOGeryyJZbP
JAlZWdS4MrtZRpQowDIzBsan3Obtbzd8sycwMf6C8ZmP0atDtbfamFcR+x39dL1C
gIKisvX74LD0aWG8B1CRN7VtwMpJiYNfX/4Ok61XKKj5oOx/O1EWj6U6v9J94JuI
DqxWdB6Zww43moRuPT65wbdVRurdVQW5TCPlzwaa9JzK1+usphQpdmvnfidztJSY
M/JVVgiyRq6lQ9JEnJq4OmlPD3UaSgSDGdp6p4bt0Saks5hYAo2tMnuR50bhkfUQ
AfJU+B1Nwch6vzuQ/JMjxPab01WflvQcpbUdzB/8vt9mZ5CIcKW0PVrqld8ehCX/
VjQVjElce6bowtA5nVZirRrlwyd9Gj8Utx+N9uhIQc6hGNuxRprKkq7nSK0961km
hsN0hj2hUzuqrXrsB28Zltc1iqhvCI0FXdXPlHbLvIOJKVP2p/K6I4gaqLbwyzkF
iWdqYTi2BxxDj+hq1BW+WpZIVf1/nI3Hocm1/S64gLMYkhordcxFny/5VnY8KwEZ
b9kHstz8j/4Z9nmDWH+aOP7UtAmgYUMHTTLY/DIWBlFbuK2uuBfCdAyNtOZUSoIg
6Vshci9P8muDUBleNabqeIjL7oQSaGT/2ofn2dIMepnhD8YdDT4Wq148yVd/arvg
5eALgmNq2kpg59SAx7TjywijZmCR8I/Ko7guW9NfftS5gauDhwuhW0qH7Wrtc9ew
smeboNW0PpdtVkKYw4g+6uF+bWEACFJHl4rOOl13mxuBYdGgKEY5ylHkJXLWGq1F
kGb6WMxuQkYMEPDJLHme2chTGzvZJaeJrRpTibpz5dQ6tZtmZvSBKDTlgu/zcYiV
Xb6gXUppGOyocmrO/hkRp2kknrruFmb8lXaF+XScRTN3aUgbZOdsuSyJ3ou1twFq
ZyX/qGZsiMskZcYz1To8IHOBQpK0Ezb62JbesO5yqZr/wxKSiHf69x9UoXS6Girs
EHTKEvoDOfG8pJVmT6IDqAp+v4+47Mwph1ZHkYxU7UyJiyMldwensow7Abl+QLjB
AGydrostupMOvL4xIuLYqwWF+koAEPleAXzH7FipG1C1bhdo7JH9+Svft2l5xb5m
wqXq5IRXeeXtZofaMYdZEtHsgoYGvjEyyP24E1AGG7/EdracnxEGnBlp3SeRP4RS
UElg86kyOSaKrH8i8B9uxaX0voA5+dAAq/qDt9m3L2mpmUlyoXBEnwH9jSU8GZ2L
iH7hnbTT61g3XCYJIuYsvkoSBJoWP3FWY6A5XsvJjXaJPNn/hMOrc6wPdtI3ORPv
p1v0dR9iq2NYJZERFQtXKaMeie4l0f6jRNoSa76pzmx7tdyH3CQb/DtamGPHgYD8
e6J60m88BYgjZKrYC4dp9vY4nJADN2eS+mnUw5/EHmyu+1pFgldXMTDtFYnj3s5U
V1LLoSqVjnOPn9P6gIHD3T70oQraRwRH4ewnS+crG8Q2HECsSDHfV7Hg+VTNwmsk
s8nMzVhVQpgNP0fuhYheQKQ8Zume1rYvQs8Zqk7OMqf9wCukwGXKyBa7gUhxk/3m
hDmoO4XoDpiPUjZPXJbH/kb6ae4UThrQY4cTvBcy+ztJHen4t1HJ7GVNPh3zjMmx
19qCdMEfOVH6De3rwO/rgQquR0ZZp5YgSuUlF5wlZGl5gDDZcndbl1AL+LXLGHrL
CQiVwHI+eGaVZ1lchdK8mcQiMxZAmMDJUywu9b9Zu4FWaEZoF+r5qudDmEpYxVMq
FYyHLbg+Z260gCtnGglReCIP8A846Hd6OG2cGxGgnQ5hOz2insb9Atj1KPLUkrMP
EgCO0dgjIwd5WidR0iYnL+gv4YzcGUa7FyYoN57YvT4Mh9k6FGg/6LLM02FsubGe
0oMxXXF7SGIn3pMKl8WdOuHjBzEcGsOo4pXJc4/Yfdjak7FJ1zkxLSRQCe9HEGa8
DJNLXye1NDTa4ubndPaQvl/t3mIhg8MUWDentSAwe7v1H+ybZ3nJ10ErEz5dCrSC
nNSuvqOZYJQLRXV9bM2+HWqxho7mK0fLwZC5ZnHRCBRVhPSm6qk5lk2M+CCRUGgH
SGl1SeKyA217+XAS501XmusanJ3a4EW6tgQquI6wH1ukX+LxkrLPmgvZ8jWLHbp7
qHJGqZRTMtqvrm93acuZoZrnH6Chr+lzI2fCmxLM46yP69eN0vKM7Q08rTEosyTa
KVcfNuv8fEtSQEY6q0LrVXvOD9KjTmLy0cw4SA5YMagsft3P5uVZtDDvzCeyCOA+
yq33G87xDNibNw9e4sgUHVR3xtUnnX9tGCZqTItbXfUvzcL6aDuuF/UHruvsJJMm
ACvy0rg6dabYs9DB+NZN/anuIF/BYXuEUCHS+MXRUNEDXD5sAkYINd1vUfI3vwAx
3wJml+OVthtF0/y47KNPs7I2b3jR0XIlf+yVraOvdgiEeOnu3owS5REB2qqiNtdN
xnpNzr4ufdfPtNU7nYjaHFfHgR65pqGu5orz7vslvFrxC4w6x9NhR5RrO0W2tDmJ
0Ce3fVuyFzt+uu50GsA4LtuAj5MUxzoCZOa2DmZ2XkLrTopAD4v9hP/PrHhVt81N
cufkzn7a7kckmcQUqzZG2J1KXf99ohf6vDJjaiadJa/4rV9zvCh9gkI7sZsYQXax
CY7syjgCZGSAWmioIoT5j4aRwW7s21yySShWooQ22drYTOzR/NI0u3Oi6z6FDJIv
j1DQWARhRZ8vsFzTm7JKmtzoqLBLkU0qH2TQ+hz0g7Y/6g/Vp8nXpUwRDsX7TdYC
oOZw9NGOqLT6cffAHJIgrv5ZMWjkTZ45QB1LByrZt55Xz4TYMADF68ELV0GciO9F
oC9S5nuMiynNHemlfjBpOEyqZgfjo/uv2cbSfUgBvvCQsQDEjiaEI7vE/YEI6UbH
Q/36zp/SOC8d8GoX4HoLh2nOT1x6HswYwLFbrimPVYWj5tDKGDoYegq8nvzqjKe1
KrYQHEs9IUxak1wobNlFTtmsbCk7BK7oDmvJ46Iz/Qd2dBKHUOrAp80XIvO2u8IN
qsTAxBrc41hlVVxbmNHk40jfufFcPbNDFATJ2PqDFBesmVezlJrCUir/qlZ7krrJ
o7dcHGS8uYv5r2QIf5/BCKntDOTWaDsiiPWg5iCLEk5VGbhvHD6iEGpieDlMc3Vy
SGpPhjADygnoEXDyFS6qI4TusZBrofmyQ+CNRePYfDfu7715d4QYq4PKZqjEUdKw
QtHwykBki/0k/Vfyg3vvNaGnoHzIcI0xZ5Hp5R/w8lSx+47BO47UtQM2FBCleuUb
z8Iw+trWJygW0jVpgKiT1rHnAmtbYbjFuAz/S+TVoBsTcXCg2+now/NRyc0u9JoI
FNSqmjVBtfjrnTJkdlWJKBk4/Tjxkhp+gG5DJG7bY4Cu8LZF7rV2/sUTEgAaK3wk
1o85z7++x6bqUoa5O3tbOFTyPlwKmMICXFXproq/4Op7INIZW1AqG3mXc2GHSWNN
6iT0Xx+GyMktQehfUCnkwBrfnQPPF3XDN3kVBMyvqZejlTVBNpHw3bRxpJAFdUam
/jURYziOHArJF+22Ww7hNBqbSginivWPuG2PukxshCc/xocsA3IRSaAeSXcg4173
W6ej3VMDVYedP29X6WaPuqpyIsh4oYYdEuBZCVYml7iqLaWWk7wC3uh9ipAFz4zr
SKFGOX7QPBPp7OtqDl2/4GqDAwD/LiURRDtugGtmCbZ+XgdbFn2MrZhuL6InCqy6
LJ8kqlXbDGFcDu2lTOByoUvtNzNvLabtUPZ0da0kyXkbA8Di1MejT0GmfLFpxe9H
j+SOwAneCianeTtpEOfHcEm//iYOAc7Xp1DfyHHti4LEzEmiXAEkRtB/5YM+IvfW
oUdkkz2bXPd5eIrpEfkK2eCiKA3JEaAecKSwOnc1KvM1Zj9qalH8p3xLTW7M3J7N
WMEA1USxD/pSDxIzAQoE0nXi6wTu4thi4yZsro0Y/GqO1SqTkP5RjP4rs9iwE+fb
xT6blQ1ddX6ppCUCXrHL00wD62C550+vfzjW3cN8zu3KHNRok57e4nm42B6w34Ok
bLm3IcoQ0GUIxm0NqG0ubKd/V77TD39NwMXB5lr3soIMG0qd0gCuqyJ+BAuMXZgo
NK+bFTRqID6hYudHVvL1GvtyeJriIs+ik26V2HBWCnC8fo2X1yB90hVFvZ6uyEco
u1x7k7szn4/urn8eKmTT3QvbM8cblMeU/9PPK7hQNx0OqAv+yWwaknE1Rxm5/13j
RVC3gSP1RFnZMots0gQevtX9AupCWJbiu5uWEbgpuYsl7+k1EFtxauAvWPFNK+Rd
ynsgAvtYIz+O/nh2shakkvFbri6scuy0zCcz3JAMidKPqKa9T1x3YEKaGJQpgGBJ
OR87i8e2vX42Fcr5mymm6QVC+6rr0nKpOYflAY3pLh/+1FgHo0AIobXMIPfhpIQc
95jNdkmnQMzaN0bBuixxWKx+l1jZG8jRzGCA1Fd91AdmTXKksm96DT0D8j5L7Ae1
SsJmYKE0Iota8adOfqOMhlPpolhyfHSoeFN1+MpQlLkcaEr9NiGLOh7D9RgOloZJ
Wy/noYd1Tgc/c+ehl3+t9vq70UHgBgu3CkGsTuz1Yg0eYJSMbJbmxcmGkINiQaK0
dYVDCn3lSrhOjbfnILjv+EtSHK2eG4jluwSniinatzUauY8I7ftmX4cm0+xmBpkm
kJOfkVu27O0hLsVvlHqnKle9rdJc7z8L1hTUrbaaS2cFhMj2q7vCZ7HJGqw4QGeM
UZiRRE213cGXOPDgJLixr8Yi8fMYxR+AIBwV15BbS7DNUJEscaIEcET4e2sGpvdB
aTb2ZbnPS+Du3IhIGY70nBlV2W9+8yPvy3a32sYw3YatVkqwmTNFxM/ZS9rMuT0P
n/O5ad7EI3hkicwoHucltqKi8/wWNnuixFTQ+gpe6Ft6osBClF3/p+hOIeBsP/zv
PtZpC3jbD0xdrDbKScbHmrIaH6ESkLZZqKetnS72XncBDS4WMDXYNNXbkCqOyK0Y
RGKULhfZdEB/icJj9kug1ly9BZJniJwaVYLCTCtYiiLSLBLBw1L3vzwnGGeX7e/a
jT99F9hj19V+/dnLFS5HYRLUcOvuEFRlSJp529PcPM/Mv+Bo2foHIOl6zaktujsr
7Xrh3Y2dRJ7HyiCZhV/YYsUnNO6VDEF6rzKImZCUHH8N1se9OYx9AWjG6+ejV3g/
pPA54Eg4Q8U8UwHminYt1haDXwS1VgAIgpDvEpXm1okcnU0QyHeVCeTQgot2Wm0e
SDKoXTadu6fEC4VZ2RTilBZaLRE5llWYrSzk4tpFc+ZqoaCxjR/ohovUltD7Bznn
QIvCjFPKrio/F9Z4jpx37LEOYaDKaizm7wJ1LGOxBrij0TfBLWFEMEDzIz9e2S7t
LSI/jvRj7EJCfG7H2llI5xTqXbu0iVQBuhmBlcBQ/dn/P5q6e2h1b3bz0rBnuSlA
BBX2+MUpBjsvoKJl74nO8rujQNYrDAMx2fcz+vgklurk0QPgApUY5Jv1GRUQ941l
T0pX19wxwbdC+z0uYTIykCYO5UYKIMlGmXSPGxILaJFZGXbUl4qEp7xX8OAxc5MA
Bk2Lj4YUBpt0uGj6O0ijcibL2TdD/TWxGGp+Ot56xhaUtNgVji9ali6vKGDV+V7D
2clB4vJPomTcTNKp5AFuLQM52dSN8sZWXgANxctz9nbLSd7B9iTM6S4aLq2HIDB8
73I75tgJYCMQZXnSBOIBwTCO084wtYGlkzoeEQwAqkgLPIrQIxvbQft5UEpWZL4V
FZIpFwn3ZMaz7z7iACmi+0sUp4TUG0g6EfvMqaMd8YkNrY8aN4SQIK6igp4t5Ul7
137QJr2WpP5dpeswaQ+r19DkEEe/6cPhQ9OvQL9l+2oQUJS++xxpF2/56JBXoita
1PEPixKieIgPT70wNP/u3MAx9hol7IZfThZr4THU/cEBRC5xHHHmAqvoiTFsc25f
kiBzh4iDiENpeQ42eEGId2YLGaDkS8xdI4Wh0IEk9dbzi4wauGvVG6EzIcZDtdRE
wppGIB/kEDWwFv03opbJXy1TkF2dgk6CIyESRijEQQwIxUmx7K2pOZTKO4uszCNA
j/xcRU6dFawIu9G+2FX9C9vL5o7ZVk8GVOeCqv18RNMakqoqCgVXN9NpbQo30YBl
D25bZ3+sgV7iod+5aavia3JQuQlf983bybmZ7HVIUOt7G+R5F3Xynpe2LiU2HXw/
QzLLMCFwOtyaR2UVV1FkdojJV/EfpoFfE8OPusUJaXq3ehUNhcuM1ljwMiY4pYbb
Tw/bkuDIm7poDwFXCUw0q3siLWrAodRatHSR6PQTYa2ymTvYtY2DvmASZW8rLvyv
yME66t3YuK36dYrDM/weeK1t/TfC7YjRInjznSickR033Ael0nYnptvX0fi25e0E
LakjZF1cCYwQkBoRRJBu36uY8VAaNYxKBOIu7C/bJb/IbHjn5wDYB8I6NTRSbEa7
+cpA9xux7Re2ubwL+5G2f6ao9phKlfix0pQGLaGxgVQH16St6/zPXu0E4FLWS/Fn
ncecE1saQUJb/NP4pj4NJAe00FDfdGnvGTC/WMXifbeqqwMVCt7Z8HULBdK6h6z5
KFUcPfzzb3122rY19jRaJrnwO2fJ/gCUk2n6LIczTctXqPlkU58qF+j2cob0G7Ok
hPaVfcoJkMzriUZhdlDAxoe4XiEGl1pUzwbsiPWe1fLGRBa7KCqN4WCOpfE8QKlA
IOI82gnHqRjqRxGEjts8ORmYnQYYQ0eSdVKvYsblr0M1RzYnpCNsBLY7EVIWA0zl
bugTv4zkPKAp1aHocL/X7Cl8f7WudOUpHYiyrTnPrwdSnklS5lMucq1NYZcp4NI5
Ra48tqvHnXVqa+i3zGpexzfVj+nDjNT1mCSW7jWn6Qq32JSr7dGsw099DYNGMJSZ
AAN5IsOikLTfTPXKqAd2Z6DUSqxOXPdWVyV/MwS6WHGTIzaQRt2kjGrKtjmihbTm
bvoGf927BjnS6S7YARdYtu7LsLlF2ebIfUFno6NS+AN2Kc4RDRabcVhKRQd7nwO1
mBLgg2wpSwDpuI8+p2OyLYPgzHAP+Q8zcwixbPHCXvYzGqQRRp9Z/lRBFrTuN74s
1C/wq14tUZQC1CiYqRxjEGbaaENjwejO+cJe7WQmANhRPod4Ye4JzIhfdLe5TLbb
hmaFaf7ylNCBAkNMUTqb8kMfdPW9wpHb+m8uT2p8713xoTqOSLdxuMxWB1Ec3UZg
m5nqbGXbpaGAV9iL/n1XjKp/3aUerdyiFsknJMhM5hVXCF30Y55N14TtoZpJxhPr
48YpQwpBCV/rwiF5J+pRdU+FYDUmXNqRHln5QxCYp7KxxaqC5djLJpxTijOaH9DC
pWkbomRDdH06WsgVOhcyPM9s+57yQI2epYPU0iKwMBKj8+wKpVhlmIY3pR58DA5w
vdKYO++0Q/jfWghY7DWh7Qwk+yyi0hPhQKEeTZ14TNNAVKfGEgx9hpVAkDoP5Gc1
E4OENW0n/1E6vE/2H4wbnSbzp2zi4Vx8e9zT8B3AqYT8yC4QKkN2YVj7Jn5ruXiD
1q2f2/c8ETX1D00DUEwOozsX++wVN7vABI1HO1odhf5Ev5SA+tQkc3OMAo6Zd9bD
bBn6iH8U6Xjm7aOTtSsR+CZgVqfA+F3xX6N33bL8k4HtxuSL+fd++5dLYrRHR5LY
/krVqJwhMtZdrV4M0+9DVQ2jUs3tzHfd5wVGidDg4Fkhp6ZrpOXSdW/0VdGGqEnn
eV8/cR2j5TYYGI+nshYlmUso2F9BcnuY2N/qGCxVgCE9tfmP6xkYOi0e17ze+rzY
JP7r8fcx2r9oKgpPJgGJlm1YDdQLcTOsG3Odmc/uMPr+aZyZO7l3r/IOkuhxDoDN
ESYd5ABoi4ZsJtgLSORX1hcbk5F6APW5NBTzvBoKgPyJwH9XpPAQQs0wo6rTwtnY
ca+/doX9OuDU75QzYnefW5wWnK6rTvLHiGc3ysSe4xOK/hhTipXZMxBtMyCTrMBJ
GAmAbWw3wA7A1MESCyqTShMAiW0+sj9E4bWOvgj+Pr//AtnYFDGN+NZwMVkPoeRv
lLJeLxHHMWCuWUhcEAl95oWDbugsYFT55isjgJkAKL0vIrzyLAhnfcSBhahZ1QhP
cYN6+W5l1yzJH/d8M0KmBWZnfwmIegFObx8vOp3Hqzo7A3fAJMrlik15q0TGPnZm
y5QYAZStb72eg54yZ0kIF9wFC2ANkS/NMXuhXZZdVPCyUj1wNnObMOFqKwcHAJkJ
sBQhM534RF3So9fTpaztHMsNaUUlrKxtqxtJ0Hvr0EBHJmoq5TycLC9elPFhA+LB
j3BwMswLz16QqhmGqT3sE8WUmDEx33O+6UNEgTmquAMmJ/QHbKjE4OOWdCUL0Rw+
06Gt949Jkr4FnmtZ/+thM/BCKzyQasb6Tg4rSQPorhYfAxR9ESKhGJVDVNh7mXpk
kxdLvb3XpPZRWhbeBtGByGs0YEMPQCtJZTwEeIxP/HcuhhiHfVAyoNUP4jerWfOc
xDiGjjevFcEYpZLlmY6EczmQXuE9cRfaEDXCNCym/Ahp5gQSQsfTFPKhOsBIt1Vr
tMOGA+TUHvsHiafnnxoIG0B24GPBFjDe0R4UcKTpDLMuG6sJuHgqFY12fzqr7T+f
aI7WS23eSvZ260hez+lFryHlwmwKR+LzdNj50mF0f4VmlSWv7Wq2Evry2jReJoa9
+NGOLsJsL0fez9Vuse2V3zfqtjKuFwOSxNiHVf7j0v99z/BQsOSwOl2hGlUgB5Oh
gTFPw2CGXIOs8EjayFZy2XWSUjOsaMDfx1PbXn1ZOBopDYKX1ysykEdmpq9mGSTD
u/qR4AXJFcA2on5S8V4f7pZY/ouWdB/VRWJM+x5yONOSnDfKIfhQkghZnrQjvQYu
FLFuKDIYcKFaFOep2y1BklduUf7px/8BS+srNWrZXcNlJ+MRZ492Unw8ZjGZIhPW
OYmQ6zcSWtcOUZOkA+nDO7p22RlM3cPIvEr4/pr06HnVHdyR1gbT15TgEra6EBtI
Nn4m15vw9cSD9VIOvr1FCd5+1Pey2Tqdx1oVlUG6Z2FWzdg5sQn4sPtCiR0hO3Vw
zePk2680F9h80V99mj32NWHukSuvlnkPtjADX9lEaWVhfFu0AU/86/hyhJ1WQTek
+XWNxx6z3w72NV7Zv2aFMp1YYuYoHoRqZrDRYpvrybXEXypZ/X6S/+F/slVY1ya4
Mv1uhb9CjZT69bEMEXtZwZztHggmTYf02VqIQNTr+VyeiKvt37SUIsYUQM5kWe/3
27eKPdtFHMt6TpBPHq4NY16HFtVVI5Pa7nqqIKqaC/0Z7mdeyOi1yKC7b4SMtSJh
CpR58xlZnEopAqaTUPJoZjguS6RnDcouS9BwOKxsY6zPqaxufM+cKZKTKXHQYTf2
pIXJbSujygolfdihZ2J0DcFWBFIQecnFiqEbqOsawyDTTwIe835csnidMgcJLND4
8IQPCVZectQKlBYQ3wzSvfVHo0hBX8E5fKF4HnAkAmW9DXR746QEjrYPOYZsrt/2
QYkpUGmzXgGKVe405Q9hUox/ORqJ1uDZgo1NpFfImwF/zr1qHcLNbVCA0tlhbsTi
4+EW52K0k8AYyo6ffYas2ErItTFyp/g90rkXfbGi9fCi8HnKCnj3mavEFsjZ5kdk
9Xx/WPnZ8KnBYiE3BlJeuPiqQfeldzmoSyxJWnFzghezkvnmy/Ms/RYc6y3plozA
jotPq3vFg+ZulKoC5lyGVae9xRRi77MdU+G+dvILlmqbVEvi/eTG/FWRVkkfQURb
RWpDm3q32SnhVkGDeN8nktV7HoIvHHcp+gG7onpNi9vPSC1qpFKWi6n3PL5vx8kN
0eI/E+CyD2fJZkhkpUIEivWqZ1zPoB5gH3CNSiuo0YsLUmA0IcNwmCt9HBZ5cW1w
V+RoH2w6jcQXwrLx9KGk3LimregivD8dLqX6CqWliXFl1wSFVpqy22mh1PY3DLAz
Yrp65g3eKU2hLSyeM3EDboP/dhywIt5PM/nXyglzRcCa7bLVLWByo85Km9mLAk98
+lcE0YblGyhEZAnwa9gOR+O5b7nxIFY5x4Jp72E6GgJ3A1EWGk2l+ZYM+8qfPomP
x6cnQbvisiuoNDeY6fnD4Vy11a8f73fZnzcZ5A5H0MUmxK3gydtrQybx4WB/itKb
4PTeFoeJUUS6IxQMXGlsy3oEst++gM5dfytXCIyslc6vc0UGBS+3abG0CTwACNxL
0LbfrJJcYBRiKu7vjb5KEPZOJrN74wZBaN4ytTWzc4g1EvB/1FYTks7wCoGLuTZV
WI4Iqftfv51FMSrGHAme0LGmA0/Ft7qrQ9idfbanipWHPaLdlSWgPLVWMVpQf/31
24nAOaaZoDGRngO8K8KyKQWzfn7RZNRruA9HbVfkLYgXNadU/UuuB4wBL/Dms+BC
gANgRK2nidFl7up6QnFEP4Ha3jKVnt0ykjYWZqKk84quoIBcKxtJwFrNHPTjGG49
6FfQVPbc0//hEF73huFiS7UdS5TR/WA7KnYe8OYokKvR4GLmc8KHe4wqMR8RmKYQ
Zfsbk1yUsMC0NjM1MJVrFNS84oiiPyKkY+IzymXbKMB3amI6yom/J7ZkljITOetB
CGNQxy8I+hcFWvkWjfjLzv66OVScY9gnQeTijimlHuM5cohVnQMTFCABz/+3/AuB
L6XmqQaYdogzaNZD7JsiElScZ2+NLAQajBV/42k2/Pv833wUR8V8FqTtrVdfbPL2
h+/u8OTLYqRrYKw5RSgufZ6AN2BoxW19llsR69lVT4MrfC8MFMuELYwlvo0dPMic
NM0n36NNRqzSiShAWEC5SceZryjGbNCalohh9Qo23HOF/5cRTwCQvsC+hc1Ftwcx
+hCOZLtPwvsAybyHryOhXtu6wPrTyXEgZ5X3puXZz038/2Cbbq9QKu20vnU9XUHQ
rLsR9jbIDIQjyHGUcwJDibGicj86ITl3Lc8N15XYUL6ZY3Eyo43w1N364KPuuip8
KVSXAxefqsF4+GE7WWDBWxqbjkEUDByS6GKo/AT06Jz2ll9AEbWHpFI8KoG4hNnz
47jRtN4qWwrD49+Isabli/aL0d1NH3T3Fr5Vs16WjotIb5XYBjB7zl/OsrVYB29X
HEWhjUJv89EASBN9dLBfwE+HivVIVl8Ig/0YzbVzXOJ3GcANmxcfTcvvEE38n2zT
tmhsiEG+OMlGdWgwqkmRiaVZjr4wKErS0664EsrIWewRkn/jTLP9OM6XOXZZ6gTd
n9253kDOCGTTwPs95BtBPErzP6Yu7E9/2y4AX9022x1xjENSO40TCZwa4JfUDjci
K8WmnGtlO4PgXWWqYSFlO7/EI4ddSpzZaa/jbJJcGwZKsQkLAwE4UENECJQNw/KY
QDYouxVp6ONBhscZDaL6s//sFx5oSQb/Sdz1ol5xwWRyXK3sDRQ/vN2C5CQFc8PN
wWaN+sv6ihxJdN4dYYdJ7yrxrB0ndkffGN6deferKbLy6hoJLKVElLXC/TUzYKy9
QMsy3dNYMC23nyo1QFwUd1eFqHPERpCwDk+3GQ8eCBRmtzCdEbfbmR0M+6ugWsn8
UK5WVsKGlTXuI2UtmSZo6dv1F1wktWceoctinUYk1v+abH6+Q7srSw4DfKgt7agw
CbmRx1N0rRhncSDrJCuMW8vE6nVj2gWyuYiS/WsqREGAAaFF85T/HpiqTt8+hmmt
+IMWD5hRMrDPMJ+FPcYFMX89rl0uZM0giaizfVxj+LW4RsLmq4iznQz9kXkqPz82
ehKqgoY/TZSoyBbKLDhZ4z+kGY/5YwzE9AhY7XYIa4DVAe//GlI9JBkRV/k+hBUR
HfZStaVTVejXAH1Zs/iw5fGhAM/jh2EVmtv7zqkPzHDX3JZ7FKF48IYkUniNGIpY
XsjzdkWpO+zB1ose8gi8EtDLddE4vyp3gohrMTo6QQXwyuTSyAo2FiNriSD7T0N4
/chvUoxAkIjGn7lzFSjETSQkVElQhfBgP9B8YKUrVCtSMXrhw0uRjBzlRJ4QsN7H
NaBo9iLYBK8Mmd4aMRXsOVuZdsNis5RDox3kT92ICfaes3uCGvSNPoqmTy/uuz4Y
5SO1QIZRkQb53PgV9zAGQAJCj1ZHtUOK5rDBHeOHs5qo3YhNIcTZZtXzC9Zd+WPn
pq0EOfduKtjulud5U/fvikkrr65oLqouy4J7njApMGuljgrPn2QEVXXXPc5LAWKH
BYTzjn/vJI24VpOlW1PdW0FxizLmT4ZZ2KwDB+zGRMktoZZp29aUlJi601DioW4u
aG6aZqtKhMrH44YW1yEnuHlZpDIrj7rd+hcZj4H04RLKqiFGQ1By6MJ/W82o67iQ
oSkw20FYoztbDKeE0WIuzrgu6bV5vtSR6dfv/Nii6g7bzBatUJeiBFQIu0IApji6
ZmbWaUCKQNS9yqfPHWPBsh/b2Ac1v1RPQ2LgfAI6CpDsVKjsek9cRh/4rzI3ChmS
hr05JubyFEcBQMTJYtL5UOFOVPLOcAXm6dzsJe+S4+Nh4e441zHH6njyNPVWG/Aq
4ROvfS0V+f9n/4t8advt1pChonHpOjZg7ZHLaV9TA7bIjcRQs+XdpBGMTeKthBBG
OhaBVGVx6heiRAr0Z7fUH/v5+LhaMca9VnY2Tp52W2plkBigDShpCPdJ2EmKUXTq
T1d4wWOzRehf+UYeIdRRfii0fpJV5d+cgp0EJK6Ba/uYvJv7ZAeSGvw94nkCMXt+
QC8BvK13XDLVf202oc2A4hX8aQyG30KQiifOzTVc4UxCsW48VCiBMZmLvmsCTeu0
scQmndDqsUkmEIeARQ2tUFcpjhx1mhRVyapdTGtPb7FQjBN4e1y9406FmukD9u04
xwRLD867Q8DFFNqJdvQxDV5xfK63NzPA4JRDWy0yWq/zqHcYSMbgs8S8pYJzV5SV
5jorewVxFk9kDyDva7UIzbJrK5ufDNbJWLf+tCuRC7tVrjaeLS1Jo+8HSQzawa25
IoXS38YOwRJ1p3/w6xG8P2bPnuD9C7JX7KCoN2OKq8VzxhO09KjDraLDPsr60Kmp
AQiAwpS2P38GX5EivMVnmXnU/2Qd3Y8mZs1XhRT2quYPNjpgABxmp2wOakbFhd9p
OmCrMX13XYea6ZaLUU/LrmcTuiO3EMGzfSzp/LJFK/+ChcG7nFVNz8R26yNYzk2O
NutOBF6GhD3yZhzGi6I8Tca31oa1BN6WJfAXBV917Cc8u8sHkYi1/2VzqvYs709e
b04vkgdVpYg/4ZTN4r8yDKxJbKDdU4HwzNeiqBlu+wCOIi/50DzFF37VME5RN0TO
wL+DFoVe75ql6i5Ud5AnB6iLqswJCzeYMHKZiRKzT8Yq6yleswLnbL/oEVmSJaNV
T4Vw96+/BWm7DEGg9rkjKsMCyRL1un4XbinZ3UP9D98tgtmdaaaTW53heN7Gbfdt
X9LAT/B8lDd1AOWk3+QnUdWcp9l4UTS4cVCDg/Iyee44m8McygR84s8S4q2fqBpt
FADY2bXJ8dGNhoF+EXp2nrnBIMPO1wDDj8LgJVEFa5SYUYcJwLMcWCE/34X9C3qA
2SuKGjEthkIul7moB8FeyPqDFbQ8zOD9ZMmKzVoccD4YNOPcVuPOzvGRPAlNr/eg
xmX+5tkU2kEBHbPE30nzpxoG2Q4SKbZ3ReyuHgPkWtDiubXAF1m0rorIWdMqmT3I
ufqd43prUjY0TQbEWOmqdnZrb11y89669aS+ueD8RlbtkTbHselKM4LRpo7nAK+f
lRkZs1JBqiC9Eq4sAJ9wsFMJb/TKKXWBmYvs7sqQdipuVly2PHKoYelfylBUa54d
ALSWk/ZxOyOtafZVUjJj90bNN1uknX2ZjS8VSrA+fEusBAOzxaV+PziWm2SxT+ZL
lzqho2Ea4T8mt9j46oNYbmLP8so29odrZASRwFPlXmDqC0EsXu6ju0OydfWnhZri
Avz7ByaBDAPoLiv0SD2dEF/Pg7TStjNW63gS/fAm/Xt8H7x+VIFGw/yTcNzpYuNO
jdQxypjzTe4T+t4nuWjdoiXrKBs3DQOVPHxeNYNDn7PwQaK/+IYNHWwWyq/kjNPz
2SOVIyz83q10O3YEGz4dRgwSRy2Z6rZnswj4gBn2Yu3wGeCayJ3drsIHWG9yvtbm
7CSZIGcJRhVKLUbACEJYaWNkFao6PNhxYkkQdqcuNxZqhK5lZTrDZ9dNql8rd279
B8DwgQTMXM3Sg8jSd+M5hZ8eS7PRylk5NqIU8ElOCzgFT/F8FeWBAhXvnF2r02o+
mRShSIDqRhRJBE14qz3mFle3euHnXZfSVgyTjeYR3CChkwEiBUhLqcF0UTKsJSPu
EilkSDsm6QvoIhr2ToMWmu2fq8VfTueSjLekGyQV3Y8tbNZC0+DY/sEC86nEIkEe
hACKej00FDreRkZEgnSIB6U+hb6szG9sxjuAhlUOODXYGhJfk53TBiGpWllS5Mz6
wzoUuCXkkYBv92yng+UWOqKvAYcBy6jAuqMD3iS6vlJcaBRlb7QwxyYZjBMohncv
cW8WiSYUND8mc7pSAfScqoOBkcpWWpNvQpNuJzV1y/Towj3oIDZwpzF/qzg4GaN9
21L+zRzp+1nsedTq+WmEDkohZw9ssAnVGUE3ONqmbTxBtFG0v7Ib7C6rMetlkUsC
9TtX/HsuZMP49W7B8SPjhxkQvu+X4WRVPw7crxD3rWnn2dVHZ7AusxrfT/ODn0XS
g5WgZJZXyYSLzFSAnYKT/MMdaugRpRzWpbSqx3gjJJtgykmw/EuUQP0tHvl1gj+9
hSKWDrC78yeBEhMo/r3aVvSvf/CU8BazlZyRR/WM05//Nv8QqgZ71l3fCjNn7qCd
2/HfGxxXgxsMHqOkOGQb7NGcdYSuHQkZtlo72HC+v6tT7F8uTEERL3ptEV7RYjOM
d80i1pUsDx83kLhImNm1cwWr9QyZJilKdJqMBYQoNh+972mGAJQnN0ZJY7KXLO1d
iIqic1MmbW4x+So1Ex3UdJGAetm9hhcS0URNX/eLhNQ1eDJXNnKYzUolig+199Bi
qd3WZi9N4GO0c9DUxTbe8ktmHmOueNtKXQshGsftNjzIittsk6M2ak7vVjGXiKDB
ExyswW6qO3FkDzsn9Jk8BCSP2dnUPyfrlWO4fPeEieRHZvZaH9ufm2jRHnIZsSky
3ZEOawF3fJiYupIL5oNEXSfsFmDyoYBAeJrGliGkazq3pKTJ7mxJDKEIi4MjQ590
07RHwkIOlatGp3kTL19kehteKIi9a7ymWzO9USpS5wt0AeaarfdXMD5+xRi3uwRq
gCEkNLn6f/KGMdl8da4ZYKlFCIr5Bql5bfH2juHvA5h8wI7tiMMyBCXneDIWcbOo
8CAm3+EafH5Y3ATQlj5wcVABCoAF8ptoc0Ge2OtU0lIwKNROHv6c5xAAAuOYB1u4
fb7qwF57RaBrH/NsC+pPxExn5dT+fYEQTGmg2OfWsRNw+nGhG160jHm7DJWjPd5/
+zklwgl0DA6VLPCYyY3d91ytsgJhnGONIr2M3y7rFhBCVUYayS+W6T1IzQzJAy3E
7/3vd0+f+CNPjZ3KH3e4vC6xyR18KOxc0qkvqOJ4Ybf8gMksbCD7o8cbr7asi6EH
TyGpa0Ct4y920ZbUpJR6IYfYT0iNATTGWZRilMV0dy3iG+2X99d0BvqjlcEra22V
AFjmXL3zpPJ6Qqn2XbC7AdywPd0CL3ZKJ9lyrT5gIeomtQDdNCvqONJhl6jPgUwY
blszz8QVf01IXHXXc/51Y0jWj+sYD5cUF+Daer3gVXRzrhF6r3NSRrMuETAGOxKS
mzRHiwbrhI5dNl+EczNxIGXGbtS4sKN5rVHqNU7x8pDfP8JZhwRj+XHF7iaPx0o+
Ty46G4Y1f/oyW0+wa0GZ5L7fI5+p+qPaSZ5d0lWDrw1DzfSgIlcjPlXTbwwa2LX3
VtH2wsQmbLX2xbfSR7pzP7KHGjQgpfeh+Ors/cPZn+DueQb6hUgn3w5tNXdfY2AN
STohnnVHxPgJ0lZovDVw/yDBG1LQf4dxnPLPHBSraLrqSiqS9E7O1n2HlvtbuDEn
cn9dX6V+j7eld3sksRKpVWfNim+64/N6WFfjXncPCEC2lX7GmxN013VQ7ADm7+28
6uvB2w5JL3MNnebDfp8DN5ZEZUNyHb/k6BBeNh5pHnSApFCNuC5eQ8MCBTGEfzuw
vhvJa9ZHX5D7xjc1v7r/CHzlOy3h68lHC1jd/QeRA6J5moFMZYe5FX7zGFDI8hna
gEBPpslL9j8nRT3QXzuZry7zjgkJD3dW4F2sAM+mzdVxChppgExpXikIBXCqVt6+
Ro+6I0byLIQUNPoYM8p0g022ZjTAsJFUMY/VN97E6N2Jfu8o5EBdWoRS5uKo7dH5
D/ogmt3daMRiQu0+mMC7Ez8qt/n/SWGBQWfS8DvXFGP5hecqEpGADjWZNt5OeCOJ
hgfSsPgoBBpkLaeWQIW71GqJ1YqVXLBbfGbMcxWor3wU3Rtnkt6DkK19Lue4+YdE
ZjNQwf8UGYTUVRaYbWmTn6AIWLTcV1nIgrwcdq+x3VK4nf3sYS/4HK+h2OcA/m65
freLhQg+N/YKAtOyc0F/cJ+mBdATNGSx85l98MrCjIP0Em9BkLIZEt7jX2XKt09c
WfLQ7YdQ0Azt/0Pi8r3DxeC7vow4gddYYxXY4paladJyBVVBa5sEpIGB7QnFg6AL
njehBh9XnmJ82qx0Hgxu44AfgAOxSRFg3gJCeZ3fPA5qQ+zBysKNCv9ffk5ccrw4
g9B3ncc/K+3IeBSNqqJXHSJ3vkwrNeSi7e4nAJWRGp3icyR0iTbNgDn7XfFnF00j
MXSYNmGyU8gmvJfy5VrNJ/SK1Ehcs2S0Hh+10o0g378bTCrtSoiXpK07U+T+wq4Y
wlfcgXTxG/LB4rN+6e+34WPaGn/cjyxrDxqgxtfx/4eJlHv9JimxBntN1aHuIG5G
zCIq1Vy/BwdkuOCHszJq+d1RsLOTcs0sQPOjNDCmZSfehbAx1W15iwMyh2cBsFll
3YlMk+mA/09sBQCtCdTZ1S/q6EVa2qdqriWO0ycu6210T6QIMqT4G3BkTjmmvret
HDtTqRRQWaXrs9cMMhq8hLkpAD68PTMmDp2KTLWbaU6zKxySL+AJUu/95O+8AA9c
tX5/7X0wbn4M6sGUVrjDjrnhYNbLz83OC9mug+YgECB8Y0zQH8F15HkP0FYMvyTy
PvOKKYGBi6g/FgthaahJjq+AjTqszjqfxeDaKmW57tggWvemYBH0c0X2WHZwMaMW
j53jeSPjT37TpCNs0PcZ7Ob52vT2KGo3+iCVa7NifpqjtKAKMnA0K+Cr8OkKD72d
ZeHNFr3a2jnFs8z5kMi73lD2xWFlhLUHvqZhbg3nYTAt+F7Bh/mdjHYi+TlPF260
j3X/UwaWITHfAAjD8jnfNPjNad5+i6PV2N4di5j6VmVmMB8pdGN3uZP5ehLyfpG9
fg48oG1rXJe8gMG0tRv3b6lsszBd7TdU9pT5wZB7Z0Dp4y7OhcVUT3PHCYE0MeDb
Wg3MrPB/yl3d1fBI2i49NMWauxP6ABj7jiVsb64olnG5Yf1VJ79tHme0TLokMPrJ
9vXnKPgBsvfE6DgabaEj0Qk95EsDZx3NUGbGCHr0/m0uLuvTUM4ovXYBzR9kR7ew
Q4f3Y7Owq9MhxqJU4LFRFnyI7XZS4JPKB/B1bjjVAhOpCRhwZgQMgZ3YqL6oi8TH
qDqXVqdldCMqKI8c3v3e20i81e+j8Rc9H5v8XbuaUxp41ok6fJyY8Z3aVPVShPXg
9Od1e9XK5bse8NW4bFefPJcC1sxThRkIxsRNomY+Dgs0r6ymwJpMooxrz7W2EhB4
kbkS4uM4P/G/orKk94qI076NtE76kZ/TtcFCpGZhQ18XZVKdUuLULQ0p43RZEDdG
719m/dvPEbaTphoUanCxptLuozexhRRDbINRV7kA735YTfHBBKCvTpwiXaJBWjSN
4hBuHOwqdPihTPPddiQJyrvuoi9VVuUUe1qv1aEhzBvDjzmsF4EC6VhcbWKOujDB
dOhntFLroUlOZ2HKyt61dKI3INDtA0su6Tx/LXS0Wnpz299kbHf6As/y2sH8e10T
+ugHMVOhk9Ug2CbJHELO/tVpQ6ZVDOCmu4LCfsD57B3OMkkTq3mAIwbrNx56/JNp
gjJKfAUOSkxietVmCO6Qyuvip9INCF3RfLpxvFvebUh5OA0zxsATGBdVHyKC9s5n
4McyzsUQbzZJXlPu9CTwv18/Za/hLEkHc2BOBY6D4MTS8rHGIOhkrNFG9L5PP707
V8ZPMWv/mvjXw5HxDmPK5VhBcdvE1TTEJ/AtcYnZS5j8f4rqq0Gz6jPH+KOiZP8y
rAKuTsGicNCpR3wvYkmQ2g==
`protect END_PROTECTED
