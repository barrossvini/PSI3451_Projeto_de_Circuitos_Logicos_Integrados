`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HAKG/zu0625z3sLbMoyzJY6R4M36eC6MJATdi3tJ+FwbItfKs3FaWDsz8hcJx2Qr
IR9CpwjN9qZvn3QJOl82U7J7yP0t9Qr7AF/yFhU7s7voL5zjZm9qd+vCrG4jQL+R
FiPHgpAn+ZgqG69wDRXVmT3cCHUfHLLYXP3jvaCrqi0x0ljywd2npI6/trq0/g5Y
tXl7/OM0d04oEbt2W18Y08QyhybjAiLDnKWFJPTVpGAOu5vFV0+KQPe84c/N6e1d
7uRiBOmHNycFp/6dOxPL9B2SVVJgBopXzkJEG4BsZCQqNRsT+xVA/qOpm1O1GyLW
wcxNHBeKOokEp3f3VkYaSDLFbRQep+3D62fouTgNFOseICh779AAIVoDtyZio1sS
iLjLvULm5BCya8fwaHL9HRXjMzoXTrPxQPX25cFxp63RWHRXfg9P8b2BKz4Zdz1G
wWelwS3MKmxTEeILUb2JDp/BHPlwjGeS/MjwqNk+54guzQZ67QQZSdFO/P/F068n
Q+ZLYgy1i66eYK75tUj9idWVgMpw3zV3miLr9wYeD6ar7M0nUGEGtcA2IS0uzU4X
paJnviZvfwhqJFf0j5sxJszVac3iAkn6f0kDZnW+a01V6yoBFxnb0DLO2rzAZ5/c
Ut1HdcF2ypyU7b+khLQiotTsfJ5bJDN+h5PsF2v1o3ZVg9NTWilMTfG7jjrmhk5q
rVxufHUcenzvdhMam4MDf5/KNCOQfD0RHuRYEPxWinwK/qmwNq9k2f/GxsbDwq/j
iFnQVTRHOCk9SApTQAkGZ85B+zTu6uoBfMPAL/lYnJ74HyvlHBFD+A/3cSRIcgCT
x3Y5WXxI2c7Vkl1hAUqEwku4SW3Juawg7vA9DRaNv0YVPUHrXaeGK2G9H+1B99jr
VS3USFR9N558AsdSBYsVMifeBn6YVx59e98eXc+oLf4oL2MQpgGnLpsE1n9WDM8A
9yfZFZ78W0v+0pOiNZzcHt222JVCk5/DYKHDJoBwgDf8fbAp7uJn9shQihKt7L2b
eUI4cQtXf8hj1fDr4qmYrn6QANJ3nZC2GzYOoBM4XMPXvNMA8tgF+IxpliAXuQp+
vYpWT+P6XujFeuXsdLrf+s1ibG8eQDVjktWwLDCGecuvHFeSt99b9PZxKOwlH/Yy
AtX+KpLdKAzN/ZPCqZ4SR8OHDBJ2660gpsi4kvVnkW72PIFGGSKr05s97krpUASE
68LDoRdPdv0LVmNb+jLntFXBRoxbrZe2U5E8zzP2xZe1YmZj8DK4TmOQM65xkRdX
Xn5b2orERzk81gyx1Nb7a1gnM0kqkuAOEEALeDGMb/vEUjzYLhYHCQqZa2cdIsaN
p7iGv8Q19jVKZV9SeBTD6H61YKZQ5IGDMJna67DdsrUBACBcsRkbpvrjF4SYEiFs
6F3hNhZHERsGUkJLVwX1F8mlJpy+VWkCpBcA7VdvFt576Iuzat8nnQufe6mRpq/K
lfrSGVuR264pIMOHkrI5qS1T5g9zRGpifyfN0LJ+9aRMbyuQmq1CineuKC8v5G58
hLSxOIKugcgEpGX0ZI3JUvDcgk9ZQJ1QssMhfEQYm3riNI4Z4SgbZgprN4uQlqwK
o6j/9Iu8CbDYoWw37gXWLJpLVoTL7viwNhGGn0cuthlPD+53ES0I+ndpzNm91ULx
d88/nUDKcyxNeWkNH1OcYTMSXU27YmqreZkQeclMsvEyIJbA0qDEPn4PJ1cVqxot
N4pgOVh+eqdIn7bDYYabOXuR+M28F+rp0wiuqR30UXLG050s0SC5d8/Q0pQXVVEk
Ya0SfDeuQyatO+CRAcJLH1zGGzNj/Ie/vwkcH0vJXCVgnI75XgrwLJbw8PrAL0nD
i8d8igfVZ6Bvbp1oJbCip/13CsuqwsxZczn+bQPaqioprMjwkfeRDpLxCSu6cGQK
t+94UfYDIKVBI5BT/XFBXnomvizSkNbIcWM87TNz5GuKLQPmryrx5Qr0l6Bh0w3n
sgDkbsrUOf6AJVZ1F/eepE3p8bNDJUBvtPyju4/o+pSLEetZYY0KKT+W34vwPTWn
2c7aOEKUxZqgeKMDsKfmC4TuYArhhgmEO//QMgD4R4hzehuFxn4SPaVjLq2P/NLY
q4GSzKpKM6fwux9/gEhMy2ARMWUXcyL00QZc3LbJBYTI7WcRtjbxSxEZ8cC7A+51
W2iVcRGRWXcGDNcaFRSWyuSo69s2zicEYP/y55DobM26F7QY/fbVUxB6Sud4G7em
2AF5IRgj/5iapBErNRDC4PIEEp597t85YLEHuYUCEhfTHBdaHK0FRUvrMjoy0Mya
2mi/aPltiZqrbx5c31Own1w7RpuMqSMJgJQDBXue/whamo+9J//VQ+nCngqQ7ztr
lucZ6ewlqC4VvG7K9omPhLPM4nwkl4uGE8Uphjl3RHoV8PGd6D/Mkt7WH0OESInT
5TUTqlaQT49gcuLvDtDuF/RWb7Ijqln3KYrnIC5jS7rAwlT+Qs7v8HkIlL9htJzC
Cf8dRJiY7HSooQf0yBANmJOYqEpRu6b9dhBKWBfHzml27YT/zzx5YQiN1MwoFlF7
ZimqfQc4NbAnx7DjGas3uaKE9QHKJ4g/V00tewNen2vwvATwqzkrL37z2b2HPuzQ
TikcYPy/zuJYo1PEiz3A0vXL3nzUW6uwYaiP0nZwMveUWYUXQN7UNOQuNEKIoaiG
HE30XvPR2tX8AzE6B9HXutnp4T9gwhvJWFVlzDbtvuCIfMxP1Yeg6ymHXQfTSQpw
e0qpKJYL8SjKfLFLlmHysJgUwlYrs3r+8IY3TwvxaReVzuRm+kgFEyzK6bXx1OLN
tUaB0fB0MIl9lzO3ZZn36sfcRzIhbhO4Cl8doxWb+sUAvQeS3o8TxNTcA+1YZmvu
11WhptWsvfuaioW9uNL6iNYFpnYPY47XK8OIKta+owPo4sAUuYjEjN0Ye0QhcaPO
ukXd036OYmonhntojZEj1WhXyH+xxpaqp3XrzDSnkw+q7vFPdeWfepaWcg/eOGsY
Gxbqd2DKjnAUBf8q032DDSu3ztxMkgef2lk6X3FKZQ4Xex5SYKF2XGx0xweF8D04
lOPkSnPVVUXnLBU3uPX/NoLPXoP8rGnlxHadtiHG0rdc5Tcpr4aTOM0OQC7WxMnw
byk6NuwmK8gPYg2CDGSGZPBaWb+DLLuIWGz86mmF8se0IMkmBITADDSQCi4g//+f
pk+IdQakRwi1HzuC6prlph2WeH2NTVMfdLzcZTqizB0kYTgeUUh9UuF3qe7E7vzL
Bx7oZXO7FNt/9Nwg23FNIGvAE/jZkJGyKoA5VE828XRlRJXCwEdVotWT5p2YitQy
rWF0ohDE4TM5E6THzqTQDsO6UB62s20A4mJN2hraE8aNmHufxMdrQB+LCqUloHyI
b3VZumTNVbDBHC3k+DKAXjQNL82oNZC/QBjR2rC/o8lfGLcGOdPSuwEfFyYZXDh+
wW2gcVtu33JUocQ7qEc2hzg8dVrvT7uNoSo0hk1VxHK2TDwS1eh3VrxUuYJ29n53
TP6UCssIOeztGy5nVisRcr+ZMX36+oNuHc8PuUEf9GrKvHZERut2Ufb0MwgzdDxw
At0TXRInHmW32Ry5fIkAEPeNbzROArVnKH73TW9ZJ5RNRjvwThwo9kXZQVoYYDmX
uSCS6oiyPI0PAwbsAPPbH8nytIAkI5GyXhT5AxK288NyWE+DvbU1WMyIowmFSrko
+zDCvyNjmzza245OMY00+Y3VC5dd+iacvS7ji7W2fEzXTYINGDySqOxNrBycWiSM
7kHkIf6cBk2VQPkohwfwfOhekskm2Kfv6t56a/5L5lDHP+wTKios+hRu4LqbVpdu
Y8JYT6RpqlRtygKRRhVVSzkr0wSSvpMCYMa6wzWM83X6qgggdcoPR0/LmX/GpEAi
O5JeubEtHtVXvuSS3sRdHqTNRmNj+vYKbmyjKF0tzEMRq3VQGUieAYl/zoL7zMyB
9Gd4CQiP/Fq4QClW7uDByUf6JjswZCDfuX+bbUGxwA+m+YDJYx5PXZIhAw+3YKok
rtJlzURYqaZ7ONaI/Wpu+K3+S9W+dTegsOZtMrOaprnInSM/6OGg7eDkhhVD/FLU
k3YNNHXPe4Xo0LTcBuxGPELMPNXXmW/R4xU7Jb+7JtwCccQhl+XUXc9hdGgUxF1E
3KvEUk4BXh/AY5ApdES2Xnpe0MIHLaOuXFzUOaHE7QZ3aYEHTactM7lQKqzdtoEJ
Dc2N79CY+lrXh0AgtF7xcXu4gjYztOsQpUeS7mI55y5VfPHxH5b2VW8aXyGXT4AL
wCdw0M+5WRJMrZ9YaO3JYMiNe80nBJQKXNx4IZ/J7WJm0HDR7Bl9Lccx5TcTaxHZ
q6cOCl5/iEZetKKsR/ziwMlA8zosfRtOrHsaIlTJVPMd9pVGu8tI3S8qD1K8/nUJ
fXQgDZ0Uo/x7bDzhDIoWM9hIj+Vj/abPn8SFfFWxpMNiZPRzFP3pJpd3saldYnbi
blrbvYUz8wnpONgsQBuJSjkXGykpkYUNa2dkpEM2eXF5+c2gZ189RzxHVAcJptiT
8XcHO+QsBa+g64J/esss9hiUNE437Rukj84iaQzuDMx4Xk3bRNl05BsyWailG1oW
WwBdzrKLupERMRHn0b3pQPN3UyzIqvqyqGHoF7KOIeIT6PbdpNqHcGQX6rCPPda1
oE7sML/TmJfS/7l4kS6X1fPHZgJHtHFSXgeRQO2gJdDSCsyHEdVtWS7lfe+0tjC1
iNzm2boSQddlIC1GOXvEQ5EaX5Spn5HW0wPqbEffMQr0V67UnqTW8kWPBCO6OLsA
NNIHadE917IjZKBBOOnNonTaR5LQX7JfgQMSA7kewzUbCnOyF32GM7m7bMVX5pWh
oFSn8LXrpa4SeRiR/e4WE3e3cSDAlp7d+1vP13p/sT8MAz+OJ5XSv8AKbZYcdmi7
X5hrMp153S9gKFsNdPA5hTtDK+AqnkiOWsIGUVSE95nKzn3agD+SxxA0YkOwpc8r
MXGXwn9Si6DHh6IhW1s7zjqCO9+a8KGCvsAqvGEjwgOi6LCu/f5k20UySLG2ySZF
/AzCW9p2DCtSwbuBN//DN+SZpJ8pGv45y6wYqw2GO2HVwsVz0GU6CORKJChQ4GNv
/ycr+HoGue+WN+caay483b9a5G2GwqC19m3IcUwVB2zbLhw++cz9DfEgi2SuCF8c
BztlPwmkcS/iIYgOfDx2Xuo1DG85R8rm/JSK358iP75RMwC3fEzGSlIvo9E2P9BI
rV+pyvEuswklXg0WwuzX3v9Ay0apRiKpFzRUrnd0ObQQp9PafmGPJkGU7EeW8ezv
`protect END_PROTECTED
