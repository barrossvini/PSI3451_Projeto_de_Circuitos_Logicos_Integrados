`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+5lvbb2iB02mmqYHwablaJ/5pk3VZXXyjfeIw30p+PVk6ESNkYkSYYiY7v34uYD
UiAXbcM2NN0DrZfR6hLlwLTlWBo0+8aMs0EVlYDoAbERG5V08E+g6GLW6uf89s01
ZkTAVDGuulXmFrt4KSQfFDef8NKOjo0O5WL62bPsL6/oXYOQlMOPGXTzJwingkuu
RdhHq2j2EhVLQlQckqPrfxkFIFQ9G7Y1Yy+270C6xxIp/BZe9jYRyDoJFED9PJgg
7Yuw3hT7etSWt1/Qs4PAkynooFF9Fpcqfri6iuaUXmd/k5KI+LO3M3BDjSm+tkbS
q5DX5iqIyxVg6F0gAg1ABbIGgDKLiuIpQCAJL6N/Y4iqkH+B9Ar+CDd/9TSdBSnT
bKoqPuUyqiAPVjCj2zest5ZYNHBKFluOAr4bILT+FnMGtvcuiOdnXB5hiRFp4kNN
4pF5MLLTdUKCEIe8bI7UGGYQGx7Xqwu6CnSkSi0tEN1O0RWR3Glg30onQNagksv1
NgHCLjCUd0viKhqVdJwf8SJ9Wh3jFU/oGXhzcFHrcRF4D3HrLYI/mH2dYhWMJiqi
XlC4q7JFwT92Dn2xZncpbU25xmhJkhYX+aTX/lahPbHLqM4D+7FK/sc422ee70sK
rErgJEc16H8Io9A3wFhNTvl1xJntcz173fGa2rxe9LsWVhWKD3ROnwOZQrzHHAi4
etcYnQd0XuMiA4cjEnrTELYpTV13sW26jXgUVXJasJT/4QA7yh+HVV0RPpGBp6mJ
yC3JVQDhtDbzEiNph5O1v/fNyAL4MywsaslTCPfhzNKksM26BdrQLBDDLc0VO5so
7UJPBykpO6NbvUClsi2OOqadb4GYFlu1QlqxjRtgUPV25aiFv+ijQq0Jy79X8nki
23j92QwkL5WrmnJ1Y2k3wR/BtbJPG+nxvmLHtG7t/nV85+ynXZL2/AxObl5IvQvr
T9CaExttKY6A4gyEPphY67kr8ip7/2rlru60f4Pq2VvHY+t5e0skkfgHarbjq5Hd
QiG6KjM0046cmkNoNmXB1lwGca08iMz1edT3M8C4vT4xShKwCKQSe9FzWaBSFqhE
KsFyLVsYoh6AM7C71A01JhaETe3EU+IsvlwFAiy/DUHGxyDLaZPZfAUlEy9NpTLs
GIpb5UHxcMITfqlpHyGFsKLS4VYgCOX6xs38MtpjAvhRJZHi/Wic4CtmHBQG/V9/
pmKTSvdecFGSoGb0TjAvNsI7WpBaaWyudWUBC3x5Hmg=
`protect END_PROTECTED
