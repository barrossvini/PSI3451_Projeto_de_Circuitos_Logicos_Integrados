`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GpvPN1d5JQ5xrJj3IBo3PrUkZ9a/HfX6suCYnqiOOW+/LVxC27vd3v+g/i8jT7Ve
k3qpUBtYA81eRRARI7H9xIzBsvaS0qqoa5d0xm+TEgaiq4YEr9LGgpR9dyFHSq4p
dWX36ZOjK/55jW+vKIVZxRyKUKAlB5qHmuABcppfWUF1/CiicAT2beXs31RePIp6
CWWqUk2U+eX2ezqsoeFjxkn/6QOoD3r+nilTWs8pNxJfDAORZNcb9x0nMtM1rlWT
Oe+Z74Dd4erVo/ppqax2GcdCFGQzu9NjIG7D5zfhB9odmGXP5CEf6gGriHoJ9Sec
D2L9xHrIo+20wMyhjY4gkbTPeHa0P6U715lQnIeL8/G+Clj+dO5l5sGqmUgtyof4
DC1dZYsqJCL+NOJ1XBwdj2Hx32NGdxVeM4pI/vxSMrKHtoJo9SjzJF8i4Z1AHkqn
ivPurtJPgYwWytS1I9Inn9/Kv22g/dhfRxQksGptHaZXdBmvj5JeDz6i8RAHecUP
Pxw7kg3zxCiHtlwUjDY9GwEB8cRtrQAs52yXhtrIVOZQMee7eWQJMyZSacHmrmCf
+7Mqu4zRZqQWbdsBcKhJNYPbhbgTBnhi1bO33dpGxgrlJNvltykOyNyxABBe1qaW
8CRWuMYZxgfosXGA56IyTTm5dliGSjlfn2PVBYFOYDrIlR1wzgVS3vnauz6ROrtY
daItlhA2tT4l7I4mXqKMOimiOl6iA7rROH1PQTprkke1CzETrpbRnDwY0rp8qBzb
+WWoo7gncj2uURxVymYHkUcjd+FSGmTFzfs0l+KvvA+8cra5/QgdQjAeD/NKuPwb
BhCOfweGHyRwNxUBOWSK5x60oIXafFLO+DbS08bj+Yls31oGZDm9AZi90jq+EkHO
xkTDV+Gm7wdJ0xxA8Vp8rs7chkf+wJQi1BgUSbZdTCvjdqi6GadEPiUb9GV6fBxz
7AEHMewXO8r+/nG6nx9YQKNOIyLDzFHY5c9aPecectE3wJPkRfZES3RnP98Tx9QQ
7TJ1afDKLJFYdTGU5eJSk3IMqJHyR/8olrk1uxRXi4YLZGHFGaCdBIfKWf6fKU2f
GaybScSJ5abYEBtYwK81qTdEs74E0vR3ji5OwSmNlVf4mJ7CC+AirtvrkreiW6sF
6+m3MXrvJ5RdzdRq9s6Rkv8raINlB3+Nvjlh2Mbdv5x8abG8rt2l4/H0Fy20Jxfb
vUAhiz4UduSTWg7Yh+Dt648CMh72ykvimRwiz8U6XWcJW9YxQCrcO/zYyOevu6ME
KIaDTFCd2lSgd7FhUSzkYvfxExYEy78jJDdzXiopJOBTUgXQJx3NOnlvOOJA6bCD
eeNQ3HP9Yd0JVdRKPCNWOCe8aMycnZgjjloSZmbXr/rp63iaBNBI3wVBNPZoUZcH
ohYNjq4S8ZyBWmg1qKtpsAnVw9Vqle6noPN91VlGtlux/QDJEMSXkSEeYEu2l802
8D7MkvOF7QZaBL4Q9tPWsux+iAihZMM3NVqCktKRorB3e+5nGfuHXVWbkFq780kG
`protect END_PROTECTED
