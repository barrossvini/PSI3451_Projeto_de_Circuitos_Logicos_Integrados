`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wjLnCfLnWumQkezimBiGTr+79RDFaYf2SRGDnEJ607DHBXMnau7P3qkF8ijHSefA
o+ycj3FTWM/qG4V7ND+0yij5Cpff0q+P34bwyUW20gA4P/aar6LAMLde77D3arBy
cc8SNl1QXBE4tvkVNaoJJGjnNq2m0r/kBLEvRTPFO/8XZQ/+5aQF5pAKE1v0JWIC
B6DTH97yysWPLVK19CP3nyu/9I11h12kCVxV+I0/C/8WsnZaDh6HHp3qBeYVI6Tf
jqo5llfWwtZvEhLLvxLeTSvQK8fWbeKQkYX0tU/PBAAqvfN8XjowuAhmGtRqWsaU
hVpDQc9JHRAgjKzbde75fAy/FTuHHeT9510Qlp7F4NSpbh8R+o6PGfRpddkUZzmM
mxTfRRcOHvnOK7orUKWdIF0QtAF2tc4jmM2g5Kr7Fr7yvPtEWvT9p8e8wL+GV0zi
LXix2NOKyvNCyRDvUTEjwyND2BS2YrE/U6flVcajIXCxn16IuaXJibjEGCrYIQkl
QxP9omyOMjc08Q//dO5QQIfbsn5Iv4ZMtV511hPYKNsmDqEjkiLc9I2zfqPOESuU
+ekBE7dis0suNOF8AXf+mAJWLbM8ei0UQ7yY9jvs5UD7dcyx3xeq2mWNwoNhPwvX
zjXF/5QJyrEZCMg59sj1bKKypi9P9DTa9RhDONtZw5Ftto8ZLgC35hIaf77joOTu
RcyGqLvXi/24j5OcBn40CAzKoy6jMPwVQXsG19o4SRFwd3nce5B+aA4CBGpofwVn
fKhZSZFBr4ZDPEf8/JnvjgOEahN80QkFnuEWlBRVKmYNUArs+fh/AWdLRrdYdt16
4xRAe8U2rIqmgFm7VVjp6H/ozDUfh/K06z6PmEgFisiWNs3oY3BoAupi8MPw198y
sAYd9M4MfNhOfml8v4AlBILEThVz9Tqc/i0n5gDv17vNzA7lefLfLw61VPxjYzFR
G8l3Zf/z0lh9NJxqFAth+D3YsB0Q5PWYtjj4AVso3lQrkL0Yt8ZICcUQnNWL7GCh
3x+zKAIRLF1rpUIN7dhRm4NDgtqzgrbic/HOP0VbA0KqWAsSlkEob8GE1H5yAxyQ
SwJc8CoyVAw0UTJHE6zm80GYBPRwfz31whoZVSGHDxYhe6IIH1VVsviq60V9c/0Y
gViFjfOd9J1e/DOFycUXyplk8COU312RSlJH1ENI48TOkWqJzVE7BszPvV1jnwmG
yEiegnfhTgvZ6kHCImwieA==
`protect END_PROTECTED
