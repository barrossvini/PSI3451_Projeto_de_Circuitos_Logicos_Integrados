`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d9A79sakcm73iV2wLNlopa+MNnM9CuzFT4Dp49hvnN1ccbfZ74YVms9F5A1sh8Eq
IM43l5zJRcvy/sejfRnLJMtCFmzJL8TfSSRDKEikE0lB/urmRAxDwpKOLTjTZFYU
g2iK3cvnZIRzbqKwxnY3AqM/ZN3Alng7mr5/NzDnbMR19JvUyWwJVBWWpdYxMmS1
zDoVl3F5BAAh4aV8BibgwfryKx7tnP9f+BKIDXPiK/I4DRz3y3e/B4t/eRDLkkYj
g4ZaJ/scvtyKkvXyX/50Jg5/ZCJPfD/kjv8hjCWcpgOqld7YAUh8yZ/8t5dIUwr2
CV9R3JUHAtRAzx7M7NBS/2FaR/FEgUFYkepZQrr7OIJZ7TNpNRVrHV5w/5OFbPtt
ejj13BVFTGmQ+RCWrpRy99TfxlRgd2QGBnHUSSEisbBqikWQ6ZmpPTL1VBKfmPD4
ihwN2NusJwdO7/OVSQsBE6/MlpMlbuOQ7V2lfCS8LIKn+q6uQeRNjrjJ5Jweeias
S7S4fF7zPtsqrSnF7dMEjKDJJmQ4KEzRQTj1wvGpnkQyqge1FD8kAObcEmg11Brq
`protect END_PROTECTED
