`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s2pnl43vJw3r+rNkKOSdo0ic6NH/HqvaHFy9wEiyjpe1Fax5vSQspord8PX5tzyh
9MetRY5HBLrzRARLcSEWVhVJYVuq0RS++90wPjTcOrY0lyQDApyuSGXettvnSCep
hf/O5UDgcusIL+fNuI9WqfKj43o2XWMqZTJ2l/hn1jntYi4H1E5vBSC1f99urRdI
wJla8cSmiRItzFFetksUQ6EepveX4ie9BH5oVvaqtiiHyz0yAkJqAyvNAQBLlhG3
GiahCVrxE2bFki97IWyX6TFRmNLxmfMaPuMyTvPLmS0+HcHYsWxURTnJQUm6bZwT
Mpxl7rhJ6g6RG/kntIrp8hfPiJjSiDJIy0Qkj8UUyyzC6U8n4Y7vjVfsIPLDAGIo
D3LKwafiEPcwLI4Kq0L4U0NEgM+SEWso/hyx89NNoF4rU8Yl77CNcrZ28mkH68Sg
WIYL0g43+jVLaSX/2NzHjqG7A1q3M7w7ib+0lfI+exoYvSxOcE30zIYGa/kaEF4L
mcJkgNwSKF9Qg9pEb4H208tV7QFwVKG6ugP3+BqhYFqMla1wsbYV7hEV3QK3ex6F
ifW+iXYYNnHiWl6voeu98OPbeLyGeS6siUb4Ewxz+e2t5OFrE+o/UIIJ+hChU+20
KPYRuCFA3ExAzLedwHaFEghPESYYhdXlQ+t8pomc5U7x2P3ZpO87myAqXbERH0lI
Yp6AHTxGZ2xzNg8q1MB2Qi4DWDSQw/AevrFu7YjCB/2+NwCdeY8wJ3GfhLKogzS2
1eh6tg38z6+Eo21oLvH60zF4foo1xRl64HnKaDSJtH3Nr5U4Bry9LHq2ht8AkMKn
f6sGkC1oBsBnpztDAjMWoXf2Lw2kwBbWoUoNNqka5H0L6+1Bdfg/modt+klu0zCX
6pUusLCLPeYG3adpWZ5J+cNyE3lEZeWJgc/y19jX4Ob6088q96spITJAVh7O7Ile
kEqt7RjCxsgOpJfDr3Yd9JUCXg+kCzuqIVISxrjTMXo6L7yrDChAt1FPQie2qNXO
p9wPXUINYIKmzeCXscCarXo1Ulwli6CJOjdfXWfEGPQnTSnodimsbc5mvZxYAAQ7
4x/mf0xI6ViBjTOuHD7o0iwG1BWfsnZavqKBd69ZjvAZ9iN/CF6Huya0gJJ0HU/M
p9A2MqKb+CHbItT9MKNKMB+94ye1i+UsQKskwOfq0UKkFoTwr+gLLvnU0c6CD2wj
J7PpyPaBI4FXJpyI3rKXv9tMJ7bZLGv2RM5p+piwPOQ91cEZnWsfqTrJ6k9i4/WT
OOrxPY414+ztlgfn9733rRNkEnJwFqr5MlueH6JVuNCo0cUAIDXXurDyuwjI0YWr
luaC6bOM/mcqmrbuQuGT2q7/zmBZU9sVxY9H2F77cs/kepTe/zprIcf6Lf9k7pfR
q+83CsaFnH/kWb7lzyvXITx//HH/QXW/HYhS0L3rKjz9JPsZXuferKlngVEdbMk4
Y1e19RBwj5ZZ82lGPj6H34OmxRd01rVWL++dFxexe6W5bktD73ZUuJ8Akqh+wFfc
K0uP8NIXMy/8H0C3LCiBS+21H68laJ6ucqEMK8wXD2DAZIQmq2OlDiGEJJbC910d
iTcf1MOfc5yR/8bJgYflW8rnPpeh9aYHtVbO1SV8SYa59EirmNmGlDxEFv8khjBy
nfT/qeo9aVs+OEVzXsPrPFspTTBzzKOhDucxKwO+yNI=
`protect END_PROTECTED
