`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jSGjVNnusP/pt96AQpY3/urR0Dho/kKAmEDahRT0MxwIkYqAu6rihmgQbeabaOGO
rDJU6n3tkjhfTIV3KwjU1/LdK5xY7sKxNmwBUExFPBILbVpdu7118gJcQBWKH+6b
sd6jaftRNncP9GBFand8OyKRrqg0muZAEvJctq+goWkYMrE/Tz6hrUbyDXwhCCvJ
SdUCzFl7FsQqci519sV0SzT3ZL9AJrFbWoiJv/s0zItH9ohXiSTYaTsiM33rYzMc
B14m5KDn/AHMhGG3oXua1wX9u+CaJgcwZshniuCF5+kurgM5eYNbGQUQSyJlY91b
7UPJ135H8bhXtU5ZB9mR/jVSe6/TmAmBeH1k2o/+vWXkVAVIPinuxGL+AJyUHIPS
42LUOtxhUARO7rYxqJ7iYwMxqpZEUiCidfiQdMnD40bED4hOLCURoOcSpmLSR2Qr
OLJTnfYzZPTA5D1QSi/dM+gGvmjWJcFsjvpdaJQt6NEPhAnMl11sNuzVMi3Ir+f5
yM9CurtVogm+Igk4chAMHCCvrCNPFodFS3Tzqct1shSaVlsdc6JSqKk8hoeTk1S8
rPLM8O6AqfoIpIQ1CwTBgVJ3PMDUjQC9Wet4YhKcwVRyVflFrfz13+M/HVQDileF
WrkSBj95wHcF75JgznKObWlFk8h3Eej4NATxJL89ziYvUnFwSA1PmNL2KC7nTHs1
09Ag+AWOj1tylKVQhvt4zdzgABPo0OOB4GRFjIdo5N6bPQRpQjCjEwqPlS0K8uGk
RFkeSCM1bgJli3wlLW9m2afOUABmMeI5N4ixqWlDDyuTEBhbZRu9ybtc7ALlNmeS
BMsOeWpyVYa1a3+qr02TF+aMGMhOaxkcWOHC20IK8v5mCWRu2z9ltaUDUI5HQ08F
dopUA27Qbla2NGiV4yIFIws113ICVuIjwfTYhGNYbk1ZE+4Lg1KYZZCQihp5HlqX
8Olri8U+HZHbErlmO5BmdChRkwar5m8ekFNdZK2gMsHwpCWgiBNoVn6f1GO8muhU
nJ5Y6Jlt1eAKG1cUVbJXDT664pWuiuXr1qLR5o3KBf70ulL+5XFmkzMkY4YA/1dz
/o4Av3HPrHAuMAdQZBvUlWtzlGtiwnTNG05b3tf+kpVUiLFdhmToMmtkIMTVRSMc
`protect END_PROTECTED
