`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HqOhxN5m8OaE3T2rzF2INEHCWY3NjWwkFs0Lr8prEASbHOm1HI2hoEBzHnCg+tLE
ULQdo4iZbYkVYmAeFRzKbPMvZuD41LX454Rkvg7XwG8iOYvZdAsx/eXG2SqE7XLe
TyXloWJnnG88GwE37AWucwfPphodpA+pVBuXjsHlog7uuxuodJ8xWHTK+TCJ12WS
7TzFlhb0MUIH2igrUSYZYJwItfomBSyDi7mbKIriNOsEsVa1vcM+h/Ewq4N+/mg6
mwptEJqJQPycupWixVKs3ohQRN6ZAybrXnJwyT7UMUMNcuwmQ+KzeA1x9EkQSH6w
4SNXnaFeUZ7CLygzXgpdd2cY8ok+6ZgOo7aj3mznrjP1T7iXxozlucrDXwCYFshD
0ZTzrUzuzqYpFQzv9cxFXPgMkivAFtwLX8TvbOUO8RMgc1Za/cgLBZb/KOOinS8A
MU0brQke0By/IDnJ3/P/RbSMIu/LQvi5bxr57Jv1UoUGIPUVbVA4IaMK1yqpBsvB
ttreZ4oURM1+4wKcwKObAIG7nBhKT2R6/6SIki4iD32pwsqxGZN+dPoqL5VvdNsm
XCRx2YXYsaXiqSTnxTWRN1i38BWo8xrGtiNoSW2J+vBwGZoG85QG35CkagZEwLOd
bQxYSyOjxU2AM5e0WzXSkLq/0/wfyiPO59u8YglCKdA3yLtdccXL28o9+5xAuulJ
NuOWzu5ChFzBwGU4yuMWGVtJGntIkhfxpx0cgjjwwQ4QgTMFO4oSQPVNbKM07NDB
iLf8yLkv86XkwdUMp0x/QZGvnQG0KPDzD5dRJh8AuFmqJK2nqj6R4K4+NCHFBxJD
5J25TsacYsLV+yURTOHK6iT1D3jhHUKwvMBQnwvWtNRk5qpKjhEKLHgJv61KwD74
dgd/eOqT04JVgIji6e23om6BmoPE/NQ1xJqUpmNGYItxNEXsiU8xex2hpUIvYghO
JGu4SrbqF8jDn+cZ5AcamwizL8tjtktMURwiW267jjvUm9ES2cnTCHkjRYDbJZjY
oJAbaLIbRPyI9wl7YHzRvP7dpaw4tpQbZVFw4ntTAXstIIPIHXJgDTCrJtJkT239
QJAUSCqEYDWUddsal4pvYvl7L5CkA2rHgt1b14TrBDVOxJZLZMB4BIFLI5M1pRVb
evMg3aaTxbewaqtybueSq8zRSalZZI3xX2D2MOwon4aZ+wJk1zyQGnNb/YojeJQE
mc2ySpskAChB7Rk8H7TCKizCi6v05AtP3rj5f9BkPE7qspNJwL3fzD/qxT9yRJjx
qDeBLvrX9UyFEP5+6h04EGmet6EIVYHIVb6cXoBfJGW7rgtwyLNUsMBWqftRh1fA
PzcPMAp1R8t6W2OdX1NwhpO4gyWlpD2VuazxEG2SnyI610rz9CF05OsFc4mHFNpY
U9m/tmFp9QgKFl6SEAqakhnZrkj1mQbNlJplOrLeCFf8aSgvY3Tx/0q0OzaxJ4wQ
BL6geWn9+s1j07JjmVIU15BNfY1a883SvsmFBnNH650OVwlhxr17gYPHYVlKRMoP
cFYA2jB1xGSkbJcN7I1T79rnaeCyciIaY391zryHcnK8nx8myHAcIq9jFKmv4fxk
W34Hw8lgKMfcBgL5cfRQcAPVrJBbrtP6FUuQpehGhK4yAnKvJTr8kQn2w4nKGokv
Wzrpoar50fDR4lTkK3C0zmakF1VjwDiY63hZ94Kvk8V4D7CRUex18CnB9fx5k/i+
nv+fsz8nVGjMkdrHKXxZ7luOCi12YjerELvPC7z7s+onLwu3hEXJvQj+eaDgwuEv
kv21skd7bF1t8fDVBJxngEuX2BGj4dvXTHcEKgjLgZsvBx3Nlkh/QE84kb7GSNm2
Oi93kOBmyCSP1CygekpCO68Rftd09MAh0osVO2XlTwK4mb7PvQfvy0HtN+6KlAJC
o17oiUZKwhpZLMMaEiDiMkJQf93gmUR98EujjpSUOPJ5UDvJX58YUf4SZU2nEdxC
MG/C7s/ab4XqIsAi2icUHc2GHs5xYrHSK+NcsLhQEenvC2HrfwhNvYVCLWsqCtjA
otX2kj2vhCss5wzlZaGMmHSkGFzT2c68GHTno2K/Eoh58psg9ebWmEYHMTnJAgsG
jOJ51fqwzj/5j6d2Tbz+rfKSR9ossKjpndjfKVFYFcF5pDtLj6uNYuiBgiN7orrG
GxOv3JtSjvwX92yYH8XB1Sq+SQJHsmSSNNdTqN73ao9MiUOF2X7AmVeKcGS8Ks9A
dJbcrJzhImRyOgHhLtd7v57bUn/9gr5bJJyjv9rCu/slkOJwNydZJ014ovLpK1fX
sWRsWQcPjRwQQPp81dYbEKdZNE7c1HIbVlJizQvUUrwJS/QM2ApgyJ31Jhl8X0gy
W+Bw0CFzSuCFFiwPL5oDayajL6UPxCGohXCBZVLwjiuiSUNbljcLCMNyLxaPwQZc
7jF+vvrXLE4CG7qHtgcUTTCMliK5L3LshDm2bdxDJ7dZGkimeffp1fy2hN15eA07
9tfZsWP+N8WJUqr05+XhclRjeAdkKvnlLN3rZdDQkuHgbl7aHV+VzQo243ir8u7U
K59Z1yp60ZbTdpRP5Yn6t2x7TYDQ2t3PzF0vLZ5q6v2/2A5eGwx3CcRae4xmfKD8
qcnwkRghdPBGdDLAI9EOnRqgQ3zLA01jD+KNEeCvn1mPc20ptUyRaiasrVuxrUt8
+YdGLvbia2STweZocrQDd/2uLDQ72ysxvpzWx0onZstnRp+PMtzh5ZxKZ7dYHbRj
sM8qtNx7Swgw49J7+PXKR0dMJbgzZfm1pL3HoqTn9JYdgjYNEzv25bUXtceFIp6c
NZ/AVsH5N6qugCQcKvEk3Xk86F47JwLZF6QyJrnhQXXQRLAHnbtTWxgvGkzZUOQ0
ffICK2G10REBQH3/EJJTpei+0mtZS56GwvFDaVMm7euRDS2EMXHd1WNGoOaL27H/
nHCHNYx/TiJlSXd6pA0z/ILq1fwcaoWAQFP5fTkW2GSCA5It63vtV+6TrnrobSzb
py0kMAh23jFYUshmBASsiMe9vK15nq0hyVp6Ky3rD3WQJUCsppoKNGvk41FpbLlp
ho/OODc28Ulxt7WZwTJSIr3zRNByiGcWaA5dtDgVjr9Ha8gznqObTu+ZjNpZ4EaB
8D33F8gEzCkFLBhv80FZJGvnCTma932sfqlSCUIeJWerOK+fqaTuS8P5Owkf61J4
Ey+VtpHkAXRM07OnGsYQp0Dem27mfgVfQMvaqF9QBiYKC5LDCkru64inaKaeRcDq
5bei8ISdrFTsgveN0V7ZZnMfuamtlCzH/MdimeSNuoB3QH9uiv3TnZglJO4WQsQL
4j4S4k8ZJj1aoFN8LqRatcMUxupo5cUVvKm6/z5gRxYLu7R2zaNHALGosak90sl4
udq/RtOrXk5AnMQwfmbNcRiXWu1cknaeVmph3OGGXXQkzRoEudSLj9avppOJTMpd
GIjRjQh58bHGbNOQFkzHGc+OryLfvTSnmUB8tm80jN8AvN+JEohckYx7XSG5Mav1
R5PBIldtzYOii/o9J73GdyYrLotX6naJaZMA/6NkRhG00Y01nYbTBkgaUiPe67dx
a7xnVO9ovYY+tpXD38VHBud5xQpYkoE0BGNQejneH5e1XLD1v7OugJYjx7cXRm8d
unxNphU911udVWReEAtAQ8PX5bmSpll7H2ct2CXSQqCs7TKwa/KyaR99wAUn7q2B
OPsbpsz1tSgVQbEYxwSs5U0po5wRmqkmC1Tp+Qx0t6kJjomGgBmrKEWgT9sO51zI
j5CyCAqGak9nhyuQVn1oBdRkvp6U/1xqUND1JLnG67ilOI6im1yUhR95tJc1VWhV
kMvlc8RwEYDS0XVT+c9RBgZY3jB+agTLlfnXVxxJ4yG4GUccMB44BFttvzqLA2Ii
XhHsidNU4A0X42iyUBxdeRyAAUDWCQgTC1vqOl6oTWN856JKzIy1YxlVYqduzp+e
CqVTShsEjzh91Z6FM7Sdv30qpOyAL+sFH9yrwZhzcZacuh13+14YeOicxnHYXqFb
UsMe1nL4/EH9AtojHArJtPKACHlLtUH1NRHuzYxXaxiQ726njmI6iG0aiwoGBnwB
oDfbEOv/svAqUVmKOLc6hyfFzqNm77mYzJ4/uCibi8mPqAReAHWj49K5cC3q27wd
Izlb0tllo4do3iJBWc368h0OT176cQozKOZ2o4/1wUaKNCRQyKsGHlMoTLVouLAG
IQRZavn0S2VttcRfWTyc2lObzpKIGpyr96nN9dJplM8UxplO7DPoYFZ2HsecddJo
Ls3Kj6ramJpysK3aqdjInoMhvkQl83aS2Qho+vy6aaFC3Bl+m0ruOYR3ql1+uxsj
pHCuEqWSi+KJkQ2EfPR0m18OxBz99qnbb0jv/N78AZst/16iv4euWqpoWqA+1/TJ
zxWc82Ln8BeAmxTw+vvxFBrKsZZ+/i3AZRB9hQcD/ltFs/EFDgT05y/bGG8s5lv4
fadrJNH4cX7JmOxQIkipTUvt3AwSoTSGWlt4A6bUR4Cqqh/hSJmLfoSIACkdRJDb
2daA3lEcTV2poR3N6Fdl0z2luqiibEw4hunLx3jof8dQBcuzed3tblPrDkvV+R0+
eGEFMbhoiYls/2R2Y+z3zD/qJX7RmIAIs1GcZg0zZXLNM2oVhWV7GZAhl2kpZW4C
PecErmX1pN20yt0hj/BuBhg1XlEcv/61JNuLOXXt8okPmL+se/cOlwPXdrGmzkGb
jqiW5g4xlliiGkjcZJ65ukRlO0zsQCeX8aT4raefLfHwfP7dq0YN1dKHx0cFWmtN
xKfUrY9vjHfSDfpQSvzTvg0WQ6ghi3yqyFiqnInQQHD3QAUhCl/24wfH135xiW5w
ZkRg08Oi1WqxpN8QGDNuWeG08AeZktEW+N33071Ge81hTDYK8pg/a7b25rDns2lR
PGGqYwFSjHLUhVFmN3srrLtAl0qDZcFyraH3erQLHWqZMYiL9srLvXVHWaw12Q4Y
Kw2LrUXdieKj6qDfeXHzSqfgzkt5VS4ELVCf1rs83Z3juNSEKhCsktnmntPCHwfK
DnYXv3M5NcNKinxgIfiAeSyx6fOaGwweVAiTtzjoI/JEP8vTpbeUC1z1gaZOOviq
/S6p7k6nmPnTHTcoR7wOIxs0hOiIyrsP+71x62TZoH+ccGCE15s5Fa8A4Qn3ya3v
qkggdK4BDt/PlLkRYwve/megcxgjGhI+H5jllu+xkIi1zO3NaQJ1Ifxz9L3nGu+h
hBoCRQLRZILgTLY731WvpOrbISiIfV4HBV2QU+3MEhPXIgzrrW8TlOvd1iO2J08F
`protect END_PROTECTED
