`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c+lXiFO3bcsphcAztTiM82rpGIxi0jTi10edSwZlpyUDh6VGq9tpXGfWIobX+SHm
SsnSTljSxWKkW7aRex9gl7RT5aAGLiynlh3DQ8LNWn7gNQcouNyD/fjNPH7Q/N2M
aAZzqjHUBdRBZH0XoiVe7xjZmFNj3uHiX5ayG6Ure/qXEzg5WlvR5dZnRCB6U+kh
3OpKVHe8KZmtXoQnDNB5o7ZYDqHgarl/jXliLuieznedJavzaokeb/2npbXRaYpW
rNO6yDK0bQ6Op83YO841SBpbENpiOSk+Ajpqba+7kgUZOWuZejvr4lnTQtF9Xzcv
AePsnn54+plQspyLFTiJ/nYYL5AfZ85ZJpcCllSI1EheE4Qbc32YJncgV+UC6xxJ
b7VCPz8rSkVOdbUDZi+8My3P/HL0sGbR34/JLwLi6LSsPaRSnoJsWER0Pu6+Xjvs
R/Y4ddrwg04vW2yFznZs67Q0DLV5M7KxExQNoYTViA3GWAKpRKNb+QbsDHMoYrkN
s49MnJYQSWUX/1GmVy4xiOX07m44u+h93N/qZf2YeYvOwIU0DpFlLR4bmenC9ENl
kozzx5FpVKJ4nOeDjkXHB2MA2Tpf7FoPICYviuiSWHwezUEM1AE/PT8uxiq/AEjG
4Nr8RmUHt9ae+XIqE1xsYrPM2EyjKMuqMFe2uW61ghn2vqAubbXLF4EfX9eWEjFC
Ozq1YbFk3o0YEybs2L/XbCxUiU4gKqzLXAtlKa8CK7Qln8pFBtVjXuGV3JL4kAjT
DGvkhl7hZHIwhPacRxUu1VN/5vzQVsHP5M/xEM764rVaNmx3c8OG2MSWrsG4JUlP
E9J1JXGVhKgFUFwmIcUgszJ7drpc8oAc6Lwgzm+peNloQZueBbc8P4DTvS/0z9vx
vIWpClTEaCZcSlNp4LW3hLR1E7MgwR/Kf2bYl8cgDdhZvPg4HRMr1LCB3W6B69Vq
abKO+AQuofI5oBYwUKGuYj6HNDrPuzLrS12gOB2e13shoDRTdGJ2fWhSs6tOjzKJ
UHQwk0MH+NlihTRDHapnSaZVRcvN+tMVfi/8G58afeJXVY0sJBRUqWhcwKqYiwUL
JDjznM868itKVEY7kqOraEpzAY8uJSxe91sR86mtT0jVmtihWy/wGFzIzHxOq3vC
Otoq1qES0KTH9Iv/ybpEyMmIdEzvzMZfNtItky6+5cCLUpylGnbUN/HBNSdpXIFq
TpBdXr4vR308p5vk98cyQfW3jooCscWykrxaTBB70kfm6i66nlT3O2PPS1/9yp5O
8VwEbfw2lc4wjPe4xouKLQi6bB5gzYvbQRjBK7ESeCN10OxL1tvAP31lpLr85RVK
qmGeba8u1n66ZTFUIYhTxEatH2+ohODAK+iHvTsYYvYKY1PMwXxe5X0awrbsyng1
HiXUBCN/8B84rQQ9XojTUcu6mbCFea0feJAYC6WlthBndP+m/EFXC6FgEDEUAKB1
cp7wL+Crshc43JHB4l767lAbhovR//HiK/J0aQIetfRyGe41qJg8aQz1NPhfm0Ii
x+/Z+esF4gfWkSrHPn6R5hz4cKMDBxLVrSo1B7LmYvl4vwAYmDnpk9Yy9FICjanv
yNxJJTeyA/B4cv1HSYQMxTaUVmUThxJswxE1TYz+mUT9ZB0rq7YUvozZJoLbRC0P
`protect END_PROTECTED
