`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KC/yVuhZU3QXAgfsrE5g232JKfN3Alnqru7sbqaGc/OnRSzM3ZHckPd10pNVe+Kt
idzyBT+0hxlMLkq+CjQqYHXLspUxiHRFEPs2diTC6ACXS2h4GEE76CUraMsMPzAO
pj/o90y8zjoPAnwzV0vTkBZHjCxXnGiL/Dtc1zUZd2pjf9bW7AT6AlXOxcxrtez/
GVrKINUbxOrGIp5p7vAwLy1R7LGfrJpUEAHR4iP5Jq1ib2XhIVz7i2AxP3xu1Qzn
CwNK+RkTULMQd6NnXjQsHTG8Nxz8f7sBhRBr791yVE3ZbZwSjiKy8Cem5H+95/LE
ClVcNd7iAVmyqtff1O8J8Mk0yvDj5FFfleo6mCdAl8I6zWDDurGX+TTBZkQ3nsIW
iV5eAtQHyi/bvz91Kl+y1cXldmbPIdIHgPw3O8OizkYYPwzzsaRPZ3mKeDaQ5rlh
kcT6dTUjp3wvG5+656baGqbd4Mkh4ngTCgpKB64SUPg5sxTBT0mCLls7BEFZbQF7
6XK/cP1zYto94JKtV0KLUW1T8XL2aWPxWFACPyW8pb52Dx2+BvxeGct3n9XP6So1
jHTP2Ju//i6CTBs2iHuopDySZNB48GbdeqoR0Rq3NVfQqVHEcAu92MJmhavYPsfu
eHHiQxWGaH0itEDCDPqpngC5djf/bzfytA3QCb62eVH3H2TdpivuzwSkRZCyqUlZ
gDWN32pO4/WLjjIIHIRPrT3/X9zZddH7W0b/s7ruSVZDC2JAdbPbeY7/T5Cc7gNk
n91a/i1NiEpJFqqiNdttGsbnWw/xQZLizzRLBLdoXZQh1ugxxK6jgWUUOXYmeOsW
toKlLCg3sqq3uLuFkUs75Z9AOsA5MyKQdknxk1yLG2UQqAtfpAGE8sBue9EaZbtE
`protect END_PROTECTED
