`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c7bnH6b9zAV+9GtAei67FErgQinTYi2Dpey2wiWYkGovDn/qzSoNu/awVvSVM4o7
G3owBtM06f0aa2e9GQb0168B3W35xPw2oVJ7rqZH8h5lwuYscdGwgJhJEF5Nnxub
N5NNQG5Z6oYZKBvCT0vdHb+Prh//z07EceSdTUbfBJO7ioE0uM4W69G64sHzzwAe
xdV3JpNwAFFbfeUiXQgkAuU1bgF2Yu3UDaoqbH9mm5WzXyJseRu3+O0ikeVKt9my
IR95lkTrpgDRj4+WXh8ddDFDlE+ibIqEbHOyCAKJtCRN0BPA7jB4nEKfOXql5Jmh
tpvQgh3oyu+oujchG1Yz2b/uHoyb9+ZjaFTJe5Qzt63t/5VktwozAEow9YX/fVcI
c3zM6i9RGqbiuy84Vujf9EjWgw9AnYaVM/i9uvLEDof/XGT5dMPDEpDkXhJ+UA3z
`protect END_PROTECTED
