`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T4Oe78ud+VAa1IatQdW0lF2y1S4KUQ+RqRswhYb0r2/u4Eijmeenm+TFD6jX1otd
33sbKbsSdiW1UmcowIphck34qdhSqfG0GRfvBc+zftm+vcyGif7XSo5zJbHgoKzg
+Ln5VoY5ugeBMnUVym1gpIv8gKY3BXME2bqROe7dwc4ISm13jOMhztROEDlFdygi
8bwDefU5+kkplpswV5cfs4zhclHqtwCLTB5Nw1vrm5BCLBS/J+SmRRtJ7PXf3Wr5
gA8swZLiD6oWrXAVksnuBTNWc6hY83Z2aKyCunmrkTLbHrex4x6UDoHPBUAgwiry
i9bP/EPj2l+YzVojpdDsVO3mY+sM0tswEvQ972usZlfBamt3ZeHuN4NNTotHRCja
+VHvqcElqF7S0UU7MvuyFCFvGXyFxs8aqmdPt3tDcXTmnnXbRcUL7Jua6dvBJAod
fdu97pmSNWvrRwmP2udVBFTQFkkcgIuQOQCoV+MChGEGM1kOMc5sxP48yAUe8ubb
EonQr8g+WQ4OOTPeNub/YI5iU0usSq7xUBUEAy413t/EtsNSTf/cIRJ/nJL8r2F8
qkMXna1iZ1YMameUA1TzStsLcWtUIUt7u0FoDM3D+KPWlNtGurYC51oKmtvDA689
4eS8rT65lFERbOL8QFpwXNnFJHDPC5CQSVClXPBROpQUDrv/bNe8nUabSEG7amb4
k1OJDnnGQMKOTTK/WNRCV7SNYGdqTiOjZAWGCa068ERTtImqbZwXZ8dYwpgqFumv
iQtnk7VaI8hMylhCcJAFQVfBauZsvbsUamF/50/NJcOxQUgN/KiWyHYkNt4T9GCZ
ZRP57AEFXEBt3ZqaU6P7TvbbUnUTdObLogQj/Cmsm2EjhcG4pQEGQsgVTC5GSt8h
PnCMSMT37FC4eW8n8lUg5SfzpL+bxEdvP07SDdcCORT3JOd57sgxxDXBjFI1vP7f
3su5FYJluQYaBc37g6clUtIJsD91O9KwX2oV4BdOrxS8I3QC2sVe1dGxGIJscECL
RyTUiVH0P21w7YPNnMUBlp1CQcoYhXYwLhUCCRam1o/TBR8diyozHvQZbcC658UF
58DMifhvxHK0AKLsYTwA3+lM2sRM3uur2seNNpO9s97VaaHN9CqgrkceIfT7lOQa
+jxrQhZLGZt+xdgMcsMvOxqeRYoSwYkJdK84OrJyFw/i7NiBNHVmUO27rKGh3xzR
xH5/FD42kmlJ2gQ2/gETUROR4enkwTZhTRvb6U+Ob+s=
`protect END_PROTECTED
