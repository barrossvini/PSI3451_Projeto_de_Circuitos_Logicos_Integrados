`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d8/WjP+0EDKFNMo2Bia14OJ7IbcpuMeqX2BKdGDBWL5SFMl5L2xToDSKEyhQ+zfP
BubMbjsBEiczF5cr09kGgqQM8QiV2GRzORswyvnQ9fGootj+JqT+ev3cQnl1h2W1
eemv8l4gOv1WIHzuS42f7JbLPvGgq48L7/NurZsF/3Mx/7G/wIVaj3vc97b1YHrr
ZyRjLsKe7mFsoIEn1ittwO/I8NQdk22r+JcB15JqCAztMiskHHKRvabRdNcGz9No
4+jal1XcWm+hosZ5fH9GhI5RPZPCmtWbqQPjaQa78V45nh25cIKS4ZeDYZcbh2f0
KUfAlIx4kzNFEJnnwfOMI0z95Kv00EVu7sWtYRsPB1ZwIf6W4J2rV7LTV76yxHxI
zF+bKb+Vt+LKbErcxnCCkaV7kTbQEzhatcjnE5qUQIAYfd6cN4lz00PBxDy1Sd91
`protect END_PROTECTED
