`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0F9Q8ZYUlIJkg8jCqH00AHpFafw5QP8Ek9vPFvWhdoFDrqiaa3rFkjiLZVLHJ9qm
PEhA0sMuKDhqCXHxQ5dt88++gyttqWk+GhEmUahLY877pEJR+JcdPSAbs+2hv0SL
6TN4KVD40uQ2wD/CDi2zTz8MCPe+nS4cuShtwsSZISyXxSJv/gu8nB4Hf5QJMq9P
FuwOHAgg53xSqBsS9l8kboBoGbG5xIfcNxm1CJUkruv9HVQmmLFpsGRTQikwnYDs
ThG3njrS30cdjVfA/0A73VlDkOaufljVFMeY7N++514s7VV7vZF8iqEWSd6n+zEY
aUyVAEg6+hjqjIjdgWeXSlC3QLs1f/bbdv2zuBxC81duGucwasV2oDtHdGM7kkrv
HyjMbnHPzgsvcTdrLs4HLtIUDMeVii2fTNeLWlvyRvxa/1Ab5Py+njzep42spDtX
eQ2mJdCSSo1QsgQZp5XcSCa9b9BNwjJcL7jr537Ck9PMBcUbnW6R5+TUU96naa2y
DzlvVjrIic9cSG45ntiyEs+GsV2pAf/jBhTRntODRfWrMW4dUlngM4EqnL3wKwF+
JeMelS0ON8YXKnBuX7qlfN9j/28By/7gm6onj8DGKGlqfh+fBO1lO3YymsnekmUM
ZMkshO8wVGMlcCJx1r9dFAABD6ennFIxWYfTu6iMluaFqreisGIIGrsobAjpwJVa
mNkyqTpJfaLInbzEB0YgDLexfpuWQ9XrwpH3B2213fybs6KKGOMHgq0biVugdiC+
kw+JQgHhxzUMwMIYMbUDb6VrGvfWytlMW0lzPfZWP9GyV+m9ZC3vtTbCvpP4ja4j
SuRbEjFE6VmXthTgx+DwjoHKkJre43d4B7LPEP7+KB2rM0YOBg8M35UfCCNgaPNx
UeZ0fWMUf20SHhLpXDjenhpU8pg4kU7II7deS7NGmii4hjMv34L0GYwvEgomLZPy
zbK8LAuI4pr6nk2KnEbcnC3LAnr6ilz1dDW8SvavBij+/IInzfykruy5KJ7btEKO
qYVuCW/f1EuO4Cu1ysXqgn1aNqRZDJVXnxtOrbDGg0L4E75OKGKB2lVvbWp6+Q6L
XeLPIalyHdpQINIESYKZE03qalrVfg6uFmqip2h7U0+IrH6VJKp+NiejddXFVVDh
Yffd+bDcKDVWanYeERBsS2PhhlI9J6cqLcNBjuUar4KfxT5eV9zIoimQX2hAEb/n
elgeye9YFXQv5vZuM4VB4+fyR9LPfufwJ1gACj+AkGec4HQMPNhYr9Lg+qzbaMHv
m7OaOBs4tsDtq8fg1r9yYN9KnKUZZV8gT/6qdnyyeqaSvHRq5uR+lQ6HCZHCELEe
xrcah7NYuwTsycoJI9qPcQcVhKgVV/Wk5PdODLbAozgtbvXi854JfxY+J/daqJw1
A/JrA0FraIKntSJZrMdK4EfdD9B8OT3IYKGtWri+0FaKM27Vh2HC/8Q7Pfs1HnOo
OJLdNfQ5qvMnLLts9xKgogJn6JQIzkrsMvmyA646Kax/Usqi0BoE8MQWdBIaXAkI
UjMPJHP1QhdHCtyrHqkbbJtcn77t5ig0VCd7w7he7ev/UG7bg083p3uUAR8V/EM0
AgueVWKKfx/ee2MaR/o/gyHmAYDiFuBhjC8fstzyL7uTqCRiYPjI36UBBWtNXsPU
MsQ0allhF2fOwrbxIa0wT7mx7d16M3j3t6tEb/0xrON9ZQ02O4v/Ah+fvTQLUIhd
O/gV9iIzsDxshd1wp/kHeLPdhVstlSPcNu+xJcv4VgwC/qX8UQ7Mem8o2XR+WEA+
QP8vye9vHmmcLQtC4bWyf7URDeD+d7P+6AKmSLEbderewLJOmD2OWLn7cmtWk23q
7BC+3RBg/pqCXIsTekdlJyJPEwr+gVd5MWl8RrFgW0oBzetua2+xxGT8vTmyXhXW
kUf6Y0PKwo8UkdYWR9j1V+BzVIrciHlaa9T/hCyMW4IBk6kpUI6co53VjqSBrNea
9d2zGbId64pybwH7rIORCFU8CX8YOrkSCO1UeXTFTQEgk3qG4NdCPbBigYH5EWcW
LoGBPDkTlG1Lp2VYYk78NXqsmFtUR4pPgPdvug7GKHW8G7u7/zAtljZ1PE/nI/tV
13hxWTHbtjraAnoqliYOQ5F5UfkRz2f55WEuQAV3tsDso1ea9EB9fbdshsSJXKQ0
pgs8MNJ4B7etjyRiOEI7Cch1rPuQ1nLVmUi4EcLYF7o=
`protect END_PROTECTED
