`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
htguZLnWIIDJfdQLHYVpEjU97KypVMDObjRDTn5P3tc83PCC0VzLC4WIt/R5k5ZX
gJSjid2zU/bkbKNA/v+TcCIYnEEbsQdKmq1yiavnvmBWfkib5gBzx6I8ip7gQj73
/91hIz2egR8gHXEiWOBTG9EOzC103MirKz35EYy4gkMcfL8AcVvjrOU6JhcwS4SI
yu8grVQ5leNLIFpaOp6aHcZi64GsCUxoZOna9BwRHJtk4kzoh8D5WeplrmkfClMj
v8ibT8ijjd31m8k2bgLLst0RObMwmvmhJjEo5lNUXygiWVRziByVqSxr6GvHtjIe
E9iFQsVtwV0DbNzct0YtPcVKBxGL4ipAJsNg7l7Z/uPwd4Lm9eN0A2kHIQpkF05S
+uC4/Y+RBZs0qIrHbmQgbvu7z+49iuTj5Q262PUWFA+WaI9i4FhB2F1kk5DXQlds
`protect END_PROTECTED
