`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xuv98xhWp2f7ok7qaE4BrmFrfveqwbg3f6FzkCc45hu9q/Q69/Jg4zX+tqMoC2Mm
9gSe8ZA7Lx0EO5a2ucsCCNhPPF3BXQu5NBRENZv1NnWKaLSE7ce9r7S1rgRAhbGA
o2qbJzHF9VjzD7mapxc6ZI3jUiPIwyvu0nTv/5BujUDzY+VkAoA3HvBn9V+mCEIM
N2iS3STdCWVFE23HNcmkwjG4SzUCuDAqvTi+0YXNPO40C3t8jeNifVlcl7Jw/UYH
7jZ7peThdboc53eyJQEV5vrG70HDflHraV4tpCWVIQHC/G8mPbCAEIJVby1agyXd
SRXr+42DnK7rscCVLu802AwF94EJLaGMpaKgr3CqNNPhqyuv+OoaxZkOxTKYnScp
T8Njt3bW/6gThYClFc1Ae+gjxIwypjuALn0vePFIvMAePixDo10jiIBueEYLVtZq
Vjvl4oZv3qWJN30W0bSh/t2IF8eGU6XhRvWQI8aGAhBMsSHBgIPmPyNzknyzUXm3
KkW60zHpDp8Wfy+FxrDkc3FA1XNBUu9J2TPsm3dp/Njx1cg6DOF0x2vcKqncJ3bp
HgldbE1pbiZAdlzsQChoWC85HAnk2lgkYZO/zWdELxVbhGc51r5/hKHfJYume7RJ
dTm1j1WXnyaGhTK2JdEYpiAodRkHBoCdrKkJNrWnmdJmhtCvB4r5cgyLSeF3x1J4
i++58ocBjO/FiaVYTqIOnERElC/Vi9HsCBZT8lA1iu8vuQmdziqvWJIXm6mKodru
kzgJ8eCm0ZFl9ORQjD+ln0xCDIafzpdee+b9hhmP0MTfElpYPq8HTw39Jk1ShAjg
mS/WmwQCsZe8PzJ6ufUxK923XisAz3HCM7pnvH37symdPktoEdBk/KMbp/5iZ/u6
J6bOGkPEyMFvXWKeMBegCUcSXItE9zIf3/wZxul/DuQjJQrVyOlhbU05W/d76mYK
dgsMpAo1R4r0Zs5vi2hKge6myHK9XI7eMpiBugb+h2RsFHvelwizlTHHJ4YX3+GZ
4LQ8aZ7s7laxkNDCYr73fCRLDjQ+TkL2Zm5GHL203CEcDMO1kAMJqRsUthdLytKN
pYEJCBDRLjhXxd7gUZzgJ/V0mn9FfZ7CDhwnjhnBSqdkvLAxDSpY5qtl/4PEcRwb
EcLKIZbSQ2USHDe/86eCCJrbm7RqlLS4je6CViw4zs4nidbUat2gz/tT1P1Q/lHA
1DWM2EdqSo+3QczHQoNXSOS60I4wr7HPai9IDbzGhOqFOC0GA2jRixVKJj8lsfTd
`protect END_PROTECTED
