`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QSEdQEiTZXFB/nsDuupkrdaWZIH9krOGY1zbRzwY1Vzt7zEKYv6hexU+rdF1ciGn
Yyx+NpoKvIyg3bmIdqbmaEq2bN22g3ZTz7LjiR2XkaMUG4Jrz+Gm6giGgXewQz6R
PH9ikqH35VsEQmqtNS+oxD60VOlREZd+oFAxoh+Ze+Jx5vGwrO3GxQReBj6b+YRE
BE/001ofZBGOOGrKvNaIsis9wYKeT5k/kS4r+2UUtIxa/ezcDxwR7FfM6G4U/jHN
6F7qn/KWU0c87e5eLpwfBjmQQ8VcHfA2AC7RZBx56JkqtToFyZ70wZ46BT3yvtp1
lAIN802AOBHCNAFenPtKWBuye/e2KmKmQbY0b3hTPC87QtMhcZipNSqM5EfA8xJO
YdryBgYypZr2LxhjGV+jDzuY1Evkh9kWk33pG1YquCMQB0lYdSqEab3IDY2uBJrl
HwDfAuPLNLF1OuYbZtQDVEQPGK7XMgMPZ5cE6832MlpfeDX9ekp6p08erALNKKwT
fDZyXjWI0yuQj0N2n6lwEtsfqvh9f8iQ2dyNXuy/NudutDMWBbMWJVA6fq5PNhw8
zIz2cSG7CNcR9t157WuVwamn/VYNlQwQlMa+8dpSEZBRIP1qQdK6HE026Q4+WFej
5ILd8lGy+XKjwkM8Qni49xQDssxxYYTx3vr/L5tuO+tSboXWKwGlos7pLiEW/dc0
VbfhRyqVAqAzV6IjC48ey0jo2g0IDEFCccWj+1qkb/bis4W0nDLwf0DL85W5kH64
YK9dltkZAI8DhGqnt6/fm/7RZm/B4BMCt/JLbNIJR5qA/FuorhVDq0at79dZYzfZ
Cg3/vVE7hc3gChHSqEdfX4cclKLXeNJxzCewnGGCV0nsr+rQPucFrJ940gjU4H50
srIEEUaE/QdF6aSp9KzGmQ==
`protect END_PROTECTED
