`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z1NmLFVoVQ3IUoh4GvxLruQZy0k6dIiFCdqBV71B4Bd+L4I40urrHw+G9s7dryFU
6z+nsqENE9iCR8AuAyD2Wi3a/w5z2uoQNGStx2IKGiP6q2lViAjdf1Mc6Ck8G5s3
sEyiOw5XN8EHfulVT4wQhmtS6kccCFiqFq+b5XWA52vJxlpjxBOxhBktfYMJAr3i
TyY9AUVnlAb4cbfmAEk4arywvsiLs7shn5J8hvWANVdxRWwnLEmW8aK6k2G7W+W+
Jdvfhr3oMuFHCcLW4bh1tof5DIluKWPozdKTsSOBgDnw4e8+eZFhSTVT/4MVtyIf
UtOQW6YrLm96EZyWNAu2HRFLxGq3DCDjHYIK95hn5jDa5yRAmHHidE2y7RiHdSXx
`protect END_PROTECTED
