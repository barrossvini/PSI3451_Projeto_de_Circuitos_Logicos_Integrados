`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pxlso6JFn9ROpGGwSEnWy+MWl+flWs2FRO1tNPCtSQo++3NbAyZCqB+hNDeSNbRe
oLLPIGOBzfPgn1oxRHOHFFTAMvLopEwhacki9aAOTR5wxlBFwHmQmulQZXWv4VYN
TrsoQMaV2YALFLG/VmfP4lBn+DMEQsJ+Gn2VrXtq85vGYQrf0jZy1/vsVhUHMnQ9
9ztUOVGoj9snb/Fic80+GvsyxYZyFhecFzvg2OYXenCnSGWVI8zfDY8zseVfKnw9
mpq8Z0KDDWJ77ocnJA6D6Ghtox2eCHocp+IemxK5t1VRh8QijlpdIkwv4hpiTqWX
A+zoV4JdYYcRjQwDqHi+6C4UyUeNymOmnyHKoxV14MtNkN6CDfpbjsB2SAvQFZnq
`protect END_PROTECTED
