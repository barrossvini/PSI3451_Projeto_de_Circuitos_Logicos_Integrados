`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wEFwWM57FhHiFShUDNirIx9qOT9jogjVR0Hl3id8SR/hpMgcIZqpMahR3XWthEz0
AR7NzGTtzfqjBcdr9qUGYlC4P1bja1s6BgJP9pJJufqQT4yCDeEdXStPQPHhqPzv
DpRps2+ivsU+bdgl57MinNy/EsEZGJICTvynhCsI+8q6RSf0Gm4Vd/nd97+8o6Ac
Yn2jwx7w0xqcWOd5KlB64FCWgdhnwWBM+L5ObxS58K+td/2Gzu4bqQtODPX0yKHu
ndIQ7Zoq1SaqaqCk9doTkh1yyrI2tlSvvN+kIdfA7UyIB04Bvv/3bNW8v8aCYoIb
hOIu9w0NaFHyHtrz0CkNYyVJgZPNG7lx9YuTbkfdH3+uomAUgLZOpds8zetEYRni
xM0/slyQM2TzquYeZdoh8xsaacdNOKJSpMAcBn63+9Q8FJjdRlt6zPrz1klYWVsy
7GH3sBpkOLeIazPuxqc9+fhkZxiR6ogTGrIaETkGdsJwK20x41tbGlo9StlgKsjV
VMM6rjBHjoLpDowT+jf5Je3VPWvK8mH7HsqJ6++dgJVdxGeE5KvDDYZrQlOssTu9
PIdAkWp2h2rbh1DrWCRxIV6gDbtj9RFJQDMbRXeY5uIqb7kai7/ohRZhRHZNRdJl
IUcahAd7wAAXYBQHuKz8FY8swY3vHlj/yZCtrl6+NDjzdC07BYN7WQrgn8CllwCt
wBEkqA4hbWHXmybnvayxgScosceatW0wAitUf/FmSEMUBAGcz+uL+7S1DR0kxEVa
zFG0k3mHmDEZgtMKTAorInMQqU6XeuM2582iqjh6gGlFHyNtreMNJhd8wZxvdQym
GNTFsBe4+w8K0CvJlEK5s/qfoCJPhK+/6TjfkujFYTC27k5wvOYJjd5Fpi5ZS/Eg
mWEuK5QegxCgGbkT1cnhnD3TLR9A3UO2r7gqwJpJfD/QqlmUjULAjztO2etnJ6Vr
nKupjC5qt+ZJOUqcTwuyqegoSnG1f53fZ1Bs8Qv79GjvNifDSSjNWkTsazlGqXgD
vannYQm88VZD3hOFjUlv2J2KDSzkHir2tKKWHqSGGZy9WScoG822CZxryEmq5Fzx
Aj2qndGMgTkOxi/Osrbm1SF+TTxMUcGkKfbIiPDpBaGgGzEyM8g6otnoE24pAl+u
kYyy53XLXacAfer53OlzxGtkFEFnJqdOKZrp5tnwAwEZimj6Vaic/1JH0No5sq3R
PxjOgeFWJd5aHBq9hLPPZITsHn13NE8y+qfeKuZ1t7YgzceRXvl1JAtjX/KcndoF
XLQQ8KtPL2dia3jJAlI0Mg92pkjn5kSTCHr4GK6EUuY0HC0Bly7VvCw8nZnEgqOW
3HycFOT1CxZyDW7VW1C561TFY5/QtBL6Nf0jOP84gj80HfWhCSGSOWP3TdKqTGNK
isdvVAFBJWe8zsOuGyaPzX8uwB3dQZbI0TrBy1xz9PKEqUqZGn1VE3a8jnNx1Hrc
kXDUK0Sf1WLbp8VpkufZHwZ4by2pF+JxKN1H9yEPCzjCaO11R4g9mXGEpEPn+E60
dO4/pGwH293CqnlQEgpxuqoSXQvE2BUM6KgsdYnsDj7IU6BTLA/svLJONipV/xN5
xPylXHREhTlWEwL6Zx5PYu54RLoxBNR7unJ6WFchDifTeViQellXAEB75LFsVR/2
ly0NiLj3PO/aK1VFefVMvletxvLxTQccqV5nH9bIp7HE7tk6i5i21Ag/13YBmdDn
U3gbSXSwKx9Kinzp1KB/H9qgdXhUkmz7801AjB3Gu/zdc/1gytZzDF9KdPmrzps/
uF4m4/OEDbRlT9HITO/OzH8DURnRUlnyKRnYb9/7LYXjWxzatpnDyr6lIEhqr2wR
NFtzZAPEuy/YaX2CkDiLINcyjAJ4LmZ50tOlcU1ScX6fOC6okafFIJFe6Vtxnyjg
BH0Wz8FO9K/uI7VKTuX3Jh5m+dsCV0f9cxszSuyC1vzXrvNV2f/TKmob6sgwm6rf
g6qCVLVGOgMckCbUadFdVNJaqEehTcpU8gmUuBKpxweldi403tf0F4hvJ7Zi67CR
pGNdGc5tC16b95/NdFidYlZNXUJWw3/E11V0wDZxuYY7V0/lV0XmJ1Bk6Ob5yVCl
YgRu7WMP4pxnsL7k5lgUet63ZTRIX/ujps3cW73KsrYrGFWZbTnL/W1KkY9i9ghA
ZEXpBFWlh5aMKpHITpqjKc4NzJo/Eq7WqePTmpsn2mHwEkmqJ21PFGL/67AaAvY2
ko/e3mB/8em4Jeto7UEGtVD7Vg/WMi3v32x8seEOlKN4YPVAl7jcz1JiscSrlgAA
xlabwjSA9We1fbMfEYcX0mfBhHVlmJ+nEu02fnL90OhRgfjgwytdslF+hjdQEbAP
azEiozv3XOIzXW6HXzQUfUWG3qLh0aJ0g6p3rsTamA0oQREeuhGKJNtUOxpzhrXh
vul4urE+nzS31N1EAQmR/H4Y9wmdy0MVtvXn7iW5UmITb9pRAcTIuSXvdvlBH9Lw
jJcFYOz7yDNo9s7YSyGdy+3mz7SW+MhtngbHgABB8M7H1FSKwgPn9bOVoiBrF/Eo
P8hXQCd919jT6Y0oSdyIMDd5NpZJzGzpVe6XREvLq2hu/ou3ggQ+dfsm6Ok92jgc
48gbv4ZDze+jIZprj8JJIAOA+PyJJxCHZYr9fQeT0JC4jeI3qBcwzPuMkipcVkcq
iLpwKrE/hNntouIzbZeHWo0sFwbWPyqkMgCZgSKZ3I6hz14avUpaxx76OFsAu//C
CNgfpGZOWc7BY32Qf+akunZ6m+jdBZN5inwpkRFKlXuaxPwrGfjG3RPbGhm2HzeS
Edy6mt/bRRB2u2GEN03YLZEPVG/CDLqvwD7Z7jv+FlaN7mmJFrTopd6cY1GVdFer
RcKWgk3hoy8pi8xzlLoXlVx8F0zpMIQznbj19YAOrEHXV+KRMEPkUgQhUfohq69W
pTiluARuhdho2cNKTGdPtG8XvtPNLzaAY58xR0v7lfC+duwzQSRZRnFdPY4HfW2V
W9KvDzISljeodr0UuPtYM/2nO6E8XtFLRXSzN7rsX8gl5owSmnBrHMBRTvXkKU/g
aysWl1zADq7uxikY8XKlYe120NdelVVJomZ0WcdfXXzQpvbrCTCASJt5u9ljKL+h
x62ApaH8yGwvGUJq0aPDVPw1gwrOToZ5g25aX7NxovcK0CUo+EGkaa3S9Ed/PNvZ
yAlTh5/ejtUzul8zn32brxMwwI72Vri715whM2uT8UKyTnLyGNMQoOvzWaA/RL2d
50NKStQKjPpvqGGTEjJInE+zvpzc9VideVWTz1yOE0/MZXhjLqXuMym2JqLzWyhn
qwSzH8qMHHN4ZI1puF3ezYPbHRHLjMnCvKEKa5l+C9enqoGjjLEonkOXZ9yI4Ncc
Uz/c3PUHycinImd128CSMb3p3Layxf3EINbq+EKPDXFvTdaMPL5Qp2H5JpZk/qcP
Mbqe8NeBhijFE9FwOpWAP7S/uarHDxLTA0ubZM2ai66mcqsYrHqv/8FXQMigoX+O
6cpVncrmHuOW4ODBB3qXrYGIjC+MQsYVsoL4q7K0SGaVmqs6vVDjYRggsFjZzvcj
VXM6YPSWfI7BALEboFwmIRL+8tKBDxnL941r+MWfStMgu8FnsXEeO66YSFY1F2dz
6cFRIN65BOWvjxbvP6i8noIeznAEcAf4Q8oim2/HFxZ35CvsenwvkEQqxtyE9KC+
jAuceYPuqAA4faFgMckV9bnbidwzM1eNna20fSoq05+OmZN+CkGKL+TFKj9txk0R
bIl+pIUwbYYr3wt2XWhcPh9PxfyHAXt5FJm5C2D6iz3YvB8/EU1AjyAfGv4P8xeu
B5Pp5avX/tPtZgMu3X2aOFRy3DZ5anPCaFbS0xdl5QkZR+RO0sFEHykFMFPYrlTJ
ctjsIrexAoQG6BHW5aFYCRYeoy8Ldh/8C/Lo1ufC+O/KBdGRVxxxAGOPb0s96bLZ
NaCkgD4R9U2kocLCaGKGqotCAn9svKtQJ/15tAivpSPLgzu3ftSVvcjsXHVyJ6iD
dLWLGxWgKregCi9TEL6s/1COPtvVisDq+xZN31jmORfdY2GItG52Crk703E6oARL
2TPv5fEcAtSha2TZ72T27Ytd0yByA9L4Szmu9fSeBM4Yvo/k3UkcGSChiGGk0I7m
9FUEl50VaxK9VoB+nCqV/fxYMK9uuVzVBnd3j/AG+aXAqjjE47+KelLq+eV4j4+3
SoyzH9MHBdFDYXzBTIW8POeuZzoCbySawnDftRUBkOgR5j8y2I4t+6UeThoLUvcX
HPXe17Ji/HI//Ez+Wqby4vU6IEdL1g1wV2HccjcfD1ieyxKOGYm2QJ0d9ivNnEpH
RQE7s+WvDfwkE630r5oOGG7AF/N6cV0fksRXl844elOkpL+VX3byuFfbHYC1VrCg
tWiW/zOTZvlyovHbC9eMH24PU0PIds71BykBfwKUXWeS9HhVvuEGQ+xUfPWgZhWt
b+OLTDyEbStCCNsFdO3HCLlY1eEXG5fUmSTzjU5qvcJxa9D3qYpNYIZoCqJX5jlK
yWjpEHAFTUSSJnwWQGsWmRuC4lHVd0PJMpAdjbZ+w5z2trEc41gHkS/99aIxFi4f
v7QbCVsJ/ViZxMjRGWgTOAdJ3m5IoS1wuVuvssgoJeoz+X4ZVFJo0iOJ+FNKsMDX
unr61STVVzBrzpcPOKqHp06rf0Kn6K1O1M17nry26MA0wpflUttJaQfRkRfY+anh
7McPDnAH5elUv6zprRBMdcpqOYbfj+4wl3chqHdUWKYTNEakBm4w9NiQ2QPiYefj
hGG1vhrfxSEPpOCCJgQBI/G5f9xpcF/VSwxsKRbCzvCqxN60/cCLOu1atWJ3IzDg
hw9CdQu94RTpg8QJaxxIZP8LJ5ZrceY/ljcDyDTzsGmJnbHg6frD+vvZl+p71Rzl
LvBJUGcHU8pwB2RJL6hGtZiStzBxMAx1w6RMcwrhJ5WXnaO0fpLLKYayVw9UsEY9
58GUKc4QonGT8NK3cENTJVZ+dIW7r5pB36iUwpxtvzh/PdnKqlQ9B0FzRrwUnH1L
w1eEwl5WLo98eRMnL//JBOzUINVtZOrVeOZXJBmGmJNfP4tU53X7VdMo5QGA/08e
TUjcGwTtFOo91mI8RZgOsUV/Vzi0j65K0GBnJKjsEREk4uG+mSdKlX/dQBdo69YY
GDR8R1QHddHjXyCqBtMq3FUIFzi5wbBNMVnJimsRal48rtes4SBFZT2UuYq9M0jx
5T04lWc4SngP2NB3IOucMFQe5wNjOWK7u452W8cBGb0eZtl84Qary/16Wigp6GEQ
uLDwJ2NCD4bDhYDjpenoksZZLo49vP4T+YmQcFBZJv/yfqUfpyUcdNwDYY/JquK3
xXZFmj1gZnn+o0uM1ADhNT2VJYNiJ4OJW/0bV2vhDIADZ7LdOb32vIpbEvMbntVt
ACVTtA0Q1Q1VpMakXQksUMLRotQ2MzYg8zmPLFya63PHpyhovL0e6kvvrSMST6KO
GhAWu4fZwixE/eFKDUvbvqq33b+20U3h1Cyum0rEwDpHab/M8JKrbN76tNQB0Qji
J/CfF18HErJsOmS41wSfmH5s/d/yQxx5xfK5CkN4UKRf9RMJG8GxxYs4FpzdSCAN
NrQmM2CKcT8/5ZK3BCteXXTSRH09M0toLA6KAGiCq9Hy1lpkfVj2EnzldPW85rak
jjtfY8yF0orPpIcRip4zHUEb+iUlC+ETSpFZzuzdWVAwBOIiMeGUtzxh/dPNxHLJ
wWUJohB7nLsDmdgq2VPrYNM8LxLnSXoazXfRryHvJ9E6bnwJx/aVlDTg6tgERb8j
SSe0hS7fxbPQu6CXRYe1wb9LyEt9xxq7SLrx0mF59hOhcFhY8w5yF06unqeyuswv
yPP0NAF+WHlmSolqnCNDoSLUBKwTflLAloowjyVrgDoEbKtyDsxJJScyzaLPh1Qj
CTktaKzlIJ5Q1XZGte2u/hu4nak4SkpgODkXfZdIi84odTWS4yMuCNMI8NGM4LX4
BK6yt/K4qpwnEqaraZdi/FeeLrB7s0SL3YJzDPQGu3ctaa47dGAfP9CaABaeO1Hf
SCyjsZbyvShVyILP/sdzUSDz6hcCC5U/AFN7V9CyhOS/jRgyaXduM64roZ460bk2
y1H22tufZy1O1lrNuuRpwzHblg1MmvZDpdkmIn6iHH8bXupgU/HIMGArVvjZgCAH
Q1yKyHZ/BVQeGsWzy9X+yTgJXpv9P4VxyTIuEVuS8KXbP9oz690vdQWR1JAMQ00y
5JptnATt2keO1PRJmJIgcyYdbk9tHfiHMPPP1JQ+ngHrn4VMt3Rx5e8opw+/n+cv
4qSfMJwMnfO165IUZI7aqfPhxmR+daw/he6gYhIq1KuNtj1Mrnhl4wz6iphmsqQk
NJxWIjznfVcwXIhGX+HX6n8sgAasGxUyIBOnfUEVNqOM1H/YsibPuXs0lK0BJlqs
kSwb9weeG3fX12P/caf7Qgva2usjjKCT5iW1l9ikvLrir+F8VS2XgMrlVDtjNKYn
vgs1uW4kBME/TXw6c7h9Gd5aUR1OSno0yEsRDONmVUVc8fi3vukfVcn9TplnaNh/
1FlQuI5W6tFFOWMytTdplLU6/k/0gGuRtZy9mTEg0dxyxLi35f0O78H+LVGt1hga
hOutFKjpkPXVGimG35qt60XYR2AoFqsOCSdI3LDmxWAxH7KqJ8r0MQ7ZoZPI9j0N
tYDAmoZLOhrDiEVz6sL8NBJlJvZ1jvhn5sbcABxpBiIllUSc/cXl4PvgABXPFSM4
RfYAC0p6c7pvxXr3+lORIaz7txjKK2J2S61aaZRtQexpx1VaswA/bv8qOn5s066f
i8gO4ILIld3qRt1NkRBo4xMaaQ7eflKwREwhuoOnf+UlloLgS2P1n/jFnCKhy+qJ
9yZtp/FSAQDQ4AGC4ZgAGMaqJbjb5V8NP6QUDqW0COq78caBeBz9stgKXjAsK2oI
ocxA9QIaVczGTzyGXua13FmJ6/u7orYSPpEMLy6zHfRnPnKM9KKDBMlGA2vi8YBS
J/oiV64AePfL3RsO3sqY8KY13z00ORnSEVVlvgIqOm0Pfg8QmjQK+6AjZd+laZq0
G6i1qhY7ImITtnlkuoGFtGie8QyZBRhZcgNEPDf9dyY1s50BugLOB84Gkk+Fw1gs
DaHV18MGFq9BDv9LdBY/EaQMT/OrnvE1cnEZsh6MJXoYE1AGHvrr621V26bEG/PJ
Jc/rYUdKWhU25C4DiPGBRHbzVOaQHO+Bueto40xbJ4AyWHG7pXB/L4C7nS4Hp1MZ
oLwtaxCg+JtFPhmgoioDigOKAoKSSN+um59Tzh6p7ADTbTYOJi/g3E3w6GPnQzt0
WLP7ERFHaKUslHF1YiUOv1Eq8IvQhvNv/qLM7PI91+AqDNn3taA/FnaniA97hCXX
yJ7LLto0EXPD4wZdTtPGFT6mtqn8exSbo6um4dpwoY9nRjpJWsv4ODxFYBKKLNT2
BZSyadHa/sWtAukl0Tiu1umLiIj5ZrzbXJm8PIByhO8ZTeIfb5Fme667uVDkqULL
y+EUyIRmQ4J6Dl9Thw7nxcUCaG3IeYFUqr034g2tUg4Qu/DUE9QUf8TEZzbx71bI
UnPBhLMoIZgGlEsIpMsnNum0yI7wFIyrfx855fHb/WWR/HJRKwF3XXz3VMs+GVgI
W6yznQHAMSD4f0N30JggKbEVrEpM3TaslyuDGDgJRzSPiUBwpepKYlE1NdpXUlbg
v04dXGAJAeQYBpznbhVhzcv/YQaV/4VA9ESoNs2JcAKuSxYoHnSMPlcdfRWR0CPS
CxctGetGY2MZ9WiN20uz43YT+u1pmwafVBNk+BDNJPSZyxE17FeVV/GN9EZAXtAj
KgTG3Znk5r1JC3OZzb5XiCzBSekDxkiFBYGQHE7Y2VjpoHd0G6oNDl6Zv5Jdpy21
PoCunT2aGmm5Tckdoipc1uhbMAZAV01lHYzWwupWcaI1r8IqzZE09vSSjTi1wMxe
lk+TV4JZwRM5As9D272+fTGoFJ+Rg4oNNjm+S+WSyI7NMIVlIg/J3kq67qA6k6hG
ieb7KQ6S7Gu6QrEpPp8cpByNNKZ7x60L95CSifEw06SYinKKMXcE8UdE0UjfJKCB
FMQ4ThgK4gFGZXUubvpdM5LgcAtdp3A0c7zcElImHMLZJAK231IoItsexUGnS84W
GM2F6KGnJ31jT7SOwk77S08kMp/CwcRhh9+g/aHR3NpRcJUHeXLDljfbLWzcqqzP
CPzOZI2WjVdwt5FqcEj0H07fezW+kjGQyQifE3dgjLRKq1uJkkzOpWRD2ZBtCNVp
ZlZDK0aBRGXodWHReUZPYfVkvz2f97gbySSMAHnCBgkUkmaGbTjHsRyFXqUfQ5NO
pTTyWTqia4gWCy8bYtrK+cBtjfVKhhuqw0nBOgaYXi2Un06ZD4jwWoIxRFednf3k
uVxowELWb/eSK7TdACraFklHxbMmSFp3d+SIgd8PCXWaNTnXWqF4If9OmNjEFq/G
PSHwIDOGIDkSbeD21cDr5IoNNgTkuJ6HCr9mUpffcSnfN+1DyjNWVpk7oj8qK1QM
+rrCNMlTXocevUfeamxlk1bs6pqFxnZBRFaXMGBfgBUWkhPzeGeBuzNWVEO5QilS
U3Mei7gjYkKT7ZlF/98tdJhcjo8hzIwzvu580CaYZgxDgoXyVquLBlV/VCuI7i3F
d9Y/jurj4xCw2maSmuj0qH2LHhTfd3gTOI9GAoOo/faSUpiClJblwid7PmXMYgNK
3jtu3aqNlqECIkEFThTwt2CVjTg87yxCQmSjEkCRNVd/kQ7dXKtKFeaDYMzoFkxV
IessyiN7zK48GkVPkQTbuiC7BxVEIBXrt6h11s4A5GHt/3C70OSf1Gf+x9ucAyY4
z5Uotk7VAaFELaqbOegrHSDwyo/31K5Qlg/AtICCK3eGxa6SH2BpNBJi4my3eKxp
O6vXKuvOJw5tlwuQf20L6oaWuuMBL5Czg/zbKgD0Cr51byMUq1yfVmWqyKQkrNQB
kblosGm98EKNMt6eetjlrbESR1+lgXXDusou2dWsXjr5Cz/8NsL5hTznkIwXYO2W
kDKE1ZfU/LTVcW5SgQcj/DYqRaqwuu9F4AC5jrqHos3JG6ErBIfDz/T+UqRVLKZ0
z/ia3c1Sa9x7yBmCHpXRBMVs+vkshr/gvb/1k14vb0xc57RHXFCWHpKhwxxRjZmk
XUpUsV/eeUMM3WG5MwmUHKoJFfAiJE8AHP+uxDarS+F2Gs5hEvyK0KJcfMogSDrY
0Dxpp2kzUVygCl3Ca+KdA1ybERwx7WXf75G+tChB432cKDdd06JMj47voTN3jf/U
bCNreFJOKiiSa1k7N/CsuQxIRj6T/YBhi1k6wWbVnH1UvNHRtg0dhMCOt2qNdvw8
4jPN+gGfRNJk3aXWOw/vlDOWwzMTycBj4AWu64vQxlT1BKnJCYs7FwZBpHne0wjL
d2GHc5Ch95UtV/3x1G9XvQlG2xQZT36v1NB1GYtInJm7MDjmimtRvy17NdBC+5tX
AgoB1U5eMLTIGoTENbQ0UaqBiNQXS/8LMa/gF1YSiIdDQJf5bLlRBp02W4t4qSPZ
LrQzmt1gTcn39BUEUVWw1p0bnUm7i8J/LyKHQOAv2pJiWU1nchvM+0hXWK7/8F3q
KYdOPQU1L5a5WDVjG84TTKwLckmJcvzEZym7x+OP+yCK4YClLIwTPn7GsMyST3gD
j5LUq6ltQnWIENogLiNym0tXFL8LqmKcs/SA4jNiASUlFuSDW9CirbzJEw2Rd44F
Q+7VjPrmVkPkbc80QANeD6NtXf4TBibe3djHaO2B60xaLcQjcuraOAyLFfqYXlww
9d6WB4UBDwZuBSTNfY6MBzbB25RGQboR32S3ecXBgd79PAduQoz8VV3A2HzGUsVT
MwEslF+IpV9JPmCdrnadePqFdKxSmeOL7LvuIB4rQ9nIyX/XV5MW7o6q8PFrXkgy
WUBDthCKnXjeWJvyw/gQ62RlUOfS2ppblTgKLTTqV2Dx7vRF4jppd3Dywsr8ulqf
u3cqBSjEmZm/dOxFRTB6wel+SfZBbVzPtZcJeas7FflslTR9E8/AE6QnZvRGBP4i
1aJbVSfoA5T1/eYQHd6kyQGLSKzmerpNyo5RmKhZ2cQcBL8rQtv6ir14Q1gSLhcw
tsxfyDacMQnnUYIvNOMaPwVQ6dNukK3KYZfgWRQwZ7ES+wXAcuqDYwVens5WPpPM
1u7b+8b9AdB2GgMTtZwsTY+QKAmfUf+5lBrt2htsdHeRrtBXsEqi4J4iShsqzAlV
IWkec/UClqrfFsRHM0fNxTVI4xuxU0daO8xpGJpwuJS6c774yjqhsLLSaCqqkSxr
04xUwyAV3s5ieGR6sOM4atqEqkqaRdtLH0pEW7Hvg3fHZ46HG9jG7oG08Ep3BwPY
kr63ktuSwCMq7DCVvyFg4bt52vdNrP+rqmCO7bO+OyUXYgBo5FzvAHmhlRerASAY
W02Y6h6qN3HCkGVFcCyVNFUlbagsUK12jiPk37zqmFA4/OPNDS6NPw8CeZwUinxo
NGPEn5XxIh3/JkPFlFU5KxnOmfOIuwI72pS+Tm1hzWfPOvYWQfK3J5WAm/bO5oAn
JFiQxouUnoo5Z0RzShS2yhhYVM4ivSs5fYfyRQA9zSp+jY+r4aTnbmVSBC/jHYJA
3LGzql77FV/nIB1bedvzg1hbFf1vcky6W45G7PesvdOdXbBsmB6wrLNpwz4be5mY
nmX0IsF7WhEZ3wZhfIsey4BPRF9tSw7HiJJotbateq8xveH0Qzlx5FSK9d2O2Hfc
xaCeTPN2hLBXR+CEA4FTmyrGPnbxlVkCfSMJ+05oxq4LhOeCDAQBO3CHLrG12aEX
PRUquxP+GIWrdEAgIHCgBSyVZMc+RX9nPLFEtCVRRD9eEjXaVFrnoLVDMMyrFLmk
sfHEQMX6qeNT0ar47Kz0kZP4+qZfvoNJk4C2m32NT0zCn91W2r3tQpzGB2J+/U7+
HUqd9GXIimqbzb3hPKMnDhAma4DFKC2Hy801H54YH1Q//RsJ7EHuO5PNLjqbo2Gt
SyiVCItrY8o/CEpvVP7JB8RTY5JWRy9DHoRqVDx0zAUnbYWzcnBFq0Y+gK/yKaXG
oS2N+K5pk6wqwPEL9Z4SDYET6+z5b/7YpHZz2G9YoOIZnCPc4gMYalztYyaPBSxt
WxFnZ/Z4XSu9BkegZ6gJOwCqnx30KtDGCI2Bjoqlf1icywLIicg2dNTgji/i3TjI
xr7s5aYaauQ3tBZf03uNRRlT7G+VOezy9O6qIyqL3xgHpVYSzWCh65iuC99BhBDl
x0VM4t3hPxSRQth2SS1sZjYBE0SitouFO0p0UsODrHxacj+hDtYRT23KgL4osi2R
gULncxtklVYdyD2nI8XbPYXhQBAm8jxyOjGfp5vFbXw0JMgV2F1eN6yqAod7f99N
xXnMm+xToQkzzWev5O0qCFgwUxWtdm4KZQ0W5gRqIzilPZe2IWD09/HCJnrqDSZc
unc/u59xh3oEqhGrWotqcLows1QjtHysZwOaI6r7HftvdFc9EOKLU9qs/bVC47Kx
8ChkXSO+L6inndOvtAf4u8PDRU35gfllURv6sf+cRNE5kFtjAUhuOzba6jIbk/2H
ToEvKUuaIxjEOpzVjQvYe3mxCpBF6an4Iw0bChCJemRNj/FvKHvCGPgg3t2C9Xwy
0+GgXtJHLWhc/++womkzZGCYwgbH9xudANt/Bh4mLkg9aYyjuxhDC59uiJOT5pLu
7RdFJUOyIOqwRDi+KfOm/FhjS/+OJ5FR7hBrkKdtv5LgkQVpIzmADzUB0XTIbXFE
4npLxdxDJgItnbVXxuXr+NAh8WZW8Hnk+pvGsFKELV8olr95jtGF015Xil6/cmQe
7bOlg7Xrk6mF/V63fE3lrH55LRxdxnYHN5xl6QBOdjWljW+WBeHY1Yp1ofWMW5kU
X/1AkhAC8pq8xdMdIKkyV3itb2HI2rGCjIaDLR9mkVddcILvxiPugMpEPd8EuZaO
+BsvxYRQlDPLV5FjUuI1BUrp24n94dbZYPeDZGz2/hQBRag7jg6R/rQh0QLoFpO1
3oUuvBhg15p9934ED0wwmMOkA2wV5Fftm1km+zbDU8wPK9xlRTIoxn9roFnf1y/t
xL3RvPGAxgrteMvLgkq6uekfnJb07HkaMpivavTk3K8Gh9f0y/z014nUILmlX/jQ
3RgV2snT0tnXDiF9XGyQ+E6cY0IvwX3KcQyM5riXtuiZurjO/Z1f0J2+UQRr3Kly
wh87fcDW0vJSvM9ZeBCU6Gj+zthJUPuH7JK2OF66meOHU78UUuC2Mnwzs06TdyLS
oebB45d4OjdHV5MeY2v9WJQhzqDMFTmBwDAycDTXNfTyowacLQJUKbJgjEvvKOmZ
QUWyr7ygZHOD0YqsXUugpxH/fNAYWfoBmgt0xFfRvGHt6q/CFFLmjaz3Lua5gbrI
jWnB7x92d78IDpUcz+kTPjaZEWlZhqRj1gD+YDHDZLc8rLe317eOV9u/eIwuZVI9
bJlchpXLaY/Feg5bargMaceSUMiIgkAPIRWetWn+45izol0SVgmv3/B9hsbAGQs8
wkduyy9wqcHZFEKrRnq/pHKDCU6VNYneGf+rAMTYkueI+SGnrNj/EKxO3NSfG+c5
6xslxjFrdLfqnOnXzkWa+jCS97BOYXFTeWJl36FZgALUGH/ebnDp7HXVHtH7mH3K
YYZjz+go3r1UoSwkj3Y2aPAFio9EIzyt4TmdIa1W4+y8Izha4w8P3knVNGrhXZk9
r8Pya6FGwu5z/uLS1u60kb/fD3+BgAdvJPv+A/JBFODdUB7QcDta7inONNqFf/HV
x3Vp8Q1bFjAfgfvus5DVIYzhCRLRqY2QBSkIWe9HsbHJ55m9/vehyT8yYl4NMalf
JiZm9Ot+SajjbLtlvS2WG18MV8Y649x+AQ4tNzwHt+hfudzMHvkgjxSec65wOWwH
oAOgvyIB+lz7y8oLM7gbDqByveqj4efGcGnwxSnY2GmzQK/Vja+LzJG6RsGvp/7n
smfgk7dJaQXR5qe6bOVUd7cAvYZPUHfQH+52mHw6YfliMM5TtR/EfmiFKmXyF4ju
eu9zbRcWEnIAy9UHAUDuUjNVbPIx7ki0v537YuyvQPB66zIUKgaFTGfVF5sjzXxS
hTmRbLaOfxJx7K7ms/jIikdHKxi7hE7ClVA1gV/123xV49DMvsFDUw9s6NEncRs8
zBnkcNZPoyuF4fFt8/TrF43q6F5h5ZXrtiF8KD1TTdUotaQakqgBd3QP5xYNjAAI
ARkNDPEALOUQ9EEkvv1Oc8mtLUbOCIvAUqJuKq5h3Da6wR/BykUXLNe4QzIfV7uG
Y2YEm074O42khjjVBl6SRO0Pm0jjtJJzxfZ/M2ClFAE85iFB7gV5zoKjmxxgF2LE
wfUUhlVgzIxqlncJ1tgJ5irfwg1LB5fr6e1aidG3Q/O9tLzZeNGTPSx8iZ2XGy3M
blj5UB9k1/IR89r7heYALoyjbJ/XXf4PF8oz+ukRWVENG2mOaQeK0Htgw8VCwlKi
ZmU4SnM8tgaJ3i8+rOPegR1nkFGg+uz72CtWAo8lSrD648uYQ+cNFi27Zo5U1lu2
/RlhiofUY51vLceu+QVn2kHQg/KtDobmE0HHDRz2dOL5RBiJv5GprzkaIaECj59v
qqT2zyi9UQHrCf/XUADoiw9afRJCxE9lQox/sEljm6bW7lECVWwlFTRhWM6or/LX
r6EfZHcRYdBCbpllR41SAFtIGyPDDVIn7MNz1rJNjG8DnvgaD8sV6zt9ECZTzH+Q
1ZJV4DlgmBO3LWzquDi12RP5go1yWpsybROQn4ugW36g/5wRXtY1fErZ2ZUjgvwm
5g0VuDmj1Z/M3pEF9Tap+HFvSmjhLiJoYMJp/TxPZkYmh+Rq3vWd7wR1EkPqqn5j
m6x7l+vx5ra/4waqhlVWIXBHr+htj/yttPaFkLctlBFjwsu1tsZ21R7/sG8Z04fM
OZQC/mtvigr+O8G4nG+qeOqGQJinDagJa/zwEQLYFilPwcMgLF5s7bgdUsoNr7a7
0sP4Mvwnjm6NT5Li2zlljwH9S3yImuE2uPxJiy7pIrQ8A5u2ovECRs6mdGsjyONl
ZNwOjWjEWOCKPmvLB64dNcf/n/K5Yhh4VSZekUp/GA1zunutJMAnPUsrmgg+rruf
8OLfVXiaD7VnESWGxwpy2tA/VkjRvxlwc055z7HB+Sd9Zk9GqwBl3NoqiG2eL3Ei
SNiyJ8nEJt8xWpKrOFQqwe900UaM5ZnRMjvrjrZ1Not1+Z2nV4r5UumR3zciJ5JD
Do41n8BvId3QJNsreUqZVJ4jTfXLMT8zbg5zHQAoQoG1l3/eioQU5SQrr54rWXBv
ErnLvpsxLqthusX01wm0isha+sxrgTGxwfrcrMGGDFWzTcMP6B7Kr7gtfiwc5Pf7
Rg+zTzS/WvKBWYTmSspMrWdSwXQt7kal6jIwHCDoj/aTlB82iUfRGyncwJxY1OE2
bNgindbtBWhP8SJ7ZPNDQmrwov4cW5VYawPGxYXnFfsRr5RZ4GBn/1bQmAtNd0xg
lhCz+6xtG0V2+SIHvgthFQacg6UruQ0vefqy4sePiESmJFPfpLc45GoDq0VmBUza
Q7NiomAbQJfh5FEEcC8Mra2PLVW5wXBpxutt2LofO9TyAPmVRHJwrl+B0YE8Q3ET
vgMtnHEx15HsmZB8J/vX1byJ1OLDnWNGpDHoYEE24lpsbZ7GWq6NnW/09dkeKRUr
cJ5civKIiFqdWhRW/p4IkFplrS8QJuMjNZmaTWfS18iJ4L4djcC8nZZD3FdJdbLW
7BIt6F67CNonKbINj/84/a3sMYDfI2wahrPpnNowJbYjREjagoz7k2e7Gd/RpEaf
igXXz8afau0tYtd+Q60frmCP5+En90q92qgyfLlP5BFo7P2ND/4Ua/bdFIenyslu
OKo3imfZn0BBX4l6KnwtDrIbfbnXe42Fi3AyVOrptSepD79+//vh2jK+Kgur4aVn
gWq8ms0649G3t0O2QSxTeym1wx8cJaTn4ghQUXxpfzLXdDtF4f5Zd6MqO5BYFdhk
Ke3yzb9E9e5YaGAUtrsNPrPv1kDuwW7WJeQ6XDX0hr/9U6h9R3G/B72yh3MshPlx
l3zvroWupenYOqYbClS+esM3c7KkKeKP6a6/gIgAE7VVcgW7S+ER/zHXbA9a2Yli
DsDQbmItktVmD3jM+HU5WIo4u5r2C+IJx3FgJhN/ac84UaXbF6XHpuSfQqKL0yt3
xqUWgZ+sObxdtbsaO2rTOTpjKbCsYuo7ztroYStPfQCwLX6rp87EAjIrHw1DxotB
Z4Q9rg/obdqjr4ngfUttgwyObmEFGuKrJg9FFqKCUJI46X3aykBtY60Dndp+4dpm
zvf428Af41Yea7AkM+YAztENwZVmOv0H1y5YmNYpFMYuPtig4degyQ1+jjvZyihv
WUN3jty5k6JlkgM1qhEHqhLbo24ApLGrQAONc8fMI/kgMUREIj0y2dVzrJ1waHrJ
UXxya0byAZ9eBIHnCeMfoaLeSTNgsn5OZycw3ji4NQVIcMEkd+mT/fA0NOBCho+D
gUSXghzxoM1SNjKeAFDF7xKtOfKodO4mTAMGyO28EgAUOIlbjqX2e2PwCYDVhMgr
/wUCa9huV3omaiGCwz1nQeqOFcqY3H8+o3qXUi+OqtR32VWIsFgnqgYPVehetI9D
E0QpSjLGipuxB6GnQP6oKKfVDu2wQbT2EUBcSoxel/1PwK3PgbYmgtVKn269eEfL
mJbzHd5YvGvnGyI6Lyanqwu3AJ36Ou8HRjjFGjR+ksy2m0PymGGd3yUIhl2TxNcT
+z+SOQsvGWdxoU0R3YtWpY0Z1nYio20cXYDknYd2H8bgjvYXA3uZklqzZ2eryu6a
2BqkB4iQybDV/abL8jYt1gzLVog742hTcL2RLJjLtJDvbaxvZSMcKwX4qpGO1ey3
apLWRBu3FLvCJXLqjoW3guqF9N9M6tRN1bGGgQ4+n2sOjl4qa6XXeL7CS9m5nx5D
WDle2Ht99jH2yatxOSSrk2oFr/AtSzGzRRsK6/UXjE5ABupDGbP5GWV13Ug8rI1A
skwidTkwWHdJy3cMUoj+nP02wao5zO09zS0+0rTsMtxHOYybNYGMNHNS1s7tH8fP
XS0EyJ4i5JObGJYH2+EXaD6jOUdDQpgSBO0LhzXk6qUOib7TglKCTkz1aVonD73r
bqYYnL2lWfJkmQmRwvtnrRK+UrMM47ZQ3o+8rnnQXDS6hrPbIw/gpfZ8lKAohoir
QAIrFHzotKp2KLi23XaVliyUrXpWWM/kCB9pGdD4uJ1xnxLj+Rt9VqUKFP/Or8Bq
nUF+09A2C9j1uizqEj5C6qbIDmkuOobDinULREVQkBgxBWE7dM6IB1zOfdupR5bF
vSGk/6Qfd5CCKX3My+o1iOyjMPbEpmqcAjkJcRVoSOFCwCmOp3QZTwhkVbIiiWxB
FRUJ+4eaIlHgelRF3icOKgbanerQIHYDjd71T5Wd2Y2lQ8tTgyxdKUZID0mr3hjG
AVUtHf3wpxMm9gQF2Q8nqjdiNpDJWe9c4JRmMFwAa8Omzva0ohsh3U5FmQ5g5wiN
CacWY+pWZBK7Cf2twqzlsoAtlPMAJ4HiIzqdL0AG6T1ku9dCCfh/RJ+JUePeye9/
HecYXQ7JGBca1HVfANuLgrA40qMyFAs2je79wKk6i2KDR792SSSwlp1Me89g1IsC
3GR61J9TGn5wv/I0s4OK+ihI55C8xzFjqNTTz/mN9UUvRgex9nzuFkJiW6POPiDi
ZUnDImTf9cIwT+eGVBd/aa923szTPi/65pcKs6pr3hHCegWhIhnUvBRDFBPh9XzT
vAVr4WpUJyJujHuSQs5zrHfbGV/21ojy3I7rdfEa86s/AMQJ2enH+FzRT8ITABAF
YzwcAiDj+j2pbMU/LJEROgbJv7TPxLWYI1VWryMj97XE5GKZuJZRHG1dDjGzCFx7
7Wjez2e5nYpKPfSIQFPBniZBKAmwMHnBmfSB4Pfv47eIWFOEdYyrjvP9Q3SE5dzd
0welWbC/Kfp9GCAqRaLyLuI1m3xlONCwqYKTrEODLqcsaWnjOI2TnWsaFj+h6fZk
xr6b86HlM2POWQ12yh4RHwrN0nnIb392BixT9KrlQf1dBJBA6dRXFYsoudQT7RWG
Wh+v4o4ma+xXYYqWfOKaDVvwXM3Zuplo9Vuz9c6wYOv/Sw+m70eKIaGGUBC5zsUS
5ni7Ld/FY1DPFVO4nxbr1WIJcGZXBOo12I82+u/hWsyCJB3NKa+rHJFOoxqUn070
95y3X3MewIebPNOS8ZepExijq9p8kcrZkkJ3qoiKe0JseUyuOcgg6VSOz3uiHKEp
3yPyJale0tmBVsdrihivzirBOHSzBJ6At3DTWOm3XHm91/J06o8y3YdjXTXW1WcC
4KXc04lYRYQ8aeyvqMn0gCgeXJTen5NoQEQZ2MsXBQCnla2aICFu747oaR6nrjV6
4z+1huwXovpZw2yYulwbzl29QtEtxLiIWbxNYEkCeUxFJjQfTRNjdInKLWdIfjsJ
oezhIwF8pO03ISje2BvMyzM/9h+0Mbk4Z4efehWUDTVp9BDAr8v88tESSAk2imrs
6iKeKM/TVYMmDJ/IKkdCqrJiaYFZByVbVYrcYvnlMlOC4a0i9PAITGShueM6V3gB
I/UZss6QjYBQ88poiOepJu2amcC23xWI0q1ci+3HCIL1ORPckkcsYojzKE+oihZE
p5qD0yd/OEZNO4JE7RZUPFXdmxXYb0gkqMVAIsw5iOh5lXNvcU5lbUzttWb6Oj2s
FNfmsbyDH/biyGaKUVNusmdQgRvFkcibkTvqBrw2WKzw65n3kbBht3vyqT+prkQ1
sK11jn86DkO3NG8ry8jvV+DBrRcM7lMj+Q51460nNyAIKjzZfrPX2bdVCfbJxssq
KfwjNGed7ohlf9hOGMGcPjq7R6pUxzRTS/Zoz6P1QfkwgF8eFn8J56KiiTYS43fd
Sbd1oCG/0Rn9y9IwrUMjGJ7EDIpLlGXKs0ACbnOaZqIZmqlieNhUnXCIXj5g9ull
7vFDjbugqifxhCv+V5DXlhTjD4zxMCvaXstpOqERyzo4kLw+QeIYPHW7+/ydffD8
IfpUUUZdYbSkkWwbCuJJzW4+VCvA2CD90dUP1dSfIPG7I7cR+munS43ya3m+Jm+D
8z+TAdS67DusYfw8H+8ImKu3AHTvddmCell8IZj9ezCia5oNeINU5vFISxzRtjbK
LrzSTsCD2xkxfr8GE2Mf5btUZ77aytQ4km74EbKvXxvCBfXkyewKNPZWv0kAIcAn
UnMWAPqvrjjtJ+7MGdlxG79urTCx5NBeMnWolMOJD1kXG8N2s6zMDXt5xKFMr4I+
bmqz9bC0IKki8T8yrSL2oLb3+dFz/xXpRV7hI4zWIvGTsbo87zPC5UStPI5sUNgX
CbnGxZRmiBoUEkWDOVgPgUQW4YMU0uYktjGaSjpY/puvo/9Xh82TAPQwt7VdVUWJ
bamzqnDKTNfDtzXV9pFzOAxaSEBPgY2vAAbxnAFHJ+9wrnvU2PAKlBFHvpJki6eO
xXR2Rp1zVy213H+U17FC/wWE1hoURN8Vkec+e1HKpLn+0wOT6X0Mc2o9nr0wiDhQ
cUZkaM5n+gDSWSsSOEb+6eRkjx02b3CaFBdtEOwr8K5qKBNlV6tc/OKFIioodMNu
fBLGwJP2QOLlflDtxqyf4aqidHFCI8QBM6P4KhZmP9OO7WkTUbaG40PATbXzI1Gb
HS2I/hBJ7RJtmGqY0hWnt9nKacfLB5iZnq9OqEXDbvHZk+GhZmftnDkG7uig9ple
FgBAiS+pjDy9oXYRGvE1JcTDNXQjYeICVh3KO3Zr8LzC8cResQnNIsVF6nySyYRT
7anVsvIOUunC7aUtUJNSkN8dvPPrie7e+SMO1L8EZCzTOtEErfFPODaQ+aAZIshu
XDCSZbdFmQ20nHqKU3vPhw5MCuivvHpR44RFKALDbUWUmzY+h7VTcXSnJYtqwFoL
I0amKv50vAf/kxyj/com3YWOlEsEdJr8rBzXb4YXrDcCdROGsddWj1zCTt0d/Dr0
0MzDkZtSuBE4zluZpbp2XdS5/xJkHuXgUYOaGIhj17SrQDG0SknoWhvOhtH2QOmf
fDWq82iEvaPk955DLTqI3SjJRVnkKvTrIUNasMrMU4rcIKG2gVtE4FQgZ829K+yQ
DfQ5GN6F189FRWkIsa3Zt5G/Svz6dIumnb/TfaOCh7B6hRCr1+SMgwZByU4GmsKh
7caliEdmj6Jz3xMssBzhjcgEiU/moGmBRi/9p7Qpvw6DSVxWxzGn14YD/ao2IpTq
ddLo+IfRGUpOcRmVslYNeqSCJnvDkV8TDjkzwB6KCmrJbgWTMpJRBoCrOBA4H9Tc
P0MAqPYZaL2CrmSo+yKKwnLoqiw+2igNl0q+km8RppH2Vd3LnfAxa73b0R7xSncS
iTgadyZjf9RPuRvzlcjiGR95MC6gmZAM0a1jAI/QP4fpa4JY/M8f/1kG7XKHuWaq
+5/Qv8i5Gj0Ju5hHskDLJtQWNIs9SMsHHO350Ls6pKtJnEMwhu3VxrRXuDEElocp
LIaHkPb7i+Wm35thUNH5nbAVnC9RVcarZZraVFcmSb89F9cy8ILjrSmjZXwBTi4I
zqKWuyek6mZ+rmUhPqOi3DrFPqGDT+SuKuEIjLBZ2Q5kPZwaZvhxJCZYEME2MXY6
5GamwVJvDlOz6SQOUURSLoia73kvlYTAqoMWbd+UII9bV2Z6dj+j8HCX9uiINpM+
QsILvXaaXvT7ukA3S2I2SyNuATHvCY7VnNgFMRwvM1AmlUEMu3q/VB6hytajNAA8
UWPO2B8BnIgp+idXWjnIAS+xFKw7cF74yCmT5frQxp+rJoOHF5P1FyYOD4xQ4SGa
OFfnZgV2AyxyKmLfoKfCmGfQtWz3esDhhHoARBYeY0tyLwLU394e7BDM2YDDTxMg
rht+8BZeNEWJDAG01wp1TrF7cv+Yw6ZQp6gQ2rMiubA2z6pIa5dzBACDhLpJ8bja
Ig8C+iCwAck1slpYcmRs9da1exDdgYQxpwInw//4pU2S6UnCjDa+YmmJA1UtTHB1
Kgm2oYUsIpgn0466FrzvF5CaSCaxqc8duCdY04uXu+q3BX9BdEQjrHHfUdt+gnzX
IV4lxT4Bh0h0RiTsmsEzLNxBa7lYvhl+kzA9pZhW1lIyrFtAonKHLEpwhZG4hKLb
7mM4uWEwIDuWjHpf+PDbMDgq0jhahyNdWdWhEfqKwnWm0FwfjeARnTqXlWE88m0n
ayjIB/3lvHuLaVVvfOJwFEzEqxpKv+W9iv7gq69Hq/D3wRl7S90nyW6byuFR3sEI
ApuwVs04Np3H39AlWrfM82V7NQ+B7sjNc0l87XQIHqW9jHhBNVnMOBMoE7Xk7dzu
BLTUrlFlodWlzk8jO1tphFZ1v0yx67q0tMGrb94XDPvTZc68JhUfqKDEdljINDMp
SdThFkj+JfueFjdaj9KHs5v7oCLpK4leVmDsjZi6zNuhdryR3l19705x+immtGHy
kYg+tCwcen0w5QUyOiD5wmLR6Cfgmv4MxX1/AkGASu37qEsJixbaH+odk2lMBvJz
8W9cQYy0fu94JrQHDw3Lbzuwho6hwe+krASTJ2Ltj+sllEQ4E4eUPxAFdlPA6bCh
QdP9kz9r/RZIL3sIOfsbnDo45yCV93dafcbgIvBKiD2n1/YROldqjIIMGVNkN7bP
zscnDACy+jZpY2v1Q3RcfKhpFtj5n2wUm+ns+y3xqnoGZvXZhH8Ylq+KqoibDGay
nGxf0cJWKbEw7AqIQkKGyKjIpURcXaxEzkw+hkqp0I4QaYvwXOGWlaXn0zTJ5qld
CmGb1lceMWZmtQ7VtHM2HrbpMhSPZCFSkqeBGEJOfJrrm+88WQGPRmDZHK4AiTYn
nU/YjJTFd9CDVW7riL01CN5pBjvqqzBfDJgyrGkpLQAa92W+fzXwW2n6saxraMCq
jBgaMUmHn1UA7XrQRzhfTyZGf7jQ84vG8BTeoTV+pDHyebm0aeXlO6D4yo0r5/u0
QMZecsx4YgfChQsB4NSSenQYDo9L6ikLM9tM60zfEPAh8KKa6V5bH0j7H7PFfnGR
0EIyDVTC+KrnZBB3/OCD77d0V0+4hxa3Hdlrk8bEE1sbAbsCxPYYFbBSf+6+M2dK
s/EUO24/vN/LL0/zsxwupHM7ncVQtsQS1QrS6r3plFGWdtiJ8J2KT6mFFEbN2+ZA
GYUFIjaNiz03E2nOoqtrdtCiPdutojic5qJlUc240Qu5LwqO9ZMD+zzmzpoc/+QW
bpV5gc0knNdbo+fLqiOehFnDlAEoucK/FoBMJ1Ops/tT/NyqLv4FOzptqmSxkWc5
pkChBGzJXsd6IoT26r05FIiu65jyZzUqcYcEG/f1t8BpMjxnkKUudJDkbOPjghSs
mVyfXjm8nko9ud/g5jjzsRLolgPngsOBJspTjFMPjsBzO/W5li3yRgrG4ZWafBiM
O+GjGyUNDpgSQ/tWNpqzFibCklB7rYR5Bg+vVzzx03i6MM0RiCppCPRYCwjI3WtQ
sc/MpAKg+ZSZKLRIsY2Ov8rIjMWH7lvL5L4X/5x9PrIabgVgBdtI1SfnmqNUYNUJ
YSgf+TEzAblVcfhb1vrQZqjZrWuNuOaxGb+/+vv34x/D773ucVx3+qnhxzFniJkG
rv/SkCBc6ghJo8GxOt8S1SBM3r62d6om2skBBxdlEqTP2A9OjYbilJ4afxsibFpI
BVMqjerz8dwZMawR6N3GPECLB1Kg+keO4gsYOTiTvyhTqkuAsCiij51QVV5LXIJa
rAvGxGGhc8L7b/sL7hnB2Ef4WX9mJWFQ7P00y4YuBc/ItaE3YzTJmeuFnuFyIlFA
UQI52iKuSPbL/yoRV6T9TZwzyiAmw1TCd0/jFXGhu8W6X6Zu4vqq0PgKID3BwflJ
VEm7BwYUKgNtlSxFEAIHXUIfN+cPyC/FYZZWeVniDF/MyZokmDIoYsSFyF9lBrIH
zRYBPDDbm2XsMeLW+Z005qeg7LfO/+0trYM97lxRTFqMCU614yxGQQkLX7y7gh8U
CCLPAd+GwK6mHwJY5gt4FUU2XnNtIaLYuQ8Ee/YqsQg1GrDCUI+2qZ6VQUPpOurV
ZIXea8sOQcOKlOKTvVnVHVTzzHL58lpzWiMUGOyc4J1WZr4RM+pNq10B6m9++4Y/
S+/4abbN3swRDDjxwelA88viefoHRAzTJFXC0nJRc9qk5ndJm3O2VG+XfVb5xKMn
GzO7dtJaYKJ3K/QapID6wyBYCeYexYcly8twnO4P8KUIDOblFOopw1DIQvNs/d71
entMIHolcqemKJVe3ZcsSn4unwKuW5avc4ZSxcfYoLUKV5bHtTxyBm5bcQERJNpx
hXQTs9L9wMsIYLxoujjEdzyiy/n25XCgeilRHtpghNyg9LHUGt7iMsBhGwsLf61B
PmpcRI1wCK9q2E5XWBGqHrhw5qKAwXTW/JU+fKJDd6Jn5qUk5XFdxkLsiSYpU3tW
Bi4fCv6rnj7LrDpNfnG5gKK6tM7tL8Hi50D0Vq429VXn3aFlEj/ocffb7Qvp3yLU
Fsujy4eZV5iItTM6HRJSMCUXcQBaYhOf4ovx4tP621LHfFA87uIgLCbvRMhNAQ3s
YTnUYcGlPA2iYMIJIQ+ABio1NLKS5FzEIb7u259uAURUgRCxvyCtg1F2OJy0Y2U9
8UeZG+pBvgbTzZSNeb9wh5y+iJCmNBxAEV/WblwPhAZ1adpo/2xXIX3RMYcRujTT
1D7mi+4S+wvtZ2VoYOCT9khhSspujgnnMJ6bai9sEucclSpt4EMT8LYFSrWME4wn
SxIH308qTZz/j2/4hKP2XW8wIqQbj6OkELU+QgNekptTfigbnHNagWxbAqf34R+l
IwyQr6UmHz2YcRVP3WS3Y+AeD26vVCa0CUdjEjiajv+5QuXx3yG/G+0yx/mI7tdX
jCj08qpUeaN/Cy3X5ESuvnsHgEpSsG/aRPbujSnv8pa83wVOMLacuTVgDwfXPrDy
+CAND5WIM4hiIXeqlkzMW5MaBCAXfvNiX9kSITDLRLo16gKHJ9I2Stk96pPDGt2O
LcmMa/uW8OkHcpuANbhFze/ug/RsCmJPzKxWohSqiO32gi+llfIHXj5pFzZYI7AF
ZPpU2KKnAPG4LF2YECWGn/iz/v1rHYggA2ltzTCPgNBdSeG5oSanlELxnedVssCd
/Ex/yOb0sG1aoTvzmXBMYsEWU1PSUPqE1dTA1gYS1I4A5Pl3rejy00jSXo+Q6awR
Etg20ZPyijjuwgWCsyJ6SfJ8unxRohpuapxZE90n8MLq9hEOYZHuyaYHyzNFBcTM
dbVj9IiD06b6N915hUaFS0/MKlsPNqlBt0JFdHYSkbjYdBd5rSbYbG7JoqQeYg9T
OZ34MKFAW+eoHEIwMYJjNsnnrWiPn7nY5bG7f58kNrwjwoGr8kHtF8+VpYac0JUj
+4ndSkbF7vE8HvC1M2Ayl+esJFk5GbavNJdUVt3Ku9c1Jv7qtTXUbbDSIrclYp2+
6I8vxPlHVPv/TozqW0T/UO/hj7y/EzhFQADpoIem0J8NuxnOipnfMVuByjrePMhT
SQQWnyCOdQuv2aNCWdiG33q6bLuwEJTooGG7jvG1vyj7wqr34G27t57Y+CDFu4BI
QvpYiCE2vVgpHqqaOXSGAKh+WzfL5pBPio0UWwZekC/Xez23n6MrMBSHob5pFKXc
rmHgxHzdBBmho/HS/NkbFFOjJvZhBwQzb/C4NxPRitPVeu3guZsW42Z4Es+63A4x
+J1t0Mfz8j/zH/+XQmtAzWucAwFmNUtgVXUVr26D0lgUTqffJ3ybWlA4Oy1PlDr8
qbTcga9r/jw4Lnia8S6NiD0wAmP+YddKXp+tTje+389I/ViwxdQ6xGUX2IsM9pI2
J2fD6uUapVOUAD7MtBHcZF41YWvalrHIqvxvU4f2v3lFkp7OF+Qsq5TFMBOk9p/V
txV8VxaYpCLBVIxYbHQQc6awHWPpjSLClYjbRM0L70zay3KbsqD5xtD7bm944/G6
1CTnBAuehhbpIfUAd26nkikbb0ryzSasRhcwA+eRBP2B42Dxw+hxsnGer2lGB1DX
AC7IBh6c4girrZNJzvxIdhB0dUON3R5E9d27J7V9OWKQJW8jTRb/U3jupigia7P0
wLmWDAp4HIDV5pqJPBFX7N6U0IYkQJqAhhmYqgr8x63VLf6IA7Z/vVCK90wdc50c
mi3u1pYo/INqCgJzRXe+cRF8NGsudJIdvnH348pVguxspZz9B5bkWOvyR/h4Y+mI
BgYu8mGpRyHVwUgxRQkDisvydvRVhRJaE2vPo2oXX+uKXwZlq3FCBvUgVdrh/dKi
FyYlKdvqaLeYT91vCFgOvq35YqvsnjRnnVrTgJj6ufWD8e5y3EYky6MX9C275YUU
4/8vD9jc9YgEPgE55NviVVARMGnsf1Kx1MXzcDpSBm6Es5oNygs1Kk2D0fbYy1mY
r7FuOB8NNSi+T4CzSDMHo34ZFetSOPsyWJmm6DlM+YsnozkFJOHcmjJjfIH5DLls
aO+lwhI+nrQXZrVgwuMKBgRs0fTH7zc3CUDKwm28I6qSZfA9rqE4RAystWhbtojX
z+yh7KjymR71lYkqCpLTiBJ7sx6INqnAfyu/0+OncwoD7TxZcumZ2PsiolyGTs13
gYISosQ7ep819b0Y/1Wo3T3GCvoceVrydILPMKhSCE6UQ6yrONCxvG9Tz1B966uv
fmH5Z5NCi5RYrwEXY3gQEAcZvPU0cC1kevez5PWfpWMx0srLBvvuxn018ZL/eFjD
WpBHg2eMEeDnzwZu5ciJ9pw/pUgI0QYlcwRrapo8gblRLCaeuZ2xq62sQyNnxApm
YFcM4gpGHHFb9tyPoOByExbvuN3w/Y+8G5P+EiLNnrSYrXvEqKsRjlzgnFpwQcho
vpquG8x/K3XDqKLPC0YNiAC81ksIImXgZ7IK+TCofpfrYHYoF6pA2feM1oOKOD/R
KcSvnPrXH9gmITGy2AFG9w2Bs5hifn6Aw1dZCRQSZY5EkyvvluNKJRq9eqSIM/lw
eoSZ38Fo56as9Q5fGpcRDnGdWRTZ0E3Rjl9InIW8oIsdHUvuvLC0vnB52OIdB8O8
8m3Qe52gzUIY1b/EHhEnA/57BdEFzZT4V5YtkIlCfc63ioeme/FW1+9GngJiRx2t
9sJ3mqWLaqAayv8MEjrdB83Z72gZLW+LO+tDEC07Wz1JmPKb++XNbF84UwTkR4JP
KEv8QBjOcPI82jxPLgTOtAs2afUo0ZLJkmlq0vpEdlyYckTl2AUVk4Ma0zl57tVt
m7PKZZXVR6pmBno+wxtICGO2hK0Aiyynd56K5sZCrEuSI+FN2EMIDcWqaXXozUQM
xdy+0h14/wv9Z7hsVxAUUOMh1hNkAAJyn2IuAKr11fBFo7MeXVOVbfSKCebHeQd6
QMq5nT9/EIcs4UtYwqn57PvnBX55RdJDbWXrNxhgGE1YtOAUyM6ijPXzOsluagzN
H5AK2ijjZW9em80soN8q4Up3foxd5J9o54hkqTdPOpJEBaITCNMswu5+C+7vvyRM
ULH+SI2B2x52mOs3iKpxzV9x2eW8NkKx4dTUHbEfi2K7r5SpZyIRZX7pP4/LbO66
8XazkZFmGMJeOZjIoRS9ycr3ERv2co5Ve0Yd+ntoPH5vQEo7VgSgLbCAJ5Ns7mEU
Q+XZroHa/4SVCJCksLZectR449UcCTyYXhNMIrtGMnG47IYirVg38Tgc8pGphmyw
fUeTZGukWaL9VIbKHkc+nywaWqSI03os4mowz37pxwM33msHTssb1i7tCYyoRbLW
9mA8HAnBXRU1PffAgaXSL7lBppgKRm+T5dnNQ+c6gV5uijwHlnwFyng9bCw8pfNI
6e1btYCTSEZFnLRKOBxVwGoVcGPr7+QG9pwX8x5QV0m5L/amMdU4P8BrOcrRsEbW
vvcNV7LkKbMQ5CFzyuK+9AkHhgwW4DBoiN507dxuXGlqc9v/wc93SolNo8v28n37
TTOsHdBaZRdXdhXSGiZnxAU6lm16Ok1OtkCAH8/hQJ6SLzcDR6KHrddcxs8yd+zx
iW0cBM7o47zk9tbtoj7JDXY8hyHMfIodb0zoD9+KjeD8VJsiDN24pJcfdbfPuKuA
AcDhvNZdMIIiVPP4QbMIYSjuCjtD7zfHUplvQA1vPyVPZ0Oz1uQpq+lFnX0NR+3W
2N2mW1z2yFUL8ZHkJWRHI7JgX7CQv+k0dOf6pharyUX4cve4grhGYH10mY8U9j7S
DuENOOsmYT78RfKpqFYizZSswhB8S94uo6uCOH1tLA0X6FzfS5XGU2aQxjIoUsSl
D/v1OZIe3UzpHe41pQuEybTigyXuhxtd/X8V3vyfMHBweoV8YSH8tTWnZHdGrs10
2A+QbbcNZbyZRsAV42pBqq5YrOpYtmVyygJypgcm1nlGPv+H3Rg6o1YgLicAnfLH
qh1h2QK5Y/S26PduKigxbrCANXyNA0dhBGEN1/obrCF8zeouBg3GuR/qNX3bg3BI
6x4DDQ2nv9ayh94AvzooWeugSLQXKYoOBDTqcB2TuCo9XmwVrQ4G4Ry69pbBTf25
SRbVVLhU7//zbD+xW6HDQ+sC2xO062SpkaM6iskbDDV9FEIT84JrvT/rhlzTPHsl
g9DoA5hsVAKY36izVKl6bqGbPYqDNZetTjL1JIya/jVbh+T0ZTXKx+wsqs5qyHx6
hDOUIyJ5ZH3llbE7c+9vgWPtNpwhhYiC4gB2JmCQ5aTJmMc3Vidd1iRtQb8ArY61
eN8hmX0hQpioHP3YVr7wghPFZslLmZOnEbKkz+Od/D59DTAp2eZ5Tvg8rOtl0k/f
8IQNELUabbgHereO8j3htIo0A0aErqgl9hds00QZfu/Xk/fTMFqouSp8rHAk74TJ
b6Bmi8RoyFsr12Sn6OYjZhuJ0O2ajlRLxJAxPjUtxB5r2ExCrHh5O8zTnaj6/ppM
4eashEtvDVOOQACSUkOc0Knopr/+QgNeaEKgSw6OcuqpEpfDO8ZUcdZkRTOawwNx
ekP4Mblk2WA/LC1QTlZfXcaBCyqPTGul/X/hzr6Tp8FOX6pVVoGFYOOfCvZ+JSd1
Gx1zkw/t/K8C64apyxKl58Onn6n5sgAPqzHmM2Xty32VGgwgt3ufNzJSlNCCvHAe
3OeVWGcSdPBe095JaJQv/76XLOdbiyfe+jiGjkA/XzTZX6hjHJFMGznxAnHuMwHB
YHgO6NY+CJ4510/LH6w+mzOGd4i25d1cjjld59G6eq0ZNVYJ4+cxU5GiME1G7S1L
LNQoiGHYSSyERTEroYeM1Mu82fDGlk0KHuPILbe5kY6GooM/dQKo4Bqap6lEZHFk
k38VllDaGPcnIK6rnjSO1Shy976F+/LfibrPxLNkolNGXcOM3Z/FqkZQATcDpdIu
k98kkMz0W+Uq2+lblp8iCDWSKvShjhBCfLgED9XZ1TFTOn+0uXxnMdJ97HGDwivs
mLN+faFft/tfVg0KK8j6N5c1r9FEzpcdNNFHcN46BOfkgB41h+WllHpwiB52AU8b
kCysrPHclrinsb9AO60bLj8p3lbhBqq1YVDKX1gUW+g22n/7Aya85esKfrELqg38
oErzklIoKl7B2JqrkfLBWnpCRxngWRXrz5bkUcvpyCa8p3wL7a/nA5ANM9kAEWzm
cDCWt4rHhL0DGsN//RuP14RkoegFSi3ATOs6Zso1sY5eKxIC4NelcC68GbQ5FBBB
7n13ULNU+qdillwsu7kwFk408I1gkbiUYI42OyiiR2l/POAhznE0EPSh+8nw2TOy
lk4LYW1nmtMgG2gHsBOLJDQ8xbvjs4yEU6igoZXLYwZs9/0cidwE25xMuu+q40Sb
E978OT7MhxdpHE6m76ETwJ30IDbPnAnxRsIFpJFqLWBhV/fov+ZcxYZFp7+v4KZV
HAYh1SSIvX3c5D2yp4oyAYQUEMcjdyZqtgmM//RGtP1BFAT3Nd2J1FAROLDdUhaL
DqLnbaAOU08oooiselwxZ/3/GLOHx8vvI5onifBftuVOSfj/n2r8ARfFGvqHp2iI
XBIDQxUydnKspQFpI3baA/Ngz8P1V09RNDXbT1yTBxwGnFgCNGpLMJJKMzOxYxqL
5bV9OY7PZUlOily3Y2g7oTr22IqfD/HBPHksS6e+E4NhkeMEWkbQlmkov4mBadIy
aVIbf+eonoafGEMn9WDKw/gmRkNC1bvoSbzAEZrsFQgMHe7xdRCS6wju2u333qL2
2ZRjh1D5DwNJxjx520rbB9bRu3poRm62Bt9dd7iEb/osrAOmSi+CLsyPYBzSRW93
jXOJU88BLm3AyjmJS6mWVL+EAbPau05AusJ44k8jVPnf0wFnL9RZ3ENGfrokodk4
Sae5T+mhY+mcJlQBECRnaEj/nZZryulMtZE3HmLBhw0WSYfJ9MevkCnSOckjE1mK
Ve0SNiYZ87ZS1+nkGmJZbNc+M7bIIZoL9mYHMUDFD4Pg3H/KBJQKdqfVEDa6P6hG
PzT61p4TJopyzs1javaiDfv5OYn15lo2EPE98UG4gZ/1RaGzLTupP2gdq0G+LLKe
CCrOLdM/wjAPgz/192NWZ32g7VdPNvoxJebGyBqzyTVdAoxS6r9KiHcbBIQkeExi
btzaJ25rMBDZ3untTvAnMZJBdSln4j/dSgjYRqyq9dyfpadCMLpDvQbaPFehzKBl
PrtXGB9ovn2dC8E+O78Dgmcb0ztwcJUCKa5ZRRtX2eHfRaVIB8C92vF9QTooAa5E
tn1QqWjf6A2slekRGh5qgm+L3IWWBs3jgS9TWAOWCzuuGNzwCpDuRQ7BlN8Q3O5P
7kHV7bdlgpMwdIDkUJPa61Oo9vYCKXF5TMicv4cPzPJH8yngPqrW4ogwUEgM1m/L
4UVihG+ajQ5HazVXbec/RdYyZ8UwO0RpOC9Gmf1SsutQCueulTk+jSG9kJD3mWrX
BtSS/sAPSMIiX3i4FIdwTS+dpBi0Vl5FkwgFh0O7TjBhZom9KPpbhF5u6trjghQR
JyMBlRW7NpT6ojs8v24tsBK2V1GF37/WcamEeC8DTgkbiPaMX44uXicVoS0cCGJD
2xqnk3H1brqQUYPillL6t7Eam0mjMf8wfFh/3PMs1x0jvimlVo0HL03V3OZPk1LY
LyStlyFIxHgwxWetOPh7HTKOAbRX4+9ip8pHZNQbySQlruQK2X3MKWNoem0AbNZz
X+wMe1+ZtxfNP2Cv4xUiY7fbzaFCKPyNVTV3Q+uMmZyU0oDsAbJHdqR6YwcVEwaU
OANqAdQr0PKrKLIdW8HPP4FNqJDlU8FQFJGq5CEgzanZlY+mqwmclMemrqFL81QB
owfwPQT3G21qbvuvHu9HkKYMg/c33N7hKf+SfkpSKkO41H2ood9b7nZ5aqBkJ2ot
QsKXLIAm7hZ/dJuXhPw8vaalbR5eRJKqcGfDTEFku6uHDKQG1ksLxUtZBRRXIRX6
A1rni0mM7TmuOQbjTYlVWxk5L9f0u3gKXfzHttaYaBsxomhDmmYW8q8uJH5xGUIN
EH+p3otq2YlHZtBXNIrum0NHMbddLz1IhlxRYMkzUbiCEqdfuA2Yy2FU79nqMkwY
yp/e+t5cbjaBa5h1wdPtLxuK28tcOes9dcKhFl702cUnMIkQdJ2UAaLmoVU4haf+
Sa9b2D85UrPy4LIIMJHuX+l5ZxLV/chR9qo0zq5awQ1LMRJPc6vF+umIAIjjHdaG
MW6OD+/+3KfuNtcUjOj6Nqxm07l4Ikeh/dCfZx+oCC7Y4nWYHrmC+2halr4Yqz2V
VdtQiM61z6dJYy/VCHeTZ4ZUBng4f6QSNBwciDxliPmpJZfqqjF60Y02GwacG6yk
DbRCrhe8q16aYjgHB4+Gcugchg9TSonirGHiKbtF8gAPSUN5aK87NkTe21npmrpf
/jD9zGcKimkjXDC9fyeH2R/g1eX+A+8xrrPKHpHuAZm23nfT4jfiyVsRKnLU0uZ5
2oep+FoFcFb11aptgb2bl8XBWURcp/V80DdejzWSeLLxb3XV60lepdu5hizVJTes
wSy1cfqL9NBQ9C2nvNmdsS9+WNNzaNtuS8rh2q26aX3f4lwE7hlhlCVdsHW+9J7G
fQp6/LK7931flIPTyhCQILC3vXdZXcYAY8mzbYiPNBcGF2I2h2E+Jw+7CPFw2AvE
x0Z0PRSdbdZmxbNmJs52IvJ99NpgIHQrZ4J0e3F58DB07cWu10t7od2+po29+geB
Q5G+mQ+iz7qqgxAiue9T0DxmQyPgJWTGTOzHnPYJ8NcAM+lRtU47DRSbZw4s5/CB
mgb8+pRjmY4MWVzdG1sByREZsAJzO4EmA/owyqzpa58qR3gQq9ggr49J2CPPz12d
YPmahMUShzj9MGYV+gsUz+RZjlypL6vCEsKmwqlcpUaMR8SwIo/5pQ/q46bI3UVy
LYEacF0R2uOHcLDeKVJj5J8cjXe/mD3SjM8zm2lMOvYOfnEo4rA2qkUa8zSZaekD
E0Xp/FNK8QX6yHNTmY8f7fvMmBhnVMThd0UyI6+zPtaM0YTSxes5RE12lCEM8fKq
TjtxwEhK/wi7lTq+QeFmFgWLC23P/BmAAJj0mDpcegv2/RJV7WZ2vQyy2aCa+6gW
lWIwmnDaDvRL5J4evmfwvu8wWWeM5rdPWXBAJKyAewePDjjNhAc8bIGAwNniduy+
UAIPfIVk1m/d7ULraKC23AA8HS9ko6/tbAlbXkulIK+69xkket1NjG0EfoBgVucx
3uPiG1z3lFmvXtvHwLq+P4GqspjzITsGi+V5tIAGyEjKg+RH9rnrn1frmbMDNFo8
gHoBdETF5oXNaoydZQpPiRZ+4s/8M14EpTqJu3pWpZt/PyeRD9OCmwMdWcFJw1cr
NbYvMlEmmMLYgNTPz4r1hgoH0b6mBWNVAiIC06DjFXas8Fr9jv3wt4b+InpF416o
t77vwykjbOyxqac8XiwyYyBLZy0hwGE+9q5sxC2brO4+yGEdy8jiZ1zClEcqffI+
+eka7VHgHZbdtHi9dOj3lCuBgzeVUhXpmKT3i/oc7wqEh1QGCfR9ukKqSLt3ZsDM
Ddwxp1rkIH7dAHQudHQYS2kVZN3PF27GF4VfPo7rqLerM35jZCThnzFvRsqJQbNp
9ty4bgyU2Z4q1ifxyR8TdOktbK7nNrhm1uic18t6w9rNMCU0iDQN9JcBJvuLVuP+
CJSDmrdeAig0U4GxvG0wdRDpmiFxQsU8xPmRDlSdLgiXbw/ZbPzHBLxQyLnxc5/Q
zGVYee86OMQhUUErUUfQpjj9eY7kiM5Nser1nP4VaTSpCKqkNGB/e8HQV8HMJMZY
Bqs29su9mSwGHUwmVHyGv9CVLkuh6e1lk3HFavypb2Gh1WSxo5iExYNTDIxEObLI
qJBp7MDaJIoXOdFVzCWmvGkUqK0LrbXRQSaslhxj4bf+biSsBPJY1IIK4Tj+db8Z
2XwGnZDxTZDSBdimzW4pZrBPLPRJZqi8hUXpzDB6FJe1/jYfMChZpmKhLWvlTAVK
sIJ6r82WpxhlYOPZhzEashbLl0AjH5z1akGSwndxaZLjzXdXAg/tIZmgPvNSgmSL
Af0Fll0G7RIwu0SJ5rTstQHT20Qa2WRoE17rvE2KlxCqML51dbFVr3cGJKGohtfF
sJ/IwC2DYGHq/XE6zdpytpgs+Vn2d9CLSDXvI0lIQeKO9zZ98J2DPJKEtpR94+nC
kKX6/ipe+i+a3fTqOAqNnqr2aKZb9I7hG0R1nTSj0sWwbx5Pkp5uFrvNmryxv3Nr
kKo4zHJhYyxpbn8pwoAgggebemgoHEBS/6oWcVYJyh9yTxFX6S4nyRczptavXld3
xF4kajpHHT+o3WCfc5dYTeC4lKfCaxBnO7J4OOt+LDFdB34xzYcjyz/JLlM48DNJ
mOF+T6As1pqf9WBsWz+6BIS7JJtwydNy1KsWHZDCqU16tWQDqsP6/fa81aID94Bf
BxDhLNfPRLZmV/5ouYVxUJWJs8Nt1psGfDNI+iakvOJSm6iZa8pPX53GGqN8TKK6
eL2O7vK2xH51hLL9hG4XeEqB7QerfYjTHUvEkKYbXyEEFb+JRHBOclkUnvvyiqsW
yzv95RgUXnsvYq19pqaPmxGXZWkjaY4hK1EMZhZVdxV1CPlpdZXMX5FX2xB3CKSd
RfQs3+l4AMPoViky26WUFIZQRQnL2n6pZ8vCPT88+QWH232ztgLELwbGRbDYtJTE
mAvP1ENJcrHuoO+T6H4jUrlrl6rQfYiNj/o2vxh8sgQs7TLaQlZluX4Q70I6yr32
sqK2EIibZMnNyct563ZSNv2OaGfYfnoFaAl9Q1zdfWj1cPnykx73rV64BxHmqadT
oGZ8T4JF1fzv6WhJLIAMs4lhMg17bD9BPLbl6fmm53CU6haAgIZx8OTLBtyZ0Z74
vrl9rtAnJ64CMQAfZUV5lQkjTtwFyPWiHFzZ685Acj6ApunLxPduqx4qpHnGqIHT
A2kE9buINzWMtOIeoYdzAcNjtPBPur4/l2x0QZZv1P98AYz40Ll9dxRQYQkMBbms
QhVGYBznPo7WB3rqlNsaGdlOb6ckNkvHAPTweNIUDxDZm3jy29Q4DvK+Ujp/RzTL
D0dobdOZpiVjgzSW8i5lQGGFXWtb9eUOf7I0q3uFce5TZAlWDpGP6KHCK7wOGG6I
YmZgYDwLv5n9NSUKbHitNGFHmxao8O4mV6dVJ8UPFX12wuVi4YlZr5l4BTUfSAsJ
8gX6P9W7LRM3gmvjBhQ0hvS5YDGXNwPZ2/hPccw3jJNIr/kpTsIiyVgTyfmdHAcz
nT6vJrbQHp2DUQGjNtBDXHiSbfoj0vcuYu6bumV+tN3H9/ddN8Qq35+AsxhEDra4
64jQYcCHG90OCU/muSEr0WcjLFkn6TJSIm867giBm4aEX5MhVSni7vtPfiBLrIEz
mGsATLP/fh2EQeu/qZFPY7nKiy2gj+uoMESgwOxWvmc0CfL9d+sJTmTVT7KV+PRI
eDqhWmJNnr5g4ebV/mmbJrpc2Atzziie5lrWGoY/vUdnCE6UHvz/ofOeC9Do8haO
BU1fze6xCOcfSyZMk73ZAJO0/rpMGoeb8TNweGkQiuvAZcjRqCPdzjOp87ozSagV
rAn4peGad0FQQvkJ5qNy8Qi7k/SWuzx/cRWlCXem4kYYUf2kADjGPBdiwJEDMom1
Xoi8lpYh4ZbySL3UtGnBagMmx5W3T0cWlN5chAtTmmC2amPyPJV9DLuFiP7DAndE
uUMIiB7cqivCRWMp4yDkVB9U6RYunuR8I6LUnnqNk5QbnPngrV5KJ9gaXPGcVbwS
Avk5R8IJ4QJ6vvJzP+ZwthD+AmKPee/dbvbSH7Fw9TWnh+NeHMjve0L7Bi6+NPJW
zudwjYRTzPXFFPcWqCT3vO99xILQFRXQhLLJjNbdnWUB6DtxIQ2lybkL+pVUaY0O
vD01MvX7Uh7jc8IEjOg8qwXD+g/K8/8jIEbffSkKXRoMhFHX8DRPXlW/hJlolh5d
yrHtBPzNAQyW2lkH9MrfEWl19S9tCOVVzyGwFFHl34QzFgfUKsu8tiXto9gixMr0
hY/llusFMK+QUYFP8rytpQ0rmFqkSkSMU1rq0abH4MjXXe9o8sU2IzqAvEqv23Fd
gsmyRP+M9xXh0aMdS0Siw287Mt0NQa9BAeI/0RU8n+2gcl2fDabAg7ToQEmNhCbZ
L9lImAHmmK5dmXoxGrQOZTWdcnea5GezlRasA2vonAd41Hmrjvzpyd07v3+GOTvE
V8r8MMFDVEefeLQlS4EM20hGmiY1ipUCK3hBOrLEAKZyh6cf/nvzr67IyB+K4c6b
F1eGNHHsw4MAfup7iwrseLgmB3zwXC7jB77soM/ukSiW5I7CsxKtibjXQoU87JDb
YeDfqdgec7PPbOX0lC0E1V0QwwyMph/6ZJY+yy3b3Dpzy8bs/VGrJqA0tEbgXe7L
RSxoMW4AjsHDBYJx5ImvekHOV4c5prdnVdtw3QqT/1fAOhm9fN/8Kw0lB9EnHJ2j
qz41zxUeMyMe3z2JEtPwwn34gv/Gn/BXNpPKbbixqg3BRBeckV1pmo4xVOUyX3kT
4H6lEqaVSiHl4CTShyXwT5sqgTGcnRHGMCsZTiue3rar23bMRZMfLaLF02ID6C9x
rvXVLe+gWk41LRm+DzXP9uoGnPqiP+sbYHeGhuEYpyZSik+goU4E3USYaEnGvCs2
hrF09+Quqax8+N7NWnnChDu3RLPlSAOoM6v/Ns30e1FgnH51G+xSWOCaUtds3yKX
/5gXpSwnTaD/ofhHmHBle//piHOQhqmzQRXgQMiCz/P9PDTQOyV6vG7qt/bWIdnM
2WnXOIC6HRLV55ohVijcjWy8QsmTb6Xi4mRfMTppeZt+hAdpXwckiOdogxcr9R32
amObyCf0UotOc9CVeAuWRbse97K+Kr1sdnObXq3OKJliGSPIOP0yUtoU2B+YLnp6
c3GO7q7s3aGB03CzTup8uhDzyVTNHCjpP8MLLqHDxJG6KjuGasw/bABx8OHs+Wkn
VnjGLdlQ1POyCCNCP0/xHjeKllPtGBJsquLr+o81jRyxgYfvP9EKH/ThFRz0BPo5
9jeN/MUgYH2IQc2ukjk+essnPYLd9p6/ecaq8VOPz9ur9v1ISeFfWt1+o05agq/t
KEiYF6aHRchAYJBchJ7ymlk+BwYjxe4jGgRkYtvmdUtvRUOdgS0tL/QQrwrFGxaS
zgEDCt/Ub+4AycwRJwDQ0/QetZMOli9AZSOoTm2phRH9mbI5Xsbf2BpWBRiQjhoR
+7QwB2eb5m88BZe9HrUu/zf/oCeWNFkIq0dZiSMvoZnxuWiORT3EcE/TNJTMGuN3
pUsb/cdGTvyzxmXr5E08SZlvyN+J3X4pLz+DGL89p1lpTPJuyFrLpxmc9C+uWUF4
WyHPGQmk8SduKd7lF7XqsS59H/ay9u/Xq7xGLXrNtf9DgMjygMe9WtJ4x5868wHF
36YZAoV330792GPrGWI9TpWhIMydjkSFvgmpqqnm5oYkNmm6aKgQ5J8QEPDdMmAU
XstU6QopMdvqd/Fww1PZniXbaKUfx+NYnuVyuOdq20ubUxNirnKD0UuhkgCENddS
CroIrtQUL3tbtNL9o1qDLX2T0vwXRi80mQrAa1NemJsy8y7avTm9K+Wzy2asqDID
6pi2L144meTvpUX3ya46uppB4aOuyxKCmmInIHgd5pomjqSHpcsIZi84CIA+eBKb
S4LnkgliDzXODV6cm03s/7FpXSgSxk6JATWqJROr7+aaGm6wQ72ujBK6TLaBH1kP
oMsml4qWYBjakl888I8dLJQSnjAgMlh/xf7zlGteIxSKpLYyqHbTkz/2QRQYW2/L
6P0NTYNy3Y8PNXcHqueWo2LFmw0deiwd+Oo7nTlQzuHgb9zk0Hp6VDXywNl6EZQ5
HG+MRtnd/KBWW4d/KkrUXbt2L7EoiGWKO9tq7LkULmwf37f17xmPf1vMhkVDuJIh
OIcDUBoj1QtWEal74Y/xjng528zv8OJ4+y83B+PmemLkGnVMTyVNoAsbHSb3/j2R
NRQtYMWon1COdICfpbI267+E7wr0/Mykq/+7Gsd20qGaCP9syHRBq5RTx/ZaN/Jm
5jjfYgn7x06PtQfgvu0ES9MjgDhOo5MHXna7cMuNaZ6F8egabjV8dVlQXDKN0Ro0
/3Hd6/MVdeqSIjilNQdURIipXSPlDQJvzYlIgZsiPhhaDc+rrJ8Kdp5vES4xPeDX
ZmLQm3yXCa0oL5PPWiC9ptc+ink42IOavdL7ZtIHIRvN9NppjRZT514Wb4EfGDV4
Y1wcMx9IKy0W1W6Ap2pEeSup8ZM12a/dn1AjAvPIzSwS/oQyjvtuYD3oUIeoWuzq
/hlP9oADhKNpe3V3+gY7+Zz45fmrjYqiH6kAZ+MslU9lZv23dy+4n2EbwKRYBc7F
pGQi1m179meZnuHeRNgN+T9SMhmlt0kwgV6W63d/WKuzjC0x+/B8GqKnJfITUMma
tnC7cFAPKqvZ9qlMhUfB3/rwEgNmNyXBeSYoiEcFy+HZ/yhE+71b4XP1ZDsk70pe
aI1FpdfgnkP5H64C9+vPWL4k9xi7DaqLQWdVm9oeXcPrNeX5HtEa6l1hoNGNFxA/
mWCysk6jBUqn7DAbbMzxlnTQQ7fw264k7ThGyRFK7kzw936zYD5tfea3nyS/Oh18
nPfNnmGLf/OqCy5nMagu+474LTAWoy4MqHq2F/ybGF9ATebrIm/Xt4a8zcL8ee2b
M1sbrBIVDeHQAX7rOswaWal9V5Io4m4N25DMI73+BKEWXDQ0aqQ8nC9YGYCCp//A
EXbBFp1A3laxxEdgZhxpmpDcU6PNtSgJqY0MDpWoJ0uripf6qc/3zVmakqPF3dV1
adTRlXAtba+Sm9j1V/DDzfN1kymssWR1Z612NBh0BVmPLP/eTNMan1P5zaz488N7
w2j4Uy68gdYwIXJ5uJSTu1x+mfHCkd6oaCrgo7J5nXVDvVuXfxLLzacyj2GJ/296
W2nLj1A96lulatELIG98bxqm1ZR4Y/xH7NKBaxTbhJf1ipwjq7mNOYMfC6aKwzig
9Jwv++zoH+dsaVCy34Wolryi1RE9VY0obUxF6K7gaMWki35Qv1JRIWAkveodm1vO
KZEtSzbrh+X+OqbvVZ2bx/gx9AUFdBDjlJKi7eJP4wLEjH7UkkDdj5TpyM9dSZi/
7+aeDjDZZdtBYIdON6Rx7YG+K/i3urgfZFNT1mHau9ZTGsI2TdNzYq8QPaD4ik51
KB/dErcc/usKwUr4UR/qjSTT5DiiBeCeZeJEZLf6opZLjkIV/LRqjvV3IYYIGNk7
2OgMCZ9Jb0Lz9fdl3HKMfir93sz/cIYLeMqK9h426UGbS7uDR0LJAs406EEqIysC
Czv+5Bg5F4TkP7PsX7Xeen6VFQrXcY7rZVQX6ilgPN4uAJ5BfecNNtP2eEcsBy98
B89N8O6Ghp8ix90o7A8szLUVGEfCeVrmUC/EP9hhTPOl2+knBfQp997rwFiz9oy4
S65zzUeEg719Uy/B6IeS0QlSwVvahN6IW4sJTYFsjnM9Np56T3bnVAyPvNNx4Gj4
lXuotlyQCOoECa5OGsLIP2/Uoco7Y2NFnbEQVt9AP7tQkyEO3ITlPhm91VgX9F2Q
VWqi9AmISvAjMpUwKEuuShx8qpwf5P1S6BKs0SozlgeBW1kKtvbjMGoQq+pv8ADQ
4q5jgGNuoPBf8kJKf1MQ3dvpQZUiqQ1FOPfjPp8phc23RNuAf1QJu9r5C18HnBkc
xCbXvG0oaFHvUh1n+go7YrPUnePe2dFtufh4spEcofp9aTF38IGWJfZHOwNQ5oVi
AqUZrX8nDlvhv4fZlZUzClmtlfeAtUQwge42XCR7r6oDgi/Qlsh8l8YTenh//KHj
PIcDDgWdVVYufGREEC7fkMPkO3u4CiY/Ki3CK49pC8db5zSDoXgPPhdMwguo64Mh
Mx53JakSNNoLFqyX/vVdLNxofjn0FULpI6lUrKwT0Z8ZTUj6A4FAYBtoWrBRV/rJ
s7DTBF9uUV21qf5I/MigIpfIXbBwyG2jcxiArZgefsFeNmvBJPkx+0AuselUC1R4
erZApuQtykacombPd3Hv9aTPfqDcGBDMoFx+H8nsDYTEWmW/lL32iwhnNExSfibY
Y09MeaQsETMh5J68EOP5v6E3gqGZHG9+3jFnSjMuSwgRBVuMSRCV2ahdxJ/05lU5
gmRlKQ7aCWcDguUiT196mWWoXfcFUH0fnOrlwi1JYsQEgVWD1G6bQWN934jw5j/1
6Bpify7A/GdVvzieI6MmHiilQsUPwQRlxoeG7N+JsYBNQKVe7bwo0/HkTvr3V2Yl
r6Muu8TBNZLdQyW3nyBHqr32T9Uyyx6otty2ZLVrpaxqiDWxNLIvyvGB4uo9+zUh
K6hNp1Qa0UNSgY3folQIolrcZUn3cIJtOX5KHqtH/86RxbCHZoFF692vL7N1zJ3Y
isPUJxvFHluO6pS29q6u4bptJUvIIBraP9Jp/o1Ve7qCkwbwanW0TU4lhd3prO1R
Fa27+U+jykHfI42OWmnshlRhmtpiBCSbXaQn3SivT9pGLuZV9czQoe9N9ZOt7JMm
OqE5WM+mrQ1xKI0BAlGUcvI5XFz/5BCP629oMgGBCD08jzFfPFDVcDFcLaVLNAKO
BDS5m3L96nz8ghb373/riQm6UL8W70SjnTG+v8zaOpAx07AGrho+zGoFJt5L6zzx
P8n7VxbEZvEwtH7kOM5KpIGrFAcPLiz8v3czuS5HYc5ETRLMAeRHDn8jxUrSqA8a
TvnJjZH7CG8WxPTwjS7/lNbUWHl/yopukQuTUEP9SrWmDQtvC9vMEo6ScqxO0AGj
HFLZXdW6rP0q+erHmJAevUaUn9MQ+h0zOJaYpE6baYusTyV89G9DPO+4PqDdk3cM
S2w32HAS5g1VruUsA15w8ktEVl8Dxwla3y+PDWXBnWyuty3cB8fImKfM1xCEXJVl
ey4+Y7q7hc1MLiUu7aA0r7CdVBolSnF4i10k2+i7pokU0gXt9gYI+Bif8o9ae6Gz
lxqqWkvTziNcNloCr8GieopivNLs8ppsXNpaAOzAnbaBbF1G0EcXTl34L4q8bS0t
ZPipAkk42aMp/ZgjYqYKXULMTanS1HqN+Sq2QLA2hRhSPAqAJLJ/cQiDBp2loEaj
s1hClT724V61bP7+TiuS58mEfJ0AoPk8SJnHeFunUg0o8PDcvPgns1QODbDOs64n
32FPHy9jznUhCFjTOoXnFeBJd0Eh6aTGc3FVIeXWKNFwNym132WF4yvVu00AHSJR
W3vR3ZamEXi5wHH4Ilunqb7ek5lwCjRUVpkeIyLzosS5+aqEroNu6PgeKaetUNOh
3eneR65oq48Uxn2GUt6jxelzs3gb7FN8LXiwY4fEZkcnHzzwtuuIWeQMScViAcL3
OnfeEWkHI23hTX2JJyCEvqi6UIJR1TywKLpdRPft1tJzstSXMim+5u4QSXTmKhWv
eDtQBDkGUA7LKKA/mz3vmmiHeQcC3L3+KdG/j8lkrxyXH/zedqqyN4hV1IhPTqvb
Rg2x5czscdhu1n5Co77dYn8Z9ubteoD0U86xuU3iEwqEyTf7PVFpkO+xcR+rOpub
A+Z6LOQDQwmZ/nhIjnnQVXK15KeAH8ifaOpgSVw6TFkE2LV8/h6bge7ajhV2n75N
FI91+XpyD+AXnkj1oAURUT0+8+qfyvk4hwqSIXoFy2hjsQU4PM8JB0jaKrOT0YnR
PqnFVjO7O2moybMenOpLVV1wW+G7kqcAMqfR610bNp7Re4mBPPB240JMC/TGdCes
xxJwjLKIbi9gqwphwIttYbf9MDruh57qUSsG3/eRo9wntf8XRPV1FoMN3i0Jz14Z
ohmgsXwyQNod9eZ/yxKyktkV8X6rEQHlHUMguyUvy4APmMWrGr4RPHOQ+S3bHSb+
a92IO1WVELqWZNW1HqzZKCI5D1TjKjrbFslXVpdc8UtELAo/UwjUg7/Q5aeH9QWs
MuEgTeIKhz8eNu/ytfrCJAHquHFvLy3FIdVg//alVoCLa2ufjxsZ780LMC/4l6ex
9i4F7wKUOF+pjQIzL/j+pjz7KzRC2axwzKxGzG9QB0eXINnIv2Zl/TWF9FSAANqI
fitbaLBAEhxqTFW4fFC4cx98C0/p9e+pRrEqHLj6J2GpPAfPRZF3G/Qsoask0sEm
300lFZWqQPPfIl03QDIeyXDCIRya7j3aNB7uESzwkHVk8fJRZvrh9+/+Ttr1VW5L
+OGd96jRrd7PbSgZ8f4/v+97fhjmRO9k01p8a8VHyTvM+1TkD6z1NzVi686SbNje
zlFzY3Vx/HtXSNDlZthboU03yBkk2n4s6clQ4Ai7kpJjdzIOvMsdhQVdhIlnNkJp
cQ+uPdEH+9BjAPB8egA8ukMR2UqKyVOxyWxPQFR5eXPo7rqmY/PFhOyIoLWLPBnE
LI1kwMrSv3FzD5p4NDYvadqqMF+xX85xIxSWUqZ7WOMgWZuQ9fGeKDQXpE2JksKq
+budBlrQrQApUw1tdcf3VlrvF+9z3Uld7y7tJmc6YzJKlb1pGmeR0lxiqMqwBklo
mOGTzzkup6N8hTauNiL1SLMG7lb9VR9vvlP4ZqxYSKWZJuViPNOcyjTCDtLTmbCt
Khc/YPT+H3Z4AkJU469qxJj73+rb2ULHYM4Hm/J0MlYeVkF5GFrXgol34jCll1H8
mSkqyadk9/LGln3ILUzTxgymxMVbiDPcPF65pB1M7gF3fc3RGuH/t1RlmWRPR3Xe
ecCFbOqhNdLFtUo87Nt8ebqjdpsfROOtSTYzzt5Xj7UYLstksi1uPJMbD3P6jB5t
HTQfscXVe8hJPYi8gB2sfZbd868T0NF+kOlNNDRoHGe7WoyIeViTb4ofJCZ88h9T
PmFELUGIm5WnnQbR2wEkb8tfQfkiFgQQO8vZNXTfFja8GUJSS5jXewLpXjoIcwgL
c6SaYHxVr3cwlN0ShOz7E/sY1Y67rUDiUZ8daiB/E7M4typFjM3Xw5AQCaiM5VCh
u7cbHagR5yHIL4IyFGi2ngJROov5P/GFrFtSXOZ+FY5i7r2d+59yB4plNphiNSDM
AKC7SLu8v+izo4XYolAgRQGHnYTxGfAq3sWnam887LOmtAT/yB4FXa8UAJYq1B5c
r+mFIifRrzxL5GHUQBw/dR3/2C2YdjTqLL/i7zD6nOaR76ooEjLLs+gxjNx4p1zF
SL5tlrhHj9zab795yD6LCitpf5gbK1/pYtCZG2HV6tj+KAZi5NoE38ywOuT7TLkk
2AvQoUPXkJgDkOnMYfJMnvTloOeIPsowfGheHrUHDORryhjpbui5aTq7az9R1iRt
BC2xxGFqorWHZoJKJa9hTlBI3+Q7AH5HJwiTep5a+ETr3QLL8xRqtXYa+D187bfx
i45AEHX6tA46beQlVA13zrsaD3Yollt+kkKdTMrjQ7FabJyCEh9DaEXyilxuCt/G
YOQR0c4R/LydfFXgDikXa9yx3YDuUtBObBdlkmewe+063eMUw3Ek52gsONNHxuOA
zUtcbRa+3K0MTfa+IZRy7zhViqu2ftBfDVHM5U51YJWBGW5QYtjk3DwkDUh3F0xC
ULnsTRmOKTYed4VTpyB/kk6yE4iHUMTOP/bMmg9qd/96GPJWTHIkf00+x0vtxmB0
C1xBQCPRLkAitZxEh4mzrkRRbWbkzLU33ItThozKqnWYDi/85hUCUZ0FK7YtGQrm
SRDxh9ZgpKPd0sF2JBHZiAhgKEayIFMRbPZIXmf1MBlgegYjpC/cexGLq0NXEgc7
REdIQQ7RqsExm5pwqMP/BJNaK3HwRhABZYoDlxfQCtvOwJCyYCeLXMZI3TsDzhca
6MRBqnPULFbfsNW1XxgDiDw5L+Hddnr3/JuIONvU86zCrwM4sYXNgsh9CdJWAL2B
SHfd6z0EGlOf2KktsIq8RXk+LzMxYEqg7c+ZrXwh7R7cwBkFqeI6MLPKNyMkUrDd
J7C1XwyYEXbC0Evyoz1FoxTz415vfda+X6Tfa8cGAr+pxyAHOjxp3ok5TzEKGRAC
qcwfmaiGFRV99U3guzMVXjipr57Wefm5eqBYp7qT+G94foHJPidQE0fAwwY56qHG
LkTRkuUjHY3yLRUio70jwHthzZszEocPUz63966oHaEiNwlE2ZfR1/xWzLYszqS3
wDKrllnOu751ERt85NJmSStg0jjvSfA2IpVf1aSYLCLUjSdlPw4mwroxd+/ovUbd
1+DbBJBj3vtvXB60oXwuS2RfqodRD64sa3Y73G8BPivxUBwJE3eix8/IGeSNkJKq
XUVC+5cn/W93flVrFF2SF1m2wHMlpQh+RWFiVP1KCQXBfBzc1/c0TwKO7PyU5guR
ViYzETS8sjJ2KY9M8w01qH/NAO2lIDIQsIV8Qia5+M7MiW+gvGDgS7PAecFCRTS9
48373PVpKs40pRLwf6JqgSXi8uG3Nh2SG1JbrwzEDFHcOLgapkI4W0laBa4aKv0h
mMvGgeYBDmXZQgyN4bXQVI85udNSWKqvzUOvOka7q0Jgj+jdy7E4Ua+gamP84pYr
bQS6blaQQ5OaV1nWnnlsDPHpnXTGTScBFo83wig/ySFuwB4cCfYrvqOfwgrA0r6H
oVL4d8WwYYKexA0kd9wx+xRcMSvIFEli5GbFP5/mQln+MRwxO9bEQ/5kWtfKZtiy
NU56/tHirRcUvSPPMhKdpcEJrEYdtHh+HclOva6+55YCzgrcjC6ADHYwUKN7CXGv
5Vt3J9F2ZVjN5v1HiWHVGrpaN/8h7R/65rwZ85vIfGs5Lkkt1w/7xE93y0PjtDPT
ZD+syC1OOqVDNLk/Vuw52Jb18X/lf7kOXTGcBrE1oA2cldx3EDvN40+WdzueQ1yz
l/YIOZ/qeaNkauYnZWjkqufWpMLTbTr8dNBoGpZWoVlk9BCJUSXN7Ku0EaiJ1tQC
2q+iyD1clMlCyGdZZ++/rC76C/Gm9bl4AEzJWj1kyuZYkveCL9nsuKJ2PvPLX+ZT
hsE3Xu6jAYjqMj1RaUM6uxgMm1BMRfdtPVMX17YKclY+XppG3PTh3qH0h7XjLVYc
RKGLcoAB7A9JjXzgxBpUPWeB1OHw/S4xl/ZsmL/o/HCfRzis1tWHvctblH2GvxU0
/6rycgHbICXizSwnptGJwzNMPArm/pWaAbg7xLxnhP3/5BUhgL31l9y2BQfbkxSb
ROd4xHCgyIg/2Lhkd1aa4MnRP46zst7C4W6Nh1+DzBlSoSc94nlC+tUWNLR3NQ4n
PrPYrVFcbtQjd0jfce88+ybughvHURWk3E2w9UX6faibjFKd0uEdNl4hWAy2V7Vq
DV+fJtI4a5WpXajcj+OORw6l7khun76Hq+adi/ZQrnTORLubBHt0Z2ftPdMij5lY
qfro0am2HPnH/ZWQDEUEkvdtBJdse85X/BCDJcDwJpoP0ysXLs9vUHxRNJ+t8zu0
atmSOsZuJGNi+iuuby/F/5iTbyRqZnPgVCGGt83+oYraZnm5yB5p0jAgFm3318sN
pp3gUXEmE2tuzHy90FTKx3WchNo1e9bET8B11a/40u+xwM8ROCY9x/L/eUu2BNKf
iivzrVK3k8h8bus1wjtJ3ZoCyB4kp5WSxPXKG8S9VAHtvSkrI2/KAhPsc7x+PzZa
b1YE8zlJ80MMd46u7j5g8Xc3nE/styHbCw+hza5lcnqjfBQK8rQ9heisu6HJiJIr
U8hwLRzn/xqmR4j0ZHzk7Cn87fo8gdS+l0eJqz4uraZjo+pyKprgp+q2YaVmUd3/
WmUqAl8w8vo1qo09RzWSHGo9bSvFjgcqK1Ay/IGdotNkBNLjgainoxeKbD1opxAO
rcM3J79UXWKjeY6iOpkGbtqey2xhP3eu03tZ0CErF/uB9pNQHASxxbR3IMb5rZrm
KnX4gUM2uJ9RPFljYfLRwiswhl4l2Reu+YmD2VWpH7PeLlR+RyX7Cpw0sS+b1xuP
jql6c/OvCtCBy+w22ybrXZrbnnJzd8jgWu+zDoe4rDW3yE2UkY06owB+5B2Auuhn
iTPZvivZy+kG4c847P1jV4B+d834Wcgs/auu6lCv1Kp1W1UQJ2jZteaOgBfkCM0N
bh2XxueGb8lDpTFP0fo+KUpHJ84aGFqftkxqR253XGMBZqc7JV/ohobQNQ/+FD3s
XABX2lIqhEM2OkXS9S6Pl2SOsWoaH/vz9lwtylqPrNAEa7FsJSEWAvcT6ZpHJavH
zHHMSbJUjNc7Xtn0AvMdM1SJvgrUaVqtikcnja3aj5V/BuPrwWy4hDzdLGV/Zld4
OXYiKiLHbjj/FGEFF0JylPNI+rXfJ/v5jgJ3WoSwlVNhUZC3rSfZM0CZIM2aySv+
BJ2anPgdoWzQe5dcksYk/oDfyOQG3qOfwzE3vrlZ2HMBdsojtN7TffC5mgrHcDuH
PCbPdrZXFP2SY8bPk6Ali6FGoeI/gGNFZRHlgMCHSR0XoKjQd5gEnRYevQFFL15n
n+bjzBbw2YBiGgLnat4ugntLKCPEsMv+cODRo3ZEZfD8618HA5YW4+sji49qmWbZ
kyWklXNCAQPfgBr9rQSWA5UCP8DNW7jPsR+5S5GgpEqzhAaAgC/m0GU/ZR/THgvS
KQz1LoQaefPvq/B7THGIO8rTEjn1P4rA4+PciSUeGPuR6q+DzMX5s6PoGgEq6s6T
G5gqqiRsn4odIFKtcTT4u+8EaFNKZ5GqrH8GISqZhZClE9v54lrg2ZFtUvjPSb6z
3RQe/woPJCZfc8psmMz830oDosCVNtm5rH05vjZeBIE3bCxyaQKQSSdAl5CG460K
XT5vjfyCd7LTRdZo/JpwDocmOqHfiiwO7ehdbyToUdx7ecv9s6h+Tinpfx9M/cC1
FcAJjZEWlbm+k/k+sKt18TO+wW7nEgYAZsH1lezfhNiGjd+G7CRhTOOX+9LmDiFQ
uryyGd4eTZ42uypO7Y0mMmWpLF0sCe/zMZp2uduukpvQnjKMQqA2tt0BcjKeFDHy
qRNUWaMGH/MibdiXiVfiXi01le2WVEbCeA8iJKpJH7b8QdRObtz6f19mI2/h+Dd+
YqZ7Zvap47My+GiKkhMXrQ7k+YVfOlemkbQsnyQAG49eqV/NoElnbGE5Z+LNGSpq
jW6Uv6meknyFQA0W/CG74WoTnJeChHRR/WznWlWC1cDH8ooZuGRssmPp0yLQrcNp
gxFL0t2cD82QUiVwxHg5mN4t21Y8nbPNcCi6IzKEB1QWA6iP0/Biuc5yRFFdizwi
xYUv3h6xaN3YejeUK797ldmhfsYHwXYoBUAOWIJ0yUUfY4udnk0oit48b8Ucxhug
VjG5MGMCcdj1URYFId0hXs8KWCzRZm60AdBNQSlmk21F679fBJi+ZWfzn65yi18N
j1I12XcVKXdQJskyfJLsY+4B39+r2qyx+sz8XXtRrmftrS8p1jRPLDKtOHCjjQrR
ypNgCKiNgFzQKjkog6hSDICr3mb8X/jCY5gVsuYouD2B2UVx9J8g7GqV+G4/JZR+
qLQn2AFeyjqLPEDRV08M/+gKIK0W493wGgn5dHUrEUSetqya4slKOdn+sm2oPNIq
Ke3NBUH/dgi4zPuA/KuOS31elxl9p+bNA/qs21dFeleYkCbp25qZPMsZz8kgnHNt
U29Z5zoExjgD2P7ipbxgAoWE2mPinzdvtXDSrBRe53P3PGOH44lQ2SYm0L9JyOKB
B7JvCyF+xJflutHmjR827JkejC92nBkHgiCor8rDcOAZpxsaK2iYMwiJOErAS8F3
CR3fHPxkTKI9Id4RFcyJWrfl0iqSvrc924LgAYJNZtqFL72yQBvL+tySO9MQ40jA
O7pKPqc0fIYwWHDkaovfLZNYxvk3jP08L7x31h8TYkeztY1IDTeYaWHj0+4t2my9
08aoqlYRr938YjImY6CLvVHx7tmau81cgn1SXv1CWpcnyKSSnDI2/i4lsEVrh29q
gyyQISNPwoyBJKu8Ns+3l4dUrqYQj2Ttz5Af+4Wnk3cldKuAv5N50P9lQp/xDeyf
8wVTDndrL/aJ+vkKygOt5q67yTRbE0DPMx8Ou+lFqxRSgEOcjQA2Q/RuNG4xfyy1
CnQQFV8FZXjxW0zPGjpddZiJKZl/mn5XEeKvblkczU3i/nZp/tFRJrbKopBgEQGO
JCjVKhUEsRHafHCsZQU60lhuMC+nnMXCn/vnU8l1cw36hhrTaWfN8f1JdwxtwteV
x/YPd2OPAnPeDzC7fciQX/APxrEGT4oKMQl9ELIjacS7+cDU+hRxq1fHC8Du3Sbt
w7EjrBsBfKBy2t/+DaIIKPc4Bohrc36weneoIZsDZYpX1yqNaASdDV4CCpeTyXdX
M01GwC0/erbh2iX5IwASEWax6WpkWIgwDwOduYqRWMbLsWp0nvml0+QKYtTi2G0H
AH7r+bhLZOeKfDluPu6Ap4KUL03w2R3Cf9r+ME/kJre/0r4cKpYB6Uj2rc4pUfcS
Bj6F8cLTo5R+QhkOrgd2d92T4sJGafZxLnoz8uj4pgC2ZdGtdGsN+tLECELvu3rE
BZpHbm5Sg60WC/9lFyduYSIqpcO8domX4StusiaPetCcy2CE9rd1NES2bn1bGrUm
+QoEarYHpw89ILgdw3g7SdOxpg0WJyMtNo5bMznq09Ogbi8WhQyePl85bb1dn1B+
vHUaq0T4Eg5OQhrHxNUh4unkPP/AGj4irIG/lLzXSq8dxsMQ0mWK4c1QAhXz1TuG
iAq+cj0YtU1OhYoanZDF44QnmVvg0uoAcGHkcpPcF9euUNNrvxLlD+JCGfGVBlU2
jAXg1q8AMj+Kcb1r4hLpq2ZoBH+xV8AtoLYMaRe06nVwDgJrCIfSPb2mm11aO0H5
LbnY7+gqWLmv8iitCG8HaGQaW1XTGSvzrm2X0JrkzFYuZ6AErgRUxiaXXmLxrPbF
ZgsTa9OMKa7J+Ebx+f5alcL/sBMTmgZuNPpK6BK/xGUbgp8TduSqWLmSy9hb0CEM
VuKf0c1SMZbDsegamCJGxbPVMB0/0fCXm4QK0+jnhCrZ540sA6lcq+A6gDxNsE+B
j2N7jRpd26QYlqWx645JrFEogFnaf6AHgUjXrgdHuJIIj50yE9z8qNaSpq5Tji4f
VbKAZMrX0IQypAn7sBqtfPIFAiQVlKj6BUOwm3Dtnv/wg4KwMLOA8/In0i0JFXiF
SAaig/7xFyPa1W/4y1ERRqT1FfMqXw0NLhAV5WtkOL647C/T9r24hMZNQdiKESLb
KgJQzxFwpL8yQRQFe7GP4tf5PWHp7eDsYfqDeDMswwyrCFrdLrpy2yNakSuYfyg7
zJ1V/wisd1PglR6HADDoUuk2nLarl3BNm+1pkqyvFiYC9DKQ1NZojPt5KsZQMjQs
qTwk0i2py2r9MiRkcEIWGRNQ7cz0wRLv2ejU+7tsLz22S8yLgmHeY3rluglRwocx
A8+nwiPvO7a3R+DG595mVROIDtO5fK8PclWUln5B7AANpdBlaxlhMrPgctZeZH0y
oKA6ABXZ3M/Zq8cVoGtYTW8/D9bh1vLtclBHQct2cyj7b2LcVdpXz0EK2fX1y2JS
rr15tGh4iSwhFHgx1gnjQbHpV3CStNBEeptwPXGuHKm4nMHgqVGLm5znZ0Wd9Ljn
bvy7lXwIAJCtvi4plbFnJReAPsCiPWzQEFbnmKr1iTY53t+29kki95m8NLcyvQmU
Emdh44+R9vorn5H6OyTsRiRVU2YAWdxn5Ts5eweIuo5tAZFMxXxJMBSJLZZY2k1v
Agvx729tkKdx+8O+S8ewJnDC5U+ztrRb/bObgCL032t2Ly3ClEbexDEYbM29v4bN
qT6HUo1Zt47hde+Xke/fqAAEfOSeOZGyx5j1AlCZxBTAtHF+Wa1H0NH+bXDYsGAm
z0wgnWDXYmXRNNzztTXGJWIX1sJLG7CcOu0+Jep2JIULy24RGM/jII1RPmB9+qQP
Sf/lMxriFtPMbQwceChToFQqHHzAN9I9FO4hN22WUSS5MD9HyS6SODdVVsIFYMxf
2PN9cky/R4AfwTZX1Xwl89vfNgbZJ4KFmAZl8hfYi/W4e/uBt03sx0jHLWzwrrCc
pZhYpX9DpxcEdwae/5XdsqSoM72Dk2R6lSDbj9bV+SNy72mwONriqeXOuOVofe8h
6436WO02cZMGfsVnjsgtKGmwI0ChxsNdOONtjDSjrqVu3Kr21ewFzOKuvDI/B1fY
yL591qm9zmBrzkqzA2yIZWaxBuE6/aQ544wnxmlFEI4g+XkEQEUrEaQYsWIS8BKj
C+wlb1I5d2KiF85HQoW+2Ti+Pl6wbjrQbeVqMtbJ7+BKrjiEYozVPSbEjl6c/gCm
SPCeGbZZELZCliCKsjh1W0wWdJPHJS/+XvynXUugKQas2MlErPGqMeBUQNZpaj6M
HUKqDAcLS4Btnm7vs6njokcTbmLHaxYEeHUw7sc6gzQqd3IgIIixJPIzdSYSiin2
jkePCphmKkGAOB+CkEolNV0fdmzxDod+ne2dAYsYybzMLFWuHWC4BJT1Bn88N5Ym
c7rRAz8DvTDWG9Uxgos+edzXYXATo3BEg6tuIKlTNoI6DplJwT2fEEC62tSE0Doq
Ud00iRuJFtFL5G76Q7O1i1C2CoWp+hMxcV5xbiKYRo/7bYLRHpIf/bc/Qxt0ff0y
KaOIRifiUNGPqMZIERQe3z+Hmf5f7EjMJu9Cp9vt19jZl7f9ysKEHuXvSB837yrH
iMG35GjAdtWPn2QOB2p3JSV+QOJoRLc7vOusNQ/blynzj5zYbDt4XJ7Svh56B30g
LRg5WcEL1m1IuhbXbNA3a4dgTZsm552ABECKyMgDenBI0VvtqVTQUEnvS4/jtOfp
nGUAWuy+/oIcMmV3LXoELP/acXSfmeccq9gDX9lYmKm3tXgsTktflRqKtO6sQFUi
7uLEWpncJ/sE16A1/rnjJSeU3DG9Ag5tx+ek1Q42uzuVkowHJANI6M62mQCZ6YqK
TyQRW0EYXp6Y35eeAapjx/eFg6fV2pZGZVogGTWsfpdDcArjUOlS8oAmRxJ/sECC
3KkeMS5mOCSwFxLM8JoeZZHVcXWsX79B//1XzX+dVIN8fqQ5by2T9eZODntuU+gW
lJIkTRufyhD7rHCzFDWbslCMKJ2XpaxMc5hAut7+1FBci7J1S/lncrmuu5Sbh4cR
pAV4Ttg/yHron/cwLthwa4O15h9JZ+XYSyJAQy5ZPzfvcHNjeTRatGj73n2Tk0bp
5Q4hVtCgpeVoc2TqN7EemM5FHkR/I10bF6aCLbGMgLdKUpj1GVjByIywWWSzmDFo
si+y64QFFkj2gCK/N2t4SS02Zku6fx0miToaplR4r1Z/VPlCXQ6Rt5V4FoF+a5yi
YdVnR8JyE03CxNJpoGQJOI2+Ol0nPbXjyktom1r6222i1pbLQv1JpRpsG6KNq+aJ
vivrJ2T9ShsMFN5QAFWOQjfg/Y0By7zsyZ0Z5QiNGjNoXauQ5ZjszWl1gETCFsKx
rH3RmaNvZmkkeYXtRCGbUEf+d6IgolatkQizAke+KXElujZ9Ekjm3+KQdffXT+Gn
AksnowKcHvzuAS8N7yu7md7GF5qykyXkE8eUbbP8A6uuRKMfIxTNfEUieNl1zyfz
4ZPGXc8vd0hYjDnyCmUX2UwFcDxjvfBvKDXgy7235ovUmv4n85YZijKp3d5C+TdM
iS8Zd3XumPkXrUHmT+T8Hl6vwKcLFY8x4+eKlD+hkfEeS/nPmAP9rLOFDS+3HzK5
B8iRklafsihL/mKpxR1LQdF+5gmu+KmrFPnYX6vdFMy8N9mb2a+pWfumnkckuG5v
4SiM0yNIOAfcw1x21ABkng2Z2chpWJATRV9mCEjq2Y2gPLqTBuOeLWaxMk68DvcZ
3H2Snv7w1PWIw+6czZqVquflxMaEUcYa+Y2TnjqE6/p/Kq4PJLequtfXxDFL9z5o
eI8MGJ39QmppAddcB1mXUlAUbKpXUShdjooX9jFdpUld6rYhVNJ3/MWRR83a/zev
lZ7SxDSj48ymQhROfBBd2vCx9bSfWdOsVzOA/Wc8M1Irb0Ksgr+3tZJNjuDcrPsC
+RoMNOXJOXR6tccL/fG305t7xMR/6b/SQj9W/O4loutFpJQ/PFnhYSPsHpY82RNA
NgjsGwlGBV6Bc9DZc8x2EShYCMOnx7cCj2gxoe7lj4zadUNrxP+F63Qq/OfQn+s7
+4sLAYPuYyvbJiejcW3ISBhHEeGMLnkPNKRvgDHkSqX2PqApYux9PTzZmMM+eH0m
RMaGScLXRWvgcumlFzo9Tz2Z92zC/xwIKdXqG7y0XruayvY6HyiS8ftVBQEeUf0q
SXHM+p9dP4PUKBi4sfPrZ4ywEirnY1zX+O2z5OidaEQTQzzKOnSNWXUVS9kqiAVi
Ttt4tJNneSTWfGkNCJwvBuZ/e4amlNcoDaLsNUhSXQ0i1S5J/7MIMgIboAbWsgM5
kMJGLv/F12f3COvSork4z25964lfpFPVUpCFlbEuzcHBI+HLUTEfbVdOfJoSWXif
OO7B4tzm52cDHxiaPQRAD+cVp0tSSOy+CdMrJJ2Je/j0kDFDgp9cm2g1B5ooh1cP
MbEsYHQxcWJPP5op1PM06aO8Br4RJboq8dzmalYUSVABbY48Uz5pQdP4Gy8xV9b3
y2XjRNB/RdxrrkeyfGNyU9yMtWU63jaQk/GTcbpitBzDQ+l5CHoXVqKRtmJsEmxh
pe8gNXqkrJHHfYBCuvz7LzB39cN3DqQVzQRa9kkxjlDeTZ6rFOXn+CS7bU8FXTX3
6A1XRtLv79MXDX/mamjYhOQjMWX8HfwDcdE5pC2KMXq3KQkzJ+uv+C1fj8UURgYo
rIcW309P6rNUM1rz+ZCB7MUKS38YWdYdOcWY4ry6SZOpFdIKb8Dmx9OqeqUXFd/X
KyMSMxw5kV8WPgSycuqpn+eowcwKSl7+kQ8Zt0AGuSlJsbAwAOXTkQ5glYqs13YY
RQVYqhpKIqhmgna2z6sHQQsEb2rXBLUc4Np1h++26bMWs749E8ZJ4XR8BMX71oXK
pyggsFORl7i63sW6yF8bJ4Uai7wzSjChzraffFISLfTupSweKyIfHvf4PjpPsF0K
5jHEWopEOWZO9Z7CltPVOu8bWe4X7AelGhj5+NHmFJwnE0syjD89EqDT+ggNfIPq
m8Y8OpO7wdBDBCrH/Sa5NUSIhSfGo+lQ3c+NYrKd1joRHCwtyI9DVv2IoaLRrh3D
QarM3CWADzroF5eBopdMptV57bo4R09jk8WssE4EMMHUUeS6Bf+DHK5lP6yY4Dxb
h2RscCDjTad9AgBfHBTXkOxJYxR0Z0hPwaZJAL2GSt8wISB3T76lsC0xUex0FoAL
tsh10MFafHcohfOjt11HWbeaK4WnmsewS17obDGePd5weB7gsdkWJPutOxzg7MWs
sX8u4jsT5X+ZgC9FunmKtfpEk69wwjyJqfvd9qNMl9IYfMVi31UeAexWdvqnIASr
9f4bBOD3A9mXBiXjpVDvOOPX8hAsMN+/HSsBHFciHQKfpG9c/J5Z5EM2FOjE+rOI
4FiF0aM4Jqlz5c2NiBxs2rOPZ8D+K5Ojjc9mzEZ/MnRuPTIlYDBbsTFJQ6NJLs4M
ZuBZSh9w/ZBpOGiOaNtzMdOpsg69GgC/KFuIvA52Lq9mUjBCNc1/hmBWhKPhhzrO
S14ImUaSVNdvDl4/30o1u5HzI/OAij110JRC+j+BOHfCBk3xEpOa1BofbzwgQQwC
QyUWjFHv8E7QQB8HicVpoYUd2MM9IDb1qRKRWDnNyMPnsJEQvQuJ2ko4jUQlTiiX
QnXtxXnPnx3eJxQ2BQNgeFxLfF4nqv27MajY0YPQxqfLO8wfQpL0UEjixBgoYKVc
kzGZD3H6BcMUJ2E/aTV0BxXyksXcKcTt1UGuFocWV3iiXBhxSf3RMgBhk/51lRAU
WT7L8ORG9s7/XNnArkg6H4X36B2ly8JBhtEV6dSXUAfm4K/YaEJ0GXaLdMlBD3Lk
kO0aQ6tVFa3Qw23+CEswI/wNxC3vF8DWYvYy9kSdQPznFihfozVbyLU9oStbnGE8
/1WvQMhUbF1pp2KXpYrYvap7yaj8gXxcll4o+FyXsGegxfQSmzSjmFsk6tBViRaQ
c6W3puCcA32ZthKeX63ivx5o/bHlY9jbDATjBrNavO6NPthgkNVpKzmmn8i6qm+5
eD4CRTjEgVkXIIUBrbmG//0hzWnpD5ylkgjiBidWV/mlCDiSF8Zes6t2T7YfWZ+H
NHd77CUgA+DtrJpaCbG2EuOKRwFkQBmne53cDRd5nOddeqUorGuGRMEOZW17AZxm
Rt5BCXd4T3A2lZUh2pbPTMnui+5QG/bEnGD2ZnbH4i280HW3XZCDXzJXoZWz+4mV
CdTERrjHMpNQ0Ieu9FXZK4vDTHKL/TbASoRDB290LuYJlAaTDpuWQcH4ZonWnoBQ
Q3RZamOclAnU4NNkwY3ia8g2wNjmmfuLC312fuXMysI4N02aViR9XwRuHk4mKrrE
aWu5OXKBbZ5hvaUeZUbZhUz0nJ4TL3mkGM1T9McGythUTxtTC9dP+tIaMiT9bwl8
m9GoRacUOldMqgqm49biVtjn01vODhh1+EGgp9O05J0wInU5c3c5mSOq1HekaBVL
aYnGG88vVMFi91f2fWyWZ9KxgVQ0rGYQdOVlxQJfvuxVmNdrQyJVxLHx4VjKM1vW
HgsoC+sHmuXxI/Vk+0gcr/sIkbgRKD+i2Q+E97t2LlkUolxrHbmCvg3t9DrjafD4
SaaF2vdxIFWYyO6sXy/RVU67oPZQO7GdX9AaCUbpluWO2A4MHAuh4iWY9SomjuMF
fqq7FFu2zZnhaG+tfZ3SsOjHV/5UAw9yXdvAGvX3cbhvof/5LgFHmkoCpYlUOLH3
i0C6s/gbswNpXqDT6SbfvzsbS9ICs2M0XaJAHbMoPj2k0dGbO3VKRZiBoNVTlq3O
jBKRMPzQtBa7cxq814qcoHSXZ8knnCgvT2/H53Gxk//2WDrLyTHxXgXPDBOnyBbQ
IzVJ9gtZ52XAjcPO77RyujNqtE+3d5c168c6zcg8Ahf+V+hkvGb7My1oAjkt6Gyt
06uHo2tShuPwjPUxrx3U8dHjohsA1F3ri5LJrJKlSIix9BsxfdMMjU6V+i8yaC1H
86QphkRSRwnUgWYlN2mEDxSW5oaEhBMh4YiPDnEMYY5Eb782J2Yf7o7ozlLjLJ8+
085y9eueyRhCEnhV5Ws+Skinhsa0RwUBtyDvWYFzg2eXp3ebmTSA4vg7tR2LqyRU
oCsAVZNS02zJiOIX2DU4wRxtogEiOZoYBquFQiqmPXwxtDP/p6p/64x0heNqpp2A
M9INmkP3sn4qkqUnPYIu8rl8LCM57Da3D3cexKnkffOM6hjQrz6PRxD2PhHfHiy3
TrFIW3MZHZ+bnJkCbtmg0RB5IeCJmxjJmYCZSr4IMqxkTRW0KphuJAPVbCXMB+UF
fI7a1CI5/XpOr3uL0G8ucRAVF6pH8swxUy/uLiJ6DuRUnlIdKOnCjRuVXFLvL1/D
p7xmwfTXzsU2I5y+zDx2cjCslE7hliokJfTQjU8IlBwgEtogkbrrK9eY78WMZNbv
THcQ6bLum7lOTq1C7RAzNSzEleNDCHNUzBwjmtZDsV1Zh4gibV5SZ4jI3ISFvR/p
F2E7d2VXREtGk/CRDBfmv67PfHUhKlhfrwmiW5LADzVQ62pBsxrJeeyutjVGx1ku
sCbUGDTlXRkTfIfc0iQ+dGQT7FkXlO+SER+p+B5/1EBDOBZIhCLvnm6l6qQl/VPG
8hXZWVBezJVMQuKfVb92SjlpdVgvYfq16jqtHxnnn2Bwa0SY6OkmNtRt4YSwmNFY
IiZWzehvCR57uD14Sgh3pwxYgkZbTs466rIA85rcJLOML2N3+gjsXocgkJUTUKdu
S+RhfsrqbUUtEW/8LGuEgKbldB7/Wz4/4c0Jfg5UoGxCQaWt+c9tq6jTfuV17zG+
VqizAvFALrC3oxOFXqmY19akMIGsmrHDAmTC1IJTMWUO3K32kAHDSccwxJa6KZh+
0/L+/oyOy742plTeqkkitYaXEOU5ViOMWnxADoYrGPK7TkVFHyq+pNVT3+ezjpvG
4oH4hDl67JoNSMJ+PLQgBIQro/LD1lU10UmDdwbljGC41hXZ6ISJnRhGVyg7Iwzq
2MxQ3vObnUIxETwYgDlHwvqHwQkr8piSqHcJI1HfQ5KHHYA7bKfrwGLfkCVJ7Qud
87PuP4k3PONyQRR6odsgerIoiHsrdzcagKgvDVT7C39meQ4y5xPuNhvNds2ZAypJ
AgKqLUKxpYpT1V74M5yseVDyCDzTpXjU9Jg1XUvv8uXbYLY21ZK8+S5QiPnl1qG9
0k8EcXDIyVevDz8uQNZvn+Kn1bkHqbniIWRnAD+ipFsKfaVg4YEmu8ldZiKp7FZZ
XArtKQj8gB4swI8pYog2dwEvbrDs0VsGcpq8cSLFouOAauSrWIW/AhsgZVzZe39w
XzeOghHSpxrZJkU7buEDJpzkgh8veV2dwluc9YXe2nR2t7ngHO6Rz5MnvdGXtAgU
djSc61IZ38Q6xBot6yLcRpVPZeswNVdBWth/ryh5T8gHG/0MmQJ2Ta0X+8ESLHo3
4LKpBmp8zmQrSbrp8g7wqy+eIMyydfGQ+S7WLr4HZ/lOAZFJ0ueKYBkQBipi5/NZ
kWSH4jGFWlfgrgRCha2SX+5gapsrF+7qz32uGPE+vLkTQX7e3Fut9BU2geK3LFb/
bQxxC7pbbVYuEzGJ9wlruq5kNtKmlVahjWS9Rly7hPNo5cE3FlCBd7D7t9ldQezk
p8dqUMNXDoEL3eP6c2VHXUEzncf3fbTdh81FTbBvYHRTQ9CPbA7P3t0R7tJZDCPE
gG1Ntq5ZGoS2CGNhv3ZYoJl/NExs2ShVirsv8enEUdUkr32uBvdC5eC0NG6vYOpC
ChiDT51PBOX+w4YJUgtCsZEsw5oNex2VcDYQ0lzRfV3NcqwfdTLICEKqL/uVXQ7p
Tf9OlIaXbDZ1k/u4Vo991wdNwmasMF3KCtr3W3wxSiIKeG8gFvxKHDDV9isrYF8X
HCi+BSR0Smq4HQYlJRO1FTTFrR1aWusXntk7LgojWMlyds7WoiV6saZ1Of6WrM6a
RCCvW/0vBmAK4H4PonQi1czUS889mgasFOg+Fs4ROSUxr/b7oPK0ik1xl1r1Tje+
V0asPrsw0bgRa1xuDSQGJ2e74RJs31HwzpuIFNq9v7SiAv7PqKYmwxZnaE+JORzC
LBgLtZ3sf5RQc4cVwMrSovd9WIiMUMO/XsTQNpU+a69BM37R0aeaaGHRXyMDZJKE
fKZpY6dY5deS8Rdh4dJZJ6W5FDQ+bS7F3lO6Vn+dyLAPBW9i3Xl7bxXLGjdQSiR1
RI4VMcej6ONG3hrewUEfUo6vmA/JgqpabhlGCJsWxX5xQKSkD+BoNHUJ2SupTkzk
HgprqnBEAsIdOVGIOYEj+MFp5opZtgPYxSqmeEQi6w5h/O2ffT76/tv/A1RcjCVN
XuPx1M0wkCjst89b+TB8jhG+fm0Ignr80iO0FdIVvbFR7E84dVML8h/2hDbwL8PY
nH5vmXSgqGVitmj5hBGMefcQLnQC8I/2FryteobTgP5asLOdJoCxhyoRpf+ttOpI
AYgCrbU5/4fkyiyrsJw0Qlx4sWnUeDHWGy5s1dTtRDKlIm7u0+99cbOSKXqQJQtE
oy76m8/B9qkj4gVwHK8pYnueHUgqvh1xvNM5JqZuHjT+EdIGBBVkO2GoDXaeCQAO
INeTCUL9CbPTLKXt3V5Kuwjn+JDb/LjHTKrs+zPWTgV9wX8+EQzpucScmoXbclFR
5SPjqdLB3TwEwt2E7HmCcpHxX8DoAYQECZuF+2jhs0M1vLMb3pXJ4OMLEUoDRB3i
KhOKf0s9B3M8OMkkZRUxCMb5ZaYqPlrtC82qbIZDru8SaZaZBx8qV8DrcOl2exmG
GGZAIlBEDMQwjhf2SI6xiIL1wCMTuNQfCMHzUPrUDS8OJQWpMvlBndlkhBNU9RQq
AJCLtdhlfsSLGDbvFMvTaFOgyt1v6mVeqad99NDHhW8e0gm6ghylLBKElh4PZDVU
XNKuXSZ9795fYM/B/IZ68MLhP9S8Awzj0jIdPWzIB64VNj+ByTdRaA8+G0dZ0D7P
u4X27NHtHDxNYcmPZkLwi+APpM9r1YhF1rv8nZiOiiFqlYqjIN+pIctu49embyPH
XaHVBjM/c3M9EXGe47DYW7w+wZcmSGES9f8mGjHgSrfvICigWCZY2eKq3W7pXTNh
ik3/m50tYZZiXnpR/Fzh4n/1GT0IaPShL/6odnquFwr7t2QcBoLI6or8Bf5u0tez
1TXxanFsPbzEUH76FU3/rq5ya5FOpJI67Xm5zwvjT4D1bzlvnUEmlXT3qX11c+Do
E3iK5ayHYhRMO0F+uHBA1aSIzUJ8EFJb8I0OLv0KJL6+S/T4I3Dtr6XPCUnwam9n
3o/JuZo8xQMFDjDkCtTOVcRYqVE3GtHr+FOgagw+/BmYxQtXuQMyDb5+HzF26NRe
EAb7o5cYCKWqtYRzDxyfeke3u4kmVDgdPyeC1+MvE/3FfisfOWJZuKypvcmtVcBp
XW//DB9zujn++PBkt3dt0GV+uLxZzP3ILOVsPPOoSLxlep7VV4O+JrYett427rKW
+A7oCXC5HbIGt9McFncCROP/Tqa70ZQZt4VXLB8H3+y1BPVySrXaTVEuLEXoTTEx
x3UCrhLnqVtZCbU1VtMWpRLSSx9XYd1VT5LIKwlPmGEMgUstU3a1g4kPkOdKFqCM
N87WG3A/ob905GiyYTMifpu5P3zbpX/rukN3io3l6QAzAacqdcD9ZUbORFp4xv02
q30zAM0pmmv4/YXT3ZdfrHQp9qjer2yxWvc0wYAOckFCrjXGUq5lC5O1T94Z3l11
ZQjU5JY2kNbvhGBievbO3IH2du3989GRfa32AgPitsH/9gm2GbR/1Bxpj8BXaqAE
7JystDvac8V6r29Myj0XJtaj2qB6yzuAHA4y8iFdJzsekjLN0xP7Z2e9C11gA3iU
obRcUo+wR3dQ2DVo0M23MKUfvh0ty4UYLWfT7835MBEldUNYkbhK6JrFJ+nHtKGX
WpHHpTKGTDAH4Rc8ZvaSfZBnnZu8XSjzMPJdrLZFMT6Tp6ZEOPRh9zrACRkS7V9s
GK31qOWYXIvQcEiDZwMqJCoi8o7+v34i3rCHw2TVxQ/221dTPBfB7piEs7j7QDB/
+NHN/JRR54KS0BtF0pFvEXRPzdFf5I0Z0rus3/ex1voup0jKG6oCn3d+GrccO8ZV
Sc73NQ3k1y0dJHTUcwu6WzsHUvLlTMoG5IowaUK+zNBSICgpZUSWUkrKBBEZjzCq
708zWCXIM9G+bFtKMGEpJFO5XUxZMs6+kyXZ+3aiKdM0PFwxrISZc5qaTsG+Sril
toalcggSehqeaKrqxRczN+Ks1Jto4yqVu/6SW9s9G70Ekfi+3ki+2u8s6PZ51Jwr
fTlbH6djm287P+mp8nZOtLjNl32O6mwXKbqRCm5OaUjFU9Rpxmyw0YSaLAxSHFBy
AWRrVA2OIQ3Q3jzOItjp8lEhCSzlr/CI0dKsNt7IafdXvvgoyL96yAR75r3z1c8m
LuDvKKwR7ajjhlA0M7I2rinIz1mqcXXHioQ/mBmm86rPpQoRcuKsbQat4F+6LmyC
DHf7OlIQx2XiBVzovXUArsXA+gfercrt9Wl9LdDwQiWykGeAOMqmeK4A24/mZHP6
CpFaoKoThOQHIfWWBFiomifZ8X+weF1UeQrjVqP0yzxUSi3KP7lDOawZvxTfCPyQ
WbTnFJS1MqFhFUytvNFToJWKdasNKzFOC1dB5zgN26SiEuI3mrKUQ7EXjDx0ZOZc
MfkO2U7lIDuAi0YVfvKMXwV69nxK43vKqztkrBYKEnkBBFuw2EVyb1i/Ij68OUZ4
dVBTBlNKhtL5BImbH8pgaO+VCrl79Lqlk+TKr7P1zgHrfNvw0GVBsWD5nkG4CsbG
B10bqQAxMhwBiSHL+rU0SjPJBQJKFH7LSjQZKlkaxGPd4FnkzrKnISGLdMPmHYWm
8eIcCMZahE+u7UJHNvYVhBvvvHJg8kZpEpjMwZu1E3skSX3iuOXuLu+vJN66zkmF
fB/eutxiDS7RXL9Kh1qAmsuplixxpcPB1Bz7fihEnSJx1HZcPx7P7ojY4l2K4fHx
zEH5BgxVjO1gtTDkK7y+gJ0PyZs56aAUEwrCFKyx5eM9vxFFkBCFu3U8YShQ0t16
F2LHnaUJRw/gqFeiJI96J3p8lzYaAXifdBeQOj395NC5Mnl52GtByBMnpojuzWAE
8i5vw4Oy9/JiMWCgU7UyjAut1eFyMqA73cGt0Fbnzw5fq16sBfD3v1aHEs4pPoW2
wuNuQpt4yspLabzvRj9DVOzwKXm4zZ8g1TbqI3E+cqY4ivM6vMQIXXK4eAiA447l
qMJ921M84TztuLEMwfWau5Zjk9Z/H5O5LurSmTjRiB7n6pHDkRIbRaHxTt1XyQG7
C7cFx2VY6wcXHkH/ZwBv8TbqrvJlhm21D4oY4e2ApSN82QakN/Q/SG5957CvmODX
hJpB+gciKF+MZUPZ9WkoI6CMnlBjdNYBR16/bwA6oQDNTnubzY0Xm+/LgYGbl7oT
QXx+p4H/x3pU/e5fDCQlk8slayEEWlwz+2Q5w+p+Dnija0z7GO0cinpr5IpCa8Aw
1eImtVmaNHJtm3lxi8FwtHQymCYqazfEm7iRBlFcowS3GFPg/dxPP9OuHyUykcoj
Iv9Yj1swPNYosSCb6RbErxzL3DUmWpAGOQFlzy34evySUFV/0DuV76CQb2mshnls
6T/HE4u+sQHi6KOY+mF8b7/D2NYv+VxR6MytnVdkuk67Zx1qkhD78KASZTkrdi18
3+nQg9gUo/cib0WulDJeQivrR6gUE3SymKqr9uuOOGlmdqhpH0DvMZPDmfbomAx4
qR5hwSwRxprj/XBoqbInXzL0WlbdWWS3yGX9B/MMFU/3YsRy1KvAA73mOEeyQq42
tTgH2t7Ao2SdbXYfV4o2p+GFeWA8sCCf7skuCyq3wY5m6N4xn627pKcZc03ykdCw
9oFSHDziX9nJfn+PzJWKMmgy7u6CKu16JFIOjFO4OKnGMKgomjUyIdOAdcftETvK
NOBM6s85lAXpHibxZTssOsVXvkH/uFASV9Q66t0t+YPfav2eWDVlDghkASjqwyyR
rl0Q4aeQIgId2olFSwF4iXHPgxer0jJd6zV3A5gKlKW8HuBEmp/HklmW63+lYI0N
WpsSnKBTZFuxLJ0Vt/M9FjysE8dFzROWdvX/bRJIh+ns9kDePqlyM0YEiW1Bf83X
b88tDIMl+y3Vvx0ZpGbnWrDdu8QEx+nbWkD+fj0ReCWRonPuoea7C3hiRqk2zC33
oRwdc31rRXpzt6V1u0NyJtQwMgtMUgzNmoWEcPmeijOQ49JfJZHIWQPpO0RQpowB
xr6la3vyPFmzomVWHaGP2+i1EeUwWpeiMfEnwkWhJX/buvUReDaY3wmKr7MuLyIS
4CbBrcyttjDxG+A2aAqP+T/F5NSfUIlRfLikJ2TOQT5liSHnXqLBxM8ZAvYqYDxU
DSwi/LtAfYgG3dXjoQzmeNs1tRwk1SFPf9r8klQMN++2RVFAAy6M0BsHQ6esC1Bd
AGHDTW41qHzG+zVbqAZe8JytFLhBs8IkeJ7WEA1CuFSriwqRDkWCMo5byEjcv4c8
DhkRkXjtT6aacXHk3+0c4A7jki+OcefcD9giM/2UgYSSOVk2m73dRKU5W0orAk7/
O5+rtWHeKATdZbq7nnIDIN1y59Icpwhe+jqQuYHEUDEKHbx+lRd7qxZux1itNlvj
AImlItRB5LuyGLD+Ldf2Ljsd1gAyad5B+tDw8BCerdD43q5a45wAGsMfyfnnxTfd
TT68hmXhQTai9+IoaxzCkjwDWSp8hL1k65TP5fDRoEKnMpA43lssgFk1Xmi+H1HO
iLQKzzoo/zVHMhIaR4oagBcalezzRp/Jnrc/zRNV5Cf/W/jumt6VV4WosqgmboXT
Fj8XJYjMrmVPgEqT5Njz9AV8781jRo1G40r73v1MESECytirK8u83nW7FRk/7Rmh
GtymUUcckcuvbM0gEJouru2oK3pBT7pq7wtlxwIUO7QghUEh9StoVQWg15c0JhWX
D438GnWs1TPCFIo8DB26u7xmHlVCqafSZ+NjmtdNR0yLaheY36DIAMkT8UlAH7U+
9aZ2RHqsZVSgudeMjHPA35pAdJo3iIz8lJxz5hVRN+HqaKDUpXwS2yumSvySm750
iU/l+CqQNXpJAlMeCQwQDrZZkp1eEVAt6DewB79SUhc720eHwRzK8wM7P/YTdHSb
uQfp62UKQoXztJxzT0U+mZwW+V5x0KI+0V5w0a8FBrn/7fWTY3QlZZYCtXM11gwU
0UnIbhsbsxguO7+iWvNNk0TkJZHMZMLX+g4kN4qIKcpS78NxXuqGxiuqlob3KibH
BHRyZQb3g1L/N6GVfqpBUZddXaAySnK27HK1mIqllO7Ym205IOacTQKYexL5L1o8
JpywttAX1qQsyYRFBA4JliBgsg7CbI/+958l+/pDntAGrwGH4oD5xWqKO8iid9+X
lIlMh2nE8mtVwiDkd6BvvZf2dZyRRCFUt2Fe8n0jkYqvBpIqSIxReCWss+56GwPe
Vqarj9E+FTqRHKpXjew0S+iVP3eVQkie1mjO4weuBLWxmBb+DNt5pigvPlrQV1Uu
GBsEYoZAUqV0e5v0RgUc8CH6OSKNhsrKBovxH3qN6IupH4Ht6v0pw+xuNAP/9vjx
2mp1t6zm3KoiRK06vF0LV9iviB7OH1C4CYwONF8uS5Vzuwo3zvMCJi5b3IuqBfV3
kUCEOWp5cgDkuMiIHbeU9AwLwJIvOtLELfxnQtm6D3HRc6pec55Ye1RI47EYBBfc
FrVL6i2JjPjVIjo9FzQqn9oPW2Q9cKsId1wQQkSGuI+bFKwpGO0x9RPmxnGEkB0/
2pliwbWmAuEaIofJAysY7YIeUc9cFnBT/BmogDrNnFinJhTh8iaCYAy226URx8uI
kFY7bcPTdNWqBPh6WXrSZ9sQz2exr6CjlHfUdV0WTWXOq0NhJeJ3QoWdWbVdsJYi
DWFvSp1dqi/PDH+zOx9Z07+QIO812HsBBgpLW1gmblNdz9vtxyB2sE18ZBfNVykJ
ZTcpWujECAHKrfuIc1r0Js3DSbtCFFUU/VT/r8Mt42UJ5wz23K+/HmLR+5n4Yr+b
Bt80sVclQP6Ff1FcSf7WuB4oyR4cR7RWfxLAxMVQVSAKVLSPq9kQpgll7zIRzGLz
KF0C25HfczSOZhiBMi0sGOsjX2XBUJdfyovvcLcQxKTnRImMOV3xR6BawumQym9/
t0pEHDpegDS4k1JipTjECfduXeHUpx9JMBCraSHrLLWY+sTua769daW1KmtCTVEU
gxtNBt1Sjjspy1Pt6KvhXLE/xLeOvcmZp0C6Tu+KIT74+pT4/nc/Ou6SrQgPMGar
SC/KlAFH19+PCF/wzhkuqQ2qlOcPFSd+yhGaOikMm+j4xRppOhqT/sNof0JAsCSn
z2zutVY8u1NDuG6blTzJkTG9jraqH7i2gCLMT1+zwxeiUQcHLNTjvSRA/iTiCn53
YHvm58+S/NtUgEaW8/S63tmjQvGwpSB2SULDKeQQG0AgdvdYM0dxNDwLi59I95jm
9GpDxelsd15XvRbQws8Gb/xsWF502iDo6/x/6lOMLD0dPpS3hGz9/6LG6WrQ3Do7
1GQL2ttey/qQjGjDo/MWZk/el/83rQAFluTSwCRzYfvN4mvybncKpKkKotonu4J0
tQJivB/rngqpy0TMeM6E4+zjMNNkKeLYhvu4imvNdP66KXCShrOErPWxkz2djB3M
gC4adyPTJqo02pHzhQfykm2sS2o758iZ9dk7ECyCHRClCPRCRTWmbokW1Tc7w3lt
FVj2rzEDSTzDDcMMqi6MlI0udC6aqSPYVQib4Ph40FB9pM2libQhvszYG+CaMjE4
S4ksOwOrlZOE+/RY85XpRAMoWBIL2vSBRDc/pPF9ntkrS1gYoWoxk9BqBcgDoVSP
NkIYZjmbCa2H0lTQgwUy3UZspJ8klUQgGaqwAF2XK2ZxBL9c89bMyeYv7oeQTJFo
pr0EWzyhtfo5uRpPYuX7btO0PW9kgYDl5Gkma6k+gooTa4ChIHi1DQ0lG2jwOUKB
5uKrOm/wjJTiEKIV97Squ/sUOX978Xb6ZN5CY/GUtgs30p4yEqyv1YFiYGz3fuQZ
kGKTDBAZOXsmdiUXoH0ZDQjbvZpCFog8G2Aww2J45jp3lk1Fef1AMlqrlJPCmyqg
sW5MdZsUZpYvn32mdincVTx/2jDVEHNr+phX6PXO1ASBO6b2AI8KPmFWBf8qRMRO
Q3QZwl5UksY9fMqx7ZHwVxNbE68uqU4SSoKzXd3YRlQ+uk78MbivU9t5j4Xm+X0h
dLAzBbUU6kssNhu9fkQM74QdAKdJUj6OIjKZ/RjOY8olK+SGE4Xq0049zt7QAmPE
igt0AAS+dBKgTuaRNTvB3Awh39aZS2D4e8IZd1LcKmRZjQF+VpToqN4+aUMkf51f
cFP5tMdNs3PVTxWfxDXSX1xEIHfGcYcTl47+yHlDRH/jpfiTdPtdaIUMLb+irEaw
Wfj1+MoXdLb0Cr/G2fM0dT39LPktUX75RrSyF5HeJmwLUSXR7IxLYxkinpmhqXVu
U0uJQ5im8ryGSARgANYuitweDiTHwejO20XdWn/PV6O3kDeMNmWzi8FLhZU5pp10
KyaPI9GdBm/waAhoBRlji18tWsGsdPETX+K5Pg050niGGtSrMpnL1hZShp5Q8TTv
l6XE73nD4V2HM63qD5Ui10UsOrLzJzkIXZvr1VGRPEA9yANuagQv7y8fonm5dYtV
MC8CuC1KDMQUxaZe7g7CBbwnrCfe2oJI93erVNc28jVPJPsRTuEN4Qg7wsyzhOOn
/Fgi56RbFnl9sfRfDVFc1aPIAVBqw5rVgetxCa0pkrSHpRxlDgGraWDnh/RDl2Fg
QvbkIYOCYgtrOX3gQ0onIYxDzxP8B4Hg9+wtkZZYDrtx82C35ZDMVK/Ve6pJBP5q
JGQ9tCj2/3FMX4CuNEqhWzNeVpOcimXnO4Kwm837lrldBWwYm7RMbJeV4k9MPO7N
xkPCmsIQN0iQb6bjaTGs2/MVoy3Qy+t6d3OKikhY06OKmQUlw+SvWZxi+v04462a
/+Es0tMu7WlS+N/t+RKseKeCTKChuIx/LqBwzQgTaxBcOnMb6b9lmE0hKUVaOgU2
futQ4mKNKyVpAC3avtA/Lk1ppRSMT3HsiDacQU9YldwtUuWj60Wzv5ZqsoCk2Ny6
QG11ioQf/2yh5eEYg/N3nCUR1PYJ4iBK/O8y9pqErr1QdAPxTeG2Dfq4bpsujXpe
m0yjMRnDfms+x/UkZppBezw1WIxX284C+WXOyQS7aB3C4qja2hRBlYBuIv5umF+q
DAO/onR56QBxuaF0MyfyVVKUkmvzuvG8tYivZdCi0l90ukxrCui5ofrZ5ZtahncH
NniITUycKxVGa44PxhvOfzJ+gGRY54Xr5S9SDj+fVSH2IVrPa726+/BGmA9GNRQa
nsJZ1hVL/SVVks93GNTN7mPqRBQ0j5FiWmiP84oCo1wchpDe78DHiMGY6YIZ+8b5
uBBDpmIEgBBIequxf36gOKJ3+n/zrHYDAojYe6mYdOHYvzQ9SFXxrRwXMsBoQEif
byZR09Dxsc5qjCbwNQgFbz+ekbhT4D4K5NjxYKtT/fCvc8aULOqpolxnVbf7pVT8
FaGFa4PZaK+FoicRbb/OKKzclQJmnjnt/k4koOM4A3yl6R983IF4yfiY52MrxgNP
WVV0Y8QW29JswaFwg4rg0jUq9wvBCxcuklXn78F+y3JLrp2e5e4JwLcUx6+S3waY
7ZfiXKNV+981XV7V0dJGBunp5anAsbQGNUHAEXWr3XVHgroHxbNKhK3kwFC8MgQ/
HyoH9goj/rLhSIcpElAUsbYkRV02Z3Yq++aKxtovwkNbY1oh9MaVwVWpGPV5IlQO
ac5juMJ00mct+woip8+FMWKgOPNn40nfVYk5XxCir0SWfGVhPjTHcc5RJH6sptpH
ML4rKWRyKEsHRZc/XiMkiOH5XBHGzEMeGqe8+Hc4ZxIPFx1ERquL0/SjfcTZ7LXl
ZzLYPS8F72f80k/Qg1PNHy+Bk5juNtd6qxUWDL0haBXZlL9Cz2kk0h7aQhAOPmVA
pyPi8S+XalSIJeMgEkv4Cm7FGD4m+Hx1R9J21Ivw9xR+ocZwKwjO9rgLRjY4zVQk
Gs8U4bS2qjMP05hikYw3Y2rQJVCQFYEnBcsAqDz00y1FZcEQNaoAmEsWCU55FVQo
vYGop/wJfmxusikiVKARPVHmJvR0XMKMF1WinbRW1OIAiXTdAG6+IuAj7kVFcZZP
/IKTw56kfm9Dfkck5e3ycXG9oEp5FMiUjfaS7LYXmyKQw93MzfvzfP6QkyOTLrQq
NJHRxoAuYVp9KplXH8s8ccVself0F+q+4h8A/Hu/cloX7/UUGlFGxO7bu5LU8GPR
lW/yLOInu+h164VIDCmYlO2CvP1fwP4/5zvcPWatZF+x5EcvcCForRJ4Jf+sBL+L
Bqy5RYYWXAM5vORKba+K8OhS3293+VIUz1pxKOOLYovEccTrq9y/pIy86BOSCL4F
m5dirIItj1xuUTjC8Uc2HYLLXsxK89WEzziHLJiS9xtAtbtpyLjtNsOb9LN6ODc3
LzymocPbYd22IHFRBLbJQOb9wAhYW8z1IpL5IPn5phEIhsB2WJLaWEOHe8L4qEMe
j6SdJ58u0G9oyVeOHU+E3uppbxg1USdhG+Ymbn4DyKVIThOmE/c3ou+Bt4lgk4z9
xCqMmH8nBRf9TndhAuc/Bv4/kOdvVD0EFqP7Fsjpo9jtAvsSodOKBJLgAsIcT506
Z9rSV/ERZUiFMPkql2rcGtO7UCpDYigpaTB5UW1U1Y1O+1NaYcRmvO04MP5/Sj0M
99lmW8Qf607W4LZie1KXA9t3xbOWVvKliK96yZgRVeydq0urj5EdhcJSHXjHAub6
sVEGyFONl0sHKsm46x3YAsL9BTYwxL9fYVvLEcJ0V3jhRWG2RxE1ppz6eFw5ZhTY
PLNsHBZ6YbCydSJHXzlelbB9gXaIgtJAQf0nwGvBqZ6siZaDrsyQf4qt6oTiRhR2
3481ItGKNbmwDWs4EG4OpQlApnHZqx297pFPAAv+M3jYmyggC6gyzMf0IBJDIE9k
ZivCPSaNLLG4a02YvRtvUhm8p+QbJQLdfvYJdGwqPsogCioVP7emqPd8TZhNpqpI
lUH1uSAldawx6MOiJ0KpcrB4TWjjT9S4tv/b13fx3pgeyQFoVYVeD78EbE+7cRhg
DFo7w0InPDBZG30E5N8Cc18esnRPmgEtQZPNBbggCQm1ml/t7h4AdaCJIdQgd9aJ
8NdSwznBe27ZTCu/HB/49JOnfsYRHFjZS38vNdhqLWQoReuYSNX9qTtPlTy315nE
tvPKF7NpPtczopC6A/elq6JlE/bQS+/doyFVZd3iblTeRpq9/HODcPXdhnVA8sey
JOB7ztqdzY1Zz0LqrglJjhqvrfCkENwGtY7XXb/gCntfXAt0ug+1ZOnCNcNmtMyn
nHmF/UnSxutMLId4viGaDJCysH1lQdbfTLTQW9BpW1x5gSV7PMaAHZ34ZQZJw1RQ
GFxSzqonmQ2HT9Amt0L0wxMwEfC+0b/fFJ6Au/bep6FAKfZ4kYbc/XYjltWWabiR
4Iam/sKoet3nsOQYue1L436U0Le/bBqTiWsWMSfBNuHw7BYxRSnysy4c6iwWpaU3
WtE/FRTykaNujBwTCK+Fw/Tv8onY/hxaB1OwVfWGH3qYaMMWnvNVay2OmsEbf/t8
Xj9Pm6RL+OybXN+I0XfpGDqVrjPjl7CMM1DWpH+bHVmTUjbvzbRRpQ99HzZuMbVR
liT3n8uc3iC506oF+KBEKWytpodZg25sWTdT3ywstXwPjRqtK1ju7Af7LteofMNV
ckFyKkvSh+AtSwIia+Lf3eMPGNbC4ZErGO4u16Ww7rV5Z4qTIYYoeqaph3BPBv4d
0PZlityd/HOMHfJNgmpYT0qXxwgezWNjsbmbR6LTqo1DDg04CHcR8SKAIukkzNbo
j6EYoUiYkmSAHbsieI5WdBUJuGxnWrBDP/fAIKKT23KL4ybMsjZPBg+BqqwN+Rgz
10H2sWEsErTPNE3ZSeK0pTFLwWpSOoZtb9lNItKpyPK5AUZtRYAITo2kEfk/lTDs
tN5c4Peu3E4BYB45gYobQAttYyimAQyYZQlB7Z7V9RRrYox7m+V5geApCcglBOh7
K794a+N62dDj5FePpwCFhU3Rquq/27NVzQqfkh86K4Bf2N+DQwQTCh+BOYuQkZbB
2mBmLJ6enuh6lKOULIymL3PJIMHZ1j1Se5tD+etVLjC/Hg27O1a6oKW34ZM7HDR/
nZPjxjZscgAQcsTqCMyKTEx82zMNQDsl20sBeYQLIGnMsYjL0ZF8krDiKfJrBnco
X/ki/v27w5eJni6JqX9eTocuMYGa4HcEyS7II0491xC4a9PFVOiZmZnYHNstBcV3
Z84GekCna5jDuKDc7S6BWuRJ5m4w4SgKe8iaXc/aAyk31+oeAkJAFWN8ym51ueR8
h0KspojHS7LVBr0apZQJFhHaCnWcyp/DoB/cLvtUaBOa62jGvcsxQ+d11VtjL5fM
a1IHqS+mbDCkONUFobpRPUMUlXj7aEpkt7ocNw9vuTB8PUgpcx8l3IT+q2A9hmoK
87CZrXuoVpQw7xOhp3kt8Q/oN9XXWa/HwlY3ytc7BPyKTIAqPEQjtOoJ9dVQoE2d
ZyT1RjvWcYgmmefJalWuTuV3UYSKaCEJmJWwzo5U3+eLNl+5ioQiFieftY9U2cQA
4QY6W0mA1QVZ5jjWgYb4NQwt/yy2PyV4WySa65cKiMsMknh0PYgLo0e+CHRk1Dc3
7dpAoFa40wl9xTtV1l179GVtCqZA/NOxWclc4qxz6/VrAZI3m82+heJksYkohtC6
H80CH/3Arg0nhUUzV+1HTrVwKbZLrD35CoYPBjTzKsOEgA3mLB+Mh+QPtHPMkiGx
bGMn83pghE8WhjUftNe8/rzWoGobO821pvZQBoq0kbi5RAITRkRMC02qhlwWPHoH
nMT6FeVUTjaOuoeOltJjURNJo0CewwInX4sh0ZLMKOYb0xVl8/CnBlCWG/EcU+Yq
yYi4ZK+LwwbhEysQ/w5gALJdegaKVfqfjjN5G086G52oe0voP6v0b5Iuz2xVYFxR
y3HvkO3z7UQtvSt95k956Nt6jE+4CxVCDx/YcACcQrg5V6Tndko6YlYFCcUvuNna
cV0rdPyTWxRR1dip9xeUt5DAm8jsTmyWv8QLKypEJM5GdA+dg1Nzoa5nmNEktLRb
QA5Xt0vi2JQH+jsMbisz93H2WpbIUlyHfbYvC8wtkZ3ColHQ/X50SylJiR8o1duz
RBoBkh6+lrSrB7F0Lax0CTd3ZVltPInbatJp17rSDOTD8qPMi/fIgM25LB04wFa9
b1F9vN3kbuc3Q5LE0a8jMp1VvzEoPQJnLgk1KjJDBu0IxZA8Z2EWuejLXreHiwm+
BjNk4zWFDDurObv73dcOxhmWmT5RZO32PzFCbUDlNFiG6ZCS6OkvM2VQIwEHLraZ
ffJ3A6fkJZUBZ2tJodCRgQRmsA2XCA8DP3onSyjQlgHNHZ02Ia1OT68gjF9YB7In
rdHtHI+rwwcx9jt1xqv1ddJKDZ8lrZWci6em3IaeDCix4QMK5COKWvhUoLV8T5IS
lE2Cdh+h3hKUKlo4DjZWX9GGo3v6mHzxNyMs7FEAOtQnXGLBrVHf0pOkuFUFHGel
L5K5Ere00xLeNTQIi8kyQYQsquunAT/Eu1X3dMHMoU/M9US6CKu6d/ZO9IzSHKwh
ycbkSBfisP0nNptOK2BhLkJQ7tbfl14wofpTjZqeEFKyMnzTQZ8HDixl6KGcmW9k
g5vd3ucxoZRtPKL1q5FC5FQcXCn0G5Acy+rZ8bUL66Fi7gvLZXAi3sx8/Gnz80U8
KgMKUSHwTpL8iGlfwAl48tQKYeLIFelJuh+3WHBaZ4UIyPmBleKYJN2plghhTEjS
9jXSfboCjaTdMWVXbB40mrpFJcrbMVrYP0uxDn+uhWfDwt3P2cbEm5VXC3izWgfk
TfEgczZKWC15HzjGZn5BdEJxoadjkMZnPjd5jcx2+6TaPbrYRWEEzd6EO8RvZOb2
dail/74CjYC2ddZ9x32g/cTz50xdpoVn4OrVjb3PtCn3xZyMxeRNh6Xveodn87D8
Gq3zKF/SVSts/dKPVkMCqJbTFLqzOvoyZ3c3t3Kckb8tpcWMwEp805+M7PC0LYmz
wK2CCnAwaHpnsy0YjrlP/pfult075f8Gr4YqAYG1v8UFbTSIEcGqoIFcXkNTVkEc
3J7DvZ6iZUHOt0VB0APJYSQTpZrddEyz2Zno4SnZvVAoBLtfwt/ALujQDMAdY8al
mnNCJz+pU1+Axa8mt88G5oxbHZWPZFXDkYJ84Pyrd26TrZKeii1CV9faaVbLs1f4
XjYEfFSei7ALyS2NyMVENDGgNc1XCuDsLEB9qRJcuX3lolS4RLCsKSTeH/ra35zk
5RZVdeEdKUImKoTYhA2LRmMVkdQrWrLlsfNyM2OOXuo8dvwH3M1WoT5RhiTZvwu8
ZUUxCzwBonlb4dkZMjbFcoyw4VY78qX1fCdrRKJ9kxDfpHejXG2NylUUtrl1bPnQ
Klk6u4ZbsKjQhwXa2iGFMmMDits5cXENo1A875PRHfxvvDTRS10xrHOK5X6p78BI
QjtbGDne/DL1GdkJ6Nn3C4lH8M6SOid4prarb3mbdYL5V0RHvSh7ghkzLBiHJMeo
YJXG8cTZteVH6L7tOrkOFaRDB2E/VUd0voTQuEqS09pnaVyFD6Et2/f3Yj4Az731
UcgdYLG3+OJtupjDKVWSIYj9H22qk0pBkIZflfACT/MUO7DnAs+J6axWLTVnx0sF
q2nxeeCNm1t3dOseoE9C+uM4nwGtLbpTMNsUac1DY3U3FLmJw59cL7VAkOL9lZxl
L5dKLgkWJaTIpVaWjx7GN/O/iLrCWpPUSq7RG23Rqkf7FTqj6Hs9ytbXX9UKvWn4
ye/eO4yETM04/j0flMVR0GFJ1UzyUiQ7xbsIBZtLs1KobOYMdAcs28Zq6Rl2D06y
M2M13Owe7tyu6t/heyk2RylcDQ+TpLIHQ+0wem+AIhzv3e87IO/oXsN9FM1ro2p+
XQLiTgxHl2dIMYjCEtL6LpTpdB+Bf+O3Ac5ta+E5YmHZxsM9pqsPj3UkvoyB6z2u
5nhkpaFT3SpHaIM66FWjUjypPiGoRy9C5TgyRQDnnLNpQZi25R9geWpbp+Jbk0Rh
Z8k/yHtbMHte5k6rwO4eQabZa1QLp2cQ9z8/dhOgNyBVrkZvJq01J/eqXZugvyom
K9IgyUT9xkH7g8G6v6uyQkicrLg/X3RGHbgLiKNOr7nDfdzDdOaIn+BKqXMfwTbb
9XBJprCuI0bOltvMzB57hVnkAUhsxjojL9+3u9tSvLk9EDD4/nUI8FSa5GoRVzk5
v5FaJVXx51YW6j+kdLEuqUQ8mVwTKkerrTMgDhBDn+BX/EP/2+/mxtUB0hzmOVU2
/hICRjSWLSfHG4ztNAPs6w8movtXbTmSWyo9qDMpLLSWg/CEAYIEGSAJL1qIH7Ul
3Lk7snoAtWZPs0MPhTCLFOLrVR+/dMqUA8HM6haEDzHuXx3t19ZTMHVwFUKsNTlo
qVuaTr6Xq15gC7x7JTnRSlj7igspsiZc7gOMsmG150Ot7F0xk/6vthNSbY/p2zG6
xNTukmPamDrxIs1nNilQg7TD1ADmwP2HTQsUZYKZcMkbqtSNsjkihaZG3HM0iB11
X+bZoplSaABOJs+JguE/xkJRM3BFz+BwLtryWnRygJomTvaU48QG4y5gr2aLdvb+
X8+iODXiLR/QoahUaa818uRUjdKmdEpqHHtktLXKwuWWakJRudzDnIzfIyP+XmMu
Vef2lIhbTZyYLr5OLG1m4JCO71heQdcVF+BeuDVTVcw2GljtPdWz6tBngT1WLGLn
f3n3usn7Vn86FF/NqLlXXdvll1dSb7CVJN4gNVUhhModRRjG7BzFm6UHQK/Fq4sK
DloDSBZcQ62nGMqOwxuNyvRftYw+IO31FkjVVC21bEL7VT1Hc62Yd1kqRTyoNjS7
2HVHX89OLEHMyOa9JhUO8Lx9YFSOxm7Nk2FG3/Cb7fjLFRuMsLuG5RwumeVlYdkZ
EccvNH1g4tYaBtPysZf+WHOnW2Zg/X+lRIyHh6UZ7EpsN/zafSQB/Bo1K4lwzNIZ
tM3x90uUBLiXGzF4wRNyBLb9xMOu1c0xazSH9yr3keIwHzKeauyOBgWCT8k7Uf2O
612GynpjzR7uVNrgqF91cr95Y8tO6+9bENt4qmgT2fHLLfqtDz1imM2MfmsXW54M
UvbnaQk4c5Yfow4W2sz54JCUO7Js6sNqXNrHDmcyvqoI2yekqMQEsCTbe4n2tsfw
C+TL7UfiqWqxh/q1Eu0sYZz7KP4urvVhFvLRIPYEKkPxj0ukyv6oEDyWg2DlosFz
Ap4OXi7ek85YStx8ehX7uovyi756QQ2LvtfPF+dYTpaK9vwWh1gPM5Ip5nZ6Q7zV
tkbtJnD2ldrYT26b1YOT5k4pAeL5UAgxuBYeD9wKngKY2LCnTuaH8f+bTX5qwfy8
LGehbYP/v5dWMO+3zInM+Q6L13BPeIQR+xcdfjjNA9Wvanyx8v40AAvfi9CpeJ/T
IPaZj+2e8caHR+X61J1q7E2JAhL/hPDKslKGnuWwAYvpJl2dmWU63vs2EL/lJXAu
LOfErL/SCioajeczNTEfbTF8plVoS38qTZNWeaaElT9DuqdnsLTTk1lyF481y/PA
h7NyMvG4IBiSqbNn4Rk2/0s2qr+Wu+FpsgjhQK9k1Jz+Ql+I1dB68molcymwHPsP
Qe6Vt9au6/1tT6h+q86Cssm+H0WHLXEZ4RgR2Fphz9hoeS3lAGbxDYaGaKcoFWQk
xVs2Fqfqu/qmpwahM8KBc29xyW4e7cvo1mDS95bPHYwSETtclVHO0B3ApY/qKXy8
JbnDp/OJBtcV7Jie+fMcMVz99tTf8757FisIIr2dMjcQZe8k0TgiWvNYM/sEjHpN
Q/Vryl71TVHJquX63PIHH/TqxDLvXZsEpk9Fpg3vORVR3LWdVpCUrSLpxV5MmFH6
jHaEoaqsp1dLSwxE9xEgVWnwgs66LzqAq6yrVYSnV9QDBPqaiFCR8DdlQh4zpzHY
3LzVhWz47k1NP6iu3geDszqxzkLh/oOE5oA3dvg6GveePrh2aldssOKhjf/GgLUO
K0kIvN71qV7insqJAJtnUns2pGzpnQSz2Y0T6APykPUropDsuk/eizS4MJLr53xR
52B9Cz3ebL5TOmXhas2CYQEqOE7w22kCX9Vj2ZwJDGV9UKFlg1i/M2CW3twChGlq
5Oj4m/hOeyMc4bP9x3OhnrXLBpA34uhkWSFLufOA4E0c+xP3j3OLjVzkGRWM8cpd
hpwhnf3UDk+nB/dzOtLTHz1JxVbKrVIOVhhV2rdbBFOQYLsNRQeRD0+vh/aMcqZQ
0G5F/bHmOFDt2ugY1LBqrE6EW5jY4SFJ4QRopDjiuVYeK8JzF6+zhwvJ+h6f5HGu
kEtSoy+jouVH3w86N5RzcRrg/f4M1JMC0QreXsieTddpP0pg1/km0V+6E7xRZatR
NyWM8RgCUKh7cLLn2gNAyMbnYbFdr2GTMrWbJmGgFDpAxKm4WmhhgwfEP1X0t5Eg
g5Tpzbo/5QPMq+ErQrgR4CBesHXht1U9jYTJY5qAy0nJQ28E0oB40gTd/yF+bNUw
yX7FfX9FHAeawX0f5Jj3/Dk2aAY3fNanvedkicQz8TlM/gSpAC0moLA+UkyrfcsO
YGtS5+VaPlDFhjhX7AWyLwzxr5o+rhHV/KRdxiRq/FjIV2Vi6gXpbXBcg0A598Y4
PsBoc/ldPK2TO98PxqeSGjPhcRgoUbfrC+gIXYfjVw7IadwV0y5mwfrYG7Qc+0DS
otWghHJIcr9I/ZYLR8rPPnm90haR7V7eTVY3wV7liJ66Lm+QQa9Kchthi+r/3zQm
VMoGRg+Hg2eIpFSvY6WWi3/bg5FHOfxROhFr6+pCswf4ecetzsYupkTXiz1bl/lk
2PmQ2jtTKfa+F9MclgaRHsf9tmLF4uLctNTZZFPjCe1in06ibBoYbpwFIYdM5n74
f6d5ERgUEBcsUPyO8Dnqqsegfoe6dI8P8l5oC92mVkrF0bhrCrR0BGjEY9LRShR1
vf/MSCN3fEcTmxs8lSjp8km/k1ZZzRToq51n74y83TuZKkaCNdj4t1LAgLt506rV
lsxFsU6GmoS8XIfUJLJ01Yfc/5bD1i0ph+GkM6QM/BK4ov/rv+D4rKcyBXwcvqkt
8DAi+fU3KwtscQueHJXK/5MRwSY4a/qop3IAT+o25fZiRc3sZgfViWkIVI1+4fSz
jKR/OkiujeRN8cn0OpsyB8WoTS5Yhbxe8DjfY0M5hqIjTkGttImf6u3mqCxCPcAo
s7Uer13HTgAA1XQ6wHfpxTz34krwg/NchMuoGpCi2WimsZ5pfTfGaCgLlpAPqKCw
FsJxkUwwNw3le95mEVfmgKK0ZC57ztOdKfs+LHj/x6Oum+NpT5qVHQxrTooDiZTd
MTFjSORnLRNElLubiJqoEtl8wSKTTnXjEdLhybjUsVIWxuvDRR8XXpCPchY6Fojb
Pk0WmmecXP7ZLMrPm5B8vyOopgrIMcBuRzuGmuwdFUaecymQuMwXWZ/P2VONJwgt
EcwDKl1WkiLAgU58XM1pITJ8z+jsay8SUP00qnmOtNuhJtLEzOO6xjn7DheTpgf3
8T6LE4lQ2ohGLVG7Bts2TMudLVDmWJgMdzBX/aKfrH0dpfkrrqLlHkWs63p1gnDC
8IvTPF2qumqbjvU/rKf5db3guTuLdGVhKBES+mxUQZL1ngQ1M06cQ52elHzxgvOx
RkyxNGdcU1SoRJgB5lW7S2Xhycjk44d1b+Qy6FQ/NKR32dQr/2fJtSAVHezr4BYi
WgzjxwjSQC7H9HcRg7OIWg5fdettNeOFWvgyjKJczjTkXfTT/UCukjxljcz2uJYU
pGfnhrE+fB2npFkt0JpjpdpMOntlN/Xm4HKhrSEy1ZOAFkUoQFMO/Emk4pzwuM8M
NIcJvF4HbKqAthlCb0DAC90WJ3xDuUN7XHP38kPpwcHi73FpOalonzbZd23YV+R+
r6v4+RpEldZOx3K4qxtjs7fUDCYLP2c95MNayPaaGhWI3AwKNGQF6Gu9BvRkI0+L
IewuBX7ZvaRsDxaVSjsLvOtmXD+T4S8xj38bhqw0M0KiCZU4XB06JaWPhGPi3CcN
PFwX/G74x1UCh4iny5Zg+DzEdhSrIS1iwMIZLjh21aaabd4EZ/UnFcQ+9hnWnExu
YLk1ppeNny9jauKWQUSoIOT5yVdi9/s67LM9MrhIGUhqm43b5LkaJK1NCTAKpMfT
LU505LugOy0iSZbJKEo0sWrboF15pSy23q/Lx4H4E0fiPE0bp3s9C8w1X0o+nqtS
B4WwNsYU++OAVkKuHcIWi1uPSE+oYyVNoFJCuRZGi60h7FBFrBVsE1p/BPnh04xO
hrEAoeMP9cza8lwkS5PWy5yb46KEfpQI6KC3FZ/3+Up7XwTN+QiJEo+G9aCYE490
Kuhat1MlKLJ3EpYVNd4s4dTflhzUE3Nf+lv67iui8oCywPxT5VAHcjlaqyG7Meno
u4akX/CnSmdXGgQCVmmlXU6OTTK6gPtiYbhWz1fUGZj68s2BA3ubxOLrMhhIjgz3
2bed4fRfO0RhqDI15cmsyO+kxj1kkPnUGMlGbLzNRwqlFEjf/kXQY+8DGODF2f3z
VtQ0ZUitXZ/oMIeX0IysQa1jjVZlqIDXSM7K04nKuqHH1yOScH8eBBhocERz5EQd
Kir2qi+CeMRIy8Y6P6TivvgGJ7Jyd31IhfMX3ofrygR4VIHkjhy6nAzYW/CoOR3l
h2OEISQ/vEsp6JXVR0Z7k75U5kgYoYvqH1/ZjTu+TznqTPu4Q7HDpviE0hF8eoxs
oASAyow7AvCsIEhnVfyNvMS4huyvaAEBlvpCsW2Hl/HzzN+rZr1Kas0CreMdEluW
nELP4erp4/6ChaZynRkjsmifMr2SxQipPezpkTFyHwOx3FqpXiJCm3yE021NiZdH
9k2EUS5fSoNnjvHNBBZa49M3wGEMatDH439FtZacpkM9Q7jryNB9G/PdQhWFL9sB
YxMrM5mI0NKfCQA7d98E2kadvf+1tL5Sn3+F4TcdZ7oC9aPEYGOPX+tE0F2oQKVv
JZ/fAvnBH8ncbos6XsVPZkqFECSK+iFfyKXMCF2nWe+nL4CIYCtlPPKa21Rz+UqP
Fmu389quhTildsgMbU+eBH2G5pYwsG6ssn8UqRST4qXQHoHVLFqMZvi53j9Z1hMc
XpYZFXcBojiV/GxicKC2/HUv4xxzHXYf7k7x9jh4Jq7OvzV4vo153+65MII2sf28
B3KIiQju1y/lHCKNAdqx1bSGnyuApqmhDn4rCV+p44PRMJGRKaaMj7jv1T/8KdpY
p5TWVW9On5aN3b4Y+l6sMNlqDEXHCD+nX2ywQJwRMWj7ENbUbWWu0PBABOtKeqPb
LYLg7H0/z2BxG14lzkIxpEcqHLZPdCkLwuRNytnzEeB1A4BfbgOaY1mO06DgIWPd
YEcnVMm5H3t4h/381x6mxJqp9nHDr/p+dkaJOwawXqJn58zpheE0H0f2M51PoeC1
IUaB7rp2R+lDPvuuCvzF6veynxOnu6yW4WfinvB8SYwOMllynbwNnpmakLtXNKNP
FpAS6okzWf+oANH7YnSe5tgfXZVDk6n6qGiD+6esnvDPXmzZgsLHkkJEpWwoBIdW
iUh9dmUTSWjx0DzsX1B/QW2aBHJWF1PU1RO3ORQ/gBSHdYbYrxJF5yiglCUEvEen
NsYyYDO6YD1okywi69VQ9fsRy0uuOx2npF/IYWfglDdSeZ8GsPErEkGQRqcJnslw
v2t0LWrrwCL+TXLodtNDkf5tSCNNKk1pkevwUC4urwgDGCSW6HIiiYPhKwpeKGQL
kznXmCwJ8JIosWqUlDtXgxa9OgucuDB54X8OokMxAfWR6K5gP5hQ3vcftK7J1zpb
QpyTTZPi647qZgWR/BNy7FmgMGSHP5+WqvkxB/9E3ySUyhI5JDbsWhVvxwzPlE6a
zXs/e/tPMVTz4/vsu10GRycRfLfJk66YWn2askiP/F2UabcDPy80rp3Z0mWD5VOK
XRygwCsN+ksMlLIyHjLfX3nrcoEPJo759uycD0U8X9s9JHkonsu93A9IyfKfe2/g
HEVjtI4s51q7IsUOH9UlGfUt1/DlMPUbwDtK9KA0fKsn7mUMXh+Ezb9BgoQru2JT
xatO3SWK8iam/Jc0BK5pgQSYUG421HBiI1uBJeHXAZHic+xC7EWJZ3m4EV58KTA9
UHns/56VAONxb5EdWnjAyIPybf5WjYR197yam2elFPX9kr9XPdGbxIbaxcWX6269
l5xQcTD1bHHn9OYfTKl8UA1HpUUeV04FdTVBL25aEuuN1qEFnbmKMOrtiiTbuu7d
wp1SbPiczKZISJ3YPPLHjpZCWZfVmkOA63UNWbt4Yt7pbDr/MMWccoZlOsELFH1f
XCmjE2bexpf/m85t+5on0XhG06qMYxfdR83i19hvZphTuw6y+IF91QKgF3leT31Z
hjesfOy8W/XR2d4R2SMgi5KgHATwlDb4Zn7awLoxeEFpS6CpnDwOgVTyS2dt1PwE
gGFzMpmcYvqUr0Nlrj6TP0Ci8n68gQTW1QhM2NbIZR2VuQEzbxOiD+IsmAqa6Ns/
g2HFp47K9bMkhtrloSfTRzl7UZ6Kxtx1uye9KHVcgkkaL+82idKF8gsW4TGwiy+L
GBFumgxynKGJRjrcLKpWjrgjdf7SCIaBIiRhKVZseLFAQg6dTUkKfiIXKW4r9Uwz
2/KzSWD3cqVFx0mTwoEhr5yBydqk+7VbDwzEF6hhocoTwaIw4PWnLqlQ25NmjEXY
9DLLhfuxFyShAobIWlMcEsxbk+dWypwz325PQxbGngQv9rniUncWMctwyj6zTUnB
5tXNP+1x7x13ND+WUt33KP6MAysQdWVJTHY+Iao+S5+LHqutLwYIiaZYSIOo1L42
Lfj7OGfzdJNgWJi0XGQm1qG1VWH6//xOJ+9zBPHogjqdnwwZOZvGf1uOP6M25WkG
SQLwhPo5F63qJ9dV5r5H31vSXV+3tYAgh/dem5wMN7CP4/VMxJRDYaPK5tnCLSqX
k1yCvPbrJ1JnEgs6Vs5vSoWQ1oduUYTae/EM0YzjRa85oyvMfN5E6QXSOCGRmVwD
b7AEcMNx0t3HE7Ma3UPUycvY5iLx+de4mXgnch/McBKkjhvYBxD61nE2feq4j3Hx
JxdSOBRtx6da8ujJ9YzFZH+65wUZWwNyx4uOk+eSlm0GFE17OkddI13RJrh/SaXm
lkpjssrplRrVQqJEp9iF47f3jsODSc1uoBr0rd9xhNDrYJ+uq3RXYabK5vFR8SIK
WWU9sLRCKKA4tG9qOUKI9rV4d6XFNgTgmLAj7sxsb3sn5eiyzPWTtGM3B63ol5TA
KewnkOIUyPV+JtAeUrzKPwJ9cCTiwmMCWHAA+7JJ2Gi8Gl7wDwOvbkp0bBZp1mlg
z8S5T9wAHvnADxDFZvVepAGcnFlFkE+iiEW+XaYL2oSjstLWQp3NuOGIFSVL43qX
cfhyN2zOr7yEHej5R/pUCZY6JxBX8Bm116AW6eT0jNecD4bN5T+F1V2kzwHDtWPg
wpzmRSHRqbuwEoFDTZf7RkhfRgtEeAtIPNRH2e8yjMNO9dsNRP4gqSeDPsfEB/s1
G0pX3J81UD6PidRXKxPpGauxGJajoAxLR5z1etI4KNYJYGw51FcXahD6tfXSQeY8
zPprVJjM7vjZZHc0xM2slO/S9TrZhYgDrEv2lW3BUWIjz3XcPvZVIChdE6L44Ux7
KM2eeEZJN014sslM5wqT+o/xccBt9a/MM9rV/75d37A6kRIzJbDSHHkcJc1rZ87A
iPSTGa/cG5IKBdDZUJatB1dTMsUjW58n/1JXjzQhagmrsjDgPW/6xXR2QrQJMHy+
8BONTIKx9BMm8tjFgSCdZthlRc9321E7gk6ouQTsgDFNrS1OPlLy44lTFah/hCve
IOjSz58sYuddLpdUhWcenPoLiSrHfTUABVBPLrkqOUI3ZfHA1lBVmhuBKwsRC2LK
wkjp9PS9f3iERr5cWgMX656PAe8/hKaJ6O5WaXuyzjxl0mcpcRyHNjyTlmdlnNTu
E3b4eSYdC5u79OUxaTtNm0jTkJ6xRkF5KIzf8xpHvpk/bQSRL4cTV4SKXH2xrq/i
+M62JObkWq3GVA1/RSmU3/ywWCCflR/KCU55YPR4A5VYxBoS9OFfKcrDj4DSdF9W
5q4vJadZaJL+KyE5mFEynvGKusDHdLOerO7oVCnybcMwMx6zo0rZiUWC/dBi5pSd
1kfGgEjdXxjdEemocpz7kMULYSkIKPkCgXxIVBeqzYXY1ZjdRWzfkYhYC8RdUzl7
mJCe0a0lzoZPWpz1Q9zVf4Be4m6KhSCiKPTrTSJ6jCV3yEzuYGWqMTPAyxX6RpWO
Qfws7dP0Mz7fJLfnyiEL1gTwxU+1qSMMCNZ4RoE2viQq7ne7UnEvTG0ESYTQ1d0g
eavMs72p+1lnhAZsYWkAOJJ2cNhkfPx4E04Sg4UItc25I5IYPBlIfFAkglVlf89J
H6fEyeXrBa9IUsbeBitOUez/r1pKUM1aBXGaYVv9Bv48/UUAax7oO0mlb+t7yQQf
LnQJ1VJh9na2zyq/OC2Co8P97Qn7OlSnGOZd/kFJjaIpQnDMX0yM8XvVg0hFNTJ/
jWZx3IkMjy16k3cZYGgd5RTX/gjBE3/WDkaEnz0yOuefvzHzzkdX9hgc2ror8P/u
C0MEpB9wJ/u/NBgzmTcJJL5ND/dDttRpOMMB81JjqzxGCbSj3rg1i5+pCoPgZ2G2
/T5pHOoecjsTUFLmFfFIaTYXVGPv56S/FVQ+Q1Da35MZ9ZGnk6V+CMsGr1X9sLmm
krnsbgJdT7VogM2aN3Gw3r9HF2pv+3K4BjyAqxot6Fy4L7ceeI4QAILIvs8RxO+q
vhCe3LTszdRbELfN8kC4UDe5rzT4Dh7GzxwQne05Z7WrxAcublLZ+4SP7A5rajU+
2+zzavpM8yUX2oomdH5dQyXjpN0dIDzBJus1Eoj+xUk+u2R6p4prVQJPn26ZgByS
v4fXJiB+bH1nTgC62flKAVYbceIXngF1+WkQd4/qMr7r0AF/jU50j2sOHBjFSSnz
H7M6+XbzaP8E6dFPT8HLtCIp4lOpJOUASdF3il0JNV8/aP01J0C1j293dmuEIM+I
0TFIlTG9/2w+555+fUe6RCAyW1mF8I1ea0A7kZRiyE2GsheqeEr/UjR/T1eAvUCK
8FuUN8etA1cH69rdVgnBUEO1OjnEYR+n3BEJ9+J9hyRwjrgJrqV/iRZGLfE5946q
/KARZlSAXu9SOGuP6ey3vSWG3kHDUgqHRcK0+KRW5t2IHroKhdvRSmWz50E8HjLv
UstEbasrPeFPAW7EvIVesCE35cMY6+jZmWXWKZ3tRWD6rigDu1eziZCMiac6Xq9F
/lXKb9l5zdJDyq3ofq265vNcllN8BMRMxajRf/rIDJHpXO/jMI3lntK9ZIUUIs+J
TasWPjQEW0YRtjP7M57inhewsL6AEmi7HDcrROXDhZR2gyb2pNrND6wsegCHsTa/
hdXv1gCP0sLKDriU+SqFqWE9UfA62XeOPYk48a80SPn5Kbkg0jFxnII+GdbleYwd
2g2i7qkJ85ROZqzGix+1objekHtky+/jyaM81r3HxWcMLQ7qkkiJrE/0MGrYTsyT
8PWv60lupOW37nFS218QMAQ4ZV73jwnx0BgP5Xsq/u4CBIMftePZkwfSOMmAtFoP
JOgKuSHVq0qbWt+m2FtJ2x9ZDtf4qwwiw6CeF9YYpffgcWdRb5q1ww36RJFxuyzB
Wei0+Amd9IIdNXXNhEL7tTqyyZ9dIxof2gjyxgb0HoAvdkhPOVf3NnThlQbERcFV
xs6APz/3totBC/IYwPSSKJB3hGCIS2H7SESQo29s/bdNN6XrkZN8gZygKJXrKmgC
aN/Bg2wvewSzp33oQxt+nfrcfh0a459uXTO48dhCj0qMbYJAiGv/afAeNegyK05G
eroXS1mVIMreLRsACS8cR65eM6yg0W7ixIj6cSzpnWGI73Pw4dGBKbv5CUuihGur
ujT0tqThph7gioxDVsh3a8NTlK/iAva6BSaAgD9daM4v3M4Eieh7XGAKTRRMCCUW
rUUJJ/HasU84Kv9TuGY/YgfuNVObx2iipEAJasMjJsH4zGItR1nQl2Xluua3KwF0
p69Y+iztWPmUwUKaW+pFSrdZLOyhCXxk72Wx0h+XlWneHjrdQ65Mv/EkcuTU5Oh7
eDq6r/cxyBZi2/8yCo1g6zUbOigb8fUg/b2ZbcyLKJ67FohhssEHoz+YrcmnCaS2
J9OEVoz1h5urbNj1GfFkh8OX/ORtUAFh1VUGug5fbNRdPggHH9It0Ss7asDzgDLr
S1s945HgMIApEpTN/6zwXHuv/AUAmeJFiSpaATjA2nOgxBKgqK9dGdyHqK/8Y5IY
wVIsV0xuDlErTpHHT06tN4Lo/WEuKsb79wVoYOiuM+g29Vn4p8h2N0YrL5G3NGzk
jOWdH3btACVuyvbxrvKSkNhcg6HhlvsOJB3ba6JywqfjttpfwF/36LtPV6UrwKiu
aiVHUtcYNEFN5Kt8c05SKNT7THdnF150Jh79KpB/zPMJF7kVUC1DqppateYnD4eV
X5X+S94F29OqV7Dqf5kLllt5UqU8iV2IrEYWeOoUnHOkKbbyPRZRV271Wu8GYhK8
qUiYoIHqI99jvne3uG+VowxHTxOpIl5pNSnn8i2WONHVJALdYRjshpxPtWCqcE2a
uG5anGtZIRaG2mhEIf38PcMDhdwZaA+gr5pwOFF17iEAFxN1fpyrqGP3Fmxv2EgH
xzPSvaFbFZP9asHd/5Q1+Xuo/AY1hGkyTiMsoMiE1ipf7FupKBuKPQVir/BSn3v4
vwbxrOElD+vMcZ5dwVKOedJ/eWGzE0EcAPA4RO1zlYRF5sF1WyoB7daXCmyEC3P8
uR5+/V0JIy5hUVSesHoK+uqwnyZ8hDOCuik3+xrCFFsX0+WzTc2LF+e71DejnUuv
llYhAg4MVHRrbrA9d5WTPSHvKwv62qAAN+oAGUiLFu2FZCnm0rcL4Eh/q9LBQlNW
zymCOJ0uGjxY6jU56uk0pL0/wD+odgDOtDIWSXQUK7XWjhs9AI2WMlHcZz9u8VvE
JKJxo5b989cS2vNkTdRhLF0fEGyeNtCR9xDVL8Q61+7+f3t49V+fruHuBe+sHrwy
x+ADsmDejNl299ooH7YbwvxLKEc9TcB6N3bRUJmHZyOyDJhECqE5wdVqrfTkCcpH
O75kzRaPryl2ZVd+/ZyjXqDh6ZNm+myJ2WHbdwSOpePR5cio+bJnxP/NjsUPgFdV
ATk6iSJhSoXQk5h/J+JDlnRKt0mtMIgsW/GNZhhsEybBHzkbt3Fz/P6mykguF9wt
hh2GgQUScpDfb5RjOML9WRE6YqbZG6iR0qNx8pWJZ5tMOld5VCXqzTthgxgldzZr
1NJfQFl1nAhBQVC6BVcZxld1TI7IOb2PLrfmuwuMMOW0/atf40ACmFofhbe2h0gb
sbz8RMusLx2pN4dgRqjWCcpT/qjDZe2FvfY4S5hE4jfJ3cYhUeb7uVZJPJeHYNqc
IkUvWPziGPV3nRMXVEO0PtZbFh8RVWyamMiqrrtwmDq3G8nl0g/7Vi1HMWz+z7L8
r6JeaLRsGx7WLoqjSNNPgUIygxxGyine8pMzqYQuIQeSf3LUp/k0RQP+jUwRIOc5
GFcvMXhR18yMe8PRhexhsCRjqCtnUpZ0za3ESfp5y9TPJcBMQ4Rrx8vjaB7Bzpju
JdkQxtA3wOP1cAmjivT1BjFHUrJPr7Lta7ruehYTKN17p+qQAaRZ1SFzt2HkSmEa
1NOoCMAOO569jL/JKLcLF9HnphM4PL8EyXCs53oTvW9/rosnA9PEl/0wiJl/xD5S
GK/mY3pDYZjAsy1DKTCNXNGeIVO/+74YtVZp+tyj+ZRSxQ3bqS9LghBEQd/WCsva
kqBmr0N3U3/n+hvNB31Su+dxbhQd8gVOZZPmAhAtq9M8YYWCw502qDthoqsJRsUD
FsfI5PXFY3i+BlhytWK4KOngVRpQuWTUpZqCtlhbufvfyNficZvkSuD7vtRNFQZe
3GlUiUTiAlDcQzUTm8Q179RkwscWSvCPrZ5yHvYdw5Rcv+CrPPsX2F1N4d+loD+M
9YUmCA+Q+VXxu2vOnbdL1ka9HKZ3+2zNN5HLxtBrJi0b+UQnqLjIcH+1nFpKL3ET
S/V6h6KQjuqtb8qduk4yGRrmHBAjomw5F265Hioqfw2MSoGTx85atrNX9eSbI1dI
rNKXAWVmkPmP7ieTjFJcLDYsUg6yd6oRWR+SYEgdWsUai6btI/NEH8rCzEZCccKu
dxs4On0bFxzH07ffJyqap/blH4dXNVeVxQCEB9fSdedUC0TMF6ZkQbopWyIsnv3b
YR4m2mkoRVgq/z5J13C9y6cNVHA1YCZQcArdqY7b9GFgcihLa+rcj++gA3FhYU1v
ZBaHrnBSIUG+EAZHB9NFu9dxhm1QQlCOPbrg+ZdrMVHAS0k9Hho5wRu/upEulOzL
ThvD2MrYfyYS4+qHkMOUX3ev/hLefN10KlVqhZo33aqi7/rqaWCUzzZEdUS0PASE
0mNZzn+NEifwh8QIiBf507NoMRuS7mtGIS+itfrcy2PcNS92vVkAGM4iOU96uHzW
2CZXxs0lsKKk9lT7qKM4wT58d7AUV7BSfXdoPRXo0WhgP4WytFxwZqbiUqMbmywT
WsKteYCgV1cvwKkXzPvuOkFnLybmo7WKkr4P6EP7gYyl5qqCdomQMQ4bWFW+Fr1M
24jpFN8sQFeAqVLwrsE4VqrBXxLS5W8GvAfoEt3nf6KRPoTjZ3xcASwd8ZZ2v1nd
q1MYVyVHT1GAMJohcx2TSJm+JxIioJLzvNLC0XBqDDyBf+4r6DIWjtznf1a9EcHD
/mwZeYkP62LfvYVVY+OWzIOB/PTTDPMm/zCZXDezMUMwyW2NcgnBOAQJ17KbKLcA
vPftspQXiIq+1jP5gPWnPh7CLXfzeATj/Ier5W2o8Ue+qguu6bo9OgqTdyiNUvHN
IzPtmTL0C/Xx+YWL1qkzj5r5VUYCOxCWz4Q5p94qQAPFobCtWEynkv6kuYiD2bHW
XQNg4dNeVJ6Hix2pxIsXipbQhzHCHLe60gffM3EJyVSDGPPu4AzSY/kPGT0mnC7p
4BX9AFymbZ6RAx6pnMIdqOPWdL6ZGmKy6ot6isHpDcczqcmoIVls+TFCuZC5kDC9
vhljsimlR/VSipzhy1IZxR48ApVvOvCk2PRowgpFzq7vHiAP21n8ZeB4g5tNGk0h
tpCKxp6wfNtR47lj+NT+ASSBbetlwC+22hBsTqBBE82ZQI4WUJhAh4oi1utqMSXY
TJc3b/JDlcvstX/BIViFQDkA9fVSh2acJ8+i8K5kHIYuVekv7hFyX2Zmr5YGuh57
r5YVkdHP1ZfLneODyNOleuclC6CTBC347/DS7WTcS5mfnUUpZP2uRbop4NgFSjz6
I+5a4awfX39+Y6VtpHokhTgAbMgQpYOCQ8qf/qz7wBRNPyMXQHmcuTv0JAGpACw8
rAz/x7fwFUtfaXBRbLFQ3mwpP1V8jO17yTBUPEof8QFslPVwYcbJGjKvyDHcDZKC
Uf0tFvB/aDlAHxEo29HU8VZez0daQjU1yZT0sBrTdX3na9ZzdvHbpfwM72ocUQsf
MFXgDjOOTq9ZiPZRaWhjR+HOOtVtcVdSzIgYPEOkC//mUTzmLFLK2eHuXEDz5pIF
Uhg9qblzlDRla9GVCyhszFgK+uTcxhZ7c/nd3Dgng+uHEEA+rZ3TA6nlVFhYwbon
UCM+jvldGglHPDv4tBCpdt0HHgSOxGxr5v5JQdBp+A+S/XGb6oNDAtL+22raBVJg
c29lqXfh07/Ew66yK/OF/Q3Mq56dUiW9dtqkDrvSFj3T1C3cjDxiZeNOCjAo9otH
OBJJCIFNOtBoeRoa8yNbzdvv/RIQTTC0DOYiftf7IGZNlE1sC8/z1RGCWIDDOd1S
nyaLcsq9tAE8wKc2GfmrEWvO0lbGg2E2+UTF8RqiagYiqUeMOYg2KHSGT2Os5S0L
q6YO0qIioWxpXkJL8P3iSYYEtaagMqtytfifYen3CLhpGTns4ZxnvkByWqemC4mo
hkZ8zcZTO+C2Gp3oC5V5SCPl8qeHlIumtWnwPxh9pBvEk8Ndi0b+zXLwyfrOOr1F
6uSkJx3uQG3AVuhVnD7OlqX90k4KHFC4TgH7gQ3MMtJkDQoxA+How+ucbYMV7h5U
KiL86SWjz+H7SMj3xmJebfiIeO2T9T539Wxe/kDOHETSmt0I6nPrx1WTUhD8+z/2
UI2VVv4gKjV+l5i255ZGm/PNWoZ3J1JUEeG0DJjDC3W3/CpfxxZsujM3WAOEzykv
ExtOf7estLsJKGQ0bgMYG4zkIpbi+NeSgiRAJS1fyjx/gq5v0h55EPu0dVB+SSlU
E56aljsqBjgLAyV5tSZO8hnH3KKxp4V0rcEzigQk+SYtikcHhlM4ojyjgjSE4pmV
8xuLDq5aztTrV4ymPfS8mGyrLswHFYDDPfB5ANKpZkYZbHFR2yWRBiWmBKzfbA1z
FkpNlGdWzgAWMcr67H78JNdZPCyUMosTjBVkFCu4wCzBLZGz11nDYEd+wWhqA7Zw
HQiN5XKbuI5E4+MKd/eIU/fmp80ysfLm5vd3Ut6Ql6lO9JxpQaqLeibhMLe6/3P+
k4ZujGTCUuJ78y9URG71LMqOdY6Qsziq64YT0z7YONu+gP+Vo/ANvGLykubX8DUD
u7rR89ZImXm3jr/KZKE59yKELEeOXbBK1Nfu4EM4q9nyc7Zl0sQT5MUSR/+e9dNN
653GnfbnUTyMGOLSIrK8Gyro3x6o0qm13AtEPJniK68Y6qR0YZx+GLrMHGz6UDPV
J8EsnZw9RGprElQmSe4vuYksww1nNdQLyifcMfQmjcOgxP5+uvguMe77RVCOh7OQ
JQXrNBHBj865MW6SWilDjU9Rro6HO3nnygfmRRNqkGuV4vrP9+UiQXwT+7265Rn4
9j1R0GBm1t/qn0XgAXXqbtdlzXLYPjrvLY/Bz4TSYhj3UNJ2q3UIKYp86FgO1XNp
SkR46b3VkNVeEq+g3OfsT3tVUTfJA0QCAGTcLcLmdZvz6HQxYd+/nGz8W8zJ0Iuy
2X9iGA3mFuVTtP/vsYOfBeKvaO7grdOP1AcVsb63xrS0iSFz5LSM3R5jqHRUHRZI
oE9HxGDj1ecqdjD0XpWxhtMYK3ecODXZunVh28T2DH4GTRZro6fXlMLT3v96amMW
cVGq2PhgB1whqaiUa+ydmrG2/YVdb6r6iptASpHamYk7MpiR5a+q5Thgi1IwI9gK
MCTXsKsmUonGvgcCv4xa0ClEJYzvfMuD+k18ptOobNgd8QZQC53mpkr/KEwN0H/o
eYGi0MGLSzDoV7waLyUohYYE7pGko2ipayE2RA0Sj5ppNGfzkG8DwmL7jNU98vLq
XvKReuHAxlPG6A9LnPxZiuloz9aVXsEsNm3qYIZt5XU7NZJ2y32/zkAWsAr8WLDA
QbxzvlegF80qQlANmZfRK+tLj41wO+La6p2iYkh+COQmcQyLgf4su9EJFlohOsdD
5saCtiHsVuwo5nF+eiaF8EG9JMeCbhIZY6h+GPvP4j/v9f2jtiKljM5fDPlkGJpb
K2J7hRNFa65qk/vas05OwoKusXpdq54bl5+8Xw0DnqXio1vDXH6v7cE5KQ2N0njD
TXsUOkc7O9plzOMrLkv2U7cG2ADUMWP2xQ3YHYPpBH8ht3/rTEf5A4ld7PgmvEWJ
+MJWF9kJSYP1YBhM+iqeweX2Pfb0E2zNyACwDf7D8Pybs9IzqHRa5FAtwtv7U4bc
OWaYVXmtGooGlIiEZCXUVnF+63l0WZ6/TyAjkE9KLTjC9OZ4ZuYTGHTH38SydB6I
dFgXub5anynVyXn+vOJTLOjY5zcEtptq0ewdhlyDesPe+pr2B7HGEl1h/M9YBoPP
roMolrKvofp3UPsfeHX/YvCM5na9pJ/HIISOQQyPJAMzD1rFMi66MvJ12WTbltrW
MxQX3tm9Fu7Y8RuDx2xOfqwIkSeuoextolnHr0hvY29ZYdBR//pPnr2joTL0jKlx
PcLdehJ0YlOEHv+Em4sl1oyhQ66Ms9CZDw2jSo/dPRgKvB4KWRc9+2OwnKJ3s2Nb
nqpQT194XJUR+N2BtmNKCEms+ftgQtQ+I2QLVaralrECKo6mMtHXWkiXMQjQKP2J
B0ZJSrqgE6YUMnfXTNJ9QUHhgwM+isJEX23/tU29iUnyWHJUTXsabcQkYtQqwl2g
2Dts2vul6prHyLF8QMHumXfDtMxGwxAfI7RrTX+p8ZTGVDbE2O2qiMONYRk31JIP
ehqxGUpj3wPS6tBVxBBchsRivKWbfZ8YRrCiZUMr03hJ53eDQga682+ffu2LApTU
ZpHH2xhZXoKbJ1dwW7H9fKq60gV2//moMXquUf5L/4j3Vz+B2XzVBs+6l6Ld5+P/
r9nHEcKjKvzKKMomEImhvYvm1EMzYha9N9HCW3qXhaYKuv+n+m18o3dMokU2YFsm
dAE5RGwSbs+PwxdFJYSi0cICA5qOaiBDIbigb9vyxxzm2A7WL90EadWNxxMAJ1+l
pFqSDArAKfq9HT+Bpd5/quXAt6d7W/W7frtzhGEYLql81dQLCcfsx/PIqtm6IaGk
k9RaSH9WwNPdmRF0M/eJ0LfWGGW7jcn0oOaT1C20+1tJZq0J5pdrFh9lNKKatiP5
DpKLiv5MLjsf9rQpzIdz8DhTpP9UFFEU1bGtZ6kNeluidnDAYjH8cgqlUIC3nv0f
oDMBTK+WvuD+402VyFcfr3hh6yUbhSwBgJmxO2Pn/7qXZZZIReMNvMRvUc0h863K
o1YlN1YYAX7/JpvmJD8NtlOVzRV1KLbMYfPqdE9V/1FMg+Z85DQnjjVZswKeF0Yn
KNpsqAy6O277ZfgHdlDuspPs/We+MMUmaZSHs48vbUdf2mAOMAK04Xmyq/mCHaYp
YDkXALPC2EC0UULp5Y+6gfZlw+LnrYFSB6tLdPAcReP+7HAO+Ru1l9onaoj84B5Y
CpjkVJ4szoXrwi+6pXZfIAYFf86uWTH9FH7W8HHj4mniK734FslaDIFZgoXCqaqh
KsfqEUvSyY282t9nRHwvtw/oE1qglYOx0M6no3ipxnDrQiGsghL8k4PNk2ERs12p
y8FcLi1d2LuFs0dj5wg94qFoOPscRZj62miI2/NB6g7OUhuS7dvDx97g3PltShV3
YuYHMob88fSMM9c9xHvIm7fu5rb2vkHciF+bkcOeBQ3GIJrJlph8iY9r3NyIF1M3
6eZb0ybzTUtwhsG9CiDfANnMaXbqEH9v7i7ntnFCT4mBPKtXPDxv4LFAt5DzLdY9
euZ1JrrEwv+dJ/B6z8zlbqqSWa+01pcdwg0eU4508+0BR27i4LBsSFtqIOHzXgx5
EulOj6Lz5CEAey4PdrE3xvuvyBAXYw1gb40lsIOcAC/4cFOJvI3jgPu0WjwgzgsL
vYwxTvR/K0HMH6kFSX3iiQYBfWR8ALR0G+P7SrfgtVQAsfsjj80uTIwJWZSsktWj
QFHmUZslk3PbXkdHrw7zrmkqd29gz3x/c10UivOt3wEqK+vwABy96he0H8G6Tber
gfXjXeCgMIhHno5LKtBnc/inxUcD+ifoNpWrQFFqfaOjoCc4FKWtN7tvnkVWo3Fm
iggW+JWXXTqi10SuYSiDxaW644YG49lzmocwIGeNSo/GIcU/nYdUin2Wof1PBoRt
GEa9SZq+r0wtJdeIw0KGdKGCFmY6jdSfGmM6QBcI2iVeRW55ZLOH1HHIaBUBjwBn
isjefccPmGw4NSuRAyv+SmTbYVjIDWYyhB2foMIT5dHSFvJVNHXSGihNzChQOKO/
Nh9UFeYd7iuvFgMMAaVQK+HHjUEx+TZytsZc1ZwI6DbJ7wQmltTTpKXbXwhdo96A
a0bDX/xWUeFOH2Rc3EQ7g1G3yW7uiStGMIR/uopGmpKP+e5JHNVJv8rgQe3xT2K9
so9HiNgCPQ45tFTI2zXlB1RdWf2EODUU5/67EE2Slyg9tW7Jz2QpOd8F2BSLGNBZ
evLkUHDC8iEonWnmilvfZNpm1kBV8wkSoz4olOszxlNC+0yRTyI+PfsfkPM3RlNH
cc15lgx1+m7jY9f3la00nX2KCSeo72gCWFpqyzfBMpe1C3D/7oeogO279HLWEKpz
E26I5xExuShU/ty2zfHdIRmB58K2tB8AciB57itv/jAUDZ26L2+ceoyDBzc11RD4
+sqO0tyFWyOR7JB+LB6yUnfoeiw/ckVkTB8J6vnocUbZQbQYjtqbtqRLglNs2qlc
k3eX2zeihAi0oGzWZxDoQItaZHykaxITkggYx/JNupg8ECD3M4g6MyQZbBmJyFeA
tQV/8MpLLP+Dcf+TI/g1l38tu0ipfe/kunqJqv/xDJcivpumt4zPuQSkKmXsEI9m
nQqQmtUt1NYcyJ296rSUDGq5JJDKogCPqHiOWPRKHiljLsY92PojJoAnl1GKMBLj
ppmmbVu1N8sLFaT4OsEUY4sw4rRFAwZQLZcq8+v0hgKAwhNIbqw+8VLfmhePaFx9
g19whxc/DdyqjXqz5H9D0FV0TEHz01ZmbCA9BRPCN31eIWiyRRC5tr1o6HQzvYpG
BvoN0wdgy15ovGsyJTAnSLgo9VvXXkN2SCAiRHCovr21oDns5ATj3rFp2EHyb3Z1
b4vZLHyIbp/Ib2PYlE3DNX8w2JUfMiqHXXOyTjwSv16reEsbrRK1KXJafKN7WEEZ
K+sUxX/sn6wxnIESucfKqft9hMa7BvajC+U8ke9vm8KLSF9iOnzrv9dttIK8z2Ne
EmE+gLcBubf26K6hrVcYk9LfhG4EnOSfa5CTcn7S/hWrn/f/cePQI9b7remXQIxv
xRbL/k8n/cXuyUw/T0Uh5cdOcY3leZCfJiol/zv5A50LYo7gLwEal4kCY4scKS7c
PELWQVuEJXTCRhMxKfQ5yX7IEibiJQAiFm/+2LlqCbo0ZzrUZQjKGNmVragFxWhA
oXFTWnS/l5i8xwkSkj3AN8RUAhCtaDquFi/PxG1wBXeqxlejFnaeJF0m0YHHzfOQ
Sbr4Ys3trx9pbKenqVvkTzj2EUQH2qXWxWHgsDKEbwdVRpl2QWzyeul8KpE69ZEB
WlXV2PK5IQnycLpytc1mXLRhPO5E3n0F77X+blfwq+kNkedlnQByrQde/ur+OW0Y
X+y+QWsto7E4B12w0vwVAHVSn6+Dn7g7tDBY16ST504gZnJ+Nhe9f1tAlP8KArMF
HfBuvqlPW5D6QD5dzrP+1slTwKPuXUETNZbLaHYdok2CfhBcgtWAthJGBIymnHTk
ZCWxw+/CE+btSNRvrRaSrLGMPUJPtDei+ymlKJQbwXNN+hm5whMgmrORVXv2Mhjo
q+YX7Gyyr/WQaNSQSVBaQbRcAsN20llfltMQOS8O9QqLpXcy2HHOUw96GcMDs04W
KZL1aephwJl7IN6Odf83RzgPVVyA8R825+/tayfaKomv7aJ1MYWMPlMedvPW0uh7
2sN6CiWHlnuS11HWqsr4yAdXRCvPh+e2WIhamal0e2s0I2QkNQqjQcklvSv5cneS
1N9b3Vv5wkUF3dicI3VFs9+AFEOJzFwTYFczHnQQiB5rTv/N5sWM1ZmdwOTxw0ZL
w74KyLBAwXJK6czv42gfBLEUROkHiD8TvmEfWtOLXUoCQ1t4Xy58n9XhYlEr83zR
kkDSqPrSwdQqvTJFU0OUcOGBswgUdyIhbMll8udYYWLcuYJcDRipbw6hlsH5KAjG
F4HdNyBOV6f33V1NNZdc0g/1w52oKS2RhErYu1EJPG9Zq0tymvEbdeH19DEHBHL5
k+y///xbIMo21DQTiYjWgR77VgflhQdXmjoiCqJPf1T8Cx6n4I5A55tSRpmyMwoL
zCd6q1sGw4Zam3O2r24H26BglmUHy6odeLmQbRLR5K8HVICG0cwc+HNhxNjQ+AX5
nw1Ei/1qUs2rBGnbjA5Fzxk1/kLySbbe6A4EPwp8uE3sHQw2yFZpZtVewk5EOkAW
yWF//3iJskdb6qb1jR5xwoPPfgXyH6yGhMUS/624hPlArwrnGVtoXghpDCONe2iK
kWAAR3Pf8ZxFDSoFdlwwEmXGVyVSCsjTa3O0PNqcHW49ACdQv+W62DN9uVLDvd3J
aaP0Rd16/UOOf805vBQCOdY+/H7GQ7Z7B4d1R7h1rMdiT6tg0Cb97h6nPBd0h61p
JZbFzFKiO2zcDlmo7CsBezQLImqsU0nNm87iqQYi+lxnEtkM1gx3vE0wDWu4KBdc
A4wnLrTSLXU2GJYRCIqX24kraVHjocJniC1MmLfzUFw4bT6ImhuBJUkVltticqdb
q44sPvIr2Ltl3xITZn8QB5FWvdVMrGamnXswovk2zv69RI97E/GNvm2WfS9unJIV
fd6Sbg6vf1t/r2UfcrmqL5DrQFl6h6GwNrVIhUfKVEJJ0WB17x0tkG7en1Vroi2f
aOPV3msGwfeg80cWz6mT+sOXAEFdo7fawEpgKG6C+069AqYDwmllDBdWXPzPyprL
moyqkEY/IIPO1BoUWUeWOSb9tPYofEmimSG1HQfkuJRaOa9zOvXyFFNHiNathSXd
0fTpNb7UQ4Se8La/mUzFVpOYhmSYcEFA23kDOCiE0ALR+JhBCnHBZLxuiEmeUXKx
ZUTzi7a5kq+tnPUxKGWdzAeN9yexivbPTPdNRPMyDavH10mTZgSuMnnN5ESzHKrE
ffbjeV4Azs+POz2dfNVROeeTjH8zCCQPsBMT6N1T36vJzrmgChA1WQ6rAQsFKQDy
QdWopk5Zu6f1gNjzFqynvS6i5kvXuFgD8ga/TVmwcz65kN/FWdyATluqX2gHwc/G
cQnfJhZCp5FWTsnPYSkKtKqi9d/PaqnQAu4+4DpGaIvTadzXq9V1L/kR/x5AmTOb
e7HRFMu39vk8UYv0tr0H4blIvEfCCP0WFmUOIQ9Fme7AI3kc1NeXCixJOCU9Cdvw
ezEf00b0kHPi5wWHZDBRxBtRx27d36Dtsz/oMJ/hm0MEMWKFlh7GjwP+AyERdMgj
0gyuN+C1F///JWttu4lt/KalR6Y+vLrgBc7PVxgBeewtVeZ1UddOi+kQaqqS99CW
Cn+dp3KbQ+C7qK8+dwMnfxhd6L7945b031Fb4Pvq74YI52SO9ah7lO8mQZWv8crO
5V9tXEdOR6gA9oQ9TJ8rgjWC/4RCZLebNZab8DtBPZldn2eNKUa8U7YjVYhiSe2f
uvetkGuAPVrzE2PSjH3VY3q95BU+43yF0znAM+wnia6nkjZ0bcAI79N4JRbqvMJn
gU5xoNlhTn+xREo7wgIsRtEHQ0voEsmOZ/dQBn8FGdLG9UNfBOanjh/eJ2Lh455N
+vh96afemK4bZ/SZc74QDXz1PFS28E3TKwJRkl2k96tPlzIqDVNbjd6LAeJwUaI1
k4JTYlQR3w4ygwrFgn5Fu2l1VWU5iC3rSANEN7xL+G5rmBcCHmwHaY58WAED6HM/
bS6ZPK49X0aXFtcoU2fas/egZRzzq4JoHcWk7FirE5M84Aze2UB2r//VRUh8Yrms
rfcx/dDmeIcTt/qbwYbMrfb4JFDer1CT1MJYf8OCiJ8MinFxDFvcenanIYR9Nr2v
kEQZb7lwMjXJRaCBnCO/Dt0bpvB1g+EyJrIGKIP0r+b5UDBPM0C1ZLRw8NWTYU9j
SnIqyn9Vd3+Cqdkjkgh31B9+rDBMuwzCrxknvCnq5krIhJ5gxd1KX/6wljf6vdep
PMqVe20HO+8PeJdJ5Ty26tQZGEiws1PKHGGzqcMAkuamDaPbHsikQVCMXm2dJZhh
ZGionURwEnBMndXwsjBY/2vkGm0XW3hp+gmiWMwpKiMwGSh1zaOfgcYbscAgUIxS
x8D7CXtoebLoHuZzQT5im9ocs/KKJHm6rcFDXozt8si01G9z4MLvyoypVhsJjE+Z
mMBpLbYkL/jpBt9Q0y0cwiZU/lpgQWr3iHMULCAuUCKMqwROrFrZyBjdqe0pozCk
1tCvWpM8gnUi0yH2Q3LH1RlebfezFXXCXr3Sa6q7BXz1qFbg4+zPWT0JJoPQAttj
L9WUhQQjKRnrdtFw69PLTF+BBmfCf0Hms+BTdrCPkkBEnu7MX6+sExaUpoV8/hcT
Ct1lJSFq+M8gPF/zn7wG6BubJJBDEHiqE4Z9DuwthTUhbuyePZobV08JGyW9/tVS
MAOEoJQUJvQRf0cF6JVowtqOrGHiLEfqVSfSwu0s11xkifxtiEDTxOHUZKKfVJDn
Hf+irqxU1onUIz3tW6lWSCEQx3ESi46di53XEotSxtswSPMX8AVRbBQk8xdFBSjK
UsKtWXRUjHSsa9/e9qDr1AEmksBxTmS3X5ns629RtS4DOpLOIXFIwWSN4zHvQIdU
flDmZ2HRrG3Pa1mH4NzByiX3LW2c7kHPd/GeE9u4IVnAUDYxSRIs/9t1AE474flc
60Dc2eg1TpFbhfnbdNOLNIO0TGGng2Z3B0TPF3L9+bw78Pq7vM6azLM+IvadInLq
lgUL/yHzfPiDKIqDNHrBMcj1UIP13danCHfwh6/pQUwpUq1SgWUrQioIbfnjW7+/
UjBbUSpnyCWmkcFvuuxVGwCFGUlp28jA5P+kkIklENAEeR1fuSwF2IkfHVCGHdv3
7PC8u4TO+4yOsJSNwIn2s45YC32CVELJE9Z4R+xlHNTH9Qzc4pKxvVkIyM8FatFs
A6VGOUam+ikl/1cLTK3dlXxoWea8JxbXuYPeE+IjzNdu9e6ss+M7yiLPYogXH/Ro
F7q1B9zg7U7v6GNw9AIQt6FOlv+PdwoV8Femh+tjAZnXzUiwbiW9Kd1BDM9WQptp
LZSzNEE5OxVchRfIruzi5nsAkPX9GUXLHZdWGEAecUobhuovferwPC5n2ON594ox
0MMUdSEHOJeWVaHuTR0t0PJOHfOlUNpzt4amB3Q7plQs6TRA8OVDW3OItNwjeeVO
mn4NbizeOTzNbmA4xnDapglC0NpGDkfpXx2jccRP1NSoUeboLKqlYIovVVybmJEQ
S5X+9pGD6L++Vvkxoo5d1WwLuMo0E+4HeJlqECKWKUcwESdh1JcMRtrX8x/QiPga
4QHmjuiO/+p4N5Nh8Hz5s6vY4Cbh4JAJlAlRXwe1mJELOyNDB9yHDLBATLu49xcS
KrpymJ2Mij9VIGm16Gz3F6uIc6ZwzESkrhIfoVyHG4f73fhasHnR1HYPmrRAcY0D
RBQIrutvrHgDSff3P3UEU3cUNZ0/MbvnTfGbvde1X3K29Hy7ZOFYnFRhbD9CTqH2
Qio2/tYZXwV2qIphDg6/10q3xTiFvwsfPkWfFyvTCkhZEZ4R+fBUyIZEQRudRyPj
XZ2XKyFUgWF+sNPniHw47mbSaMmOCY1ePCk3zvlq0/BtQYKFYf7eROjxP64i5UBl
RAXPB2MsC4tzQiZii8eu+HMbEedxYJ2NRQkr+Rz+5MTyHFa69fshOr8B54dAav3h
XSav7qc/IhnGEh+89jxd4DrRdNogypT7848JCXWbHnZLSQn62PP/IF1tE53t3cko
U6Mk6h9SLFpbOrOIj0VjsyemfL1SRmEhT2XNNmJsZtRU2Lqp3d6Zjf3B/VUKqhDK
yJelbuOKhy8UkPqk3zITA27OKHHiK8pT3ID6zlhenVDFIJTo5lYGxY8wHTod9q4S
LGtRAmj7JfZKuAO6JgHMvsGoINbX4cUrDe3ioQlysPWF3GKMmLs1LwBVWxJMbOf5
O4eodFI5dXhnLzYX2sgGawB70Gdqk3Ui6Oo2CpkWgCc7XwuyrOZC0LXyYsehgMHt
dNgJNui92oHPtvOYH7d3j+JOynyDE/a0GMrCa34EwcY9xB+vHlzr0gEEVoMAbEhj
VRH5VyW92OTd3ZJzKJWjVHsCndoixQObXlUnP1nsL7N0wDWpyd8+qKxfxEygCEFp
6qY/q1RVdhN+QXlBmzUDEWs3dEC7UB8xCrCCYmU18z6nEI8ImzApHhx2iJG1sQzv
MeSTP8JDdecZy+xOZsrsJMCt2zArDCIKWZFz+JeFht0RVYn5/01bPUAtblZmnxep
eqZH5Gpv2kPYFhi0pFvfXwXCRHuCerIeCIzpXhE/C748KKh8TRUiqQvAExo3cvyV
WUrbkkUBxhQ18U/WSVOeDQC0lIdTyuRX3c0yRAGpUHe2w1v9IJuaWrPerx6zwpdZ
/ivmjYB8IKAs4dARynqvTDZT+xVGOpYqlD8etSZ/KyO89cEjELGsM32NgB63DYc2
g4dQZiTFY4AMwBC2h/N58mMmaJSxc+uwdc6C3LoGrcOWvec6fzOhFmeBFUiU683Q
fqfcdlLkCAYYfhTEudny//QOiKMoYTuTuou2/QxNUAtvSb2vPs2YHNzKTIxSFOue
ecR85z1NDJtECO8sHu/KTAbpaQ5KPYTIZDgL2plsPI1PVrA1WQtVRO88osrV99Vf
HBVO6ZZ0GHH0+OL2l3msI5bB6pciFDL7A2aM48jwl2iXcEpfaeRaGUa02tKZR67w
MKpwtRGMpcTp7mOSSPbqjZW3ElcAtE+1HlKMridzUuO6UouVP3SmsTcqU6YOKe8a
cMO9mvTvZmw3TQ4VPm5HWaiFuz+fhl25mYeLamHVR8lwVILouN5AToEGMM+s35Jq
wO4+qzJjE0N9CX4Pb3zYQM/O+LFn2bC4TpwtqmkUSBtqofUwKM6+z1GA9Z7a2pl/
`protect END_PROTECTED
