`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2QeCbkDPCInzP3kfrBXyquLHYyYMkaNqsKfVUjUQ/ylVqpcT529JsnX71eMoUnh
zvYuvKGpr3XDetJ6KhfzQMYYVevsKtGnNQZ0UnYORbO3asDjV5ki4qHogrLiABfE
5pC6ddYEEe0RGzXYJKZp0Jj4b25h/iVcLiBh4lCLA0JvgTOIyOArCyKuF9LwNj8h
A04dylxbPjhbjNN79KwS5UFOnJgeedAxpzqq0rdILHTgk6HMf0x2OEbcF3lDU+mo
kPfUr5WMuQThmFUg0SdjolO6NWKTIBLlqtouhEgFaDlbHjz2a1IaKoHvHeqIb6/w
EyPc2BDZlj/l/ON0ihVEGUHUjHO51fAmmgPmJwp9k5bPBpLocijwR6XqCWjdez9o
JhYun+ZHhN2nyYb28njRzyE4bnHahg4/Kc5414kp/v8TC0r0JcmKz8NYGZZ/3S9k
ps0Fba8cISsQaltleXHGtcUrupdbWrZ6J+j2X5uWkrcKas+jt8Aq0xlWt+4dTS03
7Ugthc9gH1bIdNlPwTuRcPssR0nM16T3J8XQPL+zPt7hDBBNpwwqho8QGpdlzEk7
CPlnAeVnoFm2pMVnj2F0wLWRf8JPuHp5pAykKnLqrX1suU/cgoZ4lxn0nscEf0OL
uUdZRm1v9DXUVYvoMtSk3Ufpl5hkNCMogSiJjwIfNlfxqgmGWIEg/QFO6iRn2fxr
tjTObzjvS5Ma+cGf6Gy+piGRSH3KzkbhwR1HBAuiIWd3VrJYbCe1ZNXXRJGU0I9a
wDYX/OljbLQhmclusG9FeL+9rhTKzRIeqrsxCHPMKjNwcu2E+bUtNWJOM/F9gOvp
sot6/husDLpoXOqkbcCBxQ6h66JH3Fk2wyjStlPzFfFNsHc4nylMkx2NDVzuNAH8
8DWmB+Hx3CXmY/RgJkG2zOhmQ/CHwpprcs3YDhpVoPz0zcH8Bkv7xZHg+jwrF5yq
lmHPBTqpIPnSfwyjvphAB6clyJ4pMOLLSZVg64fABXlYLTPONXnbBTtHWaygVtGw
GUKOQL6coq6d3hfMM/TTTvWxRXvMjTmWRwU7j+fMNwr+ZcC2BiUro+WYKZAsVVa4
7LXwQ8Oq4NHH1lGkEpOtaqA5yqteAGWlbg/8eEHJ5aq4X1L5u9qevIGYVRE6+b3x
cYY01RkXWlwrDljNUsEQ17/RIRX56e8tILTYD13lr8I10WTYOuWbdT7xJ33e1eh/
6AKjJYTNfdRPMl6ZczJsxKzuSjqosBUoTJZ6yQw8MJZjojI6x/173R8NT7eqENZu
589BUZ2A7wCJ4fUFPhCnaxTXaA+aEBuQ1RiJQ0jdq0S/3RYyvw1ynjZ+xEJ8EajM
sJiX6qyBHcSt2Dc0Ogo8vJGMfM7snLzqzmUxUDp5zV91ksTZjZTbCjGXY3Xfqhk5
VEykEpo2Ck/7yYB+C1QhVOhhIT/NEguEnukdvcSDuHhEt5JYmawXsMT278MRQttB
iQm5X5hYDJ/oVIKdOzLatfpT+aoyvOYyNIDuDqDwifbNlljm4fJEqouMOGroT8F0
LW50KMp6C1rrWgvIB3tjw9Jv/yoXucgSU56cDJNmuGFezYDW2nXdFUOhLXCkrzgd
R4shDSpsGEfr05XeriHYBCpDVD4LG736nSnwkthgzig=
`protect END_PROTECTED
