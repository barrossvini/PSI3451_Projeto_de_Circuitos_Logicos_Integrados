`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bkTlniJBgfKZLrqYlTfm2rC2msqZpGelESf/fKc1VyycXB3oruOyiILYzY2v4LT7
I57cYW5cM0gu2btj6/JUcms/V/y4uGKCU53dUyoVphXOJPl1H8L9cDYLD19w8q1o
Op9Rb4brTir+NzdRc8+tu74aUKnHQ7yTClBXXYi9XP162l0HLKcUWz8EFwtCCuQR
fnjgm3ibNkI15hQBhxgus05tkchsJVMDEFtBeMIpwE1scBAFEHmm+K/su+jkcWoa
Ucxmv0wNcw7plx7Z8GyKxxbn1tK19j5hyKneiu/xpMQY14dG+0dChJSOewIQOCCk
3Eex6TRU6VscODjPIVQFHLUGUnLz52ieprCf9E3FakpzCji9DiNhGf1xvz1OGogH
QrZ14U7NKvkKTHHrYjogwlxC0R66bm483Sq4BHX9gu8Sr3MCKkPQQyWAFjiP0SVh
ZZjX3TTvsrXrnGzzDg6Zq1fAt8fX8AeB64gGfZXZZEz1n2JY7todHKLX7mjf/wv6
YF+9x+6S9tw8N+mSPeGQ6RfIFOxCH8KohZLI48zpC8QU/nqc/5aCmXQ1FP9EyQ85
qProWbJIDTEK/rivpIYleE8vriaNQdmq3tZ2iqeI/C+AllbjIyvDSsaSVaufHiWK
eF7tGegNKaXt+zduzD6QrbeBrvYpYtLecrNpweTxd4ofTACKlzN+KCRGLP329Cnk
0ybA6HihatvInF2vr22YNgnxJZnLA7xD9baGnKFKJXvux93pCplh1WxVRlRLfeAg
ue2tVLYqq+Bot6Yw60MsfyPY1AWT7JHHaNThnq86b3yN0mwg+Dkadr1QevF0pF3b
UIdXleSLCe5G7PC5zFqCKLjbQhKjhQafRndhEzwqDliZtwdRoM8j8erGBQKO6UG/
BOSjct7EqPYrPjfhn/mWjAnwLAhbJ/tNkYGtby0uHSh3l5nGeQVXDJrusvF2aTti
AAyqqGsI4Bdu3kFWD70bvVBW0dsoEYo6yHXzhPbvENJZ0GymDCo3bc3C9LAWt8G3
ZkXGfid9jYaA6inVy95UHNRTK4BfE3mUrarI30fnrFV8rPlEQ1nxmpDyzxHg/YsI
eXJgPDNlJqW5EjkcIkrbucuvafKcydiaefovJv3tuL/tk/3ouxZLgFiC8hhIJBNs
tzY5SZeP9LIt/rtvluxsRyw7YBUcr3rw5HJrJgfVfdYPvUHb4Q15ePBKXfqEdU86
JJ9qrWKKtz7Wl+VoRiBWuoEZmsG1j25F08rUYRsNsURPI7PWEVYjKKC9JgsxYl0q
dTRgpMG2T7U8x2ghW/IPl/A7fA8Ud5aaDgXH50fOzDDPaZn2zhYbfEq3wuI2zgl7
1RYdgdyNoJpwuFJBP5r8gSDQpqCWD8AkBYIPRSEwEklU72oCiLnaSiEgBzLscq8p
+94tdal1o1spXCAyBYA8X/bKg3oToR5lxA/GYZSioaVA/LkSONjg898O1+mGC4q7
tehWBNOwp+IKSponcpKygSu72Nq7ciK7kh2eG+RFn6k=
`protect END_PROTECTED
