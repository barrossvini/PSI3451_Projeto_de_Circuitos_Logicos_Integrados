`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7lET5mibvLWZTVIVEWbdYKg3pzLK6i1f9WlWFUHA4MswT6LBm8Li7/yiAFTccKLu
DXTB6bX2b9wXqbPHqwLjITjCbrgjOLkjkNv1frAJjCebqbDrMNbSk7csS6TPE27n
0ax2Htq0ju7PgpxkpHlkBcwX1IL/wb3hFuvV84j4Hgnm5xK+j378fWXJaFn7I+Ex
NvszNwyvnTTHV7njojB6NGXpKuQDFClzJ8g6hB/gUFRBRj4vnIQJ/Dxz5mNqN7xJ
b5BrJXnVRiGhtbBUT0Iar3Kpq+iViOmueJngX9Dn3Cvjq3DYQUTulXNHTG5WUKQX
euk83t0mceQtAwSttNJlccmG1cjLF7awKZk5TnwrDSh7bhENxWzlPHnpIZNoaYTh
uBmBuXdnjdVKTV9/rJ/Yblm7GwytTD5dMeZEgl8racBAH104N5e1wIpkQ3etWSRf
256e7mjt5qsRPugccmQch4WAFWIPReQEhRWy3YDF30UHtaElO242Y4vUp9GJwjbH
dQS3C2VvpSXZZvSmouN3vYIuFTKKpqx/FXrj7SHjT/KKLSwqSH6dD2j0MyCscOH7
wQbIfLSml/8vPRSqYefGjwSs/RpEC5VN99CpqSPUrzFsUwNn8+CVRohWrtgrnCQo
hXGsLP5sPeOTEq3a8/O6qmL8scBDWSJYwpHpEv0qWD9/sN1QLyOgkjVsoE/Kjmpy
qZQgMU/mewnmgXrBimM2/B+b2TC6rqnvjcaAQlDrYEMs3xwlNI/YBqK7NJu/Qccq
haHcQc9PC77b6gz18UTyHim5c6N4jotC9s4i3clBHMtZfFF+TJs2Ncxo9BlVB2ir
pwGF9+cWlSBhIkPIizVmCGXpDjHu5w/XnsI498MEP5CvLTzPBJEEB/biKHX1WBxR
NNhtse1df5KrNAWTt9QKxxqh3nTqMf5s3Lnd+rTit7szV17GT5EOe0rkTETH6RZn
u80wXBODMm5UngmSxJnpoY9FEWbY42ZAXeX1plwksKZhf6chfbDPwoCBN6TPfPBX
Nm1HXXWvxOLgLnG0qCTLD/+HT5MA5a5ixsalUtWoI0c3xVNdlwaYnTN/vxm11B67
K2sc7lQJ1o4Psk9XQrcDRsCWtQBdG8EUY2ATogmjKraxBr//nUE5C1wgykH4MZd1
rIlfi0h8LZYC3QNAhe7EU1Sc7uOXku0H+wON1YhuZ0ul9Kvv5y/nLoNqKbaDLKxW
pkVD1Xmm252JA+eTQavIWXckHRP8orIRDJUVWr7kxNFtZwC/ooTJDyEB8xiFhQ8C
dNHTtpbAxA/1rsuFQ4aDxrMK6WZ/+FMjSF0IKtm9GPgYqjdA6HjpuOAG7lU2blOj
B7w/jBVgHv5SaWPn4ZEPVnyBNdcI9qDVrqm+LKScioLENyqyDA5xXLD6tM4UhVxR
GUonNu2xUrRoCSOqivbgvVfOzO9Gd5EnhKJief6eeDRKeea8L6wPdOrawrxcDTaK
qTlfDAKn5PUSpVCbGc5zVxtaz67uzIVxMbap9M2lqlso+dya6DcM/YJRezRn626X
gkg4d6Pn5qLuenFKG7ChLtGfqWsHPthtpRbu0fWQ0PwXwrpmCgpXNVcThEiVC3w9
UlvJv9Lcn3gO4hl69KNPaKFN+yPJBREzBj1rpNrxs7IHe/qICNNYJp+6vqDfsRPr
ufVUGv3wWiTferXIE7GBmNwrcpwuwsZfWM+QjmL0vE7uKI7LUPBR6t6L8q991LwC
aWoR8WH5aEPrixjiSRVxfw4Kk7eLQJp1Gn4dUOP/cdlA1CbkFjny0mhSJHBIz2SD
wv3Hr5qzi1Txce5lP97qJKvyymscPT8BIT1sp1dZnmRDn5f2b7UQXbpXWhnIRzdt
CBa4gIb4Wpi16gHzP9ztso9Uc+xBEMisqsyFOCA7bZR5OGrwoQeAqOMtLPO3kIas
d6eU96qu2EnGWTXpG//awPI23a2NFo+BL3I+Io9M+rLiynWL4T8HszxQVGFFLZGw
QYFmC20vbbm+A3IiNMT4es6moYjOV8Rmq/Wp1vr2Zs0i/IpxCQz4Iob8yhLkDvOy
DApJrn+dMTPtE/Pw4sz5Rt0QZtuPKAXx9Z0P50UCsrhJlIDjbDNk9jb550mLG1o4
aCvLEn+xU4KAM4yS/z5PVw1DU9O88kdVhZTHUBjwh4ZsASgtDZ8nuWiyQM4Tq8zI
gaE9rJx1soZLsQfZan153BzHovqs1r0l8y+VznEBQnMRYiZWM8H1JsIT2dgVkR5t
nwU87C3a5aPWWlBL/OGiF2/5I2tvV7FDTEtQUqPdFKzaems1VmnYKL9dkS53rPO4
+bQng5k0u6tDHtwxd+jbfg==
`protect END_PROTECTED
