`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CL2oDFnylR80dxrbPpyA3bSv7t3PPqNI5LAp4DDuM5qhSbC1Dd/MNL3lAeCaJzjX
vIMjSSX+2Hor8/vPO7U5NGvRB6V9d4unL78/TYglVwmQNEOMmAlB9YRuccTwSFGt
QroUrxx3x57qYFCneb6ITPfSCuUVMDqh8e2cPk+DtFFTt3LRY4SWEV4Jdj8ybChs
vWcMG/bbE6AjjFpzood/fQCl/H8UrvG3Je8wCXZ6fYpQi1DYE81apBdX4plFWlIi
wNUCDjUxZ9Diia5C7Tqm1XlF9/Xd+Q8BViK1LxGZkfEihv12+nj24BoEmMQ5h058
i1wtG0zBXsl81D0xKAu7DP4eZoMuosRTL23OMfjhDsjoXnqkFPzcWBmWD3rYe2a6
l29k+yp8rCyIlh8lUT1sILgNLhbtFxnEQ29hLJT2lm1nGTCshVSUQMKR6uDaXzTk
XzZr3QeiEIK4M6YhB40kEf66kqYN8Uav4ve7xd9fGnXfoIp+NCBBP6xGCkmmzwGJ
3Y1vxDlglLBh9xl4EglZym/kuQmo9ujDZNdX+nlR9iGh1P1iD8zq/BeE2vVAx/wA
xykzzdT/K9Syqpb3mHhfXeQ0hAu4UgmHyzWYWWmvce1MzizolvM+QXVgi2DuNClm
GNCEHUAo8vA2w7IrDkLb5eT+ITkirkizFXcHDBkEMaDBfny6eyPrvAbJ6epoEdlw
rswUT/Qpmah9/9qsR+1pOpk0ZMVBIOMjI0YQW8kB0fd03uLKX6ze69RgwQ/fSKhB
uMSiT/pU4P7cuq/mpk3x3uL+C+C8O1QG+u/w/4tVhy9mXnePF8BKH6oujke1wjZK
m4/xzfNbAAkFNy2b1DcFWpqA3PkWTFTOY55mUux9TXC7saVYrfUed+HTfglLO45w
3Y8hfjEbD7sZK50/UYZ+iqpcKg7PTQEfQu1aOuTfhSbrOsOcb0zvyg5ecKibsOFt
b6dap1M7EYMWwWX7M7DdzB65wyNeY2umLYZx+617FCSMDgQyQRYQG6nS0PRbLTLv
Aw+JQfsh2oxSHREkYbmDZKWu/PARiuac06oiPGrI1o2a/QJ428BTAs3xreA/E7G/
kiLEMat//dzr1g6axsl2Z3nBr170zMEjbQ4TkiXIT1DirwtkJL3h7LEUH/8xfJAD
bFzYAx2/eoq278f6RGGl7wvmXJw+IyxpikaxHOiVhHUBSPhjMSN60fm0jeEnXSqc
+VuqJ3/5aT+wwNpEJdIXMK6BFJcfDky/RqfRSrw2GlvcD0DL7MkfpvkDtlUYo20W
pDC+8fSs2lcEhvFc82LqTwcj1xSJenZrcXnYh36Qw3guQImlk5hsWFYRHS989C23
QYXK7BSbia27e2IvVHG/63QlX443w5qkaGoWcw1be8Cyk+gApdqt9kacW/vvzwXm
wuFSeYKih7DjUVXB/ObypOlG5trt8sKK0QKKGp0JEJTaTvRj/0mcmfHoMo2YbBjo
iA92Vt0WI09gh65p6BegXRwWDPCZhQc6NIOW20eic0TPp6i+7kLQlqug12c+xz0i
H3PdCzmfKO8vb8XqYszdeXOWffpS1dtUj9AG9yL+gcB3x9xYY4oQTZen14ovsfkT
yD9HxwjMp/348iLxY6A+ZnsOpk3AzV1ZHQdcKIqn0c67XtO9cCEtX6sVkmgrHIvR
U7tjWDCfLXMXwdqTlIEa870JOC4xLvz3HAeoUzSPCnHPEGX5kWJGRo5qvnx7tx0b
KV34+/OJ4IjfapZQrG7CfxAWl5q60v93o176QHumUrJPjudRRCsszd0Vo211zLdO
yauOPtFFfJk4MrHuoi0ES1vnzwu2YqsAiVOsbX91ED3TOUPU1/P0QrNcZXsT9Hw1
pX0OAlJMR8BHWXFEe7erZkuTW16uFzu9H3XDDIpMjRJIePQ9hnThrCUUdbdAybWR
TU9VbLC86L2oLa7VgiJJOl9bbrXCzoDXs7AI63z97Pz+Xbd1Hw2ED54mSPHQPY3D
cwk3nJPwzhwF+U/c5TVCHBkDd8i8vaSS1m3oZC3QrYGRC+j96vtLzQNvsOVmAB5f
ynczyqpVjiS2AQUpI8ucUWOFj47+hB/igXTpPbonwrwOfAqiWFTp16Pb5lvDPGoG
CmjLLRJIYlmf4Crs28bd0Cnpqu030H8hqe7PLfqwbso1TlMPf07z1z9gf/h5oxSH
OIUDloEVP3BMYZbHdlNd0xEQDN+oooofgkuSOTtXcK3T2NK75FSWEYMVoM4N2KF4
9IuFVs5OlZg3cbBs+FyB1dqOZ3YaKRmyYRQHM1Qa8mVWuTBKM1pIscFy7UzucET3
qUJoYXEAr6wAWwyR88uDCHs5Vg/UWky6UgS9YoAbJRdD/jHIgFvoATuB9gueW0CV
NSOmfkakjeXu76bL0JBH623Ag62VtAmy89hUdfEdVq/wbQ+miKKf4rRQQghk9Wz5
xkfgSc22MFpa1mpPJ0phEiHE5w7bxdyRPVHCFSKl+oYoOguodUzGutmhFsDJnccc
VdjmxXlzeDlhgXi3IrC9K1PAuDlJKkzJM+LwEOkqta/9aAwmEm3rIFh54/GxUPhk
A2y9EAslShNoy0PkT2kEmKOEG+gG49qHZ2EZOim+BXGuo59SzcghQfgm2tKcna4E
15YTODWfEfchSLXoHR10hJwTTz+FKJZu+DVgvrnotyWVLWLXxPmjhv9yCCMF15q/
51xwmB32HDu7nhKFsaOb5N/kjIeBycxw8V+8pI4rLXvF2TfCl573AwRN8FhzbI1g
/H4mIWZ8Z/YiX3FljE1Tm8RSfoAd6xKG4TAjNTQ3qIFN+IsLEnYHficP0r7v4sMk
QMmTmu1W3003ArkeIWV+C3s7TQEef3IjZwmle97qsKPGpzQKKBU8dU89ZJasMo05
KNDzISMaK+kWf0xhSQ+BU62hZi6CbE3MzZyeypr3uOzeoGcK7SnMwLhOj4OPaAEH
uF9DPA4Dx4RSO61P9pZHBl62LuzYGSbGjavyxcmYVpCT8hiHeSUggc9Tx+tA7o+Z
VrhDnr4L0x5uk9quOSeTpff0Uje525sthbEgHDKoUSskLdySQgdNakInEm/rRpFJ
1NccREHMXCMx7dxKKly3EjjrAHy0fTOxgzGl3SvIkfQ5yIpATsZbcfIA2KTrxETl
FElILs2V9XEOpOtIaUFj4MpBhSQlEyWxTz/bHsQUMjQB+RmXBbKRLBjp+LW3CA0T
H236wUIXU/WccX4Lr/KpqIquORtDW680t6YIpeCNtf+aQIFp6qNnoQAEFXOB4ke6
DhCyxaU9/p3mojy4O0yb0YzaZCdNQwZjnelCjj6HJ29k5yLS1u8HYuF2gTeWxoTG
7tLlzKBYrFiMpjqCmbK092PD21tCeAqkdwe+Xf1AtRwrcRIDvQz3bBWYdyvEbYBO
1w7PmMd2jkMH1guV8qlrmBUdtWjILGg9xFrM0o0oy9Eju2MLbKADo0D/dp38zGzU
i/rH2GWYpoxn1f4zsnuuNnfkqz76jutTAGD6YOsNR3Jc0Egs5RWFuo4ic4dN2FUk
UTbNiaD0C4dA904rG0n4eYLCLdFTKkDVKei9g8GoandkGSrTYWX5q9GBr9Midb99
WL4vacIgakmaTUdxXeGCqLpXNa01exC/Tvfcz/IYSuBk4blZYEp8Qa/tz3cSDaMq
nBobqHaksTKznFXeiFWv+wGjxsshggMwGIJGNJKXD7ewC4/2Sx+AAztdGlmc2QAK
pM1ZD55xYAYZqgmNGkM7OciZc9ycY0CgpRLiOiZv1ZkTFvj+kgbdvhQwAz6HFEYV
HaNjkgf3dvoxOCTfFCxPm/E1uFYiu8sL5usLkIsZhPT35Qpuf5cwdnno6Uvlpx8I
mGOzICw8Rirjx6ZXI+8o9bpGVmKll87xEssgAxTYBHhIePcOoHDYvbJhHmHA5I1F
JNZoJ3vBCkPM2+bqlXBoFLJhyThHu80xe8UEVqG9EUNmQOl6oPgt3vV0Gbh5jv76
b1sed2Qd1lKmQxv3cS/+Py68FaR9cf4ahqvMrr28gaNjsL5mTybuU1j7qpD5q+eY
DGpds+v1RGKdEBsknGoFvPT0mXWYQ9OiJZzPq9m46/vdq9vmnbAKt62Ky1JmNb0W
5sv6XQkwflD/DjRs4GmpC+vMeKRqk1vnsxUQNxO18vE8b93fDQA7RoZQdQRhheQN
gEjI3DH9TWuszCcJDsoiOjPD8jsdmSesjWDjUhS1dvWdFBnCo+x8wnoL+cI6ZBLY
s5GApZF5HcfUZ7MamrmGpfCZ6N7j2NncCkD5+GbTFlD69cN9DEG2EimwkjWqNOA8
d9HSL0IY0/Iji6kQsmCtC662b/sNpIRXe/zJe48uYX8ObqpaBNTTn4fIZjHgwyyo
03jLskR83Gr/USTqXTdRKd0ACPeASAd953mr0E4X+aJZSaQdmM1L4O1uglcQbY5V
0jEJ/Ep9FOQqKHdnW/lSn2EL+PdaJrBm8t2kwa31gOh/4tN96RJx0ce2tpO9HfnG
WryPZykGjIDPp5Jkhf4XlyPucaM/JfdFxRvfn+fymA+PEgIjvyP3GcFEafYwBihW
1Yj3yuKeGjpHn3rJH2k1AL8IxSFP3yVIO98bS0fO4FVe0YnAPDhiC0xpXM6tcMrP
uvTb0L/VcgF8qI05OCOWIFGDXPTZY6XTohojMPM1YYQT6de5TQuJpunlBLKyMLT7
mRZF/x44ijIvt1rxhGgsJRZXgiSegl+sVtezBips9YlURYWIoewQ2UqVKmdkCBPY
aj3ubOPC6hpxBQBzxUoCZLWMf2oqQ4nbHoTpxPCu90Zf5+PBDzVwy09hImFzKFow
Nh3sUBo5R/MyUBLFHoT6oAB8SwtAY738HnqOksU9hExlNabtIRRLG4qeZYsFHm9B
MRYwbIbFVkYoEQ0nbHxWidpCjzEQWY2OwoxnA8PwIGciNIZMrXqYbJ1/Fme+W5ql
/5j9ODIH6obBQ9tF7QDo5v6NALkOskVvizwoYBxy40R03P7x1N44OWaLv15sHR/0
ernNgUYIuB50xE5YEvhV9iXWMnV5vqXXG9GLjW10eCwPvrFoKAjggEHQSrrID2JU
KBFVd07Wkc17znk/0DGX06YHLQGbBXcZj8+c8oBx2N0dDBInYOpJOfk7r9NJn7iU
tbA/vtPxufEC4021pozwUN5CLSmvynEaGcQKNQLxi5hvlUahQRvKF3WiBt+Gyzom
bpNuWWi789gI9rz6ig4AsiQWnBWtAS+prtfqKB+AlYHXddOSBvQhG4KB6vXQgjCO
EhU0Mv1jeQ6zvDWZJg7RwG6mDzDKIfitRgE1jnMO06PGlnjtBmK0UfbeWwQGzk3D
fKGiPNqSrSZogX0QhkwJ61BFwPlACDTNKdXQgOOsIlrZNccHZu9UMN7Py3apNGnM
NEVaA/qLLksD/Owyvl9bWavQ4wQ4ePIJ2VhNxxnEvqlX2+PI8bTRLfjR/SC3l8qv
1zQvzz7yyvh8AWOWUhqME0VktvAKoGwFf7OL5wlpqg265Yc2zNmCz560ZbMQ1PkS
SLa5onp4LEQUpIcyKzrNuO1TYcpsW2kwLmtT88wrV7YkfZsx6pFYXy5MrlUDdGVl
A0CNftIa4GVfxXfG6zVz4VQgcW2gL47LEbx/MWJNyjBPfonnAAPSQzQuBUu/2qFO
bszbYLWG4CtmzuSUZC+0ySRKc8gzXCYrT4kEqvUtBtjaNy1+WHLLzkZPOARHhA7K
2LYCrwiZE61Z0ozku1qozLSb+oXrJiIP0hrveuZv7336NakniEC4zKBGH+wXBmxA
AoZfwudyDyaumSHqEhyMNlzsrfAqOEjE35mF6Qx8B7SWoqzfD3aK2Jyr5xY8EeIq
Hkiz1KV4ubgE+sJRS12LTne0au2CxxVn5iwjJQNsCzmofzvceep2HtSv9AtRou8/
PxQFZsvtd4yIa0HecNHgMUshs8anLDKN8oNu0jKCOTqWSsFy4SWtxnOIcwXJJ6m/
xbhNaCbbSxE3mWIlZBy1LsdjAFSXveu/jvRh0QRUqiKjcpU2pl2FyP4TIdfJ3One
DkOTfMWykpbPMnWFZeORA0jg6xcXnUO8+j9p2USzZs0kQxBCViYpe8OiH8hbS8Ao
rc15IgEPE/lZ/MkAT4VLHWWyxL/UTTdYnvxMudfcwgZ15YjEuvvTdzZvM14GCKdf
Hdc7/uMtWh5Z4hTff878WiqxrGpSdnpFXsNFZ9vJtXZFfJKSKl/vqfK1T1Zc82mb
1F//cHwjgHHvJsvp+cDAsZQgD7GtotRIMCzFctEMKowmdtIXxolboxz3PCeIjEki
HCTKQ0zQZzvBKH5UNOo7ZpWIriEdBNOYXg8CD6oNSydj0A6gFxxfkRKb7L+UXdSU
i9sQqmisqKX8nclMIVNymiZskMhYaHHhO7bQkTgxwwEtvJLMyAlQL/rOC7LqEkKR
w2q3lrf2uDLd7XEQ7G5cV1uhJV5JxaEXjkRuT7V/9rVZSdWOb9bbwAZWUtd8uZV4
CBaGf1PUHcyOG5sGgpLMgChGSs3Q6h06n/tYOaOP9eBXXp4Usaukn0oZvU/Of8MA
hwfL00XMx/oe+TxFPTbgiUDu+82RVAIYP2kleH5cpeqnzwswi24lfNmVP7LLHIbL
9Q8wQuEz5y+229EsuSHX4a18BQ9guXISM6gooUmAS3Qm448jma1BXvG7pGr9YCxY
ZhrpgpWMP1q9YRm1GDYUqOs409rBIgL/SLsP8f389TgUG83uf1j6XUIN8gfECV1o
dVEUcDbi7YOSw7O5FAxv+rlnY/4eZRUCXnOHvsLkjj7qiXLmjSqOvUYGIhNAgy0p
o8xPxKraLNedQD7hpzQCX1PYdeFyfA6YmoqQ4FaB26eM1hbIxVW1e0Ch/cKDac0d
m2lGtlFz5eQbMsqvAn2/NKDE5/YNCVqJuzHu7zmpcaGWZKIzKPdOt77AE9bybJKv
EC46Go2kvW4fIrtIeCUXKBqa/gKXuqjcgADhqImyY+wedD39IZRmE67CoC8GSM27
Dy8l+2WoFuqHKq9HjDCze3qU185j2jjsWBwpJtZwPZI0ggDbjrUZVdM2DZjL3VW1
ZFRIY+N/32EYkTGvLDLa7Bkff6pzalWnYXjaIqp/p90IK8X7+TRdvW/TrKtzvz4c
Dz8zL3g1qsWJ+N7fVaIz0YYkptRR6478QzXBvmyd0aKQeRUGlyFAq8zpnlE213Xd
4MCz+gmOyoX7bRKCePkxJ+469AR7NdG8btnxs5pEJxF6YI8kV3sNv4iqGXSJJ9Jq
Kj3xrP8xtBs9qqPPScvCHGnHbZbi8bc5YeD26tA1UgBpISQsz2vmiqM8H1k40Z95
0FRbKl356iXIQH0UgRX+oWYFoN7S1RCZBlpLXqsEYDfL0jTM55sff7M70WjnHXhr
z2KnLwac0ieVgsqyEstaftxmy5NEeR7jKihVB7B51lRYiOsYSSnCkwUh4pIJ3dCj
1V1Bw4pz3KVdcbH/9s7DaTRmv53H5aI+vi7fBMqEY5U61oKe4xyAere3XIjE/DPU
J4B6gb40wnZqNByNYnb096VC6Jov1L4CKCDmiloDk++C+0186JO+04qTe+/Puap9
B/W7e4mxamr/921jVf7mlU+chXvhbB9qlca5Tx2v2Da0vMA37nJ8WvadIAxQDGp0
T0BFzfnwy26R/SYZSzmXyfW5haEOwjSwvcUYgXqgqJWSfnm/8JHLKe0376y/J7nC
1bUUXckbdGHvK08EzAWr5nBPLOTFTkv/VYh1Wf3x4vmx+MuU22irHPVlAobiuNHo
4CBoxlWpL9/yP7BhsjTQJFXF/j9QUtAU/0vHF/89/EnIBs4mCTF2Gu42OhbfxTa3
hGaqLAt1BpcjLWwSsQz8ptr1zaOBD5Jq+hAun3SE5YHDrkS4SePPOQiJtwar46RI
z9D5P/4LJ1HIPRjYHYJBVRvr5H6L+pBil5TAE8sCN36X33IpnLyBR2JyDI7vAJVA
jJGwmADA6xfCXMNb8WB0T3h/TeYva9gzuw1abKOZ8/6+D4ddnC6bsdsgNlftn88M
ziXIBbbnE8izkmB+CgKVvkkcoEc7FUZNHy7TKEJSGTRAAEhAArrHA/ZWkCUaChuU
WzmS/yX7Ftz40UJUkqSJ+zuq4Xh941YEWSl7Q5kW8b7dL3P2wdbsl3RCC7D4u1hI
Ts9q3wG4PpPc14JJ4+N/3TDIYimZmfKW6M5DUWysOzZhuZ18kIwMu2ZUr6551tSe
epRcTCv9C5xd8flEM14JWopXVusuOZJYzGiXJSOq7aXK/s34qj6tmHTFyw04fnKP
vN+FAhS38Q679Q+FZjxCrxgJuNsZKFi36GpGV/A4of+kDY0krSpCIFigerj3fRlf
wuw1h5d8s8gRiwhHKfgQ7SvqIFxg4lxRA8Jcr68UyoYjlLf+kkBPZyQdgV3Ydy3j
LKFQi3dMRUHU2Y1lsHg9aOZS7gn265vrztbnUKkAzi91SyBxWY2tdIyV1ntqd+TU
9Eg5Ei9fKdxCW2sBf6m3pRQMd0lv3eF98f/nKNOMpGlSQLhwfSMee0uQDQBbGm46
31fThu835NjPqr84deTflUVCa4ABDS7cVpwqJ4J7oJ8st1cJshTWSKCuahtTSFU5
lA0iUzauGWyLh1Gaw5PvyPywnONhO7o7YZ/TeKz5TIeA/VXxCyjQAF0GzKTi3bKQ
cwCr2WKiEro9oRaR6Q5tL3hYRwafz4NBLfjEYxBrJOMZ4sxpPZaIRn17ZkolQm4a
YfnaK8mkZcI+3RHL2aiTFSQmFOlnkNiGn72Vimk/zppdt45zeR7Akr4dqJtw+Dfl
QF9LHQ9X9NqIUMdfKvlB9tVOW/uV3Kx0YrCP3bEoZS60srFA1v6gtyWoIulgmfQq
PHsrj3aVYx+yvWpTKjtJZfXzfc1U4gTYONfW6qzVprHgzrReXKtGq5kzh3YR+gWm
WrqLgUCsHVoPiURIQgTBPA4Y880Bdp2usXKhd7AT0TstP2bzPaB5vf4LeO2qOzR+
HTrPIxpA08RQER8UBUx24teQHSZ0/iEekqzIqBFNW2g7SMrq/fZSjDu87t3Jg35V
KrS2dfNco8QhHaDCdLnK5GuRKOfYmx3lJJhppqQajr8+5/0kKu5pNnkb9dAMisYe
Ek4V0AZypxkz+P3/35o8PKmL6qe8cNeeTNLPLIRIJbeAFZ1lVaz3E6okqG9UUhCk
RktFTWZ9X/HHREmYvsgxWR86B7KdIBLcQtjPyWerS8k97yWwx5wc1hzJ1CTewdg/
AnLSs1b9eYFA2W1gQE6sYBDizt1/R84OX3HU5C7cITSNj6TEY1ARvS0Wejc8KR5E
YM8E2d0hIYcxVaowGZbbnIQ12fjnFtLZHlzOkIoDZjJCOGH4L5Y0dmMvWdp7OSMP
AUAF6KDX9FuaVl7pj9zT3FwNJ5KpLQKx0fOVufGbPp3pmBlrKOlW+LtrNj5gORuz
mLszo5goD+guShnlODD2MKoTj7yUwyd4aBosKO5jVUtUngLqfJYHWjBKHWEN5VYV
u3eQhOF0vXJRlI+0EJOdU6XMmoIND9Cu5HmuRs+ap/32ejaY0Zx3FW8j3tOi+mmC
TcW9MLUwn/lvoOl0diD7Rr/BzmXHgP/Ugp52CkR7Kiy6wPMSrZNplMOVl0Ab/GaD
b6cTp3Z+b36pJ5LKdJUhxlgaHSHxGLx++yhcCdN5BhA2rjHTructa5yJ22481uw+
eEJujs4WhZonXO7pcfiHBzZ5wxFV1bCy/1Ck22iT4JGiADecN5oQNeRITw7KBNcN
8LyGo7izmGZekCqXFHqSm+SVuOaQQhiJGEy19iSUQb9f4A1wTckG5uw4nX9TKb7n
2JO45YUr+2/bwLg4daujEONBudTqjHPFbmHsnLRb67mtDI3ONdlMW9ueq/Gi0eRP
fzUYtPR9C1wVa3/+F6gKR/LqvyicbnIMajFcveZSfJoNvtUKsqKs19UgRTW+6qYM
qJyIwvmp8btQ3pDd9zjwnlAQ0630aveE7ewbKEdszu+tGliUBlgJtmW1OcgYjxe9
i4L4WpaIoH/apI0RdteA58AY0hCib7/rbKRsj2KJT1Z5hx4Rt/Wt0jiPZ4V5zpTM
x6S2xiZPIQnzUn02HAZHXgHRYN+5svEGaThmE5u2SFhfARSM4JhraKGingjbuAMz
jLnIR8j7QaG9l2IWQE3wZIRo2ux//Ei4mMlOp1eYx9/HuQG6pRDc7X0AFQjHsma3
piFhC6dhVShLbHzBrBd++IHYPLuat98IUuf64R72WkAfqX2y7aGGFsqFepjerVgw
euAMEafijTvw8lDK6T0hGZqbd9OQqoLz/qmzkIHQr4gezl4YThy2GAFsK6PT9FfF
z1uLKAKOPl0CsdQ1C2v5QxmmYcYlM/1Idb/IWodSJLN0tyFs4WlatSyedRk1blpz
dOoR+V3nXGjakpZESrFTFRwXWs7duaC+b6kXCIIHOwyQD/oqHUyR/hCe93OYKcdl
CLAi5Z9IHbpx629vdbYzrvCOXYUBEAeTTggcFFuEObuHh85tRHTHZ5l/0yEQq9kw
bLvHVyklFbjE7Xkh2dD2c7CtoOefLg/LVyBL3NFLsznN7+IgwV7vrVyo1MG6IwKU
8c3/ajmap0nryh/Cl4+eU2wrt9RERJH8lMSSO9Ar8GusF9iqxy2uEPCLkqogkxYa
7pVUWBwIpXTEm7MMdcVJgXvfLczuZwm5gMT5Z2uz58jOxhb+/ys+xuQtblthB83Z
UEAqCkcjiUFM4LdMYzZdo75gS2q/M0hTKBmpYmpRdPdqhMFbhL3fHClVwpERdEHY
9EKZCM0QwJnmeGHIJhhcUKyNV+RhbQKfOqysCEypMuaUgdzahmY9DMqkmUcTvKY3
Hmep9xgvODSKUi0N/HIxifv0qzXgI/UGi1BCG6am5jCo4gfmyIMLAthedmGMWx7M
ZdmlDrgDzGjnvtqguo/Vfz8y6OAdAouk/EFC06d6qRnJUfsja+kxB7AOxlVaBzO9
Zwu6ZqY7HQEmRiY/fubp6eQZXZSuB3Az2504e8t2KP0l7l2pomMgewuSFORreeYM
COehNoHY7oTwf8JxWXBTq0lQ5YKjoPBuba8NRiMessIq76puOfaF8dVBL/WLqFMg
4BJyitTLBgU+z3QUzTmKI2nkslfEljGxHlZFhSurPtFb50rEXALhTRdkca1tnBO/
E9JoTn8Yfvpke2Sd0sqUMayOsDsWgU2e6KX31m/01L0+d6kNq7z6G2vIgsDJ9f+O
LQ8zShwI5MhIFXw+OvOhqW1t1fn9nR9i0V0uKyAlTY5EEuBT/6AElSjxYQwxLA5Z
l6SL8FYqjsqrvAgffT1ir5m2AqG+59jnJ08RG9kKfG9iNt9ecHfPgMV9M2ZLvK0N
vAOwOE2aQ7kGaqpX/VYqSSyVbfZT9wgTXoBIjUxD9zB+I+5y5fl+9Sn8uqPNLEkL
Je0L/GdG7Oiw8NhGPDeQDO9e59eFhGwNR/Ry6khL5rz9MvptAqVAB8Yy6yyVLRMa
bKCMu6NC6SSh1Bvc0oUm0kOACk0K0LtnZS0vv6N89iL28q3pTx9pGmNx7X4Gf+mv
TzMZLQqQq+FA/+DotBvI+zjLXWLkj/XWaRQ7WUsE6IXzwkmLCUrFQt+yhFN6dNiX
mIAHdA39QtryzX1ZRyZfYTeJk0lHzSy1l8H4EKyFIYny5WgxyWl4UePN2UmscGeY
7uxojstI2t3Hyoj8nQxs+1OtTfv1djmUvuGXSNd7fF6O0aaOc9yHc1/Zfq1pPE+z
LArPd+xoc1GlSUo5COo2Wg3J1nWtEbghRcZ2O6tLhw8oHJ8Hvqb78M4Kez96+kZ9
j/GloasaviVgH+aymEYyvBpi5Vl/imImkyUzLk1Grr0r60VL4nfFqSnCdde/M1Ko
bsMV4UQ0dGwpAH+v8uuEvvASzW9B3q2zrNaHVIEGJLIygTMqPJ7lx2M29ytP70m7
L/qq9Cd4MjpKYozJpqzzRulVXQiSNB3TotiHXJ6sFAnUCl8kV3qvOu+VPmC+C2lg
k6HyyFv4f5br2ut0jVwI48imdhrvopWYbkeuo7qUZ1Jd/39i0X6VLc3NabqoIi1C
/wd33nLjLkjBGGNnx9vNhOI+NTm4kLZaeO9U9TUbsYlNTDZE+Bq9vOjHBqKL2Bq+
FJMPj7zEr7UjRcLqVSfM2KV2kTg4ELUppDamONjV/TMSXuIjy1dEw5rgMpmZP3fn
RDzBjDgM0kqd66lmXwxYZnvd8k3OwmZPNFofmMBU+h2wSP+Pc6BEvnIu6Tg/I91N
qEcozViB1gGX0t7hC/6aTsDu4I5Z8C24ulFekumLM3q/UBzIBdWOkO02OCxY9eEI
4NfbMlBII/eOgMfgmp+cktRFC9rj9i4ZC9h3sw6FvD36wk3xyKQKcwmYqT6gKsOz
RWrzlqcGqicgKAG9ZsrVLax21j+QMs2T6y6cuux/w3JybpXb7AZdfcprj9bwX9ag
3s4G7S7T1TU7F5cUsBolrbNbW0ra3uWctKLBOPjOn//j/Q+VKZhfRDmUxBLsuqrv
zkb+CbedDDK5ZrsOdy2WdlsXFLogd9hamgc8igoIzhVlfjTRkOWM42hkzPACABKs
Sy8PQkWlFZKU4ffXE2olbgccYqAV3vBzDq/fYZ7anaje6xBXkUgz4Y447gMnmlIy
s3Tvqo29uk7QWQ2EpA0YSHx4zXX1SutFsmAFOefZV3ZUP+LonTqFWEDzUUrI+1Sj
c9NPUDjnbUdiJLxTf51pUKDZt9vTGApAhOX3O5hYl8O9MYemPlobaD1EmlUU0hOc
ReqjxpZrPeOFduxsPmQDcX/Jv158vkOLFVebqCSHtTkw4eMCZrVazf5zEe5XfwIq
NHneljaBNNLNFoGja4Ej1JgFsBMG1ZZ4m/3eYk4v9d01nBYPxvHjKMeMS6wPU4ex
Ych2Fk3XPHgLm6N3tlTl2GWQbkRfhYj3uWSOd6RS3onWr+8e7DkSsHQ5M007LOJF
3pVj/uI1+aky6ajODrqp10Tv80zskBuLKA2MqJrW2KGQQheXV251iBuf7cN9FvTg
c/34iD5gIJ6rGdAAVu9fvrRrIkdbi8mjZduUHtim3pqd63KcOUT7D9kkOPT+oIHr
ChTvY04NO24i3YDBFPXoUxu27YrblNY6o3w13mLolZQ4FgGRYN4E3BDHI21mEw2n
8deE9K7TCI9Dt4xU+N1bOzEsgOOCnT94SDARKskpHjokwrmA1AOfRiP70kpMUcEn
HCTFcwJbM7ABpOLx6vx4j6p3cDwUC66+FdlTKpOB/XKq4SOFaBlRMnh9GoBPPivG
wamMH1QFNKV4j1/USXtObCWoHdsxTcj81cV47SMnTFXcjCfICm6ZZAjIGy6pDhgL
mwcy87APmb4UscnIL3weRzvk0Icl0qSXJRCaJotKYsmREvsPvZbyRLfT1FeQ7dXH
/XgrCwSb2+LRyqROpGUEoICd+PHQ8a865Rvfjy4c57ljhLYabx53YDLXFFt4L2wp
3q1ooyHZUNatbbYlOKx0dXg1wIlWYNxsf6PSJMGlPD5EwFDZ7975If3b2KBIFWR0
SsI8GX/dBAm1mG1QVdR4X7N4PCXkrHniyHYsYdv6/pqDLmsdc0z929dwppGAFNAr
WpJS4RsYZwffklWF24bBH8rmMuyp22vK4//WHW9b+jJqyXiMD11oA3ST/tjyQMm0
qFrpnu0g6j2e1o2ieBzQuRmUwZKuA6M7lRo74/TB3rGZOoVSVnkG8Ae78CqTrstU
6lUEwLF6oJGzKFbm35ainDvKFLhhe5inrnfMsKPi9aRK3tYKLV5K6PiI0jpCj+zV
7tkSPjUo8kLzqBw98kwKRmkSJ9VLPjGipLL1Q2D9TmL3Yjg7eB96AZC600iFZtar
P0FiyNAkfqVdrjAGDNYX7WTTJ43Tet8p7nfBSYFP9b4G4CNNSpcz0QbUaNQpGrOG
C8earrc424ZBzxJDyOZzcQ1iy4ev0QM3W1GtXuP5u91Kg+AcPo2198xjfZ8CrXT8
fN4pHjF9iaIENwBpY33OBstY8kZnvsxqWVlh96CD7BLYQy0/teeF5zHJSYL4iLS4
N49dvYL9517ZM6chKYvRs1dP2nYCvPhlPGQSpL5dP42klkTW2HLlFta4ffVImqOh
1udHhW1ug3R55X56Lmbm4SulyjcU/z6vvjoNinYjzauwSvYIwcLhB+Ct9/C3dmDS
3uqrfhFTSnHGgoYeQ5R3ivQl9fsNIQYIFpWEb4Z3MedU5w/QK50DNZoKmR+JATRo
PophOOnDyJy8EBVpnDUmcwAEQhOo72H0XqWPPJbnLFJu+6OKRVNv1DzXdlStqGvr
c2h6lOqJmuiCwXuOsB20n/QfsjU3XuZ+FtiXs9DirjV3x3fBOZrkC5WYO60WVnTw
LvuYohTmvB27r2Q+lyHhJPbp+dr6hrpkGYWz+9OMR2ESx25jbGnFDNxQUA/HluiU
YNXHyiCoNzc/9WG3X05+xQRkhEJ7AR8Lt7MYuUNR3R7mrZ2t89DAIYBptqC05H3G
DTgcgcShQfieYH5iNq3tUdcitAS6rRlQwbtsGCS4/Sx08+QbZRU6LfkSqg9vhv1w
OD+lcw4QxwEG3QOra+yDKdORkfrw6Mud9O4J4nI/862N3TBNGakQeRZEZHP0ig3J
IfpjkHRro4pwM0ENwLM2VlkDb5vzpTCu2GvDqzgfQNHjqvGXBMfbFXE2YbKyUHVO
cxgBHN/Fr4KOwZ3vvX/2AY9W/9TRUczyHEgPpb7kJtUq/xOuZb6SZwy8V/zS2sHU
0x2Fz1QzPblpk8qWgO4sS+GfbVLvbEUGwyOlPw3fp5M6Z8BYdqNMWo0RergpL0Qw
v+H3nU/5sJMbi5916yQFKG7vJv7V6XrAbJwug7POWCGf1rRnNoS+oKFmX0wilZOe
I1OimDh1g6VmHIccQPFZYGMxhZ1Lf/HIAugdHqVT9lvOMpks6RxmtZOYrnZ714+D
Q2t8c7ZVtP+qIPA17Q4WDfNQtn3QHcH3RyMidh54RadO4+n86j3Fa96IvXbNANja
GfxWoqTvtAfiNEX2F4Xg+h/AHkq+l0KtbdujNwU4/dHtheorAvPymP7NZExWPysU
8ypMQSns+i+0t15hLVXfYUYBO5WCu6tFT9xeruQL4qycL5DQZgH2dVi2i7VfHUaE
fNSwL/cdqN9yn/IODCCkfeAy0fEW0FKxmaVQLC2VhNazMA2Fwdgqb9KDZpoVRjde
81mphAd15gB8ec5c2ohBYiAxAl2zNTV5SKFhG3P+AK7ZUZodbJswJhqVNKCpa0Zm
DcBM8hn7/BGF7LNstzlAUetilwC0Exm+KjKom7JdjMusitBP+co3U3KhIhcvgFX2
6DSmYt2nkPklXdUKrX748b2EGKgdHlkhL/XnpM2lN5flEObSIaQrfoZ0CQexTL6z
XRupoz+G+NkRaS583i/iQDd9560lmRojR2CMAmUnHYYmCgNghyouqTVexNRwtMEw
hE3GhC4UE3JFbU3lzZRTkpqBcnU7wAYodc/7byKUQ1AWDDe4jrg0g1hBEMd5/NGf
ooOg/E9VOjJztRuEDxQJyZJSAKUBl752/HF+BbhXB1ygztDVMHctzEQa9h/2pPpV
fQ0jEUOCh0q6y9UTsGqGczcs9zvtPotBITw3ZCuQ8t4tyPSm02KuQEn+CG78xK1U
SX3DIQrLqWvRfOY2N0mGlBJV4faJwwjEkDdwTBep/OWLCUQjR9pjnUhrjMecpzN9
aref3zPz/vA2O6zMN4yn8Po7zlsBHGblZiWVhXOX0dkFC+YOfn0/mi2QTvSf+9dz
2BpRdx4p+h2QVQSKt0+qi1Fm2fPkFkW43cqgt5XPPKzf0ucsHo+ACptGgeCtuGiG
CXjHuC2P7j0aEt5AxzPZz/kAM2xeHpuLq4Qh1trx6ZyDdjg+Y3ll7b21k9+hDoTn
Mk14f6u86CJW4J7LPS5UcCGNUaIdEEZ6UU+dDtB2AvlOif8A8Q952vui1Aovcgt9
fiTGyn8z1U4TaObDfBtXtPLJ9sdOscMGT6vGBYmPK3UdoOkv7Kgsl2EyFe35rQif
4yR6KbmL0zZra8HB77U8KuRR38xrD1ii/f+Qhh5d1Rd1r6NA7CL5SDuzTIMBPIiI
VM+k1tMUpq9FBSRHJaD7d3nM4acMFsrFqRXqCEN4Kdprh3Ads+sWU/kdayvyo3+d
WvA1dwmH7JcDJ2uaBnxMjHa1hPCiID/Xc71Z7LxpO82I0zr/85sn6RNxY4vBvttV
52yDPMMxEUFycn04qUkPJ8ED2TkqgnTXvP8p7RtyabE/ub3AXYyM9mRZOYxglv4y
zwWpwEEY2xsfq/QLi1mU0w0hW4qnjaBrltz8kNrQrLSGWx7F/j2KP6Ro9mwEDq6q
kBl9VJ9RT8MZ7JlK/pe+ZGm6ie+chYNYARAPUQj2WsHbaHWmgVhMQWdFbk0N58T8
hcE0Q7VTxltsdjvsFDjhGgrxo3dbKahyIka9Vy7+L1sk21kh/YBsgqj3BQ7PMbi2
7xvNtb+pY86kvPyW9zmY3yq/Ufm1pw0T8fCsRb8iFrwpSX7GaImnd+Oq00xp5TCl
rmw7kkpQd4a0+hV4JRzOg8WekuJ6WttAF2POGgNtRghcH9uEg8D882WeY8yqdaIN
kWck7lylk5W9KpMjy8k034FyamqZpbNnTKGdGdEeGR22q9Mz8Z8OA8VYpvTdcA8D
oG+FZYZTmF9JVPK7UfcvAJ67k7I1SCdP2e2jRFL5nNZjCCUveUr1Tr2LvFNBhiwO
yDWEfD6z5N2OlwPC4H60guBo2kRZCNW6Fh8FmV+8qyczJf9Ea7Tk0bAXyahTwxB3
gHFQ4KBIsyXo8BcfKNqTAQy2ruGMXbgieefgw1Qa44rDlzv7myOhgKInPFBHTQu/
+JSZaCDobfoFefK4tRO5MhNp8hFw2NWsKG7sx1g1fN+HOvIBfSbxZr5mF+aulLje
IyE6nJGpp/ySqFI9wI5dFyuZrD/wX0gxCv6/9fD9J9ZA9AY6I6sF7ihhUql2Imts
J6rH2ovlN4/r28ximWFVEOf89oBk7KZuxBd9Pi2vCt1BI0K/E04b60ZHrlU1/1PR
c8hj2dSqRa9n8MNjcZfI43HP1QJXQ/Pm0su9ZXj3fI3YOkfNtnn1LNglCjroRLeT
PnK/7zOMQsmLtFPsmR5HSmi0HWbGaJLnU4KjWuKvWTEDRqLY1Aho9bGrg/EgEiet
OZ4ff3xxInuEFPN0Lfz8rD7ZlYt8MHY0SGp2dDpMCR5a+Zb/JTMpjCGT2RfjfeIE
G8c8Z9JbTFzqDv028K8Bm58vVsMneUh7mjo899LeGkoX0sBPYdYTWUlS6YfstatX
5ThLz4PUJHgcuMSUoo/A4/2bgDaflySd0JCnUACsOlP9AeuEz5+T077p834ARlat
qnQ/sYjh00eNVbmfqCnvJpNHBdyfIqyd6zxRyjURS2zzRGP5P95uHsPBCbCAoyMa
fyS7wDIYd0Dum7H8gRCS0M66LUWHbYMs3QLgsGxkeh2VYIpKfC8lgOlmSw+q4/Pv
FKQ27HRRn8WLJLk3PK75Iomj8xYIW+0GljzRO+ZVbvShZq3OChmDChkMzrCh5Dvr
DGsf1w62y1QlNPr2+l/7gNRjwo9ao1HP8MKo0TmkMeEhAb0D3UpGShc9kXMmS3UE
tnkTSf/pMzXitNrPOGuuc/A8AMJLyKONQPzZ0nWOhhF8IS1nb/iXllblAD1HATVw
/Du+L1yA/wColb7Bt1hcv5gThB0tcQC9n9EMOUJXACK1lVke+EELTdYegx1buke7
XyjZLeiWjK/K3pkAe4S/s4uRxPV3QvJnVWhlvwMGY7qim8jX+A9VR6jhH6oBbLWs
1uynys2cKRsciMNzZOi6N2a/Sf5g7Aed4DWX4k8AnJZrAlhn4E7jptC/c3Z7I4Cd
uAWDNQtkhWCA2CuXv9SIunUGk4mWl6iV0wgBfdkmnXqD9c/j9IVxmRFg9QgiTdr1
TSncGH/eW/8VZRfPuKvvX4yjyiHI5NPb8rk9vjz8xW1yNQkZIgbbnfnc8y+KVUSU
sY58NV2yNqU6tnpprgxCGW0RyajnRvhIiviMhnvIUWCjCZioN1BhkqTRea8nyKVy
IDfwAtD5h0h9q7oRtzvOeYFaAi9Koaylgr7GUuS3hFDUiPnhn+CRyWqDOjKKUEOW
//F7NiBYoOPftpRLNEC6xUXQ5CmDoJrzCSFh5HRMNRmwvtQzmqEQNH3avI5Vrqzq
/P4ZBnE8l3K3j6bAOPM76rIdGITRF8V5DMBedeS5tjyO8T3WysOSCYS+BcgQK/EM
LmIwo5IJWDLXRxsCy7NRfPZ4OSXZHuvD3hwf3ArW2CmprkPGcaQpNEA0Nek9NS9j
qZvR7L3VKG1euy4HrijpGGAX+AjQ4DbbGW9lnJnRzwkAJ1L0HcaUIlSFNjrjAFBu
7lo8GYol7asm4it8Je+P9UJN+Op+tqTTBAmcGBp5kjog3O8zg/X87uQK9J/ZtNlJ
q9VL9HeQiPNHAERDIAd4qkVUtAGutMvV0Cl7XZKo2h7H536A8rlxYOezIZO/Oq68
2x2odfHw23eXXW36EuGUYN5BjKv/7VzkoUofVQACcGMo2Go3uds+/3bvrvEvE+r1
KcujqmvpstshB1E8kBBNr/3MjrmC5zqeuqYpc6FOHVx5RVUhIdynb+otkp2mocPg
ujuForLG2l9OEEuGtAQsWLtet7hRvnvk8/xbnzOpZrYufCnVEf/zztLfF7/pjayP
Krf62t3WtXx0LKESIe5ct9Mwcff/mWExrMQGw7ywFI19XOdloL38zDVjf8OFJtjK
N9o9ZHlSe2q3kNouwEalQhlPPeYlKsXV7gUo325NtE23VznsZglA98AYsSrJeJi4
IGiGPlGuinHfKUwUrqzIqdvggxKRXmBIAh/73NBGoZvSY7lUoKQxGqi5o6xIO02K
u6JaJ3fvMXMpbp9dQv+0k0/64uILUtGSdDLU7WGfrhmVSKZXxmCG7iW8s5moufW8
QJ/spn0XgJMK72WhBUakB2CX8ZwS5CGx0qzqwU2qmAvXn0wJksmjbllwR5Fj97xy
JujLqzKD3N2gpiLBdHBtde4yEeTBCwLioaepX+N1P0gv8F7ybNuECwcS8th0PC3g
ws7VZfU0KODlVp7AYWtoYkhYlPRZQtt/y+wRpft13m5ukJI4hMjFGgJISd9WA7/o
wVSKB7LmJjjKOMDtA+ZxEjPpsYMcoL+PFC56XNYLXcW+b+A+0qc+i1MrI0tmtnCL
D8tfIO2uAtw7ZXZx49rCVUgr7LD/pHH6UR37c1M17TlYa54H5eu8JNwAQYVzQSfc
Wb4ScV6Zud79PNgQu/upW0igOrlPtittH9KprkOh/RK06HsyRsbJD0NBT4AljY5s
V13POnSDxQ4nElF3bLI04Jkh3qLIM7YBsu6pnSAWlRhX5hdxm6H5Ugpe2fxQuE7C
PFmGTO7mLhAp2xDZswciqwj5OrZqBuZZPWQ1KDCgUiJlbsVml3iVclmUnBt/GLJ0
YXvw8q9K2+kBnHcIx/SdeKWAPW8j52V/l6dfBXA8V3WTksOvIGT53/e5HQhcVbkH
uXgqNqWLZEW+7rR9ds8ybkFbMG5noaylgvcS9WNfsB9s3fD0jtXnqt/yeYmNFLwb
d5NKW3hoUSwt1FsTw4Y7zxkIo41jKrpRK3099GjTJIZnmC9w8zV4/azPii1dF2Kq
25mqoIFiAF26XFmxACFBZDe+fU/sraybrYBIOcmmYzWLge6WKlkw71+IzPKjCjOK
PyZVsfdso3fyEyHGXfl3CSXOYAUWzEmURlUNQA113b010vAq49czN0F+GwkUt3YM
qjXjP3jlat31WqAtv8ni3szip6P67FRgx/I4HPUWVGfD8TPRlvez2uMSXTbuIamD
DFTn+P2pMnyI6jfVHfBybbobJj3guvAdzKJAtiGP26gLVVKSVOTeCwzdCUfuAr4S
DZDZJMmNK9i/I6u2PUJ8nqb3E4PKJ8rXI6deoKZ3BI1ivluoJwBPuugSyoEw7f1S
t0Hj5jcv2hSMaa40m44WzkNbSqADTdBRBPZEemq+k7Xw+ePWe9UApv13t9K3LGvr
kCvn6/RG2jaG4kM9Im3a+U2iyviKSCtfBYgW6+JRH+TnIiL79eXvCihNWNBEHa6a
mVCYwVYW+0nWdDZTxMRzAxgbqBgcqdCv/Jp++MkIUwX1hQoYbcXtcr76gP2wlD1w
dMMWgZZVhJZ5sW1KcUx+NRkcALw9k7G8MmTtdCVOpeG9dw+nKlL763TNz9JB5UqR
8eolN5PEyn2FcBceKL8F7irqJN/k/BXjvoh7dGe5Hh/5becgI+U5Yc8nUBH8spLD
vjMJQMJZvkjxR7oLALxhdC1FdKiecwE8HBMiv+GWXwmUf4Zl4KWBKeumkRbWUzoi
BOXhCwGSQYtKRwwofgD+71BY23JrDSs4aHjWTo6FtwPuZzWTrl1bZwStCgm7pITs
aBL6z031C4aXb0ep8Z10waHB+rhu6BzogFW4F33gomA6vj5xSAHa4hQWoTtjxc+X
nWUUOOOG+2YJlz2GRnT5BXiN2DmvEn1PtLUKt8051JaIJ8DqEd/DSetpvV66452s
/I+/ZdLv9MC90bH2lm009vhsW+YEs9ShVoGgj5gS1/crEjOpclSmkZ9FnznYTYoD
b3WAxagZdluRS4X5lPSl2+be++GvQg928r/yplhaLi0BDzvRss0b8A2MdEzXizyb
jjdyhEAHZSelIg3SwEMspCDYGwZhQYEwtrowffAVHOI7JDfsuIu9BMoVOQMhI6Oc
vSvIgZOmUT/T5pwjBTtUacGi7Op9+DC/mTB3tLcYzBxanRXKn9hOLEXEcitrO23Z
5PSQLR6PGzofp+NzcSr+lz627XNUOU2ehxVn+1PqCbNVnPR/2DtP7jcvC/AU23pO
t5o2uR3vPULonn57gEgnWs3F/o/Wqni0/5R3wwQIYEfhHIvw5Mw5wbQsssKyvZ+w
SbEtAJv/92X1ztBvoGbqBxFvWQ4391QNAcvnZndJWpGzt3RyCuQjnTdw078+aQox
7J10cpOKFV74eqRj1NhQcZAzAAH8gnPdifp4RjXhNixrlQXjkNbZJimcpfk+Sjga
qUWBskY+dMFytECCAgCVPJVnrmd9eSB17Q25o9kkaMK+CI3Y2U/fLYe3JDcY06qo
SSgwAtGwXVEuJWYJiIkDazzc8KHhW8BnrGHwqqGIpa/NGk/Hyonu2q0XfUy/Aw9w
pwvX5Mo1wCqq3DsP9Jc8VTCXYK8eHdZzzwBJFhdaNt42B9JAcFpqd2wYV/cFkJgs
fWz0VKBoGMfY0TE7ay/ofYOn2jlDAHLXgRyzF1aN7yMlKFeOsNDhxY13AarrVFjA
UBXjbbv1GjeoqLZaVYHdjFghdcbMjmhMjGIOtWbySOoOWRk3KCU9TgSMi/La3dFl
+/u81imFV39+Npvn2UzOallNpxYkBMuji3EjhmkgA5xRb+Bo0PwovTMg5D8xAhak
NhT94+l7rb33/0JP90+ND2n4C7Hdr+d2VShfzbxtXICRcGbGDZq8pZDbZ1WYZyVg
e2IlY5ztgzISS6uEkqn8qykcupFzqLAq74rlRDNEvUibyM56tajBmaKoitxk3bge
SjfPOmlPvEP6XcqFb4bNqfe6gGtwhDLFQu7x1T4awuihHdlTgeTLtmOFbtXDe6km
N7eddbDxmcj0hUt4txl/Ea5vhV8Fq7jTGskB2e/3ePiKbN5GV2Q2rwQpKtKFAXAx
NOmUveqP76hZplwl2hS1FheZNalxs1kqyFeacfKoMqbHs7AlWWabwEAd+WJHsSes
iJvWJ/Pvcauu8gVL0vhq17gzhkdaAxE9eO1ngkosAyPVNPejq6xKZSKY3888JzbG
p0BVaZeR/3QTL6r81wMGmipUeiSdz839iQa1B3TNfkccwUSMw70pyHmDokkDMrR0
m5ckZc+jSzvN2PaY5KFiURANUlM5Ic4ZA2tHLdX3C/SvivqQT0U7rS9XyuLwPki1
Euo/t89KY2gJlNX3gups2oZSR83XwAn97OuvsO8AHch+wOIR4LDoX4EX+VeBVhmN
EhAi1QUXZeMOD+L8N+QC7odeX1sTD6JGcTfMIjWkQcxHSNOyKdhKpR6IHC7CpvXJ
Jy3bcIEVrh2P5uY2FWync4H6BPcGxtfWSPsbDRDZkQ8JyTUNPTkDIbU/HR2WG40l
fn4urCih91KjFL5rjB/I2ssyfkSxc7n5Us9VOJe1hZCYbwSqEixYy80IMFQIrX7j
XmGxop/VqxIVnueyjQn8dZ0EkW67oo1GsWT9rTQMvrnOjK4aeDVF/+zztfAFSkXn
gEdiQeQskm1zZzCIAE+veQIaWvrIuFKT0VoOWCtCW6OmUeCfqeLaNjKJRi6d/Kq5
M3k27oI7ojoKANpUGOepBLL+Qr7TNgUOMiZfOlM2+ZomWp17cxoouLRTm8AS53/c
107LfB6I/4rDSed7mpgfO8SwlkCceazCI8Z3ldfKE3eA0U5A4PwTxr1+YFyvLV7l
sCv9W+3WS4xp2bbw9vyWMPKp+H5OzHMPfVGAs3TeArbzfY9BDtueZZGpU6vVfGrx
mrv4lKL0Zf85eo7m5RkyVjvmUHwM3iHQlum+XiuPM44NvGxRLrZT1jc2tgMQRI3x
Oj0HY6SGDeT9a0wmGtxD0eyT3NEzG8a7zNmCXZDIc2IyV7I2Qqdz4P/SStck7rGX
k24iJKiIGH4U5tBxwhE90shPtvwI/3hhlegUje67h6n6ddtQUqYSrit4+wVskPPb
Ss+T9MhfsRoXnucpO4c/gkiUMpHgXu6qjNMS8ZINchHSdpAS4SnoON5NenwP1LwK
hgTLVgO0GZfWEEObNm9O5J9S7iPI9dxaM/+q1H1TREXE1YTqSpp2KruTiW5EmZsd
ZquPJF1pQhErllJW/+aBLW1O/G9DpLBgQI6u9PLnuJDAu0kW/KXB2+7nPwQ3280M
QZHCReKlVpcGsDComWM4LTiFafFTBN2Yjpalvbp118WIUwSE9hK0f7TcCwclMDam
hl1VwM1MeoWpJvv/prvxfrNd4gEFfL1NAshWpaq9HY/woZvgxLhhoAcUsIrwop9G
uJ/BjnIQ4YqKq5zUJUERLU/ZGipmQAW7kbOUN5CVCtAtDwS6UjZQQz+SoCCI0s/w
mp5amAXqYpQafN2Sa3cayA4jdC6B7HYbwbuup/76JXQY/Y7KzRRQWqFbulYhImV1
hUG8j9JkSGqNNNGsWZVqBpKbChHoZcLADOUV7Thkw8UhUNuO2Y6Vw44BRk7IWMMI
ZFCNYWZrwH0nVeNaW4xIuHgCetvYAeMTpnG0qN2aTWM/2gkOFNj/ehJvcvyeFwCy
EEuPddgB/Qn3nbGH3RpV4MVoJnjeICh8/fFyq5VakweTLUB/u0Cs1V9IEQz+rUQr
VvaEwa0IFK5pHT8zPzO4909Wlt8o+4kjysQRxmGUqlI6XtWs5Cx4yZ5oZaHqLDyj
cYINiDoMuH5mu9AnK//Ja5iwNnfIQI9c20UBYiLbm5HIbwI7qxsazLE8QOjNhMaN
4BawdN+hvRCOTfLKYh5qpUQ2Qu/9OD+zoQonTHlKLhBSAdZkT30LpjIjd1+vPCRz
1zOA8qAZoBauGx2Mb2ToRjwlvCcN5pAOc7QoiOJSpWkWlWBAlIf7/q/VZZjKjA1/
rbVk+Mx/pyxKrTSQQpGajIILc3b1iESvB50T8gnMsI6iGWSuRL2GbQ87ANYhDMZH
Dr68xaOcvfc6vePshFHezJ/mIsZ8uujdRWCoko+u0vRVPhZAvop3e4UPDj39fOVx
r5xLGo+6nV4Bpk6oDPf/XcJkHF6gbJWz7bWB7Q4Sqrr+lcFMyRRHb9CXhVp6jjpd
vDK+5Tj0PguUOeC+hhYhN6KClbSwk7Y7wuYGHntTGT29Kdtlbaqg6pTQDYIksOsW
VpjBCJrLwwx+k3YSZXFPH0WJa9Tjgkt872wjca9A/Q9HCBCCNyEgqVcPkY04lDyj
wjIGgcc6As3OGiDJYvhiHb0PErSA24w7vad/1m0yQiqAs5VSrKzyHkwZhXlRdFbr
tmmhIv0f+UtZXgPPA04aVbzbRZUlaGYoFT5jd25yEL0=
`protect END_PROTECTED
