`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ppADZAJVU+cu8sZkfXyPngvd9mOS05DGu6zgHoTiFGurNcXu9XOWWNTcKaTQ38a8
TpS723NY3CE5oyXfXnXzByTvJz5OsFjD5giUaGLFY9pXR4btgZ7jaQgEtzV0ca0J
3K/4R2yWDoMSJGbXNl2IjDJ4Gi1N8ApLiedtJowzPTDY7r9dzOnlyH/6w4Uq7vmz
BT96zX1DO0y6rhrp3DRXzYqBDF0z3rI6/cxg2zGy+q6bU9kaHwGVhHv1tq4QLNMy
uy6V8mnobR80K5ZC06/zIrQDKxvksvYU4t6O3VbO16RmHzgekxjbb2G726wJyXqX
gH0mhdrwdLtQVulbKGW6GXnDZE3zE12P/RSrah9OiIFBeuRC6+0aUnIJFXYjD6Yk
RCb6scH96UVslOBs/ftTCnaLfC0lsxnrv7USguKSPDf5Fuw5ApNkhVG+KPIXOxhC
hfgp07Id6z7WnUkISRKMrfZM4pK/xIwsGyuebeeexhXm3x3jjGtGbqsv2rdNONMh
j3Z53H7ijddouVcg4IjS/BFI0OEbHlezmkQ5b6ZnmVZgJZfgDCSl4FDaMaN4OtvB
7JaN3b0L7EpU7rg8t8QEqsLdE/yxqzwilSAQxHoc9XP6FY57XhMcn2uVi9A2QGZP
gJpQ6Oxd3b80qqsnbd7Ut5ol+jOXCdAe3lAHjkWf8a2hHV8iFgdEbAhcoZDK7+Lz
lPV6fa+w5mqwlVrbFOtd+Ffo6Y9ijB2RTVCxhjyuiCmR1TH+mWfGNoabF5FSvG2a
sWLfEEFhklY6UTKg3Q3r3ruyMlMFFt2s4F2IDSJEyZ20fCP9tgS9ZQiHBoQAPGXH
cZ0KqGvPzXrmiJpm/rXRJcdZ2wA0rvXS8+wqnGUk+lkkRRmgZ6UyPmJSwGyN0v3s
uz2hle8LBUMGeKq3qez3JwJGFVpKp1LfSMRtOFlU9lp9eTMZSFCEk0h1m74CGjmT
G6FgGIsv1sX6LcCKDxVn0BnvebDBCt+sRuzn5+auI4QC7+qKCILJsZBcyNb93uoo
8WnwCgBJn7iBtWXAMso/BXbspWXPa696SYKYTIQDJ7lb5Tqj3GP1d7zLjC26/6iQ
LZJ+RNCJsbgvGTLpYrymZqdO5AgUZg2mhOE5U3FGIvJfHqYl5AFjE6nJ5FKjVz4D
cODIP7DkFBoiu9wRxfTRqYvlaZC5QP8WP/Kyv7KugCK6PjEqISzCWhBspVCQF0Dp
p+yTjgvwkF0vipZwsIJBoHQof2n1GL8zDmIUKbKWursEWfksD+7pjVS4xkAdtf0k
N2xZRbaXcKPN5alEOhg/slM/UHZRB0/P/xA/x4kvjhtBTs+s7MM34ej2C8EgXhXl
yEtO9CywTMjVnfUNxrnLJyKjQhaBe//FXOTWyublfsQMfLmJ4xTwyKQ2FWoDinUR
DmRS/FP6c7nHQQEjRLvX/3fqHc+6yuH7gNZ8pksNFV4DE4IMNc6EinSpGwiElVJa
rQD9D3Yd+VbFPW+gQzsMUFzBhYxTKwI96GbhT4u/d7t3f5hxqnvd4kZniDSYkdwf
1TBmoBW0O4ZlacC1mFydXkc1k3tuhT7LL6cARjMtU9BHtiRc4/SoBSSPwVjE703y
CtKTiwwm4Z5jPHCCJNtb+za9Rdf36Fky9+8Pu9XCDD/PwYgMKtqCpzLpsSWf+E/s
SBtMtpQ48JA8BpPG9gnZDyW8XBLsxiWNhfTfE4oSFXbNCh0WayEi4QoeehmPhE5r
vNxW3xtBhP66sD8p+GvBhEQBsFNJmwfx9Q0PDwnJIHdUDdi91NKr+2ze0Qu70rGb
L4VqE8LbXu+3yLiidXc66JApaOcDoTasBVIZr/vu0HBqo+evMtT9gC4njz1VUnwG
w1/WMH3kl6X1kMjyFto+Jg4T3WADFX2n8mdSx5JM7CL94MF/SmAGqBDyerWoTn9b
gt790vS5IaPfgP/OwKt1vGOXYLSo8zBJyT0M3BsnzIiB4oZQ1ErxdMlBTd6MI5tj
q/9bXCxxJ8ekkHMdJ6tg1MikzvoRleN7FpmiU6IjUGlfP0Qgw6hKICR7iIYksWsT
INCUCsqmbLAVh5c+N509WtG8XNionRxhs31A3PaxlyLTuJ9577cAob4sc1opF2uN
UbgLwqbws78V7ZDy6rc40iwoDkNRwoGI5c2n9pIrTm/cjV5iPde26ChTe3HzqYty
ExAvl3VZLSDra+ZRVfwajamYcqwUgIymJQymZQJVIQYVPcG2J9ROZQbyIkX92uay
8qnvTmMBcGEd+gArvD2alcNJhLoFcGxYKS7R2GcV1gZwnZ9U2AHtbNjwe0hL3DIU
HeY1FsIbL1leeJK983mtkwRDNZGkXVLDlbdpauSAHzGMSSz7MCZeeBLghAaP0At7
f95hey3ah2SPLo6V9eXWhRNlArVGtJUDccpLwUzDTasv/M8pAb8y/aRvQUYevXR5
g1KtEEPPWlEpWIjzVHTf+eqahG/rOZzdNBb3oPzEsUWFstVdAzp8E1xH8HbYhu6L
QBqLkRYB78jwp9JnOq7zJcpBYuIKpfyR36Pi82glqPiTzRCEu7ltFFqaBKrNIkSI
59izgyqtsSaClXz5XOLXHBOdUkE0j1tAkGmLwTRUw4lUaOxA0E3kWvF9q8p+eU/k
qP4ayVOmhbXiqsiA7Bbg9QRlVpT8pkM8A+6NKlHO+cuH8Mg2Dekle6rKlcZZW8vY
FDTeFt1wkVKqoQWBGz7CdcL33w3b62yC3yLrJ4jzG0izpF+Ks1dadLJ2RCdVJB5/
84YOljs/CyTSuVJ2w4r3kpkLEpRP+uZNkj7en5FjECvmHB6ZNJyTersHwj9+og2L
kaACJlFnhbynyPxfak2ptwH9Le9IxpAwV8gIc6+LiIZnYNOLhtrnrbrXS2r8gJWb
MJJzFoaaVDNK6IeHZKtoQ62WIV2DZ3AgPB1SvHasC02mO5ciPSCR53NIVQzKvwbO
/6CMbMcVca5CPF4KwiWjL6XGJ1XAQBbyWGnCrDLu7kv+Uj/yoy1F+9iQ0LCfzCR6
ybM74kXsvhmsgBfqOQ3nvXngqJ4fr5+Jmubzxl4K6+uWZRb6nWU3RaLXN26REGKo
1JAzlkBtJgtyPUAZdM9eblpOA1CWFyH2xGx5MMcGy4SvUhXxiUEPbVpLJU6ZVT15
x8mVZwMKpr+v1sn0dnWSyRPUXcnOdgn43vdDdTvcLrkqOr3PJ6yobAIbhJBUr3BK
wz33vhVc3FKZVPyUnJO5W2zNYSZ2IVrSmxY/t0lhv381asXLTjwuwoMDtN/Jf1gP
nSggzpejDN79UPzUUOmnA58SGHfqzUtSSndFZbHPWAsEB15dKhaiSXRUR1kJwC3o
ob9uR17FJpNcWEm2UHexFL/Xw2JQ7fj6UVZBlIvVCcTManhg1gxDHPU0mpkNFqki
xWuYLRbTqyg9ELXK/m/DsGINszhiamzlCJQwT9ooOveZY+rG8PeW9ZPfcBrcTr/I
fjzlpXP4MSC4fn91zq7vQelMWPJOTFyD/Uzz4jTnbGHJzNa16GJbSxuN8YnSrF0n
1VtTP9Ktq3zNk7tU9O91M0KDwOeMYhzaY/ULwZMgZiprSDfcrH4FlMza7SjMwBWd
3wzE/IJGHDfPo0wfS8hPgPq/Etm3mR1reTL5jlZNVOknlWsRK4xxKHVG+H6nDpAb
Ik7YQdrxj6UDNj8Xu0oFZfu2f2TIdb+QX8ua3mfrCXDWx1maUNuOjSifh2GQSHDP
N4xDeqSWnMUxtFIsSM6pFYAVOth+K8me+OKMfq+0gDt5AGk1qHx15om1axXV5SHr
9KlvY67zj78p0mAe9v4MiQWNvybJswGcb5xkksyXDsrursA5LuiUxtxgA9/hEcNq
46O/qpK7rgg6HnJjX63ERqUqVT4P56/InOvCDFED/5yTF8N+/kU6KgRqHl4UyBM0
Oyq9Cnc3p6qI5LtNHtD18lzC/JacSygbrxf2vslibXT8j/I5BKY9jd3bBANl9oa1
IyxD6YYo4SXPTG9LtzEv82xeqVP4jp3SGYqZOUJsC/tzAgM7EKQR+3HeEO1Ibj21
QCwLNt1sXDw0FE8WIpguVQm6Xmp8iHg5ZAF1tAJT2johUEFMiiZNq3Qr44neOujW
8QIV3JUJirNnKjOnc3rqNkFs6/inQC6RJyjHhTzZ0vGxeEZQOjQo1oKkij7Gx/r2
burclT6YXS3XZdWGvv0ty+6jNCFf8iVCByVIu+vY1guHXTWOnMXkztYr0CNUKHOJ
A7HPBLzqmWUnx3o0K3RLpdq4iFGZYLjjwXXq/2Pp34FW93WFUROdPZ84/XzBnCr9
FRevjrpkk/dGFBVYWFPFx5wXsm7gb5q5s750UnNkUO5guvLu3JGXz6XWGIe3cW/v
Ox8xcZsXbZZKveoT08lWTFVCPQS4vGmJUQaTP2ZWNgSEcic8e/UOG4KcdaQ5jb8i
PSfxA1TRpFQbTnL3e1ouaLDf787PaUK01zfXMmdUx8sohMTgVXYexbxK1FESKrFq
xwCRfGVHLDosqKmPY8fTNhFhvSJqzwWBSb8Bak7GFh9+fi+9G65qGvCuCzzYhAb/
LVDS3R8eAeDM57z5yhrOBVAdUyT/kCmRFsd1pdG78twTbVmeRN8lCUZoWUTqU2xR
wTxheLrRmhgcE0yMZ6OwLc2BSEKKBc82uxU55/GLFvBVyYH6xzrNeggUB+E9Uj63
xOdxyo8sQb1heMQmkv3Z4xXL6ZN570KDo3F3/PIzrO2NgSGknvEAg94/5lhVFOAJ
9GM9KJXGUn8KKGyyvwRhMQ8I58Oim8rzhTbKlIihiZQd2sz3cgRdrzAq3fxjO9d/
/H585QT7gyMDEy/m/M/LIeatTvNCHiC9U6hrBawZovHj8pNvxpSfhXO/Dj/01ZRm
cDSGAYw5a0112TGQZ6ZWZNqwwxEmS9jzAWvzpg/PpgguGF8inN2oqIgoA7+U69TT
/55gTbUEcC6CkjXIkUleNnIo8J1CIT3Wfc35+bk3UL7zqo4CHoZr2pKyvqPyfvzS
nqtDnoY4G3jl5ibfWG1ARBS4X3XRGOFfZ6Fc+70VDEfIJ7HVif8hv5kZKAgmC28y
YTR/fdL2MrwSCIMUutVsXqv23nQSbrVUQPRV1zzfKdJ8eDCw9rVfgB1p5akYSG6s
7ssVXnB2MzkUMmK+2WHHPCGB3bhcPzIjzQJ6TlE9pEWG9tiP1D59rzob/ilc5+AP
Z7Q4wpxZo35mBawshvxBQvqNUIZZO1MtwBPtrb4lN4tlbkNnm4yLcjrhiigCIgeR
y+JI3yKsrzqVw1hRAp+cSX3nznmPDxKSr9XusRCTrnISLeRvbLzjDJIFAdzpuXWp
P6HrovIxyVsCnpr1GAuaXtbPdzYHjPgWkCtSp/kSK6diqkxfPinN0guRyLQO1hZS
mGSwhRDFSwMqefj4GKgVi+X2dBA3X3mmgY2JUqpRiKSZjGRtOPFf9yjC5cyCrDwJ
18b9aofi+a5h4JN2+YyXnXApXp06dSJC38TNfkZftEv8lpkTP+B2+ZURPjdZr0Iu
pi+VYDF+tKBBctLWFo4yl0oXshW4LpABP/+b762BpGq1Zb8YI5GLWw6Gw2Mb20QC
2kyJTKmZ1FE4cResuEvWlHK7EvWL3IGP5kzRa/AGUKbNrEdIWiUzPHNdr8UwgZyR
zPR0OVpi53q3VKj3XF2eroIatzFOsP7Tk1TCYfOfds+dj2UD8XsPX5JhtZfBNjpo
uZmr0H1Mikd6Tj3Bbse7XLWp2UVDyimVhECcmZ1nGeZz9cCWxdgYkYzoxBLIGHjZ
gqVnzhTYmLd1G8VIjFALDFLGFPjJi16JD2FUbrQIekHhJsUauZxNtcIAYinWxVyh
v424fZrjQt9rwqeE8++ujLEIVokdirckvO2m/bzUh9bv88jcIQyrItFlFbIpmmpX
3P5KyDsH230SpzpiQGuFUhPT0/hfysfraGW745uwKuGSCoxtBod9r5izTE/c8XVR
uF9sio+y2QcTCSXx5aqyzuSpUo6zIKkv2CSCRPCldwDtM+LD8n4s0pxgchdQ5Aqs
x3oH5ghS8d46EB1DXE3wmb0w6CRjPudaa2mTmpoGT5/jTLIOrat/DIl2RwjSiHlD
waROM6wsWT5raFR8keMDytY81UHZavBR2OP+61UlbWw4fTy6lPkpG0S6EDg3RJ25
KtX4On2miy6JySaSviTOyrftjPYHLoFdLP1pTjvpl8BNyLqr5r1OknJmaJbbYHlR
KytIEvaDkQStKMmS6DChXkxZDuSFLKqk3dq2RL2KctH91AcoKGkAQpI0lhzZy16+
ID/ShBlWx7RbHu4x6j0GsXV4YA5e+EKwYqQ+Z31qUF5HPnKwr8Br9XeACgZJapzZ
iQR/r7wmVhSxfhyCjqEOp/aiPm0rXYZLs3r/d3sGSdGYw4wH5kMt1w7RppFmqg9t
LW+TUthAVUCFZY4fQtrMlvc1WZNZbLt0PgouY9vBDr/PTQe35PBvVrTsNYBF2NcT
xk9frJ+7QuORS7lOlLZ44j9ynhn6NE1SiKOHZIZPBJWPvwCa+GgVBDqIMFcyO0qT
sQ+D39H3Nlv8tdLaHz2qqg1JJVS82XYDfRrx4h+/Xu0actj4w/BWdyO9XE2JOOLE
BK1hn7c1XQAh5EsTvtPA4+pn/zaoW13CT9hfHfHTOGCR6se/yTlieySU6/Nf0XYB
BX0PR/WDFkZARNzeDzufFeTeLZ4W7IFKDcMGd1qPI6ug1e5zt22h2hHH0HGszcbx
KNE6MmVBNSsuamvt/b278AKcwPwhJRAxVfyjxGLCmEUAN1BMBcsPPJuowZqGLc8g
CwZ0t6gLuDiKyPIMj32n7D3hReUfDcN69JgGcl7i08kJRLNss51tcsNBchl5vVP3
XoLKKXdH1vFgtY79Wqi+aXP/kVUJz4aIrqOviLFv0/xH4G4wVzG/JklAAAHJBrV1
jkqdMRf1WovTi45mdVAL6tJnbDpfNl+rxWhanR5wdk4aDgNV/rIubOymRPNcFmI7
1vIW2EZc9yDRY9Tzme1c/W/mF6qa9k+ufW4h4YBISdrHDw6OZIZTNxLZCcGeyY8/
0sHpXiwfEO8oYfKrVBmy4aJ2k6ZalDaNG5rz0Q/Tmu4ilGii7DhQK16V1MOawKit
gkT9KKAg0r5SIlZnXWyEybalvfBB84upcvX0fTHsAiHXK4L7ZWJYIOB2FUVRzg3s
vsJ2I+G91wUTpuzrLOubJQist8ByUDUL30zJ1Nos+EbFFMouDidEKUNe7cmhMFc5
DyL+oZfFoEc7YFKB5fF6NPIUv9J6b9okdGzE3CsjKd7oUuvgUwA5xMDEWqaVEzKV
vLVR9xp0NDrA2KBlJXbSvq70am87eQdMzgcNAilCnemFPsg482KpMfYS4r4sJrJZ
7HvvpP22v3MBWYzltFx02Y/MbVz9jrvEs96B0C2YQQLcHRUbe1ZAbJ8QlbPbw9Yo
CSNHaD005Nk8FeEFjyBZ9Fu00y78waV2k1AvmKXr0mdpYUC0LDnj1GfysRlAjO4T
bccAPRjZ/rBzMt3bnrnUeRXegFK2cuiI3C/nYLixKv3oEK1GRSDH/dHvTf5gk0up
+18WAPQCUQczNbAcfQ8ssEbjIXY+RZAcErkN9L5RMeQXxWMDkgUJRZVTAo3dB5PD
8mU3YUzNOxc8nh02NL/uU9jE+PJn8vEqu8QHLcCulNPyny25xqCiUqebKO5G4HeA
MFdAdmt4dX08V8d1pSAILWaXEhFQaloRpSM9cuv4Hi8NWOi1TNFKc9XlFuUdJT0T
pCEurfPC4iLiYCLf9FbHyrcTsfHmOUpWD2KVgD+Z2bV/9ZJclsNN5T5E4V06fIZl
MuY2zROFDtr4yJ7zXlm5/Y94uSuM48I6+rglWHUsXguXSqgiQKotqgbS/rRWChav
YFd929sOvzJjStfqEAIWMITtpYsnad296bolZS6vjtIQGO2V2Mr3IxmsmwIclA7g
cvkUT2pyo2P7RgbCE0sGFR0fVUVBLO7SsiJOrs6ba75svOuzJDfM2pnzyqx/ZvPt
MckBZKOFjeBaaIvU4PcmbBoB2cxKKMkshsh6BO/hv0rlGCRs2BDnFsmw0RzSoXko
G7bpCzLNTRVVLTLEQyD0MkaTvvVx9zCnU1qFij1BqO2HnokuJngFHPcXVDScp7+Q
lnBz7YMl0iu80vaSZyM0uJSTssE/oicK6fWmH6qUVurkQK4mfhHbtTbu/8v3ba3q
EPbytzOoDExGeuw0fZLADAn5vbf+WtiTu3OmYz1c+lZokLoJu/A+3rIc3l/MQzi8
GXklZ4JhsXp+Dg+wqt5a+ri8xjy+muu/SQDGtRJOPvR3j/V1xZwRZ7OVWb9lWVF2
e6ZbMatUjnzWzolcNt6Wz9VOmtUfukVfYX3qGaV9FiLZwmR2+I4gwzcwvynXuHJy
Qc6lcsGV0gTzZDg0pzCFqZxohwvS6FYQKLREWHvgvhvJmCUj1DLiV32NKlYr4/oN
ZuTRozi8kq1h6KtZbk9D4GyBADa6wRbP1pl1OeQFTDHYD3JFwqBnnGa5Fn8dvnTA
KyAsxQi62LYXVPDumDsI1fOjg0xK2G7LSLvda9My5fNGOImyHMrpW+9sOvptfrKv
M0wMce3ODaEacnyslOw+i/z1y6UFsMDJXt72WNEbxhhapNKt66m9wASf6f2uEySF
NLHTbKraYHMlYhHUVn/v/f94rY2sw7sd/PKrPLLm4XCUAt+gCL1nyEgR7IZD3NlA
U/WiLkomso31Kzqtcu2dhaSD2rAppmQSP1cxGTYW8RGh8NMeyEcj8A7MmVSZWQoK
S+EGn+dmGNp/kT9ds0WPI/PyPbiigbIOAXovQhl+ZprFmZZawnXp2Ld94Al2PESB
wFPxmB0PAoYutDVXoctRs51ZP+ytHVjPnfJHVavOnHmVauPDCLCG4/1cxDtjKDrM
imV59tw8RFXmTw/ZBNFo/u5hFyQt06HsHBaLnKaM1r3sxcPq+7TQdDwIr4O7tGU/
nJHCnSBz1O5RSBlyguZbdrd9GmfdIESvy7jvC+jC6Z1obEGLQHJ5BP8d5Vh19SNm
9ZG39RZeBqDbsvm3JADMSYdx+ibqIA8z70NekJ0w6ijJciMvUih+3sxwxHP/12ZQ
2gn+R4dS9O4StwL0yJPn6eZW0PkLrmDBJ4NLPxiazsa0bAl2SzA2475Rubi5sTtE
JdPqbNlcSAP9QOkh6xm4x509WM5+nIuRydaWsCJdwb/lPZ60JyiYr+tGzII4djQb
jBk4C7aCceHKlERxPRx4O2tsAJd4E6ON4Qmy4lVXSBhNKw72itZTNCuCfeorHGbD
6SGTx0HvsUwRbZbGKy0gjAq2UyWEq9iSNpPJGMak7R+aXTQjuTbjYaa6S3vCSoey
hCdSs7cCWqrg1I+hjY5XgXp/KZ33y3izVL7nyTEPidgBZCfmlVHXJHH5mkwzhs/o
7FsAtmSF9q13skx+PdgQSW4j/97dJfTBIsV438K6m/U6huMngeyO1tBj+1UKWi6/
UYlew244pw9K3WIgXdzxicPTa4EOu8Bdxxwin+/5UT1LrG/+YcG6Hof/Dj7XG41x
UkvvU1VlSTdfhA53p3HeiYHmZY5IUetU5oM++T69KmlnKYFpFMM5yG2qOvYGVV7E
UqTwUINyYiEHZr+wbmMPUCxeu056B6Wfd9VwBxCfG0r0wiKmCBpeOgNR4nc1eyq3
z4k0ogNYXWL45zX6vmBFmKj48r7kG+R4zgfMIwn6nOZbYLwwSlR3aqUuaZi7rmXw
0h6lFZeM8YxVNJ3SOMqsbJLgJbMyRdVgADvGrU2xoQtipxS/lgmidm5E3B5bgRd2
zvn2GOsdORCcRJzbjtetDfOe+fvlJ+qaif3NaaxUIpxmHxl+ad62tgwJIoSxjjfA
XvC4QMIW04C1P7McCAsws4GPUwv7ogXekdnhYFK/bfxlCB0eceWky+ql16HW7R+J
g3j0mFYfrZNP6v35ajG6a4FnMTY7DXEKuxkJ9emXbTEfs22Qq501A6zu0I2Za7Ng
QZq2kOcBhDgzbRVpux3sBhhLmSoHLyytEQrV+KhUljhKsHEB+gASccZVWo/h/mjB
K2Jba9M1Ydw2TSP2UYbmzJVYy9twuzajFGQCcrZcSS7Yw3H7KsZbXMEuKMDX+xOv
nWYHJcmOoIP8TJbt1pr+h9Xo8poaYS8d6JDlTSMGVJHs3mINGlrAcwhLUVF6Y5Tx
eUBjueiiFMupP0KOQjrwQi9qPrKEE4jzaxPi24utHDiRg+Uk3WzrqzrDp9kFmgF3
CWn9jM/7eaMIqcz9dayAcWEzlSoEuhE+HBCqeBy3+ru67JDTh0rPHwEo9hh7jWhv
Xo1378iUnE2LgyCCArYN8Ua/uvxSstgEczLaBBm8t2OcFh3qN1G6gP9tLBGlL6FO
NWYQO4q6F9bm837PiFcLCsUUKMvU2Hevl3eFXzTD3wCrT65XWmsyskj2Hr+j0OnU
hWJxIsvv5ko5VTisaumxRfXWtexT/9cO4/qQyju8SGDg3B1kq0MZxTePZ/Jw7txG
Phsiuhz/RniNKPyCKm09Z/rywEK9vREmT3XaV+XJjpfT0dFV5krnXEMKBvXcnLHi
9jBhHKmvlYi9mOQoQYIH1MbbHwWCKNG7IyMSEXdjVZ4SNtoJDYSSb/te7U2IQmnB
csXvKXmu7jLy0Yht83uVmgDlwFtCpATn7pbJ3xEdh0nwQYJ/aCpicADF7665fYrW
M1F1vp0tVRBGBA5dT/awnd/uUSLvf1z6foGmtvwK64R2xi5OMlkwWgqUyo4CN9sH
B64a7z2dUmIurtB13IYx8lQJknzCuG2SP2C5vunFTACXqvHk1qYZt+5prk8N7w5I
QcstqThdkUo7kf5DwrNUZxRxukQChjBCpZux3b5fZwypDMTy1Pdt523zBR5G3sMp
O5l5ZQ9rUWXMPThScOKdl3Y5GfBoTLh9KYmSB31yYD7LcG40BFcwiGCFK5y1boz8
YaKKbNrBwhVO1lBPH/QIVaF/lGo73vb/mLTwfwGiRK+ZCILe86vt0YzNySU8Nr7t
yocNst/6oiYb9nmrLz4JmSiBCHoBY1qoXggoAgLPYBA9VmioWlpjl9RdCCxSMVYi
ouempLWUSdw+CEPs51n5zo13jgK4oNFoQoVoM9nhcln+WYbhLbZU1Uo+457M0/+w
mEj7vnkG8JZXoSo3k5O7R62SsRNICamWv+lUFrQxMZFJ2ZfoJCCxBW1eXiAvQAw1
qyYBL2Q2gU4HH3t/CUIy9mP7BjyvDKxeXEEuRYYUq3wI9iD2chJdzyhWGxc0l3ZA
62k7uu5Rh1hOprmoFoDDebqJMHXVjW1PmrPXXiEQWWNT4BXQegzrk7gDE+u4xbs7
14VKWZYK9w7m3zSUfhXnHZTCd37jkJoJLQAjDG4M6ijLwmK8C5I3jX5O0lRvFL04
MrjCtsLEPXlTe7FqEFBmkRTfO0wEjPBEi7ynISuQ5+0NNY3woOTdVaNza5S79GPP
BzPfKdwPSEXsaEUVTuvseKUZOKWbqkNIWFeT5tDllLZdZYbSF/p+n2cTgVuIO+d6
mPBAnUUf4fRwimHfuQN9nC9qxZ/hAPP0OlacvarBoIzMs7dno9xBDqjR7wF/BvsG
gqgS79+NQQ3+FNZlxF2bFTkjLr1KMfQOCwL7T0xEirRu8BwV/bG21RjD0Y0RtSRa
4rtZKEQnhKURzvqyaciHURGNHkKFlHVOHNP8Q1XNnQZWGgjtQ2O5DjiPbxy90z3e
HJfR6K27Qwnq16KyJi6JlJZuc9M7Dw1q0FLCs63ccRqa3zsXqrzFRwMa0mWTejsJ
R4s5RtCSWnRv9mzdZvUMoCYRm1ukF7RhVm+V1qXYnxnKrkFqZYrbp1leWAvJCDZo
AY+DZgZm81rpe5a04Jz01Z3oOR7rNpYRpMBZvW/7YXpEBEpCkzGSXcRoUWHfSyUi
PEAq+ay4gFzvsAS+2H+qaEkXe0oynMniDUJ34iGWOwIZc0T+ZuLT5ITTfm9Ip023
9VLan3pMFs8wLKHSrRGeqThfT5POi8RVzglCxIEaAvc0Uu8OCPJinn9lnIZDYUPU
GAwf9H/sgI4uKAdxmMh5kjuy0lfdfjprVU/7PrdUZgjt0RGEgps2jn9P1EHJ0Ri4
38wrCuKPIqOQiGHkb7cS7/NLTlmHtxaqTB+xTD8u0SfnlKcL3HMh/20GS7NzIe6I
Mowx1n2utylY5IPqi6sjnAKpUK+9S8Yat3p+ryAf7Z76hwM7G4uXdSROpZctrLlA
bX9IYxsAPIMkwBGK7/cmLLEyddhqOrw56U9cyytUYrKPQpqaSIRPrM0jLeneXOL6
3mUE9WL9sqWQSgLpxQHlW+GzEC9sqNhSqVDtIJ0eau3ZG6hS1Fmk6YD4NzGYCUsG
4xEMXlNSmKwIM894hQVEM22bYpyQbt9GtI/Au+c7fW+1k+wMIMVUJp9Wyh65sCoT
2/RyVoOynehlkrgQFiloWsNr2MJZUt62c9/ixrk+A6V7WCBpvgmJeZPX7dVcRmqr
lnYQ6ePNBYNPbAdRvNsFOxrc6zMp0EegRHqFfUVakv45JShwsB2iK4aQWdsDJwbk
2swfdVg5NEA/D5futUPlj7y+QQpSXBNDsaArQFRvv3h742s2t9lCwv6uP7itVYYn
6MH6g2G6exUDbKePULFUCi7dfeGofd/u03NiswX6c0qC+JEsejgCLbiLSxkhoEsS
KsQXS7LOpIAbH1QJpJkTHZVzctYmVq351y3phJJL4IRHNfr3w+F039YZ1l/3dFLD
wOPW52iXP9Z+J+NKyYTiXTX2OA/JLPcXVSDevch0PlWwIfTt0wmss/YYLn7NHWNk
YFKSl6puNmMjsKdSj9USPW4gt9fKD3pXN9Jara+qFvtyOJpvKHUg0/74smg/uBEO
SooR/Yv/uvUA7GNbpQNM8sEpQ+kt5qwGETs99jo3pwRlN577knttzwwRn1GOi9D9
qg6afbCwa/uQlWQ+BdwJYOubolkuxBy316lYu+qunEStB0MuRmdZBC7sD9rTS0i5
AgYASQofhoVG4M3N0JKcTU/mQcWUdoxbL8LEJ6s4KaVgMFACoisQxdvf7KUPoU/+
s1T9h7mOhd1QmsrGzEwcnXPuvx04osBlt0YmwDOLPGT309FuWJke/FmM1v04Oq0u
BLd3/deUCb8ZYPf3smFWdznK+sxEkcvwhvfWZfpQhxQiusDYP5tuanDZa25eOXWD
aP/njuGrjMGdLXetE/ZerOAXIWjilLt0+ZsrSqDvcPZSuxCoXBWlSScFuzaD3n1T
C1Zz8uMyStVsbdBHRrqmXbwu1kGzCaNsIGw30th4zcHBJKqI0SG0RW4oX+eL7DLm
mHfBgG2FGJry/8Md+kXoxrH5mgvs9aJriX16iBy5YgNv+eGRvoF2aSgLF2F9C06+
92eDpjWojkHn7ANsVSCFHnH2z5p6nMKs2sPvMxCXuL2bxAp6Qxc29gn1TQMBQRzk
J/epzcLNEbFeuMCwSth/6CAuW7+kUwzjTxekkOUQNkVIlN5hVGX73NGowRQspOWL
QxwGg5gbommM542tbbQVmqkiK7qgyui0buowbTHS2S2G17aM5GbregYjKayG75TN
Ci+9FXBLroimgTNomVPL03G4ZQduzhcacZT63KPmbypq3TxNytO9Yt9U+hn9vHV1
tJz7EOTnlty6UK8YyvGHRqeG6EHF19b3DQsZIEUK3dozisJSOGWa+ZGz6frSeCaL
gF2Lsu5/l4UW8FcMnHa9QOOV7v78RsXOWY+bi/6oIOHzM7mMM/6EwfNsDyMQ543I
143zXvtdkvKaOXloG2brspgRv73UdpI/Hg9crgqHyzOryyxhbcoootzkftdpo/e4
oa8HCKUX198LGq/IjDqe4zLQ92VhvDoJ40Dpx+/ONE1YW+j8wbMSDrXdBAIzkdFb
ZKGgCCpOh3bM9lhowHjIZ1QsaVsqodUx46if1i9/yLfZ+aK50/gWFey0ofTAzrQd
c/tDt6G2nGrOroVBrAyDdtDczIdUD5pXv9wXX43USlk780FORnCQtWoaHJjFy7Dx
dglZ+Lg6mPzMclNWIF86Ie8Nq+cjzGKOmivFTeMxpIjbk5bde2QH5nQmBhpSJpMO
T9PdrZ1XYZphjWYSJPhkW5OIow/7FVRX9+XBvsKZbDLr97MLveQRY3+ZToSI3qex
W2s223cts3Eueou9pNsTaUj59puRoaVlyqaMeJNTuCz2CP8K+VfeUHVSG2KK5gpd
U6a1XKOLpWtIduiZAd0mff32qtYNf0ySxF6qz+IBcbk7pfCZpVoptXHCcbjZyH1X
TVcFY/VW9yaKdgTwYMVPdEfxrTRCV6fW77C376+n0x7rl9Dbm9CKq1N2mnJhkO9a
BaecCtK4j9zUk7F8QJzuUTuVW0WQVycbZBWq00JSfxQetaf9gXiV/IZrJzn3fsme
SOUsVrDBL+V+UU7boo+X+Mf7ul5hKDSpv9+AXsUmHD/hWKaYcELB8gnwtC3Fxb5F
M4Gscos5S5XDjm9W+wU5HNy6nWIB+0vDEOE2aqEHbddwEfP637ZmNB0ks53PVJ4+
4ngw32XHQBRRrDbwzSvv1Rbx+WnGMzB9BEDDVhpkvr6hwhFaTKeQdtiTX0N3v0cr
OWNQsP8647LrlMF22GamXb/lWE/yclC08dmy5GSm8bACHP0N3MuCXfJrDhwodIha
NaDW+tXAjPX18Gk1hiuojEz/O2LXF9MtjgikDxrpe/RtVWwRrCcS6MatPmBUACKA
9EjvtsENWb8Cz1Vvb1i2KhPYTchOqgrQbiULZFtyES3AU6h8MEJ3TclBG7Ua1+O1
RTtYWTgnqKgGsqwEryD8PRUyY1NcBmfCg/gDnxHJ8sqCrJQscWSxjmUtvwEudMWD
X+ejjoenOIW0etX8HCRzk6XRNNUWsK5YLdNKWOBFdjdpAokwVEsoNj9JzkYBMUxI
CKHxT1ZnJLS+236JfaTExhEZffsFEi49EHpcvAuP4E7XSkhkWHmYd4uq6aVve6hr
YKjk9bzJZF6PgU1fV7BpmxUno/lQ1PdXB7ipnlvoE88xGX5o0W7s1E+ByhC8LsjY
sAmhJSKjLXsBYmhk1uQUy1mEwxhcG39/cte2gVMwR36nrROniF/W2doxlyKLVPny
9NnMUUxyZKxB2awSTc/lMDReVRIY1yuCmTbABg9sxqqBoyB4HVldsISqRkPQkxK4
54I/RI9inA4pGR9kZPJfL2e3xXloS4riWFIDvAR7i5W5iUPqtDeeQH7MUE50pprk
LPLWM6ALerYQzM/BAcqubAWUIOCluvXQtqXjs2EKcGPPdT7QNaFcDl/aijSK9sA7
QH+8zLiAB67yVkdIu6T2L/E2YRveCr/sgaE6xo40vwaPwFYVzLvKR5HSZzj+PQ+k
tSp5kkY7ZMvHhVXGE52O2hEV7YtA/C1tqJxNGD+s1O3ET0BwC63PXTwUN4vf/HlW
jjEaUN10m+3ZU4Ezd0/d2GU2PlPTYFRIV6SHcwkmmZmLAyvTNHTRWkWDXcQ9IzAT
yNJjtxhPMjGrEwuvT7sBuspk5Yzahpoc0og3m8v8vFVQu83pzteeEBpobgsoL0hy
L/nfHlQzN6MyU7t864HrJqZnNc/rSHvY8cbjbONwjZ4GsKqFR1khblpcbqCb9+U0
rZmXzd9ioVfCCk6HO2TXAM3wz4DY9BXjEq1+Lm17ihNNwFT9pF6wRDWDy/amqrKU
kz2wQkls56V3OfXRxaAQGpSauIp8NefdQiVuChlEoSzVBbblW1h/jFFT7D0HF8E9
ITr3wSs2mtIIf638UCBi7nQetRGNGBScM4oSPIC5ZyyjJZ4nQDbaynjDcHjEaD7r
coXYROyso3+DJ1zU/DKil/ZfFb75n+3eQrFYF+ncZRuCgyafJPYQu2gIpxY7iQBH
PezEy0CcFoOAidxHobCn4/llQsvbhVY2x7c8uUsTdPM1y5M9lfItav83kzN/4WV7
UecCEakvR/Rrb14VZ/CQR9XBqncncw9OrFlnI/6X21w/qENw1OvtWXRaDumm9hdZ
iUp6gFFyZuBmIZnooQXEm3cVcraMCiNrpYyzARs8crhRrr31Bp4EPnCK4SjO0/YF
0w4Kj0RuDg1aEwJMz9yMXq58+GL+FsSwLZFypCfgAYZt6Mvfkt4Gw7Q4TGY/Tzfo
2yJ4aAl/dB6E+Cff302OSK9BAf/3nSs+YSmRp2TlHW4Fcd42gu5sEdjs0jhTvW8w
6hbtWZ/5vhIoww5XP+cOrWKJWAMIQs3aFxuv346vCVd9bqH+B35p1eNZpqcZe/kR
Ky6A/bI2RfaELjS6DsNICTXCvX4C47tn/3sEya93jcaJpqhxYEmSWjbaQql7Eh/g
C7YozFSJBXyCoxKBvGLqNGwF6KToABXRGSUx9J7p14ooUS8lFQo5D2jmGLhXYHag
UCKmZnKzmab3BbW1xh35Hn+HLC+gJ0FHfn3uTGj+37NlS7Hft7AeIFe3Svubam09
kihycLG2zBc7gA9FyVm2lkax4KYRAZhmflqUu49jpmSkISZXaq++h5tQkJT+L379
Yc6G1pmvFapAbdcSga4BQ9d22SKj+lCmtZQE31vw6pltHeHueXowQg8YlT0CNxGg
WbmZZkAN6DP3S4+XXIf75Ve9fy8SQwjuXnEzbrLyLYpXxgQVuWufqbvCXZ3UB/qt
OhafBP2c02IhSyvnGDUq4ByECqDIvi8M3DOUcMvuDZGfu57ymM/MPtV6N0quood5
x2bG7Dbk+c5Ehun96w+f4/W8vzOn58XZkbV7HTBz5CEEHHEeY/DkSgH8qSXh1mvP
iaxks7Uj7dvAl6FhhairlaIj4LQziTOzHegZ2vR2s0OSyBqx5cKNxCDsre1a31dq
YFH2QZG/L1UYt5o1abLhEiETJq4wsHELmUqtmwOojrivPuu2xCio2n8Cj9ui/g02
u21lL0xygWhzy9CLBkFUL8HZpaxLx6d+hqUIBa91u10HTWAvtzyB78VNgXP1hdwO
Wv1L0PxCTgyOsjMXBXspfUle1NQxJx0yTWM1MYebybW3mpfPxHsrS6Q6s8OuoJ0Y
THS4axKR/1TwTlcj+XZQXhAXtv6IMwyOTVvZ6Yg8jtbBz1wbpjpnbhjXHUHCOL9+
A4t9Zzp1mm3PkKSUsX9McCe3RstdqKqpAsfc9RAMADo5/T0Xdo0zL+ut6S/c9Tz/
oTz3Y+wgE4Ec01/pO518LJLReeERoW4qSCZ2ruaROHEKyyeX2Ol6bwEhyT3+pIUM
cTCp8XD3Z4FG8DYnbdRS0I/xs0F0hAUvc4HCvRJVTYeT6BQRnqrotaIRHlXY5vJO
RiEzckwWMx+UAq3ngtyAlibGAoiiHhi7+PGZGuqVb0mcYLhm+Y1xUtoyjBMF325S
y8eMyTRjfnNOGpTq4kbSN57+j/csyxQBi8MyDp2VesY8+TmwebdmE6f24q+nw3Cj
Et3qor6IbVkWfV5HGz773/ImWNSXnFKOkHeH6jcNxsqe6qCy9iNpJg5kPDA+cLHt
+glK3k+tnbkDga4InO0QoX6l/fWgIdPGdnRUadSxw00LvCJtKQXhzN6GjBelLIoZ
2FkKyxmcAMjn0x9lFI1K4WSgJBe5n3ujtk3VVI2t2iOFqzG7mf4BjA+3j9Fapuh1
jSq2RfdvBCjm4sWmq5jUBA2/wXyNC69rIbdD5aGnSpNnCqrjxZjaW9mCW0lOFC7u
q1zWZba1SsTdArGPM7Ecm7rJFkDZ9UiR5xOC64YgD55/tXDJ2Ygle3XbkpdxhTVq
gtoYoAe+d+XJQbjXF6e/HOeEzNVVS1PhMrj+qruG6iamDGKefSwtX1qXt1y/3y81
mAuVrj+pO51KI8opAOi+0eaOTkstARLyR9EcNmNwZie7ibR4C97jo4gajR9bz23k
IIA6RGLJJk534gQ2MMneBibWoNr20o4VjD17dvnytCGfp5cpkcdFIyctXThhfm4s
5OOj1sKCeB9z8LPUR/EnHChVrB2i3iw1SECmKvaq7I59URBrJmbLKgOMpkhOqkMZ
xToT3wtvgPwNt3CEVaP9lP8hgZc1NfFoUtbgrr5hszUgthVnoPRAxZ0pcIsad8WP
D+nvQJv9y9d/Ak2UQILH1vRpDC0YZo4MMCAoEfs9rrOAm8fDOnzFFW79KSUH2WdQ
q4eeWt1AQd2CFIzsSnoWQA9ulbPtWfCSb1tSDtRXAveNk5xH4Q0u1cColjjO9EGi
XasrhJY46hXP09256IZTSS/MlxPsKobcyobT2IeJXx35Q0+EvLS4QGxUnXNH+9d4
0S+5WZLTWndAtDT4F2Nx3mAVtxVxGJuxsrwP7r3lec72898g/zkQUbi2vzuWz3x9
wuUs6LEd4mkySUFa1qRfJnmEsig5hMPLGWTk4WquAzbd1vHHdZMWbyOByrt1zR82
Ebifu/zi+iJjCr9STm4rpKhw97xrLsoLtmjimac7Ny1kSoiTpcaiDycWUyO/2eF8
AiSPpKX/zN7AMKMIIO2jxsf+gvUotR3V7AOvCyww3ru6bO/BeroAUgSghGRk33eE
OQ0mn7xBaish1q6GC2iwW7wqfAu74ioNrsRR7aYTmvpiqVdebhQdOQVttxsn0fmR
UM5NoGkmkcbd5adZDmTnNpBcRm+6nFzNjarR1TWvlHWzwjnA2bI+T+qWYH7xbrCY
/960S18QLjdC9288fHXgKteb/Nb3WFhwdpN4UykLcaH9AOnX7bn2IWwwumzkM+A4
iV6ddz7x7hbdqp1RmMQBrWAQaApt/4oO9+3/2zouT74vaI25kD7T/52Ntb5o72v8
jVhy+E+3cKKnXvyyu9YT/VYep/2qe2sS3iOaXN803zn5Zsk+MCDXiTcZ6D+abQOp
YLOKqEs2yBQ1ZWbTzB9KKP8nU2DmSXUYOnr36K5mZPpL2CMCm88VYgnbt5CoCvCf
Yu5gqKwB0gNusuQ5xNprxwmeDVS+v3qn8xB5DGiEe2QTWWnK8b59wfHEf1EQEHpC
+tywZH4ZzNUq0xk6sVuKTyCMaSHsqGmVntCRzcbHCjpbGeMuPL2me4dDkIkkiUFW
HRsLlV1LifW/ZR+Wl8OW9MkAr4V0EVc9ZaV417//tppg65s4JoZfTvwhifbkANfa
uYF8Ajj8Lhij65+18atWdOpXiUvpf5VLAXHXs1YDfcHAPdIzwkljnACmjroo979g
LNVrqIzFl69WAx8ITQqC5QUY55DuoqT8tLX/Y2w5sbbeP0B2Bt9duYhVGXeFbR3Y
VffzRwNV6p/sFN+gQXsuItK6K6781Tu9/ZrwFrF2E6DUP4NWsOXHy7/TtFKNEIpt
6vulLyns+IO1VOBj4bbcuzUVYaaDpikJCbKDHKxDz2uCu1+c2UH0LQoDPA/VHtJy
7MRZNSSmdFgxyk+bn+adZ9PLG/K5cyskPyKhSpTt2PpO8Tyu0dlz+lqEr49EnkU+
H4uGq4ktS/UEcw8CHwTOiDkWmbCUbXUyeUSouo4ShtJD8tr0MYviwdq4DF4Ihwdo
AtP8QbEosZzVzwQMU7KXWie8oKByecggb63zZ9//ApJWvvnAZl5rRDspdE0u7kZ+
CZ7ePCbfJnQV5wZqXdg1QzFaVUkH6PAlKUkpa1h+11frHlN97f5qZjBAeULI65Bn
UUsNBeNKSg4aLEQTqQcSJDDUZVQgGWwcfzoazZcxhFThE8LrD+Tugid5Yo48TuVD
PqqpM4Y3ml+csVOSVSCtpm0yXBL/9N5zWk5iiZcREDAWPV9B60gxUgT3OydU3V/a
dxDbRQi7+miMoRmnY7d8of17cJtWLCDOo9blT7XVsdOG7caOv07xT2JaGOQJgJ1h
vwsSVkYzlUzNwlvQNeTNecy+/yi8/mYwUGu6LYfpHJ02ISigJJentfLBrg0XBgQ/
M/51J+15ue6bRSfdUMOJYfLlfPriuVMcdfUX2E9jqOzAW3NyG6MCp7GF5LUZwUo+
7rgVVVnckgLBGkqXcO8s2icQiddKELmmAY4IiS8wYraA+HtYKjKRykoozY1SjTq0
9a1nzS68Gc8PM6jqzTFcAYpUhl0/ibQL29AcKCJhyi14WzwHJE4CRiomuQqELUf+
+lDr5b7INSAibqO9QumQ1eUPBp+KN4YwurNSyQFZpW50mJfVU34cnYuV6DvJFDNg
EfBFEF527slcnP1Qqz0UyUb9pbxE1Cs5Uk4hppO3nNILguoqmJFCzoIWjBQLLqqy
zM1kelYsAG5HFMLAepwzLfq+542L3LvW3T2MQ2nj/Bv1XVtQx5JU5/5gqiBAuPph
25aZ1dkyNxgvcc040KurN/eAFsEHSL/z4EKBXouuYAG8o8MsJ5r6DgL12TFz5eD8
baOUb+gmUoxJMMyqamMAqTREDndl4TsHxj6jg1c9JS0HPWVQleiFf/qyh31GF30t
0meIIAlBADFXy1Tt1FDh3rMq81ukClulOYJdbtoQ0n0a+0k8DRztnc0v9NFJqhGB
imiYOVs/BclrUn0oPiYmq/3TOnl5nDZSuSpYfbqD+/6L1jeTYWalyjiX9L2D3E6P
885Xa8CSgK9IkQlLUC9Jbf0J177LCs5l5bhESw0oYF9reY54JGc0mejlHzi/nHmI
k3WTEhvsQn65lN+BEGmVFlcwjchulhBxaj5/HdvAOEku4kLCi4MLP2p1o7IWwi1E
vTKY7SWh5X5TooWfjs4qcqESRArU3v0P57X7Gs2UoFqTy3oVUdCBKxx8hQMWPh4y
GQ9tevzj5eB2bT7Wj9mh8tyO60MEkLA2S3E6jfCWJjjLunULIWALTmwFvvRo+Og7
3zlL25W1q1I+hNX3lyHZ5NLvx6RcP+v/5PirtG6pGx3itqfLerXmIkEGtxU2PMnc
T79SIvLUZRYFFAHJ1N8Oq8FQw5NjldN4z40ryETQ/fDfYcjX5x1HZvtmHzgPv3jG
hAsquHUh2qJThBoSpdgAQb3Qul82JXmEEHlSM2sqNR+3YogGcTUy3x6mVFEecu+n
9zekZDKSQzyuaEzbLx5P69Actw50QDQQfsW+ZorPcR559VmPLftXellFgK+Ffj4h
paxD7FcRfH8wTuF4PYg1riNUi1WBjX/M/fRSRy15xOGW1fIEeNKdHh9Jz1E36rt/
M31BsQe3ACxeN6FEbN/X2OkiPVudgAONHMqWknyyN/NTmQgxTPQTc7ZG76zgPvbU
46P5/8fZD4evLV5zuYOl6PDGZLkhpsEIr+MJsSyRqlOhg6/DI204IeQl/A2XcbFY
HGPfJGiFjJsLUeDEaHnJvoaWuMKFqYuuUw5f45qlEAgFA7hGngPELttse1/X+83j
dRMfdfXthJheeuvZ3cTK7NPIcS8BHXUBUjLPU8PLNKxGOhis+jbk2GPaZdYwMl+h
B52A/NbWi2jQiDTD79AkGEQlbfkAJ33DFR2JQCuc/E7rfDC33uJAhRjE5pHhMZ4+
wgAndpwH0gbrVbV4cZ/IpPLhcjtCwjde6pM7S0B8inRTLtPcJW/F4RKXHhdg1z2H
OFl4fuBjn2LUhj2ugwJBLjhvR55OGxJuHVdHNdNk4aeyZLZNNYowSIXdVuhwuDb/
UvUimHgKDQdmPFAS1Fk4HGYWohd0IK911yYiNROZ3iakT7cgGM/OAqke+Z7qL0NE
W7PdEHZ+kaUb448Avl97RDgyT+BjMIKoSziDQbAQ+2uctcD6+ppaHF5crqFCJQAd
5M5n7RH/cP76SEbWgGh0RmYWbSE5r3QflRMtT5XP+12CE60DSQgACG/qTNWMReHy
pRMfAcIk5KSWy1QNjBDYPj9nROntzbnq7830mo9pk3858Hn3fYR7YaenU1+hc82B
i4zYTa9UweEBW3C6iwlVzj93brXyCvzFK0DiI2l472VWu5VlkOcBPz0H/uX6I5mU
sqFYaZWoMQNLpRFG+zU6BH+vib9TlnzjsBpWZBkQFld/2S3JzkH/vY0xnqkM6nOl
syXVZnxPZElq6uwF4ivNXVg0qFYQbolfZ9mqNTyMq5Qcs8KIe45FWw5kMRtLQg7g
II2VYGnzNp/5tqWq0ATL63ALzlxCyCvVuBXk0Hpd7AkaPENI4pmQ6OATvCyYDCKV
1pgRJ7T5bYBDL19CVJuhA0txXbobgkI3xS22d06YdBMUidlZsfa4C9U9vDSDfymS
Hhx61nQBa9YpJFs8lf5Y4HPsJoxwhMF87m1v4X66thBqDfv/UF8kVQaf1XFTRp2k
UE395VOFx0W2zBqbB3svd2klNZi8uQHJpL1JjLVLX/TEWZ+8WO/M/MkBBVEOrfjm
6BstUyzt01FsXdWvOcMYwFB576oAak4agZuIKuJCIJXHuYzchnNB8IdqzDwAOJR4
hJM7aMY/t+UXvn4bKaZvWPJLxGm8flWrKAPcsReplph29B8htaA3I8UnAlgegTUE
5fTCeLq52PxhbKCWd+qaZqCi0lk8F89378qVssQtwyS5ep068fICBQUd9miMuqlE
YwYMt5b4/dh/++5MuGwoVZ0NyQkg1StzKKQy7uxOFYYNIDJxfNb0jw2dmG9Ayo5v
ioHZXl1olJdX8PPysT+RdFqP0XZg0t7o8R6WlBCQsz6ZwserAjV86+mzy74VI5Ck
YsnpeDowptv5m/Z9dUEuYNyAuy9sM48tPllnlB5PNeIj/N/3WV8XlGO+1/9OrSwj
kQQN1krvfxJU6DqtFsVJV+1lgU197ipkMSaShXH8cMfSqMh2ew0Uz6CT6/7TSJtA
PTcRwlNSaz94Zz8rneCXVKxj6pkvh8j6AWhlunFnjFPD2WgU4JyLojEIO+X8+uA4
f6XSqTW2F6DQhe2t+fdPjjYj+pVqNda7t9HfIa9ALlIZUCBCe1d/5mOZouuAidbz
8UxOvGytjqYs2cks1IO/GCtxL+jQZz890MAV1u8NiMqAXYLjBKfv+uC/yfZHPDfM
rRotsg541mQlfUQPH1Z8RONxSrFddmSQsp7WEA11/AzPGq7tCYHGMpjCj8T2AF0K
SeWCo88XYmbjU9Me8I9MNrNvsnHAR4T7m8ZjrMryUtkz9XOjnjJ8qT/4nrqBPB4X
FZIh45qfUyEnpP3Q00KSRWSDRpLO7mPvX7dFtEEidPFj3BKpkfOS9kBv/AVGJicZ
DgLSn5ee+NqfZmyROMhtjd6/dqQCn90K0OiEQ2U0oSE3On51kBOkd3/AvrXtVlH5
UkJUQhZ/+xUm7qe1FdXVyt1zo1S9HhVrEIlF2I1BR7ScxLMmADpVVrTTk2V4+1hD
8YDEVFaeviQIauqZ5uoxQdEyBJ6vi45MmMxU9O7lAnKplw9uGc72Nf5wO4pEuBS3
7SHvBH2s7KTmlwVK/orQTXZrbNJrIsuSHhBCT2yQG3Zuv2z9b66FnkN5dpIyTN0N
jKaGPqtx2H3ClQ1aXhGiNKeYb4srkI1o85tq/KMpQqh3D7qSqfjWf1PotOvG4X0h
lvXFjxqWzNQe+boB9is6XxX6ylMjPRaTHQTPJl4qkm7f2UFrwELWVDjsTwSgpGlI
mQCubNWaRo/n5jfymInzWtqkaAadFFI0quIjetbVB5B5/IT2wTjwaaoOflxlKYaJ
sVE1CsGokFk2W5xUsquRX4+SwBhQDDWTXFikj9kf44f0NG7NN/D2tFKzRnViVABn
V2vqr/OUhqMT76W8aUP5xgnlvQK5bN2QY2bz2FO3AaVTWiawEv0UUwya4BY1gF3K
BfnbzNqbZUAXdwdwLoUgVUefMOafCrvEKqgNBG+GmSqefnxdGXyq3UTPw9ryXk8S
/l23MmB8znnei1ikA8Okpz+x86l77CsJKNZYPDvXotJflgocGkblptMxDkSPS7yS
0S1LlY1PTI88nFz0UnVsmJTSQQ+sXq+NvjFcAB7wqOPVLffYN4/yGlmjBSqWZPBV
WVCy/v4cglA7P4HOOlsf8yvdGYNcllvSmVqOhyPmqxYRurJp/SyAe6Nj4ixGhQPd
kFBRjuABnek5XFtz5UtW7A92wvZKqC8VjLgoBDad/+RWYGn2FX1hv9BUc07ZKjE2
J7Pnnv7ZYl07GsvAH1AZ1lJI1TNE0EkDir99yirBVbarD1E8GRtqt6XBSZ1yTSMN
BTGyxojTVXnkyaNt3rsK2hj/vxaPt9yFfxRqKlxcq5Y=
`protect END_PROTECTED
