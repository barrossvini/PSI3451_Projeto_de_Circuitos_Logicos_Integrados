`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y3AIOie/Xgt2wwmGgcA0vrdrEgce2nJbEDb0/BiwyZJp6/3SH8G8twPBYcrf/Lg8
BROXaL704qewvk/qsnYSba9VE1d8r6z6FVb1UuApzHnPu1qfqZYNPalEE9m7iMPf
c/cZWrsQ3gIOkZL3k7ki0K8ynbEgRuCMtyj13UnbPTUi1DnfjBX4v/PXMeRqe3F5
HQmphHAwM7DMxbZJtAX5rUM5g7TOdFcEmjbh9KkL9YQ8Qi6Or5Ck0j0D2ZwEhuXd
hNjZU/Q5voChaQpgCIGzBPiZj2IOOJZFJ21Vx55BEiULsQJeC7sn496y41uxF3Rx
qZww0b0fplMvxrZzyZVLVLYbFIkxUf4xcaNrbmCtoGrsh3YINmctPzqS7xbtQ+MY
k3E3dzKtckzOZFLlq982ygEFTw/2/VqtdYGPhto0iZTL9P56qdZk2p4FsdSQlzQh
Io6cEGZR/U0iwACZJG1VfmTW11uLPGTxMo6OCi0H9209IlI8uPwNlQSgiWoZ/7q9
zG6IQ7wWPhKqteRq7GzKG4OXl3a2r0d7xyb4ghduyyXhmWpn01s1qlDE1/CKz7jr
BIY98BoSlByvzq++zz/zz1RYLADI48vaDNtMZK6ETe0pq4jsWUKeXjgiHeNm212J
JpFRIfPshxPKGlgWB6vcg8fZ7VwesRXtbMWlZsaqb2j2eNnUDjZ808MMVRSl/lC9
quiJT0ZvTMAiP4YsJCZhGi7y54T9WFJR1Xq2Rz+ug031oIkDaowoUq/LoYYGkKwT
06LXi615e9mlD1AaRa1aVv7+zGA1sJmrV6UyCaux55DaZ62O0btlSeoPPHvRXl5P
5qmQg/Dor3QiJQKUs92qyujVhpLIZ3lK2wzCqteFQS/N8lHt5bmFaS8ir9JMwmHy
OtwRUWC0Zc4WLOUBJsloeD/o9GNGkKJV4DmkPCzthZdPEdGCaaZJ/nZd+2fQ6QRv
JX240bhU89l5R/TAp9pxKSiv3kzATlQuwC0Q42F7oH166mn90621Xpr4PzvkQbGK
mXXD9EtpkjcqhPkp81EZNijyHpJ/p5wlRPMmGZKdob2H2cp43eThWpYYIMYzrGhX
odV+B3OQxwmRgtBLEcGDFztDX1kGbASlTQLFg4fmvVKqzpDsoo+5T7yVf+fwn2KG
YXpEFTxuSei/mlnOEybSCvbo+bM/gcRX36Bl27cHeGwpIiWDe12/x1LK/U3i+b/1
DA92rLlPXlhrgNXEZgITLJLut4oCopvqcMc73D608PGvsyqOILxGwurJINM08tKR
b4zSdYuF158zClotMscbaec1CLyeKNhIH5CbCN8G+DaTFdz7UpXiIKyNsP2jbtI1
mGQHI9iuHlBRw5uO2bhtls7w44H+mH2UsJd2iwzCZvE9LsRvVkq0eCXjWIXg6D2+
M/FiR6vQSH1I02oC0yDmzovSfntFUTxo8m6Y202UrSGlAtzZ7aInCQA07ydmWAUo
hS2qKzOInkRHYe58KjIhCUrut9BKEaENCLU8SegyeR18FXb4ayIC20+D61OWfxy1
qalD9FL1XJXZ+ZeleYS7Ltx6UfOzXNLWn2eq1wXT2VE/DrX6/d9mBf2mkSUL+Tn0
NWp3u72+LA2RpV2xd5OUdB81Z3t9cJirXvNG9oMYbTNaz3d1veiQ12S93HUEPM4z
KzLpFjPp7bgriKPepg6NqJEI1J2dbi85kR9dVJVkbaafLX6U6fMhONkGCZZwbaFE
0iimvO7h9GleVsk86TB5NanFFfqspGXUvuB2RqWXE72FWJUhYuUgrUJoXCnI4jlx
+8Cu0h0iQmwtKRrcCbZPBEkBF4fGZC/glV5LfJQ0osOU4la6ejXnNeIcrfQFIDZ6
aq433fQN46u9gMZdejSEOqbskMaO4Z4GFhtM/T6DBHCJfLoOEl8Zznd/YiU1OGO4
fkHV4Qz/f+DruNabMVD2PMoUAYTb0EJjYwPB/QYIhtEymkVmaUFhxFkWdHACgUjS
NtTrfKKEM420dVoALSekNqwWjSPEqzg+JmF8ADtyFgB7cBs0ddWh+hCE3bMSmKjS
ZruzIgW8tmhDyW4RhJT8YCE7lwLPP81l9N2vAMHgaMP+MthHTeCpDrby2MLCiFKz
MyUsPQJuadZG9NwP0n4qNaVdvVM1JUEcrBYGaXVuINF+xtcP0uv7xkCsGh+yD3WL
8vbhufzoHSnJd06Dez8g4Wr/JaOWmLrSJi7ZJ/Tk55GkJuCkfx6SoLIfFXJuH0vy
cP9OfvnMLbyEoM3XAEesK3JTb0zyKOqJ/nkXUpunqSx78MUNr6vFUmFhFYEO9+3m
Psb+dLY0VdwSDrWcwVGETqUE6+PJ41QvxXs649kwysOHn1PX9XV9J72i+eK4l10e
2OTGBuRITVRzMmamLLQJsq9Dno3bKuHZCad+nzVwHSCU/qEyG4XWVWylsVdJ9ue3
5BmR2GWoxKXVB8cEiPQOmT/M9TdLhk/yF1hU+o+7MDAIBtX89gX6TE4ymBAvspxl
dDwsL39YzC3UMYGXvLNeVuik3s7SZputnbBnSVefKUqRiCj2ZUI/ljOs+ff6KJ0L
kGtCnnU3tvNweWWg8WaEsqEkEN3ZAumtKmiPNxSySXjCazuRZrCoK5VK9HxEv+Gr
tST27FILYqqHGpgUYGPkk4ELacoPNicjHyNq29xLuOpybIEeVJcf686h3j/ftvU1
OYOdD1avrOu18kSZ3yv3f4PySeUC6grQkbebs1nQsNoPi3NQCuk5UJkoRe5IVX8j
IMNoyfugSdaWfeu44kxHkPQ/fqOK+DoV0ZXb0ogE0KMpTUl+Dn8t4TtoUrYLJTbY
/nNIYkbFaEHfjEJP8PlHcS3WOf09Z3arFIh7I0aUkAlQByrzg8IllwrBcs19mPp0
JHHRmUA+lwbXvHw1iGP+sfQp6gDKrtLTC0MDs/L9i/tXbz0jgjROZqtqQD2lcVU3
l7eDNLgVxqGi0hVXMVStbGC9dpISnRKlrZ5p6BYdc7AYEk6YylC1Lykj3Q1MMPF8
EFT0h1OcuTci4qkpcQdU7dX0kWpW4fvb9Aqh7sta8VPqy1inSaX4T1O3oqouO2Qh
jgVgim5Xyxz+pOD0/VcRkXb2+oDUgmSoCOAhZEosYN+nHMSzLZRlOjy9RLKhFbfy
tC4mO8UVBp49b+hoXBqxjkNr0+LgpLdJZvohuCLvjN/YaceedE+wZXK3wHb6aWjo
+ys5p4cosHFX2ERIMpBy+r+t2T1T9qfnDhxcM5N8NNknBptTPESrcc283svl51TN
8c5NvFBx+qnckxFaPJEUPewkcX+kwCVXm1+7uPQBXhT0sBqnGd8PhrpP9Alknc+h
6Y0of0jc/5apeVOMHFvA20FdlOkY1OTjqFWZiFyUj9tyEhmCXmIy0wdPL/W0F37W
62CQeKzEKoelJ+gKm2ewTusmNFWzoZ+2RD+my2LG0Ik5GCCY72praj/lORCqmzga
QrYqN0Y+tf4LXUwoUHjF6cTPn++sAZVHSafPS35DG5nq4irmj6KmswJ3yR2SFCFK
CtCqLoYV2mi/C3OYEkSxcVZS1Xato+bfzaTVeJ6jGAYNxB9KdXbt2c6G/u8koyN7
tl5Z4pAHJILh3LEcCTdBzBF1VWLDwz7HR1G93W+zg7gKVuy44oSEiNNFy04AsW9M
H82juMAtNOYBz6gJA4OANwQSU1j+HfYhiizf1I230o2dul19u8KuTM1ynh6we0Ri
W6NOOuBSJ8sYxPz0zOGrSp3RXqS9Juvrbtc3ecpfd/g35k4BD77hsu+ttQkdkx6Y
Vxnudag5iShihgV6s+eVI7l6EZ8TH4AyMIz3slIkNlyO4nBQanCdHzlECqENKYDx
w+RbGsGXDBbHyE3kVc04MC2gsUP4myWBDJL87YcUCAEM1w7we66Rx3L4StzZR4dD
1+uw2Yq86xVIc3Ay3rwKToe/HtTkKxbAZ6bWNmOZJt6B3QqvBQMzB9+e7QvVr7cf
SaZLQEb9RsNmRM8Dp+8tXlF6DMtvedWv+Z5suTYTi6bZB/ikfSOR0VvBKp7tMpUZ
nsbLLLHa8abzByJiHh2Rg24OsnmJqQTNGuZFtVRQ5ya26JbE+ucu9GSk6y3Cp4T8
wR9HaEZ51wBcuCWJgh/77lcSNL8j7OYw7+gnG+5jYVCtVCtcgmjl7/R9XzPf/svA
vK3a9fwUKJ2637ht8lNb3fZgf03Bb7gpVocf+HNCUEm2IhzTjCM+3gmZv7LRcTSZ
eetlGcNbQWPsuXNPHXgUKkl3buKPdXPfWTajN+p875gqn/X/j0RGNGyJGaadaIjm
S9QUxurtdBSw9Gaz5zK/whWMwlLq4hYnqwrC68HdNLnaMZT8Csv11wDbF7XR4A5g
qOgn3Gwa7DZkJbAzqhmK3mFyLCggVosTyDdtYjqUv/yfVEG+dyRi245J7ZezU7Za
/CrI7aG5TL6AQ2p7wBw02u3OoTZruRmDZox7hsokZeheOmn41GL8rrW7t7k9hF6+
C+uX4WXGCA8sCAUULltmVj8eF7iqYL7wA8ow+OS2g3ZuPkpCuPLxW6I49K2mi3jF
6t3UfGVYpIttz4JeRHMM+12eWogMA8QWX5R1UIQc44OTZHyynd0ef7Wu6F+LEzHV
oIfMphbPNa4EkrXRZxyLSRA3xf1AGyMYVhL4uh5Zrb5LNxskFp+J6tM/hclGLTC2
CeHJ0d0T+lhgiC8TE9UFqC5dFMEsMOowXas4ujUB/lSqHYA+1+DSE2IYRdmlPbau
USC3bAYGsxTtIbEPrVnnFtc1US5qgon52kpASsE4tiD04ToBRhR+kN35UbvIv8m8
fQqs8EAOgJe49GCK3U+qdfaMiexVWb9ujDamArBQQD6vMoobl8HMIsfllMtC2xe4
vWu4uL74xh9sIV/nk0/NXp2++RfXY3WgDh2NCmL2+t7CSDodwstO+g1zFr+U+Jve
sjEdrZOIfqHvPrE2FxPmzJZdb2svk4i4kh+ilhzrv/dJIXWcRQxGc10nPDpV8Ymz
BsSPu0J58fA/ShOFYTyjQH9ic05qibeMX5BY0ttVoJsxSrh/dS0gi0DqbTASPXTh
ChUXwoDmRQ+plIjuOvNgGVGrBvndsqSJ5dCFoMMwZ35eMycngRQNGh3xWd6YKNEm
VPgn5TEcp5hTHaVtAB14+cKaYviIVG3f1C8EeEc2Eqm2ACLB9jLKnI4/uA4KBrA/
TSjkrBHErbG/lATD11MqssgmTKtggK333bCZWkR+nN0b/R2aC+cFjROMs+OQkhlC
w3H8zXvhKzV61GyWSpxaKk+Fk0LAEAJzCSbAPB1RuQtU+nPQ2hLa95jQ5zXpCb60
yDIJegzpdt/N5K5QTbmWXkmMQdTIS4nmn1XwlC1/4DmmUHXClKsPTI6mjh87ZT3Y
psLxA8Eozyml1DDQIPOTlMfExerGCccWp/0Xub35HsHr3n6H/d/W7hTn9hx9jdSL
ZBt1xyuYH2T1O2Gpv5jO8w6bES7IWMI+sVHTS300xPq6bOgsiyk9pSDZlVzsxLHz
Z+q9fmUuLQTbiy+3A5Ow5lDBHDoqXK/XWxNRhhRfiAJrQ7dYVqvQufdgavjnYrdr
sCaC5nFBPw8/tWlrnC6Cn2B5W4S22CfBDZPijXRSNitaaSj28pq8IJroCPUBsyd6
axmk5ofghDrIB0VgNa+c+fsjmRNAStlqkgyjhZynJTpDj5UC18cwz6ks+lKu4w/1
dTYX30zTvarnpcGSaE3mVlNi8Tr+tIIRZZloxmdhxoEDgfAGFBMUuGeyh2A7Fxpn
lJ26PYPUliYCrK7DH1HeEj3pEhhhoRXS46q7halYt7HG0pTTVP/PONzrveKAFMe2
gZxl56kjBtGiUH2BPdk19Aubx0SplfHWEmUsTFikhfvymQZqnDyqezxi6XpqWp2O
0dILLaD3MaXnn03AWupOZUfd34bCdda5Xh2YUcT+b/RfCuQqTP7D6PAm1rp6jGXH
/llPpPpqtGtegBFC40Ui7iY85YnLdC8dy7VpLZOIyI8hOZ8IhxKLupK4gevOw/eQ
H5erj8BTuhB7yhLYvMKUe29O2AIAEU6F0aJNbyul/o8zdtmlhm3qfvwHG77KODkA
H/+6pG2Snfho5okHKaChoJzd+I4AORjRQWLXlj0LY4Vv1b00ukHspk897KvAAVKn
8YtgZqMnadwxPSLhdJCdItk/K4xvbWgtAPUiV87AT/sQPzzlnSE6ONwdzio93g5O
R83J9jWNZyj/7A4dFwFK0RtlKQfNsgJ8SKbOujxRByN1264w/Q4L/peQKM80toa3
By9IJAz6wItyERgZEjtEhqTsY5AWkEzE3plXk8jZ6QWAIlFxTXV9PmQV7+mFBz8o
yJtk5ypn71qX3C2Ghn3Z/NX3wLbHemBkZOdeptfYzdX1HCKTfY1SwHZS8Wglryf/
Pfb57f+XoOHfU4ezCWUUBPWeIFH7lir7FyzaB3Vqn4xuvzEperoHwjuuECghuyI6
wMwwJSegCCD5WJ6USv2D7NXqK9tD8pXJbHuy+60iEFxawCpZkxyVA+vBy7kPwEpN
i13jPZjz4171Tv9ezhVRBzZjfgkS+yoQyCp+AX4gwlScGxpsrZcQVVVTmlVjxFLO
T3gZhzO/9/EHpYyvsVkVPbkFtL6Vt1fMe0Lpwjgl9p4D99GpV7HSL4+sg3UBBvlr
2ZpdAc/ikMtcIp/mgF0zJGptmQEhIEm3A0dr+0k7Z3SCoVUJKpkvdpEWEpVAzZfU
kyeaXzoSv+mx0odqKYfmmER9aoL96QQQdu6joO2RQ9u5kvp2UpCsVKFNwDQKLLFX
aOpFPFFo5XZE7JaWHQAV4JyGKs1x4OmGIQba+lm8s//lDUXocppk33qZqBfLNgyD
/gfOLqr2X9IhzydS1aP7/kBavGxHvJbIYQJhGGF+nMKZS/dK7TeMLm4betFubXeG
cy799uuzSiF+sBIVTVoojcui2SvAUApV5SS++Pvhi1Vl42Taz4SqSd46VwJtNrf7
ReE3oKAfgzh2JAL2Tl7RS9lPWMh4Gb2MsAHPmbJQUzlbKLNdgVFMyG5HDPQ2q4Ae
P4LLMGJUQ5VUoQg1asmuz2CJlMY1LnUKagqZRHDlv+YyRH53KhQ1Jdrt0eK4389j
r3Pk9eeq6Ac9Lyx5kEeC9Sg9JAU0M/lNq6PV3r6K+FTCzhtlvs9BDy+xwhu2xOaV
QZwfBw5aVp+No8weVjBbKeX4+oYvcZheoHck8WwL2EMLpplWkuAePuZqEehGpgLj
JC1y7LDN2MHFPWDIpzY7IA++nLKw914HT0CDwc4NUZcOYVz9TTT3hWegySnlWUJP
rrH5A44sTQkVjYip4YKtlJZuiTxKWfBFVoqJWwUIWffSYenEVC0DFKu3zVAUs3BU
nLSNODrK9XBJyATk4q4ErregfmnOJvap0EvizhJee9KC/4hutu43bGtQOqKARleo
t6bjk8iqmF40qrMPbjjj4X9NeQ9Uo7MwQsgQ4DEoJLwVttt2Qp2LYvMtIXJodFEe
Cew3dVm4b4o3675kfRUkNebLgEEXRMId3bnKaMHyJGIO0hWD/zYZiX/cIdvm7cWW
I+QsDxZzG2CEdBYHPxR0Q9vWLJwByR1NhpTxL5S9+WEY5Xg0dknHVH1AAQ5RBbve
m/TioGF5C5hCMSLwjhMVbyBD8GEnkr8eGTmLkZBiQFsGKF5WlKUzxsifxdOFguQP
lwL1xzdM8uAt4wL93D551nzqhjG4tFUn7lrziNsPiQadczjwtLN+L8judD2f+cqq
/cUXYCKzehzDkWKGun0FasJjd7rbIg3pMQ7v3Vmpmy/FeMpWx2C7aR40zrpEkbUz
OV+cKw5cq3G5kzJ8yMcLr8IICXt3lcPaHNSU74+P0d3UTA57TRMYI77WbnbBwkL9
f/HtiAFfw1rhSm/XOS9NwU7ZsX4gAHoSVhgsJlPW57/eXqQUm/4RWkYE9HtMSBsY
LqsQ97cTnbmau01Nmz5X7m2xRj5AjlWn6ngZ9k+SqcW7VaGf7Gn3JCW4+NlSNJ/7
YNN6ITlvWNEJtUTPExRaBvL/SeB8cNGmj6cucGqT/gqLHhIhZOQ2hPqwpq1mihRv
UrfVcbw4oRkc2+DWna1c2UGfk+FHFhpdhHaRnCkGW/EopCLp+9P/iot6RoUTd0hN
vgWFfytJLrtrZHkXbeTWpSMNygslisHBcgi0DmIjiA5/APtiNa7AAlo/a9cBxBZv
Xs1q4b4texWXl6Eak3QEglmzbzzDzPNg3TJJHzV4fQ7rpQgb5M/9SWEfJxn9SpXo
Ui1a/ij6dCAWNVB++X37KzFUoErZE7dCCimAwIBaj93Wybw2KX8IHoNRuAxVCZ0g
geAjvOu3JR90jY4C0V/Qab6lNwVyEtFJqf0AeMwzE2hzRP8loIpNWy3uEoDHS5WF
5RdnhG/Wo7rABZ8o9fIWp1npChC8P4eBj7VH3/LTldc05lLRReHRViA3AR0a5XuC
I/i3ZISyEfpcfGePDsaBVX6fcG9c11u8M2WfrB1ha2WJsVLnOtuuIMWYVE7UblDi
jBP2a4yA0z7DJPQvyr+nMSPmsSdIOHRMXvfFMzQaMeMeWzgM+WpmCaM+BHtux89+
YGzGU9rDkKqE79pZ6MvYWZmOXztBnkxKL/6cJHafYRV+btjzdyNHRWog8MLrwBCn
9oSJZHmp4yacIhSXaK9SkjbC3cy9TGQtuNoP43/Yxiln9a3+e2wbWTI4FX7au0kn
ugvx6dH16z4EFKW4ri7Rz7tPTCFbSHoGZXeCnSu9rpT104G9DTmckhdSw7L57f7S
0ktMCR7pmAOT7qJnFTv2UXqyHf92cwpgSUMcZxr8KWXLhey5MAnWU+jQUPtd4b83
pCRbP2ZyU1+pC4G2xbXG03bRodlaHyFBfake1iqmGwsqMamUYtLn1okYd8jRqP9r
V1tiDKYO8sKbx2Q/sZJDKJZlLGlULnHLyqYwjAvLWebL17TFDljo+WYIwoC3nqiH
u96eTNM1YU4qpyv322uOI+lozrwS3SNdSQXhMHVgRLkze5FEicjEAah4AxPZwS7n
djJZuxJTU7Ci8jv+1y1/ZYveh4ZYoCPqQapxw4Pn7vL7n0j3sXSDASNPvjv7EtzK
DrNWS0LZc95LKiL/61lk/sR5hBFMMR44GHQNic6prCanrlF/WC3uDNdvl5iuWwSP
JGR/zQhyxi/Lb6Xlrv0HXuLzwXk22USZclgcuA4mWEE3vZv54A1tVFOzMPhbhYpm
JMnOcJCEuC/vmNrQk534jrR1Gd8TTP/wYjRlRbvz+gG17gsNKg+8pqvX/ivUOp5I
GoA5UhsHj7VDctm8ln6oLphSdK5RtJywkdJ6duIdimF/dhgv9P+c03KeOXkmLIUP
/4l0QCzdV/JzwRgbhBQNrpPhwsDHY5A1bFrHzNx43VZEheV7ThuuGaIQQeaVCLI5
JJQrMaH+Fdip32LHcTZOlCxz9DyA9YZewvT6aQoLQToxiMHLf1AFzgiHVuTThbvH
gPo3PzIqeeYfQ8zR0ZhngdNd1pUdZsZMi0JIQqP587H1h8d4zxhIu3XqCNlACz6O
oP73nq8vG9NP/74Q2TIs3wnFA9BfW6JoC/9uNG5SSBGPCFjw+VdRmsiaDPC+UzbQ
yEkX/Tr9/E47qB8hlgBUyQAU6ZK4exhFr8nY+BCmudu6zgzQWGHaEmmADDkcpss2
wbD5CMEEzRSBMosfU3spWAQfzog6FZroJIZbDpZ37he0Ila5T9ULCXLHeCQ2/6Ma
87b/tG56LDytdRq2OwyWQngMzobdtTnrovWQqvoba3hdPE1ZdHEuTqUUq2y43nZd
jT/mvXvTeuMqqEizTA3TkOfPKRogEYIla8b85e9YvXVDX2tOSMFIqCdAlOwfLAUg
biUs6CNzDJTEeHGzkAC0eoj8OrxTsMmQeOTNcYlh3e+zhwiMksuGdOLWJF70Dci1
+OJsImx94WlmHOJk8BXZteU9IjGZwReO94RAmeEc3ezodHdMaq7h5iWKHVqtbMrr
vjaPoCtjiZu7rBDqtMlZ2iGEI/WZfHPodFj7njj2DfEtHm5/BuEijdNKJU6j8o+Y
BDNlCxSLNxtO2szp979AyN6Wee2mCkJPYSrP9JYO9hANZmKp19XHTQwOEWG/RDLu
GMyZySN+hsaL9LYSMlluouyPYvzZS5BgeTGiT+6RsOGXPFnjwD9RMx+oKswnK1Nl
ixzim0f5SaBmj3KojfzhrZ3OjktqL1+6sOYJu/RsKSf7DRjN6r4ZqVI8gXgU62lc
SbeIAc9AWPpZzsolbm/at1lCFPWBuaF81Yklg8o7CKubQ5zAcLn+U2WaVEe/E4FD
97/pOJhrk1Xc4Bsw+21QCQELupasXJeOoIeGwxdrTQQh0XT19Cdh+VdIb2uC77Qt
lodzCzy0VhPSpHozx/+2tBcN46SEBiV0s6S1JAnvHzjkuKcVjh0+zMFv+s9EuMQD
anp4jjdzfLP76brXEi6ZtKkyyGCGd3jRZZMRx7K6NfGUu3Ln81V6jjf6/2dhH6Qo
oji3NMVJYZDMFu9bRgOO7MFH05b99PdfvGBhnWvpUJiROU7jrSJIQ6aLZFDucDom
IPVoIk/MWxAe9vDU/2a8Ywn/T1rK9e6yokcymUs6a/ZnoN/1MzA/Cjm+OUwP8SpR
ouEeWjYwKhWOn7572ZW+dciZ3YrS9X4Pqos7YiLaqKxnRxKjuKoWvMK1+CKE4r1m
YiJMDHBGrH6W+dd8XJYa9t8jP+IALl2pX6BDUGhD2/huxiWMqUdwSsv56RBl00CX
MciMoFf+DNe47JCpVbqe5A4oso/Oh39R3Jmhfk3v2wAjyzSbEAldj/hzyZyE9WMQ
ScZpx58azJJmBmBfheq6F4ouRgzbTdHVbjR8gITV4fHVvnTH/cMR5r56Pesn9+uo
+CbZMnftPOhevOhzPCt2sLb4H1Y+I6/b3Zxu0V42tyQ=
`protect END_PROTECTED
