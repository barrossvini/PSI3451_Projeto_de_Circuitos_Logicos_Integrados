`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kABP8wQLtu4DEt6UvFsWS2bkgrQQnVoTywAzTs3HlMQ5IAGYquD61qtHmTxGaL5v
UcINtVeNhnt3/brFSogy4Lo7jQQJfsQEG1Ft6yZJzNBZmU0f9bx7xTjV+Hrjr58j
vvz1G2U2BTQDAakSA/rP+kF3otruuP164ppt5qr7dsFKeLgLHYgUqc6/JNMBr8M7
1oKZOq/7gP3IHqc8w8bQWl2m5sIEiV0JM+33OXPOZAzvBNNqmxExIkpPGv/lD0ho
49M5qikuvhWKe44rKWyNx4969VCzwcjRDWpzqbs3KhwYEHgC/8m/QMP7KqjeQW9G
bZ7dYB/dBPv/N0t3ym5p8ABzp6OCNPAMnXNW/0/JczqwtFw+6vA4sSlVOApO5aSw
8QxvtNAXq23e6NdQGyu1oI41hTVA9sIVQsmqHiOqAh4IRwkKYaVPF5mhAIjVvfw4
BwLoMPltw9U8MVVaiqLRODROyF5OJVVv9F1Ky4jm0tipWm9VoZPjqm1t9aoR76Q9
NRGx+bg+wxJuNci68u9eVQoYymkDiqp1AIpb+sO0dvVMHFWqPfPhMvUpTyhgkFRv
dtLsbRW5L0iMEeAtwIc/2Sm9Gg6tIW1/psYvT8q6w4ra2kWSX5pWrRGVO/rnMA5q
O5+IEj9meTD/scR5z7QxDi3t0BC4vugUqoGKWFmkghCMbOHWWu4njQE0JNaxcmDO
LQzr0y1hzvjteiSnOrr1NioZekHSTERtj6ryuiubdDyxZOQ+E3BdnBauzL2YBXNU
5/0wy3xhKEaJGfdwYYzZh+Jgb19wO9WX4aYhGGKqgRYLzfJIPqxUurjbUFq5dbcb
DbcqXT4tePfc2oa9kyRD3LM7MdDVb1OnDsVfbLIAtmG3WxmdTsY475BTBxZ2PLwq
PauJNsSpUfTz14HN6V2xjSouZC6kEl3lVOif4zxv/9Q0TR7tFQagsIjoUO6s8S8I
CLNr2CGmEAVtypjlwcJnNkBzM3AKS++uRZ2kpakcUR05F1wWkDSL8S+C5DlVZr9b
Quv4FebS9EvAwenYry5mxd2twrspB6VSWLjNngpsSBwrRx/vPsvzWi0T4+7szvEd
pVkizcnPNnIAkJFk2vaODuPDcW8mk2Kq0o6IpR0Ws6ne/ZmJ6Gqn4SqEKAJJXaH+
ifSR7NgiTI92O3QJJ2BDhWPikITxbLjsbZwPefVCn1wi6qUbRp/FFXSpUYsaSzDY
kMDyuoOub9aJXCGO6gBJ041KDYyVdO2RyIwj733ipuv0vLkRhzPNpWJMVCrHyNPd
jwYV/xweHa+/d5X7yoQSjh4VOOMPpbqWHBOGZTG3jqclWOWA9ekLiqjII1jI17Az
MfT5z10i9J+AxZEPn3HKFIxRR1+wDIKBBx+bj+rAF7MCFEqcuS4qrqaPt0i2YIxQ
QiurhazOJD1N3ZeLnPFkdgSh9+zHgyPCdwUPnl7N9rhvtVHo3RU77G0XQiziteui
UIyoxV3eIQCAsRVsKIzDKA0hzpiqkcA/FNdn7cV0omM+nlKRlGwXHEGXLGoqdKc6
Kxs0mKYhkRif3nhXVqybxHKcuUg0gv0Z/SzRlQmDCbSxrKEy/+/UT/wa8sPOaEUQ
aEnxumhTSUBxboy02dqGRaZA6te5l41G3zlWn/FfU8e2U0Ux1sSHoJPECaW4ZGaJ
0bjgDPIVaYcqEK187N74QfiUUAEFFzI8hlr2SLMfwMS4eoiR3m3Qu69QgVT7EnKo
sNlZBq6GJ0nKfVAcXzRypmnxsBtBH96PsU7hARvjAowWMR19JUOmu1qMu5jH5X3q
I4e043DpsmvUpjrGBsRZzPXNkgo3orN+ug1WY/OZ7LzhJO+N1G9R5/7r8oe5bdnf
l2TevY1qwg1pwlcoKAKRJz6fR7Y1QWzTj/MAwvGM74ywd6BUujL+m18vcwGjTJlT
KaLZSotcAVV1p2f/3xh7wpWu42X+DX+4VBOtDKetxH7HMN4IXg+tI2HDBh++u8dx
D/20RtztlDkuhIBpc8cet9Vh2vt35ylhJ3C1vT36mo3dCnF73OmmS6Z7AD+EEk6Q
mzPt8DV1DJFg4BPPEb1LAjnnyGRXzp+hBFamkNYtMFzDqgEYlBHPz+Eh30c+T5E7
QnR6rAkXxoa0okTvToHBsZLtIbdAn/gTPLDOKM9ta/SgXXq7pShIWv3Z+LZd/1qk
rvjIIlkM94Byt2eZAzFohA7cAVoTFtENmn3s6kS7LOLoRS98M/O0KMdiLvK0O2fD
MZMaUASLtq2Lv7no//5rvAbtQF8x3dHtOAvLUUGOcXPQiyr18eMZ4IkTGZarKcgZ
8FlGKdWRIvKFJPsAOPXlEnipFdSy4GZTvQTyqWKPAjkVSlXT/V1KhsgwRPqo06iO
ApHFSmuJzJ7pj7RrsX0cgUNd1U8CTZwrR+2w2ptuXlFJHDOjQByvbs3M4RF2LGRQ
owPpV/QOtv/E2t+5M6GKAon/I+/zT636E8GomZaELOKLi0AMaz5egyXMZEP5ErYF
JnaW3E3NfMSHrJAl5YcJGmyjxFSpeIQ57rtZ1I8wDRGLD5o7SHMWmCEeylNhg9AM
AADmqbB2BlryvyxDum9rdyvwBaILYWaatL9QFW3iXQpLTBR97i96zthp98mSwlOo
lQXTU0el46v3R8p2cAbO6BPRxzAtzYDiJu1w6WzDsQg5gILabIcF09SlQw4lHcOq
tf2zl1whUPEF1zKj3QWbLzxGI1Z5maTXZQvhAyaWq72aJfy7e8iW8EIgOTairFqr
agDZPl6iJL61hbVvEgJ66pZKDfMbhJ89k8+cdQgdLNh2PZ6gaHA0tRC7ViBLRQZq
4IBbd33z9OP+KhGS075sSyEIDHiKeHjqyjyINmiSmvGZ/YBe+3w5F0zX3OCCyOds
7GKVgrYQIACGL4An9WeagM3OgT2J/F806CYYc9xEbmHJbrtUCLgwV2z0CTKjY/S0
P0KPACYCkF0dlIIagojJ452rR+WuVk3TBmmESDB2M2oKUeNlIJMA9cdcAK2uwOlb
7Z5jsUr8hU1AXybPzDyelP9k1tQ+AYN2SqFEG4U9Df1tgVmsWKn27F9dscZylBfR
YAlKRm4Z4cXE50EmTAmy9s+oAhkFv4qUDOWZNdJ1svtfQCS6ScIlR/6bQvchfZb8
7Lp5S5UeBGixptTOTlkwN0gTFCC3e52vTYmhWA4lO01vPVOmJ8+WI3ZQLc/EaxfF
eDkr5vGR+tflH9ZqcD3EPyPpfBi49k9JaaF5ib/BYyWgUnz4FyA9Wy7BeQriCbGE
/SkYYhN7asWtg9IEjFhI852IrJA+JvugTE0KNHR0peCRykkLxXqPbMmhKsFzoVlM
bHb9/rlgQ7EHGUImn9qyiq5lT/YhWeVe7kwsnYw1ktmceNM79Bjo6AfrHZvNrflK
vbTSwN1hU4Iicgx6Iq3Ae9/Euw/FcIZ9hjJBNpuY0Ut+1m2THcCnei3yBg4BNF3l
e1FIYLNPvHk7TCF/Rw9tKpmQrbEvThC+79KerZiO6vtZ6507TvqAffzRNHvCiXei
jKoLE2wjUT8lNtw9PKO0Sa/oDVFYbrKHmV+jfJ8EOwWwrVJwgx5mXOEWL4UutJot
iIMzjchTy78F8WEbPepxvh6G4AWHxxziUd9KeUKgQqcBrkmMA51pNWPiJU/31v/W
+jFRIR9mvZpjUWK8icnPMoNLH8lIe2sqshbGu8GaCVQo82xRdGaMylldwHknVY2w
XHXsMolJP9Xu33TekxV1yzD+KLp0t6iQORwWXQAb5QyQ55nhXLsbxG5LpNjpuokJ
2g90CMMkVEHfFaw7b7yLQf+VjTnppUCcmNpYUZ7OtreJuDVoGeVjWSEfgBjfeeGw
P7iZFQ1yDblUAEtg7tJKfJmGq1FXm27yqiAWLCeiVNMxV61RFtq/0O+Pw8yEQZ5Z
6uJfSZfSpOFmxjRIh/I40fBX16xYAxTd5u1+Z+96FSzFylo7iaaF5Wo80od44jla
QHDtLU2FYqI9YxWt88FGzNtPh43PQfxbPDhSVDvO3jHPwhgTHGVoKdynkl2+yR7Z
Lrqz1PylV5MXc65tyDQ+BwPdVHOgwgw6pbDmuyPdzFzFGlj3kE6gkOFIu7FANn3a
KFKfanTEiePoN1xF07WwaUFLnAZzCWkKzf8hGTdse0+Suq7ETkNve0Jx+g0ndtnZ
YwpkVxRaHlLsE7qQOSAw/30jZLW32TPt/zuZa1Bec18AhvoummGtouUJzR7DFIUE
z0O0LN2xmsoRvKTHouya/8brTzIBL2jtemRc3Z1vbDKHKksVJ40DVPpx3XgvCpIV
3lfCAzX4+QhZgDS4fAS7Upa9Rgdxw/le9Z0ojVaM3X+TtHanVMSVoTlTC+qGW6Bt
nRwPgCQ7SYtTC706+WWZ3GA4BwO892tOgMwrqDYM7mcazZ2TXbH8yJbvoLKu4LDy
gsT9yQ0hhhB4kB5AmRU2SRRSsY2aScsHoVTgiaqbod1XzOHASaq1s2AhGh2ddOzp
+39ZtAZAtIntPo/eUuQ6GvybKMnpdaXegZfAcQXlXuiwZM9BAPCAWS06O1ARAijO
op0H/xdDN4m/GjUoOoaab5gU4iZC2h2qt5cjRgLOsWyItAaPoHUAY5Me+rqZpyDn
AYhwFGo7PhFnbXHnZgq1lPNSxdxSG/lQNskri0+xvxS7xSyRVaBO0ywaIVQLX5Df
8JBGxOlgUOFJJ1YFXZr3BNEN8sy1dlu+EqxB/adhCbbMrO2wv6Yc5za5yFkO+wrW
+TNA4LOMcdCo2OVLvbpY46JFzaXpx8TnHUn3U3jXMhmtJKPhPryLESI5Kp2IU/H5
GDmoNno8EXprY/nEo21aPD739nv4kJGPxHw+/F/2QvdHyZud/kkGv7NxHh5UWRIk
/W6AKT+FYasOsIt8UFygpigcS897WQZx4I7B/tkDbz1q9X2P2soamymb0HM1rJ0i
KOn/1GE79HlGNpJRIVgcV6eKSNTFtKPp3mvuY1SsZ6g/DMTI5WY4ISb2oJanyA6i
4H7FbCsrQ4DkbD+1uq0ixuytudR5kKv4qqZwGweBcItu0mdXBkxdNcZqDwEJ5/dg
0vcl7KZWLAtDzSFn+nGsjDSN+VEYB1jP0t+9b1aEAV6DNzBE/mQhuNKbzK3YTtJt
KXyQqoPANfgnhjWc5gU4NDQhjJNAuuUMwrp1OvnkadPrsL3b/18ZEjVq66NOKp4Y
Q6/NL3iZ+Bwze/G0AlHER+7CF2Xkz+oIUBS2OLS2R+/I7pAaGTeEk4ITHIEV2QV+
9juAlL3Lm1X8+ny5TymAvFX6qH7IKJTkRIiGV0fmXGOZWVy8lef6mQbfYDptT62Z
QHemQHitheqmctalxyDBY4p6uDusrg1fnCq2iVdrhdT4itB7A4q7lKBOHheibADY
UhJeipvGAoYoD0dEdhTCcl/3IxzuO1z9jjmg3d//2vSD8aPogWVVMZQUToxD52B6
SJOV7Sf+krmrdo8sX5PdIbxNHBLMlrc2cMZ3c2gPU3Miww/p33aaJF6dsgHle2IF
EDT889ZyOn0xpW1kxo4MHO3V/mU7I/P3aArjOPIs2n3yHby8ibncpl5qUo1LXFvl
P3XfBk3kxYM5ob2pd2kaGaT08WobKR4lhsmGXF93Gb0eE+/POKxI/LXyARFOCdgy
N/lQNPWVK8d/uLn4mx5GpEoEONa4xpmOpAR3PK/YpOeo7FsK1afYU8Ll9R6TIz2m
+rzkQEhi4gdi4kWmiA87qiTfQpj/V6NJU5qZIWWVLJAhX9mY5pwSvBDCbCdZpjNi
7sGt99GvD4FJq8sWdF+PuzgYPy7gF7rzWBpHLe1LYPakZ2rjujlj5byzfwJFId5S
YTrw+wLPyMRa6X3ub3xZ7h6FliBavqK5eiAhB4qc+JrwLyJqZjiy9MVpdgzoMDE0
6UzRHMUZalEdF+ipP9s/+k/H5vICOO2zUEDtkovHcMHCfdb+QPprRBHEu1gmdR1Z
69lculwr/tHGbRho88DZlhB7qDauc014ZIkoNXht8GghChsMiVqc0DJLrMhjzLe8
ASD2PpRQ+RxMiHmzXCEju0QEL9a9xFki6cl7QoEkBBEYt7vn0X2sCXFpTM1tvym9
E23yLMB7ejYcYvYTqQSrEOm0QBhTsiAJNhrPGtij6Q78IotDymR9lOfJqrwf76Hr
mydvw+XsGBfDkEe/4ReM5Kllj7zMS8zXwpgFaj06mciO0QYqduSapndezR+G5Iii
ortsAXCbO66h3806BDQaR43Cne/HK29HCeQNLAwGE0VNd+VYWYloW4LVDaM+lqOp
2ItALIap+3xyt68pSTNE57X58MjPEO7N2QiPgaZr3iVNbu5wCTfeH7NgXZMf8d8C
XXJmTDDem5sLCRWxq7JrFDulC9RZkcf9skLWC9CEVofdHT1PYXpbW7SUEQ/7D8ue
N1C84gle1u1qoOkomG2JPn8OvVkLZwA3sSyOc3Pz9X4drlKSWfOfH0wnIDpIMdIm
nA1ZgcrICMu2qoh4L1MMuEcy/TDH14kUaI/Xjitz5CjC/necXrg5ZnrEsl7G24e3
K/jmCcy0OYSA7clvmL6ifO+r3CpWHGLWknWQ+3BDgrlhFfrSV8GBqc0nJWo/Elo7
0ZrnF2n71MmwWT86vaPE4rq/JQfBwgtul8iY2o7nKO3GBJWGh9lZptwSAMp6xmWM
hcbE+KSCXY7gkwwsndcCBhgChLpLUnz/rfifg6ekKsAflkeZkeTkOh2BjSPVtc1I
s50EZlxhyl0fD47B8Qkrmsy8DG8yyOWJY/Q+io5qjS1mBndilvCG7qGDDGS3l4sP
SycaAtmAetHoE6+i8pnobiqf4pPTqcXeYZW5lNyWn4stW4Yy9r3kUs1PsSrfvWAR
R0/bF27h6ovdWDVM7UqRkQ0K1S5Eu9h9VvnQC6qbOYZ+GlLLrth2/vMpCsVImDOj
EXWy2R4Pnbwt5AojbKfM1zmI5+Y9EJVER3pMysTVtMmlnQKIJ+TA3XWUBiExksBZ
1jR4YhmujzChq28ueHQHufcwMEs9VBOpvDyXZQK6/xWGsruigPU+jh8l+3rwRz29
BvRvCm7BQv/to2Y2IGZqHYLekYRDmLmez7j9AZkwWMt7FnEh02Mady1LTZSybHhL
UAceXYxKQCzExVZKLZW3sX4jSixu9EANLrT/Jg5Sp5g1Zt8Evo4MDlapnAu/YSag
uygjvKRZyXGwZKRAz2W4Nrzd75oKbNqVPmFPofLoL08kH8ISD3LWTnLrGMXACaIS
g0h0BTO19nykg+vj740IGjiUHPKPO5C1U0k306yBWO9GGar5ZhGIUCsoF5S7Q9AM
PyL+yXmBnHd1JlhuxQmgH3TfFVwRvlSg1eBy4SmeK9AVcpCGQB2W6ASRbIGF1Rxs
sasWIpNtQGf8em+V1jHYC5+ZBmt9Kk4CeUxXkZBI63OrisybTk3j+r9bXH1iwWlQ
ZKd38EiZ2vMo5f7eDfXk89KhpOI6AlX0NGcJrnZCz6Wd7xH76GIT0Rp1vGwRs0Tl
pJmBqotGWY5b0FGWhY4DQ74E9hDxXGr6IZOvNWhk45yV6TWcG41zQ/AiJNpnTZZe
XYH+WcwikWNaqPr864G/o4uwanrQGQAjZgxYTzgMEWSHd9oIMQn9n4J884f1mGKm
XQqYTmNSEsWoE9OfPARrUYDD74CLlVRUPtOvRFruxvnzZ1Ng76n9w/NXQ8tS0K8H
QM1L3EF/PkMyFha4T0n9sgzpl4FtZdMUkcW+igegP7JIDAJ4zxqVogt+Zm/tmtxG
6BGQpxIBMDup1jsyYAiSZxEu/y9nkzMQMN6bquYM+6KKUsCy2rAqoSOo7WqFDN0d
OjJKIeVARxR7zseeRp4khs6QlPVevXKorcyfCGxpGEaLboJ8v19i512PEXl+c5dk
tOQr90GSrtCnLH6dyZTW1snj9qoB6/DZ0T9du3CPO+mvOlsFvkD5VSsTCJwLyFWF
97g/4+q6QlC136bsEbxvfhU5DC0vR4Ruz5AWG0tZL13kU86UHsRSbucU0rpLV07p
lZedy/edJ+7rnfporE+uulAcvke8Ceujo+Ckq1VGnqXGac9s7H03V/6YymCpKkhh
LUua3td3Cl8caCSbORUgB04PNqbHHRWm51pZSg3osxwoe+ThGSYCmrpj/QtNhkUr
9GFH6Sv1pXfOggCFyeuVYvgl+ndwIMllViHQL87Nfhu3PMczk98Zt1h/k3CATigJ
tF7gVz/ez3CuWQflNIIWjjbyAA+44YfkArZN3U+QuNGQkd4RU1QDWWvSAFZe9e+0
ioNdpvC7eU1bAMdxvCDULXV/YrSHR8+plvHvRMqJ1v4V946bi67Yomyoq0VIFx44
f/A8kIP4IRrjqvefN0gqX2vDl512OdjZKd90UazwIHV4D/7mCJeDPtg7kGTWRLba
0ZAH4CtNBPBS6W/ugwfy/DGs9BF8p74QWhYKD3pLeMU/SFmADxNJOfHpJ2XsVdC0
DCoMJwbv+JTQt9ei77ziB9azFgs8zepGR2NIAbuYUSxC4343BekJ5GoWwMZXRj59
9TIbD6MaGOLbRdZ94/27EJb63+2V8fWfNoBbCwqyDieUjKHhzTphsi469hxgTtuK
EOPAW5ghqPpCCHwOW7LUke3No3flSFMnJfxAA7ay1qrIDGUFnUmY7TC/gRSmuNog
TsAFgtGriUJIMQmxT+5IxlqAyX1lG7IHnewrM3eODoy7lvkpGnWqfVpV/cV8YU7S
d2H13nS7q3HxfNokPNv3pXzx+T1+AfV8AhCoSyonJ2dY3/4IDlKFybzwnzsajuLC
6PXcs84KWqbSTCynDXBWDyxv2pKVHPMX2RdmBh0+Z+i9hfOinXoWdJNtsBjESESg
neYnaz9WXIlkIE5pO6UeuyprTRUPT7adrswOWSX2y2MJ6ALP46thpS8zP2oh+GT5
aFQWwbGssodRbknP3cK8SYAFN2zt/hOudyJ97Zdq1B488M34FirUhaKR381G9PDh
ZEsbJXv7NjWZTIa0LrkNRV9jL8ppE5a31s2Pn+j5yZef6NCyGuY6EV1g9PuZaIxN
f2Q9I40ZkE9cz/UNxvEbNNQG487W/Q4OlOsjz5cA16u8UCHuuQ38UoZtAVZsXuL5
9JCGsd3/FaMvCWTY87y/alz3vdQEcZKLlN7zKEqPgVtHGGAmTXdZjL32cwDoCmW0
skjX72h3J//KEBiv1c0nBquOi/E1LkMzIe8mZzg1BvuVVnxCnzvnqcE7dCGkaNyn
C+CHVfo9XqSB1nFN5ms+xpHhh/AwRD4HczM9fQGojA81qrk/P92CBNM3PT621P2S
LNBVkka5WgghUeJarQzO0KD4l6UCjaJ3FWN0gMbmEO3lqVyhSXppUWGYPa9hz2fM
xsejKYaV3Sq6hQ2/S+SnUBbevCSo3o4t97vKVUV291lrA9AjNXuxrX8X/WA4YM9i
FX9bZ1v+pXsnwczsem1uhy0YCTqLTx+ZmUTolq0le2kRHAz951E8xsLhq96sjf4Y
rEwibcQA8SoSqQ40RBN2tnj8h2N3wQBZGHLnQuousUcAWNe7jQP+N8a+TRAc/c8D
MJt8Od5K7YSASxTheX4TJEG3H8HiQW9G0caFlv/TZOC0A/MtfxLWthIM85EvmPIh
nKLdulK//aNrzvju7bcyKMLLuKkElUN0vmEiSq/VVP0iKDHvCYa2AhAFsxS9oRRU
JIBYvzzvE13h97agjPZWURcx/+4fR3b+IpHwwDVhWM3Md4v3de8nVQy3mF7oiZlR
VLixUfreMYs+/+ISicJKOjY8RSLRixoe2AMjrIgYrqwMABKOfAQdfDruQvbNNjEt
1LkUz0xpIPKn6xzbDdN7otUWo6ZxpXLYeMH6/RU+gXBMB/UQMQsnVtU4JdopDTM9
POU+GqOydjPN8QC55RM704Rf/p9pNRPpaC0O6leW7oJpwUPYOBNKwGFZ7Xg9jGsW
zWB+NXbHfBV9RfVSQQJPxIxWVGA92t/RPfzpNOHsyQ+dBt4PZO8Hhkt6in2akVT/
72IaNx5bFGVXgtelGAMuYTzekSgRXLX1+yKSY0YqVbHMRNVsbETQh4TUFqStQpMR
AhMsibujVSxXL3OiXrCYP8S8EDyfjHiiQmFSvERVOQHsUjwU9/5hHoeeqEx0aQu1
FiWa0cXNHdUHY9n9QoL47OKr9mBreJrDcoHLDdoONWY535tvu9iFAiBgTpkr9p78
lXU9/lbUVxjbkeLqL0+2GiCDOFJWl1Kn7P7mumGUV84J51HsWPSfICCuz/pGro3o
6upt7kh9RyvEgJuos85DbwJihebTSp4T1a0RfDRFJmbxaz58vQwvZqpdr+n3BoOD
8XaT34GlyCK0gPlNC4Yvd3wxJq4qETse8haY5ah66VEs8HKFpdMwWkZDJWVe56Aj
T5LjGOsUzKl9QzVdkxBNU8FrdBK9ILUOv63EgJ5cHNxUx6jcehvK1qlDb+ewrnqM
yh+m+Y7JM4Jp0Z5XY8xbowFvThjlcAQTtsZC7U5w2xnHqeapKb8hxF595igg9Jcr
gJZgHknQQc/XT62l/MAMOzXo4fNeeM9CX8FqfiBE8eZPmDQb7CGsLvtxe7EfNv9g
r3YrbNmWsQfnEVBmAXZDnDSr3rCPrlznNcgaAhf7tghnZ3fi4Fm2dTTQ4Ew+tp3l
9W/NEFmy77shPHne+P14CJ4oAb7Az3SZpa5B5lN/Q4HrzN/b5AzcZTLLu4yqqCwa
jBGYLjNj+14CbkhU9VJ9EUgxJHpPB2+SnUH62WMPE+JzSzzq6tccLIz2fcaJqQ6u
KFCAFgiLzrYs3BQYokKlI/uhFrBJ2OXpglGVMMjB4W+wn84ujrNUAre2Fz3il875
zlsCHD5q0BeU4x2fLNeRAnkCihUCGrjtwCvBsVTG3yOIjnlBizFj08USMI16l0EV
untp77v9FyzZ+QTby/IrO/tASiMxJEAQskiAyIBZf8Q95vHHjUxjy4ikMARLs1ay
pnE2C0zY0EEeGg7x2hgmOgntnRmPb2uCfDIiN6AonNRW8brTrEFsaMu0Y7DNSN6R
8fiRXDeAr0gysn3iYhhfed3DwjVasIsNvR/ui2V8jO9JqR+qxgLnesXI9IfpvDyf
Q7uh4iVWWwRD2GFv5ZjHXEWqHuyje6Vxgn5SH9fZw9EJyB+ssA5FCU5RYTJZAs4K
zaerjTAqAMi8Liot+mDpMKOnWb0VR7j6v4PpkQBXkjs6Pcbf1VF6L/E+qegEFZ8a
W/d3CH/hQqdz4AvAxtWWyNi71TNrg1NbrFA3ccVPxakD7ONjpFTK9YVoB8dz4k73
rm6GVtNdJ+GN+FIOpQTF9JBidHrMvr5mSIrJ45FqVhMKHUXsDgVqC+BcoX+n3Tlw
0fWbw45BoAz4rmjLVLlt6gT3EM36/+zyDTRYUVN1skOz6iXgQkjhiLLqAe2xZw7Q
frkNt+UObR5HZfdVjjbNMtRUGKRHylKoK1D4go+S0hdyTknN1OVEMXc8SBbWK1ho
IgvhqfgXO+fnIgN4NDjNtzrJdkexo8vJZHGR+f1cM+GNCVto6whEjaNutQtt7itV
mosL91Q+8RAyv78P28vFh8kmXkoWf5Crbutjgtdiyj2a5NEvpsxEs2KX4H6R0TJB
HLmgsj7/smbLCxPcD8RaeM/whsamgSCp8HRbhrWgcbBHFhQucfD0nM9p5sln6HId
4bDfhgx8TkoAELSwxpsmm9a99KSJkuMciW35g/0NkOnlzpI16D00nGQSaTi/UGJ2
z5uYVpmocBPA3w+FF/3dh+8nff4YZ4SetqfqZQICzkPa74ul79d72jLhpjZ0w8Fg
QNX7QvmrHoZpvC0mOW7HfzR92hhz44hL9k3L4+LsWbjqCjsdqAI4L+sRTHVJ3Y5+
YrmGTMDmy5B46C58soIU0jefdy0ihjExftodUPazta5pX+eVFNZtMPlS73bgp0kY
iI0icOS2u9UyR9/IVmrZ2h2piPNE+DKKGssOkbaZwIOI4ckJDPWzotbQVxDLvSAz
g2NcRQvvGgqF8fwO3TBl2tHgOA7/D1sfmXLkUpejUgSFewKF1aS880vgHZkEIs0P
rH7zK7ILZDt+FVCVNht87A8LElzDb899VODX0PgGfp/U23FwT7l49iNelmqAd1u7
4/5uB0kFplEVEnYYCrnsbq9v4L9Y/5qUVdZ1BNuOO/XdG3eVsaarOJ4aw5Q5VTvi
Xml8UpZM+/14kGHejmhIbpk7WauM/pkU77DzASSaOqr6q1j4M5hUyhUMQiRV3EJP
vu0MaQ3svb8En6Q+DrJQZszKW0xmqYxR54bMiGce5h4E/Td7g1BFyHFYBsyCaUAO
5sif9kUOwszP2q5+f2TxtoGWGadOyIP5buL3ujp5Ge3TWQELVW4sv3d11BYAgH4J
4tCIYYLbELNIt/dtWcvwyW1v/aCh8FhCVY6JSgZ2Dl4HtkyLOwPgWtId74HWrTCq
v7wgc88YX3RxSJVYwRLjj8UzdnqBiiG3ydpxrt6GAoK9FqQdvYcYoJtrYxIRqhR0
RZg9q9VhP01NcSFeqOLA8lIGWPfn5v06KHiOddQwH9zwLwaFMZVF+dBeMthIvCoz
XAMvuBxqkbt69PKzT9WKj2BLSc0dBv/JBzJlymkC6K+sHE3HnWG/9chVoh+DTG15
fPvAaNzrctdV7fFWdwYYDhe/3XN/HByLXGfA/1SDgYGv1eSIETc3x5Qged4HOEVa
wnkiDSLd8EJTq0AiIb7cW0MfL05wHTRECKxHQ+ma3omyvODj8B/RSR70IqMYXFIl
sjz4PHwgjCiioPO4Gto0Ej9Cw3rrBYCrtyY2n3lgM/ZYsWvQNqV9cv8uIiEOMyVQ
QV8jv9cy6uGDREp4i8F0K2HMENyP0Br++NUP9D5UamjWmWTxPEjMczXcn2Pwe2Ee
Vh3SxNlxKf9DlNZg+3PDSD6F+tK7SwtchtR7hQ/KOUV6a0SENSsuCT2zkfDO14ei
r3dQRLpvpuG7qQnYOXnlM//q8wz4dPKYeo/fC6MWnTup8u1kUWQ4m1MUezk65Rf8
Wmxwnsn8USwLpt5yKNloY2r6APVDoOSKxLFvEZj0jF2HrV4pJ49JQyceWN21RBp9
xq6zLtupgkmKricBVYNGF4CDys4sjQ5Syzo2PPTlryA40aIz85JLDDIdcFGNgbzg
eiFi645taes+OeQQdUWMN9Hn+hK2rgROQcEFCeSc5vhJFLRuqQ9rSZjjSYxfeLBb
3EU96N1WrI7p3vq2qh/xJJUnl3qWrXWj4Y5b6n/vOxJaPu2T+GoC8o4PTekJOj8B
mKMv2X9fb/CX4vf+nq3Q8Qr2BwavVkdUvQ15zuD7Sk9Vvwaf6T6drsI3bC4fZzZi
e7KRPh/WTKiIOEvdRXT3D7Qjx1Gv0vuLtvFa527rkUE6W7Q90/F7Eu8SNergbq3G
ojTti4+qMvQoHQ3dglWudC21H/IQ+zL6LUERYUkuSiO8CGEmylWwIUfG/U4g6pfK
F1JuXbUxgl17H8pBMXbdGg+YbTZV02vFTxuG12eIUOZ7DDMSMPU6rx4CfN1G4vwu
3UWmFfgky9tXQgTNtHSxxmrHBHgVNXO9BIwFf6QHVDqkAyf/XN5AIcqs/kYAfn2r
a+N6HPk0bV5QjXU2TnkhhvCNXQq6XAxEFiMctfAo17SqP8lM1wbN8OUlrpN1yOfQ
o/PmmqUMpxTluOgbqiaQdpfPdDR+tOLrdDvlQv7ifri47iryEBxRfFdEPZyQElha
dN7FXxSRIuCCvgOfZtTLR+lzOPuW6DKKB5JgPc/QLIp7+AGdhRxKpSngixMEBlmG
s2Gk4L6wupDSbWNySp5kjeoU/j1L9bDBtSSM1KEfTKnEnPVCfkrpKmk9I0PfoE9L
DhN2vVKxvvNiJ1VTu/DM1XpXpoMw/0gdM4XrHZl91VFEvrUplFH3/Wgzdw0GKQiV
c8MO+iDaBKzOAeKRgbCpQMDVT4zKAwEYQvES4pVk1BrJUAZReKJaeLtUepqmsJVc
mfdh4lsGfbQMwkfkwxe1W7Fa5kZjt2DoQyAqlvfoqja/aEfQpintX5PsMCKR1h+c
xNe+WYUPa/iwPVUGn6Z7YKq0B9Y4PGrqtoY6wRuPSkOv/ADT3pb18+2UvpdEhz6X
ErLPPX7vTvUTplJn8caNjBFrGbmc1PfEc5f4jcZrqouj2RNrkgsvv2onFfQDzSzM
A6vOHdNJ1g4FKH48rTe82nQWodI2jt3JeHu9PKy+RYUU1tXDarwxzap70YH7FYrO
pZC9cm556t1qIZSkg0MIKpCr1yWYHMcb51rArrTg8gu8WLklN+EX3NZWrw52u8Ah
Sj6yHew4otDoCr4i3F9pUjw6v8yFHMmwpwDYpS9e9VwKtMuHQ0+SiUAW+ULRaVC9
Bp6r6M7zRdyiiDF2uZN6rHI4SOouzYeXmcfAA0o8UCDC5Q3i9KRz00I/fRLgt+jm
F6tEZMXTOhx7FaWxYUy3KHTDW7jT8UhKsN0s2qwRfcJXkzrFkTpPhBqvNIPBkh3Y
qySVDWUkUGTAa8BtIH5mL+4mv0YRPHj5yVVINxECSL7DGuq7hpz4Mtg0oZQuwooB
t9vwHDQGP1efjyJ75fgIbMIwMIn+UPw2tDoLYlyreR2UvTLstETwwoFnP0ZtnZp7
ah3UDj0RKqeo/jMJ7x9I1BeqBt21pQqxZssO2HCiEJMZ0lQ6z5XdEpgmlMVqpS7B
JRmIQVjgfQLjAhjStpazSQ8bDY1V6dJXMHVo6kSl3F/KgWmdGj1eG+T7fSQpLRL6
ZmJOkTCnl6fI88GJPGfR/gnUecLDQ+f5JMeWqa969X6Ntaaq7I/pDY1OoF7US1Xo
ZvKcuNRwI1oeWVNBNzRfM1QDIxkvs9Dbn8SLIa960ce93YliNYgg5+iT+KDjpwWC
z8ER+HevLeRQpOn0g7I+nZEZY7N5WemtKZ2tJkbnjl8xRKM7sV5/juLylsMJkioQ
pfxjMEKDaWZjCDPiiliTcyrawPRrufq6NQxV4mAEE0o6eB0PA/hIohbtMAiltu20
IBqDM/ae/33Vc/kHTIJq0V5H79WDACYmmWI7GeeIPfmfcwNar4mCgEhaAu+chcva
LyoVbCTbHunICRB4ZS/LvOoXvNkS4kl4avwcyALU7a53VklMBKjfcOoJEdbnRguq
RSXqqMF6bP1VN3X+6FHf5Lb/fJ/A6fj4Mkc7NxwUEFbkYBcGp5rf/g4pjodJGaah
Vm9qCR+hcmcuOjAqu4viD9PC/n8fZ3AfO2jVK2AOkkhedlO/Jd306cV3QEOw8Fbw
6m11wvMYTtYsb+IFd49lVkrCb3BmXzU+G+FuD+iqbcAznsfsYrA5fWDtanPIVgmp
iEG+5gxM1WirYo4rN6hZNlHdXc0DtJcVq6vYUmM701GIWNQ66bCqlgIrEKmn7AEd
+B0cplwU990RroWCQQH8ZB3IM1lO5/0BBFRNdxdeW/aV1PtUGY1MxN6gKKcPGkXV
/2o7Dqxnky6Y+186iU4Y/NTRHk0kJRFW5BhasUgwhy5iuR2tnV/FJRWIDxW7mZif
CT/UngBuP7wcEcqUw8H26SKEW69YMtnd68OwfoyadYKNjOKHcYnyTQpAI27C+Ddc
4yNwGEbOYw+XMJrDfsDr28wZRzCJQT8ijP8ndQSsswXAYgM5beN7heSkO8NAil0G
D/ELZiiWXMjgFU3LisVM364LJeiV/qya/38kbeiaDzhfTinBbE2cZQhloefGdneQ
Ye4bLYDijyCnpLSSqKRpZ+VHDVxrIECh1CRycmxi0Psx/+1OIVlrMkuDU4HEV2A5
q0bz+vz7CDl+raHGMWOjo5W46KWJCTDYBCw06QgWFxB04OLA3Qm33DbXo4s4eFSI
hsE4pc1zszEvTa0SeYJQH2EU++enbQ+i5w9Vw3ZoPbvOc8gG9x0fNbhBtkd3XTu2
c8VGNCmXkQD5Mv0DVG5VyLUchBztqJdV1C18exfRgvjgBSjQvoLxKkRVPqA1XUKi
GcXptXosFRyqlnmIB9zkipXEsYASHwaCnMzZVCucCKE4c3HPTrSX80B6Oed20WUf
6wXEtGTMYIXy6L9zkyNOAjXr3GGdNLZtY7/8Jxkx1siJas7CpfDZPQYl8VuZ0l71
Hc/M7EmcE2YNQtJIGK6CDtx3mK0lN0CvZV8vws5DJJ5eccAv40+Wd2r6cL96J7V5
R/73GXFolJjenz/BUeiqdvQn9TN/F8AZaPzr3mMGTYo8d13urGM0hY4MxBCcvrNc
fN+8+wMEl0QDA1nGxC0TYuXiLv9rabz6ILAtP7yDamFZkkb8vzFYuwDOgFaN0wOC
4eoxEMXOG8Pmc3226DZBhf14k1jCU4HUF7WEH+nieaDpsavvyPXwZ42+qu9PBYTc
h7fpR9r87UV3VGtnKyOAmRfdPK5FXwZC3KnW54m2B2vUi5ghZTQUted390YqzLcL
82XGrg2zW6a8LK320R0K8Nk+Go/5z0HAbRRpEAHvmkKnJwWTECQ5UzeUDaa0e082
VkA2YYAIgzVZQYT3yDpVHZwTRcj4j3r8PV3E9D34dG1Hg7a34tgUnOLVD32R78gS
TXOR1ZS53DJXMeEBE9F8jVY1WAgptMMrHsFQWQZK03gX912NUDFPLBMU91pBQzYe
19G96ihoDbQis8zFCC0V6R+yAy4uqe+mdr1GIVMog0vqTSK8+XzDF3gPgkjV1AS5
YDAiQR3zYCVV6rZgaHteL4gufTeQOICI3Qv8hwsJmKsNcXvmn7GNj55T/LPPe8eu
F7Lo/OQNjlo2waIOsT5IhsVp1z5DSgNkZBRFGykJlRFQc48yzaHj8jzF1Z52qqtr
ZMcZEDs75Pf8PJ2BDDpRc8vqsWQbyrPM7VuH8+cVCu4i9vTW3YVxHbOGZ8MycJ+l
TA4PXz/vUiQVcgMnSoHn533+UVbTn9HLIJeqtYBP9LWoNo5Xi8BB0a6fTCXwhgM/
rcP+2Q9mV5CR/ThV1yA4ulcv21LacziIzu7WU4m6o7xytCFDbXov/tQcxri8hG5d
F6gAKsTds43A11+s6nmVKvdmvn+H9EBH1+wkfxpUzw3J5VdN+nZsWQCQ6VH/D4ko
Y6ckJdoqfY58jFSVWYQArsGuZ1qicHyGWPBQMxazYDCmqjdUtJhqzShk/f/m8DY3
84OB5V3k1y80iuyxZSu7OZPAacYzrSti+oShP6FRpnvn6foGU42qS8j0FExBIIQF
FHcUi9+VzSyyoIT+l2cXJEozP5nE5AnWfqOQMk1/vwUqc7BuxwB6SpF4zfO2uNxr
gQez72OlPhOqBS9nvvlKfdAjJVvLcjLdf96IuVp/l8/v2FkVpQWPKjCMXKggMJ+6
zP5s93gOmL/FRn15xtukSRL+DPtfYG+KtO9sFcCKJQut5TFCyyz5CddA55lT7erO
akrSQ72fkmb70Dfk4XPPL1Y7bhyeUBq686jjlYr+N5m0Cr5Ht5rqK5KE83/HAZ1X
Bb+8BL0zbxYQzUEYYEeBfj8MO1k9MIIXkOjq9YCBYd2z/XK/b7j/PHUvDxQqiRm5
ZMYeGnBjendK45FmFMIQCleSCW/ih+GCd+XdgrEcVnr4AjsrCFBC3aImO9Bs6M8S
7pvreGf7eFkOBDs0nrJ+uuOJ217FHSizpMGRh59J7UkfVjlWw4yDifr4ChRC0afK
xJajHsKh4GL3tQ1eMRI9+7Z5S5vnX+98nLoUj/ww8afHLQys0g/ewNPRhid3QlSK
46ZsaHRLeEQBC1nc4EAIRfSRiW5n454dETWSGlzpJjqJx9spwXiWG/uvL9IKOxFH
ykpmHfTXvhqvrUWiqsyLvQLVzx4HM08CP2w2Ra1JErCZsZHj1lkNLDMJOqrr+lIW
Jw7WaLLvi1dkHRKYuFvwBRYwYSgiVh4Ug9rdOZIOuupdzgIJ1Xsr3wdpemMPKy6U
Yx6TMpFuWcbqCf8s6yOsi/BrEhT3QRcYI+Kh0c94gaSmEo14H7xzOr7mUeEz96VR
d+q7YCxtI4V+uwbfnJejks5mp43MJemtuEnD5YtJ/PGIEJmuGvkR5JKivA3Kh1H0
eW33koOApaKoAic0u+dQ9xh7ZsVtXdir+fUS5cZxm3VeoyGKi/UbSCg6oU6khzYN
RFjZ/8uI+LguOEaCgdThytqCRxK84TOZuCW5k3UGkYdehSQRVmNWH2W7//0HIOML
qlW3se+hamR9fh8hJV3HygU2xanSrX9uOb8S0cn/sZkO05IdRXmhLBscQjc3M/A4
Dl+oDHu/Ba8uequwBaOqXpwzYF1GFALjcTUMCxAKYcoeZtAj6uio4CYfO2ouas6M
Txzr9xN1uBYaoZK2+1gdILMi7WiBOue+fvQhosz+yMtSW5DdF9L0Gzq6KLCICiwl
99PCablZLPJLIuichHyG1kVeSNs4UzDOL4B1Rqz9tvCkbM2VQez8dRkZj/z3bJRH
fmzyQZJBWEogzzfIt+mWl0ztId/mI5ae4g+TFoKt8z9Jt9M8mC7GW9+D+JQmV1j2
BCWFe4knjrsI/yThhWX4+kx7fwCgtm5RTrjbkraLF2B4XagBwRCp2auNGnjhnCmU
ch6loMdqWw/R/KJjBe0ULU2R9+6FWQnSm3w97vKIg3bEiCzHd2zZty2L254CUFcE
LU2IA2HjitQ+/fLDNBI9HgYOx9jvG9TQRq2l9j10JxZq74kVGz1WuADxBg6nZ2Rt
fYGiq3lK3XYlKdzXrXezXhARqpMh6G4Ujs25Dqj5xmlEIeZgtG8ch+ajz9wW6WPy
LTaCVCAloWjzpAUMao2ReKEJgWfTu37802e4LSGw3VACNwp+ekwJDvmVuq5rpXht
DnKTfOMQylyfuCY/wdEFMtJiOpQUXVHm6OAOF/p7YhTGutN/v1vbIxH3uEW2OBuu
qcnX24GQvsV8F4GXwf6OOmxRQK/T9khxF034dPQg8NI2O4Fgj77lCZYhPLe1X+V5
3FnlAK8uphnymlSPZ/jguzNAsvM0S4hK7v7JLpq0w2GO3/FsX3684kVVhHyPMJtA
Ou9jFZq1p6VFlyNSmKCzkPGiYHMuhkqYMuYiR0avWedm9Ucet5d0muby6qG9nrYO
HZacG8+bOx14OJR7xT3IxOWwsBE2i6UUmEvFj80HxhPKMQ8t5Uz1mU7AEaT+y7rr
WZ6pfTUT3mND5nsV4W+4VS0VXL4qVybc+JSQgOEXPpZXYcfGARXt2BGbtGqTIlIR
3hokbfyntLJFxPQ4grBJnT7kiJr7Hk0t3KLv7CbnN40yWFt4XWFjvUmeIGZZuRfQ
b6cHV6dEggT0USisXyGxbuXF0v6NmyxkdGBf7vcLv/EtoNAYK6FEs0Ti91Wmqfnu
GytajxsKV4wLWHz1RKXy5dCCYJ+f2TMR9Q/YkLGR8IjuBzFTtz35zmRJkn9D1n4H
zwVgna5Rlz+g5uOoibuiuPHJybLs59NoHgTmdo/ghc/sWpamG+T+54AnSWLwQcFl
akfAI3dJNetWzF6KuYuOMrCC5YVaquZ2c+6t6n8HjsDCUq/aETLTAYY/lpKYhbHP
LVzcJrx7F3xfEzW0srtjtzsSNruE4RUC+Wk8cB5+DfsJfWKLT8z0xIKDmJv5F0p7
evFQ61w2Jg98Yf9zkDe1kYt6Y8ftOLOt65c5ugiuI77ShhoL8H5vCsXZgFD2uc2K
m/4ayw8i39+wdH+0wBFXBiefg/MB0xOwGNKN8vrna8hphVpWVrq+qCwkWvqL4/Yk
qRJtVGOfiasEanVle9H07ZjwYT8d5lKKbyup7GGgO/srADCe3DgiYBqKosmRUhlJ
LyNpFVXrEyZUS7Z2XSLk2W+nto8CRXDU2fzIAXrTyuk5pqILWa2PFkB4CgMIaj5K
FuSTw1DEm5e3G96NgyfzfmCAeT8Z7hdwVFPHYNwKfQrULngwAOGyIMmgZEI0MquC
Fu3Udhsz2IUTIzGoV5PE0no+McyEqy7gTsAmRHkNGQFp26KuC0nnEDM0V8fFPLUZ
mgC35dpnXirr+85P1drp/7USs4JqNSjhnhU1MOQiDh8EGc4vEN80IRElmsWQdpp4
1q7ZO3zoJNSMwo0VZRvRW2i1zPJmSq5WVOGSf9Ib3aEj57+XokKibOQ3HH8MYMX2
gOxe7OKObDvPVDTXXEZyDGDFnvEg5K7jNSWWSQRiJpBrwpEiEHhFKs5dVHKelqEm
r/dqyRGxf1OTwBN7StmqnRSjoy0hKJteFXlQsa+hEzHo2QQeoE+38WDE06kbJoQF
dliZmb3qzMKOkmhcJxYHo9krVyNihoy0IBr3Sd27T6FOSzZ0gw2q58uHaylTYMl0
KY/tIxOvztVbHaCyXL9mclBlLkIuQvCQKiITgla1JnoqC1oi8KgRcXmfczYjVC5N
tu2UOGRBFG1T0oB3Md7g7u/d0qUlnfaOqd+1JTKFogK+aXkq1pCyYi/uwucgI09U
Ey/5L2hvUWyy3eJnPFon+KAn22wIrFd+hhvekl9aZLDXAyiEuI+X0lxnTMzbBWDE
mFvAq8WrRvbbq3UwSE8kRYwnn/UnVrj0xuX6gyyosrVjZ77t2zcA6DT6rXFr1+VX
gTlqlXWb70zcDk4FoxV6VNX49IXya4BjpTk6k/LZ1d8UMvEa9R2xc8/rQuyLCv2a
zCSxmMgGa3vCe9jO8G/lVCdpDoykN9kORPklaNxUC3t88Oqp+EAis+EKLgtJdjps
2Ii2rNSKbhCFl2kfVhGc4XGyL/7ByX6dtZwjNEs3D6+hiVfD6k6xVM/I8vVo1uuc
B7QWDmega7Pf2X9BDu7WD0ovZIhmt38QfxBxnqA+h917zHs9dfMwK0PSq4Vt7AZY
Jsp9v0X8r3gi6K1GfI8TQguVIkJsYq4KBE9Wq8MgfzyDCTdY5Cu9JIVf5/qtQI+2
970ukld+d2hPHkC5eFbfooWVlx8Pfgk54b5JaPcGYawMg0mO9HKIjnc8/1wUur82
Obkff7vVkbmcr3BUQY3ks1h8c1X/kQKbol6dwZa8T/H1kiqSubQmJhz/50FMEqKY
CCdm8Rhk2kEoBoOhk5WQH9tDbVL/Xas72be+fbQYIIwt/QPu/SJfZAoMRfVt7tcp
TU1ZA7GTFC7nKFku8w6MJTyJ5P15UkzLVEajmE3d8bKhLZ3e+PFWnP+7kMrGMM07
JDN7MX0fpX+N8p+FHmn8YfvCswK0ukrr4bNZPIGsKfK64oAaPAFCxND3pBpSof4Z
z/vxSY9Yn2bIwOXOSCa4+tB5r+sKBjHjaPiUA3cAM5UB4OJJsfq9xnM2fNOSiz75
DtfMW8lIurO4kAPfcSfMgwatSEkknVYdpcl9gn1co0R8KScqMyt0/xg77T3KLGCf
99bMluIm5LKu7oySXhwn8JrQstarilwwB/6AeClEOdxtQDBjlv2QZ7PYopuxnTBv
PWjs+xcpJnZGnAGVjYRQyvyGPfcgPJNvd62WrX/WEWDC5GnzJ2yezMguE7jjYguz
2ETGCJhbauYdFeyIlsmt3q5pKLp1k1+/okj3AeZlwO28Fty5/njmrujYo07VOcW8
rR3EOXQ5+uwuR9AMhL2GeNnf9M9BIf4yfYBPBQre0eyhnxg4aqi9JrdKPAMQWcKs
hvvj1aphQJ0JUxhIAQMIzFVyWvLPXucSgmodt3xlbBgw9JE5BRc5tN9qCa9K82kb
z2fmM9j8RCpdthE7zWdO+QOnzLMfWostGlzmU+4faBxm0rQQ6SQm4iGr4JK9J4Y9
1bs+kn5dIqPRKgHPXR2nsGuGiTNRtYJJv9TqJHaXXra/3+wuC1JZqrp5tAIjgGI8
6SWJ/60NYqWn6yw0c6aH9NQUAxrGpBTW7anDRIzSlt0XVoS6IlalgJYPdsmPxm8K
9EnnAiG1S4y2zICey1ptnBxoQsLwwIZ4detq3R7SVU4ODRev1liW2/KtniTbkGyt
fyVmq+6+al6wv0WTff4jiXTkmG6PixnANSW7Wjo4wxR8mQarisgQ4+W97ar9cWm7
p+/j4566ettgIkEGUtTsSoudN4hVo/s5Gq+CzcT7wWuOeECPbsYFqOpsEbBu9Khm
WH8afJZDTqSPTVk9QaY2R47fRRJkqZOMMk8hde9Lc6Id7zZsozzo5H3ay0H6WBGY
dIA4OxBEka6gbYOszIx9sKdZ6ICA4ZsiMHYWoKeB8jcPiEZYNMOUM3anEYmAY0YW
sS/IotxM8MNmRyYYA7mgTV+F4n6dHrlFSd9GbAfcnujkr8an+a8DjH59oK0uvC/U
XHxLGEE/SrTYMVqBFQdH72KZk35yXD4Swe9flOIDrB1T8UVO9lwmF/BOhXQlrzpA
JIWkxkcZutcK7ziBkHGvcLJlRK9B5sLRGQARKp2ciNuYt8re9IhezLPOSZF7a0SR
kJYF1SlPS438DvYmvK08ICu2n/65wGMWFre4OkWepQLaS3QLmOZSMyINFWUiHRsa
fet8i1VKdPuAooH7zJnKwoT9dwvo9N9pYrPjg5SUFVE8qVnQJGY1w5k7Lyl4T3AH
xE9GKm2eYMiJHeIJISzsIdsr6DeVaNMqrvvGTqaz775uEsd90eWElyP0kKkaQtw3
onVttr6prUKAciK5qdh7YmjKQTcplo6n+Ri20EDq2MnUeO0lrb3j6tLSPJ4anVzn
1u4leAC+oNQlE4vAep0NxtEjii20UsU4HtEE8U+Noq/k+hpGFuq4kPdOhdtlB3vz
kBzj+56o9Ey0H3JsFIvF+nGN0NhrqBai2siv67pkRR4bmWYDr+CmZdoKN5KHzz5f
hRBDz+i1syc7DVSI3WpoxXWv6L1NInousjnDryawHdyHKyGhm0lcEV/WqfulVYC9
qgCfpSuoLhKn52VKzwMnlbAqFRV2Hqo+5NFygqMM/My8mp/QrAk/6PsWxHcOvgve
I8hshUlvAfsX+B4acBE/R9Sbb5sdso+ZlTuOjCnA6tBo5MEyHaeys4OLK58MlUpf
wNOTwjys6hP+NUP5kHcL9z4ff8Hyf0Ipo22VGot87O2RWcDwcygbL+asrHklSpK0
uW8HuIh0/5/qDBf+DPHyYhTXh/ojlRJ9ndAL1B2hHsakcXTakdm3MNA+ybD/obsR
yAaAdDK4P8NqWc4zb+LHTojElZadb/juAFu+dYLvvjYb8IpDNLBw1SaAUomoSDyY
NJvXmtzqst9BvDHkyopzqhBzLWzVEEuS5E7Nx8As9P6Osa3a/UXAPnWeUOseDGMa
HmM+zfNskAw/6TP1pQv0PjIYtRd4YhSpm5MpqGqQRB+FKTuiwql53DPc08WuzC8J
hy84oYUf4tB+aormufk+bQpbtEAkYpbkX39/PDcB7oF4cWUkaJ8ImQIeN+rvXz8W
BkXQOE+HwsBP3/O4kOSOlp6xXzJhqkMVhs7iikYPUo4wz5c49lb0Z2ZrawNdzPRN
Z6I5tXViYjFcDZZkF8tY972+ESxWjS11rl3VfizLxQzsF3gw5CownnHoQib26g4V
U0bAU2jBblRRceCpzF5LAT+QWZ2R2Ayov8vvvo3Xz2usmruRY65DJ68GzliuNwoP
qki1MAcL0R6Wsfal7LERhnvC0ceHw9BowK0VYv353+PRXcPxCMJz4FnVkhqi2PYD
EJXQUWfr51AmnNY+rVwHk1TWPonRRF7g2tHLfh3DJw7JfhapN+k0B2Kv4R5FPlBJ
MkBBxW5D90tPfk9FxzvDszcUWOUj1011/0ldtE99zoR57tYecVJwWwsieRBxIFJW
j+SSgSUwHPYQA3RI58oUmSHRAyNF058nmTmmXgJZKBQld8L6IqYLrrefL/qsBRPr
elKvnNGbZ5F7tc+GYWaTm1zXIr3J+lr89bbbpxoMRU5MQFhfUCg9kpatTxBKsPSO
dIOrkzzmIadUDSIVnJF0/bRAHa34iSXjRfEjorPOUrmEv/CbuaAQ3095ooYuuQPo
Wpnj3iHLRiKwn0zpZboHnQRpjkfwYP5FiirkC6yZW6+Kpk9Tdp3Aq7gK51SOohV2
uixa3z7NS9jD9q2EfuFHLzGZeMO/BM9HQO5isgaH0Oy5OK0Z9slHdpc3mzfFr8QJ
6h2Sr+VEop+vsvuuBN9GVYuZKkOPcq38Zib/8Hm6GG8wU1nZ2jgH62E6dktoh+ke
rQJ6BIGsuiCZJK8TPuqYpaZfVRy0vgeB+J7XS4HbzaBrgmk+d/bhJADTVFgGH22n
1Rd1xBnSbClqPApba5674Q7/mb7KKsNWE2GF+rsI+kWaO7qWxpE0+vvsCjTwlwFs
ZiguHyy+xGV5/SiB4FTq7Dp8sy7SRmWec5hfIgrmkkx852spMukFnhvnaQvO6SsP
hAzoYznEVPgFMjl+qZe1yDCTEela+zghSkqsTwOVuseUNZ536XJyGbuG+sCPIvAV
MNYO/Z+bVLF4e9V3+pU5Oh6puMHtyqW8mOo3q91PkJCo1CJ38WHheLedh9Q+IA1J
GSZQ3zvjHq+nEzLS7CSqogfF0IcC0F/1CgjF88Ke8GTOpdbpBXJ4n39hRCfMD1WA
3qE/Q/f/xmvuoUywy+DMSkEU7aTIycwNTbhv5x/wjEfyl4APVFhkT7FZ+M0OCp9m
muHJQQxQ3I3jQmLpwvS8EFrqly0wbBYGOtzUrRQ5oG+5F5YSRzNOWKcP581dWCEi
AS2I7nsIEqby0jyAIWazWfetudFrMU7KHehGFZG0zX4IYzgoYoL4h1GMLUeoGXk+
fvvqERr8zznq08l1JCynBofJLRy9f7vLd8/wILUuTt1FoKJhOx/UqXbPrh5zMp2w
RJqBWYPGEtHRHhHbwbwbopvhIGvNpdnj08Olj3gRBJijK868s28qRF5aFib0VVoF
TDzBMQYq5ilglF5/GymeOLGBCUx11+7tERCgQiOeaCnUbyxjPEMCshbZWDCqNIN7
/+Zy6ghMrEPhS735y6oyuk3GMDnQAblEkmldcXWOVSb6cJLWeFBgH0/bpkXiwABO
77ebOGUSBkvxjl16Y32yjosa2Y4NtV36FB7qTXRwtIbwHDhCiYmbFggkxAjxVbQR
C8Hzgh21TpBxjznz1Lr/uuy9mYzUmF0HetnWjrClxY1Xorx/WQwMG7bA1rlZA/sr
T4FcuKVA4Gg/3bd9a6ig/jYISFEI02/Iwa79Z215exgXpnAPtWcontjy4GO0od9s
2q8ACVeJFvLY7q4BOMMUgxPD50zzh6NdrjnS8z0DhwBxfwD0NclDxqnPjex8Y5uR
2r+8ShWz1meJXTHwIR9V67QC9vd9kpTetuluWk5jgH+pePzqqexPfRRbeo0T2Cx1
sgvF1HkSOVWBEmHloSRd1YOur4zjki2ySBjF4r4b4NNt4YG3Lzig5oWO/3nUjQbl
lPPoq4awYy+trLZn77Cdh7lgqhbl/JCMUEMhnoe2Nihs8zQxKkkt0K8seDieoEx7
3nC7SFyFpj350OCd7basS1k8CdHR4uxoZrkoGX6ieVJcoAXzlvuLxqYA9sSegDmY
YI++TzmAyrn4hxz48MdHB4698C5Ix44xcLVzH5wlPDuWi5achZYtHvr5Gxghy366
F809N8bxed/+EZqVEcVphasdUyZagpynKBKgaXGnN2acv/mlvL5ixR9RBLDsh/w7
Qa5mg37xqTtXY2qPTmxcnYcwVWcrR7hSLAk0b3JimebH0Ts8K/Bbd0p9C076ROgF
MN5m+9kUdcyDpLnIwUier0+Erjf3h7FQci4JSTTLqE3TYcQsjRU0b4PKfY/h2ejQ
iTumo47rO+g/z6wNPCJoVZvBsRVpquRvkmbw3yL8W+c6GfQdjCj6sq8mAtGFQ+fm
PnWVPDgI5Gobt3uPmQqXDvX0Gw/p4aeUIxThhhG8W7AhZhaix+O5jDzFBXmew1e3
BjJphoePghfXUmRiQrfdmdNMMMKZuIH7aJ1ER2eiNKeppKyDFJhmrbyVpmWNo5gT
aM1sTdnrPfPk5Tayfv3c9TKBml1nlM3LDMoW9Lt6aMsXL30cCUnyqO1FrcWseGjx
FhSscuWK4Bfxa3Sr8TphM+69GXRKtVGpwPRfuv6HWePvu2tHqoI/XZcZK49m4eIE
+IdAzgunHsD9VPU+nogiYgFtrnixOwc1xo7R6kX4ldciaklXiQG8KvI9310Z2GKS
nEaUmf9VrVVZzUtnbf4RHuXBopLeL/6Cba4PRVNiJPr1UqEKyK1wX3mkuuinT4/B
MZiHGDVctizhpmd3x9fmhOlq7Pz8sVJZMDLcbu+D0CzCmOcWj/WRPJX/AMEgsynm
q9RrTUirJKs6TVJqdp4W7K1rlLOTR4j2tuIZCyRROCoh0nBH8eqEuYNc7ehpfIQV
wefDv62JhZlgK3uvGQccEVV/gx85XiyRGlx8F14NyrS52y0YN/oCD7cjIDmwhFKf
/BP60G0IAMAq3brAkojzMoJzD0gkl1jUGzxUfZY5ygcpwn7CRtsJpV7SCK8vgbVH
E0JimdExazKTHA6BDwO5e9NI/gzan2HvNS1+SsgS8PDV7tH/jcby1IDpEjDuTWEU
gOonVI2G7Kw4h35U2FgPvtg1GUfHBdtkOx/+geb/1a5/+F8PZ5SJJ+zKnM03/Zv8
g26Uh+9/uAzwmA3UJU+fVHU7ZkXjXF7halWX5EUAWJ3yd66a16lQ9cFBUvJ6WEvS
RmsG/vsCAfWq5K1ggMOIN3Ddyt1Al1xUr5zCyg9dyOE22jaYFqaEbuk5/Czi11c5
x1q2uCdf1JP4KSJ8boobOeKt6Zkn0CjCL0mgLoIYVUEv/Jpn3cqyE2vUbzj7OVOU
rsUz1PbJbtGo5rpnwHDOD4AgQ5y6NkJBrfvrCoNEuvQ9CKgDsPu7fNq0F2Sxk+n0
kbdyR0QFyJa9nJftuZQZE8ViszGkli+APKNCtMbYx0vR6SzVAml4fxFctwqAC6Ei
aPdAdqQvC0e3Lon8Qf/MLWutL65F6z3VUSUnBwlqxT4MwlXZxbYmLpKrjf/X0PB2
d2fmUl2Rv41nIfyXkmDqyMTRNcEEr7qlvCDuyC5IVZbZOnQ9RuUz0ZAQ1zcw6gjz
p4OmQB6zLYYCNh44/7gLuXv4CrgGhbJVdPbS6YechxWNsQKDdlGVbOYWmpi+wxVf
RNdYmr8mAAGhuHUdenEXgF0iDPRYYKT/xSl7CXr7PkJbUHwj7nnhy3OdsaulUekD
ZyIzB5LZcO1as7aLXPOyEzgyBu+LZH7hNYERrDdbAGbqSurnRa/nU66PAF2gptg4
gJypEPv5wA8+FmB1O2ZqALFW+7osGy3EV8zl60/rBd7v3jIVOf8w9gv1uN8FMPv6
iiQ8iPRQ6Zp83rj2IonmFUsQyEggKskC5fy9YCDD1Akm6fATeB7BMJ3me+O5BLWw
03lQke7ddBai4H49Fmsn/4UYjw9z6KxXltLeNjsIOTz/p1GP6FcLyFZkTODbNE/U
DUhZG2lrnggKFuKIn54ku5IFTHHGpEndXSFBpmOGmQ6zUQXHgM9YNkQDUhXxM5SL
e3JUVU9+NXgTo5OpXaCt07oKY9/Qb3Pwo43OHH0INdpl4ToPsC3mE/7oBYV+MGHv
aGjGvyeMtZFHOkyhMC3vcj3mlcfqACWsygJtVq59VY6GlahOY4hu9DS/X8gW6IvD
vTy4b7eJs18nnzUGwJHim9cb6sFxAt11J93wxldnhdJTdArWo8OZ2qGP6vNED0lr
gf4jMz+xbBbeRX4083guu/r+nWit4X3IbBJwRSGB+TCxbcf8asZwBuKOHCicFGNm
6s6VuugABMyoV6aRc0Fz4Cn/uPN+UWHVNgkNGO4pHN98cX1coi4dG87E3PLsQcAs
/t4uEz1MRqHCa3TPusfWfANlDAhEBDZduPwflFfi8JcwTloqM36pIbnw5/BFcKxR
cm+YzXa0Fd18TIJUFTo/mnUkWst63+q1Gbk1CgYdGPde9tn9wC6bp8/0val9/7ld
5r9HKcKmULFH8BX7zVdUV5u251Rvo5x7a1ZdM4Bz/kVy8aF+cEefv+762nrpVmzN
qHuKGlfrO+xltZIGqb1s6FiCIPRSF7UMFc9E45AkvKPuvloAUsGtFPwU0qlXxYGb
ayES7h7nGwCxdy0RGmFIoS56RcOrLjrXE9m0hbie3FcRLt20WhUdicT46dOG8JAj
IBXfzdBggZms418e59tGowVT318u75Dw02avBNG7rG5FWFPI/5Nvs6pO7GoazrlF
lE3gSVBdf5pqIfFpT2Yw+vlQpBSAIxh66Z18bmjxfDyjrstsVWRU/4Eh1Pv6iZM0
Q2wvNhJruw8JXM57B0fw4VO1Vk7p4rtcfIczSbQ8J92SuxwpnwEyDOMsTZ6AKDdI
pKBz17LtgMHTXaz3qktelEa8sAobpN6AGZQ3GN+syZQaYsqx+Z9pnG862hAUe5fF
au/iFbxl4lmXVo+3kl+Q0h/LPuZyT7BC9SXqxyqJHSKoByIAow1K8sJgsgkFFY0I
pS8n+NKf+7qeW6ajS/ZTp3mqX1WM90CG+LNkp8MTvD32ZJiR25gtXgNrDly1P7pa
ROuDyUImot8dbsNLifBHhfisE0y95WTH/PN58bX//xS5uc1Gp6ksXubZk10eYYXJ
nDHxrDVskM/AQMFlY8r7vGadxt8uXH5x+AcDJGv+wM+ZE4hZs82DLB8I36DTave2
eig7biXqdu5TKEABmLirivHt1nLyuSBQ1saVl36JYU6WfFD2FKNNSAQGFpskJIFL
BJ1tO1G+cq9Tj3eAb4YBYCGJjteTTH2RCRh3/5Ppd4T7uZ75Q5RScxCs1in7Dr56
tWwO0kdxWDG4Wkc5CkK6uBw1A/XtgWYAD+DiPBpXLrFfrirjNIxcjoNvDW5hiGPG
Ejw1mQt2T3zE2uiGfLBU12RlvuofpmjWNMxuOPDuJrAty7J3FotVu7NB5HZuHg1R
OmBq91nZa1rrInaWY3/R5H/+APSwZkQhqwrAHGjDRTypLZ58Tp+jGgX58lNibhld
kW/VJ4cRHuls2+HG6ivaAHGg1659O26fJtiY1WmWy9anMTDOFOtJIMdTY2xIU7ZW
qBr0lx/8WxCB8Tr5hKhxENT17rvbpf11vUPT7JxaUrYC/j4l91PEhsnHSGaSY/MT
I8x2prGZABKGpcLF3IpL7ugE5ykywCMZrk81lnE96mk4D7DYZ3KiBhdxXg7CtFWo
EIpgppDXHA9tANnQLNePwKNSSYYStEfeaWKaUwppY3IXz20U3gHWUQHmPVZm9T0K
sk7u5+gJwyQT9oL2rtmZmtZhhTvk6M5jQ5xaMs8iPiqhh94CGvkR3jUZAkY+IbHp
t0cpe3BrHnkzPdtNQT0GVnyYDnL3ydryzcyKwaa2R5AWvl9LB5sCHqpTEfKG2VOa
FrkpVdxrSVQTIJqmI8wvPK78L4/LaM5xPRcw+Ex2bLzuaWZ8Cq/F21iI4thfeXGl
Lxe4bih67CSVnsA4vTuPNlX3DnZbwICcDguDSZxv/vIpe0gY36+K+x1E1IcViXSL
v2t8FAc126eazkoQY50AdYRlSzozHibNxw+MhOYAu7pkQ+ftTfXdY24vLaYMHCOt
/UdIinIHiiI2L+qKublpQnQ+amtjX8UDL2tFirW+7Iiq7ODutsHkGH1/92wKRZM3
NUuUv7+wO2EoYqIv7/9tJ/V4JEjJC/BHJ5BdtgMB2e//62v5SMJa0JpitwgIetUZ
YJUQDV1OR/HE3XUdsiAMx4i9ppjUiISBYGrxE3NslrVhBNA8zfn/i1N3EoPL65Fg
LobOiyZQZQ31SPfwBrvBZLjsN/7jkXnm2IDop3y/dY5JGES6K7TZv4b5UMnR8FrY
vPxCwMOYiT52TtpbplcTqs4/p7TBb2OPl6yx1mN01NKwFjTU8WLuZWoBg4aogNsS
pPYmthQXjaYkAs2b8rSyYZ7EXF4TP6k+RanNLTRA8Y+um2BfGuEcFTrdr6hAPiRv
CmKAqySIdRAPApTusX8D4oayJrIOTUnX2Ogv959bolAS7HFBqzcDN0NAW09O03Th
tGFZvM06dW5m/xl1vMDfEga8O2ET7k6BQmRGrD1aXo2twmGVo7PlrxWBDOuR6BYY
JQwa/9apsi7avChhcuYT0N6vS/hnQSBqPWCATdIrl3bvI2nWtc7X0sKNKrT3LD3U
gOnBoCVA0tT0BtGirejg6eo4w9oKmRt1ljDY08A57GgcF8KeF8t458WabpK6ly7w
dYflJAaC5gqdy3lyiUc/VMb6LW35ZqkGo61akdd+7n2zh6xGRH8H/Ua2eIrc3Gok
KPsdJ2sh/MjaOc/Cw/RBt3iKUbgEwqQ7AgM8EuYhy+RPRTpFe1RkLMSEtyLT35Pk
s56bR6BkiVQHX6PMeEeO7iBkyDOO8B8cy9GLvKWlOuDXDtM1xXnqfcfqwAIgNm/3
nMdKfZ8QRpK++/YMI8UnBrKtc/prmNNer38WgfelelmdmfwTBgKIPsDpCeo6ERPG
Tn8RtloXFCLTsh6vuRU5t1gEoXICrx85S6DwkucVmVAOL6eiTLP/9cUXAmg/c/z/
18ZCNwyLMCzUIH4oaiC01dWVJ+qRhwajaXsge3zkbyJbPi1MzsqlS6VXzPV4QmJC
fZ99ifg/IknaOSzowRu4huwV1GehUOPEx0LVMAboPDbCFi1QFREG2EIHUjpmLAd0
Z1E/uquBeyI8imL1KTnRpg91JZPOVvDJObIQFqTdXbE1GqZoxHZ0g5t5jlq13WIh
6CuHuw9BxS6g+ts+QtIVK2MEbA2zvKxWHX9nlCZMYpm9oGfp9HDEEVT6+IuNcaE1
J8zHuUosicNT3Gms+9VHnlHhy5gKYZp0gjZ7k3DlRNDyedqgCt18La5UnaDFInxW
3tB/bdHgOg/XogofYuoV1LLXGfQ9dwe38n8FBmwJAqZnKhFFPTQLyBnZ0kjqDzrg
tLsLyXqDmvix35guGZdlTXqUPG4+bpb6sEDWst4W0XmLhzgI8jSJYUd+RglR+5qx
M/wh6zFb2bmoFOJE/5Q1rf4ybyWSIAOR+52CB0HvP+RfmjT9TcxdLx4GtEoMDylb
40q2hLJf65D34klxD7/V9IplGGmKuMVFoWxM9bVHBVm6e23sF78/VzK8nqI3+aix
6DMhawHupj8QmBv0cSMMz0iQLgu0ziqSubynGgzu2omLE3X1221u+mMCU8cKtg+l
C6QiHMxZ/yUEoj7bMUPEqN5EJWglA3fljVA26FxqvDMSu3tkjwq/yrTmbDWhjQ0+
KLvj/LgyePGr6NASm4SUhgAfeKBqzLWPe4V0I+vY561XvrP8JzV8w3+lzW2Y8b5E
ucRPgoaOW2roNqVZ+lxVL9GJCTapIn3TWLd7j0RqBcDZrzfW0sMO/uG3Br2F4IYV
KwPGFX/uaAaaZGjb8vTX3ITiRO1bNOzlWnUM4BlYtH27NcfQFyzrTPu7loO9hI7T
O7PdmKYIcqhw71Vv6jzlZXxQkagDtpVVoK9+zc/1h6nx3gJ66GxfFmiS4eCGy088
7jqem/tqnPt2QcdOiARxyBLxH6CBHBoAS95CChxJ48KP5DIXlAtR8fFriQbfdF8V
naN8QzvLuPgQCHXXEvuERQlXSXJyqbYc1wi2LiqVeGNMuAGm8XlJVy2eLje4NbCe
wnKvBRAub3oyObO49rrHTsehhAGBKQGU8Oh33fdG3cn+vgZ0KR1U8MvEe51VXCZx
QuYwcRr9KyLZhgdtYBZ2T2YyGkTjWv9MS32iSMdwKoJMX22+tcjo2Ze4RN7H6vIu
Ea7ojhSgsRWhB61m0aT1c3xbiheplWfSFH5a1pXnZeF+nwiE+0+nZ0QgwF0unHrK
Wv9cV8ejjm/tEVbnWfF1WYTAVuhNCzq3NW7dfQa5Qu6Dtz3UbHa0+GmGLiPYcxIG
PoO2HAwl+z+tjn+Tg6huqCoCPG8yDEXgehVRSFxBMvLjZObAe2fImVOYq0YiNdcI
cjeZIBhHNsTIbhN6fn/JRDdd3UGYhPs9euTAr5ORP1p5okyrwrHYmoCoAMj4UwcP
3NGZdRDRAK72Yy6mVPzbX+18zReBsVsgpuihHcvLrFUDFTgA9oP4jiOeeCYqh7b5
EwXGroiLM8ihwJjfH6/M/rcFagMWEz7fGIWIq7GDu3QE5ydXM5vZWoxw1qloS/v0
TTZFYijolpfFqt3Rmhml7Iag49EIgbITnA8OU9ryVgZQYCrFzaqiD5cRAHgqMkFi
YD++s2upaI//bnL2lHaBSZTGUJMcICNn5COnrxPXqG/7zcVmsy8i9rsQfhE0Trr2
i7Q3p8CgljGVq04PBN7EYvR0Knmi9p9f8tbupb1kCFqtibr+GHWug6DebrFLev7H
ks0jdi35dWFhuoqzPDluHnFSae1YgsOSDsezpgRGk5TZDAgtTUkXAocASBqDZLBY
5M95KdndaKtbbyhs65hCrwHFe8/zvt6UVwrIs7nz09dii7T19upKD7h3VC/Culh/
xD585LUfJ8U1sIt7vom2xRvI7+IPW8EbsvuYWgGDAN+AjYeHImAbaHEfuE3huW4h
AkpC/ruEDEjxWjsRh71ysIE6ua/pbMwO2QoHUP1hhgIiy+HIdJAWyddY7qG6qooK
ZwNcg8Xvp9bPa2ZGEsbl9jll4tCcVF25thBX2y7HULkCJrUME3P1dlaNfRAjyykv
R7YNvXWjET1NGUKt4IKh3qaPy43RdzfCxUYGbXmyxWFXOB1RoJR1TFqZXHVNOGRS
C91/yvbUmiNIY4r/grA1Xly5Spm8pLzKrAJznqdmyfT4xMX0ptOoHkastEviwxSG
PA3VWdSXnsbo6rLT2LBor2ddBVDct41DET2CFAPtvhM3T69O5cicuyGftEYdWQHZ
WUWgTyl1phuJ6X7Z2lEJs6jA+s8JCEgGV+zTWg2zYULm43/wrsCIXOzUinWFKBll
SiFFOLyscsPVn2dTEn9YQhfHoHhKXRE0uLNThapgqx8/dr3GUbdHeSAL7ixuFWjY
YQLGOCPs7EtL/HEy7tNf6XmCMDv+HeOh2fD1KKyq5Ad24GKbD428M6YYN+W3NG8M
1WPwfXz4ez8rJe+Q737CsqlRVzL7xwo0KCDjYTmnVYl0j5SVS5mXAVP1NIcOiWH6
z6kldTdkgsaMG/PvqoTkQIVJ2YtXtylA6wAD46EFqN9Ml39a1BDpTQNC6TE9Y+tz
mFP5hdhFR7kyo8sWxDUUiW4bzw3Eqi/7kpcu3kAHrFuHuHloyeGRopNRBd0B2pio
zeBBY0wFgIdV/461tG3RLCGUi/yHwT/4Di/6XDgGTmL3ye/YwXibKRZktuaWMVpz
a2K844N3PxzFstpv1K1GA7t1fLjLGaehw+/mvzD9F0OJ1FL+0GLt3l285Vy6ocwm
gfXTIaEvQNUUl8g3h70TVV6ZmfGYlcwPNhYO+xwe9lFzMEUYlLq4UMtXiwwgRkA4
x7rEGAkPatTtCs9Hznnd0nZw5iLYrPrw4k9fAGgjISc2iEZ+xiHWYZy94KZ0YVW6
Phk57+Y589Xv38b4CbEAt2gPzSv1I4zol5I+kCXEOBAloG3WI+fpnlYpmIeyIj1W
Fb6csnkoMXzztfLQ86hDlLR2W8qeRXA2dqzrXDR66kiDmesM9mrBwXYeLyhb1kKZ
9OvMmZ6dKfjehvPXXgouM/1n2n1rOnI7AJXzPyIhgJtnrXx6W4hs9B/sG7rWj5E6
oiSd5ZAwbnsS0syBLZoxurbcKC3Cv3PIVbMrpWoPTUreS1GekMe2p1+OxLuUhJxW
JcOixCno1EFzOrzkxfAkrwOwdmuCpe6k7xzFuvZjtyRqSKb4NsvnMF1Jpk3esxBz
4i2QHxfm3qV9rmeAppKl9A0DAoDbqiFt4tsLYfwyQzRpK9c3XgZ4M1uQlbPs4G9t
OePcEs++CIgksFDGvaqucEW/FShsJaGkzh6rtRSU6gx9VQL4ruFRkp0+FqH1BOGy
r9drK8USED5992j1DtYZXch3M4OyOPrirttfrqTXvbFJiIz5bCzKfy8f20Gl4s3K
PjYyEpAsheCB0H0wK97nzop28HY0s45hI1IrqrlC6J6ljXQWgVzaSgzsbqK66+A7
NdLuou/VeQsbpFc7PfcOeKNYDY87mrVu6paLJKQSggArHJd0Mx3bYmFEXtv3us8D
iolvzeHR6mCKv/wUsHvxPyReSoMyzG9aOswCg2ZFkK+WUbzAePMwabk3pTf8YlWs
wHh0FbNAJ+RV3lVquyCOYj4by3yrXHjseP8Qmo8uRm/XUZf1BG/958wQtoxPL6i2
1Kye8w9WWwPygwl7wgJUERwiP1YazsAqGt6dlRI7ANeTiYv1h3oxQDnfupYvC7R/
zZ6+0RhVKRemv1jPKJQEEUNAYq9qAg7su0kJJxIU5c2+2D+NgjSn3cfkpCQanAvQ
dz9HBbu60xJnMEWqvy7y1dvsHbWeyl+bq5k8VPLEsUQI1icwviFFbecoWyA1651k
nk0PX0Fqpd5bdnizmYYO85V0NDQcuGqXyAoCB0AMbTX2zx4VY1QejIE739kqe2Gr
GYlAIjyuzJOQpDrZM52UXioGgGFkYfghv7Y0HDhbKVAgYCrCwYtNYXJ07mHYBV8m
lyHemBsWazTIalsg3VDGw7alQLDqrDEbDWWC/d0NtouRFen5r8ZomvHyAuvmQNCU
7XENdQtXIS6HEUtr1SvGAA9LYEncPosI87IoXQjDhMgGUtdy2G89PrYL8wcUYx3l
ikwikiNCbnMMSztj1dyF8z0hgSfvGDLSs9u9f9egcOQnR9JqgP5uxUQSpCfDnoRy
lhH98Yh9ECeBPlH142zITyV/aA/OBVCseV8/YoB4nYQLe4O6520e5w/phFeK3jCu
McxC3DB5OdrWeDLUsoWuixU3LyWq6TMeXb00jo8gp4BTr6tDrTfRRtkSb/bxxA5e
3E2xy+r80zFQfqnQaBRmn0IG2xE3vNfRln43By18E/eL3P4BUk/vOR/KLL9gLKKp
VXY9a0UjXIwKL4N/S65t68i1V13EXcrtQatMY6whCSKs8hoakKkQebf6fv57TOi3
r80zPODU/hbbOWRPh/qsiji9Qx6shPVbsci/APyEeb80POFV8mfSIk9mOmr9Jy2Y
mB9Xhcb+1Dik8Z1VEdqLOouSQha13qRMToQ/RVcb+P1tTeMmbVJ10qKhHjgGv7LA
tB/RpLlwZ1+WC3OqDI00ZoJpezl5YFEHiqEXS5b2mC1EMoIrepr70eOKCsHlAws/
hUJZB2qovHJNUyHnUcqz/OqMHTif2Mh4SmHtdYJQbJ82x3qYIMhrD4oKCVFcfQ/X
ve0v+hCxVSWhaKv+g8MqmjbdEDoRXH4swZu/Nn0mjoY5YWUefFEZyn9ZhHlNMpcG
Rmayr8A5TWmIvRXRPhTsbgCMPFYh/+qDAPC7fY2qLDAVa/y3WgJkMMibEAfAlfeq
IBa/IolLe1y7sPTUSG0QVfmE63HH0pbtsQpSsUQSdrvT9m0wJmyP6c05NipNm3Lr
14cFTgRntnC+Y4uMJ8+jKppM7xW4y620sD3AJ+Ft3MiedlvZCjz0oJwN42FZsgX9
crxvpbI1DYLG6gWaD8fgFg1oLHhXpJMG7s85JVBeoB3SL8R+0+1eoG5qwYybhFgc
dJyTT7ms6EhGWJuLM8j1i2YcSs4fsxiaxYRdoRCoUVxKTOd4PDzPK+WRj1EcqTpY
zMHy0KFhhKGi68kdft5kMyu66BJsERSaQ1D8IBA8Cd325STAPpofTGmjoc6K4sLB
XnpfOubSgn0TihR5nZPhq7Yv9n+0uBh7WVk2b+MA0XmNyQSejejqOVI48URgdCDU
7bP9tHYMRLftJMYqwdjlL1HzOuuPFygBHb6Kza2UxnMG7p/3DYpfspJ0Nsfdj2+C
Op881SIpp+5MedmsYPxYLqVD9jIYrPhwfLGZLr3H4n0DmvYrGDd3j7fZeTKODTvl
5/neNHiTkEOq6wMkEKa3h2o5zUEmJNmDgSm0HeQv3QZF/WJTZ3/kzBN35QlSX1FE
XtjknVjkRGS/Od4MTBHbN8oMul9rM7Ikw9DPXUWAhHoLkS/UkIijDXyaniiH7NWf
09kb+U2k9TSS+YhJP6u5JjspYkCcQac47sd6q5n1oXQaOvneq9herBB965lJUFPr
xVADrcCqq51saZ6B7ERto09b15PUM8MUYuo6XJvVB66k1kOXbP7rFQjgEgrXC5Oq
TL5pJuYJXwEINenqj2gipLU2EYJ5h6Q5MyMWPm+iC+fvAhjrg2kLCewaQeK89eUd
+M9qySKUwSxhdCyvFFhdLpmQr/ZU6wH9EEQg/gGwvQvJzXDyWF8renPNDGwVE3Th
aU8FeKqlEw0Y6Sre8R6wPNkP8mQP2CQR49tz0A2vMDUKe6ml6RKbAn+Flr7hmzgm
2acVCMDtlwQmu+cN1QwCWoNsv9/9oyAmFe+SvgGdMAfd9K0IrVMLHJkg5QqLAvjn
BPzcqYuUx8SV1ynVziv9SEMPu47dr1UwpvDg14RLn03r//0nVBSESiTcrVFLeyRc
rBJj337KemIUJILxKzhscX0n0YJ22unzF5hllF0IOvxHICsOZ45W4K00rT/5UYC2
aIXDyQ+Oj/faSFSTWooTcPdFtfn7DDNKb5F2r9JKjmgCbI8z+L7CFP+AYTV/fL5S
c2gKUUbw0SzVu4k9n8fTJrDdK7RimuiHbTPPPXWE2SGpp/Jif+EibP4hyKEZJJUg
xBZRq8p+EPErpDUTdfyGb4HWivCxry/FaNzaINc6hFwZOe+gsH0zOfOlzI8UzPDr
xipcHYVwpFtAD36jzBV1vRMdLMHQYgNQ+KJeoXx8iTvjT9DAFkAHbAaw6nTbK0NM
vy0CmrUBrRbR0Zje1spef4wiiLDLxgtn5me1PxrK6KdSDRpK0EIpwZk1X+1GUBuN
CSltLRTk/ecvrDYg7OOq4KvIyu4ll1O6BaBWiCrMXyXn28CxVVv+du7+y82Ahugg
CV6E/bvQogiU2zJHqEAlTCKRhrycQKnnV4c4zaYJRcrLeeRwKXhh8LMGD1l8Kq7Q
wA88JPRZBu2nUYN4a7WZD1GI3gdfZT2lMMvmwK353VNk919qu3pJp+9u7SxstSzP
IEu8lrYMUaH2gcCWP7CAarDMsEbADBmCdCNElHgMw4x2dVk48fft0twJNNItgxJE
tVA2/R6UXcdAaOTE2gBPZtAaq9GIvm+FtjfgIaQ5DNKwfznpPM0JIK/4mq8oLexz
DJ2as8oMB6FeDR2hgGGSBLyiWywnKUc72FbVZnzT0imDyyrKS5UFMpNy1mPTOv6F
7h/xzeNq34qxYhvaGOdWdL3xSTUT3zfmWZ3pI/Ve0pqThg57zObHWuDMNYMsPoPy
1691gqIk6bagfktW+Wn79R07rRghXnxIimIqKrbLPaI9XNKxTIL5pUso755k5o17
UDfqWkai5Dfb8BIS45NHXPidZd6FXh+PQkmh8IM/FjQwaIWg4MhynRh96mIQny8o
3PD39OF41pQ8Y3fThVfSvYK91XQPW4ny7ORUvHnOCoyZSBkLzp7GQ2Jvah7sst62
dxzkV8UlljBNU7JUVPYNboTQIcj5f+/37sqewphq6s1vej1qaEFOkNwVKAvXQIiD
V3SoyL3zrBCXtF1xHU8PCOCvXMaP4Wl+dTJYgcH04G233pOHm31HUQCkQU94T5Zj
ugS2WQ1UA2obf9lcnyzfiM1wmTMFbiUS2yhfIB9qfvq7MXkweqEUDKezEiCdCQSs
hjNs73Qo70KhZkWtoHdn/dG2xHmdwsJJT0iFoUrV52Swvc12NtAeRMzfb1C64IrV
EZ9e5IgPXMgfq25K4I5zw3fX1eJvYNuIYAtbMO+8fyUjUsJPwlx6DZeRcvIM//KM
IxsfJJxUqsZylwk29/swkCChVUzb/H5pANQqZWgDWNiZvQJI815ZQ+co/Ddtpxbu
kZktU1FnXqF8FtV4whD4NOtvb7DOOxifBWDcl7z4E64SDvDpi4oCjqRV53EKqB8p
2qctUOoy4yfRo0yFNTxVwcO/ZYvqJgp2oer2iV3LSIIuqamUgVFKifcw+vZz1/j0
/IzcNXChyE1NFGe8++Z/vJzvGWtRjRZ+cO9iWGMhuqUgAYDf/K2ZbD+CQeYrYy1M
G9PsIB70zTsomkFDfpaa88WvNtZylF3yRi2CE9p61U4sLAgu3051MIgit5CaNqMF
oVnGDs458q6R1V0aFiUkomp7XRVMbzSkTw+HTMPyn7emCPZK7avn/hZ0NFQIyHNx
7YRQIgelpNm0F5Nf8cha58Eofv4vAwjIS/oO7mUfKm1rogX7oaPXt3lnHxNPvzQW
UwqXI5WJuD6SuMV3xM2q4HaU/aKzI1iDl2z8QpTCaITLFkWdYR5fU+S9KdyAuTVr
hLB6CSG7r6sUz6qfprV4J5VgS9uqL9U4GMLjrWoP9HQmypmgfwCfuAt5W1MMadGZ
bVmpnsKql4lgpjDwRUjVlwL2AmZnAIj5elrhd2HgXQ1pzSAk8j3YSHXe7lr76ig+
PBA8w1g9kd65+8bQgICpGKwEdgid7bBx6uDow4Be6wPSV15VgnAaP6hIPYJ9KmKd
fsRUV+hyzB2OZ2+EI778+roL6PIEJq11bx8BAOwcJcRGoLMxArksn0zlAytbBnM+
+KwaKb7Y7e8KgHrtjZfr3pkVKdbo7XwU1hXTKmp0RBEdqs8q5EPSNrJ8Hb/74QDX
XsARkxrDhZeThIx7iSNnXFd5h7tCSQpG8awD+FKPeeMcbrGOL5cQuaiwguAOkmAk
YBG62By57Dv9rljSUnw1fq25NZQkLhzHzf7LNAKF2eus67ew9c+0QPjHOT5mUIXi
nmsrL50gDTYyTtB9k7pxS/KNhswxAHrDG8veaKsv1KkiflS1wuqTuQLCo2uZfGTt
7DvOG5sv8jIzoygdOgB5VhW1Bx4PJI3CaSgmEmXZRAxTbiZ36Q3F09ksZmL32ROV
zvbgjhW0ErZqyqbMWuCKFjdr+7gDW95/coCouWU0a+K29uq0bw1Ve3b4TZAmXr2C
P6ku6O7uQx5t0FLz+oqWwyCsAwaEInMCEglpXdzakAL7UmwahMq9T2PDEutyq1Kg
pvimcYHebQh2pS0XHYbj4NmDBLhqIswdksmA2xnatHfcRMBPKgQ2kvU3B9UAg6hz
NJfr2plSGIf197VO+3Urepz72pn+32SlW+9OtehwW+9XwZafFP6ztReMPRCSUppp
uddWvse9o3ajdW4tITatzOe9DTN45idW/XEMB9wbciyLgZed/FSEjfwCzJ7uaOZF
2L+JM8oiy6+9h5hq2GS6jV2mquIxPApYQjCyXlvbUzzXtfh6HSkSXapS5+j4Wm3Y
6gaoFkcGYCGvMPWkNfCSaXMNjmUs5W4cJr0vuHeaBXug6u0NQVXKgE/TNQhoe6xU
qPIulQNDot634JloFqbhJ2dIG2kuZapMmz8ymu+E0mxOuZt4hc8g1WakfH897JdC
L0312sQznJSZfab8KC7inDdrnib0V5VmhKM84xnsy77wJ6jjbawH6Gc3RiT8W5tj
aFaIf9LCUWljb4L8LCuDAas+Py+vhOR1ebGAhmNRQUsOgckPenjiHCfX6mV3wW94
yibGGsRKyAtlbP9oOV9KWDa/GxnH9OiNyshZuh15LNSSOmvqsICoxOlK1oOv421I
/hgSiKHy/3oZY3f81tLEu+ht2pFHje2BYzIlHYZemaOZl3p3V0iv1iqU73pr8kAh
78CWdMk0FBp9fDdYDY/tJDj737Q6mwYbijpaYgQiz7Z6p+jYZGj1kR8JPoYewtQY
Z/+7BDMh3CHtFEX8vnXdFIilFqGi4DLWTuRxzv68xLQ+77PIGjbUrYyZtgEPatZA
pA+niMjvgYOdyN9kgeQJ3Jda05B4/3cG/nRjM6riJe/Y9YDJvYc4ntYhfDAVC+nM
PYWolk4nay+j45ZfgWzeAlelCe1gPFuzWPFkJMg/LIEfojD7c+De8VOpiy7JMZEU
b3spPmh1ISqA69tmSeXW4v0petKPan4PbJ/25xxSVFdAW+PhOxcQQvJbuxy9Gjp/
GajDNWts77s9YxTLEwHQAy1RfrQBs6YGjOPtYQYlCChY6SlxDEvdvqazCIthOirb
oUlt3oz9vEfmShPlXyzjP1Kxq3HLTd6OmsSJeDz3NoC2a8c2p25o5zfMzrD3m11y
i5b64ffs9EzZhhR5ZHSXS/mlWTGADSAxegctstwyF++8SsUjWV4DeVTRi2yNBi19
deMbJBIUFEHgvdndi/eHp37PzDdGWpyjoL5W/yF0FXz8qubtK2sU+SUJhqjkfGBW
s/Pie9uMPuwHXcuETXfcHeuMahnxKjpXzBLDiLAVjlCwWKAr5Vla3LezX4sYmylJ
Yae5EFJNNel+M/VQbez4wM5UanbGjlfIAa27uHC8kiQbg/vZ2sn3wDNZ1+5Yb4n6
QEKc51osxlASLZc94kVhOSgwho0GCHdu8UprHXxSi3nnMl5GXjLvKvUFmF16eASw
LSm3hw0bIl7HMmyGHxfFhgUZoFrQWoOVGzAdTboX5oj3WnFqzBT9NZk4DcXFQKb/
bABxbK1S0PqoYPUZEmmceR1qnmyLsSJ87nBE1M7SyYlkKoHJPsB4SOcsTFjV3Em9
4btzOnvtLg73O0eo/s/dbWzhlm64FbbHcCr5DUBVD86Du14NxnHW+6YydyNjGYj0
bxZJBoUgrgaN5Q65s34y8BkqnNE0OF+TRyQoXBsSYA9z7rbDaGk/n+CXYzHgOUQW
Gc6dg4fbFr3vUnyAeeE8VJnXsK2PKvsYmWB5shuBEjU9LoVzXopsm/bNx+u6dRUo
sAgMEiM6xiOxL+iLMR+RtA0R2/hKBZ8zfR/veou5DEmliwyT+fewR5Sw7S6EFved
TE4sHWBFQUPiiFxSQGpWLph8Zc0rCUnMXF71p65/begFWNoYARR4R+8BGPTQZ/+g
KLF3IC3tuVM3ExWnPVMOoO8lJmtJR0KlIn409nJxbQ1s0PAtLl7p27n6ly8bSCHY
6fsblnuBHyEyf/0cF9rNUeQ5HUdiY8kcSnHi3qO4fnsK0SL0qgy5FHqPfjUXkRfG
BfGUlR86Z4S+SWSPj4o1YNitgHs/yAqquYvFTwSl8/KvY3MaX3AD2tmNbkUV7Bm1
5fVrRBZJ0+nQtMdrT6pQ+sDWU1ot56cEVTanetI8jOqBa0KhOqrs5Zf0ACoJaCIx
OPVP8504S0IAcNV3FvCuZAMqw5Ex4rANezmwSNwWUwAdlmn08RO0r5PF5lbLQk1R
qFxRTGAxgvWdaK3p5GLWv4gE2+/PJ0JTD0SN7uoW48m+pnNa7iBM1J7pzUPh+fcO
NcLiL3cPR1JthvarRPfQ4viA2J65pNUmU1jeKdo0cfDtTEQGMcQ/i+EfnJKOPKrs
cNgLu8z0uz+jRRYFAK4Xl4BHrn3VfhJEkWP0on1Xrmkt4Y24T/QxGWPVQQm/kMue
97CuW2Ud3feEtY18Vi/I2eZ0OclVUt2kJjSjFpYlfc+1ydw4n31m3zCD3TtlZChi
9eMC9vSV67JjBLXxl65SzzVKTOC34yZqHwllxtKazgv7VALareZR5GkT/jK3gt7E
mLTgiEVaf6iq9NCGGbx9a24I3px8UkV/Ay+9iRPgo8b4WmBaVuSGFYmv5UFVTIwQ
haEGFyn5fbX4JdMDrDgTSwgOcvuma/SsEaUz1euBATmdlLw8LwbbcGPwhmWwA5mZ
q2yMOywTO8iYIx+7d18UPWloqulvpzY7+z14Ff3yFEb/in7A+tBmddGCgcb1lN7/
JKo1A8ih2lDHGqjePQgohibM+CjwS+p8t1KMtYpo8v4Ahc0E69C8/XLrvZIVTrNJ
Fj9qz0F4FELjyqVBZ+CGE2z80nAx4bgWAXrSWd/baL2ePmoVTJC6fv1FIzFkNCY8
I0A6YlRGnoCoAq6uHd7iqwa5iFuf5PUVMrjYF0BEh5WcRiXyaPuZw1yMzLF5ghNN
9fRc1fSq9oC2JQoRx8J2dexotBVvgptJE0KIRa4/a2hNAT9rfE8bwLuK7fTBL3TR
4gldj9wMnnueNTjiBkpLotwsgkdm9FdODloFKa/F2YilLwLHZJd4NhgVX9TI1ZK3
eh3UqHX7fIg07Y6D3vs+pk8QM5g17HaVzHSBkoRD8SlkaY24iVZo3bDoRTzkkCbn
R/XRkQPmegy0Q+YFAbcUfsOpY0BnABzG5QVdfB0lWwzzNkL0d4C+hSGOc3xouisi
THDUEY0BE2moMOuDFT5Bye0HdVI2pJk30KiZEzTZHbjqd1K3gOM1xQaNNh1Jbd2X
N+Y5/zP7YVBnTurFcmNcc6LFt3fwIDesdaGaZtCYy5oUj00RDj7tiSktT/0OF8CR
18BVXYhDBPjh4O/iu0+C7cmS3T0gm8mkmmjpKJm6/2oT2yL6+XFpShVjgD/4EjM5
9vmSm8sVHXpjS/n3TekaD09vAMJjM31+SLWdYLKniOZWVVt2yZNuM+I/nfL4qnQG
lrxLO8subxHbNHjjR+6514FF+iUVHIjhovMkm76Qwvgr4YILlYkBBIbEdyITCvOF
g7Eh1RSrY+txdHBZXDVyni8x1rHc0pwpAtKne41qvP4IKaOu00qK514Eo7LEpkyH
O0hdi/vOP5LGH1CF3MoKWjHhoFijluCpBZAlGvQ6L2JsSsXDJezigfchwEqONrlQ
R5mJpYuXy59ZpBBRO5HebU5ZYh6RlYJJqulTJNrdlF6pFzf11pE9Mxgl3Pw+zFaG
AFcVjG752Mt+XHwcIvwvTfD1ZpCL0FJC3GkDQmiE93Ax1vV4O5M5ZY06BCT1Ar/F
jG39IJR452E3K511jyalM5OO0ZYUBf7qgpKJgXALoJOaejcLS59I8fH9KZVevXUs
qORAcW6BQlFhFBSG4w4/Rsp2ULy8hc+Zj8ih7/F3KbS2l5Z1en+s4U/1E/rkdhG+
YWnzQ7nO6x8hY2GCL3YJa4723aj2RKV/dnACX/21gw4CTy84qebFvt6O6hjcvuq7
a/mt+uup/nTTI0iiuEqkyzXQcqHVejHKkhL7zPHa4fym8+Z7XPnFBe19nxzC4+FH
WUWADsXo9dPIUpYBcb8TZAnMUoGRRVLO6w4j7WMVQGAM/dsKiGgoKM8OSP0ICqUw
e6oHct2eRNvUwJIZqioT2IcujvvR6kiPx4beOXzeLgaFMHnVxQ0ciHaAey8M5zd2
N6RSmFjTgvvJCsCjOSIzYA8O82asladlBevXP0jC/V3z7n3P2N1xv88BuxEi1uXG
9ZU+F4xXn23Egp54h1YpdOs3Wgw+jg72XRkmQpR38iVTazTetSZTY2eJ6yugPIzY
jT6QrVC6gCwoNA+Xkuepwk1xyGQ6i5DbItfwC8LtpLMZ9YgC/EcBNRlBLvvk827q
35HQmIDABocRLYPKkTk+es0xauEUD8BNRB42qAd2b6XwE7kLDdgxHHMMLOE0VF1I
rgXt29/ho38wnw2rfA92sclqtnnt9n+IVhML8AKPWzNgaJjftm1KKcGo6IB+4SIJ
IreImjnuaDsvzzsUAdF1Fms4ZLqLEdUu+BzZR3spK/ANJT6ZQuP+AXNBhTrlx0uf
LmCvv9OLlDWojaozdQ0ZFg7AaMjqz33TKoQxUyroM6RCwawr4mNDGumdJjK1Gqlc
9D/ai+KpNsLfdVcM20W8vOC4ny5Mc4KqKP7cz3Udy2689yKhIyexvQobFCbnlP6e
BCC2HBifSk0aNE1d1GsCUZQg0eIWtEOJL/s1skrVexcvOIzIEVKWoQV+ypY1phyf
IWXME36oItT6XOecEGCy678DSOdUIpzKKvYK81tFI5uTKApZAGoCg4FB+0Zl01nR
2iHRDoXf0MBckNVGEsmxbTOiZLLyNSJ9qXKMQMeAvyTtJkLYcOSXGf5DbcEr7cR+
FO1PxuONzl8n8odYbAIWIncKTcX9hMDmEWlLAFYwnQrc9BN08PjTBPKoMzaLaRIY
dMZei0TTIL3cREMdDNlfetKkT0pBLjiW3awwyPH9j10GREG0w9tNe8LwPZFpa9kj
TjFsF98kYo9uqQ+xwxtcAn2+LpQ4oQbRFTWZqh1tZFINUDXQgJX/JJLARMWP0sWV
mqDt64mBE5dH/2Bti3zls65AzzumYImnGxfrXG1x/+ApGfm6mgLeYoqVz3xUYLMj
+Aa6MFxnCzLjWwlQAgHI6ZzvpJ5hrYgve62tHaGGjtk9JaKFryyjWiUpxL6F4nZV
uyT+bREP3bfRxz3sTZEJXzmIcXTyF79fUGlUpshj+ILdZhO83jhmI4Y/+GtUxKZm
II8B+tFJ78MaIzx7EfhgoPDzLDwtErXuVEj2C/j621gs92lOMV6puvXoVQcs0bIL
gCuI14+D/vIAyXJXQDvNWXtrjIww6gLGjG8C5hBY0MHdAwMGj9WdgRkAAeSS8RB7
Wf1TeoFcClTH03ci4Ygx6XJlnN0k+lNAOevrNphpHl1mjcdfjrNIDSSGs3nLxHKC
tpxr9uhokTwDtNRmVJpS2gkPRw7fuWLJ78mTXORqG2779pLECOpFV9Wi8NOI758/
vut+6HyDOdMCrd5tPA7akfGT/ylvpitBECYapbx2+GOBMVqs/y+6t31tWXyaYWy9
aMJKNnoTlPUv1gXB13/Ke4gs1d/CzlSR/J4nQSxvQWAcvW0sdQosNSt+827J9Cij
0qvi1mM0yIgjpNf/dY9O4pRg/apg8FYcIqsResw+ZM3pBTC2xyV5hzOUUiIkgmTu
d4A/PX51JU9N8YovzuPFERnwpGxWWZfSXnHSlssJ9jQGDITjWy/gk9YrtjaISJRl
kLW2n4x8PoVZFHwqhYTrPN1+DsI8aHrjn+MM+rJsW+EqkqpkatZqg6NnoSHDt7Y3
22Vstaik8CIak8q6KnJgNcs8nCyqt5nlo3b6XzSVY+k6OwLA8hfgXBdVnu6D/D88
wY2ubEjvzva8eCv7BjR9NZvDsl43GOrPf1tersr9xlwRn05Y/40AtRr7d8xadEYD
okIcAqEE8YFTVBIBkFpuH1guyUtzoJgr+x1pxWbpONvAcWvCe1kMWSR4CT4zUGa6
PldJW3/OM7Elv5dhAGyaH1M63guURCcc2zu1sjnDe9f3OJAN2nt9uHQn82JP5bkv
GwnkpNkavBGeWiDp2szVjIzDoPX68Ylb45v6SO7qp8rPjY6gNGQgz16AH14PBWEf
wAUcRKU41X2GqT+t/qz029Te3FL3iAeE7Fx4FIzRsY0j0/HmXVW9wt6yy+E3sD8A
p1r0KVlC4yYTFdsJCPZg/YaJq8DWwZ04raVs31abEuKOTMH5sOIgCjsE6NLl+bYv
glD6NmBNi/iuO5QrnF/vJPu+/7wYXjU/uDpvxcJglw2TqT1NyyaItGc3yhWZNqcB
M3+9KyMX/7M+aVNwBdCZ6H1KKZoJiOUpc+4oPVyHHmPOiop0yBdCVJAXbd4B2y3I
nLinOzjEF9XOp6GfK1p/iAvXtcbpt1T8gJwonAu4ukY1uojiFGXc6R/2YeDI5DAx
IWTWLOhjGhWEEJ7wBkHEqnk+6Prtt/7tWh79Lwd3kHpnIIP+/r1Y+F9Sz7Eq/QyB
PpRUeUPPK3gUuYhAWU9OcTM1HuTWZHdFcI+XSlqte9rQwfKJJxmDrgT/Q8vkS5J8
K8Cf27PYoLl4pXr7lOKV03WjitcHuQvI3gBYgrvTRZRoE7Ld0kHJ9fP173rJ8yaI
qNSuZLy/Fd19lD6o1y5w8yRaKAkVwDDySJTkj6fHrIiLfoB1bPukQFYavfXF/oUK
SVxEOmKMGlITuEV4fQMOslyCXdNjSd5mzIHfobctWUT2Qld+PHtjQdrk3ABwo9+d
dQvj3kuKhV464XHlSRF3tj+rJ6HLevoKVYuCG/X9l37w9n3WDoZx5OlIyiQIlFqo
Ddb+ddi/MCCpfk7Mb5X/Kt9eoEakMlPuDiuGV2jApXpFCQ6QURzaGuoFqol6I/q+
Aka7BGFpkYFeCXMNDRsdHAz/ywM7HjjADwFEODs3FFCifHkyfIf4EgOkWNd+hIMx
SwRnaslEzLQD5thW9nOhb5NfplgbwVXDstMcXdATqIqMxPDkM5B95Bd0p4pE52io
5PwlZ2bKMhiZk2GNmTxOeIfDmMuTwXQwjaemnEuliP8vIEw8s4Gs6O35UgZm92Kk
PIifB+pLfns8msnPhZkKi3ZQ9BIi2zWZ30lb2xypoDnmVgmZjTpaQihMA0QNXyfL
2CZ9Wv42Gs97DNjybbW9XQAyjep7kbxIgORIaVpTapiQ1P00lqUf521vSL5/Vioh
1JgwdsbQDCqILMnxK+Dvdk1kWsozMVbk9x8L15tL/8+dMXV7zXbgIbYZr3e70FK/
v4nXjyon3rAJBcKdY1pibrzBsfT5pNUcNLYxKCdimAsnujUyRe9OzZo4vcgxsejW
QRjLvs6QBcd8AHqVyNFh51I1gRqvzyFnasE6R7MjfMzRjv5yh1Q+C2soYIWVjcFk
CAbgCHVaCZ2tF36XVVMLA2Khwwhm52ESqGwarikU1YAvMzGG2dv8PEAwjswl4MG0
cqCmV4Krffqd2dYV6nFWgI7W43Nd3iLZzHWbqPLCJ5U/+EoAOzUiizyVHXt1rRZG
ULJGFFG9/J2BypjCh3YAWy/Ssm4iZnHDSfPJ+qw1dPLOGpWYGHo8yPcH1QGA1ZEW
yl1pV67FRBfPdrRCzDsruB8mQixGCdHevpnwt55LeXQD23My27BzRW/OJ9H8T1w3
BmHR5oxoParPJUMaQlXHjcFkrHSX5uvet4HArX4Wd86kJFv+f0AgtCM7Yg/vjOLp
wOhXDtZJK/gTQNTqg+Ng3kBSTXWlcjWrbEgwc2OGVyhzWlWYup53r56zQ6vRkc+w
/t7aBWEmXG9SWSqwSEGqYUny6kmbGzXTsEf2pNWD/3N8tgVTiunUC/ymDXs17xb/
yntZ7ce49lCz3oNkcZDxF4LCaoGx0gY5vskbFa2+gFSnuPClhW8Tul2vSabSgst1
gHXqLbFHTuKwMvfy6vPQpC7LaJa8W70hZaNyx91i2Wn1930B3lQyu6Lii6bD80/I
ok6p+ZFTjvAdmYBzBcd57t31qi9HRpsfHKFJbfleM7ya5bhelxpdMgLjEbExAtKB
BcaqjQOAt8lPUAXKX8z5QV74Sm71+kZYiAL2fV9RuGRMsJCFt8ysfbj6sv8kSedI
EvT2uRtFEwJ8+wem9nFJqeX5Q+OFJL1Rg6lS0QLTKD04lCjw+Lv4Wc7NEeBsx7z5
KbcSvNDbd1UTuEiMFRLJOoZWtlkW5qyeMpWrktoJ66eZ02fIf5QMuBtS/r/50onQ
YEMDTYVWyOCbq2q2Tz5KhYyJS0KxDxPUK8WwFk3dh5sDbDTTY7NoL3NayNEz3SdS
zaJwVwHfPeHfUwnQYSAmQeN+nOnhQ2ZsrGQbA7mKvCJDYEPgUnG/huyaqQ4aDh+g
qK9TiLllz6Gfm9jYBXMSVBne4dUYu/IQDsEpYuPl8Pj4xb4gUN6U3G//6BRdBZpi
vOdvpEGUegS2eybxNNRzKmUjaj21XHnQ1o1LiB9B0lc2llhnaQCvsuLke98GdUAi
Xn08Ue9Cvzw5TQ3Pi7UVNMLA8CHNDFElW3gComyhjw/cK9iIOjrLbd+glAmykIQg
or1E3tKtUBodOitb8O1t3P/60zZkfoWsJh6TP/z3vZztSQh2kERDbMs3kzsMnSha
mu4mR9X6kN/H+tvCkZtBWcPsrvmipZsMgrT13SZr89h/dWTyrkKhgDFGelwGQadM
o3yg+SLErr7joQ06b2upjqiJALom9ANfaHeDAmIa+WDZs7tWiYG6Dc3AnMAsq7uL
z2Fhw5rKclzZpHYk8msrKNwaP36Zm4A8vjDKAezxPuP4E2ZRKlssiuzfHoDpGEV5
i5qbVLy2BacZNnsEcQMs5Iwkezb7/cxrxRCs2mVhg5mXdxFZF+crSyUtseqnjuIR
KfqQlnMhaGe58EC3dxcd7ZXgC7kba8gDiGMBFcuF715nAT/6Fd25c8UVhW02lR+n
w84k+12JF1hM4fHD7ox3bRmcyKBhpRO9r9gBYAGfBT7cq7hQc6tdzUOcz10ZwGFd
bnMFTgZKKE1s9A2jaXQdPE1XjIYZXY5JGpSO5xPvTIIj2F5prRPOVurxmiN0JnA6
X3moNC3zE8gaJLqRdntag11WXi2UcoGHwMzk/zSX+tp+b4R0VZpmv7OKckf/xvsA
Y6obTyaTWe8+K1KwjMh/Bpowv6CL79V6txqa1PEk2eh3jl48Eub+gfE5tUDHzL6v
3GY45+rzPPRF+w+y2gMEaLFTCr5jzdUGAOxJ0LPvPlpxfhPyN2u8lKOJCq+LrArz
almWFzu4SZ59bW5xKh6Wwm4IZMBTBxX0eSnBEw5yPRQ0ULWSB/14xLqPqvx+1L3H
MuTKGd0vhvf0B0iFS27NLBHbDLPfeY/0ioWOIpcIKFch9XQZQteaUelBOit6Of+j
7JQxcVYOvN2XowF1xpAKXcZBXBMoOolYVpD3jRjgs45TRtqpClD0fC/cC3Rr2EIz
ZY+CURmXyCrtjsweQpVr5Am3YH6dJA35fV/iPOTStiMDDCF6l+XMnpKW5xBTtodh
Q8s6e3xOi4xsMJRE4vsUmwrMmlbGYR715DR+ibYVfclXEO/hTy8sy7m/pBIi1CdQ
y1WivzXdbN7THtWQWXeez2XEgllJJXYJuecYoVrvfUWch/WVUPRtT54T4PNkO2AY
if2tA3QXw1RpMWnroT6WQIRAtwVVWAQ0EMmQqvyUA8q+HbGZVeV6ntYp/k/DNEVr
MrkYJ94iR6F0+jY36YgqtcCnmBNvu1BnvGB1oYTrnCrAshXnpZHkfRaTlbRJ8rBL
NHyvUl7EqmO6tqu+V5ikJscOSZ+b5Hj1w/za5UQz8rmWE/71FwbdRLOd3fhZbk9a
68/gSN0KB/AGvuHXmQ4XXegZCigC7xMp+i/qZt/dDsimqvNgHnZQF254y9/bXyxa
9beVdMVzhacnru2uzvzMCyLPCuJC2x48iSDFSSerrxwTjmReYuSBAqVFE0+izDpb
lFQOMcylGywz/lbpOkuVwZwFPJfDCloCGAr4F4aE+nG1D3kJ7DRsaR6hIx7hsG4K
fnMheW5hOYV/rUQTt7QNwe6zReSR/nmduLAUQDlJEsJlSm6B/Muf6eCLsQbxAehZ
0gygUkjCV8zmIjrefACskXjJyx6LM71hInq18b9N26yzzev37r8Vz025RD5PXH5O
16Lb4UydkAjDsBAsj7CPkyNgvV16upoYlBEmTLH5iPn8a1P944bpp5rL4M7czFGn
yt01ybiOSnP/jhjT/VmEsD+LaN0u50tKINvdVd68iYwzG7dYoBc+BcWDE26RH8Q9
mJ0Kkil6YKuznCTNRGc5imFWLevG2ovhEJ/LoSa6FwU59226cD6yEpVxvk3xW1OK
wl418TSMickax0ZHKWEXhDpBixIg4JLfKB1nTpUGPOr5WpqjS3pV4VjFZvU4Uh7q
6RGRVtxT6Ug1QUEFSQeYnzVXwG4GbeCEHYMac5wy7usgB+mD7fWIF7kpiEgE1j0m
tl9DxkGt9yk7qHn4rkvo0XhKYyDWEUq/SC+MbFHf1KSNQeYyQ1z2kLffflHh4iod
OVHENQxPjr8ydQ6k0qlXoO3g9UTOjDuq3gbKRZLf/DINt+pFZMzTa+i/RiHfd0g5
WLUJHSpH4sFZuytT3p++D8nFbWJf4PhA8JtlXTSoLoS86Q6AKS+cxmWVXxmQ0Rfc
2aFfHFCv9rOLATt2jar6UzxUtFADDqkuXUqeTn2zROA6pERNFBvqovaUwDcS+jvG
TmzzFg10z2OUkSxWFfjfpSfVaR56gHhXY+s4qFs1srq36jmeFxHYLTjLzm6x4xau
pq7ne/DP4BwGzEsEN0GV05sWDkm6J5ewG0RdWRTj3JlAeVRgZX7zjCl1+SsgSDrG
fxKcmPAcUB15Yn2QVtpP9yGmDdx71bY4UBRPoYUSDcQBZ+W1SadnAhD8ManNiI3f
oEwXnpkljoNLP23evxONsdRkNaeN9fbYoQRncHFkrwq7E+bU/g5a4TckVZPPXCGw
guBp9zOJMRya39SC6xFJakfI3qpJ2T+J2QWLLUtUbrBOVUaLnXyHvGib17Y3h4Zm
t6OnxefU2hj17aLnk5xZmi0Bbaxk/5ltYUqxq0cosiQl8o+ufi3MsYmzhkyrSKET
mLmEqfnTzeUNaiMJHECk06THMEEI3hHKWCXNTSfh+jcRpQlIiCdpmaw5SPfYXYMs
1zqIiimsh+xfZd6vVUZC0/RYH8cN8p5lD9uXuHoM4xgxWiAICK5c64fxWwNxN9sr
IWOS5NdvGit1ZvKmJLrduIuNdK8argSDimknHOtfU8ptfKWMLK3TIMLmt3vSw113
x33bICh9CoRmvA/ymn9q06LijnMog6QL5zwFB2dH4aRPTFYgIMfDbSJfGgTiLqNZ
4IAImm8PYp3f/QEdrQq8riZMJ73HXrABhn0Tw0bZ8jU54GQ9UwEo1BecvAKLeMh/
wNB43B2kV25NudZwP8dPPBJSvmIu1reyflsDd2zgFcyEvoIyg/wuCaDEiND0FjQv
ZxnGKipIfZ6J9qbwlkkaaX5SYsRaHzTiavB2gUhj/IIVa5sLUQAfg3MfmNSGMYVw
GP2j1AphXNGCywx3j2UgyYq0g5Nz4mJIYpMKk+m6dP2tf/xhMJqApdmXJNd68pzF
TdhKUldHnB8EYloWi87Yarcr+G5kFdjnvv2AF2Gey2JyP/TguHLpj0z80qPiXmrY
VILkq+QlNS21EgAchdiUVZFjQEngaXyDzeB4bF4u5B6rU58VAwd9JuTK6Q7Wb5tW
ePHt6is2xyoYOdMyyhlyvZg9wpT2aVfYP5WAJlUDLF/inHJ0xZa+NYCvVm1eJ5RY
BXw5izyrZzN6Qavs7FGEfnTCTkjB85AehYOuDGsz0C30pOUeCrg7LxgZl4NTwQXS
Dza4ORx6uyBs4UURdrNEmJti6HSb/kE4zMQ6MRZVhHgtkwJexcHKizKCwPUF7kO0
jKSslAlpJr30l1gb5g9qIWXQRYkb5H4Y7+RihtmBYeGDDqlv2fySZCU7QvjVuQPI
kOHgT1G7da9M+46/DuiZ8p2Rjtt9IC25ozwsiMsO4VRtwbLIlVZadSlsDD7WpRP9
Mdyz7yUbHG5XAZNmD0bbszIN9a0ArvlsTMRWigXb9geCfMsdGzJZvtzjjVN4dhFA
P4v171Yn0kDCsWGs0Gh+OrZOU0eI+IdeCvL84DYf7Y0rybfyeBQRFPjv02oG4kbI
smZA7W2lkiAPV84H6aD+thn86VdvP/rvXjhrOdyO+9bS91NcsVoJtG5ypVsroUu9
gSOJT1Bv4+cdweNC+05GQj4tfAlD8cfZ+3M0mmE5rG2cIO2GOQ7f9fP5XtyO2Iwu
q0niVruPTKS0UNZoHwtd5yE4CBZlhw9cWR30o5oH5ge54ZwhuVcO6A4HvqVcImb9
M8aQjzas+0aUn9eMlGc9SsxUWX/EtmS/c0ITx1N3XKUH3+SSW1TK332KZHTfoBvg
DTFFNzh8gq4puGkBcY4x9ygCJDbripcz2OVXwyEvCRL4NoX33QaaVaUbdPwuR2NV
Wa+gEp2yHPSRUZrGnJ8wi8IR4VV6z6CNiIWdQ/TuqyQcYlhmqbz1u/TGDjM3MjLq
W/ldg0OckbBsnyyv4J17NkSNZMpFApYFPVDjgpQE7BvGG/ucDkLUmbW9Ckgkspqq
fd6JN3RjgnU0CVi/2RX6x91bcjpSeoR0mfsI8x+8LI5M2omPUD99kezHI1md3JTW
p3ZEvHqDuvGl7r2zfg64GG0dWn3mThhhYJYpKWSx5kSrJ7im96jJ7ighkQxHYeW0
+IUNrzlhzkROeWlt9CiuIKEt0TaYTZaFK4CV2Y+AnsyXAPhnSbij7StEygBQYZxg
jbujh75Xnc5kLfSE6lDV6tgoUwLUeCzGECMEcX4+Z9GO9dpBG0xIWB3q8704ybqz
+hkBzfU331dUhqCtrzyPGUW/9DXGSHWZpvtcsur/dGVAIF98rjgcxdmvWoTyTHHZ
Z3nqPUWlIgUMErBebBeYiK6YESKinpB2SOjf0oJaAmjtzl5D4yKbDZ4QMFswfxF8
urx69sgB8s2Q7q8nJya87Boysx/wdf1If06WIaT18SNpRk9nto//Zo8pOG5ff+3p
zF9urAXLmp5ESnCVRH9+bMyIqpFtNAR5Mlng46cqIqXBynQ5A2RwykfL5Nrp+fin
bfxVLe2pmdrykzNeWWBYeCS09napjOvFcMyhDCa8WjSZMl5sEHIBIrdUVZ7ZW+wR
QQDX7RUd7ZHQR0gP3OR6FpS+mRoa5tt1XHCLzNUOqPXwmeiBXbVl4b95oi4f/FCG
gVYltGLen/nyc/RXG5wAnpKAoR6RLyh3XOtCEyGj7GbIo3O1jpdRqowsaVBohgHg
9815POIu8TSidfAw82D12OTzITczoajzGXDCsjhPYQFXXP1696Xvcwm10FlSMNNG
Juz0UubswCkxeYnfTIUTmGmqHyj7b1SVnvyUy+9znT8O3vGqEILmMr4qu2Diy899
1FUe/xXg7bNmktqx4QCEPt2zc9Fvy/JatP9xS1YcUVbPgpTE/79Ik5Izlu/x9HHn
mY2pJLp1ySUzLB/eh7WHj/W/BdRVtIPBss2HC9x99P+LJAVJiRPnMJpkcusmgbzO
7nKCcVYhJhO6Onzxqm9GAVXLQMGfishhYOTOTxF1BKcHsonzsvCd0AiE10fpTi+f
tP51PJVj5xNoGKMGllGLuheigCxfGO3hP4I3dh/PBhxuJlaPdVEG3RJ6w2e2GzEL
FIjmMkkmx4dsZMz52x/LzPeUMb46KnValXleMamUdUKGlg1jWrgeG6mkG1dyao/M
V0Cpz4f/c6IRTFYaKet5m4xCNneIfEQkkqPxK6QOaMw5SDi6OLF6aj6YMiWJ708I
jywBjKf4L9/yFRDt0kRtz2u2sckshTYsCXEj8qJAAAt3FJFr1CfY8e7WT3i/0Lgr
jEBqOUFC3Do5NbjPBFTGKHcRL25sABu99y9MDJZZ9U0MIVgehT6OrnCEdBxO9AMb
HI6EjggU9uwofvByePe4pAPa/9joga/mQL+LMUC4Ht9q1wltTlrzMckRlY+Ea5py
2t3iOarHU+02EwmP1H6eUuOUywLyE4FWNO8savC8xQCyDpOQrWsNfV7/pV+zLC6i
yajdbEzwwd1f+LYnorKRYlDwnXYSWiIosYkyKB0wRnsYLYIa0RFDZURnhnkUmt4s
MXXkqz+LHMnyfH2vA4WmVugoSyKcSpWgBBcLEYk4J9g2mxFFcOU4KPDgb2nW3jLX
txV7eltAfNN9ZKuLBHN38s7Q58sGLl3OUhcP2DbXPdUcPZ7ngt5Mqu8KiGbZs7mE
pzIy9whELav35EbFO/ue+dH9WJI+u1ogdifMsSu6FV1IpLx+eRnJPyYqOFUH8K9g
Hr1Vv9Q4XToPtOPh88Y9Gkm/rXpJmJNgQ7/XH2/jduQHK8wYIWJxwQVwOkxarSSk
SvnY6clARZB/ksiWE+s5QPYx8GZ/2Z3qdBW6SgKombzKq1rCvS2VJDJJY7cudBt5
wLNITmKfDgRBI+0eyVqjaAckI7JMUpr4CZRH+nFG3nA0NrAZKhPHBOB5SF8gm/ib
p5oh1HnqakWPEYQ53HtflVZW2EHVndPcdl+A9wMicJiW5HQZ0HSHJ5DDiIQ9Axk/
2f6pZWmeNFj0nlwi3r267TuXrGXkgkpMOoZHqXSqIIRifNCLDKpWaREY/CkvtgZK
QVCRH+oRBoON6rPCzrHDyOqMiQLJ+oL973WocLCe1vXGse2CrXixk0EsqCwceZ/b
TOKJuSVIwKAj7KnO6eZWKmmZP0dgBWyWPdLUCAQUTCVTvBC+r02NyTHbMhqPFvu9
f+42bjdZ8j0lx3PVLAygUktbJtVGO4MoVdB5I4SEukSe8Tz56DdWDIiy9meOjnNs
5nws9hCJt2JHnoKroyeN2ZOxhzHS/3PZpTstmnqWu7E4cDVE2ZkCsnS1UqWS5vza
W84RqJLPg4o1VUK+ktuoS0aLpsw0bXm7qO7sA38Lqrqe+aSN6eyTMMTd6kIMV1wE
DVLYs1aAtOopFWoUsO5Flb7i9ppdLAkVjMnE31UhRslDz/qp9UVQCL9ZksfvzmD0
w1EyvJPjCvA44Gorwqi2IuA7z1bvNTWA67MFdq4M/FoCs8sVfqZ5310lFZ/O/o5T
biZEkobgoFERUEsNd0TWmOUHVrrys8j4jfT0DQuOOVBmhIYa/Jyp9D2Dsv5qdIuC
h3lnqLOIeVlgNp+47obMjIMcaOJ3O1Pctx1TobNoEYnWpDGjiHXOg0RRqSt+bZB2
IiaGUnV2flh3eQGXXSy6ZKipLD8qNDDL0esN8CySo9ZbByz19oarfRfjfWMcpbHD
8oaINeJoHHUjV2C9kcOtelJ0xBLl6kM+vrm/ZituW+Ln6kFUdwhMrrY+UL160hd+
tCK/t/pps0v6hLwKCxqEv5fTHYfJnFqpZ/sqQ4W11I+xwKXdyI9oz9DYJK9L7rSN
qTiJ4jBP2O288QFZ2UiCIlpeoSPaFwgUbxFaFefQEuBZpiN9ytY6uQALiTSO9ZTF
iAna6Xwss3HzF8XK2K/f3ZL2V3HEU7lZrlVKrAhenRIv0tg8uK5xiLj9rul8zOqp
2iDQSkEoiz6k1cNgk1Qe6cc9WHkvdIysN5g/XG8Vgg0B10qVBvYTHUejJVaQqJm/
Gv/hwOfF4/rFkOPRTSCNmv11NOSPs3IVB6ZXJmdRw3yUpe4sk0AwKrl6Mh4VYQR1
PMSBG0W9woRYjCnVht/WrSwJzhOiLkvFz3gvu9YcW9GNWNRGpPlABDJEOMr8GAov
mivOKMeVAH5FcSDtF3uujrSsCHUry82qLL5h48wB5z7QHCLOH8JpRMhof1fEkyI5
T9QJzgcxVFD9OhjavyKZvoWgWCqaEFNKbPr0zmTCLwXfwXc6J9D5ZhRXfoyt3goV
lOuaookn/QpJyR3o128I6h3M9in+J2/vstLZ3ayvy809/Y4b2OcaJYTdMj6WuLHk
J416QG1+B585MmAjwqUEU/kHBXX6WwsM5HotdQb7VA61+EZm0+aJkOz/Y0NL4UaP
6MVSGgoObhrUQeqLSz/QURoWL71TnFUyhiwxEmo7H4fqHbpu4lQ1zho8tU7qyR70
oYvJaQewn3X1JJD3PuVywvqfhZ/wqZlbMfQ5+cChyf0VsA/Id3SPh5csTCJJWi0q
azZATCDvijieTsSdJSmPb9wrVXd33hHxC51VjjOo1ejnPPMz1AkdA0lRlDAIhx3S
GxHD07FNwIiyzKnZvYCPGZ/mmuDBFEX5EKoA0FkBIHUGWsBuhdVuhGxtllaYX7Du
Z7I920ZH8F/ILAYbMr7ExiYeHwFX5M07qzABbF5xTVt78b+vyoC/4iE0O4ow4xhz
mxCOiB77ciUpSGUABtnLDwVwUeaWkX9yho2ldoDH2hFrcKCfVCj9lZCwubK45ZpP
BgB1lHM+AKXWZkfPurgbykRWC5kXcmw3gSYQLBAx8HSxLtnhNCfUHnzUx8VwMHhb
S7y+GwJbbnu+ZjXALoPvdZv1HcWuHyWhkrRR0oiO+6e6qyioib76Z71Y5fvTLMRK
5JMwDbNewMcEsxIuDHs/AqSdbf8LPR2rH02m4r6QKnK2dDZaKzJj2hfhhwk4FCXZ
7uOc+4x7g84Rei8mb/O08HSqg8alAgk+/bA/5tASyTu9AaHsHrGy7hKxvwg3bDc3
FSnsQMP3xYrbyvfbfl2NVWAvM4Gw7TcwL6ur8E0hnwnrQPeimI8exXltFpNP+sXP
rbu4XES/6tsHj59vcI4NqHVGp5ENI3FcFArFDRnDl1L+rMDWG77ZCgalVqxrN2d8
6C7Z2kOtGtHzG0Y0yXkklEhRL3S5aftAHxJH2/RqBUQdBxQ/XJYQZN/+nyEaeGJR
nm7VhDWXidFWk9Q3MTNpRwm6iYAC/e78/gtF1Hne4aC4LthOHioV13prt65BAAbM
W+bcl0wCU92YI5YSo4kak6B0ChgbhO/Ef45lEyo+rnrKC9a7YkHmQ//PTFQisc1i
yfP7ce9iUwpR1MUdliELrhTQx22YCO9J0pCDQe2Hh3T3utxONCWQWZtQywJyFaX4
jjXbXLbkQPZ4FYT9w8WS3fHoQd6IeXPnTL1VPKl8Ppj7nP1lObzq8sR0ite888/L
HEjFcCYsfcuH4oaqlRdikFtw74u6l0fhJxNDVpY/8Quu1tGcPFfLoL+hxDZhHOcb
Jolpt6kTsWSvPYSaZGhy/+61B7JZF6aUME5aDSThxT8LFx+6mfIyOumUaFdHfVuR
21TAgZpuqPJdFnv1tnUCDwAtCRDqranVVO9SXpOYZyV83ftFJyB2jRiVO8Z2uBmx
G0DG8cpdUeWdtSt97EYNyZ6ZRpIFs6r0b4afURJEBQ9wy3rznoP2LsBdkT1DmYuJ
w1IleQ9QXDwN3XfHI9EdNRcgC88S9ocbc1e2W+AOkpujP/JddRcEWaihHfuBeLIJ
c+dye/S6HrIjWl7Iai4+cAaieBP0krFmLmZQoXnhfuz373n3mEcqoNulVoBYc2R6
jXrcUI49y5tw7F3His9E7+r1bz8obNCp7jdMrmW03JD8Gg7nsM3ni+XYg6Q1RzV7
t4R43qU3NwayFSOqzc1mtW3+vhe/XnYg43xNWv4rtUkFc9VDga1r0Q26D+NQMaxd
ue+imG+zMLRiGl7KVFxpMyKPOlf4oRPMvEPFqhQiBd49njeNFSmxu/otESCl0fA2
/SAOeNp/0agsmrv5dBQKrdJY5Rlu7DTfSj8RsHzcbm8MN+F/MIGVCYyTCbNXkT7g
mi+tVUDqoqBUyFfmZbnJqyj2V35xdnocoEQu7sVapx//yb6ZkLYEUuz85wi0YyFV
z2lH9C3GJTvdwr8s6lnW86bR7qb3KEBZNygOVDv+I3yftyEK3piGHBi4NxcirrXz
7VuW020wfMaVQzjUVdKRa4+Y729jpQjV+c1MFB0KGN1MlNmHQwXiaeFdAlwypr7N
PZbfWXKrdQfkj0BS35ErCRwRjNcr61iwnRzlBv86g2GXykKCj8iL7DdqO8skiP2T
rF9oPWTAbIlvfGu5OsCrXu4s3BJwH2u3U7q9Cu+xqc0CjwtaNefldXuLtg7ssBls
WbdkvzuOK0cMzyMTCJaeGcebDOEHXd9anYJTfn5x7vu+RGZDT7du2/WGSx+7N1bZ
ekZlGsxEveBAeiTHFDrPkb04ud4vtE4KYZBRxjUu7a/ASL5Q+FaaUj99D7/XXjMH
OMCKtL9ebfDlWWbYtR939IpBxO8kVzcSiGllalSDNchYUt4vwFJXB8rXM0qUE/tY
1pHRLgC+fJbaA/W6bjJxxheMUFmZmeQNIqpqgER37sAKYVlkKnTgpoWE6YOkBR4G
dvQCq4e/pBWD/CR2xG54W9QtwxfsJz/MQsF+Ewbm45fKHSk3qOC6fzuoQUDdVidN
owQGtYf5lmR+0KNQ0PvCqniN4X48kdfcC6Sf/eC/HfLH9tWChnBjyMB+mqQG+FR4
JK6EZDmYnu/b6ibXsx5QXzrxicc2ZGwhhSVQ75v8njZAq9iOfw58SU9VkbYZABLi
S0wRh9kKtvQBjPsWMPtzZiaySDMLk8PLozlGn2PNZ6wOA/2wzzZRUBvSMWZcqYfk
167JUqg3eAsY3k+firmTz4UyQWtWz6Qf+U6MwbMhSKx+3l25pEDLZSIhtBy2ApiG
XAzrXN2zh6Xm1VsoldQGECcuybsXQ3QUjLGOYm0RrSpCuIOHHF95cTH/LE5HB1YJ
uy/Cr2Q6oR54tLGljuWvAk7kc32TDe4soBOI20LR84Xi4c/PqTsN3u09/UOOP/AF
B/Xi1m1g1mayklYX2jZfyX0GvLfQNDr0f9If/iBlz7gXwMKL+KN5AxrCXCuEJhWt
+OFMNlu71cKrLROLs47+hd2U7X6PWRn80jq2/8bla4YROOKYHeZpba6MxvsHs/ps
/5J+M/qwO1ZNMoZysHPbewHMO2yjy67tByRQlVxuj48E5H+AdxXIkkk53x1fPG05
AFI+0k+67afu92R8SBhZ2bORV5IZlhIl6gatlMC0GW/ehrqksA2mWQnduHY6/oj4
KVhaeu7Z0g4/8i1fCWhCIQTKgNblvQWD6LujMiORryFe9mVaPHa9qVigGY3y7Yhf
t7za3w25QIAVv+ORKvgYQFb6mIVRPUrl1b1MT4PJOuQLa6MBMHiO20xUF96gi7pW
H5ekdZM66r3szN8eCMKTYFEsCZpdrowUt55n0iQmmLqGXjyNkecciLCjGyTfIZ72
vX3XShG/kuxpgPGCCN9gY/crOQoRlrwFnezgtj+lZMQoIgqD/CxYvWZwW9SIeJf7
DShzE9mTrpDH6hFc02WqI7VvgkV+4BG6qweu8Kc+RRG+ttxr6cnqPwd1ObkWBuqP
KxEZNtNCrPDH6HEl5KnRzv44k3yu5YkEQQgzcnMvFTC1lAZwsop1e2Hk48CnFMwN
jqlR8Yz5BVf4B/3oxAw86S5MhY/fo5nTPXMaxphf5hyCjPhUtc/DLzMvc0Jke1CO
HQfhCyM8TeL0GOiC5POUKauQjEhKOZxdkYgs6g4PXIK2A2rHNP9VHsMKjySeOA0w
0A8ab/f9dvEKhqDSSuxEGqPHeCfHy8dNhuoCLcL+uHwC7Y3plV5n3afaCESfcugL
GVl0c8iuMR51vT6msGefuFRK3hS0B+VvSv1Llm3ISRCxZJaUxT+URjBF1oOpHG6i
peJ383VjwpbXqRPfOY7qYLX64LxIQppSCKmDY5I8qjwo/LE+Y7eyYSm/iKxQughd
2hf1P7nxUnIPswwBiw95lK+T92vXMF9eNmCVXpDnH48ts9h4HhPvc/Ec2k6I8stl
3O6v04+uIFZ0FblqCpa13tOrzGShQubQ++3TMH5aeeF3fMHDBZ56q+/y/MfKNt49
5wYKQ0IkqpVpZ7iHL32c32PlxyeLiQYbQiv8M+MvNad9ou9HhlzW+cLVbLd/NSbP
KLTM6u7DxcrI1fP+Rssq8aVqDA4hIcaYoVZ7CMXxMCtVz//q+HbHyTHyQ7hpUQEP
AnL8Kg52Ip+jc551k8yWiiNRZLR3XPLaqaq5aizoTLn5rb3rr1kydVI6avBdjqgD
n903wvRTgnimaoDe+V2Z/seJiCNbq4VvAhFluV3HebPxqrNctEtuElXiuIgbSaI6
eYTpkx1ftytRjtcQISiht0zpEbKxRlxVfAXmHs3d/iuwGYPWwyJU3Jzsvz4o8CgF
Dsmj2ueu0IyH9p3R7qTr+dcRLl0cyC6MG13zro/UIp5hBffDq44DvweRdo5pxRqw
AF5LbE90p5nX4KolpqG748eNcTxQ8/py2yGrosfaHliM9tmry5jJAmXSycpl2bsi
TBDqo52ki7+F1N2pHMOA4EQqo0ipZvhSyIumF7PgbgjmGIOof6xGR9oKWFcaDx74
piWVbAH9FRlc/GBmDUL1wKP+HbbY/9O0M6HbyMLNVwyUBBAhCFMLTSp/Ni6z2Wlv
bKmgHkDcsNqSWqObDZ6IpTkJhC2WPs7i1IgTyDHUOgJX1RNM1rRPGzlVzeOoIFuK
SmdVgiKjo/93M3fpAbr/WTtE0gkKbQXOpBigrwL71imNmuBPk3lEpjRG8W6MWTVK
MXcAixM+vkSZZIj+/1TaayJ0vpxwfftr8mRZVYiFRG+suaz/JpV+vYyZcotMjGPe
g/g9avwBI2qkAWCWqMyBeiy9dhu2sE9LwSl3H46Mkm+TeqNJcU+tkQNMNoMvjXMI
odW6bKNHKL3cSIc4pE/NaROP8eeyy1GVoEo0K/9FmKq66jBCqqz3EuLSjpzdmAEH
aw2W/zlbxPkyX9EmuJ4M5w3LgcEZ8UXFBx05gHgkFW4s/T648Pl94uS7SB2WcH5S
7KBGjUBZoAStm2Y2tZ7Cj/sGaz461u0JU4rxEvueSg+DnsSCNxtJ8U+p5vzvzKS9
7UrmCan8AO5CB7ItmoGqO89DGkHDI7bFh2cjsDILTNvL0+/GOe7mUy2Si45DBM4W
bgNh/zk7fTCsTDBPk0z3ArRrzczVPPV96JOytB3eN4ecmfzCGKzIj8dnz0C//Ldp
0SEEb47EU1hQIrMQ/g+MPkYcIrG7K+uUH6k1wDaiZ2HcoFr3vQR9OIann8e47t6+
ZQ51NyHxOX99DWyQNlvPFiudMhDxgHISrkdvMsBrERrZKFk3hY4ktgNdmtc75U7A
TzocAACq22GHWwQPj/6PM8z+JgOUbh3UYAOg7Y3Cs5rDYfb07UaM/DTSbjuQDuy9
tiYiDUEB3ZVDTclz1tOCEMml4F51+kf0eDx3VIlFgmmUB+kbh34pfWVwSQ8WlXmr
q047g/se1JYVpB/sa7iw0VwqeXydE0MhH2rDgatpqaICg3+nRXxOGKeWzH9YzVsu
VDS+LbXBFt+dv2yc3k8MX4XBilTBCJvCSrhcqtgLX5krNtOZVsR1EX19buJhzugC
PS9KR6ZK0dcB17q3oEy9zjiG95N2Dm8XEOekdIbD8gj6XXw01kIlDswzp+qIBmQB
sCkYrxXynGnvyNzg5RLLkP+2qrGhTBC+pc78OGigU+vByv8rcGAau62o2zOqHma5
03PrIVFMQ+e9MT2K9dCPbfeGgYhfYUpPLVec0BvxRgqSbnur6E1qBC3YOL86oQJ6
2HwrbBDNBAtcEAuLHGpzX/Jkofu2WsJCh2yUhnx0xSiNNFGSwgfpp8sKI1FRw6rG
KUq/fRS5sl7DVZIOfXcUYZm3ca9Z2UXnCRAgQ4reL6NJ0GHguQtDeNJDTbqq9fai
X/OaIk8o1BGYj8fB5m/HBGu9WbX2eBBgwBIHIevDFpPIWqPysQhIDXRMr4eyvwsN
iZv8FntJ432zHxn2ZyqEdKGPWdh64l0qfwxEzVZRVKIbM3oHxhmc8u5wyZHCbEVX
nC90JR/yAWhv0IuonisYQiJH/NREjMpHxKf/Vi2iWgULs54+ZQ8hjuZtJQYMBq7C
hiTa/RuP2O4J0Lezio9ekFJmTZRqohcZkDeUn9QISes3tqsPUOZcZY2TUnfcmwCk
Xl8iyEXcgXABlPNyn7ImGYsbp5T3hCUyVVwlw2/O1wnDLnLHmv2hdCReYUsirwgJ
v9QtEhH6nJ7eV8NxwO2qooKmOxtWGkqSwMUV4OmzI8TyXeXSul3z7zms7a2LHW48
vDl8usajvKgtP9MG5mIDQS8lZYOhB8PoIlKv7/ZtP0AtbhTn+aueMwDiQHtlWDrm
EV1zeF4E08lunb+q2QMIMOVa6OYo9XXHEQB5loLH9i7kf9drxXLYGfMMF5YKVEDZ
dwYKAM+pB8uisJ6BY7NRRwLt/Uc4r4f0SEIF6MHqFI8ep5CbVPBsj9u+uDKO9nPl
0T8FONUiVm+wrrW2YQFTxty9xKO0GCAW9JPRfx0GD1K8/OUw6A84XKdEgZvorQhL
6+zOXWywb47dF5eYUJGJeA+qiOeTbliehCVwz5G1KzUjM3HkD7kHGbMAYjxJ63pJ
4zpmnMdjiga8P/Xu/YnrzWQaF0BpvV28uLBjDx0hfs0BPwSs9GCp2F3Q48kaX2EX
tQIpSydJ8IdC6BIse6HJiFP9ME5nb+FR2DwwbWluFESIX1msQHgxyjYj4Hc5NeTh
vUM6AseyzW9do2BHiirdDDSpnytHb6FT1QZcRtg0hAjpm5ofAO9RP7TFNnQBri47
porCd1lpkW59H+BTG6ec2Z9irEap29JiQPbNbeDe8suPzD9W7/8vfg2hy6hnfEdt
yU82tyRd/vUO8DlnjnKELwODFCzEYQnXDG0HEtPY1g7SCbC7XudUtq959w1+lTNC
BhVH649kfDCBcrJ6/e4/lM1Xieg/N3pd1EcNNqeD5+OeuH5QhfO4sE9fHJ55daLn
yKd1yJ3jr9aqy0wXElFOLsDkh2Y/+kCMljK+AxWpjW95RWlLRYRC+Ivo3Rr588xg
SUpz9o5y2u2dbgY9cMRdGSyRoj6XrhMVRd4FTC+183ZH0opfbnGQkCDxAPK0MHSl
EyNuW4Lf0aEM9xeiNME56N9lvVG1VNoNz8Tgugr2V+sG5Ei9WzjDfqR85oTPxY05
T70xJ6YbCmUjuKanTpt1L7gfknQhGImp1/0MhjBuR0vLHfjD0oKQJsUL/ZaACGxn
Aqoxvl4zNg6jxflMIOzOfXIU32lvpz+m0kyCwWjOBpJpxMoLhVmx+d3bDWe08cfG
Eqkm0aFRS4/S5muP6r1N1rCJblSMbg0eOasB3dy9KzpMgfsnZi87Ng4ehad4ECB2
dLXraQ0n4pNVeydNq5087SWGhZGjG8+gVBahpEF17c0ObUEm4Zyz9HmZOKTgOK2H
GQS9TFk5nmLXoomFtzlfnG7o6SWylPYYdLpcJrf+CYDY384h0YLCLPzqNAtJNUU8
CiLIGgxlhCfyEWrD3jELS9ww8LqZugwn5ScXkE8BCm/EGOu2m8sQ1tnxiut5GTKr
bmZaHeARIcyb9ReTwiA14erQIfJuhjWPB1CDjr/yyNut9Ju2TKsOLnzAAensT6xu
Eqilvgil3+6xI/76nomBjmIaAq0YqCWzg+PDVzCdifLBeE7934bxVsp/qIxgCq31
3u92JGcP3wE/ia9O1TvUk2Tdr+sqqc5qI82GVwwv199AxccVYc+FMxVzRZKHMAcW
8isFX+0neATU+TlY5Qr6HsfZwAAZiB3kknTqVAGk7TWQUm+QeAlN3lu8nVugiMsU
aj2c1J94wLaJR3sfTYpS0rwIb53qEPg9MYfmSHMhNUQe+HqHWuVu0JLmbRWls3P4
2eGkgA9Q9T9NugHWllqGtlmN3qK6POWxgYf6jKBaEzHZBvoNnSBPptpj7tbs09jp
jkOoH6si7nJcattIUVZK+YnvJ82/2e72ez64XNt2I7TD7MazASmGsqUMsRT7noCz
Z0WzSz72BwNcTAxmX9HhIdUm69+R4q1j1ZLXx74myZqB2uGCTTojoAo1Rk3ECnuX
a/bvvds/mFkvOoVnleE20KnVtZn1hUZ10ozOhu+UfAIPy3zxrZCNvP/pQtlJfPmF
hDq8dPp+9g5yMWHh1zwZywUA8sDmSzSULXo1q1kultz/XuUGGaHDBUKk6sU+m7mR
Iv0DeuLkaQTKfNHIjJ01JMgecgMHvc7WgQHG40kl7QwRoQXlFw2OTW8LFtuoCNtD
+5uHKmN1LoWeC5CqlsWYHCS4mGr0W9sn1q+deiO+eQJgi17ACi/eh8ZcW7DKQi7p
IEKBUB0K6Y0AYvXAiHSqJd7XU9LJlG9IFWdl6QYWPF2KW+amcaKSrmm0e6f0pCcB
o/39SpezeyWXKisHVR/QnRpAri/9c3T6fwgqKQ6ZuQnEuXdyl3M6+HyaFhgfbKXR
AjjeyLilhSmxsGu5nt4Cy367D+cuCRYvaDCPKs4yVAis87LI9XCBM1VqlGiyJqJ+
3mOLArQy2Lg2cft2L6FVsDwtMazVh07cv4cRjMop+O2sy+BbCyGN45+CSyQ5hI1s
eOxSSeatb/AOWcucu9Bd0jueWH/aCti8g5sXeA0xOxpb/1wSnGkj1F374eSOZWLg
nucoqnwZFBusoZDX6NTBdr5QwtNt01NveuxqoZ4S6K8Dq7EQkU2vMN0GFkr/4uBI
CPt7+Hu5fBaQqg4cmIcP+Mp1r4rkDhEOFxGd1OD0r5Uwa17+FFvRWBk1/8vpZATh
JFA8iBvEZXdhsx4ycIWz8jyR7WKR4lnchRkuqjh0L1+mXXQajDGzxXrVn+47sLux
s0767PunGrb3sOkfJrEsSrSDpIpRx/z/AxBl7Z9JBZeIKi18NyAU2eVhS1VlalIx
r/48Y+Y4JkjN2dUG5h4dfo072QBN/LsPGRRByQPY9LAb8+Y7KzoJHR3N96+kuSWK
yp+R5FVWLIkfXy4e/l0ZOXfxPp2LCXwClD6399QG7nyR6AM1g+oHfbMUnHjyinrz
gDJY88cn6IEzaxffEBkHz3/mktp6IlxYjAZ8VKJQXwXN4aGF3orHt6oTaqbmgzZT
0inNSDmRM6pYouJ7vd8bG6KWw80GzNvgKg7ooRfqVOwyp6d2wckJETvRmHbVouQc
lZuKst9aV3rnDdfVLm+4A7jbHuCHk1IMZuGPp28wy0TbhKPfkU1CM/vQvxQcoaEp
BPLwyu1qgy+NascjVJgDKFJqyfCqVrwiYa7WrL2apNUVl7nAGcZtL6Zvg9eYa+vN
u5GXUdP37grn/bw2F+M+ccw2T2imu+p9rueLNjs/ARMsw/FgAVNT0K349lB0+G0h
0MUUisFHadYdWekCuGhV751QGkGIJ0qJQ9ALJkxXRLfE9utbwZeTLsjFpHGGA4hE
GqTpoG115uFqMqxlR/4iKYGyIz4qdT7OcB9FeJtBNX1xK7axDob2WqLogbx1S6Du
xF6ZH7uMI1oyO2gapOnPnJAyQixBfLLNm9g7AqrkBraiOWp0dk+XGcsr0DiDHhB6
dg8i18Y2fB8XN7aFgzZcRQCNaBH/+UPaChr/62HZmz//uHa8KOpVbW/K0ofXrwqQ
+TBBCD4pu1qr5uAqDmTEH9PmUfHily9oz5YQtWtnAKZLXqryki7LJB9VGxxvFND+
6OSu4qfZ8HMVES5Zp2jaCZwiGmLpuiU5XzPhig6IyunOSr2GX25OYSneL5UeseKi
RJHoXbkkf8ZQfzM8iT3zLJviDbEuE1mwrNVdCo0F4EleU18WDeszDJWcopuv+9RI
5xJJyYaxq2riE7cTIUywRVX94fDlckUa90Wf35zrcY4uDI4VNzwXnk9yl5Z8M1/b
OWaIB2qZslI8OVDhq8cCg/q0Frwr0ESjrAnXz4gjQg9Z1GPLacrvK4gPJx/kq49N
3KNoILn+YAYSQWmIBd2zqgfPCJByTcl+qPjdVLj9fdNeyTwOqGxfPcQsOWhsbIHf
eeoaEiizwtAMFUf4E4BBiTsxgqLQa5heeaKNgIFaxT7wTldgQAKHZqoJh76r1xcS
DQN15Fvn3Y7zZbBIpk96jSNAzVR7F+aK+NTafWte6oP+abD/YLM2ChMmpyxwI9e7
UEIP5NCp8N5fAvGDQ7f8TaCutFI1rDFWcSQD8ESqmwuzKhQApN4t3mfHYim5Njdm
czzyHh2qjgAP5ZBBDqAcxD0vIE2+PGOFokd6XYWraXKNRiPpgDFJG5PdPru9ZBQr
1nYGTUUn7zERqowpzOwp2kRQ58W/rdz2ifvHmEyOZfC8g2/t+1jqfnv/Co32alNe
vDz73U6UfpNgKmrnUsvBBZzo7nFtHjWa5k3N0c2291vhz4TsqJQdYNn/XnZFaI9X
FpoiGkSPGWSXQ+vxgz4szCWij2lEu6Ys6QKqQiMryhzNCkfsN+T8D9aeMKx2Trxn
TCjQT12DFDamLqTdqZaQ6teHBlhwkD0MygU3OpS4w9mz7ebaiI51c1+8dOSMDVmD
p8ROFwct82SBNwB6/4FGxW48z2IiJ+2suPAfa7avD2BCpZ05s11w/wK8D0CsSMMq
mw4TnbyCbLCqEBpOyQPKOOoBBghCDIMMXXaHcr1Um7CzJusIJBQDA3s1Nr7ArlaH
mcPlcMo/bwU3SHzRujTOuakTevUwj4qmkJK9AqQ0do8ac4nKaB775FBDoG2Be56q
igxZrZGB2ToDI3LyYC9uNKK/KlQ4u9n6wJg7j3SimIFs43cVY++SSm5eNFilg40G
5lBD3I00/WAwWE2AsKFATOa5DchIVLAebkT9pklRDdDZ31GWpxgTsnUHKCDzAjtr
fT7hOZyur9tptsyaPQiLt00s0x6fNT1jdk2pLNiHeJQcYxvSr2feetPJ8/Iq7oCD
X59jH8GHo/xAEeAMG02CtIhu+PUWeKFwzPYLPUcln1Z1WvQ8B04Dr0uOdF5NHgfh
s2wlMicveVr61AQnawace5efJdEkxHAL5Gc3kDjX1yf07tVpYYpeo5ILlLheWmHw
Fm+bYOWwT2cNCn1dVdeh2G1+qMFWad8OF6rw0TQwIzfG2+gn13oyiB/hmpnN6eat
H8Ab8dLXVbxhZ4IWLZgANyiI5G/DO4LYaLC3P48gLWNKD/mdW4EmPkiaTq6VQ1Do
WiiXD6LMl/mWYQlECGd11OAcBuVJMaQPJ+4Plo+KrW3SWng6qsf1wnRBYtsG6Suk
uJlDvu5m/5al7WvsNLCcXBmyp7qVqttZZHN5+nXH9wbUMnsmVGRaZfhwMx1xVRdK
CLrNE6l8DdmJwvMzFo9iRVI4W6U73GThoLoZVgxMBThOwRomdKj85nkodn1luhSt
mN4UkImpH3DLHL3xyZUZw5q3zpfvnOBHj3Wd8okkxlW0dpnSsshDxC+2O8AykF1o
nAdfiOIDQOCc1qVYjqIfvbNSWGGZGI7nGt24DIVlfzBP6EFW+schUFtlyO1Seh2h
tB1OW9duDWnmOhx4J1rXXVnCtLDHHwXCQD/Ac9NZkehuf60bKBS6xRTxDuTZ2PEi
Cez0jOPvwBhyx2UiL3oGtgKXl1jT9q7JOimmipnN20FFkzPeOXwj0PoR7ym87NXk
8SRzeFn0Zxlaw5lwLB5VHK1O4e21vtWqsjgX21AmQIX6+17ePuAiQ3KNLxPFq0se
ccvjlBH6flbL5Zl+0BdXBGFXGVcSxqPbfU9k44/sFNkDdRz5VBXXWUoIpxmJDMjX
/rYJuSujvAwtAEjAfrdFG3bHgtCfIq9Ui60dYY4ixNRRLEJ6fbouxZquCbF3Ygwc
G7bR87DOuhgdkRj+79bhs/mGzR7toNvcWm/9ImrDUhX6OVUb8L34DDlFwicfuXFP
NnDvS+bhl+KI3XlT2vODRAUZhJxfNWkt1ZcVOeNYklLw5nmctOZUWH0Aej8MERkr
m/0tuMS6FDtip+B+tIR4sxUCVUVlYhFvS+acn1F8GfsR+MFNaTmmrvuf5EdOaSZ0
WQwRFBYY1Hh71vtKQmgKIs8mVwWTORMV8PiXOxEI1gow89QOGnGWr8iotBHLxwnn
5vGKCbwd2nQk0uGO5ZhdHmsQn3oASX45nw9iPc4L6o2LBBgI211mQf5QGIQxKDxK
f7M8hytvlCpdtqjgi+NvDjjCazmMXp4s7v2VpaynTAJBgYXbYNKDLjYztJu/aTBG
NU28SRjukjRjMrzUWkyvW2Wrvei082fv9f+ivqOrSYDUiqn/zpmvVQV8LZ/7wAfv
VH7S7iUKpPgHoRCCr1pFmr3+EmIckPkebJI12s6YqB95m/se7uh0+BSb6eS+dxt9
I1AaUOStTf1dbKszo2Kz4PQxdqC9cEzoaIw48bk0eyPd1wXbdDb6cuUqMns9+ZM+
F/PsLYs9+giC8+DiqMR25dypBi1CJQd+L+bQcWoMonHtjyguP4hk/HogXMiVOR5u
9CMWpc89t7P5ij7hGRe+2YeUIQJU9nxktSLQwfLCjM0fHZf6aeXtUnKG/Q9IeRUU
fYAUWr9eac7NNd+480ltwTtKzRPTsP8YXxuyaY6Pw+piM+u+Vrw92IuxiabKsA6k
BJZuLCtA39ihoaEnwkpNpudxRNBeI91+xytFOIqK7GmD+r2nMZaIPHkeyElXL6Xf
7KEIqQnZxBMpTXsFv+gwKyTUDEsc75wagVi2LrPrG8lgQ2ZXNzJ9yTNivpngNXxM
qVraoydY2acGdL7VooE+6ROqF1+mIB2Ro4fsVimfCLuOhAMxdY0r8tUa6lhgPFYk
IApZq9iJax53xa9PhX1X8YJ/7yeZ5r63OLN7bjEi0GXakGOVpLJvDaUrFMdKtjuf
Z562/Lica/OSkiFSCjojvKZUS6yz+x/8r82WfreK/jXCyQbqScXRlkJxVoOSdto7
SxswGYhfHSwVoAi5fFf9gIXq2HWNBpsR40HelozE/PHZPkzkbXpVgElTE2s4edM8
p7E+/Ej816ruYmVlEXv1K72nKvSKTlaAGfmfD+0ogahV5i5mquz4TxdG8gYAdB19
KMJr/NSmu7Q2HD76HhHO8n82pLVQtjb66MegnFEpR7db8KXapgKhR8me9IQjtxqR
K5Chn0t1c4Blmil2kgRiz0LjEtUKb8VKPOOTxN8mhAJ90iPwjyULklX6GJHdEeti
QtNKGu7nOOIp6M0n51zLe1MbjwNgzGEvSfzFC/KAwET8O9SuYXBZZZ2Y/P8Yqyc6
RyckPNPbgM4qc6Pqrwa5B1eBauXdA3px8MraFwCqBJLrU0ki6zgvPY+dUe3Mtk0m
j5PB2q6zBId0AWA0qiBoI1xOWX0kwkTbc68pz9kzdYnPeITN4Q6V+/Um45mqtfXJ
Ta2+lQxj/UEFzOal6K2nMASEZZ9pUbiEhUqGh/QJXGp+tUg7tByY4/yygAvNFn/1
wRBOywRB79PSYOGjxL6HXIhWEOwRjyCglVkdxXRvsmIhM3rq/8jAuVkkfw7TSBHt
+eFlqWIor6i6qn15SCjr9jtFJGYKijUsrSvLqMiG3EJo3A9HSz7N7JT4mLN/BJZc
EZSww/FLrU1Z+nexGBKmzPWQ5PcCskvMtRXyzvs/1hWZ/riODRgga3nbgFglDlxd
1DRyKg52k4+X5Gg54PZr7e+F7TKcouD2JL0rVyuJ78sg7fL1/IzNNsuTs4SwL8Mt
Onmc4qTf+K0W24JW5pokwDMSJIK1waqbR5CBqLGshYChPA3Tq+2a9lClTsvyKG56
WLlJOu6jiY9yG5QkeOSOH8zGfstZMBD23BxkzU1/mMBYcg3UQkQVfk9ehCbwZSLw
8rlGOckovHZLIhT5JaoGXQwhtgcK7xZvryYOvl2+eNdc77qsQs+6yci6eHkFJrzm
h7DflFMMuXmBx1W3Km6INOl6qsbvg4D6qhyOIOOBn5h2s1bBfiMLJCJK0Usvllm0
MtAZ/7IE5nD86bLQM+f7piO/LbylxUg9+mVj6H0M1goBQL8/pVkaRoz1oY4e0xxh
XYAPXG8t1yZt8/YPdagmO8T+k7imxgHKc6en25B1OrLlA0IyDob1vv2soPZTv7Oj
+ugObu8VbPLJEQEF3AuYQXd44R6AfBOjgJBdzpDQYpNWDFagzm3uil8x2BSRK1th
Gb7PnMb+uNC4eNKfjWZ4/sx6iBisScDdP07no9cDuP8L/dS76B87w0608BPmNcgz
+Fr+YFv/nDNVG6RAeS3r9tRhlP4ptAdtaBU6l0CwkWBcUIAFIr5SvyCGxlG7PcGN
Sh6n8vPxN44Ige8SYsGgEKOulhkQlzdwQhWf2jlHy8ywHAoK0SWlTnUrma6BQdsr
VeTzqcRWFCiA5zVNMQLid7tkLg5kZBNbz2LnBuyZikI77vCiF3i7+HI3FOf0UlXU
Axe3Je49r5HD5BBDXdvsQw2MIOMJagoMU5yfwpmbWUeEdVNNE9fSFY7zNEE9ba7z
ATJO3lpM1jy5osGbDxf8CfaFlMWfSxdwlGtb6TJskh0emvog0pGzTW5ol9BwUvpu
Y7XyzzDsjcj33AkEJqiS5+bXBsGo4rRMacGUiZx0LMz61DbCOL75uqWmJXAWWV2i
UWm1zLVSHyV0D38RrXRSBk9PK7KI/ZWA8KFWaNn2hnpmQHFhSQFjQAAFY97WLmi6
E1+u7LsYl0ABiC1ySJVPKIiIVPsssIuNuxW7YZNPX2tuIxfcgD9kSgd68jmrTD95
737X1XM8J7G1HZ3goi/klQTosS9wafK37YhAKg1dao9SyyQoF/cs+BvxZO/caqtu
fjCashmTXu1WZbCTN0JX/pgoUQykFeIHxq3kztmqDc+zixTGheIY3LAuI5MGCEzN
rFD6tZqB3b78PcJsS3kK/ObNX90WjllA/xutaPuKse4M0jbq+x2v2luya882/ZL2
VGd5/7h0sS6+bndhFtWGIJtOmXd6KVhZAc3SKz4XX4pApsxOdpzW/ay6AD3XWpTz
rwRBxcOv9Bj1sWKitoP4FPDHajhtEaG7ddBmPOBJpf6RhgYHwNQoBHkXpN44qu1h
I+KVOTnBt5TiwOx7cr7LzRoEXia84cViyJUlucj3DWWQrJMzfMOGueJPsu/4Bovf
rH5/ZceNPTHZqSEFsiCFyBP8qehheGwvRVQMmwrQRDnEqqh6IFk9tVzmxLTIILci
6Yjm0hoTXpnDr0NngFsQTDUCNEa2/OW96tProDP7tyfXX5MofxqsHwiXgpKkePSV
wOPdad/Uo3zTshga3t+cekUF0ufVhbAUmPM+9WGu3JnBosNeYpeq7o1BIQN1MLHW
XEWNrp1bK/pH0rdQJ6rKSHKXAP9WFZKMjxjpERV15VSd5H6BIpXTruSK6e+RHEOx
gsaRbYdVudB37lho2/B5nDaJyKbfYcl4jPjS9vGrU1/HGCIA/XWxykAlPCNqsaxq
x1Hb7cQ8cabXFe7Tm6BCX/cckv8Vr7SxXCqy4x4Z2lGSnlK0Hdc7QSCtAaAONzg9
ofsn8MijURgTccoycMaUkuqjNa6K+GgwKJjlKo4F83jiOnW7dQrCzPBQErvca2Ln
S0K3NNKoVV7lQNgdRRvUaxPidXSJZKBPB9EGlai6CD5DFSBxPIqbHkJLRfrEuRP4
VbQXHidA5Te2ybqad9L3gUr2Q31/HxGo/M+Avunil0bUsMtbnwkr0HLnBl+/pG7z
E3FSaIwD+xq2INYAjBtHtB9BCrVIxMxUhSEtOfI9eTbPLsHJC2BQva8lG0eKklvn
25nl6z8HqfWyuFtzLDwkoQ7ojzb/NFLjPQib0QvJtYG5Z+hyWwBwR51/HmiJqp7d
LAQEKx6whPkM/Twp3mNngxtDiWmj4gMAocaBU2TQebPT271TAICYR2i7I+GEmQfg
4SB1Y/fL5yByLzGBQf6V7qliP+0eYoMYyEKUHbOZGH8V+x8wKFSxEiB9Vj7uzV90
Cqqn0fTc3RxJmZsfl0Cp8TPKQkLz47zB45hLHIjtSQdOzkoffsV9XtuuV8PNQb0k
pUiY7Xa1vl5bspfwqXrTca2MGV/gvOtQYTXTb6q43EaZ3D0KpobCBe7cjDm+XOyq
TnTpgGN87azvAfXpfcCfSTWlBWM/hpmIxdMQG8gJjQ7E2t9rEkA8bjdVZjHh1YGV
1J/HuVXLfgqgmijBaVJvoU1WfIEp01jTyXZtHPN/yCF3Qy9GfUIz1rdtLY2r3YNb
2zn1p8HCjnSVKcSYasnxpeEDXJ3KIixRXnptHR4HR90my17dD3+oY9OUZYf72Bjn
lPoFovAdH/a2bJxZ8daEkt+O60MHJpN/Ky8gTbnJuM4lWOARAPNtiiBYsqUNp6DL
+lQjD66Q9RmwXBUy6zwMHIT4yCUFzQE3N0Mtpc3OXuAcM7bZTXBlx9qFr5UhwbsO
BiVu9bqnXO9LnQpk6SYOw4kD+LWRxgXzAoYRzs2wZpz5gbDmDPqbe/pP52xCDs+N
IzvFElsp0C7xMZaXlCYQoG2keixnUkktYW9b+1nTmmdGV5C2VhMH9jKCQsB0Bz26
5NIGqhRZKdMiOC3YsYyBtvd4qgdGsx57XAd73/8vu7nIWiB48wXogsSYC6/35/aL
JwLcHgk5yfVuwAfkgrP/aB5BrdbIRZGTMFRP4Wr8OYZhuO7RapFW1YFKWzE3FhHE
Fg3DRxoSHKdSLsEtSDtUHKMoDwnr9/qdZidn8FjZrPtHnnJ0MAnGURo/G9w/AWV7
rv56DhketPZro7TMz9iYvAXKbaJqWTtT3vY6NZgN8fZY/615wU1RI46n9lcvEgGM
5Jhl2RSS5n47/UgxvBi7glylQbXUYJ/JuZGpnxHw/s5s0aGUDl+dUdnEjxyxykIY
zrFRwTBry2gG8LeaM4Xm54CuO3vCIW5wNyDh1AjJIS9KbO8ZkLPhc3zqz067lYl9
Atpftcv2j/gh9TWOm3e4ozavtyLTeNw8BUMdtQQvyuTOfhy+pUGc3rplB/skIPhQ
Iw4gmAPAT7Zhkvz52QGOE1k5j0ljfOmZDBaY9RVUW56wh/Khl7LsFWYeoc+4UZoB
7aIuWEyEs+E4lWN9sbuQ7cMZTFWnwZzQVDEyJMM/js3/BJ5o1+ZMfZTLqGaPovgj
0H64cbR3paiDsAg7DFb6K0LnqJxAVdbguYjC3TmbvVFUdX4+v3SNSb2Ium5rDMdF
DFwut+WyZWnCG+FLVErFLxFhhnhQKqggABKKMetpMSrq9FcsM99pV8Y8Tdr6jL2J
2+6ejzZYT8Q3xiAtppaD3SUhDSo2RcIlF4NddmJ/tKpufWSWuU7csMS6CDvfvRpH
kwQmHRNJXpajnWYqc9sCj0U4D4FATInP6HkfhalYz321zBkrS+4gEjAmo7zirQiG
GxPZgRu+aWC/8RykXePOUtPXD66nLog3ElB6NhmqB/hNpgS8DeNhPza/yWHoziOT
FnlxObSwJagBnlI6KI6n/LV5IZr5DQnlOv20APrnP+dWRaBYRDoNq8iBcihaJsRM
nDJIrLIfU9X6sJ0ALv2jV++ANfbO6iXcOWmxkj9BkPD2VF6wnWbi/3kjRGtM93j+
otWnx0Z/MdS7sK61shs5V5JHcID25GJ9d8/GGaoxF6gAFciiLNi/XqlSWlpW8IS/
KcYaCtTzdBzeugqb9q6NkttZv6MBYoai3ENaTfGiYvBnW+XlkYf1GZx6xjxjqmNW
d9iYGqbRc2aTsCUjhKrctLLFW46VKz6G8c4gbuVHNGnx+GfjespPra00Flhp+pH9
DznRC102dpYiGgZsE32BcsX8YEaLDvQimOITxNURauDdjinsaSLLaj3LD3eZXorH
JFq85oxECSBtyrdV+cTuwspZMWuFp5sn/cNmQCHLN7i4vAHIktFIHYtE2IK6WBjz
XVVqa7g9SeQEXHRzswBRX3Qyvlr43ruRmuZaAJzq68V89zvaWQrktwOLOkudz86G
H4KWsrOLQGr4UNQJa/L+Gvt1/r8ZEaBVTEtsZzx9KeILIB1/oUg27yCneVjRhyEZ
xU6mBbHHJAFWia4zERomtsywz0PdlhjicaEgm7RQk/RApbCzPXcYlIiQtSZFY1e3
Mr5lXW3Ji+zA5TjoNNblMbDRMiHDFaRUk91zyB7XuFR8pMMwq9tR0x0IO0B4WqMM
caBanekE+AL8F28hNjrp2YIbwCAuPXOjgZ0MFYU4FG5fVcLGjH/t+DmO1wX9015r
2JV+eBJQs1+tlpVqeaRHWPpQGhLkWrTzeEVQYZSYOwaRujh7m2IhH1iSLpUDIN1/
GNHIO26Y5gxFXlhYoKiyZ5fPY25qYEp7+fs2BhY1nlIJiy+fylVyx3OjHIdRJ3R3
LUiyklIR5s9Zu9L3WzaIRbDGrV3/s6a105lxuKWlJxawfDf8epcGqNs2D6EnRiaK
kJb9QvjfLdURTeCUqV8t1DIduS1us7XQ53tEY9ec8JKggnj5X+XwRjYSi40VT628
6TuYMfSvHV9kRqZCuvDvcoA/pkAG6xIJdaUxftOFrlMQgDurQnv1XhKSRBeL6W08
8QETKucF2QqnDNMo7D/J6vDiFeQzAap+xgsFCmMgrIY2J7ggptGakQ4A6i4mfb5q
J7KP6Xo5kwrB9bX6f+9ZrocVGX94wmGz8cd+W8nvvp7iuBu202ISN78WmpBYQFWr
OXZQqaDfKmjEPcv8yCLiBHwl683HHp5OJ0Npbtk2KqWRVBRETK84ZGb3DOKJNYBz
61lnNqylEJD/mYIyAo2nbrfp+E4hQSylRrkFfEHguZ6oamgDKDVeulZ8Km3E0VEu
CUR+d0eKXUmbheXW6YZme241YfRycGH+uztneKthZPEFYZFduFASROMCl+gIzDBM
47dO1zdZR7p3BCY6z2qiGx571HumNpJtlBBt2UZudDgRfLfCHQwvN3o38hUlYLXQ
9sjB7ZVHV+EpdDKqfBf+mXE2j1E3WBx3f02YssXGEjnphBzL4ZLUhEtz/shTBUmn
zQfld8Tkogt1VZql0efN7mwAXrWFzTlQeZjKm9ZOu8uFfn72d/YSCsrD2bGmz9+e
FC/gSHmOKlUASn1d/KPn054on0YPMBZFTkC9KHSnkef46N9Uk2V8dhX9WOUqqFYr
NlmCzOhVnOnxZ5SNt2JmJGlQDqtrUQ9jTOO0+DoTD80rL9WtQ1nXAP30TZMQjA+j
KJEvOjZMU6U4oILt2ZTVlRKoZeZhlLWchBKO6UXA5Bskka8fFoPev+SOrYN1pSZg
ixjJ2yRe5cBbZAxQQeyaCFM1ZFZsvthM3PXjWqyTSFWRaCp+/O71UkedN9LtFb/7
/Yk65BA44VbPKeHBbVkb8fJbIyvlAcYMxApHKGQ7nksjBn3YAO0HoADcjKSNI6qn
KpfpviRKjKDfu1v6HBBqGtj+QK3Qp9E1GWkHCDzQx/rMri1uKfF6zwWb7Uet8RNq
a84Dd4+Mka15MBIPBSPeP7QijJEhHPy3htTWbithH8mfP+2+G4IV4wl22itZCXR1
616HkTWW/lQA2tuVPPv8rx9b+Ljjb84SOXo7n42/A/mk8zgoi9RIA69Qp793QORv
hO1MfBFgWQk1U7BEA4ZZcwRa9RC84FUfrf8tz4XNegqi+fhIejTgMH/fpxK2b1Zk
jSn/mmm0nJWj7SEwI2snA2+OypSPztTVIk99hQZ5qyaC5dCzNaafPeqHRoGT1C75
IPOeVtz0rNXEqA5ibVArbMVtuXXtEvzg8ub48lzCrQpxHS0/IK89aE3LxdF6yniz
FKF5Fd1QNYH3K7upe7hKaJtZGjykJ65a2Tr/TQjKwJbzc/H+6eWDq8EV1Fkw5iE6
Ch8Fnd9Tfo6NyOt04rIVbTWXT3yvqqZXot6mTzO9Dzo4fQ3Z+1CAGV8vcerdhG05
jdtHgkIH0SkwjOJgXPk8AIvT2GoXULOjR9LUd0itzkYr/1P1ypR8LwQ/JiXMXsKR
1lXbH5/vhuM8hxH+jeHrs1u3V5jNPpDuxGBHUcJ7VQniTezbOfESd7EMYawPKufb
RJiuhGK3rYpaw38mF7Wbkdw/KIzaPMR9QK/iDNtTnlTbp2gjqYujZ8dIdT1qMK8g
rK9UrMPkSKpgpkkYpG91Nf34aXQbGYjVehhoEvqjz2NuDqRZh80BY/Ap8pCjv2PJ
X57V0nBUDbjA534bwapiy/EobAP5lcQJdRREcVGOSgjIfSFiwcXJJZ/UedX2CLCI
WNu4K81Mu36hHmg/ze9xhFl9jBBO0Bm2QUofojk6wXArp2vcqdhnRaUYdfgvZwTA
CShGjZa4RKju+soCHJrzi2upk52//Kw8yteZ5kZba3YpMaHSSuv2YeykRcwYe2Uu
qtRL8wAvOdSUnZWPW3fY9M7IoU8kQGfvrAtis6hmGcwLye9GfLEyXOHu4b5/Usd4
xRo2He7zj45Anv7GDQYwu75E0QslwtCeWe3NPTt5/I9ZpjB+NL3sn4d5iCnyYTOL
FGRy+zYmYO7GqbuTEYuwNN1eBz980jFmnICyBbZoX07a3zJpRI9GirHiNttXia0u
HWYkVtuZ3fYMRo15dmsLPefFsGfAWUIyyTPtz0RV2cD5NFQwQKe4T0vN1oNvK5d1
E6qL7BczvYn+MMpkSES6R6/Y2LyAQOTeHG6RR6SINhGYYRJHkLBEsFxSJiD6M7kW
ZtR3XD7S96jjpXPN3jjWjN1L56dtuhATChaXwN4tTheNHkRYWS76LSvPQRZAfnph
O/jdqHARL6BhgjHdalE0ZfkQaGuQV+BPZ2Cyy0XiM5YGOLMMDvb78lVyAy6tFdI5
ZAdfXzdEbQ9MLNPgtQlRGrAaLubLdaWHAeZttDLcBnzZ8v5yCh29dYeWEzRmUTtN
k5uGgpqkytkhmccvaJwYFDFJIEhqmSvbm5WnEpriKChtDLKPXHIQKkaz6p8Bkl4A
wL0UgbKFXz7zLrHgpEwEH88vdQF+oLYiXXR6keW0Xxdi1rNzLw2dNL4h3SXD0TLT
qfnjK/pIDaIBHobRXcFEpal1uUEnzMNgRak109v3wbjIsC0rvMX8czya0p64LWf3
unHXGxegHqnwJ6Hho+SUsF0w5TXCyrbVGyC4p2fc5s6cfKEpnDJsKsBoaI6LH7WW
1DJ+KtjBFplVCoRs8Ne1MOSvzZqrH8nYWvWb4dO3/g4PJ+5fsItKoHz90HikGDkd
9E0J1eg8xrfryqrB68KCjM14bPEfCTBcM4prK2+7L8RZhvWaw/8IwZkWj0CrTXzg
cU4lz3FLYdOGEwIzjTI5YSYn8zcNVDKjewec2cu6m6WbkOdQqfAS483XDtbccVtL
biS1m3qEd9qmPyJNFxC2od/6GkrR6A9wigOGVeoETYoBfFsNA2eGxGYLKT9QtHkC
mk9u9v8y0jaffrsCjQFV/dyr7SEpQbp6LtRqYrQwXG9Unws8Goek4tOivzx+Rt1u
lb3QZZlB12l898LJ0RvTNykeKSNu1njX2hMs5gjgddEV6YC/VTn1+XWyPUczM3xB
kxHe5D5eheKypDJgX1SR32h5PtvivqDeU4rdTQ3LmXArMhMZTlnJqAg0MPQAps1U
FOzPk0CYzzqQbi75TCcOHnXBcke6z9rD6i/bv0w8nXsd/SWkA8A/C2tQYzyIkf28
GKJ8kSj45PdTGKIZF/ja8vxb/UZjKhzdiM7d6beC4xeRrB11hLNfpnZha2qrcPy/
Go5F+MXFB8JzS6PpOIKhEifSIrNpemjMuChhd8Z2jxMbgmheo3a79RIGByogG/LS
mml3moeBtuIpz1TnrKL3OzWdCCRhCGjomAxiPZKceNixPCxCM+Zsi0ghji6wuibz
7r0ZAcgjRFiz1pmhP3jTcY2NOnklPI9APArorr4jBp1N6SPHh9BikDx+Yiran9NR
lqgVIBidyvdWCAFSbrtr0XuM/Kpy9b50/Dn+hN7zFAprLJptEa0XgYUgVjQE44Uk
992MPPXQID5w7GbusCdRBRT2R/SUKkPmUjU6vibv9qfI1YX76nPnXDpwYjzJNkOF
hnrCDPhtUaIc+EisSgFvkwJsHg9qDnLrJODVBHCcTDfXfRfpuBeuiq35D4KJpxdo
NQkyOrAe5Fcy3PY06fm58s60fApNqb0BbxGHXvUCwfj06yv/HpPsGLIdanpG00l6
gk1zXD5/OMEqWtAHnxWu+30K4G50nISKiryguE0DpKUAsH2BZoPYMvXuO+Kkzvko
R1KQvnmNfQVCjh/qxkp8H6GppfsnHrcPL+PtMtpsm4tgeTEjM20hv+GI+q/PvNRa
BM3z1b+wF6sRjwEQ2HQbqUMKX+eBs7t2NvLZwCMmYN5+BNYMHyONt0HFlmWC65MX
PQu0UHqbeFD801PayydFfJIYt+qXV01dA3ETgxlH6IkIQL6DOhbL2BAzyB9YWHqp
wDqkjMSrpK363BGg43WgOZs5aStbnTO0a7T8BUb8WCnjQzxvwgzY+5wv9OKz4TxJ
bh2mGXYkkaFWoz7kTwESnIuRqbkA1vZk10AUROGTR7/DppH6ii8iTsSni5jePas0
9uZE7+oWOmJP71v+rTQxxEFjLOWpGOPopiRfaGqhprmZrmILNVN91f3I2Y3K+H65
nd1QXO3NcR/G8PbVxa35vPt3G9b0wL7a8FlqlyuTsjC2rDLf1uFadSqDUbHoFr18
BBmta0X3LkZsT9ggnH+Xm1lIhA7ZTJ0bvalmUdQCz+qUA+9xtzaZRQy7mEREraZB
O6LMbGJCXWCYGANx4JyWfu7JbnOF7w1MdEDXhxk3XQEE5zvxJdvV0R7UVb6PeMaI
eq4KO4ZuCYcjZFMBcAkyl9EGh+80dGdR52Jk/fGx0CWAXLPQNUN8QQdlGWW53v4a
Xjgs4v92g4A0vwtq4roQ3ZyycHPEIleUf3wwiX9aZOqu1Rnm3n5DTP8e7lZTw6Yr
0JpqIXvjKKc1S10nvokDCs9CxwDak14a5/TwmkpSwNGeO9yFIEmD1UiYUkk+0xAw
l5oGau2Sgy+J535f1G5ndMHCuCRSHqHH6LRWdi7cGFm6NyabbqYthUVPsUAtKVqJ
Nhcig60pZ1BwqtNc+QjKrV09iC+YR5O9HoG7eQfVwb5p4bCcHShOpZqq9jBuzzq5
ZUbWg8GwGLmBTRIrCFBqj0uBcGGXmKaY7L6H8ZoD0B85MLOTWqcDOKIrJS/JtJCM
2a17xLbJylmWudZ4ZLQbT7Ql2MGhwAtlGif9+KGVXRB1XomCEqWk2nR1YcIA00Hm
1kWz5Cln1z7AT2iGQun355/lm6PLBtCXvLGPCaXuaIoMHc9lIYLRXFYZAKgPCYvn
8qLi3/2GeM05X8SGHh91Qd85LinrveQpHnEffPfKSruntuX+Yg+KyWH/BSYEJx3A
h+pFJovIbhKu6eAEIaITYEV5O3yZKc1nZgSoT/7SHDsITAOTzGOVX87QJfCrrD4x
3IZ0lxro7xONdf8PR1+GzvWOl2Lwg90Oqme0wIGA/KB0I4Otg2DaQRkopbe9mR7S
7hpMfJ/UgiHO8Qw9p44QVbZqpsr1VGybw22W1d89LLX9vMdayquNpgipJdeSDU6r
6XbcGe1vY5EdAVroIa7nePatADFBKXMrNjRUmaCnK5F/i6UpnoyUIiu3rlmtJNLJ
QPy3VfEumTHkky2eo9dMEsW2dDHPAEYMnku5Nfeki4S6288Hh2UMfUv9DufJA9EN
7xmxsgohK3dhOAvN34Y4Gqv6OKFgi8S+j56aJPZQZbAhPe0jkFkVW6Jexb9Z6yXo
iTRPRdqMxb4gL6DbtHB4/QeA8CI/zvZstIe4mu0r/lJhLiwDMSFmIkoA27V3cETy
ycDNswRgX/JiKkUQ2yAfwbM7KDWiQHHZuv3eZiU3UlXEfOnCZ6L/meTWM+nnBj/B
Vzs0X7ww69FLBGBg6MfSMFUHRK5soTZImyGmVvofg2DBAUBfc81W6KIGiQvP31d3
WJYce7s75JJtqUX69FBhca/4l7ZAt+sYXaINWNgRB7M21n+iebvKGOfMlR1Iwl/G
II71YRdjz7Hdd6k0e+1wN6lH62UjVf8mn7wR2FmFjBR8P90SJ4KF+GrTsgwYYE6t
6FhglzkRvq8ZEhifKLL8X0VN4h6wQoxlu1FmxguqVpuKw7gidhdp1jhDNOTh/C81
/eK667ZtvW3kVUd24EJEWKcL0Jkd58QqJb07akdPIpCZphDHBAu+KTAFT43rvd02
a5Issp8GBLjin+bHIFwiUDOospB3qKgOGM+sExuD+JILd7C5PCyQ56vB+AL5Mnzl
FesNlCV2aErnBd99JtxOtccXTIq2+U6tjTOpKQfcNvIkGyA4r0fiMXSEyKvDpFRx
JZSgsZEEKP67brasDdSQdF8p7PkXvFRh+lf5EoGEzkxVsfWiZyJKk96BwawIcO2Y
8AR5ytqOcqlxcpQX5LWl2eQHLT8hw70IN/WLSWIR+7xbXqzzz8PsnLShCS6YBPN5
2hzOA+D274Sv51lP32o/Bxg+dzhBagS3x2fWnHkw8YVjJ1b6/YgvO4AIaoqRwEkX
fo+aHLpZopRorJibOR6qwUlJF2xtJys9mU4Br0DuCkRboTGCgK9dnmOQaDUPr0nW
j6ed+niL1i/KjnpokWf+VlRn8FWGH3piYcNf5E5wBJSXdrH6x2iFOIcA0JlCWezf
jKbyw3j9BQlaVHRZzX96VS2We59Ip8KIALx4XvPHdWBAUlviBr7ZZuhRMIK9AC/J
ACbL/yOJaCLtIhK7RioRGVSqWnAmdlgk/weFhUW/LM9jJHZz2s+MmxAAKIEEI8GY
EDWszr5JRm044X5jrRdW2ZL2nP+TwixOzSqrLnwMin05QQ2vk79A+JEUuHBx5BpI
7X9oFvNWsRtaQPUDetaXZRkvEuMeWY/y+JVtepOvmUyaiQC7HesmSC8+VwV5u8Fu
FwpV9j7dTwuWOvDiZCWQnonzxTfo/SWsT34lD5OMWLcUvDWYGLOHnVc1/nrrw17C
a2YcNpbSH1iI2tXRoh7epH0HzE9HUpReZp2i6olOrA5c8XU8sbUdV0JtJvoEpPCo
pA5wxSGVHyXUBtjPoTWK9+HtQzXIOcPCN5xM6z7IcDgOSSCwIONRs5O3rPxIzRF6
0JDLOdI+GM+L5p3hqb6C62/AJpVWaRrTU94WJm63z7DzNbDi4b7cikVwlIhC71RB
SWkQFlq3dNQsntKp5gGaer8QgeOXLPFYpe3qgoHutwDTXhm2YCGWWRLHelWO3Kc+
BmYT8gqRb70xzOgPwBvIxiDSbMEKQDNhOyeqI9N0NQ3b0hNZDe3cjKxR3Ww3AyII
FgXqnMx6KsLfJwbXdtheQkNtHdmY1wp13qZlauYvnSi1iOyKhvSu86DHoF2mEKHV
1eB/Ny14x1Ug12p8tY1XPYqBjFmDlhxGIncGSxQJbT4veB4m3r+Tq06rDXUTT4bH
2vXM9YkMkwhIawhfTsxQlh7wW2SlvAZUE1txG/cKHIoOOa4/vzuu2tWMEpbihYJC
vwx3VlfHqLHUJCuNvzSFCA5G11/hAibrpi+LUh1D3BRHOfn/kOIJvHJF6SF87PHq
kjKjZE8Ncf79SfJ1/NhEB/FRkfHBLtuRT+h8ZUWAyvGLfm+W4xIAbNsjIqyljDMp
n8qpGMEpwQCRXow/sThN14kkfPBiaCCjQPm7WbwNxLawCzfEI7UqtR2JpmufnLH/
DSNF9ymW0u+iXkOHI5/Z6A1ip1Qr7XGhnu007J4/v/IHMvGsMjcRyTzY9EUBtoXa
JOu0N3LFdI6Cjwluj2gmoYML2vdAgyU9qikapG/scAHruqI5V77I7DDSrQfXad/Q
YAEw1RoYn+QqTPw1M+gca7sQxtMLq4bMrrJZPajKfcfCPm9zOwUWzWmrs6t+E+N5
Vzo5nzeSXfa1Tr+UOiaElWmDY2G109NePsvv9yqCjsjRtfgtNoeCYMEIDr/jTZxZ
54fuLRAFTG2B6/PUCOk0oHoWwH8nIaQ6i5N0y0TBLs9b6+K3wtjXRkYLz/ZSyoY/
CvvQ+lphFfGE3faPX7HODzSQrQ2Qsr7nC/UN5AOc7cPYArK3WWQi30LZl5c+N0NE
mgGtGRxBbPoPXmHIJIqJCZikCNBTiL/d4xkCp2TH9yv7qDguFyfVkWXBRhUzFptd
vc2kfr2J5w5cLUy8pT5JOyGBZxNVV7EIXh//o6vPFVd4SYLV5Sx1Huv4wX/w8wvL
Q0bY+7trKa7zv5mXWYF2nSYyALU/UVBtu0+fOYfa3UssNtjRgezs+M6qJMN6y7S5
aHZJe7lPuGiFkc8e1j15Lq2NX4rjrkuTVu5m/SdPurTdgc0llGdEIzGL3xYxKyxT
PVxveNsaiiGkjMKTo5Y04qAkOmcANdId0AnxtCXPSmYOMRIq2+Hma/wsWFK9pCak
4RI95GrKW9KWoF1LiQFjqV5V0ohaGMpuGKaaCNroWR3JZ2S2S9r/2KAJE2DCPDav
V76vCbCn/bpmCchPoXW/XMtsy7kucNZOSgUrEKCyeCC8r6liN8yjz4McCPVYmtH+
mYd0N1L+Quvq1tfl8Uj6QL3HpwVy0pXzsWGo8TD0BgJ1oVCfNqLzmmrfQFtwKBKI
aUZFHT+qpO5nx2mQ2PRhUvH3C2/wgMlnwtgxdA2BEEerKyF7m84tyredISAvUzmK
XHyYe/Mmr5lCwHY8+DcMHzZS8SztHkaIFxRuIU8xHQlPWIcJuqXAz+7cuQCAfaYg
4IHw1TJJwklD8MmMsfeBhd4uXjch8vTmnl8XN3XbKi7eaR4r/2MLMiVpdIaCN3wS
TqOte5W50e28yHHnqU1785afvEvTqZxmLiIKqCjJD+O+J2lwmXWs6NtRKdkWMuyA
ARma5qQ1fVAZxX3GPp0qPIlqITA74wkuqdTdfzoZ7M/8ZPN1NVn+0WeFEX7lvIvv
0QOqphMZnnDuZiy4bJxsrP4NPDuePQN9r11ca6b6ulXR1cKIqATEa/N7QAUQoZmd
8Thl/9MS6GeY9jtki3rY8yVsgrt2zpCOYp7sy1Gs3KGkNZKDRiYuACObb0UaHE8T
X+I7tKIq7dCtwO794hi5LgwSQXd5d9s+UUN/nh+PDM7ixbQjB7Xobx3YAzURu3lH
xGWR/AiRO172ztQFmLdMHCpgwhpMYE5L9PmvtBc8eoIt1i1zONXc4VeriQRF3sPC
bRuzyck9BictvYZq10MObRl5PUrRfY5N2nIg4QjjjpU9fg6/oTvFq3K0+6kur+KD
YcSybaftjDYQzx9uOz6JxbX4dH+6XMAG6O+UGVEI1plWlakQMtQRskYko+qONeii
jvJt4mv84lnM/A1Cz3EkCCEr/Mb/myDs+/hgjXK5X3ahu3an6iVXSnHK12BDr3b3
8McwEYfACrb3SjMElEA6Xg12SG67FoEYozLXi5qxRA1OVEvKJL1DRa6tHAb5CZjS
JO8EaFVW+iVBHstXIaigrwgFLD8KHiL/scrGivgiX7d2mnEjOT60EpvPMPJAA5Lr
SF9wJTPYw0DZTXFfjWwv7W+lzOY8ochVciydf8dsAyQsnAgPOqwXH0EKqsRXyvrf
Mc7Y1fC9/ryJMVabubWuIvWkwhxJF4p7PmsVpiWOMkHs1G4AiuJvyRH/m5oiHoxO
Dq3zeCNsLlHlC8J4nI/Y3odnBbflnusttoJ/57cANsima7crS63IhajZq4wBHPGL
bbN2WtiaHa5kvA04Av4UVGM7ezwaz+Xx56v3W09lkZZ7pWq7G9+GpRqI7v+t0Unw
a2rCzPFOkWpUyJ4LwKQQJe9+tqAOvi7B4zwIAZ2hLsT//vvjBdDc9fAqtnbPzgI2
PQ5KVdV6CRvOpWSCnp5//Lp84fG+f65iPsp/eaGgQ63v+VoDL7QF47PlaAbjefEA
Xb9hmRLMgV1+yB/lESDWEdihc0UAeNOnRGxv+qqM3lChep1Z1ELLRtU2Srcwo77y
j8d/0mizn2LJNHuoatb5t+gobEIcjQootGGPoYaJd6BOj3sXE81i54lUQmV3UyU4
kxcTTex2YPFGv7ebJXNOWS8l48i+soCalfvqZkBXkHPOcdBM9ogrMYmYt8IsFVpZ
YaA6k3q04UD5B98pYTYaYfeH7JKcLcuyNn8CulCM68dFvT9kUY7x+UadSBi+00v9
RSlZ0Rwpz347m09pea1YmVhvVoMVcj0NAi1OyqMxeRNt7D0qoFHJrLWpUnO1uPcS
GQVPfPVq+4WESwiOhIgJDQTsNkzDum4vhhJwAx5Vlzw3UanJPAQOvRTzcLjR6p8p
WGM4I3+EZdK3eywE8sUGr1vEvDnanM8cD+Dz9/18gfLoIyU7Pd2W9ZF61xwhqGWC
J57MSGw2Pg1xeYVCLB57734Y0pn0B1e+g/ToO7i9QhNsq/zFcMxPHqUrzgVEfLHO
maF2LRQSeknLk7OLom+jRyIkGsoGOnMItiYcCd9puFBEzTikYKk8m1gUCp3rILRK
h2oh2KZ04ty245dzTpdZ4ZliA9JJg25Dc3qHJCkv0vF9KkvybzRl3XfvEmHP3gwd
YbqNN1T7YRzTUg70RvzjKbvOuFHPmXbd8AZ9hJrl4yqTNNgpux9Z84hAIFS1Z1Nn
z6wGD3tsAv2CCSZ0pPyx6A6SCtZlga6MmmrfkuZipu7s10+K4lhaId7P319yceXN
Nizj1zPlSUAIiNlHaI0Jh+Q29dQzTqIElCKyDQG6BTdogxrUMkMWJ6CUxfDdLmab
tQDI1NZm9gaDqTXCgt7F0wzFK0qofVxaOXHxQx9jqWJ/s3G6Tv0tUBq/Erhkc8vL
hsqR2aWVisj0azfMPMEShJTI20iSchwh/OLlRyU+1M4+pEfZclfWh/VGKw9bzs5Z
2WC1MilLs5vxLvYc3sGpV2hApl5HyOs8MOmH5dGFlHnSCK625fSisaPCVz8nuFCo
6ofke0e2e5LNSnlSaJLcy4OFgFP7uiDdPr+cdwQVT2cs7USPd4LOdrX6Iutlq4Yq
fsMsztSarXFF5xMSlf9JUEqX4WpFLXiN2aZnR3HDH9CkZ3eMNUawo2oMvx50+nzI
NLG7NG7+HBX64ek8FJpSj4+D/pWK+rzCQjaFH5VSo1H3rUjb1+Txctk2QB90bXgs
Pwj11w0FMm4m2WGOCABT3QGeOFOoiWx33WA4rl/zX8JoziZ+plVUBgKB58r458wr
W211dmpDIYVRulAFo2PKYRZGIg3Zx0LEbg2CPCP1tU/hx329Hjqht+kgatSVjc77
/nfXJlDm1KDX5Rxn2nAeOZ1nMaJUzQUq81u7ZuisHH2gfyWA+TQduIjC3S0c4Fa4
2xzTFPQSRZ8A/qcU1J+2gFMuvAbyM0JkPKYkjOUoSawoO5V4a42ueWuuNcdoM1+Z
oF/qvC5ZyZhheT5TfZw4m+mICNLitXxU25EweqBWf3Qg8kwN6OVJO084VyfURN8s
tEMMjQWJNezEtmPuBFYSpRXpt+VHjdICkOsqSdwNa4MNic4NPubv8ZTtagrF07ya
jAz9tHEDu04sFN8fjCYhOPeDOQp53J9XonbOiFqp3WZn8CL88it45DQ/rji9W84s
RHHk3GY4tyLMyNg19wq/Q2NSEKt72PIZcYQrsf9a20/DOpEF8FsLFH7NhMYRcWa6
tkxw4flyv+/J1es4cWuFiTQmSDoMvz3VeWmqWgNph6qPuhj7/kJwatosA8WKGoJj
0gJXf4SFdSTqv3Ij/hPS+U/3/LBI92bXTfWIDB3PeE6+BKZtjLHnOTal/THZPT/Q
rqEkmTIQXLn4Jh9g1+VOphT4hGihZIRa9SZV2QrcV/z3TI7i9XRmHfDR+UXuxFJZ
PzV6NUaKweLa81BU8dj657UBEV8IiaAlJpkusxFnY667Ta/QnsQeLsCieoDPDxff
m/+TkP1a/Ak7n21yUxlH1bFVllXWRjKerkgkMFwgCo/S5GjlwXZZmhQOynp2oc6G
gA9za70jq9CTSnLIwYu+K2fww/aNPNIOa6lX0XRRS02gZ8nkwPrFsASpbuBQE5G5
jVYFyUZYkgHDJzOxU8xoF+I6uOkZmGzjZ6N3gQ4EYxLnoWeFIgvRfwoWxGLmrjv/
ULi0uRlzRAZcXm08Os2SH1rdGwtys3ysr19bwk+UhjuLuDUecISD4vTc97sfNecb
IqZ98tkXUYIDfg1UcQf6/4k9q9Sfjy2a5g5uzazbUPqAHzCqoUHwQbVCwOxg/h9j
NnGh/CfCkhp25+sSbRe/RjZwVR4N1CzQGkzTXMcn+QhX+1eo2iXAQMZwserWXf0p
5lzXhWOpcKUS6usEc0c+IArSVsZhpgCTSElzZJFlq2PcMreeZIYIH9ZzGK/FQDWz
oc6+Xm8qO8tUn2MqDSCmOUZi+sGYNK/3qFgRreDz5J2FalOo9HBkyhVkSt7FRh1/
hiNOfel30yuVACZfK8TiixJ+CZv4rjcpbMmw9MYiZno0JmXwnR3pSXlJJuwWDufJ
zR0bVv9IaPYjnfK3HvdnI8yJ/9DP3zh5Cj6+sJxuuFq3S5RPJKCPheKKWNjDDcZo
WKAOSPX3lBeEA8wSs6U54VtZclNYcOCohnM6PQ9ZavbHZb7aNGzFTKJZwGS/t48C
Zq5KcvYO0l/VJMigduczwS9MM6DJZJN7uVuyMX8i9g//gKf7XNa86tO3HQbCkhBy
nZaYcMl9OqKL6wzzzjPwJIvfbIPl2z3BY6kIBRLZX7v2KeLwRecJ10eMRtl0LGvy
0SqU1RhPhRXCHhIbWiGyITTVwHp1NFGGUViG94DGGwX8Va+VGOvwbUYpiBg2+fiF
PRZ59dYs1jQWzNV3eCnvIhuLW13+1t3+aPBYhf7iYN06NdEoKjlvvpfGSY2lCtzc
y0DtqjmJlwsde1RepyC0YapxyocnFBJYFk2lyxMdUmc5sVhKwjhU+laY2Z14ihBS
Cz/OQgh+bJ/jIWv7bN1rpN3MA8pRdmKVlq6jR5xbKGRJ58kra2hxx+MrBkR1ocFX
8wKYvWD0gKHUHWittPwHDO0hYBCO/fvM/2U0p9XThU2sceTzo+UfDVYOYWEhCokB
ue/uIC8ILqpSNaXRwFyIp55gIDD7w69zNpcYhsnY2cZle59GbrOAuzaqiUgjQHpV
KFWlpEXq7C1t9uFIG4iz1/Rx27XzBbWf2L7TLaVrvUVffwfXUG/WAVZL+g4H6EfT
U6hBAFkh0VjC1YrkNYNMxICeKchpS5kKvW6MBmc3hzQxb+MfiODme/xDczxSgaHR
oWjcLX24MWmLXe6zusFmtjE1aWzu80Dp2d35SeaVmOIi0XBY8Q6hkiW8ANC7HU0S
QxFVU9z88+TTdq9Wa1svwjKAmDvZlFj8jPRv4nM8vKtj7N4Ecna3e+sFWPcprtfO
qv0aFOkTZYSlArajcqNc5+O7qJAPvtiXA5Q2vSd8MGw+LKIb4O2142PgTz03XHXx
kwFbUfdOHKmnis5AcFw/xrsX7UgMdE7N4iErndl3cfE7gKyCAqWSm9fGNSC4LWVF
J4kNb8xuMdA05nyzihcyZW4gij8/Yt8IV8+6tW+b+Hi/pVfDcdpeoT5NG2ZTOc6d
byt3TwpZZjvF12PE8G39Pmn+sA5p7Dc+GNgKEAxvdDX8JRfZr6eks3T1ZcZRxdP0
yDWJaRy6Pog1BBE50zFH01bOUhvjcs3hI02WO5qUq4X4ceojInSzr7nKzUv8HzQG
RBsntgSj5FFbKh8lppPIGRLVTEOL/GiVieMUW1+Cd8jun5/AHsouOEw6/CGT7slC
VzLxDHmwWdGcjsZB3IdRc/jn9gFI2g2BR2YOXAPYRV7anap2ak6eTIK1i/U98HIT
w+OqAU08EDZscrPioBjByPAf/lcfyUrydkRjTkvY4e8PWvupqadLKQN4Zzz7pOHz
2Rz0sc0ZeGpsmo6SvQBptpo0OUUqueBm11r36IidAL6fPEXGwK7j2kNGzezaBWsN
xaLo3CSERSMlLZtXT2omatwjoN7DDT7occbUsmY5jD6o4aQ1FTzmYnQTEnqPg6ZN
WSQJIHw1pI6Mrunvl1HHz92rcKCLSIEDkvITW2QkLbF8eLLklvJcsQvovOIUM0GT
QhB5+Q6IDoWLBWIo/sjd42q1/fSoJ4mFdkM6UDm7HSNKpkX0/3mXyweClQPLXzRi
brXjh6XGST4uri3ZOd6pSKm5R5F+IkTPnFbIcIeWKCgraw0BoxZzOv+0lnpFH6xV
tsN2Cxpmfx8RJbLh5zRt9PqTcXqh74s+dAK3s317C+5TuG4tXcwzGak62GN3NB1v
KPVK3txwqcfutgP3cBm0JVKQIQ73vhL1XHR3RYWCrW/1I4XclVr1aRn8T5hmRm1/
i+GSfsSA2wW51wFUXzd6gfapkqrxsbNSBDwfXqv+MsuYOoeHkAFRQOEINIj+wuMB
0DCoe5MSjgmEv8/IighrUL/ArohM1SA4ByZauybzcVgNXNXG13PN76M800L296ex
TThPTSHgDSRxYb8FliisIfOG93EYG+M7qRJDvxw1WUxji/SAg4rb6YKNXY8pUBXX
xKCD81Rahm3WIP/gUgDooaZ53YOeuZgTArivgO29JbhZ5WDIKlPPV87Bl/2l3CNS
ltc/ZW+Wv8tZhgNGn/6AaR0b9dBsZIjRMJ+ykMaK+N6L/Jh0ui0Ux2cE9rRnvVNI
CL+cpIga/EuVU7DGcbgM06IQZk+PqBWkXRrDeUATmDquLR5mYDk0vk2PpNinZR3b
xCf/+wsZApOK6F+F7ROT/CZKeu2nBrnLDJdalvMSZ0rgLljKTCiThxnhF4jDhQmN
lW9sUB9wPMe8q31vfzdI+kj2L0SrxgaJzl1LcQFjqCCuAAstjwm+x1COfM5LcIyr
jzchuxoP21Bo1UsrFL3IwC6v3ZvFqVSy1ScFftEUilZbeJOJe5EoAPKENaydruhb
cVmV8VWdEJlSdt7MtCjrV52h4rNaGySC2y2GQ8nBlZolsUOUt9i/s/DZwLWba/XF
pLm5V/IbwfUqGpnFEdnvCbZS17q0NCXO1kzrlbHkWEu8L5Annnc92UEEnPHs8fFU
dxW+1Abd01TnxHOH5Hxs7TAS704/o14+YSZKETmUt6bglrHxRep8wWrH9cOYPvK5
Nxf2/26O2BOQIcdPdfGjjIoBs1LMryDQ3IpQgk3OYv4MJ4Cdtdp6E+tza+VRKqJt
bseaLgEz0G0qLfDhrWGtTs2XN9MPsqsRfbO6nEe7PDtt1glfMZ6gp29pMwPe7QRu
Lu3TqW8mDReqWwWX+/IiPaEJl0yu2Emp6bAS5vFa7ObJ4DEdi6BQ8PTRilsWYTSP
FaPdj7MTEwKnKpbUI6F2F+Ibb/LcYgRcX1T5pqDwRiZyIsVPEQ69OQhIl+PotIY/
tXr09qc0i66G2a1zQB6aMYpL86zyp9IRs3Xro2sTlGNnY/8UNrvSnmWrdtEpi6dn
nNhlPuMQXcLsGvmvDTvsPIHP+Yla2IEDkfoA07hG2m9+0LVK34FbuOG1RoxQ/S7Q
QHLtIOj6dNHHLPLlNlXnUEYLK6utIZ/Fbx9TVqhWH0t/4byBR+gGNFyld/03ENCQ
9IfrslNodiVsyuPJKrzTXeiI5nBbY+ezPby/PGfxzxQ1ZujcpQlV/V2saCQUT6YG
Q6CctezaDjjfIJS2DLWfV1EoTsdOC/zh+GQWtvVmtCmA0P1RSXFhmZ72klcvQnBv
iSkfUV9juSPyCvltMP5N7o8SHunlZ4w9dqnTnIr0J3RdxHSWr61J6YGoepskEhGX
buO8Cd2A3cVfQ0NDtE2OtZ+kZmnaDNXidPqS7vB7iARX6ocW6cJlHerM6/sMKtxJ
NQ44nvZ9FaspSey1xhfiCk4SzH+Hd+4tKLWfkD4Y7bKOdJoiYVz9erEDqPdxmuzL
6Dc3u7aMEG1gPgmjUFFLx0lh9Xa+Qo8rWG9Ea/cMzN7EdWDFfyeO1wm5Y8uxqLC3
Da4MEtE4Dk/4kTNEEf+CcagwWcAsW3MADb3hCOZcEYDc66svGrs4NW4BHp1ShZIT
8A/Az0FTWuN7sZb6JAm1HgX7nAXdNCNL8dBFTjSygig+zidtnk+aUAMXSoH9Ei34
9710xMKbgtVv/2dxHkB9uGYOC1TiWWGUfuBQcFmGKJSLkDRbYUpAu1k63+Lag6FM
8OiJKziOeUoooc7S/Z5RQjeRqZY76q9OHFyEHnDJnGhgKPp5inBCu+QOmLEQfJH4
cRozO+U1RKw3AUtdi6OOxCJ55ceaTYa6U9TBBhuqr/1MNtEYqaJm+QKf15PQqe9I
2WnkCbtu5hs3md1fPz4DT7+iewUCOPXTq1jpAVaR4XW2SX1VwJTkELGzaiKi0xPa
PgWqK0NiqBm+BmeEqZ+bb9cCCFk5OXEm3hYLVYgRTFmNf1Erq7/5snjDS1ygb3ST
WAKSXZkz0Xi3WzKBFQXusTrE3h9oitYIsMbgtvgZOmcOV/sYdufW/yU66eG6b7rS
IGG+I3GbNVelZb5/BaPf9KW5Wytece6Z2kUHWXHt/ru3wxyXMuvHnfnSFmvrLHeL
Y1DostgvXAyhyIDobhsl3SsHDVMXfmxpP04mrT2mP2u8W6xRzIOIz7zGbhUB/LWA
mqAJ+IR/atVRs6Q9iSfM1KlYhs61+kJLkwyNv9ymcT2WKeh5eUmqZofB2MSBAVxY
v2vk8w4T0W56iMSgAcc7WgRk1coHSeP01bbDDIRpbmA7chb4Rx+B6eKHUf/usDRN
UfPOtDdvPZKEwCjPt1kReuWAfH2DlmRo9fvtU6YGn/oLXB+POH4vgfjwvzLnNXx1
29amE4iGc+7oG580jcqQfkD8FuDyG8FVy1JLC5MPfNYv8/pnJDb7hmcVEW1GMRgi
j6OM78UhjSL34wecvMVxXaBjUn+Z4Ila5xKz163e9mUg6ltocj39/fvpTpYccGuB
Vx/rxGjeUjTNkPe09hNA1L7U742s6uQfhit34sHoWiDBnUjnPJbbkgeFSmpFqsn9
IjcOKji/lz7Sp73I8OJ75zBMhGIFkAeiyjMZHyEjnvdk1c5IKZoPhNC1M0kA2263
PyJReH0YO1CagR4fEX8gmjREPOdTyctzg3Ll+sxUA2AXwJQ616a5URqYo5P1Kko1
7VnJDHtBpj3SC7K6lXquZmsQpiTP0EMh8xD+MshNCc8GUmOhIARJOwxQwCooZvBc
bvvNqKqc7BNike6kBOZ0MhtlbahsysBR1xIiCojbGHcYHp7ZoGAIxjEooEuFeRUi
4dGYxEypgn0CPtT3Sd/et84IHbCIuFDVRgLp2kwp0hL09xQ8Z2XuSYrcaobpwlfk
MNkxwCabjq1q95PdOWD/j7pddjYQ/91HKigMyrFb8BChiG8ovfqUZl49J7J43v5l
LVRrN5+AllwW6pLzHTnkNsHTyy+gJrsmLyLDOrFCUfgOw4PqVfVoxsxvVwZggGEh
JVtr7bIcjuhg7YMrOTIp5hrRLwmY9cnn138ZfEV2iCxZCzypQB1ndvvpkugoEbAU
5pANoVm4OPlAMZHLzq0LfiT34dgPnTIkp3UkdCtr2TBPQ1QbnhpiBThgiA4bmN7f
c1l0nF1zTNICTR7Esabs6vXrLdm1J2FQ8osEnc7wy5KX7ogawiVWPZ5RUkf6NG+y
z51T/V1+fLlFn9710f1YukFGn+h8/qHWlkv55cuTv6bzx+Q87naV1EtNhr+Nj4wf
Sh7q/hgmwAMo1G5rbvVxRWHzAk7EeIsCqEtp9AnT3jIwZLWa0Y0++UHl98VnHBor
je36wh1F/gjZ1yeLGYAtNKsZ7yshP9yEpvMiU/iaYVH0JPkiPVGjQmI0lbVlllyh
ZYWs8zY8WNyRJKfjLN8KjQdyuOVMenhQZci3gNFDd1xOci9iAokTU5j+YOR5TU+V
gk990mI3chXDdm2fN26YXpS6d8faLmjdT1PvsYXmuEGu+ZocWn7by5dcsT8t1/wx
Svqk8xj96D+4OusmUQxxmr9a8IcdfAuaa36hKVEhT/bfQjeei1Kuz0rHGlBK8/9k
3PT2uRaVSFVG0i1qNGkXluvw8CeM4kfC3RJ1xZEvnli1hzxe01GPkbDeQ5TisEKz
0hSwa/U60C7y87l/R0FumoKhNaP1VA+YepbZZS6hzO09UuaDiD6DmQqXbyaQm53i
vvnkP1Ip4RXRq2/Ahw3ztnEZN9JzRlPZJC73iFWuMq7Lhz7OP3y7T/HtzPclEGA/
aELrOMQg79/HsCosMngH7CqDE5kzBDE6TnKKAB5ecrjquwOTGo+z9LHGLJeE/fTT
O4vS5iFoxnZx4rJm85BwCt0CbJnVK96baTCI7aBQSEE5vfBnYWTkdCIhjIDrxv8r
WeX0IiZD2T7e3O30H3wbzUnrvBuo6JuW8/SbHEte+nyZyOin2tQ09e46IgFogd6A
VlB5MM6Hd4axIUPwFyagFhUMsuceQeimGbsQT73WC1b/QDtSBaoL0IuYVzyi6qWq
HCV+1gxGYVWTa/Frek9jshYhNmZNb+JXcV93o/klq2nRN9apbL6qff5d3HQsrl63
UJ1jt3VMYTVYD79WQe38o+obaHKuqibXU6R5ibv4KsRQWbgNcHKPba5mklTc50dr
OwJB7R5LkuDYIlxEimq82X6DgzIKFO5pZe8Zn7TbEQ0BlXi2Vmm/yeQ0NjsUFbXt
LDO17k+IDgaxh2J+em3DJr9f+MqrS4eo05bfX9lESwYjTqA0bv03sZxRQh1GsH0p
s30B3SdzyIVlC/koYbcHqTQ9o3tBFGZCIQLKgbx812EjBtmxq5Zfx0e/p6M9wryQ
lfaKgv8nLj3LesAu1IEtX6At7QqXd/rKLOTH/dNduvPM/PIeHE579tBR6UAflYnC
yzJCS9rbuGgkuksGZ5XzZRS+I6NjLiY026W1XAyQSRoMDHpEN8hw7aoP1gc93t+5
PGZMlKpxNaZcH/9qeqQTDJYKC/hazxtTTjfdsuoWApoc5Ajtixy+36EVU/VtkzXw
KgzZutqXtoZZDsD05OK2R6uJV8iMJD1Wb94AgEVr109PcKc/wJhKSYNtTEZg/1Wl
dBp9vsdkFfDlJwI0dMUkEaChfsHSihWNpaWhHnqyDAhOeFaLqBc55GELWVOJetx3
pMFFHhEOr4AF2tL5BhUsigj9URqwoyN4M/XcUWNFl7VR0jRHBk2hhXeFYTnCXe1e
kELCwrrM/eDDOCtOWEUdX1Goh8FoDi98l5sorWHF9ONegsikaXk/2dUPSXUOXQQ6
XAidwX8Hi6FqZkhk9DxQQqxFOm7+M5Y+DDep5mtcHSwaMh0Wo7TmTdoihjn9SB/0
TbCNbsBtuCMKbZDdW7Y3uS8Pc2nozjtBQAV2+TTOWp+gfiJEGrCSY+7lqbWoh9x6
UebHBHHEv6Dahj2akQkm79bNJS26VzYwgZGZt1+LhZCqEtQdF9hF2SMOGQU7gyS2
wrqNpXsPpLzDOhaMhPloj7dhZAOncGi7tiVqK4mlX/y/e1UcCK/+98gQyJ3waNqI
xRYozlj5c6luah9nOynmgPxIUr1YNMDgKhHceBYyScZXmJtwPQp6kRyVTdlZf6tQ
nTVOtBX4IaNju73rOAto5qYd//Mv3ei0owmN8f0Dw32d1n4eANdDI7kuaijHHosl
+o0qNt0LR6yL0Q8pCmvU7TH/vU4TgiHxa4qyJVtoj7YFwTBOr22jJNJl9bUietyE
yIYGfT1iO47bZ6jVU79odPUp9/fLM9AYxpgywkKW7RSpLnsgDvNqpCUJ6fo5E/yb
Of/HbhV3SrA725PIZ4JpbXS2UQ4cbFPUaTs0mwuuc4Jf77VScxUvwmLOS5QZ9reC
0YO1cO4I6aM/jHYVXEadd2o+CJ3GjVRzYpvyfre+Xikf0dC0e+Jgd0z5Dm0+mUYM
P8yzD2PJNuzKD5hvXyqiG8GLrSl1LpMzLrs2GFBuJg2ybgtexixRNrcRaPxnrTz8
b5nJpy/TC3poD8s47IOgDfMuU8tzt0UbpMjodC+UqAb627gaaOfbgOufM7XpWDLU
FayfA7OwW2+1vvwvBWTMd9opdXEfzouBLNRiQEB+YzzYppZylgwkqtP94OY0Y26m
Iz1a+jRI4YZV9N3xU0xgnJ+rWFcBRd7s0UXrfnd6EFd3U0cF1SYDtowT6ydE+eab
m60kFiI4eWfOr7rmyooWm1bNPqsGA2ZZwcf0VYVMARDe8Sur+lfApKM43rjTfsdT
ttUyQ1PUQ36tTN44/IC2Y08xpVKeYY+fVnv72upQ6QQrx03Idbmpofc2m8GWBrfz
tXbHoKR49DcuxZoj0DYDfZWyCMM8uuQX6AzVngbKCo+Ul8e+TZD9et6yuoK3MuCT
WxPAvsr33tinnXcmHQ1EAFjQ8FjDLJvP0Crc/C5tiZkq8K3mux/Ih6q8eh44dqzw
is/jDhQWsZjYzaNIQt40++NEh/SPom1g91AhszzxCXjY9XE6yDMQT9aN3xufRJM3
gtRh0NCdCUKYVA3mF+zOttX6agPHzpgkH4E7ztZB4R+2F0vsrOkisGc2NyFSoG+d
bjYv5zKoRUorSXP0YkhKzqisRxkkXXqmjR/up0Kg+6u9RRFtWalt62k2O5UZT9BO
jVjHgC+AStz5uXquPKI4RD/DgZFobICHh6H8U2FsFl8AX4ZQ0OQ9oyTelo2q+Q37
98DFVIgdpwsmDTWL7baoq4efl9CTWHZnAhIB8pHNHQG8GMgkqbY2L1mFjHpDHJa2
sG/173UN4/K1hPwHsft03//numWcncnwdk3khO/OGh4giINeHrDcP7vLHmBmc6Av
/n+zseOL7hlmE8/4JVhpGs3ubR9xafGV1R20HHA4D5YsHe9FpCRGGQbzGOUB2hTN
P6gklJePHK4LwkFnl63ox37bihXhhQnLEXcz7JpYzy9HwIZyWCBWOIWsaPQcijj0
UrdaFsi4su2UOHjZjlMDCYqRU68a0ssH9+XQNCT9H3IAEyIYplWgEDkrpWTGssbs
gQVT9SwNbabgtkt60oLKdbRHNPu+XC2pZdKUmkhG9+3FNoAI2PNflEQiJyujqlMg
nTDfZ5AYemT3Ulxxl7JkyAscIQ5YArRyjohaZdUSj4UxMik5dTCNktPzpfElJCyJ
fvvxlekPKHFfaprj7NiDCXgvyKinUf/k2L+Ro1k8DVQuOxmwrsf7MB+t0exuT5s9
Z8Ul4ji67Iq62WAcXTiglet1gvIFAh48p6bQJ/WgcJXH/DiLhSkOjJzVXieKTh4T
XIMmeEseW8lhvq4Z6QxFPqI1gxzOQyHCHo1pkx5PXMTO1gKCcFC9Vc9EDb+lNFAl
SKwXsgClFXCYyEBuypMm6weRx2eIJGLAD7Z6FsGO0lnPcVFox9wtFWCXPCxflQE+
1DfvCCWPCGwjV05gI2h7utXjMOEHkzEpKZ507UohUpIFhD5hEmDmQyhcqi+lK8dF
JwQymF0cgrxbLseuaDt2U8cP6yoUk7/BRU7fxNbV/KUIXcHHWx+0Z4P51hYTPJip
Rqa3+A4orgsqGJAF/rakhM23XBYl/ariacDA8mAkst5XAZWF2Wnlv7p2WHhw35kg
AzRpuDYLv+AAFqi68eK6G9V0/Tj9eqtP/jIh5OKDpfnmndpiHvumf+1PLl6nV5jb
aCXOirSSp366HDtiqDJ1sRpdUc9NB0JXP43PGWnNWH0x4d9NLaUCY1Y0m9YVkGlw
1qYbo3LTMPBvBNKXySgeVuaxNdF7nQq6qpoJndtiHjEA2Dmb6kQtif7WsUo9Yc1j
g3DieZ9hpNTi1qzEfNxOp9bJmrGu9P9RxuJ5rTVe0amJd6M4kVjgjO8sOXefo1p8
nN+an/QzkHdL21FYFyG/aP/nilq5Bj9hU4Z3Lz9RqJq7b4flTab2kljuwgE/z9wQ
EL5ndJAzpFS4lEdU7VJG8e79GwVtjlVOX7Uo4QnbTuhdQC7sgpWHS5+h9xIXXqyk
eyTuwKfYJEJmPR0meYxhFlTuSjzX7uylnveDThBm61hvyiOxYbkm0huMwYSc2uD7
xbA4MuZl3LdIakJ+Z9RTtohPXzs/aG88/L3y1Pz9kx3aTfGo4AeL0Lmmyg8BUy0o
fnqdhqrdjuFGZMYUblSzOHmljEXkYickM0QZMQyqeyHf8gTxLEK/2toxQJ2bVPLl
npRbWbwI/Bk/pRTn7kKtMsFzvp9Pt28utHEwiBTJKx97vbmtqPI/D30i7I1Dw1cf
l+HDNtRZ8HZ0gcn9yzu/Q254aXoq9p7i/PodlDbTFKAb9KjmSVZPg8tW77z8+8Gp
YgNnqdb9rDGaRVXA83wIDnEmGVS78nHTFuPHUL8hr5rhCCklJWeqDbl4+NQlCjWX
H3LnNdNTR97jUIRcc+TYJFuLbLtDyme+Z9wBUJSJYRoH/7fGKLbUVqcgy3xFvMOU
sE5rbuNcM/t4HdzKK0NTEMPQ2NLGeu09C9yIn0txMNlTRQxPuzIaknTYhsAyjLOx
nu9Ej7PiBG+OZqRoxtkZksP2doXDcK5/HO9O8ywNmvM6uP6ZBt8cSVFxSqnpVRQZ
+4jqaUjT/nxMaaYf4K6Nulo8nYDysOLJhOet6DUWHWeYzvZ5tI58nyWRnlDHVVlO
uu+EJgpSTmCDfF1Flpglrs06XIr5ILe6rN5qwjCslNZIW2MlW4yECeif18a7V7fL
GUc8oW1fTSfSKyRn3AyBNjUupaWorZ0qy1sMim1vHUjZ65CaCYUy+saw0AhVra5t
Nti3QII/PhWy52/yy5ZX4VU2DmxVySkXzUYn+b6uxEFSAklp7l6u4IXYlbT2Ha7C
81NBHFi15Bx9xxbVEluL5aDj5SA/tvtbLuBg+OeWbDYHjZRVXkNGxpU5fE+blogk
rsmhxPyFik2dHcoES9/4dbPurwlEk+ElcRdozMnBmsncH3HSUYlh/ytsvtYuuv9O
VDkAKkc7PtA2OyJXT3X4B40AU9D6/vOPX6nXnxhnPeuDpGd64h113LOTpKhzh9uA
ws160s2+uvHAipSx2DofwkYR72znXFFPBWVfvVaGUh8FNT5fy/NiJSIpmMdTCdlA
/VhIkaAfGrO8ikER7pSNfxUWjZVZSGhGzyBEsDqTCytqonNJ+5NyLMCJHBe7t5vK
/NTWiTkRG/9hvLGUoG07bm2waOzn+X2ceh6b7awnJLPtNQMTvr9CvrJSHGwSY6eG
9JchrgGrKxChxLMvSpJcf/4z7c+xkMfnbM7li5CC+MXYdSpxF7GU2+S0YoMdXCqi
Nd5pfc/ufh00E0EVjVjZ+H60281A3k+gbuUk17QXiqngsEhm87Uyfmnvug6ER/nX
qgnDt1uvTDNgJiwf7nul+FzpG1IcbyGCeOy9jPXv7UXBTwOrdPCBDaK30GfIzdFy
3geGTSh2xIlGfhVdi4/HFGSf92rr0Q0S0DQLEWdMf66fYADWO1BkptFB3WEAFgFm
hYM2wJu7+yFmDc9u3NsRxhZDD7mnzT2iVe7nmDRRSw4mx4Pql8r48MmzVoGefvxF
OBPn1T0vv8fXg+/3DL31pPl+Xwkta03v49Azd3zgQAmpdu76wltsUUQyp2m5cqAR
hEcDkWk98Lnp8dVYr+qvLWoPk2CBJ9zvZhmuU7kA9+HgcSmAZ8pNvwBjKAnVUWIL
WevpFP2c3b6pegEBKvfHHoBYDiU/IKA7+yQjZ1epgOt2ThzeYx7225S4d7Apzb/I
yNObrG5BXKdHVdfTyAsohM2m5cpHQltdi0MPReMlDs8lGumb6kuvN+YeamH/C/g7
1HCKd61pqSUg0TCjECqLVnA6mAwmouhGvN/45D4uoBtJyf7Vl7WmOQA5tHh7L0xK
IYNWlEXWDvDnEnqR48eroRnVrqskubMHu3Hm6xGw0ktOTwaD/e+3emBNVvAIdYiY
+AqzCTyi8HO18ek1fp8SRJ+CKcgYrZi8ac/Fp5SqQhyZghlLsVIZ33Eu1FBrBhlV
0+JWna+KXgOOd7vEBtQdTXd8v8uLI9zxUE/upYW1TBG+kIMfWd0+fVmSJ171EJRr
+5PtfSNF1XjKZaliJ+o2p/m6FJDfVtOQSXL1vFA1MQcrH2L9XdY01TyM1fiTohxD
vhCrLd9ybYvPaw+zbHD1VB2t/BfYun0K5iWvuUVvQe0+td/KkKF/G5YD6tNwcqnQ
farznd1eHYdEkvydC8gNPyjljpsM1IZZ+yd54hN3KDJIaufiMpnzI+ATXH2gLtyr
TAOInQylZNFuFxUapJV6ZQLdXOLLF68KwyD8j30aEGwavaM8O6mOYoxMT5yNAkQY
pAZApCPP+MYvwuEdPd+Hwo7q1NuweeK7gW0ciB1VVGJiy0+14CDijea4st4f6LQH
kkl0UuKV/wQ2jk1fF/SYXcbGeLPnL1h9lFSy54dUU8TgG6EJB4JX3TX1bAoYjSEw
RP6ezOltgD8A/UtNhz8UJOyzBUC5AM/j61JO33D3vnMru+qttd5NgRPYfMOCoUtn
ZolT9Y9OIPMIdPa5B4e5YRO7JFMzq27BYXPeVZ8xlhEsiyiK3yTuuJ2F7s+LDhv1
wuZ4jnizCcJjWIlbVM9uLbn8u2vEz3KkkbfS9LgO8AD+cNPoRRI4LQy/7lggfcrp
0pfZHeGfCKfPPIntPOynoBA3J5a1L7kLJU8sPF1D2ewJgDBBq0chI8wJe9gIsgO7
nMlqrDmuhtv5Wfq/MitgELYgE9b7P9pk/U3lDtfKnTJhsn4Or+5PedkDBQiAf6Wc
H2A7eZbJ5ytTrYk56maBwRmEzPH3mKl11oW3M3onge0jb/L1FRSYrL/RqRR3g/kn
oz9pQV+1+Dl/LgOg2eKfeDQkVAQQOmvPPfJZXx7W1bvaT36HxCfK0nNqSn8+Tsnk
xcOW/xEIYthtLORGOg16b7WMF4SCfz69S5JR/Iy+XxbKIBPxq1po3QWT6coHbEdh
P6TxnTyeld6KpzfCSQinIsloVlvDFuxlYhTqrAcckI63TWRFNVvkswufU7p2y0Xf
q0AFBBv5gn2jzeavZcHSbBiOgk8D2i07jiNC6ejCnVgmQk0hnOSqT8rNvhG1E7YC
TYqqNTO8JTtfeuwuokmo+NCMuSqdLQ9fGAf3AgDDVrH0A3/f5mv363opAuTa2ZEa
wOI3kxfQx8O5qg039T7kbsI/BUFSiXAZbpsQSwrDxj4hnUYpuouMbt1HjIcMG6Ct
EJUiZcAsJayRKMQlEvLGhvUw7Xr5s0Ne1YoibLHm4ma9m1FvbOcT9uFTs6pVXdlR
ClvEVGwq+7jXpwAzMh0Apap9jganrmjPLmaCGoxBNYZUheVAY+1EGOP2lqHffOFi
v7j3wDGFnfSW0U0nPUVpB6yC7dZdU8/JSq7w2ClniAjBbKKjdHeCBtNe6y1x2bjl
RGu5tAUXd8V8QATK5mfdmzQuty1wRdi3f120K2/juNrK/XpcQAQf0GcN7LzE0KMH
u+9ncTtUfTr7eaxOEssx6Tm1N0VAvn4BpRPJlqF7N9+k43W2l8S95+wrw7/Drjma
hG4erynTljJEn4wDalpNtRjoUFQJCRm/LsLeB2t6Zf43Eje7zamccWUsnVyQpGdU
TiqTb6wR6dagzAiV/3BiyLAfwBMiKBzls0/bmSUOMZkaP6LoI0GzBE5+RWmSv/Ek
J6SCeoTKen1cU+JhJajkVnUhSakBtg7LJE1G4F2kZruW36Yz03dtZEQwrG0nauGF
wShCL7i2YVGxRd0gveYAVgvKo0hD6AF/HDYeaOHhJKsBjiGZVlIToo68RpzFUlPK
J7Q1A7LiFu0yRx4MrdP+qxkfuY9Hf4tS0oauUmRt2wyF9tyWdqVkQlbcXHwOgyx3
3jWjVOS1fECzhqO/cxhZ+GYGz2vmhzkq2Xwua+7+W0jumP5+NmXtZtcsCJBBTkvn
EWwQtDyDgdO5kw7t3HLoErvmAEyCSptetuwzFSeTsDOQ4Ev2E+fD8cIDZmie9sjC
nhl6oCBHnGzFxAEi3YU4KWBIXAjeasWiPisYHDtFS5mhUaEVsI9JrWMH1hiGoxpB
GL8ZemH97sEEGMSfzhdDHEvMcwZ8x/Jm/AEmA6EstCETIOPomoGFVAFqr4NOOpkA
CmL2yDvmK+BpveenZTDm8HYR0FMwTILshUtB6LuUUpuwUlKsWwAZ0CREkf2VKsAp
172mN2x/tezcXzUHt40w7X/Qiqof0twGXXaoHAwNgXuUZ3orLWRtrnf9wVdOKpA7
rzyjiYUAgisWpFRbWEkQFwgfmnwON07cQ+e9PQoqYa2Qf8+1oTQ2KzfYC4SDqG2k
jRxcFpDlkmDHPUMlV3tYK0ci4ib0WQa/1Crg0+WRnq8v4AZiA1VqXWP/hGkB4/Sk
zipDZwTchqD5R7xD9WHCeVntLu3KaKjV6EOFS/C7ABb0gPeMWljr7orzC53a6NHE
65zd8DNUf2lSrX81mNB3kXsVwf3Ag1v7/19/t4k3yLpaoHN5jAHdQBQZ6IRH6UNO
6TKW2mArIF38f3UNGdAO6Ul0EdNVxqfY9Q0gAvIGrZihk2nfONEDWwH2jkq0cP1m
aG9PIT2N0bKWRUQnYGmeal6tI8O1V4bcY8YjhJkoCiex9OMwrouOF5hbyq27d9lJ
R1UZvGbdlnzlBpzjTUqs3YewPDiM+RzrBfEOtcDk6oFRpp4Uoi2fEUnNMj++xthD
ij5+4ufHTFiEVjycDiPcVPHOrjjuFnuaXVMYy4lYVMP2cJ1J3C65Oj4O5ogj5HEu
04nKYAmi/XwaKIUztk1MtMiQUkrAy556Rig/IgiyC7wmF2+pEghkNH9rh4VpQnqM
nw9ZZ0oTutgocnnp4XF+pXv5MbeJL3zr36VM32xBm3Yi8rvB4pE2xZXkRHRuOWYo
OYKvZhrMjCteNF2V/Rq3wzOjZi9nb6q9Buv7GeSHLx3noAwAV4LGkumQTrGEQ0rl
qmgPz7oAOCPdiqWW0QctIZiJ2G+GbLp2ED1n6vj+m4lE1GEJZ2gnHQvb8z/ozvQi
I+HhN3IK3N+cYV2VzLx2zhl/L1tX9A73yYP2EwSBRmJ0AaLF+mtQPyyyZwKSZj15
G51kmr/cDmsUfts02wrVZI/EqPTtW7slz0VUPnhny/h+7fc4+hD6muDzYYCkGKNF
2JkaeROZ+hwNXanZX5eN0ykBjHu4/5GAE/TNWfXShvd273Vj/ae+LuUNMj5fPCh6
EC3/gtl7kzzP5kfkDLCQDz/HD0uMxY2knxDUARGDe4WcghN14WRJl+KA0bV7wGKt
RpxN+E9B7aj4UZ0/rgk+Of5BZUvH01JjwG4iRXLvkItwGNDzJ4AXpT0bXfdWy2Lb
eLtSgUFfNKCUAxWmebmVCxwAX3HfuS5cCamU/5f+jeDwnTeyAiN3B6seLfUhByiQ
sgdiQrHQJ5eFl4tGE2OOM22xiF3obH5BCLuamo7vmRJodFi8mg5BPqvcbUAaa61/
1qaIJqNau+7pckLdJhbJtt65+HEpiIDOK6Kz97O3FAhxIgS7AmdQQID8iPfNydoc
rC3Pyr1juGdmiWIq1PhnhVQUDgARZRsPQ3+gKSL2HKDNOTOru0EUqLslBgt3YP8o
TD8sybKVP+o9ItiLx/hfqe0cbVN+hOZ2s+XW0lOB5vZxMGK6e/gvdE3tN0RmBlE4
DLxiy7HO3pBxrnOXM4UiqzcgXTtWO4b/zDfqxJr/nB+7dekjJcClqiLnpMP2BZj+
/3B1TYiHTKG2nhYjMlBoiq9TtjIC4y35I3XKp0xGkQkg6DLUr34EXY67MsPufToG
VUUad+H6gWybN+xa8W9gNUkK5BynS/P35oh60wN+Bic7RG+9xnAfowUJoi8u11hw
dgRIK/CE60dFQQeieWvZORLbii+5W6GnG3drkwGtsjAjvfDcpLGklcX1qa2bofdh
pQoaFtnVu3ffYh79zryQQMPMTUg0ch1ycVdguDSUPixWNZqgfj6IvzQnUwntXWU1
nX7e9btjeME28807iGYy5pfX7O52SfvAy1mCXteYQQq6lCoqPBbaKmIVoSLABDFb
sXNwt0dLtbS6u6Pm+kwy/sTOqrG+M+iZ4ZYIWsyXUTpHyRkfXtGKxvBDB1aCgY+Q
4ubPuJk55H60V0BjiKXWEpd4Wc6kK1G+DSOWXACumQECD8TZMv7qfjqXI5ckrkkr
hvioODNkzO8nUJ5nXOCpCzRDRJrVx7gupS2UgpkkB/CONzbU/d8+/f2sQ2wpId3g
N/zsM+cL+gah1BVq1O/p5FcpBeZs1sSEAi+1FkPl2UERPUIbRkIX9I3BppfXzPGV
BJU5DY5h+yHY4DX0SC3+2cFjPvd/tqkfG8V5ks3Jhz/4H1f8bhjmb+hOayMv/C+8
1HzUWUJndcqGiadR3EoxhbYC/0SvqIIyuse9GgVDUUWPnO3LpdGrYhMGhqC2XHKc
SZCaSq2266cDmmhZUB04TmOLE+yDAA8gU5zInLcEXU7yzrJaX1N8+7Xac2zekRyf
/0ARZHfoJdeMglhLeGkeNpS+sJeakYBYJfb7sWD3g/mylZzU6J8RtmkULMKkGOTT
vxC4kKmyx/PK099cxCcoFRLaiV/1NG4MHUBaQUAzkwnebo7EfKpnamU7fvdD2UIB
JMR/vfLqStc2bf+3MVIgt19c9cFNU6dku3x/0wqfz9fGRca/kb6HMNIfh5vOpgUf
6CVtQaFAQEwLnFMFurmTTX4zMKD7uR59xxaloZIvIATd2Edr7qCSOHWgmwOqqiZS
l/hMJx2aXTPKnfuQUkDLCvkk3d54nO24WFzxnvNpJZ8TBV7vehuV7YsifrOeq4kY
rKFHIB8tCU4F3V65UCrA/S6FNnetTH8sbBGEz1JsW9bJsQw0Vhw9Fq3oJ3tMzEno
iImjK1toZ3K9XX/r296lBFzxM4BRiknh2LZ6vZZcbymVM2SwvW5Qg0SL4GXDQl4U
5/xmdpmnKCB0DgSJG8g+y8zp0lfFIEeYYV3VV5nyDJYDcYHHfM2PcmDVzv2K5RmC
Gs1drr8sXF3Yf8Pr/afc8f2pi2/rr40dcdWSvr2JLcVgwcFZ7nB0TXvdEuffb9rB
Xpe9dqVMn4de3W1TsvMAWiW2C0GUWL2C54vdr5sbxlOTDICEEuEXS9eyASQicBFv
vI8+liW8MV53mkmnbjB3nht/fIP7cEfs6zGsH541pXQe5hakGAu5IEVV0g0GimQH
xX9ZHbd/fAVMmZgxs+IvJkkdoZQlMvC1hS7kHbV1pYFx/rcUg2RNaJqwoT+2Iu/w
pb/NYYuhoAjji1sAxydKZ+RshCEExIAn8rz4n0+LZvlC29IBdph3AI+F/9ucrqS1
CtgFW26f/cF99qvx55AaO2mLkva5701nMt+3T+PfOncT47etZCeGne6jVYNBB4ZU
9y6U/Kugpeb7ZwCH/Hr/QD9tq6SKNOKtRRNA8PHxvQ9FqRTiX3sfUIUaCgJ0ZzJ7
lZGmh4jxfrQ4Oa+vQH6y+IlTy3HRZKyG5qQYqKOY4Jc4a9VarXexg/Bsp90tXmRj
yGSGgi1g3y1aUzkoikqvDH/8IkpjQhXlfDS+P19mjzZk9U2dmkx+1zrWncjGrB3w
FP3/CqvCAM4qCXq2oV9j8XcpoC/ur3Tq9Zbyu9jagN1I4dIu8xxPSbqieehfBPbD
7rEmtdHyouURgdhPleglR/6gGpZcZ/Lhw/Z/FKM2CyluCfntmje+glGhDTHTPy2r
kSSB1mI/Cka/zQFywRHxa50tVTz/nifnkWm/jUmKWgG6jysA3DcrMiJ4GtEbfXq5
uGw66PHasOY7ZIip8TICd9arLZwV8UO5Nm9P+JnqsnHFmm0JvGh6kKBx+Rhf6SFs
fVwmWr7nhbAOKNU+uNq+BbLJJGVA8zI1sPP+WNK7tlHWehx+cFMNm+iO0/mvp3c9
WnmfwFYbkssaNxaOoIRMdAUhulSvIaptvOkmh66ndYJJS1HMy62HpakdLIL5wNQk
x4I7D3IO3+449hFAtUdA5LcHVHY+NOZ0JG1opcQ63aCv3IhOYR19GuEnvqxEcFJy
oEHJtGQYeafIMJv3Acp+AtcCXZYfpQmg9rgCxmbOnJwyQCwC1ue8l/dSdmfvnpnV
b1IXP4vNYUwEvU4VPcvOluxdSbpr0FzyMuG2mE1XvyC9d363jOGpCVbxbtzRdOns
hlB3Udg/KU8Ls0SXcQZTJl/4Sk2CqFiYkNaV3fBBBhd3UX+YJz9XdR+ZAfk3zrfR
d4+vqXyBo808NU+XjDEQgZRIehAONhUDdIlS8tX99KYauYDFVzZzA3NQsuyMg2hS
G7VWlBSGAeO9VjWorvxgzlIHoWqNquW3YAkUUnaM5sYrB3k5c7njK9LDOkX4qrfC
MJFXm53Gz2Rk+5eAnwKXksig994Nm4rFWMyMIru+JqTWRX3yitbr4A0NSVHLuhsS
4vASJmAZEdxBZ4TLJSlKi/6dFZXQ+tJg8qLz51/l6ydofAn4T8BBhY8/PRuvoTVx
bqMWwfd33Tur/YnCmWpw23qw7Hern+7mGxToV7QmNtHJnxBPfaEMOVT04hnhYbhb
3Oi/MrW/hbDguGbyQBCNSBR8Li59pT7yaOisJAjQMkgkxgW1IR5nH3BAX4eu8Y11
cZTM+mgNAopVy9YhahPp+q2SwUGU52sw8ZKjFxznUO2qU6jlxrmmtNLKCwXZCbgS
Cp7m8WcfnDW2Kgw8sNyyxdbdBkDdG71+WBLh1JG+IK1EjBVQFArFVQQfu6qmnKfr
/58RKNX2P/s73np3SXktgp39jcZXw1E2iiulAxxPnNyj1xOhYEU7xP6AL89y1GKo
oX/e4eZ6kBRyojb5wMbBf8xxOu1YCoP52e3PrLJbSOPoXMPv5tcMHVf/AbrahrZn
rtF8+TJgcZ1mW18rp9H4WCk6YxaWL40NpoFnYhagmDC8CZAke/MOpl/1T2SUuwB2
VEn91ee5Der86VLtin8nvfhrJCd6RHFEsis+iECNUsVeWRkH8vxIHXWMY/kCdjyj
G2w4LNMYPPps3ROkZQIhKqFhwZPQeLFxF70jiW40bQTk1rywaS3sdznqn/e+s8yv
RaYenGiBLtyt8LAtSroFptjajkTxv7ZYjcP4N3G/Dkqw6ctYvrVi295I2zmA1BY6
+g8u2QVZKOmv69/cEl0OSxz7SCM1c7HamzWfz0C0E/yrzuYYey4epu2Pk9HzeGvv
65GgozHey2tTbW2NhZ4gm6mnqap/kpctn3pTc3nBkNl0TThIyo/9ciX448rEbsGa
2ajXMGLC+/pC+xWkFAaFrueFkIT7z5XdUBsFl9DWK9L23kXodVNKxAMoHsBmVids
zgqPGxKU3Oi+7EpfNl+k/S+GSWRAeRgKrHOhy4jF/qaxpj4zKd6Wtd0MBFRPpSvo
LQQmlSOzvVuwnfTM6wFJW+51+E7DtUcSkFkRy5V/YXv0hQ4oUsc8rjKhy2O8GPVP
GNd5/zAoJgBGHeIosZNOFcLddfr7c5ejYGUE5isIF/glZGDHI/F3yFNJEmGHxCqK
5PFSia4+buBFzoxgqW0D1MWmA/J098FVHxs934PHYQGoPyP6yTsy88acPZo6tNsH
2kn+3oJ8/Dhh+hcxjtHy5y2SqfLxILJO1m3lAH3Zrjqt3KVXnaaArfRm4PDRb8tz
FquhfkfyljFV7Z8+BP3fjKn0/3xpGUQj83FFY1Gdt8N+ECrdBmq5O1pJJr18Mypn
0asNjOa08gIfVQgLxNI7/iz6IM49O9dDyCt7pnHslxmj7zStB7qyud3TpQeYbGxO
9wwr7yfOE4pSCX0nA/mMaqV0cZds2wPWT2jbN9S3aDRWwprsAPXapKTCvLnA8lL7
k6EPnaXeUZcaal27kRksbRgSue0CJZzgwg57Gkk/nQMHhj3z3LLyMGiesfaikUIZ
naJ+TaD+sfPHHp4r6QDxUNAOuXL8rGSFnPJTZ3uN1SYIdaP8abDB++FB9rI11f5m
CTLVZ+6IEngdoaezwJsKf8ooG4diVkud5lq9xsP+0wuo/DfVN+UYoKVeKxAbzteK
UxscG+G1gHjgQccr4ethftGegGplEo34q3roFE7/OeVyl5tXl3eYc6BtZsUbZqUQ
0HYy5stpEjIlZNNxfFpvEtKGsvyphbvuyDqZRahF9C37mO6in8OJjRAstaLKYyKY
7kTbuq3maEkZYK8tUKoROuQaQHg1QWjG1/RtTQeWb/yWobz6TZBSLeSyot7ls7zb
h+bFBUBIGoscBFcK0sKQNPKT1fRH4ZaVv/qsCw2CKdTdsAZsTr2iWkVZVbeCTQPC
aBf6Lbtm9QukUHl9dw8VVCZkAj9aoY0fU5KfQ2b+smhI0X5LztCdoiaTE2W6UUcm
V8ddh8c5CZfPvGsDJamP4gr4f5qHtsIVyStjweb+W4oFErpUOcWz+K6QCKKhr1Mr
odLlrOy9hGex+SAYqqYcpAUIeyIXnlihO0mIaFhWjN1Y3sCRwvDIbtmzxe/LU53/
uwRns0G6hlDNY4oWz6gnOK1oyRf8ERYvAOJLp0+e33aovLIR4MSvoOgtqqUH7li7
GvBtM442xgOF4Eku3Sot0L8jOsB0c96n2tgURtkf414JzxDorJ+BXTTP39f74sS7
BZuoeYuoBU+1WOIL0JpqkWTddbsNuxe4JDeIB0/Kg9aT4C+r784Kb3qKuGDIxaZ3
n1YduSJCcHHWBKHgt9fLFj1XZ9MpG1P26aetdoOj8nrR/KyHah9sLlVMH3xTsUx0
kiduVTPAzfZkQbZEH5R9tvJtfvPFM7JIdKvLqX9XRGkqOcokNJxb0IU69CLHIbaQ
7sp1E0atd66qjyqO8C54WX8vJyZgrPKGFrHfpcePSPIu5dHol+XFjBPhvUZjlyo4
hIMUMVFRVmdpRcBQysXnwygdtLE/k0h0itpkPYIzr6wOtpmkXohu2XjHym8huJnd
hR2TYwhrSkCAOtjzlcguWP8zL9P9wMNHte1ZvdxgdG/5ByilP4NgdW8ZphOfLtSl
HBqGIoA3PSrIwvQTt41MYoLVjmJ7B4Mc7JW+NQ0XOzlcfyKJgH7M1ZGLFHojmQCg
itGXCP0Oq+sbZpkHuHozQWWdkR1mFLTb5ufpqfAylKLOHDvgLu+rTzDxPFi7mbrn
0nkGUBOMRn+QAPhNBm3nzsm/Pv4cLC1JGE1Gcz6RnRwYBc0cyP7uSqAqgXJQ21c0
dhbqsXn/TgF1Kx1RR4GhAZ+rMF2rFFyS1TJeLt+9AMmBam+FlCRgFvbtnL8sgXmV
+zoniJf88wogiH4rVt6tRPS5uEX2b7ySvpQRHV57B6Bs67N3b+HOJVsDP6UBhixw
yNTL17lQ2eFRlihBju+2a+2eOmae222k4BZWfU2p3fKn14c9yGyeUubMvCUqXOz8
IAbQnJmlQQUe1eWTHfZSPFafl+2D6e1wPhwEowS/guWyQfDiizL6qJPYFKHpEPKM
PRrEvUTT9sUIeYle9TvQDymv6pFhKQkZzayy638emEg99E68Bfceq1aqX8jHjwj1
keZVRLaRSjNJqtEwX1Zca0rqgV2Huip+s2ZSD49+r1CXm3GWPMKMKJhmUTdDALdd
ckGjotFflHOPnCs5UInOG5i2Rm0GMTi7PZwcDuH6zyVLxoqZ9cxnI+2hbCs8LKFf
sSA2nEZpQ9J5xA1xRTyIsBNle7K5wzP4XFTrvO7h90QDeQA3z5nyTZcpsbaLZ0KA
Wp87AURPizlo1jMocwzTq3kWmtoFRf4A9atWR8Xfths3pbFfoGf0WgHiblHmBC3A
zLVB0vnD6n2nY58w5DmsTszKyZdJNdScM9pkIsgigC61bFoh6Tw2SrdHED5Em7DP
LgmQcM0F5nIa2PG1XBWa5IUzq1JuhM8Z6XGJnJxAWl+bDUEZHsvVfviDg+FGY4hs
MPyOOnC++SVPCPAhbTyl9v20QH7/e68HHxUFOOsBSSy9x5i+RyY8iZ6Cj0FpGUAu
zkG7pKqMmfdSI4MqoNEYMZ2ZSD9hNoSSnOrcg26uiA1lzmwIsPL1bbSOP/CvTMlm
EQtBNqCSzL8g2VvYeb/IxrweBjlR3c+CxItn1fRkMrd82VbWze50fW2Du23JVOJ1
N1QRBndDFGbRmE7Q0odzzOIdq4UniLxJDaYL9klaiofitpScBKJh3Tdt/RXQEXFc
sbLIQjdym9purnCn0+La75VHb/Tomoo4Pwv4Zi1Bdg1HlxGZx1R7KobHeVAorJt8
sBym+BN6B0ypXqCnw4xtv1TYGNcLJZDq9MrUtac8QdSnHy9qfT4nU6/6Kjx33DE3
HPwCwy/8pCC+nWNiQ1n+0/6fhLj2CngRBBOl3NzFLFZ3wSQPT18erpYeFG30cWEn
sF4mFpvKZLCwqJIJtZkBDIUDILgaO9DQs5527AflCIwWWhsgLOBCa7hZV9aB3lld
j2hUrYy6BFfWK2oOHnQZctRWuEUQqp+b53deFoRarJPyI+6AsUXcSifccSkhQHxr
yZr8r7j18HABXT0mNDkTBczetjEEbGPqJNOGtG16HED4SzyHfFIZJW4jzeDKG+3U
jbfK15q4cj14iUkC8deqhbMmAjYUuhtD7pFpwF52YLn1Cvk3cLhldTYdC2LPNlfm
C1ixz3UuPfpt8S3cG3nTwO1HOn+sJxuCGClqrpmb8hHFRmHlf7wEJfLCyEQmJ7F3
6SzceFLy9W2BlkJ3ZKeZSECX8a51YSogJG672WXNfZ/qWuWT8XXdrBlIf/oOkAxt
a3KR9sXhAXEE+brXpBpkhExOOy/MDtr6J1j48rCKNuOh5avsRbGXpxvf8g1YaicK
tSOuayKn5FIc4xaZKcQzFYkMQL8ejmP1uJlbrGCdHBNUicM99z4pNyez1Xkyrh+I
hVx7CaDSV8r1AQ8yi3Z8e2xRJICjOXnGd5GeIrk/8yHdN3BGOm3GxN0kjZCgSkb8
pK3/ibYnmHhZkCbudoJdIWIuO6Bf47pEC8eBDegZ4eEhncZWpfBgCqJ935ZaFw6Y
7nrT4hchYLx3Cbwav6mFGkULdstDMvFu1C65YKGrwrcKSbNdON3+D8sw7osPcBdC
ebs8vUkb9Ux84deBRNhfaejeZ2OP6RdcDJkZcLppHDUaR+bOrbSN5jNJwrkNUsPC
LwyY/wEu06X7pualwCnx7wE+xSyeQb6gMpcED7DEfH/3zlLN3Yz8FOOpgyCZ+Gm3
bCc26cxh37ea2bcbSIR9036n0yGOu5y0yGfp0yj7bb6GD+R/XfKoGZgyiKEOACmu
nQgbEmEOmRwiHzbRrDmmbZWfOnvQygDfLaTT78+IyfBSX37/CG2PEXTMCzIch6PH
XFUDwVdDcdMp8j/Ps7F7gQ+yrvgGpgPemeyB/Lxm3X32/95NTXrKfcCBvudMHYoz
rIrbHEkO/2MGT+qttw6Hhrok9FnaL3/5Vf/3qnyGA4DInv4TA5UZXtR39ILaVdi4
Vysm1M69MeBeeEJh1U8+DNP67u+Y1fL88/vTTvpXg4mYEsLFgeraNrZ7dhfaZpQV
bH5GQhR6cbXrz0Zf1TBRTnAcWqds3bMp+aQrHdsqoCxb8ofVubJATlg/46/1VkuO
4XzpXdIfas4mDy29gAywPlxVOEPtoMJOCkkyXI8NvthlzjMdrLayp1Dnq3ifKlNm
lJ3+7dJ846SdE5AX364FtvbGXF1G7MVoDrWkBLJP/5DXWwKVWC4kdD/Jg596PhAs
ws8hJB8iHxTXhlnRu8BXZnwIgUySjl3T2n9rkyIv8YIWO9QrkgX3MVRXuIIghYy+
VyoNQJ6q2R6hJ4Y1YtwYQ6OayUK7NBhB/Vr4GYzrMigYtgWg3HvmTnN/2FeQLscl
CPAxv61NZeVMt9N5m6sxyokFax1CE4fF6bRh3U+pygZPlyTA4PiJ8zckhHu5x98y
ZPakshHYgq5sHEMLVgXwc3aq5dnTbpg5Q5+eefu+bQkEZLiWM1Y3a7283Oepa4X9
R/ItTbJFRat0JoAvQgHrbv8u4QcDKTwME+tRgnhtrp5y15xt4FwRBCFpKQaTeh/3
LN5J1sgfFOzzVb7JiZDMsMMk4REU+sTMWz0Rmirk1LIQ9wqDo1qt2a3mXmsITL3m
AaUWA0MkcI1kV92/2o7JonCFecomUJQC2VQ5fncMZ2JP7VSnocYarOL4PRw4LN5R
utkKzzIFFcPoVXZTVnGKrWhWyk5VONmA+3w6BgzjUwTvfSPZfiyTyMJp5ryF+ePi
wIQeYAsuPpqf3Otzyc5E5bPoE9rX/e8MeIRQvfUu219VoV3mj2PLtpZoWGrorsPY
/csGypUgaKnx5isPqaphNubZK+LiV8kFbNEXm0XyKN7vgxsqNdvlI0+fdsrok2QO
8ArVUXy5oFT5BSj/wCLAjYy6gj64PVc+l1ZzSMH4BPbA2Lg3SqYABwVVqa/voI+t
jNrLF6lHLBdIaUMfKi6wbqTpuAjvXKDXcWLlW9pob4GCVnNG9tYm2OQRuY1MFgHP
NkpPmkHzp+u5YI5NOCm4yVIuXowCwyZYBZujIOydgxJdEXdAXp5TaLiUZexIjmi4
7F8fgAQaEOCRR5ukXWqC5aRf/j4NqBTVoH/yzjDno33Gbg3q0QAyHjGg1+cFLeiI
OS1HM97cfTqCRjiKTt72HhMJQwufFAQfjYma+HVt6oOwGDgZyb+tDi4cXw5piI/F
hrzKW5cJphep5KvM9KUelQcYyF1e+h0aFl9sXZ0eQ5x/7t8lLDtTB3A97HGEGl4s
G8PhdA+mSuYGQtp56vDFytXAxd92XgWYPPDXez4KUrsljkOS+y8wZo8LqYnu9sO8
83ffBUjn2XPIQF1BvSRPhPjs2jrOL1cjyPu8DX7pbVuh2pz44NgsmBr5eKxHc7Fl
0yUU/gNB6V8R/VpMw7Zh67+qrTyXEbae1bQziBfdGastPoKeddlVa9jSJt4jgR0H
LCa8jBfWwWdZyHhfNv5qhkZqKYl3UmTwlLwy/jnnlaVxIGZZVNA6axidgMjm3Pms
+rQHms1EEtYfjHlBpxp+kaf4EIxVk55uhwNzwY0G1QJ7zPtb4Qn8CNsc1pMeSVI0
4A7y01Z11TMKHtSs0o56nhkIKMtdkxEU2oQaGZeFmebBJI9WbRLmBQzpDQKCq3na
G2EtYBEB5PjH7CNHbLxquyMaZUPyELOJaJN8d6ADRPpvUC5OL75zCPkpy7McHMM5
J2Urnutb7s5fM2hPkJxuvUbAROF3OGD5PfxeQSfi89nmeWl4ao4SMprqp/1gn9+J
/30JH4c1+DZ2gPsewyxrFNVQqt/waUSTSI1ulha8camYZWclArR7TB8ypKgxudFA
nSaR1O1nUyTu/xEPJRt/MdBnvTHmAe92XXjFORZmJaPM881ECKAohpTI5m/Vq/4k
9Yy6pDCRXUwDcmbvoxL1pX3k9GuXL7rjvBuqYoVxATDJDz6oWAC0KoU0rXe10hIS
k3jpFzYVb7oGOUprrS64AoIx7ahBMe5bJuWMJltvgBjPPc+0iELBrqNUjJaQOXSy
5TYlUQq6DbfbNBgkZbR1ZS18iIM4XGkjc1ncdTWUbpJ/9uYgm7TQBnP+cGyKwgXi
6nHd9e9OwfP+yftLWNixusjnCw3EF9BIz7G6fYQ+5QU0ruJVWQHxqgUvtRledBxH
HvHoHRl4azA5bKdnd99wOcln9YQpTI+/L8tmbFWJcnRu3urpkZWncsDJVY8bQUjn
xVPBWst9sEEs7g9Bbru9EE6ASGwc8yaGSGnKPm9Rp2+vVeF1kFquOz5hbbQMdMv2
jkTZx4zXUmoQw4Clb+HzQSHFVUn1jUa+ZYYwj/Yz7LPILqstbMfQpW50Xji0/zEd
7NwyZwsxX/lpjpWWkCulmb/X6i+Hx+WjfoFQTAOP6JcO6romTVRP49e3LY/wbvvP
sSiHl6AwwG3adtryd8eldUzalZ2faPHwkBPb2UTveoixR0avCPe1ZtalfHjnJswV
ZypCbFg5oNppig6A3f7Rxi8j/HJR48QPAxdm+SRlclXe2GQIHTpCY8mibHxix6ug
dhfOLisMTYRt4uEryQX2pXS+ZDUZodZtbJL2XimX6OegNzsKdk2rCP7b8DImajgU
gwe4vBYdsP6G72xaZdBTmipeQ/C+VC1babI3jhiI6TdImyqMlkpHA/hoaIL1hp+U
fS3+eZFdsiVHDPZ8MtjIJl3AMUC1t40VQIybD4YhbRi4Xr8UUie+hIpSSViXncIZ
JtHXndT4ZCbjkpjl2mvAFryQDSpk59tLNaZEjHAbrneWqtzGqU4sZxBvbkiB+IVy
BESpWcyNaNAWvkZvLUpANoIQezWhoQZe45iPv5lirte150EL3rNGts6bsikY9xg/
82ll7wHGIumTPKzkycF/9fouN65RvjX5OSQD2ImpArTCDm/q4I3j4opGqrHA5gsA
f/Y5YsBlhxmfBzdE4+BXPUZK7gxQWJMqWxHyfe72o7PVNdKyiRaYNOyPV84g0bPU
Zo+QJLwsmEC+1dWbhkWccFeKUjL+NKYu/k5i52dKQKtnMF1ltPipH4/PONvHJLxP
tMIUWZWfhlg7NwmVawXI1Kz+kArGpFxQPIkpuEpMEzacbjh1+PiarCmM4uM6eSHH
gf3GJRy8NEl0ZHd6Q5EwUuK0Zn2wRjfqtEpZyMp9BWoL41fxbxGYuvH2cWogak+q
HE0zoS2Pyb/4T69lAWcp++o2qX2KslU4n0GFAOIRFKR/Z1AFBlVCVnE1z2IKTTYr
zPbO1T6YFhWVZiWtjDatDf3Bz8HRwKqHl53GxN0V8HAczWa/Grgw8bZTgqKDL/lr
P5dpHZF5PD1p8rE2fh7AldTl/dLG6pC5w9l9UX7uviV9xjkPSdNSFFIfpTrml6R6
mIOsKeDGcjJfH6m1oE4XPMaQevfcF58y5FTLG9n6OwL051rsl4dz+bQZ/K4iksOw
6TBl3xQzJDJiJi2YzBurfu05faCY2vF1ffe5xi00NXZJYbLjv5CUYVLT5DG3zeOG
xONFG1+dGs90qfOxZBx+jvmX054cijFVNGWH7bW8BYqxDuh6eV90EDoGNyXJQFyp
1k5jHRl92pDRud/RRQCVNGMcD47peXtUD4KTZ36zMS/AzOYiUUMHo/fnm130KS1l
JRdUPsOPH5F7sUUJyTZ34d+l/T00Cr40JFsoF+CZO9NmuB5vZsUcfKXK9im6L6Gq
svPV6D0PHg89iTkC/UjtfBpIcTLnLMVjYOpPS6Xjk5OZIREdKZ1RhMz7KPa12PmE
ETyAKvrAUbIecugKom7b3lf+BfzHmwgtV5xOXO1eeA2W9ckIIAI54euoaArw7tZk
fwr20Ibpwl4oWh6Lhy/gmGI5GroV5InYADEgXM+i0wUMN2iJATbdANpug1kHciW2
2v00j4qFarqsMml9MlDRhuXVosRMJ1tfxZ3T8FZAdLP/QUMlsf52ALKWcguXiVVC
0f8ggQmVL1HojvyMwKoIr6+1HJm0Hgy+rxekFm5WK7bB0+bCh6ToqYq+fR7L6v/t
i1xv+D6YLRZWTkXUI5Ow07oV7yzZw9nZwbfOgSUfjUb//JWf7M07LeHr/bWsXz+W
WmUrX5tFNVwqUoNXo0R4fYft8taCel9n7opQ6DL9fuRgXuNRNW9FT4Aa/14fDky9
jAfuAjN6tbzC3L7xv1rckFnYNaVb8nqdOH9fuY4co98ibu3WXOOK5ssUn18jUnbZ
k4eOrNg+j4flRJfBAzaeB1lLARKIEH/znHS7Nmky8qAM1uSrhDHEolqLGSWFjrNo
EBiO1QJuAw1JwYrwYmsIcpib0fXE6nVsrNwKDfmHXPfZC0LSzl4yipH4PBTfrmMe
oH0+lve60tZ+JZl4yQsP93kw2DSYixebd0Kh+OwML/EsDnJbv8LxSang+hN+QtqW
YJQzkbWO1RflC/9NPgVGghJrUDaurigJdHUiougO2QKw5Vk8xmxouMXI43YOvQ4t
09onvXhjs/8L8vyr2KZw7gXO1W4maXeipSV1L7KFARZAAjdHlskO5pxm4EDl6/2L
CNC53biLPAzwyxcY8TQ77RbbAsqtXtcSWwOVjBGF2hfaxV8Uy4xvatx+FaWobS1Y
/rBLKDuYILCIlNqNzPbZBXMF/WfKaaeQsohHUak969AFFbcCX/qs+5rcYk4XB199
xeLENDpjpIvCB3DtKGby1jB7peuWMQHk6S98BjYiWKFhMu87A+H0LJhoIdn8SQBM
RtL84tQJDjjFJXcPdYDsoGVCGlYL5NQgEWYmdNT6iPeVqLtLfPVuJ4NdelwXL0zL
hELxmgzZOZXIoH5aWuDQPRH1KLvlXAkVFfLYac5y4s3Bv5LPEPKFcr1WP6A6lt6X
GfnTb4nccEHT3+6xDyFjuc/VvwX3Qp/pf8tPm2+0UX5yk03NEzOI4g28Fv2WDW/n
myAdKXKjKVL2fK1AzfU3tbksU5ihohPWZ3dkNkudBZ6Ivf+JOggqsK2AagR6TUtO
c1GGuwIgN+G1jKCEqJ1YLcx5G1GYmmZyLT+MFddlFvOkuxivUIJWn8qIPg5TJKIf
eZ4qG1ReTpOIXeSJCNonE6Dh7vGnQHwrvZXPahzu/BHg296AB6DwYGZPKc+nW6u7
QI6TdrmfnCvOiw4JPQlaY75WjT10J8KaL2xohD5qVJEWekihjrx+m+DMDNAor5VI
C75WbETIA/9pGitnN6C+1mfg9VEYmBDm5m0Ei7p7bo41CX/LSsfh3BlY6bR70gDi
YjiBoIVgOH2Cj4PgxYc+QzqEHWAKA/qxbWc0Rmt20iWDroY1rsKG6usj0a0jjL4J
CF6lngdTWxjHrcrCI+/VT1tuHXvn/oJ3TBQlwO03chVNVcJcKjjFOpNtOCVFG9w6
Mvl6F9zdycr8HBZbaeYETjmpjE853HcdZ5a9SrDGQFZ1JDi5z2LiPiDfpkqPQXzv
yALRheHqjbq3bOA/8Np75u9qTvd+uXhLHnw2NHE5yhrEBUMqWfRGbd3A+Evlcfvv
oPhDlfxkeJ7f5Hzy8/Fr403Hg3e3Hlz8aSfATuvtlYn3ioCtp8ACxpxxxyWRQzML
rNXGQWm4EeZv2LTZwgEo5VOYYpQ9oLy52F8V1GdKm0Bm1sEGSqCh3vrD8AhcEEXS
U4D8D7PTC7rvEtrTr5mFzlPxT8Vsk9Gu/llvZsrgSFp+Q6XphjW8eTz0ZB9NB1IY
TJ3a/e/wsekX/bLqU97A//jCFxpNVZ6rVbSjPzeHPwEv4ujaftZioCRSph4XhD/W
yitAqfOs+BPF9d302uunXaoCZ1qVzzC1yJ4ZwiGKefarz7YvNEmP1OI+dA7Slj+P
uOJHLOkyYbYcbrjY/arR5tSH2hsrcHBVSd57VpLYIcHfu3NWXzDB1y14tG5aPGbZ
JsqtfFIqtZUXQg2VXNszCZzqX5H828+4u27Tq8TUbyia77fgVeLk2OCvgvn9vWbz
pK0s//5yPvvy8i4jtTS8/uJP2jOhvpnxmktnKkEx8KIlr4v/I/xuHP2FdlAfMiH8
tm0yIPzGbSj52dVxTrGkMoaAwfQYniMfMlBQQTar8HkYu2aMQ50Sd3nHgBuMUKeU
YQHAWGqCt5slgnFPJ+F3lGtjKgbLjZsK2T9rvg116Uiz3x9piwZkGNs0Hu3G78BB
0E6Wf21oRJNP70cP1mLhMdrpNCF9sfsLGijwvSbgubauzcCcOHZSmRV5X3KxOY61
TwQ1jZIV/gmWKp7Fk54MqnUVwjdkP74mdFVxAZ8Z4TivW+NUw/qeza1nh/IHbpYa
J8Zx1NsrawkzOR8mScQbAC9nwSfEpEEIDbiwUarwOXaOIv3oD7TAh/0lP7xfycsH
HvWkHZIzzoGWi8Y4wRoGYRS1c5aY7x9YfmvMo3WLx/eBe264XAhQHQ6211JQ9ntw
mwilc2HQhS4FTYy0M6JcweRHTMbmSuE6WNi4dsqp/MYQ1HrY/xcNiLDOWLLFigDh
pgudA1jeJCUL+nlhO5lTSd07kxmOCraWlCUIXdv5auc1IkJeMNR8uLH+cPVVfLCS
ivFT0+DIgvI+J6vpTcjKmoIbu0BHELGmPU62+CFobSafQfJN8dZed6VpllXai0iR
Y3o9gkHvPk3/e4YAKtMYUT1IkFWBKLcBz2XXNfKYmzJ+wwsLLjlZLf/4pjpPQzPA
/oHiZ0osyU8Lp9nA+/a+XDsRJMsHa9U41rUJmnH3kCsPks78jtSrU4RIw1AOoAlF
yAofjQ0VIxf+uZELpImW1vvFNwUDwJXUHKKKEonJrdPdYMzVroBvWJphlqYIx12v
HZAw6LGXY9dcUOVsXvEU9G32Re9StuvO7RmECgwwAIIgyfdswB5evK7CSeSVOwLA
qBd3lTCfB2mTj40ySCHjmQBIy8evc6lal34ZN/laDHZoxHR0qsVoX0ZhzGTcXvE8
MPKIZCeVdZ5lu+VdeSov7tVZHwJe6bsKWkioS9qX9Mo+GT3LoocD5zruNwWxyGst
jM6q/0nYGOq3R/gocdOeBQEFzVQw+WI6NE0F3AEMIdQp89ANhAm0/Set8xp6EVXL
qagQxBJzmVL2VokZUrLMR3TDVLnN47feTm9wLSs2MJDO6QVtxi54WLAog6qEjA2I
Vc4EF8GS0ZIow1fPjyNY8wrUiVedkRhE6nCN0DIrpFFolja2xd879RpYEzgMkDBR
8KEUaagVkN8tpcenvC77I0jPysZeXvSodya2GvMkMxiK4mmJm8QvP6dSpzYJt5Zb
zwPlHobosFB5F1oe+RhZJXeHwMpaQOxzRNLXiO27vieqtY4YT8Xu1IesZqT8zlDN
pymk1JJMnfJpYI/5dlqswDhNBXFrvkuFGySKlbspNW5oBSuvn7R6cqi62TLrrh1T
r4YIHhWUZ9uSWlvL10f6IXwWmQcaRRnGo9fAfl9Psx9ZH2G/e6VCnP+xRExnJY/4
GhTNRL4nu8/p8zCcd5eZ/GKrlVb5Su4muMwUDu9nsB5KhRuTbH7VOljFKk0H5UGo
CvwKkayCsFENgQzMYMEnOE7XdFsjeIOvxJd7LkpiSUTgwnGnXhnsG4LazYlzEC7H
iaPnUXVtioFLfv/DHk6EX7gITlK6A1gOKX7kuBcQ0BDBvOvQAiAwfNMZB0EPgGoT
QlKKv7a+7lFkZ+wVmJ2cnv91ybBoO04tTBqJ9R3S8ohv3b9xkj4ZHIFs1+64BDMN
5ZO0XabPO12MMMyJYpCC7ceQ3IkNLtQlfdXuZC6eR1NxY6BpruAY5zCzS2s424Xg
UrUB2wJmqKZGpn5Y7qflnKC3PzuMxLPLpd2ERJCLbz9Q/dkXuLLLqTV9hwZcg2v9
J6lQ4W8/EOoCQ6P/QnRsl9/+u9gnEv16HCPQaV9InOjusLxfzI82F2SB/i2Vljlb
7GEcf4aalXky08WXyDYXTbPx/Lk1qIakyxfH56tXt2j0CTLeUQZIXN46u3HhDVhQ
dgNREUmkE5ggTlLvoS2Od3QoV6MB2TyqBVl554lJLGAeXkmJgXFQDTNQrRJKcrFO
FMKb8nD4vqckxDbEisDLY1OfkPjhvBMSXSeGy16ARmE61pBhvgutNAek70roSsSh
8PO0U0/7iGh0byE+kQHZQ+ZViVv60z+YSoMt/Dzb/m2O87+0lfzBDTZv0fsR4MXz
A91ln3R05PuWv9WS+WnTshPsIqZdOURpa52qtYQR3JPIvj5RUg6kh/XyiDFWpOR6
nLCuMGMuihiiDvGi2ew+SYm2mZP/V/pq+rFfxhQ06/kiqduwG/1Fly/SInNN3ocw
CJP/dIKOvvIuVpiJmPpCFXTAp9Md60DCzqXLhXZk4MJpUkMXntDPzl2tg5u+bX8h
OGEPvssyu3127K47jqSunj19nUkcDEFskn4gv8DWQ5K50Q2XmskI3uzW85+RM+XG
3tRK7jP5Ow/xAL8sOc7+NyE5fIpq1VUqwkkAJNLGHi9mdkvA5csbVuMBAJ78Ki1P
TiFIQLIA13AjYjfBVTSP6iMHephC3pen6VDAoVw2bYZAiKxr+xYIaezV0ghpEDFv
+b1U6Jt5ZXu8T5NBqRMbeo/CCYPP61OoWD//Li3UaY5Zc/lh0xZT42xU342Flz+S
qoRZ4isObRTivf8seVZaZ3lJtWl8FC27GvlXMqgL3KgnlFfO1Fb07g09BFLCwdFU
xDoL0aW9RHuXFO6KSQZ7yumoiQrmOyebUsr8Zgh/KFDjVAbDiPYy2pY9Ke6W0TIa
F3TUIUyNa17eF2gLDVAccLQRfehj/utVnOFHCySQ+Dc8crT+yC280xPGP0xnfBI5
gPvMu+sP2WsHEldaMN7s0AvWsB2f305+Yg5arDMV4hy6BT4ASeQ+iKfzPakzjUsd
OVwrgEuj6yHZq1M8m4NUw1ZPtPgOG6PmeTkinHebIHpfu789VTrLVVGL3D5aqefO
LocMORsyNrqhZPIkC+6Tt4Dmh1RRHvwQCsaBahSjigqOHneFYiXSBHklgqNzqQZp
ZlPnAUu8I4RZjTuivK6VSJWlESeSnzAqgebcOCUnXAwVzWF2sTYcBC+17DsNmOjK
WfClzavJlJEAd9Fx9+08gvmbNShswEH3RuIKoRdpe0SQVXmkIXHLMNvKcOCtzh1T
YDUh5um526PDQhF9YbmiJeYrVtriBjo8+H+d1ss6gTFZgs3234S6cth2xTDubswB
3UwIKg8vAmRfqMST/4vdXUIKlc8bymk4uojnTJz4UUlUFX4MNOP2CTDZUpYpJ7a+
xl92v2CgRpnkZw0UsRIRyOfoL+Kk5KWGfVWwNqvfQqvbHji6zMPYT6WPxxtc1GRj
/HSgjWDrTzn5ye9j6bTH9DET3SfpwYq36An9ZQOHxws87mRzLCcsdWsXQz3TDutT
M2IDbJFssIybAn0aMM6a8MQIIBq9K+rLESAqFBTce3G9REeaG5IDDFvJEMaP9hmV
QQgrewrV5nYZ8Y1W/wW9NlpIrEFwBTdLBsmjIeJ0xyxedXLnUNh92cu8D6ZPFrpr
2bkyz+C3HUWfSYw63br2A/6Q+Gqlubh3HG27C9dNS9ru26r85VC2+yJHUGwqVRnQ
Cjzp/RsrXSY9yMNVonA5gDo27Mn6dhznryUc8efrNQNoj37uQlg61RVXeAECCkjl
sGWNOyZcjI0OBTzHwCX90U/2EySYKxST5ixVfXQTkj1EKxMvlNoMUnh36L3Pzj6A
ebRGCKdL3aDdzZwgmCMMgeC54x7rVJ4BtwxDYWlMAlbe3cLFxRElA4y756SOIdGG
YK4ls4Q0SQDe0Z54wKFU0v+KKM2zBjGECBj71elhTw9Pn1uJaBDWid/vW0zaazvx
3+IDQqsKO+v+cgHOkW7oOfjhpAWO+9fyJPoQ12pVxfEwabr6MBNF5Luuo5psc9k8
Vl3SYC2pkw0POyQ4DbTCaGdfXYD7+/tuO2kDWa4cP2q7dFIRnJJ00dxvnJnvGxmU
dWJkzDheGy/Hnz/9zy10gHRNJCtEJEcbH0aJSzcuvC2/ZeocSKEHxhderBomQCZt
IpkMjCXiZaIL9qlDNv0sEYn3jfAkKZbK5x4Kn5O+2Xk4zysxeu54DDXJ34b4Chgs
R1zFytKIZ3bSJ7MLB9ey83O7Oh/oZxsna38SkkGGPXQXmQOXt9UXPBatBzYHeYXZ
RokXH9qUD7qEPfXhH/17IkfCTa6sKgDDsOtgpx67ETlW8bB09nrzH9BonDvKxws1
yvy7UZnoxwyjdYqVwaXXQPBZ5apmTRM5JJMuB3dDOk8kBag0KloQU+md63uPb+Ls
p89Dlale2ZGoGbKYB4Q9IAw11rzQLoyR5YPcDMa1IjsvZAiX/3JNEbkuGRYgH4eY
MOyndPqfZrZh7ItSUy72Ih3KGhC2mhdD4wjz95aHxbOuR6AJ5KYCQmc96e2RVSAL
CzafSMXk7TI+EagcG0os7b1DBvKCtDdtFPZjNCCq+sbUVxoNg+xqif/QWdih0J1V
/k1He7R+pQvQKAyV24cs6dsZ4o8jekSfCCcgQVcgCPrIa6P7oYskXxOT/gLZRsWo
o1oBIdnm3OfBQ5UVADEeqXN33dCsoKRrFpWhEyd3TFYYYQeTwVsStrSRLEd57jFC
f2pYYaV4KgBLwdcBDt8++qH1bZAvwGpXJQERXAF9uzv6NT0VF0Gw1J1pBumIacAC
0g6GycMInXhiIp/0Q+X1nP9+07f5qTW2jFFnHviiVW9WyGQxt2zBGthI1ppO+ZgP
yO4BGxTx4b4b+ZT/+yq3HiaOcFl1W7AYCbCgHj5Zv2dSWTnX+uBxgJ9xA7DMrE31
VzlY28aXNqgvoluQNDKa66mvd903+8ZRUGXmpKvrKRE5CJqPhABhE3TgOzd6TDCW
vwIaAoqE74VC8gyLJCiGLjBW6KwaisfgUEO8A1woLNI/zp0sQOHH6fuNyCq+TEpr
usd+6+qA+jEv3iCzhUiv8a2HaIAwp9vE7u9XfqPdZZ6fuu8SUZkxSA2qUbe9X5sQ
4OYwhTbJwepjRbvk8EerPloRALN6wFtWk8NR1b1XtvP6dzt/BkrVqndsxBndwoiJ
RoXRlXgemacufecZPbQNuGJ4lSt7/82JOS8k5bqG/jjonGMosbI4MMKluBkSfqsJ
lVOLrFe1hKwj2/IpVIFT+s2XUtSY68B0UMuH6m/24b2c/pegYgTqj/IBHPGGAdni
M/s6CwNmUtrPtH3LemL4aOPJ2JjXbdXrcRUutOsblSz5WzXEsspRtAbCHd4A3Z2f
o7qw5uKoaOAF8vEUw6RQfbR1Dg0y3aEF0KV6JQynxBKB6v3aolPiuUgK7C21y2vx
wwLslgbk/vb/B2k8LSp7Mz9+nZCJE3hHH5f0EgHBziv/BcVVJ06nbGQviTOzGvOk
/0ZHmreUH33xt5C5iplBOjkfme0j7LNG7zKNDIIaAUwhPSwc1CZGVJdkWify+Vrz
A7Y/tgzSH2bGMXE+EnBSsczdANKuqCHWO1mzgesLfC9KfYgEUNRvo0lB+yAz/Enh
W1/6aArkBWb9LDjOVenJzmU03S4l7pUbycQf64eJENi7ZMUEVP+G4hYkWw74jXm2
D1fDvF3upxa6nBpdMx1PT8MqU/c3DCioEtWzbQIGcaErm+vuwKKYbWJCPR39Qzw+
3nrldLh8aZ+UQc8aH/sGjzCn4ZyIeUkMOHysxiy1Luh3KIQd70K+Ixn4kG3Y+GYR
NG4tDCNo/zxVRMx1B5lpo9BbmNb8AujAXxZjOU24R9LxXp77mb06x7qjCF1jGLL3
NhaHYcRGnYqiFPlBPByoWg00JLcAh7Lkhn/MQta26m3sKuh9O708E6zZrQ6E5z/f
pIx1X+/WWcVBk9DfR4XqKPibPf+qbifnD56kKyP73UOqqJRylrsec75Y9RGCzjQl
DtX9JexKkkS2mT2lcSHAsSyvS9et5nGuWQ2i1xAaHenaKb8SPTcehmrIkTGiuh7m
ex3qpFwD6rANZkBb5aXpdM+xvf8M8OIRar3sQvY0VN3HyXqGGGP5934YkYamV+1T
8zAOLqaNHj33OkmHRkEDUJxYEMrSkjv/eGRfKomTwdSvfqkbZhNFm4Y4BMQDYmLe
qdnMkhqj4jTi5Hu2NfPEe4yinVIC/JJa21ZtIiPYZiioighSKr4aaTbfozXXnebl
l2zYYQDOqZpT8LUpSMJz8BKTC4JTinsUNKoM6MaTY2wakfnjh7Yb2sgQOCWbKX9V
AW8sENZAPHfuOOYE4xyu/+H3snUY3w2wHGZXXJeY3xznOUXiZfKCHc6Y+EdgLS0A
JAfpgQbEDtknRc3kol0/evrVLtPF/02EwAnR9nBkDMpr6FNGjhG03PKeezoI8x0G
9HYiujKQmcKZVVTFfsYCvTP6VCFZNJoheGfZCYcq4paf2zVKDRM3oiTeM8BGhq3a
JgfY0PUAO3BptT3h63RabFZBJTQQOF3gBg3sZfAleq2FC1b9Owl9Cr8ay1xpQ5Hf
PWpzNB1XgG6jzsbWiYXxUNtRMk46mSxpcyQ3vizxkHvtem7mECWUd6wXELWQXSpK
UfZaoaqMyPTl6qq3FIh1WgAfEjKQBZVD0uBEencls5uiusG1efnOqaB6eu6EI6gc
lekp47SAWH6weybZ07JvuDO+uKnQgT+RlIlyPFrjKCZMOozB2Vz6mWrAuNTeZxf5
Fokc+6LzsJ1vH9wmjK+XtL98BSk450o5+RcnaCrdY0BKqZ6Sfn+ayHm7LoIZqkIU
a361ba+CoByKI1saavRYkvnXDCEEWA2dTi4LQr2mznhnSulrY9anjrBRFEuLyR1X
uoG0NiDRKinJ9lGio3cYj+34oNJVYgcxITz9XEXi7+rmiysL1PEl+huxQWLGyGri
vbRJLziZ+xhlbvhWs4QYnytSPlOhuTWkTWSXq9OkMbDeZs6FXSbL2vS0xnjpHb4+
nvolrtPhC9uC6OYhd6TselHajJiM/sJ0/hZLxGuTw+ULXHxFh81mPwCRAe6WvEli
z/3x6E9GW9D+Gh6+FrBB6GAEcCBS0d+53UKVyIBw1GdAXi8uB7NHuij07hAuOb8v
zPyM2OTm+7lH5RTrsvTSLqdViZOAcOjhlgRFDMyoEh5UKd4WA0OWEq9//PjYPAUW
penc54QAWXYbo0iOsUV+3zuKRxBslN+qdBEtGRm1k48lHd9qX3vcSPpxUk/ou1kX
MWxfjLCusVyaM2GNmDXN3hbGngPB0U+wmygsQK4XXJlSLBmQsOW0iv8s7G1EZfKy
syv1JUCfo3lXtUjDmh4T+20lzRJWqBBthg9rq8kOh87SPAcBbHcH4TNGNn5iMRqA
aFpNPtEQpaifaSr1+HDq4DHS7wDeXaFIotBz6H7TLE/Dr1u9/BMzY2Kw0SIZUcjS
Ro2HxdvYeqm/iJIOu/KzUBHM57hWMnff8INEks2XUs0aq94/vPSd3QQ7W9YignH8
SGE6jDsRp4B4SqAGoAydaZblwu1dMZvs17O613aPOxAsELXtTx0plZLFR+IHWX5g
DCDtJaCAk3EADQF9IPdpXYcmf+KP14pXQ2rSGdI46JrvIbdhRnkRTvrsYye4SbbT
GRdkfjol9cYOKUJJADGU62z/gYzfsZlLPrKM0vKcc1dFTQLF3qIQEtn9wS4xD0RE
v0i7NFpel1WOR/YIzIMl1jG4dvj5yUGuVZnbLhxQYE8V9OKcw07IAW1i2jt1ntfS
rdzu9MFaiVTyjhgHF2A/vwOXDOlrw3i38Oi9M+P450wEZZuyhbIc5WrZuXSbd4vd
EOpC9CrAJ0UTD3Z696ydSp+5k1GsHbLWx71IP1S3m4d0JVSDw3LVGgQRqUIQnPMP
nL/1fsLWjzFvAMCu1RabNyKhgIrje18czLagm0BOiVB5tbFmieOOStPkgpFdX6rH
qMEW0Gj/NkDP5sU8H+MusZXf8F668P6sfACjjPvPwjqQMF+HkfQGZq55iXOsLlXm
rnPagVG2U00/purvYR2Sk8aQFqu213a21geCSxdsaYF8zJ+Cr+Iuv3Y1/EjwIaMG
kSMWGRMJWkluktWTSxNI1hvHnZO1GCn4TUGuXPp2UIBW/I7wlTLsWwktJmaZP3Qt
VoiLkeWpcGFf2v+enUSMpeYsPYkdyHed6f7WFz9nmkcuLJxpGENTqiA9JpmWuEM1
Nq6bRR1ToKIcnpNOE5awMLJRCmgdt+Ll8QfcTqo2sGhoSM4qeXAMQAhYhYkrpFc4
SghmUyDS5OQ2TtbShzFw8KMEpD6HLygxOKytlI//Ozu5XCtZaDg7rWotqFkF3cJO
Yn3fanoDd91tD6fJ14LXeDpBnfjrKKDFWmgvg4X6Acd2DQkmZPOg6OSuzWlzLabg
FcaArE0XkQjLUpNpjRGJb2auO2RamZAQ0BZdAbQgn/wzo/2zI9BGskVMM2f/739m
A6O7HLZqQfvTwr4eKs9Cy3xRLcrNlHUrInwGVchiN+V04i7AU94XGls+AmPMkZAJ
MSg1/SDfADFqJA2Fdo2jxw9/NLockgXAfjgMZJG9njxKQQwsR5NkakNSBKCdUoCx
cO6qjNJZeaAnIw7v6d81/uVyF8Q01q9ou3j3pjS2cWL3JVmBrBMkSc+4extRqWN4
pwdv0gN/RMBR3RiHAyTKC5spzXoh/WanLVoC/vHkwV4/wg8w/YYDWZhuXGqpH56d
BqQpgD2ImWycP5cVu4ffdqT6LpRWzDpbcHNsTirv3nqQt93BC6/4jF3pJiKhBQEq
MyXGcioSR1OoxSsFjTHS03lQX/0uKP/SuxZwaniGAakHp72QCSkXEU8eqFdDM5rL
Jv/tglhApK2oHgaCB78Vkf2A3I0A8MHKUHduXvku9K/9gTRttsEIGVbB9ZAKL9kV
Ufo1omnskO4iM4YVloc1FuNyWZev5jXbauySPBuRg82a3iV8y6J98KpdTBnCY3Rz
BoEKx/xJt9EpsnWbVKS2MMnMyoiiH+f49c8aizHYJjrhgChq8UWmoEGcKWQgqFED
AXqD9LIHaKRp9WvJPWxpF9WT9Lc+ewTF+GnYKakAlr17AIQpOL8a4Zrqkh2aF8Zb
5pOKKE2UICP5IgUkEoPVkgE8YjZ9pKuXQte5wAznqziERVtoLt6wjJkSPeGFvMpl
GVH8fgFNXsFQJlgH+OTH2oZxB6MvzPpKkfqJ2lfKQTgh4Ls8LwKSYscsaf+EXLcH
n+0w2b0mNxOgC3UnKN4P2BQOSgBgOkO7RWrU6fHEMhkjlOKy4ITnHNfcoLbX6Qjo
iOttO5TOW/KQgM01DRYRH2/O2EzAdAlJzWa21LRu3gJyOzq96izERHOKZCvl5bft
ZA+7JDehVo3a3Sphv/9caX4K0KNk9aX4Aml7vMM9apYvuNbCBb932HXi2+wZieei
iAgm2V8l6NDlxzXVsJ9XHHOhu5rJmauXpaK1VJdHBWYrkZbkenwp0onKndDL+Of/
getK5+eWHNFD515UXd6M+PC0GmJ3zQs//VEQ1r03Xg6fEBtzFuVOBgy32/lL60Hx
/3bDiUz8aODVon+GCIMai9gHI4CF90DNTBq2Vy5kz626nk5FjtotTO5c35Fm7Ll3
8yLJUvcguF9uUzPcgbnWMRuQcyZpY/ncE4yIoLsfJXVke3G3WW2fbe7K3wJwUeJj
RYVnRPuJHAj++mHiMSpYPBwFul/LXgVlb5UzYhPAb8wfV0FQwXpj2sC9d9b0B30C
93Yidm+LCcrg+kgQRmoxkKF/cXtfwvBZxYYqxWth7syOppWDI8frCceKJ0m4k0EV
J7YpVNtmKDHWms/XLbPJnUu63IottOlnYKTpYElrdPQaBFKotbkYQzbeLwyp9ZHF
Nep7uyItcv43HkGObGZaOT9EQl/9PM29N4V+0j/2ohCC5y7DSOBfn2Mo09GdRGQQ
czXhlvaq7o/Nnlfw1DJZoPHG7NzLmTliwFmoS4zFciuw9LK6GvNXSNRd6K52JG3Q
Sq2wSR3SGnzXZDEy2u+Eb3VrCrxte1SN3YmkzZlRM8p+sPtwJkauBKmGbQdYdkBm
M8CtyeWq5wtmNQdwPkezLT/Sw7fIw6BzDBx6/WEWtEL7oXx2te/GhPCIQF/tdOQ9
xDPLUcLk/2ybo+2azHUyPlCY46lIVl0owpmPfU/KwprewFDZ6eoB6Ajo+j2dUPsp
jY+tkdnbM8uoCzoQ3hRu/WXZiQy/xRovvyJ4r6YIgBtelWYEZKrHL/Tu91hATx8G
QTUWaX4uIzynVy9qn/EbtuhqI/CGBU8kDmH1A6y7uFo4WD8juWAc1PHFyC9DRB7m
/4vZqra5rITKOobKqFT3W1CeiTkdh1e6p+Yyg2Kqalclp5m/G73WVNdvInMqbN3u
AevWKiTAhZ9MrmrwWG3uYsO8HN0F1Jc/LZewhtLEmk9Dmx2OXqEMygC2lWwC9I2i
kTFFZEssL1+ZMYv252q/ToyyimJhswb3ZB8OfRAUsfdiODSw9i6Uk1yRorRl6MXP
++M/S/uG7HkyZT8Whf5Qg6k/uDe7aNjyNg7iOK55nssBl9zoJ7YO3htEIlua8Uie
JxotgXOa9BSqUcNo2xK9BE/F0wqIB1HqEzkylqXEa7nBVDQQ22VlitJXxny9Rf2y
eMGtjyo7dm941iCAH/prcA8PMBUFmxaYMmaJEEBw1z1bVvgYVP2WI2AnjmNsKotL
wXZLmJF5qrThO6KWySjSpDpOQpcLMF9PxXOh6Ht34IOaRZ3DRbfUGlN8zENx7vMR
dYM9SJ5QKFKWnV9Q2OH/AKxI5LyzqzFX0s0OJS0INGSBUKGL5v1KEme6uCIQuaov
NlbebFu2YTAHtMYdBtJyaZgicWpaKLoFbC+2vobfcOCo1TNpSlSDcY4E6d5aIcFz
7DYtMWy6HXvem/705bsh48I3m5Cnk5BdB+ZWjwuLr7Mkaq54VBWhQertTtIugi6M
WzFLhRJq3Nqgwg2dYwB4Qk6HAbXjomOXNpMz4yErbaAAY9QAkh81+hXIHn7yLIoh
/3Ek823TCnIu9JVD/Tcc3ofBaVEdEFDXcIMeBpG1cQroI2QB449PGMhglt/sSiYT
IreXHeXwGGHbQyqyRLEefgY2ZwxSO3tWmbdnFmCu+mJ1uIXe/z8JZCdJI0/D4wdm
K21jUGapZHgGkMfrTibKZ59R/W6xsa2Fqsl7v+DUp26Vc9iDTtvsHbg+9W2zmEMF
lj5+YrJpdeXS+lHYei0oWIq9OLVvjmI4xd3tNu5fUUnYTIx39fIOKe7wlBv9WcJj
5P7ZsE9kAXxeQtta5WnFEw+7dTxSSTLUIwNywUdzUBBGnNrkgf/MQCSzhvSR/tO5
wV9jHQyuA82CnwD7P+Y6iyZunmg5hh++YwM4Zx1HBGqzJGNC8yhxwVUuRwRQ2EBe
kaum1Z6FYJvu9Ce8HF4tWztqdvPsl6DdUKjXA0jizgtUjIWmU1o2tI/8sLV2UZVm
2hAzk+PeXMj1Gx8McuiL5uoOFGMNtrqNuUtCdERSVIgF1dTiXkR42KNxWN7HicF6
X3mdfjP2clcCnnmsugmpeoXee9UN7ESgQPZUbbIuBXMt99bPkVQBJsropzFDLtQn
2edYf1HvUJ/iplrFWBePATRs5ownItxbcjSA8U6Y37v61Yrocxg6HsEqWmDtuwnE
fBfhShoTmasBryrJuIKPMiM18+pwqzQZcipNO513WDJaHjQ+qL5FUM+Ei3uwRe2I
okCxXFiqHhualjlrAcaYTDp3zHYy23bt/T+VRIdOE1uiG5yho9eNIcefW3Y9ghmy
DMsv8DYXfJC9zq+rGbp+C4hIL2ol/xK5EJlmRpoNF5UeQLb57ZOosi5bLnXUu9Ua
fTIg/82crG1I0s1t4N+eF/TgAQWSi3VyK2pbugo8IHn4hklw8iRkCeB0H6/BdyOq
ClJYgfRDBRX6R+wH7WcX7uPlT0KD2/waTpNjwt0GophrplfOHEeuSLwfOkH//aFn
nng8YqjCR5+2PZsPZKlnfm320BBI1Yr86PLO9K8bQZkICicZ+C04S0/ZcMO3EhUN
zOmEnpK1N+r8VHBwiOHGvOXBD6FTVklYZ32/+HzBiWeX4SGGE4JLsBOBknozumbe
tLmLi07AnvD/Xc9iJ1gGkaBVleDRTAitVbmlFHK3scHOAxDDgBNW6+WZnRzBEQx7
/5BxqMlFeVNRta/0n37gFf8u09uaUv8nMk6+trAWG2O0bhGOkpFnzlteX5bt4bjk
+500az6WsytMGUC/NpR5R+cIjX1djJYpwxP7W/jhghFOmfFOrF3NioOGSFFdz65l
0In6+rmUKZOzArmVwepNHLYhyvyMH7Jbn/6WCWHor4lWJEG721VxdQdO20PJCbL+
BNnRibsDa4HH8nNvM+x+yB0ocYMB2HHSRO6/X9OltbecAg1RSzxLA4taE/NAzNKp
0gcE5WCPJnWtOsFEbADc3rGQVrskAzmhcMe+xej7B4sfMkB2L6oGBBqbRSYsKjIY
jjt0uXFU8qNFlQ5uUPrlX5kISawV1w9gXVobsOvm38yZTMmFBZD7jC4kudIzZi7u
Lx0vzUYp2vBoRHdsR66S0H8b4Kw6dsNjujYw+bWUhzJLiG8kaKwHxFNU8R3RfUOY
xPApLSae5sid1r8xTCWxOrmsM3K2QikYCNBmDJy2i4941eirRo1eONM2hH3Mepoy
kMKGZi/SH2RX4OiyFCGPWQ6l7wYRltK1ynNvDQwO/u0JlpJUfMh0B3pdgfHryprA
6644eMFptAc8SNjXxRrDZ8J6KlKU+SCl30ON0nzxhoswZcJb7H88Ku2f2bC8fMK6
Sk7sKJofGwYC5HGTk/71KEXYJpBfhagLAY/pCnEDiIIV4KHqY8Z41Ogj+GWoXjO+
3VE9dl4+dtoF9fYV4igf9P6lxvsgN/o6DguFcgFLlFvv/DW699+tV8QmgG+8Rp8s
QKFEzP9RcovrgtT5EUuzyxk/INtOxFrfGBZzh0XANd4rWqeLdyTfnjtOzfMKpruE
Q5RrjPcOoIUmtFSln0B8A4GcnQu3R5dvA6crkizSfTD0ON9Re3M7/j9OXVXmRSfN
FMfb8pD3HvjLEdkhIjRaKM27JZ/WR+OIO2Vi9+S2RsmmZ1xRFCxArghI4LxUZ0k+
zWqtVNvj0uK+9Y8aW6pYOW01QvQ8vPuvb29yMEIzBbTnpv2V6yHQhlvlupqtbQXM
PeKRRP7curDjpXTdOuUsI8VRimG/ma2nmfoGtE6jylfnj04NlwYa2Q+hwtgjlMsV
Y7AqZ/fHD5MKPHsC+skzltvm4Y+eHYG1wLUmZrnWeWYbqGv3WxlbLITuOiAoTpju
nkAw2tHDUQ9H6Ujoi4LiNE3QF/1Qfl/KhqFHZZWPq5Uehr9Iq0NX1yJni+ofvd0k
dgk56k28Wig+YpP0OIkBBqr4irvacMP4jL0asfG2jMFbMCPRs7Cl5p0Nl4Bv4mI0
MwM1qsMpKbXe6cyy2YEyeQ+AMQPSjMcfMKHERSKdQ1TCtk07mI1ANovFVASqBIrf
XrqItOF42Cm/1DnWX29vexIibtTKv2U7a40hoAwoyKuIeteAf9s71U9BeTMx/D4o
wqNs/+4/vXi5Fft2nN0l+fLXEPgzLtvSR+5pT+q+zHnsVIn+A5GC/Q7sBfrfBrGP
cq/uUonNsGZaAkqhJSkMq/cjBEFEnRBFbJaNikdOWSOj4n7Y/Z7jAYPZW3O72D2v
yYEvUpSzVs6I0TNBFNxwMCgzTuQlyGPZBBLPTaa6u0ohPJMG78X1Iv5RIUau8RmX
NVb1tfUav+0fvnDKOVJ13nol6wVYoLTz5yLNr5XYqvdcD6o2F/wL0paifm+F2T9+
AWO4Tp4RnrLzAIA04jtrlv5Ze5fcixwFaRFtAFxe5qOssjGho31rXqEB1xM4f6pL
oOxhj3nV0R9JFrC/4ghax7GzpzjNTeR4piz2ifyWI0Srip6yGICxzjwJdXmSI5At
IYQhDtUEudYG+HeJir1h+ZgryIzohtWqYnqmUWdhPP3uTMDHPgHLwPjdRNnjEqbQ
DZrOV6U/mkEmzG97YC/WvC8VcZKaxS/3xRWtqCGS9Y48Dmm+6jf0xg26bWCG/VMa
UoB0M6x6y3flg6A+maLGhK51YMfoLc5Fi+SdmsopqpLefoJjEuiAoE7TgYmmwOdd
HJkALfPGt5BZngU9gLDcUx/FGKm0hGj6R4KNggVWSo3nt7iDBA3LFtOOwF7D/3rH
gyc5i0R3ure308/ro+joABCCLxu3s9KAYMlyPQeh9TLsv3XxXGM8bbNP/3b5IGX0
sgLpNNATwnVcoSZZ8qPhs4ej5Hqzv1N7TSy2/H0wTzvvQ+HJXS5EhvAJ1L1+Njso
RSX54So1X7lEwZztxfIb7q2kL/bgyAJYpMnAaSZpjQZGaAh4gBsxYRK6+MmJevCH
3qxwNze4xMtD+pLWLpz2dySlPOcRF7GPLWsi6P2YTGOn1m05pdzubQtspq36RRE5
qpda2t59l43g6FprPP8pO0xmGi00NM3Rmm7jF9QXXsSjyAEbNBC518B7G3MV8quw
/Lx92FKkJrN7lyllPYqyv7uEbC2w+LBLZk2y98mBKgKmKoceERzG8m3MVcWHp7Fu
gITZaxc91Gke8gjjJrTZX23iQa5UM+fA/KrmhPjIQPRrgCNtctgwappA/zIRtB/g
KaEa9kTAlkjZ3M8LQgjUHLkJFRCdEo5o5EWUQNHoQzmjBI56f7y1AHz0R05GfXQS
TVnodtfa4us0YwRVHF8Bsy2UXsjjWfuOkxms52WkeOss7h6aPv/43HYrIRYNNvuT
bVZd5wBUmIomZpShjWMFVmjPPSu3nNfBh114ZZyf9S0WkE6f7ODRSRIKE/eTsNZ9
Y084IZ8FGIfhfQbfaBsq0UYlQk2FSbWBObgdRKR+CJeEOCdzGhTVms4fwA18KGcp
h1zqltHJxAWzQllFcCwZ+4oBC4vP3Rio8JRY7ol8f5oSNeBoxaZzRBlLngqkgWCi
hKhOvT0UDwN0w40pGf/Jsd5+y5r+n59LXUJSuZsi3wj1e/7AurbtqU6SS9SBqx9t
GEEsm9vnGUPXqXiKWa3CL8V7T+dMlTuD6W5qp6uhN8pr37imrJIHoSopfFf4aMlT
+es9aplsIQ9btTiulng/WqHoebut5qWJfg+G7seYP13T4OThfGJPZ77QQB/c4hks
O2Gr1VYUaWF2iekk2rzOqrW/coE4CXYqiVl8gGXfT9IChGAi/zigEPZEk3NYXje9
F/RFpmmqQBQoFpx+fMHPCnnTk4pWVNmg5U+kxMWA+lWVioyloqDkwGbtw6x2HzYQ
JTDzFgrss8p4AVqjamWsJNf4GEDCMA6cXuos0jd+pGDb9gQqT7MMkBSVRNM+J5cj
VILpOrLkk4o8aWXbv/Cgl7cs9Vn+T+94h7xEWIyrptBxMi0MIE5R/i8x64wtW+Ol
ji1I+FNy1SeqA1xDASZp4LTzkt6UNS/o1u1XBeVvfVom46tOpsYj5b5twFiqnFqS
8EtcF/6sKvddfEj7/iriN89h22vrdqzpizqJ3r7GeA2Pu1kfQNdudq2rlldQJ0ZR
gqjjMafiQQT9TmcpMQRN7ngTH+dT6eOSY3ke15+j0JNNAIfH+trZ4tP12qIK39cA
ikGytAHNOZc9DEhFShnuuFl/yxEYNakQJ5coxO4wc2P/+SNSlQSpsE7Fh32Rb9Jr
0XlheuZqBX5GPk/YmeXMcdmsHnkQeKy7Tyj9Xqfy8Iq3NUTAxdpKYcaewtPQawKH
As73kjeWzrHVsINP8JK1IEjXuWNSXGIefNFAPNuBXh/PdPmj1dRWR89A4ARTZfH9
rHDtQkox0R+Rk9XBUN8MJfhpQSMBdAiZ+/flsyZnoBJ8ErFSXsa6zlEtuRRu+BRa
rEmBYavA1aB3oEJQUFGAwbqARJe2k95sciLwXWn+gAX8bp2fuWv5VL7yN4A8kRHY
1J1lfvHQ2OoENS6fa8ZXw+gzYG5D3UA10Dow8yj60grusdo6RT5dZykETzUitzBd
ex75TpLhBkfPCEx9F6Y5ZfDdjYo0ee447tHNSxinETvWlca1zRRwd83mOVHyGF6L
wIfolCaojSFdVH1TMzvjWv4gd61CjGs0xclfiwtvL19SIFhnOolGFbXCKYloZopB
SPncsVRrTYtn9838m9YNTKudo/0Ab49HQV0/502lJDt3YnpUSX3SoDj3Dhyk/I2h
Ys4WQ6q0Q4aAdgXGpHstUE+Y67fmhUi91KkywBsBPUUVs57yRm8kIlIe8EQ1Fepp
YRN8HIPlYAY6QfDAaJwA2fcNWCCTMXXO3lv1yiBtBS2jMxApaIcAHpr7R4xYhTvo
NRK071V3b90buDj0jm/q1Zk7kD5o3hVb0DqLcyFJOHMOe3tH7HIZJ4dyYNg4zHrl
RVSWG+F0utMbZhUywKvC+fZECQ2r3ACOSKaR0K3hHI2ZCLW+BgBjNVRF1wlO1lze
/Jh66gTJdbsQdYJr+fd5pgNKMLCj2Y6+VHwo/NZz6qZ70O4+cGL5b7QvrSkZ7/2p
ZZA68WiidBBImcpieGT10IrPwg70g20whWF/4RttPShssrLZ+YCk9Rl5RFE0Zjbx
zaUjQWkVxrV1HChGnB6iH9C9et9LQHGSo32Dv5G/jgBrY+qBm8w0whVeqbH0zDXv
RZmzrpo3AnqhsOXzcxbs9pBB7hRHQ2O9XywxcTN9CBKaqIDcrz1c2m/lONNGQVd8
27eB38elL/Q1a5esNsS6SP13bWIUgyDYiuP5w5umojc3Zj4fH2XCkHBMNS+YEabq
sGtSrSHtzHSWoilsWILhD4g6sLEnKLaaIS7qkwcqaQrU9hwZllsoouWM3GEJmknT
m0AukZ5mP2B9Xe4EPPpSt7ytwY4NjfTGk3SGAJUHMtsC6ETfdRJtVHi3mK6aMPif
YGzrCnnYGGjzIdgCmsghbTnsgLcOA7GqpAdQbYKNIzKlwI5swBg2nYAja3mRj8hD
8fMtD06z5tdf77KVYK/VXmjA0JCTDz7TxmCqu+xIHtGbkDGe/wiSbP7zd1860waw
7If6aFbH+LSrgTQ/dhMawchaZ3udFkmbGlWDtJ3P0ipI4pcYlhPvDUApklm7T3Ij
RqfUkMmjUDryZeZDDN45oEuOxyTnOQF2xUYgBF4/HQVcKgapK9mk0f5/0h51Zy9y
L96fDd+iRbRkWOAYC3j9mBMCg7laR8nlYhKMmp9orE0MCyJQHdOEDXGjvjgvL/oX
JJx/oCg02mUz8DcRIUSQDlaQUsNPbEK2KzGCbvrN9aRyAM9XRjm4ktPAKdsVB/QT
C1Vbcjm9OqUAyat4oDupO1XrdmmuA8tysD72ahtfobK2Gh+QAaCuJ1L/lw0uPlP0
gwX15pMf93g8FI7qF+7jMcBMrJNn2aX8vFfvB0BDkkQGAYo/LZnkFLh/fFGX1uvr
er6fnn+13udCSX5YFYXxe2OzswXiBze4/H5Vv+YNrQLOxtZT6TgywPExJ1WDtIJ9
BcfL1VPxO8JwZbnEO2HUls9deup/5OKZOmwOL7H7wdT8qAs9Wf5HqzhhAm19al/m
CfRJuvloOLVhjI0uIwtq/Kug/shu52YVbugFk8cXCmP9BP9Fx/u8DwGdw4Kxw3tG
tMdPNp2FcpiN3HwXRvjPXiZ3EgaavxwGdrsf/kszcQHPYm7coKOyo+I7IqGBNHLb
DPcSXLpX0AbCERx0E6I4aqbBR//iJUVPb267bsqj3gB9r1Xh3Le10g0iwW832Fus
226FwN6ZzKTybUF6FSd1UEv3IXlpvMj3PkagEs5XisB0xJ4dTdQDrMCrLqD5Ji82
IQ2ab8wq1emwItPVuRJcSPS1fGQm+ywiZxrS1d3iWXqGxGVbbaCbxkS4vMSeY06X
b6Q8F/VecGQQRBNaWuZzKvGHVQgUOSETLfkrRjqc+ZHzsWFPnkxIPScmb2rwPJDm
REFdxPwLytoGMWf8pmvNBZD+5QiNO5P6fW4eYrEXJR3Qie+NDUfEGPkvierVvxM2
8URIEqocghRVl7MP5wBWWZcqPA49BJjZqKqv/S8/e9s+YXxJ1RCHJB2FTumO4UOJ
aiqXhh8iYfQ/0fCz7r2xNunpTtFrBoIYmmMTLAnbGf9diyraEKxhAuJ0EvKEn/83
RN96GW1m+NRDpKCNYXuPfmV6QZ3bKiaM3fx4D1bOC1XH9VVyG+VNUZSSL2xs0iRx
1O+AD1XelXlgaSFA01rN9J8VttgwKgFFkqeoLrVXzGZvNIf4pl3h3L8khL3N9o42
qhN2M+47M4IYm6oMYQzTxGPc91IKeZNBiz9XwBTVj45/WhOJM/Mo61PqoPeAvzNi
61y7xnDBfBox7Ttq9GrLvgy7JQfGHfuC5GYGAosDvd/LTrhjQ6SXqsHiT2f/fGuO
lI5qsqkoS3KPKIP7xeNDyJP0KjqlsOfXj4vY7oaziiNlATfzwPkVoS7/tL5uQ6a7
t/snfEbb6+sPhChgTQFQLzo6IXLyBbMCQ34hYDJPWTsGO3UkuUzxndWHEeEcZIBj
thrP+hGDjupeD1d+FVzRifwd9TMbprtIkc33FL1mgLj1OlhuKnpvRa48UuO+t5Jz
obLDoEFK4eR6bQOK+M6phEb/FDctahJGgr3lAuPPAWkYwd04ejhfaaSrZTLAeveB
oNy1Sr2iL82a+MOiDMTEspprEfWLFKBNkq+LxPc+q/1wSo/thelw4XnKSPcJ+zkG
fzuYwP4hd85DOwWCAYgn/v15KOtWd+nYrd1+dpRDuyH2ilb2deP+IyE7tGcukweF
Pb3zZX7+nSZFwllFgoxT/2du5Mq0R4OSn2lcJN80K5paKfRxQ64FqckVLZD99X4F
4AG6UCX8G03C3T1nQGwsvPGryB9H1x6u+WvFmekIGumwQZJL9lxiqkTmZE+G8+o1
NbUnZNBpfbU6CSPckZ7jC0tLtgHAoRbQ02YTgUClT6ylTdfHhRkgL1VAETCf/AGW
FxcizBXIQDCaoihIjBsfRtwpVa+aMLzKVYD1ia30haPR1GnQQVjACIxIEgV9wsaZ
mdB9FjSBD86WZ8cGYkbtlsNuzF4bjktoEDBXo7ksBPFxOsrdSuekQ8nK5u1Tv7Qb
gPzAjTQCLTMvnidt/caHLKaoWt/TwO7UC0dcTlpqvQe74rrU/JefmaCZrcxTHxse
OxXFUBVkziYQzh0Vyi9/wm3GMNGgimGnAWHX4QbnSKlRrSIe7zxymYy+djMKzpoq
xQLoZV1/PPcdJcpN3C6VGFCaAECXJAFL0D2IJs+Xy++ZcELAw9LjZOXfC1xGRcYA
4dy6hX3Ul2b2W9KhVqhA/N45eJFzsgI319At6D2bMceWWc9RLAPyrdCcMfvw6Rsd
FZgUEH8mV6QGw9+FvNgf5yNYA3s7OPQNhLoLmz+mGr4szDnw2vfFttVpE2Zwm7ML
hBk4xZcE59z/v/qUWbMKLRrfnPnI/rAADPEeOtNZBOl+yj75pvjbmO3H2mEq545X
HVXUfcWizeUCjC3D2nrI0sEO3VD67Pr9jMTvDH0d7YVshvGl6cd3JuNEfdkFA5T2
GMq/W0TjknIJprag2vsCBIxMecXC9B2+DCUJfKo2zfmzDmfs4I/v/7zlnlJ4FQ7b
1tRCOb+5tBZyK5lR3Z/DSapTji0z34VeAL/eXDDQqOr995vYK8nb13KBjIvcqVPm
GHascubfC6ncxLGlPBePRLHxCdC7a/CUNE1FLbOpkiiRRfNI8yAnGQX6M7WyfnSn
P6UgPasCvK9v2GG7g37AJmqy7H+1ys/yO4WG3LFH3Y0mWfOelvK+Cpj4Q9evB49I
OdZxvN11nYmVNYmr0Khq4pTzoIsuqQKOMfKupSLDoF8cIopzDdodwvE8TDqgGtUe
Uh8MyK34/75KHv3kUnEH42MfRIvttl2IWAE2yrD0ROy8GdiGTosJjUqT+UZj56t5
k+OEgE0DwppOSlSqLa/Q4S+TnEV3Z3giDLByPP8bYRMnIj0CAxxGA9GZTlb01PP8
hAtjdcA0qbiA+CT/X3IwYQFZHPt32oeBDdU+VNpjaWYhPTmCVe0a3VCT6Um9Q1+B
/Qgc1Fjx86QTDTeBGRwnT6Fkw0nKaznIT8mrN8Tb2Xy/q4BKnn2GLrsTX62FKim8
M92AVcodGRtSYfG++y6Cfvpx6o8/xpu57y3JGu3WLvgRU2XbCSzzYEzi/DRplOPl
pAkLz16JKOAFwTrMlGbFZnVnK0bDnHgygO7mJdfj9V5TAAbnj5sscMiP/jOQB9Jd
p7j9ZinpVNm4I5cz1bxPxla+EnKASnNiww5tnUBgcLHsUZA/2ZeUUBKKdZtTQBA9
J9IRmfj6PocJs61m2jmeQWxNARjfmoEYgZsQQLRuZCU8Rd5SzapvoF9IWdMWRk4R
CeQuILd36BryfZuIx3dy+1VDXCjjfS2qTAA00dPjdKjQMjb2CQfWjFWRNR8YzNA5
ZVYI5yAR07ZZxCctaGVSx0KC764OhKp7lG+hmwirrIG2SPCXHdZQ6jpBnDy1PH9c
QYBDJE+WjbF4qoYFglI5WfMCE/mNLTKTLxESlpMqTAsIGsXembEJDkwozzthbLoH
fRsAKBHvAeyu108VU+hVBuhHTtlgWMH/sRCy7yHstAhBNbTWTsDnr/Fx4W2dCkJQ
oiYSu5Odk4cP7mwj6HClK+tOrADMLgEGojgkYmS+jMGSMgPzqwd6MinxoupTFy+Z
Law6G+ADud1xOqNn8n81ArY45n02tl4ChDYU0GTDYp1G34bnTBZRKeelb9mWlPQO
tQ1VpH8kalMNDA74sxc7Hu/mjBXeb3LSwoVyNkYHYMqCog6gpgPeQ4ShNkQ8XONQ
yVIpThN0MjpMsQsHiL+x2FZJ+DySNI60t4s+koj2M1J/MLfDf733EVS5XDCMPz9w
poJ6scvLbc+v4flZ1wc+CJ0YFNDG052q7YrWaSI/ftUB9nQlr3YIUFwfddXFBU5C
VW3mvdFENlFnFH6ELlRUt9kNyfY31m2fcLyYR46Kgb0VDusNZMNcCqTyhnK1Yk2i
e0RctHF4CwzxauLp0jE5m1Ekn5EIp8Bnu1Ddxgao2I9+T45fqGPDieNaVikEdpig
McGFVsltPkNVpOEq/obN6LeyGpian6tsbKQ3VHi5LzMW9u03ZGf5k6iOFa/NzpVV
hwXcGGTB/tu+nfWXS+qou8TvYsrQfh3Ivbxmdzet5caS9HtZ/MyCtZ5OEx4fDVJy
Rsz3h4/Cz9tLHPo+pmLhD9kxtKJc328glTUvgDrb+wny7T/dDOP85z7FntBDTCul
2jRHB+BbdOjnoXgPdys7FFq39cYTyad37krEDOEXqGbVzRLP6wXj/4m0vb9AQQqm
69vpd5vrBlTyzGgO7uXkxpP21hiL8dw1pHOoCjhXiXQi+idtnZOmgdQPp32Ys9i7
PtfTYT3gg350N8QR53cBN4/aHgH6rmOonlHSCNsOI4uMLP8HYl904Cx2EP6gKMC2
lwbqvUEbJrDDtTcQ71aBikHO7GRwct61NAks1N0WTApItAdvm7ENyqgztoNgw8It
RUY7Dgob0DDdi3qcAzYdWsrWkiLKqbPCzdJVdY55mMrlvz1MZGImefJLCLjyjabH
5OZg3BwFRNvLiJr+lAT7n2uiumF4vunUhfOc/xB7qTV+ktdSLOWsyzRrGGOjirdg
o4RQ/x9KIech/TdRwmNKrjwUNF/WO1J2jcLAoLCh/IkJNNzSmuJoQzS/APIeTLmU
0PMcbSCBfJilRl1OyKSaDHETdDkByXVyqCjRzQbie84h9IMIh8ZUzyIkf/hvt5rQ
NFJoc9n69NYOvAswNNwv+MTVEa/xw3+ybAZYWnIa7PFeMs9AKuhiTIXSIaGXarj9
97gooKcQOdaUqg+ibIP0gkT8UD5+LIlmN0B5VEOi70gy5i5D/Rd2+QSmYK9zXaki
tphuPYmrOyC/jDV+reKtyUHtiMiLS/G/I+5yJ4xgQc3Ag8OzU+k/szPTRWDt1FWw
MSomefYbPAyREtw7B7efFkMrZxQaTKtXkU/3B4tWWYBoRGSEOBUdYw60zSTCHiqQ
PJqgP/okvbHnAUkJEdXDOsNTScI/ieObxcy5IVg9XBjFh/F9ugwkyNwWqBNK+YYT
e6ViLjYGEA7J7zC6BDzRVuU0zwBIcJS7kMnn5ZZ2BnQ+sFr85Iw/MtZu9zJGCTVW
GkQvnbIIXgyFC4Lq1O8NtZE2vzXmsGnfiIxiaNfhExJQL/qPTmTQVlpVYBbLeFpw
uvl4AbYdwhx4Hpe//DeqnG4xnZfN4/x6xh1NhNUGHESJ6EA4kBFD1LVPSu2UhC93
KoznPNmgCLyzDqrZRqHyXf2mmlZF+E+FENrzzgrnq/vNvZUOjSo4dDP5iJ9S67VV
ip2Ld7hbMruGFKLtlYjMlI82sx4sO/kbViRE5LTUfUDOgROzANMM85MjooIQ1bMK
+XD9Cfvu2hvLDdZZfC4A92m9hCKyn4Drf1ITYu1SZfmjlaNTGtAK/mwYZxIdcKeI
eUlIgZ4ccEXIlqL33x5DdZR07AKujl3h6JGoS6z4vsKJt4w+JhGE/gM3zoKHrlGd
gDSX0iOTsVUWCwTehuYqjVctI13n/UODAz8y/q+sT7rJAltSM7bAS8WICQN8g9Jk
ZdM33o6l6qsBdxPz9EQXHJhQDE/jTa8wYx9ymjVELPlpF2XOxqfh3b2814w36uc0
rZmcj4wUCm+fin26M9vqWYSuTlfk7spfVvURb4lxQh9zIxaFJ9puClTGiSNWvZOs
9GtPkXm28pZXlkqDRU9HODJ8vugl3QxW5/h5ovt9kI9eG5Icv4t3qVURmNjhyfzo
FTHfPS6qNfFfUdwmHDKf24m3QrddkOY0qi0/XNYB9vcE9kY4Igq0ei6YF25gj+ZP
QLoNFrrZCv5AYqXJq+tb/ZfB21wYT703kJ4y3INZwJF7/4b6waET9etRa+o8RW3h
h+u4ZoJ5zoSGa2P5GL23uR+TpC+WpE9OdN2n73iZRYOObfOtMcE1p6O/uT9fg3L2
fpRmcy4roGoOBwLMSPX3U6E8XGZGn5xBZxxeszoAm1P7VOhk5Ls1rPBSOZgJeBme
z79IspnHTz61765H85EXs97GbEYdKLoh76Su5bdwb0/1UvPO9cwBn9v/oNHiWTJM
PMHDh9WhZuXIVu5wwaaYnQ7XmjiHxausUfzKikwzfZTt0ozrDLnZSW6BZ4raumKM
btGV3FzaLo1HaqHSvNRYSnkPFe5TFMPkIlp06EHixNnOOienl3ooqYir5ashVHuN
VVwGupMUXXoMhl5Ik8nqc4IjvoUEj4xsCrGWqg/r/wVaj9FvJ5tO9WskjdwFIgTR
0Vm6eXl44yuTH0b5+BRqw+oa1Z+DPFh1Ad6bkS/yGdlmv3gGX0QGL4L7tt4AHAdA
y7QaMRtasaz0eMdcuT1QODTXFRhdZKrAAmlNdfViBsHmDs9F1YpXSFjQPDVklr4o
1/8lg+DcjodGoNC2+z2dWq9BulGt5Gk7Tg55cVRNJTGHObtKvTzLyVRqmoWc8BzP
JS7A9XaGXh/pPUcfU6uYGILa85yeSTGqFIAVlOKSjFAYiMnuQ/T7fv6cu+mzPLUE
sw9QRpcgk94TLZaB6Awg5ECGenWx93jzTuNffHmaOI3WPbR/+heHdLa+lFchwbQH
wxjbqCqvv2M23de/Pw/6SFvplj1th3yyBHX0SnfvAX1L9uVWlG2aLZmiRiCookp/
U4aYhNfMw9BUbRYqm9TPTSvcvxzScg56xe09Wc7fLsoYwUi1nhJSP5JRIp4BMB+n
bn79ytGsdMv2FcZcg60ylrqmeKOaTIdqyTHEbm2Po/0sRC+wNfXVEIo6TSHcTbdv
TVZov7ni/QJMR4eSaJ+HIKoJjIe3ITPV++W3AkE5zg/gyeoXuHN2CaDkHIoWMx3o
am/mIOLgZLcMkrsEg9Mqq59nQlFszOfhGhpi6WSkPVbvmwtlMTr7gGRNWuVweR9g
oMM5T6cAIjwuHEVbS5Uo6BImrD5OHefyxd18NqVPtK7OIvuDP7LvNHHCI71ZMdEp
+tgUVf0r+hTeMaKVkb0yIm/tkQ+ahyvxqbP0XjjkCDlHbLnouOXgXBblNodQEUx+
XduSnsczTJZ07cbMVXwbUo6CyEyL7rkKJyqTdL1jIjWBcmPqh44geirk6KFnCV9o
XRsPi9mwpWnqQsasvJG/GtaTSYCvof1TMHY5q9DPsRznfNu+Q2cg9QfK3INugL80
GAaWgrQ23dUyIIbGm+2QXImP9EmJvqQSVh9NBbLco/lD/fXYeHumK8VrM1xvhKcj
epwokI0qy915iA7JqbBwKI2bUc1OUFSiIE3WiowuO+tVAhAdrd/z43XFXl86sb32
fGS/rEUtG3rtk6fP9NofIKl5YVaQxj9MuByXrgTR4mLmhMRry0Po5/0y3HBaYNzD
9uLjIMUFKndrxIplIST/ppyio7MCu+oFqYMj0OZyW+flZ8CymKQpvpOAT9Zypt22
l9ch5YaHp/oM8LWbqOmKn9nIP4WR4KcgIH3o0WnnwP75rj88tv4CiZV4lIYIYeiH
gfRbe3jgCpbMsMsPV8pfoonlmTkoFpmies+VbB9lAG9+byFOEjbOZJri9V693A91
LaPpv8cV1IHfrQkPP3FLuqdNBd91B2DfcGmA6mYi2N0YnW+46VMQdZp2rUWYc2w6
C39GhnkcA/bfDNxq9VHb7JICvuFPtKmfJop8r/h9JXsl4tM4y2/s807Boe3fJas0
I6lIURf3ZGiONhQn+abBFn3AT1MTproYYrWRhBmxigLEk+KYIyvyGAgLr5W6n5ir
S44zM9bgbf4jWN7+H4o3M1HFKq6W/bJj42JBFjjU1lBfnEDGWiiQ51i7d+sCE/9v
rlsEiljiamK6Q4j4q1KtTfW5vAvt/1P9eUXSERoeGsFnntAs4eCpnbEL2TvS+GEJ
KuuG6zYpOn+wgqyMUF+cnqLLEFFcoWIUNOoXiJ+P1+ysYx6GapxpwaJ7wUGK0FZW
p0fGB9K1HwQ0P2XO64dY98vEvNVUkkMWC5RgQVymM80NAOIsz+3et8EBd+WhtlQL
GOAK2tT13fPOggOmbux01mqhaz4KuzBUMfnLs/DjMjC8zazr2jjhaosMW9yhyT3q
aLZ1rIgX+4hZDNcfoYOghrFEEfXHad0wXwKdrvebCf0hLq3uvuEWf0nY3ObdXGo2
ZUf92C/j/aqIt3ikzGb+YOEKK6Ob6On4bOQUEqZhTJy/a0R823VSOCnhoWXySIZj
hOPmEMHBpfYQY8wsaBad0AUIt1ZDV/f30yz0u5dDRksVBJzwiw2HAbXeTbo9c1Lx
jhl83cDiobc3HvOrKkXw7iAqgj+QkccS9m8RsWZ9seLFwLLUzauA2zm9Yb4hZbcS
qj8owc0iC99b+qzc2c0pg1T8xmUCqErfv52s/+hmiCJeDGKYhRVtyUW5a100Ge2B
nYZbgdscQnRR78GVVZaHSJ5xHlW+VMpbkiJ9fYgRVbLBWbjColLNCWzr2uS4zun8
SD0fVWaGzHxWT+37xlQaOCISrSxFyQfPb9TRGT8XvVxPNm/Ym8Ip5oxKHZdc1QVS
6M+aTkjzZXrh3MZ34HCxm8i2lgnQftxssQOJ6pG5Yzns0Q7uOveFZTD4cy6krSnp
fWJZ7g4cVCBPH6ucUBALnX0a01Vl3s247zYicZdscPzt3FskT8pSPA9SV1fha1X2
gx8SjeO2C8A5cpbdXya69YwdpmuYXPTvEXzRLrocArEY1NkxNZfAbWdRHVz7+Hmd
mTfrIvEq8eZ4FOl6RqqsUThEFgRdgEfAkrIS8TFKfStUfaqHGA09pIsKiPKt9XsQ
/8KMIDiJyT7rTOk2qjwEqw+EodUFJbDHs2z7D4zRps0Vt943htBtsCvh1WsaqGY4
wUYBVB/K0Ueek9LoV+6wlVfyuhMRwxKiFsGVyKuyfimE6hB2uHKsn1HblFtskTAL
/RjSDWNnfygL7Bdv++lY7eL+/BE5SckYdzsWM6UR/J2REO5D20PMSAOPNdqMsAdy
b6yu7ZxUH4HKq+fL+NNf1Q3cg9le32ksfakEy+1Qv7L/YHruLudgRLWWY3NONTVo
WWemZoT13fHcgwEa3lKvJc4cCdOIomNnRcKQxg6NcW0ykqCcyOgePvqGP4M30zcT
Zo3eEfMimsdmacEKs7RtwJmnI13OGVLp/LjFsUPF8HA1OZB7yaSeKUjc0MMO8q8Q
Pcrc3cRqLmxpSM3fK2JZ0MwM8ap/gBEhenhsO1e8ofCSeyORqE77CzL2ZBrerFqa
eRGN9hilgo0njpgP20aBgRFXdBdIq38d5230U9NAyyxI+QUGNEdJLeJfH95s8lx4
Ewps3tb56wubnsCdppD7A7fMYUHzQs9QpRRQEwTfTpEfrFTUeFxXTN8l3QHDTDG6
kNoVfSkyoARuWXsm1fM3qJWISJgDlpvMrYmj/f8SIx/yehRPEp5+7+HiqS+cfqbI
WXmymZUI/gN2apRHmSm9VWM/4KWK1wCjwPFSmC9KA7F5PCn1F6/M0PKBzk90lPCy
OSEPyThOm5Bo6tmHHnn7sjqACjM0eIPV+F0jGogfRU3XuyJ5DeITEC1psPfd+Yb1
d1H4MfiflRPTMZmkoQJ/gAbu985xb+6hJOq8aAkrl35XD3kU4LZrnRkdXKT1oN5H
jEPEPOl0XZNHQ7s5MyTB7xJMZM4SxMypgT6fnEg+rNX59vDtPV5Sot5+7jNNHaaM
ogbhL9UZWVR2ozu1wv6Nd8iHkiMoNMoO/alqOusRW4fmAKzgH/Qj01tsAo6oewoT
6W66BFGzNXgdgU8sip8MxHLcdM4uWPt8Q9o3cpEPKlMotN/XfQni2MoJpBXZ4Lhj
tzm7rXi3EMpY2HdubcxWqHf72RYJW1tyhRIeJt90muqzjm7Qfki8FaqMdA8fr7MQ
3SdGjm+YRhw2HO17C0F5V7h2CVlFwUn8DtPi/eDjQmguyGUweFpS9iZvqDkdd6SU
F4gmR4mrVuqcqBGpJaQhcMluowJtu5Khyfb2xcx0QxrJqc1BSNwhFpELz5Gp6BiD
KIvf88BQuWIyuRI1JBlExOBXDfa7nvfNaFFAi1KR9mR+Vn2Vu0rxg+rLaUqTq5sw
e42MSERW90dCrDWvbMsYLUufoD2ZZnG1IFMBs66BTylTVJcVHogtJV6z5+wzwlS1
WVFY79GF6XSeeH6ReKUm8439lPVCYoPk9OXRECLYpr25sUYhGWKdtysnhiDUlOnN
JwSLPPgn9oocoKOJIZXH1owuWtIbSgndDFZsWMQq7NDL8YNqeJvHCr+awqOYHUr8
rmFBkOlHDx0nIX8CBJ+iEhGyuoLovuX4vCRzgQ3dvbQTk2E66oYngpcqVwjkelGD
QucrAYvnCa35rU8wnbXFUQA7KWGvZs52AllYMk34z6l+Xg6Y6KjTJPBcE0shIZPu
19J0wdGLk+GuHWNtAm7KeM2JOFPcbJSpaO6kvHzmJ4G31ML4aGgz+mHVZfvUek7k
6bC5/AG6+5c1ztkMNWbVkdSYsVwy4zbmPwVlZGndqFgrN+G0wupncU8jF+H2a981
R3SGP7P/W5g6cN/09XdZJcYLVhs6GqIx13j2UTPsFGgvPF1zIeXMyHyuAJ7UWsem
LFZv67ns+6VEX2/kvLloAjQy1IIIE89LbOgD2SpIVCRRfkhT/LvGOh9H3tOxBm50
hGYyHbqoBHDJcZLoL3kXe735AuXlgUcMxCOP497pJ92DLgRHhpkQdr6iaTzDpSg2
3o1EhBM9kyLcjLFTPMvfigoJlDUXBSvadRkKtjWYsXRm+GW33uHaBVzFqeE+2EOr
ZwWIulpVG6khnJlgF5HwDib2pbpCWZ6I/qzn93VHqilRnzhGbMx4ri1VM7yUTcAK
tI6RX6TdjBeICmwspXg5tQMhNs3G+GLV9floUHq/MCvaEXj2hM67Zz1Mq6a43xA5
++A4Q99Yl1My8AUdzfGJe2eSLgGSKbI68pK1W75pTD5dB3BP74xMvufhGk/r7u0u
8Ezv0/DYVdB5kuBFWxW1KGvnbILzpNSDGFYZdFEvciC0sZHBEJfwFm9mN6U53Nuw
Y/9XcFjHXYrHIkfqvuI0Mz9qkIf7pRt5ma3vxVnawaTXfLmWjMHtElipqBbUzGdt
WDcfJuRpXe9vos2uUIho8iAoGNSr4AvMCL0jmwN7b7M49Ry4aP3ZSdjlKePTMhj2
2RvorNHu3fp/fCLOp/lHKelr+GbXE7HuCIASAO9OHoG8Sxh+8ATUrcUe9Ek17Ny2
TSqQaCZ6iE+cRefAo1RHvzZkbXyihFFhLcWBMoiPFAsxnw/tYtaTtWsQEA6L+RzC
x+DRSemiPtn+1wxSxSa5tkM5T5Nn1DvQFthjPOwYA32tJdkgRgPvoVumuVtoRLqL
txO1DMA1I2YDE3RF0LvQCQB8luRou3nkm7uU6f0CRXh3YRkamfrdVYYe97D4y2Hr
tejWlBMvM/80npC1xyc2c79uYbdi681DnrZz4I/CGvPvv/Tmjt9CdmcODu3pqJ8i
bhmdTa9kgZrUGJbQ0RNtVjDR37UvInvqINHte0jIeaipwHgFTPAuJlzEoYdhHhXu
kZJ5kUAvoVQ8yr9g654CD4BRBScdSIheqzFYY/FYobXyP0Db9eNpiq69K27vH+xi
afQ3sKgJvN6dNVVVME9m1pD+c6Cuhza4046rz2YKq2CsdQ4PBvcQKM8d9IkP2uLk
jo1et9FgKJ1huj344CnN7MBGUgUyFHzHjPg9UPZLFSa+sySHzkJA2oBwDRnQeRhp
Je8bu23YiXUw2Ed9owBjbBFTUBSMrFMMqa/NJrGJs6t2Esug4OYETDa4eYQWrElZ
kUtiaXE6eM+M4HDFmb7mbBrKY5q+xN9UFrd+mo1K4LWk2nnfstvXWDjbtJNZLnK1
BWnVwHRXi4uyLbj7ld3UWs1dD1Wa1FkcH/TFVbMsqppMrUo9zG81ecMimlO5K8qN
3JeoRaSC40lp9NNJGDY4Fb6zQsM8V2k55kTZWode08fkjZs5RP9SxBVCCybqX5Tc
bnlHfB4eUSdl33A47uAHmpnB7TOLrVuMepz5p4ZLb41evMXoEUCZcBCK2e7GUzi2
dzBpBM51TTVrqTPTumBCD6Qy5EUN/JbdB88stZbmmiIO2UKhlzCkF/huPFG1adZV
2gaXcRx+mBszSe6uW30tRafaO89WzUx2FNx6tELygeeOih4LHjQH9VDrRBNUbqaB
8xYxl5XCdGKVsQCBieCQMIqPfLdRBFbSPbg346rPSCDOXEITkgYP8XTh2pU6sfA3
cSlY4u9+I0G1irDz+XJRbmUNJr2fHNVBgX2MmGKK3ztAY5mZwzo+fnjpb4oapTPJ
lS8DEM9+bTkZy3RBhGM4PVjN/HJ6BokgRbj3LernzeWwe5kB1Cyiz0ryZdFDMemH
Bid8g7XU3Dc2tUFrpug53nyvQxNmKzB7BHv5P1yZzOCadUT4i25FpsG9R3P5+DiH
vPblivc4G+VMYydw3zWyVgmGugXl6qTvS9E3pvCeY5SINDENhzaSWnrcQg92gxmM
Hebjo7/9sTOY5TQRtDKzN6mVmuvFTXyc7uoiCYEIk2LZ7rqhwORKR1a5FdWO2J/p
UXAGk69Y66pLY8DWGb5Fm2Ym81rXX59ofcVJk0q2lK1Cw3Ni8hU0ULkxsqTBk/pX
Buy4oJvEFQC/znuiCeNgdvp5unayCr8xwV3k/Np7JUwRhib6/hPn8LOJlq5B90rL
rKqviYYTT5B0TA/erS0RmFdDal/g7Fltqs3HjbS+1KgofCVeLwb7HdFjD4xcGnH5
8yzQB4qCfl/n6liMjhnugeGYtg8eBzZMvv60P/WbSrOi6NRavpmSxdvMZgm6X+2b
hf2RHBDtI04MpyPfS1upOOVcg4GkGPJNM9cnHcKXBaTgfKwYcGpaCCLoVSvURhkv
7DQHWi05Y4lcOsWAy1he3rMRHGUb4XC9tHL3pBC7g8Wqi1wdIO8WSP/KNFO6uedX
VcyE0HxfmYxeCx7VlQOgdt8+ebH6zBl8v+nLjvjttnvtgAFd1QpJB6eO9dpADYR8
4Xgq8xC1/R4SwbUn/9GizStD/uita4v3P+OMz+RSYJbe4agYNfpc4iv/fsVj6wGA
ZI50JAKoMU6J7jHfV86BPqX2GowGBpYUp4d9v/0yZ6fj4BDa91y+Rt16Chug8FBL
5uNJKlUzfi6Bj91Av6qjqOa1N/qrrDLaLWKg4IQaeAp2JatEeSOQHkgse/eWov8y
wwgE9bxQKNsw00p0aDpvOSjz3JHAT5EukIW/oYC9z4PIGdn1Zy2WZe+gNiLjQ6tA
c3k2qxRMBNWjHqTl/VHcIPVPenW1TnVbobNSDAAdn/sgUsQoOy0yWF/btI2OWG1O
je/Ewb35EwS4QkBFZurW4uui4erF548xlHQGOHe1HJPDcCstR7GC1OIyKyiBCUgp
Kyjeaz0EBOdX3J7WJf/JAn9pOEhRCGCu9jRPileaBCHtDQ9l1TSch4mzADlCC2nI
pWBfQwzI8mopDFyf98ADUVIk40Dn4MnF5o7vRyeyUT+NpCpuRVH8fMemUegmAvr5
BMxVcovJgAfzwoUbheipWAOPj42lN5ECOAwLkHsQBKoPzWWmHQ950nFUF7zyLWbo
acb5ZqN+2WXDkQ1/q8fOd30lIbtEE2VTA6DsoRz1eF9mvL2KrpMIVsW/sIYmx9w7
fAmuQ9CNrwWd4ghvHdhk8xmYSoj7IxgANHVmPpviIIyAE+E7r8wXRZVNBDmyUZyu
oLJuuk+5gddl+0goEPmqofhRi+5Ld0LoyLt60OWPZEWAP5K03kUDoilp25QJV4FO
CzrNQWvfWP7IMi7aMFDxkVXxWMomTSOXJeGF0NhdypBFuQKNOZ70lgP3Z+1sT7ca
LGpkHRs6qypwO6wZi2558JNNMR56tZH//6y4LhJlztcpmu8bv8aqCBpYmOiM2oSP
CWzRg8DowgtodChB+rhHsx86owmboz0EU142kBYi5/rpLWbpdoF/kKvvT+Bklb6v
5G/rc3rBnFECRkplXIecdUgu4HhTHWOuydEfXuF7QfOFMYsDAf0Xdr6AMwLdWXZs
ENcCDppb83AzOaOBxw12Mt51Y/7DqFM721nwPWcZIipeZ7lLWMPIArJDHb1lELkO
D8cE13Y+o7+eXIxTrw0R/PLvih89IPMeWdKVi6V9SVlxycoleyj+w8aU8buf0Oke
1qQ0oLRS8ZP7euKzalTZhP9ab3cdl7/ikevtTWV3bXaLtBpsl9fUYrU/q+WTCGwH
wVlFfMePF35YYGUsXkahKzElbwVdzWRyxV4XbYf/akeOERKFHTEzxjScGwVL4jHT
Db1Oqz81/P435eLMpEsqiuxRPRK7++wdswG2XD6Q+1R0qoimTZ7TjgBjih/K7leL
qu1hsjoQVY4+kka/lSdfosVq7E0PBOVj+NnOuiGd4rWQfQ+3F+A6gfXI1hoJ+lVB
YkXw86QLnX+guo2BnuIY4nWEvibEpjY/0l2eZoePhSQsvF/VaySY5bbkiPX5d5Pa
+TX0caMZMnhA7Euxt98AOoHq/ZPIi7gaaeacQ1TfF+jsYMm9KcLq3gLvvTZ2cmRH
5JZC1LO77LARZy+1uzge2jTfbMlVPaYvMTK0T1Su4f7vEX3K2F+zYXJQBemdI1fY
U3Gwcvd0TGDhmLZY7GDq2V9I9UfGpuwljJ1zFEWd3TtgpjOyU6YqeMGbSBGbO0fF
9b6a3zmhLBLiJTjzOMxu26fgYqQNsv8b7Uxbei8kp5D5kz/7CifsMbD6twffmOsE
pyJaUNVLciDmodNZz/52CZgwyWy6lAky5ETlJjRjFe1v4bD3WkC/Qnc704XtxfDz
b8w/w3DQ02TwmB0E5K/36a/P7Ki2AKFkCQOvuJqRVZksnopZ0KA1YGS7FNVsdBZX
WgR0Sc0/mjgZ52W5SzthYFPk9qQVVssNcEeNSMRVwkm3C1eG7KHIX7drORkIb1oj
doQghWtM2hgtV93hnWAD6TiAbt/owPJrcg6PWbU2w7+Ut6ti50NcKjhtbhOxdXlQ
sXgleSJsQjW5fLPwd+UuAmcCkFms/vsW1sUZOEFS9IwqmoD/WM6rWousuzw6wEOr
vEopLlCG6afgLzrTUwGwGmiII1VcHAUM1dsxDC3G+F8oD5aO02Sxo5vFjcXZJ08a
4a6ZaMi2ZIg0ti675kRVPC3m0IBgNr+YtOEF8QEhXBNGUX8biMUEJfzbz7siErYF
qfRQtUNPQilLvNCZqVplo9wbmGQnRZbRQ6Za+R/Jn/CBxSQ23piAPLXtzygKjrcB
BZxxy+OkbhuNVvwFy3Mt4BdoH4CixHOkuXBR9/uEneNrS5RtZmfJNX+otGVP+54s
aE68zK1pIOmEeObg5HYOM2r2ahgT9pqNRfaBxZs78qw88hGwuqt7NAPgN/UV2kmJ
Ty22p1xVT8MlsxC6u+9ZHRKlVmpAWCTGl7EuVCBgYOaYAwJJ54SdqWhAkQ6+jb4p
g5fW+GauO6TyAuscvbUbGCOavYOLENewI9ZK8u0UlyG2FpyPnXVfaLJ2bDmuH4sZ
ZbxPwjmwehZhUaYHaQMYoeJPv1qhJwLJycw4NCFO4gPMphZfdgaay5PjScu1ju5p
gZ/7bUn4zvWdj7kBMze4oXRqpTZflxIIrVwEPeG4VHH4a0U67vYgpAuyMedAElT/
grsFQDtJBTWjT5kei5AMrAjE3uOP2KYT4BP4csI/X2IufrN0Fz/powE4FpDljlbt
4dnrZARTXKiS1JxJCNcEkEkgShw2k+e+vfS9tXr00i6inL0PVr1GwnkuvFQqIXrD
B1LampuH/8TIGsrP72a+GtEgfMUxyIAU5KeGI5v0tJyDf5e771Ode1WC7FXFEHhk
L7WyVkzJzu22s/oiPsU1fZxZDgqqmmVUd0/gitwHsF+8wlhVM/7qMwXE5oS9D2og
arxSR/6ZQ97sKbx+dKfdIE+96ZeWaCy6t9ea0VoFatsA/6TzToyb24lFwb4VI6iI
5xzFoUiz7SnDyetOqAyUjU5l/kCE7NQDZ5AqkKNQmFQ9V2WaqB9UyW8FdAUNrq0J
CRgHxjTawv40NCznkDCt5xqlO/wSGi2Z58y8MA3FvVmcoIHEAY7jnjKviPZjBfO5
cbDrLx0NO68ifMi2XoHOW77i7VCdav3eEiqF2O/soMZyeIeGUqkDguAkIIRZ1i8p
V1ASHPW6gQsk7NVusjDNpW9ekUdbBlkqVYfFp2HJXBAuYUc+E1KGK7VOZ85DcFY/
Yz90nAbv08gqLJ4el1AfPR6MaapkPIy0MuXRKZH84zsMF0h9LtrE2pB6Orp64+RJ
bbSbmEOTR9e/1VAYG8mwI5ae+eqMUgF19pTgi9TNTJ+N5hHMarN1KLLOC+G9Gnns
9ilqE35tNWDddzAqRIJFG5d0GoHYa0ahFufa7m6n21+8zrock/LWmNFV0lXsxsfD
dHLTjyLf8SaWSB0SSTuYoBCyMuvjq9n9qOp46FRFzURCrI56lPZpm+2GLlpMjquX
X0R0N7XimsFEJ2yW1rVyWNBAvo26KylIm6IwRzHaQgFKktEwnYwjjh+YRgMprRNu
//aJeEs1Vxrqqq9yawkmM2iDRdQesgAdcYDTZuCkfQ2C6ye9NrvBLKPeaXFF8vLn
RoRo/pb1mwji2gkfVX/HjbsvjKxWFE0g3bltTmNUHtIqqdF2t86iLYJGLmn4H3UP
YNj7/CgZK5F7BDT72qxHVJxvDAt4InEkUolsr9jeT3HI4/lpPMNecrZRdODTdOfP
/+UOdhIulVAW9rEnlJRpDVRHHa5ch5nY1+x5oDB/UwYtYfmpy4vizpRcWRXVwQ8m
ngduKzqs/XTpNIJwuwnnNTU+uY+hDagPZOTO2gjLm/Z8gHoYDz73Mrcn65SxZxHE
GsYeIk0V6mu87uPgmxe4QR1sOZu3AlC3XwKUwlD5zFLEORYn6OWOR96KjPO94vO4
+syiV0DV4gyZ+GKAzAj+M2+xGvsuHbY23pUMxboMgPWG2rFdEwKjGzd3eLUiZIky
WLJamUP2VWTZryBjVQyQFlMusPjKKCsZ0IuT8SLW1iiWEKEGbJvmxkdwG9QWo3E6
qqtMQnGB28NEWgVtJnGw397VtrPKuEdeqY7JxlFS0K9sbuN6wp/BBgS/quX67E/y
RjOFSXqPQuP7UWmqcdzlY4iF9Vs1QtxDbNUf7ZFthpjer3IJlDpTmQTVUX4cpEnk
iXZ8oI86cobQrUdv/NiJEzZMSel+CmDfZEBbvwy3jiwuVoJIobwVLzeFBOsZnSmV
pLkQG9zFM7KKjcd0YCbS8mG+CoB+YHJ/ueSUjwEvfwUMBL5U+UiIArMc7RXB2D2g
/AVq5gYcpQRC02gsTmu/I2UwfZ71TrhB1PXP9qjrhgpR26K6w/4AWevBsJb9/gE7
5XWongtmCyT7aR3el3OH72UHf0SNn9uDnQnsDAdESFj89oM+F0ACzd5cYgxOAAB0
fy5/A3drSaVP6eF3gLdD/7DAseCIdkT4M1UYcOBZVr3w0emI9C6oelUiDgFBd3n4
ZypZURtH9PqEjITsYtNuzim5YWuGfAzbVc5fes1yq29awdyLkNXshu9HDPOeAiMA
VVNlAksBAAiraQ/TaYArLuhwSrQQWbTgY3onxn0+BH/Hxz1mGu33dlf1flEfmqGU
cblSCZGQOdvJEIBnFkH+lC9xE1r/FUpwFwLvmEKMkO3hwUPSfVnPDlpHrGoS3uHV
GY9DgtOW7Jp3YM7QomSUrDjUMu7hLjxg5lm59nEFqTvr88p4QfmkwIf2QbgjWvqW
KRz3NJkYnivPFZ/DLJAuhNGMbRWoedJYzcXvf9BTQmm7cxtViu9SLjKAI53nwbAF
Y9Vip+rDuchPFldDyW4UyyXbhubv3TOqkZZ6vaFtZzvrNtrBOBZYiudKXiqBluJv
Sm8DKmNYopmVLCQDoFCfEvVnwVldCcfAHvOTLkNw8ki/MZWrmdGl0J/Aqzt8TkX7
VhdTdsDTaN9X43J+GAnuORTjJwAunrewxUKqhPs+YCPQYDkljaOEaSWC6Nb8Dzpi
+P4nirZ44M187BuNw983rE8ficTKlcN5R9R9ZGPJuWJEhs9BrLm90C5lAlexZVLk
tntHZIQD8PPVR6LMONw656bhcJRB+q6mMVPniw8S6rg623m9pO4glBjxV1WjIqzA
EqlKt4RMdAc29ELnSOzgNRvtsDpGSOM+t2ItCi6kva7X6ha9jk3RmVqgP0bB5Z9l
HvW3xsvUJ8tlvvaCCrOFuAXo+Zax/CsDGakK8/UTALjGJXY2ztmJDNrDay814ifg
EpOODZ9wFrB0RAokjYv9muTSJxC+ztM3lk3EXKsN+ykE5ghlgHecbNE0/jgd6W87
L61a3iXI8dci3vsxDsKEEgg/g08Ysb55KKEzB+BtRDD4Rx3uYFgivIh3sPWaAcZh
c7lMdnobnMahOC82Vo5nkExv4YsdimO96jOM4ROmKZlzLp1DVme0EYCxhzwEFbeo
/t8EB2EdIIssfp4M4Ck9uO1lD3BljMCTDmAofJDPKoa4vaoaeZnanVVAuebb5ww4
6rlmm6CahMRlAY9RvPNBquzamoyx54/p+ZrGm1MlEAS/MIlrYWeNfyeESOFMVxhX
pRlV3kzIEv2gEvQLGVv+aNDMDnTV0l0JD6oFxilpz93lUm5sQpahXOui9pzpM93H
mU8jUCwLJsrjEpAkSeKQ1WThf8WwX5N6arT9rz4LojbdcKqieesV46aj/435JVFw
ESHg2+JnxmbQD3q2CGSkPhWtGnwlDgJEKgXnzI5y4rh97wCUOuLyUEHcH8ihiSaU
neJ/CxctWn4bIjz/pvWW6cgnOJisTblAcKDMbO+6r3+fpEfkfYekdIh2xY8y4dev
B738at4ALohYHO4jihBtBkGyvp9Hd/zIiKLZWPH6dbCEEY/yYMXi1UO83JBCVj5c
y7jjDoreo4TWv0SIIM7apuyRTdVw8z/gBWI8/UREDjdIkp7U75iGIAVqi0DXXJmd
LG2Eb7qcrzF+256LHpUytdCSzwKOUUheFPCNSYaKA9odxltkkE9Z+y+isBA7g+V1
TMpEff6cDO087LZCt7uRHqWclYX2/WOqvjk1TmtlzRNu7Rx1t3GALu7zPJsHLzY7
+4FfY28QD4eJYyRlLlKEzLYIxGgWVd7lrprF/oNj+vRXHm3hCT5o68Z1W8helaNr
hHMNode5yYByRJUEGdSdnpvK6Hu9IG2Tzth8TjQrnJhENJGISD3JYivl4p6Q6H96
cX9S8gz6OyBacq+lYHqSUFHvUMKs92J9m5HlFzsZtgqDC5VbpsZsp9Ahq/USL7WP
1pewbV8Lbnpo7q4s9Fi8rpMv7EBHdCC6r6OTLgAuBN3PgHRvPQw2ZGQ3HtFzHsR6
4bhjw63bh88XnNNnhaa/fUrpSlq6NbJFXCWDNCrwljj44XhM6UCHubRrkQSUsigX
Vzh2JwfyToikTIJ/3+2klitJxGn/LAcg1mE0IsZ1Gxk2AZmce+ofEIvDM8UpXW06
wTXbKFfeV3OafvVZ4xFDTFgdD1uMB8UyZ0PSYCo/FKHWH9jCfWHNPZaB/6I94viT
MYcuUS9khE030cMnnjgQG3NjV82/jyi7+3MmaS/EOUWeeiy9Fow+k3P43+jodKXY
Ii7eQ7Mi3DDf2gNCDYdQHkhF5pHpPLJqKcjsvlHqEe/mWwXuHE6wlhW7HG7d7hJw
HdtsgHkQvDtGnhddAwBsaIiWVCyZC/PTnuA7oB0IQUPFZF8xraqT5untLC22yjwI
1Y8TMDdXwT6oPLLDfa7WKtuOPgmsa6XQUR/RoZRN4QLmRo/321o/YUzfrEq6BrX0
hMTACEEXE0+j2479yc2bfcDmYIW34pVYAXYO0deqSbj+3WGt1e4SmlxG2N4SAs48
jtVhWMfsIxHBBSCspt4jZWxf0WbeNbJZLZrVmfYsQI4ilWFi/QD1uc+xc8NP+XvI
NjZ+FIgaFcU5PcFt+0M0i1Eq+BOeQpKnyhR/sQ3Imsuwqc8GrvOn6XFRwDAbJKnc
q7EEM4bDG1wuQrmDZ32vSAGwZPXi6D50zAEz1xz4IGQLLZLGOmEUF/oQsEUmhQom
4f7qJ1+B4wpSUBwEfEUssVWVXjMrI9GCy37pB1lceS/KRmdYSQyurh9b+JxPQ4yq
YZsMHK+Dr2nt5fV8GDc5rujPR1FaC0TuQXj9a3Ca0qw5bqM/C/T6UTwnbCcjWp+C
iXXGf+auJMjybMHeGrCu8jLbXGb+tC43u17zICPQNMrRAXxkCM0zQdF44CS6E3zN
/RpQwFBuqUjLPB4TFTIi9cPjNDOYlGmmnvdedbYZvnIsL7vpY2/HGFKc+0N6eO/0
8bd6npBctlWMeAk0l0fRlTneok4iKk1iq83Iqkk3vePAAtIJVw4fG/raecSN57uE
3+tjoQ0tBBGleBP4hhtUS9qS+ek09wZIxNmDowKiyVw1mu3q+VFubI2MQ/5cXWJJ
c6j2IxeKXY1pMtVlYQU0F45X8IeiqlFi1LOPPJDOx/ZHpvFuKU0hO8oqPQkqAZjp
jXSQpzzuTUyEC12kNs2x0YkM8y8eZfO8x+r3+atycV6NmOgYtvRNyj402f1rMfPQ
a3MzsCTcIV0nNwN/lus85UZWLQE1RJ7Q3wo1PFbYxlxPHmMTphlY47SB51s2Kgyq
N3zVAq0C1dpovd4pnallH/b+EYStDwfnQgpHssRj6PXvMWKaTktGQ4gYCXo626F6
OpYTONjCfRPoxq8rNq3F3HXbpr/4DORW18y8ZNASPTyk0Tu+vJP8WcS6g+Hkr4OC
ehpUKwLCBt7D8UU4Xg9j+ntZEG9YoZHG+fOuF29bCFCIE4TCRu0V4ouzj61ZZY8T
rNuMtLPsE9zSzljkiXLjsEu1WbawlJkqclIOLxLAwn6X65I67+Uam7ALaENaWt5R
g4ZTM8sq0Dps8jmh7MMgPsLbOpBCJLb527jXVjSfllwlPiN3ZZ4EZrtZ253ZW2Sf
gHO46PqgwTHCvNvZs6K5SU4W3+zwDtzhLX7VoLuptBoNJEePuc2fHlQRfwnIxrTP
xDmfNJd/CqVP6OJSzRVatvoWJmR4c9AzkgjunSAoDUsQR9LE11rYiG/6RriySZP3
BMiEAB8LPLWOM79dlhGNm5ZBBdyHtpGCxfZ4DEWBrCCvTb6nCPliRSMPl2+EmAiF
taKPSvNIeCId2TQurd0Hvqu9EOtOeuCk1eAaHiowP0dqjs4rWMtcoHQ8JPt4e01b
zZRa1emp/yvJfXeSB3HMnF6+f1eVUN2SJvxsJ6X5I5xW+w5QehsuHb+CRRj6vm36
4q61f0hVncMqxgby64hI5jRrpNYh4u9mAJHeT7dw1pIEJcr41jtmxJbPRkcIyOS1
SFqwqk+BgQJdJLJHUA3oLKcdI20BcYft/JyevAqE9+x3ztT36tVeesFxNreCdmbq
h63o9c+Xetm2sIWB4BJadze+1AWNUnQc0B0qSYudrZizpZ3DOnFAsA80J4sUxoNH
XaV1U7tA3m200LfH903g6iWV+Z3MfAulWj7AQQSmGg7D5/W3NkBJAf/h6VT4Wl41
N+68XGnWTud6wT8xI5qKZxMrLJW0v/l13+r4nBenZw5F8XiWG5tS9FL25XalNeW4
7e2SjHS2IcXfXt9hny6LLVonO4jjzT7qFErgVP8+oZit3DZHsYvhhzShoYmvZPOd
exvCdUT05VAEVGdNb3+q9TSw4t5pITEgf3xGSmYAT0+AwHkBhkZuxIAcKmYw1ZYR
JOC15JAF0iHakrl1oOsirfj5zIUveAga6zEahhHMtyhhAUeNIGpBtsLG4k3qnLst
vy9frXU5R4pmHodixFzQmUjcA28Cxbeahip3ORaOUFAdEhie6Px8vBuQ3n5FViEG
iQ2mjY5eerLbMy8G6achIVFORNpnCAcuFFw1MW3yyMs2q/kKpvUn1wqmquUQ3JFK
foOtPrIFKWl1haGKueEJTEjUT0IXbesQoAmSrI8fmVE7PDky58yv5Typwke5/gca
bzWGoI1hsR+8LbiW76qkrCM4LPsXVYUHBj+y673iQGb5wIikuPIcOgqtazdoQ/nO
Z+SHBVaCk0MbjrxUznE0ZAo/Dieo6HuZSMExXQdADmDytPZQorPFe4C7c4/Aes0S
5TcQ3Qj0pBVrAabDsOj0voFpcTkBjI3KXR/eHRIpCezMe9zcXlS7scCECrJ6EH3p
9131qcFrBx8QOHq34fE5dum1Poynu3f5TLNXfgPKwxFSWhuyBcI9948OcDxBUsv4
Jx9bPxvZcuN4YgATe3vUu9pO021NP4LHgi2hlUfGM6NwTAgNrTFWJYwTt6pnF3ko
yxQq6ZNNF76hb4dSrJMjXHqtW2QYldKHvrPOTHeZErGhHRzT4VBc+MJMgC8qB4I9
/AannnAzwTJ1D0HQmNpYi9EP/uNpa+r/rk7Lue0lx5X8aNj2KHdSSntpNeX1/ZVr
AHwyUkYT7NV0mWo9dfUD1ubUnE85mgZCH7UglqAVlJngul6EhC7M2uLNi+YL2B6a
z1FPky+1zl++ic0Je94r6H8NFCPwLSOYkxr8EiMJHU5xQ2Hj+BUUg4ZqahtXvaZO
ru7uKqpB3KrFyvsopAHnTruQLOT+wEXnLH4y64xugBfZirdGFm8QMwjAx4/OL27/
8W9halSX4VYPo+wCw4WvkywxVH1vfXrvCR/0pZfMMXV1f+530gB9nOltKwyvit+p
ZN2FnsrnMBJMo0kJ0sCBnQlO/+EuF/wSPkSTn0GPlMEkz6JFu7RzpGMVExtKfIgk
461/d0JvTIaOoYu+8xn+02pQcdEhl2giTNv8EMknLR0YdxaWlILDQwV4XkY4rAaS
Ei95aGxirrWYm/69MKmuYiRo8E+KxOggMjDL3IzeauPZuXrplj5ld6ZrlHxWAiSM
oXTsc7wJjjI1EZjW8jcjxMv0JNYP9JqW/frmffL15y28dFnkzDk40WPr4ILrulBR
gCy2BUbAzCfuSEJyawYrlDqX1IsyynW0P6PTpFGPBWAn6bLUDUK8cbg1vJI7UBbg
frgZnWmT7ubL01kTKVW5CalVov02Rp4J2STA/EcDCnEmO4ABpG65+LusWujc6ugC
mzX9pMKRLrDJowTcav0HOLJ1I06vboKwquIrD7nu7RfjXhFTQ5p8yNIaFgE/NMsc
8QZYiYrVYBgCPBBVIRn4aVkDLL4H+Ol+3xBn4/5W9LeAZe6we+6//LqDALdsUyJu
BljfEhiR4dWVZ3BKpK9HqMYfKxJbjgLTzbZJfj+qtHpmgfiyOmlb6CMSOoGg/XOt
ferkm2fs6Er4oxKy3w/rWFJDh/dAjB+tMzKm9fq1RdFoNxe7naLNceoNUFhnLVnA
XNHJntUGyPtUl5pMHdnzjVv8hpML0McYIsZ3gFADs8Q=
`protect END_PROTECTED
