`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UBQ7JA0AR9r4U1tg5Cqrc6EpDjMr+iX0SHf6NIJVKxQ4X3ihUxW7lhwCai+HDwg7
tAc2dNOcrkOFtMGXjYj/eHmuJKiVAKxhQKd/GFnhfgPEpCY532P5zRjfWeXlFkYp
6GJNTnHZEF6LASHJMEk2uop9U0UNQZ/m2NBuBU6p1gSnpvxgM9utkrKDdhXEAoBT
amdgzFJjRZ+U8oPwFXbGOEp/f1t1xhy5LvO9mzLVBYbTrO0noX7SoYr/S+6lQCY8
+sBjlNOWYXjlz3hYt+LEfzuGbFrmH4kSyOHdCvTmaQusvzfvy+gToZoHkRUtUmVR
eq/BKgI0NWGAWS5QjetkdVaXDB4pGHt2SpR57GIIBwUa9ofXnlBKyObSJ5/xRGY4
zWie9GbgNBReQLUJ2QR3fz6TNYvi7Mir0XqEq2XgmXZTWlEZTdCoDEAeecoKPx0k
3jLYE7LI1+/wRMcs8r4ZV+qw46wVUN/4BnTcBgQ4mX/XtG4k25QaxUCEys9V17GY
h6NggP6B3sRaDXp2YxENowh0Bw4Oud1ZGRQlYc2XyGh5F5bz/3SZcyG2j0ZaejGx
TuRfemgHvKhTOb+KdxizVAu9EpLFkd6M0iZblWq1tbb6/JU8v01S/UOnyHRJ5PWR
mmz968DSgKnC1xqDAzjKZ4p9wmqX8vPVV56Isz3mNx4oYG9TgjzSY2CizlU6jnQ5
96WXCTOZLzo805A4o9JghI0rH8X7wWoKKJF5m7fkene11ewykFYGZ0CJt2rzdTkK
jNsY/UihEv0yFEVt6Yz/7iLncPSHIjI9fZgWz5Nj3B6a7xj1bC38MhDEst7xpe/a
4riRuEq7mylvZLk/1MHa1j0S9zATNf3ddGyPqsUWVNNksCrDEdUvzPBgBBZgMqar
vKEybbdSU4WIpxEiuFh0qDAq5Hs1SFx9dtwYgBi/KByEjv9qrCqvuyHmlLcIGt8c
wgVcj1P/oi/b65UZMH4xHD9FOJv9plhFDPthByxOAD4k8DV3MOZpoAUsull+BmuG
K6hv6svyR1hPLuCbzKn5aTUfiYEpxM7Icm0fffku4QAfcL/tJ0NMYywCznfpBxe6
4UOnIQQJpO6OICkRdj/ONqdpLVUWv3Lo8b5WVl8GeZ9nr/apLOgdfT3nZgDOn22G
llL9tceRxvv/XTPa8II1LvRO3EFKXDogrsFS4Ell8MN4ZEbNOtoEBDxMgSaNtWcC
7T22G+Z9csSxoVYL+BvPQARNQqEkUN9UfSeBvAv1usalZ22lO+aOugYCopehGDhR
oZT7wabf81Kk6SRIsPj2fKaEK5I8Y4iz66JSpL2fTDqaUkEQdaExuM9C9rReV7g/
2gTKeEXi+oArcVWC/7TAdNM1fhQyblXX+PxfsolQ5y1fMwxnmrgAHgMyCl5CJini
oTfTtxKXlT91skGi5CWz0Bmc9dSrTHK32unoItr6Lmism36pwploEwkHi2Oa/Thz
mUBdaeLRfCIUGHgLqpora8e5sKrG56JdCCWqEhW0Wk9HAw7MF72iymGs4PmnIscF
hdD6ZdYvRBaKBIHb8lFv+1uc79uZhkMTNVbD5KysUaBiACBE5LFNjSkR+NRuFGRR
U2TJlBx63W5L6jwij8cLzEiTU6ooLlM/J7PaxdAPiMVtP/CV9XXlIgikz07C1v7m
NRVswuG1R3wrKLNKV7M61HQwVyYjENv334eIBYa/xtnxVyVTe85tF7yFcGxn9mnB
oDKd3o+V5OXoHeKRV0T6v9pffLc57ZSLpNxFh/QN0FtHIaJ6yS3pDScg33w/Gbr1
84VQIl5pLqPAogOHxbI1u/Ls3VADkBrD7qUrjj/OMMyNcSDfod+2SwZnm4PhrSGi
mRNPRbyaLGTZpQPPZpYNbt/58COYXn5PPccKed3E7i0nmkKQI4c8Znvm+mIHAPhA
xoAES8ywRvXL+K5NMDRneLpkhi6dcVISPokOLfJ97TAaDWo+CwAV8rObxxCO8btS
Wq3FllSVA01ULLIaAknFaZbCPJD+f5V/fETXrRqGJ6VerkIhA5O29JyK+KCIeDKr
ZprSeuIXSf1Em09NOCoueWgsFVB+twHMBD74Yc+JNQE7/977hgPI7uM1qJSVipid
1FjwphpNyssuM9zm2tpNqDP8d8+JLfvsrYWTkfMRe2qffMitP8X+/CpDscL0lF9s
EE7xzgWXFsHG/7OHwRE3g6twmorNCLwfXO4cGLQcrqjtyJmvLZ+Ths4XJQQ1H1HL
AmAWLRpFZ/bC3F60hBUjta8Saubw4Bmke2dhVMrxkkmHGGvXNPEkb+dhaRfOSEDc
RSnMMibLhtNcrljd5M8K9xI/QKow4fMSZlCUpB/fWnJTwRPGQmKHnvvp36Tkk+M5
+1tHisDNUr4o5fe31GUMtcg01OINR0qjZOB3Ok66Zrg/67mnMnpxLrJkpxN3LBLj
w+Jfr635vL27jFg5C2rtla2CDgDpYuEmwrhdJoBfEMK9E6vACnBbuPhm1gk5C+Aa
AqZLFYfdwO2gdk6IRWzgFVyeqh9+qhhYy1ZWZJrmlULZNNlTJF4BXxTeuquFm/EC
CAn6LsqmAClP+j60ZgmMAov6qCOQSWo1ZCJ/VDx4xFhxtT48085dkpf40+l8eYXR
zf6GVd9KX2quxi0edFhj7bB5GRJ3hNemtomFL0xif5QRPw2cV+LdF6P7mdCx0hT8
wzum8ZrRzJEBNmcY8dBjUerl1Q2CIvXvvmVsgsxNQua2Xl1G07TK7cjC+hy01Meo
O+h+jt/+GjOrPDucaXoir1Ywc6OaDOaTyHB6MJBmMZTVQa/UpjdIjQAB6dcID48x
gnGendRi+pPQhb0+6mW5wXu2jDDGc0AAj50yQL4svifdmlGhc7Dm4ZaJ0DOGh7Pq
bhlNmyKB+bDlZdPR1OEm5mp5iYENtzo89wcOXJVx1YBwHTXtrYkfSS09KAan16J5
Iojm76zqxnGOoTmQ+gPG5gGAu2qW6cUSbYMyBtPHL+IJk+L8kjJ/n0HKdaNF6bSh
j3/5bFf8USnKYRpwJq9pVCJAU0EV35+GOQHpa07QY375wXpZwiRo+3rWcHLW5Pv8
koKDoc8EpTpCE38LuMl5Wrf+vP/oSMIUkBh+JHUnlK2ERuMhLY+OZIj3XJGtE4o+
OAV1eax8VdneZBT2w4ag+qirrL/GeP4Os9GHUIdJTbmyOuoaVCPVAMY4XSY9Rksi
y/6aqQMD/AE+mZI2GivFF7MY7zd++tczJrxxuBp9Rez9YLNIgh8TnlpUT+S4FktM
ZjQr6KUTkovxTmkHnbPDt4Hi/dWZmYrTYJr/lIz86joOEFiJU6ZM2bTQR4txJUHg
ce9yCxPCTrapUq6Ck4b/5VhkBxhX/bSEuZOkl7UnypKG8SwWSrz8N3BE7YY3YMYw
ZA5+WXcZZZSRJdeS8AfcaVF69vuzHrxX6tvvZUeAEQb7WPvXFB0LEndRGaydAO1i
Ong7R9X7ff1/7IrLtOav2t4FxwXLHd8+pqfVcwN5DXzwTWmIojAHkOxb4pkLO0PP
jt064rHu/xaxO3kvMm07DG8noYBci2gikuSergW7e2x1pNdeR/8LtZ2XjcOfbGfA
KjGiaem1esvVz7Ctx5g1ByexisvkYbxlw8ZdVkNHv9CsptHERpsMRhv630hDStXt
pGqrELElLsQW8Z0ZrnkM6iqquW4pHoSzSQvJHboAAxICKvUJviAUtRZynPHUXwNE
tUpkWKSMsoezTglItzM0kX7G7/R1jsdi7ibdh0Enut3sajPl2FSX3FLlLsI7CV+P
Gnz/73v9dwEUTT5qLpUaVSPy2lQDLjVMzeJeBEGqE9InDu1qF/r7/iZoGhqDMSZw
y3JhDXiB6hKsNWhE6DqAVdbg1MjJezTi3AOpfW7Uat0x+qExnHPG0wT3c6zyG+Sx
63MP8reoAn7tj5VN5aHpZlfiGejaoUvmeFkjJ8MIdPqjxYF1ztvjbqrAqS//SFiZ
fVfI/wT0JQlDB2CWVlNIuZpdD2IaR13IUbZt9VOn1L8dYJNYMKXAPg6VGnFuNv3s
t4+EBQVwZlMHtbTbF/TTrOKPx4RVoQ2u3HR9UeTjL7lIgs6+3X5yYJVCLUz/OEte
eJvykJNiFWTmbhEYxQrkXNPCczSuLXJzDaQgAca9DfIU4zllRShg5e8QvVh7zyZ1
Uc/GrPJaU9TprPqkdK7XrlF0BEAIZoNQ41V1PlR3qKKFTHuRW4s4hVBDb/YZVv13
u9V/vyjPQyapHc8KZ3xOEYRoZz8QXdQpTZ6Sbl+ogHmRS4ZeI10Rxnol6FzFxm/a
vInc/gw+dVGTiul9MrVFFPZWibVfOAkCEcql0XKPBjbykJ0al2dnsqT9rPp3C80l
mtb513kodY78ip9ZmSl2RFJjr/72IydP395nIfzzf6vnPvYkP3zTlIOBpe3CCpOU
o86m/x61cjaxJZHPPSRdj3+6ryH8EpgpKr3F5q31RuTrcJxfcOA8bhsI6JaIH844
DUBdWeDImBoCtb0EBHLvDhESxdOPzRHGOE3ateJkhAL8N/aJYlVLeDyb2RTk6B66
hN6pOdzcpk9AhEPWjh/Nn2reYLYjL8a0iDEdVoWJOKFTW1WI19gqjQK3bG5KFQFC
w93859+/RUwD2KcZQnDOfZFhJb4E0jhCvLPB49L8DY21OTDt5vM3MhY+mluXL3Hu
cJwR7I6RhbdEFutznG4vd33cjoUxCmrJJCFIehPcqW5xxkfueoaxf9aHczZ5D5xP
x5dZ3x1KjZl2dkYxQRZHmsEylIrvNme1tMY4UPRDV8D9pze5v712MZ+5hxF9qn6M
i/aTvbLRjRofxc8jEyoy7ONDioGxL7cToXTxTnZ/6HRorvUcOkdHjwgG2YLBM/bo
j8JYFbGS9pawcZkIjLp/Da8xhS0KFDe6vPVZLt8l8f27l2IIIDxWzI+H9ZdB7Vt4
ygX4syxUHAXgQykcJIG6wYeiPCHZ/OJHtdaSOcCF0r8OcWeg4ILh5FgJb57vjiRz
t/CuUomYlmmrlAgrEUz8nBdzE+pCt7+BB9T98RKZBIBdT5ssemmD6/Y4aYrJTbXx
4or/EAkvldCyPlTYpD4/QuwOkymHwVZvTCbN0rWY85i35VmTZqb2dUTcifF7BZZu
lDaRd11gPPnJ8UdPcyxAHoK2yc16p5ZPkJ4of1V1MvJUNQy1nF1hJ3iepobNaKAV
oGGb88uI1P2+fcpNI1CMA8POSOmtTYjKbq9l+HB32FvqE7hZ9i8UomR9OZNkH3kp
7dk46AwKhlT9KzkqOY6rigLmlZoIIrL9IioIzpEhzUsQBfp7xdyBqhxNloexPKFz
yG73l7OmZvwmmnVGdfP6jU7esJvAYj314BCTHYd2q9xU8O2LUAGI8xikr/aX/NUI
FoIIdDltEO3uyaE3HdL/AV2EQPrd51JeY3OL8l+T8wFTfy9l6v2GV9iXXXVSKE2j
tHyii7ZlsokqG+8cgBKgM6WqwZROvFPy8tfj7NROocFten3pbRzcMM+qZAiAH53t
IPCyKE/jNhwraQr8od7J/uzL+bnLe/VZHJ/WYB29TwoJZrk3TBM9E+rWUOYgCZ8Z
GcsJ+ckOv3NUv1yrKupaRavDjpI8UxjsTkz6FAxomOTNcHoVWW0iGCtFtGLUH7Aj
wrd3iU1JoxTRrUyL9KgjDFeMf9acfszn0VN2bmrQvgooYDwfHBUKlPWgL2iDeYhd
XpFg8K+XsLqW35lr0zqYPGUX68Z18Z9khOCKRbqY6/9v88wG8z70NKmmMGrRA8Ow
QbPL9IfnBg4CrEV3fo+X1GrUAgOvsxfOmU7XiDYwaujy1sLJxHtHvcUN43VpUBR5
gJ5Vnl2kDz+hYwncFOw6was1CoEAzNa6QW+m121aKn7wonKrFssRZATse4QkuAas
LSA8Ilpt6WSBwem+rQWayseV36ESJl7jgA3Sb9iRFC0o01/RSP1V1HBbJTxXHfU7
zkV773zHcfZytFpKyOnq+ZkhT4l6aNwM/b/u3QWHFkqQQOnIBWgoAK2xbdkWd3ds
RgijzF3xC0MpBAwvZ98pmDEpbjC6lkPrlV+vDxyTgpLoOfH3NKEb+qDYFr4hoyN2
iMOrS6qOQI6v+0Z8VW3gyxl9+6smu8R0q8plcm1es/yS6esjr8aYanSoRz3fDiD0
9ePO0YuTjqUXbz+fO5IWVugnc45KHRyFXe+SVVGEfHHdxkQ9VU8JDn+gb9/if8ZM
tpu8g9XKGn+0vbK5BSlEhzqfSqkjfMppR4U5IJgGN8mZxwFNYQ69SLFdw8sBgKuG
L39JwMJd49WDKlLlrBpjlilDU1K0VWTtnraDCDpWVkEfEZ4mQcsu1ZLm+369uG0M
j4V85eMDvD/rzhJxjzg1+lR0Z+uY9y5fpxpHBU9i2ddnMwg8mHCR53cHMM7LW6X7
tEurzsKLVWltzF7qs3EZMIrFcKIehsVcccFIPhRTrLJPevwxHyBvp+b4xNqzijZ6
Yz4VXl88e2bBtnozuGr0nQiz2XQXcR6CPlj3J0ZkTHD66cxjxgGa2uSlYHRxXC4P
pyQXdhXo0VK9NBPMZQ0pWEMud/tYqJzp2v4y1Gwc1nOzW0Qdsf3cagEcBm6/L4Pj
/ghuTlznHE6XbDo+V5Pqt4HoTUnRMXZHqHU846Q5z7G9fpMbzEIsT/g65VLxjxF+
q8Y6CSjomPWx9gkiHxOCzpVClpeoo5PycAp8lvmeBNKppQoymWTrjrRKnY2Sqmmg
Iyjps2mfyb9/PllaXc8aT4bDQPfIlxOfow9DR7wcx7qeK/G9otlklEwKa65C6uPM
sXYm5y30JLShxG8sLWlphVZOkRXZyb/qHQzpoC1LM1ntqhdN2KOGurMKi1ttJU8i
fQACxqEo7WrcZxoaVNO5cuVEtgkGnPFU9YLtr5l4TFPcIQJrJAcOxw8YNgPTfrV9
G7yQjirPUjUPc2SIGZdki2E+DHeAApc8NH4J7ojGIVKVddboIkRqG5BKrjGCs5xl
QEwVyqh1585MDz64FvlNKfghyR15LSJT1O6oUKegBWF5b/yQ6tRe/TWPst9gSHPF
IsgWFS0bOxYBbNHPj1IDgFAS7gBD0sD2Bsque1j0C0kTv6wEJd1FD6xyk6gObWeZ
0Fdf95cpxMa0hzMYdwMxixdklMQra44RxB8IkYQePVaRKoibEcgjLIiWJeZgkimN
UpCbvwxbAbHx8kfyWzBxhK120xBPAlZIWT9Gvcc0xP1B/PCXuRaCDcY6V4R7RL8E
NzCazSCDu2DolSjPOC9is31uB1LIMOcPs1maJxJtcTCKSvNCOB+1JEEcemX68JMP
nDiyNYcMZ/n+6cTfi66S3jrDCk8ybCb5Ivhxx9WW3sgiaSVXBDN41a5u2O+KhVux
Q/jmqDLzuLuy5M2lAoVYTy6G8HkNE3/v31P6/zxUim22WcfI36FLDlVw74YC26en
MvSyqZPyBbvjk2AtupcKU7HfYf2saaYikTakxSKQ5LqScX086ZRxT8NYZ1yrr0yP
3gBypTG1MA4bw5V9rnnqaII9xB7WB9rQK90uxLMNd6WDTviugIN5scvPkrMTpxlD
4JXDvB+fT8qU3z6kpxGfib1B1cU4YT2yVXvM3sScLnRPqqF7Ldu2/OqopjCaSSvF
mg520CwEa+KIHc+R0SCwnYkacWZVjWj+MuR1q/Ef4t/g9v8qQ/oKh7LCtE4ujGMu
K90wDAqQM2XLuTf+giJKEYn/72CndJSaH8DAS6OJBJyda6WsEHVSQoPT0WzLZzLg
7ZZf2BbM+j33IlbECuBSGS83xp1Wn7vLZUamAUzMzKthPmwMR1/gIXUA6IeoaQN9
dkvdcypvNSh8wSDuWwxYrdzXUuT7g4wHk3lSzeyW2EMgXywgikb++HDi3eXtjXKP
mJgvVl2RPE2Bzjuqa5YKuZjeDNrbfppFe+yWQYwYCysJvlj5dSnrDtxkjYk6ZUKu
/cNcCO4oTc+HjhzAYUWVHTXUoLNDZeYaHkYgz2NWhiwGYnAWr2Oc4fIoQFZJ0VII
h3O0vsrmJSBgiOvz4HiRGTqcqRCFs4p5/4BPrD4YmlfmCJvqjZRiitxqnOrFdGNP
CIhz/LJETrB8n5Etdj0jBGxDvq1Kobpd2raZCM1A4Z0RxGt5H1By1lfQBEqoaTJg
Re/2cXBCzMQF14M0JdjUJms/Vp+pKNbWO+iHMfukpbSX+Tfy30aHOircpGQl/2J6
xB+/++xWx4xstW+s/e//cQYS+qM8d+r78bQkEk3kSPuIdp1CrcKDSs4gIeYmw6JR
0gnkyCya7kSv+iGtpSTf2Atdql/5HMgG7qK7Bc468Vs6ufa0ZVZ5u3AVJTEs8ye9
Bru/19MACqZtQctJOhBb65FD36ztXRL06UD26aR3laBBNLbVpoVPK4+2bJk9LSNl
UsPmBja/CaFew0Ei3vWki1io113ZuyxcNbIBt9WZ8RUNcjtA3RZbb58z7SRJhkPg
vN7Qw4m6HIifDd7T3P4Hq9yQUbGchk+VtUmLGZ7P7zDwhTBcvW0l+0a5LLod6P6D
6RPf9yer/oPuZ1eTfsRK8/eGyrIz6TLb+pcpt/dQpMdpa6RthhDkvpJFUhh/NUmQ
+RWP0wikd0AhGYnlYtzdGOqVi23TP+ZbB2eg3Sc55sjb423UOY8waMN9IyJN0j7S
U0UO/qmSM/aO6SoRwT8TVQ2BzQKsvEEQhEcWKjvDLIcmypvqoKlas1xU6ijunbi5
UYHADAuYOaaeGjhv4HkzZU5L6lATV45hUmFB+hJBQd7OHlEbemxj7nsLDVIJnzay
RkqJu1l10xj2Pgx2YPeZCxhSrZvGgskAnLKAxnPAeAf1o0uWcZA5aweHpt0Whi99
tNOv8EIGkTGE6kxYA5k6u4v2DKv52bLmSupsR07pHfHF+CXpoZ4pVsJw+XzWt2JQ
YXPQOvceWpavo3V71D7Y4nztpKHkroPSOmFxmAqa9tYoDucEKugPIbSKygd/ekXq
K5khZC0CjDp7UARu60xuzZpmVVecfL3xUUhe4y5bBdgT1OykPncOxv7jy6Zsw58l
U9lYqux4iBvptZzM5deOGSoXrQ0YZGlIOm0jf9BQrrPqrBAOfEoopee6/sYexL/9
Hz9be/NOyzTgdviBq5AKMkivn/xkaIYV+2cUqxi94bqldJehxfAMayC/Fr+lTHKi
shHIk3+ZBdTvGFGsl6IbkD+3rceDHkk0ba8/s/XdLYE4Mu9A0umoPXBMVs34k9Wh
yybmhSLNUaEnUZjeUEWrhtuaPMxBhoJ+F72yY8b8Wt3+p6OUv0BUQtnhhEnhFn8L
pe4e2eFrwe3+8bROQLdo/7kJ77Uoceh8U0d5brqSQCc17BMlBuM6nYLO3G9t/1TR
ZvoCzH7ZAyvUqkOCNhcjBDhE7yiYUprvjO4Z7IG4i7xQNTma8gPwNGO1JdCgtfKD
QtxdHDi9bJHsk8VL+g9lWaG3nIPeGHGtP42MTxv9RYehjkOWDXkInCVkjU4Twd9X
l6ip+Qh0u36L6MZS2SduxB2tz1mWR2xJJfPB8NZjMGGkltKdRUkxo5FsVHjZPu26
o4cZG5DCQ7HvBdvp74I8VCuZP3kuSs5yi26+C7NtLOqxRTv6+n1N88xbX9UXlj/v
vpE3cYGL+vljMB9ofJjXWEVHu2m39poBr0veVXoOHB9sTvpR4mVAPzXER+FVowJV
+6eUCqLs5NFs5QKMLM1g0Qh232DKPCl0kzfMsexpFfaE17w5F9q6feP3FMHGFaX4
q2jf58+WiZWCEzzYh0Bi0C/ZNy6mgM/P+GkOxPyAcSluYZ0ZfjHO4Nxf6QhGJIZE
0TnOHJgbOZtopQEB6Z1gokyRek+AjvSv6nTj2je7u3t9wyLHaRJRY97X3F5GvyKG
KrFcTqYDYBmDaVnd8RvA6NXT/z4WWr0V5P6R83ljtDIHl+9Z41JwCbZnbcE5FZ2K
vCV5TYKajPTw4I4ZkzRy8ElAMpEL8HchtezmtGfTuBx+jxUWQwlDEUhjivH4zcQW
qu95SYvG/URXnJ9/50dPPB0v81WXVxiqnhMOqAIQ3mjEKyoUDIIIr/hq9/VjTFXa
291ugvqcchkIxWvX/LMwij07d/vxJ0tSd+2U/pQw1JykJX41ipkGdGLX1Eig6qdF
bRjl160iskqYUGlxuMAhuE/RX3b5bFScLONeNFRLB88IcH2OBg9aMWz9K/o5bwqb
1fvR5Sgk3m/ZyZ+oN59dOjtnLmyf1moovgzMg55IQo27N5tSSvesKb3pUGLgrQ94
yYnO9bZstq7jCokiOwQ6soS0wRDbdA7n7z2gk4mOskRfYzu4I/opXwDR7bthX5dk
46WKxltZ2eK+sW2H123x2NRuFhD6NkBy85nZfmz/Hq3uv5rioGq07gzFr6K6Rmsu
xzkG8OlE2COGDTijWDrRplJQr6A9APXvC0pf84EBbGoeel1SpuMV7qbsfYOeMMI9
69n7J8XwQpsOrLV0YAB8xx/LcAKSc2vuOowydTAV4XjwOrrU2tDlgpD/zKKVJBE2
Ty58JsIELfLdCFe6HXhydKCzhD7VqrWNIKkdBSqYpo+LhZ5A4gafHRXqZa8WPyyE
VBDNG06z0IiRgnKOjqDSsTEM91GLZhl6I2rFrGITy9SqY/65hGirJNt6gTmwKlTh
opmjiCVWAG/qeniX4nK3qsC+zgO/xRk8e/k/uLEmFx0PCwwB7jeHTihWyYu9MfLo
tXklvnOIau8HccGeKdhrPW8g+Y5XfX4MIIKrjTdGZBMhfinojYvQQUUH+LUOTLXs
MWCvxZwUHdLsnB5wBVrpWpXMq0v9xx8DZ4jIySC/eGCegN4rcOTRBjIf4UjuaRi6
r86OQgQV9hgUXTDlBqUTIT+gWbH8sq6/XQk6xQr8wUViemeDMhM6t2f2kutUXvFn
HJEL6mTYRINtydRoBzvr57RQCtkUsLCbXXFN6oBNjm/e5JdlvYynHEvYty5S9P+2
E/eo+O0RAERCEWo6/GXvTpjb9P7iTMUTHUVEBBIM/+7/nHgUAQ97EMhtCtbvB7wU
8Fx6HKb5nCU7ArZwzPz/OO4gh2eIvFju8NA6NIxiVYhxu6ws57DgJua0dxyPhTX6
33DUHtGunJBR9xbdfbWuyYd72CmgZEh0h8uqPH6S1jm5ZmGQIqChDyEsNgD3pb3S
TsTkXmDfYqY8ydYTssragPdRlnAnDkzQVyXKE+STMXtNB9MhQ6+rs5QjBDs6QxHR
towvgbFAS8cojyOeP6VUawK2TVBJ7Ctf9ejjaL3D26Ve4qUrYtmMofm8sUVIf7wS
5uucu1o6PkYzT0xCXc4ZHiOIXSZg7SVZ4FeuwAobf1XaY8VXhqYslHJIVcEaz1sE
8Cg3e0Z87GmzuWEtY0++1kNDAxEkwH6GXRPFBEr20dekeFBaV+621MiUOQgdDbUU
pv1RPgYKZBKXtE3n8UwBzNMUZ7zxOJu9fVScdWq+vf8OlfV4jDGa1dLpsbRpkhLL
lc5EqRqlPcv+nMpaVjrKi07WD64A1ufqL/SkLCmgyB6IEIt+qDIuhtSue6GhEsXw
WJ1QCPpvdFMfCzlxfCQ9XthEQTXijVovcKBLwMrVA5Ia9v/bQnFALrg0LzNwEOBa
cocx6maWNR8j/59f8uRvrO1M+w+M3FyCMBlrfxUnKJumT6N/7jLbrVQUQLwwOLl1
lf+0zVTnisltCpdjE1nBBd/eIp5N4KCpTdBiFx1ubcybpRVkYFxBH8YFN1zwnfKx
XM8rebcVKLMYtzU8lBGbpjOtvUp1MnyxRd4B9rU5hpBOuhX68cupk9JTRiZL+Y62
6cAYm5WL+voRDdUZwIxpRAS/KNlebbiMnI2LPlwR1BsWytvNoQlk/BD5rNIPCIjX
WR3DlyA3I3KCXrECCQjNO6I58GNAJ7jumqGStmL93CHRIdA1Nf626TXCbr1A12Rh
SiMr6rCR3C3uWL6X+i1pVb8flbTBPf/H0sP3LwQErCEWx1Ik/xXCt4rgJ4vvv2Pi
m8ED7SMwo9X+j1HHCrM/8kw7hMwq5D1uxkkJtLFDchA7taQEpSXfNbkIGojQpIm6
HCNwGJtpMoLSLF2doQsGaDu1fmX4BLX1UqD+ZCZVwkujAAd5ONxW+qKf3XtfhRsP
MU/ZqGXYf0rEcjcpO0okZG8wFYMkD+h7t9jkAnt856mclv/aRbmIv/iak2ZsfdGU
A5HAcyL9fkp/3YL25ViY4078VZ2LCvV9h/yjQE19HpT9Gt8iLle+9gX6qyQj3mrs
UWPDLjui772NJxwz3O2gkIZEYwvJ1uizxzOO1DnmctmrbNU/aTGh0EFwpiXM5jgP
Cq54GBA3jtxqGSb0BIPdVbuTAZI4yyRtlfNvHcC1TO5dvZXWMTLv0D03bcBG4yRQ
69g5EN1qao4q7mesiJLnI920Evm/79opYfBBKP9pYMuFGp7vGX+EwNnv5tZYUd5j
TICJJaL/xOGA5FG67d42RMa2Ym3erQRD2dECSK4pSzbKQ0p66zlodqEkx/Hi14fE
7F/OQqwCryKyG2HomYc3L7jGv7SuSiSY8H/fSuluf0ClMz3ybj9hk3S1GnWbZ6da
txPPKG8aIlSdN/a1m8NNxjbvQhPXIFzYdcRRXpLS//GdBdmbj2g4mI261otyrgC4
ghjIseZtq/DSrffj1iOooZvMqCdF+a6eIt6rMpsgIk6FhMYi6KmSG0mLuYKZqE9L
caTT/vAFsXGRp1fClPGVESeFbc9NfTwqZ05xDyEyacn/1F33bHLkqqYDWkyLvF2R
PIOLbOsK3zHyiqZt1Vl0RkcdPxWMjzEXw16k/rr5v4D5ou0hcmiVIC8TVtfk0m21
lqvXMW9Pc7meUVWaPXg5uTFLPwXmTY1oNl9N34elfZfZB8phLgYo2gG5u3uu1bdk
sAbl18eiMj8P+4gHq+g1V6lNlgGkjoSk/GpiPhV8hNvFYXjlEHHRaOUhR39ChCff
IJ7A6vnGkGWR8FAOKL5Aye4mzrZkXDoF1ViScCfJe6MpfgvHDumgumeZGHGxGLnG
jBoIGmmIM/M5OIQENg4rUsrM+WFBzY0pChdhcCknW6m33EbXeF1x+qZq0lOwEfIY
wnUwh8cY4pInNOlwug1t3EHTXAZGC2KBofxXLS4J8e12R1U+pFyTzjlNU6PnkIC/
Q/FWR5Dne6nv0QAOTjUsYP/jfEPVtYT5W7X2+bK3s9RM+9dzdjdfNUjSGZvwxb2j
r7veumkzt/QW4zuPbIZcq1h1/+qPFGf4+Gy9vHnS3Jq2AxNag9y7HliJ4u/aFcX3
X+hNTUgpDJwoKEE+K+MrUGoUblv9wYggTMuVRWYMbJdmjFXXlhkfeODhxVC5J5fa
AaiLb9rYMheJpOHaFdP4m0EaRJlZEem+00yv6PRFfv0kcIsd0MV6fYR+nczPVUfu
cnVt82Yq6P9396MOJlaTVsz+R/yI8Kx6m1r+vJcg9t/d7VskVVdtIu7kzHiHg3Uv
loSqy4Wx/CwqLnacuOSNEPFvOQsDl+zBFwJROEpQ8EKWc0Ld5Af+tQsT/EGiwBlC
GEgstNB/baGiUvvyHAhtF8+nv1DGW2q72If54petafvBvZaENo+v8CmjXE4wkUQA
Snhj1aw+7JTQ5tga5HEnl8f3lytsvl0TygF4PXoy6efKZ5YUr7Jn1EnQN4h2Ka7M
MqepyZntN5/UT7o+qyxzo/JMzRdTkRz1V5f3+Iu/LvyqCwhanLnxITErU7lw2IY1
1VeJrZvED4HLSuEYtVafe3JSnVsG6y4pTtDsGzepL+4sic6GE6hjsSgPCxcj3tx1
Diwn1KiAJYLNCWwl4LSxYBrrx0FM5Y9ek+/EQmgW/+FDdyJkliMAF+ko2XwT7KSX
peBaG4+O2JtN6QUNqXi7iqUrqXvGdBa+nfnAp/XGvOswXWLgwp/Vt6GPPYoYclUC
PMStGXtwFLL4w0VEaC1i6FwlP5Qae041nxhcxoR9WP//J1nmNRfKHRqCTGOANnNQ
14kQgjXPZxgpXeGk8SFSQGhmJxeYoRJV5qwTv0r99TGC2KdB6uCtXx0Rm7oMdTHo
kyS0tl1RrZA+DVtZDddw75aeTZzY+lGAD5zEX3plkbS/WYNmw+pOzhYovMuf+E5b
qhfrcZcxK8uqgacTMbizhTmYKLRYzPxQgaaTznQaefC+cOkYMO7TjSgwKITzrqJc
0asSGJqOtSxgxKWO1mm3cS/6Fn5ZRfc1bEdlU1ypqW7JdwiuU4WcAD4OCLLSdBwZ
ELklI0ymKfRk3cU5YqyfzsW26s4iQmwIg+QTbfob9fRhGmnS91W7rTWQwx6p70MH
Gd3mqTeXwtaKlncJGE4i2Lu3Ot0HweIvyJFTpjIdsZLkE/vpAxNuQgZMj0i8KiV3
fhWnwVwybKNqXUqjeifiZxTUi1er+BYoIIRTzCeRiIfUqMg6eRQ+TeoX+zuqj2di
lQBFrCb4dyxW96yayJY2Z9BUaCve6l5IHXvrnlowjj/PwiaNMds3t9KMfDrPzCao
mx+WIf87cvLjjnjQJXHTta8r5JOLiPpo2fenjmwZ3fM8lusKPOzgXXVap3ITD0ip
IS2k0xbbPS/bMKRhd7QnnjNSdH47aUVqx/Yv4GT/08JFVvaoQtYqKVXEbgv5tO6a
xlWofKq+QvMFPOGVb3IKCsih89pKlzQ1QxvGMGS6X6v/gkz03uLWV9HgOVuhF4t4
dZhymuwQNbcw2+mQOXSeYPZTELI7dNrQbHaTyUcnY2OQV7wpRx3OF85V7qbdTwzS
KOvU8QBr51XfAYmbw3H7MS9Rgj5xRi+tUjlPJUfEvk2nIUyydgg3WMJgeMzLeNf4
bPcJERlLdSrkSNRvWTrF5XeR/vvFX9TzVeFsMc0TlWqJ7nja0UHH5uOoTK3yDpKD
rMzJjHmxvV/+M+qY30SxdzaVnMYY+h688VOp7LkP4O3Kqge5jVYgOhUZEnm5vzn4
94gFzgdVhPxPqikB8VlPQmOLr62jNCHKU1+tBJ30T9WF1LA0JzK++OdRmdjECFxN
L5RwTl8QVOTaElsMTItWBqTyYS3k+jBRG2egsIoRBxpFvnWQpjUfkdZOPpTPBvI3
+vZhfs3ldEZ9uzFYbrISUPl5RPH3uVhH016nOehNp0TxCjGtiwyoXQkYjP0CjQnr
BD6oSRRz8qfcwHOsq7g4TKfpCs19twOXlM3Pj5gBypRlrYKI4Ftsk00JW6n1Bugs
q4P4Wbo79abh2qFVgUAE1WoNLMGesmd3Dblu+ZX4lSN5u3YgYnP+kJEqSl0WlVry
PBblQ96gPTT/DskQoEzUzng+MwjQwO4xSwnBpNjjqvxYR4C3AwAvyys/GCIkAYLp
SvumGbXPU9EevNDZzEn4aaTXLgCP4yQV1QJWojJN5nnhsKKPDzqHOcYqhAUGT43a
TaWq2Zzo7OxacfVBthFfgAbJbDLYsnz4CvtfW8rRFSYh4vYDk+o8C1oJzedQvBv3
LN8na3kdhSZhcwLKOKj6w3LRlB+Iyb+b8CWxmAaZtZqoC+lLTuweFmLUEXvF3YbJ
v1MGFA1r2QKkrUothdMov27M/v5BiDprAGhtayuezBQs1zCLrU4AveJjz0kC9fkV
Ade1dOFAZnkTHxD5X3yB182F14h+mB7dDHD9tT0n+ZJfwOh1xqByiiuv3Uxk0nII
BmTHoChW006y9fbVZmPxsGhDP5AlIriPIk+5MEey6GAlGiNyzl2u/lxC21glOCf4
8Xa4Obbg971FV0yz0XbyOR4lpOD8C1reyPw65z2yXsGim4Gum08/RYM0SKVG17hJ
0auUd8CX4PH3u+fhXcyf0y3v0pGqGNAmf3egyHoKhGkYomtm5MR+dK/B6Ry5M1QC
EggIAabbXgYfEyZAXP5XIgcDkmnS9viXi+rccgpA8gJXRoPGfV+qh/7BL3EPZDVO
eQszSWSjY9KNeKrtzFFaiX29v32PZ2avBP4uwOshlLs9lss+twS23Ky1Ws0PSxNc
0XMrN1UPjJ8PaFjeVybT1J4yWLBmHJYsKtpai+LPTUp/+9MlSkqCzQj/RigFmHGC
5QUiXGhvXpW+l+c/TqF/x5u8KZIu4y+5NIxhxoC32XMXWam9KvdJrbz1vBF8Jkl1
zta4WMg+GGXQzdJWop/XYHqQK5+nAzyFX7k2sV+WOpS8VPk30DrnRTkut3mQ4KkU
CstdH7RgwFEk5naYDeEYbdBYLnPUeaHvN7tHAPkUMzAOqxIiVnnBRPWlDK+uIHTs
9YnfPJmt6HPU2FZACIwbXRcTFee5jMqGSx1r+LCVqg9s9Ea/+hgfYXvUxazdwThR
y1jktvf5dmNl5rEH1SqSlRGsSv4rSBCBda2FpLD6YhQIvgZHb2QVaNlQLF0k3WNV
8EjodGBe/wQEPlJPYyvnRtYBm4YZjdlYAYZdIaqnhDYjPzKBhTWMG/fPZTzS1g1i
GGwxIwpKegKQ4K0WVuKYzsuMV8CTe+EJRDxmLWYZesIxF2y4aWzkU2rQlI/+t1oi
Lrn12xyWeC12YupA/5eK5m2gWW5MRw9pPlfa6d0NnTBEGasdqZfnwCfoGoWkk8Gb
Rb5KBqqnVyTzf06PJy86SPbkmNkJPl69iTem4RvkgHY8bPTqbj3WuDYEOCUdTa6h
a/YNRKaoGAbmXVOFdufS0IYjwCeCNkhVjk/tlXadoiTUOkPHdvjKISliavg3mLOI
s4+cgTOd80X5GEnw+PxtvnhWI3EsTAlzQcKBZuKnYRpnaqyj/vfgorkfV1pPPI0d
FaiIPtfnpyaCquDtafn0VApgQjLwFY2QCVKbqrYGNkpTFJLbwc4KqQ/zp0SfOuOj
ItRXkjXWkZT/o6hjChdYvAGOrq9tcqKLEfR5qLTu/rBIVGWGdY+j2wjDzPII6TEm
qpZSnPdbZBIO3/Q5/LT8nKM1nHKv8wbNotObZmlWlVUdwBKJ3NsaIht/Vd7fYbF7
uk3HJVQiqpbCC29TLGxf+L6oYXoEGfLkkFaVNfkowhS/qXSgItOSsmfKdpFCBHM8
y2yMLfiVowNy4psVp4XQ08HzYEl+tEwnvJlUsRfrZTZVZ7gIIZyv+t9wyKWDDhar
McvngQEkRtla7apCpXUzjbBn3EjWuR1PIx7B0J0pkAH+VaHbCxYUNN04y10I+sl1
0YVq5vfk8LlCwecmIaM6SYFZyvU9pWgL1Z4UMLrEulZYh7saysXS4/E4tkahFoeK
fR9e6bpdX2p32krgxf+pLiXLPlrwBnxnaFI658PM1LtY6chytyxadAWbTP5x/XsV
QQOyHcys3sFwhIWRpjS/7hViuiuOmk9rTVAem5iH7PFzGi442L34KQtQoJCXLKJh
MDwEmSeJAFfMJm5UWYpihrRRFGBcYcbk3Gnrt+7ZaAQXz8u+t9ZJ6QOytEI/PF3z
3aJTa2tif+PYE8D6krFboWt+NHyq/0ASiDmjS9vXRcRY259uG38QA4OlgGLR0tmU
7BLyfU922PBkkzn4cUFOgSG9hb3lbhLiviEVGsxqbJrX72+DKfWFIiH6T+fKFxAd
hTNFpdwAFjCb+lto88aEj41Pf9LEcjaRQnXAMapkRRGwuRk9Kcgrz9Vq+gU0jcJS
1iXamxojsm8EPHzc1jxh5iQv02oYc8ax9ZmzkGu5hpIsJ4ECsV4sJTRIouJIDn9J
D1W4bd5Aa2wZjiYWSzVSRqgOqTJX2lC1XZvAImZjF8pZcG1V+v7bUCNacHUUbcwg
1/1oDPlBuoSHrBnF5ln/S9HWEdarzs1NmN5pfcSWJ/kNLBUMQll7VsE+XxIMMNQd
/xMSBbDw0lEdUA73P3DsSQFUBAZpK1DEyA8SMcU8JOGX50eaMqRkDPygSW+wJGjy
hf0XFd9mI6YrMb5G4SwbdpDTpOapvrLKYLW4MFGD43yTOrA6b5mSix5/gZOiobZ0
bWT6V88Q84LJGCvzGofu60xrQsgOitzJK2tGc+EvaoTJOhkImu2V/eFMNRbwQ9dS
qecuoJHL6nA6XSYgVsPmAV4WM9gpn+7vy6x/26jhwkXMxFh5kheVl6/aM1oh8act
0+ZavGqwSll3bREAcRWiYgMf/AT/bHjMwh5hWTZQ8D/74NgGV/zxLB11NsNxuT4u
XmB99ypbRuurFXpnCsmgxPo4PkceYdRrv5Hm9bwCDPMtSNTYVsZldtRjHkjM9ytH
jwZIjYqJNd729o7MG2qb/7pEbOk2pmhkc46PjGRsspuT1G08siPrIXq17P2TpmdF
9cDrn1gya2pdUN0Kby6IcBtfyS0v+SeM/zqFBFXuYOd3uwDbtndfhrAk/DhKLtl9
1NMdax+yhsSlIo3fQ7qLWpXmPOLvyvIthIgravYh05/GRsw4iLkXl8H2UssKn6Ki
AFaUqEu3tb7/a2En3S6OyrxT9auW/6/AZI8eZmPcqHuqEC3VbPE+BVp+pdcvC+Sy
AzkMV9FOhJqIDVUFeVYXoGUFxLaE51FTdvaJUlRaKQYdex9/uIU/xzpQIdwcy2Ci
vpZf0eFQpxgQdGSasOIhUp13Mh4Y9tZfEhkoZIqB1jcpih9wHyBFg0BV6xqd+4Wr
ao/UqZW33S9yaMsdJSyp6vmIPjnITatNJkmG0TkiL/CzZqI2uI2BOsptp5S7aZUo
rYg94XFol+UlRBEue+qVm2Vn/Rai8EJCuZ1g85eZVdMQeoYthc/CcgDOCrRxID7Z
9HGRgnP6M2pA/dhLUctSXb+Gac2id/U6XaB1kkG4nF1eUb/tsEzLX8yj6bwpbaEy
5G1Xp0dPEGZTUu4i0yw0MRAEI9kWZCdxD49UC75556dVgsXt0ctVaSnvGOJnpMoa
VPcJzdR+H5ELDJUgWsFKWaxztqZolr1TNGjoVcfX5fnOVoJrcZl5FJlULdidutNh
HD2svUwAgBZ21/xP6kI0JuANxjZBNljBCrYyG3WnMGYmjGs7f3LdhUdMsmgwt594
hDl1IcBX8o6iC95lVKu86FBNsul+BIXBuO9+I5BrGLCkJpGuDmZ7H49XBo1n8PRI
4sDKW5fTHS4BXop7ezKbC6txrjpddD+mLwDAwB9GMIDaJkRYjUuMeso1md16k7uk
mg9xfqhvfyWNJ76mJcbaKjO0pO6spHl5KM5EAg6GOUVxl5LhAuxtSVa6aes7AYey
B+4h2Bm3GsccOzekgkTuqV0DunLev1eaM1B/7W/4ynhHqUSPTHi2LnWI+8Oqk7P1
zkQnW4dpCl1bqfVIzYYVG8IkqO0nuJ7lxOHMMZHWCQqB4ThNmDlr8ltib1GW/v5h
giyrcaLQJ5LN9Oc44tSETUUrK13QNgWJpxl3ZO5hpB811aCBsAlfDN5Il6q5Zadc
7l4mXoSdvtTH8Hd0z21Bi+C0iI8FlR1E+YMatknQRDVVwwBsA6mGEj5JKqP0awKz
iG5wtA5Uqss98UIpEIgpMU/UXwjbDA5K6FWGtsAfe2UoX7tFTDOYGI8e1SOO+lwW
szG6qaL7OODFjLoYlpU6l7MUIXexTLlyugZ7bdxI0vSLQ1vJQIdWD2l5uqT1LlVp
gMemUICHICyPYz23j+B6kUHcQzkCHScdYVZiwCG1DosdCOUjA38vod0LyXGum0t0
0Mno7dDctTXMg6NKitLrfz9gpOKnKq/hdqk/ZcLOEGMJKdHue0J9TRA7C7dg6ZLb
MXvboPAWmOR5t6luzKUIm5bSas7cjF/z6KIAPKZTIgaCo7SjYjzo1rx5PjyVEBEf
85T76I2k19eSzzSTpweKme4KYKg2VzuCSHua9KC1cyEA+EXZL4RuUSyAmSUsMQ7J
JqzHZz+Rcr8iozX5AMF9m7i1UXc0qJPhNCYsNn37a0mULWV2KHV2N9ZaVjZx6Jhq
zFFZG8BXg9g+aXrafnrvpu3ez3aPoN1DyjGnUnNngCAwjOy/MY2m+OnZ7I1gmuqT
Df+jikVqkeTq/HMG2zVmEEK38RxXPtQ7hGMUCzttI8bmekv1gL9983xX+giiT+5m
fuEzMTjHxkXaeywmMurfmYNyi+cxaT8/v12nxKnYxlQNbVKEO63xMvkJMKaPlc5H
vhVmNl6D7pOuzAxXwMvGMmhryR4Xr8EJEYWHon8A6zk9R2PISAEaJjofOg3d1JaL
wjdHTOJ37EXb+rzUjPMeYSs889O6mioptF/Th/QeBg3vNGb4F01vOJBa96bKoo1/
D3Q/ZXwoBTas7ZCrPXkSV+5eaFquGF2jMQ1ZyHVG2J63YlUKCW4Z6VNqrUfZisZy
72tJnKzzCh0iq6vmZ/QCplefSFxrjfexesgbQGZBlZ7Ruhx5e+r3urxZDF8bjSCY
9Dsz6E5mmup7P1ORV43BwDKStV/DVY/PZGFeoxlY5h4K3R0VWQfgiN05xQzkKVr8
//+JsnDSvrzBcXQ9GOS8a59hC+2v25JEBb//CfMG4cCWTgV5gcKDHs+61/fQzoVy
z2WUAnnDDfZbSlqTCH/1KpJjipMNLsZyCLw1adKBFDuNCf+QAS8etDs9CW6wUyl8
PiKEjJe3pLFXjScV/6aEUNFCGcp8aivVLs8uw07vb4j3YEPpwRRWxlbEQV837Mf/
3rgFT34xNgGC37l9iDSbkBPC0Gm6fN40CMznFu26WpLGsLn1X258Mvp0+s6JAKnD
rA7MF9tYNcpXjrlFhAC5xK9GDd28Joeptq46Wk9MOQpLDIjI0UDcjO2+qCobY1Y8
IRWrHdVbcmhnZZxiZidY5nsi13pYaa6tgxdeG/ILM+ZKkpnvIjvaXn0S/7c/l8pi
cbyfozUTYtjBabm4naLRj/e45NKc+YLd8M0tVZPJV3PQMeTxjl15rvt4w3LY2f4n
zyxUlI/B6LAKeR4b3KW/lNlsvbA3V17BUuCSuk/5S9gDYWx4X22Im2uTxieIWCbg
vnasUQSSBssrPcBse6rUohmMaF0SzUfR3D50AmKgsREDo2p/Sv6tK3TqQwU5xHOZ
dR94PLNcPT5xCNk+6ZzLWcY1aeDVt0hrSxDiLcwh8bMtVV48PSbS0eS4D2nTw1/7
lAG5rtkHGGsAikyy1//u4NLqGlhok63DQHn6PYICOeWArWTHA51XhI92I4dhflk9
mMN8pTh6xF2Ts2V2tHPZCPbuo7NSQoIZwGrQeRvfAYGkGYTyqOy9ipgm9fmEy3Kt
wnKom3gA/J4vBoV1HrfONOBA7yEQP83UPRj3G0hcOCn5NifcSdrz7yVSmkXKSzo7
iI8//1I1mNmIPPFEW5s3Afb1UeQR+Cy/5wFjuDM5i6XaPti0N/WObbTrgDGkJzVH
o8TE/AN4AS1QniWlgqOvGhad4GHxs7Q86UosAAWxM/6CruaX7kR9RMFzAK6sd+J+
1Znb7JUS0PvCfaVxYMKWowjsu2UJalWgdz1Bmt41oaUBb0T7n7rpCKFYFjBXF/GH
chkeKUylUGr4AIEDPP7zl7VIGX9jbbKg2deOkPDtldfJV/XV1K+VkCIsgRzb8/Y7
hkBe3Qa8zk+C64r1PQa39aWtGXIDMDJVxoT2Jnt4Aa+DfYnsANRfIEXW6hKZUgIY
PYyI8dAww1N2dIcM6odngNpUQP6++5SoKdgPnyMlkhuJg8irg5/OlVB/kxRsY9Oe
h1r1xD0jyopyTiSCUFiYAA+XLftU4xXHpct6cc4i1PvRH9EBYZfI/aOkaau2v+7I
N21e1ier3aHWtiBL/QT1qYKP08b0tuFi3AHWOQu4q1/cSisFjzTvoyc+iEfxtQS3
0CdlPW1cXYKMK8PytRzQVhAr+IiX3F6o4+fCvC4g3DUglepXPsTveyjczWvZbDdu
VAZLpPcoEaQbNeBwp7/PRH+IjRCpbe3FmImm6wQX8EUMp2tQDR9oxF+TT4kyNEyC
fwjTM5wgmGp9iPNyyGaU+vdON7N5P7+iiEgdfi9QZyV1PDVhO25svXMOFsA+xyPR
Nmf1QW6QasJ/m6OFZVdYNq/KvnAzkxBgsWU1s26YZh64k6fyGs4cv7FHUSrWWvXW
ZfU4FX4Q8PHAfx3nJhQJdr7kUs94o6rWrYqv3NVLUP0xjUpsvnt43BAqoJOPQ/+/
dWivyYH2TRslelAlX5jMMz1TlzH3Lu3RoqXfPg38sGuAHaoM0VKfypQC3tZCUaZ9
PNGzQR+TIGnvftGVKIIRGkiaIPAx0PmSb71jjiA1CzVL5/A5Uvrml6GYm3jdC7vS
h4TTaINeTmt5dhTHlyf5/+EJch7wy4+VS+G7lhq39mEKUlytySmEJbjFUMMbcspl
/1kYaZn91+zYGrNBIj8Vmf0aPJK+1kMNXw2uKhuCEf+lUfQ/VX05uLqf19BC4Bvt
UgkcPRZizpAkTwuSkh9ilgkRhoalo6FEvA8HNX1Vg9K5rOyaZqTAP8wauW5L3Ckg
cLqsMR9jOEdcNmAFIRPjXONDwrA2JoqEEQRwM+ctDuy/aLs7v+WDXc1QKnRHn8cU
SEaayGhIUDiQGDl6VtNJ3pXmLaRrvW+4sdrWBj+FNvewOaMDHKdi6vPJSfTNhtYO
L3ec1KkupDGQKUH/dJ990FZ9XuS14xHNy8vNIIUrvHANfv8Bi4wAYf0ME9UJwSEU
g1ccrUv4hi1GXpMK0HOA7fvXvkQJ5TDX1GvT3HgG/x3LDPvVcNl1dAaZuCD/WTFi
wT1FPTildS1qMkhiV8qTJPXNdrKHbGMZu1FJ7bmEH7IlGqJNo/o/Vnxr9rXcJkK4
/m49aPE5YbEeEXkNvy+zgK+fVgTIil/53IFx6qJroGe2B5rrEcZafV69vdHz23MU
ynAoRfsoRe54M23b+PbJ3c5O8CS4hVKoW9UUzctt3YXL4ja+AqkPDTkLyDYBaqZf
i8PHC4Dsap/rRGdN35yBKJlrL1eUNSxeEtbUd8gCsGr0a7RVL9MwyLY8vMCTjIUh
Wc46Dvlw7FD1SEiemXormgqwiKoDs+3cAF9Jwf/f1oHXYVxkZB49z1ayyvDJavKK
w5DgI/JC8kzeHU0OUjslIaKkwnhSBRModDl9aF81uGxulpUG2gQapt+7JHlUbfvr
oCOmR5glJxmNUws0aCUU8ve8MB21/UE9efwetl3KubQLnLToIo85Y9ckRQThs7CR
g7oEsqnfI1vu0IkudeiEhknR+xEbQ8jhN9VWYp5ibPiSNhA2Ab21ufYReXfwlHWF
2W/i2mvbwcLV2wPLORay5zlI9R+Ed0OoqQflmQmkDvZ8OwswAd0Vvbj787UEXHw5
HJkf9N+DQuEFi78ZV2jTirer67+5J2ItR5iyIG+vX+7QGdrg/o6Ulv5Ew9Deo7qH
+8dBOQAECJXJVjYEvWLYUIErniCR58KkMFAjflRlUXRsYFmkaME/wvKw3N5TmZqZ
PEnn4xS1T14CUnw9umcxA9z3IMv3FLaT7lMXkf1S9G43iBk2MNOHRTKM0om5iRO0
+ufd/7+Gxog7jXX4sBkwqjzVUx4nu/HCTA5OxKRzm2c0AgerR+lZTUXKYeGQys38
Otp7XN31fdl9Yl74bg3yT07SdKBc9yhbaUldC+1Ihl0oBXD+t8lYqxzkU1rJK2kQ
hzME7mKfspxV25c5Cce6t4p+6IDyyV8R9V8cxQSVC8PW2He9ul0hSOsfUPsJuTpD
Z58LH805DHLEMi58/Xg4FjwoekZWpEiyRRrNLuv4QyJ6bHaMsRP4iZNMW8Tm1U+c
bNEEyObSc0J7SP4+DKNTytnSeNe/mVqac9bCedHNrSyS0FsshKqvwFDt5Feql4Pv
Pwgv/iX/2Fhcz7pGuBgRB9UXLkX0zRYo4Ut61v7tnzgeGAu7Vg7tOQP1SWxBhbV7
wBVmtcaWI39POOX+y5ywClqrJFdtCq8VKORE+ARgEDtCql4kMmDc7a/M4a6SKNHE
/q3CY31gguRNNUqYupmKtmZYp4oztH5gP/5zxA/MxMyr4EGCwt9HsMdAI02+YNS5
Cv9hSJ0w1Plway3+4+f72eNo6hunhH+/6nrQc8yUGuh6yDJd1JPjrFOsEtiBM3FJ
rbe0DiRzMQLA63kTzEIg4/pMHYBONhvKCu0cKEwJd3hwHCcBkGcvPYaMAeULp2Hl
yQeEybd864sNpAx7maefJYyyBlOZbwgHXxfBcfXAK5rN+UX73DcYEPMFg2sX6/O0
la2MIdGTuNZcYgb6BB06IYMou7iqnI+JFc854v4aZNWY3vEmJTWgVhtjh+cDzpbc
ZEk5QR8XKKudEfu6xr8dP3M4iRJl7n7Ild6WWU49n7oNX8Dmf84ALEDyRKWWgIPa
0xwPDAsr8Etc7eVXplNgaIdy6EOYniA4LcAZnsOQWLMVwUTqNg6G10tM7pTPl1k2
AjNJ4zcquxqreZsJ06DQGHk9bRTeOfozNWAGHXARSB/iQEt2UIqzBGpeeT8LYqC6
i3TNGzTMSCgN+RP+4NDjYp925VWMEkO9LppJjBsQ9SK1ye07D6Vz378n0k4VvcAY
Qs7Zsb9pSygVXNdKA8ZoYInk3PR8lrBnPHi23eR0N52k2oAtivqvSL3gHifRJfdg
dPyhr+aqQvcDAeAjbSDi8OE4xx4wvTkBL2PR27On8FoqQ2MWBJscBOL+0xLf3WZr
FDNZD6W4iYP7f2w9OIaAburQLfGTVtzFcF23TtEmBKi+lO2hVN/ZzLb8Gzjc3aCl
FrMkxOKlk96fSrCyhGwACrerWiAIZZz5tvmmRqFGk30RJVipPi2DKM426v98Sqe5
1wnG8tunf5K3JCTGMeojnOJXJXfUJ0NeK1EJ+cxrNhdNNzqjrayulju6NTvEtlaP
Il2UJs19PhwZEqeCn3LVfdQhBqPy6WtF0iS07dDJhdUg39aiv9g4cjtU7OYvG/HM
qm7MsCwq3lhQtqtpf3UMbDKUZ2JQm94XmgYfwuRifwDU1o0fbS6zcFdzFPuzo3lb
4l/n7qZpEFo4K9eDSSMpjg/za3WE5BhKyPzNnVJy0YQdyeFh9XbvXfsmLANR7gXz
MGdYizgjuMDC8W/+5wQMAp1ZVhLNFaX5Vd39e82DDHrll8iJc+RAtdi/NSiSvy59
/u3EUw0EEBTAX4rFrWaWXagVvRw6SMKaA8HLM/YbjxL/Z7vt+sOiTxbEo6tkSlXf
bCPOHs6qlr3qCu4Ou9Jr3yx//NLCWYkhkgHZW1v1HS0+IIw+gfjBl6WPKTJmDVuh
qcshJ4NUDLhrPggtR9c0YhOAXJJVYgAdO0nR1NiTYFCMkKcapBAI0h/JtOqK3ZBT
AkCtajtJK8ophyigPud/R07KvuJAXBV3bCGcx9bKOSK7VC6Ks8sf3iS+ikrZWZ+s
iHXzxnImlKjY3WD0C7x+yCBJe1Dj7ZoAGIEM68KqJBhuJG7aXUZU1GDf8hImySIq
eBO5tCaC6bNB++byzTATXpXFK2WjmAjr1u7k3zOVEQpm/6sa2kwlL6hD2MsW8405
RazqQP8wDW6dOUx7bTqqsE2EjTOcRprw0PMxGFMPgLUocG/1YCWO4X+Jw1Qrxyec
Y+pYsZi+UHS4fF6GTGvJOLnjx63RXmDxqNqfjF8ATjFMG/3JW/tjo+lMcL9Vve70
0cXbGlHE2rvalrLqicBsVZh7EhpBeuvvXgGQ68d8iK53canWyeiCM+fCnQPB6jXY
vm04K/VJDRFZ/8gnT2/ZBEQA9GD4ifoI2xLMqZ3RPi9tmOvEIi6forIL7HbuHijG
lhDoee7dh1SSZmwXmTjwR6mayhsw8xxlO7y3eun/ZoRvtJ6ys6zwiVf0nPFW70Me
cYvuYDLgO5zsM7V1CORVYalSOVI5LUSkKL/Rff+YMdfayb5GPbsY2snzcofJ3fee
k5Zg8xkeeZEVfswC6FtcZoUhYCuJELIdNu4MKF5rkMcblf+S1ip8sqHFx/tib17J
zwtNJXgPKg297piBfB4ZpiEoRSFb8seFATo2QpMmybhFFGiQCBmIBAFJTIS09Tr5
yDBIRwjJJsMiaKyjOv4OZuUe84TU1uJrOu8v/1TUkHjOg3yhlJid9f2tQlFqYvtv
w6PT9k8rimJWJqz/0q1CvDfq605vSSPG68vj8jaL4Go0WmThZp55brnNuqTuqhiP
YGYVEOPNM0q+uKKqK4d3s03eoorzzb5APFhoYj5mDkpi1E9vAPIS/EKInV7e0KBB
L6DUmMhUTpiosX5bDZ4SdNyQjJj1j1wQaZOZ5UjsJlmvNewMZ828Ip7hMIRAS1lJ
2zCznXb0w7OgorliLVTLRYlGRr51qoVr+Ex5ZpIjsWjWX2oiDPDLyRfBW86tIfET
/CGjTU7JSraMvY2g4GBs0vBa09USuO0+/Mp3ixW1VrxZbBo07TX4YHXRB2gSC8zB
/txQ9dEMleVu1gAzJ0Sfwu81DKhXX7hC6umFPNPD1n8JG4VUolr0jdiUHsX0YaeX
7itGBSE+x8hgrmGKO3En1OjaA1XLyKPSkrpd8nkRSeSfk7ReXOCz3dZ/LKkvgBCE
Gtbys9ycTKUQkq6BK7x+g3zEYlkm5Y6gBQLMVNdT988rVMtNU57tprt3dRuHX30g
6XZtCx7ssqUHzZuxQS5OGQD7wbXTXfXajBX0Y4K/lk+kNCofYhQEu4SAd4Y9jI2e
uGpQCPEGBAMQttFyPGwzk3FU5lyAaGbILn+347ih51aj/AxXzYJkPUgP/lDxAgca
O1qvWDvYoVR5qScftMm9VOtKWcZoRyff5UjybnFTUM8hDufrdw8t9NBDU527FQVf
wgQFOAGMKYlgjMze2PFtzBeYLRd7Z9KBVvtYL4AON3rbT8NU2ICzi73KwoEyF2H0
johMkw2YjiecitXrkNutj/gZ7olSYC4UwaCk8X4K0t1I5ojiq1GpURICye8CUOx3
xVH1ja+eINzEC+my/V50b8sHtRBdJlRm5ilOz0CZ/3l2FaDhmqOP9i35fsIj3pid
3XzPeF2NmzbJwgaDLP87Zm5Uul7NOg4gd4nl5e21XrSlsSEVwpYV8qe4MekhcFa1
eeAJ2cqkcD2E7trLngbfEkumA4Q6KyujEjhbP7uHzSwF72UpsHBOJ/PI35VcfNkj
+KAmwY5Pr/cN1eVP6MCH+7aT3NrTiFBVbuVpvDYlAQdZpGXVgQ1qdNDRFz7cciuu
R7Mf0YJ01OzFdBzc8k0j523UYtCsZ3I5yFvzqNJ0UlqudNrJ0bBUWIuLCetgcKsS
2yTe+q8gW6fhTMHYL4KO2qxAQiHCDh+NVZGpjN6gLRAVM6LwEqVSeIaUPnqzO4dx
STLPm1oTNLXkAwXSvfmnMmQhB1Lasz++p4zUl2bPNU/eCoIBvTJlfMeODn3pWFsM
lmZgpsQkuVQ6dwJTWLKcPbiES2qqzRZTpB9qRlpdO+QlWlCYQwA7+57o9nf1LGlc
ja7LpoEVsY2W3DKAo2bQZBf4CTwqmgrorjvti/KZkMMPgDBSIV4jLemHv0XiJFDe
cypIIf/+uIPNdjUi54sFhiv+fjBxGbqZ2i5XFFzSV4rRPO0kGqgxfXvEowYkYCiZ
HLV3ziupTZ8QQxC/BNe1jRhhkeJhLvIPN6dc41AgOADIia+TIg0JXJf89T8gdo0v
LL7Vym/+CiLd5UY0rd9D8DpnsEC1aliAZv1gTgSp5zxaABYczXIv5EZGh1yhAryv
48fuLwwGIEX5YcL4haXN1bXmL2wx+jVZNqizjN7fxobY8u1lKzudn3V3yuwLXqPn
pPTNlvsMrcWqDJKV19SDMmHuFMyw0ZXW4v8Wtr7SlSnNWlT3GEo5nICvtnXTE/gB
e+FSbIphnXTwDJm2FdPh1uiQbmX9XjrQwnlvoFFccRanFgxujlOI5W2djsp1DRXh
5FkSumb1NPcjBXRWM0K+2RtmPzbFCeBKUgP24tbnZXrg1BSyYoUsCyHKggdt88pA
kuu2uSK0WNDthwMycL9KbGXOQ+Q3bdleWhB/H70IK6CRi+oiZ7niPD0GZLWaAOIu
2bjC6+wB+VI/zJySp4ymtF8FBkDlPWsu9VsBZZ3ficbBERHypLAXeEiipvGGCsL1
oH2LF4T/wzRuhK6rlvgtDA+HP8EY6TWKMmaWfWOTnARcO6GxJdlf5PDt8uySjzi8
cGM4CDIUoU/n8VIJEAr8hOMqcbPKzI5eB/zuK+66RTCgTI0UIp+/bPXicx5B1bQW
I1b1bRtqve3E+maPSrAqvvSAq08OjgA/nm0kPFoNln1EihjrQXBsuz6GiSbta/My
IbwmFgDJd2Wnqn/ePMlTCvyz7CoJUWuqU65/l9wFsRyATvAw5zHc+eKeMs1kH28B
hMEjWCGERBSsNiGcuRkeylRAfQmRDt5g1uQ6rp6VBkD/L7VFSOWGZmtAUxu+sikd
ltbSxbk+qePernIGKPFe/YA6qSkbvfm3/3uwfXCdQUBIYwCVbDUCOoiS+9jAlWPI
opf8IWuIaAz1hj3cgu+/XznkYlnARG4En9BBMN9/1brhmtNHZB4sCiHxQyyfBBxH
iew089rPKCBB3UrVLac5xEwFLXw0XitPGy/W4qCGi0OXKkEpBpbDRccs8McMu/MA
wmT+USZCZVJm3/rkc19ekKWkmCQeX6vGY++Q3YNhNhcL9ctM/ZpStzRqf/lL0c7R
H38K80jSaAxA+PpJksNww5s17ITa16J/fipQffwoiLva68fZgu4L5Y4ASJsnbYSh
rgmGgIv5S8csTJ6+a2yvtRWSzEp00vxQbafbm1yPKSBb1myWLTo8RGpx95NUiQ4p
GYJdfjPq1HU9P2t8eV0hfIo7znyicLBUYLy3+9Qrv9aZAK3irAM54oaK7AGgtS6t
tYxzwm0N0qbtoaV23oTBjnAVxlCvIPmqhBot5X2l3Sn2xNNMMXNsxJBIfksiwTM5
o3G4l9UjY7XUjiuWA+J0w/S+qLXt2ef5fV/GtNaQjqsJI5GyxDRFDUT3DManJ5uc
rJ4LNqVWKMPlepLoD/x2v5NUBj4+dBIgcw5wAG0RiOnbHnuS+2tDXY9uEvxTu2p+
q64uva1x4DLV2UjYSuGt5JGwHaOB0a87YC4qnWvFLoyWL62+dz2TkxpurJg8mUC+
qx5TM/FgXyGXUftgnYiDKNCSwIHTLLI58wQ+VhT+/SLstdN1kt0KAMXsCUSyiC91
OlrI3htRYjJP/nBLSHuu8fLuDD6aFmVj6huPS1kAL/SmOLsBh7CaVt3EYxkmOggJ
nugr2aU/uPgjbmCKm9dDkHhVXRmmayPveYvSltTocndRK58bGYRLdhMlubEyi/Vn
X52jCduHjUw0X+PSg3hH2vlS0Nn6IFc7csjYefTvouibL0umUtYL99ngTBHEgSEt
z7J+4amAPd9aqY+BQc5NVMJINOUlnH5UDWSfYLGgEpuL9baG+St9Sbl//G18GP9C
zwcnHxMwvSV6Z9kedG+cLKIv3BqGcku23S/uXU0s+shdgGBWgaqBxgLcFQV+vWPd
P4/jGsAPmI8zxhh/GbEFqN8KSMBRCbfF5hlpRCCUrGS6A+pydfGiR8l/TekleFES
ToJCFbyPptK0p9UhvmKlFkKl38uMbEKV5yuTIJ4JrRFUvs7DH0dEjBeQNUBuxLw2
RRklMac/vS2XN8buf1Hq565PxjCQy1UDdh6h3nSHB8VCY1oVyVBN8C+sCuBTCizN
sz+lqHGYxziGlIGwsE8YMpYkpq+TbedSb2ZnCNiZymuwm4j/5mX9wqlXzyx6Jc9y
1XGURv132aa+u0EjNt5s28AxQClxmo1ZTqLNnqwwo3+Ir5/DU2lmksDTnAGvAccg
8pCDuF9QJa1UMZi0SRdIlDCe3U9qCW1U4RD7isNyaEJrV/Kgy1YyB4NKzzq46cpe
ZLGZgi+1+Gd9a8KTT16OyjpqCDI+DIITpqlGaxayA2s/4w1yZhDS2lpcmDJxxuGZ
lyOzvwHuN5niIYbSTofC+s+SiKbnjkUaPyPoA54b0TznCM/ztC46d3Rg6RMZL4hK
kcm3aGpabPfe48Wld1zhOx0VFyvMTW7l6I9BXBc08GeL7LIWmf9E/91oW+knV7VM
wnWTGg3zxCjKTDf3FbPUstyMgCl28u6a7ieBazG4LqH8f54TJTIBjYkG93FjlYrB
YNX4eSbdxca/6UDj/ELOt3FI7bxfsDsniQlZXhOSjGlOaKIFt0M+cSF0UDtdG1N8
R+9sdHEWZvYXOa3YRWdFTOXPMg77ijIVPN/rU6pi6Vsi8ynSlNJXsE64sWvooGdm
9DcITymp89VHIgVvvqAM5FxGxGnX79jRiCZ+DrZhbAFFwoYLMDs4IBdhxLAA9lfg
7f6vWEqIUe5MtedvzhS+2iOXihxuwhSUgSuo9VnCm3HgZQnasxa8BH80hcDB6QPS
dQW4BYPFe8bi8lsvR/Gp6Jf39uCt0rEhgiw9WiWYlZRLva8QPcdL2hFh4RyRdKkB
sc/XkSRO22rI5i2aItqVJdwGVTrFFFWQfPr/xHCcVGIpw/cbMyVAKqNSOywEBQcu
cQxddcRhrOWnAi0/An+cvoGyF2Aej+Dfor756eFPEESdxHKUoBGotTMCZ7q/UDZc
C1ErbFBVdyL9faDEmKy3qgs5voD6ZlmIrzoOC13zu3RtmhZ+b9xi+5mGxFQnP0B1
+zzVjfR81dTA/ekixNtjmxWkLhU7srnRmckxOOT+KMbJg55jI5/B9cgT+aWXD3lR
5QHAuold+Z+1Ss71JlPwq587nLpFqfaD67zSkhGFBaABt5+8Ue/m6GZQZRBKxkcY
B+UM3sZFibPTyT6zabXsGhGWFgE2XmS6SSzluUEP3b5FCKDZXtBj8j6gDGET8ubH
EOrdo2zhshxaLGo+8/RjZXd7aAktPzjX89N0A3Uao+ea3ullhyeKTf7mzxYboNBF
JZTYqxm+joop8SPzq1jgEnK+IjxQWbrzHEb8NGOTN71w7goscC42CzBPib6sf6Lr
1Yx21VUkDpZFsIvXPU/ydDATXOGmG9ZtbLJkV8BsSX/KKvAcM21hNEUqncyjEG3J
Cni7PfkXMpmXnbMu/pd7nQZJ7qgnHUkRJ0fvX3I1/0Ia6KYdccMwsAyEvGXszfzu
fr/VjwRC7A+AORdaOzqD3OgJyPLymPfB4PVTjeBEcgDz+5lADdIAQMgD5z5FhHzU
EizNDJdoNcGaIwowL5LFEFLgXgTbwZudYNH3+jGcyOdzdq+n7jSD5kPB/R2dye8z
LTWXAAyP1s8yggTHsjFauqv+sHeX9oz03RpsxpzXZ7MCZCa5IA9xuoEUWvgBRZ/1
GxKfl1Z6L0ZjzsFicYS7szCwc1fdoX5fX9Yx7nwUiffqQ42zd7xV2pGRdZqaXDkG
X8TvnYUyd9tfqRvd4shMTCgXvnFLFg9wWhc33QYVjCSm/Ps36lrciIUwREOvwofC
/qcIeCKi1KuIBanPe8akTNZwY+Lds8g99A+sDzw+Zms/YD2PjOBw5tB9X4ZqogV9
ZK+AKYWVOMmzSsMBJEAEmTTLYZeE8jmxrrsCqiOwDd6YeS6j11jY1o1721UJIvkL
VC/RcxsQV72DuYf7MJEN8gdac5p6wuujBnjldndwbtPZUawQ6+TGM6i+TV6dEoOI
6hu6oDwoxn5YxWqpwZrPKOw5rDN7wL3dTKsZVMUkDDNtgpW1O9OYW3bCr+/55c3M
nfcnHOkQzOQmmaAd0eA0DEss6u2f8gZ0XOZGgXm2xkioNE6z76kg+vc+lyyxuhXd
kwsLI/ckRf9Li2nwsidqTRCZagm8Si4HPxQf2CIVwWV87BYVhjewVuy0sJSMAxKG
HI9lZGtsMSWwgra/Dk8bFlZyB9jDkKVsbi6raangRTUs0XWngQ/bl4kqrig72hCO
uaMsslu3JKzpay3wm4NG97d+UhC0mJFTPsS+GDFTVORf2F7fCUs4rqFaWob+n73B
s5iPXc1Ip0fCaM3KTsAKuD/r4QnFV10fPrWBb2rjcho43TPfO9+U+M32VRzJH3ig
yXuF2QGNqyDaTBVlGIgWfAmtbs0pS6HhidqlDtbqXSPeybWfHSrEps1M3jMYEU9I
f+cT2zDrE/SgT+suOd1jOrawOKWe8cCgmxYaE83H+PDwaguel1MBaL/AdeLvEmmG
gu6hLOjUhUuaZ3TCZ0p6Hg/q4BPmnYUzurHQTnfilb1iBVdZlZYXY8t19Ji0qm7E
NIqkdr4R4Ce7RkZvzbT+9tdkGvm6KuD1s1oNDgu12TaP0Gc8LPySgFOhl78xyzor
My0J6LTUZ1tUjR0AoEupMYIxqlsgtSB5RKkTJZCvOUCVuHmuQl1pWVUx+kXpyxBD
8PtfKkH2NRjXAD4/eFnA8G24WOYR1OegTGKXfhWcSr2Im8Ny4fPS+ZRkj3alrhWo
p1I67fS7B9JVqJ+GHEGf0jYsNZPDKJaYxvgfI+N9TW/LxHdtOEgRjLbSdOz7ypWW
2VS0CnhHgBFCBczrbbBH1s0GPTOowHx1fFLQTabM3mvNFe7BMD1bhoK7mWbxkPy0
n9kxekUa48d2IK4A0JQjcACFKanqRe0MWJIRdfTrnzW47HZzI/dbM4AwADdemJCN
QfYvXGd7X10/f5WksYsxf+LnD6S1VWfZ13AM1BAQVQiO6OurwPukvbSfAa26ETit
PMY+bQlnnESLa5wwkZaMwwka+1sMBwhtYX/M7fAZi+1RKLXXMHePGK544fHO8lvB
zL5+3B7NS4Rvw3Bx5dfBbKcuO8AuDXCbc9L4cpSYMNUaOi8BvtKigKnuQ7iugMX0
iOb7fOpGP4xNem6LikSOcmN4ZknErHPf/ak2V7qMlJ8uT0f5EFwMZWGb9QxxuJcU
NKJ+ZAV5pqPB6dAqEY1I6Mdr3YS/vvyp6bYW2fOadHKCYJshPOFSs8RT/119LEMY
+PORnR7VrKCjVpdzU8G/rqUYnVWunx8DQ0HDh3tCpFs9Eo6WwYM0AmcVFJc6fFNU
Ptw7SKK+/Iu/o0DR29EnoQ3IMnAKzYhRfTCR7qW1OXltU7vAFNq1Tzp6f4FXM5H1
wouQC/E/rVY13nLmfinARFPTmjpEmWOxtq47IU7DMclRBhvJCCMcQwmdiBgx8yoj
HUCULU2IZMubx2wvs4+S6FuCldcugIQQ97c8/eAJz1tJBPOK2XKttk+ly97+ZtY+
w2EVJc9MjhL1eLP46NhB5ZY7sc6xNu9t8Nyh+P4OUrRNO7EIA7sDan7kY7nvSFRs
MliIYv4hWXBnNM3zTc4aDB4zIdCgf+F6lkP9B9BqpSggB7HNOFzoG8PPPB85pXYX
+EvBw/XHZ1V0H32pZ6qaB+rFCh/O5dIy8hy8a2JLsbdTzJbJ/xvJJDzOAwWCcVBf
bvz3aZsXbY9ckTPBeq3Wv5/C3uThivu2SuwwP42Tp5QLPh4m2J0GEz6Wj8E3OL53
0ZHdljhAVo6Ox1vQXq4wR5BYaidqJxZoAkdreV0LGyeSyBvzyh8Ou0Pn8aMxgYI1
38D7Onu4werzS1REJRcQEbwFkJ6l6Y5duYcadg1zqMb59/7ZjCR1qaimrGz7c/V6
SVtHctqBFswD24YYV20Fj2DEcgauqGPtqqaMzACXeDgf1zn02xT2nl/ATMVKRSzm
U8AC6OfAEx/7yr+UvlMTDvmqQdYxLd2CRsohKbLSqJlLa/f6DrPllu6CM8ZTYw6T
uG1DoYRdGWdMrYjFKWWA0j4OdS1BGDYqbZ+DNQqicTxZDmCgrfBm0QpV2nWzX7Lt
ewY1srd1lEwQqOdYv4msTG32mGPJb2b9n0a1xqSzB45JnSf+9kO31uVr7aBZlTrA
qO/TfSBeerSDttl2pfucIupgCk1xpXTbVkIl36xRdY/m5CoyOCIGzgS3tQUNrqgz
p/KxKpF7TEmM4Hp+XhHCdLOO/Ba7bnmENXrh2SLKuvp4OhmwJqUX+EyesxNMJzcz
YO/KnRsqdAGKxG2ZnFsfCOL+CtgIrBP3GNPadwcJsMUJHoYPmlznfgiOA95jAb0z
Iohvc78cFXLs1JUQeuJjiutgysAKE/1zGqUnWz7xelj1xH9N9m0ow3l1IXW6Ai3C
XscBnnCGxY3TpYV28PXQHEM+d1pbzkac6mujV/NKvO9yfWNw5nHKBB5c+A1mNauq
HJ+U+DOE1W7DmVfYStwTJQEICs3UKEbhaWDznJXRlkwwsI4zbFbo6Xj6AhNwXqne
nfL22XX/AuTCk/vq2ynIKzVWjnRDop0N7Se5C3bcLWXKVt677FjzlfXyw8JAzGHK
6f4gDhbKFZ4Q5n88JAneeaWonToMVzehPt0Ou2Yt8BfIlWJtO+tsCPmxCU2v7hPw
b1uwinEMO4C3lLjs72ouTjM1XleOTbaWGuIBsSu+M1lgjri1Ht5MSpNL5WZxw06P
INL5L3JIwpP48WKtE1ixX4Mak/QOPQKcvlJJO3uRjkqXN3yBVJ7dlVbY/bE0fgT/
U7h18kRxtLBl+U5iEVcuCJUHMVJxtQa0tvx+vpd2S1q0yt5iKSO4RYf4SKXjxR15
Pi2CfVmrFYv3kZbgnjJx7BziiKYio7NgZgpDYsKj8TuBztLi4yHzm/PivIG1zuSb
OG8wUv5SnPJtMkm/Mm6i2IXItZndHM7STyh8aDqyp8Ctleijqr9VEdA/ejDrXh5x
G3NwJLgbcedk9F5dJyDm4ydgb7aGAXWv+C272lXyzc+Bc6y71AY5j0ZnWTrs5xDS
DnRt352aya2SvqKmiPNQ96IxOCNcpYly9c6Pbs/HYcrW/HeWTha6cEMkolkUdtrY
5vcHHKRco8Hj8BEWIzF8wfWD4NZDBZ17za1zYxVPpE/EGutU8UDjVUcR44A4bKH2
MBo3BpN96OvtVEVm+W2xpJyR0jYbVZT4M1N307xxA+JqNCdkC4BpNWtt8X4J2fwr
3dmD8HCJ7PVw/URyNx+38r7jFyVjRH07IeExKqnlnvWjecO66YK/h8a1gj9YcFJU
7DRzOhQzpsucKzqDI0qxfMXTDsK1jxRkbl4CbwcRUFVLj6+hAcjTXxirxcKQGSdB
Jh3d0gy/6LNdflas17bC0MfLfZlAyTVvD+0O5oSbJaAFtTuMW0wRBqI4QXbrm0ep
pCmIFyC3usMYDDQTJDKLnyDd3xaKrsk64Eg1zdp49dKdMhREEeoaME9DyJ2EScLa
9+FFTySHePXLKsoK/vZGD2FUm9xEUss2S+YMPoH8mQZt6QT3ZNxMIkcnPKSy3TON
H7iNTIGbDUxXjD7t3oCzGkCu/JjY6WZ9/VmvdizuYHshP/MQc2wqyPRatot5T7xr
K0QdV1mqlFRVgnBGH/fAWt67xj55LGGWF0IEd768yGzps29qQkz4EmOMoXlmujUA
oQMDppb/sK57h18co5+XWmA5RIjV4ObPY6r7e1wQGTDtYWpxiRZvMypSBcGFum16
Sfc4+aA5IjTBA1wQ8/tDBl3SrGQ01/sodxTPpb7RZ9zM56BXGQ0DXN5BK+NbEoPU
KhDSbEOtUI2Go8i6COum3ckZvwsmIwUpRJKzXbgNE9rjgN+OoTALNy4TP6+KBqSV
HDdR9S6PV7JBDohGPRn3vLP8f6sjoph9gJEN+oi/1bB6dw8Vtn2mlpGwp9IHsAbz
Tqrw4i+U76wozAAHljL8/sfND2uOQoWg4K9Nq4DgdTKtQ/Y08aOeN9nsHw6QTwNM
l81ok9CzGuoOUo8jFqkmrNTta/+cjyDNSjikap5zdcNX9wp9Y4SRJ/+nj+myXXfo
ykeUGi9sMvOvrQTrpRd/GgykqD7mvRsjwLTQ2Ai0TdnETbu/M0s4sJ26gzGlu/w+
ihGqM4irlXTMZhx6cVmwP2j567Yavl34YDy+7IPFUIv2Ou2rkDpgVJYk7FHvT8dq
z3eWKOvG7ZYSl31jyKdSn1kcziYl+4JA2j7fiQGVbT1Hwu8Of/froLyHSl/qhS2t
/XETZqKCrU0d6JCQ6wM9Hm5nvm9u3/deNZhsKJ5B8jxas+D3Qp9A6ciYN3ed4sSg
ijxgVG9CC0tuHeT7Izp1TEviQrYFPUlP6u+ZqgWdU49/sq+xZPkygbTNyc3N5tbP
eQF1J7GVVL3WuFzEwiRCcc+lrpeEDLPnjjNl/9BK7t4KVQRpBwHp6tOLaj8m7WcY
bJbhS6FVmhhxcbka7My32gpzJarSoM/jTyNvB0yNjjWErsjqGvOuMDfSzRJeHqvk
89gCi3toHJpnjcWHn1JnZGDF0s7r/t0ZNszz0zTbuYkc9H2v8fol6ZCVhaqPEkLm
Nq5FXIz56QFTN1mjxFfKPUEd6mNHTe+WIfg6KStp/0CMHpafM2F/y1Ai48rs33Ld
88D0AcCbQhR8Z6fgQ1a8ZUU4QenBcBM4ETL48GwGXtKQR/OnJ4EV0W5tTVVVTGoV
I6vyT5Ba8dZzKQe+Ud3LMC88bjgdzE5e10XiObrmuftmXDO0OtS8BpbH1j08q6TO
iTc8vDK1jxVLvGn/q9pxe0thsqQkCsVxLLA3LBl5DELoVdPyJI1u7Y7Ams2112Ea
x7S8LqF7Xl9DjzPlEBta4ky6cuavEUBDYlDi2LYTtg5hmiYVY+2bZWLMokEo82Qr
Zef2pwBtZIxW8q5vOhQVoKMN3SK2wUpu3Iv5UzwSnn4TEZAhDSrx0mTTlLrlK/EX
TAA+1p11BEjdD1S2DGVM8MJnZqTMsGzWhxRB6U4gClp+Ls3ulpV6ecBxfYAxxMRu
OGE2sAxNPr6cBzI4vIwMZl4AZzNuhjad5Rvy3QYyD5NEUKC7U2Kow4nrlwl3nHls
woTfkkFCyV4lTUVd8NNZ7sFkQknJxZi54wZOBLex84LjFQZ/6nKIZHszItj2cC2H
/IaDNdtA1lg0f8I2rxLmp6NPVtyogu3PPL1mhNRsJt7A6fz7JgQ1PzoVtyFx3obb
OzNN+pyW6udKeTViTr1h3jr9dtDG7cXfVFnttfiBnEY+uz15NoQ9kTCUxjiO0/Zi
bv8HtocV7LJU+Qsw5JaAODmzg0KsHpjBPqGlV7LOOCYRWtZJBiOUOOuX6NkjNRXY
wVZ+ko4KmrJScXZxYGWnticOehkxZ7vZkNSFqoEb0OCgEfMykIjLwFmTMWDeaJKv
8Dq70Y9X2oKPcdL/1xAzOkh4ZANA/c8FzKuA+WzLo+TzHmFClQfkaHwK4rqYTlhn
E6Homqn0hjzM5GECFZ8aDOzeAWmmI92Zh77fDmVf64GYNhARURMFpdlDgEX3tGqY
HQAkjZnt98d4Jlz6pMGquICkSugjDi1UJdJmJodiMk+GPMH/qGl0fzZ6sifQj3Km
JjBoXkaxQo88SVSqAsN8QIzVKAxsrEvJeMWbnc8G9NXUBSlO3Uu84AngTOM5SYcA
yqnDt1jsuThBVahmjML+SGDTKHg7VhNqDVK64aC/PH2wDRje1oPkEFIqeMJ3Mkne
3UpllelpELP52p5xv0aZiF40b/F5nHj9+enl3WzjG7vmHKz32eaQyc12fhnkSGUY
fIoe1saDi9DHaNQLEU5XFiN7H6aR3xKV95DYrNMCGlVNnxglbNoMrd2zoTXPEQOK
3olkk+Mf5XEw4mLzH72OX/gCW9FYJeBVMaUtVLGpz6GTyreCa+DISDFHV7yT8S4Q
/5ks/V3GyJaLSKBcZtOwrJxClz8ULQojCzWnnxcZ88bJAkNHZyJQj8zI7DKy8JdZ
+zZJq9Z2KRunxfAMWeevuxVTMRhaTLf0DHTirt1c1W8DGpTURb1itPmytAmTkXRc
1lb/Yr9w401NrrdFz+zD521XTcKrVPtLPYw9pYALU2f4hp4HeXaDYgnWM9T7lMBO
yU/xBC2iGxWwpTDiGGIgOGbaH218jZYdWXpGsJbzj7ptqKyd0TYQXM44dZshtDjK
SBNS9cNM2+1DI2L/pBuKYVNN+CuF82HLomhra2N7N5dwxxU6qh8RWdaG8G5Yc6Jv
HzqMcBB9R9v7rHiegcxFgm4jJg8RQL30zOzVSbhdfDD/0lvuEnaR/bYS8mQWvUQc
kTtXUNKKqxY9nJzgy6rIl0AMvnylXo1wGVUjMVkaqhRWwbVZuS4vrya2sIbXYfe7
o57q2bhfS+QNOgdIgfIXFXHEuQtEnAkA3LDAXmYS9XhVG0eJGOjLCw3JjlLHJ4m7
0CV+JcZHc05TxymWI5ybbr5M/uAySLkyGUK2crziwgHXClGQC66B11gFxS8m+ni4
CjpR6alaCm4+heIfEXd4eE0dr86BsfnHEMX0NvA68ovAbxg3ZLtnnJUT2feF4jl7
LqSdY1UheOPtE92RaAZMUeK0qip4WytXuNi/WPohXB21FT9d4almGcm5j4mxRUjJ
EI3zt48vFURZWAaxHuA0uzQuD0LmngueDM5RUZMit2iVfmsxI2iWYMRRXoB3sQRf
Dr8dhGqgNDwKvjv7jW4at9qbPyZ9LqS3a+YtmZx7DZLWNYeNRP5VhNWheNgmpNVw
/0imng28SvwzntPRjiI6JxUwSCmwOYkwZHhS1A2WAEQC7kr4KJXBnY8Fd+KR1T7N
Zoh0uPZ5E9dOryMzyLuTcYSajEJXufbH/rHeu+jyH0Ztx2YuGvjzPfZ06VwT/CFW
c1ajKlap0t652n4r9tNwFIxhSjJa9ckordTLz8J0WQw0bHI+Z/kUKrihtGjSJ20I
aAKbKoKQYJT1hl9dHvaQKKa4SkICY8NaUHm2w1q2QYh/WB6dAjDmXgTdMkwhWGHB
IiJABks773xh/LgTt6Onhu/7q4vSKwwtUj+RI6u+4alRw9qx1S1/e8qADJF0V/c9
7SQ0a7Dz8yxjnGb81whC6OfWUq6Au+YnvqAxNjpQ28SD5z7JjzIaZ2izPGUon8al
sPPLEe8ojHqIaK4Kposak8J5pZnWUYzNFgAdcuh7+iMMG0P60dDfPYNWmskpkS06
AaRJUGISQvwdJys4wmZvBPp7wEjVHn7FxS6NKpoHBWGxlPuZvMComWhoevj5pwHI
59sAMP9OXLIn2/kTtuuJAg989F6fhnKRQ7Lf1g/C2SGhTvJRZ3dQOT+/SuAXPDhU
mYoPy0yLUil7aCQy75A62MrMZ8F3xW2MOcWB5hqgYqFoSEdUp0/zQNYPvM5TSqHv
QsSZ7g42psHsLOHCqTH34zb6iPWLcHsoj3gHPUx2fYRMPeg4AsXbLJrb90DX9YXs
xZ1VdkTeWoe6sLzQc3IzQJjg3ql0OEEdmau6hj3Enka7u49W0lhfhGX+RbQZbCEc
ZaOl0II1Mh+KJi14Ptnum8ENTCzt4V1wgT5GSyBGLtwTbYfsJvSJWC4ax6H9tcmA
Iydqrd997BzbxboVP3psp6Fuvtjz24mecHMA9Lcf6ZAKXrKDShOfz9nhp3kT+P7E
Cs5MWznKoGSWr+PfbkGU1yaxnc9PzRDMteYF69miX3mnRJ22+/HKLYH3YWuyFALP
p8XdLEIa+aSr6k0bhGzZJF/hSevjo5X+ewlJ3WJ46T7OJZOkOHawltvUCdVNGGxP
VRxOImlW8/NbPFJOqU6lajqs4xdsp+w5ajrNGtGoEi/BUNTVl2bhIjulmuarv0hy
hOLT5lrJGziVgq3nLTBij44+Vaa9BKU00PsrRqlOk5Fm9tKtGKOjSz8Lm1NPB4Hv
vbfBynEemQQaJwxRIvG8akQ1JpL/L2L8/uFMbN3bpc08sBYBO3cfkWcNXtTKn9nO
qZhAZh+n2isWuvOSqfnQkpr02BPF0VLZsTiubW1fAnfx6Nhn/RyPKf+IAZjvRux/
keJ2YRbPDjIJW6N05X8BQuDosL2ETJcKIC1EhG5jF3idGKfw+/6rPK5D6jO01j8H
C8RH4bI16DRQKxz0PF4S7FJlKZRlUY1eW8czfs1i3XTwI9BuF8/frvJPgxMMVBwZ
ZMB49A5cte7HWh+xllwy4w3XYsx/q7RLAgW/9uGVkidfO1UK3Cw4kppETZCJ83YC
GHfH/4Wlt1m1c5HQP1h0wL3KMItcJwr811B5ZzNI/+SFQWW726QAO63uaN07/H1z
x5SBEFtlNfzu6AFQBHkuYq05UBl4hqqgpAWttZmDRfnRno3Mn+jPTIgv95SU4tdU
YixzWXNL3yVcyJKlFONGRWot1wtIb9C5RWUWTDgmC7Mmg2MLcx+j/ERtNKXA7oz4
JpmS2sh+Mhoalp08oB6rEUshO58GxwX8YYXslZGdlDGv8v7OEhyitM2Qp8X7MVLs
wunm2uXQ4wGBLHi5KYoKf72WNknFsqGaIOJyGtLF5PJ8RTYjofDdEnX+kxLcfud6
5mW8y6vv9OaeuCzqUHb2kb/BMBeL8HaOP5NzT3YcjgSA+A13OD7r2ad/0eACGo+F
xVnTcSG062ofE80LjghRV2OvXt7GU4SnVckNYFl0tj7F1y7oCmqNW9lSZiQf4bB7
/1LfjlmT3l+YUOO+R5e3KEtWPVW+M9hlNI+oKZivEVSzIXD9IFNOzymynK5B7KNS
M9BoHsfWGdYQ+s1+TRA5XcrEtmF86fO/qE/OivBKY4RcUhtJGtOMbm8jrq3QB3mP
/7M7yCseba4NE8mag1NNf+LIq4rtjkiJUCkaPn1WFs81p2kA/o8nSboRI+n7tyeC
e/iUeqbShwPH0PJBINdrx6jtY74X3aIXkK5gR+vPv3ayGwLjL7ZkzH59aP1PnYIR
oEatqv7sgH7q2yCA4WAMdM1MV2QCSh9uutdCo9AxLNLAIpWsA/7R4A/t5jd6bvm3
3I7l3dKFEIJt5Z0FXW350ahMIP4tGCEgD7Z9AqDWHnZuakJg9xwOOkUrrhCpOQ+L
6twIIZHbBj/p24W1rzq2EcIxJtS/1VRA5Hz8yMVC6R4H9AswLW2O+MZGzciD0knG
Zbj13oztEaVNvOwutBXcc+U+dxf2pGip0NkHVTRU7miYgpPkhnV0Pdc1ogAWS68k
mqqwgoATo50WpjpzuozMeDaBeDj6eljDcvWyPU+S7OSif8XeBxSToHFUOGYmv7pB
+uHk+i29HlxzGAbXCwjH7nh5G6zaIEXxdTXWiHuIVqSCF9QsPunWlABwV7sC00iv
SxxUDqy1WWiM20UtvZoAXm8lKNNpuMcw4YpOq6ICymsFlaFvS1s21UUnBS9hjeme
9RwIfUA6C/EgNiuZS2Xv41kaeX9Lkf1ZW3GGgns2hI7Eit1UhNMPmvtgOBD0nv8t
b6/ypP3ttj9j+Y41sEgZZoZTWo3PSeR/kONRkVNVxKnjATXyq3UYKf2cqGiAqerI
X72PDi54Gmjm1lE7k5P3ScuZruf+Kp38w0cCOLdtlEIUEScptYNWgCjelot/Evux
HNZKVTf/rJ6bTsDj/82Yc5/d4+9P8daN3GMC3ufOG+CV5eR/THdKzwCmVMC7w/nh
hydUdxkUwwe0wka+EY4q0kvnlECe5bLAp5qKZwKxUKIx9N1AmCo634P1wFm5lVJJ
cg7xnXWjxWdGQ/acjC4Vu4Mt72nJVAA26QKSIOQbxRYzOwMibuVlqaxz81yLvZAW
uvEcHPfa5C9D0I5j0PBp+mtmHifg05qcTYrb4MpUeu2pNZ4LSoWeJRKkVXZX223o
ZeoN34IEg/PY1j76Jtf4bRbm7q2eyJa3AF3LEDkS9fO0uZuMbtAbO7CQME5hcxSD
uFsohtfosRSfxrHhwesTdhgeiHK0hcEQnLbo5AGr1zU6vIhZl4p18hil1+UqvRNi
c4q5OgEmB0rFrqsAt++sjr8Bpodvg71qyuxInYWEXH78YbdGPOa1tUEfR6waPKpr
mOtjR8Y/R8s29UK0RfSfrm+7y0CNN0wo63lyojHIn2sJP+h0HKn9X5MojJ5mTvYO
qKHpkenkxznb3FeiZrlYE+OcYApVNP/FZA+GnlpfHw03iB6SgNnDXgr/efCSS9YZ
JWcrmt7B+fPSnwUZd8LqWE9T7EB5n35vXNFrzjMC9GE8DOuIaReHvt/lVGs1bJEW
KUCRW4vv0kxCPD43uRDl0FYHjjEc2tdhPnFq/diUuTeeCyo6o9Ai/qe5qXGqDcb1
SWSSCeqgesB5R2k2gPaJHzJguadn+QchZVzA+DO4nw6bghISOYFdLkxKEhbuD/13
mMryUK2FgtKSS9SD8cO2gOUWbvaQm3qWhiVW+NGZ24krmpXXcrnirk4S8zOJZMhc
PmlvvGkKkJKSLYpGLWViSlAlh/UnQX7hOWEcyVIlC1SqffeXgaXXzzxcIQAW7eY/
tJZjovVcUM0c9pfXIhOPHdEGjJPdRot9WCfi3YIufDAyyAay1+LXHs6auB3OZMYj
oTgw2ukoFSHqJwsogj+b+eFV++T5kkhQfwQ4EUgZhi86KDxgDwberksvvFUbvcct
kHc2qSMcbFTU2RwDX9ghGZFLE3FnqByvGf0lJOq7/2/VMtKJa0DkXnIJlZAB9YTh
kHKwqAmCKgEEM7op4lnSCxNnyVdHT0zc4OnY36ftx3DfLnxfXUTaNiAUiqaH9khT
tC0312bx6aRMEauSSH3zdR2a4EftxB2A7Q08zwcCoxUCqRxmR8oJSuj3Eh74qJ9G
yN/E5yYL8ygKhgyB3pHuhBsirET+ge1bVw8ZFrCUfByvaEfT8415YdtY35tc4ikC
a5d9QqTOoopzwMBb9v64fhK8xlNVbVGn4+diT7eN3hqwS05GtAfB8yNilnTnYj4D
+YmhTiPJYBh3asRlblm/Gi4z4Bu5sOs+LOKRfnMWaVoOuXk7PGCcBwThi/r7RHBG
svAf7VsdysGfPbWz28x4f8v1Ie/ObS6mRhoasvqFJDpBXc8D5GIQ7bpX25EJ1sWL
tx8VFIHGAKtInaPZVRi6/sM1hPa5QYPft+quwdOfMn6keVSnFcID/d2mvLwhNAlf
xV3fscPHAWUbYmqJxnhMutt1PUEAkz76vsB2evOdaBbarJ3CRZDJVDLfTxefr7Pa
GKWAObM9Y+4BJfREAl+MAWgZ/K5YrrHeI4utUSxRoTUpLih0MB/0G5hqM3R+a3sw
OnaxyUwTUkl/x8fh71V2abxzV7MCkbbJoBQwOaLgGdbG94P8aJiVt+y1lml0KnON
2zruTzg7wHPzVH0I1COakvZyqu/qoFcJr2/dbjB/amojxa6zGL6FxCLEmemrzhhR
nYCuM17VogYIJvuAQoHm653seBbpzIyHvyTMhKG7Af7oHiJkWdEGvvvqQgT3hzAJ
SCheNn4qPvmWKXQ6jQ6Z+KPotjFbFklM16ATn3VQeWWfJDWKH0HdUFye0ffN4+39
MPjPAzN4zlX1WSosLVzkveMJsitrsw67YCLTFyuaTDCMQRXu6WZGMt/rgY/q9Xeh
lzTmd+5beGh/vpzWXSAEOVNk61QuVGutgL00K+SGrarEAFMfcnoMqVLd5gvNAgtR
U3e9YaysMmYS4JHkphap0KtlfdWjDLORGIs2j4xKJVKAOkujL7vpPHaZ1W7tshbz
0CQsxMuKOv2A0YWnkyW2WSB7G5KXXDjaLmJn50cegIjzQltgXtx73BwfB5zf4P5Z
2jUhCVSfpODh/fVpvKWJtrCULCJIANveu64F9B+8M254lSPEkBGR4fa7WcMbOXN/
txIagsUpGg6R6QwEqNF5Zsq4FK80kjzuKFTnajKcEDmXWajrD9D5JdDhS+dBDtnh
8HZkmx3Tj3wEQ3I4gTqJQY5zWeIpBJn2d0NkSqBKFQXGOSmBQHHRKridPGtRgMSR
VCMVbQDYRtxG4C4AcEoQMq0hw8nfUpoWc5aPH2ERFP7zn/Dm3mnvIhGfapwSl/bR
85CnQUHMCeTjIm5AGcboLMRzzaL/kTFJLfkSXlQYaHp6EXYVuTb6B9o6hFzTfBDT
AScQPtZ4yWd4W1nKZ2vOUWmHvC+Ol70xP1sorQxoInoT6Lps4IWzpyF0oxxydV4Q
a8d+G5Uyydch5/9tzOajlPgcJQACz82VQUeO23Mj5F8FzwSKJ+xcIb6NtRg1CwFH
9KdZfjoFoSxUMiIo6gIVZUC8JIIJhWXFDkOrzVvbWWDMzfiHVPgjvfCoCUTNYZKa
iBqITdg8cANPGn/fUL7uK3ZAWL419/v+G6cErpGOtYYvpl+EtPVuyZBYpoUf/bgS
awEeuErUl9/ZG5R8Z2TJxuV761YGiGbjwn+dxYKKf1jHYiQTKgbg7Gn4VkeDLVaY
yucZgecML9bqJhDOTOm3kxcUNiLmCXSPmnNbIcK/17A9G+ocQlqLi1HWofq31jmw
w3GGzD9/SJMtSMjW6/jHoTEJMeyrGawIU7umf3RxylX3fC8ZPF7FR+lxJk80jeqp
Zox/du2Scrsufz2a38owJK1Ip67Eb8+s57s30VnZP1SzxnRrdCN7DRDcYRdOytdp
WTHqkmFXfTu83hVyPI25Kbv7aJ2IUxCasxv90wdX3HuH0mNx6VKDOYuJTy+pKhb3
ejeDAinL9bU9OSzG9vlco+o+Mj4IoZhFMtdEZVIv0zc1lhsux36cpztcZwkjWDaY
7ookbyDUdT2k9OE01XNwzsJu3yE/gfHTPJbEDWJN9CYWjKU8/JuPS/u1+OXqAbnf
du3tmMVo2u00//mihr3BJQ3Ao2CcgJWe0KZTUtznpoxRMy83GW2LYCVvZyLfCryn
gHBvZ5IxIMBOk1jjuHgbfDJq8es4ZADvFYAMWBUC3On8Lbu5XJP09dk6s1WEoir+
We/KJuhrzlqBj419EkdCj+40N1xsJQdwelby7jTeZVIlJAATZtrhYzwtE3HYJMIn
Li9IiXyVJMrhOjyjrtBdjyWmo6m6BgUbDQZtgGPXLYGuq0+IgO3NeDnRNbYFYNfK
dsV7ic3kMqPq6Y7QzvdVkEt5eAAO3mo9K98yCCcfhoGWTmveekUh/vxQVZqrdxzc
Op5aYFnvFjtKjpjg3aKRgMRR3K5ji3iD2VvmUN2fj2sc0qKHMF2PCc/yaORL9GSY
2/sxXHQIGM9jHP3Hajkdaooqc6YR314YrTsBDoy4hDoqv71hr9aflLUsReKlFuHL
v+c2BfYzi7bVgnz4ONlBPyAevBdRHQX74djqLniWPZ6k1bE8sYmSjsMjIlZS0/3X
QRkmQLCxPc8jc7EsrB6l3f2cfc1t2J0SI0gcZvQhS4LywMsDmKh468rr4j7E7xs5
+M7rxjKwO0AjXplT1QoexQKbxgz2ag/M+L4vKGXPrU+vxoAjgHyTUZGnIxE1CmKe
y3yZAYy/A0GpiOlboQesN67DiD+nUAjT6CN1EAoTpOcA8fGiIxVckKtMCqQ+YNXH
/qU1o2etbAmP1Q76IwpS6cLtlmZqdxmWUG6gIjizFgiKl0A8ruitVydlVsZ3H3cR
XS32b9trPtEuWAcUeGzd68TIhomPwctUdyDAlR/1zH8cX2OstScgtp1TKV2if53h
jD7wpvGS/LprrJKT+33T11CcAkLIYT0IAY6MXx+d/PPbSQrdY8x2fI8cnsRJcoHc
d8Pmd+FFungbgFpwdp0qY4Qqdoa/JvEnGLfhM7cfOwk6R9AR02V0wPrQl+Laxh/i
wg6umo9a6+G/QJ+bmlggwrID1SeWhZ2ju6BfaPDfSpxx2iUmsB9742daZpSobJHF
xvbx6jL6OTDL39Dade6dQTcobIEY6N+6lfy+ITe055uPG6jJwPXITS12YdaDBuO4
HIrC/3TBmDWY+p55ac9T/NQ8hpLpp4pQaJoZl2oMX0DtFHtr6Xb6FXAwq2SFakLV
jrneqSokhcPzhJy8usEdgVvEPwtNTWPkCGDCBHxFXUsLgrG562r0n8YRgwqcagSA
1LLHy5Jg9QJZefxLLnVmlv6CrtVwNBr3f+c0CqGqWM60Fsqnunxl7HbHW7RISh2u
84OMmr/o/0spnmmAdHd+lATWnYf+S5KQwLRKbz1uj94WEGTH9YuA1Z311Fmh8dMo
9w16dQwm+NWyPsuW+tnQDfiI1BPHSOoNjjXHb6GCywnW444FuwdKO+csZq5+rpHO
QN/fg9t+0cxRMxAwj8uOp4OfB93HljUukzurMVSWDvXChVG6vEJoCAi8wU19NIJk
VwSHS5B8e6KWOf+ej/BeBp0hB3u6oafYFJodKFD+0AeSWBKdZ57ZwIrHGaFJdJ61
QsOWOyK6guYjfZXigZ1kxJ0/VnGuOP8teNW/KtkL4ppa3JS1fQCOWaVaXF8RNqRj
tFwQCOZvy5YpXnVmVl6O5gCy+VdP3ex7PeM9pSyurPqFiwGB5KYn+CTdQ4rEtQmd
taYoCKI6MnCDh/h9k4GC/twxoGL2GIBty0+TWxe7Ae7YyDnD637m/YjPtdpm2QMx
6FZ6VWe0Ipa+X02fXwbgYbjGvz2+3FqcwINhPPVaZgUxIjxK9bhBNZ0mcBr9upi7
PapKZSGlgkB3ZNDznVaGRckoYuvtYanjvAbDwgysKV3flBQ0o68iS3S2RvnpHWaL
8fTfcWtt2JlFldpRbAdeg2HcfQbSnBqinzl3R1dK9J3eMwJ0IV0vS80X2zTULftc
AViRTHzWmGi5X+r8gcFSbnl2WUes2XE/4hQa9PfF678mcaoF4J7BsVBJw02jvU7d
2NlMTH9a0c2vk6Jr3Fu2HaU1K912+2cLmTMA953GSQdLdKd6iizsIjWrKwz+zG4Q
omnEEeWLpCkO67373yb6Xjc3bkqtWHZS4yD+zNRw6qFPx2C/4lbcUlaEhD5x9hMm
5FgfbUvWCQO4dsGMXoAaHwdcBUtPOh8iqMryAEDMVeomzU3GU89VWCKaUqS2fe7S
Y0Gm6JqWd/EOLqgpkJvlDo4HqviUqXsCBNoKiOUQVMhTGujvSpqwtoi6aHS18/k4
UF6dxy7YLztoN9+e8Wm0h9WTryyCyGQ40gJr72Jf+uiQph6KSeYKljwe/9LFmE9f
FV19BAHNWoRS8caM97EOLnzxm8cWUFrT7/OZL28QhTdjBb3UAfeMKYjGvXZ5wJdv
Zgk7x457ylVFAX2HjPTWAsEl6Ycf0gZ4pVogRxtJM+Y/b0lhHCvquf+/wy9jI8RQ
PX1RSxiaFJBldgKV2f2HicTb7uUDYjekXi/yJdT+HrqMctin1A9wGufvCB6poFrr
zcw6OfRe58fKW1YQZ2ovMaioj+4ZBbs0g0XSVolUEqzSNdfhQ6i0TVwIpfj+E1LM
2g3pWkLvUd3KBpHqI8HZwjGdbo57GNK9P9t1wXOwvNLrYJ6qIJ4miLpf/hbm723r
H0AToJasPkdgCTRpX2FGscwXeT2Ap1hgXZpDwKy3sfsWFXWYK5LUiCQb37WNFtNh
A+mYRYRSIWmNzY9zfy9MwnwDBt7raua+h9+HFmRAwHY1jEgYlPFZX9wbvLhuJIxY
z93VVhDdYByOx8+069H26lqKBBYUoxOt9rw0pVjCcmkovDI/H7tBAxuqBOANF+3A
cE7GK3qy8kqi23vVHl0usL3pxsfs/ybMBOJ6vD65+VXZWq+dk6x6sM+EUDb1qRje
wLPTNKxYS08W4370qR1XBwCtRv8ozj1TgAvQhwrNTE5l9dDApeanH/PlzHi/ejx/
TVxUTqXctILL6N5UBEKo89t6xFN92518K8BBMonAGM8uM1NyExlAyS8HyofrJrjc
E2YyJvkShU3MxwqLF5o82kzGA1NXtICJa0OJs3e7qNPi/J+YCS7UyPPkFUaOxJCW
JIavdrjZR+3sDlDxQBkT7OO4IowH5UwyFKZfhM3zBckNZ0aZxt/wHxsRYzVednri
pkhO6gp3vFqeh1x/h8HlA3dV4dmHFlATRgDfG/hkKAKG0lqRESxRQnEoLDC5Vege
5uCmfHvdU/g+ZyvwCiVdcatLnNUKpBX4iBWB9JGJFnxSed4TLtasz1PQDr3w8uBs
kk/YTr6yqjQRhpK24oSCAiBLpUc/Wpy9z/yZzFhZxLqmYe/P1J37p4ZyyyxzYB4E
mN31uiYMH2Ma8jh0PQkrAL7PheOPpCLyoTPco1TSG5gtIR5UIvkQS34jWd+OL0oB
B0NwX82RGYM5r+VEIob7bI3JocHATON+lZXFyrLzB04OWpk4Nl2jFrZcj+ODsi54
6CEZqVNytFB02bJ5o+KUPIZW316BFQTD8eXdxYoER9Ryuh1ugzz0IElYTRjy0OMk
dT+Nno52PvdvIAzBaZdjryV9OPLNgAIIuQdDHPAWwY2HBkqBCbR3S/tJB2aqbHAJ
jW//IpZUWY9oDXTP3CScWTaFUH8qLCdwutxAGVCRRh54rXQdJ+gVP5BjBVlBEBey
HAN73M6Df3dnqP1jnC6kI+EC6cnDlg6WKuTaev7MPanA1y4vGygw0WWLEx3Cbghq
qISYrKAfVl3aqtx2Eb2d4mHCUX7TGEQ9e8ev/j0Aqf+rlMT9cG6ATdBu2Dm4oso3
shcdFStLpwlkK0dU/TdrBN0DbGQTCcABZlUzxKlr7u+dr/vsN9e1ZiJuhs2tT5VK
pYEg3takfq4UrXhXgVEcvQtV/LHYlcb35+ruVdl4sqF67EaR+F/lCrkoE0rt0phU
J/iL7RfY0rRLBS4r0aIn7KTsLoQg/+4rY/zz54PWE6yNUE7P90X7R2N51Zla8BWg
BeBjvpIcMgXw34CzHpzlBB1YPlhvpcbdK7hos/NzIuIR0mjoEl56igS67LokMAtv
FsGGbBVmxaS2uF6IN6PqKZzmMzQvn9QfMRxOZg3kAKpRUyrS+K3b+UO/eNLRJMFQ
2skMgmPpMoHnYTkdj60XmwRtpcexAkFSYYEuIkIHJH9poy09zPXIvSpXY0Wf0vyH
ex60phbWgUr5q32d4fuQOIKBy+gHwGLg14fBTc0nEi5465nqFMVDp+pNvGv7EpUw
IBCjjI+WITZ7AlROiPtnnTLiPJ9R1x4fRkQdFuBlm7C66OGIYhoJpGNkJUqtVbLW
nQwRWRk360hk3IgfavcHHRuMzZztSveQr7Yf2WSppnSgaTZvNSbByRvl29kCPRZt
pie10lHJqXir5am60uRJDzSki+GZP826bANOl/+mdqh1ETmELj/hnqS5Wihf89ya
f/7VCgBmYcXsJIjveLNnkmmI704St7dOpg5cdryRk1Z5W9YtrLRqhbi/R1pM1Re1
pJb/ARBxGtJB3dfnb9mz24U7IqEf+UlMHdKdZ+N/x9CtnZV6iPOn9Lgb3EsNlrl6
xqE33BDV+p0V07vaiHETBatkONH35m6U2LCaaUxNEuT4qwL7vsBYe7slu1Ja1vDd
y7so1sKfDOdv/tMs82jIEJSymwcVKCmqyL4+QXyw66TsNmUvtKTIaEYcBuSqepkE
oX0BH9ziK2Z+XRRORVfhqdfz+TneWC+Wadov/795sDPWJ7BS0b7juk3Lu9CLRW1L
44U9qmSVyARYL+70SpHm5ryOSrECV5PBR+ZrTDq0GfaGYya8amtyrjWPB93KO3Ah
sFAAA4bLayq2FLDkzmfjFl/Uik5i105ZPwGuLdrZ1SaK4cjGzLBUQjVMbuzqLf/b
CJ3Fu2SCQTGm0Z6JTS2ITqIhL46iDTWyJbKJ7TOkOz2alH0ASwpC9IDthw/Xgj18
MTPNhe4DOvE6KV9uFM6iKKeIqHq7jgtSKcJBEPW5BJUvFCXjqtA1j+hfivYT3tt7
fEs6zKXn4RtoOiPDDAhXQq+ylmJIqDDNoDlyAPiN65dv9kiAG7jcB/rcCXv8g6CR
ZmHGaK3wTNLWV3mVFGE0g/D4j4yW6+wrHPSOrigBkBmMws95QBfOghzUbHd1Qs60
j3Q9TEAjhy5r2qnwoJtlqWEBTPClXWrMZJGGua+edmYYXoHA6GhW1mF66U9eDxTF
kIvnHR/zkLDYxHhyyxX5ai4wr1GP1MRazlf2t5cMBeFsNxQSHU6wpo20MHZj1VMx
Ox9aT9BteESHleYl7+a9D49Odc2t4jm63xI9+JC9UTC0JjIetxeJ1NWoWKmF4VY4
80w6ztwjPNXNJPqggQZFrKscPqipKVveMxxZCUQQWqSQZFqU4wLZNr1S0aG47nrg
bRoEVHiqwg+TWbKCVh3Ya9DLQaK6j0v3DLwIrp0WH1wIFzmAV8+XMyvabLmqu9xB
2NGFFAfghUO8tiF5EwVjpVbrm2uKiCmdiY9qBoGEZWUfVNmtToha0jZ2XFZdvBHV
TutlRGi2dUpA+635Kfr46DaQWTKTZfS2Rtcd9tvirRZrMJEC4Lp+Qd1G+HQz7QQ8
/VWyk3r5Bb7ony4qjr7w+NsziWpzKZSFFv1MJhF8fuBCur7PB9SFdcA+nXsmdl1M
oA9nX3xYaHPUYlEHMKjFiBSmw77fVEPMahzj5veoTj/ClSRIpBjdrkbnXrSI4bRu
3qaJYSNhJ89lqk8P2BTeK61q5vHXjIPZdzI+GD8uVbZL1kkErte8pjqjPGA19LRq
xPgLNAJUogUotONDjDcFNqpVP1Z0PwKeJ0YOMz7h51MBMhUpO6K7QZS1n+QUu1r6
BfMFt1ZivPaewhKN4bOOEGLTHCxlu8OXJ2g235qoKK+bmznLRmXFiEw1UIs5Imms
7Snz66YdCpqkhLiViJt5MUx0Q6PetilUY5q8atPL/PGClkjCLUrg/JHi4+WJywBT
aNhwS/qeZQyr0VSIhHSuTjeFgjdEo+VWYqV2HlO0DHMhiuCmplpphpEySkqLvp7E
AVPPaIXo09CwCxvGyafCBqoY8EYTB4KIfWVmQ8Q5qdSkp2U4/lV2DHxVTAiToBqZ
G+/po5BUnSE9wayIJCD74KBMa/zpQtKFZWvYHjL62f0OO3YnfFFPnLHMaOdSUI4c
VkufOfxaFJBPeMmZ5HX3Bej3mBqWzB0xv4XSep26DkAh32BxfoCBBBviuxJ+SGS/
EA2tUrpuRYU6DpG8/gyqfTRrzZM3oH8Ff4BrCOWhRNAWL1zN7uAtxOHVGmxnKl/q
xLnR20iRiAqYUmkxxYzZgPC1tUs1FVR86lPbltthvQlD68jnXOUVaSFgPV6+jc5J
o3QqC2X9oRbtjGY7Xoje5zq/4u9J4oofWVu5ktkZKvbUjcWdY6WKvMHeyfsovoTZ
8TF50n6TPFgJmX9sRZG/NMTnVK6HIc8dT5vQZ7NIHXLaDdxa/wT3/0+PNrTxYzK7
YyMeOXeOSsaG1/xU5fowd20EYrZOsMwFNTmTPEJCgcE9nNV9rt6DISO3LrCA/uU3
MQ9irXanzqMAeeI3DA6P5tdJaei3tyjwwMQ0Py/wA1SvXFhkif4Rmp0Q74rG4hXt
Wt3/7dVIkBUe5T+eYlvy5ONsKeNCSsQIJLY9mxwxgMebHP6YRHeLvk1RP11AEo+7
vIMbYHvfXlEcQfvCQgxfsWPaVs9NlFxYmSgzMQoCRJZauMQjDZe6Hcvnjylt2yzW
ji21qIRAFOF3FYYlrsy2C4asOZpZDRIo70CGYdwujukMwZbe2EPQPHBQQrziumlT
6tNAzMhFcDrESWkfhrcHHqXFKo83bAu3X77MkNC9zZsa876WF1oBDmP4IL13ZZc3
wi2zkEeknIDJBFRrSOFqaGEAyGFhTEotWvjZYg2+S9cAe3H3oMO7tWPp/SuW8HQo
4E5+711PYl/3Jee3zuEltyNLuqiGw8fOn/zYxY9RrU2ITxkdbNxIC0Ea2rOuIzP4
m4/7h2SzdnOeIGGpK8epXGZlN0AKRMPf8mZkJI6kguESaPWoysBZIwMOS5zaFeYt
6/tfp0X6A+ocX1ah0Fq81GXhX7B4Kpb6B5SxhY28rNrJxFWQGuBZgvO6+cgljxsJ
tMjQrgL3dXPXEbIy+aYaeAXpm/cr+VNiBSpApam6oln6NpsJ3YuwR0bXBBh6ZGLX
pfyA+hHH5BE0SR4OYsm0P6PRDqK7e4eYkTN4bzWT3uYO1eN0M9hs0me9QpobiNa8
67k68B/94wcPaUeAwlcaryeVTC4mMQ0UKh2a0FuhExlTuSbwVEsMhi7rCpa4Kl9w
d7yGA+svhDF/UOAC45lLkf3xX3xaOcW8Uc+EVi7qtCfGLlPfu7id1z0MvtdxQMN5
NVypnURRXCY4svg7HZAeQzklIJcCzpAndn2gGMF3eCCz8LqXURiaoBH6y6bHDNRM
mDu/y8JyPlVzI0opDF18+Iaad0XYwy085AOFYRhB3Ga3yUH8DFs7m7sYndOf0j/Z
jhEUucfTvptA8dXLXl6Ce+SZ8kF7GQm71xUPt1SWssE2z1dKJHUK3ZsohrJSKjcV
1LzSBmecTB8+sE4fKJCdDYP6lsJ/DxNWSfDx4NpeccVlMQIiAu8Ub/fY5SWeeki5
QCor9LPe0weVXufS6OLTvPpq0B226U3vWztxEM9+qKt9x2K8RVE9EGKdg2aIcI/f
Sm5HSLBd+jW7jD2GpNQQu4W37KkAHrtJU0VjcOfvdwwHF5WN8hZAEPmzvyo30pM5
8Ho0DZzbnP0Ns/E7CNwyONHzFC26j5cXyTg75I1wDmjLM3hu/9XaxTi5opW/p3GF
7CeoSxMpL6jWrvfCJabj5CW2tYCM1UqOZN3XuU7kw4kyFcGzC9KtNtGhWiAzvAQC
3bgvNAMy/SgvnzV6wfMDHDpe90LAYNeWresajnjWiDcjWzzySx8ZBV/7HvCZSGSz
0R74cRH3VsrV16ugWE01vd7gj4ZJ1NdB567np13wVvnIbmCeOXvTh/Bc9Ta3dj4J
+zwi9owc03rIROsMM8my7N+fFXC/eVPphn0+EbHpbS3IboCTIWAKit1W+TItsRMz
qUKFGgXxLUruHoafAWJqlzkzkmmYHhKNylWR3lo2arUmGrH29uKbRmgKbePJ1bmG
QjCTPPvcYs+TtAouc3k/urp3VNciW4GQtKKBM0MRxK7YyuR+RVdQZuRdEwm8+wl/
NInzxO7p4LekroqzLq+6uk3alhpZP+kqM/9u+v1T7BGZ/8pVl6UZlo705VTIMSwj
JulcWFaxUkrjOQJWNaDQkWgf2zaWCBISARZqkWgn8RLzftThG7ODsbOQfFz0wn0q
K2+CbGQyz7jcXXAIjuB65+gcAG1yNPXjzwFQCKZ/4+/5qwVnrsVoFz76Pzwbn7GM
8xjg8i7rb+HHlIMQ2uRytyqdIt5pokSFxyoREK9A4za21q0d0WKNU8Bc7zVvdk+m
dWaPUDHkWRPtGqO2HxiF6PMHWfvtQr8wa46hbIGiOTiL4B+N9q1qgRmLoJyizX4z
noKKgTYzj1un6dVP1CHnI4lZHzFe6Tb2KHevA7Yr+ngROKDsaTaB2Soc476B8eD9
y2G0vDTOmZv0BoxV1IDCXay0FzpV3U6LCBw1YU2yVaqZ5BjJr37r6Pm8nQ8Eh7yd
QP+3YnvsBb7bVvj8DsA9Z1wnrv4q0mxdWRDStQFrhfv0aCJket9/1bGjiq2yRref
sRzTD2t91XyLvvH/imK46zsgpEHE686uXi9hKRJVZ5i4P0h5ZKKUjle3LPTfXjwr
Ihug4eZ6IDPp7Yhvzrvo7xl4WxXm78RTyymUrC8d0VSOryBRMtEp3J+gy/GVT0hW
N1MpDb2Irm3sPdY2sEx2BhbzIl/3xYBTcN6wABbOQsSRe72spDOeH9w6OKZtUpgY
03UAoDUCJ/1bpmbupvUalru/gwaArrBXWW9N0l5Wuffyl8ahqvmNs5v+IfGI9X1E
1SQVtTc/ynkraUlzVh/1SgIzHT20pROCUTej6wHjpjtPGsgRbNozAEtJolRAlV8F
ewMvyPLkv6bL94riQ6rOOW8iVuY7aGcqSmzGnJrfXP+1TPh7Plh88P5Lh0F6824J
5lSyGkXKomrFTEIkDbdI5+5mxxN0NuxN2ESOnF5frqEzD38QvAC3zp3b4p0Vd3tq
bhpd8ItmswFeSPmrRPc/5cZAKrt/do0dd4nif8VuwKwPiR+HKYA9syBWTVim37Z+
b/Fxe3OC0Jh6F7MzEgoHsZfWo8T3dRSr1dscmoJWhAEHARgjf8AxKLxco2PSYvqC
RP42nCIie5ZRtIpxO+pBzFpfwSixZwy36FsCx/gGxywC9hVftrLGZsUQizlaSuXf
XST3z1wpVrazjTUSuM8LAHjb0ejingtbdp6tJXWEkYXHs28PSMHCcZH9asnQUatm
QzCw/4OnieujkvFhHTtiGHEihY06299imMHoMuCCXXYGHpdc6P5E2n/N78xoIQLh
/SuZK+MFXl2HsquxTBSNOCMklfTjw5Th1BMvqsZJDR7Y/S2osTwBinahwmBlwJ5v
rRa23+Uwf3FczLIIh+stluBn9rSwdtUMhff5wOVc2UqfGkfRu5KwfTFFfr7ktFcI
ng2KykucyMNA/7fDHyjntGWk+wdU0a/SnAuvKsXqYwlQaZozPT9POTQyTN+RUd7V
j4kb0ZodblSiA4r43CCYZD7s7lcX6RhDVdykZuJuNADDcTsyHESFmytRFbdlpckK
ixI0biYCWlZkPe3bGbfKi2GZ+BfFP6q/QisWIoZn2vCGaz1U/xOpYOmK5vXXKig7
xc/r12+LMwi1ogBVaF44ag7jfi60zCdzSAkq/b+pfREj/KlnhZgZCtKkyjNQlqtl
6RFg6LNC72w8z7c4TunOG2qgLtGn9aV9sTklDUoPSyIW/X5vmyQDpULyWDJnjbJu
ODVI1fY0HrIG/EqkgdFst8EaWoggucc/XA3xkuX+zMv32uztAXj5f5w1EZpQNMjv
Dig9TOYd2R3uFps+0Q7NQ2nyel9eycno8MmZmizPMcXY4WEJ4OQPJIKv/ORgeI3R
h595RFUd0a0Z/a6pBuZwtyiRjfGq2D1nVhO9UiyBgqhCSF7SOOHd2vtzn7S/zank
qTHbsijlFK3ZAyWlyAeeE6e07g76JejzF0kboGKKL+JFdKDsdUJNloqzsRlrzVtd
llBm3/pZK81jibVsh9xvkLuQaLq/jCzA0UACvRoJ9tNbCLRMbN/SFiC974nT3zf6
CuA6tDtQJi71r0ivTjkVI6yqeSqqRWeBVzfLxGROs5ddJG+sVSxq2wBeQe0BEPM/
9alNWlLxSuqEA0Nsl1i2W80WpZa5ZcCRekjRjDl69dZBgLtfdgEleaSdF2hLHjz9
Mn1AocEXQ8k098DBeD7YttOQJcAybh5UQ/rKMXWJNATsRTDzgNNIzZfIq3Fd6e8f
M7kNK7Cr7iwqytigIPPJdxMJN038TMYG/x7vEfHy2jtbT60cytgDIaDT3XYqvYy4
UPRgVx2+b+5kQs8bPnD/13xlX/c+FNbuJ6axvFnNZ0GSFYMfyZmya+tiEmcWdLrg
5Q3l/0voX+zEnryN8PAgRE4m10B3xMZQuHk5YbzPF5GG0d8lnQspa2D+tKEsg0OI
UDh8MsYrSM1QUn2lc4w/9iy//L9z7o7kSYv5qdZtCdLEgUMYNc/x944jIbb0RagA
UU3FS7k1dW16DAkCfo9G8T86Z3KYS1Vv6d7gSd2Xf/Un2AMNhQuTILn0R1tKxISt
hrVhqzbuG3zwl7ESlXFFiyEPmH+ss91Q3ZKIwhLC1yQNkfUPJNGtGlSOtaeFsZx6
rFb+c1jJOu2z6djTQHihlQWTzZmlAf+Xdz2WHfPvJXEWkG59ml97FI+h4+tvg+i7
BxQE6re33xagLWSAYDpSJ43h+DrLSvd3J8A1pPuKEh/b9+/t/lDIqkpllbE27psV
Ml6TJQJkDgjk+GqNXtNxYjQFK/CcMBRp6bpYQ55JZAgafnMgoll+5/Pe0Z/cEmki
3YiTQ2d9xYMPQJppGQWPmOPuQwLS9svPxZH/9DPX6HjqRXpuu4yr1e3azU4ANJ8A
bhkkWFlwd+XsUAhkSCUHwyIubsmx9gR/j9KrZb4YDldDMpmbloMzpBhPwvmDK9DY
j7tZuJNqOU+3fn9bR/6JW7Jve9RW3quQdcKEMNamjTFbxfDRcYBT20zmNV25X/gx
a0sbGo/Sv6iHhRh0yp/IXSvCol/WmF4nCcPlzWSL0yclV12ofEj5AVM5QYiMK+dz
sPVCmWTOcRCTn6mV6y7S8rT4QfV5djd56F8CV6Z+nACkVqL5R8igGcIU5Z544nQs
OJQIOQPvQ/Djdk6XjNLCaovZQykQ4o+dwe/Inw2UKGjWKVyv1sMfHWujpe50PZjZ
Zf7Vyy9v3OB1WdybM4J8ycbnGiTn42/Z+odtUi3momysdW8SAitq3pjDXrruv829
EbXNhqxtNIkan39IOnwAiB7hPGT0r7BYuIeYE/OVszbJmUVNOjItBU0yCTAfZtcU
q8Q2Nk8t7JBeOjkh4vvi/SG4myjeGmDZ8X4vAZ6l9QhgG4gfC+y5WtHfe8TPE7Oo
3wenfji2nKWGqSoyAwRVFxTJtzj4F5LvphbEkwt+rQOrGdsQgyHOzultmrFd665S
yHxjwOs4pXzou9CBtXNBDmGk3TC3Yxly3J3YxO0AkH19IBBeiaJm0Gg0cXUFARnb
URTheNbG3CV2DBJz1/atGsmHqccfQq5UfBKCSgSC/zatXE2lTOrt2KIHm/3rae92
UXZ074f85Vut9Q+ENHRhf4vq/do4shmWTR4ujLskQgJX7qUtYCsimJwtDyOUTHTJ
gFdsCoWJgtBLY7+G7IvV14AGBXThLv5x6jAnl1JZ/srKW+Cd14gzZNbADDaJGdE4
HYEDVhaghai8hzdEsOwYleMOYTBlV1mva0r2qELgtu/4mF0SrmNC9ehua/gA6l09
mMQU0fAzKiDRbzaYl1vGHeqVFnR3InAus2qAkjSp2y9MPUizN8L/ChuueQa4S8va
FCgnFt1VRle9UgogEutp0xY78oMN26dhJflUzhSfmj22YSL0EycqK67PXHrhCxnB
hG+pF9MnUyC/VcyG51wrpmU6R8uT1eZHAh60zLu4E0EP5Ahxp5Ygn3aMVSZ/kR5Q
qUQ2J4+g0bz3csfp5+6qJakAHWv3sl6HWi3Im7Gi5hD1S0WUuIglDbPKoUAN+gA+
GjlgJZbWuG9AqzWXe3Xo1FBq6nmiCDnIKTtw0u5/WyuPGkWna4HyU3msZcWssZZ7
H/etA5JFlEZCGgyEqjl/oY/QUWMMlHpt6ElNJiDghhB3BOjwsH2R9gXhRk3dzviu
/CPOzPhuBBpTHLoF7lFhBPVbpevHl2oQ9jGrVr5828LaaORbKoM9Fq9bu0yXgo+w
0p+mJIot5QQBtfcBqZfhzudu72Gc13s6RunFyAyJITHSsLiAnq+LETbS4pYXDz5f
EkWVM+Y2BxWqiDV8r/11OUB4VLwACDutPeX9MPJKzE4QoxjJm+twOtN5/YMNKXme
mtIik5LkMap//q4HpLnU/giFchGllzPC4TpoPhHyQ2CtrevygfKRAf+doZPiYO2k
4Pu2NLnUNpktln8ER8A3Lm588PcYy/WVChcf8vZy0pXsY6YoUa5YMCSLvf0RmImM
w8Bz25jQe0eiZ81mVEFYeVFmZO0fARlWAAI47uG1D0yP6zmVPWUGE0Y8mdog3jkL
4FtZXCKxwNjjEoNAA0poslavf5/j8O9/neM1QV845u5ve0vBNJdFl8CjCsRESF6F
fxnhsv8J+RhtlK4fFPgKq+evSgHCGQGNQT3YnId1GdfBDLW1iuBVaSjj36NQ7VXl
aAqRI4fRwZEDDay8asJEUm6tT6UHrkPDriTVngIZiprK0ji9CJx2qA1KsJpwW5m+
ut5FGvW4Hh01DemNU1PZArSWyVK8tX7n3KFO/Td3ua/48eYCOX7dVARlKMBCBUhv
M+T4I2HtmlwtE2b4yciNnrRmqPN9wWlMSFYd1yR7n9CfMlmcsaPng1yMa/dXm6Ff
/YCUJwsA6+yrBgwuMGr8KLw3VIBf0uAT9RICvugR+OW1qNIOYM/BYHbDejmQAv31
ypp+eDp1KyHZPwxJPav5w6RH7e+hXuN5oY3/wEkClm/jmMgFNmBoOE+lQMFBSxOP
oSu3WH1NLML/BiTeOR0/rdtSl5QHKmoa45dIJKA+R1WmSaSWqHV0YvvbgH1dkCrU
sznJTxyTPMU0twwar9mUiGAFZ0H+8jGnzmERb9GVV+exeDhMv8pla9CYtC7fnfLe
w6TSp9kgpSSBOYAC9snSIY2Lf75YSsfWqPbIY16ISt7j25fgD+SSSzaSXL7Qmifo
FxaXXfUEjJp+d0tgz8pgDTyTPEiHU/Jl3chmns4/TbgJnnNTQebdg6njU4alZNdl
zhXIehNoP0x2V7hmYOYkgzRNX8gVXvBk1nZoJVv3Jk1GtuTXw1QH/0SeZwEQhp8+
BwS9YeXpR0qwm0Z2CCGuUvlGhAiCGIXGe7YgO3VaB0fIHrqv/yV8sq2E8JaDWcKo
ziSJOdvz58qpS7W49Cpr1zyBSsEKkcLUsEoOMc3Fb4csIlBEjDq6QIHRvEJn1WzV
YIbjePXm1Dus+9AKAkaohJUrhY6itdCgdVTnyQZifJg3Pb6sVhhku+7YrCcNdCXP
D1NBcEEhZGATCVI9JJg4fYok+yPrBbhKbTa6AaetWRdhonO4/SBTd6eBdCIuWX8+
sxuVkUF6hYvDqqZwtZfpWmavVG09kBcVGVZ4wjWGB/vgn8XhRE4bA03PEZB8zkE7
OQQCgOZqHrHv9ihA2hNMutIYEM0fKYLwRq5cZx11hLoSsdf1gKIl82sC01w5B1p4
zyyROebCr5D4KBEs4SzvDD3G6s6oA6QmvTUF8JlKc73/DdVukPCOEIAXjSOBDmgV
ymIRVZduh7xyT2OSYRx0BjJnMWkVJ0fAb48DqVe+q3lcuzWce7n6f1Fxib1uBa2u
cKonbK6jwVimo9aEvnl9pMQiNS5fJPjxKuAZIyRueuEupvpETIEVKlL5ht2s2NH5
H3IwHu5TDnF4WzeWKyVtIlx0pWrntsLjuD6i7N4xmT0xcg/2mX8yrSsb5aMtOXgZ
IrZSCMrq6VkdsDv4KLcqnHh2yZW0ARGctRTtRrKT/ub4sDgDodC9CUSplAJ/tGU2
jjOD3UqhXFSaXZjGDMcIFMCYCK/Pr1t4u7vf0KrIuJC9gSh2Czv7fKms2BgEm/uR
gAKuy3zp8y22nzBIQ0fXMjfvpUbHpeRzUHZwHet3YoG5nanodVitkxCIFAJbEBuT
CpGq3JW4yAswjU/W5Db45RVznSZv1F/f+5m2Ng+mcOZ90r3J6EkgRazaXfC2JosR
Rh7Pe1G1wuHfdUo5Xyh0O9aMlfg5O3W08/hAW5i3WKcVF040DeWVAv+u13N4PKjf
XTLrRafyyCWAmSKAXWqm5JBNSYmdku23DqqgBZ+LEfh2tUieJszeA1S5dEnBp8yb
NUHIBEKs2skzlim9inTX0E+cfu1jMI5isYFBWOSNW9eisCQu24LxMloziy5A3MEg
M6hlaQNRvdCftWG4jd7iI/JqWuTWQir1wi290n0vaq8OdV65iZz+tFCuIVaAL6Cs
+Th8PsYCyO2kXc8OOQr8POuC3vCFqQ8sbS7H/FfqvU9mDns79DSbqRexxmVaXZIN
OgHr2fcPbZWmP6XZATfECSpeR7bNE9oH4jpHIOuZyPRStlHeIrHIfCp7nWaiVmix
YM8TT8NDdynq66WVRgxAjRDk/zkuxkeUz0ZjfuPqvfmvSgt/pNIegQU6S14TyeRx
vAVKL+RAG70uWdY2qob3xRw742O9MKG5/3sd6Xv6HmhaIKK8PMR9qJ/OCnrH14mZ
MLb2UghRyxjEVJW9uUQBipsd8QabCW6juN6TsI+7nHgJCGMgKpOmjH9+WbBU9wBy
ab5FTx8xa/Ctkmca5XB0Zy8aMAv0G0F4gOmpbjUnBIg55+ePWcaIfTTsIFkDTOi/
unOhYivWZhwh99iCpnEfprNpFflUkP7bAiJdWhlcZukpRNKGrMshEu+1clGyEhOK
TbOhbwIz1ZuH+2jnkLrybCcxPjVSPPJMysTvNPGyUquOBLDXI8qkObN9manWu5Rs
EYcsiy7OZz0+9gmaPq+JsevJp2vQUxKEodHCzdgxEo7R72emL/4TPzRSsYzeppMM
Nro23czckcUGSgftIBRbxsUVdT6pQQdL6ma+gwQJZp7G9N1mp00v90WlxIlUa6gb
8UMwSShUSJthb9GJY0tf8wJRe2Qirfv4EnEZRwOa0Gd+on8gAqhNxQgGjsUVZWWP
So4FO1gVjNhOLY3zNEAb77QTwOgq2FzZgnaY7PtqXdD6x2CBpD6lneR4o7nfVJu5
tbt06I0YkwSzqucleqChYAk+LOIVP5R04G/UgMyHs3ojXzfwFvWUcJZWfBsNFUPq
oaPshbl04JV0aTYqHp1lxRWVdLS4xlIdBvIqu8jP0nhMm+TkZ627gS0BwP0pNIxY
vYmlUeNw4KYjel3NTBPfGY1eRvQZYmJ4M3JSfeFZN7oRGV+rTp2obCcBYd40sG/7
HYT31qP92u+XkY4C9N+vklKxwWdOSSuumVfamlBKJ7AUUGQjfZ7G8qkgoaGM9mpk
xJvv+8xH+sVGJKMk9XJ5pSMRtHyVYbdfSEt1CQSlMAaMu1Seuo7KSQ/TMui/UD7O
hreydf+YBuRdKk/m5xEs2YxbszFtVWFeiyEAYpptHcaN1hR4DdJqQ8hVzsXsvruT
w3fBtTRUBhUvg2QqngJgg+JbK7QdROXGh/eIhwgjZ1Xj63EdaHQ7Inf1ElLxm2AG
5dPw8YiterqzGex8VJkt2cST11dsbDHBLcRMaqkbAGZIX/5VlPoCmQNm/aYmTrWQ
jbKPiTSlPjFk4IOwOChMF3htP6lcJVwpVNB7Pu3vbSkn1bSQNFeP6N5CQG4Jc2dR
gbTkHtbS4xfYjk17aVL5aypjVwbp9s9huDow8uvF/935tka82cb8O9JxiCqq4G9H
bmYmmjtZ63YTMlVTyiAquKnC2k8fyy2+upVoleymRaSyRDJ1JCwWUm06v5Jk0OTH
mgDDQujZTbVtRH31XSvBAC7K77AraAiHvg4YoEI7KczNWGxQfOViwUpYnSj+U/oL
WcXnGhz+Tpu0nDaom+z1a7ZdTpYG177kn68ecuTcV3IqaiVM8zl67lVSp3uMTxJm
uuu8oG12I2ne9/2d+FfQqNTvz8LdYb001jb1WC/GNaZZLIKEBW39Wj0Phqj6Nlcx
AbOh4CKOtDlmmuZWMm2lTenuPZMyKf5RZucCohQc/vBlhnwNY04MS8PZOYPreA/T
kp1BvWIQQYLfvKsAkk+RwC9bLdpipWl9MtEe7XXZoEAwGUhABtZyzzepyXGFWoX1
qA6KXmOWXUkR5BkHLnHoU0fUMxjWJPUn0J6HnQG6VUa2B+mppGniq4EVGgSHIs7/
/mOuRVQBioBFSlFD2VCEezxi5RNSjdBRwrSKjYZ+1HVuSWXrO73nzSUKLizxYm5v
YhMGwREJo3hVXPPWpp/G1u0kg/7rJOfQxM6P4WmaAaLNhoBouhU6ygT0mgBEwDNf
YDtgqtp0v8uRtWcLjyTWX2giMb9PnWW0LYYghinoweeeoaDNuOXcMhKaZ5aRiOgM
8vKjOkdhaPmDYkPdeF350zlnETokxIQkUsrpAje739I2LYwVuOI7t5T15/oeXI3K
JEoHnDL6H5+Ax9Vq7kKy/NFz4pNeKF6/lPbrBLJtbSuqHDfx1Oh8eOW6Wjn2T0E+
9NS0rAEIaBxPzk2TAnuy/EmBnxxj3lTbUXyAFoRbzshTnwyUZZF8SgZyV2ILaGBZ
PLEPaRSq1SHMO9ZFjgguzX9A1u8pPabgNeK3tCxuCOCs56xlD1jN9Dr3QZ9mECX7
BD8Zkn/2MSCUtKZuOIpWr3u79hvjFt6/Wu2yqzUE3vVpMow3lTz36/WjoUdqtexq
8U+Jc9mGF0bOn5DFSip0likZWlptxvlO5QEhhFXbmkkHDNLqX1laNWa5Edk4tCyP
gkNKxxAerWopSevJQYjYAyut+iczjwHHOeaNVFXZQtXeu2W7J7xKFmv5ZTiREtRX
oYXiyvHJEHa40Acm5Gje6Ed2wdTNDtlsbG1GC6YZJKNojVeIMaf8Fz5PycWcV+da
dIg4vfMfU1/OvKGS39+zAv7O+ZQfoh5CWIOWSB+XIxXZb/vOpgQFbbSphLkT+9iq
QpkgyiO8cHfpym+B3/9OqZAm1g0UBhjy9h3ZUbvxX2dA592gWzgqx+cpknafyWlW
dgckM+62aPMp18eoOODZ5aBi2OwaGDGIQ1lAGKDDJQdttORuXHdxDaKPPXfIHlbJ
JFWy8XYflt6FqNrgUjNWRf/7A61xtDFPcOH8Z/Efu9upGuuFFpkz62RnDrwjzOxu
1FhbLpukIbwRlQ2JrC8ipZjGeeKInRSedAPcWs4+xqp5dX15kqi/rAk31Id8z/6E
qeGFJ5BaJPC8cX3hnh4kfZrkgakEE9YlXXTWq8AE+M8AwzyOo8CrBKgcSCQfz9+3
luZnN+Oc2y4kFnPYqW7PlONi08081pYN2JJmbxzS5v3rLwIFs8UVpG573tuJAJSq
1Y5BSxvsAWDRJIN3442UOPO0yol1WKdDFgdcXYTD4jgoJHwEQ/LpgjYwDvRu3CFH
PW93y9/oYC2hZ7hzi0vgNYMVsLcAg/FKdMHYwSTyL+QMcSpiZmoikspOp1rZpYVR
30wO7rqg0TeIwAqXhsNWQfWliTIUW19NKvSCOAPchliX/1c1pC5tzPTz06MyaGs7
JYXaKjToC9xr57gnHWSI9HiJGsWk0J0oK+lqngpn6X5R/FxgQYG7TaEw2+uNnqli
JsU7UEgCQRsQsQ7jMpktetZfQmr/9qF0rvnsRXVx6ls9pGoRbPsVaXgIUhqVFeA8
QnDKAQxy4PdMvrbR6TvuhdczLa41FUvS5NnQkvGqgUFFJe3idydtAZLSxwULF574
POF/Vq1bNknj3NJhpSXhAg1/uWZP94BNuar72n/RmAvfJE9hRMy0k1JR+dFGzVJi
aOfjTxFkqB2tR6Hx/CTF9gmvKU+IoRKX8mmcKFODctyZtFH1ly4NNt8+/tIiV8xM
Rm2StGzikE+3fRoN9LLSd490saCDbXP+l5yJhD87rAj0CaQc5E5oiC7Bb+7qb5Bg
q2z8vWUwOZRVCM/XdbUUvOWy1vHzzoMhYI0V059wwEncMuvtCW6wMGrljqtjT6Af
ISJZZrfw1U2QFPiBEsu4p95unkYks3ysANQs2bCeWWk7NWYmeEFeSnWJIeTR4M+Y
RJVL/GL9CP0CL5vRiPQSxBY56a/Lg4lQa0L4XCI5iEgN+/7XUY5NovL6aYtuMQJD
GS21QwMni3oNu8SnKoWIce0G8cgYOWsn9QL8nniZVZ8lEVE3BiELbloeeI1GC+VJ
b5P70YLEiHTTOmQBHOyt5++k3bwpOzHepSBKoXlAohUd57Od1eIrqefkZBgbrkPi
Kb4GC+Ed5nM4xICh9WFbX5bKGdtQjdh2tJQ0cJYYOxTNFEcUDbR4j7VlPvEg7k/3
niYfaRfV05jpEMpUwfflz6RxGeOJQKwrFxz92B2rXOhXmQT2zQ4pnQ5sjlrrikE1
h/i0btD+l+oaxlfa/fc3ta0mIRYkcuTjlP/VT0bIK+nonSyYiWdp+99Zz5Lx12Tt
vQLw/WKRKpTZbRB0Ur4qKzEmks5g18nPvYwX9xt7pLxIun3bZ7yDvLk5iednLR6M
4PkwRxukTnlKgOR55MFfzznXsWPRZBJgkqvVkI2QxgE5TNLCU/Sgz3GlrhUY/PZx
drbL9NuDV4EYreOXejAcytzYiSPRq1/FqMOM77SEaQqmqTGmu+Tmu3WBDruk/dOJ
Ai0cmqJO7h3JkpD2NhWqQbLOLvX42KBOa5knAJAR/9phHRB298ZVDl0GE39Bi9TP
XSoEHGKxybYvrJrirWNiImBv35C3AvQs4KDZlABDfjQ4e5Y507K70QSNj9i1lG1s
i4OtfEquZiibbz/HOaFjRAgeX63Stofbfwj499OvMtrFi7NN40Aod0QQ7r9YRVMK
WUYxsJNNMuKEdlL0Z1est7qEhlalW/nHNk7GASyBWlUJq2EdPtaHc9kAib3urORc
XmejZ53YN2cpcqLqsX2j86OturD/rd/dFKEattos7jurCV4AxC2W06lL70euFRTo
ta74lmULq+yCpZDVfz030M6HKQb9BAuuTv43tnGuQgygVJW4uMlbjjUpDYyb6dF/
TX1MUYtF6ixrKztoMdu+tdQG6T9u3PPqHyWNNkBIsdxEeiAhOqJJKs/1vgEw5DG9
R0hKqwCswoxLFMNSPvryTJcfE6ppXBixogIOTYWLP54tBQNBi/ZHoI23eyadeBak
esUI+pIg00FsfMwBp6/q3cx7ZI06AKRUKWN0PlVzUv+OnA+2amriEvu14dl+f1OB
p497wDp5HDbUitF9RqzJJbGTGMiOitRJZpKmIc0Yaua4wIG5LAS6hsWasUGr4eWl
/E/LXshJET8v/o0wsN+rRyEs/NswOrItb9sK0iFl3G9PmCyFJZd/iAXXZWzU9JDb
HtmP3tmPSWAVVt2LpUJmi9SRZ5pKvwzDRijSJEuqmx2fbWU/XBOkCUnxwp+fEHDs
4OLFbUNfD17zG74DXG7L+KZl3q/nfDxjOWd5xqnrE83K8LkTZT+lbx+cs9Ijpyh/
aRGwAvNPbLAg2Qm0pv+H2d09lxJ92M5keGXaCgA3XGRWgfyV9bFzL0I5Tx/NTOVj
fMNANPhquOJHzMTQza2SsSvVcRMqMPV/u7ORb6hkfs6jHoh5tYRQWoZcRU/rT/a+
39BR7J9AVZPSVXvMkpi0KS5D/85n8D/mAKuTWC/k3FPCUzL0uNwMsSgteqgSqiUl
+3PJvkptevEioT7iBvIAugbBtL33NxxSf9+fw7Ufxxeu+8tM3X32xTsfT2RP7+b7
GVfvc6lS5DUdY9sqRNbeYLSfGTFlVcKE+4PCIzbx3A5L0uM7Ph/9cp+FqRMpc/r4
e7Ulxu2Bo5DlQHp9qRF3caQSYrV67OpLH4k6ydmIKCrEIw3+7mPoS+zT1ZHUuEyR
Wblfo/cOi3h91ngBcu14F7eLzH1hz9uhrxrXY2ca/LNsJs0W7PsXa3sVM3/4ot4k
JMH0xIlB4vgPSG01YIcpT7TQ8tiElWuBHNzHYF9jE7hSmgoMrHhFkUm2Uvc+OWSw
2ppAyyRvJXbPSg4taSXgF6RCj2G4VCX0ua9y8DGzWFcKMhPtnYUERul5fc0C2+p5
11u6ZuQW9m6m0HpoPKAEaTaLr4Icy+P5nEyw2mNtcHNMy1MvdVWjR2Q0iCV3AiZ0
io+MGlVu/WcnFxfHBmk58v/Ooz1OE/ugvrGjRGa/qG1ExS3J+FcsRQn3pVS14J5C
0pzn5bdRNJMWPT40OBnNLVZyKnAv0XQk7ep8ulbYog4hPnewj33daVb73XtUlDLW
e6CbJLmNZIBlIuYWrZNd17EV4r/cwkbea5bixqUxUcQLCXTvRcRaYmF71yPKGU6b
FsnWX98OEAt+gFWt3mYpq+uLTYbsvI68qTGYG2ozobum93hX5Iy3gkgzOp42AMtY
U0bXG3KP2eeDwgBYRRX7VSdQJF5aMUIs2GEneSMELJqQI17tl/y08Jt+RzLd+ZbL
3xB2j6JYASs73554yRjiqQkSMmEAXnEwOPanJBojN8BN8jXK5+TjFd/Ac/Ak821R
06+8HB82/Q5guPf9ol3T2A0TTrMOjANb4uMyNomVFoG0qVYU9e4JBc5XU4LfIFMT
5KakDMAsf3QBjM2g73+4fuiRj1pHIxjiQ8G7hDWxWQtRAVhOcNPyI5yVlEDz46Hv
YBlNQurKlCxDMNz2Psbsqr1ahOtYSDG4pn6/PGIcZ2OCyoOnnuC9RxE95H2tw/gS
9K1aeZv5wvCadcR2+ofA5xxiQ7Zbger9W/xYx1Ojzzmrrjvu4dMaTHmC90bIJ5Kv
2d03GhOkLOWRVQHdS/fQKLVP82WXbIlFj/HsDoxqggpuhLv9WS//VELjScFaPCFg
lCfJ2FExjDIgMuJKbXgpDr4hNX3AU38bplLQLFUBnYl9OkprzP9QooXpXAadVICg
ee5s3+IsHjEaGFdMNZkPvV0MN53QCDUwqA5WesXwic5A61+q0gRuzRVxuNd9HU76
TzbL296arkoKd8E5UJynp3TOyjwWgLNjNZA15J8sPLN2hJ2xlCnncm0p8JJQVqLJ
WotdqZtMx20tR+utNuFOUOF8LwD86tebos+JIzpOhni/kNgd6Xl1Wiigekw0+bA0
kAqE00324WoUs0/Tr3gxnu3DjoxJtNsXf3GxYZikfN26AJs3hR1NWZjBaND50Dsx
vtjEZ0o/l4AWTgSQDrci0qBOXKW4uTel13zO72AFomaT58Qe6bLWmc4RO6tiCTY6
X3NGFE+Ww1+ejO7MIYbMeB7iOXuWVdz31UUYCMOk7sZCDEAyEkscgGoAjnMfbKep
dZw1BI1k4AAEm+LYawhdRn5kC6GbeIXeHEn2Cikrta0MZZ67dq2BzNKSW55hgRGM
Y5PBpadeskJH78C2d6NaIotEN5540pnuFHfV2HEsYvztUEahehs1YIg9WmyaWilj
SZeqdmruzO5sHQVVWBeoUa7SedUDakjuARqJ7atO2AeC61Y9q/sejBSYCTuTp0Be
fGAbzsnOP86srNTXicSKR/0uYxYCPaBjxYlqhp/UMlVjhWFiamfzPm8Hxp6N+dFl
uOCKkONPLFR5AtO56ZW0AJP9hj5sygzo+UyTWwL2Rjs7K7Q1SBa3eXpFDXn1/5aI
Py19KSY00D56aHxsd/Z0SqDNAemWoXg5l/UxjRqAVqZUPrl/9rMdp/Pi6P+7Ik+9
zLF1Vv+nkhs1jkoVZ7OSqCm3mqHCdyTYicWJY4BKb/U57Z19rk9/32mv98Ff8GRY
CLNGhatNPNv+maYKBarqybTYXiDH8w95Nb1v777Rw02z5/W9xRfx6nFbZS0pDHgG
yimmj5xrglRZJbOjT/PNYuK9MXodEs31x1GzBtATPH4ogb5EdxZJNUx6sXy6Y+Eu
8N8l6ifGbgRgbtaQjeNGIzuojUHUKHSM5WoJu90iv8ndlYH/cL3YfI2Me4hPA37r
OHcX2RiwxLOSlHL93h3RKamxrmaWxn6flObcFJ3WWgTzSiRO+fCrNle0Ch7Q7hUk
ew/m/fK3RJMytw2ZBViL7jTB2q2n9Cx9gwjShaahmJX/iSloheoP+AXZFIZ4+kZJ
LXS0zz49fMUYv3JGWVscHAz0tsTqUgL5n0q8J44gM2kxisWFXDBH7QuGJrP2Au05
eYYF6JhS476O9JVauqcMjH2chTTLfw+ot/ZAwdtZynlkmX6XMAgChp32kmO1okOa
lca/5h4I+HdZJBe1RAfgDKEze4I3jYgaPmO/AFP7PBhlFTVrl9zWkHhlYWpVmNMX
LSBU6e/8F+cYkxArn2pI5kuNlmGzGJOKYRHR1deLImJdtWNxZs1jcNaHfGPL8Gez
BUhv+PehQ44xXeleZqaW0GZMCvhpjT45wxk4Od1alzprJnZ0s6u1AYNG7/QQlHdv
veU2OFhTaNc/Y0zqoZEEUnWwi0JMtrK8W2Iqpo+cUb4On41kF9suYhcmbDwiHP84
tvP5Gen6U/tRLazpd5asOT0vg62vJkwhF3PoNUM7TYyjyyYjdZb1LwJKbbRFALfY
8lp2g+7i+Y50manZ1sW4wHhULyiEsYeUpD37GGO1whJ2dJsSgEMnm8AhHiOMThwS
Vpf4r09jwYywCpc0RK44MiSvr4GPyKGY28Hs3R/HKrN2wwJsP4WswBwQgkeP+esl
5ctME+mxx+NQtGuTqhy3zqlt9+Me4jZpP6BpSB4EDlM+3z/cJ9XsX6ptK6ySmn8V
kcptJNPhm4OhqibhszkQwxEVHUsb5jO8fp1sbeQYfVsweBASopoTh2MH40H7a848
Pz93akaoeKFPX9VT9IMcu65bP3J6ESYgv95NQ2eBbXYVta3ahXjKjgDlUnbEI6v/
h7291EpS79pbvHysQpyt80NSn/WRfbE/ZRHEjJP2wGtKIQYqz511tYsDWoArM7g6
6LDPW0VYFaBf8V04OjyAQRU9a/CE/WouLtLZQbM/i3azaH1/2LHARvLFOx1EpfHw
rJffCgrnlpmQybaRbKISvcFEgNOl2ucQfxzjWwcO2213qOa3oCLGWtfVKmwfo4Pf
fK+A0dGYcs8b0nmp6SqjHhjWgAJ1B59aIRCy4PEM6pFGAngX6DviBZcbly/QhWGk
+OMxOoPtSKNXWh8k6ZYmVXQzG+CNtImb8Ro7uQ2DhKkW5VfhxVsIGnKy+FW5oerj
tqHbgpf0aHoj647oLvTWqXoHkud2IoBr0NkKXQsbX5C/i2kq/CTtU3axazmetJYu
C52bu7CtDIgag4U3Gu8s+zt9Md7vG0lCmrXLVr6zygolQR8YZaf/8ilf0nCLpVWC
yalQH+CCwc1yfQqW1QGC9hjq/3VjUIlrDYP3k+IuZqNonTYwOedpAzzqfC3ya9+D
8YsRMMhOURkvsOpo+0DevNqsP57fqRYXhwzMgNGU7yo/rvh8E15gnxpEuy/90ieY
n6ioAYFZ82g5+BXEQ+xlomHnMKmF9cZp4oBCfp/u+yCq8hvXq9h8qh6HrnKa/iOB
KtdCHysjEkrFKav7n7O4wJI1AKzoFedtjEUKgXJFVwv/RQt/JGQr8MdsEuXI4Y9R
sSaqLSA60Ndqf/OpRCusTHQjSCoAi6l2m1HE0TwETe/1Fan7wfoq7HxBriLeL+Nd
qfWBJsQSLbtt8oYd7kP43shjVrdB1S6JBZdvQo+O6kr6JPvAutq4i+2X7Dpx/VkQ
xGmFaNunVIC2Std4vcGgVIfL/JF0kBWVUUereLUNexL7oO2i5ieDlkMdxiYEzAYc
AB+7IaBXLl6cSJbDQ2VAG61joqkUGoVQPg5XVL0QNt4Hz8A9GkCCJ/Ia/pudQyf+
TYJFBhPyf71FGKMHz4uJDKc1KirEgyE2CDnJ6Ofw8RqUqF3+k+dTkjeqwG/J/r4N
KuNTMUCmqfCggX3o68/Q16vBLuU1stct48vepm6nQmgTskt75KtIuy9dFoN2idmc
y2nUW3aUQpuW8XOaaQinDmxLECLlO9zyW39DIac6ofOAAJVbxy6N5ongXyvSKT1Z
bxkbG6XyFjiP9oLrPmqKzkBRR4mlUiUOToESCIKWJskqj/MzESPeGylLVOkgfhDe
J9+yhcTh3w3AnAUtBJrO0NhAJWhIV56/M7OG6uXhbqwNEmyDxGKS+7p+K2H7QZmF
yo6sqFLQWS5hdMXEyDnb+MJqa9FdGwWc/WnqQO1q7YkgRImrm5NIsBgg88cxBQ5t
G9OpbZ+cYzbP+TnsdAlIQHAVJqpeqEo/tpNVygwJpY/L09jT4p4HeFBxRsgHv+XU
E/VGEVQ/PFF9+w6fIcyFbLVXBss68Ebw8eBDk8RttRMwEttckB+pgsaf3Gv/fI9X
7nmesNX7GCNhtV5fJ5+Wxlnw4LxsgNMcbmgVq5FwkRpykW+GcEohU7e0alH2fspE
q09GtwMlbuU7Cji2tp4LsFYLk1GBTkOuVroblkZbWUbvEReo83skOrTCnaqrjD3p
cmrgohNpdXt1+XzELoD1E4Hjyw7zdTLPFb3Y3T163/KXeJVsrn/gRXLv+tH+ZWTF
rurIoFXXZsJ+buL+VTRUUqcXmYTJOjkdRnE9L/96jfI6BYjnv0AaMsR6hSywnF/N
iNatMzJZGFOL9UgCSnlf65cMl2qUzIdrzq9RisBFrypH2Pq9EkpzYMikl4fJG+K4
xhahCP+Q3zSKKsDSVm3vP2lXMZjCS1u1AV2QXX7xOwjnkJRCilnOVNd4o4RHyE72
KuinrLqfxcgnFP1QrESwK9KciyJf/bk0Jrpq1BeLfdKa9ZYAGXXtkjVUL7aHT9SV
3Ps88Q3nujikAlyrp41/k6QmdyU+x9him22vymc/5H4vpFfGW+mD9Tajm+bGENzX
RXaqlfS2ItnNiKmpdYv7yVAqUfdiOBDS7vdO5Ezk2cprHaEu5e4bKrYCA2r3VHHV
fVN9vXZSVnFp4iHmjzGiktN7xvzb7gflaM/IuKz5DSQyQ/WrixOXwG3FlqnHuFND
RcxVCOaxiV2QS+OXwZfvup9Ywb5ApuLbodCM9F+MTD2RxdjT/RsULk/cuatI3SCy
h5SlMn+zSiMPATvl/DUED+VpodHkxWbMjL1qZbxzfk35XWLz0toLmeZqtaIZbamb
0Yr8JUd57nArHYntR3CaNoIh5s4ftIP15/Sg7scIrabKyeWzbzuY1OnCsnxcy06z
QbNjl9i2FTMwrmqUVfxrIGgzckX2CHxsZO5j4A+4MxGFHQa3EMBFWHn6TXOBMXru
mSGXlp5j376maONDaCRJ719vxY1MIxemoHrdR/gBAfXRiMv7A/g07ULGnsVuxT4Z
3k3vjApD5xGVlUp6BjpM8dj1O9Zj3Uu2H3c9WVU3r+Pr77IyO4sCw6v5WkGliGkf
rJYBulyrv2ogEi6O+btcZfDYU2uthxURcg+ue8YUxVYa9CRo0uGLSJlMmwxBp+Xw
/wCSW4685nLjJ6VZiB138gUbxToiKTyqyFoVVhfX7pjJT3jG+QHpZtBPA6F+4jso
7ci8o/W7LX8TVLfHsdCD4eo6f9+nunFLRfzJXXnBInl1Bv4H+8vcFqRI+JovriP7
nTJni6FwPrpUumr4qDVu7bzi6Xeh0wUCh5O5SMLAIpypY51t+hJZUX2fY3xOtxYi
7BuQY71SVci4X5yD59KW8yLTjBc4l3OR0CUE9IGp3NmJMFKHE1mxZDIKJouxCNks
nx/WvqzN2yY3ee9cmnCAoik1NJk4dvL4chCJShSwFZilWx21xCU4lAXmNGbkTGeQ
gpUpzCyzmE9D5ldODMHc0LBlb4kEG1IFOI+TkW6tqY15+wtc948ev9fUB52EF0o9
Vcgo1YjOyDrWPErIQA8IGqU9/afb6LRLy4oMqNnIeDShFjfcUaGzXQza+zcdy1pa
qehuHyMhDhZvh1QhVdHtEuSUAK13UUq0HMENdzQjTxZEnMacy/9nNO0coZLcBoeq
7k8xuTwbIzL1tsBfGCST7eQK3LpqJK8TOMQVtJ54wdeQra1Zye5HfWWOZVSJ+/pj
uqwmbQnLq/QUjZwLARtZO9O9N6VVEEDt714Y2Mcqfs9WVuOQFqKhvf6s2/xAsBEj
qzbE0EkOwdJxzn/d9DRUHBQST0GC/3lEAR/nzz7h0Uis4xMx9DjR1pwiTLDK45jM
f+kb7Oz42Ddr1eIEXlxgn6AHPNKVDWepZwNrpRxfRotiJ3avysCSwldCEanTsVKe
feYDM8dvKEjKlp/Rhl2TeX/KQ2G8azwIEYlrbtCYE9O7czyOgqnb1e/Vh+i9HXx8
laIZSZX9PuXRyLsOBO3h6GlOdnzBwYbv1lpP9JWFnGY/PTZANXPo1UQ4hZcmdRCu
VJoGbxsYLmUoDLvUSHAOTzurEA4DuOsv6x3ozbOyTpsQ017UcdFZ4aOT0mm+ZV6h
TzHbQHXO2llahPieWXicF2W5g0ThSIuzuk0A2b6iMpYr4oB6iFBGBZA/vVzdu36V
CZI9dva5wYDQb0g7lX0IqqOni9GEuEmewz2KdHVnKhntGwT7LYGHLDG7WOoyafgp
xpPZYUHguq4vZAOHl9G639xs8KipdXcDQwgEM5AA2N7r/5KkFu6xdAXkZmn6wwF3
LxdrrcLCztySbA+/TAO8AJH47vKgTuoCOW4K3pBTVp8kARheJsSompqqWVG9cKdc
kx2vO6tyLTMDHST5M3q/Vu4W+QgAuBjaVZ60xA4WprdVRxRLwq3Fyp/iGd/uzQbR
8lEQa8D5RlskfsKqf2WFj291pqM/TV6EosI08LVOvgWkDdaRkdNz3gLb6PNNfYF9
ALBEJnEV2Fc9osIB8Zx8j44IAP5P7fpW3Dm0tQhcZZualiJMyq7hhFRXqDPGoLxy
Vjzu4IRzZSQB0X3xojnPqjHyqx6dtv/9FGXTbEca13JDiqf0UK0Y/sJ/8J1ouaD6
zyU+9nb1B58HkHEPiuoiWUHlPKmgjbNFtGbX7Gdh8774cgILQzP+0dpK5Q+44354
HQ1J/3yckuWhyUBMgn1whG0w9k8pO6BJbL7MNovFrqvQMaPeMvpR2gJN7+xNZdQV
DteGZBio90l/UR1sK2FU77zlefqVidvRi8OF7iTJv35Jd5FpaJMNnPjpyjkj1JbT
ziJ6BlFMUU0iSV7tXZLmWcz+tjMvss6Q7QVjFUB3vz8859wkqWTW1u6PUw3OWlJs
SoKhIXWPtLLRUplXDeXscyPVrm3z54g4mT37gwsKWX//S4LDIbDL2ydB32J25TnG
zLsaK3DFHCu54Ds2Y7w/Eh0OO+TRtUy5SBnkWOoitIyDEmTRhwpE20LzEnUDnYK+
n04zwJvunPojOnjeRq7jXVWAqBmKyCtUIgfJbdUDpwnbUf9KbZKni3IRF6sMnW4h
9UI6675BGKTFLBNCMp/jgy7u8+FYcig0WAJReZ2kyftZIHTBsUPLkKzGxzp6TyKx
j6SGGa11V0LAMeFZUgenXbza4Ss0UrT6RVPk4awMbla09VXyryLQ4vsw/FVNYwMi
ay3WJsv6Zui1UI34VS7wPU9gpisF0+VX4Ufdszf8nbiFxMQX3akyDOxM3tqfUz+X
xWNWlllwXrov8WkIGWvYZJ3NNzXPfxTLJcGwUZa37bjc8hobLJLb/tUppK/Aox1g
veXOU0JAEi6TckpO/LGi/5tD8SRegna0hkJx7+kVIpPMXyach8M+pEH1aV5jDbG1
EZtLpRM8E2H1o9qPiEJHSIsQYazG57ICElvG+hRMPFPdCJWJpxTBaFpDzQuFjzch
ynVmNlfOBhEBxwaqZt0FJ+l0Ragr9wldDZguDNA7ZQBghOhsXdodVdcVqXtGb4qV
UKt95Fma0eCGzk2DYJOrVzniPOxDemRxdgQWZPWG2+j8+toviI17xUN5w5cL2hRm
eoITYpRQSZIs41EJOl9ZdypvXBmcsq5Xj2zgxDVFHPlXf2KtRfHM5wTemVC2nFKE
loP9hxXyWYvCk0cOfZZ0q27fjObA9AgKLQBXmzZUmerX4cla0J0k/O0JkA3XJaX5
P4L1fUPFbFRpuA5YQWlnaiZ3QI8/DrZCtSItMCOhAsFLpKaTqEl6Pm0SJipoM50r
2cCkRDu64qDS8yizc/eCMbJI3EHKogCjRLq5qXKQUnbbvH2+qS9JD57AClHM5Gxx
JdZ3dp0anIDwl45bGVmljfLqo4Ng+aWCW9f0WDwvbEzozFhXrYECvNlbaSU43+So
olO2gDDY1dGkSuBjMlzTAEHu66O7tk8SWy1CaExkjiIfr8YJfhbcWSkq/iGHJgPo
azdxldHZ+l8B2FF4YgEsNUKdzXNyByoVsSIjEyu22zmBJjI1Y/XUJvQ895IQI/km
ioGVRsr8kAZ62UchNdim1eISF+MyQZGK6sFD+tmZurxnhSYyXr99m9k3wWar2YgY
QhGIUVOL++xLgdTuvbi3IX911nYabPH6lj1qAuUcWdHqnvAQ+Ik03Dfa/aXn9jMB
njjohFY/lHeQqsOu9C4J2/YG0yKk8uh9X/XyytPZ37YSZj8HiID45xCH9pcpn/N8
o/BxLaYPnI5k5JLkz4kd1lWq1HEL5vXg80kLHKVbwLZIiwozJBDloaEddCGPYY5T
6MMEvFzJLPrXg4W7ZSRQNj0LHBFCM0fJ7X3d0CtgAOV02X0W5xCsd+390x1sRiqs
o/ICNqY9xSsxeufh0F8HqUa6EAUbkdw2Q9hfOYjC0S3sJQ2gXBYTFYV34UZN/sgU
PP+aQkfggpNlat8FO15zwGoZd7EUt40xBX7SNxaYLDNlAkpEjDr7SuISTjuIjiWZ
lUC32ea+f8+AxcHEpkk3YKZWHOxj5emnqt6IVdxuOGfXaxvNMe6kjw488V8lgsgf
v3HpLERvljp/FMVoZDKRzaCpPY9qHXesJhTsGpTCGUJ0fHcVoGKtyvVHHDXrmPFZ
lRdagWU6WJGZL+RTxU2/vopvrWLa/qprxBJOeVB07ard2PXixjwZ8Ud8e/DBuMwc
/SdmAFItAvvgDYBrbCi9qn30tSBd4Z1m+hU/LPIY2zY32a5q5vZvbQRyWMetrctI
m/pvXpCYPnQVBgXe95w4G1wtCaDPnOtNnfmALOB4DNPRuuQA/jtEaNEG+dFGnWX9
ScXaqIRvEMgNt1VhgZbnWkMcyjM9nBHgfoCiqgYYIoQDbkPB2UbyNb958ZE3kOAN
FFcxRu7d5UvDX7sIkR7vDGe+7rnWHWLG719ZUwHeqrPc5vL/NGhN30ru8ko2apQe
rGbAdGQ6/lVBPadQwuCXKE0sWO5dLnGIhhXFcDeBAl+JD4PnyqKxMA91rkSOzzlC
nHS6IP0H2go0mw4pc/cQJSdUaGgYhEhzjTdj2+elOiXW4OwHv3xwy92SOFqUyt7W
/2ELtYLZiQUUKvZ8unGYUW5coInosveX4ApM5YdNWktbtHxhtAcMdcfqyFKtoBgC
zwftbL8TwsXgl1nh4IMhAqvVlC+2YYg7DI/yh/bYW0raIFk6vfpWo56rOZQBGP41
0DNYWc/vMwKkF+0S/xnr5/DBQeZEkQjNgWW5C2V28S9OmGwu1REQuNxxUcCuiTBS
hAKWKfwryddykGDa7QzK99wIaAsMUlxC/l8mlHfHuHnEVzcFVldC07NCKhn2Fnf5
ysKhIWEWBl2yDPZpRvHvKYCpD9lORf9BXAn0dkyG2daxpw0xE5jIlIVonRPnCeuu
0qWzC/3jNQfGx+jy9N/6xZWVQbmgTYroQUDaZ270lNHTMQ55ldWU7VIGJYe+3OOF
Kz6rNGOQprB6v1Mrwl5sbN/MZF7x8zq46jxYEStRueoQNYoB83Q63W7a/7RgOaEA
SKagJ/GX3sYGL+M9Pw0LrMQhmJgszivo8hla57IhLyHeS8oT4PPTkDk2+tXknY0j
ZY1i2RXw8+34AEfi6yOimhYQ3AwJQFuyRiL/+wfotayOCUWM2URjUtQw8vLwnEB5
68169pDnMDi4pGSxHFgyi29vMIqlgC+HUvR+9eKk5JtaE6GIJZkf2L4OLYlgKmUJ
lpGHH5maBTs9DDP9HfZ8ZMowvsvuNLvceZL1g+bcbQ7+fP8EvQaDaLXyi78qJaaN
UPm55PfZRDkIrXTU1aDZDTlvVGsgSjVkO0KePct9V1pbea4QErgBtGxjY0gDHZdu
56pruD6QzRQr0nbj4DedqetQ9P1In5AHKLtI+qrNvUAW2N3W3GQ56wothOAwC7J5
ClvzmbGnVdiCs7hYT7nMj93lTxocxGpsUiDmgjF7AUNdsaZMMLjwg7ricXLbNFRx
eAQL4qn2aq1Y/xla/6NcyGt/OF309N6ptPo0Qp79k4fqThBQdmqt439u7hKFWhBB
Lgz/g+40z/lsVllEyw3C+icmF/Tics2xF7hRqElDAaFZsBC6AOGNvX0TOwIWojoI
A3XDLkEoj5cEWj4XafiXPDpOJ+x+fOv35etuBdkUm5FCbRG4kr+0jXKU2WYNtYHx
HU7VKTXKtHVECC1GXNLWsEa3OBNfSv4ZDP7TO7BcElS0Ln4tQKrgpUrEqFbpqP+2
GEBl4cH/i+cZ2wfl6s3CwtkFagK0Va1slntPnfBx5pDL+weyrhGM9pgZF1baMRPC
gePE1r8AcLhyawRRUrGrf2Qy6biXuxafqQccqgiJZJyJCTS+Nz1G6xU1GkNPYXAL
T+irkjW0DjqJO/gSFFKqR+OqKGJMwdUI/AtrsoEFlaO1l37Z+CIr9DzSqLfbXaOE
BzOfs5JAs0rEZEiCuFa4FkRT67Cb0n6isxa/Amj3jzb+YkNP+AhF8nPx0pCXtCap
yMnpGp+ApBcLjBiOq43utG5gYA1YzM7AEgZPmnfTYKUOM5bbABMuvBNypV84wEck
9sVZ6TqLt0B3dDxn2fn+y6U4K2hKjMPnef9LP/2rHcWmtbh0LaztTAYk4oXVFU0e
ZbH+qp8ns4i/zIcqGLIyh2DNAGMCBdV5Pz0PiGX5g+VLw5hlGJP9F0OoPW6uojTd
6FX4ni8hoASqjxJxflx5ZszoTE+Bvvp8ITgPLqEM3M26nqQDN+Wvg67zGPzB8Tg0
ukIucXT6tRaXACLN+G1Xpr2aWT5HFVrt9XiEljlPKcjurFF/sbHrWupUbiqwks7r
NVvceveeJITeUCONs5U2PgCdpVG9QPTdSDdhFxkXH/LjM20k4gjyo0y/eTJoqxWW
/I1YVEbjb9E9pgRYikNJZsqIGg21TPZkoIZRt0Mux0G1TfcUsWL78TfFM5wehI8G
8RB7/lrTpxEAze26bdN+OihbP7OpUbnE+7+ATtK11QUIYcwc26/qq+XW5dfuNBU+
ph19L45HrUm9g9jumMbN+s7o8HTZEabPOaTiw13EMls0b9TZnbWnMsDH75Z0qcQx
3cpxOTzDmnsMaFbYnZmf2zgjCBlh3K8VDNGyeeGtbmvUd03JncqRd3mv6+j/Ud6C
vunnD8KFpL9YMJW0a679KXhYIiDEcRO4FAysIk5j546H1ARCC4qdnQyHc98w/I2i
7Ef+hoiQ3GMV2ZnTtwYNnGiyDKPzgGFT+JRBLE0mGWKFzYO+NSsqiaakrR+akTbv
XIFzbPicx9UL0HZ1EjRG40/qkQ7+v8KPaLbAwiio/l4LSXo2rdheAQ2sW5VAt3QI
sPTBdDJ8ypbuic9d8hNuD/izM0uivJgZxzcO1+95rAEcb1Tdgy7fCWuKnxy8NHxL
IMbZBB1cqU+sRga281+BWFJxUDkdiYrFF1NUYhloZElJCDwceZHOtnovNXgYxhD9
gczkRQL53wvxtA8G9rrJ5FqdCIv7OOwUJLAJhkyf03NJHsjgTQJeweOlHb1aJYzu
MRWp+at8on7cMaThcP58HwmIJKATDNuNskT1jPQoRIQJbcZbjnjpmvdXshffKMLK
UWbeQt2xJ10Gqbzh5jnyI0uuiyxFeBkNdQWKS3rJ12IvFaoFpc5RFWelrcOFfsTW
iGmffAXsjg7Uodxkls82EEHg4aT3zK2GseXOeXQlcziPy8DIZepunP8ZPpEJKmqa
oAaA+h8YchFzQ6AcyNxB7fyiVGYlMfBHIjJDCuh1BJmo2hrcKOxfmbOyxj3+MI0P
wYEoDBqMvh6ZgIeLltquoqOBVuGrE8H/0lM6KW2vmkadUJh+w46QDTIRQ8kunBhu
OkKS0l0uIaevJ+prI9Dult/vz9TscACQPidQsjnji4bSXY8M1RRhE9GsOOEQmSwl
IH7pu2Gut3pQq7vOO6GGcHo8XZ6kXO7zeVPYPAHJL79fSRDtNBCJ0pWG4/roqc5w
ZZsvUcxKZ4VahgyjwloC4+ZahLZGb0BgXzxjTODEUZcMgWW9AIZoiT/+85mAqcMO
23W+kGUU3idPm14KLl+D8xlozDOmFfTlwGTG0WYUjz0eLFbwbgC1qB4MvoX+feS2
aYAWZaNVehjValBmw0Rls8sHH+x2ENwZaeZPxb3BiklAnpn9BOjy5i8SfEKtmjji
gyI+0uZSw7nWAa68vclY54nPIZUIgfA8UqHMYHOrMaYOsq77pfmSlWfA6WLIQERq
X198/D/SCr5YJSky76vAQm8GteTnaU07HognEz04GnSFcuTOTHg9LsDJMPG3itjj
nqyfbcw2YZecYk9XJFE+OBHmlraTapvSLei1n1D6na5Zx4bjuefpVYHUhvVsz2c/
DbfaP3f1VH/04XFWIA++GlT3SnV37B1Ydq9qI6+suAd0wbVCwa5l9RSOV/4lUGJ7
+PLM86/KVIP6iUNrpj/Jb46MJl5wmenR8ES05vz4AK9blO6hmuZqcVskFnkZ6oFd
yXIODHsze9NcpYVRYV7zdRPjn36I/me6UOpbUvbSN0fUWKuA1XUgqn79u626h46t
aX2Vc8HCSwsPnU8R4espsZn6Z//U6O5RciryqTSsQGCuOJWkf183FKRhNV+tzlg2
oGWCRqez3R7T0SDrZW96JrjjW69+nPd2+0YQm9BjPLjeDXAyiFGzcc4fu/wdFuP4
4vKYjkbPkWfHNawMJv9bf2/4H/SVc9xh63MN89+5N18hl+soaFqF0P9UtquFiVg0
9EbCN+Df/NvnOseYbmyXG+CiFUfowbY3w6cpmgKHffpOcVa39x7HR4+KRt05EAsy
M7wwmrfmZ1EgkD73Zlk0C/8zuunORYmtnWXzOoc2ONOoi5Mpx6KNC+MR0r1cQZEt
Evp2RvVDBy5e1fSM3h0uaVcrLuolor0rsn607sijHOqdZhq6tpEiiiKiDNhHXa3S
7/4DKwcPhTyYP9XGyxduDnqhUvClPxbL/9J9A9rdv0fjjaE8CgoaTh+GqVOl0zY6
WVKYOy86rAPzrF4r1HQ3Y2lhWK+S4eFXNYd/LKH5SiUX+izeelQ8GM2Og+siplt2
aKPEnUC03vz6NwiH4nmDpCUpzEdL0WDpp/6TVwV2K1Luai0kges2mMfKcIzLgvvJ
oJUpzLeu6hZ8q/lpbxudIlVxIAmg1x0CfUFDHu7C13cyh4jo1IFfEF3K+Rh/YKQ3
mbC8MQvI8eTn+F3mjjihnsCV9OQfPzCmta+6LfRqRmfdjU8rgPRHOxdafD6xKFZt
pMN4at8VQvrrf3YttiCm6XDB3XsL6YHbnN4ea9AiTJwetdHGY7ksNSJSqxfVWFXL
wxmgGqikuQLG/f8TbM0NejM8abOR+JWf2QTAJ5vbiHjMhVfU+Ur0eKrSiCwfhPa9
f2KUegyg+uM3nHNixWQOWRnOOj/5Hnh8uC4EiPS//dFQGy6aW5bNGDbnUpRWwMmw
EMDwNL5LvcSte9xAEDy0gmPyAXg3rOeVP3VWdPDG6rHDV0RHGdPZvQ2EAtyznp+b
rrHOHD0eSmVJZ50ElKENUphJEbdXuV7XRmOjPGpT4cbRa+01UzL/aGBqZrKfsP0a
oqg20Q/5+ET7i51Ent0ApNGEN2quNOIa3ul6O5iqe5gIwsfTJTgHgef2KAk+1AnI
A/HhbpTbPwyQuf1YgxwWa8BWyr73+PGjPEzgVv6lB+QmKRMrh2JER23nbOVdYzN+
lZJq9TUcCxgRaysIkMHbrcWKEZb7Kez5+K3xfP95zSYjCPsqUT2Iu8cvaon8gmL7
5BwHBbUs1IuUzifUUBQoYf6MFtB44HQWRXYbxXRqv65Bf9vKYp+F4L1w1ukCs1gt
/vhByYnfSi8er0Kh2gsuPJgthFXJCfW2REl18uIXm8xViN97WYZtT/RzCNzIFPa1
uQrYQzhBgAoLvdDfDRhY1L4mqN2Sjt+8h0X12tOm+2qD32/DtRa/ZHdRYVe6bUG6
dBKdwNzlWx7woyYpdLmfM0sRovEDdZCF8W/KxUUcVVPxcPZ+hAorNXKBkGOMvsBs
8jV4HdHN5YKTIJfCtwDutye/FHa1XozZS1JpEVrqRsq+8NR+KW30tikoT1arMcvB
bB3OY01QGAQciZBdT1jGcJqHCqfr4SvcbCxesfuTOoBVVhsC6sYkJUx3/YiJmpij
PQ5ry5PEO/u+ivFG+Ipw6jKdzt1Qr2lF4hoosgJ0fxdPGB4Q2E9C80GRQb0JNiHm
KZbuF8maZ4QFt8baqGq3GvaZSdX0LGFHFF1jD0e9VB2qWsd38979j5JLuyJtu0kO
OUn57ffKGeQmDnW+UikouChE1oEs+VKs6l3ydVWDmY+H2M4ihn4iOB3vV14/GuPV
7XEhuo7B9poiYlFzpYeYkYaEwM8fdCH8Au27DFwI3XreTmd7btnjkQX4xsXWfmBL
gk0mMKSLXfodJs2Tm2GkIy962OETHwkQthXGcH7lvMvcfKNPpmZZlUYniuhYJR1r
m/fygZFOdJLyyCjQiwGmCoW7IBWYKYCrnJh6taEYzTHXZzigXDfvcrEQvG0kyJMz
fTboaJbuIpE6XCUiPbTYDbhdKlHKaS5ELvPvsOMqC24xR3fSLR+wU2d/xE/b1tWO
YpdvBipM1IjhrAVtJMuCr7VacOlCA+uJ9aYIi49DdET3xfR5rwSsy8WZmaXv9Jug
Z3yt4s3jkdl0DurgbQ+n+CSDjt5OkooWTAa7sPctZGRXE+tc23CnCxh1vPEaRZS9
A4TRZ3cPloMHiUfTicZgid8yRo6XHWY7lMcC9XaX1Zten8U6qtAgC1n4puZZZyKL
FozhmCJ92p6ysVMhO5UDdTal4YbRSx3JzrQxHtVuTPhjxFAZP46shbsvuD3cT0ME
zLUpYhQ5d5pR52giWDEDXcpyHDGPaTD/82dMKryIuTiRE/5hQ72Ey8/MBEr9n5+v
PjASSO6sj2Ui9ojjjI2LpQ4vhxZC4p09jgyo4Gk9D/Hxd8flDLw4h3yAKE2Al4rq
OALHIcKtJxCJRfwOY23HeW11dxhghXHYc/19uY38tPmcQRbcqtKWHCfODcDQsF90
Bf+aOMh1VOQ4pn0nQCGUYE4HAsFthtsnRK8G+9gVDq37mSYBA55TNRgWW0vRBcYA
SNpgNK3AUpb/1DIyDj5dKC3NyIUQbxkISG5HYwevgj5jDL6y2DZN7fKjSLw2/JCM
zWUWYt8T6YcpWAWifbCfaqIcVkrek052MsBXGY6xJKMvZJ2RK8mKHbkyc2tQysbB
Kp9qOzrrdM6Gtsv9zgMQQYqL6J+9BG5//YHC1P7fYbFv161B3gmA5R6TIVVcOJDQ
0u5MTJjNE/qS6fvklHQCo8bKkqusyF7r2U503LepKffmt2Z/PXQK2r/V0dT5WBQn
QZPiEqrh2gvf7QDEeehADBV9F+uYCRHD6jH6wpzt89dl031kDmvxwdtj6AI3uUDO
vOUbRLgwOkO/B/L5V5HMxwVX4A7vulh2V0kvijob8LC3SDKpmZ6pmHHAzmyF2lTx
9Pu4y3pEREqGYh/UqXnVVR34zTl95xHUaZJtQILLBCV5yVKwJt8GbhuIsIqEa76x
rJSc/NHE9OBJDQKuA20CgbomL/+EonygfyGefFF//wPKG2hHvRV2QbQ7Z+pQ/fpP
0MruomcFqk/9S9Hg2r86sAm54FrNMHjvEk7KPMUGFXqh3nXJcedZq44QI600Li04
mbK3/JSVgR4qQfaNJ6Zy+HqaW+yexbQbO5RIT5+H1iud7FPs36shP5nU61GozCKw
e7a80Vq25/CSc61ffeoszWuOTBo6fkrFStpt9TKUPlYFop8t6dLSAb9JaIV/TUjG
ytKHtmpfEyVcDOl9KaAkQSRRA1yOznlquacApv0+KNlEELqa94jJDaTC8X01kcrw
nLbnySYlrOaDqAxkRYF34WmoT/x3Jng++kVAi+kLvbX02K+N5MexA0LP2im7l8X0
X9qO9QW+8iy/3zbf5gpc66kN/owIrRPb4fOQRg6DTYyCQ8G+nr985lITAx8AGOU/
Ov51GhpZRH+pD7u7gSulhGhtdH+A41wQimavIkLB7ctIdkMOzNhNo2ustoB6HRam
aCiCPEVrYi280AF5k3OSTavzWOhg3KTskgR/wTUa7xwWi4RozjeH9bhhBd/X9rU4
yeOohWQi8gsmI42vorN1RJChwwnm0tfH7O5Jyxcw25BmJDNfEd1Khj3zEQg2awXv
gWYhsCH4yst483ZSB29Ai4igeaQPtmv/7U9mGKkODgdtBtrRfd7k+LwEx/wsbFnt
ENSs1fx2KnbdNG9FqjCRnu5xkSAG2WzDfnlyf8c2RmqepA7uV1KmffFpb+mzKh6m
Hfxx+jgKDGQhd42odHgbXtmlaa4EuHzoq5aaLetwTQ6AjQlp2bSdK9W5VWYqq8NB
l8OjnRQprQXsPC7QRSYhLTQwM9CzE3GXsciq3Trg9TAPgYQVepQ7knb7J5RY1cex
4E7eqAVo9FN4I+QABJzXaiY5CAyFlc0LzKVwK5QoVdjcRNXoiyVoVpuULEHI2+a/
yorfMxnVrKaVCvPXFsl/R5LO5o5E60KxW4zBtA0dthR8rt1QOu7+0AZeOBZHs4Ez
eabkAlmUXjqjI9cHARt5DfwoCwqEuiO6+n8rfnV2wBk/5kGJUIV8NZF0DBw+AJQH
zQ/CIJhEYlY8Xyfp2ICiEYGEc+irHDQ1200OJPkyMv4voSLzAESSUJYhQB/Q7AO0
yCoG1EUNCWGPEiIRRneawhSs7sV9mo/ytVMQ653RwXz3ygHfvmX5l1cWPMisLSV0
E3bgtJQMIZRuRFplfMWAP2ia/ksXh85XTSD5XEgOLHUDJdV8a12usMt+MBdjwrB0
NYScE5Y0cyha/LJ9+LV7L1b5VtOmBdRqMMoIMnvBROg/CvMETHqDfghtbj0j3XaA
sYx2X19joV0og221+EZIpwSotPfSYrPvmvlzZvoiJWoRpVz7Ix3gzUaMQQkgnZbU
Lr04t95RIrX5zhNyJo9ZXMx4keHQf+1MAgASZbEo+mQhgcG52J3kCi0ToNOgAwDI
S1r5tjbrMZ3BngCBjgIw4+vptSiiF2ezY1VrE4IsUfgBFQhQKBJP5lmlCoRAfgV3
bGBs0Z2r3mL77yLFGXuwe0DwHFDyX6fMPTbwO3sUNWoQgUSgC+nm+Slje93QlQBA
aeK17oYf8OHPQee+tqYGPMLXamJx9xEEDTfJS48LkXYCVrsqfRpzomFfhvlGjfP6
Q8J5qo9n302Ys03nIErEQcMTSNxDf3R+Rl4I9L8QmyxALlfPWPbx1L0G9WAf7JCI
dGky9LCfhjYYtDsWkV7OW2kV/ad/j2iIt3Qkz/ujq/Na1Pe1U1TgN4FMDX7ogS4i
/j32rj8qV1wTrhBsgYi8zAeMzGQS78R+DElrAgtySAAX+4NfLd6siQRIonNI4JDa
4mYp4isVTo+b8PGBis8WjccX60tq77MHuCX4c7MT+ywjX1DgxQFALAhcwLYI0pyF
M/T5knPNtN0zCF3vCkx387putd8CPbLx8RTiz/12pX94TCplj7FauLRvttzW/gAR
RiXFg3rIx5nuYLF5pxEIB6GJLs1mzkBNVgjY9nmlDCpq/iHpdpExo+KUv/H538ES
UmVLNeJlBOYmHlpoakPcU8wQ7pgRO01+Kebu+FcQH+ddJFFWYmuTuScpOjuMopbr
28Q77CDTA8ZNWDY+CHLSk2GVWHFa5ROqFMbJuz5iBRA5GHyGiZeFwRWuKhMJ3rzi
8G6ErsRZdv6yZopIEg1jO3KL8qpOLJtqt/ciXLujotPj2CLoR8X55qiS4An+IBYs
qNpjkqqRsqZNoyRw1dFAUBIYaZ1QRTZALD1Dyat2by/dI96TSeWmIdGf9AlCYHyJ
tnsBZMJ+mfM3qggmIFWDlbsRS9rci8bGduZnwcdxHM771PP8yNPvkp3n0xslyKdS
26eo4fzuhNiMWL53qOjD2JIyQhxNIp3ADClxWBnOkc6bWxTUMRLgd+EGGpwhIgWa
9SvrXDWQOjnyge/09hZJql7/VAB+zvpC4C3gui0WpHpx00gVxmH4mn0mfAX7UFwB
03lfDJDsdpI06eA8+M5mx2XdJu7uukL6nkD0cA9uH0nTOfQPKhXCz3rccFhcTYRq
n9DkOsS+ofS/VDT4XE1oR9Gf2xm84zydoNt5qk33G9TqoWhVkBR2C3iTm8uUVXfE
vBD9KEs19dFPREhsRMTwAyI4352GHYMsnjpJWYZMYJaFKoemgdT60KXLcCdk+p+v
o9+ER2J/xA7hj6kUw52kN4zl/VQ3rjlXJPrht1WcnZRPyqegNKy/WVTzVqykFgH8
t6B2dgK5clY64jt8mC4Zy+S+LnLX7T3V7QILCIF528UsO/uTIdjfwObtY8LHt3Nm
gCHBphFtVN/SEGzQGTy7mKiINxBZQZQkE+z8FNYlTRSb0cp54DkaqSXO+cyBpevf
NiCLoryu/FT5Us2Uxo1RPOZDwqI2sCGGMevZrxzw9m5m5xXeDmwKXtRnXG5n91BF
Dds4zgtylQcq4Nd5yXiaRBZKyPhVbJUT8JwIu/xQ6oOwm9jb9Dk+3UkP+Kr4GDzB
ZBu74zOVFe7FdAhfVUBqySyJ4WV2D0D/eIdpbRg1aeWCUWCI152gkxVwbkhjf8SG
vPIalgwL0GZvx9tP0DR3Lsv2gJqd8zNnwm8uEOa5cImWBqfCQnXSpqsVyNiVB/U1
viPT5BqZIwae4xmWBlBVd6f1vw4vDu7bk/JoeIJprVCaM6G4l3e2Zkoj1PgFsg+i
o46F8NhySIQ5KVkO7ujH0UWDYhDOa4RevWBJqMmYJzPswkZt6Y9iDjPqmUCHf5to
2JeB6JI5gba0AnYerZknl8REfToBwjxDxLash5fY5PZOo5wm/DoHrycgbYol4tqg
4Hb3c7T5o9vTfYQV8qP7VKiIUu5aWH1rg6G575XgO3yrSttgBY6TBcqJmRvcpXeF
HNVz/n4nuiAYKAVUWhMjdLhDB2mw9z8RZ6Of3DhwafTVwDqzlMVqcLyT8HmjMHMg
kS0f1TkEE/Cu/9hj3p5mqSKyi8vqAbuBtz8ePJ8fcr7V0hQXocWHLHGOdR4o3Ht0
KncqQGBcz89KQwPguDXGdKjjMA6e+ySJWcXGPXXQJIWF40ROVBPvF9I63bFH42oL
eMzu2b5aCy6+Nx0mUW/+c/9HrZHq2ykak+IaL0Axrti8U1cNQy+jUaDCmnL6zJDi
iTSXz0uLWbOZpW8Y0udqcDI9d7buQqdA+Chy6mHQ04J8iVsqUGSOW4fdUpMotIg0
KaanKgLxclZM0tPu1GJII6Ejx/C5EDbRODWswcdvaMR3u4op1QvQ9uYRyTksfv5o
PBOJUwp3JqLQsV745Rztp2rqRIJWStosbv/0ODxsmNQ+5ID4Z0psjfzYKhzmANX9
XTn/9K9IHXSQAz/UpeApQoQJUbGIs7NcGZSWx6lUou/FnRNcJJVQUJnLYLOTbQ1c
0uaSMGG/GAHgZie3XyomBQ1I4skT+q/1QOvpbGZuTmNvH97l/xoVI+74o69RSOef
4eDbj74g7ScCZYL748AxNXDH/VMTJ3h/mGNfM21BCZlvE8S6Ol9c8I+6ehr5+DDN
/RmUIcPJ/y1cwRwe+75oReitxdyYQS3hZ5GRDd6mkhEybnAAQ1/hWHJ1nhkBBdD6
jBQyggMlsm7xiYZbwR3Y+fJJ66qJO8cos0UZnmVHwGztfGki0GIVIOgZUwXacXjy
f+L4v51g7H/bh4xJvFcPiW0oxyhChN46UxEBZtrYIDwv5qD5XFskDR4/N4dhYN7U
SMGIWXsmY2Meez4PVVnFAQJ3Ij3GU6fzeIdvFSDlyNOSW84Fnwc3EtU76cLa2t1e
lfzFgMvQABz0Op67cXIROe95N826uqY+Ygw6ZrVdjVooq0WNMGVgCAuybsHUJCK4
xN4VHsE0DxzyuTNbf7hfyE05/+7YE5Se+bJ62SwSn2nsjxSnOVoXEWfKPkpIAqfr
F4CMLOJTvo/aIG4/ZnPa0SvMkgVHlx+YpUjsDT2joPI3r/UrPIVd+fVFxpDZgMlh
+6wJAoN+ABzkA1ejIW6bnmtHlDgFSSHoVUCPl5CNr5jEfyCzKCrILSWougeVH2F+
hYIMhCzlmbPXWTXRt3hxRabb2kBb2vNY2+n4SCN5o+pQr94NSIatrdLzFORkSQt4
UYFzP4QspGZCEcSDNu8IjpQi5PP0C8jBTjyMSVhLnjnunLQCnCO4rHsj7Tz+1g89
B8DliSOPmJtk7LaTf6E1wea4d44Z3SOev/CRvamx9yLoP1IDvxhY7VmyO227IQAo
tmHQ0fig4ziwYv8PbFR4FCGSkLiSHtJ85GpzRq0izzGD1MlkD25qgNWSk0ucs8Z0
l2TnjGWD27WKj4micUWyF5jCvPCP4KD+B5YHb1ucuXhUl4rr+mr2cCVoK2UXlphq
ggpfcndGT5WwvIMH6qqG3iUJOrQjpmjCOFxKMicnyUJGhFe10wQcZeRtPU61Khml
EGe8gfwKUGUe2yWon09CO8qzPKap9Ves3Ss5GOCpMhhoY2zF3QSZl4HMlLEvFkzi
GM9oA3WWUrBcS+5oz6b4LLs1+XDayhSO9sNn3bU7iSd4AtBjycrYyK/D3UDc9N51
PsoXr7vAFRexoVkVMK6teEmsCCjD7pfAp4sGTIpYbQ5QcpImKCgps8VCRyZAWJKQ
AuWDM0y4qs+pnNQHIlVMqN3g4XjgwxxYzhTHxw/fhNsthysHYYGNJfx3FZAC2xie
ZcoMY/l6BWDd7jfrekk1HQlmLx1s1uELeP0JUZTBbu2UVMKlJxhSmTJ6Ed65/VvO
ZLvpy9QHTvez3zQaLMD3E1nGr4Ci9CwxZ34H540z/rre/Th639oaP+w0upgwwRsn
yt80L9ubcKaxXPOxv+Dylj3MJdqIqgi4pslongCLF2UY7SyPhCckwynw8DxHvXVX
7G7npydJoityu0uhaMrIGZi7vnb8Lkxvn2IWztxxDzdD5+2li8TiB4jZI95MbEV9
KQKosk+5kX3ejGDFadgma0lghM+XuKhWnO+jcoSHlb88OY88HZEAjHmgIYvM7emV
nyR9vDZZTNALcxmHIiozFY18GAj+c/odE5Mtw5LU/ImfdBvEDKJtV4rGcwVxDcqG
X8zbOtUtNyBDE/gEI8FEtnEKNzcHp/eJnraQG9qeMviVDUHGB9i96c5Iv00TYflM
pwlhU0uHYk1Pt++V72uZFk7QMWGM7iRw24u6OaR4nZYhetOXMH7/Fy/ta+LS5f52
6XZeAPBzw1ETopwA+bwuPPdTO4F2i/jv9WH6P/JsmT9dlt/o8CeQPQ0/QBlIGNR1
etTC2B6JhB/LVqkHRJnUpckcV3GyiKspbGK2PyRui7GJqQg1ze6eeVuVoAOXNBI6
kVQVOuZfLzXMXKWCyXIj+eZs2koRaIMU2Drbd9GUQSv28/nDEkbNOSDqhY9l65tq
lJvJNotSx51JMwIXnU480K6u1Vwy24a8K7LU0mJJD7D0EoNPSFSVPjbXN/XX5hSm
cGe1tKyXSfqe8DF82d2VUkN7rM1fdb/HA0A4KXQcUa5o/bYJ3YPiJZ6NLMMF9VPC
fQMVXpqr0gqsUva2s9yrGSTRE3U0Iepo2RO5JWFMmbhXSngA0WGbPdNJ/vZjoKKB
HAUqEWLNP3p+tC/msVXPjSBae+RE78ECjytvrjvJMVKH5sPSvWTzA/lFSDbfq94F
8RTMpy52/JVDioDObGZ2AintYmJ/KzyBXNDqCj8hLOvx3ajMg8OszPYjo7X63wug
ReO3TwfI/+3VuIXigKepMb4gxGnn2H9jynrgtQbK6KxV2pBnA6BoPd6HGDJ5R0I2
BHlJIkXJBnNKpXccR62FVCCiOlxCoxWlhOtaes27qP9F0/ZvA8e6cpJkWyLZVnt1
xBi9fRxzd3QfrXBn1v8G9W45czrH7dygwU9vngkOHPBKfqiKmWPLjj3xW9ThQV1H
hiiQFESJw7ENUB6VJAzJU/K2Q12sodPuVMkECZdULUHqTQXL8SArqnA35/LzECXQ
tCYFO5SaNj8fpI29lMmJbieBVRiuPz/oBUwrw/8kUG6kGrX1xANEw5cdYyN49+pR
6hSIIt2uH6ROFJ4Fknqi0TbM1GcU0C+jbZI2LJl2HMNJZdNaZjcuPtBeXk4dqD9x
FAtjPi2KOouPNc4YPYWaxsCeaRd06VVV6FnwxxcRsNLInAt1rkN32QWjmlKK8WDP
Hp0RUJMMPT+gOdfEq0FV0AkMusqp5BPmpMcq9Nw5GQJQwAiWPpqVvO0cmO3FfLhp
JgWroPNNVLMOknBgHECuFjMBpmtpnHy1ghbAJBxNghTOqKeqBHeZ3c9b0eYty5lJ
13GmgoFGq/+D8wrh2GuKJ7Yihgm0DPzhYHepBHNpqtVtNghtfOi/l/pE1yQyGdPk
LDSD0NSIfjpsNUGZ6XeUT4oeRSAxlU6VEpsEGU3u2oiwlRyng04QZnwIoqtlVHWJ
jc/Wf6i+5U9wr+LEUxXjb7tEXAFoldlXGldMgdLkIuGyKPCTsTwNUOs8OOgzAJ/k
KahggyktTfhhn+KJZgxLhnk9/T419k4ESEYceLzwL3UzwzimkuFkiLbwLIEwtQw1
sMfFMiy/qLzlvBGX/uscWxl0zQoBI/DGPbkpREmKnsBa6dl2N72gn936XveGNhPz
R2kRJ9giqUJqXyM3O4Ztl3KS5zjR5re6013+kJ8dryZBcuRcJSudgPWz+J+qF83F
7/nJTw0Dk98l8zurFGawF5gtNsqK7/GwOkD33U6V/uL3rpwQC2OBLhODLpWCRxlb
rptmRGqVZT8sam8tLDXhquQMk/z9lqWzBFwFQLRY7+tPEAMNMuA4a+Ql4DljeG5R
uhRMOwzOVKLfhP/6hgtImcaYPoYaqMLFZZSDTlC7noCHLVGN5FcivDF6cOlYjjca
MNG+dzfvG4ntx2E0wPhNrHsCAqdPIleV91Nxw1z/4Bqb0cgfP2g7oo4jzQDpgqcW
LRYQlbLR1JWjJuZwM/gS7CU7CauZIO3si5dVUfx4Qpw7hqLJ3W9VJqqkAigM5DSm
nFqKwgVrwSK/UVa+rBIKiu9d3Nowoem3bhYglpXc5pHCkKSfpGwGA+dP1OJH1fyk
ym8f4fG42c+bpy1/gfEU7VRRF+bitJKl7kB2Whg92xQY6ajVVXVAizv+D2idFuY7
+DFzS+F6xDsqgA719PsGdYWGHvL94QSkcZUZrATWIqms4VR8u4lCcV/zyPJPJquN
NFSChEXW6ugWPAWTYZN4MlL0+h/yG0+rp+eG59xZZrXn9NV89Zyrk0OQI+t1x7uO
f/TV1IQIEEuvaMGjmYXX9WQK9nXF1AKa9r27fHp63A+VMFPIlCQLfM1R6eAg1UlE
i0hf2nk06zijGtgqNs1EAvnz7X2Tp4pkP0lsJYbKB4/I6j/nchMWcHIjGjmJvW0y
26Vcqetm4X9yV2ET7mDS+YLnMwBxHgilnDj0Nx1tA8Xm5vHJdkej+iBEXCf/ar2P
pKU0i4FWOJlelZgpiVAsaiOU6ml7vZYtKdd3/dTTUzURlDfJ8/xBkElVgd0skG7H
VfuFXHQ40oiiWF1ysU7Nyzm0r232b/vk2V73yqasRi6nxzcGBidJiCGlaSbatByV
JfR9E4Pocp8PmPjnIiwE7TZoHew0GS1lp32XMhKlbiiD1GxxD00XnXEEQPipzyVD
CZZSOUlEeJJr3Iz5jMtrYim7dZR42IB2+K+gbYLQNuM/7ll9/t6zaw2MpHw/gcS8
2f2dfbOhATmbbLagDUNaJtw41oG9dlO3mbFxaW3Bgf3Ycxgn8s6SpBtokiT7e4Zf
u+PcA5S3fXMqbfW6vfeODSx5E4mwwkG9/3eqR1GkaosPxuu2jLJzBOJ4rv2W3pGV
dAtELYkAOGS1zwUVVbUX2d6BX7CukL0e48EAJvs6pMf6dsZJXm4aNVoRZ2KXUW0W
5jMlCusqpmMcdznnYXp2fGQOkr5AejGIzu3gc8Q0Hpon7QISsWU8wQOAEAN9n1W+
0GsYfSnAjrBHtN1YzFh+gk7535hN0eitEB1rEsqZBnytrZT7uwr+Na5BJyn0T2Gf
aOAa76EurDCA3boXgBe7i87HaDYXkKYY4XP+wNcWqb3LF1RFo7vsEoDHdrxIKIsj
zAc6KtJp5hh2WWABx1qHFQpJQfq1YfvX4o2PZSVr6Ur9czLRzlQsDmJdjccJonnf
H6DbuVTAtu/HasQqoTa+k7TnoPEB/4qxseMps2hXxSWPJaYTvbhafEj0h/ajxpKF
uVv7uIB+MMTye6lTaT6dj+O4IUvf0Q6iTqiPKo3VEfAmaasmjJkcTCsMzNJp8ejU
xwzagih2AiG6qF4JKRh2yE4bKoQJWDgGyB/lBOswrO3Bo/ZO/HQD2G1ejRUI4zk7
sDA4S/ePdgA72JVXC+/xoIqWGPzNpc3Pa7qQ/amxgscWrkrWLQH6op3MBcOcumyT
W051ANggH5cUHFomsGIiD99fA4Iy1kNVs05HERQBUELlBK+v/bhGEHGHHkBhRs0M
E4n7OSn410kgCXSm3rWDM3RB9+DwALL8fv5hzF+0LoKS4V8Pp5lEnTxPAn+5FKt9
bt27kxnygAnG48Q4O7RGzuVC7RuCPGFxDaCSfZTtTg4tdOdIGVsJHqlPWntZCgWZ
H0N7RPsUdhr5I8s+/3CBjtffCy+by/QPAua08YEif98x8yjip4qGbewXPwogaim9
R1zkhUH7VvnUGcUjL7sHX+Y4DfALTl/mtiXt/+3kHv+aakC4kCw3iNq8/PDfv5X0
knI5VjfzE3UrMAHbPWnj+Z+tvErzYeBBjz1PGUvpqYteg9dvXlLNVve2RhUKepav
I0HNMu/INukRmBB731CXc6kIUpd38Q0lMGtcAAGHy0Ub7xxmPOBquokfFJvrZJgM
K9+k94Qa7Pobhs1bmhiLtgR2LsSwXLdup8eNPtLhSgaaNUazqYO/n32wCtt725D+
Wb6ybJ4AjxwiOwvek7NAbqDw4DrR8iPjlcV6XQYC3fXNPEZldrseQlWrTDsinPPq
MpCsdHV/iF4RNVcI9bSgbSEz9xE/dnapfU6bChu8owwtV9dwkpHZYGgXJNj5f5fD
IMfZlPkLashPtm1f8KJ0oF7SiXgXTy2F9qXN44hbMwWYBF+gpQEC5LDxb1i3DTqp
gjVitVXK16utIFYODJ6bviJsSDuGNvH3CsTx6QWtJxrKwTzlLQQl0OiHqaE9TLeW
Q73MdK3N5PYlrDQotPZgZ5f5DLhaZgDxd0oPoKXWFiOcK2JrcPgLlrPWQA1HdxZR
ojFWOgGgj3cR9R7jjMZE2U/TZzUl4YXcLxUS1ViUgBWLeGEjw3jY9/fxoPbNPj93
E0GdfPjjAHHq/vdN1CNM2IC6q+DZ2VTeHVtZCgcq3MB54Y6Wo8L66ItEzW1Pa5IY
U9huOx+FoYXkJEqOLQW8VhX9MMvfTSvhYoiZqlm53RrenDcqb6icttVyLQOXAxo4
h38FDwiE3g2t7li72atK60naKmYh7yhDp9LHeOwmHwHTQ1X8lgBsW0hCQyR5aq79
nM6Wi0EZMo+R9o96CeDK4w+jEUejDsFPzPONjwg8kCKI/p8jjnMpnbCR0oSHMUrw
E0xhq58ETF2TVK+6GoU1G3yFhCUO63IDgz5eV963nVh+hlxf39MOirfnLj9SDcao
RUMfKoksrJTWBwOBhiMvbZ203FI8LGgMXdzrYnmGW2mr4/cIcLuE1/OAoGvvxsZn
j2Ntq6TZ8UaTWOGgQFO1LMlI+L6TMIWU4qV6EKVRlbkY/nZDjKlTIq13z3ve5sDZ
MT1kj+1II/ZsyVvNrFq3TExWC0FpiAbvOyZjq2G6plCyy+H2hnGeYvPLj0rfNnIh
XXwTSTzgxD9VC1s+PngIG+Iq7lQuHozq4ot87qEBEpR5LSvOVW5X/SMLbzbyc7cx
kkuojq0VKJIgaEjHNZDTp4Uvcrtmy7FULdf2i4kTTIR5DHxdvs0ko9+7oxKJa27f
hr/xklSmVCseDRlIG6Hn9N6Jsd6NzgHd5pth70LInswb8V0RmKy6K1VCSbmaNFov
jj0QGCd+i3OBfo/fbqgokEAGZehXeuJvuF9rScpTo8YBsjmEUYrlSc+Sba+XgDHl
1N8wlJrKLjKXnIot1L3y84TTOcry1A2/DC+G7TzEU0C2q9wFtZ/4h1uKZIeTftUv
mMvinRHCwIryLnF6ZOyhp6uvP/oEQsQOSoQ3hDZnaqcpoc3XpMsXHuCZSjeQRLcR
sHBwbe8vPztWp8GRb0KYSZTGW0A16t7RU/U8UxN+s0jqOYeubhWg4dfevKRYDux5
lQgb7qTZG1LWl8JdlGMFq4NSIqF9LX3wi9Lp8tri+ziMlT/vSg1cRappYQHWfEVw
yt7Q6L/Z6Pf4q9b9QuLnteVV3PG6dLLDB95jtQm+mFo8IHxenNC85+IEJHAJ5p2y
qBM5jwGxqhin8+ydRfJUrlwzK4TGG8hHO0buMqfIYhqkh0cn6SoxaCBn3nM1W2Ae
t1L2Qw0x2JrRB2pkh/KIBqYDSoXH1dK9rIYNeL0lOLCN1G3v/CQ4DuC2mffJk+wA
ZqQyisW4U/Fiaxqvi3oDtH8/V05s+qn6Mt28rNdF1GMY5o8NiIbTgwMT9O0jYEMR
bX/uzI+Oc4J+D4TO8jL8HpHLOb3UKeWcIE16x+tS7rfVakYYPsXyjrPwtxJY1WaL
8YD3MyFLDvK1IQyzcgr6IzGYS2RiVHU8A9Y3j4Fa08BDeIRlRkKPNWd4EZRH49hQ
cKg7Pe6YUVytPKGKjOsS7vwMt1rutZWGqT6Mu4Hj9idrB9YriEPhTy5GCc3fmwqR
B1MvXAi/xWIhJNqnqrhC/fROtkPIYlK4mRFDG3lUJXfGtDwmeqv8HgagPp11Nx7b
+PjilHFYvE+1KIUBYr96vCnEAtPJ6quASfKk7xk8ndvT7LdyICDnPH+xEesSJmJA
+dH3EYQLGTf69koBW5Yk6tulBa8qAaLSRV0lubX/+5GfgmOBB33mcyXCZO5AucUA
mqBK9MguzI61PyX+DrYMDAWSyX4UWTGVh88cEagdxOOe3blCzFoxx0j5m2eqDMkv
6Y5h93YvQLohYYLImVIRI4TMcNwLtxPnONvSgpRj3p22qclSNHwS3azrQ4F6kW3p
jXk9KyuQ9X9AE0ktsRr9GbQpynlFZmjxhqmIURQKJGkaz2rHBmD59lCa/OSytj0d
tCMKJ7lEf7EN2dQYABRcHjGr2J985XhasuWgmDYn3PBns/3QShSAlvwBS4ST2veD
ekmHZJNmgunHmrNuA5EekMPcB2ban3XMGeOSI2mn12veRS2ZhVe2myJPnI81fFbE
PTTNIIWmAtcCNLRwkWZM9CrT9QX9Fj8OYOU9zsmmcmoZVzjNy3g8Zyq80e0Ke5Ww
rk8WXS/QtDWxLm46FRfx3FzFzt8e7H8Kbrv+fHOyZbLPeYiJlKLsM4mRaIOTx4Pp
zpuzCCCjODEgxEzPt589YcvMu8/7UM81CuYKl8mF2jzQbpzbLdocowfiVjDDBZSj
qHYTLUYnfSYqYhLhChBf5F7e0htVjSNvDjODqU+1W6rMDWfI6NG4TZMopjhTnQHh
3APmTM2injlWn4PIxYzTus7FYMjvOpQBzDa3h3cu70wjr8p189tKBym/i+QTNphn
S46HCpq8+Uv/vuemWVWIu7bUZh2gRNmfPBjOW1ipgN0CjYWrNGtPKF28XzjocY9I
XGmL5FlpA2RwZPJDMqcJ1sWlqkV73fAg1HxnXNQR1KCVlVwY3k7i/pj+ZVz7aXLi
S2a/3SQvHwk2UIXC1i2k5oNJATvR9/5FF1BWKb5OP38A8vA5dh8eYQDimAw/ocHt
bZO8bkxGWv/2hmWVO0758dJInzEfUuvS9rAk7kzJ4TIjqLlIccnxyyRY39OP4IiC
XucY9k0BppSmzPWOsOIeeJ1L/ElXBoTdjOnIYK0tl287aMSeNiedID68JZ5Meg/a
SekGoiSH4gULzmddc9iIPiaJMQ3eouNIZFmRzvci6f5AvmYphN+UJ+5+Rnal9BR+
Dqet//KQjzN12t7xksrVYW9tJoJXI1NcTZV78v8RCePC1eL+sYEsJwwUoS7cCDRt
aUlKYBvyrPmhsUIv6jiBBbT/xhJW89Xv5s+YiYLpRSP/4xCzHonBz/dVxt8z9lFH
kRYaFRHniLhGDg66h233yZ51jbtf5BdbxYbJMnvkWa/+yb9zYEX9z0a5nwBTJXUM
1apt3/evqsLbolCyYwjyYTg1Df78kDjQXS6V4szUBfSaGwGjEKjZE8IUcoCMlu3W
r5bKF74+2MkOTk8xQx4Vw4l1gC5AaCCTSUSIy3d8CH1Z6JDD7UiuLwEAF1X9GYyB
i/dVBbDqwrRlvNlKjfBzzLT0ycUDXLzFYPgWznxxU9+405bOdDazvcfF0NGIRPZ9
c4h9KIeMFbT2ig4kZLiuNj8EdM6xtZOeOSLHNyeFQlSeLklg4+zdP/MYskeynF4H
jKMxCc3GMJcxfigdxvxJOHnviAt9nkPC0p3aoVqCYZgKXeGhTkemECLRhBtPi0Qp
RXBBYCyL3FJFHJ5lRIiUihRj44ir8asji+uCSF0elc8kNMzpdrymEaCy0HsvQ6DL
iibJZ2i9VIAZL/cwGFa5z/78nI/8AMP/zdw36n2f9zlflkqbCSlhRyra5LOHbZ9k
BCNDpfYyW/Y55VliKdy0oDyiO1XfABgl/fi2KOviEYFLE9RgRGuhG+fXhV6KAemO
HJz/x4AEdb1crsl9SePLluKauwCP/fKyIO522Lpjp0U4WK8sUKRPXh4G4yjkuC9z
Os+hbzwLgtsfgYxKaMILsNQ8E+wdOjW5vgYld/aFSx4+hzIDfc5ii5e8FQnEm5IC
nqztD/x7JYR7Q2nJ/roYnTt6Lct2thHprn08Fuoun9pY78c39i0iZAv2EuyP9YWn
46VLFdJS+E5Wxsn2J6eYzS9xVcqWZjogdpiWcyMKRCvXWCy9pVTdObI3XOKGQ0Jr
TjQ2ge3jonMV68HtfO0s+/cq1yV4/RTdGvbG1UVq0aIS5O77Oit44nZOayHXJT1w
uynY6rAu+/MdJ1UckJNZ5eK4bPUMhAgrLb4c6uG6kC2otXwyNWBBwOR0dcxl/RJQ
`protect END_PROTECTED
