`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qdOiJoQlrVCK5BV3k8oiE3ZHK8kshjSRpAJICq8IZEkg37ggp0d/0ebg4XawcKxE
HwQN5MkQAUglsETPEZsJtFABXjYHI09WjXP/FQiU3rdNm4H+vCvJTAwUrL/GE7sZ
ihoyanGAuiJ8Ix62mQnHb2uGxINck8nmT2jjwjngxGI=
`protect END_PROTECTED
