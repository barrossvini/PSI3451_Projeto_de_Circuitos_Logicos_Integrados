`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y50nJXLzh+hDItDtiuwCRfwk8jvuafpMvM6DR+mxL215klTOAAl1ZY4fZT6p3/iS
STPFjcyENTl4lYpiM15hhnx1m1+WOEj5W2qrqNZuhPoo6ID0rprSMCq0ysBxbt/3
QaDg0FD80Adbf3rFr4ZukpeXr/u3t5NesOsf44Bry1jAsMO6HHWZ1GRvJlhYnyhQ
1v2LPZQuTu3ACkhfrPIHHXka4ADl+hKcT5PxB3Cn9y2eUgcAbEHDy/rXh0KU0SW/
cizdZBkaXYnYphmAXXqDIy9MxB89SH2EHcajTmOAiBuPrpyx2BYitHe1UOn1w7nN
NzlWH8r8ZyYRkymFS/g6SXAsJOWLneUQysuo90CDHMHwfXZVAiwFS66IAfIppfUd
1UXDZW5IZkXA+fVfy3brV22aTYwETcoeVZVfVtMHUXhud1tOIPW/lvt0L17Q0Q7T
q8X9C4/rkYiVXgTxLoMD0x1DFZunlIdQ75v5CzCcoyq3b6+U1asxE7AVtFEgOCU6
aDRL6RBWfYzHSwdsj2ooeNs9PgYWZK4E8itCje6lnQYLuA/8/Qu6mTRaxqhFv/dJ
sDpnPhI4pob6swtvNb+1uqI7otngWvoVCCbNFvNMW/ngIyNGxL7O6hxb+sKdUfYA
9r0QMfKKwtIQg6YAvrhKW0pXecItHgrkHtm9kJiA2PZGzg43gu0ZeuoZofSPiWB6
9h+3emQIfagCelHR+pJC3abhr9yt0yzYkQopovM1Uo+C3FY5YRmQ20mjT4xJi+JL
dQBlWmgfM5gfuNDCCEOHrsmggiPt8L4c2/5MRTzYi1bCiIX1SVhy87fuXd/q0yHp
EYBhpgBbawveQMpR76sg8J/PSOS32eDlXzwKHPQNXDvbtH4o24f6Y/Fnbg7r4Gue
oJnEEvMFrcSGP0SR9uL3B2irg3nTS8dTFb4eMGGUniQ7XcIHiKDIoGBwsWgrUq/l
wLBZmu7J4XV9XYvsGJeafE4hMGD/G0o4OjF/Pbn7sSrSNizAxsaGm/xPN8SmUe41
PimZH8fuRYHTrwJZbFoie6dByzX/u/lmjDQRO+ySFWsR//IhQ87MxGbMtpovZul9
V7r4+SWyPoGHa1uW5+NxoJNlLONqvxL6R29U0ocvlUYAZZ5c+hNnI/uBYp1GKB6V
XFn3z8dVYMnTkUiUvRtlzgPDZyu/Ky9lKFkxMqOIXb1qhMNcktCc2WOWNcl8DXuR
Ufxn/y6MCljJpRUPlfbbQObCkuH+9fdWz26PMl5FbBbhw18avYHGdIE7Gpd7HVeN
zLkwPxPV98umZrx2XvUDPahesErMksSdDSla1zHRKpIxhB4+zoegqIWUqQSwA1EA
Cy63AUxH7Ox38JhX1+nJ+lN0cm+S9IoxgNSv56FKUSpLdv3zshrZKA2+VjFYbcfL
QD0hXqREtZNQhARczcuAwfe9/304sLiE+Vn/ZpH9M+FMVKQDuuCUwAeHGth6f7T4
nQS37eK1OUUxZZX/d8WH8G0q+hzICV4FLvyUOG2/MsCjCzh1Ld2eAJFzE2j1bzSm
dxxPWbYDamV1V9N2v3qlIKD63w9kuOJv0m/SY85zKVGl7DO3guLQ/Xo6P5Sj37lG
/JsoWdGBmeWbvd4nP22n6w==
`protect END_PROTECTED
