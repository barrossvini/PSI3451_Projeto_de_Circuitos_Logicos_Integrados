`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xeCVloZQYbr33sCcQDTzkYcNQ8GNdOl2LFHPM3ITvZtCpx2XH4qHg9hH1J8IsCZu
pg8ZBHP8Vy4N0VHdPZGUQztsD9kqplGuUr3VAj6Oo2Fq+psEBS98AdmaxgnuTbYo
LPcJSAHfaQVGfnN6idJMbxF6iMyjZWPPz3/XqcErEf+oCN7axsYAW/C8DQ6A0d44
UzRB645ExTtL0f40HHrhdGEBp3PO2Pg3aums16k+IWoeL/hzeNnYZryV6CdV+H4F
s+hogyFFFk2VI8W4+b2+TUrGWNlLvtFzTrNKReHb4vl0mWr4ue9tOkzfOu3s8Ew0
Nknk7enAvo6I0uPs9nGgMYpoZemkHQl623os1od5PKXzOCVMb9NUY9tjxgxxF3r1
CA8DkH/tdW5YB3QdBqRHxUsBbBwXllRRlSLwkdDvFx86fPJBveKAHgHyz3doJ6s8
DobxOp/DXt0XWCKS3fBhpKiXYaoTjs+gNBlGmsxDoGDgKRBtuQQ1gmuuNfq9yGGt
M10sYX3TJQKL4kUHgC2Z8E9zOvaFzgXBsZpoyxX8dNaVulDGp9EWqEIfi/ASDjjw
CLlbaPLDyZFjS5rHnwZzfTyu3zxb8PutJmmQr8VeftUAyI9taBLHsp8eZyMPITXs
d9F0LIJhcn2b4rhqyZh4uSWu6bghqYddNnimwXqkE4XS9hONUaw9Daj+ziRugO8+
`protect END_PROTECTED
