`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dWhGZ5ARQDuocbmowc+/551BL8FATOkp6faYBXPv6hKq2oCHy5Sj684fDxGlM8zL
yX+LQlczuRnksQmSuWUOYkW6sRIMmMmCVN6AWC5fOWT/KJBSvypsl721EHZdwiGP
pBu0VTAqNGoWG2EiNmmQgu0a/EF5RN9Fu5+dxvUss9O5IKP/sXkccBfRs/lzaSZv
/YpAQBFL2cBWXB0ZzN95EFd4vraIFB08WKwx3BFuNaA1SLZG2NQ5/GJSVi7MptNt
mjJb+2mmRbsqZGCgY6GeMuufZUtd0IyHcVwP5kc60v3kZUWAy+Vdmy82WCJ6ki2o
rCYw5FgRVdkfNL58o70N0F/6B/x/gtBTgU3cDbeRS0LO5hPy29EQoGn4AwC8uL+c
1ZfDq8s070okXebaUbxA3Kc8lx0ycvrdFbWeIKQoum1NdEtkMkRpfzUQORAe5vJs
tydJxKejZw9cKzDuLHU9IWmHyfNrqYBoSXOYoRrSWfdJL9dAhSeXc+Ukd9W5oFC8
luEHyCulMNVVcK2ZsCRmyUGm1y4+Kst4s/tJsMypypkmP/eaU1akX5e07TMXwffO
Er4jUB++dWkEeamGoQAgBlY4NYD7eeKdp7zybZs+UO+tswvKNIRfZSJmenm1BA28
5N7865Y1mpgtmLrHO7IL1+DEWS8sHifCcOsdX13fjPHe9Xp+j1qykXsI5NOl7sCv
Qid6mJHmoXdHKno3JiTZbENoV9cumv42wSMJ31AwSLB8ktSFylyN0cBnzcsowZD0
6/hz+mXt72JfMxcbLTpjjpcuA4sv7dNNGyep4b9DIGxLkt54rStGrAC+yJBYfn/B
M09Kw7etpOBx0f3cULs9+9PfdjLsQrPRLgKaubfTH5bADHk+Ek9TJx7gVrMelKxi
VodvOduPJQyx3XCUe5LcG4q/ByPtmfbfSpQ84TXJnzduibGm8qAOil1PY6bxfA13
smAJuDeG19J1zHxUvmH9gw7oGxaIcIVaWshxVw2geHCbRKxp1goMcNxLiR0hxR2V
dOciEvXgLgVrrEm4BUCAblbXCESk20HgsmxEHMdNlNUdfQTyt1/q8TU8OpmbtXUv
W5Veg0s9UgsV7UJl7wXh3amJ4N4t5hH+vsSilMNjH6kgfi4CI5nTOgYhIU8dbLB6
l+HYf1i4B/pElzao5edKYeJpuyz8ZGjun9NH2mgOKoKMuK1yMPwd4Yd8Qujtd53R
BMHnTbEfxJkMcNjCGxRh0BZ1QfJ9O0d90fDKh1yKbniQq0srYiL+gk5BzTS04YhO
Y0kX8FhEmKetAsRx11H+N5hp0soPy/Yoxm+mtjRJiF9BDfESoVYzIx00YdBjcX11
NTqtHgSZYY24Db5Lv+dbEA+M7FIo5fv5gShMr+4pDv2naOibzqklCjnwx414IO6+
+2uByT+d9xoqhBn5HRKNkN85Eweio+xpWkchBKQYVbtdp2WTdxEqWKd2BtVPjGle
WQ9xg8MbGIm5+KXaYEfT8pkvyskCPnMVvpIYIkO7hUeKs+pO9RDn5dM96YhYGpNA
RTUkcywzUpXc4s1w2WC8Cu3bfEb5ZTaQZ4n4OS47mHFQ6TojyNrivxhkHHoqS9rz
XzRWA8W7PMdZ8nLgzzjH/ZoLIbkH1/x4MZfOkb/6IcV1fHuadj/zr6wsEdzjxL8e
JdJ7tOCAeWuilRvkSqO/MeTzhr/4lsHwi7urxg5bFu6G/k6hgThCl2o5P2dEQPWz
/jWpqpra49MYuKz7b88LHb0IJqjLYMMNjyAG3iMWmJs91fM5j0lp6TjK+dZ+fZbA
91N3wTISP5qCgUeX87VxVcmszqS54vD7dbkzZ2Jvo9iHNyF7y0E2qNKbeS4ikv64
iTkM9L49if3cVZhQeM4sbfrI3R3R0TfPoGeu1/y4fYmjvFZ7LfNyQ62qJh2p8x2d
4ASY0rnQqpA8ATDMtwDvnZSuv+1Dme9RUY7wTKzZ4aVZvSSPVR4Xy8Ei2xIWdZIy
mRmycr9hXRgBAcWbKJUPkyY1TVRzpWxOYc/hJUJb7K/7x6oow80pLdZB2ANZ7/qq
GM47QOrnutkdPqSk/CsYq7eR3OgLlGPVAOharaOKtn4sHwQMVcHddNZuDfdgQsnN
X2rkY+Xz/dhD5TGtXxnhWHUrDcc/cXW37hlWwtXvDLj/UfJTU9GiUtQUV+3pwwNM
yqY4JBtkcSqGcDj4B2bGXzdBhxIluya9r9IbAE9LQUU3lLLHFAMD2JgmhhjKIeBf
R8YJwXrxGBKdSYLr76Q4/G2bzORqXaiDm4ElPc7XVr9hx2l5aTMaCNFq9ZxvOqzk
fztROXDk4K+h3FjiM3h5DqCOOFLewKDWXrfs/H3T+L+U+it4Pg/Ia5TPBCkCSZZt
6Qj6AmW99CbdNcrBxS6tkKB8Ju1pTaW0wriA264NwC42lwUJyZSVHsw5qQGYrX2B
YjOtRF78TowL/1RETVwagA5KU2XxlmpVtbJ6Xm+637gXDjO6xfy82QOpADRFLt+K
gBU0NF+/RYImiD9jCceAYOfUs/9YSF5SpbWh/ArHndz5MyPB/w+lDUbX16ww9gd7
fmuZet/Vgr8roK2dzsmxNmp9/D3vCJh5VzoBomy1UePrOjLc1orGsV4az+lAmhMz
xtSVBsYmWe/CPpUWqQ2Kg9JOvJpyVUDV5UiaYb2fBWAFc0g6mHMMKi02SMR6pTM9
LOHSRFHIV0DOdXVehd030ua0HgBItaCfZU2T1Y0oj6/Dl7V5hn4y0WFz+tuuzW7z
lsHOnukd95cRsTp6icfixcAoRvNXxOitjUENp4W/UJh09cIbOuWwzMQD07QAbm/O
rhdF+9PORYnuINCoNk95grH5cFEuzDI/uCWHgsBNErDyLalWZFZndJENtJSE/19L
16I1Smh3Cq7pzuR6B9tTqc9kM6m32keUtApoctzZXIgPv66dD9HxTZVGruqI9mLQ
N3rp3sUlqXnzpHTR9Dfl2G0OB0nS/X0MsoSKYwB7ZC3K5vCJwBrx+rcFW+hYAbZf
zhYQ11V0adh8wJqKC196KyTJ6NptUDjErTDiHXWE6yIQs8TGGeQX7U4XXv6v3r/A
cF4TwSOYyLNQjCYi3SUJfne4mv9YjMRwbl9+5jLe6UDrRuvn7CKz5hkKOHDse2TE
vm9wBNQ/IxHulXaxseQyb1IYX4mDPOPMwxglKTHwaBqhDtkIpzZ2eYOsWxV/epbF
HEvFFeYumbGaW32RnF50vak1lB4DTw/IDKR8uQgBJj0lmuLB70ggyYdfl4natxVP
UZEYh7zTMf73AVRiZb5DG2g/iVoySGEPVMbqcS2HtGYsErDXR5XgV5kFmrPBahzq
WQesqRG7XoD2MbOdoXmXH/pq37w4LjQozlJ2cMlIMwSHAtxHW4Zq/7TxMwTnNh/3
HlDcJmEm2piegwaCRxsmfXMFOFxiXx0mh4ee9h2wyprhHUthxu2wIFd3hL9z3d8L
wwTKLWaPV+XiRW89W0apjx1oMXUgflr3NOQqVV5Ix5qqRGL1WztBrmZNZHFKHBJ6
2KXba/3MGA3cEFpCDYUXXmbyUckV90Tv6QXZM/BoKANKbECOJpe2T4vhwnXIfB9v
vlpxTifwcu14hujaNDrlawtdUTLuamZS2Eb5L+WIppSkNotV1IcLx9V8pcJ2Fdz9
kZT+pm7HiMFUSZpPU61FJTdFwljMsw0x53g46NpWh5xCsf4FmWCVMBscq1/j/8tm
1SRqW65Yo2dUopAlRi7sk9Fiik4Zt4dViwFsmuxPW5FxQqybH7rGrvcbxfHEaw2d
tCaiFtqdv3TJu1O/0yxokfqi45zcKYJ5T8BVHK1cZkkNRI/S8aBMHbsEtrt7ZPgD
iA8Sk9SWeEuKd8W2/S0hMJTP/IGhBhvkHZL/C3fyQ8CZ4SWbuKyfJgQKf8hjrbpB
hiKIpHzoa4IZJrQf1hm9hUhE48hZFrRG90ZoytlxtUs3fC1Zux5Xdm2Tjay7hO7v
v1ZHxGHvJl1AjfB+MvcD9XDrZnYR2xrzHqmtmB3+oE3jPReqB3dSdiNsbEafdDYc
EGZe37Jfb9jl4vkPueaudx3GXZ+4dtD1T7HQsfkRiZv53LTii7K9Xp9YtwtOTn1o
QzhCJS1e3IQlFGxG5GSOEtUY0PY0XYqOdvp9yhoCoz1TEqJy88SQMv7MzAreXB/G
0WOej9deX2hXJNOeDF+aWIdOokoa81KQCNn0+HWnk0Je5PE8X4SyenYB817pg4nR
fNZ0djUvilumwEjROrRY7+rYx3vlOtPDkLo6bPbVoDRQUbMJo3rmDN+3PofD9OK9
R421vcBmPqTq0zdt65jDStgkThgdmYm6JFUxIfU60EcCzzwrg8Vc7pZBo7w5TwUD
OsjQE1UiNUFFrtmdi9ctxr0225bBsspOoT9SnICHsR+WCfMacK4U40fezC0TctAi
BaT+nsTdRknBD9lRfYxdTs2RFYD9UcEaWQHEqu6NhnkWejvFKCW16vbYTD9CQshc
Mw6P2Jc9ktJl+/eHyaxM+hp6uU41rNpZqJawp/qMmpD4SlyrPbz7Yli1kKa+ORc+
2GMqfSbWn1L2jkGwLHEhITo/+tIElJtUl+SqFUrpYK3XLhN1kgRLq/Pwj2LMgTra
L0wRfQ7dEO5Yre1ym5Xwb05bp/m0sE5A8fu5qtGcShAsghPPEkLhLXt1YFTdbcGT
VDR/fqxGfjJoxUsv4b6/CCyO9OZ4lzqBneGhiKpJIl6xkkxHdXgJCGs5Ochla34H
8+H/9Mior65j1JQ/zfSQiVN5dQ7C6W2nHc1T8JF5AidDpWxYMXuxd3qDaPo11Elj
vvi375bAIKlSetXQ9l8DedDjE1O6ahMuIv0IAxH5IpvTSvg/zDN/E/SLmlhWMS5t
iZhXtsUiKzDuZ7gn6cyjZqf5bwKxOwzgiHg4L8hALL8nZFlHlz2XMI8y/TDIScvF
4Vz4nFhQuD/j0Vq0ew6oHK3XxQsf+YQwEZBO47woDT4n1bj/s0WoC6umo5aTdzIb
O8c4GGqbqcu+mOtQpUbuHiHvrUHdJX4GKKB6/i1TTT99Exzq1oRVgSOamNnkA+Pf
TVZKOc/t8Ss1m3qSmDC9cFgptqquNZrNf1oroHHkao1ebflULolNMzJlGVS5Pp0f
1yHVH2L6kW99WucKEU46XqX4FJJb2VOq5mFc8imI/B9PQzexrCZ52DLQicraU/yc
MFxiCJnJelTrng6QgwmZu/ImWHksGqO4ebb9sGiVp/cwDtxVA3bGaRsNS9C1SNQR
3fCt6qGe/83bVzC688GsKLA7Sz+5susvDD7wlY5rhV1wRDnQ+EsOT2WM1YBgdPI4
fM9AUTEo21Eu8eKIm9rdHKQAVzSWt8kpYPQceWuQEEzx5SSKNfMDqwIjBsGDIPcp
iHhq+eeCK3XoJB3Z4rEKu4uRETn/IBEv7KC43ymx23HAsqzGdGCpPfubFlKxVET6
MJjv3bRNdQYHHco4MnCXC1GsgoD8zK5ThCGzpTozNvip5+pAT3pdl09TFCtXTf8L
FZIgSS7dgd9STCVmzsvzbbiARghJozBvzOP/Q0tXyWMCAlAVrye0GmyRgVBnjtlh
Av55x3MjrhcyO1erz2Hif+nUhSOm22zr1meBdQsnV8i2fbuQSskFkh4LBPa0NjBe
ckOw743txpseeVlG1ANkcP0aGFcngwlyaw73Cq0Aa928MTezFp9PTY8ac3p2bRxZ
5tm1t4ozq5sEuWBKmGslW4dQaIfsHkLT6xn6fwkb4Q4B3hMz3DZK4YP6G8cpzs6p
hrOnLiAWqJdINZRyz0JTiGnieETKRpN48igfQ1e9qgQaNozEej3lOnUwymGhBi9Y
AKI2bp31mKmyiy0s4cRSujEEa9yc2RSId9A/XD1vnvpoRirjqlqJg+qy0y0xQJmR
ZT430IX0nGXH3vTQKt/4SO72aTA8fJ/Z2pLCEiYRZhz7IBXjYBUiH3mkrXQF36NL
KJGDUKoTVoBsQLXLhvst+M4RVTZz2SMFUMdS6sZItCzIxVQZidn080pbqciqRVNk
rjhv2AkNcEpWEXvc081Ho8S23jyTwhF/TdsbC3Ok3Vl2yqi65jMJ2Cl4U6prBKIK
M/KYiamBKJd2WaC7JejNyDxxXOCIeDF/v4rJtlwiAo8GGCDGa+DCsma9S6iOLCPQ
cEolJzSFu3KTgIbbg9DL8UYgGTPhXIy9AFj2lBNI1uSvamZTw1SWhQm1yNMbPXmK
IGTr6mB7zpdQAsAl70LW9zW+ljoB7EAwch7mmn6+mpgj591zxK61IfY7gLJHv3wJ
nI8K1dFhHT1TjW2YOvs+tKJsCPrLzj7IMO8uvlbAh4bwy8faev2fppVrhVKiPt8n
1DDQIGleEYHeHRi3icPCIJhDM6BzNGL4d8HWL8LWeHA+zhdmERk0nwRRslhIE1gj
8No9NIs9RwCuXAb4BMrXti/R418ILyAa/igj7CR9xyiX7v/6TOJEAfKpJaSpLtF3
YqBzAT1mmt5DgG7XgdN+ZSLvpUYnlryl9lE1s+AzBnK8en5AV4xBDnSfqEgnwhOA
JVd/m+RyR5ay0xMMHMrYapRV1oq2uWvvTBhj1fcbOuYAqN1qWtoX7tn1i6M7csTU
BbVMgnleqRGZOP8HFjFP2zP6NyK/kdSoVHXv/lKydlzZkTJAQYfIOk9n4Q8H+ru7
ptHG44PWkLInaSMxhS70IFrlSPMBcQkEbinzJ/y3FU9mIjkx2huPsSIA1C9GkzqR
TO+ASQ9L+nOMcT7aK77hUOLIQZSO7BoaWKdGW1uR1/h4TOLIc4Kcuvj7MJSgutJQ
g/PB0YqY0xTSXrzDjaMzAcIUqt+GUtb5mpK9kVby9KkqhCan2P0acTu2NbSF+fRt
XZglMoD+o2glpHsLZGQRs1lfPVHcG5tvPIbzTqV4+lyiI8NnqyQvW+ZinjX3rNq/
vrk55E2hBOAs2US2wnhMNqmYpYdFQcNozCmc+Y9hfRRmemCFI65/zXjq58uFDWx2
MHSLoVNhHGtZ+7ogOe77a5Vt4PdvJPQcWzLr346MsCcjd4zT5vW3+H0Fo7Onp9XC
yvjR5b2GkbwZdANK5FLuePXeWI3qLT+vDXKY0s6CtBNS0PNvlvHcDqZabBflfDEG
FC++Bc66TslQ3IqcGkCrX8wtQiHegPriBeWw29RRaRERM3cYZhdtx1q1obH6eRpp
OWbetjkoQ7kZ41u26oQnWdomqdKUpGLDZwp6c9rkR9BBomLqyF9O2L3IvHRU/n0A
fK/MdZbNmMtRhrYU0XOedAtAsdZeTo92kmMSSHOpHsXlbdCgm+xO2lnwUkNujHKT
RUbSl4J/EkO5PVfIN1bpdZewQNx+bpm8PmtHRED3+q7rw8jOR+666YUWM4cG4pSn
m+QhlQoE5vFkEJ5tOUmbgLVTvzPk7xNo8J7rFR7ZfhkiHVEGqiRHchpFDJ6i9ryo
am6dToCjo+wqoeLQJ4Nh8A1Emb5TOu3FRWNYMxZ9f9F6zPnT0Gh+51jDtMBrmEkU
g3SSUILNv7Krbi4Ojy4fjVuO62JtxFmnr7fla7N0DmAyZZeEr04Mf8B5JFRgUGnb
SpJaZ7THDuz2nTWtZkE5dd9xqCbIL7wUbj86aQInDqIRoU+iP+wiTuDwf+CapJlg
vUQhsAczKuAeLI0dXAdsEgtoeFkkplOQKoR8BeAIKEliBTCdr/b2qRGlJ63oiTkq
AspDZH87zrnvuTlIn6URWG2SpunO+PlcTsBYriAqNVue1XGyvwXKDDVZQZvH2dPm
7mGUqB0MgPw/Sxtk01PFG7QRHwuzdJbWubRdQdk+GfwGd1KW6Vh9R6GXfXya/DX+
tTkPwvPKNuIE1hUkUvZiOV7k/DTMsQiV/HlgDeZdHIgWKz8ALqRgCwqS9hnTJ4SN
gCxSiE3/XwjdjgfdNQEepXcbBAx3oLwd4IwxclN/oXJH9Fqv4/JGuinDnaRhEP49
0BSaaDoa92zYf4Wb2PszAiUdKhq5xprE6gFtDAhn7G10Gsd0so/IcI19DeqElZe7
4p9aHojIQdpvrnqYfYb8OXGvsCVLtsaMrPTvSI/EmIwwE8dn1voEMJz9R7idE5QT
sxmKYDpcBfgSuRxyitWG0b/UsIXDq/r/RMjByZT5WtK9FRb1hgIUvqF+WKv4WlCn
anwSkT5AcXlVpDp2gzLP7B/iGyuGQPKzDroxFTbAVJ+rfilHV+XrGcxyygToWWce
m5uGEf5/CQ33sZurmUOCVtZaxJ8IujXf6EIoN+5CAiBqDH5bw6VorxF16FNQbRYL
DfxFbNrcN/mX1Ae/PSCqQqo9O4R5QeVvdHCbF+tb0Hp0b44Qb/vUn7uo9ouHrZLu
xJc9ZjX1DOvhmJ/ZQgwAoJKZsosy/zWsRxp2harY9vjb3daXTNlF2TdKbJ8N9kSA
w9X2DJvdIJC255NUsT2pCdLaSX32ywAy9OE0rfhNcmJv0uL9o+6m2/OwB44rxadu
B0nvBV70th0iLjY9sv3OzCOdyuc9GnfmaXcZMMTPIne7T01TR8zrLwev6+LQjIwc
UIxTkM40YH8sK5NS5jppBWeFWLvQ9FKW3vKJeu8YJtAkAzrfOrLg+DDUStQCjcRR
CiB4Q1QLy6zJTtJDrpwcGFmNl4YZ1h0pnDDGdLzj5TfqLQeXyvDLEeqCg4FCah27
M86ck9RqiBnO0R+mTBIKCtLBnnbU6r7wijKDxmjbfXl2DVInjpgGChu1W4COb9pe
FoFqxAAZ/Np6zKMepiJ3a7t37iM9NTkNSYLWlz0kVNr5X++blFfVkW/t7+6LR77z
+CD6ovotYXxBgBVqfh3DY2Sg+JLgAWryxb9Xi7EgqHrbYx1+xIKJbiqDOqyjSbRd
vEom/RxG8JJtAwsCZlhP+pifaXB6jR9GmDxopOl16N52bbpJnrbK9gSWu4XyLTWB
nyJiBFOnv1XFtU3/iscY98azrGFWorahaU0z2iiMnsC7h7pQoBLZQJsOH+M4BuMH
5L431ZcE48wi/lfJkgQtEp5LFif7H8K+nnmb5sdQUIKK3MwA2GtweOtEex2IO24f
0QFnnAqVk9fqtZGv19o+d6DeJsCDAStzyYVdxveHe8HnGGq5y0O1D6UU+SiRx7wG
eUNSEFxWy1YWn0dJuX6dJF8dr0YIRWDi8szhSygyPqMFUeEXzRHIKQS7yuSJWqCa
HbWqSpJ/Wt2FlNnMChW6UZ7HiacXun4Sa54YSORp/ELxvHRZyn1isikZBvCLdqa/
RGui9z2P3Rhsq7ddxFpT9RVyy1RewZ3ZDOgcrWEFXdPxErX+5yJznLd/YwfIOJQ7
LvihX3swBoppSjA8tHl7zVMnWq6oemxzOVC79nOw9X/eviO/I0SJ5YfnEBAAFPf7
elmUlJ22Xkg2bIbyrPUwnWaGNgvnnkHNE2/329htJk2rvJdi7x8RUhlrnPWl9D7o
tWloURTlUPewS04M76zhFuf1GR4xYSjC/T7+h1KLe9uURluOzQwi8yohH3951jOP
2WzK7rjdYJwAoiRsOayRDXkc/7tcSBhATnGe0P2JFYN182FGAhqtc2iowOmv74vL
g4KBGPFerriioTwySp+7/4VLhR+74Wqbn4Z8Pev11xMYTE7DvoWQ4Ag/1PAuaiEg
8Fdch8ZUeBVQHcz+KLqvBgMDmCq0BbcSVPlrmo+CJvhH+T9sEnt7s5/KPXhdB94d
TWuuESo9s/GbasKzpJKDS1piq8y+9ZSjAkZfeIuRX/P3lFwcMvOwAC9a2zGepP6o
0KLl5o+7Z03ugx8UBFE3LgujT2y0sSaVhOM/wRbCFERkz42mdu8y1eVlmJENpjax
y7uDGnNRRyzMD+LSrsbonvAE82lFG8RJkh2eDJAP0jKx0x7NR6iXKt0tNik2NUBP
eIkiCHQo3eeWYhIDcjiWx8gD+BCYtRAjquTl3S9tews98kQ6E1ZB9XFBAATeeLUW
MlaTZ9U/JbtzLq/CAFGDpTDrN0DChz189tXgUKnwjH7vtcpXkDGrL1plT2Bro82K
VwixzGgN+zE/O/skWzA6LRkcDdWzOhRaVcynIvQl5+rsCOYzFt0orZG21ShXvajh
xIQbQwysVZ3frLfZrY2uxDQ83Eg6SqGT72qry51H+GSq0+LH+Hi9k8ks+DfCBYnW
nDzVeBI+zqowkw32KBd76n9CWZtI1hPP++X9ZIVMgzxUhJB2fIf00Z0fKom0y5sF
b/yWktvSbATG4we2Na2sNR1uKgplTaYWBmnJr5lTFJWbL7lpz/7AnsV4Bid/a/Ei
516r7e1kqoXDlKHYoqQXIpyJ53a5hecVZ9NmYfXW/AGojn74bEorlUxAkJQV/XxH
I7Pj1PnL/sdikIjVCrQXlEcYA6ZCaTxIWaQ8ILI3ieCMlP59Dp7b852NlVNPkLv4
4+Nfkb0d2+gVkW3TlG907nE3GJMfvGoLVyH9x7dmicmLJZCEEALAukLVbkV87rXM
dBx05J5AmVIVRtdU6LgPfXEMmFqSEWo5vHtevuN1IQrAhyu3T8odW5kH77Jwh3HF
0hCaqHvp5epEbAJapwHVPyml8KlrUyUCo+/OTySwdJXgxgMQbrzuhfof59UnzgFh
bwAZal1CmKMFbhBsDsAOPo7y8WcR7BSoE+6fsN8ZFJ6YcgCWGC9ayLZVLRno7lHv
eU/QId9YTHeV3G++7TlQ8xHrT+Pa626gARINRY+3r9TSPK2kRziRvdfwY53SmO3c
rX6KbrtRYH2LFkxkUflYtNmHzEI0YlX6eWdFxDofSIXNv8ZN7QqIJy2U6EsbbdP2
T/ue0l3eZXZKeQyoaKHpXba+OIvPnt8aHqTCpj5uJs9hbWUvkA6IcFY8cju9sIx/
yEdagzXxC3kpf/tUb5Zbf2G92Y2HTc7/nnFWZjDjmoa6JJtdEK/ox9slXV6INbeG
2EP8HjZZo+k0hkexSrGtuhckNW2LVWnBdsFYmaREffM7rbJKjTmjwSIOgODOCrVR
k3kr+WIo1NSAIk1h6eN7baWYT1AO5x2Qk9a048VZ1X8OtHdS9pYQfrkLpEAC2Gku
P1cRLy50An4sJLVOorSPItqkXV6in7BSV30Ihckze8Bwzv//HebLKsoP7Xq2nC6P
SdcnvlID5ADaYtRA/F6uXDL9UjHJYGDhPw+OuxjXH5DY6zbouIC9YT+k0wi7J8Og
5W6yqEQJj4kVVmKOSklHA9GCIN9LYkyvEh7fQRD8cKbuyJLbg4ntOuC14QvtgMVg
KpCOimEW+3zR5njuk6aaLgQtcXg9B9FLYy9mUinuGt27eFXPGkod4qDkTpM9k+tb
FgT2rNuWTA6glSBzPiKxKu99qXnGYfvBuvQG2d6mEs3i17XBHJlc4FxEqXaXenFG
IW6/RaRxs6XVMNoEcoEPnYSNSQ9vQ7SWkkIisTnq4xtv2SNSXraStKrX6mO0wVJH
NBXS97pYBvGhCLh6gaFFqpOGkaIGXFTw0ymusxx66+8gZbc0+GJYG2QgCXentJsR
5Y2bwAkgWsoV7GnzVwQ0ZYZH6MOwBo6knw6oFqjBBcG7xUoRg0ZoY6lnAAXSRm+C
V25RKcEHfj40h0LM2Pl04jmawjPOg7ZZRYDMbg1lkJT3/hySS35Ai7ymQ8zGvQth
M4nNP8BHaVmLw5RjsOQrQ7UV7p+/zI1ie0z2u0Nh6p+aKOnijPGvU+/265gGX66O
Th7Jq8QICXfsPqWGhD7fd+3XCqOFHG97XQNCGPAXoU3RCr/yiGFnkxpvvlYstslG
NV5c4I9Xm4gd3q0j15k2caDU+hH9LbQXkWfX1HjLjekpwjyv9lKPvWwS81ArQz6G
Nr5BtaTkY8WQersFK+AyAPtC9K8S1OsQeawXVeUGj+mdUWxkZdyCNPyTTmcqPpNp
VtW4kF3HQAOMCjp567zdOGXNxDh/Rjfu5bj/0geSgvhB/QFuGX6CHbBxpv0em/vH
0tmSfxObTr/5mKCxzpZXbssP4eUQ65fXS5O1ZsRRDj7dhJH2IaK6PH8+XnV5pkWC
KPPEoTKR1MTvQ/70c+wqwhuf1KjmJYjF03XrqyRXCp2Xo1CRyCbkOXMJr8kiGkCd
/Iro9c8K1D+8ykAMe0sAhvAzht9gPIwYQmbPu3Yys5L4qCho+xq0glQUMqEdUmxp
owWnGoO1dSV96unpHRzqCnaWgluhW1vtUl0WhKbyRGXlgHxiWTGxx0FCxrlvryyA
ytFnMTKnnQNipH+bQleh4lVjW5v1YGUmy9LhdZlR2Zx0Yy2YD72jTp7QJCrqlYG9
IIEfayaZGX0+f62XXR53FUvfhWRBFqiq/wXZRqiDnv7A+8o5Jb1D+5RSpF90bZYW
0J17krbg/9SdgXUStI8fhpfZQCkKmhb6qTOTCUrIYNH+T8ImI72xJ1lJnPO+Z3yn
9IttNY8QJlID1nFesiaWJIIV98G41/8ZLZdRc6MMWMVLhLixaArAHk9/Q19/G5S9
2zzbAfuyP/DZqZ5BZH25XTixscVVQrBPr+FhlG7oEDT8JDu+z1zB1P9f4ZmKcPX0
2f9FsWPeqbckG8EZZ1vb8x7h5Kh8/vSJiKD5F8df/MLCKe3IB4iSpJ7R+Ds3AJ0h
rhwL3x0uGRg1dbV1lXQ5ZgwSnbhswJrE8EHa1Y4FZYHiW78NY6za9IpwhL2iCcWZ
dM+zX7FNb36LsjSTlO65fdIliYO5YUyPKk/HmYuI0rAn5kr4ebaCQ9tnjJ9I170L
uTwUULdLebcqGnOLOizpKs0JhOM9jKufRpeZWEa732v3bheM3kHgu0fPbPMf6OVe
1RfAYUxaonh4xg6HzDrY/6uTr6OTJOxHAcHPIXe+FTzGkF1g7ELCsvmAt51nBk9F
6uoZQcDEKKwqJ5o0KlFGXOO92WejZLvD7M7PNlHa+CyJ5JzaQFXLo+XMLCJeuUaG
0qurIiKFJOCYfKTST2oBU4cyb6IBIMxZkMwcFQ64VOWF/m7TblYyMck6jAC9wl3G
e962m4q5SUI8aN3FGo747iVGmStzEKLjwKSpF5bSPsYhLtWKVxjh7iq6dk0D1duG
CtTHJDQaoMGZ/AeaNYzRKr7w72DYoo795+DPo68anHm4gjAjXVdt+xxyo1t3lM9O
XIFbHLhi/BFo6MKYrBlVbomgUOvullU09F6Po94HEnLhv5cD8DiOxxL29Wo3fVVS
sH6bYrS3xNtORmzP6A6NgBL12tB30deEpjghnM0zYE9NFcUkAO4gu/VVZN9Y0Yd/
KnBTHsGWqgkpifQobTF1Z0CTMkEqv56Ll7n13hSRGSPJt8YlhyM2FlFf7NlPKkWs
jrDnR3b4YuwcLf8q7blBDXL/RXxwFjVdyEf+w/wNugKctUhwQz3D+v5SQlpX2CLl
socTm1lih5t9GhuQEWACUfztLqgHLG2jFX4r6ToNmuZT8uenLWYrXqTVrhHokrUB
DpJZ6Go4nx39mZWvdzvz79h1nRrLSWmd3bdqrtz+ygXZv+ZcZJaFqoAR1iixPoC5
yw7QMcz3gH1rqEZtK7Te3bLblE6h/Z6Zd8xmz+sUo4gS6kehZ3srbkcv6BtrIQRw
X79AviluPc6ct5ER49TngZBlIDiU0VRSnJK5QY5zHJ77LHVFBGPv0ikF0aVJvy1n
OxGWGjbwqVjoMCs8WoJPjVXwywHY+5ND1sYgeXfiojPnOEwzFmnGu0ST9qYBHwq9
RbW0T4S+i/OL8rw5MqfimeDJCcsDE2d4w2+eZXtLMapcDpyLTqapYYOXc9ZevEHZ
P+vqH29WDNTKduxzGPf+Xy8B23QCS4dm4GUzOLp7Z6L+L+Qyb2X4e1DXe1DvOgQk
NqOpG79LP1ujzCrk4JXoccF5xaTm/dCeVnUUAv5zPAXwTAVn82PqFaZhf9pNSXUM
zw0LUlrStyLLdOu/BlX246onVEut9oI12HMAWANgEo/u4pEStBJ6Dvx3aowNSHMO
cIpZ5MIlDvPPIwWdlpaTT4YrORyn5MXpL9wY7M98QaB+T8OfmLXUgGCAOTwLDDnx
6LLx11ZIdCOZlwtugKnDCB+1j/QJQO1w3+hRVcEENoeJR9C+qnxD+KXdughk3J9i
HEe/MN0r8yPRuzBftiu/VosgugJmS0DhrWKOFhFbaIZ8ceb5qMsHLxtcl3Q+Ul47
M45XRmN0wFi8TBpJv05kx97eNS+M+wKSuMyrBID7fNPZy4iCz/CADLlNJXrvGnaN
cQBuQCI9kdnNGdE0rf1+xGB2Vf6kqm0jWTjm2DQx7jXE78T1bZhrOiDGsWYRg7eE
YQeyd/82nFhHkGXOYwpZnXVzNAwf/g2U455jAPYS/2/J8C3Ra3Xl7xICQx+Aql3J
U+d6rLroPtJLy2sKtWixzPRwNsOTn583YfUGm1VdZsMi+etN8qC4fqK+XdvliIgk
bQeow4OkCj+Ey8pR8W41XxqiQAolrcTYGnwtO4z6BjFzODa3hIp1jo5+W6UdkXow
wTDVt3ZZflkfke4Sd/vf/0IoPzya1wjcXSvotxjMQg149ucVZSswNs3aN9XxliIZ
EUPFll+aWGnsQjSYtbVyAJTnAdlSYdSpVykiQ3Vb9sOsFMJpWZxglmkzgDayVX3E
raPU5Nts4zZU3f72HKKrl6+TPvpCYGqF56af108yklqXyVVKSyatVIMTX/iRMF/G
ipPkgpbhjBk5XhRJFXipF2iQAwpx5dm89kxlZZ2E8bNQaMQJcS65J9xWkfZE67T4
W/1VzkyYeDIonZH+QXZJhZ3JoYKyhn3Q+OD5bd0P4g5/6EKin5P7LvVjwo6PkQ8Q
ELmNO+3dHTz22TQR4zuSVXxlxtTHuXetJhB0CiDx9vw7rqPnvWbmCJpYc2xlcmbY
1vxOlxIDcTpvYRb6yQMkpvpD1de3gGoPiA0YK35neMxJyqHXoSGPX+cRQsSUEux8
Y9RFvIailQlkEBYzlcaQkcGAF1DgF2S2ikVGBrql9Z9bce/5tSUbAABr/DcVIgjm
3tOTEHO7O0BLcR1XLiwVQkboMseiwT+UnpxM9U2sE/8GyXFmpHx+RPA2VQmFaGyV
XTkfJX4PXwuwiPtHtmu6JW4Z8uHsUJwYJoTdhJNMiZbRaMc5+1RRVBxG+Fg3N/Qt
Sr/OLoMATBeGz3UNLXu0BvDNOfHTFLGacnAv9CydOjs7WksMqBv2ygGVnUmCy9I7
hOZprF7MeFwzDLi38Ll/M0NDCg13zhgk4ZGG9wWBQpLEW/apk5Z3seR8N+jJHpYg
vEVJo3omQAs2Ox/Dx0I55V0Z0xdiSaLxMJBlAb3DSSA7aYLvV6SXuLmV5XXJLjA4
oFSl8+xpMqcmZc7/Hzqhs1afRXVg86jQitw0Y26ykA8PdHmB6fN+yGUE5WlMEwt7
xyOcvdN52F3SsAqlJtMAiWGwnQZJXLhKsGW4dMslNxrCANmF1OPxDX0No2iZAtfs
+NsN6LJl4iUxd4wIHYQvfRhHAW/dwCa/fQcap0aImZfbx6CmlO+I3ev8QWkxibzS
cGLDBUBQ6pPK7QIIAKjr/4j8uvONttdj0WCCtugClhBNybQ1nMPgllC7s7xCvvtw
xwmHOyXf62TiZxld8HmR0EOYtpSFswSKjPzTw3+tO03H5wtpc9+qXSB1n+2lqRAX
9e26lXWBoPg6PdJ1VXAKMqEw7BtQOgcBMqPN7lkcQzwkwOCHunvB8M9rYFRj9tVw
qeDHTg25Xt4fhuJlNkqmfPpmUxXieeAvw2uH1vTYKboc4lfOZUamfZook8/Ua5S1
TiGMYGifN9dPEArMSEHEzQzOgzOuqWwhioYobQjNpQGYMNTu35j94SXoPKz3KdHF
TqDbFd/ehwaeDexsV9ltZBouCefczeuEi/LCdAGXbfp27f6x3Ml//hXNe7KSBulT
Nj+LBB4uQBBUiDVyOmWoJ3xrmFTAhgI6EYkTCBxHL2nHBaG9oAoQ48I178pebtC5
ewJg/7pPVeiOBUkja2GD26XSUhV0yiqp+dHeJLUI2cdkjmbWekGBMVbd0q4jZu/m
MmaMX+TZkelZRINNW0QAS04+JyAtU5f0z+/SktpoY/qtNMZN2ucv73FTRFjfHLtM
CcsnLzKOKbDcQCTfWz1yaRYAXIheQV7CdLf4mLCeUbOqOJGwrqH1Ap4D6FTgVD/w
bjKIaQV21w/9fJ9Z+pkms3DJ2P5n4dUQd2pABUfJ7ylNPbmJ92ioK1hvU+QjDxDm
M5GEfFNGQ/v4RQqxApj6KExbjmGj6YinXFkJDR4WhoBqpjE8lk1uhpVUH7Pf24c6
3/A8M1s4gnY/e7grPtILn8wzd37o+x7uYpFeCTpYngJDSXum3KA4UzqzGUHD2mHM
zaiSKaxy7HU8l8feCtu7p6iF3nx1BMxiPNVUruYa9yuKsy6bGknZKOCqOaA4twOD
+QNbbi8hnOCT4dyyV97iCaW9Kl6qdZQ+Wf4Gg/IDrisbfi/gCphtInqUkH/SGsP/
IYAc/KWmhlz3etERh65UGJR1P+Ofn9400OwO5kQPO8Ov3bBCbrAVHdlUEF1raCaj
DIqCBwfEQfw6GCmTXQYS4BYn/ZmMZl0GRoM531cftFCdl+UuvM9Ta7PVap9AcdXE
IIoil4rADAFElNL8p8uOkmamISHU13cNPwmQQUk4wYyROHw82bDlf0GXb+aFykXj
Fnlr6XMzLNIxIq6z78nviEW7n2ky+5/pOEjwvmRaiiP6pz0eTXeOu3uWrylQEr3e
DwSVeSo1qMyKFTt4l3iA6IomLB4MTPDWV1An7lds5FH/9zMvcWYez+x5lsD4dFDw
h9Ubh6qunGQNc82qc/hKz+VlZOBl3QbZAYQO6lHcQbiN1UiNC5WyDUd0SlhRZVrO
xlvcZslJbKJ9bYcvz4QH8POohDRxE3RXBYJ6xR4yDHAvVEHxbENtq3MKFyW3apAf
iLOybBX6HkHS9T5XnE9TkkSPhrClrJNTYB+cNlSrVLhu0h4c3ssNR37j5YOzSeji
xT73fFGcD+aWSorRnSxGgKul3GUkYZL3nCnkmsIkURQ7+mVjkhRfErtTbCznCi1n
IHceD63TVuMaay1UTe6qFugIU1NAfFuSnnWsgwMI+wL1F1xn98rMxZ46H76+2WoC
bNYKufVLxpy6vVzPPblfT/xQs6/D8YEG0jyM1kjphqLoKccY0B7HK3K7pwV1wgbG
0KqXkUUR+Mzc+kjJdTDOxuabwXXcAHvAb1tRyJ6nu1XxLqzBwTCB0B8gog8E+bGD
KdaRaGPRsZ+L4CtdXfFEnr3hdxqRIiSt6t5fDiPYiWfpvVf7uKGVc+waUIQM5r+I
aEKOu6TAtA8FsACFIbqccmBi48fPvQg+xg2+2rSNo11VXkQNevKyR0MLT5d6rBIO
uF0Yuh8UZ0rJFUr/UQpTEwW9QofYsocMSR0Kk1ntcOU38fWZSIhYXKBlHGn/IM2E
QU+hh5WXF+tbUz1bMg10XjdHqXbloMVhG2zaJlyCy31q51NAzNqdraKUJqQnVQk0
uUQXLud3P2/fGFaoajL9JdYXXvd0MyFJ+cWjvT4HuK5tdlDitE3O+CRvpLgszURm
tfOgn+PWisqFs7t/z3zM+oZ82izmvZJTzHTOdKZfsc6e+9NIFG2Ce9A9wTfrlnW+
5VxpBa5wQ4GARlwFeNjJa7FRjNtjeWAqwfCUu5sCKOTX4nk6cpqUST5Ofb7wTWEx
RumKH7OwztzSJ2SBWN810/beT0awterG6vryP6eqh5EG1SxgrBNcCUU4+7+95YLz
4rXmCy9nbA2+ZS5neZcPbzJVfeoYQwOu1vCcB/TBI5l3eI9zlkanrdG6ye73WAzp
1yeDLMfYoGgFYWykCL6qckGHVseeE2UpsnkpFn16nNec4TWX444ByN1uilXg3eMt
Cikt+H2PzxWcHOEq3K7ncSIxL7V/nkf9OnaTe1df4jtxNh7zor/uwMe8Alht4WXE
rS+m0q3owfRr194hoxgKicCnKmikxXmeBDSvNsxpIrNo6tB3pq7q6QJHI7b1t9gl
1fzg+RDA+kdX15aO6NdIf39Zexg+rsg5ttdFtwPPdAXZ+MtMRqX+Zs9Vd0Z0EpQt
EMH+CMA4nQmxS8fbWOg9pmIzun37NTrkfcZxyt8/UWFUFeiSb0Qvn6AgKbmmehdn
rbQR1SsQL1/jAJZd8qBNfKvOg5QFxGx8yWO/n1bja0F8jQw2sZNqdJ8UAxcWdPGw
mfDtwkupL18Oa3tvdKq+wUPLZrwK7cF4IvSFIav/ZG+sQbVSEqD+EN/krnTyZTWB
inN56+F/BrF449UsXwCN9BnLyUCkfBT1L7FUKd+0e0jay3H+k0C0wa/IVtrGecxI
NQfX0y345JmZV5Z+pyUL5A+zcVigCFibQIUEfIP9ZvQ/H0AgrBkoGoj2h3VGaJGW
pyd+m/3V/GBJnJl2Qve0AdGgnUgnlmJEnBUEmY+0wL089CsOoyRsquxHaqzxZygu
mr0tdCxguGRWlpiZS/ERFzMn0otGvQLcBmL6OWNPyADZ34p6HWPqJXVZE14ue1Mw
z2Qf/6cQ6he4QXWpFV7ieZhzw5+hi7FgDD8DpzBX/Y5qMxWoVBS1OKmlu6s2Q+Dk
wBVhx5jTkFRI3g6J6h6JpkJiDzl0XFGb82yBgPJ5HKOwegQdbFfakPcqs5leETgc
KU4xSgJIjzglOKa6cRKKhZI2GiJTrpfQKkDBNNqBVWr3BQ0Ve9IaRmEp2lYxWXMq
0u3m0S3CqV8/Qx4BO6pEhsy4n0XsuNpXs+QYMfg0IDDOqO7tYoaIHdDp6Ofpytz6
wtiKaccXJ8rTWt2Z+WcOtv90nHqOoZGXLJQDytMaSoM1aA+T+kU2j/kf/UaQvH6t
JljRmwLjFXFcbDopGZzR04u6cTtCTJi+jTO8HQiHA1d98XIFVhIKIqB/v3Z/YbtY
D59xBlFLokpeVlr27nBQM5IW16lthKDjbAz0zO6HereAyHRltnqTNNOYwUigEc3Z
P8YU+VjOvORDTUtBywgWOYKKc3//Fvc9sq55uheai8BTZG0+6cfcY2EnlztYcWmW
w9/D7CTS25x+bfUwgXrbUbEBs/gjreNn5s/mS7zSAqNemwDfFnOQuaMP/dBOBn3B
sSswSO5M2tLJC/zbClP0mTpXaElXs03SNHyoJbV+uUOr5YPIhhDu4Uev6+ZFPcSI
XU+ZRiL22CLvIj9omFrnatvly3I5AhY2+AfwqBilW7RJNsufBmqeYTABkoZUPh+v
swkQz7t+0G3hYYs7QLiVY+e51ky7lxZktEMgFi4MRtxU2eygHUcjjjqspgbjGOO/
Ozxq66cuUozkkqRWmEQcj7V9TuSSt4fH1QifJ4YrE8lRg6k29Lc+w21ACbMPkqou
mwb/HwTE8t1UANu2dMNUTFbKgz7QFGb2X+LWNMih3oo3DDt1bFdnzT3TogwGCGme
SRLS1Y8NoVQ6/sThN3x/X02/vnjd8xSUJe0OOZGpLrHOXn3W+ozAijYkjqTXAz/q
D1cSkPf1laYPGX65gA8m+h+HKMk00AWYxIJfBUC4NqrGZVrr/IgzERfxoWl6GOEC
llz++M10nn+tJAmFm4eEY7yqvGpQH4PM6lpbEtpBjpuVuQp/zGNeYasKl+mOm6XK
42ypPNyNdiPVDUklIEfVmn2Lf/sX11lbMuC5ztZngGabIAVKGqCyS3jE82/ZXk8v
tHTVeRn/01YH15eUSi3puyDE7ksSLW48vm5XXqM+6DZ5JY8uj2Z0gPC8T82uHUGq
KJTp0oL6Rb2wubHVW2q6xmnDRJuOhYHFSUxEhQ6g+J9tN1uc0sovqaTQk5oZBZao
LrYDDDOwAgJlFMZGGFFcq6Lf+6BxU+l+2dAVBTKxmOqzHdj+Ht8jTRq0L1cMutmb
2PSsloA+4Op5vuez4D1KZeCDAXIj/Ean0gQ6havYDz3Z/GG7GQI7Yn8sh5CE2Rc/
kK0Rwlqr8SRSggh6XBqSP6TvRNEHn5AH1pfoiXkAhHL2fZfMs2D8X3vSjD3KW4kW
zk8M0AnW20FKFsxtpz4vNfv0RMOFSETkORzMcQpPFzMobB+22ya9ju7O+RUejVyp
lKIaFuA+c0JbtwU8LPKhxFlARbEWN488OxBXGWObybWtPP9iCm92JDd2IhlBK+GR
ie9NhMdDkvX/38OymJwF7hIwItylPSMPWtZjRBHjTpx3+2eCHo/1DEPCRgMdKqGc
dQcOg5a5o9kFEYzVYZMI5SpCCs+ycs0ZlobJlN3vGRRWRyDP+CThZrBeg6VwebtE
TIaGWaMjlXciup/K+oy//pOeBShotpZf5YcWO7zJggztn6TNEw+ITyQpqQLUA0tZ
+NW0dBaeyDIkrOzuZzWcUlYowioiI8kRWhyKjo+8SsGnXMmBTU7WJPGwddzjmFbI
xRKssQKOSQtpWQXVZhwI0WD3amFu6W2VTAOXo209TnLq/wsn4/0MoK6ArZzIlEfn
RmvKszTTh0/csYZh3ViSDCWhGn1qkaVDOTQ8/0oM9vy75yrIAI4uBBEmupRGEpu+
UkH3l6rRZF9GOJv7MaMCm0RHL0dwKMxUOYgoe4ZLhgy/R5l/eVABU2DpM6S5EEdG
BX2Id7d4I0jaCJMsXR842gqi4Gz3NhV45z88BKv6219vZRTNUq5jpX1PMtTb+beZ
NSgDsZIVzxvwXmeoRs1hd+6KBDXWnosP6YHX28GjM0OLLTO5jcGSliY/5H/QX1eN
MyElSYj6xRJHbi8EELaFQFzwRNMciDE4Yy7LXLHkXslepqGHKBG/6dO8U0kSPmuO
NFyB/j6gB33QJNrnAy6TZXFadC3Lx7gV3qospt9xhuM7NK+WKNQyaY3zDYA/BInk
+znGP3/r5yqUnAP2HNugHSSsw/oJbN2ouHKuDrLGFJ2A0WETKGWqwWP8qzH8PFkj
L6qh2piyj2cl/kk+smpij3FpWDVMy3nQ8g3JQ68tAlGkHHGnerowv60zjxi+TX3y
euVKrjZU0Dxx10GUptsDYFMovZJ0qgHfdmRHeNxi3z9zkZB1ZM4InliHXNmPWB33
DA8BfhU2OLXxVX3p1IakEJc27IyncUYau1t13VPg2oYA0WHF+cD++uvWjqgCohWl
ooCVKKNYf4fWYypocBKvUHG8OSsMuTzgj1m07RSj48P9GoCw2FzkVDc5LGMw2A8I
wzO76eG60w4pu8rmMFzdRiI8FR0qMbgRiK0Em6wUS/ox4W2RXyQET4G9mC1lJt1i
Lr07esnqdu4VzsUD25JMcp9CQByPYa0gznAEKIyXRtc1l1avS9updf/d8opK5Ubl
FDRBUpQSpTUS7w95/hTkES1O0F3V+6QllGF5ErXHBu198nBcv3qpTrQDl0lcIaSZ
au6a8cu8NHq1o6FStF7YRpaobQSF+ik0eaZt6pIC8QcAykz12epyhoVJGAXVdEoN
gMLcVsC+iahlrrdMfdCJh+5f/ZLrjiUWxVWYQrg9S6A2VZfyyyI/tYJ04YkV7Ltt
GwgPfKR7Eu7hydx5d60f4ce2T1bLFEm7Ro7BAX6cMlO+6LfKpwgEBbBPQ2+vaFES
O6yvPjlrqLnPXtbfIpCn4l7/cEwsnvAPEwvHqV9MQZibgcpD1+7rxU3wQAJw0DHg
kUzGIc2a8APNClxfDLUd1vgrZ7Lt67X4bxIdAhpfAmQGG52gV+BjCDh7/gP6aIlE
CQE6BwXxGzglWA+V/C+nJnhR6kYiaHgIX3dN1DvCl1vRAXg1o4Dqpy/etgfQZY5e
+Ce8gu2RFZqsaxLx2aG59/SVWfm25TznMSuDMxfGCyVjvD75BgvxAAdYeT68TtC7
fJS1WlBSr/X6G7pBq9tBBunuTOI+eRSWxMoYJ1xs2VnSKeaL4uWQ5dohoIr4RrVH
SZlF+eachCg2+RbLBKzCTo/6gWi92x4D/Gkj8JecECJfNOksTtzXf51khlAafQIM
q1sKpPdfWHEpJ16U7eoZYUlml9rturVoWeQ82mqfignk3ZSaLxCEPw3EyjK9FnYT
hbmgogtQU8hpO1zGc/vDq/vHEi2Pctnw/tDUEUy70UG8BYL4rNAuSZWeWvuP0Hp1
NG19P/R4bVmFa1z1245Nlw0t61yeW0uiWUEIBfYj4Q+auXqgNql9I9kSyHKc5TTS
QPGotZ+GfL5HMvUpy8ynFiiH607rgKyMFmxWmBLN9DroUUIZiAwLjZzKD9V0uPv9
Vi5XK+U28Ff+EpiVTUBjKficmplaQayKArc+WJNNjBT3bEO6XauDETPtsbCIQlEw
vRXOv1p78pOUis6HTtD69LihxIvnKW3oRh2NRpHqPFdGiREWoUU5mRmuXTQga+fp
Ze0opbzDHb5+rRZqJsDVWJR2KiwWPxswES7A4+xDlyjz2XyhdqDFNycxyGmTYhns
bhCHX5S2NBsTVy3mSmtwTj3cWb/xX9h0RHvSZ8dpVhWwyy+rygUJEWnBkVNKkMA9
plvdWkxNWx0ORP2ZoAk/vfX5uFwHBuURcZy5qOVOkLzWiS9Um5NMNBMFWL+oGn/0
PQ3ASKqKYSVjolKydcmoJ5M9SbMK4bJRWlRRhZiy33LLQ5mdK2VPCYMdqYw7h0bO
Z4dEPSi4mK2NmQ/Qf9XjEInxgeUvXfY35EhbdrypI1U4LpLuA42i6oQa7li3ixaE
7bOI9Jy05bs9/dzKcYJHTUZaMRye6UMbdmCdOyzAkuPDgvoXEdd5RPGYSJnM0TnZ
yAk7G7s+GGP+xBqJzIwLRVnrwBM60QAXqnjJRDFWaV9bCuuXLLUumqMY6yBlsMrQ
ZYVyqp2wcNz+r7zbn+sUzP+w/u+eBT+VDGkj+f1rlTtWwHh+tJy/UshlE2PrNr05
F94teeXFt3ePcAkq8YjUpm3IstS3LCbukjFNUT+Rm2xVk/X3MCngt8MtQVbEllgM
H24z3se/y3cDXAQgHLsVy9JRHzBOfLC/NCgzOXTGGLHEa3/+Ikmv1j9w7FvBm6DX
jySEdgA9aCpDjBqKK1Xxv2lD+GjniGHsvFJRymSN1QQNVkuyPHYW9uPkmkOuJQ8i
p3MkBxb9J8+ZYk0E4AcdGioDixAhVEExesTPa4ijn8q/7Cisd6jmmnedz7A5BG/V
9u1lGLbq4KJ6egLJKmbgDsSbMmzsnTGBAaJUwYqE1/EttZuEGcb6ov0s2+87lDIL
bUy+Q/ZQZatHqr6bs1IF7di3TZsdgftGoEJRl/Dq/JaKWWIn7nMuEFu5KHBopMrM
zgiaWPNXSgjssIRFR/yIsiEoLlQSXwE2WYb6Z8fynPYAOoOVlnxn6LnvlxcDGdJ5
bEuYIXxGjvpxvRx9b3ZiJARGRjuebw76txpm40/myex5AfDoeklyRvInS4WwuJn4
tyDHnNNRzO92rlEdNXdgx6FtIvmmq0BuHLweyf0ApnApSJdGAUuELlbScPCrfqVE
RLTBrrwQlPXUQ2Sp7Q/wwwY0b3JxJw41avYzoF+C1vtz9QHolOYLk7Yvxf46kaG3
SRDM9unPiM1GScyf/psLXi0NohJ75btf1i8KYaXy6F0JLMrBuXNcGyMarJEtSs1l
B5U/LVdoyjAlwXAAY6zbsaTNWBUOhzE2h79fqkAaHBWQDLrPONTUeCgAkHKaFemE
gI6e9pgadwfV91ulZ6eo1j7t76gX2lzSIGzoOtuF5TkVWiEpxlmFWlk4lf0heNiu
emA5Tk92liEzjKvNHekqO4V2zV8YWNvTP1h3fKw/M31IzprCluPtCo7tCX2xNovx
n5MbKlRW+Nw+xJAVGuzm2S90koyALgaW95kkRBtqOTKua34l7HBJ61fKMp++hE1q
YuizyKCy4sTCcZE9wVbFCwVw3gx7vRf2+Bi3fJ7XqaoOWu2Gm5/gYOq/7aTTbrc4
1ub50FyrZEy6Ht4TMEjIWDCCHmw/3dWlzejQBex6FsTG9snEb0U+rXU1FHCMFtop
DVkADasXWg4Y5BOQd7jH7KXrQJo/dYbuY1wRDKl8co4HdIMESBpFKqLRjHNZhffI
xnur7JWH9ddX5+9fQjGwugXXB6AqogWPUHQq/Vi09RyBLShEMc6SCs7u/Sh35njn
UjjdhYTY70p5tYbu6TNPLNB7Adw/XycBnGzJn8QjvFy45w8YhOoOUJrNzCLB+Cil
RpTIVssw4WP35kPf8BAFFwe1Ms62uSnZnKMAOPyboUrsjM0QsgsKkgXi9J/OQpJV
7KAAJdyXHM7SmQnKCK6uyS2AV07Mayzd3lEqDK0WRcSh2bJR0B1xPqeV1BpPLBjm
qaaOOsM2Nf0N5YIeuh98SiAbJBvMkoycE6Q536an+X/c9QSn2RyE5xk2vcO9/gqn
5EHnWpodHBrqq5xO7r7jwjczDGi5Sns6C3E3zbhcIaA06h+VWegxVPIV5SK191Xl
I3vhWeUvwBZzAZVsCT2GmIgR93aTuYVWo/jrwh9J0ahL7KtqXSljnJxRqogieqYx
Ty5O2cGqnAFBGB4/kzpRABeVCIuEkzIyh0m+U+6i8VcEYCwNIqLBgtwpJRH+2kks
eWB/MEglqX18Xsx/WdYzcXLF3j90ejejfkAbzsud/NSxaV+Kw5rG2cVE65r78p4b
laddpiS5BNynf4YcM1mzgDo6zNh88TqKo6mSfsdrlNg6o9i347LkvpQjAZutwsXS
Q6dCoES3Z7pTnpjzKPRs3z87kjwyWYrrFEi869noIQ3c8SjEIOi6CggrLc+oCpw/
M1t+NeloyDcZK0b52B9A/LUWmVsN3Tu5QqHLQnV4o9ntZZMO4QDHFlXf/DcWqR16
T6Jl/ugopUC+VgubliGPExQTe2jDnuR53HuvZejkhSztZgPFVI66fnY6oQFAE9/O
h0UlCUIdb6PCNKKKQVVfANNfR+t18jFVYoQxi6hV84BohFMmYLrTmu6v/DSLwpBt
buKdwmR2xKYpbA7fKK5d6rPNERwPHfFDvLrWw5q6NU0U1ysLcYJDlQ7pd1LpfTe7
HmO328rosBwJmYTuzZnm49giPzrx/+bqh9wHqSa7r+VFweOlPPi6kMwCnNumfHX2
7lwREUbt1TtXZ8ha7eJmQ2yzbdCeBhgfPp8L0roTSchliYRvaaV3mephr3QL3jLw
hXulmNhxwa3pZIleAcnlPdQGuwIm45il+3Am3AxdP2zsZ3TPVU2U9t5pQeL7voge
s71Bta8U+9rSltZl457oO28BEpKMnU3yNYDOxEqXNfBaaFePmuQkV/Gxl1VQkfMU
tSuSgzsqyD/Gwjl5K/oHQeiYoQUmFG6oId6ByTCuWeMRGTZiKtpdVl5oywd1DMn9
syDYM4agH8G0PE/f8OYi4gFYhxiTJ5ENsuM2mVu6TUVaiuZat4Rw5EkvUAZKGK+E
52YTxBqIC/U2RgEju8Qg6zKcePTRr0a7XmS4SN81wxisxn/zGTBBj6AON5yTIEba
8RQW6EKlLievTJpMMyfJFGHMuRMMvrEkHPemKfTCR94xYm87gkJLjQv6nvyM45CH
BIdYy8PtzafhqS0Wi7I9kVmJVMXY2kZlk6/S8Ap4yeONgmdcsMgnCogkEHDnyYv6
FLi2SyUFXpc7De5T1bND+A0xiWmOOcl/Y0vuFrgplJ8aAkv7eAbQz/xUxb+5ZKjP
2ERqLEBSJjCK6pUwS4/kBd/e9wIPlUSb0o+xBD4fllYQVvSU9rM9nbf8VJ2JdSJo
LhM4OujaJk3LNVE3lyFGFt83RMP+c8HRokVsmX+9G84tv9urF1XBnPVPrCx9Ff8+
EQq3bCSzrbfHVmNcrdF9s+EhyIdBK9oWD28QlEslMIZal7SzNQ/mejWdf1JKtcUS
QR/u57j7qPnLj+B9TYEjn5Mwx/h5mqbsP1XTXeAOe+QLTFSjEmaYnAkzE7rrZ4uw
ZS8ceDJzgGtIXI3ZBwdB/ZcSb/hs3cjpVdKgjoycCGYCRjlqhvGmQ+XDmN/nRqT7
EGbNPlF03oBQSxBAoM2HOQIHAnDIWTzoMu1TFInwfVx/chQ+7MGi0pnqpciMx75k
E6Tj8FkGj1G/cu4y2Jles6Pk9SawSn8H9NVVwi7URb5S7FvMuD/PbVKSdikonzpf
ujGgeOeECRO+USpBdrNMonR1D7vWxoGqBxKSRKVRxEWXuoIEOANBUaDEsLodzpLf
PxQmnaGtp5Ssm5NZcZ9uAqsGvv7HAtLUqHKDkBfuoLU5u1oKv3N0iB3qrAsYki/8
pVdHNGIo0bySLooj9hNpXHS9119Y/5mm3VtyqX4D3FpCWm2LPYYIIOnnR5pxRvuL
mAUYnq9faFMmibjz+VCJfuvT1gY1RGrqv2wprhV+ST80hNZpTVuaoQ6ckb9tpj37
YVQ2Q5JMLyV5Ve30Py4+nuXUS/DLqxU50ySx+035cp35oozbqZDinYEwlApZZGn3
VjRcQhXAqifeRRhwUIAGBfZmT/qM2qlXE8Jnk+G20S5CgxI81XzW/c547puNekfW
JWOcDeyNbP9s/m+3SzxfwVRaeb8h1mlhQ27Gg/OfqIpo7HDKUb21hLUeD5WCmhqr
vnnkN763rVkPsLahuNS1tsctWSbbovMLLZstK9sDyuxFZgXzknStV1QRvKM3d6YO
JkZdpFXzEPrCWu9YHcfm0RLMFCBgktysrXJ/Bunp/OnIK9jgp39p9EcfxPR6JUwK
oNA6yX6FztZfWFONyaXkbLvz9rXCZ1ERdky2Uf6gRZI1EZu5bEAXa5UuH3MynRCO
OW7+FO7dPjsA/dWMex1M5TfBrazfJlCOoHrpTgW/oK6APQGM140k6KB32h5mz5g5
baFMIg9D/9ViLwuf/7+O5RU4r31xHQlO/6TKqkSjEDHROebuEfZCFGRMCi4iF2/6
k5Zr4kEc9tUGlghW8U8YQeG5fyhkjk6L37IsXfo8X2P+pfHAExQvo9wGvk7/SQ+s
iAbUdK8EZ2obUmBRpUFPELooTptCWkhbkF0L41vVnYY03PmJ34Od1hczyrGtqm4v
VO8eI5F/dYb3CWw6jkBCkk1loJHL/tjrqWR+V1nvQum0vJsBae36iaHHc5H3Jzam
Xtg5eNBhZzHYbZbhfLdIuFpnnEL5M3iMVbGNyVInom+bIRyr7qDOTq0OOg/1Jky+
eMlsIxAmmBFZT1J8h0CoLM6JG1EyvO1kcuyJqk+Uc9VWtGETwEMSge1tuH/gff+y
/LaD05Z/Lij5phRc5KJBfNR7+paQ3q4vW2+2FiG+kOboKG6hM3kag6lwEfC7Rk2N
s/3r4jZO9fimg2DMmzc5ydxMJcJB0HX+b0PqIXGYyDsCo0M8eqcjer+28TcF4efM
junbRs+xOHBmlzHS6ADyEhRan2j7uSgD2lWbw10+YiBWTApE3pA4I0KFpLOntbkH
yPrPnxnBiTY02ivbPhdveR51UNm7TfD5+6xDqgpkuy6FNg86AeufJJGF/CMJyuyk
6rkBBJG686TY1GQFV+ubx/9hx9eIWWXlyc5OagWykwixwOLQy1CNRlvEkcQsIoW9
Dw/iK1UuOa/d7v3uPchkcEOymtyhMuMkB2VW/kTI4kTclEdOpbJmD244vZcDcGyh
4ThjYC+zIoyDEcY32XR7RbdCPWkMwnedxmFPSK8loKoQaodOn10IuWxkkZeYfdD/
7wBksZlTFKpI/Zy3goSyKWlXk8Tin5UsiKjdW9U8igSf5p9UXhcrUuyBqg1E7P2H
ruJAokm0XNSE4Nuorkj9hUjfBcVuYTsBY+3eyqKUWuYTgn7qSumuF7kpBpYreMjC
Z6GTKkGuu09aDyjrBEay/5AsIFBokfLy6EhzW46GY6GrDQP0HR+V1e4eo6LQaPgh
qbeiR2jezT0Ex2U2nzz/80FqGBrRBQKEinhVR6apOcEk7A8glFaIVZ9xc5Pwu9fo
66Duyi6zPwewf/ulUSmfDnOUibFLk3wrIxiuKyZxl3L32u0p4G9RRKM7xgMJS/pq
+xEE8uAt9cIjtfeysOLqna8aGdOnEFqxz7yB5tlEoa3NIi8PjUr6Mj/cfX/WzI/l
IL7pkKJ7K2koTbi209eVeZn1aY2ufuIM89Mrfe4werX9M9xuQI1OaGme8ZhxpwCY
oGG0qmYxMdMaF29+JwWJ0kbwnO6qIR7jLLywlsZYymGt/OJDnH78hytdUixfRNDe
hS0A4bmdlJPSF5sdUkL/ioqzc6Gjn9c0IQXQQHYo51hjTOinkk/lhOhVd+3lFmYe
gEKAHaPgDcfnsv/1R1MSPdcVR7KEs+/Twn76o6Mz57pdyFZyF2SIPfcCtGnAKROD
Tl7ZsiO0qS1ujc8nnzhQ9+VIY8+38bEFVeM0k/hYlHIdV3cVbywYan+MdSPDFbKI
z8fDqAQ8rW/5mF8KtyjDTnvO1Ky8nOxRioZnjGGflJjW6NbnOTBRI/fgv9dLntJV
ZClbu0F/aP11labcjaPMVE9tASzJHs2YES8LQZlXkQ8pP3kR96UZsFdLt/Ry8apk
+lk1ty8TvmXhrY+rq30EVH1juDq2L/E3oEDLtmUMijha6KKVwkXFfkaJnHWKQBMM
qPo+Dl1slE4jbOdhZPBjYxRwtCbOM+Utn5a0vHPJi1uWOttVWTqEiTo6kcUN2KR0
BBZw5IpjCEiSaUuXDMym+T82YmMzLmEq2KsFlVTGSLODmJlwnRTqjHFKvflKpdp8
bqQ5jrLwE+aERgSmjBluqrZxx+o4QXYM3ywmAtwYJugz1kmpdLwBItqELxsq3q1a
MvxW4dF0MSGshbw1T7tgnL0stTIFigAa1tpLPghF+fikCw9EJhGYEy6XkuBvEY5q
kq6UZHQRsqrF6k/WKgxQIMzIiW9GL2o6Qd9YszCikzRqXHcVuxxUgzKnxJtqYAMd
boc1uslLRSNmxDZgjtV31CThX6MHDBRrFiVrPrIb7N02XIjSWASAWXTB5tyTkhIG
9MVKhtbJudOMjHJ4JzAhUWUgN+ARvxFCJmxJW2IveTgjysO7X0+HE9w5+UtiRrCT
STbzKBxfcnISqcwtLJgP9sXYzvy6ql9bUM6jGmRGrqLmsppKQ0Pt0UsHNNzuFXq0
R8wIMmPQIsmRaphSXn6ro0As0/VrNCoBPOS/tUf4qUsiA0muDijuePM+8/Q121Uc
lUfjDgDTDprKSzHbvfR2+q8Dpkip5H0dBUeaZLF1+DADUvdEz6UCcuHLa620PTnQ
8+n9/qbQ2Z/qHwoLDgHBoFFKD2fnzY5oHilzhJt+ZtGzJDozsPwSSqwHqO0efkb8
6Z3mCaPrSz/vYPzsx88o++YAnckVrz0V9oUQN+HfmBCT0r6ccBImS2ReiDFntBtt
EfyNpnGNywPFDipE5gmoPnItvjUG1rBNC6GwXXLW7rXFfaE+tMso2dZZ8BNS6nk8
0HhwiGMu/NcPa4Ek80Cq8/gO/6ifxpMNd41572vCtK1Q2lwHSrcibWWarf9pxyXk
OeOTCy6VtLNqO0ZP8zTV4UzYI4YoICXDssoHnIqiahtwk76CCn61RBKl/daoGfr8
/LlOQKyQvh62qvjPqLeDgQX5R5mbyYLyj0Dxo5PgJKXH8i9W+uNTPCo9++C9O+9g
a5IgMRlkosBqI+wisck7Xa4qTFCTqa28LIqar1RCgpH6uX6Ipg0+z30z/FPPMKmi
e09UWePV1+Dpo9sMQ4Mfl1m2dzunjIlM+ncfHAGsGVb76Tlidf9RGRKEYBg6P4Cs
W0ItCnb9ErTE8IRXVIFnXxvahfHW2YWA+drBT/KQYeyEgY4TxWi3d3w2ESrMSli8
g/TnKycycyoRlylG5lHBbQPY/Mntp1hVpzs+Z3glPMvOtZers9u2O+m+0naSgbm/
qLKjQBe+352F3nUA95YondkNGdLIHxuUDEuNkoL7ROQgdlj1epQSz6YJacNAYmLa
pr4s+7nVui/yLruoclUBMtmdBeCh2kYYexy8xh6+JStDS8hNmrTSwtiq17Za57Iz
+u6ARiP9OrYoUMEikdVN1RW7Po3mY7fPNyv4kT3+aFw6vzxeNu8/Pkiy8Z6Vyco6
fFxqKzEq5qBEVSG84cvsEQy4GNhGlJGwDbUBBl16b0Hwqk5rQLeOen29wD50Cy+O
0D446TfRkNBPkkDY0cOnzmn+C//mpaNB/UUagxG1evlaTu/pybvInxulAcmS8UoV
0VbTCO0E1t2Rzhi4KAZnur9uzUC77ZIoAiUbeg9xiXK4SEC/ev4sOtaLVeUJVPrm
OXl2x5wS1aoiHMGbVd2ynaQr1sGdw1aqupyibAP/u6WsKXhL6ZMxEuCwnPZ397wb
uH0dAuuje5RXaS6LikDUU8hlX2WkKUr8KGE0KnEWuZOPSKI2QoMs99m4ep79xwTH
XOrhCN8Sj1Q5v1eApMmdY+I1DAyT34F3eq8xDLaJr2XTRiN6bBoCIaLvyq62P38z
hZJBSq7TagVpVCh7GL5Z7OEwJ0GOJOOqoiZ78ODjFLb3P3aJO8RYR7cjAks72TAM
Xew9ur0Ku1FB95p6VpTvmb405hMtN6tpbACsW9Q1zNeuZ/ixn3emg62PGgEnhMpS
zVly+mb+hYkjVhrwuBN86gE1+9Z12Gi+fIJy9A64U2nbAcJ62AHXLYW51zj1ClVV
teF7eWSocPr4nHeE9ZouEzkMVbbgFW8GII10eMjYqes8ONsu1+U8TKKUaD4PcTel
ZubYEslkLbl2h8Zvt3tUabucwA1J1wBowtT/XZ/RFA9mZqy7b2M1hpwUDCzTw2yW
SRqE6sB5O/EYuTd+Ghvu/9GhfwKDAml4Lo5sTybCkcK/jEYnYTe4BkpC5W1+cvci
cQiK4R/3yH7hdIbPJqZhZosEAzX5a+xGTNFQFhZewJzKQYvFSLHeMrUhESfEJlwN
cHru6M6vXXbEoivEu3jLmFRoEybrJBwcKswUG5IP7Pz9Mc4snXhYbQdg4HwgTCZk
yCbn+16IoZcqzxYxSHuCtT/Lq1mEwZ6TFqgstBN/61lDD1TvumlU5LivX+Qjox8R
0joYJydo39Z60osKH8otH/6gdNTnHX6CoYHo87nm4Jl3bTfJEUzp40rAKyRnv3tc
PErDtqJxAn23pvX1H6JAVB6sqLvjBrhtQxmjE8w1/iuBWZU9srT3/AYeUlbbtbyw
QOBHVOfytU0Q7bSKRCJvS7zs7iltLkRc/lI5L0m2mm5gsqjGF4Tyy8SvWnhVhRz+
XEkYFjzD+qwwn/Cuk3YRRTJ87d+LGOBoLliFrYJlT0hKJ8z3J/f/37TXrAGdSCg9
ls3647k9YbvvHsv9NrIZpM3p8G0HB24PFOWDirbRcVhxMVf5RTTM74eWio4NNJDD
ZoQyVwaUT805PTn3Dqc8SpD0Ezntvs9hfgxj6UYMODJ7agQpcq3AUFTWGzfjD//r
CNSlCBClDb6SNj8tc6kDBWiFGWXeQH/0GWkGpMZswUdCLbrqAPkAR015bGu+QOBZ
xnhdGUVkjS4W+tZ7ZQrBriTVwtdip+bmeT9aL0+DEL9A3HwN4cBCEN1YeURwoBU3
8MUzhgHK1Hq9JLAggKR6G879KHodA8SUPfuQwx6hOH2958yS5TsUvNUDlKPUF4CS
E285Ndoo49rR0TrTCHZjKhBa9MAzoPitaV+mNo6pH7OElu5DC9jWGH2b60UkZMyv
GGei10HI1PvsuU9nc/6BkXWBXmo9GAnRSP5ITfS9YcJLF1ue6Q8WMxKxZGcwWPBF
w0I0cIjPDnB1LfwP++9V3l9EYQKTzjeIFVxUrOt8Y+SnDRnJ1wQ1pG+7bNQ/IG4u
0Cw0hqcxcuvVt+7Ij3NBqE4l6Fcsh13Z3R2dI3l97LxfLdUWBAbF62JMnlr65uo2
mpB+wAwevsF3cetcfxVIOmSpUQR1xxTHDxtdp7hEMb3BbJ4GZEkeGWYm3AR3tpIc
raGzzEgZ5p10tEH6NJcV/n0MNfiNF/N3lk6QnV10zHk9+Ojzpc+/p3VPt/jgY47c
fdxo2STxCD9u/NHhD2eRX0H7RE4zbsw/Leo5P8Mo24/09tAumTGnU2XufDs8g6SK
DHuFEGyFiEJC9A4D4vwO/NIdTAcB73lcCxrtpHz1pCrgelOgNO5zzYdb4pYoukrC
E8PADqc7WT2Zkl2WB58WhafIyoTEkhU9y2Z3eHw2lScPWoiyyOSWPkW5qhkXLYo9
6h6sBaNV17EHk9V+md3eQhIusLccFXblv5nlkz3lv0SCYkV+TBl5ULms3W8wxyFO
M89/JfcRz0Ox7Ey8SoKub/uldpqySdt2JDUp+ycBnOlKu0nRdvXHEipw6bDaJ5ck
mDUQQct2nqiD85D8F4gt1W+Ffsx552KjUQlcg3dTTpjRRuRVUueB8180DS0nI2Pr
fo9BaeBRHdhF6IN28j2Q8fwHBGYBKLjiaf6yHayGu++WQYNxi9qAyXEbtVqNVkVs
IjkIVQs07psU4jIXjVttQWUbFGxI5beVxqkLxdYNsAU489FC/T/BR6+1v80SYw+a
ymEz2WUI0B9hC23NPdwwSRWCm+/agBbdTUd2IUqKhY/lYPyswqUTStBzLdZtfwAb
awHE+UcTiR/pYIgwmEGMpt9xhg5ZDIWC+xdJfQnDcX2AW7aiXw5iU78TiBvqq1Lx
b67owBBdAlEyqtX3mzVaPSauWvRtpaQR8LQilanSBDGWF9PGLl0v6gGygt4bs0Lf
w/cDWn9/LozmflvINlmdNXfUNF+zv4MRQU0wiUZyvdqe3jYt2Faard0tbeV+VxK0
PI9ENpHiPUlY0aJwjf5b37mZ+BsL6KU2emWgUH9nryODnryuv/sAzNOVouqNQfi6
StDT6o62gHgJO/fJv4tiSGiIL1yMJD0T80a/23tRHzIIOBkOS8fo0RDhcSZlKLzF
fNMlZtHuzhzzR/SGohO8OqUsO1vbi5lGsylkABRrTS85hmb3xZ7SomSA2EK5WuHF
kUxcyBWfVD+87DfnALtZJLIIL8lhx1vXzZ1BLc22XaSZSZQJXzn9Grh/Bi8HUy3N
yn5cfxWsTiFmnItB3BuUaEpkRKKfX60j3vNprHK7d2vI7UKalTOi+6/OAycL4SPx
vVwf0+tdezWiSq53LN3/C0t3inQWS36keFS2e0b9FjfTZYfEj9h1I2xQktzIaZ/i
JHbWnm/JX9o0kHcWBNKxdUBL/wpFi8fTD5oxaLXzb8ECOk5nlJ6O3Iyn1Npbmwhw
JmUV27/3SphfJwHfUPRSAbwnshWy3tCuN0GOeED/5HRUofO3OKqTzs+XRCFoxiwP
i5Lgj4D9FDMQiCvpEIgVXEj4mJbP13kh1W12xv0wlnAQnrpl3lhZgu5gFfsYgsir
O/g+QNl6NgXcMVoVfPlqjfP9XeIrADl1oKv3VDLRHp4xjkaXrBLDelEv0nqv6Xwp
Q9i5UHdzF1BpMdirBSJOACHOJYHgsq6xvKYKFKPz/YGtHGpYW4KbsSb4PXSjm5+3
N1T/o7KLggJ5fVzWs0wj1FLgF/Rlky4S2mak4wU0OY0St1wyKMJWqlsFzFSeS0Kr
UaTKQOni8lNwmbYTEzOXETTY31RUbMfCBMYOyfjywKgnDONgegv1N3ZQm1JPY3P9
TGWa3Afzc2EKQzD1+qBe1uHjB1B/U5JZhRUaf6cpuv5+bybQOoK/8IuvWgwdgfhb
SATR+4du5HibhuMQmcnxblTj6AVSFxYg0qeFDD5/lolg/QJavK8jmfkLkRZmUbnZ
XEQ0hbXKeZBUrcOtJ3zr3VO/93YIYg6Lh9k4PDPjUm9SZnK9WjoP6jkkeYZVHk5z
2ssTmoHGwtg6Y8qKrOI/0I623d62aG/6R1j7peJ72+zXeOfpZeCsFpdEHBNQywyP
xznguRGYSnBZhrQdUxzPXapDsmgWaXf5NlBl5pjIXSUR9LIzl9bUYJ+L5WhIbJq9
Ox/0Fdkqs4NFs74BVanCGLjmrnsYbqbNfDBr0T8sy4Jc/OvMaaYQlorkm0yz+Ya0
6E8PhWCgDnZVWYIxRVYnl7/5+An4GXlBCZdaWEmv/DrEYZuN9RP+0XBjUZfG58Rk
7K8sgBvc6j1lkpsw3anVY9G6/TCuA4KDGm5O5LqxvR8WMlbkV9YThL62QwhCnEOg
TER0qNQ7Z7nzsyBGLKKe3QSWXrvTRmo7MRQV3ruQph/iTWMTyjUy5ypZgBwL2Yji
kXyjDVnSDH6FzY5Jmi59XGo15vPWmdHNp2WMMHekGjg7CuSCaFFIUjmBCDDhdb7B
flBmYrJaXM9c878tImov9InqSSvRRqIgvRLQt6qWujznmuyStofZqSAhja8eIL/r
a3io5MA81tpCW0jIyv4ehJ8zW13BAHpk3qUzPQMFPwKRBHJFa1VKW1Myw3PELhwy
pjrGWTc0NqTjV3anWbhlyb0RLzQco0fnZnnTx3xtpvGnWk8+UEH14Uq0mEgUFyGq
FvgrunChSaIRC/KgFVdzNlDzcfOo1dZIxBrcJnonSeYIkIP63W8GjV4Ti+I3e4gN
mC/mPgG21wd6+tGDVBhh1kMjmbYqYGFpTX2/MLp6wzc/wM8MQFUuA8ia0pMPcbQa
w5g5G4VpIUtqYT2JV2guMppcE/8sJWi3PQR8m0JDqrer6Vc51Djn8phURyAUoGKu
MhmaJ69xIzmP+CslAHDlqMJ80OVKX3uVh1rXe4ChxZ8KlkILKSiYdSs0PG6OgXCQ
0oCGPD3CdLxBTpuzrAurCueh76LfGApJ1+MqsAAOllWsNS5zGgc9z7AXEtSh+kyi
xKyBh0BjzAmba15NUGvcIIlTMbgoir6dMWp7U4agibPW7G0hxgIJ2+SjVYS+SrBF
UeaM1BNxOU+WHDb3rtMJh3kn9+6VQHv5yFwJBuxOt1Ifpg4/mvT7dLP8wirdp5/x
Ffl6FyyoFcUi7cSVf/PEq3SGdHSbE+e7SGgaujiQCUsGvru5po/3ebU5tSuylDZz
1aW3ZVplSeV013vqDaPvUK8mmyhVBkY34Fup0m6koVWqePaf7sqUTNhc82+NLEQ+
RL2X4mrAP46CPoKk1wFfZSx+jWguKDVUjigXvmF9XbePnGNUOqTgwjL6Ml2nxeqQ
MpBpyCJrO24mDFxPV8k71nRbzafEatj6sU/V+noOG9irahjhEzbH2fsGBm3Bz2Ti
UAGYLVf4SLItnX45QVAvhu0vGQx3472Li77q2Ih3BkAYVV+zyvJLeeSSS2j7BRCY
2KYKdKbjBXIAzh02QwrhoZCzwAsdg1Gn1KhSvrjKyZVfMpWtP1C7bOEHYwyEzFwJ
HelJ5RBvTsIIpx7EV6LbERu9tf4DcU10Bgg+hetvQzeCqd3+sWSGm1CO2ifccs6K
O4swZCdAvWVuo6AwabieiuMSgS+mgs0Q4wLJdnJgLAnJxT58mj+c8oCl74TTiZKw
n8+HuDnEB2/37LIPZMqoqJts86cEfPsOOCdK8lgy9oo6PLLNIZgDetPjGBG3gbSB
mWdsUoDZjo1A2PFkxfAxi8Qb/JgFLsm2FTA69pGAttfq6+1Tg3MA2vl+f2OzbZ6V
q8OnmnGpG/paJDobVM9wYfCxLkSTume995mV+6vCXGyNbDLBo/5SNjXT073TNZ1t
nI53DW+UhzTjGc0Ks94JJD0KOX14tMXxdBEaU0dh+RXhw3jufFFUnlAEXefEW5cY
1PVS4DmByI9H3QZ3ZNTDKKLLiCZANVivn3z7vffmNcDxcsvak0cYlPx+SMl++JlO
nVKS0BE0xetGm24oIrthmBSfjZl5DDDmuumLoQDlHz+jp97RTD0bXF9qObxlKddr
Gas20yGB1GfPk5jwJVLIagFoNvLgUbM1DavjzkpF9nJgnNW4bvGQ9FGFfGXvcgqv
nBhOym4dy0ngJ1Os9uux17fwjX2YiY9RVks4P4ZtYnc1hG0xRFI4Zy/2lqiuAG33
lotowcV/D2W/gQ6ItH/wz9Fc40rmBmEL4KV87VarM8O6bQNbEW6at5pbMBUI+v+C
dbVOxOqTMQ3ylGk2jfu9FsPi/7GnfQckY6WeVW7lqFqdvew7N1Y+WkPElw0nay/+
VyYP7NNVqa4bioKBmvGLzPmJP9U5TjIhWI+ApIDtMWf+eLUQUkhAD+Ki6fIO7FiS
PnruxYv8X8BXWuHn0Whmz+rx3psVjhwzD1i3yxDFBhD7ahpS1nC4MkhajXAezDah
sUJRg64wA0Q26vMczUc5/OPKOx3CSQmEorPuL3JC069cArFsouOG4L1AgCAZxh60
N6qSVyTdoNLENnafv07VnC9M6YUCJ7jxnf4p1gMoO1LRQSR709fGp28sqrwSkycr
NCnEjmHEpW7S23NoEZh2Xg6WGBCmTRlVcpPj6YpFL99qIVQ395OAVeQkYZEpjWAp
6fEybN2vLYHXvLS/5WdihvKI+EBfd17m0WJFREKMtSiCYxl6yaoOGzB1KVvSl98s
2gwGV/3kZc7NjAn+YNezHlTyl6MX904k2MGWghIYnElyPDTLD74SX+ieyKWoS0lt
J1zDgysWKP6NJSnIMuA3b9u8I2gdpyfezJ7cr3Cj92tTlFhXb1g+NhFmgbJoIrBD
/no9YEIyhJWqftvvKetN/kbSHlO8s5fLQOaRCwNrODIk87FWXaAEZL+3J6+3/s2U
KkiaGptvaAQz95T0FacTKG0q4DCNKeHCRWUlvH/dZd5LzWo12AXunXqJMaWiWCXd
e3iLLSR90Qbo57dvYkeWRo012sxjnFlHkLrwwsvXctAMKG85Yy3ABSeSmt1uPQlM
yfLWfE7rVjwxGI6wdVPYSEJhJh9mG+iX5XzmAPqpSAGOZv6MOxAhoWg6/mytOkq7
7Ck/O9zcMbpQBW7dzd+QrO4MTdDPHopuQWuFyqZ7Udww1g6VlVal5fR4viN8sAzt
ePjdL/DWWUGxidZQzXAp3zksyXc8h+7L5YlGrldK+qPDLOGVSgnUeg4DPx44uw0q
EdMKJueMnl6opVfw1AoHGFd0fGKJrlrbuzBhQ8AB5LixR6hYAq2x0LOddjCkI2oo
olUwHXqJkhrP1dW3SB05LMuUZ/kAxZcHDPa0rji0n8mkZI3BOvvYMlifJLXDDqgU
fnAm07XFHtRCxh+wH5UexF216W+ea/NuSYHIwjZhrdxiSqpFIuz3UPoPqgyU0MCt
4Afa3Z+WLUrCxBk5zSWXSIMS4ZsaFlGH6JkOls5pKsrWuVQY84a8QbTQYBxIveP8
Z0g9K7nAtlgIwpt3Y6O7hOBNFjvPCcmSfGRaGh1C2bW6Qr5sErFpNWM3qQu7bseZ
/dpPTi9rQpLaPHD1FHLDrJbZ+ustU/jW7s36fybEPFNEc2a6HjH93BYckNBgKPJ/
MQXODYw+WwY3TfnReII24hy5XaKW89P5xqOsuaalsOfgZ0LOxjQdY/RCzTjt1Z5W
qvAKuKHwyr+iC47dQeZcmj5slmhiNCpScoyoFDa/d3UUE0+TcfypPSH0wrR8Ws8+
cVTsLd3RzcInUmok+nS16eIjNLvXdvzy+i1cidshrvO1CDYnNK8kmXkfWJ3wfAUi
rqF2D73DyO36yk88xbppeZr2T7w5D0hjBwhG4IkSorHSY2HLZ/3sz5iC/p0dgb2H
3Zy8u6NME2NzJacEo5YYne66bBQyb+OQR/Hmp4jRENw9XBHFQWQIP64zT9+29+9a
n1pIa+Plworn1qYwxbVqDlICRJ+0k8s0fGw+a3HBv3FWL6zs68bwJB78p6ZccH3J
/SzBwYXHvx7F1NewkWm5JGuA81GdRjhvsQpZAyqtEp+8HcsMOmDYdwuV0dpET3mq
ZFKFn7R1hwSj/DQRH3Cm3mNQDF1lx5jJuIR5I+zwPh0CwJoDcd80rEjgT8E7rs7J
nKBB5V2RjWsoOCKMXlWmibhTTyhaPO4UxoGiawopYFo7TyWody7/YBcERuYcwVmg
IVB+edr5D4KSezqfSwl8wNo6exCj4h3L4EtDlsRHPG6piod4j8eX2LxMpkGcksLp
0HE2ZeY1l36ihF/Iv1cPEm+8Kr2YHMJCmuIuy3kZfzILhviMtMljjsJtO0QLzZxr
DBtol3VT0geTn+iOnifRnFnlltrK9s7lXD3kNAopk6kXQcCecNV651s0GpKuR3xO
bn1+QeY972QfzpKNv9Bi8FmVfBRCRsBt07VSdEJoC2ZePWExMwCN3tmwnagpyhEP
mHaHVTifng+qf1I0+BFc7GQxp22DmUBfjSTZZCkooIOncrFb1vVYPSK1CyS3dZRw
gtIYugcUWRDeKdD2KAsdqQw5hcEzbu26mg+gJ4mbUHXHzU3aE9hryyqGpBqsH3y6
TGyQr2a+5GgTkdSkxIw3HOlRtJeUqdimqOtGybZDcoK33ARfVQ3kALl/Hbe/3KLn
m8ox2jMCwi6ekX1TDpCLBco8ORAY0OZHK47s/onSeKd9ZvrmNAzWomlrnqEb0Ndc
nwkpdOQuARoK5YhLmb3BRlj5kxLReEFP5ADGKj90ZX2AdhYWpmwNYw35FV2iy4GY
NHZ+X4YWqWMM/ZYL6//8eqnJxHJdckx4kLKxTeFTY3TxBhPEKyJwMPsiplnF3T+y
uZa0ragWCZkoRzUd5JNKZx4O3Wu/S8I0b/343zfrGad8HFcIk2U9xenGdYvM+Sv4
iMTbJMCfClDjcJ7Mg+EJNqwkLtpA0KlVihzSXywk8ESM9hM7C1VMNGlYe7SLV/sw
76ntwrsoxNzGlL2ygQtDwHEFUAWvNNlSv3oFf1QOuPeonZRCgsuvLDaCUGS4wdg3
alAOXiZHCWTkPnQ4f5pQVgbbqecQn/sKhPLNFWQwH79Y0axdDhUv7Dkkto4UCI7e
lrAv+9wvnzBh1beGU5VeA+ClLIqH0yEeFLdkYDsB3/mvA1DDbGQHb5tjtF5pjj2X
7JbNBWhssipO7mEO4MJpJt+zmx4npMDD+PEPtM1h3V7kTgGgIJw4lgwe4D2hKwUs
vbqri1I1jLc63VL1dSR2E5jTRv3AHebKTZkcPdA5JejF5Feh/wWRKiuzpkLDOUEM
xXHmpseIS9iPK1J9Or+0unIViJdjOM65QQsruA9xT7PtXnmKkYmwMywrxSRwZ8eS
741/rudyIeRKY3eTyOyArcJC8EkDg2TeiaWPC7Ve9n0H+pBEWcqXcGhZ2/w0mSYu
MUn/unCnF97iM4oXnak0riypBdZL9wphHzz2yO6ZznSPaftNKOCghPKZVjzOCVFv
4cMNNB6Zg63kypQX5KyJl7/i2PioYHyCF8ezj7vGaztD63PbC+oKaK2hgyTdE40r
JKeZb+3F9+zpU5eecunx+LhofWcLonR7MP2Bdo9OCcjICeSC0ef/ELtdCqtDEheP
HmxokQMaw96QoEOqln91TW9M3f6sl4C18+uudjk7+gNs6C0ZmAG3GWGhaueG5Lzg
Gq7l+AUcK//DCqDmoupk4BfECyW86rm7I7I+TyupaWVv894o9uw2FEc97enGeWjF
llgTt64bwtlYvhMGC4qcuZOb9aASgF23RoOcsuP0UugRPceUOvAQUu2F5gi0Bj+Y
uwSUam+btzcRT0hmVDD6aD9xQqdUzrWUpUexufkFLoDlW4hCFcVB8pdAYwj9ZfUI
J7yvREJpg0SAb0noS8as8MrlNY4bMaVBPeiOP0kgcRHyewr0fS/aX+8dxt/5OZDx
jUe3aAOIJWR1RwKunSEfjrE4JUiqaJRGhR1wCJz/9Si3NqGRlaEplxsQShRs/Vgn
MJtGyJDmTdJ0dVpA4NbOeDtV9PTwrw0+3bHbi+rIYVH04sOsJtVOqyWY+gl/V02p
bG9iepfqkGfRONafW0IEqUwLAJEnKzcSAFQ0jlmxzJQeEpJZMxF8xCuLeqhbkalj
KCHUoVUiWu6308/USd2qagfr1mPngG9ungFOEh8Mg6aeZRkZBfPNHGg+kTCKHcgT
4mnGnkxB316NwC0zqSwL4jgDVwBwjumUyOV4SiNatEOAGQluiTQcR94GXupSINZw
PGLrh7k6EtDGtQnIwYbOAzRo3prou18eeinLdRqtNoJhN1PRaUZnHZu4H5Ke786s
3VljpiHPNhyRkZhB1NDs9ugEFj7JHxFgy0CKyW5mjxHE5yg9usjgk1eeFmtNbcH9
CDA0NeqpAb4UePuMVzvx12xxCVOFVPzL/YOsUQNiYLP8SS/yRwpm9wSXbVn3GuG8
RZJUnLsHD+s4PpWCM2kNiuW+uYu3vc8nybdPd0EpH/JFUEJhLo0l78QOwb5hYcr2
EwxP/cZLGsDC/uBqRceXzJHgKDsQs3p+Vo/ln88PWtUyRMq3+ve6zc6vikCFLuXP
Zo4xQ9xZei8JfpQhYHkYdH9wuR3spwcqHtHLoRmYkytpHfqI9YLJD2AR9VEM9tQj
Tnrvx+jV1idiMwWTkb2d1qzv4lihDEhueD9uQJk3OgCJkNhUlE61GoI54/70xNwK
z2n43V/5NNDGReORsmn/9Qs3ba3TSpN3yA+XDJjjzjzucV4kUwHR8y/m3m66nvaZ
RPj/Ykd+CKRv1koxjHIS7i76FKSfibi13rEgFnUrQqyRMmgl6TyMcCFSfbX3dpIw
FMJDdal9MFbeDzj1aV/RI4a6sRf8PY/ZcX6c0fkUQnK8Oh3NZi0TyGNdYejd1eBO
W+MdRidq3IuQsXofKsseDD1q6P47ASRxiQbrW4zwRPDXFEBITw4vBKeXXL9InNSF
8GOALH6CBmfrzDDVwvmVvhN5xogtJutZvqALVvwxSPdFnURKDekdixRpIgM1dsdq
q/v3uneVPlffhwlGFW7RUbtcSjsG3DQnGgGnQSyXxBIM/uKJzwp7c9cXNRwJv96W
HR5b3w1b2umdA+cyyG6TYC7zilyP2In2gkC6YCOiH8VtBiu8Jzjb/12cLUqRWewP
osblLU6t0LxZuqBGcyj+tMKiJZXCfrGgo6hIFqdNeiwwbwAf72cS2yW6fJHVK7dQ
4l9OnlefrU2tJ0r9iOjK0DM9tPyxHWOeac7L4/0JyV8xu18+Fi+wD+xjiw5tUd8W
qcNthps3lxmedF1ox4lTY/E0p20z+CSdT5JBG6/CEtE0sB1hlMD1GBjbGzHTFxZz
mTYpP56iq7Q6VAe3FI9fHgYYndp0aDWEJ1ayRSWCPfYR85nYBFytWhgofYfzHECj
1EhRcNjLUe+slE8Na8yaCoQFmiLNxXqQ9zB/lhifEWognCeRsX7vOLs2q1VdhP6W
sSxkf90VSxHs/OyAUhssjAAUNLX3zdDzf/w+uj4G0FsfqwtNWxJnyw+9szwHOofQ
Z7bV2WGB3jHbpPknAilLJcxvc3wvfrF+rb78m9L+6asDItQlrwjzrToaMUc3+2cv
wbbC4VRz7WCtlh5JRnkmsuuDjS43EvTZkjXKmNifn4Z5GEqd0N800KXNazGRYjYq
TZo76k2BZWromlrCJIes8G25JLdl/F+z4YueqAxvckNamn4/Ijs2O7G2L4dW9Kg3
lJ2BlZzIdc7QKhwzo90ZT+xbf0wzT4VisLc9DNt2cTME8iHOnO8e9BRD5wpXJGAt
CmjFm9o8m1486JA99ledQDMq/8Ub1AJztOG2B7HkGsJpWu0Qeb6FnqYJU4yUNxl/
D+GFIsnLwofxdrJXXUq26VPCc0jUJgifFJTxzHITeDYrI2b3+rG1ie0o9rsFHj+7
t1RwO0Exn7pgYgaKGiQdkmnz7Z6H8H5pyypY5OdBnLvv3foZVsL3k0frMyZv0eDk
5o1CfJufY4YsuB8sWm8nO92C8kYNGcHBPmLjGprzHvA+iP8O3jBpx2/84qJX4p7n
Qg1i6vYUnwFECtnjRkDwVKpnDq4gYW7P6V4U+cHV41VamswfPCTVI4YIlNajniA2
6ptL9xCEdNT2dq6xFO/GvKnOmu9hrpGc+HfXJcHvO8EKqv+ShwRi4mZEEiI7Z6xL
pqxBE27m2jqSmgpaya1YuZuzA4Qf/08Y1SJKQ1SLY82xenEjPXJCKqd93+hqZWGn
v1iXCqyg0FVztmWfeLeu3/lxpd3psAiMwYkbqbzVqfCIWJNpuXG7/3SnKy/ay0EM
HRKD8R7Y+8Sm7TAQP1iIryncBEurfgfSrVGghyYxQZZS4Y/7d+JccY59uIrs2kGZ
1cXSgHsP7ysUL49g3DLzYpeDG1TFrkJgOPPsPYp/mqESLwyrwjxcLDpLVF7uYnkL
tPredN85jSKdrIjqrID/tlkqYS7EVZbAS3IYu6WZFQBnCG47WrrMJndfSwO/ZvhY
svKhQiEtLhq+Hzi3htA84KHY4BjUHhsNBR5LKGgkE2YqVgCeOZeYT6dVb0Re1+gk
s1budhvscv+1jb9hXi99cx874qq08g6DafnBW+Ez4CVmSZQ/IftwgsXtDDfYf6w0
zd+UNbpuu+ARyjeNRRZtlLoCs2NSW0Mi6Vp3+4/yVZEA8o+F4dKYQ2r0RrIk+1/d
v2TwalelT6xYr0nQn1A2k44QHCUyYLNHEPkHi9Dcz1mV21gV/Dzl2Me94HTujH09
e7pp2FAFH1hv5JNR7TRguj5bWGWx5FBBFN8XkHTNvHHsoyy8VltaekzMYZz4AGa5
Wmdiq5biP6cLPazkrbG9YbYVJJpFwdQFCSfIwoxLeOoixCMl5SpV7OIDrWYK/fR4
1JrRfkYD+mcj4Uwd3htVl4Zv1zNql4jF4OvjJumoZizF0g4F/rR4hruhgALm0hIW
ahHTTFMqbWAlFU9941xjHxYdWKtXXofnqX1ltmpn67xMHJI5/mLbOYK0Mxn+O5lK
DKG4WqgmfGQDnF0bg2/AFid4Qg2Xl9BpZ3z2Rr5I67UhPMDlZrqKGKkcRnk/7zNf
piExuG5SW7CpF8lkyholBBuFrQXS7Z4ueI8B7hOLJmSbjq2Fu+y+0R1UF7FhHa1x
fmwT3z0Srqv4FVavGXv4jFNRCrsjAUL6SOHg3EOZ8jRL94mwm06i4WDKAoeXVGxN
wo2rMQuBwDKE2ZxgO094XAilWccE2r2O8NdVKJzumJxND98JsorKe04NqrNSdOLI
093T3EePAS942YSxuagagW9EKjcQu+31KyxLZg9WrVlSDNu2RywH0eu9/murhb7D
fBZTBG5ALWFmovDfSemYmK9CAEpoKoLcJLvsCAN7d7WYJx4YSOZpKhXHSP6jNTop
1CQjY9h2RDxF0wl/zzOapwy4HCDuANlAQtaBma5jB+320Bo77PM7+l1KCnQ5mPpW
ZeuCU/GHsF1XFX8lggMvEBZPikKfBlqDX0Cua9Vx4jfm7wNfE/PIYUWxBZRfJ8ba
4u8Y0yeKva7u5cSj4rYHZgWTdCfHPf5dDHJPcD768/UAFG1uFibmWf9gkN1WAyVv
muu6SOSmn4KTITcitrni+dozkobzXK0RaDdYezv8fXVIAjcBIUXW/wKZQ61YV480
fG+bAGTY2qd76mih5IaS8l1jwyEbriDXytKYlJM03mf9woXHe4mIVj5hlTflae88
joQVDyqTvv12d5nG4XZVFqOkEybctMNb3DA06sah5TuVo8FBoBEGGxhYOuZBfx0B
SKeVWTzRiXVcD22+KRxgUgoyKfI3FwlBe3069pBvvXVf93v9i5RC4c640ZfceViE
T2a657PxtAyr3uxgpQzBTMmhB1gKjcCMgTS1zFd3P6DNS4da2mPz1rZlwvefbvQX
Kkd3NCzhk47fG6+NX80ebL5/fS3TzzQtLSo0Zx5yMw2yczZHKgzR7zaRkdKKhUGo
FDB1sUpXaGVBJq70T3iuTqjEd4gbRYapdGyCv6WLWgH4KMjoO1tR7lr2LFyJvK6Z
WDZsSRq5UjXt9krdyPbCoWaqKPsDUanzlSSR2wwXg7stv5M+m1Lxt9+2vah1ZAkg
GzVL+tu69YcwCTBf5zjDVXBZk/AzzONtJqNRQoNn8eEyEEvOLbUbZO/k8fM8Hm2N
0adONJMZM83Sh+wV70e6w3F8ZCf8g2v7Y0mXomWMNWrtYbrtStmmzuNKhwXEDC6r
0lk4z+naB6QLZkWdpxy24Scy0/7hOV0G6I2wbz8+MVgqg5bLx9NhsyEMPbpGb0+m
wPQhCBtUbjvHuxwutr+b6mA79WX4ZRvCyYyAw71P2sWWgV1zhdQC3lwX6caXsBgH
c+rNxvzPdYPt0OPemUqc0g2lRaeladg8NOJtmc5pvUJuMJi5mkbcPGZY9udxcpK+
QtMGCIFiLh8t2myhkc1z47llKttDD+YR/zXqSc+QM2dDwqH1s0MnbM+CNBosiRrA
kb67ZmkEpuwe9niII1VYzY0oWh90/OHghfDb0bDr6bgd1RE+jAX8kZJzPL27XWRL
ScnU6Pe2G/11EkN84s6UORS1pq25QRSrHHfCT1jT5CCjWibvNRtqPqL0tyrzH4JW
BTi/mvizObdqUYJfeQflySz5RwJuDifCMbhuQ2xtqnRABKUHt/Ctrie/wfXWBZut
DVZ1N02kKb4yQU0tACjK7+v/3/xnl2HLe0aT5JjZ+erO7Y6Ch15+8OfE1tKOf0gY
tlbcap0D1hXuh4hJmjOghFSja1H40+/kZNgnS2qoFHRgVW0BhaAI+Y0NQBOKesMD
IWc4W4uRTi5632ncvz3oaIzeBtC/73SZpV1VOmbMuEprHGBvtZZHtYnpYo9AWsLn
KZe3v0HsX6chGavbwYnD46Ij8qTg7Je7Abc0Ru5dOa5ogabyT5sealAfFcKBYa6j
xtrolPxCzIUPgCglcE43FFxtkBPkr2d6+Tom/L7wFO8T3jKd5LIi3EtvEZCWhj0i
nAf5e1saPYjXKxGrRuxFw3bGTyNjATlSglxk0UkLSpncRpPpf6ilx5IZkNbFfeJa
ukF3rr7pYdBsH6wt7aTQ+RpnLKdAVA5DYvFnf6SIMuVoJgZVGg4a8iSl6r6uE2LU
2uh1wxjGqGH2wbf512vna4BoCkz9mH+50TTGo6grV/H0FJOqxsQseULyoYx7uq8L
4O936242W7hRmVJVptqCBTGWl8H8RAhMvGzyOI8l8Obd9sl2kcRTK3n0xNn1IrkD
YTYVtoLzQ2PNGzZYY8X5oa3qQJPQTZ1VxsEuUz62jjSzyja+xID03HRnS3q6d1W7
l0Eh9/WO4QBXL+GaBqLe8pUFrRuyplIO/qnhKVtS/5DJNE/Prz4tKph/1mt8RqDL
AOjPyC13sO9qYgLjrnTLKifbL7xlyo2wEl+Z3q8SIwKRbJRBFv/j3c5csV63YE4W
KuYOCredPEi6Ri+MF4AR2m+4UA9qlrS1Mu1m4XCdhxilpxY5ySM8rZtkkYcNBVhJ
RFufDk8E0DY6ZQ4yaBW3pGElbtlcPQ/hrtN+ggqdhLb7uhhRXkKfrOLKW86wyGIn
eUyaNKCzG8tXrZQe5OirJXbvaY8S8ExfjV7V2eNdgk6rLAiwNMzIOcPgfkePJKnx
KNtLkeVxHv02oTT3e6moMOpYyY4KmAoFxrckxJFprqvyS5K4HEVfOX5NDJQsF7Qg
pCbczejP48XtHSWf2XAz6XFrTk7wNR1osXEEMiOEicK5F9+Tm5rN7gYnbn8HAePJ
w1rcR2X35z7fpQjCS2GxEHsad/ji9nfT91IeHKmRBZnz46sLlcNOov4GOA9/qxkf
K2gweBm/B6KnZptuEFdJbEp1TbgY1Pp2hBfA4nQVz1t3pdK+4uu1jjgtkvObmH0J
tMDDw8DGoLkMIjhX6MK/xcY5TxG/lW2B5g5XKgVlmeqW+9HD4fIXnV+wtLn2fsb3
YWj9TvBuM01j08KvMLrha127lNVKkaBL66fL+NKpa7qORC/uWA7pGYjpoK4/sbXP
LLQnKq5rG7cLWw8ohvwZ5KKMs7djtFn1GjqJRLeUNjNVhM0zo5QxFHNZ4VZV3xap
ZquYZdjxNpqI4P0yqBVT4EoOMoveTi8/wECRemU90JVJ4NIIoNawKFxhv5mV70cB
2Z/h29lWvo0clQwpxUZDfRS6LMU3XKc1NlQV9VBHSXz/g1p2G8RXC3uyRvrAHgtc
bsUFD98gm7H3ck1nGVM0WWI5beq6y5JMjhQFq/9J7XykgyZQDsxcSSZP81Hz6Sqp
JCOb3eS5oxfeqR1RHf06FEn2fToFRyLarqTk0UEgQRq3bJzdCe7T/p7k79g9LGE2
sNqq/8jioJiSldwNeXzHk8MAOINWZbCnBAzusr6Se+pdLDLzT5d3z7xBWj5y2X0h
ZGiHgfhtrU4xuxFPvPhVN5xkJbtP1xAE/qb3QtbJgDKelX/tQI0se+snpF5gZyXP
Hp5Iuy4vC5PQqJcDXPM7ejsTmdXQ34izBOXY5XIyChM946tXe0JFDB63yiacmAni
N3R5uA+U1kvO+vPe9uwLzRZ+sFBOUMYTaGj432BTT1y134zT+PJ+NbcQuayk+Eza
UNk0za9KV5D9Zgv66nUhqMOM614C2hApH4irDF/QnUPzik7AeV0FTVhyeFZRcFc0
jXlsj0C93yFXyk36CSK8FWUF9RtEJNhmdpeoeQq/NVHFrlPfVCHyVBjH36E2VXzX
YA6WVQOb/3J7QmNgeyViRoHjhBsw1OHlVWKXxA3Lkgk5sOkHXDgHMrZwhS/j90Nm
lv7+9MXv6DeUnDqVs57/NAI0kSAGwf7V+LYUzX6+VNbGA5qjNchTl1jLYFpNH75c
bHvAmdzvykQDUu6vlsE0Umjgk9SEJgK0L1YEEGPPsksSG2/TLPLvhvgRguquNx1Z
7QEKCQeh1uO/xQ7qfuogPseJa7fVDGpg0EV4MSKnvGGyeob+EsEXJTEPe0MXbxNM
RtBehkdcwg2MejjUfJCibS9D9bnAAbmChwGZvecwvMj2mEMAmVRicXZHz9XCUY2Y
rqiyDWOtDpIDH7xswPhJY1tCf9aAwT8z6p3JmSNu/pkIxBxy6FhCNvZpVVkLuI7A
j8kTPdgu962M9GpUjwbPCpeUONsvjpB22rLuSx/m5d1i67P4yP6+CeTpbHP1IUcp
Scd+RbYW24AayNe3th1M8geWr6jn7Y3uENV7OfbUSyxGSkPvM3auKNCgahPpi+h2
E//vvx4W7DZqQQ9OU8aYIZSetJFe/cYtzTTOHVOAXZYlDNwVqV0Vi21fRtIDNZdG
JEdzcEzcNUodBwmpfHKac1vYfJGKUmfcetcI8VE+g9xIBcQlc3stFo9kj5ixWDbh
iCydCwWb6W6jzhQkF5DeD35F3QQKAG2MilMf3dDr1Qb0IS8cpnTuzQ+TVQ1n4tLP
bgQdR6iIMS1UK4Mt+OtC+tlV/7mUctvAk1PPV6pVxtLBVGeVWs34a/8No+ibc+aU
eCjPxAlXYK2UpCW8dH9kR+BeZ90vd0deQNyLlEScc8UPyjJ3JZjBpEWm6slO9yRs
F6t0Bs8avCDAlsvqKzC/O1HfZ3UIxfdCgQ4Xwa583H/zd4k3aWGIT6aCEXi8pkCQ
7vsWSFsWXq8sFA0BLS06YaOVigZAbhYemtGBXUPiJGvGxJAaxhuSjaBO2KaFoopL
J1kkXLbFZaOXXd2H1sQyBFQBk4HilMRA80kEwn1aeXRz22is9bpY8lQK18sdJubM
nlBplk4x4PH3HY/b4MBsZHg9tMEFIl/WI19bYJFCxp9lYjfA4UCcMeLMwLyCeAnF
yWJkEhQPqdqkKcdgFFhUwJspJUVLoaXQ68rsvEVKuQfdatEs5y+z7HuQktdsxK3P
JerZ2qmFU4mWk/H5hJxvL5Z/6WpdBt8ELEWXNjfQg/FFegkQEAlaOjjJIA3bzFVw
UhtmRBLqM1smrlYqlkHW3uuIYNvBhadqQ0SmGnHDQkV8BUNWm9SrBKgl8yp0gh9m
Sv+e7ClExdDkZk0gPBAawHirNjtNB83BQCa+3Kg2mXnDuimFnm3mxfO28H/BonLl
JoG/H32fuRLBX+DhWhOTuE4TTIM/Aqw++5dsbSfrfpGgSJ1kGSx9wVHD/4N1SZXk
Du3cFhx+HpLA4Rsgj0n6z/AixOxiuMVgYZ8qKmdzx9vuh/CvgHa09gWmpAVqAD2U
oLmjtUzbAADADGCU7dqL2UuHjYYbHmYWDSivH+r78bekAU0Bu1d4HOJKQ+VKlB2i
zHh7MMoTCcpUhY6m4VJfCo4G8vAbwvplvvh09+IBAWtLKWI2+5taCGrIfRYjO3SS
bewJxEUt8BII0Zs0twySYledLD1tjRI+GHOljrxp2s99kMzybcrcMovXd4CQD+di
a037cvZnM2IHEPZZ9/xXcXibXJ4tqY3q33NKVhYxdN7bLRUiqu7GY14gVXymNZbX
oG8XerYd0ddnmY9CAlUWQE80hjkrOhoiskVf5CxpIjkSbApZ74yWf+UcxCKRLOR3
JXsBYXLDX3vIziZo5nRjBQSVxQcxFYpKWuJGTRxeR4CVsE1CkNngUUP++joa+4a8
kIDcVchIDzvB12SHN6B5johVRy+uw9Om2j3MyjG9EsgsnY3rGqhR1EZX/57O9Z2R
oBCRxkZF4ROeCmY5c6qSADiQeCoe2IZIXvHAn2WEA433JyZpV+LqA1Kd3IdjqB/y
vbXG1HGvyBVSajCyVbIAlI6GNgIrfIzoL5ef3+nnZTeg7aBGoctzjxL7pZS3kWo+
uwdo09WqykTWRsZmAF8ZFzb2AHOWEgwnt9FdDtMF6htnzGvEITraEc9fQptUtbd/
e1/eWBQf04s2z3fhLSFzq0Bh2UUI1x7AWyfS0DMGhKG3hxqNRJyMwN95eGTa8ve0
GyjgojDP/0CEN66d30xUz24xkjijuZSgrB3J5u/zQcAmeG/uJwbwTR9D/8otI4dR
x1z4hGHuIC5/ZSXjp3mLtR5uDpH1G5I5eEjkiTOK4qJyjAWTtZ+Of7lFR6TZRLFW
Pe0lF/Ms77DDl+cYjK3RU16sAU/kjAHGmRANhA2hJ0h+oV6NsJRFFe94EG1rxEhR
RcX9F/qqotqmUrVXUbP0EHIrYQQXbjFsDTRp3weSLvpqaGOLGyjcMr3pt0qvjJZE
Uuw8SbA4J27TvrV4H7p/q0fA8gWNAnYyPDp3TYkeJKT4iKY/cEmN/zZIuOAspi+T
dSnArB1T7xirn15GkohDrpLIAUlf7yfiOBZSS13ggdLcK7A4/U+m/JW6SulVxF68
2iJKGTS4VJKJOOSXvKvIwOJIPyMBmFdTdtn0DsvzOsauGsE7DWajnZiaEDHDT2yL
xYFbHv/V+mAf+tWu+fDp5gWSRG0RHHzzr8yGP/oyOBp9HHLB8+PQVV0Kg3hoyita
5yPVtBKoYsWJKoe7x1NbpkZhqoyyFyx4xSOScYOvTYQlfjxEdUGr0qGYSoRAgBrA
lFjWIpgj3DvkwT1U/VELMqwIAUMiu/MlHLlroaI3rcGfNlMdACpmhm8P9b4qBGG7
6dWPDFXIiTRE+hXaoBz15cNkRsTUuiVoi5a5LgIVz09lhdWbaNiahxdBm+u34IVu
N6YxPJNOGAhJ/gIMiFCNg1GSL/VyQuEVs7VYRmh5bn5ZfV7xp3n5LOOFblwTtOSk
K7o2fbD8Y112kp6NVTUsCXPXzlt/Jikeua6G83SRbGlshDBMgB0+0GEeY1xg4iOv
ERiMl+l20l1R0jE6JrsayDzY7m9AlnwQriYEzWxDsZJDbxhZCkobME9OX5ScpD1t
Fz1OOg2Of2Lm4dBEWS6npXRIpwGgX2ztHDxeJl7gO62khmlG/eCpODk8Hjakjg2J
Doyr42BpW3kO2HmAwLgnoQgxAw9GDtexrLKE/Y6NY44x+3nFpPxXS6xtq8e7Ckxw
fsobRwWwue2UT1LAL0bYF8/WKeptJdf3w5RaRv0ARbszrvAp2xuc22IBTSJJagZ5
IlRmKvaXGRY3Y718WYcSMgLJMxnfsGLyXB6xOnbZM1UDcBR3E7+mgiJM+y+P09ID
XwCxafR8k1bh4zPW+Buhyp5hqbSF2nEe1d441SMNTgn27a8JAyf5aSsmytplf74F
q2Pu5poE+n5DzPYWAPNytXMj3mHCDO1X3JwAfAjdJfnhsu0yH+Qiw0ExkAJ51D4K
jFSe1YdIy8TwrNyhD76Rnfa6qCZs/TaOCTaFV+X/+CbsFQ+ExglRX8qCBb8HrGI3
tVnx1+liREg18MriwP16v05nqmYF3KD5VorhdBi4hQmvy7TGziFrSbyG5kTu4zhN
GmdLcohkg6vLqDPYqvvMiz9V1121gV3aDu9BI/o4Btvb5gzuwrltr6qiLmhDzzVT
jqQG6RWJPbVl1EY9vo+ThcBYtT1pz/rXqo7sC0rY8RkMg1r+4d8HSWPJOYocUQFL
w/C77RpNvPZS1kE7yatDgRVbKCj28tVl/G+YzE6x4m1KTXyhbgqqI2Kzng22SJJ/
KgCYkhSdUlXxQrMMlTgHPBz+Kh+MIm7rn7jq2NkZ8ngEwMie1G1zZMb+i+6jQB52
PE5IovPa+WUQTD87kYXy0Q3sHGhqBhAUtqiFyAIYSTN0ru8BDWeiGhdk8TlkcfbZ
Ba3MK1PK0o8eAXRYc6K9V+U2VlkguhMdV/F2ACrJacO8VH/wONOV4mOZQEImehVV
43+6mlfRYFRLxR8uwKEo5350jPH90RjhDv4h4W0YZ7NrTl+M4uW6HyWqmA041IPO
rWUh90aVl8epgHNDSFKmU3DFIUzobddQRfobEFRqssL634xRBJr5esX3lHGDu5ba
8WuMXSKJ/U0fv2czGXZjLxzGtDI6qBiP/LJDuUo/xM0gLofnyePQgfemWNgtwE1J
4kWeyJ7DQbvfGQqK0oAzjHgRx8KZqWgSlrwBAVzOGarhgHgQssoP7yfECmnb9R4y
zKIVvcVfpeIVImpxQSunLRFZWpKmhvt50cQ0/ludqb0gTP80NV6bDRsQXcHodtPX
2CU6eTWX44fsSNStiHYOjwavpr+FmvUWuKnZEec9XA0WNWRpfnSDO7Fb1lYVLgi5
B938dRUKpIxP+dN1C0sKHoI38sOaUww9yhDlsNxGk3UOpr9s9oJ8A6htC31FmjSc
varQDD5/0Mem6UjZ6IYyBIwkOmNlaT+kUJ99T4II3Z6BU8BVsOopFtywsiwf586d
ESb1mPU0UK61xSgjqWFN79SR/B7A0iIV8ACQIl38qQozbPpg6AV2vG8s2syS+Aly
p2uoW5USc+AjsOgdeDeONrWtxecCaKuY5KZ2fJyvAd06ySGPUBdk0njA10mXNe2a
E+Q7JsNpRHdps8roPXG2jAGkYFdv8BLidIej+m6gVdn17NszulxcdzUAwjg6k8zu
FPBDit8hWSNrOxxxwf8UBGlr6xDG50RDKNb0OCEe/OHLGE86iVl6P3O5eM7JIvmQ
mkONM+OHIddUibc61At0iULhd6NDxPPLzGXmsSaBT1r4zkDEv/zMFR6Un4DmFvHI
waECXxpi7xqx6lUqNF/1gBpMIzZLQrqpYrUVRDXXsqbagPZDbenSY8BZcUEyO0CU
l2EL37p+iQtg47cQnhDxhlPKnkvGjWa8NfJ3cNyyn72ahyBBSoiuV5GFA5mL6vT+
uYPq5P+JeXDyyUT5z6jn3jCq+evTbBYYMlRd1zobXlNErwupLxxSj4Q+bdZZxBaO
2lrVwaI5w5Y+XEYNANbEBZp3HabUIVhuOYqSP90rLU4mpty78zoEH6ITyUSuGqUC
PclR0sY+OLhN5JjS2Pqx99gd1/+er6MWrCqLhwhinvEa3BEcKDCc7abFwah4Z2t0
a0pAAfaKP/uy0zAwuJLeaz68YG6zbCur1I0yjxOKNTXMQkMf68oCP3Ov9Rmy2fTD
9c9YpoYE6tC1ISmpq+9VDwoxDZvUpKvv1t/wSXakrIb5iRtS0oOlLYidJiPTYWDT
rVdpIpS0U/jv/Kn5vY9NsdLLBvTSEMTxT0letpWbw5Ue7Toyf0K/DbeUXNaPcrLQ
sc7ndZn53xWmeEpk6qxBpsz+t77Se8OEIgJeDwAyA0q9XXhCkgrXFYXtp/wo04EC
Tof6uYTcY916zMLxHrPb23PvC+WQVyYmTNKD3qWL2TUiX0jqGcEzw9KZZgCuoTK1
W0mZmDTzPQr7twIVXl6pLt2W2hjbWGta12Ua0KurlDZls1xAd1u93vEIZ5c75V5p
O1AvAfaGcXnklzBZwi89CT+gZyLie851gKSn7LX5FCGF0xG3QQVs4XT5gM+GYF0R
LT+tQcDs/m6MFn+VDhIv11Vm6AX990D6wQLyFCE7a9oBHVXsckV14Y3wqzPXgehw
eVZgEF7VtTGyxqsNK/eZRbVFloLECd0G6G00Y5Yt1USN7jCk/WU/J0V5dISfRkhI
Fe16DvXGFdpYlxAZxfvcOpXZk2wNDjwdqgcV0KXqeDQgcw5FJ6bRm5VnGSlZmBB0
6npObJZPa6nrmxEG8yJ+5t9TpPU84ormcl9RsGp8E3fCADZ9sK7R7SovRPqmnWxm
vPXXTJIycn+ZQs0xlfNlykb7dMzBv+IFqlYaBVC0UjnOK2NAbAmsm7okIXdeIDh6
Q3sDULjntHnh5Q4GwqNiY6zs+Q2c4ykPLp6uI8uXz3lEJv6Mw5LVrDTL25CgLZlA
sGDYG5zP/VDR5bk5H/QBgTGSPF7PAEDYBTfTr0MQ9JJ5i920LDgZi8hQ8tCo34ig
U77PahxI0z6sD/kdNSAT7wBlTdAVA4JqH9VWgbnv9XXyZI5RhnRInHaDnGVLk/RH
65hWIfAdy6sFUqmUHxsVTy78ILtzQw+nSB2f5yk2UQ4Qq+lm0CqkI3gr7hDIpEs4
RwSEugrqpxNQ8M77sUhRYLdbLOlaKbQRapnvO5xKN0Xu7503i/pX2dTEP6X0TgJk
P7xJYrdsZu6/AW+6/0LtWDB9dqtP1tI9mHLLwPuqADdXgGxNzVSGTcLLCHq/Dli9
g0iJ5dPOS54XkuOa+4KXSHm2t7c83VG8Jmnrij7BL8yawmRCTjI5rfQtgtBcAZf3
SxiFQNH8Dg6UjtRiG15OZGA+AIrgApenOVI8R/La7PpVZ+4xx1aj3u8ESj3QLDpS
hKjVvCbdnpj4FO2SRTYQ6qmgN3iuHwKPXuRyyP35arZJPWoo/fGA3/mDq1XyacQN
Wvd/NMbL/eYB6Q+gRySWWhMDqFdYpjGhr0RWzlpBZFyv0w3yGdKkBqDhRsXpU/aw
ehJBxQQZk75gc2IclNKQH5zXCwiSh7I/qx1wP2SPwZPvdT4Fx+T/M0ZpbbDGEd//
jZ9NJm1Q4CVWQkFRqqrc5YeFevdB5r2Ev/xFy8HV9Vd8/Tma9CUgjouSwxzsU+7x
UXebv1Zkp0zDkAGm0GoPpO0vGCMBfKIygqsNERKucTox2dNVPRNSyhoHWQJuY044
POvNOdd3aC/nQjYM8iMo+z5FDSqUjKmSKdm5DqbeLy1sCBMyB2KR0eVqdeCw3dL9
38IMvWKV/C7THmoKvMj/L76xzS+BUyvxZQqtxgmnl9Mt5+l6C51Hnw9Hgfr8+gvM
xIJXCLAcg70jdEjZ/kecDo2PQQUE+qyG2WTZg7ET7GZNlZAmZEVawyQeoDaVUUbj
FZwNMoVgtjMbqcB08K8CAmnNIi758THHwGmpqs3eEtceMR4Cxq5uGTjTmLfuYX6X
HSeVULTyo1Ep+R2Nr46SYmwyfJh8jEky6gGUS9duB+Z7ayXCEAE5FUWfKzzd7C5u
q97s5ZyApVnCotDCpUAm14xEdFYwlJbIdaulYCZ93oywLcrkFKBkBuSslUbTlnDt
jJhR3UQ0hzrOhw7V91VXxPRvGewdavc3nMCTjv2wk8/AsKrFwFDiMOtVJai69RwH
VgVk++TduyUyj7p+enyh7L0aPGJe8kbj5Vc9txMKDkBiOORzHfLqfQs4LsBcZPBr
WAuKtHNrsIsB498uLK1UTsDdJGF8wUNMGX72PZ8gyQbKpVovrqHT5XvieZpi2Xhw
3vcc/xTlD0HuWNfrXZvH8tityphXf6PD47kKP+NlxHQO1CAPUhU9HbLgW/dQWLPu
pzmPXI3OP169cPC8neY5Ii/d+jVH6a7yOCQ9y3moRGJC2dWFU0MYNoFtw/uQiJ6W
x1TzajzJiEI06WZ1Jx/K+lP+S4TYQ2XN1FqF42FQmLpc2KsXwG/sUqx8j1SNIyM4
rxcD6+xq5n7DQFvnbWW5q+fPnKElnb8PEtB6ZTXbiw3/zLrImDcEEilctEuOIjHC
i1TWluC1Ceu7934FNlbsI95cDwsMTXd7j/otiE0vv4cz888WjHFBwRU7Mtm3mIzJ
8TUXztr5/z54jX9sYe84hcsylp26pTv90dQIocMRAgk1OMzl1ywRwB80r/zmpJ2O
Uhhj0P+PPIXGiTXhA7wnDF7ouS4CL3URnE9yS/GmGfYh9dw+NEHZaVbHD6DpECRk
fJndeb05KL5LKBtQGiK1Cc8fAZTFlZ/zJx26EFooxks7R0ObEe65iTIS98iR5SVK
5icXZd76hlmpoDdFP/AptrMnADRCeVbSSmK68iZkCa5/jobb06BNnomDuU40Kamt
wMCuJUKEGuvsPNTeWUtBonfry/6Mo9bg92gj0m3XIEXcN7utwQHbsmtKeMnN1QHc
NfvF5cwjlVKx5BlS8OeRY/uBVbIHtx9vljRXPZIcWAT1MWZVHYSuLap3BgPSwkoA
DVvIp9iyXfKEuxJgZ9tbLPhUREkUry3e3Atzfenryp1A6JGRoz46vEua6cqBNDlr
EII7A7r0bkMN6/jbM1cHoBsuKMYx973qvuvjuGH7fuXY858vLSstA7FbhJGS/BvZ
n6FbSpHEOtR3ZNN8vuvHlCnsHjsyFibBeGvyhfjF0k+szC3GUYX2IprADPDsBAjG
`protect END_PROTECTED
