`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yA0cdKni2x2vgbCYYPcABomLwLDFGQVp9ouYrP4hCsVSB2vxyy8X0j20kNh8CHSF
A+tronr2/tfHDoRm4TvafFXlVUaIZB0/mvtAXsrzBYJiVYEsOUGk2+6QZ9842ZRB
F7qB3yq/NfDtHQpCT1NB3cDZhUYsP+e0PG1mmKu+Y6QKKtd6KU/XUayXUahG4Wh+
NK06XIIQmP0l2HKDyUDxQwBQMdohWZBKcKi0qXgfzhxR2VQxuUx5qxaXZYYxV4B4
s+Y7X9+XJziK1uNOsp1ysXFlDpDR8yHljtHUVj6jnhGMvX7Cjqs/18wVGvE3JjPL
HMUUVbP/rP/8sSGFIXhzzT09IPSTUxD8WMiDj7MrPyeyi082dVbUIxpYYUVdK68T
BFPopzarKYlfUibefSN7eOBafQVzGHLQWO38R9xTve6qQDNYzM0Y4my3Us/Jo1Zh
uds8tQdLWujy7S74fp9cdM7ZlOzYAoAb2Sl4yoUhORybpW5c9DZtxPVwZduDuGFq
Z1XopMXL5/qWoBuenoAzzkV9T2H1oreNYYyRI7rGgyWA8oDItCnid1r6cnA21m1i
DDvoEici6Psjq6xj9aj8JI09yWdVWbIZmcnkJCsuWk9ufusIHZYXvlq1leoVsepp
lUgZmyG1VmpRLDKEqZERBvZPJPbYNb8VJyJ7BcAtlrUrChjAXwYLsR/bJWNqyMm0
moOr8EmkE17atxRGQXaxXzzkMRe38u1dDXdGj6vuqJp1AhqMh9NBZi6fk/RlIn1w
rglNT0Tgx/8PjSgnsYb7hlEbfpo0TvEBoIZm/mLlb/Lhtj6McidH8zptDA7TC/QF
4pt/2BkQLxEYAp9LRw7s2esqTPNq1Lr20SzbdfhGXvrgRDcEQl0ZOL9BvbQbXdIN
`protect END_PROTECTED
