`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qkO+BZnIjYg0JuKpkO/e50QYQZIiri0lXl3UhMd++prPO2zKPHmXq1bgxFGfgbS
m02OS2mXsmq5LK8F54exR5nkoAbiwFF2tk8wfRfTv7HYM5bbw0ZzxX/e9+SpDPlu
JyrCuf61y5H+xLDGhTfDIAz8+XMsgSt3JFtpf+BDcKJuwm58L+AOp7uSW+6YQwjr
DktdQBhX7oQYSg0Xxu5KA+3V61q7Cl4dC9/wJ41nJ5SzGMypSiMOXKjynGiCS0Uk
igFj6X0yUlOStwG2LKe5knVlITLNa3muFWuoyrNGyyBZ8FyQiJG7icGqEvIV8C0K
X9N5Fpf/Wg2Ye5/EAaYtWz6U0mDSe9wTW+NH8/yzCVKyPGre2zqvdtFHYoJksp/n
2vGeF63UsWLQQSHRp5Qq0hvPJ5rg5vNvubOEdSpwftndpesViM09GoM1Fx7rpPfd
QKicmYqYMWt+U7ak1uEIoCdxCRP7hs6B62catYoA56Ivv5v4WCJlYHQGmd2EUpr9
lrQaF7xX6n/LcGhay/ZvNmIl9z0MAjliC2aCg5i26Mh2F9xBUkEOc5tUkEYeTcdU
NuvFsc+MqCgoIkHCL2e05EVV0ejKZYTvlgxQQd7aHcaTHiNlI0SmLMPQKmVPwJHY
Dt6L/YsI3zF1iGQo3v/YD7u+LyNxprsnW41lNZsT6x/5UKAyiX2yl3m46kD4kRwx
9lzuJ64LN6z1XEnkbZaWDpSDPgNQM2X5oeO3hl8YWK4NEi0je1eZtDsQ9XYH9D8B
Avfd2+4AIJwL2tFKfjvwGlpnKxHtmg0JFRfQK/ShJp0yGuKVLW7sJNUMSyrCAf5m
BDgGZ1zCq1QRh8rWdTE7QlJJrKEcoWLQKnlFIPBTArdQRVmQMSdsm472gA3osfgh
2oNY8xZ2offf8jR8I4G2Aiml8AYwHn7xw1STfnXOS+I5Pjy+f85hiVgJ+qaxuOKw
EqkJ1jolWpSiZheKo+hVDh+LLoogUbTvup3zSJyi96yTLFflvn6gueYpdJsJPLDp
xf/bnX1QJq/clvZeAKbkTh2jzqMSGYU4YLavob3oWWeN0USoudKEGfvT2weX7OV5
lPtFrVl6XBzaHZR4bz2QJa/KWld/qDp5pV/iGLLX5Z6JeI0aKP2Vrbn2iuZnwqQe
ybTtKxbI5d7bvlqGzB13aC/HtPqLV3echJTmA7r9e8JwvhSFDxmfyJ8eFGXf/uJq
TPnkeUtauzAEReh+f2SQHCl7mHoCUsgJQvyO+EZegwhLaWEHn/XXGGbxokVwMr2L
speF68vqsWoqbP8P19KV8GOxLmP8IsVBcE8+9ObLGZBMrYVmgytKAu/fHbz2eqEb
0vq96n+5l8xx2S0+dYEiUS1AJInGQuek1ZuW6kTGI5XDR37ZsmG+dYWVpaxzHHzr
MzY1AexbaTwBku0pXGIHNjszlTPw7l9k05IdNJFTicWMQN+an1RjxmAcPC2F6CvW
J/Wxe8k7cwrVE/wHBm0JG2pRNa9sK4B4Lethsk1P9UDfDhGTlqDEiO34ZieY2FWA
bd24LbEvRsNt+1UPRgWd913g9m0ovVX1xuo7m6Y8WkRhPPIFDWK/I0HKTm2DFhbh
4eqzSFHQdnY4U/Cu5lYl8qYpwgywndJk86wSdSy999D0H8dP73HrACwGM9Nb9neo
VwZQckN4ou5Og30b+zq6bnry7ChLMt4b9AC3Hg8zbHnToXHsnNkRsDoUGdQAy6Mh
opWge9gHP8bA1nMa8qpvQ8Z3kQXVj3W/174TZR34mR5NfqLJQT/OE2kfq06z6Otb
5w948+AccnPDgNCtgeQZ3VstF9COG2qpRY51JL7QV0k5CReIPe9XUNqcPkSBaKQA
IAbAV9+oOi7xrkX/OmNP5oX8pQdhMGkZKyYypsfh2bfDO6kPGJM9S42GCBwilVkT
C1zV/bdVEN9GFi1+0NXaDQjUQ0uZGzfcqLGxc0CFqBRgJUh1tpngF9uoPsHXI4RE
4RXoookyvpGrFkfXX78XjlPRtvb6wd6o+1QSUYywgk6DmWlOm09l0MID+nFynrUx
XbI4PXfNf0V5cpNF7uZ7NHvHrrPQ7MNSYGnVUk02TTibsIDzlvwXdXvrw1hUhVtf
VEUQF5wQlDAd/Blr6xZuXmPzaz93zMHVoX47fOlHdf9EQHvFuLjJakew3H/X3aYM
dW1yhrt9rsuycMLRxUTS7zaFsYHDUQXgnGHulxxDtA7H1jIbcT7uXWU0zxQZxBpE
jm2CDX85ymxXKCQWm5q5dDdxGIc2LaXeJp+GhjYiN3Xw79M36SsCvw791aJ8Y+oM
fIdD/fctsxqyk3mKWjgVQAOj9GMI+dktz0ZCSjRILP7VlQ4vyLr6k/bBwDpsFDI/
JTtYscYK03dh6DMMSLykvsyGd7ej+zOT4BAaPyq+GZSjAHmJNra1x8ZLBEz9x1H6
TbFPBHdHAZhAlTtU4pryCj0tUB2dMPNJVd4aOtHbYDgtz/FAS5CxfLZ4CBeUgHtt
aAdhW6MU3sQXj4/wB1i1123qDpb8fmJR+HpbVYx+xmST1wjRyx/J4GnFW1iPtVfK
xtnwvQcTcS/aOUUQ4LUmXeTHlIF6lRRzMuxHSd6Vm8guJf+aXgOy5zYdXdfp6xHh
WYXUPcwbgncbJm4/OC4j0hT6mpBFcniBj0+J0hwQeyVmqBjVvbTjZoXru1fvA0AT
aOFXpEfZwj18ZPvZf17mf/QtNKGVtrMhZj1SQ7Apg2HuhKCef9TBI5HmTjVMHIW+
ME8d4ejLtyovqjWaIY51Cp1V7zSmU6m1SJSMQifTSSbR/AbeHDcJyRLnJerlSY5K
U1quosQud8HcDIaFz0Yy9LlczgEmhvunWeVL+Tq1Hy6NUL7Himm5Lw1P8XVmIZSE
74784vU4zwQWhqtJbt8yix4uw3n7QHs6aXmT5e4qghRED2XhP9v4R60Bi2bE25Zi
91hQmFTInPRckTsvCJiM3/2NyzPClujve1++2q68cNDo726K+7wOeBQUOG+MW7Qk
mq9Av26IhbmbmZmlU+RHHtUWga/Ewm7wvlD8SK2pjlIvC6ck9F5K6y2l9kcwOfD5
qtxBfDRf/6itSuwTESVTSy+sIKI9b3WH61zpnj+zgPyabFNZ2sIOezafT3wkTS+Q
4c08haS6SERZs5xmK9TESwmy5FS5O10rJ91nFLEmduPCT82Eu2N5mYNjmIaMYC6y
biQ8Vc8GwRGWMTYeh1jAZ0Oi+TCdc7nN+JxqARGYrOKmndG99znOtSwvlXakaOih
H+CE/q3J7qA8+IfJAYIGqRqS93amQa0hLXsDp5yG00qhGSLCIsMCEDbWhgOM2SyF
rXengf6L3zlpi5z+zNUIr3SjzNrnpqPXk4MwBiTt5uhFuDClXOB7F5dJQ6LhjXlY
S8PTnLEnnZvAk+X0zVeGGm971MiU0/28TyR5s8vY8P3jRt7aIpipVuPmSwwcfoi6
r9nTW16ibdOLLusd7Ejd/SLRnmGmlqBdWBqKTMI/AKc=
`protect END_PROTECTED
