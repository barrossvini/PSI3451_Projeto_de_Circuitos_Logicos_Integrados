`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mbxq+pDO+1gQFBE1JSuaEwoQV6t9Yg5tdtv0MugsIAhxuMPyOrLrQ3weVHwbTzJy
TXV2rj72hTvR/ZLAg5+B5Ou0CmWStyBnSbdHfMo8o1vL0+RiRrRj18XvLNiCaZ0n
0rgOxQ+JpiPINFcfzJ73FH57gzlh+vsLEQZivnAwDfkniglGsYVtDcNJEYP24bWw
3QShstlmTYP1VuDDHFYD+YEem/SmEV/NMcq8IUMA/d+uGfb6BGL8D0qthTz/3qJ8
85Dq5KlHD5jaH76b4mfF6NgqmaKRl2fFrKNpPD826Rjxd2gU3rwO7DeShxRLeCFy
IpztJxMKe9/oYWH6AdSuqQXuYJfPNnZQpUpYCB5Lwu3/SGpxHS0lqOOfO+Yp8Bfg
e/v+Va7vKUenSYrf/PP+16mOmWLE4w6AeHB+uGIDu36rmF2yAB4zD5cHqHO68SUp
MhKZiI0WsZ6wYL5GCUS9BsBripGiQzOKiYxAt01Dx5P0rCRXvvXchKkaI4d2Ubv5
YkQWKmxUgMaKjPQ1ota9Dkx5rog3rPxiQ3aRt0by52vZ7TbJuMSujoo1gQfy/oJW
NDim0zkP+CGJEn9j7Mm+BsrazFLxSqATvNXvls81B5thqWHBe8HMqW0z587ZrcyJ
tNKaE6RtWa/JD6HGDxiB3X/TUgUpahJoUDeY4fRDz/fj6ZRlaeji1LNBc1i487ti
Llq2+BzZG8MhNwHSJ9MWRfdjpQc6gwIez8ovhYKq01GapXHH/e5uZf/Wp+SO+CWI
lLyTOG+7VjSf0/2RjMl8bukN5aV2PjaYZu3f/iW/Ab3fcXDichUNkqt22pU59a9u
0xJsnDSgHJTHC1+JXCzWmRxE36e1MWWq0Moi4KVbCnCVWOdOoQDIpx3Y9fW8jrwR
66BOoADYF/kbrjGn7/bV3dAipyc75Z/RMyEo/bczjOlHr9B96d6HmFS5P6EZP/VM
oe+iJsREt/VqH72qQsJ5rOm03z0UwKF+c879ODY0m5OnIE+bv+K7b0Zhd8damM7U
`protect END_PROTECTED
