`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R82u99EfWzgHRVN1W+9YXbsA6el6/Jz+6w4Wj8GoxSBsJ4rM4s5N7M95xWAwrxOC
4KlKKaBvfxvqp0eR2W22PD933COBrJdQx7knHgou2UED57KyKcw4682BTZqociAH
Sew9DOkkFRytAGpP5zSQLI6GD4l76BHjWoKTolbSej3wc2AJik2/GdGAHH7N21tO
dnCZn+9Pq40XfaLW5uMMchaxHSCmMmr0q7Rr0v0JGhhkF4aPffwm8Bzm0buchisU
X+9djW/blLuIO4F7N0Axw4f9kTiIgff0SLqOB9Lfq/tHjHRWbef4GZUqeukWQaJj
jpTvofKaSX2qjf2wBv32EG8Uw+gJ6jvWkFcGc9eLvxR3d0R4cSc8VEHbg/SKYlPP
gjzY9yCPVKugDp3nFdG8VMhDtgs2h5zQ6kVS3eKgOuCJUiJL9MjuZq0yNSHK1U7A
`protect END_PROTECTED
