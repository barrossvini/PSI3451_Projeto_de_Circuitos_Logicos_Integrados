`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WCr5PqZPtN+oUs71fD5uszdygUYOuihppDx8L8nxzNOn9Stto5fVR7Fbdibi6bFB
vYop2fgOK77U3pRjiZea/7Zt49Rre9x4rJU5q9CKhabKgjsyZDfKae7s7WBh6Sm9
5w8QoOH+tMqVnyJby3vS71xd+V0AXRXmSXBZmseS3RvYJQo1xyF+Q8bAf6sfN+yt
SHi9rPtesNZ+ygie/8uNWmhKdKTdbaoONSvOpYvHzV/p4O5M3L+zHlETvFIBmBJW
MNqkeEJzDuJhEoGGe8oHiaG2huyaJy+7b0Pjh6Pis4RGyccROVL1ut9kGfB1PYfr
Qk+5I3rJAuTSr669NoH9G3Ywjc1RbDiwbkLjtYHgPtvLGO+FOrEm7uargy77D9wY
gFCnAOMt+X+D9wiNNPCC3Wl3kI2SRS/GIrtVfC3Jn+W4WaVJJ/lRj/1np295pcjU
kH7mcHCoL6l58EfpoluM2QC0lWQFS9nH1FdwXF/iJvYKrBTMO6Y9BtvtKqaKvIQe
il0FlAj/erK24f3n1WU0wPLTercwpyTFLD3UJHIe/vjrncP6VYmpPg8pEDYFVnqq
oAe+LhESauFWUnZJgWL4+CScFiCh1gFa6cODu1f1uhhOpkoML0Ht+8TZdCGhxEVS
Ezrt1Zyzrki+tVX8RW6p2oXf27aYwp3fDebrNQUmdzcaQD3tzGS8w9wUW2vrt9p1
7JrgV/EenS6rQ0OFhwYhPfTsZhxgnt5M4JQVzCIuzBMaWMPVP3gArqHToVUEoteL
o2t+qDweKqwQvWauYqpelzGABDpm2KmCaBCtkrTPFK3j1UjipjTNjOXx1w9uKPcN
qgqqMbs5dwsrea4ku+moTK+xeBXP6og4ES/sh1eGcD2TCTQLLKjrQVoz/SX/i6Oo
Zn/dlvNMHxy25H5JdbUX2s03cB2dhedHvrIJndWJZMskQhHSZIe12/kDT9+7bLf0
I9VyFjKqyYduNTpuVK6r/G5zFRjJ7vXQhQPoVWdcLw8ydB/LE1ZfX96yPBt244wL
DvekyWkz2f/kPoGRcOratZPBCdbwPitPAbcuYplNjgUCJlv4BrOwBm8+bFsVn14c
YiY5Y7yp1QZQhm07oAVHvfZyQRP3hshrnPYIjgTwiqW6gV+j/+2ugSEY6tUyQ2gz
MTbSZa9uL1vUbLMfbvdbNC4nJwIaKXmv3mAiwpp1k7YaJNAmcFjiFfUTYyrybYsw
GQIfIwdMGDNYmzFLGzhnyWoxNYshUt3hijvpQlO6tT6rdkFLeGaRih0SHR4QVOaa
2YGbh8fe4ZCYXiyQI8zUCm27k2ZuDVprKOizgSXhL+MbPif1CTAPpGyRsFlel3EO
tsrldNnocpcet9g0jornKbFXgFSeeAvOpyqSGvBDmnpm/IGiNHqdSKUnuGNI7NFA
0VpdnToUjbcpArTtHDfos+ZYnaPupS2ZggdnfPLIyUU+1UDJdeL/kVHizoJa1CeR
W5s9oRYc886W/rd08BmB366PmIs9zd0eZcfPZK347QmMySIo7HPlLHdoxvJpBPPz
b9kOiGZgfCaLJX7njka88yAEnLglAKRsCX0mSfIApzKiQKF+v9Y1a/pwtgJ7+pyZ
8MybLHEaLt+EjxY68BRhMPfqERHjzQiI+8zMVyrEh2dza09+DFUv6bf6gZZylXh7
azQeeRUpaYiCU23DA1JowsXrdOTrPixI9boFt4V78PrcNrWEQ2BrU3LR0TOfkyUw
oOLFlSh75iy6j+rUjBZAUKL6gGROslUd0BARO1Z3K4ZJwaNsTXIflLk5aZVkpSfl
eaBHxep0Jy4qqXN7B2+RfqgTochimg6k3HgjuhlpP6MCXJ8QbA5tdHQv6DkLu7dg
RViVNTIoe3uf2lt0TkQluqFGhhz0Fk7Ktohlg/INHVm6wIKbA05AT/kM1hU16xTb
gar4kmMoX+M+gTDf/R5PlcuSOQinTEdhlBvPFn8zE5kFKG/1Qj3lpOCm1PYzxmTU
P4LDFmsUdNUCj9HGHm93XQJUsbIr7Curfk0QYT3zjZKuoF7vQZ6WlVgaC0f/rZU1
EhcCGxTDMaXKhYKaOXl00nDlNX/Dqg0bgqdrMSFO7V76n8lkO1bTY6AYUcpJM2j6
4ewjbT0RUKq1k6b3n0XSvUR+lO9KmhD1RquhWvqf0QvnPEGSYFSl3ISQQZAnZSXb
MDosE9zs77tRS8KQcE5So5nwbNXdLkTA/kybP88pJwg4Q65KxmqaIe9+CHks74yV
W9Prr1az29MElTQrKgkS/PNMHrXIC2Ou5YFcXasT6MM+SYNo3mgPl9goL0+FyEnK
OHehRzS1kqWheZKj2RM2ZedbmaX5tpw7R8KgAL/1tJ/X5L1pU74yg+HPHFKZbJ2C
awrnwBe3qPeIaibXd4IsUyl0e79OONHUAQvn5FsqZZLzoiWj14VpuB5bSN+j3AiL
jR+F3ehqhzsFZr+PFLne4FxhmTWKwILQWEwkPj4bj+7z2JpAR5mDI7nocd9V46cM
WznM27sLjmNmmLXUDEB0R16dLr4LpBMEXnH1P7ALZmljt2lnMPj+jlmm3B4OOWHy
YIcBnA/ak2zLHuqF2xIKC9QMODmNzXzI+0CNQ7a33XEPqvPL9Ob7NbY0Gu4Tt2/V
1WkydZI22uIL3gXArMIcXuTWtKSzkvldKO+xMq29n/M36/MtprOjI5ePeWB38ekG
oCe52cgnUfZxlosn4weZGxLmq/ZIMJ5qnc6QqsKXz4ZmR4L8dM2PF1KmlAl5aNF9
R86stSn6+Oe66dbosUBOZbG8+XhhrLRtm8ePlGd/wZ0zjMM3Z6kvNLgrETHzZxmO
sQH6vqzPGX+g9PhmRu9aBdWzI6BQAP9NxkRMtdOCD5vkFzApH92MoWnM3mGTOt/p
OB0dJdQp51cRmf9aWkol6jNG7QRGu/9N+SiUNBBoiyFanWiTXvmiMtl+/H5JcGKB
seQaZ0i5fPkpn+I8oNq70mzoIRgTJiLpnMujCHtOMjTiJ1x3dwylSIRNGhoAXhmN
wNMAStCE29dBRTW0dmCYoYK5z0B8zAhAty65D2mSmP+DMAuIZ9/5HkbuSn1UJkXH
zFps1yBdgpt3nEx+IebJQC7+dZMDaLHwEf5W1/aHorILdLfRGlqT8ka0MZiYH/N+
A9/YA5X3zRY9umzKOP3JvTHE+bKriBhyZ+6/B7XC17JTYAlo625Hg7G0DSsC+KAx
h9nFXnUYVIWR3FYHJaygXGLrcuw2eA/+ip5PomY38OuBNWUKG+eCxguxJsSc+Prk
P7PsOu8tViGVursTfZvO7QdH+pDnLFE4EjxvpX0wJeFbbfrVnrzUAeXQBaPOE6um
DsH+dv6v7C5cu0QqhQaxbizMI8RjZz73/ZJZyIqj9tLz6P+3ymurA68XxtnbUeC+
DJkxRyGOQI0TWyEM8R5Y9b2xdWXnhwApJBFk/5gzNOwzKgBZfsURyqHFyzc+dfn7
K/JtKgY0Nlk67IEbQ6XYp1kmv0CXfZQf1GDs/x9jemfYTpnuBqXno+yHgdVPIUIZ
8qS0t7q5pOlKM0XEk/rG8E/Ztz+2Zthqy6BzhX81fPvTId3Z1sOGvr1Bs0lVkhxG
iJTjtTTiwSEVXqoExImS1e/Go6iWN19z/yMsf5ZqgemYblSRYpoZkjKyEpGnwvqt
VdZw971nZO1uA4AGomsoNlWg+vMpzQzmK1QyuWJzpcYvi/7UPyKelbtLUOAYbJ0L
UJ/w9TfWXSG31Jbv9m1W44f+00mja3zVVTAMPw1juMq79+Gf1YKw7kAaMYiqFPjR
FqnCGofvIeDKK6KbqM64tmFBBd3Fe9qxCeTpCgarqRDcrMOQxaQQtu83NzaO8epR
cvFe1x4xAK8im+xnbEYMHAsJiZB/lqwY9sKe6/0mYuhb6WFnAvgKsv6bSKVlwKl6
D/Lu7tzLUpfguT9jrj5yTbq6pQzXkSCwauPHp+PFfWWxeWqZCDliL5C5fHQH91Ae
hZGZI0RvVtWrwRd8Maxdd7KahVyEHgJkK1V1MAtGwcaufPgvvGDTu1Q1cCzFucyO
yW9ckBBrnluCsh7R7J2vao9Vjs8oYqMOIZ3yAXHApNzF2nnhcBZMqUt99Rv4y6Op
wXEbYsm9Qxa6XqiweChErFivJLMEelwO9GL6Py9V4f2ZgJ6j1HqhVh+sHVpBqXvd
e5raU9ZipSATOcoRNrPLHaPc61fCAUYPFK88cDsTPKAzMF5hGRlFcRY7fsvo8lXS
TdmJrEbOjaFP6pUGtWhCPgAJAZq7qPVpoRsEMigEIqIjLAIE26zbH/hWUn7M56xu
jJ1sv2E5g1VUWdj/07AZ+fpYW9KyTQ7dxVRnx3G0+sMaymyGkU4/Kax3MKzm5p65
QQnj8tZS60pGEcPEO1lVSUwakXaJUr7YZplAZ4hspbvm4g+xURaq4HfH657QtmB5
kaVE35qv2gIAP9R0N9yS3Eoej/IoQudw1xjkQtLEgMq8ubKBayBoV9OR733gA93J
TMUOVFcbK4mDiC4fipBBUsp0lHsjKbXveSk78eRyACnMx8Q0qb3amFaHajY5fC/o
8NNgx95+kw7pPd8zpZHtMCeAZOPSooABMG4BqDGbG7elCVwn4B+hCnb2iyQiAz8/
CjLrJe9PEm1/uYQtAGENGhBFtthb5r83aVAPUCrvcJknQ7rEa8vxzWednGPThbza
tyxn9PoIMXXQTAYdZsYkmABYyouEuXwLrhSdXPcD/YS0GNtfqzWM8ongTwY+Wm+1
EgUFaivIIKT3ST2im1Figzgc53pXCNA+eNBRhhhGa1hnoeKGm1rqX4M0hI1tuuft
bfiv1QxLQiQ0u837SKqtVP0Zwopt/G93bB1BVe/GGThuHyg+6UUud8nDW74AgvuU
4JTmnc/cd/8IiQgy1M8S5yHsR2AaBhPAmDgvf0qodacPCa+U/eYmo7R4H8IfH1TE
b9f6IzXNO/KUJaKoyVScftyJUZ6Cz3uv9CemyknLBRL+6azDAYQIzBLe8jdKwqNV
CkB11Bp6Ze7sUnZF4zFQYgA3gTMcQCiEHoB+/oQVbFEjPK0avEFNhbwFrSOXFeyx
+Qf0hSC9tucAy+lPLeuf3ZK5L1ontyykF+Ru0TcLIja7wIOCV09o9xSDz8adlCZM
hHuiJ2bUzUxDOsm5Wt2OAi2Udbgjt2OXNrPxrdnCdXWAN49WxGU/xOZOdg2N2rwG
uaNcvv72Jzr6aL7O0yg7dtOXb84kw7AnGGL1hKXmpVDq7jLXEPQmpCdMjRzTK/65
+Otwb+x4jdZF/pwRWAKULPnpBYmmh4Gnh/1vpN3KWZw0DJmGlTIS+dGZdzbA0cmJ
M4TThfhI41Dxvtahv9Y3Pr6ewxpzOZ5HcYGB8tzZkftbRfBtbpHm+gVyItCqlAwd
N2/fWZUrWKQ3NbN9Fg0LLmCUlzEBE2Rgeu6N24VLMsux2IB7EYr3n8E5VimGZ+3S
o0aW7xgchYsr0mq5CdR+xybo6ba3MtGBvy6WsaJL8NMsxuJnOM5SwWDoSejWy0Bd
aUNmYh7eeNUOJGAOv/X6XjieibBppugwvBPIl2stOd1ZBDnbSiONykiZ/NjhAgLv
3WHbq2zsjXGgeO015EQnEFA/lozMPh3rjqQas1jCQqlLnq/wy940jwDdoZxi4GBC
sujGz4fEAjAjhQKD1LgoDQI0FK909F+E/NWigRYqNzDDR6FmxhQ9V4k20nHEi8BQ
Zfx+sT4roLqDIDlsnuyCNDdMGt9dzIczovgK8JdazrCaUoCZ82MtTdbY1fgwIoIk
ni0F6VR0BXIbzRZEyQOcN70wGi4ztDzZucbWGJN3VLI50Mv12Tror0YEmEOHlyw0
NEYiXo7Oc3kXkI2RquRjhahjwzwuV5sbPor4T4U3rAh9hAmbemnGcWcC3vaxR4qx
E33XVVUugkmsb3hf7T5vqvDQpOoo/DqEZd1IntK24m+TCPViw6i9AllwzO0ENacu
bj8mEv/t5NBZTt70czxNT+wa16bPG1cBUwp/sxnewQ8pdaZOLkLYYMhtBIiaUanw
pOwrp2kWbtBphIA3l/LlbVZrhbsPc18EAsRU9ePflpZf7AilsgJyT+S7WRyQxKKi
9PXCjWfCEF+nJbrziIrglbzcXQWpSzmkqdUumQ7U2ZEcSToLL+0YDC/J5b9ogRs+
iCYlNofHcjtN4uNPltWedl/ymNRYdOhiWQqVl7g2MaP7vb+EgWp+OW/pnxrnG9jX
d+afIhUOxjGjMrIs6wkhNsgvH/ckA5GLJoEyzYmqvV5dhX+ilpxsUst2hjhVc646
GIPGIjaA9wv+ebgr1S/rqaYc3RNHZTtndwN+hDzb1YeMvQ1MoB63d3Cm1+RF8+MD
wZPhojcLnup7zh15l8AUpBAiOBT3i05rDM/jjfI2s4GDMwuyXK7PvbgcnjlkD9WY
MrSW7PQThqTcH8rOfKkyVsAaY4UbXE5NO5nK5wvjYAx6EBfsEzSmn3eZBu+Nj3Tj
liXPjb7s/0LlLa+bshAKc3yaC3VEndx3kqsgrFs+xj3SRVcXtQ+xyU1+Wo8HcbDl
ZbCBRUqgEzRet4bXheOZMgq1V5XKpDOTKCExRMDFxbQy/DaTJt5hUsLFfHV5Js4B
B33x2pyMdSOPSIZNqjv3qjFM4y53jBPMwix8hrZFEorfWZcKpFM2jc80YTXKmp2x
flbIHp7Y1ITvRpiAIQ4ndnayqBEPWkIEr+i+dsgQxvHstKpEMd4vrtO8y9258v+Q
Osn8RAfToTcHtrMiOagmymSzhmRqxqxJXmPo0/ncmjaM2HW+2nkczYrL4lj+BEhA
EwDBZ5m0/Y6pOhAOz5aA/4tJlCPw/YSNu6XkIFDYzAeXBUrHP/DEZ1wwxOkzOJ7A
utapYX64N/ycsHejPMNAD4c3XV2puI4SsJ0F/Y1QHQYGDGDg8Lq2TZ+jI5dqC191
yqRi8qebmZNqMQ/5b79keAcxtJM3k7JbjMQZVTbWF6xvn4DJdxoOXnnxQlRaB9wn
nJsha14Obywmy6Dc1JCOCeX03degXq4l/4zDcFYKox4cp05IeI5f2SnlAPFzRgld
gq/t/umVQVRuTSJE+3Zf7hIli+nW+MkTBu6bSpphcSIEIm/vWs2WgoluvTMxkNbo
cdjf3FGuiuZSfTqxY8+/sI69dMKrqaquIoyCxyz/tLbnTUL4qqQYUkXGGRJWsS9V
PMQxsExG2XnFvV0vWylmJ7zjf5Vtcrm18zvPy26Q3Uv3QKybYayhmEqtIw3kGhJT
+r6N8boonDF4QL+jHvgxgF8nTZ4kzaFXU4Gohx8+MM0qe4kdTn5kyZg+mMABG/Px
fSHE8ZXmD+D6BnDFucLF5UXXX2STvW128hfeqaBRqRc7tmZj4SjMh6leLSOmgelK
T8/ezbqmgE3BSorwM12qfpq5Xys4fmwGefmz1WGNW7/D3l0G3/p/MEX6aswFC5+G
vt/StnYx//OC6krpWsuCd6RciXKjR0w6JqeV4R+jKYL3jKE8w1jJfpy8jRPBNVXs
WWITZeXK2nbrWmdtwHh/52avHvhD4zGTtXby2kOa9EmMxhNY+eNJVPJhRgadYHnR
U/7ETDPY7twhOX0yxRCgtl2USlGXUVXRA7UCWQckQVHm1UlqHzTXWbHiD3kYzr3B
eNYBokLSmmC+S+yL8Tzk2cnl8w8+yugZLMX4UIFvySZRgPa9x3QTWPDooLmxs/HD
Ishr3rRomg6DDGvDsnQd/x9zyk7qWGV8HHOZ2iaYZA9tlDQ4l9JJOJtE33p9/HOj
5dBEq+s17ohX7tyxYuO+J9MGncol8ZWbXzqkgv5UgG3lTsNB8Ami1K3NHEr1KcTS
h50gtqHLSkleIvkRQAkH3x7wfIblKU6wE8vEd4wfZgziZJbY5/vQQ4E6q63gE899
7rhekNJI/FGf2De3IwE6UeBFCxxDr7NZi/qkXLAsyXcCaZVFrf42xNZlR6OaUoHX
8LZI561I8U3pna4E3uRIAph8lIJHN/9Vs6dHCfvhjqazB8y+gihWMvYgiwS6Gw0F
B18q8h0mUp7qYHgyx1vmabKfLyEswHex44K7vmkFkt72FV3fHKoJsxbpriQU+FTM
CfaQHqJ/zCRBD9xmmC4HrEd+PpAUsBE9oniu2y9jCvQZimXpMFAAVh1FRe9lTWEa
c0z4/Eo8rvvWwEtCd+uIlnjXbj+Ya9DfFuyyCnP9Pi8wCzsUXVqIeIRCWt63Y1ht
sxSmZh1P/x/NDGWxinfRCwZ5NYHoc7rEqqVgtVBEI+Xv6jHK/EnDaiQZUoXhxbYz
a3KPSkM7D57/1lYQgIia4kxS5Bs4vSwGuswkGXWgaWFdfe+z6sFzbm/YMx7j9dNi
YjzrALPhtWePu61NKbOy6opiMy8Ho6Sc705jLOgjZDfh0H3fX/HJzCh8UycQVgxl
wX6brD8pVKI3Fi3vso0MvRAI9CQNKLENjORuNqOAyWw=
`protect END_PROTECTED
