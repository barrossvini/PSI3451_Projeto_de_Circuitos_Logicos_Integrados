`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pqvQsq5xAU65JDveUJoUu52hqrhK142JMJ2nMjyfuw9y38npxcaB9V3DulafgBJ4
u78cF0WzMzhlwEoFaioLUY0G4KsX8ChFLjUFJX4+7FLfyMs5RLjC47iqZxhmKg+A
zOThmwC3P3kTfFNbpK2+c622DUiOmUjyIqKkPDnNR+fjE+8fLpPTM/rEIGrS55ty
DmWjwTXieD4itC/YLhjiuJ8iuU1WgEPBERgYRIhT98SBT8Eb6l+azSiX7Nimt39g
yyReKWOnFN0Q8ys7mpCVkJlr6JX49hAnBSa7apK38PgyAoXMwzadDcYI5iwG1Lv7
Bc/coDEoTrD+RbKa6m8SUZW6AdpqZiWZytYiNpuTOpRH+G4SD9W7esGyUsg417lo
lN38LqUKPS+HWoLPVobBQDuZ8NoQALNcnkpmLtZxwgf6trVZculaqL8rUKfXndPY
v8BsPFTv8ELw8rBQQu8OwKleRoJxyA7jPo9gil1BXt3Dtu5iWZQEzvoTiMLCUirC
Th739u2Y0MGVHe/3f8NIC+lqsk+T9bF/l5qI69xUiQbrcZpF+TjWIl5NQsyM9cZr
LzPFrGJAaPKObPyZTrzT1mcDdqAULOKmOU7hNZizqdsszhwCgopCP49JTCOM6twc
aFxMpJ3E3cdhDS+eJOH8n8MUAqaU3FAoOeHCESQqCUFav7hJTv4NQJNqp2OGvL3H
egd0EXSKE97sG843Ql2fngBlLMhdyxnoapQ9HL3NulWwPNu9XpEPHkMT0JsYX2RR
tpt+v/uDBfMEzVbbAZMGNJDzRYJm9x2X0wbbxqYW9th56kT1FrxQKWYYWhdueY//
rDINXayjrrgEvWoSIql858Q3iO6ovsefJ5L5Y0NYW8nL2DxfZ0/VEfP4Q2fq0pnx
cHqRXO4NDYPpn+cbxUHT1HJzsKi6jRikRolScC8loUrjWKAe7Fz+CC1gy0TOZ8vk
Ebx3lhrz+q/xcCKVi1nCZMRfRPKBVlQsFuUc2OcPjVBf0/t2otu4M4GypQC0g6i+
apRnLjyH1VBy17v8OB0bu17YimUd5j8mPTb2wqglBDZfu8C1aEIM/lyOnYzcYI3J
S8FLAhqqLyjWLc3DK/OPO5MbzAT64YMAt2T4ggEfuoc3mPlJHJakcIYHrw5dmdem
yOZpjBzsItBjMD6hk6xc+qm8Ljuv2tdwTiaX91w5LL5IJjkGh8LZ/OsYuEtPNbUI
WYlLIdrCpUVZcnJRHN25DhHQeVLvU14LUpvSWElq2Qr9+rUwyFFvw1INO+805fRh
zZ9UaLTBFdn8o+w0aXMT6tMQ8nzJRKZ80pKobeEFZraI6ltBu/wUhyWYehiru9XP
oQRDjRizeEJvexxfd828y/X/SJKTvkYtIvaWWX2Du/BzayUS8psgAEwJhfayWG8i
pjPGAsnR2ixcgPKHWlHiRwJiBS4Q/19JCRmF8tSZB+idHt/zokc/PhlDR0X7qLIr
YV5pZBkNffnKWWHcdryla/TV5j6YeeR4xcmxicrJaHUNSGsGYbUgdgoIg2jNBrDy
PUeV0Gk5PeCCRMKseEe9RwvISGO1NDzC01UtoKPFdsY4GNjVn+FlRy07chVdSOim
ecSNmGpSO4lW/BRma2g04QpMyUpMgEQ0yj3+Pk0lFBL7SEsKaDH4d3xG7nGJHY/3
PFhFRMqwTHmYnbGVSsxI1oYWQ98Q61ukcstUMIG+lp2xkDBh/y4fXtIPh3+zm4gY
6sW3ESZYU3zFa16ll/PBcVTuLidOzDK79h7k83g/iKRxiIPxMG+0V06+CjAVe99m
DvWoukE/ytJ/dxd+UhJJ3DPNa0xpfkqZ3ozxVQ9TQcWU5iGZ8vhvBFxDVJsORdji
v+X1XHrGcw1fVWMACWBEvGiALd4+R33TJYN7u/z+tE1lbHCAv6PmSEHygZpM3Pgh
syyfbvDfhnPzZ7xxT1ejnx4X5IfNvGtN95jo7QG8YLlSMXg2BtqHlvpZA9zH+rDE
3NuqVlkwDe8CKPrW1rZSnOxsMTI5AVieX/MqHJIbCl5y8eEbaUualjuPKVkaQFvK
xskUNEWOYuL9+HNkxkaUjmd9Hu5fXPXjT2PlhNESXK7s9G/LRAZ/XHCxG7EnoXrj
uj1tJd09v1f0fpHWPrlWdeavva6FOKvwoe+EsyTch1avGu9GQK6rLvKpXrTmK1Df
0Lh+wL7nWn+Z6AAiwoHzKB48jp/IwawVCAn+lKnlIWiqEP3oDnN1BUBNoB56ca1k
2uaMgkOuGY3HjhjJo+2adpikzvZi5L3dndR6BJidar9KyzwsCo4vlTKPMPGBqAeB
2uNJVuDC0qhxoBhi12vPdo3LM2GXasYeSHem/bq9YB74/P4PlDvI+pdo3eV/l1c+
MTM+JY8R5uhn4olu1rm8olDBoSbRB7jFSVFC9bx13WlpH8bpgOEmrpc15OTzPQB2
3Oo//pP4Yvj9EPp9oYyCYf+nUYLjsZmmZJOQKAgYd7RnJUHglkwEFBhqKolGgaVN
tJ6E70gJTcUebAiAwYYOAJzmrCrXIZK+KArfL3n2ZRgpVi73RuFjtAVkX5zKdN8G
2p1niy4LkrpK7nu5uZmiYLBxFGb4asXgVXu4dgysI/bI1hi6RgPd5WrB+5hw1CG0
sjsbS2OeDIFsyXnXz7bqLj3p+bf1NbvNSkUgMpxyYBoC2DzbqNp2PV1XOwpwgZIk
nxZR0O6mh0lbcXse3jUNUsuYRACKP4BC8RkdrJ5YU1dvGH96u395LKlLYibXMCTB
Ri1ZUTRRNZHe72j8XsIMMulITYNAsnlC9HEwA9s+DE307bZPte3DUscAB1Er1kgc
eX5Q3xMXiIxCeDjaHTgDm8Ocu61plXfHm6nSMJQMM6kIn3m7rzeKGLktwCBkKzgi
r/sPnLwvkdg7YPQKlyO77R2+uTyjCUXXXyI89hD3ZL/St4jhMGVPsm020r0fV7rU
TEzwyeWCfHpU8U1eiWM8tXjYIO3Xk4xekkOCi7HNx6CRdfJUNBWDzl44Dz2Ft0po
pb4JlDh7GvETzqgpV+y2IQVd1eKg2NOMIgmQJ/MRfBSZ+WnHFtuxvoIqL9x5G6v1
qJ1s9OIDoHwO4VrW8VT1f/LDUPv5RcYMjWaKvNGdc6Ir7gj9sNRxR1Xacg2X6WH4
/PPXbJ7QMR3VZ3G/wUK+ae8pjIeUkiTxdHBIepNSn+/pyJFuEEH6VHQiS7xZuNc5
bqvfJ4L7KUKdAzKUmbBDazYXuL7/gEUFwk1lqoIlLODCJ0ViFkTgT/EdvvgFETvh
CCKCZHmmWRiZ1IKtu5x/XA+REesb/jg9oeJL1UoeeQUb37TnoBUdAjm1EoWqINop
zN+l8su75+ABBt3bf0y+x2jfeE62i56s7WIFAA4idUQRwXxo5YD+kbpgUY94xhB2
ud6cIvNUnPS6VKwYbnOJgXFZNZeGziJiST0Sc5MOVOWPZkGTe0RK2dByBDH0KQ6S
KztMvThwoIBduRdWXy5mZ7FeiXMm+0ABgJnQIqiceNojzHuKEfjdujQoc61cKLZ5
sXXBGRilJbvy9cPFjEedOryDQnalUZZgtchBqIspibw82bcsnR4X16hLMqJHGOKt
dpySHfoNQacHrxmSqmfbS9BZwtkUrQ8xkwhJFjIZxNHPFLUDK93ifMsX0GIwGW00
vsgLaNeA5tbIe5qhXWBfi2Fn0tzVeIh21nO+oQNS5YLiO2iKXjl/TzIlv78Ncdeo
ntZaQ0cy6wui/v1xj1K8H0wk07VU+CuDgXMm07Ar7kkCzktV+4CTWJ0z/wzRof10
oW4pqLcIv/ISOS4niYxoWagNszBuWGzZQ8QrXhEgf6fZtQ9z1p8EjguOqytbujws
IMrbxtb2Q9dTMTIq+cuKM3GLrVVhj1RWi6s+SwtER8hKepGy9BZh0MsnGoQVo6TC
AOOslGIAIAX6aaDAa2sMODOcNJ1Pjk/JSbxD6Tzof6O2swH3rqI3JgyNYo3UK5ue
F5qPBJSK1YQLe1MJwMttUJm/qjHVM8KQROxmAfXi9G8MxsC+Nhy8tU8jEmzNYAKQ
vix+Ba9tckvEFAGDwlAlgM/q7TtgRglDLo3MROJ+mF6LuxcwSNsprbODXKs8k7bq
Xksh06u8VVgApbiM/Z+VMaB3CFZCN8jjLY7Y7ukRde23buovJMAwkRNtt9f3hvH4
CM4i4sw5PdlTi0AEiZX/psjbJFx5Z6UwL5QhwbmK+q2dSafHmmmRr4Rk+fwutGcd
sGXWGIY7lmh5skox6ynFJ2wVyh4UvNA8hZWVD0Lu1nURIUvXyvfXdbSKzu4RQa4R
MKSak9BcF3FXvscb+spQPpStuOugkSmOM7ZTlCMV1xYfOrAgdoNVqmI/P1cNsNea
KHVAGRr80LSUykp1Rrzdx49JUbiw+0UeO5jAf9wGyvcUZxoS0FIq/5H0iLhABgAM
7iq9acY+W+8UlPjykphNIMjvmhdT5x0xhBinYNBrroVScmEILtoljqbvUx1UapWT
gYCzQkfPee+eAlhQXTO1gNrjw1cFVTxjwmKdjrOiP1fLK29PyT52jz1cWPgINQHB
9eqReB+y/1YZyZlBuUvI3vYQPMyTM52KvfvxyZ+qWS87iEv9BPphDIAlqzG7C6L1
tzYF1nVOGGkWS46CRlOt0hdo84AVciUTBz6TviiKE5KNUCdJpvXwMgQKbEt8B5/5
1IVALnMVmyYPOIQ/MYKjvhxK2mu4wDbQXrTYN0gfUR5jLYcdhOi6/N7zRK7+Pue7
W/sT4sUKtFQB03vsctxcXQNQnR+AgvjVxkMfv/xNElc6TRbnRSnEkmbgJ+a/K1gy
SiR+Ih1938+L441zh0OvsoLWBfi+DAqzBI2/1BHVCy018wGjJF1AzMgerlkITy0u
PuSjYklGbPISnFwbnvqCo3xNkCoOfdReZ4GorOzZMDwDA7Z+sg3D0iytzQ02VNqW
J8ZbK4OIBFDszcwgR/2tKk5b/HRdROyZeFOL3MKA6xCGjS8daj/nMxB7OtMYFA4r
FPrTrUn1oeflsY3mmyVXHkAJ/WlUKIwkZ1TwYKz2dNuX3f83DuB0oO4A7aWuzR7Q
HHIj0gq2FiuD/ECrroragXqnPxQbBzuphYS8GxjzZw/KvZaJhGVDkRklTKv/bMiu
rLgcZ3ouVcURZIcBsMNL5HeHQZUiKQuIESDTcV+3NTeZxPinbCizQOuTfO9YeRNH
BWnBfg8M6xL1dblynN+dis8jrKxvAkJftWALvgV3OYUvZSMUx6Wny/iGLzdeBrGS
MMbYRBzsx/vsjt40kYlf9f0N8OEjL5VVl5A5Lz2U0tkIFuy53xZ5YZ0FzOihwMb9
zBseIkSUJiYUiPVed1O68CflKartjx1D0aLYgZCBJqSyzHTRBtzPAqFc6r7PI+2p
WC3XRAzd0cEm9PE/DA2W/1eyFbFnd+W6suD+7emrUCJBhlQ8mhFfkJAPsphEfnx1
JBUPRHfGZ45PpMyu962IAqmIS4We+WpZfrFvkAbjdZsK8pIdnuojAnfLSi65RhuT
Kf6le+NnnFbKjRyVyNKOfEhPgAb2Hy35eQPOsJ0Mqtac0QL3I3f8lwcZKJ+8QD3E
fgu4KRteej1Mmk7aIy83GpWANW40rXg25VhRDYfX9JX7jsOG+ZZihSS7U1eXplNG
0ikVQetTCyic7nwV+kdY4N9fvh+CyjyyIGvFfCM3agT8P8x+ff2gc71P9cpnV/wz
W/Ahbx3gPi7LW6y7/fH6nDPBoI4agWbr+5XgI6YD5DWZocFuvVJlkz4cftHYwljy
bf/9TwOYvZtnMvdYbmhxMPKat8J/uqIyT/vI8TCBzfVuf3Ca+1SYV+f/iG59jwG9
wbP/he8aGDXbIfyuMCktC78OW4yb6f3p8coDttpuM3j6w6+fTPOboHyFFUIsEdVG
3GJG+Hk/BRkGv9iqGS88/M8+M01T3Wq+VRqufjv87qg7G5ExfDHDxyc/d9L2umbw
z2q80Pzz+bb5vYrzhf/rGkVOr6/eu3wv63gVmwgHTbbRGSdalF5mvn50h4qkaOr7
PPJubuUTM69nhZLsKGGY1+Fw9R/N078Y11nXa68mDxznouVGXHfokiOOVEoDmeGv
Q2s+xAOci3zf/piz4OLU1uLfcQFGMXoieH5ildCdbtX8b8P4g38JSLlD/XsLLGyS
mtJ10WRftx2KGRito38xl752rOdLWxxBt8IKx+PAEuwkTuBK//et1oThvcS8De/X
rQX/czIByl50E8PBmHjC1qsIkuZOvmB3KC9W1xjsF6J3nRjNwu9gndpT9FVJXUo0
lFsqVvLtXiBlto/hzjeD0fHcIrg6WhuwqaSrDZw0tr3RE7mwBFfY4GB+sci/aYKW
NWoLF/8JGABGtd8h+Hd8CXeGSymUqueVRKAkj8p/8HUdqCobwED7JLm4Rdlh9GDZ
Wodng2PHGjneYUJg5qkrsPORwE3cQfxVk7N2pSoaOmQAnpO3CJP7q8IJ0O5HGRK6
dxQ+/YLvGX9dv4biQPdWNVswLBmW3MfUueKqg7Fjk/HNFpc2wUg+5r6g31El50CX
4naUiFptJ1M9LDZbZvi5gab1SUJ7I41kIxNmON7Ul84I2zXCeYwn+PCNaH5ZQqDF
cI9Ew1fQqwRbnz+MSj6+PcelqhWQZIbvj1U9GuZ4IYP41v/z0b7r3dLUzj1lzeFx
LpJd8SgjCyMMv7L1IIMmEeV0/V+kzBz1wqubIZy0FxJm60/g3dpIMI7qhQXnK7KS
ONr+K5tHHr3kfhxOe+ibCBzFodphnN3hsOjhQdpadrD0vUntgGOGQfFjCsJ6wzef
CbyAdqtPfoLsIm0lHrt29WXIDEh9MY+XZhkZf8A6Ofo4hXKV2mVrnJOgDyxPyU1/
y2j69Ph7AFA4QcXf8+ZEprozi+E0iLC+vXeoh7kKbmxFUSdYlhmcUdYA6P8NyJJS
hpZoIG25VOBZ2znhHyJJ3NoUk35zk4UKpX/YZBPVLoAYtMSqkqviVDqkJoTbJFtH
tnK7iabRQzQp/Hjn7ZyNlC8shXKkbp68CH/qlC2OcIXhChgOHBBfO7EHbjLrSZn8
ptiV9gVXFFjkfwAjoIxRJi1chpK98gN8wlD9N+9JhaP4o81mvUtkTqRSo+MsGfqq
rAfwiGADK0ZryIfwCo1/VD7AUiDMmxiekzEzMDtFHsmrxME2RzNIuIrIDGVM+Obw
yhRxPfsPb75QG0qbWuVWu4eo6W0aZDKay/2/vhTD4AhzcZzmhJ2pNqUgvdn5u4TW
kzOKNuk+9hf97EhkSb7QS0LHLHvdPjMUCtQguvIm9T7bLdNLBjKJEcxgfTwTwg85
sWIFv1wZ09AzPXIZaYOUxe5uh5MNyfuRZFoth2ZSXXyfdZCAVeUYlR2/qa9rnxby
w0wpSqV6rLS4JXPz7eT5wvZuK+mlRuFbb0WajiSP1NmKcWggarARn2gJvWH/Bvp5
+QagQLFQUU5kCgUUhdJ+D+rMHIeaEL8HfCOlqOBS2afb5csMnrlRCnDDxg6tIUG+
B5nSIFiWM9yIZ0iQxRjS7Z+mzFgwWtXvXKVf7/uDZDmicZQWHydxEzG7oEl6gNRY
Ml2/I9LHsqf776wsEAzPQV6Qpa2IWzLnsfQq7lSm6lRA9QO8Jb/iwWdgo+cPmg8R
BIPrXdtWjGxO5wLe6jo+XkdEa6MjXfd83ouzIbJCPgO9xAnZhcXOBADIzhDe9vN8
b8jzDXCWat+ngTofmtklbD1oAOgr1h220U2Tuyo8bem8Wbe0rp7hcq/OUnjM17VB
f5m9zXXsghtmVQgiC2t3/l0GAItv4wm8Avjsg66VuEfSiEoMzIYx37+3x2Qw0luq
zt1oo8hsR3uguvi1TVDNO6bzz4oTxHKyOCxxTKRp5cAg2mZ1Bo0SrJHewRkyBavu
8p02K07kg25Nwh0jSyxt3zdWv4SthINDmLc8HTaKoLf7VcmVG2WKzdmxAzOxbkAN
0ReYp9iJzjbNPXL9tDM77gwqFH6n0m9myHhKqTHtasMn+er256Lkl4/WnULpxEbl
CiWcxOXGZ2yTInlItRTJkcU40XBCbGrWHpaDL2jW1FLCmIBgfIyUanzkz5MGaO8f
JnzdjTg/L4qoyRF5QShjMyaYC0rjOrJQWO4LMYTPTYrB7LACJdwsWsLBIl+B8Uh1
qg7uVzH+G9m70TJQqQDvOaoMg2eFYc5XfWLvTFoYzo3+AzLhI8NT6negHus3ZV7G
7wE/KFWwTRhsQVJTYrheoD1OfdiWpvIrFvZnYiDFyTcFTXexf7y6/fyOiteeQZjS
xL96clUk2kzGUY7wtbzuwnFunSd/FtgeyG04+KI0pgVOUxwEB3Npq7PTBzgbSEMc
ugdHZolPjXKm8xO2Filoni8Ov+kNIykAtGJQcn6BjQoYlWY6Lz6ouo52XFi1mvpj
IkQZ+MTOfRFTgBMDOOxehs8QvBcvPwhB+2qtz45sOnHUh8Y4SEg3TUDO6nHu/NH9
zEyb/d9M7UkquxgPSGEq1RZmGhwpBSvk1bpc4gY5f9Y9aMwCXSop/UnXUyJ27Mhk
Ub591R1FZp8CwmFK2LPNVSuYdDMUm9cILJYAqcRE1TLNWIqvPRT9HTqBoKsk+qJy
1vLeZVBIroG9hJ9+42VCwsgePbY3h/jT3MPkGxJOlqjTEbS8pt9JA8pd8v5kVXIR
qFrHjALSW+w0dui4Uf2i/4nfEbkunZTWwNKeWJ0Ri4EIUGReQz2t6X+qoZ49Bap8
O+IdS4HqiekZM8wC4dxKV4wrVf++F7HybjvRoOrDtM1up+und8O+J6C+Ush9SoWI
DIXXMxS5TauG2yZ7+gh1UlD9l7G+jB0wWr+mwq4Hh17r5LtRXXiwIwmVqyY6x1Oe
29PglSXkqWJUVWYoQkjALhHcsNFAEoedFOUP1neNMETEbUHjaUGmuB0CoiWdoUX6
8usG4OanRJ18EoaCpZfVn0J93dWPjlH4W03ZeAxQEP8VRswANgjjDrB6g2NgIZWb
bcp0ewq4hCB1I5jdv7hhb/erPxwWSem1G2EMw+4xKs0Zu7em2looA9aKJ2ArSNkv
iyBjvp1ye4SKadrkpzbJkkeipi92Wa5cV8G0vZYpK3nNM1o0DymsoK76W67mzsrk
JDg9gom62LIuR4AAf7XmhwNkNX2sKyaiS06Or2YKQ5ka8IcuYIH1+vmlPU0i23C0
JuShlvM/KA6GwyBBSZBUE/gmPy+PstY8kotA2RHdylj/X7/8jhjRgHt7jCfbUMyw
nGd/1wuTLhIvviUsUOLyp2U1tK7XxwYk+c/6jZMk9nzt34TSzWwZz06XwEjeQylC
xcZRfvQlA3mRSPmM9FXF4YqHCUGhyAb/RQhb9YNQj3mLod2X5HZwAha8y/FIFImc
GjH2YjrYPy9KwoG9lGGJ+ijsjikrvMM4cIyyDdcxswcFsw4c4BOyNoSa4T9wB5xU
/9hYSuLni5+i5mzpX3bl76CizzRdLuNPXYwBF2vQVKZpgfYga/brSlX1pfALC3HL
j9vUJfTlr2CKGUJnn4RwITEQbFLEgxDTRbTcjetaY9UKIOfajit+bLfEvYmkZ1I6
WlfkOZmm4wDGkrQ41viCgSmIf5KCFv3QiYaFL+laF45ts2SE7yTc4ZKNbV3AXEHJ
dzD9tMOqGJjPUKJRZWoKoVSxULlI53JMUEe4vKyPOgABnwlD2T1Ksns6/Ol8j1X0
FR3j6JkTmMnxKQEd3PR3miGZN3gGmSWqxvPKR5jSUJ1neF+BHUh02PKyfE1QWPnN
12VqgyfUny5eodQzCiCZZ8T/nKJ+Q2+kavLEk5PMhXMIqBFuZzAHpxQGpFkwrGXN
a7/kr7SZSOS92U0nMM2WHsrf6zrTMg5ZxL19tdmF8MHi98vzsfzz83Ln/fiFX1Un
sYgE2BxOD1989yPqif4krMkleozSGikJ7dWvi85Be9qqBrDbs6JBxZ96UxvzWMEU
96fnjbow3CJUEkhhKfOCbS+UB7IEMNRILtNHjcABPsYRDFkjKppR2K4HotmEuQZx
IGygFRv9UtTdAzS1b6ioqQsA0W4inq2hcRCMa1Ogj+JoFOeh+GhIAlIWki9L4Dbg
h1sAMG3DG2u8OpG+21/vVBs1WpFnX302+LrR0IiGqzSPX6GT1OUwraMK1QyI0yU+
UC79m1zO5brIed+/t8miVTzpyh9xQ4f5+mEPoXZMf/q62oD2Qf7ffhpdUnF9RX/j
wWhZlWh06EKt0oOZQT6cFF2FUAdABSAmITVA58JF22U3EEGFwUaL2CSVRlHah2VA
PKBKFTAewX0zmyneZdbSXHZ9U93F9MtwYMXJ9nAmdsFkG4uINIQi4ccZ+aXNDzKm
cxCgYgaXHEBXJxYCnvnfEqsruUdmDE+E6qAOsw90ZDQ1hjPTIQLOaQmQg2EUpkcF
8K6hRRU2IzDiQMm7NXtP87gq9BpuCIlI69zHJZ6/OeQD310yCofeo7az1MWHCzQ8
p2rNjps932v0crELGjgmNzZljI83X+PASG1WZ6nxJ4VgQsk4uzd6k8gRT42+OwMN
AYo7AkmJ7nnFO0oSL6UfyE3bKYgnsYE1L/OQ00qTfPGiLGM6mKd1vnehusTt/vJe
HX9Gjsq+gUFxqg/fXSrp7OwmMax7uKhE0IcEMG4WpWyO5wa1ssdh7P6jUoqxFHJ8
I6X/ayZ/Kv93asHenlJuqKAG32rbMGcG0Z/Esv/1ZobmYBeY+CSAoj4g0kyCRS2H
W0EldVI5tsWatfXeKHCpNp87WkFkNmGstOjXDR7EkSMRaAxRQLzLX4waSIN7ZnGR
ISKvGSEC6Ee2KcbWmk4/bCbdwlqiwxjGX28zF8BsyQxBe/cC78L0rOX6UhOWTv4e
ZAlpBfcTH53Y61HKmJ2txyy8cd2ucEsZ1ezZDHAJpIbbe9MWWdn3L+Yaxr0l4H69
M/BsdrqEX0jcBLBwlt/48J0jRxoRtE0lOwZ1Yuw5mDfjimbextGa6yuUOlAlOme0
VoG2JvmP55tG75mNKGgcd85vagFUBup2hQZIhATCxHCyeqtvWKHojlalhfXHOxZ2
LBz1xyDL8pzTw5la0mULLBShfWKKtCvg0pe0n85xG7bzeE3YG1Il0NRDcMaMBBBk
qX1ttRHrouTowyGfpznqfmJwk4nJirZVST5bxDgP5uXhZiH6OTuME4PXHgYwBaAE
E2OEDhYNpJ00HmsiEQpCcusIPCMaL3BZxH5IbA1YHUtGsn/KOTq/XgxqxDNlz9X9
J0ZRz2Xy/pbg6oz72hkJsr+kb/RfYXDU4nBdEjLXp2dofv6nodCINLpdYCaT2STd
2BcR8G18td5wEAS5FGSMNLO0XXM1Xx0AQpFh1n9H1sIC9ScSCC3inXAkZaSNANNY
wGFgrbBJhtdz4LdLI18qzbNPh1bADFZqBxPZu/HsFKNEXr/nW91JXLSZ+v56NdTT
nwzycfzInOVtZuLRtY3i29XW+C5cWmediU6XP+gD5tlU2C239S566uKLkw5P35lV
/TwotmIYGZmHrlW0rWIWlkqb3wmUbAFELZikkyZ9aItcT5AiGqLjgUBm9bL8Cblo
/tOnwtFFsLeErnbw4nnmGbhbrpgL/b2mVCemR84y7TvPicgDBw3xJHjtkM9h1aYy
GswdCIaQKis7tW4KQPUtgkkugZw6JbpfBdl1lTEdgE6OEBIjoGOFJDTS6lzTy9vp
SDj+dVkZ8ZBsr59eRKR+NqfyKwNa0c5qojn+FfGSeaL5lln7vPsWR5TEc+G8Ed8W
tibyGtTpqXa6/+Zv5sW+mZEkfp+rPKnffx2VXERoElxO6dXTeAphC4mOpyysV3m7
r4xDecZdtIEWHgWuZ3B0/809JrdkrYav8zqGh/OMBt8CzrZL0xXVuejXWfFVzm8K
y1NTew2fI4l78q2eCxqnVOaAwD3xkDX6abuESyfdjWaIyWeuJ7MZKwfOPrhJhwub
pnqsLlqcU7p7NEJzLFoxe9Fa0JuhYq2RD5zYSMFTtXmPQJbEX9L46YGeMfEyQEvp
07mqdnwoQoYWMXELXUWO/Hw0io0jgYPju4cidgSnIgrMnIZH2s93c2OOAoJWl4zr
BIAeuBAvOg3FVbDbE1y3V7a9isEwhqwnY1vWc13U1MXYP/widAjqdTQzbtgR9sIW
Q3N+PtUi0UEW/xE4OHcy4ZUV+MyFE6MWP83GK9nFuc/9kTG75g7swIk7eksdEQOC
ByNGsp0z6cmUq7lKKsbSygG99xFxVZxi9e4dwPRg0TzdLfS/gwZjy/dA8JSEcw5d
QGGP1yU8ka+FuyuECIM/jeIiSWCytg4sRq79bcyWTZS+R8QNzaBmdM3mEmtcBQ9K
KcxoYhm2bQ33Yib3PhGlJK6Tl99MITJMpxZk0dNkq9n/EKne0l9HhGz/HJdIYoDn
U+V+ZdrW+qMnativaRQFBccq9oG4Pnf/YIMZE15cxPnT59UrAPdeCFpWS+fb3OeJ
AmClPr8vUvOn6JWXP3k3Rm6IrNWMWqs9Olhif1G+mwHM5dSuqnCuwO0g9h34jeDv
INVw0qVHSp4jwSsGDJK2hqOEm8F2k18XUj/r07lLUTTaxqHziikdqjZmAehFwSEa
YHUJLJGr/19X0zZGJOiBxgkwUQcuZ/FKDZBAxO5nsWqP0bh21NWryo3fTBjVmScQ
JtrD9Zlr7SnhfQyBZ4ekjACBYxuUCVDkKOmk2rkKam+rphbJZW4f9XidMZL16n6b
ziOJnpc5czVOORbkrnM38/OK0bwSETE/iQxJvzrvAQw7pMaD1gYQUTuk/NodpwcO
6UJ/RVGbHKTG6i5xLMQDYEw5YLiguodNZksdb409KeWPi/egbH41R6GV4Ao0JZ2Y
fP9h+euWwrGvC7BV7zEFYGpTDWB72g+nGZmtchot3zTiEw1AVuQoUf10cPILxHOL
K+CGFE2jGHpyPvYDwlaa8VYlv+Jv/QnF5VeeOa84S4MzyCekXZp2P8pYhQQFd+Ln
LkCwCQXTYRwMhj4NeZIv9IM87QqqBCxy90eOS0uIK4xdEJQ71Ws/yNFKDS8+2htK
eXi5AI0SuBxAMUxGlGKrM/M59E5ayu9HgjKFp9zpx9eqv3d3l6OeKokx4+/klb7/
3RgkD+rM3lQaFyJ9PcTNQhvqyW7HM5wrfnLH4ZDzYv1bl0Vgc1Y9LyZJCsjXDU9p
7cWtgLj+lt+xz2if8d4JPvkLQwvIK3UXRzBQCwR/KxhNPn7FT7ZbFZHYrwfHO7v3
VnnUdgczPcWkUkq+kLVe45Bx14WRTcDNoLUsw48hOK1qvdSCJkM6ApJZws+nEHr5
gh6Arzy5nb2BW0xEI3H1enrlLZX0H9y5Zy4q7OnLGfF6MIjo0PXTnEYrXWMhRxJz
s+Q/hsUs+bjNZS14czFBk9f7HDORC2SZPsBTdxGmPiH/BXVTkFTfBnhuV5JRXQt/
CL65261+MzCmr8zHH770IJn7djrqHeh4AYjqQW9bL2zOdzFwqCbm0iWfGX52eA1W
RDKTvVBwJeIOwbyeHtOph6KosvNCJ83OMH950sNs/5Hq96vYdkGMxyfriLJIX4fn
EvORkLqjTVUBDE7fXpCeU6BYyM6W2d9o6VpDiKqorh4itE6JZ8xZjdMyaqEqAb55
c0H00/khw8HKo3CUaM7AwcSP7+wxZomTpdONmD/dgplGKSgoDUoGa/fK5qHaJWgQ
GXQvMlnD5AZDY0UF/Uqnd+ZewELjXvtlTHQGhsotRG/h/yFOtbEnHz8psZQs+pyY
n6aiNXIxVgbz6izpTpE75W77IQ0rmfRwwLcYeFgKfkTzClqRgs2gcrg4YdWa+2PF
VHKuprDp3Q5sMJpMtfOHQ0PzK8ep38ztJ0DoUjRsK7D4HFd9TQkhMD4q7Ws7CDF6
2wKtV5YcEwU/irPVOmtiCruSPcKjKg23ZSDYAGZUSyL8yjG4brQgp/bJ7NgyBtjD
utKDsUj2O409Stga7iXvLnBytkhZDUjei9yvLKDEnfKSe/Ik/wJZjrZwxpnBM5JU
4PolhPSJMHf5oT5mWTyTTxGP4689GYiud+c782TmE20S+A+WWIXKv7S+XTPXksBD
BFzXXGmSKn7lIEJDlLkdHEGMA5uF+uui+RWttq88TdsaxngFrooBFMLmAu44nfRe
okrCDm50lyEJhlvqKQPUJEqeSvWXrSinsHymhMVhX1KYIfTp42zVXTHRUth+La3e
QTEm1PqWRk+6YGg9tGjG2z4EtYq88URc2l6SurOyAfemot2AYzWERckTi17UKdLt
Jjpppjzs0HMESz0Zlc8wNsjY+47kdWOVXkPtIo1fcNHKF8Rc2iV1dnTPiMGQKR1i
bUHMYmD9nBhDd/zhIzJBs53qe8pkgW4F5QgwN7f5Ck5/tc1x9ahS5S4I0sNlZU+P
gpqf6lJgM4xijvTr/NbjZpxFZ+EXBAllHVIYUMHd7fL+TG1vg5jKVjbZNUh/7VC6
B+uV8ertmq7+CNrxzQXgrLlE7C998BTHRyF6BXXn+qJmf1/N4efAM3boR/JYPuiM
w65fyj4r/GuLxHU19ciobSUff8/wUgzIqA/ZIunoa54ewXBfYU3XA7GKo24vOfPR
NQKJ7nhBW6+c7NbMtQaruUShMAe/TDzFfSRwj6lx6i515udRZW/Gl0aDzi9gnC0N
VkuNQCU6D1/YVixGG305Gl3n0WdnecVGLGdy2AZr5Vo9GdWnfO/V5JD5C/0XgiWK
Bew15fU4BfVGms9zwh1JtKLObtnTAVCvUuR4TMNRIZbBQpKJrWK8hOiJFneUCf3+
KArTlWoIXASZtZNMFt2znuV68i58NLHhu50PCQQi3KwcGBWgvkF0b3riViovEx4i
qovP8Y7UXu5S7lFBEKVxIBl9zrOzCJBt9ye9daBm/1uy4TISv7SbDf84lD+pTvU0
DpoMXGw9HAzU+XpJmdl3MYB3Z8ryM/WyC+IRtltHPqhqqYeFfPKsZIL3pbGuJBBF
yyLrTbpoEqav56JhcbCCmi3smXeeqilpShj7w8ZuJ7LrVXutPk7mB1YyyYCJx3jY
7F9pPPWCwe7HN1aS/738DEdLWsa3gDz/nlWcUPPwI1Wlj5U9fZHe9PPBrLLmJrlK
Z81he/VymC9h8c47W62bGruNPyLCF68zAOcOPyindu1G4ZylL8z9oEb+RCoNQKus
nNYodzu1ONkb4KwQ5/UI7O9nXE+lFAkmM1JRBDX83VuHx9tYXnFiDutn+wX7JIR1
yyD4xXvi8X2fFpx3H9BPKALoFjj+kIYJDiWvuGOFpepBp7PBKGJFfVh/1X0zZK/3
DQbKnzQ7qrvWawg3PNr/Ib5aZlND3TNciF5o0qjMPWcSE93QQV/9C9Y8u+JXNmKU
M7Q3T/ds0DBHYl4MO8qbpLrnFpG22ZhqZhopzNMa8qNnl9gZEomPh9Od1/4HEERp
ZBM2cLbVAKVMBT+EfB0n59FqBGHbsJBb9xsJvkenMBM9HwxkQBhhuVzkDamls0pk
11EYh+Cn7YJwG+vBTWSxGopKCOSXRNrzysN1iFkZcKwkeeJhbnVM/lLy6XrvMkM9
mC8oOcqvwySs72oltVzRTRoXeItXNBTIP1Bc/jShItwE1tWMc6C6CDN0L/yhHy3e
gNzgqiHDwztMkfeKgVIJEgnahyWoYzO9DsG0WI/phyyaeLTOSn1wLEdQQ+DfPP0C
gLp8ZCh8NnnRkGQnUY/cnwGNiHHZeBzvz0Zcy/kRe5NyF/ODJr6Fi/F/M66WwXNF
gV1ty8Z1P2zWwzp8VfTWb4Rc7IwACmPfFeIJaFp/33DsKT/QH5Tzd10UiWmd3qh4
1PVtQeDmsUMNa7I7HwiOzvSeYXDR7FP9g5B/ysbDF/0+Uv0Q4FVu7cL31jbzjWGg
LAUQ85J1UtFMSFJg5tl8+pLxZGwkW66LlWun+fP3QcyHwwWgILsBpLko9VLawGZ0
rtmsCDhFxo2pVxWMxDQHF+mBASP6sppqacxPqXW7Ay33Ikgwxyz+KrxQ8AsOlFvV
lD33HnUjcuLvz1QdrN+bRWAd5EUnrO3jrKC8Z8dI1gmK1ETslH2L8GGfFD1FZldu
9bDb+SDL/PhGZvxixKRE94INB81yIsLJxvAlTLeqqlqBfH6v6MMT7H293tA5hJcr
oGaPj7rJBdmAnrecxChTJ/MmaZc1dDrjfeK/F2rzIssy8zi6VeiL08Jy2zozKk7Q
fvOaHsOEOpy+BVuW0fhX3krlFXOLvMVZ/HqMZQZZQ+QzA57j+XEK8uopba5IoKFw
Cye58ds25Kf/eF10csd2Pg3WH9ImyOHXFYzR40mo0VelcjBRJ+A89dymvH0XmpUc
8aOOpKvjk/zWWDiAN7i1XjORzPb5v6lsEavHZJpFr4lWRSBq92o+e/AJqAwJxdWb
5jScWX6I5RNikCMiHpZ5+WJR7pBcazodZ2Be12xRxCLTi5HPWyFbqmjjLPRCJS26
bX0lFfR9C5HpmiUuL5dbhbvWa8xaVgM9pR8IS97Pu351TwTS7Wgcugivl9OaqgKv
hP8+03moLbuCKNH73NWm+syOhn1foXeZkMd/IxbPmBKumIcc0RqKBeMn5fDesYeG
h8FVtzxd+RjBERifDumxDWcttWk/uKkZXUvShGiuX+eSgd5CvBOWixu0ifxee0IG
U7Nz+y4C0Mscv8hUtsEdhdMRhPY2rkphX5PI9B05uQbRZdxawIZ9HRbIK/4XGTx+
w13UPPq2PiJeP4p1+M7+Svc/5QfpvcvJg1cufpSI41mv6LgfYGpMimWkNJCXERwS
DjmvrplUGShZZKTHSeaqK9flWHgPc/IizbzCfAF2gDpW2cX0dQr1OtS04X7PifVy
IAzCUUty+qSC7EIo2LI2rN4lyvyiAiTPD+RfIaszNG+NUZVFrjZE1jyA7/z958+Q
ciis0vN7iRzykPrZXcMi+FZpnqVQqBPq3F0C7/AsDzVMe57GeAZvcrB0jP6kWFaN
BA21fcRPVwOS6+ot1fZgJXQAxCrgmV3GERyDZbRbGhi+gh83V4KGWw7RCHGymaCo
VSNYWdet3C4ED5HFdkat7KJvB0s5vJNJ3EMPwxItYb2bs0Lwgf35EKtmgQqqT2F7
4HkjLfrNKLIeoJFl4jNDUZDavmlLL2h0yTv/+zUw33Lb2+naM7vReRVtoOnj0+Yy
vpuexygOs8QoqD+m1H8a/6tIuF0MyuAIPyvJdBwXrn1Hf437H+FO39UnuyxdUCQL
AAJsuSNzCmsbaWvNWpZ5odFyR+thH9ZlXRQ36VD71b1VwL1kwOXh7OtZPjbNefk9
s2T9kRJ3gy5pBJQ61cWGWiNXdr3cnK2HATQX8GruYP83M203T9cbp4zhlj9iBWS0
BRKx8TY3ChwM+ja/dhupzV24akOn79Ymn96Tka1mO9xAU/MqaYV+Lir22MEA6SVt
MugKWqGbOb0w7/DTZs2mws2jW0RY9xllrlja1JGc72fbYB82d3IETGJ4kekUhGtl
pU4bcmW3w/g+ZrOm3lKUOHocnagccD0rmRrWhtXChuHY9Lqq2V909AeeEU8ew+gE
3XMJLsBYtuDAuTPR9iGRuYaIyx6l6M+1mP9YimKDUDphZGk11v2eHF2wMEHTfQ1d
W5vJT8O4vIMOpyB85d+hkdvjCu2afsXHx8Dah+tsivymg3qa+CnENOh8J6U4kKwr
fJWoNk2a48igv55GFpM3gvSztjaU7JYGNOj/sKjXhu/PATvniDawP32NpB6iQUzP
Ek7Fklbqd/CdDsSbdpERoVx/WirtVjJLnOT62j4e1HvFlIQHSNY2n5phOSvzvFkg
0dionAl5X5sgl2J3U+x43yOc8VKjjYYLhvkIYX7DFXPvZ1GNVx4LILRy41xzOj/N
BzB8nrWEseX4Ha1rQ4D8QGPOW9sk1kQ+oKlLxqH+Ks4WoSdAjFn05I9Q2DVlU1iq
KRu7qXIFPBwmIAeXN+a3PZgkWpy177F66E5blceIA9CK8VBs6RcMKKAN6Mwi9jcn
aampeDCZe+1O7ESx9Em53HmOUFxnh9Aeuk636bjMlB6MGUjABDVs0f5CPfZJcLOK
olR3uuxzb/vNkEYE2fwq57gbLs7FEbUxHwW6WW3UiZnkfuaCeOKjNWzsFpVXZRdE
okgX6DPbbwhBBn8Qtq3nJmrTCLlTaATnrdYnFT6gfgsbRDRy/lwioQ9dU1H8OvaI
lN8syUTtTvDUl8D/qX0Pwgibpyz7+ZN6yf+fMq08fTnUX5Ds+l9i83Y4c23wKbio
W8LJFO7CD4nyc/XZhGNbQAJ8G01zzRlLvI2taLKiVeSsJmOLfsHfX+vJNpnsL1Jd
YgzwcJ1Z6nyIMOK9ahb8+9qb8q5Dk5nvrNZ6C69a/WSzYfI9PuCKQx29g3GF/Hld
JSMbo1jZc7WuZMrJd8DGF/xhRxVciRQYpQ0wvrf5z/sAiWpGRR7APqmnYuVF4Xw7
oDux0GcRJTZgRMDFj0GN1SRG90WmoLeAAZqsJWQEhnQ/bRWmTWCxghdjstLCyDFh
fh3PLEfP7gkZUUyG7lYFfh7zqC05ZolS27PAPqVJCKTge5qWBAWRgRniowUno5O6
6RS+W7vNVogRDztyMyCjtdcVaJtco3NZ6csYQsWbkcZEwLhGy7gJuBDa5eeinD8T
YppSC7LCw4VqO4j/LZ5Jo+2UU54CEZ8/oZey1WVA8uXngheEHGRakvXBvkuiEQO2
BjRjUziVaStuFaMd17ySy5DtPV/UV209VuySU+fdc9s19scjLXxrBCjZRbSZqlDb
WDIOX5h5IetiPQ7fJTXNKGXBnqDBnJ7bCOJx9eCuFokpwYwPckTFp53G9xKAvInC
KhVDoN1Ib8tQ2ACsyG5XMEKe1XCK+JIKUE6SXTnIgqnIeoF/y0MM83vvrBqjpp5b
d8ItdUXcYlPlIcRsoS1CP8dc5fv+FBAH3Pc4AIMxqd1QJMJlHs7TjO9l2QPz1Jv0
/7BtKEiRmnh8YE1M6NU7CaOzsb0F4ag4asyhVtinUP0cugEe+yxqD1Om8ZjBEob9
8xf4zT/n4iySs/+XrgwqfKdKM1RMh6uAe3vxKVw0xO/M44opIexU5RpgEtO2x4DI
KyTVE0wC9JkvYPe6OIT4viNJtk8v1Fdhb0WyzANBHfhnT7eq6NRsbLYVmjVz3PAf
Jm7boJFfOfSXiVARaUuHvoxZUdEWM2D+mp/HHpUtqFcMjhg77FrRLchorrktlYov
0YWAAib9XQJK0OEH/hGJ8Io6TQPzLVWJxKNZLHLNHG9MriBiWep8IyLxKH4pQokL
GGE7BnPWRcx/ukdleFcvyKiWqJm93gI6TtG4YuK2I17X6taBInK0EbCqeJqHdOyh
vt86Hx7IfBDD6biBYV4txN4uW6yiNJ3qBQ3vjztTzo3QyC4QMinDB3Al/1dwrRCu
ZuK0YxhTbfOjx3u6SlU8otuxIPxyTRpVx/WmzIPK1irqOlhZHm4Qt1DGHc4sbP+R
D6sg8o1oNSGiZspgUUVKqpfSW+YTfDOAF4+uJQlfQelb4GietMyegLqrm5mdC0/1
ukZNniaqe1BtQvDL47NRLEFmANNsh5ST0lZeqUnT8ohmAJE9YH/qScSp2jdh4Ajd
vTXKo271RzXzOHDuQAXhPA5cK4UMSvpbnFi8rvvrBDwEn6HegDyS9tDqLshcmZhR
h3clwXIdrCbouxc+2QDYGJpRsxqy/oUolqJfJ0AwS4JYZMObmdgTyoda7vDAl86i
aJK9bJQpVM6KqEEQn/lmUJ63RA7fIjG7YCbuLlAN+dI5SRvk8FcYuQGy85Im8MMk
7QOtGJJeR18Syz+qptVOPN2gbE3TWIYGwMS3X6F06J/76OXgtzqex5EnjZnSY/D4
ETNGVz3iZPrE1D90Ki0QhSrpBhn3c0mWVR044+1nkVBAUGBmFn5fVEYtD3jelFd7
3VXD5Qh6OKKXvGE592N2e7eyw+b1ot4LRw2UfY8EoM0O439TXN7Kr1WvMPkxLJVV
lD45BZpTucgarFU+E08bodplpNASPDqlGHDjOuXj0n+pq2DjVid5rR/v604kO0HK
cbBP7Cv4dEncHa9gnfhM/AeglrQ2lLiCHVuLku2qWXUzQxPFVBl2cOx1G7XA0Juf
acLdb7ucRfogPHLKVhWKUMJSBEnSYYRdEmog9QuzXLqvgKLjortK5qU2NU3Y+KtF
A8AUarxv3KY6Lw6mAWW8PS0t+2c+upr41bwHNMVMD6mvOusSnIVnjQR8BWv/6lxF
/B0tr2Yr/wmHrhKblDBkj2sH2auuHsFJaevyc0K9LSDqUVx0E8DP2dKJJh8Pg86N
KcssUWsKonJ1MusjwUVKBKKeSLrfoNCFhHIOr2zHCNL92fuBNW8rDo9DTOBuKvDt
ngfTOtzqVZMHGhSHfCYYPoSWtd8zKWRz/qk8dld8q+WoN84UG8gDOeHFXRwi6cJL
LbkjiMLoyw7FPZ4TsP+hZLu7Xmzd5uP8hUs+SH660fEpzyk4NLUD95Mw1lY2vJfY
NEz/Kp/ZKRh0b5EhEuKyYUWm/LI7aEC43qGe1Wwsy2KpDsVzJj8DYFPu+smyvsL3
RKPlPUSwuPewj2DriHOMPm6DCuXp4htq8IYa3RfFKLw9SzOG4hxJxuURHRwXovX8
yZNUdOLcJ1/R30Wv08qsoU62H3WTEvkEaDYvXa8Tg48rM+xgqF1vLy0mL9Q4xU3T
dZH1qkAyTAglbCQG6X+K5L45bxOA2ungXx0+CVuzaCfLwvzqdvqLuSWb/ou61Hj5
XgfGPnqCur95fG0MboiQcY9pbTGxvdYpYurtshDFnLsn9rAQCf9MKC2HsVECDQ+K
cmk0xKz6+Mxu3EXbg5XPPQ60h/tFdAihBQKTTxVU9b3VAx9u0nYOszV0ySJg78Ws
PmGUlXzrDZ3tonah3PnmkpA41NSdVoUHV/MMucpLnwWbeiaUzBlyDbvYlE+2ni9k
IVmy20SgcLxVRwB52XJ2dqvo2m05JXgUahA3+qvgf+03/hzzbTN9g4xTjoq+tiJv
9BOZV2zxdafys5cOal+UuL6SMp+KtC2RSUFV7ww8kKoiVsTYuPcg1PlR0SQFgu4a
pLa7EV6tMhrJUDB3/drvN/+kO88LlheiI/t1OFDnEClW2kjaD16OEm0BhqiJHhHo
MhOWNmQ9lltnGFvSmMJrvAutjfu0SoI8Vg3UT4hyWyvz/uhspklVaTWeK9sc6ZGi
OTbaTd0kmcLZyWgq8sPUQxW36I+H+Ia8YhXJdD7hjfgTRYNrDD/cO9X7M2DKHpyf
8t82tQhOthL7+TV3SOLdkYfWOm2B65QXnDp44P/WFtOKU34D7vUsFIIhRHm9Zf+O
SR+HccgVJvrn8augRZqfNwOizkhsQkzCvBqeUoi+DJzDbfdrKV9IM9z2ewwt78Q6
K8PRHJXJbo/E/fMuykkLfTntoSIXGtQxjEXEMrKDtR4mjHBIc9JezFIPJvJq6x8V
MpthCiHUSW9dTwKYhYkoss7yyb7cPO0gHUjA1ZDZGUb8HZlrg2oeebVIyjnVIIIr
oSA8zO4aq+1Epbg5bRzmGmGLOAeSuQgsNZmyJyT39zTXXR2LwInFFMaeDPrJkoYP
v6shidfkZMtfm+YSsPUzdx0fAbj5UY8FR7yJJ9NJbYWQwAxIBHIYVkAup5VdZEmo
c62+0GPO/Pov62Y2oCWZGMaavqfHdiJIxjcUtRm/mBaAVftbIWfdqT+TW80fds3j
zOp+YjJCaC9eIxjY43R2oroRBuYvn+ryLGhy1swgYcfztLiPLIvfq9100pcxkvM5
FqS6Bm4GScaqdnbq7gDbPepZUT6i6Ranc/DnlGCB0SVoBZ31rM950ba/iTPz95KQ
ccwUx4m8KPQZPt5oQn8Az7V7HW5kJJBM4aXrEZz8cLlh/Uj6DuXcD9qkwqV9DerK
3Ii6DWEJrXInvXdfaVi00x8jj6Eh5tD7qNugSXdsNpHns7ERioTqaivMAuvgiKAx
Ai2DiqPaG8DfsU3tf2SJrMjNB99UlZCeBSisBwfZJfozC6c8+uftk/S7iIIlbN0y
xqXdR0dSiUlTZ8u6qeXXOX/WmfBn3Jv1KEJYKB1oH3cNUtGCl1Rsr0ZKwPuAYcGX
Zf8EPl28MCnI0Y4FWBurF4grNRGMaJaE62LaWzQm+iEGcjc6Pd9QsaNDb/YrUAKR
U9bSiozq92IUX6JMmFvu6eCso8tx9QAs3HYghYe6sr+SO9r4dWgDzW91TO69O3WD
U0Ny7K9Mg2dZjKgp7gTkUn0ckiMaZ8gparEGOecb/Xuof405jL+ill2pKHwSUTyz
muTUHyVNrdhYUMc2Hq9A6ERUCMqKsZi4pbnMBjvAhqh4F5I2KF3AvN+j72U+CQu7
Y/2StCM8JUl1hwSP9yRqzY8UaWxaxYRjZ3RtOc9QfIT1ccRfyjH8PraJdEg6F39K
x3JTEMxujNMO4fY4InEyBT5aWqXV4s0qv5x78r/DG6hFz685okZV6S1p/VU7rDBQ
J9Dk3NvkzGc3YZo5J3aIhlxWb1xErUdJH9ERuPtYaUKMZRcIOiNyaceAW1JU+FVj
YyiSI+exZKqiNVN4k9e3l285J+ezSUTTsp+DtA5g+PsBQRrixCJzQqe3oyyh4AIx
CKwvp8hkWeztz8SD4cWLgA+jQDxI0ps9OJuXkp++drDkSLWo6QRvpriDrv6iom4R
KL5UDNbDAzamnUNfC52GFJCc68HoH7+hxaYduLYnGvoATgXjl+OT51QJm457B47K
n23LkEOvhLnALX1hTk0OnGDj/RflshFQaWvjktok8hvu4cCec8sEIS9p01HwigGm
IklPxdxN+45fWI4eL4/YXjDgho8atuAk830cDlMk53YR7q7Quv63NpP1hrIpIzet
di0mVcjOmM8cQER9lk8C7/5osjvSo/gnzNDzyH6AD+UEOaL0pSqq8Ux1Ob2pLcqj
0zSwjjaoB+RnTcR/tBuay+0w9JetBgi1NYF7BExNrvV0qLs0G8IIsUWfG0NotJi4
gRv/GGVC0vDlKHcoDgZ2gJwIfaVBxjmy2gVbxmAmoABFAi+EB1w9AEzSDhaQC5ad
GkD5U+f3pSTfIl72oV1frqRgsD6k94UGqL+41qEJlhkwT7Jbwml6H3cg40enVBMi
D0TIoO+PlFZFwPKBAa62U8ZkP9EYdB6GCkMcTbJREdr/riLpV6tZPcZkXLkHREM+
GSeIQpa5rs67i37KYTBMs+HVIJUOo2Y1STv2/rMg/1bOsy3BTg1Tulj7A6PGyJBy
HGEdPjok/MZNO1QM1bwkfPyk9qr6l24N79TfaNs4x8orkv32KfsDD3NB5BAoSyOb
rSYbdIzRaRA79QhoPSVXjdC37vkYyhZ1y6zaTYylQCMeJ3IxUizRujhlfT7juwK3
No7Vl1F/2pOO+ZwVdmnkZ3PLll8As5UWLogslC0QYFHXpTlC06Y2X1Eae5xM5XoM
4f0cTYEMayzw5Bz/8qPfy9tFNRVV09BVNpX5pTwukaVXqjDXutSzYX249/17kmSk
SVLbuStdLam+Gtva2grkI4YXPfHwHEOpHqc1qhypBjsKCjZgcDX6gCNgH0y0D7gg
DVcN4SZAimXVG6i3ZeC7VX+bhz4vCeB12ckEw0PGJVyYmhFNi7z+SdIOYVLkr+SX
TXZBFPXaJ0oz90p9jQZ29WuLpzeSb87FqgcM7kiy0Xy5D42g4+IFzggremlHHtiU
SPeAAZUlhRID6yM4S/UxrPPODEzefTX9tX1OaOl1O7eogzhkC7E8qYjU7HQbyyAN
m5qJUbQzytIVztWYunEH53yYdO+ih7/7jI+B8HFRgDNhMc5vEc8OWaff6SdRsrdG
/fzSZPNLn13FjrRp4hgw8Byi3fipVpdHdBU7qd509sJt2ugS6QzdTfp10CDB5if1
ng4ttAQCIHONInDlyIzuZhsMpXwUqq7gSigRV7J7/sPwqgXdh3skYkjC6bk9Ld88
rSBsQRPvldjvsIlcicM6UUt+7hZf3X6220pve6GS8vSfZbgplWg0MB8nU9gWHxiT
JrG+kIT4u4Tm8eFR+baJkm3JUXuoy+ymZMgln0m2MJyjNYzkHjx8GP0LYlMBg01P
6NzH8Zcvrt/pxAhW6KXqZdh+jXUorn1khVodbWTrdll2pyp/AIUNDg6mzILDI7+G
mt++W9+MV6VTqlWuYhnXArlHqs7aiPzf7ebbDiNBlEj4Fg2jR9jOQlLAw+yTTY3T
UuG84QGzemfOYk1qNI4hiQ5sUUcR5A26TqxURJ2YCWBVtj6Zp5qWLVdyTV2QrkU8
Ab4iWPllFka8nrc0g9wYp6Vt5QPHJmgB37Me/KznbEemA5mL8DsyUJIdpSf1mp4w
GquRVz4PYWzObacoqknSXMfZbmgu/k80z5by0RsdrWjUkAbU9TCa7A2sa7D2790U
InFNji0R3Zlqty34xn6wZBoz9whc104Bll2yuaXne+4kU7tc2nFNaxkvZ6wtDNKY
N+HKQJ4+S2pnfMM1BhXAHhLyuWp84iJf1t4ATElPAGtOgmPbCuTxjps0yap9FLvE
TuDXsNQFaf3GpiQ6KIMf25Qmj2jmCyDwln4GFbOpORqy1YKRK5tJVZm/YDJZFe+g
+1y0cLWFaui/+bkga8Ia9qFDVI5bJQaxJodl5OGDkDF2Bktj5Efprg1XNk0W2suD
H5TAg9pxrBHTyUdMcVbTqZlX3guBNMw9kQpSRXQhw5Kka0QNgy0/oTIrmYSk9EPl
0Mbn+3MZ2LuRwQgZFevIVa9+zx6LUkNJ/fa6P+vVvszVZQ+lWMCY0wC1tgAiv6bd
dSuRCputbChJxV0FxmJ2V9RF5YeMKuxCZ23Mu5myEBR2L0HSzy23cWysGx8EtOi6
5XhIkF6m5sYPYnAE6TR5PSwrJj3nrgy7GVdVG0BWfTjyVTej3QYolYpHGOHcZZYQ
i+ooe1VU2LDnXLuwSASatwF54G5CMXkkvwbaLivggW2KBNsH9hx95PZC3AI62x56
4LUmueVynF2BuLviU6HAiA7KG2NsW7OkwXpsY+6vRWPIY4hTUxPJja1xUw9WXRqM
5xGyaxs3rqnyhjouAjnpxrFG763e2aIzeC7v2nbYdc9m6lkM01G6mF2B9DL2Fbzn
RQ7oFAvyk7IvmVynvh/UTtjPQUvI7BOAMsqv6dkerMvnbU/vrXgTwsQ1iyMHktRT
+XhpN4UQDshQjjF1HDx6zjkqGZ/FVJhEshQtghrE3+UcTez0vebH3nkxrmP6McS1
kbSVGSxTQiCOY3HTsqlqtWQjzlViHCSkfLm0l6oabjR+qy+G53qN1k5aGBWYcV9g
sHBm0z4AXLkizau4DIUMyVRHU2GWQUFhAAqgghsXKTAOyhAw4dP1yu7L5oOzxhkE
120orvInleJVNSDANyCaVDVOv/0aGnNYHOVOq89GWp4NX6zSqhuT9wMkmNdQYTeq
RHhWRb9CAmPDV7ZYCWUxzoZTJgBKbC4/A+NnKhKPEbFtm7WKw1cb4HMWInQkWRLn
6XWhoPxH0G/YU1atEbhTiJVVilsi5FyiJytIaLp0M/E9X0T+RW0EYl71NC6GdQBm
GtkKQIJRoqBhTkCcXnkF1I+D23QAL7QJLrF8lhOldyprfKymzLOzS1Qv9M7jlEO1
M4HAEQGAFlCGJ/Uk0a0q86plZHQeI8yixRfrT7/w74WTJ+r+vEQsN6vAyfFV7LK2
QtQn1SCd3icdcsCI9mXF5eYGotSTPydYnxhTRpj9eIoVdFaw122wsm2eQpx2wunk
yQhZL6tUrQEnZlim5Fj1yAkvc1xhinNhMtRU2UUZtxhgCfJZ2E+dUA698zCpy07X
sZJ9ktN/9EldIHwzlPRGMOs+51q3oDlG61dp58dQUnNJPg8TFa5o9ExFvjxbJpYD
1NIkssYPclWsi1xKuX+PEo+XKnlI4+u18e5vpMzLMtccKO0WOnNyOaK1XGuufXNu
nT5Au0VOrQU9yGNd2C095FnhcPHjmGc6A2XZ3zwdn0lmZmzr1qLhpXf9VP62CwxR
Js4+xK+1DxTGzulAVL0ThPa6YlW0E4xEbAwzh01u6hWWxEhL5THF+0E4VBXUQ0i7
zmD9I1rdh1nlIYssxdn4BPibAZbalffkTqaOQ4IV0ycWClgolGJ6EJWiaHsKWc3w
TWeGm0JtSApsB4BsFwCwicOoTY2aUrltkXluEoMv2yuI1mnI0ctduu9mei1g4BfK
s2tSOlYcJPSSLi59/L/NXr4SOZAiIeh0MGVFp/BwUyrruN+S++AK2D6GhTLbWW1F
AKRMTvnMzNcmtDj27gU+vbTu4vD3walEnh/B0X8THIDAEdIKhBht48Iih7IaNuvM
zWz4AbqcjgWZEvsdlqUIqpHDC3EXnM1hnGdbDqnAXXemSfGMdJJx9cXtVFWREKUB
2i82n6fjlEkg7rQaH8qFOWdfwBWsmwu1TW+DxSXSF70kBn2++OD1Fs7bxtJzZoOx
+8xXJ6E5s3juInuNt9bItdTWpMw36v/2d5CPLfLFv4Gx6G1dNwMaVrgK65Obh9N1
EFSQQgSIm/Sw7HQrOqOaiIxeCD6ZtL0cklUFfOoXRGJ8XPGbFoubx/lqIQjxwChW
lb/tSVcxqIHVlwOWIxVujOYJMg4imHeuMMIb/IrfSXTm3b2Aoez938MxvK7aKrHv
oHL+UQrZa0xjYoqwp96dHxHD6kgJdr0IawmVfg8kawZCUIqWZDAQLoWxFXD/d0qz
tIJ5EUarx7EvTD/prGzsRFwzoDqNpjfZT34a91DerjOH+1HF9ESXXUi0am7sXvbw
45mUYCIQr9qDXQI4y+6FfE9jHpRKIBFEeQNaXs5YMpwPI8XaFtHkf3M7cfLxyntr
8E33/I/Vt7J4tXeyKXd4aO5i97r0hjVDlF6O5K7OFKUQtdFP1rYqqcN4XdnZ+YLc
sDodXxzZeqWBFUBTJVi3H9f3hP1K47DPkiylAqJWyeAg19zUh723Cq8+isS6wr+U
9DPZ6gDjCn2LtLlhKUDra8eX6cu/NtjCxdGFUXvTVDCXYO8DKygEb8qdbh0MurWa
NR4SG2A7iIbSfNPcLa76++b+G7/Qx5xdy9FmpEAQe0jgHWoFnVKL9LOiisc0AP6z
2DDOTUjzL9yW5P3tG/1W7FXDsSB82KvvocrvMgWBUox+2hBe4xcfQPzqAItT2OTX
hfYKjPJURAB3/dVTT/LfBihCTk9paFEsW0FGh68fLkwKd+ADVLjWy0nuzLbXGnqg
gZbbglh0CEfkZNcsDBU1+HzEVLnef5zyQdmvs4psETuVf5eXjB8WHKzJ7S93tWO0
9GssmEQYm/G6SwG6BbXO//lgdmzfg4ThqwRv3SsJQaAdOhFyC4m5TWWk1fuW29LQ
hyiz0y9oW1hVoYvbl+5LL/DcKaUAXaOpw+okrzOGXQ172LbiIEpRh58N8jWflN9f
7uHUd51lTfUa8f3HOWgCmUengRMaoFOtUSK37DBcK0XGb1A20wK4GfEDCSbhw18Z
FKTGnXkRh9KtugQQza6uvEZpFQ2lwfs7NcILdJH6raQLD67/G3smojRZh88rT6ci
fOIOphmh7+6pkS5Q9i6V+yFHXafpVqWCNLtGF7XGKuK1QYSwTu3mBxob6PusXmk9
w1yjDZVT37mosFGp742QGeik0wqgWp3kiCNX87IT7tX1ZsDXPGzCRjFVohD/996y
rOS8L2Ym3QBGSJSTI4LyyH6U2itcWoSFUo1e/2i1IFjze69a0aFDOvJjlfE0+RpJ
Cl9iPoI/HbKUtEpwISHl/xMOKe2VInHluE1WELw3ZJn3m+KloEdMUrDArpNybiRh
nxPJGxF9wjmdW/nuOeYcCX889tog0iZ7nNKBghF/3T+8JfbpIhhKUrFnAlPCTb2D
6OXlVBE9xNoVwkwy/v+VaDFAuqSJ2iDlYNQ463WClYo7qmmnyvSDAx+5ZA10LyrD
tTfcXp9sk9ubAvlp5JxH5vbaLus/TSLvJpEhDuky/itX6oEKTvCnlFb06B6P8qIm
f9UaMup+oiBc4gNi9W092+6vGRy0g3Acv/SB9Fw6Zi1bZJfoJBU+7NYlTxCioMsy
z0IzOWtztfXTycq85stumggd62FRRH2fNrtTK4WbNX6XwpjShklPaxK7YXt46ZC6
dCHVvnH/IkP+fCx0AHAF3MarwoWLjYFyaCzIqW5nLk/ePluVecU8MnVzRZ8TxNCt
FdmGzKRd4A7eH60u2sGucdtaNn7ysTgXIY6gQv3DdgzKHSUhtjcBwJxUduO322x6
zDxMKdfKkSE+gSi5I9uayno+ksqtUyjtRn3thIDRixGqROqH+dsgTVpfFdJVU1BE
EfSQYLOBlHlSktBGMLsI3KHqIEV71VdOG9nAcuyc/uRh5SRhDYVO33PiMpG8yfmV
mvKUGX6Mi9q1XwMbY0p6xC5/u481ka8hSqZe+HRsxoZ+Ruenvy6GFXiIL5LY433G
4f2/nHW2S+37GFeKWW2wTBLarFuJFIQjZJ9nhr+RsW1cVPiPSw/GSdYFwshf9GaR
uWSV34VFr1IrdAZO4bZyN3DteA/drquRjHAUPyisR3ngMgsqZlaGYFwfVVHlrh7K
KqjjWnViT50mqBEhWolMCzkDFZPMCJJwNJupfAurFNAI8MD9pvkd4sX9IfL6+ZQn
46roe/9T+++U5e2YyNyf/GhbO7AGKrLfqyfYZic9MpUUGSoREQaXOhBiJyjx8h4L
AsjvU2o9cczQnMPsQadXLUyOR3w5JJDjL6vs5J/t87pLQaV3zMyrMoZ6osNiy5XS
bAInnKRa/yceqBd5tolPSmgZ1SqfGV/lITIGiVcIEvS3lF9uzguDuXSzR0ZclVLu
uTOf/f+sHq9pmtVBOCKhDCTRVdKVQJXJUoqT6YXJmeXR7rcxhQaKxdtySWr+e1kE
gXAQu8G39nU4qAFZEfIiMGknlZ+XkGk53XxdtXjpyGZnZD5OfbF95eXXfrlyyS9o
dHL/+3X8cOIEhKEgW76/79yiwzWTL8tk27kzDSS5eBod5M9r8zL2uZFBUiMIuI+A
h/yDVkmGCeOND8E1WoHw3XqxdBavmAsw3mLTlroNgaO8Ee7ju20dkcI7S0uB+jc6
e8HUEEcaoXwI6PDHfd6dUnQiX05xKudqi0vythPOyasz7+EIA86zicSW8uDlt/6C
aW26shLBN33GDvJRt3Oteg0xUAAME51TzyFZ3ZJNUofXZlHnoEovHteRc+uaOE0y
YSPAH0WhxYj66C4RJomOXE/LPkOBWrwiZrjqaJkE1ZBQPeCRYMBuISBzhWmQo5ox
OKDVbRNVul7ZLRt3MqjNLmGDP8/3BeUFVjJucDknAvvzRwSGTlzWwuimaqEp0XZr
TzLC4BsPuUktRCrTB+Dhxn10LrmhiSE5WJ2u7d7vS+pfYZNMv5LBrFtk0SGwIJKy
CQU1a1Jo7VkmUMNBvz17nAwv4u2thWlDmUxcfEj6pgbz81+E5Jo6f+Ei4Op+fg99
toPw3bvOsqtvV4TFqt8eajDna/uZfK3hKQN3nKHRmc8O2kDOAchmK0fUoQ3ivinD
POKCc+g6sxWvZpzHhLnkcc4fgDt3Y85WP1rLrVIfIO7M8JsG4HW68NdMuktrAaL7
vX3XX4lwqTz/x9U1TsX1gKc6F7De0JrQh90dbzn5p/tAL7N9MwEfLChJaXdf5yTX
wnTxnKzanVLzC3Kw59j7seUvGDHbmtz01/abd3IIY90AxCR6L90OoH8DXaOBIHa/
J/qq9oskYq4ENyf+leXFNjfuvwzSDXDOEIkSM2eV0bAB4R/MWeaKG81iXHaxertH
qWT3xqSTPmVQTQzVFlADj2I2YefrtmNpUv6hA+QuKkeaTWUldMTyGNX2g/63Qmcs
4YfF2F2HAMSwzq8GSsLFJLLN6i2EtbnAUheZWWHNbzzR6fHV7I/UxRhgC42bNhRl
qXAEzSkrdHqBT/gwBrG4+LOgVOywckOp2psbeBfsDFARgC2Pwibt3g4huiyvPfva
zoMnBBKXgQdDKGQYWXC4fQnrfPSCexYZajSjJ4sKd9EwhFmvalP8wfIouZUL7RLI
5OoWGIzhucaJPVBW2DMFOZifrYdnIq/n4UH88AljUDSVvz5u7MIYsHZ4DqWZc2dZ
63/5oac92wkCCFkzEz5FGAZk6ndJenAZHbPLe7XQp1Q2310xeYUazV5/09sdAPn5
VYBOmz7Mnr3veOKbHy9DcRZq88HMiaFNodsxAFOeA+puC4BQnwMbpq2fXu2Rc2/S
jJV0NH7nnq5jl/faZ+d/xcAUoh3vNBeBSGmfeK+FIj4N9pes5wkX8XfLfs3LcAh+
xCtRcH5ut6IaiLLRFCAlXxjRHqcyK5jl2vmJWH4jG/Zpmpjv9wiaKUtjzTBi/Hw5
3/T3GBXPJAucMb5pe9JVIc0EmeVwjCC3uVvYObJCTR1DBK9h30sdg157CVCRciRL
pCODCV/8MWD8iSX39qN2p27aHdeX0fngb8vyrJQa7ed+Q9DwN+obfMr2UDxSIrKW
boHfzWqspMhWdZjpQKYoMDaU2ksJGnc8RXZ+WTC8BK7KDfkaQvwsO5SPUio5BR90
PBO4h1lBKQqxaSm0cLCy9JYHwYPiI6x4sTYhYhnaLnKbLbkw2JWYzhh6AWh2F0wb
amWR7yuN5AyjwK5jCgBYaTmNZQHvue5AN2zXKCO0pIIk3q6UbUZ/NVHsN1OehhCJ
B9u+EjFbrA8WBDl9yYlZI+sAFyCTLuU8kM2YUj3uT1JgDzk2UwRDnXuJBP7efMQR
ZvOB9jMskKoYT5UxG8MiAjTiuk6CpJ+DPVX29Cj9C6+mOvU03IiMvXQI9wexI3Ta
0kZA6PrV3a2z6w7w/TB1mimbhoPWMT4BHoaC4AH4UAIHG4Ok82VMahGDsKGGe4kF
wAn1hnB/ttmGmtmoVSOXo21gDIH3JLG46w26ifBnz/Tt3Bi/THKhBEN37jDMlLtl
3ByEPKAF7vS2Yqg9sGbJkkmBCfTwy144TsuGKxMOPYnmZfhOxzdeZaVyHHVI0vpU
Q8c7D0uLwt+0agcO7I/lnzu0DJ/sD0cnCdbbGyKABYpfJ1vAX0RNbQqc+NQpaXNa
hzndJYoGkmMAU7infJLdhN0T+ZwYGXtW+BbL1k5SdbMg/Lo3Q8lo+xxtQ8OWbUwC
V20nGD6d+U0eVULgdC9qxrNu6+MayEgGdApc+5mWNGq3yOZi35PKKITeu/pSbkYT
BrsqRsvGn8ci2z0kiXjrq0wDlCjz+SUxZC2Gcwt1rkPrLTy44ENpBx0A6yFaTXo9
2EWlgLdEwbhevPYJRhn9BqOQxtXDhyzk2N0wRQ2eOraUDLa3MXjk8Y56GS1Ppalg
mCWE976Hz2EpfuCMbAiy5/1KjfwWE/1XvkcuGnkHOa5Y3ANABnHGtmnHAhmRlfvY
koIpIC9GILbghKjbL/PhbH9QAcHRlaqEvf1j4uTIG6g65tLVAwm0Uzd/Eoz8SWLV
2kNOMIA3lE9sYW6RbhUM0Ebx+EqGXAmgKoQRDKVqde0Nlib2y7dKL/zFVOlY7BNz
He8QbkBLf93eTftTtcXPv7yMpHnz1c8bzEZU052g4cxgKacDQNDYG4iXt7MhB/zt
fgB9BiMfg/4jp6MtEoKX8FcR4r8GrBsDjPmxhamrnDSys+FxwBRxkEclefQRgOWs
CSbqmgNaUzCZaHDJswi7a0sdP3E1yil5AvF/kva70H5+JXe0aP9FN4HkV6Tk6XHJ
WXEWW1yWsICmKO1/xQg8V6ysmWalH/StT6NKvKL6mZRKZM+jxCTXaDchcBv9pf6Y
ILqdKaO9mP3YwYDDsxwlirDJa2z0q+u1Otv3JIZPdURMDBsaUvUqO7vQp4AN5JIt
2xpD9JwqjQXuAk8TZq0CjQ1QcLtdlctAOeZp9y2YLcTe3t2jr7cBvcy9g0lBhm56
X6XjsFZFvlrlqvyHkw64tpse8KIRl7jf3R6RTU5mtBcVpxY5OX0iRDeTdukbn0/E
4FvoghYRqi7J6y/nfPJE/zuC9osGQ4xYGbr3cLqShDYWXdnjVWKl5Q5b6NLLW42Z
prqNrfgwzzO29HXx3EhRTxYNNKpbo+llt1AGRou5MZjxhAL9WUYgWP4loSN7CXGa
pDdo7yBYka/3LyRfUNdXEGV4CtqchbsFRhm2yxyZqU1LLEdX5lwLx8p5IQWT7MAN
us2lj08j8biAfl4WOGxWrBvvjXLneM3EUnsUo1itOWsn7ZbgnaRjFz4cYMn02gWy
tkhqydY+tAvhP/w2wddJDSMAT7xNR+s5AwKjvonBffS6EEWeoTiYdkpwDqJG/N9L
RME3ZTCcs8TP+/DxCUYnERn/639G89fy5lHDbdGUyf/5kDFQH8gO0w9+BYLeCi68
w+8E10ddzpqudOhXljjwV7Yds47pS873hYWcGOmGu40l28Ohh6twKSSbWQHmI7ox
cys/WMW0tunGXdlsc8xrYh1y6K1CmZNgtjc7lNwYiJZ+UP9ozPxDUW6XojffP4ZD
5AX04MCl1ADtWFe/tO7KqiXDbxZocuOxIauiPp1RDIwcyfAxh79zC/3MJ9uu0sCS
B9uZfwysLoSsC1RMFrb3Aq1QXUk/wJIbVdCgD/MP/QbkZT9fcs4lp38jSAeSMawF
FlWqOPUjnVKbe0l1Lc9KfxCvi4lw/at8FOBJw9hiQdL3a7UCQvcKlnbDfbnhhAJf
5p7rvlGeWjaexau7YafpTs/jRcSGS6UzLo0PrZUHnGpQKO+fXh/XZCtMh4dMaNhn
5nz30lkXoVEtVuolaApw9aSnTifjSNpe7eIqghg4JvohPN8YTflREUAh3DN2Dbwv
WLrvBDU43z1eqAyaNc2t/lt5jJRfSk3mINOX7XvyrUNQyMu8LzNovQHxW5q1zu8h
0IQNfBBaMwKtV0DJvcyxBH+ulICVwujetulu3EAAIQN4LvYgMsXob6771LRP02rY
hUvwLASrPauhwBr/8MlhCWWX9ndo+a2KrFIzwYh0tNSwLFNxvXLC+UTubdqiREIi
1ga2ID/z70Yk9FcR9+kfyD8NAECmQ0KJ05VSaSpGIPYMjs44Qzv3TbRmaTsjIRp5
A+WyFb+dfUwCgRl3zyQK/bPxCHSq7HY0Kmps2B2MibUzRpRUUfYXGGgqLW7UPzwa
HDtSxS3fjqYoopf130q9gllmo01uT4xyQkUfmPtQ85EInWSxZTWr0X/1GxZ3mZSK
X+L/FJG29AaHkZVr6LAD7Rfgx1d2stU5IjpWQenN/zYAcLuTGE+XGCSzKlURWDie
Spr8rAyJF9yAUaacIt9PTdSdJJy7RCNaIV7ttS3DX3WAy3QmqRtWzTnsNz5WarOf
pTPOtDVCvp9QThV3JfMG8CaoYZfl4gPWb7JLWWnwvRhqOOwiO9oDhtKVPdKIK3PU
JZVTS6ba62jA6n3zbk+QG9W+jx1kcKua/rXFfYcQNKLYS2FVti/HpUHwChUrIMtd
BJtI9RC9te/RLGltIFwrZZYelaoDMC/q78n0SJlGke77wmBMxPUVR2fGEwXRtvpL
MgMfgX9bjh1oPGZ1yqMpa6RNlvJblDnhMfjN5Q7UyMFBG+0t6tKJ92mteR2N07pn
cLv9fQIZFu9NEvsY6OdR4RKaMra3X/nkXNWagQp6ZzDvFsPGGhBBHy+IAXpdHzLw
EJjAajvxFqrPxywviE+Z8y9quQWalB2D3DcAkMSMEhLCItWUvnsSdidcxQwqYdEA
pO47cpG62zal7L0ZEUTHfm9kDJkUkoSvtjHD7cML824Q2BANZcfkZsUYFilZotq2
rke11UKFrk+8nPhFPExUVWTYFWq7juhHmTKIFJzX1w5HKhol59jtGgDuJ/1SkLay
oReOxs9eozHbrPHdzx686yjY3pzURwebaRIgUyO/XCZrv0bv+UhajwclpJ9anxIt
8bS3FZYyM0aAcNjmZMhS6o7vW5kees382o1N6Z5BH5gXYOUP9+nueM43MXjitTN9
HDGy/2e9+QwTrk+Jni1cHWAx2BfS9dWCAduJvX8cPzT8TjhN3f0jxGy4vBcQHrDT
ScOI0N++aTOfJKnCagpmfn7cv8h1ZGzWbmXrSn3ZzX8KqBCKj+0bUcVJI0rEV7a5
oWrgn29CK5ojcaSabm5LZi9CwfBBv+BkWUBtclYiGKx5OXbvpiz4enjoC3GzOk92
2QZzjkAW9AF3DjwRBsbrKIVGDw4guy1XMTOzix51hZXu7N9GmXcnMSB6GYVBXN/Q
JHdmeNBP6oGO2IhZIWiNzd7QXojKPLDhkg2MfshBB2kdMZuzgAl79nY/Y4fP1Rmd
8CL0nBPdcUW5BulZwf+ltbZF8OJ59dH62/JXXnYVf/KOFMf3FarT4LCrvmNJ5XiV
KVfI/kU3NUFw6KKDofgE5laWRoB3ZitziLpUCIafL0SqF488ADvJxrT95ZihOxH3
u8wExc2L0PmhpkzunPSKb5I6Ua/cwETgTO/TykiAn6mnkv3/PrEh3C2NK23CHJnf
631kyfTDv6SDJ1t0jJ+zIqM7sehn4fv1RqE1dvMzWrV0XZBr3ifkDSfLykNV0Bs3
PswbcuAZSlAmF8dSvGpI82G4szvVjfJBlKWAi/XyHeE1OWTfVy34ZV91AbfwI8Hn
ozsRUcogALSaABBYjpr6Djk6b8+5YBHzUPpINKrsDSXVZx+oVUIdqBxjZ6NBjFBw
fR9dWvu6pqkDwqCPCMALjbgE1It883edYC/R+XRtnjCHaqVXHoEWXvzsQroimJcQ
qVdjUQ8OE1W7cEypSwddJoy6jEmPNmeLMZAX2yNFF6YwheIBWXRUM60z6Rx+pv1M
ushXXt+i4p8u6E/om3rtQyTMfg8B12QnaEwnoqnv7jBpkwU+xGBKY0d8Pn5yTqFM
KJezCJQCBcWpAUIrYxEKwgE8eAD3eHHBOGyTAEn/WRh7ptj38ynNVGeT0zNs/JN7
J5Xc5FA/POG354f/Fy8zJPzUs+NhC9RxdOhlQPuWO3l7pQE9ZIBz7uQrGgCOMvZL
AAqPnEhPEIwZeBUGSMunBu7Ao1Pu+hd+QvSLzGapgIjjh9pp0zJq6emiA1g7QDLr
siztoz23+J3epCWewmOk57dqa5Zm1GaPUv8rQV1DE22r5PNpWM6PQNKCsQg50eto
hvnvDxSy0m6uiOE1J5DoTqdi+89cNQKndhC6R/qlneH1sALLPsjyZP3pQtFKQtxZ
8jura17VHTqJ+qji/kTtfCWjuZcuKoeCzldvI1qzvNezvPx14pA+Hl8Bu57HeGrw
sX7Rf9SfjCuli9C3rjQd8dyjELW/J4bVoUP874bhaLYred/6WAt/4aAaRu7r16ui
Yuh2slLgHEOe7RXWpMblMv9AfDUAEoW9sIgnh/enIr2GDf0WQ7LGQD5X2hovU2tP
2MX0MKd8qLEo1+zFWR3fBMS2NMKxNBN1xHUvKFGq9zW5F/JxIRq8KVURVzW9+oYv
4CrVb88RmfuK6q0WjZdCSfSOE5Cxcty1hyWAExOHWjaFs9AgRGoMrj/7v1XzOhob
CKe8XDFeHtiWbhrEjRAd/fv1MXlSrLc79VgkRb/7XzbGQetJGNC9tY58/nAmHoJJ
RdOo7uA5hfspndLegTHcdMcASoR6t8u7Go26f0Q9fYP21Owy8uQmUwrnZaN9OE8+
1kCW+VOqLhLoinbDR+aWbq0JwbTIwjP/F9Iw9dIAViW0qS/c++joZ2BRgVV2tl6a
LoLY/MO6XbFGElxXQStE5G1qrB3GOYDgCmQdfZvRJ3G01iaP8dmrQgFouABnOpTU
cz+nVeJsKdr9kNhoBT4oOPl8FE0IiSSdGMvFb/5BpNl0u2lNQRFBQ6rJIf/iJIB5
4mhOPjOtqsY0FHQZemn3p3zfpB8hPm8x1UU5+z5MZsx+1JYlQMxmcuu3Qg41j75t
s3fX0uaKLfP90ZpLQSbwSu3tL5c/89puClM37CPPbxArM5Gl1sFNy2uLBPCqW8bR
k6vOo7x8cz3BGdXyc4ik92cSPC8kNQdLghgOvCqkfQjtnCJS47jPZYhFpbTxDrFh
ZecaQbzg+zmo3kLlo+DFu0+h8+fCcfO3Y6ZJKdIy9w0P9nnLk2CgxHtksDynMxgx
r5TJsMh47qXTcbpXM7psyRNzGOOZ2sRSkNXY3J6RJfrNifTp8+yRSAOwKi/TH1/K
0izeCe3pZIia4HYh9fHiVFV/AQ4wDd3HEb+TOZk6nc7EKFvTbECUr4vTtvtlO7ir
FY+5FYFPbAqt/6Us6MDFErYL08ILaHdTO9+XFbuwnHUKSwVZ5rFIW1AE1UsQ7cvT
tWG0Ok8bfb/T3BFpU2tp1/qhLlTB9aXociIXtkynEuKPsMjORAVeujbEXX70skKv
No5DuC/Lna+28osN5ugq/e80ppqH8TzzHO1p0gUCCz4kRarKHMQh2n/YZ7e6tLKb
wcwHaBmWwI0OmTvv2XXhu8fMIs9vSQR/1lcpmwQLUeVTLZLqwBwEEiOoG94yISOB
dY+IN/l1BLLVXGxpcuE+H6Kg6EgX2mO5tjh5IQKrge4Jp9JeVHR/9KOaB4x6YI4Q
cWAOj6lmx277W0YWDqSaE78ms4ZrErSr6m+kTRnsWJBzS3dUbwvUgRBtz6TAxlga
h4yU9rFztu0Auz4Qt++c2kYEruHQWp64aoE+D3jTHnwtnakRU8IwNJJWSnYPdQgY
0OX1sIo21HYZhtlVILcc610bqV/vSru/Wl0R1szrSpDg9/4rxCShZXp9Kyo1s52N
qm9XeXeNLQ53P9+Ey0dJJj8mVCRwsCmLko9kJ2Pg8yvoIi0NCl5dZGTJODb/1NLm
Vqdbff6Bzo1RqMlnMAxMuoc0ZZNSP/lTAaVi18OIuUzuxf3hpQ+NzJZbOvmv+bRc
tIKG0WvFmwi4Wm9MHgGb1QFhAvwhJZF+cRNSaHcJuEG3LK8eNJBk7duiKjYfwWF7
S+hGc7MKNmisjgSMbqX1MupP4zWaC9/UPLybvNBZzVysUlMmiz481682dXCcHwxC
N706s4esI0Zs6chtlzPcP98FbYre0YmJlHQMwSKtDxw0q9jjY6RxBot2wo1ffFR3
fbtf0jwwzOtv1XeNUf/Pqy0VyRQmcXM+W1Au0lDI5Kf4aYzqyQHkF7LqjO3TQd3z
olJW0/YbnwG1BYNmqSc3mJnPSTTN0ocC5Rpi+KdC1DBJIEWlKi0i0koZzVcL63FU
ObaO/JAZWW89atSjZ2GF/rB3MgexZ6plDctCOJZue/OMGtleNegMaJAK0rsFQ3/Y
C5e85LK1/04VADbFH4vpHZQrpLI5Mj52xLtYOHtQ66OnI3HxxUgtitzT71no7For
2Jy6YJkvjb+D4MkQ1c1QptCk25B246zh9K/N1tosA0Z7DdEddfBXkMaM9VR/cZMM
qYToo+BZ/QBBAgMLgX9OJ/Ktopt6e2T0vtODvboyFcJoUpMFV8KYh7RHofi5TD25
1el6hKNpMlB8haUkr+3CXJV1hkrEKlqBIN07OhFew6qmz3LoA1RxWm3cJ5thhNEg
jYPb3q7MG+SknyEHSVoADhBjqPhAZr4ZI7PTceSYPDCJNMj52jowqg+L0sT2LMsq
Czz3YDl0hvZvlr8Ck2LSHrIraK28nrYXJ/JFLGjz0+ptf470Rzd5p7asjQC8UpHI
mQPS3WhE5GKrIBUALF6K4bhxQowszY07wEAThZQRELyLnqUmBIj7x4wFX8v/HFPp
Wumdg1Ry1vSjfM4FpVINGUtjV30RWUaxS3LxTiyKmSushlt+XgKpqujOEcU1AgYB
drMGw263yYpWHP7ROqi6cNBm8knjcF43uFMZ2MvWgWWlfSbMMQ+fzHmZa6sTND7x
3nusBaRRckNpGBVEI+uvqrqjLIN21MW2yb9wi3MgQa8E0px3ezUoX3DRW9V63t7L
S6V4R6V2IVOsyMqeKnfbPrVCy/IuLfkVdrIx2hFD+swwlwrLn/GX6wmoL1gT0C98
JITD9tMftGpWkI3KhI9kEpeB0fmZpycA3p4JkWTQDxowdyMfgyhZIwBPGbQiPraK
x3Y3CRp1RbGg1fXr8ny3kSmd5jHTOeI/+Ao6yvTuQrrU7Yqo9yG5qv5PwTTfDO4X
s2sepW2OlBmrX6LM4fX+OXtExFgbeKM6iuC5UoS+OdeRJOhd2ZpvYmVQsXZHKje7
ZSf+GYe+exlwegFos/qowMZj8kgPd+xDGeeHrwf96ZEDOHsTY7ePlyXKehtBIUF3
DfSjvpPeSMvXwRIlRbwy0sd/ujHCyNQfvmWwtvbSWGa5iJ13uWySFxf8btZfWfiB
r/q+tuApajmmATrUViCiKzI+uxYWEZqoCPKXWZDIThonJX/g9zjEBZQNrfNFockb
8de55GOJvKJMX64H7YZKYOin2QZ43gGf2zuCyLsWogcCNUq9yOLw5Y11zY2uS1s6
daGH7kGkKmQcn2E/momShlJVtAvAeKj+IAdC1m5ShFoBvW0sMSXDo+1nZc9+dOoa
CRLOB58L7cIGWpteEKFU1xCf/Q5/hd2DFKaDFzJcvOBCDCC79lVYfk4eFPFUmOQa
pO+Plc++kcGSpAPFGSvV13Ha4tw+oy4NA1lHDb3+o48UrAQzbbPcF+QZox0VO2y5
MW8V2IdgrKFl/zwPsbOi/xG/itcUEXQUiANt0N5VBd440c6+usN7zjV0pP5vzKbx
IW/DKR6pVL4Th9pjgijWoCiZTRF2BKa84USRFosNNJ2Ch0At53cuy+C6zRBlx89t
qLaxu4xdGNC60kAHZeCHPvjWOAzcXM946xHtVFQYewDL8BMQMMJ4/9Y32hZk/BgV
ztSRcsJb1kIpJ/GGna/KoqC0xYaNSOE4CQZ9BhpH5JJzqWGFJsm/KokoArfiCC/m
xqHzvYGyx+UNL9RN1GtKb8du9d8+doRKc5yTs3v4PycescnC0jyFKT9zn08SbLF2
byGI4iA3PAPWRauiNmGPtfE3tF9Ahj8tQsHWPD18yDyN+WnGPdn7lMhaEyPnmmrp
sNZo4ZD3Xlz3sWhE6P9ScKR+zt7Vod7TGNRe3nU+5YZokbYx2J3HG4iT2ebhmsX6
fW6aEfaAaoLae8iUtBpob4r2BRAzDJFdkVJGNj27I+C99Qof2DQVMG+YAD/6Imhv
Qm6OSceCXhE2cA8dALLztdn8Cos6+2AnvJZkPD/3qUjCqGsuOcIO95O+DJwCGNpz
YeDcZXdkTmsHj2L7w/1XhfWOUKkBd3fiKh4/uEltjgmVqGrjvuHTHniYmjHUjLZN
oVEs4OELcbzkjDsgs0U5EfnBkadkNSZnwJckoOuajYOigz+GgLD4X1/HMFsDTQ1Q
oX4nmLT34MgpuUnGFUilpoya5WmzYHDZmxtispeBDq3TodRPRSJoP8qt9AeFhuut
Z6mXHIPS0UYNi2Nc4XO44Y3slKxj/9OnSggCOPqMYAYMZnS5V8sFjBsZiaxOYloZ
jTHDw5uokJqkSLONGNqOjFjmWWGx5RoCjeL8Ch7Z0T7OKICPFmLNRgnW3qoQ0/rE
kEJj1Ps4YiWnWEtrkZsDk3DytZ8BPhwEkBlvb4GTOkXg/bYDeWdFUM+wN8EdATg6
qNVYvfr/U6XWJTrXTh0cAKNd3JHO1z0vwXI1C4kJSccR2dbDHdUgfCnkdogHqe0+
TMvozAX0zLy/50i6MwmETllTPHkd/UkhkBBmlfR/MyfLZ6FtOaZlD8PQ1uo2Qnwl
Y/m0ZR+uufbjatUfpyzdu649yq0ld1qkdOFN8Gt0TfU7FqwTjoDrsNaciSBuA4Gy
R1CUcvFVQbNbQsqjVN5vijguaLhQ+ZOTXylCrCb2NyCZhsXkbzdpov+TRkmXS8yG
zM2lcQaYjdmeKuWkV/XGA2/iV8F1o0Uxn3lBkovtfDEjfOYPuCWQPJESlvllTdWw
0XpBCJS4coUgZpgWRc7Z04BZBcEejk24bzk/58Sk1BD3QNLNDFYeyvc+mrcELLxe
tAGwBAMIYdSyPjYlBgOT7wJfL67Fe2/BMSvLftIqIytHKmEyp3Ynvw0IR6pLoBAs
/vERr5p5/bRzTYDeGKy4sO+67zUre30G8Ayl7E81zzx9BcfjvjJ6PFLPlUolTWGq
zaOTTMo6FCFydiVMrfbOL5EH5Uwahs5cB7roMVOPbTr3fHhrhP6e06nz/6x+mDml
ZBAk67dMtlx2GEvnRCRE+Y/BjMbzNkx53dJd9FpO5ZcXMmGvk5mjH6e+Ti1++44l
K824ipuOvW6ACvwbs4tD6YXozyTVV14Vn4TUuLQnncGelpNTtKuaemnxXSv21lco
un+T7phLaVG4b3s/ppi7e9uG7CcujlV95MKJi+PD7mde2VBEEKbI+Z9SXPFYiriz
YMfuOsIKE9eSIkdPBcMJDwVmRpqp3OVOW7f7VqLKmXI80rIqTgOcSH9KMxsXCfy8
aL3U/lY8cxW6j2kMcphk4jN7XNgw56py2qPVSpCKgiIzSXdm66Pi/f+7CBXr28ZS
jzwSZxyEKm8QmMPalkuyBWzL70GXWteHhOmrGvC2cGDX574mJvvfgVGtgqwSJmOT
tMWnGtBVk7VfR6TdY40GuIYCISe3pVb011Q37Cd496sF+hUTnTt/cyDaXnx0+mQJ
+uPxjxIw2DSYCrulNq/092MObvvZ5CC5nYM79CEJkMN+A4xLNodHoNNUCvYqxeJo
GBNtZAD0tFSSnQX64nb8vxPUclplgWhB5JgC9nBd6mF0fNLbjy9t4QRzkYxLBKAz
dENjcXniR6NS8MbNPttMgzwzX14YvFDeoZG4OGogeeiXH8E6GA6tVl1pH1Xpai0H
R09p6+cK6OrmLgpMkYiHYSU+8v3V+HcDmm3DqU87TdStG26SyvaA4EzLmzrTTunr
IOgy+P/x3AR3hq1wWp8s0sBal2h2FWPh/DrY8uTnatIpZmcWmcVpp6Plfl3WiV4f
bp+ZX619wCgteDb2LlZDLTUCL2nnCJ3SXgFWkn0bpG07j6M3urzDEjUFfJ6OJL/+
HiTwGqWDAne8v6cWFoWODkpunIyUyK8Mg43TYmzuzfoLBb9xAPbVgubvZfCr9bsX
vLREkW7lpsVC3TMWEs2gn2QECB+kFVqe4NKaxKMGxlnZFvmIV5AaGC5o4uMqLIVs
F266aTCujqupE5E8h8iHVBNcQvmcZeX5/E8TeK+uj+e10zUVuXGkDYDNy5auzd8e
9yfUwzpYCdpQCnrgGRL/EMmuIx+7xWDdjFh/eZB9BwjQyou2lrdKH0ffO21BKY/S
DDJLx4+8a2EAyRDkelZrWHEQKiAUUgYuH8o8I8z9d+AXREIfWe07enjPd1dNszzd
Vcy3KB2Xh6l2v0xC8cDYCd2TiB3MCpEwggqO3OKncZSBUKz6scXcTZqGneWzTenC
h0onQgEvTlKRoZtKn2W5nC20RsCNSpTzgi2M0QBO067H2Ao2OrF6kVBolx+1vN1/
8fGGGJ1q8TEAPsYHBj3/zmRJQCJc0jmbPiXEKg6F6OKGbq0e3YtxZ/vDoc7uhwjj
62G/cjLXtfFQuAoVxnFjjfO3N6vnl+zOAxHdau13DLrXw4S0mb57G7UcUIJL8Vul
SJV/lSzUMlPwK/lnzgagx1QH1idfzd7qHxwokEwhnMrKuHAamHBvisI8yLhQJXT9
prW/O/q9rkEDUb86eyaPIJRbrZEGaF/+UBv2kp75mE+vuPNsnm64uYL413ZYepxU
bwlbgaHf7r/3Rwgr7gxHZUYIbWHSHuAd2X6vOiXLZbxQU2JK0dCXPe0ZhlFZBc6/
6KGlZ8p2imF4762dhJ/yml6XtkwVyAGYzwxLawqqFUXPatKoOHZLzKVEz4BwBmQS
8H4fPy/xM5W3SfpDaaYfY8mXtbCJs0CHHbXe/5M1rFmSx9dpTl9kEycmbxTe+5S4
19rBLHcgo8dph7W4hn64i/5fOl41na80hKMaMDAOu+4f8JBnjm2SrPXm4cFNyAeJ
yF+goXI66kxZzOgc/WpEO/UlzerUv4qXrpY+1JpRJvjLYx7dZhnOffoCO2KJEESb
4cHTRg71pxCzWchW1F59w/uodzzsoJKgZOimdYo+V8dQmecPPk5sg/3qLqAG6twW
8xf43Ilvj7097i+6Aoiud1zHEhmdBMA6hkszOPrd/6NLpadOgB03MWW91pUphkrg
naBau5Sb7Mt8obkcYW0an9K6vjWPqOgGt2JUHzT6cgwFnTc0exm+QgMd804hNLzE
6eV9yCthQr86HpEeYdHc/k4FnFmmeShbKDjdT/m8DW4k5TZdJdvx1wDSxKX+0LCw
7W7f6Auq5o3msvD3nke9VCmlwZO3CxjTGFFBHpPbRUO9sABkQXCls9a/fnskeSaK
dqWc26Ewv/2m/jJeAaH6pqhNx9dVOHxFCX19194ShEpodqQIlXpURaL2+XvkpRe0
BXiedkGPICpeFU4PwGZWa+07/0S10hVUOGOVt0/s0oZdmDYdpZRm1vxvdGQmA82R
+vAIfXGbhjRn5PEPVELF1HMMkrsLb10PDOP0Nk3O1AZ8Aka6wKKn2yGnWdMtCqkO
9sxMLLTlVugTa5njgdyw1MAPosmskWDycgm+zVws+Tp9x5eSOR0RwVtVC4pKiI9S
ziLfLkzEn7vmcm+3ZOoGIZfFpD2rcIovQl+26DERaXNdQFl0NyIosAPPNN8NEeNW
6MqmMKYj7uM8ADGEl95ikS+WMcj2QU3flwomOd1iM3e+pY4uiNz4be21vMV1Jfwf
wFHIrqYGBZfUYeeV0mNGuVNJ62FNb9VeW8aQQN2JH/LE2DVn1/9NrUBDSrckqogZ
MeGbnxLJyzphJVMrqvbyp8Mzwl+P2wHLN4fs3GKrIhXJgdoCRJXNgK3IPfaw4mch
gzwclyAhV6coHhihr522/DtyilJX6/1LK88VdC/mqpHUKh3WSEGoqDhGz5dsRUEq
HqIV2Mg+m3jcPGC497jCqgVW83sLes0m7mS/ax4k/FTFM77iQygZzx/BHn8aHQ5Y
nceokCiXe25nOcOrUZAGnckphYJsDE//jcj9jD8tJINziEaYqikAzLprOAzK2Z0V
tgd4uETLi5xgOedxyxFYMzv2iBPixrk/7f2VJsrXWFfWbTEUpmqb0fjyNzZF5iuF
yqDvBnCrqf5mP02HjbxTAulmiuvZaM4NuRe3Lj+8pRXZUBPLKOAE/CDf0rCJMemP
3Lw+gUAw3/rq3Ft0A0BX5z8m93+3xwKSvMm0Nk81kdzfuKKVjrMNQWOi10WvjD1m
JK1pVMMaEfND2DnzGgcdDK5SRrtmREhBFUiwxtW3zk4DxJ8lJYhezX4eJZZM/ZJc
vowIvYmtVpjV4BuQzR1TreiW6BWvQsbdlFScpgc+/S+wjST0p9/jb7h7TI26KHaJ
F0FLKo0Et+0RbcnN19izxmd/CGTTDhdtvc2BS9R4xrkoAZygQONI/YDyQZoGiLTa
m1HuT5lkO5wWI2O/smaB3AK8iY3ffRM5AS7P3PnOuDFwYX/kPIajFQBPIH/1GWHf
/KPbhXT3G7Hql/xIoUuHZVfwKalIQy+4V4llocvv4pYDfWwMYyUd43kUcTzqRj3u
MDHUdbcSIM3Yk9uicLFRPFDoXTxEICHbNM3XQmbE52NTdwVFMnyMvYzKa+iOB7jI
YZg7M6gVNlhcVaWKs2wtleKrpAGdrtqjCYRPnCJ7aKzEhcWt1uLb1egk45fs6gO3
nLh0hF2GOGGjrJqS4PXCGApwo1/6tcVDEyB5c5wIVGLQ72/97mafMIYRHHClOeE1
Vlr3RuiqF5z/y7L8ROKQZBkZKbwDtH7s8oYqmoYALz0HLgVMf7D5TQjkFA0XEbp8
i06+Fzw+ZjNr/Q+W3R4+AmNBcbhpUeVlctDG5kf4y29e5AAvbR/YlVWZ58nYlAc6
y4pVddBU5ygxwlgOioD5+wqOKLsBYSMdycsiq1Vqm6pa5sM/QrJBj52W5bH0sqOX
onJCb0h9OP12GSjiyJr+My/j1nihp0V6SUzeMcqMH5kC9P1THrA+cXvZMYQgP5Gp
JUXabnrN52og0APKq/nfVhrMDLw9OUx+rDZDd8Yx7IgJsCo3OBEd5h/zQEJdCBB8
Z7oZujempJDFnRnB/8zVXelEoXwGrlTXowA6Lg8REahX/wVi6r770vrsDaCOY8LW
em1kUN4nUQJsSpcen7LBgOivQEOgNA/Vgz12ZN2IWpDFrp02xOt7fbtqeqK2q63s
4ZRSIh6zPifrqJkWs4pOCuwROCc2biN1+gBrsdNqMX1hwC3RMND7bQfYzW2id1MR
QWs/gmRcg99/habN6XZS3GAEJccDauAeUxWdurk1u1S+SsHaZf4nvmjHLnhIVKmW
kn8GZiMVuLQf39YdQ0zrvAUs/nKCHIkcWOlOanEZPwBDc22iqe4sMVCtOdQLm2+h
660eTfK8WkF0ngVe5swzRAt3iqjRbjDBDZ/EiGJOyOEnDN0QPgnngvAbc3v4mbGd
u9Ia7ykb51c9sehW9LmCXWS+XfOAaa26RuEQfPzmxxVU+PD9ibkY1wTOqX1XJDaQ
aK5hBzeORWWoIApatGWdvq883oDMnAZ3L65DSEy1+Ky6eKYExHljPSJ3VvabnmAZ
AjmMYJv/yA54mZZIB1DxALd3FhqDg9fSKYhYa3cql3Y9pQ55rTFqUL3lLCsrs8BQ
CaeRGDklNG9lDwYb17cLTX5Nw2TbWs5xXFifv394Nuq/HRyWCFlNU9wUwqvqxUFC
G9o8s34hWh4lr77j70pY3xF3QvuPeLImy4H1jKuWV8lEavPWe97poy31QjUndKSV
c+fErr8YUg4X76i1TqcT86IUNwmb5cdz/YoYTaeUU/aeDUTPIzesgGp1WctvARQQ
ec0BjnaJszwddOGoiIXiX0R5/cL0a81h63v/xiwCH9UG/Ax/RtEaeehJfnLsVWm5
cHzbOAMzynOQM9aHEo0WjWxyF3hyPubogbosAeDlrBFKwj5KA43DI4aiaja2a6Hz
2U7HE8DnaF/38uQueQ8DfnEZ8h4yQfTgncBqLqfwVl54eXhRV0BUpW061E84zhE/
1wwIegtzFg//SLPg48ZLQeHXe4hasO7wvEOHk3/05aDohV9wBXtpre2GK93TUd/a
9jmwq6dteEwYg6yny3CkuW9XPfujig2YlrluES7sn6Gokye6N5KD4IEvPlA5vpYE
fyE+5VzII8V7VAOuFHaHyMenz3IuNrz6uFr4FNKl4KhbsD/bgX1NHOXaRugMYDY7
T0h1cIfiS08jFO32Ww8cdmqmFW7/WSR9sG+WQprw35YlkIZaX4EwepmVYkGb0i0u
R0XXoTz4YNN5MDMXNX+uY25Z/gd27TKrbfEqSYdpqRRMqOh4rlDLzBQu1HcmNGWv
yXTqzkt3Ccz+xl5LrFJg50rg7OQnDhEBsDC62JQtw+q30q5GG4NUeuO81kqt4bpX
c8VfSkkYTvUVhp0QrzTykL/53Nz2Dw2qVS0PDsxdmU2685/hLfcSBWHZqlSUWQ61
lpvJJlxwlv+snhjRQADEbOwB2RrrgfB6M/AIXxQLLAI9cL3bCMSuDj4Ifsb9A3eL
octQaRZ79XUBG2ZYwEuwuDeQHgkypZyBdZunTAgDlTpEa1c5dHlCQbKxSXjKoTMF
svXRi0sdEbaxSIuNiBfgQnQCJrJGZmod7FKWycNI++zmClSN2bAdvo6PElNVDS/w
CZjlKNofV3NjWAF3zsoo2iCP7hbKPApAYMxU3FTWUcSDXETbea0U6WsrOki8BT+R
Wrm59FGi3wBIAkWqi2DpJo4GZPhdJR+9vTCoHuHjULaAUgGGbbeD329hJ6dchm67
g4ci4Pq06Gl/iHBJn8gbUj3sNztUjVqHmEHTRQtVBCc5n9ec9G4K43HzvqLbvJXX
HFsoDRvYP0Z4BEppP0bl1+c3LHSFxxszyOI54HylC+Kq1pN58NaXMsIRbIokZtw0
tG4tY7dTHjL6Q1BHhGy3mnMobxZ/xL4XBVMXevkFeyf55NrqZljcvVYVgQd+wuF9
wJdJ99rnjixoajzycvRIz2onRigNlhHI0Rgo6ai0lElVSaoq48Z54UqGZJR/oObj
EiHb37vdMcPkOYtyV9VCIjVIVFOBQrR6PJzBtZsKnkirADM8h7xqQaZTAMJsKfgk
auSNsVb4aGe2B+tdqOXeOAc23e5nSHh1DpBcMulyDyh7eqABIkMu55uI/NwEPKU0
+IGs1WclmI+9c+NC8nmdCxNmlLSLlhIKi+lIBcdjfsa6648HfMiTLp0UeEDsBDcB
OQ8e0BLH4XnEHe6e0S6uv1aXWd/4QAFM/idmjmbGBJ+crry4nMXBRDD6Nk+WOZms
cq1lO3KZDwzjv8RZSxn0JZaXqpNgXQd2/bptznTxjeIoIpG5BUVVNM9ts/lfgvBg
p0ubc24YAeJWPVXGgxnVSJZggKPr97P0tNt2iFydAACTTVRVFoO30+sQ7Kdg9pUu
6A1ge35jkWwsF+J6/oCSclmxsM9vHrr2dAYZDlKuohwitQg/pSTT71VFbV7bCFM/
9Zf13OsJnnr2A/LNDxwVHeJxBNmDEuHS3tORkNnqDrV4CrUwnAWqDp3iV+mSGPxL
vxDdJK6HaHF+qzTTliLTkV9EOV3rrigS6ZIxJ/4doZTS7BduT//Ob6I01reYPLVY
Ut9j2/kpXqywQXXWigO5t8t38Qv2/CCsNi3vjwOxge4EPvSXxwAEsJG7eg8u2SHi
QgAQwWz6UwQuOaSApVtruSzTYNHAGMFd/FtQsUAd5z5w5b8H9JnYu1312QjkZXVd
HlfPmS7usmm8ZsbnTEZ51ZBX4K+fhm/+7+UyTcMrbeU6TzZs1lT+LTIXpyTIJWJY
wd15ipJ4rPeF8Pk2/mGYbn4n4DEGCUYTP722cQeS3FrDeJQxrl59Ynl+uBjZs4ka
5MXs9quIJwErxQNbbEFmZMN7O7T2rGoS8ze9q9PPdXpbC5hrvcC8S42Y2PjsD8ig
eq0J23HyHBFhWpznvNVuQ47KRT07duPQE7Ndiq8IZX2HLaZ3XXM3tizR0kz1mKb+
DPngg2t/4wlIzGsDtfaA9qmZ+sM+blHCb/r2atHD8uvz1FD4xeSPEq9hc/5H9srn
vlAGIYuDQyZUgbfGuh4Pe4jtc7G+8K5EMSfhRJ3735Iv1WAkzU0E9HTeVIhNp6sj
KDd5Cxgc/b0viOSAYiX9mO6wjDNTpBiaj/3J7TxU/LHL1I6nHTYVowrppKURdWhy
3HT9senL0iNhzPUhbsUjbOxooQsDQQXoG/CHIpJRkncM3sEZqVCkoGE/ce4Rcclj
z6EATBNmKHYVJY9yhA0i6wiIXp6bXpis1eLw+wN581q8SAdqcRqvr21pvkknWsA3
75QcuBF3MnsMzM88NIKe+fkEBIVFwWqdWNRPNAWYSBI25/8HXz07+/Aw8GOvCtXc
omYSF56041DczvdhhUiNmAWBsc8rpAdXb6qaOcTW08/Je6ZBY4xWTaQH9tAoFuwL
XL0HOFrgbB7GTJ7Mn3M/D1ipykl3U0auC5S0gkj03xKJbrX825/wutPn5VYLXhJ6
xPzwho8w2R6eBqzHeQaP77CP/SGzCojeEAF65RlEtZB9I9tNTipi5CdsF07LVFWT
60LpjH3J0ts4DrMC3goc9RchLP2rux3EefoolDTXrPISBsPg2gy8HKaZqZ6JjWoG
d/rKQO00alo9cGqoHa5+pKXjfEqi3a+lX68SgmubQyYbl5lsr162O7YAEhp/2CSM
qVDU7rMhkIr5409SD0m6mu5FOq9wNzL9oxTHXoB06467M91KgCIfuZZbynNiBuNt
pCbn8jDd09BbfpfX7eXGwTRYMLk0naNc1szLBoGrfwWbe+EOci3fvcNP047+ombu
U+0b4ev0Zy56lU2e/PWdojrrvWiBJ6Oy+Y1Z7Lq45PknSHRq3Ei1GElmeWSKuIFu
Q5gGl1R4nLmGFUcY/0crIWippYUbC2wdzImbf0l9c8qPO1vYOZ89ChIJMR3XPd13
ah+DbvA/YvQknd9w3DpufKH3Ew3mOWfup34K2RtMxemHdl7I0E8ayz35ozz0S2gW
/C09BsuWguwUQPw8ZjAOriUU8wFzMik9nJygnA3zpKhAYIBrc7CKSj/lmSSbqL/1
jeB6L8gWIPCoTpbL7a+kL6VOlEOlX0g5EAIaj2AtiZRgvvgwJQDy9p0QksdMhzsb
O42JinkWENYo2V2CUHG3hSUCdqcqvG7Fg4LIFfgxW6aEIHb7js8E/CfWJY8jzQzl
HUYRjS/Rwj4VEYrsh8E62a8c6N5LZF2tQbPv4wMqdpii3o0gM2BjprSr6ATst6fe
yThFZcIoy1il5fzur+HexQNCxjZO3cZlMhTIkereWLaWcvdgG5Vbhgy5gDpjegXQ
nHXGwPSLhOx99tbjhT3NQ7tA5KGZYQbl4/WEsEkWRig8DrWexo+MqA8w4vSZ8Eec
gK/n+g1daH9JaItVlqQ1kLzSAKVMrAwl42zu0E+3vLQA9dipTjMFgiT118HLl+PR
kSw7XOipVohWXtlZ8HlRAGoJti87UFfe1yTzEIsB/v9Hb+nj8ssWnAdcskUjhyQH
9fZjNSx/qT2wWCZErRujs3Dw7cgqgcqOpLOF50tH3EvuJrKiD4Ttf4KOpg+2JxFu
hemkBc6pStimjAdP/SccXAfhX8CmcUg9mAbK8KibppZHnAKGzwEK6P5lqOSmKPwe
UBU09WAhKyAftjn+K10QFGrHCWvZHAV2sK9logrKK3HMBjorPqvNAo4i1WMaNxEb
JrEi7Z5d6N3IH0lXNEnQ9Fi8+M3/C+lu/6Xy91+RB2Z4tzCOkeNeyKoVknn6Vn8h
wNqodyFkYXv+4f9AJdgDIFf7FdI23xpSM/V4/sa8BJxeKYmgQsqD1fQmiKjxFWqE
SLMyC4MWsWhi1lvgjnRRCb/S1LKwWe4nK53wcUbYGOekNKnwSGZrEL7xPRAsRbRB
RHUyWEulHrU+Q+h1ym7yo7yR5X+tW0dpBc5wUN+3l5RLCAqFQiDG1GAB6+rGcDN/
Nmchr9gARuZaMMp6iknDTmxkNx/tzJVtxS2pEPTg8f1L+n7fwv28iGdakCBJ6yXo
rYVJ+ekNMzNG+AIQBkYC60OI5LdPZ2KmD09ke88VI3BIWFYyfcHZAEY8Ll4TGto/
USQIIIiiwnhW7H3cvC5YjAm2mbJoScDXxRruyz38v3iiBK3nIKFVBJlUxufns60I
PmWSZGtzeMkHfx0tKq1zQ3An/kEV8ptJWsGDRIn6SiQbYPqgz9jGnBJBooNDRzg/
cx5YQLMSYA0/8nMIHBvptOHN4ZbS+qHB1l01u751Z7kL/Z7zoaz6w0IduUx8vd4t
40WN59f95iIjXev/UXHncX/DociMaKORDyQmf9+ZvtZaD7FUX3c3fD6vZIaTsGoL
tQwH1ov8ABviPUZQ5OwVhJ7XmUSx26WwTIY/xAnGwIc76ftuKY5gxNFMEK+BfU3J
/BcEEcyOKBkv7TXS+g3sjtPO9XXsdxrjKvUDn9wQSPB5Fjmqxynjc6W9yfindMy5
xkVuRTK1IIQYW+LeUycqmqJzAAhfZWzAOSmNm1hzvOxwwII0ts/4MkykHZ32M2e+
wFVlCYjTom8Ap52iRaqVQOywO/MLFyMCRIwg/ENf+byjKdD0RNjWp1bs3bs6Y7C9
Ui4SDch5o/o8HQfj5Hr9U1IKKA356/zGrbPOTJLufenihXEC64iyqhK7H40suEBP
fGSoH3QqheqosAtUSydXvzf9CIrfPadZlgfkZYFUNh4qQdkRrUVSwFQ+x+SHZf3M
lt1UCI5ONqu6dIxXGPuFyAElNaKKBzmaFnwyCpdIu3EBFDrbwbldEffi+gSeR6jZ
NX0Z36g/TrkTnqMNktdJqsiaHL9bPdQu8rZV60btJO+q/HpSFs8gbNppJB3zW81S
4eB244hi7Tu3Dtnc+PaIgnJwmM4qsvbA5GX/L0AgCjCeCbdyQouipBqwjynqwCIG
mCn8iZkf7+f3HmKzxr1xhPaWmGk6Tx2BZyxw/tVkqsVAbOTcIW0gvKqX6Rs2a0cW
u52ywLSWjoKoVGNUlkLULfUWNJLoT6u7nypap6YHS8xc9iGIh8+febE9Bi7k+93e
ow9GiHPtQ1Ia83b/DhfvPFh9H1Lrl8V3awr5hGkYICoSc1A/9qdnS3AZrXJ6T+V+
Mj/vnKSba4AqmzIKosqoD7Vn35959fCERYNIWxlgqsRkH5ZGU2YQ5pGPN/Wujtyb
d+6t2ppIoctzW6mbAxN2P/ktsSd8Fgp1vsyGwKzmRX3uQ67My5eF2StTHmKX83vd
0QEOYdKetRidJRY1Sf08kS3/X90BnB5ApOxKgsBtjO2++v7/mQt9xBgDwjUCrQFF
zQLalmlD+2N/XMjwqDNyHXMc1Pr7XnYNxi49NL/vKfFCwxldk9GoZ/AHz6iNs9sl
Qhz9FOSrvH8NSHEXDu0L230z2urgHoSFRkdn2mQvfMy7ax1kxrtmFJUx6MG+D4NC
uXMeI51Q2dFwPn190y++Kj325t6AMvdxJ2msB/iAKzcUV4cmOhKhpxoOI8mmgUEG
v0jPeisBHoh4R6vzdw4dxffC1uxJJiTawy3hyvHD4CxDmfCyWhpx/CeWDO6bmd13
ruh3PkFydAsyMk9OiLKl03b50t62iFhnk/QzKDHBxfB96HDWPF10l1WLNe/SFCnt
8iMSCBhO1wcKtbpLT4xOiF6TNiHzjWImUiaLT8EL83FRFXRT2lvKnNB+E0enevoR
heu5dfPjNIrvcyoi/TmiupKMysCFkhVCJ5x5etRk+gLcXmpp8omFcwiz5hAEv/yE
AFRtdkCmOigAZ24g7ByoCH1zhKMDTjnONCucizGFSzWuuTVHw6wvV6/YvSy9kflP
YdcuiOmoghty0S4FWkLq8PHbcI5GBLvSFA0C+BDVEQAmTAu4Gy33ask9vXMt/TfS
MDpgspGAXxaK5n3ExnjYdKlSvOKN/R4mUsvW1UCo3X/g/MCIAs+AcXM1KEf2hVX8
iakCPpvlWluNxfV/yyQVvuaN7jY2mFG8a5uvzctb4t+nNdFLHGm58JnEJzs6EyRI
EfbZW3Ho+BXGqJ7PVmOWCgHzF9Th/5/dYz/2hG4n9k/XPKH4kAplu+NFSzXh4SYj
CGFOYckKpNx8VOjWqRmJpBplvp4wEfOUmM8OzO+pTgkZK9diC8deIBgYu7cjz8MJ
gtNoRf3BPCFvQnhS/bbUM51RN3h1cSyHA4O2nuYAOQv6PymI7nbC6vSI+h/Z97TA
bTRblEz3kBcfkmUVM7cIjZDIxuamlqBJRzJ99PHLO6PbRbVZTfxRVQVrMUlpg/kk
I0GDLDKsxcnHFs9Ts10eaz89yAqv+UjFHMVui/Su/DSnT1v+xhFp+xAT0aZksZkN
NqUkdIVpVc6Iau6xa92ImOwuv4gd9jocYBZZTohrYbPkM4SmonY+APObXuH7S4bU
2ekBPbd/oUi43nSikN8XJIb2m7TJ0FLdV4VFkkjfnFxTVKrWD52wFIvf50petkPZ
n8FaSdYgePBzgb+QP066KrbS3gDulI+pG1/eUSFy8j6vFQ5hGOEdthLxwN85BrTZ
E4gXNZyC0jawbW4EZxbx9P+a6psgiGEsTHzaIR+NxScGMjwL95hfNucudvjhIE6C
PVfS5p38IREwjRy5RGnjaKR6OEMqLylQoaSzHA2IcVeRftyZdgHFV0WJKl5r98rr
pQY/YreKjgoI/aUQ9WEIVR8FjzX2MEqzes0T0pUBzVILuGUa21BFl92H544C7xU/
B40mSi4qdfPICK26wxXtT4nnlGZIl9T5MT2lE6eqjPtECz5zJp7EusXIqZ3mScg8
5wfD1Oqhw+leKjS/ZC3/KPjDP4JtujKmKTn79il6v05xUd5Rba4EzTPAeYt7mMkW
lPIBM4/ki7DfZVLKDnzG72xByUWCSs0oRRe5wiwtMNRvA5V35TuhSdBrOpAI09rg
vF66XBFFDEz/3AUmEu4/RpLDGQ/u+ycL9oER6HX8n8eNm1WJG9OIdgr70oh/mhxv
HbsgRXzUXgNaPqVIYDS2RiyvO2lHKl38jo6aJN8HUAcWuKcCmGfRxJHba0n9EikP
iPiScH0ZUxWRMMm4vLxdDYjSx3iyV3HNgDA6EgguaXH+Mkm/QuDmaRp0B4hx2ONm
vAAUxqHmdjU9gd526zJ+QLC23OVnGGW1pHVWC2B7/BKXoSD3zslZRL2fOw39YlHO
lMJ0aTTgdliVcPPDinjZtegjqCastSP6DdIUvWAMVU1P2M3E00FzKjKVry/qQKKg
AJKBCId5Y7B7mj+4OFnUanXHy7BwVEoa8RJc4GEeLZztqOhKo1nfQTggaxGV5380
j2olHWokNS4ROBspVAz5Z8UMlOxZCPtOrRXkjMd6sAoYnGE3lT+nCwXvwJ4YQ4Ae
MDVHpNxTXuZCl2ygB7Lk6AdZVN41+6D02iyoUrgRh52dC7xKwF+JLrIrL9R/Jpai
Dav7xcwNOHu39yetP4rJXuav8ERMB9UoAz+2FyfZUcGHKkBWMfeox5wSVjWZcoOx
i/O3q9griNCdzpi8i65VY5qbhetsZEwx0rRiRXm8mgzzIBiKzLKSRcVrAEPpJNYe
lhvFra8jR1ZhBA1K2GmcwWVjH4WCNi3B0IqIcsGsRHQjd4XRpiF3Z2Y1F6Lp+Njm
ftpM9nwziYgS+qWICBIcJxOMNUQ7A6ymAxrtcqBwuSpPgKTrHepkNDl7cymQdCqd
ChnfoKaehX19iDyGFrv1xtWRC5E6q2dtSKp8IW4/UogvQRrv2wdEdcrRuTnZ4jYp
kkIouzwLRbZLMGSR5xNKaXKYslGbNordvXMgq6yULqprqGU0iglhfnHuLQ/rAcMf
SbotoGXaQ9ZNxAooL9qZydUL3eXkrRKkv4bR11LmoB9QUwYEsjVnqaGATOMA5Peh
ixlA/dpYdhHb6n5LSqprx5SjgN++SlXvnhs+UQrJRBji/IDsRj2C471jSo32FS2J
faMICmtl4qtqkVgzJgDz0J5VOfM25Jg+anVqvq7iaHRSIN4gvHGBpx+sOzM1JUTl
G82hWbTOzdpGxYNp9VlnTk7DPLw/jcN2igU+fD5DsmgKog2ayQmEfviGiEvEzXr7
xdxE61+haYPwSDuPDeGTara1B7Z6b0Rmbl8k3UrmHFrM/w2q3CIe/D2mXwuuXiXn
kB7EuXk3w03zsW1z+bmVZ8JuoEpDETYa7Y6RePGzJGkaamZzXOX2J/rLW3CAGw6w
gA1nxiQpuUEi83+QFHspaGCEydSQyHmmH7/KS8GlH9Z27OjTnCMN9m+QjgNsM34Z
GaKEz2TdqY2bY5pwkLmdCz+Q4H0oM5riXrxyqSR4+R0mVE+82kTNSNPoHFoBz4HO
048Xdaxrwd/edHK9sgQbbyxoPURoFFVkG17IaLrCFeR7FVUDiouhGbVvUJBHjqcS
Mn3Z2MWZYk4Ui7dU7cPpZOdDYzfPbOWhlxG9BSxXPLJCVm6QltZIccX5l+OyGtXR
NAiTlFKEjCHIag1t0yD5O3fuIkI7k88Gg9x79prwHYQ+OE5oW3dVXU3VNquV+4SW
P1N/y1lmAqXkf9rERXH5JLZdexbtg4z50m0dAiL134+32Ndl1+nHY5Y7HHLzg+FC
der9tHI3MW6xjlgVP6UI9sNDfqfDH0QDrA/B5tl/aE2sdvlJ6YnedRsiVQ2OqptQ
iAqw5DgIFmS01xHIQ7EeUSUyEHXRpoL3pWuA+IxAkIIiVY9J2q0NdhHW2c7QN4lv
ikL2kXuI7r8WU2SlUJe9z8it/ThtsNt6DKKx68caHbwP4G4ddmRzz2ZqI8Tp3P8t
u+u0jVvVXgRlge7E5Y4r4bJ/NatKMu5t0QFIxwQIf+x6jPIj6dGhl0B1kAfbD/21
v7LDz5zrLH88M6D6TIQU5xRp7FlD6jPyzOxJlEBYTG/v+5+pq6IdvnuOp9Swc83G
VRC49Ma0Gbm1/WXx6Jle3tm2s2G0yRStbHY+57TxyNl6BLxECU8NrpLDNFNAsdf5
+/d5xFq4fXKbnKmwiHCJGcMooUMkRNV9VXqmf3+0nauT2QXCdCLUU5dt6R0Yjx31
F1WF42+BE6eDX84E5alqKZIGf6eCagdDdFP/9u+jFllbhAiILQhmDP6+mZQqhCPf
RJqDyXeZwnW7aNqq3SqBgBC8857cmHI3GjxypsFz34B9qro9HLERi1gzplGTQdTe
F+NJC6Uhf3LPeZivxl6JmUKFFhT6jTjNEo6Vj8TnUyryW3FbofIx+mKk8qTB639S
UQ3PfXB2k4jSwzlNuwXQhNlnEKjqdYSFIdHT32uBWR0OiQ15n3ElE12OJ0rKYYlj
r6Wh3G4gdMx9Uwe9AV3W0BN7Huus2+YqEIzZkR/j6JNBCRxS0kgeo3t0cfev+mVK
kjX8UfnC9fGKX8ZuXZvqVbzOl3K4UbwAzXuJl/ZNsPAMHVjt2Zx/T6fv8qbSmNZN
+uCkqSr+l8xxVn8Pq1NNN9XsIszo2P0ns+6JrH9rpdC75/rS+N7URabEw47GrXof
0lzfsLlIgnZm9Qn/zeifLKtg0S2pIcTL2cFuz7opSDFWvcp0nfjeZUnYJtQ3Vmh5
xPabLNsUEWTMwZEyzNUqdSUVblA2TL0Ot02sfyRQ0IEd9KKPqwoucuTcHXS+tDNy
jZqfUY7Wx1krD/QyFjfe23LC7WUPqok9YS0u1pCx3S1n+oWaDOA229K+BYllYusW
axCNHo4xn7Quu+hRFfr91Lki0uqBki//mKeXWoarZjPLHXz1gB0JKDy2mvH0tFCa
hG/oYCAVvJYea1q6MeGttDEpPJoSfV/BwU3c59va10fKwAl22tdbLTMXdvAIT9jw
RhDimQyKHGlhdEAJvCW1pB+gT4ITq+oo+w3tW1xqGkFSc11PfH0tJ34VJotXfg8H
l7oqLMAMUeglKo1LmM6SsWaqfDViBuuWwfQgqO+j1DRRSaAfngKEz6hf36JqYaqD
Ofb+6J07gmSnmFyUp31SCEderqYYCoVOoyCMfAY8NGNQZHuJ34vDQKediDvuaWua
ehA1i2G7YwTrlRYCjimA3EVR19Odu4tj6sOkXG3NZJsgCWi2jkDahQ2G+h701CXE
JPCg5iTQaIxT4GO6RRzVVmWt1ksKTy+lKx90NsJDX6RfUMi2M4nrpJseySP0oceg
8NWRWnO6XuEvpkELHNTAhCee6/D0Xnu4jzQOsXua8I29YC2fMDk8CoZb0xqMl878
7immWFkn6KuUt8Xul+u2NIenHv8kOI0Inq3zLSuIEBbfXLRvNm23KFWWYDcsiXeR
FLv58xpNQX/20I6xOrc/+vqp12jlH+Cd7egzZaJYQLWYKiFT31qDHAHZlTnwBfPs
DW46AD6F7gCrrbaLwrs645wC5kSTHXzdoRMNB7LK9ZdaMXQinGCJdeC5IjECy88S
5Rz8zMD1rIb7uQD6xA6O174D3lE/kj933D6oAcmV+GG1xoRsXP0iQfc0iSMEO4o1
4iOCp4MyrtoIqp73MI2NdS70HFpaRmAaV/s/pUcgUi01vW5jxgK2W7Q9suYdR+mv
n+gDTa0JZ94L3vAVzY9e9tw1fCifhHrfy3z9Sb0cm0hK4nPKhP2+sLLW50dgiN7i
/Ap0DC3qnyU1KXw4rJfnzIhFTg12LjHTyDMeC604Und8DHhz7v3kVxPnsdvgoxH6
sJrMmFk2ERpAU1DuTU6fxWyU/GUHqRANhOv9sYDnNmPuXHnVZfkG+U6BK/XQNBKy
2aV7M8HnOUCnKP81q3+E7Ik/sZtCqYMF1lVGNWFyoR2O8oO4FDO0cLz+NSkYXhD7
7fi91gyEgwEV7edU1VS57SlOFgADw4gkkDWoxwS4KdJYT45w/r2qqAyAcnCFxW77
3Ne+RuVzFGwQV/EHf2URpQQTX34pzoMoD5Jg4Ln0wCJ3hwf7RoMlMPgxKGyhYl+g
v4Uti+OgldwDGP1Sp8kvPKkVnGvOU79sLJJXJZ3lP7W5hp3gxk73sL2DA11c+EjF
qad7ER9e4KBaEyhDMZg/uxVZfBWSMEecDQWhxS6iWcnbaH6z0lW6paVEfyH0O7Dh
CsRxPdgRubCVeyf18lXLyQYPFNzTMk5tI1q8bgnPhvP14HZ2G6o3hjpaAOC9wvMy
pznl8Mq3MHpo3dhBYCRjUj1FiY0Q79IM5k+Plyh5Uv7D6QE7HRSp4Ju9UIl9aYXs
XJuwfTo4Rhql0A+FBPK9TUFaT/irQ4OIL7c4nmQX5v1WBP5H6ssHvYow9I7Hc5gP
AhXomfcFnYvacrKy/v4W/HLyxKH24L4S5NZkn5LimMXQWJtfWBJNN8n9yD4W28rn
oZAsnowSel7uYMfultetpMnP/c+LT8gaHiuJUtIsEAABt0Zuvxkg5b2KTg3oVreq
lxBebuKgPzUCWgR2s5DjgUZI4nHzgfqdNCHcz1u3WRRFPAywPMdN2LMiE05i3BJm
sciNCwoVDpi1TE9rVA25fs47xN89JgeDttVhQBqyvZ2oGHHMTvyx/VfpJE5z93jT
yXZgiohDhTsiC7BWSYfnLZSQft5n/r75vM+ceFe8SPuqLXy/C5o66GzmtbnXmtBZ
h1XroqEmRoweZyfL+R4YPTBZ0mMnuixjYqlHpw2IDI15B+lnqzP9WJPlHV8sZsiY
MxHfl6KTYdY33ZnRA05O8THO/tM9FloyCNv/CoR5bJiCrPz/MSyDH3gxX2fId7JL
h0b5fgzHdlW0zbG6EvguvmqmwPzeJz8wwYQQ4JRq1axlmDm0a2zuVDp9gCui6MEb
tADIIMbpr/pmbbwhzl2VtXuYKj4T6j586AN9VFKh3z/QrkX5ITS2XuH6dZkWH2D5
tHBr6gNX3LEEgNo7n1MGbhplG5weqIz1rwzuG7z0z2cJw/r7MLI3uQvIRlIk96A+
fCT61cFRgAlcpERelpV9Eh4YHycE4hr5jncBvCIEX3TllKzjDE+7XtBkOmrKHIwG
v8nxSI6Q0v5AX6gyZVJbxc6w0s2QA3SmNeGvSWepm3eEtgKvkKOnIF17KeSD9O2E
cmD+vAUADMoTRtvpKDE5A4dyJhbmycISUMxFS2qX1KR/EkomDwNznCzguFWnH6OO
+wyN5oQL9TI1Prbp+JsmTeep/fELHnyfKXuZzGqsqIMhcIi1wxNkSmDnS08oD56J
ujL7eo7b3Uo5jTGFaI83C59wBdvOi1y8kF4XMqXkZTEZ6oHF0WJgqPZQzEMCoC/J
ybnfap9B58H9KZVww8/igbeFJPo8TX8a1ZTpYBEreR252f6TNLkA0T1RsnNOg7/5
/MnHcI88bMNzD0TrqeOCHjs89JKetK0Cvij8LZwrNg26li8mNnmR99z3OfFTx2M2
2puqO9N/6hPSxISxrA10itHalz216IMClgwyJupeGCrEBhKVW8fbOBXi/pGYqH3H
3mMM8Ef8sh5nYsYLNOTKa1NVpSxT7bs07PHQjrhm0k5ERJmUTfm5wLn4zcwV3eA+
21quIN9W4c/KcCDByPZgG/Pk1gRd4tO/2RRA1BkP/5REZl7JsoTGM/Lf8qk++GTJ
794+Ftdg7aFDI4BUYvFzSa9YFsHNFeCF3VThFDb2ER2Aza+tWB8V1mSSkz6EDGs5
VdBiXrpH75bs6+GlMVQZrQjLkfRTBHE52CjG6ivzJEwyV+GhOcBoqP2mtj8TOcNu
/8AQrwk4+0qwn2K4jsaLnoiVCzhLCtZGR/5t6E174bSAVagHalXwEr9LEzlh0Six
twDK3STh2LnzpWfJaRssXncnPcho2phd49ngKdBsi6PcAmo+5U2Q62ZXvIvg6p4a
QE7QDiATaPC+8SBr4ovzab6JDys0DCfgPsJPxJljPWjNNsNndkWCRjr4jFGJifFJ
f1ZTMgr9g4dKp2kemrccBi/wkOF1f7039qhqk4F1LdhAOehCINCzizkRlczx9Ug3
IgQjfF/uwKWqkCbVNE2DFzJgQ0a5xhAktClj/Qy3f4oTsnnVqTIDfEFmyBzH1L9D
4lc5qQbzr3/d1zCaIsnXoPEw48rzz4vFKlj0wZLpRzugfmeQcHa4en84OdPaa1UA
QKiLTHsVxzEAStY/s1cjtIABCqvsw/leMC0iGiJ9ZcXHSRsnkQSqEIKj90YZvN2G
wT0fOKkhWSLsnJ68VUsGFIubuaWDfpJRNugVXreeNMvepz9Sc1GZJy0M0ut+MwW4
zcq+1VpqMC6xOIKx6Wx6Qd+g9YPwHpnP51Lj6yPWnw4MJsewLXSp5itsiFMDsydS
pJEUVhaBXt7CrZeE4sf4kXnNSGyn8saKNkuhkcovmbKW+XlYGljm4SxNzwBNLu8I
25tHE2VNMOtNahsQEXzSZjQwZqtBzzl3EevacwiGNgbkxb1et3i6zPZzRE+0oVpv
vcSStjnhcAEBCez+qbuDaEhbbnc6UgVPuv6w9uSfT/L/RofLlSal/zZ8fJcCerM0
LEUrPUdkP09KoZOIoaXY/jpxwpOcCt66mYBfZEKyYLtMJGjjpSkU0MncbAqpz1/I
GUUbBHmz/jOJoJbuM73vbIiVrkry3NcJy1s6tRD021MFQn849CDOWznk+3sqT8Ql
T6lxxUjafFXYxTvw2JyfGT1qXLXB4uEtdn5WQGCrxZlURaO/Xxbz1b/YLnYf0rkK
hldiEpm39TlosyRPbtAlU86J4IzesCHV6AeNRycJz0XgVXskQgkEHdoYzRyAxl4Y
xPmSqINTY8mpjcwR0Xf7W6oGAHkuBLlKTqxjFDN6YCe2T4h+dJbj7ZSFGB4p6IhP
uFuGevNEqcHVb5xMmAMw05SmryRe0rcDM7yLMjTL+MhYCQD9faZbYjeS1iMYeadk
zNZOeujIM1mlPDTY7g4N+4zfWYDYPSxfgF/p7vwu2f1OvjDAAAJxd7tgxD4LfzUZ
HTwrZgZkH5tel0LD6u3sxwwV/eRMH+RWBsLd1euodqDKy8eqnzgvbxXr/jw5xnte
Vya86B0LgPf+dia+HG+4MDpVHBvdl3AK9lXeIN2IO0S4JW0Mv38CeESkQMuc9MNj
lPILX36eZ0kHxu20vMaJxlcqiXpnZJyNkOUG19e8C7GSvXy1/bzHb2TcJFobbwCv
fWqaupQIU5KGRO3/zigUrL/5x+M/kr/AIXI9Zxu0f1rr0fZ47oYA86qAGaL77lgc
4nodDz59h4lC6nox6R+02lUIkuEj3yGh6Mm73ow9Gp5ANlbtMKmJR8qpxS+wnOCw
GbzoHlzObAwRr2qq9dj3qSlBNTYCSGlMXKhMMigieIO3FOuLbn9u8r68a/d8U3tN
VD7UNgFLNaOsLVsN6eDFpJM0upeRtuDrm6w1JD9UM7qmK4blxHKivMDT3YilvsBn
83pa1gMWT5cldEHTnwO6Diha2m+oXca5MKx53eV6vBlGw4pkezRjXng3SzxINoqs
1S3oF3RhJN4x4A3v0NsYJoCZy2LxRr/jINWonLSUSsdZymGT3kjgZic+jnSNaF/f
jdk4x9Fb8nEHCvEIF5Cg/9HQc/WVAWpySj5k2pdpzY/RuTRuJ52OCEX9XjEY9YJW
bNX9Ru37YQyeekblu1sC8d0JWNpWozaLD70sLhEE1Ub/PfZcD008JESONhLoprzs
6aqKT9UrubnZ7sKGHYkcyyhugc1b2+Pq4VnGPOQzymupFABlu8eBUkWK4gwtJomA
6XVXC8lN9hQtkeDGF+QTfHZ6b3MzGHaO8Ly5WaGUzonpWm85lqZO8HO0/xJ5TVxn
2wsqRmxVavYVdJWMF5XMozXOrIolHReXETjrrTlZrpNjvexB/+U9ZYwY/0ReVfnj
wG6WximuiN7K2DSQt5YbIJ7uPTmaQPQwqCQT4nO/19/9pDhEdaHOv9Q+VJC4W8rb
Mj7NyvHVJoFLiP1SYVVpREHyw8YVCRbSJl1aZjDfWIj4OjQVS+ScSvGNhdj3EXal
Z/bYf5T7A1ZakcBXru0goDd5uUvAvBTWhMU38cgXW+K5SNQeYC3Vlw45RlAgt3qZ
l5NMMgjW+fjogvpGoJ/2RuTuJQUS4EWWlF56gjfPj0YnGF1WaEHLpuZaNBDjcr5M
yzW3WoKrp8pC8Y6fFILJf8myOy+6t/+9eAT0s7pk1xTaVbO9RTc/GvR/tTLbnhl0
rmkXyx3Hh7QOMHk1jazJkB3AE0Z/EWv/8f0T9AdNvtjpUJn/60aPemhfkhbnq22b
HyPgpiMb+v+z1WuWFZrFSono4ocIwP0kNRWJfSDFGGq3a7lLdy6tUQCbVE6hOFPa
iG3xHo7nCCKnkD1fd8v0Bpry9+Y+3U2xtGUBYBhIpVBweuk3Au+oTeSwb04X6LXm
HCozhutuJHhqQlmDEHObmgwSd9fY7F0/uIw6V9qgFYau68q553sDlJ1KKc//jaCH
yLblkt094Klt4HdiAjaxu4PBrMDwrPsWldsgVoTd2nbwI+Qdxxt6iTt3qVMDIleo
VFOEQyMEfGk0dUy4+jirI6kxJsYULTUlqJObabIetWBwa1tiE0zMSd59aJSqLQ/9
CNjaZkIfGsNor9OP1DozHhSJKHM5eh1XpFQeXmseRNUqeKk1Bidd+jEMaNN3bhyT
koGN8bWXXlanBgVZL5CunYSV0QeVswFrudAuC9CF2q7HlBdU9ljwvSzzHGLuZ/C7
877g3PKwvD1S9ylSiwaFHxt5s6X3xPdvHZwAIdqCCvQAG8+vxbU246jC1bMpyJ7D
d3vEQSBBvuVFZKrHmDLTe07IIp80DEpbdlHZ9PK0r8TDKDxR3N0mx/DqxZyIYzVC
vj06AxUC7KIeWSKaH7A0uvAZ7LOdHDJm/ogNAJTaNZ0v6FroIRhTeY22qe1NXVqn
8SIPHvyp3W1+sB7HKcjACgMqeC+ym7qW1EG2tqiJDP+EQ1cmXK7rXq1OFlr20ySe
3HHz63NvMrb2vlxLiB+NcMRoZukt8IMdPjneOPmBSCLGBhZZsBgHeUJxwgCZHVsw
N27iMImgjVfBRi/t9ts6pH4cWUmTElA5PUdRr3abnm10q6eURmiMpamFSgQlXhK9
22GbLLG9wOMTl6rjz0V51f3ZdgPhVgHSv1jaF1vCYQLAdGcQaXM1DhydSp0Eaq6m
DXzGELHwlHi7vBAOQ2gi0sZusAAokOjlSqghV4cyG9Dm6al4XQO6nzszK2f/Dj5r
MByOXk4lPbv9xI23v925S2ORCR+IqkPUNHDBeme7t7umbeYDeWQeTlmACJG0O3Mg
myTM+5hWnDZsAXrzRS9PV9BYLbx345vkQtE72Lc09GJPVj9sSQ8yqYBlkn9BppUh
RaV3bgx79kQK4MLaOXTEBrXS2tyTques9VJ/Ex3VLZcDNA9gOqFhgxgM01HlKWdK
0MySj3KsW/4Vaku/0JJautTu5/ABBKfI4PCI291FxDd3h3bBcDAqiSk33xPXWak3
fmh2SVewjRgB+vb6HQGs4SH/LVlmr1PTUdhMaRbqbZCdBspJ1g7X2mp/Rh0DhnSn
HNtWRoR8ry+xOY2MVFvxo9R3PZlBsFvOdd2+xfKswI2+DmSUkk9Kl6D5vPOhTy8c
w8vZG5B3mE/iN7JrQt+zkdMzUJJPv4f4EdBEEkj/ML5qXHBW5GpdTeCbkfNCRqT0
5B3OkoMNntAYXYFQ4k7lOFGwvZDvmBHy+u9V5pLK7F0vRCXorearwsWkyfjuAU2X
f/jKDqJK9SCtS93uchhhhUHE8ssJY28E1McMaCktPIF6CGiquv0IWG/dPHy9XIuX
dBhDgznf1Ba22QMbIQSmWFLU0Fr252cS6jR0eD4LYNmX5vhuCIoV/d/yAoOsJ5gM
CqlSjCTXX5/u9xb3OYTdw/i8V14lX9rA1HrxHlhrsMZMbeVVAhP06N1y8mwgoi/N
aDkxEPE5sU8wcFY4F4MDyKps4g1ef8PjLx182lnX8NoLStOw1vlgENeBv1V3yg8U
r+J4Jm6B5IqCeDXeiEtG7nzuCjMyK2btvbHHYBVJfAbv4ML1GLn9zlL16gCk5LGc
Ag4dpYYPtRFE/1oQXtBM158p/WeQR+mM1fuhwCXfCCkuOnBM3KoRxAeb46thRbDY
ZfZBVg2JLBrs/Wim42nJFECSqAgHPb3FXrS0gptl3M7Vmn0M4hhkBwJrFHtuY5d6
CPYM9C2PHqWGqSQX78iUm8mE5ey6G4ii1o/TvmxnNA6KJj6nGzX76RQ8f2plIMgb
4/8uUt3IQL3g73Y+8yfprdlAIjfPnmA7vHKkugHKb1jitM8RmjA20IswqwfZ4kr0
XyGEIRL8Dv7VlbH3SKlay2mnWt03K4ozf1fxdXJkigLgmT3wPQGYPjXClQ0Fm9G8
1GMN/xal3DTSaA6i8hnRcuQqnrLjKop3SqQKwfq9Sxbmfd8L0mHwjOWGNPp2MMd9
ODSfGJOdL7PvJvWstjy5WVhnUa0VdMoYlp5HcwvgMWmNeUETwTaktri2Lk/PvNS1
+TdTJXbiBs5Vb2fWdKm2YbdTp3Ak9XCLdvUdXsDz+2UYt7ZHETKi6U7Qr8NzxcLi
ziVIIO5mF7nzqE9E5N6E/hZDem9u1T1qgnua2zPoyqMtIUukLFtnABH8T0wmE92J
k8tAxVeXmthf08/XxLJiX2D9j2UKZyc79lrwBzEvCPEhp4fqbARz8KUGbv9KEjTs
Oa91IVAFNV+WBzEfPLuvBZZe16fS5l3H+0nrFrWw1t7onT2/Rdqb4On+Pn343hw/
zSN2KBFvalW7UnGZA11n78d9EHr1Y5feXWq6QrZ6bC47Bx5XCZeG67uDtyt8NkLL
vKBwOh8gJANsSAcRyA1A1LcJqzlRDo3YD5K8jkqtcEM9ERgFO+eT3I6Qx1bQ9NnY
I9C1cR3bC9SmN5DveMg55BxvMWyEXtlbIozQpyf4AC9/C13J2ruOwMhosveEEH0r
XmVlgB7nK82QCUvZhrKaOOCZwF7eN+c+HdwkfFO7WOdDb5g5gxMDQ3pgfE/YITtW
4E/6v9CapZ4cNqoJXycnrO8VJJxSC+RoFNN15Epx3yMo6ZCcf4mONIRbSDziSw2y
7j6DEFoAgXIeX1V6M29vJwCrUAoO/ExL+fa8QiGQdjXUCNMxpFVbhdVjDIJ23dwN
TuuZL+QEYlSUkvivXZioUN3WvRnP58PMc3nvgsge/QwVS4Gg32BPBFRNvDxdPWep
l0hHPiLfMP+9mMHlUP4GZ1znft4sXw3HmmuOPlX2BYy2q+VE85Tr4hxo4c0GYbsR
MDXJaSJFwf0vtOsWiYg43140pi3sO6W7JQK287FRvK88fZ77Q2Iy96V9s8M95qzI
4+3/oQtpTme08HUXSJEipJ96+wHNajirvAxhkI31w1vnX8eo4UwFkTwxmkqckwUG
St+tdBg4Wa4rCLYo7oCR7DZ3nVIl4MJC1+a+7mvTg5l4R5x3QXnDpVfoAzVpwnJl
vaPMlfslKRaMzkmqILBrpq0B/8gEDYXz8ikaFRNzYwzRjFCVABZnjh0nVlNqwoB3
JqDq11bgYcVHx5o/IEcIJuQmdGSuCZE7ZRzJX8yP4isxcjt0GP2sdQbmENTPMBaQ
HRFeUcf/2Yt0aY/0PF1CvROdLamQU7PSEVAnqfCCAVNQHSx/We4T1eTP0UaQV3mi
+JVh/QOFRheEc+tv7Mqv67EMhd3Ww1VU2yIc4ChkC6vDA6/9nXhEYRdYO241aMMN
SeitqcUALb5riwq+bdS19l+M5gKVOm1Uwvf96GBu+sjBhPdy/urHlclgwUiuCySO
O0DATUjAiFWCo2ii20I4zMysbuv61yY1VfaAC+SlAm31z91pDH/rReHmmpGgGxLP
tBvPBIyClH7+iZ4fbXLni2KsTgXHCm/5XOZ4kfI0nvW0DVGLh5NB4qbLMHh/F46i
tMuqco4p13yRpfdEdn+5DLO+m9RfLggc02EhDKeTTZlEiLA5iSB1j56mecnVlYIv
12qRh8tP+M/ZqUrTlTuxrt+U6bIT1yt4TGpSYbeHaykIFUEdArAHeN1Q8j5T5h0F
Ql0VbodIqNP2RPHPlViZy13vY1JqWm2PRiaBRJ97pSFaZcIy3veNOy5lpDp4zu8V
EIR9oXyDE3o98llQ8XkXLasNNLdM2IJ36q4SQUik8zK+bmk95yv4Ltl8FYF8nQPF
uZlhbpYalSPUh3709ipbW4ZNK5xTKp1utt8hAJh1ESouhI+r+el6/uz1iRh400gR
D4Y5+7qeR3iqbK0SXBO9XxJHL+c0aO7kKwXHVIo2WQxRE3iL0c0VPEU0R06n68y/
tjT1A00CHdhJNGF5N05Fv7EhrqQ/+TeOOqw4I3QVObDpv1hHzRmDyZQTiOpT73/T
UJYyEEa+4QHjc72CaaUGvFABHKSq6RvnXGj2moiFdXEl4ypsIm11+40ZeXUKJLKQ
jzESBw+dq2mJJ+DM9F2qPwXefPLq3F9aRV4VqptZMxzcK2BGMu2xUkylzG77shXt
dBCRuXe4B5q8yQwlhxEhv0npCqj7zyGZsL7SRM/fIaTQgyKjArlJhl3LXC41Eudn
Jt2Mrduicg8R+6B6/Gy6SohHLldzCfmPYEUjej04VkpwJ3IBadfC9Jzw7cN04fwt
MsPqQ36jbMERM9OKUC30QDARsN1I4cnrhy38Og0xBSZR6rxaA5NMeWlp9YMh7k74
Pc7anZErbNLHecujnIV7Z4qBdf4SB+YS3YDfJduyvgn4luOHnZmdmfyoQzSBtLp4
b5JjMPH6tU8lwSSBKcGhAmAGWRgdkVG3pBPPZufDJvnESRMsA0Qam/rUFKtuREq8
4EzCZ3iDR8DtdqQTdtB+kgsBDvW7WvawoXYfBSns6UtJzCSIoACfVRjKh4eJ0r4/
2rU+nh5wCJSz/Nv45BQEwCS9aps8u72SNYXNccC//bxdY97onU7X2W0MjgVjO5eJ
8MfqAQYyQYe0CU2Bf9ocRNVVF2Hh1J6XIYIVQSRfy6smr51Qeo6eLowUskAeH4QT
zQpLX03m6krp3BLUOtvHYU/7E5Fz9nMweqhq1xvw8a6i2L1Zo6+LpKf0raCTDBGb
MfWa1LRNVXL+Jfh5CIkKKJTGPfzAL7MbMgHHktLgMH6fxLYwxPXReuFKRDtOBKbD
O5McdcQb4gygy7iVMgMFniudjFRWen4uLHXhjGi3e60Kiax4jPXFlZ0OzpgSLAed
IWqcoafNtDfv6NUrZHDBsOf9MlKNiYkQL4RkIIv6huGNtOERjUPTz7VYfkcb/Ec5
TpjSem74vqgLxGblGtqQrKpu1saCy5KVjFrcW/svQ+Kdrf+sFBSulow/RV6W5D+M
SCGmEpgVnSHlteCGDIKqDFlo1oHZHbKGbJJ7aNC9omAaDINkWd6hq3/89xrtItX5
IGMrGh05dITKMo2JHgVV4TEG/Ahm9lEzuxMLAx8r7jbE0Q0PONgq9bQuuB8YVUSd
xDQQaTnbvPAjcXKkDlMRKPc6CKW/hGkcqK+veJS9R1ZmM5qDEW9xeJAu6ZcsVvBT
HR53CgMqCoYxoxZygbdMYgA8xBKBnIxnJrzoYXQTxnfD03Xn1REOXH4YGrKyPXOD
AXwvsb8yuHTuBrxLSSFqUb5udTN5GjCyMUtDW0Kdm3NasUl9xiyyCht8a/m0f4p6
yvxU1uTaKv1aDNf2DkZw1g0wfIyTqY63Clx0l7iP2kmuJykfEW2x1aGOxBJVQ5i9
Q1NhVHV3vqw4zTLjFjYymR/w2kfiziEG4neVRnXNFgeHf7707Hv1ePpQasYCJhA+
cmJphNmQkjybA8IuDYlwgnR3VkJLdV4vZ5UsSs9ApyOLEvWYQS66Q6tmD5Y4TA1i
8t16DmGIkKzTFWkeQdfXm4nEXdF51Vk22NOsbEgyhtLb9lLHfV3Pkf2DNAK7fgaY
nyIIrg0WDnU0aXs+YSAux8btHLkJzYHQGVQvZmKvH+yh+N6wogwVnm2iVwhDTC8y
HAjxvjsKxHFXkP6fJNH3lpbKNIE0kiv6jFlbdia4wcYIkbFBAonsr4u/EJu2FpuI
JUMZZZmlgeYQxb6NtTh0zX/jcBxoO0AEoqE50Ous2GDNzX6hCrlHfugwW4T+zSvC
qfUqaUkiyJBfTO23d9fuH72EnsM7Dd62U7IUzo34vL2d8HU1hvTYMzwzbp6SGLfp
Eiu6Z05gJMuYlqHjKySPelPgOQK02f6y/v6/RZnlSDNKGg1lXEiG/WbDRaMDVefn
sWJ1MqJ8BMV7UYVACk3dM6TtYOZc9DIbyNZgP10ke2fvXTxLRiQ3h9XPG2GWiVda
+FavDVGduQRnV2gJHIRryPtC+EGQgiQTuygVqQLsochhJ8TcAvjTakUcjjBrsBfY
rzKmi3wixc5goM8fR2ye+pCFSapm9ODCRevPeVL2yiDI90+xaNXJ554LqaYP+iju
s4t4iFUW5/PQyS0urk7i1k7qYQHyvLeQtWIXEN3GFeo5iIYAvwCvv7qGrCz/D3Ms
anSBx2yOokyZ69Pa9MlDSaC/8b2ACwrXLvzmBq5h9/wnDy2zxgO37HxeazlYjNfM
dSFi8YdvNktp8Bl8xpGcJ5cFWNDrW2KlxaYirAi6S2o4o9lSm7pUHfEzfJrBZmvX
tqrBbi5ZrluTmFSY2/U1z2OZ5uSqeffan9VHJsXIQoQamAUkGLIOKI8itvdxPMz1
Pik76JXl4+pMeXuUE3xAxXiYmHTrPgPr+vW0+jEu2TuMFLIBrjpx4/UEmd7T2ZcF
zh20wZIa7B7zruJHbrh4Ir988gy8837Ckp4W8mPgR5rq2YVaMMxbCqQcpjFfos0t
HtB77nOXtA+FErYk5Am3islWvVunNlnLf7eOqrzuUgtE+hmT2kxGXxFrPxm8f8ub
Uq7SdjSi55EkCMO2gUTG6VJ8/5VeaHKDQSPMDhIR8ZsCdVayyrvY/ie5BxKqtozx
JVfV/ICHEPKoeDvu/RPdrTyOtNr5yCGgc98zdCyDYNPsrRhUBQYNCVhQt46q50aI
JGRvbOBqePy/eyKg82d2HyNyjpelouxXQSJAzs+/wusF6WRVqm3YwKOQSqA5yErG
HGQIyyCFcdZiupVeEBjEydu5QgNOJmOTlNGHe9ifgAMHob8iDDBd2oMfy6QHjXPM
YLPDiP+3fN1yJUHMFAIz5Gx6GdoCY9Gba8qn0PW8gz0R4BBbVkSBM1wCGpOXBZcC
Cm1v3RghZ95QPHROZf/7S94Zy2uU0GLQ81Bst1N+eTaa8l7A2wRGpoqMEPGt8B3k
H06iQ4hLVpEZc2GR0BvAytygn4nwtxtavoORvIrfEK6hiQ8oPWpUGb1mNOEioIX0
lf17xwA29lB4BZujxy4hWUR6RjN0+U0SaQ4ArwbDqR0S3a6nh51zRTUNiXeUqaNG
X8yB0eRBNLVJvgZlAgS7R32CroTJ4pqnZTa9AnrzNBgS0IHJYRUmNQ8tHAwi1eLx
bvCB9HRiS4CAmr+TD+1LXL1ljA/MHKGf9wvvTWN996FJ+TEr8Wf3VbF+OMetF2W5
fI1rf+C2OYXCVJofZz6lwvB8dNFA2IsuaDDIVLjTEY0CG09dzEEuIwlZpbNJqJNO
0dmmVZZl7wKUvNImUy2LZ89JtoRnJXiLHPL0oW+R2CTwrIbLO46vTswOE6zyDB7x
JbAnjwdwdeBNtBkRgnB8YJhqyJga4xQ3j4clFmKnPnJBp6c0souwDyAo0cdF+j0l
L23SWOjAe3dI9crppCZIZRn6NZg5UdLgfQcilkjKCtG2uVVB964SKMkAUAH0d9L7
PbK/i6WsH/ncS3ETo5AuA0ocyRWbk+nSthpQ3yHUutMIQmSgJmGRMCi1Ip7013Ua
NZbp0NehcagC3MiRT/NVwh3vF9HQI/tJVELWFlMGpq0EXq84HWwNaCorw+zGFrPj
IvDeaZ4EiMwHbQuBGCpS9EeSItloZYh73xedHJXGkpzTnuA68yUJrY9EIka3TIRN
Chdi2QiES4dcnD1bRZJ5llz9JWseZud/X9LyOsettL2wBNPyyXTubmb5WinZ3LDd
1D/9kgIZNcMa3/WUl7MGcMlp3GiD38ZbPIvqjW0TPtjU7fa+wcaXUFzRmBDcz5+U
VGdUsyhzA8DUEpeSRZCNY227RT3Wzm9ldguSzLT0KMl/R+cVK+iaXiIl4SlFqUTS
tCC5kBn0Vc4t7FsWDOKdQ+jVzkc9UNdyKuG+bidQdplb2n5vbDA1YGtY4BVNMssA
KXu/pIzxl86wiFqsM4F8hyQThs+VK3wy3QFmbm7AHMumMP69hnLfXo/O+fWE3EuP
hnU5Nt6wrVyc0+gLAPnui0ngG+kL4D3go8UyEBj6etwp4/5lWndEQrpg702Ow9Eq
mYd/xZyw2jAgGp3I0TOG9s7EMS8tEHcJAkmz4YCyTWAS+oBu+WlJRuuYeSF7lik8
PLD6DW4ix5XhqoC5kKlFClZegN/eSb7NWbDieEhBu3wTzd+ieNv8A58b0l7rJwAL
EUUckSshm/FZS2Y/W+h3LSV0QLD3mBeHiOGk3AMj6An7HNjRDgAZetrByB31VNCy
vIYpP/V4WSGRFUeCoXKsjyey62sOjh4vRaKkAX/vW9cHwkTxBZEahN7A1k1k+g3Q
ekLtuswz4ZSNI3pIa0TAbuZ5PFjy0i45cgsIyU9/kfu6zc2oSs5DN2rVtBfsLmt0
vilAaylH72IQb2K9tHKIlcMpWFSbx++oiWyM9QVXWCpm5fHS73nCmoTovFzr3+Ps
9/oS6IWiB/N3Lq4fMg0M6kIM1RJnab8a/rSZJV8zmZa3zD2s9w7icz9bNKiNjWV4
ffXcg/t3TiSFEztlOm8AlPlQf7sxcbIushDlzHhpIErbZVYbQ2fy1TjUxCsdYGWG
y19CQGFZoTMu/eZabZcXgeP4Iwjr5SXRhMbt5lYn5W+oIrLKAqIqvCIYV/iibQ6k
zEuvQWaj0VWj2CzEKjSr4AYcyIMxAJCgqs0i8+YlG2sRtgmaDcy0AFV1ty2HwaQk
LuPBjIlyUQ5WKFdAJYBshD7gW9LSRhW57m8aQsV5s9t77Bky0d7MtCiZVPnrUQ6y
6/W24hXqfdmy1it5Gbh9yPCJNp+a0s/XeiEV5VN1tQasR2R9yPiC9pp9Mjfft+Zb
xr9Q+jDCTatH8jP63Msg+wTF+ELKzYhy0dY8obOwUPWEjGvMMEgHB2+i6TRmpSvw
yoR9qL2znrSk/LpZkbQOHtYJZimNBBlyhu6pzqVrTLjHhZn6ZPBcfczgITDyXT4Y
YyaoNYrd4quxBEq/GVP3CwyH4226j9Rvi64j2xSWiNlg070iedTQ2lbgE1ak0MPa
Zjmu4Y3YNjAVviYqOo68WQx73Og1u2BU+iTf0SPsx5U1/yRKeje2OztL5+2py5tB
Q1PX+HXmNhk+ZEMNxGHeOXJ0LzrTYrvIP6SGJAr/EArNa6OOaVgRfNz65WfOoSR4
i0gAnfuv6Vxjg+gkvsyInVyQPVJHdPSKUOeup4LyfFN405hmU5r52s6k+2d+pozj
7HzvENJMOYBv0EUZ33PRmWmpE1KLcaaKwBa27KAkKgx6fP5htz5FDEszo3JhVGBj
WEiK8dUL5pCZz9gehJcmFuvCkQ/diCGk/JFGJyndfqhtNLGKyl7YNvFks1lucqPj
evNJrs36WSNPULslciyAQs+0hvWMVD6oqZv7XbEN5Xk3mqlelA5XqPDr3glaCLbP
kFIvTHm+JitFVHidx6P9+Dbz9HG+REDiA9wAyO3yNmbnoNG8Yxnd7pElOLDIBg3S
T3Q+NaEN1/43lTpbRN8ciY3XHydBYapSUGPVsvE8ybnLMxG2ijxF1UerQ5Raz6xo
+5tyGzCnQk+b/F1NKxhP7+hGlsXhyMW/T44JoWE5f+Au0PrME3dHXsicRT0X5JHe
qePk9FEiCstKsPkac04oB8hlM5uQCiHUlIyqqTLrEfx6eMGYsRN/CXz+bqgjAcBB
9YryYHcLRAoSqLWuHuQS6bHhsgepTBJBxyzvqWd+FH7eQgeXyEV7IVBK5VdRt3KJ
a9WZiPIhjCvqfgybQFBkSk77zOGRgQ/uH7ipVR5RWoz67r11fKV20EnopmKmVjTz
/4jHnj60LbLd1gfPgTQesxwnFNuOhdMFJqGwUIy+bqs9p8y0o0nYAwX5VwTgWCLN
D8KPeor8Go17bF+FWvdun1PJ4yAEWcy+Z6gfNXL0bB2HxNIJ/e7GW/26y2MBMLhl
uLQV8WDca6yDLGk5hPtZjxmZ0CFIXwytkECSmc9DXF8KMsfrX7VvCf12JJE1E5ds
BVtzEW5MlTj5pq3Nze3I+afasPZck8fuUdJTKg8yf5mlxd0wYDpnOYavHR0tJtzd
6myWPCP7CgBguzwAzjQIR5ZmXDFjJior/9BnuTkAYt1mpnszcf5G+3xxuDPSr67s
Z9kZSmL0cUWfz3Ay/dteJXJHy9zYOErSSumg85iYs8FvwZ2a/slrgY+rav4PCbgB
8664tM4AlgEmE/NqyIxPmVCw751h2rPIiSguZ7bkro75mBhTRCFwJHqq9CdBHTBf
ICHnqjnClizYAQZGPJWKdwEEUJBFFZdmNapJVqmkeTBRdVpoAjlho66+Dz9+wOKE
Beu6GVVdofamlbgRHv1H+yORd7JBT7eCpQPmSApuzlcRqVlh+kQb2DGR5ZnwR576
qpb38UJmbSdZUWuwROLptHg/H8NYyUIawmmHegKwJTfqVXfQdCwnWXILjLM1HHG9
tHUxXmm/K3mpMcMIs3xbGxZ5lNb3rbG63dCVrP1rQGbse4+nO4j/FbZDqEbFLvf5
vowgPOEZaGqS8oUAuoyp44TDVeE7afPiG/NUY1BVp/jJG6iIGASzXK55b0vrXeZI
W6cSFVPuE9C5lluhqzqzC19ifE2iVXxG1QmoOYt5k0MLGwVpBlFHuJrKLILCTVP4
ylw6fUubjhbOaZCOxnajGcF11TUtWU2Gh37OkafMiPSGrhGnG57zbnbwkDyKegDl
iW1AIRkqq/yPdAQa2wsroZyTYEKe2SqSuoYD49D6QwrH9gdGYWaUv2pgOYHOHtWk
S5X3Snwpf2vO6LMYMpUYLDfOrFPatwpmD4lMbrUp5g30DaNW042sP47JNFDvSs9c
Q7D+3yUm1dg+i2XdW+arWdFvhsgUw1iKZPEdCyI7CEnyUWRC6XJY28RoLuqoz2QK
mgcBkn2OwplhV4U/6d9pY40/tRt0Zp8zBZmbTOzx04nug7pIHMaM3zNZSqDpYdWx
eJO3SauwFYOPlbYPAfs9F9eHITAUGCJDrF+55p41EEXaL/+GlRkGShYrdFOpMZG2
gpIMtix+DiLPkyefyBVbD0VoUYtICMRC23uGHWVFxnakYUy/2kALtW5MqcWD9/fS
0cMffCbvR5ybUca/KanF/8OQxS2DOxEBD5+uA5KFIyEmnN9J8ejibt2tmDdPzzEw
wUN1x5OGNkjPThgpagwFdHHPXQ9Sn38i4jZ1f4bxDa62MBWSsWhxTw3ddBCkOZnE
bjOJ/xdaEben9vO9BQMQwVG8ot7OMoIVs9g78UESCuyqVwT+tv8OPdGfxrIrWehk
0MOThFz52QgKjIfDdkzgh6yaGrajOrvTTERm7h0DgoHclqS3+++ZejZUhlt5cKxD
zGDdnAVOoCKv2NwRRJ280P6B9dA3J9uv6fx/JmAMmXjbu3nO+mWzvz2VNJxT5sQK
g56bcSKCaxud8tWJOLWKruTLBBOp7EjOVhgwbELcVwG5H7i5tN59k8uRibefmKMJ
XuRmJto796T69jNbUez1TuWZX8iKmFSoewnvpxhKLQY8m+N+0RjNXuRYn4f0auwL
vxodE0g41E1OQgYHhpGX5PakswtPrVoR2AQ1GjTB/Ugv/LP30GbklT489OYg8imO
EjfAg/8WpmQIjh0DjEin9uHXdam9JwPUIqC69XeekOETe1DXoVBp5zjuDHDjtJ5T
j0i62kisQLB2VGVz+FIOiJZiURq7/Xs1PNpaa/KHB1T/wUorFg2QYYCuZVKsIEZE
FnnsxWxXEo1hMip43abdiwYFGnv7avT87TDtChCcGDxYkFmlme4hEEkJFuQlS6tg
c4WqOEZ1CfbMVnlgv5yX32j5q5JWTROUhyEThtSanqsQ41kzCkFE5K1kLrVHYEBb
nuLz1GblMNpOedpzGiTRMtv3JCOHARyEgvP4yHZgXRvTu+/fxxy0Nx61rPcBCLkc
SN3pqxM9Gu4QA26ZMtJiws/cBxmaF9GJ2RKDSoByOcK7d3wu0yyhlww7ADOT9I0Z
raNYqei7QVkiAjhfVq69XsWOLQEMYGKvakKoblwsdGQPTWgSXQM//u4WTiGzzaif
ASHp3n1zpOHKmP/Hcxc1JFOYkAEBbKLJImEaSOi94HdBzxWZtbqnwPVjBaxzLSUF
zSSxCZmU5NbfhF9E+/K3SXZcYNl948jhMxKiyJVA2y5RRfObFhTCENTjrY0tlWfA
47o9Ii6ucdaezBHMZeE66OE7nWddli2pnEjFefHvj1BGK3vV1Qf9zI5s1bDlLl6w
c1fTe3oKOhu3GG7QnCWJ53HvLb8pqqXFFt+6L9bVfQY9G7Y2bXTpViwokABa8C4F
NVCLeTHiaK+joUQtCZorbtw1RoFUBXLCTUmwM+c4awUpr6vc5heOIkHgYls8cxp9
gtl6AtdA0pRouWuB4LLgb2kdQWqzNDnsZSvk/QTNSHc2zChFyt4h+c2MeXMROtb3
Vsd3PCLjRRVYctcNI4j4gG42zlyaAjMmsA9dXHlvtyt6Lj8uk5buLS99x5KzyL+D
10sRXzfPIAMuqvzjR5rhWQyh6bnrIRWmIKOblxANrMvQ2OrBt+oI0+hMrd/8Q2Zl
QHk92cFb9PVP6xRuYqyOhvz7aqL6hspbBark8p4bBP/XjRT03oPHPLUvzmvSQpL8
Pko9ZXDTTKWtL9GrLLBSFsOUvb9ZW0hvs63d9Pq/JiYwWHWGe4cOgyePijMaJJgP
i0BaQdBTlIucNZ86660qb0epjTgq4b+pWfozy3SkWWosTZm/dVSATNVb4nHOtfIj
46iLE+LHt4RZbtxI/vmrtMvzmAihkx42YfKdO/TO9yW+RLJTA7i4re19L60IEeNg
BkvNFN84Iw7KsjoiLBviAYsCd/KfRfjvNI4fnKV3pvl6AiigxEZx475yKx4wcCTS
SWmytSKTK6DnaPunClr9AHmPWnVEI8SYOgygARiMkf9vsSNWC/S/K51KWZpXG7MZ
aN4gplmrxVzYUOfuxfSnVNJSkopG+2uwaGIOk3UVpwmQpMq9MKyxcU/p38sBRYSP
zVukHrZlCvfq9uQ0UUA/PNMbMBJlvKy1f4Mw49YjgoJuIX3Qv30joi3i+ocXHAVA
0Ja/C9GwRyhhgt7pMjfMZf3NBMe/JMdGuzWDEzDf5LJ92oLjre+NFbKZC0T9db+z
R6xtnHV95Eb7pZWR3E8pkHVSErD+5ix2yYO5zc8FOf9uqoejIffFoadlLVq56hdA
iZqahoGGc29y9BX6H2yeKogC1OMlGxWh7Mksiwp3reSs04h4qBbSw07Eq6i2XJud
UiXeT8eeX+7VaRCaIc6MgSTs8kYNHb8U4kt9SPbTxKNlQAeGBwbpUGkeIkes1/hk
djDgf3wfWi8Xju+q7NxcBv/rkLLzofWxIsX8xZzT8gmi8wxH3WaTjU8e5Fy2blK+
3dkpvzGCtToffVHwgVvmipUT+o7SisYN2e+PSeyVz9rburED3qKCtOujYmIZsYcg
DMAV55eUD2vYqkOM5G9CoWWq0gxgaEjepDbLSvdfCfWsjqjhwPbvlN0v58AwbpxG
C8YqsBTdHz27JG3OBWUpE293cGILRCoyWjahlMqQusQ=
`protect END_PROTECTED
