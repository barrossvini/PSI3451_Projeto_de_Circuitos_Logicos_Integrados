`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mf3uLdxD5Iw45vHdnZeAQ9Izha9BgXtxnqFbdsCXXDGg8/Oa50Wg8DYwBXMjXARY
brY9thLnFZmhd03F5lat0IR2eb32+6GzyGR/zpNNCjU0+MwEr668kthdddtXr+bY
pQFpl/kTpdWIl2oaIzgeUddURbj1Qg/96EAPGA+8D/S9k1rNQl1ylo2xhAVEplA1
UOQFKOCSy2Gf+1dYsZWSmySCO+Lm4WIyr8xQwQVEaVfSzdkCl/WdyTmuq6JpJ6lS
AhBFggnqE0Pzeuxqtnsp7C9AlZYuHDbpbfINDtZ4aVCvjnNLDIbUQfP4Gw98P7VN
zDQmhMnSSUtcopyi2CEJXUIIUDPcz2Y8blqRqwYxnvv0uKJFzJDa0irdtfwlKm5K
CYTgxtoVl4yf67BQZsqQKMfKMwJ6kFEQINEESL5gxxQJmpUCELDjeDdbEzfq+jLt
TIJKO2Opk28bkmNpemEnMZfkq/d4Tg9mteyXxfzXKbRKvOCTwC0C0OMjtkHvPbvk
0RzUtdqczW9mprCCpJJT/3k6TEMOwgvg0kVWM3c5jFkJxE67oG7o8XHktKLCW/Hf
IbNZ77OoPd5qmnLBCCUuEeEfUpBxpaYL3yhkgDg9xPxVZIOFNIwa9gTOds5iTSRs
w7Cz9YdP9cO1sirOFcU1Poov3/WkKwRrTalvebCn0rqmlB7mVJ4YtxIhDafNnu9Q
RS8KPpp6G/vTWzqj0tyUJWld+LnOEYduR+vd/eWhYFk=
`protect END_PROTECTED
