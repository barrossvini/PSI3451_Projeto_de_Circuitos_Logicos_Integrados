`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y375nSkeO89ppAJ/ReqSNj0yn/xL2aAI+j2d+H6bxSZFjWlj4oOAUxDeT4FeFCC7
6Pdb4VypaqH04CxxTSJpE8OUMQyQV6EUd/JCbT7wE6YVma06CNP9+xF0BDRrHEBY
JHXMtFFd9qVdCvYXQlZxMkwu0coyLPM1UZnPe6qyZeKnZ7Q9lMrX9TYVnyDmcJd+
qbty3Q4P8zmL5vdlsLzH1bYBf+kgxFr6ApQ45GE+QaL+cU5e3TEwuTjY5UZJbUrI
bkJrUirpv4bqcjMYRswH8plb6v5PjRgFFoWFK4TQ5jvy+B4H/AIKFesb9ij9UpA2
RPuM3UppWWxNrxkIP9D3D6OZFcY2WbPVs3Lwh5zl8kXpkXFazOvRcngN2aVteOjT
/HF3CsVvqdHztpYjL8v41B13rNLMuU6YvmrwNETAnSskuy3TsZxllR1sYTNujfG+
CWZNUY7qggaypm77+0Z4DOe4XoB4teT/L2rbHBLb1BJIXtO9WWqteffhv90cssCZ
/zQjc3dNU9zAXy41YRaoc957IHaoV0F/JP2uWvtOHy5XZ/rPTgFakuK6ADoZggoq
F/JMmXpS+ZNM27HxhpmQSuJpdyr2IhRLYEwYajcynKg4pH6XP5EegVJkpd58CXgZ
kfWJ4kK+GAB4/Gkshso1+foRjK58tjHV0I6pCDLsjR1ZTI/zkANVrW6NmNxWTabj
sxngBknSMXnWswrpvF5zYtBiBrsAjGppmK0UfW7T7j6YmOU6g0HZZyO80XJUEg8w
BJXn3ZqJ6F6RrGVA9UT3Pg==
`protect END_PROTECTED
