`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xg9gSlT/gEgaBNuUqGXh4CEmNI4zDzTQxgpcuCy1cKNL5HDeeulN7hgW3xRVJNLV
za6IU223jNyy7kEefwcoDAcbRK3gwUkG2lVhCACAeOIowr7A9oqLiKLfOhXRSXtw
hxCU2NKZ7jl3s+H7vlM2baV1qixxXn1WTIBpK6tPVZSFba4yxMdbM6DsFH9ITjBD
ST48tvjgJgUXadTwBjI231Dz2Gj0t7AxFu7OlCO69ABd6X3h7YB5V5ZeMentCAfE
CU823NMZ4MTdPlJqRb51+9jgoLAh7S2pFoDXaXNMBvW/nrhUEwta3EWpbXQiTyAB
MzsxZYYk+QGROau/mM8CWZR+oQNLODW2QoVwhpeHJi/NE8HG+bXDuu+Yfm7iOiGw
dg1aeTiPdLxBFPbqoTAEsN0wquQH2kCIHR/hCR6EudVWyysw+wLBidEf4kWe/IRp
w9mFwr5K3fEQwL2ONzeQwb8TwXGeo0YRItPK+wqoN88ddlAOXp0PkSMQQp0Z2mFT
qJWEK0TvzAf3mBYDpINuAzDOG416lqDVAgfzzLV9+Uh31teHuu6GmQMBL/JBkikP
yjv852RF6Jswhe5poLDC7q71eV3ovldWe9C0qkILb4XMeBk9UV9nrMeze9bujbuw
oScuzKMiiQHSrI1V4/Cr/07YOzyeNW+/XAPI0awZRO6sJAj29I/w8mvOoM/fI7ik
YOGt47IQjxlkhc1wC0hm3CyUyy53qynMt+dd46FVSGQ=
`protect END_PROTECTED
