`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t99kxexPN5FLRC3CBJhBt5S3ZYBM1wijym4doh+q0TKHmaLLmgeg9PzFVxxBPpbc
01/eLblTzj3zElhi7aDWbnDZh6e4fnubXAedgYte/O9L0oZgXpNbQViEYnSFwqL5
LyvmD9yygA4LABGLikZQxXJEfYq9sJdjYwGmWDkbpqtHPxSmnf15xTzzf+6rLgJW
LZS5Rwjsd1tyd1ZhTuXuQMjOK94cECeCzuuxVEgR6c5W17j3u2QfrWJut4knCoAL
QGEKg1VIgOtNPiG7cuAPXQ3Suo3gfW1fTcMusT/xl//HknSaP6B1z0CZswmMYIKf
UMkdyAODdXisMnarXdY72eIZ7qB4dCS+1J+GGbR91ESfUn+b2do1HHm4vOgKxgTp
09DfWjjWf8zKXoKIukNZEjNeU8dRYSzPpfYUzqgpLNAuasm5C8GpiTN98+h+JSVf
iCmt+E0xXb+Cj+D7uAiLrxHIqAjl4+ltLu0am6p2ePfj+a7Mg/xScYuBrlXlyQN2
UBQb8ZNkOkblgxagH53ahNhixD/17X/+fRouK/BG6ppFAuDhqbuNczV5rea9SV3f
/ea/DmA6jnUCyTkGVEilLfmhyRvl21z1QUqjhHiqq18kfofuqrQOWi4kdo0ZoFhi
VL6b/QJuwrf9aqZ0dkvavmJCWs76HcJE1Wxdl9u+JFf0JcPAZgcLjTdwjkljFJEh
SzAyjWe/p9N1QGhJLoTM0STqsaDMuaKuOcUYqJqsNnpx3kpmuNXztKFeBUDQ/P0G
m4OQl1Cb2VKeUv0vIUvkUjdufulgFsfPV2VXUb/pG8qgFO/MbBWkVY5zptknZ2iu
nYlXQfQPVnTLMO+GfXbTfeWQ/sQTYLwyOAgVCboKoHj3j+hyppcaWALfnqsMi315
Wmjjc53Q6GjPqOP2fskAcgG+Z7UcZNZZQrEksvRz7oQzqD0wgGk7YhuEg4mGm1v/
qm70QNe8iR3FYghdhJFvXITFfVO6KZG1mTSm46Zzap1ZZOCjfM5IRgNjheiI0LMQ
qV1h+HTdqEbpAbliLcX5anJPE1TdJO8ou5c8xTbzoKC7CkFaOiD/SbQJBf/+/AwU
kn5qssghKf6GhFRrAEFGrIM04KZIISThGMTtgHBDgcauymlWNF6MHPtDbvQDGZx1
lGeqyG7Ew4Mnra3lNLjBK6nSCcsfEkOIb8w/SJP0M2n5zbrMy4aOd5BxB6vpWEhf
p2FSJV9WHPw74OVCYc29QAm5ZVGFvXFSuMso7M+6zaMxLe82fpLGdL6LtVSCfIUx
RQjE7mhtuHYJgmpncwuw0I5L1yRSPOxd7GJ5EjvfRb1FJNmV+UDQBQIwmEh6z5ts
GWgvG8K2TKekwTUnGa0Yv7GXCUCJWacxPI2ugnNaIGN+W+jboinC9zVJNVMxXu4S
R/13S4LpqAxsoJ6d9W+tWZn1GkZqrAmS9NSOdNP8oEq7y51McSPE9s47BLFgxt0M
vBUEzI5lYQx9FZFJifJorpzNjipFOPipQ6bcCNR7AWeP4jzakXVq5bf2AZRvs6eU
uug21Tog+20XINHif9Q53YR2O60qIhBGenIaLodJ8uYtVT5u5EeRofpT3EC3HykA
sfJOAq1bQZbjSckISbIIfqDof6NVQkFQdx3EK8xzhZz9p6XUCu8q14X+OIbQ2cSU
WQEwXXSpCLTJG0O8HJ8xmLaR+7YbUbiOGFEtrlcpOtgVfdH8s9MRNuGjMRN6oYnj
mTqKqXBBottlVYiGCQRXagOBP/9HBGznNL6UmExOX8b83JHNOsKj+gQ2BNYATwfb
iRZDk02h7IHwk7faiwZY+AR43+FnN5IHQd7PB70bLno3jIX5kzmQ+HI+eMuL1z9/
w72LZzAbYPNRBaLon2JsP2/sLXkBLheoQ8LNTOnGiQcgu7f+ZQ5sC3AptbJE8M4s
NsaHz5/ilYlltOO27Y14HECHKnRn9XC+yfN1XuYd7CsQKmBgZrQV4Mq75qowbwnd
CibHwhu9hi0/dYOvtMNP87fwLd8wS16fJ0e3xL5n15JB8/m51jbXs9x7gdDNzODl
poO7m9kedofTwAapVuY39u52clQA8ZMOYNbmfTp7gAzYJj/TPnRCQhdabdyoemFw
8mHqMSJLxhcE4trFZaz8/kr/XZuedS8mtK5AlBXeDQBdg72Be3e0XDjRTlPdKb91
lGNSDmmOHyL74wp/ez/QjbxmlQOb/Gvx4S/VsANSRS6mXr5ydenZQ2G75/EsaSHB
OR/f4HQVttkKKqTResHFIXi92r4WCUFmPAlmnImvcuoqOe7X48V2+Rw7jLuIu63i
qX/+WW1dfwrrM9BD9ix0PKHj95GIHukCkJvJMKEpNCwuxBOVinKfLQZpmxxrWnAc
R5QttP4UlZVlctV7JCY1DlFr5/FWrZerzx8duibf8AGNvYUYuMEGEqQ6IX80uYIN
LrJp8xAg8VW4CoDL5FRtTlUK04bwbVUlholJ+ijJkmUcwKdyEU7/y2GpMn562p0+
tznyWqevijL4/VYZ1L3ZE2QyRdxvyKNkQOsGey8P6tt8s7Zu+0xFh5Lla5YwgMZY
SqVdWCjIQSYhL/H5JRlN2rP9IZzX+AsquABws/tvVbuCShHA4bcy6bdn6/HbodLa
R8Ze+r6oV0sYGAHBM1rd+5LKrq3sXq00P3NGDd2ceCM/AlY6gnPmtJfl7gVx8cjb
MzJMhCBwPzBdG+SCCY36AYjREYXUHrTgF1b7A6imquWdCSPPzngH6xKZv8tWyzNu
f7GY/eE7pQ0tvCAXH6Yc9ZfKnRN/cAEXwTefaP5jJf0D7nAIiPxCWTXtq+Wul8Hh
T4wtPGP+c9ezUxAiXrto2n2rCeDI2hrF6uSXUisY35/08J/CfavjdhwAPuj6rS//
q4HAf20D6+i3nB5Szpvvxv3KsDbCNHjkgBItjMMaHKunSdRU/GdQFgXo5eRu79x0
H6glkdmhQskhEa7PvGeDZ4k7buxI2Tbu0lbXIM8kT0Z2CjU7Qh/APhmN/g9f+B+F
jTtIfPx5aWGF1SSB2DGgyzquyxWHLzlQU0CsPemdpi0dArsBd9kSJBolXhCqb+eK
CIxY8x8yluLW3EWu0Dy6g3ufVda2aq8W25gi/+BxttqlqDevsMdExE/mjccncoFO
U1JGKj6o2zviru5xqZ5828jXLnW03XLd+zz51Xo8dmZe7nGHepS/SRF4yg/Ldl1j
uD5p9Ar9YeSzo7GxHMTjaTmUrzdNqEi3T3baDfwOEiXmcdM9clhXgPbI4DY/w6UF
r11IskcS1Kx+y2nrFqJBismjGvd1RLgN9YrIXhZoa7q0TNrfDk3HzP6V451PTrpN
PuhoqGj2/sA7a4YgMAmobjx0WATY7J75VKdAxuCjz2nZvDpPx3ud7MDXwGmm1od8
K0yE11hXt28ZLvNj4VQLkkkSDkInj5zzgWAPcByEFmZb3+SETzG96aUU0Xihpu9A
nKuD4ZlRlrFbQ3QXqcvxFSrJeSEqCsxedxrUstyy3lrvzP+n8lhmfQIq1CKR1mvW
swZ+lG5zqeQ9/fphqrOnyoc6qZ4BvOXTSNKF2J67UAazpkzYjd4xUzDGMtSVXyL5
e6ILYr3gT82ulycZpJpIPVksOxp09cXSs+RWx0zSsI3mw7emxnBNCnZ01Mt2cozp
n9eD9Q4GppJCX5mwl3/bbc6F/JNqwdx8vtqssqGBJDmruBG5FASxMuDpFPMZCLJF
eQwZO7I1Z0vgx5GqdS8kzCafcLTiivoMYhogX0NHVLV9pwxkozPrIrf0vNqh7noY
sgIGTpZRCHSpJZJ6BREUqWYc0AlLXQp/gIyYyHnWECs5M1fhSXrHeLXPK38cQpQg
M5ym4QLPU9UYOc/E4r25PUPaPDMIYQAFji0snGtac8CUr7AwD2A0OQ5EnszoZy/n
wjCGebe3u1hz+0zJwabA4BBdQnLPr+1rVd3o545bfBr3CkKDWUEdwE9CQxEvefJY
fxMz2q3F/lnYUazplTnY82KBIXthG/2fOxnW4uJYtLrVHKeDKUaBL5CGcleemUSV
aLhkbr95IG7fkhSoY/BXEioFUdScDwxxvw5amfmwwHwI15BQLkUreuN9bn9x5USg
8QC2frt5/O1iO2wvjX2xwQMwc9b5/27bB43Bfmif2zrAR/nuZMA36Ga6wof8PxpT
lLtrSR8hMuSqvfq4kd9D7KNYA7qZBRV9V0dIuA0uhj0NxKNCGYv1TUVLtND9ptUg
RgdBSyiSZyHCGCzOkzbmFCARNNwZvGhUNUdoGdr4XiFyYUZTOE+gG4NZo4GyQztO
Hh2doX5546BvJtuSceDOaOCbyPcyH1lg1x7anmnnZ4rNDOrsa6wnNAJ/dJ1y+WCZ
90RQKhK9vN0/3603rYlo63PJ/jBT8hYB/UX9cocLNrq9AX61ZvXyovPvKkD7fglp
vZIMrVttF83AcmC+NEwfYrChJIjDOZijh++fn0D0Un/vxI/t8E4vWcut/UIeyxIi
Mc54cAP4HtvHDB78snYYAuAPS081ol/01q+bt5QT10uoUqaww6AuuKpAcglEStgj
mBLbo8YyE6GItjnQXZbrp77CVrdYs2piP5Ej/W1cH+5228Z1ObESuGPc63bS+wz1
PwY3wp/fIE+H1t/u6YjXq2UqxYiujFi1ZGZxnE4rgERxuVooExk1TBJ93rqB7nxb
Q6ScK/Y1WFjWuFs7cS+5OJGsAfThF53UHMVBkahbISgGNthMyJqRf5sULt6mPn0b
C5UhuTSRlufBvmZ0JTon7pOT01iegVr4VP9G7oiFFRs0j6yAOl9KWMoGNKYZjosU
+EyvmfQr3y+M3ZmqLiuhYqUm6jlxFdZxTOHmfWRcU0cJE4o+FfV1rnCvOrI46a5m
sbdWAeOm9eEMbZNlDudfw7+1dZy5dtQSyeRzNiSnZM20V7dfUzOu882I73UatHru
zk8SpL65GHZozwaGwKw2MMspCFzRKw+HlqY/b0lPyA/s7QAOC47Gn+B8JJfmNbHT
ZjR+qrX/CL/QdbC2ShHLFzJv2dksT/0J2kIh+Zh59m/xHcOC8ibxbUWFwweiMg8l
ehnkmMD7SbMI2rDdjxEF0AvErCUdS8cmrhNyfk+5EO1t4d0u/oFu2IA/HM3xUksG
OGbhGLek1IUSaYBi44xCNPzRz+0YvO3tvM+tt7hhpmhYww/siUmgqU1/3MYYEaF5
SNcfxwMaujjbn3caoredW9DrRE4PeerSiaOtAEU2B1fOHkoEqwszI4qSUXtdwMTI
XbfzoyxTym6lMlBmdw8xK+lfkOe6j4VDVaXh5ZsKBlQs26RRYdDNLnbHxTQVHR9j
VC4/RmNuzHdlgaLumy2IQdD8Nq8thq1YsPci10/wL3I6xfOBbD2Vc8hNMsvQSa7J
qkD5Xuc4KZoeGwxMtAvN36A+/QoizyIC6YGK2l9Sd7RCZy9lP78cJ0fjFN9ZZhKa
vK91keHpVKOffGAjITmiVCAoYCq9HgWLmCGFI9Tc+gYSrvRGqFRrK5svkrm8C2LC
ZM7PKX5yiuiTuBFPhFkXxQ4JxhadIA0GeTMQJbpFU2nFXV+vkoT0nfQo/8KvHzyS
jgb11xwLDILojNMdtU2ZO4du6UnO/5bWlkSArkqCNR3HdNB/g0t+BNfYas27alP6
rD8xu52Lqs6xkp+nzR8k/gPSi7b0H3NvwmXlQncQoc1qxzfSVlt9B1ZnCCIMSZtE
pF+v5NQj8qqRAfUy5/I7v7GmEAMZh6FQY29GEgyjLyJ/9nq1t+TMgpmYrwEeAOGL
Drqig8atSba3M+5ICfv3zbmxIidP8+a9X5M1iP/Jam3uKDumscPxNJNm1xTnW8o6
k7geA0PTxziUGbmTBzugFx1BBgBcA3tGxsGBb0lTPvCIeTs273WkzqJm6sYoPL1O
CUbhGOVhjRFZEkj8KPji3i+0lYQ1UfQlm3VwhZq4Ur+pe2oo0Iatzq92VLc6qV2o
GDYuI8Hq/0hI56NeCik90Ebinr+HndMFFEZY5F4aQOz6Uct06IXmGGd7Q/ddzb/z
Mob21yvPlhSLOmBVuVfmy8fUI7kEOwQXQG/hjHLuxZ5ZvlYU3QWHpb+5iCF5da9P
gaNbZSHJHYKb6mAq/zqyz62+GHyr2sNJjsenh87doFS2tSoCQLgYsyYNLpkwZcsS
DSVrDx3JQ4MV0gqTWvUfnPCT9fYQdcLUGti1GNSpDQ+KCPIC/x0UPhEeK0JJKoXU
ZrfPLKrY8rY71cLYryQn6vkPSC8jWj7tVMAg8GKPJ2GAH/6pU6z75J/BoNT2+KId
uebi3xzFK+r036xLl4/EgzdEUa042oBOk9chtMJb646EjaMM7aNd94lGA7mi/Nhe
SfxnqPwkarZLmczoT+cw3RFoT7pwU0BbKTHn8D81rBhOHbalFNU9jyu5QaXu8ieD
dh0Xf/Ly54yYwGSPg1mScgPj+fHsZWIUu1tVOIwjtKHHs5poQY0MNp2SCJiksuRI
KM6tSQooCryjolPdiKdam960034i2pfZ2xlld0KYqQP8c0DRWdRPdlZ9S3dee5Dq
xTysyqtRio0FPvNklSxDvG7yw6sd1LCbZyzWQeGZHVOIBEjDtyLUD5FDcLK1MuBx
nc9a3j/yTs813Zz/3QrSEFEM5MEdoz1uomHUc1iJi8oTGD9g5WnKQX7jOUaVoANQ
8MYMKjxvWGZRQyHayM7aDaEQcf3n8lRMG2y9hrWNgWF0GB9ES/Rf5Kn1GodqxwBn
qpseNbtiSzFCQwYNULBChqwXuu71fHFnGGD3v4iHnn1171Xysy3NqKEOmprMpuXD
mPzCrQNRNYU/gGNF0FJ/b6UjDrNudmziJgWnLwU/dgigAe13JlLSflMxX3dyrys8
gfqobd0Cl5Mt9cXF2nnFDLxygxVmPmcYIL8j3gpM0WqXh4R1wTZUVYuFDi2wqamJ
Vm1dnTLUZUyZeQ2nbwuzCdaDbVGyTBE8MMY24BFS8AA0pQju4VwcePjtUsBFQtRq
G7hcAUl7OyIA6MsRg+EZdd2qQbqFGgyM/pFNWkfiEP5maEhVizx0NZFucgbau0W+
arEGrcQZ2peML4/39WclsC/+7GzdIQGGHRNP5vrwRbETu6WvlwvDT37FeLzJcGzf
DN93I5MovUAawZMUwmXbGoLax1m9EqesNWVkKItXIJKZ5qqLERNgzORclYeFQTeJ
j9XriQthKih1H/OQ7mptIXJ/aqb7Lb0SnANLk5je0Lc2Bi2cqwap05wv9jE94xWw
6u7VLdF3xD4LFnnTSmpcSYcaLlbCLMUhfWWgv1Pj/1tACkAci5+zAg5UUL88EhEz
tCTsB4l8Krihniwiv7EUIxWLDh2qcfTyO9RiV7Q6pyvtAa9g/Vieq6CKMHp578xd
pGqkbWz/0rFcmQ6izxBQxb6YV53IClzuTTQrU2zPbIENQB1H2tmLkQYXDQvX2q3v
EobKT4qvqN26SRypxKVxnAkDqaBJxWSF6wpb4ceZA/hAW0990bg397KOYVBgTQ/M
wiTAjIUeZaMPnwDnsL2z8oh9z2QR+oUkCLVqFI/qV95ztXTcDAf1HYzU6/jB/KQV
+Dusrt6yvPhsZ96MV0i86+kS/TA+p8j2aL5T1Mf56tGkgY7ZtBTogCnCl9j0BQNd
TOCAs6nVPLPM/tho3ojOjPX30g8JT6IyXng7T5j5//W4a1YIqysExw0EfMnAD21q
zwcD+5JWYhGICWkkRMtYij+bqFZW5txnj7v4O9TzUPej4OdCTfOgYTpatZiV9WYR
Le3FHIp30dA02MmtGzuO5K+2SQydiEvYae/v3+FsHZLOBev7UNjX3PPtXXxkqQ92
NI3X25mbnQfiitbU4aDVMdsVq4PLXHhpmqJfltme+0nJxPjXn+i2NdYC4AP9Oq7s
8cqMXPrCFMVqKpsBCA6TfaDGMtETdwLjoT4LFWYXjP48OsJHQ7iyUTu7SGR8kiWT
lCzli4erEdgEQ9WDeFdhxM91igXptLQJlPJgUkyofBDpKdPpsFUktH9TZHkmZ+2H
KB6IDs9tFbuyvTDlE+YAkwD1flRXZUC8TVk0YJi0r1bod9yqa1yKTnNHyb4iumc9
MHYOb8z457iOIxP7xEccrtz4Bo0EJd9P0XIzH6A0Onko9BEa1011JxqT0tt98Oe+
57YGAcU8kWgLenegHrEsHQfKazyt32+iYvsQ5Qdj8t6szqrC/fFV2hBnVHDOVOlc
3L/GOpphIO3WXZGQkDyMdXJBWYUHkU3aQ7YL1IaOXDs31ErmdsXl8BsKYaVcAu2J
WXFDOVcD4LWGygiPSjbUZHvLVAAjhnWZE7jidHcx4pudXwaAmDezwmG6s/aa5jZm
vdTKqdiNYt90JBbcuIZ6iQqQUx56Lm8cGAIlz1J4mzmxauDDjtHHJF/bl7Wb5/y3
wyfzPm9XqBoaxSSRM5DhbTkAGjP4wqu+pEsWHWOU5AdHgAVmcbYflItz9SFitIog
5jHcJn/Vo+HVJprSuPkSoj7X3gOXpluC2PCira8+LF1QBFRGhPyDsiuVJ0/yFHFT
2DySchoAXJZOYs11+5OvAGP4NbhkvXt+opq7odVFFnpXdzOb7QVsbCmp1Kdxzno5
omhAu+XTiu8xASSZCn/EuMik0uutkGxvrQD3wLkFon9F1Xo/8JSws5hTafnpJSqb
ee58DB3PefLTuWgyAX5QMbOULIJHYVyyBp1UKqbWazbRlqORaumMGmuxUrspTico
Blp3VbLzukSnWob4MN0QiJgdpd5Xz+zZupA7Pc1Z3X9+xNDgzrMc6yjqMP4sYAEZ
Sq34dl0QGEBRrBZGKgYEMGZJSKwcZYc7+kcSZhFUensmQqTQJ0G0HjO2xzu4PXBl
YOQgr+c/3JnFD6pLhcWND0CzSmg+o05FbHQPxevmkEMOc6/siKyMf1S/K5j5IHnF
7nU6rzWioz0xB7mLrOycA9NboOpFwvg3weJaD+Zy/6M2CCNSZUGxjAoIDQp0vQQZ
wh3bJtKNB/conECfqosz5iFArPwXXuPUtmFZbVj05yPJk/DFmLYXy89MMZkK3UgW
BV2PkOm0QUEodGRsZsqg2zBo6QL5rlDxHLTGLudzUSOIa03cX7KOEV70P82kj2Jw
dMxzup5u0NoPwp2+9tDWOaohvVNb66iM4ZQJXYk95ed8350s7FTPy8uwwAH4gRvk
4bcjGZIA+gzRibx7Uw5RtMkV1h3523xof5+iezojsTt37GBLpTD4UgZ4UpAABkhX
UwcwXb/5L57alunDCJCa1gTBkOhId5pEELIvSHt1klYWunfYfX2sI35BCm6YTOW1
8jWHz5D76T7pFywYYkxZVBY5gsYlqeBXFjhEEfG1HrOcJB+bM2y4MBTWPeb5sGFJ
VPG2l41ujzr3EdAxmgRep41/I/tX98ZFZytuoJCn3wZKAT7mCEZqRU6B2eMgPTRb
H5M51Lz8P9V6idHTXMGXfdsd5fwkeG3lJ78sloLQHdBtAjyP8lIGAZfuFSr+9Nuq
Fe77b5agnjP+naadpDn60GQW0i5+vIHrEPXZ6lxPOD1kxG4PQS+o4MC6iTfZ++Up
FSuNGBvKRQ5i9XvcjEB4d7Oyu49XkL/qdCTkBQ09Ked+mZiZooZfptHCVQDLUJN1
r6E8dexjQAFTRS/bpb+XmYXe7LU+qbDZGSKUFBf1JCGnKCSOIvhR3AJyICxGD7Hv
EBxQmMSkLJQucmNxTJUBkLJDXB6uPAEVr0ObpNW1/zMofO2KgO24dETrRfkgoHPV
ufUQdIrMPg6TL7w/qt+x+1QA52Q85fUlRLT01NrNcAztTxSaVaj78HaFlvSoBTuL
msHZ+LYiCMV/dfAIvwEAlIC0ZhwhNEFDHdn1jHG+uTRGMkOfPfqQyHFdFM/Drn2M
LtLZWohrgMWOlXLl2BjTPyBwq5gTccH7e3fSWMrje/ZSR/LUv29uPcbGqkwNQku+
Iavb4tZWGo+UQAJyBz2abXPT/ii/TcVQdpbeD0ZUkMIdNfUpZbtJcpVWEnLUjK1C
+M/Vp+YzWitDhpgfWoQsUmuQ4kxjY8+hEYphWYmgnrZkmgKbfz1x/82L5YOwDggL
o1wkcRTo2BpIb+IAj4ne7dRTy7Gmy6qqRNHNwhElYJHcy4ftfqTlhQqpkH2sFQYI
kfLHUCxX0vXFLTlFuSfg4VHqkeDRrsN7WvIQs8/R8yPFCpv8DacNDGNF9fVhnrxi
IIHjN+w+vZDenR6hbEV+JyniwGeUET00fAiYnhYmKmy7pC5S652+E3nneH+ZQNGR
cMRbzL/ifK1cIePXpV/IZK+EZU5sI2QxxvaBjDL7mggOjdTnjkBqxpjO4EEOxWPW
V0GDda38ZtsFqaki+lOyZrVmUub2JCPGhG1qH5eBJOZxN32INhXDWYdkQFq0r4Nb
ObtfnLFAsJjCpIhX9UnzSarXk3gYi8rW3avTnUyuRQMypX7iWCooG3d7u5v+DaBg
m/zsBgrbTf6X06C5F7VNP3ehfT9CK96l9wr5c16bHHMzz1zJmYXJbT0qp06NuGIs
VDX0K6LNG59dEoW8WOHlZO/CV+r6Z7IeL0Ro81TCblZaV1QAsrq1tGH+00+aCs3L
gHLR8p6iVJGPkuGxO4D/v8Noxt3S4eRl9uo1ngGDfZZfuifACcwIwdAKk+NO5hUD
mlOO/K0aUOrvyIs2YCYgQXWGcJkz16pck/k2WgTE8qIvzd9cGYFjuf96a7u0EkEN
mzC6ehmpliQCco6QVo+RRGmwc/Mq4MszPwu47uKKnFrn3h06cTF6hP5r3PvIIyqr
09fLEOTfmApyr/TO8D8HSOrdFr4ZvEpNz40HHHPq9DA7pP4WI/5G4h2/CUIm5x80
wtNHxv73/anLMQd7W6C0FF64YHzqQnEWvVL8K4d0W6WketyImm/sHNWSC1HuXM/O
3xL3harxuIJd6QE4jYkLNlKtnfxDoRShXATcwdoU9FGO7YLJy5kfilSTuZCONKvN
6Ke2QOSCVKuzgV/pA1JrDkl/t8RlrKdvOT6PURzV3tl9ePWRGLHjlXgP/C2Ge8d2
l/gRT+i2rp1LaVDT1Vc8U8EAMVQ6GQk28KPDfBF4jNJEVXjffwNNS8G7thvmWW+K
oA3uiWS/4K+A6YL+m8uFcsyg2r2ikJMCXxO19le0C0zltl+OtifHvJRaf7Nw2WKJ
psXu3CXF5IEPUSBAr/dp3+l+BZ1ctGM+MqxeNUSp6vwoxlTVsNs08FsliYBqsPn9
sVuJCj3HewnZOuNcLHTTJxkbv0brmbZHRhCnkC4gzJn4dwaVIhlxSBPY1ydsgzEA
hVnmZyvVP01XF8cV+xgaMsXInzT7fLoHDS6EEWhj0BPpPffqeIpbIYE2383gcL/E
YihJYOfxhrbQAD4g3jUwIUWBq5NRGerPkpLqxljmjdZbt5eNZnN8/riEZcIwnvhp
ta+fawLOGYls8DPkVA2eUaBLiq/o9a29/lVDxzIu7wTLfRSa3HgJzde4r0K9J/PB
gGAnuZDpccACYxTgyS4YOvYXJ0P+D7qkgvvjr/5Wp0AYuHkyz5QgBUi/siTcW1v1
G0F6cGAeCBUwIdeMjngpxc/hBnF8JmPTwsTZDx8vRczYRUEQWyonFHdZBHJQVYsF
23nlR2FzmRST4RJTf6G+7KxNyM7ERwmONWC6nos0sGhsSTzUp3/l8ycJ40N8JsB8
f9+ZQCQpfyFpK0Qt4rx9b7IrO+bVdb6GGRQOXKCWx2ZIquvuvrODs6vyWkT9mPtr
mL+pfw9TGd5kzsfuMpcFHETr9keAeZ58JHjuRZmGMrZQiOL1u1kVSLErJAtsIjo7
0yYwdJNzXZy1yP/enhu09w59RsieE0MhcSMGxSU0Q4QvpQlcgt+UOBue4B6VKUjH
yD/E998LhKtefSpo1U4keRABSAlXJPFxymmkj3nsRD+mkzy/gEZB0wFAh69PmeEd
flMP7laIbov1jjxlMKqvz/OmGheUfhMIbi4LX/1EQFAooTf0l43QP2OJoc7e9F95
itzgintymZ++6qDn/CcRFUG8IYbxAuiIhxZdzHpx/QBwWXGkQk+Decqw52HIIigE
O5NpvH8/UbLGzw/DbGYMMN7USjzjIOn682r9IqYqEkrIps8VUy4vO0tGulqGMuQf
HpcIaV1NckgQ/nNJ0OD2YhaQfZ9TuOvJ5F011DAEXhXmB3tZpgGEBEKhyfiG3byv
huQ/PTjb7+uBAI0vDFJ9J2d4OLVkOSPz8GRRkxDe5Z0ebiLMhgWdlGITYazDtCA7
3cXidlvfmL+ji4m/TEcEjLQ05bLAPNmoyAqiHc4PE1ZgccPFkOq1yYksC/CKxfkV
mUTl+zDOE9sc+jqt5yjmXtQ0M3skSH/lL+axKL8sKgi1k/vau6uI1QH2JkICFtyB
f0IIZQcKA+Itqu0WWjzW9wyITizw1UI4Xh3IrAFsz4R85cssUD1paKN8OmXYARvO
vZjWt7WzHwUDRS+3nQTpfi7vbU1nhLBTkFK3Q7x1GWGSYtdz5iOy4f92ErL5X9+O
UFCBSRrA/SxTRiEC+d2K0Asg8tPsVZnUVZkRzT69Xm0=
`protect END_PROTECTED
