`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
54QqFFipyM8M3CwDRrqai3hPtC6im2+63vHioVChsQKglkuwZbPG7V3Y1GeNmSyD
9ck2Fw4PGUTs/y/Fim7XkiJzQLdooSpIPzS0jmh7E8+NBT2+oXeFh7mkq0JggVCR
17sW8vEAc9Cc4Jeq64OzbcMu1jDnoSaFfu9GPZYx7At3+DqlAqD3oCkZIfo5ZO9o
S/43JIeE61p3nDxExXyv7eUw7rkTKjVgbrRqbx+vrd+x4V1hGLuaqt3BzQo9b/CW
BmdGdoroLD3kKtPIPoGLDi9PObumdHv6j2zXulU8TpJcUGDkvxXeDpd8otjkyl1l
GaVqf7B6/Hp+dGO4DulSmumjnuBnOFfwPQ5RVtG4dz1diZndy81p1ZaVPp6EyHTl
Z3/MkwybAh3p0pgONR2xx7YqxbLjDOmQmk5stkJZlA6ju2aTxa9alQSxY0/QLf/t
SmjWfpjGeTTVrpqBYuaoaLBQFnnzFYldhp+SLaxVEVYfgVa560yezs8xDPhh7Eg/
Q2h5HL4fStD0rr5z2aV5d8Ar4hxZgEg6ONQ4rZHYwZKCMAwUCfly70xomMXlMKah
ZCe3rzut+yu1rY6gSfuRhfwzAahfgWDQwgrbP2JPpAdfavn72vwAYQ2XgyTYG7pb
SU2rjLrtu+575+17B9ytQW7uWHiZ9tlM6HonJop4qM0Oc2W/tOGPX0N5+bilSrb1
Q8VWaFpmabh4bVF9zRFPMPX0kanf4c3b/blPkc2444LVAaCrMgXQ3dSj+PB6U447
2HIoYQv1uZ51B1AURGR0lUQSi/T48TtdsyHsSdjbEVWQ3loLMOy9GUlrDxPcWB3Z
nwUCWoN+YEZ9uMO4p0ByKATQ7UwrSRkeRrTtTefwewzncni8l8a+ud0ApWUvdtzD
vGjWxzjpLg1dA1IWe5Ow7PeS+H9sN5aJuBISE8r+Ka7E9sLxqomOWpW/au+VsqFr
ki8DUSc5CIYzL4F2SYT4TGPCAMbKCBsE85idPorl6EJYFVCGSTSKqWyjeO/VUE1L
kSsN+B6QZdij+YRM9UspQHnR1iKnb0KO116AY8wlAox0KpNwTWGslfCOP+s51/gc
`protect END_PROTECTED
