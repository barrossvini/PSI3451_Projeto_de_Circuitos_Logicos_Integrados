`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mYVde1yfyhFu8GBiqm+ks5GKtUzGUhckPAOGthNjvTfwhtEVBI7Mtc/5wj5YeD43
B6NOY4Bz8/sTTeZsvrvr589WOe6Qyh/5PVVYXgU+S15+RmQ2yCcZkuIdgdan2Zph
7ctu5rMyZucFx4oCdKtEUftd5N2Djy/BmzjAoIglXrYwGeib9WvyE67XP/IouZnH
5hSj9eiPnYkseQAx7Mb3JbqpcvwiNlD3/fxbYLx5LRfZCKlwWUA1CHjeiH/+o4qG
mjrMg/J/1Nai0eIK6Fih504GrzAeXOEaGnGdExY8VKqV/QQs2IBNlJ2voxvquNzg
SZgfiRgDEyDEwrl3grZ7Znvy3Uv2pYpEop17rshT4XE8XHRKEriWt7V4yBoqWEBi
5M6VKNhRc6FTIaPGJqJipdRXySga6P8iezclMUGZOMmoa7N40XfFsYZsEUZ2MX0J
H6lnMMqLCtfx/SDoxI/QEzdiNEi3SmLtBcdihTJ5XYNrWcoK5xjVa4gFo3SUWP3m
pzV75OOoFmTCRyzwOGEf2nPuhHi44OoLdvp7fNZPiCmYzBYHxPfNM71Z+1YTAl+n
p33CnXSPnrcERWNgLCDC04xzsS3tQcM3DdatKCCA/DeS/NVd3MlHKZlrBOyPKkrc
aqrCgB1728iirSXcyJTa+8JpSOp4tyIgiu+QTNeX6zMx/hNTMX1bzp72pvRkN7V9
SWCKRwNkifYwK3PmLtLwug9XnPPD4H3nfL82yxt+sk1YP3NjDiOntc2tWU3QRpIa
fhpKhbe/jLNoLfIdiSNnp+b9+7XIbJ84qAP2Bnw5m4gA8nn3lVpO6LbRkOAh2KQ7
RaJqkJ7UVUl5H6VMu/vSFFw4dyKPNbHI/eex9WQ2o4AFzc88f5euEEmK4JOEn679
baldL5yzSXo43cHPs8vsNX6wSeAXKwodkbXIREOtXku19PZBK1420EpIkic9WqzR
p0pVluMJv1h9SeMmG18oK0qLcfgX6k5efZ9Ef3irVAYwpVluUxwm1LDpllp4AXnn
mj3d2rcOGvudCxNR96W8kEzuMLTvtId8kLjN5d082kFMzrpdpywmwm1PtvDywcSv
ptuPc5u9ej71GcXQbTudhYDhNXzdCYYsF16uD1iQ6/J6/KX9s9LYWeG6uiZhOqz5
2RzcA4S0gR5u+jsNlIal/qncntliGnp2qqZ6dR1Lm+5f9zPn55vaKKAfCVfTdI4n
nSgLIHYMS/zrz/6fU5KDE7AGtaE5xvu7qeiquXZ1Ty6BKiPiWkyCinaXdiQfE75h
yR2Y8Xq62d6pQmAFBNRGDsIhGl3JuCAntxsUH1jXvq4kF0tUgg+3U2SNDpf/JnT2
qpeiSnZHXa/S8LMOI/8NLETWbXFyW4CPznsoRvBRfE3C6BtPDRCwlig5Ihk8SxAp
F4jrpka63YIR3YHHrHE5X+EiCHraY4geSoieJtgySWYKkT5v+e6WOWzfhNNgPhwl
u22J6QvnyMJ9vhFglFxxKfE9SodxEK4UeKBmFZqE/RHYKwdj8sKxMnxhgYBxNZlO
ml0Di3PXylq7+3xCJgTWILobN67P+ta1rsBFqx+5p/Wjh4+21XVDyQ9JH59lYUs6
w/P1tHQMj6EeVAcs/UJUjjuENTXfgFjt5PYWHT0tzbLrv4S5RaiPJKEUY2KRVI2i
Olo2h95rjmKU74oYNy/EMeT667Q1WS9luU2fvmyjtdD4xVv/ti2RiyQUlCIKsjmo
y7U2ty39H4FcnGervcphVwMt9TFH8jzzZszgCSCpmGA6x537OQca3m4huwmpMLg6
nK3IbHXBZY0K7J0dAavtvphxKnCOhJSxn9qkcC/A/zGWxpgPHt7VAbjRN377srOh
Iht1TSZE+Qd89TaFEJPx3jI8+dFzJKaKi2eUexPFCmVx1dFHl/5tvatFLIYbM5YC
pVEAzv0SW+O6H6p2q9RJ6tokV+KCMt9iSoYDjTDZva4HC13RgJz5kU/BG2bZQT3t
9nkKkpQ9XMeWDkC3rC0EXFJnsW0wQWw4LE7mwFnYxpGun/PxHBiPWKNNziRL82qO
oPkORlwyiTsaWsq4Z+BNNGpUMngXml/702peRgz5DvmLSd9UQx0p/yCC33DDd41b
XyaP/ncq06AyqLM0M9qdFctusBnmV/dC5DrE1i005J7SjQtb6mF4BIQT4To23itb
iKRrT+TBmejyRF17WLHdaV6bX2KOBXCyiCGhF9xyGJMveY1jvBsVJa0NNC+7RAYo
v8va40eWRYyYdTwHC7pyRKLCvopMFBUK1BYjcW7cy185fPHUOTYmWUE+PtRTGgs5
2J7jBqR09Q3nkhEzahayy924zbXQfvN6+zI4D+iI15dQR7W//wTDXcMYWNBU6HHg
Ysf+bwEJNxyvWbEhRVINV49Bwos312fEWhfhHyfyQgyvrTO3VDszp+v59OUCpg03
UCarkvn31gI9gwn8Bs+Y5gvVPjRb66lQBZTUuTIJaGwbb0gc+kBzcZcQAxPCBp0O
4gPfvWE5dpb2o5OVUWy++AqFpEBEmPav5L7C5JnaiN+8NjM2ERfSV1atZlZ7jNyT
lxu+k3kzWfN+MAPb4U6fdmVxEtOjC7nTybnvFubMI5Fbrj9AIafymwjAsI84QfRH
mfwxnKtR9Vl6hnhzkpsZW3UgWsmQ9Fa7TSBtsENj7pVX8/z4Rman+gpNcZ9j6DIC
ZNFy6jG/2yp/dnYjK5IU6JR5Y//iJn6CHDHawZaM4DVBVPEchWQ33XBsPLi+DtX2
6p+kQRROjmfsHk9kiu3sDtDfYrxE/frGnJkIr/VZadVCyWOqJRsRr8KlUsLsQYj2
Oyi2GEb/ADszcos8NRJp8AFsJkeBMSE71CEX7mhkH7PzV7wXdoiFHD76TLAQ65KH
rq7pdLMcmSmXRMOTd5smIaMCCZnunrC8AwPAY4TmnZA/9lC9FcVpLiNMm5JP3Jq7
frZJiKTG0MqmsQinRGpuQ+wOGnElHJpCa7CEq+0JsH3G3s/M0gpjpVaFgCw4gEpw
DXAse6b8ZL88dWmK5WYezDA6NtdxitSNvLChSdFWImQaQ4Wla7fE13P2xEugIE+D
BTAOaVPZoj8SFlzQ5Ns3EvDJZ2o6Z6En83g+h8Cmea3SUza8WUgygVg8gSmDeMpS
GkbeZuzF5vN7omxSg+2C90KaNDt9Y1i1wvIbtU+tMvTe5r1t+WnxewQYmsvnr5UV
2MbNOMftUomVvgjMU0Z3bfg3lExidw3FUFaWSMn4a5M5xwaVh3pJpc6r55+qfPW4
1ZjJkJcV/eNJ/AhIotRqCgXFHwACdJOTkVCSkxY/C5OUVGEzjAScXagK1ZFsqP2D
jJ0r15RTYhySJh33ulT7ixqxKo4J+tXforNz+s966bw41ENKD9Qnq8Jo7qVoK5Ki
G9UUzhqgjVzj2lRnOW57Doh0TI3FzxfpqYnfpAQwiWXFmkBCoxGT6U9S12XXZNlS
PBjYJ+406dGwyFxCFXmiZ6j26cyCpApLTvEzeXkvHqCuP67DpCPWJg5pWhkfId2j
DQILSDUY308so8fs9goEbaQEqytumiH5EvYv0a287AtWTOhcP0xMqnnbZDhzIPXv
dpDAjC8dzM7qMQDWVYcGuAr3InsDhT3jEOUR0QIqg1bFmaUszaxD7eGDcSfCJ0Ms
KMgSj/KjxclA1DXBCMwOwhP8ZH5fT/uRuFcxdY7NxH6XlPPek9BOQArfxJiy/uPC
hh9ntCk8ww3U9ZCqHdlXHwV9tfb/8qeYbr9u152d8SCtHcHwReAUekt7VdaJeyhV
jr8JXydnuwurNeXzTDQ0ZIvMwj0n4/ez3r0vOGOS1v/aBx1S3wkrKGKwsLFY/bp2
p/dD3G9QkEAsWBwRLN7shxrihVjeen+iyBszNp4Q3oUVngFaxUhf3OLqzfO6cND2
+BEgE1e42bKeqTcUaXk0CkNDHc0U1gBuIXglUDyElwSFjPDYe6JIOC4engd7byPb
FGnMUG/n4nmM7rev+zW9WA3FvCgJTmBBBO9FcQyIw7zLG8HuO8JO5k9KVg28e0q2
1VeAew8Y/4vaI87yLc0F8XfEBMDpzMJxmfxUt+emFagp2uvTUFSsTE+inK6Qxyoa
tj8xj/nqWCL7+XzCCoyPbCtpLu6grBi+1Yn8DB9zlD7sqa0axFucNAHxo3bt5KXr
I9xCcsQfGT5QbiYHO0qaxccWfj0QxckfyHQkLtz59StVbnyBqk3TqHQuoGwaySVq
izQAaDezh1fnAGZTgiSmYM/zmEqaTsuXke+bw59q08P9VLHjV6lbTTnVEGdZuetw
Nut9hBIbZma7RR6pLaJi7hCtIft6jaltOzI5W6+0+eoe0AyRA76hQVkA+YYp/VvJ
HE5Yz4TLvdG6zw6ej6jlXVyx0/lWottyFM4FeIvaJfqKSz5oO9C2hb+wMiFjvaJ7
BndSqAmb5M+Iruo0bUaWDQncWEe8m76vzwf+WTrqZHhNcriLovwvkT/QHTgDEKVB
9yOPaQ8j0mJhJZztdKI+0Isk5XYIGjLVeN4EgDorsMcWaaFSOpEc1YZo9nKLfrIc
yOV1Q9yliMlIUNoyzFmCx2fqOah/axmDvySDo48PltO/ixzLKeiUuifvxiShjy+8
JJ8g3jI0W/QmKqutTK0A5Ioui2XH1xQ1WOqPGgPCiGYv94/x0NVEjQyCzjWq9mCt
KQrbFOJokwivMN/1YfWRnqrnHDp+BJXwDPqh2GJbvCmJ0F+gK9Co3Vhfaac6q7XO
foaXY4ZerI0uvPSAuGPNGt5sHObHTZgcaYgYUo+yX2JO3hCVn4I5UwFATpV1CdBn
qiU2EYZYfvHMg3QTvPQ1hjAehQ5OUs64tSXVcZkr9iylEXJFjPug7+tUVmsMZ2Zu
Ycr4I6ER5rj8Z6UnnrxpyMRSkv6GSXZexYQ2GZ907q5NzzY65diIjYCq6kVnWEyh
P636SvGmEKS4fhULR38UF89QHec7KuNAC9mDmWceyFoNz5LEww8hGY38iQbeC8Ws
gzUXQjN0237y1YqaxgPs7MmWSG6JsXu2NksErdoOTXDpbOlOh54sArIAxQyON9kG
MS+Ja8nYIvJbUOALw/4yyKL0M5qNJPHiC2cjoeyzdvZSx9GlmVskqxvfOBpA8Sj7
FBW5Er+NR6v0y5HngGXAH7xZ973v73aK1Pc1+1y2sruokfuN7TvmSU5QJjZoxV3n
eboH5c5MrlrcLKJ8SodXkMSfpujqK0wGthl6LGVUf5hhyvAtA/jh4M0siS2QJDe6
0kvLQje8U7yj46+lKOTQ3p6Q61x/68lA/nNZVgGvJjeyCDbcKdpGPdlAiY/QoD/0
WyOOSzY3+s49I3sgpPi/ET6I4bXfd57mrj6O26NJXNCGBSlc4DyZHNb/6G6w8y3R
ZrBhcA/aCzTKlpwxGeXfMkZPUmAlMXFYiV4x2m3AtkKLrBdSBpTP/6n71LzMSwPL
CO7iK5E/D/Mb8m6UI/Jr7lgGa5XqbviG1bt5RoX10UQJ7U5jcrTFCZ3UqeaG4AJr
ya4sKohKcgazqlJaG0vc5JYE8C/rTmz+SDPA8xxQZSFkrSoKBUUNJyi8BLoFRR/t
ENnWslVUKiSLdz3uZbMJcXy2h8kczM9noRXsGE4bCOyskAa7DgqSDNeWdX2FLSQD
x7FOPbNIsRZuOQ8MCOObt6MbYNb/WTNRPiUMYn04durKYUfht8VWwFECYxbu4T3a
SPT5sA7ZUA4hjrn0xz2rBNPR6Aa/ANehBpEtqvukqRtS1lvVRq9GGYXpwrxPzopP
UgKcbxrq7ZHYLsnoOWp9pVxNjRB/mubXkXHtLBun+Xd9QW5nhactiju0DroSpj7B
vLipJmyaxaHXXuH/lj80KU3kpJnHGYTqOQK2JBiNvkUsWnlDn8nvE76Dgz+kfdmG
9ezW3Oeii3M5CFdoD13JRr39CiO+xo6WOOlnw/ja01zOczlsgkcnIANMpKVER2mc
ZA5whWWGrMxj1lHFreNHWO7npvEc528Q+3yTL/KFXccJEIpFwspoA0DeiDqEu0nJ
ma3h9picxg6q9sxcwtUmXOpzWMSJ4x2C9S4Jru1iq4g4Wt8AsfK1EiX1h7XkpmQu
PR27+8AQTKZwwp71jSTCDI/run1byoXrnZO5JfjhPT6/0Y7/5Sm6nBRgX6QPReXy
V7VowTF4+bew+Y+Y6amoJ+CpxoDHc+6VqNnUftIhaUkHnVxssJ67j9eXUuH779ai
CvF5do+q4GNFeVzrTv09TOeyxruRU0QTGQ+B+OefPbCEmSHVcS2FgEk9+7lcAsao
bx4amLz95F74o7pY/GqJhxFwAzHzy+wRf8GQEWxM8KJWvTFpsf4H3lZFZAhKJTb+
0DFz5ZHKhFTKGypApJtvwuB/eZt7x1LmgN7kWxzLQDAkObuAvEVEQ9pKqjtW+3nW
+akvmZROOMwRr34j5t113wAnYWT59MQyZIvc8idkXo/rDnX4EZ/it44oBzeofuBW
gExuVyJ7XapkGEOHKeuU+4KScjp03PguPFT/zfuU7mXM83q0OfIGuJPwF1A7nEvt
6Eh5peDPIPitaBi2FzhRI654nAO+1QlFZQruBc4s5O9Kh/CDcUQSQ9GwgkmbhmQO
JDDqn7mAAmssM21V/MIbYnClq8nDeO8aplu39DFdragy2jzsrNU2mMHJryUn+ixJ
HMwN3oeMXpyxp0lLlCA2PJaIskY3zDrldsCheFtrcY4bcoYHvd6H89+g+l1Z2Up3
Mrz4PbG0RYfNpzIezDIghMUXggvzucvEGdBIEeBFrWU3Mfbc58S2/+S+Q++ikkbe
tYt48BMMGSnKtTOXnAxazggp5yNNGlChiwAD5R7Ds5sCm60MrFyJn+0bHf6g4arN
UZA2/wxhHX/l8yaMLq7A4xwOjTIl9gSm+Uh4kJYaObKPPwUhZnKEqPZfh7to9BV8
L3LQBbaQKEV9COF3oMCOukH/UrxvMbALDTIRZss17/qZRKJ87jPwQVFa9bYiaj2S
fAvMgHj4O/EHbpmVKZl+L99dlCJq0E9AGvXGP+Dxa2vkryf2M1MYHERAKnfY/tJ8
XDRiXBPtDyW/FW5cjgk3pxrKdGVGKEn37Fh8z+PY/MnG0BBIEJmQnrcxOYexVQGE
byUOsB/4aPyotRLYfaiHclvfzfqs5XCPkokBZ/xOV5akwzVD/0PU0rKhH6VU3FV4
Vc3/3b9DSRm5yuQTftK13vTnwtlraxVOuzMIFEhA7WPK714Vh8Ly/BBWEWiZOk0p
qu5XAirI7HwnnI36yAAUFQa1s33COA063d6XIRO35dJKycZWxCPiYtWB1wuYcMK4
EIDOC2wzC4jMUs3j96O5lbjXpLlGmeagN9fenG3XtrkjzlqfRoIKio6ql144ybhx
ssO4/+aqguo9yLgU4S5G7c2hrL23U6X+8pO5+JfdV/nUPhjgtBrfbsmsPHnovvQI
XINborbpvSuyHDUiMY3uzURKUJm/1Ej7xfZGeVBRxJ9a5wnUrH+KNsGVOZasjT90
R4ikcyZnkyMq4Fe6SEa9fGTlWn1S00aeguLd1IDmHNXDXc0lLxurO6h9kn+76kGY
6AA0zDODVdUE+BD3MapC4J5MEkM8l/PGCE/4xFglxPA05ttmwSfaw36C+v/JfcBp
pAfZQbdJnMMl9Rdyz+2uxgrCoJRMYvTzBH8rw1AhBV7rAE6dqE2vBJOJRk/nZwxj
HV0tORG3Bi60MqWzVbogwCa0OdmOz91lfHBt8TuBesWyF8hYoIacE0yfT04TN2ea
kyDRORaLaDklKPLulShzpywhitW8DE1LKEbMTWAHFwvpQ7JIBby3zK1HEmd9/So8
n77P55a+SIopJkZ9SVt7cBLAyJh7BzR3ZhYP7ij3r0PBMumhjKo804R3XakIdf/F
IX8ojvYKYC1LPGnJrfJ4eUbvcnGOJHmYc7OyrvKPPSg5P6u/2Q87mkYjSykn4b98
W8KaRWRQ5FHJ/F67iCBXEvw4cxONK5/8UPQi0RiEx7c1cEyWLYnYzI/PFlMdnAS/
eqIjAYnXTBXf9/vT3GiUUQk8ldnTy5euJjbDWGAUNFfp4UvJgEMQiVEjycZJDs7n
NvhkuzrIV+LXivX/FdbOAe+KeQRtX+TQ/YOjy2FAFvMF3WyLaMHuTyxtvzjlpR63
rNo/5+lnGxWyKz2JN7twF93zpFh5dqoHAmwCz1RLNsvYTA2Ph8bKZxLZyrRlrCpW
J2PBlWtZwjlB3w57A+JTPVxpi+eahrdAwc9PpzANzrmmbNaXY3jbwbKmmiZKPxjG
32tO/Ou1rdrBpghJNwjM7ILnJMZUfU9TLPPmvvC2oPHX7hLIrSae9zA8z057dI3W
o6VtBOD9nGk74Zb4/VJ7cCmzRNX3R2S0qRwOs6KuvCfHgsO+rO1vGIu7Bx2hnZYG
lCDP2FymRELV3O9eBMOkzCouf9228L+NWTyWKx15mXi9Q5jNJ+hmmPEk5QHgYKAQ
X6vDB1PWhmNHqmooZfsSbhCE/hqTVJO10WREQWAMwCPiXs/c5ykSLsq80m8Qkkw3
i78oFLe4GdpqGbxMJ/GBldM2QS9QheGUkP8WLBtsEs3k1a6e01lK/DAOf/yjDyJj
VoDwTBh/0mOwBYmPmLsbFGU3T0vbtt/sIypriZjf3mBhTfLfTk3FGX1nCgYelWwW
2b500UkhXkSWOJ8+O/2hkI3r/LdeY0vDNcIplUwkDakhNNiQwlYkipHfSWx25xqy
GjS5o7lyjS82eu6w635WcwJuuvzkQ/dOTgihSNUmqKPAbVRZshkTJCHb7j7tr0rg
cy68AgOb9ztM5Eba+6ZQuQl2x74x11zt3h9LSddf3Z4RQL8gbEdM/i4fbrxfbxlL
tVnGSIl23+BwHn9J6SN2XEk3JgITxkhbbiPcWg1H4uqzkcyYqC8oM2fi8LHQDj56
31FKjhFX0Nxo0T9npQQp56jplYiryKJtrMYD5ls7VIjqshQtzP2hZJX1YZZHuj0S
+EJq6D0DFfN2aLOW39a3SyqAGy0GF/4NTLE6GbRGYPTX9rGV0pZJNddgP2LXS04I
CbaOjCY4b8I+dRiQa/HfAxBfnjjzBKyOnyQljrIggf3mTzJJzewdoX/26MWls0Cr
80my1MTrH90IpF10aflr7ZwEo6hmNxMe740tx/lvX9NcHH3rZPRl74xB2MENlopm
lb0VLM7uHu7Zzgg+rm2q21EaJqGq8oWhmSaXV+DMvICpix8rW7U6ysoHZutLc8mn
waqVx+WnyoSawfsdSBBBfzgU+tpuWMaMdA39JUBUxh7g7QmigwABXvebzDPKd0/Z
ksVB9acVv1p4/MiwoZ7L1BsvR4nr7IeW9UtMZit2Nr2UPrFtHJQpYqdAkz1lRPsi
hsbb8+tmqAOIFdJezWvrAO+B+dbpbN22ziklnUIc4H48JB/6lLHalyIvXgLgUh19
84X4ANtwpyCVzZeAKFr8OlMh31F/9Tm5uVsTUV3f9/aeiWHBXk0FyZy0VwXzGBEh
nRUQnomr+f9zqS+cN3fklUZ3aQcaGdwRZEgNWIMxUYt5Bk1l4i3uTzShE5JuJwXh
/aayrpiXGL/HBpXBy7EVDqctakDjjbtmf1ei5KjT701N4ttHLis1L2MIjEmkls2h
tO2driilpyK1PQNztt5ieuc/94jHn+roJGwy2+E1aJxT60V+Iqoh7fvMblcZ4o64
xhJZIoW7L9GiA+gbFgo2hQkxSDc8Ocf0x3XovpHCWm8NSo+4O20N69Ahr/qcA+iZ
qD4vMcjoeeZPH6SurP1/fptqBlRP2U/VvEyuP+Mw+ckLPk2212cSDQJ1bC6Bq7mW
8f3pYNIo0JI4wVjUejypjrETOtcdL9XyXgBmMzMkYMWbjKHyOPaBp9djervq5hN3
bYEl1emfWCMUXWwMNZYfoRhhYeoyujHTKfdvZw37BsG6fuKNcClflNEPNGX5Bbsl
VCD/yCTPjLnboL4alfSfVjUr4rETeINxYLM0y/2VjJwPPteSZsoeZyygijnP9Gv1
Z8aAi6TM1NQd8qajCEFVYtaRo5GuxiupSDoKJFbRoBGBcX04DEJUML8DDfLlDwBO
oYIbRLC3KxLqw/KRvn+OK9Dypknykac1BVta8oMwqxV4vGri6A8fRWvnnTQkPMin
sE3rTEGOBEoj9BH/Xj6+makDK3KO8a3SjEGu3PspMr06gPR13pUu+yp7d1kMvkM3
rtY1bzr74qTkUgIc2/gGmKQ9qfvPlblOrkwZQWKK+zwvwOcf8Ag7lYdm5YDOhiAU
H8hBIH3p1Tuwc/UAklNgDRvigop8GRIE1KStTIW78HfbEL1A7FAFTrcKJHSMjkHS
+fPYIxMGwnkan+1xZhxfRMljoTznBi3jDw4jQsTQFG7J3vS1kHpUQWw4cC+jL4Xb
+UT3OgdZ82sKf1IUyE8kDxERVlhzIHtO7McUiMi2Z6I7M4uZjC+BwIXCDxRkzslT
y9f6EiNEyKLWjavPw7nD/j6IzRdHoGHVlm0nUT0PuzMdZzdSqcfW6lX0NTvvHTOu
YzICR5qN1knNSzk8uEL398wEDWLg1cSfAj4ab2ijJbN3eTpXkoHusDgvKvSM6BgG
hviLE1gAo1GAr9iqMoTuN1sOzUj1B3NA5aiw+sj9pIUdZcPrTVXCIcCS7OmY1kMq
W1/LHAKZvyHeMRocIkPzOd1CIcpbquiLbTWPiNfpFaEfanQzm79N37Mh5XuDJPme
k2/Lc6KC6LPkXSu/Q8e1+6rS36clgWEzRYK64hXr/2w3S/rskLXwpVbMPCGMOO9o
/qS2g5sfr8Hr/wRFvuhRpR7AJJ7NxrboXrvp/LJKh4ewA0OioP5iwDMYC6xtZuwv
TRwB7yxkhqqVCJ2Lbd6sJ3AXbvI0R0ihW336Ty1udzfyagCo/3N6h6e6fZ7yY8PN
AQqQZZn3PtA42kE6sm0xmexk6v4rZQpp3P2ZkKZj38/3x48MHZMyanZeZ7poqIbv
+0RGpX7cano0NfMAqLtYqbmbynhvTtUkDMHmRGWDxinhRxvAV7puoDqDpvjRdgtm
RgCPi/RD6ws8eU6URtfWIQ9WjKSg25wQMRC5XcvyIKGFY6lSj2mxnsA+f/gM2ehr
SvtYEAGDxNx8OVlWeE5MLEoKsR9EvxnpIdjWt3G+SjzSGy/E/kF1u3I4RmJmlYQK
/+gA3k3BnzCd6oF8sQvIZk4V8LmflujAQ2AYsTDYTJL0JD08b5eEkWyIoNrgP4R7
fyOjgO0f+FcO5Hdhlsbw1ms+5YqfhdW1YuYBVWtP3RID/d3mx8wTfv39iguIzSx4
Y1tRtsWdzCJ2wU/evYcJi21vHWgrCto/OSmtxTE22y6QJdgTZ5TvjSdDf+kdEt6D
i4/DaOHPuG2erm3eTH+O1/5pg+yZEjz4RyqIDt6ueAoC9udlAdD9gX2m9jn1UNCb
dnh5ftR/6gG7m2YFm2fNJgV11INwjOz7ACIRmoydjodWHosmI198PqaaWcavEb8X
fIwOlPfF4RkWt9w0aG4JDCPLd9pKnjYhmfBHk5Ssmnkfg7WBAZn8pzLpjr4LXK79
gEWk/+ka257q/Z3vLES7lrLyEst/F0ESC19l1WlcYVUGYBDIYuHH0JaYHpTUk9Vf
rOIypL5Tye91wh8EmUxf3GLxA9cpsfXLU6uIhvKpiq3R/M+e7w4tZikdA9g1k7IB
38jH/FMzdo/xiNiRn20GzpQJwOlMId7vbny8NcnBJGDyCWGYS057t34Vs5My23Zs
wYSLktmRuBfYlYeEcwSBo0JSin675sIg86NdGGV3diSKbjQrL3iSoqYQroVG9OBn
AipUu4g0h31wiKG7yEo6xouJSibFBkIOqE2QjYCVOlRppm51COtiyL9Kqp2QXwA0
udfOTh07kkZPDS4z9geiQwhUhypqd1m03ma8TX5nuzGYsu1cDJUrWmmuyxS5XAzJ
BMLHgFi+ngXNxGwzCmSu6O0ipiomjVOixrhkMzWH7v4lTm0fBzA1eSf85gFuCPX4
RFcEnCAzlFP0DalxVJXEywcklXm05VrhILvvjL5MH0GdijLj7mln3BWNssSX02Tl
TNlbjXrtVv+egiAKbdFiu0k+QxAOzMtDD/wl5LyRJaHhmgJz9fHqs34e78Qhyrer
p9JkIWIkvm8hj+FUMH7qUtK5gONuoG7W3pzXp9n/ZJwIi0qNO9IrwmwxLPyMW4yr
vxdlcM5REHxWzCQiAh/DC9a2gOQiDUOdUTZyA3odxUIGZ7OI5pkmM86lLdSLAPWw
gzY14WdpwVq5Fug/3kALpVQES3Hl6/yW2rXxI3TTdZZ3lIHupVz2QR+mge9NQzIr
EHgb7Bf6ydThiuiQqPZaO2GxuPhwNbqMcGdIezMitZftFH+jr/DuqHC1JEuexhEL
n666wP07W6f2V9ovRRlpYCYaOmKv4//uRK6hv8zfV0nEf0jz+Mk/g+lO2kjcp311
Jouv3PAZ0CxJHzTlNXe193tNcZ/nSlGA53kLJBqL2Et/eU1nBGxOzGrH1VGmISpW
9By/kElBJNDjC89nin9TJHFQqGEalUenFnTsQ4/zy95F8gRurwhM75zvUdz9EiD9
92SBnf3S2dK8Acz8SHMt7aH7kit4hQxC6Dne4K5Bs8SSf98J3DAXEjhdT3PjkWUH
XGUEUDaYEH9YaqdYoymIHNbQrjE2KX49NhyQLJarc/0YggxDImer1ogimaDoFuk6
USdlngym7LZmEecwGZpoUUIIfuOylamvNqIunaHFFpefUeUsBqnVzql+YMsSBv8I
zJHn1cctLYCjbJTC/ccFe+oGo5B4ycAEsP67TaiJ5UnsWZgjtkQ3mN1W6WHPeQls
HI11amCvpPgKlo8cr51A73f3FsUGEyQ2l2kwzjiPfIgqR2voCn/e2yIPxA5GTaHh
VOGMRdb05xIhmqAWPEGnxAF/ExMRlCV1qUctf9PKP6Lb8dJL8XlQoZbGO9St0XQB
5rYY10ilGEC1qtm9hzsvJve9E4rRm66cd1umekJJLc+bHNDYaIv+9TdoSmRlkTNz
vXdTp3vvrVbZFWwd890UmhuAGMJt6cja93D86sBN1T+htSglMz5/bP4sHDf7LzyH
W7AiU+jO3nzEWtnB+jk3tCL3+S3WGswxbEVAIHp+BzqZ88Zbx9pv8mNCPTWYw6Sb
3RDQkuPs+qFcg/W0hBIPTjA2ivJylQ5TPEAzYL8srM3ZyEabzVD6HJEPG0aiV6oy
AxSDUnE6Rx/FPI3zy2LLtlvmqxsZJCN0VL+XOaFBTuYYjpRk/SH0mzmNlfUgT6s7
`protect END_PROTECTED
