`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uyTzV+Po0PfHGGmIdu/8Xoq2Nit/QxLrrTDVoDQVeI2JGdtIrQZ5hO6OtvJZfB/m
Toj8TvLrm5C3z+V3HBt/u7X6n9SHmUF11gREir+OX3NPswEGGkBMJr9ZMQF+rvDt
xrHRg20Bvm/NO0H8OkJifGNRbqAeMG5Iif0JDJ5XcryDDwNVUO/SA+mUeaJO1E4k
lKe40Eh+U/FjCrHxm61gnptpWdSkN71nFWUhVOBlvb381VoXhCsYZ56gT5Xi0CLd
A9k5t9z5zdaFbmZ8g3K1ltJMXnrsWeaR0sy6R3Dlemieoof+8adLA+0PuUGPUPs5
S4c5YmgViqqvkpiJrBHzxp4XUsi00dmHO5H5goLZ7o/6t3PzjRwO1/nXzUDg00nH
lp691PiDeYEDN+MXzJchSbprn717K7/w5do7bj1RgdnIBdk8PFyVCeSgMpVi3zvK
QVovQG0xEUWe4dxQWCgD6QRD687AmGjg3vsLzYL6725XO2IRoMT9VqeGrOh2iEt4
Q5XoiR3yMOmS7OBVe+4P1cl5y2aNG1auCvup+h6EJw3g4N9ZDz/L/J3NoN3yJpen
Zj+fTabFJq6PxXCKl+mLfuzh9Zr+edNW+ISLIZhmppOEAIFo9e3aBaOn3ankMNqi
/U9CBNasPkuNTrb6vJ4pEUoFVrmNAscd3DYOWo8yF8mhBYlEQ/JbrlWIxfWL1iZ6
+895f97/UBRuCDKSYzJrqjQFt/xex2zGEgOKriHuPqAhhW6ggG97Ucfzx9dqMVUr
I1GAT4SeGb0zaQvIJ/+aYTjcQCuIDiGILBCfsqSt997J4XM3E1rzk5X4hZVVhN/L
Aluh+TEAKpzlIUQY3fWMGdVoyncPE5MBG/zx2R4WKVokP61Yd8/RaecQZyTTD0Ju
kQlFfHU2MDAZtRKreZ/byR4MpMwY0VppprITEB0CbBUt9jBS0dkX/bNvDpj6UN3h
PPX+gq7cHKDYKULvEg8IlLbHwrsOfxtR9Mi/N9gYQSVRBX/J9VsBDMbMPuT2djqN
9RI8E/8Vhl4N3r6G2OpyJf2jSAl+yzvFBT6k77T92/LirCzqvdCYNvIXUKoYtwiJ
qJY2LnWNzetWNW4Ihkg/TCCbj3yAUdNGy/7yGOMQoLimzuQE7OtWaOiojHy4+Sl1
yb4PnykU//tMZxfHAZ1ABQ79Ntho132Q7j1efXiPLlpUAsSCswBCd75BsO2ue6mF
eDl7HfQtCMf/9rCWi2cdiglre+Qa246ZPWY3FkkpmyzN36wJi3XOiZ6GR1AlVDQt
dYJhbc47zmvbAzLeojPWMKJfFQdOJ9eVl4FzFhlNK9yZ2WzQz0/7Y+FP9HU4jATD
m4cxwKQlo3FSTNNG3ZBDeLVRFU5l6uXvlqqAlJvVXbLzlaqDgHOD+P2VzrtB70op
4p0Zk+d48RJUZrq4KTkIRCwvRAuI8yvCqDXOTrxA4JGfTVLGLjc1yGLLMkPrx3Et
zEjux0bvF4QU8qtnG/eNwq3+w8LClR9kclORzxX5qXekN+NF2PiUb4IlFnkhkzHC
gFTjEIikMfpAS8SjRWfw42P8MNY/9DAkqwFIodBDZBDLItYyU7AR6T/Vn2gaKcPR
N0FRtCxTcymeljZDGd4FZBVrquy0vv8awNrb+qakMgufAgqfOGKq1OM1981LNfo7
FzhfpaL7xqTECJqrLgF+aushW08uA36JLlVyg2vEkdwWF6lhKUiLNVslbW98IyR1
EwTu1+ocxrWqEwHg7Jr4Ck3+XYmL8D+eGsX61d2s76JwOSKwv8G2ArZ8H0miDqmk
vJRu+Vm6+quaxm6PODXP37mJDlixqFctQTavXBn6T1IoFWYimVtxHc/ag54K7/Ka
8aLAz3NEpYjCqHCfxa1X60f1rxVx49XxK9dfpdVhAwFnnw+8S8Qo4GtdcxMUBwri
PP7/wXmWmGzNW2iiPz0cU1j7nQBQ4LuQKKFm1uB4te1sCglqWFZxPyuZ42rb/p2L
6/n2lnIOsEAy5RddQqm89/iSK0P3zlr1G0GK/nYAkjWhJmc2RIw39Z86pV1QMBLj
aps9dpk+fvm6GPjy/VSV6enczsOAUJihtekkuZb1mDKGitfGqHDVytt0a9qE9GZT
g0UyahCf5qfrrKl9yk+CfFYb/xswnL4eE2K9oapM0FoR7q3S04exYkQATN9f79iy
PKZtKE4gk9v9t5zWJryPdW8z0hgtfYLeOLawrNR33dD0N71TWeDlabXz9oHJzofu
/gg5DoaMkmhYa2/WJ7B6xrb7u+TaQvseeXEiXjOWtc7ttVBqTgQJX7U0zI4HnzrK
qSWJ0uTdlmL5OAeX2rbOWAHw44oNFORUY+RIiM4AgYnjqH3eLfE3f7rk5sIW/bGA
vMsPW99sxZ7vaw813W957ZlU2jv0xXc4XW9XTEiFjsfWllPPTp8YdpA7vVnEOTCZ
xcWZUMHMeRvCkCwVTQe1TnB0HTYPVxzGJh84KidydzQ0hkbPdKcn719R7brel8+w
VPmJWYO/7YQHmeSz0wkkooZRnopEWC/XxNpOZCzDxokwJNgqvfOxoibCyKIF70Cn
JSSieAUj0F+b55lmGx4HWa1YlD7+Nr21x5egjuQMqppWw2GeLYBPVUAoMhdOkvgu
muD1jPvbugdcFC/LRQlTT1HcmMtlv7EhEaFKcTV9jeb0pBblMZntZE5d32SwGO3C
gcKVceBKHQh9f5TKeLyw2OvdSbEDLHOL6qk8AoeF1ukZ1hyFD6ooJ4mixRVw91gu
EhvvhntQ3NJSo4pOkmTvpnxs5UqBpCqC+davN8lM5XZ6gI/+dO0rXnSTKgWNzpLq
+mb1je1LPZT16+R9vSXKB6QPhZVgk3O5OTbC9vbUKXHdFmNXGNJraYMrsPT6e2tH
YxaEwWt2ot6XPWFo6WxypDOaM2xqpzVbon3T6wY80jgZdpInaB0KV8lcc9jDgelj
QNVS5kQxQ332oH8xLTs/4F0rMUrVBiZUyrFBWYkJR3N5g/Sg4dbtO1muy9P3nshZ
1qsLfn7Tafj4/Bs5m0NfPDS1DML2jEtaONfQ+SeAjQB3lfbX2aPiWC22lYwDVAEJ
jBraeTF6FxbovyAwbDpIdNj9+yCLgtwipIGJraHTBQt+SSCtQUVCXUKSqWUY0fND
phO8HBZH8ad2gKP8Up23iaPZlKsKD+eIRiqOP1DPi761j/A0VN5itPwt0DdwkaTR
0wZqE0qQY3Dt+QK311KkDTUPraQl59ACOts56EB/OTpoAZgAuYZ8Y8uZlnFKKz8a
Nb8b6xFa+XHwTdTLFGnLEP8lfuy7Lz/AfA8PsOHdcPSgL5Maa3trr7x5A7dvtLP5
MeZyDetiJtVWD4Ck8/awvpsIBH/p7qUU7lFosDIxbur/JlBRxz4pV6XopKdnHNBv
vvDwziJmqZzdFqTwVkhp7N0iaT1dvca959mwfCLwcM4Cj7b7llsfV6A6ko10N0ME
3NazlfUG7IssCzSRyA1T+U19fnEUZsMi51Zkws3qBWK+yVhwhuaFCeToqh/tl82x
rDVVYusSCDYJ95hSEgP8uBPfAY0clJ2tT2tx8PVXkyzfiSAWFw45KudjvMn3sCyF
9PIFIWjt2lWuvHyVQx4IzpRzSjIMB/YpM7pLpUdtkCVSjFzHlLF77Vkjhmdh8Rv4
j94c3PqEBlPxduNq/KWnUZ026xUhTft7YJqdjp6Bj605RWoO7Mhpktp7xwt6JmV8
B4uwnkJ+sxHLCKNq+SlwkbyA33Rmanm3vCQSTK4casaP5w0kg6PKKOAorRvTuEOb
ilZ1IzoVA3+JOeYkDDd6MP+87QenXF9U84hhWxkhFkUV18iS3TXUSpHd41IHKCzs
SYArGDKvrc8SjZkvZkhGbyUgsg+jaKRZBzsrn5zqRcKqPf4z26fF5UeHo9yY3xjm
dNxlOOIiW6cKtYIe6Qix10/TFfICRWlIKl7hlyPSfTD1SNIMDDpCcgDW3RVEw/C2
91kZqv1jvLv1rp0iRksEq9LGRw1Q50YkB/upXrbgvVaOKyGrhfEpbJoMQokwklQC
TGZuO8sULFLivaS629RzJThfuuQroJrQUYdTIb+YQ9Pzx5iUiXQS26XDLSpz2Oex
j9LuSzquuh2lKJcdgqMvshF6PGjGVGM1X7j/qkJ3pzpukf8UYevfuTTWHGVvT3FQ
7v+Z0hp9pXYAYZMjCFSKlPOPPlHQNBjlK2SPM6+HdCzZ444LTQbKqD6/xTsFGTwH
Cg1gdjVd67yHbgFqHcU34lNa8P840r3kGz7qOYfBHgO3mZcOVOnb0NSbmPoJabTm
Jk9qjE56PAIuC3rd+l8HFKxL1t3E0PfPQ++4lXxA0Z2LlPWrjpVDR1wC+vEvaUoK
++zQBziAG2zOkCZKboUEgT1GTmF+QQxFe5P3DqAo4JflooD7Y3xccKa9k5IroRck
hZGMEPjvywkW1bmZSWjw+XKEg3KKcOvp55YytyGVlusD9ClyjRMyE581lHtSyjrs
yqHERhX8DMZJgqFTx2CqLHpONycrKd8BZZ2uA2qbQP0H0x8aK9UelhLmYNJZCGW6
p6/Yj1nuzsJZtyJ88n4ov3wXd5AoK2ZP5yQ+A7vB5Qv6m64R5Fxna2tE6EGF/Ls3
7tlh+Cc+Owxs6GtvnIa/wt5GLWUSKdIBZKTjF8NNH9SRVZeGJKJQaR0rqPaQKPuA
LB1Psrau4YY888Y6OgXC6ATVDRuRXUCzUS1fCBjM+7WB4PkC4NRXqEHuXcxhDIHE
QLmgGXNLPhNxLA2bn4SEk1Yeecqp/tBm83fLDZ7+6zMl+iNhqUfO9vwbu3satLWt
E7ymQtMecj3jOA76lIR5Zc9lEGkrgJhtxljCDlMSF0iWpnfDdJPVMoLoDbar5X5K
fAbaY2HNkm/6rsD4rWEhDtgBwihHcKJ5Pr/Fuh8NKjBq3v/FzpQ1NOZWuqhhitab
wdiOaXUyvQm+/tgHUh151lu0tCodV7wHc75Tc22yUwtZLyCg3OucdBVwnF0/xjuZ
c5V42Z/rJlWHTqlnHf8x6i2/Nt6Go3eRZqjtevYlCrKknGp4VI7hRCaVziSMQ7+h
RcyRG3pVU18XnDw5Nmt7wB3pzKaCo0R/3iCiYcMXqWhFkZeFjXO9Qll+kZvio/5j
8i5e0HT0730kQshw2PQh3BhOfnXOY8NJxM7GgH584YdGnPal8QJGpBIEMM6asHoe
I//J3vhYTp1yQIZTq1RtPrR43EEicub+cp7QfOovuOFJD3c9AJDEvK22gD8gT9dk
1TvMNC3TC6qEupXfjeE0G7JEB8SbdalTvy95XhhSK9DZpJSsvcV6LNPC4jPo3wca
r6JYk7oeVFXeoJy8DpBr+1yDr3XUyhbzzIDs5Xeomkk6qnk68zIVWABMrPrL9LGe
Wd2ihCPgWSKtziye1YJ5PfcjZBJs7hi1k/q+K840Ae1LKa/bPpyfs+r58kZkKD/L
/vHdobvc2C+QQqdOEMeGQ6+iiC2uYac90gqzBeyzjt4CxdlNAqvfy1Hn79aUN5C/
z75tSmbTnIDoeLc1iB7E/uVkkj7mApuwvAoi2NilMo9NaP/IIwTD0tvGEBvYm5v3
m034iGpY+svNi7xsSO9StcgEro7sWciEyl1xIzbJJ80d9hakjjwiVhuB29OXdpLj
smi+68aEwBT6bRcNe/ZydiJ5s3FvOjr91l9v7Meudk7WWjnzwmVO3UgAp6Jvy6Er
MLF6Mf3vE15qEz2mCEzTN5ARKVebfEF4nPiSGvGptN3Lhbh1fG9iAKmkhxxZeNww
GKDEau+Cm769EF7b1rWFUcKvTZtjN3FOmlxzIG/nhnhJyG7xr0d9ltOf1VFlTyCm
syIdtip2SH718IX4pWIl6ZufFF5Q9wFYaiFn7X7ekUXNDDk6/O2SeJOeoIJS7NQb
l9OTO0gbwIfLqdAkXp//pNIi7w5rasMYQFnyMhk0Y2Ee3iFIWtOqG5mLi6AwTfgv
rvQmzOguNpv9NattN+PRAvCil16a/ZqUhmae+t1byO/QXUjjXhGNMlpPScBwdZ7l
/eDXazu9OKlpf2SVbQBSN+I1A7R0EfMypkLiqHrQTckrry29eoyrooxKzRyinMN7
v7ioj2hiE5Ca5Vw8ZcFtoU+5D8JB+GtiUnWVZe+lvM5tfMlS4YqE3gLH0s2rz41+
5wUdxEpBs2BMD2WOHw51tAmDeawPsHzhb/uXeOA2ZRKAvLAbrE4+TsfZWI6KmrQE
E1i6gB/0r3bTCeIdLaUXPb7p3iaHKk4a/PAAvMPhjRIwaRkQJai9+i/MoNt4FDU9
CuwcIaqKpAUSqgsGDfmudUPIQNuyXvf6LEsxe3C2VRk5Q1p7hQAJu2moK9yZkAGR
0L+SEN/Nwtb3q46VLHSZfH2sFcAmDyR1dRd8iR2Lf8Y2wZO+O41/4Gr3b7+OYXNf
sY8kX45LZiC6w+FPZgtdWrHh2Ez2pcv2wLAgDeIrt0aWFTTptoqU+/CfV/59eKGs
fJ0FtP0Wp3vMkfmRq6lhnUB+MPh2j05T1Clipj5mc5QiIIhz4rOyD8oE2MfBvPGc
2wOk2Of260B3QN3hbZFcDZx2IsZzUkj3EXJVIMw8wOHPhdVxfAQVmd/FtVz2fCvv
59ZxI8KfEaS4oEv/nQS0ztElKT0s0fa3LCx9mCbjoXEkvjDfmISdsCuN4t9WY8Jn
NbRGUXJiYcoWnzY7W/nxFDv2D/zNLxNYqJeMdnAmdThPmDde++x9Fx2BVd1B6Xrm
oU7ZKFipwJ9LwivXSVazKVrc6CqVFYohUQ70kfMuYnVOqszW3gLC/w3dD0PQwd3y
3rXke6WIPTXe5ZMdZ0dHfoCaZhqW8xO2o93Ee2TFeAahYaRwzv0j4HS5b0kVmRSZ
/b5NUgWATXubA2kjrgPS9vGb6H283JdyaGzSjrMT7PKjRaIHej1OGt6v5PyFJz0V
15fHweRz+QOGtu0sqZD3qJVU86AuSpt3oWbcvUJuXsASdDms7uqZSHFzl/ffl0It
cBc4Zs+g+5AgZxv1FQi2dvu7ZNBnp57dXqi6r7sijD9yblH31WUeayzXrk38iFry
KNKS7GQ4iWv6kFjY+JVAepXRzyd2VnrhLzVJMiWlyifASvkuM88DemYYboFayZQ8
ZMkB9fHnVXq5nH5koJM/xdVXjKXjnkd2u35RM15HTfqCwgkdQ+L+ksyUu7xkT/r2
9TUgYmk1wc/JpSnLda1cjtbAUVgyS4oVSLSyinKQaQbYPttJE/UZSLk4XLmFsyDu
BzJPE5ukEc7OS4d8cheNWw+iDuxQ9/aJlrRAcGQgZGz2X0V+ld8RGfkGv6325W5x
GxpegbBmDQGQTITJBv3PId8REaxc6mk9r3EUyKC5T86d3G1iQx8mGQEKkFfrDqvP
NIvMqvbYBCj165vaF7d9zyx49aKn3sbEHVI8wJHTU3TA2qjENbinl8t9bXztRDfs
mzfDJyUEfsyinsAG3peTMHv1b28x9ktATOyrR4SCvMUmyXDl0ichPBMXANzr5BOk
B+gFcqOZT4NpzUN8RM7VZinqusUGsRuIRQGgOjkOO59/WfFvYTbOmq/NNKloyMgn
UVJ4GWi8IAnt2B19SZ20/pYKt9aRSX1nbjEf341H0eJ82nW+OxQo73as7KtR16KM
P0LzXBrfefsTxbwZe26RgqgachyE6nBgpLoLHmprISs2M74XFYeAt23hfupFR0jM
aRs40pyp/lgPq/X65bgduar+e0hTR0h8Y8PvehGS/9op3C+SalXvudXIbVbYclWR
eNjR7WXAVaoFL7tipoXokfwJBdE6tED7uED398dXSuUN3siUDyj/jqGXN23KT7/9
m2QTzabhGWaDzq4CPspdviiowsSQm4xceuwyrEQ9Gm6RKBLGf48o1anOPQX2WfWd
PScluD0YyKMwhbcd+P/WrOP20q6s9fUvvmd5aukp1XZJKntG31gaC001DQ54K3uD
rzP6SopL04A7U+UsJsvG+Va1YaEkNwjo2YBPt9vAdM8BmXDrQyMlg94sxAgbxett
X4RuBHsP9l0HxKFDtIi7p4ooY5IsHtO2o2nvf4E1CsuMYOxZjFfljvIUWieOa53Z
hke5vizfUjA2h5h1g37PvRNpDnxVYJDJkLUZdpbk89Qcb6HvCKnRm6qHCQi6NV49
l/UiebLIrdHykAfFQQXZazaDYBSAqLhv2uDKcWTUynMM5B+H7OLYVV6ZcJHKhl4S
nzfWE5P/6znP3Krdv4gN1J2BfUIrjjzsgHScPQWVWCbbze3TFH9tpCGZo2+BD58M
5VUX/IkhJYWtA2DhU3KFd2/NY3sXgsmJiniesNZq2IqKW3QjqTKx7+FtJlmkX+1i
Lc1MuUxFyCVo6MjT9dyZ3krsEELdyIEB8ketyTrCs4+C2YPrd8kQ2X2aBT6WZu95
H9jsTuChPf0hWPBbVshARj0knhTQrs25L5DSUdCXO5YIFfHvL+jqFb+XUnRmzY5G
a1M72g3RnZvuyZ5caRbm9u7jWCl1gpK1xrvUrrOk2ywLiXiPh5JDH2tf38c9W6CN
eiJ8JOxoMnHH8XX/sgv1KxfznCkC3EwcOWpA1CqrFJOoW94JRnf36Qi3AUWYZ9P+
XdTyRzx2vJ1x5velCw1pXxKhjfDkV+uri1tUzjr6Ptb3ecHiFQpYJHGuD3SHaIFf
3CbPBqmR2krUDAsCjM7eqJbhspbuULbWMJ+jDZdVukuiOegiQw38AuAM8/PFEl8t
CwaUMmXKU3Z8xpZkSzxWq/Hbh2WSmEfvEO5HGHp8vEci2P9GouyZXK5viT9OnyBN
bJ1ckUax0RuizyYrpDPXfCC0C49a6Ak8sS7l2NGsPj9KyZ8APdxIH2eYGxtNP1d2
pPjIG1v1AjuAWa/dHYPRyRwuKYJscRB1Aq1TpoKcXA8XBM/E6hHdSFwXgmYHXAEt
JdrklJj4AyccZoOI4Go6H3esU2KN+fKsYs5Op7mds7RO55yXprtzt6kEdY2EzpB6
kMtV8Y/EH8Yy16iTU9JoVdO4BVp78arkbVnUfsr4zzlEZr0AWO7c1wTdjsDB5Jsp
d4oD2GhjsOLgCeQMFc8y7j8DhwwkqokyykZrR+HUGfC1iiKUm3QJe5peETgyyAzT
7yQCI97LK+LfzMoKi/00G4gjiCVEpkX1h2xDsU/UzWMpX5VfnvCuQRcWMbcVHP+5
N0ZzXy4kxVDIvuGWu0DShsZ/0VLBBnWlwx6Zy+e4uZZ8HT7OW8QtTpl9tkfGYtsY
dtnOcK6SrxEMToWELdTYdHZ5gIYMCFSp7iZCOYi6EzU/+7J+MFslmbIpdEiP6rzH
CLkM+b73opCHuYe9TSNDYfPu4Yvhb5C7IguqqEUs+hdbyRJyhhhn6VC/43+2SVZx
xKwN8rfv1SEr1Oez+CNdT0tIlpC2Y7u3tNW6D0XK6m9HLjKKhCoqVTwnoOzdSpr9
M0V2k+WzZRLmEs57kvu8NmeOxxZOfUHtL6OBALulhNgRAuuW+EF1YGtm0hAAwbXY
eGP9UqD3XzNDppTY2Cc0I+y6Knc1nYKZuUC1BUDj5JpaKeiEfCATKeP5solFRyY5
UDBL92kt7wmK2bbxrn8FHUIsTXCPqTBPo2nO2ZDZ623SbUNvt3RJ66iZm0Cdw29l
lhZICxX2zQuKMCyub+sDykUSH7nfJYLfmCgqwOHvkO8yOn+GxiQKNN+SGUtlF37Q
DGFSWNBGJcP2D6RHEEZtftxFPZWbWj4jAqG+OC4AlO0+QZ7Nj7xUtfQHMAZM5bDq
adZJUkSqEfTqmgQ6sjoW5x6y9adw3Zuw+kvXVkrPu2Hd3Tb5jehKMwjp3iTCS5+i
P3vdqt8dCy3mTT0ntpPx07+e2XOOxYfsTbcGgwD/OEUfNTwzOEFuYt9c+SJgdUps
5ZLtEZv1nlkIZP5iFqt5aZCbsked8/j5ZE1ccwCr/qQTLfsqTdP5PiF7N28pT0ij
KO1QhSuPdqqEPtdceKubzKo3/FbFODKFR266v0HduAg+gwrdXtnUnFzXaPCUdlcl
3WZ00SXe1w2g6SmU23//GREOm4XDonoDrnYvFSxN1hitE1GT/Seg6MZCvujdFqJf
rr4YvfbX9VfBIiXACa/4f3BULfDajp92nCzwf/LUdabaz2WeU0hs+23tT+hFGoac
FU1w/XH6NwmGgM04yUuw/10cjUrSfZTm6Zkrf7+yIQI0aeRkSnr0JxmJhLBdOXnr
rF7rIc8Pk2M1zyBl4ScV+oxuV0bp1K1LNVA4o5iBOiMKHk+IbMTUZt8jIIOH/EYA
dy6GfhqbHSJbqxQwAwyxSo6bYki6VzAXN2tUkKMVNaIe+h7buSjPuyAPiawIheJg
JH8x720gRR2sqRKO/bHb0fBf4CtjhoHgn5jTBc15Q/ogBE88QW78ZlUy/UbFZIxC
8aTFRG4I3h98WKyFSNVepFOqmBAbw0L/t/IkpeZcTgobO3SQPHFl5zaZzzuaLurA
rmvaVdnR0+xXQoaJ9bzmEkkCU7Op44sV+5bVUO+URmasILQsVJWzcoiTvbmk3kzg
ejh1UEiiqdMjKG5H07x7QqgBxo7ZZ/oBxwXgoWRS07vZf7b84wkuTPkihZrUzCoq
iU8wbXdhrP2nDRIcSTSMU7Yg9dzXoEL0xRbbNGsdo0K0a+S9IHO9smUnxnd1SNKv
L55dHNt6CEgAxwDCOJyXPtGBnJeSr9PTVmAlV40JsO00RbGfzOq39zWPLaP/a1Ki
mzHRUqNEzN5ErFZEfYZfhxY7Y1Y0H18uTxfyePiFI2BtQNkRq84rtmgFc1sFQNp+
dB+RCUkO0LynPo/L1S7eFgtabAvv/9JaQ7uDMI9baVrnhJ6766qOP+/V1T9AHCOC
rq5vBZ7E3qyLtt6AKBUZ+na/v6BYx6xau0Qm7j5AoLropb47sbqDOs7UM/kUU8Op
vD186IJahoHUgu+Cal4IteoqokRDKuIOH/iRvOCFt8Wl+u5rR4n5xDTxCzER1QCf
QFuUmZoQAk80wx3wo6NnH4hOnjICV4VDsqk6fybpswdr286JQP+iB8Z8A8Ef/Hed
ENtTNMCAjbHel8RgyEibTMRUqwM/ZViKBxitjwJO66Iv54qKLJRl1jNiWz4/uoC/
ERRTHfzLLr/jtq6Qwn57Jsb7Cj1N7Q/6L8w2H+7+vEGwN/u4/8J1fnMRRZ2+gF8m
7LPUkRApq7zKWVk99KKuow2Unqk5686SlUP+RGV/Q+mK+rn+V7gg8TPmGSx9q9Qx
lYwbNHQn9B+bpfe+nuFElvmA+k8QfMlYRHvvT/pSsyoW8CKApSlcmXdjKYn9ep8/
rvjSmaXkJvtxsRzJ74jmxyetNoEZwfDeBJo4K05tynOTZro3Wl034GCfYjpk1k17
udlUKU7bFk2GyrrmyKPhMFRUe7mNvfTr5cmcLwIN5jBfSjlUhBxlOxqbkGnx05cA
UCQU8Bgb6y2jhWat4Uge1zshJRVLpNESNK/ul+xRjhixk/gntsRvAoYhFKQTO4dj
1qFFFlBmA/3ShQVY0qcis91xjoFno3DLLZK2aEhWhCXxmzWLdvT9/uI9cEgCQDZh
GJYNIHEX/Q2ooZNZKH0b3fMwbRIKuMDQAhBS/bmBt7PKTGB3jRZJuAPh+18lINKC
UpyWeiZnVUCsS9Ucqa8qYrOHkcAmzhjvMKrNvCoWta93rULChDNqhTPe2sdMNAdO
QZhVa9mnbyV+K+3CBIoQPlgRL4bVFQ0Vc9cOQSjNA84pA9iDpL84HWmuYS2N/NzR
WnPjGZpJlQiGCbrgWnVBs28KgXX9bmFKaUZ2yw5oRprTaHXkuVbnVhq9BlVI4jog
R1w0rU23SiSduMGmEpYENCVngJku8b1Z+nF4KPWg1cKl6IbVEfQk0j51+7ZHt6ZL
r+uO6M48t/GXA4CluYIpkOyxrQP35htwXpUtsrT8G59p6cNMrI2e80CaVj7U1znD
SpJIpvYhNCFdhmD9qnBR8aNpPK3WFOcdMCOVtFCHIXe6SKI2iqVPmkZNDPAIFsR3
fmAIUtSgk9NCTr1OUZgPlFSkui/yYYX1WzLpstz1SuDDyFtenBA2IITrAaTY64DL
oQqzQbgTjR4KYpPYh6uD8Zo+6P3O4JMfSF7JAw/etDpQEXIWs2vbeDuWRecdK6ei
JayOtyb0h+eEoqAgOlVmToP+fOEN/G7D/HmZxfY/LuFegxIOO5P9+2VQKsk0CCOi
Dn0XgmYhN+g6YtRVZ6isno+Xz4xhhFEwWOVlUL/UN6cQUrgv0kDAnYL1YqMJxvUI
1W+v4WL+7ls+C8F2oAwdUxk1dDs9cyl2F/yuN6hZIoTKfhsPUlOWk1nsfD78bIZY
vo57UOy/fzJ1bAlS3wq7EXKJFstUo1cWJFvR56eDFGTC2VIUQGiNK60DXSXlSwlY
ohNQMSP/0IT8lckaGjm0Lj0GXUhw4QEIXVw0no4f+n8/wnVRNW8VPixjjwg8V4aI
8eDtRJbN1fV0aThqLzkEk4DgF9foF5x0+1yNxlXox/oA7MeHoQPmdSlCEuhYmltW
BfdfaudRwqPCCP3TCXQ6PaUmuPciVtCUt/33GKQbjW5sE9l2BiOaqfewdlUhXPHs
ibctR/GfFwlDDL9RtyPYFesEfG+eF+WirITYewqejLrX6fY8FqwLfptYdktUb864
JMTjI0FPxvv2uu/TE/cgLnooTvJWxxi/B1gPId+xnMFy7z1unn9n56WVXa956+Dx
VrE0EMeoLxiQBxubTYm+dYS90qP0yr8NNxUwWUmKWxYbtaD34HZ+bYpcLdYS7gr5
mBDDOYg+SVb7CSSsORpPLg39kaWXCZkfaRYA6Vk97AD8pKj8eklNUNi/IidBK1lg
QtASmYHwrIt5pPgkwEhtp3CkjBiVi1IjEWlhhq1KoF/6SPWo6AGmfiVpW2OyQPuT
MNrqF141D086LR9RM110T8QDEZQntzNT42bKuF+R518sUxTr6kft+OlOUMZnRmuD
p3BPVLBMC23FSaOE+3Tdk2LulwRfxnmNuVF1ToLTx4VI3+/j90vAg4dkIGMKXaZk
k+BDMSUKLsDUKcrv/KXH+HVSl76L4aOT0duq0/fzfnp8IABbLWQNEZPq+tYhflRv
81FwZdbUL48wTmtPvGF/ITt5nk1smaSRPhQO7A29pL+KLLfufi+60EJJQcQcL9rK
5vRvKUbgyvT92tybvnbIoVZEsmHKzk6WZJ7E2Xzyoge0WLtXP3fvaMmHMrWCR0Ow
uUtd/TJB7QfZfvf2kU9DqVmvZVSbHpEtt7KUCmEO6QqhkblcnYF+TwYtVGxQW+Yj
6PdI+tZM3IYj5RWqyb7JM2ReHKnyBvZ02Rw00kNi2FcpXGJBE45sUEm90ZBswsEk
SPvstuJHTY0cmyRP1CBScGvX67MpP/N1xUEs7j7KtAWHgiamo8PXT2cPAQlNk+7S
lE0F9DSJbdSexuLmFwjvnaxPo+iMiVkrLwIvxDXbOLR40tU+4/YUx1SbREw/CZ4w
qhY1782s/NvKrQBDqaU4ZgjWjHzIikJfL+JH8yAp5Y2Vv6ezmvRfmMC6RIYruquJ
92H8NiKg4WV0BT/wIWXUbKND/1b4VnqyUnF96022PBd2nhMI8+r4tN1619XXjgYO
q4JqKg0HJ+4VBuyAgoogjx4F4ZThnxW7AZ+G7Xv4PtTODcfoRWjJpP6P+n37C9vF
+eWLRoe4jeJSUU1SnDyFDeHhStl53FlOWc4Zyko0nVRdmbdVM/FFUWkvIfM3/gBR
YY5ZlFbVrzZG3QfqJ1orySXc9KJ/ZkPPiDr3lRo/CSzISUFLNQPp2IOeYykQ5u1i
zheHS3YxbK2OOohUkhUPtq6fOjbnetpZ8BwhLfJbU3t8oLX9jpAgdRDPg+edLjn5
u42O/tykyXIQz+ryyDqnxjWTaGD7US1xnoDm/6MAId+y9knG+dKDeedsMlA0z1ig
NRKK8mn4vLG7hYsQJuzOBEdVXRO50qeDvckwq+TFWx7aKKLHZXzrs68NPYz22qzy
a0vxtZSqfBvEqpv4GcfyHZZbCTQiBTMs32tPXxHGtg7bLYpwHUjU3VZ+vxhyPAwB
NMEn6gvfSSmvU7WCr+nq5zssIVNwVVdRfGJVRHRG6RwrWyBU8mwDn7f8weIakMxH
nzqW0D4xbtya5+so3R/nx35GIpYrYYXHJ7x3SBGTWu+g3ZxNqBlOiUbW0DdtoMv1
Itoxss9tONiFgUGE6vQFxqBico6FQv0uWh1vqVlATxmCP1hIfT8INgGOuozFQE91
xRen4ZKUM2FgWMoPvmUznblo3d4hvWpHeALorFjb/T3wcjYVJyz/g7OyO4AbalZx
KP3O/TfzGPKcrlPRnhUu3gWmtjxtevEpUNGJbwaPKD1bEu3i8TDi886vINnJi9gg
UM8zaA9nNIM02ZBYrsj9Xx67sx3qNaMpcktP0WghcrBmRbaBmUZmKD0JuhNG8e1b
Xf7erLGGqO7h5wKhqvmAO+IAu4NA1Z4cf6m9FVFmZGZqKNF+ztTlP2PJhl8bczuI
IBE/9fAKkaIWjISkNGgH/It+1eBOBRlvIHKrbHs6BlorULaeC5xomkBtCbtYw9Ih
gFY1MQrKyFvcP0psGVs8SwExoEnbCtv5+cRnSsLAIY/8kyXp9W7Nsuo57UGajeAd
amRBInrmpA1oG6Ru2tW0+QNcB+UcDJwBsUQjKJeVPTN93FVzSe2RLsuZ5z5Op5r6
ytfJ8b/QGHeT+jBTgdQ+pPml0znJBK8GPVw1nzDKZxzzcobImpqk3N9uX4brgmTq
sxZJcCc8PpKgLcG737yhaEYDQMS4tpTdLn9LbVbBcigafa4bh4tEfER7mOL2XWRh
8U81eBkpVdCOSjiYT4KFawEDkcLY54sOgzXYbki6rwOsY0DyrHEwwWAZPKenBvEB
noIDcp8Wum9BT2THRIuGnUjqXSZG1IlhbN9Hc+JKa2d0LgGjYTqMgmmFn3hzgYV5
hRuUC/SCnHji74PrSZ/1GRTzyt/TSv9cHn1apTgJcz54dXIJU5W7jSLnifZjfE6o
7DqqTeC1Ux0Pvzn14jRPez3xsWn95+HKRSF8sjN3FWQem/qHX9U0M1slXgxBPmwq
a7B962uDdmcchMz9dkXkZQVLx1/6tE8UNDJlnILYgN888cStHW8EMI1diCQhiVbE
OC0m80IWdjYl5x9sVnBZ8PUulKJqUhH3YajgrXUnpscGplh7k32dP85CQd+AleUi
p3PV8KTWSSbK9TkTU9Weh22kgM7LhPvMNPu5LaUuN1cvdqvlD8C/sD0bgq89nSF+
GUjOA7b8gy6qOqmVYJLV5YQrvs70+944Kv6G5Ie2YbhPvIAgPLT6CnHtGJVw5BtL
lVHgm/bmLG1E618h59vzZnN7RMRqev/GHoUaj9BJiNvAcOMUBz6B/74Vd5De03+j
voNL8GSfbfOZWrJ2Wbp2a2AQu7UMafku+e7NtnVHFBr9knA2k4o8Ovhddm17Bu8W
KPAIk9+EWmRns/iFiuiUlxRVVdRWx5ZpHgrlFryOLt5D8S5UiV/asujG3Kua8W88
mxRFAN+02zbE0amlI+6aPNr7crFHhKld3HpdipgEBD2u+cPaeTu8c7XoMtkLLTKW
FG7R6bM/CLK67MpVqqOT+dhsoyCSsNm6OASXmEeQTHl2YAVgkh4ADpys1viY8ycI
MNMU0/Mn2o9ArdEIifb5IGsj+9GXk18t6wAye2FbUJPlY31tpic6RqQkSCgAULxa
mIuayVeJlmI3ZAoHy9z6ypW1vq8iPKx03AY/ziqacagvc+2gJlN8VydxYBZJoDcR
ZPPLPtslgxuf2tsI3ZdWS5CL8Y71dKXvrJItbolNm+r2Xw9RlT7qC23c5dxI+BYJ
e+eg9Wy0tCq6YIvdlU2lqWbg8iDRJfiQtLUzObquAz8id6Swr4q5D9OAOrVbmkpk
/5p/0dpQW1xKwsuijVugGLXphePR1cKQZHoCOReGGoBVAiMWk+Eb9UfrKuXfuStq
abseW1JlO52Qxs6sNPttWwnchu0oZNKFH65cmK70d+Il6KbbiO8ZKB2x/ejEOOGQ
A3RtYywgo/cRBI7i5mimeGCJLLEe+bnS+A8LbB78FRw3R/mRfj+aFRxc5g/3U0tR
dtxHDaPpumPrd5RNdtjVF7dsx1bWfWR+Nd/aCFiTKEHxhrRi1rTipf/WWVsUyWkq
MTjwgzShJVXYFvRTGotxXvhPOhcoY+W/q6hNR6PUJuAx0eUtWt0F+BSYCIWs1tuT
oQe1cjLZD1QZ5/UAd9nVULClICr1DxlHbBPqsvmr0K31Idbvw1GGZShAnz/DCZrq
qnlnXS3WB9EBtoiwBnCF6hp9w8cw23BdCG+4gdvFopE/kd58N50fycU/K20Gni7d
F5KXZOTTDshSJgHhrpcPO4vl3TBL0DEUI4J8AFq+Djmk+a8svc7B29aam353MMqE
vxoazNMSCYpRnYXXyxG/OwSIMhjWKAvBMLmcaddz4FfKhtsk7IOaoc91QIhojsnV
VMN2ofMhro6FW1RiAeWR6p34Y8MZ/r/roUyrvJn6Hyqard2F+/9K+fAtwhnksydF
WWFduhcQtJeiaSMa2wHGu/7pIhjAYy1MEtfGaUYsOeSbygKDbyi5ofuvFE+7kdza
Rf+Q2xOmixMNQnjFKQdkRZq9XIPrshAmuezp5JcLCw9tos5hhFw4qIYiNwNNd2c/
+u4BQ+V4cE0OHU77msf7xQV7IvK3khCkwNzT5M0FonKzS2534iR3XK8iaI3UIqcU
NZLQYNy9EP3vlEL/ce0dRa9VhSU2sIBbG7+YbGWXUO7ZiMiqviCl5UjYfrk2mM9p
89h0h/CcoJfmFI9+0mZEXUI5j6ArtTCM9ZUxY1hfq/pBRUTTjGV1V6ow+RKx4ZSY
/0wV55t5/a6hBsaZt148kOQHQRkLNb9DoUt6gfCTv6vE9s/vXWQec4A1T3RXuI7Q
ezYXISrjrSYXxViKw+bWY+tpQx+iWBFch4BxR9LxWlDQygYLPbi8vG8QttcpNzlI
aQsUAdAfb4aQBSon+NoCDL1Y2Cw/GbvIbJpGJFWb4KyO0YDYx+YyG1L+Fex7e/iq
PrIQ07FP2QKnGJGn1yDJ/tPxFmAgki/0JoVbxmMnyskxZijkslmcDZvplpHu5+Rn
Wh5Ra93+UbWvPmQQZpWz8htOAVlV6f7bgzA0CAL90Y9ZFmDqK1H/sqBiGXYDATbE
SI4IpRMRgoMJbIyyZ6B2tiP8kab/v2CnDQm41keKU6yUfMbW0vz1VyPg3kLJR2BP
JZ1ySLgjDc9SnkDwgbhJBdCQWvL1Jd+xkXp6tF+nRkNh78M9WW2+Tk3pHzkhHUdW
Axab/ki5DezXKtpBvqZ4Axurstv92oELjEBmt3RvfQJ+zSy6e0P3g+he6msGrTzZ
3Vdk7tgezLyqMNzTf45Hz6SUOT/Ph26ymgqZldIiBYlmaKVz1+ujLWj5qh52Ej5q
WvHY5Cpjjdziq5lZUxZB/JChPnWz5RcUu0p9md43+8DHkTvEOpPGhpWDC5kU8O/q
uKtS5bCV+TlTF0PfkGSqfPmQn7OpBNUhsprjWka1xjo7saVrqRfevjRz1X+DPpGF
b21x0tTYZZFqeWYSVhiHirN/v7+7Q8QfXS7cKkOqkst+ll5BiY1UZ65eHiBL+sPG
nTlpwWpq5VInsW+D8TTCEX56hDfPOtwJzXZuoKpkzUsKXw3XdmF4ZiZFUTE1Gb9Z
DahcWg0o6SBZ/Fsk7tF8DCWB4adWCed2TXohoScO6RZebyL9qiuTzyxF5S1sWty1
q1Az3R3xSMthwR2p4jNH8jMvAL+122uRN63BK5oy06OPZPhmxuHdOnTecbO/3r45
4C+EqMA0ONrP/1cObtg3lWuj1hD6yEkkNUdNQ1uGDPjRHntWyVGVPtXXkNmkc49y
hXX3D8Z/AAf54+tToqPzZZckaTc2QGm8PCaqqul3E9NwUTyKo9Vxpn4cz0cz2eHY
Msg44KuliNIuM5TK7v/wQG+e7mWY6zVuFKR0n3X3YkB93UXYBBotGw09WoXOVQSb
Ba6GYZBeMd3vuYpusm188ps1X/23T/vNinnVDTb8yGSpCw6q3TVwtYOUzTQSyCBz
8wQVzGtWDFQDgxNX9mjOfghTJlWLbfn+8CQ6MuHo8AciccsrA0jYlSA6so/0r9T6
7l2kwukcViwvbPncMZ7eDCRXivQQc4gdU/AhMeWusWg/k4OsnPe64cJ8YQ5z5Wfa
fy0IrM7lTb0L6Vw6fdHqXNT948gosnwLt5ai/XCMWlSfPtquVfKvUhQTYVmG9TbA
bE4P0drv6O2c+8BDCQyaeDOmSji0113zU0D0mUTN41zv0vATpujDaV+JSruchRNm
vRFdh1mqYgktte03TMGS587KlMO1BZTgwaDSc8nllq09YxQUjl0CQiP4RumZIPLc
2gpFw3nXVowkgnn9xwUqXPrcbqC9OGVxIysSQTBmZaeiDYbZeHsjjMC28mtjp4cf
yCt9pcqpfdGyFjEeM1Vpw/S7SVrkOrXYUhMODhDVs/DeAx/fzHXwrwK7ophTB0NG
4E21DaIDBVFJDj3mqJBxV5U4Y/pxaCfcFBgR8E5FLUVyDdHdfZ07apSfHrtgtrKm
bFKXvKfex8DDxDSEafMrpsz9mRE/CJdpDyu9snaNfG2d+kth3Bwz3c3p/SlhADhs
Zx3U2uF/YQ0bBVnHedPyJtflalxWbKCEYGMQbNRQUFN1t0xEjRtGJDCH3ROP2gmf
dEdiNqbsF1m5qWgVoN4og9TQ9lfWaa5EXxczrgL68nzyDN5B+M0XufJDXW7XMmDb
Z/L+UivTc0s5Op3URGOPmMyXchHRwkGeBhw52J+CBnMddIFoNDs2uE+WXHb4g84k
bFdCUm7Ulq0kbYkAi4Ctz0tDj+t94TWMBitlEkc0z6DmHTT2WwFYCcycSU05dXdz
dsa7ZAUvN9/ftHyOFDUFLenWteZXbufko61tdToru/kzUAUrnZEF/dVa/zNhUwM2
Q9fGc7airpr5XvnKNVH8q4frPycC1IY5GXVBgz6XPFgE1EcfqSYEvwdFu+rkGIof
TE6b+JJo1D69WwXG6GmAFXv1Cjpe+T3sYYbm6U7WKHvNgifceqxJoOnpgWE/refj
k0pph9FknHCrCDhL8nRVYtl9mBqSNpZjH0DhqArFsp69P7XXtUBRLD2wprxSALJ0
XsHr4U3TjXqwM1lyV1w5csocaFFiKhK/WF+5kSLWrZkhUvx2wvVFlqTZnDb0+KnY
N3SkML/NegYEag0pPF64jZTxbbmMkNsOsKz2TZNY5GUvhftbsEokkkDn5IBroWYS
6CS5TMYHV8q0EIwBZp/s+64axHqYTme8CaWfTJ+vowEmPd/mLFzY4ITpvtcE3k3M
xjZakvsvP45InNokN9bpz+MPQESRnbFiXiR++uMIlIv/1CCe+uAuBLXkmH18w6p1
QkMmXYiA4lEnanmSB9R1T5XwJlMF6CMHXDPTP1RURNiCAROEqlxbcJd2V30EJA2r
6KfmIg+S3ipWxVO1QmTvgBjHZvSnnQOyJ1+aR/yJhxsXYo9gY15OKZbucLEFFe6l
l4Ti6cwSsM+bjSFdXIZwJ0V9QGT369G65Pqu2ydAxYROs1fxoyXbyHxsaVG9/Kew
4h8YNPZpVZtnxx03L75o8ltXg/HkepbssJ5O7Q6voPlqAyP85sRq6JMSKQTI1WM9
LQ3oWJoaMopGl8YjH8NM5LlJe+mZY9pcTG6NYwZjXNRSiyx26wEXcnLN6qpCokfJ
0SJ7OLr2sypJWzEP3y39jNvvisG4KbLUk5w7ldKYqr86yVuas+kJp+sYCVLxnVYn
UrqyEwC98BELj8D+1gE8HxBFRjf1o72t/aKmwhxym5Okhw61cPStRiD/hZubesX4
MOAhe2/AznzV8HrnMbWiXdh7F37vTA79AbmfTOztbgBWtDHNGeAUuQDNcXg44w74
5R0brtXkV423fnrajMNWcgRwJ4rBQzlz8TnWasar8N+GiZFexke+yl9r84Z6Ox1p
iAhQs5sstntWvlYehYlYsPpmdouUxOTo5wUG0QuvrH4+nFCYuLqfXl7Gk1KeCsco
1y5QSVoLPvPnEXdZQOePvGlYSqJEOMMr5yFpkwVFrhxd/UQttBaOiIzdt4LN6gvQ
NJ5I1Ak0wgCiG2RzSX3C/JuAlFh8yuNZkFxWlqIAwzaGEl3Q86w+az4ZztF0QCx1
1RO/c9dCgAmCsLQOdbxxrUly7X+3XLz0e890d8A40ozwJoGAYKaMYmxcQEK1tcjx
HDwz348KIAgusZZ1XGK1JTkI50HiD8q0JfZuUlVEsfJYnKRp2lB4fnIc51pPsVPG
3IZ6QLPecrS7GkDR1W8xXeD3Fqq874J5fgadxWpU84fk+96U/LX0dcXIsgR2dcOL
ujENNUSAqW1IH/js8Ye5bfhyPH4SGQDQDoH9Web2CZE0MYDqhOufI3uKl+tYue/R
6zvuGlBSeFKSQZQUU/z1b9ownOQuGZtLiuFxY133bG/yHqh594aDBLCyEfuaznXd
vEaEJYks+ftvb0J2faN+5lFwri7ZR00u5QCORbA6asyN9h/EPHuTkYB2oDYqA2XP
PrD8DZAEqIri3PFVsSVLNykY74ZO73xXzg0kvzEyUuTw3MTD6nXuI1dtf0a8X44D
tqdwnzZXGHyQl1enqoEKFDNEkUgNtjxaDvCC+57tH7oynbGpIVqeU2WgzUFSglxU
YJ5cqhuUoIA2dFru/BL/msfK9Jr1UpTkPr8JQP2Pi8nO73HpRUQKCCSGpSBKqEWW
+n95ZoL0dzG34EprAfFMrR4KrmkrJHzLp1JQogC1/YIHK1wHuiEkgwkdiXFM3lFM
vvuO5QO1972FKn9HOGQC4T7IQZNZCUyCGBsVIHNQsH2aMwERawxdo/8huZa2MddO
JRaDjCgcuEJhVF7MFGXd2li2XhG2YNNhAwZpZLuTytrx1uHrt7JcbOO8ZbN59akd
oCs94AyV0E4VR+0e3yVIM/cS5JZwkjnyqs30iuincVN/adJky18y+vyBcU2L2P7t
egE2IwYM1xwse/3PS/q4U7AcdcZqvffpibcmVHijrkPsXC09t7r3ql0rvq+UBWw9
Nvf1beaCJk1wZP0h9juTWjbO3wfJCaQpUCwwXcPaq6qis+fYOL1FH5L4YupeT8Sw
Vhfu4mQx+wE9ZpKaBXIikCrmwdEqSXPnW+OmD22OyicT/Nu5gRmG+028qH/70ibo
wSTPEWQtTp+yNcd/TUco+3pP/HSooX5oxRGaQlexPuYpLeuSP5WT/lpR2lSfe7n/
KO0W/7IhMUI5I2qRzmV2dlk1RHxYJvnWeQAqomNAxNr+nIoT7iF2+ujlSMNCPp12
I4Knwgm84O15cc7ybGkms6d+YgjwjVJa9H0Edl2oMDrdZ1qAmhFKDXcWvMHMPM6r
Aegmfd/v0NXVs+B9h+HErk3OQInwzABKq04Zvg7p/5nOkg/WnvOY5esX8XYGdWyY
BqQNprsSK4NXFiP5asWYOQZWWMPJeVaumq7MZEytE2UHQzoc4E1AvAjuUm2CrZwv
ZUIHijvQfERZYBPjqvHx/c2tvatzwkupJYtfFl97kDazvExP5pdnaA9G+a2+bRFj
NrOgq+pfrFr3+3MU8tj34MKSZE5SWO+P3aUNixMq8TpXq2AWnDxv6Uwm6Qb8/XOD
EnbNZbVUPZR6qTNRk9moWlCSmvvxwRFXLQKmui/XF6X1j4lNXopw7u7PaOBvgFyc
ewKqWtOJQPNceskXA22BXL+i9v5Ba6ivay8Ff4eB/rIvqwgR4cdaGc6qWWJzEBWM
4iGjAA1lKeUQ8HyNQSmUFufUOY0nGINfeyP48NGikPDp/26gsk0QUMUAoFIf/Txb
//FAGO22qr49uK42gExlybWYR46S75BjO9BNxFiLV/tEdND30W4caAGwK2BIMdCA
VqGnzDdtX6BlmxMan9xFvRPFNEc1aH8Rpq/F4V7zcIJ/qiKuFsj587vYq5ZXsEgo
XgFYrYc7n1/NjFxcyleaiwzY/BxokZZnVtJd6HTycgMYSPs0VfLDt0ckSA4xOFTw
l6BLMA483ZC8zTiYDFYOQDUp/3gWfe2krDy0mGOQc5+1+b0b6ahnStJqPiV9oGIU
X3zPLKdD6L22LLB3bloq/2zexhePjUrQSfqa7gj2BcIGDU7HgFvAwwelfvTOdHSK
EcpMtsJuoFjn+g6UTRgyDjLLd0PD58tiBrg/zXLrEPnQHfxXv845QTxlTPB99/yB
nImnfQsw5NyKjrnlpE8dc7prhB+YqXYrRV9ySdlm4mc53nxZaTEuaS4sqMc+NcCP
gCvDM9QfglSrfPymp853Xw==
`protect END_PROTECTED
