`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
etcMMilJfFIsE+et1aeJcslO3GSHtk3MV5xyqC4XC0EkM4RbgSHSZ/aX22YIGq1o
HJ5N6/1NhA9mLCKN4keQ8Bz5o6VklYAIRVEj+TKvsfsC4rQ7zlmSO8WsugEUJp8x
wvWb50tYyyQixZJ2zd3KyCV6Or4IfBCWAJqs35L0y6+trqH6IuPlFQLfUeMhIewV
rmRiPD6WRVSYngLmB4tugp0oG87WrOFWhHExkVpyOJv3K7bPcm3cKLoHd5SBCwuQ
n89pL+hNq12sft5VQQH4ZimUIOxPP2TjgTK70CkpuPEiG/kOgK/hxsBktoOvqbqF
u66yu9WWp4kB+f4fF/QoivYSJoHaNuy33W7I7YRWfH9vMDRSpN5UJyZ/3El32odW
OH7Jim7jv7RZBx5m77OAQaYkhqnEWZea4sIghW1oe+g82g5sgfW6sFa2eN1018aZ
D8L8W0W2V2Kt+Mabp0MoOw87OdcC1SgTcNbwaTpMfnzaAc1b/sQ9C2ucrFRTMOVq
flw5Uyffr1A8bDvbil+tIPuRSvvxFlsUqOqlo97E8gGjB7tz9tttvQzSHkRHqB1+
pwzly723vEU2J4vWkYVPje9w5Hf3pv9h/dc3m6dR+ny++SvSHdiKqJkDnWbTkjLO
D20ilmag4L7caSom6Zd6uXTE2ZtZukW+XT/XDPi4IcX2w5j57X7GY0ywW3E488Fc
`protect END_PROTECTED
