`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bc+LgI2KWGen2Tnd4y/IYlssTvJ1LLezuixaX1oHFm7mtXt4NC5RUeiRzUWjyiQ3
qVazEMH3xZ4iUi7KmSffQ7ZrsRAayc6b6iMQnkDjR6L1049HXx7FeG4Cz6JUFR5r
O2WencwAKMOp47rOY2PWq0MqcVGmFHIiBOXWO/xBMYpAj2WpPums8Gzi4MFwNFtc
8xb8e6DyImgTN5Jqqw1ESNgOw+4XOkMf/xzH+GyiddMjZXNyMVm7Oa5CCJAEWujE
ITDOiG7kH6nbB9w/mrTKxtyUOlCw94gQtXxQyINSgFmha2vz1cScn7KEH1NqNFw5
0w2GyKC/YEXrm+xH5qXmUB7mR5JYbA8Ion3sX13FOAN8aKU7JnAWOSrFqRKloewJ
HiM4Z23eyHZkqD4dNssYG5Jrkr+K5N6RxPVbs+j/34DlTdcH9UGxjMrTIQGxrl6K
`protect END_PROTECTED
