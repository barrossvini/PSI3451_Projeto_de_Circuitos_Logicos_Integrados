`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Phtu1taxtYH+T+EIvyTnCOBXiMoe5jpbRY0Thp8tLhRtkmhtRK3pcF9fcb64qYFJ
PRlHJgvUi5U83NpVQU8s9SYIHZceUyosKD3Q1r4gxEXwWnOj0ncDFA1EVve9hT9J
XhuG27Ig946dlkvkcC2sXvBhT3X9GOcIUm+c/pg45wr/4+MKi6QYxPeWD6D01EoC
9ohx6tm4pnOxnorpSI4AGytd4Kkm1ym90VnHXIRw1Fs3Xi2Y27tAS2gpVdpWFHx3
HehaZxnCMs4d7W9k10yPsNloNJEpL+tFvesxWZvgEJ4aB1l78as5sWc3447lROoB
1U61ON6gTG+vPFQaey/HhLZAyAiKyKFkwEcYQ2fCoCfjJITI1Cd52zIXZtPRtKAz
B/aFRDH6Z88nRttGlfbmO1aUg2zISKY4VaFksC+YUjXcdUobyKZCt9wS+bo1S2xO
1TOlC+6+VWagVYQ+pVgSt8vMy7TvEvK/nEpM8asiEsSlIoL8X0za+ViKsGuMRKXb
epfaNqHavLNQYFRNf0Zr6gyJ2GY4wXX4bKfpW9zD4juma6F7tvCVemfLYGNQQ8f4
PJ24lJdrMvxZxw2ZnI/aUqIYhAxv3szyYkSO/zKu2jhJV+j/+wc7MQ2CoQiEumj2
LYXPYC8LDTkRa2+yPalD9PksZCdnsqsZUR2PPPDz7etpSuCOf1ZmSVi8i5JLOYq4
CmsuKEptsur7+GRGVdytMqziG2TVBR0pcQhOiSc0bWAFkufdfwYYWIs8FZok4vy1
MBWID+Flpa4Nx1lmIIeWBYfxpz8cjengCkMvE3RNWn3z8op7ebgD2TnEWFVRhKug
NJx69UYBW2KJtJ49fVgkQA3BV1aSbBYBkzpliqO/ZPeiRN7PNfjiqmjhp7K6AJ6O
Gm9/hLHiWsXgD3EsG7M1QyBDVL+Rsojl9/9DHWzlhG4KCkGdfixHMruPMBMjC6EJ
QsLfSXAA7h2sjQQM43lND7EOttFpaMPoJYHf57hXRzgUBXu8hjcERixjYAyxvy5c
LIFSab+VsobfdsjPOFHzyg==
`protect END_PROTECTED
