`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lGHYtGHb0+aSV7lbHvXshU2c8d5NzPElPYnsG9RnKhjxw3C4dIUYEO0JGqWjJ/lK
zML68YMMf5qUjDa8peKU4JuaiSXCpJOrzBf9bvjefVuj9NwFieVxbOQVzL/JxYQO
uQFt81kO953gr28r7RGnVPevtj71jS+Ai76FiyrDA90YFUnEh4ZH1KXZDJ9+0ZwM
HaRLH1T8vhtyegc8bQYpiWDld5XFVVZZYfQ8HRJ7gyIIOI2a3nn1eC+BcYQXFYjE
eL3Pn/iymzlmX+gldfwH8AUJ4P870KGt9xhdi85mkbqHG+aT32ymsE8esNxgwj/J
Wi0HR4DKtGfYC0W4OhwKbsyx9/UiSapihPX9dbv5zDKvH5WRYp/nbGkKLubVq3vs
/jz7TwrVb7hPrmrYgweqlBxoEA/E6SrfikrvGQHep8EBrrvwGiP3RR0O/cmWLwFx
LCMJq4JJUNt3uM4MK6oYwntSsgBjwD1n/RmYM4DhUkn27zAKDnsuvGfxuBM45fb6
yI69RwXO0M3BaIYCKTWarrxlHwvXYhxUAueK6nah4EjlG7tuugmpqOrDDjHrRYD2
UewKYPqVKyUO4YD6kwEbM4NA+8XonngNhlORGcG9Y1j1TChGWvpuFvfPpZof+1AN
vdVoasgfmE8WSOEgXfhxKgnStcqjxMRwOHWVPjcVW9PqQ7XBvnmGKvtVUrkv/1PX
Bu08qr0gn48A6QAYDxYeN128AJF9lFKJfdLnrC6MBlwA5bP7y+y9CeTbNEF705pZ
l97y/MeFsbSh7+9JN8gJwRWrlWerc/JO42W48Jb6eoE7vVPiG1t0JwF6QBMiTfJU
uUp6zzEnicLWwseB9gT1Y6+fkVzzRrJOZwlr/BTYjO0rpeVovcBNsBBF/XHvqY78
Ga3kLe1cRZqcgb0r6gg+vYeeT2/EBPSAEnWkcG/Rg6fcC3vxeMRhbsM3/kjdRjMb
kVzaK0K55JvUOe6O9RbQyaRBN1AZn4NQSzn79usKX/lWhvPcbHJMt3sCHmm4mCws
z+zhem8/VLHBjD2EQmSALCCaYKqSk1riXuDkZaAka+Iz0STlsAymz+3dzuNXNI0r
ZaL7z6hX8NhHDJ/e7lMQcH+6s/i7+hGCqCU9KUD/SCIWAWEdxu78s64hZCDlmnnF
3cQccf5/KeDivE37lnhTwyaOYwGE6keXJHtWu1paTsnciuma/3GbT96whv/nNwBS
9jZrTuybntM8iQEEoKr2Yq+IbtLyb1Y3u8/ijQh+q7PxXQtN5nNKOwa/XoPY6Qcg
`protect END_PROTECTED
