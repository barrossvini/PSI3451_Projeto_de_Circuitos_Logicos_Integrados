`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7BnP6vPE8dllbJ1eK54n2QWk4CEXfXidne/tU22Usqy0Zg7BisKV2+191Iyq/TwM
Sqiy3RDYDKBysG3VStxrIRyKumdZTK99JiRE1CeiL6HKkzjKk1gEu5eAS+oen5QD
qBlpCP+Olsrl+PGzNQd8JG4v/dORhxfmuN7RTkAeItYRwqeiJDBHe95VkExQIJNy
naWsYv2hKyRpABFM29viZju/NY3EztrTD8kVPUFWtg45RGWCAVqvJQHi2W+/lJbL
tmFV5CTWwusCSAjP8rpRMB1GKZF8X5UH6kVuFrTXN+tZXu+Tep90DnWQcOIvGApb
d6P/nrSalq4A6J7sPe91jKiLAzmJa6DW8L5i0telPd032hIJNhFfm4Be76UFJ3jc
+LssDczbyVBahYTauEu4wIcdXS3TtHY6iRUARPzRdHAyR+3auamKiaf3wdQWcBG0
EvTVg2iMLW7nQwnQlM94L3mczMxKoM46TpIwwzlS6+SvU9SK5Fl3EtGefhWefOk5
ZtDBQXb70oskiuRWcTLD+xQgFCs0be0iNRChQzp8J8M9s46s9sXUmN5tu5a2UCZY
/PtbJ/Xy4Y6849CJUjJxNMxW5cHTgy8jZ8nj+OlnpF+CNRVDiVkkcf/YbbOBISH/
Ts6DmkbEthsWSXfwPAD/Wfd1Dmp5+h1usFByGH3fgEgx6vRmfhYOP83vRfhHmZv9
Q5+YG+4o4+Kj8fVxqdL2inTE1UniFIjoYuLHUTg5E1EcgO5mEnypzMMj5JOT+cA+
5fKdCjM5hOj3RYcRlo4vjyJSuZzc7AHNCOkzduTrLPxAK6kQWpedzJNHS3VRpNUb
3GnksMGUriY12Q+QPN0ebk/+MVrJhdBi8A3QSrAQR5IKBqF8cGmiijgxh8So7XNu
3+eoXiVF9uLrk1pI7O+nkfoXeVeDZgm8jeTbwc36rqZ/s3zCqB6zqIuo6kFuzmEX
F2KeTLDf3125FAl2n92ZyO6C2+EsgEAf4lfrxRF8rC8GuCxN3DL8/85PBAkDT5Yo
Inv8FoGYaM0zUf07AAlcD9Yj9BxUokem4VfQeiYUzgs8bgfAYmohrBh0/veW9bvx
g7H+E7sp0L8V4pMQMMZ1TITXQ+dSxAndhG2iMJJDl7vhFiBAQQbvT9FzF7qi9SvC
nkWn7rzgx1D1dC+w3OSXnorFUVZwDtDiQpiHd5aVIJCpoIsqJZuWRD9snWr62TO+
odmRb5JCVqkobVHLa3J4HD7G/7mHT3vBfOfCz4JwD6V2XhDplA35Zq34Ax321/Bd
NsNZ7I/J/1lDt8R0cGDjLwIOWtlPEMnoRUuTJ6ZmU9nWxQ/1NE2sGPIheijmfDnE
l86J8hDTkg8zVF2VatbP3vtPridFstGmQwzCyHz8tkBoFgtT1mUMwcS7e/jNpUhB
nlYBgtiAWjWt6thWDQtT+I3Sf/ygbSnz0TM9i3iaq3v0RLvh+NXHgcieLH2ULC24
WdYtryyN25fkmNzoxgDT8ejI7Bkz8dV+kPE2uQ2osix+tg9zokggL7uZ3q1RBwer
fXaYh+lk1bsi8zQ8MzSTfe0FZ2ndko9Hctir19DhquIy9oCq62vyLStS281fF+tk
/DPOURnqVWchU9YZaszTt8/UIP6OQ3n88FzMbv6Jc3WUnqQskagj1cHpQgpFN26B
M55cNVqE4fVArn2xR4yub28zHErXpVe3dOPX5V2cxsBxLU2Bm59Q6b4f717I74C3
iiFA25W+WO3PYgLHmnHvX144Yk+pgN1NPSEdkf8/uHYgIwPntGMwL62j+F0foWad
S8EAIN+tQEtxvOvYiXBVqYBNTV02aL+RWKw8LwSbwBxwgbZ8mcoEoH3XlepxiG3E
zmA7WuZ6075+svlHiSbJxH/zmI2eByyyNdR71FEU/6MSzmhYEUX9MoTdyb3IPPM9
IedTYYFHbjC98nInhEmqanPA4IxP1NsQWv7WK1oYGz02NEu/pHtHJBWTcZkyiki2
QvwOGRCvZWa6yDgEAikptUfNDbOoRBgz621F9CKx0CwWa+TtEHCgYV5fw+OFhwux
Y+cYURPvt0vpdL51qzU5ETfhMo6QvcNIrSap8tIovyPa07S4qtORiegpG/BlPT12
6aDC4V+yS5cfmTfRfmrbInA+Yrt4QqIDJ0DMlc7MdSn6JYoLvMVRkv06KAKZAdpQ
hfC04lzdNxoyZ6LwUnQebj+LzA+Ch7cno2x35kPNCfPWRxdKbsfC+AUfqmELfyOX
D448ZjkAgNi3r0b0KnvJlgOCy75aGJXB2epNDGMNnTZWKa8QFHl/bP3nCLYy1F/h
UT32Tun0Cvqaleb3jwhZ7sGQLmXAlAenillKlCf+c71QZi+hJUIMc144KZvrcWza
Y2Rr972fdLLes3nRcqM/Tx1Je7OZpy7S7KTp2k7fpQ9Z0u417PhtiBREqee9bomx
h5Uynv/zDlo/EFrDO3t6Lzigwr6aQL+AIDo0bxzNWoxus7KLyYBmpHbqdahc3LGU
k0cBWLeMB/rswyWnUIjljiIpiPnE6Nl1fevDWCRLRgpho8UGFFhEsAe3N2S0HeAl
2orAOIN2VcI2pQschq7XFS55I1iYZlU+p6Cj/dFXIl7feJCf88b/o0sieWozOKWE
Tr41UjsDVA+8LELNNoimrandgJCvGlKx45QTcjt2drD3lUEXQwUKgdbmbJP1e9pp
taouCeoFvVVa1J4/RXy9OVbj3OVAFv42OzmqAIAC8y+/rYb4G7bhkgsefZ5r/FwB
qOfkkK1kHR9S0J0hq7nWjJeLwcI3BGRuq5zPMx0PX+NVFgzc+SUqRzeTZr+Pog47
F2YqcPiloUUhXecU5UC48CZtoDO0a96/9D+yyxcQEq5KnB8NhBCK5Rr8RI1QEPOP
DJnEvmCqQyjaBLyFJHJG0kRxcA4UkUGRnJVhCKNuIGzZ2KFyYH2K7PkQQpcqCnWf
QRdhnZqSJEfH76NkJ2iFmb7J0G72LHMNQIfYVR7xAcNyjwmDvdVzxGvuZORmOBuQ
u0YTyANJHz7m9yF4m/qQtRvbuEy50CXDPQAbZSvZZY4rveDguT3vNogZjb6d5QWd
2Uw6V4OW6KziyCFnup6ZthygWxBvsTIKxPj8B98pEfAxuRjzXuY3DertLM1r49Us
LI++tq+b8R6MbwWpoHUf1GbzM9eBY5i50IMMglAtsJEk1JObgg8fD+Q5T7xDLaQa
tZRN7xfMa5Cw1/Q9OZ3JvGnCNTdk5tPgVc0G1hSIXmPhnnzIhmmk4a49yOmA2R3j
BRM1Es+ZVwDRtmQxhMkwsYdzhdIgYeYK+zoIt51AAFqy1DX2+LDvmijMf8r7lP3y
wA+A70zIo6pRxkevAieEBoNRXAEwzt4AeYOVYqKQfliFofpml/6LavCp0wVl7V4/
gWl6JiOtVKi1poeyoOwDUVGY90/YkgeQXLKoX+2Fa+phhHpmKeN3f4RUex7tm8uB
lUwgNv4KYsGIJHlmY1z+RevedHGUU8cokOpM/VDemH7gq1u/e9WlQBImkRsI4zXR
tKxv04rPDz8JDdeIg4W3qpwSLbE9FjOhiXHoohscGrQ0iYS06mQeZD6vb5Onr626
P3Bo1UsSAFzsD7l3kacQ8JzON+uBzkoGNLHRMb4CHnoUZn7zM5Ft1PxMi+VsTTMp
4vLvWTPs+ZNA0xcnYq5xY1d32FhscwwvfUHUs1CUNBz4UTILHEpuw9jg8RHjHEf5
G0rKHZ5vE1HmeBszUcTJBbvyMtAQHfRiKIrKF2+DzkxIva5NBIerdrj/eIJdUAJI
UFsmfgeQPGir/urlF2Q4oNCTjjpurYm31CaoepNw9dMYfePXyHkWb10ZYOccYknq
+UzBzf+9IW0k/1yNHuO2DvICkWzVpjPG6fnDtFnEH3Y6aQmzvxNTHIgLyhsrB5Nz
dp9wg9sJYp6oNm/G12HUJPcFnr817PeLJfVEFtcLZ0xBIXP7BvYVHPIuenCwCTxw
PNMlhbOKAZC96J/Adgnk9jFE5SECKuYxzENO54gaJIMdN0EX8/AWtVnGPu8gMMCh
POccqxlkXKXAsffPHbAy/+6ZtOc3P0ggd7BNsP/pcfdL2HLVHwY3OAl77VtQqjpD
xeewb7i2Zg+ZASM9SV/hOfKzucm284t1kmNQAX/KRm+DViyXVPRyarmt70PAiTUO
jcJ87iSH8LSP3kQir/oJTr7SuQnc1PqHh4wXW7yf3fQjy9x/xffJk2bJ0XRe+PHc
uHV2eXbwnOeg8kbb+UrpZ+QrhSTqxuZsw+VhxhB3sv23eMbDDTpUVbUIkVVMwqmu
c6ngm1GMEMRIJB+tPTWh7Q0qnrQASzB/5rprL2jmEyTpJkBkUyK8AvGh2q6Cv5T9
1vGPZ1ojc/65FR9+cP0W3P1VCxrpARLPn0rip2SaZXcf0Vqhqz/fOvt/GO19Ldye
/Wh5J49fnv7MRoyvUTDUeu3xeo2lS9jvuRFL5YrJz1BDuewPh5rIodFbyki9VAyA
p8Dbka9y6MpyKvnYydqWzSaXCyF7yQk8z6s3I72iwQjPczEm09h6eUtCSsQdcTAn
LoYahjaocfp5Eq93hSrNQn4b1BOJTutb9Tb4ANPFabHQWlqRO5Jp1BNbMjEFf7ar
m7MnEji9ATMzFFX4+dJ8IaO/+RN9DYQHR9ONt6kPeOc/Z+K1vYNpSJ1cDcnYjL6c
VxvG6TUxeY3hN5LlIyxIdfzPvw37rjMw78lQj6CPqmzAqRMEOvhc3fvrxPzjFsti
dEGlrkUZ7BJnMLfcs2CjLDLiHBO2E/dYLCPp3GQUv32WXRPhRdTjyUmk46UMO4yj
KtPJaSMiFLiOOGuwwaVWr7+n9u/CWGDAOeQmuVB37AlHNXiSNn7N6Md/4uez4RS/
ZBvG/1VE2QychYejqMWcvnsaUsg3b4MCtz16VUAvsCVNSc0J0w1i7QNQkKOlgbOa
aP5AbImsIY7WLvvh/vRoATUTdeq/Z8dYwTNoroE+iptUQs6RvnB9pmluz2cv8Qt7
DVRBkIdua28n6My1E2TI9xzsKDbMjlvu3jyEuB+jlbbF0cQzaCUq7Sq8URBJ2mmZ
haz5XhYHI/jF8jrl5ktIlLipZhlXhKS3uDKMUCeIWEZRY67eZ1TdwWm8rCwqXMKy
L4VPJgzaEhEgjvzD1vCgSu8bVr8zQEf1iNIeqWbDVNxhPhyU+0G9Kd0P3pzeMSxP
PqbtA/tixajRsWHveTeHGQOdj+t3OQpBN0IyMzvqgam1Lh7ZEpCt10aHktMqLesv
+NyJA+net29Zgx4eLAfsUE2sJ404WjeJL2rbrvdvKeY2th6mKR8kUDG3MZdzaPdr
`protect END_PROTECTED
