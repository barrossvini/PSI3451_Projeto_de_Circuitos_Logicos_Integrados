`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zNOhAQtHgnVzV/ZcT/GvP2Sws55s/EoJKf03omCtWCeOy93PK63AkSI8w2B5Rany
nv+8z9t86PXIJ3aHpBX2xe8/GHrsgr01/Iu+DpeoLF2Zpo/ZVowrLSNopr3mAxNG
QcWMTlCcRPswqE82nhSf6AJx1EOGACil0nwzkemFm6LOelV8aKbPCBzpRmVTBpEy
e+Pbyca8wnzfN4uobOK9ltOZm6FUKTcS2Lj1z8snwC/dCFalXxVSoAbVX3iyAgI3
62sGRkhitsjaZu0UO9rjaGVxZYQ5TI/4N67MywVVUVm8O566F0wBAhybWr/uEPo9
n7dd01HhFKpD/49N1xDKj2nySxMXpUrov5myzOJdPwEJouWCMIUMqlKpuaoSJl+N
ZsRco47czhAZXAbg09qIAfmYMyVvyBtVkGCSh+pI2Af/Pd0mx7beDl+oBYy953nG
7nhFeG1uHR3pJjsengc5EMK22EF7+UR1N7cK/FtxGnda5fWkF3XayJFwqpcVVkMp
BtjiHb6EtebAOteG6NqrVW29il36LYITkcJL6nSVwUTvqNgwBRIGMOU3HssXTWVV
ZY6uv/5vXsgr32TsC5HV7lc2GPwTYlmsEsAs1StGJZ+lULo9GzNHYt1765aLp2DL
F6xlcF+ZJvEJbf9+58qr/aBifhfdMWfkqlTCCcnZeb2RQ6juma8ciQB01dMArT14
/WQLe6UPAkJlPU/v1JLi8x1mgjgtP7ERYsuU4muIDfX1rMYXW1T4GHmSZ1ISgPpA
oiTajCBK42OVEHlgUHEV8gC8r+xuQKqEwUQ3B1ZeuF+Ae9gOrY71FHoAyAquuW5q
xrevv5tYEQ/sviNFAoKKIdMutol1GvjfBkS+GGeJ8YIx12PrRVzlLLSYUyHMW2OM
lQOR9dP8ng6b/H7ygHdj5fGuUIo6mO7vkuYYbS5QrAlXCT7Gh8QOrn5WNjfa7mCp
DJ3ydWWuWysbtt+02EnR579RwfSYHSWPxlyhDoXtNqtk286urDKN5poYZal8vSSY
WQFTq+X6VEcROUNaFYpbzCf5ZAssK1LEhckIzQrQykI8uKfLNOUQb0hpsx006hSh
Prswetal3l1/Dpl/lZn9rKKmQGt8wOqa/lfV7hK4DA1r+JcCRT22DVSsWYkvkcAa
GM3umbHW2sjl+S0Hr1rnWqYnHCsn3t8hCikEjkZRwy/Wmingx/0EUmy3UTvqyxbN
AUfuO6KRS0/OSxea+cb7qryYy+4vvW6tx6gyW/wfhvlrk3dxYoue0uUnCLICb+uI
Hycl4cryny64ZTr+oH2/CLL8O8j+enGYLDSYHPWh/EVu3C6Rp6GGuaHAP4sr2lu1
sOY1+elpl2i4wH0Q3zZdRYiP2NAHJEKqPCMWlv335oiwGocArpONaf1xElQNCiQK
+bLQaPOdWq28rVShGug022x3hjwbGZYsAu/QBGgzuVn9XarvQcE9S6h5IkHpwEj3
`protect END_PROTECTED
