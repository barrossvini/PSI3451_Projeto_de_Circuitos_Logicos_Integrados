`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDlnf0kSms1fBJP80qvqS4siiWnyXOx9lkBWzRv1O/zQy/eJpv1Slw5P2Zr0icOT
R+LRr9z9ldMxFffOLd+l2zWe/LkbR8v5hG4EB+Rz/D7VmzHIY50jp+e6ozPRbtbR
1q218VUw/QwRmxFa0+OPJdAxaP8BIOMaAZTbwJlJXmGs16AFXPlH9Je3bObpQ0+7
IwDmaozqlVjWMgB6XMRuLVUFZErN5MiPnn12PeBdCf7QHwAJ/3MioSksbUL2GfrT
X3yUw/S5QhGQpzn1YkY3ETBEJhRhAKLarPbzyOiHinH4jjfllEKRTqiytjvLRVDK
26ylSyp8XW9kgQUh+s167J7jvsLXWo2Pc+wsumTcAlehW+jR0zH0xKM6/PVwN9CN
7NQzGiEHoVTfpo7+OWjzg77melsLnWsBHntlZ2lySL1dADEwlB4dXBUo/1VI4TWi
C1chcVc8lkjNLWdiwjVCfnfRtODsw3wiHgxGI70wvQTMeh4b8ub9UuXoT0cOsMUP
f5c43NSddn0pdX74L191B1ZFSpq8iFGQcSNSCtMYFwap5mCNpPh+baG0ALL14oxF
8gYwBnz2tp933sZW1Sk8VgrcufbAjydjMuoFEkqLq93k87p6XG01ohZdM9AEVkBQ
x6REP61NgsXP2IHobaOUDEF5FA6+lk2opOrBAC0Fuarhz2yPaO9Q8pD2s4bhHicQ
wpRj9qG2zq1S1UEuhJ7BlBza542oT36AxsNO8kSD0idEsfVD62TbiT5Swsw0qpIa
4WwR6PR3LDP086L+pyE9EUMO3IHmAcKN5qRItN7Rb2SsUs3JSWuSj9RKLPz1PnEA
G0q+drKojhgCrjiEt19MzUZyxEhw0XeXc/JWgThhPNC+A9NG8f/6tBXr9LodxKNs
EQW90nLpC0y4eLnCDI3fP60tpRIp7SsqWfdRZv0IW5FGLc6SpXjg6b1AYH0ogVpO
IM7IaIujQ66HzO19YqOig0zw+WBwWMLKF2Kyf29+pzl4x1HdbZ9A1AdTH08L6n7W
mNy/5wcNsnq+q7nfqUN138raESM02rp17NlObPSJR22LoHvJdeW0hRLmZIeFoO0c
/iiv3UvCs+Hqd9gKK/V43qLqsUtWWIfVX109iqS+CbU7EcMhM5LU3iZ6toCgqZaQ
OOdEJd+v8K0S90Q50mdEZNa1eeY0nBI8J/OsupklJM7hkfDW7VH5Yq9ePuTNYXBg
mRXfhgTDKKKuuxrMY1eH4OFn1nf4tO1D4HmoEWcFItEgEY57wSiitkh0NpPNIP5Z
`protect END_PROTECTED
