`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lkHtHkNcapk4biunIz/GowtKLGf3CojswG05TZ5fQfk9QYjToT3onsC2RIXbjmbx
eCXsyFOUGBPUCVI2UxZVaS6G/sHyntlcPKqImPFSv47aPcbSeAgqGY0gtu3Zih8M
/bABLJX9MMM2Ee3aJkXrZwuc/fh2kSQMafEgnhXfcXZZcNSAC4kC6wfZ29nJbOfK
7LcAxn2klpSKmIJffGK2xVOto6XZEsJAV+EnWPVmA2PXwAllRS94uB+dNb5RdvfP
XOBdp42H98LFMxo2vIN35nZ96KmoccltW1nRutbwq1mDw7db+Ef0n5O7DvFLVQZS
dS0VAQ4rhzTESwRs6o8WVdApDR2lhsInOgLsZMTBuofcTHIdE853bEPEnvNm3OJb
yLZUAarOA7Q4BIR+qh5CFDMQ+vJlDay8QWWRH2uTmj0rarusX0UIC0M+Pegw/Z0p
2Op5AzgLdFmzI76bi9SMdKvT1PZYQFW6GvwRTa0zFu6uxkLzpMzMIL0XeFERaJCc
xcR2gxdN2Nrk608PEw7JWykoBbzqC/O8L/nrc43VBf0QWIOB7Da985jAJbviFBC2
qtQHmsxes5KFWiJJDEpbnMNzcQ28A7aRA82y3ksBttD8fWuPGqaHAZeM257l56y5
ZJFG3XoKNuqcqvMWTqRPfxowWoaJs92gRRU5ILw/65vDSWLF9Hfysc+AoFiyd6mI
hyPPIDurEFcp03GO74zO7aPSD4FWIJNKRt1EQ02ic1auv3qWfOHx2K0neRUIoYEs
uELpI29DU7HQmdXbnhILzdGWANjMPd4P7K/mUPfFYzv6zDwAr1a0XZVO1FNOU7c7
9jpsYnFXGL65zifxCS8MndmKpJM8Ir29bHzR/VOb4EiiI6RkaWzFV+TGC8JT5jB2
u4PrfFP4ICARHGdf003Dtvk/PMjjXuLyc6GlYnFc667U5aPkrQAH+LSAOFlAz+Vs
bn/kdY07O1j0Dh3bCiUE41o4MIelBWXkVNu/g9TRzxpjsMKT0iuEeVbjr0xvTWzx
MeUrO9ciqbGs3ApG37Xagyt/gklq05nc1Z87P8OBZHJS9Nc1iCpr7kyi+d8DN4XS
YlPngx8s0QZyV8A3zhzfQ6qOzaIRLfjuBriN/IZfYYCkdAJgBPOAvhpdF4hFN3/i
2U+GVC5F12D/wSGWppYS5AszYAo7Ub5d4Px/UIk4QacTcjSibRfSKUlhPbSCNPhE
cvNnBXXhx1rPj0rkVTDqu/gLNzoPa44oxXhq+pYkfKYZyOYgZF23Z6maCqoQ/s9M
u2CBqYEEKJfX3N8lLAoajlyFJavpfIGhe4Fof5Znh34HBzvj5/FzYfP4WMJxfi2A
lHAhjHyYjixYDMpyrBSbgGuciMOpCaEq523+xXgjXvNrEYwPJsr+DuGlNufaH6vy
dQxSp4dyTD2uOlCSxBb5ioqv7pw0Zm0U2zejFdQ8S25hm6u+H0Xf7OZ+z87C1DKo
0uAFB1WAcY28V97V+M8pz3n5L1lmjEf/Un2nyjdu9hsZSRW7JvS1ddTymjnVyeVG
HtViY1ttlpPt5OYGr1zNLgLvqhQSEDCaFIW/k6vl6C40yt2Yp+PnejAD7dItPDrK
vPb7aYdOsCHJZ+96LgjyK0T1hsZWk4v8N3gVKqZaazyPw/bh67d6LRII8zLVzad5
yI+Pph57a9/IFh9O6S47z/IiUG5POZlXTSGrLYx6oa1UGXpp3CaWdLdgC/qC5RHr
`protect END_PROTECTED
