`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
leENbwlWPJlCouR0bCckvOMTCGiwunRZL0bK5Od69zKoTWhyNNhzEdkVn5mrqLoD
4AkscU7SRuiEy9+R3Er7s/usoYVyOIQasd+fxH2yX33KCjAcSleORmkZA4LnVXcJ
PgC8UofE2d4REsrt0EWxZkQQ2X+RVgUQ37VwZQ0GWpKsOpq6SVUG7IeZ+bfY3Z5b
Lo/BuNJn7nvrjfVZqvYfJVbehOa3RmwdsYLkSza03tJlTQO4a4hL6d7nydB0mKLl
88C4szwOpVqMUQ3f0kNtHbEAzR2m5BGUCkzWqa/MDZMRU0RNk0yYSJs7ZaReHGyL
e1zo09wrzwsdsx3qaqKXSIFhoSihbypipzfqYsBQTsoCKNEuTZYgwXfrIRUVSkzF
pVlo0c3mUnItT9yMox44XcbLxIs9E36msdF0SMuUGzKVZ4b2dRNUKhBFy7BpeVRZ
LJ3wprPTEv36zUkquaLed83Gqx7Ie3zb8GQsegmx6gnHNV6zfN2yeMooBXdxhl3k
i5bqAOSGXnInvOy0Clse0WNZbHUaItiS+kv1E0G3kVlUxZqA9cHYG0gAphFY5Srz
3gl0lIB7a6R+TeK0xRLQp48/9Hu1c0/bJs4dFZpAmCXJL18XwTJuNirASfoYZokY
xecZS9qZRtfuGLSbfCr8R/NCb9tGHENW2bBFjRyLe2Hy5EcbWZ2GKOQYVWCnnlo6
5i8FA+2lM+bnWRnDAo69vlEHQDJpcKnPre4/q/wvWmo1har9dDQuJYC300jDvbfT
Pp/qN4ScTAASn/BBfoQotxbeIPLztCW90Xwur0MmX45RbfzAa6RRPh5j8xLDk79C
ALqqPa89FBDppZUcOZhcp6PFymGbM0uFi6ch5FkDCfxEFEKJjRL/Ll2HVHEBdt4m
PwGqEQDTjBZS7p6U4QttY6ZIbrWHDUg4Ftu2p2dLQlrf/rIlpPkPo9p8a5gnOK32
tUJoG5owPlsXi+dtQSj3Foxn+KdG4nPITuaJfoaO8/aLyEsW7nMSaeBdIv6qwKSv
qGA7c3ta3pcusO2mUQ0iobn7iWhlGyKbd1XNtLPc0IQ0qarwiAATrXw5j+vkcBvV
V4y7m6WGTYiu2DLPYWXHMu+EBw3OdFWp8GTuV1Q4OwIaNpgh9AIXlnIeVkrdT5kI
KfGWrOKdyHF6JXxrZIIo/nuAlQXEF8+yP8nz0F4cH8vWFbKS8g3+YwRvuO7KgC2k
XNRJzzsZBRVGvqHp9hMFcfxto4cp95ElsUrM/b7DkAvYk9sqNxn4fjOwvu2sZ6oR
eQ84jbfo8S5y7gUU7xTzN4IoEGbnd570wvODM7Il7RhRdxBh2cSEI/CmS0gCT3VC
Nzqk2ogtzqbtxLel6H6K6w1lm9vtrO2cg1ESaI1vdihZGppxZTqzyXDaAStB+vut
zLgqFPFfpXfSH6vgkxSzPCmT6kCkkbaxIK23FXiScwMmb71dvQIaDltlrtd/OfRJ
NtOSVso1I9nhdFo/LfDlMis4UB96Iad5sqjYd2HwHFLpAONcaS2QBt4RyeD1SQtY
abkz95X00Q8CSSlReehPlthF+KNwahEoYxXVDMYgfaFOuR/kADP/5VUl9jpGDfNM
wfBOCcjGRIcSCOzl9qLjxMVhXPplvWPHhZblznvc+bdI++Dkv+4A9CwtnWK8KrAD
aow81mcq7venKFSJnkkkEXDcxhn99QEfK91Rg2OrBAj7wkxVwy6pSnhJuVeZtx1M
J2IAsamFGTANb/uqfye6A+h9BN2FkVJ+zjslrH4DrrNv51SKlIEi4cz7p0WDfUBd
7YoCT/rjbPJua3ogYnsVAoW24RlF71KkP+q+sBH9C+LCt6d0N3ZZGPtEI29+BQi9
qVa3Shau/FFz2TN3h+20wpws3/DlMq8rSXMByOAJB23qJN1OWY51a/CxpsegwGCw
y53OxNr34WRuPHVeGYVYFhKpB97dqt2bEZSRNfEcgl8sRFzXwZ2ljLiyDdJlu+u6
J4pg4Vd0gi7ytJQKlV6Sgz0ME9W146tnLfDvpaUC4zNjz3tub1lbYDgkgSda+aOM
EOdswxi+tbhQJitHYhhElzDqQWIeAk14P6yLXLJKgK9fFU+9h6uLs7TcFHoCFma9
/TItyK5aPveVlkep7fByNXe/qDgmnj7L/M1wqGth2rQ8gP1nGLQeEP5QmwytdFt5
LCeVEfPjEC0s9a4U1w4oUOCHoLDsJdaaPHg0lOnuyReK9EUvUxB9iMH5Bj7xXeKb
iaV0RyQJ6dSCN8xCLCjRrtf71JrRWDKuG6dopXFqJ2uZV9rsMousoKCPLRPHtezD
2heIRsqx4scqwAKWcajwDTIZcWzdPA5+9DqO/UP5JQ5EtRlEhgIa4Smf6E5VCFTP
VibDFR4hloGtzUyPPDLYks9WdCJwBL5VS5jK6QhFhplfbasI5wisfunjBvHEq4AB
Z06XW0rcJEzTwNWwKMH045XwWHGuZNrq/WVobtHaestPLh6senmewNS+rQLw9RHE
NYjXpBPpLeryKJXyulHGTgQezOSOfIcBNPqiSZrKmEJIXevAivknVkKsd0k4snCr
jFO/QNrBU/hJ1dYIhotNMo4JoDsqe3+7wGuhsi1ARKFHbiiqhJhYRLj+I4OxBc1t
OJvYpLjPNRS9g9U7RSopZ5JWsxS/Rz5i2Xt4bZwq5mNR7Zg8bnr/CITXArA8JsUj
DXx2Rf7Oip9DvQB4FbYdeoswRMnJMcCW2o9iMOzTL8NnhqMIkKLWI4NiQvNysOmL
RmFRdURYeLjGsjbD3C7Q13pDE+Hz3aK/xrkQc9lZpEuhvDTEv6SpvPLDSh2rZqTH
H/1XQDE5IgOF3odQ6ErziLIrQj7XAYNld9RzCkA7bActkrfYT/LcFBM6a8UNvo0s
LQ9Tr80FayJAWIWZ9Jmjh0egjtrvo0SGwptLNSK0/duxKsk1tPRp2xV8XCBJuQ+I
wIiAtxB5g3+QH336zGBFf7OxRqp7qGpBM+w2fyVVXc96CNpDiohQd5TReTJOjqQv
RfBVfO5Kl3lM7BvLjkTckycwmeMT5T3bn0QXNCfUsk4VsYJL0ummqXhc947b/lej
8BgiLduN5rTLTEEITjKKLsdxuNVL35ON9ExUrM8IXhSc62nK0DZMYGjs2biL7Elw
LA/KQFYZt6BcOp6c59Oavy6Bld9VsXC/emtUAkN1pHQyTbfszeHbpHL3GN3hlyf2
ZDmdxrB+fbzTxNt+35QKiPds3RvheGmXDDA2mZvghConUDOrwbihS9XfxgJrwgyX
6KRBI2T4Zt9xIDqRHETlyPJoKPaIl3Lccr7qDGC9hGw1XZ7M0pt+4G9dDFNoHfnj
FCwRP5/zwFCaiMVYOZNKK/2/6Cc8Q6Gej0f3Fg5dHCc7q3v47OcV96WpbQHKOTbG
yW+9923h+JffecpNfyXp9CA/3W0u7kTd6qFxW3s5XUIbRKIjVXHpOHyxBW5ihIp5
lgoxrstQO1QVOsg4rr8yf30vEdKOVdiBCz4Iml54g3ilz4yCjV4X1YSQuFVwk2He
mJE6zBtmnHuLLorqEGyMOiikqc5BH93uX4A8tn+acONlJcTKIIExjIbMWfAWPV33
gFLdN1HpfbsuNN8V+CdPpZF6u87CIPY7eupr1n5k0ijjy+BfBTrUuPLVy/rHYGc7
IDzgHGsCMoogMgMEOLGWNAk2AirXNgzFmqr8aJ6E83qXNlH2j4ejNc4DnFFvzmNQ
8rjLLcDtzqVbiwFXU6hqi/mlddgDDrOpvZoxBTTOtS0o0UfRVVwwq6JZRDj84Tw9
pDbln4op8FcW7Pi3c7dNbc2PiXdKnrPWxOrHfteGjp0/xUqZWz0MCvliHqTxAn40
8h7agt7HPeraba7cjc7HHg4An7lHU7gupjfzrvz+QijKgW1tP5/mJIY+PDlZTlLc
2l/8Zmvc50fqTaxkNem41btQNSSzPXFicEVQSVS2wuO23glYTKhzLaHMnqfRbx35
OqVxCzuwMF+uvb4Ef1BJRZq6FkWIIAodZ0a1sRgJffxWgvFJ4VyqcnZuN0o6d6F7
RrscUyoDF6co0/K8H019GVHr+RHa7r0wrAcCBTa89KkBTpOxTwYBx+8l/Tqokra8
tq47cmtIYrE30dJlx1suPGAVoxzRMpagByQz7AoyoBD6DkDQ5KMx1vnSISXE5bUK
gD+cRfDETl9APirBZtRzcg2f/a6NiRmhkhOYPNMHwlrCLxqiYUsqIzuWO/+cdEu+
CK8kIl/e3fLv9mHT0KHa3MGt5n4Iinfn9LNF6nVCv0TpVYNqjTZ5Aus5G2OVpiFE
DDWxJ7uckh5eVOoVxJkJJ+y3Eyvv477v1B2qOpAhd/zSDE0wWNw3HCKRU39ZXdZp
Ty4LuwJUDdmLkt4G/gZkTf719JjOcqiwQwYS14kAhOwuSQoL0uJZnURs3QTe2ro4
Mf16loXCvRkKbWxjn4oqmUGZDG70rmN82aFE/lHvecae/7+gDbKkdSTlIbEh7wNg
O9IiyFwnDQ668k5E2T1UOW3kCL1Khc8XFC7ElZDRehCG/PMUw22e5E40f8ujYAKp
XO65IsECyLCFqYKnwi/+cQiJcG9z98uqBuXt2YDrdKns/cOv581sYN9X78izp02x
x2XcdztiKxp2D4709KrF3PJ19L12X1EaYOpJBDMWAsLyED0bcyUKdMLzpI2FJhtH
vTSJrDJkuBeX4k/kgQ9zGnfitdBJTl0PAHLYA5wlDYNzeOnmAjno4GHWj/QSwSm3
7SXV6wvBZd0odceCCooZQiIRlHgsWQz8lAelHb6wAGutUwRCqXHqkfeluX2IO6ND
nydvL4ugz26EHIAyHDi49TBcdgYWFg1KYC7BE3QCAGvw3vuM8LR9ecSRXvdYLU8k
X8tmOQDjIrY0rpEo3d/BAIkPrKPgULIFgkG+1elnXN4vMQ1sRiR5xeNNvpF+m9LE
Xjj3VI4+Kt7jkUhjVn7nweodf7SLQhqKgPyuqyOlw+RcnvgMyFBx2/sxX67tYwIM
z9msIP1SfEccAJP9hBJ7h+uYhywXL+WgppZ7q+b2+3HYyv7nBu4onP5GWyNpLGL2
yAbAuAqzFDOrEuShA4OZ3ZtXKqwkF7Fv+OCxXlpPj1upf0WXwcaMXDKNi1Y71w3Q
CyiAHYMEb2c7JF0rPyVHWavbAEFcFAhmA+FN31vrIqThQmihiXnu83vVmgFAMM/j
SW226IcMkMbXtBfAX5ZDtRvAFP3XzyuEwDE41rAP1ys0MD6gEIPwn5hWE/KyVIEg
0EV/XDKpLW6WprMmuA9cXR39urbXq8ZwqiLg6xw5PQKXCEwi3hfQgxf3BdWaVl38
B455wYeFzbFwUrdQ1kBdqtHNaN+UCFc+6+ST664/n7o11r9NhjNG+Tuv9wpOc4Ve
wwuk7R64RJrJxsRDgVRN05LHbzwQJM455nsTVPswAuVMbC8gIO75sllynkm2xLfQ
h65e9ydsahvvB7xzxD5VGaP4yuT8+/oy5Zhzhrc8TEvNrKQQ5fhIqbuRx19vKYPI
ncPjuSke6Ez/dvUyP+G+ba+4bqXpSWauJv1C5bRTDF36iAa/zxqmBmLCEDcZPaUD
fZ5+BGoHlF5qERG9hZf4JZAgsxicm/zfLwAb+MhU6iQ4JD4POOrgHDBNe2XiHHfF
sLcaRg71mR09rrr98qa1esz17GUqs85Y7+PtiPeVbJeY4nv4mngZ9Q4YvNz6qwvb
mo73TQPZsAAxQBkg0nXzTJ3BTgmdN+OUjflclTgJ1FEY9gvFvegKQoG1DtNe4QON
X0u7Il7JHQ2+dc1EKAxME8FDf9FJ9w82atKuFdGkjRx7fWjrG9BLQnQ7UvDbXX4u
J3qqh3nJJQ0cJtsO7Nxr2+GDdKaxeyXheF9/3uSella7oYb757ScZ1+g7OXRaY15
bfKs+7y5jsM9Sk+FBJ32lYa7BQUGRoOaN8rZSlnWHuy4ZWaBdDeVMXs5BBFTyHPR
dlv34tmmG8wzZh0vtdAtKGnpgPEWh4jLhmPvFd4mDy+/j8cbQhsb4qVMgOmF22sG
149gJvhWUqNh+Xhmneutjo6Wy5bNXUQrWI66yHMz5Us8aoaHfDE7fm4ZmmOQ2nyG
wNMnIphs7xG8hHCfi/L4knVUbGlIkbB1Ugfhny4JDx2ZolNQy6x+ruj8rhx0BFNX
W4gu+1Q6MVpe1y0TD//JXfGO2MQaoGKLYWYc8K6oOdbtHZFDWK58IM74xa7Gvcpo
FCV/iJ5WlABf5Rujk5SnCR//8/n/N0t7h7XPIWIXThDasxMQRbvLDg+AZDR/QhaZ
G/QQd+fY/2htoS9qeHHMFGw7DkeDXbjpqUWAJ+c0spWFr3auOVvVFYFRjcXQsGNR
BL3S7+WZ9UKXfpGwFMYqyvkrTcv4mvXX7vf1GSmb3Xe5alBlVarG1WZqoccYDcc7
5AJCoA9Fst8ev1vuhyiansBjo9gBXGTlkXwwdN8y1dPFX1C1vTo+qHA6kfpPJ397
nUyjDjr+T9hUKqaUPBUYPkkskcxpZxuebmgrBdmvwCJzCznUuoEEDNyejwfnk6Xf
Lw9SXCqVwM8X/oJxdAnq/JfuCpOu3l+EWqZU5ulQCAasqugRliTXXoDtv5rHx0QQ
NGFPBr0/gkjSqNgwRAkNcZEtnlLXfnpXQMf8UKeMZaHNhtVSg9Asaek7STyH60sk
61qvDSvGzHhCr85fxH6+h9E+NcVrnZgpI7niDLrKNllE5xVRhssGSL0fGLgeBsk0
0nCRhbClkjLh6IcK8QOHTd0Cb7SFIsevUmcGNnjNFX0xYtppcvTndiSUi4BiJqER
3z4K/fPeuappfUohuu5BuKEcEEnTuA7W6di0MeJ1UKN4DoP+hQ4dcxDjgmSV6Ds/
`protect END_PROTECTED
