`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uLtnjjWBhpS66+kCEwdUDs2jFeH2cNojpMJ/1CMpQhy/kIyhpAiQdEzazdcGgkOO
bPIEG1tq44OmS1Cx5CQzFht0/DDZc5CC5F2H2zP6ErhI0zEAr461H0yla6p8eHJd
4L1kIF4onp4lc5NYXn94NK2l0MnICQeoXu94duIiooiR8Ue6I5197AoL2Ojr2TAr
SgqSiE5+cKRl/3uCffavtyLebrKoK2hmvrbWATjCr7ou5/hRPw4g7iXKg+WV9Y/g
qGRvUQeOYoJr97sOsOAgc2LLFnOx6LvFmCdnWuJnTsT96UQbhY6bSADJ79bSquRW
aTMF6FqgNJa4IZpb2bB7U1cJRjmQ0a5g/hLYMZ7P5t4OvBXKSSMy6qoU6BYVd3hX
IdQwUAh+hJYUgADAWwDfF1p4hoxU65KJYyotnVdZM57rDDDTn7pU6rHNriMlR7/K
7ancn9UteR+DW5tdxOUZls1KqvCArUxAWKkD0G+Bf6HH78KDYU3+71FLlz2u5Gca
+/3kmk8mKI9EjCs11tQnMyy6KJeNt4C9RBptyeW3VhJVJ4QOBIR5RmCvKIXPlLom
EKZN/IAy9HUvwBb5UIzTFjZdTtqInkAhQqvkN0I5/n0gclJjUzzD5mbgnkvvDK5r
9s2Z3i1TGk9R0d/BbzBE0WtWmeCNGr+ww10hGdUOpBRRsA3oxzS1Hop/5L6q/zBN
ebO3+lxpiq3nQNPx3YQqgrDZu9RA6xB4U31pl4CTRfIrdCQQkrmMHQ+EKy2z6pas
YIIdUYGzVxNP+H/AQ2eHnrb2/gt0OZlLw9ivCAI6PbaDXfIof1GNHB+UxouuWDEh
Uuz300PIMpyn2aiwsi83CM/qwb93XgMIZwOaYoq0aM3BAzAgnO/vuOwFf26GRyhh
BDkTTiRxSJi55KHuCwTyWQ9fdoymCHOLV5Zbu5EdYAE=
`protect END_PROTECTED
