`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hN6608+8bK1jspvHvjcLCJpE9Xx9RBwoKBo/teIZ6ed+E7JzWz3vQAz8gDrcdjx2
uYlQdACRcYj9EQ1vteVdzcdAZwnM9vuXlauuaaN5MhhQgzms4EgQALfmOqC+LnoZ
J3cEThNY9oWbQ3wfN7/lcgd8a/hq3LpXvbAtG66/DiilmK9NqqmetLL90A6DC7Xf
9WgJcSicEflTEJZcsBR/qDJf7wSDR8/UUWHw/xHj04zbWi6d0gox0ZVfVriOqYI1
wvXWHFeR8eVBJgKZnp24kgpH+qThcfpRxXbW+pqOrLHfgaDZFFDYiyQWYE3/a7DI
iM9DPYMqqwnI/JNVfQgcOkeSjnmiRG9vLcGYWH1iG3HMMktHe3bTEKpPuUi5loDa
yFy67H3AdyzB2Lwxk57BGn5ggc6xOverJaP0d11hbVSr7kAtYamxyGSR0MUT5nPa
fBnzqONrbeoGl3AY0DEQJ4rf8GadUWWpZ7R9bSi73rMQHg9Fosm7Op2wgMsgt/G7
h7KhAUKu2xSAcrgW+zY0rdwzX0C1Z+JuiU7mrz1LLVahwboEV65jOBVyGQxt76v5
L1bt//8ZpJgUSTxdpfxFFhR+u3Ritn1OVmPvaJnjMDEn8da9S2ObIEEPh2CMiS/2
SD28+fYzgXp5Wq2/HgaL0wDBcWMSNZeeyoaQmk76oaJ4dkWwXeTP+oxXdrtT8hgb
lF3Kbt0xa+suRqNoTP6BcJ1aggf7y3d8a2AqQQ0QIGhbfcuKbwu86jpgTMklVckS
HVeWkqR7lZEK6HptCmYfKhoBK0xBCt+BQOEYBnpg3Btws6IFQiDVM4zKMZIC7i3a
GR/F6xD8svX0F0SJLY61MvOOX/lYJkYN4m9uL+7PE0hdcG7F9RFhtz/WOXN9LwIm
dMyyOwYluyXNIcYehjWr9YtQYbmK7On4s00wYUL2YkcP9Ryg+9WDk4x9rwB4aY7h
QgXc0qg/+S2RqL5CxT1Kz2tPLRJlPp+tR+lLS+wTQ63bDbpIvtueAPkS5ksHAl7I
yG93yWL4RhWUGfyADekLBY+NjP2qC6zDEwhXgT1NyHEuZWqW96uuXpHi4C/0Z3fF
RRYbjfS5Ewz3kmICXSkzCv5AGhNHCTBzg+5EDUGo78ogXxRUBPhTZp7ilVCt5iZy
tQxat3NGLi9EjQ8GMkeBRX7Yd+y6PqFksSLdaBgxAzxSKhXsBMd/MrBj0CfeIyLn
YsLRiaW4LmcbAT/v8lTqrujz0jLnDiEBJ7a6DlM8Y2UVlj/CFSNsrK8XNZoHVxER
TTVlkWxlqrlDo6OtPpDiHPklARDRZHii1/2LKJhvqg0XGqb3jkYCX8G17mpOo/EB
jj/BjWqvDCpxmm04g/I8Kz3N9mtELtJATqUeP4wGFlq3zYThIXZrmremRxDD3Yd5
w86nDdtg3Kz90+a+vPyyn8P+/eAfQzD2OSgQ0gM0smP60xz3gCn7NNIog2A3qGjS
3U67EDVNwb/nRIxVYCvWtZq81YXCJVIlGYo+odhYVudPUF+RBrb1a4YXsllLo9xW
zyot7kijNeNJ2F4ZBakF7oKUEKVrzxI0kfKJeX2VEvXFee6www38SBEVek1vZn5H
ck2IVc85yjH463x4a6Y6oLM55OdFR3H4iQtd3fREizGLtXvlzafLtEAo7Fy0Bt9X
RZ2kfSgJdRzjh9CGKx8f2Mz+seJx+G8YHF0R96jqPJ0nErM/UQbXc75m6CEvPKEB
DujJNJNUbipm6TsWwY3/4l6qPzDbmT6qWuAc+bs8Hb5asmHpGS8tFMheSRmYlbl0
NefWFTf1kvhm+VWRL2NTJjm5YME1e2o9psKSj6CYLFT4cNYUkeWt9rbCNVJZH+P2
I5iJREVMOPWdrCkPfMTReFYoUuATGpuigdE8YEWQPEgB2XmptkLDCbptbwfui1xz
knhW1jIaBd/JSahzm/4yvXyD6g07IEQJc+v6EAgXK/smOERmdHGAUg3HDe0DxpBx
dKBUqJQ3xr0soWpp2tQEWtlGAxfxE2x3QE2opNd0hrowgQ/Yo3pdoQRyhZ1u714g
rhoYrjeP4i490nJYC0vboT/bL5mg2ysMyx8J1KINIyfiFqTy5ZPfseihkQV+UaFC
Pzq8ODc51Tj9VOxnxft11lFBvFoO057Gg/d0K6A/c7vcUntmuNPWtbT0roV8uvzN
P5QezsNfdLYkjpzKm4Q/Ho8TPhN/3vgqnIWba28zLrqc6fWzwxcLpDAaUT5TtJbD
tSwg5nucbs14IOTMSV32Up6IEihqUiui02R3rgUJuqfi+bb52dIw2EfnQkA1zU6M
cycECH14ONjsYnjfZv/wXqIXLuvnJ3T5GiNZ3V/C6MI/48KFmX2IEDSlBFGh4PGK
mKFoAYgJgpjv1scHjl7weyNU0YmfeCU3q9AkCUTamQhOqi9cx8CL81ENz42HaF3c
zaZdkuAytja74JvIypTOrTVJHEeLpjtA2YMkyERHr3vGOvQ5hlbzHqj61rCdeTkx
olulE7dmuM3pvf/lh0QaoNhhctqLL0GvzypJVzPOlg4T+kI0g6a0Bk2T38rZRQMu
77WQ5idK6pEgOyE3wpRKw8/+NEX9Cu5MHFNbEArbbA2u2Xnv+ZihblyTWXIWRAJ6
CPH+Dmj7xAE5EJaPDVi9wMgd12V2H+xMeNxw/cckFxvtQ2VtEnsV+cdQGtZpILQZ
Clf2tVFfQeNqLiv55wSOkXJZv86trMLYu0akA4eZ+u8cSW8OIdWUgr8f0e2RjwY1
1kwpmFDCiYRlW1mrLyyBUgN0qcuisWam4Wq7bRsxS+ZaHLB7PQDmQHIW/GPb9XAe
3QM02sAEeQQZAxNBU6fo4xp4lbPUTlpXGti1dn9VOjixZHuMYNH1qfPBZaWN0CP7
46cziOmItf2Ud3jryx+YJgUKQnCjzFzcGqG/U5uKvpJWaC4hv7p04TApMbXFYAAq
v8kTruE3MK83kN6PzF2iI7oiNCogZLxCZRpSB8nUmaZPJoicSF3IgfSB54L/T9Rt
40AWZ6JxmK28GwDea/Au9NVJK7HFCV2siTjNBiFuf/a25gZmau0PCE1P6iNLmKVj
20DpZXFjA9Y+3b512/cIn/bbcgiqZmrXWDkyMSMlZBWcrDXWkqXEypdNBQ6f1HK3
lObyc+ajapmLM0mf4ETmqk1n+sjrnWEJ2omJKL6uQT4Ci9LKYYGgostuj8zRvP0U
UyBw527RKxbZuI4dRcP+ErTj8FykJkSGAK6i6uLBiBcxScnz6h+z6ifum1tcAnVx
KfjJwCvyPFNbjbJun19eAo+6Xb8rlIvKIrct496VgHb6J6F+R1ATZRYafrcqJgX9
+YK6yI58iZm40P7OP2HK3vkH20Jw1vN6ZSVKW0TJMkFu1i3JxR+8pbeTWqOFZSIQ
y7srqgSYH/xtZkFBx/axqtEpqJPo8X51jP+uHE/bpDnd7ngxQrTbFWGLHbpuTXoL
xHpxfIL6oaKYPLJLOWjJG/ef/97xupVfDXJwZDjnsS0feVNsTldhV/hml8h7+ElD
Gn75gTYFkHHGoAtFEz+JM1Al/9AS8T5tvzmAgW+dntbDGyn5zOpGRNRVO2Rc8xbq
nlRT52xfc3HoqyHKx3scuNr5PbNZWQz6vXwYMeZf0pSpOPZApNqSj7YsGoGy+xGN
StfgIE2mvnuK3HHYPrIkIsyacWevRHLz1HdNvxVajDe51iwf0lw7dy2oZN3tEIob
CZ0bMeKaQGaf9b+2cPuY2lwtjvtZnJHoRuEHRsVy9yME04oFw/6/OHGqm3sRhhGL
YCr9pJ8S58W9fGtrrUqpFHq1PRXXWgE0nytjYdQK0Y0cw77lXgcDSHzHd7PqD9eU
8AjxfYC3m9AKkvZdu/l51TpWzkGxwoWQQCJtKIy5S2ohkqVdpzMT0Kh5Tv3kwXJN
A1G1Cw3i8OXWZnReB4Drye34yVsbuimHh602KY7hmaL2iJ7yZ9SKJoVPMZa+TeiQ
dmzsJX+6causcPTCnUWUFrP27nQlI0BqFPNevwuNQGBpT02gmvn2HlrvzyXjrK5k
M+NnmClHpplqNbaqV6/CCJZfLHgPZpxLFUek1wsGMaYauBA7+GDnbBm8e/ude8AY
qS2j9VaG05cDZMtBx4pqz7c2msAeJq4/VejoyJGfRAMdYJySTPZ/It/uA47dYxbF
9SDZF5oFHd753Ao2rMm3CuKtCs/An0BIw77UFDnROcOD5ArJZCC7UxIuQ+g1VLU9
WdNxci9sr/AKtveRFClPJmIbFN6WQO/hDbqvCT0l4cZ2FjPifuKtOOz1RhDLxGp7
vwLA4zR7YQ9OTszemXVRXkPfZ2KV3PeZFb5+Zmh1nDRFzdlr6yrNgsdAxW/LbVv7
SfkthVBq4feEcXT6cCk62QuhPS2v/4cIgiSUjq7RK/PIZZ3qA7OVz4N58H/ZQTul
PwblarwIY3clREmkg2MsBAiT9FDRpWSe/naZuA90zcYIAc4LTnewMDS7Xe0VJofD
xSjACwm29e8rixQu+QcSNEH2TsgI8RpY1p5yENFq+dO98XKeKrekQGa5n71ucqUB
1eU79+Jyk6zRerIxCJlkfAHSU6YoARn4qtgncFJqFs+JKEbgCSAUDsL2yzCcENgE
OnN889meQbbl6E5PUXZ345IJCzi0nBmfnCCnGfn9hBk5P6R59WML/hwMx4t80NIs
0EjB1norZCu3pUG9uKSL4aHi/3t5n5HuXpaB9q2htz3+eIpv8G+jvnoXv9Oqwd1s
jB/Az2Vbar9HM2WWnTsFvRz0Da4IK6mXC8AvmlwXWANfY4MChTPHZVVPLTAKA0Hh
mf4G4hYlCsU7ML9q0Xq2PYrf4dqYMq+LL0FAFOKxFr/iuoMYmQaZcyvLpO3QxY0+
Af18fp+LamxGOAaK3PYBrr9F6hHg0is/RZuxj4+huUU2UN0aeqBDMwtjtd1juerT
FES6yHjqsMXXgKDhLaEjJuOrvGK863WdVeM0Vl/oKg3KHo2E0YRlb0ZGhYBpLTie
pnVbnSGZmAU+9d4sw+0dmMkhixlvkXf29Patx6AvcbGryW6gd3LEhqUxM39udS8+
h/0r217v7e4+g3paFmsodV5moBkrLcD24oEEv9LVuO2iY84m8Ye2BE2wfOIgkGbM
lHzxAVi6BvZCXBRonqIW6zDJhJvn7c+bVIYD5CP8Phr3SmJTK7dzVFqNT5VymvV2
rDzdlD9ByjGAaYWTSCsSEZuAr1/mT6+fLMSGrUhpp4vvklgc2h3SLzsJ6RvakVzS
pMNDEcjkj8p27NdgwNL01bt6rJC8FUtOrpVQRTqjzf3lX8StzBJ/RTmHwrB/2UQq
AWwvc4LFVwfamq557QOJXjpwr401znXi+x+Y+Y207c77/mn6j4CzDjIqQuECwH1T
moh8wYl781ZhfzrI252aMLCYdCMff9YA2Qo2Fx2+LoS/QVCe5HjmvkWwkr48MOyz
CoftNduUWR142WeNuaMNWQRaQEr0OExeyMtx8U0q2u/TJFH4wAGBojb8yd94fJ84
wmI+5xNrypGG8CZJWCpeYf5EJuTTtpddT+9hJWb8omYQR+28yADYLQi9Lzqo0a5b
sM3pYOo4GxQbgYkXaDPnwr1NcjEjhQrkFIGKOy7RLqmJ5Znfwnm4td4CuuIqJSek
YL2i/sE3tkfoFgbctj3tiB2jk6ta/v+Tw0FyIfOnuLp5QTBVkb+PZRbFdONbnCmu
72lb8W66F/+5gb1uo20BX6cQF2/j4+kXVWObcQT0y+W832evoP0D6Uiw+2+HvqF6
y7aEFo00xDp62xFqZ4uGDryoQe0SqupVt4lRuV3lvniguiRlJhNnHboZRZKdL5km
054pdCB532CZwElVvDTiDtximu6HXPwQVTU0Q+QGwnWeMJPX9PnQ6mEnWRSKrfnx
fvdn5XN+CKrpbjU8d43KzDjibolyvRqy/o4vr8nfBDYH+GPgdiZPOXgIxhehgOl7
vVrIacEFyhEYAO64y5zF5F8QOGFLuYmf3pJNJUVd+ToUPAOYHx1Xiixl4okzxRTG
EVC857/jHrGLJOrczC19QFVHPKvb8w6Q0cEXq3XRJT0mU9AloEIVawQ+EytQthzc
dyZ2Thzx9nmrz5poXzTHR4oIXbc1JWbTFPIPIQHNEMkGhlh4JK9xwzqgHVurRyrD
LEG/fS6wRQmNq6JZWQT7CZkqnq6kjsM1fk6KXGJvo/VbrdjfQIEZOhgG4+PWG8k7
WE4KNfZuOh7WtlM2v7a3i8RAfFalNtM4AphyAf4xJAVUqdMMzvsT72ZSdchGUpEI
Zhm/WejRaSbU1OJ3UiO/N07tO+jm3OJ9JXHkcBMRi83FZmxDbIIGnZcgWr8jXbKm
ZtNUzludOQyBTFNW9IgsCwbuBAaY4HTcP4auOTMCurEVPyOSdhBJ6Kl3LX/DXBFI
p7o9H8TXRWlgR7GPeFAoYqADBXGeaa0LfphbBPVE6qEWKgPjZYNduOQGCaI/acjv
Z6yIrxZG+igCA1lxyJhWGTA3WASZRluhRqpPeTb41s+JDxdANTZ8OYzD5kETf8yE
lehqhmVL4yl2dLrEHTwANe5Y2aXniFE2AjDMS+D5p3Kyq0WV8wkVH3VIrOg9dxO8
fYIF9v6yH8xyrRcAbGUD7XJL9tTlhaXSI4y4USpWzsDRtSBS5WRhD5gxAlYvaV84
eUElcXoS8xFnMqXPOccZCPNj5ui5npzdANOv7v2rc0peFytKONQab99M5PCYbZGO
l+S1K3ICBoB2Ow5yzz0QyR6J6TeMbjEu2OVV5+a55gFyVGTMTfwzxK4jCRseOQZC
RG8HGmCK2rg+U1PwDhCgogKJeqXm/oh3BAhRilPl9b6S+HjOmqo0XN2VQt1CJ5mN
GtmUCX2PRYkseTnaCA2XWjrq9yOl1Q4HVZoE7Oe5GmVQVK7oslAB3eA5U51dn9Jp
A1+CEvOTwjkfU1f4SPOrcPCSZGy10IITRyka3Yt7qt0egiR01ya+InKQObGKIyg5
bd6ysspU0bh4FC0jjCFsrqO6NIMb2FuFmSS/+tlHaAp7++/ZMsAQ2H4Des5I+RCR
IcQl7QtO5jEd0lv+dfpv9mt2fRJHeRmiVJyf8b9FB0zZpx7GE2rcam+Dm28oq3zY
g8n+m7g9bd9GUB9jVIBS3gGLQ1/oLcgFYQGj6IiuCCrEmD2NSWzj31ZR4cBcGOfM
hcU4wOL6v6ChQthngOkNpzZMH2BBwXRwwmKoczRH5EZMnwy4Ol7jW/h40h1Qua+S
tPkdaq3Jlg1vE4TCi13AyQ5LVaC4OxwpaOPahwE0spFXI93kD4d6aMYEvujTPDsI
cO/ZQcseiFOJ8PVNE1//CH10bPT7M+1LpBvDpvp98lEIfk+Vxn0Cw/OUI7Syd8iV
NOWHvcOicrMfuNGoEm+uftMmi1oWoj94NvyW3HiBagIjxJaufvWcy5rGnFDfnyf2
++E2Df2/krOtmKMNlBVCQmFn0vg0FKrxVIVH42IVvuPrL1tIGEqAyjQL9frxrVd0
C4CRyorNNaesncg+OP6XhyPdZp3OdejZUt/6RtEX3SnlwO3NxmGbSoU/pLXM91Ac
AR+I4JVUMoXinxEY5dLYPRCjilL+xaJaKF/jjFh6gCsc4S8rlvClne6lRYHU7sc7
8vmeLFyNhaW7hrDCmz/6Hdd+lYZAGcPFg+oa6dGwyS0A2Ws55bJagIfrtDL70mYn
2uuEnI0e5yckv3b0UMfFhJUyz/rz4ztiCTvMLbd4EprIWeQLkdUWuEokzexW/2XM
Z3q0iiRwrb5eDtTTTDer87Vxjw8eSrlpmd4qBNaVTt+8XjjMm7gTP/r2rRKRTkPs
7qHQoUOKajOsnpi3TcTooGPV2JBlEWmTnyz51gfIp+Iou4TDCSimjqQcD44FSM+F
GW8OuEKSUABEV02HFLF3vktmccrvaF5cxVer7c6G8RcAOSK41hstoVtS6oLar34o
FdjoKUv2XS2gUws25vOcWuq1bEXm9ZiKMJSRJJlPUr8VGsdrjMwD5IBDSzJyXttI
BLujWyyrC1fEc+SaQPrec3Q4b7uqzqKVO6X7xUQBv2ZlNkqrN2r87b0sfhFzDNZ2
qmdWokoljZBB2m/QWv0RedK9EFKFSgyVOOPmwqRqW0l3juKHiG0txQMdpmvvS7iJ
LNv5BP+Ua8FuGRw5KXVZKwPgTyY1/VLs3SUpA4L+TumaO4AvP5SDJib4TUdixcN0
CMKS+JEwFtF5+CzCt6vN9b71KmCTu6WAYx3Dn6yxFg7O6KmiystINBMB6qqmgMcR
vRnSVF5RSzi98sOPsiE8KZCcWtjSg8qPV+UKAmod9WyCI5JFv+Yt/281Zq25vCZC
4FfYVcBbtJtNIIBdmbbvemzghp1PSx6iDnGxwCfrk5+EmQeFeLZ7+LhlG6pt/HtW
dG1n0aetWhdc5sn5LYsWweKAqKpNzK95MFc4A/VEUueDeiNuAbsHDnN6RMuRK8A8
E0pVwgsN1Ps2wCOzjXU/x24LsPBYr2p1v47d8pc4KbZA4kMB74VG04VftV9Gewpt
ppHY4UX6zGSuCcLiu03SKsJ5vwrHMfCeJoMajZh1Kcweii08UN+hGOKNqIjEfdKM
1vv2sX5FYIiAqXL/8cIVy+AN9Eva1cWAzffct5pGHot7BXZBd0oFOzUxwqDn78Qq
5kKv8x5c1RrxKDYEAyVDOvjf83dBypcnp6S0n6UvQgOSC9QMHs1Xco2rInKX0cWl
0qUVCZfiaUzpC5gnC0r8BnU9GhyApH9hJX27p2pO1Qy/ZoEi3XHlHdxKeN+eKDKM
QM/U1Whe9GYJPySbR5MkQj3S7bb/vXVUV4BG2Iv9DPVPRmwx21+fN2/ZjVGRvYpn
pti8Wh6vFA9a+mn8OHkTNFdP63Eo90YAxfIeXK1s02ghwIY75nBKz30bvBxp31pX
1JU4qzz/rmsqmbESAkCdW6BKr9ehzovYMfNn88eFYv9ogfksTgs/jCgzIGf4x0fO
3Dx02mCGywBJavUn+Sg7LB2kTYNz5a5nUIKkrbQcg5oIpoGpQCySr3o3PO+S3m93
lDQZTy4BrDuPValcaGj+yvF6vE7C2e/6fz72fTrMNQ4BA2CWrDBoTW7O11LrkeTW
OhheKFfVGMiijT/71X5R0m4Ty3K/CEdsHQCQUhzagBHXUp2sBhARyWrwtEF180nA
IKVgo54kggGZm05jpHT6bpM0mXCzsPFcHijaGE+Td27FMSAS1NbnslyAcOXAuueT
IaeeqTIZBvBRp1nF1jDAVXGKmIHKr2plpK4k8llSsLoUy+vbWj1cja+jf90Q6+jR
HJo6KL1U6n0ES81kMaKfJlc1Z4534RV2EVtlF2gKrTAvkpduIKipA/YZazFqVakt
Vw8qvqcEIG1lVVaMLZ1auAJX++urvs3CVlvlXXSmb7ZLOGiRYBzdWyHzhqzpj8CD
ZZM/uctTqML9qWs9ve2V/rbSPrjhgfw7g98gJjkb3fCuZvKEvr4W1PqW7aAcRe+F
muS8EvDvlkhJfs+witBLBuA/xjwuG3mhKRw/fKwQ1Kw3lrGFGLCRQb56JfGkzmui
jY35X2/eVV7XWnpDymFfC9e9QGJP8kdhXWGLLXXosZhA5W+JZbj7kP1jSONXfUBF
0wXf7Y2U94oTrWCginAaJZ9sw7eG1g/OkkUpe1J+d1ZOo0bbSdKE9mulvImHWsq3
S2jPvA81v6PbdbMYqeyuq9NYYs0YuHEx35PfYjJl+jnKLavgoeqdXrFS2vY6vTUW
9uR+UFtmIHXEeT6b9PDrc73I+QJnLvQjvFXHrYw05aCAukd4TmYwOVJpU06XscSK
1EC+Gqo1Cp7Y3gngpECi6BzBmWxooAz5+5pHBn4eZrH34ZqguOJTk9+4MkLvP1lq
1dKvkZHaQSim0cb9JRrpyHl5lRjyeAor2V9R47V0PgCdMO1nZz5IiRm9FcKMAz1V
jIFOOAcX5++56zrjMX236JggqH4Cfz6/y0iX8gIGqwuGTsr+HEthhy6PmR+YuFqJ
oJgDkG44S7EnlNKoGM0LroFH/ueNoNTbXJ1rQZ3FPxAfBLidWBk6kTIV+KgjlRci
ownB+2gxX2d4sKvFMDpNx+/lnEutWrpzc5nnVwXwdKh84qcux9mA6rIcaIEzyOPT
Z9ebNMlbZkmfDEUzmgK5QmlOkfLHzOwjIqLTtmKvUKi3uSmDjan7R3GyCW5o+VEe
4ICPOXfJrDkOlBCb9UwjU4zENfIEUp4UvLiUO0TM2ljApsay9WkLapFMSsReORQ+
30olnLUJAzaw/rSQ9JXE9XWrScaiACzexwG7rexowiAmdqYWTSCa88Y4vjfXgjum
/pj4cmtY7rNd1Q7r3fbnaLy0O3ETN7u6NDYBPrQaWfk3szoU0XoHFys0FHSqkjjq
H1Qcv6TaRPPYpGGk/e1O/vk3jNDym4RV+soTlv9kiwTZx3T9jcKQjaxr0Lma6kF9
Wfqr/Ubzz4uiB+c/IiY6/komcuueC6bWY9cJIQLK8sCuJRzPJR/GWk5L6FZdbE3v
cLqxSAHWlm15/T+fxdNReQJoD3LGjf+v5D1RYtR9TxsJeICcc3O91krrPBhUtxiK
k4MB8I841xnhYNUzR03b+Q+ziyp0wPL/iGsyfOSfDTuDyI7dcimmzH+qFZpDBqmt
Jk3VGl1cC1qhw7PW9RVLWMr2MMQYZ8EQvlrne1n6J//99v76XLUX4qsXH0FIQpsu
gkTdhwvPbbis+t98bP0bhhrHirIrBhaxVxWWthVpWQMt0Cob7VvOZgC8GSih+nZl
2qzQXnI48IfQvJcB9uaA10pVIvcah0kHvFNJ72dd0Qqv/4WAyd/lXJrZjroGukD1
7wv0UC5Gv7lhvzbrSmNXr24vkflJxVQC1+noT0t43W8=
`protect END_PROTECTED
