`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
stn8iGwXkOo4WGW1lGjg+XBYLNqPGI6C2EQyKKo7Alaoi82ESDKYFxvwMmA+GDmf
V9u7dD7emzesY+vEGjx85Mp0l6IXwfpxJ18T9zUGp/N29ULdOQCVWNJXBbdIVj3R
/IDShfrL9wCYVgkYm+3jI9BAVUTvwqaVBJ14nUS5a76k5I0+DbdQc0hM6GaUsf1d
2n71hz5DYA9mxvXgRNadTx2E/hxRBjH1CC1kBljWZXE0GBmGCxQEPo++cEHQ0fVi
gJ5MGvmz9qIDCx6U6myy6Q0t2xqUAYGHjItzMTdk0caBwMk24W5Gfw4JpZwuDKqV
DVuyFZVq6sf9EF6MTc1F1Ib6J4FlxMfCe5TRtthLwhp2VFp+4ZOhS5wrI1Oym4Er
FriDMP3Nmb2Hr4I29luVFOTh/ZWbnbvP47SSkD1eTWRzSOxzg+LYu5QGBiogdPtF
g4Umyx/CU6JC3AsVxWgxnN9d/JK1KcGUNFn4tfomSfVMDC5BRVXDSyWwjEjLDovt
Z4H10WYznwSLxhLBQg1bftqW+UbmIS8WoIxN4WI3Mr20/IcXR/NiN5zMd6SBBzgX
qrbzvd4VDkW53xpKL7WICA==
`protect END_PROTECTED
