`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZPZzaVAaFJyJCLB+z1Y9R2nz9uPgf+iYmblV4+F3TroAvJ0w2UN93x4Yms0eWCQ+
cYPdrdSyveL8/aQby1Q2/vin/o06LgZMmVsE9CaVMLIwo1ZqbVBAEWF8+8NJq/c+
JBKbj4QoIQbLbG9i0lskmvB/fO3QWNHgP6j7huoLX0jDnAFz6w+uJibnYQQcolN4
4bwKGoyl3lB1qCLqTSO3vifd7aefkDpa6g6D9tvJ8y9CcUTyEPK5M6T/1HgIsKdG
UukPsKArmSed6up79bzCINIWkn1Iy84h5/eGo2OocsLDriV3EVutYVGtOmqSGDTY
jpLqQj+b8YoqnPU+O0BEuZd+muewkfOCZsRIbNQAvHlQQphdlDpxTQ8h8OlF1O+E
dnZG9gBn4iYpqsoBMDBkMrO8RH15GinVPhpkfLOiJ4rjs0NqKnYs9xOXlZyJHYhE
objWtZm2G5xke9HwB6Zwe2nJxHIOlfbx3zeNtwhukXbFdWfkpvi3mhuHJiWaKwVm
1fTA4yzd5dE76wmQprH+0rW4U825FdKUI7UDCV8BgjyeL4DpDV1yWadU61xsJJDH
z76dGFxBk/OvmGIHr5yq/du9IezRLWt5/+sW4AKLjUrL2PQJYMSPH4pyA7ynOQhD
2o2TwCvWREmK1avgoSnPoLSr6rOiGRP6H0zEgIYxHjVubUUcyY6jyPuJ2Jv5ZVsB
w6i6Xr98uxlgofwtHJs8pw==
`protect END_PROTECTED
