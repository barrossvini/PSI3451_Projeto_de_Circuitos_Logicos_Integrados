`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nWwaX6AtwQZX9TTkmw89xtcVZGdPAikc3EaQFsN7h5eQbIYY2EHoG6A1te1tfeYU
QQFff9v8cE78KbhrWUfP4peYt5J5R+UmO0jPmgD+ouK9vGDWDNrnY0kmPdHs71H4
oNRjE2GAa4yZ+DFsFjHdStR0wP2Z94fq5ib7nz7m5TtXGwYU8XLuAf0neGFkjQxF
PidJedJ9f9MWhgtTJUBeYBx5i1T8IA6K47oB4zzc2fv0nBYDBqt9HGvB2+gIgIeP
w7AyP6oRSghDjjuCTpo93GLMYKfhwqwqLSHGW2ENjVhjlzcGj0pm8w68WZXvRkvw
F6R4T7pl1iIUJx1EEnpohZqLmCRmsIX0+JWTRcm2K0v0Pa2g8Kit5rvUF8qUKj8k
6MK7/SZ7NPaKkLNDRlV8v2qyhhWlhXbx6VuwrkAQHeC8BEjMZYjMuFs8ITAFnmoi
NICyA5un/NN133QLGrFA1w2a3CrfNeNUEIzR8AqHATcwjXBkk4Q9uzYqR5fu1iGa
czc8swKe6Jo7L5NXqk6YLfEfQsUhfTpLXX86LBCBUyuUEq+bgCbm+tmPO6JWF9nK
HQeaUj1lucX1+Y+6M8NsrkjSBZL7jv+aTvEJNgYVNIpwkOulNdY7YqeotAPz+sHx
kDx6fFwrox/ZO2rJYiIQcpiruZo4aRz5jAfP5ikWwD4bDrsnqUYln0eJxEZIx4CX
H6UtcFA+Wjcaz69npK9pXzt7W/OFBO/51l2JFkOK7CuJt9tMlqLMtBvPQ/J387fl
sisdGEFanFFFsPs7uCv7aEOqcYMtG6EOmL7FQio94gZe2p+Xdn+NoIpPuR2qrBBR
jzk6wp6xtjrzQ1RgbUuOlbTtCQHME7UTGJTG2Y3h9QIY3RGqkEVNn2fgNgIq/CFI
3dJMpuiCIGnNjbsxl5Qrg0k//xUZqzx2LLAge4s7WS8yaebeuN3Z/RnVlIb7CJ/8
5WEBGGCRPGPqKSSltDuefMAOc/LvB/fW6NDN3wE2YWoE8V9UB0VpD4LRwISYv9Pq
NA1A3BCdsvf99R3zDbVPhvnDrg5V0gsHvxOG42I/mWsW6p9tqceaduEoJGhMKycz
eGPOny4D/CzlX4Ugrf/LF0h7dmBlr17qELL7+3/gfu4HModV9EWspG5y5shSHfHO
2McEa7zAobc6trUtPaN/2Ehq5AzdZlu7lvKCI7ueFi01JAJyuG6MFNfcoBSM0qPa
R5MdHN4ZhajS9SIWi6upGIBEeL3nXUw7jtkW8sIklhNWVjyfliJKJPwWEFjtYD9/
0EhzkRb8kTILC990Kc4iAFXXGnBGozNUs8brW6ykQWSijx4ajLT25+gt2S3qDKOP
I2p6OovQFXD2olUuieXl6G6/tLiq2u30aZ5dmQv0QA9Xhb2VTVCh5gzxXW4ZjTZf
TBfBsHMbfO2Um5d1Z1sKqKgiAUHELsFOhcy4KnC7nDQY2YnzewVUgu/QPlxAioLH
FmnHcpmNHR8GSefKHugvxxyRU+B8l3scVAgz8c/mhs0XAjyPI/G3rpIYMW1vyRry
LWn9XL+FHURcrLETGJdLHw==
`protect END_PROTECTED
