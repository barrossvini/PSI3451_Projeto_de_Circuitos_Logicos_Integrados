`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9l+k/DaNOnd4f1WAvSYpa+Ap1Zl4SSd6FUtwZR3k5KWHSCaYZAuCk7ff7WkDf4H4
Nc1Ri0ijhWdWOHRCAN0nN8aNl18Jw9w2XDTjMPh/Lppk0VU5f3qoF7ZXNiFeE2FS
S8N9Wew9STPDKjH/MIPBE6dbIIEFOKa71dK+678NUWUY6I7RQ47gs5jbTo7XeNjZ
7WFaWQ8rAs1+RLHb76wP9Ph/Ic4yguLCztpSUpgN6W2TMGm5FKE9mc5S2iyp6QMM
ojbaimvccjInAyyh3/Hxm9BQ4JVkcQ1aX48GpCujFMyiSCVfUMjm9z4PDcgejgnr
5gsnRHMi2M7kqqIRCKFKPUavQwmhFegJvdZm2yML+AiqfdblY+7YDtfSqMBXRdUb
OaLZdgiYh97zuKOMy+wv/INEYGM5qmwXC6sryreQWRTFqk3fIk4J990uPXDlOgUt
EnZ/sw3teZqijGwSi0M6HbOSHXZbdG0Pg3ugeGAy8SpCqowDNJ9xN5aq+LFBbmaz
EhT7dovE5nLDPL1c/uxMp4m03jbx2aj9jq0WoWzUmWT4yjeiSwSFX/L0+PkrdkyD
Wu5Mihl6QofGZkOl3imyp2kBeaYfUb4NfOKYuT5iJn2JoN4hlVbQGjIuOzwNOIzb
FU7nnzf4ZERhaY5ndfkYxaZcyB/HhFnN+SQAkvytsDIBz7dUeCK4prtGkht88eJs
5wFY0LGHnjpYbO6B3AKneuow8u0BEGk7rP8p19Mt6LHPba8UpVVvPu1+T9lP+Tdk
5OwoQTsPdSX/oFt/5ynBOBboziQ5DjlJylrRk+ZpxbOcF6JBb42O74JoDFcK4d3W
iIrbzqq4Pj8OMvqe/U8MDyTbWRJqVw2q0vsBSNINfUBgB3J7/TUJ/ODv/EYHBaVX
oSNQ5++RgVVNPq4J7vAge7R15cWSQxUm7OpZoT2XYi7LSB/CITWwLfV/2VirYHcg
C5fP6mVtzMKUtue202V3lPc5ZX5T/RbhpieUg8gHz39IPKSclAUi/7qoJDRyuIu2
dSM5pNq5hop1g03VgPLz/+Ux2JY3eulEpKTv6XrLRkhwqga/Sj232cDw0lCr1Cn+
dveTdgt89zxBNcVuxxC7iwgH4wgoGhA1r/EfBZa8psGRbE32uRUrC874oxmBJJZ0
ISZIQXjVLEraGb2QimPC8fTHT9aRewh9ShuCxkknggi1bNNVkEfDuJP/udgh+FGu
8zu4Tmd1V3G6HHqi+hS9R9cQOIOqdKxX/0EdPQVFZ3WIWNesynWa3hcNJrvXiARp
SoUPkMi1bvIo/t0nhYEUtva2E+x877RQpX9JXbY/fwkwYgF80wm9dhdyX2rMdXQh
ublKpkFQ7XTaFK12kaBAzhDgA8xHV/I07uPn56kYNA78hoHVN//hjSrvlnt5Krae
Il+XathzA80v8WCJTogY2PwZUq/bJpIDZS3CJW/0liqA/cgImXP6Cm0thUCEvf1S
OaOTL59fY14bZpRx9nmL2M3sp2DLZasXgwG/eU/qQSMXWvRNPOSb9VtsHG7pRJlD
SsxOlscw5dBoIfv/IWLEKGgLP0AxVZ0ILbjP3uV3irFh29ystEti5vOzYGrtlEJJ
WL1u/h6MXoLO0XgTtXAduHIGgzoVqIRRt+KHTJtP3ZxXG+U0CfVEzfgajaqke7wz
oIqpQAIMMh5ci5Cc2IZYoWNRsoIySO9Axwip7cHXr1O5Pd5YSjDKYdqWURblPPCf
cp14mGxlbErC6B7XAoTViN2gMBbpbHm1he0kSluDa2icPUbAwJYnL7GkHLwkqEhf
nvqdjUrvi+pxM7DoWNafyi6iwMen1pqKZe5kwbIFUcMxu9LEUyHkXbVHJx84ZmPJ
UojyKgSfqunjUKAFE8MUk6/Cz7q4U6mOe/TuM3/u1zV9vw0yZ3W/72arOEfRuYEI
C256QiKmtqLd9GPWHACRUrhAgAdM0z9+JEFJcRymE1jIP0B0kbr3h24lxT022TFR
OLPDeyhCiJldHSqu2k0ea55Nm1b83SqKrf3bTXKYg/zlMmR40CKoQecKdaqe/UlI
Q30C6/rK+JZEA9EhqH4q77ZLUzX4lu3+cbRKOAVlscYx3P/ObdTh7U+H1qzCOOlr
+OHWa+kbxYY4NwpVN4GdHgTxFkm9eRkSwDWe2SDUlRdNbrPXqboMRoxLs/HZ4uOx
zVMI8gj7aHWV5dvfMcEU2yODnEVCpnNh4WmDry/L7XSiRtVDqux0L+akPWJBLopA
EXUmShCWWoBG/SCLwWoxjuZkZAqTNyWPI7dQ41zCoCPpL3J1HWUZePhKHIByNbf7
04bVaKCCw4kH4LX27YLUxFwSEwnGXiTbiY/MyKd4jbxCfuok9rN4KeSKZM1CAN7d
PrCq443oBlMtEeUR+43exfpQQqRDhL4QW8IanQJ1pbonWLmmF7pvjYjSNC0aKkeL
QcOPia4KWTWd5T41Bq4wLRNgF/+5VCvX1qrmVyMzhFqJtea90blaiIMCFhwNdARo
+3CkUzfvV4COa6NOck7ZpRh+9WrPJmDCE1OgPylEvAT2SQQjQBinrWbfCf6rBudx
fU30cOEARANGijm3cuEaSeeOmDA9+MwJYiYPC0128uFZyNWJC3RenMd430aYq2aP
/4IJW69FFv70LdNkbcM04lQ3Oe6IE7hNCL64/0LlYld2tdJZSM+Dyld5kPLHWjps
eR348yz5wZjb2MJ/urZHNCvAOsSn9dz1XqT0YbBB5E3Pyvvxk5aF9cZ3g3jMJ8mX
4bQCb070qF0TQ7DdbZfO9ubSS/VU0vMvrpgaTyfxIn274m8B2dTLbCORFqxHgmXP
kiV4w5fCxweTbF8eouV5jIW/4HWD1XpLov/aCMwlOPx13Iwrx53T8+YvxsAqYNnY
8GfcegDi58jN1HwJDXB0EilAa7lIoG7NDwVdeP03BhmRNZMDhsUIbuoxOdLEIwnp
2Uiiv2cAJNBW/eGbwC9ZpAgscFDkH+zHZ9KU4Jo9XQc3bIkeNXgdvGerzRcXGmBt
xIQ3HmlKszn0YmZ7H8uzbjk8CrQ41RK2ytV5tPD/CImOHFEOPpchSKgykWB2pJ6r
dVDiZmdjcYB2c0DuTWZ3Za0P0rjaj6vmtknmDV5nvFbdFg+cyUvLdlRchRM5iQPD
ndkHDrDWnxXH09egF+RqDLoxEgtZSj94E5hkDlZf6rLUIFm5h3MLRJvo+rSwhC+t
KbBjobwW0op6b5mCxfT31W7KGFBNw0P1Onr1iJq9Rt/RLfQLZ39OAUFY3MzD2f/T
d7twBwBNY+baQBr5VkmCwJ6rY3pT1MeYCCelviQHQQ07xX29zO3ot5OxQMk7VKW/
ZFf9dkeY0WE3m+mEm67eFpHp8+/bfuh2a+ocNoTQeFOiScrydUBh7yDrTZAjHkam
1AZxvG4KAMb7e66yrdSOD9LfV4TeoxkA35qyjDvZxMG+9SrH9VUxN6fJnR8jgiYd
H3fCo2F8I7ZI5rOZbJ2727cYaTDg8k65rET0uLl+cF0ToGVlAWBoE2G4zNyawMdW
AwO4pI0Mx4sjAX/XfnbEcN0oaOs2+c+FI2RlVB8qEWNV+G4uP1rXbIe5P+hL65zh
GHduoeVdlOcIT/D0r/eLlgr+r2+QkUfDPWN9XYsKSQHFm03PEuUbJCa7VOGywGlk
HRG8ZBXKnpg2k4d5vsv9DxkZTmy2U1wC1H/4aOIOHGBksVM8EpeikBatD91bIZ0D
KyDyAEiB6BVdOXD9mzhvl6EZLR1R4BdsEpXXWlP00AL6Cz1R5rT1RhGGLoGeV5V4
EsjPS1dWOhB83q4wl1iPQef6MQX3d0E/0boDEsLN07FuXFjQWVvCgx20anEkt3xN
QeLSaS2S4AUpbhjgN98Kw8WEbCVZQSbeAvaRgNMmJ+XZrLyjBbt/yyknO5h96aUq
FAxD6/Hl84IalyUFxiICrplCT0rm26pxRUQTaACG6V3c2gz5iAYK0aBqLwjDvq1l
E6805UIozcdW6K2Q0HWLmc9cxoqLsJmezaayvai/gBf77dzlDrDwjGv3qqR9IcV4
Vy49+I/IdJExu/SzH4dbp3zgrpNnmwLqDoS4NDz2G1IKMzVs165ohTQRO4zysJzK
LlGs3MdZJiXBQS65GYea/6/1giMkRDAjRWv2+GKZOG+kFJr7pVLx9gt7/jLqDggj
4iuVUROAJjUDe+3CG/YAGZ5YG3nhd/ko0z5Bln6lbCiiJCVXHeqdJl3r85RQGRJ8
j8UFMFg1uwAx2vtzPw/vH6LesYkjAMKDJGIdbSQ70X/60A0M8u3rCS+IH86Z3fpv
r9agDPcsRIRYWFf7HtWRPUjBJXsYqkQRr0GvDbI8e1hZcYqCvk8yu4YBuX0aGINT
m5U13c9NVflvUH4ZDKlLLH5+2HTArLQYCy4lEJONl9I6forZRYAAkWK0ySUKqUmG
7a4IjhNnhnIvVVjvnwNehy0NNgKsp1XpOlpJSgqmMoXodlZkI1p1SriP8Eh0ATCq
GvFPyKfWs6bdZ/f1L2c4lMG54O31edb5O4xHh2v1Z/VfmjBhZ+7vqbt9jJaplbLp
IJIjj0nhw0ci7TmQ6QLrjbuvsDO4VcJ0ovQ/TdVp1xOVthiIIPH+eYxRZ8F9W1/a
pUbkOQjNlKrdQ1qkBHuZcV80ACBMRg9PKZ0u0yeavzX6FtRsNx42j7FVxlL4FGdf
8rl4wqFU7+g3NJY5cHiFJI1foEt0wN5SgGwup2eMA4XjAD9V0U1xxD/sEALe1aiy
kRExmkxLPtJ0YwxvZtBgfFZHBGyNORNeI48Hg2n8AKljnz4NFGutUS/F0j6rlmyI
SCx558XncpoWkVhvXQVC7N0kQ3xk5wHt2WHD71ldZYk8xNsltNbBK80MbANBmlM2
4PoGMJRJWiT7GpFhvs8d4EYSBKj5CLyRHr376WO/jB12NfKPR7+y0p3Vmkh0pd54
KNjhos1P5nFjtjTn4vdPjq1HbW3DFJuUgnzi0PqhiDiKpPj8EPOoSrqBEYKzmtLU
tjq96F0J44KpFmmXYVLvnS8UfPrzhsdkVKp50fa9G+WOGOHCmQShWu2sM5R3f+dZ
dKq1Fig8YIqbtBbjCYYC0lAL6OvX6AP095tYfwzw30K8OqblxGWDmNsYXHHkr6of
ihjFDUayKwSxBrjaimFfTTTLRendWUOu9jwAmTVLHAwxl1hWpgiog8flAhHf8DDH
YHtBNCKCuFTk7EHMznuG0O4E8T9V7nHDtPOj14Sqq0d4/PUQTzoSkPFGh9MkcysG
ZHtH5cueAjKbK1nOQqfLlUh7EtlXVXGcPBFy34kFUQdhWWPyIr/b36Zf73EvSeoV
OoiiPzEempUTLcfHR5Cv6kfKiXuc06iehnhnm+1DUwJYR/EV967i0B0Ac6oivpL5
LIk92/YQezFcjMENm25EE9MbXAL3ou7p4uL+/3oZKFYgmp3TwPusySxNXzAsqrwl
uyJ/8sVe0Nrpb4lW12Ij+WeyRSKCMXmcI3i4x6hXSPw05/9N6WCPBvmpnGlQe77z
K5LWZWaBgEkBbul6nHKzIHNDJ6rFdhjSnfPN/WinrJuZt0DPNQtryV0pjbO5E46U
Fi6Ou1PjDwXItij9FH3LRo5y7ho4ZKF9HMZ97mYEXBkhGU/sL5CSGcn5ALhHNKcJ
+RVoNII2BPk7vJaWvosXCchriLlVYtuy20FdS066cNZg+UOB0MmstwPmuCm16/ww
LEbqhvQIaglLZIDqOvQ18GRMuU8Z0BNN1tZG5DP2l/OeTXV0uPKUVKrdOUIK3xyF
SRqL8l6wtwWAKYzcRhnbEncQ/cVmKFKGatUL7C28lPUYNXnEzwskvxW2IGwKmq4X
RMfdO6xh81Fxtxb8SRhABQqupXnXmO7+I0MoVw/7KheOwQzk3VJ0r9uqEWQUKoB0
ahSJklW7MI2L9B+/8Xh3jipfbb4wysr1tnj3swIEAEsSUs7VowUAey6TW5RRNz24
e/u0Eg0+oa8lQ6yYDM2LOWDPbXaQQc9KwKLZqrITaR5gGlCJLvXkIq7k6C1pJ6Nt
s0GgjQ+OSvkUbNN/Ep2deXiNkqBwpt6PDaJ/lJ5iwWLuOm8S7Xxl8EeCEFGylbNo
WvOsCIKIcdzpTBv+62s+X62KE1Iv+ZTkigM5P4RqisXjAGF3pVEovxnNFpvpJM0c
bIX9OF8dWJ8yZq0UFz+ILVkxBAAuWHRPYUbc3YrzRyutocwqRNe1ZvWbW+AGOK8z
vcSwDV2E86ZGtMD4ZYBFN7QiwmahxouHNvUJXN354F5QiKTcjT090Wrc3A9/YMZI
Zf6kevoq9Q6K58yLpf/FQhd9hhgrRd9o/OOTFB97tzXckRsfy48eaIzfgmdQMGFZ
xWO2iJyX3LWLCHHTB5glww+QhjWe34e4k4xf/NQJt27zF6wiNcvJywt4YHarZIRy
q3I2RqB4ILIyf9uUZo30xN0zJlFKI7CdGFxMSWlHVL4Vj5vKQxB6EoJ1D/J6xCTP
9hR7fbTo9qvp96wJ1rf8/4VVJXe8gQOi99SZFxJybCvaS/G9diK8laja8M+je7NB
Z8Q71H8GN1+ED/EKb+PPRHRjPgFelkivcow1yL5bDW0SGQVspAJneuUwTnY4dN/s
utYAWhaeB+QYH1G1AasQvq/Yifl1jPyRKsU18d77BU5z4HJ6JIbkGszWDIkYxcA7
9zPvqnxiZBprHu50jKBMyZyt+RJATByoXJywJoJIO8q0bjHV8NZDzbTEtCSnHJTI
fl+dbg+QhPPsoVtvBmyXPlnIWBB9TsY6Z7jxkaZEB4tiGsnyxopZYFbtldvRcyJe
YJap+s5pRHT/E3oPI1+0h0D/QSCtuQl7WabfCXOFxF5QicNBgZ2NAvvovB+DOvga
XYy4yxnco7LeqqM5TSEONKikwIQt3tOwoDBcBLNklpGTnBED5+8b0Dyp7oRf0ruf
JsAEH5UMDRYOB4DCR/uxD+zK3xQI2vhUMJqYezQ930OXr5JjAYHdii5ISXCCTl49
f9lGPF5USOnn3Dl9ATSnn4Ux+Cr5xPtsHbr1wBchhL/xVc+a+fA9VFkDnDK7bYN6
Vlc7huOANyC/md+fOr4LkUwgDlrQK2Wz93tfWNIOgErjwBRdR0M7lm1s2eNCHNjb
XDutaf+FgH2VqUoYZ4El2z1cd5F8nlOl6FlU1Bulr0niahpgqOQSRyby5ntaMqCJ
InAuXyxiqVNCefu+dciUnhp0/VIhs6B/uB0BfAEe5KbgLPKRMGAykkyQ6roKt3qV
MXrsUCJxro0Vqe2IvtH1BsZwqmbhmpCUJXpxcEffCOh8RxiwefDDeylPgs7w8ITS
jqyKjhfwQJPm5UqD2ot/JjL0sjjt/BUYdUa4O6enxGY5dJ5L/Ns5jVOkGnfuEooK
LZNR3oXEN8+eZ6Vk3MDTTg/5BhE/+ljubqP14ZWtJkt8z8OricH1DC159Ouy8xik
eZwAD086NUdgiGN0OcdtR5IXR/TD6PfERFp99OolU1Cxq4+SnXwCTWbIrobaDLZY
JHCi9wjhfayq44o615g5+UJCHo0huT9knDfSIon1tUMTX9eTtaVYBTNX/23E3dYM
HhDBla7O9jETr56i9ccbHq9NAMADtpXFW+D5za8Je2MI2sUxNDdJ9b7yPa1AzECP
Iq+hIF397y95v1De8Ppx0bFs9Ka2V6+gJYTVreL20Dp00FJHHuSuQfy+hWfyLLc5
bbpMCZAdbG1ueep1tdeKnc8pvp7nIgoneJk4ALcjy8bVzj6wKEH8+TDy747T2ZCl
OpdKK5abVorm4dKii6SdERuBMcQuNtnOc6/+csTkfO9W8mifrOoalIPfIB2ZfV41
tcQ+HapfWt6/LPsboB3y/hAbUJ2pvXv7zD1N5cV7/clt1Bxn9OP474ki6mO3y3dv
8BEcAPSkY7t68HJF3jbcz/mvgDFs3QzpoyzNCl2hi5p5QRM/V7FYI/3LvxgPU6LV
HNun1MkBgidMAr/aeqQpPbdRbTbXO9tzYkmlUsh6RaQ6L6hcFUdMtN7kkazhiAH7
Ljg16qg30Dq79+rueXLYQQKprg5z6H3QB8vwqiota0kf/pzeY3qIxjW61BRmDi2j
Y3i5QwjYNP6sRBAj9HXRqMd3kGyXKYrQJ6pfjYjT2DguO9jsP73JfwI54mfjpalt
HzxgO1WVkZDKePbZGQOBwayJB1oKLrdinePmaFmtm2jtITk19lu6G/q0dtxwAMBR
y/b9bHtQ0VpcowHs4q70WR0CZC1RDPnDHqvF4z/tSKMtpKWDLJgV6rrcbEquHc5k
WCtckesJYw9hGCl4B2bQzufhmMn4hgans5GZSWRt+52SRfJHbKdmUn5w4A30N6bs
KCUr/cixDwvLUDJQKfqYNZKJKwL7TYN6Escpnwm567Ro2JNvahkk3HStP3I45Ua9
WTTt6mm6YkHzl5lJ+WAPv6m1ohrepuR1Ti64Y7hHs2wvzuSlIJmpXQiTICgFecUu
6GSiAenHxYNozGtXdxYcjZ9grLSss40/JO3RBfAic7/64Fy+W4qddoA6NFGQA0rY
5CSIGhZdUYyFdGbha0DwAwZ6VEnbAte5HNHLZ5OwXQYzL4pFGUiL8TeXJRYAxJQR
MeON8+7okMZ+9kX71pegoG7wRohX4IuEEyMa2NRG776Jc84xT6zh6HhVhukzEOjS
5cvZapK19JuFDu5B12V/b6vrRmQ5Pd8EPDdjJBPA1B1g8wXhJ0X+lMATzOP18qlS
UNiIijQyD+lNkSJ2hnR/PrPAlCaz4Pp9HN9XM1zDqjNg0s7pZX/k1KfgPnsnajU+
MBq5RqcfzhfTDR25QP343rcwAZHQ+2FP7fZek6i9BcsTzlC1yFg4158ZjE5tGHW+
/W3MVDYqCnEn1nM5cNdTEFuXhGNlv+zPw8fU26DuByvz8+xcgiRQaPcOnY7AVYld
odZHVZ7ObibJuIzqlM3MeplwiW6U4/LQRKy1m2TDlyEpo+QhVtQIvboPzBzlLjNf
Ov24wvCO6YieTFKzUIRzCaDZyRdTqb5W4lA9Zih8XG6NLTM6ysZGb5BG+q0KtxT/
J8jzmyG1uApcBKUVX9nosQHIJFdZzhbdX3jdJuaOTSyt4Qd5dHTh7GlVD2daI5dI
cjDd4kEsfqiNCgn/NuYNXYiiv0xe/tdsOe+k2s4B2T4df1ZTsUw9zyek8VApoJTW
EDAfPpMbexVB9WSXheWRH7tqdbJhSXdfx0ts+KBu13O764kbze/BOkZ0FumCoWee
//EEx95p7+NXGecvWju4Z+PbtKuVjlMjaB3ayUCYHM++njF8LJaXZxCW2MlI8oLh
PnfG2W3vaOQCmQ/a9chTpIQQMcYT0B9btyvlEts7BlCyRnSjMavEx2miOO7swKt+
9M8eKMCuRFETofZ8iZhxrZ8U8CiyeSBqLTTuVwS0ML3sz2OmC09Tt5bX3NJ0i2Pj
Wh79gNtleeeaZ5lSsM8OFXB3pFPK1zXmVR+kMznqGj1s038BX2U97yaGZIZrBKKo
JDjnG63yaosCUqYPQDM7JAuURy5PXxM1kEWJpwgF61utkUXP9rsMrmpPf6iq+0Pr
QjmYc5mj34f7SISL6PrrEimJe1wEiWwRqqjCOgM0QvzfYiUUUbmys1AmGzRZ5qVt
/3OT8PnrSLf0TO+3T18wHn3N6pNMIL8gsWolB44w5nnnB9UbwmIgUsAYbqV6wwoZ
djygsXzJlFzkXYeLvDxTnIC0+Uvx7VO2tG+3Y+eWjfFspTANDqly6JGJX9dnrzTQ
6x7p9T15X3nT8Imx6X/A71Iig+QLxORHXVt2A6TzOR3TnK7TorXzIXS3e5jSYB3b
C/hdVmffBrnRCPsScvID+rX8iAdjP0mNkOLTBB08eBYTH4QR/TaWHFyH52yEFL99
msYfsuFhpfyvIHntZm29cX2TLLYmsSKmYovNs82c/UxXpSHC+4gCfolACRb9mNxG
DopOU4bcXkI8YC4gHZr/5XikVy+KiDrrbKgzvXm7qZnl38WkrN6avFikY9OIpqUC
QifxrxDDueqSt6b6qH2HBIotKqTvlgRdjWRL6D+3At/lL4MAqJkBS7MbAw7Uh85Z
4gjLaroY8CwXpe+Bq09TvQdf/Ky/SlIyavBB7O8faBDnddE/62Jr0Y1C4Bb6DovH
vXcDzIRzyNsxV5tpGB3966DN9NlPGBAVvT8b5VSi2REGP2TFoMPB9MRqieDy239p
Eyq1fZQC5q4s9tO7gWHJVLXD7y1ebRDilLVREkv7vbdMUn/I56ICmK2Od/TjGY2Y
lE6zgSWr1WUiAj65OByWPE9uWgm+CSfI99nxEwW8COMIUbZ63IPFwTKWKgsTm+XR
UDs/SGRnPhwNZQaAMrCQRnvJq5yZHrF9Jc5s4ZL2RQU+7j6y/Lr4MtdQII9U+ERC
1apsJEbrk0tl7ETyrIBaEErRqm30WdVAoQoM/L1iC0nilu/GxslXhczkv9dS+2Bj
0niDWpguEekV1ZdaofFDado1tWPlFUmWgYpKohF0LeGvlRswE2dDWXpo5SKktGqR
rN380Kx4jxeFFTp+1ujQzOIO3cbczvDecl2jQoi5FWIi9P/i/1rkjHQ6EolZmHle
qNaPhSPflIZJLgova5XWDySP6hOG26oQgbWQM9koUIBIzt0o2JsQzg7E9E4HfhOG
v/BbpwQyj0h73zKwCGVylc5ZTN+u99Of41C4ReDA3e4b2fdvmcTUAEjIxQdoYa9n
mMiNCAkIcnl1RrPTnZetT3t43x36yK7UC1H+9RH31NxEhXukY0WqnLRkaLdL0N/y
vs2kY1wpCRuezbLTUQttoYOGWR0KfLsflET6O+nBEM8zxI0Dji1qfAMfeiy38QsY
S7T5DJ5gkZxCnx/bA3Rcm7v27VWdYx1WBHZd5NmTiRUBXLMX1aiA0AeHGBXd+hiy
OKhHNYkXZQSHtQIhWq846PkP2hGpy4Jux6REljuOZDAdTL9WFyaOC8OYTrrcsGk3
h2mVMjHOrfYzj6XXpG5oBhCxaQ1wHWMLmSVgYcV9gzvQivbKc4YwfwaOCqoZVmjq
KSxG6IE0iaaUAw5lzghWagSOgQRU5y/uO3U2oah0St1Kj0Beh4i73pHlPo5ORsQm
+ypljGE0Ri5tFBdgRxo1YGto9MuI+UxpMXykrMz8unCT1QhisFDx+4j42AUjcr6o
TOxkuswhugrRIH1ijqly6zBCiHNfnRz7bAXmxnraX5meIScu3CnTmt7/14I3Vp7H
NqgJPb6x/5/TDafyFT+Pk1jjz3/CReegP4B1eW+v1G0nHF2KHIuS4gUs/ii8vd4h
zLWCGp8i6IpuQml8uAT0BHUskgKAJ9K42YOhiBAARacEfjqnMS9+tG4JwyoajRFD
J8TmQ9hcMZcV8XIWer+qmtYTlnAYepCzV6p+J0/FgkBqYMSyoQt7mTHuqU81/GmV
DhCwFeam4CjdGctN+lz1d7IEFxLt/lQDx/EZWVg6prR2Qz7t3yGOKqiLSteZxHA5
8sHbbJRXnE2YRnSTHTAJkq1gCkMkuG0PxwXm7tUqTgB3WSl9Ys7plKAW7wzvggUf
ctBAsTe3TqmNnWj8+7mCds0cSXX04P1YagToDVTdQ9lT+jQeGlZGvgvObSr5kgcW
nUj/p9ksihMp1VN42nnfqT6xcRkKU6D4EXGRtPi8LzpJI7O/hVdeIWypntpiykHH
Olf1SZpiWqUxwatSj1ZZ9+Mpw9oWGijR6jNkKWbspR+/fJ00Fjr8qvZ+5XDXX66+
Lm51ehqIvIBhLPcPgdnV5Dnzp5DgZmzQgyDTdMSAIJSzLMEuOqaOd6GxnLcHuimz
e6huCCwZCTgiO8q1GH7ERBKkWXw2R+h9K1eXiw6K0GLt0wknMpTVWCEP+u6vGOXe
mRofXZOCYFajCJKQaTVz75kf/Luo4nvxOzg1GSAxVfRzj3IVeS6Gyuo6vRKW9UHu
j+NYW2BSExe64uEz6uSTr9cunN7KjTgKquW7ZkHdyXEEdLgmmRmYYM5XKh+TfZm9
q6QyJ0JhBxzWHAwTjpM1cOQOCnEaL3eGaU3L/YXINz4RYFM0p/LbIF7di2Zu7GPY
LEu8hfi0+yPXq5M4BKZLjTmv1RPqG4VTklpvvXKc3320msDlfMYLyzJprlh02SNV
EteG5YSXwaMgI0RW60Hvvs2U7Fgx4YSDHZKLNXheeZ9EQXY/jy2SvHrX6io92KE4
/AxcEKF5gmY2VIe1HHMzt+IigJvp2BwuLM2rQYOUqML6ewIjNC3sXtOEY0jTdrDW
f5Y3pi7buf4h1OJwE4PWAT/TxSiobAhvtx9R8yMZuAGuzdH/GxPEeXD+g/mdGxo4
vwyERRIuOOviSrcBnvMNmnAv3wsNJWy54I2/Y/duHBnD+h8ZeozCy+mNTTbKl3o7
d8gEM2d8Y7r4jvYGLuOxxmEgWa8BNMUA0SLxN0jQRltkNt/tXHUqGuStWkYAyOxF
b7wdNfiNCRlRryzdVvoTFFZfKDUvh5Xl4N/EGRAJ5WWF1a/bc11jqzvDploQ+jCA
JULRz+kHKnp9Xr7w3KVKVN+BbEsUdfD95rcdVI4/rstoFIoiiZylh03CS8eKA4NF
ceT9an2Kq4JDc1vJ6aWOTfIUf+7XDv+CNWNuvIEpVOOCIoz13GCYsQIYq/QbJDsH
gCH4Hfpn3g2xJp9UZoj3glsJSOkDufrd+oXnXZs1/PtJaOkyQhL9d5KYKkLhLzTh
v74hymT3meFBNDShvzuoahQes5R2ZSBDMIWIhzgAmZ2xbMhIgZCGXXb6jg8JIKq0
V4Zd2Gssrd/wVzkpVhJorcBcfGjW+A+nSErpZ/FJ+SuJ5L9hJVYaTeASEYgl+QcI
qDcKxGA3KtpyZmzBugpTwqn4Di31ENjnyi3bs2MI5o6mzQ6dB/l3fHHQiBWdRR3o
0TQ9G5ck44+pz8KjtiVu5r9DGSWwvToFPGMdFxREfGXTGBGt6T1BURGzK41ybD6O
AUfyL158gGaO7cGKQUsPXzYloPOH1u1IJ799t35Uly6b3GzwIZd/lkYT6NyG+lBD
2mxbtiVB2CinvFsYPdST3gWwbvLZNkoKkfUEJDWmfTi+kC8rmchJ24zser539M2u
8mOaDta4CArCHdLE8zhtvC9B03LnLx97S/o5f9lCW0dSoUtTzSwAkO/2ffaTIzJF
5cWCtC1GRCWqZVqbZff0hAVzZWSQXl13sTKq8mMvQnPxH9I0xdbp7pd02vYGRKKx
8SRlr55ed9bC2q7HrkKGsa0quInGU+RdfopWan+/KNZmDB/y2UjvW3QFsFvF35VB
60K8QOFnolnMmolnEHtwYk+elOJpGw7AhTqq0na1hdBBDU27XsTJmUIkUuMlgDsM
Or/nGs160/6IbtYxOu9VkuZd4EQg6K9x1Diq/HvFe9akj02d6ikUq7d9kkijZxVP
avb4E5JLJOSNmF5GMiobYUFnQe6SvaRFN4GzuzPYsTLBKpNH+sMsQVz9BjQNaBBP
Iai74bLneXiMNSxDLJ3b/KNnGKw9MFCg5BZr7oHkyq7Fm7Y/H6/guI9LI+zz87cE
tOu6ssMlbyL7Xy37XzNBEivrRa1lVevfDd8t+NTayVTLPf7IjBr0TtzjHQYqoMxK
my+n7lYmYMCfhO11DE4sU8TAq+nzmeCAuNolNiW2Gzr/1xDU9g6UfaoeK/gKXk57
xUSYozv6Q5okjqlnx08gLvBsq5Vvo0NNyb6KcccfhH88Wo5InOhprrliEHY7LtO4
yvHADQgsv4nVFDwf5euybiW1e2lLCXP0Kdy95DZ61+zeA7FLP0/i/ohrepXKE74t
mv00egFf6Xa5nply4FchzBkYoFUHVhKxdd3OVHaDqCF4KCzhhkvBIGzpdv8ldltu
YtCZ1OUYQjHj0ocbAdbKKcVNmtg3CE2cytoARJAhH9CZkQjJ37hrGy+1osKrRB3v
LvY2adQK75yvZlCUpxOeMuAsF9gRYDuHPL9EJkhWaGdicVaY9meRJgXgpo/nNTKx
HaBJ/Snrug6DlEDmsmTZVwujp4nsmjF8U+HZSqvANCcokSO7Qzd6DINHP/XmAqba
kawWwIk8UKi9yhgg9/GebI4V9mN2w6enNDIPZuY8XVKIyG2fJYwK2fqt/vugu1RW
NUaBDBxb/RNtVhefQExpMJeC+LvAbw579mqRKXkdOjEgRseG5iOlEAu/qdoLKmu2
CRHLYsrc7asPGlvjNzY29pGR0b1zRy1/Yv+UHUuEVpNg+7Sb3Q5ovd6un0djGVl7
6Gh0RLsZFS3xHRrNhcobosPVtKAaRzoHUoVgxcecISOMKDMf3sS3hflzbSw1/1ye
V3MIeX0Hy2mG9xn9p8QnpBzAvR8L73U8/piTifFBJrTpB66jHSZIoTaGt2AI13HI
QkGJ9sHOLIM/bo3W5ilrgPJG0Y7uNfFJ9Eg+Bqfl8SASev2tr5G88oYa3+3Jh2Fy
ZK/mArt0W1KGNCv3SiWkRqTEtf+quQMaiF199656itBt9Bf6SS5dC8FXSe63X3Cg
EjmRDHIhGw8S+0ZX1mujwa+Pja1AXu+4A5JLkRo7xCzbkX+GDRJ6/iA9Qf5GHiQN
9FggLAnlydJxxqpRuMPzebJe0wWKacw//J2X2t8AcGVt9z7sGwUfvEMO0Sdf3eA/
wOJSGhrXUEdhsdQhPd01bN4J/IhjEyNHPfQe1wn8uABQQ+l3aGwXBRT7v3TILjrc
qqPrep8HVBlr51wz+EM6uInyDw9OzEvNtC5hH94pDLw0jTX89H4hWNnAqxCG8uHP
5PtVTGbZtZ1/kLHg0HAKwYVA9yjM5+es55KIM0GKfhfmV46mYYlybmQV5LoY83fB
fgRdJ2KSdeSNuPWZnXGvpvdy7vwFIx+aM3dtA2cPNVDWw/T0M5Y6FmcHvT3fpZZF
tfpSGtUVc3CGe4QBU7Lsam8MP7obE9ZSh1RMJQCTMirQU6RI6O5gOJhKAdf/W3ev
VMxrva4Vrj+ORrBzlcivuRyQwGzAkyrM/JlO1ag+kD/MIpqc3McSJTKejudYElqM
j/GPBGyEcWsRbVRzBpJ9UQi6bLh60ZTIL8hhvZb50wZLUyUO/JlUVlWdInVdhJJG
mMNCKMEdau03TmhqtQwXfdq+RMZ/z8rO7JhzqPFFhemDg78tnYnGncx7Os6I+d6k
PMQfhY6MlYh+gfZ84l2YHEfWaJ9GPl3qUvI9HIhq+i4V5eaAzTYJhh6NUZWbJ0A9
58xJdmdvGpB+A65aY8Cm+BUKOw8mJ2gJsvlJdTRR3JxT4TZaWcvlf41s79flbsSe
cawtmyA3zwXOQ67JtRSw3T0HeCJhkr0cj+IqWBXKT6leW5NmSKX+O7f1osyIJVdW
z0tyuyJDR2iGi3O1hIN/cua84lq2KND5KHhNu5OutKSXgnIhwdRhpW7W6IpR0sl+
zu5SZxvrMaHpYMpmqarg5/4kA/OHcGzh6WDKf3gSorT8z30fbxO/PksDVk5uD2U+
Z1qK39G0h3Skjm29Cu1uv/WizsZjWm7ddN0ABlM6JTk86Chkfpm5SzXwe3w5dLyd
1KO/rmvrnbRLqIFf6jM4uS0FZMwZnj6TKzDNki68n4UU+gPn8m8UnFHVwmoyh4cr
4nIln3t6Q9nzCBFhLrPPSEzCgGj5LSPiFjJRx/uAEmBfw/GK1hLacRIpG+Oohf9B
ZNUooDBCRPm4Z5BMBM1EpUK5t18yJnQE9A6MCbErgshavqugBzQx8obWzLS8sM+M
1hdeIQxJULy+o97DNMmssk9i2yUu+9ehU1IkZB3N6wnCrGP9A8ppA3PoixbFb7O/
fy+gycx2mJghfUgXDjCXSzv7v2vAIGpfuXB1fSXwI6n2ZR4BZfC5A/7or/XyXh1m
0ifulHghnkJNpQca9fzxwqAYdp1LBeisAkekiEsbYVsd02GRueeJcaNRwSwiLnR1
gfMTqSfAEcdrz5Hpf/wWqsnOnBFjVAfA8OgLF0lXZQ18QPBSHL3jZLV6F3DriDsw
BxaYgeNQhpUYVGOS6pgvxuM3P6v4RLUNt8A6GgKiaTAASzg3E7k/DQxrE7TNxxWt
clZnRE97ZQQXAJAzEj+fqix8l3sqNoZOUTifXugjRYMkIoL3SY8iJJrhmJ1GSSrs
sCq/hS4tEkTBhgf/VaNLeVwtveRSh9V43Vas77nYVeOv0EVPn8zVNyLb1sPr2A8+
w6u3MzF0lgDD9uSkPEfJOuyVrYFIyQQq0gOhcz4IPbBEfAYBhoXwmsLQXNr4zdLK
X6OiRBIHkxTMzfzWu/R+ByqOK6o33kvSgJDBrnssIHsib5/26DFJ/rrWBOhc2vQq
zPTHTYocgYyV04d+bMDQKmPjkicGOluRwloxBg38IwydUi2qUcmOfoHMYA4hLgpC
OO7c479HZjqnN1i8j9ZoUz5rLLTcV5XbzO68XMxIzBOOtWy32lE4Sq7ZKi4V2bV6
3KRypv1lfdJ1abPpuelZjY1v8i3ViVO1Ob/7DkdZrAWWNY0s7pyEIQmeljcdrYJP
arTqAg6X5I/XlaG5ssW0hLSlOilqAG+lPgXpT/krhWlxHeJbBM+zK7RDUW3xCnv2
4fJ6Urv7n7SyIWwFHtPCZvZEZOlLw91+mJ9CO0o65AY+K5ppoErhEkWfdNvkGZN5
RPXwql6c5lJGxFEhpdHeuSnBpFxggumTMKIKCZayJfYXKV9WRn3bhY0TVw4BAYyS
YTdONMFSLoYa5uECOfhtPsdJfGc6SmbjPCFKTa+vjNLRQXeAKRYkGSfZldw80eh2
FfumB+npbKrnJk+JtP5PTw/Xol5BmjtGBrSaKDj4fXrOX0JEdlEzRFpQ/FBKtdyS
bMRIpSi1VI98IWqDGSOha79G7VuTIPE/QHzFJtANFgx4NwHVbjQAhusPUMuOvkP5
kq+gbgB3uGrmrtqqtaSCjovqSCLUDlKGraJ+TuaLxA73E086+Al7l9vQKDTz0DqC
iS/USlX0eekbrpY3BslvA25TfnPxX/lcAWQb/beNIPmsGduCZn0S3J2/VjuMm+IL
9aSM/0obT6UGBkznerd7WudIpP95HWWm8VwsAd6QdB2H/Izr3zAb9Hf7bzaOV2KW
DgpfhtTB1E51BHN55sfT9B/PP8wplj4BjgRjcAYZQpr/jAER16UWvTlayrYGB8Hj
B9UmrE/pRxUkma+YRP9OUwFsjmG6b6wrxl9bbG1m84lCWYMcEPn/s5AqWmEOrAQj
1lwOL16udmrasjLxOkHzeiT8mFdcaAKzE3+nedEP+Wwi58HXULacN6h1XxdD8hoG
gI9PJ+nglaFClRJw+eb1c8h/8RZ7A7yr390xRDC749mxmmj5p3j5By6E5mhAf3G1
1l5nUItfpaxfmwzsqxqNRPCTHQ2lb/+KFuMZ+SAiS1mULH7Do8Rx7wwNiakrLkt9
cj+K/k3AFbkYhc56ZktwNZW61zY+i+OVzH2yiYBP0xCBvmq5G0xx/aooLOoobpMJ
WXupdJELYHSZzDLuYcM41Ohs15Lz/3wMdocEkNiKGqTrLrb9ix6wqc5xPvH5Eas0
WfTbf2DCcUooWtCQWENu2X+bLoYikZn4jQ9MO2cGQ+lCMY90RRDqm7qOTssF041K
Z79xeLZFJ/akm+/P83TRxpG5TQDB0RFJ6ic+KvrA3vfhF+xEkzIy0mivL0Lr0Tjn
AZaS7q7MoF8tWhIayXw34Uo/Ecs+4UFQgiB+n1ivO50c40BN5eQv9xViW1R6jE4v
46w42tbuhIP0rHir2QjNC65r3wTtEonK5ijC5X+PgAnwczlBK4zPVwIbP/xzskTf
GOkKFaTGBeOug/WWIMQBgVDx/FSiggoeYycQmsmuZk2fH3Q059Bk8zj5UroGBqbc
nM75q9PB+zzhO2gjrlFS6pXU0dyKDMenoXxBcpPy3ky1QE6428TqLD6Y9sXYeyac
UYnWaeqHPCqDeHG1MRkcjlir5QkWI01gHkNYXADg2Bp9Y030xZRAybTqWjvDFNQK
bHJudYfnevmkj8TX8t4ORpmQA1Wk/flXwc1cEtyN/5YL9p38gr1YEE8ipNAB3QbP
mEcI1/6oXVEvN+W64EN8fRpzqeD9Ae7/BxxSLrBPlfE6RMYrs7IHLcMiYvOU7tGq
NghBIsS8T/wH1Ss5UielT/CiE0YrNw3dKkiSlrEABvIdcH5ZWkRkwyRv7vZ21t/n
EeRMeAvaOGDP1BcxOqp+OinaVO/fOaoegVpUxzM2sPUlTT6jyYgp81A/OgfUaPYv
SIbHEZYH5qmQJCyQ6VHWnf188W/Jp3CX0DZGemj1y6qYcxzE+7Yb6FJD8pnwgeSi
zSSCwTAYC9zIYkQTaJsDVnCMKjJZLTGQ/9qPqx9AyZK63rjklnXkwJ+oko0W815j
YkCXZiPxM2Nksgqhr7QoRwJTGO1DVsEyYVqiOzqqJ9ZLVoLIqLqW58DPi3ZKErxI
9pc+8rpvmXKqxEDgfZvXG0rYP8YRgVoAyJgV3/oFYb/Zu2MrT4Q04iX1+Ur09jHu
yxN+Em/OhKmCkZq6ovNYcrPDqHTYN76Nipwu9SUbCUayRylIWsnMrA2IRmHewoPJ
asxIqe1zz1sBhDR0FV86HrD2vRlLINl5NqRnUN8Ww0OdNTlqmxwyyfXuo4iSiyFb
C/9AMHwMcJVMD+/SqoFMpQMOUGy+eKShhTueGZaQhWVk8AJRE/NYYodQGN4MN4TR
Q+/YHvk2MVRoWvNofIFHBPSARWTD7hdKqGD47b+mSgRW6eXmWNP5cqTq79jok2PV
P6NoIcUgc5OMo5ioT3Ow1yZV5QGD9CUBQNqTJTa0jNqpYtQHnXSAt33tswVmfguT
Dc+mO+P/aOqVOLpOMlbG+KtB8fvaGeofcc2K6KRljm2lwGDjvnfTfAINdmV4E/Mt
17aqZTbjyI93pQU/n3hFao1IsTYA8JEM9aniDgFidyT4F68FzmqTNP1A0eZ6Zmh5
+9Bslsvv0tZNR1IB6Mt7duPvzh1kP4/d6oiWvPdibg3tQPj13SJuFDbo2YuvaGwX
/2PH8BNCFaibVZ4u3Z1f2wrZUvtROe91eYJOqyHgY7L5LlazT+wYSvxCeX9XXlbx
EMmgmjEAoleqn18anJb7heTsoaSujB8J+JdnLsxK2wRk0ejDLF42i+5fjG3VIEdH
nkwadQQqY6KeJv5LDYyW2G/w/QIWmChBwM0q0JaO5A1PdFuNHplvb+wyvtOfaVvF
ITHzHBDknL7FXtuom6kXKxzYHvZ/Ppu6eY24ifUfkF36lWCMSi/7ryqOaRwYuCSZ
tBqAe+yHENeN7Ogiiv1A14FUMJtT6Ot53cibY1QukwL1Ks0hbDneVgdy9bFOpvC7
qdAgMROS4wPgPV6G1Wl/5yMpCUhuTqg/OQAOFqp6dbCotyT5M5hl0rudMvPQJK9s
k8f2gYO40y13SeNe6Q5P7EFrXD38jdpfBxPNiJ68Fqr/3lbHrm2dUMp9R1kAKPqL
6pIROX7lKBkGkqyDkRvAcA5a83vnxinxolO2WrJP82UMGYd1DKBpjEQBCAm1awec
yIqvNZ1xgihnRAdTdvwuPV+UjqrSrFhZwgx2B7hRGGEjL9bK5iu567rkcxTbxjbr
WIKMHzqCU9PS1NGIEjDLm2CcaEvCknxx2Vy/+tlBH+z6uXnr2VWkcOcE/IHtDpF0
Arye++xmaRgRQ1wGMIM6vngE66UfevjTwQi7G4xvftz9xzaO7UOe0sLPefFf+rEx
V8CSfj77O/1Uraca22D7oZGy2C30TnYzSmz1eeBJZDeVgteTTXLqXV6ZV7u0KhGZ
CVIjOY3ks/sirs2j/sLIgUmyevudexvEfKmjUihscCfyOVpIH9meBWYPnhnGx14i
ySL1ksd27wEEoO1giRaz/lwIUu9vXVnO1Zk6vrg0r3Lze3yqpEWpQVvAm141alwK
Nb7XHMVoI1It8L1Jvx8kS6b+rzz7B2NmrvEGwqpZ/4IzUwLxZLecdpl57vgkCWy9
vf0DMUhOlcU6AFTmpJ29/kX5tSFmo0N1jdYZSvdDHiVJuzxqcXKmVPIptQjQ+3V3
YstQAw8Q1ThjvfX8nqP3jc4/2K7fREnXpQl4hQ1Mtnl9N0Xlvm4+K/8M7nsSLQSy
TKAOrkY0ZAJhosElpwBUAI+rSMQUluAiDdoHe/RRYhyUFPTPqefiNnZlGLeVDFdK
UenuseaMj6x84Ztw1U0CRYK1dvEmRk1K0WUtOm+MxA/zqfhnkgtlA9Kpytds9YHp
yw6vG6d0q17YwLfe0qrDNrc4zqednc28f/Vfh7AAq9hAea4QI4PKuGCsa2HZVAIQ
IJWr5Aw+68WZFR+DEISqxrQk+K2cRMxDRlcjmnqHzl6aVl+EDpZx7NGsLELvvit7
ohDtePBl4NWmGRPBEjq+scejmwqqu/LYWI42MI+VmphLRMVK4Ib+zLAxtHi5kV8r
aUB020MfEC1Lxvjd2jqcN2N1FmkpLuFLcDip0xhvEaOt3/mepxYWR7MON2bQKRGJ
9d1UDtM72LERI5irlIvsRfv6cIbDJDbtdScFWjJ4YiI5/zht91P3G6Dzub5OiCgO
0VF7ToHSDvfWIfI4cGuqi+nwdLvNw0Hc3xKx0L5pbtpTGczrVsLSLFarKTC/CcZn
mXsUQafoYRfddGiigZoyvoD2eRrh6SYBdZfL0bQvvsm1nusmbkPVwPrIHv8TYTFj
LUaxo6jJLQJkNZy0+81PzzSK8aAsTL438ArvgyRM+DisAAFTXgBRa7/cxIMluWCc
3zwjVu/cPkhsgINUxxV6WAyYl8nHDbCkKUvYxLEYSdCw/JAYMHFSSyJ7bhxOO2aF
m2hCaiYfqrGtAedrODfc65sR98bmfzcf1achv54szsc3uB0w04AfGSyNIm/WemFk
xeU6ORdnThP5qsr+kM+1MrVv4Z4HvKlrqwmVxeNXfZCshh9euvlqqVWJ5xJjWQ9n
S4QjAI9ktQD5zUl/IrcrFXo4ajJObQiVBLaSsU39labcEiCEm3vJinrndvtnR/2l
eQd0fYMx/tsxrJcm4tfGn1at8FwMFNROEelCb21Jrzttq1s7zUXUe0moWAVxNFx3
FxbS0NKgWlEPE/HWtPpr9c3Nk9r2uSB0jApcyPYNzh60m3rhwBbY0Y4Wi9NkZROQ
8WMA4BKKv/C2ik3lx54o0UxWODeyu9GPtWbRqSJQzOHR5tIITZfLiqotm/3kiUBQ
EqHJe8hScHUT9/d7hiI4lE4IMYtLSeJQRv7fnMsqFV/IjjE2Ns3Ui550kSHRqBiH
NhgS+jxBzSpNNfIF9Ix/gYaDihqOmgFjOHXWGsT2i47NfMAU64uoA6rVVJTsyolQ
N6/41BiHjUyEdXNqDS6ta8WRX0I/aA7nlW3huz4Ay0MoB017mhgkOHVkCgoNCPUU
fLhC4QZpapZziSs5ptXWGah3q/rq5QBb6HwSo1naW5d0w1X6/8dtIfLmbTRgHTqZ
6X6lDJm4BgFEdL4MtjsqtNK2/z0angkNo68QfYROorBdlgDCK1cVWFWunbnJgkCr
wwthSx4A+1Eztq7mU1nfTNK+gYpmTyc6m81aZqrmqegW0o+R9RzoJmBqx7Mz6epz
Rf8ftrEUca+kVeC0kLPeXTPGzvFkRsXO4FEzs9j+Fj1jz5t/lntd+D7prCS/w4zy
cSn1jolm1dD5itcVPFT2xjJLWDalYBHU6N4R/8vahrV4EyD7FKtgkBTu/DZJdRvN
0QlbZeSqWoQSq4hEotNIP+iRU1r2YpPRlq9/+/4zPlUneTIpnJUYRbQyDNLzrIvT
5suO6HMErI3J5T2FKWRknPCsQOF1JKncj96to75LnLtwUNpDr8pq2AaCIFdxKJa6
mep3DDWRN8V4rRRHhr5kUGGTUtVJpvThv+hKptgSI6uT3pGZpdjTKxE7ylF6EAyq
7txVsPXkTQrw4X6ls+g68YIS6FeJbhEmxJ8FzwnnlbbSp8iW3022YW4xuCcqQDV5
sKn1dz2ZYYnO9CV0+J4PuRs9ThOgxC0zYc5pRkZz/b2SnjdEMSqfLwYrrSMBuhqF
SdYVo4IMfniFVWQmAPnfcV6HDj56MQo4A8hmhUXjB4qy0lFC6FrK0g438S7i9ZKQ
CDRLDWL5QhMFroOPMk4T9SV9i6GTh6Gl+fWvBWz5Z9xFsB0dhObuH4jRT+E2Q4OL
5SCHplyumrDP2xbXq8OForRP5yPObDT++biDHTl2GIGTR+GcP8Gtyiyo62WIsZRA
/FIP+1bO8mE8GQgwBvSjUx/tU4AkbO1HvyZf8/a46LLZKmwufhevBBRR8NNAWDiR
xQJLYHTG7qFk/cv/TyQdM1PG/8hEkxSfB50k93gKkyQXX3NlWI8RsOn7OIugDCT8
g6ckktpureuNpgEw8N84FMn3yUCqew5odDkcP7/wQ0l5nUVa83IIcMFkOxS/TJBp
myVcZWxwTHC7LKVbz+xbzs4+J2j5X/VGN+NiOB2l8i+gZd09JjlaM2x6HZFSyOCr
nNyczD/81sbaGlkTTZ7cJC1lKknWF0lfWKOVweaYGKas2xcaa0d36g7oXLuL9pGS
I03aSaQGTAQ5ROS8Ls3jxwqCYzC9/9PZCm+TEUCmenPF3Uw8Pw7QrzVRdMYc+QKb
cNJ/yydixOfpu87RQyWXrpRGnt2BP8JfZ2g2cgx3dbTsKAegJkZ19HPXeMVb/q6H
0iWF4RGv8vVosXitBWBbclM9WCt647NyjlaMWpjndRIwpDfgV6CQcfGRktgH+0RL
po6EzvgG3yHavdpEPMU3APrVKMvZKuXe8GEACs8dD3JSllxV0yXVzFUEvZw+VDVj
ek5FcPDziVVnLQOfGFKaJ6RhWRoY3Jkr3PEk8K1raVIInqI7h9xArW1kKUGyhnhO
QIJ22cb9ntoa6VSUFuY7bS+Sh86g61IDYp9Z7bmNRBN5yqywLz7mrO8qhzAr0BXL
EmWMiboLbH3icJ5jg+tPUvsxIX9As6dmcHlxJ01M4fe4Bkpr2bYc6bVrRzmQAdZc
/8whbWjjtBanVMS7QIvpytxuKUR/AZ6pP9HhtZjTPxhCWpOtxyKmbo1TS8gqauad
NryCuJIg8tRMtijgz2NGNpjN8DAhbFmh0O+RVcWGnm8P0k8KZweDRhagDG6VBrzJ
SP+rGWeKS8MmR1YPBIcry5hFKmYsOeF27DrlNvfdCzzS/QwZtSGWhZKLoS8luSVq
KJtrOgjenU+FhapHExplAid0WKYQhWwO54z9R6Mng9OSrKvp1Jx4krkiyHQhUIvI
uMO8KNv12LF643SbbpNymcbn/We5OfBh/SOJzmB3qf5NH6QRSjAnfMlrZf57IKdR
ezJEqqTt/auT9u0L8k0W/+Te0Zwx17B59LgnFTyKIE0iTOWvD9U6hUURG55puSpY
/fV9mfwVyrgYS5v5NlgfTCsl56witY3d8V43iUybHw7ie0NlN8plPhqtum/vpwAZ
vgEEGVmxSoc1uhkFkR5yv+O3F9fYkF6nmb7kY1vOtdr0NW05t7DnVU/83JW5um/E
yR2+IRmkA5fej7fcL56ZwgB7uyFIbB6X6CeuCMSA/leSu+RVGd+FdVMI4Ug79ltk
5oM8DxnfaqMmArwLCU6Se5wT0BaH4LiEkllwhdv4tlCKVIli6d/F1dYdg5tLyXtB
qDS8l1khM9Q5/5VUrvy2L57/KPC9+rhY9SUH2pv+LS8SOHRL8PXcsN61Ekf4bAPA
g5O1WoTjD7+1Ani6N9HpoKqXpL9PsvpaQlTKTKTFpP34haL2hmjVPVSbPGPRwcFK
Lhd9ApBRt9Ni2fIJifwgtWFTWNPMqqzLCh9qNcxH54/d0PyreVaLfqGm+fRRt9PL
UNbP98nDdPIkq3qxllRcmeZAQXV6zLrNJJ3Nf3FQmD1Ln/EW+fEn11qhw63ABR8M
xnbtQq0zJdNQpj53NOJcECuxjVrmNRmeyk6aem5uDnl90RhWC2EbC5lOIzJKMGNy
frxyEuR9tVoFter1DjWo+lDImb5yYvuedRANjS3b8OYGp+4Sjkzixu9xQtEJs3TW
EQabu50PcWdS2nphiUKvGhHDg2VXnBVbvIl/mi9EwJLvYPRq54ToBsp/b+okCpWx
iwrE2RdGKD4g/CwCI4dVztLVTxdZtv2ipTcT1ACKU+oDoETHmWk2edhNQlpUZwHb
DO2EzILedsQ3Fz6RYtNuItA7x/KHhbWTAFtt1tqOdEZ9iUDOZUEqh7JJqnsHlylp
4jqZUfkYmTI3r1GqvgPNqHFFdj5WwGa9Qm7PVW2cN1xKm1Yv6ozeEqwQhE2HTV0B
D4QKXo2ECHHGN2V2SNDpjAbun4KH79eZcXRCvAV9uk1+RcgnNcKN36Nwkq9n7WVk
kzRjWERTFG4RsUgge8zDu0PSRNoAIVDByIfowhzF90kv+IjWkYDExRr0+rR9CW73
NKE8lPPPstw2R54h0TSTZc1Nk+gXmRy6JULb3EPIrteZhl5q7B0OzX8Ki96ejPE7
uEka9jkS8OCnYwXRK9tgJDUgHabLK/LSGXMHyC9ZyRbRCeUin1ASADXsxD4AxZqG
6OKcXBvWYfd5S+p/hAzalgxnq55QBvt6OTxdATwh8sGVpvojFKIKpzVMSjGBIWYC
J5a7WP4wqM6yT2cd/0kBPbfmiJpgBKZZMSB9wKxDkt6ATCuWWtB3lglNWN9VJwaj
iCx4Ok4jkHWf7whKxAqnHvB+8o9Vmsy9WfFFCbKybB/QLGo0XD5dNbAIpWv9I/aX
k8M6Msa8EtgFVzzTkb9dkSt0y0ofwBCrzi5VovD1Nm5I1pq05AT0qQ/kyqBDWnkl
p/jNDum0egmCWK8SeXvXVVP6R0G8acXm2NTl9sRfreHKdISWNmP2eXcUWJe6wVoO
5sMz58/OQZuXjoDzdw0R3QevILALRBPKpiendsWI+hyB+ulpXukHpN2ZDQFFQ1p7
ysFTxIIG51uxLL7PMUnv5nXodLflVWu54csm03t7pjUz4IM9FSPvq6+d+VCLlKAt
6BcDr2Cve0+eaTNIOscThb1lWUgjfmmPMByX9ErxIJcovbr0fOl9ysPWgEw1OIFI
cSkOb6G/oYQFHe5zEU5qOYOzB7mB7Isf9N4jqMEIUYiJm4hleL7pjXnc6WL8zdPA
2pRL7QVU1d/fbRNntyU4RwcAaAC/u7fCuHUzsOy9SBVsANwcgLcquy3UeTuXe6ZS
kyH3+ALNUbhy6+72/tD7xj0whPELsk6j14/9IIhY3t7l9qPLMg/pdiypEMHN1bbY
g78t4cS2GhISJfAntHUb9xL47HsTk6tyRWg2pm5o5353+CcQNolanfrZQrNMEl32
JAj9mCRAoFhEZm6sJqK/7UhMhxPxFzofwD6XlIG2ifj15viLY19dqtQvwxJ9B/sc
/STa0qFow6YsY92dAM4n9o/51yOAEy+AcmhqU1ab5PT/OS2hS/hAJZSocx+TXukH
swevhnpwgxZs21Rx0DTVIUNnmgMqtlseSoRW3NwBzkKfKAfVezLKNlpXegmtc4AT
QQrj4ICfIUF0BMO+r87ZxaAnTdk1ILefAtuy7joBl+LZLo+3XQYTZYhU0cjrxVW7
+OPCQOuR1Vj+nm60hqsWo2gGoQj+fPlwXLV/GbVP2AElstmBlQe7fgCUpSqXIwIE
zt6T1hm9NO8IH6hdlmZAwjl+JtIagfA6t0+ZNoGg/r2RaUGOp9whKd1Q0eQ5uErn
hMBD2StonwEsXtc4h1dSOUjUGSc4bC7zI3MS4TB2tlqFwCKTpBy1ekcc+qTw1Gxm
Is1zTkBVQE614w/9wbc0NRRIu71mmCJKsilZOHHPgyPwJXpDm7P7UmN1v5MwWrXv
BI85AVrKfGqTn9qMJx6d3OUN5B6GJR/H3y4fHuSkZuBp/VqOnrSCeFGh2M0MBglA
5fJZFlA5Rzu9mkF7ak1PJiPkOjNQdc/6CyvfEsAXebBvTnGRxBZ3NwbXcojciKEF
QjgpuHwIe0W4X9ayLlyENcaRW1403rIuAFybet6nK7mO4dGX7NpLmLri+rr6wdqS
OvflgONzTVrvfwZMeUDibXSQIXvhFl1jdjGrE5+2juI+wMmA2mqe78uHY30jXGHb
wzzj2CuZwMGARy3pzn+kWrtAPyZcNmg3AOCm1/IOUT1NTCm2eQ5qOTh3VrVGvUfl
C0VtxkeSwAi1O4dzY6akh44WlpUDlpAXZ8qObvgw0XDT/fZofQwJjgvL1D7jWcQ3
dkBSxPa6mQVyRSfmGcwf1IMrAYksZXCiwkPu7vbLY0jGOBaHTJeEDyOAvLfvFDR8
AdYxHqs4HMzwlTtpyLyVv7HBS6JO2bS/kZ5kS01Qv1Q35LDGST5ImbOvH+qzZSNR
Pv71E6hKFNFWLRSn680aOya1lUX40wR6JabHMhCJ4fNnTjNFS0/R/kpJhkHZStBo
+3D++iNVqV9AeQGApKdr29xKPJcXxnMehmZRt4WiOZkhT5DPdcbnGrLbUV2E6KsA
x4Z9t6S9hGq3mmZ2bF+SITA6ZBfVV5rERi6ZmCvRrKHUmbIS6b5MKjLeaAXlvY3F
G66T7uGaTu9BsSHX6PmTI7BzJyYyklz6VpTWRB/JMBU+yK80BlkHUOEknwrQATQ3
sjJEqm0XLohPV8yZL/lr0vlaGrXtFBBb+Ym9/8qT+CPmEtg3H6ISuFbO9dXBd6Qg
XJkbm82kyQPfio+IqOm23Rcet4FnuMM9d6iSboVUmLjjNbaqv3N/0j23Dhd6grs2
JkSpp5OW2tcYuXVNjZyBLFqlqOE0s+6dRtegLmGUG5/LHCQmI9L1zHqNufCMaIQy
3KCAhOIzYrf66PUtbY9BF30Dyc4A5ZvcZPAOI51V9lGqEq116LMYBlloMCIMHqQI
6qgcPDaBfJkbVXEyznvUAYlHmYNQRFKiOhBPY/KoFiTfD4G8cw5c1R5RLSt1snsz
odv8S8kzBFuILjmK5UkpCzEgfynx3a/QLLvh8oTRmTTELhkuKfMnGipm93FJcTVl
Q4dPOFC1Bkjvo0osaJOyaUC5bNdX7GhcA/h5MDOC2AdFoUYDGU0n3alvW7XiyQOj
esoc0+dlb/nisA3DMZqN6RX18EONnwVuoMFGDCO+X7ZkG27vjkcorOdq3w8nW+dj
Idy+bQuCBFqOYqxFHTvCChl9lsTFxu2h3OOOK/TQRYZu0DgIrCVZbI4HAPVrQd6l
42Cw2saiONIaO1ZiHbNMlXhqm2TFM46A2v7dU8tsYXGWzN/2zM2Y9FCg4ucWCkQO
r5I/nydprjtCPfi94l1nMBRfSBsHNBCqJHeAHxgSNSzlq0iscE+1zMy5zm4G+9qm
nIhM2LumKwZfhOrSRtuBp5k36BB++ujAXKoU+mnZC8Go3bw8i4S5HH1oiAFFL9Lo
9IQkturN6HvwZ8QKE24WY3ai9EIGpNNEQ6Kjj3HApMYj1LzWPRcif7zmeHkB7R+q
s2QdPEvMxRBMtrYmu0ZAbEz5rC6HAB2DmyVl0XpwWt1ALaJkivXCcXgiZSF0syUp
Rdiox1mrqtK2SOm49/F9Bg5GRe0G8urAkVsM9MxqFbrtCCb/Bth7NF82kqorobY8
H8PsidTytX3hA54rO+qRHaB9jPiEcMnkXZPLKNgKEFMNascVipwivkkzeByOBqbh
9TUwjRw/0rpiFGhhfOrcoXt6k8xfaJGxxFU+mHhKMhyAXrTtgnUWMXX9ub2gkZKI
0pv33RPE2ofz3h+akogCoFs/ammE27NnvI7U3Qhio92pLQWPHBziTw22kFtzE8Zn
21tP/i6sPCJNhNSk863s41mVKbuod7tFEsGXVzJDCZIuk7Z4SikHHguRox1As3Pj
8clt4FmqCZbnNVfDtW/hyjzDDxE5U/1R6boVXBZYb89N1Eo7zM3N3MYeYyT8SkYm
4h5xXsfchNT9yDzHLtIPpM3pGX0YO0Di9IMDmfIlHf2W0xnxW9Qd9NJSsbmMZAw9
CU1gqJq3YckkFeNA8OuAVHp5EKh/NTZv4Z6Xg8WnEX0QJt0N999M9e1H0iehOwFp
DxfSjMIjXneZdWQK/2WRPVcxJ40i8BgtN5OA4XlJtcxOsZFauGokTKaGLGeoUeLI
OWLfl4yyxYeDUmrt5kq5BpxubUZ9D8qe1SygfSapvZCGcfYz75w89Vnx5VYpmF/q
kn0g4Wiel70bPHJmPKOermdNhJwZcWLCiYPHbtFSkErL20IGviUn2FobLTpT+Of+
mZQAZXXAvhgzbn6sUtE6/M/SRH7k76D5gfm8N6RhlXEYSjLxHBoLp2LeSRGRmBEv
mJrIa7jk/gN2Y0Jy/ISoNHUielo/6xJ9N6g2Lwya/yfn6trmvbhzl3HxGgf4djP9
XoUGHAttidw6ez8i630kt7xuAGjSitjvLf2g8tqGauigAypNMogO740RvaVJ7iq/
vAZeePHO4UqqVHw1wk0+Pj0ZRG4hjiuc901bLSmgVdtgGRRxVd0p0BzkGGXqc0ny
RlL2kXeVPZFqVBAfQqefH1KgcGdOgc4jKWanKn4sh8lv/fhGBuuxx4Tw8SBgne1p
sja9PZp5gNjy3kKCIiKWnNCfWPzpDHFTrvL3g7EhIcjpIamp30exZTh0+iWxpsYI
o+E0+braKNT0r7EiikSOFKa4+5+cz9MRomVHggjCBfv3w/U5invSvCllL/H4oLIL
x/I6JpWwSuASbe2zc5HCcbMQQj/2XFsRED/MWM/YzFbPVL/uZytWrKfxTwK+DOpJ
jbPbQP+3bAiru+RftNME3/725C1dIOXjCUb3UzHYmRhQoSp9AxjGZ4W0tLd5wmx6
FRkfhypjNqwEISNI734ngz5M6rezmgrdbJUKegu8MmJ5HWhI77R6iZ0wXZlideCG
J1PCsUqhPgHNPE6z3SVoC2tlQVKF1+OdJK1OtUrKr+Q3tJ1krsKbzTCJQYNcU0MY
8nAfPCihwxm2etg90eerSVdLhHIWf/5rXeKdAzt5TMedLIPqK/IMRvwM7JRFPrw6
2JST6v4MMDXAYn1wuxqXVFpjimJjM3J5+UxALhQoYIpsDFxVFeDJoo4NqBwcNqtu
aLPD94iECAjJuYXP69M55eVGCtiypCGF6HEV1JBeAmeSJ2fhDuPszw+lBxYU4Qa3
2rHrIa0Gq+lmAT+YGI6b/SOW0glzdElTVNChzgEuL8nEm46VUM9+nXC7EY/DEatf
ireHH9+qcO3pQhzFpNMuSRa+w0ZxndNVJJ7C8acsKnJXpevxQz7LejDsGY6zq3u3
AN990Oi5YDyLsxo60+dzh2PBHt946UGfVIOd9289SGyUgljlcfGviLtFun5FqQFr
QdcoTO2jjyF4Hybhxs6dBMv+Xsm4wYbZK3cuV85GLEWSSJebEL3uwzbnHgQB7jsC
5W2Df7E+4b2ygbjLEd+AZdGC9mPB4epFU/GvS9EyXr0BgBzyoHxPsYq8bh04/sc6
pESva1xqqs6uxoo5Ts3lqRMjYrqsz/mOYE/hnR4LrTZVZv6CbAvVceC/6Rw55gyW
jMKLROEyE9aOSD3Ej+edUkAIu2/PdKXIDDd4QuhLt71d+ohNUbMorDCBPO3eK4B4
0JEgqHXiEt+NZ3dFfZJSPobTlbhEhKJ0+pp5ngKGj06/o4KeY8srFbMqT4gab9gO
4tazboeM7OyX0pdiEdWGua9+ZJcdrnracQ1K/PwpT4V6SohYfI4KmPZzI5JW0y+R
dU7d28zTNfFf21p0LhVaIUd0W5zvTf92cHTbkBGlpDHvT052oaFhkVTBjhyOxoYc
S9bWbTAQ8qyvFLBfYgZ5KcgvBsVPpzpnQCARkkiMk70yzk6kAIEOWxKTe6hpe/wg
R1GWMGr1RH8N8oKAUal6if7z92Dgbw1PXEqYkkCpUVZGzyveYixGoXiSUUX1QNDW
/0AllnuCKSpiHgkUeYHfM//JasozX4umqM0cRmobSJxIm5Wog5sfZWFS2SoZtUxr
e9/uU18wPVi6+xoabQm/KXUpJFH47idskgUX1+Mc7uzXIWUJHx6XJnurrMQf0/eJ
4lhYLC/xC9gqJIj7UqAUp94oXB9vPL4akEltK9EucjS9iXfJcNRyPsa9Up9cvwA1
E+X6xyyX87CS4ovAMWeDS7zxJljfO4hoMUmZE4c3WH5tr4j4m3p6Lp2PCZ8Xa9ZJ
zbmw/gQKOlOgT49JgkMmSfDDxkCU8S1tn1Y3TscX8cJNd3l42WUynRkczazohcsX
/o/vvB57HvPdguP7t5LD3BzubjnYVMmIF3RyGjLYpSPD/ynNiPmAAkC+ELzMLVmG
b3Kfy+hmxVAWZMsuJn2lcKUr3c8asPPR7eTMji+Ds10GnV5CG2FTYkuPOX0URLGE
S1oUuD237ejQtLRPTEZuKDgE71R8Us+7jP/mX18rBDzheb2Kuh4aAU6AJbTvdryd
aEycDB5JvmKZv8HQE/A2Y48ke64dHS0VWXtygtp3Wh47tC4sjU4B6/vI8+KA5QLL
uOGcRWhAyZ+9fxP/cGShLQWxCbvll+nH+79ymvNA3Ejij0k5ZBVgrJa4XjqKafkp
bdg5ZFI6wmaOFMaHmR6zElOLZQwh1raa+EeccxBc6N1Ha/xsS7YyFqdBVi6uQl75
h41b4SBkwdwx+SNbXQpTLk+hodL4G2CZr8VCyMo6sHA9Ho0/frV7TAdLoJYNtRgt
3XBVH+bLCTsYC0UFnjNX3XMAIGnibLGQ7sz/Cuoz2XaCDW9QeQZ0BTWWy1zUGb7w
X9FH5h1KDcQRcd9A89s1kH6oLsHeHWBh8Qs5OxyQzygZtxks7uxDovC3rEaVA2Xd
fkEtIqOiTBG1d8zmurPhrXWsz3+y3DpHMIVoq4O3OSax3UQwPL5etQo+JCjjnla/
23d1Hsq2u2U8/L0gk3hlfda4vM6hc4pkaTIRErCXb4tIYD6p1dVYWGf0yn7ny0+S
tgfpu7Ajr0OcRkz8v7DMZX0wUOfPjF1wa7XPJT98ZQoXIgop+T0JhoP791M1es6b
+Efpxzh6N4xwLXyBc5NMjOtrysFKdh5YPE5LB50VH8rviVduYoeqzg6KmzjK4COw
v513DJ+KIUqG5idcMtYSzMm9S9TG0WU60ZXQjTTAje21JMGq6bAZpxEdIr6+E3Bo
/vgrnQ7JoOiktUFyn7EOg1Sn7qyzPs0hJ/MQ+8pzzosShYBvXGxD4TUD7otWyq/I
30qDffOUm0WuCHEWsju6XBzh7hIFWdwum5bK4ns8ksyasqCOqROcdm9p66Y64h0R
0DRzLPoS9mGO+wjRD04jbG4yljoZThioH7jrUBHKRdsqueUEZqYuzDjrjauXD6Id
abkDUiTc9eEmHRIDB12lTGPAAXJlU4Nhlk1U9MFWvjbgtHLX/L0miklC/8MzbDqZ
STH4N8tt3Q5qcBQjmNxjbHKlhfDaWD4azoD+RJ0yw8X/pfZ+/MO/eeXtjhOG/6ye
DWikLV//qaJB1kz7+x5cRbjCZ3jKI3BjYzDMQTQd72HSPJD9ztxqdijJMTUFLgXK
GHNzpIVBn7jKsbBetcRWRpnz+goA/VeeOSSanrfTMdtlxtyQe+396ua4vsguQf9f
y1PjBE7modXNg8C0ZygXBEl90I6PRFq5uFOT7tin9HbiWR8OH7VmdsfLn13UoGu3
0T/rz73eUqb4v2VNSvvIPxy5rKvib1zOswe6lAAWFJXu0kN7NEHTRdTjXmypLIn6
xFOraLiP72YlZJICbn/u6K9G1Vq+B0QtEyTaZjDqUFSyl/17hmzespGI6c84UIJS
AChVME/CWOUYNd0MA3G8Ku6C9HiVRL4bg2675oRl1mJOxcbK98w39u/9ykyeRs9V
9YoKahBbvIZ3ybD+fBn0+joo0HpchLbClsqTuMB82RL7moVpjbGiDrFg8pn/42G2
mgc3XQmcawfF5ejdF+sHMNddilx4HumqdeXTm1spl+aVp+Jx1mNrDUgu7tfsU6yB
gGGGn8YVRvCQKGexfzJN7b8vGLKnrW1PoaUYdoOSDAvV/AeYgfwjf27uhymHnNVq
AAIA/32qHJQQiJ9GRA9K7n8K4WBks2Aym5jF1NFQe5dybuRhNXqoaR10/rf7nifV
/yIqtYqMCuKI71+1VD++uQ86A8h8IRCyIn8sg/DmL2cNxp+pTovcJYTiY6rVf1eb
RHT/b2pQetD26CO9pUhoSfuSlPzOxlHLdoA87r/b9uP8o40uC5uwjSM8gWEuvZL4
l5OYEJDOYDPGvvUWasoall5nOL0LknivCocVl4PZeBYF75trF4dc0vDticUsV7q5
zulNf1+mGCKUaM+YQbLRYODbgLSBcBRGg23ks6ihuZaIIYu/p9NjjjAJIiJ7gq+r
pllLv6qqxKZ+Bxb9j5xO0njHO06jJmY0X8ufRbn2UC3UPx75Q/YJl+8Qh2y36l4t
oOiHsPqga5VJTsJemOgvvxL+1w/qanwduOILDDoY2MchWOPVu1JAOa0t26xfnmt6
jaGGqsBW8AqeV4L2Hm9PXOpFTx0J28up79Qa1xwYbHZl98Ucl6uIzFtM6RphL2Td
npmJ92K7VGMKcnf5ARRrRpq2cu0AowCYoE3UonAstYDOQH/UqoZOXAf0TK1ZIEAh
9KMrpcLQSoqJsGeV9IRbkjCIIwvdpBarB/DDM3Md+SsK6IKLCB4Cgn0krOKXVQ3Z
SctyuRtYId3XHTPlqh4VW/uXdntkXC7K38WYFIDKI1oQ2bVofzEMdWLQGcK7LmjH
Hfa6RRRaS6of+RIXAQyG02QPalmYH3u2m1wsmC0gfuIFRbVnP+g8VUrarjzbe0BB
uOxZ94q56+y3Pja21t2ZBHtflu3GdV16DSU/578PJ/NAD92qVkc1ICzt0CJ9G7WS
BYSZnofxgkimpcxhAhtPvFYecozUVJ9AvupJ3wZl+T+bi5aJEV+K4QpdexIhBnim
XqKHyiMFCuq/ux6ezo7C1YKHF4AgWl2x60enuXv2Fvz8Nt5Z4pwz6G225340iveO
tewaa56b7aWGjaspRSDY0ropcwQHTXHMAmVOJIKTKBzInCYyOnKr+OsHRcbt5uEN
Fv0XZBz6CJZczI/z6sEnXKdvuhSfZYE2LD/OS2U83sKgE2QQ0fqLVmh9PsXPAg2z
eqmpA4aTatEIvjzN4odYTF8vHnf89ovo0cDay2OUn++o5Y5SnrENXrdJ3DIymBRb
ehDP9jYFDw9CY9G7i7nqBbeZyLfuiCvHDl5fgNKHptTK7LqB/QpgWs0o5clHOT1S
WHcv08fn70jcS4wodEUhFSfWP16XVgyTORIxhF5fW7+w9ktCcgmCWljAbqmtf/M9
qeCJ/G5daTmzBNfNAGlwb8QKlTQDuM52hU+8BF82nrBsW+Tt6bhsmBAHdV4Fm0Vv
V4ZwrqBoQeawpfIvRaSaJrJUU5C1MyPo4GsxIwJ6xLbHXfNvp9HXHykKgcbX+jaP
6s07iQULVP1rDUn28SiwI+u3ocRRTAckOLinkc7dbYNKBufdDddv29A+fo6xNcoi
RsesOZGJ3JbGQTqd7MnQr94fLZBkJIkKCRYypVp57UEC/Q+wb5CfJfu0qigElm8R
TFSHSDXw5Muyar4nsEALMStTBRYQhmU2qhD7RsW0VlzOsPw3NzRxDWGznSy4eJCn
bsPeR8Z9zspB9hFDKIETtr5ZwMREUhHW2yvOnX16mrzNmtsW0X2tCOoqrfqWZEF+
VawEUy6derxMNyQ4NUmu2aCk9J81egB+VRy9q5IMHluOzA+RYH2NvJXxIeI1KWF+
tqxNp+BYgr1DWSCeECzWQH/MgsdHv4ojUKGiH5vF3nTUY32gYViwAiBHOEIDDV69
2EbJU59LAAKtFwyyGOj9N9hcnMt1wSfIiQgdWEj3IPN2ScD18v5yJhRw8LPPU3hz
v8MkoJJyCFd6XEeeVWwdFFFVF25ioJG5QPHBwCFzUEt1VuHpUkkBPaVW9V9CSEnD
5K4mMLGw7NwVgKj6TA6/6+NnSlTnLmPNXoVqM/BWhtYqTQFsrV8X6X4mL+sGdtMJ
Q+MiymTUMy7eTyM5XjJ8niYuH3DjujW7eITUnkQ/HMvHQ4tyySd6/poNlYlmQ/tO
Cb9URZ46qtLYQ6WtwIPkzjgHgPABbfKucB8pKnG/qlWvT1L0Hdp7TMPXL6DLFH5k
6hn3NoNa+lF5snjMe8tSJfyCNi6ZrEfW4cyMSgVygMKpfgwnS+vAb8uQ38K8nLED
dFgmMBZnSNg/GW+7trnMvh3K+hX5TWQFIk+2mWJxBKDDhW0c0UR8B/RNyTvJN84R
NhgJUmIfjcvrw76b54HHxXlGnUF/SemqiWP/+st1XcH8ITKYERJiSk7rncEIIeoj
a63FU6xTD3zf5TM/ZhZfhXD+njQyKo7pJ8ZnMNnFidOQh4fdrVfoJxyTNMSmOkBh
RbZm2Pb+LpXZso7P9pGxWiZO207m9CN+4ODcq7daS8s13K3tZVY5fwzWdzZjCUfU
NJMGFjwrjonj6g8z4CAUg4TLJJLCNpccBz8RXCHmTHdeI9QLk+edbZmr7LYVM4cy
mOhKFv5D75W+PWVR0ndx1BQiWuKr3Tdrj7dRT+CoV2RTDkn1/ZB4xa1rRcMJUd5Z
/IHQzQqCJU9PZF4bEDBpbgXIksqgcxEMRUddQIU6kBfgOuRTVqFmoNBEvPUl6uNg
Imikw7/P0GghJ9wpFI9ql/M2IVXhC6XNAF42pQw0oxHihKkpckDiJ1E6uxJId6sT
rkecqeAOGqHvHuDGX+/KuI4yRFlmPacCo/Ww00aUOn1vFdoSLOBWMvWh7VDmDJa8
PCyaRAHyixAI7Gek0ZDlTynR0IHOYbOeCSfmPL6HRq82W1L6zco7sUwzncmnuLOV
d7SNRRN0Ciuivf51/aIweJ3YUEvi89bbHWYHGLOuA731bBaAlvEfvCaLTBCMbhkx
FqsVcfs809pLcm3VvvN99edaQWiUoNqMKT9+y8x9H5Ba8izL0e89TI37zQ+0oQhu
WvbjVhi9Mt3i//U2Wfe/5SXozrkUbgaq2iQ2YLo9Wb72nOhIeI8IwGo0DSL/GGNW
EM/Nmy+BBC8OxPDcqlf+zPPurM+LjrBpUM5F9EvbHEAT+jmQVHkiqPcB+UydwtTC
JbE0ydk+LP8JxbdyS2MESByMk/xGxxOqKmctK9Rr6LxMb9j3AU5K5K0hS/yxhXR1
e6PhdaylUUYIFmLAAkHIG8p55XZVj1Tq/rz0EYEubNdqt72cp2BZl4qXr4r/FDkx
4uBteqsOYec0ZGmgn63/47AKYWTZvoYR4ccnnH/0i++KDcnW9LHyXd+K6lXVeZhJ
4T26aJtUKdMjB7LRK793V4ct41DAEA4Gmf8tPI8jQBOMsgu49n8IDWZ5RzQB2EqT
oqCuL1wOoSuw5zU52iZg9IV0INp0kaatHzBZ9H1Hf9yHxLJso1Elqmk6k0Nw22iS
OVpB4zzX6OprMRPfDPEOBFn2VJHpNc7kHxiDsHTUWNavygwfV0mOfdDWH+iBgxF4
yj4FniHLJ6vyjFvZS4SJGYzGmOIwjNPqvPH9LcSGvAs1HLE/CO1RZ36RllfEe6hS
2WPPgr3TFvES6cyr4kLSMiCpEA+mND+2FDWSc2AfFjIBwGXaQbc0oB8RsUvIR5lu
4lke1EVoBUM/b0Ib9Kj7O5DFwFvRpDt1815PXYXN+FQ9Kt9ZGC6wV6tfqxRf1+R/
ZQYy2JO0O0n9YYh2n9Estf62r8iIoTD1+m1c7B07dHSaTK6/30ujEKIHOtephqF4
ByHOnWmnDNxRMR3WzzEEewY5If2ZPIzAx6klm6x8JYNqSpCX6vCDQj3qdC6HKJmI
6fy3Bp1Ub+Cuz8PhrcZeTNGrGVIhJaFriSnpNntZHqeHq7b5ItZ8OACJ9x8xzLkE
VaEPs4mnEcTCGPjuBJmiXHn6x85RWUir6uhGdgKgGKblQf/mqyOhzntYr7VSCPRn
SkIJPBBvLL2nVJ13r79mJdACTrlxvZqO/Ss+sU2q517MDG7T9TUv5rSfJtmVVmEA
Eqvnj2kZ+9ZRlVUYscsBat3A2Hi/+pq0vbPWAZvqNk6Rm7ga4Ly+55wZd6vRg3IU
/4BU9tbG6XgeBssnV/pBI7yDDN8hwqGOeIgmVL0h1NafugdZY+M5GhQQx0gYKuN2
OK9bagLYwAREcNmcktvK6pdCTpnPxrKT0ncjmQ/EVY53fWQnEsm17tIuinDW5o+K
0VfFJBGPDdvth/iOE6xFMwk/dBvABoZeb7eWAuCGkSLMIaB2fChlSyWqefyhreG0
Qnqn4gVeSO+k90elwMgHK8By2R8QmOH6aFNXkYuDghBcSpeOym8XFoTv0Q7pigb3
LyN5sY5r64pRwncd/LYJu5FGJHo/MHf9O+3usYc+ah5YLSjHSVWnEFPXiuSmdEDS
dEjoPPTQ108CgqehdzXT3HkxulqOycOLwbuhkSRgc0aA3eHoOTxIwVWtBbAdbT0V
75JJLcZGBKIO2/4eQY08ny0Hufoo0yg4RxMO5BY3vOUUDGmYTo7Jym+WPRIk/H8H
gd4bYPqIfT4sjdh2b8+WhR9RdQ65EMzqP4YJt7TZGC8PCWT7n+e2MPseBwGzUo9h
bMwsQR0Twjrihv1ushsSngoeJch+soM/uEhdNzHdkZfzh1UzWP5jaxjlKajHXHOD
QIdjZE1O/OTQ2ZxZcMw/jGy7a0fZbnZJkenIIeYabMwyuRZMirKNpXTI8MJ9Oqed
Xq3TimBGA5lF6ZyQOjE1+lzdPtcYqD5DUIrbVV+U4OO8dvfmXfIaIxZtn9pj0QZo
34frJmPd1ICQ+MGfG01kqON5gkGGhxG21/XaA+VZoYftvvwnP4TPACgJu9NIxljb
Yrn4Y9s6XZSMv8cpagnzObG83prnLau5OChV970nyBIknAT75NDap042qKOyR1rP
gV85fh4RuGCzz7m19YfzGRcjwTXyrYy0DpCjND6IM51SgCIKnn+OJQpO/UXHwiDI
2pXBvoKKK/IQBQdSL4B240xdgGstXWD2ccXstzM+dp8ISDyHPkk+mRq8xOFnXkk6
7i0vHm02B4vx4QZe5vXfciapNgzKh2mr9R6I8seQD5gvAjtRxvI34gVqx5U0H6O4
NgcT3stbTofGFWO6sF1KKDPLdxhkjetBjoxx+pIj+TPPCCWoGIdU7GVsqrGA5Qxn
fQGI1592WzcmXEKVIUH+cWD1XI609gXEXUVZdP7NdDKNDHOG6WkBn/LhjLw9CC3H
VypehfA8/LuARZGiXMnNnj/TpxmY1U4uFacj3JEDd9ZcGRNHNh/X4tTZ8Kt7HPMS
wAH6+33wzRLUyZlmMejF9ikuP7k+KvIeL5kcx0mMiPd5Y66nrZImlnR3+xL1YRVC
xu1bGJEttt+bjkplFYF732IUYVCPGLFPfkwahd/H/84HrJFiFhOoFxmAQUa1GaNA
ojbTSVcrzrGaBpSwmDQeHTlfm0liWha7AN4OVUjkVgtG8/Hn5HLGLLgwWObs371a
cnVoOPokZ/DGZG1VKzisxj68dInv6A4QonnJamqtQizL4ORNYxadfj/9s/2NvIGM
vlXZ7MAGCFQ0II/KDZ/Z2g6vysmqukTnkNSsORh9l8sMByWRa57zxzNRDnSA2Xu1
r2/nDoK1yRjPZFAHxeeUKHjLEZw0RYGTi93krFlxbgOYG38clmqfGCdJ2AUyD5mA
E61O563IU6JUj1g/P+Dv/KTFQFX0cWx1cSD5Ui1UqRhkhsFRZMWwILlJIqg7Rbrn
zGDdx6ihJt5MWUPLtfu8HOUad+3SjvkhyvaSkkc7IVCs7dZVoqA4k/yP0mJ4TU+L
qRTcqfbeDeBMcEz2AOUiePqGkCo0+AeI/8Fo/2fEjEIQhSv0885ySzGDd4cWCPIV
Vv4zE6XrBNFUijEkWUh8L86zdGcVuFNZzB/Q72HxHICzuLgYlkwA3XQVVoB4mG0V
kU08kyVxD8Xt41vTbaFgh6DVq38rJUPRGHHI/nJFBJcaofssNfcKAW5xzQTET7sf
Gw7V5JjpaaVT4guH/pVL4qNq+qbCcpfGeuoDrnxEGOkq1rwzqpq5Z41rCqLJtBw6
nAOOc5Aop6WP+UqVTPr20IqM/V5uBYAJSPfuubI0PkbdYJTbklNwRNydIRh7VQoj
z3lwgtqYjJmc5cKjnlHbUC5DM9eMvudzyckJK9WFUeiHIGSDqU6rJrepyjXdP82C
ppMRY/DzG1AiF/QjbD5InVDUYzBGZrZMOYaRTvhg1lQrP5xKTm/pWPkDmY19nNdU
LxwA3GNVGM6oYzTZbQmsV5sOD67dSvvD9i8qe9gYAIch5r6nqdbFnphR6toslsDs
orMNj8nV4R2xs9GFMGjQ7Eq2IR6jMXCM4I0U4I9jLxEaft0QLpyl6lq8FQQRbt8O
e1Y8kFdTsS2jjYA5pS3jRl8Xg9ORdYRN69QgNZWFPOOaLCoHX3OTChjDr6GmBb4l
toq6WIykhfR/1nVM1yGJN/zRvZEbDp46Zj5HuHA0uNczXCMJ1OyVXRIXYu28LlhX
uTfoLutB4JzYLfWQpafOZOdqc8CyshWWp4LoCDKHXnQbHTLQPBbJpwPJTYDxoEdl
NHq2Gd4hiSCGXMoLD78W5K1hqMH9CiNBE+PicW29f0p1RiA2qjc7uUkJLZuQkMI0
CcSxiLiyitu7Sh/fQv4ukm2zb3igrKhl/sbAGJsL//XYYgil36qFl4bUJsJFoCKu
4gUCHZRwWFpodHfmtTW81hKmIR/dqv8O34QTkOKs07K3I/8BRvgbKjTgUNkQOIxW
OnhlK33YctKUXgRqchwOF4FRl5tg7dQyO2pjEpmWhxg2z3Il7D1RHsQ7n3jIAO4x
emLDgAS6LA+0+lExL0Q91tV9DzLCBT4GWEYwaXrwiiCHgXiX9fAUr9g8durBXO3j
yDlezPrnb4dnwUAVAUpd14wSi6eYYTATmLBn732ebvRnIaop8cp2o/iti63zxZfW
62mpilrNFAs33BS+N0rEp5eb894s/3NeVG3oGY3FupFsxw6osvQsni4Anf3W9WaU
zboT97ZFDazp5+xETLZ4iXjJDzgGoUnTTPOfKKLQiTtKsVE1gpdE2kkXKBRqzgxS
PYKwvQu/hzbAF6tVtZ7sG0fz8TqDESXjSx1gwfs8rx8btl3MRUP1IDND0y9kuU9w
2zsB7dHoXuApTwjSon3fAFvgSQT66KD4ZMPRq8VZdv5xxjkdeOL+hp6feCu2JSTj
r7jcIzpcOpAMPQFEH6Px8K38qbEiAOvzZ/WoRS9rENQ8rcRJ7XA9E4yE99QseyhG
rJJl1FF1TSf/NvW9vMAyAlmNg+g/dnCTVbPla2yFRWksaq8q0/hyFP1ohl37foLe
MkoTtJWVlJb8OAt7CtEuGdMJhvnKGueorPuWaC7TuvL9OHo4MN7Jw/98K+ovU+8E
Aozg2J4B5O7y4jJLkZWpf5uRmJKvyxF9g8U7d7xQjYa5dSXgo/cFByTpprFKbpub
30nUmf3jvseF7obil8OxWyuvQGZTwQrGKGd79HYCJJws5Yl9ptimD1lCo3TWSzbZ
Ni01ZWvYjUlolRQLu7znlHlK3UP4tIoO9GlmLj3qs4EJM1Xl2M37kctmP+qDVgVo
ApD0lU1Kb+94Vu8Xwnm8W0kzZdywSzAJQgLswbopQpctgm6lF5xTQhXvBK80wP9f
cwQvpEmJz8ahr1Sz1tlPoKuefDBm5Zd/Ym5kqwM1XeeN+igUVYgUaLH7JQakAe4i
tXAx5ETZdBK5dNNVVilP8ifEFOSXkwQN9pPQfHHOg7x5mx/1NUWzSh6tcT8yqFOU
I2PU26oenBDF0XktU8W2AcazIfn3pK8xirLPZQBGD+OZnOxQE990f8K5FZgSR20T
g3Sz+K1H0P3tVkECjoRrAE3LQV9/xfROcU7mmP830eY30pKsWmn3hVxT28igrNaE
N/L4EG8HpyIGbrmiLoh2fRptJAP6xydgWfyfXGYMfdW25oBFatjUSysw0y3MfJnh
/0x77OXEj4CcSZ7g6SxzbmOT1Q8CVabOFgSJ6y8aqtWLxdrk/YrOibuSQ2KRVLNc
fUw31VPR8Gq7PB+LEkIH/XEZOt3P/O8+Ri11pY0PM3keJQuFLxVQQd6i+krI6BF+
40/GNrcmNXBBsLUOAot17Zu4uPqvnRA2+mj8aKJJBrqlJ/1waVIvHIR+DmVpAKtT
io+TRRLKnc2jRpjBiTDGBTa4auEfEvTI/AScSivgTfM3TIz3WIU5QiLObvzTJ7Ux
LLl8LZOhEHHxRfWplj/omo4t3mrgXHpvDxMA4DXLvnB8wqhbMHVrYrO0HK+Q6wPw
9lLSwTI2htknuiqwn+HLUop9IRz1Xrq9c4tm/D/prSu0zu0FYX2iDoJojyFUbk5V
Pxkcqs9wK1U8ILsGYeq+p14J07cZVMoRGt6/iZGc2qBLZthCduealPTall5+UnDW
4Ma6qyVIifVJFrVRZEjz7MF0rxGuZt/m85eFY5+27bjQOwSHARex+YP5cKGWG07W
P1Mis5PqqNRQUhNhy2Wz3U2TRKVc5ny4Z+Na5y3WJ1YAecTPqET5TsA97i/Lq216
/YQZ7WyUgfKvzcvYr5qZkh2Vxts5lyOulEOFgVe9ZuyidbwqjaQOtiZxrTSEztD5
gOS5E4PoUm42AtbbyQB9wUZUqLg+Xwqnmu1bsOJnIDWcE6S7M9EzfapbfX0D0qFc
QMC//AMCKSVBpr1s0zDn+TOYA4dXyRoG2C6U9Y7RttFNxcA/jGnrWftnSgRz0np/
MIIQqKDRLqOl2uJOYLwmU9EBtOjdBhpnWUuL+rPB6jLA8i/jY7TFCCh+9C0CjwyY
zpvb1ZP6EmX2oZongLqIYqXlPZ+Fp7c1GPUhYEJBS42SH316hmh+axl8Z1LMuKdo
W0iNTkDvgDj2VS/L+zaMTV6HE+udifPXV6CBHBbfJ5uB8wt6xCLXv8pbPwTuuJHp
ttIAJ2TliHvY2iYpfycPRBDKKOOSSP9wJftUOhNGsi9T89MDHpjLVeiuA2zA7etq
jAHVPDspzN69e39Y+jxQRHJR1XfhreaLUgWUoF8gIqHhvQB21sa0bA3VVJEJIXPp
fItNCRWmEOpq+gqLhJrsxGrEr5vfDbra/G8OV2xM6GnGeHeXKzYY2V3CSLVwjlf7
/nB7Q2/q0bK/J/UhwS8sBU4+RUQbqwEP/aTCogq3m7Fxm7IbSgMATeNltxQhL1Va
huwFHcQsbZ7k8hD4eIr0zThFpblGW9m3C/baF6E9Ue+hPBjuiCo6HX24Wrq1f49u
53jgYvDxQykYKrQBWvuFp62IMZD0i8C7/SY3Tt1wO71357w3MDQzhzLSx+h0P0mB
Q95e1Dpio0V4hs7lpM56oZsRAXp1P2jDKPE0cmtNdfB9Yt0YMO7oXBFYImNF23Af
C/wJiLU4QmahbTg+1c7DapZLJMPf3X/dfNPG/t3OLV8rzN6oX4Ha3e7wYlL+4iJU
YKNLSCHXgNXL92iKNT1G1+vC+k7DCVXHKG9DAVyIyKQEV1HFLOR/LdW02badN6iz
vsBLE6jUoiD32H8tMFIQwbxyDUwiNAWd8jKVGbQiu1JlQwhqYlcucGZAj3GP1Nyq
u83b6oQoQX3YjHwbhWw2IFhRT6IwDsPmFMBl7H9f8aY73hqezmftbfJ9nRZ8NJ4X
/wqApdr7rlnvGxg3pq28pe4QpvMN9hXcYNg2wWgcyHux0ur3J/KhcyT8omlIYfLj
zj4JOIbZ0CZc3OqKo2IzIfIJj+cmKAisrzeb8UQP/lUy0lvQqReQMmJVAo4rqSgB
Kd6si8QrbRSUtPh7UniPPE0CJ2RgnS38vU1hfh/pgygf1T2cpIzUpMAFj/cySD1/
bmJUPC08Ayrl8qqZ43ccY2EtQOUHArUZfxER5kjko2bm1nngyKTLzB5ohxbGstNz
HgU78QN6e++s5YM33Sm2OGAVfl4Gu8xaasYhvwgXHXn9zJDrmy4UK9qNrItWlpPV
ftebtOhTXaXruaoW7WYblV6xS7LancklPaTT0ydMl6w/I0vBRJLb5Aoxou+0kTHr
wDOfgFkfb8tHkzwYdcEUvC+JzthV98aV+LwBwQGASIcJVtAP7NeNd5FA/iskS6Wo
UQ77JL27RDZmn92ZA3AG7UKLQqKPs0j553gq8Q0CF1KYT+qtKlI/tFYwzkHcAJxq
/Tf0h34a/OXaR/UmzuxUJ3d/pkI5HDJX90Qw3rxy52nBht30S/ibPL5nAESzOryn
AvFGPOuwdVpr+zqZdN1mh6gizjXHY0IU+bOwRkcX3490MzIytlFm8mStlvV9GTe5
dC8viBRSchRi+SwD+Tl5yAZx0b0H9EArOokK1sE4/cVFnAALzkjxxZZ4yMT/cJ1I
hvFTA4OLSqU+wCt9rnIZ/zwS52Opc18IG1iYVXjHv3qtdyJ17zYwpoz4782IyIAk
quWmVUmkStICes9c5rucN28ymRhW1zlI7cvSBuzinD0jJnKeBtEi8Z2y/aBCGUYx
cv390I8C3IF0kVVrN1ylCW2PT+EtwhJdfq25aDp0KzNGCogZ9Ydu6WrPH6ckW2yZ
k4AqJPcHcStIaUUojMvYOVXxV0g7w/gDY0veZ5c+t/6uo5EVAOCarTNjCLDdw4sw
ynfTvUF8aEMerdfiqqHcPcbOMqkKac9NFK60jEHe5w1tyRIBDTf4/oTpIvSOTCH6
5zxMwetpolQfODiuv3NK18J6JQqTeaFX9s3C2P6Bg85pEQcgmcQLqGF2OT+cvgG3
luoE2GspSgRimwGvBD3wzlhuk7UAGreaut2O1QYhJJ9PysCWxrBpEqfAsAw8faG9
o6A13OQmdGP+pDhNUo+KV2CvEAYp6xjtBzU3AMTxaFP9iq5qvgR0a5bL+CnToz+r
3xPQT7cHxIluz0jAY+8IVSw85ZCnLqu6u2fLdnfR+9vm2t2wVbU2Nr6/cVBQuujd
Ln8lSqYFic0RfMrX3XqDNx1r8MV+UkUnTP8aTJrN3Tsaa4YFuK/qjEe0JJvyRRuC
i6IneDwevFmIga0e7JTWQLAFiaoqVxKLdTvp0pfuKF2C4Ytp7D3gQ+ycvA8APrn+
IYm9pP4RcTozR6GajAkTFe+ujID4ApaIp5w5dbVaPgIECZT6EipOlnrjYSfucPWF
cbHPTR/Im6vA+MSfNC7Y3E8SdxRkZdWZvkSuj0qwBo6bWgPaHHzr3k6sC4B+wd/2
yT61nHtzdnP4omY1GFMcwPkRhJdyOt8Z/E0ekUTy/1B4Q2wHMUba4784zXoDFJ+i
N4DZ7dv6aBQrQuaN5tQtWsOI/y13lpv8tV6Ok2Oi1IMtQKcDrrDQsCJD+/9PWnFd
aK8KAhP17+OPbsAToXEzwzyjFffLMsrhamBLIJoajITV2gZcmruIB/HugfSJZhZL
3zGwa0LIQZI1RZwNmj4R1tiW5mP7Y1kEnlvItHxrwRqOPIqWq1zip9S0mAoxTkEi
pcjAMMHVpzChQS7ECwdmuU7paICHusyA+cdjeH4N4Ek9c90ipb64xEbCyzkjZlwR
OHCElIzFqxHvPoTnnZVmxCS4cqLREiPwuddI2Ygc1KuXg0NRNTC5Prr+G7gAtUx3
qAl66mf21EqV1naFylB0EcbdPBbTidrseg33jUk+XDBEjOcMt03R+PK4ZOjEmq6e
9oK+qccUoSg6WJcsh1JSii6+lphw1TL2W0FIfYRDX75JCstd+O0O/EFBEADpr4aF
g2QRKr1uTtlXyWbuo4oqEcZQ3VnvvSPMIlJIZcaycfus7/40+G2yCMX42zFCAiEh
ReWQIxs7S7o6nwZInNyZFq0ayufoaEaV5ZJsEU5Y+9m5PvaFLewa8bNQMCupyIbp
wisOnai/ecRiyacw/rB/Kn4oA1VKSi7SdHuFHCtIkrfDhCdYXHUZDZBSEmcpjE1K
VY4FiAlZnAYzJES9gl1E0oYeXbQFBc1ddoZ5qc5cuXjR570gth+tMIxf/L6nPxAx
EOHSd3cYBOhaczrQhYUtcDr0EJkfcMa1TapNZLNaKRcwuO0wnV0M2M0dhCumLiI1
ejLokzUlgCOZHpYP2BKxx0/qChqUgP89KjMYiltbEIzE2xJ2cVxIa1cdbUzsHkdF
sCrYNiZR59QfJiLaQZyKMcp9PJPgSZa4ja7CyZdOvo9TIWq6DTlBjlAup1jFLE0A
f9y9Iz+RXWleFPsiGz+SpW+2gO3se6fa/LfAaz60CvV9uSkik0BcHdSBKPsAJWjF
5YhncfFmGKP/562hD7DCEp/hhTWqeWlpKJnK5QS/OAlmGk/Ujj4MhIvP0F69aUV2
oa50Lrr0M6WwU6vCPRzRCIG7uUD1vZMHJyRn5pD97OFdeZDJbSHi+i1+IMVsrapk
P0+kenNHq+Yfds7Biwul5pmrA2nmBggTEdUw01ChMzVXWcSEd9PvWshxYeQhK+kE
quZx+jFiE0c87DnyTZ6rCNVI4XO2mPMugunD4uBHA5088qxdD/yw6uuGUJZueAJp
oZCn7eFUajixhNBDASTbfaXJk5W8Yxh5FNQcBSJTD47du6JHMpY6YI3IhuZZydN6
BYdtCMOGxQ3YF0y+Iii7/QgZsDgDrl5iocWmLHJiRvlUl2P422C5KdCXxKnHw80o
Z0lK91WYGlG7I/NohFoxKlg/cuAa9vNL4SQPR23ZNQR8Pp8ITtb8cHPB19LGCWPg
b6D1q2/tHcVF2v2ir6x8J05oCCs4vaJs2rnm6loB1QB58+S3SgF9atf6qOH3ECDP
fdVV6WTwW5GUNRKF53DulAxuXjwACNulYLhVCRKsh5DOlYKF3CHDNPmCv10c6DH1
tgXHXz3fFcDFpzKLOX4INiQKUULKdMOuz8Tb7mH21CeB/lOAD+Sxb6BNSaO/tjbP
vJhTr18A1O5yKZzHMZdkJmsmEp58BrzVEWukJOvfbAhvE+Lp+wPa/j2nOsU5lf+D
NHo+9juFozAnwxrxqdhZl2NOVXj8/k8lbLDZ71Iz4+RCrXlzRq4gz2pakQG6lx+V
VYk+4p7avUARbThvFDNaPw12C3Js3VRR0/BuAUKTkoHDPqObw9PNLFztPyprZqhV
NOagPON4oWIDi6pWBvh5yD8yrNOrdX80ib2n/UVw2kWOJeyT8B07YY6LSnWDvg2v
1krElJrnEzOJyhN91As5G1Uqa3Wan4PHRohQdTNKpDbPI013nc4lBTAE+LFXdLKF
Gcwjx0ucVrysUWM1Ve986P7dFKkLMNjNvsL22pgyqa9SsJcMZLLTz9jbZDvv3MVn
hcVOGApQVqDZfkWg+d1xX9I+3+Mtp0nDTGGVdzun5ZKwFLbzqcqKBHwicY5sSoJx
t5RJkCkI7sLTa1yALXTDNkuHdaFXN/iUXqhxEwVk7vFvA2QX8MsefGeZdp19n2Bb
uhlVjhzBJ3z01N974B9QVTDRlejsfljfW/oikYYb4bgAruwBh9tG3q8KgOUnFIV3
uG89L9sYillBnc27FRzELbsmwAmA+CXZRD754qZnWCKINWXZcrPv6ZWPnYB1YZOL
msDPjEi9Lrhh3A4nvYOj7e1JQDaOT5JY/FtzJBcbl7Pwb9Fu2M/qooQzsLACSdUW
TSznpRWvLjTpun5xcSbpiv2YsbL7dHOeNOE8Dj8p9hPESRqJeYhbUpaDw9HOERo7
f2wfNSW+Xq8vlvssY0ETf5/j0ecbzFDXrxNwY0AnS1/jdTTJFWpAsyuyQiTE6cva
f35VdeTP7BzI3rSTpfrrBig6umZWEQ/SOX9UTdEazaMoV8bzUe2lf57YzK5VeOC7
FpzuhpnobLi1Ltf9j4rr2+LpITtQ1ERoYjDNFIdzCsSicAV6tZweOqv9nLmItU40
jeO4Rdr9cjBAXYqsSp6exf6tQHNjm6otm7FeyrLz6v5Jxpu0IlUwznLheuu7xUDY
yCKsrlsJm+4q1KtJIon8+LA6kHQZRcVwjLKcqndg8YO1C+oC86tbTg+Pi1z3YNcP
SIeYOhQ5gI02gDcal5ycQfB0FvxgQB+YO3/KinBhVHnDMJ+9Jfh2ndG/qs9pL/fx
fp/uAfJNZm0l/dhTN0fH5/Ca6/GRuGN4yw1jLJw0o0EuESHkswJaC6gTaF6LjhVn
YtMDDiSj4p/IAcIs/RSZjSLguwi+zsit5GuPQuXTG+kJO89EdVx+xGsqq12vhpTS
w9wTctq2Bg/gt5MXh0P16tkrKNChpl2u4mJrRyKpr61AXLtZpBqLkDvQ6R7EIhLG
Jv9cY2S2VVWLhV9NeGKRKPiC8s3bhfX6+g42X7xH+wi1zNn2DgZcpkDfLVQveiqB
xUh8Z9o1eaeZbuhAsmwfxQabdKOx2SGTKAWyem3qichThP07/3z3VKLkbcqIyYeT
VQ8XlobPIMI+S7Fah48YfKF2/iJEmLGHBEk2zmvKXBAbsDJ9WNnu/Fhw6kiurQ4s
pVs1DYSlSHeTBQV+Db9nxlnGZUmcpbVPBQJ7xjwqqIal3KWTN+K4wyyt6qxLhpHD
nI94U+IBLplugwMgpKTI4EU+Oh3rOhGF55kwszG7agNFZMc8qxYatBTch/K99pXZ
JGyai0dhCPzu7eO06gYpEEst0/6fam7kVBYnOBGZHe0JJRoB0iBm6KHqxQvFJlC9
8dOBeOTSOPaN75RR7+IW1mydBKFVFDptt1rsKv8q/qk+KgeC/R28O+n9Ptevyo2V
nZ1ShZ9Y5VpcZb9wHl1v63Q3nS4EXD5tdqf6ZYjfvgpILTknyk+cX8y/ZxnIYyoG
avVTcO1xOCb03fIxro7/E3lqP5iIUkkaC3zaALr0AckcdePWO1mGRzz87y/92uex
8JDNwNbjaIx5jCYr9WM9fb3c6QzCYmaE7uB9dD9ilqP3KvsnDzPijekMn8cd5qPY
0ozMhX+RMZ9VfcjfHzgee48UXkNrPB6Ve9YZkwwTqvvc9q8BXk1mzRQ3testfCx9
DHIkFVtmgOgbVW5CnWB0mQg03yUqlcg1cFtdFHA7gOfZ+VvBByKg4KTGY90m93mF
ed5nVvG3gPe2WHIuHpcP+LZqegaTInVXL1E1jfJbsTYAwplUpVNSqPyhFBKYNTmu
aNARa7LIvJs3cv6y5ft2L+xVglLJQxf+4BVMgHu4pXbGD1A6Tun9fxeuu6yoS+Tm
gCdJuyQTCyCD1Ei7KM5s6ueznejFB5Xpso7BA6+8Bl4zFUX3F1hQGSgzX2V2IY+N
V7C+wwXsphyQ2sXKRmJixr5dgefvJ0ZD2AhojKqHjcDYwpv2i9S3nDkCuEiLvJNR
2gev7xHvQvuGMIwCTmtdcruCovAGV+KcdHjTvjqE5F3jyMYy8iBU1A4NB3L2s/vb
iY5G7JW+8NaRF4b+GWLC+o/nhj4pN1OKl6oGcbqzYCjrphfMKZfs1An3OUV7ohFt
PEzF5zLGcYsm68Qs/DLjige9Z//+POSAfpUcKCmGBkl59d9xLeNaHG8E1e12g3EN
2tz19ZfBDtK6yPYS4o5EyirU0RSb3B24TDwR8G13fRvmEk4+yqUewMyTxFzxBda/
zCzG1+NDXaqXt/RLx+gYeMMYCBYAv4zB3pLUCVAMsJak+divJeFrr06LlEl4RcKg
vmFL994Jj8D9QW73X6r+dgbLySwBKej4/0Ae+UGg9DoKv7k1hMr1mzYwaSf7fDMG
oXg3gKc9WNp4vjM8rVZKcHpunZWXd6xqGnj+qBstIIqufdR5+j2GzQU2DHzweN4i
44nknbXenxmKgtkGNXNeZWmLwE/7mTfWe7+yhNF3beRdwyDgKbHpfatdpbjaseD/
riXgziJGPjkYdQ55u8tDc5cYZna8Xfz8NwH6wjiOvMZn8ZEANtMr9HHvmK3UOFda
P3eg0HMveFG+4j6+fRY4CxxiuoDIC3fuy93z1gSqAC69vwJ6VjTvbrWWhxc2h3SS
N3pQdCQJOnrI8z52Tg4kTIWy7nrDDrlDeC58XxwuNPwpFdZ37DZazykx+h5ABVFD
C/AJZatRa7fRCV7Zj+3rVP7kThyGt5tzeOcDpe3yxlbfb+mMbfYtKFEImPUIPnRG
Cu+3gCqTF165/FLhs6R3eaRz2MtMuq98rmClk9niBLW9R3CbeeazaMrZQZ2LgsTC
iagcOfVpqqXxdyu8dY+kddmShnDD/93tffVH0Pu71Q5IQLkhdMsyxgc173JElT6/
KlKv1NeO/HENYBi1QUWKk3/j8WlMZpW81hd03nd+J4gKPruo4vXSQoGf1u1LeRTm
MuwRvtmkQYNlBP/a95SGRb9GGTvc0WwytyuXFbWXlKcMDv5Qj2H4YZqugR07o2l6
sVLXNTkswQxkrT92bvtmYiQdL89gouZqtFXnFQzW0fJhKYRblx0psHPRuHb+F7Xm
JJuFfbZ3Bf7WQqHteS6b88kR7w5qnTZ+57E/xByAGJVJuQH5tjkz1Et/VNNiLKLr
F4xeUExbsDVQXicjdBexpcsnSMP6pb1caZ5yaftzk19vDMIa2rKGKACTPqdC9R0P
rGEULT5/erdqJoBUBcyMOOL8CdaPiNTBhA7YOy4roE3L3yeBzQdvOiFjSvpJ+rFq
38yfb4mcRsBCoO+yXJ+FiYMI59daLbiGnW0/sxsAjd5UmP3SdUjKn25T7yHEaNRh
5FDJleM104BZMdsWNR1GUnpHKdrqcQGqByhhhoJeq5EDhzAGdX8Sal+bYBjgGNql
suzxa+jZJXqM3gqX24ROhusiDrn8dST53u2t9VH6pAOtTY2yJom1nFXMn/Vsjdk4
7n9iADk2j9telnWCvOPFEXtQz8yYNe6ZoyinVXMPUYrv+kzLtFortEE/5uarJ20p
CiqigGZNY4Vsfv89UtO/5AxTnpZDO1/Kx2bYJBRNbvwpDxaPrWrb4mMeMV1WOsk8
Im7qk/wrzlhhd1KNF5z1JB7PSVEXE/D15nB52rw3LyXwIh+91enyJn5y+AFi11at
vtwdOa1U+conMp7EEztv+ekrz9hKAorVzsmQwazqPly33CxUL8XVZy+/vksVtCnk
EyeXBar5guHIFzTvczN5ENajTmVnfGh77t7/uvxMqu5z2i1AQggM5BXGIN/CEkDf
iVoyYrCNjAvMGZsFTM+wMYF9qpLIw5hPe7ajtIqBtbTj/BuOawfRyVbbuW/vsXSv
qyAc+eK7jhGePq3q8nUdttFAjdz+rX/l3FYE2wxKDKzkPGuVAL+SM9FezcK7W7ty
AxmOM8GRrnsgJ3t/y52mhT2wg3Q/W2TM4xS2/kUXSNQIxiHwYXHMvw1+DwtPepoo
hhnttpIwguwQVOQRv/ncbpjFaQhF+V43JdGNa+hiR7ol5NyMesDNi1noe8zNhpTu
xUMYUP0MTzM2sF3+NZUHTuFONrDEn0CMkUXOs90buDW2aMZ5K8T+d3QgG344L4Ol
+mtx0c1rgHSJgbCfIySLzkQ3SyNGZeA9DiitoKlEhR8ouewLpOL6ZNInhhF+THQB
Ly4pu3xv4JzcH1IrrtTsNqL4RiyjgqDPb9kmPHGddkb6yepx7vW71YSVfT8jAnBD
qIrKDa2WsX3MFiT9vO+iqAE0x7ck5dRlBc5K5CQiPLutbotRiOQ0CuNTgOv2G2re
2qDTom0k6B6FlZ0o/d6U0M7qXyfBCZahKksf8S0V0VXFUaNJfb33k4JM/cN67MVH
jneTMoRzm5+D6Xo2UG4uDZyKVszOizyyiobzykst7o+UTqDl6eW9E/yFiaaZokih
xOIZZLVdtSVm/89npWdiy3OVijsjgwhQek9jTRbruRRg7PQsOnnIPhNOgPWhFQs7
8arrBs1CKvscAi2Ns/f5+5rMJbzhe1jLu8tZi5PDKaBu37iFGoo+na5P+QaN4snl
zJCdyS8HrC9OoOLpVU/gx1iKTWDS2m/sN0mOFjzCBhOOn8UR5RnROnpgzPuyHdyt
xN+x3NPYbKmy3JFUrBwSiHePNaMN222Z36LQp71A0B9Ak6tSvSmg2WmqzJ+bXvxJ
n8UJGVt8NMrhaMZQvc9bx2ho7zYO+pgD/kOhBQqr8f4RhOy+rEQscRU0zOo/jI3B
NWoCdDF0Ed0VrPX1alDHd0VtkTdAt4vymsaTUFx3Mb/KCyzXbidvDjh5JO+VZ9XW
dzSpdbrunnuS9YHHqQ28qaIgq39WmXG2hIR0s6ysARtlCkBMzCZqhl+xPoeuXlgg
iT4JGdu5uF91839BBCzD7QGyIFNsWXCpm0rPmBxAgE6pz8kzGujq+kY1tUMDZ8Ue
omKrAvbEvp+xVDvPIsHZUg7Csov60DJs34zD6UmECF1dciI1zKpvBwmVPqAIjRk8
jOo6F6FP9O/2Jn1/JTl7zwENjUqtbmuaZioZDZf23URO/7VgoC1YQZPITL6zdltZ
S5OXFPBP8bCfwv1aSaS5VorzWwh2Rj0Dc7SCvMrd3Y3/YeU5vOCmCUdGMk2ewUNL
XgCA4wvMsbGFQi20wz5+XgXqgln+7d0BrpxUNIYjsnrGO1QrIWE4GLjhqujfCBPY
Vj9FM5NgJcRD6cJe74j5xzwuF2WKLY+nz3mNFi74NKbJvhvpKPXripxk8AOaFBm6
oV4Lh9LXYTy+/Zuq8XCF+RAfY7aTn9jnxokMoHKEGf1N9nKXl4AjI0LOWNZltWro
9+80HU/f3etj5MgJ7dTxaQ5w0y3W0LhlfcNMjwplkgyrlW9d3AzVsgUMyqflHcv/
9q4w7EUG3MqsgbxpFgfJYKBzANYdJtsqMygCgb+S5vVXS+KWXA6nlB6/85vT88Ao
QczB89Xy2m5T9pIX3V11Gnef9r+Mte+1ckpdiTdKXZBw9ITAr2tcgrg4LPMPJiuv
0QHZswkTNzsFVbXBlb4VJCvJV0S6DMVz1BAunArWLKTLhXhuC4CT2C3NQEeG9P4c
woKueEScOkSsgRHOsQwkgt4AMO1wsZfHAwHYg3hI34+dYAPWRcUopRAq30mXN7Ae
4c2/W0n65mmBvXkkx2Odu/ezhko/U4upzTdR58e1bwA4ZieelcQwPI7xl4Q0KigP
bAlT7IAeZfJo46rgeegZsY0oaUUMMIqOnR9x/Yw08cL2nltHnTvwVDlX94f5MmZO
XGVp04d0uA2t2l5HVnocNV9hfZw2e+lHjmvLfoPzkwg4GyTkPdYEd1IpRYhYf0+E
AxtLfCZCoqFaNyJueYVXasbpokj2X7Zxb+00hSbJsk3gege5CmzNjmMeSO4QSaAy
p75cIMZ5Zjm2WatpqIMJq0rmw2OH94k9RIWldINvJIo9esR916vYimTQmCt1u/Cw
ulqeJYeK6FFTyzhJXrUOPd35cENhD/sB6bW+MfInOqUfy3teB1A83OgPEvA6EwEm
onleyah+hz5pCDrnDdS7PG8gacIUL0cUm9JtiEaHq9fpok5DRd7O7H7gElu0mpoT
7aBNNyWSR/qht49m1xAdvE8H9U27fa7uPrrEsxZbWIPORRMPnL58DO2OO9yXraqr
VsbIFvs8e49r8evtMY9Zkf5f4xKAzmiDY73qQ6uPr1cCBiPMiMKZ8fIPXDmlzUpz
Lqw6S39i1ubEn7d7nf0b9Xbga/2dqhdw9f1GYmlvEHuJzXEZrTND6SGIkjdyE97y
S+KPGNJWOmbWy9uYC9OwgcOtQhyi3MHwCmo5cbjKzlQBkdO4j5QsbpD+NPhO+Fyj
qwFEcSthM1FkIPTS19HzWQlUgV81Cf2JADDSRVKWf9C8eJi9PIF77fQNbzQnn05d
f54b6HF8bDdwcca5E97BaciHdwI6sFxDglT6DdyCTEKzE8G8RmZxt2EDRYSJCYha
9/2buFolQGqzWqr+8L9hIlPIVBIioZ9LM0Qx8i/S8pjVwxQeDxDdTHYx4m7FZeHQ
Hy59dBCHpONr7hYWc0RM/ossg/6McN695jt8nQLR/UiZXKOHXc2pbMfon0joz+ox
exXJp5tDoZa6SKYihLwUPWaOFcGJQ55gpqrYzuqZ1foh/9RA5bmQU0iIqx4ZZzmB
u3l+aOXudR3Qk7BRPS1vu/8fLnYxpUbZHUoUo9QuA/tSWoGx5tsW8dHErQAP3P8f
wF72pyqo1MoNdrvan1EendmpDFvxqPpeZmZkzGDofXkEQmKJN3tZ2MPf21OMvEio
GgDjyLmgjNFwZuEiUjtg38L3sD0/3qP+fJZ72wvPHKp+G42ExuDddVLy1bvPaycU
aKMn7X69FmUbkzrzNyeIU9zDy9D39pptmD3XC71EO60a70EV5BOemWmS1TsjAEIA
EKxggRwMJeJAoArZd3+no+h3bhEHhxzcpAHGWfXgw4B/+1gSMRHHbvVh1NMEJRft
5OmKG6fvHUvjg6XODWsxnzW9P5l8iR23luz1NM+NGLsGh5GMypBX8fPsQf26NC/7
4BZBQv4KPq+xTy/WyoL7lhoeC520ePJQeuhhkEMQEwx80Ihiv6E3ua0oBcQDmy9Q
VvN9IwbiofyIn4fmGA+VSNqWpTJG7TwHk7FXKO2aQxW+hqOeYoAoLWKuwcXVQrB2
3ssEas7uaaP+NDMwNXu5ajtsrI9OJ7YslmPklDX8YWe+v8e0osAOeKbxRLSN7tnZ
H0xMJ4qNzbwwjnqGMi0XcMWxgGsValMH5P7s/xfwubkuMEyoMucg5kJIcODLhQhW
a7UUILyNdhmRXu1m5Lu3id9Uraocfd92dg9JUegaRls8Q34+O/rxQRbpBsSOxrxX
YMbpgiy268ZzS3HmuCnxoL5LAwVy4x+vkPjLS/CbViZCrcOiGymfgAlpE6G+iNgS
eyszH4vxHpRkRBNA+jKE3MlS4I9NC1tWfHKJ5lzx2LV8lU9f/H5se9zhI0rUXhI3
1Vpy8PyzusZx/+dbmI+6qbqHn7Z3m9Hwa//5pmwwKrp5Y6Lqhq9VdzgLRugTt2Ho
8vP8gclincwjigClKm+kUBPssWDN3WaR12EPXqES3LBQgGvEHFoZqTGduR8Pdrv7
IviScwTMqlmMUr0pZtx/BijJxr+TvtM26h2/P02t+ZDAMWBXu1NEtQLxRz9NtJ1m
8OA4vdGNNLueRI0cE7vfEO4zneqQmu8w/ykvMMMYLTNydfXSnDyvH3ryCRI1vEKd
MnjdBC2tlKsq1JGaPOBPNXSnrPcidENWBK00VYoO01bGN4fPT9vgwafx8grSGJFa
nCV58pzlIXPBkGcqu7kMMNDFCjx0ypyCqk+82VQgS84E1ENINkz6ohZeUTgWTAme
xdhbgDt2U+HRUqwD7hCxLMMIV2C77RI/PZsa/H1+BVRBPA8NYYNn13mZztFQWvHC
IjA+xCiAu262FlZdAzkQuwdGJnUtP6Ect5ezg7119JdImDfaKD1Nr8N8u1h5sBif
bxWSn2ZVYo9ldNFvuv+y/WHN44yj6PXH9OpfRD3rJzrqOoNi6qg/BpijhrKMKf6d
r0sxKmP6GbHuYyZH9ZFZJrSI7RxgAdv//5nttkXemstvzwrYpL1HaCyyYAz4Knnp
eZaSUbyywoNrQUrkHpWHXSUv/TRetsl4IrcbnEDssu4aPwoJnZ+Oyn4qcjA65yPw
jq+aSbaiQjzjsjIjaJIz6rYl9AKow1IwwDMLj89lWAKyoORWwY5biQxbfvOAU5zZ
5PyEfYTTvGZcU9zsFqhLtRdUHMScrr6vWHBdppjxfNhDxi1DxOaWpeGiNelFFb17
dnaksmtJfdPFchWLMdNZFIBeuZ8jyQMt7Wfz8udDkX8aq3V1IuyTjIGUr57dAIcH
u8LtT5UUqyKZHogJyFW+NofKcnvGFHONy9MmNFj2bPhiveeqZPdMYPrUcqufU1BY
+/wV5tU4P7NTVhQR3zUnolTOuw+EFrWwRuq5zJT36uE+99Wzu2oDAfNWdVCMrlGu
jE29EovXyD3Iv+gy5Xs7A51mq7qiPp8LymeKmv4JCky6cKLU7+MU5Hv8MRxFO6qr
A9KecWxHaUbfdlp0THn1u4bPOszYVRe0n2nm1k89rvqFft5713Jaacc0+mjD+Kdt
34zzpL96jILgtrVXdXedmlUZoF0grMC3dw42xbatMKf1GfiYVS4gI1nrPNJSqI+J
OIGHUIYU7+N6PTkz7TvweLJr74FnwjpSYz8fOj+18hCO0fYBTGm/yUqBqp7VetbY
MjDXkWtwIRwRPXyAn9QFlhJe1z8zVwURbPM8lcNshB+Xh5CshUESp8BRgO3l/nhs
tb0WIgF1759FLx7OqNLqmLDpGxJQHYz/JhgnHdTUS/UOybUpKfgke7oB6uCj5Tim
3gceTVjGP1A+WlAK5cy1AvYxg+ZVsF3dOAbBS/bi8I7gIyigbfQGKVdNqy60pXS9
qIn7KwKIzfSiRW3zHuUzv1ckCTMz25UOiNoybB5nJvnR3oPHtORn0EUfv7TYXmiP
HBcIoL8Pd57qrqEf8MTWaN0Q4V0erqs0TrMU+0Il51V+2n7PUT1s+EDhj2UWFFHL
ao9H2sRp5TwqGcdfZFdViricDAFzWMMfRAJEVMghWcnCVJcGgZZNZ4xq9GLVQ4Nh
xTJKvIpIC3zs25a3ac/RrET7+0jeULxJjTMFP6Ra00qov+PT68TC8hieivXS6fid
lGTUVuTviY6aM4Pe2wpG3T4kumu4e+iTMs82t0YNmIIj3HF9QDa6O6i7qMyoII0A
`protect END_PROTECTED
