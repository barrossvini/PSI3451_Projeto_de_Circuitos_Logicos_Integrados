`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e+TwLEREqxrHDfcqg95Nfk4gi8OVkVxivY05xHV6DF5/z18SXcrmiwc2L3Iuh60v
FOT9vIKq7mpQA7GAlc9JY86t/hrolTI+WnqSd7smQjl7YrxB0MI3S/2JKwvdQLJ1
o06UJuCRYXyjj7kqUft4oO/pxT5VH5WcHjjVf+8Bj7XGqQ8q563Vy9XFvcxeaBW5
zXP19CKpkJ414iacG+X80pheEh+sJ9mMru0vBMGPeNlxwOp/HAfykCfUl4QXP2aP
IBNLOkZdKcXDFaRo1hAQ6udlweMUX9RJl6hVxlaFJLlUBoXKFtCDzZaIkMHaAJ8s
+iw8Y6lL5swDm+8a7THF7xSqs802oJIqcq497h30YjNnNOpaKVbqaUI/breXF+zl
m6I+5+Gd1qqOMKW57rdODoC50ittOg5A82DNmyehu58HFLO6h9ERtNHAFqzBcMhe
voS7fXb1o6riLL6pRknqpVJXI/GTw4QpJYZxHvQvw1Oy9j/23NHbZkHJtH34m41b
qhIrx7v1stkcGYpbafxCDB0oXIKBm+SmdHFDHGwrrsH/frww4UKv6rb198mw8xYX
xTH7/rY2GonYBke+yoOPbZ7IBPZ2sy56Uu/KHSngUEwIk4/i61dg9cEsRB+Lgez3
Dl5N3AWrp3gWR+CZa8ZiHeNXZqrxRYEplMbxjSmt+Dqo9TrPyRy/MY8qvwKF7ydd
INyDBcfgDlIrn+SaiKvifWVfvqIL/JCLnQrY98pE1NXsdUQHMVMspONkX4VoIo1G
dL9Ga9wjzAfgn8NzegG3hamCWCsglFyI3OWsvAsEDVKGEPLO0NVQbR/e6vrEzgzx
JS1hYYa+se2/+3bO2XbDhfmOJ4j7AZRRc534/66A36sgWrR+uDoOEs5W6romn9iG
3V/M5XR+R0tGqmonCOA0mzwIbWqX/q7sXQtB9NsGVfwsPxKATkinj6SNVVYl2W+U
VgMImpTR9QVSh8Licjb3hlnuHvbsdRuEMPcbhCvkNoziokQ6Fb2XMsXv9a12AJmH
RaY2m8gmmZnUQxr5W0raFQ==
`protect END_PROTECTED
