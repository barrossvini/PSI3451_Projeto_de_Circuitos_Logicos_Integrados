`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MBOw6nKeDtbmuJJuOytuRksZJjPUJLDbnYJRcMnMLDT5tTRIWpQQKFd8LemH0DfV
Dc/1vzF0+knQxPjfRTw0lYPJF8ydHAh6HzSGao/LmsLrYBPndLd7Kt9RiuM/YDVw
n8e1zB+bBLaJr4qYSb8c8uqS7WAvzjWlFukY/zE3sOA1C4K/BGNHVDepv12R7F8A
Lyxyu979vUCx9Q1kmdetkJJkJtXzrG9+IYh/JjhQz58pJmzkqKAZmOjmpLfUZFJL
5+hO4q8E8f4rIBKP5f0ctLVKNnYm3I4vli89iL4tzT6+Fq9w350QPjBI2dtdwrmr
XdNt6N+9t0SIFAy4UaiVvxYTfd3f5Ehl5sBXHz9qhgb0s+EM+RSoCqQXoHU6kJol
tst8GdtjQlihZ+8/ssP2txn56vF2rCnVTaiI87WJzSapJnv5WYIKM17Gg+XW8GOW
NncnHSJQEJR0AGfN/tuLJUZr7IZ2eeEi2wRAd2au8E9xss3GoyH1Hbd9hNCaLGha
eUNSLbBeP91VPcoDyt3Pxq5LmYOiGPQRX1yWU251OlGz1DJnnCFUxDiLpKlPjo/6
`protect END_PROTECTED
