`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WmfOFReoyDRDK1sCE8ffgmIke9qU8oM3uoNv8QKiSFqHjlgWNYjoJYqJSZlmsvL/
YaaJTh1K2Whghq4aKcnNSks5bkmfsqidL4Qi5JaIH01ioIy34gE72Dz7N31GVM1Q
i81MK4zPsnPY+pH7bhA5MSSqNJeAUHddYaJB+MaZ24YteGvDQEvrlkC+olZPP/Nq
QbuO6W2XZrwp7/1OyaXntkj935B20ZdMWyUPW1UKOblz7Cq5qovi1RVBxx+q4aYe
ZZZ65xQD9fxiEXeMmQNcl6+Gueu4jR/TeSFFYoF8exasJ+rggY+KZWmqJJJmGBse
UTah2Ib2NRVx0P9d7cTX9dflZbIrMlbgmqgX7ccmEoWaXM7OxTmBi0qXQaoImyAV
o5nVSjTWaEP4tMcCG29ZDS0aQ14QNe/wtCfle1h0js5Tv4bPGosiz/HJ2b8nt45Q
kiyknIsqTcrD+I8Wr7dMrSzlvPndTkAR8wHvIZ34MlQFwPQ18+6zLO2Q8eytn271
rUrVbxMn2IRazc1qnpDVZpBT3dIx1GqvyhQ+N/IeCERsEHsxX50DV6qhAOsd5hqF
PB+N7HDlNVY99WKk75OqIxycJVw4HKeANqf27HC1WL8DfLMkPeqZ23HjyiBhA8/L
dx/aNou9uQGJlzsOa2/Eg5IHw4eOt+5LfqOHGLUPdKrN3B5aZYNgX2eVr/tEfMBE
45qjaEf2E9kSWUQ6QgKBL3duZ4QmMY0n2CMvPoiEmQG4GqscNq1WgGbWulJPpFBe
EQmckY5DJs4KguMJHNCMXbAN8zQuLvUkrvKD3QX/CYxfuOk3k0cVz4GHsLBzjIb+
rgfuVuKFIqWowIQXLiU7INLxC7wrYme44EcX9814FNUbXo9HqvNtn30UqHaqiYKs
TqRKeQRoslp8MbGxsk+u+EEqWjc/tcTgM0vYOVsj6yl65NQQwrZg0YLXd92Xzi9k
fWpZ38to1/ecyiTtyl/ZSdKViVSGGHttEgJMw689IK2p4WG3aIbhb0Gzu0Q4j9/y
1ovTgmDq/Ir8oZK11enRAPJqlAVhrLAHLHGEvdrLxFJGwJOsiwIYfAecmCAmiNFb
T6P+HbvJOlMjYFmN+s+2AoJamqmU3NsHOd5+y2EhwcD6UHRYpb1cFcnuBXuP/lTL
4Fsfz/lVB+HYG9DuC0EO/TttL6HkjOvgFI0HRuz3qbHbHGqDHn7B1c78dlm5JgUX
5G3VnDCMkgcrvKDGafOPECrBuV4qtk9xxfHlRU0qaxqpV/4TbxTygruxl9xPBN4P
ZbN8J5zaG5SoNoLW2RF60Y0o7WFfUcOBx6LvRJ4EjpeGgDVUyp9k8IKyZx7EyLRf
K6SstCo/Ob5gwZJrzv27f6fWeQ7GC1zIiPp1jBvP29dVdiCElEdhIIPKBsUNLm1D
SRDoFhMNTVQMIZsE61PeJPXkA3JA78d1u+lTkiWSc6U5YIwqM1k8jTv4MIuZXieR
CPPVZqT/9Gc4tuoG8BW9cdWyNxqZSOQ9gFY8/EW4pxQWoprtfq6fISv5F9w3VUa7
bjyB+V+DYDJ1+I/yBXRG5819Je4emI3hFL6IjDXtlGRjIBGQnMzmJl8kRtMRQDjB
HyrslAXZwMSn7jKi369W7x7Qt1FD8XjFjNBGLOfGodN9sKiKra0hdf0BY+/5+Z+D
QwsnFO5f6h0xz03JmM3qjw+29ZLnrOpKq3qfTuN+SuBU72eWIxZ9jjM54Mni7ida
6XnTPnUmRmCYji6yUNuQiU9FrICxgVDDsWFr5nGjIhTVaBuEqSXrSGo9mT1udCoT
WbIOU4+5TrARBk6H4RMRLql4T70eUYHF6ssgx04UjBA=
`protect END_PROTECTED
