`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pZRLOHpD+2BrdvHFxUbtG4azqRVezYpZVd5eIfxmBGRpHCwCvVw4DbbcaDGI8b5i
KDHbOQpZcA/9eu9m4zuF7p8wnr06Ch4FD68s2nIgzRDlRp0Iv4UujcglHTf+UVMd
WlBcOPO3CzwiJVG5oHeitSMKOkdlOE7VQii/VrlHOO2KpmWKG2iR2mgSBd8Lc31k
X06e8/z3yiefcSrcBILm0DcJn4qbZkGzPE4NMVZJESNwlNsySLlb4KsCJHPuUXbD
J4MSWnYlK6OVd/8XBHXQ+nxqcXMamFu7Cg+dEivf3twp/hYtH0+bzSjtwjgqt1Gd
gfqhxQgjp7Wh/AW5ZgFrHCr/UJf4itQ7GaSzDMcIeg3bSrRbu/M4076vl+do3ILs
LBjJ3qIUbuprkR5auKQoHo+YPMGt+5q/Ptiw5+gdZHtQ/Li+8jQVWQ5kAFhXAn7J
tFbg7wLr3beNjlZS+JDcSS3IKSbArS3eAhozreALUXz6a8BDNqTRNF8dJsY/pkUj
An/MrtJOVqmoJemzZfp2dxsOQJqqjRkZYvnXOkmLIrMVWRhA6oSVdtodcaOBECCa
COdlaVZ5AnHOvkCNGmrxR0t+0LWCRVf+WQFuKfp5A4G3/Gj+gw0Ls0S99i6IkSWV
BjPcsubPNp5xmvtgaETG6GlrZNptZNwaPhxwfyVGLBSv/RgaNPPqoSbF1QPMkJAQ
vR1ekj/4m3C1cD4AlZlfXhZNT3GCL8XS+DtUBNUppsnm+tIIdqvE6DnTjZnI+g7/
7SLjy+Y57APXpEjRJn/0Jc/VxlPx8i1so6zJzVMUPm5qZrqaiU/NENyPFAdIILvl
GI9b+Z9Q97p6SlN9JYt/a5YUpcmcFoKtA0MraVY5x/tzvfI5+6tVhNA3x0QN8UF4
tw7bRXLcGc+7KRs3PNDSqiScVBKC5FCXC0uCwNfEA/b4OGQnPWR9YMvedb1R/PqK
NwCWzlyknDJq5T6CgXkZbz5RYoo13Zo6oCHIYN6Lfp51RI7q/SVUFiZWqmNKE2gw
Vwvo3wwHJptaiWXr3TGwOgjAcRP5xNS1RRJTyUj7ifKCJMHMOe7XHzzf4YMlskxm
mqwfEHV8n1jPENwc8QjBqGF5q0TUTzl78xMhMUjgcOn17hWtL6g1zKilrGO8rM6S
KmJ8aS+UqfRNQji/Z+lmTT+fFtrnyemWv9HsBcgp081XMOfJTxNlolyIXLgEQ65A
aTNNpwwe1i5IgcxMH4lYkd7jED/0A1XFlUdg3p48n7k=
`protect END_PROTECTED
