`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
171Kj++VT5Zp9s6YBhfV3ETX8p8c4Uhr27ZvVi2KyLtUzF3mW01G8S3410N3DG/0
WllnMcQOola16RuGWb2AWK1AFdk/7DZNG0qdHRTMoo6krfFKNddJpKZYt4ZqVyWR
zB/BKDdcH/lZizXNiYiCqJNiIgKF2w/4t37TviM6JG8RP/WUKzbnQ6/5k0EgepM4
v8mYQ/1HMNNRxc2GJaIPNqniEEHcUrUAWeP/Z0oqjehq9NaWGr/v0M0wAh6v7Fu2
0okNOEpwJxvDuAEj9JRJKr9hRc0jiLFVZb1XEZfcjOQpN/0Ep75fJao4wa72oxyi
ew7Bxbm1jQO/s86lIHA0jW8EP3UTk71dkYlI5qMNE7Zxb7lXEh4nhqL654CUqM/M
TDNO6lRb4OByNuCtur77BITiJT/6eg7fLoYEuBzSVq33oZaibQdaz5GzZWsdtxaq
rhn1NMXFZ775Hp7Ds1zEWGpItxGJl/0AQ5h1MQXPpIs/h7y0ijKGGKQjxHeNmPMv
QFq4N4nlghE8oyR1sP7uBMBU/Qs76Tqwc3KaIk1oh/vn0CVH/Hllcz8xZl8ExF9e
sauTNedGXKds0nCptjAGL8kEa+FtaZRxa8Bt6fJR1/eVwXqHrpCXMTQ8KdQ3AtPn
x4MKkV9fVT1rajBqDOcy4Vjf5ZGiVKEVgfylxPo93H4cTK/kCovsG1EW5kW/Ljfg
C+gO7y6xcvPyqs1t8p4XS1URkElpoJCYuO9AFjJWQicHyK1ftB34TnTt+x9vOgam
Ym0WZ9cibQaMK3lTKxcotpnyYNczNv+BmlfFPVRG3CjROHc2Ki8NAsLkuGWXebOT
w9Tn2qbYWBZyPCNjppI4gyBxC8nzE79O67Coo71c9g8BjnbAAUo7AULHLfNpPzm0
WHSvZpxWpd7sUG9wvQM8WI8yd8YtbW3rtql+Izb5G5RQgogJ2vD61wnusZDobrjq
j8dFU+1PpIC5Mm9d3yi+vCJ/nh7c8NU0k3uhAD/SWjvWmYiK5ijd9rqVtc6h/35W
+eCnEdhnTnUKsFqLTq4aQEAgfLWEIrRlvrWkWVy0A2MoRJLbK23F3LYym18Bxl7a
nye880O0w7SICs16xvYkZqP3cX5sjxvvUWfGHCh/siOFU1onVLnuEqWRKRNJE8YY
HiHwoCouIHiRgaU7krCF1g2Y2ud2J99E0TgnSJbO8TQvm2pfGiF7fDD4IHx334Ch
b6Av4mHw2kob6eIIdEsvKPjJE2D56Ti2Zyob0MhRNbOYxZ3oR/pp0y6xglm45SqG
4mdttTsURXydo9x8jcxllj2V5xyNTEmybUCaHom0p2zDm7Oq5E+XeHUYjrHOtGfY
SEwsyg4RSkj8HzWYjgexpXWMJoQDb/VXZlEe7C3JWFeMDkM0ZdrEZaKHABejNy5D
LtAU5bnyQ7V0RjZpe917kcFK8QtL3pWr+XB9/crL0rn5cPzWcJsXSZaRFoY+NBQY
9kxXILcUMUGzzbCcoT4Q3MmrRqf8/wllBUhBo2rat78Wr0cl0d8qWwuPLh+/3z4m
uxI5tNsv4BUVyrnX4Mee3psUHVXd4gssLjj163XQ19Pm/JWsdwWHF50qzO84NRTZ
iCMYJsjo1FzgiNnZ/XYgm8wQPZliZNdctfagdbPABwa2JppvClCQ1HV6qH5D5yT5
rUfcyPuHaKBnfJfDzQmQdu0D6irW9y4aBnu9jyfmxAXYQ1wAlHGPqRgFcigCgI6b
UInJkuSyKXhCQtMZR7FrprZuhEFcOUzu92aIgnHxYIo/34nSUj0fqJH9A+8H1zGP
twL5DKZzzWOUNDYkL+UwBeUzUTlfSPN12aX/4DShnXW/XlvovUvjayttmTbNmZ99
guFD7qcuDiKIt2F0AJm1hckhaNCCpzy3ERPkEilFLrvzzoeXtDv6fj5RpiVJZLXX
snzP8rophgMMvZ6qhL52C3QQ+/YPRUDFf7Gt5mauwxQFlP6s3hdDrN0vF/+htQ56
ci8R+lXdwm/uV61flOdU3RbCcrAab8+lteOJDmewtRfgN2VrnteqLN2/9NBTkUIA
gd6j330pWqAjgbfAD2ErNnnPKSDEQaR2OE9Aro3/eupEMYyIsj7/AQZDJXC+doWq
K9dCYsZaAr6OOFpHePttkVNGZMoUPnZK6fjTaM2Lw0LKcmxgsXV//pe4wAM9m3YH
CklKrRynSybKRqkP2FvYe6C5oD9DGT1RwPJBN5rOkfUSrJen86oQN6DLqGw8VhLh
45EOCNXSoaKrez41lIMS/JT9tUCTBDc2wKFhdJN8UV7g8czqmo+J5V81x1LQew3N
u4Phi8832OiVfQW4YoY7XkM/RHo/AKJIpf+Tz4mWaz2x0kwRQGcjd5+xbgY8sJ7Y
hBN7EPuG53k+AKSxPz/zl4Iza/JpzjMsSQU4Fp8VANmpicUcu7K3IPIqoCVz1I4L
EqhRquhJXXsxmDe9EZh+Q8hNpErfSJjBvJ5SofXUZkNmKojA3Uvuya+/8RC/FFE/
t0VzH1t1u6PsYxj9Gs06Tg==
`protect END_PROTECTED
