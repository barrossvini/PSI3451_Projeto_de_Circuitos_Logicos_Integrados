`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UrCMt9Hl+OkTNAWh6r4PmJ4prAQ0bc4b1IrBV+khnkYFY5Ib9DxwV03m+h0ugdiU
qbygs6teVk51MsNaUumiOb2/DRFSHChPx4FPig05gT+YDxE4UP84h5i/RCohG0uC
JxJ6L4wGzz4NVnjLL17zuI45DE11dUvp7yaU1Fd+WLMl2M0yRlEItVjoORKkSkB0
Bwded9Glprwt2yF4/enG/5EqNIli8lreT3LWfVS6CtJJO2rwhQEAhXkW4yJ6E5F1
eelUDrVnGYeD9ItlcGDS6gKv1otfmrZ3RVn/3OfwT/U2c6Z0fu7ofdNMtj1mVg2n
a9sjGGjUa1fB1/dlaYzoC8DrdWZYlOu5mUaYjZ2K+NtlOvFOFFt7+/oSTxpA5XfR
nZ/BumRZPuu6JedM8SS8oMn/LYafrsFUM6Ee5Posj9xP1BQANM+2fkl3Ijbo3j79
WS2pKOu3PYTdImvIdQ41Q9Ea2pMPxDuRBaSlbwXUqydriUC7LUeOuWdAz5TUWTCD
OtGHDTx933M+N6z7aV96HXPMTM3jos7zAZ8/5ak+c23h9A+Xx8+co5MRIqM0ijR4
BSGVV/lhdnxuChby7n+Mbb6+3m+EWI2A3R1jSHJKFyvjSGLMfag4MgMohBaMyJvQ
emxIpu00+jPiFdS6FnbLm8ZdcE6aTOMZ+w3KdZtFVa3QU+YKdoWN151NPfWE1bbc
ZHPJlOpHbzjKxKOn/x7u0mwR4Sn+v1829k8MNLcDThgmEu3ePSikac+xY1A+lrEh
+4CfVXzKeo3oYEj/3sfmUmdosPo11WxhG+zpVaBVwhH5JAKSpGS1clxqsRNJVgRo
OJ4sz7JriBvzEZ+J7pntTDek0tJmuq2p0wcsfsgToujigQE5yxByI0ejmOKF7t8j
Hbzd7SzMAt0uiA7L5UVtNlr5URuUzg31BFOxMDVKaJhDue0Tg4txboTrhLqlC923
aubABTXhWY5BYh/hUKycVbxfoxRgY7ROFHceo+j0mMdT12pbwM9aoYsukdPk+8FP
zc3Jda2FTO/KmZlRkRjR1zNIdJFNXqOYySVAHoSfjrg=
`protect END_PROTECTED
