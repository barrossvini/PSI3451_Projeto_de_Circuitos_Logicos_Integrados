`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kEmi3+cBELuiAosHhnnHnY0bizPWowdDq8jJ8oRqf1otJ2mnEA5Bti5tAcI/oBUy
fH7lJeGFx+P/b9cS/DjvsksCu8H9ktebd+/U2uiD+9WbV6LAIDAbauiDM6BGrMvw
5xpZsChENcOc5K4/7Awuh/9pBtz8Q2TUlig6bpUkL+VK+cokwwTcUs0UiKL5viZy
BlPyiyqhq6INAWZ9LNGgX4CI9sgLNZYsBB7D05IGvXyqXrWCwOhVN2r/Qy96W7F9
T02pevRPnGwZnFLNX+fRbDWUkOiGOHXFTLF/6JePT+Xnc3uogbn2L0YwxdWpJQvQ
MONxctVuUav20/WvHfxKcq8L2qHZd9ONbr61BUNDSFlViaa/x4CnAFPWTx1M5q5j
7+3FwgMDJJNnXtAmzhcUGM4WxmLlGPWHEsRONpa1OOkZdEgiZUEwAs/re/evbMET
GKnSTDE9qqtYeF7oYfPHtb1tU+eYNQ/LYvryKsHHHhWnjF+Z4G3aGzG4vsaB3N8P
vDpQIEP2loG2AkqtxAm3tQ==
`protect END_PROTECTED
