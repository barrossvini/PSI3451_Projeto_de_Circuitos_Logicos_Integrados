`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DiKC94OH/n458KI5zCkrc10MqprbVzfJEx19qbOK0/ypv7ahB+eKWtzTV1H7WSb+
ToKlXxFwqvTk99STOdwuhqEe7aT2ayRroNDL02wFKtJJCJxQhoPF7BelIxaI7BJ5
c1fFEFImM2x+Z1Io8qHFHFnLxN1x+Cqt1y81+dhO4bEi9g7PGK5b54azdRsVfh0i
UFOVO9UBQ+hDantOd838uS9s0wC5lD8ChexsmD4IWqGrbnjCrhzAb/UcTSzZIAqO
q8PzAa1uZh8vSw5KnM7UDRPEl1zMOTMLRld+iku49bZmsaiIABic70KUr/LpL4pM
p0nejfynoH+GcG6PRDRnOUrYu5fe6V0qwtdofzLloqtA6nX/THaJzMfSZubWJRTk
/X8YBzG8xUqJmGmNZHgwJaaCrPBKfLMDp1Zrrd5GdXX3A0vW9aqM/qv6WmEykSF0
tSXzwU6O1epWc5w8ZhLAQ4eFJhIN5nvgfvj5mHQDDVQnTS5QwGLnoDHIulEj0hkh
NuDVxq/CFlKZNIhFTqC4ak9KPXP0kEd75zK6RF/Jn2vTF2vd8tZswd7CzKHOgknP
Vb9Fx9szI8CUf/2dYdAsk8FIydtKPDaEimjNSTeJpequTbtHHlj8Un2RVWcWe9D/
a4hfY8RjSw6W4s/1BhvoTosIFYSBRD6524imZ1HWov/k4SCsb9XasuKDuP64wxXm
9eFmJv9Ampf+I4ZBa2HfAv2KjotlEIdn2daZ1elCnhiKKkbStguBS8jnZ68Y6Ask
3zbmO4YdXiAnRb4WaTWFPvYmT5zGaudone62ErnTYYw7fKg2P4JP2KHGC07RiQnv
jOBMBSb1XkAiWYfQC/+49IOtOmkawJxGBsPizk8kvJp5fhLKR1w+uSnpSNFh2jnt
k6ymUjLRleysK16njCEKvsoGDYzCniFwB6Uzwl0PiTHylV/1lSClu4Thhr3vgVFx
9wkzoRtuyzzzFS5UqY0Ville/dbVcwEW996NVTBhGRPQMnSojko/Kg3Ms6dmFexW
RzlTs47FxMf0XKfYyjnafgJ1BrnwDADjlJNJRcRkefh33pV2VjYMMtHHEmjAAC9g
8+O/mYlHxfnwrr2pLu6HQOkqSXH+RMDYQwtcn/nxXHjbXkj9bLF6al0Nfwr/JVxX
LPQeuKZ8x/UOWPpc4TGt4wkEsnKr8FM6lIrZp7B/otYFdg58s4e9E1a4Mz0C6Fe3
nVUWSA7pvnWEYVCdUQfzcP6lJhuvdHv1vHbft5xGQKMh1rhSYwG9RoHWKxxOMu+s
66Vi9CNd5Q1DVlx3uy97xkE7Wuv3xbWsri2+H5pE9Im5AImCLny4G2Fe4xnDK1JM
9jMRiy8hI182SgB2M68FBioPmDOUXfKopOjSANBNzuHCUgAfWLR9mnxJm7OISZtW
ns3G2d7Z3LLctHl/iaNqm+0VmmkgZ2VUiaVd7wjYmyYAsO7rn/eHHVuF56IiykAm
+bHppGsuHk1TVKDIAq75fJWhh+pp1x1EpaHx4FQrqlP0ZB8+zrxECtLhUuf6ZCoW
gsp0x+wskGSl9+UQR54NZ1ULcxGa/JyHXq+Bb9pQFiZ1lPRu846YW6AMly9fAR6b
2ah99XzrPMaA0hdauyzMsy0mekzoMvBV/1XjBzD1SdDp/xIBBl4GuBfTFrBbRsNy
ioxtZJZwydgUIgT1S72ISYyycchtLwHls56EsmWxsmsGxX5oPg7FK5uf6m/eR8JY
B/USgBuX9YFcljP+jMlc3cxGvCJpcTCByHxWyI1F71AKAjULZUSZE2YmsUXMYU76
HjzRlmB7tZ2wZR5S5SXQ95ZbLlz5HrcG83rADKPF0jqmH0o7FCXL1mzPZZHTnbZv
p48t0nm0cQpYqSrgJTDT5NfQId8RRx+h9aK5jQRllVK5CW3QkusQyfN4rnfeHx51
oct2Gl5KBFsf9DFXo0e/yCMYEqOgTXQwKmYJKhuf4kPqmKUtq75wawxfaf0Y0VUx
xkg3C8mCrPdlzKpEOxXF4gb2StZYRAarZY/5DEqhcp629YfW+QLTVuTPxKlKxv3c
QwcujsFKxEDkHKpColxMmoEY5+UM0b1OJ+VHgQgNq2EszZOshOMmm2Q7y8lpQKbG
1uvfwe6LZsblh5qTCRqlyBVHMJ5mI2kstYzTw6n42Mln/w78RMO28LeAxb62lLHs
PH2pLrBd9C7Wgfng/BWhho03+HjvzOODiLPhgqyDa7ida9703vFLMfUQVnzCMDC/
FeEZ9mi74yeKrUIjx+hzb/9aGb/XFk8rD2BAV382ZD27lo4z2/VXMoOh2mo62kul
f6duGZZbXaoG9fMtYIBRPhGZWeDjHL4wV91z+Ca8XtpELLlw/bljLKaCaNE2euvc
2ss7/tm1s0lHeKFr0OGPZ0QqqkYoMe8JnfsiPZ4ZmVDd0KFu02lkz51LEopB/eal
vr+wJgfTDkc35qX9kSImwdwNRaLPDB0StVR94/X/xbTnmhT2Q9zNHWq97KexZ2rd
ZVylo88BekXQqUE7jtt0GLWtwNQhnlfUNv7swG48WYxd9F5F2s1Dg2D/1RZNc7C5
rdQNRxGtLbulKqSxzrg0XPUkZmCewP8/DW7k8XobUnhbPBkJRTdJsY9sCtL4Zxum
BNHCpAYrK81gQ9SRYFozMW3pWO2pvAkT2gw7eGIrsEuB1rSeWYvomG46wLgM3cex
WiUHaH1G+J3W7jiFcgMvwUSB8XU46vhWPM3IuLCEbJzSyIxHrhelUASMHqoNfZiy
lNYLyS5qr8HqJm2Ml4rx9/QikMRtDHIpX/WC8feGeQQvsD3/gcVz+dRXlfzWBGuD
tyjZ3WwX78/VhP5gEQ2JUtiQxDI67qPo5P1VzAa8UyRSlfHTSphH15X7PbdihcXZ
553OyrkSZZihOdxs6wNydSLadaQqCIrhTXvyYaOHRqGUrfQM7vtglz6bIxH49sBs
OpvZvhXyVs7oAFWz0VkARL1+To8Jlh/YfMmNxYmFtvzQKPGIFIFOrMysxFx4uavK
RgCy3bBPhS6tsx2gsfNqp4XuyPNw4h6fh4dsUOeVUoIJaGC+S6TufZ1xu2KxTR+p
S9jpRHKi9BE0Zh/L3wbZzaajTAmQjXid0wVOcY2RheaVU3b0DfKrX9H4jEVK5+70
Lhpu//tohm9NdWYfkPNXvFYXvbtEVGdfC6KyhKhy733b46FJGQkUbzGXf7KJHnS9
1my/0MCM+vA2MsaPwtBQke7yUQmYorbCverbwNHUzmK3iS3EH1xIQRxQyCzxIU3k
3RRfnsN2DUHzkYW3rdYOb5seoovhXCsWB7nnX9hP6t6lohxx63x43Iz/7EaeVXWt
bfTzDW8pQAyOel0fwR45HkeeHMORH26HRHMAAQ+3vwmE5hGZsW2S4Ita5jSTzAKN
6H/zm8i+vqlqkjzrt8aC67IA2SQgJ2KOSAkRGKnXCG2cz/jmIySjeIg8vM7CfmQE
u29iGwE1hYQwBYfhiWgpBe58yf/ctiURx+EvQMsPylvy1I1vRkiz2LCOwePOkXoZ
kK0apEkRklEjIvAgfKLHYswNplAkmFl1HDFwGKuLMC9ih3yhaLOVbxtjutyEaAsg
SOWGFQuLJVAOJptULG6LRggqp3ND+AI7n9OvOsPPsWDPNLednZVTThoMmWUnnaAE
UOnaQqd3b+QFpgqpdiF/9wEw4HCW6Xd715kBRmbBIE2Z3xK6BJRKlw/HGnv6eDHs
zqOGnhsL2ZBjjE+rU9liuDEfF53D3fZb5Jrjbpa8sdZH7c32QOu2tNqGMjPU0i8q
6Bv8zr6lkdp7N6LDy9g+zi7isUtjyc0ZDb+Ahce1YN4MInn+L8/iDwada+nfsfGg
+5CcIfAY/6essCSJXGWiywlvHhHraS65xTXit8DG98eDQ7anTdJ1B7KdBs+Wfx+T
PTJSfB7cLGroFzc3GJS+9c0A9N8iVqoehHvRqCngHvcSreFsY7OwK6LxmDcLY1J+
tjtlyu/04PxuIZ1YXNuZ3VYzdW8xCd4X/Vu4UR7aibIW/hLqEKy5DqK1xtLX8OOI
x5gIGgm8i4H+ZHdGepRBWE9GwV9q7/k1nxi4+RNb6CgZJd9vg09a7kTrn8o/oJSR
+Vw0MI2F76SVxX/EQBGLZtH245K/6zUn+iWXnCfI7yXMYn6/TPJqLYyjH52wt+zx
8iddQVmCVo+FAyh2G8mSzv1L0Jhjn8sER3ESgh28TZTLOq25n2N2ug/qFvM4lPyX
+qWvpHJkcL2dUApFz+iCR8KzT88HuF+vVCkDUBXS7KfyqZTTRohhiJQEeM0KraDx
Br8lt2btdVGwMYDG8q1EWXC7tt/zMTnXRsP576sQ4hybLML5zoJEvXa36PH724r/
KNa8WergB6ah7BdrQAR9w6H5qY4m/pALqr1YOXFWOC9+eRq0gMLOIXudB9mnehRW
foqEDVoPLykippFsSuezcc+jwc57uom+5AWMMVd7RGjSiaNTSCdwURHqO34WiD91
uqHs3wS+wBlQoolTFTQucEJ83fqEDf28TArSdB2YVvHfYdmN89N4w77k0dyCEA+X
bkV2Ua3YrJjE0Kegl8QRmPEjPG5t+fsf+3s8PHkp2G9RC3ultUVQxYsuNDEezG6v
VhD7oXMZuMGEr/Dbc2RtHnEzIcfRPaEa0dIt4tNowfAnEIVRZ4RDdtFtuAiWvvTS
hUghhG+SORbsQcMgxCgHzR7f1zzeLDLmtemj+W/r8CIm/KGh6uKvr68WfBfWXQXV
D+yaRlUNJjW/tyv+3IVHswXulk58uQuqPD3zoQEMBDK3oH6m3H0ufDw+AGLgnQ+J
TaHCwQZKaptBjYj7VsZ0OCu5//5tjbywuSp9NL5ySZ5eZ+ApkAGELMg+S9iht8Fk
4BXiM4BcmtIIA3+dTS5fZw2/JlAUfXwPW3G1q8KHl3bNr8S4GJZrEXxagPHiOSmZ
LW36EwihRPFbAEXdPVbgbLSXW7TcbPPOCX1zFGypkCtoSp2xnML4+k4ydZpThk/e
e8pEPX912uKlLkzcqhc6K7HYfnj0+ya6rAZ9DOMSQCv9Gt2JaMgMSTxTETET9YQg
Iw33QlB8OgfgJtDIcglvcKnUX6QsFIi6b95K8Ng6S4rYcF3ZDIlmbLdrQrY0ZG17
H6qjRW+wpRls2SeTJpeFhWkygtG9qh04KYCMhyRi6IxnXo+jxJed81NSzlw1cwNm
AFY61nVHw+QRjgBWXQlsbh3/4wldrn0+/OIbOug0yAD6KEQEYd12OAWDfMFnCYwA
QZTV9ET0MjeOqMV1TsU83RamH0Ggv7yS2iGtoQsj2mbHNwCxjFylLvNNr+NC/G4D
SJzq84rJxo4CIA/4vWUN/k+gNrrqwrLMf4/iXQb/BJeCy/GoguwWfyIDyT4nS8PN
sf/fqeJqBYnpybZjwFVhMP1CqzejxW08yoqBaAH+oPrqhArzSN7hftONFA0Dvd30
8LWl8mfuXZ5EkI4rQWxBLR+C0mFC9cIsD4+Fdbuc+H7lxzLuOVenPPk3Kx1z+4Gt
zlYYqr2F3OqdUNKTRkXzr8RRduXH+sQ4zvtt8CIM0H7FbGm73ZsmVWzf0UBHKTcB
mstF8TlVnpryxGE9Nbzb8PuW7eBhHU4rWM7Im21pFTcygmPbb/XQq6dVY5oYnpdg
TirVxGCWJY/HWFIb0uLM6yXhqvw1y71RmiArkFIwxgsa1BC8GD0AEKjPTa/Hk/DS
hpdFIKQ0NxeojcP19Mu7isJZ63NeF3bPvgyWjwmmlh2kUHIX9ZGYpy2A1zeq5R8N
9TGHZzv0RLgn4ulgO3wBw6Zv1lPk8rXsXRfjPbZ/kX/iaqmPP005h4Q4ecj2n6Lp
ebwNlaP7l1AyofW26+2InRRraF3sdci09DnqDjOtLQBBcRvkw3+KPTa9WjG9tnJ0
Rh9Vdr2lMCkErcGtbFhb3UT2jM5aWn/FLv3bAiePSReIHvaHHkw6B6/E7NXnW/mE
5jsGbe83DKDVgZSn1hlqkVeySZgj6oG1TSVMLiw/krzJeKA6LBPNRHqA4JtCWuKl
73ZzADsRlQiY3TwCwTcD8zEMGBanNrQERyivvxKK1gJevd5IbV3wpmEhvhe7Jo4X
Z9s9gj7GJ0ssJurp6nd+mQ3eQQaxuPAS/HS6n2SIsZ0TUc7f4CTpxBrQYi4Da3rJ
ipvSdQNBK1Uu6pLX197JgksBUmGmOZqdmMYdLnkPV5J/DqfZyd8yja47KLa+nvVz
I1pZXXgMNEOqKMBb4I2vDK2uc4EzkURjfE1kEvPpWQ6ov9w3VYtMqhYys9TljBiM
bVDA4VwaelteqlRdijWMgndczlW9BxrMr+iLFwyAVlj3BujaHdg9iKP9Uu6EQRqk
qcbgm65UDH1lTeggeZqjlBBRR1aCA35nhMsRrgvT/bh/zDCP/TXzWJ+5/fOc/K7b
l+IvmeIvjdf+XXA+9NrwrOJ5XsYX0uJFHPKqBbBjzv3G4wmKUCbJ+itK0JQkFYBO
TlELpgVgRvwOg2hISydX63xvy6TzKKNXK2MzrWDbqOY2rEDm+qhQtTZEpvsxW+c0
3HFk9b0AnammKivNP1ArCAyzFJ41z508ZUR60RS4PZhCaUmBwRdicz1/NjuKG3UM
riC1EZ+I6rOeqdnSu16k/ADyZOQJFnMWBB8aVtJbknigi3gf72vBPHAevnOSBrLv
W6EFpFsyVRSe74gsSysAGo5G4MKm2GE6f3yEYzIyismVQ+AtPDsQ3NvZeS6Wii8Z
BK22fUhi31uxq5Ky+wqDhpkrZSJ6WZKsK+5Vl/e1eNIqW9l/D9Nge7gUf89aoUqf
G5qVLOR73CjeTBp/FFLYBE1YInZuMJ2KkrNvrpfCcITaFYryt4zla5ADgOAUluPF
PtUWCaqaSkIo8Trh6e7JFWIw2diKtMewKRRDVXUGcuWH6LY6FvHaT/suuAEkqN47
QKe09NpuizWjKKuXqENChSk/FYi/auCxJZeHpvFZzCI6kLS94B30chcM1KscSUap
qrIDCkXYwgltm3ymG2yOZ+qqV0uZ5qmy6q/YqCAuZpU+FXHUuIFX58TtAkCaCOeJ
CLjiTGSF1jAeQtX3RozBVA29aTSxgcWP1xJwwIfJ+S6TnKbZ8QVzdo323teO5SH6
OhxrwzxuyLWfyLyD3C8jW9sSd6tuRhUz+pZSGy8yidXMbSB+0Kt1SLDhVYA8DJnE
Tb4bh5sc86Jw6W2ABOBQBnMJwcFoSrPs45geDhdleavgkKYceuwZ9XS7wnAhwm+Q
SbUxPIt0M2lXCuTa799iGQGjx/v2wDJ9qvu7wByIZSVWgeAKeH+sXOq7AgR+zaHC
4/lVDlLvb3ZtM3wi9AhLOQ65GzrHeTOGVe/f8hrMmpbc7bSiHlFOOXWx0M9J0P/H
nMsiKbf+5W2zcZUUCkCrI8vWmR9qZ9ommxDIN+rsbvCkOQ27pYjQNDqpaoHN2GOE
VRoJYqxADgjmgbSAkNuxFyQpb5p235hZczO9edeOK7bqu/VSv+gOUoXZ/rNZTm+N
d6CUWkrm+riW/MR1FmyZyHH9wBpYvo1FJzYkdDPgQ8C/OfznJusF7yHZ0rRmcanf
IrH1bOXlxL9Cl3I3EKXg3+GASAZHtUuxKfD6KHdozSFZ470y2JjeK1qjYALRIAbu
a4BUs9J1Bze9G1x6XCIhv4QNb9cZFksUaVxuKrrBVKjpJoTQhqqFyspy4jAlQLQZ
Dz+Me5cCkprGp8pKCdKNO0FT5Miil+VbefKL3SSMyW2kDz0BW1Ir76BSQLR73wV2
ckiR3cG3z8q/HVRHZKryIHyu1pvcK6mKe4fxO96ZEM/smZV4bOHTk4JmEeCEumFl
+9r7o9aSEt0bAKkcgdC9r8qksC8xAB+H/o9ZpAp7iPilSC5rvVmHLtJMHl5uXv3m
nQgqOmRr1v+bqBxQDUMkRluM6gaNulQuPt/nJDjuhMU8IWh7FNSE1PaQ8B597YnA
rnXmivOKyvngXpC0tyZy9f1vGIpVWx9Rwu8LZpEO9+5xjyltqcM3ojKYdPsE3tKw
4uckl3pdaUSQ3hdmaO1UaJ/KT8pKQhT0Y7BdpRcxv20Oj1KxEYuGPkGjiO01usAB
T6ok50tkcs/WyY5L2elqyi7uMM24NKB5MX97Z1OA8zmn71lP8PPNlk2oK5X0jWQt
5ctJ1PGC/uTu+PMnU4xaEmfM5EmE/ltOTQpfgKShscF9JrkjyHBgympqBhqe1OAc
jQ1oSRdHPfDb2kG6E4ov06MFO1aMzDu1/CAb+1SY+KTGVl+PJrceX8QdFI1pjCst
rbw3rSwzweCvtB51TzLWdXlH9NWFJp8K/gAlLPJxdo/YY8s+08NN0LyLSuELK9NR
Hun3m/Wtfu2e1l0MAiWFixnSFGWub7eEsT8JEnI1ZiAgpMqqUp4SfU9p1GwqZUpb
BYmdx3TVTKcBN+2fdm9jzZHL/vUQpSBgj2LQKwe3NTINrHPPc9fIRXZ6qSfxDqWI
lSI1ctEMK0AXeSMTIViBAEaENblkSNPYnNFFJY5ZoWquPr3majASC1f3EUwDc+8L
itEUwjaVnvAO8ipZUrbD19mA9VyyWhkGzC+qsQTukRtwzGZYe6DEcJrOFbTmEaeM
n8dNsG639I4dj9g73tWIpSg+uyjMLBq1cXHQqwRpVtcprpzOYT1xbHXV+ZW7/rhB
UZ2vl4GRBgQS2DWEEE/CNrI2qXlijDhIVYYcR5BJiTINCkROwIcJWQ7FTOvw9yfy
gG+Sb2GhpAvmYlFS1XjOuS9yKdZfj0nH0bGACpp7u3kVpDbGcGcO0f8s29POglXI
6zAD7maI9VH55sjqqkh2zVg/EtwBAUDhqutG6b4XDJu/DsPtSEdGq+v9YKpmOKya
v2kO7J/Xl6FZeAp/hr2IjQSc5pRZSkETKEuFXCSeP+c9/kZ4f7wBeRJWCzs3w6BD
xMYSv6e5193ygcgiHYKfhi+PcsuTAEN0gugnoMfCtalMeum+ksBVn/dhqihC6gGB
JqA+v31udP743y2BULRXdPD+1p7NFDPE8Rilq+W/155M9PKeF9ztILLxeF2ndE4p
GpKtqWCmW+Ug81O8GD7jcRHpeZCx5juHKAiTcgXJno/sSFHEGKMmheVLEZfLXBco
TWS8QSJVMa1PHZjTzUiUPuzikkK0LRkiyY11m9MPwc3dyoDnDq06gMYx5Oug/KiA
GAat6ZAUxd8DFTZ6bhR1bRvTLT5ygkhDfM88xmL+iqLwER82m5Armexr7PdIyc3F
6sdzwN/7HVS60MbovBYjSr6wb+rXrc6QJVRLQRTAmCwZEhBpgyUMROEWqmOika3Q
qQfr5QxJHhr8LKz6ZBxCIUU+N8y7yPHype2CgipL8mYXME8qW5t1p+tju8tgQSid
tObSZnXqiEawHtvl3Gsya+hpJfDAy1jQ/JyA2zu2ezz9pkNKkdZulNXJzCE+fB9H
CLasvFe0er/XDybur2232BAa39Fa2OUGqNDOmHf3Pu6QZ2zsU9o29liN04uCrNot
e9aabZdHE0x6LlxQajb3WjqLK+T8wgZmfhBdn/Y3XtLni1dWpCbY/vCkqt3Ilcfo
BT/LydgEmzpjkVjjAdVdI1pr003sVjWvkhHKjZNCGgCCWm11R7FUO7B9iaXPoS23
BaUiKdm6umODII/uyFO6JRY0xuiADtHhnZWJcLSzylykMgZMlIXAkLZvkGttkC8o
LMZO8fi9EFTPWY2nA4PT76PmZtaSgFeY7bW15U+VsY5o+Oq86aH0WBvs4XrYPGig
3ka5N1ZNxO/sVy9e1uctdkt/BcnN/O6ujSzhy6d74s74DnoEvjQfCZfY6fGIK0XF
Ijt6nGeyIP3mO8D4hjuHbOoJXwJbDTUSmdQ3A9lBfbAZCT6lgGQyr0zZb1P74mnL
8grS7ct2QJNYlPwxdymqYG8TadsBCMTG4omXb7gU0vyblvoWU2LVG+EuvbpPc7uD
kpP00obIhsOYkU8Y559bsU3mAVisx3lcN6VrcRGkJpCEpqyNwYgH4EnVeBtBx628
VxJ7k3thAd2Jl6l0cpw9Fz/O1PlOLxr+bKVSqCNyFYMg1gL7vssOu9cwzv7hXFQO
3E1n2MsjpgDgL9hIt24S7F7PHBzdYIS9xOHq+CB4PWKQ4b0vHKg7N8WjdUMV7yla
Zc/yoNpx7zZVc5agdStEckZGK+/EPeUI8CmoIqdtFr6W73S26WswBBEkHvcCtjH6
b1gW7TcMJt/RMv7esufYZt8kzs4ZrF3DuqYmS5Okze8ji9zmt6ms4ZnS8TOYm1Bd
jef7O2dH3ZNXdbFEzYURH57KwAOZfL8idZ2so0f2OREp95qJD9q7lAbgroFfUJ5W
nDjP0ABrVWu1+vj1/dDjMwVg+mlp3XLC6roowD/0r8GYUSR5feg2eJamgPQeIrRj
uYQJtORJrwd2wymtdrFmgEty5dlIcxhCEy2lR6w567UnCU6g1QUf3XKvXA6ErqBg
3+uckMgKMSyv4uLWniGMbz0S3m5ACEd72mZK9anJgll8UWosI8MOnpylJYYX9fMn
Jjz3hmYrpDIwhXST26Pa36ZSufDcUJhBVGO9pnFtmEUaU6d58xsnqr5yGonE/zJy
PEynkWl0rR+R87oxN7uc6f5JMRf5hUcJ7ir5jqJKOxDX72//JFswucFEO+ZBUpy4
BEs3f/rhjIAkReYbq2XuI749zoXhAXgv/dcG7HZFzOa5gnFknmRCEHs1KYRw+GDi
aHbD6HeZ49EYqeXr43TavbQQXIqNI9G3p3xtZDAvmZm0szXAVn8ERqIBv6PSeHBH
ASeiZNywD1vYE5gysFQh36tz3/wHYA1GxdXhTC8sMQUj2Y5U1wV2nAndzQlAOf4A
AlkltmhYlEdDKPiRP3fYnHZh6Fz03AIa+L7JF2Wh0VNMIuRgaeADzFbf8L7X1pWh
It1nxwUpmZZaFZfH7Y9TPh7G/+Thv63fyH184786fIK4c4pddHf3bQpa8e1lOTG2
p/mOmplsknTKPAjoxerHa8eQzhc9H6LAbSbpwHEh4y9DojnYH1NRAwheg9ArY5Xj
YmQZI7rbVVLQfxuzyrYckBq5JF/WAPBSuMJzJf5zAcZTotfto7GFFASyuAowbNiY
ekhcjpYu2NWhomeUJmcwBmA6ZFFQh7+SKcvyxO5/m2azLyVNoMHQsseUw6jvPJjl
ygtE8aSiu7XpinGfB2KCxpLnnDrHC2kaZm0v798Ca3fHkVtK1shf+BBaW0tQezr4
tr2ZXCt1hProhKfzIZZhrd697Lblko6OMa9XXg8w0NH/jZ6oPwHnGIUcvOXljswY
NU3IajKCdigyai+nzB7QZ3mvFe+nWS+Ts+ubWbtlMhtT4o+aZatvgiLnjRunnXXE
Usir7mL7X1EnnC6uT7LvOcBeoki2REVcCb0Ei9NBBLnpfozCsx9xtCHcQmyK5PTz
GFk9W6s4/SXL+mJ4W0ezoo2GQLSLiD7HgIc2NXx3vojrdaQ0z1mZqbskGm96Ru3X
gFh9LJEe6Xb2upHAE95IgDuFLuFer/jRVzQd38WZbIQhnfgg9P4oe6KGH5li9Rri
y3O46QlPeJ9hpR5AQX/BtK0mmaE4BBro4qcnNL7GC36QXNoCxoUL5OeDZuaGocAJ
FjFDtg+3ErGH0gF/s1wLyMmstw7gPquhf39JYRe1C72QMSdtnt3EsgvUeVyDxYsC
3GEXuwZ2lEsUz3bRGOqx3HpTDZCOO8KyIrrAWaGq8vPYdftvpxi2rY8GilTh9J3H
/CBDfVyXGAMqpN2soinrK/hfzsPZ/rCwknB6o9th4znvpVLOKB6QOIs/L8ayCtCK
VisnjlDoa26MpFncGUO3qslv8ieSzmn6p7IyfE/X7z+TqrKzueLbMk37pp5SVC1u
ujvzApwreL7KU84JIWZTe0So/iDB2orV+ItTfv/ra/zg3GD0RCsmMZPw1PXR0PC3
ElX2fIl6IUO+4FA4H8mjSVRUbF1e5hj6WRQFZY1eh1NCiu5o0LP+jEcyjh+yOiL8
3iuBKZ6kUukEVwCxUrhBwnIfzWqIXLBIBCzovzNTHbUsbvlPbZUbCePkF5VfLqjT
iwFigR/28Dr/uiWIq60wdxBiE6aLDnAZSIPJpkuqZ+l8YmVnZT2swFt9yQSMKNf7
WDxoVbxB/sP9rQoVDvXJ/U79gxzBpOTu3qdZKVLEqUHCGJMioWaFs8XXUums0WMm
1UiQ5fFlxlfMC8AkTKbd6J/O+MBoO8vq6TjfcSwlhV4feIRdB6pJAyQ6d1fHQcl2
AYwBrqBn5mgcSFOD+oAmWrC5yruo7cUXmL/sykzySQNZPOzwPADcNjI+eY2yIohX
+dCgRTqlQK0w9IiDC/hQfC3MCp4Pqjnfgl9WaulcZSVpW3hfntTwoh/EmTIE8B9f
8Dlfee1BfHq+6UFOBEk5aRFke2YTDsK4cycHwGwYEW6E8UptoFjXOxKKUNCrWstC
OckYzZw/AFJSS1Z2lIFVg/h++Ex3OPb3ZE5kvBM4WZhBERyW2iT/05byA9M3DgMT
MA3uM0/yEbqSbOYkdLCGTDXBaKSnU6qZBvCANLYH5k762TWB+KrrAS7KNi6pefic
NsNE7wfINaCoUndoKkvhNl0QdEyHLuNsNu7TWnD5LiRc+r00RKybkF8gLD3tmtU7
gGgDUaoUIg/VCs54oS+jSJZFF10OY2PQQSvMplPDQb7mm0sgvCjrGumyxnzrlN+D
Bhl9irIZU7kDI4RhENmjWre4qvB0/tcBCoxo9Xfg7Wv9U7jgzgeXBcyjB9Fa1lgT
ATwdthSOo8v2LIHVgYpCu8k2jOga06qyjA8ocXrYFZOMIyy+TxayU9v2zmt0KvhL
o5q7kSlLb7azXGewRUziKA/R0/2c2DQQQoc1Sa1YYboen03bRW6aLQEERxjcse6m
M8zk/d4I7ftRQ8RKCdGQFdJmwmMjYYDp6//IzQJbiPG+FtBoU1QvTVtJ4q9gC3ke
F5azAtOTYNl8mumgZcDZ2weclYxLvPkFx4e8KB0/fkHM/6oV35r3takfZKR/UYix
c3yRSK7ncuuMyfaS3Tuf0sSuJCkepUOnRVwYigesOZ5kkGh5kOf/guwd62xyvwMo
AbANZBqCMRjnAnZxPrfpEzuU8y6O9rhPkwqAs1XaJ0VHfXcJzq1YDoqoHDJ++h4R
4QLa4oWyIkOS8SnmzQa9YbyJ1SknJceG236iVkIamytP/GdtBe5qeFc0+UReoTJz
vsvlK5Ojn4D6wAr01tTy8ZvUoRltaqMgJQBaE4fK1QF251cec/G5CiK5jGysAXGV
ZqtL1TlGusLv6p5q+/gTAnUzs414+Cf8pCTtwAwfw1xtwUIzAiapu9CaZYBvJKkB
xK8RaeVr706qgDuee1bjhwCpXJ+5m8P08w4UoVddRgpEZpv0Qv+p9z6G04QAqRRp
RHnwvUDWtBzVE6llxwD4lrcpZbIuTyBJ1Gsy/1pyB1G/k4HFjVcqtbmabHmTHBjY
bAzOqTtRkF36AoNSxBOhiZjVOigu72DtWmVuzxcPmngv2IqsVbj8xZ/2T6UzgPIG
qjqz/t981oKL2Zm9FhDRdq1zmVnDbOyePaTJ1qcjMMBQazG8ynl3036SdvMPcDjm
Q8bJQn9pagmKD8fNaUNpIWvx5h1W7tCVBLcZ7h74zWix3zp9FMyce+llHGWFz7Sz
8PS3aHs+R7ZdGB3/CezSVrYxTY5FDqfk1ExzGxUo2BF1M6G9nssCi/GniDsf4s0I
/Q1ApoJaT84LsMhn1+KHnMOQrM7PVj6ZMSXGF1Cta6EKnYyumWKqM+uPVFsnK4al
/3iUBh2nRqorQV5rTM2DOBGVunoti8h/jAU+WLoa6wNGOSqCDv4BwVaon3MTmeCu
tzxuUJ1YLNHVZvzym9K93r/hUGCznhx8DUMvqNGpCLhYBBdUXjK5xfTMoLp57VYC
8oypCCzsMQPm5F8AeAPhq023aU193rMWDqGU3Eo37degZn/onTmG92vRyatOUMQX
nQ55Fyvqoj2oVelmdXs7ybFKpQM5t1mPaVOQAv7V3CqU+1+LevqFkCtnjZRx1gVX
fGPIQhuaPwl3ARPSJIQzcjnPEUOaJLAr69FnlYwXZTy/LSq/qMDuHmvS950OnH60
/XIDTcjoGZl9OBwlbZzGrmBt5j5nZFPPOh6q66e8neJpmZEVrBevAtAjJ6c9qN9o
Nc12gtP754nyGGC2vZ5KsyI7KivqQwdEAKV7fgaqJmvQdwFncWZZtzjolG/xiSDf
cdDNOfNBkWiMIFRQT7T5ri9IDybN5no155nY3zdtZnIAy3gBg+3Hk1jn39jyAgIH
uZaclSny46vbHCcGz4qiUS5uw1WNhLspUoxw6iwI0/dB3yZQU6xKowcIgnBNoAZ1
xWuUlAnosME2jlQ7S/uAco9Aq9QfNHzZziBxz61yneW663w8/YXv+NGQo2PZUa6b
N1D9FLtsQEed4HIsxwj4rYFMpD/1moJevhag1VFU9jWkysfqd516LtrBTZh38YVs
3wP8a0Sc/GyYlHnGr08vQX/LiA5jyTfU6aJDrY+8Ts88G4lyqD7ghPSyCge4GTjx
vvT6uElvWRN/cT1kJhlxrKxtdZkG3lkfGMKxjgM3bAAcbeu1plPiQMPCF2afEFy5
YmO/ePdwSfnfYRSg/Bpee/kmY+SQG8A0skTclwGpoH6Xlsh3F7mVIl5liLeTraWT
5idd1pb+IeB7GLF5ygi6exw4SJZmAOaugf5JwdT89UsCkGwoUKnWAH1Y1uR3C2Jf
OPLKOn32sTU2ccqXGovtVXQytocHXEltfYT2D+cQ2NqEg0LfPWSJCqJReCmxwRr+
g4XzixVCd+nEEIY2OqWUoOk8toxudxyHZJSGNdV8YxrEW7gQU9Q0PlTyBZH9JttJ
ulLL/Zf+fyA37mBqSsky/I1oqiSb7G1t8mVhdT5pEWTS4zVit4IKCNspqvTUd6Go
skdLur2IfquJEEEtQtXyI8mTNkwWT2wbHXSVTGy7OUyVhVTzIw4ypLgJ1zni2irh
kVdfc6EEaMp/SkMBsM54NNcVmdDsPr+EElnIQuUNhkyX2nCORUDAOXtfBOBMWxEO
RB6MF0U3Ohe/z5X6Qg2oAHokUCUNJvKP8VklSqkKj0dyhMtugFGqvvFeLdA+nesT
Y6SXgh9xzM9lD1znmfzNtOA5P86YW8+nN5I4sVGDlr5jI0X1gwGLUVl/x1gGRbKa
A9KzD56K0hGZJ5fAXYCxiAMJEKR/2bQhggkqjKT38Yo5Tw+zsREBb3SRThxxwf75
aJ2QVLtjaIuMXC8Qb83xzkmpr1kGEMDJM85BUkZPbC6pTlEZ83z1d+wlZC2Zq93O
gfF5dhTddYgn/KPqLpRTnzyLCOj2QxJIEdRgHh9jEM2RqIcRTwLDrenXmMc06+7B
88DaAcgY7kEmlRReR8Sgu/Xb9pGwjXNIZ3/j279Ix3thVuYs6uJy+e4jNc9pPfYP
E+CsSDnksFyvDySMc3g4z5Z67naBNNxiakw55kZQzUMbUYBuRy6qbvP+kZU1kpaw
vUDVMLzeKSygyC8a6nR0b1hpFwLck7rjAJVm1e3p31+KlF31uK9oSUfYVkSDDfIT
gMPZvAQ/I7+wK90RuzhaznigJURkew7OsorJaDXxRZI6baA5zkNu5vMsnGCwG2rB
Hmwnid2Bw5sIXn18bTQ9bYx9GFS6aPLuxNCSP4Rq1cs4yxvixqcab6Cf6J/sM4ez
xhULqoBm4+cl7tLVDxT0YR2vJhEWYOYcSGw7Eq8K/SEdgQkjPcUVbsPEmbpwjm81
By1S6kfHFRML161e5ZT2C9NDlTupfbd3Nvx9QPq1BeOZteiBKXHHr8W2zUz4s5B7
tqISbTdYPTEH1J6c3GfRV28zP298mN48NXWykN92PTalpDqDhK2WBtIYZRkLlh+9
TNL1yRvJXJ2OWT1uqGUGLo3XXd2VocydgckAz/ICeb4l0+CZT2iD76OfFG1CqLFl
A4BW8wxK6KHmSsHHxltv/JDiKbI0/EYRaawIHXwrqxCDSag4fWdlda+kv49PqsWU
v6paXbjkuTcKrCS7U7wZq2BMUNmDvRQkNcxmw0jxLm/95Y3JWcY8ovNlSHyS1ygW
gvHnsa6Ta3intmv+8spn1ZShQGQlPNg/Shvfx/lwTmQ+Yz6yXKsIxr048KISZbFF
zwPsbMT522gebZ6EExgWusaL/btmTHtL5dNHqdX7NOJ+t/bmN6he5MrPXruAhHbk
fumhCchGNZSn8iNGgau2ET4H+02GIFBWmMOl8x5p6ynpO9BtA00D78h0QiR9/QTM
BZ0A/os9k3E0d7y1I7Q/gmfSV7KxIL0b9OImijrs/YZ9lE40n7JJSh+lIwGwJkTK
UO8x7eGtX+3pCb5evroe9w8skAKdYUnQyl1nFvS+tqjbjYnmll8qKGr3XM20ruYW
6iJgTUob02G/rtBsFtQQv58DMKmSF3gJA/eca+Adq5Hm8YvDZ3bXp99k5gqCcnPw
99xhAlkrcxtfcvcJT/F8srCeNvBpp6a5q1EU/Cpd2ZLnUrG+fdwqWAsvWl93RNFT
ZMyH7NiztQlz1It9iwZMpm6ocaiRwmptXnEpQF+QL3th75nbK9GMuJC8YL3kKjBs
Y1Ms2t4XjWQ7uy1KOQ7DdH2VAYwTH8QIwiJfrdOxwPcEgL/fjLf66jEg3y4ntP8i
XjD+Kr875mETQVcb67diyDCD7Pc+FvGiDZBsnduMqWuRBj1QtcVseG8TLl/nv4ez
FpWhvUbTEGQqhTOMgpYtkvh3ytL6jHi2mLQDaOMUVVb/NJi1bCnurcp8lH3ncCRs
1qDS1Yy2ErN53euzEiPwLC5xSPGXMikTvH1znjeYd4j/I70WN5AXeuJlUVS7twCH
5A+ESlRAAMSEKSIgbQl8iGJNCLOhCPN0VcL8YTBKn0hz+qB/z19nzjhCjf8EzJqt
nbqRfqCTXwFmILqaW+zu/MmECPdi5HAyYw1y8V6sdZvyn5n4BZW0Qh3JxFlm9gXv
ieN0hT2HTlI7wOC6cmKZzgCYBUSMLJPwH3k5eMWJeHUCDWnZ3YKDGbT2xA7COpVV
odspfv6k6ltmPP8UMjZ5VgVrTjk3fbfaJdx9YyC38SIHv7wd2RhEZWAzvFa20Hr/
GGiqt8S7cV3tAGBJVNZMWdxDSPBv78Az2rXAKe8fbD1k2zLtxlNdtBW/3sOHoNnl
Zoi5c2sGDynci5zNDxzR+gdVC11Daf1c4BNR8HzlmGmYYj/PtkkmWwoXlcuul55O
D4DUzc/dKG9PMVumZ02PXOaAClQXqcf3GiUNAUD38R9m/jj+ofdaR5PKcrrVIj7s
aeNOtvstm+9zNuNDVw7VJW/Wwzj/7hGoT8Zo8XvhFwhrILnCnDu2VZjU8l77A7w3
59e9gVuOv1wydsAbKA+Np6lPxo2wtqvzuBj7D4xK5kJ72gACfdXBh/7s6qKIv/8w
NlhDH11oZ6lG4zT8lMHe57iIS9FNaTWva81uVoXR71NOof0AUv4oSBjz2lIx4n4I
smIpUORWl+52ogB8MFDHw1PlKKcLfsKlg/iWCtMPt/swynsn1e2egkowctrermJt
RSZbUopORHvRAwXhCLrRTH8a/I9qbbYEH1QhmPfn0HgHETNm4GWPiXfEViyEjqpY
OLNrNtmCAc4kMjcj8iQpelXOQCEr7A66GL4VejsHpika/m9fYS3/UxPg00vKCTFI
IYJ6yz6YOVXa2w7454fvAw0ekSHmsnrE+CCPL9fa7ksMUbhxxLLIvoqzAEnCoriv
suReiN89ehUkoRHytFTsi70nAnMQ3Qf994xzj/9OruHNNrr2p5wcHCeSz2bwNggO
p1GRAV4uSD7rZ9GO4E+GxacJyIFreqEU0ep6HXR3mnR8M8VQV1khbwkgtaIt4qZZ
EBHNfv1xomhJfhn2s0GFJf/PtBde1YVE9xlCC/k9ipPoocpKTw6jVEqqKbJ0UJgh
Y70GxiHcQKQceW2M9Ifwfh6j7lnSfWUxTAkAobCLdjhU5Dm/AormNix4SCjZ1Yst
pWXXQx51X9JfW1pE4pWMrc6vC9B5djbkFVB33hSX5uOz0PvZRdQeDoBKdtvYVEmQ
hnHdD2TawGrUCQNpzCuI4ZZzpJh7L2nyxJpwUC3v4w0W4pbE+ZSflDDI2/Fa1CvE
wgwT6OUARZIeBMsBD4dnLCkyS6RhZV8AuJbGqkHrnw5Y3BcgURzXWimyMTCiaezj
BxeObKJwRyczVAQn/V7tAgMudhG/Ddllu0lav1gvwx0Z0Ko4jqVCRhHRf/S462tJ
UpiZqMiG6H3vLHKkLNAi/2a6LXnf5wq+U4fsgCsIxSuQfgrs3vFwbw3O5QHvCOp3
jLTjP9CBoh0n0Al2kMNszL1dUHjnUe5QyBcHjk5+HeP/Ccgzq98jvM0uZZ4xNWfb
pRTUJYwCEeRy5neb63S1sXQ8WZTUXFhzYG/w3lRBiRYiStG5UU7uKpeRAfXLdJiT
8MCdFpsA3J37GTx4F54h7rxEJQFtSp6unamLCWHWLTK9EE1iWkQwIVtfVa+DhO3c
ZeG+sLWiTNXIlOiafJmIR/sQwuszuRZrkv1+Wgl5gwW9bzGC5LZpQE2ANxlWxkpB
CloHo7dRydih089lz9nUJQXgT1p0XMMqfC4NmtY+qig/OZHLJNSVCO+WEn6eHYFe
sHtsGaogF7OqZjFxrDYNrrLZ1qjbe6KD7NNDzggb445owlfFl+FnOPYzoJqYsK5O
gSkuyI6yc/D0iFBCZPXW8+YmJpR3suoMuSGDCtLImfy5qTEGE4BqKHfhPDl6fQHf
JfUtl8m5oKKwLW9KT/duX2O/m24HvZRN+otLSYvbnH8WWlC5Qbdon81VxRPBErd4
rv/Qo5S01Z0odafzDAYmVm6IPAQRxCuo1Ue4iAUgaUyRS6v262TwGnBdmUSMKmZU
fkPvIkK3EpkH6zGg/en4ZVJ3MvpB1uGHypAfLCzRcu/NiV0iRW8qk7rszAipl+3J
3iI3SDD5m230PNzVorDN1uR1tlE2QyKgbliuBWKTivzhydfF6GB8eJCJfcAyzquU
RSS/XQbLvPYSj0cmZn/Ivf89wpGLuNLD20wBaDYLP9sR6saHtC75gcDGr9yr6apk
s3SNAiA/31w/mgvlsrk3rpdyjxGDG8zB810548LdPrRkvH5L5uptdOt7CwdQqr4e
sqdElWbo7hy4hQrB8azndKYnMAnJv/K7PBIM0mTCrzKd79FtLMx/2rlHP/ZLLYMc
LEqzMqCoZIG0d65ZsNr/SX3uS+aSuIuWEN8yjDjoZu5Y5KLd6l0GJfjRf3xklLQe
Q0aZwItO39GjpTjdHRfs9nz8YicmwMW/kY39pj0kwrUqndp4rrXatTS4iNGi49b9
awc+jQiPWiV2nuq0MR5YBXSRNMveuNIBCxfRiXLX6ccuUe4w0ilqc5y/XUTAEdx5
PSWFyB17uNuxTzf6SE44vNRKrf9HNj2CDFeLrMlUy+sKYM9tOIIL3w+jlldCfNC2
ckt5e7cZR338zjOqTT6BJeXYCeFzhxAxSldshWgU4ZuVbHe0N/iNHsIyIEuMFfCA
2Irv+BmPWobteH6kwnz85APVG5MZpSdY5qGjjLiQahhKoC/hKBxsebBHymAkj/hN
mN7IW7k8xt3L8jKjD8KCycn35clFoDzVjU7MiG8Fo1Je9o8VkkuM20w1FStrE0Id
beRl08OSEMs1s7Hlb/o2cc6eO0QrrIwbJ+qR3bzyicFh/EiAQjmn6GGKYEAuwUis
ZV8KgPO9AyfCuYTaZjtSbil5xbcTm1qoqsEN+HCwtc7OOEszToWHsOueYJpDQkua
+1dj4sY5+ly7dUJ4QtDQvjV2FbgWOySaaDZAp2l53aAa6i34mGrMVUa/vi3AR8Xs
8rHZiLflipb15WxQkJgNIuw+5NhxYYWCrT8rm4hqqAOMHBGYaeDj30vtjlh6WzoE
O9bDbF5mLivlaM9Nrlftkle//LpEOJwPvXYU8cVIoOOB8rhzbR8RLlhcpP4HZoWU
NzgxjFNcJ0jMnpPJ9HBwBHq0blQBojv2GfCm+IMMpOB0cXNJIn2B3AHhDkV4ehC5
237VfQF4yDcxyYzPUlEUm1YoGrAYuWVawHhMZTrzm1e+iQbO5XVFMB3AvnNeDogo
S4bb3acG1Gtsu1HBLvpqyQWfomSeVV+FwNTaXkF88sTXMHfo4ERFeeTiKV7nykhR
BbGiP1Hfh5cj3fsnaYilU7W4w+hMJYTo+O5UWRrEBHo1PCAwj/CyVxjOfGJQBBSo
RpEATLTMZwtD88ZvYbDJ3aHTb4pycuc/XAWLQ6L9ni6qvTubeOg1ZcfLz3BUKUR6
CdmTr6hHu7H2CZf7ORAnVmUgfLMQ2o5KH2VMO6Cv3tSaNmSWMdkmQ1jjDAelVaQ7
izBzOz+orW8JCxLKK7CR87rUy09hzOnxXUFdPvglQCBGlhwRrQ5rHElWq2lS1KaT
DRhPukAsxyccBZMo3vnsW9VUmERZhRapSPaowilBfHTzU97EB7B2OPDBgNrWp7qU
VbcH24+gPKOVWM1ia4C7m7EWpiYP7y9y5/lpOy59WYm00cgrxe2Mcd3fCAOqxCKl
0k00HhNxCHpQvOKddVU7dukgi/pi2AAxpVWCn9m5wrUlI/OYgZ1aQoR5GlXmk9UY
ZWaqWDXysquTPI3oZQOEk7WfNweDXyG68gD4g8Jjn3wgVOZYFg9U5UegJA7okvK8
SNLtItI8Lw+1gq6Nvjq74/lXFCv7ecZ3Cj+4dT8G/mg1jF7RE4BzQOC+w3fYkcoq
Vipo9gueSYoEyyrj7WGvKeU/2k7CPg3iFRjA8jip2CBYR2PRauB0rYzVIvSH+ba4
KHQMABvS3s3RRjcZpEX3vKzeQUT1fZIDaxRLGToIo3RevCJUkYSl7QTyj5hKJLdj
7jrmyKl37qQ4pjChisx3aIYXZ0/RVsVDpm1kPMKVTjdcf5tYSs9lVj+lEk7QDf/K
h9ZMdClhNJVjzGvj/UMIrGROrIzkgflL/o1+iSmwuoq4pKnTYau2azCXQekhgYsb
+a2I/QlknkHmVE1MyHBIOFIf79HcimGrdhVVkWNnyHZ/vX1dRWVRuVELFAgYDHwP
CCYmRSI5jyrU7jSK+feN+hnMxgzJc0NaDLSscapceobMR8XLMkYB4oA8kPQeCVGe
PHeyCqZQrToLQiKu+w/n2dXbpBlp/iKg/aensA9flSutQCSQFo+20g10d/vQCBMg
zaPruwXwQaJ1D1Wn0VbgmfiTxGoLEDjwwBVhceABPZ8xaXKqmzxVJ9WY8U24yuTp
jrJejv4vf2m4PuchXHn9xP8kgpdNZ5HOJ8GnAPJ7WEbg1c+8/PzlS0/Cg/dYpVJF
kWBxBAtxpvS4caX+Yt7IwfgrJjg6jMl75czgcPNXeJFL6QJMDOU0DTvSFyLELqPM
68asoDn8E+8YJE1Q7xyW7zqHhm9zrPCLg6TZIh2ryY6WmtktjCtEzbf+Dd/M8LAC
XoLgE5Ys4EsAiVKRcqjELXlp7jIJIXovy2H7Y6w60bGDsvsTTVT9Q1pq4y3LwKiE
iCamLIFURX4mdioC8KoEUe/9XjZorDGOE3yVhecqfJGp1FDBFl86b1+6Ek1dJMex
bLe8RNCl01t9uvpAffklJKFMlwkaHxDKv7z0B7DAp2Cdun9oxyOO76EMpM9Ed5fJ
GslKcCqpQXKCutW6oPhHfMYh+p8xuiOhV9vg0RMNxIeY5hbPoH1KT4mwa95itLVd
J/IRiy+XtFQcoRIoZ2sg/ef7+3Ayi5gh8xSM2vwA+nNjtSAjWCz+mgcH2RtxYPdt
1BgVcB6tviYLMqO17dXSLbyqbW9SgYZU89DDiOIi2EEcr+CquptE/+28N/I9wYhS
BYJhs099wEbjnY/DDxFonXwzt2pmnryGs3gEfXK4fM5Hb4/dJ5OwPLNBPpmrMrov
CUaiEyw8C0Apo0JyZ5M98oIMA1Vc/ri7W+Dilsj+IBwXjKUKx2ZdxH3rwG98lU8u
dPP7j56b+2bYt8eCgAGNY+P8LaI5CnUN9vKkLI+JUh8rz7+V4URhadMX/1n+obk8
qf97XuIw8Zdm4icA7r0Dsz4Q3sIXZawc836c7roMJWoLE7tpN4JyQfpjdooYfzBc
xKD6AslAF4Yms1g396RXED9ZopDfqKEZvBgb+iDJ/Mr8zOJunYYLIgGEuS6ogje+
k4oMJFPMNLjUEwD+k8E93nX6rpYzfDi9Cbefrf06yYC84WR9tIea0qFl/ZeUdxkX
kSVyO0cEjA8Ze2A42v5+1Ql7xobAVxIcNgDPDpqs/n+o/FusWzm+tdZq1vV17myS
ID4JPN2xvoPMcmHTMn0vKXBsWyXVH90lXBVsoYCj1n/LLnmcWaQ9843aHJq2XveX
czBaV3r9+0Fnb+SoUP+SwQa8cODQKe4uCRAD31xv0Vabg3ZkWCrlnoT+NxZlnMNb
dh3lPk5lElQKC60CF32TnwzxfZjysj1atuShnJOai5iODxdhj08T3Us+w+Ug5lDR
TsZONoPg0fk4Nox/UdCt/DCw+iAkBXfOBR0xjhA12U9aLskcJuriM0snPqUY5jwv
gE9f+ERp66cjRnfufqNNwTjuoPCX1X8HIv0OMZi7M+D8qDGAPyb0BjX86dmpvGzJ
S6+4kijf2g5CcRYMv8oS6dkuTAEvP/rVm6k4OvSLS51DBYpvLlCCLaCpRao4SK5/
lovJtSbHKt2ESsA6H31ViEbgopYWXqOZn5N+NbZNnUtmLVFpNTzulzDqaZ/pTJAD
ZyYLQTYqYxhByKo4GJFWSeIfBDfa8RAp37khffCD2g+43DP5sZ+1KYrkGnnM6A07
qTOdr/TfVpZvw3LFwMsh51QXIL+Urf72YWL66aht8Rd/at/px1yaKGIn0W+wAMMN
ytSzfRB7cVZ/9pYLCwj+gwhMTg0ZUTKepby8tLVhkspfd/pFHzsCSZHUVsZXSyQI
mo2B/24Y6joyzqo0Xg/MGNY2A/qt5BI0wd9uJIKSLF1HhjbkYz3pTVEgB0hVdzdZ
K4PBfnlHvidijVgkfgj076kKZSzqrRphChHFJa9GRTuRljFA7PwgRyFeQfDL9NLx
a0NsCZA1725DnVEx0++hwg/8qm/56SEfRLw7NslisJP5smAP5ZGshtV02ZZwrJVW
vUCk8IJi865Mht5Gm2tc9GtVqe/RfSFF9cVAwIyTouIpOdPmiDJdbCidtdPyyeDm
G5XuW4SHOaWEgth4C+qTePqvQyR+UtBrN63566dolyxzbqb8fevHS9EsedWzPcpT
iAVBKaQdKgMT0+mljKRmV/LvgcHLyhbrdUgKMZu40iP35yaY/2zkfdibnEAsr/+P
/L/mMM5L3al9JshIGSBW7fiuQG9NDe6V1sS9fUvQtJemnyqC+lb6pGJQH+pGQncF
emkaFMhgGOs29GxRUkLJz9cBsPFvO/hFX54SYbXxLdvnlanVy59+NRW8/kfid9w5
igrYBAa5dtITPfv4sHJMnmfmcxA5Da9STs71qtlr61Pe+mRcPfh98nvLzYvQgiHs
XH/OC9b2f2P7wDvz1C9wcMm5JDwGMRLOsQFg+DGwKOfXr+NvTwRKPCl9SNXAslR5
KkSw4GmzSWac55m9csArj3tCdu8W52RheIh0r0L5RsUIGAHo93H3xkgWE37U8njj
pkVuSrszAnRFJXqMF7ieXUbhvhI87RqVcJcYU7WLOVEsyOiT75KnbtQnojoW4niK
ky3GgI9JTZnHOmkcldVQnbRqRvvoVDbHU135H53ejlyuVsMTA3n+jqRGu8JIakTU
vo0SGQkM9jaisAYoiSHLynyIGFGFMHpTftGyZF3Qp0xJU4ikOpaOL1fhCXcw3z8O
KUxJzx/G9Jobwhw9ij7xXZrkfUej2yZoAMI8TCcmU8aR0YhYkIRWaRyq1m+H3BBY
F6XOaOKldz0LmyVO1fqEywLZF5BVoIbGFOxhOyyrrXB6vFhhlRIQppml3LIiU78k
OcJBb54ezzIlHwMep/nba33HHig9WvvHeDbg9RYWPAZVb//XHIub6dkEqt95v8YH
EQEuUgZ5eDYEVnFq5k18hxAUgzn6LdCMDuTpq9ZLIQ7GUQMzVlo7+fAVnXkP/GUK
D8y4wRmYlgW65D8c5YCAXDxmFbORD4EhbxQQpKasZxRo2aSB3mXb9R8ZirBupQ1e
3v7SKvOIOwJ71cCOm1+MU6Aase5YKCV/b9qpsoUnxMNlcEKctBU5w2+iad64RwlY
AfhvrZrJDYlZVp+CTgsUUdOJzfnXA170ukgdHb9cf7Pm8vFLJAFb5vn1jA/ql1eG
Ze+gN/t0dDEtaQbcGLQH8osUmxLq7MsI7Vl8a3hi1hszoX232VoqPOGALbgzQhkr
G/BMqhdwIfUADQjDxQ6+NFf13D+wNeoZMFPsI1RBtgUVJRrthiKXz7PIaemABcVT
XvjKZCMNrSVaxUdpOXS34YSb2HdOq8yTmdwKHqCqFzAvZF2DXMo76rrc6FTTGv3O
sWS4dWu7U9DY/f3gXPFFUnJdN7QwfQlk7xpvq+jXPa/Obqj2LgRP39R+aTFXNnjf
c3XUb0sI7nU8/ZiCSwFiuaug+jR05NerXQl0JWO1hz7PzCn0n575lfAQsnIQetIH
/qtYWxSatcv+4gCVkHMMI6TqXVYy+tnEdpaNMdrwTGI+hNvbr5V2Jj2NmVg6kqv8
jIxMVfsSPO14uqoNvqYR/I4CP+qSnPdJ5Vv4idILeOX6XTChUJOBRH5gPTYYkJIg
ATLeWlY3Oh6PmRFYjLz9eaImCX0XQhuyQeFMKfGkZyz79lHBbTc2xZ6BJZtJ9etr
6AW5CFUH7WL9fCrNkKu3X44wADQj3PDuk/j+mgqcxYxT0NXut7aDGT8F751TsiGX
TmvyvHsAMMAe78ia+fTJXuR5x2HCt8X8rohNR9Ltk4x6NO5epb5Az//x0e9zffvh
PeZ9a7nW4yb5jdKHMWX8h1CcI4TnH6Ew+R9Oz4DXNNhpW67E1yxPSJsx/uzPAjoU
h+74+k2j3BXHaU1XucbP0hwJ27piKbgk1KupIZRLCbiJLpqYouhnERL+sbIK62W3
gvLSkSM3aqGpOn8EX4A0YUexPOVN7jS4vuDlbs09sAfgt36B50dT36sds712IiHa
LrY37B4jwrVshaiSsBH5uU6cF2++7SyKRc5toTOwAZoPcdAnm/tUA1PBRgxKR9Y3
+eq3t0xlDxzuzKFhKNGH26I1jCgjLzN7rY3fvMvQRQZlKSVXLU3c/f9kJQ1fKfZ2
8f8b0w+QEMqHXMmuHVH/y4mabnbQBSFH3yi8Pn/AFz+ktb3ms1uqlF6JALl5+CHf
IsIXmb0LcZYpmDFmW+Q6PMLxdBM7l3QV2kM8b201ydon+042z/Cr5AKcwWxApyHN
1O/RJscO4uJyPElYSkJD50/3Bd8vtJNk7FyjFM672/gdXeDxw7zIWVih9f0Ds4m6
KanQq4y/qHMxX07RKB/RSXo3K7jUqsTSpYf3VNT4GYvHQ/MB5gHN/Ak2Y5NHAvIB
Hbn+5h92gQ6xiuac0rfdXeB+wqeWqcI0RAXsoKZjkIYAc4JjVbx4/pVGgX9Vicky
OYI7HzIvgFnV2069BlcgYENYSHSi2VItGfQaS0R0emqLfRULNgRuUpA2YMyHmSxh
ylW4CkV3wxzYpoWPzbbJd1+OMU4O/1ti+Q1yI15qRrfb9jS/uzmCzPS2HcmCs5GD
S2b6tuOw0LknmQd7JQxFKJRNOnr9ko6kiTs1XzNwW4Kh3J9pTbACKNQcKEKGQnxE
z8gY1lSk62ucKq66rJ9YI0JPTY17+ak4GUy/n1Vp8NFkQdpoh8Oz7CsoqxcAhUlZ
XaQ2nm5pIsxP4fgSEjXP/BEExnTxVhG/Glk3iQTjR4nsxABAuTjaTT3JQzTp8h7T
Jfbs0fyPtOC2dc/X2xYAZI87xd7Sy3wCi7qSkKu/q625sCCYXdiyYiQzU3TF+D7r
7RksLvaKMbK3yDBby4tde/E35G++BuCpCtf3pSzuEBdKmi5eoTirUe2bXmYLgZZ/
20oFZs+JFEPez4pW12xZJx4jTlOG1E0SWpq86m0arTpAMo3DRCrMCCtK2hkiU1Oh
svEzPZFdqKs6QTHAI/WdSMRGr+5QDIVNkDlKs35ZB8/TolPpHlE719K2oAfaZzgr
PaLzDVVvcmx5uDkAyNLQbUP6ohOZCrN1QVao5kG7QP8AQ3HY+xBzSpSqzzpzpUbs
xUM4WE7V2XI8D3XeMb7CqA9KxKQ5d7awjrqcou+ILQCbbRgJBlio5BCRiTpxpfK8
RW36ma+2a+fLAbcdDG4/HyvYHbxTINUG77peq6SGI3ESKWr4cfNykX815Z/TWoWO
1fMMc3+UrFLUmuL2pJssAPHWzZgm+sTn6OtzAykwN7exAy6IFBUYjd0vMqsCiSPR
4WB9s6F04lK2SC3/8yKYMHm+uQYB3nV9DqZYJo0TjcK/rPA0DPPD2uK2ncLkOCO5
7Y5icDTjx+tZT2JB6OLtgKzPQ+aHppslk8d2tnJDylbvlV1xaHADg2+ODXOX7VUG
cU6z5vGzCtH0xp2bhejlnMOyE8YgXrGNQPcZLdMbTEBtX0fL4/xg6ea8o/tQDzu3
JUtGkmEUx91qLX+l97i7ZbxG2kib4jqUNDS1mYV+mF5LrTXEHbzinJLnHABTvFqp
GJ/QAXZJSgRzoNCjmLDwaLShY79WRjQ9bRbInGf9TM+Xtf6PbczvH8zGlSsAcHfP
C8bkZA60KrLPTuuuA9sWOtBKpJEYzvgEsvdPcHP63ScClasf4VQFEndQvV/nzY1t
0pamcgKG1mne6VxGqCkcVVygKmD7owDaaur/sS80q6jz+wP9pHkdNAzHa5vampe4
ndi876NjUwW4q8b+cRW3i++zujPQNPVgepGmAQdDpfCrNQU+BgBq6e6hEBXg7vVX
j7JnQ8p/2VdWnIODHphHWkItj34BZnM6Z1YbUN5vqaF4hJSxkPwAxH94NkAWSnit
vkb/AweJLH6BmeM+1ICKSoKqPohzsGhEpKdiu0PgRc8XWqyuoNBYTLi15lGrsZfo
/8+rc9t/h/EfVCjUf08MIYO54vGxy6AOZYmK6kXMYGwvmOnIdqphsQTLHzSaV/E1
mHFZ5Sb3xVfjjcfMnN6ECjvmfsTYBOdLSKB5o//CVblMmE1gm+8VoxhQ8Mk9wK/1
IEth71BMisWhTWnPAMDmzjLt5mvMlPIDZL9Ipi2F9xyxaj2jryyCbppsJs3/MR0k
YL/baR9c3NmkcJJYFCIBdsUadOx+sLH3RzuUhNXwLtqn4pCGMd6wjcqzP6haE9UL
ECrWgc5xFCxUhovR1dnex5/4iTVVqgqJs4YOWWgBz3u4LEpDsH1HH/gSOOAW/dfA
NfJsXBXXuRijAlP2geDL7A5f6TS+g2xZ5z0bbq4IQZIjIgFcnBaS8Eg4foxbdh3L
H2N4weGtJ+Gf6uUaWUv3Rar5V0l2t4M1IxkoFac2HDLh/W2HKJcYHL9oGDeg6KkC
zbf0hw8YkIZYo3Pd8fZ0rttoheVCstpQWySg6erG2WwfmBIDCxHfV45rvlaZyiAe
Y9eHdZhnH+PEok1ASn8ebxhSJsikgYBlcn+fGPjlst9uvpx4ZRoMVP+C2nm25DkL
l6dZ6rnNyzSq3MHO+rZ0B4+B6AdEEUhMvdyW/LGpDowNNA2kpIyDkFUljPq0y7rH
p0v8h7t7xQvph49DhMob94EvhQ8R8a7bjkmVUBFjeF52LH3n/tXdms3/qrFI55bD
5l02Z8bn1xQnUTzrK4yYn+ESMYSdCX7hU1TFXQ/mPn6yNRPpyod4oXmodJwb6du4
5NMRODhpHS5o6gnAjjzc82odHhULl5hci98C4fJTureyExtTJJcgTet+ueB775rO
rGVWPtnjxquevmQakDMhvZpBsa1I74GGornRYW0FeNK79bbmaa4xZuANCwZluRYr
rQMjFKc276VheGuAO5IcFi4guMcpMXaq3L6wN9yp9B7oEoEkux8u5oAUEEv3nzeo
lqp9GKZpDZ6luu57grvzpx+G91CXYyJVxbyqWOlpihkllQpdejjI/C1hSV5F3T04
DPbR/uuNwnIdNK8UNbpAFWiINB0Jkw87R8JSqqEuCtiqUN0NIM15oxw+ENGP2baS
w7ZnYmDf6tXFQtRy4cTr0GcbIMbNjimGTrzQaMjKSCnr0xxr6YiMZsa7e0SxFxfR
/HSqxZpvTLM4cxOZNcMZaoBniuFldtLnZ4euN2zMn/0dQevWn9jvPYLtg/zTHQPg
xBbOJEtxSCtnuyQOFcGOcvI9zm/8gmMVE8wBpWcJC+FgJkMidtoq4zwyJ77jZZrn
ytBFxlN4bg7q7GBjzymkhaB7QJ4tfX7XWBBuig7yqtw73BGmlF0ZGd27vyU70FeN
OYPYeXqzt5bjyOQxHRTG2z108JN4d4iygMbOvxf4V5wbLnh9NH+KOLaPE4miW8Fa
2Sjms3x+UVGVDNMWF7uR3XXMCwWR0Cw7Lq+4qgwZJcovRSZS77k1Ebl9fmbAVLCS
F8CJu5TUwgn6p3dXQM1VKhflNbv8WAeDJmSEsStbfE6Yk0+pO+BKu/e/gepblu5F
+DOD1ok0uj9ULS1K+GYaOVD3dFaz7LgOmNYF4geBmYkJlEVC33ZoL/QC1WIt7ZTN
l6sPsnGfLryJbYIwQv+757Fgs4773izNFeaqSLdn+aLMP81q2Vok07cVePOSlino
eUnu7asWvt0wc0NcpX06xy8txnN/8JpOU1omMNOmHXReA2go9zjJJs0oR/TNctIC
iRXTRmrTKS5PzGWOBC4twmajoUp9lbIpNzqrXAmUSsOCJNusplXUK0uIZALYk3ov
+9TsQVMfQudz3f1ddE/wWHS90iUI2R9Bv98ChHxdlSwVT22k8Yir8PIFgrjE3jWj
Vx7lFSQi21rgOnUT2hRAXqSf7nsOR1mb/A1okjoQMOJFZN0q/5CCRQXtBssUANu/
55CsyzIj0K21xMaOslU+f73cIJ78+DCpePpW7tm2/2fKpgidDR0tuK+wkCDKg4SB
GIAcjuu4DeM0/o65ZSAuGVDeG1gut7xSMojVpTkGhx0NH42QN6+wNY8O7T3/Wc18
uItNeTcOhX8s9a+irp0jz/hehao3P4w9FYjmVU4B4sCYXIu9H1fHOXNrkJRSUM0Q
dPFQFj8ZT9rJLPHYGgnMQuC00PL7U921ZY33FC5hzddk9lsFYbsOyYJCDCVWPg6q
q5vYUpB2RuBaHKJNJm/wSWyrGV2aMLlajDydiA6RUzabO22cO5hVWQv0NbbQB0Bz
9/O1+Fhed4eyxMj7s85Vwnddv1TMe0p/s1KoeP/1M/ruGuISpv4MpjvatPa51koR
QjnmfBD08G+Y0m2zZtjKI+cAzZsWNWvaTft0W7SbYhnxwSYp7oUeZpurHdr4rH5i
+f7GwAkWh0iJgWWloiNEKEsx1nWu72Ge54Ym0UhIvdEZFl+v8n+MNTdVq5YK5eFk
u7NpbpmdcdIKiLMZrO4BVRyG2VyW2Wygyg8X/sX+63B5HCq5lcveAxbjv//QOkvQ
oZg67bEXNehCf5yE+eAxyRnaCS7SXCqzxZfMpvyKmj3enjEbatG6HDKP1N427hBS
du2tLdZswPttd+OV6KWlUbYqb5/obDbFdA1YVoty56u5RFmYeCbFggXzLDUbIIJz
QK3BFE8ARjYjnDtUsi1mfwe2/KL93hnLT9fP/a9fmmqa1PNwOMZk3oJUu48v3ui7
hKm0J+JA5n9tl9IjJEMQNK4aFNovM0MWgjkr8ZTyDpBArKhryD1XM1vIP9R7hAqp
2euSrtQXXlnHISLJ4tjhqfO8viRAJzWuvLcx3AIPBGZ1NQIzdjHA1a1zs0CjQ8uE
mIEJQRRjJEwk1YuLYgeILZVIZIjSxe8t/oTMFWn9GZKxroAVq+Unkm7afzkTwQz8
joapc5FZSGR+iY3kfRzdR7Xr/GrRQAqBCPZ6Sgy+62FLO6zTkSXgV9z7uNrWvPLH
rGZkHW/roP52qEsulkVdSqm8baW7u5UhPOPg7Au077j/e7MLCHy+xMZ6DCX/guwv
RNvhdxxEy3neFRJlkZ3FHjfJ4usjVJyIPv8XJ625ygUu9z10E1iKUF94Vx0mGp3C
NJuuBq5ur07lAC0rlTkcaUJx9vKttsiF1eQ7zG1J5azl+qrQRTkoNA1RkJy9eAoA
8WZiWQRPBGj5CrQeW1xXEUTKej6bwoHAVzYx9PxA2O7ngQsonxPvMkVoBsuE9V0p
j4BDJpn7xSq+N+ja4mJzocovC1BbMWW6ERRfUBVdwi6j9LkQcH3R7eaFVHn/R87N
VGw1iYjxJ8dlgT3TdOAMpjB4fQwRWRSQaHMaqaQuTGJEjEFa0cZokbYpXaL0C5yM
uc+1pz3gEB10rf8jgsncKm8wUyzEG/9xh4SijkMbu0xEAwB33upUMZ9rp4bhL46q
GkVImXk1V8KXufX/tBpykpqdCeXVx8eI5jJQ9w61+Awh1kJMPR9v6lODgXSCyrLJ
8va+FwVJJt9xCgI6sFq+CaK/zySBAwZjdoJp6lwpQTFjM7m3AEo80nDOjvI5pHaR
uvxB+RnqjoPT1TuKsuhvkBFv0LMiHCkUbe0bGHsj4IRUNiKS5m/+E42ilmxM3AGI
OICVN7WqBtpJzHtDhWby+JpFyF0SAL2HOuK3TyOJFXyvgHTMFp9ChyOQhgm5lJnl
Gw2LV409SimVM5fjtznyiADxF8ED/IsYvrdG/Okkz1qr+8JzAHvfhV0EwIyMbX3d
IgSfjQZSdxwOOTcd0QR+v/fP+mI+1v02rGMoYGHT0fVIVZmIoSSMSSoW3XFoGZtZ
cC7hHWhn/xuTeneoi7ygwGgpgf5dqM9hKkt6ndN3kL+hCyAOjzWeqkrJ1KIUtOAK
G2LbFXGC9SQPeDYxTLgmYLHlMU6GH0shFuh/55QREItvnVIdqE6O2uuaUfr2O6FP
6ulLx8MauOBFacrcTAhxu0Wv49tZzy+NgEIAXbaEeJnuLiRPug7IiG+V8BJpVgos
apFHtaI8dmXLqqyvkjsPw/aBGB+xllVGuBuszhvx2Z4aT4YA5FhzsFvadRm4xQ1q
ME4gVdcHlftECaV555MEVnrUlGCjIEkuamR20QfmHqwo+dIeyjk5Oq6aFvByUnZt
MCDAQ2yT0+i2P+xtuxhc1dNMDZrmiGHd/sJ6HogS0o3EVcHNOEIznYM5Z9U3m6ck
jWXKT44JNkkyfnF+Vpdt3vkpGl9a9IN0EdGy1qaxTLUbK8jXWPFK7F//WUae8g9f
5A2BsDOdLJeRZWELqV7NmT5wVeUv81JsGvRVxe1/bAE+pJ/CXQO8MYJr3tjQYCdw
3RefAt4FkCpsr/S11SflxSjJIcnayFrotF3LiexhWBI8fyOn1VACqs5qe/c0biNG
SSiv+k6Fyw+MG5fdyfadtsMZz69/grGJjKAEFDAs/SFCqfT2VljSJq4kxgRY+bNg
3hY27BXPcDXz6QOaEa2iwTWG5dFtXGyA1VozTcoLm9mgwOeMQi9pyml5clB4d8NF
mefFpTIOHaF30uLBoBbTSw2xr78FWg7KidxfuhwBF3ABqnnOJlNG2Ldob11ncTtk
mTyxKKFlbNzWJ15v0Yg90qqObcJRV81zzaRcmp+cqC/RRtA8mU1CItlLTW0g+nzB
1CROLFYYvTQy8X4NYS8wqFM21OOz6zTU/sCIIxFHk9DtOdeWSGscjYazrxGI5g/q
WAEJB+eZ/7h9zFOrT0+jc3++i8a9Z3eITF7PmuXgn3a414Ag6Ww9uHJ1sLT88yAy
iKeGEVCIj84isGxX8/QR2k/4LlDaFfK4+XUkD/2EI0x08tjthQnj/+zMeAPGsfnT
sBrDy7VMtw6CpHUou4/aZJUWF6IoYbbeakMlJ8MCZCtV7zFtIZBPUi+J8k7udgKj
ur+d/9MxR68wgd8XVsF9HICUa7QK2sHHzJ6M4xfKuE2aWTyRzr9q6ix2/RBlenD3
EB42SnNpD6Q56GeO+E55MTNtTJ/F+S4bRvp9IXFxm9/WeZb5UxHTsRZTMR9WaQz7
3E8KRZyn4K4RDbgxajtjzak7ivwgUVgglGIdzKCG2vGHXSzgbAi8iJ8JRAeCdFwG
Iu/9hmhm7J4L8MtTeYYXXIURQmas4TLB0Imu8DLNeqSkkqESEIxr+uRsx3U3+WrD
Uz2lSWxnceR4bqfvVz1reJ/PPRAT4Csj/elftDZmFnYVW3/G6ugm05txAy4D7kA9
oQF3jTRdNxPpTXhOg63m9pyXfN8DPfNyyqhusivcCoGulfjgKxRiVw8a1vONUyum
hAM7up2Rp7ZnhQ/P8usnsGcC6toaWzj+h8RBeWLs8K12ZoWmSpH3Pq4WYZb5XAiA
MZn95SYenbaRap7NWumgNyCE/qDryvax+z6IXusjB7hAubt5JZeRqzeCUJW+MvnM
C6YG406SnDI4t99rHcnMWwTx6qvee0V4hcgTy4L375zq/ex3umafBafePBIbJyPt
wfRgvWG71sF0pZsSqBMG92z03rvOtCzPu5dcKnusd2ocW4pr6nNCTo9hRoB39VKo
v9bzsvk7PDIrvp3m8uGdfDepxDSyMxtQehouWu0h1Jvil8xt9MBuaPDIZo0QV5C+
Xx1bPzcMOzlabUQZEogVaXz5qi8p/XlX3QnMvKbF44qvka+JHSBZdbjxPgMT1/mg
Kg2n5PFoQNIs0TJtyLSEZlfcl5CLrYO8hZ/d4we5Vqfj/rFokmhd2Ov2WpYI8ePY
8NMJEiVyYW80Q/O4CoslhV/S4/pq6J3otKeeNfWxcnDf/zcP4itfxCvuVwe2w+sx
CFLYY0I0mYFFGdTRVLbXgwD0Gir982DgUk2RHVuoZpTKQY+49kYeTRy5Vz9xCgkr
s/f2OwXFITIg0H6kn/FZSwBfGEyt62EuA0FfG2jAb8bOdn5FoF8MvVUo4t9pVfK9
sxBheDSmHCnMomA3qp9PM0UR9+fbdwNeP3fj9z+4xKdQm8U3MN69Q204l4BbDYfY
J7BqvEHcCBEXmVzAUD4fzjoiBpqJ5u6kQsMIMjkwwiZsCwmyG8Nzp8K1XUjdgAfh
TKqFgpXXGHNmhxoEvnEQG7obDrtZUH5tz2lqzh2Hg8B/9Lm0Mvb9r96oQoyqGk1V
uz5MzHDqbzLPPY/pgBWS96KJPbJdts/YKIqybZV2mUi9f3l6RhH8MVS9usaw11tv
JiwYmbzheH88waclNFO7JNiAeV/y4ea0yaNHkleTZ2EG3LAyq5J8QH9DxhzXYMYx
KgODkxWVYTLqhzFZtcsYdSgqBOM9uBVGO1Ai549oJAF8B/2tBdSry31hZ2+DqRLK
+jZw6bG4s2SN0Oa3ecq+W16+nsdj8T+VILOcvUsg5oscpVVKXxAftZt6fJj0JXjx
KfS3Dz4mYdlLaB721IRb5Af4PdPFY+4cdFCcj1gB+AndeVmfE9klqh4zMofcuQmr
b1NvfbyW2pthbZTGktKujwFhNOgDHGs84nNsBhXgof4CNaTGPUyotmq2XuQPd+Op
6ispPMteyPoFjOZ+PfDmvD/rIPiO1Xasm/LiJQRMfYsgXBiZmAG7R/xXQhjAhHma
sl6EPx6six5s4Qd35NIk7jZMeBHhHux8wV6g6XN/5oV/A/n/wrecMvSocwxlk2+T
iQ4gm8MV7FV1R/EZuVjgCm76obye3jT5vJVJanoztB8HpPZJK8LpGDZteqGAnYYm
qWabG+EuGdx3klEWkQ5jEc8uhvBkb/0ga4eKZ9A8l25Wz7hG5T5kS6vbynY8dXkU
CkvzmO+TAr/Lbk40IZEfseUpX1+Gy2T8V3jtPCLEzgFFqxZ3oPn5RFkav69E3SIx
tmHxMqjrL3xKun+QCdo73cBqusQsZYx/T9utdsYDT5ytocyhxWENjCuCjrdjEJTx
+GwCtKprOJxdXvJmC+3G3ZCvc8/wl5taODCUBpuvo0LDyXW4V1T8OeQhaBctexdu
jwsa3/UaYynHc+dDI5JcFpQuTdkjhnrYfHTUL3OVb66Bvi5uVrlAbFtqVNfJMbVe
yNcYmv4OwTmyIm3IoelGZiMxvYGEcPxl3GVYaCGyqX//AoLUxrVYBIclQa7+n9iL
QuPEw6rFJCVqPUbrMEZMAYSAQIJC+BbRLPMCve/5T2aTVwSJqKNb7XzUpQP5bSuj
H7JMbGp+OsdDInU2KbcFEz69nSGccIzEpq72rcBfuh6orMwrSlWhRGpByl1JiMd9
Gkn8LeoANeua36dBvdhiIwUBhMgXyjEJMAH+4qtPrELmTab7ttWhAd9W8kiaytSI
JfCHnE8G4E1gfHOxDgQ/1rJwpy/Hwg+rTXlkjnrtcYw2xG7J5MdWPaiR5jR+ow0j
zSkjbnfUrUPBAV3Ge/9M1HZUtnzcSblTeKwmbuHsEkCj+vONUDCPVgZiCX9uuRSb
34jHZzT54LfYHelXoyq0UyIa2/dumo/yAdrKSoDyglKztm9DkwGLQk4zgQz3Ys0p
AL9w/Avu0016kPCawNUr9MRZ6QS8zVJVphFuyMDfuZC/b+OaiZsKomd8kQm8gc5S
NvlKvoBTIEsUaeyLSzz6BywGou2gipxjp+y5JpspuLrD0bLpodAXp0DtAQNhbOsS
E55gd6sBJKR7IoQ1mWBRGyZYgsGJj/bXge7yvWXs9vDjA5c9iUASVF97l44zeupD
EQDWqUVBjmZR6nQOqDepEvz/vhzt77m+eh9H/QTaM5KVR+BsCWuvbELybtruBzDo
gjStFuNRB/hchrkPaTiuvCbDSmNIuq3khMoUbhON6IE/VApOt5+/alV+lGUsLoHj
o83wIFeoXtGhHmO9SaGgte04PCtjFlfOeYxm/CxIeFetcLx2QmniROt5IV10R2xj
dJljymROsbu4RhNy1A9ozxzmbbO3foTVmbcb/564XZV4o++5f8KYBwPQDJtwYhD9
56NHRScilv3n+P8DE60mb+1spuMA6lWUtlF0H7dDUrgXqZin/m2WOARyI2KGgOXh
nfjNs5snliJmYxfejua4tyeCw2BO0I2yh0ul72l5D5Kec0ahmdGWbkehmNdSQUL7
/wCZTsQnnGuDN92cUN3bthbUJi9laxkXBdsrLDErTWTUme17Y+0HLnzNFZIvQdEX
nwWw86nA4kNrramchWcG5bgT1cJoi+iZvz5apzqCSI7D2Tnz10vX5VPzKHd/Jypp
yQ20FGVnEhPRKX4ZH0pbYqy0iQ6Kh/o9KyW963ySmY4UO+5dgJ4SnItmQEZC4wkg
+uKUgKH/kylFevi2v6aKplw8ghQD9TWBiU9Lh0h/RrKO7npStVsWpOlCERF0BLDm
GKGHjviVfnagCCnJ8BqeKdpsVDXr1x/6WEUXAsrdyh/qZr93Awk8AUu38mqLqsxN
AcrdXSQSEvIDFWLsbya8T5BXYV5I4UmWDxXqOAzgRB6KCnWbgzUWJYI9uns/49yM
g+v3511HmbiCZE/Q7oRv8I9pP0EQufGijob6M2Hv1DA9PkhK0l/kHib4HsGOAY5Q
n+WW+IsQDblRhj8cLhy3t13eEWNXtCavoziZUQOMEt0uqUf1HtD7+ToFhzg/2TZe
mAueW+HU4zMTTYFSdhLCPKjtd728AVf7wR0ZRCGPFFFBjGXzCj5IqyjTJK6nYUjI
SUWeNmMOZ6LhArIaJzSIod8QUBF5C9qo/1BCsZVqLUePxeRPWhjZub1GKMbsV35s
lfMi6Ltt4PgzyqwS/5xGfNap1lJtG1xI01BrqpYhjkwuvBVd5iCSwTEtINhxPcX+
WM2qTBc0cuh63yZyHfwK3LR67zxTFJqyf5XTWfV5Y6l31OZJpvZaxvnWt9hYHCew
ZeorWxsdjMVd1P6paATMy0pvbyNv4Uki/3qXMC48Akb1YaeeZvTw9kT9vPBh0u7U
qc/0ebPfOUnusvCq/T1oPiEuCF0p0rjjdOP4sAnrj4bdlD+G+3cP9uN4FvGyNx1/
ge2Lx52JaqTh4FbLN1y1UGIRJcTIOoel7vJi/JetnfJ84VM9XKhqxrRKJ8M+WQS5
TRShQQvCfxFjlUNxpj+AZpdmDfL/yHkC4mQYH3wnWTKM2OujXeZnsWVsD38u5J1Q
ZMJmFvz+n/7tle3/VbPD4z0pbZHigCL0MYJa+mem9Q0YH6dch2TGIRqtXAMNoLP0
aSmLRImIhbZ0Utz6rwtYEwMk1tzUJxll8iUP2nyZrAvXgj/9vkFzXKejs1xYCYKR
iESoKqWRo++MwI5vczeafq0Vz9W5Kz2HP/BUYk16pt6DbpHT9PBk6QmXJSIDyoVD
gVGFcPdlSokf0gzWmNu8icMh/hKws/tOWyXdfoI0PJHA6cJQSTn8ewsy0W8z98SE
GRkqJENqjjLOYpyhdOgGwmDwhDyOmtFJpOxf95ryzZALhBHQREJJTHb4A3yGFoCO
UYCYR0hpUDlkBnpU8JNeP4UKNRRyVw8Kea8O5wkbtJhEeimWPQcRpSVU/lBYRfH4
m3N3dgwI3ftqmJWFQCrWmq/Y+w/tB8HpgfgCHWbGKN0kIXzbObtq33z+XN8OC0RG
9LyZ8spYhBIS7hfYjpIG0FIO01XnQyR8npZJyIL0QJejf9M+n//zpeI7Y3/99FCr
lP4raiiNOcMmyFUzuWqnrf6wSqo42JcAEuld6omIAqwX5eAKTZZQzdmfabxXpOlt
nw8OhC/NYGkgoVR/SsYtmt003ujPOtPvs7tScbTs9QXtNByEznShk+vOh9rPZxYk
kLyOkLD8RLTiB+KHYB8pQjvU6lAK0LWAYe05mlH5NXXkmtkE9RR2k+WCeE5QJVoO
FknPme9q6ZeWbS83iRV8BJ8YcVfqyoTC4T9+a7gjsAZRCMB7G0O0YJWMifnEOE9+
wT6EjjqSTBRkdYuiPfMweDzspU31j/Db4Z1VXAywTrosvnYSOCtpkzLl0BXpKshz
r5bNT0Y+55zkE9TS5c3wjV5riMUCXGWSzP/o6mkU0mchB/zyt0YUWbrE94Verfir
s8fNhwrka4wgF9eENAjBzxrU8UZWPRCmHYkBgxQCWi1i2PTC02RUKR1Qx+8Mz+1V
67Urhc9iFDJVsoV2opmREdWlOBi/rk4bcTm51nUrmROO5GEZxclXA9F3nDDEwKux
OzkksYQuq20ov0SP9qyxZhRvlmu3mu+P1rlRbHDX3VqnoyY8UJC8Z9QmiIgV7ue3
2fE1MdapbsHWiJ64vh7crRH8gF9WdAbiL06WwNJc009GUXKLqu/28jWDi5iUBPue
mLIO+hBZ9coBcb8J4c8V3jB2z/xWtqX3g0Y0D/4VNzmLRdgAvUj4u5NcjBohXk+q
o0TX5uQiTjvvQSAVi0D1eQTw+AqprUDhbpdxh+Wc404ZmczLqBA5WzSomKG+BqsQ
lpAA077JvIRyj72lNGgGfXpXzkJauyRmRr/OqIkqxMHgjDEOSjZQEacbwL36nRTY
okumbQetLSBC02LapcaQB2mnzC1rxaLVNYjfZrObggFnC//9ahNsS1KVAmPbRGh0
ysmeWJXlCKcb5YLZnNcMnUm4hc0zPNs/PLs7VOYuFdT+RsAObTc8JENfmiQu0zI4
G5bz4uU+2gdMOp7rp1w8QOxDz03JbeCKIGBgt6srNI09ZPgfGknW9SpCaLmqLar4
XT0afU+1QQfHb5dU4DhbR8IOdvatkrIrZoLle6dckqtoxPF3t4dxN6cEq2b86Aoy
PuEdqMVNsDQru3EG4UZWFfMYrH8oeV6ny1bs+eo9N22fMxWG1TKPheq0867Ll+Wk
gHdctczW9/vu0Vu2IfpuvHZUxkv016HGx+xBAab6Nobl0hFldVb8mJ+kIOTNpxFg
RlbQir6qj2OYe+wo2TFslebBK7cdHE1jM/Litj6/MZj3ftFg+yWCThK/sVXZS2tA
IJW+PT3kC9gVTiAVDHWxrTJluwJYpC/Zlarzlmy0HZqmPTNATj/BZHbhnrCp+y2d
dO1+UV3j8HU0IzTa5e0ZiWhcY45WyLUddPYnxCkn/KOz29D05zHc1VaH0xfl5e/Z
2hJ/FGoNkUOYWHHnouHOcvf9+LgGMaA2WryLMKeuw0ZZO7RFKi+zRyQldJl5L5qZ
LAEWvWCdDLEflMJOFkNiqk5uZHrBpcYBjwB2Hku0/v9DFZL2UisuCoy/VrevTwzQ
kEh6lfjP1TMbxKKDVgJhfGI/X02Uhkl3YRogLLH/bUXK9f0AllFk/6MLtbscGyUn
EsBKcf+VpMBfNSHr51+zXSk4ASIq/zMDSDfjccYvvYeVxwvflCjdcTK41c1yban6
653XMn80z+93MM0Rx9gjhQG+qupeJsbCU6dOKC3nLdE09bE0KyWQyJdtte13Dfgr
OULnO00fRBnt4DEwvqIyWVW2MzUz37f0QqQJxH6i57TqviM0CGkKvOkJrkzl6dcg
rMxd1OH7Te6SnJXTgs3Ir1ZBYHJqEZWmflOjw8zVCfk2O91TVr1+sZsO6mSGNdQ5
/QHZy2NC7x8l3K8aXZ06IYaJB8d0EjATV4o+3DgSLGAhMsVnBidv9+w2Y/A7gowt
NmRLSqw+sFwtwZACHnP0vT0rOIzCjn7FXiV0Nv03Pgj+sW+25honKUg4jsa9igsv
vAbdSMWc8E/wNcR9Ni/3jMojYy22Spx9HWk2tZwbiMgSfmw4njG1mPFdR7iSe0CD
78hi7uZviluw5eOuW6LnWWgr7hxS1KNi94DL6Wj2jZUROSDEXcoAX5N9M69XgBZy
kfHJofrHvkQQtwGmuajwLLJGkgyVh5DW8GDOjq0NfqKWI4XFoqf3Bc92cyPmDr8I
KhnZc4TRsLjLeAJlFYYPFt0recSPY4QslMUfhQLWOvBPOWR+gcJXnhg+RaOU03EX
5Jc8LJC9zAxiSnKgICqBsmSVmkNjH/aJaULJMGdd0agbh3PV5EfG4LjtdddWEjgw
Ee9G6e22asWqhbxnTv9RBwATDlPjW8bwEY1NbGtvRyHtpGylGXGDOJkarGO9nEbs
YaUjEcGdOYIC04MtlHIXkm+dDprqNOdvwvfYPMGHsoUPvsAAMOXRrVyjs9DOO3xW
ue3XXd9263IzhUBaXw9KP1vE0oHh+Vc3GOdTIC6UU7JBJlUATRiwYbOgjhT0f0dS
PsyaZmWkOa8uWoyuSthIFzHzYAxl4ahqyF8Pe56KXGLeL0Ye0YcZOEfuuaqGSC+F
dJRF64IkTJ0pzxtwNuuyPauh0RFK3KhW2gEmo7hT5E34aqM0cAhUnoP/vslW1ILI
h8pXzrH4y7GlR+JnVXCcJCTp5tiL+nppidVNsQc0sYPCZJ6LWTsgRrM8pGV5cgLY
s/ruB1OLuxPEXEA7HgTbhhhS/71XTRs/B8HxKRdcZnm3Tvrowg+0OSJm7GEr2gBC
/n2oyPWcSWyLQiMkjSofQuafA9h0lDA25KbCuvo7D1ONbqG/E0peJmECmjJeXvYV
ugKyaMpqvEswT4gJei3AV+mNyiXrNWGnq4v0iw5FX3Z/krx6I+eEmzGZYnYNrgQa
1+3Osy9LIML3m+AI7NnLh4rwY6IKpU4FwnBezR9bY+ega7J/L6b2B4A7C94aJEGr
TGEh487Sc2Q5neGPhtoFy/M4Uh/pyeoJfCvKgziC3OtbAhag4RsSJfTHt7dbW2re
Bs4rcY8wtvOnsgBOLAgbwj4vm1W2qD2cTvfy8geBqK31wOTZXx3eSV7taNDAuHfI
LVmBOWZETpK/OzWRzbyKRl4gy3iRxf0J87C2vciruXj849ycXHnrabWR13Vq577W
nirvag/y+JjTOhRe5r9lHrfAoMlc0zYiAb4DnBn9I75pS/ysGDiLOaMgGQkLVJXe
aFw7e32DnYnjKQ3lx294OonSb/7EdtL+fjDElDHN858kuTXcyCUfV2bm2uR2hYs4
oQJV6HVFtne9nJO+lJFVj7IwQZNF4I7NXZGiqQFJ12wk4hHXw4Wn/B6qrBseif2l
0A7zxVwBKrr79DrLe3dMBprMUYe/+po6qGCvXvvnBL7yfkQFpTV+xMe551DIPNdD
4ChWkYGhKJWexf8eDxIFiAuvSYVDEHBG0JcgWHJlwtxD85wxZvn5DDYEeju2+yi5
qgSsPkJsuLB6r9mFp5ecZUES6pcOWV+tQBVUcxRYQrOxjuIYq2Rsmmo13/HOlph1
TVY48Tv1ZTyT31FvIv0U7WTQd6K7N08FBcVYGPnA/2SycH/LcieCtMRkQI214dup
AIp6MH3zb4GJxmUWSynXdmDpgFzXVy7B38tw00dKJ5jVN9CffciijMy+k1G+Viqc
uoiWi15u8jnTmvIEkI+5nun2dTXAux0olias+GluY3zEBWm2wVqe/ZhJDUA950rU
H2tEINjMa2tbvnglVbQ1FaLI3jbR4At8F325m33jNXwUCuYPKaHlMSTMj+9YnvjJ
1oF2EYHh8p3fthdGr6wxE7ccJA2Atte/J5Hj312ti0PV6gkZ/iNrRb4ZXujs5zXx
JvC1xpaKWcPw9+2zQ7qF2iEAtj8yfj8EHj2h1L7QdB4DX2fEBfTXxNH+UnCrUii5
UdeVXlOaPROdblMeNy1eZwleaTz6+QMjD+6sUpNziy6wVDniPTyVXcbNhYHSuLM0
ONiw8GWjt+aNNuPpItx+FuvpQ3kyEqqOFwk/BTigdg8RhcHwrlYEUjIcDB1qaiYj
N4+H7yz63/6Vl2UNl8dc3TmV3JcDPDwnGIQIT4p/y8VUdrZFXXMKS8aaua4Cd6j1
SBbxrdPb3hjfJpv2vN2ZQ45/LI5TjsPF7NHPcNE3GRCgTw/LroNg/pp03wgmYoGy
38QIdJEIYgmauXv/af8gcvtMYVx42NKTCNzEGbuzgB7dgds0K+mw/u30hkmMAZ/P
s/0WBUtr/5/ShkQvwUefqmn5VVxJlrW6tUA41yr/1MFUAQ5XiGkMEYzsJA60pVC3
iW5lHS3qJkZf4BPGawdTnJ6hPY8qhZ6AddkzfdySiX2H70FwDw7K9IwbEP3m0qO8
zXJy52zD+qENf/mCjOc6N+vmlD36h93U7kpCmzSWxnnRZBzfRcR1kX7YJfChxzkp
loOFvlLSvMqGYysLCDYxwmldbKEmcNc1L1aoTWXgl4zex+YDceIgU2em0awu4B33
VzbXXR39KCNSBfN+P+93oS8uNJgvTDIMH8ced0YUc/we5bDN20R4OIyzHXN12tUA
yDepStudJ7fubjQ3hbszNK8ylyG64S8iwNfL4MgZpnVx8n9btYvEFQuoCDIsgb8m
nC2Rau0woRVi3HsTFPxlLzNkgjBhok0JmqtuUvjzgO+z+zrOj8TOJ28poLVt4D3w
SAsqrwUW8abqKocb0Onc7q+euQmA1nFjKBu0v4A1VC8v5j71UPjqx+B/bpngdmjQ
zrWa8lIXVx48hfQW4HoLkEgzyB2MeqjKBlTNBCwrPt/hhPHsRTixJH99fsuIII0B
ylC21+D+jH/HgpSXSYF2njQ66101vZphQSUbHpOgp4C826UJvx9y9NsfCwHFpZhZ
h7D6Xhr8MmKmauhaigRPiT2qGQGo9wP6nFeGqQabb8hobn+C0dOxjWKEW+3LfvoH
PUo8pYY1TYvrocYnjUsTbuIXbct1BCuwd8WHOnsYvTi9m8AKiLzNkh/JZXrYuGb6
9o33YIL+nIhdf7Otfj6iAPwMu2tWjzA8lRorOkjYLt77VS925HVLmcB/EEvP/nvF
JsTeEqyb3n00OblkSZpZZcI/NJ3i45Z9azodS1opjpYs6lPKmI9QBQvBjY/KGNNo
sOKAaP4hrOj8fle6g7D2x++sGmRv4BWW831XMpzQIctUeUPnE7HijiuWgn52fhNB
a/sir4q0WI4g9QIqSmoW6LPc1Yv9CJ7+SWJuaQEJ4/8vm34/6pQOWvBZRvn9/CAd
4z7pFLfVBaNTMtbIKbqnyosRdAUNqGnbGZ5ZpJuQe/Fxc9vge5DhmTH3SIuTBYz3
VXBlF6v+p1u0ozzLdrHfpwIBYXKDuj9h2M5FtHddmPIrKrMg5TkAUY0baa0yowsX
ip+Ch0kQVrsnEF47vvTzdoKmalqATKngEzIR08S5ZQbX+NvWBByh23m0Xlo3NRBa
0qTVe8lEIHjoXQAuJxYVO8iBwas3RWPU1HrbVJjgoeCk4g8BSg63xbtrG8Uowqix
FF34HneHlQlcX8it5doEqSyNfNZiQD3rHxC7jggm8YYrvvBam+SSm71seTwShVgW
Ptv/4AUPfxJBPNvr7yn8r6GF5ZvcvGMj2CS2vM7D9uD6uAfMTM+J5AUsSpDw9KQJ
UUhoXUe9qk+NYGmtEMYIei8qLpxbN42BMRo1/m5A1ISiAMR3Rvd5iKiyhIc1Am3a
0dSal2tTJJdl40DeMFBr01MTMk0TWqyMD3dZgaRh3JLoxpFfBY1zNgchHnp8BDV9
AtpmxFem5GaGIcvGZFQITIVPZo6P5X7/3aZatsQ1GDGiPStnwEF9gFL12K/IvQ1Z
i5osCZF7eTmMC//w56xlqaLEqsFeFFLVbqvGHIt+qfOTUud+zaCHKRqHVEzKkLRR
/SiGffeciPOQDG6GgtlT+Q+A2VUrZtkQ734QWyzcsgVYg+NqkSxLY/bsoVKqvNwu
Wvr9sQGTuGS/qbBYvNLJli59IVSRodKRWpYkm933gPexwPbI8tnzKVrkMxGinzn+
+5YuSI33EMWu5QTMAWJsu4adpiKD6oAEOgpWxQhtEVh7J/dueHx/J5t8/4KkdFB+
SN8hPnGzq5qT5jgN2L+dojhQ0/ocoxo/p34AWeQTYIUg7RY8/zU3fODpTeSX4JM3
4I3XnGIboAEIxONt7oqZ3PoWPCjpUDSuxdU3el9FlS+TJZ61SAXcB3I+vNAJA1h2
rK43+xn2s+iXfWyrzmyWCxV8iefWj1y9sUr+crlj6nVLQRGy1dpriJkgSzhJpQdI
cgeWUcEJnG1AY5DPPtzW9x316pzB/9u11F4DWEFSSb+YtzeYe0wLrs43qERZPfsV
QUvfgwfznifbgGu3P5qTCJ0OarmbOU/Tn2mBkciO5FvOCn58Moz309a2P9RH7vsq
LZYXXv5lgVRLiKH3R/65D76W+PBMzop8RhekhdDtzbCN79hA04wucMX9zcOgeV7D
ztHvjHJn6xZJDXhS2vjPYlq6S9qjjPOM/r011jr/R9P2HHDAIppyKwt2+l/UNO0P
+UOIgVgylcrO1ltELcl2w42oYav3ygdZLv/cCzK561z+71+6/B0BUpHKX2nKWAmL
sUXG61BHuC518g/vFEX632QI8EKtQmRYfQOVVK568me/w+Evcosao6sdSQCfDfMD
gWisYV3HH2fgrGLubUrLB3Sfep26Ty5mNQ9SMmLRed1yh0q8YN5EblJdinMIDyZj
i8hl2Ft73u5NoWx9Wz8HI++lDODPI1CnIBPZB5dxAJmijrED4b+KXyX3KZTHOtko
aND578LXdWJfXVdFx944w8qH41s7FymoeZP+cmN3+xBtyiKQiUASp4kdJDNb2O6L
N/VA65CHlLkJ+4A6KFcS5zS7vFjUtn8E+/rXPd6+jFQXVbKIZ8ukFL8ZRtGJ9XoV
4Z3ZOj/N/m9aP0g856idUfORHAykPXG+wVcGNy21+X1d1g+TrrMa2qGnOTp1DetW
K/fdoDhJNFF7ScM6rBOPKcyfB6bF8UJr0Ve97kcriJLYaWnGF4ZZRv++mOcZJzzm
aEf32KB+5D0HYmfv2IQhF0dAGyAUiB0tfWb1ZIxiTB1fYgb8hmIndS2wIfAJSock
e6V4WQeOcU+Dj13mZrvHQ9qd3k2irQTN34ZyFBIMuFuqYcxnsEknN44reVYq0gSZ
IV1ZaijvrQuTsyM1i6eRox9M6le67Aug2QgUey47o0DJPFvBPGx8tq7nwB6YxYXB
t8q4XFkhW6FkgXcURUxeao8eFj4cXEg8ZxNud5AXzN0v+o8JxHLWyu2KeGmFlhct
WJ9gfmTGyQRzcSqtdI/OsF4NDuUlnJ9oVh62VCioYlkH1VWKfrLFCk54EiBOCab+
RW6bKD16UuJa01FQtGDi9knC/+Ncl+brYu8/ch+BsKWa7gNj9tDJLgRBVJFOQTVH
9MSKVmp3BXM0TDWXhuj+pEbOlcRWOKsWu27aiFdwiz0MAo/S4raUeOtWAh+6aX35
1AJhftOClygyYW8g1P33KExoA7/Wez/rwDsCBHFbuYh2ZH1uvbtyj7hUHaa2rOAL
sFThssUWb2vCs8IaKnJVbOLC6QQPn0FdbK29caqTppyXLPlivNmT9THHsN3yFYXW
bNgaq3B2gBmpafMxly2Z5YuKU+jpe10lp4jabt4mZBXUA6uJy/HhkO6QEgtsl6z7
OLz4VLXXj8MxKXlK4i3Voobe+R3GrDekdlLi5DWlNo+L3+n8CzThe2l8oMRBzT8i
+wvh0wHziCGW4YADVIPkoq2r6D4huqogl54kuKEsZuLYX8v/o5vrFUPOmXyC4k25
LrwoDeJGq0FL7RgE+GR0XNZOvWex3tyaQKRA9/pximRfVm1bQCZkhZrmC7/TPR8S
x8CKx/D8EfbVeu7m0gjCoTYLkGzjRNGSVkhOaW8eMSGoM/3tg/XWoTmmB29V0ws8
2210ouYB1WBoTpNSmA2yVVGudua/iSZfKWj23m1kCm+vJCYyuIWjgeNlxFYIjwCc
3QrfIMLNZZfEID5TkdB6rV19h2K5eZyDGYEVzzIGIlui8zxZ0nPoheaHKKBaQPD3
SMYFgMTiYV0ZTN1nuu0hdDYy4hgdebS17wpVCwxprO5I8jedaBK5MuE/kwCxqz2u
o4f6Olp3PkSGJTkzGCd7huj2zjr1Xrp1gl7jK60jRcbFkai2g/PomEk15XIrYB/8
yom4e7H36lbjUQp1k59jfpkACRCmhjfB73I1oUWFtRRlSWVrQXG3uhInosEQfPgm
MTwrFl2JHbXoih4i4lAV6W7hhikkXGyarhuRdk5dDzQNhZHkvAO2qTy7YbAVb9FV
t8czPmFJ9UQdPa1Zf3rI/O+AhSdohYKK2rs/SfwvoufEhfGTC9hivHGyHI52cP1S
WE55IxSHjAm2/gnr5XbZEZqgJUFtW0OhzInhPh3mn0PdJbGebKU1nOi8KZdOMGV0
zr2ssfstl0SuEyvYPQmWqV5HPoRC4xpilgO+u57dAmf1UswjZ54M0zquaARBPXtk
oYx0g3mf9IIATj16YFbu5aYIhpEVfe48MngEpUFFe1MAio2jTjfiwpL725r+opxz
s8KaUIjsCnT+b+7xlqMmiGovxBTdFVIWvRLJak/JUHtq3B0kxffJpc4zptZiMZNg
Q3DQKRj7bsYPmsiC0LGgDJj2F7XwNFtqVUeonQsrV51K9H9jWCY6CZ3m+K3Ib9q1
hhC4n48uydaTdmSg5TGaJUi/ICcfHtwhGJMs7XCROqhCkGhlNGLeGzgiCpqY8X/Y
2yRMo8Khf9GowtwSOumzqRDk6VKvHKGQvx3Qdo2WrXYSxvXh6WihNyHvEjOp9UUo
rSVqbfljet8rmV+m8Rk6GvWsosmlDbjNnw/aj1FHpKSScAIBnN1quRIDaEwT1Uie
NLtsoVSqDXZ1snxO2YWOIyCM4tER8ZFTmFh/ecDebQx+5c2ryARRrG+zBWu7c7fL
ovBC7ZQuogLAWDXBHr7CwqK7WAXwM5ptBTj1Ss9DlXPQyTzIvDUYXeYpynSC9Bnk
3VozOu3a9nLLgwrDvq9TwcdRj2S+0sUPzl70k2kStNuMAMnaZ9/nc3z9RlHi8xkx
+h8r7qiLkr8/mXxvv7GqGN54VMYbmKCNT/h/nYxlvvep0t+lK/TiBPjJ+SAg5Q16
XOlyypjzWBafS+pKpG0o+vxQmBV2LZTLJkjhrYdSbsBQKA0ajhoTW/LwtvaSM5MW
SKtffIeUMExeMt7id5O8LDJNzbUbvUI1JEpzap2kUdkNQZhbUX2/FJR3197qfNXF
DmwfKUe2lxoZgWiJM9f9OyAl/UL29g5rtImAtr4Ckd8QUKx4jL3v/eR4/UnV/YvB
BeKQA/3UdTJeGZb6ioH7kHZ4A/VgOcmQ/a5c1e6nVU8e8TBdDn5Q16qMb/POP2VY
ky1o1TUjGmtzHrAtY2NEeuPn4ckLD/dQWfzypdvmoj3PLv5nKU0h+vCXj0GXqkKj
a8IZ2zJZ4HwZ3Fd3vxLpsiI0GOzpQs1rEr6Er0taGBEDpXe79lgY9DEAWfMn4atZ
f/uGfy1EnsQ9TLnABmIpzqQeDHFErrhU1wMQR4jWuDWLOw4Fz8zKOg48deU2RTxK
6O450vyCmcL5QG7M9Wb0gfmSjmdUFxd47eoXh22Np5WYU3pMJUyn+6QXYqHsefTD
pwaQ1EPkINU/p00XzmaS4zaX1n+AaCrgFWQlv3IyizFq/t54I6Cafh/RFjCs/+Ll
mmnJXMBw4MqM5nhyWcr9trFTMeN1XYLokmARBVdnNVnOkec41u88dsGZwAHlW2SD
nq6hh420m5plIBRPTpSvenjmqTIkA6pEiCRw8dIRi6h3VVfy28+C177FG1NNcy/r
RKBeErK3I/smEwm46C1zVqAMAKx1lyzQ82EwgngAIVI7W+OTN40mT7xyI9NHulSE
sBSGdADeiKgMtcr0KzbjEXYpnGmKBZtaJ7wJ8cHQbrBpm9NQ82PrKo42wpmoQaDw
/jjjbrzStEdnFddpB7nzw+CysJvpLMHF1egyWdC4wKzoa1rDNWgTV6mX6GWulzHh
Tpt17JDX5otxn5fN+CfnxUQllTPjaWK5XCZnE8Cu1bEVIvyziZJCx7CknwfxEBuQ
FmEUPnzoYnPkE2KM9hvaiV7UVkHnb5TyyfkZNIkhUdZj3FbqyGmoEvraLjPBtRE5
hNG1guSTz2bDDApGPamSZnAaxfg7xr1KF0I1yCVdDsV4K11TQCtksSl3jnHAeMhE
t8nnPF5juqK9F60D28ZNtgBn9jFNYKWaKcEUPQ1AFaDNa25sdGf2SGpH6wGsClmC
mptqF7HnjN8YrOicZixgB+FsDfllf48jxRKvA69CjNWYZ8rnW5z8Toshl+MuJXNZ
YJ5htIjKvYo8kgHDT3LKNnFY4peAmm7wFHjV5WNi6CMgQqJQ+OtCn1svx7Gce/d8
f4xTcFkebAgpnKRowlLcAP1bRqHLj+2QePKcYZAGDj3Lc9gee3A9pZE+hFGa1eoM
lmCBUO2TzPpjFXS7kdPn6EpnQBn8yptD69pDLV6RUCwDi/ls/IgE3rhxb9VMH6Yz
sIhsuIs25sYu0mUj85eif3MtER/f9dEv/ACsiwvsOsoaW4p27HwxU6SiOnXeGN1+
TlG7MLQ/8ceP0huV4lVyiPiCqs5++I0xsOQMfgOUdyQB6fqkBok7ZKjmx1HMCB0E
655YFf40FbFzC3AVEPO5x+myM0Q6mSH8kTni/ZFEESAC4BOtVtvMRtcRHY2e5r6T
2MWanb+IIKG/PpT5+1jav9zjISYrGkdvFTvpJRr2NWdcdU6X3N09exEeZKbWEeyJ
iS/0JpJb4o8o3VTVjgdquckiO9YnVKgBehKma2C7RgLvx9DTJzI1umzbBM8UNa2E
vyPsDjxFkSUIZTVGz5FRZGY4y0APZuLX+DbO/YqjqeCMhhgGiWi0BVx4PBHYRgr4
ihw1Hhv9b31WwP7ZxGSNzwvgPVgdiW62WjxHAzbWJd9j/vt8sslr0A/+FBoYYVbH
uqhfz/7ueocT+FFeitVyl4o9G9pKVdadq2tJgv5Qrsy3uFJVxsgiExTgih/omCCF
FlCPMIIFmqDOuzjb2zWxf7DQBjpLZAP7TlmawwWPiOK/aYTg0fdvhUmWp2qDODqa
NDVXkac0lgF3Fv/DVFy5dUQUOvlUrhFbZmoMK3r79sHCsS31kVbx5dKrJ07Pbhrp
1zUtvJv1TRY7OLkT0et/VT4hI5ba1VF1qJOuUV6/TliI64FIYB8oeCK/0NJk8RPw
ZJAsw55glyiswazFAXsF4UwuO/tmEp5xv13SYmVHWjKMd66O8gteO32HRTeiJvhB
jHHIxjN/RvavEKbwAvhkWzcWKEWQbbV1q8ll1hVy+b6mvi53TygDjqEmKU6MmXzY
7TyKvdrJ1s1gA5AjL+N7n8cWcbPXeYR/xv+aznv3iqVGuwZR861TpiNfZp8TVG+C
CucLFCov/rqvabifyxkKdj6ILA1viHCOdIeakkkX5/s3n9ykbV+imSHTvllW21K7
YRu+BVkY+rx04HVuhw0FsGnGiJmd3CJV2F/S6KvfBMwlETvwcKgE3/k6pHViKN5x
ZwcBpcor8YannjNk1HN5ZhtgnwmUjocRQw5meouP6BgvrO2xO55KELPb8jANCP/R
S2i6RghnnT3DOpzgx6+HZu70NWXYP4vi+NWCZoRa2hR/Dk9MdHEvXMKXVM7w8nCy
9Dl0EEeGGfXTsiGg3Wua73qit7Dtz4PclV2mEpkHGBuyIE4M+5+LjtPVBwE8cWVc
A7nSwaX2yg8Wp+QASDckN2L463oajXWvt/QsGLQpA5PCnwKRz/QA0ntLL2UUIpvJ
gqVGdRfTmbWCMYwuLQ8EHbjG6e1JLils0GAibfOfgBzPvKux1TSeFvbtupaDk+Ch
eznwkMYHtrTBtwIzZrfMMtbKtL40aNZMg9fYWv+6+KN1Puht2Q/3C2B7tJKrI3lo
uX51lLnO4dNvxyZj6hTazipn1gfyd8p4hhULsUW8V2qcqJkbtxX2LGMXeCeLq2LA
z0lPkAWgMo21x+TqL/WfTpKiOSp/Us6yKhe1lOkCFl4S6o+BeE5Gi1/JvCDWAq28
0LxIyFpbzS12XuV52yd3NZe8bDeWzeCPdjt6+R5tXWCRkUV50hyngOX+YApopVQY
WwZsUfQjqXa6bTkXG8Us3xRPmf8QlQ4UXOue2PPhKmszae80lW1z9hebF5n57IUy
qQ4K+nF3yca7/2UoWGc8eNqmHG/tfVp61nHlywc4OVIoELaXfeQWzwFoGGhV6KaP
lSV58EaWZNAkkf7kU8kFaae62i/J6fBSaqc2ZbvnUjjFjR949wdeJ6jkItcbv67B
mCM/U6jU8uYcP+kdMx21OWHYkPCUrdzo5OiL4g+JHGvor2a3Jg4z+sYEZPr3tdsU
p0jN3UDErVjMzm9Bfvtu2B7pj9+Zelrfx5bUMCFN3viVbL2AggJ7E2ZN5LDMcKDW
VEiUuFgaaMZGE9thn2y7dAEeIz8t5p7qz165GoPxqcO98PaImg94EI+z1lJ892rm
wAQFyI0GK1cbfQgu6roX7QUXBhuZyNXVfnpYTIG4rQtDXltdNE51bcD29PA+BPH/
GVONm6AZACc52fo/DqkqwOSXTg4nnUt453wwBkbSpCy8ginX7E2rxRwvPVxJ+rKm
R7nMIdWfjWerjtdHLGVnXiX0HDx5dFGgrmawXgK0qYwbG1RlfyMWfjh3EF0pawIU
1lX2LCAnyCb2AbDTqlbLqkeRgw5E7ioK2dhxq7Y0vnU798Z1eO9evquYlgC7OiF7
M5qxs2GaOrAbTCjVCsXmn76wil3OoLiyJSdXV5jPkmjZ5qULzXoBXLOkc2qWdLy+
8bO54Fcoea0jUNlMwECUI8aCr61ajtGzLqiL4wls9Qy6OnFb6s8wLLXc+aRmqoFa
MTEmaPlTZiIBDctQPl3UzsRSzwTSjsapu7SsCqKnMLg82CypPf4nUOz63bTNL/L2
A3K6hhe+AFT+1Ycz1j6ur3HpzDlK570t2rlFXvfu/HtMAv402V1EHVjNEiHbeS7z
UYEULO87XAd8Su6WDK4IjKGGqI5yBNzYg+n3hl3tARPVVykXL6QQyQLORuhIvC1F
2G7lzCW59mSJ4GP+UzKdbqvOpSPHEriPD59lDiiGGEidO+0krqSjYETcWWA7ZXR+
25c2N5dDXwDXgT0u5HvC43+CWNiURs2lA7kp+7dosirETtZf35c/v3NlLwQ/xcpf
pfG9O7QBNImcdPCtZHWoJJPdG3vBtM7XhWDJemrT/E5TnmWi/1up4v3gplqEi9sD
p1ZczckOO23hHhtIdhPXeLp5G1+fQcZp86vTQlb2aSxGnWdIeTIEugIyEVK+3Dl0
a4rgjvUCa4VypCH9xany+QzWUfXf5xyXBa2B0ObI/Zo4l9dVSSkJc4UdzlTl1oPY
N+aw5TNM4eo71SAOKLEkUl5ymflbIaS8ezoYZ3A15y0G0pRpIhOFsbtf4b0FiGM0
PONwprm4I7xvtmBMgvuGsAbCAn85NZrsMN5vyIrGLj38iLMqAl7Y8kH13iplfRC9
8HQoducDrPNzpw648ZAmAYLdKH80mFJTDmauiaviOWFQ7k9wHC4aiOLlQiwMZLCb
Rt7nX99icu9aE+PMcHJQZb5l22Vt1zCVR6Di7RmdyaDNEcsQqjVNPIobnP5Qz9m8
TYO17gVAFJQqfvIimShF6MBm0VE1MKjZCXcIMUMymRxcg4e6N46V/7um+1Isaibw
effPWFKhAfbYEqTXVxA097ACov55LR37cQSRINaO/a0bzrDEOiVZ36htXjQgC/Av
ffI78bKaOF3Y6QqQjvy6yRYLPL/lBPSMKmHv7l7DfgbToku81UT2omCIWO1ZVVWN
jxePtijPTS9S7o80MOH4tMOoerzpAnBAnz8Ij9+zKijYiGestoJsPr0MXWOgb3RS
EEpwPutIc3zqGPirS2ekmLWjrbw/uEOuFS5nrnOInBEE97uMqMw2TERNb6CjS6q8
KSdCyt6+FjQshBwfeY31adLAOT8/mKOzkwp5VD6zL+95e3dtyoq8ZgzdNAQTN0zc
8HANbwXDXy7K7kPkOPj5+aM3v+GHFQxY30O3kZiE6p7R1MXMRQgajleYnV29os3h
+8fF9uMhjVz23b50slnreHF+TZyWooDRWcBP4VNmyb6oD+5iYsQ2qf2jytfDsALt
frgV8x+zSdTWEtKLg529UgE3LS3hY6JKTPlP+wfduRh8PBGsucfUR2JPG0H7cvhr
/OJUQq6umY4cZOPSUaZ5Mt7jc2V0sKPA75dyWQDOoNf7Lu3m+soo+VVfea6WFux5
b6u5a6NGZt+glNBSFFyWtmFCAkZLf5YoCxeYe/Syp5vIlfiUhVt9pd5oR/IAlHJb
ilkCY/Lbu/FjL0v5L2zxs+0fz9ZSeUQ4GC00y1i1H6Vo5KMxIDUj1JwKEcbf8HCx
A4s0Ibq5FMZU0heHvA/B7iCfNxD+1Db9xGm8+DDU+wL7SGvZYtf6q3H7y1T1cqmC
19gf79J4N7YbvmQyaxbOTZipcCPUVDwwayXYazWZ/eCAJ0DIwFiWZI9lywhEii5F
x05xPHkFYQ17RRXPDm5rvQBZ/NuUe78JlPu/PyCPIJg0fKnD4LCZE3Z5vLwpmcMC
qbypTNNTfNDp2ylFWFCq8PPN6NEzPe0yrQWbQOMJ3anvVik8BJZ0XiP5pW9Vkajc
XdPc5Ncois6KEIzzn8hWihrUYkTjHeOTVyofDWUv3FR88arGaGXW9aokrk94PJal
4bY1M+t3JgIE08KjBfG6sGIih+3vi7vQP5HJ+/lm59yI9Ulfok83QRDtH3JVGDA+
K0rbS9Rq+fgnJbYyA0fhaDGOpxp7houwjeneGHsxGX4St8eHsc7f0x+Q5c5+miWZ
hlCvkM8sVjscePQMckmhby6VOHe7xb+xjuzeuFsVYTDhFbv0v3ZVZaqMvB0gaBrY
7mBnQT8SXSDP44a88+2Yt34Cl26mw4/CqqBY67cYWPxK3hnKzY5fXPMhi19Nd/9X
E5Z1dmuZQNwndd5c0Nl1PCh3Ftkf02ff+T38+aw5ng6oVAmdS7Ti3dd1ZVktyOGE
O1pEYs2HVIHnFd/IzwU+y7FwlX7J0Y5NrOV4v5EGK0BWM/zxL6IRhFIRsGK7dqh7
MMvQAuBpelAFjvgCKV9sQhSIRJMOXRj2uTxsqfC1nRXGhx3+Piso9N0W99SUn+sf
iwOdhjQkw9n+d89BlqwanrgU8AVETrKOXVw+C//o7qXJr0Rr/gYFzglTzKKa87ll
+uYfTOLWHPfQL1jI63Slhu7Zj6o+gmRnbvn76LtrURHigB7cww8HEUmQpH1v7/Lj
K7CkaxS3eDqJcDMGMWyahqyEAzSmomJnzOR75T+WDYvTPPJNniiwSdc2ohfhCyD6
ilpng464zcM7Sv8peFgf+6OXJrkrKsC3UNQFPF7M89cUN4PBhGPQaSGCXcNGHYhb
fP/ROO83lXu2gVQ8d8Ml9LY4EsXFIEwF+l/Pcs8PAXMfJitoVuLrB54eXKSvrg8r
IEKbgfWLJr1KTwgTNhqqzZS22vBFVeXqER7lQD/DMf+Exrv0zrOAxA9Tpg8VzNqU
cPAoR6dGNLtglxYJvpimH/LDCPjximGhBwHp/nyEIKCgpFNGHqNhJkiG5WUiekxh
ZFZuLrmB6JT0ZXCYhVQbq8rErDUuV2aAueF6GpIR3dU4muLBCUaC3H6bwyZMP8K/
OpdLiY710C5gVmJZVmsCJdRRGDvKythUGbxPxRv5DpJVjWus3myvZyIgoHIudbFa
4Ryh8iAn2BFJJUzrRmPvoZneZ/eN2JrSwtIHKc1Fw/ToZe6FBynBVbx7HCnFa1VJ
G7KYwJy7T7GvvSK23UAxRZUDjVffdED6k4ELYPcmdmB1tcnncvi/jpwK0qsIWG9j
SOLl18+ixevyX2vUPO5Wb6rZ4whuDDSZ4l5GJCgOc5ZGmjQFJu7/syNv49uzbhpv
nD3shofnNbSGi1nvyKe/0lpzvkZ5dDfqU2Kwym02p4kCnGMEeigaDOPGmyfAVNBT
OSywRTXVIxWx9cNPybNPD4mh4yxnefZ4828/h0DBVPXU2MeILzxfcslMJPiHdykN
+E9h3x5nK4s2NWQPGsewcCt7HBTgaJ1h6rl4DsNMa6zcs6YXMhrEb2sQ/XNO5rqd
v+fxkHONpCYdzKEUztfduUDR0Y5l6sRBaYCsafCTIorxNlt5S8izKRPIVZL6GURH
fuF0lWaIXvw1ZPoMDAv4PQ92dvtYgPNe08GMwkKENRrcBSTxjudsk60aYVjn5MrE
6MWk0eApDmCfjWeJ2oXsYP6NzSxlCUZ3RX+twMt+75KEvfyrWpCnYjHxAoYxGB9K
hyny6Q5UaF/JE5pG+TwuaVfOvKdJEfHEThO08cFz1Cb/FfRwhVitbO0RGUozGmCJ
CXbgtSTGBaSoyD0GqyjA5U6fLrzKF8C3dlu5gD5ja9Bfq81yWBf5iI+aixvT+Pth
D/9FZh5QWxyFAWqWqKjTId3Vvx5aoeAEWTgB+rUPe6gZ4BIGPCxtfb4FWMoCAqc/
vO8dDxfnvZaoKCsu3lJbN7mBBdnRPbGQ4X38PDTGkwXniLqhtaHzh5gmNJpkBSfA
vC8z9T9m40EH34rOsPdAvTR6MjtNqLcnv+qd1iP+CzPFnPmqK5w6BpfiPFKYw3Lc
XAjGNMI4gxyhmLSMOTTwuYb5ECI2vP7t8HyLPZqkDB8uknDLtVVs8uGHUwhmHZrw
pNZuoorVN4rwitvetxg+9PPLHYxHpA28InSsJYNx05VcN77mridbfQdpT/X08zLd
/X0K4MA2QiADYNq59/waB62nTr1j2jF4W8pcEgzSGGBl7V+azXnu7YCkAegBaCMm
CfF1Jqu1+0u9nrt3VhR5LPlhu4SilSoXAqEJwsA4LFZ0Sbs3knfLpAe0DCyz/LLy
GFnDb/eK8rNlHt9V4gyZEHsmJST4NjGpAwZ1fWgGV8A0Tfq+442OI4trtw2KytLS
I3sbul1ZModRm68B+oazpR23Q6btroRgNvjOslhWFLFdm15KLCeVXdULSpX+UVD3
MJf9ijP+CWbLBg3+zsThJl4a1e8dgENW8IoYf01wLHiFYjeHtZwfuYzJN0vY5qaF
JiPTEto4ovEbnJuI2e3NTB5wVlgYdpyIS/mVLbC5YIpB5VW7tul3CPnjgcFaIHhE
lJEIPJCRYaNUXcau+zvlrivN925tqBwqB6UoF64HDjySFfBPdE9kEIFrVLXIXMs1
sseEZGaM0+EMI8FfYsVpYmyWdPgLQ3sSiJTZ+cKP0GY1oSmwN1MIVTnJOER1MCLs
ouSjb5NF5jqmqxVnHScePLQcxrii6iSkCdSMWsQFlnpe7I5Ut8D1MSRR7CZVWXJu
vegiYu1Mqn8T/Tcamvr/vcQnbM0BwLk7it57hIFgImazaEfJnUX/assfFB8ke3nh
1rYZLgiH+E/jDYV8EI6px/b/ztQ36w6+VEFbxmz7GWyk2bIG2eqbK4hOLASkVlvZ
NW9/q5jMMlbXKJvV9WCib4sdYQD0pvfe6iQoAe/8y9t70YW4LqCuQtB/Idu7oHMp
Zk0rfVWh8rEDGxAgCL7x9HPXVurO7Fhso/59odNSU1DJx29UsjMixZI/he9LTea7
8oxEiBOFljVo7SJNP48Sj7Vzw7hEKOdQDwyDuku/UJSaC2qAtJqr63d1OR7KX8T1
P2jJ3ay+Cljn59YQzt67cEAVKQeTljlGmdYBLq6zrp9naiU4RtmpYrm0Mu2OJjQF
YHkc4EgbQycX8htwXEPBk3o4LWKzUcQVHYt+0cmPvCGTrrXwNi79pvAnUtBdoz9d
Qe5MMKL/v6ZFR8i0I4VgczbjPB0pi4NQ4KNr7FHUDNDYITGuA+WzhnqEX54JfjwO
V4Md+YLUtmQYqkcnpAUxGYnYx+qgn/FAezLOtKkl4lUaqxxiqAzRQL5PwGZjtKsb
cOwianqm6jSrdQ10N2fnkErn2w2JQu8CID72P0tNOmoQ23kT3qEwb4Ul8aZYVFNz
G0Hbr//M2BIMyEY0DeS+nqrtd/VgiKRz5qD2P7KZc8ncldYlnAVmYhAuG6KHG9Pm
tF6xXEvlXRXnsVXiSjV94rH5Fw/TS+uUaV0qQC6/dwLIIOezNuGo2ah1XAgcTIVE
rGapI75fDNLwV98CgKEQhN3XIDVzxlnpDof9W/X1GJnds5shzGCFrf6kP1FkkiJb
30GRGsUThFjxAtmDQ6r0rzcW0M2H+ShR4fFCrAeOsAxRzae5bz3Ld0ZcFKKgkSG2
cHNgAx8uDHTvy19hPeIOC4ed21MTTjsM80tn6pI/R8lpM9Ym4fcrJiwf2wNO9OzY
ukntxHORdFi1Q3LtAcyH9SGGmo2GU4l5DEGNutA3FfsGATK/M3LOVBuy5b9zBFw8
bWD2xYMK75GMBt2DmuQ6Lj8j+yzQJhyONVc1MA2weYoGdETHt3SHk+r+AFHJKaO6
Xa6ABeBs3dVaeuUmwWhlB8lxUQ0vT+bCwBJEoNTGnyFLpGC/ippORhqbY4uly4lF
rganNhTQHN92mf6td7iH/x22v9pR6X17lcWgsymtQx2NrZNVbMpm6dMsaxfGvXE2
2VprS9/yg5E7CmacAmRTJrDREuY4W357K3b0yPyShvdTzKnJJXV3T/pA8eapZUL6
wawfw67c8lVy0IDUAbz8a1AmTr9yKAOc0+uuMi6/YRK5lHfA4l/Hp2OiD4TOiVbu
LRgfRhVisZNRNoVvrE9Ne74o9M94rtGThva9aiDmf6aoOoSobQIiZoQe42SbaLrj
zAz3iFruTfQ6GVKHmow49UzYYed9u7wpx5qr2/XlB0HN5RuHQ9Et2KRBcYgk0qFK
u1n7lpHhfI55nhUc8rUQoM6SY3tN4K7J3VvAcLnB9HDtQivJP28OP/9E3TyiMhRK
QYv/AwX9rsiRVhqCUpCaaHw/J4VtF933/jBgyp0hWmTavjfZjdf7qCgNwnjx8Tn7
5D78RS588lNOuXnwTnsvQZX8Rdu3b/vOvR8IjAF9gQxieXMiRq7KtaTY6w+4KyWW
pDn2342HLBbVk47vnZZbUGZkMTtqdiFE9APZdTqp2AoXJHDnrV4fm1x+DtZlrRbB
OJFYUNVVnJc/pM+jz1/LN42io2UsOlXzrIYezMYDa7IKfeLP1f/F0qhflhThG8/v
RSzAgDCLiMfrR2FUUV1YMtPsHxXziOCXAg/i327dkByo16jVtmQJTPzBNBvgBJD2
DKQ/vIyKdk0CReSO7MBewiLv9l5MKkhvdv2qwvMWbR1/OKiVSZRdPXW/bRKTxOBS
X13DD4TSNdDh/yjIiDIV/JDcROk4n2tDn3GsgeiqMyYnabjCazxB9zTjyZrGS6H/
9TT2jwK8oImQvnnW6yJXSS+kaXSAHQhQ76F+CAg4nOmCyq8vS69MJSIIwzgagwHM
0o5MWWcHUMdocMBU3yiEBOzGAnbVKC8nICtWgIY/fWzYDJ48Mi0kHhJXcB4xFcCr
o0xClBQcdHsvyKYsvU+PlsfRhSuco/b2v1oKviT5RRobrtnkmoj0he68l+/ksw+y
/fXcM2l1Bxyr1Ow1iovjggjqyY/khPmQILTj90hW39FEBtMiuntMfiOu4USQ7B6N
EwUm7dSvj6AKGGWtHLzIy365nWuzRW3Rw+IczhvvAR1trEqMICbepozr/YiNi4yH
nzRlEtuKgutVbBbEYdBj6lX9/r0JPl5KLWbqU2gZTNJ1rccCknvmwj6cs1mEixOV
CoUrX4JFRslvLeXGZWe5anekVDzKGCli1+gvhT6TjQ0fbr25foHrzZ0RQSw/SGdK
iDAHOrhLh7ZhZuN1SchRZmZ3AKUHQ3WQUhGvyY92kCTb5BLlXhgx1jGJsANwt1ys
9pjU8zY1pM0VC0g2jnI9snfKad7SzLwe+rN2DpryC1dF9NTvFIaVKqV3FKYVC6kO
mBXfJLgr+9x+zLG1pSIM1VBLg0MjSbpzgYL0N9S+TzXvf5+jH4PNMvLxcggP0Mer
mynLsCvwU2iAnYSiSxZwNXTtgahaV/mU5Ffp60u2bZTg9OYqh6HdVb8u3DIwPaLH
VJ5SC55dbXUo6TvPqrMrygT25ziHzPfdUSZQyr78lZZN1cvvwb6oOhwjN/6emQPr
ND+FEzxceDsE0kVaEk+lk8RgaOxDNW6tVDdJgVc/wn4a0mugQy6BzeBQpW/XOaj1
04IDD3Zph44BXwQoCowOnuYuy5TOjCya6yfoVohLipvDUyxnMsNwl3Ax3hVPKaHb
VzbBBl68aiUN2BWibAnR+mC/RDWZvWxgvX6stEaqSdCXaHXHyM+QyelI+mRSJHVE
vMdfAPDMIg61Dcb/C44KzTqGdKOgCxvAfKo6g3Vzo6G0LRk3H4Wb3Tr2gFoyUPmX
hPvGPexmaVyp4d+KC68kMiucsLpYFH20sifaMryUNEq8MtUTloL99zvqYnhRFxwm
0BAI5cupV4/ceMMwUedyCbPyIH1itAJ3cZT239QjwGj4bvkvCiwgbPzC0cJx/s1Z
vrUOrbn3sb9V6Rt1rkC7bEjnSYReopGITYhZfzdkTlil1qFEqkd3V/q4vZ2Zvifg
u8niY/01U2dm+JYT5+lMvTCWwwBwmYN+9jkuk4jSTu5qyiVNkVs5QXc/Ft5flH+0
gh2IJfwwkoTRv1qtK9spD6YnQ7XfG+ldy//DiZmMt3Bpr7dBZHst5Tn4rDC7K3UX
kvI3rKGCQzE5XBPgEw+faKk58igsOnXyJhsp+lUFngaLwhoruk1QOt/oL7axdZDx
CYaEUF9oJ6/htcmhLF6PsGOxIEMG1ZC1Lc8zabW1t03D8DMR5sgSMrnoHzeCD2tS
J/1FQe5oUkv+iF2FLYR8gNwBZg4QcrltJ5uLXTDNkz4aRNXsVOMAt6WfvxSR1eS8
UavXGXQyJT/Ez4kfFONYoND/1Z+gQ3npOZ/aclP7sI0tcK+Yabqlkc2A5YADH4nI
DskgXVq9AGy8UJe4V8WPEccAN449YhrnUwVcfMx+mpfyu8SXNMlpTvfifwgW0NiO
N4rp30l4/sWCIiI21PqRmH4f6OWK/Ec0z8J+2EYHqXrRaNfoizQS+VaQ3jfMPwtz
vmNoGmkQQovDvZTMFOGg3TZfDNgP1bpfb0xAeCdD+2MeA/1vCJ+pCsMiyKvgjaHr
y+3tjNTGF7bsSzUpnxGmf9z7xbJ8ZHKfK+opQE0c1LLOL1w13RiWFOv5GaX/CjhG
lc0vEnQ0v0ARLCE1qmhlmPjauBXEDvbZDnZ0KwHGOkj589eBcYCxBx0X5Mg4yr3+
tYuksiZji73LxmUF/184XW9RaIk48MGFYqtu5RNbS9Df6OH3wrH74HfZmQyR2tK2
9NNIH49lINFLu42Qy8afP7osM/pYdiWsFthoSmGzV52rI4AXcAaUbSD3TrjmVVBn
iExft9oKoJyGHolLu2saPtvBN+IW9TRmrPrmZYrEk6AJK9XEb02ofPvsD8EVzpnG
6oGd8nn4bkcDEAXNPYmwXrtuOSmXbXaiaWom3E0wbATfz2iFDXWNnmrjvQyYfCZL
CqxHYNmWZs37v42+WgOD0dPwHg+QlSuo++6cpgOWChMZ2hCaafEq1oXEGlfkcGGU
ITFS8gxSL1CdIS+rImLXy6IG+pGfpCdTqGi6Bc0ZB9lntaWzwVmUP8QmwF5kk5Ge
q+nxsgs9VHXntGT5euPq1WRoM8LxrCAEOdJ4+wSo/RKP7OEQU8YwkuCCTr4+ny0U
iu4Mov2Bo+wXS/d48W6oNdTPc5JYbpdReLFE+yCbw7TVCIpj92GbkXnhK0VJeGfv
qACTHGdLN0NxFo6kOENiL5lfZKuaUK8Zw9i31TDgP0P83VyjXcbNAdzFtyvz1127
wmk3V2C6+M7b1JixsZk20kZKRL9FUJttm5VhEYNjdsvfbPDbfNpaE/AqRGjtelZ1
hwZyoiXj6gN2RyQpKt6kImBlu7G0vp9Mhii1qWbF01Ed/2X61JgRRbkHwt1geF/o
uUsXraK4mrGpu4/XTP9dy8dKuZWqWRmi7eDwJndYJzT+tA4ReHnApeGr12knCvlF
dDB/gXz0E54WuwXkBgvn665prr91OtThUl0znfv+QjVcRR8PmczG+8Nt0D+v3EBW
vYnqZKSFWkw4QsYsfca2K+gmxm68QwX4y0Oi0chE+4jk+LdSKNFGnu+7i4ysGSD4
/n5SO3sCcJKAzk5YSSeVxihm89yeTFmilUPmaznqyANKf4PNdqBEMOT4oKj690iM
9JImVdl8TZ4hG7TwtUojyeC4jvOhMoUm4XMsYeAUkFQgKoprZ9xZkJ9doT70BtX8
JfZWIdj6cTxPdONjVAJbqh/AqX603ApP2OCDZark8YP20OXRnzyFHAtJriuJmVVM
0+eZ3rRJqeSCxQJCSGHuDliiQe7jezBzcgmKGWKJqztoRolP//WlQIL5kykZKCWT
WBi3R2qW1DZCW1XHqwtdFr3U+puYpL9EE/yOBMxL/uMNt1OXWu8Q9y6BP/ZxtfTM
4/xOyrElR+htiV3ziUFu4QYW5psOOVP/UYv64dqWtm+BpsuFwKY57Joib1WwxezJ
ldMH6nejCDrRxd6nRVRKO0u5HcS9QFmldKPFUKiS96dQ/rqJVzBDV7d3J+TyjJc5
R3wFAowiVZC8tzfVw67XVgu9AIarjaReMcskyRSnohEDTyNMYTDoCfndVKEuIixs
CmfGdAzQXR4UsanwbWy3b+w8wuH+cxHhkk/CG1A1U8GyS3QtLSTSf7P+BE741mpg
HiXTmc49c/rGMgqvNfzYNAYYJ/tKM0cxPHpWR0Yk1N7m02xZ6ekGtv2AEJpT7SFF
lwuLf7y/RpstxXPfWrviY+vzV5LyU1b8lM9+zoMRbGwTsK1ZdKHD5XcqsFM7YznY
1a7JAxH8CgrMx/sExzoNPy+BTeOcgTle96J5PfAbzogOrtyKlu+R5rHjLbiogPqZ
C9IBZEJxMnMr/sdD46XKIa3R5SY00D3WRYFOzlxeZvJIsRlQ6yYdEAs5e+YHCxUR
mAUbt8PUwx3pbhnc1VWPTPfqDMPKgp2gCyDj5qj/k/BGT+zsLZq6khP5VtUo/isB
+2kFjG8UkXFE95BKcKqs/ah2lZDXh584ni4dVxeyvSTkADvfb0u82wPw3sZjgvBL
Yng7r7iuKKTCQ67lf4SbTVyoNGez4oLfVnsPMKX8wlV5OttXf1qFHEbgTeDDz7Dh
bEXOZKqT+hTYLZqOwcbEhiiO97G4h13lvbv7ONL7Fxn/CwVOq6UzhXiSfIOqbsGM
LUz9l7qlgmB5qprXu5ZumWS0nR0Qiek37hVxzaqrVUU/IjarUNFsATNwJB6FnCQb
3YiaDbXeFx2+8lC5iT9FxSV2h5VqFxpijH7PaozB3wWRNQESw/fn7BtTt2mMEsJ7
WJFPAaxJBOWBocIzfRqdoOJDaYHdxl2Xq6RUO11Ve1IF8DeRsaAToFUXROCYYmdy
3Aepavrwe6fbIGtYVjjdQ8jkLHAiGltYCuKYVQ/3mFzg58GoshX8BVFVn5KsVxea
BZz3nt3I7xCC2tbwa6TRF1pralZr9Vay9hD1XprpSNwfck9r7rnah8yKu8L5r1pk
NSlAzY9HmydlA/6ppc1M0am1l8+QEPk9IN8x9PuX9h3ghCYzQ7RL6xxdqcGxU3oY
ABlSjxXLIDqidBV/+0aIr9atVtZuKn/R7Fokg92mDipZAcUjyBHiFTex96EmykrY
IMp+rsetxHrfzkQUJWvWIalcsbBWjNcNAhZu0vn5nxrCni7rJiDqeoUaHo/uBxQD
d33G/PZACl7T9FXh1B0hESxNqTaVNUXCdGI6E+ZEQyrlI7ZuG4p3q1QbivZ/UMzS
cRMKJj0kaEbEJzD0fxQgvOhTJN+wJKvbkCDZsYiHntnN3ynAoxOWSn3AbLvrKlhQ
ZwPPxr5bNSqmF1T0nMEvj9wMrQHyEJxFcjkpp61oK+P1k05CPQOOjqJoZcbTOOkk
U8VKhp8rkIVG+KWPRb1T1tpzI3yuVF/PQ3pyEX8s1YSEmKlo1JRT2XS82EtEeqSa
qzCmm5DM1fLlxcQUgtYZk5fl/q+2OM3040VkFh88ClbKT9LIUY3o09XEWajhoJgl
LsBG5+npFgDxYyeSDPj1w2PQFCFPg8OLnGOMqVJPhYQgX66CWUSvIwDqC3wktz2f
MPw8iI2Pb9gluwI4ABpqZHeIkVKvSELoQSEkwvZch0x0AysMNYzIeJDTmzOK827H
4INFlY4B6AOJqH1+Nv7c64RBpJgmMW5mHbCvRQ2XC5wwAvrHqRstFqBzDmOwUnbe
LUNsLN+rapExVHVK65/TVkZxV55j6JRrrWQHDD8sQIjmMJxLDwNmG5g+MIYViUQq
+PPm5A5n/9JzJuzFJLoqO29hiZ4jvV4x1FDI33wfaNPUWPAQrN+5aMi0wI00mNRu
pWunU6zbdNHJzUL7vwESwIvgSDLCNSzG4FVmgjSp++PaRtkHeUee1h2nkmSDd8h+
nKbCLyMrDBeOFXHQ42leY8G0/4VpiM7jtoJFPa4oPRoeoS0w3wDDzRugurmJvpYb
zKWtDCrweCTTFft/JxfaD7HI26HIW2RDcINT87KjaG60PynhqwjXwFbSJDI1TzLQ
UTeuPahldvPLyFUIQoUuHBP7OXzTGo9dT+6NYR3xCrs7/kcgV16UlOSYXz9A7ktF
srKtrt3TGPhDDAjBOpTpqr6pLtGYMVf33BHdUaf5Ingy2KOY8KtnER9lRwWReMoN
wBv7T8w0PTAXqHQgaY8Uefvf/ZWOR48+9Nwz68xhaD9yQzwmxK3xFqCL6NMASEzk
ZciGMCk/axgQtoxdYgLjOq6Mcci3u5qKU3cVVeaghsPLbUrKpakVmfx8OtMngo1l
T8hG+hWY5qNmF+NBRPkTeiwasWx/06Dc7egMw5vl4dyQoYzEEiXOJfKexbjj0PLw
T3+sYU/q1EZp1vsGGxOjTW9aZdATMkEJkIt0DgD1H8r1SLXQdH4M0jSwWRqG4UJ2
CxRA6gPVhFkP/3+FCaTHLlmcWfLBRco9mK226MmGNAmVjn0PFdI9GI2fSrUMG40L
f3pzu6/nmfPl4YF87n04Q68DJ+cg0MLcaJkgS/YMki10J4s96zHyzlI1wOnX8fwI
snBFYSBlUT/xpbjP4K0UtSVcV6K81H3TboRMLvveGi0OFjCMPO2dCCMREjtY0Xt3
t5a/xSYEJ7nSQ0ghRCtdHlAzoGutKldMT3Mg9yjty9GKT8Bl62+84OhAPmL32ed5
CyqjHNBmpcMCF+w6Buq9K82K77XzVZfppsSgIhmKZAoV5jx2d24/lk5l+2ToZby1
5S9RpIH72MqWAmmgBlGRGsV8gmrX4Urrpth5x2M8+GnBeGofRIDe0kJZk6VWa9kX
MgM+FhOZkDbBv4ers0NuhvWdP+hlKvmedHy1HzUqIcMUAeZc+uHvSvohKkoAwZo9
+734HPw5N5JBsRsG0i8cByLyCdo7zqa901mwwI0hEPvNWHXypuPLQNyViHTMeSDO
hVEic+2BXl2Is/frL0iHM0a5ozVgqhFsd8qt9aBziOEz4uHDsQg5TNQbehRmkSuf
RQ/ZUtT7UlctjBW5/uU+QJic2GN4xVyxB3ytxnwFs28HLcs+Z0crN3GGqzpFUWG4
OxivML4BtrnZbOlMMiigg2y4wQKX4W5vikRNjJ2xJvRrGj1Y2dGlyW0lcer9b/5C
3kd/DcBS1U7pA5ETUJ7Iw+YY0ZJIlnnu6MHq49GetkzqJTVm5HcmIB07wZB7xw0u
sYF9UMw7y4g+NlErGeobVL6AAAIDdxSroAeho68zKfqtGw8HTDsimUu1894GJsQB
BkA4egrjB1oZivJNQCLkgdzLMW0kQSbiiofV7GDlxFKbp3Z3OZtIc+MC1f+wdVEJ
O5ReO5USioi80s2gKKnUHv9axST0sfrqxy2LP56ckiMGt6cRm38kjgrJV2n7QToU
DjRClCiT2zhH05KtlzyVKV362HXoNASOylejq2Bn6+znCGQqMz6xNojg4nX7fRdu
hvfFIWjM6QSsoANONmW67PH9GRWUfrUlBgu/Qp+QsUuo51jXlMValSY7u2n2MBU+
p221GvSxq/VPRWZc3m7L9p9kl6D/s2IuBReOEXVPuFGvS2v1H7NbK+z+hDBdnQmD
pC1fH37VwMTgynslT4SBpE8OXFJXtTjTRg2iSqRkkjTgShYcjMWaVls8eWOCIDQW
tRGetqo81TCc1XqetTQR3Ub+o1Sc4EPoGZK2iPle65owGan3JQjb21tBam09rJug
gt+0BVmfIGHFKK9VSH+EZJdsi6tISswKbbCm/TXxSajWBYZnpHkH8nhBwbSmUDBq
lLwXwvSWdY4L2/3QG4I2VYCuV4plHmhQGqB+mueER0AxEWfznrc+FXIOKknJ6aIa
Qy2ROCQp8W52LbryLY99Wo2liuQnyhyZ8cH1tUk9DSIElv+k4N8Wu6IeLJEhneCX
RAmqzw2BBjnwQbIuMRmaQH9Yw4y39+uFV0LRs1Buj1WtGjZGOGz0F4Bf6RinjOHd
DD5IvVKBZNljX1CXtLW//iGoqhRJr3sIu7nf/OgaRP9zWht/x/zDIOxMPtu736bI
UV1gM05OzUkcqrN0k1JlTc55CDrShc2sPcU8PDzXMWfxSbSoNqz1RK1ZeDdB2vT4
KMrzSZrLet6OR+KLMLBaWwjv3bwXF+8swgzqVc+WHoqgImXAHCSMhnkyQae+hp+g
WmdzGqp3fd703sDUwyatFbor/z+e3G91seD0RS80JzKzFpUtWsU3pDj4wxJGMYWN
A4IxDRpYYIhXfa7jNW1jUx3/q+BQ7+3uVQtwbzzmmxmP1D6UHD9jQoGK05Ls0c/z
CiC3OAJeMX0nuefWJwekrJsaZOOlxClbxDUw0pjbmT7Z7dJL6wBOEKyu8X7zxxzM
oaAwUpiEJGhpCDmdcnOaawgBc63VcUDwnYruI06Y3g9QORoARaoZHgCWuvONlc1C
TnL0JYkBiuSublG/bQpAyZVZMMx1lF5eGcUGKSN51HZTQYK0hshkRek9y067+7YA
c1uabKJDOPzHDpmzbvpM1xu5/5UUbaoaBsnohLkbrisC8xPdISYXMmWkRqYILm66
sqdJOMQo/DIv4sJtpNTpRc7q+7xbKzMWp9UkHIlD0S5H3NS9zdgXUZS0904ZiEBE
+8CZgpoYeXenqfn4mEmxNSb2RmcfFmmDV6Cz6Jy5oa8GTTJ2oimeQuEBDeTjp2UL
Q81VoBzOprr+RryDSrkUgzmTy+qEDyJ7Y8alG1ffiWuixFEdbbJt1nvDe3IC0KlW
/Smmket0N0gsS6D4fThhdifTzYV+K3XQsZyePAjqJNp/s3cpdzAIUmsJkkvazj7a
Rbjy7y+g9g9byFNYnLDe4MyFyiF4OSmcXGpNdeVpyPwOh+mo9NS4HPijfq7o0QFa
MhwJ4sMciuoVufUuc/i67s/P+Mb+FVk91nhIcGZhOBS7RYZYULmnpES6LRRhTkr7
yCBtIcVw7PzyVEqtZ9krKbKIcYPgglX5loztBllC9z9pmOYowNm6G4fJKi0nJIbi
XQVji5YLIn4/3aSz7trT/y/6/Oj81ni1s0GJdjj0y2HaDFhJczXrTgUJkLnLCcV2
LxfRh5jhVAuomfEKLjRiVK7egHh2GiigKkcokcDhbf9XGXr70Dnd/GrQkqpoB8ce
rjGq/1zF+bh0gDA7jNdBVVdMnxUwTSHae11nwVMuZdcJYUqf7DzBTfjCqLTtYkpF
RxvXWR7BTTVfb78sFVnHtoxH2EGWAivCzUjQ0vNUG2NA16afyVvqjlYyyK6Z8AmU
lN7cQbV2AUl2p7Lqsmy8pXoTkas3y4bhh+JzPsoRNmVDNl1FW6JrKXSOHfWavOPw
MIASVBymFltLbaagXLOAK/NWnSUm9DWmhF8L0hM81wdC/lmiIa0RLQcuKcFlAEP8
275AL2yGvqxNOijt/pTuiFLrO6aHotGXYS1rVdmxCd1UrfMm44UizHDxEbIGSAb9
kXRFxg3e1LTAcQ7vcaLMoc6yg+Azp5h3wxbfnMhCrz1WSKAbUFdWwZRUO129+e67
VQqVUiIoDDhENSQ0vlo74Up2xMEsZWB2Ru+v7avYdfphCfT3q09VyVr4ZowX+Id9
hTKsPUx1x581on8FKMuAOM+tqJrjpNPqT7MVJ2g7JDX8niKvRb3vE1jTeSIr7yLf
sON84775L8W8Qe1dguqSphwp05xv4eahM/9uwlRad0rgTCIBJJgFivZcdkYLPNLD
HfwEMBsQZMQQKzBqAmtXc7UwElh7Fs8vPUssuLbd9RUXklNovkcr+NWBQOhy23Sb
PQfK100jsrMgC/UnSyQ82rjG39ojyLl2rHl4gZAo3aB40W0TekxIXMYRsIQIDcDJ
oYbCy9ZQrFZB6y6qr14H7YKvZJNLuS5hApmTCnOwzmwLMaXirgdFcnBUI7lEPHDq
uygpMdyLf9rVSyDclNmLV6YwNLI758EK3+ERq7FkRQOG1YViK7s/6AfVxM3n/pM8
siw2zr/Ggjr1qYLjDC0YabKxavV+p04eNuh+Ea+lPAir4aHtYoSygxxHuYyWFqzG
T9WQDpP4G0zkpuN+hSMRftODCpN2CfTDgGwhS1TLYo1wJczDVPZnbxr+JbzozQOE
PYq3LGJSBdokjad5ZN+5Hq0b7+aFZrLOfdupWsqHwa/0vM2ZPXsQhsYDlZm/FaeF
AsCYKNvNdHUAA54DL51yRPxAFzvFbfznhROpX/eoLke+fIzpGv1tPmtdl/PBbAp+
IsdunOI+fLdt6m4O6wZpxqFhs5BQ4Z6uouq+Sx4AV0JBUVNIuxsimAVm2zuRfF0P
DpqcnygtjKltCHXfPyKTJwzbtyRTi7O+qF9svh9u00Deq8vh1Ye3uOhsEY5JaLIK
K3AygK0bfdFyAX/YjxD0VtzU+a5YorrXNTjS7Dbsu+gBh4deJtMlrPt7fnevdUGr
k00W6LKBiRKyW0CaDaL5Ffyj5i5yuU0HtPvEmJhXF/I7tDJXnHDp5nxun4/PbYU7
AzCCf+9tDGp6qEMlqKJeGADwDwii8+asG+sRTz2tHXLfy3GYQzYHZUnkjiDyMVP4
9FetE+55qTUPUMDfT3sFDTz3RCH1lRfjzIjlSIOVteELZQMV3SnWJBRwpZdWJ6rJ
sUrCFBRtDOsaR2RT+SDmDHYmD2pUa3LESNrLpVUxywQeZtkwcs5Ga//zK584SGG+
LNBykVawXNFzJNXyk/Ztn6MMtFqDfIC4CoiXbVrvJk5rT9znL6UTf+w00RsH5x/f
jNUplVxT4m+hq2uMJ+lvg0IiHPkefZDAFbpG8yAW2R3YGa1Rl2qByEskZ6wKNjNi
KlyQjxkdUVI23YUG4nY285YpJbwJH2dpCiPjCV2fxdVL23q+ZPricycBDu4JAlXB
xg0cjtTejKPcakUM/T2dmr3SEqxnpf2eAwyiNUR48x+bQNbc5WPYCnc7rKkeumQZ
AbZxKnD2ShvYTxk2L9JddZwDych1BfsCa835Ghn/FmdcKE8IuF2+lqbmAQ6XC5iO
qH+9kSi2SO0D3uNEuY3YcbPW/8s7pLAjfC9IA8zOXrdsW57sW+WQr197r5yHsurx
jlNosQ83A2oiDrtDiRe35jkpg+31GiGo8Vaoe9MOygrALf7tJWc8j27UjjwvFn0L
pKyK7J6MK078GsCCpdsatZrKJ+FWAmdcRr99Hh3CAR3f2vsHBbD3XF9BPud/zt5R
c3PtpYI7mk+BcZo9y2JVb5dFmoFKtPaXPnucgR+6+R9C/U0WQOcDYEvRJfFriMEx
+qsnQQ9qbP6l7O93LqSyRwtabCSbTe8XyPwp0f7L47Pit8y98krNYOJZt+R3mPr7
gMXFVnWm7rSYJhiNgmeMwpisKbFhbEOmzZauMcuCqPb6k7z5Rvy65iJifPMrpU4/
x/XN/0BTdX6N1FTcVhXDs9/fhTzVuUV8IAJ8af0rWWwoEqGnu+zfyQf0wglqU8i9
HU3iqE2fC7hkdE2wpAInjwV/ip+PFXO4Pe+CVOIru59mFCKZ2XhjnzKYQIuDKXBU
/Fa/U0Dnsu985nqptuUQGYr/l+1D5ld3qqyotQIRrs+hLDjy7v8Za+L+wUHUih1H
KhSq7IwVUKFHFK7VZhUAO49BM/JJ3Ozvo+0TbFLT28QKy3IgGm6Z6/RM1DiZ+0+B
qPDPeah9E0NeXgqxUA0hyip7JhJv9dFwbI1ibuAV+gj6Yek0L0vYwZeQfcWZI2mG
UxOC2sfZuuTGehaUhR7KQcSCWqlJlAgkZgnbaHzLIpL5bmYJS0h92GCNYa/Fsm1A
+BaHQKiNBmPcQtaBMydLg7jA4BToLzMAkPDs2ozdZF9AZfuZiqQGm+CKR3QYGv2p
TNHYA/ujsAx/MfPtoH0peiw7De8xdOyxQP/eMrt9t0Ljbqi3DxL4DjXj0cck+9Na
ZkAdgvuS5r3rdpLbqq6NyQQbHrQLX5jrEID3LTh1o7pD5qfon+YLgXhyTMQf6vfK
HPSye6/tSm4jvN7PenHYieBUCrAWMUoTm6EhJNflk+jKpT8cmc8CXCMICbc8yrWb
OQG1mzKTjfxvlqZEluOe1aFEZsa2RORKFwIID1pmqv/d7V/Al5azB+jpuGKbzx40
rAfl9ntHbu0G+yH0vry3TApVFZMr4agV0rv1GM3eOYgCINt338IMPskk31bxSTeZ
gaiKilbXOr8vLhyG9/43/yDAM1EIGtyUtqTVZAwd6HG/sdOfLCS4vUTNxQ+IYXkL
q7a3fgH3Jhnrznpu6E/AovHSw3koRyq95uf9uaxXUl0GYiXkoPuIhWLkaSeyGQhE
LR56WTNNgqd2KjXMsRUiiKsT4Iazdf3UhcOzdyl1cwLN567AxiJolR+PIj+QbVcM
hA8xWoJzH616aV5NZ7rSCRstFafvmrh8FklnRyv14LFnLcxtD+Tu+ARAbq1ABxBH
rwupBqppiYJElzPe/ELF+7RAzeyyilUS3Ukz/e2j7E0TMLNF/1HYMisgrsBgvpOk
F+aMrDtGvQ40jL9sYl3bBQvjlb0Vus37qXRnjaIIPhNb8jc8P73969pnc9VK5CMa
3ajs49qVythNm+Hnt+UfbqdUGm8dwaGMUO6XdqSgbK8D1Zo2iop8k8WBo36nm0QW
T2+oRR4WMdRfh/S6vaZrkaVzpq1ciZq9596rA+2MUqkUclvQ01WlpYHj2MgjXqNB
YpO0s3Ypp75JpqvJt6NF2XqTc8ZdZr4ThiRRDtqXvV+PAZcn0KIN8W2tWssMql5e
MK5hccT/2Yh8wlebkvz7YXZWSPxhWNeH0P0IDoorqjkQlI5fYuvJUGI00+D/LJ/V
W405QvzBgavmHsMfGjmnmI5lnoLn1aAbF/nNrDhdrgrUUFA85Vtu6yYlTlXJYKgS
I19GzkRSI39SZu0JhKYJbP7Gnnt0yZHGVK5XsGWzxUm583JESZsUMYMALX47YZwt
MQiqgAU/nSEFU5LbINy1yyTyx108oXF20A3Nx+/RThSPenob72EyHvX35FkcF0Nb
MJe6s2sAgcmVajA9NHYc/NCSuToZldLNKI6F9/JjyHarXrL1yoBx45zwTCHD0l+v
yMCYY6tz3ENk+g/51kRYTe3AUyMIM0grVPuKLSKI3FpRmIkCR19nYqDKSfm/ZykY
RQcuDKVw6Z9y2bcjnE5JTzox2XIx0X5EPk0CSSpAhJAQFJuJUPb3Aw74EL7PUvef
smPOhIEWpMgT3Q9mX1wIiHugbXXiOxLwoI5Ll0oOsfFg4+NwILzOmZDP5CR2b3c4
Dl5ff3N8VQUGcyfWGIuxKKf6zqtpHPCRE47bagz6zYMpDrdhtEe5YSA+zrwjgNdH
cIizZ7xXiGMQ8D7EUKSK4w4kwz3aveLyZyrbsz6empGsEv7UNK5APKawpB2tHKO5
BQSl0o8aPy1tMIzFkhq0DFvHyGoiqFnbcQpWXIqPpMn/7iILDZz70pmsfrnbVnuA
3RDzJXF5iIbwRwJ583JhRip36+Uyj5pUJZ5q/5jkJXfIZBQBold5yJLEaeBvcpch
IuusSMn0/8ToG3vhdZYEI2Jh0MXq9FKCykoMyPWFjDFcr8Dj28v+eF8CBdYNGrBJ
u3iB+BtJQIeXGeMPT4s/YUPC9QzGARSNHmjkh8lg3NcOy2XU+spv09bDYX5idO9Q
yV9sE5Mn3Cc/RiICClVwToaixIAqb761Q/fLB+FjopFXoiPFs9L3Q/lPSRcS5qJ6
uuZEns7aQwhWLLJ+jjwaJYvZYZAYP1NaxIGlEutC/bTP/8G8GY/mwKEOij90c+T3
uqoTJOBB10muYM0ZFuWbP16sC2kBhXechlejMaNAJ2rDyoI3l8dWnvkh05r+sTAH
E4wU9LQxT6uIAuliDNY0E8Qw+dCmj7XC2uGG3yROK679cHvWsS5vj2pRHvwOWLmi
LsK0TUTMNEoStEWQv3F7ozqVGBHsGXJvPU+Qw5jSxVItg1486jdCLYL8yiCEKYmv
jMuAWt9u8sK7o2uWuDpcIhOC+qcr1zCHvPxn6DFy3Nit24Q0gxU9qu4dR9gVmWzm
kSmYJEZDU0X057W1IYqdszD6VMfwbyNa4RpWt7RqqKJJt0jIs6hND6aAQ2ooL/go
Rnm1bk5FtQkYke7yW1i6K0NZ5nEeHewdUH2DvIhnfE/3hbHiOVkKF2laJxW5Yn5+
np/mS9n+nf7OfqHPH617zmuMGWu+rFSRuEhBAyCknlt5Xr6dYGVumcDI6lzy/e+3
ghVnhdDyupyriWjPNCBtwOk4+rK8epSIdfAJaMq3FWJeOc4QOMThx5jmYy2Q4QIB
YD4+aUAwt9fy9eQLzDcXAPH92KHvm0Zh/OPka/mb9edOKZkS9WfOvSUF7MsOJSUn
2FKgDfzWlZ2jtxTb/tpVGoEbBbGwTtohZ98bIaE0Wo8JJeomeu8lGhX52gHjuWJz
XP3YlcH3RqBf0jLA3YljQmWDNmMmT5T9/3IqsWZRMa6xI46aJeBiTrmFGaqR8sXT
GQ+SFAf/1hufZmNLj+5cmYz3N2sIK441C/bkS0TXuS/nUzN8/e7cs60JtloZhEsh
mZoipvzsMR6FAr3L2Rnpz2zpA+7KAkh3pE2kZzSyy2YtRfhT+MISA2hPh4w2YDlD
ujr6ovNPBUZabq9TzjiIuPBnFdHybBu4hR5DBNFhNn4txrp7e2C6D/+7zoPZS1+E
jD6YPNPude/P3ss8QThICkctlH1x4+IDEdL2j7Fk+q545EWqTZMQZJxvSETLnPdK
UFrBiEf7diz0csFpl62yLxJMAZwQJpd2MEyo5eAqYTjYZSi37csIwMMfUaIn62Wv
gZfDdjvhcDU3Tycsbs/Q8+ecHPtDXT0dY1wGLRAOuxgMPluwoc2JLjLanEQrflC8
us2dCsyXIlojuc3dSxeuJFIWoXuUxjvFM3HUN4SOOK1rRAUeBb8N6DdUrit0vVZx
ZO4XgTXPAnuPXHrgCF2NOhGmVgxN+75o4aysp6Dv6WKsgG+Q4diCfhV9ltTUGlZ4
L++NzxAFRskde9e13FwmFyRsOMG3zyTPz2cvj0do+A7SubrGqtgLT+kZO350B6ej
dOosdrdjxW3x+kA7A38o0hiQzNfFZB6vRxFGy7wWZW9FMxnwoGpKScLaiVR8tPCu
ll3OfD7We/56wEcfMFnS1ojYS0k3jCMdHQSy+xIueQNn0viNydx6Et+vxSpzXV3G
2qKUMRJI9fazMkhjMTZIjikMI5ienHQKcw6B4eCEraGTc57dmG9sdR6fJjXu0lwO
De/Tc5PRWg3bpnpSCuHFAUB5kkxNlFyn4+7m/N1SZRm+nCwKtWk5eBeouy0/wiwl
fTBilYDGDRvad7Rrd7XsH2KRtTwlFtJeP0yJGk1E+BRyAoxxwF+wichmhmZFoTm9
HaiUqpV+rWes9jvVKtHcwbtIoJreiGIZ96NzgzZIc7kPVp5IeW84uvYl8bNvtu2K
le7/lcdkSL7lvNbqzRItZ+v5NhF2rDFNo5uv9UsKLb93yAxzVHGxGnmeTTVQUirN
oQaW7hpI9owhKmZnOT4BKaPt8dEpKQQcNzCu/UGErPj6YOkRLvR0P6awvPv8Bpcq
cg6ff9vASXeVs6KQXKraX104nOA8qT70Vw82JRVlbQLJGPCDu1zG7G6cAiW4yztS
ndPX4GGpB8geOBo/83TMiD2GEt2tclOFd6q8qj9WBxtLlaEKzlofkHmO1UyYQOJr
Kgoq608W2fSQGo7SE7YFoiHQGHvLHfWhOBbyewqIM1KQ+yLp2BaZddkbYP+dnZpq
T0VsqIxidc0hoQ8f1Mz2RdH2D9wxTAqabjpa2xkuQ227qlnZpl+sA05VLFD+tyCh
C3qUxqcIJKNb2NYJDPYb3tYpW3yW34BhtIW/AFNXB5ieT46omw9/U5uzK0ziW8Ij
0ACHWpVzdGTqTAZ3nKG/cHikIbDT8m7UeonbyaCgy3nuAM68Er8Ee+efJTFnITii
0q0QM76HbSJ25P1Npb+fx/r3EeaJU+FKn1S8ReVxuQfTlwzB/PJm08Y2hRHNMi/A
qF+9ZQ3bU+LrIxoogM/XozxqVQPET9iz/ofW3LdloRP4SabNtEg7R/bb2oirzN1r
PCLPdGFNVmHNEJ0f59OzsBy+Vm/9vqhAmHb6WeGeuMWnhEPz4u72Q1Tgo5Cq2ZAw
pRY0bwlVIQext9CYsQYMNYzdN4pLWGqNzs3EJTeRQGqXUTIGQlYwWUQ7T+7sziQB
Uutlzm/mbwPFvb/pRLewzzTnBayBg0Mmc9tscHCRX15LYs8AjEHNtxZwrOil4lh4
o4RZjPxBt3SnxIC/9gvhgGuq3GKOxpjJ1F+fmxNQue4cT+oSFpUM+iOqk73AAEQC
KsxfSNHl7eKqDd4P083QT6WgJsQ5G7A0Zdd3i40ujcTL3y29wYwcBYxOmMQ9enTZ
uGO+Rqv2wD1mrrdNbdBwUch0EmXimB8dIBHBmV+EARIyymo3yRDp6Sfh5GJpHSIa
yMvzs/aGhN9BxW7eHoCFle/EZcpgtMPjPuVxmFOUwX0I1Kk7eN3up2dD0pTDRFt1
a0q+jcSg4OLp7B60gUftaPqm4w4FUp7Fdo2o+qQWXKuIjfiGmo29NOcpnxg+7mLH
hEDBrTJ9sNWlSu4LjwFyeeyYyriDfO2ywc5CwDojdVrygsIv9PkY01lnV192XYWF
wntSqdcCsjd8dwOEHktuxSYuQ+ybQSMBozOH2XrofIyfGW8Kjaw0sg5mI9eAJk9J
rgdeEWmbWGvBsqhCs+C3ZrJclbzhfUBpR6oKzEkLMDToGLL/In5iGoFWYdvkkrCA
Yz8NmdlQrM7/q4U1uJvCnsGiVR0IG52Hpig2tOMYa7r88q5Z/XXunAfKNhqWi1/B
+k6LEiNAbZbbvJpoZyqHBcfjiXD6BDiW+4Ez4kgXG1uo7BzeETMDIUiO/r3nOLsQ
JRXvLTJGBrh8Y7rsHBkt5HgahpSVayldkfVM8MREe/ai9sHQxv2coxnguUr/9zS0
E65ja96hvsScZVI3U50F6VMjEATydc6Cee/l12bEk6FAhTzPtCiZvwsPzw5TJf25
Mx1BVy1BFzDjHoVq+TTAAVjWoGz7hVQV4ukOykFgeHA1Obj1Znv7NlXvv/xh6Ape
bewFj0R5Rpi4z+OYNp2kLmeHf29E1pfWNv86zP3ePxwpLSGIhKL+glmM5XwxgY2z
PwKXRogfvZFWjbqORPEKz7jSCpvg/u066hqKXk3RMoL8/ZzIKHxFiFO7G32CAR4/
KrRRAIHnsnGZS/OYbJo7/xX5jA4RSJbcpdR95ZlPFwgMUKNINAs1fo7/LBe3zKvq
0jaWpRltzCJ7wc6wQVbxesmQlTbuyw/6GDLkMxEQdUqxJBnuhWq534Y4pMO4c2Fb
lOhYChIjOwftRcNqnNGuqWrrPihKiVdTeR/UHkjORtua836gW+d0POym0zTRizvQ
DpeZSIF596oriXuPRmTQwxEa5NAj5pHHjKXCZtrO6Haf4eATJop8BxKWzyFH3Mpm
hRKfNK3PKhV7H4g6aHYBdRZXbwTLkym46Deob5jyjuEyQ+X3+d6htgC/esP6/wV3
xinTEyTlzoEPzk25guEqLuJGWKdQvMXKAWbZMP9gRE3kk+L+ipPJdmEnWIJusTfu
gh+yCKLA+2iKC92ViACBobfyUXzmB0l7NH2RlSP1eO6IbAs67wMG6Icg9VMD9063
guVmZ6EaMCUn6HwxcVjU+BCxxLTsflzikVsC5AESGLG6vNNNI2wQerd9Ku6aoZI5
FJK3IQ2UwU1Wdv/+QX9xL/KtwlWuc1HxvpKMDOhvLnTCAu+x73o8Fj6AQM5OY9Gy
nvp38mkAB5xsBzFOLIMF3ZJ+MiGhKkhICfepp15t5liUaB8ymuI2Y7XIuNjMVS7g
S76wm+Pk2kEY75qXzIDtxww/FFee2GhSVEqDYypNdP0dzEMfZX+zkpcIDwKW/IRA
MkLtf/6mSXF8V/SfY+WR4UPNxTyPJG2Cxdn8RrdDVb7IgLd24JMvt/p2JEHF9nzx
SooqBNiXuQJR99oOlbRZrmmL+dIaSZDL38+Y6U6ZV9k8+97dEfB/QQBs9Dw/dTD+
6Jh8rHwO8a+n2GtbJ5Kh5rE1eJD9cO0K3NlaMjHC+IihQ9Fa7GMpHAMGMSoAiD/8
bES/bxhSgRefsE4/7cymaY4AP0XIONSt16a+adcBeE6lQkSRKK/jiOctX96XLZpP
QZM97gAmFyxxpAegnFBbjAtlDzbz/oMu9s8MpL6Oo9/B2fEbk1wXDXKQb/Xiiumq
jwr8E4HNKxu8vcaXFbAcRN12As5WkCxUPm6qwqSr5w6RsOQ1K4y151LAe3H1VhsM
qENhY+1Ajnw9njhkAqLEqKdyt6mAxAw9Km5XEj8yItaK9OVB+Mc//GqCs4lPp2r7
mzgLtz6yIsGRWvVnZi5xfNhZuX4qOkg9f/RfAgYGZndLB0bCCtXzH+daNUeBNTrR
3e6bJy364icCt7J1d7eeivZ2gJ1expsjDiA0bd07HXu02lk7mEsU4xZlkX4feAzq
8GwPdRvbcZDZFbYkXUzzDcA2VxdoHOjIVhr6fM9rUHf3tLAbwGtWQG2P4ogt9I3k
SH1jZlXWH7hokTGJnGq/m1594s3isox3NN9smZhmiyvCeVCEKP1MMCfqxOOdMuvV
uYQiCSQlTEKIpyltVUIbhHQuJeWxg1WhGOqxZoZ+bvrnYDWJLXDhUwcHsACNhqRb
W5Ox3YKZ3Qh0bqj8fEl9qqpwmtjQaXDmrI3YxkQtAw7T4ismgbJiHI+tQVbArOTh
ypnoTAg0gvPsQYoBPc8BBY6uLPk7BkYQQVXZQ/fR7RZsf17QvVsStYqqjwi/Ei33
JF9Wh72CDTNPkQ2LbCqAAoCXuZcxEXCWDD2Cw16DI2b2U+npUjZ5ZkEezDvIxp/L
MfKhJ867ux9yqYJI1HjQ2QIbR9jOK6CGiPEKfo+PipN1ik6xKrD1K/sqQCjx+gZ8
i+DIclpjR5HuQ9jg96XqPGJAXqT9s81A89avv/2+o1vkDu3OecIZUo6LIe1EXOhE
JOyh5uPeuOm+GVgOl+hvDqnVq3yoWMjc5EzwM78Mo7uTHG+FG0pQ7FpyJa4DPU+z
y0Ws2sdis0RTZjfLZouwxCOwjUZtdRnaej54umEEzw/CSCdRZDAVVho4+/w76uAJ
XaCR/YdofVeXw8nFGKDL05qZH07rCy3btxJo9glE4YDiAdzNwHAdCdbezMvL/iJR
CCSlDcV4udDPQEdoqwKXm7Rv7MVuZnZkQseSACkMWbIuNPwgDccT9TQzr2aI86zf
I8aGD+1S8HcxaWz1+p5i+CPKd2HSCi3ZUYMqa+Pk9sMYX0tt5WguMSvhW2FOCJ8J
BuiT09nSIfcnGP5aMutNc46BnQijbessCDi+liPNMvaMgexwLL8lKj/FB6DqWJ7e
j9CT6yNtv8YIf4hURCrm558xFDMCJiVoQBef2wt6/zHf9gQcFDsZkbbXOHdWlAdX
x5Hpz5GCL1JBYEswjKfc//KVpqBUqXjEY7zWGLhT+AHViikBPWqIsi/KUhUP7pbq
c/UvKuRv20lfCI2FnA18cxU34a0vXd6f4LhfuVHwSyu/1sG3oF9uqT4wfokSt28+
vLCm6k+BE76N4khtSGc7pwp0HUKsn9toXT5fQuk6ZaY4JpplWjMi4kjIRMPSHRdD
lCP4bBNbcRdXpmay5Djr3XNgYD20A4l/U2dN+WJjUEBppaRV5DvORctVAjvlN7c0
dFHN9iJdgWMnFlRkIyT1TSvenPC0VmOyjb0nxk1HE7eB3r9n2fjfNrOV5tfRC7SC
aJLKnHOthMnujzp/0hRQl3bxRI9wLa2w7E2ZuprBno38msJsjNZGB/NTyIbS5/kK
64kT1go0IXN3Zdqr85uNxz6B7TcJMfd2Pgb1Ld5sjuiLY+QYe2YIySIFA22Q/4BZ
UCVlI6LCRqDHXlI+MiP++OZW8co50mVAAOSpjcxLQ5PIYGVfzyCPpaM205kyReAG
8KTCYhHUf4IqAYvasrYZ+7oZMRoV0EU6wSyJS11szRaJoH5NtmrsEe1UDMKzRU7m
VBlqGifZFn9gfsEJF3XkmLWpeKVtoK/lhV2XZarJp/beBzCP0NwdTx2rdZvEQtoS
qERPqdT1ihnh4zZ+E5zht8BlEpLAEt2FmfvSvVi5AwdCwfAe2SeKOxt/46t04+fW
C7Y0GLspktnyeuX9yytTUqrCQoxGF9fAOfv0ryx0ispZmBz1qbf2rdsgPf5csuLc
6OdSwrg4MW0xV6zyP+pK/v+lpzUO60nf+PXPlsNXZ8pORVnUvnJ3mkfFfR+kratX
lXpYJboSGr+qhbgICFDlCl+dklOBugaASgDz/X3nU3OatnQHv0ywx/HSwZdM4J5e
HXn9lvjej0jhLTlSufQOeQUqbGJJfEO5mVqjxyPmVytViGtGT6qRG8kYYUF3zfce
iuLRb+aARwTMp9cDTHf1CK3JOQhueyzv8YQ5uDbe/seh2DWz7a6FXoyJTnk3rYS1
sWqCohED1cueklHoEuqv57W5yHGWVizi9fM5jVeXG+ilbdBrSLsWAZ0M2uWGonqN
TCtVbf3VqPzPIpwsvgcnEPVVBCHmVlFbQkDEA8QpTxmgYtakkbe0xFhlF4ghIEzs
CNszO0iHnquC4UpJUedMHnn5YaZ7iOhlWs/payVV4Ib1iZ3cs/qXSFl3eVW2ki2t
iMXX865y7Tmax/f6DtOjrlCK6NbaW8+d2cN0LiylQsQE2jLBC1hp5foTxK5BNo7O
uU6QfjZbCnSChAobgadSwI9HkfUnRwknuM63VdkTrJvF33QHukJth+5rGlgNYcAy
8akht3td0QpB095UqpEByE8Sr8Lhf+R/ZQBwrASapGLVEzJsUYpQ7e9YxY9Q2r5m
CJzj+7mfDgJktbY8Jdt9tBeVhD6KPyPgUQ8yszZoMmSPRNfURjRqTk6/ApljlQcQ
GQcmvvWCeT1Es+n+j+pkj5jxM+OLRf7Qfr0Dkv4tIInUuAzOdA5NbHwBXawuI3DA
TQDzZjYe5zEXs0OLjBS08M7LyVEC2CpCB8TfLLsNUgFbwza2xhcg0VBk8OgjuZ5d
TuRzgGpZXS8l+UZRJt2Aug5e7DGJYF5BMMXPNz45WM+9GiW04jnSgdlqa14tR58e
/I3I+dSXnInAYavOePeHXQxLdT5HIdjnDjJYsbdZSMvFtQXViBnunp0/B0WOsGfy
RpPyWx6IUvAIuAGhLFNGSJNb/rOanym3sqYwkbixY15EzZxmtiMQOCKf4CufBFls
zqlyg5mJWpntzkoQzB0grEMvGluUorZm4nVgy19Q58ucRA5xYkBucoeKkXBmni42
Tf4e3iiC7exhTLdT4/VZRHkFTUI93HIP8erqNZzXg/1wufACqf/X/qcwCdwParSv
EYV6Ypg0Xk7bO89ZfgMgyvNHCaHmWTHCwIy+Ugzs/CSH8QJWhmG5n/qxvkM4Nrz4
Jyk3BTuk3bb5wg+/gYQPyo75k4/jTAIDoHgHs9xbM/wWVaebW875OlbRX0HbQ+Tn
Uw9ojzUsgPQoLH+c81KJEhl4rt/C/vmv/MjFggji3fOKAKiQTBZcpfRY7wH0xLfN
NrDHQdQfUwalnTy+LAovl5GR8pkEhsBvNB+nbIc9invgtU5G2NmmBN+9Rdu+acpr
VG/ge4MLeLjVS7Jczneecmd1+zj496CoD91A66rxHJP4zXp+HPALXKM0rV5kWyQS
YxiKJwkXYmZ0gnvNuuaPi/PbG3XKgl2kk+w0gKXYaA2I4vh0t0PcHOGuv/QIZ+IX
gpJnmAlmIk9wXP7GerQ54WNNoOBWlE5Jk1/0JROPWEMI6WW0toYimWVCirEwJio7
WEReytLI07NQC2L9knHIQI+RZyuCLrTw43btAvAGRrGiSpbJbgCOAL7P75w+loL4
R/9cEgIUnUcql+vgjZxLVQdzS4XxLo+TKVESz1aod8hkhHXWa20/eNE4I2GXc/dr
yjpxKtIeLBOU+4VT4kZXQyCC0c34ltsoV9MzcFhHfVdVQvLjvLSaH9K3TXNkjNDM
s9vNwhu+WiroUtsdq/VCwdIUW6L1cq5/xPHQadFnuNrB/xCc8K2tkcB3EJsWgo+M
kPtrso7yjNMSz8n9L/8yQXY+nQXZm5LYVWYN4cHk4VUD00vWrQOhbJTK+AOQsAUa
/2NLo5ypmx3sZYFo2BU/uptGHlWUDSmX18IUU1JhmbrREknSxd4QjmfbjfP3NI3v
pCDw6W5W9H01SMHw26viqT/duxLvKdLYOrkUx6dBXSquD5Q3wqqgmeAmKd16co01
o0h/aan8mP82sU2kukS8pkzqqFAPy3pAf+dI4bfPuoMCK9kDtWMwW+qfyleEz6tC
x3DqTW6hOEf7TQjf9xRvs6ai2C1oexhaL0f+ZOe++lMK/dq5SJbCUu1BHKKsQv/U
TtXjuqXfjIjkpY9zzLIiiE3JWSRaovoOD+GyoZhRzEeeYU8YYBBnAbu3rPHXK4KE
0pwWqrR/4toulRVrm+DCYeURU2r5umXVp1dMiFMWWxV6AOVrofOYYUPQbYqSqjvU
TFnDtyJfotDjV+dk42sj3wLUWlIGk4geBpoW8El5Kh2cVg2Z/OFUEHFhJXm5AwJa
TFdNoyR2IAcQJVke5JgISMFr1qJETT/KuYgBKyRmsFEydCRio6Poypsgf4kKlLKX
yIMhF0czMA37i7QtrralUbPItysO4DueOrObWW3qY3945LsSG6eFf8QYYJgqoBoQ
/qOmUnpyMnemcTD7zcsdVvVc/Sp8KGshXmoOoldak7gqVira86YFjMW+oCT75hEX
ywQN68AjXPXBVvgTA43kwrv3PQSImO6zIIf9N2nadfctE35tgewlrwDHlVPBobMQ
KbDfNFqfzlk7SI1SmSOkDmgo7udL5UJYi49+FUuGdEoELH3TjFMn7uBLxX/lN4QR
J/1pP8ZPqZtPqUHXP+nF22Hauqi5Gxth7eQNGLNIODndJGhqGujFQI6irSzWkaWG
lenSZUdnbJMEoqyqSXHQCw+lrmMPQmKl4L7E7AUPl4NVsfZLgz5l/ViMxO8oWypO
k0vJ3KcVvdAb1sr/i9ah3jfsnMZ9sS+gsXQ5qsWEhP+lbTwLgwhq6eDDQGw9ucv1
Tctar/8kryYd0dY36++cu0rzmglucj5ZbaCRzso2VQLrnYxggc13V+K7X9Kb3pec
AWJZEpqXcXbUxo1fy2+8qm49hZpT6S86ZJ09VCAGGWwX9HecRdMBZhl6eb8UfegA
uC+WrUU/CqLrXLlyxP26nRSz0mCdBcaFfivC6ZRvnDKSj8rFEse8yKzitxU3hdez
Pwu55RWp+XkzewN/UAv4d317iDB5w+pW4eQa7UhXRXjOUxWrhsMr2x6PvBmcjsD0
QrPWiDfLKIujBBvE1tKWDPBC4ni493DT9bn9SCWSmc1uL/X90ZTpp+a9+pZReJMn
RnSJ3QbNUKi77M0oUuSSlbRpa/UXp+g79G06mhTuptBbJY7YXPN1ysqtRSciMThK
dBXT9sztW967JQ6sjylReLqVzSTZpP526BCK/MwxKYjLG6zT8y0PnP9xyEm7C/BI
yGEHyAQVVkK6mjeKEWxXaEuQy0xE5KN63a4Jkv65QrhqAm0M/5ocjld7XSn5dEID
9xtzQMKdgWFEbMQr82f9cxQrtoGqZniJXimV33TZ0cTXUfaeqkdg7E2trQZedWKt
uNCd2rkfjyZNY57o63D9FlZczHpFvwPnuEHPB9hUBkBfCKgWaEx5JcB5LyMGcFrK
emwUQ4xlptexCXw+1u6u4LQ9BhSf867XIBseVUoqjPVD6RuaAYnYcZQQHuCAJiiQ
B9pW0AE14z0KQBCpoLrR4fcUI78g0meEabkECMAPdGmGTJKxHOPg3u4RG3o7PEOv
AMUybPL4+HX1ON07HvREybuWcsiXg5LbxEWc7YWdWP0uEz3v3U8NeEtWKHY4buwd
ahFf2HDDjN5EH9GRXzx9pOfNJa7peewdLPfWu+kU7S+p7QohARhOuy0g4dbhb5kz
QTcO25xrqNlG9nhkwF6mwTIgy9VxtGCBhYojl14LkaS0xht/zV3wTcSf6AAwuNPJ
OMhhidtsFtuwG/rh7C6QDmi5oT2QWTzGTGfyn2RRXto7u3ndYU+sYgISpzCzrVlk
8vQhTq+LFau2aQXAi23NHx3Q/tLIwGbuns+lzFrDG9jcCU1Bn29w3tuFsLYqtqts
C+40yN31KfJgv/FoLEmXXlMaq9PyhIX2zrreOTxQgCehw6COW+Y1pRu7owCl0XN1
L1DPHvKQJaL0F96d8hjrZO2TQYCMWwKk1lVPNZZnqvK6UCiI5hQZ0aFRm6s6OTCc
ohLOcNTlwudMy0pXYPYcWWDVH37kAxt7kuZBME4vOC2XfHcgZeAqwTPNhwpRemyn
MRePb3uo1OVH5hngQ7opJ8E0tsLa0en1h13DeiBgnHKd1CUybYO2hcLqIyGandVY
hHkA6Kh7KzsNvikUXN8GpmF4tAvhwfVaHgHu3AarPIU1jIdQpsk3lTj+/3JYHFqx
+Ns4vH43X8LFeOaGI9SnMyYhnonLqtEljZlOwWTpWDFmfOWatkM48Uy9Fuy2vZSq
hybjwgh2aj2TzPZdBKzqMR9IGHXViOYxgILDYecUT3i+Qbqx56/y0Be4gSllmHJK
FATPndIP8CwM621Ry12Jf+bZjms/41jkWh2krSDiNmpClx9sRd8M4i2J/5wtdO0w
5z/gbUU0XwxpY2piD5pHrA0+K/HNtuuO5MibqBBkbge0+DSfMfHoup8ZBt6FzzyE
lhEZBYj8wFWqDd7vt15pXK6dJfjHGNAreGLg84VSnLUrUEQnu85F46f8nK95qWle
EROhzAjXbzTo8C/WeqWqfrLtWxsdvEhpjk+suyPQXarcreRXmZvNRM5mCNivGz/k
T+4B9jtbLxQ7XQp6up53xa5z/kSwZtt7DFqCNwivV1Iu54C0mX3FniiZCZAH9m5F
UQU0ubbO3LllvucXSgAqW6vRpZlsZIEGWt39ysyc7FHW8LOPD40YyjYjHT3bLAH3
WyzpIUN5k91I++nc7ag5hL+RfjEOM9GS7GT2kdo0jc5VrwdX0uGouOJ201ZO9adz
ZFSatS/SVzA6Ad5t8Wc3/807CfEHGjIHpjRlDQQaJ34ToDL/dUt1quM8bMYiACZ7
9WRWBX8pfGQrYGN8KwO357Cyh6z8m/ovHQy4tIF77IEEAq/n3IWXGanZLO8P8W5r
EiiD+kt1jKVaOtz4/OhBz0VJj0aqrH/nRdyaV40Jx519xzHleg+7iz3IgpDSpi0C
6VLb/vUKK0ACgb+1zf86E00lwQQWtGRvkZWkl9fTmq96qO1fNnMHWq/F+amVAcFC
aTbwk1/JFdBbteyPNMxxPlN7DBo2MKu5BA72LHEuSWxhWv2G5FFaaxaGt+1OLpBp
FAWj94M/RSDQMWdD7R0J6zHAxAKXe4toZuf2F2USexz5193XY8jExrhWi0RTWPf3
7+EJEtDHP+PNNNu+XGKgMwCokNfI+BZQl6rqmMnXcrSL4ATH7zY27iPZSjnTi0/1
BXlINOalELNN+wjEKMNOsVNCoyBpzMO4aqlNV7gxnEni01sysGyizedkDXQpDK9F
FKAoJAbznKh2qa6MXd89X9wBi8c7HuK12RelaKozIWv1d7YCqxlUxDnkqt9SLWV6
e20zym4jVdjTKo8nxgCEaRZQEOAWKuZ+70awhOh9edDqoSGzkeHSu47hgd93NhPd
eRi3Cypb2qaeghs18sC0Rek53/zQLAktS43XzDEi8Yc3SPD6uXVw00DrRIiCI8VY
NtPwugknrDH7NZb6Q0D0MaCs0bcBYezkHS2YnJBWkcyOlrluN7zkqsf2cktzEf8x
YT3jW+6jgdDBWOJLocV9sLvm3wZeIlUPtIr7aBL0b7oMCRaPAsiSKNeDl5Ldfecy
+ved+/o5BXdujR5TMAtBXEjld1jvRz8dLuoIi5anhB1xuOuKi9+2QYoX1pNwxXJX
Rb0wL39BSSSYAUxFB0CKiS4gmeCoa6Kx33c1egNyPg3mWixysezl1UhMdUoP6DeS
sNF5JFPu1OJuUf2LI4bqYoRQSl4kG4E1yezb5XbUBF9x7Q03fej1XTwZTbHB+f2e
FLr9kF6il8kPstD2bUj2w4SBaTTYqgZACU6CCBchaAvsXXeOBpbTh1Nh2Btu/e2W
EP1/0ZoLsv3VC37CnC45hOCJZis/ORz3fpj/G1hBlTIRnin020r/0tIitNKWUd2y
Dy+822F4agh+CVxB+s85UCDBF32ZHL6Z69j7hZdavDC9EI34DucuqyFsa2M4K9Rl
39zX/UNscpuEtnh7crUe5jyy0qv7vPw/gw9lHrMhWorkpR+4BSIwuca3l1Bj1d9T
AYYELPQbiLRxG0+eRcUOK4viWOBnQC/PgM0+MYDQKLZNClnDd+Urb33ebwzy52ds
aTnM+YLZaYJUjgIIgJ/L2DdUymxT6SFiH2zNuhf6h2rMseRiKJFRcOvqqZ1HJ0+e
Ymp8A/FkZZiuTsCByTCiGdys1NzP/dYrIAWQw2kjwQhatz0VCjOWHycoo/b0T72L
KpwrUEk0LxYmrIwwpZsIA9tV9puXo1rc215aSIyJ1V9jgqfGovbqmLT951EG7/XJ
/NC3+q8+HAN0UTatolpv+crIhCQwpEHTpT0ui8Eo6+gA3C/jTLTYtVPZSEAp4gF4
Aly/JZH2sS5qN5fz6SSltD6X7P1akGUGwsVhhEaPB0IqqsMc7SEiLH/3PPCZcK+a
XobeSCqg+Jx9jpXWM4qM6AL+gWSFmFP1xtB1ICyFAq5UXVsN61URiRhSVq9ESMC1
TTrln0LA5p1lHA7VTtPtmDghfpjRR7tn+73jwljAb6PZvX/0EQBBYAN84s+s8Luj
UfN1U9a+SIIzjlI9eWGctdl/u9IFRCH4lWH8UZ0k+uOg0mVf44WJVD33nHUE/t1p
ZCEwfGgWgtPsRd3iW1HWuKcw4uD0B7qt+yduud0i9OdgbJJpb5dC38lAjGEanLh2
dA5MX5IGhdHf7iq1rj1BFWvVN/U1BMoE+3sDVElfg/FRCMPt4eMAUMG9FUoHzPhU
YttYbpR2egC680MNM4hT8OcDkj1i4KAOnhjtRcaDhSXCYIRLtWS80mqMkOGbtwke
Ei4QTbipWRDQh7cM6XAVHBXQsEZ4eXxRa+wCNt31o8lqCS3wRorUTMB5MomvmlkE
O5daPL1njZ8vYjCU+U8SWgfilm2AbmfvN94KiFrF9YFlA8DeLunFwvQ263kTaTCW
8X32Wb+3d1wwBMfN61FRqiyUQqEGRWQr947L283GL1Yrh+z7V1eCuxufWmaNW7XN
ASrWiu2RDW52VQJ5NJvvS6NZDM6AxgMwKSGSbDZf59uXTOaCz4cVwZN8RuJuIWrm
p2rojzXhzgysMeHwPyw453BfrpG+DFFElcAjV3Z4WnWPTMhZCGc0TvFq9x7qwajV
5/XaMIxwnNYy11BTtYcAeMFT4Cd6ZJNpTm44M3UdFRL5SDtrMbW37QluRushEqEQ
qwAKdmoFdaTIU2QwNTAq8rgV3EFiUMf41ug7iPjV1+9ljRxkxloaGdVfgMRFHXfc
1K8BX8tBfL0+ESJ2VHtPCoye/2lpSyaglovlAL9bo3VPlly33uThhCvYih6gWeNb
vBn8543hufsI80d8iyLklPzjE0SY3M95xLkq396I3b/ujMJ1/7NUeqLJVBMiCR0h
5gZEtn489uodkhydRMo/ZNZUcg0NYo576bC7pM0rgUxByP5oPSXRSK4c6EvZvlnc
y/D8nGjOrN+B8EVAKvg+erx5SAPKAOP1TyeJwxj7BCP+OMCzr69/c6aCRrLaFCeB
Mcky1FkY40HTGl21cuVWulJzLftI9+Gov4FMmvO7/QMCMJLuI1bBT0xIUqnZQVQT
xsG6129UnKHsdYiGyuSMMLOx0uEWP4KlsoBatDVVI7CVl1c8it8iJeI6OBgyoxW/
LZJ8BI2ulcQQNDkUOxJKHeooq4nMboGAtTxZhI15OHLdAbwkpLFeFMu7tGQ+GfeA
F/k20CIZ+vl0M13g8kWs4eEuHvKw9JmAM0n/oiwhFvvLgiLyjkg8jjoS+baGecqG
R9K/agb1bbqBDsuIKHmghNLjfNfHl9d+KenPCbM+XH8XTRBEvC+ee+WoX3OtE6Qp
iRbgJE8OvT9D1XxHGH/7SkPN8ES3AC13f1hnbho02NnwQ1w36vObT7sZ7sMVmugq
8JzP2uhZ/PA5zUifKMoD0Hd2bASGWpWkGqUj8Md/sqqMda9zcHaLmRTDoXCXBUlp
W9kcUVxrCm3e5yaaLQPeUCulFBjhFSIdHmv3pHfYhOYziXq/Y3BaJsNepRHERalR
UhqmO37FajnOsO2g0cJL//1Ac3W9XA7w91+f4kO6Kq4Fsj0drO6lfcR27NvwLIqt
TcQh3aPlLcYQOfweaE7PrTwbbyntywDZEjYpYLu99EjiGNgfhaLB6f6Yt5NJBCI0
G7CHGdj8IVnbpq16vSW1u72A3f3SId9AQHzJe7JZ6yZATstuseJoQ8f5EwmelN78
Yp/pmadTeWw/AAXdBwVIVD8OckwAuKsu5zqTkG+gQ2pWa2RRM+1FnpIe9D703wet
pz3s+ij61i/jVUgXlteZkraf9hbAqiAPptu7baMlU3ny3V7czhPCoKqiI85gRlKD
ernqyUTRM2sCh6jLJ1KN9metkq45mI50mdP8GzTO79yyFolM5QBfuG7m0Uh1CF4m
bQdHWMPCcjnFDcqVYes8BuxdIJtpIJ9D+p1KHHqAUPwAeIQcMixdRuOJnVNaxUYN
BsKGSmiJkdOzOSaV0mNl9dTb36Bn0ZEZVgsCM2QaQMySWA/u16Zd15fdUU67USvR
4OaqPcPcRE1S1IAf+rzBT9U8UZiAHCVYSg2OV3EXX92yOyq6E0yileMcf015Pdve
oOodZurObhLgYQum9c8r5rlsFUwe3eFTJUfsMwmtpl/styObv5hdNjYUxzRi89CV
ddkUDBSZtaljPsWkVVr19ivYKg/xXiuTjpWyZGN99E79z5wIrJKGGS+dC+kASeqW
7KHelYrWYHAPuxZUqkoRNZ5w9e4PwN9JX5rvSbe5pjEU+npfdrMggmX4YSX2aN3C
FSFyRmtD9RC90ksJ0aqEVZL4hnpKol+zMkVETo3+7LILEuHZMBpTNqoel/tKkmK7
EuU5SIDKlCyISW37C64lc0dYGRjL/BGgpS6+A4ak3j+bH3Z9YKo/9DQTt/FyGrdA
INAo7riWUzu4zEa90mNCR7is8f4vZUviNz46NaFadhq1XTO/jZgTEql4O0OL1ZVp
bazP4eBeInohGAHayAiodTf0tnnd8S4JC0KTaqn1sq5SWuf9V2ftEXCi8tAK0cC2
7xZ8Ind7FbYoSlUtdajvQGo02iQ7JHbJqPh32sOMVYk1F9ZGg8/Qo0PPzCSIEZ8a
mBXAGnZfXwJ/dgQOAIJB0kqb+sA5TySytt/UXmo+ev7rLT/r9qM0uvAzyG51GjAP
uOxzokm7jS2mrAgGAnpGriZ2MNhzh11W+/LmNQAZSrBKdDNUBVIXZX+SJTcAQZzG
iUyeiToFtIDZaEF3kAbchY6tHoQIOjZxli9v5t3ogOKmrrLiaQbA7m9Tf+h72+Bq
Z6/CNJvIJ7bxyCztOVQvZ6/0zN/r5k31QXQ53bQhb71iWL7LVC8ZD8FVBA8O63sa
b2oNvlHtr9ZemRG5eG6ULVCIHS/UooUtDiNyeroMaXBh48SVWlJEdESsXLnTWYaj
QBxmR1oqq5oI/bVow9QcfEQqV80gW9TKzRsMXkfU2QMjMIO1gqdpKGzUjG5YJXyA
oOQeV3zKHaj7EnuzGvfOodlC0OXh2zpIBhcjJdZPHycFxOlL6CrbaXXQqLgjpNQu
2iT70GyOA3XFFXKv/izMGi+HPVT+m2718loFJVzO6wJ+xyGnToqjyI6MsLMhMX1b
rf7QS0aTkis6gFPdFaCNg3DkMutGmcousoa+83Gz7IsrYT0TZj/n21MdX96xTsYH
jRMDu+6h3AU8rUQj9RxDicSleSxwJG7BVwG5hjRH0DZi73rbMGoF8312bmyUNpw7
QGCNIqDF1VXLWA8NRSx4JTnNtvBF+DPTiQerP/kNummj1ISrtD08n+jW17tPaa8R
uebAIIhaV9UeL10uZ12+IdwBMqTmDvwohqPdCzwltE+2k/ZF2t24ZEOgEOHcYSTB
VxQ34LH3853m2BKCTv/mgvZPYPQsjW5nCpIUf38wwdlWxb5llPOomGA3ykw77t4J
yvPxSRypMQqH6XM2JFgLKKPPdbLGno4ObcaxeUCj1NuXNLchsuI/UDSOgOo+jPR0
Th21P9ZLN52TSO3YU0MATbSVq1i5NuQGuOXN12cYx7MzSmz6lCzyYhRH+eit9FVu
wpZvHQZ31VlZWGtj6ZjYgiB4S1W7L1wXukXv81T+Ih34RSnBSfIvxH0vxwHpjXl1
TFgNmc4TWwtOTN+1ScYLuXq2dzgbI0XgSh2pC4U44b+l6TMjr4Oaft7twmJLsiA+
Av9j+uylzx3mTBjolCrQdsxVFfrsyoJUbHa1s1vjdIxDNgmGAVSr4Tjh8M7C+soq
VG8WTdOuXT9bbj165j4epCIbbjIZAJBrTvX64uqZ7NGPebqowGJ/Ykmqgg7UPUur
U8id7djCZ4uMSXgD2jKhvCfH8mMXXKyWWPTgY9pZw0Lwv+dHXzb0FTY/OPJrv52P
bw5+MeN71uoN0O9vI/W26b/m4hjMlT+Rhob7p+NAf97SOrnvlXeiQ/pjAjWG6b2Z
PyXE2If3kfnbkjatu6mRTRdJi9RNRqGxxMNWdFImkt2w2JRntoLMlpSe4iX7fScZ
zHdZYOwAKiLUvj3MJgRIbuJJZtORO8ZnP97AHOoCCE2o30awv3zONmMoauAIEuyE
Sxd8B2J7qLmg3roO5M0W3WT7AN2PWW0qra9xNGXbxkIaka6DoFy8G5CUVvFArbHG
M/NfLrGcmshOi+BK4cBW9O01tZgRiGNqp4zjKwX6hKyxEWqlttL8nkI9veW3eikY
ZE/tx74QVElXL+02Y3+r7iTLwA1o+A1xMZ9yhWu/3OVIvaxhhfj2pv/nygs798/t
CNKLhrJfeuI+oeBexxUwQmqE2giBRv00NVMG6ZGoU4TXop96IEvuhqzIj1Z1XfbX
gAdL5Yc9xLHz7Vx9/CyoMk+VIsgHU4ORFG/aeOBsoUCyEy17osJllpcbrZD7WzdR
ZqRv8ELKC/MXuoubdOJpmJBfGTMza+h58eIiYe5yPyx459O+fsjMVOcjlUMcmfAN
TwigDfWrS6+p+b0FwU8W7/eTAsPkO0w4uuI6cmJ3M1fkNM2u5Yew11/tFHZbuNyc
nmbyMjkrTSP3sifaMYoguAAHWcTItp1dFaLDxuoLTTtSnpEPYajPtIreHf5Z46qy
eSPWFXM6g48x5DvgHE+fZQQebcPPmnbBTa2F32881ERHmhmm90YATCDUt6FliSrv
Y6ksUr3kL6IapoG8icG30ZU53jrZehwxtzQ45eGE26Wd0SvZVRHfS615Us57mv4/
n8Y2etI1ps8Lht6txGrn3yZpN8jqbWwQYq9fT4t2DpbTIzLp3wTbF+14fg4hWd8V
Gs9LH8adyFEPTY7g82qyG96aWIDmMSjgKr6Q5x7s/MelzBUNz29D8UZXhEIPmvcb
pZGCoW0qtpogrBg5s7pioBq8NsfusFi/O1G2/lhYO6OBFnojNXbyWi72lceN1zt1
tfIzZPAZfgHqzORQ2ddJwOaMeFbdicFY0aZigdLIi0Xd9hV1+wlYR74PZv5A7eh1
nnrSNgO8nHU6hESTVJoT8F8GZ6YSokBzKMDcq/KCTQ5TTy7ZfghfEX2hoP9YXMFX
qwdOw/5TfK3eBl2wFNRO6ktn23GwHOWAGwWWkd3Wclp7KYZNB/wn20gBmstatga3
GDPLUNdhU1nMCoK0+CTFkjZRgQWluVaso3ELYLkVWzXrxde/16v6yXx4Q4rq7qWO
C0TY0kr3pX85kT9Tuvllis1iMyzzPsjf0NYj0lgbFns1HUEYdXT/Y+5MojpiZbNh
479jGHdCDjL0jh11PdqcjvAAy4a2uPw6j4sVP1c5Msmyc+EBEja3Uo46VUTzPitA
xZtWSFh2pVIPCJQIT+5QQ+MotQGqgD6SUOYD5WlTQLobbjxr1W2rYXfLYllIKTfh
8IexsptKabuhWuZYe4pFAhzQpUHc4ZEVe2C8GquD937kEj3gmjO4vSIIwFPEkYwR
yckdm0VejKy7+xyqNavegP6nJCsr0LeIrP4CuPNlHRwjwSR4lCDQ1ncqCa2OY9fK
5gRHcJqPUPXztqsFmwWAVrT9C8tirv3PCWkMvMnmgz1WuiPL8Bnp5HLbB4QHRDGr
eqnqWOmV81GM7D+JhYlsWD0L5fW+JZVnQjHZDySBqdaDTEfs7yynWDnAmlemJpP5
hlVSIXCDQLFPW3H9voPATJazKHKaQk2Jea9ywd9G8xLxjLwiYcKkptfNBNhMYTAm
7bQXM+cYgLTXboqdMiIGo3uBiUKs69NhcZTE3hsjetI2FOD55NOvhvA/Wo/5Up+4
Nh/30w/b3bgEuMdKssaR8bij5FJIAoDZg7bzNUfn99h+y1QI5pY+0YlhILLq/IxZ
fPkFkuWQDi7z/Yn6I91hOL/4JmGsM1RM+uAbJWzasd7VTA3fI6IzNsNsDisRjj1N
syoD2jjjsNcTMBq+c4jVESbrJBwHt5jdnv+VNC4/qdf7GZfWCjR5HGKH1TSEuUXt
hByx/5Whyf/+wk2HCsR0Ohgmp5RPoJnKE4RUg0NunVtfhe/4uvGtsaApr847GYEB
7qbZ4FHYCSQBiCCbYe1qzyd1/WlPA+eQphuFZ/iPygoatHSrIAzJ15rd0PQilkRl
Qn5lc6bu9IElhgH28S7ucJLJcmRa1LitY886hnnaNkOaRJmby1WLju7M+1Vc6+mg
sjec6h9SjK+cqjpa9i/dOkupFP7kQq++MLCyd3lijRHnWlXXvDZ+gzh6nTHrkK68
d9hBm+PV7Ia0vR3ijMiPElW0x6q+faj1Cl7AIEwcEH1BUYqqIect+hIzjzfqRrS8
jzonxcRqFGTPfQkBD1SmLCOldu8GeOh343Fp8uzEggnp8KmUBwNAF7gZVLvKRxre
dx0rljd0vDSOPU7ve+yLk7sKxCQyq4RwoKO1+mHxdoZuDpWI93XiPA+JI+4NCdvt
bWX41n6qykxgBpHqVJrWICpCUiEx+z1Nv2na/WrYXPab/weIDs1BeOYVmfLzN/iE
Um+xSsIc9FB4dwR+68vE+kHiAa3q6hVSlPY8ClcZicDVVqKH3hggy+Jgc4wRvXJm
x2yQ6kM21B/Cn2y4yfk+MWR3HzsgP/wRyR/qXTr8PeurPlE/cbQ6e47RRDvgeLXg
aCwF0mLw8Py308MHwECSTjFG8YGperX3VjBRhBPryhFAAKkwx8fX2pnHdQlytqGh
LDpqhCL171a7tqMPs6b4fIS71RJvTYJUvsLyBB8+rVL+64rT/MRhG2XF+dlKfMRp
8xoIDANF/rZD9LTkLTpUCsTpJDLygsPp0BNA3uwbeLXgdjLguP72O0Hf3uQAp/4Y
MKx+LfJQG+hMELPfVHOyJ7JYSkKrD5guUnDp1YWRxc/lxGsqv/2Tmw1VMEwTFlxr
e2a1FV4ig+TmMGkzzZTHs9xs443iifSyyMnzmp58r+LDXuH0nyFvHiM/vL4tQXAO
o3OciGnc5F+m1OmJJQgKLBsgVYYjXniWoRId3FTDnc5a40H/r/AJ6+sGeBqmvCZ9
Xg3IYJxi2drUqeUz6FOuzlc0sL/GLtXlNlVkOPoksESf4jxl9o6LUBvGXcBEifwm
jIZWMoUfcQRA/NezOzKDnk2V5aRIQKTaxmNB66JmuVMx0RdQ/E3LAfKZD5izuQDT
aJhXgNHtFypbKNgKZgpWwwuF4CG4jyy/txO3h+6jK0eDdaEUAleJNXKw/3Fq+KZB
fclX95CiRccV/YtAzAvX8pVKZU2W5DPgV2YDURUvy1iF+OksXYFCSIz8AHE9dvsB
NGP/ml9VmR8ByVLtfDUZ+6SCo+kL5D5t8D+FQw7TQPgMelUNUukBej+29o7XlPKE
hQA6KfCPskQqGjp+wvMFHrtRFy/WkB/rP88hCSqewRz0wcACP5J1rmLSoHa7ECD4
O/85U+EyDRea6kSmXggLS1+pPsh6dW3+6mjpq5+mZqIuqmrWsqSMIlItjSz4l1C+
Ucw7aIoHqCFowlN3HVsm+zbITh6FkKauB8neVprYiwat/npFG2uTNdxCII6XXrcP
R5/nQzdtmvi0YEN8/qF0zJfQrTrOptF7pHwfetWhbKqV813mdzrXvEoDTobSuR3X
CknsgR8oSzmz2NptqKtTwZO5LyebfpiwSqfq0w9EDIs6VaxP71eg5RW00avjMrjV
6oGLnGTtOMiLOgEMI7IU9HRwupUwvH8+2X9X2+3SrDTuftgcDBALMEToPtJnmenr
JdJuBnX3dW2Oej2BEBw0SflWmq/Wfm3H4rNQCWdO2IFGJF90NCPLVP36UsjeGlmN
RINxvEjyn7OZwq1s035lPrdcNPuuA/5Gd/1aTLLEB28c3nhRYwegpz5nxa4vSaDH
1vqNQGYhoLxNhK2CA0t1pAw9Y6VKJqm20ZvULU5isxpNBgjy9Gc7/4CKeucnynGX
Mj7DS93h7pJfVLPrbj9B4bbKdaHzxHf0MjAwRuEMfTiy+Gp+NGqwE5UNqhSfluAz
1AUMXQZDfSzldfMnqPIT7ZHyF8uK+JmSxZ22PNAHBwpfBqu04B2J8ISLrtRNMzXw
vzfiuc1p7HT1cU8arPa76mxdmx/Cz3jIBTrb0F6d9WxOLtcduIhiIqaZjJOvxV9/
h2VoVuijVmYJ2ni6yuFn5TGL92w7pI3JrurO5R7rBfBw6ddI5WSu5QqpDnpcICKV
meSo0Ks8v1rO2mortLF9jpajGEfFvF9O4OE+1Ha7ac7gLjjZj+4vliiiLRhAd+aF
xTuoOcW/3zyhod2qUhDTLg1nVe+1v2BhC3vPPn2IShP364vi5wkxizqXIn+89P78
XglSM6aDUdTIea3RPKdsDh0LkTn1Sbt3k4njWhP8NCv3FZ4C8GK5AIkjgnqlHjnB
w84Kh9uMSNbHb5vvpV9kn1ByOO5d3DI2+I97B2gSFvdrlj/xLyxUgmIH+alK7wr+
hoeWbKEWeLNrU9xQK182wNl2bu12BAASoVGvuj+GyvRZe93dh1nQRLpX6tIPkXhC
cDtWgh6SrXbyAa4ySA18H6PfMYAcC9LQzMLdpAui3YIatuQdZyaEWWY+djS1zPjy
Tl17ZtChMvaYnqKR34UA8EO76yDN0hIBi6HGWoFs0Armk0mtgS+AGBObdrCrCmGz
1gsAa3/Aq+/Es7AIsbN1GTIZAhCclZYB152QgQaWP2rEOtSqKNP4qMBg0vvzOic+
U4WB5smojiKybHMPs5/YTz9+WzCTCNWLlKYWHqs1zz77NmtW+fw6KN+iMK7X5x5x
Cytw3IKZIj33i6deLdEVT+/KdfdPoCKiJdy9AhNWh2U/yZgdnm8bLR/aY238ZMH0
XJLBzpFSXRNv5J3WneqtKlvVzrynIWaeuEPoZhIQnRBw62tfUHgl9SK/cNAVNNkD
+zOW5zDbTQGBLfP/Vn9gqm/coy9LlD3zm0IJZfvjNt7ReqSX7jztiqRIfJoccwt7
plgmve4c36dzSqXv2k+oZDeKTaugUmJwkXD7Z7vpe4QV8KLY6nbAUO6NwdTeeKSc
CmTKmOQ+BsFctNYFdOI8ziZNmyh6FyCXPX3mHTyK+tYs94MQ4aD/GfTRh9AvsLJe
Nmiiz0JginSVY2K9hbiRl1kaa+pjz95bIQ9EV+BHDvUdINBAhY0a0m4cKfPUcw2/
wB+uzD8dLh4owBcPAsMR8uoLIFj0R77sYXsBH7KO4FxT2dTH0SkSjGk5JqQMnVe/
2N7s82/RpG2MQ+EtMjsXMcGObpcXfteskcHIJytRf14yCfCS3HyFEpOL6s57uK32
Ew+Sy/2mzojFXVw4vHJfnGtx2G8OIE9ZYmQBVMPBHrndYNU16oYzYID4zSk13d+V
dK3Z0OUfSG26IE+fySE/jL5W3w0jDVvdVJSsHpKU6CAcKcqa8mq55hmBKLlu2izp
whBALj8IyJ8RZADroccGkJDoE7iKYDK+H6XSJZDBVQuDBQvV3v/93bEJEXoWVrcb
bwCGDkRDxySFU7xvnk6t4RkUOpLLO+wpK9cxMsJgtPrjjpJFdC804N4vhw/K5pBA
9jfoq3tR3axoZtvzIs/7zjDjrN+gWZjtLMjxkI7XkPhzQKTAs9XXe5zGXrkctLDc
NUsW2+0RS9CJ2rjSGDJIyNhBO9QUzS72MAmcRfztmt/7K9d2iBqT933PFC1x0XKI
P0YWPcuvkzuuKavPgDt0qL12+0wRpluNJW2yiRYoYdOe4it1j1YQIlqFfE9ATJAo
WwrSDuSA5vIpjvyhUVEJhiVCNOkh8BJNDt0oAazIWq5yfMYFrQv2BDtyQC1sG5tT
S6DoJlF7LGz9lm4H/tZfum0iFjP0EiXh6u8Y/LPO4DquaiVJo46rSvUvbw6sh5VG
RCg8tspwENfGGJna8gZPAQyjiWD5aHMr+oCcP4tgcw7WFJiMbtfNnV+daQrT2EQk
flbaRHadcVLN9dFVQx7AlHVDnIhFDIqnUGqnr2UXxF4s5rfx6FMHA+4hmyMZfDt7
3/GelygnW7iqDK3D7Ncww/q+b7KYmJ+wyQt/tAqaFli5TvoMu1NGzaOvPJ3YvvuM
lhb5wRf3oGy7BfEftAbTy9HBb8R4x4x1smRpj3a027osxbLMYVIVfCx963Tlst2v
4QHHajVH+n7wwc5f2ssd005aX4miO0SWUcGiGD5Dw6nnAlp4drcRg5kE7HnA9K49
t6vc2cRrS4zNy5ehyrgSu2Z828hEgNgRfK+pJ800l7BGjsSJ+S7cfVYNFkiIROl5
2wXjfcGrA9n1y0DhXpJ+DJQNPcdkxW47ATX1TDfeh9PMHK++hNe6fDhCVtgE42Yu
6OTQa+LpbsSGiHW9uSobG7Rrri4ry53H+/i4mEPEdDXF/GQ3ucNzbR6VnpwspXQw
Pfa/eLjX967deFOotgVT2sIB9yBUmQAI4HVmSaBLEJJG0842dCT+aKKkt+qOVaef
8LC0cg5/mZhcHTyf2/kKwwlKjDaKu5hKpUGWnvdtpBAnexnAO4aS7VEdomgDM43i
/cMf8jndBWGXqtj08s56JhYQOOgPxOh6D4prERvc4xEVIPQG7wIBCWkWfc+Yi5GP
zjVQKekBucCyKAStUhdbusuQqtYgxQEC+C5KvgWI7OU9rxaBoNoW+q/DaxJGqvt/
1/B80sVBixdN+8cJBQNA3XeqcTQWKK+znJhWQTZr9+VrxXKwgU2mNIOcITYg1gjQ
cJfor4zP9dAEIZY6DjiEVdUSP/z8jorJWUcHFsblYAZB/BXDrKtX8xW7AwUJ6Yxk
MKym0Hm0pRYkkoJ0lq7PSpL/ljIvjI5YPrh4+vzbJ0dD7tMp9rg7oRfA8jFCkoMt
obOjDN9FHxeHuPbC3k7ZHltH9Dco/XSdq130i+Rh6UlouvjwUOUS2nuioiXqR80p
CPB/DQ748vEbC/U5TYAbwpguf7HoDUx3XxoP8bpkJPVkGCMuQuYCncWli1kBz/t4
JxKJG8DYPFCI9NlXEi59KtBCG+FCmq8zrkoflmjBhGGOatFAKlD8/2ZLkWKRG1Xp
81zYVm+swz0iWlnMvFUEdKCrCbMHfWzr/winRB4kEgMJzwMQxg0F9KV+UYSy3W8O
scvR8rUaEJfKFFzHXKXcIVfTj00RplLcTNkmWy98t+CWwc4UpbuTsWIOKW8sGwWI
yXa+MklWq96PFw7ITxvgH/J8CkrXyO3RsnhEHYS4d2Zt5klOE+iWorc6q8/Xhs2T
ib9OMeO6DAk0175uecvaBjP9Q08pHmNB0NcPBlO35jawopy0/8LwRTQ5fy+oZxNs
nVFf1YOYTl/7WiHPfBYv5jP3VSNTW79jAQa3xHpLZ9NVgZsgXVjJvoShRJKIvfU3
93hN5pw+ZmYu7sXLzI7le/yQf1Szgqxw/Ia3EoYNUaV5hy19OsOHzwsYZeYqxZNL
O5IikrOnpgcqioJ+u3spt0JJhbBinT86FCIWGex2L06K1gES91JTB7OVQbwjGLNJ
bi/CcU/DQ9f2oKhdy3DjGWnIoP6A602apMARIHXOnbzq1fQBF+NkHgVndqSiEIT0
FSR0+Hl3Sgz1pmL23yP4AOGdgrQ4wAMBQq/tuetZXAyTug+SDuptyVRL0oK9Y2kf
cIkVQZoweAgSjUCJX9MdeaaIVvTFoqD/L1hm3HrycaRMEH0MTHbSf5pUbuFkZU9U
QfJk9+D0sf0Wx3kKRUKLagRnWejZJzEvFV7aVb+ADw6p+eHWRblodE3hfz62lz1+
gvlXqyL1Y4lfrG6/LK2Lgs6NxmksQIUDGLRtrVgd/FqpNbWZDKcVKM70erbD6L0K
pgzzMr+63e+krKQTf9xBYDubud+d9eQul2k9D9SvmCfveffDmvy4/4UFJLiC1YW1
UERHxZFtF5zMESRHW1tqucNVEFWVGnGbsT3pFGnD4AAXmC3WOdYfTzkx57gOmedQ
9rsYSU2we0ewTYSl+G+GIP4YXKOuqf9/Pafe4XQhVLoyk7pvDUL5yhRaMHngdR+z
MVtPd6osT0FJNVwZ/Incng494OGHXakrqthmfVOG0glB96xPD1IK0vmp//KDT/u5
k2Xf1amJRWE+CZGzH5fah4bKbHjveTuXOui7ZBVw4Iwhta8kNOFCK3uxY/CPrVgF
BEPEUAaUrFVkeRc0knmJ+UxdiqYvGjIhShnr3i1x7URn/mUUMDnntsUOhzuG4aqg
ToYvgP/BXwTSjqKk7MoJJ91/MdEL2tT2Gp2kDeE+MmcXboUMOaclzQWsC8V2ansr
HDIgvHVRSSpPBs59yL356r0v0GmdpNjnZDUHVxb91pc5EAHvObN+KCzYfRD/D/6+
yox9r319VGxzyWCwTN600s4kA/fmZTlegSiyQRD+tNQcEzgCFwK3LA5ncFYRnlpp
z5KYJKUIC4Y24Qo+lVtFwdnac4MYmeSvpTy/jzlfMiB0cgvg3WAHVlE0sWg5TGq2
r9MnmlzGrihdsM2lyuAs5NRzWY16PfNT+z6hyLS21SNyFsHkbOXVoGrS2dyliLRf
81tMx7dANqur2KwzsHe8Qyt0BmpwlMclqkpOmULMgZGVYFwFfNfeTA+lhsAJznEF
/82BgdXZ0Q5ksUg+BVeoFwTL2k6g6MXjWi85cKMC9g+jwMCsAn0KG3xJxIchR7ff
ercVzd4j1pLgIMrjGp1cTAlhx5Mpu6+t5ShpByg9vsGKmLqfBDm8IAzTZQmLJzXT
5B9hTPZZzwLDrEHzKFQx+S7+ujwVfpKsKlN9hhHnv5Qj9LHc2qA93lnh8UL18cwg
VbCEtOJu9JZbtdOBLw8dOUorF3W8zXRV2wsomqaNtyacSlEkkmKNYdt0AbfKto+b
DUEFGpkzmZAUrZtjk5ThbUF/l2UUUugS7msIv+u0c6r8zgisSVNzgEQSMAYrda6e
kGJlVq3jpDG+ng9KWKU44+X6OncUes/iPRSDySybACSjx32pWhX1UsD2gGhF4avx
1YnijrJdJsQ+2yHP5DPrmPKhMUG12ZKWbsICI+hjZi/UhcI4LBBFiF7hJ0opS9MM
Bm+1Q+aLi8vsUKJEyELTY/Thj7pc1+AekYz8byR/Q4RjO/vUReZ80k3svEKfimp2
qF/2w3GyDMiweSoO6Q18kQhP1ZkXNTwoi0f3Qm5a7Q/UWLQzh3HWumb65TOeNw3n
lKrWEs20j9rBvvT86pY7SDGCWqQvqmS9vxK8HSz2m1byMgio7j09nL7Ld11cs6TO
WBo/YCGN7L7OuXA1ojsVhmxxKPwvey4BFprmigkeGvMekStTHN/lyV38NuW5AV0D
VqB5tO4tg+wlUd+e8g7GKMEoo3GXKSOvS2FUGV/H2ZJnsLsoCbb+EByjcZkDeEZY
vkklv9jlQvTdbxKqSixqZD+BQtkmaSBBarP8VyOqJ/a2CSYhJoC3zlWR4wNQGBjT
clrwiK06SvI6zckDT/dYv9ni5NpGQkHHoUXHFYXC7VqjwRgFH/rRys9K9SBSXAGx
RLbyYBob/qNwVtzh7xYuVcySJI6v6aYa0cxUBWNjijfvZar3kLoSZmzBq9RHpOH1
nrodGCLDtbhAjR/3yjywpry/O4babmsyq1CsFxHBvdSU3KnYEEBiAl5kQCeuRIMg
kHYtbb0qYyvt2HmRyzpMc4smNjmwGx5aIDC9TMkSWtpH3Gt42fGtYWnjCiZsqffn
y5OM/oe9OnS/jQ6M3iea9ZvGEeQY1U2z2eP014Ym+n97NX0Ho5PGRwgsukP7b33v
tT/JyzhQFVeSzvjDnD6qzmJzd4fdsNGQ9JAGK4ZCQJFNdj/O8xkuuVbewEiOq6TX
1yJ0iyFNG7NEpa/oUSPMkRCzt1qiNMwQIMOcsKPznC26Jtjn7sdlV0SX0TjDymqq
gboNegBycTPhF3yPV/PlBiV0/rDp1squ1eBYhU1fuqSYwPWeJ3k7bSYifTWEKKOa
UFvMjLT/Q8RL9Yj/CaIbZjgBk1nQ2wTIpBVtxEVQe966g+xH3DoC1r5XsIxzrVjD
PNMFNZAXcvVcanYhskEFtR+O1yUpQJ2s9qi2+LIbyJ2LeoLJzCfQrqi9oi/StifD
8sMneOegyrAUyhVd3JnYrxkyWhfJRi8cbA3t++eHBZMBU1lEFbvx3539/k1XJsqC
UhTDXiqmrE7SNWpyBRUnVbDmKXn3YreqN6iB583zLfkns3H1MoXxUvUXyFUeofvb
OpZPZnD/ayNDyD/UGvFlIvm6ocRMbBa3Hp3lQZbrNEr2B/jSSNVQT3KD9GsbTlmK
pcBZmRwtyvW9m1XhOGcU9FaF/ft/YptqUYHIR8t5W53ZskGGN7HQQdPdJTjaG0Uv
zHsm+v1U44Khw9PU3x5rOqBHCOAC2DyvAhyzDLGPwY67WCjE5byLF06hQX3VVPdZ
XYNklR9DS9+D8H8Jf5IUXX4qgjko6VBVkByt64gECDMcDnWRGgsKqKNnFmeJ0T6S
cntd920vkhLxv6fpaBAzBgPR4pw2K/XsqWK0Q0dmRBdBejmXwQPkHsuqQ9XmI4cN
NGquzXXS7gE5SXyRKXOFCIBTc4/gAkCOg3oVZGOukw/ZP0vKns7VdDOvNwqb/9ZE
zV+fO0AbvcZ47GXEfhxL3SSBbjVfOKRcsp8lZyyxdltrpIhD/16BNwwWQgslplle
OTE0+F5I0WyU2+l1HReglRvMdLCUAOnOYeOA9bS5HIa4tHSCSS+oAwTGNSDO6rbE
pSYH5fcuuX/ZQndzPB6jCgleH5rVVaxJBqKSDkFkJ3hiTtsBK49IvtXOUWT0K1/+
tHJ4iOK1iHhInSnoC/X343Im+VUq3q3G+5pd/QUdnP4kKtWDPldl9ZyOv57rt3Mr
buToyfCpM+a2sBM8iiCCteUf6EWQAiOdRiCL4Tolngdp8fRMBpcxYWjrAojlrgIW
n3dmrhlxBzlonu72G1E2HKDktPlEP0Z/PYMbcPv0YWY9b6jbA6TOJP479FSHpBYI
+WOgMgCLzQ8IeID1HsXTKMIx3hhwFAVMUg/xBuMLdv+/DthDrcQJVjweWGFzJftQ
YFEi5f8AhtKPEt7d8Iw36OGoxzOF9QmdDM/h7AkLQYghVGvgEfbdX1tg2cFFhzM4
77ubNKQo9y7y7VOSbqHC5xepKaEr1mvgbWnlLIKJN8DUzSm7nBNy7hn/geugBeeH
VhvAV2JPxJVU1udWinDRz8jdXnz/hPDbpSBwuUl9JOMN8Z2cbfUlhAOdWIvTC3yi
XeGn1aNL2TJJfiyVgJpTLwNdGo68y43jDUiuh5lU9HQM1F5e2/xzufsBzUkkK5RI
cjHQVVvCufOc2aQIK7GqGU9jFV4U3oLjmRFd3nhMeyTu0/fGLziO2LGsPo0cQwl1
VJAGtq5wXpqF8c/4dFs9RUUJl1PsRNcPmN3dtC5mUtLmieHdZVhvFitPpZTJ6Pb6
J8B4AMXImyvNwPsYWiMEF1ZtXGJpIxPdzTbl/RsD5zrj0b4YLD/FrQ3IK6tZBtJ8
Wi0cICBpdvKHIHOaoGOFAhAX+Hh7S0UH2LsDFfv5pj6JR8szo0jD4xEEU/PTXhAY
acgus+rGCovHxfV7vNrSaE8EhQJ0GEuDJBQIU+h5ahXzyzLv/lcVlFT0hBSHiE2c
jc/4Lspu8Cyu3E/Yo9EcV5HZIxCznvqvbRJK5GxK4dtkzYgUTB9lrChh+usmlHw2
UdmXEkegcLAPlu26SV/vUIV4El3TUFCyyPpOtL4TIbG9NuS1Dhy+8Q92IVphnpji
SBddGPf5ZAiOu35ftuasC3mKZNTniSXyXEn8Qdn6/OBas480BV1FU7YayOfD1m0p
cDJNQwnGWpzWP//gcvt70J8lFF08oXcmrE8kluji4BBtPWmu/+ctvYiuZrJVhKyJ
6oCifn/qucRvXbR/ezlhil3UjVABAXfQ6iTMrqARqXAUfWkzmpuNiE5lvA6Fc8mE
Ml7+xY5WDkcYXZ075L5E2HqBZFNrhzUWmyLvca4vXWUwhhjWo3hcC5ofGP9BQjlr
mvUZu5kwN14OMK0EB/oM4PsPzUXh2abx+bVaKaLuSCR/BGlKXQv4mMhwt96QbEy/
boeNyHfZeSChYhd9Y13b/uGDEdW3Gz0VptLr87/2PsxS2HrMPox5A7i+HahsAvw0
zrfxWSzQevSN8GVQC/1Xb8O3XOrIYLgIAHohMiglkJXUSNLpREDSLrq7CcY1O54I
nPjGr7IqvnWMSVI5/vnOYh29J8LBFPrWtHbdJ/40s9g8lzSuWspHZP3RFf6VU2Bt
XQH/VtkQBkNRnluBvau1m4V26CSDtuMPgowFVqIwG7Dswu0a93ISiDL//629ejsc
97SV1yWvj+gpC1Pi/OcAOChAB3p+hky+8wUCRu6b0IbxUUIogzh4u1tWbKHB6icn
gMk4x9MHgO2sRsWqmImCnWp6xiet9JNxQ/Yzw/ivvTmSGJZqTLO0DsSTGBJqSvxo
6q3hWvtzdkBaS32jTmpr6E1/FZ1FMjZY5237bN+4osBA9cRYlRWijZLs/WS4DzRT
msTz+Chn3k0gxiD4k7bIb7cLZeEMqeYcaNjq1LY5+C/tw1oosvkKsENZV9s88P4T
Eknrc7V8wzyuzWzFAYt9DZmhIkksuw1Cg0YKyCokP+MxD9fJKR9/yfEre58VMKqQ
SWTQyEW6uL2FyCDxZF1yHM7d9IZtpTfBWHEqYRs+HfkBv6ga+tN3A4sA4Upc4LoB
6oOj6ZL0CqGrHo3hWeWGbBZdITTZW1/bHjDukH2j4me2MR3/MVA5JKZg+N0zMwCQ
pyDAMGikBj5Z3ZE7TAumoDzxac7NO/UfsCJp2tfEKMzc7Z2BRholjCwKfvKvc+ZO
MSbKOgSoEJntC7iLF2UDfiMP/upbP++TuYfBOpQi0KVw02s/jtYxvuo0moeyYN07
frua8bt50THFi/QQzYKSBid7r3iCxhrcol9Eng0RRbdXkGuClMOP4PF0oBvlAlVo
rlHXSqrmYtZDErcqyYjN2wasdfDmaZRiC5m39s7t8qTiNBSusk7zaE5I6fJIvysZ
5+KQEJWr8LBnGmjM1uINvUHS3zOiED+LNqdjjSontE3BeR3SXomHGqIY0nR+4GU6
RH/M+Yz4yeGQQzEN2S7ug+SRMHsGEHeCgpRvD/iPwwhQsKMFPGYgQHAgbmggAqhw
Jv1031UX/ebVyqfsU3Jf5gs45vt40+gXInpUe8dLDiaximqfFLO5tk9M0Hf8hS68
LTRa1Qt4DxsMEom/5vNvG8A/4cXlMveyz7E2hjVoSqKEhhEHwK6s37RB8zU34SrS
0K2sB13yDxP84zZTDEjbsjNKZVnAVm07xqG+xEQ+Ef9Va3j8B3cKyERcT2DTdDmZ
0Ni93oemdlmlviSwkn82UZVsoI0/kYfqMRq2WMgfJje3FsfVcn5PhPZa5llliZOH
LRw7pom8fPuV0anNVdTYjxIlksUvmzKaW7F24Upj5z2jdgS/wmI9F9HVJHLB982+
yD+yQZjCnJMEbqtkj2PTtcYGzM8mUSEaSQAA4OYqRVcCohBF6ISbl96RRCwBSIm3
9lih8/j7HBB3HwizZwnzPB7ye9SxF1B0mGy0eKVvW+ZMfJF0422a3HjpzLQKxBlz
uraOgV1Sj0oXcbbVk/CQ4pHi3hbP1WkkE3r3br5xrz9F4M2+DeczNpauPwfJwRMH
VeTNh/iun4ptB0kw7T5RcJCtm2WtnVrzBpz4NEBZzzHeCcO6QyvTT0QF11vWSepI
M7u1UzSNCWbOr1LpJ4galfnKopQnUlnv4Ch2Xt/MkDJxjC/NMW/rS+dA+z4qQbs4
yn2N7kyW5qJJPL+nz4lhUcQvwsz5MoWWUB2HEclthFeQDQe7NLpk0iQG0Iuqn5xw
tJLJ5YXfHwuZ5CakoXTCgQfO6lSsTaCnt9L7OfyBTdxeCfK+UdRHBsQChz+sRRLr
b4QkDZYGANJgl3yVs1w7lj/2feAdMLC3MStlwpdGX6AxSunYzvL5qa9g7xZWlYnh
SP5/pXA2AUW7/I+M5F7O+a3aWjGqSvd6UkcL5j1xMdivcFJ7gOsPEUVuM9ztxbaW
GllDQyw4aUJkCADlwAyrTYHOE+90xEHTicPSsWj3z+/vWwhvabpyo/ORL1cLpbpH
gqZdJpxQrla9Da01XvexnjI8foGzU67FCQExxg+b7R4YxSWYuHPW5a8kR1cwpyTW
ek67LbhkoEFvWojrRyM6KOd2EEwfJXmNxhwOuMhhN9g+Ho7d4OXz6QY1FzpDQErx
y/HXnQeMCoL0Vfqt38tzq6dgUzvRfmFbkf9qtyb0dUT9rCh33utyFIxVOZkzk7md
k+DTyvnhP+47B3YUOsu2QR+cFhRzpKPo7cc0UrvT7rA15vOVlXyt7ssoHMK57Lxb
gV13aRMS4wWnhqX924f1KrOZbey5uWQcaJTNT17pnT58jDz3oohotdtl0JhMX6a3
bX7or9frW+zIr47dwr7TOFGhSs+n/zwPXGH6O/nhTLRZEkE9AS3aB1P/ObklRHmk
DlOQHlMUD9jryeZ68e6rPEId0z+BjH+fAyH4IzZeYvg+n3RPTn1mNVEm7vJ6UwjK
RB9LtTLwmzWZr1niK/sTMFCxxtMKakk5mgiKJPLCBQtA+5P0qBRZMUk838FGa2Fm
1IJCfGdIkLMcGkgsLR9sgIABQ9Go+PR0o2FVCtxmsrAuBLdFvUvMQn8ZBW1oDgz5
npUdO9JYdARMPOGu4OA1LJeA81gm5IGPQovsVDJHfM/fN7g76cCc5yLwPqjNORLw
Ny04BWMp8nbQ6t8/faEEBuhxPrl6xqnh0w5B0acPAgUOJjC6j/fJHOHNiUSB2J+Q
9VZRSsYs5aDPDHo4ShR3NSrBTffDZxoDf/6Uo+X3FN/VlNQNI70WG/SGtXKiPlDv
rBLopEZFadLFPrcEGOUjF1T30PXo2w/sxcoNACN59NNzhHkAL7SjZngv2MjPyTWq
mNrBnHRXT00cYBm2rsUlnxPPjyVl6BrsqERjdVFaMYZn+F4WdEcwuJf0nkAlLBVZ
HVSE/4D8vz5Ly8i7YR6uOPz4EKgwfgvM1sBMbNz6K92rvWP1Df7W5b7h0iE67JGu
cQJwat+lA1+HVAX8glTl7eZiWXZ0iKtUD2KbUXJIlEMNvj5mGMe5Wj7tI6qEPq4V
sMo9OTizQup21oEg3C6LLastB7Hezpk9DBV0mvpc4vpTX5Qu33rDUEyC2t6JksX1
9dFE9ElNb/OHPQKsG0e8knBlVMqyETa1BUy6ahqqNB2Xk0hXLA8YoQieBYRJV/mG
x+2ZJ8sM0UW+gyllqf4o71NCUON4kc5pAHOlpL0cHNzWpz2Hzec6t5X0fPaY56Qe
46JxWRJjgCyh6n06/e/V9ngwlOdLoPmo7NOAltZDu7bD3K+E/99EdclwS/8tSuti
9XGB0zVhRwfWSISbR67vpUOUbGU309acucxwcIvXxpPnO36MgTeVDz61dpRQ0q6n
csyuq6N5omYfsl43hSjnpFS3ley48lOzKY2YVEX14lJXSN376vYCqAt5K3hiH4yI
LykdHHabrzDj0PEEoDckNHiiRut8UeuAW5AfkbGKQzlMBx96azIYYIsCR10dYBNJ
Sdw7Hv0Yw9/RABMigmBzyI+4uMxTAkOw6Gjo9+jvuelg7ycRNYVUz7BonQXUCJR7
CNegYqXVPHkPHm+K1kE5DViNcoPuocXqTynVyfNg51bP3cTQp9pWxksFTyXIe29A
2KAAeVORR0B4eyAurYdcdFPaCuJKVOxKU328NxM6SUOMKshvuVnXeebcd9nZjNCf
qdwEFUADnLizvZxglE6YmxmVFn/1I9KuIxnfH37f/Au4AJz4iFdb6vzbK74WDe1N
0SNwWyDH5P6tCwO4qvDcWOtzn3EGwXzKp4ZzxYNKgixFAhCT4y65RZiC0PBD6gMO
fd5hNdruI6qyF+uQhPDpvKHlhtf3sT76SNtA8KufSKP3I0d10Vi+HUSh6lSMT4pF
pwWM6bTsxtPf/fDKldneDolx1PWc+R8+R85svaccTWfLZ336bX7F3q1rPi89yoF3
l3AAMiUsd17X+FNr8ReWEz7VDHz0Sa8uk/HT/umbOfG5mLhefdQQ3edln6yoJh7V
F9tmE7o9GoV3ureSygFDbS4hDJ+w/6kf9nzbdmol1RUMZZBjUN5uF4KEzQViOX23
TVIiuWgEV03czjuz23bnMh6JsKZWX3gHDUbwSrBocpmymdMvahaKNlnuXohJg9Gi
Z5EyUfierJdbDFixmupxRMVBdeNOeGZ57PNzI3adDzNrP8RlX2Dxg24h5LLYkXeb
FcZ5tHpUQ4CQywUse07h8i/0UKFsW2lzma9LFR+rKh0dgmmI2sSPxoi9Gb1QZ9We
RGC7rA/4CZ0Z1h9Rq/6x0fWXk1cidgOSnsKeIlubot/G4B7cAtoPP3J59N7uieC6
C33YV3wzp43ZSvSxuAD0ALth4yLYXKmK0RtsdcSZe80hlAfmvYiQII0urq9nY7uP
D/WWN7+ceHYpwVsVRCdvGNcsYFZWI7bNVeFebaIkq1oWk4FHyzysxLuaL3v1pUxy
+r+PpreY6jpVjG0itCmaiFysK0b4N9qO2oAoYUnDcelY0gJYMA7WL2+jsffvWaq8
VgSm2Ul4yt1Az6KtUSi/0wUs+vwDEtBtHuw9xJXBkmuFnA0H1vqO6RkGdXf+uFan
XeoHsmvb4TiQ49PB2owEvHZRaioFNifcW9fMAhnl7thWMwia/Kfht4X7wMTCbgOq
Woto3fbVGSiOpup+b1Sf1QkI7ksWPp0TcHpO+mCCwdCVnYgtAmZRKRREjIhNYrn1
ENVBdv84N3RxQFSpfNRyShQmq4ETcufhQYywD5DeOcktghUrWECI/JFimclG6+ZR
Nm0eUhCrXA2tJDwuVUyjsTGPM4oLpsDgSkM9jJh5a2J9fuqfvGkVxYBV11uDVnlo
a3ogQfR6QQQFfyVaEUjGi4VAqgdF6DwWG8yfMYlHSjcpOJ/+Bb26UozV6cQgnxQR
tqDRPN3dLefUY72knNWehAgPu3JMbnrYFoEamBD73ykrpZXdk2o5o/jBtA4+I2ef
+Bd5dT20xuxeub0Tp+G5f3rsKsG7luEPnOatAZnXnFAQqqFj9lzCCrPaZ0tIg/VO
6Fuc2DaVSNeR4hcozIIU6DhbRXSG6nXCo1YVrWBOK/nBfrWy/Cs6si1vA8U9AkcA
ZjCz+8jDFxIu9evJjLs1syiu9uL93APywaVPgnU6zejefrh3hogr/ICh8OO5Z7O3
KEizdXDocOUBuXZynwGPBu89Juv/t3nAkul/M+Ma3iIRecAhARVIakWO4wePTKg/
B0wvWpZJfU5R6q9yW7uc7BE/Q0ZjV2MSip2k+p3vLBwJdNe56BGSJnywMfs/5Yba
AyzP2aMa6JUrFTKsb+Hg7rO4nuXhyrRdlLhyaEXSP0A8oE5Xn31xOmt72RL63xIG
ZsQ1skkp78bKDk9V720mkP4UHMFqoo+75IcSi7yPyS47BYmhFgN0FtTTVziJO6qn
wvcYXE+awner0kyn8oGZO9BTsEnqkHLKAqyjaNjIm23HF6ghWO570pY9CADgKl0H
FtI2QUiyZDESPaEwFzVSwAatvLv8zeK2+ZphcC08N6hpsob8JuR6wkc37xLOOZov
eAfT08KlFFi5pfvYUEfvBhLPx8wfvKWS+nqN0E308vDfys8qchJ7ZkGdnLTGcjqR
WzpeV6M8fKcG2CVoikVmLz2knPPecb9XMlcUB2vlpT59+b72nmx+y3VgxAc972F2
gT/OXO10BeK3QtRoO10/YRMgncv7uYVr57HtPrMJ027J2UTxXewpk3l/rumKoDxd
7UF/jrswupbedlgwv0humg3TjQ41xorUpTNvRgMpOX+LemkaI1bh/8x8B22ybPCt
iRdRHVO7rM9xx044w2KXxQDeWNbLN7wWo5JM2M5WWQy7aRGGy7EFpBSqlqWee1i1
e+5CS4FXVqYCvtZ72GEuPdTNrJlAzF69x1FCyrNCy7Aw18duWezUf1b157ja9zhw
tN+q2AfB+Ws2q/U3UdEHyDjnX5D265FXHMGGvVNunElU3zzTbUBljzIf0bRlP1EL
8xCw1GLmIXGUE6bgpyJUSgyRWD2w5ZaNYUUk8LpVAg35C3Hp/vbZjc24jy0XLXOJ
1+qWKpxW5gIA6zgsmgpRwmxb3P5fPfIaOcsmPiLaGwH7cR7xci1KxLqgJealZard
B093ofx+Zpv6eqVo14O5s4NBI4PfR64mvM3yS+v/YV7WCir+dswPFQvys3DSMQaH
+yjSHZctf7ttdHa3I4Os8KTodx3X/lRoMOOQq6/ORqQpxY8zILbu2RhDNiD2wPFn
Ecl2CQ+A4pl8e/sg+alvnLOS1g7xWUpasgBhz5ri6BowzBbEKt+qHJoS41BCDRff
uND9A2a0dHyghbEMObITtjKTud+Ur0llBUV2UVJBNlCh0/MYAbfpZuLbmOFY148e
TrEs8f1ZJ/3vZMpokyAY3FRJM3hE58x48DsqZ3e6x1F6gfYQjXQ5vMSdTltimnHp
M3OyUYF7a3J0aFxC89AghDVZKdQzw4Y+V4RMe6hKqzjCtC243BrCRfQF2n7BKt1H
CVIPqa2zwW/KugQo4r4OEX8emfMyK5cYfYuhOgyJ1YhzTRr3jVzjiJr78s1DaPTr
YFKW8f2R/YFm+zfxZU6QVVSD07RKTgbKdQWswYryWpdpaoLJjz5l9SmzjGOArxNJ
Mj++bAZSW+GtZ5k4dtJsEMhoj+vZiIZWiOteX84Yh2wyMbq8xeoRfyBZDqocmdIS
QZ4U4ngr3BY31gsurgpkq06XS/BvfGGrIiq+NmejLxgfwQc4ME97ACqRqiBAO1eq
JA5OujQ1nZv3RRbBLq8Q8PP+hajQSaFudbtTpiUgPM5aDwaXMIeZ6snnai9yre1u
7UGHBUYu05KBsCoSwO1BXxwqHpEHEviShBeL8ZglS7CZYRDKXdTRJDzk189XMrpm
vAbOib+jqR54GRn7Fb7MudSGsyKdHRiH28tPk2DOeUkMOcQTMu2FmzUXkoNcp9hk
BxEoeKpcF/eDAeJ1a6taD6dBZ8lbABkHZHlNMD+qXTSCldVHTB3ZaSHdDyBgNxwS
rHUl93e6TxSLBzwM3iECdmXb8/3EdeQP41LvqalQ2gnsPzDFJ0X7aR/fMqA+Bxic
TTg3FRlvm3UNXXW6FTvwvz+dWwocI3soBx1rRvh7RR4Zwv/5vMLxRh+5sBs1RHlp
0gI1b2UegjVFiemJiSLicCe4ayeb4x6IeDxalXeVZhVyZp/dNv6k4fAIzC7v5tFW
vcsterloU/YW5pdhq+B0KQ/bxnHxLyekhoqNzy9p1N91ob9D4xKECJPE2SrG0SC3
6FPcKY/XbFXG+7ThZ2dkdvuSOOS8rNdzPwaMgxHe+p8ctRA4xsg7Fnn8TkSZ0hF3
hUIKNo6ggkazOgQze7wXPc7a4ZUFjZ5Sc6lBrsdLos7As58jj7LvQ5qixloP45eF
Ii7BJ4wDUEhQrQ3FnbEvq8cGTqCuYPr09c8OPOah60U8eE9m8nj4koMdnG6a0ObA
FJDXvBFLvv6Bylefl6KJtNQr3vteVu07NxQxz4dHa5hwxT0+Ly+n1ztonrKVAn2f
vShdp75pde7h30iOWwtqJ4rCtRwyZK7CXJ/ZrcpTDeohN6Wo3mjvEArXKvKznHpi
x1EJ/BuyEd11LGnbAs2oJAYrHlMzZc/on8+zr4C9lDJc1XwokKRLDWucQAS8JrNd
fMix87I0Rn3fkRStYHtMJ3B5vu6In1GhwVZxXmos2hKQTfWKs8naZMQvu9oe1pGR
oNN2n+M13qkbpLSl5VmrQDBFZzHTklEPJqijE3FXyPDY393sp7b8qJJxhrI6l1AT
36IRIE6zDrAPYJPswi8/BiqRMtRBCpVT5Olk+UfVp4HOv7lQ5J7LwFhaB1ZRQ7Kg
N2Eg6huoxvbWA7U3Z5Nra3UcZKljI5STE6oqebOVwnPQWr3r4pslHNT4CIfp11IP
I2m9vmrhGj/9klnqnDv9YdTtLOimBjSqF+YX3++EC7bNO8QRnsrPpYfA0A6B13Dt
E8IH4/r0THYHydb45MBvb6ynogH8haRIsQdIHcTOzOIX06k6o49aAFhl2kdez5oT
a2VlVKfP840NJbPBHzXA+EUf8WtEN+ug6vUr9LQ4K9ItB1N5AIgIt5Sl7ibH5SYL
udAC7J27wQRGxviDqM9WM9O6sVQVCln8/RN9upiffbqpAsXzeqsFy3x3xnHdgxSn
x98SGwIxoZVQLIRZVe3ERFWPTZBGJSLW8mR0KILjYyK2RGzSCwxBfut5X6wKnxh1
euIj6nxjegqPBZHJ1+/Z9t8l69UeGBnh4FgFe0Km9Pq1/pkUdTcTjjbX0TTQlAWo
TWt4xEZng1zgnzPZ4Zg+ZaXoQ1R1FB7ho+/27MFpIXp3nbBQ3T3xGm2GeIQusypP
aZ91Fvcqn4U80JT5VYwqV7sSzs2B+8zdBQAxnKiDl/+c5jc6FtlgaYz6pxRUKTvj
Wm8LJlT4iVIWYYX19XOK4CYYkHX8IrqlJKx/aYHieXxFEdT6jTUktVzS4wOyovLr
p68Snz0D0v+eMYImB9D2WYB+CxSNxuUgvrIqaTnVhJc/AqdnXWKm4LHdhV6ky8Op
FrVkWDuVLAgJT54PSqfIRpJcC/FwT+WdzdlV89st1p33cMO4IjUhOZ58UAcdrftr
5kmwk27cMc1/hyypj0HVj25K45s9vtA3nPUtVebS829MFL//ru+EsAjokeJyA+tt
coQNd9PpXnAntfa+BZQEZ9ohpyKliliTXdDwAxIdseMMsqrLpr+v0Nm5xwmPEHT0
O54G40tQ0Pb64LRFl1esxoKn7LreVsvuxv5iuMQAnHLELJLctus8/VbCbTO1nCXF
6Au7BJ4cUscgdJqPYdZddljm60PDFksbMLXwXbVN7HhtSud0k7CYlG+gKKTnBreY
g0lPFfIkEhCkOeH1+/q2jocVlirIT00tLTocI1ER1uN3IfRDnqj/iK/YhinZJUSh
lMHMaEE2fM9zbr+njhCnMlUcC52gU1xmBsXBpl2BsDWp9OkiOogjlySypKL/9xDJ
XAT25KteBJeiG7HP+g47WxjvisB7RzHnGAfAzObYB7YOx4053VO2Dfp5iPJYGW4F
u3kdSoziNvepsJekGHyyhuCdiuUMLTliV9V/l3tG/INFGt7SvFCVRQAb7VSYtoDy
tsciFOXqLqA3HxaMh1c5rGpi8kh4nfcccWALTsvR1Y3KrT65K/4f3nvClnCSeOBj
G9Zl5/izjuZ3hLc5wLSl4HaxynZ0QqIUDDBFwuhSJsTS7VofPEHDqp0HhlNo/f1d
FM0fTRx84wkcozv/7awoFGjS94D4eKl8oUA4lLvzGFhgGMw5TQEXqBF01rkAfWMb
9xRmD8jkoGiGFXP2YZ3ZR91AT1FmE8++n1wrraldJPf5u7LUHe7qsnM5fFN+4yRk
APJRrYbMUjBa6P1rOhstRoozQ5RGYjI731SjzCgO90wEs3V3Z0R7XTBGOfY4lvYm
f67TW03hkvmOZSdoQRuC5csqk4jppVibkis+jlfN0bKeY/fqiYsA+omV4ojKg6Kn
EL0/PupKBpHsT7wmYQjiQlWZ/QaUHIJfplScaDFvUixwTRrlQjKNikTKhZoQaMjX
rdPeQQ1UOWbVp3PPH9q5iFroerdc/RwOAEfHHa0PtuhHlPT1XguPJ8UagRZeY3Wp
D0VwvolreP8BXnLrEE1DQqIaZUCk84i5MCSLyXpdZXoRdfH5Wp+6RFgapAYuuINy
KRlspm1mqHHu0qFx0s2MWQ6e6jL6qfWIkSa7C52Sr+QzrruLh5a/9idQrQxzLIC6
d/yiKg/lMyadJFgMbHX3JM5qns/JCpiqJzkIrFgDDS/uHXyp2axYHOtupCHcs3Cj
+OYVqmppOjMgpte69qm2uCFzwH+U8YRfMKrjXCFxuhzSLCEoOqSl/TlhkuyH1udP
3qeOfEa7fsfyU6FdzRZAg+aGKT0H4MumymKqkeu+PD5KjuhnL/KRZvHshU7CYQS9
/Zu0ncAj2WtRiqQDgopKmcFmkDAquaneR7mi7XEzm3RbFPSzPDLRJXtxOdsEpmoW
n7kG7o6rhmr0X34iAezKdCisEwn0X4NTBYc/DrzVyDopDEGJgPq5Tz3nekJCZD3S
FMEA5lBgs8J9OnWL4SCnmRHUHo0gMs0QdBXy0LNd9XWxmYi4NVbp/6b7Lb16NXAV
M2T4G0lhRXOy4VQTfUQ4RHsCgtIl3tqffJ4ew8kY00k217ZY4Li0CP0SVnGHeo/W
udb3p2uAMRma/leUw0zy55pjQ6Ls6G4qeAkUpmOxGDFr3ZSrUVjNivzI0x5xyeam
R1q3T7XG1auvslmokz8PCw/lbz3NcCmLBIyFO9tlHS7KA0vl3zeq93wuzFt6s6cJ
YAj395dwN8lhgYbt0FKXUV5CtfGbTJK1GHuhbihLJDCZ53QtQ0MZdemQiinYbzpa
Q8Tt1TXAaX0T2JuYWt1dY3Z4nZQzNtFMia7S8R3T+nUXmFLzDzUmZ/h5KB63sTns
9IuDcYO8GPnO+f02wcadjddyhzJsHfert4D+NrbQfOpr9TPURfygon1Z/M0m5NEj
cLEN/gF/KvVW4j+lrPqBq1OeP5Of6YEuly4+I3dwplOK+80HCgge7SUu9/p5y8Z4
2JFAUeKAnGrZTpB0D8CfrxLKLvlsAowh3OozR+zveCJOnK+13/fLcOt8y3VOE5BE
bsunq1E49BGDVrVSBiLcPCKVvAuiunpeH0hHBnPD3X3DzGE5NYVTa47V7+fzzp3K
FoMZZTLe7/u6pSzqYg+SYX/Yxqa62Uw3mukVGMjiYjqf3S1muMsN8ZRUgsDEFR7Y
q0jfp6XoxhzcFsGCbT2P7wy0OPRuf9cdYeMo4xpzuKEcvWpyhWShNhNwZkklr+xh
u64ZWBu/lJWg17HKNoRS+piPtOuyxn+aLDmmaJD+kDFHJxvmSP3OvVL9DZXTPgbo
UkLxzXHIk/XUhgDvFfciCNbUPgMiSANrj1iaQq5ZKtGNb/Wums0BbqTImDRRalvb
Z5w/xWqZAAr3vnqEbdWkI8kmfSDJzbNGB6pAorz6wGeGfEgCqwdLBMtvOBAyanDg
NlhmUAiBa0P5SjWwxL9pyMm9Qt2npMBQoUhr001H11vNY04KuCNYx63wr1WaUgTq
jYKjvVAilBTyXAL0OhgfVyFcYR9j13qNRAAnPIdIBhV0S0MTvzPj+dFi9vo4W2AO
jle6/l/nqZKyVDmKwvc7BZ0QX3JET0LEDYan3N9Q+c2W4l/6UBrkrPWrsu6CcYTW
CNVsL56RMnaUQUgo0tbroVd4vQLgIDZxIB46VlxrN2j2CvkDKWmV27IY9hvzaBOL
efDarA1avvNDElDHRoi0qiJOAXeExHDSpd9vqpFzhOBjbKL8rdpKZnxzOXjqyzCe
VXl1jOc8dktM3hkdigd+bSYXsvrrwSXr6dQmVVfMNxXV2G7ks90dI4+Cf1VhtlPP
HYc88cNvPyIG+Uc1SoIJ4woSxY8qzggDuGc+s27s72PgugRPVawfoI7UZjAsd0hm
pyKHbGR1cqBDpfhsLem7+iehn0zKronj8KOiHNIzIv4/l7r86at+bxIuou0RM5xN
3peJkmNhEiT1eFVF7AoEIRFXha9vNAEpKMDLOb1hIOK3wWZPVBv4om4TyKq84jgp
QImtzT2CRuegEgX5vpbmebfq8mCp/5pDUoUN6iHYs/Zk7iojJ6lrl3KZW54nS/3t
+Kn4pNRmc1gt5hAZnQWlO3Iu6ggl5G4FTOg5GXqt6Cz8L1yYFUsKIRqXbc7Qn0+1
mxescrWQekeWbubozF6707GweFFblstkpbziu7iC9s916HOqcf1pJmLEJke1pYsh
cZpJO/JefsDeHNGPSXDpyQWYOJsl5er1ri1m1nDn6e6o4X6gc+9TaITa/g7MRnTo
478URxNLg1d9GRgt/E77xz/zutFXg7m9oepNfxGvMzAxrPJLjZhrZrCKvOVNLu7Q
ekaKM1VXwg4+zL1UDxg3xDGa8l1jlJMLrSYBAHy0bgbj85kUkpxIg+Xu+TmUxk6m
hMx5l44DjNvFEYK3hbCGYongNvcihLKdiETYu0YhVJQD9D4oi3fUidwC26+unBrN
d3C8mPbEU30ONC2aaeBeb60OZTRg/hpH7tQuOurhISQMnetlqNx1uX4sx6gWBiZ8
f9095nlP7/Mbx62sHDJsGRnwZIRPyDGqGo4+qNRntzo9vnIl1kdLBLSQV2cExvFG
rZxgwVALxRKaDmWS17efWXP3clPY71HVMBoRaW6e+kNlf09vWbWpBGIblJpu57TT
cn8eaB8cUVGuCF7j9HjcRaHaE8Mn0AaNzZbbNMZ+T+7peQyEioDv+7HVu/oGoqoK
a9gdI+gNP8gMJr+Wy+0LZ0wXV8YdGVMrKMGC0hd+6kK4DMY6gLKM7yYUbu313PrR
mpAp+CPw0aYMNpfDt3y1vYDhBHvJ+SbbJSESnX4sxKLy0OmUKm8i72Ryf3U0BtDx
b+93eH3GoTI7KzlRi4e2Kmw8COfIIAyqA/0FUuxLXudZBpVnClPVQtSpH8aSFAZB
YrmY+uHSEaacUuv/C+JUF84ozX56C3jrwHzQLiQ+E262tAFpvXB3QzjtMSKiJoiq
w0cS8jFXTzAs3vcepkae2RCgBaLXMJ8QhDY+TICdROlfPhOsyc3Zw1SIFxduC7h5
X+TIVibGP9zHZK3vMfIPpwPvjP3GOr1ZEKXuipI84PZJ6TSKV5u1oAdBzkHcjayo
g04tVS/SBG8Z90xij071qpjRnnc8GrPGUfJpEBmdAlmSzmxvYcmV09oWnzzQgFYE
dTaHdcEuF3uLVSZ2nEA5+Qut0C48WGik6bMk4jpSu7mJVHT3UHETxb2vhhfeIK0a
p764Xa8edTybvZj+QrbcRBJzzlpRnit6H+oe9IKe9M8WjffXk/1OZlf0jyvG5f0R
M60VhOgXSwwckOP4Znpc1o59FOEQIjx3xlvpsTYZWpHJ/fWlImW5Fm0DhMAjML3a
P33w3Iel3R1rXJ+Iybcgdgu2ekvoxxq+iYpULIKgNhuUBrPlgYawbP6aVnWmyiNe
izxByCcfvmniJE5GAlhuq7adFFF1DPCoPGlnZX4PWj5lmfPLMYQRjb5XgoURoBJP
d1VvPEBRghA0ExyrCgvTFqtsTE7diIgKYZZ+mZchJ7xXyKhG6jxZgSGf73jWedG3
7NbkhfSRFp6rjzdSuwITOXdGGoHQISwp+PPBotDt4QIxaZ6Y0h/nwcdlMbyR5dMR
P9bVnsFnBvB9FYlSDOHha7cQTdpTCJsuXwwStGBEpOsyZzua2UXWxJZu+QgVTIP8
PNNyAnf6wnHMQ2Tp87K7SAhD2PIeBf6A+HetC4nrlMZYtxXaHo/fxym0GRzd9Ejy
L+qXq9oTGj0oSC7BoMBr5uDOIqsGfJGMXo1MJY+hxnSuKXc7N1Ut5bukLaWiRXCi
RuhUJwKlEiIzyMNGlE45t2+01+IqiViS4/BUmWL2Oble4WkHDERQE7NjkJ7VBGzs
PLGpuDhHV2171ha8PAykwMw8LT6eCc9rhSVTMrSn75wzQgixqxMuchlfBfqr12Tb
QccJXLbMCLRV3F7RhL6JK1bEnlstoVUak1LqEoColEtPDNDFKNGXcvBWh3usoMfj
VqW9eKcyUTuOObAg8CmTzUNCEyKHe3Tyl8Ot8aqNgsswKT3oBXDMUt2A4y7ZJ4v5
3AtfbkWI/FJJl1rDhuqh1ixnQ9y31Yp8CTxdoPtckf2DgSPxwTSFEEldZOu92bYB
DOlTl5wvr01eIFS0b2a9u7y3TuEFXxs6RUfcjURVyGMYRezmtHUATn21rtynCZ0Q
YYlZrD+uUlXNfVKdc5Xhuvdsmgq8CsCo4twsjgbmtcxpUSr24OyLnfY+EPKi9Ck1
gFQlEXOaccc7KOD3aT56N4bEpvAE8GIRVq5NHnPlv2RMBMitpB8x0rfYAq1SRpVN
ckQDPNlbrAtiZRj/qmU03QN0HghMZqgwoKCbHhCWUXGR5qU/aRxgu5xtvLQnkWLe
7QAflrD8BwpNiMvSGEwtyPoUGFdzZwL3DIvnlPyvwxztXais7AqlGrcXp8Igruin
/0KAQ6ptif1uAfzzAMQEDfIRDNPageZypVmyTLE4ycqqEFx6b3TtvF3L5ZjtEZFF
qNPhhl31jxuuk8/t3w42rPD7PFiWikonYoCSasGc0CckicAhwzRL/N+V7Sqx1qMz
qjgKMvzuEo9mvIIiPySWW23cSCXs86aPRN3420Yjqcf4+wbZEWEY33U+0UTfqT7s
m9b8QzPddtwuIwI5QYLgnB5CJc2ntgRTNsPEE5cwkCRKtfmMqB7x+ake/aCntecS
+c+nP7X5dnweBzpz4ayhkg/Xj3hdMNcTjBRWHRzvUk1yxhaKieB5L8/XwwWJw8sD
TyAbDD1xL5Fv8vW5NqdqqB8GhgeEQ9kCX9ErYnL/UdWzpjzA6Uk1aq4kQITzPjrU
2G9XejhUPnChKWWujk2H0P3miaCJXavFen9vadonzqBKtsHuc4PJyLHGTtN48lBm
rZ3WiUhJgXSMZXutzTbf2WRJlaSTbQZf3Q/Jqp08QVrYE/5oGC6AGC7fPSqqdwn7
O/Y0Vj7ueVdzYmGCHKLp6FHe3TuSYHwowTBAUgTOcCBnqsoRlubHCaMhLh9w+vPd
gl/bSSod9uQMaHQqnp4KmUWWvDw0NpEw7AWD2Rn5dfL30tQNeg2KjAzUSonwPfm5
/m2AGzg13UNqFg7CfGbRi9tAvxVxTzlnnhqrCobJX63fCxBVcsKNjq2kWI0xf036
8iCZAGlBqKW9HrrT2uKzKcoLnMI5lrnTtx5yuEEjosgOTq1Fq7RQunFJx32ZNjWv
RZQDPe6BmF5/z+6lX7FPQ9qfZCAe+1YmeX6nBKIJ8tBDFtvblI+bvaPVKvvkBc9a
z4qK3ap79qH4tnvrsEa08XwrW2oT+rRKt446+oppejB8wgSezGdEX01vokMPGqYx
MnZis/lFeTcMJ6Jx3Q33pfK4DPKFV1AOt8Jawk8rLtc5TAUk5nIvUk/UWFWw8aTp
FPsQMlH8rruX7oFEEkMeZ6HIGQZfLhIlknpSH3UoodXfmx/Yndj8yvHSE90GPfrt
FFVt9W/9rt+fw2ibuxpwQrb5i0p0K6LNrXzGqrAsrSifCacrSN52mvazj+hPQlC2
dLFZqldGY5JERvUllMOvc/4CgvM77Tl+88B/hdcjksPIunD22UceS1duGawJ+iS2
BCqc23KA/jCrVqjG6eJO2ZbAOQjCcHnhag+J6uJ5zcjjUCV1hDwvj3YEipTz02dr
h5E8Y2m6JOOprVhak4Fsj4b608hF3/HwV4E/IiT3loWoopbdXLWZzuhYNkrurLhr
ov51sxlpDl/NzYx2HNtcrzGr6Nm9AiFvQOxA+YhKN/dfHRRnRwAXJj6E2sOR+iZe
ijWEZ+eeQgU+Lc2t+qITHtcKGU1hEtpFkw2gJfIiYw4XKQl7k/oErdYI9QCuVY13
95nGx1Qe1G/ZiwpV59X95zrKJoYi59ElqOMWii1Fl5yzLzNw2r7HN+qgmjISOzzS
8aRVDlC0zDl4CDPcp41JA2bW8n0i30YXVZJKG8pxcbsVjoYq4rMwUzsj5HLp8e+Q
p83XQpidu1qtvJwqJYRxFVaa3n86WFES7iKhSVOEknARce6BlP4T2ODEOl6FDEHE
Z4hSvM/63uzqDkvsyTbkkerxLPDpiSrci1jeSnIfto1EO3hBjXTi+2LNAfa7eN2E
Z3FOuizhXEC5ObeNw8KXuuPLvkjpNl4eU/I/D273P5BUCiwjW9jxp+gYyxd6V3pe
UmjhkviToVFHpmnRKEQ/jJv6YYNQHAt6YeNVRrZm9QBFvjMO70bxtwMxBwgjsKIG
Lj5lH2H70fwAOTCERuijwXw3eoevsF95m+hm9uN1v3FEbuqc6nEFl9DPskHfg5PV
NzP6brzZJzzptIX4O/GapFO6Uz1f0deOb6EWVAFbNejcTilOju+sJOndCRkt/v1m
BkMOiMRBmwcWyIESO/0oYTgFa5wO7K05iG5r7TlHzMGoRv44eO4Ez3rZSR+7u84Q
FVV9T9AkB5bfqJp/QVzjrHNmPjppcUF2LNgL42qmf/LGDyrSOf/7YKnMT7ROQI4B
5+Ounlepfx20hkNTXdDYWQfb221+g5SPYMJLcfgwwtW6kyLbRemGPElp28WVpHCH
2fYB4dE4w1E1Hvow5BSIfvYv2jX/qs9s7i4JtC6eje9NBO6mx5HysD/4YpchcOsm
vLaE15ORbjoNHKcenw+j+tVgVE1ebbPbg7lA6JmCNdcddRa1JhAXFswq2BUKy0wv
Ag1Y0wMaXTajYJlEhht0gUCEB0p+0mGIufiM53T3rnOW0ap9BWJyVus5cIZejaE1
wht/NpOJfUnFrJWn0NU2RwPBv/T/332IpU1YVlsktzAyAftZmIwgVmFpHGnntRzc
1qGbbLET5sdpnHOo5HCHBmd0o9Z8NhykuHH9uT2+340BsWAP5BrWRcqkIgRYBS8r
tn7TReon9RwH4jUt1uEqLhsJmLL5q9GcuaP1SiDEu/EyjdPimzxfeKX+Q3uY3RV2
18GFo1zUwt+GjFZafq6mgjN24iP5hwo8t9RPTOYCFxJTXE4T/mH21atBw9Rdqvbo
I2SLW68nRr861Rxg47oK8qWeQkIh5IZpRsTztsVjH6WPamqW6sS3MKy/AUO2bc5B
nwD9d1Mj3UtzUKifZVCNHhQWPZ4ZsalKYjbJ0dDxF4pom1ZGT5LOuppt7iQKySPA
EEL1GWINC3B4xwVUaEsmGniL+J+paCowLsV4of8bOpP6cGGgpRgUqXaaO1H3Vhr7
H+YzXGbjOFwZDBx6vsFFugXucyVjvCIGa2G3CvE+lXDdAnXk+kgoiWNB0fPiW1ft
sSZlRAyK/Men7QqzVb4f7D0WBqNnYELrb1bHQQl5oB9w0DaYPoMOKgfvrNuJg8jt
05VkggkquiF4OXbqjIuRzVirrpXRSqZaplScZfzWiYjKjZt/+UgG2ocUvKuhV3i6
egxgxAHjBvpi2BHszSe4PIb4n3tLJUbiEzz0mtBSrdTBGBJCNxrwIG1noKmHm7MR
/O7EnWJE/FWKKd8TzAlLRTnQU4ZGxc+HLaAMMK0VsSR3sQEh33V1J3iszARi2Zdo
+5WwVGlydxBQqZqUznxIw09EzAfBsjpI+prKukE2gJ51ZJ3RK+3SVLG1A8Qxvj3R
z1JFAoUC/TcEIePNLH7frVRbO2qGwmLNbPJpdAUX7h76TNrCiA14cCkAxwhqkK52
bkdA92Bu3LowIFCq6Cpb+YnIGImHbleFozxKd4yISnDf585qzRKlOkl3dAIRviw1
6k3qpPlrCpqS4eLwMdZpj47jw7FV+hSQlD2xP2eeOUr9g2bLqEb+Ip3hb5OB7/AT
YJcPNsqpES/dfdLxGBrlMfR7csYnBB8HGT/QJezReu7b4OSti2uwihqHa61F4ReK
gYKVC7FgLy9xZOPdizgGkhIl/EAKKxFS6gotMbFlqdpKby3LIZUPuQXMRqvMSwTC
Klkh+UmzKIWSAg6kUp49Lk49bk5Tfm3pj48DDlV0kUfxwud7HDYRPzBtnOmSrP2a
sHHbY8MCXyRuPECdqahQYSPv875CzXaYQS7Dwf7uuqe8JeqhXaZCyb4j9e7qTFl8
qczFADRgKhKjV5Gt3thvR5nNw+CNpwaJBNU8JXMbiQAHDBUhG52AC3W0kQ71CLsY
zFrl/cOVZ5ri4zjWuqXk/kx3JB97gH3lbXUWVrLvn5l1AjFHYmtk/xZoORvFayTL
Pr6vmyWAssAzI9WsL1eSyazovP156eblBwWuoxUvBLgu6EY4VPNtvCGRmk5tKe+0
c3P0ctsk1UwS/enjRBsOFJl3i6PiMoYhygR4zdlZZWFJX6sKjCCrAISpTzbEtIHr
VLekNYo4BP7+Wj7WBPlg+Wg84tcWd+/vP0PrGMG3hhhByfkRzgp+oYD+XWE7wilq
0sh6Fq+2PI+HSm6LlFDzZ/GYpXWm9IzgcqBDiJCqyBN0LzDpEBn4RwIHFb1mp+CL
x6k29spi1/HwSI42jXYeU0MwLBZosMvVDhUmUNDzTedLEAP734npjSTXkqKWkyYo
LD6zHMfpm94t03jVEc8f8Vd2Bh1qcGTWm8LoxI97bNEDd4e6M6Eq1MshQQtUqHFu
4whgGOrqBKg9tMi+Ap8Q6PhJYHxTiyEW7OICOpVwn0LYHCD9evabs0kkS3sE/b0H
3vhdJYwTGJ+88iGhKPGLeFwK/KQ3lJ326Y37lCnla+5LxMQEiyBeBcphx1ikq5Du
Po3WdJhl5mfVtOHBO/nWIiAhEEIehdILbR7jAJScO2/+i7+O9ZYLOYLJGW5Mmh7w
Ja0PDbc7zgBEcCyW62Epiv3XkGC0/VjBl9VvFi9Hf70V5hI2I0SAqEeoa+NH3DRg
kxX8XhwLeZAZ9z6kYH4OE8dqnU9F+EyWOMPmCQ76urRvzNXSeMLSDffmZfnRX1CD
F4xhI4FIJR6sn+g5EJFCFbz0NkshkVG9cBQ61FDsVyXYzvf2NPUmQQaSioNs/oxI
LLXsuZ4eZ/nK+noN1HaJIZliyBNdsYOaGPvPch/v64LNVu+Axs2ZZLN5nQGi8/eb
4flhoHtjCepzpWCHqIRXqCDTWwG3K9zXCg55qCjzzrqYiQRUBfA9CyRtJp0ATCc+
7Of+Ccaj81VzhdVISEbwtckhrAGzdfemAEUxVHhDEPWod7Oameu34ROcgaU/PI8n
JswmtvpH+2j4Cv9C+LAvYR6bWFAaboq1ep8L+f7wxFdlP6WUN6/+RJWFu+//RkI6
hFna4g8K/Tw0KC/WWPIG0ltA90SmXl3T/cs8zfg5JYLHG7xmOUM6yr5PHYUqdBAM
EkWmqAlxZA+Wce6j1VK+gjxoeVpQpkL/yqLRKIsKHBLlbwpuL7zQkEGeRQjD9PKh
3RtH3C1ZssNyzRQCMAbu8lkBI0olKW+CVdQssAiDVATZdvGRN+PMcYKm8JfNm/Pm
M4Yr5pe4Xkrh400LSu5hMo4q44WSCnjmJ29EQwsKc708lRU5g5UQyqblAxzQhqK9
MQy2tvr1hEvR+pPZk8cbbyxr//kk83NfRxwqFhDqAVkRBqrSl9gh8IYbRIK6uAx6
mmarhoSufvkOYdZUFjCsmI0zkxFdaJWa/hlgiROHPwuXZz31H2DxBZW35I1dLpJj
nxN/gA0f8twovJRFBvJadEpdJDJD+pTAmGUy/mwh28viJLbrshubeNK2+KQej1QY
sM1+hHH6LWZKeJNRwpH4zqxIeLVSUdpUkVfUF/p3nnHHyH1wxDTLyOtrwJMR44+9
KYNIJDt+TZbTE8FyApR+yVcTbkNiS7JfbCsN6ujrYjrJtxrpOC4QrHIP6teRUPep
bzsJt8FhYXMtD4zM9akjNiIr22vdyXrmYNDTB4t+07l0YpKm4mjgfrxw0PmR015A
2hOoqOG0Bop0IrZfA4wNQHFiDFxoaBOCl6TFh8v88djvWvTCmsE6jWZB5jYLN8LJ
jMi6NM1AtXIMGb+aQlXfiZp3eDMJRJemTwzYcMJSIQ3MCtr2cK5LRnJ+y2g6FOPZ
xXBUmLywljh9kjDpgVwNVwY+4THGNZ8sQioA2mZCzj1H/nACPXbuerpRo0ZhEXPu
nLOQKwz1h1jzW1o6Xg3oDrasbLfFfAnemqz6cjcj7utdlJyASuQExHT28a50tagB
3VsnvZ0FBCiLT7hSgMlbNB8rGVhC+a2yp9EtD09KKbDJFHhSWFdyYyYKMAI5wEfB
Nxsgbd2BV90z81Xxb/gjjQC/V2kzjc8jqBG1da8kUI3LW2hi2K8jVeGgceZB86Sy
jy2KxY+9KKb2UB4hgiLJEceXs0kvB+Ytvr/iUKVMsFetpHlONiDtpK4CRhxK/5a9
m4P5ghUoEWNvP2/pqYhF6tMUl0x+M0eHoID/PIfinbAevMYnppxEFl4ssULoYSyd
R/ifahqU1FNOqY1wjuR2Hc34j/anD7o0/5lAkSx0TVolijimy7azOf55MZhDlbr4
H5FmHufvW1C7wqnJmvUtdAY4MzCgDS3an755cQ6fPNQQLZVsO1Ot3hkg60sVu+/A
E+mOGpqWhwB1RSryssVTK+zr0/2q99Nn/vVnt9umlA4att5a+HaJdRmBlkSj1Id0
MA9iHqFGKc+I+Cvc4wEX0Qbi68DI5ojUdEKT/39O6dziIh78vGv/zKcG+wkmJI67
6XCszk+kaTyO71BINc2A2eSCDrpmK3bk/0v4yFsKqZTZSq5y9nZhDkAnQUYQoWFb
wWR/YilrbBsSUHHCwwmsFrLiL57rKIYkmV4QVsMmvehEoLk0YzXeCEzBHJfgIpwb
xfQI7HW7sjcxtcDW/DeHv9s9B72GJDnsa7/NUBmR5qIXgjhU9KWNTnY5vIs1J2Bj
v7L/PDVTWgM8sEf/cOUZPE+xpG0gkbhuxnuEvHY+AEkmE/yoce8zxZgaCfZZML4k
9g4jbLVeSrft4Sl7PZUM4qDBfDYO3hYKO099yT1ig5MysqSWM+JyRV6uYz3YEws4
2oviZfcUMgXAtnO4CYpTM9AnyHBhnsnNa/PRc6zfsEQnIoUYTbCefYJj+f9PKyGc
77PjeCfU7wrNdoRXcqigVr7tKvBq3X/LWP6I17e8AcT1WKET30zercMivYhBnj0z
rJveQesGH/IxsOj4ETNXPHdYNMfme9qdB+9oAr5MyDXRCF3cgS4Vu6DLZ8vh/dYS
YrDOYadLBj3KEsdmmtBKh4Fw4coqDkg97jj3T2lB/OsrJJeILA2lUCykI4g4keKP
FvE/Fa/YWAMHWXVYPmFQQaGeRKwAa+TBgQVKSTnj5pxj1W0JBIvt9cAu5Lrq5f+v
Gkdt8ZGg0/fZxWdydYRtUvPrbShtMP3onNR2unXzHgvGpec7hsqBgOqQQeebxaNA
6gvvtJLwt4qGmWeGv1Ycffc1XXfG/TCBALUM5D1sVf6qgDLa6QYlMUXLVHVn3KZx
PFVA0zJIu/VOorav6dXR01tFcNGoVJ58nEtRsa+owYuMX/CuOXt11wG/4HHCRSjJ
ynmQlF0GUjQxd2RcA4deUpH1n9uJf8kN+CSGNn97wQRTfUtn1/461kUg+M2NXhza
97mC02YSb9XsR/NJOicmcCgBU+33buHmf/1H+HdanAdCb8OyMKKTsYivBsmEq/gI
uMBZEXAN+4poFIEvhUsW3NM5zCBDVJmuQUuU1M89FWS2P9HwGkjvx0EUWM216IxE
C1wueo5FTntkvZf9cTMeGqjAzfUBB3jtg+r0RGmM38WmOthfseFi1ov7dVHSom2f
pUVvpwzkwU59Pegt66E83GDb76jfssghe1TW9VRX+eLOoPn6muH1vCHHCvGOd6Ig
7fcj1MYQuLmCQovTIgYsQz9+poKTa/BFnHm0NyVYNE6rSYnfLKEdj4AhkB26By0m
ucMhpOCsbLSxnGujRgUlOyWoeRJTAiu8XHN03lrbfYhbIm+riIauSxyABPyO7Me0
Bti/tPN+FCAaYcE7RCs50m4LFWX8Q+XAwwq2utmubn7rnJSvlkIB2nd8YUPai32p
P9SOLbm/5SrbkvihNauzRwWusOvrkuF2FReac3L4Ha3YUeSyoKArAotLWnR4iIYE
EGR2Bw6B1pcVUowY9vBCvuVV7w8tclpou/N7oKg3uN8LajHhpMoEPWGUE5pOg8Zi
wkCEzmso5a7rfWTWCNg633Jx9fG77D32U0CnFCOwsMswyvkMRxOfhkN9RIn9+Tfr
7mkPueW2UwI9xt1cjkVIpwFYC17RZQwRRVuw+SrLUpVAkhaYIlhhCjbrzlecWmDt
Ys8oMzK2751Zg7OVLa2Sf9HMKhT6FvwIyaIvBsIb2AKy6RLJnX/X2/HSA7DXtECT
9uDync8u+MBuzmI1xavF4LWo9KgYfeCS7RGurz4dxVEb29mqZ1XgWk2MMqvvLacg
GfR++1ZJXgVAQRTwxSNiOqrgZy4CvbNcJB+j9F7pUdqZ+VIPlLrJcbrWTkPC9rmJ
NOjBu8H9LsBf3IUZDOai8efnoRupxA//rlY2dqKNEox1lxdOwGX8IcEHgTfxC4qn
8e9ycbtZKOcg2BJBjEsX5Z8iuDPPfgSH9j3nf42Y+JBh3O9yMR3QXqbf9tFoxh8y
Nj7GBt5ZFt8XsQrz1XZR2s0DWx9ZyExvnvnf2kacjnEB6ZCYP+Zv4vvuSwurRODA
j05fEHvgVVyAus13WsOsGCoMJDkaH5GchsD9hz56IETxvDpQuoqS8l+BPNJfny5W
wUgkGdQLLWwnc1SpHT83zbwDfOxp8e5yOaG2vXr4IQ/7p/Ixg/ptnPpjKM/dCDPt
xdf42pv3cyUCD6xvxVu4iET6vSLXClNvLDX+lCRcKMPgi1Vjl/SBwGVNHdw9TfU9
+5qGr2c1FfHlGdXs0Csfq4LB40POjP0vKkRTZS1yALATSH2UdvaERroRTha7e2Da
eOqTJpE1NbhSj1dCHkUq3KVwh/z1GgFTgUiMcJaFxwOnZOY9+3AUFURFXUYXZX/Z
oUvxsr6xp6yo/W6ZAeM2NYxHfl4Odioa5xfmOoSAS7qWYzG1q7stc5Gua0WoBW6S
3LAYoJdhxqnAghFIXbAcEPmJGpTUPhOOTbQqFQg4rjyhhJFiIWdudwMqBBWi/Y7d
sUBcRaNv10JFWtIdVQ+6ROC+p7Mk2Gg6BOMsQRjAQPprhZ+lbYHDDjjcfQ7sNny7
xgYfaiSr0xgnn/jwFs3byCqquyppCS1jLIJqbIBcvTc597mEXRLDpJuHGaEzWQr+
oN9LlCEUGlGhEDBqXK7OmNTWvOPHIRAHYas5e5aDqeQJ4Jfhdb0Pbx5DshNqswBJ
CHEkOakDff/6zPrgUQdYrFghx8BQDeDlxaHOeCLJzUXFz0KX+ca1hKlsxVjwoY/8
sk1fXUik0nfaBYCWxB5d5XsSK6ULQazbK5OP0jQJXkb0S2gZ0vE4buTXbJrc+9/+
yFJ8n4mrVNvaXnJAMcxrOvcV25KS9z3j8fAEATbDMHSjXLknRh0iDduH7RrEHUOY
8tlwUJ98wE5UW5iuRUu4eEIDYQ+igypNp+YEvOEr+0cdl54pne3pWCRTDDY/JVst
xA5L4HxzPHvas32yUUzn5JW+fOlqGnYqt72qRxGa+bEurKyJ1JaKgfM9ZAfUAIHT
Xn1fqSh8bjoGNmb6RzUjrF8dEk5QYRL+5PYqS4WGx/LpJWzDMRh29gRRytHedYT1
bihacj8bj0pu7mg/9LZYMd5WB/XXKaMP3CMUVxNcbLfSIwwg13fbVbmcFcBN2RNn
uCvdq4Mclavbn44kV+LG2qvhSLHXwIYqz7hPVDKr4/byRqNO6aTM6987GvAzuShn
AIOUNClK66qj3OLZrV4KroUrx/VQxF7FKI3G9su0/GjjfsCkn/uKCEs043ofrh0l
0F+jPtS+fs0sds7zrkLU7t5KcVcKY3vGV/NHdZO/J2oPXMiw7G56BYLwpQ2gAMhg
oT3cwGdRRcrgag5lLP9YDCCcxxMVbsJkhU1voOIMdGXXHBp152RlCIub1LUUzV7o
A9OukTJ7/jICifvrlI9JhNTNtnf38a13DUagNw3fOdDw7Ptz2j93hlKMvcAyB1LF
j6k+KGuA3rHb8RRjVNDTXODdlFURAITvagme5XVPv+mKFHM5ZIobB+SDv/jdVdaA
lH0iaCiBtbifKlvzGCRDbVm1Z/ApueL287VmhfRFgTEzpROWvYugRugmnVl4exmg
2cLqRyxjahRgBT4TMcrTZ1bsWFUOEKMVI0t0b4JLiBYX6JxFJdkkZhnj5nwG350M
DHM5DhZWNuj0ahDnFhwm/RWEbgHTR1/v15/4TvwzfDGGf0XjYHM/YW+JGMyAEkrl
F8kHiSQk79mBs2K1UqfgFg0tHaiAv7ZA2m6jWRcjcAs0Jxv6mpf6GDhzcPqeBjWJ
qG6SpImXrSCjIY/eZ+kwZsQ5vpfbt2/nz9eF1d088RSoNBW6xo1qFH2hHnjl73Y4
wXzWiLQw70jaquOwhJQahW1MroUok1K9DWeIKz4yLc9r8lQFCmWuEZH2VAr+JaWh
jShkoSiKDgv0XSRNg1LAnteZ77F3IK2JNce9wZFDxhovAuAfkMHbyJ6LAMTPvKSl
9XivQvA8da/W2yHZM7sy+XFx8V0IPxNNXUEv+yAvKgqo69uLHdziod3TL/mnAu1V
I2lYIm7BLpttIJRv2jACaKbnDDacELonDnv0TCCQ4r8rkKG93a8lee8Gu07wXEcC
BPQgiYsnmHLgyeunBnKfZuPvdaXY6AAFtta5vIWe1E2bg8savZKoAKGKBvVwTkAr
oFAZ3LbgrYc4U9yACm3QkxSF5wM5H+M1AmZz3rfEQ4taQB54cvNXIHblucSThxip
BDW/WhAcM7N+XDxQQvEGdxLZGEL5JpWlPEfaoxvFaTOgrn4GBaViP/1vEIO5yqsp
a/RmR/pLE+7trVwOsMnhN8ByhEbr2cdqZOkSM7dV9YImIH1D96chPxxCoPG38AOz
yA41At0ZwtMVurUTK5O4B/jxyMlLls6xZSOJPA79k6EyV2sksJkyOhg4ZEZ25OGy
JhWcf8ujTOOgE9GE8jgezjzgU2pDgceFwwSA12Q2GB5tL8TDw1pP3uu3G8PHYfax
au72XeBhOV827pa2Dae9ToA6wxd4S0sp+BXWVf/+ZiAf5AYHjy2gvB+djvIieh38
P0hF1euLNTHxi5tXigmPhxMMl1IdogtwC7pys7/6f1HpOvJyhOxK5o/+bt2XNB+L
IPOeIpZFPCgvQz0VijhKZgq1shfprM6V1xOLPpkzADQ76C1BKfOlfDgITpM09BVw
lPJ9BmNlD1+kxArsFlGMHQAW/9xSt/nwavQD9NvECPmXUPB/dwJyc1OrBe3jJdTl
9y63FcjtA1I5/9/zjH6RoeC33+MyZTK1dstCRR7QD02SbRMgcfOTLnB8T2DqpNTj
hNNh68Qw2r4/QcGipJKUK9Si48llWqvdfd6Mocsw3OV8n2C5F5oarE6E4rWilYLW
xHIAJ6rUf+BSCkEU3S/an71mLNAzje3cJA/daA6LfuNerOUvnNEBCy5va9DFkdLI
dVHaUbUeX0FFCdoUmU8lz55jQjUEfkV4moi5zRD16UfZzilAQ3nTn2smwTZWtmLU
FntJ8nzKvP/BYQ335pcBvLdnDJfe7SR0NEBFD8EzpwFBa3+Y4B8bvoWv42n5cquD
Ogxuk9u4d3z4pAJ9ztCBMBS1sHeNTDYwQ7QodxK9Te1n8Ws/5A3hTiOr23lNNwvH
G5kzkj2C+a0ZX2NBggig6DGa9CwhhgFhNNvn7kFlwBSJEsFrUtSxfuOZ914a2OZn
peYhTic1Ygw0Q+x9oUN6Z1ft6anotfuGi1OkjB6Q9ab5hNgEV56gRzp19V5d8xPg
CWKsQaz82s16xb6od1XYmXzcAW+AT+sXhHhaEDBzHXpnmcHeFSL8sbbPy9EGYDM6
VTBNZf3TPon4HJKQc1ZFoo5E3AOoDTA3Jn33HWRW9Qjyj52D2kqxeM8Xc/6GOXPh
7G95WQVkW0F6V91zj053gAOFUIT6hk5D+sVrbxT3VjwhHpxsyeA+AZgKnrJPAGTo
VLFzGpOCQaR5xfuOg0lZFEFlULJd7zh+9HO2gnOW2BkEQoB5t98Q5NNO4atQEzUC
YaN62pYhHYx+zCeaRW1zyrWk5/mQM3OCoWjvp5q1AD7ocjmfvF2iZnKgQX4X8r7q
qon3lUmgbNRM6/K0wjkIOesBzytAJ0rbUXBGNY29Yeg9JTpKKxJmTnPJ/Sus1CST
tzM44Vck0W8IN7ZeQ2/zVP+y8rfgs+nRsfs1rx6wUSW+Qh3dqzLWCbthrMUY5T9s
9Mg1vcWmpQosW/i/gRzYc67LxNvvKOWwNLXB7Pg/Dh5ybdpUd5OHE9fq1NubyJfL
REXSiPMPqjKir9xlu3N7xy99kZ4trvyWfmAq+DpQLDM814t1QKxdkNobe8eyegPW
siaa/93VHDT+e1LKdjSQpxanVaIfDPHSKWirSzEo4YbxowXlZ0bqcavtPhiQqfpC
BdiqzzJLOMGtEWegBBByIjpT7B9x5geGso5332iQ0oXJcZlDaCrLPhe12S3VAK5r
85gK5I1gXzVeJfLVsfAvj1Mdxj8PmwVB67NYt9m/1vZcK1gO2n/z1zRaiNaupOXI
WnKMS0qdGxpR5ZKXbcnrpykM3ySHzRyc9ESpKsLAeGVyij9uv/5DZyhV3zcjUUSY
Y/7Lv5T70Yst9130XC0rtnCXtkiU2XZLT7fT9+UoqFMUnx3KGEH90B+NBooA4wtY
T1lbh15xpuDjiysk7a8Uvst2/VOy/EEmroWgwoeVXCh2xXTPjLkeAmiS/uHbfIAV
/fMnWTcy0IlmRuPHzdVQEVo3/orC5VPR3wbGRDkaDV9gzwlSv1F3Ofkx9dShCo//
Ct+UYNOq16Jjhg+k2sXnWcQwxRqupXdqgv7zi16+rYN5n5n0auUh6cqFNShXdc4u
CD+rpSxz83mmMSyEbUfTrUgg7Ajy8hMG1Rm/Z6qs1D2geIOZErlfySzL2/8b9cJS
Vwsu3TfBQBt2CbwX5zFKUQSZe4JJQ7vX9n2NP1v1sv09s2TdIfFnDppSHQH2/9IR
oiUoTLYaU852TBrajkJLltd4xoSkH4XxRokjb8ib1XVIPo8Oz4rRaz0Io5s13sgh
3eD5Rrt0d1XhPpz/69YAyrre1y5G5fA3UeVHRFU2MsRhCBOEiq3rKLu97sAfRwlE
osdiLs5U+acKMXf0dyXXoyZEpY81BJZ7/Q0/cC4O1RwipSKsVWem3ufJDv/vgsYw
rPojD1GbqZenScklXyddyZjMTH9LLVxbw6VsmM6qCPcUZ573rToV3489dyCRrV74
LfzQ32+suwwbkOlwqghVCjnzxj85D8deA5unLaWoOa8rRNC2F1R5dfyIIyI0Ton+
XAqljSJTEkKV39fVN0YODmdSaxJ8QzoAzcrDCyoKu8uS3/oIobxbHNUAw/fv3m22
q7DrATAgn+FPNGKNcuPAHUR1WZohNzxWV6YgJdoZVpoRbOX5/WnaGbPwV4g4JWUr
lCSI/kBKq4zXLBNSFWc4AM6jXXMY5MNcgDCZaLlTzkqijYg8vLuttC/ra39VlmRo
2KWsxLXOUMxU/W+NPV1kpO6PK2b23Ok+wAT53Q8bEiDeQGHMU/IhihMLehi4sfAL
FTvqNepII/9EZwMp76Rr30Dx4/dSUfl4tqYnWelGtLE+ePn1JXXnJxbG2kaKSHLq
FcqseH90Z2hEnT5BbyKn/JRju1bDxN19VzdFfUCPW1QlKG4y7yDuWlwu07AzKES9
Tpc0Cu37+04l4Z7KqJ/eKFm44mjhzPwje6izVGg1JBRHb61mKyOA7ny4VlodcJtk
9bRUK5loWvSaLAjJfRXAgropXuXw2cMrCNlhOipnkRHBYeysOjwfyWmI5mposfaO
y2ZkAMaIfXLFgd9gpF7bFf3Fgy9fSoVNJ4EhmcYJsVYKEas63wieyAFZS+PTeqFe
we1IJ6UASoIjd6npfEqN5Sp23Lk1WYlg3OpDeXrYE2/SHmJGOoUllxoNNpM+G/CC
1JhvWA/snmrN1IhlqkKLculug2Vv25/sfMahyBmCabkY+KhzlOw2TCjagfk3dqBl
HBYl5qlBhV3UT4iVxb+nrLVLolr/5ZRvqbDu6uN9Pu/MO1BBE6qlXdMUboJJ456t
vHOKyKNfYmYJvg0n2SVeFTvyGcOaNkzhY7yfvBpxpOcg/uBLGK6pyqlZ8Vtx8bzU
W8jbBqa5sCGDP+esDvQrETkV4P31H/3xZ7qZ9q/xxF3qd+VTFpebxd9RVxxedG54
FqgC0gi6NW/2qeZUdxPvJ7mosYRF9jprYNWd/aoMbaL4Lms3oJS3SEdPB3saevop
trqdrPi6CAnWgBJeBbOcbeg9wXmWOQjQdpGmg/4vnxmVkuDRsvOPbglb5GPL1OW6
CV2jwiwBQI+qHCR8m8sSILOe+sqg0mVojth6xvXzcdNLkS4qpUfYx6ItYGrWRwhN
O7r+KuxzY2m1FId+yC/AhT6XXzSpgCdSQVATEekxjVo871BPhkYCvgRFOAB9MSJv
YH1PBvolj1yjR9N/E/p2TzK12iCJM/cPjj74guMzPFLccN9d2TR5ZHCjxYlhsQ0B
2N48onYokeLWV6WOFBuxEg/+SxMpVtbLfH5Egc5pGosK0TjiBR+mIDTotGYcUC/j
+LSGRTNX03b+mFdJ9tQ62WWKk7wmsckC3N9fgK721bDdjzIid7eMk23nbWhQpufK
ZhcENaSa1z8m3CPQi3IVFTs/70ge65ZEPjUGyNo70ByLIKxnfHFaQM0UziownRdD
cnrraduPEA21fzX6HkBvoB6q3Ge4E5fb4JiZZvtHdLRkCTE0i4QOJt6DcPw6evd3
/g4x2c3WscE1Ics2JfYHElnwv52Zg4CXK0ytL+Z48iTJS6hLXBd33x8/dbnk93tY
s0QRhQhbc6t+7ka2pOgVZsQGihkwAFiyyWDx/DMBo6bx8qh5MxQNQvOjGxH3LbU7
NtZdQ/q2fIeIWGFKjErv6OMiWmstz5Prd9zHc93j79CEHKR/rXG1NMukWxWrGvIs
w2gGJZs0yWJkNpHlRTEqt/9WdcP8QEtlohyA0uADElrYkh3ObLIu5TXrI80BdEWq
peiQiXmy+AmBN4NoxQpoBOHdi4BbOVzxnuaGLO2pUNSKKO8EvAwBLp31OSNk6VKB
vCE9nnFE/0L+b7048SSbvguvYJTMyetGVfKvZW5AsaK15hoiLRq6XBG45xiuQL/e
aKcSnhbjRk6rrbMfVTO5TM2+k7YxUBug9iQwPInOmzBKKfmMDdXzDUj4vOSpEaFH
5se5yNxzLHdSDpgQX1V+qr3tbyseoZ9abFkMoDJqoDGPhFOjo6zZISpnYAooe34Y
8Dj77gY5MZogtsa+/ooIbM5yv8J7NfKBrDwDSoTOvrwq911tIEknQ3nLERI9Ssen
96CHW2S/eln6wZKs4qIBWR61P+ofPHRY26WRfQn//WBmtty32eaU4CTip8mq/D00
G58zyE4B5MrFKHLPSM2quMcBw5ttpSM11dhG1yPi1PVHfiDSlSiwvtOW+BY/jv4q
UljGq6TmAZFiSCTjswhVNT2XMdOSLmJQcbN/8Dv2Geg2R0zGomcCgyy66FhCABum
MRGe6th70aBMb4Y+k8Go+vjgNxnyKPqiCBIZuePoCbWmNOyMRXe3WuPBkpSeiJsj
G2CaEq4/trOtdTmECv6+fiN3xXokCxENKRC0o/F0uF79Gd7vKCnbyXExaliajM52
lGrR+6v3QfAkfkoFGVqdf3auqoow589aSWAHYJfHgHktHXW6saOyAP5BDCXKxp+Q
SlQeGKH+0Pl2JZapHswI/NejGzjGdVFaCeC/4uZ8Flhl1ofMMg5+VBd3pW3sq8K3
1IAax+1f9Mpxsuy7OPWIUSLrBl6NaoiJYSSj+1O06N6viw4QeA3BPkq13EYfaJk9
om3RfIiSRMvh6dXSRV59E+Oj5HcmSTb2FQugEiFzYd7Ksuyfeu8XNhkzBe8TND+m
xHNMCj+DWXS/6zb/XJ1jHgDoTewVmSkxS7kLgBmlxE0vDplmWFCgQgMmC+OeRVpS
tRUMMSPbqVRlIEMCf6LjGef6F6z6gfTepOUUXrxmVmOMV7lSbDcWxI3XDaA/aYAD
6++76cOCkvfPTb33a7S5EUp8pT0yZJm+SneArRLiirZtXDUXuzvTJrJpG1tRUZZV
VVrsxOgdpdLpi5PgOtKiLbR+vcQa/0fNY9req7XiC1XQsGNyO91iVDztwt0NU9ma
NQkzthoyrE6eIIa3kXySxWFH7ft9D/ST5wddLuPBxf41UIEPPhZQC1FrZ1aopXgV
R4KjzfuK8cO0sE+kFbTAH8ns7kbndPEZ+9Ce8aGyDvuyIJhiQ+y1rilW2kLNWs3f
QlVhzICNvqMnYV0w2Q/Z1Kg6LG8Yqa6YR2RV/y6shrE0RwHSEUgMhsXCvlCrE/sY
OKMA9fQ74Vi9vl+/9jVou0jS1/RjVvs70KVNakLAEhFbas+GIsV4FCTGqlsDAriy
hRgFO7P6ywgT7x1+x37cO/in+dTN0zG2v2hrAzYcGkXfaGaHbaDMFaZ76gtlgFaI
9mQO6CWs8Gyz0j1SLJa/jQLetcWCG2S8q5unSOWV+rgsWh1NexNIw51Nt8Xoyfmb
SFOUhy6zRrGNO/sGyRPhgskZwd30DoBSsDeHNt4Q1UvVVLe3fsmm63BS5MF70ALx
/mWbGppov6sMjmf4AvzYh6VN8LbHDyC1qIE79f+JQaykZhkisowBSXSWhzNGAuQC
5H7Z97MukCPCWFMjBvqai04a5mRwbA3oX57NYBsZrKsm4TH143mk8/i73JTB14T5
BqKk7vysNWsUYBe/FPefE6LoQMzORLgq1MttBDNYyW5MbMoAxl6J7TyS/rA1V7VH
JTKx1HisKR2kE5FSSX7q1zNAHcQFDs90n9IID5B0uQ9Dkk1Q97FNIYCeN164MCF+
gt9oin8l0b//RfEZJr1zG2kUZVfsLav9z0P72mmJcP+r8IW8RitQbhF3qQ+i7Mp9
0w2XB5GQWrnL93ql3Aan2r2zZk0wMbfagRUL8w3sFGj3mm/R4hIcBXJ9V0to2VKe
QJImSK3Upxow2W/HZzw8TlphEFiETiSbkPhXVfB465b+yFpV0cpWwmY19+V2tmt7
nHRZwPex+gs3qTdXj+MPR43fQ5W6cdrGNsIXD1k4lUtwpqHOUusW5v+mG/mESgqQ
p9l/WnR/cX0uRcegE7Tg5fKuhIEK89RCMNLjG84gqtBwHx1HnyinURDgwNY1tuQD
wxobZy/9C0jIB1tOEWBZLAuiirTjWOohHoDWQM6it8Yv5l65wvVi7/kfMCfLlcwJ
++gsvrwdMqRWAkMRLI+uWG4Yo1hIQPFZX8b+TKpt6wEIX5xMwHau7ei1nE3OZDhz
dL/kOnwzAlxpg76Q4l4R91BeeTlMO5cUaqUqN7/NQ+SxNMJU01RzKidBiwTrS93V
am7S+wfkcA//NySJTSQpnKaccy9QWhCtnTLV6SExSlt6gY05lFNaL0ywl2Cmn+T8
Ik9SxOspY7COH+DNKSeoxur4IguNbJ9owt0Rz3lTkRlId6VwhSCKk5CfrFXjfh9I
0WWGvFBnBKtHmnffHQz/On378L6HinvZml+0jPmnpjCQ09nc7vV+l6FipQmgj05A
oUwXm7zUi9CGChx925kqn024g/QAJM2fdFGZN3jW8UuWFFztEawe2B4UJbXXhKBR
ZXd+6E/fTApKDxO+t6+CGW1PQuo5WaWFDuPy/6mXRoVFbpAkbXk+BCbdUK/XqIqT
kyAqvNTXoMjbbWwIppKOi+TyRURf43TaI0WhD6h/ENlQ1ZydKdijO67qk0ftXruB
y29E74A4sSMG1fJQWp/wOJvAc9ixRhI9QBbnl8wpDmh1VZGLkaNr+DvmzEIfcDru
1m2+LlRh+kSJtoj0GDaZ4x8wvMEE5EJJVOmu+THlT73NQvmnSjUOoIfs2ji2PFbM
WIVlkzSrGOeCAfn/9NPYje0mrVd6jEWo30xRvQ9KX4MH5lxmYi8uoK5n0BX8pslD
dxiHzSN3kmaHNs7mykeXbq/B2YbhgnuRNYZkM5ypQJz7Pd/fnVuPYbvMFCNLsMEC
X/KleT334YWVcx/ri2beh2nwawQswJBP0d6Agi/xK3ToK4j5laSm71wfxRMDS+3g
6ahZOCV11SuUgFS0SRaPB1NQBPWrv7evkscgmGhuCPiVBiepRpokOVXPb39MV17b
hD0snI8mpGgl3AyX0DV+yDEUg/L0m2axrJP0uO6PripVUU7w4Zr7phY9jTMzZ4Sr
5XtVYY3AAIO2F3YAoQ3dkeCv83g/koBA900/xWOfA1qAPxIv9sIysbk5JsCV4rF/
4PqG4+ct2fUPUqPTR5dYa8r5S/sdzhGM6H1LRXoyZ2a9HIaKvOk3P0GCCKQAQGrp
rKV8R3Q7CxutkbL7KiBHHkHrUUrs4uieZD0/d/fXw1Hv5uNkQRIKGsuV3Ukdr3mn
jAVWewM6LuQF8AM0r1wl4QBvUIE8QOZnzPKm8tVk+sGlwUfaTjgIWOP5AkCWI8sR
FqO3z/mQAe7LiyhQHeL3Cok/ekLM8owON2UdxXM/kGIuaiHOE5o+CgrTxWPobYmU
PJFYr1WCm04AKEbObOnOZrULsTnKNlghpkikPJRUJVuXK/WGc12wQemmieq8uMwu
b/I1KYDgUKQlz3UDnBAwv8S9ZAfYF1EjR2/QpUFlDmp3mtk2H5MewczrkQQPAraI
w1cuxlcINFRcv5S1uS5aBrpcEuKsrxMBQmCoJdWSroNIkSIMcVFGT6rOnbipeFN/
XzvcuTcnsTc6OcJcQ8HVNwAKdQDi1TRCT9gC/S5Z5Yfh1FksGq1xzCIz7/G0VMxR
y64ztqS+WRmeOiAajKP/Pf0gvAqzD0xorON/JT3KLHHUGVE+DskXJ356ErIRalE/
lB493rmFjcJdbtIx9Y05mrfIg2CIt5i00kVpbgpjTrVhlO69IVFF3TEfkbRkFNqs
mF3dAXVhQiChRRkwVcHF+uar47D6sVN0TlRlie8lCC6+7uuW/P6S8x5o2iyL3Utx
GW/5JEcTvABxsghFJjxilAODq0CNxzy2IXWtDpnB6eO9hM+CO0ZJI7DCZBTfFos4
CzcLMUR2TdA4NnSPOFaImbFmh2n8oRa2abfT/0CTSCdlyZp6qr4uHnTrmmEIgccu
kPHjoPaNKB+B/5Ro3O+TJWm2wRiQsfOIoVdKDg3UF4ZamALo1VbsoaiNgTGA0icx
nLjUgmJICI4jpQAZNhw5recfsaajV+asKKkAsdBYZaRDg2QEklvsueyy2bpSNkBV
cp0x7cm0FDps6dQQ9gATEaVL057pafnofQ9LJBOt6EqgwikezIuHX8td4UoUtL68
BreeKbjKMp07VBMMXQ3EA0Op+eC3CwnO/vR5Y9MTgmz/ldHARyCM2hwUyWL9fqt1
S1YfqWdHddWo2MK667WTEdrr1wTk7QKA33xJHE5WxcX0iINg+iStJQCDoXCJS8EI
sZIgaHUZv8avcdhgddcwpZK+QDCHuiG68O9hMRHyqcCL0M5o5OJS/cQfd+zziRXc
DNTwIVVpABwDB6OMboc+e1GRdxKPsV7nIqeofOOf5m7JKiPWGZLQtrX+46BL/N0V
w1nH0TW0hfl+ecW9KEYGS8IaS5T3SpF4b6TrPw825XScV3CoYXENVIWgJOwVcpDs
cmKg9Jcng09XJHffN1Piy4DkWpHDvyb1+ELGhQLgx0VArUX4ftBydF8hV/CbNKdX
p5NWgwGjWk6P3BE2X2XKz7P8x1Bu/vmdLnr16Xh/hVf8wiyK2pZh0Tz/NCeizErM
Mqm1HbDPgPs5tc56Eutt3UuDLApAMZXMbtjh799I9qFh2cZ1amfYmMn5U7wNROrr
VWPVjRxFy7Mv0UKY37Ncv+Au+2FtfovCb7oI44oSU6l2aeF3ZX9+C7XiZpXVht3c
kjl4GTWG4Wc55z2dzH1Jszl26xnG7U+33WMd6NH9546ueNgVVr8kRO5n/N/NJLWf
ARhd2k7ELNkURNOnjdSToAcjYPy8F+QW6xP+dpscY9lp4BAK6qj7mTmyipkQCT8s
3+YbYU8T+UFBcgpYoeysHLUlGXpYb+DB9108Iur11LteedODeaRC04qx8KAT8LSi
LPP1mq8PZC8N/XuYnGCYIdr23pGHjCBQRHLu5Kwz3oREf4YNkBn/x+AFXa7n0A2y
XQA+9nciac+WaPqyOy7/+0FzWJcK+SAn+hLsoMev1SY4xrrlkBGihrcPTIub1q60
QHb2RU3BQ01R79X16h7E2dp8HDV8bXrTiFsnXk+s+bUpZh7fD1lwyURTr1vypv+6
EGAFZGq7ZivQYxybAU9xJwn+aOnbK5RI6J9QH/M5ZU7bUHOHoH9xDkFIu1+Jhdzn
twbBLeCg17bA0tgKnlCkTr+wWRWOqvCTBwKV2jQFehr/YoWRjmieLZhiYkBngcQU
llJbFGEvCE0nP0igACNm9E5417Da+d5SHo/Rh/bUVcdPAwmnr0ZU1FKZtpyZe9mb
T+ZyO8Ov+WZ38iAF71SfBnrYSY4qruISv1lyRREPLKUKpIEqNuDSsknDrWvmMRU5
6tSLKW5P3dS3Dy1a2PJDdjKiOgPwCcTm5Eqf78zaIMvjnamiAzTjXq0vEVe6omdc
N1Xn+W1Gj2Xl1op8GeaENxiOqUhaz9nx7l2Xc5wMUZu/c0SolX5D/SEmZwkxx0WS
Xa0sOkZUcXyVKsbkgMn4EVdirI/na9r9pgiyxuBzMfD/cLRCLn0GdelPrbA39bc4
/l/glRGN+LzsYo5kizX2GKGvuTd1D05Y3D+td1Uy01RzYROIh7aHzpwPuAuIy2d4
EcpL5IuQsVEtq+wa5aL5z5ZBEtxXxYeQ+wOnRH7gGcDESwdSxSk/q/qmTxNX26ZF
3vDlDhTF5wtZy0YY+twxjXbRV0I5ckoUZhVOHkGvKV6ZQOYzZzC2QqbKPMbPaQm4
GkTVg4YBPPoQBytGQEpT2jQnBRjDaInN1P/oA48bpRz8Mkq4FrGypGcWVHlTurUP
mk5pd5sx+Q6Ckz47RYjUzl+bm212TShNqfbdfdIGaKk1pr1MQLZRVBDmSxhKZKmq
yxmwTFNXaITvXDPbe8HSiqXG/vvaU4f6J6FZAf7hoB4OMvyO87LqjGjyXCHfwReX
0GUvs3dZNTj61HbuXeSLdCFYgzfL8PJUJn+GmdmDp1lpQ9sibRkh5oYSCm4AubyO
nr7h6AjgVDof8C/KG0nog53/wiUpEDjk5pdnjcnky3nvSOI5NEV709iaVkOJOjEJ
J2si6gTFUr//KDE/sHCBEQlqATD8P30QNSsBbedW6JjMbA8SltOhyUEPuYzNDvYb
SKxOZD3hGALFhtYf6hKO91HGWmUKPP91Juxlilt41ah7dLPaYTVpzvRn60vGjZ6a
4il0/xM5wDodvW8eBSTb6SuNZ1XtjamRdzhAuWbHmtJY7DGn5rdb+yaeLrfuLcbJ
uitJTiTksTHoVszVeOUsthJd4ATdofioSE8EO8uHGLunJhiaKvtRb6olnfpjnFmK
mVy+oDSCZffGsrLNgL5sK71YALFZpJkYDu+NBuqQA8x80tH6Dedfij9y+cDzWwAI
nRR7N80NPN7bJ/9UyAMDLYBG13ZVQmLCxEF86vB0hIu+VYklfz3y5EkpFK6xYs6b
Aa/cS4Y/6DmiqKU8QeowdrGMF/CWLM4m3CCc84IGE2zxihkhqVJ9K9NKGwJ8GZuV
SiOHDoUOfKSHiT4hC0r8if/wkiuROJiQXmvKlzXUuCzgRpsrHzsuEMgu7gj1l2C6
P1i8dT4aqcEdQB00LA/6YWdL4JWSiTFsQodFW28YnOR3Bhzr7mBVhyXlft6li532
m11GOGPVl0RwLlsN6sUI56/0BifNzUkXxjK/wRJGxmD1GkY4mq1EGD5Ko7gA5RAt
89a+yh4gSfMHXNT+C5qJvCT37Z9JYB/tEnvxkZqPfNg+eH3r7LCPJRwxptt+6fsr
A+Eiu5GjbCE054PR02cKLqCIwoUsgJb9h7r0rriY/iClbwp3tXrPTy5TNl/Lr6NT
IJV2+iF7/T+J6GlW7TxkGCk463CRyp/giMxFuNXi/K8JliOLcke0u0AzJ6veTxi5
e4Hv3NeKg4XvOTNuQS8C7m42jvmfmImR0rt7tE7iuCJtn/L3hwrQOKBptes7WByE
5NihRcNWOjSgSWKU8Nyq3K3eDorAx0VSCyquVgC1+Xzj1x+vaf1/6Fh2PGVk9t99
05zPJl3kC/DyHNWSMbSTQFMZIFb4yBKfKDgZbJEL3xqedKcRCVj/4v+tmKL2KYSN
rXIZxI4SoeXLjUcQQ8g5cOi9tZCRgrYszuoszcWQmoPAG9bEen1QwU9Ii2dYb4pS
TQmgpUiMaW/il9qNWSGrvVNFq3fyh0hCWBP8b4CuaCZ7RImZ42IN6hfVG8l1pCAK
etjtla2xLJxlzWiloGHIO4+g0/Ni+QOkHrzmwUIFc7hiRWnlohzbOBo+ZIcVOYaM
QdYGqk5uGH869iMxGt7aNaghwt+/5B8mTMuHKZe7TfejTR22v9NhaX7nYRfV3fmc
jtQanAHDA2ATCMHJQbyTpskPCGEWBGMEbDVyCJ90RzUrf0l7v/UhmQaaa4CoELyk
EDtwu7NKXxEApHRKu0SdAPhPmFgMah3Z3f7OH4yxuNFcCDyHbULa0hVtdspPX/Nw
eEumNp59IdLr7kVP2d8boxq7MQqyfYmXPlTf4GCanh1wSJPjQwhturrUxx1/vhSv
MXK9+PzyKQ6/Fpn2NRgqKokqnRFPfnl8rpOXxKe2X/2IsBvug3ut6qcXr3qNa0gu
47w2GidqtG8Pyk/jdisyTMRR09bULKGWmybD4ByJRU2nd+/THNE0ZC4hSvD6tZAf
y8GGSg82lZCo+4LvwfSIzNmxZ0dIoUV1cIuw6P2QcmCoWf/lsJXiqCSrWOr1pJT/
95Cwp+Qdzdzt1gd2WNnVXzljiCbWf/fyv9MPkpYuiV8wEEB050N6MX+Q7vR09bov
j/2SXunKBce3OxoJHNZcoyFFVu+9OgZHE8/WZcIgH2I1wuIJ6fdYRtTPr6We0wHL
C7wNGZQcNzTcPPB9Zg2DK3fvUCMAPNAgLEF55asHTqyZsVf5Uy+NcVNmi18hswwH
bYJ0bcy+FzIcdc1sLP9KRBgND/drMQDw0/hAshEb+8zvVNTNbjHIUT0DI/MdNkZT
WpGGXk0tqZXTFqQlTXtTP6Yse/nl0Lx3V8fwVZUAE7iL8bzzV00FjLWbxLmpj6hf
pi3ZBX3+QkAtaLQuMHZC2nNwLtDIMwJDlH6p1miR4rYhpXeO2pceqDiFE+ft8VIU
st398rUZsVWu8qJy57fxRDX4YARQ3aIxWpONdxT1leKR4l8QMQLnL5DDhbwfUHgt
n63WzfiFwXPgsJMjpgrJVQMLJXeOe9+Ta/GhudTyLl1DRYk+NJ/p6EJhf7G9hWAa
gEDIYHgGDEHEPfhspJqb9zC0bq2qfyLUWPG6J1fqUQEDQAFkaC+ZHf1xabQmHfi9
6mOR4A4QjYDjK3JccRYXXyZS5TD7v45pIwGSFbYznk7jnJtffJDc9XA6BpIdr18j
KxbU8x0uqeQLn+I26iilk8hRFhg/Sy+jsNgtHrYhcX0XaVX3lB/peozQAQvfDEoF
/zy5nzMt/V+3wj14tRnmJoAxzFkkz64UR6ejvgpC1vmZoAHJj0yISmzoI++LNcSQ
TzWhhyUkN/+Ym6oOWJCPyMARJbKhFc2YSkMIAWizR19/WHHK71lJ5Up5fGDDG1gw
LBJ9+YxNZTqF2Bs+AfBlVdGJwB1zWrEaYW2Fg/1iAxbt82lqJHds6j7mItEQi/HL
kWs21Yy0ZejtpWG0TymltvGiDrW0DEN8JnFt7FesqPc2ZX8D7FBkq99RbpD3B2Wb
lEgQzy2jJBAnpnf9uF7P2HHGAVk4GVBhJYnpjiJO3+HM+cROvu4SqRp6BN//A7gB
qhrR66rL8OXjtQL1nt7qWU4UrwZkbnWo9rjWlYZg6oKsscUEjtsYKML3t3J27CVd
ZY3BxRjmy8M0Ya/ykpu/YBOPmb6PC1PCTc6RNrqCUmMl9HnosH2WWeicVS28AZC2
z81/m+8f8BZqA+bKD4VPJD+OSbJBYnyO8GCiX0yYBOVtIbA1GeMG1+Jdb3QnprTs
83DnGMtU+7/ltMI8O3qZCVGMtSs6YynClok5GVWpI3GPzQizmwaT1LSbFusqXAe1
2a4h92H7g0v/xKaCA39FRH6nKXhklkVk6b1WBs2Jz9S3379m7zv9zbvX2EtfuAyv
9o+Kgc71Uhnap/vA1g5D4Io2qs70KqbxvNaNp+QWGZt9Se004KJXs/+8W0EFIjTL
b8zzvdeEoqQErfkgeFYN8/rMvTHFnkA1HpknVONfMkA69bNeqSzQ/pvE1JVw8+Zs
DhpSnD1ooyjJb/lGaI78c6DBcErHp6j5XZ2b2JKjEl4QzerBJqgNUC0j8mrYE+Lq
1G+z8uloFCsClodmIum0VRfFCu6JkdncdTiFKHzA42TPAQhP/AUST/rH8ssCqnvZ
F3mpEVrqD4F7Brs3MlujXQOhEQVnkmIYW2Eyo1KfYJ3h/X++MWV6zHJ0TZnUaoFz
fi5KWuCt0AnpXvcbXdnZuXJTXGTkZSGPs9QcmOqnyqX72T4y1B+0t7xmGSB3KpcK
uaxa9k2s8VlrfLi18Yg+0YsrkyB4GjeDJAulcJZ11iRc0xIXxLbVlsm72pb35kDI
DiFpGryjp5+Uw3uAkEuuugaHeYjb+8Fp2xrFEsx7PhiK12JosFBjOcGJAciTpQAd
RLWtmDcGnjB8f/gVXTy6iDcJMRNMGVrtF5MVUwq+m6OBkFP7iVMKINDowk8qavd2
2Tjc5bGcSQ5lJ5MKH2+MW+mfl1Y0IeFZHqBYy8Il9QVkDnZZti9989T4pPg3yf59
e2MkJDb3SpDpKU2CdH9uHUglXsrkpIMV8jGQ6A/eDvKWUtt/R5jJWbPCW9CAStt/
crDQ0dpvmcHyOT7ZaAbxDiR7gsvUzBkqCm7hztrmqg9vTJWPwp8T7yYoYVLw1gNu
MLwLAIWjDOHfHEefwc52pqte9YpMbc0aAhE+sVhvleKLzDJCNZ7BjnXIwOf2+SPc
vhjeY+oCjQOlEToo0TP6QT8CZCpIiv+OLKIWI9qN25wCaS6d6N25TG4hW55YnmWr
NoTwsiu52H4a/L7KncG5MaHPk4OB8Q4o9Z3xy9n2EGvWn35e7ffyG82xPz9tm3GQ
keiVxDYMikfGEqb/73xyQqLj1/E0CLwZsRNd++VPrCBUCK/kXhWtqGRCINB0PYP9
4GAWavI3B5WlBNSaweu/4nzeHQYtdb6Vz7RSaBVLp08XDKDFZbV//Pt9lWi1mdXw
5zeB+XywDWXJqFaaGlw75eoKUvRad+dsqlfX3vfHWESwgCHnIOF5Nse8RWXZxFK2
VCVQE3vZiLn3UF5JkbA31JLHus30lv0GrDX6e0WvvZYe0obo25IgA5QYIs6fF8NL
K6/hVcbIMxI6XgXS39MRgtWf8jeqZmwcna8EdB5LLHW3jALBIFv/Vo6AlQKlSLS2
PsAcd+HX2sSie9o1y/OG3m9yDCfiVfN5fB2llay1KKqNUo6N0uXtZ4mH3ERlQzyR
8Tk/8rUf7uCYnX3OjMNxNi4DbGW4A/kUIRV3TpTjBXFJtrKFR+q2Ib1o10VZk0wv
Y5+heAjwdj68EDcXtB/cskFfgAQdat61KoH37YMvDrZX1yu1gO/L7iGAGrOQ7X8j
wqgvIi4UDtyArz6rKikX833Ml51kBd4sP7pQmkP+3/zh2xbpFAMuDCkA5ocIWczP
2YiP2z1AzCEp+L9DAL6iat9m7w64xuRTSV07VRyMiZfcqry0Pns6ykyiMCldFO72
C6Aq4GFwjeOpf4CHQOLVpD6kh8P6pF/hSVE0JFxun/hdbCiMZMWGUkAa+UYBcn4i
XmZN2H3cBgCoc/dxJaB4nSYnfrkXrl7IymBW3/vpz08ZymzwIbVHI+bNMVOehKVs
e6FrIGSnI62SPZ7QS3M18sMyYV8XI9meXMYIZE6OtERdDsz5mHKZGAta3pDpHHu6
/2d7yImYxhSzEfpx6lKwgfUz3My+HaHD2+Yp6XkLMTihohYcblQXZ7h1t0q/GgtO
udgfddxXoXrap+jhIZOrvvzU19NPcoldEi3P5sn5zDL2TjNRbRMjX/DRDkQHbRuL
DZ1VjCBsAkTS88qkfRVwoW0VK3A2WXe1CTEcn90Q/MoSMDLcFFFGA2gmPck21lLX
BiWOsNQ2UAqKGlBE5pNZfHVTDZ/yk1Sz3VOxu0u+Ap3kuscSazPZnO0sK7J5T8KG
39Y55rFqGBzWmQUNHu725lYF3D6Oy6Tf7WnMJKh0qbdo7VN7Hq7mHTY+CaTzyanz
ZVbaM0FmVy7t1xcBTskjkbxahYaizqB1sLYiI5HMySQwSB/zH8wHozsknv1YMFWS
pDDnmD34xK+AoAqGjS8P3MoC1JGV4ks7NtUXCcy7SnU5rAIvfK2A7fnyG7+RwLL7
dnWHlJ53VPx51R1bgEEBSq0kzcZ/lZMnpJ2o6jQMqaD/Oa2tpOP37sPJmncqFqOT
w3v9tbfE5ZEDfd1Tp49OtSvX52U9jR/lZ0ABbQKgv1vMaISN2pujYItA9Zb9cbsQ
Vf1F9i4zm/yjyeaLtfbTCJhnLeU6WyySS0mJ5wV5VopTaUv6lQNwVDdNuiJxfM/B
Iw/qClC4sMospmQZHK/WhBR1wKW8XkJJT5Finxs1pXlsFtl6mMhdA3jq4BU/EhsG
vdsgZaBOHuz5z8PN4HTOHH9VmEo+XdrPztWT+JEnTRqeLfJdQyztiPc+dGGNPnpz
LFxFKMHSadYBZnCnqayRlKRokm6/QEPZ+93VhLwZyfw23Ps9w7WCn2JWFEF2jJDm
hnySQl9oUbZwSXGD9x7HibqcnaYSktVuUheqcbiBSkcYTEHFCqZT/exL2VmcKXOs
FYg0ky50RpIEGOYNzSJLipQpoKsMiAZGDoUMJQHOAaCLhXBnmzc9w4tpIhA93nPs
TJ5rlHoL//JUSoUnEY5l6HIDLBsTGnAnXu1TVlfSY1gqdPvqTVHr+w0AnZDuqIXJ
YE66nPnz9puE593hzxIuyK9Z/NfnZzXEZq3jMrzsLWUdfqVucvNEPcykL6VfedjE
1zp5niXpj2QOwZK83vaxqaiJx0VQkOkuxTdnS38eeYht61PrbusBYg+jG1LJfvDB
5B9q9f6kU4fjQYngZlU6xqXXCyzguN/5W1wfk+qkumIr94lzR2Q6upriYKkPmDVQ
Gz9WuHsSSXsdiLeA3gDK32Zh4CSkzG7cjTRwT0uLDXmws0yf0KJo20HU+UmOD0M2
68ZwXooJ8oPCu5Z7UJssZbepxm9VGjWuj6p7A9yrE0Tz5Fgum6snoXInacwX+C2t
BFsbj5IIXjl6Sr7Xq087BbHOwgaI1RtvarbP3UbUmZUrSAtffiMrCOFfL8f4O77o
Ta1A6omxQLSXcR5T4KWhtkWKNg7zaVIqRSxBF2UkCNz30jUTFjHaRg6/rRMnRK/x
fYkEQVFTMoFTLHpIV4UEawFNXy/TSBnnoWAki7c7vHLMwWN7a2BmygOBZt6eNQ4/
MJLtJ/V+ni691iZXjty4Y8Re3ZNSG0Dtq62ePGuS+9SbH/Yo2yjSPrpuK25gK8tE
bmU35M8VFjwV5NanSghvNB1GoP0p9GQz9/cD2Fl88cv3yeWam/DG5IZJSAD63eJ3
Qm2LPEj8R6N8bUu+brdnezyO3p3vjKFCKbu/Ii95jNwjwsqM+qOvW2wPzzOa53F4
Hh0PEfpUr5HvVein5Q5R6L9ioEWAqFfnzaZZr7tqUuJxSbeBpVA4cW6b8pZ+5j9E
0zQ0rehbIlFIG+MCyOR8HbQUg0+XACd56UAnLgLu9TiRAV7x1Wt8W6vlsWX/x66q
RMVZNrvbW89JUyMIB2Ql1kq+i1chMU4BrIf2vju8cmjMohHt1FWq7ISuO6SDZcC8
8ry/G1jElfOYZj7+pxy8Uy0JOFaJDaXCTuGAoEXOs+Fokp7w4NJJdABlYjKlNTWE
vhfFUlAQ4tN7gDFkyub/KmyNTkfLxxqKbtD1gNH2gH76dUg2fP/OZ23TTkagkJb9
ldWL1UXp697iKDn06rNKP73m/cr3Ae21NxwKkKswoxNBpzuvIAFwYBV8sNdE5y6R
3CbOjx+jGEapNB9RZIIfeGJzIy3LVWnO4+/Hacx6q+kNcWPRYvJkVzl3/mB2jqzo
SUw8pqgSw6lWUN9ylfI9O5u69IO1Xg9Mc5u1j17OZXkHTiIf4pZ6y6Qc6CtRm5FR
nScg0F3tmDYimrXhL1xZ9Pu6NqZXwZBy2veBxNNEK/Z/oeUM6SXaJwmXhzXuWON+
6DJEeqvomUJoWi99XAju61XZHxidqH/hFGFpNkp38hQkIv00PBpptMadH6l21wdI
gYBroc41deUrPJ41Xb7WSpM9/RvFwHn8PodHO7fODxLfKvmh5fTtJmQJ53jzESmD
5nvZ4iWFtZ/SrbNWs8bPf6n64Hu0JeFwh5oyjcAsn8kgj00qm2eFYNEaCKE3qH4M
MX1fw0+UAVWonBDZfZiwoPW6KOGsmIFn/2ifSx+UqnuAaWvLi1nLFaOJNO3wJv9I
9AZENd0h8MXFcEOLru+Ok05s1LMDliCXzVNDXf9OnVwLAe2xoQpF/L7DNffg9y8C
uI1zDFoKNwoiosyha862PtdKDurrMOYih13PXqgjiEhPtC/D2+PHxp6vQXWt7MOV
yHIEDyMZfn4iqczT7XzZei0mnYTD4Yqa2NnqH91jmMxstuPtSH9CiChm+yjv08pR
xdpHNBrJ8BDX7hsz2GCbH7OattpBKUUfOhIE0s42IV5WJtT/JwZfhzogDvnOcJrF
P1fsyodX/YuchBfkZwvJV1HrcxYzbf9ga9euYZ7PTysTFXBMPLrwf6tdEK2xOR4s
dLFufH8Df7LWq671vQcKE3DeNP5MuDPSurGIcLHbaHvL2cnBoocE1JMEQyf7M0qI
DsmzerBYCNn4EXUy/5f3E3fmbogzVQxXmQblA1DOR9rmxnOPr+vuQrx7qkVmZ2mB
ztGeCeQx9eAl0zAI4QhL9j1ThSaogRPjbk5on/O3oe6i3PBOyZio1GrpPW5cooK/
0C2E1EB3mGeEHSOgdml3+VpSrhF2xtb5cVeXD+80mHQAcJfPxPrjtaglz5YLu3Q2
ZcB4EhRfLDR+xCOCWAcfRE8xh2Lr/7P2o7cS4XZwEB73w1u6c7kAoZVGxA11+7PD
l3236atmsaIwFapceMrISjtESlBAnucD6c8IjD/wLWiQuMAItM6Rww0JZRg853hx
1Wqamf5ch87ly26S16cZ3Ha/N5ED5SYgaNRD1ruC7mqWbnUmbBRliP4fLxAT111R
JKPg7bzHdw6rBkd3lPze/byrpAis+pDWWS6/f+2/oDnvHVduEVXmknciJkTjsTwo
G6E6uLWkUYOmsQh+TVNnxu/W4GG6GybzkblLijPBTQcNkI1rwF2Y6gU6BvFep4YB
xlIPvhAe/AsHB8AhQ2OVMGerswB8C+WC/9zUDGNfR91sruR7KiNj1E6iETQS+nn1
aanX4PXvXWUiiNCOA1ayGAV37Xp9C/tJljEL1N+k8Wk/WkZAdRyJ/xs3xYo/Lhjk
/RZ8juH2XSYigBeLf/tmZehoMOWdXDYtfQaGAq7HXu24Lgx398HlH/q4j1FXocVY
BlLkV6NXkzYIB6j7YTXvYNPU7bN9jdtM5G/crgOf3KmvBXVlxCS+daoLKiCAxcbE
kQq5QINfLyR10znmqHDF5sHujTzRVJH+0DNMzCSbLqvJukabFytxvQqxDLQTpMwP
gd/2Y9zRJVlq63/KECml7BRUQH8C5bcfqf5GhDbkNbCKfjmYrS457MSfbiMd8kEI
ndvkgyeGjtao23I40QTBaEVKC9MQGJwAacpSXM28ETNy5Kh3C55HIVp56uFcapmQ
l5G39Xq+YJNA9+Bnr7H2Fuw6poBgzoUCf87gnvSqUCyUJtC1RZajZfeISIJlDHy+
8QerSMYwMOgTdML6pKWY/nyDhlm0aPP/R88uevNx4FApc7t4ieT6ydvWpj+L2j7L
whFYTMhJCyyPexnI2+UrN6x/zoopF6qRHRxS5LeFCMZ7+dZjSC6t8/CbSSMAM4Aa
uvtoOcJ93JEtp46p8R4fUGtxvo94F0t6LnI3kprumsz4Irg6zyF2yDeujye5mL2t
4FBEslCijuuGVPle8it8LOSeD+8fpw7Y3SSPAmUfNhP3hAebpZUgBkOw29xT4oKk
IWyfeN8E31ZX+BM1Hx3iG6IR7MKI8YOYjLPtK9+dYO8C7jB4Kb8/dkeFzViFnkTk
/IL3FI2Q8rpuHxvpXNjIH6gNm225gMPJzNBLXJKqreESbdaii1zxQCru6EhYIm+s
jZrMFU+IGtqDa0hOpifeezEfFSr5ko0irPQ6HdbuTEK8x7BYwoeJA2n83J2F2WvT
/Qd7VLcdSoEJjySpZHRiEOjf6LJqNieLgnBPO1YKwOcsn1rojuk5icZ5ZWPy3a4k
6pKJFEZeGpKly8Wu0PXCmUOBNky/NnnP1/HmkNiXtXUmu4KlNEaYgVpBzRNs+9gl
fWJJWbGQ++TdeuOGWCGoHYheEWTgFnDgqyWdnrKA1LkWx9JeHwfEbReTs91O6QyM
N7YSHUUgj5dmNvT6flMNLq4XkHviz6hoI45ji1ilbrqbK9zvBio9Doh7BjcyR56n
Qat6jfPq3t/cvBujTYgX9g+RUDU5IdCizFqY19heF63RkClvviPBxOh1p0p4yyQX
Qu90VS14f896loRTL7gHz3B7847w7Qq68XI9AqV9tI3pUMRMT1DqGGQn7YuIF9lA
8XwlYpVr47eP8CJPf8gx4Ba4FV22f+ITKMnYb+C1PCnwbonQyjn3s9HD7mRENVKQ
Px1bkXM6XZOR4FpJK4wZ29Yu+KmoSypQFNjmufMQYgFmZ4yhWaVtrniwTUhGcv9u
HYlTOboasD6r4XfQlWvIDhr6UAYsD55x07/N2EY9TNjtpc1U0Y/V1kVJAmEV1Xsz
KHuyKY8J89jKsI3GVu/HBer/oH6VQY4lln7nS9qbh4ZA8J0LM0MnH7FL+wcWCGZX
3NFlqR8PBdPQ68Eqd73Vp5QyQuEGp8gUqxv8SSDCtKycGQeaGUuyjJ88sQPJF/DZ
N1b8YzLeggnK5KEoIqIqnpqyCpQ2l3rPwT46Lj4fycVcsjS0ZVGZpGkq87hWm2qo
oapmPnYzHZAiD62TYA3relbFE6nca8XwWdaiJVATWuQ0fGoDG9KiWtgtse2i+pUi
kWYOjaeFB6Oe1WFBkgX744vaZsObCfOoXZFQVrY+lUDm0g+PS9WXve+mHL1Mo74B
W24MF4DZ69Jc0T/1f6TuXxdUktoDBk+eCAJk50NpvcSZ5XpvuAzr0Fxs6SeiYRy4
LlIc8o2wHzwhQNHaVuNAwAslGQ/FZjaqE/h9RSiITxqlQNYw1wU7RghqACiwzakj
kMkZ3rnKltg+V2+UbgfjllogBOiUPZmS+/ppjGuZHhudHH6wDzeYHQYGTlFymttk
3mqgpAQu0XHg2F3XWUEhDuRCvw3BU8pRuCXKvln0kyY3GvJPAz5J2tPDXxBAvMZe
05BN+7Nn6+khippaB9knzw0f3cHH3X2HSPZPdI5hUMew65WfFYpgUPXqPiVPZj/f
TnTtB952RFUSh0DLNJ/2DuqDhUJuiuczQw9JeMJ9WA9tpvkoBTnhpPA4yF+ijsAR
XNEiaqBwOvfwTPa7ILffPKc2EwNsegBw1/hVe4BjuI1waGE5hnHHbBrL98+ZVI6V
J0LqSkMngkn8xFSlXY+0xOtYHAhwiRJyJfGeesvYOzeEuzMy1JissZRgMkqmnvwo
iMGHzEY5+GIPYVHCbmeQ2QiIhRI5rvZ5dsUQm0DLWRxS4onuCo0l+kGAy/+VOhVg
D3WR3OZuIFJ7hH3F61+N4pw5FG2axJPo0X25g+rrxnpgfw6KbNB6/F1OX56B3mri
P2ROSxmlCd/LKLIX4bdJOpg6JDs/Uas6ccnhAVcMGgM0ZEc48B1sAYueUsePKYBw
YmAaDl6Cn8G/8fuGwM57rm8Eh3z+njWWamMIhNck18n+aXYRq0sxG8bqYOQuO4Iz
fHUnCusTi5AXDIDBhNLKwRLWtzEKR1mIT9xtcJ9y4HtfGlGQxtwGWEYqrpLJS8Rz
ZPTVcyZqAYaLM/zbRtsnh8422EU7lTiNyE78uQA2ZV8IsGgolE8RR959+grkddvS
8VbJN+fl3hdhAOpdL7ZdViy3u8DjbSMsUNbWT8/U59CVhAJ4kkZz0nyQetDDT/4a
N54Y7IlONTqr8lL5rVMPKzMBHXh+/syka1264h0q0jtoijAEUinP1y7mZTZ6rhMH
VVAT7hKSCvkD5+BAe8GY8NFlmOJyWQT7FldmCcaGss0jaUMYq8USakOmvexm/BKX
ddk5MLeT1UKrYDaqbXBv50zeFw7h9r3ofhv52zkfXGbM8HQv45PSn8g6xIvf0z61
SuiqyMKjexhBNA43Lofifh5FxPQ1Jvc2WaD5MGfW2DkBoMwcH8AphBazndZrqZA6
8Bliz8RSV4FGa1qWv5DWkJSfuj3ka/ZMZMsRRRmihlfnXlOerIlNfXWpDh1bXixP
O7FErPvJhX1EwOzZXPl7r7oQU0Lgz0otl4PoqDwfkJ5J91EMHD34MQXv0X1NXel+
BzgGl+wfgHL3enhT+C3ybTL/+5ATocU+xgB8v2b5zhoU4sX7MJ7OMfjzcCUtofsT
i7OLN9TED20gLpQOCRZvtklv5kWwZAd8xMZ66BNmbBtglVHma/Xmxur5aNiqx6mt
og+uVpLOXHXFWifOsciMtfEmjm2IUFn7ofNNybLQY3vItGL7Kq0BLAT6Z8Twr1mT
s48y8q8UnBmCwq7Dt83Ll8oNuGlOVo1KiFNQuOP7KXHpTOZOO4ZqsZHS7D7qh2Xg
/cvygjerz2i8SztRtfAtz+S2uKHlks2knfUUa2PF1QSmmZuAXE9bbEoDyMyStM82
mlXl3/ezue/HpGy+8C5KCbaPGMMp49l1nrHiQ6ag2y6aG8EWDIndcTR9mQCReSyS
2WEKuS+e31kF3Uz5w6tKfn7zeP9OsIeRj+eqR7g5276nKc4PRrT4AW7BZSaU5Snf
EVX1Uo8ksrcIJfDv37uZi5dyY5mXabIjfHTAwrNMdPSJFRu2Vy24E7RO0Ph2zETx
MFI8affnfWJylC0u5Bhs2okIRLcbFBUWdpnEzm6CoDE5OHESTtZnBwWWIDzYzeET
HGutOlJXjtlb4gVEgehBdhqTXocU3AiDRxo0pAYdwizmwrfYjMLwzdceW4LfVDqz
CHBaniyUSEja8I6FKvOQYf+e1NWkWBqEFJWrrC1smq9OfOCksFKnPfirIDhvUxLj
g8tk4kH0+mS71j4pUgDvW0uVaIRSzy+92rwmlMAmHrw/8rwqtXcCbrudfqbZ2aKd
+JYtMcvt/UORN7ojC4TXUEHOfLGDySeINXewtIe+b37mC+W82A3UwAUAuOppAueJ
EDwAOoCVKjgjGvjPamuWKXqcJ2l/RaOwWFQN4DP39VnR655vpU4029kUubLFgQpS
UiaLJV9apvVHjq+MYVBPPv75lvoGgJedWDrf4ZIdLb8TCEaiXSK6BFFf/QBEOe8k
Pg/oBdc4RgktalMRDFIMjqSzRkpqOKYFFsbzYK5yNOGzriQqWenSUHY5txi5nk21
l4cVk2oa6VmwcbYXD2FwFhIYkXW8pR20ACMDa/1vK8QzXvJqUQq7uHipQnarmuxM
S138sP5XMmKxLpNAq4hkt/366SIMBTVmcK5sW1zcdcL8oulBKI02Nxg0NYBJPAuS
d9FyVS1NvdF16ue2/vta8FO0eqvi15hTbG3LGvHLEGDJxENk8FxaAzMyfPpRetzF
5BDOVwP7MUCOOGTlVKWEqcXp2cfSTN/nu2E8FgX6iveYnE7Y2eFFqtbWPqOF2PgP
A2caYhph6S/h3STMnM9aE1RDg/LTmPPInAhUT0ALhC69GLyYByg+Z1C/Rvbsl1Mk
FrsfNa8ltyRDnGqd9CxKY9Ho5Ll9xVaEjEIzVqWhbfsrIG+VL8Xe/4QflYDoSmTN
R/KtZ7qNZL6k83XdE1icYLUg2qhkDMumFxeUFxjciTTjCSecfblk5xCfJvk/39Zj
Yd6zGDHCfJoA6+YRPA+/JyJ7EHJploHyEof0/WJaJG1kil+HLo1qfnlSGdNPJC86
eLsNU9MNO0qT1HEy/NVPliUVpcxPrzF9IOYAL8UUBLBrqSKE4bc/XFcC/gR94r7P
yZO07y0MAplSAGTtqFMgxsU24vTrCz0I96Pb5figfLEXC5BIMfiKTsL8GUrpKS08
uE9/Ei1cuM3HY9YYU072WPYU+JFWNfAwp1a9q/g3KXMcaAfCh/H0rwEM5qZyJks0
qgkXy2IBXHfPvJ8lhezj5jCiNRPddtwxbOd5OTouJ4IlPK6NIg0gRdH9ZTwKuSfp
HiNdV3vME1c5c9jUQSc7ebhObE+Py1vCI/WjXe35FcyTrSwh0Hg/ehR4Hpnipp14
+7wubw2cwiGVt2bWUcM5PEUei0QWIn2YJjV/srp50FuhwRYlO1/3AzA7YqQ4noxy
pZjUMXKzDYfAz5Y77lf6UcsW357FPqyXZ+0BRtfD6jaA73vJdG1SQ+kAUiEmsy4F
B/u7xzCCkDPj9jpMfYre7lYHe/5gZotZAX0cRL1gMOtc9BkcT+Ac/rjV8XJN3tv/
5quGz0WtS/NQHq0CKFMET/shutIsrVbtiX1/OUwhWWFkk/TWSiMLfMvllY0hXyPo
p05MM0tnToDSHa0xBQ0CJOd2vAoxGB+7MPOspjGrmFdn4nE0u+5x/o6e+/qcHYlf
T0War3I2c/GUiXUuM7wY/9nQVt/8S/2TdoE1wbsSEheehLHiJL3fZXXYeTy0VlGs
DDoWxQCBhWIFnPPcTPXVFN+v0K+TuqgzUoQiU7D0S3+B+Jp2mqfsJz8b5qkTbBjY
saP3bK685sYQB/1SE7TkMaGhrAJQ17ka5IBW2YUPnmivNt9gjZoF+fvNLud5F09o
8Xu9M6hLPx0RzyPTlAFlQYGRyWMwVOfR41ZesQ1cILHBbIWfohzF5HC+6jMU8E9s
5hVXpOM6W02k1xyYbIHlH6X/vq7cFLT0S/Cz1Q6go22N5GaWQzh5rqm0zIbZ/Wah
QkP5WRgZvf+5Q9yF2sEOfV+y3SH6zqRCArJnaKnVuVT+mPZ4GlcgdpGCyBLXHVpK
c8tnHXnF9hIv1aHWKUREFYTr6QlPC/d8Jsj01LRXMPgfZv0myqWZqkisCiCaJ2A2
VOeU4IwnZgQITvnDUz3aO15h//V0DzzA5BXSFXLUhFCQOvJ3LrJPEeHiUhOo7ckL
w1BoncOxFKZylmritBA9FGV4BHJ6cLRzCgWZbBK8CBTFXEHPRFzEjyMBvqGusrz3
++OAk4PmV+e5mA8roelDqX5hcErUKzfSLX6O+5cpD/hEuB+151il214iF+b6homs
F/JWhx0Ubl3g4P9Vh+vNCE3iZBHMzi4IkiMm/pLrm2ztlPwraDQvPgb6m0jqYZp5
vjoFeWiOREbl7e38kBT1/BeHKcg0y9vgDCdAfo3wxkFazIvWvp/o5wSjB/48Kgms
uOqfujgU3Q6jsxCDjA5G54RKLrvcDD7YLGZFRF9bWRAlqGu2VTz8Jga23SwxkVJy
cGzBY6b8T//AqbVsJaf9/iS/lOgnFilO+f8cZboiRAeA/JUF/rtVk1YH3DwAuhuf
e2jXZfIa6rh8U5660TDslXtuRxeJ7x0Zi+ZwJjWpne4X9oaY0UmW9yiXEwlaetLW
Gzn81QqveFeur8CY3KsLzgh19ELyzxXl4iXLcfv+3NtYXXHNZcu55slDkg902O4J
jYEOr6ekNuJWbBhb+0Br6tQeatVJme7RGiVAQ5Jcfy8ecELPj2hvGCdh1eRYE/UJ
AZDqU593mt8W1wS7NLnLRSEEYP4gUcC0j+hNhdTAhrVKiSvkoSfFyCFK88HhEigF
OywRw7f2JH1uKLU/4f9LIQ36uIBFvvHMGy0+jq92RrkX+8z/vXQGUJDM/Bn8Ar1H
gHOQJ4Qj7qiraDRl3nYPGhXYaoYfIjK+x44hkHuQMixKFC0akqPgvwdp6xamlkZ7
c+g7e0mQORBV3cvsLscTFX1v/VBAakJqidKEIqqyKyIvAwVAhr8hpe0HtMxxsIXk
axnnT+VNVxvpZ+dvCJ7XoN2gYPastjvhLMmyzOnU1zh10DA4nJB3dGlNRfyjpUaO
eHz6Of1ma0fpINU1pQ+R+AqobqEZdHyCMNnmMj9zPrHq9y2cHigY+BFA6fQd8aXH
KDh4grzgms/5uWw09s/V0gygMUiP7KHlra4L0aEY+6Q/hFrO/X3BOLw++PkLyNje
CHs1ujysLs4RYLeRhAC7IWLz2M+5nbbDd5E9CTtTqfzc62IGxcJQRsrgPIQ4/ydx
4syeKSOGS36MHS27iftJeZyFDcUVx0EJPPmJuHdJOjdiIqMS77Lt3If+qiNnKrrn
Ktaju96axE6kX+IB/D8B4QmbQbvO21kdagVzII3ku4Bq3+G6vp9JJuqkaLvc7jH+
EaGy+ka40vQOFIHXqO5rz7qC+BTCgEV7GDea8EorP0aeGVlWBX8P4fWrocsHBh5J
8nqO3dOQlKJhXD8unRWK8TYYIf+G4vk2CWKdycW0Ix6LSmZAmeNTjn1wuyzBOgci
xogsrWuIlvy6HEMcf6yXFvR8KCdVg1nW7zPz8f/0QL1sWtiWdlu2vFg/AFq88cGO
tfgdtwLk4sb/RdHc9W5nDPWUOixjWuGVspveCG83mUbuqmLMJNfGnAYsPI8j04O2
1t1bqoXe6bJBsoI29y5C9Z/i8Xwk86fIOhwwhu5XhzsAmGtTYObfV8aBKhpR3xOO
LFxVp+luo7ttmnvq8bbNRJ+ILL/TcUBhqjFM+U9Z1efX4M71NQiJwDODGX3Yl6kT
XTLivwU7xoZZXgGnxxLYTXtEUaPnW0tLJFk6jcvC4VzQL8DcTUvQHSvnO2OdIz2L
u2aiWaCHn8lH4iwFVa7DPkwI870PB3fjqNxf0zH3OWLpoPNMst9ruJiY5zppQ3W9
7WthUQeaY1H8/OEjWEsKUNb+/UxXJJak5qqKApTTrcrZBUyK+7NYF9LN1offNgvC
YP3JTRGba5liP1NzimsWFkdApOlxNedfoIBKrZtKnIK1RvdfBxn2k8XJuUzUNESp
dJLnfboFluWNZ9Cetnv8N5UN3dasnKjMjEI/WDzSSJkUnVvCIP6EquLXRIo1BPhH
JzR7K7t/cZ3YotkRti3+NYFEtcaZwIr22GnnAuC2SP+bclRjn9Z7NJRhzIEwKqsZ
qsLOgOkeJHH/Tn0fYhtHjliUTWmMC9TEhb5ZTmJqZOwFZa25fRumSEWqF/HdMbkf
cLuBEnRtIoMATVEKcHSHWYSNXgWA6AJWKuu2OedR0JNf3+Bc2OU28ZWEPq/gkq0o
cGFC2G6Xd2QwbCMaO/k5aBrH0pZeoX4ANNJ/K2/nRXzi6dfP1v++mKYqA3fg3Vtb
FRMPqijZI7oRSbArWmYe9oPQQdXQOqkoDUoeXaLvoH5GusnDnZ0GTj8DFN3N8g6s
EFY74ZOzXhJ4uQLaeax5mtVqbsSv6HRWtuJi85U3+OjZP1Ho6u5rh738PAxq77Od
VC3P5ckhOkk9xkujNELSI/ygfe71bhCNkgXDJiLy0qeOQEbQ4ThORW183R3mXIa5
viNq1SwnkgjWOtpn9NwxF3DVZMEkjFe1HR0Py0UVEiFjooasX6yDMQDCuEI4/Vpq
9KFK0j+qb9cFSnrhNFDxXaYF1hRuHi/xsk2Hgu3eOzZtKQGYrAOYLuelrQlSnxXg
qhvlYq6voOtFyad5ddSeB667cLrCwVC0fFg2j45OGIBy3XDS13jegxtfRvkB0phi
dB173Z0pRk7rtVtfmRKzukuzrRdOmuXUtH+QUmJWDJ9g41Arn0Nw+jNbuv1sNkc9
cJWp3BYoyyGU+t9upbJjmW/zU+mvYHxOOLtYkBUdBGwsOC4UZdLugksrqiQ+bSRL
lS5kGefx73MMH68JF+afjZ5HYQho5AjP4cVlUWz3TZgHAjVscqp7iP+BlOENbKar
f3KAMo0TI1efx7YRd1ME9kunce9pIxUKrIIlKCrJj39DGpKpZAzjmvYLNk6ehRt7
W59JXDaw2t+bHCGeDGDi2Hq92cna4FlCqCNjX1C7aPurHsLu8V0YHa8Ev7S+1uA+
iJAS7GoSGvD4AszHmyvYkQc4hQyVXyZgM+i5tpSHaAKMf1frAh6WTVK10NFgHgHN
K4MdQ8KYqY2SkymJcnpvMeeOQxmDhO48Xrlz5UqMQ6b4RntpkNdekQjy7HZ5oUq2
NDR5M/koWW6BPKzw+yS3Qw4sV1jbBQakEbr6no3f/BzfNnDGXhs4bRoX/m0nHjlt
GXWgttCjbUrJ6oH7KWqe5KR2mD8SqT9m7r6hQVq9BjY=
`protect END_PROTECTED
