`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1KxYhn7kgLuwuUPHlpec4k/kFKnfuNeILXKGI3a/e/4OjE/KaCmbCXcsTc5j/kR/
xDblWA0YFfvkYwbzQ4YaNxJeSQaVxF9iKLP0RBoHYY/xHLzdcPTMB8dqceojGVTT
6Yl3heqxFczn3wdlWpfdjLysIIjnTIJpfSrZ/Igk03s=
`protect END_PROTECTED
