`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bqma1zixYItNa01Vp7w4K7wX2UlQhKSvMcCnuF17UkziSNN3Z4VKNL1sIkdNUuIP
wg4rEjizobiRwiVOfxqR48cSY+/i4wmf9Nbh68nX1ylWL8UtUKEDWzTe3CVQL482
Yw8Wf7jJjKI7KiFEvM60/U9iAuUzzEmZowrKgOkvGN9gx2e5fOjPH+3qiFwjDZf/
dN4CTqxbjZq7sdVeCBNEz3BYZbtDVFQdQ5tZ/OlEm3Bbhfzo6L8QcbNtxQM+gCXf
FVYgumpxDuWBE+1eg2bh0RO5mCVlRPKqGhcDJR6+s8m040tNyBVDUYKMK0G/KLDI
CSoj/OJPbZoTvhoIIGsNVJwH4hNBqVYKOITSQ+Ltdb3BW/o/QfXalTI7AtP9WQuk
loag66qLCgSvuLgYz1PpEe9McvAph035rjb4hcBsiZ5RGm2bRrhnmXjD2D25b10S
`protect END_PROTECTED
