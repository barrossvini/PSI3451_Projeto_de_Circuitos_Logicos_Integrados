`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1lDI4W8j5ToH4WQcfCtVo9NYdRTCCgoFeJ6o+MAbE4fnf0k0hgiHQRzFdeObkFIB
QIpUTocRagaFy10cuA08HntJrJDpJtmTqw0mXIRWIVw/KdLDggjJZVuFeKWKtWE/
a5ccAYndyapIAYcSgF5wZjWCOJXw63sr3PivN8K5LjuwVY1Kx2UNmTPFmX2qImVP
OgvSBz+RoHkB1+fOB3uD0QkOjZCzlAn6Fz1QXJVdIUSDchTNcM94ki+W5EnYrqIl
S0VxMvNP3TQTjreBGfmM8CO5hXzYZNrXdBSDrG1esswes9TBuynEMRdfFdoYxDRk
vNFCLckJhZHYs1MJtJnt4+lPf+9WCYFoxrRaiOx00W8MGfQVIp6BeJG+TYYjDEUy
lz8UZlKi07xLBUQEZGI0xSS99HdsDFMMDaq44slaV9+mDz8EtUCS26KtJsuN3Zh0
QioIS4uaJiH6MEP5V1yYM6KABk7haxl4qNQD25MLnhhf4FrAF1kkV+fe5H4kJVIq
wfYEO9EWb3tUGIX43FHttTjamKeOkBSpMoXSE2jMCRp2Coed7qMcLKf9VtOQRAlR
NvqzM3zH2QLy8jAcSxmE/XPNVCo5eWWxDXOkTPSrB84r4z2gcJY51Uy23aTRJfBc
76qhUuVOAI87BMoUEdRrlKX7bdSFjdQZ/ajWY7+2w67Xj8FOlDRzVeWdndCglfDW
651h+K0BA8mIRVrfpntj3kERkX5RoLzYPdg9q8LJOqTuLCfx7+cm1P5vh+QelVa4
k5M3k1+/GWIXED/tgu+TlMzgkWVo8ACgO7461fqBSHctAFQjXMHZ6quzsdZhw5DF
Uktq1Y6T313ztKTav+UQjg==
`protect END_PROTECTED
