`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9aoI0EW4Y48aNGYdeLsMKtP2Rd8PmNMzsqwlCvseNQvtpUTQNw+s64+JuXRHfcpz
KJW3PAK9Ql6efsbbvGKiFiZ0E8qG41o3TkCljqm6MyOMpK3wVviGoOE0cL8lUocM
9Al8Rj01V8sCN1qU/wAGQ7TST3uqLccKLO1lHVKtp9I5AEvGMz2SC+3/j75S4qqO
hpEpuG/Bq02BYLDcCn+6LNgAcBFx3ZqZo85P23e191jnntgNIs3OZ0Nw71unPGub
3GjsnEasHW1IaNRT10UuDeciwF+0TCUy5oAHf3es+/mHhmdF/AJ5ShE9YOkrVWm1
6oLco8tmdNnsYBhfIRqUuBbgUkyP3ci2dKyf5V5XQNjJP6Ori4gQ1hjMawbc3cDW
2izQIneFtsVrMVdLF+bALiyLnyJ1CcGLd1S8k+vy7W+Df+cIJQbjGTvHEIECQ5/j
3jBSVaupTnFI9Q3fr7YGrLB0hQP5MEquGHTAcI5TA0Qd5CErz+JyCZib8QL9L7Oz
2NQ219eB6z+E7u/5rP9q3+SJwikETgWOiDNeg01K9I1R7DrVDSpG3pAYAN0J0hlm
C6c3Zk1pNPt4pB0yE3/EN6zcN8KFm3xLi0GSTT0eJwc=
`protect END_PROTECTED
