`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LqiBVaCweD6LKHWVKZVgmwt1XfrSicxQJBWS1ItiHWs2MdZoJ3bQRx6XMAPeLmQb
kIai8WFrDBEUDAOXsPmu49NflTDTIUJjd/rfz6hOBcATnfjEBplf1NHOcMW0J4zi
oTxCUjSPjBLOEwXdxjuRv5ofTijIHOvY7s1IT1BtDGRzaM+1LNXoaBcOxx+xTKNi
0TraNsg7Au10ps2NV0zSG/21YBQlgK2iGd3T618xiBuX8ekcp9BqJhY7jCO0MdPu
8lcHYHPG6s4AgGt9P1IKi9hlf28UTUxZov0jGDMWx6WquqBkDQ8Y1bYBzeM0+Me2
afK1TOY5hUVMmgat9BnuxA331RgGULdNYDHvwxVUvCBKouoSq9gUE0wk4Sdz1tWS
hj+y+E2Xbb9ssyY+A5+NOAwwT/t/gHSk3mPHLYk0DKdotiiaNSC3cXrw56cFZNUc
8nYK4YbLS4cWJ3+bciWM0MvVCVaDygK6v3bCa7qtkgoUIMsF/rfEvrS6cOXbFwxX
WwA1yF8HwlUvAZ5r6DhmaCF4/1uojyBlb85/6ByTDbwk+d9fcAkXol9RCBvujzo8
/5LhAEoF9ouod44O/WB/WGJ4qOpQ1vdu3WWdB6XAjVmgEuWw1rro9WolnwHxxvQC
StkedMQbHDZqlJngD7ZzQ8qTZNRIYzf+Vguky7GZelMuGfD0QyUnHY1IOFoRLf9y
22jlN/dNk+NEla/FbAEj42NEPuA/1i7O71nqMx9AwrzCpyM9aJWPn1/jWY5MgxyM
mXHP8eGRyu86ywZQjR+Y91Cud9265m5i6c/p/s/n26NpvYxIA7giQZOsVuCJTObi
eX6sBIuLFzCOr6fmjj4N13KQ42GoVI1aE4WcNYzx4oyk9k/A4NjlKkQongYtb8Sp
Eh9LTwcxqS34rxMAPToM/a1p1HOlyYH+3Pd8JlLxPOudTSOp8DKHnL2Pdf/Ws+me
Enq/NuQobspaHsNiDqCBPyTY7um2tAMllCT5CHUeENCxWaWCitSDjYETpHpYLMOn
aJJYocmPApsl18pZZojVyDs9aoyF9QpvxnzKyr/bEOG1LmLq4A53GmQv5yI7uOz5
4gsRzh/oxJJx1ZAgk3pMz/uuLU9AREkm7lMbLQD9PNuPXg1HdwYujEJGQukzFNUw
jZTLy57GfRbr6N/i09Rf2hSxwU3ODV/Q6isu3FfUC6Xat4KzexRxH8BgJxoAaPCQ
9K8p3R4YOUKHA2ObdQo30O+WdHjaC2A7vNTYDqBmQAapo9lIb4013Ut0dtiaAKxD
UF5NtJZxHhktFGArm6C3RuK28GG0WLPoc8+PA605gm7sSheh6bCFO0rEL48XIkfP
hGSpi8BFrC3TApTlA4EGUmUwMgulm2WumKI9dJHOIEq9mzgaTNmM9uhHTZCN7PP0
CtRP4JyQO+QeieHzC/R146QqnWXwQqQOpO5IkO3zaK44CvjdNK+DT0rUb8BirJ5y
RgHAuq3jBC3aHno+oYkcWTAvOEl5uOkbzA7H4FeXGwz7fAqDC1NLkq8FcJx7K4RB
4Udf6C/SFqbUsJmIMGrBbVNaEWKEaDepopfn9JOzgra+Rbab8rfRPXLpUuH94Eml
RxZlxNCp/Y6y3oKj8H3hHTsN/oAK0DBzLnS7SogWjiP/7mlhiorkm6lXMkI8u4BF
cGZrB1+B6Z/ZoDG+0EWi1neY2GS9Fy2IXc39ZwOUwgAS+ROww0c98RBa2Pu/QaGC
2XC8hvRse2HHFuSceAdCJ8GVvNPxdp4RbQKo0D98e0dJeSQ1pEj9EYlT47Rzxbeo
RmvR2rVESrkKOpbTp7XY16Qo8Y0aALgaYCixXwu/ifspLDEC1m6ICccKmn5i9Qsb
lxFhooOhw3y6ydNwj1sfvceONnw6BHzX3r4e+RVf9oJyCVK5HWr21TEX+v45jPX2
ErhBBw6YnfdijzJM6kjSjt+gmfNB/rwaSelrpn1122TwYlqnyvNrX9ehcT8PFKdj
MAlShGGswVK+FYjAlBrVJDRHzTegISwpYMlT2CIvKkpqBxweYyR3RyOMoUqurIOv
OvSBFac6e3fq0PTKjQaCBLeN6fSzIkTFyahge/m933TaAqC7P2YOamxlzxHizjDU
KI9mnFRAhi83jm5zYa3aLtLiMWY3jaJWAGDsenauajxYdyG94CSZG0cenBI58qKK
502r11Ael2Djhh4Tf4ByNAn9nSj4nxhDsUUGHuPo/Cf/rzkmwZxwo1bQM1ovmN25
eblmpI6baKzPT72NkcXFl+5hZHS2RZmAMjocUFSQyYASBogOzqlKK+hyGuxXZMTd
KP+jBfZQVz5Z72iZHqeT43iPMjDCLVpAY2//0cXlUXccdBFrW0dUefllybByg9wo
k1YUpt0umlHRsTrVNls8P4jdGGuusEcoJDgqxcjf06/CvZNuz6nAFXUO+XFasjLi
qffjC3htWuoFO12XUAjZ32O2+jR6mSKRal9WBbLiuNK8b0UwPZ80RhR3edbn3Yxh
p1SRYjyNEgH1dxZdZWjamNNSo7x97ptJh1txeWCfAiVL1yfQwC3bwPbWBWAZ+Wzt
Bm2MT82mcuhod658ReTqCfzgZfENBn8E5V8D4A5SsvHpRroiD165dom0f2grJdwu
Tjx0LHFT6+GrQH0hbuRe+jzXbry7P3aebYxocnFu5UrXPiwbNJvoa+lmlSerTkrl
2Ufvy1ENRNGH9325W061uc8oSquvR343BYNsMXG0YlE1BtdPvDy8+Qkcv5Eh8ylP
e6cC0cI53n2fwVo7yBaO5DKy3c3cqT6NaNHMTK1YkOyJTJaqIaeqaH61qebkSdie
z/8Vgv0ScH0hiL1Cpj9vNEA8ZFxF2eAh+CeYNDnAU1IUopWmWa07DiJjzDXoIz7y
aPB2JvyTTppcilAVNwu5PI6nt/K/ixsp/fGFI6lABfqazUgOf9u8fERNzY8uCX6E
vBZjZJVeGwGFknvAkXLxElNlGXaoM14iRwqeGMGzOpghiLXE/lJ/gkTd1a//A3BV
1oULViF4WGZ/0R9Wo4PqoF62GspDNOHh+/oLquA8QEwWdwyqQxOSYYkVA9fQAHci
IDfLClYT/TIrtqrBRUfKxmIar7/SkMaRpMgo6Tlc1ZCbw9h0Mtp2l9/ozpSj+odU
p62YTPEzowPEUTtA/jPNxEQQFt/qNebVP/4rQV5k5jeMu6EHGIyAH0pRBThOGNwG
GCyW8QHOj6ttG7Z1WloySUy9RiU3WL4xFHuGie3+GDDyivggzfAWy2ViXy51IyYO
9VMeMgNQxnNwY2589EF6hS+DVpHCPI4EazWI6Dx5+bAn4AmlU6qdMxY5ykZ8MDJP
RooPRBqiaXdOS22mspdc50MM77lwQXqLIGLaDK5BiQ6AwOrfHAfCM4NMJ6WLxqyz
S++Y3f8G3dNAZ2rxy9Wv+yqOjcy488V+AH6NHEPab5hsf0dt6XILbUXcascnx++I
pVsaafSprFzfTeHOvimg4DMVLqs7pC4WMLic4JeEG3QS0ymKl/MishjJOH3N3lmm
4v58txKPIpCOTgLkBMgk4A3Y1VIXS7zURzvheRly2Zy1RfiTZz30Xp2ffLgkcATJ
BBeKL4J/KnSMti2xsBEeZtURsjR9KpLJlqqY4yTj4zUlKjXQ24IRwk2nP8v6CG0W
V/V3ZpHWAwj+1Up3Cgd7bcW++bZlXIeiqE9gKg4pm2BKoRH4PE0y14sNw2QL1Sdm
oFIEISxY+pihb3u1XY0dLUpr87nl+9sScOIOIQnElKk7K+K2b6x9rvuy/zteVV1E
OVJQf+h33P3diYPgXq/YypM+7LcE8ejcyZZLmTfPjFSwPAgaQVYUV9ceFj+j51ZO
GLOZd1O9+ArehU8nYhs8QQAJn2dxShOM0jRCcGwfXNVYRpw+p+cJ/l6Sn9Q1hYT+
H3h4dExeBxDpr6VfPD1nhdke+JiqNpOWNSjydkgQXgyla0DJ9nIWAAwtZFJspOsJ
3qBnDmCfhAOm/bUXU1jANew3ERrIM2XR8kcyhHEmJG+07IWZH2j265pzHfWrIHs8
QYkXRgP+qxmFrKBNLytcX1/IX92PULM/ha//LkK4v+ffJbqLGYcytkWU/KpVeoZj
wkVDNEB9ed71r/i/c9s/MClQBvZ9jAPJuh1Lkjl//SWyywTHvgmuo3PXs/aep25m
FTJih5rSre1eMGSVPvsazLD0QV3qYjHxLL96sovr12JGeMD/NDbx2cIsqRCMUsi3
q5iRinjfvj1ee1W9PL4Wxx2ieWMkYByr0M0hl/ZbEGmFZYxF0d6ctbotxYt+Xgkf
/FkqX/DCO95JX4nL6Txld4BdmK7wBrrah8DYZ47JyaSYLyyqk98yMc1DyNAx+tor
HSAoYtjVK9wgLBrInr63scQh5r9btKrOHByL0jp0n+RVX+S/edrh8DysXgdWUa+a
wqkhIkHIyGtKT5yvQk9eeSiaYHlvj9VSrpvTIrS4wQN8RWtOAdDHw+q2qh27UtTc
lReiywwWOJBaBVrQicheJTGcEJbizC6VcysnFZk9ngSe1KtWb2IotN0ddFqpuXUV
iN+rhLO6y9ompVYMoDFA2LgQyMirvem8AfihnqWwH4JKFAlQuOhJFDByjN7cuqHi
WHfoc36z+Ok/UWvCeTFdJZQT7NcxFMkJ1mmZ4QGqMJsp7k++nVVhKXJeM/MSkzy9
Y8dadLH9Ix7G0jS7bUm+nsgNQxZpEKon7jnQiV/5eJRKIZdiugDPhaSYWnUtCCrr
rqLQ3SX/9JJMmasIPx/SoJ+0ZHrUKcX1E/0JqnKwfy2WATZ3qCsISyW2FA2yE620
iD7RaJQIRyD4+5Po9l7Ay1+9zqEb7x9kVDwCIHI/ftEKoVjzsyBfLiC8w0ivT9Vu
EH3hrX3eDaiYXj2Go7nIIBawZVEmwLlnP4ui0vuB1w9+ZuIjoPsR09cXCzE3of95
v/qDG+KeUyDKmtducqJhg9SL3pCjyxdQdfw9bT+budeqMU/iwwcqULSDY5biYWXF
K/DY3HgFEx/OAlm/z82jHZWddEMzgz7OkyDBge6iaBETqvbaMslZAxKK3cRHK4pS
PhwYDeMxfY2k1jEmnGP6WeaHsB1IlnnTNF1aYQXgqYKA410utZWLrcKXr/G7xLwB
gX85DohYFfryG/4QauDsZMAnsvhHVdKkOzJp9u12bBRuYWc/2BiYM3mhOpD3sRt1
GvzMXlcQde2rEOy4C9LvRMI60vevRAvKEgSyeXzwmfd9CdwZwAr3UccpPmX1uXVV
ZbN3OZ7mKgOkg5SQoe9Ak1jwyKsBSCF1d5TQUp8H7IoK7+tIoc6NOqNmFHvOSXlK
2+LStt3bWqDAebMh+P7fMvwoq6lFL3nlaUfzEjNMEq5qKrfvAUpzxhbMqnDzOUrt
U7Ql1QUY4RpDBRSMekWYso6LgIANarN6TkymDouUYVQtXOPQFLTzUYUbgQ39f/w7
fw18YxdjjujoRuG8fh2s8xWPQ3R81C0mrKlB0H/2Uwt1s6ldRPxlA/c4M1Rd/441
XsAELngZIjUMWtvUROyPULhnh6sVXGe0369aPgBlPwGAehwdTJb+d0ZucGB3IdvV
fhSebpVzbyC7KQjKMNblEBZylPw6IhGXEPf0oBIyYOt3QqXIjt33uOlJ0fkrMAxY
SOHfWAKBYfjFDFnHQnNX8zq+7QC7MbJR1/lAoVNDPYYtP18/WUsmNvKOk4KucTY1
k2Zz9XGWJ6HGfIdY5wuDrAG27g3oKEPkc2cQpZia9Ld2p5J2TJdvt45OIHaSYye7
nBGFRUv5We4gT5i4JhuqTOb7HfGsJcB+hv3A6z5X01W/pISYm6XrRLIA0nnQwPQC
5dKvFkp8Y7mCv2REe8YEbTyyqDMu3Vj4Y1bqug65xoYF7Qttd9/kgm1Z8QsrFTfV
VBnzn5EqBSLSAIuxC5xPwlgzjMDLylu5Rlf6MPUBtHanEs7n1r8nz2u+w8LCONc1
4I0VcXZTKnsyUxYVe+9IdZyOTzRR3c8Dyzh3omRYzXtXn7Mcdc/vK1qM+rsemRqC
uswhm/RVlhJ4RF710pWwa049hfkKGjDSKptXNwjqhj8Dsee27jP44yQF9AlOar/g
wpiD9xmny5XWFi3+S4CuoVPcApKexC4WacOdsSTZtZiKLfVFdknhaDa9l1oTB+Lv
oK2X9PEJefLNFEStVmKU9CwIq+AyBp0oWccc0uLlmhfdAer3LcVDgU0hnJtjLqMw
wyn7U8d1oUCdx6F/Ns/7dBRJJuYeefhgxyiZorr6o+Mjta6+xsAKMdQXAE2mZ6Z/
SpvFr6eZVm3pu909WYQf8FHkKx80PKZ2H011/u3qe4qLRiWfGb0kflGGciSK/vdQ
xqVozTUz7hil0QZDQJCkqixAmoIxg5j2hlePkA9KlgRXLGMutOtC1bg+cudetBBF
5xpfxR76Rir+et4G0KKNshJdAzsugGa9cPBW4w7N2iXfZjINEtUCJn4ddiRpzkgg
Butvx+6lxfdPGuXYIP68B3Q7gEkFwOEvNxsbRaxWoKYrVBUfovLNC/iC+bIBlBRS
0sBdoOqs2GE9umw6VwDQnGbUc1UWIeV+lDWDIZBsBAOYeNuqX4MFbYAv/AheivlY
D47vxwVOdFBfss6aSNmEU9lc9IAVGI8pjaEbkrrwBnGD4qwrIbTp9lGWX5GuPqgF
/c4GD0Iky6IMWH6KIEw0jAKoeBh38NHEnPKIwzslwD0QiC5rghasUpX8Yq2wAQ+i
jr+eA2t/fLF/yUFsGr2vzmiEf5uTVrdnYibtuqHnNm3xmgtKs7V36xTCf8eH6jJd
C8sCJ+9yjAaZL2zcXD2a6O8GrFz49Vm9VzEPW3E/YGUjn30M7AGtNFSnQwD1qMAq
U4+002tRtqD7LnLk63uGOIUgVDl0fIIeB/ZaNYZGjqBjSUV/v8YoDHbw0AfznxrF
MbYKqrpVT3iOf++ObOiz5jiMie8D0qi2vdcZdS4V7zDGGRWz2yD4Aocvyom++B65
YZs0eoXfEk7F5MWm0T4ChFueX2CBvVO4d0o7Szh25FjwscwR5vObMtoH0KX31Gu2
6rEH1vYTy1AmVHDd9yEexswF/xGKwzriIRXjCMa4E0JRVQbak88AvGRfjFv4a0Er
uHDX49mFnAxHEQ2S92F9hqtwIExDKd08vCBgCrCseAOX1OalnC77L8Yosb08PpFK
OuyIsH0rjD8S2xfJTMjwbGfBQk78LTmD6GUgdJXVFefp+XB60F6ZG9Pr8+t3HHry
UrCnsz2gJD5Nx5YtBMUex1ZWveV5EWrp4U5bvpx5J9ogzhAYOFl/tdNhF9cVicNI
cTqQzrVgwrsWgu1kTgzijzOk1ePUdfQmefWGtZKKJ+9YzDFQwZHUtukC3LxOeffC
VFJBn7oLh68xb7/OQZsAPj6SroqPUXDNIcfwSn9yaLhUWC1Zl2CQudVbsiXIQ7BV
kg7YwPViOVHeqwiSMjkx8oopz/ZL9fLLsJgkFrM76U/jxQ8AKxUj58HtBpA0LsdZ
3n0ec942zhGONBG17/ezc9bhILF6qLWH/L+EDX0DPSG90Nah5MhoHzNCcwREmQTf
IQLFgXi4/F6WqbIcupbWw86ESWUtSl4CR85DtoI+EJx7fEstFKXN+3rnHUdvfGHD
/b6SD9ZlNVPEA4CFCQR8RDXctLezRO4qUx3AMvLqoBwIWBewdGUJ78fKZTwzapJ9
MAsEJj8/GE9cCxcjdfanyjsfVbkuwR60OO6pdzJvO+R1DMctHkxq9iRrHd3dIdhU
5GGcvBY8EXUmMFmUt6Db9ifI/D7iCNn88aiS5J5nJMk6XZORfToOpehN9x3bXE+G
PyfZwRT2DWY6g8GjDRHKPhwlXmZWl/GxZ4xGFQjHq9fxbzgaqEfyCgablLyMazPA
Hv8P2U0iUxWbjhnvJiXnp4SJtKAWBlccatjMkGWDfP/bR+r5vaI+K6Da8WvYg0Ey
usCxCK+l7Tz/9PWDiELFogAvNBsXu63WeZRCpdmgD2gs+ZeMTiMsksZTX4gkeK3F
XyEOf5RjoY9o5D3D13wROsrhEAYOYBUhFPbsULqGYPEpRipJHTvsallxq05Bntd3
Om2smsRxEGJIVNkri78xFMLeqt+haW0LUlP7D4Tllm1D1hA8VDLuTri/GQ97gYDg
+4Oi2WtQGwSYwB6kKdsOOgLVDoZb17PFXMfdJImKY51ziIgh7q1CaBEB/4ndzwzz
suPhcoXPo7CD+LXzYrscTfAQVIGVKuP7M5fdQ2Igf6bZQamHcRf3op2MV1Sge0PK
PZHiyQH2HTAT7MDLJZpZTqKv53Y+2CrgD90EKLAyDN4fwIfg3prBJa5pDCw5xF2G
AqeX0oBU9piertyfiuGHVzW33gxTiFBteaEnAXnyLgyIWMLldXduR42AWVC9gRnJ
whutt0YCMpcQWGggHbOa3prSJ9fq8Z/K2KF3j96dFruaHLuYLPKluiBSu5T7ksez
q/waz/qBsFvDZ/zL6YSRxc1preOTNVIT3fcCt63FXazWBuoXUqEwm4cPNNxh069w
IazqgJzyxp5rGQzrLH5NeUq4UaNmFN1NNqePZEXjQg6of0zk16KxrAp6/EqEAt6L
DHRnao/3ucOM6M2pN0XLCreb9JO0zMCj85NPoOCeW89pfXsUA660K8XuQMRrmxpE
JC2yyPh8mRiQ4diy3qOKzZsnUjtRhpyr8c8Zsj+hCAxK9Q63VKOelpInf/kNfWiR
XRa3aHjigiQFEs+3cyNgsCRxOSGwGd2f9FxQ1Q6Q9VT/TApChOpPasxNbX5+aDP+
yMIqzXeQRQAm/cSPmS4Kipr40MUlvwvlSWi5ci8wzwVnP2w5HlYDVec8zbO5cBkZ
dwZyyPeHlyd7kK1KY2pUdJ70j+Xdf95PAVViy7/puusG8qbz21GPGyDCpfIfsGsl
Jgbu0N3OEw/FvIEivpIBss7TQMQo3i0DY/rUhNiQX+e64QXiPwWrXAobxGHkCK4o
SvEale0h6ZquvYlHBay9IYBJ206d9NuFvFE/LZd7rlBa3aJANI8SyrtCNsBwZehR
i13SvXxidhZP1yEXcHfQXuI0AddvAP31kxbiSDmFQDr2EVMc1EqJtsqObDghKGhi
DFgGsYPd1Npy0mztvKQJ5oF5jQuhKPlyJOOi/x0oCdLdjXI8A9Fdio+DnMVW1ZvC
ZEzXvjQdumyKPo2I1S2WXl//5HKD7f+YqzcwkS+SFe6sms/k7ifqI8T9tV15OhXy
yK9aGnM47xIN5UMTrkBHc0UMO3CXZZ00oyaNrwiCdErWy7+gtNqQ0+llz2ocPUDy
dRRTFU4z3l6qOIDPkqDkEHtxhS9VbQX1Y4amZqnfkC8XSKOisOHwh/+X3tCg7K8Y
VhNrDn15/AZew5QWD2W0sZs/npabHeyLxQ0UfqF78YdRen7p7iAAi/gBVar0zp0d
HpWWtlYyJfm8LD6dfzsDkDsprAZ4ipTe7r/H3/1BQgTiYfJculyCy1YYBLtkvmqa
uCdaPxxVC0mrzFelu1jaZZAoOH808FHKXLoG7y4SgU5NAd2OtR5oGbjRdnXTLClq
qq0gv6nu/MhewWHg/yqvWfybQ7j7CNO54qzN7QPCOb1a6t3iqE7cEHvg3kEllukm
LyWCNSR5SWzW/GRYvLHD/nDCw3SpQZ+ic20ZzpNF1bS4nWAb/RFaHioRzbQLY7Up
52gvLVG4Pw7cc+0EKgf5DPLgVg8DS80UNaXLbVscfSAigrwyAr2c6OhEl7mDqHLm
A0YGGBWoyaPg8SbU8fwAHg+6feBsuZsGAVFOa1MMyV4kq0HViewajE9es8qGuE1+
wo6xcxVsGHzjMBF+Tt+CnRRpzwWf2vDAA7/FaWiLe4v5YCzXNH0qpCWc1G/ZjDxD
yCYqhSTy473icEPFjItc5rOOuVT4feHVthgrN4aCOhciwPnTMahWBGZLAlfcmHFx
347W4D9+LLWvt90waR8ACwYf1W6Z7fkpXaAzq0t5rfGkKPzId4VnkAwtVvQM+mkV
MgFPEP0nARfaZff5rzb4tflo7DpvUo78H4r0etw1IEJP5apV1tUJjMw674LEhoBv
pIdYMKjwK3Nmn2vdDkLUlGWG7f2CQaL1zy+Hh5i4N24fPqI3MZZhVN8m96NRV5wp
ibXf1hTw/O4Ce/E+RXPjLTiS73sMfGQnAU4uSfoIcN1QHkM2zFR2XxAu1LKGXDtf
hJE9Ndsc2vv2KR3OM3mEYu/wIFEUitQQjbwbxkn9r7Py921lRqc7bLcTL14K8ZIF
XbiKQv9sB6m8CwbL5khGNaRBFw++W6YbTEBpaZWJka5maTJnhs2ndFASfnv3LVsG
bt7LKXz1Pj8/8eHS34b4XR7w1KK0GoMj8dExsdU9dWmuZA+IgUiQnYEOP4I99hpT
XQi3s00FKvpUAm15NcEAKDLIvvNLTJ34rVu0Kt4lnu9Nx0H5JBYcQ18FTa7DABTX
xp9UsBj+GJqdP7xrIXWy61wwXKLnF0AeQz1xTXQ2i5k3NrpBFNIBSSPsbKyJi9AI
NFc6B1J5z4GtbK9FM1UN8VYB8inXm7VfJtFZj8T2tW1jAob+2MLltLMP1H/Hsrxk
Afuh0ubSF4OqDcAjua2Zq4fncQJDb4mLWK2siEXZLVov/gK3hYGsPg4ZD6CRwhwn
A53MPWKfvBDkmPXdrlw9vouVOv1cjknAf0C9nhoLR6io3TVGrxXYOaqN0Gtw3+Xa
AvY3FumcijR3NqGDCec5RkjBZh9/9ReNTarXx7l6l4GWTbFdtd/hnf8IYlPWm4K1
NDaEm2c9va6xpcfq2lZHxpAygOREsPnERKZUbHQjsJqm0Js9wCvdexlkyMQYzcIw
upe8GIGr7Sg1TsVHXylUHET5eufJ6/Yt+4zl2n1rG+Tty9RpejQkrpckP6wcWFuW
Njwmwr+v9STyJ5x1hQ8YtiFT8h7bUk9mkDlsFhFxtxamx5Aid9bIAk+X6LUjANqD
Sa/ywPgTjmP/Dvm76NPJjq9BBOM7bBHjp0DLLAFYxZsw+HG43yGer1N/5gzvJ8PN
ruLGKwhz3s/MkwITbubv+PmbUs9bf5bia6GXPm+PFx10A26HEURCSbu/ZiyeQsvi
j8Y8POPZf418Au05Lov60uvwiw+FUGa/eElBsnzY/EAGLdm4QqZ+6whkr/SLYkM7
t7CrburBaCvh6fwF1NHdYycQMf/hAy6h+f2OgYN2J05YwSNUFctO3D+dfO3orAob
9fXRKaTLa1kon8S+jsd91sTft63N7biFMqEGipafTFMeSd4pVczWwkEWmml9/9X8
9ue5+3gnzbVr11X/1A5Cl126AYAxB7i1gUgT7TFKon1CBno7HlZD+NkT1aysD+Va
4sCYNlNumgk6jK68mr69OqaMU2nPxDOtSnOX20U5W4zweK/YdkJNfv/AEcmlhQI3
bd8DdQTiJ3Nde2ycXfnbWY7J5rzimk4gVvtIWQpeJFcNhfxeqeN/PNm8P/2/O33J
nO9gAmDOxYeAlC6uvOuRZWY1PuSS/89Hxr2mEIvMD+st6s53j7HMpzSSxKSgqQ8D
hHNS0xtM9fH0qq2aYl0rvaUa390PfGZQ3mHho3aTcWo2kWCLW8lLAqgzrug6MGYo
5cIIxXk3jnVyoU3Xcy4UJjphqn17vMh+pZ6bylhka11g92ySpeG9VPRlzVV2/EoL
FqC+iUX/LAYSggaj8ZB8mZHKLU9Qmm1/D2pScaL7N7+CrW8zSDBfYnr8z0HTDc6u
gnWZkgyUBWXUwofwyf/VcqTpAAm3BYxU3xVBWLqmRq/D4MKuKiaORqTb1ktAUYg7
TX0AS1dmeeFVQZNlyyuFO9QEy4PF1TWK3x4pIu0QBJpO7Zu970xYhsDWX/KWY/2b
DKhr3pJ3gPfSBXc+0J+Q+6+olzgECiZr/MvdwprakYySyw9SNAuW39eI6hRBpN5Z
Hst/fkd/xn25zjzfbjFV4CwZVAgurbQbeo6qbTGa50yVQUCnJy/Sow91QqigrGzv
yHbh0Mq4DeSKaKJW+GJ+y6X+1TSxK73QgpMAzZV0g8JHlNQtuPU1UZAeHSuLgWAg
DlXoXrqQ0grDWkGzWQ/GmqZqikTTdFVeSKEgfoC++p9i9GHB6lUTP+FeGnPfEJ+d
j8S1lP5ozfT/9dTo14DdE3Ul2yyy1aTKwcw/jNYVnTm3iHiFKgK8tNLrN0qqFkCz
7CsxGAlCARnmyLwHrZwQ1JoAPZpgcEZm8NKYQqCuDOm27E5lbwKCwwa/bPRdWnj3
Uud5j31MFvNUDGsclrua5b3uOe0tMvvky9dkJ6yHj61me9ayvIQ9Q1VrA8MAJWXJ
uHZUcUqk5e+8YbSMzyzr5GZ9kMBkQznhEb+Tgj9l8fQRiaUtaiFle4Af3D6W2Jlo
eVEl8RA54FV6rBIhVZHk6Q85I/P1Ax4uU2YQc3N3lNa+dFHGiWgwauZvxmT08zdv
Tg91vB9+nvV/UbPpZukrDP5/gzyKERuUXWkn0IyvEp9S32kAJ8fOLQKkJrrZxn+X
3gUkcQ6si+So9dGa8bHuL5QX7p9bPo74S36QlNxdwOK0jNERizALX9PP0jQGwqcC
X0fCWfVSp0C6aLevAR0lYTbFzIp5Oq1qNUHjGmbgFKNYc6taOgHfn0DUcC1d2EIY
scvQSTiBaY5uXmsmCmxm+Q5p/aHaPsg58aykkkG49AAAeUz1RLYMrgJhHfzmdqw3
m53KcaKwTwq42mDmwCZeaggEjmRIWW3Dritt5v/KK6A6erezCoz79mwnFE7gnUMB
HTBkahAkFDQ1k39yOGo0UGGpf1I/nYUcvOOuT1kMlTKlZx47zamqfIN7mqxvoiSr
2gWFpSoi4N+vl/8v1OCEVprORG1iTb7KT5povdjf5x9iAP2NdzGcT1TVL0bcMzu9
2ZadysT5csZkaMij2ErNypaQfxLQIhjRd1Z4+w1huI5YMNLUV1UF3IVLD1TfjnFc
xur6SxDu7uUYLKvgUEzu7mvSA7tZGdoF/NTVj+boBYKWT/W5iLgBzFTGLHjBeuIb
T874+ch4XeaGJXKQlutI6o7kaVbznm6aE+6n0F1J3Yyc+hUDbG5yDIZKipGBrLAv
N/Da7vo2VpPAQEXe83OAkh4Df/b0YsoSDxRfSRq1yXuEkM6l7BUGGnd07pDQePb6
MtLEdsL9WhV/e7LAZm6mR3P4RnIpwMhSWoeq3ucXubO5uRm4CniMU997JF8s9o52
HFGuR7kphHsAKQvnvgRE/5H4nzWbDeaTpeNgCCP/ppo/1opkrII/B8IsUv+VXI+u
cnRSkJi4UZCNhhK7KNukmfhc+G3aXiE89uWTNxLGeWL+tuIoegUbtuKzFJwCywka
8Wq09LpPhU1pqrexlJbvIA==
`protect END_PROTECTED
