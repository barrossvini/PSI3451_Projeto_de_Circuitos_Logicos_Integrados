`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1wNXkGLvIaiNZXTP67x3heIJMIFSbbeZ1Fs0EP0cHlG6jCTadmhGmMGzwAUIsZoF
LWUsGw4ko+1EKuzihNLrOkGW5MdatR1d55/UcyhF5jaYB2LjBh5GbwmcWnK1RMrG
1dU22Fv+f7wv95zVzzCbRjRP2SdxgyNtqoMiMNkBZKqW3zlAj56Pt9ZAaJ1v75mR
d/ARtsMkBNAwAnR+tuiDB0DQCWaTmlluF/6DwxBiyfTJmvX9SkZ/iVSC92QjbJ7x
BXp6xRzbbGCLfj7b6ZcYxA9lMj+rZoUWAVzrmII+9LrmrHZhm78ONqaWejLoGhgI
K2bWmUdj+rMv/JCEYpvRe8b+kaHOIWisu75dv4xbNUpdwMLewOeeHNsOGwPTataD
q4UjFndmgJHZJzAJr6+uaMaQ41VsazWthvq2otd1AVOWpYnoKJ7UsrnkzWEhOjAo
t1Yt5XYncSiem2hSKs1E/W8lXSc2L7HnN6Qj8cVAjT/OQg7sOz1piD7wo04osXJx
DaXLpDA6fC23NoZgQK66sGwGZ0fNmPLGOkzKV5qKarPnvSLktSD9V6u9QPyXmNvD
3aaUcHlyL/gn/bsCIJBco8CovSWCSjFFk8F1RjQsqWhXqySgASYidvorE8agfLhE
0eU57a7pG2qH+kg01595ff7dZaxy3ZO66GBLA9cDt1a/hF64FIoT+gJbQ6goKyYW
NBHko8HaZxw5VCA21uFMcw/fkPKo8cNfWQO7AJX2NbWZM7s6HQSgCPWjFX4h+3pB
qTAn44WbBVa8D6CASUWdHtityclpwYYaAixSRtdAYmpBa+LidxMi4nFoZ0Fe9RDd
3YpgMvLxo8pols6YRyKCEwAYt48BbUrneF37pl/lVrtf+cvD/O46BZjIAgI7MOih
IDLR8S13x4ro2lVKz8lG4Yk5R6Gxk1ULTXM5RrD4bmmRZ9iPeNA+0haSaWUVpU7/
tu5WjGln08SagFLKEdnShBBNzRkeLONJZPcdk7ZDpq0xidqlzGOgh7jVe8+bt8AJ
Mma73gWDcb/xUmL6HYlSoMyY6sDj99UV805l4Ltm7WCsXzRFgo4Yz5DkVRHcuzs8
76MnXYveciXvnJUrr5g727TZHkXXt7WQUhwy0d1E9QeoRZqtyvbT6J/mEDf2T9Oo
/N07N6jYUOPSswkC3OiS53PAHa/gPiGvZOf6xJ2GVdsuAnjrgy3VvGk7PrbYpMC4
744XgiOn4G146vHofJayp/rVMdYbRJ+oapeyt5lVBZmmsVsh1FVZBdpp0zUAJCt/
usT+f9yfDH+E5tAWsRdKU2hi2WCqT+nuUTRiKvy+i7/FVNRr+ehQOremNa7vLRMz
70R07QnE5DzPdZ27onC5EYiDplH/eKC/BtHUpOqKo8sc2Pi+vfuNTBTZIlduFYA9
XKwNZqyqHzhUD9UVJoRtG10CNw9jSLZQmhM/pxM2ZkVmXuPoeIP55Ylkdk/r7nhR
89kjWgAejSe5SuQAZsYyomMy1e6ygTkqOKZdvFEgWGNHq/7ECLRgt6UlT1cc8R65
iDGLt6Iq113ykFwJeJEtQmP/COOBHbqIJMQgisa7aZQADC/Jv0vt69vRuO+z+kpD
RueY05lwD1tAd0dA393QBD5DuRLLkF0DaiBbI4KTDJnPqiT+qU5ekLKMma9CspnI
owmEh+OGBNKyxYt0GkjeNc5g0UnEQzTgcAhQ/l6JtFcYaRKKyfvqJtOYLdrCM7SG
nMZCFk0+wWBolyo+6w5n2h7k3UKGA0FA1skSpeQHmFnUqY2xk5Gl1Q92O6T+0rkS
l1wKXJPmCA4CoRJPmfMW+8plm/3xyOhmiEfAIY+ffhwgOxdqBB8dPB6XC7Z/xV70
jKRKEvELUEiRr61AMqZAJTx6XrYv6QqEpWSd+Ux/BoZvl+a9LKv0yzHQuvWJorCC
To2EiBpU6ExhxOeLolZ+ZBtavCi47937g68i4rMkXOqmhqaOAi9Ou+UG1W3Vul0g
GCgaQ42b9KqbQ01gVZebCNQnkUZ9ThA4fUWMyLn1EflPg87wOhzsEiUe6YcS6LD7
S6qVgqHcnezUfGqPRDF6v9cSdXOzwhAUZ2P5z/9nMhcDc8zeshbodU4+DGFMvAB8
ZYiV90kxNjfkjz7vTT9a6fI1hTzMgLZ/QNGSMwl44hVntvF+xgYXjfILVEIkskHR
i0vayBGxdLepB0+Fig8tVouvEeJe74Ho86tAhVks3NK2sEzQqanyBQdbca0sFZra
9ZhnL3LtvResRsaIX/4W14RtcilR06HJI0f+lst8kND5m5P2DFe6jYNzn6Wl0aow
ACMem8b1J7Tyx0qs68pB6jIW2fbi2tYbGkvup7FhI6l/ls8yNZFXrrpiT2lOgAcM
xGsgDJLPUVKCzlZcVTH2G1zbKkngpMetEXkzX33xqagMePkI8xCRyVhHi1HaCPzY
Vvt/bFuPoz30dtJaJTPdB3im2liNW05h52HyH+RSgVltaRIS0ui2D6QofGpm+i3v
DWqEj2yMmYSaqouVOq+5G1h2xfKLfIfzXaiGvrIshpr8SabUz/U7eZfkJI4sIj1I
h4au8eDeSjnRL36py8cB14rrkiC3I5e0+czr2wWH2Iv33J8Np7NjylVf3PH9KaT4
Iqwt0e2J8jSSYsnobJMwyRJcyglrtIw/tYAQ3/r5W6g9yXQ7w0GJJf/NQKbl+Nse
4rs4NxpTAVIeVuNRYdLkqDJC2K5isggBezzhxEdDKIATzdfeaUo5TbyWjTMiMfnR
V8Qr7HolyogEba9ptqzDYnT75yk5Gb5zkXcj+ES8I/Lddx/9GqvN6aWeAFMiW/9j
jbL1efsF05wL9WlIJfSuNH+Ir/4MTy+pt6vt0WnwyrQrv/ElfU1enUMKv2Pa0L40
OqsDxbs6gVe1vL40Wk7vbK0YHX5Elud9ra0R8HZ3MCM1Q94mDyEn9Rjyv4pj4wHj
YhuafNBkQJfNQg3S+5MG21iCmTwxQbBRv56p+bI/+EuLpPTR9nE2Nxy/y+Og6UDv
QiolhRiQiEGf167/IzgYBVCCwfo/m+xea+xM36ZdLikrL6px/b1CkdIrPpdWcJC2
ogBlCvoRTRszqPFoT11TOrznOMnoQwN4twENymWKvIiol4o/gYvhNl6IEQuIQM15
IthFmjZYl1TpMwZyWLbqhm4Q68Lo/jfnTDS15t/8EH7r74K4B57iQMxo4L2Hqoiw
GkO4I4jQdI5xFMpt1YVaE6Hz5oK1ZCA7ulsuTuol5vC+xanydUJal06d4+IXJ0cX
/L/ScIM8DLuDrbHiCykq9UvypPowd2ABgn9zfJsJXLqIW2avmnSHbif3+MN2Zmx1
6J6N/UWCk6ScaIr7XdWu7dB6A5dybG4OjSs0tM4xiIHFc+GmjZ+Uvkm1H1+0oyaF
pqvyQu/vnS9Yca7dxg6pQgY0WpzazMZbAX1LeIyb2Nqvg0GSqmxcAwzFWQojZtaR
vI3xaWUi+wbE+hMZpE1eBiS2dPEOGfFUvC8XDAQBnasDRfWL6hyAiE3ulBaRcRAG
df1CTBRuLbslWX8HASwBUuzEtK5yxPfkhhJlDAmUIQHCNs78rX13FGFlFykwzUqc
3Czuj6JaThtbPAbmGXLuvFttM6eLOjouHUE/OylsuBJ1WtZS4Qk7lJ0YfpFmcjdk
dKVwqtkzr1pBui0gRroOSFTui2TIq3s7KAlvUMB1WMPKkpPk+nLhE56zylHwZPr6
RC6WlvD0RK/mZi91wKRWDEE8PxHRViiOzaqezO3DRSbVi0VmhFQz8wu4C0LBrifV
qBHiEnV7G+n646OeryOrvSqEvSK3m3Exr8iMbEUIMKBvQz/gOnqBFcmrZvlDp4j0
5Y8PExJb2sCVz//USBMpYLBCSpK8Xqcl6QBeUplb8U8lBR62CuKA9G5ESVBhCv23
WQdaji2d/pYStEcNucOuhi625IbZ1QKZRzeCelenrNT1WlND/IJHW8+ZzIHdDUqv
jWtG/QJ1VeBjggGaQL65AKsDqWZJfzgMQSJ6+FW+aBtQTfTD+ui99oMt/vklMkyd
S8ll+iHOPMmiQlOkb1Av3NBZyyejCudxfMV+JyuYGGJZBnKbee7sk/cdN3VLFlme
hRlP187AfOmeT0OaRDyNe7PI+KdEcKTDwItduUbE2jLrR1efsLX7gbm1rTUtH+Mp
A92QoGeJFVyvR91qT0IF3hNDu5ytYfvtUURoxRJajsb15ye3ISskb1u2kvgUXsJZ
2WFN3kHRymHBerOAQZzgsl78ExUblFM83LPd/k/yqlWfDZPMOCJmOWLZ/9QRoVH+
RhUwStzw4bikhStEs0dqgoyt6smU75+x0ugehAzTdXugkFHKhbLhso3Z1GM9VA0Q
8YRIVLiO+ZMzIGmmHX6poUetemi3tgabUTdraKHQL5m6OdWpWD0/XTNLD2l0l8PB
YGqD6LasZevYa/BHiUo6D7DaOxC27oKyUSW0pJ9IK6BuUoe2f1z6a8YxBGhS8y3O
o+RzuJn2+uBnHOpXgTC59KmY2Td5nvsIA4ST1/9qHIl3CmwZLoz8SCOt83aKbbmP
BKCFNTbPIaZiDZ3QRSZvf024Ii44UQyjq/LNhuJigtyg44yi+9RMg2CgpsnH0R1+
sv/wHVCVlTnXM71ROpBlwrnoqgHVgTg3IwSFw5A7kI75vpTB8QtQ1Nzk2dli701H
k9pwuWGTKKbelA64PYcIMrebnd/gBDjBpRc/tRXQBzckDsD7C+D1y+tmWnPI4x35
m6roON5tdn+aAfwPHrxrW0JGtv9Q5QVxO0FB2wiJeT46XMN9CKnlDoJWvsFYB4sa
WMkaRDlCHWc0z90u7mTTsLcgBlk15FkztGmibzfUtskqg4CW51MTRppR4J7n7e7K
WnDRDeQ+glGnKnTQc0Vtm4I6lj7gViLhiolJBFV0gTAZRg48QOehLhi+AjfQ5myu
sNBrI/8m6TAEjV90cN4QRHGoO1dhCTxIc+gtMYaOFq/eRmHReqznZE37NUiMLCJ8
TiZxki5uDuQ/xhFd6P5wJ5mcgxHOGKwqMtnpExDmJrRW221BG9lOpvmOFttprpUH
ZICFCkwl5OdHT6ThukhTQ8elqFcODyDCCsztAi5LqYSfc7W0SJVbhF4jjvorqjTf
W0/rVSNaSQ1bTlnVbSSco5aEKTnRlA0evcXt9sW9Awc+hua6P3RU2B6ZJrZZ+nIU
uODW//G2mJStXrevsZ8zbqGcat9ceAoyk/NbtwHCCG4LapeZMBV0A/cRcb4poD90
5guGEpJ0KasG4t5UkfANfTT5dAVWKsNvUhJnFtUh4R2CJa9YIw/zVET8mSQZJ9Ij
va1+xFrTxqFEU5S2Q/JvnL1/HTfUxVSKXnO+aeTafI+F6L2nIOWVXcoGzY5eYz+k
m2RehM4T1vE5KxuKbGTCY9fgHUPqu5hDZqH1m4Bqh0AKju/7UjneQvPLRU8zhdfT
bXhZUddCRn5QeuBbtTB0m8CZr47pTOvHtPi+EHL0gNwkaPAsbsKVB1SfGmOvqLji
nw7gJyZnxh3D+fD/JJjS71XZIAWo4nPiw3DNu+CqaciGfr21hsiWktF1oqFC8m/K
X1SSBS8SJwoFJvUyb5XKWaCFhKNfqUro+fP4ttN9csjwajFzlog7UsSR/dbXRu04
Th0689z67jrSr2x8rdlqYYFW90KjR5N78C520EVd9TAFtUWoDQ0wSstn0ItE1wHS
1ToAKRiOg6aKy2HKAaEFySWUNm/mn8TbsUbU8Hl9dUrVKlBq7++FpqGlYZ6kp81D
P7HC2eexdVB3Jjq41zC6O64YrH6+Tf80xfNBD7AhyggKjivnBuRDsM4ric7ZbTbH
951T1cnpcUD6lmikXfQRSB4GJT0vpRn0sKxikxuWVYF0xheykgMJIyY8QQUdu8zr
IaSPATUQqEDMefrohN3a2YvSKcZm9wooCl6Sd+7JoN8WGMIfjmGVqepYIwlCNTQ2
8SQj3IxFUNDtZ8jI7TrcUc7G8yes5mr7icjS2wHgwndENJHa/wggMF24y6o/delm
JhcBlhDomG9uP0ZlpTouB8B8G5HeuNjPHibdwGf3G5/ej4RwBK6qJ9qa+ME2qcmS
ZtW44ZjrW373UIJknPWqBCSVvQQ1zqKz68dWAGBEUIWcH216yUAxnc3OPfVehd+w
DuIbEpZ0SqNux0xc9bhhTrebReAhBLN9qdEB1rTmusZ2t5qgWLcxmeXU5VgpKdb5
95MTdbsvfb1dqaOSE5enMch836+18OdUSOKT+vvQSDPB5De6PqkOPI3owe8AeYHJ
RnH3ZZaHNcvXuAfjliA55HYSqJ1lZLwkiyQolribd5aoF7u91+04IhsMZOELdwRh
6+4VoXf5Eg+j87U+O0+WN2YwNM9Ibu4TQIXa0zjiLZMSJgaaNUriLR4YqQPvVxHX
C7ppqCoZY3c60vqKaIt/v6RwBq4dwmxRZMjYj4n7aENbTP+sFNemSVKshdu8fkpA
dDrYOICCfpTq0nVhwt6k3Uane9B20pE6pRwYMWamf3kUq3FYMsdOtJbT74DkPHFL
EbPMOtKUsWwZGLA5B/WfyqlLveNgXAEe8bYyrR9d6W1I1rwDv5/fy6uj2OVvyRmi
LgSmtdriWgvwgpSreHlBLTdRacrIuqikMSEYM+SJIt9YIa+G8ArShxVXUKDUCXHn
OhtKH7GSUwttCvU0Ko5c0QB7DQ4G9x4W7rJvW2v6KonfVeV3BdRn7B5E6KCtAMII
2WWgik3mdTX3YzFcP1viPE2yekjfAZMBS9XWuCO4sjxLYIYau/lqS+zPcN9t1HQP
wnJ5hP4pIb2a5LfJoxIo6+LVUX5/M/ottkmq2kgM+TOn8kdR26IXYCfe8LdsDJyL
wVZb8IhqT/31Sr5mJ/nFsycjDzBs+UPuOnxRbW7mT9LguG5uA2kXqaGZ4hv2cvz/
VdYn1Pzq0Raq+QOD281xuR0J68DwEHH1XqxHonHRqS4+wDc/VCtdRqhannB5TaEk
xBTg+unAlg0ftGhkkVGtWZT+SET2jKDHPIWTacud9wtl6rt19trF3skJfmZqsBwh
q47fJ55wORgFqcsW5MsQpW1GIQjtUo3qwcj3F/+skqCGUVqIvhY9S7KMxDvdleWg
LcCOF56ICXyhrHcLsF9knB+mg4lkWWWJLkpByk2XG1HHkbD6d7OGlcwY3eIHZkXW
G0LBuDx1M7lbgS1u+TUqx06fFQtStdsTTtsitFVZaVF1lf4O1LfU2TX3OF28naS7
z9eXswAEughNQMjeJkBZez4WHdT7LnWGA+/y3JQPBXQOR8XvG3JC5Y/430dtM2dl
S65uiMLkNDC03uEPMJ8t/2xZvm+mjMF+GrchyCNaKg+r5+jrg1IcWlCiz2rGsMkD
XfMMSIFPf3oh6MwVm2SBrvjKRvrexHKhGwj4QFGAejbwLFziWLFZibaaooJmqi+7
C0HQ9bnDRf871Qwrh8enioJ2DBSvlPKE2qRDqf8deqEZun9rbxpotgRSTRxYpUiB
MMEoNmgDn/JKedx2dMJI2vUHUe48DdZphJOrp0tGd3JNEnHZ+UY8bKllZxxQlGxy
X7dp9ItOlHgmDsx7+BOYhQ+s/o+XtRpmKHA8Hi+13ti4hyu5mB4m4Mrj2Et3EQrJ
2P6P/ntZ8ZJRX1H7bOCrOkAxNQzxcYL/1nHWYyy2jkoWAm8jPTnzgW/6P/X0TcrK
yYLtTNAX3tB7JnctcgH6fSaqmbbbWPFMqIMe9ea90X23ePF/r+/AZNjyRV7e539J
ZFAj6fm8GbCmPxDrslg7oEdzQGInA+DAfyybYcdgWN+eH/JGNIpL/Eqy6mdzXvch
bgFzytPLAQe4iM14QoZjS8nbAMyv9uv+gmjEdvaE7TbmAd8vkuzy3svNvDrDVLTh
B6OBvdYMLf0Z5+n33dY/p0xR1wzrK2gN8Yu4x1wx8y48alqXmSGZupV8D4At7/Xv
T70BB8g5bF11SZUsYlwHzTzSdAqzUZMmvPJi84a8+OKr36CFb7MX04b1hzzfZuC6
50i+Os8InaHXZmIhd7sg5a3mhYMl6lecw1Se2ldOgucfQW5LkBzOqKIqi02Pr2Ly
p69Nj1gkWH8qr6EXspEOgDwFwJ7mOD4YtZLFP29ovJSL6VKZTWyL1YmoOKfATwBO
qJqz8lbmeXpjfbPw4YXOYpSRkF76xaW/oZwIgTElmoO3r0TPMIGMUNO23UiP/f3X
n9167Xyvysag44RkPasaXpg1JhaWPLM5zaa8mYqsaRpX+h2eFoWAwZu0ouxt+Thg
vQDO11pUvqdZoT2vMtCyLBh60AD4s955OD7sB9J1nOl/CWrpusEV4RRWfDsC0q2s
QjrDTgaeUY/AIMI1Pzv8AjsCuuRDLNDp2oCkwAeRYh0QuSAoWTMkPFEaN2rHholp
laemFGab6VwFkHTWGRL3PWSC6iiwr+pPZApwZal+XHq4Tb64pcod/s6TnyAPCUPj
uBsY6b1jPIfQLPN5mqTuwV9mWazO5vbBeQDMiK5RlBoKxTS9xNSJlvAgsBpejjWb
EW5tDE+Qb4QHubDT15w5KMPDvlruEiaCfyp4KGTSKv3lMYI2ZK8w++80VotxaKgR
S9ebyPEae4jrdjnRoJgdQat7bBNFDmDVuOv7/Bqwkf+pqsACgmHzPgkTVaoLsjJo
Gu7jTzVuuVWw7No1DlmjUZsgBQayktrgHVSBfDnO4KbpO+2e0rNNZGBR0uNf270R
7N1FtodyabNdRaVzWTo9JNcwAg1PQY/YV7ycq4pJAtYXaZneVS6U6HRH+GAWb5QN
Trco3VnwpnNN+6San/n8UIMWj8JnFlBAE0wGU7F4J2VFQRFWtXitwXkDK/cY1Fps
qVFvi1Q0JiMjzA2vYlJyYzxUz8lx3Q1r415irJvnH8hcxIUFXkrgLeljsVt1mJYx
lqqlRE47B5V71+gqEjdenBq1e0NSSRopzDqT8F7ac067RGYjYksSPAvGEU+TuSfw
euLfsVFtlFUWYZmrAbICkoJo6qjYiLJ0lnw3cj0MM5nMn9oXn5vqx8pzY9b+RsVq
ZRMIlGUkgcSNd3iGlLF6gxm/GyOjbRBWOZQ7tmEHll98rje8LypPjvgFYOfXZhVi
hlgw7Fd4XniXR4tHeqg3AGt4nOIizTpFgAE9H3RDYmOz1tzAnPqqU3fRZBNKv2sT
FR342DOeYOE7Sr3ZyMsZBj+ghC+icArsrlxoGaQHKbh4faAUtpTZa4rBmlJzeI5G
RzIEGfJXcyRbXbhKQniKu1Bns3yMgpMoay3Z6wQA1EDRrjIWqsNUX6KXumXpkeom
F7fYrnHEjyEOticOoTa3zk8FctjgI21CjaDs4CdF55JyHt3dn+JcQWja3fMitb2A
4CCFKQLu56NC4brkz0UrGVYYxyprgztp/do6yCLnnhx/tRoCYia2jQ0Dor0pW8t4
bM4EeLlp7LAJaNC0hL0OqOJ5ic21emv/+EWazaqjeCkEa7m2eNledfTY41tGjW1y
fYNx7aQUImwWNo/CSus74m+Z4Da1xZ6ZivjrbrNVdV7eB1IEuLxDjYUPdi08ISAA
6rftreeVRWp29Ye9qKG2G7DwKiBhnMxTsHUFXLDvoy+BKhjFRIuaZkAVX/q8KBRh
QtMh7e/JyH6mFYntfQKaw3KlzUz9Jpx1n2HniAcdQbtY2Dzl5tFGZeBqzKpIJJ82
2kn0piajEHwjuLBTgSZ6JXIM3f/9jz+7Vj/9FqCLJ/okcRlXbKN4Lzm2HK6k5/al
w8ylmR77RRasJOO6j0fDnjdEMVGQP0nHEN0YY/FZU1nETnQ+2AH7f3fi3shMkrzL
zIsgkjV+4qYuKl0ZuRmpfwijH/3bFdMIx+0Q3ec3L20+4kKG9zhxywlf+QaZZ/Yw
6QAMEka5d0+nCMd0AjlKPgX4QhuiNZR765DTFhJ3v8gFspAEokdqEfyzp+qcrILD
2CBCmO7nfhkY/kNBzLxGSnkCu0U0ZHH5+1IMgsdMmvyUToeLOh+gX9opkhOD+iH5
1dOKDICTqule8oKmiiT8Jy6qG0sO34z6UcZ6agYgipMkLNS06NNphU0/3DMZ7ABf
L+OrAnGzTI0OiBfB2wsg9Frh/fuS+T+ZALUTzSkKjeDHgsfe/QID5nrAOBfRzFGz
0YYV7Gn2UJpoOwPpyShEAJ/ycw047oTMaW5QCaDiItJm84QLvPa2Xx4I5kFqvNAE
QrNBqxgiwx9bNMOngMR7AL4BS7gmJPnoxNjIPUW3pMzQo+Df376ogaLJHze4Ucx+
uI16shfLRnhj7EUAbF9OBbAP9lbw0NGtQBBonSEig01Ea2t7Ov3bSsHLvLr6J3Ng
ewoWk1W+iEO1mh+fs/qqxEBKZ12eBJWwNlVhFN90AzTJt1l+aOo18a0YTSVWfG9D
cERz3zh4eZtOCVrgU9hdUhywoVooqtbgWEnFJ1Z9UgsfqvYERSmFyNaNlEa3zWt0
RpBzV8OJZZqxyexPrhtJ/TPdi0lWEu2Zzuv1og3AV7FnQRyyFT4oNiy+9h1Z4xMQ
qFklMvE0bvz/ub62TulqSgz2GEQNzS+qJfa5aafA6yedNlA6pYAFdsmcLFgAx1Ft
kAVA1VbAjOF9wo7RjwoPtYlUY+pOwhdf0rSn+tkjL7vCBC1W41mIeT5E4BCDEYpb
ksr0tChOfxtN53mHbdSJC/Sl/+T1mpmELOb7sOqKAqg99X1B6pBA9i1cyBUuUMn+
tTDjwNbsKmnxw2xeM7+uXgyssGtGlNms7P//p6bjHA4G/+Hz5ewD0MEl4vplGaY9
GlnveyF04ALylBIjTDZfQcbhNFNaZZOp1DCprBa3H7GcPyWZRatzB7pbbf4wCduO
zrTeUhp+26RqbUqJ372zc354WKfUkaJQbHvZrp11nv1pIbTBYP1RpRBANh2QMd5f
jdAyYDNCqpQ5PSHPYlHxuP9kbVNGk+6aAvuoONQVylAnqrofL1qg0sTXn4x9ZXeH
op2XMbGTTrPTPlJp8RkRajACut5MWkjIc3nVPVgCRCq00koexmfmS3A8jdhIYzXc
XjGt9i886CUgqa0+pt/fxUe3FL6c3YPL7p6TzpmHWXGQ7mQv3G1jf2oM1PcdwCoX
Uayva2zsBJylma4AVZESqW6jEQyUTZU7A6NXWGTOPJXwjNtylcNaEapoj/+osNXT
HTx1ipUX1qNldClHKIkAlap1sfty1O6Gl3pO13BI8rknCjOeCsBMQ2PCqW7q5xS0
ap+5QH4H116Zw6sR4trgfO2zqHqRsYnT6akXafbC9CNEeDjI60JIWB6xn4kjXcMU
XA0OBB0K1ZNaL/xltbgMDyTzCy1aV03ukNAgBih9KGREi+rw3u0UCMEoK3sZm04t
ziX7903ab3X6KKIsNVn1Dql4gokK4DMd0jX+imt8RJWwTyXBc5FuacwYcn00cpdQ
kyyyrubD8VqV3K+2Sfa//0kUeiJH6f7qREtxKYxWxT2tF9l2DpaV/2JBwIrXudNA
ZWUjYxZPayMTWHmHVr49hKtZYpXsPrm5rc5k5ZO9c0oUpDUBkYz3QtacYEzyQ9/L
BE+KhymtGOGYbhu8+QB5Kn9z/4VKux6aYD3VAKc820678rIhDtmBXrTk9zPZAYJ3
+yVT0poibVGsbJj5Wv8mNoKyVyb9i0Qq5Ltihqw8C9ylDo5c4Bp4npbDbPq4MhYC
+WJ4h9Ban5KyfJjf5FSe7tKxkwvp8ko2SYo9UiTDObaNW8B/MS7Rs/f0VlbMglbk
UBxAx+RXRa60ZVNgVUKYB5Al1IRMqqGgedocKmibdUiE+3mmri68eYFeSesDoKgG
JJTmRKOV8df9ygSZpChuT1smdwtgAAPFGPAEJjgheYcWg+wcYE+iFV3sCVvd0szg
P6YZkyFhc8Vp8W9aPn4zTPuS1IeZm7kkN55JYp1WTU3OB69IlTXflFZt+PpNL6Oe
S2YQ+6V3fGRp+nduyERaRJMSKsqYNsuTLOk1ElDYxYVns/W85xX4Mk0iNSAraARN
dICAg/x+9ZEOg/fg86bPC1ZiAA21uYEZyFTl0CFYipAYunGrES/981xKnTA+1yOS
uOGE1Bi4cFGsAA+DL/gPn15p3Cvzeq5HOmKl1wf13PZiYyx+g7i4sjTZFgC1YFjK
8h208SuoZQ0fXrs9tKaVHHfI63UaQrbW+AYxZwCIhPMCAyfS3gznIrf8nx3PYLYY
Z6/bzju2HaGyE/D7dv1vIXYSNM8B2TFIzCOzVc293Q0Zl2JVAO8t+BhFMgHcdHyq
1TLyJpGqTHxN8DQ3c1Cnpk/WLD3RtvVvIDRi+4bS76woXpio/kASk8oLGVuQMlt0
A9CBZ2jdkia3ZWWQ1dOtkXM/zam+Thvk48jeX2lSKLeHUxT69necZhN6kqCEkv8w
+/9UpAO+J1CK9XvFBnR7yGmQ7bsg3xcq/j2a0L/JvqLVs2pnUfL76lZjUPQwjh4L
8WYk/HZBQb28zgXpay7Bgysj8RQNy1lgX/iYCzcVpHAQpITkDT2inIiba/iEBXMc
k5xU9nA7HsLiXCpqC60jMNgF+iBTH+UOY15dJaGk3oN+8mv7Tk5X+KubK6v94Q+h
zbvTULyqPvF+fSYcAjgYoYyK1OU+oAjLJEOPQ4nHZq8C0YgH1AJNyTdicsgQYJdB
riVIMAvXahdaKhZJprvgsSkyp7sYd/p/2dwfvrIBa4AEcQzQJEVNmAHspVm2u9bm
8BMza7ZHltqfKBxQSThjz9C6XgfB0o5uxdSSJVTiaeYF7k5BLa+KZ75ondGtzGcz
s6EXExFSkkdJZxO29I0cVyVNlq390ZDIupis4WBCKza98k+pMGolCKCE2s4MfiFN
UTdugYHZVK1tt4z4BYzReYwMfZNH0KFhFAyCohcTYJ62uKd693aOb6bArdaUv8D/
zZEcvyWWSkZb0vqwpJVnPEnPLOS3T0V3SRcVBqDGim+RsF7Rabope45tkAuTlA31
2A70qBWojPIPK3fCldmTyQz80w4wdXWPB60CyNZFSx7Is9m7RvAxasNspTcVEwdJ
aRhfLyp+TTz7M0a1TiSDhln54isQSJx6En4Fzh9kypiqD9OsJ8aXNipJdQu/wvZU
2CoEFKqMRbdY40vbWuXsMpMXd4ySRvZZk9Ffd4e7AmfuZEtl/sxRhvK0EYCFuva2
SN3+lK/7/S78HBAp+3vtYCeq/lKJ1fyGz0HHPmtByNSiv8viVFJ1fXij5+2MopJr
+B94DtPqc1OXuSJdKd8BCN4M/srVmJsZ+7lWxaqGdWm38ELAodV/QKLqHPcNosOh
m7jhISQYWmFU1u+DOTJY9LKMGGuwhMKX96SCFWzN304vv3McERCdsNwV82EQL99P
164XZqwALlLsIWJS9VEyOLpqZkoJ/JPACqqyHiuGl9DXFRqhc8wvbBUB0pLbp76p
veKdLIf2pJW5SV/VG0Jn2/zrQ83ZsIhx/4fyfxfboYPWqJURraYGGKArh9dVsTPd
xpbbMcnunqXWHWM7CBkkwfrVnkmvSUKnTboZ6be/sr1EEQiNNf8GouM4x8+IdQFg
IP2ywkNhdUJJQrHE87LFHZez4m1LjBehbmFFZKpVL3plla0vUSg8ojjtxPX/wPBm
dlnhVBDSocICV3WhZSiBAHRBo0PuPS2sDiwXPaYxv2QLNrNbX3AFlpB2RdFnaCG9
s44yT9/o/5ProbDnWZU/Psj872YqUsRw3GeKQSeRkztN37SK+XqcrSxopdOIBeMh
6uRgDxn0EWBcuBlvDWLUZr3lYbNWWO7zK8oZhCmUyRBpQ2uOacaHpUflxlugNl6F
taxQ/LH8NdCnST2ZmD2vFK6b0x2BrN52ulyNjLX9jEBu4edneQcbVHAFQQCzQsoC
PygXwIHvgf6Q9KlTI5e5HE7ypidf5O16xe4qOmXr6VkGv+MiQdjGCAlray6hM32/
PxsGXx90tktW334By9kTCHvzILZIMq7yLwFIahPTNYpBL7vTMxWzxjQHL0T2Fp2O
Ijo6cJhi91EPiTa8VSlcABgB56VL1SmZShSMA3NaD1fr3awswgPKlZ1XR1O4gEFu
2sdBp0o6ky1tpPHxQJlWidBV1MfbONM2YFK8qVapoCy8bM/qBfvyQE0w2+pM1K0u
bbM9S7e51ySPKqFcSVfCPjBtp5LYvzOsjBTLGu0PIxoV63ybipaVx+NUp6FpUADB
nB4teiDrF9gj7Zbx3hnKecnIdXYYEs4Q5bH22kIQtGfcEgp27x1sumTCp95QgNKX
8WFvPHVOXHiMxkQ2+sW7rFvvXYJb2BPn565maxbUMy1AeUwOd/AVyDCcqXcAPKUH
AWmiEGaFa5UsSOx3cuuiNLuGfJC7uusxOyDe9D2ThXiGcluKC6QzegWSNc7f+gUC
N241YWC8vNHH7FW/eeZSwuLbFbhZhoNs/7w/LF377PJaKmCQaroYhvkp0oJ187VS
5UooWSlVK5/CVO97Lftp5Vcdtph0FrnjuJ0JQAdwDZ7FgqILcXoxPGVS0cOI2LsV
p6qqxPa7lp95vZXWby06yJkFPHPK3iWpRQEDJt202j8IojgSJv7F4mSNhs5N58EV
Sj9+pdu4Hftib1U6HxqO1kbGiEQwxyWdq/Xy+DnMZg1hUK+UOidGwQEHqAjK9IOv
UFa52lCt0SF5sYe0rVuoo2co7+ov5Lf4bocNSqrMNvfklLMK32mumXEctB4tz+c5
n++QLCnVeKahy4NPyk9ll00fPJue+SVP6tDwe5+E78ZmK40SEepNb+9c5ME5Fbsg
J+dymQx9VTw2kD526ZzWk/s8LS7Wf9pwwlogIdmhHb+En0O8rStEh5PEPQmJSUQu
8XfNuBpSe8UumMFRxK1UDsC4WZV4gFz0NMNnVoNPMzTHlEcK/fwefjU5ny0+w0Cq
JZWLoeLz9CrQ2V6EfzyUVgKVATiI9bGNuE2OwA628nOtU81ZLMGjHro/FZuv4Pds
EhYqcwqbrHsoXoQWyStLf9fsIXB28UY3NFmjxF0t0E/kWmb/t9bj9gfS9U9jsGuS
ncAHh/kp8bW7mifWTSA4RwxF1YFeEA5lFbA553hJ2MxVJNvb32v9d3fK6KwiuqxL
qeEGkK6tsqciYd5TioIoPryRELDvlYaUkoKwrWkBCbpx//fgTQNP35WmnBcjivya
gfmrYAc3x+Ops40iA46FTpn7dZY4ZRL8RtY91YBDzGP8Jp6jBF4FuWFZvODKwUZ1
rVOJaEnPUENQFehgm5Z8jn6k1theVOolPuf64B8MrMrNP5EPzc5XnCDPXnWuSEL5
fZNNsdHocnWj9HwfPU1aTF7rz+YFZDFANY3YAPQNw0EflyoBaIh/qQrSk7z/WSxo
KG5P0mLxdaMgYRyB+MA9zcP+0o1QguoLFcfbBGXh+KD/7CG6fWaxhvvv5PAKqWJd
0u7V56KaL2NZGjtdaiR2qAtAzqMMjmwbVeVhwHQ2AXCZ+qf60M1vQ3EoNoV92gRa
a/mkh5S2yC/3cyL/+BhQJZCL8lVNHbWAWc13x8RPYduSPE3rlQmvjlnTypDba1iP
A+QAA45F3vW14hzqo/DF0Juzt9BRDEAQEm3U41x0lYoFgFa8/BCq5NklE+iwqTQB
xx/f9HXgl0ytXDYOSu+nVOOPoKvSTUyXFV/n8HcBopY+kNWsuRO0/sFaxkI62sY8
qhsTcMZ4Zsz+yuXDKTmQIVE4z8mGRza6nq5biXwQx4icg6XgEzMQ6byJsK3delJ3
ycdkXBihgqCkbF1vYA/SmaRHcCmm6DFmg4cWqbcNSu9QTKx+KrB1UBm6ZDPU2Ixb
fRvnmp1UUSi3Z9e6/kWX99QxsUwb50Wh5cRtzTDeyp+EPT7fpSCBT6FzT19JhKQS
3gIOd+ap+iOEWvWnoGEp4Y9YrwUlwTX1PbBd60fID4xhFGqXMmzGGIrwAZW/qYPv
WojlXgyhnhGaYieY3dmhBC32+ZQGllot+AlWI1wApJ29ovC25BkaaRYmhb3PcXHE
bStEtf3QL+TBeLD5030HpFybgvpjMftIAuIX9Usri+M3ZVTe4+m4SyjgRVWUjrs6
YL2FEqQSwL6kXVl0XFVZUL5Ar69mtSuqHK7ZUPr1CQ7IwTmKNWzkuXjGBKX4j4q2
zG7RAiK8y+ZsYqHj32aVpfhGrb27myvJNi8p2REg3qpaQ96JY1FommHlok9+uDWG
VSmeuMxn8kBF0uu+4M5azOVnTVFBVUkFFtbPML0hnRwp/wrWNg0kXL/OD3Zc5+Fo
g400qFgW3bpSj9VSrEqiDKwI8q+UCKCFZxuumSX/NNZIu/xvAF+GZnE0CtFqGt+I
7T4eGY5+R8ugUMUfgIafkRzM4CmY+vg+VakRd3tvxCDQSp/UaCQdplw81N0VLq81
F5Oko2KkahZyEFupNFPITciGI1wWJNAM/UbYRsh55lx/j9UPgrcmzteq3tKhCrC3
T43zP00iDCR4JfLOtaiegB3qR0x8D6QqtMMkT48EO/q5GY55zCkhCKyafUWmuWR+
mmjLLu4EXZfwe4Gz57b2Zipp1i05XJSmTkOiv667drV3NPXHvngp+5c9PPtNivar
j91Y9WyvyTGsa8Wpel0C669dk9YB0GLqiVQ/sjDqfh42Hwf4VWDcIlnp2lUVwEq9
UAv7BfKHSO0tqJQ6oDCFzemVDCbBYZ8mfOkuM3CBRnBas/wabFA02sSTWy2vue7B
UDpDMCYkVMINs6p0Zb0fPBpXJC0jIsfTr0VRSFvobh7K/N5IlXf6xlMT64rN90np
YdhL4aip5wdeXWwlkiwwYKCzgs/68q/0ITyAdd8EJgJ5p5k5P92C0AwcmTLa971P
X3KYQibMnt/JpaKlMSVQ2qrNbn1fgTCLuVyrEXZqQeeBP9LQbcs+Cp+O2TfQVITq
JtkZdaLW/w7gZiFwggAeNz2Lt9fw00mNjp9dKD3jjVmGAB7qE5/ama22ljY6F1Hk
gKE26GAa9AVsAdEPXuRp6gJMkquDls9trikvLueUasXF8PBDbGZGGfVRh1t0MHUp
8WF1alSZD49xjeWhX1zFB/mjuizCMYgjbfQCp3gZJp2sdl6YlaPTjEf5B6WxCBwE
siq4P2cXGtnjru9s064dqxzbBXlRZaGhFrprlwe9b17Y1rehLhOJnwFTBsOgI4FO
NuGJnFlmGI/dQLa1Cc0ShkRkgZ6Y1akHwmnNSnlJWRE4eQy/2c/WCz2v9Mux+2MY
otrPqg6rWbdQH697RT30hiNgyulsQ1zr09oZL9kZpo9fbvOcT+SRLcivF9wJWb8k
VCk55W6WU0S5oGN+x3LH5Hmh1PfigdE+sbDABsXAWmk1/ZBhG/JByywFCVKts0GL
aFsMil804Mud3lU0UtZeLlcYOKhb4z6Dl9hKbqVta1FLSYkWLl8/r9XKKPyAOdzl
2lY4cO3ehppeYR6ELnk+A/iEV7VM4eCypaSBWGEfmw3z4q3+B2g6O1KM+gLcm3hA
KmPfBhP4bGKlKC2YVSjLLPWV26ZqDGvaPj+c/bc8DBp5flYoKIHq4buXMt0FrcfU
HgXK8Gmc1ywysa/J9/N4Z4ZtDFGkGwF4mwzXcAtJ6O4YYCE8v7GcUbgz9TBYWONp
NGfInW2oZ/4Xb0O0dbXzkpuywuWglfdX4lLArHsJ59e393OmM13KdxJarTvKPohQ
Brbxf751RedVSA0X30Bt3N+IX9SEP8vkyna7bCmIZztb5HyXJoEHs18gg9HHPfxk
DrpD8XD8wdXVk+Wv4P2xinsFybxzjxGxIwSJlm35LyjHrNuK7j+lEIEXe121I8Vs
rAhMWBkbv6BKlfks67ekPP+pIIjG28AmWWmqB914+8Azuj+ybg6yfcEm5I2HwRE9
fbg//JowN83Rv1IUps2VvZbTnUTX+4UayQxmXUHmjsD5REGC0RSJbe6OadH2Vv/J
nf4G/Mj/ZsnIO3yUr2WSRKIGDa2ZbYxLV6OJRhhzHhGe477l2j6dANhKXBYmvH7u
ClaAIWrZLG7pn0JMK7fXsLM9/8RNcIexCRAUva8684dzimhsKHUx72/WUJ5Mj514
HdC4aSXgULObe4xlROfu1dygNZqz4wKagHWkvhtcYWDCFPbmNJ5Fn1j6JR3t8Clk
7Dxe0mcwdF1cRtSAS3MD5wPNQc/LJzFrbGbH8xV5/r4jjp1ewEg13shYs/3mxcSb
AisuoCeO1tVQ39Exxs7BJOGG28KrfcfUFrBrA7Rd9Svub3HtvxUcezCEEd2+maQf
UMD9gM5p/mvtolZTXpBv06qsbBd2Fp+O/Gas1ehjIGHlgQhDbKZiTfVo5HG1Zo0+
ibCOYOFNMqAQfwcby24x3CbG0f+zvZ5Fd0cPjbBVPz8DrSBhA+J/7TqAP4FynLtl
zXTOngYkytXCukX2ZOZML552oNgcQBovmTn2FvaiHi88/mgJsQUicyy2RnUxe3GB
DXDxINPO6n7h+fHYFKpjCtMQ9mD+VBwuOIIReVqAQtFhfbd4p8kP6d3n2Lca4om8
j8aFY1JObYjU8+HklSfD04ddgyM8nki0bDzIJXhPdCRjrtnFM4b2Bs13pnRqTHMN
KFLnMVTKEPxr2vAC1Akm184SIhUjb+HmyZW5sNZcXog3k9JG5vmkLREwoqb54OPu
xKkrmDXkzWg8BXqRH9RDh4xh6pTY7iRcSe47NBsCEBzZqEiu21+oECs3g1HKZzFd
5PE9QGc5RNj4Yu72fuIVPMU3fUJpGsNzazqYlUU2+IE4nZ5El9Z/mfftYPF/EBPN
5VBeS/aGd8G76DhWpmW37fIF566FkySgUsrgckaGLg4jfoAt9DwfWi263CwLZ64M
BkjfxADxc26sOf+a2alcKDIME2jlEUJv+VgHZ7VHDI9i0/ngDaHaaUqutJll6rla
+nimv/4zpl103tV44/C+9zn2B/8C7/Fga7hzHpaADfRMsbebWbIlleKvyk3UF2d6
ryJpUa3aCkqAJoZji1zBCLi+ymHXQy3SfRa0ykFYkaysvZuBZIfrY3L9knYKhycV
EbQIIAmDlyKxrL7gMuCjQS60q13oKAJd+JGGlCrd/Z1o6ACVGKSlPKUDWzRaYADD
h9sHOBp/CVXNKyM+826X+ZiW3csD6sD96I9bzVJHaVGKoHAcDyAJfx7hRGHsQMXe
mHF5A/zGskkpB8Hh7JMZdXd3PXAYONZ1miI80wCG0Z2Qrp+oe7TGuk9QhmzGCE3L
75QAAlOPUZ0jxtvHxQFRsNIZbU95jBy9BwRMvmrgN2cCMoXXthSaRdTQwa1PtkGI
M4oWMIIXZlYkzE7glH9si2KHNP+BUEvLJw4mixytAujKZu0fRqwnm8XByeSiDh1y
pQkdttOc2OF2FUn+akb7xoUic+oxgOorlzBXTXDE8cvFMOOxUnsoJ7ClVT14iGeX
+1jHtxMJT0orz6PHcYdA+a4t1jH7broELfT+yS6ireZ3TbO+N5XQyhTDn/EiImQl
khKpsMSnHxJQktHABEbcfrBrYM2CAVY49qrVhN8AUklCLTkc4voWD6N6osmKSieM
gPde4IqBuSHYDQHH8ZTsPJyAueR6oXOKLmk8sEvedWz6gMVrN/j5tpRDKom0/+Dr
IziOzTVC+C7WYGe+uRyGaDPgXT8YbsXXVTJIEKBWI0r6K9FJWbxEPJM+f1ixgv4Y
j6oyrP33vVsSSYHdtu1PWiKr6qHbMj9OirGC5Lp9dOueGitSFxpWYTRB907bFE3/
VtYBrkXAxOcU4ju2gn00reC16DJ7Jsw/XV47h7mv9Q6eSRxSyq2yuX7GHc7w4ByI
FCtJMSeaj5f3d+uivXtF4Yx7M5RBtnEemflIGVv7xvVzFeLSSxNz+0RzBVisd6uu
xK2Un56mxdfUkIicb4eDp6kkU0ez2cB5UsgBF7aV0KrKxoHVUpuqQIi+JaEIc6Xc
XKVklYPw/R/dVMR3lvc20YkExAx8FoYHDqe16L+HhjvY7YTLHU97cQB3s3r8mg5O
ykqVOZDMTh5E4kaHnIAcX2jtm4+2aIJiaeRWQkFo4mLm8lbRoaHQCUQatjSg6Fux
DYTF96afRMoe2I0/d0fdAbNxBnWb1yJ0LlYTotZ9E6MEcq83jFwIptyNMfB2469D
k/c1Mk+YbTKeASmbnQWZTqeqDeJeA/uieq3HG4fUrXY8EX060Z4Z6BqZDK0BH0PY
sVonzIWu8wH7Rjq2LK6dXL6aTtkk6zVbd/FApiebMK+3VX5UkP32fm3vh20fqeDe
Dm6CQVQvTGmsr3bsrViiA+UmXqCkQd+hkUL0yYVMTIdwekhCdVoiGG+SRGAgL9Za
r2JDQpH1yvDrjWp1PYtQAy3ecGsOnN5nAP21dVTmx7QM/vBRqQm3d8oJ3S19+ZJL
2zyUKlh9VvAgxBRheSxGBqnVyW7jbGN4wtxV+cpbfcb/O0wXHdS7B6jFLyc9DzNf
qb/JBny0S0OaTTKy7F3XGHa8jwEln9+Q2KRVILc56PEhvWekTOAS0xcCpD3NCrZ8
1Hyns7hgStLBENkZDRTjRmil2k99ipOHSXF00KNWnumAfJ4RExLWaKBjW7NPTXPe
Rhv163PewmxbgszMUu4AGDsd0g86jO+qJLoKDH8ZdLnpkhde0iJY4OgnrByQS2he
VORWIVz3OGyu2qIeJ5X2SkY74wGw+1CdPXHRpCWcDedpc5rYuNDiuoL86mUkp3UD
/oVY1TkPnjgRDKzKyAuUIg71qye/00AxPquW2rlZB5TQnSJWMXyA0x2L5klOjoAA
CaGqipfdRdafXcG6Nt6vCAXjEpfYQW66s4CqIn2qK2FxWyPOHvvpIVwf8nXqXbcO
Ak3AOzPhUWoJwlG3sdQnugn23ayFCrjFq5gL+F607ynBiSk9iw3dn5Vkk2Zr8x/U
BYj4gyfQb2eTNGWHjJWl7QZJTxLB3UvMDAJwzkYK7PWodC5JpJVuQDnHJ+yQd5Yz
sldP0F7Mih9MDdw8d3AT8STIDbfpLg8nbMuKyVvwH2TPoNEs00IhLPWWeC3T91QU
FYEcTTZu3OZcfqO41cARoyScFBW6w4HyHarXcZCua3QxTU5jHwxGi3dJTZZa8azX
s6WduDPQpAfGBrQF6r/uYPJAzTN57XuKFJZ6sK73uLKoj5ezVit4uxEnRnwd42b8
LjxHeMTifbLuPvZBQa3lVxaVBDC+ynIWOXJG5f0Y3UpXDIlSfYvr3LeAxAmH088y
HeEOSDmfkpXuAEGZvc+WotMX0/I+XsmhsD3GUPKw2hOETlt5HaZx0q0fTEroeshX
FG982l7jRRcf95m5x7bZtQC6ixxNPNFi8My40tvMBPcgAJyLCR0mCb4nryd7KzXZ
v1NQNcn9POn2WBdPMdKrzGWbmuMRZWqflZ9HyHWIZKloUbX+5xDdyIfjUpifvq5l
ZF33cGGLU1OsXKJtyW9dZeavyOMxwe9crd6Dy7oByVMLFIjTKtm03nNgJCtMsOyV
9ZAWZ3Ecs7wcw8Xb4uWnIemBuES6acmhflkw7Mwwbtp5cTm3AXrDYLQiFhaQAbzL
wb10KzHEKNTVGcZVypV26psc9Vyl8775u93+WYIGq2OGHkCRrxmP0DEDaVZgTgP9
BaovLGMz9at4WgONEbXBmdBjvCUflZjj1nPMHH729hnFqh6wcDUY2e7+wFESG+ey
rGh5hDCaswp8xuUvdoTE4IL3SkPT0ZHOe8MxxLvFUQ5Ne6ohAzL0JmqlBgVOJ5gn
Z13WwCw+Xauv9/k+ImSQB2CNQ/Qqo2P9wFnqrNWQyNqXEifshpkPnwfyffVIx1fv
xTekexNFGoVo9KycJGI68mDp2+EHR9GRon9+zcBGPWAjBod883m29U8p1DvchyTV
fpADjjVvZv9KgHTAPKmmuys0EPqt+zAXs/P7Q/gOxbJMXx2CbNZ9vyojhJmlfI7X
2PioVXL1TBiCGMX/yutzQ48zV5MmPzybKYrf9BYJ/ExvqM3HIKtCfqnECAu3e5LE
ITxVEQpuz+EhB0hjrvwQZ4nH8rgEFVAgxtKMe0YLXp2rALRbOZTzkJ27+IMTBipk
3NkdccJM4OblnmnhpDDuxn3HhbMMBsK6dTzWsLULOS6lerPix7dsWYgqHw3GIFoY
90qTIypXRIwhZTejOvhZg1QK6R3s2YPYj3vj2RlocDkK0xzetjTh1cNNhg15nClx
i5KCYpGmFJRM0KDebRxSTytA+Bz9MPVcgtWdtWjGG354AxrGU/KiJ0iErS3C70Or
spmOdLadf3LRFimnUWMAzxaQlE0E9gjf7pav9ZwQ6Ge9SIJ9v+bYiqkaz/U/9h2Z
3pjbukGn53bCV7zWXstN5r+mUgMeND7eu8p9O8L1TjPQyt2YiEDdPvu93zTZyzk3
kygVDoZJdu5SLT0Z173mrTEMbGDacax4fnR1wDwjSdC/iikzShThxW6k95fNahYr
myh/jO9hheVzRJuiIlFa9TV5sv1pmACwYikpYrzodmKstMle/ARCGYeCwDdYHGPi
xGuijk9kSLbFEr44tX5xRr1mSzGhgziTc1/j7SNiJTs87G1qeX4ZDSpiRPx/guKJ
V9d9/BjubKB50Y8UD7Zg+u7xhygPx76PJHqxrh41j2mBw4wYnOblUmnPqtWUXwlw
oGhwOXINZ8nUNejNSJYaEf7Xv7WQKQ03FhcvM3c9DnLOv/AqaHAqN83TtDhSMLDU
SVxcLSsxKqgv2ujljC77Pj8oyPqMaJGTuDDxExKdT67VBG1q5tGoT6IwOrfGkrjQ
LtQbH1XmvRNazj1tIazB34mHIF7AymOwR95I5j321/lLjSxBi821MdBCInB9/jMR
9YHVfiMh2MGwciHKk4dIQPGTNRHG18juv2QGO5GZ3FHfiMbLwn7kuhDRZW0RGxAq
pp68bz7dYDEKJVMkGZux+Wbpz/0xh7sqEyWL3kQxVeYkoewU6wS4OXQkX1DgAVq5
9Qu4xE37/ApI37Zm7xVSwvY7GVo+iJkbyVG/ReU8rJxcg1/YMy1rVa896kS89OsV
obfJfmlsZPaOcC6VSMshFeldgQqssyafFg3JMDB4rsXvndbFPo5gO2BcM7MIWWFu
OHamzn5JQ9mGhIzrwMzRnaGmQQoKvj8WmGYmskeU1KITFnZKl1Qe0YGRgGYnIC41
m9n0LMn7VB6RU9eTZr/4eZp9gIBD4BGdXYIfyxNZZQbDCjp2M5s//zSXCPVpJxg6
UMSkzxVpmav1k7NHW3X2SOSwQDlKNhI5Fa5zWdSkvHoTXZRujfWNNZo5z5IXyLxG
7VD1Ls3aslgoIK8cU+E58Jj+6RBSFiNJINixFXaj/zZXtFEiCS2AqGK8kr8LWhEc
klf7oIzvoY7xcNC4PHWNQDNQkukLWOl5iWZlrwc3M7JgQmEMGg9hxXiOyg9N1oPC
fOl3xpvo4OK/i79lNmDB8XkWG4tuOcmk/7GkiBwvpSH3jiiCoys62Dj/j1Ur7ZQY
5skKw31y4iTquYcSDF7Wou3QGC2WkuXZVUu78B5TAAkL0Z/v5fMc15YPgH33ZDxf
oUm2FI9uEo/4gNacNUhujE1KIv8HNYAg7Cdbpum/eiHh3eLhH6TKOVmIwqDARVu2
BhVn+xeUHl4Z73B+A30bRGTNxj26XCyMk5ywHaJO2i7afsXTssR+1xVMPENF/Spp
1SuX3jQcf9W7OJjG3yk36Xn0uURmxzZJG/EKIscSrbre+mKwrPZ7iT6lTkzUrYsd
IIsdwPZCXBHRKy/IJbrPqiHDqkEnCgEJJpghN/F4GGykG7rFDrCAh2UiTPHBP47d
hfbKTKlKe/UQ5BGhC1y61Xe7ouwxjTKUvzIfbNrAboRwWsV3qG20Z6UaO8++CCGL
66MM01jvtr2GWBT/VzFL9hCi5JOCp93R3KeBUh/v/MwXvbZSL2U5hFLA6hGvPtaQ
A5kn0qRWNLWKx1KlaXJuFGeaofOufuBI9J7TFGZZk/QYno1TTasiQbt9ObvKARCJ
VwWxq9T6ezK8X4NzlpNqkTl3yMUVFZJrCyaIY6qdfIb2G6ss2C/M4bz5WRryPAc/
4G9fvTyhXX0GHod8QgkWPehh1v4DTv7UntvNL4LYf6igRzuLLkjPawqHfVC62JIZ
YZZ0V0nzUGvJ9tRooe9B6GFsT7ZqZsRUMHUpOhWzTnK+6NQs5XHSJ1i3N+/lDOsq
AesViV2QRSRWmW/94PnugQkjrWiDf0J7Jjj2sGeRd+BKYTCq29MvmNUbN8BhvbfV
Cf44JN5mPCZHKu80kCFC68SGsd7Z9mkYJhFIRKxp71zuRFAyE/wnmL1w2MU6Ipma
FZM1aEHBLhekcmWE4WBhQXA7OoxP36VbWI0EBKgSsgnt/oQ4Qj/3kXP24NwdMHTq
lO96VXdClloP0pY/0rkFwe/ofuAhlEcXWK3XRsjkzvf/EXHV9lQcxBkCuzOH88jy
trUJaW3HUBEsBiNg3hn7OwmId5R0b0jlOQuSavcom8QV92lyNOBlTroULpvknTbl
t2hkLYYtOPsAZ3ft/FyWoBroGmNGMjQqTfJqEeZUR9yN/WT+fnE176w2DofJQbVN
G0Rn9PEwkR9wnQzKvna7+oUN5tAqVmOcoYV2gWx4fq5Ke2Km6XvGn+QMecM6BwzV
9Gr86eBc2KYeldGroQvhs1ZO5JD+fL8THNSQyUZd059YKzRZTU9L37TM8ReghhYs
NEQIe2YCM8mhEOvybKMOK1WzIvhGooxjvSwP7DXILKfxKiuFt9lrk/A4nsazjlsv
VjNn6kGnkXaH4I2YYhNHLQmu2g39wGetRWDRInlSM9v18EWfyFA4WyDM1SSNfxfC
onmEbFZRqwJdhCWBIstH7MjHxmnhU0yORhj5kN9wq3rPEBqm7usCSFz5lVTmZ9eB
Q5hzLacxR6rpQPDix3xAPyTpM4G2nWnDT6s+xpKJgRWZy3xoaCNoKIXGF7E6U1oo
pZP7JeaCwVQngP2Et/mNq9tFSpkuhhUZY1fB9+In1KFoklAfmMqPar6a9KKwziYG
y+do6gJkFrcgBp+wbbtyo6vqcTxUPOKkBf3QXCdQdWI5CL0nREED1oZXPS9sAuxa
ovbMPdRMjWWXod3i+mNXYJYNliRaRHN1jIgNy5g38QGIpGTsEkyYSl0JOfIcc9y7
RB3k+o5VWG6c5+kFaoEVnP8ay1P/0QY9sxUdGVLwWiS53nU90Xd2rTaf5IOaJWme
New8PLCgYFeN55t31AsgO1q7l2VUr6pys2ovihTtW3d2npeiL+7mRfJcHugnmidk
skHTZwXwhsVlXw1Y9LU6N74XyVwWjw93ZfzCXKN+C8/+CHsUtj82ejaIcnUURABV
iJLT9t+xAcMFsUKNYhPSyekovDhm7j3fXA9cms7sKN/MLaANLBST9giP3TJWAYiV
cPmPSmts47lWG767pc0sD0avhfg1E8lzVX9LtDMMIMcwLoD24gonBjUZ7lzAnIRP
XIwYv1UdhkOob+gIAcxnHF0uQSXD4ApYqV8rZJK1yecED2McighyuBGY6DSZkaK6
gZmxQCAZ4BxNxnz0AjvTxH1MOhYm39lWgGRunNv1VWaY+JBETr6OtjajK7oXhPBb
8I1otJgslZRfsbU65pO4FHTw3HjFc61Hryl/otU+LTwylH1QbV3lZmgwO1+BrF1H
H1cVSo2bXTH6lznfzJHzufyIg1r37X3LeNbBOIQ34bDjckcxw/MRMAoW6NzJG+xx
T3ZDcJ7Lh7CBqYuNXL1GZLPEKZOtWBEy5Deb5DMwVUGs23UQn0qE0fLRvZQZdfA+
6rHXYlnQx9fQF/2tIuJ3SPSqxR1AV3idtfNWiVoSwPdwEmjt2OUDxiF03Sddu1Ec
aIpvgUzm/bn/gVjWHdk5duRCPCVwZdCAtXXWg+p+wBEOG1A/tU+gFovR5wkd+7UF
AqTX2jKmiu2NXaDVKu+WB3OsL+R/C/O9wpEPY+oCsaF5qznjbDPxrzKwm4SQRVui
EWv0Fv8XhDoxSNl7Sd5S37TZWQvucdgrrQ6r8dBjFgmyVPryOvvf/oxJDGHGwoP1
5/bKZ4bI1e0sn0VGE+xheCuF2EaESdMETXCO9ErjoCJv/YaLmZx5MydgujdzUWpG
ykzFls+HPqN1f5w+kZswAryKeuUS+gV4TNHkDsifZGspYtYzmPxAWdczDk3qYR/6
76Vhr/+l0rjYxWEMwAcExtHySKVkkJUYF/379IOQpMBDWQ/lGCdCDsDJY/WSXB+k
ZaSw/ZtPNg6enmuPBAq8s9PzJwRAbnAD+elgBTgwJ6A5Fk1ZugnNm/MCIHDpsykr
SA8K8NgUIzKyTPkN30+Uhikof3l7P6Jp/ctpd6Z35j4LoGp4fnvh+C6Bp+XTvnUU
Pbolz2TUDsXCeX0ll9ED4Gz/YIly7nkTiW+gUvfrDfkojBL/MEwnwAhG/fXx7XZD
9/5o6CfBVTiGgmabHwMFnTKv2SrKjPSGZlh2w8P88/LrnPDY6eV06Fo2LU57j6Mv
OA8N5ZxWJbiwF5L4JYzgXD8cE6XRlPL2vE7bpUwicWTTjtjxNlooB/PIV8qhEP30
5WxR+RNLhcJDufB80peIU4f5fkWVidQueW2Vfq7GAGBhQldzEOapPS8JFrk83olQ
cFaWsnr9TRJhr4iPcFFkDP3/TqsGSoLvfrNb8HsNrvtomLb6sEoVxukn0w68E3LE
e6aR0aS1HIYOBDl+Ex2guhszBhZUoTbHDbEwo38Mzc0GV1Uuz5UEVflAn7T7+kOY
jLm6PJkV0RE3dKBj4za4xI1fqKw7o2uUyIXAxm0xrXy+xHylPuCusx7O56QWOp0j
8blZ0+TIOnGEl8TucpdQqkojcFxuQ7mKEbIbtk5rpQxpm/4f6KBZdrtGqQvddJRT
CWGsWwyAQwqkUrntB0Tr9mHyF7OX5X0FZBhcmCloj7CJuV4MeJCizCJshANr7paP
Ger8JLOL+byB2xFGaxdfDU5c9A3v+BozY2kiJQVJkexYSAldrpJt+a12S1dbD4Bf
fbAJYzglSgvvIWT8DQ/EnWMH2MWZo1zBcwC0cAh9fK5960GEJAAvwvyoR5fKiL4X
2I6doS/eUDhVlfK2rarWyEItW9qNcMYz0kDQUTN+GSvDe+qoanGgvaw28QeG9IJr
BFO2xkZg53trFlE8hI3SI4YjonuWUr9y80SgWh4QQ/26ZGWl1ofFufeaPEVqai7g
9qwupV5ZiC0HowrYtWWHk9ysnoI1HX6Uuau2iuRP2TcS3kxox2EdyoQay7MYzHzp
p4vA6eRitzeMIVq/qcVsnXdmLiiAtMahHxvN/J6GLHxJ/WgFtG0HgFBpFTer2LET
1SJMI/FQcOzOQc97VM648Iic8lPZ1sDCKLcrIBplZmpRMWk49ZH/KNZ7eZOcq+i+
XcB0l+03cbXDDCzuGXs3mfh8O8HdtYfQDtI2ttYDD6ZtaxL9NzFvrKqSbRKubPeZ
hZNeSzBfeu/IQldj9LNI4RGTT1dbzaOfAEzSLtZ1RVJnxmXNg7dBV9izXZV+fLNI
q9QFOqsR/DWNigGQX5t8Jn0X0S8JHD3Hje7YNpJpPp7Oh4d59Sa9oMonV771MQ1P
zSSA/dMUKMRhe8Rxk3wscAgZ1S7tOdIYzx+VubzV6aFCwSQFCY9OieeOwYyDzrBi
wDEnihG8zOX910MBKA/tpsM8KUoIpd4/V53e0RfHRs4saih5ddL6p0JnMlG/h0hQ
1LWnA8DHE+3YH2ix6UKlLPDGrLdcoHbTDjvP+rSqiE3hlvGdNjN5kf4U8JUZyTmg
KFvTB+j+bvs854dQjPm2KSpSRa5ZAI7vYTqbWaCnRY/jCXONWYXDughZWvtpOYtP
CXMpIBasyeUSk+vDdAAADeCtYVbltCug/H8Bk2lKRHvmmBNxX/xlLyWkiObYmE3/
pyu/CQ6dcdP9YABu7OjkqfodzF2rO28o+D2YZmSl1L63WbMzeMsToDjKdozQaMUf
DMkF4vR40K4ODqTz81j4vAteyQR/t+DLuf0eJyEYPuq9HIymkdcGQi9HcY1xtby8
9AKULw0ozUZKfgFOgMp9ztzkX6VRs2AuTT525XozlxLGfe7JmHF8ObfJFR+0o+6R
A3S9tPa0Cbl56Yv/8zzcQ/E2Fm4pW6jRYPqLb1oJM/d1PeZ8pyjUi5zoebFuVBsR
uk8irVXBbMH9+9p/VI7yP6QM6QxAVk1RZDvBixueoELnj1ZkOfQDVAXHb0CWc13l
8TrJC1ywrSeo4/n3zPLldppui5fZ517QqXgZ+q+oXXpt0ySccYGC9eRmEEMJpwjq
HIIh6qegmQZV8RZvZ4Ld5uw+SYtmveDFb4ye+aUuIIh+jS5kC2c5IfnKry7fulqH
E7TUuAgxcy77AmoL+pOQteLG/69GNVXGKq81wQW7kH9Tvv4cjMuO+gU64BsL19O9
mr5qiOkF2BKovQOYXEwQVQ0J7Hh1u97nNhgTSpLwqZBK14oUMuU/fmJ/YUEqYOfg
wR0CTwkiPoGVSpvyNQAy05v6n0A+HdKFWkq3jK7i9QBn9gJHrpCWIRpcPfmISWr8
gEwUelxj5KfzaxSzvnSKSxqNC9baUGJStcsn4NdzoDmFnBukYp+hmzeHcZ+FIYaH
XIrjFaBNAKx6hSb5dCOqOvUO11dmKip/qudXI833yuDQGpNZqTOgl4vVrbQ+Ir2q
Hh7lVprdlZYvDHoM407rR4f6hkEXbXRNpSkk9Xbm3Xt4MGc7tVJzur+9PIw5eXkt
gDQuKh7o6a9+nwd0QoyorXRkRnlHIi+I9HKo5LJOONIHOFQjeIhB6o9k+78VnxC9
duUtu+GYxx4VSpMl3z/fsyQXYOJJEzVvJ5Jh4FUSKCZQyOIuJt7P1uV+/SJoh2z/
GfHM9WAqMf8u88tBvCR/0ih2GHzAGSPpz46hiUcY+Zuvpnzswa15O0fvx/gUB8vp
MW4ZTrMvh/2t+vSII+Yu0ggkyX0ZQeINI7KKeEMdZgjR1eK0++ULGMTZtKTdj9K+
d2q14CjnfMnkdezbHedAFfXh0ESKQF+LM6fjR/eiO0iHDRy5EZPKR8XQt/30MwrN
0lGO3RJYJoemFogKZN40oFbtmNDF5M5/+RXXHKXCBsf5LfSQ1WwQfBcmm+Qd93kW
Gyab4u1L4SClD2FRhOpI8anpgUspdEC8DZClX59ciev3kOyZC7YJgMtujDAmnOxc
G1+FnldBlQvafsPqJcPUv4zXSm9mxAh2uYgmzEPgddxlYmvpgHNjhdqJEo3w9uX5
aGAk9aDGdLnq2B7uIuV1cSVuxImy96/amDjyiqtj1nG4DJSq5lyire61TX14kUZB
gtVQ3h7PKIBFta77i0XTEnhAhfrMNIERq4IA1XSm1BNwjQkcIj09jQLt7xZrpvpc
2Ca7HJqVdNklqNrkhpDg2mn2ETZ7Ij6KOPL9rtQGywRyVdo206jwGAdmjfKj+dOA
KMaM9DWaql8LPpz2bhHC5CAv560AHrigsU1SIfW1+m7t8FdAQgb2nsSJkmgITNkY
ugFsAX7IIKpyPgfPvqWftEmqlJc7QswLsgNd6Tkp799XxsmF/16GqDQZo5UzjDWr
Zu/1FwGC4xmcyIH2Nvj5Pst+0WCuJ0TO62xYteHezsRL3M30i97RM22VnqmVlLXk
K5xkM6pq3d6L/COWv58ZUlktdwK7rtUk6gT8Kvb3Dkc0OlXb8FEPgjQo7P4nO0Md
WIeuHrBoFubQt3wrQlAlctWdYi5V8u9bYCLlHpZnz+E31Bl48S+9H28cPT8itrHk
OJT+LnDjsip3pg4JomuFt/bsy8lBam4yjMUHzBtrWjrmGnokpfPSuIz7KEm3Pyg/
wE6zaQ8BqBv/vb50slZB89H7ltx4gRv5Nbi9/cUWAUVkvNuWCIA4eMYrk9bd/tyv
u+ET71g1X/ROAwG6nvs7x2Zf1W/0xkFHuCEQT/CIC/rMsjN6fr1xbOk1WqN1EV0k
FuPZqYM6Z43R3Kk9dzqxMCY89tFLBsP6WZWxpx74XJC9nGeEpsfvvctTK56RkcX9
ABNWSrR0/5McLf6ohUWteXZX40a9XZaNSeTwt2F7rbb048GdrsyetMu756h1OQBs
8i0aeQv2qIxjp2qk++keu0d4WGMOG/32E3gnLbrK4h1whROn6VNjSimH5UKitsbL
B/NByOJfoGgs4rEYvjjgJ/LPnALEDyQ8VY0N9BmDSc2VxTFSMmcNj68/8hJzJCpU
wJWMjgNEPz6lH4e7VqZEp0IjwSb0AtYgHpe/lBXhxTDxE3Iy4jcq0jpJ5+5C/0kq
gwh5ykbmZD6y6A6yr9/8AfOmBfuDqoHSd1TyW/k90OTlPpzXt7+VDMjf4fvfxp8O
ywmOoZIgbHqrXsWYPhaJ+NQffw+bk/JUdJRWj43ljpmnI1lEjWDfaYOlNt1VAU7c
DEnwxMrTaa+UUWIH9Jmuf3rAWswCxzlc6MW4FkBnvWtAgWW3hy5hsqW71m+ikEsG
69egQS0rchEM3TdwN8Iy/5AHWWA/wj2Zy++qC+pIMzHoXfIlt5qYfMeOs5dbJRfJ
RnCDOPqGrGSCcPotkXHwgfrHPVzJmV9u+xEygtfhLdY8XOAPM6lEqdLXgD79ZEL0
QCmOb8j74dCIEbDfMRFXy9OU1dCry03thUSLAz5PXriAD4EORm4Z3c/NTPra3Zzn
QfpcHeQjLDTch+QZeU6+Fd7pY7AyogpLkXcyon6n8K3dYpjfw3Dd/L1Nggtq9m7D
R1jhYzd1q7fjEYrPjBcT2hJDLwO2kzLzgvZbgCMgFZR6EQSC1jf+WgG/OMKtSFZn
qOr32AqUuUSISE7M4vx6L+Nomt92fhwdgu78DWFAwh8cE/wm0RZZePIpH4gArtlp
XH6DYqzIi+M96cDSfY6LV7enTwzLVjf2BAfks3nWQbefjtl2sxDJyaJZrXGYgQbR
Vg10r0Zug5NCIJh9gzcoybUCKfyA27TFpqI88gikMzKbIma0dDBg5UpBp/lDkXgu
dRThyO7/7wXbYAekKtFwl65+5tgnx2w9fUsG9LBIR7RixQDNUZi1WAtVg0riYx+v
5fqo81mS7fAS1iE2GP6wKPU8u9Mc/kWxIh+GFzRuWN3dmtPEIymm9y2uw7cS1775
wEZzioZW1a/iamUImJyfpE8Ir/8+gPQ01rzdEGLaToAuga2i2xkf8VMeu0BFf1EU
7VfnQ12CipRqFQGJKjHj/6C4cJBebJbF5eGF5ePmsParb5tPNOZb5KikJCCM0URi
zKqNvQ+A0Bm1wy3WDv1GSaWnMtpSKdNbda6MuT7flY/B04KN7buJ1JIZRT7bdKGi
ZCwh+gE+QDAxx40OpotIr3dSeHvP9jTWy7px5nt22jQOdJcV6298XB8niZjEqhCq
9mHr7mSRdEKcWeQ+KpdeynN/NMmGeGgUxwQbVR8qHllse2GeQcAdnQ6WBtOyegWA
KpxEimuVOO0VTDiVVY1oWQCgzbwDu4VT/RuIdCAucjt6Rlf6mhpOlCfutpruaHTK
Ur34IgkfN5gSyylw5r2P0DnjdlO3JwKZAUpRcR+qBc0/lpOl8j4wTq0elg6hNk3n
bgqUI0xw0wIGyMpi2Jhzq8+9jwiA3QfitKbo9upKBd9VPtvOSk0KIwMUWcO33lWO
jNLxGjP3t7ZwGwKmJZaMJZxUnzpcPLZIfqlmbB2SvqpeDKqRcuhDmJwUu7svWYAU
yshlr1bq+/nHc0WPgPTVJcrWa/vRRuj/jnIloVe+elsmz4JrSKJqpQXP9FCY3qgr
8wPFGzgT94ZxfxKPLShaqV9n4hnHDXZlfNYYH03nM8WGWEDwf8rn4hXj76z68rS2
7haTcYPgioEWvGdUcOvKlSqtvRRtJPNmMeWUXOHn8B5Matj7avxOrECOD5a6+G9x
tUMIhGcALGaH90BUE9jmt/XDT42D6orc04SGBtwbMBqXBax5R1JHG+JlM3Vlfjep
T31a9stsTlEA4wfQ3b2YTx6XXLDT2eLMLXk9yX6oESkN8JEot07CBkMvzC9KK6TB
wBMwDBQrGv9OngPm/HwdNuqh56NgzvL/dHuOMX7G3NivwCsmAxTDTOF/iJk22zn0
wQNqBTsXSTIxZPm1MkxtBAMCQ8ZCGhlWS42EHgK+Tz6ymmOucY6K+WAO9KkYqmFn
2/tIVk/jifLkgz2xv7RFWGZaRkvInaOwYp/iNKG4GiViWzi1uwtkvpEGj0Zbrng5
r3FNZ2Rew8TvQ3wraXZrpz/SxfW054FCFD3B62CMdjbeUVXcMVIoYLWK2TtFDxSc
eB+FQrls7z3CrmpFrVfYfR9HxJZIiDUwPdVsPomSWdmr/W7wy+kGyel1rarT1kFE
ULpaCBrHsoIP8NEbn901Nr8H1IhR224hHnl8mteREoksdK0NDR7w74FHy37e6LqC
hsNkQmrkPciojNXJEzea/g7yI6IuUypPMnONjKOEAmlVmggiR1OCiX8SHL/Rg9Z7
FlI3kHeejsveGTNacMgqtFgUT48bDjMb4a3O2e5tD7AVBRBc71rN+NtnuGJOhPy8
4OTCjxFz8S2tQhayxAsZX6i/fmldW/r6khKLrrEn1heR5QN0D1stYh77/2ZDdzEE
sNtat7C217VGzwGeRWtEnum+ECpqg0FFh6E5vE2hgbnUgqdn4Pwm8KYPU8jcpQRC
SCmuvmaI1qBL6UHi9997nyRg6JW0HuZ05l7HPYe2vXpJCluESYUmEIZmo2icrXQN
Ova34IxV4yvSRes4WaQY7P+qR3F8xCj/fhwhAG8y4o2BVCE3TlYjnTXlyqNW6vAN
O6tAaSqASk2W/J3bNgo65jgeJkESYXz7AosnYPLXM9QUuukVFn2dK8X4Ipsp9dzw
dW09KBZBlyU3qzBItFjj40vmBI2yIOwsRImSGsofwyEu7K9eD/slmygQh2GpibKn
rajUYELJic0SrhwErtaqyuHtrrdd1cxR/Z0uGPmHxYu24AM7SrnkIn5xvaHgrm4W
G4ImvlKJvhPg7sb/jFnNXv2j+r3f8kvkiTD/aXWuZX8TkGMnaqXWkqCsGnZES1X2
mTTRvBOa6KpEjY3/kK2HAHUqHTPW1TR5SgEezwgU5o29EMtrEBNFvJuqaP6Q8/Kj
/Iu4azieX1xdSNgl5ZbKLTdApMlPtvRc57JyFwYV8ya4DWHGxsAO5mBucXHEP88S
pbNUVnHTJ8zOgnAnNIYdi69JmcxCzbUggv5nmMaEmwrvVf3lVCXMi8fmOh05Oo0T
FnrmUZ5y67USqtBdNa6hEoSVFRzArHcG7pl3J80mH8TuX+qY/NFbL5HLupCOpQaB
qTl4CNf3SFrp0T1FDZtnddcfiu3k0lGYbRvNedvFI2Mi4NrytSNEVSZtKPs6/KpP
ftKTrAbOCdSCQJB8I/VpK2vTNAEnprlYIb9L4u+bb9h1lE+4kzcyzC1nQewQQJpu
kek9CI+b3fmryp15HuDTwJ4oLAOaR02PUzRwAiwPY0cmqJQ0lsUfF7+rAqQKrjIw
7ftYDqoyWhdg+Z47D3aMIF42qV7X1pWUPEltlA9C4zIFNXK0cWNC9eEk8n2JbrRl
gdxL6V6Hys5zblMI4lakXWVspk5TU7MlatDrlZmD+gJmymzylGEzcD8q0m8G04fB
EuP5yLo1Z3fbPctWp6+3jCifegpuqoIeHmiLKeVFcjHWOLACRlCgRQ3V6bG84ESU
zJ1SP7PnDqwBJz0AUm8uMZYdfztgx531YlgTD6qGa8St1t55Qq1MPOjas9jDdbhw
diqk8/Tl9nysx8eNKqGKCynwXcz2WdWCAqMh2TMemeoW9lhcDKfPp5Boj646Bxry
/DHWgxyTnQcoqIfIRd05fFU/ish/EPc8Lcoxv+03zUqMp847lYE2i+oi5+iegcBW
1gjWMT7Ze1+g83kn5TuV2Odvc778nxl3A0m2i+T7Fh8RZwctUqUkE0fZ0eUtE2Bj
M6hS8NVNBCNFju7dhTYDR7gxaZcS5Jpge5BqGcUawHp+xp6/q4Zqjnd1A0mx36Yw
PdVV98czVzYPlnz9Y7qtu8C8hPTf5MMKNS0A3fyY8Mt/NUDtjD1/zRyGoNqEdM5S
BKFBBtnct5IynySdAOk5lW9KoTzW3dzRfA7+dlr2jX4v04lUBu6ZTL1BGRf1LGP7
X8S0zzcRmWhzyvR2K7E9PRHoRwUQymtgTk4lkN3uwbbpYNLCsz9ATCTv0bQ+TYQb
w0F33rw0MXNFTTelBYONLnwHCtL83wAxUdeaISZeYUOp6pnA+P/rVgx66QXgYYTm
uhh4yzjbN44D9YKzv3Nd1WlIh33wvRmng9aRp0DWbuiruoBxAsBUQGs7uc2vFn3M
1M9ZKcgj5c7uQGPML38MifgTJrBJ55q7nkQHb2mrIr6J7PyAdUhik6GZfU6HfH/E
WfuBrRPaRhZqXbcnnXl7K2JQMKc3rBoXBq/vtr6GVrfs8aN7v0E0RC4W9q/wCDQZ
D9PvqfHxJslaGQKdAp4doZE7RQabPYqZFHnLNIllQV9Vv0aIc8LrSZKZFqMnGutB
5qa8fHoInIyCqFnTcnJMPw7l2UwPHaIzHaCx9O4nsT3gKL6VxUkJOctr2cJTFshV
16ySkS0UvKkT/JrCQBeCzmJMYGRu/+xWUibC4vD+slgTfvSg3DTNuHG7Gta0A72G
IXKsLS/jQ5iNy2CQFHNXQ+9kdq7hHb5crbaFXrRngYqX3/SkNNd94CGaE3mNo5CT
uoLArYGyUhzJE9mEFltgGpiOs5I4ouVuuTlYXVgQeIzmHQ8oDLN6aYn6i0SSiRAc
3aildt1/braogJkfFYHeFYDYVpR7VJCMox1RpjTtKzt7D0BlYhSAjPOhj6pBd7W3
fnWbTyCHX4IxpfqkrLcK6+5IHoQfyOZn8i1/YVfIVklMveCPU6xv+Pl5N8saidGF
+BVCkqNn8lztRAkdowipLFgd01CDNbv1QgL+re/065dQvJ+yvir2YxETzpU2ELDi
sxv1gwwKV4QX6FttbJdimjnd3DUErTOjLjC5jQwmfba0GFDh84ZkHRk5a2veLCr9
4TUqe5/SA3cbnNoy0OkFAGwlvjk7kPMgACN/pza4acAx1QqvUlpMWB4WtAzwFrvw
m7v0PbyhNyjYuihWSguvqn4vkWYolOQ4gpgZQWfqLCLntn9o+x6PDK4icjBXOB91
jQ7v4q0K5j/z5RHEMM03wOQegQosGzAcmfXaehwnd5fj4b2nP+4eC40PDLqcf/PO
KeeoaKorSxy5sMceq2jkzUmUCjgknpRFnqm8Z1jAt2uYoVWN7b436Iqo23aDmZgN
38alxxMb/WETLioIyPy3MFyV2SpuC/SgAm5mZ+ZCwLRx36cyeR8R3WhZmfcomxAJ
gG+R7h/kKxCu1YEMWAxTnr/v6OPo6rd7oX9qo509Uo3lsXrfwFCaSTsDQvyAMpxo
rZXFSSBIgPM0cgDYPTw9skuZ6R/RzjRxhSJqhMFAuOWE5Y3rYJOn8PqJML1i19YU
CyTUZf2M2/uZk557YKfwVoYESMrdWL1KoVKGzK8ZnFn/aJ0jTzSdK/D+amdnipsm
YeDpA86HAyNYawE/1OV8ddqYc7JMyDlHv5S96MWwhjoCnfzlo9KlZeUxSM7Za2xv
YFan0NPMgt8Jpx/ZuxlSgt5mCD6uHLhhT+9R90dvV7nIhgbEcLEBoRCl1pZexvhP
BVh5vF1JX10+4L18TsEGBFvnXUjV7zJKVgkZY3H6MeIhVygXUASC+43Q2fE3C9Pi
N6fEbXUJMXKAJ5NoHbS5R0QsauROYfoA7ZhdDW4narsRBJDkGmAGXLGL/LsaZ+5n
QySMFmEMTH6iP6WNVWErQp10a6G7EUwnfd3op85NoavKCFgapGyXxnm52g18EsyQ
bRtDDBnCwdTNmOeKF/bSQdNVTh0zMSibo4a4QipWSrE4Q6oDAkUjvaPp3HcimloN
03bbLJxLyhziXx+8KP0j7wnyIC9vY+bCbmPBCWTGEJypRz38kPGNr54hteA5tuIq
1h4zYGGAnJ9DRyhxY9mh9q2m3Upq6ouv0SATPx7bfBpoUUFnP/ZEt6hRCNcB6Hki
X9z16PXad8B28G3MfilyqbWsQrfgiR2YVTMCnKcYRO/OFc/4qvUzlZGOeMHaNKam
qZzyoKk09KjOQ0KpmhC12uMX1AV4PrTyOdLLlntGZniwVO0wD0R0nMSsXIrmY5Ls
XXBApVgNmQMDPqd0edsoaZXOYvyQIgYua9bOsZ5JOqgGx1697Hvy8PcIpuGGRHAv
Mb7O7XxVU7uvBsypTmOYCSZGqWHXzX3y0aSxKHEqBYVlFHZVWtwJx9XUGmpiBe/M
ghcXUi4WGjwLV/MmyuyqMC4kDLQ3omnZ6WeCiFrKiLzAsKYUkSoGd+Woq/grZS8i
BLFdSYSr1plkSLN7Zq/QEW/gVByIwy86kSjyo9S00i3C4EXBA+Pwl7fHS5U/MDkh
RXg3jOECaUbpZgK4ZdijxxKS3+8cR9jVTUxNIYsIOvpcLwXgYkvmPFnSj2pShnVi
Lv9u+72d9WEznuBRTn8O+NUJDwtAwG8N2Eh3kpVYPpjQzetiJs0OSpRfe0V5pF1q
EmPjTYBSp24GLGqiSYKF7nW6pSTPKKuV436JTlMe2f3jxmfuXhHGxMhtnDLe1CCk
LEoBTqfobC8qo5RTGu4pKR+poBOJuGS9rvHAtT4JApeqyxxcw204qXvazOskwQ4E
DOcANxgu8mZwR5hMjWyhd3c79OzPu7dHAhCp1FpTWmEjSFROqxko7biegJ/pmYue
rditQKBCpojv0fgBiTWtNBbOx33NRsARpHFEBh5on0pGx7eq1giCKzdbDrpfoZvd
pVZimzXa3RfhqLbnlwmxueo7b9gyd52iaT1u+/avFT0S9nhv8zSI1RiCMyBq9F5W
C2RqPrBzA+OmuOR7KZGkem8OFjbQ5Ge2jtX/sx4lB4CliMWbfnuo2mtK8iv4Ulgj
D3SZVKh1Epk6RFTXJEaJwYam2RkY7DGDD1TSStbz31LLD7e1WTGFaHJoZA4D27f/
yHj4yRtcq2HpPN3g+1S3IroXEwTLwvfisqqyK80H/U5N4mikLzpcgLytAb3Tfjad
4vNP9QPhmLMltR1vb5Iaz6KLAVB2YYmLCBZ7/wCoy3AFt+3OiCf04ddeLQ+eehio
w4smcsdrrd0mxl4Z0v7s7YGK+2Dk+mVxWR+ded0L6UwFk+NcoRWHI7AWNYPREy9Y
AvuXlafswzu2XmY/gW+pwMZbHbPpZAwU/ZXdUCQgT7dESBTCnSTngxE9R/WCqI4r
S5GP4fLdHV7Vd4hdf3In2TsgvuKqv3deU5MH/dvtVdNHFUuPTc9OgjpKvPRZoseU
JxvHz5o8o+jHRXSKaOSAMRFw+U08h7lZk/ZmmJTB67rrp4NH8mn+jSuWw1VxR2JX
rd49l//BIVydIPMxKKRrPLfbBrqW1D070OeI8os4gXL3Y2zBPjczJRDpticbbzEa
MHntOESQfXyePwACTjQ0XrxEvVcvSrfpeZopVqh3YJb4VNh1eLbF7NBlvGEi0+bK
UaRVrbQ+Uy5gH4kmRBdS7ZSh8IqddibqUe+frHWPpxfjYfm5G7v2EufdWL0AGaxg
x+qhxmVmx3ZQFuhHxlgFKmPn35Mh9orp9EGtDnB1NYVKS/PpPFLbe//NPNPN3eLn
2t7VFUB799rrYtySvX/QXuhy2pQheoGxYOyX/a1QnJTKBsZkoBbVcnLm/KG/qlCg
hraKaBA6FrjQwuY7BaRPmoX1jhWMma12z3Z9YkpH8LeVkEMHJGVSZSB/bSf4iOow
DAd1GVa7eJ1IZSojpidpSwFEea3LRo/1cXcTSNt9HTPlOr3Cap45XZWKor/RFOEO
gy1ZYivIVUiGCUr3jCw4/snu7AJN8TzFHOzq2BoGIk9Nl7PbxszTvqp4Pd5D56vr
cxdAk/0L+5vnLKkt5KywlNIPz5NH7ZoXpIhaRAHcE63ep1ml67jgMlsbsGUV2r8V
v7opJlzVecyYagcdvsa33en3wjlflwfQbdqi7ErjBcpo0DEXb+kTud8PvHv+mI4I
J8eIW3ud9vZChJpdYzsQwNyv0AK4S8f/fqczOjKZ2ylebBAl9aMV5xNa4Q1rgnmq
FY4OQrRXVrRJHoJz0Cs5PWrd8jWEzUXqGoJX3ErdDLSIhO2YBBqyGFZajzXHM6F6
s8Ees7F+lOOuXhR/uoH4nC6979ypYO6k8QCY1871+sytpHEQs7arFw0k6Ce4dpgk
uxzx23JwzgOA4X9zQMb8x0hy2asr7kIrbjC35s/W2VQKs3w6ovJtrVxIH15knd36
KHY+rk7pFG6iY8PlEZKVh6waTWx8lcqx7OWWlug9ZA350YLN4pwd311ADMlUV2oN
4nnLo/sqO9/JelCJs8wmoa+JMfoPZ8p2wtf4gAAra5CUErrucUjFp8i4Z+scsTGn
+xn2RyTwBu1aFwgA9ploKohM6XdgGNDSq+I+LTF600E13mABjl9gD1DgRVoKzUli
HwC0oqikLlHQsex47PJ/1VbBOzoQPDJXlmu2tbSQ7f8/J3to1aWBNdvRAwsgJ8Jq
YQIlsC2oMVGegpSWldiEsMP2HLZn/Fxy05WZcK9iHaiM3Jgv5oUxO+KtEBRTJ0aV
EQAqUwFugdCcJXG/CDsXGD+u5bG4nCsoCyw4pCpAv79RXtDBSymxJ8d7yTOHTkkq
3FSV0D+tJfHs72fLKmTzPb3XJtyaYd9/VeLhC2rXoDxAzJ5yKIij1Ay0Q8L4dDql
g5TXBax33QccUSuWXat3zoiOO7eAGkGRvhX3Hnn0uEmJDn7B6L5bq2MltWn76R5u
vFnRaut9HaHc92eN5vp9XB3kHTZCvH5Lb0qI3yNkto6icFsxTtIXXC0rMpiTGvtz
QCatY6dMDAN6/yw7TGxQK1cxVAgobkzSqUFVu9cKAWHyPffetpGzS8LdWXFN0XJc
AHxIUQcJkOAXVwoVp3dqFXZ5ZYGGQTJ3RuO2DYXvIW25YzrcfEQwBapDLx3P9NJv
KlQyGW6um6TNMcRS5+4k1wR8Qv+iKYgL/IJUx0qUflakktNwCcpBCdTklX3zA3dJ
Er+FrzAwQnRgqotBPWtYQi/xDXJbO7X+TpBOszZ4t72Q8IhhbUw8IkEv4fdR4wM/
oQCJeVeMJbOkCIoMOOAurC9UYZm49a+WaC9soP+yE5H4SaqGswny0+yFt84I0auU
llgSVI6R4IU0Tuc0ZR8+W0obQW8G1jRTHbk5r9EMBZUuoOGC8iTc0ckHw2oCDIVt
EbYgBqzSnAFvSihRBXu0ToT2TNDynpTL+mKRtrtBOv9PVMqh3wRe66n4fIeeiQQ7
I9nqG1qEPhJj74bZUPzSeRsnK+WVYgeJDJRFO/MjK1p7wlH4GlT+VyDJ1+E52aOj
wwYnbkveLBHSLrfAm9kNE/i0iFnXOnCcinU9cFlzmSu4ttV288FN6XKECPkpBgZa
XzfBnb9DmKhGYSYmSh+06WpqSvgmGrA8T8w63SFTZ8538oJv6UfwSCbDnzLqmfJF
Kn/1WPEm8I4rqJ0Ld6WB68eKN1WIamZCaYCDn+tFLuC047j3L/vGDKAhelFarG01
94/D1+bdWaWRuCKK1NHJGAjt7mdkRb/OhoP/Cn2Y1z38JNqSWkFOA5JcuPxUV070
Xwak1/1CBnMPlUYCOKvCCtg+wQ+udyHsuQljc+lUS3gNX/Md6aO06gN+48pp0IDd
7P4zf7get/xLXehFhYXOMqT3h4AR4st5JedOWHwvw0ATRLdQjTtWudzZW++YPLqx
G6fDlWEql1ZL4Vej/BdSSE65eQSwIs3pRTJjnhlGA42yGc6bfZP3yTxlYo64lHxw
vYQEu55TSoBMwHFa2m0C6ejTCBXEDq60e4XcqJmYMLxkgLj1/u5pL+kE4O3bIWg4
NFTuycGnwYPVDOUNZtGdH7vOHMWOm7DRXA1ZxDUqa1Zm5uSojqOe6kb4IdiiO0pz
H2sI0q3kxHQa087lB3OF3pq4vKyl3Mw3BCkYDQKrY+HipiKYGMuhqk/0cEWRdXHp
3TtlPZZZo6l7ZFOt0rm1w93Kh0+ziVKCRBW15+yAS+RVox5BNcq10/f4caFXsWvp
vM2+pcx7hgBwAM76vfQB9xrIT3UXcN7TinZ0pq5m+u/I3CLKMQDsQEcEdxWSm3Z/
Haf95twgmjbsiM0k211wDE9NMZHpdDmBn7v83UPEaXwtKiVaUvMsUcxdJ7gTpW6M
0Kah/IwXKQfcZO6AfbabQsMjv5MsODFlCnhP6pXc7GPoAM0/DjtaAACzYS5mvZAK
0PFjsHSQqnMfbGCDl/e8OggqQnvOhB8iminh8LzkpnTWZzcyYFMeCqA83O0emSoD
gxnA1ulPGJ4j4eu4J8FvRFPpf9TRh7kgaQZtYWxRav1Yjni9AeEDS5gvy5h0LLIQ
pJwFZEJIlCUB4/3QLlGYUuK2bjC9D9WN0Dop8bwZjjtyQJoCMBi4Wbtqe0sXhmZt
Q7CbDiHBMQAfFlA1pvcQ6EpWW/ZqhE91zedsiLmA61vomiwJnjDXmdqxZxHvjtGJ
9oXUh2nE2G7yiqfm58B8u67GNyC4kO7DbgNkGcZ+CbJInTCa6nCEsdioTu3uYOTJ
ENUMzIFQtyUKd1hrsUBf/t4t0rsEiGenTCb6PTj9yFvJ0pesiiY8LZ5RrvDgq0Xq
R+0E3WocjMO2wC/Hjkw6v37pst7pTQFiqq4pfvgWf9BTZZeR0aNL5XCXP14UWqFc
sTupfxLFGCt9Ahx50ZFt2YKeXuYhO1UErqEGcbwPQ78xZ3RwB/HuAbs9QEAZEJKJ
2ck34SSdAxtB5fbdSRU0Ug4ZpckDNqxjGlQO/U/rzhlJvims5mcABDRShDvvzZ2+
TvBmXBvWmAzxkO9hsoKyNQeUis9gJGjlutzgrglh4fP3X04Hsc77ol0tKsxZ18Co
gLeL2vgdf700RnzkcWXrAwpXbAYdm8AFfR/vGJzrjHoaHJBdiWPLdmS7sN/ZDhrD
dRxaBWl/063UfOrzd/z0Xi3LWgRDnkvMdkGQQ9sdWqbR4tmTM141aysQX3qt1Isy
RkjfdF7x7tvdk/xNLXnhmNTGTvZV6ITK4vatBumVNBnDeG0nH8lKQqPD2lAXxeSq
c3oMB5sGqcn7+jgTrJ57zQznZt9BZbwtegXR7cWNUA4bPbQBSHJYFQszmfHyIN7V
2mG4a2ifIMBCbeWtZLGpvXjndRpKzJJdPC1xcsRSrayMan/h4aKrTkjzm8IKBYZF
vGYPhgSdEvv/nrtv/yX92NHGSA/LRDvggNWH5G/v2cmm37ehMkeBNdhzZ/SRs7oW
nQGHwTBAOcKQpr9wtv/KpqicriRTX7AdbSOBGYS2WeTRG2AbCWjHKXNXVf73Ug1e
j5SkPANrR5xEk+X1WD3k0BNv4h3wj0fzVwm7FOtgGOCo7QRYLTDfoI7LoogV12N9
zdltWQoaRaXjFLqC99hXPCS5u9ZXhGefg9ASSigL09DodxxltAixyhaF3WGNUjuM
2ebbXicImDgpAWN6UjaAmlg97KiL0iQoNUaejX0+0CcHV0OJQ0y2/SUuhUXIqx40
78I5eGxjzHNFXqUiSZ0d1duPS/LyH00IjVUjh9JIAUFhnN05rzBQCGHDAt96L+rK
cYX+k3phCslw0GQMWYS3znjO4jwJdLhY2CSkXYgGkciH7Lhd8NZMpEbTAXU3bof1
ApVABCZyXzwBqtg4rmI+FU42BVVQCnKC53IdmAORLOScPqExUfs6uAdCsgFSV4W5
XiVuJEZWYLS5hmhoQaj6e0y8gaFW4s+NPYWb1S910fuW7JdCdXK85MgNxI9HbsqR
y/53A/LBnmETxTt2s6SvUGmj5gINuTGembBTagsRGl2410pGN8mEmXq9dGtoxo3Z
q8kkRumESY/Q64h0TTuZ90HzK+NcSSmqTLhUmBkTwGXHsIBN6vILvP3J+0aNAKRy
KRRGGoLxYvvzGQ+GxRnzO/8gZCeGu73/+LdpY8tQPsyk75Tq1mCz0N1ltuRzn8wf
9TgEcay1i0WZr6zvrFpey4baqatrqDNmclpY3EPYZAdAhKrPBZYtuVJDYYcEFaIH
9urMbgphVpxwOWiXcv6TE7cQDNQ0FGXwSsyqrlb7BEVag960Sq0AIw7vLJvOgWm4
xa1t+9ZEZsT275xWTqL6HH/V59ZNQ47pRod6RftmzCuTJXhX67mOFMMorVflm1BZ
i+Gz7KYZM0snyp4yNfgMHPHmAkx3Z1zX5GggFMCJatV9lHtT4eKq0lY0nqWfw+yO
RLv/ifgtqaxWIhZI5jLDobVHAnB8JO3VCCCvL7EF4YFrVnyKvxvdY9mcfk/b+nqQ
/vpk2d3O+u3CCqrosBhiTVDq6opPUbWxm/vq31K/u4xH0Apic1fvBIgWDG/Pzvk3
Wdplxy1L/a8L3nWrct6OT0kZaxpBR1I9FiMuThZp6ewiDsUE11o+cWCgO0auUc42
DV3H3FGo0CWwbiprRrEubLoMF341lXUbkloa9Gv+s9GtpWfMrE6XKg5Kxg149D7B
KIoI/2KQM3laB4gXjwR9e6hELJfWouzTWd0ieF4W+teNgh9MKsBBi2dvgtQYM2CE
efeb3uf2sNUIZzz0zi1p81trm2q+esrXiuk5hq34ChJh2SyUNyJyyD7FiKKKa9vu
Bz73gfOH4HBvek5hB6OOx7Qt76WV2LIVEqbB27k7oGkRYTmt6OnLfrs+dP8zmfuM
NxzCwHF6QWqurTlJaJ7LFKevGyuZYUNmW9HAt++0UC0h4GjAFXDtJRL0YEVNe2T0
u/q0d+6Ouy1xUZov3KGekNFxneFxJ/Y1cEPOuC6OXLyOXVQzmPzLYJlkO+lo2X14
TkJSOX0VxMYItrW0YpZUkJIkdShSB8urIgy1ss7YlfjOZv9IaJgRcD9s3bB/nEIE
qDBO1UkayqPsh1RAQCccyoXFapgCVWN0WbQgHelqWS2+wdwhSofZYg7H13hKEyd/
tt0uIETdevMcmF458fA7RJtCSGyOB0muFeAwXzCCvO4yrr9uOrX4eDnw780YYMdx
kr3ZHnR/S/+p6d8+myIhkNmfSqAqixAQ3x4AbOhwY0UgpgVbxSlkiKLIWVeoAG+k
/HLCXx6pOpNXWU70X/xq6Y6D8FAwi8MOS0ee9BSHX2+Ik7ZbSEnLfGxHQpyyBLiP
FOmfM/EeSOHGLXV4WBay53Gx5hRa8Gt1VnH3S6PD29V36d0bhBfr0YqN4kN9cfrS
RLfK9W07Dr7Skhe84kG2QkWD3Y2u2hCzaMOY/+oL7ShzWTtSkqhR9+1zsqpTnRiA
IzLHLlAK7/VnLnY4BFn/CJeRj1GcMVWWaSoUqH+NbJBT0gOPU8RSUuo2gU7rEYm8
FSYsMwLFwu9RgkuuUcLQ0RTrL+W8R+PjMA+3q8l70DLWAVWfFL/B/6hggJ7JjN6M
sIdUJk/lI0R7Q9bcf+cpu3MqsdOYvYhdf+dEF+rl9De9CSitLkj+gLXeHcvaIuPM
o1wlIEiCFtaowa9cWZ5Kj274deLfEGenroupikqWOy4y1+RFjBXdfIl7Zv1R5S5A
nIbEiOgHU7QGDCDygm/VqmkR8RHKW9edscg0KFZmsabsa+XMjjLg/JoezEJtq8Y3
EDrejxDDiWsQx4sIPGkgYQ730KUkG+Qgv/UX+3Ads2saEtHkf69YIkUj3Gfhkh8k
Mv4l4cd7OrJD60j4/KipUBwrTXIXD6nM7E5zxjwPM1FwOstBOfGEzMlMKLb5Ct7P
SpM0P7oDDRBFV++TgPOdMIVTdz7PKsWYn0ykiJe5L8kwcijeCBGlG43qtVY2DRr1
FEuoimsJo6yEqRD077cImCcGlyWNkGL+v0fOTW5B/xfMoo6oOqm9t98of1a+7t8t
WVDqivMtG6gW8kD2NV7n360AG63WcYmVQf0vc1M3USWwykovoHftd8Mg1SLFG5tT
IHzf+TuOaV8Cyp7yHn/nycyL3A4OTD6bm+LpL7Nlna0nclWeiYuFE49ilyoD7mLG
K7sU9D4HM6CkywB12RonzpoZP5XRz4JOndPilGdwI7UNsv9vbWVZyNzJDHi9pU+Q
MRNoFE504vtr3drUF4K/B2y/IflrvBnP1BhkTthrz4kburtRLTOeiYRDN29wrBxs
eC3yNAmhwiZ/yWDGrToQPU/u83TCHIUFCPwd0ECn17zdO2tVnqOl2ZILFjX01BvS
pxlRPkgcD4M5a7Nb07x7hiwv6kkQdI2RO0P+B66i6o1Y30rycsxtWEXYfaEBxFTw
kuZV2YMI1ZhaWTUNeL+RH7j7lvfXwqOPpiYcm7I04IJ4izp9zaRBbYzNaN9YGKR8
fcc7N8UK2D8sfcRimJ7nCzs5QJFai+l14JdE9no6IoB7ZH5JmFGguY0bS7MAzYsM
hQaIzH+j686EHhn4eCbhVOaMvnpQLlVlcQWoSdGmf5EaVukxSGs5pbzWJv1SqbaO
s4rEEo8YyUUaU5A2mhWyVDV6dEk8+lO0r/UqJzUr0pnicz90Jz13mJZRgbT7tfmI
Mx+UTBx92RKRl47cvjHKPY+qXfaDYreEz2QTYd9vCiraZ+zYsUWv+EhShGmF64Hm
g31aRujStVtDi+VDrYeLA32OyiMQD+82JhKhbKrXrrGdLRbI59YJcpwBq4GbzGvs
ooSzNxhpX83YdVFM07mH0c47hdTFqESyCRlFI83bhEaUz2kOl0AgS42PJ68AxTNP
Z8xR8hXvF9w4U9zFzsYbDOr65TsRyeJ4G4Ji8h6zavBmA/upRMh8Y/8RjHCSZPro
UEUQeNEoqkLzsVFzHOVLg9HaOhUnZe8F4rzON0wa7Zm1PCGKhpHB5p9k0Wa5057t
OrlSLZizNm7XZdY37DTzt+p08WtmAhEzYhKeX4snvpa2VjvV1Z3n/YI8Y296IL8E
wBnbtet0WsfeQrZkklkCoatm2/9sq5Y859IKc2IZgZt6BfCme7bJnaZFClXmCzjD
l1MTcOcX3zlOmr64vccuyEbEIQ+XesL8Av4Yn5H1xKdNl69nTSFA6Mo3iByZ0aLw
TwgPAs1HEJvhhGaV/u7hTSdohKYqMoQx/cfm9igzG4kliMEpjvQWDmRyUqw9AJmr
QTayu1oYpi+DN5v8MZow9Z7RSdpF1MMxjUOWOltEBw2YRLIJlc4ryNSQ0l2Y2Dmb
TQnYCN3NoP+4R97zuLfrfTd4PZUL2Yf5kcCucXOdz7p/EVQI1r5VKL3e5UpBzsSM
zpg2ewNBGxCDbrTAqe/2BsHmICdX8e2Xo8wja3h/UAgJOYo40tAe6miltSlbNkCu
zrCL/gJWKcsUZhcxssEuaWAyBu332Mmd6mkf9ko30roHi9V72VJ3PHea7Gv8hrpW
pTN8zslXVkjBEZF2Yt05Nz3w6n6/9mbDuFyoxFpjSvisOVp+aJe28ROyhVEs5sAQ
gxroWgD0A/mOkOVVghRx/w39Y1XiNOIpOFUjAJSvd6q3bJo8z/OGtyjJH54D/VQH
/4zNVaboZz36oviyqeUPB2CaN2shDRw2gcxJMISc50sGeyo7N9BiLk4Tn5U/h3Km
7JPPp7oD0Uym5KpkqFdgZCpeCcxgDLe4elXncNq/61CPCSF99NmQoA7zOWzCTSiP
NigDE8Irc8KHlD4eOwQvu4XmDnHRbz1GLm70nW/crcRL6TqDASlU2I1ONFA33eXU
Hlsi5K9/5XjSONx8Mkfm1BmqzXbHIv+wxbcna1jIiQfLXwLkBCWPq1EZIwxPTJuM
6EIkJ5GvEF3pgi3aJciqUQ/8ms+SZjMgbvOP9W0cUapKaoFdEaiuqK1KKzzC91oE
K/4v2c570sLlG+AEJ82t/aS4H6gXXmZZY/Vzij1pl/OHqCcFjpihqECr2YvMe/yo
Nq31hredSyVPIkdYb+mGOaRduUyAn+w1l5R1LZiuEpIWRuTIX9QayGjABK7e+pcj
3PCYwWKTpXXnyrqcAn1pld1FOuUMlyUj4fAS8fPXuKrnziQrjexINrTbcwMlKuj+
7sHdqXwZwUJekiHs3UoGxB01hk4grH9mAbph5XxrnRAskeEETVz7kC1OH6+IiTyw
ajuUl5oQfSZaqoVfsp/8Hs9V5YQJEoqwSUGIaBf0ooJ6AR70kK9+EhWjbHbyOJao
OVISVwYR4K7+VKmBEscmBprKa7fyZLCOKool7tFH0ND6xWi3Ou1RSIvgCFn4OaKs
Pt6nckGeEkSKsddTo8Eu0YasUIRAfodrTCqMHN2jiEmuNWjMCVKN1LdKzqDQjmHb
vIlWwBybmM2bUMTQ5A6Vrhfa6YauoOYm581fDMUIXzDhq600O9eQH+dhna6vaZLE
TKBnS7a27rLqjSAh2SM0a58vBqKRfKRSoiGRUcc4ZuiQ0DybDMyw25+drRzo4YyA
OfIkgBbKUzPjBP/UkvlMKCEsUqY7nh8i87mtMnx8tC+U7avfiG7N3KSr1TU8rxLN
ppjC0K5a7ZRgzPDHbReD3v36gkA1PdqkARjIcWc3OcLXDAZyRtiTbjxOuLw46BpE
fS0RdyoP2AGtcOZzmpLDJ+q4Y7XACr76HlK8Cs2xKHssiHkN75o9sesTXccYIBrK
5QVGcRfPol/24KL6NPIU/x9NhdY65zdhRB7pZC23AkujjSXtnV2YM38OhWXOf/6z
VLnsKuMNJ9JiR1YEuv9D2mBuke9xDYPJW0bTEJEAcTJw5J04QD3jCIq6PWMzgm2k
+OQU3EYsZ4QNd5VHZEUveqPH+rDsOSoVcpmeuVxYNFjGaEsm3/urvKJbkwkOTngx
3DB79Gq74zbwj33VlcCl5DNNO1NkuHxbP8wtx0U2++rxUKoZuR96U1s53UX8foOi
8tB2P1G8mNHwMMJj7s4mA2nvCwBMpfueX1oB38oHws7nmoCxF8DgdXmgt/ezHy7F
4w9jhKoY3nbH4HKfvDWDwE+RZjU8ybtpjVjBAPSp9+JHnmmQOIpKxPGzKKfTh2Qw
1Df/qhh3BXnnI7PqZvJOYzDy/PPMV2DFK9NuDyvchrFmW2J72SXfusinb5em5/JR
5iV2EWGv3F6f/E3OjBhD41JRabyRaaIYJezY0rPNnRWH+W7K2KsotlnbficfsQDH
0Xs5X6gmTe+H+YSx9f059F1X8M9Sz7Oi5yNnPoHgTEUNKa4t57QxRLorc21FD9Ig
iX/h9Vz+lAXUDOPrfZeqDj8vlI29hnqBz49+HBSn5oWNbJXuJkXKEPGASmTrExBQ
MoE8M+H1/1rfqHkhDB09FlqkRD1PimTrXV5a82083EVNmlaESMn2Za7fNytvNPdv
/aoUQhr8LrjtXLy1VX7MxfAnZlJ9ltvR6/nKvyody4iMsF3slx6dvJFuC+y1PtgE
j+Ly8BcuqmSdZi65qiBdUZnzEQ3yuEy10jg7qfKvq2ExqUHgKce7m9qJ29VTy5cY
F3NfvlNv5/yElCGbbu5/uUx5CBv5HvGZWAgcQoVmAABt7HsGTgmZOzs4YYZWHpo9
pO6jADyyHpRACglZhnffDro767Gfwoxl2czZbzgeW5bCQAHw0LqWUZHZVQ0dsU/l
pOw427xdY4PX1x/tdiS2fraE7LLTe7isonfiluA5t4xpHQeznDxmRBbzxrpK995X
2yIUoCT1uNF878OBPIrr/cSkRjSWkoa8sRqpG5I6giQg9kCG6u85fxFPD0obvIUz
TPg23+FNhs+V5TapqCIhC0fA1U/0XnEBLOCbcm2IuH8yoAoItW5lG9dXIp0Cv4SS
98i1+EbCuw75kCKKaBrAc3b9Atq2xvm+SPPQ/umwKaS9QOeANvFj9tmWkPieDLje
SQ4ORULOq6trlNKc9plJqsh0aLqIpfIQyv6sxw/L6DBGRkLydczwjLz8JuULGWu6
bVN1eJxjjRqRMvOsGSH5ymkcQNaJ/Jzb2Qq2zazVPXMUV9JC2BZbhhN4DZFpFB6k
IJg9Es+LPVFmm/nCBRNsDhetR77inhUz3VD1wyTrj1Q+XoXRXXHUQDuMdwOdyqaC
61CfuGvHRvH49Oi3tOA+lgh48OzvbY3175foFR9uxIUBwLhOG8egxeQioD3NqN5x
+XE0cTxeEs7Qvjty9j3LUCOEC7B9QDFH1VqO3Bw3dYTQyeMuNH89h5Tu4v6nEi8k
7YWsZoqD86Xxk2egO6KiTzJilsUSugKIFkzeybIcuIY8S8nBs6uG+97subXqvqjQ
okeYAp9V5c4v9Eu8BKICfZNn2swC8aJtk5pUj+qEA86bxT9oZ7OBUdLqcf1Il6q4
Cr//0kD+aNINg1aOj3pmc4f8gYzztpA5LhYW2pg84RmL/i+CWAS2pUKytg8b7doQ
/RZrbbrptX4HHTtV9J8N7vqQ59gGZA/kYrZ9WnR5sjG2kHWCWVYlroCu85nCG2Cd
Zs2aOZdHbErZu/rHeA+rZ3ULor/ndRujhzukpS0VghtnF1qpQdPc691r0Zs3sv+v
+M5FzGSe95ml0lf47NIl9cJVIHiTnAlkR8orTZJhnT1WGwMFcCc3j+4LIVcm12NH
f9uDo/W64JmfZMkKlVDr/OZIK71IpzVQoNxapSzFWz4VkFZhslmrn+73/8NsWxQt
KFRthgvdVNgr7LcMPI6sh1iiX3hcOtwV4nRA4fhxb2mrMVqJNTLqzWZ7dE19LgJ+
sK/iUSeBkQ/eGANs/b6x3j3XxufPf4gRiejexsLU8KzxKZjUkSOt7/69kQJ4ADN+
QOywTcFqpQl/2CXVY2LdpiMyskuPPQH0rTDvWpd+9K/sN2/nnnSLBqquqqx8Psa0
uhfk1PljatvnmbYz6uNx7ojgXViAQfaZ7fKCMolJ0aCXLHgew3R4F0NFYE1nUdmb
z70zLXI0/PQ6khQ3Y+ABUUGS8vBDfipY1h4fl3DU5+REMqKY73nRz//sROspAhCp
1AlThrBeDDTH26U6XRiZfyMpzW42e6GCNzvhRYIIuF59uRbmgQF/z2thbnnQC6n7
E48xgh1vOIlcqfjFhggxx2rCS+MO3OMiOnWU4WfW+LQT8qnhCQK1nD6CW8myucB5
71R7zvH68M9dmjSJPwt11uHFL08q2iDJzFDHT1RtToKZFAch4sZoiGgvK9HBOU2T
ev7qIjYB3Nx9dWqGuB+/dYWHkq3uVsp92V+W+cxallrlK4l3huGqIoTT441jhnXf
jcAM4TpQxuMsIILL6vwdCGMbNGQ2uBgs+F25FDhSxMsed01sVMsUObwSHbXiaD69
u06wyGacRpz3iDomp08fQA+Kfk0bELONlUURMWwEpKNCn41UIaO7Dbr/BgSFeZ+Y
VhGFVqZ7m8IKhvkr58r+FHjsh78vlSInyFfeI3rNE6HPxLzWeRsY/gieC+GqDLsf
sWqN3GkHZ6dDpKIMLw0r/vHIAUFzuXUT5HltGBmtHpYfFBWG1tQ4DUuI8niAQEp4
3asuFMYDrc6T9Rf1xPhehc3LwQeLFeXrqCb3qByyAewGMjH0YU6394D25uZSt7aH
Ul7JndwGxa+IgIw5pWbQglS64PQUQD2uL879YrDhYpTJ6s6h1osfvdorLo96o28g
frEiYhnSNfasw/43StUBfKfwNvLJ++TW4zngmokkc5fbz1ETdZyyJAc1H1L43n9c
JZoiYwzV6IwAJz490RfGgEQ2se0hhCsNNb7UTvIQ4UbLgsndR1492QcCUsbGR7Jq
rtdexw4KT69SJ9rp5fj13PWfWWSBECOh0Y5PqEusMobS6daaHNnw5utqzhclH4vs
jTIeSmcnEA5hHWwj+dBoAmOLaOuCaASZsHTpKcJicKG4SdN2UcotM1J1p8ZdUskU
GpOvHllow7bQ+ilnCCmF3bksI70KS19kSWh3sMsQ0YXxMEbWdMC/glMfGYyDDTFG
ATBqc8cq6VJ68e4HTHlJA1oTHZ1esMzfTowlRYCR5/h63cWCN82zH8Sdi0EE9jSL
ZhGzL0LsK2qWUF6PNtThPk/itFK1n1NMHxGJBlFO53nRvGVPuNzzMmo3vmu/8nca
+jNKw6IW3RfJwymPOol0lqL6zFcKRlnWqP4I0JP5KIMZUyTWUe5bJ6NXxrvoDCFV
7hIZTD/up+ul7VLfTAebHFeOmr/2cHwrqmmPvpe6ovL+ffJTwQpwFNtF3D6MJMz0
RKXx7+CpqyuKVjxPuEIUOMSgtSixXan+vasKpssAclxe6Glh4NUzJE04mHLetJEo
iNFOeVkdp/VPJYtvflPdYYRzkkdN57/cbIwtY120snjTEVg1VhVcnfbHfUvCQNU/
z6sCHvJryBV9GezaKcAFj/++tdiZK3sVU8+M7BU3uheRgyCmvvoRsT9EMJMGB5tz
OFMn/LSqR0AHtOD5igTkqzi9ujzHKuGWGMN9342m6UA+3knnLbZUdMoCm0yQFUxG
0CGwWAnSDXQoub9SZhnRzDDGeghA2cvpoWo0ckuvfEQGg2XqEn+6coNXRxFK8KRa
DUBdMRpoBgeHF2gsdG4/GsITU5Q/GMSF7hRg+JdqJmrP6h5obZNtzkgEFSJOimxJ
TpAgeLWzC0l8Y9A5UQR+FKkZRKeismnUjWVNQWZxXfupDJfnz/33oAVgBwQZR5rl
CZLgFuJPeQiiJFZySKbDruTX8qi3tw839eV+24dN6bg/Jq6EB0iJCK+X0EXZ+qfI
rSmAgv4p/BMa4QaRJ54SKKmtefmrZ//1aaKVssftog7Gcz0NvjDb27D0Fp4kVE2r
hKBZkcpY5NZ0Rgoqa3qHSJOTmZcgYqjcfgoTEv6etKx7gILi5GnzEUQqP2bu3zxh
ymK/v8amSL4gSug8dqj3DkAIoVvmGhb2HJ0REqv+clkz5r6Q2l6Y6BBqbyU9wZGh
sgKVhzECF5pKpkgIcr/HlCtuXIP6e6d6elIgyDlPoa4qgDi7ghw9KYgZP1V+QC94
F10Df7BkJzUS4zM/Om/pNEMA3R0gVo6FV/nj94b9YMaDryYauboYdaJQvfkzJET3
YQDDF670K4jLccbVL0/1j5qyNloXJaLeqtDc085xe+UmhreOkemDdBc139k1PWm1
i7GL1AbBYvgpI+r75f4rktDWyztw7mMIf0tA488aDPv5Hq3hv9F9CH3eeW5drkiz
KoDpZP4mwx6ndfG0HVDGZbl5XpxSkebRr25A17odaNp7OQFJz/R+2fQ0YKo+avzH
y0XISCvk0vMh/TLYjm58qEA+cjnFY1YmXITvo/n8de4tb5ghSqYECagB7nJudSJM
AibBAiOdpgPeJwjMxdNL/fsOC/PvDT9PKVmmnH6/ACNVCjILH6ZGtxucHLvCM3q1
j0uuWAA+eE6Kok51bUCvrzliUTnDOSJuy1/2ZMYMxA5EukvavoJSDb1eN8qUYRSF
ghmc9rrTASb3rr2mgUE00SkyjpRUL+V9YHsFVyDfo+4t3g18Bj73eD5wDEWKefv6
BJb9pqDn5atK8EIWQ1p6stuhhuPbhYvse3TDio2g7EiBmZ6AwRtJAawr1WDpLTTi
xgOj9fgWuoNnOj6pGo3VZdduvrda+FPJsOy8+n51Ck0O4wSZb/Z4ZizTDafNy04Z
vQylt7D5H9tukBt4ShllMqMy65e8pzAoDUjK9E7LFLU+D04/e2CE88awnnpNChmE
wVaSaf+XLnTnWkUlnsOR76Xc+HuEyeK0FQYpvGzkDeq1J+5DY9Jq1sl1bwBh9DwU
OqmOi9lR+6Me/6xWu0+Oipxjfk8WDu+62fZK4KyzF+Jx4jkkCBAu7MA5qLiKxQBD
c6BpHmMkBAhV7X0//TfuQY6OnpxWzqmCtDQNwudpVfrLuAFlAHQOHwUmohSUCHVi
8Eh0TlMB6d0ZnZiVON6AzowMRCkQn2/aLpVFPu6K1R23aFWpuflJG/eZnSKNEjdO
Mvu/YJZS/IauuyGU22WeTlYwLUVhLeYszPZkvnj7RREdpMRlfndCZXg4TM5gbFXz
njxgMpsklBFm2ckBYawhbJX57sBCLhNp/I4Nxh22tXrShOdEaL5sq/lLW7B5Xu3W
cqKeLres89AbEBV22SaxZRwGunvzV4593h3qpBw7qPM8hJCutdnrTfWlyS0Z0jaQ
2uCZJ2zgjt+e6oDtHBpUVy1Tv/+9r2fbG3h2MVHpxJCZgD4rpthjv/vwARStyw6V
Q+/COo/pBA/DXT6d48uWvS51ZOFA5J0RsrlXmmc73cO6QBA8HweXFPC8VJZxxgUL
sQTfxniZO67EvJab/rtufOvTfhmjn7LKMiwPB3CgGltjgVOUum/igm+2lO0fEGJB
nCA3K8SP6lzkrKbwxbu/71CupEDuKuup+Tv7GRQCnHyrpjiIFEBZ6oNRoqbAr8az
F8/n7mVMubE++ZGh+Sm/BpW6zNZZM2ToC9pPplLvn/0DuZzdXl8Y9v5Sw4VIv9P4
yzmsAPsmjLkqwZp1ns35dJdUuoTjTwxpBSoILtSzlsa+G+CciAdAdHidCVLzWgoU
AJjWfgBqNgh05mIKqXsCaWl5iL7W5ONXRgpVhuoxNBOETKzzyAIHP7hjfSdY1PBd
czk4sMeofECT9S3iNOBlMMSNcgK6I/px/ooM7GttD0lEr5XcNd9Lc8H4pkWcikN3
vIpihHcYMtTVD6TJm5oWTLx8GYxW2V2ocuUOGJ1vDm0y9W3Re88bnIAMqeMXhbhr
mAkxWkbd8e0FY2YNIP2qLikTspIJRPTN3/oq7BZhkqmb1nB3V+vB+CoNNsG8q3rd
I87JJAyedr14Dd+3NpkPsIHSV9k+gRr4FV9vmVYwccQ5B7n26JgqKHiUJ93NmoqF
/O7UNlJ5SZ3dQLK/boFO9RHQy/31aKBhO/hjKqdbD1Zt8kAgJ8hHmM+XtKF/akHm
qkL/MPsWtHycyMBmrcUOkYLx55OhZ9LeBS+GDVqR/O0jqJb2cRR87k+liztz0gH9
lyeC+ugFJJZeJvs2+mJEiHhEPqk7yoSXaBd2WQbbPsZHHkgf0e/5oCVNPZhHAYis
gM7tuleKHTMF5+/TdhxRBWgl6hYzAWHB55n5dK/ggtp0BUG57UtiySFSP7pMJD41
BVwWIaIa/sWvAJ0oAbXVmc0saeMn+nuR4x0Qq53x6uoJ+r4qY00E6IU3Jkx6tXDa
mzl2rOvHNyIKAYwwuUpzedzYXBFhs0kHstiSA1s/ZBRLCZE+bM/E426RE6ZC5y0i
6wVxSxOTKySucw4vzOo/He5FZzcwZn0ef1NyLJYknMCosx3KcRyk7Zi6UbI1YXo+
F8fuXkEK3HsBAumfcPuKxLjmtKQjY6i5OfPaf4Izsckyo0Y2Cm0vj0ctd7pJkUWY
06ojrrEm3JuQcIWL82JwxJT/faDzUYUumwn5qxzh4jCUDKfvDrzskuW9/OgRmoVw
BV7VWTtCW8OdVJkWRYsNO0cjQ60STuQLqaks9zORpOVUqxQL6FtdcB9VqQwQ71hN
FcNAS45gdwvIby7N8clWns8R02n1KL28JqwejOkjRztw+UT72xeMcQ/fm4LwCOYB
xPq0d3a14CAzqP8YdpT2lTVQP3p7AB4C9od9lysp4oKQ0VJpMPCiABuETK/R466f
PL2gMfIKtPlwSR+yLCzM8YULTKS9D/XZ8E0wlJonMr9oi3cdc7IPld4YJbUPsddl
yMWPNgJNu2K9zO5kzBsiORY8kXcgCJAf7hUHHRFu0paugdKWNyz63YQ7TM74WN4J
fjEdQARGZY/acLBSNQ8iDAEurGiNOk+vSy8ilBr1gEgiUhAK1DdsuKQ8oXgkMX9S
iMY+vTv+7O3bLN683GF8ynHaGQKrPnBobAhHyDNs6aZxNd52wpgmZmJWAfbWuYTF
heZyMzutUpoVFHPDKtGPWHcjyUX2L3gPZGTyltUtGToAziMdzydxt+2uLr2uwvml
I8fMBz4jrjSS8ijmnzUXIRBvZz89CHYmhHBfvCNSr5aeztWUshKT6luOJNULHzyI
uDRjPVUiVlasEqXGiEyscV/KaRjLygJ4AlqxfMlE5XtWxWIjaGxJ49Q2e14nQsXG
wGVWF7uoUFF8qDtn6B0c5PAFmYd1qrtfnc1EV7D9a4CgJF0+bK39+aPeVxUJxFOc
fNSoEBZIrLO4o9aedpbhXBGDHl97h/9tOKwr1iuUUs6Sltidk1uI1SvvdjAcJcLd
1tXkuY4kMBSbgeC4Ip3ULp2C8rMy4XcUi3Jta+a+8hbtMT/8hTblr2y5MrHEpwtp
EvaV01wp64wdhPzHQrT8+bZmqOY3+ssXsDJSa/zMKQa/Z01iNXew/FGes81YkYVH
EV7jYZ1bW2p1/ehI7Xk/KuNf5T3aqMXWSqfATW1YszT1bvzTvSdfdTx/9GWSnpl7
/kjT5Omae6gEoln5r0AqC5SS4dPxVq7DK+O0wyCTryQINbnPv4xCTo/FJYUrTOPN
yPXuQhcQR1VKqKdRXiEHLxmPSLpJxiOkgBjSk4AFf6XaI6gjtZkToOHXeHXNRlx+
VN4236yW7SbOSL3PdihKeCa5FEO458YyCC9P8oYuEX0gX5JGBM22pqF3awxABfqx
UvV5n0486avBUupfyU7JfQIWM4U2FQplW0SPBVQmiMkCKdtXnWiOmudMdDs5grTL
tIUbbJCIbtEjm7sSM6Tsd2Q5VKQ3PM6n/qUFuR7FEb49j3bEwVPfOjYTUXLwKHOc
EvX1TGBi64iZhm+EWZkNIJQ45f4HBslAv/xP1KlDtYJGx1/SYdYYDsJKIgun3CKe
t/l80H2NzDl/4dYCHe33DXSxnHTRGUJEwujQaK08GZ3j37XFUaERnaxh6XFhUoXC
PBM5aJ/KzvK4OD/rLc4lOXgAgf7qPaDe1kXoYMWnQRlrOipySvkkIn94q8oM5wHM
Vf7YsHVO8jIjSxXdE4tJ8jr+s4PXcWQ6EIgBMjQ06rYdtlDXsl7OwhCL5wkJJ20Q
DbwX67gZA0SCQRNE60OhLeIOVP5rtNLR04fGgpfQ3J2Ui+nuXsOofNPOOCbGKfGV
++6ZZfBTAsstidzT1b/Kkw7fQ9Hgabm8miNWRRWgF1KwQq0l7J1tXWpqsQ7tcZmT
iWp7rxm/Qc+k+HSHYYcYtEqItbka623tH2ir/3FRfqFuiE5b707lhgeNYsmdVheI
rfNVczZkoQoRQAvQF/1HyQvAH9pmyIAo94mD+qe7LpbLjB8OXtlrNFulxLFOF3EZ
OvLgVU12jv1xYr3PEenfopxPr3UjTaVeZV8OKg/w6FieMVM5MJyX0CQY+GtaCdot
eiX3Ck7dMIltwmZwxEK9+eQvgUUqYoNhzxd8ZI+ADUYI9vl4+1HjdnTGRStC4lfE
1nYnsnrFpZ6Rmvkv1tTqqrVN2Oxr20LgPfzL9/DhiJRGSPiVmhcCGJsOC9io7lUc
zDQiPbEvqeUdWprTayCsEMDtSPERh8hMYMnaI+95PeDaan6neVTELO6xrbwRPKpa
O/orLkgG6mDCMffcbO9B03yeNyatTe2JTBiXy14JhkDzj27/iw1lg7KUInAqIxxn
emzhNWk6/fDk27vsOTl/jY7ErvcMNv0J35gYNR2kwJjvgaK3IR0c8GUFQYLJcDJ8
Vq3gosZuplagnmT6vI+k2BXsXPj8WD50z65n++UUJGfD/VNMBzUa7c6H4RzgeSRm
QGrKigQcZNAHVsW+q5QLYskmB3kLGHxuOw2DCd5pM7CFJ7HWBHL5VysHHZ1MswhK
guGSsiQaWxQMln0SbrafCSSge3VQurdoTA177xIrVzm+xnkSkFFdb82RIye5pFdu
88WJrtcAYWQ4ti/5QdwRNjEJ7ds64vT9fgbfINesJogc+EnTZs4eyCtmiRvrE7cy
2maJdQBRBTvw3E9P+4+kDSjvnk6IiRG56UZW3y944x8KQpqrFMQw0GDMq4Ty7ygw
FrzpMXbVvCEk6wwMJArduTOtrJ/ydKCAZpQt20GX6hvM7G4NGteUQxVOtC76wdxP
RC7mwxwF0y3p/imcfSDOpeEjqDTkRLOjc6kGIx2CU7hKUCt1kbzo3jsWM21TtbIZ
xURHsHtBZ9RsqDcrqnthY7MSKAm2plIFAc2QiAzLCUxP2dUIbLeevu9zzeCFor9F
x/lG6W/mj8bQUZleJ+SZFneS8ogdY707ueJNQ4fNKmrqJX9z16vKry8v/AM1+yHW
jDLm2Cn6sO/QXcuLDLuYtBFuiYFLyMsxmjoHstBN3BAnoKXh3utuqFK9XVStTApa
1cWw/sOYQOHrt+i2UQo3/FZbUyAHWsvw7I4UXyFQ0r+JJULCCiGz2e3ujRXz4L7s
NAxSVmczxahNb2CfMlxGPghwk3VEc2FmS0byv8udE6QXbjnr+sS4jZR2lfqgKU9O
jI19fiUsx3P4HNY5vVXeE5d6TMwh1W3KQ/fyn75W17njHBj/CvtWImxHAa6hlFyQ
gentx1r3xRuufUK7/+Qb6uJV0K9Ue8CVpFt3UcQZYb9eP2Z+ZaHGPZtbJpaZIoM6
5kS6iEZAHayw7iT2wDJ1CTxVoeOxNLirc4UQ6e6Mi3ECaXt9+nHDKhrS2SovpSy1
7AI3HOkwonoDKbSFXmnB5sMbHP5tCH8PIqPTcSfTdowRo8v8ki/zsvRlqIMCcDgI
5gb8OtYo4BkaCx4UEz6SHOn23eX5kkr6cW43BHc80Q+vRexOJZLGnhmaTZxEnsCA
rH3SW0vn/hbgnMLIXmvYg/X552JsUAEbIOFnaCem4r4m4Y5X0POuSP0m4+qYBv1r
tRh6z0i+pbIk9GXa56rmV2VHDSCA7fS1KLF/XCAv2Ejla3UTg2O1KPj/25hrTgFQ
4CtbQdKuW1CLUj0C/0MnR/w9R2MdgeSunAeYhonnU8kz/eNM4BulkU0CSodwoWRM
K5lOKc5JBjQcrRNptwYVeAQkqUv5DjfRdH56JYd1qNK0WIfI4RWjJ85RSX3hFo2f
pcegUu0BKWb0xEyYfsQeumjb5mnaHl7Wma+rftz1jcFY8Hfl2iOLJUJILrgoVUxL
nBl6XnmjV4GB6B3+/PDzh+Bl5KDduUt2B+K6KRZtegVgftQskKj6DtBwBa9mWYye
GA4h1YpIeBDxOQ8IzUkpghPzn+QjDAyiAQhaAwb8S95UJvWj++SyRz2fyT6MyHi9
qFE8IJW124j7GkrM8WLziCfEmEKSV4ycKMwz+kXK65DTMeJ0PkAmzTdb7zTHfQ2Y
IVnxh62/viHRltT+wY8vQ3hX4FgnkzOkc8bnS4lMDBiEWfeJViZkh6CJQ5SQ7PcC
GFT0n2yo360WF4NJ6lZVNCJCB/juHCPLjYXNcxgk+OhytZCTMVKKipYj/wTcdJ96
Us5tX0G7i5hLk2QU+h8pZ4K9/IfzzRCi6yRoMxaTBEPPzBIB12GM/F5FX6GS6rCN
VEIlpyhlCt3KePceKP5uhOs4Cs7F8kDLqGXUoj3FyJwrY3OdbRpHkLLSMmsXvDUg
iEqp/IZL7gKI5b/NkMc+YbeOVHvwYY6U6n4W1bTnALytU0tmqqyg/KExJ6Pk97MF
4n1uEqskPAiR2UgLzuVuTGtpL8PwBxzo2Lj40IbF15tUAU91GWiFErW6Uyz4Mp/4
vkbjXRmgz/bGx1vATfehQQwscjnNTTc9T8TnwAdhgsQulzKGzcroM92URHdNmVx3
HxG0sGLDeI3OW9vwD35v9JjxEjFrkE4W6CcOFs0NYgqW60Ll9ao1/NuewPuOb5hV
K/d5aA1YYXPKbq7W76JM2KBGVglWIftvICrRlEnNwbw8Kznw6czhZD5yRV0Xj3AZ
mHqpwNNpkgQvYKRAXBJrd0stY7E0wsQ6dADc1FHWcIgV9pnnSQvOh+n84ch+GCGs
0aMttjl5QN/GMSOM2itTCXqRdQgWORY0d0tmP+Nn+U9bAAi8bdPDX+WgK3VPXf5x
8P4WKb+V6QPxS+v4a4lN1bme35rh0cOs9fozJ0Z3zEeTIWaguiaiuGybqLX83yw+
dockvgGwIztBI7XZG6+g7AMLX/C81jWgLI0y1pFSIHRBfK1zxMW4JctoY9uDGuyD
xS9p/jGcRHOsbLxwrbDaaWsP/elMt+AaEWL7He/VHRTLTgpfTl2AWHlEqlGjlwzr
algFw9CW7c0a5aKNYQo6zgT0fgfDLnQdggJOAD2BCsudiVfPTcgC6X0gfFTwbbWC
Vb+owS/cf+D+cQbnZ/C2y65dgE6e2k5gnQi5w+xUzbfrIzsTOkPxzz5r8zBhGPWL
F+VJPT5+pbbAun0FHdp8azVaMjpAASNqDMB+2LlQBdUv1ubJNgUd6Cpkdw9t1GV8
hsjnTnbspJjlOS6rYfTXyqGrPqGzFAvml2qI2aB5dOO4MX3vn2qcj8L9GzjCK9JS
2zrIpx1+Q2AYhwJUGmqeKT9XnHS9SLfJPT5iOz2YYBnTT8kyvhTAz0xqbVGKi2kh
dAyEDfIrKOCMoan5BV4hATF00OZm5zERiCXa8PwqoqRW27qJZ+W5Jr/cdfirrJ8k
kP0BJWy38lbMnwIX2oAPdiV+Rnwc3/1VG/V57kCvbXyH6jNmxznmZRrfqYiDm6C3
2iaybPtTHyPTkySHOjaJKrre7YM+CJuvRziwzh2UoUHfm6t1dHzCoCV9qjhxJHEp
4c1GD3In3COdXsReXMt9NcESLS1gpwcQCyJPJr4570XVzECNpP3gXByeFeQLfmH9
cjo2THle9ernUCFurQXThSHJbzAemqzUFea3oqXI+P6fLcmJgNyl4s6XT2oquXfJ
NLMhUc0iZP6Iz3qnH1mcque+etDd1/2nNRly33wt2M5xndC4CPHkdzwO0EM10zDx
exNWTakQHZj92r6K8ieYNiEDumbbJ2CHxUc14k3yMY1QCSaRSQfay7QK1LqBvBG2
epuGyGCHiMjfzkp8H3oyCQq9n47lrYD900wYK7YUSOcyg5FhsMDfnIhEiAsspD2A
aQ+enTmp32M+XOcmHorqZ5O+tfJVYYtaiOgr2pO50qRAfycnUEP4aHS/XokYnDSU
o9AgG8ravc+raD9nZUrhtQxueCuVhLGkhLEG+T2chFZN5lgMt75J8DPT3tTb1MLP
1Km+GrNe7o7aZs+9rN4QNdFtoG2EB/EdAyYnfa2rYEMhlkOEsAJw9XSZu939ZSz4
319SDTUgR9QlEBjz3E8G7czFF69WbE1Vt/jPyjn9f+i+FbGDja/5UBBOsKMXs5VD
W6/C0eiBnsVXqG1sd/v7FzG+eLOKcXCv3UuTg5zmEPF7LhIkhWNNt8rUh0cIL7lw
V6dqXu4/2pkA8/EzoXw4llGMQ0+AeijHC7FUBakuAG8iR8zQwgtqPJUjeNFA54Sg
8xjUoFfu5q+L7EJspvw0EvJRRwvnMS5dlou32vzindnpSjI20DJsU8qo98zXau69
2HvK7rX4tRrqAUMdqRcAfD8yVCKh33SeM5e94H8s8DjbV7Mj9E5y62ECDkgI9sbl
fd7gtIljqocrUgGk/Ii5wy2NAmnPIgi94+VVI9pz4eMA778lZnMnDX2wXDNt+GN+
hLsSN4FGGY4ehhIhayqYmERYKKgGhNZKZkLSJgMEFBBqUBPmonh+CHGuOsZkZybv
W/dlarUPEOeVQWq1it5RrwNpdxYEDtXpZT0av335hS8TXSsUBNmdYa+yjgjmvGJ1
6i5dGjEBvFTK1ULBqb0Y6vuyt0k6kU4+kD48jwCPHr01d4CXycGHsDUkdurB3BYE
Gmm3V0D8SpPqgPQ7VYpwSHaX8nOE7+1w/tiET5/qFburn4N/PlWBol5fW9EDt3q9
wmFWu84YDbBVXWD25pNSzjblV+rt+kHMcpCo9ZRlcljeOuSvchBpAqkSy45phBcm
4dnvxtFvglomC7ZEPOdTf8S1qLp+VhnAVp5bRuaCDJt0x2va6eNp18dymekbP7XB
TqEqpHTlBc6tyjjutw9/j98S1wzqfy3uXF7oPMBKZ6j1kE7A3Scsq5yL/zQXcLuV
xnpRIHWLX/r07lA4Won6Jowq6H5bTRnRgMgrtzyArZqOV0eiE0G00xtvJFVae1IZ
GHQUP9jV28Oq/w48BZMeIhd5ZzbdDGJVfJD4UiyDa+VwiVrXV+16F0b8rTvSL/q4
zJIZYA/jMBeQyp+RBfoViz+rv5XMyYW6OkP2YQ/JO4MeI/2jSePX4YFkJ2bi+ZEH
klcrdQNEb4YgyIFnU2u/gsBNmii+iPcDyBM4qI4r72oIFBwwH/BuZwU7VPOM2pfQ
VxxHzFesKUQ/i2viTJvpvlaqGnI6SybVuWjrdIIHx/pChcb6SMUC8JexQ4fCQA4G
s9NJGKfzPQf11vDXanZSl3jNGdWsqqpwO4zT7nld5hqKVpSV/llQfQ2bsuSH00Mo
iQ3Ygu747jSCtWRopWau5oR5B0/KyYGawfCLAt7FyOg0cy/doUU5RIVTAOfj0LOU
v2aU18OkZYGJrrwHWbx/TUIFUoGtiIwp0u4hF2ynWsWiQNKw8H7yx9ulOCmOuN9v
/giZP3oti/fI3eXlEjYIbny9uMLKpzZ3qVfo4T6cAsosOcJhldT8h0fSftJV0XD0
FcTXLAbEQEeE1CvsToGrZC33eNal2UJjI3O3shHh/6O93dcDh8l+1Ajf2XGEPPqY
BnEj8cPdXueXaQuIFs+MgIPkh4Ob1LxvXgpr4U5EZDvzMK72dCUwpB9WoYAIqpvJ
pTCfZDwN4ThAgUMPO56U3UkwOQMLgW+bJ2Dh5ke0EE6vQzHl3tdC1yIbyqWyDIUU
XwBfh2jUzuEUZEKBZ3dwvMlUbUOaEUrAqQwDExa7vpazgszGXaNvb+46XARTgaTW
c8krCx7NIpY6ZIvEcMnelvPpkJjObgPTYPlHiWP6pq5A8J5ePlqfwJ3ya+b+789e
3Rrc18xqwh3QPB16kh4PfDdubJG/xP/Uuv+BUV8QbzDnFCrUSXs+pmNN9cbFWZoM
+ZnAUBiv2mDZzl0PM52dHg5GUWPaUZBk5qyifQBDFX4p9LSgvBSIQNCWC68224EI
qhEDDQjjaN04UzA+SBOfZjTnrbJwsqtXOfsFCp7EZ3/XxCUldPuvWkLY6kTXngYY
lF3o1WtMHazvOFFDAzliMS0Pmo4qzMO0VwVSA6+hWU38kgLglH7dCSjjrMZnwQOi
qQR5543APP1pawgix9OiblOWA7u6qGwyWRgkAOtTvlbBN7QeZGcB61wJWOSh4rRV
JS0Xv9H5f6YX+AI/O52mdpwsOS7IK6HoW5CecFFedw4+jXOh4AI2owPVy1e7k13u
zww7KO/dEpaAbJA9/PHH2i9HLqqOnRiFweQIK0aj/XT4k/B4dEQu2S8GEOTEHmZW
t4IHPzJBeWcsX7kaFJXdQTxkcIK7u48gt8/7DE+CNqkWBgu/dTgbbL6pMZLJyekA
lfLvximz5xSW4IJSLYVoJWBX1puGwBpO7HeZzJcZljGnFwXpSsco8+3efL86Q/Rf
F8UxKr+5yoXYi639LcwbebsCYo7ZgMnn6WY+PpffzAN0/br7JavwTpcHKYH4TS15
GqCjp1WlFGuxE+diNaZJgr3J84whT9QcwarbpTAJbjr6JDy5PCO/FNuT8p/nY9Gy
AzMJk1F94AUIFW5klIgwPlGIg6vb/A4qdrdDzab9qI0DPsZzGHlSGEvY2tdQQT/e
KiaimMPno3MMdVOBRJjRJYEIMb1qwtSWY5SLRkrYIpEaJ4kC9PVg3+SCnOnJr02Q
Rssjy6qhLRgE9ybMKiisbObPnLEVbDs81jlf7SugFNEe/az6d8kqUI+bSnnZeaYZ
HjyQhzd5DheLaT6g4X+2EHdLDdMIkKv5coawSgeATImAAF19NKEpZDSYQkcmus/+
TTGu9rRMYzDw3JiPWNtTv+6Um4e3cENbsHlcvD1Xb45VwhGpc3WDS5QWm2elPxpW
VtZnfPJ+sdUgEDBQ6NTgvGMIDJd/EsSwIfP6gOOE/LWRZzU5wa1/8c+Q5omKB4i+
xCegS6kQ4oToZhjbICIaTz2aO1cmj1KEEwa9CE+mC1XEy077PH+Ef7eMh4gHT/UU
1K6jKHKdCNehbIIhhzlZzUuGQ+lM9eNQT1Na93zltIEfEuh7DlcybONg0aEwbrgC
t521HEhpwSQQHuI6QoN/sXM4Bups68cTNF+y66AcE280JGdn7OI9NnmyBZ+qRE06
t2mwxkZTYQfC4Lcq2gUo8EdN5N+0x3YQUa3DXzq/KHkopIUZ+dcmZWjP3Ixqfb0j
yHbNCEEedTxz5lxNp6TcU+XcUkzOCgza/WImjs2Qoi9Id6eiqqXzPgFQqvbtdTYA
dasl+ecgIL3AFJx8kMZpICVQYAqQTxw7hZwDf9+s2u8iH9WyjsvBpHutTjFHaWy6
e6AuGMZawlSjgndK7ojMlKpghf2+r0qOcbHDRQqsfrmRsJ4rHt//C7lRNkfEzPwJ
tOqFhSE57NlttHVh3IdaM4vcp3yMRsRY/dlASu/PRMMB1/Fy+bwcmAUiXVwg9s7C
Urxh28cVJMdcg/mKPY7x37YpF4UeQEyeDwYog8V3peTv1rX4DqfH5XeG7+M47Z9Y
7Ni70d3zpK/N3uYEabclMBgIfkkhc3biBPfAU7zDNTOQCAgrK5Fr/VLfj2+qyezI
/fxzOHHadBmnQv4ko5TbqZ86jaVMcNyRQCR2lilLgLp3tEvj36jvdLSyGONgHLQS
je8C1bY8t5NBz2+9xVmyY73Fsq7SPuAu5HBl+GEl13DurAGpRWopCiZZQLAUVGZx
Tav87qx7td4f7aju0zGeolhHv553M1G1qVyGS/MBgkUf/MfRe82rcVII2px8NNW1
PAqKTE2n8ZjsSJMGyUkDtMecTPS6N1zzsi7UVMGUE0Fx2wplI6gKxt5tcPET3lG/
YxEOTmt/yw1dJfzy6KeHx9Gt8vVi9H0fXgeUETij/VRwowUvtuBDgzeLaPybw10A
XmbTlEnd5XdaYR050lkFHtdubwpmKYc/qk3nOKu5BV5cXZR6ySZ7lf6JZSFN6nRZ
szgRV7weejgipgwryIrzNVyOWUopvXgIh6Avq7qIAVz2qrS+4fgbUwB2BZHgsPOv
KDiLLM/1ElO8ibntwIQ5WGaZ5uaJgAe5r0U4G0ycPQiuGI759ivbb1+el8j/mj8I
ZH8D5iAX09AkHA6jkEKnKuUfwNe7OZvfQQ/LigMlACguE1PiYL+gS7UyHu0GVJyR
UnH/30kUhd6IAbzhGFsEBP4p4P+bJ2S1L2W37nq7wPEOodMPIAG2kBF6oycha6Cy
EDkTAqgVMKG8DYypIScmL2xdPKq8w7XIojld6VEXf8xue4WFYCm6Lqnp7TYl0W63
2RM52k5nw1RLrRQFkIhJZDVbKMp14f/strCwvQp4Jb8q7/Ts8H7Hn/ZaISnxusIP
urTQKVrisLUyZdmauZKpolQOOk45zmIdlLIyOiDRXUSrJPgTd6l5n7jHF8YiB84e
nWfYQFMsXMrKua/QEPnPdZN1CpZUPef0EvbgDBamnhJJuczxZULUlsftS9ryynjQ
UIL4mumHoF6wEROT98us0FVc8ho0L7wilAo44rATlCS1RKeH2SucWBHZiqBVdluu
YN6LYsTP6V1iF+sl1o0PoMNxn9vE3heIt9rttnBx1alTh8ZzbMtPWiLDY8kk76fa
mdy24wh3dVbnxF96/sHuYe7Bq5/nwS33DiaTMUVrncC2z9Pr0P676R/maVu0zP2S
mGi9TaYWyrLAe5kRyTp3VCiBUtKMia4GEcVkbAfPWbR+A2EH0uFPCkZF1d0UV7Im
USSZHDg5FDDzY4pa8gl0e5pFzizC6HKKcUDnZGO5HjWjJizW/eFPU1P2AXWpotBY
/Uh/d5MbZ4+MmjaJg6UNhcjZ73B0itvWL9+JVUchieXHr+LLbB98OQgOECf3f258
bR1dErU4F3aVcg0OcwXd6giHRyQ9gznP6aaloVdsF1QQeNod4TVwwcW9TcbL5CxB
XUJub9dhh2Ed0VgJLPHIJhM7Clw7uQYAHkueY++V7arzD7xnfGQq/1u6ufQAgNuj
tWO2m6jdI2UcwKYF4Pu2qwAEeXln670hDarcjzHhky6ovFMYMrbyHfVtjY24NjNt
/j6ipWzCW6OP+UEFcDKNwIjm2pwQ7TgxeGUawiZWP6lYetJFQBqEgxXo1tUD0QuZ
EAjeV2sj5xJltIFuYXONm4bNOx5fzFj1ZpPyjypQ/Y0/bE6K78c4Oin0R9KyGqtn
5njh8+iy6bA4RZjCylEI+3XH7z2pPouBIxZgvKL1VTLQj58dQ/RPXCavNwe7nkIv
Cz4fjNIjR0i0owgBxbj4DlOGh3ZctDMbRnES6wTnWyf7/q0chJP3UQAS0OlEMf0l
GaVEyq2h/KrEKtsRhaeknjMOi9XJ33U4mxvYKIJkt3r0iekHiMyVzXnyz/2WiLFI
YHYLwHB0jXbjY0I5srtm56AmWHUBm6ylXbWXPLlWievKWcVkcBKt+vZmQ0srwVGs
nRXukg2xUg3BYuCzYndGcWegY0QBvCCYn2INZK5cB1SVIaVowwJNZkmDz3eOGKmI
BVW+kqGlxJC4lqvv4uquq78TeACTGafOXXpbunqxUZwiLR0M3KxyzAmxhXKXIBwE
ypYow7nUF8xwkMWR08x9c8ItUdephHtqR9InwkqnWEr/ge4jakb/U5afItVjdbzH
pRmWWYmv4w8/vsCkQjqWf2/IzWAFXi/j5FZ11nIgf4V36I5/5WFDkmb+Gbs93YA0
HaQ+AK5OjEaDy1EJBFfbVGSu5VZr7cnDp3Sww4O6ThdmnnnjAAMVasx8w7izlNQm
/Vs+eDpfUM7H6LQmbd6UxjcaDCJoVRRJutDLyFHha2ynEy9LIcEEho/f9rahuNVf
JfGol2hGNalevwY0EmdtYrxD/kIjuziLkwm//63q3WDcTyKDfkxXS1LH7fCdB0s8
Sv4uo8/y09pfRk+JDT+4B2zvffdHdqO+6fp3c2gcARxPRt89OjdfIyx3UfgjS8NX
mfYoZ5kgjiDXxM4nnzrO9JZXpmSpwy1Da9e/z7ucczZc/rwR4qLn0SIPpRBdblb1
k+OLsSusSIF9k8daX/Qh7IL2vkN9zMBTq2nYIwe7pFlw6Ljo+YxAm0RA4SCg7PFU
CJ9SxvjhU/k6o/gjTQXJaGnz2hxyS/NRfXypXUf1IMb/EZIPkryt3m9NovouJK/U
WPNKx13d+EfPSUb6QtRVfUHyK1L0PLFWxYyV9CUMYC/0KqFjTuwQJkpC3H+2Pmg3
NiBjLIbidFacxIXjAiwrjmBRel3cZvqwykTfEYAKNMowwXj9raBNX0qgSNmZCD7f
RbuqkQ5DmUiUrC3Oz8ijZjSju153PAlq8U2hCHLCIOnvhNdIGYs++ud79YldC3gR
WXkh5sg5572RSGoUscsenwpyH1KvIOFX/QbEZ9ndP/8XtqGswK09d1ZgO6UuxDjY
ZJZayu28lT3aa92I/cGbnNBBDM9OrHhsIfOY5Q8gV3HwjYtdOQRlZdoKuB9O1PAY
tFWrNSEQco5oYhaX+zrJ5jwTrG8wX2kZ/mvHBj4bK+Y0Tkn57rDOS661ji5oZx+V
iG/a0tLphN7n/+Fv0dwkPs6LaEy9ynkqchsPVOAyRHFP2pZQY7acMlVwV0N21NT3
Kqhp3sEYW0SooZImnx5cNzs8u2NN9h5L83ZO4LIqsx2KswhvVq5rPyr8agLKv+/K
O21tdJ5eDyC3nVSDAGzlxdH7MSlG3L9t+/Hp2AoZtQJ9rcf289EMGA1XrL8bKxA/
Hf3GY6DQtsHJygM/Mr541RGWB4sidof4Gf+Dt29hqEuqkWJ/hGlCAKM9JtKREvmC
neyYefP0h7GG+PxJJ7WVDbH+LdnOklFq8zsEY4EECURzWviGl/hPc8w+5fb2eO9i
8XW2PPbuuEAjQYtaoyMEGM6qF2u+Rm+ZIGpDny141t1uZcnrM9arqZ9856/vinWl
nUFzshqGeeiD9DILxmnGpLEH3662HIpG6UXnPbLMcIGicMt49mDsnbWs1D/3BDL9
w7RdxxB7z5yKr9VbVqsakqLqMrHlUUFt19xq2iLi+RdoIyyfcbn5/0HNvoexQmIw
eB9Iinl1py3wO53kg2ftyQV2t6mVqg/2bvlFhl9LJ+jLDRj4xbQZ3pqDRm7KsOFi
6srzWrji7ago1KTKzKKd8Yk2AJsnw1ZYc5WBf6xb3mz9VkRuXB9iNHlFrwFyQJWi
e9gUKOQe7SptQd+ERT4/OHzyjAmDCN/X37Er08WLDkC2AcVXigoduoERvb/GH/G3
tM54bp6HNRfV3P44F2675/FX0ca1DqZ7L0ypuXyuwppU5Y4wWBZZ3QlfwuadCEJ7
4sVI7j5OzwvS9trvbYbrAuxMESVUeXUiRBRW5ddL93t/OWr/sxH34W2Va+QrDImS
BI61BRkLYOKDre2MkK0gKlea3H3Vv5R4/VurMfJOQWopQhZtlLB3eLQ8gJ4qp78H
xNbfFal9Y1BO2Bm07iM85eW3azWftd3g/E3h/1xlxVc3vB2HF6iohNR71ZCpv8Fa
sUroq9l8TsRlojr5Dg394PmYEqL7E4aTjK39demn3sznooR4fuDWfrlVlwFT4yB6
/n96IYtwj5Hj2URUps2x7NFEY2dZYVWlDRYSnmK34IwpkzifzhmwkR3XNFQTwdUv
Sercv1t9RkzwxfzaxfRdbWfZ6trCC3AcFU0d4AhVqu2gRCAXb8jRLTSJAzCsn64z
z2EVrVTgEzMHFjo311gjZRvyeMc0Kd5Wl+yr/DvQReZcMWmk+yn7FPDyJXv2XJlT
tWMRNJNW0xaL6hx660l8OcluToOkxUcNB9FT8jYQn+bNyE3Bixn2OdvQmD0TxJBO
K2dQM2p5Z5B03mGUnbPul60QGA8XtWAjILXwIXC4uW5hPlbjcHL2zndgNQcVvq08
ElZBseYWiXlnSR8qB2dDihskn4xo5ihc/YKMIEgLmPusyzun6AmcKXIbqr/DUZQ1
K/Rh9vwtC0oenVGYioCCgTUdrJp6l9Rtf/8tjG68ixi9lu9mfEp0uPc9fG4NhEkI
gL/cCRuAuqMacOW5CQhqgc2FCsS+G8kJO7G75ARXxuFSaHCCvS1QoXuiMtt5S1rD
dyktpigYDzGvctui8qXDJaAA+L8kpRGiKx9jMjFkxJ/SC/9dXHIKijZDsrDOxfue
XE8AaE+wsquGoB11B6hgC9gJWRZs+CbkHPyiloPtzWLb0+4nx0IQt0mmD7qb2CIZ
lC1wBH8GXhlTnPcZAPQlh2asW/BSuVUQ0g+1rkDTvZepMRHsuQqpPJkEP7SOqTUz
4Ep0vLKHI+BJQ7h0XhAEDzbeFEmoGD4OFl/8vpy+5QMSMrVDy+52ipI5yfx42b8c
UimFzJgsFNPNNJdOITpnltn2rmaxjoosuKennn5LC3eW2lyDckncuxOe9aFrawB2
asXiAHCOaskLxgmtq03nSVc5nTX8fDs+Lu1YA50NYVnMMjyUWxHhFjUR7jyVetYk
SoEdnnFwX59Ap5nQb+Fbhwzt2jwrvRWCYsYh3jyg2Uv3WexsH//7j4gcX4dE+YND
1Cud43sfo9GZBwAZrvhARFwSSArGi/J7GBEOtCwbHvEJ6vMXVaZSmOMufrljoRmd
04KZBFZu1KrVzMrG1v3w12WPwnu44tLdes9MycjOKBIRZUuMiHJu0zftYmua5TkR
uEmQkQUH0t7+uMeK6zItWNqBgGfm+irNQt01fzDcT2l/MbyYW2yQwX7op0Dz3EIs
QxRp9EqJ0A6psYcTUU7kb7Y7zYbDhmi0ieshzL0RfKCppge5JHOzkzDjeBbYmyWX
9AMg5Qwes7pymjbORVYsg7VBmtQ1Ni2oVYbv9U6aqKT0RMlUXQwDmDnm0ir+V1Q+
ufak4V1GfHi8aWjgsck1LnV4cbejy52jWTsdpgJXERg8VVL9oJYb5Wji4/x1PP7w
+4BBYdx3VCueS7F6/OjruCnrYFV2DrCWgqDTRJPmxfPZwkRIfN/VYo30vxo70c/7
jDbitfwhqLfMuWd5+YAOVJm5n7pPVREOeRmUW22H7TVvNFdEiQXuHA/sBgdZsmoa
myJvLH2807G2QouiO6xtfFzOldAMXNplgTcxD118cKWah4yI7oLtCRpBAcH698ID
hE9WgljvTaBnLrcch4QZTJkIH+lGuh2XLvxy4LXy9/pkct15YCcUJ4euYL99YQM9
+cDqeRBomc1RNXzD5kcWToGraAmcs1PSkXUBdnFus4tNosUZvssOR2q4f+wpdxPw
VUUoRYMaVI0OXuswo88K6/WmjX/vYucFVNrVMc4M7s9dXh24kvqCyqZBzx3TxXg6
aw6dsof4PyUTsLE5DFvuNFRTdHBCRa1G1TWVm3PDFlmVlqP+D64cfd6EoYCEGQmn
XPZRGcrwzGHA1w2yPyH8aiGd2toOkfflbtjC/RePn1R5PwrW/7+OwWC1azWzgOke
mljvvTRDyIfutX2vhWvgbjJ6NqeMjauHPFfQEc/i3lPZaoW/Nz8nGkfG7v8/Uu6B
80MjQK1OcFiM4I9WtYQC6T48RTkjRkTj/DUI5shWmlqbHQizETOv8hbjPJKrJB4L
O9hV9Qf18x8xZ7B1WBvmLohlFH5SRO0afZ+w0zS1EcdVneCD+Daix58nX8OPoiyA
1V5nMdSaw5ZZt2DRyO2U6lMMaQ8+rbQL5H6cIL+sBWK8PHR77OVGDZLTOeTqURBc
V+0dUSNK2hjRjh2L2oOYvSAUTQOcjumqVKZPvs4C1RCYtbqv9z/8z1nmnVYpShbz
uixXlkGcRY7WM+qtkqH0+xLk9Ko2iRybP7hZVgvgyuawhFgrOxK9e7weapkP5OaZ
Rij1HYq0zI8/92FwB4/U2KY94qGYn9yYmiwkjJp16V5xa6ZeWkFuL9D0jfMUm9sV
om6AGq/jRWu8gi8mr2bfRlAerMmFhncxS66/kDYjGHBMty3N3vahBVxiNlXHf3oH
eoKzCx8P9d3cISPYZwYbUKywlTrS8mIBak4xynDrSoRBUX4VRzBWJTlDSWjeWKjU
lZhd2iMySgVqbnHm55hsIDoiUZhkW3t3wayxyToggJijMRDEODWV/Zz2TAnXKafN
CaydkVnPnGI+KyFedwx+GfYwXAjpD7zDH5GIXS6OxJzgpvR9i5S5hEtRlNJ+6smK
nANbB7NPAq82Coku6A8I0qaRA+KX00T486gdWRcOk7R/fG+qVr/HIg5mftReXbwj
3faO3FQOzl69M/p1mlsMyeAG61cMRo0Vd1oB/FuBk15Mhz3eiZ4nixecr0uSe2Ay
7ZhB2ly0MPaIqhaC99i1hIPLpvBCQ01VCbFEFO6T3h6OCNusNMa4IUtov8rMvo1s
btn21o++K1lHH81gCyCLcSZCkdzJlXmfYWwzRdTHWU7itkvRde+3P+LJTm1RzKWF
+etKFTk4fjPOTVBd+CyLspcCaXPRUH1xk/jVhg/k2gTT6YxAlKE0f/I+xH4BqDQv
z9p+95SrPqzgpkCWBIA8t4FewGwOsgILmERl69Z4fmgCcUTtpRXRl3azZCOtzIgX
NmvNC4wUpatEtAeRJF+O/72pk1UD/JNQyZ/hKNQ8X6YSSjB8lvsMCqO0o3KW/dLe
n1QZDitMa4WUMqApA/semHRCs9Ea+Qa7edkH2kzYE287OKYV5hqYLZJiS4XtNUyK
WiesRjRiVl13w4RMjiDWTXbuiIoLV99bliMh7cTVCQE2KASB/ckj6RhKe2kscUo3
QlREUHYwLZSp6HGbIENyDlY56CR3lSxkHTfsODZRnqHpBs/YnkhU2R9v4SzIzqSL
UFHnvW9xx1I6jziIydBxjoB3mxdb9LtURxlljSegjY39OOiH0HtkbcN53vMReazR
Y8MrFqjTIxCNbLqfwBP6NuY5i9d6LWJt23+swfIQHED/oX34MUwSkZhv6l+q4GqW
ci+6lD3E2XIqJuNs8g/VbPGDIW9DnMC3aRAXjTGJW0dpXxHkZGU6Toh7Ry7vr4WG
bEw+S5jgoHHIGyZ8Kk3K/0E+9fZqxZDfbxIXe5oMCWJZZ1X0M0DTeiPpFVMGTfnr
0rwtoFv9jWsYi9m740Shs5Y07iiniYAD665LRq6Z12vakFXNMQg0q3FXbladneAx
pUC++Lz2DWIE7XbPw0X986VyiZS3JuNMVJTqw9FKo6ml/cEIpUPMpjX9G5oWBnDZ
0U5PdvbZAyqE6SQGNKV7GduPXQOpwT2aVelkwifXzU/PAJLkugTfmVpOLTEmP9D8
OR+D/VnCTz3+9/9Q+oACRc6e9nA3vEjcnfrHHshQoeE+nhD0ytE1FbOqCTMEIEYz
2c9xEeoortmSzk2i7aW7Y5awUVo5rwCFf/y3eRD29QxIVlpmY4FKxiQtMb1Il7wl
GQw5evBphs8FpSDsRtHPo9l8T4G7KrJrq/3iL1fHVGge/K8Xy6duErb7AZWsLzoY
mFBSQBefW0naCaGTCfOhC+rgidzCBXwm+QnwflFs5gbjC2RvK9t3w+dstXfFGPJm
uPic2oVELJtMlqjmyPwcKmth9kAY/ux4RqAUixPcazNwwe6/c+aBeEk498n+lz+V
u/ofgFduerKMf09S96cKblAA5twONvP0kNQJk+HV/1nqoU11hWitumWCvZCwbn8u
5q1Hwdst/1GXOvdTcDaEwVpG8pQ4P7xKKBlRSDB1v7KP9I6BFSV8fV1u2Bwue6tl
ahd0Vj/vN+7HmeGVX5p92Yo1BjQ+S1K4UZ1cdiv1EBTc3RhU5JvBlBQ/iJm7yH79
pZxTRIU3n9V1XnQ+V5tG1JTx3dLGr/MO8bd5IV8I5dcNgd13ceg6tMDyVP/zTFTb
6BohDQ8A2DIwMpsERg3q6ApDu0r20qx54Ncyg2MCl/DvtxVh3U63JEXYPpZFUsex
jfriBf4c7RkLQbtVBI3lyrOUtOAd21XC2sl21OhzWpdFmLAstYpPGxqdU1FTjNL3
HNdutV7fe7ER/4Br1w2F7kNWYX4gleo4cKAdVYtSF3mzYdbtmxLCOfc3uyACENGS
Qhv4fqLVeaYL+Ajk39MlRdtBGd3UQqlPoLDaW6uCApki7UhzPvxEQ/rYk8gBmoeC
E0qXIkkUr50RPciFKnoZjOS+1t3BXhA39++iYK7qEXlQ+eZdroBkwJNTYAlJ90OL
z8TR8GBt/wPOBeHjmeTK+VJIJigoA8q9VCV2Zrl/Fs9cyNW00Iqw0tq7OkDaVV5Y
1zIfAjrBf4/lyxNL2e3PBRCr54hvCbIrnB7ulnt54+eRQ/Hzgb/hsaldFn65KRo+
m2/c6Cd6Y5LQz5zySvabpjd/vexhmLtphvsK7VfMsxe8KliLuZbGVHyqM7cYKrWJ
fB6z4gPDYKnLQG1yOstUFXyK8GeRp0JyRO4kY+zcXZjXszp4GZ2y6X+nsrMxvdEM
GHmTYFFf4Rbe7CtC6QgwmsE5Hm31aBUmrAdxpJWA9ztnvDB8U2g/kagUIMuvbBcN
zcl53vHR9tUMUg91nCa4bVnVBb8l5PBRNxUkmfLlBeKJGtl2BviBIkjSzbPSmVRa
YVUCOtEejBQS781T0yl7GW/OdEDhpwzqd8BecfwqrNFFUpvAUeUWW4lTNgov3ptu
Mm+FGX0btBpfeTLzlNRJW6BTGtnCPekAMd2sL4uQQxjmo0b0H10VW4Jvm3pDJwgh
DMnuF45i3YP3oxYH48qsjFDdyLEjczLzgKstZkjp/gZJODtoG+8bh2lVbTdxetkd
ALad+bnOTAwA6Xd0fTGyP6vEiXytRDZKW8JEAUTw9i3f6gosMJM9+u0NUVun0Vos
iwg0l8SVnbDPdpNHBNYgf0Zf8E81Nmzu1XCoQI5YYbD+jdVlIuttxf65MinA/Lnp
F5vTfz1ics7zCdbdObXeeQhTF5wIgoDWM5uwMcs3wvN0YC6TC7qYDvLZtT/BEVzT
tEuHi+W+3URdyJdN0n/hhwGhZ6bUA2U4O9QWz3Abkvhraenb6aTsoSSgZQW2yomY
9LjvwYQrRyjLwvmM5M2m0i+eSBk64U/Yhs0BvX9RDRM0G0di933I2GLeZFEgmo5x
TojaNTRBx/eO4JI+IUQ7ljGY4Su4gk88x1a83/tMyV+WvtN7q2031WXtLzuMx6Wg
10ibVuSzucMj2Ws2vwYBZ27tO5etLhXSp/1emYTC3F84yH9AIQhMafqQ4wg/1LnV
NcbPw2gx/rCTaJulz9+cwRmxZw/Q5up/JlrN+J4fqoBK6/BWAWS30XzxkAXkW3qP
ccLRWQ6cDmRddxieYL5gOGyrGNI/i6ZlaO3IhSkuiTzC5o0vLKs+ulKgHRTOLSOV
+0YhYZKtgxoDAxDxvaUpxYhqd+UlCjS7wSkb7seM+A4S7nQq0lOlajT8edtZ4dcl
a8PSdJWLEYClLh1WeM3YV9BsglGQGp2MtbQAdcu/dsV6nLePDI9ereIBh7yc84r2
Fy9Yy+t22U750C8RzQLuDKm3OFPkb89dHHve8PAm2r59TiahzK/zyYIfudR12wJ0
q7ec9bIotm/EXifQp2RBWF4nsvtaNp68cKyAS1yaW5sEnjL3VpI93lWlIziNuPuU
8nASsQp+jOfK7RHdweb39VUYAluJyQjXNbc7DV4vcZOSmwTUPjjxMu1Bdja4dWQg
aZPTBA5MszEUpWhJmlS1+MGTQKWDkZA8yUdmOrzjRdnH8Ce6uWe6PHkmNdqKI7t8
sxwt88JkHC1YzaN9I1kVn+8hFXFq0nIWC2OFeYOLnEVtM28qjGicvX1wEZReK9U1
AOhDPNw6W5rW/QFCJ5NemEd9Ng2ZbFixpifn399X54mXUZEYpS7sekpG0Ix8EfC5
bkrVVjmm0TvPXRbcgcY2mgt8Tc1ND/Zt8NWKrvy9kTDpeT7lr1s06zKCqrh6j+aa
K99OB/r3nf+ETB/+XIVReMlPV04tPD7Vy8ec6nyKa3LaSp3E6g3nQcT5nNJC8iWl
0WGTgK34zwqThfAZYRoOKBtiCif9d4p3Vr41su0QDiMkaP9nBuXLYc6OJoKjU6IN
oxhmnJ03eH86mnfLWwb36wOnUNDF2Gd47hsD8Rwlt0HARZhjMKjCBJ/JvNsb2kHW
bFsIoYxOrL67/eBGrJ2OkpiCJ9hnGhhZsWgNVGcJ6Fsn8k+P8WOksMXwHxiwmXct
T4GkKSTHILg4mMSRLId2i+gpGW41AqIbIKFuNcpcOyh3AFljCKMmvT5TkZgSJj9V
tI//EHkXAVpuf05ztSAai0FkCyejDmmYhxj7rTZO45PaznLJQuz3c7CVpkr8l3g8
5+Fm3rFUzkjskY426lCrmWS9vJMoHV/koG8k+4doCAh4aSdhv3JDrSBiOFM8SRe+
TZ8bhJ5AB8CIIN2oE9dAMCrpkK7t0cAaoKDN5DR697IFaZDc09PI3An6AvuIR0Pi
RoDrOdWUXF5NbRJi/g5r4Tabp6WCHzvJCFhQb8kYxMwkZHr54AmA0at5DN3riKzv
ykNpizhGPj31+enJ7Vn05ZkYClNzAsoAdTpITOqquz2qDhZWeBiIfAMn9ns6kL3J
0qRRxeG7fcSNW9rnvslrX00MnT7OgCeR7/wLBbnPBCvQuE/OogAMeoLmdw2jHzY9
S5CXfVAAvBL1X6CH101BA+ziLEwAOkiYoitK2c6e91QIzMPtvakpBHSbaThTNnqF
FLCphgx2nCUx0/6psxzOXJXQBtzODhIJv7rNfEa5H2ycE+7d5SxtKdc1VOtPW0gL
cgvVqELEY8TPVHJlr5hAdKeHo3gd5OWufj4+eZX0sBU00CHZvmxBRsIzxKGHQTUD
63jkleDrlAd/Z/sQfvjZdOlLy8zcvN3/rxkJHGD8jplq50QVxjeL3wsIV5XWaGHt
FvBEHx8PrdfqaJu2jG++YWc1nr7hxbJEhNiraOiG2MM=
`protect END_PROTECTED
