`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zX5k7B+ycw4J43dqzgoozW0OnNjH6ophyYSfx8Pj3L5kqSkExfvH+1Md4GSOASxW
Mo3sc6U3Gi+EnlOmMxH1BHczSYwvEzS0GEVkWda+ZGf5p67S0rSWxMBj9JtyF0zl
WZo3b6mc487wYpORoyvgLXGMK+sMeimICnnMJCoQmOaW3gxvUUvmSyjSt4OcmLaz
GoKZ99WzTNCRqQes50B8TN0jOmLANLNYn2syT1EExI1kWzM3n1XccNe5ypa4bBMA
id/v1EV7s7NGpzEsEALf8ZZ2hoPKBgo3LiMDhiW7OngwHkcZLj1erahOj4N8ZGJM
btGLE/rKjUuCMZDmBtt0yAeMuR6CX+K96t4ZvZeHetbfgJ2gCvDg8nenjWrQNvbS
vmC8Ovr7mWpC6XGHzIvJStpzNGw2bO4g4LI3UGP0RwvYlc6JLsR7ugqSOujZatfs
TtkssAeZt37vXtQlFSZSjs3572il32qQsMjV6aq1ZOh4atgzvCf7FtiBlDXlzyCj
JQoiO8N1ffj/N+b2YKMWBSuRQ7OP7Zl3t4qJyy30h5aPv98NK5lwpY/1KJfrpSWB
BEgP2yuzkQNTRJxatDLAGyBOK/gsy7Mdr71NJBkO6f3pYC4BGQVRlGFKibJWMLB3
sI0fJMNQPnpbDkdRu3KOlzTVbgpKWRmct7c/RWarN7Tl8gOMJBWnwYoeeSecGPmv
7vPKgxwt+kVveOu4c5DWWzS0nfWJJLp/bD7uNgaDje5rLTNbrUXr/yvMpOBdJN2F
9KyAEpO7IKODPsnldak812+jwe+KxtuXql7y9FVcWZWjJIDKe1jBl9IIJa8R7Pfn
HHC4erA72sToBsyVLZ+aDutvak/JcEB7bDbu5uDUNscT9EppgGpesfJP0xcktZua
SbAyO7ARtro7ky2QhqzW6DoLP4yg04hZ6j7G/f7OJ0vqY/MWH9SDYtlpkTLUbKJx
WV7LZ1MAC2HH9WnqXimdc2ALR7SP03sj69xPZIjWpdhLI2anw1uLR3hsTg61rOu1
nfZ87CInYnyQP42vuvpmvsU0MfxpbjnwY09MTZrxzslXH3ZzEh1YYHcJx6nwsHk4
rqP9T7EWKMGuu7RytmBSddqh9UvusABvw/S/yNsaZIgJjQHZ9Xkv2PEGU0UZzMEI
ftr/LFTv6Z3pDmeFpms2DyA17HxOPCnlmT+4bfcU7IybON8hDMTDMjIsL/LD2jNS
l2ZxZCQIxcXFGI7VBkdi5nx5H51u18OD7GUgsSU17XwJl4Vlxx7YEMDIMNQwY8uR
wB/J8lKmMqyg8e79jrvHyX3TPB2OBeFTze+qvNab25PPswEVMlfMbtgHQMwQMmL9
A0LQem3apad2YGO8XV6SjRlzWpg8BkTWvbKWFFQZFtbiwquaVrtg0m/ex/o4PTyG
T09C9zZQ2iNgldOrwNrkxBjywi7I3zbH+MA1MvXVrDaUOQL7FfQUmfoz4Sif1Ja+
cMMNFw5wwQ+okY9o+s1jNbr+kZdhSqMcSj1o3vbkCI/9tg678vCrjbpBAdzTGZkb
Xp9wWsXrXC38HWaP0i+Gdw==
`protect END_PROTECTED
