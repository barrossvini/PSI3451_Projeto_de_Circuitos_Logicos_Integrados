`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LiB3FqI9A0k0i70CKb/uMUTHYTPfbK3lhM8U5CDAFJKzBTDwS4qcsZzWTTfcodwx
fl6lKyMDBFUpILj2CvhxCYLlcacyxdTc5ATsZwW59HYkhy70xq+quE4k8SDQGVQ5
nnyANduu4xOwe92gCZScI3L/ybRZzZb1bR+4D0bMP79NicryD9Z6vU30K3Uluevz
eLSd6V9JlbU59T2CApSpaiWpsQsmQjaLKSsyW67+7nSMeKCaacjavfms9JIJ3KKs
eOtnsQFvzggamvpd1NB9XOTOo2bvCo8fVr0cy6ZXyAFN7wJ7VXaVUPCA2cShJKCn
vMoY+D5n7putiK6EhG6CgDRA2sg0NcjJzg/K2wZPUv5Zx5eWoOTmsT7uzeUoolT/
ymDfOHsALCnNvRCeuzgoUdRsDRk3ub2lv2iLYoquHXUR7RKYrRLxZw/E/CV4fJDN
MRozLBGLulhQPH0h5fnT+naNTxrqVGCAcm3Ua3jGw1oNrBqJ24rwqWKcJdT1wpmc
mezxX6uYRHdLu00pEqAJ1I4yjYtdBFfy3JYo0fIVpJ3XfL5nBVP0ZMNlPrm3zhno
yiqClcNub8g/ReeJFHe1JP+10ONvU26cCwZakJojCv0J3im9BuTtPSUH0ASMu/r0
n9wJN6uCKDFZX6cmujqOdlVmKPAOsTcPJpImyh9jqGqsGGeJQk9NszVJYs6PCB9s
9DWdMvG/2Krd38XXxuIklDiF+hzqDXO4lk9BDdur7WTnsL91Qt9UwglHd8yDb7bP
zc4zt2w5feq+KtrEo4ucrFUqMrGB/u9R1NoUXOL+xrFz+Tp7glOt5jb/zhXixv4c
XM3kGXV7nNiyTaWbqOsQYmL6e8q2iFYPX3T51dzNNvTne246pcjFmiWwmFOfd+7J
fydm1C4EgRz0qxd/wZ8MDoASZfWSpP3sKJ3h49OLOeLRZ7YpOLe5bY0cdkhvhtp3
LACiAjFsuvcA7V+wrFE5qi0lTlnvRoSqCzOOeb/uiLZCCjSAcRubv0KFT8ygC5KU
OURLNjisMSSkSGiUi9jJsGge5/jBEVyhmhRejDqrZ5jNFmzNZx1uWxMcCChuSFNE
eg2T6GhuS+h7JSVdZ3/WEkWJ/wvpUxZyW9ph0j8C0NfzsstAdkdkXPANLWSnbfRR
LHVz9dKMYpXA+GqIQPTJase5qlOFPoNzxRlT8+FhFAbh28LJneGxDOdLfRbezwCU
x2QyEzgN3YmjYwCRMdpPgf2Xa+sPOTjLLdZTbNygbbTHkB06rsinKgXZBoUD94Mr
2ygw3+zKgYdEzhzzWRCqVvSdmwUzgVSW9CxZ3GDdLUB3Pyc+tIDdbk/i5MwAadVG
cvD9QN+9xedsOliehsqXIR1hfO3nmSRGtmMqUmDfZpiaESrPmIn2SKLqz8r0Zfk7
MSABPyn0NhVIcm044LIywDnKf7D0EmZ0IvwTdXCw1pfH6jfq7WgeM23YTPZWGKmF
b+kvTkU7JLponjwsCzHqFBBEbSOkR/KdyzfQP6+/BQV3G4XRPR2CZHnRnd2MjOXC
DYgegN+xSQdlKERBP1Cg1QtQOUdZN1qgq+t/hR9OhQSq+EIxgmCsSQ5nTnXTJIV6
88uiadNP/U0EngbDCvyktsM/aynXEe+gxzaN4vxk+CJe08riyo9kg/XVVErANQ9f
H3ylvMxWTGnP6hFlcll+WIS4HvgCYWt0v3mcysD7PEYzsGZFkt1w9SsMKk1Xro8H
8TxfWSCQoQJWmkG75eNlid3QdOUZ12b3JlJO9KM9M+qDSTRSxBpy/4U9U2mc7A0i
RxEYOB7c2tK5DvOdP0YDDrUJ9iC7n/l5BtTwyH9CnwBOF2DI79UBAY9dYyYMlGkE
mseqDGz18A3ZMAu0gWfvZFITY4mMMkKxiRziG75Gv8DP/bpRprI06exuzskSzXb4
ZPsmn/ToFlBA2+ofCNgMH2sdhSuF3dmi86Cj7EIGK/okXYF1D9Y/ZRKzokjSQpcj
+iEsuFrHPlyq1KyLJwoqp2riKuP94rvlvqvPRJVH8FMIfSnCmvo8FTHCnjljmNSJ
Hdya5jvZ7fea5Sz/OEedC0rzPC6uHOBsk9t9+2Rkxci9DR42TyrtGujLyGLMU32d
hzBijAFZr70d6x0GyZve5HH34bgW187w1WC/G8CLvIVyeX3/T9xjIytUDkVa1NnT
Klx36WjcpAPp7mZpiYBoXhosR6SkCX5u7GzpIdLbnpdf8WPsjV0cjkHfjTlZujfe
X134L5E7i7y4fMPt+iJR0sH6VKDKd00n08g0GZtHnxtWOTi3XRrjCPC8PE7v+wGO
zwr40AGI3aNLN7sJsxB5RbFmpqoaH1BtwjrCif+6+7asfZrMpmhErsyhKaHlhC1F
OPy0tYOYlC8uaWZzYMKGvM2tO4fATPtqHq3hsL/OJufvUiggH/XwSG12IZui51/g
9x4tJ48T6/VHu/W52Vz8rR0lBxrcsT/HOK2b0vh8fdxBMjYfF2lLNbFTFp/M9g0r
9zB11Gcf0zFj1QLjhogZxlvS2INNVwAyR9ET2Ta1ozFbAFdefvJ1Xx0BWMXEHnWa
K0TSlQoCEHYTbb/L5tm7IN8gwD4Wf3WgfVhFzzplkzqcB9ysX6lcEm/kA2kCZYYH
Cw/L49jS9fSFy9bPRUqgWqy/gKL8vEMI22hzDL7Xe1aLabIS/yo1GNK8Sp6gI5ae
/HiFsS6gJrXSSu+udbJ44lcUbxB5wLrJvf19uE8BVfoksK2nzaMxqR36a01RQP4a
OcZCKZKmU5H3q3dBR1yZmwfE0Pv70s7SCV7vjWjkM7fm0iXWQaciRdqINKd7+D9Z
1tNq25NKleScJL6yIaTzvphPea6hLkPkkNLxBXz9l5Pxg6vf7AntKD7QR91Ul97Z
86MJ3OuNjMsazLl+higiHbwAwT3f31LhVPX4Gcky4nBGjU9R4g/bkCIQYoUhQ4vE
NkxoLZey2fgl03yrJYxKOO9ZInq1DCj2/zv8oN5vaoKaNS4dViMgAAUIMHlEYCB8
VKc9wwUZ02fZaNEKjIDDCxwaFHq9k2zGTSHBATvT+6eWsJLdsMwhr9XenfX79+m/
sBs1JxTqnFXfhFdZXEG8LP9zyVXi2AOHoTJnHj4Z9zq8RwZX0IJYuQkZ+dbGUaqU
UkDSXNGWGbmVkRpaJ2fGEmcxMrd0MH4w5lfwzG4TNP6ljHZ0nRd7LTHxCpUiI5Hy
IH16hjPvcLLrtlO6RV5Xc0wcQ0qL/npkwCb1upV+4Y55UR+JOpilzH3F3JyxgaHs
QSGYzo4sPMaJrvI8KQy4MJJ7JMlYYg+NthGMhHqK10ZSx24rEy7Dt5XS8oytmPhR
GDXRDDk9EAUb8pYHtQs6gJV5ELQNvw8D1I9VArjJ2m+FV4OwQbj3YdpCMze9hLcC
UX0B9pIvQ+3NxyLmWiSEkKVeS15tFgf26jdCKnGYdSWD3OFaXyjpxp4XT5OU0YA9
2mkDSuktqlWJk8SCztGBsnCinOOS1GTlEIJytJYsbrFNbcSURSQK0N22JYnV/IsZ
BwNVcIPMrp6tOoSHsaz7ev7CLE52/mH7jbBTWwGFOIlhA809AuRM5wMWZzhhY87+
B2ut8wK82A1oIHem7qE4DIOuf8+lnzhBMkbny8QgXFwXikFCPmDZiVNIMN3lS17h
LMUnkFM2z4RuHO4DtsI9o80Nr0Qb25S1nAY/NyJ3aupgiBLUaMhm44TX1h44r/RK
9tvm99u0vDkqzvpf0eHsgWPpwszpX2Ti9MpkAeQXV652PXpk59x89YntYEB3v5T5
Yq3wpvrnVZlRZg2SOVhrlXm+GIJ78J5yMm/T6gj7Par+D87z8C/YrphHNxVuESgd
w/+7PeaVBJ/cFTQr/mNV1ggw1iDAOJp4hSQyAsGQDcXSuCl4/qmTSCY/H4ZZuf5c
XebJOWuz1vqPrnCff7adHYE97CD7+LX8AxVXu7I4T431rcTVWQ657K4NtxxEzyHF
aR1taiC9uIjRa2/E9ZKcvg559O2esEoH/JDsb+97pPJV52BW3YNUlZ6XKJ5jiaem
cPwJfwGZaSfwOX2KEZkHmsgnhMF/XKRKdCMpqBIa/GLQEs3eVhIY7PrpBfnE5GnW
bOS+a3IDOuAFF2hMAlnhPO4GGaYo99o1zbQTppUWK40wvC5aSm6DBgeH3bnEMz4y
4baJZdDFRNX4pm/kPP/pHANUpOHg9k4LY6yaNaPcfKN9clWzQeYMTDpzE/A2CNbX
TvSN6qlYdKlBDiDL5vPHg2HqMK6Wwom2GNi+fjumBJNx/ik4lRY8AP/JZY64ZNet
yby6gPo4b3HP22JNimPldEIFf+8hcEWJQ6iKN8FLoR0cHSUIiNRWbB21soe/DO4e
unOo4K+B1yOdOmGMmMZHQdiD81bJmJt+9Hh/jKsecg0VZ9glaMnsYxzM04H/7atP
2Q6J5b72cRwgPj1K2Gte0GmCfHMAOo8DHWBWPncCjCQJ/19Q1xx1QxQsSAgUsizz
l8TOe7TbK9XIbjStN3lV9i+t1kPVboXdQalns+2JKeHBO+jdgZ93Yv/rHnGqeK+8
gjCln/l3IUGsES/WMv6q7eE6QNMZk31eKqc8HkCUBl/VyOxfO2kEcaBZ9w29Xsi9
xWCMWJ/qRv2bh6BLuTEsJAlFJkREARZ/fM0IPwKOVBT/1K3PJJOpuSRQGe9QJFqk
JMLNV7IO6D0btDMI1YtmTaj9nmUI/nJMk7M+H4NbN0Vojc9K4cJhGISYTcjuOHRY
8uBRWCUEszbU8UfxT9sAE82NDbC3BbBKnnv5vy0bBJ+IiJEpjWwI1imkMhStBF0T
2KhAjOeCuSIdEzcMdAMQwtpU19l5jls6S/qagenE60eIyTG/s32lyWThqv3ZPhUZ
F4reaFp+dUWKz02zpXU9x1vBOhdWNyw1cherh6FV0SOQSHKmGW/TJqkFFJ4agdwg
qX6e/pV9c3gaRad6wLyVu0c9851QQi1Y7HVYV4jYWxSEG6IHFWpVKDi1+wQLtd4q
tT8NE8Y7nmoRj8Wos3D+CKLca1mm2aFkEF6iTrMEGj9Iwwq2+PKixP2dCOEOYi91
LFVGw7qzKQQBl/rF5xtvASE3QOu4y3dT65HVtEM3j+lTnq4K6iESX4lSE2H5vOyF
ja4m33C/OEco8rKcYm0DJY/9j8g31OrqWm78o57k86NpUVUbe1oLjx8hxAsWTLsj
9fm5akEhPW1dqgUqknNgeqNOhuzPt9tGX/pN9XJWdRoR5Dw/ZmzukDSZKaOUZyCM
uH4FEFIVB478Ze6LGthk6DGG/4FhPj9j915eRdGQb6ZGhoX+13GOV0VYiBbQcly3
2ssBblZmRPKYj9Ydwkcw64RwhIlfyA9WN3tBF1iOelrbiWD7eequb6b5Adx2FXoU
BWN7OC1vzMRotbfyZLVXz9rCdPUL6c5Pol4+5DiU9tBBXGZOd1I+tSx0ExZc7nSl
bTOWyyxWwi9dPJfjEGiGHtQ34QpYLu44pYLleGegQ77I/UP4vJUeey81tP/C5iCq
2sj2QlXK295Q44c9wxp9z0E88HvGEBAbQ+W+fdpsK9a2SITRwPvcUdP+dmD7Xb6J
mg1UC+LyuZM3lCdBOeXJj/IPbtnDTBJgp1Qf1DqpUe/0oepK+mRTRWhX6FJf2Ry3
RsaL4VFYUiynkRuco/hYmrTajSqhluVp/4somWowuyuksUuX6XXSZnZ5Drx9Krzw
8+ebXDescTkNJhAeb19wiwl0i+2hz7JVBA5xB49rxCtKjbkcSphwaF+i1dT6rnNG
T3V7YM5Xe6KEXHDaF3VjPjz6irwsSmCM6PrIK0kBg782jDQJ4X+K5M5f4nUaO6Bb
GTFExzpC9RN3VUbXyzrGsMnb8BnKqTI7nTfeHTmMlf4obg8rS9nzLgSIIxi7CYR3
a0SfW+zQYNk4h0pqsGjUa7h1XUxUzBRFJg7A6ANL7o6zoSMxuXS900p3Ydka5VHH
gEN1VbXTtvmXWMr0mfZI8JFkoUZvlu2qNV2wyxLuFVBWdlisnwwEtBSOzpPu/OIV
ceExUKlYKhvP96JLHJTGJCnS89vdqUhj9kf2NSaodbQQTUQBCINg2imPY/XKwUQc
OHnz83tuv5x7ioEM+qlA7ukTe/AZXzTSKTPy7ShuWORXQgm+qMPop6QCaQ5jjR4g
5E3suxGLHGY8R+pqQWAyl1OJyuPtlNmi/1j+eI4dHrZlaK4w0k1ayAtAzBFKHbHD
PMF+P2f+JeDIjyWA/L+bAIQo/T9HJe6Wv4oewtdiFWgwdHyFuSM1t/qlcrdPRgOQ
j9z/Xiqwav/a66lZWCy/8hJm/5YucpZgC7VLrI9+vjPavyhJhR8E4cXJ2irLLdZx
ygtfuoVDsqbvUvHbLw1fI8DEqcFAaCgsnGoTXFty+T1NY5T64S3dxHd6+E7U7nLQ
LUONJAhGeAPJAmN3rZm2P8+oPQubcNNFE84M97EMeB/A+PD8jyY5ESEyt+Nr8Py5
/VK94I7TTV0D4ZUkF+YUvmp/3zec7ifqQ1MbRkguLnpgdLODbOB3HZs4ez8p2/Fj
BbcyMZ41JH38QzkolsWfwGlUP7PrsiVVcUWl/FMmuL1OuRzPMG8Zyr+muLZboZZV
RYzeYtCTeMpeQUa2XyGzZHKnOrYJ0m1APYnmHSmE3W+lHJeUWas2CySRgmMWS0SV
C49tFgM4wpt0RMaOlA6L06sqWfoFTHwgJAtuXtRnFBwTljL0n4NQwjo7Z5rz1fmG
QVsnKZsH1copE4IzotDCRhXuYrwAlJa2kqugXLKMcJyKn+1XX3pDy9QXn6U+43ab
/kOYs7em3go2fHZHatWWhfjKuzjooFEcumYysKso1HZmCdH7XRW3nSJEPsv+zfGI
WVjro1IkPxU6GoXr/4+BR6jqJo2ZFrrCIaKJVde3T4h86cZAd4aRf9YIIfJk7QzI
6FZe5Nc9XRrp+ln4J7GhcN7CbWyOU60jUQLK571RfGQr7QjA33PAHOn9ztbzgo+W
BAUgAbZBtWuPnjdwYxtOwxj6pY0n/OVGxeHypC8qDZjf3VkgX7WhxnhnUPQiezf+
1eYqMHL7EshTLOYQofuUYeTdISHNdxhHgJll95shRgbm9u3NqAy6qrSXmCo5JXBe
JtBxAN9fr14l6XTU+uexNLzOX/oMcRUBbgTsWbaCH4EU8E/P5lZ6QJNMUX9THzPm
8neC3TDTbuhzyzQaMimGe+IFoKS7AUvsBpMDUNjT4pZd3CdyF5REOX8AUqiLs2dL
Rw9rZyvfxS3hYRgt0KCyoMSe9S0RDPRZhv97WmJ0eOA=
`protect END_PROTECTED
