`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
djFegSuvYe9TVfq8nZixt2TW+0k4pmK3AYFpgwYHpEPAz5nQSlLtNm1Td9mt4ur4
lP5MJrO0U/2ekb/EZJM+G30Ojy53BSe3H2ktVUopWZ2N7J/pvEp+XTq9fP4CNwLd
yfYGfe0iUpz7i6yPgk0Az/KsRZXEGBuG/HrXQ8EWLFrLtPeq0gCthzU10tAjdQ4b
N3EOrndegQFx3TgSHrZO6kjlBiHTMZecduETjotm1RrPW5o4EUoErEHcs4PMC8LB
EpX2hOX2YlBO/8YPrLjDkX3K6Z5rOzWEIbiFI5b29wiX5eW/ts2DCuUCewqd4Qrt
AsfzxBYvGYiSlfyH1EUaSzMSWPRs6QlhQOSTymQe1Gn1eH721b9CAAKEG7VOsEEN
0Qfv4K8Sl9RVw0Z5EZpwf5v3qZepRaX6vuuSSlfRrWnNTxvMn8AELzDfjeFFj4aR
cEexcHMyZbjn1fRcF5wkcI+ZOeNsprSwKhEUtQssveALN/euODNrYNRniUt2ij4A
7DVBHiQX4I4DkPtIz4CxJd5BBbxCr5d4xF0vYPLMhtPK9Ed/hVAWg8BKjUtnNqSl
X/SJ55VdDMTkkitXCr2RJwU9/4h811R60y20nd7zzoykCh5QiWxYae9uhbMq+pRv
f7ZadFo2U3pwN4ITN1MQbEZlr3mmfkNfy5yZGsly+Q6LWVzpyUKRzxol2LDf0ReZ
V2GadYpVgJ7qCgEkQbe45L/bwYO4+uCoYKdpODBoIKBZRaDZkbf5NbdHx1CYBAws
uiNwedYj7wBhmSZVdyUjWg==
`protect END_PROTECTED
