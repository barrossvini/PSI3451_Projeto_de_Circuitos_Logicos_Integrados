`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Jf+/gyNeIt0ZY8LVej0gkLgtL0ftHFxX8XkoW/Aw60gpidt9kInjqKhQST+Wt9g
8FNO1hMt+20bqsxVLITcEVgyoQPLihPNvkzdvvbAZzGlYoo/8nUDXp99LBEO8+/d
fuLAIRrrkee0500x4OzMks5jUZFdotfFWtg05BcQtEDWWm2jxMk0B2dg4/0IdLUe
vx9e57jk+AbDenO95CV0VTsUGoTdcGZQ5CtLwqObzsXR+EuzJMymNA9xQuMkpZD7
J4KH7jdcdhtjRN/HV9TdIVhIs9I6EQA5UhYyOzkfL6mfENVzlAPgwVJQP3vBO3Bj
7ER9Bzc7Sl+0FdEA3ClXhHlErCiIeg6Y5HVH1xuQHhdyUb0rQqHHxMNfmFyTZBkf
YW7gEf+7o5sl8ZAxENQkWbgd7wzBnOQ1ABk+8R7m47tkavqJ3Mpu11xahU8EkS76
pSmxSIXtqnC71MV59WbGJvW9QA9iqLfKzxKi+3xZjx/WX3UfSs7R4jTuuKvG/rEf
Gqn+f/B+2iDeHiCMP7U0FTOVOUC88lt0APoO+4Yx5MlMy1lZ7Clv+a370hXaISCX
UYxr2wSjrTz9byifOKJnm3Ystlcp/7UFdM4trRwejAhOXQ8TcAZjMLhFE9agsk+x
yhMgpitJf1qk9SlwC5IjnyQrTy+JeW7+JBQjYFB99JNznQhmu85dQRCqo1UI5iFP
DWppN0dln33Jayx3IJ0he/sUaugP5UZqDNbUUTPb/2TcD36gzlIswFqOoi+a1dMy
p/QFQVq3/3c80YEelIVJPyIqgHuGAv0EIQkHSW76aGxAuhjF37FsF4MCOFyWekkM
DlEv3LezWcEkaG67UOR/XsjLTTqJtOaVfAFgTndyXCw//RfzAntVyDTssaC6LRxP
dXZu2hn2nq5Y5RHtA5dBICZph+bNV4NgxarF7nqXAJiKQ1IxoAnb8khOkpIuBx46
4a/0HWSrun8xEgaRQb1K4jYDF/jbdhUleaSHm3KyTmzQGqEGFUnHPeDlEBlGcil6
uQ+ZBLTvi76ZUpb5KkqWvJ6vQQuGP0DkPMdUzBAJZqWrXm459IGopfFiCjbgIaNv
UCPaVxd6QuN+CHrpmOagL2fo8C7G1pt9l9uLM2Oe96Tu4TLrm9Vc2bsbfVEYL1eQ
0V6pENsTdQEkhQHkGZMk6G4mVVd8dEb6g4oks6oMflAcd2gZnBGjCjmrykcSumrz
EOpZ76rhgPcRhjiopEMqGJHhGEhm8+ZpjKdjMWJ5T8aNRD/KbXMtriooHWFLA8Me
3P/sa4wfnzZd+p4ghQq6o/01FNsd7fxFmtZ9XoJVBOfo6WpjT/7KpybdtgyM8tEd
L1wT9kWDKioeGWds7IkKMBZ0Cj3ychv9ElYBxJwKOSOetJvdRu5u6UOJ7CECde23
R84ueZPxHfjWL75M1t+e4wMmRX0B4TA4s2QC+s/0oyJeR89iXkdPrIcd6VHkjD2n
ULJDwgeLSM3AftrDAbxhC4v2v70GB8Uc+IGph8oRZGG5HOr65dgwxlDDZtvth3ae
1gK5ZGf7pFZ8jQ3xUgJaqzFvXtrqQyw6TLWelGmRu5FNS/IfnyqCzAYA0VUUYO7B
J/Z6RYwSljCqrhaWPcMdmb9nipB4DNPya2496aQ6sd7pC7D6tk+V7qpzn4Vuw8JL
rglggRH2LZbWZqR7/pnqkqlff1ao7Q8I+BUxG9iQt6jTdPYTiHuAq1IFQaKTf0ia
MO8SnkVgwhbfqEFh2yACsHLkiw2IhGu5HPV4fJmFt5T/a9xMZzlHmtf71O3DXSbE
oX6hiMsAYKg4yWwCfsv2IdSrPlXWGowr4MIMvQrXEjhQQEPIuVu299S4zFWZOzG9
8WUKo98ocaevlC4MDI0TNsv1cEd5OYlquoDIE3l+5kEFDf63vt3eBV71coP7Leod
2h4NPyMkvJRj5o1ogUpYYS0zmkIaII5G7d++VsdmgFGQK6oFkuH+hr3Pw4+/VrRc
XZzv8MKbx3JURJg6mNg6VCAQH09BiKkADeFiE/y2WaLdsk8pDrQlQ/LDFcO3B2/e
bCKmEIxgQF88mxDuqDyRal3aGePzw9kuAmdNTCBOeZD8yijljOiTVrAxf7a1j3gM
YPdGaLMCiptfnysU+dwq1fteIt/go+ikkbE/nCb+0UKBz4JPiRU09O55N0p9St6U
MIjyZqxQ1lzwdTrdQqftTzhURGCpXM7iKjH+uH/ppJsLtbABYsUrh1yRW9Cx0Le7
eZOhimaaPjhnIg0Cha9vdA==
`protect END_PROTECTED
