`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DI7/C+4VzyYMB697Xt1aCYHQkWlz1mBp20pZi3DEF/0uApo+ebJDu73S0bsboR2t
1CNNV7liqoi92Yziozn8JjaigIrIW5kIW57+ud92sM6gPifrPpIF96l1qxzGIXj1
Lul5TVpo3zXSwCa7fbqseskraeeStHSq1gvyTdpHCeheTHd/W3UH3WrYCRDUTMJ4
TIUqpR98MwmQ0nhsJvVWj1m4lgWCScWUipK7lfo+M0phKOFl0cQpx3kF7V2VR7eU
xFge3L2sfsm9XMjFqBmiKQf13Fgx5CHqGAu4cpDkSU3VIfaJpncqBfthyzK4WqFe
vcYllvwMpqxHX/jTg8M84JXeypd+fKfgvouIURkDB9CYDBTZ4Q1L4ImHC5Oynr79
K2Idbe3cakyb4p7QQAtNW9oU+9hVJjUl6C0clM2+XfQO7C5hn2NRDbZH76POynHs
YicKjO4UPcrp6Zb/LluFRNYi3/rPlgTwXcpsZEOPjtTiR10BdfjA/8EpmPgTBKRs
aEXsTuewgpa9uj2iy68lN7Y3N8HG2BevtPA6d2SDZ0ckAPYwCBOJ0sq7ZGiWlHct
BhXWcZTV4hBNypYCpGAtbhtLjeK9pmAKqj6l1/9n0hVXFy+tfMw35nKl5n556Gxq
c16aJCcCjFSSleZL/yvvPITlTE1CoE2LuXJGrN9/xBabbckBBsn8FqxZhFVY2Xs9
IVsVFEbcmnPY1vMWtAyEf6aVNnP5HqccFqGyiTsYS0lFvPszL1AnXYi4mAUq7b3Y
KvYE9g/aR9WaJVYXOmgmvsk9yn2oDCLXBruL3iweYEYvFD+4Vs0oej0NbOPIYulh
94TXJh+/CgtLwhFpfctTLpL+gGf2PMBxUiLL4c+2IIAJIcjSBRdIqzalrkkyZVmn
dAqwMMi8ju3/aQKIImNTnKRr7EYKFoEBIoz6r41ZvNGwEiTq9k46a7ZrXwUqCbAh
6/AJXC3n4XZIRxI718GktPJHEWML7xfvGXv0bv+X5RjXelCEqYJR8SVEyl8C9eIf
+n1Gl+Yer3bREu6Vl0Ae5Q9wDOWP6Bhq3znGlGYidgbClthxfgKz0i3QDxoQluXq
+TbamSF2zOmG+BESz0T+2P2B4OuWiV2W5NWcsPZpI14egv7eihTU1rVK3cLBfitt
EudWNx0PS2BHS93ocCf3VznTq/Lmsab9u4I4HMLYEqvrwdTiTVB5jXBchFNZ+pt1
C4rBjlPMTpA22MmkHNlXDPfgIeQu4/8kj0/GD1nfCFgaUq+OEXfvUVoR6Sz4kPlT
SoyN2dhTHgqTibAqFY7WUXCRwCq+N6gdfCp4zM7hzKd4aycToMmzOrrjfXnLnSLq
eXs6GyT86XQZl2bnRathxQ7ue7UptWo7sraU7d7ZPkj1Nr1+HO8O6TzZQ/phSdlU
I+5VvkCHjT6y0/yy5WOGJ8RoclePPVtdMhCrBRYfnCau0ulV4umQ6LyPGR7dTC68
YX3eBVUkHaUjfokcyz+8Hzo22d+N+1UzPtv8A2iB3ubS9viipi52KY0ByhYIg8hH
bY4SIgTlTZaAU3EVtCX2Qis9pUdSzSuUY6JOd2e9uhO4MQ4E5zJrr/Gm0c6ov1eK
PaSqCwOUmRaAV1tlaAK5s2/oK2fZs1M+rMV4uMEkgOe0RnjNKtrjsPHvSWGChq/7
IVTb8rPlkqsP1UYhpxfdt6x7+25AYeD4zsu24Vp8uA727zXGB+O7HdlVdJw8o5IC
VO9nqRTLcp/j36EhKJiThqPW6KIJPbyFmvbIam0cgx31+RzXdW2y1f7Mnb6jyBn5
BjvHGpIAPOMSaV+3IZ+KT8kYEMMw0NCbHbzBFrXsz/HQxBRht1s+22GcWCqPr3g2
G3QMAAW79xFzoQJq+YSO3YV2lkIohNzuT3VSW0HXqaFJ4FRQ0r1CfvSfhnI87Vhk
QBYMJRFwirbb1iVEcgwCUKwnbxP8T5mTx4DPoO4blvY0Jc8pCoDS6TE2CP/lJP/X
XgyRD6wgs85df4XU1Od0+MlqlPLnLeBU5x8MIgG0/RlCCmXThwxOMqTbmLk/ky1C
mCs3U9Tp3aj77u+pKmKz9jv4UIX8AD0TxcqBfGs8OxLNHcITjkaE/cxrwlBfoJmu
dHzIxXbUqf5x2nfs+agK4cEJl00Knr5WSXDzWMPepbVLLi6mcZsrWWxHF6gYP1bf
KPv4n83N15jWCUSuCCfCOypXioNKNoFLMF2P50QrCXNds4dkYKoq+baTyMDjyL4H
+QHFDTR2AAEo1lLui8q0DGD1soJM3OKXM6YiHzrP7IaCVwmrlSvZXAZxOs2NARkR
RHKQf7/g4SYsYbn7Yl+mhEzM5OhnfR+8OcfaF+2RQoyXw/tj71iVPRMKn2UQ0cTd
e2Mh64huP9bj6kCpRZbrdmVyhaX2Ou9zP1rk3lRbKBLZKzxKcKUiFnr+LHsd/D/J
b173SmwZQI23VbMGsb7HU2PiejoF6D/81N2VpYD6cS1cq6TjrH8fNdkOE5WgdRHL
PvbJxEiI5rsMMIecywf3DVcu455Kcqm/wX+TU83XkGlm3QYW6SDR8EFQlG28SIr3
r4ZGTkVCruh4+ne2Rqkk/W+0F9wBEyE8Xbo5im2NhGHap5wY9h5zxFuZ6zzeKzuS
Oio6KheM78xxPMexwSsNk+OpdnUQ7kSlWxMrJZDICVJYWBbvB/C8WXYOGE1XQMFQ
NiUb3eubUTc27MX0Djou8IXYFYGr4ia8NI7VCfCLXEe9a/xyp9t7AZOOj7LZ+k72
XkmcapkjV8T+4CaoKqCln8X7rOTScnC7fTM37hs+0B/04FIS98JZkYoW2Dq5U/lB
0EBc2XmJK4Iw6x5KrxhInsTDQPxO27v72JLw005xVJ5NrHzz7HRu6dHMx3EF4efJ
i2HAdvyacW8H79n9HGvLhDtk9oPuaezyLz7KY7H6ewbnnWy1Yo2bKqxubQX1Nfbd
vsKk+ztO05YGe5rfaQweCYhiRNohM7ewG0/GrXQ5hf0UNCR+K8vYZvvbSVOQ0m3X
dmFPLPJu6PSWZCk+VDwlEPtmcXoisepIm2wdvhNpVJTVMzrgkwy3Vs37Cu3zrAj0
xzkL4KsAsxzge5lWicjmE901Ie9km5gZhI7qcQ2E5+tPbwRD3NcVrTvYjgbGfAyF
5w9Rks3qXUc7FE0Z61ESuS2z6G11OF5l+obefwjMNLEfPvQduBM1dwekJ+V5tGuh
p1ow9lcnqaowSJsV+kPdhtupiasrvCrTwA5gt9PdiSEfftjH0BsGFG4qorEHAh8h
15EKQactHdNw3NKi8SU53mWBnLpuZd5pyyYkTcnkXnqQ7SytPHQ2ZWsqZq/hc3wa
hZ04xMlMvog2BXUZoAQnk6XUkBwS1D4mtxPvMzQ0McFtjno0n7ohaCpZ/gBqhrFp
bd5MKsE0qsXZLm8psi0xoJzReobgo2AUIdjFSGU6gxXq/KqXbVpP1PP0TchzYftw
7kSNUqXnEhTzthmyK0cFPmR5ONq85acqrS8TOFMwjRGZ5cTRyZKf15mVVLB/jrTB
yUIYewMtgBlRUSaYyuMOhXBGB0ixb3lSKWRzlOv4rElU3vSxH5iU6HyGVdek3hOD
fhniQB6tpFtRdNBXjtektp3Pa0ASc7Hy3S7WwArUZe8HP274MUYnxDKFUmBhLl3i
YhKyGobwML2BFye/dySXYg75joodswObAZAeimYBoyqNqHmFhsQN1ws1LBcntAnz
U1XTLdkqZZIlJPCWSYPdybK+4lnDVpURa48sLXhY9kykG/kIzOUt7ygrkS9cIm8w
XsfnBc0+Y0PY/3QDDV9lTklWQ0le8ylDFphHWZDQv4RdZvs+BG4h/2GY/vQCVxy9
sQnQQxMO8thRC+dwmov8m6YSsySe8Ph5ZkbB20mn5BJOSbdBWHF+HKADS6YT0fXN
hI1XgQoOyiMhbCGinZn5RskrOTPerrhwmjf4/gOtJzKZYacZyd1PzSy13cPkmQ5e
MuNNSC6r8rNXSiWG5ga/t1r/OOEHyupuV+/fn88co5VCEDy02g67mbmD5nfixCQe
oNHxAo8XTY4Q6wo8vPL0H79ZYvrsXO6mdpghZXH1sLukSHT538/SytfNjPSpsuYD
kQdqJoG6mOcmYeQpNxc0V5hLxw3SFtM2T4q6fXZQNHDRtP+aPZzVFg2aZflkA9hQ
bJQ0iBPhZaW9i4CHsiEANgeR30OBARUsRsM7fkcr9Z5y/w5Qb5rbEFgloloNmVSO
afsFgWOK94P+XtUX7kAqSoYoGXKlAUKMzkfHaJANt49XzBEjXsPdVNXb6MPI4dqH
v7wc/Uzh7dv4dh2to0gQfrf5FYC5dfzgwH2o2FHB6+uCTSWoKYjaHjfKTsXs/sZe
0u9yl9LC6l5lhbZq6DC/euklGyNgThe+AxJIXV28lsKddxCAknrV8kd4MifHx0Ud
tnDPGCGWhp05U6D6eLDztptuyuLRVYoc57kbAAVQHuCLwNHkRQdxWNnc6NTxqREW
iHv4TbctPSsRC3q5urLXqlp0PSQp3n0WECzHBOnreQ6MRajrJ4Wl4+2AmZ2HT0x5
6NelnITPMlICqo9HsPn011uEwPhBIeZKOPylG6drx98E7lAkgppOCEdSykNVpLfz
6p0USonVYTP9wRRVsZ90gnvjKxFYktsI8g++wfJ2eaa8cnpmsvdN4BQJvdZp5IDQ
zOPnY04nmSysXusxK30k4crZZ9xze1rdMPe+n82SJsgZF5JRLDSgCA38w41eO2tO
I+tC7UDPjrKK8Hg14u9CZFUlcQKYO2qt1FY6QSHVGpe12CGwQRMNBm/Zqtr3Uc57
QfDZhVbqnJP0YinCtRHAF82DQC6/FQfcJIqSOGyPvKp4PCMswt52mywcP4X1hooV
vMK1O7v9os4hajnltsbPY2ra3IG4AOJXrbut3it1EtsJjqkam0xJ6czAt7SS0rlt
pWd65LfPOWN/5tt/V4IScxNzZq+/vZeRzpjgaeVrxe8J3En/7Vq9ysso0TFqTsOb
a7WHrJdlloNNjvxSkDKErzPImlVjIy9DtS0LwkHyyvV6Z0iPP/4zb9KKMa51Y/1b
JaCpf89weuQlBx5nqNpMJHwbuf6kk1Y86nMXKK+NMI9xY6RpPFLxIvERTiNfALet
zIEPbQLigt3moteFuK2ZsT3i4tbmTRlgjI8Ppn3m4CGu5I4JeAUjNeeieNNnGbNm
g7SMk6rhRijpq+dHgUeLVEzxWboIV4VOGUlBD9b1U98SVBwACnpNOHpshKSrI9qj
orcueBHnH33XHGDVHenfOyr/JxjZaWaxkagAuw+aUs6qjuD/8JH6b7lfNb+gWWUH
FOpcxb9AcxD61Q5ouCda4LOlnpAmlVx8ZjOcIqvaqjtSzRs4PeQdyy/8RXEePAaf
o743C9rcTUc38eARUTLEK6uaU7OSPewH3K+mZwOYvcnNP8B5q8ctEYFKdIYkSQuv
qrk1NfX6Q52k+kBob99chHgyjPCxUoez/b1wYXNqKN55ZjHkymaDEsJarnB2alkv
4XalgNFHnlWhbSWaNE4cJF2igstKoglT+HzoFVXMT5k4NHIvSVD8wkRnN1OTAvAc
2rS1XWjZoIegUBKHVuAs76YxsE8dc/dd9UIhU7ex+tLnNr4NgYUjYDSLN6b638gW
OB7kpwgfardlypRnz7+lQuG+THkJsgDJ82IkKYTQ86f9iobbr/M+BCwlKQB+V0Bx
QOFmB0aTNwTVKqe/kH8KinC9ORR7HDplmB4EXpyuwz8vS+Nw5zjTemhEnYveuViA
Z5sf9pTeN/EL7f4lxCmdZxyrWO9g6Yh5EqhStcyoPrhpgzYaup15wj/hjp/VgOBK
cuQ99MvD3Zfam+gzbw7VeNby7dkqudkPDvZxLFuxoMsMotSKbwf8HEYicrRkn5ez
IA3d490PIBorfRd5jOJr/l6oKvJ0qbeAWVmM3D7miq97kiYF2lX/L5DC4p9/37q5
VZmzT2dymd1nw8aisZkl/8O6MpYZQ4DTfbD/uE5S7vZqhfqdS3D2i38rMLAyHiZ2
bo+Z4CvCqq2pe3WjItIoDoYh/9v1dHiGRsvX6N2P8a1hx72e5opY4Y7msC3jjRJ1
BZjMjGCtRwAm6hKYAEPYeXAvLQIBSU7FEL5CwKoSNAO8UGMCpvPO5u6tU+TtLb2D
j6yEMRBwqvNoRv3a11WGtAZv9F66Rz1DJzNeVkMlcyhpiRz/4BioCyfnP2oooB1Y
5NM+ZXXVvR0wh1KiMKJBkETAGh+CCyBofuA2OYgk2z3rIhgKGILsqohWbPfqghQy
1R/b+s8tEdZzZCe4Q6pfPz1nOAOpXRSJG6AZIhN3xhMK0cW2pQiLlTNK4gvXeYqs
tmMQ/hYHuYHGJ+upkmJuM5D3TukZhBMSWifvI8s93qBxctUfoUvYFAjdXwh7arvT
yrkVESYy3iCYkDFEmgvAoey0gOVSsKJKm3/OqrThUGMggRKM3N/MdQhEe583IT/j
f5a7jwaaZZ8xBxDM6sExxStlrkEMuZFklC9atqdgoEHCZ2349HsIz59MNRQLBfp7
ebZDRE9/i5bMY5px+/10RQIuETPUUoI+HhfaSNWUz/F3U+4hvqBimqP6us4Jx8Dz
iOw7TmP7EnqtRgD1YHihXsBJjs1viWwcpds4nFV9JCmwjVoID1njHDmXOLG8qC2r
V4zYDdpOGyue6D8v7gYJb0LlQyE4+Xtsw93xxCjORa5AoaVDgch7w2a9sEWnfomG
aby6XpwkZxiOacXs3pTTsKLLvzJq28rJuF3V9rCrFOGWQBM5omHGcDCIXedzJlA8
PtGNwVCzJCBMuo0TtcV3O7T7AbQ+olyAJu6L8XtgubNcIAOobujCy+v9vM2/B9Uv
UXG7i0MHbtdukGuzJEfDwkCmXD/hBiS4ab3uuE2Nr6rr4r6Vv+O4tJoZPmOB1Lkh
vzRnaOm8KMY0ESlq6vZ0vFCg39D3J1hCfQwEQZIqk31t/DsAt97YOmVMxyIZXXrk
EYuW+k6fwGx2+j8atRXFhxTd0SsN9Wy6KXOpO7uWz7Y+mXtHMViNXqoePvfXGKHO
ZgUKcllHFOakfujiZ6Od3zaVaSJFtVFjgk2u2Z4ZbOGWhD5erFOD+24S6Eze00L/
JkNwGfO7SeXRonR98E/NYJGZQXEXBxtQTQS3h8nFDkzwjE44SnUDgO1jue5K7dbB
YGNWEJ9ST8wJwnhJuszBnSh1ENhd0LnSM8iu6JQuNhmqv4aqGjXzLXuAvcFytE+F
moBLTAehln6zx6luTw3xoRKc3u2V/R4HCvtM9V858TqpTMcnwhaw9PAJ7byFUIx8
71NGQZctgBuEWl9zLX8auPZDI3KgzVI30ToxReIZ7+ie4+lz4+w5s9gNj+B8bf+A
tll6x2waekSld+o8GmV9Vk9zkI0axMrhxCoPeeAEdwODDNje5nCCYNeKl+7+qj8m
oVaxoK99aI6ELg6liR7ISUga46ma3gGWZiygaHBsPIQ++bB1hjx5Lrp5oXPc/J/S
rfZqPBhQyriDGQXHYglA1rgXxEKP98a8W2GdZGW5MVH6Id8guaS3eJNHZ9otJWLi
LJaFUpAZrHoO4zkLdHZvMCfz/Nmg40XWTj7XJZC8LN8Qoeuk9a9Vs8z87uyZg28z
ogqIEl3EeDjQVGYveXLZT8jEzFXYgznoQq34TgdY83U4Nz/iNzYeMzBS4yiTvUjD
q02JRQQzdUimfeMbGqPiFqsptfRlpgG5Bj9byKDdT1WUGioFcHQTnMeq2mLJ6WJJ
L2D9fJ1lKOxqhOrcjU0hyzsbns5vkBV7rqJNqhvve6VGYK3qTQ7C7uYePYBPnv2A
Gl5TneN7Cbgr9glF274WncRW0VTOcL90wSvSi2EvjG8KOaTwdg2gLSn4QnN5v4MC
ZEFHkQpwqBi3Y5Hz9leV4Ui+OIB6FZ4u3NEDJDaBwJ8Ad04fSvktpKQ0sy7YTuKn
7ziVziAQrfm2so9FJE3McGYOVm7r9Cmnc95+3Np9erR1USKnEfTJXtMIwfx06r+T
yWM/+rmJ7j8i42J2cD8+ov3w9y/7xvl4BPMhJnA4i7fPV2icunOY4BT9NAZq0Qwn
t29H3Pcm6rs8ZDuyjqc+aSKrvQgjdMY0Vt+nY06Bc3UuUWe4V0CIgQabmEYIqkWX
tqd//cHTLtqJuN8GmU/7hctcS4pkMJKZNu8pmzBSUcyCHpoDAfFSF+wTcqPbVJJ7
SkRPySrH398pVTFlf3WR+RG+9oP5UFGLtj8+ks5ljzb8z+nQIUlMJgF+6Ogv0P6S
boQLL56bBqKLF+/+fPZErgxGx1aUgkchFzRwtpvOMCagvvmeJIvFKFihpvownhV1
J/UEcQZkDizGAnlDcyrULSzhOFUnNll07QJ2eiNIkpDMx5FyatTzsJ0/ASSU5teR
F4Kt0UQ62DlNc5XGPWiwJDe/tJuVUpS5H90lTNthV/a7p+8LtrxlhaeGO4bv02t8
PQE0yJugFx3Y7bET5jmEtnLSzszPDTlHh847F0iFym+YJHCBK86V0AzrWNsGV+I/
Vked6Cum5jAaNOj8P9TjmUofTKBs1h9AFiM2OsbUAmqfH9ZjrTNaS+ZKBRmrGE5j
Wbbv3FwdaHvctBI1B43um5yH+GwO+hAa30Sib9vy78Zl+BepNLvjojp1aH6YYONS
3GtAvRCVLgAJpdXSJtqSUCI3tm+nEO6iO+rQqyK0CAXpU5F7rZfOfF7xe6sPkJjQ
Pwxv+Qit7P/6C8W0Nv2fAs7mKCHeDpQzYSzODQAaZ6fuek+1S0MA+xxWoFOzUPoQ
Cn3+XoyG67yrbuxPmPzyh9TgwfY3qZvBMvQXP21G6BukLQP80IeK6RxBVFUjakz+
4+XrqNB8K+awGSLmeAXJXGBPX+B5JiWlOalFjAfJU94PVJqlshWu99a5KY8fPGJO
5+R1/dUsGYZWkr3R0C03ZVrou04rWVvXMVwcaf07RDrIMs8aa4anH92DjYM4ieHi
7vaRsHmeA9bzwni07dLecxDfPanBM8jSzC5vLQEtw8WI/fzwv/KwbMNSdOmCbBUw
A7r0yl/ogvEwcySX13oxbnDgj5n7Ed0FsePa2CU5arHj2YtSe2bHhSlaRqBuBLz6
kNlEM7yygyLhAdmUaif96/tyk7S+NNeQJ/rM7Q4GRmbhTo1btAWjCiyhFWXI6ny0
QU2/nnxlpGh/16gL7tu78zckNUyFOGdIytQfsfd4Oo958h39t86xbNHVGH3QxjWC
J8eBQikGSCdFb3J9iOTrn2oVCJVTS/YeWVLBV0ZNDRmV7GoH87lHxk7d/jmAkKir
rEMf26uZu8jdu9uLE8E0pbFJNl0oWMY0bjXw/CHFNUeNcmBzsop95To4Z5/ZiIhm
I831y9c0JdGmlbR4m1xVUyrER0riI4TW0rBMEUFf9q1rs9olG520+L5QxfdE2Yv3
SGP9Oaxc53Mla81TQNb3S1/4aDR5giI6ePyv0wcru255qKBZdAhUQR89lS+pwHdE
FAWypom39m7m/74NZUdL7TGsq+tflnynH3uc4arOp7oOUDVYO/Var4xEvtbMhDW1
LEdzd0D38VRYtd/i6OpFenpFDXFVqCu46Pee9dg1FtD63DSGxVqF+p8fTKw7QqEH
lSYanxVEizlxVVF5FPdFizGVS2j730Xs0ItTh5R0gFmFcsoShqaXPkzt1v/J7/mJ
evbWBIqsQNNgfqDatwxhun+Ahan7N/Xxco97fEsPWeoFB2/y3GmQ7tzmSY03mp8i
eBMdwhEqQT/AFRZgAhYP2M6SwiORcfD71J/YOWWCzWXK3CLZHtuvIoZYuMt+Xm9+
CBjsIox7uhsPcTyBEg6r/mZxZbpHzv7b1vDzUW4jPUippY2TZzoX4feM2p1nBgDr
pF98Iny2xGFUWw3IeLq0xwaENY4J/zfGaAyYlGgVHzqrJiATxNUz1duU3Nf1Qh2B
N1jmTI/BsYDaV9qNLlw7XA6dpTGGqniJyQz7BTl069CLvAIizj+b7cePk4jsS8UT
C6nfGfSFNqOaRvMkBHZZWY5YhK9UD9CVY4VcMGBSQf6CdErcNCDrJQJMoI2IgLyb
9WWLP79dNylO+KYqbn0v1joa028J3xu51NAxLoZxhMolcpEIJXLJPDPcDY56UIlJ
YzERVqw7CRgeQp0wsX7/IaSAlHVmUyA20KCZ8fg10thmhNVu9yNytcqpGESrjTHl
G9Xh+enkMXQ+0iXsaxO48ncUXhp/Tkuc1rguojsQH92RPt5mVmelnIFth7O0L6ht
Y0ZjUzzlv9HHj6SU9Uw6sRWUQkn6vv2AcgKxz33deeMan/gg6SxSzuQ5c7JeOBdp
Az52RGRp0PcQr21qdYa0cb0VUzpWmQXtgHyJXozoMv3SAezDZxy9VyjhH97Lehlp
y8l3MGTq1Hp9HIT+Q0uJN9wLuBUdurL8OzwNIia3qvfFQ75lnNUMLoOvzMsHVxI9
0vzLPQ+KK4D/oVhnNcLUb2FTmxiPD7OXAHrdXmSN/4wtTPqsqqCJWVIMS5f4DPI0
w0eNV5PdkcsfZzzkiFVjoDNZtKOCqklbPj5mhMbAPh6vufqfUJXV7ent4FPU6eHg
8rH8PK33w6SraRoRkxOpABgHBKm7P/884AYMJeCI3yGpr/HAACStDhyyiFi5n6zD
W0BnEzCkYfQW0D8FbYyvADNZzPX43xZfkHus9JN84UEvtBySqDXh+evStxjuLtk5
wT6HEsOd+33FKQ/HznRmraIaVjBvI+qNlOgcFrxKrnIYKwwGBtPr5QL9+OXMQAf3
9rre8Tv6OFckfNO1n/h8huPH09lujdkXQ6HuahZZ15lE0FS7zBe2LGlSekOmRiP3
FFD6CFpeNQqLRjPyskNrCl99vqHK6wjQVGcujNbw96pcdjdVDMNFEUpJ8/iQUbIh
NmI2Y6dn3FKTXZlHBSCyaH/6hVD652kuBMqBA3ObE4Vc+xibJx2BtoOLGqXXz+rX
42ny4sumnJpObkf+ijiUTE5QowGN6oqVptUHQnRNtHLEyUYhKJtXjBF6xE9BczYj
j3zAJma6yywHvqDTIyhpVpotTdpkVRE9/ETweChLGTTK1H1GFfDC2CndomsCkMiw
6VlX6LcSxhwz1efrYu19HPssbwJ8IiMc+LTTTay3KL91I2Ma9JGbeZtNvFXAWsFL
R5TQKeYepz2HQjwQwiCjGY5SYT5GTf9Tv6e+Gb5csaJbbe4emuCRSVAjJhgTx+Z1
Ouc01Ced1CE8nqF5wEFkYe8iV39kP75gvoRH23smO7n0jsQ9KIoaNtY+OJ8S8DZ5
nb35YqETHTk2YQDcna/Fsv67IIl+Oo8XUuGfhqRxF/HXgDN9bKss+vFpWy1njaCo
wk/Z7TryfxGZbXuso1ngaA1a6fsm8H/03Q6/irtJvNO60/I1grTJs1dN/gghQICw
CKILTDR43vLcqgfncczrrepO99pr30vMnb/8nZx/Mc0XyC54O3fopUx30vsWeZQ0
6tkgiKuQgfLAJnxTySO8mgRhuC+6PHaCntkU9H18ZmAHDnHKC6+KIz6UpphKapPP
CXrxMwb+CLLaiOhmYwFNkRHr65N911Eg7PWLlseSYST4reXsD659Jt5mRfTqmmCX
M9bp4MJjYOm41vgGVnBMeABXd7VklswG+hfP8eKebuQQ//29riO2akOZFa1fxFyR
9hOoY2decIupFup6vRjzTqoOEuJzfLLSae0A9jXzHKyAkXFf5+FzqvR9Kl2Nsa4t
JSXstIIbS2FpbPH5dMiNJ79PCWV3ZzPf7BGYzyfKZUwe0E3CWyF1tlvTQuW6Q2kq
LdAvfN/Xj5s97a6ZNfLwwBLviUFTjZhDbDElDEB1xSJ8Fg5r4WcQhotoxrV63DXy
tYRiOUaoxXdkoWiBPxx5T8bjA9L0Kzhd+5+03chgXCxIM/v3VYQxMo6pJjJHYfQD
U1YXLnMCs1dFPuh/m8nQqDWfyOO9RY09gs49JfJX7BYL8xfrOfeY1fvZrNeoJWlI
rQ/iXxvEcHHZoOu2ZWNdlhSgq2yZTAiR1pRFplxZcEo5CR4rOueMI8UvmFnJHFAu
0YP3rTRdzDv4yV02TnSQ/tlJG4OaSGMZaPFKUgggsRDZc0bOBhu/+0WME6pvtNu1
Hb1yoVtLw2lkyuxpiAV/+EGZxiHR/nKIGNeWVu0LFRhtmrsVIpOyQYGVPaKxTea7
12DGepPFDKW3IBEmNITYDEP+HZWMJbKHXESyOzguKgZExSNUD+4jp/WgzjSdAEWs
odN4nHIMFoQXaO5XvSo7HFkf4eJIR9MnzuapiOd6JVw4WoKIWkEby+69tnF/A8sE
XDeXgJyeOv6oPi220+eoBiONu/BThjcgeBbdcQaJD6OhvsF4vHJylIzsXZgcjBB6
4TV+VnsgW0lP7BnBd3kG7lwDgK7Jl2YA1ZY03cd9p1tK5q5fhFFaMVotycHEnqI/
WnH0lw0rSdy8ROcJR2hatdEu4x4vX+hNZCqTMqrzUgXQNB+KPlJnKMcL22QbPzG6
6fr3PZ71Rz6iYT6p0ry9AWuKtDAV8GBHKS+bVEYX0MAy8xceFrmPSyylSMq+Zx9w
LY96cIkAZkOIO95Wy81q6dNb4kMIG/ynsPuQMIqFDBEV8nYdd7ZKo7kHWh16mNCD
Bfy4dxcjcMrCrHeZZXR5C7HVXR9BwK2vdmzziicWiFmCnx0AYgV44LVRVsoIz7KM
rhwwN48dqAZqkqv7aATLA2eUytAQeq3GAvMS0yQTDl0nyDEr0ZnexgGICidrCwjW
FUgX+XatLo2M4C8ZNeEQ1RZT6g5z3Y7bR01kZJedJwzl2dT8afE00PFYdWPvekNQ
Lu8DNOTJZ1NZbYQzEpHV4te6BxH0AQo9g+8cJq0r+2ZpEv8uCHC9lO0+BAM/SrCm
xF/wDe/LBr152XP9x7HBP+8E+6e7uEbzlWUzJ30mfQHGnbPXrSP8Mwwk+Dt3ii3o
Jd2GLFVtM2Z2H/r60DRY/Reg/TDJOAJ7AhfDBjSbPImBsGDJBPn01JxuYCUI9Ans
9C4J7hd3UCAVFbIr2mAA1ldBXTvxT0NstvwcL4pq5Mlm2KoKkGmaAphBVrx7ywpA
QggipHoYv3NvOzAKCtPYUGqZoKUhO5qNSdjEsHGTg8cadlPq5oV8NlH/dOXVg1I7
yjuxu4aIthtBlE+kwuxGN0zrYDvBXlm1+s/PBHMEPKY+GEIy24eF2kl2WstJpGPN
dlnKmLoW28r7k3l+g3RoKzG7wdMvhs8KoN7wEIcMsQvZvYkP6ATLNQ/m//HqTEn0
nIxCfhWzX47VwzGf+EZ3HkbAcT6XMmXrdV+Y3EXTCBDE+3rBTBewWH+1dg4w0kju
1uGA5rfhgQEGyTNbs5LUzDv+yPAzsuoXpzpaPxVEz1DUD8skXptb0nOgl+/X8//S
S0VY4SDCqR8yJd5DGS+sg5hvz3luyLsZVRoSvs9xmH9SBw5vccJIIAjMyb9S/Y2p
1GTUADQQkVYHIEs6g2sFPs7BBwa7kuk2S8TlVgAgQWDKo9MvcuvL5mtWkwFHLzdA
2BnKXOgreAJqSwuW4nEWFIRdr/03b02nyeWwuj75qOfte8Yvw0zrAFRpv//artgl
tELnzeSlLd4jJ6FF3YOfIHmtFz1JOz6HWJiLSsJSMIFs1RkQQQ18hEWsUXJB4SvS
N2UektoziSLpkc4P8i+zU61KcaPZ/LiJVIu4tK3oKFr2/3Wtzedp/dr5MZuonP4M
8TLrJKGw1gM0f7i93UhRtQ9Dj2iNdcY/4xk3uR5FiRTZ+pzMqalC2fGFENMvDW/3
hLHL1MibgJQzVP7swM9kWx7rwpjpuV/xWj1oT1ZFJrxAKHsCU1TVDbaJWuhZUCIf
Hvdq3avaZLsP7biQFHtXX3iNNUEZkY1PEEIQZFdDN3cakZPzsfAudOjLtZJhL+3S
uq4jCqlJniWzaauWFfoqGvJ6c2OeERjGdF2dpzY4BDStVfAy6nK9SZTBtY/DBzGV
TD9lQ1trQ0k7cyfQwEaZLxaF6zXXnsgTEimRwaxZqd+1cQc59eH/vlQ1hez8Jamu
HJQZlaXEWJ/XGCceG65O4zBYqTwARu/xIsQGLE+K+l1EbU3HH/9gnSi1SbhO4l+S
TZtEgFnOtJqPkv+wkv9nd1sfIGBHSwQL5pnDDwhyiZthgpINqwBk5WhRC1DnmLkS
dn6E9HfamOXgxXluKoibPOy7j6NFqcV8BoU/0Hbm7vvfdkmTmtTFZ1GRQc1r+1g4
wP1YxcKiB5TI2FLfA8XoCWnGy3VKrHzm2UVIML/eS37eHk136viviC4fxQd4lbxS
fOTijXwdmwqD68DX4I51vLgwB3VAc/4cY4euwRU23Ii2JqS3p/hKD/MuiYn2/lf4
Kr0m/IMyvKSqtve0Mst6ldWXj24O+glEjtpYdJrK6GEsROdYb6qmP4cSH2Y0diWb
fmENkItB5HQFTS9bmfgly4IfDiQ0SYSouQF5+AdsNms/rKz3TZQgzS3OjTPb8zW/
hJiQxXlUawQrIZNjXdxcbX7QjhHcNI2y3k9UPHkKLL3meZu8su6t45++3wqjjRDN
qRNfSMWm19y+AM26l/M+8pS4ii5vLoBrAJF4+5VV2hicHe+XHtDQmEJnAP7rd6sx
UwM1hrvqv2DB3vyWqaqmqh+0nXfFFeSSFvMNvrOLAajysx94okYoi+c9Avl+wm93
WL1j3ntI726/0jChwrCBhoCP5jFH3A+V+XdZo9TWTL1DN0OCqO0URDQUBOXQjV7O
9ztLp8E2TflpR31fwxk8aM9EftoakgfZDVdTW/A1hj2JbUbgwa/hetCkBV+wSaYR
cwEoTew20k+sOxbT4EyNQTNLKXPU9v2x70dtIZs5cfeMte/Sjt8XnwrjmIWmNxbp
Tglz4Cee3Hj1PJ2edX4pLNs8pSONN/pgH+ayAbL/tJ8jRNzo0iP11+uWRMww1RXF
o479B3+Z4yYSlfQyEBR44DWdwHxU7bZk8ZUYvUCQhOQzVj5LSBwMc+FAnmgp5+Gp
PbpeDdzqdnlq07jlug0EhpQyLKNUAslTCz2VomX2WRCTKjUsJWHhQn3zma0j+zcB
+1IcjFgkwOc1UIrNjz3Fkwkc2Y/37AGLBjU10AtrmgJXVVK13Y/W11NZBcMO2rkF
I6iDlBUEQ90OK4Rbb34d3T0uqIMNr97fQcrYypRAbiMLcDLhYv0F2CRrol1t8Kcc
Dkvx512Dw5HhQDBtDmzQ1oRfkRRUsS6jC00pX6muSoGZMUP+KJjmx89NOHEMMe4D
FHjwZ095Z0NhHFJb032zQdcSCnIPpqWlMDRNG4PwUQEkERH7JL5k7xdHRUTHNLCy
fMtKKkTp3/SvFFz+I9Xi4AU0Qb5K5lrtABLa4IHa5IQSMlaTLsNm+rcve8Z64WlY
vnbA0KkKSXjU76i7tCYwOfH+IaaYaEmZXMKJVS0DFzYcd2NuTTWkuMXGkZoybdTp
LfEnbrEsIRYNE/g3HSk5IXvkIUTUyFic4cFYb/c88GX04PwWeXHDWQ/PtwzWY5pE
73DhSpbwp7EM/4DcKYIh6vY6BJB82LyfCFPR/igmRlg93NfQLex5mUPtQy5MF+gF
fH3/tX2Dz+KIfq0L1rg9nhSJplkD5LjE7rxIBcG3B/nrxl53i3EcRCe6OI7srkjp
M9f7ghIa2wQhbGLoabIXliYjVNMRUSUAtUjj55GSmoDbmbuSlxn3aecuBUOcgNAF
E/1znepWsmhlqoqaWf5eg0QgZXqIEUnQsdnSFlxwzmw7DBSLLFb0S3R6IX+SyfBV
qCN2RreOUvXR19MsUjkT389UJx/IfLZ86uEU7GxpAlpRtD9bHTVajVVFSNWQIJn7
kNcrqQw3Q1blgVix4SMDZLbf/pwHG9mxmfIMb+rx+h2C3K65tc16/LOtjp9UPYxU
qy16upi2tdrwBSCYoBVGvw3pw66z3+hrvMRjpcDsaXs49z6GwsyedwykLG8T0qWf
8RBRWtiqW5XEvnpxKoApov3M++blP47KMuXqcPKRdJcdtYciuxAsOusbSnyQLfPj
yPB15hy+FQWD4alcXEvOHUQFf5RDsYytiIId5mg8vw2XvLptPztFIXFUu490ZmCJ
lvVuKl/hc28EcWA8IyKyx8ZdDlFB0soL3f6AbjLnw0BfxZV0BHoQpjcDlfgUVNod
1IzE/vong9AwHXvOcyhjkyiD2jYsacCtmvicvu764KvuxUe2fD0QscLY300XPXag
snTgrIuJH6/mEkzPv2WT4waYXlLcFVZIUnWZkWV4OKMM8LDau4ETH7GsrxCPW0Ug
Qr9TZJfn1uQzSckDRczqLx4d/2x8wTgFMLVJU6isiGVp+IAxpU1zmADFfyOI21YJ
j95OUNVaneVcCNDa853KL0yENYd6LE5SyeJa/yzINq+pxKn/TJCF6KN0uNWYU7f6
1zQRg6CLi7yp2phqGicsk7v9zA0Zl4CCG5P/xVsWASSH6fFanA8Jkha9mep7r9ix
KMErSMXx2E5/cwTSYbnOzKi+8gOYH+NyEhQLkaB+Wlhz0nJ/rcyX1FbY1zJGIET0
BOUoYIzeN0Wq06gSkYYodvZfCeM3ySBCf7iWsPfxbwyIheOhYCpTEzYfkSW4l1Nd
Fq3g51PXuJnSf+AMEd05CbpKzcYvu6+3whZTyNvWJPFuH8LCIl0ipShePX+vM208
4roaN1vVnX4rLZURTsX8zlVvTRdM2HREUa0pu7B9Z1JoAHEsaqRcUze5LJEZN6hR
HhiZJP5uRU4T74YPeMaMBN1KD9AObZPZqwsMi7KvM09CZAwJdpsOQ+0wCDN0A029
u2v1a9gltcBUb1KdG4RjNYT+BS+iXQyhcr4iaZWBj40ECsmZm3Afr6uz+bLw9K03
t8ccoji8cOLwTuC8z/tkDf0KLRnAPNcojuOfohKIL7BbX/jrdOEzChj31MD7m1vY
NM+yhyCbNKNh0K8itj53HD64OWzAy4Ci1Ak2+p/2b4/q10vImOw5aGwawP9ayeZw
8BxLYF2HOBtFU0pF5CAa1WRJM2pIhlhV3qxw53Bul524ccXl8S1mIarZKxt7ZDz7
9wVGM+6RK4KKB80yg7w9Eq+eZzvLxQISVO68f/yAEo9ZYtrsNKlYG/ZMjYDzbZej
IJIExKmsuGOyiQxi1wvO4wDX34lXHArt2l+hplzZyojr5mf/vx5z01hccbSaSFWY
RcEwP1k3lVPoGg+NaBXeOFQFdJG1dKWsRYY0iA1IjeWv0x7yOPZE6NnQn7ubRbTw
cj+Dopy+N11KhOuVDf17ohZ5ng8uDqBgPhMX48qD2oAtNk5qXby7wCgWoMwfdX0E
KHO/Iav2RR/3UUR54HDA7NRBSLG5Y04es+zMiHnJ2+HCGlCmLllt0vlzR0fotdUf
QwIzprDQAEO//lp8W7Fo2+nw6iu5bWRGD1ajeNmDOnGiNNNEQv67f/m7+k2eUJto
mntqDh+wFM+OQMAuDlDGIHz6QJKbh8NIwxH98tP6MSAm/0QYXW8Mz34894HyjQLa
Cvn4EzqUK1E0HKG61MsS2my9lXbf3XuNyhyHBxD9Mt5TwTpNjwlmSHg76m0PxX/x
czdrYXcypqIK/KwDPldq0iuVpF+7esaZlrZxJAXcN2hDJA9asJOuF+LPP45Pq0/A
RsSiPLOlFIVHHIL7Q/X0KF1vmJlEGFrjWXNAXj7poyBFOFvScyxgf7y7wyT4MWO+
2yD6i3RJ0n3OjGwCg/Aq0OGghbWBze5fuAhhi5IoXHU69G/33BHCY3qGNknYwd1w
EJv+AtKhOfOTH8kuL3iQ1kkzmqBxJxlNC2Tpg11lqQVZc//kLcxQX0hBre3uyb4a
xDNvzcawh+4YgHLquqVm4rjJxO8/0Lrl3Clk0ZL5fpy88prf0nToG1BZJDEcOz8Q
azXCjmKI2YosK+XmK6gopzwXQQW4+aPgTqXjyW57PkBETzFo2sFmhs56kYheQznp
034qvOqrSo+XO7kC1NTMRdzblRfIKvnX3+N7+N1hGB5DjPIlXgbj/XWiptMKG3Ri
viPiR8d15UQ5XBdLufDCgzkU4VSqE9zV3EuukUCH9/6Z9lagbbImFxZlosaMC3PH
a6kSxf8FUTmcY65649zjuHkrCESky1cdrcLBwyyWRf99FehO18grkYbLVvyKkaJt
pAlrIq0TLEgdtcGBCfSsU7lsz/KBlY9xv10b7emCskfXApUvayGlyUSldpXEyjNN
1gg1n0ILptZuc0IkiyP60aptCG8pwro0uAViy+ZH+cxhRNSdN4GL2blQ9+jnMh2b
fBDpy40YkKKqBkGWqKdf61MKwhrZVEmepekuNcRGTX18lJvnJhfO+chimD+SOh14
7iEb7sg9yo1mRMaQpE1+HAlOO1/Rwiu0TFnH2RaHrecLHqzAQL64ZoN5s7MpbAli
wMzesyjukvWx+QXUl0n9fakxpFV0+y/K6PF4cntpkUG9ihJpa5WTDX4hwVe7MM81
f/5cgR7sNnRkyiwltBeP0q7cHgyNUuS0VlGeXlEWhtcxGIKUcaEjiK1RnaOIGSDH
11EI9rfLlRDrzEXoWiW/7SLQLBtHCCW9DpJTC+2p4yHgaieeNNeLSD79J6yXBTKB
xmfsJ8cAHcdtUluk1R8R/JZxxypzp7irTlgD9HArO8XvvoauWORluWTiBvlItd9j
0HA/Q8AqySer60Bb7GQ9+dh1+Y4IqlOwQlEPx+yXoOnWYZeu9w9pvnNH8gobb/Yc
EcvHRjhkfAATYeMwbhGj9Aiy/T9qllz2FaEh0zRsis9GF1rIOkMPdT0v40qDRaaA
ft16qFMunvY4w7iPjIepGJKjeFR9wFuVZP+HZ+FG4oM3sTKZfYe0N8jHosfaETz9
jjOFqMoAj3EgrhHMgw1pZ+YSbpxNtrPaFPKHX1iGhe676LC5igsjcJMbXA7BLBqU
LjQ31BE4KBOSOXchri57VUwC1K6PZUhIyUkpIflJltUp0LrI1hQOCL9ot6nIOPl+
m/+HipPyGm/cpaBKYwYv8KuvZxiBcWQnHYji6ACKTjImJ6xsYXZrwdMc2o2gIRvt
0MFcmPRldher/xHYWbsgV36xE4DJp2d5UVz78gGcL8Hw06iKmSKVfyCucY7deFr3
jBiMnPmWGEM2t6gpsilEQ5hpHMft3bXEQwH8Tugn8dU1PYe3bYawqClw8VJHGjZY
xWuWKanvesl9pooaeZsrNkCNXhbwJ86GcuIcGFsecHGyiQjcBUWf4gcatMNEfOFQ
qT9zNDuCbeS9xp5C9RqYvyQKAJaSpKCQ4g+N7l0iJS2I4Y6Qjn1M8cL7hc83aOiM
VBp8Pzc4qN9W6w0Ib4P+mYAfvliGDWHkihb6c7BpXGDGwJmGkgwQhugAHzTTdP4e
CsgG+nU/+SKnHXFgs3d5rjBOosNdRuC0gjlDd1PHuP0kEe/LpQDaIGZecOLKtrZ4
D7cAWHUGCwv5efgFiIuOVqrowjUhvNIwCqqYv8lZsXKEOBDmUmoc6sMsxxvDoDNn
qnBJsi3lW3Z9Z6rxI4hCjTmoNR48/YQYmRKCBriLt9j6KTSjLloaIh/NX1/22IKn
jIlsE/Sl1lTylB3Ry2Li4arZxTNygR6vJKAtKJsW7jP/lGPk4Jk+b7J+1Xg49taW
wfD7XD6amFTPa7HNz+B8GRTPRrq0V104p7yD9zwmZaqt802J4mI3b0RXx3BuM62i
d9vDStL8IViXo/5WE3/8vyXT3wnvTj3lVAWyWlrR6PWuOKBJSz+jdnurnX2x+BF8
7M8L4V1EDptjoV+ODHRq6hSw+ryha41X9ucCrF2GGa9CbjGauo9mjqoBQ3WcU25v
DuCBO5XEelwLUd/xoxR9UnU2AWXNGuBxyckofDxLhDtAbqH/6iFGdlfY9jTa0mDt
GTgYlM7ZmUq/jgERcSA7vxmIqbf3jHZDfLTP734bebAv15+zErVLbVYUifYg6uzt
S6jCH0lZLEOMx/2tYkIlgStl7AGvDVcl2Op0s5vxk2fx6/+vZHfE7ZFglILh+LDi
12z0pG5uimoAYy2PV3H0fwy0wM6UT5kmYyE/+vatbxGzNeFer4xO3ZmUNWTohuPN
fQ1QmGrXL2+NK+HE4vizDGwXoGiDg/Ng45pycy4I3l+7f+uvZenAXdIr6v+yV0QL
gmHRyV1IQsXMvIZxHhkguHrjfTNrJrW7197lYfxjXF30QwZvMywKlCeSZGeFdMdF
w5lBpf/EAzhooU0cGdGcjVDhVKhYgpTrflFys4Yu6mSt1iBz7CPVF34NMmqGmNr5
KwCYh+98eCJMKoTv5ER9UH/J+g0ZAoswW+jjXLk2wn7hXWoWrHddSiDpDs1qw13r
UERr4ApQgAf1OHS4rDXEovSWuID6uIlJ77rfyTtq+7NJpxV9YJI4a2DOceDlyeIr
Y7vRNNNUJZvxc1p3xESgzcnACNrv5bZpwxQ66FERg3mhepUHCse9/HPZQk2B9VQu
cl6agGt3dUkfj/piv/tnM18NxFiOWGB83Oub2nu1brED3PiG1UB56seVk+UDifAI
NNST8/vAeX8gxf+YPtIV87T24BfP/KgbIXc6cu8bKIQgQGpsAt5MeVtyUc4MTK3f
SSrmjge4WgbkGcBFotcvwXNmwlVvn1YetOWdBFy/mDPb7UxTOJMXUgKwpqaU8kCM
TJ+bLoil2kxM/9b4llqZLE1YF3ZowSGHPOj+cUpA1ZuqktWSU906pekrDHq1RvqG
TBIokLinFwCuSguehs2gi7Hkx/OZQ0dY1z50ssV7Qrdo5kKX/iM14/MuJvvwPsDg
Wei57bK55BNRiEonVYHwvFrhFTDAuhjJ3aWbH6WeppefAR4hDZl/SHBbX717xIEr
W4ENApJVplCjP3Dvaq1eHO90xOP9YP5ShtRlxdP0fuq21Cs/V9REiQqG4eDqzpan
UIjPi2twxOdDfPmFaYuAvSTigAFyqxtXi7dIV/rigWGGFxXflr42VJMSMqmOtct9
rB3QRmda4+ukPJgWHL/sy8DfXwb6vhvFKBhDpHBuWENHXtsSMqZAtfbmPAs3BA6J
OJrY415S2Y7IiuF2Itt1vzl9UZ6B4nhCvTl9EG8BLAruZ3HIaCnjgIbXNSlyjSwv
cQliJ28aT2PXHE+Xy+LUH4ORs4i9oRz7z4DmQHmKOWbtoilvCCOcaXUMfcC7fwvL
vQKUderH5kKjHKiZCR0Duf6kKOPIVMESPvcX94SC14T8E14g5zjEcZGY3wlz6wKV
ezXlKDjGsOm32DS2+tq4P6/o8foNh0bHDlR7sqjDPGqVnOOGJEQrvZ1IcAY8adwm
JXhyzkOiT0r3pkknug8pYbVuoIOG2/2qY04hc75WmIVDS9uT4GKzoJIIp2Up6Dt4
vfhOpjfdo0fT6xdemQdHdqEXjTYsPRnd7ZE/1zd4/gXi/c82JwyDDcUTKrK4ZC1P
/iJLU1Cuw3yWL3D4hXavfFbdVa118KAd4+OsfxnbrxS0KPjrNwvQrOmW1MBHwnrV
lD2W/EvzV4Se+XFnndClOTIE7kHCGBt52QQ9clKmtQ5AyvNZuMBkmb6ZXF0JPlA2
WQBhcBfduYAYLpSt5aGdSruLuZI2Vu0u/Ncr1/lB/OBNLqMUc19+Hf9+/th4WjC3
QMNgQiX5tew4wPNGe7VMdZ1aDCtgSNVN+NhImhrNkfdEX4JsNsnch1xXQSmYvc2t
nf2/5lI9m4Q5eS8QbCLvRYHF1+0BAwpnsYw/TpG1OtDhYf61y/z1RsIT7VOEizWV
iXLKrOaaf1SJxmOjccfk5DzqboBY7K1BKb9YqqDQs5MXoZyJ+zum6pveC+XRFVLD
qDhEv47l29TlrSOU2rDlwlKJJw/Js6VjHlWjXZ1hzmCv1wmo41oKueAj6OTi22yf
wXmFedoRmhsTs5nQZCweAxI7k3qPj2SAs8Gjn0ERydYmja7rOsPZhgRmNkW4LFHV
tsP9vLbx1OKixjMSVMLd1QsBMg80Wiu/yHoOEMRcOwyC2z1Oryvjfq6jkxejOVLF
C5+i/SjxhEJnj4FZUYBD7ymCqPkf44njiJsQAfQrPvVbzv3O7NXgHQuCe1NZiA5B
cDBEneL7MagQnZe1mtP/Z3KL9ilF0gwB1nyxM/iXVUc1qWKz5iVXfpEfHxBamub5
//voTS4eAfggvsXtIMaoue+P2pdg8IEGATEbr+phfdC4eZqBWdRJPAgSVKCdMPXW
1bv4jV3sSzodwoPQM1F9/l/sXtqDGG4cCW3sz3xW9msZdvjujwfpV/IjL/cvQcEU
NMXDn0N+tSEG6aAZGk3MHppXZcehXsKOvTJt/nvgG8qFtpLz4ylGqjyLPJU9S92o
ehtY4jqhTj/9IrYfIdDG47E7Z43ss2bMKjsxOl/3GVxHob8spvA2XPY5fFEPldMz
phPKCuutf55bsDgeoFe+p4vBtR1RWP7FynNhpXSJkwqQzj9AtUb97mg1EaIlgo8v
Kv3TXTRETsKsOJ4HbRdHBjeYm6XXiAYi/KWRXmwO+2wxhbxVfdjIO4U8r0ZDwwNr
+yxEawiT1inUHBL99EbFOAqVYjdE5t4Rpbt1Ar9eS1URIMcJniXrjbi6jbHUTG9s
/S+AFEdgyzav42fIPdixTGr3H1v2vlusXyCCwMqiZygT5ig4neIiz0jhz4SImFFl
hhL24Z6BLP/WyYpnyhwwEtxDokQIuKtJKLTgRzNsVQ52pG9pVEpjvAdM1zpM/pRc
G0VxWmRogigW1xr593K359+8STbucjRIHIwRxWbF1BkrIcpAeKPytt2b/KMxTQFL
muO9HFmBSLA3FLssrUIRVVVEbVqBO1WeT64p8iJ/jMZ/7gP+aDzru1o7X9u6KuOm
7+gnwrJoAciYgyqQOj1tzf7gjBzt2TT+QVwsKGyhhQY9qw7tlIIon429HD7LYmjZ
vZZCzAAy0/KA6SzM2VMmcCZ9pbZigNd2S07P1BA8TKMhbor1jBklZ2px5K0bpSp7
UOUt9x1JgG3P9SyDKucXBxDyRunyphULDWWM7hKWEo5SKxVrZ5FlFzPnEljLxcex
NuO+jjsDNni0soVneUs3AHAk6vJ28pubW+m3BHc5QXT+AXqoHXGgeXw/OhO+1Vh9
U3I3krGB6Q6QglayMHLfmFFrP9c5z33ndZWzeRl5POhnyYVbilorpz3BKMUMBZBL
I/qDAUVnNmTt3TgR7iCfv5441ewDlhSXA0Ys9QNS8kfFETKRWv3vKOrPMXvfzxMq
m0BUVnIJFlZ2gioxZPiTuyIdoko/LOsYyIyKSg0w6rBUu5OT25A7jxiBKoCUb32y
qkyshz9SwLc9MQE8RiAaGwQiJ8Ubifb0YVZ21T/New4LjJfq2Tjoe7ps2KceoAbI
Au9+s2vbt96kpG5fDawW1rVjKaSTDU1cc0tW5yH/SKfIRa+amg9q5hN96SSlrWH4
IXmede8QnZUXveBnivW6RLXlaVAalqMZqCMptkz2Jxky4fA9F9JGckPJQjTPViH3
9g06Ja6gW4qBf6uzxcmtqMICN91HFI/4A1gTCgaW8GehW9EdNNT8/TscotxNOj2K
5K6k0jfApgwMCvKwoI38g1cklTXqOmuPs6yAb5XnwKgooOrR60dAiCBJrUl1C6ed
QRhckLjsYR+a5zZyhuRJzlnjg1HgQ0J5hvq3kAGyWu/+oSCi3mSru448reesjiNX
oyJOPWcN3i8rRdBYad9p0QtqMQS1tXRMSlCbc22ctU6yYreRya4j/hqKlZVuXxWA
RKiiZVBRfidbmToXiGE2tggqCojpUcY6MyyeMyvGZyan/xaY/voVUTycQjR9+Osu
BsMN6ITmzL+cdz9j4GD/iaC0rduF5B8nlbSkMinuz2Hbla5FsvYByIVtejeSkLK+
QLwkD273OyTlUp/aqJXQhZzY8V+r6wUVWCx1YHIxQKYs/teH7ogYrwdCMzLGB0/L
tfTU7KyopedgZZ77rguDzBmHHNseP50RR7I/89XrCtzoUIuvZn3+L1If62aaHrSw
1StVXYN7n1LGOlFemsxalOZop0E9jzPR6mpX8z+x1/7zT8hQINYolLN6nVAmb+GO
sJSg8XVw67sN4wpBtEUcv6IjdJn1CD4cslX4Hsh4GTg=
`protect END_PROTECTED
