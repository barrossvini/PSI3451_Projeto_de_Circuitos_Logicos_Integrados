`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mExad+xMeEmJLgb7X32yzTq8+uAlA0V2nA1UIGy1Auot6zwH7hDDHl5F13jAXROG
GKpxbgi8uJvbPw7wXRblGLJtOvxdI/ZCPA1No5w/LJAELhPJh8ZMJ9p6s0KskTQr
Nv8gjNIUtpO/pBGYgmz6hdD5SliwRHb6H3z1/gD06Uyoaj097m/fp852ob/XntMl
bM0TCzfIoLherI/TWjPUsw4bjJHthJY38BDeHZfIezWmx3fHzydO7hW+ehhnAZlw
Y67BRp19PynoWBI2X6hlCessByjWZ+D1N8MbQsedKjKzgAy6AI0yutPugxrpZ+OK
YNhcRDoxfRVeRc199ihMVc63TZQfZQvTtFrpGkYMuH4IHOWo1asr+Fg7UC/RPtoW
b7MDfek7d7WLSGn+tFPI8xsR3e5xYwG0Rvh9j6M2vhPkhNKBOdqPPACepvTFFU5k
4JsgsWxPtGPmxpRZpbO7IbzOa5Cv5AuQvbG3tyoeMcu6dD/WV7C+akDMpIyUjjbl
/17wMNK9g7JOSPBgz4TLDByIha/qGn6lHW//ZIgbVfnViNdXIrAGHjl9I+3YVUQX
Tpg9J8V2Op8DZ4GC+piEvJTc0J5q8b2pTyn5Mc5QxGUWv1N9v8KIWJYkjps2ol0E
qwuB4THSBrXBkTUpFj2daSftPE5cZuQ+xDG742QORLbdNDv8XTSjE4QBTbnrlyq9
hKf7Wv/XPB9jotq99BoRYACdX5igay6YKc2jiSsFuGgLLGHFg3De4bAN7eW/JFgQ
W9lb+hemGKiEKHkW2lXSwDuv/D64XGrcC7r9wTzt8qUDokzWNLBuyLAELR5jEIh5
Xuf/GzwgxCTJ5dDk+Kug5jwvvQzDJoiiZMmA2VTC2Y7XNmivixmb2Fd0UE7gtF63
/rpGo9C0R9RfiwE/Cy+kQRC73XhjuUQpWPBJf7OvZvb9Incq7NFO6OZGxf3isSAx
Vid/N6NQ5MEUzsl/rWKeBT+fR9uzduRVbCuNCk7JewtpUXmOPrCIVtBx0NN9So5j
jFRdJ3giSeBpaQ5IXb0D3kMqqrAokTp1d5gSDCGGXsYQYLaWJ6PPZ2BqjXbh/4d/
T+E5H9mt4sa6SJdng609lNkLsbTjDTGpgV5EqRTtVQ+Q/9iXdab7cl0irJ/CwAba
kNJXlUY8mlDueF1qvh5edOaRESwBdLzAVI1veN7gHTy1zqy1MwnZB5U52K+KHXLG
965/dy+f7AbTuQGK5qxOyxw69FjVWQUrecbTL0DhWjIg5kCbVZ2dJjRkVZV4O17u
LsETPDrK2xEDwSrdbZkJMPdJqb/s//BNtDDS7q2aBywYONBqKrK/jxyKCMZi8pod
d2rb4V6P8F6luxDOgg8I/tBrZM6BfUGyvroa+QVctIv0QFt9YhI5eIuRtOvTwHHA
1yRysxXaa85BSqZdiGFPYLwHOXoaYr9WpVfdGpPJhtaNSTiUfVv1hUEWnelFKfns
kgS+CfF1IlymPSX7EvqFXQQnnBVkafHRPDQgajdoGSSVQsObXv9/nbilAvAHhoZ7
rk8k65C9jNwmuVsr6K0CaNbdlT7mao4DGgl0DPXIqNxYrz/58AWjfBicOJnwtbf7
5CDRTEghy3gC0KNT1S/XLsk6cIWXyO+dwXmTv9yRPopH8ssL+yuf7XwN33OLMxEB
If6CnXM7VAIn5eUzETrmhHQK4M9lb45AO+KM1CS2sNo3XBqPlRPjz1l1jCcr3Y+U
RNpa2E6VAPV0fjH8FdnmriFdGCFb8kUkdBEZUpxKWGchP+MCdSjdLy2GZTfiCr80
oIIEuSRPbOdsv9C6aACAnvJIIEfNWrNGCaE74GELPx/w9uMI4i3PHDcLTdqCUYf7
CMFMiU7DwBT5qDJdXlxrEwn2YVvrm2SSoX9Kk+ZFPXm0xBQq947chM3HuN4KXCR/
wGVm/oLfvQzoIuOx6MukLfy6ht9GSlcu/Q07MnZ0XY9t7xHwRtU2fnjtnFePjJGS
317aL6uxtfHqHPg0j4d0hzoeDuRx9CPADeyFsO9DHvjCQU3Q/1/Ielzk+gDkTm2g
75P4IhxnILaQtAE/2X3x8DixS07Ce2p5Mo25HAfZS6Jh7rf0p4Hde1EqE8V5zONJ
uVfP09JqBSMW4sa7SDvzOWFUDQA7tJQTZbf7vyxMrgEdmmKc9Om4FdjMDrW5y47b
vMq+cNJ205XwUgeAazicFZYxibxWcOzbkwt0yFzYJG9aJvFeMe5LSgNilXA4n9Sq
KGwAwRTcuuaRLZLODBhpoB/c+IygTCIRS7imGs192Og8SdTkUt4iQ3G+fKCJYE9b
BrYVkBh1CMYQxwKzwRP/xP6J1tq1m/CEnlRtrnJ1i9+qMH5oC+55Eg5lxv/C30oc
VngGK1cjBNvCwTWJhObB9Qq8SbZQeBGn7+xO/lIHVNCKvK3hfoMzxp2vyEGUdhwU
aMeGtFwxmoehPXyhMhsQEBFD6+Pyc+JyNDtuzZNrSorSodYz6DO5M7GVagtYWENX
kPkb7T/tzuX9M8jxcvXZx7TnMHaaTkwQEooKCevNyiHj+C5WiAZpiKab4zcVLuSQ
eeUz44QPIN1iuvdHIQnnv9mxAd23lO7kF7DC2ZJoVow5h8aFW4AV9e9zdC1PPwiO
8aYX4TLEN0NoEFHZqa2ubkKM8DbHY8c6cnBeH4PWw9RwrFzkLe5nfF8iYNn2YEN5
GSiO9CqTH/lgYUu88kp7k0ixmIW/YwMcQjVHAGniiOx1k0pPZrDSzXmmO8ATOSTz
6NiCCHWomr1y/fBaWNC3biY36Dog3H8zF3Y6BvMg9xd5ICx/GJezkw1MpTuBFv8t
pk+JMIZF37PoZ2h6Xjz027lHAw4MKO6gW3tZl83yHiVji2mVXzhYmhm9hdEAXBDN
NyRwV/NOXHNoke0I8hP7C/+nNcWrnEvKOI1vELmManle/D+newi9aofCMwvkoLR2
YpeHxAEiP3IPxhySzYp5q0Ap5g+vIj/XVNelroi0VAq75gjqkh+8i8TRenBA/ejO
+iVBz+aVwfdkcrefg9272pdjaeDCJZq8GYLYtpbXpAZduqzDV71Zbdqi8ycRSfSf
dxrGJb87I6s4HOZvR99YlpFIanLeNg6Pw2/BxtLkOoaBCO9OwG7rSGZflOuLJKFR
7gA8lhj8KQFQNZlpdAyakr4fnuAI56+CmzKB/VNpCTWe+9DA/RmadRYpbx+4aoQV
9wQrx1zcNvpCQP9oVYiKIvIcmTrNKXcZPHdoXCOKxyqwLqFbSCNshZDCZ5ldoL4J
aVnz3cuCgoQoCzcnWFFOm4m73arBCGZLNTdK/XSD9vDZYuWLYvrI/SoxyI0CWoSs
+XpW8dbbnX+TNVM3Dmc0vfrJ7e/uA2laHLfOLNrJsU9aVjyf7uqh12n1bZdjybGv
s2wjmRNDl1bPBh5wqCFN7md+4uo4J/XdNtz2gOOz7U2zn30tXttWhDynCFbGB0vU
bBdwZcUfx5Xy1hNik5wzI3QzRNBGlVydLEDs87ZtwN/7ptC1m0lV+lO4apcyrr/N
MRQZJAEQ1nDbVbNOMUOInWkXiuZVCmUeN/rTvMyktSwudrl/F0pGF7a/jD4XsT5E
GOGpYRi7ag/WrOYRFBn81EPqmYlerCyPzYlaqkbF7ZcEHxZYXcr60MVh6veX+cZJ
F2TGzB4fTlnCR+kFN5CuF3LLTVaJIutuMN7pQXMR2QkFWRg8OqUkCDMkkc68abNG
aKKkIq4bq8wLlIr72i3mUPQjvjfoG2J9fRWX/71W1hdfvzbXPh4DcGfYHw4ZjihL
dFkRI/CEx9p0fndZ3m2DJkbOBm46goyXhZ/NxLuKhf4qJGT3CwV1siymwZYIu40F
yK7MVOEEdEq1TshxW2h3julrxaiWkEF2b3Niqy1MHqV28BK92fQ7CjNr0jx/EPpS
zjE8AZPwC2yJm7ttSJ1/zlKop4Fa8xM+wcWOpIZ1lSNOyBNyvor2dV9tH+KpOexx
1K7x2PacIs7NrhS1zZQaeF53q9TwlPKa0De7fDVvSzJ7FQQvvUBgeIt1HVkzXmVh
sVyfvyzG1aKboT8oaNEsxPtq4oduVZDRZymIylX3yLU+Vg6/Hr7v10SyXREUXg3F
LUzBoDuVNrc3XfkBNyCQ41HspvoHfJd1Be5CBHUqi6docWZhtJb9AKrIBRT7lwJx
pm6RPI+8Fge+njW5W3ulnz+7EsrcPTSHOX3atQDMSRfLQ/8uHFc/SK7xIdgHB8at
rtHnmY6hJONKr6zgxNCuqs7Ia+qQaePGhxX5DIWNM7CQ1PTBZMXbxOJ1/TYShxLg
iMHLnTTOWcSTKwxtE3kEHVme5bYI2X00Z3bQLs2RnZxrmqWDfFtk3pF8uhFbBavm
YETaWZgrdFyeXeKrn1G2UYSsaqfhVzlXP08Xvv/tsOfVkUYj2kOtQzCo4jV/3VuA
lnZSOKN3NswstwjApu5cKeH2PSoyO/UkBQcqvybIWurKrVJivDthLeBXOqSzz8sH
X0xXmhGGBlVmVy71M0bS0FIkxx421EtL66iBr0OLfrHZmhjxVFlgxzntt2UEEf1Y
epRGDv+J/wwvCY9qvlPpNoUVBln/zqagjwo5SmftXhfVozktoyIlVB/0BBQfUJwA
shml3PGInwYNvWPQFNBVMPrxw9YqmCAYbA0QjuQJiTBjZCVxIlXwlo/zM6CGHCxs
oChIyuoDMI/ndfUgN65lZhCPL09m8mFwQ+/41YTnPhE8UPyKMJRWCF2gL6/dDT4J
oV0QgjCSf/pYO2U7oXBYY92RaADPwIh6kHdcejAFcZdUofVNz45Mt8vEbkfw7KZA
A/pjeAjMbOaqFvmt/DXfVzU1VuW5mTLIvuZFMsf+SYMiWsNvVHFH5esHtjJF6chm
hGZM8Zsd228a/Qoi03ilCzr18JsqfD6Zs0zVkiCBQiY64Njf+yNvZYksmF4mPTD3
DVNWUiMIK9i0cnr5lIZX6jnCKj5+aKGbr5oqzRRLry3JWUWhDQzAcqvF2IqJ4WTN
0IgjHSjhSinGv9ra7AKJK8MCAjGvswz6RTixoOLjiA9MxF/RQpGfAeby2oun4Jey
fIEpjWFlElC2OxgKBLZmpF0Rs0rzvBxRCC846i1plBLdv66Hwtipe/j5Esrpbk00
msMWv1jg0s8nzirh+yBrM9eVUP1gHrO7hKHC/Sif67Q3DgWmwVZi6zKnz452c/tU
FvC/3MvP+Q76izlW+8LTUSpp66TM4uq1//K6yydWJwgSCCy6y7x5tK0DXZDSWL1u
Nhpeq6/eOzFYGM7SVb54OXRRMqHoUk4RC9L6MUm8TjB0TG3EawF4rTripG9BDh8e
V6sS2xselKVbBGeXWfAFHYhQHrq6eSz6DRsgMR8ScKWa4TlNH05SFmlciAFfzo8O
TpfU3VXxUqvZxL1hUwLVCflF59XQjM4Oh6nn18Ytok8BIy9j57d9oWHaUSQIwXtV
ZON3tpesIsTqVx+A7Nb42JMzd/ff5CekIjhm1+HMNhgdSjKOBYBng86R4QGCm8Mh
aiWLZ371E9kxaqMFWbq35c2yO3p6rjgkEoDcM1pso0rhpianQWOYZTC69fnoK22E
lWUr84OzDYq4ul29C7AGgP7OYJOb78OVa6MDxM6KpWuTsZV9MUakfTyBpcYL0ScZ
CHK0g2UkJEUNemcyiAyTnMBXrjwVf3VS0RGStWOSlj2HZAteILQZRpC3lSe2bOb/
Gh4SaOInWpFTPmY/4ksfisac0gqZ8he47NjwXqywG2RYPRxIEOmMvEwgJyIM4cs0
CeWrv9ZCDFnTcsTEv8hOm4enb27b47TSMhmcf2uknjS+19X+bwO0KYldF9yMmMLO
eEe5Ve5szKXzdMemskuwNENjVOn/x9j2U8xqkf7nVbjGIHfPFGwtR3B0SZSXnz2l
cjmvBYx86bMnCDRdA7zdj5RS3wP9IfXdIpz7yIQQ9aoqr7FsczAEWcU+oPEABAs0
+ixZZsY+Ala5vE5oRYLDuiLfokor7/Fv8CuzXjF+UzxLlPX2jBFthA0svpu7AdOx
7sMQZbiYQK7JuA2ecM5OotATHmUZxP0OHTiENcNXxnr2uQ1EnmdnLWr3Cc8n08jY
z9avJfZSJsLrS0San8htzb8QXwLMv8xCD9d1xBCg70pmL9Jy1EbeunsgDAATSVJg
MfjmMAGQn7HGvqF/VvxQhjhWYUwf7VmkU9coiZNQU8VhGge6VQfdxEcgkNbVasbr
Wqu7LX1LtbjTCKl5EZSmul0bosgx07sN98qQJXl52r82HgoOwL5PWiJcpxFr0NdK
s26iXN5ozC9umeZuIv2NcelBYlPgYItT4s3XuxYVHjqGm0LAdSsAk6HxwI5SQWtt
u4Ix2XpjCdRh5nCPngW/zcMeCMyr/0SiLu9UFz45iqXywZOX5sMYmmh3zSvsffkC
rhlyaTDomWgOedYebQhVxSUgrZhDObhZdbozwhq5a2s1VTg+qNj10hliehe7Lb5o
WfDNcKkFd9WGiUIR033RTL3C3yBCY9UqR1FHcfoIG+kMpcTFLpJHKwbgDqGhFb0L
ByXwS9Ai9CUyimeyiTlPwUWqDoxlXipS5+DTKVUJQfQbwoEm+Zxm7KDhB8dcXwgg
FZAcMX2Dq3YQNBPKvyoAWSrtGByFweo3LEFLAIWtLLHz7OWaM8F/OGBhHW8lUhX4
aajIfE6bEXJ0CnG3MF/uRiC0PU2cK6pNVR+6PZumROsq3GkToqIRPh2zxkl0ZTsJ
Vik0YiZeG59tbB0NKxD7J9Rt2j/lGNQez7SSLUa0jq2LsEkfTvaOuYb9fCBjHbGZ
61dOh4PbAQmKOJ7z8P/eyv55nUaJqGmw1CvA96AkJouLMu0u2VX4hl1VySR7ltCN
bIelfE75Uwe7cYunaoxahCs+G7HA3DSmt1AjabQYJ4whm+fUKun0icmfxN5YfQtT
y1oKBVM1iz9Hh4B9liaGDXgG+ER1ziZFTvHH8yy34UlXPcUnRdTvr2Updfs1Iiy6
HHUCBsyGvsnxjc2vhTurT5Tyll5l/h4GLzUlpopvuZVeiXAQVc/k5BYGz6PWwVl7
Pu7C8kZKSmOGGUCmSd0sPJanHDlVNQGKfVwydNnjMtzngMSv9BKHS3omCTvJkVcg
VpzDG8GCpEuON9fwQ6Cdnagoi9o3EVqCAr7OVe+/o6ifAgmbZWFAE0HaEUL2awNx
ABhScROgawR4IIgNWNDLXZD84qFTRVh9hu4564ChPkK22Tr3q+SMRIbzzbqEXB2l
6jQXHSbVfsUW6DRDRvjYIHN/rmvjq4FlleA8qJnKM+AZrG/PuFNr0oL86giBHXx8
WkFZ1HHPaxzHlMOJhbbgTcNk2kU6OuVImSnccT2btL9FMURRejPYLLpFPVjQQHXl
ADMT47IWT5FFG4vrSQPGVKou//wP1PBM5mAfkebs6ZLyIxREduMfZJP/nJgkNVpp
azfhckkGpQuxE80xrp278pbD7SgY8h2pXBeRWnaxycYCEv0+cYn3NF+Ef4AHAXn+
f/VFjg15ONtVNQ0Zhh2N5zfo7xTF9BbZqOfiW/QPBKgaciXKb49SfkJ1Af0PALlg
wLNFGLUGaFBzq8zBqlCWndUsYh77seB8IVtdFRjCfGY1TKs2gq8InxVfCmdl9/Nl
buINERP6J096Cwzj0+t0cA16hxTRdTOLqqqawNbY22Myk3JxPpn4ns3MLE/SvVah
eljmCiXGredIXM3D2Ng/7GDYGQAzPvE6f838d+Lfb1BdKBBm2ZM0CfcWDlRr0On5
VkjPnIGaDgoW188tOplo5Tm2+6PkyzadyXFCn3icImDPQcWeeBBeY0wfqQe/Bizy
F9NkSLuMpCHbgyVQb+/6b3SXoGfa5GLNjHPJ9Z3w6prLiplhGcfkG5+W0lrRgBY/
2mGhAFUKR0Gj3WUOoR+COdVnO5EVngzoIN4lfXwgp0+7/morhOzKMPjQk/+g5Ej5
c/xdyVptJqBHOU+pd2qj5DixhruIK6YSMltsZ3L6O2O8FVswSHsBGjeiuzbSygYD
jmMCsWplLSt/aRjGzVFKte3MW/F3OUCoB7awozSSw4NeNQiQDkl5GT+dCQJw4egz
br/RlhZdbXPpOBdM+ldrsBzfP4UUL8CFnRFb69At/Ah8bttJ7C9vFgbJFLLrBTOc
hmOtajegTz6//5G3psXK1+d4xvj78SaJB5lWVmwIpuMp7HPmf5Y+nb6h8jwss8X3
tvnK17TRaN7HNATtbvVsKnc7eH6LVJ/brzYIM6qNZn2flwKO+h5T77s1NdBrX/5p
6i4W3vMx9QcmR2nbPbY7iOhVzufXe6FqNLPzO7ZyAODqi5X9RUQaBK569m8q7RoU
YWsukeT1RVY7UQbLSuT+xfotDo6DVdStIR9yMKYgTvTfV+dTQ/fJEEs7RsbU3rsq
0MBiBE4cNWfbluq6yQJQLrFeKrRNixlSmHAKM6L8P/0BddQdPjyUFPMHxj7YdDVc
xgVrkTz2Qb46YCBpIdWobr68RvYhsWhfR9Ri1ZYE6MdKNku0pyTPdj1Ej1ADLbvL
MLcokOXy1d2bOW3nutdE/WsLAi6gDB/mWcEZJxx1WikbYgcW+xntDxq8OBiCnkrd
Ux5Q6r9bM9Fpa2irVQpIzYOw3WwOst6T/N31IIZhkjRvKQ5JUfBxn7XZb+5EGBmk
Dz8Q7t1URrus5PVfUXJe2YLiuTe0/3miARLYJhxSi+JRXoQkoAbfCPYMs/7tQj5l
gCKD0FusTZvUrlw1ZEaDeK4SyOGw2Obqh6lDVT4IMHgik5oopZvfF3PUjuVBGKPM
UqzWba2u2QsufJ4IjPmbFFMxB0eX49ea6jXvPP5Vd444ylP+mThsNKiUQcyDSVyW
Te9unmnc3o7bEqJOo4K8td6xj0CcONE6ng3de446RVVskJHmSPFGAqnIdTy0tsk9
QMmmPZwWY8+Oyp8JXw1RU4dm631kM5lQSsHh7vsPOUizLFWkBMTYG9xAFb2geiN+
rG6tuycqGTN0vMSja49Np1+d0IROVkNsYcgLEusTXSokmvCu1OMb/tip+olfjtK3
B9W3poWOznUoid4cdxb68kSRt2peoxxL8puSKHNM6gKu+gbBLffATFDt1jprP8ko
5OBYxFg9s3ZULo0yTfI8fhUCWwWrFAPPniLY83cYc/AAXMd0gntx6mOLFSxKg9Qd
6ilYhjVilkwE7Gcd7tELO+n2To4o+DpcvBa0pe2ao7/9CGok5LpJdC5ZTgUw00do
/SRN4FWxtlFtt1IVrayVLd2h8knUgho8vERVICJEhE35J1m69x2Le82yPmYQ+kqX
wyYxsM/wdhuupiQ0vtR7rj17sRzdUrfLsipM3SsdtPRV+lyOFGQmLooBp39DvzWw
QMs1JtBbz/uqVhZOlXZv2tCgx5wE7cL30cOhx+KekLIQsC/PyHGuCvyDvi0h/DkQ
PhCIYeYE2E1229T4mffWurx018jnJgipQGjCLjzEFebKNzBUFxNcPBxH+VAPgC5M
x41nimLlcb6CbB0X/roYnuV/g5xtrZ7FtmVUOZ/j1Jme021YxK0vYg9BgPOSMS8s
gtPffItGcHXEJ2IfWZP8iFnj8BE+z/M2sKLeHBpBuBfQcpc44ECcscvUKcM7ehlg
gDP69PzymwxMdikVRmXYAUlSdwBw0WrJLjoNJEb6WyZ+OgU9LHN84SoAlQCA8WUb
gDCQ/YD72yTP7euXTSxS92Z9p4DHabRxCM7OWDhepHx1+au/r/+S6vM68UjxcgKR
wZv0wOTh310x4g/uG4eFPUNPk0KsPB5+vZWSuu5Q727SOXTPOgsd7/+PDI0SAkji
xjb3sQwiUsA9UEufTf6+UzwuvyyR/Al7bPnxPmp7A8mZMnmambBck/NcIDnHAo18
Dtm/GXtxTO0NFvS5dELAaFdlSRuDF27QronDaJhPcXATSUlaeE5xLXllZvyFT5rn
lKzQtopUovCdDAzZrDZphFHwqi4mT6L1WdqlFeHCAh5zqgP9CF7mNxaX6GDpNeA4
eMbmvwDJO9n3VcHE62J8xpaEMvgw1xaj1sHiM1t2yfBI51oFVTBPu9iQkk2zV5HI
uIUcOtKWbeALi/2cwi9IRyhAQ78C1NUIPtc54+mw//8yIetySp9usfWiQuyC+5Sb
V3cxzrd7yepi3xfsQfopoNBgk8ftjShf06ygEETP+bu7FBGekekyw7py9TD1UDjd
jFgSkMx3csuWX2NO2ONEXDkljmZFC1sTuDcSPNebCiESWtsOqEMu1M+WMGXkFpBl
vk/hUukVTyxRMeUtYxUg6IOMKa1i0tRU+ZSCyT0SVZCkS35CHD17Kao75KRdY5wC
nU8Xe3KUVYvEieehyI2xQd1hKPsOYbvgXKYccYcUXoCaf6CWLiXsNngFCYhTDTVv
KhYBbiifE9IDe8cc0az3irj6/0iVpgGl18Kor3BMwEDCunD9N7xE837HFuF7zTas
jvv3bm7eUyyEqDX3r/SGj3xkvL+jRAfsJrJNri2Cq4g7WM/swKOddC8tF8UhO28L
4wI8yC++RvFXQw1fMxsKngxM5ijXzZl4ylPcAkF163+p/cuiFqq6XcdYsFPbBSsS
paI7VjASQ5bpmrSbSUF/cQeU8kkDAgqmhVrNpaeMrBS504oYZgSPP2dximYIquVe
2LQIeTpVvS+iNvIlfR4DhMlj59Zrir5eNTP2AXDVbsWru9KVjSaWoohog56CiIER
zMX/Uljx6BKBos5d8YteRSMAse1jdFSteY9CIAX+Ynr9rq/vHikebIykLAr0wIiS
Eie+Cviv4DPZyfzdUpu8y0vuCIekj/8cwOAYBJZYOKVAAiazb3vBG+SgNMuM4pzf
DndsH6meZf/XRwsIY4g1it7llbPD6I8pENRyNu2TwwYutMXE3ekTtWXiKR9KIHja
AEh8ZiH+FFV1UQ1nVLm6E7FvJ9jBYSVs1H4aU04wzHodMgC3zgRspldVuygowr4F
9JtX4RsK3p05tUhEeTfED1XyWBIkW2ut6kVIKQY8Q2UYSBHjTFgW4l92RBSAvknt
ffeMIsNQD6/YHMVLeq0LqrWKOTfb7yVocZBP66WeOSVXuAMgwakWD1ecaL5lnfDP
PkUH1dn/3EzXNPdPwr0Nlbo13Ji2nTD6+b2RH5NbDoHJCxFhACKnGb5wf4ew0LkG
LY2gifkQOyuV+UweaCbjhqLvhytYa3wrB2g3fEjh/dBpG/7/CafSwyQCUwlBiqbw
U8czU+/n6Xuh2xEixXrtyrj5dPNteY5OO+go/z0cpT8y7CE0J+sVXJXNtcVRPvir
HrxFOZZonimyUaVloSWpCTzbQoFesRzz3Q9VDvnvFSB1OqL+wqUeA+9tSBlgfEL5
0YOQCrRXJU75dy8tMX7Rr1UYvVT7U30+/psYZwsbzJj1wYvfWM9Z6DgAYWwupIAb
ykttIVIy0gNjnptbn+JdiGASOz0hA5J6mwYRqG5p8pnclYhsaOCd1X7cqmh/Z1pJ
+4rik+hamEmWNJxnZFgtYa8mFernExlPTDXOguuWzlNToncGgBG9gGr7oZJXv9Qk
2oxXIa8dr/5nTjmojCPJYg07HfHivO6lgnCjciLYlKqiBAINjXTo8DNT69xDu6za
c8EPMfXHT4aG6YegmyHYOxkxwK9gD4r+r9yaEVV14qQ0F3M9ZZKInhRo0i7DxmVw
Q7IRwF7ZXKzBZAibnfqZlyXQ+Aj7RGTJD6VCGhfc0JJJIpL0oNrFU3H0JywBCokB
gpSkr/7JUgDn+dyH3rm/nIxd1GiWZ5K6/SkK9Nw5dg+u/PUh8wMmffaJgpQ2dSj+
hyvKxpsULwcx8AJIL37HDQTak4fZAfSuCD7kdR8uek4Dhk6TuCokaKIK8zmLwALx
5cdJ0nO66dTdjw5fHh3HkUdFQM9zYp7lG1g3EbsgICW9DFh1dQgFytdg5jHLM6im
Wv1tFBDCaUsnwcxB5QSJaiQLjNfF0SqvDznylarmsI1z9f+06XjoTNmRKCbNSm/s
OhSiHq9NOjLU/TllQl/cG/5Bt5VfAzY+JY22bsymUO4td1ZkR7DAaUxUPRpEHxGs
XvEwy9GbuVA+CwLTMg9ujLn8gETWOF9IIKduQclfATo541juU7leLUA0Lx/nG8V0
6va82GL7vUycLns6AEj2W4IhWVBjpFK9SEIM70hUp7kDvWTiwLSH72jfOc5PHNOE
aSEY6DmvnKKZ3ATHnsMy/ZqY3oSSGiik6sPcXFerpqPg+rtFjDx8jgh0BDL0FDt3
/gMsOwm7OzYqNQzprqVpf5pgwf5mIdKm3sFgGNemuKFhdkEG8IMpLhwJcSSh6MxF
yzdubBt0LieNqaYt5bEKGRe/fM6c3VuvbtZTdjzXZzZ+rbfCOzMZjmRMZxtqxevy
I0hsbKjbolKINKWiyCxA9xyxe2k4/mBA2UCDCTNqT3jmrI+i22DXerFvePsKGB42
bMrPEABXxWDE7H3rkUZqfTggoPnH12imvzqUUIEYU8FwN77roQZkYT6WItACsL49
9MxCyblaooVTYEyRuUzRarJWg3r2ux+4UNPK0G0fxDxHCtiV9mxw1kEuBsDvb5do
RcHOCYGWJ1bCUo2d9vNtbscFHYvTvXwxhBbUlcZ3yJrav7Wgs3iCKyRTUWMeZQiy
L39b8BtUhXBvkSnfazzeV0OwFdtoE66tEOsCQEJXmhL4NG5z8xI3JV3ExVZ2vc5k
PU3EZdSnubhOjL3Hy8bpAk/KpSTNWMoDrM2F8JuNZ/ppjwgbKwRJIANnjUomPLC+
4Kd0Tcyq8ePEyW4eG/wrqOmF0Pb7CIYYSffe1mj3SMeBRDEaxYqI/DwNhYQHI5Eb
956701Rw7FaYgdaS2NUf7iaOP2B39Dbcevb7lfbD+y21WZAYaLioiWH0SSmYd2Yc
20Qe/yfp+7hb2aitTLl+rjnvaPVkwarJDSAmuIBv9Rxfqcf2rptCLOVK9SysGjFO
uqVMvqpJ+l8gJbmuPdanrBrkoYUVZtfeQOi+w9aWzoRKyMiA+FJQGRW/p8Ds5pJD
lh0G84OUPZfgz4wVuRk8yYq+B66rVqQ0Ruf9I2kwq9xiuKrj48Nt1/rFXJS/DZgD
htHt/CepWVe4DH7sOHqO5aEF3cyM9n4W2WXRnytoTgfNmgahTNiHu84TMUaWMqMd
U1oNYogq+QzfQMGKnuk2TnjO0gwnHwfKNI/Kt3AILmCE0jv0ScIrToue7q/gZ4Te
ZTvDEmpqFsf5itDLy8R5B+Bz0KEIylpuwdYCd6LZPoblI95Nz8A3pJwk0GkVG8K5
WMJ3WWu0SgMLd1wPD42opRyCAmZGuyErtyPM1ffEbGlSWMz/DOJ4SRrzbg/d+y4C
9CFnE6kF7IQZ1POhW16HElIn2FyQM66252Z+JTormgEi4xIy5W8AqE3BcLHrYrjg
/cVrRh/BRq8yC9YJPEklOHafa2a3zO0EBmbC2JgfVOPZOQEdL3WVSukj1dHfA9Vr
q+bLehrYUTWLZAQp3f9P13gMBUY4h+HP+SUJrSeYPpkV81KC8/o2nygoied5H1wu
AIzVdfKsvuoSZ9BeHSe/xPZqcIgysL1+gzw0cxzk+vPnTaM9tmgdM8a9yA7WAxsd
hdzJf0Upo9aA/GU/HzP3A+YfkUAVO7PT5x8k5k0bh3IVPB3Cu8llusjYaaKl37sF
XpWhNSgv7LRxavPOYG/JvWeEVohZnJklLAUFDHyEzIMS7GaVXWLGg2NCOZ9S1Sxe
191xutqs9dbts9F6pplEzHC748FABwwy0xK1a/whQLzo5XtlvMAsPSUjPFoM7Bn+
j4Eujw45sYRnDSDJzQLFHKKXZHW93OpZoBHfefuv3gIvir8aQWoK9vg4K502Tmnm
CecjTr297+JMLQxwHvnL/Ms54Ca18x5BIebzsG+o0sSq3+bY8OYCwG1rt69GSjiM
0SJvnmagHEyeidPGw9UcRaQ2rEy1ROH8rsZ18P1nhCMkW59fC5Pw3rGtfnXxc4YL
WiGwd0lcCjNOqkUrtdguP7+kk5HWjNC7jU+TYi0lrleA4rUY4+yGe9rv6riweXV0
Wn6EGVIMD6dayUD5NdyH0kVVLVOPpcSFDINicrcWMqwmDWhqWbbq10Rwu/IBAk+0
IRi9eTgu8/e6QGoU7k7t0gDgwoLBETKZZweg7SswxHsu44lCw+DBQREZRkj3c+c7
qijMdnvk7KNXznEL9aSVEICELuZuLXXGRuhhj+q7ZyKZ6+29IFGVVuUrNWTAg3sR
5Fx9oSRrCJDj9ZPMKdEgp0pvaKi+i0yORGkYAFEu7L/MoKKvRep1wXgbprqZNR3Y
O8pWg6P00HQQ1b6t3XzAUIoYYY4zUfUUfMf4dw1ODy/QbnmkQ/VMlhP1qBU4esg4
2/G4He21UpEPQLvSCNH4PNQw9aisTV4S4la3qIF69EpZlRsvcYcDanfTBThSfAmq
KFQfCY7MFX3SdRPTppH7G55/VPYUi5Uw0E3PntDaa1qObgF+W81/rOhPMSIUw9is
ktQe9C5AQYxQ8q09ISaKw4Q4l7YJg0NEhoMajK8O2MwjbDVvAVwtiOFs6/iNug6r
FqxWbyrY+1P8yRDuLUmNx7XkXOMHD7+n51TH6lbysRhWCg1kk1uZ2Hq3sO9ybLgD
FQFZ36+LxBWG50OoUSu4K6/RsIbclAXZIHtB4GJKNJFT6ivGLD+L74rTgXFr8C04
BxobDTja7SWrj30kyoc30rcYmniXKBtvAfHK4xmgxXIQmb6otx7UZm+J+qHeavte
zHkF7gHHqrHDbqr8pHGItqXT5EhXg6KfhcELTQN82Ua2FsJFZZVB6+8SyFGWT0dN
19namNygDE2kxZpfiLNxjMnlknCTVpAneyK4thU8mg0XThkL1K7Uqgf3DWe8JauY
p7OC3TqBKSHB6XGM0irnqQeNu60uf6gl9GPDVG3wTo8pkO1ZxUujFiMPUrWpfmSL
ErYfI7rtw+LehhRBbb926H6Lb2wVZox7O3DJwoGQ+IX6KdJAJ40tnF94vAKHdPqE
flE2zEb/KOuNhj968J5vyBSiJstSlTJnJoFVJI95g8FAhyML4xIT64Oa3S5/W5Ry
pECafuMSylaafOKr3KUL3xSY39hN5U271Ondls+MIJcwFpU6G/YpNAINGYOXcYzQ
qHVFnUgNz6su6rg67x78ACoxm06cnCapYyRd1xnO5LW5jsuRO7o5CA9CmnlCL/9c
gZXTBDMPGmpq5namj4bTX6s2uxr8zpNHARm6VXXNarSnSwm9hDR3hnRHjN+8A/jZ
aikrGcy9FjBuVVlhUwZTfIZ2yffl5QBp9r4OLkegHPv6qVCeerbOveOnmaNen+cY
MjAA8+RX95X0KwfQZWDW6NvsLXsv5KCXqLlZQYsJdg6ZuYWNIAzx5GXI59DCZLL6
/K2Ws2HAscbzpyh7pTwjwyho0Y5CIs/VKguixgQp/P7ME3VQSstrxrnk4ZtqC2td
0bCOd1gZB+g7Gx7AnjS8vr9tO0ObMd28nbfnkHgtIbZ6UGGyJeFx4XEoj3bOLEpr
4/Eiq3rqz7TWfcKD5F8UQfQIUXvSNa/c5Vz3DYENZYRjRb5faVK+M9yxhvyLG+zJ
QNxaOIyd1VW9IeYmPLDaRnmT+rz+fa2fw+GvNqbrjF9j5jZX0oNoi5Xc7DAwYmgr
Z1Jq8SLhtlrUWvnsLVSPZ8dty3Pb5crbSkCW5qjOp0jXpMAv1fperl9aeSLXX0QS
fDxw6pUgmzNpdX/bvfBYfxBIjY7kktaJKKtXhTTdbpHB6fF5Zv7BKUdkH7sGAP4e
qbmmS+A6wdnU16C0/ci8hI1T6jQLvSADOElngZ0uJ551JxXe4CKIn4djSiybYpo3
D9S/csapWUvyVO8rxGnjedradhOH7+sdoPQsjn3sv+Ou8kFP2o4Wrcz6DBlDwCHT
aeokAAqNbHO9UYiOQSopre95PpOrdDadR1W4+snQiCcn60djbzeQYoB1mfsLT4Fo
IBkh/b7eqnenIC+Dj+Pc/1uxvm6EFxTMPdYKEeWnUKnW2qSr9BKSkTBq2zy7fo7V
Gpy5fwUooLC32rK4zIr4iRS5qsAK6b5kXx2PU8ozVn1CNvyac5jAS4HxznpYtp45
IoZhkhMvvepBUbpUAccsKUZd2wXd/nmaBUa8mNA9w64kTxxuvoEXalL5Oag8hsjV
I4oRbQR9ezgjrY8nwTDqcewC20MymtD9PqfwMhMpVOi7L/BRB1HGVpVsKXDic1Xs
knpXwtD2UvCxdxDZM6erF9kqWCt5+GCXNhOzyIa6EOqnoEnsjFpaxm0R3RmeQbsu
nmk2FDHBhfCcN9s9awypvIvd5ZO+fK+Eej9XMG19EYPWporQTyt2sQ7JvG6Yfsvd
EQj8xlgrN/MYWbQ6UTrcBiMYMb8U/ZuhS3WmDdAhfQD3FcYeBz71nIv+wZUCLtqf
kE1Wj7hrnlnm68E09CGw/Jq8NrAsCVkZsrqzihqCtJy0VMorLAnh9tLc7Ivl9JPk
qSQoY6zPeoMlQsMj9tK9aLb0o7FIxE1zRsmM4IStP7DIVDOK7q9tOKOVULt06T6J
xXCYuDQmMHY4V0e8oOBEUYVXksa6fo3YumzhA0tmkVlOt6+WTnd9USPmcY45ERLh
z9zjojGssSi6MF6lfvJ/Irm5CNo/+a/9Z3j1cxhb5ja/d1UWfCkQ70Nj/mfn3qsR
vNLK8oLA1mi9T9Wf7j7V2ZNLRYvge+rJq9jyrs1RyVdA1etmzlqyfeOuxh8SQX8B
9yxzXHWfPNwyIsrDQbzDeNUCAYKe5BZPKAtVudzMN5ktJjAlsjeT/70Mu7si7QZe
p/IhzCCb7lKkaQ6/tFIsk7MiZczvtSZHA9HGDx+u7zr0nt7us33cx+QVBoR/e233
7TFncOmBlJexa5rbvZ5n/qMTxpKbIpiLCBZHEQA1mYTUKT5Fn4Vhfd0p2hYUEdZt
49P6xoXAP6uUhD06NyJhCczke3+thfhRau+zzGBJds5KHJ7igYt9VJbu7Uo0O5mx
7/B2krBQRLsxXGRzBldCEXRqzOzDHBfRktp95PKnLul9uXpOJZnG06iOh2SvzJ/0
ZFmm5tNWKqBhTtVPbj6RfBv4XBTO7DD/fzOI2zHi4sebtlT395IIwi3YR7dinr9s
gACj7aPRGEy/pF7ySOdFSrhx8EoewreN/IR9bOsmvBQB99mjyVam1KgnHDKwLE5A
/rtiY2iO6FFsw6hMHRkTBacNailsGdDreSTXiq5FpEhgNjo561FSNNFfjtpXQeXH
VcOCcJBgghCMnlNbU7hvLIONoBrOnLForpB3sQeJ0Gg4lhu7rxYf8sbd5UOWsqs8
gf9d+qZ8r4D87WjigLj3aaRl3l2LXcAbqgDB8c59J7CRPH9kNq05ksg86466DjfV
ZN5cszbWmBY2HMwXskw4afIWnnuJpf2/i2i1nWO3lArSLzDa3vThsaAdNlO6Jk0z
h3Dr2AlmVw/JMB/eF4CbASSwMphqUKeuaWgLGWJSGkhHJHS5HuBBJLQ5UrCaPwTy
TsaV9ou+j0PMYYc/w6oxfuyDzPqoQh3SErHHMMdchj/R4MPmOVg9hBPGckwH3AoV
ydZ+PgWBvKhUxVUDJE+NWtqXLaeEMl+XnxCHrPRiI95BYeTcsIDeUbXN5UVRzwwP
rJleQIi8bAPxBAXsjOb/bBW9tqXPBkwTs85uIY3wu9Uhh2NS/9Vw1NHNQDag//us
23SzY6DoHMSBMjYcvqqLnVgANXY59n7pAMEIDDrmcff6a5jICiCP096IPA7pUudc
xH18ybpnndvvEuNrl2QlEhoyP+qw7ReEhJIKmaLsnqNbcjRqdCon1jMwM7rsSSvn
rJ2KttesBnRXDu2X7bd1N3qY0z5HQVQ9VAK9uPPjIgG7RmysO6LLJGZmqwoXKYFn
VOvw9OVVaEYhbU4GKPnG73OjIZ7UGdJUQdh1fCudHrm/rPtukBQl2ZB//OKURILa
bp7cTsKHMEfbshkwqPaCTDZq/vVsdDROCEn+yBfIm6h3NdWYkA4MzIW1Yqzwbf8w
lUVDcimAhR3pl1/SwA+IkU1YGVBIXscRBtJvtFIyWadrQm8kSXTAMHZdeIY42S5j
Sd+VndjqqG/ghLjXN17dAxoIlMJAMHC1UTysom5RbtRsrkQTgBwF/c0j/OI/oNRe
jzQDKqgCdtOdsm985LA1Kc54RneVkX1xd2ODEd8emyQd5zKYElWRHilkWlZiUF5Y
wo1VvYVbwis1xOwsT+PgWysIho7hf8tCqudrs4swCrD1sq9jv+7yh5FvtRLk4uwr
vEWTrRdBXkuKK4ZVj4/S/djS6SKg2AnTPGwhkR7hbW28lsxTIt/wlqBqaf4tFSiu
yhcESsQIB+CTyxx9b8K81t1lKsMWeoYbTUgjrLtDG1qRbXNdNnyN3041Kl1wPhbY
kycjjj7Meu/ECaxSNzhUabuiui19emf3Zx0e9fCtLJRvkjs5y3+mZsazDZB+gmkH
vtmxaUafzIUeO4dzxu9F1VUwLtwe6nCCXfwpdAgaimD9OTJ4bDEav89hRogoiXi5
Yk/1wtTunHGETxypuwtLGMqfEbXNMXUoG1QHvavLduVfSQQmz7cWMCv0nVcIadze
5jJoTWg1O8T+TUHOK5gyRrBdaK5X/e91loXQn6vtYtV6ulmWK98NpJ1qoxB4z1xI
NUe245ybNp45a8cGkgZJipbUug3kMF8jT/ZeoJbh9jbIIIYyqTN6Yyq0aetSemXs
7cGocNXELrtQY7Z6zxEUt/sFbGEb0QPobq/ubuPcnOD3AulnOfXm+AFzv0jUwym2
KHymbScRzpYyw39OK3CkcWNB7kgInt5Xwa6d8IvLb+WQsMsCoSypywHFOhFlnrQ3
2V1CkqeNYNhSuDHTavkn2vZG+y+s+AJvl4oEv0p+YmWFSz6wJaCsoeH2PkY5NmW/
BC8/PEXxGK2SDjtyEVymudmPljCBgYD7jgxkystKJLTYp72De5E/6t6TEWQEijT1
/BgJlgrLwJKSdOluz7EYYsRw34rl/PEMdXb3mcdMwfZuGrTNhXEO0oInb4Oko09X
wzXQ7q2t4nJKniTrrxaIdv0Ccc3n6o+0+IGurE2bXjqP/YM3/9uV1in5W5ovKQqQ
Yf27drie5GXwR0e0enHUUWBUTx/Gcr21HFnH6zRnuzppI8/ClBFedP2FBJkMNt04
Ta3Pt7pUNjqulZdXBQQtOP/tTiEuKCQlLgf9dPMObBF2XRgbZ81c2uNLK9vgdwTA
5Aq5HMK90B1GF9f7c5ZnskMGa2Vj8AO04mV0wuxeG4mouSG56xOftcUXgMFC0tIO
wSDUbddIx+J1Wlj28uam1pcMkXzln7ERvuI0Jh+c0WKyptU3NMwhN4EX0s8+vP5J
afkOVJIGp2CA8dMCKs7ogAyQ0O22tamMbBL/Pcsdfpa5FzdOR+IsQnhgrMFSMiG8
7WfjKUdAzlHQ9MXekj7puWAukd/u/hlt0sxL+vd30tqT7rIP3zOTQPsc32zPqFjk
aDbRfnL6/VI0p+2f6M/mcHxpWKBJWOQbvHQuxUj2fpV7x3SXIkhtmhd245tgklcm
wOKaAAQABKMkQmWOP32HWhQ7gpINGS4V8uFzs0Fz6ig31Cn+DO47UH4MWUjRl/du
Fd1GuS2DY+Ajs9QPYbkgFP/W9vCFLJYjenI+RKM5+YCcoO7VR2P5foSFkJ4VRJXE
2SHbaJzRWNLklgvJBPb1JROPwTZ8rr6c3bBnv1H1icf7d3ofE2s8ei+mPUjo0MES
lEwntYYL/LOhFFwBbvG7aBGX9cI7Y3oK5uSm3MfAP8j9m9CDrt5MjzBtTxsNSrr+
8VJZKzWXreVM8Vix1I5oIgUfLPfOs2Hno2yC+KQiMe9ypijXOjpldHoZ6PBz3Rt+
3BAoKMkzaFPsJ8zXFcbFpY2Pxmpdv1EiKAxGV+tGPp4vHJTiTso+Fblmrm0qgwjf
llAqKlZ/4nDLXs9dwUD2kBRQuKrEtZGioUSZhey9oF2v2Uc0s32Na+FHST4elYgF
2LRso8AgYlUgHqsM6tXmzje7qZ1fGXmZl5C5AoymHAISI4gvi3JPohhf1C0mO1oU
OdRWL6hFkmvF3zDjJeboCSFmXME5FBLSECduLA5Ln+QWFkBRiIjYMTdyB9/clfDt
j8STgHO52ljAZ44ccSnnggyQPtus3sY69+jTFU8lqxOW2Ox0FgFEOA43bEK5dKdf
D0JHZYw4yCgX7/wU2gI7QRGgrJo1c04XvnAZAUvXTXNFzQ4lCdGZQnE2yJDn2IlL
1s13nxAQ7H3iN24YpQGgRYC4OdOckeb3CHZo07gExYh5nSa5aI3dgkBQ6sIz9six
jviJF7M6NfmyZgDNYq3QE9mtNNe6ktn4scmFD7AYbIw5p7kiYoBh8Pyj/7iRWh4e
E1ozfkAyoAB/Qmw+tGbYkEuOULUqpUP25btfw7YEW34duWNVMIfI08iiXqQ8m9KI
9CnCOv5Ys0LYLQ31zdBgtOrlpbPyM0NBjKS2gi7pEOUWuN5CWBOBHm6VSfak1ihY
s3mp32J4JgxINVavUy1nMC0Dw7BWqfzaAHVv+LQFkx7oxRTzzoozCXkxNpRkgvVs
PXPBNkb21IN+ATKyKn4AaU1jbhuqiP0IdNFa0ekgbpDhlO8BfD4yRd/KhOYWiMd9
yb8AT+K65s/E1vUq3f3nwkkCtCXquwiwy/lA7Vp63mOKbpwCmPvoysC23HkJ/1w9
/gbvunyFZOY2ttyYw8HguAOwatMLIkgfJ3ciFwsoqX5npEljIhfyvDbMHgsi8Z49
MkSdB3Ip10cdv84MnHuszldWmNssJwfsW/jb5RHvsM61vVr0yrseUqK3CLAPDRFg
cL3E7wvGzJT4aQvGzqrSKXk/AfEX48vEokVsi9hY6nIdkKU3Thr2gcYiaWyFJSJ7
4c4whlMndt1deGS4UrYVgK5JPVXMi13vJiXow8R4LUtjUwDfItYDV+6ykNxb0BAj
QOqHykm3Sn1Wkl+IdNJxgWZxfXHzsebdirYugIbbAPgahUNhjTFp51gNxqiica9y
eZrYO+PQLvM5xm+q2PdXiyDzJW7SGGw6pdDkGWqbBtiS6kRjtGNFxf76acdh8HcW
iRJozNINOpeH8j+BBW1YT1tV5NOeBqhQvR8K0vhJzbt1tP+GmPNSJTlRrSwaeJFT
+62Vc0tGY9TKWXXbtkj6t5pFRWMfEHEOYI4DuDlZr3zD5YJzh1raYIDABL21aZ3O
Etdpox7toaLUOhqWGYEG5aWfEr8SfPGJCQY0WaOydbVVLqiFaJ+sE0oc/bir4v/X
MTnUD8ncPpfoXk1MMGYyPkiHr2RwdX/Hqyrai4QPZrSiael/opjclDkNkH6CZEOX
ZgN8L2yGG6ZgzGbg5tz1oOio8BmEUBI9+cj8/qEsPek+62myCq7KciTO3UcqFsei
ClfScqEWlTuAomBtpSP3EU56phWPbB/Q77lWHlPqPsk6vm5B0chjaCaHXsaUdgmA
QzKlstD5DOfnC5EfvtTQVOtpcrDtGumxpJaxkabdDgiGfpiOr1k0WJA+61SHKznn
j4x4NxVfVHIGYlc45W4RWGebTdb5Il6yEGpSK8MHwI+7cPRPTjC1AgjEOzdcG1/8
ce4V5GabMEJ1msiE3wsVjqjeloIzyvqtzkExv3vfntQlV8ZJXSMXLwj/gcbhdT3j
6NHPF81d1ZhgcnhsHMpfcMjeou03VC/YysF5YmWU2ghSUs+jD9fj2tZpcJNcjuWr
hnzjOENnv0Ec7BmbLoyYP3CQ+ZqrZEuMIVrheFCHjaoDE/SZ3a17kM9J7WGnbKPT
hfmMDZzxbQmPcKMJi8jkhkoZQQXk2aXr04arrm1mMnFZ+qOCys7R/ADUO9AF9Po+
asyttZCE9odcC68UEeqItaVR2Fcudh5DWq4kdczNQbkvgrs5w3QgblVZXYgt5Xbg
RpPjpfyXDFIcy0jZGMmVxCeCUExfqVsHqRupNL6tkGeKn7wZsJLF6OBXMbCQeELL
zadIcqWRN09U02NcnR6WIKTFz83mC6AaPyLmm3OIaAZWAwGt8F+r5pSCZYXqzoBD
cw0/U9DqXakfWcdOkNLM8FLxZMrxyGdSx6lxUifMXHVwDiYxcoC/6oKoKbsIV9lO
sRvyoQ/ECtJv+DmN4KXbGqewscssR1XzMciFx/42UQWt4P5RCJrZ4HN7mowHOOvx
oQhpXOos32aqOBqWmSKyjgCOu0xSjewlVZ01P5xuVbqeOsxqoGq5RKbPTQQpIl5a
0UaUPIYpvSDFzrgY6J0BURCAJcjKCkEZE+6PS4ULGbytAHUK3JsYCvOBJrGq2XM2
ZasQ1J8BieikGZh0fjcxwVcMtZf66WXuAb484PPtVlQy/NlrLWAf5ZfhOelz6u5Q
W3wcOPdz7eXI+iYdpP52IiWNIxL4ZPDY/j5pOhoSCaOYGWne3/FXLiFXJn1yOFGh
UbEgXsBG9MXMeIfzzGZY9Wd2hPgwsCyGI6ne6ZbPw2cCSttbtMqlyFFZZ1QzkYBP
6ote+IM9JvS+QaCBgCoXzUM65QhngH9G8KjVBVjOTlpfYZl7Q5HDJ96JHBcXadVg
X/kmMW8vG0D2EcFa0rAKH3mIkbE9V52w+hCUCdubuydM7M/5TRQlvMl7K3NM//yd
lL0gJkpL9bpL3DJ82VqegPrHDnlSd5LcB82xJHE14k/h+M0g0fdtvNLcJFKDSZch
P3n2TV9nkAQVpgxkEAaShrLdEhIsLmNFrXkR2mqHYGB255UVaGKLxcM2Nzn/flMN
WLxivLGaoPuIfFddnFZPFqf++5gs3de1MCefhMEY5liCUD4fr7sy+BZgh0on5KXw
xvYbCQrZvRQBpz+B+vuLuzQ7pJEQXIHznS49VEqhv2FlRmAWRkqkw1xQaPoABtxt
HuoPSpeCuemWMYWZ76f/N3k2l6VFsP2HqHWm4OSArGg7G3QEEXpYNZS3o/8SxeHt
8+pgWcUHpRnSWe5YSH3IJMle3ZWKxmjVWFalPfTpk56+TxqEt37zpc1pFcDbUCIJ
xkC7dlMg0UjJ7Oo6wXo1L2KV9968UdIrUsRVVViSi2awDprJFoHwcaD+XwXHPa74
0kTexfSA2UtzungwmV9j0m+pmhceJzdsw4AAqlb9H//vqeDQwcVPO2mErL23kDX2
socqPjq83gfyNpZN37d/IkX/eZSmf1Y67K1My5/BA/UrSLxOruiW1GAj6+KBhQIL
glAkTHTtrU0HneT1prEemkvuVBSOQAObreV3sXmNAOEUeFE3TXPqSJmw56Lnx3Vx
pckLHFvnyaIaWtJnAJV8bXgIxlvAWB2YhXsBzs3rI9MhOPHRg9OPZckloJ8dow/3
L1AK5y2NRBJvf4DAQ/ZbS5rxDMgwM0VolstAV1l/beNRGz7s2v79D8nq6wvh2hKx
390dRr9v5057WZStSkXveD9I23louMhwAvXra1IVzELNHFNdoezeS5Lsvfzk3csJ
ofPTQp+Iwm2WOVAHpA4vQT0/MhTNr7PoPB5MQM/zb2C0JyXbWQUQswoNvwTRALku
MwXxcbcZR1wL9vWtesUZ7bsoISyZrASLx51wGkMOXj8/Mxe4F4tYGl/hIh0PAt/d
MnZWwEW2l9GrXmMaHbSXNk9RyRqPFBvWbIAjOYOThTw/ujpIzr7yu1e27s2o5PUW
GpFP5E3Z4awRZ1PpN0ocbBf3GgKq7x1EobZ/09Ud7u9MKzfkotJoxu84zM+DTTld
BR32UY/C+B9Q/BsMeW8cvgNC/Ek5FzkQtleGw2w9Vt7DwUGxE4ySsPVz8N5QFMeu
4YyRTWoF5uFqXU2JK1JvaPoTrnwhxil6gvc/PviyRSUCmneST11L3lZ6rODAS3Aj
IYcWK5TO88RrXZqwcALAXql6PcqNjsLoXvlS/QOe5FCsYzmMrtuSsViQdraHcLdo
2PTBkpnQ7PAM6T9cNoXMEtWlmupcPUn9poAn9q/hH/sUb6XQ19TMUrpksaiv3BJa
4ZHeUll+8j+CioR+h58uFw5Ax9ULU/NXtDAax5EVUdXIGNciq4WghnmjPrRTRILK
cd39cw2zs0W2A0SrzLKne4cEKphI4U3Z9RqkkoatA9mDq7K/Gyi+fvtnNxQilXWH
Ri5TvxtEa17+Kue0/0t9GRW263m9UaN9Kyfm4zrWgNzUNanZmQrRaiqH4FZQGQPz
S842/PBbNjEqq2G8VBKwaSxrL+JirNz6KkxgUEg6DMY3/AExu3NooapN8CNCXZql
V/k59gFTJ8Nh5qpBUzOjbpXBt6wO3VIhq0d0KTmVyTjx7eMY6xao1kbuhAxoMQv/
Q8Ccd9X6RmR6pWQJMSTIQzR3wbqWBI9Ktubxts8+BErzAvvApfJ8Rxi1LlJAG/Ag
WTTePs0YBT6b157dOeMxlRb+In28EBCpn+QGk+gJskvQ7/9gwd6aZ2NTZpRRHADK
nkB56zgSTZOfcrPSbfCd2D7kp26uUiYoYIzouI5eLmObtSryV3FUS6nW5EHmsyLJ
vulhDxRXLcrPTRTcRD2BqJGPvPFsF51aSwDvuBXveofuiMDW/P6gNP8UkQpNaJhm
0cFg4G2G24C2/Su2CTiZEmng0tZs8hPn1/hwXdPlfveZc8sRRoAgRCZVt2pkFJiz
IfM6qkkEwMHrX+PBVPoYKGCKMOLt859znkYV/3kTF6EGe4e7kC0NhIbY01TFCa0e
HQk2DeUhuPSml/u3bN6zXaxchFg2NmbZZyfrhpsXZMQEQCSCd53PAgNW8Vv5RSyZ
6FxmhFFEb7TlkDv3cjgvEYBjshaJF2OI4TN0A+PjFF9graRNLDN+Sg+FenYqigcl
Zx3YZGaldBCCLdXuu2nVsscJXudx9GasfFgauZQ0GcV1hdlUESA/eTxUXB3+o7sv
M3SgfmtmNfPGFVMpu48DTfDtYa6h28WXMpS/RKA620XQwZq4qzRgzAVzdkmi1+z5
v8/8SDa3ghrZPGIQobOJOP6ronekjuByinWPkfEXxvo4FVK2qVYx2IS1CsBfH/dX
dQHhCiqJv5psIkC3946VUaE6Fzz6s5IO9NpcGjsjkiNfyrVWzFOmK+EDIyLy3/lT
9XcQi58K3iNyyFqrNI93bvem2kCTlTzhOcJu+rK0NMQ6AVzXLn7VKcVpyqKidJZX
dzm313tpN4xDsdXKwJMv8L4oKs+yG6wD0//fiQn6XtYaxbRD6vfdKHW9iE+Zvoeu
rhX4HbkI1m85xNezo+S0QaAOpRL/fobSykt8ct+pOOMuQJcMC8Op6N0MoSMWYV7c
9Ep6il1SABTreHBduQSkfqYnl7iIt925dhWz3O1m5Eo1t9DgoGZMptbKjb+yaaus
lheBtCd8GD53sKZyF9++p4XUNTb0VtVdTSMIvYVoYENU8Vw3ffwqETtBkxP0EF0y
+JPZXi3mkSXxjQ5OcrPH8AkwQjVcPFMCJAPBlQxMoDmAjmt4OHHGq22FT/lDYsjk
NAK27qYsFa+zCjKxG6zFyc3AwMjWvRge4Bh9FXJmbvpFi8+sYT2uUCsfjKbf/AHy
tWO2XGuauwtI9LJIiWdXi0SJoJcnHQNvKqVQTyOGuw00aHwlXn+P+L5OlEKKA4vr
IEDYmaYLa5dQN9ewG+64BIfBZuXqOHkcVs6qay0Wk7C8ZIMhrxZpt16EfVH3Pie+
OjPcQAl/sJGNwjx33Qe6eIMbs8sABw6SVCs6HZcSScjqtN7I/Xs5MV6AvNVCxx0d
mEuUZ6zPQXmgocjeOVg2jMApd5R0danZLZBt7VHQLmyc0trw/6sl2wIGVCgbZL/N
vY4JvgXbm9OgVVGgB82ZLZyuNXk76BzYCwsg0KPwIBSLobX/gM8/NEK6C/XTtM7C
ZlRTxD9Y3ulnH8mFlZd7l7rortcy00PxkKnwpeYFuJpHejHFzHJLuqyNRHQuyEAL
8keX10/1wJB9kjMb4OzdAWCIalKrgEUuX3TcxAMTedRyPr8WZL9RHUIA2NxeJhAh
flekKJ5g5b53GXJgauewvrccIrQMbA519IwniskiYD5o77pzindBvrNLXte4vdRH
rLjCiqFUEGbvvrsNCAxuFLXiqjQ6gFXM6XWL3MlCdyB1iUVmoE2cej57rtldqhgz
2gMonaclcF2I7XHAAPtogAPdC9qaaKvGSLrUTPBTZ0eLxML+l03i4sEpcZB/qaNQ
Q3u7f3ZYOvk4QgQ+ROBFY0Hg21XXdCGqH07pnBJ+vYUabzgjspV6L32UOJcgjQ2Q
CwcIyfHfOuqnuCfnzMrtpdlx9xUclzsxch/wQQhj4Sm0dnMV8HCOP95dlP1eHbbf
ru8t85zJl/OWvGwu1lgn8TJnW+0I4zb/r2V4u118hTVRh8fOWUV52LZ3g9miXCJc
sQcgVGJjrSEhTkYVaL4/D1MEI4zK3YVEOYtKp+EinvNbTJJBnOQnGZU+kyJNltqg
I1u8nzq79ipIecLbyzpmq9wqVxQw1ECitBHix4Fxzdl+xYJ0CKR0/GGjONQ43Pl5
eKAHHeM6WC2+qJDbcGlkFMjgiQpHXFFFnvF5zwNcdWiWuAYq0q7KlBcsBZUWumrv
77TxvfBT0IrjILuElcYL4jlYBJBoj1Hf4CSI3Xso4L4Uiup5TV/mdtM4nq/pcnkW
dah4IWMmG4lh9U+UQ4o7jA289UCbAsBMkY6JybPgLbF5FoQTLkT847uOiG4SwKvb
SkU6pIxJvzbnZNbPnsxQrUkA3eTij8FhqvKY7P+3SJduqweul8gCd/YB34+En0ew
emDtOsJhacPsC9agkm9Pi9tTF6U4q0NuiuMQxZk5QIHQef9BOsHn0vHqZLBb1ImT
TdnvZMhHFfjpAP11zhDjhD1X1lGHGbhNNnU9+XPg5+LnE8fmyCVXkxBCRP7itPJv
hSrIImJwhnwSgJaXbOKi906X1RVjUTeDBIRbXy5i6qFRNHjOmV0akONvw+iJnh5/
b4/MF7Bkl4HytZ7UcP9S6DGzngHIypqlTQTzLn4Vw4LaaBTEcqtyrc8YNcAzUYp9
o+kqueFKcTlMh3ZqhPHTB/TqEU5X2iklQq0jbsrKdgOd5J93KzcDRo9UNUKeCKS/
eKQxj7mMf6tWF+1NUbeQbhtMd2N883W31hsP8kttlDb1hOV25ijIbOHFWoEWb0ge
YkRpXXsuqcbTi+F85SMoiSFOs8eMjsUMd8TKDPyUOPSpgiH+gJZ6Yi1AjLUAMdhU
a9dcRThfR5LrGJA/YFfR8CHKD6mTcRPZ7ruRSOEnCj2prBj+UYgLsmqUDwakyqAd
+GXe22QXl7Mwlgz1CwKF+FcJ4Pb8FfVo+yHsCmR5XXH7Scwp3WhxxDvxrkIhydSv
EpdHMdwOIbAcUqZZ0WaU+H0RaDvS+YUmGu8z8rTGU1ehI4Vc3aS3AN1UA9trj8io
4rPBSMdtBsgmEPkoCHcGHMwaVggN1hqH+0ru6sTUAOk718o8ZkZFtP1khTyyLBw9
1K16EZiB8drYCwE2YpzDQsm6EjkQiyX+MLH5m7nfwg1wXqWBeWHrME31vpLR4JXg
B06BLoWXQC3beFGf3b7kuYdvY02HIWfmPjGspt8QWcfXfmI+V25XBID4qaAMPXoF
6GKZLZn3QUMaKjhuPrGhJwg/fWng9qL7GstED6kgxzrD4dtR0e9rv6/vDdFw9Hfm
+xwoZ36X8tAN96hgUUdxT7hJqoj9xjPtLXXWKuHKbAQqVOzGHXsGCPUriuYh6Mke
EdIFPjngCGaCRFF4NHDXf/iG01NsniJsrwrq0tdcQ249/6mjLSSy/Fo4QBnVc0sE
zDYmaY8Xn8x/MMGErbD2skF8gRu0WpQQm18CdsfL1frYJQ0UitN+sb8GriqdXVRo
nq44P5ZPp4tc+Z8FL435zLzHl0kGIBBtM8p5WrqYg0xMj/BQWGd+M97h4T3zb9wT
5s+rPSPuHEAhf86R4iUnOVhaFA/QKF3teIj29fuUYnG0ET98mySVwtXvMBkmuiIt
5G6vxrfVy1Ht7Mgcucmp6Nu2Vm7LfQ+4r6pdIToS1RCgfowSAt+6mp7G62oZlbMR
8M1fayAOaT+TpvdTYivpjqVGnOkSES+jyxwswWmpoCbQ2N052QjF5G0UkY2e9wqc
6nwwQayHF6foCqhtdKmEqvPbRuNZSd9cS1K38wmZzd+R83GDo0EPH9E7VgcOVLfq
XkqiTHJfA4uJ/mPvp3clPZsgTGl2DpB5HY6c1KESruSyzsfBARS4UuUThkCWcZTV
N8t6pPRje+k0xcXV7up4tvWHFvCUfnxolb8E4ubIkP2slZNci7YQlp0E8R/HLpV/
7XAQ/IBkMMjUhiFw16Zr1YvnVHlwAUm5Rugk7hUBE2aMtWQ+I0EUJUWRPlQzrlG5
ZikrXf+4iACu+W8RWqsbpbQqKXsWeOGGLuQ7ieBrS2JUO+ZNLalfj3zEZPD7rTpH
Sy2ZZy3c2Y3GTSEN1uveZmZFexRNcIN4EKEM9hAvOUsdJzIAu5f4gegdhMTfmlQi
6VnZ4QvFVhMNQnfvCu6C+/lwAsPorjUstaGEZoxIVANBS7qL4f9HJSQp8ajreD3c
NS71orVAydAKLpzhPnxOoYcns4CErAymnCn+Rf13Xp+FDBlWZPxRam2c88Xo/uPw
HnvaamCLL9TiIwRQr9MAXDFpFovoHR24XR6+bBL5slw6ahNXawG5fDnYDltwMua4
lqS9MKGcb6azxFlSupT/BfjMgKezoo7Eic9dvUeL5AMgigdO4NlQM/C38HMYtoGP
HBr0IQugf0/cOofbc7Bqg9ixIsMAZvEfkFexYCVjUekc6e7YsiOlHONUsiyzAcdG
Y1qDPtK1lTItbcHHZOrLu7C9m9qOAMAVuj2LMl8FAXBHr2Dxd+meM//lh4yJJy+0
gQXELh3GcctAoF3tVIH0MxrlWfT97qL3i6o0aXyw/0Azhdc37pJiMFoU2Wkx8Mqx
a4e51gwA1vVmUT8jiwAKQZnmbxqUtFibHxWAajHw3ym2Le0+pJopKLtxL1snvJwm
OAbDWD7sx/xDfCIIg2K0yn7jRzMfvqDlJhDeT+DWk2rwRcfnCxuG33PlwRuaSHni
3Y2rNFjcbxU7MWp+46v/3o06b1qqfgiWTLCMTwuWcrijvz55mYpuFSxuFJm99GDB
TQovrtBOxiEPwsEFvfWLgvXx9VseujC27DGgXVYcJECRYz544ofFLQDdEc1NaP6E
sjF9TxX2rcaSYf2+wdsf1KVLSPbLCBsxndnFaZSY9Eq2vRmetXH8gtQYoifSmLS3
6KVCzWUomV2lKoVvrDR+YWz/4eDdztjbjg7NMhhVX/xWYjShmThb91bvT1Fw4V4M
hF7cl2iayevl0sx8Fi3eSlSsaDGUDp5Ukd1/JA2ON1g4KQHq+2BCnj3EUPCjCmxp
GXmkzzYo1RABG5GD8bNkhPveheILu9muHqRI3rjZ2RZ10gaPhbgkmUnMDGCuoa42
BswNbJ7ZVSsF03j+HMLEJO4M5RkiUaHV6Gj2iQl9lpuqW+QDoqgzxDh3N12Ti9p+
qjoAownsrorSlIux+fdYUtaCVNCCecZLkOkCmaqm9NMSnPByClC9JpjAx4EHJRFI
wgBYtfwElpGDdB92j/0yHwsRDrFi+HXCwQVjvj0MljXUSCsez+ugr2kQM4h4AbKs
89z2orqglhzzqEkTMsaDvEhandBHrZgxF8jJNvlctgKoA3QxNCLQALS2lbWd06Io
w1VZb7FhmjpdpWBq9DDN0DduEt7QjboVZqXFIYFZgcdmFcVIryAWtBzPjR9QTjKN
ohCjbFtJrZj3M9GDAAVim4GTw5jx6QtSebgKBFDgXBysDyst1/5yfL/vp0ka39hT
lE+3kQ9eLZRQ580eyBT8iTOVWYtRcu7Z2tVJDVqQ8c9o8lPu0bwpkeEyTJNdhAqk
Gpxrtjst7O52tyF4nG5NqzfRMxwhtRaZrQJMy6Y15F3nqbcO7+zKraXtFLvw8dMF
W46+cSe7eDbeIxlUiPLnEZbUMOyswznhf5BcDxsxtA4/NGXpgH16Vw7xDSRsSjIs
CdJFSFKqwYTDZT6A+Uuj3TW6qGaFgLE8rtDDfcUWVRGlRP59DcykpLUx3jJ/Rbtr
SAxeIe2j1WkYKUQIMhISX7F77upjYpnN4CB1Ii79RNnuuM/tmF3hKpdwIL+pOF1v
R4H5ErZdQKxxWHVmCtpIAEfQ0U2JgWKAbo22W+OExrLGrg+FHprg1GZyPf0ZTcfx
KS2FZ7mPZqBCwnR+MJaAQWfBCbtrBTTNgpgfyk6Km9M3sMPTe2fKi34cxs7GYp9l
XOjkFzK5ED0hhUdnYX0edSLAE+4GnfMjiXqe6YD4de4X7RJK67MLU4QAs3c86vrL
OdUsigeTPZUbjRgD5RB1pQ37VQm7sZzk+wbckrHnXlos7yZM40Pc5ZR4z0hhwdVz
itQa8uWMWsLk/LezlXZ1ZRMoZi27BFgHfqbXjFjbYGbSBFj49+7YM+ldwHf8GmQ5
rZaNPP4HJ+Hmi9MSSOnNlXfv9lx6LtARgogrm72UzYM6YDYXS5vjbGZzkpU0knUk
OV53PzmuYsLfWPf6rgFzLF5fzx33uMYQcxniWLqIrMo9Q03PBSnso4zNI7qQAjLi
vWI0lNsEq4TSMGdqpXZNg4Ft3CAdcNq9eZp+AB8XGNe2f8ymRaaIzKhLMJXNc948
PCYxrvbSf2IHnNKgRxc5zQ2n6sMr5KoEir9RC+TDcdvx5K7tBAmce5YF0ZdX0UVU
5wsp1YvEVYCG/hnNvAYDnzpK6SBog/z7T/SrFaCwLnbeGHtqpRTOG1uCMRMqH+uY
J+lQAScK0BYISZ9WJ3tl0xMR8dIbqnfCLZxTdp49aLm0/C0eqpNZuLSajXvJ+x5R
1wgu7OBzqntgKEWvlD3g7Heo2obNdjpEbcMgMd3mRtEDo8e5aA4gdH8Z6n+2U50e
j98J1/YvJcmPh/7FV7pb4JDA6TpceeMJPOtUEkV7yQ2rJzzcumv9cLwPuem3LFDB
cw58Kf7WbM/hNz/1rs7aXNca1MWdOiH4cy8Ja6xfXJj9dTaVRY7b3hkHvpvM4aLf
IAWDAoMtlsyReuQrwimR7Vcrorv0MjLlH2HiwECjj7M1a8KiEPXRjsPLYSZDlq4a
aos/wQs9RNCTLh1IcgY6uevbpK8jhZaowg7JUzD0W4kD35WGl8gZt9/ukHZUZxiT
UXFvLUfucK8GI4BdhNdmefIk1gLn4akPp5947aNYUszybtnzfwylXO7OntSDHrkn
velDJ+o6wKF3Bd9x24csv17Bf9bxn29Y3LfWhH4GRFIlO3YmzG1zhVXzCGe+XvEi
R1O6tLhj0qAj0iWRkJbwEKc0wXM+cGg1+pkGs6O9KEYJTL7TsugrxJvw2Y4w0KkT
z8TYmN9YJPZtkXG+M8B+W22MsVgOBIlof1KZ7uSn+6OHmmHvxgPRdiUQNwi1mx2J
DSfqs1ulHKpN1Uajuq9isYGwiihzCx9PjYiQ7c/E+IWjRGI2xuDJN4xnrwD9TfKG
PW5vDUlg896psaA30pjA1BscYGZSMjp10jWyUBpSXuhDJlu1YXC2jpUjY9aL7uHy
O0291G9rcNfRkAqK5lpUcXVzvBNQOUS4QvQHBOJKMh2lPSKpJeYhjZMKV4B6rcka
SWCIkCeqknvxpgrJkbjFZfquruKY2XVZLynlh5cEn+ZtbMyNyeYCLcCBQi1Q6a4N
I7BT00RI/sRPoAOgejisfNQeJvbOqGz49AuWU/z7u24pZsObhZAvEDKzorvJ2zVh
y6EtpjIMfGfPCRoKn8J7/0UHHyiMOvYxO4PRqxkoolT5qAvrCkBTD5Kg8I1mmajH
9tT0cgm/FZI4m9ZkIR2cVnBFi4/F0K+ZWONsdDY9QKi1AReXqYqqzb1Zl83RmmaC
Ut7lzXDg8llJ1e5C7z+Zmc06Wp8HUMR6TnZVx7bJrnwF1Lg/pXK2yCNjQ2BXjuTb
ZCSs79ljfojPY56WKwtI44OkR2P6IdpMGchmh1F7NYp9EHvL1t1JkCSiTU+Lyee3
pEjodTmN/iEyljTb/3KZoixdEidpo2CCoTz97DXCRQG0fJ4WT3+kmyHLTplidY2w
BGDTTljJy75ZnnJH95JOXA9UcJ38bWYbgmL82MuTXddXUiS0cqjwlHGUnfKrFgOv
BUwZ/Dv2z+SFapJgBzpjHn33IPcWwsuE+4F30awykJo/EP8JjCYqMVdCRWyErkX9
P/EzV6h1cyyNVfiYP5MjWSE6IWLxFUfWkfhcJQr8HIJyPCtaodr1CxgxZO16YFP5
6KBwgRK4H+f4hkUOQzSYvDX5It5G32+ZTI+A4a8OL+jcVKz9EOqVIQac/5pmsLe2
LEKVeSmgN3bIO+fICeG+T7GG39TZaFm8izCA0avpnsfsOK/mNfIMqQCsjPax3vdf
NyC8NV7T6AOihESNsptiHSfrxAS/lyk7uvxThTRA7RfkqrySv5znMQCcFyne7Nr7
BNrbXfraXKwUWApmJ5JJUdaE+l8UfZNB1QtiEXy/LmKAgdx+ptfcGDNMIvb4popU
W9i0WiC3NdT+3PBskJPjCHnJ0NayD2ITgMczK/k7lALgAYI+OY53Z7YZvB4XdLfK
Fm5mclxpTBz4fyW1EfAvxvnmqt2zfDO3l924PxhDAiIIVb1tDCwdv7p+PqTTBkO0
h5fOodMnV4u5xZGIxxc4kPrZGzpYSPt8IygaOiDaLjXQLAumQF42Fv5bgjZFk8YL
DRHeH5VYKlh174mt2xdzPRAV/Ntrqvdss1QY1Tiv+XTocBjWVUS18PkrfXnmbPND
T2+sblwCk1Lg2bUQA7+j9Xc3PaSq328R+UlOYu5y4vybFKXuLOz7pLhlilF3KzF9
zC6CLkQlU9JI7IuBXuHflEJHCZT/tLvb7/TonzI/gAXUQbEjb57nnSatiC6UV+jN
Z+9M9gU+f6rDroVZZR70IrO4CQuYfN/DKf5i04EmBIoKqtmDprGqpCeCWSgCZ5w3
S5SitPLGMtIAMimHufHUACq+8GAo82sCIYrOikcSLRDguGGIa85jH3gIp6GIevQo
/nAggP4MKtuOfjGcXpDIO+pSFCltpqKun5nFDoPQZp1y8WAPQ0xnOkryN26BkcZU
isfq1UQ62p/v1RX3BcGlkIylub1090DJrLrKbSzAkx/mV99wKe6MG5TOeV8aLUiV
WLKRsl22GuRU3s1dgDuTBX6WR1oSY4WUS4nIUHymaS+0xel8DqaTtcCKbTV/sWOB
5fT3AmazjKKFWlA3YCswl15INtveBtPHqnt7UzvDqIKC5FvrJLrr2PmUHD5MuhiI
h6perg37/hs1Cu/+czbs4cZeYu9MgPwVkllGeaVrMQsoB1DfxeNrooBlxLNBJCMY
3JyCcQwYW9c9144OwsYY72zO06a0Foj8rGZ3Wrm7oWTy5N30BUyxgjob5MARmeWC
uQMxH7GlbQ+wUIOOQjg1JWjbYJd/+Hja+bHnYfljepi8vLpuiCoTt8vD3kOyqIka
i7F78D3Q8KPl4JopK2a6WwQAmmmruvCw1wKbIom6E2sj+RWz29QTGh4oAFevOnv1
D5JghMdoF0kvDY8aN4AR8Q655DC9gP2WRau4q+qzXJSnV2N2GvVGrX0hl9dpLJX+
LZAmzVnxhFnvLaVAT/ZGWuZa3LPKBGijL1wj+28X2rWad4H+4MkSNw1rhFGOwl3b
4Kql/IgHFdxqCm5+5xJtkj9ajvVaJDPQoapLyon1G7HXh/MF6pNubul2lXKqZQKp
T4Aj8VjNAJsO/OtZHo90HXgQ38Na1fKN83QKgClbhN+SOVKyEfCbV6yXh608a02a
uu8e/nlauLsJKuxbKk3oK2CWDujQf3eyKVkkN3tV/8WfzXHJi2LzYvdTJeGEef6g
hfqcpt8o6NdesSveB4U3JdtA0JRLVm4lhUZcfXv/17qzPXn/WZz9KDW/uOKrU7J7
GSNiCx0rMlz+MntweMV54c9Qe6d7zhXO18+8865RAWJuKGnzpb3tibQq6e6I+cuP
q0AeqCqnoSaZeoY6+js/bLpPSxAqjlMhA97s6HYg3KsDOHlQ2wLgUWritXou1TIs
ha4mv+NRN7StKBke4A/twHD2rMoECnYwL1ErdK8oRsjKufcY4MBAAHMsoVSIUl6U
nM8+n/QAOHfizNAqc+/JbaeTiqxTsK+6kKxXNY00TiPyskFFrUPNGKR5lBQtNsF0
mwNSjZ8pSuvHTJ795OgHpXpD7lLHvp/5WgfJPd+/BpIpnhIeplNRNt/W5QzIYDgp
n5XcKovgWzu52oAHFoM6eIQrGASX5GDZIOK+KC6l7i6CkoYHX6F+BK7vBUyV+me+
SWbF0WJ7qURL+cU8xfksg4izmmocn1oVeGSwKhBsXfTA5xwUNSEMVErUewg8Dq5K
YtPe2/sZFQPMS/JQMk1f+nFpIfUtCgnSr0kk59929J5IB2WinbrJv7SRU+yBsx+r
ffUrjgGBxhOjo9Ty4gVU6tkku55/oznxx8wbXC9nfAPe4hOCzvrzf8Tk609754Oq
muVj21nfMXAql+0e3LujSEPkOE7vIpJp1qbc9HazF/fENwiz1NUup3PjY7Jhz5Vu
Mkezd6Cro3vUc+6CAP1DzmByrnVl1KY6qdvGmrOfmPXNc+OcvOtS5qjkcpHBx51+
e0S5z4nAenGRyTUM2ZmKWKjAomkNKdWI4GWjsBYhGp9K5ZkzGZY8aggeYLzysJnj
nJZEQZKyjmw9yYwrPgVRSBc+RQieciWMxfZf5DWYByFd06CVCDkNfIdO88Qvlk78
TEn9pyMVg4ZTCVZgjrtjamC/ZZEw4zUPUCYzKmAjxyn3DPdEr22gvE9hWcdPSt7n
tIkN02EVoeDjwq2ToquOALTumeyFajOI2FnbwkbLridmjFomnyc4hBMlEh16SdqA
4fUd6QpK2dHwbxT/5MB25g+OeiAOr4Sup7wIxeNEkUOQt+rWlIBXkKZbhiCIm2z3
hMhCrmqRhOnxgM69XtNoD6wfa/zxaLkh+MYkLePCrcBxfhQPjcq85V2fWCKHFrH0
O/tuLbco2LARdh+jACHXFvBtHSZSZj0GNgNycnVU/tVHrQkMMqiESLeI/u27OmEC
e0EEh5RB0705LN2DTJYmicF7xZsnkdLNS7XBVkv7Fd419TOb6Ze8eJZpydR+zIem
iXCMApeDw4ys43U0GztiFKW12Ciq33ZtBpV4q5raTG+J1lwL8/ctCVDl5x4m//bC
V++1vGhckGLI6/4G8IRVq/qDZkz4/ckdyccIA1MqzJK4WuP3btZAavDiIoMYFfyH
lEnCRXSJkksvM/OMZV7CVMdL/6nn7o/eLXX29d299JqzC18YSbbEexu+Hp6NJSIU
UYuf+dUJ7RmblsgHUY1EqP4zwJL2pW51zw/Qjob0XKStmPWv9h370YJcNiOHFHU2
rR1Ui0AfOV0tkb933QseU3BUv/R5RqkD1Zh/EXvqNE8x0YMzWS7DibsHQN1mtSye
apX0cuD2SEG8qYhemI4+Pyaji44TeAXRQmWyQj7Go9XmoChIX5WHiXG3B+Qgt2wO
iZN9f4N7Mxx1BSsM3U5jzAOX/FaLxdxsiNpsUsoXJcifSueu6aqRYAgLJbZZj8OQ
9EUz0GnvpUJS8vlaZtez4kw0GBXKdl9SY9KlQEf4EraY247rdqlsckhLejPsu5ay
YOHq1t64FfFdrFDfwGZbO/VK7lovebSLdBWfZtx0HE9SH3j7VA7XAiJocudokMiJ
PPW2PsqFgFasSdkU3XMjZMhGWJ3evbrKGN0u4GiO7uxOanz1Mk1m/KXfWmkZAtRD
70peQUpGX5bVZFmn8lCCP076QXtZs7jT27rH5jjQ/HfIBIciEajaY2PSts2W+3MG
sJQOE4+PBGca/ZDPbkfGlEiH+u/GiFhGU3DldK+jHIrboexqswxVJRMvFUokLqrw
oUtb8Uqait7k3Dkb9jfakP6gvvgwyq6XPnYb0UU3mCcIny5wAskHAesqgDLjyler
rV+epMxRO3GdaaE2ZVbgk9vJgMaTVsAVeRQ1HQXQMi1okq/5VSS7Q1qvppS8+eJL
rGoddRT6jT9r2gEfxoyWtJ3qVByk7P1J1pX0vz8TGQ8tkL+2AoXAaNX6TMce+3YP
2AlXqP6QHsnYxYceVlWplFAJVD6AAjb+V7k0O/HhQNjywgjWMuADdv+F2etnzjw7
yP3t6R9loC8qi0+CHdvmy5nnkqnT0RVB7KuwDJgcQ5SaI0S5zDAWleoX8G7HlxFX
rer4RdnBfZozrLPnhw/DuAriPB/rtNtIpemmtJKglzBLV0fUH94uEZQ94jTDJOZX
q1dhIiPfj/qzNtUfOYHOYP+ylu3dlZulftm1qAQX3qC/Mrh8I//NXv1r4mvdF87J
ql/5CoUPflIP1tHI9R/hLk/o0rr0EOfp5OayW4eCV9/km4/Hie4NE0ZYKqkGdyr9
cSPCJrVIEyLEe0htFMibNIJOzIkLaH92PlOq0f3+f1RvrxWYGsaKdABiKZsYGKTf
uaH0PaIrYHe7dSQ5VC801qXscfmMym6OyikQ4toFRFPEsIaPkx1S8cfda2mutegm
De4NlhG3qylwUtXHJEdSlvMHxhTsux2CkD5wydhbJUJ1YTtbSncItLiAktu/bPN5
t5KhWmBtFhJjVyIcIxkRJ8snuu0xYQ/UbttOL/UhyXK5kC4i5zWV/bVYpasgAx6N
T+WNxWqV3M+vET+8s2glSAgTIykeRUiltNXf4NmOfoSQHZ17ArjliSbYHIVwmcXI
uDKBrA18R+ahq3UYEIULTbKK9OzNev+wffeXcfq+Hq6S1OB0wsmu2gCbbskjtOCR
i4qkGD48WVoUoPk1E0h40yGzrnognvtFV/bF2e3XSsD4EtNYQ4VVOj0lJY766fqA
GYd42hODqU3B8YqxjeIYb6UMGAdo54BGBLUBpWiwn8AcJrslgY40yhXxCItr2D7m
Z+SAlMH64dGRE8x4fps4kw5r0THJR0eIz0fU/YhGcHqHhw0ciGJYMDQWWVORaH8Z
DCLyQ4PMNDysDMUZUGB5YRv6Wz3bJcW1A74Y9RNsneQITad/OuuD2o494Am55WOW
TQhfxhxS77m6VpvOtMGHG6mLBZmSbhLCd6nHDek8V3Q57gy/06C/E1o2I5F74Tm5
LRYbpWgBCE9ZJwCbj7XHqOsA4yY245CS8Qqamfqf5KsqM9RGlKtVbzNUjrUiUsft
b1S5gIVZCinhHeSH2F+AjON8XQCBdayCIDhjmTfckCLrs3n4XSqqt9MClkpNFK86
WEN3wiZcyu8EbSntjwO81oH3tt5ov51eGjoDxYHcHDNmAokCt1+LssSEiXlMPj8a
hm48nJ7qa+TbuBy/LP1HBcHKuL/PpLhQF+ycyBC/Sd5B8q6lugsYKF/4yZuahPAo
WV2X+MJY6B5sbkid25i8mJf46CXYULHcGUQEvFnHXiKmJ1iRnB0Y+eOovjSPByBY
wmINuEKR+SO/c0yguhPNoejINDkbBjQJPws4/dmca6E34IZBuGAReysmVZF9qvuY
gE6LQPTa2uJ2armhAXjmKb0N2QEEtuoN/IjlA6fpxXlSNVjxo0I5oZLf6u4kkbNv
lLnnqIUGLgfFjhiR/G2h6gkI2WN5+xpmz2JkW8Np105R1jE8r/d5JEqputFBG57f
Es53f4utSrwYClLE2OIjuanOdxzmF/Sfwpu3n4aTuKsKG5i8vuaE/A3Icsuw4SnP
K3EnF6lzTy1nMdT9Ij/DlsTGbjqJXNJDHiWv4ycjsjZDl8PhncT4ybfsgrXfNlBY
+YQHytWy9F7HGqjFit8DM9yAgEADsUqi10/s46cna8/Tu7edVy7dsAlyKO2uBsLV
96HB+kQ8g8XZRMeShrlTB8MV3q7LFAD/wYfoCPpmny55UVxZFVM42dYfAeMJlQlh
xoQxsV+IUQrVKB5Fn/ShYsIvUXxX79kasxy71buJgrA7Qr7RozOeXLk2SBsJqgcU
pmocZSi43aCK3PNwp74+m9jx3No0cgYsWmx23jnplSGPul3Y3qhkO9AgljOEWZBO
ARl6L2oIqSpQqRD4tyvdTcXbiV7kgUVS000MboMy0/iDqHr87PCmIrqsm5Bk+qx2
1HK0yk7BMd4UVq6SP3ZqR4/BwvpmnUGNL461LHg6r87JIhnZB+62KcsyM8/Dc33r
W0om7mA0oWyUt/uNX/OO6iejBziNZ1uc6kUAaerhCRkg9i61zU17SUbET0A9kPk2
GqHX2ij7DcuVrYTjy6xD40sROq/2/qGMLNg7UL/MluN3Yy5C27IiQXtl80jo7eN6
P09jt81SubT8poh8E7BGExu93fJa76KsAB/cw4MaMO40laLtpdsTrX+dF6xbv9vX
wnwqyt3lE5bGKsoUcuedB7zrh9TtF3jFfnOp5wDSL3d3jckWWIH8w3g1xiOOV7g6
k94Bg6FI7DJgyBjF7oSyqOu4beWSlro2HFasS57q/YBlObB2ETgI3RkQX7sJG6Hn
do7+MliLYy7tcIQ50NWOK6Rr2ZI4tolPNm6HjnNsMh7ky7CZ81qOx/pqFGwz8NRB
b7H8lgrH+XvkvzLCHPv7eGXSs06AX+wgUF9HprXdsFd4fKj20IgsPJU4dWNrEmGJ
1xZAevf8rDvCv2q6yX//enmXT7RPZhLfNVSXWRfpgypEnD+IA0flRi41Dq6DOoTD
SbDs7s7Qg/OalcT+WbpjSCljnSU9/EDjqxHhfaMFtgnhh2fM/UmyGdG1MCf4aASE
N2lF75vRrCLjQPv902f0QlPcm0HescGHGS28ztLT2c6R1D9XI8cTKWP9MW5mu3U+
CHccpVpzjsMhCmz3lBc1cYfiquoE1uTGAOVJkcl/rtgDEkM5euYWod+gTwOjDlOk
umI3nrzrrZnXUpLCSflGiwHRXaPicFky+6rHjjHBBDjKDZORdQ4dYiF9lVSQNVMs
f3v8IWvfEQ+dkQQv/jOnV3eM8BeelvmQKPz/IzI+rtIQeYpx9tr1uGpZzIxvb9ND
WAM352mpDSgMTkDF9Z8oqSDQxmhnagXOf6M9kOj1ehIc07EnU43s20o6APdnIBqE
OBwo45DCccGf5RJnIEyDaF0BLp0TiMiX2i4Xh/+yseDHsE4PRlv+1Mr5637hJEuH
rXrpeHEJx0ByDoB4C9uhae7lO+9pDLGt3Lm+YP1vyXxYVQwvHm8hHoz+/Pa9e0bK
ejuo1RtAefzun1XGnFlmCAY2gVx6Ggyj43CXB+nMSuVw4Z31tvnz3kDfPgFt4QO6
GBj2WjyD1A9YTYzYhJ0d7uk2h8gxIj8exUgpVqwuFvH9JfYV5q9BAQgYVWrNm1wu
Q9KIARuEbbjAn+WOBjsePGczaDJD10wi7/mYcM8c6l6+v72ATm2pkgk2mi7cuz6j
/5G08R7IPiGM/kArms8YDReb3cKIWJNyY6pk1F/y31AeispkhIAEfzIMo0Wmbl7U
UzObMwUJf22J+13azV3x9xSHesp+Ok24/dv3QJbhLM3tVRUM5kBLq+7sM0PJvYSD
/El6MGWtcDFs7KL/OqFrkLG1JaxAl3Lfgz7LhDx280oMbBVmO5QBvbL0MfIIWYG7
irifcNpCrpfrUe7rckd8FgwA0/2Hn9bCFBUHqZ3GDJ6hf7l5HFsSrrTr2IgsWEYj
CBUEM3fxIQl1S+OU3Nbr903zEDo4TtY0EngEVbJQsJqoAoI49P1quV0Mun5oyFG6
qdoXtyBmy8da96cPIFkpeE94aSuzX/LTWSn2Mk+QMW8Ea1Qhm3lN618/XXhKJEGy
3zGgftqr5Zbeb1gkH74wCj72MG3AreJnQNFg5vWKmx32WGvrqsU1LFPLNhk7NrLP
1U7YNXwSwHQa4gZEUjENycf7Ykro62KCj/eNEiHUNQPAc9BxoQgCzlKwPRRmWdeW
h7xNy+8NWPjt0lGtTBy1Xd4rivTAyY8TDezDpy/D4QinGuRQqFuwTZln07xDHe3E
aIiSTKXqNNuk1wh/OkoDuUV5HXSixksttd6z3nUinaZZg0Ap2QITSplXndfafpfU
d1LxZ4Bw+3HivDGJsmcNTVK9/scw4avTulwY2a8mfdC4RLnQbDNxYZWHsFm4Q/Bq
nMDKltXJiAyh4hoCTMJOCj0kCzxH3Ms8xq486TqTbH/tym+y/CvkBLEAJIfvYTAP
4K4aNNyxVo8aUMKx2XK5hVCNA/5a4HU3kHmmJhFwo7365LXw/7geolwvK6qSK68K
tYdLdlzrKM1YykRuHQi41pVDdkmxIxgYB1o4QR/i1zPS0qRILa/uK/6Xd2cl94ss
DiuT7cGDoIAqn7TpX/drLIy1XOJXMSaKNNH85L373auxFUef6W9FTGRI+Cum4TVz
V9yZD0CGGdSPU2WsLRD67ZTQhGrzvaHAmJP5L71m/yWaw/kvotTlNh/m4pzr6iBO
dWxoxZHxXwdFofIrBGB/3J7vQgUGQ+qKmBdnBccbP3QS5PNgXqTQoVdiHIVzFBwW
3wx7QhDBNKmwXavXzQx6OEP8czQkP+pyxjvqMTwexDsHTrOx75gXXnSZL9KbMWiS
xydMIYM70bsrSv+ObDOtZyCTbjE2M26ugeZvKI79bpg4ibC/6eT0iNTjWBiI9x8W
0x7WSraZW3FoWp3yZlaaYSdWZNpPcw9TonRL1nQRpBHjUCqvP95PiEq1c/oFnvwh
0tNROVor9rpUuLKwXfJDcTOj601nqxVS1D+MVP5uE6hrV2CxvT7cfXDzu5HthWxR
SeU8yBVsFMV/dPX91sm/bbApC2YG3aC61whA5sYP0Mkv4YAIudV3Q1JWmh7cjf45
PDBFyP5xSwlAY6jXvTU41uhSwJNMDa1JOV+Aelbv/trS7CGphY3TZBIdf/+DWWzA
XFTTIsbJAKJJ5shbmaAd5FOODmRI/IEQSOLFvfRrgdHCrrLbinkoiAseXdkAduDl
sym1YZzz6o5Q5awFn7c70cjpTxXrxediLfexO9XAI6Zcp8zeGRWIb8cZdI2whRgG
YXrY9OPrrAS97PdQVxHywJ3L7VCdJOFuozWAb7R5C+26I7E5m+amQd6W7MHpPJh9
E21A2nrMtvlisqyxMw1/Rz/9mMDU+706rlh1ADRwL3yS8VFijh3hwCuIjbnfHLNn
gOrdRfWEmOvdMKMnQLTAGYBuZJVoX0UKV1H9PTAf4Vy7Fjufb+rUPIg2LMxjhf72
WED8mRBlIxrabVvqb9Q4J7N+YTPKDVzgUskNcckybKxiGbFnqxxqyEZddgKKVC4I
irAmkn9TxMqayy5zmMUtn7I2/1cFKNmI+UIHYw3QCv3pKRAlX8GPvKNOkNMXpAhB
NbaKlAVMQZlY64Rh1VK1AuKLK49mivoAHZkPFwBPIrKRib45TKHigh4WMMW9T+PE
lU6qBd8spZHa3PgyxSh1zAcZpBXvZ3lh7vlp3h7txWHr9rNLJ0DL22iyG9cE2/+6
/yRNwAF7Sulq9P4RuRdT9290D6qwqC8LYp+KmrqUfET1u04hGqf7P4erJZGIggnS
LLIwQnS2DfvyOws2ZgUz2idACLDACknY+etJGFsNOihH26zCjdQBgu1SsFJkXE00
ymEvjHVfv7kkC6Dm7x+cY6vVlWPOCIFUc7UZ0uayHKMSv8Y2dRrwVpf10WfaSUb9
fZBhOOCUnx48m7RizxfFHuEYTbYG92OlRibITO1HBe2/dx/ZCezboJK+4Dpw1PQK
i1J9Jm86WsHCv7exxU0UcjpOESDCb+TDr3UBVS3DhlqNQ6v9yQuF9H35GFDaMNB+
7gZ7GZTdQJ5cIMBsspKiwdlI3cQ9b1kx36uZ16KZ4xB2aPrNJwJdC/A29J9RfRSo
oUSgY86VxTYN39wHaDt3HclNbnh0GbTvdw3nuwRRBKGbviNnAVv7JGlT0GEuNbVD
Ked1kHs1nvH/DQ/SS8e4j34u/TJTKKGBXCgHNNXh+kqSZpkCVz3p+l6GdlII4CpM
cHgolu3aqY3WseRNQ8DFbCxznr9AsuunJhwzWKF2ZN0AeT3rsX+FM9PwQQBx+s1+
TPKqK9ZqFe0GbupuskZK/oOLU+JARfmZMA/+UuaRobIm0UpuHf2rDiT5JAqE6mIe
QIEPjw/wBVEwHkE7dRTYgT0RbCpNruV4jmSeM1o5lgUoN7kAolFDDT0ExMpz2vvz
N6ci4GpF3YrUsVHuiI1+4qVxO/9k2YA/tvajh0FbqJ0W4ka4XbnR7zPuJDamw79d
tV+GiJt+dHJaIixJ5ex+iJlacLmQJhNTqjeTv1/UE2eK+ql32Z6m3Ew8TFQiIp4s
zdOysGkuaV40j9gGRUXAslUPtCrTwUL05nh+q3yNJY5k/zN+ccSkftfYG+ky2Xz0
mZTfekythWm54QH+oDcE8IuAQZ1IqNHNiADG2EIjdK4+8g+pnPxAuAMfz1zQYwqV
vqf4bxQkh4EDRNu0BmtStkVURF9hcXbdEbI3PdUt18qAK05ngL7cHr96sj/SF3Sk
iYnFSvt1t4iGQEKGb6WfSUSgDtVyqm9Bkaj14crLGeDHKELws3lZoaTsd933x1N0
IBInEWSxzOqTDXqdXS8vwvmzCSIL8wryx/2QREoJxY21ePG5ll+wstqL3fPNsDqp
IAzwI8BQ/6eK6NjeWntR5CHhOIG+WFEGITo9DA9HNudcTSYtlWqqjoAJsQfu6c8x
q6nCD1M2JZ8fb9sQZsonJ/s/udRsn3sxw0KtOcYpgiXMAi0IKvIdgHKqw+mNgxb6
NfXlyQPx3wjYHOWDI//WDIN3Cmy7dpv1+gOJ1uiTw2yXtzhHibcUqQErtBPLnzHT
UtTbNqFp/jvz2QDODw0v4UX4yqY1LPChI9/SnqxsovfHtBUYo0O99KwBUG4SwI08
GAxfDVAXF4WtFyB2nujsFPAHMMIqKVVZiz1HAJelP0ev4YqM6o+vcn6BXsWAafdt
jdSl4oqRqx5T1Usru3NDj0xLsDmv0fsyWrPHG4rY4KWWvpBXxNr6tVtMsU6qZBL6
vY9XmRNr+QVttbtk2BeTtIb0z7Zx3AoC6HGP8lBeT+LoQSVJLQdSGod0HNr8pdMX
AtdntPcVeO+dAQcrS7iAPoOHx/E/1mDECh6k/SkvIThlPpUTQT602RVnRLnm/x25
xsITf4KtpSQL0XMq3f9SwH070Tzz4Hd4MzGO91609QWap34IRe9xv28Kl488B4zo
M4FVGx9ZRyWIgeTmVrWpU5cdhwNSCjtmRI6V//hs/5a7LzYDWgG0uVCRyPGL3Nm4
LTzdoYV/dSHd4guuse1+UskFP4TEeanty5FHQ+VG8LiSpAg60hj8nPSpUHUQ/k6O
JvmFqUgPF4hfikIQX8hoWlYEnsuypkjC/D1SxSiygmAJT4TQkrQ9GBRx1TFEnnRN
+w8Va4Q7fRsJTnuT4GkLTdMu9vq6rGa/UIefn8iUniXWdYzj/eIteKU6dUqFeR4J
MjLlGYm/H4pt+Y6h3IRMiGr3CrZo2Onbql2dVVPlCaqWY5KlbqqqpEtrNSHsBjII
ZJPG3wVbkl8hh9eU+Znc3lQg/WAtQ6LnxVpARkhRJNRpeIUyFdQpJr+3jowp53Ax
5NuMIc5EyqGVZMOvgvPMUtv33bLuh/JPFF4JPM0GpNfKuaovxsrVQQUwZ/jAI1+R
r/IJJLSJ6Hs4KXGer3cx/FkZhPisg6mt2J6A1E9enPD2Ewe5CCMSj+t99voYjmmE
6uYKwciC+Ma1YfaEh79UIgHsdlOLMSWUXlSdrr/4/IMEUED2ZrxLcyMhAD6yoFSh
vlHAOz6TQqbzOH11ImJ6S145ZzMf03UYw1VKqVKRbiF/dDincXKGS4kWBDIBET/2
nlZMD5YIGi5e6Ur6s4ry5+I4krhZ64GXXGQhnWwqIOFbkG+tUq8NhLgCGOmzq0hf
4PImxuhhEothCageKeerO1A4rpDtMD2cPj3RX2jNvbrHf4V9U5bE1sC8rOg+6uFS
PXDM/N+8/F/POb0nx+26M2ESDpobxV2GXUiiTrXRUevxM2j9k2zQeZPJbdH2I1bz
/b/nklfNtMVJqKh1RNTgJj5raSvvPV+NoNkupJv20IUx7hOh/P6uPC/++MhcydRv
8oYM6oJLKePoW4nWTMZbElcUzVNtlLme4mDPUC0uEr5q3Qox87xBGJ57CzF4pB/M
iue3qbmKgGyNl1SJzcq6pqc7GqOoN0YwQotZSiVSADk+glDYEohMlKp62iN9i4/O
cA0zitbpEMzkihGqrhUaO+CiJvjAfP80k/FVOdacSFMc24PMFzWWufwZhkudRn8K
A6uhZi4Pbb0iHfarI1l1gZ/rV/8bwfM8QoFU/oFq3yFnTn+KIYrhSE/n83MD2EbN
UuI+0OnJSWJntn9JkpcEapRtQuwB0Hjhx3zY8eUujXLcJNElxpA3qoA3Gpfmk/va
weJhJFC9l1rjvWJ/r8RJ2KMAw1P/oO6ElceBH5/3eE9q2zutWssat7xVziPKOoJH
LK+TjhwaGuOHui7JQ8zvq9MMtaxnnkx0h5yqfV7xdQBKOIcMEVj6Dxr/gCz5A+de
MHc6IIaAqzDk395sv4qfyt/MwjYBgano4kxk/zoOPAMBLaVFKbmQYGQRMU47NzTf
WJvWvlihC03IyALLltbrqbV42JAxRovonuT3+5QJlw42P/z3NQNrfD2e9XQIwpcf
sk2GH4fEDMHt1beJz8UVaX9zymycM3xAm8DsmfiOJ6Ln6mhOmURP8SGZleGb4sEo
XMYO43GtUzO8yUdDff8XfsGHybY7zZdaym/dLP2xd6REp50bXZrBIJ8+6d8io2y6
fAjuHDM/ttSOx4ZoSJvUfWNTuMMlxrZZ9ePYwvG/Hpqnl2POPq4Qz14/iUxbR1LB
3ITKsltK0H81kx56J2YLYTcuzzAWAv7S65Ho7db/sq6tbtfRvZ9Bsu2JUwIVt/e5
CNleLOI7L5jp2XJa6o/QMTVihkCsszq/6h67WeP4+kgWvsbhziGfCZ9oG/2Zwqqz
IpqG8TiDEZojrfZumIFWCPAP5zfFkPX6NVDVLAdJJyMT1ZHLyvErq4b2gL1OHhTl
wqTqo6Jfg5080nGfaIeQpF5lFS5AVL8vT2AyKv4+cUXsCbD6TnX8NyEh/P5efvqy
Rm++Mo7xzuTPl4eSP9FOR4LgDz92BlElgzePKwkKFHq1i+I/99PsWKjYBzgdJuht
yLyWn+PZxgSkLpyE/LodTBCsz9k8jt6rU/E30g6VyASp58NDqh1DVXi0BmFlu9Eh
cfg6AJOX3ICh4EpD0US9JZvkn1eY6gILJAaP1laGqQqe4H6aSaqi0gtN4WDXnHls
XYNK2hlAIvHl3LMaQDNj89NjJg/7FAm3vmeRu+vn3Sv2H4QhxcX8Re3yMHrPSBUE
2/ocTZhsOcGfxmwFViKxm+ZIjJ1iWy5vSz6XkPN0ZFQ2pfqs9H3TKLeY0MVB7wuU
qbnr9sJgtmjXNEvT6ADJiYWuB1bXncinxIyXu6810YDdTDmnpAIVr2toZtEHb3Zm
Vb2VPewrHjh7zx93+h98Ns3tC7yXhVLjwkJOr0PrkAnobvTLc5ShgfWt+WqHW0kK
U4Xkh3lcXl1xb0YQNREaCQ5VVK06Dz43MBHewcWHCgSae77U7DPKey4gRo8QftwC
Pmw57K0BUMGDdFUN/RXkh9O5+Nzjkx2bzHz7YChAk+rfD4Kq4c39iqGuW2KkFxdX
x0LGiFduKkfYHFvUZlMC/EM47OceGH7sF0f+r7m+HP42mBydVZnbm0HduSv87rNq
QLj5CzBmkIttPGVSehOJjcFcNPKXgMtMSkGZX6n1By34wDfAIVqj/xyU28vocvsd
ZxPngMPwNMtCWCMp+W2fhXGOaBvfVASUzCi/6KCXFEqcBsy+E5hqa1a9IhpAKCTY
KtuHIuMDSGHGk10h0+tnOOq3eqEpzwjZRWbnrnJZ8K6HW9P4DRdNL6XcjFvYvP6+
VfaQJpEf6GceRtGTSBG6ulXwcVYjX3htZvd/SK2fitYwvT1GbyBxCAy06BSd+aPr
4jmB8cHdy9YhESQGazGiFbV3aID+3OPm7RahjnCRuaTicODMJ7d0pNCdkOPeXqwf
eB3wOyfTYkwkrV60rUkUjaQtCI/hytZxwp1KlXgNZy2o3SL1gYI54I8rC1E1qC+4
xgidI5qvwWSxJNS1ZJ36lwpbnUZBlkmUyWhib/RyZcuqEOsTZFfTjSmppC/acRgO
PoG87FAeQl6xOe/RwWnTt580PtCpYZFkr+gToeZjssK98ulGNuY35foxzq+3oPlk
bryH8qqS4IYub+7jiVE1T1mEMruPzNm6QClDe9GxepRlqfVFrkejRbqOgYop3xra
j98tTahzAmke6E+bmSb34lpQX5o8xNNEmLnPj1+1s0JoP30Q9Kh/FcRk1gTNw68t
4vfPsXmUzABAS9VzRcpIgws9z+wCD8Ua7veqIGMnq2OwI96uDTI7BwUOfZiWp45n
EMMcLosg+Eepv5lhyxgB9eP/s10WBj9v8ES1K0Fa/v+iMpHp+sn1yN7YnLgi2oNw
lBAotUplxgjyssk/tYiKLi5CWtoBKPtMcVbqEbh+uQyCej8UKfIKHBErHafuS8/0
I9TzFtJwpR+pizqdcbXZnnuitMTXJWehzHRTRIDUTO9SQiRRJj8hR5Ii9NVzjlUP
KiP19F8yHikeP8J4xWmrun+EFdv6z0tEUgZRScHogjVn5U66d/FvJacLKwKmlqoa
20ChPb9ol54Q3HG0tLiohjlOxvJza3j9unkwQWTSF7umGxkksa6JHIZa27/YYxTx
imXRkEPlIfmNvQkNgQDqMngfLJc6xG3EvJOUcdTX1mNVI5MLt2V1ObPRVEg50HDU
eqr4e6A+uBtmW8pgbzdN7pFdUZsMex5m7gjDRbbn+PQpgTIbve1oFl77n8mzJW4M
rzrk2inRfgC0SuHdWp1z8rr74jhFcsQbn7lg2u40enToOjNlT3vt4r2xneTWKlyZ
4DVxYNSwMBVHn8xjwFDmDrhLOiNqd1jnrUo63aWpSxa1N1OOwLSRRxEXAYIpg7/5
IsTV/iv4X6w0NlCCYXNbPOx7dmdgFzUjyiC5zWCILula/Ds99gLBP0rmwES8sANk
CF2vGzWD+Ithya5gV8v/BlFlPwTgssgCGWEspLPkRCYc8X76PZu0AMTA19lvsFE9
Fm9D2BLUFeB9bYUv1mfqB8uBCSK1tGMVAZQzH45md/HMDbGxjZWiFLLpuI6CrC2I
VtY9GgVwb7+9rl4rSsK7GZ0BcjFNIEwjCXok18wqglAiIhvTSITXvHrDWz972mjQ
ndh6o5uUD0N+6alz5PMU33mXb0QvbgxWl6/WKn7P75jMtJ+mEdKtaOTxZQ+ptdCr
EtmA98UvGnJUK8nSiBktodM7DIgthjXgMntlQavkpeZ+YoxCKMnIDXZDp62ew0ou
JpLatGsQUYnyA6uDkZ6LrS2/rmgHKz0zZH7A0uVBaTT8+hDIj27isqwPdKQ0knpK
rvQ1PtRezMhjqUgWHQR8EW6j2ND2InDzqNT0n2jEVQ05MJZGsKuQa2OAz6CgbFbH
hbqgLyLfaATNJx8dSdOWRzls3N6RkXCh57LuZg+oCqIlTiJmGhkOwHx5jzGMfYPt
BH+Cp3IaKFrshu/9D+bEvhFdKHhFa9+sgkGm/fM6hd9zWDAyMwJ3K/SmFVkD9IZP
fOlKQRyh+00fpZiXadaVl9HJX4tMYNGuDUtqwiXjyYpXd5QKXT65DoIS/g0n/p2a
8AGywDnGTtzSd3RrMwzeT2AmBAoF5Gv3OLqY87ixux8vkX/E37sG1vnDbJBoxCvS
MtnDQR2fFo2TtGwdoX+1FdkRvRqFq2zgS+rx0SbDugC25YahSrzvOJQ1Hsm7MB1I
CUSdXCaoHPxvHdyOXaGYHiAIqukpqNFThQXB9NIYPlsnSGqSc/ee1IJjK5bbd6dX
CYtbPggrKt45i991CRnYAe3nOg+hKdebRdzzlsjnoeSfylvlHdP13Io/dY5t/daF
n/CUmgcw3D2WKkQCz/Fr+F7zBPuThFEAeaFCBgW4LunOznBcZSp825RkXymHKrok
ezEl9IKCnKtVdlwPnOhdIRfUH9KHe9FdmIKC/JnqgIgyCbfBmGKHKsegqIgTTpXS
K70orPRDBJkHC9kMcBkl09j36UVuLzQRVu0fgLqhtupxw3rR8vAzy2gCtd+MbyD4
JO2R/2CYGyWmKIy3si6PFsGFhahAANOxBHBghid8xTb+V7Qs6x/ykiIZ6OQO0sOn
ez8RUPPoS2u5QjLhd8devatLMh7L0NxgXweVPBDX9NZJ+a6Hijw+bkFPfyFlvU0B
vXluO2CCJakD9aX4D+VT9YHEonwX9lrPWTD3gywo4svx5Tukcf+95W2vHxhFd2IB
ZL8wj2tcZU5oVsgOrR5s0JIWDAYrTF11FdlM3Nh9cNatfkpZWwZeb5aAPTPUwIWV
upMW+2muqEC1/v+J9l3/+/6mL+KVUFlw7sd9R6dn2xOt8ZjFeBin+1TmGdPFu3KG
+sZ5lIZa/hyGLO7Dlxb+FXVGX9i7nk86Jw5ZGKPXKW4djdI/xKAClSJs6JCJHjxG
naljS6BMdw41arnp+8W4b7brNJFEFD11v0JJgG86O72Vq7WZauJd2PooytKwK++g
UlNNVNezjCkBQVphD2BINhi3TBrtkuPaIqCLgE5QBvOuSO5IQmPoe6HlXMqJTHaj
IdoghlPnIUT/31q87u+FWIMq3iBoqTquK3dChSKPdIFdywOevoVlE1qmB+YLebB4
ftFbiFV5hUbrGL50QI59vW2yqU//76eDlSMnn1rpjxYar8giNPMP4m1QIeL+mgzA
nxyXvml3CyesgOuxEENmkSkIPtPibI4l8+mr9QUloLNRj4ol8Nqxl5x+UM+enfk6
1iA+0NDhn15yJxzKY+aYLKN8b+/AAUe9neADyg9VYFx6ji6sHtDMDPRAV2w39gzq
PJtAxArRyjrf4bJkYWNseT4pFpBUIDN9HuDEJP+YLumyYhjRqrID21t9h+ALycyd
f3b7m9ceO5FISkl6TXVdByvyud6BOkA4h+KOpa4VOcZhDkdc56ymLpuxW6H0/0+x
ZA/wwG9/A1goUybKQieLvY+k5KXSrx+bQORCwM1/pn9z/zybWX7VVhOeN9b3Z47l
e4nkpfGGUGI4SoShfvPgYhLBxN/TwvdhVMePIKZd+MCd6vDUlh0RVvCu7wnf15Aj
04n+dImKu4HLmy+xbzga9tmBEsrhLEk909kPGPioCw9DVD7q4x4gBwWvjfygrgKF
aqM+/LNhMxlRpxv+kAtG85IeQNSdf3ixU6YoDB4ZkId1YfDgijSQRT3Ybb5JXHyN
SaAWxQK4n7eyLCdK2dQjjzqOcNFGkUct1f3NwHh9P1CG7L8LnpqH0R9sGtkryBP3
xtOo2tatidz1ca1xyYjQqzOnYNsP4jxhbEmcAyBbfrTkyKwSAD/3m/3DFooQrGM9
lPLdt86xh/qPIQBtoXTG7Y8caHYeP4IZ3fftE5I6owfVLmWAkNH+5f0i+RInpMhH
6QBWvkYghOsxDVbwvkOo3LeI58XPwL9j9Y57p0PjXSJvKkamczCqz08Ry3ZIeqmK
qjNUd9BgZbNSxtGkglykEXFWyrAxJgG8unPWBpCWgmqq23JdWiDVTDwKV8dru1rj
zPNw9G6B7DRf1MEGPQYZF94NoDy5DKCDyglTv3HdAAQCsutTHO5zgCvv2aWugiy8
Zw6Y7mrWoi90xNBJO29paUDlxlmZCoqvETBtPWrAOwIl6WqfXGMlaEhJ72Ocw1CO
zQ7eAaq6Vm7UpOttr9lGhV8pc4S8ZSlUBrfm+Ht+d3dHjKkDC1EFHlixA1iip/CG
XPAt+KRpq1soIndyDRKDjKQGQGxwB+vspwoW0OGHkgX8HpXBhtwOee+1C4Yf3ONL
HtugtFNwb3PedX/R4ijPdgR+ZyXOoIgXkYIWcuIcX8CunN+oZyxkB2dcDlilLHht
MKbJhepAQXpLmeKbjLcj4qk8NdfXg3S/JsW2kX5Ge4+HUcEV/erRzllrL7RDvHKu
aI7Y0vNEUrxtFaMjG0B2IRhWRhVVip2HuD3ixvjoyLDJQrnR3w/w7gZR6AVtsVPo
GsGRZDzHfK/YcFZzIaUHEWm2F/QJbqp5U1WOLzQ8dYDYQOh5hlwbi+i4bGme7B//
hlLbYRETBiESrejunfvn9/1PrQKFnfLMn5RZaZElEmIVSLASzJU3DZtBwwHLPPqA
D0VnQEeBlb711zB/omc2xVa/Vnnax/kFqr3nZ10RHItQWrOJd9k7kAI8FQQ2qTP6
vYiuDxyrtz0Nwp0pAq/9dUUzZDdgb6qi2mIlTIRRn1+zUVDBaftqq2x7uXAh95ul
Zo0nvhdenALLopy96dMwWTSxNViuFvu+uQrqzH1yxW6MDZ9Tac53KcJ+9DWBAwrA
VgnPFBhNyDQoCGD28ZgJZUtjX/+GxC6+f4IMJtl7TwPy6L2PQLTABt3hI/6t+0GW
7F9YLXW0FgHFZx3mJ/Ube5ciZn1GNIf/6GxS1Y5NiBx+fGg9mvf9m/92RKF78lMS
Q1Ywj8I/KEJ4lpQn/eIZ6cwmOVOmOFWdiTL0HAgjufdYr+/xjA4hMdaM77LDGnB0
1kKYXuJ2BQ122zHIwnDrwkPZM7g8KUpFlJGOJ4cCPdkUk1iycLifsm6DCVImWmbt
4BpQbD9z+fJqEeGlehvMm0voXM1tiU5f/D0JbSdP/x6Y0XQtnIp8FPavWHFF1n/o
SDqWJqiLknMPL1ouW9gF3yrMAWv9UqehsX13p3gIg+nrKrkx+i72a6YUELF/bjZs
iybIv/4Jm/VJS/624m1ZyYR4VEVvOzeLtjgpgiAOsJIyxfdkkQgici3+G525V2Ch
e5Qjvv2aeVcYl/vKV1gG8V5MA2MKkFF3OPNoWZ5FdRK11vBuaw/UlTMsGuNv4+hF
1juPP4iWWvwC79V3x8NNgiADhkn7uwlPX8/RhuXb6R3bhjDLxiFitMLuChbiMlhI
kGQ5fGNsyWf6R+GZQwyRcZ/xVQoHC+ZlEbmJnBtVI0qrKm7afIBy7yC/T1fBX1nL
fakpdBoUOcGct/j5eIp7Y6E2u67tBs8eNBbIdfCsyfFNER+D9ohv+aYV9Zoi6xJd
gKscXGr/hvTFHaamv3DB8l+bShS9vcmRqrnuguIKa5jeOEygjCQBHb+or5Xlv8HD
fBksPvzpD+dlW9JMvAkkaMqYHI5oZj7fHOr7YUONRcyEItMBhaJIr0H+BrYBds6b
T3ZbCnxaORjMMCnl1/rAkSzhuHoPMk0i6gGb0alaemM1JpI0pBdS4InEpVAElIsW
zDHoUJEkl3Yt2AbE5J0xMwZZ2I1BmBDg70DCsjU5guPte4oAQgYvYsvx95hSyS+L
HSwsq+dDcEzCaIO590sZWyAzRdJlIiC+jQFNvF6KDgKpUfN0Jp+OqnLVm4dTH5Ux
8kU2Uu1iwbp3L843L8IxHukcz8wvFuQTXlOfHI4YZXefA3kTVfc3sJsTSBHrLViH
gy0cQpqgAfa94ub+7kbDym798/Y69H/caK5R7v0XPecRwzRYA6IA7JJITzGozftq
0505c476XnA/H8kh+ybe4zdDTaOFT7jHdfBhmcVyK/H7rmIvS2i/AUe7o90DSExV
WP91hiLB/dfmlBAqWMy6RewNykrVb2H5dOmAICrmneltDXbtftva/JRV6yPACqX0
eJFdO2Wct1IzGdl/dan7SxzXGcGJR2AF9F7i1UNWKUh1tBx1uZIL6aCEma7bwOb6
iDMaH3msRLx27bZqivtYUz91JMeibaP4Oc7FNoXTQrOr+j6HcABuRm8Qrl7Z7m/x
+frWR69h0jRLw5c9pNrgdAThnyxyNXOBx7NsFIojL/QiMbMo6oUNgaF31HQrFcnJ
/G6ws4TKiBd1UaaIdNBWqK3Jr8zocFwKdG/wOPb6IdfIBlxI7exoXEwzC38m8XtM
5K5J0rW6zNNKrgq1XukbKcElKgkO8W46JS6m7vvNzOyV+19FZ+dlgULA9SIk/HM2
gjoA6iK3waclddtALcRaN1TeANZ568SeNamo34QN5kcHuy4qko1/0EujkKrk64Fe
H5+XLxUCRIx9iY3s6aY7co370woR81Ye1yJw444lhjb1Yeqp0QT9ZKmYT05YCF9B
QbcyDI3ZanUGePqZ87bR4nTy3paGqtHoGMsgnC5uk5llVaAWjkWMSlMKxZvy6Oru
ZzMr/xbntzKJet0ghzw0I6oAVTBzzUPNr1tCLDWvfcJSoPcwx2Z34c4qd6qXegmC
tYQIE4Qgah+5f558Qt5fpnvtYDUPhO485F+HaTExRzmwWIRXNM6nEHKXaYKw8QLd
omlgwY28lP/gbwcNUVBdll6Yfp8pQRMlV4ohzeHHfe6dg+I3HKKONBUr8AOMbWMR
OD6yodRmHXZp8SkWiQY2yiIygLA7+Pt6Dxqulguc0cWItN3k8zOgTYfA+l/tHP5y
lDfqPCE6UgMXS0/S3O2hUFUfdHytKFIW+Y360GOHS+z/UCk9PXi7HjrhpPhT+2N1
O3UQb48Ak2RzKq+CC1/H4nN7yfmpXRt+sIBpLLx5BTKsIlqpxQsFO8Ozh33Rr0p4
pp3CvRL5HFIgb8qiQ8G8uBH199wdu8FFuVtPIcMUddrEYMxDSjMBvAANsrwUNeSD
MdwJ9Y+CB37Qqwrz/MKPV7a/c7hqG3dulT0QFwAiwpgEwE6fEe5GTkk39yePtzpO
4vqsqlRKpFOFz0JIuiKvNo1VL0Kyhb92VnSLsFdEJqX/vIeVSv6BOiKad/fxaX4h
0Ds1xzt8UNLFgcXWvQYL7powJf8DNvLtwElzqc6rst9h08gXIZ3mzrevr0Mubn2l
8o37Ly6lXPFPnIY8eMe3P3Kj5lXFJ2yLFjxm4+ngAkE5bXIOJNa6EBQQmk3VUQvm
dJsPKvoC5hZMXAShurZ8JXfG3nyVahDKSjryR8QrEaZ+xnuLW98UEGHJrK8azLV8
z6N936BUiPTkB/3RTxwULC9Ahnrv7eu8nUGVC1yVgBN7QtMV0sRQcyqrCwPA25UB
GXFIx0JLXSYiUt5ZNKLtaqobpRt85z+szxS6vHwaMl8t/PrEr4yudSqLXrxIhbZK
nHMY8YrOuc8iRyNt3C9Z5kgsbSXvOAX2WHsmRiqzMdwu5CYcAOrz1Rq0Pt2ccYY1
fldLbJa/AE1KBhuxo2p9GRsV513/iiqMHxqT08FQj1JakOBElccGFtptjvdKYFhk
CuXnQCj64YKx/KwxB2oIKS2IkLt6I1BEjiXHwRSdQYGMREoZ+gbcKPMp2JYBLs9y
HFcsg5KxE/2imRgUHBJonj0g6ZYMw9GGUc7diH2LYQeC4hoGCyQjtHhuyQZCzkcb
5dUDfpj4doP/iLiFi1mtqKmE+y8qTwNuP+oY09ok+x5w07KuK57zhYSfcrVw+G2v
lwMr5M36D+IV69pdD1b3EKC1yvU+RydBjTt1vWz5Oakvs+IBIJ6iI7AhFmAzX6oj
FohNPNWMjgq+bkaMed60FAaWrlQ+bLiH5cQTbcnchOXV8krqn5OEUjKxTQMZh8U+
K5YlIP3aO3JNWZHa2wls5Nz2e3xLH0c7blys4QFUGEB0asYqX/vXnruiKPXrlwj4
GERGLrqBR/9Ex60R0D6mmbnjxyV6YxFThxZRf3ejOKNgacG5pP6wGhyMVAswLWdu
RV+sT6NbyjbSH+WeiCBfWVWrDUrmxSqy4DhwId2GD8NrGDdadGAmu2GLWTN9vL9F
Pd1lBxCsxhRSwHHGtZZsGmMzZRVZKPzMG9XPSuFCFYFdqoyNJvsXSfZ8SdtdhH0+
UvojBdum4c6mrhZ3WpJVZ0BoRgjhse0ZaU25vBMmj2ztJC62Gk3JZ/HqppHAu4LE
um/fn1sf06I6uzhv9CEAa/7xfsuGD0IT/sY3GP9IrrjtAqAUnQ4FvzmSaO4p4ZoC
zdNIZnYSQNO5fuGVB0UjR/e1CjdJFgWZuj6r8hKDnZp2B1kz3/DpjIeaaj1LmuXL
5ujz/V6f29GCm9r9i1fdRmTSsGEaR49xcfS4sGH1MHMpBj/Tw4mrhAaInm6WdteG
7OjE02hHkt/8r0NQ4f8qvhXbB1gtiCLkl/Ls+oMx4R03PmUY7XOYENfaKoZdBd+3
T8QjxMg4DgjjgDYuKytkQ7S2PM1KMFws+9KtMNrXWZ4rXn5QGakQgVKBG2bdUGsO
qMNwjKRUPznpkINO8n1uELilUR/51QaC7e8BzAhYo8JlZVa0j0Ncs6fVZfzP7bXo
qTw2dacpASKVZJHA4wdciJy8hurw8AGRnK7bHmfwFkYAcGy7fJ+1ZCgqJEBnjnmx
6SoctiZDEdqtUu4fdDk2kFqyuQ76urRqnVIBxKoBkj8/BEi0xzwrN0yHi9tXQDq2
FVtB51wxAe4kdqR1tP0Htczy20SK3p5GpJTMC+iOqAh4H/dkMEBKOvG/fiPrHBty
`protect END_PROTECTED
