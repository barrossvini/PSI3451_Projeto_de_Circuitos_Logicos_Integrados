`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DYGtQ6l/5ir0Vw/BBdAdG+Dhjlqz1WrjKygP/b6l2SHarVWKlOf6XLSC+PMKN4HH
m+NBLtwzLvO4esvC/9ny0yvs9OiZq+RtflwqAGZNDhtWlu0GPCFcSX2aTzVDyK7V
pXEKwXpbYXiQfsN9PTp2tF+PX3QQ+sF+G6c71ToPne3Xw7S+2LhiceLMF69CxvvT
h8bY74AvfFhhUSu0q7Iafq+zvBstSh+NdJl99rgO3LCh7iKiVGrMkIfzO46XgRgp
ZqJfRc7dXhG7KxuF5Rkdlp0eB5a9Ga/SgFFE5+tXk2TTg5p5Gtrag4Mb9OKSmuZ4
5TrwfjmV4s6N+f5lBWIVe4kZbRTrJ+R6xYQoUHcRLvc7XCYX/9Iot7brsfoTBIdk
358/UVJrZVRUmjH4adX/37JWf6XJzVy4trT0A9fJmSsJpM94czILxv4XHF42gwYA
`protect END_PROTECTED
