`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K2JTK+lW5QBd+/ZsISez9iCKob0wycMQKpW/abou5na+wI+Rh5CnQ2mesEQfNUNF
/T1ZjEWqIeZVibYsFBZ4RyoORiQ9NOYAQDd+GSbcA1hW+xNbIYsoqFsj0JA02AdG
6LfMG1SY8/kqGc0u90wujGsF/VyVneSpGf4hcSipUH5/RWsaz+CG++0bF/149EXD
x+e9meZSPYwf3p2RiqiPyK+NPIN1d70ggiYmRVSKb1z8nMasByQcizoHbywzcLgi
JHifyhgH4cWFpgIIbXOwHv7w5L8hJnxr+PFjmuJpOgNTudS2DMx+d+gw+nvpYCE2
PUKizCLPcjK1/u/gMGanVZ1VwWLp9DRUeOtwgAZFRiU0+jhe+ob0rhB7/PSucV6q
r7I9CJnmogr/c/6VUUjiS8M7qrKLyzFipcRDksY05nscWseTSDf61RojoUHKz11p
d4fSP+4YzF809WOeq/am7debv7p43KRhsBeynbxWlxed+q6kr3KXW3ksDlXRU6/X
FLo04FmRNjLCdHlGlRnfaoq2djOIbt4oPJyGMMzZrQKlDJrKBzUw6wqPm7ozat29
9IdBuF1UnDzIkw6FdwLnObL/tJJuZvWeLe23USEd2oTs4Ab6w85XDETlzvpj3F2j
7PKc34UtM0oYuxhzywq10ZWtbC4N8+bRPaimeRLsX7iqb5VCws0kqrizdnokPV4J
9JW2AEn2BbYn0mHR6zgzGtO8CvDDhuVYeSdJpFrgTw3Z/VHGbpRxcsYNiF6derOe
aRxn0FLDZs2kQZsz43v741/56bEaTG+c0dfwKrLHhsl9VIrFEsw3Z68MgB/VEBNZ
1CRdkBJSqE/f0+RFBm3OZWg9gjpLPJ9Y5NKZpJgxUZU2UE/f876PxNi0/UWDYOmF
n9Ak/ben626c+umtlF9Q5JdFASMEDgDuQyzMCvfuId/gdFk3tytsZ3MyfOstvRkr
TP6kobpIdE+8Wt2TkKoxNjsHkcvTbctbzNNygyvxT32LD7v285HEtbMa6qZ0UCPd
CBT4OI2tFZqbI1vshzQGDwyRQJR2H8GRAHD/1fKm0wSzqftelU/lz0xYjnmhb7di
HM5SI3JKqFiZRhx/WL+CTnS09hIm0XdTCU+z9Bb0nsVsxI0OrhKBkjISsV3WLf0M
1jmqKBrffc86rbn1FzrV2P/nsCRGpqSllc0cLPwb8NZMuMoKt7SkKJJxFo2uzEi5
ocHTLo/1qctH//nFpQXnm8L5GeP1hF4zbi/54ck7wCfTW0gjVzoi3YMSMM9Eh7BF
F9mZaiI18v4UZi3mfLyLFcGHgqESbcYoPi/YzZOTU+adlG0xq7jjlGSoa1/4u0q2
fM/VT1gYZqE7cbE2Sf542xsy6wubfMTgPO5dR3zOv0g0gC0lmmnfbwOJTPsJcdz3
Hl2gRjjpPq9jEw/FGqd0KLzC+YgTmr5kdK6OIn9h5Qq4VsuF15jZpn+IlG63xi+K
m/XF61dafUEtvhavmmy12JuD33I20tf3uMakPuMDdV2IW454/kmHTZL4J/61SNRO
40qTj5xmvvO7QmSUWC4cF9+O5cHdpA5Go1KK1UHDV7kXlgHL3cE1wBpSQBn9kiiD
EJI7CLPWySWRocmGlDqQGZTDQpwfHVqrrGqpEWT9uZG5aApbMaxRN9vJKJHKISl2
jPCcpnNNNN5nx+hhj3/KLqOr4vfP8r0zwIya/lmQN/zHx3xGAyhDIvQM/Vm4YocM
W+wBpwudvF6pgeAvYtVTXRK/Yqd7Eo2i+XX9JWProanGYvVVaL7vrk6BKQlcXHn+
G7BnvMavaULMMzK+T4T04+UNjpna+J3LhtPmfIAxaOCitkYOmUt4fxRVO5Reel9x
7d9ubYWu64MDfHLeFAES8u+MY/XBOYGp5Jvd0tDo7WZ/bnsRPRL+8mqBskNNCOZt
qCpd4GMBMzx31iwU/x3MW6iS6qB9exNo8I1SiOOwEr2y4jt3/SGcdelav2toRLi0
HnOmMi3wqjPQGXBZvHo9bqybjEtPKwJRm7lC4goYjLEcSTRin2QFN81SUt4gT2Fw
Kpm2sqFtrkZ89kOISQqL50j6jPnNEkF5Me0e+WDZrOF+7vH4EyR5+I9uRbdbXEpB
936zN0gxr66bIR2gAzW2Ead57lrSRgnJy5GavKTukXOtX8vCdx/IoaCwi2S/ZYKv
FCqxyJC6kVxEC/Gy9K8r0fpvMWDIwJQK16ICYbZAB0aU5tKiYNsis6gZwGmVVaTO
4sw6bQBGMhIj6e26tE4wPxUciH8ir/8Ox8BUJaqJ7GKdY8uDwbA4YUDQyTReo/yc
vJf0S/bh0N9XvN6h12OxOi+bfOImZ3v6ZbprHT+8Y/g+BZC6cZGUWogkvnXHvO3v
Z/1Lj6uRBCeHSChpyaMJaFikTbyo/knWBIzoenaHzhQ8VEOOJw21CoixK77XeeIG
6ySP2CqoglkOX86FHGgUBbFqFcgrpJ9uzZ8WZFNjZrkcSS3oiTwHGmY6UtTe/BGn
IuL/bXKhNd8RTHxz6uFHqy/9KEnr05j0VT7P6nq/QzQKjlkrEzdVLzQ/brkxASNQ
PMQ0NHTZvC1f1AaC6xSHu99vcBJ+B+W77t58xyQ8g0+z8Q+qfHFYxS/nAzB7o5eS
f0p/565BxTid+xZggTPEFuDQEn1c1kGauvqYB8RsQt4HoRRWjxfebqQVU0RqEDpN
p3P+WOw8s42JD8ylozvgD7ltiqqSVj1FVlGRxQ/l5nb4andlwBjIXsRqGoFLDZ+i
ijmy2Uy0Puf0QYMGoL6qfed4lzthgJHonc4YuBKx9xtYq/YXFmzGJwYQiFI/Ex4R
OFRWGcKY1uYh41NzdjtYgoC7rvLZaqXvESZg7UhqAitmxPtVefenDm14Y8uDXIGA
tfNxuIQpmU3I5WKYQ6XIPa/puk45suVYkN/5UU9wB+9etoEE0WQM6VI7uEDMlpEd
4tJ/ceJfKwxpSQF/clquHDBOFC8J8ryeudzDyK+bfHM+ko0NrRnLLXWeLeJNMM7W
vK7phooBSlYspTzLkChlaVW5Ub207TYqEz4Xd1QqWRAeuSNR/o/5qG+xW84KP+6z
zl17ISEAw9d62j9jOxMfdfDbPWFJv5IrGrjK8QqHK+FxyUdOefKJK6FCYmUmCVHN
8yx28pkp/F7rKRwjPPNddpFOymLgGxt+nLrgcuIlEQ1Fg1BrWmwpKrXcRFHw1E9u
T4q61Z846ow+j5uq7bmRsyLtoVKqefOtdUT3plSemvvdnfecTWID0WaKxP+uXFGt
9kGImf85WSwAkJaDS+2ablhHvLjHJiGLx/00jVIlvzRUjEQTpnHB7B88N2gLYTpf
FFghVZpvv8w1fb/PjcThbgoQlc10YuJ9/C2KhISENBloZFipHF8kidlUMjrrxjGL
eVLYsYKQEuJbFATkDAe/nGiHys4QMK3erAkFZOrUe+THHqAm5e6EAvQq9Dbk7vnw
gaTBjFYwLelip1iHik5BPwEUqPdYZqi8othoCuGj0alFOGotJKUY8l/jXJ7gPoRV
OSFL5MotBIo2nw880Ndr2JXn7a7ZLJdl1/r9r34m70krspa7AjGrRg43CT4PygKT
uAdedlIkBcaUbV9i3timZhA/UjdWQTsNoGj3KqfUSzNkO+DC6Gv4en2mLO9mso40
E9eB87c7+jHE5XhgVOll8sCDHglX+vg8QiNAzf5UUR+KcWU3hhzPF8/RiBKU1qE/
viw9SpqLhIxSRQ+ve200lrpZx/ZJwEhDlZYfd6SGglJBknK7fUVfBIJEVhhDjAvL
ZKpeKOMAMXzmvr83wl5bP/sJ9a/Kjq7BYC7ROiU5IsVuaBg7n8cPfxzOZyO6syB2
7Do2QYqIXg8ZteKhkjqRgiYV1lz/M4sU2FTQitljE1nEGBSxLSJbgPHI5euuCksQ
1E/6LDawXB/zgcp4Cmkbq/FCXmIBr0cJSgYjxrx6ReZ0cH4Y9/Ab6UOtT/AkCKhS
HNDHCFcaw81RjEN52Jijf6MYk1yWvMqnN2XGZpe5ebnv5ncmMbFf8vC/TahhsUu1
18BygolImIg5NgOL38rvOzUMGovGkis7elIylov0b/+EmBFjc44+loXNjWqjAUP3
yBPSJs0W6tAgnp29VEN7y8+eH2v6mXK7FtnWfk2o+TMOevZ0/W6oQFSTKIPUS96+
azl/yc9SLujFYwvUqg9N3gao0fVyMEbC0Dlx5iUPw6+Tn+7ghWVAl1hlXm5Onon2
jMl6r4wu0Dyu+j40eti5GdqIo4d2KMO0C/jv1Y80jLhfvflomNPMAhVVW6AHDJ0v
lYEy7Ho4KlncJ0CZBjQFCHcS3vXTONv6U2X6ohnbKD0hHwXc3IriJd39mSzRr/ha
Nw9P6ktAfYSoankj7KAo1KaGZ1dAYJO3PDREyQpNusYJZpuimHwNm51MCZ1qbHOF
wwOF+o5nj9YNaqYRyhpaBJl8dKIC4ofEEN1A6TUOkruiOhMniNVtj76i8GYxD0kO
ynX1eYs0MQJpLM9mdQKIa9e0oVLp6WIex2XTfD7g29o8rssYLNfRJ0NfTykp+Djs
iWeCBD2KBgNgSTnAzfx88zFElBOvChST+wVIafI5rxhi5qDFIg9keS9Y3m6v5s2A
LEMX3+Ypm++Im8xSlJqlnrLibAoILyRK8S9/CcAMbig7Taj98GKP26TMS3yOuX8L
mQF9i1vadKFDBTQujm8tN0XCDs+M4vh2yDDPM+DdiBzTe3/pucux2GQTXWrN3b1G
iV454FIkCZONgQyp+SevNS09rcPKriZey2wW7v1DNMzA9IVwPkeZael8Z8/kcv+F
5hLezUtnPZz4+PjwdrxybCopJL1hfP8WYHfspaGlawZJ+To4Q2Co5OcSq6Z/NLyZ
ESLrW8DBw6tYtOanuEE5jBFA+4SKo+wqvWjfr7R8lIjpwiAc0RGcgqwMztlc9NkB
Nob6PYy2GOeOIOL12LmSP6H03HXFJOY9JFco5cMo5zGe1a3BVvPzRAiMzr9xwDCA
O1Va/FL//gyQ0yBgqV6uUB/zuVCVq/DwzptCFr9svsB61D1JpsDUo8upQf2m2eyN
u6h0gvT7xxX0O0UB+n7HcacsOyBDktGjkxcUqUd3hftXsg9KQ23QIhqjs/6AV69h
pvFwd4wAcTrFVn7yP+aFQ5u9ndgjJgroWZlt+HGkrvWgSbzWs0W6323ofPr7deBt
+SQJ+6Tzy8dMbTbkpIIWci+whqfp70oxr16XfILCILIhKq+PNOpQCLmsM03fUIYo
81ex68cd64qeXaoteUa9Oox493zra/izuN8RMfu/8Xj9soPYi2VSOGUZJVlfseKA
le/61W5FB77h972NhetF2tasMg5+lt5Zu2FxsiI+WZ7pfnecOSUJt6T+fz/MxX4h
AISguJ6HSdezDm02psU9xmiy3idZ/aAkvzuTbno9y0USZihxFd1LbtfsmPv53zYC
8fISfWTsX1YSFF7XGJrZfglPZ+/vPS9IXo8ZZxytG6fdbSPY1lhFmdQYvRRJ5CuG
faVzkF2irRAHGfJJdTchur+3urQZqj/TaXMonCj70e7kysFKFDIcpTyHILF20hvX
r+9b0pJ7ccPKpSWYvuR0IXQAvzDd4hMgQED1scCySqi4eWrnDBnM/RKlAMVMOBT3
v4U4VASaE5ey730Kd6SjUJV05nm5owKaEXTpOXdr3D2kwXWG/+SwnyGiAy9MmGHI
0DgYkEIAVb3gziAs6tSsczeml4ykxvYHaFvN851jaXF2QoSgbIoYh3qlbv2k3B2c
PqhopI/nLVoyaQ7mUr8GzoOmAOkbaqRy8v7xMDhYZtuBT9ws/agL1EPP8/j9eFb/
tChj/34cHxIIBSZAiRjs/xR0Z6c5jR58xk11dARnAWgDwLP67tCAuHR712LieHgF
RLvUzbGGccxqT2TSRGM1pG2Jun07CXAh0U969SQeqGONGO8MJs7LbYdHb4vpOGb+
jQY3yzMFDgrggX+T+Z6N8VXSAZ+JF4R9bSXsJ7ridBpg/GTdsTVTJPvtpsVgrKKU
HJUEYjkPf0vMU+AoN9anPSoGpfn7mHsdVzF5rUxXAuT19geyAnr1MQaBVxqf2/8y
rguSPHh5WgkAqhh97lOkgcFZg9twiXXWBJbkWKDuPOUmJD/ycuBGEQLroqSCm2RY
ChgjWGHAZnmO+rb9bd+j9g0r2n7+RaiJm9aUvFPimCUaGJ4dPiq/poFiETwxOCxU
CVAOrJSWwjqk1JmGbsx63cHNnBwCYu0ywzG5hvrtcs8p+ze7NNridU/cZSr30DKV
SrfnOJBXL0Pe/7GZRFnDcQDV2vNmBKeyYFpfMe7ShVbnAdASIT+fN/73YCzoYfyu
KqL0/WI6kXebvDzAGkLmmoLfEsNd/SOis1gOwfLrEm6lYXoOwSF1aePCe37AoSFB
IyXMtICvmr8xtcW+LRkaOsPT56hJMXicosqjJ8nXUtSZGpfShiPr1VcfPpHmjl+N
NJQecCA2rB6/zsqToNaYJWAPx+6EpxeWA9TP+3ZBhIW9eSadrWKEFA76VU6R4Y3o
C7CK9BHzQJL+pYsippE01UmYDQSd9PyxYY25HBeRUmJ6H97aUgyk9ToxrX7C/89F
dlMH2qvms/h73iZAWVHhq404+heqVfmT3hPzD8hGAmQQmb0G/IDgLFtVP2mkmSLL
9IBlvMZ2QZr8i57P/f4pep8EOOm9W1c8IyirjiTj7QnOFXk26WbsbgGV2g+ZYh7K
9PYHPQDn55UVhwpXu5lhbTiT8UtS+HWdbHJpkmozGBvl4u7UUDu7Sh4glGblZrSg
582/7C7G089zUVf1bi5EfpKT7QFAVb2dRR46Io0KNY3EM+hraqMRHUqzNocSNiCJ
eRqSAwKidlbRJMA8PmdMFQdrCldcv9ldJQZArDykn0i1l4AfbDmt2xgNhNDMNWli
0ITlnbdi6Tn7/eubVgUhPByS5wfdC4THHfTgufMy+BItYRooxVQG4ELZfbRznbTP
l7m6IhP6t1yiuaAnSJqILa70O0T/sUf1/0z6ftCG6F3pFQhY0EDnCuH5sQ4CqvzH
6KSYx+uAyY/7o+FqfPBzs+OmDtPwlCGaTlclkUjb/OBzC5816Wx70AAZpf2yRxws
wSPc8jojMQgpURFS+xnCH0f0wXF4cihr+1B3J22Lbj456S3oPzu/rylGfRJFwGca
NH8hrYZQ3gWlRSBPary35E6TkiAqRsv9+XeqCU0VnfVky0PB5d7H5Sblb4PyPP7s
4E3JkSydgv8ioQcislI+lbwMs/haix1V7/GsjTEWw/EfgX7Gc3wyi5T956emxX+Y
pXuuO3MZVnui6pDvQvaGguwdC0G1tFsq156QlFd/J7b/RvO6tBmnr5q7nz7xzZzI
5XisXVp5fMZVmp3I8xabG9DdiOYen+uwVhdS3B8cXrk3x+TyJwsFHS5oSR/PkowY
cOHQzdBWxqnCbT/mPr3Bq2Hgp6rj6+iKxTWfibMoZw5bGtXAuUkFPEdBsfCwazJE
2Z1/tEiiXZwdKHa5ZRx9ntGyPw0q5+yFfhVJbY/MfVCZ3eyTZXdalrFjkvopEZnl
ozc5Sn6Bxp/qe49/89nuaAhlWj+k44rt7i2bAM+jbH6ePOVljo2VSCdpqooV5HBR
ueLeTo36QcYzS/JZlrNDywbX/mW9Aee0vXWylGuz7//mnJc6B6ryI2z125YqPqKZ
L619mBiMyA/KHUL5RQwsnu4Yn3Zaz6qYBPZcpobKvOUA8MjH+RvD79BA+ru9dnvj
9l38vBMFdjamCFAAI2m3ibRigD2xczzLtmTRlY308XWsOWQwToo7a0EqW03ykGMz
Xe8F17EynTj//mfUWzI2ktEeqotwIKIcUK0XU5eSbimfHLREz2DUx/+gWcWnTnCO
2PRLomjZjMRakHHMKoBk47dtZbKy5QL+YrPPjAYrQP1nRROsmRPdZEwOkoWDlnUD
6292FcaykL7V/GRG4JQkmAcysX9b7PZy3eE+Lo4OWsDZti7qdVE5nFPpe9POutOY
qEJ/s1E2PjxjVB3cLDbSLV4wodCF3crkWpNELbgM878BGwTLwkBOBVEaQJurIxrx
D0qaZAdbQfX8hiH6I6ZAWahj2U4Nd75kPzJG1tI6r+w0k8qydnhkus6rOP4YutX5
UPgFh6S+y2y2RFrAVqaG1G7fMw5QQWiD5G2pWxiold6WxyaLkMGrfCGQbYBygyJ1
pdM2R2SSegYnVROAnHJFc9JMaJrqr4ZB84iPdTvUJpzLBF3hbmHARSNsMxk4PSd1
/SR14vxEakv55NubCJ8qLvckTL7CIPVuMANYxLW4ZpNkIjjXeEyhvGTrTtcqGo0N
5OcIHbOT/WWzujTeLklHiMS1L4AR7jrjkSGTHGc7nGkpRRoJfpvQisAoE53ktCXP
dwuSUjao2UL/w3mldNOaGV2egxqx2GXLZ4eBlwMGUMx0tfy8xoAe1pTDuai6Rp4k
h8NL3W3D8fX7oyib3BjbRxm+TJhamoPAlbe8emJiGmo3JrTxOmZu88KqzOyX3Tca
Dvxo847YlxNLyoEByIwHi8O4c6ZV0Xkj7AKPewi2B7OQwYtVF2EMOPMVgPvV4Xy6
xKrOYtWkCpYT7Z9VZV5Lpkkfi6jo9lz+wWIlGQNhkqFFxtDbgRRzFwUGMzmFPcsC
KoD3b6sBgHO/uOhbg7tM2plkisTu/G4p3RldSG+UVSxtt5bLtYYc4/Vk1/NxdEMB
HHLxx5v63Q6CpX8KOKuaU/ovNrnvrPG5CqZdzmVaJtMgiOv1C9B5O0/VSiZCrmAE
DjgypTbMp8J7cx5KLYRMzWmAPMpVM4dMmrlja22NGFJHGp2DRlOUDozjQHXqxUPu
ZOwL95V6aFCKaee7NUVUGy2zzzz866iu4ljUwzyHPnEH5a7pn/9Oh6whJX6QHmT0
u/Gpt0Ph81912PhmE82kPlVmE4V/v7V6Q3RRrY9oBH3LfipB0V7j2qwjupoS6wva
POFTT/D1LsGgG3gunH4KdRXoQkNREjlHxLRd0qSmbk+1UlUtfryiAFVds17Olos/
lzTaCQ75TFlD2EdTrEsnBaePi/5zM8f6ndYjHKgxTl7NoiWIzvMH1Qmhj4jBQT9n
coBq0AjY2n4rKVrVnZc6+AxKeisMgEidyYvyyG0c/dJsDueigh2imhRnGfSD1pF0
PL1e2EPPPjB+s3Mkc0QNXx65YMInER2ym9TC0kW+L0mmKpokj2bm1bVrydJQR8DF
zBDNodYAKyBwLWy+tbAcypylgzFMBLyNDgomW61PXMTec8afKBmFRQkw75rt1DUV
oJaOTtxSRGZIwu4MZx7Gv9dQ+mxt81l3nOxjt8yjb8GohxDJmnlXaxZ43G6UAw0q
owhTAhu+aOApv/uHii5konCq3HjHqERay2CfHRFNXbJ58jtc20x4pcLxcUsKPuXn
s3k97+PeiFxTnlPBYyeyDy6DT+UiH7RJwkYhK+83SjcriWskvaZN3LZtPnY5Fe61
0i3cp2VudZfaYSYapipb/lPa0I9qwxFMFcA6/1YWeRoKMdoqW/myF5q1zGDM6azW
sYSjUpW8DtZV4rOtp/E9tmzoPGs7OuG2xyma+pn6b/PovfTAkgeAqj/fL0acjn3r
QTJJAEQ0rGQiw5oxj58aEg0wbYG6unCE6jAIUT2ZxiGUQ6KnvMjhqNLfMzWA54J8
cvYNyBPYxEWsH1PvXbbiHQBbxIAi3ZMEoKACmMYBDe2lxAWcyiPUy48RUB3DLzIT
y54reAZ031CuX6tmF11l2m11hO4oLvknRmrlFe6iyh2GalMoQhRYfT3aJjrgPs0l
1susEtY+haHAHpgPvMdphB1UAs0eLvopXHbJdLX52eROuL51bV5suIOPwSb/tI9o
pasw1ntA3OF0vuipMTAFUn2sTHoKxGI3OWQi7KGfKmMINRUkrVtBVOF7pGWMzslF
Mh5UbuxO00pTGilOUgNSnRdXsP2UBKBXjg/rz82bV3D96bgco+l3rbBEeaAb274o
5op3Xb2tSaMYAhtS5FoO1Fc1ySUufi1mVL4MmIXLlXAxdjcy3BWIHQ/ZWVzArQIq
ydYRpwsjS7eDMJPlvr/ZPPwvRs+23Blf0vGZXLKQxDABQvAGnKmiS5sC3Z+wDCQM
DgC4Zl1XpXtYCtOgtil0Xy7YXt/79NZaPcX7ns0HqmP+XrJE6G/WZF9TgBkKWJ4u
uB0w74PvRQ2euRbtPf+R3g7IQMQwi8R5xnYHGdIXlsKxo9MdMqSR42351yovnouh
fIubkGnAugiWQdNJ8WwQXAx0h5faW23Si9vD69wGMU02zLL7TV51O9uYxJL4sFjR
13R/okxf3oZxwtSXjxny8k4oVRy/LZBLFVw6Bz8sah9984LlFngzyonQW3KLOwMY
ZE6pH95szkkxAbj/ROzvIFum0x3U7iWfT0pXJRONZZ6ykL/RR3t4ZqyYJrVG7Smz
r73GzeDHNiaKyV+BDWljnfJupYnNJ7e5WghuaXftFDYBX9SQyQK8y7MPmhTJ8e/3
HQXH/8IcUA9xtLd7dttstC5B5fdsmAR0SZIyRhjYve33Vba6TKaSQDWm46F7TlSF
9HLguhg8hDq0HFtJ588MI550hBxKU2Q/x5Pvbqw+YBNy3ib9oUO6nQ84/QAWUzzx
6tPTje1S8jmrVp/8kw0ROBs/D3BqYUTm1WSvJul2miLW64PkHlc+x+m95iTmBT7Q
cqWRZ0a8ymniWvhdvDdwU3pgb3Q1torNJVP11Z/FmJwaY/3M7devqZsSd2mwyALg
LS2F7CWI0+YM3OaVvpzcyDe3WlWUhF34gexDrepfVxgG6kSYIxZF1lynXOdYmJ7D
G3Z8F3teKR7ka9JchTRVZa6BO0g/CP/WsBVtbuYy3W0Iymbeg8p0Qo5IxGMmL/6D
7AT0GNCPKG9W8j0i7F1eWFXfvgQZrA5DIE/zvzZDu/uxtIiyoaOVGiXPdKZ7sNI+
aWVgdFyVzCtNrKJ+qFAA1hC9x7SQoErs7AOyoat63m6lx+pIqDAUSH4ouI5qHN1J
9wg/aUc8xHtm70XnE/EYFYhla1uOFYEF3HDPNv0XCfekRzuBkIR7pU1g3Nx256z4
dThhgwvGO/3oL/X7IdYpO+KaqXtXj/psLEndsRkt7TUnoOxzLzIyA/1l9ZmII6DC
7LsLDkLVpBZrDaE0T/Y4MWYwvhd07EteUAJMPlle7ZWpD0YaoiYTUiWEcscQklDF
i04I68PfXJxReH/HINX8wNmBf0ok3sWKkOB43pfz2I3Wa9m5USgDVJtnr/jRKf1V
AbgGlT6eUHNJ1eof4/h5ZMEX7+97xiiLGqMy/kLFyt3iRLrViEXKy7XzM9KEpAEb
jNNzx38VKUu4pecei7QkF+dMAL2zZC6OjFwh35J0EaZjmQylKc2nfZBPdHKDddhO
9RKbizcqjMkO4tWXK0jA2iH0piQ0NjrTNARKXkJ9XqKRXbTYePIflz/NdERmOPsY
EaNnlPz9du5cL3asXoQsrEM0mvv7AdmPx61X4vB/r9dlXcXhsExVG50de/oQ3oeL
YHHZnSZePIc7mkKkdKS1T8pTzkg2uM0cq7szZq97Nb7U6DPKRoC4lTkqc2rilo4+
ZeBz0y7PSD29l7rIFTHhyI1QF6XPnpgR6NUw5ClTrAPJWTBxBVzYr1zf1iksFX8+
XevjpB5wjy4F0r6GUlL2mMDo2TxaCN6E0F+5CNcutFK8wH8kLzbLxQ0fyR2GCU9o
AWkaDboJQmdz7mFB8jWrNl90elAmx2EzuvZIBkiGCXAXsqX1pNHz3J0woXLopplf
PjW0azauW+V8ncRUECdhzTXts/5jgcorcZ0MUixBGT0TyRFrWoTr42lZAHMkVQuP
zfAxv172Koe3lLnFSE+Ofa30cfT4h0CmW57/Jq1Zcn6SH11v/xKGxTbsUsMB7Rc/
XXCgLrcMu8bghMpAyJ0W5phReVa5XQ5KifXxUP0oFvSltXaPsUd+EjRqYPg6GOQn
j64yFzNfhxkVcTmJ18Gcw5IMPahZOPxJmpRUMRvsr2CGxiUnzS9HHXk98P0q0CLV
fo8xZb0CHowsSYLNxhKjVcTH0R2/bDz5g925eGJr+9xbiary4U2qUcKBOMYorMrs
mTXfARbi+JOmbxbu9caB4nCvDStdf9amNQYE23/+ywvP9GkVpYpt41tRz6l9Ok4G
cBFWkIBO/gnIN4ch4gxcD31AdiqguKo0SVuA+At/xjg20U9RO0rCpX6DvlinK72v
Bbzk+pSxTFWQGYEU7/LfFPqal2ZiX7nLUwHhGRhJMrkM/TMz17JVKlduf6HZCa9s
K/650TcZL4WGbXIXxIjoHTBKlfeGL3GerYHmmhjnQNVAGxe6Y5teZun30h+PPfwM
0oyNXjT5FwMOTOeaHwirYA9F2o2J/s3viaQRGAOcr7L0wXW0WCVrChCwTeSzWz6z
TlCskVEnddxxPR7kegGppTSIPsu3mQJSwvd3yhhMuCIjh283wdQ7hw9R7HIyBSNj
KYCpEbw+ERmbd05hQiAicOkg/wYNiFK9PZuJbZtX4n7WY8dLonuuL1CHGgr3VhU8
sVzLxhhrma7LoanQia77oN51dAW620N9Ft4EL/+2EC1XsDI0erki+mwdnXUGwXpN
L9536eM8SkJiol+4O7kJ35FxIA4punkifb1IBdh/Sp/zRV6FHsPDUBiTP34kLDNm
+fduAALUGPGeHTAWxE7AIVryWod7Wqb9G7MKARqYQ5Qa0R8CcsO8/kD8Dvnxd3Ks
iyp3jnaVTy0AHlZ+q6MMPRbqwRqojhgL2s+m96S2YB/UN12yIpZS7z6f3ZLd5sjx
VOoNAz8472umPbJN6ohASHWw/GfbJozg0CzN7qO2STg/XlIP9Hxnwpa7loJgQJAp
0Q3HTSeLJ0wg13zLR+EvwxrLpdWjb2Xtvld8nYjKKW3vcj8PGNmhpGSFF+DkeylC
eK0PotzadyWCsc3Th18Nq6Y+kOIOB7b5ex8LpZO9lUwHUZt8oo6n+n3Pe/XSMA7F
G0UO1nfJCqB8nwEA7yHSY4OLuwNFjGxRh7eSPCzAdh7etHYZUWcF+Nf7kHAaTarH
qHgsYOVypIV6HA1GcbafnSfV2kwoO2gvBFEkj7CpEvJRCW5elV3y9VUMrOJM7sz3
B5glJZpl455rGA983cFZjbYIKQAzx7qL32Eu4a1XtRWV8xdqR/26PnaTmlF70ByV
kziBaZMHZ7Mt7+m67t+YQqgKGvlQ2j98Bi9ovlf6dk3lD323ip6fGJhwrhsEMiku
cHMSXwf/jOdfkPG+Td4xeXMZYdlYMcgAPWBOKS7F7D+enJ241sh1ZAzMyYoWkmiv
+Wto9lTOw8smkZmF251znZosuKvST9PfV5WrWoMM+9fylfyw8tui05t+YSGykel1
SlFDD0lIsQGgSDXTRIyvzaTtCeXRv/QV8ryXvSmH+w1TxNzOYhrmRTdLSvY4LUmp
C6h78V/SfbifhFaQRsteRONGhR/PXYvSczng+q1KfTvzrHSlYRBRXP4kIeSU0F0V
FXzLr5+jGVKNjudc8RDosBPvUzFvB5KavWO5XuNqNGgdRmEOyvBLNkRUn9Fm/pp3
0o8p3GQnHGJGMrHp9XElmvseJ51b8//mcq/eibn3VnnKotXtw/JDmajEIhoTAmco
OF18+PlZ3uudxD5Z/6b9fwqv6o7D/5aRBe8sU2dd1RP6nz2Uv+ZDtlDkV9oD1/pP
4aQNUhWert5JKf82bCZtGzhYil2i7sRTmFGb4AfG8dLLmtcs1IqT4J6BbycyPipz
cUs7Xf57k2Yv0pGM2mlcQM/OpzrixbxcXihThH1ZbVlyw8ogOj/DbbhLgluutWke
+DLylZR8gCEXXP9TmFBIv9YOHq7EafipL6N8iSxM7n4v+VVhkXIITRxCx/AqTCJH
HQSa+3+t1aS07NxcCJ0fRMfmZ1ioyJ1K1yae+6iQJQzcJxQsJJcPpSMX2ypRpbkQ
K1GSUxIaI3Kslq7kBWknmxpwJVAl2w/uUPGMl5rnYQf5dspW7jdf4KgClv12WXS+
2O/NOP8Z78DHetkSVQNWGeKw0UY6u6OiKCHOLieXIrOd3OnGQC7v+NOH1GF60H43
8g7srai/hggRg5EwSOzPbMP8FX0cNiJ5yj7Y26KfMJ8A9ogL5xF8GPLKEJ9FAjzI
FFo0JgovhcsGoII2gSC4hoS8MkF+HdD1QEEKJziR29IDo9evheQUb7X0Iu/+SmgW
KD9+dW/d3kr616KbH1M/qAiFbpbR5AFrn4QkXb3WRVWMnThOl7HxtVuhy1Bp/4wA
qKt9Pn439LxdQoY9x0kFlB2GjqYbWan4fgkPaZAsZDjSuba7KcwiIIj/E4kdNeqr
XAX8EFMgtrgDGalHBOiScWSyeaS9mXSLfAfNvwVWIEhxzU1YRpIA/lRprx3H3F2F
3bDYLOu+JXKsGSst3fbKz3kCbMwMKWYjfmAfl3ZyHsaNeVqxp68xHDeXPSAcmXkv
DivgDwGPz+SEWRc38Vfrs3mu3xoAv6moxmXyQ34qXJY3lodPHbQIWcyTg7dgYGzJ
8L2AkhO2gEYrz2hLsgRdwgyPsVfqcMnR0nmDbwqHN4EF4Z/KQD51qHagINCh0RVp
EbqeZBMHaXDK2Usp65QYS67bAIeY5QiNxXO+f2TovNUjFtzJMvt/n35eLGdsB1ns
lUivXtEAvoSRuVHLMyx175xiYJ+gB3TpVDb4oPSpmjvcW49PsbbTi/GoazRIocKX
7vFCxXYo4ZLZHSbrSb5o6/MfVzKFjwcggCwFur05kpIO+u4iCaYiLhhfY+tzyNzC
70uGoJ/9EeA06+FlVYD6/6xrGK0gUVSUI4FuwEciPpjJuAB0xRzDbphO436VOn7Z
qA2ZUVRMym/EkvAVzLYdcgPT/vP+8jqgWxjeyzuI4kC7j9B4Prd6REPK0T+k7QWT
OCZFWx23DZAnMiijiOIEFNbIpaos+cvNZSqbc7gWoMS3MBc0jmM3EWRZkeWs4og4
N91gWidDH0PIcK8nHNf6v5OftRDNhKnZEvVff7h8SvxMvBZ+0YLjAm1SORTHt5Xv
twolT2dwSAE/Da5lD/QeAbIkYqUlX7JTHtEWg+k/MMxvnWns4UlE5LecewQGvhh/
AEebQpl3xS8F740CaTXidBnwzZh8ZHwniR9fjPngfJY3eCNaYsfpr3K+9kLt8smA
qzmI8ubr6knRlxtrC5X0GN2pzHi8vUzHmFzVu0Us/5Va+z4/c9xklX8vyPnAAJMr
fpcIHAZA6za4NZwITZ3c3ZYBefO5f0CgMvvu7qL+vexA4wUvXuj/TeS7Ho4GdVKn
vMftjwEhPkm1dCQXZTs6uw8HfJeYwXr+mO4Anjq26G+SOpIqFUDDXaEqbN0bfcBt
K6SLC7C/RKsfv1N5N8sHZVyifwTQUBTdBGWQQMgmKN+JH42xZA8oJmsIIN09BZRm
7pFLrlTxamfPNhwrIWMGL6qVLKQPiGui1K3B9n/ZxK/kffA8DrceY9lRFjNOfrRu
AD2z5zzSxiJK3qkfOBvVXIKSLtwaFEbtzBUh420FjBVhOg6wGg4E0Bid9fvt1bUf
dzEAnMLl2AIry/dybN0xDl9MIQkeON8aJEjmiYU969e9Vj0r1S9WCgae3GT7a46k
m1CVp7tvV8uc/+P3RnsEDrSxihNjYp3FkYTXis2i0zS0Zm7UuQA65TFZAdx1W+K7
+JAbGEHL/mr8s5NBcXGlJcNlXkUZb+8Q2NSk58uqgzbFWaMHHy7hhZqmpOQ+qhWU
BFLZW9QtvHL146GxfH3+KigstmEfT8lp002z1+3GhilNDb8wk9BSaFKDChGvUEB5
AVFTJJKL7IjE+ZOMlAlBB4QJjCik1oZxHVDnpTapPiiSYMQKxc5nnsV2YRLAPnYo
b1ZctqYFByGGkq9UUn5FgxaMAkZGppJsDRxqWpezbseiZVZvGqE8j81Vx2eh5AuK
W4fcdYVFCOKcQ47XsZlhxl2RRYnKBARUzxszZSuIXIaSgWRiMVYZFn929cq/aBr3
Y5roYPHsMTXSD31p1CUMiHi0Xq1Ly0HoA+aONX8DLqZXgQwWquu1dgZt2X+nXbvw
7FDQte0OcOdwqyMudvDgVGDIddWa984Q/VKzajxgczXX9NHwLmj44Otdyihg2t1p
5ERVbZFlv3zbBIukZ0xWBwCWEAEQ7NxiOWLrKYQibrMHfnVmPRQ40rmMDyQxcx8m
wOe7t9cIujQh70HHTmmgnexOKoSl+HgR2NwJ/igFM1lruccIRNre7mNT3f29xwDe
vcekIIgC37p0cSBqoOFXIz5gU1WGnoR8s9swee6r8pIIU/NYF8K7zfOzGT8toMOv
0hNQNZmR4YAZzjltEJC4ESx9ZlWwW/9F+3dvjKb9RaCnXci7w9MyrifbR40FtLR7
gjGbtH3mO7x2o3/KTAVHKQU2SAv5Vgbw5ziNPebeDkzsoHSj3N5rD0/e8HMQHXMt
3O2L6jx8FuyOXdnvZ8l8rsAneH+H1S/p/P6+vs6/tR5LJuX+DXM4MKSiqx1UMaTx
gpD47l890Xh7SpdwsM5/fbJFjt1uc1Xtu/V+j1BlyEVZjkfk4MnnSwW6znNcMaiH
R+kk8aB/tnQBdZoogllHIWF2gECJKpWhL5LJ6tyUownoPJKLaYbx4stbr1Wovj+8
A9GIZ+xuzPAMkdvNXom4f49CCEXBH/cU+h0b8zD1vnP9L7Vqf5O2TQejGU3bhRwG
ItJIgucM7MjmG78PE+9tKFw1mxgblQzFxaNBrEluRf8l527RItXOJSs3EEVWrob2
sgfj4YhQg9CbGYaIU7oxu/T1GT/jchCPHlbK2daRvhVSBFxLEG72Hde5BkE51ni2
iKmXQe0Xlp67RqqV/FdSH2YGXlpCfq8O389Hs61rxQUAFWDt5JVL2NikNtoAEFvt
siXCww1KWslXZeXxLTnfaOSWUL8Fhd2KYyDZqQ4LLqF2guHZ5OLinEgduSWj+AaZ
yuu/DvtV8szgANE2bVNHplXIK9QRHolIEwqvtH9LLh3H8KLZ4S6Cqrv+3zgZp+cG
jXdIFH1OvUyhBbVk3jneK51FvGVKPT4z5eQII+PHsBdie/nC932DwXdbHsRYqM30
GyNbdxYZfK5/+1x/I+kYjuOJLkfZECkBPAwL6ThDZ9VlCocv47oTHb/Ve6psP5gZ
L2vHk3jrzBmSwqQ1Gprc8jDcWIVt52Exv/auxZrEPFEqzabowRieCMq+L3oYq5Nr
MoFBjdx3yv+/CBcCBJmZ/xHVWA0zMbhJp++RRfKQjvIOqOfWhbnDOmAkM1Y8CAqa
4iVFw+9g/v53qovBYT1jgGxQ5tgDUBnjn8o0/eY3+uqwDjRH6rPorxOvG95hyLVd
QTtpXnml1OxmmY7gdtM68QA0WUDy7QZs4pvSHSPoCLa5vm5JbeUPLrjQKknG5wBn
KbfGNb1uimSUAwvQ0lnUvzcXCD+FXP8Vl7/V4PYtlwDTGrFrFGMY0JQIVllXj22R
CWIoYRTDHn3T0kby4XuXEeNKrdRxeOa72NjfG1fZ8Txu+CB5QSOCJfgiBmmabuec
Rvm+zBt0sfEXA3fnQvS6yG37YqgOehy+NcujEB2CklNDvoX1CUzuetvc50EuUu9t
gmr5BpoFfLE6ZtaARpdrfptXX2L+Xz9N3YfwP8l0x56zqEUr82X51fJcgcmWQybU
5cB9R+B/8NjqEX11ON0W+XfU8JIitMiTkJSDxtF2KWVGhVYsvqkLUv+HBxIV/3tq
8RaBx3yHwwN+csyejgprc7amRBRH1xw3jUTCxH+w2q0LUzvdbjBEcM76ujDVW/kq
DVbGC8kKMUk78v59MOnE9lRMM/e20zt18JPrGtaK2oztpSLedS/cDOUhZaIY8eNu
eeAa/UB1L8TQERrv3J8OkZTkeZ4C+iKPMk+1l1qTN0NVA7C6n3xjJVwdvdkzovUq
MUOYP77b9lqRtRhMcu375EAbjPWBHcruZK8nApWap4OEsGqL4JZLA+72kWReJyqV
7jG99N4csYWb9IZDcxgDwW1RgIQUQaEFmApkNrWdTl22v5gzzYvlU7jBoclqegPR
SmxdVnnZesEgr2xQs0Y91V+xOwGunOhT/Tl5JnxChtVAq5rsUd++lWVPqWUY6xs2
XItJVDj3tys7S6gYnx9gRgjLL0y0e11+5O4TTyCLnNpLaD2e48wHXpSFdjmYQuXD
Rn9dirDYcwe+T7g9/hy1aFP0MHvXagguz4ZJDMcqtprNKJNDYbMqADOB7K2VMO+6
bmh07f3Xd6Zz0WiZoAPV+dCLrF8yKNafoAwNL0TzrJqTWvI5wEJEOFjMjRxVySRa
sUgTXfc6gKKJKBGapIBXXC3rdNOMeuBZfyaleKG3sgQtaTwhYNmACtlOCVUkK17s
FNxsSw/Gp8FMpcfiOBghRdp1voS9xilHY6KcFuu8bRBXM8iLePBtFlluoXaV3j4U
GK4AD0Iin3Xfexo2r8JsSvcwpCt+cglwpVLjJBi5NWM/wzl+l//iP44cL7UqUiMp
F2SO7lhaiuT1o+4Yr8x4ycaYiUYeezCiMZ/UUZ4870CwWZ1ZB21nVvD9mH8wg952
bhOWkUXWt530DSS2XWW9GXqArx1FD4yi/7bCwHO+YKwPCLZL5DK35zrITYkIn+TO
oWH3Wp7luBv5Zsf/uo6SG55mhwQ6YFKw+buqt8yk7MeYuq8lT9SDJv2+LQgX+tV0
W6mq35faSuWCfgprRt9DJBq53E5ZyNI3NhhgYrePy9YL4TaSzemze1XPZCyKNFdy
IEd6Z37QYpmLXCJ9Pd/Uy9NcmcESBjuVrrgbqgMHKcpQFalBasn82THtDJgRIsVN
tBr1ZXzwYrQqKsecJ/IRnBPjdU39lJvK3xw9VQ5/kZbGOWZkMtnk5n7oTgdzo43p
RZC1y4mjaXF1u36c5K3jXZZ3T8DS5VOl1VVmW2MN7s0lOJSpoghquh81R+uzo0tk
991KtD1STMG/LPPXcfi+I0x06/w6WSqjktv9okc/izgpSWAFj80le/UhHH71zzol
az2IXqv9E6f0UkDUptXizO7e6L0x+46EBLs6kzMCd6GW+RBUNykLTnxBRYiLTogp
6k4x+hQjhh/fmhBZ3yo73Q8WkbgNx3/fWoEEsBBn8APymMa55TMcInd2BYNLs6ZJ
Pq5yGwX1RNVIdadLbJau1NIsi9LIQVgI49VAjzxv4J/CSCqxCemJTaIYHGmNckah
Z+DqUXTH9zeX56P/PqBwo0mDD7BmuWAfOBniJVQjAy9XKql24nhGGR14Dix+5qYt
HFDPjMSqmOI2TDIES9XklOQea151rdRsuedZ933PXZXzSIR88y0aD2bPCAAHCDFf
ixFJ+tBdqlYbIpphi7ZtZvJbRaB15pizkwhIFHsLsxjmgn9wJZ9LxnwRha7dHNKg
nRxVp6tvjEFHqOyP00i7FxwG0uVZlz5VvZhb05bsiORlglVVj03Wg4ESIiZP1buN
LV1TnWMdboeFeSovIl+RYad/aoFakXAY0GSYj97rROwVPZRj4an4vPSEcEiWmPE+
QFYnkAXwiLzy3LeHu1sdo/2UOqmHfq8bg+4Y4atH/PF8fQZUeYC9f3n2PBCc8oBj
Yt8iNpm/mnJj+HycyBwOvAtVjygJA1D5pEPDuFt30lpt6X+7xj8IaH9UnUTnE/Y2
c/6NWSF/UC4fFvhNeo1D9UYTmNuQP7S0nlar3rCRB/isd83z+XqZ1+TJq4DKLNSP
dkh/ceR9uB+CbPMbOPVuvZAPSo3jF/zE4l9Br1s613FHvn+RxhfZ1ZgNCWA8OhDG
WS5XPoxxoIdiX3y/bS61JdwEg8e1Z7UblsE1ePrCxjBKGKGhFRU3nqGYHY8aIbre
Dcv3V7xOUgxeIMQjej6MjItAELzBghVR9zawQA+5KBUaIXQjUI+k/tgAGSnBkpAC
3Zskmtqlhbish0VFgvODzbkAc2NlfYo6xKwvuFHuMTRZauGkx1F5nWbwrwzqX04U
cHnqvy0kzBeyhjXBS9Dlya5CSNfJvN2eBMF3PLmniEmrly6q0qkbAZGansmUcCNZ
+PHVJAAcXBcNWgyx3Ya5pf8Oi9Cr7MGkjFgV7koiap29Rf+AcmKgRXC84ZAW0Z6F
1nWqq1s9VFrQ3fBPR4TcYEQgHjQbs4toZcYvzB/gJ+fk8ER19jt8t6HnT3uLdNHb
NoL1uoH47C8avdqSg47pJUExXanq4VpPxdp5mEtz1WsUgYqc4pHv6mjVNqHJUPSd
2PI2lZvkr8GaaElac/pxyd26dCzImrsvRrEUjTS6Gu56nobYUmh0bbePykh7K6DW
DC9kQAUiff44jyOcES2+CmkKm8jmujutyaVMBEx1mOKbGa0Ks1n6nCUYa1i5kLnQ
Ec92Pk9rvEKZgSRxvb1q74jHxQ3BhRIhqq1gU0WOMfMHdku6VOpkFJhAbXLUPP6q
MR9efNoUG2uqYUFNnlY5s5jrgo6ZGZrSkO3ZgQJ9NbbwUmpK8lIaxQcJKzNxDgFK
F9GWHjiEylNnFzgtcXIeVERmDgajcHG4D9m7dCShkaEQI6lWOSk3Y91XGXBL1Zjn
yqgo3vBTETKK5AkMH/iI5XfyicSC36pwN+JPiebcvZPBn8iTsQRO/8AdoKPkbGNP
BjMiZGYS5FHuyzYSWHMs3EkWa56blH8qPh/RIZNJhjDFko++D6T8Aqwq5I04CcbC
BUgyua+eRPfo8C35r5jZ1OsKaoyoHKL4HsEoaFADQt3IjhSqKueKotWuTWHnC0LM
tgrrEHdfRYfZ/fr0cZY7E/gMiTza+UV+gTG1HFk8j6ZBC7OjV2+QM9BGEb6B1RBc
IpcBURd4eUj98vS0RascboSmVAHs4UMelxohMex1SY6ePnXRR1+f3BeoDQqeRB6G
3YZAQdUgfOe8zW2opuSgFjZ5Te67ktZB0ljC9lvTMwvgcI22rwoGYScs8jBr7HBs
IPLzc5GKKPYUNbBqQqs+c7Qq6fjctIq+JDN1BEzTBF+uQi2kfLog40A3/DAsg45k
/T++Kd4jBO+WW/In4zKLIai087ydhodaVsPuGP7u1KRKSoE9mc9qdEUB+HBFrrdh
+ws7MybCTjMUWLflx/818Mi+hx1NwVszPa4mgSglxhuSR2PQmew5OwueEXM9er+5
PUyBPJlCYWDuDWxg0RLxpcURFpnr/SBvFTAC7/sTRmb23oaoNoO2JclLbfBaiv+E
F9mT9jhlG47f3oBdQMv28cAu7hNRDs8T+25Ydf+eFsAfScMDM3QGLVdjahXBjxok
L9q2O+SniHsgczayMzQWYSFpIgTqVBIYDdf8SrO2TABdyuPrDd53JC/YCcRd7U8o
eBD2x7xkCrRk8Tm8lqaYQRB1ePUlZ/0pfrXZ7F4Hk8VHkuMdDdUaVxlp+SBXeJXl
SsyPQYJVZOW5iR5ynXQsAR/LyOhgCiY7JSArZGpM89FV2pgfYFnqm5UbToVhWPuH
nPJmo24HadaE4PVRTSBHIecCe+DgWHb6BkweUwVme8oljMKudfmEE1xVSggJLq42
0457U09OpVcQLWIB21FRi9bgBeF7Jd//LAiYu5w7KnZzZ0bRRyeQUkZUVmFhBLVE
k81SeKEc0PfGL5/VT6mmv62bSXeTeWV5R0qZRjJolhFoLoF8CivosCCwnSVcD/Sc
RKGHfLCxwcVK7KY6oQiGRrR0uYhZY5qp3qapIXdsAyDqhEno8ofUHrvr0yUAoq8T
7Gu+yEHPqpudmzdR10a2Yv6nqpybTpEEpk/ldrfjHjDwr4SCJVH4KA+YYFGcl9+G
C/R2rNF9oF+9KK83lv7lK2EIeA/mJ7uRrd914N39VNvO2tYb/Rb4adbvrQ/kiqDT
HFfQnLooNFoaS/1mqbaGbcA6+W/vIz1aHQ7DRQJruol/YaLW+2UjWCreK0ZcxKHJ
wPMzCa8xaGfJ9RSi/L/fABWDUK5xBf+8sK0WsgtQ/4r6uN796NoZYItpB+dJv5nU
LIWbHuJAOhH3M4dGYqa0zS2UTcbsinuBieHbgeZ0kkZzIDjPHWv2FXXYwO6fq9QZ
Ba021d+KfXfeyvDuMzeHOZRyGqrCYmh4eZmsuuOvbQ1HtbHhLP1vGW9f18ks6w1o
2WlS/5sqaxVyV6yhMtIsvRfh3Q/cALnkCJTjjCwW/BfZ+khTBjy4xSYIVOdKu8ZO
hx1Z4eyVthS7fNyXwy8yuMiT3znE/MSBnx7N2F0ggRysuNSMGMC1aqkwgGZxwXOw
W5Ma5kmHnDbxPp7BJKdBCiboIvaojA7WMF0ZEZLrUY7WihhNluJ/C8qOFmQ4ik2p
p1kIbJU3LdIJH9l6GmBeL60f3WhBLFzvIDJjUQIluvy5qwirGcP7OnDGuhmRKWdp
bI1hHhgN7afj1l3Ued3FNNmxDbWr+m86cni728U9of9FZ+RACDbxb98+S9r3tzmK
l5LXRIpp85tUszhv5CB0z+IHiQR1V2x3o66oR6sFst949jqTs59+4HwWRkJ6Me9a
533r6vOEIClIvJ2MdVio0UPq3pbSQiMBf8ZmD9Kf/SmWDq/WeDNf5qKgLOikQn9U
cvdyUjPaB6IUNV01V868O9nwbqWYH02Z8MKhZIg0+zuaZJWHKUM887wUT+b5dAtv
xiXD8LiUWrOQEiq71axXwQLf5nz5ml9KQ9lmCpsaFvJ4ffUezT7v/VG5XZfngV1R
Q6+xqZQJxv5+Vislq48jSx6feyzbSNMaCHP4rCU+5cIj9mxKoWv5eNq2K6VOuPD6
PJ/CdTGDfOZ7S6kM6MXEPkZB/iAkP42iJlllvGtZmFa6kox8RiRaLTbw7lYX4pWo
WFFkbkYaQ3LV5XHplmv+PrwQyrF240dWaqKcQ++Xzg65RqrKV9tyMYRtUMB8NN47
1veKCYcmX/RwQJLPfmL9dm6YJ5Uz+6F+AFfuR2buFfMoMT6FeA+3a4S2JR/++YHz
1sO9nhV6nwIQ+0DgdNjoy1Jb1WzDq/G7aLqhPN3TGzmdVUAMLWlZWfxpWGnnjX0R
O7pQZI+YkDyX3MrlrfjfqKrqS6RgsxNJBxAe8/MlySo98Gos1i6KM41k3nSFXGx4
jHkFPOM+PlsnLWu0nNMAtB1O7C79yBDbbengtrbqMsLLYcl8wbjqAX+eaq6FCl2T
Vsj9gF4e+9A8/xSCjJaTr+tcq8Dv86gFMXKSgs3WJWVk4HbFvz+7VIu7I3C7HTdL
fLvtyxVuH+r1TYFmEX53ql2Pjl2FFxEa3RoguxCoIWpAiX0pL3rrTDZCQwZcZLUr
UsAcjJGYZXAuS5sLgy/qDu+tXRbKcg3Fk9W51g3dvlJ/mEW+lFhS6GiSGBQT+jqc
oC3qdyyfdzpOSu3UsoC8Z0anroWPRe8drxCGpifYG4qFZiNGkXdcY8qQ2/ZDqwph
sFsmcwp1+wgyFr/J3eFWxvAmPbyJ0vUINymAUdzK4h3JKU/UQJvnasRxrmm6F9F1
yFMGzG/wGcCk0Cfytpga2z3zR1RthpemoT70wGQaI2cTla7F4T/cK2xiHG6fck4h
/7vGcBEZuqa8eCYg6MWmtHABUPRAVz2+jrTPteF3h6Tw42K4NWtVrGq+FOsI37Ey
d5veWDssq0VWxhLl3oUsTtnw5o6I5YWF6nM778QlZUA372h/rAi6YIjUumsa8BaK
mpbdqHhDQvsCVgaiZsXsE8SklDfnyAcPlkfSVMnoEfEU6o+Z3RA6OPjWbs2cMr3c
z8oNNpwBljgPUHpcGJnwEFSA07JIbpaSTluQSAsMdxAJo7tFRTQxcvmrNuWFx0n8
tMvvO8kUTBC4CPgUiT8S3Rm4ForQUKG1yhDtasIQvRkUd7ekLE6DjHxkQvvBPADO
fUANJPZVOV/aSS2vmCWC1Jxl/cIxVw4M+yQvtricOPkTQ8SV7TuGHnX/9Ao0tgyW
jgTUeTPox2H/h/zQ4LEvbSu/jus4iMvQcXp8cdnmgVb0pof0nCv7HlZJXkvX4idP
RVvxw4L27XFH4EDlt3FbYERT7WEIzXT4GwjDTcScD21ehhIztJn47I314zjFwVAz
HkoIF4iajtcMBTySumOPX574NUkWW4sTwm8/1UBocdA2uGQC4L2ZXC8X3qTwHUes
hOXZ00vf+3HmyLnNKpfbYF+nrfVw9kgiY456W+U0zG4mfA+0fM2eVXT3IVuslgkN
q4jb1qNXAaZwKExAbkHTSaaQNcqz1C7phXnXmc5ud5R4AN9b27prlHaPxrcVhIwk
Vu3AYP8txM++2edOYPAmvSK3r7fUEv6im5/qhRUC6TQWx1SIvZXlIAQFd9EJggTJ
YpnFoMv7XMvm4mb79W1xzk6Cg7u5ZcfAIniKy5MazPoOuvLbsXejki9ehnP/ixMQ
iKxL3AwZnXnp+O4RivUWj7XTZHU3GDObeQ0kq9pe/vmcXsVf15dwe/H9Lxudx9i4
2tmrapo2/0G+L/rmvVF+ktIiGAJhKzVmD/0rT0Ifrt51iPnkFoabLI7JWM90OsOs
3qlSJ7w3etZR52o67GAQlhetFwmBEb6dBgGIoEkkH1NjFVdp+IKVHODlpqIus6Bg
/4Nej0KMHNnagp4tJgYtjzD46/EEfIFhyVXDJqW4s7O2RwOilImcdUYDB97P7Ree
JSFKy1jHFqzmJHp5tfz4EhrCfJcut8cCk2lbIdBh7I6K/1sJ1wes1N7u1pIgxAWJ
QwWvqZseUZbZNdPcdDoe/bbC0geqoUaSpRdMXaPCUYem/2luOi1zt5p18xqTp4Wd
Ptv55u98vIOP75tUEhRwqGx3bhYDyG/T/fEr1YDY5rg5R1fikNjRyatIxQJv8gQj
UQTw6lFYMsFoqPkk5oMkSZvtarcGjvzTWUNfPdP4Nozqo9ckBmv5xjo5aZdqyY4H
Nivj15wK9r+LPSKSlj9Om2mpIdeOH0Z15RBvTiWUI1WMZ8g+1ULuB/9Hw4BCna/X
NCgxI0nxDb25yeKzhc8bqoJQyVF4LGKCoEV//tFws6cFMzb1YgBAQevDI8+QzsCe
Vo6aQxO3J89rNIJRPSCqLVxEdwFsg7jcJFvlXZSDJpXjTh0hvnYJyIYmTbJc40H4
OUlIeZBkL4F/ZB930Ytc//P9lY8Zrr52IgfkaOzaJvjfRzsHc7fklVNhQW2kDxJq
ntGc/WwvJmyILOPauW6oOByXwvxGHEyyK8Vx02jEzLC0WopiZgfqs+YOxAqB7jzW
LkGeMAn1sUDQmPYF5l+ygp/40V4H8YXlt9PQB7ymlYa3lKsZnWfu6eAkVVi6v3wW
3pskJRKeY2tblQ/Vf/uLyh4YMqYEX0qpM2QYV4dG87NSLL8s5J0SHw0GCTY+ukID
+PIDDURH70qdH08ERS8Hn8T+ijfxLvRJCbrTUT04tjulF44x3L9Ih+uUrMLcUfzW
azDqjXpLSxV5JVySwPZFF0EHcsfTb5Qt7UVmI2av4ZjEjJkQySxC6U72MAk1AOb2
ZsTcZFnKXza9MD4aWidF21pkIX+HGEGYBLbVCh1cLf0tv9VeheT7o72J10gORsyJ
LxC1vp0fqcK1Pe5fP38qmEM2UT1WjSjQdF4UujFZpaTkQhufqMJxPAyY+NmAD4ud
cSFPmaNXT9raMWFdXKC3x4pUHPFl640YrPPxpc7HBKvFS5yldb8AdiHwEPSuiqiD
Wo3Ee/0c1d5ZNb8Oc4f+/D0BhgSoA66Yp9pr1MTVXCQw/FEwTsH4LnTp5UzDVoP+
gWPw7DIVOf2jeUDFbyqULixsVRyG9NbYXFdbJ3mvjQjByJWaGTkWO3uuXKaVQt4G
qUSGX1d85C+wjlo80QvlYnLov8A8ARq5sa04jb3FJsjzmaEtfGN1+GD/Ch5KuUB+
H68+Ltp9gfF2mfbbGmoosIJvBOh6uDEOdylAov2tIGWNlytdxbgOH4LEssugg9Zv
+FQ1hEl6XdnsYu34WEYTL2dL/BQJyPA8J/Mb1p2nUcxm2+tRpjhi3RVq/l+3KP2M
/2vGIBO2TUhsd596JpbjVLn/Ukgb23lpaec/L636Tx5bA8cSKluKgP+7DBx78CHE
zA7/ogjN8HrAYwCNaYMmuj6IfybXNknjQE0YoivG+bTN/JRxl38YE6DfIrLpicST
XDDbOrFaCNlMsbAMdbu4XNBd3hM4mRrMEU6bzBfUyR61SZfDr4yaJzWKYj/8Fnmq
z2hp6D6lJeRRkuZBTOKky2A+xeN42mHyx6Ct8g+Kn3Pl/k4jhJN2kvGeiIJkHRv5
cUXW+fglzoy+qmTHjgxN3ep1DYNuu1Hb9GNUGdLl4aqm8SYN+yHsFFBHNrLBU903
zxq160xjZILy4dH3EWiHVrFZX80GVuknaOezpo4RYUvu88yxhUP7N1lSAvpRsQ00
JOUK2fnufd33K4/kJs5HBkhdVGHZRM2bD75YiSBMLx73mtkQPBLvDSoFFOuf2Psi
b225qVoEqVSfteIgwTRAeR+Ozo8lz25up02aWf6lWJMjtQDi9BNF4Igh1IYFy4HA
Y0/CIjzIuLMeLarrxt4HQHQqkLqWpak2MSi7jf5YKBwXCFfuje3FwhVPEKsorjdj
lwNYiuZ0rc4Wzy2kUdSgzu0E1NgJkJ9iJN1xm4xRoXN1TtdiXwUKSR5OGTDgp+Pz
x4Caz74+vIXYqTTbxTakFB37sgs2IIVB+ri1GgF5Zxs6SU1BOMrgL6TYXtdV2vYU
zS8LFJzLi5fx5cS8i5ylBBEcXuhH7AXcDEfveQKcJ8gADkToYcf1ukS0125bV/sH
9W2sG+wPkplJnT86ZimKvjeIUdW+MrJ3ynmO05eyzc/9EvgHw3U4K+nIdCKUGbs6
+ezvO4mScErrxQp3cx+D7nqqCEt/anVKmw5dIH434jDkMBdRhlckamUmX+in1aWN
8bV6FQM1OGrOGuDYFPoxOG+gaHWdBmD7oQGX2SCli/qptuRUsxxqXS0mNQ/Q/7OQ
2wT6En0yHWprYYH2P3jFChRhHrqs/uMRIVIZz5ZV5hLwk4QZFZ7ltoMAbq/XpzqE
+FW/ZWgKFg60UJTbPOPVfhsSCVF0DI+4slg/dC20CCYUUy1mGOHyQxqiLXzxK/K1
Ur3Vy0gLMOjWKI7kPTp0xRHvzlpCZJgKERk2KOKVQZXpc26S9DmVM679hGwMlbwv
kdUjUOMDAgw9r1349snwK+MIlrXDJV/VvLd+ox9sERpZb2OjGMsQ0oMdh7K2PZe2
51Hq6XXIXQnlEHoqdOH5gDKCe3AMS70lBJxKsxzqZBujyxeQRgKFKfJZrLzVMlxv
Q4YnkHJEJU7mkFFoqAy1bvF0se/zyo3kLk2yY0MuN61AQpeA18xJ+jiPXCJov7SA
QfxiWVYsdnP/ZiU/SAWfF6MTPk8mEpNAd9jEFAP8bAy+JRXw03jZseYNcfz0YsjA
GO3ZVeBAgEVw3Eagl1ELOfYrTyIW4Kd3K8Ba0VF8gVpFTTzgzGfFOWljvC/mGCwC
8I/Z2zqV4IT2G2rAc+m81CyDyPAYuK9n/s/S9UeUHvhp/ziz/WifErFrSf74VAW9
yH89HiQXlqLu+JVDr2qGHpL8c5LSYqNMttevvXlgnEni63QRrzvzQ6olj54v30k8
ET1NUScutqCbpscXNEGcOFxtEJU+zDSIJNhQu6BXuwbZJlpdT7GqYMMRofZWwRDx
QihaXbX2Bc0TmU+rmHzn+XTbOSOUtoOCLmcjCb/77GmjxSc6A8vO72oNqcNjQD8n
aW9SbVOS8SvLKtpTGMV0hX6zyHlZmvDD9j2W52NibEjDn4vMD/VwiphgFLKZici2
CV6zYWWY3iXTIAy59LqghxmQNs1afIL4QT6hpUFHQaJgrgKlvW3y/gau6+NkZ40x
HY8OXVE7mb/kow2+UKwMECm+AcXsiQUaPfq6Hb1HA2BMHSK8njSEQn4wqeypXzD1
GpHDBwSkNgwCUkcDpW32xqyN80rrR0jt9GNjlcIIEnwiK1C1je8wmMcQMhKTJFZu
ZgGCUw+ZwFDzOf7dtSgOAluETjpuR5t0a1kLeBRb6yYNShXxDj/JA03WEoX3U06m
StL2vgqXixM9GYBBaJk+OmtHN0bD7m4o/Vc1mLfFTMXxl9mrdv5WpaaCwiiyBzjz
IzqROymAmwZpZ7jcl7G2D4nNFK022x6qTzB7ta9W1i9QoXXrcnRlU65V4BStvQOt
mhXw2vL1sdS/ShcfzMWRWV2oju/ysdmBcCXwVytMJb2jGgL/T55RhCHvhd6heRXE
Sp9McpRpbvsrrClwjQtUowT4fUwlcz96dxd+NfOTSesYSMnKfhuQlDnYZx+pwGB9
OaI8Ju1JLcSCVYvgfxJ5mmC1FH90w2zvYn31kBSgunu6Z7ler0LZQn2/NAXUefd3
UV3Szdba2dK6Ydy4erNXkABdW1YiaOkaHrNAiLdKAdHmskq6PKb95HbJIAuRh3GA
xh7lVblwEcNQeuyWkCAnRktT5e9uLrQ+vzyFArsJInVLJlny40Y0+1N5H+5LzpqJ
msIlTlhBGWYC8pMApQuVkyRnb2aIgOe5ENPeaxmnns+lZ858Qwd63ZCfUQVrlZ/F
CD7rmY/Yz8X5z4egMyuVKGm4e3uNaJOouWlo00QP0f9+ua0TxdJJIPs103NSVdxP
l1c5VDcamYW99tDexikC/+syeXsDA/k4SkDbUYbo5z4fg1c0LKqdYrgKPeP/VwlK
7+Ibxx3V8+F9i7L0CVUm/sZqgIYjxSquMiEVzDhSfomSX87SLDTMW4PZUa9H4IC9
hCVm8tirFGeBeWiM55kDzAgzswB8RR3tsTMYM2QAVRTOLtNoCGD5hgoc9lRElkP0
LIsKTtYcVbiJqtvr8uZ707qXQLMrEDDsehodvEkEHHxaXdxq8mexCFii63E65j37
FaVOsvn7xKnrIhOcJ9Ytrpu2zrwQ6pskBs/RFHBEAJbQoOFiiKr8pjvqiDG3KvkM
5lPFcgngsTQPQFEHvDse5YsfWOwt4iNOhMtVuEEzoTJF6xv1EFCwctgoEasrnD5o
yOU7Em7kEmEy412n2xH4Pn8Tr+Dcdr6V7g20tgf2/8Qre4F5ihuOsoSWzzm0USZF
DXGgCxuMjiRAaHOEucG0owN5r3WS+dH5B65OhnpUzncOGqJBgL23GXeSk7XQUu8t
nMB/c2+CuyYD/8N2Yz7sBH3KKezwls6N2BQ5mY/uoe5lM8Bg3XThl/KzGdfU56zY
120Jr/haSVPmDaIXRhe2LBrBStHrzPStBVrhX/Hhsiq3lXawRq2qYYNXUvO7bOWL
LUn3rzOAhW+dAyzk9dN9kfaRpkYHzp3BFWqW4Yqqmppz1iNJF+UF/4LQnBsm+CVp
n9AZIpnH+axhponMfcnH0S2FAEXIuqXvZAgAZOiaE/VAl5okZ8+f5OKmlq5j9x1I
dwOc1K9sE44Sio2sh9Vap0lNpQ/a6n/fsf6enJOvF4N2ff7qwetcamVvZ6qE5WzH
U3z8ftBQaoCFru0rBHiQkM3MLJAJfQh3+zJsWiwEMxEqmQ/oBaMRJ8lDPJhBW+J7
H1om0ie26qYXMt0/+O/dBmNm6nLG8LlEIiMhMptDS9a0fpKM1/QqW+4szPMd/JDN
05O6jcS9T5lGL8W4ywQIM4Qlswub90sZ9zTCkWOLWX0f7TrtxWhdMJQ1BKgDfYH6
efVgYTzz+Y9fSyg7LZDKNAeuT6gjr066cZfIemu+NU7mpkA46FsYRCg4CC+znQrk
HH53YVx655ZOPNcWNAji2VXNuG2QbaZ5r6AnKsDr8+QeLKGeKscRVS3xcmk4QjZH
h/3bOUcun/JIk5qVpb8hSGadMl0PfnwhfvTPFZLu3fb2vuud4gMiTjLP2RELY0pE
1ZqiRaVaidK8uqgu4wkSJyulT7MZmXxZdVn3EpLjne9P57845vFyZyReGKPsxxAd
kjdy/X+6NswjBV9jkK/QlQglQgcfcN6GdBo/iHpJdCntj8ZiPz/8fLeWd7oBmcpG
jzyOE7D9JKaGS29Z+HIWFvNgHldtktfdSHiUY/WXTzFEfRtcoL5c65Y8SN9l/eBE
4S5DeVgQBTKxw/9kGNTr7Ct/tkwPa8vzDkHcICfNX2nlMtdBnI1qduC+cEJIFLLU
krF0uTMBNZCRMhdIRbL32NMExzJMLtXOjn4rdlVmWak/HCXNRF0vP2CzgpakHJoJ
OgJq5bJ+bygI+V39MbU1F6B9d1RgtprJE0EqdLNqfHsnZhzK/IZvkXd+g0iqUNRc
XVYGhKwlUCCFhKhLrvgifYrIwDuIYxqwISba6Cw5Psnua7x7GiUmB4Sk82+ZdIo/
o8HwcUrJDowFpdnllWue2eA4i4nMPnk4D75Og2+NKr1pzvPI2RBYzCRiO03dObap
lpQt28QsxhIBCJ+isik5zo+WJPkR4Hu1SuZeVzFDfUgJaezm13ajYPCe5FkdSWUv
R4dJBFeFwLOhDtwXQ0zOTD4gzvDed7JzrUuHVJ+fY7iiUBfcoCQo1rnG0LwMDYKu
DI/VvqaJPnKQaMXUfR1/P01jjsAUh0BU0UNibo8dSw/J4mWD9BylabtFCCfSy4lm
IPylbj5r3s3t3B+p+HWPQmqooGGmaGDxp8ShgBSAAWKCWLIbZS6aA8BlFvFHSKuU
hVP6zf/yWjPIKrkp3zo2hLmOi8d7EbQbI/Fw4NcxOH0C748m+GyYGDoW03DucxVW
UyTTFlAQyI7fa2sprWqzohL4c2z5iSOCVwZLMITvD8Pk1vSg1iLQZbSlqw1jH1kH
CiWv/ekKakBHA2SXTcdffGVq1RqZR5R2eoEIcrgWv2ejw5+juemGucwq90383CyK
Fp7+D8edBYRyJCGOr3k/XMg8hhOdQW4TweVTWJvR1MFF56jYduQ2mskO6LybV8Ne
T3mLGH8tBE7m/79GESjpqcs0/LovqWzwcYs4wzVSPPmEvguQoNOp0obvUQXw0orR
gqYdvcuj8UzJko1VN3mmz/uoOgogOBm8WBsYKrNMbszPiODhvpTmOPpm83uodHN8
N31xfneqAPsAmahbzrWBaQMLdRvQrTU5NjtvYYOEcf01HqekdQNGha9//TnuIB4C
OCYn4ACzk4XrlJUf2d2FZURvrpK8UFugFmVHePLcXrArzFU0RsdLa8eM6h9PM47n
4bDDjW0aZX9B95df9gDGLsKelF2pjlrCEUTgG49URBXweIanHHhYMP2jSTVCS4rc
N8mrbvY8Qh8XJg6DM5rn+cRakb4tDTLPyy1fYk0cJMuwfmNPDfkY2fwFnhlQ2Grn
mw76fOZXGJ6kc5ExsCvZfyyiJHdx3FQf2jjLZlb911MzL7vYSsNalhBZQb54hNT+
EnxGs+SYovntJpZXJ4tjNY2kZUU37x70lUtsOjyLvX0Vzd1r905PQt+YOLJcOZBG
crlVR2cuVHQqskyoBr80+a8ao7o0cXNwpgTzi29bHBbjOsrEDWeMkmyhCpNrzoLR
jdGV9nu2WSqVBD60lgkyprp3b7i7I/VI7vMOi69uTXqy7SPPYF3FZMYnJGfVmcpL
jqKlfKoNOYBCu0LeVKF8tWjH9Innm0G209XoigZGNgjyHggmdLh53yFMiKeMfwlb
AuV3tylzWrQC78u6x5tJlehtDoR0M5Jflgoih81R9yh0wyNUW6KmRbanNSGVuhIe
TaZzXMNZJQk+6QBWO6wUIwtSmNDRaD0OITqqaGPevPuvct5unCqPqvuzM7n5+fZU
NdSjaQlT9TsLp4yFbZyeI/M/J2Px6qvh7J6VIVrXC6Z53ho+qotgqOk5W5myHa1x
4xacQZSfy0oYhfxbDFHX08kcao6ISoqun1GgMoyjDpsYG576gs9bjZRmARKgzN0S
L7OFFJagkZA67n+fmtLkDIJ375TYNRrPeH2YlbgHJ8FSyI9FXxmiqHkctQPo46t5
MZ6nHXpZCjv4MZ7mLZW5lXNUFpaZGbe4ffyE/IZBKUM32ldjBTU2OV+3aMAiJLpq
vBeu3i6o2AuUnnI+qr67468Ye8f2wjwYaRg3Arta0OIjkI5NbB13/bI+k3VBua8J
Hbv0F/Oc9YERHMqO8Hyjus+SIb8/n0oQ8Ad8M6uCY1YzL5QV5NxBkJrtQCR3X5h2
YqrUfy2GOkrDSUr2GO3Y1GGMgHik9vsqi9Z9IpxDY9l9LRATBtR+xCnV7fm1TsAE
7WjCzAO7zK95AA6dexb2lK8+n23nugKHzpP8KSADNN8rTWteIBoBGJvoiZqP4BQz
9ufHUo+MHkHJ7ukJnbSDRJ+4bUUcf73UP2wd8HU0IFZkgE1zKFDjdNQyod8k2EV3
oL1UcMfVwC9pjhhmxJyhr2LjyGVhj7Ehcq8nAgI4tRMdmX0Vl6kH9CYVkI0tA9Tx
feBh2NAQyhHirwB6GPXPcSBIevE4aiUaLnTkB+lYkOVkuvLmQ3+J3hyMqe5T8tNJ
x8VgsZfNXak8iHa5jju+RMlltaMcCQEWnv23PWcdVPCVJMOFGaRgIyNeEBayqCTC
Z6Zqh0+uJ8xFYb3M1yTLd9JCExbwI/NBM8MtJTZxlPCu253/WmIdwD0ASSuUbnAM
3/AqQWRp/6bwaB18Wkp+ctSawAZajnO3GdleIBH7wNnmXyFIt+LkJQ8imGCHcUrf
sUvTF3E0R94bG4rlu1nLDiZKen8aaqaYawfNgkyvIEWEiqQYc19Nff9erPGChyoi
WsiDjBp7mdvsiS86G1uyiSDHbTrnQt2owyjPNw2dmPJLUUvPzs9F0waIvItS6HD6
wbP57dcAQsI7ZCgk0tHauSn6t2sS9uXicUAwvvM6rgOPQc3YQZk99Axl06rptDX2
HJLQjcAorqa+sBM6vUJr+jvQTrPBOPfl8fw9jxFBxzGbMkTMsePJsfy7BPkW9TFF
rW3NWNeqhQ9S/oVUMbsndjzFs68VXGvFswW/kvm9Hvp4aK7O9erQXYjSlSo1PeKY
d9jVjOWryEM2ugbOTtuNTN8OaQlmXWqTFlJiUC+jfFHAtyHSC9t2MX1TtcWmyFxA
gSSfgN1rIde85a0xYyrduOnoLqt8Par7Jlqr/h4YydqL7MyyANq91cqRvvBgClXk
gzi/h0W37S9GUb5463NW+zUn7nrgcW3IgYze1ERYCCh4pKtNCfzdFXxWqAqNzq9n
Im+LWK3cMGslRVpUZfa8CjF084ypmqQs9pyIIl0qC0kIr4Cn4IrbL46CNDWaistN
Tfbr2IVzpTYZD4I1dHlt3uC5k/6TnZNVIHsmHASci/GdNgznMeqtSE7/qDmfc+yW
nzXvMx49onSYd8NUXdiCFuulh2g4AMK0ka/7uJY7U0EigfAx4gpRFeMp7Qspwhf6
2vF66RD3DvyyWpI+nTBjfWT5058iW7iTBOqV85dRc2kXtOsB5mTWON5OagFyiVc+
o+duyXiGfA1S20ARTCmWsbPV5sNoYNcJIJ1f/ry3eLZmZJVsrPDIYCp550oswQir
rH+Qj+cwMa/DojeWIGXyE46/SQZ5c6qwoNcSDxS5OSZUT9l6nWtqZM1m8i19o46t
V5YdxLG4bO8kP4ktIZXGr79BY0IuPvYy3yQrUBuzuxGbxo1e8jOLTEChqL0Znpvi
fwDCFp/t50Wulu/CXVfnYEmboAXbKZ4v+0MTiUzGA5uVReOpviaHL/u3TY3Psyef
teQIVyY53czwPH7BbKfRLhiyl4A27txjjcvo//rJ4AihEvUihnB/xfC0WjrpjLA1
rs6Sz2SL2f4VBn8LFBRUmNf+IdPy18Bs6tZ/GOgkDinIn5zRkzRboWXhI72Rtg8m
Wk9PREjuQU+h4WBl1eHC1hiv+qr9+sf6aESy26A7u7qjKk5ggpT3dn3QdxMC2hSW
zEBtvIsrBcYSxlb+2TzhdCl0fMYY5xaTi0WcHE3s5vxSCH4MAv9Py7lF8dOaJ7Bk
WsP+c3DF58pZ/Z/9+Oqw9msVxGq7Fpfn57iAspp8zEaY9yblPUuBqEDmn6nAJx9o
bFmFY22nLoDaSwtTakidx5kufxro7F7nDqRAZneebzwxGvv8C7tkc0ebrf+09ojR
JGWUxpOOlhyHG/u4ZUF75k+Pl7Y4ytNxBRgGRiaB7SnEcyLEcwaCVlQrsrbw1qqR
K63YGjWVsSZDkz/iew8OjhCKAOnTN1ikGVKX0WZdTWf7T4yOr12DVqd8rznp0uC3
PLOy6aTNmzYf/RfeKOXaZtSBL+63c7x1gVK1FdePb4NcehhvB1+7yEsEB7v718/j
/MliPZspx5son8gBF/rC+RAaHC61T07pkyD4P5MfnUVBVoyAZCjokORXMFIP/nmp
3AhHP385cCeaYz3m7AaZ+CohURvmh6Mu6KA2fD4p60SxlYUJXK3TGTKehk6xTrpK
BurirwaNzuPgz7031P+HTcbpUyq1SVTcJrzWyY4ZVk0SlRAWsIXgFBENYiQRfi90
r6Y8c141q4yb/RQClPO4GMCI0Ou5lfncLTthRniUAx7OERO0Pgk+u+IgGXq6NcaA
pceUeTNh1IkkhXl6RK0ZaQOrt0xGsYoDIhRe9AHu8Yp3feq/tAdZCldrc/9jjkNR
7NwLMXSot7pkaySBI+HD/MSkEjQXNZqMNLXLl8Z4H77BwewMt/DRD8EKh1NVgG5j
nawFWurerlaqF4g/jyCRITweI4rb+uQGYRllsdyxLi4vEWg8eRsDHxUAVEfsyH8a
0tThXu3/tq34Ff7ZlRqulPJF5/ZRQMx/6UZeAb1aia7xFYttZUyQRRdmh1Dqrk72
bXZFjMwGMq1JExclVIIAmKw8zf01moFKFc7NT0A3ThR0aKDOX58zvvVpDo65gl0C
M/yF5dgzSXcamZMaKeGgr3sHFqsTOtDsOgY6ZSDm+bgFkZ613XpTsI5G7fY7q0a5
rLGR2e4l9zKFMr9hHGHhrU9cuu/d6/Lxml5BOGXDOiHw5bP8A/iv2f4W8r+vcqA7
NeomVVJ23z2XeV6RwTHR0CufRsX7aB30MrWQ15WqZVFDI7boC1WJ46MJauzsg6OL
jn0z+Fe+0JYnFYm523o071kgUb2DVOsT3zSBMAdTS/kp1wyMXUgSslyQng4s4ctE
Ul/uedrqccWDwf5qS932jdDXlayN1nYLH6EIvGi1dQM1bXrT1F555UG3kRAzfN5w
fisHLf8TJTmmQ41Wa/6mAlsSEPvhFUOmUGZmKroAqSYoBgKpZEPH/0D07PJyuXI1
9GxFavjtzn5AysAJ0Q8SXVYh2UgGT4c7mohpnpCA5hr1evJOViM21qDbRwWExJC2
7iBibCZmusonKMG5XRZ5Fhcuq6O5oBFscmDNj+lxK10+/uX9zke0eQAfRPYvTuNK
svmMmXNuKu/wyI4QMT+stU6yEbrwZwBd7Rc2Z61ndvXbdIEoP812LTHvLENC51N7
22UBIzKTVRdO03+tAC35rClg4QCNIgKIeRW4SS98UFB8m6JfR3erqoUEV+o2w19g
H53nVxa1AvA8c/xfJUc5DTtsykSibX5PpjS+/DhEIBiv949Q/Htbqff80o+jdTJK
OPCNk8YLG37IpLxoJFFjY15I9+ZU8dfA0Rv3iwGYRcmtptFBjfh+tDFHnO46dNdF
3E6jxNDTwmWXpffyAsms6SS72yy1kS1Y/MjkXfp63e3J6/miEevAXJ8Vd7sIZWZS
LMIHRbSJX0giYIYvmN+cFGjH7Egf+4Lk8XhMCHSWEH2J3wdBOtKMm5rYn/CtPpw7
6fb92yZhrWpZiu0gHCT583MfpoDsjPAuOmC++MXqImQZ7H0kMqYEuaVqis1RdS5q
Eo4F1FjVDgs0CeIU5YmQYYZEDzqOhLyxH4t6/Y7p5WYtvfV0YJvAm/z90bo5ZGfA
/6cLv9IulQSo1T7+US367n6ojH32RSGncE3uLUo9R0EZextpRkz326sXMwQHZ5zI
O+8DIf9KXq+FrULo/QMICWJ+hyEwQL0YwP9dZ5KgXjV/I8eilYWwpm7NL+YQAaUI
/tTA6uP9fV8VS+Fd5xEumQjy2LnV/O08sHAL2J4FxXM9FPhTeSVK32t32tAFSFT/
wNtRXwUE04PDUutqIK5J4nIyFYiICY+MPOl8R9SHjL0F3zivQpfPuP8srZ+12PcB
xA/3bkr815lZObM+fTU/JmzvD9yzqrL865J+0Tl5Ldv7GjzFs1Oef45kuUGBNHDX
6xwzlz/GgILRfAbZEhjtzRWZQWSPA1YGcrOHTjvL2b0wwBtdn1aq9HYgSeFEfZ2P
WbGoj1caiHNz3IKzPJ9fga53p2pimWxOFyPQ3PjZMEj6BfTm8ZlrUlLcBX+wYNg8
sqnne6Fr/lsRogMhJHtghcklCsYAnWciVTyqDu/+ZLUqBI80mawRXrO9pSDNTcaE
BX1lBhzlvmnCosZ8pDnZ1l5FP6ZB+xVZfiPNOSGEhkMrWqAYWD+XvmeG9uCBQ1Tg
6kfSS0bryCWxA29lBAT+6bljMoun175teacnPbU9q42hPrn0w77dMAL/wmrZ2+91
wa+14pvKYNfpXssTasTImslKa2yzEbwZD2H6Kv95YEhrMniJKVMaX11e0DAxG0RU
kIX3unyACnJYLZlRbBPxf47mHeACwZMwb2fijZ3X6M3vWlNO8a+Fn8kaR1EAANUi
+X23taeTgxuEupH9bQw48oGvxr/5MOjwlrc+6b23C+DHOvzdwWLUyDyOJgiaNcqs
MeSGSpfdtkKZh1nftI+K5RB7AG4AzP+RBxXMTffA21wrzBlbD9hh6szfHBoUcPM0
8LVMdtS8JMWorYJ3n3TvxbbVhH8yWXWvTBWi1yQvKFF7yv8pvYVoDZ+XarJNAynX
Cyo+DtAOhiV2S+TW/lCa13WLi98/1iMq4ADb/29ePWN8gvm+3LN7pvxosXPaaKkP
kSQra0BMQOBt1dsThRYR2WHZnrGCxed458YEweCjpi00rcYezwv+MziNQrEMEWof
I162TL5Dx7R9nSR/N9uUzARwqzpxNyCEGgbcOoa5aTgsNUzKRFcXBuOlxKRzWeOw
lrOEdqWaHMeOHIxTXR783JsiYTUhdQngb8PzGg9xKYKlHNmhAhPkKzznJ6ZtX4vX
3+GeQsfN3l1WvCgHDymRfiJZLsfjnb4Vk2bbAR4R3iOPqIXq8Ib2LdFiqL1IbPcA
JHVu2LrfAUUtltR6L87lHHlonXpH7hh4X+1C12uyhV4h9dqShGr8lNGEKbd1fIZd
pbbjHYLorsaf//xw0ScAaLtgFCO2AJHScc58zsMjiM9SvYaayy4h/RQ98ajE8Qu0
q5QISckBycH4Yz/QerESUSM/1TdBS36Rzt/TPhI7Uu53rnv/MN4GuQsfB0Ap3tRM
OoQJo1SihLLG1Kno/cRjNIopk/AZNkWpR5DpSZ/OoM9fLNk4AbL/qxmb9qqXj87u
hXQqC0n1BWVTfOf1grdpF6pplXZUlS8UCGB7R7+fanpcECgwsa+TJ4QaddgBCS/d
Rf19QK7FUGOChAZUfUbpi+l/skqtVgcONZME0YPa10wFUSFG8C1NwlCK7NhTEuAT
LVtwT/lmwF2C0wHlX8aoJJ4sL6HGmIWNaXg0tvszXzgUDqELDdkXi4mJOsnCJcap
KHO1nj+Vv8hmEbDzcCZ44Pru3YzKzuzYqg+w4oOcuvpLWdB/VyoPdabVgTnjRwgJ
qZJpFaDZcAzTjLiGiANExlh9jwwa//y6+ekK+NReXRK7gD5XacYzCsJYWjTAdg6J
92b+2lHviJVGs58opRFMazdjC7bugsupm9FS2WWCT+5emVeZLIyEIwgd7tvoS9iW
Ih/OEkYq1nAerXZgAQIB7Bhxd0fxNuyDep0pgJ27iwmR/1GOD7l9AdE2ADLZOC/z
+bJ0MZOKP+GPxJNVBwzL11sYe/xlh/i2GkP0+CSKncMntai++chDdi/M35mdGpWY
LBf9nIbMhQv5yRIM3dbnKUZOBKzaniVrL1FMGqV+dcb6Gh5y0lzO/WzzUKKT1rIo
ELtt62v+vTcPsvfk5vZSqNXoril2l4nwNki2tD46l9njTu3VuUuUxneOFjdxy0At
VVpG+GsriAPRLAS9a7lpuJODDHRW6JJB1JBPoKQpPTRDEbS+du3f+cR+71Kt2hwL
vtfhOa6WkvJjoehA8z8MD/aZlYe0m2gND2zdU0fNhT20QY8u4shqBaG/56Fo82cc
4hoxAuMnv6Zp7dE7CA2td/NxS1duoYl36I/RaJXLT6JezYh2PGhVrBRtPnucLX00
aDJhqvcy6WB9t/eDcH55/sY0MW8GfVHL8vWmLknKYz7vNKdQRwSVv5VbLqErWsha
Ff5I0pdaZ3Fj6HZdfu7MuxJH9pydiet/6StWNjCK5glogJbKFad954AzH6pUcsqY
caZzGIlSkb4AxVBhaiG4pxeasCCo5iVjTKd9dXMAS63jwSxVzQihI9L+lYZYAzxq
za99df8OX65+sjzSM982jYqA8rW86232Zf0oOIJZqqAyaoXvPJUFLRqyDeM2SpZg
t05HOa5EOtt2sgsBn4+8zU8WLVvyLepaVI6AKQrbw93Es6MIBvtfV2bAK+dPkaaY
HkGTrRxqnWF+dK8K/Q4g0J4faG0PhHGCHyY5HL6DaPTeDBFji6jPUjdexjNcX/7V
HdYSdXZB0v7MZaWPcTp5xAsW+ibH27GHRi1ld1EjiKaclcjSPllrSwjm33d3+/z0
zPfozVPZMWX5X7Q/791tYXJBm5e6Qkspi6GCjCKDp6kyBQ5wNmQ/MIC48d8O2Sh/
KWTtFrL7sNsMYiQOFypG701oJrIQQbfDUfvpqcoH8n5PhCFLb63/v/WKqTGDoXV8
rHslY8CNM7ozdYEFXUtz4C3vDxKBs7d9NxfQATpI1LmsSXYHygc2buTLzJ4GYquH
kxBpkXNT7slkfH4vKWGUNeEhprcnhlPtB0b1Ne2wTWdU/Tx84yTmD7MTCFwyBehq
uOId5f57GcyIALkST1Ehegug0XBxfYoiBKOR88tBAePbreXW13ttf1IkbUcGOwll
h6gdO0NtN7eKbIYtHRDeKbs2lnzOBpLBQKuj9bmnIpk9bwwEMIDx9hblzIygykqU
7kYwkbnn799CaEEYCqMX6AFW9cgmNAp8iAUkaXY9jgMf32KWJmH2OEXJut5rc3SD
bz2hQ3vDl+lzkw5aAbcfjELfrJj7zG1JXe7cWvMsqkWh/knis2TP8DA31NSpjZaD
oFqny83VUdWuUWtQ+DP2sQFbu5aBOZ1747s7LAPS7X6tud9epU+Y6Y3gI+mw9B8k
8ZE7WomrDfaB5hzga6OFtite2p6e2n4y1RArziAcArSYhzRcM1WlSl9SgA8Sd1R5
r+LHxKamTKmHhjG5xiae1P3t5zCzSPJlOtok0WYb+IdwOEyUcUsJf1fOTJ9GGqTk
DB2B1S8tsZNhJO+5PUbVC0AX+e5/yWzpaWQwmM/bA/oozif96kuzVOMgtBtAjfcv
BdERipomjcMNrRuicjcP77SqII6tVFdIIEmk73URKUG9QYfKgJy6xLrr/Z5FWyoW
fMGsHXmOKUrMLM54SRGYS7D9IC+h66RgcvoP9+EbW31OlzGYiAUqOaIAqIc4ALzb
UIbaET0arnN08DALLsKb8j+22OANUdTtbZtPgDZLdynECp9U3OGKn9JulWn/9v+1
rdQlQ//xxUOWWfr6WuIRKIeBgPbpWQ5joo07vYHZIct8rYA+48lreFSTJoOTPEfF
4rpX+BfDbN+nb5oHyZixtTKvloAH94G0I4mHptm4fiH1qJzaiJfaF5nAeBOAlL4G
A+9pevGCO7JPO62U+2gWaVN3rei71GvRIANOO+9RT/z4hd2o0qkcoKjsBb2FHsCM
7jrLziUJ5n22Flyi+y8AHz2ub1H9Zm40aTDHaYvyadPpRx+9aEj7urbXKuQLkyMe
3MDKM5i5oGgrc1i92G2UwoWLMm3f81HHkQjcb4kcuaPzSfUYwku70yWXtR+sA29/
zG9pjEsg9cP8qjQrXf++ey4knFo02j5y+ILIQRkw2WT2LFPsAr2xowje5nfuT/Hk
496Ypo0T71JlkshuE6x++DKstDrDp5ZrMytSrqNMgFwxB778n6khsArHmmHnbfyk
vTg2WHquIfWJhk6faPlqea8kmd0ftox2u5cR04eLjKhaYpi7aNedLgAfeB9lnJAD
JM4Es8320tSV/Zm0Ygrb4ofzmJmbgi3x9iCxn7R5O4nrwPsDPMpAy7aBToANszp5
uj0QpVsOay/c/T6ERv5W03Q6gQDTE3puHlKb0ypNln9RU6gUq+E0pgVnM2jGOf+D
+ZzzCwtPkGOPqHwUHrAdI62e+3n1fS/XBX+zoDEAzu/adctFVDq7meICd8/W9Ilw
bWh1gqInTN4qxRRWcVINP3TGLG5uWqnLzFyeYD+Uy5K9jvindLPgAJfXK8Md73SF
sKRfqaf6c5y/qCHcwJlg7p/c3wu3SY216HVeXuhzZde3/T7WwHZ21o5h8w5gwYxY
817yehGmiSzZTuAr33x0bU3VJ0B8xsoaKMefed3kKn1BO/84cvywnrjEutBp8hga
u8KYsZoEqGFt+EXBdaKSAbhN1GQJAtEtlmLnQL7Al3KNf6sPrH5I0iBZcDksNa2A
sGnp9HPcioP47qVMbKaZYexMJNLpmoQNxgdlrYwwFOLXfeH5BtKSVRy7k2sxkQ16
2/22NhPoxOze0dkDvTg6l+8OFheK2TugedDFdsFOltA2fwXsiqtIXNJVmgikdau8
z8iN/b2DmCuVgRTJQSnOYzLD2x+feLtObgb0RswG8AGANWl8ArKg6139maW1nLIs
NbinLwiDwQUH5zAiZ92iCRTFffdvehID9YFevh6s5XRqaRCuadSg8feUWkPqY4Pv
4TyTW68msqM13Pjm1NITBtVYZ16fy3AS0WMG8oPqocWNSg4R/WksQMQQw++MWFju
xvtFonheKZaitEmKGJzXUQLFDMJXukEWqAW77wpSmhTrNmYfbH5s8wnckU2o9nGx
Dxk2HDQFbsLoexynBfR4WuI8FpG6vgETeVAjxRHE4/9SJihnNjLmPjguZrTJvj/H
anWpabvASMk/eEaNRUDJ7ohv+qCRBHVBWsWY56Ohg7c4ZkmXYjeFyEsXMs5ShqH7
fTx0oXFwE4EljMmpXwnctbeECCQ8uXWxo7uH0oWFa1XAGztyRAX0zv2DHTmlTEzQ
Tt+rID7HXcJRtq+IEDZrCi3y7v8QZEkCzwkQu8UyHRhU+tuCrLxbUgxGTef4cic5
do0MgTWCcZaTHST1ftmkBklUikWadeWeHadnGzHMFx7Urbl9AId1pQnsEcpFJjdi
jnx8Qmoonmo7F+UbL3NQ2FLYmZC04G6YsBa79JD91mXKtvHqte1JKcvkwyksC3XD
h/mBBWpLtdqSEzcfwVejIrapG0euLOgqIqIvqbvfOB5Nj8EL0VVC7dRaDG9s5Uis
IWqxxrMxGt96wg2Woph/kYZPK3OvoUXoXSLOwc8ZY4zDTZQT3cvjqpnpmTXEuPUr
madOXP6f2Wt2VNtVbithpW6uYE6OJqpicl+oD/qI1ZNjAg9bbTsbvJtDyxn+xiQ4
sW2udwR52Fc1DjLDj7m85eF0C1SJg7Sm5XCxv7pl26FeSIeGD6CA99QlPZKz6Uob
jKiULhIxanYdInd1JDprMmCpirDVR3PlThRFcDHYmwVCz4UhTHIp0dbnY7DHGoql
2s3g50VIyhJOx0/qGC87TI84yD+AqoFkIq7Lxs874vo0OJctsji2dlvn2o7PYUld
eY4W0wviq+Klh9ir/68agwkqZrBevOvMmP0aPy3hJSXthaLsdzSex3B+iwgFKiu9
+B8ko/fFzAzk8KWvnfAU8AQaXkuAkROKHqoZ/Wknyvp3CZCWxiMBiAcuhxnrclSx
r5kNbBbu8rLxgEGNzqNQJa9LPhqEFkXK/NdH9BEOFV7xUYRzF6wi26BPE3MxTOgv
CpAMtDGjU+DCNANWglMkV7Zil9jsY3Z39W3BkMDM9IQv5pTZzwz1CFJ8s+yAREB8
DHQpuQWTmd63LqlTMMeMdbkED6D2KtMMYQhJQTeLgGXPmriFEys2pppl2IFjapjA
4jRiinFDheG+wQrk1q0YVQJs78rTsmTZM9Yxdw6txbVbJg4m/6KP5S+1/wVVUJ7D
IgzlRlioaMCCKSeIaK1mFS55m13BdKYnHAiJa+NXchlBNLZ1wEcGuyd5m2r0cw4r
Fcxrf3BHP91Nw5d/Dbks9eN/12YXQHKLVxLNlffmFmSJevuu4GzLn5CyvHJBCXPU
S2ELCkC7HYdigKCEneNsQwwynV5Or/ZyrZfyZSukbjce5y9Diej5A1cERsB9UdPA
0TU1gAjwqz5GUr54kGs+/SZGMrGn/yDz8Ytw+CnFEivunQv0u56p2xriKLP7gWV2
jKu3ej9SjsX/iO43L3k1d4TqgHiBgh35A2bmThHENl/8LZ6asoEApPyxJqSItl4r
8LtBjs/NvoIMJkTR96JFcmB+vgXd93Of42I9TGKS/ezZxZ1ClRfxFp8I+xTAmVt7
/C5hZy7fkfsUaM2CvF9t5klKrosnNMGNs+Evm1ugfq44Y+RdnBdkK38ZEFoLLz8q
xdET8glCXTfbNPbWpKCuCWAszpU31J7IDJJ5o87s5Ipnm308ApXlQg5LhMSGqdN8
9lvKLjhMdXGIuLjGgSoX6HF7or+twNY5bokmWruE3v0JRNQqFNaMRu+MUXIzDCxD
PjZDGmUWoOd7E0vNz6KeSi4vxGXS3gunnLSnolMANqpAV8DQ0mYQTfdQleyNCzQM
XBm3Uxw8jNMdElFfWWYFkdFxP70BD+oQj7mkiAth0r9QMy6Vj78hI4zrhZP9NFMk
xhAdPe8Bk3/dABujtHfCB1l1yd6E/sCTYgiD6giazA1YsiGFlTZfhZ4oGGJOC2VU
toG+kWLlqQ+oXY8p01TdOTInjvkLTE4evdyIfLyhMm4gpFXhc8yNq9xDjCgr82Sh
621nA/aAZgUu/RLJcP4aiXfuZPI+57Hrl6vnJlErPTfp6QEttPDya4RyhNDfug5S
TI5Sli2NywrivggzeOIIGmO+QJujPFom1wD6p+22B+WlO6Te7D9qvQLKyLQXT2QM
ZT7Pr5G8xvtEOd687V0VSWsmyQW3+oeVxn88X3CKhS+Tw5bvevUNiquabQE7xK4C
e7Ghl91CBKG0GI1BWQxHb0C+FGFZlPTyJvsPfpduaiAmOyL2umb3KAppO52tjOrp
r0d4ECcf3rsHg0mIvM117ldZ2L4OrzJoixJM0HAw4Vy+Rz/aahsbzeEZTu0j22sO
ah7R5LA4wESyRx9pzDVXg+nNqtZpthITG3/NqXD2sH0uWQbS3R7gOB+YkoIEXmLZ
cQYorzNOKK9pycB0SosFsmIGNYGvK/n9I4/9ax0euyBn5y5traOXbIB0WOC+h2OH
zeJ1YrzFsBYCPAn4oE7SCPGS2uXECbIvPde6Xz+/9XdxJbozBJgM4O8WViwGfxoH
GsZ3HmYvlBcGYEaXi0dn8UUjLe8QzdiI5e3+eXJIHYN8mSchqIT6DkJ/lGjRi9ZY
9K+wSQ18hUIUMWEPi64kl3nv5tL1UeIYlHJJyB5NHmiQmloFluQTmp+hblxnrv+Q
Mzq22tp22GOFvXW5wSvaLZjipUVJOAxwZWD9yYvjs8S3s4iTCXg5FiOXC5mYX1Om
V4b9Psqs4g7zKz696oazC8Q126N/Lo31cTKEFqiBp+ohvlaIP/5rK5bS2lNk+haU
y6qRsur5b8FrDYB3ZWfJ3y3UU+g0CmOXyELJagV5ASqZ8prt/t3gXcaiqsX9TmZY
Lo+D70pgrdJA/20aZjbTGJ5Ko9iJ1PO74OS2GOPPa5wi9f1naoJjzvdYPXZDUgUy
dJuGtZOesrek6cjpIKW+IO5U244hwMmeyD38MDLPqyn9SinRDd180U85d5pHSwn/
kXKh/nKEU1ODVz7c33yFNtKYr2WZcbsogP9H/jcYY26PEW4UVyhpG4jCppo3X0Dn
RXUnHcy3fzldmJH+hzec7CAUK1pdWVfs+jYWwvlE4kHNB3y4giu3V3pIy98d1/qI
o9otuL5i0KiX8GOFsTCMC5Rbxd8pfu0XT67xHOcXjiVuITIdcuJG6OY9hkb619Nk
PzV4Si2FGdDMnKhIY6oZDKo/RQ6Yv8TXLewQM/fw+jUETn+MJ4iT/cYxxHAmdP4R
ssarc/RalzjrRzRet9gPQD+mkUyCPu2Xo+ncaaCGzRoFLvDZAfdR2KmZAf2o475u
jmnBtvd6cAkDPBbFpurXuYPQoe5PMcFswExqPFvb09tm2VKmJ2gp6K/sMyxFsu85
ux0jT8pAgynO81si7XUXscF0cMGGIhpf8I2cXtvv4vHcku9YKqmr0d50vdq30ElZ
Q92dnOFxJwi5i2u/qX98hFMw4Nv4GuHPMVHqQ3+YZ8ioI+RxdMNXmodYXHa93ZsT
xiDjXPPvhWoNZjqOaBWbNKwTaYjdhG8kb+9oWxCla5lgQmmPo0mAu4LoJmccHdPT
gBb4P17KCqB0VPN+pSU8Bvln4SmvZtkuzkJtQUhj89j+lXoXEX86BZwg2fiuTHEk
fwwdCcN+Z0flPdiz+Y4Pc7WTam0p0KJA4ioghJK53jbZbAub1TQ3NTdOZ5jbBEw2
jlON78nzrxGG0rwWtUl5H+s4Jc1My4AfqurqSElIWuDwdnSJpQC5TNVLYy4BGgYj
6eVq8bH+fVWfpqc/yHWxD1sVjhsUIUZ5PwEUJ7KfLSqOCoOHY2o+wvtAks0QdwzU
KuargoqPgUsiQn5cmshfaceKPpVGY/o5yL+bp2x4kmk8gMZInLVsr9RY51LukYm+
A1bOxP4raxi7Ke3xb8zBYP72bqXiiV7cMT7zl5ndHS9weKCouX0qOYvdM8V+UNyj
OhO6PW7Sl5IQ1RVw9mKcNKYmPe0zxQBx4YOpQSt5uSxLnUSNKq+G2hXz7SM1EiMJ
iffC2HzW4rU/JSwKSHGdyBXF0lPJHDDnllAgngAj7OAdPBTEfR0y4DIkiGRKEqN9
lIGHEZdx1nAUiP7o1Yy9fCoVnBX+lhJM2pGqJ0QA8uS47/4DG2PvuTYXVx1Re/Uc
Vku0vrdYykG5uCaWgRJDtGctQpLBVIaaYyTvWOGqWJ6aDmWElPFIvdKxRi3G/fFq
WcGK1HawZIRRJ86mU+grXx9e2P+M6gM3O2M9Mpr7QMNpa8SHthREeVcUp5butnGA
A6y3ywD6FZfvsCs18vvTyItcjcnY6ZGd46mD8UUgcUU02dKyslx+YdJO28GJbMPv
IaQP21jZmEOxOD1sUJvKlr+78ArQv+zwNiriBDY6IdHXN4zDwZcBpGGUH1eJy0Pc
Nx1LS+b93Brw7UQWejm2axwTWauipFfLMtpYYT/xjpwXpbYvUEJuLWPi0lwkpXpq
TCfa3FQaD9t5gAwg4Kp8cMIJ/2GaMzWn8J3ZMhNv4I0/oJYB5lVL4O9md+5UAvXC
Ro7dewE3OZs7sb8CuEL34DYNbaTAktsEg7TpXBUMobYBFnZhUGCTcdRPvzkYAimr
HhzdUYe6SuZOYaWdQSKns3YP4obXSEFChAzYpAxkYybr0huFKG2jyyqQzG4Txn9a
TvAmRgN6CQ5cj5iT9ULYHDWfpZzeXV0+KYcA/6ndaYpDXvFu2FKPbmK+w3emxzGT
gzoDn+1orSUeiYtXKDcVDbFUooF1B2MFdbdQkaBnaMo016SkIDQn+pql/TLDlQS/
U0qgA3N6cSHxIksisqJHOESSwY7jHMGAuGaYyJfm7yNtukwPZpQP9Cj7ky9fNOFP
Rqjqo3g0HPo4ZYBBDG6nIVus/M0rGcrw5Hl+oWy5seLFRwdolJ1LfIiiIuOBxtnC
IkJ/G09LYa6fcxxJL9+JEpyWzKCkCTScdjRdTcmneN1cJTby5tyxpCG7r7FHuPZd
pUZQVnaeE3vi1vV9cEdRLM7n0dlGnpuv9dbZd1mB7yhOqiDMTE01XmSmHmdTpfX2
0KSqjo6AC/HCgoP5olsfxfyPtZrC5dmd0CmsBRpgkM5aMtCg9wAd58ml/Y0yRsnt
fsx2Zdl3XrwxXSuxRl5rCTy+1mUH06IRbpzY3Q3qlZGnWvfpqOGBcAK5DtQ3/SW1
JTGcqFCJb1A7TBTmq3JyL8FL4WUpOoQ4dBxgzgUz+ce1CuApKDDBStnepw6brpZP
ewE3qRMdkhVX0UcyGrmUIiEclhU1MNfLhcoztQv0D8AEzW3aI0vhZoTiPo188Hrr
FaccsxDucJ+BxgJo+9S+razwoTJAws1IQfqMAmNX6HzMufco/mwsEB75bS/0GUnt
cn9q9LcDdQCFzWewBD9GFrFGnWejgNpBE0ayUQ/7PW2jhWq/V6fe1YG15bvS3rIF
2FIPErZFd2Vpgk03KutIT8/cA5546iU6xVqfOEp5n/CpRZzuMlhiH9NjiaMhPy+M
UmKMQbFkv4tBtGHEbLuvTUIF6F/IEkO5zexgubN+V2tKbSahWHZxhgGWFF/+H6JP
idDyRmNQreWj+gXQNjQ+Fua0Vwl2DQcpHEr+RdhMtpyZez9xJKIHFRyMxncz+BBr
Y60qYxL8xhvHrbcGROd0bXrfutOPM6C9aAy+bhKsQZTno4V7/56u83z2DpJP20nr
fEJAXAz78Ve79phDCT3wO/ppoMTCbhmKcqgEn4UOPenUA63MktD9B2EUGWw2ju83
rqhxr+qYeJsKyhL1ug3/o95FXi+V5jg2UDM60bkJFf2IijhR13lTGxGHmMggdZiW
O33pYLN6ro2vA/Ua0e3NekLxwmwA1jyHgRP7bY1XRgBPiwuibnuGrhqCgm89Qv4P
hpzpL5smREgKz2xacgAIAl8jG6M2wLrugH7roycSG9gh0EJWXO0wKxwWLTtgclVm
Eo2sxi4nvfKPF2Hjtlxwr3KT+zi7GVjxA0DAUMzbeDmlBz2FU6hK5Q6kGIsFeDIB
Y8OLwyMRXIpb3YMRAToUHrIqNNGuacbRyKF+Sp0sTqOX/RLizP7xPFG4bKWFwwD+
YK/rKtbaHbn/fq8ZyGS6Z6ZRY2q69WTpzJoGEvBPo/i71c5DOX09YdEFBvJ274Bb
HdIgpqcqMXigduoKAeCLX3+Jo3IlYn3zpCSzpeKmBjg/NgcQF/lnR4YYag4mPyeY
VrvePhGGcqspUiby3O1BkWh3uhqJh+j7ATAe1OEY6cmAS2xSuAWM1+thydnjSz2S
ZWrb3WUV8I4mb6bkE4Sda92kDxSCnVEutDgsNi0WfBBeYVjAqot+EfghObyNOr86
h7a+r9IomSUEDBwA/YL7a/lyYvpeo77mTl1lzVvVMFFJzRwPYhlCdzuQQoluEiJM
tUlCY+udY9qJLf7BK7s4JlPoVPIlqq9urG7Dof9SVVZfGgeJXhAeV05kNURu7bUl
T2QiGRDFkFCO3h6otGP8zchGfDo/XmPeC4ZwpvFu7Ejw5Jz/9d9az1KbBaqdY8Xd
IFXrgOElHVMjgpTbC3KuRjw96RVLKi5YdEGlRcuKHAKXVHIM7IlJlv4on0xGntM5
hDppU6HsOB5nhdDkiX1H7TcEVPNh9kUfB3wlrmk1OQC4TXfv22zr0TvcQ4sVG1Z2
u1AWnjOL1DwuY1qkE6ykbWL4oVcTH7DYlFpySbuWXLpFRUhht5TF01nx0lXfBq/W
Kh8pZPJFgMLM788c2jkKw2YFdvgjD8TKuLKkv/lxVmANFjueco7EKRw5WQOOenoz
bq17lQTTTUp6sN91E4mITWAnuWWeXjXwKw/peb6xPCqlv3pV5PjzUlDapxyOsshi
GhUlnCbO0QHj85ZWGCrY00sOdcTzpljKg8LXKLZfNitPvy9tSE9+zSj3SP/KhU2S
3tOzjI9duMIzQxoXaRlEQFd1rywUTNdur3o38zkcxEf3elwgBpkTaRMNqSUjgSDm
hcmHFgGuSwY8erFaazqhb6nXHn3dq02CXTaGwFYKcrG3g6EkQcVcVE/V0BkiepHt
kiYUluAZkl9ahxw/mUjZf68j3s12+xgeU6nIcaT7+QLofifnCKJbY9ee2i74ob2L
/2XYy0idfTv7PUrzOKWIViHvLibvAmyCMjHxLQVtYGpM+mXMPBNtYM+PACncDZer
2VerRzFjgXmNDpWYTlO1fxX5U72MUILHG/DjQPVckwwgGvg34U9Sy1oFahKIanx0
IxhwWKthnSIk5mPtFte5ULlq90LByb5ilQ7wbE2D5xa3UlXlUaSR65zJvTZO3jEM
jec6AWe2df+Q4+Lq0j8nOhX2QTh8ZMjfpDcdIW+r7cKjKZ1DH//l1BTtu4w7zcU0
foIGTwKrBDwBjgUNgmuYYpkFglKrfF/wYG3Dn4/TWLxQVWpDXPGo7UMPlpPSnfsD
Kuzmdm+yjamg+TR1d6/5Eauo9MC3HhEW9/vH4vWI/eaXmDpl/fagHT8AsxcTmzb2
MHEMKzyXd50dZusHYr4Zu9NdkhJh/tFYqXAvOTYVB1cxPRUg2dn05QIukErSiHK9
qarBdObANfAx1tcsuVKQyjimMvruc3leGOoTDBLxlcrn7ZnVKOsTQeaPaQ9ueY7V
vMdhAnwdp2TDxCxrbETxI3vKEwVA3UxRud+ib/ew9+dRXdG6HC42KMHolbssJdst
MT8VluDmBs6i34AfJJVgHv0SkbCUkdD6OYwbOmAo1OjjImsqBMQ27gumTAVD1GaI
mEkiA63NpNpGwCMG4zFIJiXU6yJa3x38JuYEplwtzf0WvHMDxAwU/OPo/0SnOQZu
AwhiN6DfDjwAqihPJiPpWt7aMD9D1UTQsTTM4kWHD9iWe9v0170tmeZvJHM03mNh
D3WogxTwWax6CMsWm7UPN43TidyB75kS6S9/vAgSxe6X317a8S4zqbFsXD0Ll8qR
0fl4YKlGs4sEFmZ4OUpqTl4Ab09tW51NmL1KdAuSOkgOTkPo6B8xOepndgKd9/wA
1lV1WfZOfq3MYdvQm6kqfTJijruns7B73KMilqCFi5hj3ETF/zqzeeycF1rKp46H
xqTl6K8PM2jq88XwdWPIKBXL7FQRgRHeZy4Yih18xwvVR1OKl8krp721kxEmmpQV
wcvhwCITLUaa0GINkEjYL4amdOr2f4sdKcfgdRN7wxzgUI6sTWVdmsDdFFAVQ4sx
LWB5fMsOwMbADTgSIk8enRRUb6sH9N/f2qo3TJkN+cqgw3rP9JRQLcENO7qHbzUY
4NrVs3zg+b3WBGwODMaM8OHqbzetbfnUdmiMFj5J1zisNWtKmD2/lPDxrW6nSLfH
TQ/QkMMJrzFE2AMXNM+zhIe20xVlCGXYKhk8wm863BjOzo+6lqstNjMEKhLN0486
AOwrDbpANAveOYivm4U4FyqGZOXvF8522cJRcM2r+76CqwiCNNVk6FmdjuxIoEMe
qIN9sPVjWIXCqvweTzPxJFO6oD1wCyfJBLHVbLCObfkzZE9vkxVrky8d/BkN+GNB
ISEA11v3glpj4tsHjm3jXkYrzZ6ZZZchpPCtLqvKH9dq2x4tFpcfz7DHqV9g+iUO
BnwpCyKsPoizpR4Yb62RY+sfSJf6x6jWz36x/XdbcGDW7174JpPsWpLiJ484uLMd
MEBHPvaeO5lHFw0Mtf5/iDU/Jcp6SwfQQ5ome7N6UmA6ovsMH48+Er8nLPM+UHVI
wX+DvMhsFB3DE2TjlaF6047l+YDjnj2pAgnQzQI+spXPL3SazD9h+6UNjysoE3In
oAJ36Gxl+/tM7XQAT5+kn3dYQDwOnYcTS38rwfMrKsBdqzDzYf/52DM5YrLIf0hk
oEmuvnK5n2cmBnCRmtOOEYvdcfMWtSKMOabAv37YbKDJssawKHggJ9tAn8SI1ZTs
ywB/bhPt1oSTSPGi7yZ7qOI1EY363cnMhsbXu5gaCOd1UJU8tbIxevqLpf3qgSHm
9trnA2g8Sz/sR1juUR+ZtSOO5OBQEA2gQJOEk818yyrRsKPSJlPkTK6B90RX/ynr
tZQ8J0NjLNrxj2MZa0ZsOiK1t06NJoJ/8NgpVngsh7NHcFmzeI0Ht+c6tM2j/kuw
z/Z1OPQbUFopHHJ0czG/KAv0TIDkoT0C32qvTZZaUwncvhqD/2+lwUaNY8YznFuS
O3d1IW/XpqOCgFSETOMS9Ck01kQL1oqVMkP5xjOCN0T3MZfWO92wt0YbZlcLdeHC
tt28i0CoqY2sgnrN7tAXVYIIpngxGe5hq/0ijy/A48g+mQKxLWtgV0tKfut5D5ql
LWus69eKrdTNjYm0eC8LomNPZqzntz0u3VJEV1gRANX9j9r7Oc0ApP+PObucw9mO
C4wDZ9AgOiHw0WBHoPVCheJXt/ZAjAXWK3F/bUIZReYj6htJfkxAEtBnFJB/VXGT
Nvztz0x00KU22mvYaaTPwkKQtjL4m2eij76bliLmXA6tIGWUqKQ5+l6ymPzHwekN
trq5hN6SRIfS56X5+VGZLF82b2pjWev9wTArv2s5I7Xj0t1Z666I21NIeCH/CqZm
jMnNjAUq3QsX3by2fHlV4VNT27l+bzeT/4SFacvZzuLDq0rOJ0qO+FGcRNNZ1tm8
uh9Wr3iWL8xdMIlDud2o2elqb2aTCzZqW6HLWQd2WZKywUf2YgRolSnm/MhEJymR
8hm/TzgBxT7kVkE4cUHdt6ShAxybNZAwZZUGezvoY6fTwfq8K5LI/njZKREf/6ab
hFcLNvRLcap4BMV3eW0on4UoxnfGK+/pv+qQk0roSza3VGslU3RNPtjs1rELkBun
9O4hgJl8297zJQj5rgCSZDnGLqJPWA4NF23idsrM7xVICkBxSebtUdDMHP40F5d4
F38AMRruZg+sHH/mCyj5Vg9hWcL6cZr/FdGmvsbW34uazd7vyV7q3hZd6G2cZgYD
x4ehpJesy5udKCQPoFo/Kuw2xOCQVvsqYoGNyDBnOdsnVuJsdjDWY0ZdjVGKsmNk
qlIYAh8RNVXtdc6+rcKAYB3RvV3mTVXYSHYxCAkBbr2Sla8yvE+3U1ifPecEnJlU
H2Dfpk3Kf25Q0hD/Uawc9B+bR5lf1j2b4lu0hR5Tl8w0vexNFYQzQRGM1MbHEAYZ
kJK8CD86gQgI5Pq+HkVAMeiGODmVRAGVR3qEnfcyYD8JAlQcwBNtQ5hcHFDQOgzV
LX6YETM0nb6p36TIfQWAw3NIkee0q2sMPHOEi6DDZaNy2b0Qi6IAeAStJ3ofRodn
QvLkUoO9V1CFEDGJ8FkRC9c1/4M7wncfisbYqt7qm9FTrUpq4u9PeIUU1NrXqvHY
l4GiVn2M9HMjySL32tIE0YX2Z7gwOF1uCK/AlzNBOiav3pVLapEOuUaDOLsFp88M
13OMEJlz21k6EcgVWdcHGrkq3DrZdQLKzTYcIVW76HlzFFrEuF+galdXKaYIcIDu
wJ1r7kDfaLHUsjyCRQoTEk4yKDk0FLh0sWV//FUUkI1XD8P6obBfrcWr/yLAi1fi
pSh9Q1CC3Bma2Q1SzGFRIwrfCqhxXhKi3h3IAwuamucwt0cTgBcALRytImf/Eh5p
bTxeQyEu3fdqfNJAyM4yKSQlJeQ2tnM1WmY0zwj9Zi/fog62Gt6Fv7I5SNR8OaEy
TjT0vgysZLpMracH95Y4VEE9J3pRVUUNJFLk/4i9ofUhnLRKt1uNgHHKufHwFHW3
pH8lw2hm6CW0hnB8jhwR88CrQ9JrWF/FIdAHhxHMPRr3dmbrk4HTp52opIJgtplD
UduKoCDX9nyd0THPX7AkIXCh5VqFOE9/3F4SEaPNQRH7G1V5GTPgsAb9yeh7JPp4
ckBONpkmQzdBQwdClfhRfcNoAVQT8nw6bh/NJ5Qz4urmqZete8z+4yXJmqw6Jf/4
u3MQIDyi1biMQ2W9AZDOciADVbReEBcKocDbBWtW9b6OGoeJmXX6BGfZ8bFRc/08
QiuTEOCaTZ6bVL9KZNLnVmLubyWKXECRTGlR7q0z+JPR7vbLOZZzHCYiNtToSzCL
Ta23M/dFI5/6rTVCRxyjvqxpWU+uQYIotNk+4Dq8kc9XBiZYX4h0erf99+hlztKD
BJxYu2stN6RaR6cxG3pa+f2Ujm/e7Y8ZWcoaQEOPl22tfDS90PGhrXu4L65KvKPU
5nFTxPV5/FxNPvborKpIXPaug69+acHb5Q/yzZoxh4Xls8nSheJhZg5JpBkOzXjx
+LK6GZuNghS7FDGYB92HcXNbNUPOxT3kFu6hM2f8vZhz+aiXITIE3FQ9lLhx7OQB
thxFI4gNq+yJPKA85FzzKHhYArahg4jEaX7e3uj+CP0srGU5LQnoQAHAEFnRAe2M
jdVtbnsAUgwKAWyeLpzY7F/qDbvSdAn5B9wYoHYLUg+nbOIShhx/1Cs6+SUpn1Ji
O8k+x2X5AtbmJczdAEW70MH7yOzqc96AYN1NZpikOWcOTuesD3bUdn7Md6+VhGyV
5z/o3WrNotANuZFYzejROjooW+q3+JY/oT2GN18SFekiak2Roj5OgIYzLQNtJzCy
AQTyVOHj0P0krdqwrYufrnfuM/vSysSEEjPheNGf2flRqmCqkG1GMzS1mfI6h288
iWx67tlZVMZcJGmra4pV3iTTlZcrqLV8moJEk1Q/VLnmji5STNait+AW2wZZviD1
UVeK+TfAt0bnc76o2pOV4LLIXakVYVHbTu/QXkPOkg49o+orD7P+hoe2E0cyRS21
TaUAw8zRGGnj03iE5RTzdQ48b05Wj8ZDUay+B0x//ebAs676DaFONnjyk60wsNvY
KZAjSHTc92C1dMpg2k/DLQWm0naPpR5ZF8RGGQulY26VpIFI1ErfPH5sikPze5MO
quyg7lroyP1IHLO4CmW5ayxRl+1z0nV00I28w1yUfPP+yEzoGV/vlxZ82rmwj536
ylD399GoJih9/l4PFUJTVPbsVzNCOfD1mBc7X5GHegC8OouApbNXmZpNDPAdvHFg
sYHaWF45YgUkABE/1vK84x4DYGz4fvDynCKovY7AXUkWRO5nrvo+S3bh5QhNEeLz
LAelD/hbapu3vNoAJ2lgI2aVlw/wzHZeag406/w/w4j0zc6/6J5MGC0+8W7uH/Ep
gJU62HEHqtOhFOh5j7GWe5j0t+7FsZCH+0fr2TgX1b7A93HaW+esHvbO2Pz9ievw
UJyt4ZRX+Cxc9bIm+n/4t0UehfoWpoZ2/p6LKGaF2y7k/10MqVF/XyKpAiUXcI9L
vb7OqAAmUbghm9SoTCxxRfDKigrUnq7AJjPb9hX+TcpIX6BlmNU0K9tHjJoThLFN
u2QYZ0O5PetkKjz4hAuzzAKRBaar5CuqavWwqcD5AY3qmNZY3rR9wLrqNgprZwB6
wv300Z+sCTFjPQS2d1gUKRfBT2kSuJpFtH0tQaNSfPmEdCCllJOFWpDxLMK63FdS
G8HIes4u7W7C6Vgm5EnujPG70nWRPGYvaQ4nHjyQGpl1lSroJtfz95kN99cgovb3
FcezwlMIBf+m0NXYWzQVjGGXKvFyyHluZfm+SXWI4mQpOn0iUw5DOiCz9Ws40QRB
2tomx0LXFWQ9yrLAWnjH09N8cwHmdjaRR7hq/a2GO8kjhocTYEZF9Zngp2lIzrBK
AYPdcBNX8r0z+dJoKcapSEOQNYU8BuIsLE7oE2rbh74rBzj7gwdEZ6UwvNxyj14+
Xv5cedmj4YjaKLdsAbjhxJRyXDnlVFNDMFvSTVMzp6Dah80Lvb1O2OzJlF5Ccsoo
loMPWpSSdQFnZx1THuQEfILtFMdwJFhbxNCo4cMb8a5omKGPEYI1bsubUP3pDJ1Y
gCFZvxjzpqkk7eMzFeta1m0rAF4JoPeO0HZv69FjSB0y523Zvwc9D8zj+GV96oRO
CWv5Loy/Agt5/6zObNML5ZyOqgyVkD6oMY4H/FHTinsEe2tXicAD2oh9FOezxMJp
Dsy/q08RxvYru5e9rlSybS08pZuclNDQyWRlWbvE5bJxLIvMqcL99+miQE8Nizh9
wX9QsSL2RjPKTdQaWawcNrbUUgu2w3QQeGwmqF7lhGkPc1U8ZBGWsqYgAqRNgLcR
ymHTsYvdls8be4Ak7DUtU4vilQZ0D4scOggq8DKfWPhQDObNbRQk/McNoN5e2C12
6LX7rkL9Oz1giVmmGlSK4nQS2gBgb6qYTCuXQ2DGBRLOXye/CUvDtuzwZGNiAYeR
lFYVumlyVSHfXy742dEPaChqw9sksSpgnFtsQiItyhY0ejiW2CL/1nMLtBKzYWj9
Cgs/hdplodGEWP/VRpnwt8N80ZLiXqCsmA/DgAD9MMIfjq9pJ7MYA1e6zGGS7vdP
tw4lvR3eOufx4vpxAtXmI0HpuHlPY1nPlNSDq8F9BLM1cp0FdQaSlO2or/DTsyxk
6a8IuA99uMkwjzcBSPyBQ5+aSdftbbyiMenqikjHu4WBq6t0LjGBE8W3QG86AEY/
W9fKe7l32Hsn0dZXgjtktqaGy0VmuG/AjlQ/t/DGuOrrkxbUnU1e+KNyYl0wM28I
I9F4bS+/leVn+cILlLm8NOc0cu/aFruE9Ozafo4PIqRA0SuAPq03A5ZOby/2QH59
Hq0C473k3SwY8ucz9g2VbaVevnGSeNu5BsYtpBz7BVNOlRumRNStTFph2KB3YgmK
yS/ndv0RuNdBbSyj0WUJDMa5e9u7di1TM3S/bhSpM44ElAy6dV3O0yZsV6rh7Hba
dI3aphPT8NQbpJDDt5qXj+UhFHs9CWTif+GN2JjjDCoCP4gBf6NKMgSU3RJmYdag
awDKFZ3lXVeJn+g4lnI8uwLDF+7CYUtq48FFSj6jq29hJzbsUU5ipqbfifscssn+
zrXsgIGI3e5xGD/0u9yYBf0pgVUIX5lFQkCCw+pR9kBC2bC9cv8PHRsFc2ydjldT
SRZ/V33qMPIwiFCfwHLi4b3J4Fd1nJXob5oNgBumQHtzPnjZziSrdwkso2IjLHQJ
+Huyrh9cAmHrue7y47t9XmjjUdRz0KcfVcezdzx5xD4QLBWMFEEExGOMzYouqn0i
s2/7WQFo8heAuWGRkcXYiyczPPV47Mi3u5DMiPyshE3wrY7f6bf8aE6Kw03vGwvf
4aQaHEwupd/DAcs3ruDyEWZrg7BIrWzQPW56eOMAyp8Vco50yyQNjcHjApWkOv0g
E1YwsicBsZIJBbKZbUlDFH9FXtg+LcKxeLFZFOvX3lAwFN9BI1ibVZ/+GNJUEqmW
xuZ8ZO1u+BPXIkunYniEsC/1vw25nfK6ZdCObHkget8gMHjiUYADqCIAFwBFj3oO
1b/xzPOCPuJGwSJZQXCkpH29kYPvo21baZEM72swggouDUU2zN73Q3n8P4w4wWSK
/3/ndFldjETIQOdki6hCmc9DGQ/rK2uCABOZSCjqymMArUad9StOQKPaXIDw5hi9
/Vxqihrzb/4TZxbJE0hyxzezjy4VUw+LbIQy2qfDolVEF6uEd9hl7ZkxhaFakCEJ
RChhOSXQBhNt6YhPozzVU8bKfYfWFIoWvCDPExrFG1llnllGEKeN/wi5UCcd/MRA
loFjLo+2izJlnvUbLsY/dlvnKm/wBHSw17QzIK22ALbbOuECCqSSylVtwUamohRD
3BFusTr9XNBdeo1TooBzW4PtYpxvojJ3YcZ+V7twbBN8qRhy7HopTI3xqEmqnmT9
0ckA825U3Z3vxIxNrqqCrZPj03GCFulUtwhtTl7WHutW0j9xE3Y4QvDwllJoo+66
HLE9Uz4iX1XXsqZecZW+2aVvn7IzA3+K8QGwBKlnoetzfu2iYZHp92tUg/7ayu+E
RQogSNhUyo+zMh4Tc1IRLNyPGXijv5AB3X/ubRBQX2tDZ6pnHc9EoR9wN2R3Ch2H
TGyX+RxS4Q1nJO199u8Sx8FT8lHpTz8wQQlfO2lmxv7SF7QAaMcjN3t+eLOLOv3J
d7kz5yjKjMzPL2p0JMhM+0FUmVdBJPBUbEjhpIXNkbIDbgLWz6dIgNQccNEyy75+
Fq7zU1B0g/hg9cZ8DVFxGljQaVW+0oylPhJQugo3SKvKN1h/OZQYlE8JshHoByXQ
5Q36P/5lysGS3MbO2YRIZFqhhUa5onzKyXNNdCeU9lU4qL5gF3dUEEGYNVJbU7nP
EQl3guYz5289zoS/vPs2krwPm/fjYC0cvPwMP1seL5VpEHNAynMz/0fzsPsK6gJc
ov05Fcad/jjz2Qs0XtVe4xJJXcrDfEe9bDXUaMBliYxeesO1BujkWTuFBQTO9VX1
fxO1RRXhAjtp51eSZIcpFw0ut/lsOk9wWZS0Erw+aGpg5aq2ynrla5ZOn6Ld1IRW
UQCLT7ObWyPf9IcX+rqKKomvISQBdIDmMQhtgh/I+BYKIj+xaYwx/FPUn5L3cGNN
w1BQLcVuFFe2FvnkZAXrce9WSm19b1Fd4IyU4UK/rEmjHeQk7ecihQrQtSl/Bsbx
t+EnnvZcims8OoZC8TnlMZBdRodYLjS3nGzYlv+N7yzxFUE0jmpEIyBdCMwV5dmL
Tv/XnSbMwHn1NXwdD6PA16enqOv6orljNquivc9mHxo2kDIgioi+DDtagRwoB1sp
PHpAQ+pF2GdrXXNvp15hIPsFtwkJI07sgC9Gqt+XH851kPzFTg9vT7nG7KhrsKn7
52hEtUIrnQXUDbdsEziI6cYUGKnjaoGipDzY7ebcQGktA1Yw+eGOefArQa4eqovl
7pVqVTfjwy0W/p/5c0VcTpqdDOjMoOhQR5dZPd0ElpIVJXWLaf6OCGXbbvGZE6dP
r1H1veObzxPfUKBj4jiFdAuzpn/4b9/E5cm5QzHHFNWae8CUzB30nO4FDllDYvlz
9T6WbwUU0mninYv96k4bSDtkqjRiuMtislJmHcVpu8iH4JuDb/lXk9KwV6rXF0Fr
KHG5bA1M01iwHSiMjSICYsd/zZLT1olFasRCYYE1rI4yEbLBoS/NjGkmyrb6smYF
4m/R9Jj8A8dDnMb9srAOR3tYlmBmHb55kJdHCDeyH+CoU1oPpG2LR1crq86GnE/f
eOZCWoJfpHjK29BXLSqhXDOhRKSEN0pfwspc22YzR1B76+yUBBpNfAId9LBEunUQ
KyNY9OblqlNMewvPnOekk8c38jIwKKUpXQqWR/l4QlPgkAt6SpnQCLjK22WeoZGw
OSmqhLgMxfnGgmvCaSqcqhctk9L9MJxbfzX9SNyJWsuybNY/tZB+yYbviYysmEU4
lUaRm9auczDQIpR+r6V2KtdUHdKGUwwrtmSuFroRejDstzaNls2wjmjH+mjZ9YP7
XzyzvwfsNwF3O2taTH1de8QMJWG/RHHpQQQtS4ndoHlvC8w+Xvm792QI1EjC1/L8
0lhm+oJfuxKZs1SVvteD1oq0xAseu1baa3quM6TIvfbZudaH6MiJc77Ad5W7tDGV
sokpfQQhNdyAd5EBt+j4Mo4eB+IBMMm5mX7ung+0mEGiquwBHEDJB136ghYDMiDg
1k4VkmCY7N44LVm5Y/kSISKj7ZqKW2LeFiswntDEFE1fOSb8n72xah2bvZ8Y6wNP
WcHDy47v8g0bcTtcQR1HKF+N3e0B3dCbyRu2o8y/PkrN3eBfanwhLUvnqvLy6uYY
99qh2ycleQNQNSeCLs0FW9FF9+1TxzmnUDl3UVV4w/cW0t2pZkOGsl0+817jVohH
2pSdeiQWXTGvhnFWNoe6pFvVidJ6h60b31oinhye9sKBOyvoPmdQKNRFicxsPqxx
NjSVb9mXjFxmyLdWUQ1KFqBLCsgwpgKYNClI5HCu3l155cGG0pFOxEh8vECi03rm
OzRyzTKh3Jt/95Zn2PWsOCCpJp17TT2LesQDFlm4vL35TFeURcuDlOe1DLiJMFQo
NZE1UvVENzx4nW9fIfv9KnfsQvATpa7YlX7AxNIODpkkvWL3RiPyVhkukGJrY7IL
+Sp0/0rRHtDTcmfyWG1Fh6TVf14nGGoOrUEWURzRAZgZnsZCCU4Jto64znUW/1x5
JJNQGBF2idHCds6mUvzzHiUpJmZs7IVScCCa2I5o0WcR40wgLvOzL6IHgHUSFJY5
xQzTpFBXXBGs7PdcdDhAYxbicaO9AkOuiLwIirnrGSKV8BXpymDPVEZqTUmergnL
uIKoDp1DCKS6DDtQy9y5uIQAfn2o1QZruseoE8yoCDK5NMGoC8uFDXdqqhdydPom
8pqIVdRbdqFBJ8cyDLTxlK584SbiHDo7UtCFe9NG5v6J2qsyVxavCi5DrQBo5XHi
eD1Yvj0rlA/03LnGicm2aJeEBNP86lpH7BtgM9Tkh59r5RraN3g0BWTC41InLW+g
fzrAi5+LoQREahcWVzZMVt1uuObHtX/Z4+BWXtodchx8PKXaz+A7w6zvko/J4Qmu
hYu9BJI/b6XgoLFdDfTc73yZ1T2PBKzzyzYl5MXb4JkiRy2cpTZ9D+oU9KuUDeSS
oX8yYJtdjuc7Uzp0CrNx6BRkpjzLiPX73gwG5k+kylmIDoNZ1gwbPCaPcq9Dq1TR
B4k0v5AebpuCyPnVrKdtkGJEJR1YMMIy6bhavt9273VfNu4/rOs5nGG6c/cI2ykF
gJ9uCT75tiQXk+8zhZEGyqXGH57yTcwMtUsBFchz/3lztHFC3uynmzflbeMjlClI
cBp1Smx4Bf98NUHVhTprMVtCh1ZH+3imMLYeWCD/QujTTGOZRtI+467yM3rinGmC
ec6J+KCVycX94HvGzkQ6+i70MtgZpRJ6gOzx7OBnMcvTb5vlofAi1AfQInGoCS9w
O3soWX8av/bKamNOuKblBvKdu0adsHedIbZISlX6lzEkusBav28DaOuZHEyg7Sam
0aptcNbLxZk0vqmrxQHQkeeHYJbAU9+HR9lBoMyQeNPvMpzUK2VGAIwt6ZShGDga
0HTGM3XfLOcRg0QzmXmrQURj82tPD8R53oJczjRKQeytYert3MBnNJ92V2stKQ7k
618pKmEorBi1/2V6mWFN/hAUcqiVtycG+d4Ln/CBSCgOFTkZPiNuBeo8ZmmbM3A5
3TI9wXtOc2laoLON7fNa1lDm9tz26vouV3PEHmAKZFleRLFKBsERATUyhz3mdFIC
EudKDuyRYDpsj3zzfcMX6zU6yl/mafDLbfaCch7GhxWNn39+Q0prsjNERTxK1zMe
ojcJLhvKmqMAeNg4fXJ0fLPuM6Nd/xBTOkya4EKRBWcF7guHp2UTRq07kAYJaJx5
doTT4sherWaVA5XU7MkWLjkTzxDxqaxfSCzSdQGxUJWadLx7mCFgHknlSzCaVV/h
MDW/CoDnv7mk6yFoYAJEikNob+XMSi4YIkY+UOqmmIdk4oFxMUEQ76ZQ+VPM9iCe
THm/HKHlRXTxOP0TGHy0lXRn1DeYF+1XxzkpV5nwkeRIbjNM2ioZ51jTJvaeh4Vr
FMLb8dj/At6SGplNdd1MEGoJjNCuyleeyduQj1LxAMp+DddiUjN6ZJKAnehImHvt
laWmzXx3zErtubzwrzvcjWZYnMEQoYeETT8trWSNn71/yfMy/E8kc6tvbDdrwAVz
Sf3ZuEdFqlxKVJQGx4TRMZKwsI/O23uSj/DtcsKlKslj8wcfd3ourM6WvXn62LyE
NbF6s4kJqLuZU0mB3oDZGUw0zjGg/jK1y0AkWTIUeLGUlpRlUJkbmUC6/l2FZELU
SKbCgUiaMMzZYpNs2tucc1IFSL1dtjQhPC1iVFl/rko/I2GrI6g5r7PjtoIPlswX
vHImsZZffrZVhzFSptPIBOw1cefQFrcvCVDPNsYf0MQ+h+wotS3cLlE/+r+xUlBl
st9vUrNarhOwruHXLBQhKdsiH7LWGxwI85JcsIFJiB+KFakcdFtetSkO6qg3NDvx
YXId0sfGb1SBIRM5K7oKXaq4FUOFOzM9Zf+etsBb9NSlUQ2iFSyKyoLyzPHbQMwO
1i6/i3Vaz9qWcxYsLIHNwt0S/IhB7Ez//r1UXnPPNBtVDETSBZ+9aSudKRjnPMVQ
cBZ0/K5gXZcKwZLOWaK3H7T/SyuT066Ts59LcAWChdlcpQVWmulD1Mk8qYkXE6Tj
fKANfECYLTX9Os5Frfn8hmZXb/RI27sfBb2H0WjJA4AVIgdjwaWPHmTw7oykCL+/
YLwBeFvB3bg6kgHJxR2evuZMnb1r6D8XffcSFIx/DIT1WxUUYqsOA9Ed8Q4j8kMd
4TcWhzQftVXiFARmMJlmgzj4AgwSp/0HhKXXjXQsOZY2qNZAi2Dx0qU0wk3WoOhv
27zfOmPzyXi+RVN2jHFHFEujbpsli3n2DxqwpQQXqWSO6cm0978z0+4/xEklBSQc
owenDoWtnYBryOz00JbJJ7rkSUop/3yrpuouuM8u1ubqh4UFB4HA90hUlFHFo9oo
mCbDKiiG1RdH3BpAAcMcmcegCQZjx9BAnq0YyZQJ42B+yat7QTLZVFPiEAjwSL1w
m4KLU07j7ebHAfBDEuvESiTh47xZr4h7jfgtkHqHUwGUuXsenNX+gt5oocmquSl7
Jux3wvZIryYIdGp5TC8mcEgCuMSPoxlYS28fkAFkg4ge1n1sG/T3ScmoXqofnD/A
4jXiTEjU0VUstXtNpuk6MZ3KtBPZT569C0yn1IVsZbKEGlOSCqTljMpHELR74mu3
uS3KM7WUgg9c7PenPYJMUnHDr9YvCY5FKeAo+HMVDyI+lXjadbtDg4TmWx3/MiAw
5jv6fquAoqs06hYrlYPCEp+dkA8YRdrXN5q5TEytbWkE+vPhdXCG49lpCPvSpIKA
j1JTjAN7cGk4garDRalg2JaTb6IpYzZxWYqjSqjVbkZthNyDA0XwQQ+altgPlnjh
Y1XO6wI0BpHJJ9BigiPB/llXcqUtdISc1WZf51npWv+ekvIUIUHJGb5YK6CYgeX3
2J9SreWwLT27vgHqpM+mD15TDnL6QIv3VsNfhjag24244XE9h+Ij0iKihFBsbNex
6RRMQb7+pHxDvNP8JwQ3yboe7DOTsXJJnuQA86P44cBnUHmQn4zgGdgmfeag2vNO
8UlaaaqIk0W1gXVrJsXq/jDVO/hATKGSMWHu7PY8p0ngO4FgBlCBAxAx+tfA5yhQ
W+oL/86Xrx6XLrDwbNVKeQBNh/kVxYMbtEn262m5gDfHWXzkezutIIuSGTxUe/K0
F9nbNBqpZqPscZEQK1AI1X55c1JoBHcNI+tjm2wJBjK2VzoE5EtUDTjeAhKrN9Uf
YXn7pQFCpzJql5sMp/efqBPCSBp3ag/iO7dV9AUeJ3vI9XJx1IeDdKVo/yx8dGEs
fuW/F2EQ4hOQN6iLf+Hvj1CKZdTPVwGmJeLKJQ7t/Girg5sVuNZMxWOfQil/lNQx
p2nNBpIID+O81jYZraWc70WiUI2vQ4dzjH/3UxeVbx8V9vOO/gnfN3vfB32Hqdnz
X1qp9Kxb9z5DViQgIKOFJ7vVuWMzosuKx1qFyUbaDU4sNqNukXdLr4SqSIgixhr0
V9W5gG2OJm1JtmVaxRkiVCz6UITQoJDhGHDji6EQQZ6NzGeirCRwKYcl6sn3DLHM
aMiAqFQMYhPCWNZvTdfJS304mQ5fxd37I6NHjw7UxacSnecccTcIIhfCNPQOmZJ+
xzxr++PJPOdAprHOjcHhEqXVl4PZ75uCw9MwVhlCGC26EQVCF7vU+Jsx/XCtOAJM
+I4yISoXgIpb0fv3jHVQB8wgbF4me0d1mCKlktKCV5+sdX09ICCDUUoutyBCTL7m
QkpIm7tWuQQ5jcYWFyqNO2je9H8aRZrORooPbs/N0YeyFgQ0dOxPcLmGf8gcAqDu
GOImExKLlvyfx4tIZ2GvQX/XWpBp1lB61qhx0bfwOzvOxQhThvYOi/HoMDlib5mZ
yndTPmTx/uMQ6cSOKB154Cxd/XAF2Y5l4VBA5nQCLk5lU5S92zJjax/i+SHgMLgi
8WgxRZheT/EwJe/RUj2FG3XTpnzzbFg8xyqxeEirHYE6rMNCxEDcjSFnoy9OSVdB
KM7oBjwshEOjG9zdyGtd+CHsc41BJianTYedJLPH09kvNn3URo6G2q0pcFl8uWEP
6L6PSlh4CrQ4iPx6iexp3XFQ8T5BNfGNMq8fpEbLxzcvr00Z8EWQtjtS4Ua7B4wn
OWoB4M8MWkbW0pxLXSSdEV0yc/q8V14H3m+gVi+89GEeQQy8HqU7pXzujcQWMqWa
yCO4udc0txAeA8g8aLJ9bV5lGTIdsz7KJS2hRQI1yehpc7W74uFhkgE8cwlHuxRB
4Mi2zH8uToj3xG5/pBq2EB6LJ4dyCYUpKoFarD8yUGbsxyC6imDg2UBycHrFXZlr
izTm0cHKzP4AOed6cP4GvWzCHr3EGd7rikwUbSolOw+iTlUubfsAg1Fod9nayJZk
bPgl/lFTfHCLKNqX72yW6NYQDUgrOvJeKnvihGpAPHG2wS58yUn8oDZxkomH9Wcd
iImCQUYxjtrFgZxffo/KQu20Yp1hWJ91mkeD4pA0tjfhF+aPdNOf0QPIxFvxDptK
U9aEI8gYBw6MhPYc6yux9iWH+/zl45EeRv6Ngazg92x3jCEtDskXbv7e9+L5TYD0
7Bq6Rx9/LhLgbVuZP0g2HGmL/bwisDTL7SNl1n6U9Zid0NHU1MJpsyJ6zw5pHL17
yC0tPbshexChGWt3yNqCjB+vJfvPfIxo9StkKJyjU40d7z+O5SAOtzAbtUtk3s9w
ipS7IHx0gHC0ByPqKJIaNRUJMdQJb3tlzrd0+ShxJwn/WNQnSlJIDPV0XQNyRt7E
sPsSgDS2pp+MTkS94zpjwn0m2Wh83f8JITuC2/paE2YT9PaBM+BM8f0aqxBAIyYM
W2g4VrjPp98lVJXDQk363nWCjTR/lmDKM73c9xOYNdNsoy/K+uucUejMHygBtLCx
CYm6PXUV/mkvT4smJR2n8sz8EG624YZsSMrpfF9w7Y3UOBL2EhSGnEzdJv595Eiv
HfAWF1sMMEkaHM7bs0cX7IApQDiEDf0lJzj416HXA9CaCjvXempPYXj4M0wLkVkV
y7XJ83BkTMrjpAlrHKNBse++Qru5fcPRzoTQ4o2xwzTjIlWvxOAXyDZrbB4nxrCL
z5R9w70kS24atx5k719/rSj/iZp1Sp9VNQAvPBFbSFofQA4TjWtbVuFDMEiq/CNH
i/BsnE4VpFrZDeSsQdZm6YjDCZmV4IdFU248hvRqLqwDP6kt+KjSEA5mHMi4WCvw
GWLLdNOZs/fhxOSM/iKtRm83tFWe5gENPYlbb1IRy8iPYKnqSN5pfXqVjJ5wsAHR
+saTAFpb9kf5gxKMm5QH6/i/kZV1Ebmjw83mBst0aAV6LshAhiqtFGNjNAf5eiYA
NxwFm8IzITN5WMSyyHAlR51FO5ovx33ypT3tvLN0zW7AxyqxFzJ1oe4RjMmcYK0Z
O9R4UFuBOZtHLDXkI+1M+6nPb/H9QWTFDQG6Hms/hAKtP/fzt7DDIfNISu8TfJWs
hNGG4tNdDVqWapjdgANA7qdlLi/lrOWD5IS7QmxHcKOUIrHPpgXdr04ApxAtiN5w
R+XY4vC+20WN/mO+qZjd7d+D43dnNtth4M/gt90/iBtHHg8IWRWbthstqVLzd4VQ
H0p5tcW4oF12ll7VcLlC0R7uWivZ4XdKN+KKtZ9Qjgeyrjg5b+hC/CkW2PIEd+LT
ZRUJdCcw8f72aLUIjbn9U4tlVXWlaM9h0kls4iB2CBuu9fG/xy00RdjBMMIcCd+U
VY3FFoOFLvHxJcWZXIwIFxu/C0LIOfpHXY7CC3G+5zSbyauq/IK8ZbLJsD2NGnUN
ArX0hxJfUBnQ25Wz5enxFQgVUDXad9+/DdFVD0cqgI5+B5o6dy9gWsuVCBhQ6bOV
Oe+RRxOfIuz9kvCeDzdQQHAjoRT+5rxZGR3+aBj3Z+LZit3RwVUm/guqYmEGs/M1
VwR7fODtixb+JQgpAPKENBPCbHEkk0u3JhoPmKdaWd5i78A2lK1APYgxKVYQJdSD
w94j8xYD62obDglnGpD5qeiBU7uHKhXLkw9kZpypKbeoG9PD+2uJhOCDIfvE19z/
nvww36a5J68K1n0OSiuhwVcKqZO0+uXWsr4AC+KOkR8dN+3HLWFOGx0JZyw7VL2t
wYc5yHri40svHGBgZzESm87ddz8nbiyjd3c5My3OOHzpxpueAP9EiKvwrvKxMVAk
VTRajBsxX2LoR2GhrYxE8mFcqD7bU0ojWvHl4bkDNBoii3iTHXu/6su2AdSeNi2v
6LFEUbiiCc+ageY7oOHf2Q/z/LCiEMQMYaTPSDtOhBR0M9OtmadJthlN73w/O4vS
X8FtHPPn0o1Vxs1Wl9Dq9GTsclAcSM1C0iEMTB7sKqZQtQUhoKg2gdMKhWdnZuqu
J6fTQq3fHsFCbaTSDjVdiIMg7ROM8h0KD0m5kDgjWz5zA/S2Ki++myOd7QG/JqlQ
lzTFMY39sxXy7iSjqeXaWoQNkymTJE5Iywj77wexPU4+96Kz5qHCQ+7H2ctnvfwG
0bA1u5fpbwQLIURiVSLb24F1p6fuNb1U7EWCdtpHwAo58CdNKyXvC1V+QtE7zNmC
UebmwRBMjA7H/DHky6vlPuOVlyBcAgdamPCQgnJr4ujzIkBeTWOT+2kzGWgWBj9u
5rwj/7Zh3CXRZmnQUYiRaAuC4d/jWTHMehJOuyLPbauIUnrqgRmK7p0PcZWZ7U+k
H7bRZr7nTxpqCp8kaAP0bYdnV9P+Dghksch6+6nfNhC99Rgy1MkWuIuf1p6wz55a
AIHmV3fLVXjnOFlbs/MmivYVP+U4MivUVTTYhjoauhXzixCTe9Fg+YRvFsYRCEUp
9yBAtLtlt98eDgbJXQZKLHyKFCbr7nFQrZjgKCqFh2yVdwptJYBcRE8YfbAYQztp
DXhW/AsuVU3TwUOQfM4V5uOacbMDNBYmF5FlP53pBeObf3wXFcisychibUKOLB/P
5JLwSH1TO/Plcuo5vu2bXNA6eWjYdu1pi3BIjqREixWwXS++zqUepApo5xc/LXNL
wpi1BkaqLfz4v+NIgioTQeZdUpDaXQIubRM0gDJuPIJEXUtTcXkfsMlaabk/GE4R
NLJOtfik9RLFCW9Ru98RXflORHDANNJdN/o8oXHRnCEboCzYaWvYLmL2C4IZEwti
Wm8n+EJceOcqIf6Mn4/kk0o0r3wS09NgO1QZ+lsAisWrbcLFYRMB9BWu0tMwiPKw
FBBH/v/lsj2tOwZ0hcQcafCREtt9GOsRwQZEfuYU7OtALusZqtw7L4GokNxazPmw
jppKPYuQjSGnGcqTrHg7+CVBd+NKir8buzKjxotKf8str7RVCX8JjA9uMo2H/Cws
NGDJsMf9wEO05A57kDkj2AbLVWqUAieUPZ1mcucJARzCsALAUKrlADKJycCmacj9
d4r4lV8D4/OVXV1USBchwCGLerhgymVbJxshUXt/y24Z1NjlG8ms3hpQdOR5XbXc
LhC+XSq3b1lV3BEBpcYrTUKhezBUx/i8UGdrcGIcMpOjf1yH4/SlHJyLfZ/l8z30
v8Z5HXU7T51Sxs8BNwZr1J/tHmZYCmFWr1MTyqAHOI/XjV1fXknkRC//FITbxRyo
uKE6v4cb5phQ5XwmQHz909v4gLvjThLXZY1nRb/j4J0aRbzTmf80aqZ3bJubGUIF
P3TNoKUjk8x2YXc/L33ZDuBce7wH5Wk9eDPL2p/JjCePaj7OvHDEqq4bLtb2arK9
+0UHnJGvEjuQA1bdspF2FOUSSd52t5bfFA99JhmZm3/148vqKybaAmfjbGS/3wE5
iCc6/licpb56Xrq24tgTtEY7HwvKOW3viVUC3PARVK6YvuFVDq7HZ/vr7JQanOqH
B1nNavIbfBWKPp/1DzdIBvY/ZV499g+tGBfgoaq3qXPHxk0hXuAO6ZuZeIvg0RLG
VmR3zEnU9bsemYJfqUOVMB6t3EUZh6rN8AN6pnGBUuzIR0DD+EBCkdTW+u8RvWRc
qh2XWvM3wPgE86xBU+2p/9zt7jvkOEnYMeUd8hajOX4ARuBqOttV2nZSHWZQ0aBp
iZmVE+zeuYKVjcUPGbMv3sGyCmApjSB0Vu13mhxdJPgd02NhgEnKPPXcxO1zMf8Z
ZnQRxgLavK13b2lPmgutCc2V6sAmrb5CqMSaXAd4LCIYlIXnzms+uzOa8V1vQztP
Z/gASBlBRBOcRwj9mjtl2JDNqhGW1qlHcrizV2uA6aNDHSa1FutiOROvECPxGUWL
/J4TjiZdZSqdhCb7v3q6/ITRrDRjw+cd3FfrMA5f6T8HjP2gtHkRDFgseco2MhSO
/mqW22Bd7pDiXXceZRs68BImVlm+hhnR98Kbc6fnRnXbmdgqYFG6SS3VpOGzbdc2
u37WbPCCoNAsE3fbow2le9exf+7s4DBR9xMW4c0Ko3ZJij3mM9vEkx2bvAqkn492
Zo3Kb9MklkX01b20B7pbB7W49h7riWLnLYGK4c9ipaU8J1vyl4GxX0ak7sjkCHoa
emOLFT2qGUB5uauGUPYS1mD4n6iVoVD6YIjNQ5dRPg0l6vCUWkvzgyJkdgG6eB0c
uDYFIB0/pWxEnCniXT1fYd076FzUyiuyRckfWxcDnNuowVD5slQIIjM7w7M/ztaQ
NEzxb0mJRm1lcG3o7D+BcHY3kvOS+4yaEMsyIBuCVBTZlmWdmHwS/AiCQvt7NH2u
RSEiGedURhzMS5DDsYoM6avrVUcqLsKiSTBveI/rXveQ7SEb1OmpP+ZP049BS3SZ
mRoczawdvUQNcB0oVhVk/KrROgQyV3TGagx9VDuyxYTHFzTvDtfsWKaarz/bn37S
/YYT7o81vBpaOnVClDtSHcSr4ax0Yy4mJysKqgquAGk7n3io3Z59i1GKyUpMh9++
xi5or28PTJ4GDzSM0QXriRpxYUv0WAumI+JH1JAb5AMLzPj8KLI8k4UWP/iyolXQ
Y/e4QA6iUPTGyg9DakAzCAdGmRAHe0O+TcD036sx2iHCvesrCoSXVKZSGN+JxS+e
K+a4o69TCahBZLdmjIZSI7aHyCQSO/eM+1cL9wx4xuddXSG2PFBiYALaYAtws7A0
mdO9RXbt9B7DFFI7y6G727W20jyWwZrcobzS0IclOszQapb2zpswm9xk8k8aoZpG
McbU4BfO8y2uG/CsITTTply61kBiARHWm4P5lx4Zgwfw++qMTvj5+BA6LLr3pZX+
otoQH1hlAVzpy5uAtZ3cMKHgHRcp/zDRdt7vV/DxNIYQdCvaFgzE5+JiKepILutB
6hEPMq0ul+cOKVfgDIhpuJyJAgoQhgECYemwamV3iHtuDVjKY7fpaKxmsAQb8+wh
letHgg5xMkXyc5FGCXIPu6LF+IjM5WBUoZobj3jgYQjddscYZPVo2/rYvpW9woGx
gy4+N24yHG7rYcmypnWdECksldFhPKC5vyeMFERouUqG4tH91Qfv+x2Tn12Kbjr9
dCalyg4GJoYuk8ROfpeHwnEyDOK5bpFMX7yeSktLPJSKMTkHAUK+UJyoZRRtxp8+
clfW8xUW58S/f4VJ6vayM/HxpEQp9/3iE3W7YWeRQHY85bV35RRxdLknnD6DsyQ0
0ZpXeTGj3up6STTdRNxqWOgvOBemGBGLdvJJpYqW0WMtHMNZHeFAFGJM3S/facpC
IlL6wgFymUMGU0CIIXSHz8M+r5NWNeH6pUXFMQsALgqhwutNTd6PwVyOIwz7QA2Z
Ew4J69Rpd1pS2pEn3BmujiiQpOu7E3shFTpzNH8AlL3BRPiI7hV5YQHrCHtLiPgB
hIIthZGCXBVTmyNiChudVbWQy4wGLyiClDkkRNa0GLDxJtXKRoq5b3SPPg6xSiA6
8+pOs/eC+RFKtJRLu2vEOPi0J23H6B1gz3kAVAyWfqANWqDrT43RJF5LBNfqxa0a
PaP+qC73XmrpFimNRaY7KVl2QTce1LcdURj+xUHBZ1PlMkDhFrhFuDQ3PflkkFj8
TSX1m48MfMYS/aYk5FTS6aUyatLYtR6GOoIs846s+qKOhUB5gkojhV5+HQt8dKPv
RK/S0512dUCqL2SgA9qPknRp4B9pl8ivYtBuiz0mI2gQrfyl8hFgcAUIryObWs29
Ro/0hEzyLSXq6eIC3OOPxTUjfCBQBcHBzwsdHH0jWQr8xgKc5ZSaOgackOzV8jU+
SGAmQpGRy+EXX0fAGfwpT1wGYLTo/JORRjSA3y4+sjaP3ghwm3UlQ20KgWlPsId+
ZUjxQW+DWr84FkEkA19+jaDAnWhcviYPdFPIaBJWGJ4rQtNJlHmUxrw572mXCVt3
nvsdaPzktAgu+uqSQ5A+8N/qFtkalLr7jv2anGHVrbDN9epUyUgymSApN5GcAEZn
0PrPlfbFKT8vpI80OsUrKGZT6PZBBYbYpZZzZZnHwWbCQuvNpH8ckAgVx1TRxayO
RE8GEaWx99qFbS99oW5Qh1cU5BXxOw54WFd8cw7mG6Z6CpXJ+R/ub7Nuu0IH+svM
7RrR1jy/t5DsebxAseoAhkktHeZqZV6HGLelqgHviy0Z80ePinLz/ZXOHKb27/nQ
Vd0dNWaZVGd9IFkctZqHY8vZz8K0xdymnLoaDlDE06U/PuiHCB0PycgafHYueqhW
L4ZoEzU1AxpJy2sc6Y79ezPUoEOu5pP38mHL0ydVUUuRyNTfYAkRN2a3ITKOK2M0
jN1bFoe3SKjroXppWSuK/WMAm40bUA4AunYVjjYtGA+JIK/mTckLRT4+5XgbIJtL
PeYcQPTNYePIU4bSZyS5Uit6sLBJV8KeD+qotguziY5jTnQgU+51eNMAayChHu39
jSrzEX9Rk0SwB1oTXs2KifEhrnPXvyig6jBnfme0KZmHpfyTue3qM8CGt0sqR3nV
7pwOfiVdZ/qCdNXiIk4tTDaxUvUrgZbcEJKhcIHbVkDO0SKfDL6MvGvuT3C9dvpU
8DWgPf4USAxCzXeMQlLdJdwAguzcU36naxXDn+NVq9PcaJS1ZCj/otP/jBW5XTwi
ie5YEHDQMJ+WiCBe18PMXHJoOoanQnRLkBeT4X+oGOoQGZjsa41Xm0wJuYOJ1VH/
1zw36No8mUJKwXp+tAcsIqCV4uZkDuLzfS/s+fLUWV++8qn3z0N0qhB7CV91mqyP
iGPmoDvPs2q66sLmbLC2waVY/2lfclzDJiPHGjtUIZoDWXyYrD66UczF0gA6DmwW
bplRXZjnGYErsUQjZHCvSpeWM4/fNxUG6ajnENgoCCOw9ZkGNqbsWCFELosqO4GD
DDL4SEi5nsiZ/YSrmS+buNsVjelocExQdnLzO4Cl+f6fZwLlc08kLWMTHX4cFFwc
kdK4CYgA5OMfyywS2crbrRIiuOcnChen2Xn6RzQbEAv6aaAT/J8XyqtvFxWZPS3j
a0+cr8vZhqKSw7NSm1AW/il9vJp7j1iC4maOkzNbMpCWfgCI0PERwZY46qxOnTis
bkr9zKtNkFmKT8A+bkxJY9bU2pRECSOBsndDM5k/S7sK4ybSefsSLJ+kzvGUmEZu
EaVk4jOAKydHBD5GtHnkG0/je9laGwJTg/IOwiDiO6t1aEOHxTJYAAb3bodNlYuS
H+Xaf/ZzNhKMQieZxDGQs/o5ImQ8KLsdiOqJ0MeDtTCXZxdLy9JmGBPBlcUdKIRH
rEdOTWO4LG5CeBygApWOycdHckWbdJTGPxEzEW6n6+kVspqH1KxJXrHva4jI5e7x
Bw0wd7kmDWXB1RbNSuxdi9LleVNn/BH4gtFFdUkHdzoPFGhfiMCNOcWJf/Kao2yl
FkgnBAYxfYXYI5MuD0cLnQdBaP5sUW1icraDdXw07HrIaUrCeGAnZUq5eK3ZqCZc
VuOJ61zUMxJA3glLl1n/sBHIXzfGztxSoYZmrl7ZjRLDxAzmNu1rbAcJOTj8IXcs
NUMl/YI2eCI5xH68ZHtTA9/dtM00xAErbanewjMjVVaA6R+MS5u2RXIF1ZTJUPHq
0zMNZIrt3scpXLgREvdJEyEAg8r8er01s2FqWkfocoAZxZ/O6bp8Yj1kXPGZqX9A
vTNej0psp9C4pdpR8FqC/wTcwzN7Jw/twrhTjdlyz9a7rn+icPWf9eANt3Xp0hjE
2dzd6VryjVChH6eDWIn7SqUFwtwD5tZPQOPhkOQK0Kxq631DdlmXMBmZtEevOwf0
dMYFBJCL8U47opJgi607ore4roDzL0jI6jkSG/hXXEqq7Jhg1A3WpDQ8g04lOaDB
Y0CbnCBPCmKIaMPYLjS+7D8E/luYqDiRIyFTsdCK+3j0c9YTXFqKZprinVHg4wkl
r6IR2hfimj26CmX7yuDFIi7Qo9BSoKIgOZ/DYG7zwowVd+yOm/IDg7fkhSOyJqmR
Kv/kqDS/f2y1diysrDdCWFWuJdqN0562a2ZGTyhWbnmnBw/BViwUS9OhNtGEthNj
1leS6WZZdyfez3S89bdAY44Ds+saScQhES/zcmiX0K/17rP8N/kSD190vJ4Uc70i
cpzRitjZpn2k2yqyeujlzVdISul7EfnzbgjcmhkxT2xBzh8RDyde7Sm6NwzMgGd3
8mcyOUq1mADkO371ePba6sv1hju/wuCgM6VF/xR+9bhOgi8Yi0AryqLDxObfRWCt
UJbX2EwNuetTIsBJZIFxVRxpmWnC/ZsQ3W5xiTbUPh5TzBUrafWXbDkiCWWkELLj
DP1pcHVcmhskFhTDdbqs6emnVzLwhsA1QsMJoqNMqOxSLXP/YVlT9MKKO7WFnfIn
53WGnTWHtOFjgkdqftjaoI5kUiwhh/lmDIHna8YHkUrZmDO2AtieI8WFb0EG+I5Q
qX+TO9uJaxRjyreqUwKrEcisrjkhcWLFA60gqQbt+0b4U8RbOi7UerrwY0mxrJpC
vMhtb7d6RWE9DKkhG1AgzLV+ORAu8XB0KmKj2W2YTDIKlE/lhOC7KirpEKYx9pMU
6E+tkk6NOVa/0MelYI1me6Wh5mUA/KOxqgxe5iW2/nBlHmoXzlnLnarPPRDjqxeE
eahthCxBjKaziSGAxWO3ZGkq0qkrIjCbKZg0wmpdYBoSYp3xAaZjCY7QdH1LE1va
UAXthLN+Ey3Wo417+T5si64bknjg1XY806msqncFhWKzMP0LUmzOpWxU/K3/rIo7
3b6+sFGOfY3iY+v7n8o1nRzqASY3AgJTsdiT8c3Ut5nNsUDANQLyAfLxeLECwQ7F
MJnW0v4iLdP7aXhc8wZ8IG+NuiMRcyoS3SFUgIyLLPLNT/bUAUL8nU785/WDyZym
dVuihPeCL8zHV4v3fiuxQvvtVNRz1lU8ltvX+Yr3BrtjFGFoBXUBr265Wa4DQmci
kxC5L9TkEGYceZSQX26GQyHCHSBJM0AzkF1FNnvvRN8/h/LPRIyqtFidH9aGIdRL
TlQrM+12dCJifyLljOlRO+yV6qSJISm5U4G9wIScP1CFHFQPRnN1tkbKD4H/GfD4
qEjSG5KV+JLMCwaM9ob1trAiGiZhHDIXy3CTtlqWh108rFxeOQOhEI4oiJMmDE77
emiltA6wXF3NSKQgozOCUDaDthiBrZppooeiOVw7i1eLeh3kPVV/MeLYUShnxisu
hG8IBTIFrxapzetVzcx/w83rLhFrZYbBIkstD7tsafdbWGQzLFylEIOGLW/kPGpf
SCaJKjEG3FprtriVgWKDyomDIq0aWGohnjBdigwDE9XKYjStSTFeD3N47M2yvKCe
P5iOziqKp78rzWuALJQcsBw2VBvuZ0j/KlTgSGIc9o4w3DxV2GbARxommQSgm9FX
JGy2uHjd2R/yBF/PIooyQiYPVwlDg0g0CXRnA9WIYhukAI1JUHfB8xsajpnIhINh
dFgPRDL/QStT8Kn3klDSy2LIfi9DL+hfzkLTD7Mv4i+F3xWXtkENkYeU//nwoE3V
i7OQyaXAkB+4paSMKMwnhtANCOTkRfIDXZ7jwRSmagOfcR/tIKZMa5/UXxEbv6Fl
Yx38wPkPZ5mfCO6UJMbgukziHCMxMiWtldRqQBpH3AEMNm3PHceQGj7OzqwT4buO
X5o+lHgF4YykYiETrMGlE1B5SxknoemmPi2xRFWZNbvy63M6EUvSWddwK8r4svfp
CUZ5Y03oLEx4FycYSC6VD4yQqaIBEdMep0tcEV8O6PSRoMBfvVWC7n8tsnU/c22w
qobf7V/rxYEl85gHBS4nbFMT2PxIGQ8mp21d1NijzjMFns6mGNyNOGAj84Wy659m
Xy0WygEJLnBoOPMY1luR3cJNzXwVLGh/9l7rI6AWJtNbA88mAGrSU5pknM96ivgm
42trmxmc87Nb8MrdwkVlLR7s4TEZtJry1xxZmy0k5+ArJyIkMha4ch6rRHA1VICz
5FO1IfZeQv+LslbPRI3UhAGNrZdQFR97fdnOViJE2fAcsxyoqqP99XnnTUx9SebL
neKy+of+oBWUSIj3UFheygG+V+LcomzguUTnD+5C/nGN5vSqleZrRxgZ+A1HD4TZ
nl3yTWLLANmHDiiflR0QU2SNrBCq6VtvY0H6NpBt7K3p6kuMFgV1Ra7aYsCwraFD
mTx7jlPykibCBlWS5V9sFUiOkRoJs+Wt58Z22BX/OD7eQ9EHzvxKIR90ZEGlOtsk
gDCjKH1fHbvpclcvVSWwKoBh95YwAlrsEAlngnGCtN5vT4bXo9JwxlCMNKwpQYXQ
f+mcIRD4v9xPXz0J/jh01/vv/ePRxd+2JZQH5Nm1dXb0E6PulD/7IwFHuFwkuBwx
ErdSLINrkTlq3LhI75lknA9aDwoE5SGHouJZt8KvjWt4oRfQvbNwX7oW7/bs4JGc
xz1sDLgmW+qsH2nROtWpNRVW80McexK9wQIFa8aD5r9qfXVg7KhxTX37l2LhpRhN
DScEkEC29bXHlvtVOuUadFS29+r3WztoZAkqU3H+ekFjKZnnw6OWK3i3ib3knIeM
8VtY4VoE+o075hkNIUV/huOHbgVRT2HDVLQd0+w3ya5xlVi+a3UDv16mSCMLoGsY
+uNFWA4gZv/SZV/m5f5Z1n2pztWm499podrw9aMilgWlza33zeOqCjMrnGQruqcN
aZGw3j1vNA6mKxZ/hzRYAVwuAJa+CWPNeHrCUzzclfK98tW4PdiyXD0TjWRrd5zP
EcedkvITrWrv9gnlzUnv7r6HfFUSbYdHwuxxOn8uDTirSupGSRNXGhDbhD7iiKev
QwjrHKi0gKNnCyORuub83eiDAwOj/VjTIuOCY3negzjmwY2oeibpHd0naHHpH0lS
0PWg5Zsr34zaHXS7arVScRQ986jAfPnVqaX5/Sb9DEYLHa/KFyHSaJi03KuLZjyu
nYbmDIKnPzloeM8ormwfFrRvE0NXVI9g41SZsIKTHU8itZJxDYfeDB9pI9E4tk34
K6OznY/MxHYQtlpvzPJvWaxtRhnRxfw8MS8LgkJ14BkDIb7tqfG9op+txxdEeXGu
Per+GIH1GoDKAjXtKqoZTp6en3vSWHYRqIKGmCnXPpbyWllqEjAMvdlEd8vFDllY
48x+lddaNMUG3ACO/O920KnUOlimO8Ew6Wlqz/DgPw9AcZsGGLutk/1Rr3QKKRZ/
yTYQ97d4FOzwSZmmoeCyQWHA6X930c6S3D7uuONsvDuDGWk8hFDo2KF0mQAo58sU
OQBMPzCxXKMurTl06KpOvB+LXHKeJTyJvyt1IP30iy/z8IALGF94m1HpWZsTO9PG
1+tgvjLkCEeVZgGHKlQtroLhbHvhQjJVY5HSeeoIBJVGOMuSyYtSlOMNnDTrZViy
qUAEGaNRiTQuuMmnIVwvW562OckUJuKATdeAb0SZVzFreX5cx/PaUC34oq4c4Smd
eClBerJ0LYkS6WDDirz7rMQQ/tsLbEfqD8GisTVv5F7QoQqsuJvzkDEomeBu9pHE
3CsVjwHO11WgWD9WOIWdzoQ46TR7Q158K8Q5Rqo2TieQfMkYNsq9WWZETrp8TEuQ
3prv0aqlrhtrZ345Z1+I8MFs34K25Ply9Y4/FLnxf7yipG4NPLdfWmFl1WkDdnWl
dvyrqKhY9IWol+SsIkEx4meRKRdq1/Jrmr/hi4Jo9FgiFbzvqqp2z7OhqdTrEd0x
0q4dyzbcDn9FKwX3xdYwK2U4pmSlIZmKW7Hgvv/l5DAvX9SiiXLK+VRRsxwLVNJO
KO36Cg0GTSoS6bcyY2Ay6fp/ptjdorN/rserweh8018+m7w8rPdI/xt5Cye3OXuH
YWj+YnDuK5qJA9tjmz7npc9mYaPOwUn488uTy8C9mXUfw4JnF9cQIxncgq8IUGyz
7+by6gFLh0sr7q7+8+uejdqBriyOZe0G4N/GFoAgIp+9Boq0TjX/QYn1vRl0H90J
FBXuidLB/l8cWSE5svDvo4F8xIHuRSM0EwWMXrg9QDMHh3DILtYfDJpuH0YN8O/c
Cv/9OeQB74r6/bgr6eNQUv58rgHMup6P3/7wBF98lso6skbfkWU+DZc8aPE8rpR6
OiPtohcsJ4VJEJfnFDNTAzm9AsnsqgmMWrhM2QhU59W5ZbD9RGC/lxc0aJ3ZflzN
7L3PEYaUAg/070N4Ph4DFTRGyBIJjv+kyZTMvpwTqywTIxsS9sm8C1xAf3hnd1F1
WzcwkICIodWrp8vyD8YzKr6BbZlnLJpyZ+i3Bob5izs5wiR9jzRyGF/zb3Ky71RB
AigfamSMwN6MwpPkyWEWKAvt/guahm3ljLY/xBZeJN2k70aH4J95je/qELWSfc8L
6GDUynTt8MSXpepGlKwabvjjHOgrg+j/JWURxvX5mheoRspUHM7LGr9hFh6N1m1R
fUJuDOpb7l74rlXd45FxmZl6Xyawn46FEFu1vjWn0VAP0WCNInCBt8KbLAUkKhva
7tLNswlDSWl8jdpJLa4DDe3nf9qTg9DzU9Phk/dJoo/lQ7Zxk6MIEi4oYsoApyc1
xL1tzEO18b2cb5c7nYO7vETnf7TfAdEBCQ+VmwgTB1NQOe84VKxYPapM5E10cmDY
2NbQch2wP3dvtaC8GOjSIfWBeEvncMsOZtmpJIymTqfRcl2ttfd+JiQrxYDBmZJn
3nV4CUMiQ69jEGYLVmX6GRT2vqCAepk3rzYWzp8ChHaagp1tE+D8K8iUh6pOeGHj
MZG3XXySyfSpLit5ANcoZ3AzjyARqNyBILbTDIjnvVrC70oPH/rQM2CpBU8vy/bX
+BWnLR+rCqS2FywB8nsbEN4RSx9oIocmxE/ZYPQEZFBaPihj6vgIcmX1ZJakpPa6
9JSV15OHIagZ9+pIMGNy5n/2j3vC0ayhlfmlsDLy4WGqsdpesUQjfy+cm2yL01H0
TrBHXiedeyNlK+SDnx1ccPASDA+wJVUHeHcB/24JrKVbeKXZThHQ1yY4ECSVvrA/
MDtOVTq5UEOTHAHWC445ShV3gjf+wJxRQjSE8w78tdaxyr0BctkoPvL56ErKqiGy
Hpm+n2MzAhujFJmOxu61l2RrgvYjmqZfsMOY/mxiIhBk/JY4HClGdgHdOPF5ApSM
41zQFuUAqxkWTxO5sOKJWuShOxZbUCB/W+YyWp7e6OmihORta5BQ4P6CjS4Y0r6n
WrNLgapLdpkIe14ojlyIYwG0i8CYnFfQTFhHhr4K7Xm62ZJSpwx357DosLdQQ3le
yZVtTuu9DVSGaHRafJMIpVDCjP6aaRcEAdYopKTfeMWtRA9rJxEmrnN1LjSxUjTn
grtai3Hkyjj6XNfRnoVNddzvCPhkkgRCDT7rSThU1UaSBGycYxXn9HkXFtn+8ufo
AmoWTLrXiHPhXzbMaF3Nw5T+mixJ377r7xiqwlQz6VnEZ7c0nKsFpH8+HYLfHRzh
qI0veZFXzH5aV9hbAO3UBV6gB+WOtAvm3Ua5C5AXsXhd2IZeyVogD9HVFhtMSfSq
0YM6PT1mt1ZGIK5OkyO2I5a5y8em2clVvoSHem1RGM4twDPJSCBQlyX9c09pc6IN
5n8vlcoxLyf+U0IftHg3gVH90cpwqP77b5tKHPQLMkgcIYwd7NEksH0wI8kqPsMQ
KYLIW57JOE9hbsbUS5ycUaEDg63kJnS/Lo7cHyruaMNb0F5Vzx14wSJcfiewn2xp
ReKTvMUtEfu1GcHthANOfNVAaDUlLxxvp/Y70VungACMro/jwHNppFRBglmqBATK
qJk2a39RDUVvq1jHMC2qzo6yYJ/UqH/oCsBhxvSQJnXv5vNIY06E5pReomyJUPuO
/c08RQNdk4VbxOfBVF3xTphCWV7fpJ+s0tO3uWAdW4plQG1dDilYLc7fIFSvMIP9
9dY7i9linCLW2psyn/UD20FXCFzP6pOZ/rxDB6zaqxgr+XsabGoaaO7kiK7p8Ui+
2nwcWcppxE3YyxTw/+jMtp6GObsDA1Bce0VdJoRZ+TUT0P4HjQOFyRdV4Qwj2te7
XVbftlJ0ljZ3VNsIYsRVI60XybV+M443AL6hhzDckLFTHNrDuzX323nydg387TPV
2on6OG/hetAlkzdFq4K3tV6BrEPMNcJUFfgDzEZSxNGMhzi20+l3QGBbgLa3lxJ4
6Yw+fvAWocC2SaYdgLv4KqNDQThWBw7ag9BHV6Ae957hqFBFgOjYSgR3tD8wx8yk
XMVH6m9JO6D2Y9AayLEdsaJr9jH8ObYNXhvRhYNo+sC4Nc1cLTL66COh3vInYUDn
Xam30jUfXaNxUKP42eVOJBiTaFRHCIwJAsAFvwEt9xRUJYvcS+0Cafa+pKVvVvvX
lknfqn7aQvUfmzEMMopmBcidUO94Pqb/+fEpW/42WLWsGXecfkbUXXR9WuaKZviK
VifxVwMYaSSWIl3hbCNxy+wfXN86F55tsV7au0GUj4gLXHN6iP2O5ZPfy0k5Fbyn
N9kzOFdNbzZUaXMm8W0JCuSLVo/e0RMIKRlvITd5+f5trAvxeLNzy9IvNvsA9WrP
hxcDkiuiYIR7GWC1zDLwcQ+JmN+0FcsJZH0TepuWhblsZ/k4EEavlcWOJW8lCHLF
Wq/VjTHfkp73NJSxacJ7cxIfbK+GAPj/f/MH6ofPopETz3u7vMdlOLqEwpyGU4Jp
DyAwjDZM+ggQipxYChsApj3oyB3qbJWBUgXiFb5uI8wjvjqi4PVpj2i6oyO33Dr2
NF2l1dPh01TeIS0iaA/HVmItLQWgpsyppcE+ronZ0cEmThm2vxUHpLExOfRTMA1I
F1Si8Bp3ALb+zi1t8kTtbC7ajXQD4XnwAb/t/yXss06z5qTnIkYNpWJv4Q4Cf4Ox
PRoo40ok7BHbeIxbrdJmAVlg/9lNPnEZlmfViKihNVrC4TyNpop9pbSos6J4gUIp
d64ZGuFSdeNDQu+7iL28cijoJOTbJWtwxQr/D+peH4HkKyu1QKqhbTGrZViQKhr4
A7CXIo1XbZAW+Rs4THbyHbbksnUVHxvx/XUg71s4AKe7LcIPhBoSkZiIqnorsx9j
XdArHoJYNCLSEvqXq943dtVpP7kAKEFYuBfR53h08Xc4P2SAcwvhl35Pk01TZs9n
Prd78rs5Z0C44RPkRUdErX4pKEajezr+Bua5xzRHFUJHk9+9bpjZSPfZ5LB/HgJK
vq04X4ws9bSMLYyTY5uCy+2poXPBqFFxljAvTL2Ux0aQ5b8sqs7W8obwCA0Kipe3
lrALgcKoujo2Dc+sNilqjwtT8t33ehFhhKh4VxVib6IwSQwCYB9ZNZVE+oCgdaVj
ir0fXPBUvlFtNvNrvCMtsRbaXNUP0ZWp9GaNBnFmCnsK3heYUaFOuUAqvHl1Nt6U
ZEVKrsMlNddVOlI6WtGFTCHU8zl2VvRn5dImQ4XQ7STdcijxLw/x10gDT1+umA7k
sLD82rLEBxWfpPd93SwWm7VoBcYewrfGrNYlO84rC96fdpP/z/FnRZS1C3Vz6rYE
u7i7k5rvdOGYNzLgky40bpTvTsp+PFMgzD1Fp9J9edDrBz3kPITe79UgeNYP8zw0
CmHv1k6E/TgurFnXmlQu3VeMF8t6bmWbV1Ut27nc6g04B74x6mZj4bsvg1As1mab
oVhSUnM7xh1rrTxcuesrYdlSmUfqE/hIo5Y77UIHAeqGv6mf2c8I1D1M9KDJVamk
JsXfAcqW2d4jZxwYOlMEPS/4T0CYzUpWBwL1ADdcZrj7ykerga2s65tukLyTWdBZ
qygGYOLu9fXtqPhf9KnYFzqxZIZbkxgW55n0JcS1qLnluyEKg2WglhQ027lNfJKF
wn3BmVkLIY0I4UPQcUa8pgi611yfuZrIjzi9JCbyiW8jQgu3shZJmUSSpuGsds/Q
GejnycJ2t0I0nC7eyLgnEskTGyV+5WbhNFgw1benmIDADzsWo8WFo4qjERu1ac9D
3UIsDXyOSrmOdirHoKi8T6HxwHLyClPzjh2Xc/vhYaX6DaLEmVaeBIvpISoduHF7
hbBiC2e/67N4g3sF1DCp+N9yFWH4SOHpKz2CpK6Y/sQiglK1aepbH8648oVhY+/D
lPDYqA9SgI3UOhgF5ntIGLNDhqqs2Or1EXy8zfMRgIKMQEPQGTqJCfbiLEBnhxkL
GxDLTle9siPLxwGZRuE1vCFWWXjEvN+ZCUYrF/2TxgCxMUdoZLkmt3TCL/46kSoZ
4tKXC3C+gDN89mxoi61JqNtXMk6nv+rtVV3Jnv8taitWpiOxWvkGOwzjfF9/SAIS
ivd+gH9gQD04/nWQ9uflIl2NXUQ4RDggYsseTnlx927l+U7cx0pamfzjdSyx4GJm
uWmKPDKmAoePRldzx3xLJ8iif6jUwC+tLSXBZ+V7QVX3hURSqt0gC0MjuDilTt6Q
ULsIV6HjB1an+hvAb7qHSVXpuRwcPqbjzJHkGQoV9hg0FI+g1l3LdSwMt9lEJex9
6t+vYLeL69K6zGGqlWIT75lBjSN/7JXjHt5EGJkqLi9ftkBBUjdmtF2t3rJnWKEe
a2ClqpmXOLmNZfgZJzf3d7SzzhKEBOtDQDVVvzULXV3mFYxNlwy5kiZr0t047SqL
Y7fz9EuDRDEv+nlf3IR4UPB+CmlOFhrJX3TpuosOgC9xEFpYVocTSmG+/mWmWbvW
WQb2YNEx3pEGjjNhrzzMUt43Koi8UKweJg0rZjjlefENqD0asnHotnVS+Oy4+SnK
ucqsnOxx1nvUDD2xEhK3xBSrt/EhMPeSBufeLxo2CL0Z75hlNiEJEgQ5xdJRxX0z
Ztvc/D+2cn9CAm+2JT2YRfqv5Hnzp+aG6SnvpNubN2jPbuA9jPTe5zJHzv2V66xC
VnEQFTqU1dVRqhMIUB+9vVtTNS2o2kWPi6dTfk9IGNwxw6nIsKyLfiV5SKWZdYBQ
RDGgjYpQObuXQKPTj36mRzWLqA0P7exUSn2WBXgRvm8Oe+QdInNXXfKwoSwiqaOD
NXRXU8coRPfSY2ddlxoWGbhbegk3Xkr9+fKVA7E1OZFRhinGdhwqBrDlT9n9FqCq
EDP24DiuTLIEYhzzsgMznvCqKmwJiw0pMGjfPnZj6ZXQn5LdWYQfHKPM2MjC4M/j
icZNj1Vb77MUFAFU6NpsfYbATtmDumLSxkd/r1rV4Aq2ksCxWQjy5uAJU/dT4XXX
wGNaPAbaUuyheZLn1BKNynlFTGcNv19t6qyQV5VeJhWnSaUhhDyEPR/OuXW7K5SN
gkV+40jzLj4sks07QBWD38M4K4doCpC0ZtueJR8i8bmqs+u01jiSDP+msWSeUuhZ
jMOZWj9NNs2hkSsSBHvwVN5ANBJulDbAXgL/UNqP/v4CwxP+wyX6P15bDhr6rLvc
KARvNtoCOi0NlJFBH+32B055n32kTX3nSx3q6eV7Q3k3jp8GAuaEhjR2QZqQUzMc
JR5gkDIYa87MR2NgYlZUNg7H5kQPUBsMtAArEbm/0tx8Zzs39yhMamwiyKacFbyQ
CoMtC4akaj08wkNR+JuAcCmksu08kiI5ZEJL821O0ew0B7EA7NWRDSChVK7/wh4t
69/8WvDpCuVDjpetkOIPqcYEhs20XwcMKdjH8YYE1ou5ywJFV6Dctzq8fI63xmBp
8szTcoL12DplwcnWbjGe0sGFVRJIX7xZwqZ1+TRbuLihWAvbgXJnzOcXG/wcl51J
hyvDg18S8T097JJFKqwsKyPVCZ5TQODnG8vYyE9X6udWnlwU6oc8uygsayip/t9k
L59tozdFApLIExWCrd4e2E/YRJwvyzpSH5n1SK90+ixPdirEophlDV4MvtGbisuu
taWF7RxCUWNRHxp1va2vS4gFcL+p4++ZPxsE6XNY/C1zHhIHsbGF3GVuxN96DARl
8dm28dl54nDFNY4KjFNX37Wt5ZqQxPRoRqtvdOPRGcYfMoX9hooLe/TBm+aIHCFO
dHGGnlvV3Q+g+JZJI4N6MoeBNHPl9Xvu9I1MvgrJoCdCwNzlGSKmv6J6NvOTG5sF
o+2mS5jxqsg+m1Xb2VL9JlwgxEqCnxn0HbVaDLExZ3XwctJxZKXpN0lR//HrIrxp
hS+5j6BjK1F8F5iuMUrxjM4m2q2ioPyg/XKQHasdkLoujt0GyiUPbXaogP7W1hp0
Cp2lu9Gx0q/mbS82BGNOGiKE6m2+U5eGBIkobHN5ZhVZPet1P4OyEk6n9j+E6bqk
360d4X6+JcOrjRoWeDGwPuJ33GOvHGrQQhgyZTSecXNLMB6P+W0PPYXHiZMUIfx8
rJQ/lnujMFewvr0FXcul2a99iRY1uUlm4bCvXbZMKua05oKuSOHQarrV66+VNxQL
AU63l1LjIWpvd1KRDScmuK0wauBsyhrsRkkF14QvzjMwoYa2NBMX+o2K3z9lxH8G
TgX1J5K+M9FWk1jKyezbgWrbqVbRtkcNvPVAhshEFIRwV0HJY4h4Dzj9JhcS+dqH
AR8cmihfn/QM8BTL/jC9bVYP8IaVcTXEDnJbuBBT/BxE8QnnfDEBwdPcIfMv8BGj
OS6WuCISxMQgdDgKhhHduHM4fFMc071eyoiWEpNDinJKfdmA1LklPv3vPkvmbN9R
yxW2jTe6qvfKSSXdHoqgiwJ6BwUPJig7oNtNjIHiU+nsBy5VqvB/Kr4N16NU7cQZ
F02nqrhPhbKPU8FBfVaCmMs90KrnflspSVSiX6RbEcDRFOyy6CZpPD6DLpi5I7ty
1gOOPmcahBmNKdVacFXk/V8X3C+BIYeSQAENZaV8e5AoQJoKxZ5bczFFAKoqGXD/
zbEZpmtuG00mwzZq1ecsziQoSym8FqZsxMgIrggv3NQQayknS80SGHXsl7ie/uYJ
efEoAewFS6n0aCt5upSWWoLdOGjs++5uWcDR3uf5+PauYsZC+bv6lyE+m564t8po
D2FYvqUDSrDN+90yZLL5Qg/rxN8TGJP15Mv+C04q0ykZzO5hFie55afSosgsHpel
Ky5UxuxOTsjzCucWQ2rlZuzLkHsp2rgl1UHBow10rkQTa3hrCNQOD4bTqdp69miG
qBy/Hh14H7T3SoqOBCYkCotXZUNZGbWXRYNdWlx6rSSBQvW9u5+tIGTvepJiQ2yr
Cx28O+dBUc6ugwr0H82+Yb9Vf7+dqa+a68ieTZTpr9bt+tPvQHzLNx6ogHhfGpdc
U6ZzR+D+rBg7QyfQF7/WnlhxxxHPM8z5lm8Kd9bLUkf8vXnhRBHRfpOAxn5xEHlo
KdAi2zFhjX4LRzDyE3/HbUj7yePktnKAE83XQ4d9B/6iz1idzTs3hF4pbpQWPCzH
3KmHXr9sEyQS4DV9DnzckdONyBbiK/UQaBx2ybrrnt54+BywAHP38jnGVwxjnLYb
Hw/CKI9OpTxTcVIxgS5DeH3OqzJbYqMFeOhy11dKbBoWa9yDA1FZaeuY90TD1jZX
eGsF3+F7mGMp9DhWGXzjoSrFMsurs4kVtMlc5rXGDjx4IBbi/v7qbkYhgNkEfMTB
UHIyuXPfjHzvpxUMTlxq4SbkOePlfEwN/DNzBTgJBQgWm41KSo1m8IqwPQ8fGT1O
lKgurusPD2uc/vsEBYpMxvS0EZMr9UiMG36jLThoQtPbl1ARyoeGnP8CzZhllXwf
YpyNDMEV2yObotgP4EUQrB1hJkXBJz41mUML7Bjd7zV/G2VaowLf9RQYWX2tTIUh
GCvJ3zbnKieHmrb4QOo5bBRS8ZbqtENHiFajuz4TbgH+yfsjwDS8IiE8dufl/HGh
jBugH91A5iQqAtO64Pz0OTBVO1adLrtp0tcyJ6xsLVJqm9LUBtHTytppGR1L+lEW
3tiAvFuxg3zO+Gb++1B7bQ1oL7qhCNP3J4jPbpVPyjaWN7/RTFQvBs5PTN5iBQD3
7n0yx8zetIe53rhgZWSaNOLM1pKCdtu3GwOUnXHYU26iSdFSb/A4FgAc4QjBJ+5V
4uuL64YIMeatBXMHUbCRJtXGusc7dSSCydgZKvxHVquCG/4NIf1fW8R6f6jUrHur
0k0B7I9GvYTV1gzCdVqNpKWUbtkznQMfjrW/XVNBIjSi/ar5XoexS2XjirlWxylu
b4N/H4nTrIsZpkwo/3+k4LR18uYzDnQM65op1kXHq+3kUUzXd41BbG4SlSkUMCH0
AcvjWkk/KDDFQdbADWZqgGXg/qjQNeFCKchMzLOL4ih3RS0X7vyS2Y2OJZBsDgnw
X/oKcS2XUifMYe6OT42r7GsWjAY5EiXq0guWaHYF2VIONfgjNqcyihN5TVUvC9D/
HidEdW7R45DMuBzUKpheEGRNQYzx9iYVN8etw4quGQHZiv7q/pWHb7C/+1lnQ+eK
zOthN8otKPkrgjqcOzfYUauE/JEc0ewtpvo09xnTR70C9OV3TleHxqh51A66jh5v
4+g4w2ccQSWuABGjsCq2DsTOzO0bzRIa5nCDl/cJ+JdXFXaiyMTXqiFwxPPL2mbG
4z6nV48setQg9gYkrziZQMzdoE6F3tXyBRCEPePsBslFgokKeTJSMdI4G0TdlNTD
ms/81BZmFKo5n5DwZJhOsyJeeZsNlWUHqovt4jX+di3G5nqyUZY+JpCt8dBZKe5q
n3J77yKrBvF6cOHvPWgae6i6Q05eyIPUKp9X6NyCczf2TGtzxAuphxjdvUg9EFtT
VF55jaRd7VlGP8Gk0xHZHeevU3V3mMM+pTnx84Izbb6isXaRcrH3TH23EpTEa0kQ
1aKeF0CIcUMZcccJ8bxKnjcXfnzXLDTvft3TnbrirfnUtObLSDW46IoHJ3DSt+jl
0DTL6W4/+fP48OZ4u1aFSqDhIT4MFdSbA/kliO0C4W39MoX08KXeu7C9zc/nBYJ7
41z1ouI7QSihNb58SgJgLw28FPNcA6bqRPu4SwB0ITtecE+MGYPwic9hLOkANFCw
90otK3f096p0H4IWwmxazVEjxEGughat7MeEHNy15dL1ddhY8+/ozx25vEBVL971
SdIRnJ5LdleMdI3B/dOsmzoXus3GaoqZckQbasJWakupmpXIe4UKj7IdZiSFdnDq
AxgFap47tWvuHiLQ4rAasZQo2kPI1cqOFuXJSOeOXdlEZ53Q+FvU8CBfh4w/YhA5
cdVHiWSG2PC8iAfBMJKiRWr6c+Qu+NwuVaPChd6AOhY6+GhmFVtv+Qw8X9XsVsDP
+4fw9yc/EDzWoHl5SYC39fbqHr/05DaiTZCEvB4OjtoQdyluLIICW39BlW5h4I9D
z/nwHZxK7JeuQF+/Fh4on93dtU3KokEebB2TvDtKm/eBrFT4z30KrQzt97T4xhvC
tILgKiOoVwACKiy0fSfCa5hx876iwe98aJSWAyt+nxFTZYh9AvQOZ6Qr53PXWwI3
6ktwsvIzBTfTKMr+Jpt9TP0KHv6ukqqVgLKCrYOyvddQFHbrds2Nr+VdBAo6JcGy
si0xriFOZXNndMwVhDJe2w4ut3DiY61FhDFq6X97twI0XANGNhk9ziPXsc5BxmRH
ej6A+Brg/JPJHlGabtLTblMjqcJWssKHedu6yCpMvYuHrQ66RNeHfCc0jfVQD6yn
GRAyzQ1Wu9LS5zl9QayuUFUrLGVRadZaP0ZiteU1EnfjvKwt6XXmUM0fhfAQSWap
d+HCdMZXOIv74XR/iGKeLN4UYPMO7ReRV1rG+GLcFYuHhR65O5qBFbZTpaiIdCdG
ewmD4mxzw9EjhbUdS3Sjw66ZqFTVSKLcdEcS1zC0eEJ80gg5wdNR6gt/t/wdikNk
XsGKB/IkPHqQDx8KtpgPt3+iBt4xY6dwJwH0B5Ix7PCAPprPtNAJmeJxt+nNphL6
W2S76rbAZ6/gOaKlk7g4+2qKOh1lqsz4iWPXdyzFshLykmlWriwgqnOb1KW98n8g
+r1bNfWQovrH8t0WIn6+D4IOb77IsQBsZgJ/P5XL9pt2sJhUnJm3Dof8DMKgD5+I
UiC45McaXV+8lfgF2lIF0ejnVvBeNq6ZIJuawldN6jQ++Wld4tvm+gSNH99sTXkN
7Y25rdWbj9dpaz1/X2tmiQsSDWmcsXWpjlFXeLBHzAVnLMfKmzV4lSWLAyMdHoiG
vjkZh/xk8ABaGT3hQwBJtdW/NTq1YBezqfE2jiyDrWvZDRDwzXYoPiY4zoQCi0pJ
/e5BTA/Ex9v7jd2JBMZRC71bUSOTVTMQ25rW4lQ/K8QnIqnjtBpxG5pYLJoSfuxS
S++5RLubDnVz1yugo+ZNV+oDGtd7nQkaBYlDrBiSEDJBCIaBOgTTKmUd4tmRRAow
5ttG/zVY4BtPlsYpfFSKqPnvi4M5CNFB7VhrOb0N/+NDDAM/P4VV5EYmQLf/E7BN
QSpWmksJn/M1R6VbPkrrqaymhsGsldaEjr8FtPLTp4hHNEZIM+5Oqi1/LwpWosD7
+LWH83akWT1qY12zOgwKJ54GjtxI3X7qG2HqD1T7bWOYOshOegSd1XwnJjNENRPc
/2ReadeRxU9D3nTZFzfADddZbviiwae1WkxYIQKPmbbUNdfKfG+7xFVz2am9fFXB
GnKDtqaalqTMzjkDtdKCo0AvZPgjNZDiHy3UD2lPcbRuKnLCPIWCdUXBWVS/5qxD
OeKX3ZTPB86wmIJbOYVXjKkSDDlFKXb/8rvHIR83IQwmcT0IfKfNpspHw5hN37LQ
CwTiSWIeWUOl+tFrpUHNMdO/Aqq3RgoPZ1FHw8T4wxvmNkk0mruTr9LCGUQ5yrC/
2Qc/S2IPjl+n2qXEHg1J1JfuarX/uh0TdjycpdV8rCWzQeCzeh5IOhwNKvibkAVa
kcRIwrLkjvlpmHtejyDw5F3RNsXiMgLpTXuS9qhFDeDpxQVbpPWMIF7gu9bPaKbE
+kJiuMnwFA+ddUENPpgDw5ghXgEe8lEvKVjZJ3mfAXBqz2neMJa6H3AP2xfAYjdB
G8IVqIFKC7Pqf984y2Uo1tnB787R9r0pLBQxC6DDPNiPPBEWaXjKGmSKw4u53FK0
PcDlObvFo7EXvMdGQhNvqoh5I2yUv29+lSjaSmUzrv6ISQ2yz9rL75qgOSUhL+hD
eO3nFBOpWsQW/97FQdGjNsro8zUEyEcSYto6reTBxsY2mXLmntpJfvyi4Z3INBPm
xmEY+NedkL8QV81s6om9v6A/PAcNJSozl1Id0WarwY6gvwEp6jLcngyvt0LJ9OHR
jEt9swM9CfNgz4HiELt+czNvgTJCX3NrbzovXFtU2Aq07xeJH/qxab7ykQqGCfq9
naZ88Jdh6sto5M4agMbRB5eFflQynpUk6IYdLaW/pSNpvdHl2SxhlLyYR31KwOMB
q/Od3B7ShwzcJx0HBpJXuQwP0pXapMvjck/11OA0r/DUprNpHrMpbK3Ia8/N+Jk3
O+UFO/TECgaI0n3QCSK00yrIb2FUOtBIY9Ysyfd/xI5jjmHIipNhxxqiF2pVJfMx
2dPb2XMa90aUsGbRJapEyl0kNljICo1mGIpcdHBEEmpTUEg3NjOp7+9CiukiQozd
Ooi0K7iDjzw5axj7CchXC7UZqpJ73wbnJmsRYoIQv2q46c7LJ6Cw7nzmA9EAeAsn
izWx0TVs1J8XZWOAiNJBS9wqjk+tF7mNQ5JoOVHOziw3Qb8aL5Wee+aN5V6OQ7AR
DQuP5G7XAFg9N3FFPmWIRaslJDmn5e0lu2wdcth6fAKd/EocNc2Gl6I+0ODwydoP
OXKhFe6w2wMzf2awVzfq4SnqG0RFePzYDjgEaaqMCZBppj1kFBNLBG0UzqQOLfW5
l7J44Z3bEvMlOHpuQUdp0IeXHdHwNlRJHmYe8GhDRM7finbypSSSMGkVwTqg1f9W
mMct2Rm3Xbc0hkl/F3ox3+BBSSZEfcU1mXUOZ0hcpBMp4imVX/IMWphZIQfkKYQJ
XLPoHZK24Qpnv5+g9b+GbFahlA7jhiP21mif8wwONkXwV5acaLF7z5+5JAjRyspX
Y9dMcP4k4iCAWBCAmHxaG6nCUITBSPpSKfdztFwM7SYiSidzUpaTVwqq7rn5g6B8
cMyS6QHUpJm2QnPYz8CC1ENYu2nIoYSVenAjzxwTazdYGdzFLT6L3l/NKYyFWGTN
F08wt2Z/r56NLqt2h3ge4k0QpHm6gbSIkhVcrsiK3SVyd584VpE6xQelQNzX4Qex
HTW2XpbAtv6/oFbKOvZYIJZRBpgn0ko7I5zahdhNUemJoVo6v4n1OZR0cv2/cOL/
oh1eJ9uL/6v1Jdc0enfupmPMq4nSFTs7mYcdDH++/mAT8zCb6RrzEoFVufHDWc0T
ZXy5UXXd7q931qv8SxImPC2u91Of623d2xoBFkuKIaGyBWp2CYLfKC4Hn93MXRFA
ZgfOnJZsFmFYoTAOGhspooex1XuJEp3FrNMR68hEseEyRcWUNAsrsxB8xz7FyWTp
5qujh83Su6M03osAf7RAbInnKMlb6/6iNmeEfjuQIaCeyFh8Zbu/nkGKcr/AHS6L
pVFBu1Re2oBa0T3EnnYBQ2ZnZpq8Be6Kg9IHabh2L4wTkWjOR11idlHcgAu91zsZ
OFmiD3DhEe/6C/WGd5wckEwvhkMc8Hf/XfBNEE5NwVmQM93GQmg7I66NkYNsNcJk
ZC0A7zMdTBf3R1aAaNRwBlFI04lF4zoNFDVlYFvM/PyRkC5uBSPpNmksshsnCg0E
mrtK9yVPXzuhwU7DV8E0Sb467F7oYqRw8voI/6gKFefJTp/8FIxcQu3ezhOIQvT0
jftTQhItAfhy0CLec/Dzzmwaqd3A3egSnvzADyTSSklc8LpqT7LYugP/B1uepy2g
pw7TU7R0uLiCH9iXqu8yon+N5qknp9DYSM9xtf/nyo9FeWyMMcSM7qldeJxUd4n7
3ljxnLnJ2pdUgSiLzIc8TBuJN4B5vRacZw9zSQB2qi5b35ZXMPNOWUlgy8IVJ1Ev
VhQ6kLRBOrBSJVBibxQnw0+jSEsgfW7O25n7LrZFisywtEK9UQtga3+NxQWY4W2f
gtFNspTwG67wIk8aywk7jPWBcLJWT49u5fBfKi1s3nY3CxTLsBbBlduLotWFu4hu
bwMtUxmyBY4yx7Sv2VyLr+K9W104rpOWSMsVspIdRhwwTM+rjVz7Pnbo6i5kZuEA
SvOeyn6+8zyPaENv8LG7IGUK79A1kpJk5y9hoTrc2n3joiA1UTEqpUgQF2l/GvEf
dAi9bZHgszMKIB69utA9IvJypy1r1yQV8o6BxbOniKtPhkRNlTlhN0AC+ukP2C+H
xS/5W5AjcWqa53/LIofBccpJcpldtRdaPFrJoRkz2nrthkVfYMZBXugldWqBMyzZ
jJaDjid+7llp4tVV8vbvDiI5wYGJqOh9I8TefCqm/wRc0NTL7KsVih9/8IDc1d7l
qpos7MxNmdDCLY9llvEgq/RbDrIbQ7Fa5XJ/1hbDeCdYksvuOdixYNBajO7zKkhc
RWrU+BQuj7cyKX4QovWaFijG4AVa1lO7+6FAPoZBPwQhFqi32brCMeqk0N2mHz7d
SYEv4OuEFfoIo7pHiuDA7XQiW+x7VAibC8p+loIxAqA6TNWve2otMjJpoSUBmpyI
/c7Q5z3WcBLfu3yp6TX09bIMFFKBVksEpNsKB29LBG/KbqPWMJjNhQ4Gr9Hv/IfZ
0Bra26fcvJGMKDpTdv3FGDuLaw694/hTsm+iOt6h/nE/4DkPlIjCEpUYsgJH93tR
AxHRx7PdyUzMunwajQ5fLlIJFsVyNa77pjBhNrl+1aQR1LGBBjilJ4O9nzyJSzb6
L3dN4S5SyXKsnoUoq4qvRJbBdadWAymBlAz0rbr+dpffDfEImGCeC/nJVYLAjdiQ
jFzXOxSTOEtuYK2wzNp4JR9/iG+lIrtTr+288/sYW+xMDHDebJwz7i8P5Gs/p+Qe
le3fds4AtJQh80KAov6fBu9UpJ5P3251AV0BGcEPBEYyL7fK+FsCZrNMjyCp9G7y
hj6U3IP0fJGsSyccmAlCA/xjg+e4BdMiErThJFFkrmz9UWSxonUOxVYPCdNOru3F
RJFuNWF7RIFygdbEA54nLKpRWm4J/G/eG6nZ0pXPbrDWsDgrTHWiZN/ThptiyuyF
QfHo+GtXyML6v2KcQVEGlwDLNKK6MS2O5S9hXBg76GMneTWvTOe0r6R2XYeXTQyJ
/iwdJsWEC/UKRFTInYe72j2DT1lf3fUcbFGPxVYw0+hOnFWa4RK0paP+3VVCz6cg
O+gI37t8RAyTUH5+dpckmuIuuIk9TUY5lRDxb9/oJj643Q1s0znrAQ4Cc/ucJirC
JCLQn8HGfVR5AJ+gaDMrIjm5RA0NQauZ2RnA2IscW+LJRznAunBV4CltFwxhkhF+
es1J/Jhin2jG5ZCp4mOCD74tJ4nhyVuA51UzMxkmOWnwH+bhzH02qQ3jaW4Hild9
n8DmZgz2OHo7+RwxN/z5wVG+Gsmt9eYIJDGv6DOpbPXniqBu8Oiuptg1XOR8zGl1
emqDRCMTzl0o0kk/6AB1ID0UTmT+zGkLM8l7Z0uoj8C+lesi/9ZZSRxYdZQqGUmH
Xvjat/BxVYFrrEKFsOZgsC86B0STmsIZd4Jr7usUb35+fptVgvdIq9VMDUDda8Ql
mI9kd9ou+VtzDE1OdrhPs8Ek7D8D9qHI7n95BKAwaJDHaQjZjnvbOhjD0oXa/OTI
5ywR4wwIKjKZBkkZUio0XHds8y12IEiPADCEYTb15YI8oTJ/s6N/tVqRFy0nta/a
rPTjMkh9CbdUiun3hytIUfu5lOE3vAni9Gd7eLo3cC5hvNuX0jy4nEAAsBaxl5wM
DOXDugxjy42NTmtSIulFGVWMkGiVPvQbs8DauPoZjrU1HkTYK5j6cn1J4pHEviZP
NpY/gETJCVwXivmp25Ca7ax3lN4p1pAHBbNc0TxQEeqV75fCvN9LgiE7SAYxT4t9
V++vPwSyxVCBldZaOsuZN/2EeZJhJ+z3thTYzD77Yq5hXmDdW6rltSMu4OOhr0BW
iccMjQrVtpeGQ82swc+Z1teO37rwGggfDVNT2v5xbXTun3wrQEop/ZF1KDHrC1o9
R0loQt2UE2IYIUUxQjTupsrczBCmknZRUbY6pdPCb1DX7iidROuZpFMp/ZgYBdU8
Usg7wKwQVfZ5Ezk3/q+Qnt2aBFx/G6OntYPBeZrx6l4InY70INPxeK/npLJrQWAK
L4VuhaPV1ZpbgHv4emlJmwoWYaOqpQgluMt1Z6HSReqYiFWJKBu38BvjUKqGCKyl
3szwRuxMYJjxA4DBDZqDirIIyI26T3kjfzNPKDnU6FCcStqEeSjsCvxuRCH9lPhv
UtA1w7uK10322AynC3q6LQEh+4PS4vcZj4yDQq7JTqTynqaSeWU3NLHr9HkE1oET
r5RnBEbl7JaYb2XUPffwhz3OMWUkaur7Z3NC6vVErRcDsR13b9DCBtDv2YgFipsy
Erj8TNbaRfvgLssJeFqn0FoR5CgLRzgXcA36XK6hoiYsDp3SHCMuaUvZbseZ0m/o
G0ci0b9AuE97gPpSy6eTgAgRYIa4qhRTcttSptR/N02jApdI40N58naB/CRYdit+
azGUx+jDXS4LT5DSO9QOe2g3m3Sqk3M/0k/qEU766oVRrPnP6M0RUvY4HzmIRRW7
F2IQqrC3k3lgyDZXA0+C20nXh3QP2Esi38Zox1+I4LQqluyx6ynu84mwj9FCYhsr
dwcBzZmnTlp7QdLZYiOrG3+wKhvmGBT2Hb+tkLUrRpE5JCLIpk2oEO7DQdm5uVIM
kP+xDtGUJpiM4Ov9zKaAZjtvjT3cnlOzHNjtUmp4eH2hpaxClGFH/+xizkgoCEdx
aW8dJcyY3aRE8ecTHh4yMnKQoTErFLVlvMkzQv1wjWiBIhKfQLVpR22TXk87Y8o2
TW8jl7bi9Ux0RWmb91C1lmybc8wbHezzTpWjfqk4CKxRjXNxUlH3k42r127DWilM
bckj9Rq2mh4vvkD0/WM6FckPoi3uIe1AJVcmcCwa2VA3880eUhNPZSokx3QaQswe
hP53GUY7vrsoXALdjJ0vNA7x0jTLlq3SS0a38swtPv8PEp21EbOJl5VUyFs7euCR
PMYam/Rx90m1Csau29npaXXutaut04U/IwvwVi0bqITAsY7mQfJ8n66fHFUz4pVW
GpP+LM49wYwVo4zjF2whgwgYrIhViPUzjbJiBkYRakFNxcBjLmG7UXtXCAT0E/lI
yRDZhBwhW0ZzPCanuXk5dqJr+cFi6IWOqOtkDJHbMvBrLTKWLBjchchd8ca8LnAa
+r5qsCQURmXMOV+zRd8SUSXeVE2VLD8wMMqMRddlIqURmtYbdIKpSqm0GKl+Y7no
K38fg5JhWlcVjPGb5y9gtUr1SaTx7fP1osIlG7RhIv97U+VTVaqwUW1g1HhGgwi4
kvV9dPDMl3e6zSHd2IpStghyeBzGd9CkMgYnQZ/mlOrUrtlgd0cQKHKhi0hBNZR9
6AvVQuNKFCELwODmWWCsKRUvEoBNFxVm/cTVpc4Aj131VUMpDtgceFgM1J6YNqDZ
acr5iiWkD7W2KnTNSqVQ/zDtes54VspA+OCBgJZGnJqNntg7IUkMguDW3cxT4kHG
123bJ0KF1gG3VmGzMjT/F66cz2G5yZ04F/fvaeihj2u5Oxz6ibGuDGamfERwoX+M
azFFZ4KHjSckH52LeS4nRodeR7ax47gOzyAVZf5zflvTG2AvBfGtDHNvsuRlhD06
+tPWtbLVRPt0Gcj0Gtb9WKj92Vt98t487Ihn0Vk0zvnquK4J7rw871vpra1TCQzW
40D39RnwL0QiDFQnXvxagCnTwxcRsreI/qUXQK7IdwqA3N1CnkhV3sJzdcpKKvSQ
vMWfAjmQip5Zt/XhqW6Sk0mysnQjA2slT0HuoenG0hWFtMe5RuQ5yp+ngqM/cTc7
1NnupFWfhrFfetvjyQ5gKanJucVwoA5y0TMKx+zctfdMRrneQxo6S97GCYD/6jQ0
bnASpy6aNRtHdT/VOVzhvqGdiU/nn6bz6w1uQ1AdFRt0vtQskEkdSJOuIOOYu35T
yJwUtusN1O+xhn/Hg1/qXLLG9Csmzo4gqinUEVI2jVqrMNLI/LVhcxHArOP/Am27
7MeBzyxcMJaeH0Rxo2/e4NtBt3od9ox1kEU4Ywt1PJ/+zuR0CtbDLtIOFFkSV1F5
tPDozNaAx7viKXBqthJXOu2mBODVWuf5Rr8Ahss++WooBif69bgQj+RUZBROOUB4
3fMiZyCgPxCVThj3pVRO8q6x4/4HPgDyVtTjSyJ7IunNr37jaxHnmnsii5fRR0cW
HyqD6UXUkTufBxbmShFB1L0i+ra+uRhxg8dGlCyjAF0DToT9Ztf/oCzvGutNpHhu
CRhip8yVtfDNhU99HDe4EZhhx2FizWBK//r0Z/jd+6lvYUdCYJLZcwSA0j1b215X
xxm3YBbLxibVVlEOQwKRyehbBm0AG7vEHw5NZsxCwuS35ENKtAP/q7JuetN1UFvn
lbeOkn4GiGF679QKor84xyRiJRJyRYBec7YtfoNMT47mYriqQCpzVwJYPbfBXVCF
HAsPSKueBFjhcV/+Yd3ciOl0xsvZ79h/79xW8yx6nnM9R+bB1bRy1PdOmRcb0o0g
DYFNTK9z+ONl8NbAzQH4nJrgJYVoso8KDnk5nJo2lfF0yDvHJiEKp9ayqpNdXMMF
vvARxgXifTcKriQWXzu3hDQ6iVST6MTKXnpIYB6Uhrxncs5pPingdokEUBNA7r6S
vBnM6ju8kO22NQedSTkzSW5HLWTEQJ3XkK9a2nqf9BCF8+ejsUnMbEz/ldSkj/u5
NyFWWr264eDlsJgPT60py30YrjW/6RhwbxAbdzFqzLYZd1OSzWEejGo3q36FgR9o
Axt0vMd4ne3/YtBMZ9En4euw8+juQMtpgymNmh82qif0qNEuwi9JFtQ9vXjYmkMl
Iuaa1NvvOaiFLjzdTfqtsxq47jgnHbblBP0OtW1OYcqBvjmkkUSSFmiCL7vm+pys
WxvMZNpX8iWsFY4DcnqUSGhGnnUnQs2834awrqOIpqLrX9bdJ8nXGYXrJf+3wuCb
KjeSDnBdWT0NyUTQLhphlDqvVLy4LyxgkMXpQfowtJp4gtFNfBspKdfAcljKIRB4
cm7N1+8U3/2l1eaymJJ5ODq1UHCr9X1LePBRPboWd4m1yLPVNnuxIZ1I44xf/fok
CS890hQOvlyShsD7JXCzWCboZC/+tAIIXDLGOX9OMhHNHKb150r0lAz7tybhwgrD
1URxrr92wDzYOqaAbp0SBsEX9EO9s3AlQAYwYys84acKEUoxxoouNw5kCoWs5Tiv
XC6ZG+vQV1cGR8o9VPDlyBMd+ii6kc6Ir2ZEX0zbbQJxn+tg3vVSZHsS/3iaiR2l
b9WVsQSfdQZkjnNIJJMvKWBv7xerITJT3kbkpjCMLBdezSSkbmDwvWaipNtB6QdM
hE+O/LW3LaR+DUyLh4dsMqfn7TutSIfZEugKGgM4V0Cu0Z8mbkrvqNtQ8hVvzhBN
XX7xU02hKt6HIH69jrUHC0fbgOFO1Yzph/hHfwF7x8ftaeAffNWVl3mnSP2WQ3SG
CHTzN/MISj6/BLY/fcoWTZQAeTF7R77Bn+EsO2Op38qxwA4U7ne5vN+/3HZ0cHP2
U18hc+jUgHd2kKl44Q/nIHXj1oc1jc6h2T8ILzTpYhdRh8TxkS08/OVjPLcIzytc
ea0YDpSDfjWcbh7NLr5nZby3cvEI4DE0ByKbDk+fep/Bags1aNRHyTdOWDNC2gut
OUxpSZtSlTf/S9MtNdaX7vy5zQ1Q+ynzSKKQ+FWk7rdzaIPO0UcIBW1EwYk2ZFUw
cwCRDzLIhUZc5ZA01L2aptbktz1hlIFlbHzumxtXzhOeGeamEX5ggOu0l+sX5+9F
RJf+lEJdIyBgGT8m3hBWyMacZKyvf1263sxZoTKHs5RKejgTJKERmOwRy5Arz9DI
8YBSTF5rx7SAshj5ipMWJnG9XvyOa0lLWldIugx/LWuzCn4aBcmezqD4AijlJfes
fw3yVOzOBH7tfXw4kFrhd5kGYA4YcfFjPGV7hAjUKvhanaqGOKVUKvKw4xOHcl4r
YSIui/7LetAE+xrishnQTJWGji1o6hUfdW1G51uKELJszoA+GULf6oZxpMlJ0kXT
156XODipPtge1r6R1Ldkg6YMwvF6f6qKrjL9jr+au0pF2pclc5Ws53V6hhbREt0U
lV9WS5MHViw+9eWbBRnvmtLF3dt9AnVrGMiJ+XznuAj0W/PdJDc+ZtttiyyZPX6H
XtbV9CMGykOCIbaXBLS4RmaXxifGtQ7WmOV2XApwFvm4MgHWmY/xOja5BnbmuM07
3pryyE8nSUoMMpHIlFl4o8T+e8WUmBJn35qMwAYhIgvnM1upRG73ujpZS6YpqdeI
dR+glaFSWWBYBx/lPaZp5M747ec2MuRPlrYerxGUMyAG5unQFQvpKoUQXC9qql3o
n0NWyww2qtCOOJVXO9DbK4jJ6RMP7ZvQUqhpESLvu24Z10g3opMdHQPTdD2Ic2Kl
nfhymRL3fUUXPadDMJ5yO4omBbqCnv973q/RtmEttJx8aeHLFyLJKa8MLf4+3LmN
BtrvKe1Bdw9H27o1V+LfA1vQCsd3oIdITiEF++7PzN5Pt/f/RBDo2rviZ/fL7g+F
vQ7fNYn3+XGdtkRKkUqoljgBW3xNAK6DTn979XrJ4bVsPipwgpNvJGEDHXZWlBQj
1952rm//oXpdv/VhbHRxV+6clcmu14aznupLm50UPeEuyLACR5HaqIJP1DE2dlU8
cG/RfSomGoXUCYaIGPUsbA5A/lYcsrSn+q55yxI6O9ktpYk9ziHgANhm96HGPmfy
`protect END_PROTECTED
