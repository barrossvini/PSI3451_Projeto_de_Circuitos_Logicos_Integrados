`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+3dJB0dc966iQnDq1p5lTQ22qKgoB1kb4x8akeEt6lF/SW/Nj+Cv24qMjG6ZNQDq
tDhrfyruwv7RLqdzvjhLJiwT4biSGqYImp/F6ohL+VQnXDwnu2rpY4KsLU8jB4yX
subusbw4u62pdV0e//jBVd4Y+zjSpJEGnSn4CZjDRsQ=
`protect END_PROTECTED
