`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jm215sLdzls+zidDH1avbFmGIWTqgieFjFYgqIqDjqRdX4AXXQuL7y6nyYn37DlZ
o65uxBO8zzfP0pmk8yiScxM9Wyu89mSn1ZdYg6GP3ftbU4ybNqqsw2sMltmRT8kt
eGW1svjkKyP2xDGcXDWPBl/wdRmYO1twUrXuHxBDkFn54Fvf9iP5g2AnUkTWLPFN
tfSq/U1EmSY4vTZE4MaT2W0C+y3GLYBLjImxf6kZBKLzFOPJz1DgQ+VHZfHK8cz/
cb386vEZCFWqUt+O88K/jqjcavMPDDrmB5SFDsfvTZ+okbv84u1BtrE/BSijJv2x
ACYA3QR650Yry7DNOrMAB3mQooZYYNdRiMR/8YVvEmnTF1Z9PtrmpMfP8Nd3RvHQ
WRBnNcfppKIdUTj4LeImZfuUDhSgHRQd++NcD67/XF7Leb13BKBhxS7gNJacocjj
39c+m1Efik7MMwISh0kPCkGx1udkXTt2d79+BGSCTAzVUl1Ms3G/n6skCAtJMtMJ
7Uxk8zjrSG8hlVeqhIOR3lTrXE+SfJJy7kooURUamGP6slHg4UtTflJLEkKQpd0J
Jblka/z9C2M6kRIuFNVlhsAy/+wNUoBVKkg+pc07nr7K9pfvnlW6szHHvB48Rqc8
+brgEoRIjHHtb9CNyhHcPeLXgswMuSIxrDE3c3hSZZX3DuDNh8jcHq0FW26BtQQa
pDHkyVHSapb1VweCvlhdx7MG+bh+ZA1NA5Xcrpvsax8VC3umE0rg9/INXlJ7+G5G
tJjg9nhWpg70inkKjUz/qoRDLUL/C62/5TPvOM+v2B/6NXNgV/if38un/HU5Nlsh
sMz3W5Qubi4KsvWSkiTPDA83nCFTJbtb6AvPjgrdIMMhOREEIYf79WeGwcIxOAiL
QppWauvcaR8pipEE3QGWKu9cj9pPfoOi+Gzn3mu4XvUo3xgcLY5DgmG+6dIem84Y
TnIoHuWjpFGdwkkFhxDUzmfIu5/rwOO7+xFB5eL4pCt71Nfpgj5MN4dKj3yDsfpU
+UEhHpgILnAqQ56JYsTiTxbkdRXMS3sF3XuqHM/oQxq81l5UDN9wu2ew4oedXb1W
s/my5OkqVierRwTuZ/6jhDeKdwClyUBaWx0LUFaNawMb02ga3qFh4/GCU1FZnh+9
L8nNqmINkzamJgWPCOKaJ+JzRsAVA0/tMFqnPIXJaY46LNkC2/Jt/eDnm9r5usKX
S4IyPmsCJRkOMfMiHXvlvFlNMFVaExlodXPM5g05YDO/1M1Lsdl4okIQqbgHqKfv
IXwKGq7AvlLsNj+iaqUWf6aFUOI2M3BBzwCoaECI4tUPmWzSpS2Ewy9XZYmnkvnT
lkB+BWQKhQlO45WszN9fP41AXaKLGndLqNbsWh1AI4V0LpUuMP/mXPrewlhw2OqV
UREekb13cGgyoI4dNc9kU29Fng7TtykqPHroJUOxC986HCeuggeuxd5HbTcOh1yI
c4jxmADfukagBYxQagxUNsKw4TWCYuJUd2PacCaUSv/uRzmKKQWcFS0WmL8TGrlH
Vcgj7MkokFiAvb4DPpaQI18ul8qHSvzwXRVxCC43EVkowP1WZ4DrdaXM3TXQ5h/8
4U6v4RD5jgzXtNDr6FIwMDWB2WawnERGulV7orVvc4Q=
`protect END_PROTECTED
