`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IdKpngouOjBeFjPhLsg6K34w/70qVNSnHQsK+wpj8HYBQTMqxiBMIpa78MDchaq6
KxvWAgRmYlaRIf+eE5W1Q1yHNZC/g5bKW+PZ2XktYFVxt+TL411iBGNnIFKyVCzq
E7d5PLicYtbgMk3yvKnFUbg7vT0ohMpsHt87q55mekNIBivFx/wQL1D/bzWa7W4V
n2kEI75m2WY8r3PnjNn+BRLlAEvoFXqCt+K0jO9DeIptr1+W/kE3PKMIft/8Crvt
enDTgZtGgTrEZWW2JYVvgJ5ksdtsmR4CtQPP9f4klPVgCujM8zmej3HyOMsk9UQ5
q0iTp6Jvh02u1MA06kieQSN4HKXu+9OBmmGERykBvPdGPXG9bSZOSEFNB/Yp4EYf
9lOZJNHD2/IdEDIZWwM1zgbRG2DkBwgcnrwucdJJ7p/6a4sKjTyiEIi5Hc3HHdkx
q5OXfGH4MgrVbguYJqozMeRi0SdXxwLARcBmT58VVkIQ+7YuCXTt0Y8/+LAFm8gl
FNIKy6KuopiG1Sa7wyKhmTRQA52qfHoKxzZmc5jX208DtJHzWR3SLirePP/HUESK
0nN2sax/zpewWJy3lH8tl8BGEUlYqKXgqaHk5h8OtpV+o2V8B9fLsiImB0p3Ayc2
5xAPK0pk8x8hNVZ/iapHvzApAQI3CW8MMcxBLMNURjwWMvDToMLsMjGE++KDTCOz
YqNtaSGrztU8hgjfp/8queGl0492rQlkUZBucAmrXZ9e9fgELAR9ld9m+vQ+Q2bO
giD//grIdmCOEb7SsL5OTFsbAsIR8PH+qzBV0gYP856ohrEBjdcCFSpdLJ+ivs74
Y13diVE5gygE3I/SN+ctaur9oTDDH/dEc94VdoYUDnLAgtNO4yYGiTkgpvaYSdC0
dlwxWag3ICGIauZHsqlU12GYMeBWrxTvEHW2+4G5iZWCK6geDOgMvugalxHZk+rP
cxV8RwRTMcT2oWjg69wL7yD1qI1KY9bcWTibHVTHRzzS/hEyagM3gMk4ub9n8Rpp
s3sPylCirwvRjMfHwCFHOgXutK17E75vcsJzBMHOAFjdyO76ilO33pIL1YWO2h2N
DqCvZm19QArdvXiJTtKZUhLo1amKHj95Ro7o4KdMxjXd/22C9xbRg3WeIPWUvvOE
JZE0+/sLOfjqUXJvUQSbxjxKmb/ayNvJefayAQ5Xle4GViSmiA05/TUaIYI5S21R
QDa/o/My2fl0CSRVzJRK15cKymKsj7Yi803feXOFMDzWgu8GqTOJAinv7xexwyiN
Wvf8Tn/H2d/hj0/h5hyiZHhIaMltGnz52VQqDuHHAgyJTiACgummkxDt1GVCEeyV
dLPrpQM0gBM0GPafLr/X3fBaKvuXLx3EctX4X42DLceM9PGJako4YOICXoArpvJG
tNR6BgRkkXo8QZPVHawfLA7HaKsPazGy6HvtHreoFhnlLa9HtR+PMq4SqsntjiCe
w08YxnYapeoOGuwrTtd2gG0i7joLxsjLKq5ifvn9wLnFjcFIrs4GmegyRKslS0t2
/EaRN4V6htgYpY7ybPUG3qF4O/v39tZJKtYkOz2iyftel2z9jwTRONtzrIvt8/Ua
Vt4KGbD9ELTCCDGZRY0zDiWbno0MQg6ScjLCv8qxd5JTcHdNJQCWH+0gueqgXDI+
eneoARyCB6yauIc2lZhzpvK7fl6hKZfpBzfs/b7UJtHfLpy9MKFfpMVhOqzX2NPK
R4MPoPHvqgTW/KsmecAO7vQvrD4NJCumxWV6zdl2WaUAqv1keA+LSNF8+3n/MoeZ
RMN03y/K6kze6C/JDknkmSMu8Xdc0x3jS1UNrpqMV7FlljZXXSZC7qAM9qnB1fiI
P6lZWYywr3RG8Qp8VbitJwWGGyXZAP+MAjib8DFh4+E/DAffvfpB0dwywYQDHzRY
Ch7ueg3c5JzljgqkgOd5lOvUlm53eATKoi0hxWUD0FARwsZewFcTKgC55LgbXE0X
Z8X8hBdxAvIsAb4a/aL8aZiKri5m+cYF+9wgvIbw/5K99tzkinZEfWu4MdogyGc6
+zHrYY/SUZ5j2t5w98RLNzmNgZPij+u9JsZ1/ZLwHRBCVnohO4g/TeGGc9gy2bCF
+xKZ980eElCNdxXcLFkARJCveV8onqtVm9X+2Qdap4sm82qSLy1aRufe4WeqyB9m
RU8DGr2xt/xyyAt2Il0PAQ31JlgR1A6AO3jEla7XukZi770YtNtxVbPygHfT6xdP
DjCefqKFrg01FfWWVP5Lp3iv1ZFP7UdGKvXJ7mmimZD4/bisZasLifS+g2xa+rpm
T1LPK0cvYf7PaQPm81NmSitVPZtMXboHKnSmBWmAfwHzkrNRzZbUTlNJsa2Bcs+F
cSAjoOs9SP8Kj1PgRnUXeqT0D96gYbSP1qPlbWB/DXU9oqcouDbdoFMse4urhNNq
XWIOqmb6vbIxizDBSUP0uJY0ytMCZzhFrA0r9r6FX9ITNtf27xIkOZ/+NHOA2Zds
o7mARnnbW6URAphHsluUPiju330L1iBifS3s+zoEikVXKkXucR2oOlYAk4LcTZ3c
YjWoSkN6wZ/jETORbDbnKOFCJwFCth0sWxqacv95LYkmBTyjAaSBWJ86dR1eUjX+
M8U7NaXMWXuW4SZXoUl4fAi7iiVvOPK+/g2SATHMcC3uBlwLEs9p5iG3lVnJdcTE
y7tVPSFWOdHjOoFJYChJU1CBYiVMBMkdjRxM5JYRBROrt7PSxrg0HqrRSOUBpnxS
sFbcUzuC9pxQZvpBIuyqNJAPnEBVhDJYP/rR94WvDarax8pjUxlHKuIWk4DzYtM5
uwrPTXTtEz+CxD0X2yCP8Lre4lvXHY8mstpE8oUgXLWbKYATw2S3iYHDkHMmE8tu
pWGjLbiDAqPSKXNLIP4tPHGZB4cmNK6RBfYCIQVE6n63MyBsoSaP+bpgAEHsjg04
mDtySoDkpqtEd2DmWeD9Z7JRdJUuUTaAiJpNuKet8+hmvRZmStrgOiyDWfyH4TXY
3G3tUKBxBIVC8fpEjOCGVSvcd5Vw4Zk1XNAXtuK0huphDBrUtk7vxAGphzGfY4v9
OGiJ0VC//W2JPcLjJLCNmlrbQxlGGUKD9ZpPrC6/aAsa/ZpuO9O0MWk1P/kVC4f3
dt1xNCm4Eb3aXB2rDh1n4J6GRAt9bVPlq08LXzU5FfdzeeJyFH94sAo3rIVuNd/w
GDAZ8QuT8UwCxT4efeZ8wcvwXYwGDaf2x2D8OCXT5ygRV3u3Kadwnf4iIdYLVGi2
f9q/HxoUcWpSApdFySscbyTXmnb4odECTEkw4m6c76lkho5J+sUkKmmk6cohfZmT
UWL3M6ax08jG49l8I+dy02wuNpoFL/QLYFOG9kYucEYOvaDMmv1wTCl9HHMRWVPc
YT8+BI1lyadjGHLySynrQXWJCU4cvrbAqSCJkfaCs2/y+H0+ssY6rw8H34Ujo8CL
sz+whMAI0JyzAYZp2VHcuwTyJChBtRKzJOQi82HH70R/6KLtGPRHyQq3BEJPfYGJ
2qJ7jtxwvyAH59S+qQYVhpfn8/GWoaAeqWJyp2uwgNOOuqXp6gq180WXq8XYbzEh
xwO1Q1un6hbGzAveEtSWYYYXYHNGmWZTEFxM0fI+e+bKUIV/ZdquzzBmr37lBxDu
WCZClBLC2DaA3/iNsH/5Yuqp0SSxgggpPioD2IYjrsRrey0035/UWO+u7RW4d55T
UzYy0TgUQJaapt5DNrPj0OBg4esQq6MdbxUaM8+0vbr3bjtZc/i6d0X33QuhFRIY
OaLSK4GUa33VNUKpAQb3p79TL43VCANHMKQqflGrmqe4qXu7wK1VsggeqaFmh57p
WThUMn0Jwj/6jhT4+sYLKwQbpCPs5J+HMC2YCQdCUWmtELrmTEFi0NJycnfuSFtp
zRAFIM3L3cVZCwm//6HPV+Vh4cGOCZLFHwxUgSuJBNFCAR5Z35XRGvU08Xsba/gK
xknBlQacIjN1OTQE2Q6BqI2Ti5Bampx+4o9EGvr1PktdJuQ7D46vSyr0BLkokARj
kT8b5SqahFpHa3EPJCk/WxcOtrEogFiilE1I8dOepVKZKeefs9aCTjmifpF4E4Fy
Z5NMPpZSSY1U+IEDhbvwRuO6VCXmSMqRvPphAT+yAH5NySwJP/9NHFsRTML5W0sA
ufSjW5zH/CWfjFyOuo1F8KDth3aYvAoiqVAfRiQ0bVWCZPFXW3R1LdHPcDQv8Y47
yN46IodYZ8a5U/zy+DIm3J30NaY91QnD4pi2wzFJWoKRAu4jWBtuYd5VeFR+h9iA
0zhEF1dp2gsxAJux8d6X4eklDk4ZHXPRkAH0cWt+UAhYJrzMK9cHnNsOPByjbs15
C9rD35RObubuXQ/muzYKW8p4lY70lmX9FUUjBUqDA2BIgpwU3EfjDPkQyL1sMvdM
vROTJzVUXWTg1BnZg3RD9Xlgs2PLm9WhI7JTpgMGRJ54l56GIFDpPOpRcGSiW8Cg
yP7Xt6/1dd0YeE0t/NrACRky4SdokQNiai8xCUR/90LVqVeFmxvfmvcdOB2XUCE7
tAu76Ou/IXzLDUBuNnJ2fCkVRz/9XJswuGLudzGMWVj13yC8g6hGWgPE6tdNvaCp
YUhHeD/svXJfmeDw5UlTpY+IIjCbf84H9nFgjfiviyMVb1E2dnvKBFIvk0Y/dcTP
3kq5UOgGtsJvoTD0yVMw8ua8GHvSM1Kd8kTNbBa60Djng1fliwTikdEPzBVSaAA3
QgGFGQ2mV1zhhofmzCET9iVVidQRhziZg575L4Dq84PQpKaSINlZB/UDKufo7hIf
`protect END_PROTECTED
