`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S2HbXR+sRixEB5LKu4xLVVHzkPVlVoFGy/+m0kn5SNh3kBBkzDrSx6Z8zkHvIxbf
eE3XPSRMcJOPnpaGIRCGVVVRpVTZqcTRsNPDcgO4X9COQIGWA8usuh3xm+wzNrRq
gNf5nr9orQQBl+eKAdxZNmtkva1BrGwOrReFsROCwVgY3fG06BMd6VetmMoZ9nJy
OoBWxAtb+nAZ5Uhv/DJdYCY2f8OE77OY5h3SgmgeK8onaEAkp/ZN/RGOWOG93qZu
yC8HaKO2GHjwTYCwfbWAFBRUvPWQ3znQjZaJrgde7FV4EtH/C9oBtIWTGlqJQifE
Ad/RCLU4NctLZUrDHwotqIRP+EbUGvEPSBl05UoJLI8T3OrwDt+Ix0zeYhLZNfuD
`protect END_PROTECTED
