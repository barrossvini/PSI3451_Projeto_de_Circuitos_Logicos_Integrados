`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ylsIuEGo7LbWbtOQMCG7ZfpxQUnK5FLTjJHQCx8NP7TaFsOYoBOw2ObD2IpAc2E3
M3zBNICGTLqBqp2MeZPt04YZbSGUQOZKLdv7E9Rvq5wCUQgzcdi+Y99C/H7iOFBX
NoHedCigz0s16JEJi0TIE8+1yc3paHqHgGLz0JuhgG8ofzzsXH2dYWtvYUYlEkAA
G696ao2+rD72D9E874orepAdZV6MkH38EkplBkdd+2k90EboUaGXgoMvyP1bCZnc
isjoKQ0lsA3/z/Euxb21MXrNfCCIV5MQOjGgLCoi1mUlkB6tkZQezAoCZK+tVGlh
Ccn4CIlIVQztiCFPqsVdovBWwEfcfhhA+4fFWvzm6K9IBzZs8ghWJT2NwQ5L8q+v
wHJ779sI9ejOJq/yWhWDfNOHSm4LeqH4Dfiinu3B4ZSUOk1NAwH7GhEajagZLhsr
jU1PxowANPsIuIZ8JiF3z2sFNz2GSJuJz6vuRj8MrkFgmtgdoyZ6nXNwVACrnLyG
z5s3nkKY+wbsOFgPVT74QxdchHzUfPUgWXbyZfbVOPWZuMY0y/R48a36ZWMavqEE
YXXuxk6laHGBMMUDljzEOEhA+RHnTO1QVGq5/unY6utPuwNkLaPvt2QtrzetVGwX
DWDCZvuPlvJ8asRLtzHhBpXQOvmLlSfSG7eoQc32re04HGOrWPT3r0WtYYmvGjsz
DZS9H+4wmBHKSXPl710KWJ/u+38UyqBGtGJQ5l5Bvjd+ZEvBOnojO45VjITFf2HU
uCZHaTZ1eNGGZYex9q4dCCS/gYShv49ymgCDBKxOacHR9FnDDCnBpPAUOIs0C9/8
pNg4EcHmD986Rw0HGCY4KieKxEllHKOccQpXcEWy6fEmsgVGcdZ98sCmonz34cv+
mQMNy+milP97B+rVLJk+yoEZRa0z7Nm5qirmZ3uSGrdA986yyXLVJx/cP7piPqsf
lYdl/vh9Q9CY1MDYUeixCG9K3LWW+k0plthRjCJmgUep9TtSKQMQdJCeQR8zOF0d
zSin4gJJQD0Ou1LBuxSl1Q==
`protect END_PROTECTED
