`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWvRT3zwmA7je5KIL6Gugwhw0wdU59DVXzOq46cceixjPGU/LQL8Mi9IX5IkaiaF
Z3TBRbSkZxLhhPt4SZ9PX7VD2eFNg7MbtS7OKoqc85iHYRzOecOnLm/zy0GUf4ef
gyvAmbg1kHTsd66Zk8W/YZ7rkPt29afPMTVII4Gj458guKzX05SyaQmHw5BdahCf
Etbc3cqrna4zdiDyR+yCtGJiepw2tUphP7Lbok0xNI1LND9CrcJXHRmoW6yursEZ
3DGquD/P1AUivrev1pq7uICRla0f+n4bigwiK48mImVYXLLX5ejfp3hznWAjHANG
OHuBaowku43SYHnsernoJLayorbvQX2oCJAj8ursMxGizK8jvzjcsktCSqZQqMHK
c53aw1Ai1/RRqXFdUxa5Zlg7doluKkUnWcW3ihFuduaCa6OCB/7eR46OqAPwcu3m
hF7IKuyzEMO4T+WotuSSmFTjqedYtYL03HPbZW6OLl3wW4InxJupq0uTZyB17ydA
HzFbjdgZHaX1OD2g+AQYADDacS5Pwv+mQ3k3pqKQzrusbi5tkRZMyi5g4oU3vel5
MHYZdjlxhd4CCZMN/sBkZl4x8iTyvKckMaUhS59grwfABUC90UxPzuIpALbHaiN1
Vg1PlFen6eqWHYxGk2pQ5GpznJwz6sNNZfXxDAbeb8JfPQeOQjtu6PVk338QbBGp
DePJIjPzG7pE7L1rbMOJ6gvApD7lW+yf4/tXgIUeDS463w+QhZq3CMbLifLcWhoF
08k7giaMHup1qBN1GPUNnD9dYsCeL74kmfMYhUWQPpWnR07sBWcPKIvjMNeY5M7y
qgfO4G9NANQfqLXCLh1sbUV5PG/xoDBdOX3dSPQiGdE=
`protect END_PROTECTED
