`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WXTBxBrD/ClpQGlbdv196Myf8ebY+Frfsu7OedFJzZsg7WcOaJPK9LXqLyG5YdXT
YEDNIMhZew1hSrkQKJNAiyKBOyVHtIm1wTekjQguh8B8xJPq6U+iSGJRS5vB6Y7R
3W6/U1snMOzy8NSESvDtL4UkdzYBRNIinJuDIw795EgaUEQGMvmTxnuOPGkD3xh2
5LMU3w06KpwkpNusBc/ZxxYJS1sU3H5wKbWl9C/ee6xwk3QmLsObMdYLdlJUEvi5
zOrjQL0VhKlrq0wM+kZbXkS9GOTC87yRVDuiNXlRw1CeOnURrYYbgU7qCiBibo0k
MqHAIIkympvYDZ94P763RNZo/DV2Mf6fjzAdK+4S+YlbYajFbuPPRPcflXmC0oJu
6ohE5S1QXX0SwZsEHC/SawuPd82277sb9FqTzLxCeuEiB/DKOFFhl8b9zliy9/O7
f6RIgMwNw4gCeYOIHHfyizhkm9ZMS5A22R+MICRZwGU6RCB886Q6NTgVVFmCQEFW
8bu4Alibh89Sb/h6MI+0DAypK3l/xXsLROQkl3/ukOvKWa4hhaheuRqUi7SqCo8L
ZFwbL6XPcWZoDcA3qHCsHLIMEDNaWCkrzgRNm2JHVyj9SqJjWN9g0rAr/YgP8k6/
LJfWjZilBHrtyzh2rTaaCNGAAKKhHXyph/9PXa8JbtK7R1FWzL2JaHfkBUshKzOB
Ipew0FfcmGIRL7huhl+yJBkYqSIbanmMxJz2VxDow32RkvTuRHo+sB7dqH2lGVo1
BCmcJ+uBP1SKcEV3/OykdwNNoBsOe2FzMCfDVNqlcEiBxzV5fq4HGsFUWwW0uaI4
vBWJHONvRkCmUmlbuPQwrAI0s/aN8M0GvAFRXhXmn99gbrSwI8uHifkYQ3cyikq5
e1kuNm24UEKXFmdTuQ1XYUH13laQLuj8r95UR/mqMZ66JDxZsfmIUa6WDlUVxk8a
0GaY9vULPPa1oCBD/nda7vGVlPDIU04smQ9h3INAvtgR4C/pcI0m2MiTroFN8yax
uiO+hW13d/LzDWkMAeQ0aQ6jhCt0BlDAqFLNwGKgf6oyKuDsYZc+mmERzZzCBGRc
4mWJThk11pLXr+jwP8jfIjxLmCy5P5taQNf/7+32eF/tR4SLECjch6a87t+3Tnsx
s9Qb/C/3wfam8d2ntXN4EPX1UqGMUw2u/desVqU4zIQtxVqUYUip7WeNP66rQVgU
KUKx4xfumNoXd9bA7c8xPBTjRmibWkm6LTmYTn4GZwbDN7VP7E3lnfQ4x1/4L5Bz
kEwDgvviAcL+G8uSseH6faBvraPfXrOkhxPx4D9/MGSCstK11Dw3qBxwqQvijHZU
Qse+gcEtIlNMYEOcL3OBavgVnTmuRt9LwHbgwZpSkkZ3L6S5q4ii/ghic7EU47UM
uO0XMS5l6KW2M6eOx6n6Zy5/rgncnRhd/BenkC9cXoqDX2joib1sj0BOBSEn+yRC
wV/IM8DCX9sbfMIg8qJZkmwxJMLByLlOrW7mGIf9fdGiDILanmeTUbblhb+Z+6oI
5KPp5/fOTZe/y0pLOn9oU8Kp2Da2qcMUTqv300At8DXvTPKXDquA4+UOcivPAxN0
`protect END_PROTECTED
