`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EbAVauGSaHIFJ6bLCkQZIEJvs2RBLKLPN1nU2M3waMOG6QjmD5xwFX/vy7ClnrUW
yx21iEL2GPO4qrZdUhfOUtugO01Cu1h5XypydIIXbNGGcyHY4CMc+f8iT7s6dSCj
lzJp5SeXhte09eM0RT7yIImVJuXpT1NnJFMHsf6xvS4WAqbbWrvSx/K3cG8C6YbM
O4H9NQuTJFnYMWHuepQfvp+Hxk8B7hA1TT+exe9zYdIyGCjHW4OnHiIGyxikfUeo
K8mGMyaieYCRSMXMoDVeCAoqyXnqE/bo0Ytl2Dx6ex5PzI8Bi7IK4H94Ux/Am9iA
rD7cJZZJF7hMNdomB1lhUOcnlhGUC5hZ/DnryEzbe6TRqBtScCTHRI3FzmWgzlg7
weMtuuRIu8Rfhg7vsFLeoHhzc7r5febVWCewipzwujhPOajroulddpxIuWkb1mKL
AYlOrGmd8dwBFFYqm/wEfTIZfephzlm1qmSTrX21GWfgLp/WXYnWGCjtxGj0IJZA
Jl1WKAyPstHrpd5dqJF77bWlRKzA3MC80cXeDdAPHAgfpIHvtWd8i61fr/8OJEW9
Su72nKA96um0HCJzWHSnQUkz1hcwPawxfXHo3og7tW5toAyo5cl6yYOf91FXwOZ6
C328v9GBS4g/k7ZdULGnWD8PQwFf2EsgYPUm1tK6HyInWYccFsnxKbtU12XdAimx
Vo4NLq2q3wGV7fWFkeDKLrBAVt+tbnJJv55A9/MY1MX9zuatGA9L6l3kYNsUTreS
qF8OL3UWVLKEEUXF+i2/sKkAR/BmD/Rg5HxnUAB/K8d8oZbFQIkLjaPyBXBmVcDA
iRmnwcNEVdJZN7Haad0FwwkuqW2ZHo6vkjknpMOJXalfx7PUDedUmUwuYUuvXemF
WG9LrcHyt8+9j3GfKvmVZCtGZko1NFB3t/Gf5C7If5+rCfv4FxmmG3Ehr9UMwKhd
`protect END_PROTECTED
