`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LEbc+hbHu1/JQ72lud6W+1Ac8YL7Jh59zPJrfxmUZkzJbMjx6p2qT7vSMFCwcPFd
L2GM6yarQUJGPdaRCAWaJq6wswnzQLqBcJ//aJH+2m+JhmHiXUEq9Mz1gbbrv9MK
HHyqQJbi0dWw/Cl5DUbd1MSY0vobVD13l1LVt/C6G2WOdKMMFzy+ervKmH66oOoR
PA8/U0VaMXdQv3W+ExFxnsbu73H2crLykkP+ZCqrdtTb0oyIL29zrZPIZCaLlGZs
IwWdHP2VjOVtw0WvULRpH5vGO7ZiYTtDJ0NqWClNpqtnogeZDVD6+3BkRxlgKav3
TdRs4tc7xu7iTu+UstbfQvyLieqa/NP7hE56ErKBGp7jjO6VpNAYM3TqyycVO5YS
2hu35Q+Y0gTgpXnuNzK7g/FPg10xQt59dXfl52CHfGn/gSe5+pWcd97z3doCeXIu
I2lyiPVhbnMGjfX+HosYzB3dz0pZIB7J6NQhxB8/tAmebkN5lXev7WUjn4GL4I8k
Iq8UyzLsUcjIw4TwRnQueJzMVmQhopyg+t+AZk+Eq3vzwQtETbK36KS8XQZGxYxY
jFFvUWtv6hvi+W/ddhtrDAnL13dwcVLIEUlj9yYyCGyCUqiDAsKmTzZMjkBg9AjN
ZlB6MwUZqYIq1zy7Zi4KK+qQhMy18k+hmi4YzrFLjxUAbwgZLdST8MuY1IupzFLf
Mxy32fYgJlnOo/v2XTXIkTV80mVfQbM3GMZUJc8midxv+EYhPUHSH7zR0pU1zy/W
v2YBo42L1DiGV7DAMk7gAqmOj40Z/2DlIvQn0ToXli5USN54fSYbTOKzXl544bX9
GQ8EpnPq7LPfNkYsw1TjShtoCtritFmbYAMaWp3u4MJhuqKH9SSNFXPhu+vzV8+c
hZ0a1CLFNg38XWQpTrPqInsXirtrIn+KniLCnqe1FvKWadMp2myKsp2yWvarMVpm
qZA6jwLkQXOKTuDDXP0OA20quiEVyPvNvoV38NpxevXrVClURQtzX+R1Ee6qY5LU
2mOwzYPhiIBd9k9qD40j4kLyVkdSdLrFoLoLDxT6mZChW8aO+5hiZS2aqNVG0q4u
nzEoj9h+9EtvJPyr/nJH2axxU/2v3TKWl7sf6S2lm6bXkRX3dTcnuZ11g7bVwbSy
5dIOBb6V0GUm3Q6xJFJTEOL8hNYQuYaweZlzf1scw9L9sZk4nkPfNoSaj0MlqsRE
2rXbko2eFap9/5O/kpcr6a2iHT0YAbWJ70n1rP651pIO/QbLK05mvMXYHpsirkXl
ORYlyG7/pF/A72Qd8JZzcvvxpT6xvfOKclmlJ+aaUag7v5kEkRNQXtQwfx7VcRW+
XzRj/lsmOBq0rmYeGu4J7dcjEBjP6eDEBVhcNzwjv6tzHgka7xNR3QqWMBKIMb+c
rwxlJTFWqf6cWBLhwfmr+u+fSmf1Rt5rOWqyTE/Gnqa0YTD6PELOZia1/zwiw7IH
OosoJLa/+Up3ZLrqLsZSlObllRBES3S6CxzBcKUIyAKsX83WYSpg2Kw2zY3z6wjA
UMIL5SVfSO/cKK0742Ss/n6ixY3vbbMC4nNNDIfk/EaeePmROPVUJSnquzMddoAH
FKxo1Q2HuHlh7sSMGswX7lBBNat+381bdJ+GpWB7LgazyfGzSYraLdbxMSnwa22a
ZnCRFMcnhKaGMPmlj5rtQkAPLz5LZuFRVCEM12yT04ls9bC0ynEDM4YM1wdaJfce
4wIJi+eRZvaq3sxhwkcRPRDUgcyr7ChZjKr9Hi676gxEAvKgiS0o5HC1xgB3m/i3
7RSouwtE63eEyh8Ld3A/fgmVGtGugr3+JS0YdgY5ruVO7EgUDQ3xQaZyBAlQuUN9
tfJpJWVVRPGOGNHBuOtVRteyRRbP8U75pB1QDmSwAEj4VSbOoSPfbjQWFKK7PUmV
roDvO+hngWKQpz7IQj+9shST+wk5Av2C/Gar6WO42VTeHP8Rse1+xz82YbZqrtO8
4KNN93tJjkYTW/gw2lbGCq8UaNKbkil3DodRDNlp4vAzwlGMxQHGe8wDRJXzcsgI
T6zB/0cO2Q3QaTHgLUrJ0sa9YqWE6elLzX+na4O3Hy+ySCjeMwujiGXRSz+pGbdi
WOWrRyFYZr+G0g9rCOf+/TNXAThxob5AsXAh/Fr4TbRTLpLrmtfzkoyLb/x5eoAs
p5WfftrCRkAazjzsTuOXMiL2pZs385uFm31gtuccvGKyjs2FvMAc9ZIfUP5Tt8aq
dxAaDKP/2w6qHE5D1EHqFsZxfeV1JqjTrhNf4Udr4CPAQtQr+9p/xrsJ0XWs+CJq
eXL9dg84x6tHk0NCWtbyFns1cSjAie2b2esEu7uUQaF1YiQYQTYFjlqNRKy+rAdo
XZwEikZo6SFOxiRkG+KWuTO+VBypB1zx5Lso6iuvH6+6w+a/lcJ7WFbIaCL72eNR
FKFkl81D/DJENGnZNa4JR8ydhz/Jcq+iCqR+z46ZHvh7Z+Iy9/6EF+jFC8m8DMo+
MlVLOPNpVfT3vPNECUNixLJP6gjEKMH24NPLomuehnET4lJdGyrXHMsSc8fd6Xok
BHgboHinPVxmewEmKHoVqIL4/Plnd5NcngGbBDB590emGFb9bNjHASt4Hq1Gyd0A
GNHApnapLXFy0JlffUjhoFQLPWCRRT7w+KEGUY8ZzuybaliecFDl/GKecDvBXqr7
weJwoq4Y7C7mkjjrNVL7gKQaqoZmqatmSA0YCuKA93+5HY00jtma1pG3djew11zi
H0LpY1ct1+tMmyj+DCnzYeQ2xrnIfhf7zOTnm6Lrg9tHlCVpflIMm4ki8mT0OyKJ
rZYQjo6rBG01iGU3mYmg7GpIg6XSOjUmcjT07TXBgMQe0klVYGG6h1kHx7Y42qrK
FW47Ho94chGHbuOKO4OFbv+K1axwTL8f+ivNNxx+2T0dhJOttjmU0Vb4rDFqAxpe
0qDpNFjFBB88Ti1GFKIDLvhTLhHWs4p5KGcFaf94OCzcLeeQPHpRFA1zv9tbYeaJ
IjbGQtsHg0/KOohuP3jSKLLpGNyPkQnRsvt0lKEtZZls97g6mWg5qCUtkGIGXaH0
rNpqTPyVZew0uB8pB0514ZX82e1Gml8R0/h16KeKhPIOSOOA559jENaLJB33e4YF
V+0zKphTmPqZhM4ctNuT1brfnfoJ624IHVNnxLyjJ2GdguqcarClFDXu8Zie209a
hpGplexJFKft90wiPUBbeHkOXpQViGp8xlsZRgf9pP7AnwgfDC0VDTbyyKVFFIJ+
ujxzinwv408/kkU1yS8Cxbcm3PWasw4ANMvF8MOq+CxoNR0RqmUcXLmr//xnWhHD
zTcT8v3sjsLnComyKTd91QtcMWK5wiCmfksJ/bndnNiqIH7/jBEwS3Vekz1ygcbd
PiMiZI/9bVkOrU8aLsJuuYHYmfb3VWNTn+W5hZ9GngP0uM9Z95GuGiwIOEBKV8yB
LBJ6Qk1tVhDhcCJBkIRm+FJoVaXf8HFC+xD7PinYx1y/iIDoBbbNb271fb2v0lKb
veiMbbKB5MuSr59tUy/qwLWZsOqHQqK7ac7XfrEqDo96UOmJvezL7MPRV3ntDFXv
tzTvDQhmCy2vd++KTM4roQqly+1vWhUUdG1IygG4MLtRGQ2z1SRvWFZKP/bIz6H5
ADub7gpgynuxnmkxZI/hcByAhfL3iOLUAAJG371+ZC4fJbV3Jy567GtMXwsg3jGN
yKufcaplOE2vXyNqUxwWxg==
`protect END_PROTECTED
