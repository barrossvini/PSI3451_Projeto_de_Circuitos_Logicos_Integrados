`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9QTVpEtNnzirTCv9WbD18p85H5+3oGNOEzSr9ILdmE2V7CmZWGzYYl1TveG+OhTV
HitBYXZFHfX33SnOZO1pIrll0WA9tu5eh/YW6ihEopUv/EYYkbd7HR6lf7Tl9vg/
EFOH2uQ5Cs4PUY3Yz2yuVQRyTfRUgkq9UI7jOizgfXkH4ks6V3bizr8fGgffAq3d
uGMRBJJzx3/WQaVvIXjKBc3/OiEMnNZs7NK2gBJIj0x7YLRPMXpo8Y5Jr/YVzjQE
H8R2BvoArUhrG3s7MAyf97lz7kbvZ5Soo7n+I84YasVIegBFWQr9bkhKAkjqPg5q
2qoQxqVw1pE6o8v94zPlhBXRMK1Xr3eFki6ifgZflsW/RfYQ3LLPQ5OPZXngRXer
yVY4cGR1gv8x9BsgtllQBjJAusQcRcNGsIbqu597q6fDBgGHrhMWa6b6zxo7lGvC
SrlAGeJiFLGgyFzznSSskAPAHQv4iYPNgR7AGFLhSulXAjsho0wnOfRLeXKj4qf2
lgP6PldC4iqQRVSqZAoQoOED3YWeuTgcASHtr3o+b+mNcgmxHeqnUVTGWrQRkIwx
s+IH59v8D2KzkzHFfFslLhJYO/4rwP9MmPsH9wuLLt3NJEXQaWS/BDb8xvnTOz5Q
7769nllfchqvJDuD1kSOyNnouhtPyeD8sjcZfMu07lG9MGj7i9kakCa1tsgDvCKA
59qYMjB8Sp3etbZSTuhB7uhoZzvr9UWWxbcvZPeNFhDCMnlJrzrb+Ixaspg0XCTA
XMhUBaBC3EzxMhzpQ0goTvUkp+EJM9AcrCc02EFhBzi617EJcSKttMF2FHz+Uv9j
fvpzthXU1TikFK7L5aVdvesjQKeEoPqUra8w/c9sKebhHiTHLr0jbx3bIzggkrPj
RBGqc38sgLO4XigF1qifqrdQUkLTjYahYQkI7vv4Drk=
`protect END_PROTECTED
