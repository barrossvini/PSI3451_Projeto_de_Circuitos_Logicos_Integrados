`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+VkLE7A2HF2Uf7F1YemPvoeEoj2qM5LwMj2h1uFeCVw1yjfHtD1fE/wwCdbAjkM+
LbGuYPPSVfY9qxaFJC6yNz8LGLv/Sfeyto3gR9H9XYt1fpWN9aW8DLceeRReuXAU
x1I1dYQrAKw9O44XIp+Q6cK8Wt8NqpJH2HDWDqbinuW8cGrX/Ef92bG+1z/T7/KU
TWqt6+1SGPlNbofDnu/quQNfzR8VAaiRuZfeoP/bGznaZP5tUv6YcBtsnQs9p5b4
Ame/BfIkvSsaODYbNqR83MMXYjdm1MFBd6eXwcKU1CegBHTqKDZw3QdnI70x/4e8
akIyoWiMmrrZMRMLnMPwik7czabPWAoymOiAZSOtlU7PWxsf9huNZPjDHu9yq5yb
BGTS+9TB3zppdgkWaCmAoJhmudvEbE3UIm4PGIQ+bmhh57bN3rFhTNP1Ee+WnWtd
B2RHHomDmBKGnv1POcWiKCIFbNf1GIo706/MxcER+an1/RebxF26KKViRg9A6lbD
64dywL9aC5vypiLyzd+mCFtYxmxqIaNwgtRzKEPExPVTNp9g399wlyfoFRJRQLYp
Og04hgUYGPti5ZVuTRGMaW9rqmVHKn3iFlqAR7I3rOqYr36vboZpaYF8vDoDgez4
EYq8yvZmWJzL5qjWxt9YFG5SlMxIhnRECzselfL2YW6yh0yuGq2XOjG4S4aE9XRF
M8VDFbQSxpEuYVN5x7/+z3HmjVs1iNEYj7Wyg0l894eOLB8Nrevy5480jdW1jnj6
vpwFW4jhEXPxTXEK9RkiOBeCFAQXIyN0MiZ247HNJrfQ+dk1XmuXL3vgzi3W4ymN
lVJGTVg8dTCt88SymR3bIQ==
`protect END_PROTECTED
