`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2X65gJDUvqcvcaJgEt0z4HzuzBJuCqasTEk+6bvarKdnAzwkBR0HB8iC66fYzGyo
mZ+5ZJkf9dc9xJZpAbQsm4x8+1JhDVGWm9N4h9lWgyI6OUBocyUnHnDCwtp4hjQY
4xDJ6x0t+ONBWZ88tbKznNGBGc3v84kgAZnOcA4rBX4eKTdgSgtDcSxYx5B7HyAI
u/4bVFu/EJrrFLv5fMb0y8QIC7BE7Q0GUDdrx6M+3RF7u5njzHjor9PNyMzQJzCo
7PkdK4N8nVMxoPTPQUxXEYkTP5ZNRqs/rXp5c3M7VEOuyzuAI4DetAV9tC/BSeJ+
nqMuSooig02JjX1Uk6Dozu9k/BsCO/lU23E/UTEqDt7IM6d3T6UBNPchF/cl68RV
R5Aaf8u2UctYzafghmqEmdLzS8d9oj5qnnRiuvzEly3uOmDxmizEUXx8urxvTYBB
lw82WdLAnZVxZoQujbbswLGjz9miiKbRzpJx0WmcfOqcrnNeSb8Jpp/o03chc0vL
hslurfGRSsMFfzIaQNYHH7xKK/pspvoyBj+8XXMUQCtDhMMxl6I0bbiUfCz3VDhv
+GDySm6cDzg4623aTxWVssKHxrztqXKlMwHkfAyEtHHvfxFJjbUsYMW2WEvi3AVw
Izi/o00j9wrqRJtme0Pfj41SsKpEcfIqyDAMs1UraOrpJgVbsW3FZnYfOc8Qw0Yy
HD5uuaCpBjj0ZZ1lW42c+yG3Z+YZKWTPai637j+BBjx9SxU9+dx4V3s3OTCq52Ro
yzHBUeUxE/xAlybdV8xnV8fKktM+GSp8sFUYjhqS55jKSGLTecFD5dYkH8p26t5T
tRc18s681ZAnqnLYKoq9PXtQT6BHgXtQOU67P1kOGW2PXwoqoPE1SVuUGpbsR/Ik
5QSWBHJpNdrYXRzDI7uEUaWE/fN1NwSGwdq05QnGhDzDliMa3MBviBODy10TMXsn
+KpAy7ZU9qyRVvTWmP4XgkmTZ+wnLI3jmVxOY+QVrZVnmZ0jzhX9rM8a+SUZuy+3
vcNryqETwdQypbZvWwcIWA==
`protect END_PROTECTED
