`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WEBNOFi1q9eIE4tB//0vfbIR1I5MkoMpbB4+zLS2PmSrXZFQtL18BIO0L3SpFfKl
87hJMpiLidMc0Da0btU2aIlCQmJW8gEBQJaUeGwuinwg64tmSUYhRoyzCUsOiEFU
QLj5tT2IESNE/r+amIczpt//Mfj4No+jMRsCx2uQgNz2btyzW1byZl6F7l8YNMrf
dU3vF+ZQeIPOEydeUig9Vy/6GZBLRJYv5yfs1wkCFOMIot+M9mP1aA84VZb2IreP
onBkU9LGp7sozgO2NoKiG/d0MfQ6MVxGrQQSAP//t8xJpVBjIbVYRPZCj4+GpI4R
CL1x1Bxr7ZFNQN6LBMEkOaO3wQp+FA8CmiO4RacwxSzoOPnZ41xYZ6FtstlTTtGl
GNgMo3+kgZSsTaEoLwItBCeE9PVzzF+7Tomqwz3LbXtjoGRWOVWy+GsEXrfLHkEO
M/N3x32xvxwbMEASj7KmvmwYPVSy3eXmGzZjQENVXzmEBqb73afBU5QK5fgSQrd5
NIeAvWLVcrcvCMJAd6VLToafviPhypEi+ma5Mv63seX8yiiDIQGnVT87KfldS6tl
Yvk4uG2QA+qN/rizQ0pu2fv80Ir4Nqw+YoiuUCEo76h5xwOYihACrzOdIK6qRBLX
iSBhYF4tVyK/OharLFEpGAT7uoON473fybDt3AvunESHUbf7hqFc5s+aYI25kpbW
AS3oI+yf5JBc6Qh6ExtecmKAMfaDLy2vxnYFsYuuKp84o25uDOTzSFfU04KYJV9E
vENSlCMXk8HhVXzhtecNX6GviYfnpEquUwN7BvtN4eE/2OLoxTCxhDmDfg4Gb5ro
`protect END_PROTECTED
