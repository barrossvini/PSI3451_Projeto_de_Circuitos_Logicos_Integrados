`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EOq+UiFBjWa8BfarM5q5a3mJu4rJiOE64aEuvy5In9snj6GyDh4m7FBgs2t9tomT
gXTXkRCw7bC1A3t3LNhRk/eRgVIdYb8iDhCAADIig+Nvrrg3G953VRUDl+omzNzI
b3hAkl0E1wJDQ1PUPpDoW4AV2ONag4LGJH17XHm3WDu/qJ+4ApFFp3W+wIpI1Ou/
Vd8Gwqne/oSPsLdydZhF2o3kICLmLgj0jWemPyNiEsEI3p61ZBwaN+5l5ekcTMw6
V1+kMh0dUxPoTdNPdHEEzaUdTpM9UhLYRlTfn93Nfzmbq/hNZsSMz42caoaAcAtS
qKN5MNEvq2QOjY7E73VnN61mgLP0WwebMBmsGQE/VvnYGIyi7DBRIHQjTrmGl+9u
4UqU943iCLnxbXw0fvsCzMUWv3s+cCMHr6O1dwo2YQ/I+IWXfrH3/h3+MizGUuKP
NeWrrEnTk3z5/jhx16FGikJAmNVQbeYk8EOTaK3wNJsmHOdN7Q2SLOVf2AyFOXz5
9a67zb7xtd3aSxpZICND406SwkOAz7NleTmdbuf6xpD7MQp70zJBASy7nGkB6IL4
tjvZeC5fbJyvfIv+lUQKwyeamf0gkY0Fu7Itgya3GB+1BezqF/sAI0moH7hR7AWb
m/mjsGEdwDW3TNIy6fa2E0U+eOsZ/faz2sVJl83MeeZppAOpvlDBErH0I/1yQK4f
z84rbb0NcJ8Zz6dyArOQgvIB6dKTpXH/Vye9iHPTlFva9CMbd8hzsn+8ErnV4YQq
5Czp+DxZG0K/aC2hKfytTjrKCET+7gNKDIICWcAMQibLIvDNEhcvR/7S46NY6uy7
xBE7mQT+7vwKBGws6WNRUc17QCGNIsolNyRLpBdf0LA9b+g+am1buVD42o5x+8ZJ
`protect END_PROTECTED
