`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n8DYv3SNDH0rv6vN4ICpA/QBHFcUt89FfJTR9VaPPMj8cE7swlZQa+Ti9I/1V9ZQ
gB/XJQm8Hs3LCszzG30+YTKPOdyV1ip8t6uTlugFzt4u6DIADn7r7LuPbkl61aWg
yOoxyX9l/Kcx7756Ld9d3wNkkl5YJ66u9X7TJQuYqYdyyoKZhmGLwcuxSc5TJmy5
hqs8QE0fbSUesowQuDoi9Ej9LFtZky0G/FnMDLuLsIbrpNTwYzOOxvaSfjQmWX2v
kaMEW9WDbVsvKM/5/NUbZx56OU134wvGa/pE3+GKrPjZqYU2nHo7yco1AqwwG1Ql
dRMzb41WDgg7ccujB5pxoJAarm5LTuC4QiKRZaMHqvgtM/hSIPangs+69xqpB9Fp
GyxM7pGt6RVH+aki6OtRVEiKWs/uLZG6V16ZL8CAaSyOtgd/vWmQJPnhowvsvZTc
8aD76RazFQZP/dmRJozCqXko+TGKJiKAaG0/MA4flDCZTTP2TgLGy7u66Bm7VQHn
YUTZcpnzFt8Qg4nX2uIC01j4NOVTgWLl0Pss9dEcG9VUB+WDiPwWxLpLfVO+OVYC
32ExFRUhtekxQqCGAbRLvz0WTbcgD9b86D0CD1i09k9N4lA1CqIcd+FuEJcfeshE
VSN/hXnQse9tvG5QAvO/gLHChjL1LyWMATPm/5ACvSdgNYGjctxJyOkUxp0tUnVY
`protect END_PROTECTED
