`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cwrc5Vwv7S8FaTiwecSuAQQC5zuYaKg8xz4pJaK49KiRTrua4vW4usiyGI+wW7gi
IQzwUkO1C9c9ih2sedh/vnbSXFQa3/OhTL8iKWkN/2o29mSITXcoOoq68b9JXvYb
vBcZKg+UOWL6hubWrJV+lKN+zIK1gqByaRER8Cdo/W1X4979UJsW6c1hZPC6qFdz
O0j1IqRxihECWSmXAr9+c+ziqoLYIAfosoyamMYvaztcPXIdSWyFbI/k/qmiKce/
7pqguiRVZiKNpc31s+9lwZ442Xh8epq0+ljqfNSWVe1wcpjiHo1FKYoSBQptuU2C
VsnxT3Xe9qcXaD57tPZD6oxeYuTVt/A1oWIPMYfh6LiClqVdY1lw2NK+c2JRVH9B
Q4LjKsm2KjWdJIAng5RbPD/lfoZASTLJzh5tGHbLLVt0v8dOoIkfqw6U/doSifYb
8GwopLxirpjlSe4vUyAGXsSBI+91lMkomM5auXSE2U+K2O0iDj7qMm5ohYS3Jgtb
DAY7uLiMK9C0ublTfSgZ1/maT71cKtuoKxaNsU25GRU0ev9aeJzQJ+ZuJPvje4bm
aKPic+pfrmWSftJUXavIiDNZoMqn9/Oy4BzjGX4giUvk/a/45uHeh9BAcZaSuWDv
x4yVpbkPIGRWbcVudiXO1WHpHn3fH5KUYJ3dVXCTiUUoEVRxg1ttaRw6w7lKSd+E
1tlcdrqKuhWt/VA43NUAGOOCYOT3PPPIbxmJCs0fi56XT5CEIkYdryYGUsyU/XJa
0OPl4Q+A9ipnqfcE1t8nwgBOls8sl+5RPpgJQfVmaF97PVTuNezJjrRK3hSl7QrJ
gV89qeyNtYRQeKHu4wDqSLHTW1aH+0HVT+IiGZPkq5plmPMJO/P2EnVkhT06GbdH
79wPskqxRSbPUFd3Jg7WqA8xeOklX0No5mthSWkPJo+jB8S6wh/zV/l9WNghp875
/zMx2c71lP9/ytyp/0fjcpSwEr3g296sUKv01TRE+H7ZBiipML6Cu1oOd7EEbowE
DZYZ7GXbwEJBxHKNq2Y+6mTpFoBWfwELR6/gTyyFt9c5Yuytd3Vq1eeDEwFL5iPX
yuQzLhYhLPXXtgGSE1UKq0ohXVJ/9L8LyYCNZwplP8Wys7d/y3Egt4JKi0caCuQU
jTK1cj2Xi2mOLrdD7w79b4zdTdqC2xkcBnbsSIBLK1O1lDvFPr3mWOylXNNvqRmZ
5xbzg6bCmDXp6W7qlgEGq/R3RZfebAUW494g0czKmQcjpLNSuC4oYo7QcORpswuh
WlgbXZPj3yqzcCeWjmrWkBU92+rv1Kuv2ffOjscJCNRz6YZmofn1LM8rm6S6lFNe
OYb8/DuLakpun714Ey6TLkFlJtHM72YR2louUIHryh0L1UpNCrBDfPXYJbjryBHl
WhZLmuUF+GyTtpwUCewpqKovipOS68j1OVNc74cOlnxQwhXTj3TktLPQ1hS7NcRz
ntxwWOP+QkhBaWV7dI4ExXEymVrj0anz5AddKWUk9yTZEdbwJVZ0Y7dWE8tMT+vz
+vL0BXozCmighrFEd+x890hDPqRFe44b/QvKOQVQ4NImozqgfa3TmmT6bwoB459v
HSy73FaFajemh/JB53gO9CRE+nXTHIG3Ngtp3p9bspGhJWuCZaZk/B7s5NEDDyQd
m5Fsi4ZAM44iDc7Nv9zfu2f79DIM4Tovw+1MI4C3HEdka+5dJwWNY9hFqA6OFeFu
mFC24uzUS7ALIcTKl7kXOnwEoh6VfZMs3Xqq94mK2DPPWy3ofKaSn2VXxpkVssj9
MmzF/qqvEcf5D2fDHlZ21drcWGk3/KfFqs6DaJcA43WZVERnnRV/UwUn4cFFjaOR
BFdUluPRYkyeWrxEeZX3+eAFETCJkFRT89mUxrVDZCVka0x4iDccmezeF4N9NqBd
xsMlpCsBTcdGG/FyCa5zxzE6jghNlPB5kblcDV8d4ZVGzBvfGvscS/UvMTrE86Rq
LFuudL9jmeqRm4+Zu+8ITdr/sAMPbWy4lLnYT3JV1x3wCzdLjHJU94lpGYQDkuEe
TkfNdsgyPVPzp4NyVGcGvlXp8WwiIWtsY0MrBHQQJdXma38lkYviNysnbVlm9rTo
8W+WDMxK+FPCbBlH8525yZ4jdyXYQ2F6f/n1EZ4jGjJFp1jgRCAHx8Dzh3zi85fL
jgc/5czeo187UPSMzs5faGISkgy3cshQTybv1THTOmZ2RKKZUsP1fMmdXQIdld3K
YBak5WnKIUO9OQALunBk/dbmZC5TtiStP4bv2Wgt3VZBa/uLe2seXcFDsXHucjJ4
3ZxwoTxl6sMXBkykDrQxfywjXJpFyOGqc0+KfTlE6xHZvMwVu8ELA/6EwZKvAold
xrQKT2RDm35SBjG0jyOUcQgLl7pS0WmAk3fDUB+/gANGbawlMMESPmMIsKrGJigr
otvN/+ym824rvSHqEvV0ZbvIVOvw0yp10KJ45aUll1igC4lmHsqlUaW9mXmh55IC
bewaezPDdrJzinzIg695ihAkcJ3xxF3tYDySaB3CXNoJkdY728o097IaCOnKAdY4
Brqd4TUaaCezKF6XX/2XA5giTHCmkT5rZ+TgQGqbQVBDkP84v8kmCiolqqaI8MFp
iWD7w2IWqNyyatBTB5tZY2K29ILObHLAyNiQdWDHtuIZmNom3PU6kKxtZj03ASkk
uqlIwRPl0IRFBRg6wVcIjgs4gwrobRamslucJLRmNGRPFkh8FwBGFvA6sEU/neIz
yhy8pbTHhs4TBmhas5yUR5TaST4bFCR3DcH54w7cds5Kx6xx+K/Em+br9Xae4w+S
RDhcYaZnS8Cvps4vpb3qmUEz2U8s4/z8jliC6gqxOjP5FU1drOQzej9EvE0ialTA
PW8EAVzcJ9G7dEws5Hym6i2+JzidBMEbo/9ySfpa1AXnvjvNqFsd0Hg1UR/sCO+S
E+w2SsNrn+QbHRJRMNJqT2lgDudlaWYnbLfE/sjaWlK0UCT/su5HBkE0MhRJJRvj
+M2yKw1KH1whuG2HVqSYDoL9qXlQJkkBdou21h9JkzR2rBYtLY/cMzvzFbADDO71
OBqbhL8CMTpXk3M9oPXBPsLwhtn3dmq+CmBHTNCjJ3UdSuJdJCtdyAXJSqUJ/X1u
C5xLjyVWJyKkJXrCYeiUHoZacphtH9o37gIZMsA9UlAUa6HnFZQ6+wFn+EKaY4q5
pnnoqM/2XUTq2hpw+FzAxAkgJlGSezNB3ROA7GEz1cC6xQbpoJulZgJzaRmjOpiF
EWzMFk9kgQbNmztuC24GdKynY90sL8omkEQYvBHkDGQLX23KJdcweWBtx+m8Iy6j
ojrPv0P25dnrTSeQhsrKuxWoO8ljEJO6Y5uKV8zXEZrc1AwxSdVaRynqgfDjbeJI
u9I2C//bO9LJNsQnuc58fCdPGxkCMD1FOWlIvMashNUTmJkZpqj1KUNyOvSnrxSW
j7j29AUkfMdw4GxvEf5S7O6NAJH0yM5YxI/yYAkDHlmmkMVPSOWzjF+rgJDHm5Cz
tnwIdQEKBJzPmJ7FZLMrBhJXu0Do2iz0vswLXpU/7SaP+Ihre/uxfSLN/Cnk7Pi3
K+X6OiZXWhlhG3YKiUgYDu2A2kBJPVsfKPvcTZLV/53LEjXzLjUgB2GHAd+/7Hhc
FbiDQW1Ers1VYiI1iYQa/5xUNy6T0C/FtpwOY7Z+3e/wFIoMgYurEwKtk3yTFrx0
EXkEIOJj9C2UKUf86QfTYAXHziDmLtM8Xp0uceZUD23tsaFfgfPJbyDgp3S7JTeD
J01pDs7TJ4ObuOo9jHDoOP5MEfgmQ1ddv+6HoQIPOCdU2SB8S7hMAlUgwvsOfIot
642WFE+tKv2iIzXcWUfzoqSb4WRS8PojGUa5wXIVmUXtZwqqVUXArbW7PFRjKcTh
sCxh2/W+g72XhsG7rAMD88VOHJqnMIRLa7PVsk17igFzhNpTqXvCNNL/LF4FQ3Kr
HtSDly3V8BezfcrH/9DQ0t8DePsn3rWT8aFUTCitbTaB7/FES21JiI401tff1wbz
2EGsiIM247NzHpCM8O2JKvPZSaTv7SUTbVLANq5hYRngkCPnDDaAXsYPbtpkrvuB
4OPrMBtcT43LXFj5uiAbtozoBGpUqExYL0MTkARUeoj6p1yPDEgjYrTRG4lGteB3
gss5XRSJy6pzhLf9TQGGM8EjkdWiFU7fuX73x6kuutpy8b+u20acREeSw6SkzIul
Hz+/o9E8o0mq41NV3dF0Gwlh0v/ULC7OHWnnsTvz1bt6FlSTCBlpwv7CeYKRNAeP
hFXNTgEf/AQ3db7m2bJagjP2CuYjfFgwzCkbs3GIefXOER6MHl92KZjCi34osr8T
/HEn2nbpxoCPN731Y0qPB4DW83sxnpikoRgO9XgaXImhzmSDwHxOD2m8lW6ax6gj
rezUdN0kIssYe0k7nMvo9YkLBUl67LLVmFLQiqU0Zba4/AVwZ+oqixw0jYF+7eM5
wWhba9/MbmJE+GwPECAaMwRkiYwW95go3duWzB4kibp+JrJxEjiiCbTb41ozyAmw
9IwjHVB7O5zGxw223rzIVtDIZmPNCckivp6krwNhaqrJJaXPawZ3irJs7xfVWCsn
g1UePz1PM1OFw00fZll2yfuXo3U9OF4QL84eHu8q3bQ9PqJyoZ7qoN7JL6duvw+B
n3iXnPalnZkYrk54v0WD66q/f96eFj1iLl991RXqW4WmDG3ngrVvFvIgvdk6mg3x
ehe/VATMCo0FCiuJBu2TdJm+YQrxNjfU8nXBZ2djZ6TPP1mkGWuQpB+k6N761kuZ
9MiRsF/gl8eMFjTM6TCzv/3Dm1Pg+kcV0KwDd9S7UWXDqJCpDmFDFwKfigCluenY
KA4xdRQg4anx83bKEZ4nC7ohtGOOYzB1s/RQWXETxxl7/+y9zLeV0uohe6Fa1KTe
HXUJQxEwspSKf1lCipaWeB5lryKvKfRjC1GtMc+cN66JVN3GQA5eY4D+XeuAEZcT
P1QwXqbVLmjukQwmYmEruLretZDU2X3ydbd0bEjCOasj8h3a3xwvC2Z2ta5j5Pgl
nXdKDi4CbJure84UBncxMQvm6rJBmm1iV45XbsOruF5xW7r8c1S/Y/rBc/YTWj4V
I4l9fWg5FwRwoJfpznrQVzysKeVeLhza/9U90BS0spU7ahm0RMYJpuUSrCRqZrKJ
Kf9TYJljSoX2uIYXoa9POEfrw0N1MhVB9TvrECVYY3/IAa/KCRC/+8BcCj0t65Vi
SCwQzCewZciwj6lk8tHG7qJ/ZZsera7MdEny4qtlvg4H6cRhXklEKIfop2OVCuFB
E8HGXCh2PFUUU50QkTY8DUL58C/67X7Ke3mO5TA+KuCditj8R7UFv/sAX62wc+dk
oIYAAzoxoxnYXkWTRytCbHJ7RgOI4WTdtlZgApww5czaOUIPCRGmlCy/6YKGjNdr
FyS/neNcPYFlnCgBEVZIp5SBdqLaVfsMpLPgLo5yV52P/SJevDYw76Oj7H9NOLW6
hMLViJK8oQrijlqHHsGULqxYTHrcT0y+HLhad/zxUmAVe2ldFZ3NF3owEvrL44+f
2fQLwhM991jsnsul081/yLfQ4wPNBomY6MsKqx9CaAQafViK7NHIkfZVMJ4XNvDH
FAqKfnU5AxQXsJZWte7XVNembiEIpqDKtweufhd9VOyaiz6a2qJEnwq1P/7OJaQz
K+YwxSACTiV4cU2HwRSQTIXgbFVDNDn5IsLqLrnNx1NISPqQ0S5BVJlBkmT+Mxxx
fH/M49v1zw/Yu7kLDo5TSAmZNQIGNJj/wa/UuE/BFgZgoAhqb4GgxKLEVms4CUP0
4vUf29JyIXg96ZsKROKPY5/hKzIcGwlCDev5B6aQhoyF5TIaJRJlZSlHHeLovGoC
N3khymsKvqGklOfptZpa/8Gv/2zSVBfg9YkJvjFVvG6UcRB1Y3RBQ4KlcXWEMu3k
+7SkatUz7MdFD4El4alJqcgtwec9UXKxQfY6A06Kr0LX73AM0C9OdwyAe3QX6oyd
sOEoI/V2dzISMdw5iZuM7jZzr5YrdwXRiHDnvusUTkCGsIhMkP9aaFu+03Lh0Zxq
jT2pmZpMi5ib0/DGH+G13dQe6FT/eOrsVlfP7Mux4m+9UZINgAiB6UhAADU0QXLK
3QeH0lGKjqeyC0Pgc+8Na7B740MGzARJhK0kP7VCJtjofhnF1pyBlEz63l8lRmcR
mtRIChQxExewVgA/dQdxone3hTA/oXqNnY+0fspKLhpusUVo0Y3aQFgAREvVNmrU
4LwfJMsbE/GtZhO4WLoqIoQS3d6q6P0xFUcBqXWyvGFuUnwkC8+Q0PllmRTwdLsS
bphy0NV56GvSN21fUu0jp+7wZAHNTx+f8O82iJv+B4vQA97q4CKn3g9nQzWKjMke
uOywzYEw4YzCG7lzbpM8Vz1Say+bZkiVOjEY899oEttYDHDad7Qf+gB3CJ8SGJn6
IFPT6cn8uYlN7lLp1fiswv1+AV8BheBnHAmg9jGNnu+Zikz+ZkdWUyZ2qI8A4gTD
RRVVafTpaTbN4EWJ5OMUoitZtNrebuRk/FZyS1yMOwdMm76sFVqpx9v9RxkWEuno
tkh7MLbjIHwziqgwY7RGMPUa/auoObB63IryGXDSi55KTUYhaNkEelaC3NeFDQS6
vKjZpfEG0Y+DscO2GashqqRuBmATgtBCOMQUok6Rf6BJIXJHD5TOJvFHpJnZTjS+
O+GIyyKLmQOd1WJsxi7f1+2K8N3kLpXg09Gp6nOc0mIvv3wP3rUUdf46LDCbHUaQ
18zICJlCAucUq6/nuYgltGZzXiIjLYTVbyNn6NHRPnTp/EfJXZJcVMZWOo7dr7Lr
EOAEadpIr4SR10rrkc3NUnmCzWb+aLs4CQRN1pAebfn5gpOfqlO5rQn5nCIFp7ZZ
X8SFIRorbOmcIcuFFsI3TszLxIhr3+0Nqn8zl/75QdjO/sI335NuvV5yGg7NWAJZ
SZFwkAfYyW6RUCVVkVzu4IaAj5QDOkmrnOg7nXaFGil5/l3K00vrGoP8zCiJv4dv
HlPmJsPc96LnbaaYFLc9e2kzHnt8LoLl5RaqJjddABTy5FasZSHqjfAf0B0++cYF
7fZhp03198Wr8wyRHSWQAhpd6M0IMuwV0MxMR/LhSb/RMhPBMOfKsI60w7yIkUFf
NF5LUEup4dl4GlUDPDY2GSHaaGhEYY0UYsK5GU9keLloOKWHCsmazWLii+WJPM1y
3fAc6n/QMR9nn+BdeXTZbS+nC2mPIbgzhpnAk4yJwqvgxieVcsLWPnVFvzvexAWg
0ESIjbj/WKQR8bPHxa2wXDfu/nac7gOO4vkA1Wz8zWEu6J/ZjDcvXxG0pET7sn2B
Hu2by3sCJi5j7F/1dqBSOgeTBw93QEf8YPO4d/P4rZQaHgYzri3IuXAVGBm7aAFc
JJKP4fzg/tuIHyoRWZ5b7a2HB7X+bWVoGPp1q2kDwtkLs1jDNz86LPWYHKW81JrU
Wzvdiv+ZFwdeqK4tDbJaYHwji8YGV3hb5adeTMMNS6tbwPxY8UoOvGASLGxK/09/
NO6J6ZYwQay1JVjeXKluD2lw9kTxBIlktLEHfz0yUpSWAEH3sYXt3WyPkftGXsUm
8vHndFs6gLgbYALlOW19kQTH4/KBuRR2LOsjvGBNFbETeuNpYTIJHw82jJXSPyGq
RdBQC/kXXLYirbxg+HATNSvwzwdy2jSEX4UwvXyG7dnuC08B7Z4fEypXVHeDM/Dg
E6BSq/QJt+dOgyGmXdioUuHxjK4dSzFhUnR5JpGzywvwhNmHhfplyv41AaFHdW7y
/yPUVQcpt1yHfhVsNFLnFNpohJC+XmVLS6ahoKev0Ej6D/O+j2FuT9pskhuduywO
UIU4n8SavmEkQ1q918Riya3pjwkju9eN3pvv5PlqgVhAgSha7kgb+XcWIRjYJani
PaJQvxBbz3HsV5Lq2pK76HJbjJmeEcGHbcpAgv078+8mW3fRYEkzg1da3WD1KIGL
W+lyWh3+vgdxgCpvzG5lNOcU8HgmIbVHTnJyfcC1rpdhJ5DQDWjLnh08e521xXpv
VdwLKD31a2hqW5XKsmpVB1n4TQh5pByf1MmOO+LJoPnkx0qIzhwd5lhT5n9jeRvJ
7jS9MH8Lzr9R0npdmx5p5GNYZkvauwjch9RyUsF2peaGWM5OPb6unryOhGU3wqZt
R0BI8A1D/EhSjWownjZKHMe3TDHbb2tiQHOkNRHpu1t1IObiwbgV9hRbRgiMbf2Z
2Fu13oRBdocdwV4QrpsQX1utUMc1w+w2lnTeo3gt58P6TpK9St8xNHyekqiZFa2R
yb36TRLdVg1+LDhXleegV8JoA01RYVESTes7CK3f3tmOzOkDgh+T1BP96o2BuCTa
+qX5izvFUn37EqlAvQgL4X3sh3qxdTp51F4lyXLKUaRMsgXTTxh2bv20jAbf9Czv
YNpxFAQKrNBsBShnn/b3p8c+HTH4gbbzlRPvBz9HdPN1qrXJ7pEFUhoay1erCiSm
5BQCeYGlC7omDMbLIq+dHpZNEHmaHN7s2HdVBVp+c1cSRPz4jIbyOA/jaLRFcsd6
0d1zhAKRUw409kGXBORY90Wh8HcxrbNK9UZCOMduFmOg380jBKMA5ybxDHur0JK7
BqagXq24iSQojQVbe0JlOA1Kmc1+8O/jKXxAjwET4fnlwn+NfViIUzoeGsdn08nX
TZJIlKfPgv3+10Q4ZH5G6GnHJExW3YlqeiwdhlyI9YlUIP2AN+06y4scr5NmlvJj
UL1UGAcadZwjr4ndDEKvBlLGf0IRzVcb3C5OUJmYuZJBfMxzuWMtsnaauOoUcy9h
P1ikRRfmtrryQPF+xQEXIsjVlopkz1kKmaTPz9ciFlp7Pq9lAY6vNRXr9vxw+zll
NOBs4TVWLEwHhu4OZw8KkKAPb4ItPhIUAfA2IObF2MB5+nVsd3UEHC4xjXqDLvvl
vUnB/8d0NuBom4kgFUBMkQ1jyrpxq7MqFvEdwqljWxQNkV6GYIHsdryh5s56IMvz
rIjQNlWCPLkb0Ds4ox2pNphG8dE37b0fwI2fHNVhYeNwItrI4wxVCvtRGDZu0+Ho
3y+9e8+KXi9MVjKXGzqTnBRS5eZVdjrZjrBvHU0uQuvV9dXL8Ay4EEUXo0Kru0uY
b6OyF99yah5lxBJWpe1SRiOS3AT7+tu/Y8uDyxl9IJQPW+ChA0L6WHQNO8sr6XRZ
BBUEVuhU61QYEuKlFU9ELbLjBoJu8vdhuhTncM02DSr8vTlCS9ZCZyQRbPjSggsj
WoFTeEaTLOBdMWBvYkZQK27tyPeKqXMyR1NcL9E8DBWQ1bKZuwp8GhMIcpoKCtun
+FdmEPd8lV3QqiRByZzJY9YfF39lbvNVKBgv8Cq03hNO6OWbYxMHmXnOkAL2uu09
lxhJrAeAGUU5R48VZE3OOVTNgVRaHy9g540hHj8GWX0F+LKjz4cRZb0one0U4s8C
Pzaj6EYnlfI8m6KHinVinWsCjeAUS+gnzBrfMl9tUarlIvRNR73n2WA6Z+vc/fV4
ieSiXDQrNpww/Ur+Hl0uxyAy5RvXoEfcQQXa6sECYPLo086wG2Y/ygQOx0q8sYtr
peuqbyM5oSgL9UxGks8Z76WrSNRnhyYQe1io/ZDxlkFC+OZVaiJdTUkwQmBPQLE0
XO/2fquTMZkuqtjt8WOJJHO9YU0i7vn/dHEBhJ2LmZSRKjZNN0TrKZUkR58NdEpu
vLmCHJvfn9afEBXGp98VfwtvkYFAR+Y8IfqtH+nXWDgloR9o8KgA3UJIeHPqR52r
CV9ivg9GYvp4LrqV+pt3pNgTej2SwieqPNOviOEB8iNN3IB7l9pLqeWXuF1WcnQb
atGJOoem7j9UcRO6RcG35a5F7R2TsmhVZaKlCVp5+nCH+/4/3DSCsi3Z7ADRgXA5
IINb+efJdbhGo9tMj/WbBQmbc6bysdrtemH8YLwRcrqJKH9mANdGUS5O2Fp1JnOS
WpbBgP3EbFgUxwF3WvzYU0lsbzhCoqzXvLgZSIOak+36GXptGi6IPEuTOKq1tcVr
RKQcHI6bGVHVJ6v58b6Oaz9mGY2TbvtWk4tNZb0WopYG96ipjLP0YIiDqxIDBdoo
r0LfNxDf6BbO/ybwowGgcg4MC63mUMGwhTdKIsRyqvp6vgJX8byHuVq5mr9ujCyZ
cAB4CMyQqeZF5GeKfHlyQiKftIXS6pdDf+9b+bqQyv9sfpGG8XyD9QX3wbhY5or/
vEb+CbMReOB7ZqIr7MlRYVDU7WNGUBUYokiPKfT1vHz4MzbuWmu1QnIA14RuCNRG
Dc7XC7HYFk4d/i1/XqrTvLkPkbrY3LWpLT+tgQRg0NzQPdoPtdu+d4eAlROCowj9
w8J8r2rZtmS9P8DUsQEy4kmZXQrnJRyW2U8Y0pIJHwxGXcMliYqw9D5rZXbvSQi1
KTF6sNzGrxorvovniGmg7ntaEH2xi1hyOerOWZWZv70Ms26xw/LmLh2/dOeYyMUd
oCDcqdwF4n+nd+nle+iPkvtoQXBQF28WL0EK7njXOYHAVv1ptI06TEZO0W6s09wa
H8Au3t71oYjrS31kFO6hrZ3ND6GUvbEhaBVPxBIsVaFDaMY0o7EkRii1F1x901vP
es5BE9izZkTcRQWDwGUTI315MT9zDT2oExTkVRY33EAGLyrLUPicvVnm7hTKfXmK
YcFqaEeE+tdI3pAaLuKWDs2WvAOVUAAp2pwHt+UdiBwk960brPsPxDFWK1x1kj2+
1XWtkiYn/K0VckCZpi1unje7/Mn7V2dNSWwbjVsyrSZfRpB5151wyoPi2KMgMr2Q
JukFvdgo1LG+Kd9sqRpzI829uJ3hwsU5t9nhZ5Ej6FDLz3i+U70Iki0B1bymo2jS
ojzdZqDD4YWo5UpOHzQYq2EZKwk3anebeJ6GWWEeiBOFPPSAfncK2wtzazztyfHN
wMpYYEbu9HYbdfnARqPQtEHF5SkocWN09QSOhwLigzwEHDgGNVsDDLu50+vgoGT7
oEzU+HvryQ8MxEN/Tp50bQvKupRf2upYxR3PNn5QJ/DY8/5STAk0AjR2V1bnShp2
XUXtAGQaQoPBNPj63XfoouxDUzkov/H0Z0ZIZJXNLHaV0VDlTIL4e2UH7XzQVt8P
0CipptUZNc39MuVTDNnlrzlQbOGerIewnN0xsLQB3lBTfJaa1PGAJl/vl5wLDdVD
550mq8NP2Z2IIUwR8dFqi4oJ4BqljJzJM2wLD+AfMZsBNsv14xPLiLJYOIMM0H+G
1U+Q7K5JbALjsRnp6vN+iPz9T3J+/R17h944f9FGGPlg35Dr9A6Eb4KvysNevtdU
s7xS/1HrB8uHjQJV7gkHclq9GRt9XROWDvgGEeU1myQ0PgN9Lvgkwa5Ji+PjNJqU
oGZccomt5HletZI980zNhvV046YZTCHZFSh0u4AKz1DBhMhKUL3Vf18dbZlfzAA4
49DQmd2rFxX6M36S60oqurd7goOwDs6TWpeY+uEAa/D98pERRos9O8CmmFJa7Jbc
bynA4BUpsDyTjEu9jVVXt2tTpzEIRrRWiAucSONL0Zg+HYe8ctYUxileaN1bOLTe
l+z1S22JZ+jDxUSwAP8V8HaEtSlN59JAvaWwdMwY5fZCzq6hRUUZEKhsrPFZ8W1D
rvFPSofLJzZzF82WNXz6CJuY13TazdHdZmssCG2w4kEjMnnFFh3LPzu89F5a6AOl
hVi6CminEKCfVpl3/2ns9wnSP8H7XwVGervS3lSni78f/tgHLWtpHAWtYCgrdSfh
JRWzpe1V3az8AuKppYkUKJ3XBX9WfKM/zcqzewaTHnNcwQbvTVQicJxynarm2GM9
9p33xcJd/vDIGtJfc0H/nMl3pIOlADUziEXotaebRGH6bUGmqpc0VHRBs4ahABIP
330PAhyUtsfEsownLKvrR9qb14uF3iLVuyX/+MfmjGx/eiKETF1rNQAR9H6/Ykqj
A3GeobXCCf8qbX2guS9c6FZKi8jrM2nbFQ1jB8zkardphuqnwtaq9hJpdgeptLg/
rK8cKJbj29fLzeUf9O8g3Q+9uwSdVzPDb2d7CCvGR1Lq6LgzoJobvHeI4O2FZ+9n
0z6HRiHeb6Vw5lj4KorXm2HnwTNcTyfDSZD5kKM6d+UVpWBNNCjTIzjdOKOjv5zZ
Cp6PvhU8eGPQ3IMx8e9X5S+1QcHHaEqjYlft7DRU0ZVcyv/PaaCpao2cItV9S9qC
zzAKmFJkURYrZkuJRVHs3FxkY9d/wmU8vFcOc/7ENtuMWxwLvJ0rrwnYczOnHZCF
R+BsyWNbKl3Uyu9a/nDdDhGUHPq/1+Iuxoo7M2QKXCBnx2hbpzmwUO2/0UhbNApF
M4vzZ0e+WJC2X6zl8sKaISKevxRYRbPu8OO8Gj3NV2KZT3QXNROADApGcpRnFamq
UCc/unm8x6vzIv2DAvc84BULnCRrtRR9tVNERsuaPT0MwmJF8Xz7+MPxE66R7w40
l/MDh1LNccxBVbeWbHpi35l4kuhJzl9CQ088ioNbnno01YBMskHnI8jDx2wxdNjR
EK0BImwec0U5Bw/WKmU+EL9Gku23IskyRgHSeCGA3fWLy8dfAckgVa1dANWMhO1r
WPpBeFpDcarpo+Dc9jOD1fyXa9ycP+Sf2Zz1JYI7pp6V14rb4RHJzKQQyWVZEk5R
tRuRff3wZF50ySE+KFtkdQ==
`protect END_PROTECTED
