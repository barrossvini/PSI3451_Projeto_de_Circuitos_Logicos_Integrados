`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AXWFmCbYxvz6jkPPdrHYGMaT/mjf0Ye7aB06adouwO+fYvoKUwegMOIp/4pQGiOr
m7s52XaV28S5ySORGYW7hEe2WHF0dl6CISW6sMKIohGNHPPDo8x+S/Xa10p4xuoG
g/PzBXaXNaafYzgkj6nEDk/niX+Xh0fZLeJCUcTaGwqmQOXorktbp4vn2EwZs129
7q4n0pr30WKdZV5MD5XDhsnB1D2gVw65dlLdPjsMH0kEAAkTkwVZUHbkiBP1cUfe
WgvsxklNB9D7fRL4bVJaWyJSVtWY5WbN3DgzDCYIT2g6JdyfX3l7iJRhFms0YcxP
RPKEUZf8jHpaqV6HTSDUZjlSAFUHwZryCsinxzYz7lzeqcYkI+decGaSiCkJfxDs
GnpSUH+cjfFmAa+SmwJ/saj7CxEnk6wJ6GDTsdFO8vWoyVzM0jfYwldXqlLzNz8l
lRjuCaJ4yFWuxh8drUNuvvrEpyldNjp9H+ZnzW/WgWDXs0UGM9wcvpdr2+c4s8OA
42Eif7VqVr9SSLrvGV9rpFCdPYS+jI5SJG53763nbXG3h2b3s0ICY0oR3iQN3TX1
+Z/6A5eAmCaBwhIr0DUTKFxQIS8Q8GuipDZq7A/G1JOpmaJcr7jMEO0Q+Ngy4TPa
EE94xwYL5XHsTNy2Qdf7B7I7DcKOrNZXTd+fL61ukLunKSrCNthKZMOpFLN9lAeb
CEoCYgSOinT70aZvpTaCQNpDjSRVZ1sZaCUPvE6Z1azr+qsx5/TlWE5YcAznM65t
JCpdPvI+3wn6HWt5RW7zLBWuIvmp5URUETxYdiltAroS0aWkj6U0F4RlqZi39kiT
DMoMNjE0BNOjjv/RffcBs1AhUq0QfyRqNpTgXtu5Pa8/FLCJoXaxQwjE+bDBhsl/
KHjqlFGgseHMKSum9pJkW1QzKUebw/DZLk4dLEk0ghA=
`protect END_PROTECTED
