`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dsk6W2GZ5mRFqUeGlON5v5vAMdYEexYLzakyS/WZg+plKCn7hnrB+dTbwf6uM3dO
4KAWbvz8wvFxBEGXa6Dp2u2rgIRYWRwWxmejgrWMBRqZsM9Bp5u0/ekc9VmXPH7g
j6Imt1oHQW0ttBb1+BY7PuAJcw06cjqKX1LpkFJ8VIhsIB4pzY9iau8juRc/bG88
FPf+lPYYYrLWni4HrqBOw8UNH7PKQh8oL4DF+Ff1x8WxWZgsD+KCKmToHnMpYwd0
1VHEiq2p1H3UNgsxLDEn/x0Sn0/Zmhx5J9riqy2W5W+vPlAbS+h3mfbw3sKBm2q2
4NEZ2SZ2zckBijTCTia0viwKD6ThbaxijUvwEwg1q69fgJYF5O9ioj8LVtyhLb2U
cFNCeGMyKMa9WJX4GNkykGVeJzFajHe4EjR0sM3fppJjzmA9suSXebK+TwfpwG3S
xwkMng7OM8wS6yqlnCW94RuMtdZR4It6F/NHNh4jyOyMTEb+X5/YE6T6AdnFziRa
HVKTlCIQU02dql/EBin+QzNX5eSVo/7C8GI6gLp+OHG6NUmCjbC1ko/BGWVVtC1N
pigxoWwbo14zfcRTfp5Ci9L4YiEfYRTa24q8jPdoisKlhWR2PRuTPGPHU4/WXp8B
Z3zVpjfyboFWwUs7qIBbl53T3YNB9JoW06B3XgxK7dBoBcUri2T/9WJSNaBu4rrT
ygd1N2aWRaOU3326eUDWoJX9bV+uUKWGrnnlGYQc2B6Ft37nHPnGC/42Mc8pVrlz
p2KvVE0UzVIIF55fbgICTOt0+5qNSeJbEBNtOKOUsaAdTlo1XblZQkLX+RjHOYSG
mtzxzVab0fZyguqvL8UFssxja5OlFcviwSRwvWIF70iy8ZkWNKmAb2cwDgC85Kx5
02PsHeJnr8Q9viFG2WLyKl0yJ5Ag/fJCkhhLoG2dEngEVNgIiHzdSV1QXXxp3jHW
1JfqUDFabsHq7bheUyOUpTWKBnY3FWhIYClWBGmirP0XET2Nnux1X296OHXPoiIz
0K+Cj3lnSTvCrHkLsvbR4wO5hzA+eAcuJS0FdnrrgRtJjI/biuGv/4243OBvTC3m
CCuVhm7DVMvzThkfAjCFdM/2V1QdFYLTDC76bdEL4TtKKPDq25JTVrPHHCbyljPP
/e1S2uMayf/aZO+zdamnwWycxC7GkzRVZh16GoGF5cp+h6tR/d17bYxYIf/dOViX
b1TbJCDU1AqV0bP822i5z1OrTlfide7FDl6n4wo7LcAuPwUz0YkoxqzY/0dw2RSS
ejQu15uWVL/wmnE+jLGwek3jxbSmVwk5htiJF41Zg50dJN3hkzyZAX+5WmnW3uFh
ON7St87DRD2MSreHqr7p1uGpJM0EtLzfGQAL4DQrdSCU6oWnaFVIn1ghVyQs+4AU
x1Zv91AOvdEHepE/FYlLiGwteo9UcxrypBA847F2pvQs0ju4IZKO8IzWHEzEXs68
8PYeqlsnS/KjnEieTo7fU0iEiIU16dAaMH5gZzKEUdCBol2nxSbAGf06EaBw8LLT
gSeqhTUKxnFhjM33mCBsxPlpjDT3zyNEVtlr2yIGlhZNCbKInxfVGv4WBOZ7sfqv
qiv1PMBtwgsrUAddZzArh82IQ0xcUF4BawwtfKajOhNhCw4TcSR+QT6b/yrCojkg
zS4lDLl4FsVwLST7c0b8YPMKgHx2EDohQMe3l417H+DaO7dC6e4LrNogdpWuTtu7
AXuQNF/VNMRqEXSQhqqiVdicHbvYnj7XEWja6xEJ410IlqwH7lt2yI7z2uI4KLUC
HXJxqE4SDxWbnZIiD61LgzRDTQWEu6HWknQ6Y5t6mbNpWsHHpkcW0O4vBY2HSyQH
drvBdo5Yn46g7JcTiVM2L1KtVjSGn2/VGA3EtZbKrwJs9zKmxXrtifIawykDnN9v
nOLy7uFDAtGjB/c2QKtm9sxp5v5pwktvlX2oUB0pAPlyC0vrnx4aaWoEHfMYbsFt
cdyb7ANvItTa2pjcwLJshEMARg+wpiMBLdZoUuIpjlYfXyaqJEOS2uiK2veDWfhu
yaNI225K4a0JpNXpgRi4Di8SuqAI7EkhfhPCmr/DpI2b0VzIFIWHlICkFNLMvejw
uiC6DFBpWYjLhdr2nl3oCwuJS981ZgrWDHko0Xg8CRn9o9tG0KCPvUEE5uoRwKLx
ii39W05BJEurg6Yvi0f9D1kBWylBt+tDxu8DkPPnlPspddq87Fk1L80ZVmBBJZO+
M7Md8IcVGH157Nqpx0uJuxzRcc8ZLh98VmZmAkIIw93jUzE+A8255NJ1YQOfwNnT
M9qazb9xgaLGaf1irWTDyEb/ZmoNh//6hqin1nRIxN/qA4h83jaGfmzN/vgMp3FW
fImttp22bujyS/OqnEC8CagjFkSWc9slZmYEO32rs7bNUGnZpyxX14rx0wKFS3eD
wnCPwFKhZq3PPL3TBQ9qtOR/pVV4GvhaTT4ucJ4KLeIyeNk0zMzGay6lWQtesw2L
F2QxiauB54dgn7myY9xc0au0sKm+sL/1Pg+iRLNmjp9ioawYTlTHBy2mz9JYPl0Z
AtqRG5DlNrVsAjTTegfzh2q1+K2KaAjbzR7ESfY/tGb+evoIKyRiqmPniQMYgwAf
LNRAHALgGX1K9CNu0WyZ25e2SEb4gAiowG/x6VZ6zrtZeSftjlDZCpNwQRX/SwV3
TDKOugi51GbriRmYug+isS2fLtzZx8NFcLer+i0R5DQj2/VQoi9vk3Vtgi809b22
f9x0MddX8PvyKbB6SIG2Rqhz120n7IWO2WfwPDBtl7t5lWCamqkjcO7LavbbbDjY
zCBFuN7EKPSxKYk3s4rSC7ryYk1YbUXPk/WCQMoAFqnGRcFQ639deps/yxffo6ZW
vnrxwcf6jNU3/aRavhsYmo396AXhzzpv+Zj0YSQDvEg+4v2tj7W13bgbpTEevj3H
C8Z+gKcJvMUNgTWJalVHkQjTLq0G6XnDDcAQFSGq/k3R/JRhLmf12BMqoFmyJMib
X8nQLrSrtRWk+O3sxwxI7l2/LR4a/0IRzZeQ2CvB+VHViL9891PrGVmtC8zwAYov
lGhiflPvbUnA+xMt9MvNqNfnXHVhLzdo8beexmHDMrod4CP4jyyrTPeLqlFt6gro
6l+eg6iN4WVSS8i/J2/uRqtDsggTqJeWWhmhQ0O/FQMFRNbKm9B77vFLplgm9G35
LuEmZ2S6jCARuCSMYoH7maSitRMT8P96JCtytCC9FXfGDzqEchAi0Ibcc3If+TXf
EB7kzZtcbr8gFY/1I16dApGRkirFZHwb9lyOXK3G0yuh7wUMEoxCHAUkIeoNUjwV
EnctkbaxgfvRqYbeJtbVPFBCptYoCe1eWAIJuY/M3hzo4o4h4nHTIiJ+rdlefFJm
KmNyk3axml2rKhlyuFUDZCaLMyHZL1/wewXFh+h3WD5FJMwoqt2uSqn9t6MMRVaz
wYGVud9j3pVymXo+Ilqi7CdVaRqBbhjWM3bKsy4Pbi2NRoz56C44rPRIKP4OScur
0cVgzBxdJuMr8Rsi27bTBWqMK2q5YT73/KR4EvDwb0MmY9uCbku1aUApdQeOsGg4
Cislpo7Sqds0dBl4YyJl1HdITw0h/tss8LKQtCs/QLk7aNUTQ7TqFsJq7Foj7c/Z
bYtTXbWhnxyj0DCBuZVuxpBq68j3vEVcA88TB2wPCBiDT5gywz6oMGT15+3/ExM7
gyD8RO04YdNIXDbFa+xoYWMicsS+4hWoT2BXb/3hum2dQZeq4voWqiZ4SkvmPoev
Padz+gowsflWLucif7oVb1ZrdcZrXRrhGiOuDEOS6hWk3XpEMuO/V98L4UKWqexs
bKqrdrniyPcv/VHZIbIVBuZ10bGYH+oLWmd322SQOijbFfDqaGdxt/fH8yMfHLhF
D/ETiUGjC5myiBGGfebx9dvKe/ZL1L+rN6Q7TdyAqJ2yVCC6Uce7uW355KcWBa+j
1qKaIRpOsbV6g2k4K/lOmBaY1/ug7+gu/AIqXdCkfUpsIdSdP2V49grBCfx98vjn
YGSKbN6wNEsJO15oka9axHPXpdJMFSDD7KwhxufoMZozNZos82cmEZr4VcS46S7p
+OUbCzKZ27+aOBaIWIluBUQELnC34ve8wcLBauhtgQRMFv0PH09IU9cZcnFOFBFh
fVSUS360gGtdQjMStRPocFBLBxTmhSWf2MyhcbDVE11hXD3ygTHLyBLBScy/IGja
gPdVX5aNrK9QeO94ArMlNREF7JrASlAZuiY4ex3JOFA/c9DtfdzMtoAH/+NAbzE5
ZcS1ezMue2+IZ61N88nYArVJWxVtnLEWu+i/Yg3BRtbzMXJq9HveDqYE12Kzadq0
c0gTG1ZctDBBe7UiMbT4EImf9IVq+GjJvBYqKd8mKK7El5BKXMHev3rp9/CkV1/z
8Nj81sYqmLyQ/hV4ttNTBk/2yiOeZ5d0v5FZeUJMEg8fktN/Ba2mMuVzuBt9pPv0
muBbOilXNKa0HFWEp9oRfXJpcB61dUj4ri3gCyrWQfgf3Al5gvA16OZaEfYxTrAs
fK6VhlSVpGZPB1gxXD7jNgMW1eWqi2qReUWJH3ItDw6ZOJA/MZyfMyPBNAOVzpHm
3KfSI7IgRyt6HIKdTTuBXcAXQkKrEW6uukdumaANQhYM2kyRsp9qcxx4raMqdsDQ
MQC01B5JHqaHpVolRI0MIcDUgliaiAbyAQhwxx7A5HO7FQTTitjvBxUHMvzd/O+G
S8pdDC/d3jH29UhvUrxzW7S5Hh9ymr9VmQKDO+WdHbwPzyDZZiPbs/RlPTX6D/L6
+3qm5qQDND1BCjX92YOTIODv+6F2TfnPTpi6Ww+Ab9Co0VgyE3VdlxDJjKgF+9gx
ni8r/EoG0XORKoQsMX7JRGfaUsi/xkGpaVzs94KgdebU7VbKotS3Rhz3MB82B0sx
w2kr0Q9E1IseMEChFr4ScfvkbIKNqhF7XLLboM22XPAgFIq6N3zoL2iZC/l8U8tZ
OCjksiGpFzpu8gTje9grcbug2katqJiBmSv8E3SLxOCCzx/pz8gAJx1Dz1CVF2pD
5VlJNZVJcly0gG0xCOmeCCKeJrgbRM9PuM9KGcabcUdC0VpCTqjokAC0y1tR0L2S
go2BOvMilAVGf8TXEWlxgQU31IsIpmMz7IXnJQZosCFtmfCiNSMbJVbKPGijfP5j
ETFncY/uzao6PVOk+q3wrX40nJUHGv79sNJH3XWVJ58u7vBcS5X45ZUUJFYc1S/L
ceY9ITdO41N1ZjKpJhfQNJ8it1u5KJOwTBZDjhIo50vYRHXqiBZrLlO2dV5L+FDx
RqCPdjF5agTdE0r4RQYWWpzDBA4/rBcrjRGmMWKwFi1opTJlyZEwLyiWfOlPbgE3
F5yNvkmSMuXjzlD2KQb3socon2skGmhGqck406S/3y4yqHr32zHXE1ENP/SLAQ3d
xHszBjOvhSFRX+iCzcJYhT87s/6lw46n86PzZtxSiaKq8zGQmv9G7peQ9j4npx6+
yCX9oDdLrMB+8P14tueNnZpzE+OMgyVXmHaf7KuiON2DRNUlirfn7+2aPW5XL6Hs
yP3310YrlmnnQorx4RTXCLi1uTGUuW2ZHCE7QvNbI94U/EegpyGH8QaAoukLxT6X
SclmidvIY9FwAolF6QpiCxgVoGGpE8DMr6eGhDFuPi0GLwwDYR0A5m2s5FJjiM6r
qQP0XJ8GRFthmUKZQXSRDendtuNUfTvgQ2pqMLurr/GhpI0wXnuPLpVmw3Kpa/ID
4C+q6tLOFl4mrQG8hSl7A8weiAsxuyFqYZ3YPkmXu2qDdxb7/FNmUSFKMnT0JuKO
mDA4/iq5NyKD6BhGxIZ2HNNvxy/9zqA7H0aoKBcJzSMKkLmr4qfk2Lhw71MdghwC
gKpcGce9aJ66V5g/rD/ZngTkeQAgkbHlmmiSgVH3t0wePWLHmU1HiZ1qC8HXpeO5
QNLRZRZLUP8kXf7jARN1G8ekVkLnYRZjEbes1cme9bPdxwfyttPY4qQ3pPSc4elx
MxTNoyKA7KLgk51DbE7oP3AdxtnnKGOHblACg7UQOQF90BjTbOQkIqbsXGxhjYoU
/hyxuZ6s0XmQBhazGPUxO9cafoOvTLUT+efFLSWocjKi8aLqbUbdW3WFU0fx41S5
sT+xNTdTyt1IYl+wt1Vcch+q/agetc7uwiuvZ38VXpVONNR9mZbh1XZ/SoehDlcY
khDyB1PhSh35RNqZFDbbEOND7MlWi9JTq57trO0u2TuriKN1Jq6nkK7PHPaZtUMM
ENHVNRKgyeTHRCLhN3WMwQ9xP8JMb+kBcbse9wmTrh2Q3d0Rwzp2OeCE8q5fHu0E
oLoTnSD062/9K+5f0e3PWt9tISfWvz2EeMU/yJItxBHafaJL5ZW4XUugDeHLT//b
XoOm4SUTXhU020p9eXZKFLgZofnZCZx/PEsunns4XKiNnswP2fM+71jGnFvINltr
Yi1zXXHAHvx9zsdR1t/CvCJ2oFcuIi2RCyRKOBSYGnZXC+AXqJ4TPb5Q+QKYGywR
Ats1iCe5X7FbYEdMmhvLh2nNYG1X7xKdF47ig68d2NyVCl4gMcX7Wn+FfQQaXBfi
Sd6E4rIJbqykh8MGqwnSIQxk2l3byeC2OFCYlW/SvecJkRlLYF2GY4d9bU2kPG5j
xmimxOwqowKXmaVI0gYt7aNUixmLGnPUhAaa8Ixnl1DHimhvOqw/G7NW+/Do/cZP
iiKDaZ3a1IWOEuhw6G4bYKf1BkAbQLrKtg38Za/T0xPuTcFuvWexXIgrh6XSLHnU
+iVV+gthd0moCq6tthqEvzN3VsRlCM+86hwItTz/IFmtLth/Rnpb3AwtN3ZFCVtQ
cpLtg7yc7rTXtuOGsQot/Zqx+kXKQvCpOokFjCwWOqzml56vE2SDuWXeXX2WCfcv
59WlGZiZ8/Xms78wKfjzddS0bOrBjimYLkuVYcdS4p9OyCAL8VDOpe64jHX8KLAR
p71G+v1rTPd/HeBh7pkebQnfWnPiJZP6ZAoE4k/B5AygASUJ0iNSMCOQK9wreZUf
5eDWfXz6VwWt2Ahg/Itd+IiqCJ5HQtKQ3Cej//k7MLKDKi6bIOHkZ9nTJ3IS1RTE
/YovD9WsTIU9g4+HkyQwEz/1W8guvZUEZw92Ys/Hsvzsr7RJRt7JWNidLVplDzvU
3S4Iq4jTWjKcua9CINjIiIIMob1g4xmmoDiLd/TdsmoEaiSwqe0kQfLH/4u98IP0
6g7vh+Xrqy+SEr4fU3ZnfN2N1u9zE391z8nnw4ze956asWapPn9whyw2YJD7aMeQ
D3xtbLh6k/npv5kbrZNk+cvDEjjrN+FoDjuK4zyp9iBlHasHQBqXELi3scmOdgbR
OF524nF1lmchzfqZv8eU9tUCSX6UjepV84sJ1XRPXVAoAu9nnqxXKWpS6OIHKNIc
9HqXhKPhp66rMERYZu+vXhBBXVNCZyY+Zy9fBZxmMP92ybg6clvm5fJBjDDqASHO
A4WbR5F4Qxo6QZQcXVwYMDahNFcIjxfVK7OPPDkWGF4zRLZWQfAB27Wso3dVetL3
fufW+PCB95TSULcKXdjWqY/4tEtjBQpQ/68Fawuokpw7e98C1fn+DUAeazuageTg
NbZGoj3iv2YXs2Ea7uiHABPUUH4iCfotS3awQh9/G61vqu/dbXnCLSSBnXYgk8+O
iFDDj79lDFAD+Q93cb+FvkeZb+LDDQX/4u7zveoOhem9rk9MzDmR5cT9eETfZUuu
v5akHYbc0M1RvlxQsWQvDeOMeqXXOL+sq6eiRlnfCE3OaQi0e0KHxUEsfApgz9Hq
WbKKTHaI480ciUix5/AtyJkmiwQxTMPK9yV6J61Y2leXZYASep/XyChlB6lBCOLs
ox9E2X3NwFjU2OIlMTfO5JrfCnhQLo9s1cBo2aUlEyTVjCOt6htYWYJsbtpT58Xr
XusXMncsKWfPCdLAU5j2Dy/UWlhadnNThR4hiHWjWLnQWZoqmZNAe1X75fVvzNHn
sD7LDSgyPd4FH7P2ZFnWnL1oJNu5fxdQZ2gDyM5FvXIF8b7z8FYX7hum03U4A02j
J9HxMm1wWq+BUMPWcYGnT+i6XypRcBgn7T0pWAP36rzrWXbu3Uyo4Vx5Ro2JavMG
dSAaF9LNGyzJOedKvi9vtPDtMuTBVZlrIssDVi+AiQiVkWtho/C4FhD9UN6FLWEX
FWotHcimUu4B+90DOnEya4jL63DaeV1w3fPxGcgi6lSjSbHbrqu2Fn98Dv7FCe2u
iy93fyt3qdp/CfJr4diafZwk7wkVv1+WtbGqaJK80fHhiNB+ph/GP9hYYskmibhz
vLJsLrQ68dRbImzEIeNRVNRbaTUHQHctg6R3FyAgd06qQ5/7Rk23dCEzH4T8hgXj
lBJCMqwe4TJKqLPwwfYYc9IzuEtquGNn7YrhY0cMOu6iqwaPYe28r8GuixduV68B
go4YvUt6kw1ov2tvHit0vfXasJJAJyqHEjikx6GmwesCF7o0QotbhhyhjVsauoed
AnHyZj4cPmpjRrPKg7iEoUPw15D8jeKYyvFT7t5pmZd4Dih0CYqPPmKs+MlmM1ay
QRA91Uuv+LOh1qEVxdnDaGRq0/AkOI9UVi7kbyzA/G5WrVuedpLQgaAJnW3sWLed
atiQ+6xbW11jB4M18RgklUQAGmqfD6YPrwBU6RKh8uXJ1OeCQiaCtkLOPXNFzFes
xA+kbgNOob5ox3JgvHT77ljHSVtR9LAeJvM48S4Xm19gfOPh6GztuQZFnaGP3rgo
Ps6IU8CMW89m8Gtqxg++Eb2UYQmvlSu+KQqJeKJg01aCVKqKEMTJCGV7m2rOHjON
xe04r34uswuanMWATLaNDzuCplLgOKyQASRIvTxcRYDdISKFZTNYXMcLx98UoVOi
XnynyzMOqDgRD3oEjMv7xT7dMDAR02Imz/RUxukh7U7FmumoDmibIykftUHXVvxC
FfKzOD1C29kRCSOrE/fNCh+OVFTMsQHigSeNbJSEQ/apQvVMn5e9wbs+OqOSEpki
TY/9LXRPzm6dO/PHKpDiEiwhRm0or7a9JDtItGru7+6VhJy4wJU3HUZC0RT7wC4z
YhoXmqUruvcg8WHKBcX9pDGX3jaqL9S6eK6C5G1LR92GxqfF4VoBrlfooYSGK+2m
AsFbEnZKH/4bM4QrzclvYCo5/iyHEE+9uWCFT1JbXMv2aNVHLPWJvyKQ2eHcjLMy
sjzTTUsRmcLefrp2U4RARBFiEFSfAKfNLkUM7K6Dy14pEc114k7pyGRJk0OPCDWZ
bPk2hp9XuqVLRZHhzF17PA30U6115zH5Sce6pnxWHu62oG5vwV4MqhBh5cP4GcQW
ftbd0ZpymfA+CX4ENwPP6cyf0fEbkDwNa2dmQpKJK8jfrJYVfDZmXcZYO1lehRZC
3qzw1o3bFH460Vn8cBxbhBMPLdBce8rO2nqi7yLNxkJeABaLOWdoljvDc3TEUYF6
AdMWG9OQOMngv5c+d7N3bADLFpmVAsdyDtjFpJJ+EZ+5Ffr36ey4Wx7HEUon6ldu
HxdrJoiVef52POMO2JIwFyC8UzXPsPvc9KtEbpDfvHrXIAzIwozLGSeT5INqMJ5r
9kOy7x8gdtyi3grxQPoUPEWSCXJ3bPGUcKsmj6jNYqpMqfAVfqINdzjhpwzOfw/C
JSECCSW+9ABqBMBHByuTDjzJFOSAiTNQo0L2IkrCOyPBjhAZ5rDcHeuagqqJCCBZ
9doCV2uJ7ULvLC/C0R4/+M45IG9eRJR0krnwRrIhVcrITazDKMgqGIFdhaXOQTaS
/8S6Aw2utpTUWqbKJ2f+G3EFFDP7vjwjD8j0DbhXh9rEwdsg21w3ZQ50DInbzKmy
GXshmnObzDQNPINx3mHAICYFL/W8BdnU1X7eRkYzg027dUTkCwBj/mzJdlZenCJB
LXPkezc6j1NIOf5Uy7tqkaMY6YSCkShjtPH6uJU7Zo0x/k+/iDstBNq65DJhig5g
NJvA+BoYG1kkOGph0KBlBeGlD7eM913aTl1wkFNYNNRNklp01vuMKueeAOvL08aZ
OX0tgWM8vrlZgmTcFQ3XZNAuFOr1omx48j2U7hsSLcSUD2Gz6SxyCVx8vW/SIsKN
qweBmU/a8qFPdzTdS7db3BOR4mJKwPEaKm2iop8NwQA0I7MPupnMj3HqNlRttTl9
422RZs/scQBMy7SVq2Qy7UNRzqLWmZTHqRIqGIv9yvGH330Z6qGrTXTkkchqIfJL
2UvV5VK/gpuIERh3YlbB6fEsK8TlpZHiq/pPOCCaH/oiG49iAKp9+xAh2DBLACrJ
Sut0B8N+ddkWKmv7/imjdgqYIs6r/ho5foHM4un14VzaGwWw/YNbJfb4XylMbqTd
ixvVZ0ymuuSuIKgX1RDLoFPrnRPkqlvdeFj1sOCppDB6v+YldMjmRouWPiQncbBn
5HGS8s2OoacfY+Xv7H52+2b/3zaTBF9Dk2mgugdOVvAkJYXLHC+ffjxthErrqnwa
woJimxQHdvktqQ65b//0aL7ys666k+qOHJqONaqBagCHoA6S+tpSg6Kfd++3rZYy
WR9BNZkKp/JrsHL9+utF02p/GgqdSdxTwfySFmbJlZMw6Mi0EgAFnRh3poOK4Q3Y
jcv/pmNwZfqHr/MjSpUNbIB89It6PZ1WTkHuwT9s2K3G8noe6s/gxxOxHO+G63la
cvzhbAV8jZY5dHe43hI9knU5jc2rnXkN0Plwqq/63fMSRg5YZ9Kh1/UfuHsOVrbJ
qxiLLA1f9GfaCW4ME7umAyDPjLrIveNXwMl+d4oeAJFtgEVXIWM9LrpwAwMZK8Us
QlR1zKJXe3FbWPHNi8yUm1TYhqjJeyEd/jy0bBMzmqPszAta3Xw+HhIgO2yN+Klz
Te8irijIIn0NXheBk0GECLfoLfXN4jWBVJiijRiVYRU7BBnePy56PHVrzHnf0MQr
h5Yvy1ENJ5EGemyfj+NW0yg/bebh2c2BISk7//LdgCSzhTG01aiwr5L/6sxveTmr
23N2DACAqoRGY3cd9rzxGsiVouSoLnLovBg09fLYa0THGccqQ+TexILGEE1ETV2g
6iZk3uW8m490Q/U6RVpdmyiwNDb6ZHVWcAaDbIT77oluzjHYEtsFVTFwDp4t+mit
pIYntKvnkI4mClljB8eGMPbbzB2cfMGO/hWKElCyQsaZ3b682VZo8YqEE2ynk8Ul
FwZy6uPF8fIh3wySwVp59X7dK39Qn31fAZEI3USO14EKcko5znaQIIObitQNtjpH
Zk0/MTCPY4GH+XZXG+VNvZihd3/s+gD/IMJdGeE7toG/1fRwbg2qH9Po6HuIuqeB
4EYU5nbGZ41ARe+DUcffLP090M6iVY4guEonX+yR5T/5Q+sSx44ySRGtCkBVlmR0
znD5Aq8ruhMIEuc92PQLkmgqfQ4FAnu/Unm9u0UHtij+B1qwqp+JSvsF4IlFXGqm
12g88vIVD38IBcfdN809lLPnaLN9Hz+rt/NSdMDX1H008cDJ3ewFOmQljQbbWPvv
AuzYCw85yJ8pBsYQXRT9BwM3L0EyiCTnxexHIafe9G8CSn1x7IDpwDPzNbp9XhGV
R8zroCmM5CRfhXWshOnDM2iRAttFX6Nmc5c9q1nbxeW4fCW+k5qW7t+QX1Nm2E5+
kKroF6A2luwtEgCECrZHn2G/uJV3x7MZJxgHGqUqixCahujofPWo/ucVsgYAyN3r
kkSy7VPNUU0WE9YzOYt4eXYREdO+BwSFWuNRY7/rCySY0pYg5s5FhCqLKB8Tw9TO
humcShHtAxizj7AVBs/UrXaN0+c6N6kPhG3JQ3I8VMlI7N8HX+Q/4GXMC9wTCY13
i6UmCQy2hNO8Zy43vZFTxaI+mfcc9iLhl9rN9Aty1dh4tcJbVlF3tbxQjkNMcxj6
Enb88jF/2xDwhCi25kFhVxd1CEl7alfPGXVMN6haYejFhins6tr1KAMiGx1NlHtl
oL+nKAGzMGqZPgStvPlDQ5BMXkYlGj8579nFzPeJXU1qO8alm2/owp7yR8RwSHDn
QgYvoWISWfYLfyOPgQD1DdOgpOSyXLD61Xe7/kgL7NzFLUaqG4YnPGI2eIgkpkd9
nvOigWUjih80T6Fnk7rXAPOQhkvU57DDgIPCycDImt2KAkT22PPqfJItTMeL48pD
Sbn8XcLz89+/fkEs/o4tQvubIlYHAB1I6OsAWAoghwUSFJL076R3k+16REgczxse
3qsnh7VUAg/iiaYFgHxypvFtwaVxMI0+GvBB++N6Xat3OlQdo9V4M8VT6gZHUsBx
ufu9N6bpCp5ZwjPB5PO7vGqFjPnL3mC46fPkaINmf3h4gUVv6w88G/j0ufeSVjcT
g5hRY9cVz1kAw5yE19TQT6dD/y31X/IbGRh404S5dqtPpz3G37iwVT2joLUqXwo9
cazkxfIabCqTznYHx/04jCvQXqk9SrFLZQD9EtnzpCC3sTKsOfm+ANZDXZrQ3Vhb
IeKq++FLGkWuM2ESkdYTB8kCPwRNz957gGhzyN4tIaMEFIekwJb5zNCNR1UOVUKY
RqsUYv8JPtmsZ9r8fvioZFUMnU8Fw+dMJcXPo1fjq45yGysQ8dJFl1n0efSi2iE0
XjTy5QP38Q20NJbUcR4OKhcALOscKAcgbGQ4t+Any4j6PEYs2QghzR5iu5Y8m21o
hunt1+QgEXsVMMzFw4uGgvu7Ia/ND10uaq1lNfEjKmx2CeK0SGslHgGhwysuSo8n
2Y+Ton4Juv6GLvjHdQ/oVp18T/FAp5yFxtZuE3M5Vi6Eg72rzGJ8b3XvzQIZc9VL
CWXx/tfPdqkrAe1vSQIfSd4YRUdNmAFPXmBexeuPDR4JX+GXKXgETdhk82sODWoJ
WnzViccB0G8ldqA9qyrBWIWj2qWZ/t3NmIMRGCqxxl4Tk/khSpm2hhxVraVTUACp
IXRq43iLwlJbZ8tn4hpl2GtZeymfjwcoIhRWO+leOs7ATpRt1WBtu/to5JofPbfz
elbIY67DJ/jmq2Yjn7WiQBahLLRO3Xt4TDkPpM+f4GhWccpAxz67zhM/q4XRRVWZ
j/bC3xsAnOSU5qToxcWI0l8crRE6Xeg91mLfPPUUlD2yeo7OWmvj0oWc15t4motb
qb7ZvyLZRawqfEUmoT6kdcVPgadPGcq/nXaiby2n8WeohiJJ0AMwB/+9Q2eonkaf
NnPlTnScgUKz9pVUFgg4SGXhVPjrkP+OtpPFVsI6WxfmgKWpPPqbBbeMn8EQjG2V
TlGF/zOQhKdoixyIKn9cqkGIPpkPEnhtnbiwWf8fjnM3bbh4PrMi25ryW5hlQpw0
B8tujBtkXQL//4foXkdxNXBNZK0aap69tdfWBgdZJ3Iv/ERaa786vNuAopD9/WQC
7/7wv8tyoAyoXYgrjtx+r+piaCFMvT9bXXsaE4iYtKCsuH/fotYsVvFsJUoMH7kg
kpyqP3NFj/ipUVi89a8kj6D0LHvI0BB1H3W7akH2PjRx8mMpyDRCMozFF4l9TY4i
TcQgBecMYWrcSNOLsqAGWO0SjUXDBmN/S8Ay8fU8fKQPpjArQwuzelKDxXm/t/v6
Nya8srx8OnWHeSWGniSij+KbahGeYPcjBU9jpXq6+3RUwq/JTaieJgOn9rm+NzQG
svBzWwWQ/qnQwd0dXlqBd5tntED0tPb7dHECujG74EKZaAKMylYuxKImIbNZR87Y
z5psVZphIjfBRqo5oYwJEzCeNhoRemDez0Zq1ExniyvxiLLchXO2TRTEL5qWxuBm
99QpS/iS9QLn5So1mLx3TKVOkNyZKv1lIQ1+xisiEvNX4IvYItC+6l67vAujHlgf
3xnR0+wKTSgGeCFo3mjktVptfCWl+ATpW4uuorG9dXoEsQUD7gYSr3ag92wKw1Cg
XxGdmwlpX+OYHkMgi/awUAnm0v6hlDwjjZe3qs6D3r7EKFz9wzyufvK5EZhNVvao
wFT/4tVnxkBUDPp1Hf+AQFRvy02NCsJn5tKxnUlEMP2oKdql7myeqtzpBsqNvjZm
WlcHQ7T82LOr8ESvXotwtMzhWyUjdw+yjP7FEBpAboYB1EekJL/+h+Vf8im2ZgSV
vRrMbJ0EgIVpmoQV9E52S0YzXvsM9h3D6h/G1fygbZjki7q9S0lT7fBT60ho6YRA
02zQTmA6bmCY39V5d7rhplqLqdmhgbv1Dc3TyCXbQfZBUlMd94qXikE2IMemjN1L
B+TjhymdGnM7kggnil/EgDBMkoIYH9RIKFbCJN3qhyl8z7gYKNwT8Om96ABcPKqK
1uFdXzLYiZM2u2dB05FjYA6JE5/aXKxt+7lSgAsC+rXtR5usyPuXpONrUQOhVHNN
ndjoGRsciKoua5opJ8tHNXgSKAwlyZZNRpMAwaZvsu/+n6mfG6MCZ0M6rqRe88Lf
tCGJafbpMA8Xa4t8xps/QLwsvJ3nJizuht4f/6FS6Qvbnycm39FvsfVBGvnVL/2I
5jDjby6lvxXBjnRTd79zZGrrFr3jdlLFbqn1m8eX3paFzEYpyPRACjeoGVAfZa/A
gtTCF/0kpxJvURJOjFZ5U6/HCV+MoSbWvvHulr47Zjh+UNKehRxPq/t5F0VR/5Bv
oeq7T9Yp1W+QTrNqmQm4n5AXO3h/A6p3qM25WEY0IzGoiwHAYdyo/XQ38rs2GCQT
Q5Z7J2CTljv5Jl+o7nLWBJwTlLE8dxo8VRDY/nSrGUJk0AHbeuLqqjdyNPrxaZc1
phuFkw7efmzXAHHgoMRWylOEuuvZaGEjaweDO4d6r13jjjbsAcV1hwXIRpDowuc5
ssMM3pltc9+WQXrwmn6QHbM7E9mO7YxDnze9KPnE5lFldOal27FQeaMzvOivoBzF
j1WtzeHr8G0YMs1L7hS7PFknkAkN9/lXi1fTnqkvi5Qbiglns/dKyOqgoq89Bxk7
V5axMGJE7miZrJO4INHW41m/16WIgSBuNIUwqMtn3FG9kx++NdjnMLqR2+WJ+bpI
2fN7d7SzdF+ax6iLcTUlvhGNNBXVQ7uZ8gljdtgJgGHalR+W8i8xKG14mmUr9QGe
Gbltp8hbWaxr9pRtAHVjdzj7tqJXNqZRcKRhbQ1djAA6cRUfWSz304xp43a6cnH1
UYZ4Eb+I06sZRFQJTKJbV74WEBTYaFJny1bz9D0JtC4dsqjzkLG4VCfoSoFpotrK
KERSsREOYDQ73q5czdxEZjffR3xx9p77kdxF8oRg0L0ZO0gkQaT8LYjy+0L5t0dz
oihYMYR3R8VAXgV0ppAsOQ7Z2NBypRmiFJKs2WY/xUJDE647RosU0AaOPxUJcvoX
mFiQ+/8n4izgrwNg8ALSEK6YId03sXUhKpAl/F2asijpub+Rl+MOqs1fDapUNF7d
2/XwjO62C4iTjJtvajQZztEplTcfFl9yzxXnODsTCnHoiTL5mmC03CJjf39p/fRY
am9zvl4oZTQAYiIWwt6LpZ48JcCPtqKD/rk/E3k8jFmp9Bez06y09NR73/Uwfq1C
ghkWXillyiWCWyjRzc0BcvDuFNbFZXSdPgb3uprgHe8=
`protect END_PROTECTED
