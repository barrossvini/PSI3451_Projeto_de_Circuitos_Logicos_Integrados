`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LPMyD84S6wP7NOE653cZhlj5t4NizTOIBR2oGR25Supw8xMQW0s5WuEbLQijWg8/
5bm9laBqpd4vEQG3ECwLuWE/X28szN14oTwuXwWZk6lhe1oH6OLApViVF4EmMcX1
C0uSq2dGXiwCT2gWpG+Ipi7ZJxHUqFs0LcjzYC4o53/ToRs7sZCX3KtpSYdJOBAf
l67if0gEj0t7uajG+A7WXeIKkvGhOMs5BKku8b80TG//hYX8n+PGV9PRlK9o6wmp
f+4Ev8sTh5TyYmYM9CjgEu4/fhvfsPLATnZ78XtNf0Ta2eMCC6UpVe/Q8FK1Sxar
IY5HqfmB3EkWO3QwBDe764sQrDt3GyGLs0kzBtx3Sn3fJm01nUWGdU1mSDXdT1Hf
MQ0lj6sR6rGzU+eDnknYcHdzOtGCKRbaDD/QhJaFpbblA/Ix4cKOcjzaiOnBencG
VejRceDpXSz/50TMGK+n6fm5JxRA/kl+9p5tRr7bxGtn25xDrU4pB98+5D5kUeZh
e2TfEvBdJfHMliMEZuRvuieCCttYYXaZ4McSI7iKqCxYyrdns4zPrX5tlYPH46u1
971r3UUhsg+Hzj2+Mbjuhk51rkYNjWyNVwN2Z/9jXnEPtOls9oDBWxZK7u+qe1M9
QNAAHKQr1/jUGHOQAh+SDdKQi74JMAu5NPA7DPfSphTrDjD4m75XVIXCZzFc7PC8
DpQBFzQCl91EShV3dwktQVEk6yBtft/gPYsLyQuIhUKtkAsWEfuNpjhnkHJGw+ru
FZW5xeROMk/G7wpw0BQCeTJ8off72osMRBObyMzvZ1u02rkDipp2LcGvA0PbjEcH
fLtQK6Jml8QPKbulMTwI/zQYwX9hZ4mWptz/dXrSL+4OU7/tHsCyPsdwGkTewc0I
pJIxgmJvNNfaNOYXUaKzJ7BnCL7VyJ9CWPf3o1lhQX+jE4/aC5qzpcb6L8g9Zg+/
7eQmS5txx8QbNQF7ebCrLSDJ9uj72eqCIvwk26TtHDC4gKuBCatFjTpTwyiMmlIF
dgu8+jPu4Q2OoD5bXCW99/3+x2sHUcvvVCAtMk2WTc3iBDdBEyzJNJqdVe8juUWB
cEUKAwptrQxnInR9n2utUs1WdrghaEOlzjJ0wkeAugxcLrx41g3I4AoSpYTTerpl
Sxetjy0Tnw07soS/1aDXgrTAreuFHg/O7hGJtsg44oNk/ttsELRRV2uROF4ysh4M
Ziy2ay53cDk6HVyfRP182ZwCqqfHPtkpL+QIyezQ+nvIJq7qVe7ahIqoHggnLZ4i
ze/MwydsftUcLeNp+QcH77MNfkuj42Xu74cNLakpmJArjvY5WXfowONH+TT6NYVu
Kf9znCOs2su0i1dHWRvEkmJjHWhE+BQN6OBo2tMOwdOX3Jz9nWLcigc9L3vICeOk
cXJzCiLlmLYh9Uj++qh88kEo2Fdu88YelO2hfeaHwB9KbcTmp1qL8gMCiRnaRc+t
xvIo9qyK+ry5gZfx1MinFBvMZJdP2DkXuM/R+jZjIe14DYKOaIvV8IqY+sNeM1Px
n9tHYXLddB2xAYEQtxKpGnCnvthitEHeLgI39ptWDPonFH9v9g8Iyt8h8R9ZdRc6
PnDSe7c6KT2IrnnOm0sBR2fy1gBkd9m9+CZA8FPEAMEPeOLwCae8tzHa4SuVCZIc
Aq54+lysqhVzqtjSpFYDOSUMCqtZJnGwyw3nkATZVx5L96RInHYgnzQ7St6MRa6V
gUOvurbfMyEe4hIR58UPkaKvzVoUe7HSIgTkgJsQFqARO4X3iynNdPuFygqG89pC
xERP6lmQHwL/TzmOjWATn7skFubpvFkoFlNjhnM6yLnCIf6mXrDm9McGxiYyr48U
JZcerlO5IRsLNesNpnbwz7Z+5KnFZhzyDFG7xE6mMxNd2MW34TS5VWA7sYAjL3En
j8FvyRUSSI7CbOJEJlJJvc3T4qy8LLUsfcJ9CfGX7cuCEPrTkwg3yAiuP4/eEiYq
figD1XhyC4M+naAzw/V07MQ+1XUlvF1h40uf5pu4Dz9Hwyk5fuxRrBGyKuBweEtw
3fsE7EXBSUmZWpzixJawXHc5bJ5JlPJIUzxBCLBa7Jfk0vp9Yscj6qo+T545FFAN
TPe5RHWd3wnNarKaysIM36/b6Jjrwt9pawK7eNET6qkv0XbgVWV+8+cQv/XMwvE3
0ubCy+rj6pLlHbz2ZODrAayYvPjx0vkZFX6JuQj9lgTsGkWMoc3KGrICUjDzY7Ki
+C/eC5Zequyi0DiapADlOlNVPw4PyyaiKmUP35cIIn1CKbfthd/T19SRcs294nLo
QoKNN1MuQYOwRthKm/EKh8JJFcwc5fZhj23TsN1G3IfVfTE46drrvEjyu2XheQhC
YUvP0OtceLc8WnEMumVE/mZqVgE0Wl+HJtZi4EpCmrvnLXN57mHUbjyK0sL8Zjaj
LfAr8Rxy+MM3Nqx/H/ApelSNZQZk3HkbUMithlzTQPNVnOurW5+hba+ApTa0OrYx
oHXne9Y5jShUMefCoCnPKZNF9KbxQ8iRdStTf+284OvRFdQrIzEV9Fo97NaL6mRc
kMTaflFPGUJt/z0JM7MO1OhkCHLPu5gT200YKJXIi/Cn4AV5MBUktkTQ6URTrc/3
qcolmbuL/0dJlJxSBLy03vgiPleAB8jyvkwYrNl5lM+1oIyVg8eVdKD5XqI1xnX8
LiKjeyad3jzwyDMuqvChEGf+Cp9qvYK9xE5ZUqGQbU32FcNULJTbgFeKDaDiRMvz
kbWw5NrP95PgALLElEmpjyRDsXJ7s9DqyGuIh5vyD8e/2QnuVYWrMsQEzhwg2Cn/
CfFeQHZ57PbR1MoIjhNa0V0owiWITl8SoSj//b40Aa8lFJ+IQkTghiNG8bUcLoNW
wi3ai05x1WT8qbxN21DHTB5692CiF5fuURKoinWI96oeFilHU7yhBSMp/0/ljauu
j/d8mBQEZ1VRnaicbJWAEdN4TH8TqJhjTScFcKk92lwHof1GFXlmDQUUPcFtENZ7
x3UGJZAkgybqv0ZxxMPad0yN5rcfTItlQC8UxakXArnmp44RUMHxLflSL0N5llDg
nqPMrBQ6nLdr9s7dVLUPEvLVLg6JyC9aTWcSRvLcAxlLN2Hx5woUXNKjBrqkrGJ7
jh+z8/xMDzf/2JPBvyhkXytY6Kl40Ax6J5F7eW4EsyWsEy4rFKeUUBvgbTAuYXjI
GwQY88+S+7AL0vCxHUOMxNCaNKlno7xlY/wkZe/maW/cs+iEYDD2MMKk0fG3UTC0
RVAjJlftEtQ6MEug/+SqT+remxIyQxatg7Ey9KVS85U6bZm4b74zjiNsklrII5vW
cTD3xq/qajHAgUjutfrQOtBX5MOmYB9zzxAey3yJV5BPHdUVaKTfRnzXE+g1eX7Y
GpR7q1J9WmRNrFBvoRx2hbXNdtD5qaqpUkqN07XWa03ocr6qlaO/lu+IlymJyVSr
O0jSq2fb8a8pwU84dAXmQIhF121xiU7uAD7d6nrHyDpMjaOKFAZ3T+3FBufXuUll
wOILaKnxS549QHFqBOXFV86Tl0r/jkd2hEscNUjhuw8Xe9GD908S4uRde0ReraVI
18pvIhpKRCvsV4Rt0TpR12+or6DM/YERRoEH8LwUFbCW7PtvonU6hVkLB2oHobjJ
iBbDOOdFNJNo1l3dbhn6kJ7GKs0cS+MvYCyzChBy0JdzRrh9NWJJOrM+UJRhiYOT
8I0FNieIzXf+AazYaRykCrHDdIgkDJKBjIs0QqvkE63Ovn22Mw2Q8cQTmWOdF+Rw
390Djj6UIJ9Bwsy3E0u5NnnCkio3xbxXyLUEXJk4BdatMUh1k7DXG9YlQrSdmh6K
fYvtNCpZvkKQTyHfV/9dm6OYtRmAJeE9JivZPaiV0l42nkCmVTXDjgfmqA83vlxV
Jd28hjNtS7kK9u1tgyJ+uoTvkQPc0slBelYDoZ+mqQgudQx/szs6xBTgOrBHF59m
5ZWCR2x7l5lV82zBLkpDI8UD8mYl/op6CQFXPg+tvr9U1PyTC9WlDgfp29Y7zdwL
x7Ps+0sb0hXXU+5o93+FxI2SXVlADDFIYjWRKGJPmh5Wsn4XsoW3VW4N+gFPjnMH
cIs8Fu1wHMq7ZJ8rWDaQrygyJSQiHCYvfRqJdpVl0VQLMIw+9YCJbVycso55OFiq
BDceqUPrRckedbCd6Bk/BpwaoSMF9qgh5TWGmOiLrdkjIrIP63FvnnXmDnjnuts1
cgjydkUIK6aXTS1l2Vteu0eVztdS+OKpKjdQc59WhxmSu1AkIEy+RX5j7uETJ4bL
anH69byoYQHkc64c2pII/+Ip8ao6JRVJ+b4F7VvZ0gxD+6kZZywmqGMI9TKdPTZo
R8aEjQzk4bJ8PhlGrRR8Le3PbgWdllh+Tg88N+ZUPUIPFwG3YwXAlrh2UItYvUAB
MF8wNh5XpyrVUq9G8LqDd83hTv52DsQAhyvmp0ee2BIbit/vVWB3ctszkJejIQSG
VNeyuKIM+pMqDAidem6XJOIv52hijD5apR+HyEAvXigclrjLfGF3/f0OJQiPDfTY
tugmSsXSHtBdx4ol1GVfBBo4eUv+6iA13EwxjnCppT7ajBQfUpuUPpKL4H9DnsJU
CZZiVl6F1FmKAfnbJZhf1lAKs2HZgA/alxGutizrnTxmH9EMEwLu1P2fOU10pDin
UXr4PwDyAXI8Lg3I4FWjW7EgLC+SOUkkevQiLWyyDg8dM0h3Qr+fbGv03xQAPel5
lg4daRdiChGheYTEq83Mq/w9tHIYG/qAR8C2+ivEi3aqHwxhil0ODxVogGOETZ92
`protect END_PROTECTED
