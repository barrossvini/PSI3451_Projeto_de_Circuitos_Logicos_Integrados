`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Q4C045YnkN1aOinFClgI7GrPv/1QuvpFxL3AHcnnNPH3+xCngoFDR3p0cojROiL
2EFlv/9b1PKtoxSJAgrLZ/wq8g4b68tMU7g5ABthf+g9I8rVIXFfQDT+YJBmJTz9
8xHu9+xp5WMkDfAvh9+5Id0nywacXU2RCUHemkG1rS4srefiWQTOIfrdrBdOg4aR
iyWiwuvXvtTYPZlhG7ai5/+ad/TzdVe0pYP7l29drCSpZESQ+QO3f/LhR80o5qCZ
nxhKMlA50P/UmZgaFUY17K8ZAKCI997MvEvfpmR+djuLqevsWnywKXLzetXWoDl/
3tlIOCBovSPZhaTnZiWr5S8kKd2AjSdd68e9s/L3x5dWwiK81SeLWWANJJRT5woS
w0ngubEGeia8rmIc9hAoegwcSRPbhWsJlIcnLiV9kKSE82FM3aKahLcjstk0u8d5
h+8/isYRenCcLC9m4QUpkILVfZc+IFHGQK/Wk/KKFX1eVh9keVZHOtso2HDx2QJP
TDbk36kXxGhGhtOsfv/bBE0I5ICEngLcvFDvDrsw4+xex5Lu2Bb+sFiZVMlKkXAf
4T8ZKMsjgzKlFY82R/AOcUmshePmfl66/p7qPtvmE+C+mrvMvYCtdBcgPruBYnlz
CIo2uchuqXPDM96zqBn3veIL4SvVUizG+DZXtInz0shalC48p2yEhIZa30cD0q/N
Ip5eFyfGbPoSBlXprnQLBBOFzpFrKB+cGjoun8El73is0oUXnELpwGsX8KEu3e/w
JXJUmY00jIMaFWc3oF/bzQ==
`protect END_PROTECTED
