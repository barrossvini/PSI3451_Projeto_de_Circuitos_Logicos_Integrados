`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E4y2+xNEbviZklQD09sqtbLORfi79oT9rXxBgXm612okRrKaJK52cy92TWtf6scS
vYt7nby9A/rtQzFCRjLW3IFTnINw9YHEUhJSQ9QcszXsywzQ8/jxMFLrEabqIwy1
5fxoN+SXgDibBst9+qqkeiTrKTn3WsHl0fQuU6KOsTHTFllay8+0tBvYMLkskL1G
n1HC2Ev0ir4+KVtIriuYeW4ke3qVtubhvmcgokkhie+E4JLmu+NEmGp8Qrr84zqS
4Po+bdGFC3SgfH3YTal+WXw7Kmpzb+5OUadSS0NXRehVFlIGgffuuesX7ex1kId3
UCVa3VGbMc4v6glB0dAWtZcOgPHmDKBQbAVLX5EZ5vCVc+p8SHl7fMoo286VPhVN
6R7mPzDctZTLM/vQuvxImCtRnGDbcIYQmn/bZOx0T1/zFfMfzasUP+E2eKbNvpl5
4kokA2Yh4Z/7DMo7QakRfsPGjW7X5LXH7lBOcV5km8MA6/Nxffgqgr8m1yP+a9MP
o+MbAaNDSnpSp4bXDT4BKIvFbJdpzHcFDLXmFwMO4+1MZxzOVEj7IGCVlH14Sidq
skXay5Eg6rWq2IwTO7CpRoS3tVbDSNNc9Iubf3CqjMV64TQhhyN6PmLYWEaH1RPg
z3UZaCj8TK/CYm0GNkpJGEcXBnirXVMUl4a4ipD6kikK+4XkAaWX2L0zsPc3T0u/
ua6MWhoussUUCgXdCHOVL10CSYJF+tkzAWKsb9GINTADrXSqYGawLZfOx+kMnz6K
ZG4yWNe7W2/DUBnjCGP5FWtIdx6Dtfog4S1l2bUT76lacoHOfYc6E6MHIxJ2Z7PH
Pa5p4QxIcg1dizKSMP/ls2iyqksrKike2sIYc2n3K5DnL/4OZrFrQRNfWa43kP3a
0BBFB+BxhCD+b5++shyZKtnPStjO7WlhBH1MH9IVwig=
`protect END_PROTECTED
