`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ByVP7MmVYpxuGBzKW0bcP9bA3smHyvOhSJpK3nrQCU5uICrxufo4UC1y/E+r8F8e
nrmSH8KMTARgyldsZzhqgqr9Ej/9uIKbukGf5PzWMS+Il0JIDffMUmITo4X4p6zQ
LJ5FhRxJkPA+vvfn5PUFv2K512GFa63+WM3oM5MvJSsaHFB3/z4qC6IV++12td7w
Q+rpGHUm4PhNn5NRiUSVA9PmLLpOpoeylDr5B00svoO0EWhxABR87cGkRZuIJ2+0
BBbMVrylCUGVnmtzr/kpxw==
`protect END_PROTECTED
