`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VCDdORVNi1kU+KJkYuRcWc7TXLH+4WdkMg/kNa9F6L4eaq3FU9LnG8XUOlGFtRfG
xPlMfsUflFtHWBhI1UMTa+9PlcEcpp/qPxG/IBP88v5PlBn41EBJP9LJze/9nk4b
9b0LqYFURWLweI7DeaiXos8YI7JJ6GOa1yMtNLfJcmv5A7xW8osXr1iXTvo7iy0c
2GiA/DGuLWPXhBmOX5BVnXuZ/aA5BpgjlReF0HfkoRUStWmLoku/cM+Uv8JTT6Ct
BBe9ZISESXraY8Bpv4YSFoApEMTvY0WmuSCO4sa9FNT935UzvjkbhUMsUvM1WocM
9W1xlx5FLXf7DmhoAftnpBMsR5N58E8XRsLtvaxZoegRjTAqsdyL60y3KEPuSssF
gSZsTvO7dlYBD0i643xT9pjHvGzhqROVE51lPsttDPRdpCkMtvN6suBCwi1Rxr81
fSwTYnqv7YdlB1sfNimLCG6e46rBEU2eWIqfja6gb2uOQc4vDa/z7Yl/paR57iF5
nUrAhCYzj6k4syfrq7NGCx6tNgbIWGH1wDONQIFh+wF0oXRAXVPVH8INfgF8GLCM
RotpFe7kU0fQiAEiKnFlfflaUlVjQRdzuOuX9syGMG4uZSUAbp25dpzEBeM2InX8
v4ukSWYz5Uq1XFxy0yGvLxhgRSoGQDcP+M+Rwjjw8Otj1llWchS+PMg2mbJlF1Gm
qwoews9k+wyB+eAJH4QBFgkUeprmqiu4Z4UJx1UA8x3JlaallB8ciQuYQ0CaNm9s
9Ps+sW+ufu9o4cyZQg2rA2+StpvYQ9XXqF30tipQ26/YtYeoErFvs+do6S6nEkfw
HnZ5p22HquwhWu4IZwm4IWO601IqsTBo8Ij4ipg4J08MucJRFGXT84P+GNUd4mt+
ePj5y3zjIZOmxtBrcXYqBfP0bYgQProPPJd5ZrnjC1h5pJQ/sisLHRqz/f+0Uvow
AMawCYEjojMv7IEA1E65/Jj+qFyF3aAZd5AWWJiUwz8PGl0mmRbOin/Z5y764xGn
8NRv3+TslQqxl0VgkSzr4V/PVEFECk0yKDKzO0AMd07Elvw+QiKXmYROSqXM+7rC
Ema9igtYqXuQwaJ18/nYkqtHfvse3Pgf/AxVzUwt76T4aGjDdrlrX7dK1XTKd3Eb
O8cTffokZmb+fT3SD/BF6hg/l2Cp5AXAk84zgPOZslQi+uhAuOVqmZp4B02oQJit
qTLD+ffKvkM0+2NeV/sHW+cYXoxZ2SO1K5nsNYh3F4LzicVEnVTtztpcr5qC7S6G
7cRRr8hpXNeivEBOLhxRwNtnNNbr33ZrzZ2u8bt9r9oAGJGU2K3Kvre7vu2LHHlx
inMGFQKx3LRc2ygUkUnj7rP8NJEZLp20XcSDmF3BuBUF74efwEsimS7Rsu2jhG/E
P9Vsiq3JmwoLhmfDLz+7XLZtqfRypzO64exM7xWy+nzKbW5leRCWNSC4oxG6Cpsd
sMPvb/7Nodq7utrORWe0O+I7t4vh8wursGtMxE3DrL6YXoXlY+7us+vnjbkcBmxi
EorfCskeA7B/MaTGUkv/mXYj3IoV0LUg0HWsRXPATx7Tp6SZTcW0aNC2u8gQsoF1
NA+HfRkrSaFxy9avjsr3ez9dLwWVBdciXubhTtklWQbo6hXMcPNprGIlokVX8eKV
5zcstUgCLyAwL34g33DbIA33kpm0Dy9V4nI2xUwsKuUukU5QXinSe4PanLGXZKJs
5oKKg4gVjNMaYRF6stDSTG9cFazsF7k//bf3+8khkWBSR5+c+QHQ/73/NS65b8FW
qzpaXScm5RNGsdV4KOWBKPLfVBt5Jlahs4e4+Z5M+ec=
`protect END_PROTECTED
