`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rfKypQssGB3O3Wc2a+hNrhi1Nm87+D7qYR2rOoScDWRFvAylcmZUNbu8H6cYGKwT
ITWGOaL0eZa9BYgYgLHqBXVkQRtun9VYaueWscZ67TEKm/n/E4vcXbVwdUhKVkVD
E+B1ikV5wamdf6FNRPX4qbXYRTW1VWsc6aWlHahBLqWkIvf6K726RnnUW8xF2o2K
OFwLW/5oRxtP4gFMEjuBn/ThTcP1Y4Bpe3VgUJVk9sskoIs5fw2EF7FFi5vE823N
fpMbPW57/EblQKqkQD0e5UR205VP1mQYEk42t7ShMBtR8WkJ85AwSy7dTKX9d6RY
9/eoVuVxsvFBqbiz7W0giGpsSYBC4e1qCYia+JVlnurD4kQM007UJ8pi+pTtMmhI
4wc+DpL5PIqgiIwIDFuhx9Te+qEXeF+cPeljvlmq8Na4vprcMESv0LGwTlKMl6zL
9ppKg0FPpYnA1PKTQ5iwY7FYmuYFKF1VkskNflAiBbP5GSedBq/CS5I6tjPY/+Kf
EZdkk3+QVIPVZOt9O1nCpMp66TSh+5vYSD8aI1/UE3jzi2TpfC2oyhcFTQu8fuo6
`protect END_PROTECTED
