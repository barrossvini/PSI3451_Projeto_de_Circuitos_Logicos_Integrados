`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dfg5AYJaiNEgHpQHAmU60WsBwgZ5u3K73Lj9MTuQvrLDnq8qxxP0GEmWoDrPagOe
Mb6uTjhxoEnZPY5YcE0XPyPqwiYGIPnTvcNcrUB3NjEPWcVaiR9uu6CFx4KwoJqR
hze6q69EeKTZVGOcZZe8VpLBGZ2POg4WbxNACeHy4jBiYFvsc9vnE22Ij9puNIfM
dbPPyQk9/tQAL4n6aJhHHjDfe3WBPF2QEXQuR7S6/JoSNmhRfft5HT4oSJHg8lAt
DXpCQGHLw8bODFl1ruC7WuLS9GPDJBZcGRjR4a7uEgFqNlWYIMvoMPoOzyikbiJO
SV2HlGvmHQCbNxWGV5ABG7y8WJmOosx2XlfN4RzlA3IiaPQFqkL4iDrFWoM2ZhyZ
skCByIf7MDuzX7r7TgVBEQFL6XOUEMSJu9v/fjo1kPmXU8DiYSzUwOBg3ORIf3nn
Rm7ebgE0bgguamsDpfG6kj9EnnHwZY9Fd5Y3aVeoYn8jrE0ePLjKfU0kxx1q7brU
1VoIRPonH9vHUVTfFfOxd3l2qgdeQUbEeBY3DK5QjMgWsZpAenOxMIpsZ5d9wSIg
`protect END_PROTECTED
