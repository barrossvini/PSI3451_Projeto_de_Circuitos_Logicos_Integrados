`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UYtVBgpp6tPAlj8IsB07w23lck3SyG61zTWdU+DvmbCoz3wQ9LctS3arrjhiIyqw
rmUttbKiCprP+dSucrzkBKRiMIQ5oJ0OrbjgnM91QBq4LYmCHDTLwN/Y0YCBVApy
lWQZvu/skVahaxSDUjtOIHYEp4TKRvqa/Yz/pLnYYxyDeCvJJTahpaZFugEvdJAu
6T+rfvW6jn9NHVuMn4LEQRHwP6+184CQhvbS65AUS+4xbfxP0NlhQi6JhzTKSCVj
Zos7HvUCldoea329Z5k1GuPGaymuhLMSsWAawbo3pvq/wMmhuU0yNW+y0MSVL3ai
mD7Fe5qMbZLKuxNBfCmKxb9wlwOLZIOIi9r7vcIsuliIi0gu9xFuBpzU7b0/lSB/
Bc/Bln0G+jx7tcqsmnr08pWLQ+TbwC+QGTtzjXj1edexGWzPqzNeS8TEdTDGKG4e
urNptCU9iSCB2n5t658fkbyFUi7nrZZeUM5rBhF/JPzxxgwaEa1uAZGN4ZUtJcGD
URP8d+0YlIU8sKtgANLisxwXgdLH9MuFra/uXTZ9QnsQnMLO+kUeWxQAekNcRxdZ
bxi3wcikvZ9qVW5VeKIWDMgpN0lP6D/mAG1GgvmX9ixk91lo5jvlnyfbB9Q7zjnT
3LT3Bk24hOrDOeTzHekBKBODKCEiLvV1TnTrWmtk1OARKS2NoBlIpwhqTL0fpXC5
Y/ncePPF0yZjJcZBGxqGXqq1jwWgZxvsX5T22/DUdeIpAfXSrExJEUXR0Y8VmPQl
ttMidtY/5enFGLkvuB+cIb27wII4wECbbGAwC+id8ib8L5f2vtD4F1hJR3+BX9bF
JLbLxfpzyYtHtt7od1XUks/kfR98ELkknVYrzWd9FlzfoAQU3nu5BU67aH7zYuXh
GMTA9lFHtC650MEslxHAB+6ggCOXh13nECKIDLo6xtlnHTVGC0UYwcGyI0LaYkR2
2Y3dh1nWHlO1gVo4gxKOcEVyPj/um7VAeFh3EAn8w/FRIG/NNdJ+VPJlflB7k4+o
W9ngjSq6Jz8M+Sk5BfzzvptTUakxk8cXXou84nP0gxBIU3VbLVuPsMOnbaMpLHwh
XE+vjNXFlfdyMEtUdcnax0J5ezJS2uKPFaUoid7t65BDkD6B3aH2JHLjaDNri+LB
24de6sFLNqcllrSvN/uLeLKCjfcbPhcUAZtLIAaSSAz45zhxXxiBMON3mzhcHDid
Mdmsrd4Gnexh5UHBzSnIColvmhIE6/X0VUSJ0rh+EZgIZPafibZCF/j4Fv+BUgy7
ddDRAA29bEEiZO9/GfUR4EqjKKTCeGUZ3tQckXoUNIN0IS7kwSYjxSSOp1judusd
iOVEZp50nGy7x7kTLwTkgXR+gfrRp+5cqCTXX8zdMdO7h4e6JEkOvB3ou6M67Gl0
1q7Z4Oczp4wuL9lBsVpqycFqC03WPisIbcvfPqHIMwtm0vFBOuyiJVWLIHC3HFRf
vMpXu4/gktBvHaGgDsjEQ0k92lyQ21afK7hX/wDJ6o/IHb3GElQZ4Ih/2R0gGs9S
whlnwT7AMTy7GZDyMYZucKcrPUwpqlU/dBnEGu3nYZxo6EIOPKA6nf43aFNKtPyP
qlcLGcbkgtpx/W568AbX9fyARCfAdXN7yir00IPOm9pzz1rPbJgKiZiJpcysuTMV
kqWCqOqLAUSUJO8c0DpxTbfuwSASuD2a0WF7IA+GmCnwDEgB24gwVcw8ZrHicnm2
pHSQx1nWhmcayGuMhaG9Li9E9pu4jrDyZRbtqwzYXXoJvU/vJs70mdSY45Eaqtla
mNnpZ+aghzRi9GZhCIErijhu10nwfQQBuPeLj3kVrs8i9FvBz2d/Kacppe1kkp6J
m43VqzIw6Zdgg35Sr5Ukku83a53OiP6Nii3z0MMMHRDEmh6V2EaExfAcjhTllpnh
FmKWTxMhYmc47QDvEJzJ0LV06+97wMe1uuqpaTmB0M0113SSvMBXFAjUfrrYlSco
B7ExZz1hoFVMG8pRLzmacBfYB3mvdRaFRrrGCVBZcOe+Tk1AMDxTZNmQrS/xhhIh
PFjtPWsM7aQi4/n6D0MJlAq8bqoQtOadZEDdxpvZ68mG89r+kxsROUTpu1nwiVB6
6A6qh3ZqTOnrj1sRS1Hd9FB/9SlFfbWWRofKx5olRuz36v9BNffuYbnC573V6J90
AzCBGotGxLkoTgfh1dS6d5Qsa3msx/PmRYT3moU+OD83EqQpwIcnhzf429MPrWKP
XRY5pgqLx53U9V/Qc6LG3K371RPvMaLWMbx198tkrwTdrRnKynnWhJzj9Tx5Sc4e
Ctm1Ic7r037yCKczasVubOsfGjCQ4FLml+LylZoAVvUgv5jWiZPNpAYBr1wTEn4m
cPZMNXgvGNJxZ7OZ3zpLEx+RFiWsU95dswtDhcK7tacwULtvcM5qxK5j13Onxem9
x2HQlqFl+BUD6i73mxi1yERt/rgrq/wvqkzbVRr2O7LAk3u3mpXdHosDjw2UP0Lw
/kBsbF1DvBSyZ8knCIVGw/yPkWkAgxl4wbVM/rZbWVQgL1TZXhv7yBL0O+nnJaFq
GqJe7v4TZg6IElnmf661iDTH4MwWJ81JxOEAegYxCizwiyhNzYIin+CfIHT13RI0
5YAussD/hpQNS3mdaeCUeyMtspsmYmr6P8f9t57RFzJOSd+/tVBXooLtO1Ch9iap
fAn4YyZzmuE9ahu3xVhAKIN3NFL6XwXY4fqWCCk23wUl8Tl7In+cLmu+Lh2Gv66T
M2mfbSy/wWsGGADRsvQ+dVsKJ+mgjMQtcxLsB+N/CKMSa3/TR8+r8Rph6vmqkuaT
xB9BrKrLFsFJUAzif4eTwO1Y/u5tVHmjO0wOD+l4jSQ2QoI7+ZIVcO/kv5EtF8sE
gNzBGE+TZHZwcNZYIOhEqf9bHQKj3xCVLfSQD+vt04EaY/r4+jHal5/1+wd/zNwM
WvQuGIZxlFisPsE3zPCw3sWAyHrK7nF1g+2fBKiZTtWQTMMR1SWjPBDZfBD/7Bol
fZRsQe24Tl1WSMPszzdzx/ultvFW7SfrqlFUtNRVkYWfaQrORloazlJP+T8BOY+H
hSzTGbEzMu6+In5ug40Xn14zCwMjr55HZNW6LLsxNQTi5ek1PBGVDYSgah/ef7GE
kSDLEdZ9vkggy6vtzWZjaaLCDHtJlysRjw5+MZEsz/XHdB19/dIZA2UJw5Q14GTU
EkP1GhliWwh/ezOGPnGrKP/valVFuzjwG37CYqjKYNzMbA/4UEqkDShgiUlhrCFJ
b73sDAm4TaRT2Jq9uiYNR5X1RbWOouLJTDgNEhmvH3OE4Sdev98dPMETAOd76jjs
JWVAK2ALRVX2Dz+3m/rWgoJaOhqJVICC+WLHGqSQDD6BLnxS/Gm3aYtx2Uh2SKUx
ZuEj3Sw6n+fNyFEzwZKrDaDVNk6rs/wF1rROttH2YCocrdPH+YNFwEgPxCniJ/Wb
Ae/EKPetOjQwKNcYMgVsbb611scfGJbdzk1vPQj83PDo3oImQGNaprYZPioC0ZxB
hxzm3475fRMrMpvt2fHJ3c4l5dMXZsW1lVV0tshyAkXfp5pBMDwphwcvF4rq2/rE
vP6PayPqzOcWSub7KGstdyxHZlszdY8QeQ7uqUsKjhvNGmdjdUFwm9cBe7ELNfG7
nesJutWPJUUWLiDtRTKuC+h7OUwoBdWAekpZkI1AQw1DbLxky4xcgoe6kygAjXQc
fvsZU79uwipEvnQlY4nz1iVmPVS+QrZkkkuEXyIB1F9wsTA9vYCcG2p9TSTshYJp
+x880OADxNjW+5jFnGPRpKsi5WDN7qUryl4isSMvLP0eWYy+SXAj4xq92/4yLugy
v8r3HZV2HKzYa58kZnk9JcwDsjY8Y4sHOJXMMP/0ROVK7pGXfiSGrAJt+BIzqAbw
/GT1K/HYlA78RC4v43SGqJy+PgaQULx1nX635I1VnOWikiRfHy+MmB52svAUW2Qq
a7VtAZlaw9AR5TLyYLKHBeSpSxZNOCoXcz7AEOcgVQl1YrAPgOjv8MODl5gB3Eoc
PHdKqimfgFSN+C8Ar9MTJFxJVpzM60tkc30R3EiN/T9RyW9S4/b8hHvSrHPhk6zs
3IRNG753lcptoiE7BZPouQ311WRfQY2zf6dugvFy9Vvu3nNDzeQOP2lRN330QWMG
kZ0Yra0e9Sj6Spk5ipI7pn3/Rw1Q+KTRAH2auQUg7VuaOu5HQPfjewgUiTAjVRHV
sujaiWH6Rln7eAVKS0yqou9tzoZlkEdIm9dlmDW8Zrr6EuNcsDwl4jgS94A3JwzK
3B9uDM9nu90jKQ2rYhzerSMAgG+8plz+lQkK318mmSYnT2SdnjcprqB80I9ixFBL
tEXzTCsCkA38Zc9TsnbKaO54HvT0MnNx0MyXIfAEQhRPpMHtfJVB+FkNkAMMb042
MQIPtFPcfNLCflJj4g4j/XqwbLGWTr4hMjuCt7tvFXnxRiNVbhxHx1dDkpD3EKVu
Y6t+l6LjVvhJUi/nbJJMPFkwaf5/hyMHqD8xBcF3PO6crFxueuc90dLwVx3dbwvO
UvHra5IdA4vncV+D6DsZU89lL7UykvLdNez06Hja/0rtUcl0DbqulnqzJFoEGS29
sL4ujqjYNXKet/g6sEmmcgp2YpAc4D+2Dlj+524ZcWO4mY/c4LK9LyDFm7YLlkTU
6+Z3V8h4RnuqwMY5SzD6He6ZdMB7+EuHAylZvAD4OnL234WypthJpwe71uqwlXko
6CRc7pu2idR42i2FZp0FGT5EGBDWYAocCbAB9jpPEl+LJoowvDdD+YMncmG23l9h
0pyPhOe7htd/fsK6FNe84wPyT4FgYQN5+towhOK8uWXMxZHzZZXLSat5ueLSSQcm
WGF/pbGhgE6IT6l16etBaWSWQIpOubeAIXAyrWKLSJIiQ4p9lwl7Qx6IcHp4txJF
RyqXhE7Z/d63FBTvLIl/owHqROyq6S9IZh9IcFYfoGNdTwE4cKWTBophoUd6XfHy
Q+69rNHqiv4jQNRvJrAJ89CM/wQNumXEx8gltJplBACam3x6CUt+YMSLlmVylwev
fcnwV3lJXGaCnMGiNddOLA==
`protect END_PROTECTED
