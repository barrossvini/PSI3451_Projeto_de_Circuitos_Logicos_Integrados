`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s83XSmIw+94Nb1wWqtOW20FDiY9S0YDvssY3phFm0vsYUP3n89rq0Tnm7kSL0Gxh
z+jKxYAEPNtYOsLN0ZjAiAsLScScBdH7zKr9tRTjzA0m+uL+FGmQxrvm062mc6xB
+LDuL09ha7u4s+eL/0d3mToM2//DGc5ob7jzizRhietn6rRe/yUfjQl1yCVhqdVn
JzySLd61apP3hIQEJxs28rGyQDE+BNX7Uq3n9ksYuYfVytUNxdD8UKxSrGxG7h5y
gQcNIuhF+6BhajcpT1AEbgQ4JRWRNXerSjZvKz6cKniVTcNjFXjQXKg1KO9jNNad
5Cjg72jxMc/XXU8t65HPYPBNWWf736nWz2VUKMavnCVcOg647M7VgX0e7fS3H7dm
17eD9POR8a6UGG4aJH3gWMvo5N0sTLb60tIMYtsKpHzq+buoocTVn3sMtarv1yjt
Rz6Ml4U+dOt5ZAJHVCLHLgxvlUIS23P6t1Z81A+++5OD//f4HbVRqSh9/KzNS5q5
zGwrlmEZ4bZVLi8yxsnd/oBh892C3OlGynmE8QiUxAB9rCtr1l1NYP9UzT1sPbx2
NZ8zc88JluT/CzqPE27mfnASnYTidN/IGC3UB2KAK4rhYtrwLWDCC8FWH11Wjnyl
ic89He8w+cZAa6+0m+CU/YSxkIfs4v47aatUk4SAx5NKimLcieEqEkWhUhVzfhi3
EgK1Tzp137nLarWRa4vHjBhaw6g9OmoxomKb1Mr+91AkRtK4b7Az/md99INDxpQ0
kJ0EPyT2qoJwMNnS50WWqA==
`protect END_PROTECTED
