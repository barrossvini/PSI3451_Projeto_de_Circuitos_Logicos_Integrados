`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uv8KSCz4yCVsoau5m8yrwpEjktRauJYy4b/T1tXy/+sQ5aDL1pMB/6xBEnIZTlCZ
IotqKqqcRlfxiTzoLw0VMNVJHfZkvx+ttFOhee0tJ7W8Oq7X91V3CvZDJnv+5mAQ
1uWaiJHUhJlYXv+/LSepcq0d3ODYwz7XE/ij42BZIMdaWbPX+23NZmLs+0GsOhUq
qX8OCrWYXP8uFgvTVn370bafbdh0yPpU+kdw0jCq0zcxQWqoSUviqfHR7upgXUKk
MQxUN0HEacJNaIj/fk7rXV3i3UvbLQPSP6n9NtE9BWQ2Zdo1UmuKB4jhYA8d8Wh0
BR6012FS+OmJvk5aIqT282o+jktjUHtcodZLkVPq8w3QOfTLOyyvpa2oltFK0P6h
lIjB8MaEH1nF2j1XDAJ2rty0jCMEmILYJecfFPsn+IT3Tqe9vqvd0W5VpgHBkOsC
F0M850Yrwh1L0Zc4teSTxfp4PtUl3mvnMN6VdxmOWtci7OjyqNtSjehkUfia7qOy
xNif777RWklRhDIBdYdN5g==
`protect END_PROTECTED
