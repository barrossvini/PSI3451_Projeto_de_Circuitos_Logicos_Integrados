`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6M8y98bgTCDxm/6AyZboDpTY1vJlp3Xw1kMSxqkeWX5FJCXjLrwNTkg7IOCvFeXm
BOlSKBzPsqgsKHzbjt+olsWQ8wG0lqME8WJomNtQfBHcarIrLx5By/e2cBNO/yIo
ADM14VbrIdpPiR+IHGg057ZBXA+6A3NvKst1tjOq8yB5Iqg7MtOJT5JbtOqojoFO
d0jQioweh7+uAm4c8YSj8UasXPW5jI+dWZ59dgl/DhbzlyFZxS9S3LPHeYN0v3AP
e9KsRTNdckdbBycZIUl1xCqgjXReTX1YGwrsvj2PdGzzy7/PDBcwFahLgyqreZfK
9I0ul9A4U3tFOdRHAdVvFkX/ZpFR8KistjtJaGAQmw8538FSidC6YiLC+ibWvtES
Ff7jrvWemhVaaSWiwkz0Nldm8vEtgMptjVR2gqqakW/4t1HucLgVi+YrA3yuhg5f
9D+l4S7UCK7c4aXskfEA1XTeHJv9JvvZfZY/1UcNUOA4egOngobmvRsftYQdU2Sc
uM0lX/4CTS0FkE4bQgdbfbS1sKMdM4gpw6ivn9rWmq0YIOUAU8W2dxcNfscW7XrD
Pk6jU2n9c92I+qRn8uAQijn45JP7TH+6OXN//Zsb7JFTsmu8yYoilGUCze+dyT5o
wC+K2jmQmnlzXRLwh/cIfUT58KY0V/Sm5vn+ZUppBg+Q7083P9skx8eS2BqgosKS
AU5F/1q6Q4VSnF1itRhUEDWiX7Scn9xNIymzTSCD8qeI1D69d2cbVNZYYgzlnKGH
FAiMmaqR/3LULuObNh67EqMAwk6iUBkYm0PpvHVlhYNktszROmuC6rv+lJr1YP5F
TCT/ZUgIPuBWTdh36bHgLWasJhgfZKJr9b4ex3lHaTlX2jAtqGFo6qMSHXLrs3Jk
gl8eCjfZK9fbICvyts3VqTLUeSbnloU6WVjaTg1SACZRYy3Rx0HHfbehpdr+vcui
4WfpvlK2dz2M9JpsNrAsVua2V6IJRmEvXDSjU8MvPBxfRWsBrHASYDUk0yK9IaCZ
8CLS0tCwUUu6CY3OZDEBrlF1TrPcYP137IIy9pqMcAS6pAPHdLOfy6yv5WSNp96Z
y0FwPMaJUeichHt4RyY7omouTQkoC8hJ62SrLpBpMUfnGabUmUUzxBQiHDX0tWFY
7nRTdAmcgNeGn8Ym/V8EZ/o1G0KycvMcjuAyZTjr92wnVX1a1auuawvFml/3e36g
A9Yhsj3/iNrZ6TbaXpCYIzrCV/9K7darq0PfzMIisLO40XyHRnFT83oy5ngvVrgd
6y7cK40Tgl+gS/6H2Ha0RqIE+U0/EUIhkeQSsnCtG613uM+0io6xArC+yMI/fc4H
wr+I/AVCDsY9NNsBZ11VsJ25Wpjq0A0a9ZOxCFg8jBarMyI7b+8fHwL/Y33zuRdk
lFXvF7leGo4z7sjhyv6Zg9/DuOJx3tJw+Z0zubc0fOufTDDJa93yYfVrn+evShq4
EOpDYciJhx9IGIUu+ZhHTetVFGzW9U2h00xf/hfiYdIheXbiXct28gsQgjF7IYgo
aqUN21gRYjEZ3R8WAKrgJA==
`protect END_PROTECTED
