`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/efPtDAxAgZQt0nLex/BiR9gyfLGfSIF5d2CyTjbXy8o4uGGQ0n+pw8gWM8t/419
OIvi0ugvDl1XZi1asadUGgcI0zzrd6KjyXFuyvILQOnL+0ckj+8UN1SV2v5kqO1C
GG2AO1wA9ft0VLx243LvSqKlBJb39B+U7GtT9rpydeOCGGDX85lZki2yvEVnaLSI
geSmf3DeoWxHt1XHV6bwSToufJ6BBV1UU+wI/4d9hP3JrVSY2O0RYFnQqzrwfOpp
FLdQjchf77qpuKMsRZOjNAnLLHDOoLxbbliECwJJBGH2fhVavVRR7w4UBUykItxV
iReNu8X5Yxh61C9K+H/SrgKjMyXEouVp5KGL5G5QGyhSJzggk+6OBGiT0ncuQRUP
KDNq7amTa8/h7C8r49R6W4zGwiuUJ44sr60LGNp95Srsr4ZHvGfPtxecKnpRaguJ
`protect END_PROTECTED
