`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nKpcDJI1g3AFfGckScLdAOPZi11hHJiqZJzWxSLqkuGmiR7ZYiyZCDD5xOJCdlHm
WdR43DpEEn4WA6B6VAbft6uz4za4KAwiFmb+3OtfnxxwFKIb0v45F2n7tTwH0lM7
SHnBlv+YDADGPGNosEqu74OBX6ako1rI9qngoPhLzNtNQbM+JuuCBsBK2R68RycT
YiFUQeNUyhnSY4+6HECYk2K+oGmNEqTYYnBDWfVpcaM+1kZGoNwQXrVVsSUP5JGV
by6K6+gWWr5S1vewEIbqXVAC2pTJ3q0fOBFyNwRleXibkRwqpcuXK6N3PfgBxfXk
9/2v2P/69JT4Tbr/sbJvFh3ADqKuSCKuy9h+dhpMgT36G/qVStXFPRpvx7KCXv3l
nXFnxFKwpvvLU1uHPJ4p41dcOVK1OyghxT8Q2p1gMp7HxKyo64JABegp5f2Uml5B
cy9KAG8MC35EgotU9d5AEDVXDqjfcKzI3eUY1yOQptMYiT+80ZHfkc+mHTgiaPIz
rrTq2ubeCK1lF1RM+SUwE59o8afHNsNgX5XKtjiFLXx/YnsUBheJwfgm0vC6ChoT
8fBgFvB3bvteVWHoBtCHBZrF1oON3/3MNtpfqy9F21cW1nab8JYUHKiszQa06M3o
iEkLlWrnHuJZwjHfLj4osPAk0BbK9qUn6ahp/nm7dt9XsHTJDWzAIGcSjCmXIiVr
kkNk9ExMzV1DCqcjwCdlO3VOHKtwHj90kjqNCfrxHS5dGKmiweozh+T3HpOzcQuJ
3B7TSuEF5oLTeanJy9/MIPPAR1Ow17FUNp3kx0i7Lyr2IoHW4EKQzJGfmhKDe3kU
`protect END_PROTECTED
