`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yavLQ0cdN+wUah6aAQOyDIihuH6io0geTPrd15SzdT1fAzQshiXiHYiMQoooDWjK
oRKJ6LAJ4iUD7SyXMAjMY6N0rR875ZsIaRev8X0c8q2uZUjTbFHcxTtOgezsNTEr
A/uvtkBvSVXheZdmbvMqiHQGOvtxtU5/xvYxgMJogTxCCeYjdqxmUh/Bv9NUe/Mb
pL/2Qm6p1sNiefaN1sxTFlyikdgf3cu6ZAQDTJjmmSzJht/gD1FMuM5un2XgY3Yh
UHdxQIhGjBtA4lGYTRRbRWhEZZyVY/koB7d7FeaXhiLjSzEOwNog02at8PytHzKA
CcIg40sq1uZx8I0zhpLl4RGvRgHwA67LHAgo3EDIpRtU//wuc+RUQnHMKI/PvpbH
qy/SwyNUsc5zc9XfxTIVsTbiVPFY4MCD4iW23YS0WjESe8tIo+sMylxdLHPUC4Pe
hohRflw7MgjeK03+sHLCdZdwnZDlXQpQStNOzazfwtTXU+XODDGKtkzlXio6LyEM
mA4HPhn3VNKM0/jcPi05iYKor8Im4wMtkTQKF6vGtiB3M74pHdk6CY1E5XvglE9Q
ysxXM7JwMf8mIV+uy73WQWNzniLC9FZ1elDl68jg1tCmiw74HZsQPoGL8Nwgwr1h
mbfas415JKKFyzHPksShZ+yuLotO01rYT+iQoPEV1gFK9+MA2RXlza29iipB3VV1
Kh5wgjOF1Z5WBtedMncGCYj1ArbZxowDz+g2f2r3vgmxhIJ9/lpE3ZELZJnU/eZN
e5wguYEQjLHDFaG0dvnWOCJ01+V/QovNZUQPxcJP1izOJyyQtbwd5QC5Q0dWHCLr
eexQO/PkDIYE+JiUgryA42ZKYYPHXeKo4UY60YVZx0E0NUJCA4zlpEEV2AyIaKkm
kCJ/CbX0wsAJ0aKj5y+0OQxef9aTONlnbATGcFmOADCEcrcYUmkt6Mf2EQNvAeqG
9+qpO2bxY6K42xJBOJ5PKlJk8XMkmBcHZA1lumcN/GnLwlV8ljvTgwuKcbg8BY/6
3TnlNLC4mViLRO8Hk+M0hyMcCohKffUzEuW1t4P9DN2t6OMaYrxQjlIYJ19eV3fZ
LnBmpSIdo8FiDeBanDXmONYNOWTNeB86b6ZKBUeZ2RmoY4ikU2cSZZ239qs8dqsB
ISNm2AdwXRJF+4xc6zQwdrD6S30N3vxkZ0pBhSkEKCUHRJZi42x80WA65hglPSRF
kTPEHNmi4sPyMQ2o6TdDwxQ3UNf/403dEeq1JVkSfgdpjqfWnXXaAJBnP/2Qks11
vUwSrhgloyxohUhxzz/ieIwIyR8q1HYrtzTbLEMOryb0Zkc4mRkKCPWtP9HWgXDG
iffxaBACIgRRNjfd+yErylcFLGqbbZ5LWLZzP4fzL1pdtGhyiE3f0w3qXY577NE/
TbinK8QlcCwB/YNp+uJugzs9lF+YYdoxkfC2FIrylzezXVv6ffl+F4dbbCkhWN+m
5JlJR0Dkxy4WvHyzhbwbTMPmpcnDp4FivaTumXh4GLuwNSNMMNpgrDYzDzjGaaGC
fE3Rm2KL+JJuNTqAy85GZHIvWt+treHXuGG6lMUrPtgUwf1AYXcGcP0mYuhPTC4k
sX/PgYzg6le7tT9EqIEOvZMdydA1wBEzUdE+M2SfRWT+FejgSZ36AXlJt/ALSR2j
9acoE+X4xkMnl1JvxYAWf8FYwS0oQH90Uhl69Y4fS07KTBsIKEU2BhS75QozLnI3
XqccqchLOrdnEVOxi/cHgBtexLoRYPGOPZNFRKDw69o8ZN23zRGUCzmh9M9cSL6p
ik2rOqSHKuoyp4J+f/4nVH+PDvSmItFZJt4NjdPMO7BaGqpgdcaDHYMXWm+G6C94
cTu2VydcdOAhPiem6P5sWkpSZ+RKpzQF7r/bf39IJu46oQtt1w+fK3kB4h+7jiUz
F25shxFtaVfDQfvvBbDcDRVpjN2r1/reKeNOCw4yNjyQaJwv5hGY7BTnOJmDgYl3
hy7kKTiRCwzECf8bwefKdezs4RltDbGLEeijsMp3/i1jISUyCCtrhODQnMa+xTOj
vOlIoaklumJ/zF3pu3WHtnrMSVtVbq+ZUrJR+S1j8ExjGiuC0Kz6vb7nQEwJsvbS
uM9yLqiXYyUdSkkXy9KnS1EIAx4t407sd2vEy3dxrBrrlj1RG2ogUKHqGoDu9caY
SLr6qIx9q5nBeBpdOamTuH0rvGpIp4/z0/LylQZ2nnWX2iWx4vByXGWpgpvzqYqn
+dxHyHcgcWRs0v/gKnVzdZORfZ1jPRxzFR07YuMjnGTcy6i1wjPh4Jwc0D1LiyS5
RtejNmobneuW9GjAwMTpgp7NsPhA95k2yHTjsCOEjOU2Ck/7SHUr9NiiIi+Y9yXV
nkeFxDhpNaNKy4sBxVGNJuYHgnpedfUuu5F6Sko4FMTWwfypU5FkQAMFbFejrmcG
PKZ1WbuR25xascysavK6DCFZ0u5ilSl/j8JtksUs2pEtVOgfmBnci5T5yp+19ZW7
7yZL7wu2vkkMuTM9nOdnzLbwY7KwsanHRCv4JjO+DS0Ptd4pe198l3xYC2r0CJqh
vVL+m6T8dfKEkDzGHBvlFDrPyOfnrlNxo3Ut0HseGq4jp8xq2sYyEp3LllopH8el
4WcR8vthMDLhWRiBZAtFjDxMuWM9QmhluWpGuCKI9FNSjPSoBNA7ytbSPZLaxEQ7
v5aPIl6rcSSKQgKXduiA/h50GFIhDfB6xA2CM2ZR30xnpWG9GhXe8sYqGqig0zxy
Sta1fAhadfcGFApO5gZPowa8zfr1IE4bHcOxMB+Ol5A919tJdui+DjegcZbFxcYW
CF1EGIcLPftLr+n3clQhuDqzBx/LlmzFDf2XzhPUKU2QO+MRmlRCmaHNCl3CmNZa
0HMcoq+hc4ARtXpJ6i6ms8y87BbLI947AKnwUzBLtl2vgkbvpi0Rh0beCfmGx7aY
L1GLEY2ck8dt+3ZV3Cvv3qyzah3BBJ7DuTEh0fgoTXTDK5UUvsStIZ4KFBigvDXd
iW9Hw9zFCkDW0dEEkbvE2djGmKOvu2rxSVZusAPbKI7sX/Ry5CEMJKEn5IAk1Iqp
JBW0lYl8yltRzsqDDjhEiwBTssXh3XHLx04vO0vXwW72IJfycrMcvFTX00gREODw
eWp3o6/fkqT/c/V0XyeZRpgdau3ZOXGrSdSiLBA8BS2n1s2EZezVr9m03YxG5oh9
58yyK+ergLbfDDK1kbeJJRG7LdoMKCbgkdYvpnyeqVew05UqlmyGullIfiJEBlxX
r1JXVcULmWUwX/oO3SOklh7gVleRjyRn6DQgmHQ8EALPvqISjt5NC18dsJL7aKde
z9VZB6u618toO+wXpSe7i0GTEn0TFsP/vZxVZcrPTMvAnEd2W2rZi25sRPFNb7RS
0P6itwlWlrtlGrDT5/0fs6np7u8q6MP9k6LekPwdMPnucsRg45oxB4APmfUb6zDh
bTfmBo9tphLXx4fnM59xLKQ3lRtk2kGH8yU+zq8vrNfYnuNMujfgwmX3+dq3OMm7
D0c07GKATjaIkbRwgSjJvBlcYJLCkH3PvsCxxQ2hfEdOQgjU+rLFLe24i7nKexV9
On7WeoCuHS+EoPEc0ZOhHrafGiBFc6BCg8om+VQUDIoS+CnjghQ04tCYFTAEV2ch
WcDJ6YG2rQRoHXiJXzhj9Mmq4ngoggeY1iduafBD/24uqb36s3IeNvmBdEPHQomA
hew1torP3DKKNG9Ucf2JMe+prPQ3Gbnyxz1SlWmz5Cd75NCFD/vetnL8LqoNDBqh
Iy3OCXdnhjrQ/cn1sTZxkkniTOgsubMp7gbHvq7NDOHenkRZ2KRe3P28uWopBByz
fdcvwsJ0EJR0O4BwjmjPf4xtVtLNeVh+rkBfkLPeisKFKjKh580rin6tqSTMEbDL
S0Dea/dKkAPF4IiTMxMPcrtFTt0z4IRhGWWz4xPfqlprBwkguBJYBoyKiuxvc0sI
KqhnlSziQbW27bYaL20HNr716iErad2p/mla8wre2GtYY55+gsNIvzNRDMxgekY+
/5B0aTgX5Ii9lVkMnxE0lAPgXpwR91EQKfFvR7x3hsXQMZY5Zukmz7G25+otFVzv
XS/YTm0OJ7FjWwjhxd2WpNQyh3nf3baM3HHyNub63L2+0hOdx89ppRVm33jnrVHU
OfXdWV+YdztVfidtbZJiZ4Gqju8TCSAmfpviY49vOQ0zAXMhxEomsNBcKYCyr1X3
zUvC3romBd2G571jYCJNxQNEWQsoTvn5ykBiKbXiw21EQtqFE8UX6fgTTpj8bQR1
gNnjxD2NQoGNc/AURgbAUxgHcdgrFlTga01ICKyqcn5t/liDYB6OqDL09U+dMjqj
aiGIzIKEkdN6S9u/NPscfZjh/qMvOKT1bGjn5CZB4KtD3Kq//pjnBE+/RaQ8q/kr
vUUCAThSuc7ZnS7ZTqdMdqTNMTZ+/xToP9Opfq5bSfFRNyGIvzBBV0/U6ydQ3K9L
qzrefIZFtK2reqie579R2jAyOuddfG3XucfCx77xsknQwGKUern6lhD4suME427o
HzxH9SdMVMPjUUvTNewZzvmRzGqyla1BZUrw4+fFcOIql2Z8RM9QfZoZqVZH3TCP
JWWR87S26Fovv5K2P1GQWFOOPTJfG+E9EcV9SBM2bytLDiPaBvFuldL8X9G/4qlO
4zB16Kea8Ft9xxRF0JMmO8OzJPbiSQ2bZrfOCHcquLg+I3ZilnENYU04H1iSaXGL
4rodu8X0/B/ILlEkLsd0WNIVsqgu601udL3j3uDdHEp0TCrTbuCCr120EIitXlui
DVDik0rndYgxY/VsOU7/trQAJ421qGXH4Vecmd3hcnttGCrGlgkuExBGpakUeZFo
Z+mb4WM08nwAmi7Xh1BT2lx4c2Mi41l8KpwICBm/P6jkgXA5vXtWLJD+MbgE66FY
69RmaIxW73oKGRlO62OgwI+nDZlvff4N78H1QrDp/l7xtLslRcaxAh2zrhRP6M4u
wHTPzvnqT5yNtYqF+IqM+EqRGRSJpYuaZUz4iJVqL8BRHk5dAqEnG/cg+Pc+jIJk
xzqUh6meiP7FiMfzuLHZiLmX39n7oJTCwN8fHmRj4KhFYk0Jzh3unLUbUMn4cjdf
CbTIsSw0u006qreAWf3QeblRwvA/ZfIv0MPAVAtst+S7X37X2DDqhQju26Idk0IT
vr9ZwoykoIDbiIH36n8fW6ir8c9Kp2bQUrDHyKZkCFRuJJPY7T5d+wOm4W7zAx6A
2a6VDQIhHYi6gt0jDH1akMTlqgXeBxnF+GzC+EgXt3JwO33nQopz7jg3Fzl2DXFk
SakEKrpIY/jHKVVUiO4PQMEmrKK5+ZQBaTLBxfnjO7zpsS7oYU6EwSI88IZR8lOY
2LyjPUzDbiNUOtfKqe8hCyThqYs2fCbtMC3Zq9KHdQJT/xzZMyGIT1kFX2gO5Tsc
aupY4I209oRzCgSABDgBJd8IW9/m5EN6J274zsM+m6StNseJ0B6TlOruMKUxeNCn
6e15FaM8QsngRhh3ScRUK6V8SGcbbGgesK3OAyb9okBZPuqIkAyk32CQzLGmSqCL
EwzcUpnb4Cvvn2n7AQrbOcBYaN6IstqyFUs7+R66CxgbYgqyfbIGR+HbU2O9k+Lz
lADKbTR382id4GlovnLGPqO5xiAUMbBRuW/0pDSvw8g4RZYEG2DVOlo9+JOyl34b
mvMP3CasTgPhVeJBGdq483+TtL39EIkQ//N+TBDslPuOz2xizl3JCmwvcSLa0/tr
N8hkkjKpxgzEjkXd7NtzduDc282kroG7JNSEy4Aq121w170NZBy4aBGfrvEldLts
ItmJDbTNWWhlgVD4rL4UVgZTzfEMoXgVChp2dOCh24t0anGiCuFOqO24GHgrxXnC
wwurk9vRUY7v1UbaMzb9ujGt/ptuWAc0+w4H8FvyqzYtXcZUEFWmWLUIXM6DqxRK
dS5qsbCRRMVXu7trOIv3R/MPypyUsxz7bTO5hGlrmhw=
`protect END_PROTECTED
