`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mE9W9mwiR5GAUrZ4bQ4yqlpoFOULvG4DsDjrVRAUuYNZ9UrlYNp3crsPd0J9Kph4
tFV5AbyHW2fM8FzeF/IJPoDLzocLctkjr8C2VuNJSe/pktxMlvyUq3lxXxX/KLP4
8iYjkFVYU2Hk2PIewJYqaCSt7BFER8VO98+dWYnRbhwuc5UrXIQEREjy2NRY0uZT
k0RgahUj0E1D8oYb1tNDLLSYpYRLHl0IVHzdU0x1uEDYLEEQdppqsOZ6lo0OjrLE
Xh1CEajfDCdfThDFp05oz3ZKyweWz6YXa9Uzei+y1hfHwut49rRq1goz9GgS7zh1
Vg/ZcUogLnK8UN5vDwp26d7FtV901y+ieZ28JddmJDUQ23ny678Q3zQBlskkn69b
XLzPEjBQ83dtRrT4p8zz+gKhvZ7NL/MRUVLsHtYVAHrDMZ8jlP65LaOi9SozsAsd
0rlvSkbeAkpelHHbGrvtytx6Mvj2manHKnf4K11M/P4tvi0U9pEKiMybVsVblnbL
33GaJoUVHPUF3jU2xAi7tJxG/6zfmKwGzi/I6dgnxjHPO6fA/AKc++b044CiRk8D
E+j5/bfy/JIR9ZrZ/vK7P/so8TdMCSejBmGxVGI71SaEYfOgFqS8JQrcD8it8Ee/
Wo+qblocRRwXxNiMDHAtn5HmjX9hk5/96B8C+LtENs3i+BKCqwSNKILCH/idxH3F
0LgqMGcE+5jK7d+R/AGiL89Ip0NW7LfLSvMx5vkjpC4U0StiC1FL2JVOfloPHMGL
GzixyjNVgxYtHLWBJSMOOuI7uZHiDgMqRH35LOUaCqcPjqwyZ3BEQxYGIH4GxqI+
fcO2HwixZwwEjUESdIaBhSRI3b+4xTDYWC2GBVUWqbelkASA5dPXcPCu1FUih2im
4BYr+Yp9eNfA/sgq+oAcZIMJQ4HV2trGUOk/Far1AWzFwo8uKqJPA1bBFhVIBQSs
p18zPk6GWzTEqJU4dthkntfsoKFWDlpNyyPdErJeDpk9NNYSJuk+Tv0ERYGL2qkD
8NaZmCWpxvYAovfyE5K7/JpG/ypIFPS5+mQEWz9gPK+Adn5c9elkS7vcWsA+7nwL
Y3ZInTK6YEtaJMfCE6KBZVhtNo9KHdr24iCf2X7o+7CGt7aRegHlIjoOq9XgCeXE
2LZVS7KQSJlGHU3Ef503WOCgmbESZFurX1r1Vmp4RDBWm6Id7N4g2DVuxLUzmhka
c93h/dINFAk/Jd45CuuznkYdITbf0X7ltQErETAndP6GMJX2+fOiLHHEK4wBM6m4
Mn/17VMkmhh6qQHdDVlfF40oOT0XRuOqTRl56hpeK7NmAkEYRp/nI+MCYm5F5VR4
xsO/i7ZvU52s9Y3Ja9WyzoysVT74ITNKGSYAFdk9yOtLTvmoriJ8eGJVs4+/Jo1m
GAOtzEPmsmXt8jxiRfQxtdLKz/1cMK99tAogUM00TBVAmC6b0YVCunGcB9GucCX+
`protect END_PROTECTED
