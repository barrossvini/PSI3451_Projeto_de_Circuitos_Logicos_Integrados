`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2FgVcxuoA7fGku6hbIJm2gol6Pxi0dvZl7xu/Cqwp/ehnEwCCKAO0K5zgcAmN0N
ySnlJE3IOi+w19n/WzlwR47WZwTbPesMIXxG3kFeasYZQ9oDqIUKf8xJ9ri83SNg
1CbpTvTBxPmBWMudvZxfPJfMMyZkW18K2LsCiWKDZ9gZp3W4zuyTjC1/BMoHLB0/
LgBT9MjOlOR8Uasm7TYjX/5rOEv5mSh1XN+vhHehsw7NUiVjRX085VxQNFfqS/tR
k7dlISl5+TEno7l5A37S1x08KtPOyUITnOmaCJ5+hLeyZnCPVp+4YlpE3tHrTmYS
g9+B88NToiq1w0b+vvj07HASebNlzQQvgU7P8nSigv+HW7sf0Ffv2I3o9OjJwHw0
hhmu36FgjTN9mqaKm2ZyejScB5GDufb+9x2wJSB7NfBBgRxA19Sl6qHQsC0nvA3Z
kgQIGiBHX1+FeiJEBsNXR+muhjc/PuE4OCpbb+xV3OuoXZmnpVtvrsvx1fmlBbWz
WY6NDio/6yIEVix5Db9TJe6f6Z0hbFNfZx9hYtSdq0MfIZUrgekMPzzdl8ijbk9X
ZE/lw8FYYjSozU83C+QMiNci438P8BLNNkUgRK/K4bfpjdcqyX/o0l905osnxIuG
XfOj1cvtDPf/8Za35p525Yc7uolYS5yi5ye95b9twiWbdySLV1wi6aW7cjcomQkw
ZbI4ejnz/tSG7pwtzgupABEWRz1fatn3xWFxLeBgDt4DCrZBRDWHQr0L6oSF4jmR
JP0l6e4SODG3bNrIwvd45cYdPjrG8uyi4PPjzNQ0oHz5ExoAL8Jf+mURq+3iir+J
i7aVRRtzVmUie4zARuKOeXlajvbnhYSqQNhRh2FNG2Dm70PPsqbm4yNpfPbsIyDH
1TA+M5RNaapraJn/GiF5LTYgPBk9EKlwv8IYfyUiqZvfTZaT1hEEXkB8JYz2cOj0
rvHHIypZIW8ijpj0uusrPAmO+qU3rcLIkRmStqBfER8ZBEqPNCNqH+wLeZ9OtqB+
+PmTk3uEftyk/VaznmsbpjfQ0lt3sml45nxtQ0OGsg5kgcqaaLYowXLmpS0EvK2G
`protect END_PROTECTED
