`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Mxn5AqL7AkebfcB+Du1xdi5pRl0F9Yt1VpADst1OPn3t1dPDW6TlNcmtYZ5d3AC
5K0YxffrnBeKrqamXSl/3BD2kqwKVYQw782e2VftpAf5DkDjsuV+v8ceX85jwFxT
nqE1q1GvTSgrjCPSKQEaZFRhytSNfrK8cIf5i9oYbhnrQvqB15WJ1nPSGxTkts6Q
2/vXHxvzCEeANShOJAk3D0QvuVeMooUFwsKJUUBz1JZh+Av+YQiHzh1fn/ibdWbe
VCedJElB3nGi1s0ch1rVOtQN5+i9yIoRar0NqwdVJsBbEZUf2IQCUIpM1bVtTZI0
ICpw4662mEAmXFltYGTUOsw4gQf62VhBaj6bux065zpI0oqZRoWm84/cEFU5+/qL
zqKofrA0svUWRRbCdInOW4HBh5zspNoICzEXVvhLzkz+uvU+EgkbnyRGiW+pDAvz
7hm2JJVwQ+D8utbw5WoXakJjbKIzKaIG1+g+zSMX0zzrOnvsrWMa/kVvWmdUJMs5
ladbahDSVyBV47LW6s8+edsj6d7btRcZN+n6Vxpj+x0gBB4i5tvaOuYIp9yXtN9F
wvq93rA50lTMN9NrJyl9C+MODftnRviLxpyaB5hvxRTxyfOrUakMBYlOYBXnQo73
PdwAeC19DWZpm1QiLmjNyR+2dHQxSdX6Qm2izat+uKHVwjSZ47QgO0Gz7OBtPwBC
f41fbGtheGzu1zR9NEKrCdyspBPGHTFcEczFVyKwI2rHTYQbjmGqxreLZsDrdXry
zPlPBZPtSd6ys1g3H/F4FQNGEtCXO/9SF8aKSOMVkGvQgAHDQ/lg5rj04qg0o1I5
BGoid+Nu3qTpt6mmXdoJWoSrsck48I/22LsRiSyGTA0M5ogplsGYVvS0CBqTYely
y0e48S5woorPOy7JbC/FG8R0fmwNEbnD5s4Nh1uh5/iY1fwN5YgQLas4qrczK47M
JMocZK5ShX0QmY88mPSzw0ObxrGeZKWhLHd2HFVTsjt4/UKIYsMpeN1x/1atoI/v
wqzsbsDV3lK02sQknMK1Qb5QihNCLBRpKW/m5O5bAB0=
`protect END_PROTECTED
