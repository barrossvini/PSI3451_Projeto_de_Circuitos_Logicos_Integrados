`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwWpMrJJiTrJFSJc874VNP26brbS8t/IFVGd5qrnCyU3cCHPmKfCLiddfLU6nqF4
kOmBcanZMSWPMKhJve2UAvANvedZyxXIwi6oEdulqw8GqpbXwFUiThWbkAm9hZOz
pXdzLRlT9V8NKHvXly3kRpp4avilrHHkeoXSV4zhBrvRYMRHKGnEE+U295NUEmJ2
TCteDxuiZgrAHv1b2mE9yqJkkVNsX7io2GdkZsRn69woX8/K4UnL0m2GRzr12pYY
tSpX+PMDvYwyn5nQGgyJtMnaZCyiXlGC9M6jlbkJ6wMhLDTG0j2+2lBHO0bzofP2
Q9j0ye+d8Z8ZsNZQVoipwE49NtPS3SWR92qCNnaeCIs0qx6qC0DPgLMo8syagAYx
SAOMN5uw6WV0JbW2G+9N/J5Ls0nds1uPSHxjq7Il3LLpR6HulJmXnV7Vsz4/1hOD
sNGfmR1ytGzQ4HCUxnNCi4UCdwXCSCGWah7kRkp+chFvSrAZL9bpjZKPLcOLaqpP
YAjXv+8CX+K+rx8j2NsPcENUKO8nfMd18WPiXejO9pHnLXWOUrLy7p8ubb8kS3LH
qcvVAy2ZFVYSnnvdZIAlwP7nrutchRZFKBkL1FUaP6J0f3mECG7Ybvd6nbNPwDuj
gu2nT7cU79e6k32NAbdS802ffnXpzoROEfT9e9CtkmN73nkaN1gQBLNjRkKMb8Kg
BbHCJVwm6WnWDn7duEmlbpmOytoogEu9HpzvU3Tu36uBMCX/tr93u/GppP9uUplO
FY7LeN9vdDPGUeM2BCkPOgbeJDLGgO0Ojzcj8dbCjGwwr+wFzI0OsZZskZ8cRM19
ArM8vT4RSQtCKj7jvugVU6cya1vZJKGEEKFK3t0yOsYvRRjaLJH9Gk35dW16S4qX
YvC6xKiLdnEwYZse/GunVGaqIsmVkAPYf1ZjVIqixC8zROhH72ddRcitLnrw3/U9
lQrn3/Mrx2RmUuWw0oTP29FYEi+sO6SgGIdVDLqnOQ3IHDrO673nH5OWEKc9u3dK
XZcMZ2m6gtnm0uuyWS7YoCle9B0z+L7tTX3xVJge1PoVjAuodpiOb1Z3VcptUoty
QemOdOCplqNU2rgsVKqzFTtQWTtRqv9+uTOBPNUI25jEKQYYDGvuGtPrwRDgyzoe
Zb3LDw2SnA8BOzElcvQqdcM/aeDnQAFPZSxo5NxQtLxrmyLPDk45LHPzaayG/EQ9
7cG0fUHs3/PCQeJnYk2pyKpigfykEdPE0gtG2kqSE3FRhXxA4gKrpIV2Aap1Wpg/
`protect END_PROTECTED
