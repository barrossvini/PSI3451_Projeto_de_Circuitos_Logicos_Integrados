`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HwtG4KyH9kMYnsySxZoiUBYpsRIf/2a3G74aztAFL7niLLrs3ySSzy5aNuOCYlXo
reh2rPYrIiSH2CgZPR5haubYGDiHKKkddHKK8h31MM5rPiqwoAovnYdtUPCg2O3N
X3q7WKsoj2qbGuqOaa2ZFdAO5zbMQ4PcS3jxQEjQxJi6KrMREKY67CPkmiLIvCSZ
rro20AOelSI2suIqKgkuTSVo+HB0UjyDDJ9rE2Cf3jQStAm3nT0yjVbWkjgq4ppd
tg3EgGLcyh16SP+4YlJ8o8mzY0W3pQQ5fNFsRzZo5wuczCacvdrS2z+5w9VD5eDL
g6Igf91ib3hKRmcAmZS5Omni2DWG9pQv2Zwv+dOdh/bgW3Bc41btPclGeabbLfrJ
j9dQIQkuARdwjp+Z06yyHv/HCsoUoS7l9qgAjrWjyA3zysy4LOtpm2809FxVXirB
JC9Xcplt0mfDc6ZSi/BUttuDiTVwTiXfr+M9nXNCCCNaonUPQ6BfNv3uJ3Mvcqx7
F5z+cRsA/4Z1XJVn+VI1uJltJ1DhHT2prabUMCR0pX7EW8akOJ3ePT5nuoLSw2+2
T0k4qKsj6NxeLzjVLeNxRI7gXeS2D4X+ifmt4uCEOvpnMdlN4WS71PeplLWgMmzA
kfAmp+r2GczMeernpe/N/t0TDi7ZPcnePDN+zvppV84fPXWob7MW55+xYeANelIv
amGIr29RCM6rO1zaMwMA9FZsrV1rNblMq8BrDfp05HuTtKApSiL/cSYUxl+Q7Gjp
2VATN3ClmlaIv0mNYYVBHnA8ubipn9ll77TTUdSslbayhlwyY8uEgRW+p6hMMXnn
Qap7BKG6HEnAVSiPPh0yu1Kc1royaOB5PmMaP7ubtzlHSY30MQTpgvDEDZHzgVde
8FFl+FazlxU2QfgzghZms8EGAgZI9IA07apoW/cNlmROtxVsmaBo2JVkVDH9aOU6
/rii5ao6Gcy4IuyNcN2Kxd+jIvQZ+sfPF0AtTzc4RNvzwta9UavibZIt1O83Q+tL
sdwE14ambhMV+HhZT0PQ2lzfcNPFtMug+f42OI1WVkc=
`protect END_PROTECTED
