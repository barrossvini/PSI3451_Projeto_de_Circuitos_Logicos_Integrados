`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJAJg6M9e2+INjwnC/foLD4Aop1OX4aANsfb9FfVtznLPdp8db02Enpz2qs31Wh5
8V4G6Ju+lNoKh7peKsf8/AJFzlgzpOC1pb8VnUvYg75MvFJVB8qNHGnxoQfnSNXG
CNkMz0TJn52Kxl2VeRkIT3cj/NDBFPOt+Er3M2uiiAEUohjbYfnKxopKfLVMljLe
QQmEAACJOCEA4KCHzNcopU/niTX3kKy7YE56QsXtulYU/BUfya2JWot3VRMcycBH
fBiOCGF+wK8KL43LzoD++4FnhNJ2Dinh4tIkp6iZevhVpMtEgMaoIKwUzHkLnpxv
LGtKGiHw5gyEWH5nFOxnPhsa8UQ06eQD3PzjTNfCHtpZnEkEXI9JnAqPpxEc/OCM
+Jq1fbWsQijJVIP7dmXyCJZ0KDyzkRll4E532tKHWHtuE0g3Jma6cQIH3FCO6sWD
oxIY+59mUe08zIOe9IMQdMDou//YuBTRH15TnnUp+vsDDt0/QKstRoFDgNJkiLtG
uYumxylE5YzHdn7nRK10h95Om/QpODX2YUQCRVooMi23ioNy1ulDejKFWnghwZc7
1aqEHuViPCQqvMiUkT77Tp0KP6PMgJR3kpJSQqJweGctcsnDVKa25rAJnjT5Z6Bo
jHEIAxVACSf//56/3Wj6ezXUqATRXHkgCU0xQ8RwtZVf5I6eWD+qz8XyCF9XV3gI
QT06A3FJ8AemO/KHc02m/zSl6Yfr9mmhu+YIgVIXVyAMKyxLFwyvct2behoQ7pem
yt0K033uBcXijFJNDvtpIRVkUcLCxpmZ8P8RbyqrbLvE17rq4rptIOGxXQv6BLY4
`protect END_PROTECTED
