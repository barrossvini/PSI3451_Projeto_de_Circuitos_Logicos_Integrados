`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
58uvy1yC2yn+vv/ZY+EJ6O+YVAhOKBzFnVJ5qAxBE2OOR+tAqXAgaPXjIzLQJG81
+q7xToBuxpho21UpE6NUXk1gRza1/pTYBv0FJfPPrGwRdsnfzqsjt4JZR5tsSNUX
3k67E/HdLdShaPOU8W41pkd4wn/6vUunfs2rt7+0WzSpfGEzmMaiuIMO9CNZ1KvE
VKLv+kSxwyg5y4bGjSI6naX2nNvHTOMIez/jMCVbPzlh0hoijZ3ufUwbLI/umsCU
BTGrFtuehhB5nGsbdeQKnanDqSbbsflT/GvAsyvc+CpTTSPUpYANUAB7x8eTLG1m
/TXveS0yjk3XztznQEeQxXr8kLgCuIY2ys/vHpdB0xbIKNVn46V8x2e2aNAZFM4F
zlZDQXfCQxRIhZuFzxcpbwN0Na+Z0V/V6zG50A5XMXwnHyqePsJM+Aj1cOShYStd
R7gRDZ7ScIKWn62mBp9HtTlGKLtYmzgru33DJAXU1XDkSFx3d/IMK6sWWzyBL8vi
MFE77otitvvc0N/ktA+usWdP8eCbFmk658s9dDlR0HdqRyZk49xFUlWnxAdWfsz1
qD59+pjDkmO+Ye6YYz0pvAZA0ywnkopwtm+UozHWacf7li4zci6d0/hobZATdGST
02ayzXZv4CrXfyeO6E0JxQztb+ug26g9oJeYHT+gbo70paQ9dgyTfK0bKyDouYgX
VAV/ccsyyJDNXTma+r6hpEJa6sbv993+g7hoOvB4ERPNBbW9tz0H8bX9pNfRYmVk
U3q1afnWwDyG7h1/5ic4Ij4PuYY2wea0qlA6FkAsHQpr4kka1S2PYinFV/8Gsfyd
Y3Z95ajtYE2nEPqgfCF3MmXMcrCI7H5rN6HnXuubrO+5qJozzZbWzKWCRTA6i6Gy
bPXR2bqonmvehWElFh4JZZyxjXjN/Fxvn9SxxQwVWwIhoWDcbg3RdkuusKSppmLm
u7Yo79LUactEeQIKjh3IOYZnUzoJuGfPtLvsmCymUP2vk2SNs1jb/tDCKkOi0Phz
oC3s8UBCT5QLGWH9D/z72AQLL4v2hCutF9W2YLkjAYASSHxelleRj4o1if7p3qSV
smsiJQQd5jxlRX4jB7oWHiXDp+UnXd8HIXXY5HD3OOmnuL3ZPmLOPAjyZn+kWvX9
gJcitdtKzMW7npgAVRhqT+VD1PyCupGyN4QHDoc+pz3l+Rsg4aBMgSB3ED3fVF51
T4EV0NaRaxG/yy7V/BlxuPLksx86L/RRQGW+es9mqRFODCvI8Agz+vXsY9siyqAd
WuPIFNhqTetYGuQ9RXO3ThQ4CKX0s5yhalzNtGNgxBmPWk94YomFhKQIdqzl+mc+
RTRRv5+7PXXA9OiN8Nv/y3uK+jrz/KBRkKDYO42Yx3oFsYJpBVPmuIXBZ82YlKp6
eBMvzi+7500APT0KWLGcEO72BjtIUUFQvm3L0/JBKHuScpWL8OYlyWVSpj8Txm/9
QbqGgSS5/ZkzydrB/J0nC050wuPKu40u/jIwfJY4MkYZCWPf8fvLhlBCNxWSI+15
9P9J+A0aWzlggYKn0XOAuG5MH+RaU0h9nXXY3rIxS9ARGWSl2CkEmiJlwzcN0M3W
Rpljl4AUKCQLNVbgY+eIckt/PWIFqBXNx6YVJ5mnW3HsgIOymUGN3MCuknwY0SxB
HlRviZYFs+UphYUzok7Y+OdWiJVDkXNrcxX46m8lqEtlRGY47Zjgvk6hbCVznDF3
LpKBPHr4JFTx3B7y2k0xP6lbCs3lIxCzkXV8lwApOndf0rEJ2uGQ2R/P0UxXoDYj
gq1SFjqiVRTS45gVLt82sTsIDBhDWx2cs1rdFt9o8YnxHbXvl6rpPHwHHTjnswYp
O4rfv3Yr9xWQjLUXM54jx4uRAPCMSCXDykOcrF2B9oAFE7XEcoZfFVCw1EUoAl0z
ht1gbasbCGJ6jF451g15H3fpBl3zGnpMUauCccq8xsiDSWBRiv8rWkUDowOaaoPE
Jkm/OdDalos8svEztcEaPd1N8QdyjKq3Ge1ZyFu/IWZ677SNym8ERtFyXnp4WLAq
KaiTLyUrvNIVcM1LpYkCN1BEABrGHyHHzAnc+rTzg5X9k+Jj3H5ArPg5isXYje8j
gABUw+Aq+03Dz/RApqpM0DThtdOi7rKuisofU1kO5zo7MBNdUpm77kTtIOybCEpB
GdSZdraeYJkDp0gjLegtiZ9LFLXTpYuwUnPl0zUPeH/Alf+jUzwOPpcVpuRfshHO
L3BXUa1xp2uiDnj6Xg/svjedv5l0Ti5UdHMSFr51g1NKM+gDe4gcGbP4Kyi/y7tk
FBnC2yoDTPncUi+q/zLTwhfYc5GM0a7M4S3nToQy48Ql8haZO3cuiTMFmw/CTCvG
oyQa2IE4+ezxun4tAEvyKao3lan/j0Lx7vdohApFnR7tzJS7uE5JF5v5DXP/bzph
nxvj+By4aHhsnX4Mg4gGb86StvillwxpMzZ3hVqiUdQwTGb3Iw/xhC8+32+KTq2v
H7M3hr0Rg7UTfD1NpRFyo0i+g/Av8CgKdvdxF+fEtLU=
`protect END_PROTECTED
