`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpUXUb6iT3grBcv7iYCKAUBZVeAhaTzdPi6YErPBIeMXZ0o0X30y4z/U7CNg3OmG
DSICjRrmEWOl9tQOmLuWUpt8rO9JfGQug8RMqfgFitB+DFxAljFeJUBehNpSl2ZY
wL0WCR4TVMfj6d0dY0l4CR14J9mNNn/71fXJJGxlWR8vhbda21rTY+g4P1kNqp5T
mPc9OAygfrJuhfA2vtBRUBQ+/m/yPQiS+E04FnKIqFnyy9FBZ79U6tJ5Ei1RUX0h
rnrEIfyM9FaTKgWtZEia1F9/amdL0FWLyLr/ecJj9Nx4fj2yaC6+IVMWVH+6yOZp
eWu3tuza0K5RyvnO1shcaC+RLirlPo5Hc/doXPQbc8uu/FXgmNof0fe42u85kedE
iALP4wzvUiVVMqQt/nHyOKHVHldwIiNP2dZpE7DoN7KEoGeLQZcr9ehtB7txNu9J
xi6C5n6+fvasxjIA2/5pWuBFPKuZ0N+ju3dw94lIIt75myNoiP+odbr4I8MHNxqT
VwvK8wsrvHFhRWX5H1cl9IsYnaLAreRqLW+Nknd+Nsi/xlYSN+axltmvvz8VjByy
vhr1dv+SMyT7FqFubQHZNY59GedM9vEtnDxdNewAp9DNxjQsGlHUfq7arjWNan/E
xfrgfwl5ij9qoAQXErllP/cZ27kabJA3xajWKpf1sqrFnD4B+r324hCZtwVz4Q3u
oK8Rrm3ZmKnBoZiuZWPMpD0kufPK8Lphb3mOkO2jARWHiHEP7kdg9tXZrDvlTxjm
tcoQk2wwJMee4cqISvxoOJ1VLofSpKGbTi/4hvfVe04YbYsHe+15w/3FZ7k7wM7a
oh8mDOxUbtXraIdZdGv3bJ8bFwpU87rJJf3UEfLS04IVxL23d5+RsFTFxpCYFiCd
3eKFiNTDRhJ4HL09DUouVS3E0r0z4znIv/AQmavo/8wHWy0mkbFQY1P0+kleqe9/
`protect END_PROTECTED
