`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H0MQnI7Gj/lErlNRgM2iZjT41kbGNBtBM3WEoHD7PM0cGAS3uvHyIZKxkY9L7RDU
ok1Usl0czgfjULjV0l5/Djw4KXE4pgV+k/fn1wJdfu8sC9/vf/epYi077FzbVNPK
KfPdn8LKoLDRp8jLixMoTS4fpz2VQpI0hJNG3EL6vlXaFhe3B2njGzPlZAPxDae+
4HPJEP5XpnoUov7HAl5ORkY5I8rEz/w5lwEyIliyB1+QW6gHR9yBkKJl1JJN1t1n
nfOIkSfGqYKC7aniwOW5D1qV/DugVTB/LUaJdUQDeMB48BWE61wI750Gr8NR2Zs8
K3QZbPdwIo+sZhEbYLuWYQjy9kcopeYK3rx5F44/i0IuvJ4np3eBQW2pjm4C6ZCw
aAMeAPe9SUkUFqpHEZ+30zsK4VRCmgGkDWTlNZ4FLwairCd1m/I2z74xCdcHjyv4
z9QP2OzP1ZxCkJq9ZiZ6kg1Bydr576PoQ/LKpqcoZqXzK05fbUrorgNniSDYIozT
EmnuK2F7Vvi7I4BVz+ahi8wRnwqdRX2iCm6pe6CCQ8/Rqc4ZXUwHo6yDlGgx1erG
6k52bRGgELddqWcvrmI5UT0+dzHVrnTgxJHyu833rQ6k2aXVV7Xf62/7Zm6GIfC9
X1NFUTl0O2h6qGCq/lHEyoHDowplNe/oFU9epRM+GJdYl/k51lpxLE5Kvm9MXmlS
VwZFysXr/n7yEN6qV6G7NRBGFMfqXN1KYtNakd1M5gMw8pNkRmi+8Kiwwtz5ac0A
5Jnm6SagTXgIoY/Vgtps3sT3vjw5VooDpNgL2OdwK6P4YpzSN26g3PARnTaBJpLr
Gq3gWjJ/9AjeHNIz2yZJy94UjdFMq1ho0wh+MbM2ARdP4CLMm9uh3T2S3SYY3Zcx
`protect END_PROTECTED
