`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qBFYJ6Ul++8a04lZLDsLpPOnUVYiK8kDTq/clKm+61VZASKAQzPX1Af1HB614y0+
gv2gvfc7kmlJYcZD14f9k+QnDdv31FobAuYuImLttpx7YJJiPFwTNR2lJ+LmCso9
ZfjfD+V0eiEi8LpPLxLSe6Smdb74/yL/OH8xlFtjrZAJGENZWZ1hEoTyBM48jzG1
xHcePuR1aQMJ4aitAKPGj3MzQFptjheqxp3eUnA87nTSG4yQIoJns+gTcR1+8Kmn
V09aoWk7biBcVdo9nO3Os/21xw+zbGzxCsuNvA/K1eZBbE/OEfy+2jtxVU7IKEIS
4Cqr7ByX0f4JBkB/F6B5bIL7DZiO+nssEZWBPZouFnHexrer8ev/wq0OPVdBeROP
oCd6/Un43BtwbbPBwzXNLYT78iw2krA96HyGZbOqdvW6euupdDz0ZbkxRGaghE1M
A76yNODDMulrqV1nzoByYVzN3m8OQZyA59oD1RRmnit09BhrG9j1h+0CImtDPKDQ
QL2nQo2p50LJ4m5868sJU4XO8fCnVafIK2WLcgKlIY9pr9v+1rE6yIINP0zLOhRt
Ire6bm4hFq1Lj/KVzvuJyqQOmzBmp52OqKvV+uyRW0o5foUl/8IrtPGFU9z5eAZt
SvzCeLgA/vMSVFeg8viE0YmtVpKYxOIfp8DHCVTVXvXqrDF1QnB8ImqO8muQdki9
Y1133kNYSWnIzbOzFtdU0tFN2V4ku0K4kE3aOgwFx/GJ/D3VZxH9hwrDXoiOsEg0
NrZKBbpVU5ppasEzqr0xFJEEDHwPmRWNAlqXpFmIQf6ooUQbTfS9ZLLr/hPM2En+
J4Rjgs3Vu+zJz1QJ1YCMfJ3vUnzsXjVp8cmuiE2QI9U9p/hx4ZPyaNGciTpI84o/
HkoMdliJgDuhukGaTFrpBjq9P/hmhVWWuuSTnodSO+/TFpwIJvT5mT6QFDzoPLo7
m4XXnJst/cybJW/8KExR/XjDu6Kdd6on2AaPAttUbGB1w+uyMRo5zNRB8qVrJmVU
q3gq6jJ+mc6k074bIEQfZfxJk+k0tUlVSh5uGHIvStOTDADN22i3U3aOE406E28N
LrAFJ5IGncSkQJqdZOVV5TB3QIlI9LZfqRH9FExteLOgEd+PTu2Q855Mp/q+Z61o
5jRM23tOMZ0NmmYlLEIxQ3abEF+s6hYB6PLgPZ2uqj2pb8qlt2W8ba2vtWbcwk6s
nXb+hjsAWyx0kitFVmq7iKBC2kRRmfUDFSfG/goj9IVcRrK2wUjW/B+YAfEBz6tx
YZlVrSyg+4Klil7w/DtfmTtZpgWQoSBOp07/IAcd+tjpSmxpHUk825MjuIWaJNJ8
OddtMwz7lQ+JCOMnl0gm/+fGkiXt0gvfp8uxdqEvlUJQFYKg3G9wjwRGR8hfaEh3
neR/eaTH4w/QsmYPccCzTaGyEMDhb5lmaufJ569+9fVg4TqoDIVcHuIl8TGgk3DC
kZOq71w+z4X7ciu3ZNs75MEc9YsCwrj8U0o+P7lDdbxTxPrSLQYA4v/vNkxWwwbV
NNsHpaDUJyvi9k9RKWnUR+yalFGM9+EvebpdbDqLyb4Ni3QTTi38t69FJt9bn1zn
45lF0w9XGU0LPyUOuIeFlqUY60KvLpMeNWNwWZzT9psJmka85ZQfPVuI2euwMx/4
8tRqHhft4uF1aGBxBSLmfTubACSZKrOxF1ZuJJ3MA4Eajtulqvdni9HqB4+uGbet
tVj/6Tg/ko3H6LaqGsh5jra3+dfzSU5T+yfBIj2sM5EVwx3luActK7tzBO7pfXjo
eTEKNFHw07JWcQrapYJCUTPO4G/QQjaf5mT08n6MgRJFuVV18vlh4QQMbYur+r/f
HNR3SZlEWLccCgICU9jNySZ27jtVqBjgdMDwNvSuDBUxp62ZC0MHsjazkc5n+8Ur
Obk5PcFxrLQQjvvAuXOYh+isKnFLZKzfs79u1w/rVmeDYxSsf3ob4UICLm9GleN+
GBpo1PMlXRkM0QmjtFKLq6fSe8RQ9jEe6QON1AOovxlwL4Ezmm0JQCePIOU8qVcK
R0NOd2JZtXA/jYJtHx7KUtI/hhr67KPz3oEtEZNPz49viIaT8/Eh7IgKsBmo1BLC
nhTIOJO7HRdMcHRrnXjXkqwhTgWjTWCEPLulmOyrq5Qzq/o9Pk/YmbJOl6efV6Lt
XF57V859QECM+czhixZ1GTIuF+P0TLtBBqFRKYW6u7oQDN4hKuolVqE2C3L1pXnz
4nE2lgDQ22neen+L7lrhqHoZFigQ6BWHgTXWAQlsVqoTuxQ69v8v+/1dh1B/mrvy
+BE+v8JevvB3yy+mpCxzlhibP706jDXsCqsJpof/5qvY0cqNy7T8iT6nOgyLrtHy
euL1L/wP6maouLZXmwtIPpnQxMB5gWxE2ANKqJvCv0Sj7Spwkh504QrzpV0dg2TH
XbQ5lB0R0S6gqzRPGx08z6cl5J6SHSu9j5RMBLdprOuOHyg7xsUihknWTWFvnIC6
COUDFZnJTyzwLkDbL2zaJI9gi1Z14qUX/6QmgKuRiFlXL8F/juzTzJciFXiYmJya
/bTzn39ZPWMrjDJY6WEiiHVlcsNFt1VPrZD3vkm/TV1lQBKzNwYAmtrz0xstQYaw
sDPZHFkEviX9iEHuZVmIqtn0HKODzH3AaL2l1oOqY60wN8xw7gZbUjx08D3yZ7iH
R6SMdmsEyu+qrzuwsycaM7hIfuBrKJDPZ6C4XrKNNuIFvmEUCB+jhTPH9Asz2Ftu
f1AXMQbGjas/YomwxGIA4GwjWhZ3Jw4g7FqY5Sp5NbP1uHi1HubSQOY47rdQofDn
O+6+JNeZUetI+5lDTTdbKW1nxxutjFEqgDHw38CgROsOLIgsQYpfZPKYQ5i3rKxD
3BzlC8Cmxs6CWhpcDJHC2Rvacu4GW8TqmHXH1EmX2k8vKUx2P/7XKx8msJe4997Z
rQDJOcH+whEpCOsIFdvuK5lKxT+5o2HUjwWvO9yWaptbDs8cr2xli6uZnPhGydyK
kT/e7/yhyJk4dDIeRoK2THTPNmdlqi61Z2FjhF/uGCC65HPsljyeXb7LTJjdggwT
bRfi5hoEaEg8mMf/5JoW34YDsCR482VrbJ65vGqi5ksnmeH/XfFirwMsjvSZAbLQ
1ZXKrPuEtJA0z4VAjL/ib4Pep+eC5/HYwS7HRf6j7hgt1Svpcm+dFhpHjea8q5CZ
e0SpUXpsCgQh0vtW0VuHiYX7sKEW9KoMm6q6cMGsXLXwLS2pNXO3sk/l8MheSIv+
fV02dGcqtSQ7jovPbDGOS6vxnI4p6jsZMFB7um13W5wcc3UY51HKNQeltvyxoNaK
7mC/RNajT+b9i3MINPQz2+Ey0hgeScY/5ataQq4icnwNofZ1yDoTHKFf+gtsgibc
0C8MbYh82gW+suv9WTRsXSNXT4qAyxPoDHcgKmIhFMxtdpRSL6FzZ2j+jjl3F2AJ
w3MkCy26wIEafdHEg1oK20qE1+EJf2GYZO0e/JeBaD4rpUQWa45uhJcVqVu2q8Vw
cZPn7Bu7w9ei6c7dk1m9f+kULX0BpQiAZV4aDbfMqAfL5T0PJEPua7sK7d+dtBwN
kWPMiOah4rZDLS7NGfkt6SGO2iaEzD640PyHP/3c/xNUD4HoFWnZ1o5slDNJa6ck
ULb/w+Tx5+EN/FEq2iEGspHzZM5+ED0TF3E89dJ8U6bbEeS6asv5B3O54WtvblNT
Q2x9TtFNG4czqmdL9S9rVSgUmEf8VtpurdG9MZJgJjlWSiAmhxq0V+MC8xVsT/Gj
3MZWQOxHVzwnbJxj7RhczGyDC32Uu7pedfSZxdziW2KIJygysu0fjTx07mECjiV8
F0OBGBUxrj+TCzpZfjZ/OUQYqF9qOm1mZkgGu8W3FJGtc81yIeGLAiyRCOm10M08
3vQ9j7+q9tfCihcrE8aBiY1wUk3oZS0/xUrstgrr8Nj70YAnp2nvAg/uqrKOrBSr
ANgDDnz35m1QjIayf+8sYvz2hZoCQtb+hay/00210TeQ2SAj6T1YqlcVTbUxpimG
QO86F/mIeNyM92Kr6k84VO/VxCp+vmSmZrwRLV0S6it9eQJ9qJRlfTKh9w/bh3WE
nhLY41HQkBSZajUzByKSYdaWLUuFC9r3jqTRdodPgvCez/NeIanNInwXHwM0W9NF
ZFiFWjqwmua64iAUvboYXDd/hrLAs+G+wE8iyawlZ6kv3s/L53mfaOaXZwLljkRC
ePiRH4Pon9fBlUzfTlfurBD1CF+IERJ/htrCu6r8gYnQtCmyLJObKYaMvmCibkDW
KPmFDFNzBteWvyEelciB0WGwWAskgNdyFRABPtS04ANxwMSX6Z2UHta514RnUprv
Z7TsJQMeEXc0nYFL6VipqykQsK8KGcqKFVSsfcpXBPyXlcnlVNmggq/7NnqhxlOf
iehbdNhDFk4PJud8RTmqy8eLZTzxLXFGxrTdSq3fEz3ussVWfFER6HmX5QDttMMz
ocqF6f7F0Ri+OX2XcfWzwg/QrwedHQw49c7VFAKf1Ct6VG6tStFQhnt9ZZHBGx/R
X14VW4N7ZgeWAVt4pkMaCK+6j2MxZpfMWutQ9KRXNXMiyqVmU6UWk9xkLGfgxxDZ
7T2NGxpo49zSZi0zGEkjjWqwSKeHsFFmICR2VNqspzYxQ5gi6SSRSp565An65q3t
Ql/A8/emNwo7tV6tgA0C9DJ8TwveOL3ieEPP7t0ydk4klVpglUsGw/DYflLs7BhF
U98OZaIHdf+XaUkH16yZEwbG4gO+v1XBOlSleNYhu2NveC1T19FRX8+2AcYMKRPX
Gm9ueUiYL8TlVvtYCP/JnoLYZwd6kHAVA6oFfjxqmsoot9Nc9vOGvscyQJ7Lq4Lk
MORrPjjYjx2liA3ykqP1NsoQ3vdaWdC3baY5+mE4OeeDk/zjRFwhrS8aYknTUgeu
icFRT/Zn0XWtYV5UAH2BmzujVrXtDTMk9dKh7rDYmQ/O8RAxzmaAnXZtiIibyfF6
RgU6ye3yL/iQSDp3IvaY/XKFFLUHr8nY/Wc7aRH/vA+UBgoSq5PGX9+RkPbI6zh8
ODjzOwY5F1rk9PvLtHGUXlhZKShg844z//BOeuszxft97/jjP9v9uQoNK/wDTPSK
a6dVbcGP7n5SIY+N/mm3ed2NIoYNTQPvlUuOxJzl49I4mqxb93wece+eVCNb/ELX
rhQER8SCxO1TNtHe5Z/XkHc4tcmRElQpp30+T0V3cvKIP1l35Oexl8aVg59KjsJD
+IiormktTniPy9DfmJN/6gIHr3Kq/70ZMlKwYfAPzfgXUXAkvW01bMhrwocfb4sR
r9YsReGUIZ77atVTR/ztYosqMXRGCdp2AbtwWHyaJkKmMZieUAvd55om4PPIEqK6
+1D7zgR0wCJaTejdUFd0VkHcpER+Ttva1vm87hNUHHHxu0OV1cfCfJbhDGhzMIe3
XzcxFJnFhYiyc1LO/o42jaxxbcbxpBKzTpwlgcEDXGt9PBPpcHxDsj8jn451xoum
mYZL+ydUhu/tCaRaj4swSbFHPWYzAJR7P1kUNesTIo/OSwZFI2OV4fru1gbHoYvs
rXl2pl8m8goDEIPwclHXykCCs6KOm3369vscHM6cHC94KvfAOTAOIJktQOEoy24H
Zac8X4qxQz3ziGJARNhRNKIDECl2BtpI11qZ1YvAbGrdJQkQ5OA35EmvrsrM9z2t
uCe7JElyVmVGtbigdROPGPFUmPO83b36cIB14Sl59C+U4MyPKpw7ZVRaM3r+K4U4
yD8QjvttGYD+Vtlx3YZDAaikFF/ojUUZsOmvAxE4ADZoJ3iz0iWi5FJKUhgR8gVI
4cyJr9SbTn9M2FEaPT5vmH1WvZuTr40j8f9MBF+e9Crt/kNgYRsE9l4iT+xmsTYr
kfDyAbTT/y/7iBvRF0tMyIis5kqXypUKWGf2zzd2be1h6ZMYNQ/CY/ZhAS0vzw9/
/GhHFdR3SIqj5CQzZrcCVI4QZBcVO+WwC95pjMm4xidZKD80EI6N2FCi/58P6AO4
rJI0GRBrkcT+wJDH8C0oWHfgjuIYg/OwSW+KGdNBKaPPxRioxedk4LAA3PJYuUjV
hbltgsqF8MsNnfDCzCKdmLaFxXFugmpEV501FXIihGZzJNqLfY5jiH07AEU0g2nc
uxWM1S1rTYCph+nc4AlqXPwZeZZuVBHrWHVhVTKr8Zk+AflE1wfu85lSE6u+S+AJ
BM23MdWpbWiUrcFrRuyYEFTtJgdSJZgxvKr/zKfKJqoXl5rQWapjkl3PvYvEcEOR
bCqqKCaHNjK3Ajr7sCAZ2MxnMPQL/paoq7qzkswm0KAa2pbV1vzkdmjGnjzFSEIn
SOSOOOySGKcmZv8bNOfnb41OQBTnn4ARJyor91IhGU9FxCLqxrn0qYTUzYy9kh/Q
XBb+BWnGupQMyeq+IqKaZZ7J8nUrgWiHvmVyMF4t+qgqBTn2k9Fs7j+3SoRicb9Y
Vq7bI/IWpVxsUR9/9P9n1jyY7L4L0acLi3UeY1nC1n4uFHyEN60yk2if2GveoshY
mZETrPcwtw5BQ0GOVzGFrnBFIm0RGlqQkopkPSISjbWkavhgNNRSIDe9A8iI9u4e
hCtW4KKYK/9w4lwTHg3L40/hDajQIsZTEn9VdETGvdSNFCs8RknK61kcgmcitIBC
42n02y5yKYB+KaX0085ZfXA2+1j35RDBK//6bz9WJ8eT+Sy4Lq4UndONqqRBtLd1
Io3oOdbrzei9dEgmT4mEWIJPTZNl7PnxKjVscTXp96e0SfgHdmaYB549kCSdRpS1
kP8dA97vEbbxg88N4jnsnawDf5TPm3KLtbUQOQlcq2WQT/jfuGociPVf9ddQZxbk
+D0LgxmODphXaC4N3fi7HofM3h6BNb0/+4qoOKWo9zMmcWHLEFYafn2st6gJKzeM
wQ0JZijBVMPmVrCpCBqVAqCvhOk5+rYbj/vGigP98x4mbCO9+JB7ezo95KZuVOtO
4B3WFkR4bj5Fx8QAxFudsoqedC1/Rh08lPXmCHxuuycJC8oasGPuhmG29Zv94dPJ
b21dpIHbuRKXz3dwJcBkKKysayG2fVehTKrtazyiqMQzTZ6bTv3SnDqCY6f0buLL
4xFihpF5lSyHUG/prFt02A6lTYKPc6knApk9DM8kB+TAQXQMg5L9v7ppvUSvC2Cx
nQq9BWMQ2ijfv/xmkSDDsPt2chzb/aDGxiFhqGVrOA/MI6UJT3E49SogwVP+GVGp
1KRgtgrqh3PAMcLire9OvmZbj2JSD1rmBWiSUNZeAZ1395WPeoqRQunKzIj2TOyJ
1e5/i97Ttmoiag31RwmUEeag/YO+7nW9uNAmFTz8olgBnvMg4bgaI3wNcZkO0sb8
2yYAXbWpeX/IUti4bNE26jGja4h7EhLEIukOwpsXQvWwXr8XveeHak5+z4PznWM5
VxUrrgSaqfTvvLwA8TMt0wQSZ3dckOJa0IkdtdbtmxdLrpU1DD2herPmTN18U/bQ
mqPNIgk5vFpKRbPn3SGLTziZSqWQ/DZi6nmOYh5m4Sl/XXh9CIzhxdftAZeTtrqZ
Neiss1ZujhzJBUnk+Akc0XInDzdXYjWjPtVjyw3frL/tFo/r/2uJVbQOduvscfdu
PuWLgpZzyJi0kQy0wbNfvIBUSHS+xDMmp5fP9qWMRDqcf1UpxLPR0C5Egq1m7rzp
tcSNJ3atcKBsrsFWoO4Mnv/IKtmiaaTQLU1MhK5G/IK6zmgT3MrrfyUIUY+P+lvo
3qf66kgKIkyB+amCCbuGnIK3xRBUDqcP21mBjn7oTVYMwG+pOE5O0uv7WlHUam52
kTtJ7eqNVoKYkBWjN/vl9ge4iui5ShT7K29TTR9EP11UnT3D08rYFFCH1A7KndUP
uDe7p6x10I5FBBUxHxQ3xwkWt1rRUas9amosrLeKdAafxQNqtmXPllH64T/qTfhu
DTPq5fnXnGgt2R1OL1RNREitAFWp3MVvHom4NOxFwIZcxugcC9nPBLPVZ6mU+aJZ
Bu7XOp1Fsjlrg/ugrvt7qXfgqg43wsypZqoNOI6egxr6E6KOhYTfw2iSzH1JgPjK
ZBarSrUp5pgA53eqkcTPRlQP1DYsCkkuWd2GDewwfQcThU1r2ehmE9ebNBmzsXGS
PbiPrGR22R2qqwcHmWtCW9aeN/cIJDAdirUcTvj+Rn4EpR4PZskf+e8aGtgbbmmq
Tn7keUPL+r1zl/0Ku/LeG0Ycjr8k+YhdYCNYQXbLXyOLjdk/GC6jBRQbzDIkCQB/
cJE7tyrnc9+YQsGXIfMEJGzbnsh4qGllIivzOqSCN4KHlXeDxXcnAdB7M+F/Y0O4
ndtr6YR08mscPjx5IAM0F2x1UeAwI2PiOb8NE2XC8BIxiZLO48Q4UT33EQ2Kxs+H
dkzuKyyPPPDMC+P1sKN266QCW1M3nEqpyR/hBfAJZcqtM9ZeKpatW0Z66TalBo3L
TT2KihyJpzKoh3OZX9fY3lFuvASG02CLxyD1e+G6yBAcnIlQ7qcyJoy7gl0V/t7i
tnzOdywzMADFTsvDE2d4ZExtxkQld+0HgIZHm1iKa45coJKwi4ZVYhxBqKOrD2mM
2DjNp9LmnwP6qWPWBczdcR1y8MXb11iPwKh2C24rhp8xOz5osqIUymDYDONL/qTR
dTYIAFhUBf8dV8oschvd2PgCeIjvc5jQpXe6fXtgGHLMVGEF7InE/4LTFR9816O+
ct7pP9KR/JdulgtFc/dQhVJrd3uP49qGymwOd7llSTS0O0GnWiuCnorBJAbaUhnA
MAkNc9ydYBZ/IlbtYbeOmyUTv/aCOcK7rLm+pwVcuHs/ODbtYQ8C3OXEMxM64oVc
kK6kW+WWw1TC2WpglNJV/0g+/bD+gpjilCqfCSQclFOP5arDyB4g6ptVwXqqeJba
bzwwyroHb812EaKwu2FLcraRXPup8pElobpF0rEALOjr0DBIlNsNtMfhnaJk/9zD
BCFzO9uaBBjjdyhE1sVN9kwT7RbXH3TjfIE3eLw0gzpOS2VTF5ewmgZQSWZJR4Ad
Mrn36xN3ye/hBCfVrNVP8LBHLGUACQxXYjU/5NcBBEx1bPFkECwLCWT8rOdwvCTm
rOjOhktCd4yjkhOPcwKK+s1peRyh4wIHYATy4crzz3vAZdnIlh3lW/gHRQq+V1TO
Mv4tuEYmBvyfaiGes0kAszuPH61iyyI603JeS0NU/mIj30BLiIxaTpELVqCUuFi0
gn5dvgcIOJv2Ht30m+pNRv+OecLj9RnQeaL3jsK9k7dmfPYEj9PdYEa4GUvWYRc6
GJT0sE6/nYBcUmKqbW4dCE0Qt21iuu/H187X7zBZmIEEKRvYwt9GyGZlJbXqU1FU
eQb5nj+Oivs/WcFXy8ygkttOHNoL6HYUz4XtXEukyhY7m0QDLtFZRxhQ72RvZvRB
SrYr9zh+DaKSG4G8NMSgtIkrJvgWpHcjElWlQ+oVyxgCcsXFymgJX3KKhTOWrwpB
zMvOjabEkPEpT/hQaeeXywoNVzpWqVjciGK0tn7gXl6k4tDr9ak6QhXs8aGrmaGz
H3apUkEKvSRmKu8DZV+vuZDbT4D0k2AKilJynEf5X0t7lsfOX8/bYO6k5yrkid0S
06WHsIUZNzLiakP+SCxKcsVa4nA1epwFmKb1s8jisGH7AJUl59Dyl7p46QaByuOj
IUyTOJVWGg7FcvF3VBEWaekPtM191ZsA8x4ia2JlW5/uHNPajs7vFECCQy1cMVnU
pY7oy0NSJ4E3aDglAyuHeZ1soRNImc9NjdNyksvJyEDONRyia6DThCBYp2wCeSMT
szu7xRj7/k3qlWGsWQaFoI/BStuap0xC5lihe89JPnMrvHDXNoU/UXTL0idzjr48
b35W/OuLbt2uk/Oyxj3qK76YPGGjvgQzfHOBc8COzMRz3lm+7fKid9gPMJQF/J+h
X4ceNvby4sW5d+UnIhvK1Djh4BMKMyKCO9DY+fcQpOhcrr8smZZOWwt9oALY4HA2
kkrpdcwA1yB0uxKvjD7uUcrgZ2gSlJtIADIjq6g0zQru8CCru2hfy3/BHMZukC9h
aMgDC3AzrEC9VZ3dXhrTsZGep0hZhM6TZc5L719fVL7mukp56U4YVPhsDCoMQejI
wyAtmDmbA/1eE0h0Nmi7uNuKKSFkAyBw9Sf4ns7hVYA7/XADhN20TCkMs+1EL1bx
rgWdMKVnWGZTseEJ+tF8rvx+Jw5QCGrVYTbRs5Kdk+CzjBJv1LWIjNfa+/KkQspc
HejiSF8ZcNkFtxo5NPGZ8edvFvF71kAT12mhwyYzJau1Hkty1ZXf5ahG3evU53cw
/2jR8PRUCkpHLl4+X+h+qqeELxmIcxOH64hdH50z5fhABk9yts9PFtaWTv/dq75d
l/o7+GiXh2B01qPslaZ1tifsXCNyH+JIfqwqGRIEDnc7qYG4i8YgJ3waLSMXAIOK
9PxywrgjLnaVbrJi6MMdGNqZ3c2CTNmmHtgYWCWWdk1SYoUyoBYy07U/zObSwOyY
BYnW7fonJNsYuVGc4SCiHBqkqei8w/XKh5bExQv1GGJ7DKivW99ZM6tpTrqBGhRD
az4KbxtcgbWBRhw3EXZ3mVw5YBcM79rOCdfJhKlmbMItYavKGzwPjpaqTILl5dNt
PFwaulAsVvBJ68/9XAT8VhPCTstwVgwMXEwgIEw9inH3RreirtlZ3giMQbGdeCE+
NAZ09qJYCRA8I9ZBuJ0tjPwV8KmK0tX0FSwYOqQjP3lLvwUT26JhLWUDGHtOAm/S
RdHYICKaVYbFUmWEH4Y1LJEqeixSoq4HQa/E0ZYZ2uUYZEpR0wRkU0k9RjJPo8WX
0TECrhuQlDFfxDrH47QspAs7ofFnwfZ5DkLT9SD/gdpWfPq5O5UTDomza4Oi9Vfl
0Qn8M52X7DHXT1NlnNrt/+9qV2oZQc3TG6I4Qh8RleFyqriK55FSZgwjMn0TMOdb
hPjLg5mQ9BlrsVRl0Ut9a1Es+JXzqvbqIVhXK3uksQIk7821nWfJPsfI8P+yg885
9ENoYQS1ESZ6nGh/Rtv1cJBroTuP8f+weRioJBMcXM5pbvROsiLltL44ockB6Wgp
cILr8iQ2AnhgZtFGrHZ+jlT3AntTWq50FK/glVDEhH7XqqSs98RMWInC3bAeHiha
XW2T+shS21CArATNjUY4L9BJS+n8PLrYpKF5PktDIc6hVr0+ayxzjYvsOnFkCS/z
t4rTLzlzi+H4oJdl0LeiFh8HHjN7f8u/jxStYUYYJvNc/bjJaRx2tuJEirOMJIln
m7TOXm8FC4riJ8gRMZiH2gYZOsHhyDHAKUfj20wb7SSKjFHkAh2eLxa1IXX5gvnN
zian0Kc9boeEtDb9ut7/bA4Si3oi2XLAvUk8UzGQz+SeCC6WWhYpV6288rVGwNLR
U6pKpQmIp4NW1s0O8m4YHKyISPNZPwEZTXnRkoY0HyVPKYLtt5lJSKVpNjL/+z4t
UVOuNUSqpfPtoqIizhRr4Y1GcGG+ct0Skb8tn8gT7O+jXXa+iRrC9pAxdubu3xbg
m8lEgIxAqNrbvlUINGRQi0/kP/t6pwo7oNF3ZSIGe69Pk50XRf/Wm0j7trxMxLK2
K37j0RiaPsWznm6aKDvo2rgAJv7SoqYLEWT18zwVRIFULzKbBk9Q9adp2kiVAEni
CIwok7ljkgDWd3QVjsl5KT5mBDg3OR7y5cnLrWGb4kdPPsjV+vY+tn4eBPnP3n9h
FOsT5q2cQmQQUAtvWnkqxR1hSES2nD8ghBg1fFzSuJnOBTjHBeh+sn0969NwPJ+y
bDmNg3Dzjjj3MeqEEtAwheJtcQK/R+kT4+FpcRiryo9suHLK0tFG4qgYWQXNgpoX
4TeKuoN+LD7znI+jOlq3JOOyRiZWAxFKtkUuB1KGFcD5p4AHA4OffdnR+T00dvMQ
YWBVLeXXaA/BWCCsCjFBTi8OZmrzNbBq2YHxokTFFnO8wgGVhSL8e1sxUj19bw4f
rMRWODzEHfe0TqpWFo/J14zlG1/SBeVwY49IPR34eTjGEry6JO0VdQGlu7db8SM5
W3yyKCmQQzJsKLuGFEB9zq+71HjRY0sOHPyy/AMAZu/G/I9v73jUwObdpTqsI1Oy
kCyrvzmwfhwm2YnjPBKtv1hxSi8BwRVOTqSRlUJSRWppTsLzgrtaugzH6Zzj8FZc
PeFu6pXOFoTmqXX8Px0DwZbWyx/B0C9ZprjWhM6DpOz+iLG6aKscakxsyUbwKGv1
aX+SXHik4Z5mcmN/QlBwhflJ13FJy8hwYgqv/FYOpvudEFF+0S05Cu9Gb17xy+XR
XYR3Y7gFfnxHs8Xay5cW/PIsmjKFXixyR9H7CMoyy0XXqcoQQbMF7nqik54pEBg3
JFYAqn04qk2+iHnh2/Bfa+Ty/5YK0Z/Q5Ljq1R8d2qf9YsfBxCBMjiNHWEALOz5n
OoD4Hkbl5m1u8P9E7qqEwJISUJ4uHC2pqy3CplumixUfANMEVsg6KnPmLLxSeP+O
YehGYE2UK08g1mn2cHdDQC0s8nMb5SPvHpygz/+l8bK1n0TtXFjW2rLrVlrBLJg8
vZPd8PT4J4+ogYabZHpRKT2OFx2o4WkvaVeyLL2nvMKGLFZdC9jR93oY+9gPxsw+
Q9eaMJ40NMyl4JAxkeeRJaRIPXDFjGPIDvPKeVBvEJdgW61kxPpwHPrhIu2rINMA
PlugZ1eI6C60kWAvP5L1iHNGlnVA0tM5y70wL2HtsBgaCr/kifmfpU/Zavik8kYM
bDyUL8JGbOws0DwfJis1Ck1wKIH+kFmhkJSBSK1eMsAz19JDsvsvtBF+vhAtJrhl
Cj9KiQ/CC2UBoh/iXDzA0tr8ACgnHKTAQaxpSMOEcTgeC5ONLhcBHrxYZje01xAM
sj5ags+p5u0hyuCNYAeGb7260DwcQixt4SWAmF1eY5t0Wz9YdjkF6tWrSZ+wtrs1
xAhLlyDG68i0zHszEXQ7dgPohXruISNBMyPdoVUuD5KfD2/XdoINrn7I80+CEeWs
bePZMsL4RpvFwSIbf8LBGUpSEItAIWQeYU0tQ5SOr+ZifwpE0oYi7ZGXpeNE0c+6
b64kD8juhc8b23e8ojeseESYbfpwL4xp2+BqrIobep7AkxtlOo2Q/flop/v5Y2TI
0lcG/L7U2kARCFJGcHFWppkiKb+jzm675sX627hXH0EmQKX0qhnMTsxWrNdfXc7S
YOkr8MiTJLWDmL9dcY+VU9xZrdpsM0iMXBslWlq001ISaljDub2gauXMJufj6L5X
Eb4+7M1fctx2ouTVNQcTVvNjXlhULuWbBf/sHlQXoFOBTQq2HKg8ajDg6d4ctI2B
Rj0uEmf8idmb96wM+7kdJnjfoJLyKCwGCh7y+LdKoDf6gpKmE5fZPXC9z86JjwUB
BYyRfsMidyvUY3efeRS+/WG9bd21Aoxlrmbfyb4YtHfMn7By0hYPg5fXiw4RgKEI
+pL/RbqM2UAnc3sdl+dNy3zaMiQdUSXx7zfB8EerqS5Hvtlrn5sB75rTxDkNvO+U
06Ox8fQRb2Ib0Yx6l86Yq8kS02/CWHa3/tzJ3RiQQo8LmNOQIDDv0UvfpdCuSM43
3zws9W5L0tTvkCIj5e+NU0Bs62K9W6Ec+2JKP6Cyl2qBNs08J0DNHWkYFcAyj2Q/
70Rakojv12w62Loii+xbqtUWSomxpiJLJEcqKmW+75ZjuFd+L5vxmNo+w9sRMaP7
wQ+FV3knaGVcW5y4IVC2KiaQ4Bg8/QsvSC0Ie/OLjI6GZpZBHyqJOrJf0AdgRgIt
Ij4VlKuSTshIAwJd5eTAwCzgoqutaizK3fzqZtjgSxqcuK7I7PTNYonqlSlh4v2K
YG7QqnkTJQD01bB+jQdRGzOEnsLB3PjYiLmPNerNRlTCwnl+bLwL/SfWjsAqP7aA
YrQ2CVtg5CMOu67UOpKthLDwVYKLD9bT+tcaMHEK9UJKAD/MX7n0oAVFagyL0Q5W
0G1KhPe5I5TaM0tmu4wDgiiAK3YZOgoR+onjFWUVa9HrzFUs4G1mGlbY6DNhk1RX
4UkN/XMh+nhq0uQ9wJOlCSXsmDt8Y7AA5G7E/u9LjKbkRodToXvFTJ6kLSCklHV7
hQ3A8psB5Rn752NcfusOzdDUVvOB1Mclmthaf1LG3OdS/kCWE5ZhfpFtxx0k2sX8
isoELwCk9mmQLD/Xzl7U7DErRxd2HXwK305NVDu8QOJGxwEMOtbY/icCGGjGWVmI
cJiRzfb0jFp4IJBc31K0yeISAGleit72adDemRyJdYcIS6viaDpR8gLAsOzDdkaN
wY8BYHBFkhU4YkIaNTEPJpO2L9dEbB0u3p7Yqhuhyaxnm46Y9fVhIIVLz9VgeHeG
cZdyYl4RRXd8dE+lVqTT9lYW92GlftBdU3lBe14TKFeP4pLc+fi2/2zChw/aqQXP
hRFhCPSnurxTdPv9k+5DR37xEsU3KBnYvFgfitDlcmupIEOn2W6G4/iQITS2QPX5
7wn64eGqe4NECyV22LF+rNs/TCRZVI1y8KPBZ7jHx2hnZfiI/TQ2snHJLI9snUpJ
SLFh/DpBfkjG7vtSbThP6QMERB5egUyHf0s3wZuibP2jgz6tyoyQFukq6bEiAbqe
6ErYB/FhFhN93uHAptH5odepSPBMuT6M/QaBZQJ1Jhvu3MlYTrysh+scliwjQCfa
/UjKQl3VBYPXzp94jSkJCJ7DakM3oe+jNoDvE/fGOXEb5g5OA799AY3k5zspyofR
rsG7iEnAgHpns5rGuj2V0u3C/8ZgsbngntpnjkHR5fq13NLnjUCi/yxVY9us/tBK
QEtDuZJFb5UXFUv1cy9Mvp0uw3RbBbBaGrROKlm1rgOwi6xANkrZcKj8/kzQ1fKW
Sv8MoaszqIW6ucJXaT24a19ChEBqBYnNKoAk4lWyagA+kc0dnfsNZfYby6Egl9Ld
CgIOhC0Z1R7dsQbIUdP6dQVeDnboyBXvIxwXLEtcciB69vLCAnzm5FMePf6VqeNp
aWmACQxntl8hDvctwnfFMFO+siZKEzzPmr1Jxfy/eePzwxNIyW+Ok1hLigQJnk6D
Fjb/aRzSAE5DwZaJsStsQklRkg2LSB9rvCw/Ddl28mm4ye8K97tsnvyj4uZ29WS+
LogjEBe8FJiAvM1BUphMRiO/AIoqC3M2lif2DxDfNciJ7v7SXFqiyXVwycOB4B27
fMrT3Y/tap9TlWfUl0cnd6oZpGPCXIgYH+gpAI7RMjJVKv8x+HkxvqaAB+91Uw9R
Kl6Q7F6YWGpl8Y8snrW/tjrQZvmIQVze5JnUDjSCbIHMSlmMOpt2lF3zprNRff4k
qpNyQJjiyDuHVG6mmjVz5mpmyIsE6kzPlbuLQmrIJ7TknqTzjwM6oD0SFn0/aIs1
7+GWKRxRtjVNBmyHbR18aDqzPdU8idQ2QYMOuEabBQIm87uAoaeB9BJU1S1Iiqjm
9O5PZQq0mu7JDsWVnJHnvdDbxtcyVT4KZERM4g7nYZND7WCZozI0LretX08HLhwe
mg4nYmEcAlidv3/qb/K+EZqnJ5tffE3TRMDUBqzL5DpUqC3pkJCqoxBvDjHME+8i
NE66yFUzmpmLao2BWQhKVKAmLRszfYQK8dJz/XoRrjazKhIGzt+zrtUoYSlYYgAj
wsxqggi7RnQ1h5+Ws6H46zdmbZ3fNW6hS9jXhC5Hv6UUB5jwNFlWMd6EiH8BLbYv
O5YsJH+ft4s60jm4D+UsGqVB2LWbuft/G8ivoy+0EbjaMxXalgKcUzXl2LVBTuhi
l2lIi+rZ330gIgdQv8OpoXDZDszXvbyuk9fbMzCCLDLNJZwObdlpC9M7YZzHRcBF
HEH12Secq+j085/wgAoEia0aChiv7BY/t9kuD1lmGjIztiCGd6+j6zTiRyOGBPYJ
J5ninIG9ammDobzqn4bdrxb5W9UvKK19ECPZLXwJDQjM7VJHrNDeczm33u1qkDLq
is5fZ02Z2fTldcgl5BzthMTOU0FCakpkp9NbU+dSM6dRQVO1YjeoyRSoXLKrQ+pF
oLN1tMwprXVyuVI0bPJeEWE9ondRZ7pYC1T3O494e0PFLOM72N/8QXJHHmfY6wVS
yBYuFreONMVHqedaa9qk+zwIYFxH786z0SWZwYwimPL0eKggqsMU0EDjQg6TlIx/
obEOxyOOwjPgqCHA2M2zALK7G2TgLR5+G9TbusjXyAlfCR1GVnsfcWoTJBXuRhmi
Ypd4WGqtxKU73VBmDim41LW9/oQy5FnKZ/MDq3fs5jsL+doNgm2ES0UzO5ITcsDx
M353Hn89yHtUtKypOhqGitGxUgnFTzhyKllBRw29gKMfuy2xPm5l0XG16U7uvZf2
IDX6je3gm/AjSagL6XQVJq5FcpDGj9+2oiUW+1CQoCpA0wQTvK+OJ8iCtH4GuRze
w8Z/aKBXTKpUwe2ln2Mr6LIRzfNA1N05sk7fchr9wwcD4TpefhGcS5FOAKT0ZjIL
Jc4FiVwqOTxn91b9Rmp9DuXyRylHgtsEG+1CuOQeMd+OWQdrqL5I6OnioNTK9bke
rO4yP0lUhlJW0+e0PWeasAoUjUN0WOYTJsN8YXZor1KMm5sFrQcNaAPE1gvKCvAc
y2UbHBVcMLFmTezgdys66xnRIKLnA5FwjGIIViCvW06bJA2pvQ85PN4KcINmLdkZ
2+mzw7vHT3hmphZPsPo2w+81hFZG2sukNnxcHwY2WgHWP+0ZnK+tA3kGeuehj22C
MtJv0Nv07u5ra3Ld29wwVhvsMy/NDUn18e9FiZYlHQJgkTcz03qiMMV7E55nJ+Xb
FwOo5QOfmVFHMbCqN24Gbpud0FunxigsSMDVHrdCKUcvpMswZz9HfCsj5wl/+dCj
yQLkkpnGOIpc7he7/OmiEKGq2Y0FU7R5R9Ht1I0khJTQFZKjz27ZCcY4tExmRe5h
SQUWlm47LXwGJ4+cAyhBo5bc8HkWA3VcAkkyeRh/W3nUEpKcQKpwJXPbw+tsbGZh
YMFS8BHkoskxOrRpOz3qipLsoEg2MyJ4sPspoR0hv5JkasMhCJI2UegXDm0Rm1ez
Hz1rE2cq/KbZP3lyTNzEzcbcbryPfH/m0fL2GdYrcbJOxhbmQfgNji0pStmAnZVC
7ECxOHOXpLoo9MIOzz4lI/l2YwSRxNvgKjdnkKxZ+wBkinkF5Jg7odD9ohCR4ryI
Hdtii6bcj2wN0fEBmiSwxUrbooP/tbB5SF3h2bTmA/LchWY0guLwPBlm4Y7EmsOv
PeISpjUcAYAvSL0s7tdzklu+N1SakJI7/f77v1QR/dkIFCj+Ki8z/76kj0HPzr55
vATNLYErxuhkee/3hnN1GpsrO7KnArLdPPU5zKd2HXvd/9l4KnLowAfdA+C2UBfk
rMPDEOkHRqYWn/mBZOP1hJgoxzZcjbm+PozzkVzLGwGK9lc/RVCkuF8cwPPG2b/L
DZU9o1oBfJjh+WB2bwUPNoJqUi2emQMp3lNlGK9Zz4MQ8Xmv3NZs0127Fz7XDpiw
xZWAr06WENzAF5ZyPXpNVkbaUrh5DfZquPlYoxE/5pP0/4LhGrdRApOxKxMECihb
gyCzanYwvU7vGTyPzGlrSyeXevQ8+Hp0eB8hGyHFA5vECI0K4pozsmEx8iEzHmH9
McUkmWSKe9T7bwN5LVwuazvEpzjZOGePgNj9/Hf2G2Iw31nazIf0b5IymdbpXgDG
f1DxQZW8OF6CJce7xYbFktMMUy72yxNrEvHfeicnMzWrbHKGgWfwb1lYAM4rWW4U
sEA4v54NBVGTANBbEEBgiLF2KG3zqGupPOb3h5UbWS+5+yDbYMxrnEzmEBanRV1D
lCfyo0sJSUTZ8N+sHTnxQwy79QTbPnVf1MXIqztZpGcMjaThq+GxPIYvyVEwiKd2
yJ3HMMgOSK/i2PHMyfCreXRTYlRLwqkJvD5p1vE0B9rssHgkXwX7RWiben0trf2s
WXb/mjjusOR0Uo4lBKOf2eFVo5IxseffNc1p3VeYe86itgPZ3MauETFnDA6m9zcO
o5iU5wZObozh6gZuDIsOyETr6hM0JgYl8kKSvB/ysrApF7e388WOTVjWZz3GDPzb
qGCtplzvYOQIneUwHQYVcM33KprnqxF2PnmrDz5cTeJtM6PDgp1R1xNbqRq7e9aS
xPV8f+oZXzv18KAGJp2Idu006Kw8b+SOF7fM6/4FTwvieKmalhot6vttob3VOg83
9K4NZgGEnDapLj1VA44IoROLA873I0KNk2odOybumPj0Pj/N1K6g9nHqGA7Bipqp
QbqdE7tZh5nO0+9U2NzHSFIwxx2qdJJ3jQBcKf/V5e3Ol6HNR3cQZ5ZucmCxd6MU
/egK8yEiQIRlyifkVV821b+q5zT+cOdEdC2KY78IK5EQFgjDlqGMxhjYh3C+Xos0
a8KOeow9dh4K5LsMjSM50OyGcr49HIr1BpaYiX4ueqpZFvGszRTh0n3n9x5cU9j5
BFg6MtKp/ftTh5JDuhO460sX/ZDMwdAkFOLcH5XE+t0aS+K7q9ZM6cmMYMgM5SDn
XflNQGXrZGroocChINxGV2Vgux5kkMwtauEhl7eNC3XpoSs4c6sTxaNK7QZe/1bz
g1F/ig4+rLuOCcjoQhXaD6mpxhCZkx9EjetlzswIQMOt1JQpJQoVyfbxNnbyn8GH
1xVOa4eDQOvDPLD+zYn+3kgNLDO3yYntp595JceSGH3WDc6Se5a/aaXQCX2K+yCv
LdcDpxCWM110EE/ObkX5xiIxCW3cnrIEDL/ptiA4Eu6h9xr4LQ6DW6WVwoehfN8s
nKGrH4Z0Lucwx6c3zH/BrESOqAm0wF0vYek2AA6ebOEHtC+293npT/0nNvzYgyfu
IUBddj7M2gyjX2zjcelO80tjW6k1Jvdi3Cq/8H9mxz+ifPw4tlcjV4slDCkS5mcG
YINTCx0Sa1gxI7WblmmrzChpR2IcLJ7HGt3tWpS22xAtcmXMfONI/2Ngb3v/KBvd
cdD7VLWps8dVTMAc5ttddgdskueOW8Xjjq3CC4iUDrgiyUm/xQABxm9xIXci66Jt
jXCK/Shww457ptbaJnLLzvZQvsWSVxR0qbS7U3rYlnJAMt9tIoMUmXFjMNX/BWSq
clZ5dRzLO+enx1s1ac4b8S1vvuMdvXlmMNLLg33xeX6wU+eG0gHsGvqcZ8Mese+w
1tV2e8AqP+tudQ00ShgroTmFX7SpYlXRyZOFrsPrvMTpoJQ9c9Ud7B4L2DmvwetW
lgaVOZM6l2XrPP+/JftYt7k6QqGK3TegrUIgxatH2N5Ivqm9ZvghVe5Bb6X9YrJ2
pZsGZUZrxj4cpaD8OtkFFZBf8BM8iR/eToQ505i5ua6ExWN51Dd9AMP2Mb/nx8+Y
hLV3AT+JXc6q9An7kFsDKxYmRm3SgavrvQl/iViw+Ke8WhGzegYmIWkANF51yxoj
UKCWQ/jv1b5vcZrCWu5O+MWGAm7K077bPC5iKhd/yMO6FidOKXI0cZlb5DEuOY1A
k4UhIzGegMIHFL/sHrzHtqFR/vuJpBI8bQb5BkTbbSIK/IBLod43OclFuy1Go/VS
XYw+KEun/QjxCiS8zyEcqfT1jeXDdD2/rOi3DQDt6sVNaEPtpyrLufwTL5P//DNc
ACzdMqBJWTDYn586nfpKT5R7zucc3mLzsheGAMQ1UqrtAiXhxzSoFVxaaoFXq+59
LddIW1wDdWdfo7Xs/ZndutkI+mMBLeM9JN1h3bsAsFiHWhdrn8NPQyblsTF2qTlp
/gpNMCZ/pzKRPEO0uN8OE0eYLzWyTcOVFZ3dNJUWf0cHyz9eWcpMD86vM1vciw8A
OO3Hon7ZgoTEEL7fcuxUwwvlb4INBlEPmVLDLpbA7qyQb2EV3isHF3KJ1idAxx80
Q9o6wFVBduWFUVTWzsiPRHZ5HMefxDArYYJ6/bXM39mNBMpyrAUQHiXUy6n+//GP
G0zpbaF1BSc5f6TwVy6wiRabSU+raCP+nSBlKJtsKJctm+QyXL55ZTgXBMTURbFk
LB0xuHHXjY/ezpQd7UMizU/iU94gH7naTD9+RSOAfjbi3g4FsfdKI8kEpALxpZGQ
r6tT8czzLeH0WIVGUWkoheKKHJPp1F1GQ8wsN9K533k1lhej5g5SlBRwOXrX10+g
5hQ+tGb426y7rdPJLfwfV6dflMwSs8ohOMpMsIM5/DVTzIONpOSYZhmbQM+3rq0s
gHTcDmRw0Z5I70iY6XqsNPrjy49d2MOxYRekWDbExLnTp+2fp+txoQusGx1ic6ax
oEc4RLZIZ0YgwG14nuF3mQ6EyEojz8HNikJgABQ5vag9fJbzClKrxx8EoRXHN0XQ
rR6/T8dgY/2MZcFfZ7YobkGj1B2yaea0G3h3nylfjD/IqaHdWhOqqMl5tBgQkrZA
cDlTU+WuaZnRMPziC/1LPx0f/gtyJiT+QQ+KAyHBgO6swqmS9m+xu3Z/GcctUFqO
Q+wFPpfnWAgEPM+n1eCPL77Kh4vQJYk2f/W/7cEI2zvm3tPAp4HaloKgFJ8g20VK
uK+MoO1jy3WUvPwbnyNNUXDwRbO7RhHAYYEcmZq/eUgXNt8Nx0H6l2KViP0OozS0
AVpZqb+RfdMoVKQj6Qh5sYoh4t0efP9juS/IMg5d6++rd6EJtTV0TACrTlhkDbVt
wDDbtvZcMIM5JjDJhp6+C/GD2wMV0HH0bDBzbRyukS0oLukrEPaVSiqD6eK0C0fa
15fVmsZAfkcJRuYhpsG7ZVYCdfonG4Lik1aLjoiJvmKf+/i3G/zjOClgLRvCPWEa
+vE2xbckTYB6Ix+c45GK3qFYLoy6FCHQTmWOOmC6zbwHvpdFgmSpV/Gj5hxzyubv
DhnVWHv+pQc31udX7oNbO8vHzjwAseOvghH8tYPA5wQmxsDTeK3BbzupJcAC4Pkq
TCTZtdKIF/dRlC1MnIDdvhKV8XtAYkJJGcDiyhrB6HFqvUoLyRKDE8/lt4TXFNmN
7fI+aQQ/Cz2XQ0LdYQkRI4iXtNIFD6C0bdsYShpSg/49NCp06qvl1dWsBtDh3y4L
x4thW8Pdt9HTaGypcbAeX6TdxTBLmFMaugbt8UjSs2p1EtyVSQqEVs/BZeXbMoq1
ZEg3A1EsHfRx7FiBCCj3fjStOJo5uMoey3SZHVaZSSNzT6WMkp6hxIpKfy6pDXnO
QdTc33FzUQHcbX1F1IQF1YVh0pPZiNmDwjbIoBFUtS4L8xvUUsR/W8pqC0AinKWY
FNefm8ECAeu7tS6zXZYtuMFzr6M9fG8OVfDRJhIV6h2/ab3DycTcDAu3BERKCGoe
Wz1DUQrf75cjZ4dQ9Es09JZdxt/zxOzQNIJs7XxajO5oRbkYXt7UFD3rs+6ZR62K
Pm9ry9uxJvZPoWlLfmZNdjUxrIGGREsI4+bqaLy9Z4UQBZZB9zrD30DlS58Fe7Pn
W0CDr44iJW/66VPLAJnPd3atBOSfPwCjSfnCM6ier6mOUs0ztWfLAGR+QLOGTpZ+
hHk6m9AK6KWTwlWjN+owhLQbEyOhaKyCUpb7AcZff2D3ow/AKHWkdES023DdeJBN
apcZZevuGn/UAktZ1mZwN09ndh8DrmDcHL/V5Ep1ys8f71DZoRVqC7UgybIMxy+R
rzwrdNXcdNUb9n6pp1S9UdR4uWdVMKqVALJdzi3122fvGFtrUuVFd5r50Gzm1RT4
fnRC78yQdU+wqpAb6BJpBs2uWLEkwjohC9kOi1LvAXQKTjftleUSFm342LmeAiIh
6/hQ6RkVcebFPbwhI7/hn/5BUL5RFqNH5MPPkZ2Xf+5i91UAYYN5KpJtaGSrhU4m
XmA2IBYqimRvyPhi/P1c2NviqMMdG9Qq6Xy8O1NpY0xKl98zijm2ARpGVrIoGOxl
1O8dKSmxGYw/Z+ilEB9HwUafF3j7wDfAEsjqRIV6rWqaEUx9qrfQRPuc5IGC39vI
0csPRchRqtEYGwJeBhwGZ6iCbAd4nNRLoL6tZMiwerK2POdZwS+/FVPaizDxw2ut
0l3qL8l9ek4vfbkat8QTblPhC0TiYvw3R9D7U5gUadnlunRyyClxG4+2S4LRtcBY
2rn4N0Xy/d30g13HEptkys47GDTEsYvVK4MH1e9uFZkyTSCpMf2n8bbFo3hOL0iW
ebrCc8RdMokz8Yptrz0TPqJW1SuNuvPxfKdCPYK24Ujw0jSs3UsG3W43bT1j7gBT
SW+b+pecHGWwl26g/f19PRMBWP2L4nkad6tRJHf5jwNwYIwhaVs251JZkJBjoiX7
v9RfTPcc5QMkFaXsPpl8dUmtavfIUvHHg9K/Eh8F8evbAk9ThJ+/rJJZR7KJfMvO
xPjhfM/qm4wPAD5zAuMHgpS6ILH2O9QZ2HthMebDUOrsskEk74N/U+YMze85fZ6C
c59lb1GtQW8F/0ELP91UMRpN6AoEceSO4vHYMPEXw+EnzfJZi/ifzu5I/7Kblmji
JE8vwsySWCykj0fm7JxOzOam9WzTDqKaqN4Q88Ok7OFT7t8bm2icnSou2wTX5Fp4
hpoF830n1uoI1erauUx/Dps3DRgzzRJWGfTsj5AlYKUICJ63QxymMXMM+teBkQM7
1NihfK+ob6zHT59lfiRPbWIufz91SGKdt8ceXtyv0DA8YVVAtGOvz/kP/qvO8PEO
SgwZANHWeVfzgmSfAmmiCUcZAMwNl3Q4wdkWlUpPASZkjFcRdMlnbLZtLxJX2iR4
dyMkauXzVOuqgblXyHoJyeeF5D+iCtJ0/YKpu13+Nv7yMEDYOj9XLukFK9FRqFBJ
epVvAQr3vnKdEM+/iWb+3D+Qc9Rj+hgv3/1BmmVvHx7vpNFk68WDOe1Uj5fBtlwZ
gPpKdF3eim8BHQdWdflICPscmD4odGLXflnWztpdtpVtrxKWDSf7hzzuva/FpC/S
pCwi4JQXU2ucH1wQkzZKjIfb1ZitU4cT5wHOEcO5f/bVKlIcc4s6CdCndBCBFtIz
+Xc3v4uHHM8D/4Bp5FYWIYQzOdwdjxl9hXUzhw9aAMiPek6aY2F4MRQRlx9oyAlc
vviI4aoIJLdFU7ITOaHRWuI5o8HyYzBSzJ00NgR4r4PRNaheT5LbVscrEhHlTFnA
G1ZjBqYCI15Qh7UM0eRKgReuwPGmXRfs5ztxFg1GyTKq4XXfAQox1tOOzAuW1LBB
Hlf9I7b4qnh0yxyjrNAaNeq+SI5O+rZEkTRRwP+uyiYh1hqFMkNfKTzUIRPBUmNJ
79EIE42Hx5BC3WcBHPRxYIZA1DHCAOVXjHY8tLBe1l081QOgFMhiXArJDsLyRZDe
sj2qgSZBYCodOI4eCasqEMIN9SrdJf+qlkCexpwaIz4E+l/Cy9c9aga1NSV5UPEF
2V4tNkmbYjRRU45O3c+xgAd80z/T6HNgG7rmGFGGAYHpiYq0vj4+xmeKpXK+HXvl
I+I+yZUHuCn/Wn8wSRYrsX1/eP4LstRMYe8C5xwb2Y5n6DlH9aIxb7bC8o+U38G8
5FsdChtXDWQttz5llR81cU3GM9yvBHvIdPtPuNIIJpBP/La7RcW+ydLMjKLvGJOo
mffjptIvjZPKOg64x+LRYdgLWbTjM0e0FtoUiOaE6ogpN+hIq59b5WCEd0Bapv5V
XryALM1NSgO6clrU+fZLFqTRnfGr6P2xcZVmY5hT0TGOVOAefj/tsgmlrwsJXWA5
PsW/3UeV+Q7BHJBEFDEWXeVE26S/POy3s1nYTgaRUzwEZ5j6dLnWojlsFVFI1r4Z
zyfTkXS5SXX37skIHt3Tr6bgUSS4NOEL7MNZhtDV1pj+meVxZA1V2DdR1euriwm0
VpPmSZALJUbSZzJPrs1rIezmDd30PD8+tBUgp6GfhVA5CxUUQFu+y/1SX/RMtq80
C7N6fI/6Cz2NN3YZfm/WUlg6WXYi3SLuacSou7X9cTCUxBCohcCcdS2U3h3bkHP5
FYY95/qkL2912GLKeF3CD1pUHaG8npLgZCQIIAZFK/1Qje4Bde3PlV8le9sxjRF5
mL6s9Y9Q7kNJpORRPjBGgQmWSvYkEMVma6xOBvwdPKw0QmGUBybosUGmY7OQYHZ1
+umPLMsO3VBnLz18GHPdbcVQroDoJFesm3OFOykJMt6/K2E047jDruI809viAk3P
0xtlbyX8D3GbKjNccfa/MZ2CcLLUIrtB/No7gbfZWTHpnoMP9/el5bHyuquNvnOO
OlwIR6daAZPvq1F0W/SmxBw+YhttUmrYeIyJ4JsjujylJ4Sjat/yuxd9/4nRU37G
+lwmShqW4h+mAcCXUqSY2CHv9G2kg+zqwGnYxFt+sclrSJxwWn77sAZOQyRoWOVG
aj6pQV9FRZ1b6fqEJyKMRonvHxcLFhmK6Zmq8NX+kRrWJ9EwBnSp/XR6Ph7Wt/TO
d+NKbgGULgk754qjNulm5csulFUTp8K4n0MqSw4RBX6T3LeyCD/jQeDQCaTOymBO
7wu74xOFwTXaf0GK1LOoCzf68+X/j1SJ5TFk9GUW35F8em6I6JjdFDJL5PpqecMf
neIb4UJySYcB94PF5//9A0FJR79DZluueWCS9aEaIC6hJwGd+VhxCaQR/NSvw6xT
UcPh3YGcEgshNqLUPRQC07T+oivgyvgx99UQzMRZGfBy1iuoeAnyG/IU7vNfa2Wd
fXfZydXYkqjQ9VdzRoUPDxSKR/cXS/jhhQDiLOIGIp6tqtrw0tAafM2Qb/ikU+my
UhCoJOypndYqNUri1oYiiXK4yVPYxZGTR131Hh4+0oH5i2bBBhT/pxCpbarrx5f1
SPK8JlRKwo1HFDBZvo8DTK6i/nCU8T+vMS1nFLYP181FTL+mGgYHstM4yGlyI9d4
Hl+YYueKM42FK6bUE9do4fA4XrnLcFgeL/fwLEhZUoO5qhvtkIpS1GphdQhs4BTt
YJvLy8cnUrDftcpQFQ5m/KbTBLTcZh2JDChZFJnu0D0q4yAFOsYAMrDVG1bRLKl3
BM25gT7vMKPSsIUpON9d1n6VrgaCOIKg1+v4AW0xctJ4GIzRDKFDPvdnbpErtibf
h9KSjm0YCj43+Q0HN9ERaMdVYf92vjFaK3cx+sZGEop1H4gNGQI+gD87DbLqfyLt
LzjjyRutShesfbr3T4hnBcfMkmiAha1F7L4tmvyIerfZYcFetcHzIUV32h5/xIjg
0GJrbprhlmI985sTT4z+ng98zK1ZJ3z8wgTZBcgwxZEenKshrFQtGwd2nlX7zpxg
EI3kS2Pm7mCIk+p4tTCINLfAxA8TMYQQDr0k+mp2YtYbUEMbG+Tso9mezWGLo8bR
HRiIu2KJaY4U+aS+1Ot9fSqo5uUqslkwSYjpV6qixbOdfiNH0O80BNUXp1Hi2kUL
HROYx5kJx/a1p5vs2vUYX2HbYv2KyXkH78nqGc+FAVOjRMNTNx3qS+L5nGCOLC3X
Re1DpL016hCkV+gHD1q4opX/KuApNnHt71Da4oXCGDncphQhIYlXE90hbvr00Qhl
xqjhtl46HLlTla9GRBJ5VFcPS+FjX+KfKH8WHMDl9ENeruGeS7ngJVrWpihHQr+Q
YUVg8Ie3FID292ApZEMzPXdUlUnF8YAhiTDK8Y5OiIhZIrBXVGeKlJ8Ic02OB5rK
1Pll638APvl6iAKuEX0Qztxa7Ix5NjS2WfW9uP9qG8vxiPRR1fuWPHJm1aMwQVZd
cwTlH/+Aotst8TZSMevBR/ws2K/dOIm/2lJmNJaocCOTPkgf8DMz3YH3jhqsf2JN
W7M7XvrhPXN7479HdBjVY2WZt/hV/M4AKk+5cn03+/9uAZn0d7zMZNW32qRHF5om
jfgSb5WeKQDN/5TWvI3Vb5InjPukhKxg22n25BqHfuAQHeQerFS86jDFi/Kl5xQO
WzRPEjP1yMCsspLW2fz6LOGl8P6iAZ0FgKIh+tIqf0pSh28NV/U7Ijiq5a3SOgwD
W2OxulasoTAZmpnPjRpljZxPcN27p3dxN4i3taUzmRlu2/dL5NnAHoyX1Alh3BR+
yOukDHW0jcjEHLqDr6kMGfKt7D4wFW6H7HUwuNsIkqkQ+MeJm2GmamuvmHBmGoEz
v/Gwc+2Po8J2y9w/ydZPubpZ0/m/A9v9x7j1F/QOjR3Advbuul5kqilO/9GDIrDT
Qu/RcwDozavQwelcqsBgEWv8jONsxuENrZtJD5CmEI3urEOLrhhYnLviNOmgphSp
6xiJSo2RAXFTu157QFfSHqqpLEPkGXAd7PvBC15jBslFPwHmDn8WDOFCZBczXk5q
cQuptUdGcvSGANGuARG5z3XCaL+rTzz+rkIazXxJV0QkuHaz/xoqgeRZeRwb2cM0
a3qh7NfCJlIQXUOU3gy51H4ft6nj4UdmTUotH4kn90rY0ZngUtBfOFJ0zs+dIcec
/mN6zoxUi2Xa5DhVNUzF3oobaqfHqbaJ74259J+sy0gGP4StXo+cLxHK8C62hSgV
U6wOXU1aF+bpUQSVisA3x3vxxlT6UhIlG0SvWiASdIERk+VTrgENUyzh46JmHKCJ
P31Xm2Pz6AEmPKOEp8JREtszaUGiaNVdKaYReWxFh3I9L+RyUrIWsi1oT24yOzA1
DIU9uJx9WyqMxJFMxN/hRIDFy9N5p1UNVgdMSzGbLXt39KymSK7WQ0r+6kPb4R1i
BxbHEs4oWGPIHiienD8Rfh4lcY71s1BmC6DPix0u2379MbKwYe4/wdXEDAhF/6nK
H26hnbHNkUzMFVGllzgpXrIIlgnymXt6JeJND7gUOJmcWMHCRisdj6NaPiukX7kQ
LCv+fJtA5mGGa8lttuW6h1jScJwg6sYwqSTVIoN+oxUoi3362q7O7BAv8D76n4wZ
P3ovjT2R+gQPVAqQg2M9e8lCQ1is54WA5ao3PIyv9act3MBzJBb/BJ15QpbROhm6
q2pas43Q0YuVlLPK5b/AxUPxm8HEIxKnmENmOw/m+g9LOmGTlFQskiqSu8ELVOCg
wXHkpBIf0IfT1ebsfEy5ISEUkqioK+SFojQDrHCfkOZk0Yfk9ZyXYnrDb6370dJ7
ZrPG99dOWefZLXrt9XfnyJ3rIwy0BV0xkMmVyLXQPNM2JWnJeNc9fLWKFnKRwibT
oK0KWbHE/2fFGtfHEvgq+piDFwW6FNbwCN2IK5yyq/eTes1/PJqGepW6M9u1rP1I
L3wm8pFSndZjy9F0Tn4mkbfVDusvCG2+b0N24kVJnZ2P8MBlp3NfrkzsfTm0WOK0
4h5du2wcleXNrtYvBp+Vjn0uAiCvY4Z6hUw6iQmIHEGDiyK8RMqBZuFmtT8AssHO
un5s/NqmCX0EoMCcBTlil5f7u4XdV2aAB464cD8EfZHC/CaU3t9jDiYiDnElHypm
DL07cObzjQqrEJBFa5pUXsPCUIKiFjTk/8WCjhchP7a3GitjpMfXGx9BqcKaGCiE
TaozdhGMiiksbylJQNT6gmpXcF4JJH40xog/m5Ufr47sI/anFHF8ee0Du/9BseCv
cjL0h6vjwzCbzGoPLLWMZyCGr91LKiOCq4IUGRbWWt1AEbH7LHBXXeaKXKqsYDJp
l/hGWM5Bi3stoON//gcNv+pTlD8PEhVIn1J1EAhtDUmuhI4auDvO6CfuBxQBWl4g
y4DrerB3ULIA4HYylFrsQOxzJgrV3oV99RgNiDrAlNKN45K5BzTceXv+Kpa6g3OE
efYbS5/MnKWvmDe6byt1DzfYnj0c5kCe72hDKZcfNuPgydFPkm9Wb0r4Zhzf7Ak7
cUQZBbeJ9lUMXIZoKHTb0dXjU5dgaeqNtEB7rCFEac98N+2PNjUROUF1XcL4oNKi
4E2M+9dg+hDAx6RBT/6S/VoSsr69NMUx2qgDSp32FgVozDKy+LfQXRdbSOyh5aBh
XEr2IRuzg1+lQqu2hmHJPBNS0YfHX0Fq6D8DcnRcxdJIQmlJyQRnoB/wDFLuZK/4
imDnjiTl+hLxlKrufiY3LrVDq1Lj2Vo+UxZQs4jRkwpzdJFcXUr+sI/kY5QSDKjT
w+2JLkYbmo9Jpt23mXnE2wODh5eyXtUtYaw3xEaMoTGizDGb+CUiGHzNhA7VFWsL
ZLD/jiky+lwuFFUJ+h64pPArL/1o54gBkeAatvekT+XtBnOkpBpPFz8fk99JbYkN
1MaCuS9Do19YsR1lldqH9EUo3weQH6zw4bhplioREGrmFX5rTsEtIX9cZOc7J+Az
A9hMZHPrzV2cBZCn+/ITdWB5+jVyWEmRLfWtTsoscHWPUaDlYqc7wkU/SodfzOj5
oaIYxExo7JqXs/F74RwRK5sCH21e8HPO0kir2a5rHhIuHN5G+FNrbBwrBsGNucUL
RdHJIdiJhlygzmM+PTHpWWgXSdIEeqk+2tt+gEDR/nNg5JBwp1nMcbY/eWwvOQsM
XNdIWzROjHHXSefnHSTb1OC8X2SKT0fb5XftmZigB1FTAHsG9CNhAKfYZeSXEBE0
WWjGI00SHQLsw4HGMldAVf9S1y9URQDN4QO9WIAcIoKpBVH6li4RbVWpKtWDn+QI
tAt4XSDHFQVVucLfFv5bq33hFGufABcE1zz5KeXQz9ILzLFHUfsPytVOOh6VJoKo
fmj7XLnsQdBYGYpoQ9d3073pEXKA4vmvWP2wHHEkdgSJf9HMJ/I3oTliUEmJECxK
wt6jKGrD4s1hEQ0fZb+6IrcFuXVk4GNgKkYVr5SBQ1oP3lWaTXn5Crtupxy1GaVl
yenOKidrv5seZgwsjlMgfydVSd5dxCIwjKpnkEg7++f7jrOcwTmXrkKuZNMS14gr
W1rlfjrdPi4og7pKZAXxf31vA5yhYIJeH+/aHx+tslGtHn92ZNJUS49X9G9B9php
9UtPBWVfr6eVQCs9ANivVz6M18UIB8z3NyGqil/qXs0lEp0X87e6bybvuhsGZN7t
N9I4mP2WBc0UX2MWtGjzu4WFzkegT+SlkWzHxUNwY1Wtr77W6EZzBPVr+h8rFk3v
HrmeYzeg/JRJSIvb+AvGivWuQP/Dg3YL2XcfSNOKA0mvW+caglf/P22vwuYMIh4/
tZypDn4aQGi+4iCzhPABCW0EGgH0Sw9jCOQCVAosmrhIL3gRDMxeCKttwdyvQYnq
RVPc4P77172U6at/ZQ6X7zkeojuZwEG8h7bu4WavuR/WghR54g+o87Wq77HtuEKV
8XJ1BVWPbGdRoZnRcKWka70gVe48KcABLDIvyMHCJYOjV0X2aUibd1sOEOYZ3v8X
H2mPPwExWbjeDdX2j/eqLF8/7Of5cqMDtoV+4lZzp45iqFL5TjEbPfGgQFIWoIgG
+QE0aLa+7ZCgG2u29XLGAoam8nDI7G5eyZQC+/rbNUEUsNrbhYVuHFnX48jBW18a
97+c7sGvWI/ZNzDk6uz0WTZ7mJLnQ2IOGrTHN0lkwElLcq2tm76a3S0AFihDYtgN
/EAyecimxxYKND8kuXZrRotPsB2xJBM472uCk4++B+FeVhrhvRsZ5bU+g4AD33nx
qzi+3PRHcC3VuN4EfMtP+JeqwAiYcZ8gmYUfec9N4cWSviTqZTOhxZivJwSEtK8f
tqHXDeRB25Plb00mSbRuo9lllNIyLu8ZbxqSKOzkyLN/6ui+nnEQwDHFeInme39q
AIeyxlbqCz4ahtf6Qg8Qqbq8b4+iC/QTb+axWAcmXWVkdpbgI4k2/D2uMNTymo3E
+j6SNegrvCc4lRyBM4OJfuedcqgGRoDCl8EyI2bYngxkc5HvcZpM+IiA2asZ+5j8
G45g9sTnYaY4KxKoYVudPJwMwU6109mkQWr4QJbJaSfK+5VFm16jsiewF15l45yr
leH6f48XVW7KyvJM5Rw5ZP+jCU3Umn8NmpV5iCAX1H7Ek11GVL6YN2a69R/EAhDy
8czC70WEuuHE16C5h2KPOz8ZVzIVWj5E9y++abAkNTXQqK0n1kzFxbAiPTmJFJ8I
Ph+p5EPGmeLtt0Q32YH4gxa4hgn80+mOfMKXeLwlZo69a485r7Z7C+5Jj1vUAhRs
nFK/cn0X4kYpEjRVnfsyzOcIJZBj1HatGKNqoQrL5pUi1oL/wWgwTtykK4NyBxeX
4hjsqFdJHq45J1Sgv0VQzivqUfWa8FjpB6kzQF95vxwEkvEni5ovzbGOaMJ8ZwA8
Rc9s14miPL9SIKWlXnwqJSJ1R+LtWdljErdwSla9UIPCP5bFNF+o2YhjJxBEOz9E
r0QCMPM/tU0242SQw/W9LYhuy6XsTkrAfmqqBA/SuzQVvimghoL64AmGebhV+qzM
/KDwxqlUMrSoXPj75EWZ3e8ItjdqLYZBRzYheh66HSY6Z4//pRsUDs0J8emITnRk
2DzuzRUn4q55LphhSuYl1IUmPUUmbAaRrblpglbi6HHJwtZACXEoMjz2dgVjBS33
iOxZ25LZihktScaUzaH5FcmV3uxzJnSn59BftwYo24FDwpHJcJg+rViYstRBOuL0
GuLURykKmt343BnGVClCcVCUHSzV9ON32L+mbyv9a7b1cmVWDXdRfT39eGVRzTox
p5ZbqRSerf4YlbBmu0Hi7Y28fRVx6jYhV5Curh7BwFOmhdsQa/qQEnhxzoJjVZJo
Z/hQeZ+yeD5tEnH323vMZrSslLYtpwuBTWRvLiB56+uJH3cPsuJ9JB+F07SWEUwl
pAaVAEGdZvJ4a9XyOeBTgPd8b7yYESMPecKwqpaeb1Vf3yD76NjTfzeeCLmvs/Gb
q/0YpBh/YQcVUmn7zjYsu+6lO8on2aSPdy85GDCb8F5XSqrKSvSyEIKxj3qCYebV
gSUy7M+Xz9VNiEDnqzDWkDTuPloj7NXZJNyjPlgIwq3pYNOuT58K4rH5sKzPp03y
6UADJ442q17VIFI7NoQjC/vgMtG1bkGVzx4dmlleHbu5vO5uxMwP8CMhL4RXHu10
micYZQDJeBrN22jKFGob7xSM+HcV45HeupNGMjNnLy4TFNCaehBF0spZUELyy7Xk
tjya0BlQ7RJR/8QeRc84b0XqAjjdq789HVaHijW8QGJ49Q44ss+3/UsN1ScAQAFR
/H2uHelXviIhCs/4QyJ3DylcVK7zxKhiPycsCEFWfkpmbK6O2mUlEpjRO6OFQCzW
d3t2Z+7A5buAqKhDKuPw5nXdZ+tHlb5q/ClUaMcc+4f2AbQ6/obXrUw58Dt6PP/e
SWKVHranpSmLteWaLUzRilr+b0VE/MT60b+NYh76X+/FuJsQbRPr1PVTZWGK8hDq
a1AZQgHGC+R24oEze9sgNM6/zvCX5BhlLYrmrK6Yt7kr+pOTJiaJHs43LYRyoOzD
RLHjYAOKXUv+YJWK2wk5hWxeG0NQ2/pWCjWXifhR+cV1oYiOTNSAYPxzozFDdT9D
OribDrL+cQ/LJLcl4bM+IxJ/peIQUrml43mNM8gcbQIR2DchGazWWjBf2Fp2k73X
rpyV1tbOZwf+OEGdK51NO3YiIzlN7wXgNzqaC6Xtc/Hk0uGliiEU5WZ1fSLRZSxV
qBiKe8TZIZ3iY4iToAilkA0WGUmyYtAfkTfOqw6XB+3Im2kce0PS2StIDbTRcBIS
Gy2q8xgvOdB74bDEur/nAFoPrsSDOF8T3fmkT4EauY/HSLJNHAaOGp4nRS4x6MNR
TiEb1n2I4NxD84TB56lyaimoK/Mdux5iWm3w4ZoaCTAGtEo9zPb4w2w32OnhJiv4
D1lT38YZgu6R+vcf+BVI5fB84myzElmg8XuSlszBmPHwqtjF/m7wBk5aia3lSMH7
TRmNDkZANBGwl6/QH4vPIxddmw0M9BJkc0qEqDdFOl83Ceb4NdYS+Pr9L97L+ZHE
ukFqa6jOE+u0m1evqW0YnbTtBxE/VP3XD4P0+wy2+kTu3HvB8uiY65/CFRu2xMs7
ak2qo4Zz+jdrmoldig9sDuFaODo8A1VmQcL2stR4c6GCnvzlC7SjeOpJizCAolI5
Itg6m9kkX5mpVmX/q2Ays3Xmsw1I3XipKII7WnxTxlrDeDp+u+OiZDIU2ox/RCdF
upmfai76LjgbRWne68D0+cr02VxuChfboKI58xG5SoqnGnS7i5RCxue8njYrYI+s
ulvi8630LPKLDy95CgPGMqR7XpXhjqtpC4VMoTbP+gafdqu1hQdbM5P9wR+97ztP
xedeI6UOR2NGXMY9fDCqS+xvEzjQSgU6fKGoaqkh2rXWTBOgDtKI+sYSUDIEUmvX
wJ6b8rSnJrhVteMwSCaZNKWRdUIWxhvFUls82/O+HJ6cSsoOdJupiRIOxUfWFCYj
ohSpsSD4MAko31SqilwwYUFSGRdQJL3pnNTeuvG1e9zaRz4iR23TMaBzlNn7o1HH
BNu0Rz3c1N4WaqE96VzzgGgbLeOelmOHNQSn5oo7VUjfLuvpgKNBaVa3+/jsPz6/
cvlxf97a9yaDha02X77JfYprnHZH0d8L1wyMnqV1LH/BvAx3TZk+Sc71vjx3oHy4
OMyuGP8ryOf1j/E6FmeBekYOSdYK0XWNbQsB9TI0hGmstf59DicQ9xTB3cjoMZ6N
AbBwIqBFXaAOsL7kwvZx1fGm1p71PRCMIGpG5pCr13ukMJlN+g/eL+uQyVOvZQ/p
jdZj8+tXsaDwke+FgMh7K2bbVceJX96jBegGZSx+z3D3EZWjFzMwE4TuRcoFZfM+
UeXpxpN+mS3Z/oY2vG8DouXTER3LU4U+oNl5jRM2dhxX6vItTH75xq0xk1ij8TfC
09AIzJmsiMOycaz9/ZUmqT39Yw2PeC4shX7R1Y0fSfRyDg3qaHG31v63XX6j6WBu
zX4rT1cCGEF7OOO5F+Mfx/jc1q+HG6PXKguHVqgbQAImv4RX1f/zkNsvDEF+4hau
PzWmkd4q5A9ymvsewu3lh1wHQxf6wAWKPLexBXkSx3wDJFu69UN+DezV+QsiMiYl
sL1PZG5td7nuJQpaY83V5zx54FV3PziriA488XweqJryW6tzrbyeubD4iskUjaER
USbbdH6wkIoDFAHRa4PdiKqmcbZPJIElgtJ7BtuGe8sGYELMADw75KU2GkQ+3L9N
Bt1RtzQSXi1FyHqnyGgNmhh448yoV8EEo9t7VH8UlGpH28Cex/MWkQEOi+i2hcYZ
HId+SEPI5cbHcDfghesmknp0ScA2hJVzDeIXh+lOSOFcOI7VJs1aGV3gBGtAEOy1
8cEBo2Qg6X9tntpU3MqaPWTIElJQVgGKbfZeQR6Oq7komJu4bJdaajGRvzaI8UZI
c3T2Cs5Hcid1TfMzXKXuuECuDC2J4x3uL2Eu45tC3Pcb6un0tuxTpkrXLc4bNPQ4
MR0fmH13z/e+SlAJ5Oy42BVO1Re5DMtzaUKEEmLhbWDH68WT/mDB7QJ/6vWEYOQV
7OrpPIhzoVHv+yocE1n2XUeRxksPOG7nvWIsnB9ZHeTlUGjoKrW5djrVz1T3DRPd
9d48ju6aKo89whsR4Aq092hIh/ZBT/br9LgNiLYjVN3Op8IK+PzK/BV0Ri7LKkoc
2upLWttEfbdIFU363Ls2xuiHYzqL1CwYp+Xhw70thmNxjscQYiLjgCVKtPK+/R5r
QvO44Xku4WGWobUxfHCvX/fwmyJZiku6Iqbwl+O2SY8Jo/4RtVcgs6fDHqdUDRzN
OtXVNvjvA9bcw8m3VYnqv91yV7DLxK8l5xoQ3aJbxAMD58mpM6I1WcO6rOaaB70Z
uNfkWuorOXCQgIBmUtlRbPtMJdKQJ/7CB7j16trW9PuSXYUnl6xLKExzWvWYEyWG
eaouAAaWHDdrVXOGF/k9xNHGjjyNLDuKEnpwmb9uAfgSFvdRyeVa0Zm2DJdNLgIV
LfExtosbjMa/I3Onu2WjmDtJxp2iO4AyVKyoUQTjv+W53bqZSmNbwTZwRnthjpyD
rDJPDEIK17quvC8D/KRQ0XRwrdMdsHMU6GDpn6YlMZ5BTHPzszvULjDSTFg3w4z7
DjIiPyf9NHz/NThe0EUs86EaFs8HXYyNOlVQgGjJEngwYVj6yLnewVIYuSIOjpzy
eBxjleUidITJLXGZGWmAARIcD5Iln7Bd7pd134JB3Fckcevt+QmiVfw43lGbg13j
ZnGfWQ0PtzWC6Kz4RV25KB1aWn0Cmc6lgbQbgSZ2i4qJQfL13KqSkZODk+LYMco/
Pxf9FNXDemlOwE3AwxNVi70p2JA6aPRUrK1mb5sCoyvLHRfq3dHA06bnTxPTpfja
IW1jHm9iWm5S1x++h4N0iksBiz0IVW0Yh4d8AZVmpQuRuMcxEW/V16pDzhw1aIdp
GLgCgoBLrXrfPnAYR/wtFZ9bj0um4OJcluIaJCcvaGC8RTHCHvZM+fsdwBi0/nrX
TuLO42ZcLh5u5xEE52bsXs1bgyDQNLF5o4hdedr3i/3mNGujQcMjKwl5pDZaJaUO
Ugd+3UpnKWigASwwlYtaMhNbAQmRbY/5X1H1Jm8sFbwDMH7m+54KSt3P9zTQFpWu
m2/ljN2uePn0AMYVidzRq43wbTy8/QEndF5tuCZxSsl5cJ+hz6h+jyZG4x5WUvlL
eeWf55xCL3Tuc/XWB0G5rbS1Mjp8DUE/Iugg14oeJ5i0BFwFkdZ2vqBexJxT6P2H
n71zSJN1FQtOrVs0wHJ1o2bMpD8fb+7RFDLEcDuSGL0o/ay7VZvTtNVqSnSdQMYx
Gpxdux217yywGu2MOz/FYzxHL2C+DDNKCPu7E1nJM8pGKGANWmFjDeM5rxFgYS05
uTkuVyu6s1weY4KTnfM+eyWqGN5+1jH43mtVY+HYioWg4CoBqPwTbKEDchKu2zAc
jUdOXcul20+G2Jbn9AAbNrpzw51BmrtdHhDK0EEDMUvCPzEG4sUthtbIkBqa7LDX
80gJ5amayv0x9SeoleO9/VCICiJM4enJr74aKeXpAmGVJJVzU2NnjcztmZ8MmKIk
crQWTT9OTRz2cGzmmUCJX6Z60VfLO+H8vdtB6kHz6XjgivuVgZHjpobC8rSS+UcS
vDU80t1uG4qmmsOpH/nPwrgJ0+JVxyvmKTOUfV/zjrawPn2aAsWDTl2ZrTLSEwad
zF6KwshS3ikRGQSSWUf+bdhTSM2f54U1kT+KQM15RGcnwPBOGowBRbhVu55JEXur
vVoVWUaUyOJ0oje2DmUhFd6f9bQ7UoN+1hf3XSqZPmrc5F08zK42dDeFIIcQDHDI
hhyHhRhaObdWXgKb5C142ct6iaLEw+cxYguHgLf3V/dk6Wq+kpV8WAVUfLZnXir4
lU8pMKU/qhEp+zN7VEg1sz2UcphGJzPeasnLT34b+JEK8SR5fsdPIpJ01aI28dh/
PYxXCRFpeA2pkSxCdDm5G8lK6tJjuUnQh0sgdkD0tFc+9hx/RMB72iupXYb5hRHR
AObFWVyLEaM8296v/N8H/r0F5hyBUwP24yyuv2cBp4m+DPVeXyOKX5sFnJgw26qn
EL80/MRa3P+qW23bouWxg6VcmhFhrfuEN8UO6DkWCcPhuYY7hFhUG63t9g7PLIeT
5lIuptNcUdZsUdP6XwHDZkhCoZjmyOVyHnk0GNWDI2gRW11q9ZEQqqFH3b203+AC
Pz2fhFaeGEKT2Kth524rhOKNF8NyLhkHiPO5PI4Eda8khT80n1wPCudtPLc3/gJ3
rlFo8lHfRGhkVW5tCVawloa+jWBrpqc+MW7E5qSGpObmHeZ8IB4rYLbULt7VMQba
FmFjXpmqZiXFQUukdUv6Y5GCnLYOSgGYkjJT2niASG6AeFb2F7r10fLzSXmLEGR3
4QmZsxSvvgPbLHE/WIzepcCdnz3wNoGcS1o277+pK0VSbqK8X+ZcG9pl9KicolOv
Tude7d0+pFVrPe6R3caglznUJnTkJ+VN65h0gq5eKj2n4jYTt+97fEMo696ye3X8
ZKzvRD8Uafqf8+RLFuqltob7sZfwdQMjHcF2FN2F1htrPJoeLQ6D5H+y0WPly0ni
ej/VwH+WOwoEJ0UXHdnJqP5X+cKtGPMiiKE5sDBZncv0L90/pyCihP20SPPZwrQU
avD0NLaXwpXzgcDqPHcYd60klsunm9YDqxyqdvFoRbi7c3dW0X35rlvOext1OIhM
ok7sXjgp7Q46JvkO+KNySI23gqDXQb+VPmY/tFQao8S9wNijXF5XnlMwHV9jQJBX
0wtUg4UzuN3kGQH6gFSkzt19YoIojR4eBV1kMTJ3xmG95iV6LUB8aAZyed9LdSsw
66ZcUGZmsHyjjUgzlcNJXWWvMtrhWJ+hzCCLyCaQ5CL8AcXLyc4FlutIB+S1KYeP
MUyfZUkJXOM34YTr/xZSx2gUAQRZhZGunI85xaRX4U5Ew5vqexn65PDk3Wb75dsr
WPUHetLetdt6pErttzzDCMuit8XRxQVnxQ2I/2N0N//7BdSUMcrj7imyohQXn3Up
VLJ6W8svqnSjxWFdYmau5QoP0psbYZ/Ede+kxz6IInNOZO4GBdBGVNJoq4FFdZsX
mrC3pdKRdOC+8xmO/1j8jU9NbYLY6OdGg42ewpzQ9rRLVzmnsr35I/SCo2JhMC2H
G1gNjs6/q9QIbxOmpCtl2okqzLpSgxq68ROWe/eXjJsLnf0cXUN2AThVGjb8QKER
ZjueRT14vbh7bm4kgz33E7tiiOwBrw/SsuPRvxDa9+IFY+0fvfLKP+l20GlyeMDP
VlcJl9q4Qzqz4YFZrzRAJna0N+ylyd1mrJ1DvkH6KgbvGkuYkkIBCf3A3mUv2FXE
y3ukSa6wZA0TFV3XhTpAsVGBToMVFb8oebONGNDX7NDI4habHoLa+tpXsb210Ou3
Kzjz2O5bctBmivYh/tkd9BDhYlys8YiF/Yk7dbJf9fsaft0dCIjjhc4K3OVoJ3Yg
dffjHVdWLROizIe2w8zWsjRqKU2id/cHZPWp2BNuPakp45rpqi93ksuMk9HmfVDj
5uS1s0D9Aqy3Psyay0EPDGhDgKrq6E1a2VVhi5EiHoOpKovRn7feiZBwb+H0tdkH
cxEP2WvzsHXY/JwX4SF0bGRYZp8c4IRzMOluWIjrdhxxpkWKj1oOYKxd6uFtKObl
p3m1/fQx009Ybxsf82C9ECxD/WPxH0lRYTaVIWtMrQr0fT/gJUnO3vQ4qs560Fbw
IYKe4MZTrrmjZJLqx+0iKRHgc/u+/l3sYf52nCy6vlzLOZK6kyecNUj+93As9riY
YgIQYiRxFCNgKeQ4mGFYK/k+egUIClTsduh3KQZs48g5a4vYpqSVg0zaKkTHSGdk
lBOSRwIXvc8QaZgmaFA2PjVxwUcSuNRh0+9U7KTM+9B8dIn3/fZWNV5MPVyiomPg
cyqAQxAysRORRaCwPPAHGmvaq82e4LWD2rqAxs9QQnLlQvN+fTGwErdT2ZBho6hL
qMsR24r0DEOl1mu4eaBdS+yZ+RqIitlo93AhzZZnBZBJlEFfS+TRjHPiXXjGFqcm
a1PaXdynfkEXCsNIh0M3/8IiyadiwYc06iSpkr1fhRcCqMT7knCl04fEcL8G9b6u
mdn8WdqVv/4nf3H336wUQOttABUYdOCCm3CjO4vicolgPlREJxXKhy6C8L68GsOm
WHpjRzfr2NVZHee9xntvYdfFgKaeWDrB4aSi5avNEbmM4eBFwFQWS0BkXKHUWt0i
bKfhnbQwT0x3pJ/H4swUdgIj/sRw+w0eBPBuhezmM5GOjQinzM8BYP7X21j0g668
bh+0RxZNeuiztGqmcqdXcTHzETS4kCsDAHQvzmfl7ODCCZma3Mql9v+KrhhQ9q5o
WWqFEY4D9hWCcwOqokWpzLN9ct45HSQTqOKvHAFiKdVoQU1u7Bg0EsrwxYAWxsyN
7xepzIs3MPPsM5WjVadOoLP7vpqLHoY8MrHopeHKKDTMHf2BFkdJExORqnEgUcbl
eGyz4jA51Y3NmHWgbRpcmkRyl457n5mIPh+fW4w08uPlTYobVlRPxAuR39ktZOBh
PwWGd+Aar19dP76h63JVADdhGns4LO9i9gpj89icK1JjtvisW+mEjzHicMj4kdCl
h8ZUFKAQFv6KtwKFIjLlmvvOFk5EbmD/TqKm+YfvbVFi9eGnE1p8J4wS5PvHZUiu
7p6lZ+sKnkhfJL0FFxLGjIWSZOCf0oJkxpTVdZU9/2ItJtCBDAoib1q2kTizsDAE
uZrf6uj+eJWZuZU6c3fFkYPcrMlZdjR05pycrZmEStlKhCKS1uVeFZ/3L8v0SqS7
6XmBtAOdIDfDTnGngOMZfrUfI7hVATeAoay31IEJfHAiQvZc/U2bE2dH8l1e9wYy
8I1jBi/CVtQXQnK5KOdEAYnQJ0tALu/a6svZfp5QoPqn+usNAFhIzuSkGuSTpHYK
O98JTtaX1yT5GWAuNaWGp1y3ZJ7MfdooFPgvkVokEs+LNH7cHdY9Qhl4lwFUqdGL
nzL2DDWAdz6LJ7zYG6tJVqWTDu2i/s7msZy5vH4YlFZSIfGzL2CijfH0cgu7NQ7+
dmc8eu46Mn6My3ulxgZu+Mq4eiNOaU6iP6huMKdQl4vMCbtJ4ZkG9z0dcHAI5v3b
PM88ah7NkCWG1KQ+a1VYBGxskkAsq/oI8Q18NwA0edlzgL++cRKLQEVcGi/YTzfP
98SQR9pZR3sp+4sH7yyzcAccalytZ9bFv6wQey19CTdnkzDr8Ry44yeh5uEclfTQ
NEPcN8hCygy0PzJOp892BcwP601o4PuLBcEqocwnf2a/wRYG2QHZComqKlpl9bKN
tfynQZFs8wtTQad+OGToeCnta1PbJIlNHEN9xCh3USx9m9KhcPtXRLbhs7xMIZEa
yYh1ewGhUR8C37Gmmo0Vf4wXY7n4dsoq8WZ+K3cdUVUPjAgCGBni+Rzd6mFHyo3k
zlKVWFurCdzBpMH0kQQ11D6u6AidclCkLIr4qj7WahpIWiDFhyeAtedzyFCksqfW
ZJiznMzMZgbi8VXVZWdsqVpKbhwYLvZAjPzxyK1EbOVH+0CQrb0UAFlI8zZ5rqpb
pimveuPJfWXfDPYwv0itUdhXUNU6ZBcJOn8BZTSnrFct/6dxZIf/CImvY2A/cG0C
J0NsfafFQQ4/jVUdRZ1iJYgF7OC4LzGMwGn22yGcxwapS/QDBIqzdQNVhF7cVDRJ
jneIXxuMhNhXjc2tUMfNCF1/hkk//ZBrG8xEPe9ucbJd0/ZnwhegQbkdMYl1ONO3
qapfi990E6+hsLmuWK4ko01DZ08FxcAvQaKuV1s9d2kQycW0ICYIEeOavfv56SNw
Mx5nt4N5vijiPFl9SjF1uLrKIra6pLugpgwa8/QNC1Fwhj8T8to6zq6ifdDRfiUK
qe7O67coYEnClz40ZNJnxK0qzhf3CA3FG6SiwTKAYjIiLO5n6n8EW9RBo3xsuMHj
c4NHFBJ0W/bvU2sqPxwqVwlG+zEeKMinVgS2plviGOUgWxCNOzUsRleRGacgLRa3
ibUbF4J6pWo5D3pZLZrijaWPntk/uOi//iYnhSy011dpMcxZqVae3Rr4MifrBjfG
i37DlONQ0RZz7UcGLG3yGU2gO83NK2PwWzjge8APlb9cXzJrM9brLtI+YuE1/Jny
T+L7w/Ov4UQLfTfeUp4IH4KXv48iqbl+EpFbfCpXKbEo+SH7XSVeo7Wn8SdoGW0K
y/O5lcUfcZrJHe7oLy5mwi5pIyb3r4FGgd4p0kkKSUhPNWuO6flZuX0g3JOciioA
hKZThlPO30ktf1MCAdhYxDleGeVTlziG2Qc78a8r9yOaPU1Ja6X6u9DYrYp/Uud0
PFqs/EVOLOEFFOktzqoy+5estlid4wVSHSC27j350MFGkkNQoTU69PlN27yIdcOK
PB2Ys9SfJ30cHdYXggk1Z3s30InYcqD74oiS6yg9bIt9BnW7n7N3GSfHgTrwmy3e
x1S8E9pKfPhbjzxeipNvgR563rGHsXXzMinTFVymZXBf6a2m1U0bREI+YzdTfrIJ
GlM025r4c+wRVFze89IGddzNciCLsdIiNkxJXb3TwptLKLCKifxq7ABJTEJxgCzL
5zwhkJWmvfOYEqNzDOrCLQtQN1UwzFMjp1qrVIjz/jwqHEEMNtsvPg8euT6icWGw
a+x4bjH8FJy9Qn6wCssWzTT4FjJS7P3tYV7mn6Hm9DzWuoLbuySQQaPj+GCDRpF0
IUGe7AHgSdkDF7564oQ8TOjGTj8uqa68P+ekDCtOzCojmEUFeW/WRFs/Ag4iECB+
X1JQgxogrmoj2a9ivYht9sIIjFS7pZHijpO1rf2bW3iZitFDooTpWERz1NCRR/mu
4n0pS3BQTkFftTsziWycFFdFUX2U/5IyUK4ALbe3YP9aM6TSvXGT8a6oQWtEDGJ8
ljYBIRCuj/GSe0fVU2cdF/t879KxQ1QIDUO4T0r7jb4RPcyPopFfSt5hAkGiIHJa
B99S50U5wTXeymTs/rlL4W3/sjwKax1QJviqgexm+j6HA2wvPXdBu4YWnVTULxOc
VegA1kB6khN1wMk+pxM81+cG0Mxa+LoFY6/ipkfgeoLFhQIJnRGWOOrIX9G7XKpr
bx+3sSc03JBk/oMK9i3lViRgLbEo2iphhG9jTyVwweTU2qQ75vo2UVrHwx91WK0H
1Xs/jd3Z3ztRrK1oUcS4Fsc7xZhmGSu4n6pb7CNjhL2S+fMkndlkLAtzUVPvr46E
hCtrS2IQuzSffap1WH1pj82VFa1cx/p56qZ8/VqiF8/lN1U5xDz8xGHdnXZmx8Oo
GdD4g06ACH+CeBT+BS7HrXWrTyjuKKFX7iq7krbpFjzpEUi62sD1PLNhDIiERllW
P2ONkIGB00L5rIjOBCg33Ld27Js/wLqXRsMwjlmgPzSFr+4yjyqFRHS3EPNaL52G
vyct/PhaNGpLsBgmLs5SjTpYGicksSjRcxwAs6n591hMqpjysLd3LT8sSpEEdvtE
5UaUyXFxe99Ytj51eaB+dESzd1xTsKn+cSEAG9zQxrgrr2KY5SzZhp6VjTljCuJg
92VC99jWVAb/zdo6SZh9Fs7KtL2RyCbzuZ6qPYUgBHUwcvwPNcgBL6pi6IpNLgsC
8Ym37lNuWup2weawWjw1flKH867wkxSxbpSghne3dZtuJABt3hXeRAYuKfoOwZ+Q
ybc9ULzyTKpt6UzBsQQzByxdzi5VOZyCqWO0ar0+2XoKcnH3hLr/OAK+8QllJGUq
YLBd6c2skR4npoAnXBi4Uh6M2dpvGupfFI+dVToHNN+DXuAwDC8nekpn69zyqneq
ADCM361l8ng3nDw+UOBV5ohEOGcwf03dNvyWhZ8XOIjDyZn4HftNGfmF5/djlsBR
naw5YDDakqfsQYV8dgUiOAtl6IfkgAsu0k8qv7BuDAbB77w0RxDZvRrGbxOzBGbt
LYPxv26DyNhXJNxVf0NqS2ke35ODixhMPnSu59S7JedH+dpapVPuZK1Uu6QW5bba
20//DwUMjbrjYWzBXMRqtVPqlRqUARBTaMyoDe+/UekP9X555sEoDh1vTC3NaB0Q
R0WgBsS8t2xVB4bL+FJpOAZbiEm6H1g801+oyI83sRdr3O/TPZKpDZrwen9w0ev3
3YevLxdTKhfwKRfIXzXyxznJ6uRUnKg3eO8P0cp13gvUn05mp4c2swUKZQILvIeV
2se7bKfqwO4zZPe+fG8h6k6rC6iJqLW+lMCzFiu1dkXZ6QerRY95CEA6/F1fIqIq
Z3Y+XymnOnowUQUixtsc0ISNGG7Q2aRyvMfJjwIUXiaTS2xr7vcBVudu0YrhHLyp
uEfD0obEB8VXRNGJUXNribvcVlL79ebzlzhLPjaGSlqVfeYdSQuk67jAK2qEfe/C
CFG0AqpGzlyaDouO1SI14Dq+EWQCbF+Yi7eUDgbsPxZ816SK1RdBLWDIZZSMmgI2
qUrslgVZC1JKisfycwsWRPWzJG5EwUZ+UfLT0RPt5cbLZVgUxlDqW7/ffScpExrf
x2yReKlTrx0UVdmEKe3ei7DpkCMZsOrZTLrNmDCWU4g3JvWLsHVRo1/IYxPbVh4R
iqOG5Z+SqoRJsj9NoGdg8HTWgwMSNrrTSPEM5FJzU/YaGRG+SUsIGj2MSy3sctv7
QRr9I2bd1ew9I+latdDDoD/s0bsKyrTohrAtDwDimHf9YvNMaloZTD98PaKIzn1t
ZZizQs8mQ+rv/nME0SnXhXsghK+sP20O/oM/4sehaIh39rJPerPp1xn9qLU+itNQ
TY1Ws+0HhufMrWxI5USdeWPj9rcf6i3uCLTBFjdlMJmXXYuFiwqezW2UBWp4tMYp
jMspDGWOPSDTUfSx3t8/Tueg/9lfSg9wRwTcNNrMyUqtz4W9Escin0QXynE6Yp2u
Hi1s04WjmjZ8GVgzNqAr0oxPJyV6hq30PmMiEtXK4Rzmee48+VQgwdYO2lf0YFA2
BYTN7TtuRnYpQj56UCuhLXO+R/IvCIsbTPL+UmFxML/g2Y1He9gXPO359hawkJTE
sBIOTiQ603ZQwe4BPh6zzqChWALuAMesSOiBEAD8DT3GmifmqVLZM09d7La1+KSp
aBzsT9uAZ3VTN/A6usXShU4s9db5QHTDcNgfyrD58gDOablTLVPGCBtN8Ud0MtQQ
BHQL4vR4LXZ4LQDsAR5q0ks6thcXdUcWBy5Sf1Yl32OnKB5Hk4d53LQJ4BZreUmz
DwQ8sQLb3YVMxMfSsjz+NO5rlcn5E11YS3QjrdTkHJTfRuCD4OF61mFO0syOoVEQ
D2+ByiWFDjE1C7leRyK9xW0Dr+n2zNwDs+weyp87eXZ1BS13UlVG4b4dQqhfXrva
X/asVDo4EXewPq7JD/7NKcu8an1IEHZysWkhHOu95ok7T3yrfYDi/pZwDJkx5kkf
vckTTYiek4R89qMhLZhK5Ig57PlwWOf9uoRMitOeioIHsztWX4SOifaeKL633ADl
q9vvLtA0KwFp/SVJaYVO5sJGDsuUIuEkWFzEXCclTeoUlRfXWMuQ5eadEb/RjEiR
iP7uK9XVK84K7s2vSjBNqU+119GrMRH+7g5SWnCtAb2x8qwFBgCjYaipbftCcd+R
BbMHx+ZiQ7eFyslGT61SxuCu4iilKu4cYQ9xhSSkCwgXISI5QR8mf6nJY3g+q684
tnzA3V2HZ/uLRjMzpg+Keupe9pqvFn1FJbrWN99tuB67gSIrsEKczvmc8ze4AJ23
FS+xoMxcs336w5sm4GCpW1+9F/lPgpQaJ8QJTUNgHYFrKZJo3vwZvpZcXeOckO2Q
dn6bL+thgJNHQRP435OkeVynT6TELum0ULcr1Y07cZgbVjFyLj6jJdkI8gEbeaO2
EreeH1S4DJN6+yxb921BZ40L/kLyl+6azO07b1rgfzczrWCF8Md00dCYrpwgE+NE
FELVmW88i+BdzPR46xqYIP3BKa8TNe2VInxeHZK1KGYrZLbdtVqIbfcL4XFB5cML
MBTIPjhvfGKPvdu0VExS3dK+/7khps2/Xiq3Z+0bfX/BA7weYLSRdavh5UQEuYOm
voKRDdQa9lcghluIU0O8kWVPgAwvgfXjH7zMiLWcUkMYQUoeqmfx9XUKVvjtspRv
CE5RsGjyjyVoXsdCU+wro7kMNfLioGz8nZhizVyRwSBX/+u3QRhPjjLeVbkmosSo
0hdoC/a06tDsEi4YywihH/YyJJyW/7xFPu3ykOLjGDBuzYRPtfiOogcG3jlxgIOE
n/ua4FVTT3pW581+LX3rKJ+/YhwtmtLLmGqVVAKuBTGSsaceSJmAtc7vSckRWu97
Jz+7o6agOgtis1AI5sHEHd2vEW+/FPQnMMOPoITZ5JUvM52UxY6TErrN71BQ10QI
CFJJQiXBaPHRLcjxNojINMv+li+zbtoHfFf3y7p8iLbFBGvFvN/Adyq/SzoplfHY
5PvIXNnTcOn3QF8NBSZ/2zaAFKdr6ZWo8gYx9nl5WpF+Gs8TBIRFNdB8SsbJIzgo
LrsM5VoukEEp39nY4SKUBwhGUUvEqZr9gfYa+I7Hp925PpOP2I7ZB5kbhowGecVZ
wulIaKc52BPWUCjloJCVjhuRczJ3e9lYVO97KUUklkB+HHNQ0xN0dmJxKEz9B3Xc
GX5Vib+M7bJzV+5/YX7CB+nbvS4mwAn9GT8yZGGx+EQUMnKdHo+372wO4CgH0C+O
DZcCuMGuIF2+77DuS5OBQ5tWXDcu6zsXypo1XZGA7IaEb2y2kcG3yO5xg0975Dyo
CL3A+PERZn8xmHITuf/SlaBM4qV3ZwEXI2AZOdxBMvUpr8xejUmtcpMsQnKLa/Z4
01O6yhhYD2FM80yul9mKS+JO5aM/OmNcPmLOiRoNXMi6ggiKheKFUQxSOdL+uISn
aigc6Ei6AQ/jFaO/Z9P3pvZj5Wh6veXL86PCAqhju3aOXE108wrao0DixCAFf61Y
vI8T6/34ZNLgvFwOmli9OFg3Don3kdcMIY4OWFn/7ksSu4PFXpOg1WXjw0dw0BvR
llsys9Wq5thTq6ot91pLpiBvQ378456bWwHLGdsXbL/LPjN3Pj+43JuZLLB1hLPW
hhEJLRbEKnT7UzziWWMBdLHz2U8y1WXSD5ScmS+COJbDfoQOh9ZkGn4T11H0h2QC
anS0tW6ZiIpmQJ4SZ75h+W00OVY/cXzuOMx1kNEX5XiV6gjxWj51Hdac9dZzEYZ2
LlztT+pIl9Ds/SLgIGD4mJpOBthheRObJM+BuHwoACim3g7ZtRIbNUwRGgf6gR9P
vVkGHf3H0OYfU3Z5X3phMbRol5pwl5WQ9fOz5jfrjTghVyXPXSI2kFJR4zdfWrEN
AP1Acx4/c+Dmy1CKTXGvDfnE5unbwSUjW8wAnz7M4vO/GYcV7hWKlS83SsbuWgOj
cpqs5qPnMCUajsKu82o4D9w7Ei6r252fO/xyILkOgVjQFSiBTcl4W/qPdQT20JbE
CaSkOPu5N/dGpot7phF0fDHD6TiqAOT+GYIvmPo2/VdtOir/E923mvXLet4lI09a
1+aX1lxEUEBWKmdFvsgUBC+rVn9Omj6WK+OkRmPmMEfs9WgjLu+u2UvFNeUSrZLm
mwiwZfry+sPgGpuJIjVf+escaTEX0LOy3OEFHJXynofeFgi02IYQoCiii4j7TWMQ
lSQd2S6/BEAEWdZpdhOWD6jIy//hI4bbaMB7sxp5gSVoWQJrHHZYewesx+HxIDi7
1+SFOjyqWofz6GD6u+a7NjKSAU8K15IwT6Pe5u9l5/wK6a1FmZuZhtvK9iCohqUF
wTLKFTF5xi9HVIx9yl5UAhrAFZl+tkwex6H9AdzeabHP+0yPYFqbl618rTNFMvYC
9Dd4s5t4T6EU6Gpb4LhuzIJgpZ9xsRhH6V7aSl0c4T73+QSDx/KueAr3kAr7+Opw
SeuL/OLoHyHoo2CYFSyNuXh/696qV2aGiXqHA+U7Ba87oNayppaqIRJiR78v0Xq+
rWnM1s6YFFt7s1oVbSKyw3N9T41fLucMShoMDyyoMwtQF1qKBSJ9DMJIM0i37W0L
F+m6TrMiBgSZn5kR4Hr92qbcXd9wQM1CDdaqgQvx69Q21c8ZIiJHhOvDFwqUQK24
evW3dk2l4Ax7V7yxjjEsugIhs3JWPBB/rN1iGOrkay2R5cuZypOiifNJsLS8W8qY
cECHRIE7m60CJ1kvsmbEGjuNAfXORcVy9BE+32i47JaoFv6FQ2UPlXD0GSfJpLFR
O9TD9DBBcDP2tV0llNRE2wnGlSo1gJAMWCiGuTuLV/4S3N0tTQ63p26NnrMzBvln
AjXBF7wQ/9+2XIaluDwQWV2uCTM1kczFF4uCtqjyjDgEVL2UUerXtnCeusOhKNmP
LEjNHkuC7oMJpZKMxq+awboDqYEscRPJPlKq2zYPF1LGCr5ocNc1XnSFNXK+FKjQ
MAf5dKp8VXlIc6X86Pg06paTTw7XVevDiC1880//Xui0XGPXhHGM0QvC+5+kBaz7
6Xyo8899kFM2ZMUp4s70LlNwx7NvJjDCWeDmFFlMlXlHtSK42OQw73UzoQCzkPb/
0fVp9wDeP5n5hfF2U+mwNTAxnaRPVyRv74ggRoM1nEugkdQms54jej5AjjiiyA1R
+rLlr2PRgKfJSBmL9xVK6zwcoHnvlF9Rf5i8QDhfJW/vFtoWNhwXsHU8x3H5mgR4
ld68oDwBsAxAYghmH4iGYgtAv42ScNVr3WsFQrPBjLdAUNMp7JiErlqQREM2hVAe
Shkd/HlbItNYPM0CUzBetDT+aLmgTgHfFVZ5LAgoe7nhzXKm30UiUI+VP48keFRz
dEfrxor2Ehax6WkXxYANrcH1l530BJz9ZjzB9XNRwg7puEnDcLdooVEgBHvTSFY1
PFnsF9CEWE/BRVyUuYnVEK/Lb98rwh3MnNzoWRD/dHb8b/BU7O8GZ9RU/1EjaEU6
qCiQS9e1w9ZfDMg5GHlcGQ6UnCm/Hk98bRlqCyg8/3ynwJPW08f3PXZs1o7hZOXz
rSZMPZ/1nghxrnJEB1IMY4NcIcuKNRSRlfZ/QaP8ywMhnP4SL/JxrpvB8yLh6XNV
soQyso42pP/jTgN1cvDzUKsU9H1JM6w7gduQ//qG1Bk+nY+JAw3yLMfY0PbadQIr
4lLgdRiqMINdMyrqxa6xabJz5SuL69rYmd3/9/6OPeM8e2wqXf0d23W7HBu6mpQs
Lv6s0IHk1MBVW66jWKdiK7uBnaPnr3ve0SYcbd1jYd+qQJlQZ0KHz2ozZLGJwPsI
nvJHC0qBHa7VoLPurWypy8FbS2Vr+hG6OpgxmrEXiGTf7uYXzNeiJO258D4tDi8U
5iCgov0QYY8c73bDJI2P7tI5ItsMreJIxWRIaXg0RIkDl9+CfBPK2978doVsu3IO
9OX11d8eldklH0jmLz0tg1kSKFLEPk1kBlPuUlefaXtcVcfW0ZRj/rB3SK3Rekh0
RfjuQdKfs6BNOTqoHdH1zf7HPAUjobX9r2VXKU0Js/ip8b3VvHZ5DMoxl5+yGODl
zjlAg6A+RnJ61hInhX8zvCmg37kvm/YOWlTWTdJXgpfYZKUzn+jL7C0BATHmPpYn
iULfvuZZfTnbOpTArwTswssZX6cmWCRyW3+HatdmBJci9bBKn6RWfnnLScY79hHS
G3rgzkIzdMnJ5yQt+EdDJbuO0hmow4HAiBvUjQnptYaFqAzRVfS9mKzBmXyeUChb
WAnwKG7RhU6k6rIwbPl+H/AcgUzjI9alnMB3lZQlZqqQ06xWFabrat048OlwWbSv
ToP8JETxz3YxqpBkJIrzuzQJt+pECc6vygJSycGf80dM8TatgbLZx+D6AsQQ0kJa
+aP/3Uw56c2SCCkdE80jAi9yCSk9+FD97YSSi3jC3SeboZJOcgI3ycy9VZivbZTG
cw07j70Ul69igjfBY5uB745h3ygXFL72lUU0kwQt7aic/civSwGnq//oEg4rFCHn
e8kmlLczewax34wmFQTSTkV90BMja7zd16rCArNcS1La4wElGwawjEMPUOEXA3cF
ZxxPviHf/vGiyXpFwzMQUqCjfS67lovGGCnGl7iJ2Nrn3HEbaw7rKHBBac5jUE8q
WnD2j+u+F8ASdzXntRqhrLZ2J4eJT4tR9BK+G3uhrjtF8lmlOZlgC6L9hvEpJmYF
jF4jpXTYHCWxpLBFXPjpwQrQ/3ziYOqFEP9PJdcF/5oeALZ1iqQyBSd4LQNGohq/
cdRm+TxHRJHjsignTtOeEkpXwH1qfPzwbrlGMgoI50MNqpkDj5M/Yp+acMGsU8+H
O+AF3HzD55ULqhmrEI9uuGGxOs5Lfx7INgv/0hGV4lFkrLOXr/Ycu5tRX8wlXkDO
6lf2nyngTeClSAq7/7njEIUiwsWJ+CriRAh9lMxiFZtB2sV+ggkbd1nN4bGguZrI
ZAe7qR3T5p3XamWqoiP0+WnnLu2WDORs5HxxICAA1W+kw5KANpzMmQVrjnh8TzIN
NYoas8SHVt7XPUFd7kAXuP0kiEVzgGCoi76UyC8ZqXYyeOuWYUpgRjVJNrAbgnT3
5x5VgtfVX2LNG8p6FUIvvdjDzBSeXNHA2mRAA5VPpmIyyGwPF/g4GYQP4dpc2d40
AynsGjCUI5P07VplsONAERzxwUaikGoBJ9WqK2y82w2RRIyPABlcuyFKpn0gU/Fu
+ciBqG/sg4kf+zY05apKkg4x6BHbGE8CvvmmWIUQGLWw89Qv9a+vRhLdMd02fx19
S6e+vGnhJ5nUxS58xc3Q9ePQC9zJNe3/ou6dF+xWV5QDRChx1qGAZL9FDpgq5wWy
ro9B/U2/PZeuxyTP60h3EcJpjlG32dQolHtKD1QC/qjHVrxxlEjHuf4nemMnCDqk
JkoxutQl4fPGaQx2k9rttT/W2a40ZXAz91eXcHSJiADhMVQVsoKmxuWtPPKJJNdl
a1KQ2nsIuZ1g2/DN8NksfY5v+uGjg5QgEk5Si1W6WzhSmK0a+nFqkNNfEC2P806o
SZWTJ38AAOPqTzo/Z9v/czb8pwH36Elr6sDjy3InLkKhG7bBk4+gj4gr/XKfla74
5Sz2fDDrt8c+BBZTo1IM7wxJVBE/cFT6gGyFPJmDY/INGZ2NtNC2VuuiHit3a9Kw
Bua3Z5zYJF27SBj3CFcVNy4SnnLPHTyQ3734O1TbdMIM63rwoUi2+Eb658ZNBEJv
A2j3L6XE34qZlF+TyLsvBup7fD/sqbWV+QRjPjiMr/y6uLI32LUcd15B2hcm4bGV
FgjBrgEQ1Nj/uUBngpFCPDlfD87ZQ+GDty9yVRBDdnDcYUGNaSuUJOAwT0NCjvoj
EzrnQfEkva+7C5WXAaSH/ESvC1DqDYg0cDJOtZTw5oph1Pp2iICUXjHGKMdP9tmq
tXVI/OQZJhAQgGPtbR1gZzCa8uVYjPSaIRPcK1Apr6+7Ca072FbhPICV3FHr4R8F
R0dJbAGMpCH965T26tlfCA0HgtzauByLVQVGf5IjTBZ9BcCP/1gni/ykTWgljDQt
ZbKKxKS7r7D2MTOElCyNaCG65go80Rg22UYLTyyZOrd7s8oRzskUyA1zT580cSD8
KTBq9GCUGAmyo45ogF7f1M1njhper2sjgpiw6nogC7D5B1jbnOoQBFyjTiKbcQvA
B95WoHj5W6KHYCkcPvODnjMUuK+Btq/QPfXkDvjk2j6QTsSlCZ0UF+sEN3ey3hz8
vHLrxI7Vd+uYPm3iX6hsPJUoiHQcE5wis2PcfRPLOpBjMIKbb1Lq1zH3DHVMvWpE
L8dozf97YbjG282ZufWnrBrqHoVEVYa523vM/vRk0NQXaWWuUpiBEV7If1Nk0/0B
6bB17tDMre9JsntDf3D7pAVYTalM/uaDBPIJr/lHjTIsTztEQ2pJi8KSErybCg2Z
U0k7E9hTWW9iJRLi18cazlSDRoboSEbTy+QYYCTY6TvUEKoNYU4/1ALfHZZwjVsr
EPDq7ONDJn/fuqh6qc++YIC1IGNJBVpvEMzkErbwkVb5Muu+268YxMk9K06x5F2k
NXHbUauf9d4+32VMaGewR5jD5ZZGuM/yM5xkEkxYzwQ3nH1D1hJ9JvcnOtzBGDnF
kf9ZTwXVqOEGnlsWgXbQE+PTv6FLOND918M91McoVYBSJ3yE4UKPEdUJgg0PFKbw
ifIKKHA7QEZGrZRxuBZZ3eN3YvImOd3j5vYchJ4K1CwmWLXsgvYA9yzqxKer2nZ1
zkSXom2AxSrAhFQIlAzZqnksi7xaZ5hn4T8XWcUwkz3j+b/mJKzNolAVZlkoiA+P
JJNMDxZAOaKYKGrAA4fMDXJYWUHuI6j+AhLBqo2chyaGWhmOvurnz4UJ5i0ujFol
/t9gwrASLIXD4739Xcby0MQExrT4TuYF5bgnf9KKdPOj6fdd18IMK4iWax7xjysj
LfM8CdvivLdqqxcwfB/Ym5qRqJPPKiooWl53130shEWBBQFyie5m70Wr8peqDFJX
BTj59yJv1slqzkN7aLxHiWdnKfC6ysaJNojXSBvAYelkCmibx4VSNnbX/Rz7qyPd
8XaCQNKMOO9nIzC7R0P/UnSj49J80c5NuKd09G7y27CyaSPN5bZxkbylv7I0fTaM
e269MXEdxAN8b1GyGtZWVTOkEolXNXs7g7hSkVsuixtNnQjaomXOfyPaiAWxl1Q6
rIRDS+icG38gDnh32J3ZPVJ8YOopHz++VHD9JjYa1vuzeK6MpZ4HSJ945i9ZHGz7
5E63ypZgecljsXBZXpTklg2akm7Q+Ti7+l0AMTn6egt/hj63guwLasD9DxjLNDfK
7i/9kOHDv0xks4KIzyExR36WA3bpv3aZHbno5gnYgMKztxAX+YTWFnsaIQ0C/+RU
1SaffkZuPvJmKm1Yf5VH6fXAkvVNI82gmmWl7MXBva+tpNimUHrN7K/yAYGLgVPv
J6m4qGjkKstL1Qk4QTOqmYSl5y+y6AY9CHXqO6HJL+abGXjt2RuHyeK9zKN5j7r1
xOmHFmA21pSy13gPJDUWotoOHycX2+jMIGObyjLoiIq1qq9qFgjnr5T0ikTNgTAM
TDGgfSFvXP2vb/acQJ6PG6QN3ZjqawROJ58alqgNGMomMGZsbF2/GWlMZl8h9/KO
sZomYBQbBIaHNEOziYpQVsysfFpmNTesIVuWhzOmFGacUZAXGFe8UYARwmAMRlfo
LKqi8e5w3VUGJij8uwCJxK7B3DQ53qko3GNx+KlNdl4eZrAAwTvsedgt88EwIdQY
vpOX78t9zj3K4P5HPTjpnKUOxOL1s/kATUbOeZfGBtLkNY0SxviEiItNXJJ8Bkfe
nMjME2vm+DW0T2W3dtEIh+Ta4hvSAGQ3LEjkoy1ZWAP9et0XsRVJ3MnM5LVs6U/e
/VuAhryjA3KcRHYkgdPFetqY9hpUTXWgmqlNdt6W4fIJiZbynqbrht8MyCeRUw/M
94GCZ3KhDcDLOrYmSsYWzCzhFv27VUpP6PeK87YixUJbCNlv6WTDjnCRT94tChY2
FL8CcBhIa6P3Fl5creVBXpiEfhu7yhPLUhay36ubW5HOAN34xyMVFYlkI8pIPAQU
LYAhixFLavS25qV+uivH8uvnHYOhdU9581pQZRUHMsC43KrVPsZ9D68DHqFr8MLa
pONCBUhCLRwljQrBRL4sKUzfxMCNQGAXL9sfZj+PNp7IIk7XCqM4sMJiAMgF3EmR
4nZMNC4+C4uAuBKXo0/e0lQZyaQPxTUR1g9HQHsXaw0TcXZwpyfQCGXqX8vpJ+wX
otCnKtTKZwso7ypSwxakrvgHnxiSPx2A7qM/KWEXHe/q30dn7RysePg+C07qERRG
T2gm0ObIvfDw3KEPziQVMVPnY3LHS5BCBDQ6NnJYg1ynOeLLZ/CDke0AlYs0mesj
SlebCbh98CI6tYzqlo/ub1cTni+OWgTtS3JdXbdaHHoBUU7ane9kO/337vYKOuNQ
ocKCFj2PQdDCTjp56CUIMIcYWQwBLn+lyE+oH0JSVkX3mXwcf8+T7hYckjLqNy7C
9zb57+AMdMOMnG4tk4UtSx4uK3gOPwqAoQE+O4E9eC1RGM9WLmkW6HfPiwvOxLFr
ezfShNj0KGxChi9fZdpaeYL0dRUjc96+RF8POL+3sT7+xlW5YVy6cQSEAhRUhkik
h3D7dLiQAMVkyjxBZK5homKEC7XibHa+YCFvLDoTlNEMTS6JH7nrLtGNaDD7wL88
JoNDEJV46Wihln1T3cjlgykseg5MD5qVF3ubyyof0A1HcGBs50AVHIcAlA9TYkqf
SEKyPm3hSeBzpGw6JAEakfQJqxNA0+m8zP5OWMz2dGRhXmuD1twT05wktBbdQJhl
LpLs7kqiGhevQK5WK6scP3gv5hMYKnRRWV/2vXrnrXcliuwvtwYwTMa/F0y04U9q
teaHb90F3At+hO/mCx5Sg5bS4tM+I/sFf8R8O46BtRa6j8rtFl8ImGIIHAqQsT1K
guu69xkhCFJ0QA//0430RHN4V0QOfBtM3V2ePGvOVI33wjnxQSWsEM60AvVng5fj
hj60lZuf8RfZJXd/NxW/hw0tsu27oBB+yDui5lBAYQbxUt+35CHh8moGUccHJaNj
aU5z85rRDj9V2YlNP4dwMuB8WMzPvqzQHZSeUQCC8s9vDQ8MlqsPPwjb5a/bBGxX
bOzCDA58HvVw+jYlIU6X9PZP+XkNurPJw9kK7L7FVkxsrMDiUU/uTqSxNSSops6/
1fQAexgRinjYGPUE5FNfLoEUT25Zajq0X+s33ANUH/XKBYE4VjrDlIyu/2xrFAAy
lHfx8erX0IVYmpTxyVjQzytwiZdkmEcgsh+AQP0CU3QJOi4MPeJRd6pVkSiDQZqj
0fORV8Ea62o/lO8mRCsTCmxOEV1M8oAXVHFIAHS/n61rmpOydQA8zirIdsAHHjKj
84P7sBIlSD+CcTOqU/lDVCvQS67e1mI2hdHJ4n8+4MuSlkuyzTNfi9+rcEMlkoG4
hjL0UzG6nHhVdPxOaCWQL1dOb5kJSdnNMxq/lDgUYyETA6cRUVPVuQ3XTBzrbWzL
9W1SECBabhtFw5SxIil2sX8LVXClrA30h9uqSMakUSNxko/K4R8C/WnRYHH3xJ+o
OTn8BTlb/0Jiqn1ckcAx1n0vP0o/yWAsa+GiDCO75YMBr1z6ZKZu2DoMNreZ5AQ1
lmwp4RiGtqZSQxMiGEfTOarz7BTcsPfup6eEHiDq6Qq2qAaItGd8IP2/P3+zfzb6
AihMer3irb8aO9crukDw4H4Ra/KBVmUEbXH+6zmg6guoQGt8HVKGYIcGXLog+B9E
POP9ipVTTldZHfB3M6PlVtKkFxzd1n9cTHuB/vYmyBXPu5b7AQicQ0tkmRc4CHr9
iZHteh4gKrhJYmSNJa85AruccdoJ5f0jPbFe0zDCQ20ts1kHg3/FoAw9JyIyC1tJ
RhKWqJS7Dq+Ijo7tLGRq+V1ArD/4wJCo60YoRROVAfcGl4/jdMmQM80nMlvHhqLo
YF4yMEvZ3w0Gc6TXcLuVfa8l5rMc7KW+4Wpb6EhM8HyMKmGpEeAS/kfbnnEn4bpQ
JL1D3nASqQsHLaVX0/Lo14z7gJ4m4vA4Z+C2gXyWyO3dkSNMTBa6AAhFp8FyT7dy
7zzaKzeJH48MKN4qXYR4Loyjr/RHIGuF7HBJQmXDqZLi0EKlUFkagrb9sMNYQoyc
JJTePuwxtp+aIxDy2g35hDBfM4neS06Yc4geunfPIMO6XqzZqAhoiTR5YQ26Eu1o
K94pYKCBhiFEnG/J63C07k0ho4AGM6gUx3KuSnlGEp0ZkARx6DWfDccYf20TBx6U
JhMu2zXAWjmALyD/Uq8cUmAtaZ0jq/2izIBWopVlaFp6IT/hqkS5/Rqrenipc4OG
kC2OD1Co7EnmvlQj1msAO7tpIx1s1qm/yoeTmCLp1BUWSjPaDNs+70YOEATZagJU
8cg/CjkStQF2FLKPBhvknhsQtg1E4aoaFuoFAYqcq0Fk2KNqKKe2i7dUMGSz4AtP
sMuAbiyidhRmXJG+RAQe3ZYoVlyI4s/fvW+pq7UI0GyEAfgQFWBif2bct1b71e5p
uiTBjx7aZvchDWYh/YMz7iHTS4eaEImbe55KRdOHjG2mZZVqbzt0ap5YeEU2nglg
Ym/Z4ZMNsmZsZb8qkM/jgzkB1+MvW3vhEaFDtzxtY+wcW1jkgARG1CbUzOl759t4
0JQPuXsO1hmsqPTRIvpfgdFI5cS+yjv8WMp0aic/r3fASv/m7FKn4BPlVWfdtkBh
RWy9xBifLQkNBurwcxHsy4u5mvEjfkoOpH/eaKHsjrw8su5RgXGMMhO8vyzf6zLO
7PD+Bmq/K7Dh66Eki6KQUkJdyyK5jyK9c3CQbGNXGuuLA5uinbPnrnuE6L/+bxR9
VBs+8NHac4LVzJI6aQtN8hHihZnPwgOXPHkMRZtJ7TvgG3gjNkMa3Q6N90REow0k
58nFZVL25Q24XMnsS+on7MZHEKYer61T713ag9rfS1razQC1eQa9L1Z3j7kmn3HT
x9Yuk4b1RXbSiQWI/sWLxeh8GKEEWMEJlXRf81XqoOISeiBy2pT24b+e0hScQvYq
IBq7hdnlEkk4GYwbEbeILlGRHkC5NOOnPU4likQunaHUu6SMJtQb70i7itNJrcBK
r8YrMOgLH6jCb3hJ2u4uePnxZj28Fn6t9JaeMfaZHO4m2dkTRboeRefPi3exQc4t
3oKuOXGruoUjgpgYS2NrNaHhue5E/tPsSH+M76JO4S63xMcvXTRZD7nsfKg57YHE
cCbDKGEYIwz7HD4rY5I2GyPNmTMjAefEHn48+aoHq1fbC50E+Y69UFbdYQ2raKV7
+UIe/l/u17G8ApnoNPhwtABrwXQ32sIPjDMTqN5EcMEc1Pe+q6JKZlj179l9R9EB
9LcUq/YaxkECBEra/n4oDkaTX+DS2pwGaKJke82WxnngXi1bkcahparZ4q5bsF8w
muIct9vCmjMR41YcWHoL3tEuql+opPTWf1sFFqlFci4T7EF59fyx+cTcRogBDmi8
XeQY0SDiRZKN5F15UilQRBkUAvdiNsW+ORS0ArbsngA1GGde9WN3Z4kN/ezNyAjH
UpK24/Wie2n//0v9muA8ozauzRkJXObMDWflpVRKvna+Uf1DkuEtW/fZTWYDM0bc
SzSdx3jWcaopjOVz9RSLuE/sfINrW0io2Iyekmyq7/J3rTvbuiw7jJF8QdfpissL
+usx+nzIRUfFLnbWM/4kKUvbzFjdDBz/Z/X4gsV8CVrbEhObLHqx6fGMQYxVDZBI
3StfBDl61enpzjTS3T9K58VnUZy2P/scKIvb9H9EtlkpS4X+lfFgyVojrNcHu420
p56hXHvpZ9EuuJgI+r+/a6fBFRZOutG6ycG8m5qFGWmmMgIZoJlrL9cGO5+k9stI
qIHu2jIVq43nmEhrZNF9I/rA8RY8NkbVm1L0A7Y8PAAH6Dpvjay6K0j4KP6yldIo
vi7FVyRlUroxq+RTlnIhiaJ8AOGJpo0KGtmqLJtgMQ3BOp/zhFxa/dkj9ylNjycT
0noAHqbS43HJ5+Zg0NkDxeuc6IDJc+Ys87ZIpjPd7htRyLWlYxbU4k80JUVY5tGc
wZrGU0HqHHYYtdmXFn9MVEU3C9hJXD+Y1CI6bLmgp0X6tHzQh758czThqb3Bzmw8
JdTdAdmgBEZlyfutCMB4DhV0bAQbhrr2BaO3EufHSd2Sx14bYpWKvvY4vwdlLayF
Yd/jXzBsbYQbQIER1y83mOyZ/OMv5IR7PqR3c/1klgTCvn65AULlpEaCSR2nQG5V
asrKSwbZxZN1TLfSyCQ3tG3+Qr344Tk47uc4Bqd0hDiCaf+NTmiXB3FVlS8jWxYs
X+Tte5CAdnZIlGL5bBafvaBF89y/V3orbRkHEDiSPTRwkn0d5kYQzXgJmc3UhvBS
MzJHQkSjCruzxkf8lhemh8RcZqZBtmdVWgRnWHyBOQYEf4R2Br3z0SUsAG6WoVHq
QFaNAnNNTDLxxFeH8yfDD2Gr/MivCKw2/iUp96TtKY7a+AvUK3evYSvxOEwEhgGZ
XMOm2W3hqI3vO74ImJ0j605afmkvJ2WFoQmVru97WNnW4IMM0CZYQY7+bPpxTKsg
uyJKSC7zDWFnA5mZBEJKpqFijVQ1A3igpUXanVBHmwhev9FRqRIKuM0dbK7W/7l7
SWhY3PzIPDmpDC0793n5s+JQViSqyKijFZTQVoW8TD+iPRUbaQFKqRQRjJI1KNnA
2c5mdw1zVyqEwJkG50F9lPAsk906CDXt4auXlKAs+xKPSCLIs8772xdl2Rx6O++R
lRvfwHbHj56wkLTbsUf1omdU+R5qMHvCIuzqR6+/e117H+qHOxMKVL2UIfwHJ2dk
miXRGnpTd2WTsRJCRT5OYnSWt1xmTtVZIC221ds+Bg07oyU5nYDCZqqd6LsM+ckg
AkqLJR0IQ0gERbea8qj5G0TQV7d/knp+RT1Y+mNzqzvTafTsYyy7CokOLIyK4BVX
V2IzgoL2XD+ShFdwxFR81nZCWCtvfhNZIH7qeuI2k0F0wdLqrBAhKT5B9qADNmdw
2XodMR1sKPl50BK13cO529YFtaIX/wwX5BFvyzt1sEo64KJhOYmvdcvdF6NxkTwH
y0N18iP1Vk23KmhuxrFnskhDsnlHA5IGeOdOhI02R0rVw0K/MgGtGbiPIGX2WKpp
jMWiX+fJL5IA8t6R38qexd06w+dWHadIYBVSKn42KSDdkJd2FkM2CZL3wzF492AW
CNHaXDWOlCDwY7MV6fNOYqz4Yc2+6s5hLhQ4ZssUbEqA2yeOTYKJjxI8NgnvITfC
Yg+FdelkqXwO0NbfM+SYMFbav6icVNWOWr3mJgkFEJAE5N9ZkzkkN+Ksqk1ST1cu
Z2pJSPuBWekqIbrIJqelUc94vGbVg3z1BWPwNF/unUQuM2uo0OOoOf22GkpM2IbO
nnH6WPz7m90DFYPwp8WMcAY22V+ErAMNRN6QedQ1ngyJMq6Gcp6iZPkoihZrhFYs
8ibY1Jv2h0e3SZGlNmA9UwztRzU1ywyymLpbq7qewNEuOPZAGqiuR0VS3xL85zbZ
C48fz2Lk8DWJCj2tOwt7ggmih9OnNFiGsoHufUKvWRsGrCrzFDZ43LnWk0GHXjHF
H01N3/biSYjHRQSJzw4Jeb1pOwzBEo/INZ+AdlVwmt46DqYEfxekdn5FvrVRDx4Z
6CLnqRhUWmUVRlP73ho/gx012ng0IJdeCtobqMvuOzeaZYMoE3iYlEVDuVAlwZMX
UDxB/TijvsK+I44nVv+j1MCsuOk1IddvGAd8SUGGNU3y8Xj5Dde0d5l9bz+PK41B
kyHUDDmihTefZ8a/8qW2jVQkUXEgihv6+38dXFCWH1BX05PNQHNHj5Bm6ZBYfAfE
M+dklSbks22YCwEyKlzKM99GyWoPwXOj3NwSefKyn+gYHoLBbzBNg+PXgOPr2dux
ghmea7X5YMviMtWUznPgOu+YWJU0pqaW6BaMNfKSCVdM+TiQ3CKvO3riUVoK4RkG
u5vUVCpa0OsR/ERPBWe6oO12hsgcouU6st341FHKtOGkepaEkqTdeKIVq6sNXKJK
6dDhktOn2rhnehZkoKOk4+D2HSanvG9n1mquNanckiOtuXFM4b56/fLD/qY3JH5u
gtuRTnmB83WnuGT9A2K1AXMyzYiftvAi0Ug3lDuRwt24vxVn3b+L5NB31kA380FE
K1CuPoMZP4gfgxuit/n0J8B2kMD5lJzF5SootgMJy4JXfoBJZOk5uzLOkSv+A89c
9ijcMcfuEev1sQkPNsfcTI51E/aDPkx82zzqeaMHYV87I+O9E/LF/aQ9iaHrQPH7
buvSQQK8LSkZD2oRIovUIaze/vCO8hjNi8VoYxyJ3onEKSWcFDiByab3hf4+kHNy
6RATOgTcxtdtE8HMUnH1o/eYi/M/0TeUjfgl8MT7PI85tJmi0hR0zEACXIX3tzM0
mFwtLJAVQvZf9YG4GvX6qRdIl3X8rp4aJ7WMMcTDk1hvyAZksEYdGBXJVErwDzQe
T4mlR8edJ8s27GnSE7M1FI7RGR0J79KJiaWqlqtr2zg6ZNfMrfoY/om4ZKuqPT40
HBUsXAtxeoPYmAzYfn0ZhOYVixUl/HAJ8SYgFsQTDesZEg4kia9hSlQc2WcOY2w8
bAJjVcv31v5whrYgcf1Nhw/l2H+Y391oKx0+s6Kwi39ENWo7cVsG9ohLaiBan4NM
A4V9YczA+5FVSQLUmahYN9TA/o3JK61nnkvQh1uLCu2p6O4uuFhsoVLIoK9Yqjxw
cXHIsxrm4aNzsEqKjiD9nmQ1kgvnzsmblrSySY3pRvauU2YcPkFKMEngxWrshr/m
M5RHhvwoxHtUuYFvWzRqqsOOgM1TiVI9qbwsgky4e8hwJ+E+ZFb5jcDmP6RXfk2M
7QYoCy/Mu/OxTRcb/otTkSBMmuefnEI8Cy6Vr/xn6qENE1yEquHiVvfoiwEWMLkI
v64LXhrbY0RbzdSXi3iyh+mADKrlYW3Vt20OUpZLFTRKvtcNuxn5TP4SAC/wrlU5
BEz9/8U501i4m734A2ff0qwEFRXWo6iUuUP53PG5Kpm1GPncj6S1LvsI4dFXqUnF
VyNDrB4NfJ8k+0AoEwyihBop68CFHT0jsigroEZEQgMO6BnH8mKPddn1pqkxE2fU
uuGhxHSn2UUgvlJ06kKdSVsNkhE5x9tbS3GR4hK8zMnRE3tW0YLBmy+FukQE8swz
cJU06Xd+7G4BwDEF2KlIecLsUFD3Un9v6C9ITcL328N43vwILdqqmq9RS6AFZQy2
TEj5o3eQc3bdlbmDCWQC2iOyH9yyvdRPIQ5aGNMp6ohiNfDCpQNHwJ7BdWsBYkDQ
sIvGmngDnXmYFCLeyLMwOZlsC4En/j8NzRAx45rAsh7hRtqBYf94WB4YS3HMQGh7
zaXYOIGjCDyLdh8Rl4U6VNGMuaa33m17tnRjHqlB3zmdUQGCE/MKdiEsrB/T6+sE
b7NZkRIkSGwiBMvFOeSBlumyyalIIt2QO2bbGFs8ptjKk9hCEoLp2gogITOCUaIY
pqBkELDxX5t9ubN9Vk3XD+AYZs41jbiH2KQw8K3FZAPzqpj+kTgVReRK4TfJ/6/F
+MIaBd0M+yitifUfoeVlxymWYQ/mK6DvkifKyxl0qS2hkuzu2a2lw9MF9Y8UIJq+
dH5EGyvpgPwz2XOhwJkX/o/38dFmdiCGAS+YxfaR3wKzSVgE+RBFLqC0E3jp7eRZ
sZUcwSsl8/Ngb0AAWInWFBf5n6AlUistoOUyA1rh5rgGHc6xJcfQMH2rpcO2MzOQ
sEHpKC2ZuNStPmdHbvVENhCjSCTjHD5TTQIn63og30OdagxoXBlL03SKwM8TV4pI
pg3QN04U2hC9V+1yf77x53Y8t8KVOGRD+T3gS8w7jE4WE+BQfNu+H3BAkuAYwo/P
7w0/Noq1aLnWqDYONQZovqyJrHU1v+e6bLOtBruu5cGsi0ASKUC8JMWepSMk9DZ7
IYWr7RV2lgCoUGMsNSMHWNw+NX+MIzd/nbuLCtZ75gOQVw/FpZTFpmOYLi/MJTj4
f9Urli/o6UxOqlZ7/+JFvlYPoLUoq36RZEWcGF3H3cetMgQ76SRMAB7qRvHA/PWn
CbC5WjJK0I4S6W/MHKwxOZjjy3Ra2778ngNwg9wduyZp1y4lI7NLw4W/zw5rBJXC
UKdCouN9kSNV8CSGDf9Nl9giE8EiWrL/L0Ud1OSa5suuwc8Nq/q5DrYtUgctWw7u
7DcBjH9SDuqO/jZgLHIIgMyGhOtWbRaa6QYbnceO3ZUhe3kpeELu+J8hk2QEeGYP
hvcqq/GVvG2i3RFmMFVDoQYLGgn0DK+Efpwm0IkwQliu0x6zPwqMRnBqDklIMRiI
ttt6xIEgaOiNsowKaAy0Ad57+a96wa6wYTLj42UBL66HI3inZekYpfBrTGWgiFDg
iSvvtYSGms//QdoFG0noRL3Ez9frqxo0E3az1J4ZOD3lPx2eI9zuupA2cEosy9yp
T7QrDGOttZ904CUTSCHnL/d/BOinTZfLVmBZl2QxH+mKh1sOz4SH32NalTLvTtR+
wA4Wo/0pHIqwxdF2r9C4lWscEGxLu6L/d9E2yt1IQtMtIKzJszxjgnXJs5EPwF3E
dVu2SA1k6rxfSGypwi+8CNIPdv0lH1JeTvAJCmvvRL3PviycSnDtSzowuNYqB+tw
dseTsx49ZAGq/JiK8zQ+LkOirmFri5VwAEewoiNKm7vBxEQiY/ewe7ciF89jw4b9
4RVvRQakdzuV/mxlOzUMsHLfv0vcYkBcxW65fV+xUfosU1HIFihNHKtHuaCmybDk
xU1LULGRBl4fgzyInYTeTUQHsHxuZiH6lRd+iGNPeHCEBnt5tVVdti7lZl1Y0cWP
c/ioLOtIa6YoWOvo2AupctItPuAJ/KCdU/I+2TaR0L8UjSvmafRWUNiY7GH2nluQ
7CmxKVxYHsnETR4kM7C20HzwlMDEtNQ5jRqEaBAFFRm4xQ/BNM+Qe4k8laa53YGX
3moYyYWxgNy5Xdg97xcexM+0O6umdRY2pDztuODjMPmDp1IhAz2+Ej4AZfGpIybn
SQJ5VLSGk1fUGKhT9jZE3FYWvE4MTOegN5Xxx2PDtGOSXhK3uE5italipUgkixV+
2FIM2WKIdAn6PbWBZXwNfa+84rxNAb0iDRWWY9v216ff7pVGtcDzhsJofNB1yJS/
4b7SIlW6gbpVZzsqfMrTZ+3fUQ5ja0u5CY8hNXbmCjJ4vMQxIAvuZzOmcjRWfiAa
0LBWHVJIKK0wLxPbzHnKcTjzloB0Wzh3Z5N6E1XrAKJzX7/VwM9tshhkDpxLDKu7
IdUWm3TuoYHnyfW7KYQiq20KnD0VRDF99IoKo7N2TSumTt6L/gPtGmLBKTECXZxW
cqNVjGtAxPfCRbo21kckYaSuYQF2vzQ/2QYTPSN8ES0BOa5I4FAL0+pH7gwLH6E6
w9YJ8PaPDb5DP9kJWo+lPMWTad1cq0ig+f4rIMfYOWJLvqLTjGIWANGjwZcdzwtM
ayVBUBW62g4F+0AQ7OM7Nk7VA0jZ/8ICNMJXaBL41fCPLpyu2c3cOk+UJsCL0u7u
nvQZsNtnBdDA384okaWHiPFAb2BO+FSjKKIgjRuGumDwVE5ztS4bP0ZPziU5RBSy
NohHedwNtXLS8DYObZOWn2Z/9bBRKST6CC9KvvGp0tBcGb3YLWnZzVuCdOiQ5RBS
8rsmDkJFrlAAaifYjuTbjGNh9S5HvMoeL9Vibyq8RKBY/LNIMNdz/ztFrLSGrN/v
EtKOkQ9P5tqzE/f/u+ATvkBIi6DMoyagi7OqQ51bGq4GQ1dXXqsmL2Z6vyX8Yv8g
1oMugirtkkor558VUqlx5DpsXG521dPSnk4KjbtrbAqMzZkcnLUIjFDJy7eMhyyM
pG1XS4RUH11RbG/VJe/rEgP5G67EdJikjsHjUCSbNGFvL1SLNkvvxn/LOhNfpdOw
uJHvY780jrZO43h7yiv38R/TIEdrtaLYva1OBG1fbFCacQtyRnEkQ1xQsY4pDhrr
mfPXMCs2YmCGs/onsTuHpAPxizOkeAZ1a4az7bpZ5TRT+at/q11ni2gGF+V1w/Bo
K/x0EMtmEVUj2TFb2kHbLCAYWECSP8eoTunb1VtHLzphLODtTR+ifQIRSnP53X5c
cG7O5buhL/Nn0LZYbbAy8HxyaBMjAaGX7hcrte0k4gN2rVor1V9/9NJi4Nf1uafP
gTxbjJWxsPr9l+o0Maglr+g5AUfjgBmmloDTOZhmdtg3hQnvdv/9oSbyadzhz39b
OeKbeHzfttQLOBm3hoxSwOgqZLCiT6p6zI2M2GD1tuR5Mpm2ZABbihc/0NGNXSE1
zBxuW6rQ6PwLxroiB2XcUIGYosKoQJav7OgFOJoSTc6vTV1ohnPRIkaSv8hKi4N7
/F2kVpIZBbDudymt2XOr5BD/EumFR7ri/AujmtG7ldi3u8TTIlxHd1r+y7mjUuLA
iuveZBJngOPnz2siue9xdOVNwaf7eGjGXcan3lnAZouQWYDINT8QiseLVOffiU+3
hhrGUmFwwKiIq+DH++ND+9NRjL3hGiSROO/5e/hBQ27sjOY4TVbQ1ZWeMGuX9lob
WPrsLb3iefMU5CQ8oXQG+h5KmHW3pMz9RsB6RDgtogsqThxhfIKbXzHNGy3QiPeR
osg1yxmrUy+LPfqTInzN36fE/wAQmkcHYBOItjhPFOvfPVI76+w6GgluT3oVzM0x
Yqf2BxWxws+Et77VuJiObyEhwUaOCb7sRVIO0Zy3sucZe9uU3s/TRyailLyOvdnz
ZYWf3s+M5Ya5Vhi711DHGgmPeh09xrtc6yDh0/xeYV90NZaID/4bHG2LTQMiRIHM
H+qVlVp0bUuAHxgel7ZXxn68Fm2NCnFDmcOl/YVNY3mNzQjRgz1P9QuJcb5EgWFq
vxqR1qxPuzTDJ8VLm86kJU58rCSb2DGoSrHkEfW/KUaVEfy0GlGtp/JCrXSBnKUH
8n5uMs+e36potH1RTT3BjzuZDUXnZ4H8PiHpANAdCPLDxOEwfyIu7vAWS/QinOwL
6oPh2Fp1hSFwkQHjHvm3MGyhIUVEoTg2PXuUz8g39bqzb/vPxl0DXILr/aazwbJf
xGAWALaYUMZT5Lz18D5+/p0r4ZQW1ngv+BCOz2IbRLtyBJdRFJCQaZQOK03Bv83C
4JF6GQdrdEtqaJG1ngkfHVS4ysXZ8Qs4ayRvPB74yZcTmiG2+62Q1+orr6D5CAsJ
T2HGjfquw6QD17SFNgwyOPF4PQO/UqkU/p0pq95S0XnuCBmh01JE0gkeDTWVpaKH
RQB7Q6MTsM5WeONTEK8O2Q/nmtHkdWN2NCzpcKOax9PppmFwTBll5dPqlLvEi6BH
3JuF+nBPXfZFkrf6AAihqlIB8+DSu2Dt8ri8AP6sRC40NNsftQAB2kxEz/APzkSV
0zkcstNtWvOsldd1cL3Q90U+/4qrnOpjC0+5PF0DUOlvhm3/LfbQCAeb/dxlxyza
MD/uA0uC0zufNVP+4kXc5wdE9Ct/qB9rRqpEr/uZEi6Ygd7wK6eoZWdtygh5jxNg
f0f5yRAHzviRqQ2t0t4n4M3Lb8RyPbPHOMln8B1+M0eKo/hXA8wPYTuKfhR1kJDk
JB1Xk0u1CAjEDKYSeEVFfSOtI4Pv7afpPedM6zCBiq7/KV7t/Yo2uVDcpSEFc6yF
6NWsxM6uPDJFQZk5N6hX8RIV+rcWwUxyYP4BDMCha7v388MhZNUpSvZsJlvLheLb
ol+YSpRVH5tYcX8fZOUc22NZD+crALWFg+lpQMnPM/PzEI9CKzXE+DkXpuqOO9aV
fsnIZU1wIMfIsB7f8qlX7MdvIrMLNil3jmEzG+DVLmayyz1QkjxIUvGfda5X2O21
wLwVQjI/t3nKsrQ09T10riBjdWMCCKkNlqk0JEJJ8dvjLYpxyxirOtDi+5yYliO1
WapB98fTzdAdKT9R07g107GRwHDphq0A8x7327YtuZZzCUc6SXlw6R+jVZlBizPy
NgsBWtuxqjRmTWkXvysT5SLMA56ZZ0rsmT4Tp+n/MzmynAno+JZOg6VPASHchnFj
qKx/CQqkvwAZNbW/YDzBK2qZ/p8sywCQtrqs7Jp3jthtgLQyLhYbCCPGg85ai9Zq
YsFFRYMONTNrm6+lp94AHWA3/0TeNsoRTR1mOVKlHFs3CtM9fRKH5YIfkj21MZy/
G22gAoEt56FJr4aIvqPCSZeTa3ndSdMU7JG6Juk7QPw9PfqdeKKkIiaVUgob4nNN
zbEdhOh5tmOwgMVEbc6ExNYuW6xTXQ6+lMUObYkKqNkZtqCTSjX19bzU3GOP6man
CPq1sed8OOQz2Epf9BSBOy4I6gpVKvBLoDlqYWTMb9whmta912NI78Tt/uSDOIwy
CAE9BjE8kXYaYNaHwUUr+sVws+z+okQB41lpjXg5z7pG55BtsaZl4TbWFMJsoefk
C9XzXleydZZspYwb87ZXW3vu5MyE01Bd3AyIQJGgjUrUgu98nY74a6eFGFu/qyej
UjsJae5Fma6hOQ+xDlz5MDFzSlAQ6BgYtQbcmH05YynlKA+wxhxehhcbbtSQ4/zM
gi5KLC3tJu9rxKL6AtMwKdWM9PZ8ON3sgiW5hC2PDC5G/bxFD4uYp0KEDUJDDL5P
7AqRhtv4NVrWYxtjAhQXjI70TO4PEFKcGGYIM1ImNw72rRPT2YSHoZMetKGmYSIb
Svf3AuAknZFr7lbbrkOoUndtDqGVVM+FurjNbPV5KRKH+Hj74JmCSZAbZpFXsC/7
+l+k0zq/qy/OdwVlO2j8g6IQvh4EtEO94qmmMifpFUMNAO7CwKERd6rqswRwkIiw
SleypLgdzAXi2LjoUkVulQXVzt3IKio9I0e5/KqG5RlCDYfQOb9lqPbz5Bwxt5qy
DIQP8VVxol818JqbpI8HGKHJPEjewRcfd5mAqP/jPX/CWhvaX11K+VmEwO9CZM/I
7Mm2RSEnWaqSKa9eHz4uFD8lIX13ZN8712QfslUtXriwBXvqDPXGywpQX4lfyKoO
1+7U+Pf08UK71hJ9KMq1WkYDO3tq95jdBrqjwDHsVsdLzkSWYS0cNZ7YUKQH2QqF
8tovlnR3FfJlp+sWJA82yG4TgI5ZJZimMzNV6IIYEtSqCUD7Wf2nUbAW3hOOycp5
ThRxmqaRPOXEvGgPfkNuWMfTiEuSDkozJjvUTYfInumwHURyekRIzny38jcxepcQ
sScYHQg7toHtlAkeWDvctzHsOFvLjlBntl+hR/2RKZINxXCHCdSJKfFoQ/H11/FR
nlfjWCHvzcp0dOxLUUSpP8NYDC1IXaLqwwJHYGCxa8pymmqYgGNknRKQIUhmA3BG
ELE8TA2NMTyoKaYDqpVYMC4HkIZqo6qJkJWEikKXxksYFe6tNuEHCeE84uAllSPV
yZ+Y6Fta5hJ2gpXct/7QMkjuMbTcB24zKXRgi4yINnqnTC0YSdFBAZ6uWeYQ0VY0
SjNyhE3lemiL8pxEcGsd37bV1D5BP4Dpx9izvX0mpXs/yAznrcJaTF2vfKbRlUOS
Mqa8UMGdvOJN2AH1GPPWwDXNgybxIIs9/aEL7nlyGksF5x3TlS+2ub7gpywY+iPN
Q+KfZQ3gVU8A6VDxUzYF/7et6PrM/UPYUn656MCH1iAz2Fw7SGw2x7I95LcAXr4K
W4pa/zei4ylprgWTYJV/MIyO9T5Sw4TX0ZG4rW1yU8xk3hDprTtQ4pyUMWkIT40e
KUMv2Mi4IqG7HEMmb0bE5KXVIf9zSl9+f/8Edi/KnAComeMnFKhp1TbSvMgki+Fe
oyF5lNYEnTLv9rvhnusVLgaaKX/E4bQ4tZkWtI14dwlQugZr3AHWpDrOWJWMVK07
h8aOLEZil6DyMBZEvEVGzoHQo5FxjbrNpMtwmpZzHZAVoRoHLVvJWZjd6mGKksYa
vnFjbKdp8YGvc8LHFWS5H1FnCCPRe7MNJ3eS6ljoPPNLXx/QyMins93st2NBz76l
CJphCdtwvyRPMOnP9eJS2+40Hulp9MputhDbZb3AuOyZcSOK8GHO6UY0GpUNjFu0
O0vSFHKVBo6xKBwps3aLZ7SLtHSHHjoGYBGykZ+uP8jn5ud87fFMGGMIUot+tn56
+euJOT0Tazu7zwNk6RNRTwL0kbgLK4n5SXLc1N9K9w1rr4IJeyTy4xGPsrjuhVzo
wmcIUN9krL74YnHXYYlLC9YUfTyaBakEPndLJisSA2/Mcm87tQVqF7MejDOcfBza
8afAXBAsBlmgfqUCX9HAAL9rWH/F6HFUwzS4qugShEcDxnSgsck/av0vg5ys+S3u
Pw9Dq95KqfbhUWa/98il6PBp048AE+zjVfNU+dD0KkvFSpPQZelkROJ4vX/vIReN
DpO9pSvlsFQH0F/dscTIx/qz6ZGTO9aLeZzyL7ka1epam9RPUfGQxHG0KKrJH0Jz
4HnE1ZE486wqCgFaMhDFmJZSgbJ2mciaHyVgotURXCNCTLIzoD0EmFCEW70TXZym
AF74v2EGY5yqyK5EpMYzEVn5r9ysXBOSdcgCpxViYoST7roR3R0iINo88iu+CNNc
P68T9+ZQlbFxL9IVF/dj4IaWnCwqkTxEQXBHw73/mlkqco7S+CWY8z2LrcRjt8Jw
xWahNVPTg0kukIEGVLc1lE7dsX7JO6dkRTzoBDfDUuYXfkj9tFzzYXx7NOeU8Z4L
ajXb/k0ka9/tZe6UnnngJMOQcz8FVaCd6nYynBKHbt1geCytPtvUbvCS6DOq+/WW
GCLurzDZFMu3EAC2Jt6lv2iGTnAl8OIE0gIibKLLcVla3/YIKMu95/Te8lOBOYff
zl8g0GFfpAQVkfY6wjJdXaFTehxVt89PNoLDl4oUpP9QBkGmLmTxN2Wo6YNAUr/H
gay+uRA9elZ2xXyJ8GsT4SlyQZr7rfpMfXmj+XuA1wCmhoZJYIVurA3GulzuQfPY
ITaJWnnbXWY4JPoosqh74wjP32htk4RZ20X6Mn2r8JYkppy0s5KPB8MEo6MT+cPL
lwhkFQAKYrCl+APjbbnZmtv4yU723FnIxPwJeetNydThdqvY9irNpBdjyccpiIal
yS4HSwtmaCcKr+MF+bIOA5vxZ04SmhBI5ImhQX0+oUmWdUUjgFkgb3yvUmgiiQKu
Zxw+xOsEGIPZKtUsiNjwT81CkRdpHSbx/GPVACfrFHBTvkuOFkkzhuKmNnn6iVwj
3/c9YoJsvkon1f16WKY2JWga62N2eyCF7ZphEXopOu8r4+sM9nksttIgTcg9lwAD
5928DwAm7dlH2FzYB7MbhI+MrZxz2IMp+OLiM/vWCtyneO/4HM9dAKF/5udYbh9m
eOTnxndoTVD3piQAFjiX4LqnL7loSnjVznFtr4TJiYNs88zOG2N75PHnIBc3urRY
j5pTcJALFKAvivIrVehOEW56kLqaAHBAZ+PLLOQhD1WlNosRSezdIic04HdtZ18I
T/r+pCmeOw5qvQ/d7k+veDljgL1C5COvpU+ZHwM0JEMBSksjgTDMN0WVz9t/9zkm
uS6kktjrgpe3/rFgXWuWA9jF1KAGuinuDC7cL7qNUr2fGCHdCLgTrbBly06DoyNM
Gkg2qnF8s2bFXluNaEf3YqQdJYex7K5gN6rQh6nHBGhZYNoKiNYkWnvrn8Ec+KOD
BBq4A1KhGibD/NZz4Y2OvQ0ojInYf0uuJD/K79qdfChzQlk/WCTcPor1E6N84Goj
CX1OdrswNBYFchByS/pYk5/cHnMFYRAZM2TOJniWGYYkMZCJK/xFk8H7C/ozbEjl
oNapC56O22RmDGGvm7VKOIopR3/HmfHtm0qpsH91dDFos95pbCVOfrLywxkVktTy
nxRTaTuZw3cn/DZ3I25tFshc84NyFaEC+HkHUD3of09gJ1A/aTMBSuifqar1s6Oh
9W/71BIOxP0yGsmcym96S0iongHauwUhhCXIwS3PmLTQ3Dob3lXiBVHXFGjFUaK/
4/PGDUNbkadavT5YJvKkF9rndFV8mnnRU77TLCELsZM3Gzqt6cHZruAEnPmq4zdK
wKla4QxIseSGCZLC8j31rqOoHU7wJ23bX7DML6I1UCLtSm7xAFhbS+ZwlwZ+96BP
84xPgbCrb1XW82K1tJ+OTbmEgdiZn3w1tctf/TTDhgMI5txIoNurRfESRR6lgyFf
3EumHqyd6p1k9//Z0hiIT/0ziRfejezHh3Lg4m/VPTn5iKwe4sjA2jVgZ46Ovr6Y
ERGtdASPr7V6AqPgDOXHc3EUjUzQ09Nb04/QBLzIJ0zBF9DZObixd4QyDPRkC4wl
ij8ZSxMMWhrGS6pJQ5nAFwiIcvMh63JejbNoauK84CUpmEJKAT2e0Cp/DSQYIoTM
r5Vs8Xt2Vs3QcF1yknisCHQKUgwDnKh58KmVJ5busi+S33MlhzWR/Agyedr/C6p+
3GPyGtDB7hoZG9CEIRO8nQCU3wT05gfCMVM/FFq7o1fge+Gjy4YFixED5H4fdOSj
CjVMQ9VqoBwDF5CxueUGV5/UN+Okhch8JXtREJK1bmMUiZNTPzLSaXgagJrF2AoB
qwAMsq3Bp1+fV+CYamHEt+H70TbDsxbZmaAjOt6AWZ3kRDejsBRlWMXLx0d+at34
wLQ3tf3W+0fqJ+SBWCb7xQgzR1A/Wax9fwk79/BsJcEFZ2rA/cTWkfxEvgC5CQzX
O75g7ChfuCQGO8BF8+Nw10XA6V79iI0I2sy+amjtM2UlgVZ1fVaDogeLKnLFZZ9u
t72XRPU9QSI03ty/eZEnsTwEJlUuVtSRZ8bajRZIWTXw9FNPu5IYbqbUXGOAp7LZ
mZH3c7pF55uXyxy1D7d1NVHqCPajsdWeP5PBiSZs9nQ/taHjlf2sTnehDEii/i0s
UxQspnj75fcWoUqrQLUVKsZqosEmkOuJFCC+Sjlp/ddcPr7UIqpM6g//H4Sx7Tl/
DXn2ce25rNSF/rGD7kM+8GoKlwPmWgR0ZCnNvsZxfq+2QRpFPoPlZPQ6BV74HWpv
woVsDTd+cocI23QBUReKEhypkqhpVEdZAHCZso/rjQGJP0oecmH9R1iXMzRrAhJJ
tiotgnTfGcoE7+B3H/EhZ5eheomjliwieZYMbc9rDkselvRUX7alIEaPsa2vydDk
MEVX7ApnAvxwyPV4MHPXgU7fRUQuUz8QryHJQysIN/e2z+KZfU+2o8ZjameUzhMF
4xXDLx240NmsdCTPRmsWIKnVjUsmLdIPkJMthdoMfIXH/zzdgp+CEPdm2qz9+iRZ
jMuHFm+yYYVpcEzNsVuq26ikZ9mvxVJfHucxaak/katoUqaK4uAkkdSvBb+AlnDp
j2+KPB+Fe5KmvUgwPbgpT2ZUzCL1ujc0sd6BMIi0V8lwFg2FeCFYbt1ErIlzYilj
P936qnQP6ioz+XaCMvm7WzVCIHr4SbYv8HtdLrveiseLmNNDOkkos9TzKWyaYOoR
23XNJG+d9QQcZqYq/gMZThkr/6R1HzI3yU+Q5tio0mc6oRclulkSQ+sbafaGjmyO
bpa+YdavpsMtW+Lb6d3dtMDMRW25wsvTdm/7zJBg8xrzG4ss+ABFec0/JFFUaQ68
/yOj0kDVmrHo4c2NJt8U4/wOqejDD0bMejNXBWAK4nhrDjz9grTkluq17GvF4ArY
ct9w2xU8XlxkzfvdupNKkoqxtz6kygG2adS4L7L1DLpkqQREfmF7u2f2Ljv2mOYR
NICEymApcBHUeMbkKzqMV4ToCkfUsuGbMsiif67eHRe/AGrw+JDpBDExxgB+4dq3
uklVmxAAxGH3cLY8j+m57lIhzLjWF7fZNaUY1utD51Zg3iwMueax3JbyZtnXQybZ
3OqziQJlhMq6YdrCmTeSnx4BqBUzX7vIARP+IJKrbeCyhLGxrdENB36FKKqDd85M
Zy+3cGsMm833+ekgS3O5mfUlQJNKyvWTmWOyrQEStgH3Lu5HLXdTB+TpTSOEFOUm
wn66/MZoy4/bDQT/rWSZxIHkCTGMOTP98jP/ROBKpbSqPcAj5bFz7GtbCCzprUUn
98pV/Sw6XFMOSwcOMR7oMSJD017/3e684noDudDM5/kDcfVRmqXb8LBvz6QHamf2
sq03q9iDa/Trcas6xO4gJGr2CRkKmEmkG2pXYCr1c9AbpqxNTQh8NMSuSWnKSkj9
O1DHTxBjpeBnxYiwd0fqYr9/ikzIL3P/upok76elhPHrHct9aTlTi4fd3lc0N7ej
ilIdwngLluJmX1xs+Or+2veCmRtubTVrQ9gSkdvKDagbpQsVsR/ihy6qm29hzQ3h
ACpKaXTlM6B9oxc8KC36JB2Wt0zB+Kgb5EnMzcJPbE5a2KikSEgmo0SKvm36He5m
3qmjFUV+HuqqJ+btZc9IFuLyHh1fScn03s2/WAf0o1TaYk0MtIrS/BkkWR3XcU2/
eVhJVLjqxZTi11q6Th7wKFol789+wSAwhD4muhnuG5wrbDzSUCDxaQv18qe8h++J
THAJROeUIxs+rTp2Plm2eLljB/b07VOHHt+An9aZNIEds0gtCGufKJAWdo9Xgltk
U7E/iUbIHuSjHIomFxVowCtdyFS3N/NkeuugyzvIlPXLiE51669MqRgWrP0NzC3B
6lKnmX9mGHdSooEoTyCnFzRcOdnOdAQawOkxsHtAIsFmME+EOm8KGEynj4pWoRof
L16uYg9lOAGYckAd/3LBPINsCwQn6x5kirngUDEkXJLGGC8MSL3Id+UDYtmdCKFD
JotfhlRNA9+SwXlia0+8sPQfmfY4/t1RGdn8RaQ7o7T7peIxVRCz1E4liHidQ0oX
FPLjnETv0GehmmkgCat0FV9NfR1G1cgUYh/iV1eu3nYs38H3hb0S5EZ2LaKB9RxL
oc4m6LbeU6likaNrgAUIYBIWKt9dLC4TM5UtTJu9oH2PYVSo4sUKw8VwiQWcESQp
v8ZSxh9IuAgAVklH8HJy5iFpfomVnWqSJiHrajtBO7jj9u1yK1Q0SycchN42w9pT
RZAYZNTe6k/5KsbkHVkYWy0VlJloI11Rj/dqeN+t5OCivmYqd4Oe1kT/uTQdA1Y5
MXsg2CIdz0Wb74iGujdI1/WEeXRueohfwcUzhfdwpk/MSjuvnEGJukQ4XMDQrFwq
jFeYgZVEV1R+KjgvQ0Gp6dVdUZl3LFwTWSZiCho5i/TZCoqbuPL/WL05LKm5CvBT
Co823Cjw+rBPreTOjjgcVX6z0j9uNVub19FGkwklpGRjYsj9E4NWA88RgtCzzcs8
Q7+qwqa++D3aIJ5prfqwgURY90zlQZLPQlggivf1fOLqeXIQxIDZD/YUNuf4x+L3
IoPD/fvo3BL+K+nUcKXG/ho/s4m2HBPt+KtWCZcDWlSrRjp+0wY64Tgri2QLvBMD
iCagZxkB7XUMEUCC8B73cNX2R9vc3apiQ8lHQfNmqW19eqoh919p5zNvDqsxDqrH
flYFYVP6Rl4NL3m4Al39zir7sRxGcuosfrXmelue4VE0QRkpOyntc5VejyulK0cl
tA0TEyyCXCBXh0FUxP1ApX6lNV8rUJIhFBAlp4ChkXUD8WFTplxAaFzkFnR653Gv
OqF/1KfoabDYyvrkaVpIHzKP8y6193a/vnkFwa+ofLb4QwRzgVPkJrFpbYw14KZL
+0+Di1qHB+t9kx75N+Nq+FdJBn1jDyRB4sSc5Ls6+JmIo72F7cBM+HXLQ7TZrbfM
TQHgID6YP8okJKq3xYZ3sGS08khfPVZ2ojMznHmn7CG06vGPgrHyp47B2Jdf4VI+
ymFRnEW4OVB8DZfMRkYEDXworbJFfpMEHfl1HX4Ovildy9l2S3X4+72ffQ35hW/j
LlvsGMDuqhQAfW3DRVwtMoEIqN2bUzw3LtzG6niQJvtFpOlDJ9zimquK+6tN8Iya
Tfaen51siZP7WJe60Fih9BQnKolHbJJmV96UNEz1/RHB1DVpBVhXHwV5Xpv0kRbo
cr6vuw/N+XI8h29ywiRYZJKw8tY7hT8grgOZOFrA7q+JCMWy0KiAnyVB+t0BWwH7
CCHJCIgIM9iivLZHcXSabiAwFugUadfISiGh2WFSsfbJQ8wfkTp0OwM1mfMjMls8
zb0AeMdFzgtOlDdnYZjSoJOq1LhdBVBMKCCoULfLzdOhvAQt4QrD+gUMV2tDPYSI
bTu85gVULgR1wk7byHj/09Yf23MIW1dk5NLIdL6ETHP+hzXxvJZgeLcBwrj6x0JZ
Rikah+WrV6rF+dG+YBAkomKtxQkhywmQLdIHcBblyFKgjGPygFKmc/Y+fOEXI65P
x4sFO0Mp0BIRR/IBnk/1C9XmYst2mGjXIh4Wp+PRSyOiITer2PFDBIJ57/nTEbJ7
p5D4AcPA2QIjZhaaFGn8yEZtLg/MsRCOBdV3/xffmPRpeQ6d4WgJeqQ6qiyk5EYY
2nh5j/WnwEGt/lWmQCaI3jSCBnWqUQTEwCrXL0KwTvIh3quMA/DZrkqhR9JZBYSm
E3cJaHiUfjeblRxvQKhioSdwBeey8sY2f8YQvZXJBugmbdNAik9oONCHOMtRiPVy
68XEGMbCxaF1/IqCTDOZygf/823G+CrJHZHgHdlwGsIcGVOkLGuhcnII4qVSg/bF
nlimrz7JLN62tk0C1swoBBzdkv/qVZt38H9cMvv95PmykQm58Rll3f7p49bJQyKF
jrPzM9SbKhoR2Sim3NM7TdgxVWNp5R6WaVfywr4VWNrAIyeUfvzX301qk6xbm+/a
Q3P3nux1a6JnzU6sIuEkWj7lHI/ns0rd16ADz6ki/PHl0DQafjQXMuVZDdooEf4c
cK8wfBIgTsKZmeMsfalqI3qjqJFzwD+gkC1yaZGQGbTGutrMYvNP/GAazNApy+hO
MFk4DNY2vege2bTiQ40svvEhQY0w24Onx2pb9txRWjE4QzMhrvtNMutRkifI6Lll
rPsaRf2MlWNOHWHyMUHw0UV6866AtgM6PiWfwSBgpxs5M7oVOQTtMUkuFBy/JWos
Mx/ZXZY6wnwq/U0qUjhyMPd3vccgejEFV/Hcu7ItSqcRgE8Ps0lXNpxyCkgAdMVA
Xz/+UCRG0Zfn7xGogxTARvY4t6rrasnUSHbr+035XJtYjxX8vHcgNC11z31rgmcM
odq3V1LSa7zVx2HAPZFQ7gZ6d3uuItnZj/irSS/M8JmUNsRcC45cSzQG5Bl3/XVe
EyFvcClBthmcEycYrwaf6riY6FljjCYP4OGWVlJjX7/cMgoWJp6Q/jjQ/tiHw5Jv
fYwxot7PVzBsF3ovwJcHwARS+4f1deOE+gUlgoeE0Z6/Lg4DKL5OnPaPe3fer00B
AOFm0FKhlDfX1d8sP7+VtjW5sqECfH5PbRJsGupGfKRs0faNGXeIwMz3V+V3OvDW
OV6H8O7BR0KcGMwQCw3bQSENFrcx90Y95thvNo/w0tEkQ5G+Q9vp8+hu2mIkUYf0
0ztRH8MV0rzX5VUR7Hmq1DU03lwV4E5iXiN36VK6CAhnDfdzNL7pn9CeJFy38UCv
a3xehizdCWsJVd89H1biR73PASZUi1Ngwmd00xybWJkdsL7/UmBLVm9sFkASct0h
HWBHhYmrlUQb3wMzOuHIA/TTpFn2lQyBSNU/KVR3sZGuhdU0MbWqpKtiMs7HrBAD
qNIv5SM4Q/KQiu3+TpyNEd0dGHsseMIY/wl00sQU1YglRyUEjCriIuxCGpwAyFt9
oH6ZcFI0VEjf2VtCOwqwJX258URlsTzpPn6BSmAsaZd50dRmo4qCz0r6SXagWxuV
H3Ya6MMIbG39HzmjSTKATGWqts8qpaQeDGlsLIs2NuJstWD6f7mXEK62iHG5VdCk
uV/Stt3TG6+7OADPeDgCpstfJXXCUElH7k7pi+/Jbpm64A1h+52I00Z1kIV1IwhG
ZO5qiiR6/x49wgyoFCimaSS5Xiq+cTCk4To/LIshGa2hUiXYEpGw/mr2UuTcqwIo
+fW5HMuxO8Eq2VKOyxzmRlWEDeYVbysvLTt0kGShphHra/xD2G0Eh9CoQbodSePz
LLqagvjp3kH0Tal7r8UWUDaYxAgBAE7I+bHBwwKOeXXnuu/UTNZMYYA7VFVtu6ae
zG3jTq74MLOttIKzYbKb+LTAMTogX1qdxYxzkZQo/30h08lixzBPJ/tA8Nu3CJQC
fVY4DzusUM+VL1yjEnAneDZVaoto9xO/AKW2rFXdIrzRKupNNGvMQqYmmR5xn1IM
OEhv0Q6l5Uw5UL9IS0IpckeAFp4uBxDyqRBSZ/SkgmhHqEElMbOb7XYVIENqL0LC
mKBD7L1vR82Wr9n+OrI/unrItDb1KPLfByEWhiX3Mb1jrVTNjquD3TVBOIWhInva
wGYsyNwwkHWn1uV18aZSzr1tqLo2GAqUMqzFH7ZEEQqphh3d8BN1zeWTmpKD4N9C
O9nE+Uq9Y/JBmzPHE0jxNdal/K68xLry3THafUZhKL4cVW4HyPe0rA9W2uutmGMQ
XrzuiaWU/7ry3FIfIgMXNpJ9Mu8mZOWjQfEPQO5QEYYB2eJvuaOjC+TKS9S1g2G9
JsJgE54xAECckTV9itlXiIaijAz/Dh0vC1encS82rET3unX5ifs2FJIhxJ+1OYfG
zAiYRhJ/bdoBOp2RGbuSHbGIEnNT607kLjdWIJmSo5nP8ZpYEMQhLaYQMqLNjXw4
pe76E5hwLHgpwuj6CMXIgkfpg9y+W6EeFBtwgDEGZrqkojGPWaylVV5z9oEWGtun
ghZzJCMzSbXQNCT1hVhivoG06khSiUhjYSPAdpW4wKmG4V+InJiJTWeGECMi3rCC
wQfSSf/TsrJZQXWPfbzotcXL9a4Xy91bRDW5MzQ/gm1mvVYUkC1bwO10oHE6gNSa
8yOJl0pSn6LqKzT6M5ziKaAJDqfvtJVE95DXEvRdi/5H+8We5PC+9H+ImMQIumG0
cupvyR3P/gonQCGBLtm7+3H/NJ2a9Wz8240ZIdJeXVvlmxuNEBHav9JBEKICixWY
PWTmBAv4IqS2h6QrFVQ/r9CWXqXmj70mUb/KNe0OasqH7ECQzb6B3Q1YQjZFaLN0
FNNWbhR4j0/W8SO58GBaEOSiaPYmch28WrsAdE1tdPEo/cKmVjtH1D2LNExUz+hu
2sCAoQSexq/Xxi39Hu7iW0AqcS/SapNLvCSwXnGoS2/2wZgSJN1UK6GVESj4Nsln
L8WGtaJRhx+Ip8duHVA9YeZTyeSdo+lh2kPhU4b5x9nSx9xDz8VYYOmmM4sORytS
OQEoH7cv9WVT4ulOfdxnCC/S4g2AiWnHrFm6iv6gQ44NcnuiNb4OMwMNdq5t6xLx
n6dV9PtiC2nPse+X22+kb5CnBlOCl75UqZTJTwlqUxtMbn6+e45vFVZFdfkiiNqN
1Oc2rGfNBr4KxJcyP/CkPTxLzYRue3n11VSwflA60vTlGePnCpScaZX6kVvxhJ7H
Nqp0G2UEdHn/1yM79NYtVz4rAf5gQAAvToW7CWBx+D/epnTkWNeoLx7amx19gu6/
VxWlgUyrlWAFbKQwZOH40FwcDoNwzCO0PBapTnBXaJqJVUAfhgc/kIsXARlUiivT
BZzQcP+/AjWvtqJ6KjWW+CeI2l4BcPnsjUBT0Xw4RpDczm9ZFDu+GyC17mpBsQ7/
2y4JfX2eGnuzBhkmf1FU1p2ELBxD+P4SBbWmRdNVU68vlv0y7Cmkm+61OXKBo5+0
cL+zPgMBe53vWzr+91UHRGFRfpMzrPBUavlMMqSoT7ygVuhX7tMBM9CgqlimCFdD
MmIqAhVDDuUkCs3p71XjLlaN7eXST3XEpB/0OtXpChpI4qZYX/UbEwzUmjN8/80l
HOprS2tOpOZcYNlM7wwAQhG4VLkBJnygc0fcRHh9ex/JyXAfFEoxmQ0kgBYayK89
a24upyt8y4doGXOrsgfH+o+ApmqPSQqff0kZDOksSIkx+5H2uZoaRLwBF4pxO10T
kOvK3KNxlsmPcvend7z4/AfsIqnkEwS+3UE+duS5GXABUYjetlpanpvs84RWdMRv
UfJpq7ZJcrxGHtcz00TUQOYOq2LbawLHOTIKDkkeMZnEgzbTaLgzvYchmrF0Abww
3EetS/xAE73jSUOUBjPhHbw9AcjhRL5Aofx2VbNLl1N2C5ihkMmFWGoRI0rLCPVb
NqugFLe4TOfNVF28viTsCYqCLz90+KQx13i4WlzYzvQNV5UTzUeQ9MHp1WToVxVE
glJGIaEVnaWH3dm6nzonapPFYD/Yjnxhg+ZrK/ZQ1XcJfvytZHBjhAljJhIgW6fY
x/+UId4YYoHCGqwE8PD1eBjLouGpQcmJNrRQecv7MUm/zMFcd5pgTq8Cfje77dHW
5aQexmOZ8iue7DBcTSf373XL4AhKWY+iyqK3WPe6NOEGFNhxy6b23oldtUb/zo70
0kAQ3x5RdohUaSZCNhAaGhaOh9BoqQWW4xsAAo1dozMWQ26u3CPRMdg8415nDIzD
RVhmu4x5B32IGQ20OYmLMoccEBb0JMC0jn4wTCB/CVxnWzLkBts3LSxanE9dgiT6
YUkf+ymm1HRQ+XUZc7q/p7U6ZIGx7ulI1J+14KlWnwxIQ6rndxk6Tzr0QVaxmnCH
IX/rY2/fvmBJNwyS560/t6XN+Pf0sw4yClfCeMllmDASDogfWgxpUTXAsMOk7HdH
CMzFu+bZjL32E7EVtSr1yITQGca/z18cqvawM/imsf649RtoAzbNV11zQW6O0asM
62JIyDTp0iiiTSKauKdXtx1/0HQ9zgIwvNLq+GGP8sZS0Iu8b/hkQ8DivaNjGXb4
T2+J72xbecX4B0tlDlyZh2SOno/D8e7zrTCxmMMaevzb12MAVzwcx3jo5dsGspGl
2IYBnZMSgqD8dM7zTmCCe6TZ/7MfJu/D8z2fz7nDSvUJJaV1Tw1cDBNhHbgSA3f1
Biis0MM9tQaEcVjQa6B0Z6mpygLH+JAgPF3wegTEAKYF+kdTBJyX1ZpzcWnO7GmE
kBqk9IWiV/VGB2AeJLs047eCeV2RB/10WEivMzMMrkq75YRh37jyEA07JYtJrC18
gAXiXlHw8GW/ojl/D8/gXTDEAV/KyPGzv7z4VZ0JPG3QZICg4K/cxpxPmNP6Ctko
GGx80yweZJ+WWZI2xMtjv8RKQSRhOeWv39JZE/e8QuE3QvskyGVWazzZRZAZxE65
zeFMzLV/X5zIFBYwf3SAwY4uSeBM+P22TOZiwchEdwdNN1r+BMV+5yX3wlwbv5Z9
Pr82o9lSUyb58u/mE5J+i0x5f12twM7UcgjcxkPIjsBGOX34gXe7Gd682zHO3DtW
dzyIGyaDkDiCdrfyoePG0HXXN+vi8A1roa017MkNmOn8EqgpMTZUb4bVWoO9sVBR
QynQiWOPaI+/qJjUAw6JV3XCRQOPdbtT6G3OtEUYDBq1DS3Sg/uKwoGScCLQN5bL
pC0XNTNGuW4zjicPa8L92N4L/Lcbdb2yGdM/phHRUBY+Mkmrpe6sAevxY7QKps6x
HHiRFSMAQmrdSZFPNAxtjQ+zHDImpvPhxYJwlF/ogOTT/oE8NtwS/5I2dSS1JbkG
2ivN4OPbe5pMtKYn29R29dld2GSdHCgSGlYuwYrpdzpLW/VGL8yU5kl5QSgYi88X
Nobz4dKzf9l5ZUluZpNqwQtHH5yuTY5Hxj77wU7jWMFZxYBsMEsrIRKYTCRa8s1I
/ARQVcQjk5HpFuV3wk9lLODdYz/iWgn1O80NsVihy5Zvuz5BNy0FlBQbcGrSqa5e
jnKx0kiLIXDt3nNFVM6fV071xTAu/84jBxwEQ68HyQhWN8L5ty/XNr8btP7CNBSN
5FnKsdzT2Xalnpet4SfZvwRnaXe0jeMln1E1C9zihdRCv1vyNCim+XVEoF2wok7+
N5I2HhgXb5EKkskjv8uA2Aomvc4jtNl3GnDMR/ZZisOpMwlSLSJ9K27dDwTegvHx
OCAz6shWm85jk48bH+45Tya0c7McDoxtNcgUb477Y85dvALmapjMXhyfPrXJf2Sd
Wx8subNY8qE3oyJMLv1UYdtFOSOubadcqzSfl66l5+g8KQTi43jrd3L04PVqsfRq
JaF0oR30xd8zmQl+UzXRxdGZz00jqyV4IX98q3aobrooPAKz2yxmKunNUv1b6zwo
jMDI2IggSiCVIeC6jXo2mtXnYsbXlUin/b35lomGVbVxP+1UpUZ4EGjIWwel2YRY
dXVEac3LKDbZjXftQbUiEMectOT6FoAkySo4rnZNYXGEPNaLoTWodNIe4fYqqPN8
TiIawaPOz5qaDPoJElqScswqYX68U3lJ0xNOhzDjPDHDnikGmD0x7EVc2bYS4BPK
Bhp8LgMNdaI1323FcSpViIZ59PBLANwlzMVnf+jKrNXwqvynWVXt1VIt+FXjzqBl
vwJWdI4fMWhqVmBPSpnwt02kkPNo8ltItDwrDNxw84d40IRlXhNs9dW+Wlro7cLF
wJo65J+7wsPqrhMmn6kFNNNsYzGoR39rwYgITLX3nimLlqO1+w1B8DllGqv1ngBQ
zsRWXyzYEJNnHcdolLZJdN1gDPR1SacjPdxIUkwZAFyBt7zoszL8q03qB3DCBtPC
kU7bas8YBBqafdt2TWj2Wcl3DclUz6HHdq0IbZHQxDFrwyPDYW04b3YZrJVoSvjO
wiGfmMzGCrQf8spBpb7r8JqMMXpy5/AF9X0zKgDl7zlU+WHNttU5j5VP840DYi2U
yY6XazPHr1eNAIwuVx+Dtn1SmVArvwflssEJURSjqjNQeDkVGcTuALjR2UV+Em3U
G+dwNv4mFj6GqRpFSkgQ27s43ptGQDCsxaC1O31BWORiFQr68YnWkFFQXdBbjSF6
WtVvKBpqeCcpQ/8ftEW9ybvDX1ALB6PmPPBxOJcem3c5izYQZogiQAtNxFpe0muG
QqljNnsBFQUSyIpkzKp4oT978ot0PGlToXypuAZdnhoxH4de9MTBonS/mnZDElGS
1IeJtzowRFPgT2jiD6iDNscLrXcFLoSL9mkxi8cnbMwkGB8kMftZVpWIWkJRe6j/
H5hktqBSniQayOnXR+OHVoDUWoolL2fJfj9lvgvKnFw67qK7eLuwg9C0QBdKtGDf
m9KCxYi9PEXui3MFUizfh2Ls1/Ct94tbTnc4hLQyvvp4ElLzBYgDOYH/SJsZyJqv
2q4WZyTG6AdQVJg6oV/Pg8C4tVMwV7IFOrfmLQZXXAhmGRLctmTH5r4dr78OGfy2
UhDarDUG8hhzD2DK137J1Gi/dPqV48RreZaztjIe7m/53fAkDuvSo4cHIXhXWBAd
qHGQ9dwm4v+UvjaFO0Uv12QyanGiTUKoxhwdayBUEAG1HFt4Lhr+Bd1po759/J5v
/6zbp9GXlEmyeQNIzMREAm6f5SjhjVIOG6AVcRQM04VAxYeJu8mSWOltSmdHWpuX
TvHwECycNZYZ+aSWdPMxTzY2lQpFKAvIegq8fxy1EMGAmeJ50KyKPrgpUgvPs+Sz
oHYLF8YMYw2PRgTnBAV9iohYRUrLSSK3l9gA9FQbxbvJxFVnwewMDFNry0zF0lxj
I+A8Wnmbsa3dWLEl+exGugWMap0HNHNHkWwopFeEezm/wpEPUzP7vGMVDgoXQgVP
2e1rGMUONvnGS+OnbuULD5d55BronfEORIpo1DDHoA3m2NzqPsYcGho6q7vvm9Ym
53BL9+wTTtFFyR01lxPRzIp1RuWvZD8Mq1ctzGxQIEhNQCrekCn4Ar4i/CEf5SQD
X0nAMuC4jBsQQeD7M0WGwd6vAfWFsyYUDnR43zYQw/g1CNHfmJn/slPnAMdqlpCA
Ifsf5JH+UESmqmIQMbxMkxsZd7D0JRO0fIOPYAIvKWaP/oUE9xzGcNj8lpWM+jEb
cKWAq4TVqQ6Y1on4TgtFfmF0RfabHQ1inERnIe3gaup1xWt894Iw3tARAJJCGTNy
MQW7rT5YVMrGtx7owip8hHY/SN7SlhWhmf3Hd2qDaSYFeGC7l1O/uhAdGoCmCubA
wnf/Y52GvtyZp0oRylD8EWaNNDr1+b4z1AQB2QGHEHvgebSZI6/q1CJSh5UvexyR
IZvE9eZIjNBJRpAwXvXMhbLQ3OOgrZuq2gUxqngsNAnJl7xFo1gjiVQPmvOHk/QJ
BTxFO80aRJykMXy2TIHiZDF8k6Ryqjl1UnKT8WmPumMQPg0cmI8AillN9UmIDv/u
BdiP8I8e1bOCXTHQt++QvxTuDO87tKoL6QAo73i1YEsaHfabIgJpHsQ455os7DpR
rU3qUZVs4HR/Y5vJNqlFrOzFwyJI9yH7CvuOQhDFIVNAhYDsaY1XYaXK0pTsEGUm
yHJ44GKaPQlEPI6auFSUnSxaggpJ1+zTBeTZk6hPr0gE96JZeRTmfD1WtyDU67og
w7EfsN7w+f5pevAaCkPuOV8kRV2FbCQs193TZuKQ+KmY9NW4M3Ka/KlnNjFGjYbn
NhPheNpCRrwB37EM2hjJvTL17MLSdb/MmNuUsPXEQ56P3RdryuUEa2oKCoJGRffx
S/RB/0OqSgGpQDC7pD6L/nWbfQPeRsi9QyEHEfueXYurI9yT6xklCtOGgyBZWLtH
U1Akdd0jfmxVTa2rlZbteZDAj5BgU6dlojRNGpE0gpuy0/wYjf7HvXQT8hmL4Ddq
bPuTH6Ducr6oMHtrWZ68K7zlCx/Q2lI20FcaAV620H2mYfNoc4HF5dMzfWuRdhRt
MS4PE6ygVuQ8t5DEVzh/0lZMdcaIh30KXHiUqrhyO0AITzIDEFaOasrLMvyAoGnZ
TQwdx9FdngooE2mCOAGAl/LgINaFRPF/P0sUK5VHJ45ISYIkTqEPckdeqN5/MsZW
YxmGPN1aqQAAMPmESoST5x02ugxaS3j6A7hFlBGxYdjmxe9Ptgu6qct8o6CxtcAf
9U6GK0rgRKVuKWsWCvCyJaLvRRW4W4kd/PoFleIQGKvk0fDzfkRoM1HVp5nujV3y
2xU7/W26HYoqghd8cWNOgC0stjxx3NQCDQEIiSunb6aiC7MOiZ80VuU6eLeA4LGq
I3PEgqeruuMLDwolvE/tdKQyo5an+WrR5xNk+S+dCJqhSZmMqek7BRLkdsrrakDk
UoHpuukkoea1wViUJXisIk0Fvx2rGFwHR6uO1wEtiHwe1SaHUh8j+Yy5XLZ6G8xS
kl8rrL5AZEXK7yeCJ8FssdnId8gZ4Qw3Vol7NPFT+3FbMsOxyE8xYXhp95Tn0g7x
nhIv94XWjUnvqzgOcQqXnm7ASU+cpLJ7geMQ8ILjuKJOfVF3d0V93J38gG4JOcF7
lVHDZEONek7B/qf53qs/QpFPJ6ZV1sLyt7vBHfbQz3PvrdEbfSLGL9sazcOCd1UR
nD+XUmBm8ISFncMDbGBKTPhSwFeBmbBFArk7ZSFPzwotNFbOyvsItt7kGcejmmDb
l776X9qrkWRoPEe+V4amxk3xvQt0iCXuaUQTa0QKVDHmebWsan/yCqu9UFkoIhRI
SDP8rkGkiuuW+DSdl1JtUZ2C0Gz1eXB6dikEJzI+aPIKW7fNDbIroVGKFlX54vx7
zOFNVVxc+5KoZa4Sfw8Ie5LFc/TOY3Toze6ycpXbHMsidMxBQlXFyja5bV2exuxZ
i2qg4w/KSrCyF3uhviNjqQOO3rV52r9rY0/yWLS1a38x88YOikX11l3IifoCFhIF
F8nI3ud9kAdH1nrAzYE5fE69NrKUDOfe+zFPdy24PJYYG4JBIAVzW0+2TTps7mHu
P5f/KUNOgKwA0LNcx4IqkgB+HAX752O2rGfBQAATEbWTv3M0O8bIAKVzv90mC2Ke
7yWbkpMACimmpaqm34piYBGr/OETdklDChtT0mwPeV53yirtiIJdcKGiKSfgOwZW
HbbqQL9x0bZ+AvW3C8CXkXwTcSn7TQWKRFFa0rABBm5I1ZRMYw0xnVYIHmjvTtsa
PSw1TFO1JgUOsatCk0Qf8LTpC0LCw+8ZWgzwiBtyExhuU5b52Xt5zDS9VN+UOzJ8
w1PVjf81uIaNnWet2cauSKVsNZcTfGSbOMiZudDHTHKehBnaLPfTpRjsA2M2gevR
5JLA+r1+u7fKmW3qzAJf02v5vCID3IEfG8GJWelYDSP5Fsc6kBG5HpYP1vUGN2iF
S+9R0tBDTAd4hIuDZDW7tPd3bXzwGHxWNeDcZnD6aRoIrFomuEVSF9qNVqZpv2HY
LF18F4CYVZtLLOaZkZAXtbZ2tDBcyRaKskOaE/EdJyPwglzHUI0z6p6GZVLn3LCW
vj9fMH0LX28qA3NFcMlNNFZhKIThXQuFge+8nFe4zJ1vf36AbuFkmIJ9UZtRgizE
o6GOIxjKp4uo+4AP22HqXD0MO3TtEovWYQaZad3+HzhPqti1rdPveaXYtbBVMErm
qMtVnDeodL13mQFhPDIs7u3eGLZhS0/InVQmTS/LTuxe1wNfi4nCOk/IGXo05hMh
pp2hztO4AjW4NSX+B6YVowU9jiAC/sn1lgsCfOC/YHOrNi1Et6A+kyiLyXLT4ZXD
Vk4VnGlLlGOarZ2HYTgxqbVCP7AjR11rv7MrsYFX3+Ns36APV8fCOWITT15hAShQ
8eKGn0OYlYQtAt06TgHT4HFD2McmMhc8jU8eGG5vfjNuMW5mQeZsYJtwyvxK6FAX
Q1P8kQ7kxAK+BmdbwwGrtIHRoDZheazZx4+PtVq/E1ttk/POQF59RTGSxdznQjQL
7TIGCHfa7aJ05OWxtoNzPCHRZox8VjRN8OEGosE1nZ7y+NsG3DMmRwIdKynH37tB
IE3lhAAsyl0mc7UFp8tOYH+obI9IOTNoh/sYaK1p+6T/S+Dj78mHbkaWi+0XUsc6
7e+VwijmyyNgHnHYE3jrU9ygGhnMVO+q6/RksfDNUTBIvnHlGvrvF0sVFfFEQvdg
NUv1SY1cL8WJBIHvzAZ330/YHDiu5M1LKaGq02ziLBcE6MdmHO1rnTv5XGV7f1G+
c08FXrqKMmyO4DrsF4FuWYJXIZeRV8lBZ4rs6ECu//rQRPy/W4QC/YxBUS9Jbn67
JBQU0lcFdaYUZWr+fz43krfp1tDu2pdPyQXUSW8squwFvvqtDz8Wh0o4CvWzsk2B
p7Hg1kAR+DIvcHu7tOTmwJltuNJZDhwQkUy4iDVScgAAyFI25v8djQ6xvbRJRtd+
iUCJ30HbYhG0F9Tmwop2q4M/Wo+sSSoHZgZwZbS47bWjz/T6BUlhFp1caKcL5lNa
8eI1XA+SrUMLHlbR297oIT+9Ao/8G9V8jpYQpLo0vnnDImsfq8iEHQRJgeIASra/
wEapJYTsgKWMelUnCZbiz++RCsKeK3O1kBOUf0WH4AYhedVVIpkRbsU9UYeGk7tF
dJq2H496V6J4JgvPSaVBBV0PkCQq2s2VSVcHHg62RvIOHjB7rxmXg2G2CCsZbPiP
dU+63tmcOZmmows/1Gz+XUl3GteCwDC0UyIEmBMAZeRvJaBf/pVQHpWlj/e/n/cY
oAfJQaKY7xIIv+eYP3Vh6fe/x2AsTei441iGQoTnsKDaSsba4wo0OuE+GeZhe9dF
VAOhn6NL4onsGIu6+7/KbugIqCcijaeNs61Xd5rXmEzDwajXUzaIlJT7A5tbu0DR
f71hXTdZZdYLLpEbmbvMvf0AbmfOpIBiZ4OIxg8wXyrXc1yUrdaUqEmdfgLa0uop
zgP4Uk6/cgaObIdvbfT7GIELeeYCjwPZi6OSaJ5F6Yqy2LMgAP7qVyFsbUW+gkOe
cgSIwtJ+jAYdwChR0SJc3lDPumtRNA7U/mukqsUtnl+JAvjXXja28vGrQFlujs0q
prN7HtEhHIvh/fSYm8Nx+Ox8JqLQeweZViHBPiz4be0/uWuj+eVcUxH+66iPD4bP
CB5DFQDxF9a+6iMz9jzUlDoa3pgC24qeLJE8c4C+EaKCgyUq3ineGVpWK4PA2zi5
7NjoHa8tO/MEmuYovjLKUvf5bvabuTs2wwYF3oS/z47u20hE3bu+dXOk29qc6zIR
uC83Pabs8hzW2Km6q3EjIRUPffzojWbmHIhG9xI1qxhTn+oVum8OgbTWWTaQfAMP
/ExTJ1wso6QJBtcPXPvev4DZNC+RFkWlA4b/OhRQ3320fLSOHmQ24M9IKtlNBxcs
mYp7D2hoBuUIXOhhj+vZtZKJK6U+NjOyZfN8j+9Zyr+rkklUln64OgSZW8cxS1za
t43uViJxw/stjsf31wrGStkW6fA4lBLoSjXtgVyQggmC1PpEZOTsfF8yDmRB3Xdo
H+653CHra3rzivNvEr0iVKQmGq2J2pWnOD9snMmD74VZ+VADiC9wwP+NV/u2Zmou
mHdGvaHXzegwCuOuKNT/8JniPdbCiu48e/oaZvLRIJzzsyRXrzWRV23xx6goiPi8
grmmi1ud2l74A/AFei1H4Y6dJNAGoZ86GJJ79i7YOpF6UTI3DHJVIGBzy3leAqAt
+SWcpGF3aZMyoTRvwWtYdPO/6FvkSgw0y8rowplOqvzQzDLLt8lj6gSzCWohQPBo
+3yiSs9WF12uE8uWnMFDtdk+PaGcYJOuRg0277X9sruQUogg2/Q1Vx3UQXeuAOEK
YQbwvUH3oI+xIx6M1KaT1TW/hdh9/vh2B53Tn6WePDf6nyvtDqdDl3+xJY91soG0
Hvj8ZIRnehO5PH2pbCy89S4jRqjWNzj4c79ZNtFtJPuCsKLuRGj8YBQXPTKzv7M3
qF0bAbh5Q3AVBxYihM+MUzgM+S1rztLUFSEgToK6b2rmCuz1ypVFUnnpoM7+VE/k
FNwfitaN8NxavnR+pOUx+yvo+FwTTIxYhyInpM1Sws/EWiDEAWREn3gHB2jWagqj
DlF04mgzMTXpsnAO9va0zI0L/weO+WivWYsj28KirmfooVxTKi9GC/+HD3CYhY/L
tybYoUfiScdtQJ/rnQ6ZscepyyQgB3fqsLz1IZLDlwYTtUQu96YcS95rqvtz1M+g
HEMFPE/9U8fxg5iF6LvliVFNOysTwazLzvbf3epy3vBYQ1fWU272suy9bAHz3tWg
6LnE3N9iV7LTNTjLDyPoxL8IjS8VsbAjeztivcSxKEdEkRZeApXWRvLpA2UyXY4n
uOQu/ERYtD08xie5FF2XqVNOlGfQ/Pm+bkaVIy7KfeQeKOc/TTFjAcrybYEa3NRp
/B2kQPi9DWfUcxq8nVBMTCo9Y2vb5LBOQe8Z1Et63yWucQPg6sMvOPotFKg4EAPp
ZlwcJ6ktlwqbxAsh30s7VyRX/WsPFT+8IkzfmYxiGJz0hyJ2zWOLiU3Y489igbJ9
AoKkqWalhreXNltCKat8ndcKESA2jI9vQiCWrvKQqapNbkYmG35WnynZqNNU33XB
3HWg8Bewr3gjLIS4hFgB1vZr1sOjxYkb5xzs23PoRZV1k2ZSL64CNmCbG8uaGpiv
0AJtHlUwChM/99xjsRKe1MzbG9kc45hr89/vPsf8KmLcsFdvHx8WRgpIxYkxlKfM
G3SG3xyfpEP4nTPYqMyHatl6lbG4rdtnWq/P8tt9lNcKMHeOGivAQsdMk2j+7WYl
8tdr7LZQlhqDj+sf4HfMKoeG68ArxCK3OPrZFXAqPnysrdjNKXy0WWbCog4qoNuD
kliCuznBD3fhH3K5MQtbYEKM9ZPG4XXKW2RAwQiMrJSNf7WwFILrXwhScSBZndgt
Arim6wIpq6JUSjtYnzS4JzS5QAclP3ypMpif5cXRWpthNPf7zaj7EW5hZICedYKl
qDcItN02kEURz+DXMTFhg7RM0iyPT3gaCUCIBdsK7vW+fp2W/YgOLT+whtEa/mHN
HXQaZlMU3rstWbLF1nIzuCQNaV3H2K2sK18AiNz9SKLXartNKEsLJh3J6oNuRPfo
JJBJ9rxTbEAKbE/6BIH4X1JCQPFy0Tsp0OSu1prkNRheE+IxiYlNlwIXrrd5RPLI
SNybWepNjaCopmHC17xqrINBOlFYTdsWUuaxwIhoZa9rZa+bPBXu0bXvMHU69lad
tbNOwrCo4ehMzlnJ6EOfrN8XZ1flHTxwidrPxL854m0yV1DNGZ8B7QeAgQVwN0Yw
FrYtZbLfOc8y3l7Ej3LZ/ukyAqzca8NCKAkv9vNegXntST6k7hZnhVjo5QJeL42p
obZmdDLnSkqfAtTptCdEV/fllkQzpqFjrVWnVvmii+90OT3jJ0FQ5chAJB0RYJ/d
dgCKHT6zHOSU5OQATYMiBlpcAqyiCMkqS5XKrscEuWsM1jfCuRrMdzQcJYolSDC9
1PbrIrrcPlmqEGkDYWN06oGTmHZ90eYcw3m9o0f3VC1TJr4GkqT8SnTKOQQ/4ywI
VnDH2ssf2OrymcKUXhIsr9O4oxWP//xZ1MDmM4sgqS53A3B+tkyp4cpR4lumtC+K
2rCmydMDzV5iYtU1rB80v2vMX6/HldmrccaaPN/NgCc7YjujHTC6nvYtcfDt8c9s
De7gKnzbEqmBwq8k0qYW14yJU3Gy9h9gym3Nae1d5AwVMHsowbQfrOLGlcbkdbGh
LHdgx4567cvz0I23Lmd0MIWyQ98KiBqL2blZ6To4SP4uiK0UCVYzC5D0Oa8HpxcX
9XWaPGb0yHmo0A+OMdvctx9Zh7DeY+8RdsjThtnXMusgiDmWXPYEqGboaUTFriDi
hS2iaWu5FjnQOleHllEQDQCkVt7XcEn7aJ+pB6NkrsR2Zkz6vSarepvlLgvKFHKa
o+V+bsMLohAOOc8mWZTWapRjdatMwY+V5V6eZ20pj6tkTrJ2x6Yj5SczJortEnJd
duK7TUsmzqvxY2Z1LUo73oggCoI/oi/M/qyUJsZjfnP/iRysFFRqdnEDK3S/JEI+
dN/gahIKMFFMnFC6lf92U4QXXupkARlyASZVODh8/JeCIj6Q/WpVSgqmoExCT0E2
cdnfTVQcKxnw0DZAa6jdokGuxvoq06rzEJszIc8hsIqOjwPTht2Rs1Z3JKAxi0X5
uObsF4pFxwwRqBDcMSuRa71sxcR17VJOosjLq8m9ibX8a+YPj2OY3cnIka00UNVk
5uTcuRcKwRmn02unSARPFOBGSa9kf/Ojp1KfDKj6KUdxnEhjsZlp5FfFcmH68HR4
F5Nm6sRih6y51dYMMuDHnhgolv/Byq73Uh4dwSRQQ4Cf8KtqgU5+brItvlTDCbx0
nTyCnpTdIT7rwjljrAwEDHxF8J047Eew40fyC/7yJtrgfREtK/84ujtclfA26DIU
2t51wLBLpeNZbYtiqepWlIuHYvU/ar1wrYvoaYZUVtPDhnwHqvW2IEPADGIY8UzC
2QqmFh8JBn7DElXB6LHf83yF+LE7av6vT2vhzoCZHQ3sSp2hVEbiNetn1Ryr4Bry
cMJjm2oHf7NHKQ0S5Zyv8tzEXMDWsvcKfQZ7NntvKwxQ5Z8+fUL3Aorc3CNVu8Vi
6GcF5ZmV+MSx8Bs11wAJ4jQIjYlPJYyhQ9uJBXaBAfC+gVJbBwAZIGYnhPaL4mT5
WCsqq19iJsmLpF6Az3nxPi0Vrm8a5oD1NkffdkNFSKAzs5+zQrkR7hVx6N5O7qYq
Alxoc6IgmVTsdO8wqkjCGZJXjgnarNjlh1RDso0L1BlaaCke3tA/ovLpRiCs0sHL
q/sYN0hNQiyKWV4Z0G9I/wxpg1rqp154gSAFjMi6LU+wrqUI8XA+YqGfp86oV8g6
sd4bmkGd10dqDjRkb3B3YqRJbjvdqv6LjnQ4BdphcPb//+DhjGOUN+J3MuV06zq3
cgn20JgbgvDkoW9ZxGo7pXTxE+PwOAwpBYPE1+Z9NbZTpyCSh7Pxyfk0LdjmzA5D
lwM0GjgdU3UqRupLnItgvGYyEFhbgulTOHVkMBCLH6LJq4lB6U+ixARh05nzqqhq
KtceoLPxnAU0BH/Iv8CCaqsPmvRK7Cei4xcqF3YK639YJWqAHkBW9dpWjAPUS6b5
ZulnZw0xhNq40BKWYs6J1RpZJ/zJOjZzzLdEr7bbTzJMdRMqI1JXdtn7bv4sXDTb
uTVJgndpINglzlekz4FWa0C9JJe7dMAgqKK9mHULdvvY8W80/TbajCCxtozClN3M
EpCnpHHvse+Tjddql1sgLzck/XxdwFATIdkhwuqZkveCRqaORGuiy5j5FElj3yJC
gE7dIqKLE/mbf4RSi4Gm09Jjpq4qsv2fUj/JtQbjjKXGU2Cmxe/rwg36UdZyeG1h
rXE7+V834ob4d8+6qcGgiAJ/CzmHP0HWaCY/D8WzVfDEt1imH+gPRHBtqcjgsHLJ
N4jlQIBGoM5+ZrC8nQ2ZBtkY1uHGwwLmGKB3PWwJ/urqbMpeNNv8nPS6EOIfLdAE
4TjLE7mWurqEYTAkNN7DPtyR2vSlczt4S9a1ZBdkGJdQDCDW7/vDecA2mE32SKfs
AH6N/MGe8Jt/BBDrz2hpzRi2XUr2Li0exXy37ewNX9hqK5OpPuU6I0E9NcEwBz/g
nRl7IAssQy25JsK4KNkQFJd3wmKaMXt5UIxXVqkXKKCIib7FcL2iY4N/3C6eM51W
FrBNqxs1z1iXZzEF1q3qpeNji+Yxknmx119a31WPtrqQfGu0D9i9Etyx2qkfHuDe
mKJef9kVQOgjj+ngU6TbBZAq8pziZ8o4TdEng0Xq5k2ln5B7Zj6/X0dTtWp7OOkw
E+4rd4IV5iZuOOnGQMFK5XnRYmcEF2jbsvtc+qYbSiZh3CF4VL1optg9JhlfUxC3
zPtcyBcDstT1zdRi8gydgrxR0NdB75GgOa3fM3QHWPFuiYf6mQSmlqp4uIh/F0z9
jpbBNfimT6jC2A+xWsHgKK535xhLXaPn0HXFViPBbKMbO0kq9OFjKdVduqfcPqVk
GDllWjQw/11otmWxaywzng1HVRc4fmpZbfjEvk3vBIOQUc/Z6RUcrAstJWBhfAPW
RLw7IXThnfODz8reBkJTiPArWwJiTNEnKqwli01tW8zaONUhjlga8VSAXh2YheRP
pIYygUdING+iogsdZGrkUZF2/GbaaqBT+2s6DBUcQIKAAR5vfZCQaf4DAllVQOfC
izpMa52DBqXyRRJvvF07Gc+QcF4OUD2q77S88FOLsny7swhWhazR8Wqagev6hkr/
7fDOpAwQiQfzdbLFWUvVOGPFAW/xk9IHSsRPhtbr9qyWjO0qLtKcpxxonRM2jb/Y
6NZB7sVfkHCNGL3wf+Sg0/mBTITu+qKBPwI0vCj+uWHZFliEzZMqujx1h5prkRaF
H0X55NNUVrNZQsp/o0ilGst8hgpPxZqqjAg2RBudQ/naX4WpU5T+k+iZ9DZuttGl
3z29sb04Bcqt+Dom2FORV+Ni4nA+URfoGSQAMy2V+velZ5MUM0IvhjX6bDpT8VKx
nvRJIP4se6n8XK5+3cgIOrsvtdGhTOOnfEGmQGfGH5SUKFM/GSpb6utKL3reXWiy
8ti15DV328P3exYRdBJ343RUThT3I+YZnCM4FYvdq6gx6+STqDly9yUrFNnqzxH2
YakNct5g5j37CeKS3LHouYnDihIHe+bs2AIUGm/GNEfokzpHuaDiUusYmyl7FFNd
nppZ5jOOu2kS91l7j11nFKBnofqxhtKWjgV3nsEbdmgl4swu8hl2KAsGu2IlFFTE
MKqSemAoqydXb6qEg6nSq/kRCse9jAh2Yur5/iVwKzPCJ0Jmh4WjY2Na10L67Eui
nkH9AeqZ3GjGQEdND1JgqP0bAtd7xw0Z5ubW2JGBWyR6lCZOvWkYn4UB9wihH2pS
I1Xdok71LKNp8B81qpWKJPsMsA9TV7SLdQRTJATJI5v2mRpVgyuSndLRldDMSyRr
qVaY5oBlaIvl3/La8ftZ2kxXd+HTaJtCIkKjqqFVDy9rDh5AvgoFC5AGlLvpwbmX
piVvumac5z3kv16EdBCejSv5ZXwwDytzkKCcRzKJTTvoxN+HnWSxeKN4dR1CE2jK
wcDLG1b6YdsjeGIS+tscXDxPrHM5ZlQjchDd50/sQJR3pMGo//i8wTXnqHkpkYpH
3lcVfpWuCahQpM7J5L5ohqfxQukgvRdN4PBvpzCpOjOpGpwP1tShc9404jrrpqkD
Nkp0P5YBLqoV8y9hDpfwpVNJuobhaK1OEQth7cO6krCPleQN/qLO8ssTfm3oe4cp
n9Ek7t582q9efaUGRtM4CZEe3SkXDZGERFU8q+uEXS8LXIRuxWH1mB148sqdKp4g
JmkikcIn6ac2lGSfhFHTFChql4MBZULMMDdSyY9PtQe52/UUXokJvzrRChuvGDg1
6C+ktQvsm1onVVMGSnui+1LEDkhiGb1No4pNV7YAXTJbYYP9OIJ3AM8p/X9RyqtW
tFUe9QPP4fdeKRYeJ9xogaD1bsJrVlLxt3ZxdPfIAtfQcIcnSxkCtX4JMXCd2NGw
QMRCN5P2lExuSEJcjOiATHFfb4mpvE5OKnIMYsjWgCnuElVLMM/WeiD/RZfpBf1w
ErqpVkpPtr6GhYrLadMmPI7Io//P5WsbSujxWilDdHN2UC+gFAe85TYrbizLuPUk
uuLdPY5ZlzH4KOKcI3vGb94b/FLpxbkeYyeMIu2aeKXLAiOEmjXSUc5D/7Q3Oyxf
JF4p63ykVS3XU2Hskuilc4zq19EcUPBWjfzPr4Mv9drTnrs1u7kLHQMMN8gQ8zN/
3bQu/1aFaY7CrtnpVzZRNJHhOntGqszxkVpph/VbQOGqwsdOqHPLj9gZ6hIhFKO1
64OLpD9vmvlEWZh/XPoDATlAg/1Y/EkjZpr0OYLPNbjTj4VxMmofxarpyolIeGHT
2b+R79dJmGgW+O8l9Dvfi38Bjsr6jFULSW2txjjxw2g774u9GLCI0nylzMDTA5GP
aGuy9PSKeFciMw+3NxL4TKZS6PY3GTZ4pT7B74VBT/3+nECK4AJJV15zk4OaE/Q6
cztdiitVtVpPaGU1odHRHh4z2xprTUnXpZwd/zC4dm6qhnE9W1hKh97uyUWvFBQO
PgmyqOHr4OHF9C2zyex4z4YzQExmVTAg8GGUzY4BFOW2x++mgvw95UV6O+Hd0i4s
cquZ2uqZ2lqtDCKzWXyoVlvFGqrlSIYWoPuJ8z2pBpxSe9zgBrhxYth2UBRLNHcA
y8ADDfYjv53bSG2KaXYvANTN+ItqmKAZVSIc6lbgrIkaP89UEuy4bLNHAtpQDH0F
qauG1zfX7LOwHZqVXgpj8k+z+XD1+eKKAkwdyjroZqv5DYZ0ql8LeG9rEcJ2t+YS
AY9zuNv7cUXozTXYZgM6PHY1Pw0AAPfWAmR234zuLxbqylQ2TMwKGDVMxK0d5itV
Eo1Uw/v4UDQ0sFTuWqS2IsU6l9v6LRvJdCok7xhB51WclI4DR7xD3w1FzWJTk+Fz
O1/la0u+tFpVw3NY+Lw7TybuhHm3N/POH+IN67I+oWL2B72Zad0GFaQwB9GH2OmN
tzH+pek7hULGPRkmPrZO/9Ms3jF6xSnjsAeesfpP4bbyvB9PffZlJgzY45nNL7j4
5HlevsRJyvtHAnnjJryHgn3uzdTC3mOYh9DERW5GheR+ktp9hmH2mRARqbRLeZRi
BBYEqWYUCEyx18sWSSwg6kZxNPBKHinsEgLQMdkifBvrgeJZtRM1Hfb83UkfspIi
vk0KKW8D2LDKuP0gwlTVoBJbVSxHrYt1ElVekB3at72K088PJWfaGpSzkKyLj0CN
U84AmKCttLK2UmDfgi/tIo5i/i5LG3R2eIwg5D1YNF75oCYdWGIYp7esuXpYD6ED
4yWhu3RuMPTtMsnkAbiTw/+qzYSp9XiU3VNGM1iQw5Yi5yZTPLZYLQkXDTHp6Uhw
kArOgV1wkv11yeVWGjNKCxmSrIfrsh4Zv+t7iwoUEKYZBZAQq0r8n5roiJzrpQre
mNuQ0HXoWfCQfbB2hFEYui/UemW3MXDGYlYuEYcPn3mlm83etxC6MaFQS1afcYSc
hy9dO5sffBWKka4eukUiTci0NmOxYSBq0idPRkr9KbJzsI5msGg4kAm/utbWUrXl
ju9w/Xe0l0vMP+ogy2p4HYqNv5qPjIspWhx7zIho+nF2Er/5fp6W7P/Zk36P65M/
cj0KaP4kBTrD4ONVJjCeyCBgpIGioqqx1WlZv2zC2mYBSf+F7NCD5h6gqRxL+a+B
JlZzYDmKOoUZ+gHvvoG8sLXFuL9RU+I82x8XPuuBQFKe6Z3zJFRmJcmlXD7MfTAl
Is7RA/wfwVCKxRyXrtcLGJmKE5SbgDuP50gHRfaIELyyK7q1HtIIvvwO+8CdP6I7
JTXbRnZ5UmATg8B/TKlOOIFGOFEbq834JdrQWH1eMZbkgN0H82HIdh//Z62q94Kn
ngFeX41eRQd0USFSTVZvZqXwy8PWwiabZ/cBHq4vHx5aK5cSxqTJqXQ603XUfcLk
/O5DsjL1VRbiFob9sRruYy3+rh1WqFYI1JlEnCXr3zHiiy5/eRMzzOIEDbwCntYS
HVgVhWggY09/1jNY7f66l/blZTGhUCx6+d+qXTKIaNYpeszyZbl3GYJ4Q1JLRC3u
ykttsDbiM9NqJ/XlylQwLo7rIvRBDHe4DU79+fuvj3q4wqhvr7HY+bipZKfglg3m
hp2m6mm7ziaTRjNa55ftBD912IplF8HoAQ8GhkZUKdsZz0X370RLq5OzEHEEa6t4
aTeIhtEdZ2SQT2ODWd7A2WnLpK2RTOpAbYow/UI3d7T9OYPagsttpUBUQzC3wILS
hnHZUyFAEslwawFmUcPRsHGnQ/4qEPsLJywj28x/Kf9CqK8sfbLzYeR5gf+tqDop
/g1lvTGUMFonjAojygCUTQ+3FQy3gaRefPNPspAB80PM1wpB4oU1ZawrTJWO7bru
ltyMQGgJ9ZQDXiMIPqVgjw9uKH5/YcDepD/5yNIA/bJj02SFwYMlKxrsa6Nk5k+v
IdnpufL13EJZdTJl6pFNZE7DD1vK5CMlksUJ6+bX2Q71AzbO2ZXt1luduSW8I7+X
rMbXjp/Enpgbj19Iyoih/5C56KipciVxDm0njRamtOVm1aqRbSezMsah77DTTYGN
RnQuafTGs9xWgE66VkS90heVerwh7O9U49fbRLT9L0/2PHrFmVIYBS0VrHiJbIVz
vmRmGpDfGxZFja60lopiyIdoOkyjZAiuEWg4g5RTw7G4J0cqi8ogXBd0aQRXOZ/A
FydodECCNvH4zmWVReJ9K0vKnLJTdN9PRlpjPmUQ2wIzSAdqRBq34fEVo/L0ETcF
A+vQAAcvLNQwctgGvSl5AdTjknwkMKMPIhe9PUJ3nvsVpVm2aXKhrkWoKlKP1/Ed
s7U73cWbINoBxGgKUkEghbUmssLd26vBJT3sHEkM1QAGC8XEUWxB1q4IAgG1oRqe
/Wtv1fsN970ATsxgAgSY2Se/2GCt+G+4SLANh8q4KEb/dIGbZxbKTesZyoMnIpur
QOw7cyqvUfqszQJVv1ZiOgC5R9bDcGDwQya55AlxjU6pY7R9Ef5sVyq7qAiuONG3
kZ/RirfBwhl1x/v7YeE/J4TmcegQqsh3JOxtlca7QLN6FBJnRU0YfZURjPZoYiRC
sQMm7CMKi4F6h9Ok0Ja7hly27Y5iXyFJIMOkCg+RE+T+KeGQv/oknAKMWIIS77TJ
94mHDxZJTJiy3Nv/B5Nuf28u1Wjs+V7d5UhnpOsPooMfjJ4OBuFxEOkyz/Zyok30
T1WHBWquFKs8AZaYxw/QB1R1mFmgAaKUabzzP1aCGWBK5Z9gIp6i7fQAnGunLp2I
9zDJUees2qJ3VsQ6lnpovbOhT515eNm6EHhW5/03HtPedWq6ACWmvdMGcOJfH8+R
EmCDZzd/Li4UT3HPlSkTbkgbnIvu8NI/iNJYT9l5nFHHz+UjGNS9q+4Nek6z1h3J
iWI2+wpgtPjV3lmZT33hpW0P52ivCMBHhzwdAuQp2JEEFcQAmTI/gPmeALCte2G7
vxbL4qmpn3rUYBM2AZRfF2pHYJDm0fKek0uliTPB4P/MANhiou7+tiHpMix4vARq
H1GkHNtw7Zg996kqxLI0oJ5jvMpNUK1rQyaBEu5tl96RLduQ0CBP5qrKksjAIsqF
4BS+d9cMiNxz32Si/EzQfja5RIL/YXMBOFxMyNVwPoYkRcBJRIphUJcgP0jgNpBB
SvWYn9Y1dZ4qK9C9PfXdLkQBWoMwECQJfbaPsn+2t4yPlt5CNt4fX2ABEm/6OKVz
No6ZxL4tB3UrkQPO5yiilmbQZIy4nHzS5OchAmJZ7yHqCkwVwobOWw6IHyk+QrlC
fd6Dx0U0hNYXM03S6Tkx80Vgdby8FADzw6QhRKMVxKRA3PbQ74FtLrxtsYTbV9Kd
0GAdxmCfpWLQcocsqVeNMdBGgzWkr9BZq6UapKS0AphPYuXGZyssaivbUB1GV66C
thSt1TL27YhGpi47D4rj9W0WGDI2BW1y6Lm+/gTxKt+NAktd2XgY8rfO4PN/1B+b
VADUiX64ZCPtKhb+X6nmXo177EyubeQ28DryJbvVrjXGDhKLXhtcKt/geqBJq8Pr
tYb31+IDtVCKPxE5bj9RryviJ86/VNTddIMv/DJKelPH3+URzGiX+s3YmCEF89z7
ceaO9kq/ES1HafVCeqX34P5v8enuyqxC5PRz54RH7AV7rwsUedMdRja4miT1DKmC
XF3VXbweTgo13f5rZauzhEKKCWa9c6UjqZfdWU2/aSjXQRDu0lnzwQ++vPikqZoy
/DHklgVgoYgbdgVJcpPId/W0YLAjM1+OySEuwkkbUL9t45WxCVsobZ/U2JoNu4zt
u/4LmIXDpd7e5p1/JqTtl/I2pvzCyEVI60ydrNy7ct5D/G3A6i5nQRtbT5R6Wzx+
sfE1btxbGt/j8b1KIx4yA6Una2izEJLpdpWvLgxjirEQOE3/weLVlZgsfbErOqCH
K0ZV1LI8o5r3gXYXlfIiJTykVU2QUIa4c1j5fBgHZOCyIT2FVGQxV1Ehytjy3vdW
+VmtE1QZuuiD9+Hy4/tiWN5JwO3fBpUNelzcBKroPPZQuPJyJoMJ6L/CiPEwCfIX
ZmLIaRTIzo3km7kszqmJajGCSsB0becT5iIpPU0RqkiWyoZrwtoEL17tFu8nSKuR
lJr6VatOGMmxYlqjMnhpzTDcbarRPtMxnFdVyYVel2NPWna0DLWrt5K0wyt0a8sc
BotJg4RmgvYMdJjzXKUoEYcepg0WO52iiuE/mKCoY7dhpH6bX8jSP9VGMtbMY4Ls
q5Sko16bkZf/RbwnwciC4nSbWZa8Bo4zPheDCSyBnsYUdqSjrBPjkkVvi6iR5YqQ
YW15EZwGuUJSCNGVBZww5qsewlS9fnJRvYeqFbKSjvUX7gIqIOLrjrKB9AhHsc4U
4H3Ryb+cqWiBzZt8QurPYjAxDf+cthTdf5RYZKKzKxD/VOH6st5UiocD4oVaCiH4
BHJsLPrk6t4k1CGLeE74szYy9pjoPJSFahek0TER8A+3oZGei6IZ4KDhV9Tws/q8
goixnKEnS3PV/4Zy8j+SKUyYGd8/VwjfO1UNEH07ct1zaza4xuvzZ1CYz6UDi7LH
eTfLeqqduLgsz9tUeHtZ+TOWjO00ateF9NjF4C5Bu8rbFmTFBMbSlzduKdGynlEC
w8rMeTxDTU5vrte1aYGpsLMN5IVjXlNGLYIw+WehBw4pVPBuEI13OiRzbHTifPu/
Q+CsB2qqYsahDEKuh3+bBGJCo4mkaKGp5ozenUuT2qAb0ZFwYKvsTq2pP7TT+dvP
XoY8JqmnD14aA1a3EsuG5W586plOzZvh7x6dyt78eW7PnKYHa52TLd67pPcALB+t
5eRrmgzRjo0QSlPBkq+xfytoi8EYeGd06JCNvqsINNPaqDW9N6UnJevAPXfUODlT
eAtfc4wr7RuIVzMyqxU+QN05wwytAWNrHv0ezArLvA9PHaehRAVas2SYZfyRz/v5
nPh6MLmy3CdZGLvxo8e9zvj4BfZxSc3ZshfYK6GAybH4SZVTgfHE5IBBfNXsBKXj
HPjoKoK2SE5CdrLfPOXCrtwRqU5JrKEI6BY1TfxU4peN00XLavkmkMf1gZHDOVK9
8fcz/gDHpfkMvzay9xE0mj0pE6EbgfBB0oC08+fAbd+O4yE0n8e/OCKDHlhTJ7GC
lNuLwafMI/dWp3UjkSGHMBgRJJuG7iTlXeg80w0mvGUT/fKe3Ava4cASYA95H+UM
SkBfH4370CLps4TryM4cbmhd/akHwY8XkZZFS+ymAEe/xxHiB9QWublvKuszp1nP
P9x46EFEUwL2gUkXcvMtiG06VdNWkWvrP+KNFmTaeLbGryzujnYyqdkInOD6aVrc
tb6SXn9yYa5ugh9ixGHdLfSs80nPH1/1XXIAJq31dO/adMRqN9Gna+lxEu5mQMPl
qUoVcfI7mi0/RnkmNmPdFnIRxUFyPmpG68iBroQceI2LOM5PrRsvPnC2IxJCXWQX
evXXMn2L63lRFLOncu9uQFipAT5tNAoZQdnjcn6p5mbgU8+OIvWdBKiRcgiWScC9
gK7EPsNo+6hbdDL/1sgkBpbuKPZ1BlU+/dZAvZdljv9hkYAVT827l5BtnHhuQeGg
gv7NjKnHYzANxx9Pe1yo9WSHmlO8YPjd7fW9fn2dMRJ2KEjpBDNKpvgbxZZK9G1s
rFxooaTI/fA/m04MNLFnLkbaC3RLdJ1IgPaotjZY1OD70E88HDXTE6bBRyZpviIy
9M0nPjRhpJNlP4Pvzh+S+cE0+fF013JTIWaN9bTByf1ZphlG+tgSArUfnCSQmFsU
LBho9X6rVcdJQY39Z7fT7Z58lZPDWC9BVi3mnnHOkD2bXZRXOKh4izjeB8qsDQwi
AWqvVrekQH67tHQn5LLqCdTAzIKPP/sZtNcVRHmcCxeJGXMv2bL8MNM6t6TU8Dos
9ogZ9+VGjU4sdjmv+ssbZAJEwfER1pqTCMJCRHZVa220wL4KZhc9SaeGdCyGqYJE
AJTWJf6cMF81D93TEEo/EUmD2HrqAMaS22QVJvay50zPiPiQYXlPOc1DXnnTUEAe
RdWlzlNqcuMm9651yzVqd+3ym60QScynrfpw9jmRrPiK61M/5szSlk+s4gL8Lz+P
NRBj9nXIE9ZBO6TzW/QkesnI+iF6ZR98zUwytDhfZe84Sln8h8yulyMJsVZdLjMt
Y5w8M617lnCx6JmrM0IzqjHI2syWKHtdHTiiDfHiOcWRKGOHZMgScsP10T+enrik
TMOQ+F1niKg/xuwNroUtm0gT5S8nvAahpzuOr88u93dx9Wio0ImQhuZgDkDlSK1o
4hcY9icofbL3wRR1uYhWGN6kncjSh+N3DWA/AVD19zNZNRiT0QVnAdKlCVPPUxkF
6S3OnYFc5EZ5TWiUHv4uXOiwvAyEuG5cuiT5Rmh1iu5/UgUAZs2X9QwkbHiOi07x
U/AYZzuIdhcF8O1DmOO6oDE3Pqn8VNe1oT/ZU1cBtuxJauCSPJtEElM+4HSHgu3h
ZOLW0ZRkco9ntXqlbqg0xOIPqrLddWpP4eMYLyFep7ChqmxGbWsohbUwgS23lj/2
OYj4F2j544oubE8jucjwtTwqrs8NLda9T45dis93miS5RLs7mD3/jBkxi3erfOnJ
e+/hIGj7djwe82uwF1jET0ET01k9k/w8f+6jO4wiJAMOulWt05IRPninlN3vjmLi
U757/BfNzO1Csn6PMWIeW+Jb1Xz/Kyy2u0uQVDk1t6LNhzNDDhM3XPP+1QavRhhs
mD087SVouNrgLqLMwFkWi9BbdSTK/vISOqa8wm3rXKGFg+2ie/ft+P4eYPtMCasw
DD3wGOa98DsOWUCHnBrYy86YJpwdLpBcV7CauSmjS6JfVQ2VCXwEfltn3c2GnxBY
k6VmM2HVDcNl5NlPaIrYKZA9oFnbo2wwFw8s5qWyK0iKvVQwQVd3DPxD1CjgOv5L
X5yyZax9Q3kO5N7avuS9yrs1mQI4wxHVWpTYirACN4S5/+uuTMN+y8YiRtZdKjwk
alxj/sI1rJf6JOCOcRGIci9izCwRqPf6UIRK/vELCpuO+UJo05a76idl4yjEMnQJ
0XgeDu57qB0EbbZ/WptWSFYgE34VycSb/BdwuXi6HBTdltxVEHuosN5neBUv/egk
k7d6CJdJq1YS+rWYft4JVrnZSzvVYRv4QIt71/w4kO6VPPb4AiS14zeFPE/4ZjYr
Fko8pKq/OfXjwWHd+mOkRkK12wDT8n3AzM71SyTmO4+BOF0biYtHu2s7xtzgEvnd
OY26g3PJVky6gbCO+XNhtTFpKNMsmOjm3UPTLHvfRWun3L94v0OOve8thP8O3ggk
36xoHY0F23OL+5TZY+GyE2x3kvnKYyVrkmElVTmXYqHa6SjbAPhrvtC2chr821ZP
PrfyelWEElvzoKAvXNGVSG9cRoCOLgPyLaiKB9LAZHwgOSGza2N5ARkv5zdni1hX
PewiOoAMqbYc9KY0F104f48gaVk1kXjazsIhNMmnWyYpNT9lWIdBRgLWFlz3wKqW
gRGr1B4XZPjffguwnUCBALv7sc8pA023/wmHYdL6p3iZDGWUbwiB823Xz6HItKoG
jzgTMAtuch6MX5dYIS3LL2vH/oanfASQSNGTpGJOv9/g0H3fw8Kl/M1nV5ITPQ0/
ecxxZ7P8Z9Wo/JZq76/iDzvp45BIGPXmCauR1lTgjm5ULpM2zDIQ9IdnVxCNAD7E
6KNSQ3ssaZ3qSK5JYlm0ZAo9uyxu0eUIRwXMJwQt6/zTBmbDCVlFwa4/hxMmiyH4
RchsMMXLEW2H+8lVkI2g71mUPUuQno9GTFykOqMJimlmTIIfPZP1ycAJM6frvDiP
HRFmA8OPjWZqq4DBRZbtn0Q9mfVOAnv88xoCcSfYut/Xm9rJi0+xhOTdMBXoSI2t
aAGjT+ZGugusyaFrLhcceEyyWxp0qXPG1CQjtC6IbjR+UWv7PDGzSZlp+3fu0MIn
oV4speuzD8NxT522otOkXBcMpajJVbBimcShkQA8Uhh4A/9I9VL0OacJ2bp59rHI
WGxYXVTFspxrnE0cbcvjkwK3mkrx3dWYMTsSUaSUvggoeojRngjELQjqeBdb8J5u
cF0cfYWH+wml3YFhYw1jPO5/r1hzkpxLGhf/tXTTMSHN5why/VRR3cJAoF23Ekey
igeZkfPrZPfbqiVMNyfgZ1bePzdM5MMf/blZm+pncmTIJc23rddsuPJhr5Ele0zF
u3dxS+lk058C3dCpqgWmDmgUVnISgYTFmjlnAjzsgfeDYVjaPPAzTpniE0B1LQsZ
wyA8yk/0m+YdY1XRPdfdCTN9Nw4lbvDJA2WO01uuNyEFfuoIdRLH3BYJvlUmMoYy
57Wu8GYwwqUFUOa4tggFmhyabRWtbelAlADMB1lefq4r3fvjqWk8892HpAXHTUCt
t22S0vEFNY6MfVNCtnrPJqMnDC2ake1JG7BJ/yzY7cJ0x7K9EIzfJX+29U/bZP12
nA/xfONkq24ZoxQUE5dLU1U9T1rmgsNch8iJ84RCSgOP4sAI+V3w7Lx9VBOBTZne
dB5uL3x61ZwMslQwBAhuRbgaOvJejUhS1AFCmzmnLpR0iC767ZNcjT7s2FnSq8zx
tV/7PC6U0OCAooRMbktr8gh9hYC8pojsNZRHQEBR+/x0gP/UgwxqwbhlR9RlI1T0
zCrM9uE016tgvTkGgerfBCptPDVOV7L42Ef4Q8pxgbh1E662N5YfvieJKK/NUvcR
SD2/z74XCbB4xIlRkOjVuIF4M2LVS/iXRsxBO5I9qLjEELvMF4XrjFAxy6j01lYS
w9iqNbeL0rNxx+uTIk+EwRVBsexS7kerTWqeSxxbD8QJfwCS5cI5+Fw43McozZXz
TZPn8kUwsJPX7RE/CwBq9kY1dZZNtCABLRu3jhwL5WYhoctrncN7scd3rlpeXby5
aSlg5bXREvZYkF15T9EsMG0qShTi66s+BROg4+4T5yIavQwf7FyBRlAuWcJNQWNn
rmEtuTjyv1Mm45tS30S2jrtIqlKCxL+DWFYEpkkN4k2JyCLenyct2syxuX/wK//j
7ILkKJAURoalx7ZHvHX29uMWmIP8t9WLJQPuORulQAvD+2fErBhZScQbcqV/lg4/
8A3dRxzyfeU7hIApPkkPiRt+sSso2wWfLaiFfsV1a7CQ04U2p3Mfi4sghr6dgqC9
5mDtI+zHnqhTrFk5f8mcYtad7pdFqV3JeC8b5TCmFsi5NNnAgA704n57cZypkFN2
9y0caYPkzktgFegUolZ3LWQYU53E1RdXzx3T02YqBXx6MTOprkKL0XugCw5ri4B6
dj5QAbE3+o7Bzxouchme/iO/+YQkidM+jLsiUKPtOmvQBRSHXzzkhypyd8swUxGW
S6LBHrWzQM2y1j+39tGh5PU9fmXjeO2OyYEH/OpWYsr0jvcir9Wa1Xisy9paa7nh
pKaLG0xnhe/nJqcKjnuyJ0XobhX0fwkPuayRUbB48Sv3i8TnECZDD3q/Hed4vju8
S8/6CDSpwXPyymZFrm3uESBTFiaA69mY4fHftB01Q0QL2vLx8KmaEWVdU2REDQbD
SgHBeGqBRu+evP37aPl2Pa4ht93dVjZJw2j9KdjGIzYTxXD6AGEzmnwvRCq1+Qst
4BSvKyPdCUrnVuoToqMLRVvYbgg6+HYdZzlR9BKBYlhsZoZHMjJdTlRpDY9kwlzX
xkOwdSfmmeYQ8pX9CSW+NO+JJ8GVWsjk3r6gjWABsmDcN1Of5iEd0jRwkVO/uOvK
eWFT+brxqxuuYJZh3EnBP41hPrJnxYMTmyCNWQRaP8upiDBU1iLpUkY6KYgGft1U
65AFtIJBzw/JLZqOj2upzhoCPd5X5rVgil/jlULvNKD+WWh3HupwQC3aZ1oQPKzu
BbBlszf9gts+WPAi4zozjPhC0oBibIn2yywH1C2ea7+XKMGMavjaHRkbhKK7GUho
82txnP40pyXElhDr8ymY7p8qncJN4qsCLO2RgyDZXfDnUgRjXhx6egaOdbCGEkOU
JwpbG7mhOl/QHmoz4EmZqeQPXnHaRKR6cWMoWC7XXdf8ZhfAkMiW5FhPiYDGXBGK
3aT/L4Bs5HLpEfQAjrL/m6I2741q7x2ue/1/Fh+5zbu7axAKtn9Fmic2KYt6fVU1
QvrYs5ZxfETNdxtkiNRHMRyE4NJRiFlhUZ/h1wsHgTiI/3n3IT/giy8J2lyR43Fz
f4MWbobfN7iTf9BeHKTFx5KclkGZWecTfiD4xK0JCftHTJ7/9Uy5R4HqFP4sSCCC
X6Q0Oh0CMjlAewqpJoBJT3XfDXMPxAxcPJcS284sgniqlUXNS24YvHRm28pNZnmU
EznI8QFKS+lePKxF9ZsGpK6TFfAU3Uc2W9rMoE2YGl+qpLXqfnY6bWHJCleNOtGH
p8TyRg3fOuUARYKP9Drm+x06fa/+RfuhHazGtV/Sw84PGWU/p6J2YTRjRn8J4Mpm
2Y5B2ra/OqFYx77S8mYOjqNZFkbDCoCM3yOkqNQxROWSMeaFXM9mO85FxCulyL1y
rKN/mLfJcykLza5vG9L0Muuhpevx5mL/5UMeA8vLP0UiJAZAUsQjEz3L3A/gs9mx
Ze/pnp3PEeYYMf4loWmigbCmuUTiKeX4Q48wleCN5+b+JjbCtTQvgDalmfCjfjf1
32AgBFKYi+1ZtO7g0aMA3+PQ17GZUimVcglJuGPLci6ZZnNXx5Vchhc18fUCo3W/
/p/NfOVa7aYDhMIX3/XCjdK3kcUhL0+fD6rgL3UCB56t2eXWoP3NQErFd09sm8bq
SYbRhoDly1q6jXXHsu/TYgJ4W2ohRVb1qxhDhlc/PK71bIC7YKLLXvHDKwEV4eI/
ylPoMbbAAS38rZq4zdsvkzSIKVxBJsGeSsSUoPhwmgZPRuRVpSd/wLBLgVZz7H79
ePqZ2hc0hK2fYe9Y3wIE2dXC3y3g3Kx2LSUwbcpoKCO9Q4pOOmbMAj4YBXasEJ2a
UYjgf6EpgT208BH2buClj3wVKnbCdOy/qgwRKkPMREkiwFpGiRovZJ32klzVGfxD
g+hLlMdEE6BL7d4vCxnDeqg5iM/TBk+GF7xr+60UIGbUEdb+ERtmBBguOBA5wmCU
3FCrccQIsvgry4O5t108eI8L3rUXeMipiiAeBfaVHS4aN0rFubslionzP+iiLuDS
xhefPyKqnhnvyidexpn+ZF6JU5xLH3ptuJGlVuRIXHk4BLzG5ymzjnrCDx85dLbe
WYEVb+hL+e7MX8ypM24X36rQfK195fg98ZyfTLgvuMCbJSYj2rGunHdRnclZ28yb
SXW81+qhTUSV2jxZALQDjrEGxeewbC9czTWzvZ8Y7Myo8s7ha5Lxtqxyi56OPrzN
X2KsYF05RAz9NcS5sL19qwGUDzhblagBKC2ASgB7PWMtE4+hIkXFtIMUdLAxdLYE
p5ebN0pyaPDmt763jjkS++aT2HxHQ4K0fZNhbXyvXimloD0IWjvSnx/R7P70IbBq
Qgr9lGL++D5QyzvZsPf/vrd4+WeLdz70QW/cOep7RsORDqGrJEc3pHwsyJj7BpI+
rKDmP3+mlbPAnZ9/lOSmaOPI0jvQoAY4wZJPzxSbzgUjlzfXd3En1jLYIVz9CR5h
hby1d749s/Ft2TUJPIOW9z6br7IM67HbQOiuVbdf15Ol/yo3GmEuqRfOiIiKpLMx
EgjL2WT9V+3c7mCbzRukgRxRvO2hjX8NoW/4zNZl016OI/9K6mlFX9eTx4E9sU4Q
h17o1GRGoZ/XwCUDIYaKztTu0B4eU4Z5GOmRv8zUDQjJalNogjm9gTL8tM6NYbLz
i1oxTBoi4d9/kANLICx+2TP0JB5tWxhSO4nEDspQp7cvZxVuh5llb5WkGr2GyA0x
zvZY1O5mxvOgW+HDObg3oe+Sctx4bdoElf3VOWgyW6KFhkUdsUV+nanWB0ZNXXTi
yJ5RtX6HCKenQlQY3ZaN4oblB31dYx4sqHG76kUhereTsBkt2pHmwNNGX4R8MXi0
79fp9mSPKhX8Ki1MBuax7kPIuuVp/ddasUxXHhOA1kwxmIxTG+iL5KBX1NScNtbV
NM47MwjDwFDFwN8dk9AxYq2Iq5qAgQX3dXtJ4jOH1RqgCSkbnwcDIFK4EJOzkBlA
gWBCENQB7tz1WodM8LYpM4K8n1RtPYoxVoo3EasiOwkbrIaQHQbQXpRqdehE91yK
K+km3JOFDO081YaS9Ht4K3QcH7iVztSKLj3UpyC5M5VSQ03uEYhnjwyeM20mgIoc
vG3bG/1uJbC714zF8xR/JoWehlrMSITe21F7OSPXGUEsGHbJCooPUDTUqbcpSFZ5
8zXhbudt0yG4lS58ox710+uV9OD2rjxe43xb7UQYYIf4YVO+GVsPNXYwnL+U94YH
AW88l5H2W7cuZDBaLYschbZA0NUG/ZgcpZuQXE0fwbj9nJt4A1HbzB4ovBjc2mtw
KW20StZflGQrJiZ5grejN2PCVT3x3zjPzoy2D1RTMT+ECCiF3Q6qKgS7mQMjXFWM
xUKPocB5Jjb4RBSKWL47Xn0AeA4WTIHlAvHrADInbTTHBVKYo/pcWQxQAmRp6ByM
Keh5AKGgs9E4lrVa+jcnhmnJ/W6vbjPEgSO17lhS6SZkQkGHoxAQuEkyHrHjh5XA
3q+IsmQZwgk3wDdr+lYi+BbvJIcBfAtpKbHkWBbdJVhvVX4NrBTF/qCBgeKr5+B+
0PNkx6739NcTG9Fpqv3y/JYyusoEnsSX3flDKTdDCP6wVEQpKiuVB7dpK/kev/5F
GjCPnhM66XA65Oc/jEFxQrVcb7ypM4wE8LMV0si6L2o/pEVU1B1MH+VO44Rr6QcA
slgaeRx9xCPQT7FQHonOt34mxGKwIlmWuKUNa4Q4drhZjNhtrGJ7qSPRMM1nqV4f
QSU3wiQ7xQ4VLFNnp4Szd84Y6yV/EtF08xSznw9ZgIbGvWuNpnl5QjmuLHsijPEi
ML9KmTVvRrXBcSuYpjk6oSuaIvelLO1HCXxKoPgcPU4DE7YDcwq40s8UyxbaSRW5
nSveSr27oym1/4/PmHKhHnATLEFdRhP+vj1zg9997Y7GasrRH0rviZ0d0cQM3eQw
iG22vJpMxP298Ea7yAePG64xD/9BPCT06GjnXDdA4V99kt3HgOftwjPloaq/tf6S
2ZPEa7ezsBxF7cUEFs3PaSac/sPLhUa6S/fIdVM14qXjn9liz8ybc6wu2BIbTZP7
ElSaeDTSpr3bG2356piBlgeUm4xgY6IYp298iXKgMgMndWgBC6iYL6uSCW4T0G8o
Oc336GiM6CNX9FmqNFbp/fHazuZ8MADxLsnF/Fq83pvW/1UqVerCyQ/US95W6EoS
XcpIHzRp+M2roK+8cdockTE5bDIV4QsvkT3/1mdqjLD8LDsrlckChTUDoI65CZym
pZH8gbX+lDdGd4Cul8NtaIB85SG5shjYWiulHXJl4KTFEOZZBoUfAWwv5V9920+H
Kp1oQfcEYsVwmz/I3Ct4SupI1XJK/xZ6ginfYRPEY+LBZ3d5PrUDzbC9JKwYcOHs
97CHTyj5la7+e8WdUfVTCMA+ADo4MNCrdGL+Al4PllHbfocYoUSvHAoc+XRkTuPu
qLGWTMxV3NqH4EJgQ86UCsOn8TybERV2syxIg+U/122WQZQ3N/QNwIrIZpCjRPj7
gCsoN58N7ALePmUHCx++yvijSKq3KcnPuhelAfdjkHGlzUxW9dxUyYTJg5FyDn8q
6nRAmKWvnAPs2uyoOL2ibVcBI8D6XEfZiE29+wigMQ82rZAx2eaciLv1IjChHW0K
DKoupnQDgW/zanuJHJ/bQzPSeI7KxykV1bPlGrtaw5lNuHjEtGPWBvd7zrr98fs8
R4cVJyXtVlrFpopeXWVgkiGKRogoLXe97rdGzNK0HKwt3nXGnXwuh1rtLIZAb9bh
jC2lO9QMhnbFf22BdC3xbGciLaqjP3/xJ8ujt3xkvX3q2fvYTiWRXnjTrJbYk5rR
tNKacapkXE1K05wwgJnjsD/FweN1jZZ5ocdwmxMB6GUqOs4Plg6DF5mpSHxS0jnU
xTij7et5b8SmTEDHCCtDaknwBEP58DZFdc6LItj0mLugN7PFRq05jO8TEbNXZhKt
ncPVRno85cG32Jk6F1yCSkGxOmN7RzzL7/oimCq2Zd8kl5fa1Tryb92p2dFoN52Z
rtS4RoffSUDrlLgV0SfQ9gvopYiw9nbCat5p3nSAwQfHBsk/bI9sNjn4xEm/XwpI
d98OsHkGfxR9ahdKpKAfy37FhsvsOcnMfh/G1PzPBKK1eNVG+NKexZPPOeAquyaP
MxkyB4BmzzzaWQhSQZmfJTypsZfQ9iEGet9DDPcLlclxAzls7+OTNRk8kv83GB25
jHl+lOixdCsHP+Wjg47PH7EWmCh5Zj7RHAIURFCEPnUjyrG913cGIH9tdn4kBK6e
HIbop21086D6obFWrHO6LI9Dx5F1Ry9+EIQOMDI3vMutgRhX1TQYrn9rQeIcqKPe
9Kq+1HmA0msb/2aDS1UO1+mYVRKi3/YxfDFuQR4H/NEZ5f9UvvfSJbaeEbhuljX/
rTbdHmY8vK+lAoYK6lFPmfAIt8CIncrbQPOcOHrin2BZfmjUe3HPYRySAx9YTBVA
kPc0xwlIKsV32g2xJ6zPBDXLI3xFBEFRqXrjlc9W8EuksfDt9qY9IrlaVaABZvte
zP5KAz8iMkJKlEnqm8M8UiT+8/ZtofdD7wIXoGzD5p6sYFWwn2aj5b2q/aybZLms
QeH62qm4zvpPjN7OdB23iSZLNExFuIxAUxF889PcIez1Rgdq4MwYgtgTUfyIypVc
xm44OvGJg9yVV+NWgU/p87TM9LLQGEPzdMcGZNW+tsZMXmne6Kv2OkBz1NMLn19E
mP7sQh2mkMbdUv51SdLPAnE2Z/xi467voGRF9E8ga86hGeVCrja+CFQVTGHfLsxS
EXZl94F6XxqnU28PA7/VrtnzIANhY4SjtDobsgIiOtRriWlriu3mCCjIMAm7KVWy
CBWV93uHUhg6B3b4aHAw1yIfptsxkwu/B4NxeZV+NIW21unyF1+bcrlyWcsM0+EQ
Ekc5aMUoxLXobkmmTKz9jb8n4codEQuuHmO5h8zk5+mkgtS4/qZXg+P+gb157Mys
yIvNhC0FVWSFJME6N8j8fipHLJ0AECwZVEE4UAgPQ5p0O5aoMY2WxThPWpOA0jtn
mcYgcfwoSZwCEAUNAJXeOEjfodH286xKIzLkZcViWh4mSy2QrR/xyygVFFSxIumY
/fFQYm6C9+OAoPE78aBWpSxG/9d2DDBzEl3YsVv2o3YeVavOzi0ROwHeI6++IedV
Lrw55MQuTmbZr7I2MdZVFd66a0k+OV20b5XV4GzoXK3RQ4oAh2DykWDCl/lw87Lc
1Q0UbQpcn6z8fdp8XZwsrfuFarT8QeyooRdY3Lna8EGA4HSrjpK/KyLD0U/9Zd2j
3Vq66LXJY+ELJGBMi9TuviD1ZpTEVOw21moN6xVrvrKO3hibcSehqYHFWaUaDehQ
Kqd6A4gzYFUxepw4XpKPJXA6h178FuYjqNC2xyUh8rjstbAEOvdv1K+oE2EnugBW
TUVaHvNhXLGbcNsbWEJTs+OZtBOJQmbI86oFN2JXXuiMKwzAtkC7if/aHHO0JXm+
k9iM6prcGOhHY2lwU0UGIpOL6wpGknNyWw2GhzRslznVNMsqNM8a/Q0f/20D8eh5
yPiZ5rY/CCJJRUjVTIF9rVfimuORCuJSDQwj8O8f/ks/ep0QJJmdkaXs7HDtz8uQ
P2icCt9QOw7UO1WIm8YTLDXektsgRLvaYMH2heozNxccxCzCZqGYqxB04kEAAcfE
m1CbU197TI4SNj3a7E+Ik15QOUucN+Zw4QX7qrOzZ5wimIo3FmFjY1gYvtSRnSiw
fgtVgiXTB+17G/U2Qu6u+27ZKFEHr5ZKAQt/nRLCziYbOGhTJKSzruAv/8crfSk/
fFdCZf/px8ykYzYeKA2AQ5svYLQGKg7JU2THhoxWg9UaIGPlQ1OoBjET7R2Lb5LW
i+/qIATe+AQHRH/3X/PRyEGRIkkGvsF4XSN1y9ySO/jhnA60v52hQh/kzTvcEAt8
2/MYi1CPNs2jwgcjbifQQ7mEnkUNsfbN0OtkYDyFe/0LGTLc8JCKURp5qgn4cZuw
hQK5jm04WiPRtWEWK+bTdQcNY2pLsFZAA+um2aF3FMCoA8gITjxwaX+JtypDVtzs
VsWheCaRFpCHmh9vy4IzqdwyQt1H/oZ5s2206LO3/PSEmWFJ2XnSoVD87X8+TRLW
7LpldAZLzx2/SXReTVj23/Mi07yIj1l9RoKlXzp9lFK1ePbd5WDl5+nDk66x1ndr
7o4q4ePen5W9eVRDaJbFO1fYNIkkEBZZvt7lyYdE7zB4z22iIrfD7RdCENjPAMOy
kT6LgmL9wloe1ppo1n4cneT1Bulqoh4IG7ly4ZVgkb4+fMgFw/dAVvkYEWaUdgPG
iSSVZxv6nLgR/5qAKtIC6Qy0GHKLI1mcxt3NvSvHNEmJO3qavQPi/FkT86teUB0Y
4wfbmF7pC4ATsUy69YtTh/07xksvHHnTk2XPQqn1Dmd5PNUjbvG7xyEZskj61adD
Rs1a9oeUURStwGEv/fupeebDdY/RRbESL34AhfxIlWFnn7pqaCYvC1KqTzXPXhoE
0yGD3MJR1lkCFr4GKbbLB9kmRV1ciEJQwA/CmGlI6JINkGaFvfnzQTOEwCGIXdAg
7ykAHMrQcK89RgrkymTYNLSz/UWAu3Ixz5T0bk3Lcel/AIhiZ2+q+rDx+ojeSgJc
oofz7X5ZlTvOEnI+YZKGQv3pSD5GU5t6s/4TJZoMXWct82zI1dXTHz3oC1I8+hF6
Ui8Fa3NIW/M1J4NXztfZc2Wc2ZoWgV1NI2yoviolwlA8ISQ5dadfO/b2hFG6CxVy
DVUrjXfZB6kUTBLHASin26uHTYc6FexRJTBkf0tDW48fwXOvkulEkO64pb0AuL/f
wv+ibVNdybEIb3azZMD+VAKYyhCHIuzg4k5LnaSEtIQ8uC7k31N4TRRMIVB6k/sB
/oNWiGpfJj+jo9Mu2Iw0M+NzziICgbS8IbjyECvl4F7VahOQnqb7daI3dMA1EOIT
lXkA5f30W3gZ/lv3moBgQt+dN1YU8Gd3tk/7dwRlEOIwUOICl0TL+2FD8rMf+lqD
ShQrJu3RGV9Y8gR9ROH/EL1jF8hmXsDKIF+iCdU1drOoH/96x5EvjEOE6Ma1zZPo
2cVt4GVhnTMyYm+ZaC4kRBTrnQXqbsS69PE+Ix34c2gP1UgGSPBuRgGaNnk5cPXE
MkLmBPRrB8kQisPA3hy6QOx/XU73FPNeE09PpSMUh2ri9/UvATsl/+UaHFQHNwnC
VbtAzvzJAbNXUkR7mZzwPew2iX0nim8sytWeKwciZR3bWWqC3I6LHR/uPSaw6mEO
pYVrwNwhGnqoGMYmncBTUEQf6D3flNVBaUCHfSN1WMoHn/yzFrfiSq6yrWyhCDT2
1jvMH6X4nU3Cuu7fwpfVVfBGLcAcno63hG8va05ICikjoYVYglq+s/HoDDy7kZ/L
OpyAptsQzqhjhqW91xSQ9LXaWAXw1pVBvQR2zGaaKALYR1LUdHfJZMhZ+bAEuEXF
msH//zE1w1EI6rWb2qSySiPXTP3JggRBS2K6ApsprobcIskwtUtzz4jXYWJ9X2ah
LpHYLOR7ZXyoMi4MoKUXaGhX9q1j44+2DD8nJvOLrhx6r8kIk0VyS77LZ0R287s9
ipuoNvRoRcEEtZw+Lx/Io8KeNoDZhkOvXpWBl3vir4krK8pwnJZswKfAIV10qnqG
tn7lpe8h1HVIFwvtKV3wedJXYTrgymDCZCspTpNAAJ7JUpocLxG9DStyO9BhzVoZ
SabXzpzs9xTpNnlzNIm6db+ce7N/Z9hopajAMqCshv/D7+W5j958oR2Fhp/pYH1I
5RT11T32bvPE2A09AmufLJz1LfjhT9gpJFarbYivTYpRDsHk4nA7bxFkEC4AKpcA
dq+i4GexakbxcqPMwUvUDrf3mWSX/2Uc76AYPZJAeOd1NvYuccPjN+o56tQiproL
QYTSdXczSIfBKGK1sw34YMKIhkU2BAwM1qtBgCKD874oh6YFFA4VUaA/RKL/0aik
wnf97seCsJu5fqfEiL6dG1PUlsrkxOZUACuI9StigNzIjK6GfLUgcXB6NQ2l9EVz
lfMOHT3fIfM4RrNxAlzwN0S3E1e4VoFJxDgPiQRu0l/pC1DZFxQHZQ4sA/zk5KhH
ALUfsiw9gAd4LrmWLWCllUiWO+cchpWiZx7roNsu+5eErBOAYeJ9ofwAmTqMZA4q
I3carxTzOtJaCtPgiGa7hSv/EbeSA5GLPzSBMsue23h16f7S9iKoeub/It8OX+I6
byXAgpqfL6D5x0eRSIduSGjllijqngYn2X5qHIZRC6ih6WOfnfUk/btw8zzHCNfP
SPe5UtarXgl6qG7Xp3ykMngXOJjjbql14fLJSiR5T95B32KLtsSZP12U3EP6R7rx
++z82OB5zuerseoIP7O/kDW5cEYXrS2lIuF6uambt/cRDPf2V5HC4QoTJg6uV+iH
mmaAiMdKGR7w+xozfEZ/sfzbPSwZ6MACQAE9NEgWxftKQAJVtU7jeK5NfcjQr25l
pivpHQ7dXeLZIF6PARpOsesYi23c/8n7kzw2W0G6Q1EacWdeDyqpwAK3V3gy+gLF
OwyHiLCI6MMXBz8VfKGmvAXWufO2o5ylxq5sdr+hTLYyFcClG3i8vbfNqHIlMF1w
KM03B2sXX7D8E505F9PNOPotBnmR/O+lp6/JuZtatYGqw58b8hE45iK6p7F/numM
cj/OqPNeKK6HqIQgyFLA0YiLdqSUHYI+TEUyY1APlPoDmpCO7CBVvs6nHDyVQ7dC
AvIlpp7yeyJ+rus0HQgd/dE3orC5m5QShMViLV4lthw4Rx7bVUPXeg9XnbvaF/sd
icU6YFkJwOHZDcKPztj/nYgq2R/0SKSidIFm38+0VGLr5Vtd9JUhSMwVkJsS7OGW
+z9nNwtVpr6b+ZnwA1cg7WyqWoLoGXaOEln7Lh79gG0vXSKCb2MB5b6cGvBpTbyI
8TmOsg1TnqcklnapYELOnhm1b1lG1ORjTfVsfz5vE9hamAaglU7mEgv1cLl7LPAc
L6ZxEgAeux7K9jj+b4v51nr+/y38E/+HawOwe2/wr/bmY5nMGKXOCfeEPYugwFHk
6MDCsFgkatdyKltCz3Y9alqyxzT0kBDNX/uzSSlPWraSEgX9n3W2wkrX1VGFtSxb
KQRlPpuXRFcQhxVK3NGSi7DNSME+iUj5IJdh4QU/iIt+A0Mp4odVEi8M+vAUkI+W
rKgeq4baR3kAmixfA9D8/dj+CkJohZGYQTW1+1anC5RgsZ3/dBuG1BQbc6DI5asF
9pWNYfek0I9ekpiWE1z0oi0eMEbcstq6Spkg80R2rw6QwCgjp3uEzRPKOKHD2FNZ
kiRvamiXrd2ybPvgcp9g7LW1ywcWLIcwkRF9b5g8U8fDAxswbo85pETztDxPalHC
xuG06YWQ3Q50AkIwa/i48QhXBiYRMJ34QMse8eh2PrAK6VZd1/HwJqBWmMcGKUuU
/rAbeDBlas+RIx+HKSGQPuR77GUhhFlZe5zRLPA44agAfbwkByU/NuWofTKAnu/B
NCHb5ad59hNQAznM2UZ2wTzu3jeEfOR86HD9WV/AjzJt9ukEz+3SEJLdiUbAbjA8
94ShVLdTJR8CJMXAUABkj3lXV9aFPAPrWXs298gNxJzZI+xY6x1a1eWYpsulv6Gq
NbQmvISRp4x2fwg7NHVn3q/9xPHw2ViPpQHCBK+ZYbjt1jCw5cE/eBouAokILAf2
RvwAZuu0xqrKaq6OxOEObunEQ4FOoGPmnzrDO9rLgSvNzfu0LP7M4YCSMtRnwEoy
5yBT19Ue9r9bnSgFW5xtQ5C8RLa9MWNpwWm+I4J3U3QCoDvc2vHQPwyAvj6DIZCY
m9zc108uyjLWac1OLl4Kx+rDLRSrx0/jID7nLfETFDWWdivKAKy8/NRHkmD963sh
B2StMKzQ1h0XvqSAV1PaKEfz1FTIfEziOo32h+gKEGqAWrgOHafMXkhCgoZ8veTS
+zLyrucgLqDMGOH10FSAMarSB4LblZQqqJHeh161zAX0IiEoVoUqvog4uBLh6HYj
K1OQy5LJtcKc7p0REZQxY/4nsR//QKtF+TV7QDcvqvkThxika9/z6+FGvZnr55Ym
haT+EcJV4Q+CBk88TVx9b6VI7baQZJidhP3jc6iOL018YH5IFsHV/0wznmlZkD0P
8/V9UuSjnu20QWIecf0BeNGSZUPV8wq/LdbXLsz7Uae9w1zmNL54uCeQGCKDLt5d
j5LbBcalksUyd4rdPwxTAvtShHnIzMVl/aJh1z5hBczfrUg1spWa9cUYhSrX0Je9
ytpiRt7SnaV8/X0OUFKkLJmgtQIgA+FqMI/xcyupvR/ZrjpvvZfkW+aQ5SMVQaFF
MzhvDshO0kxfF55LSP/hwfrcGDJWWBlOkNxXPLs8tfOo+cjNz4f9I+l7ncfVWW26
vqAS3Je07hAF0nVJc9dlOIMaA4KUM882K4tPhQO6XWDDZTvKZlWiiDEuunB4Nq3B
3ZNyQupk5oqe/WRuip4eOg/qyDP6FGC0AgUaa78LZPk7HRjdEKdOZZvFE51nAPxR
y1x8tiXw1s6oFwyCv33PvxqeR/hKz25IEzCNkY4R7RmvkV1TtOdRfnu8dAd4a878
SmEq+x4HfUWG1GQKMSGdv/eN8VO/VkLojKfvlPOTV8CCVd/f7nWQ/XQ/fVgOJfEz
Urqqc7MEyi1CDpFBykx+ViaVI0yKgDAF8xRqgmcRfSTGMJV501HEpQ9vRq6ii8gd
oGH+x2PCKk5lroNcXsAJmPlTfFnMRJ8PmrDb2Yx49VAs0ryb/5vvewYomFTwOY+/
r/UQ+oeLEyH9V/n5uIbJ1TsVYFBQwgQPw0ZJBuVs8NB4xAheN9xt2bOWBbKNfAE9
CT4qO9ZGiQrFsnFlrMhQWEU8jxrjiBeMJUV8qgJywPxCTIOZg5mt99qzJ2jwYGd+
ZNWdeWZRVJDckpfXaM4A/JwfpCCnD2R4dZTMzs8NDcrZisqcGo9YAKsriU7oiG8a
YmpqhHYM4KLloTjb85NdgygRCRP8a2nxHUHCMbaCIpTs3uygqsD7OSkySKvEBBNi
twcQlMAGpjxELRFcMgkLoft6g7ZkzoXqGmMnJO7oeAqe0yOOhHO5MRn4RDv8xs2i
ibeoy+fTaKyacawaWGKKPGmNQdTbeIGedanFhVdsUpWESHIEPJsT6Cnhcvxg+LIO
IWRNksSKohVE0fg+4qoaZOhylCdD5ZUJCSHj4D0zLPoCwJ9d89CxDk7SvBEq09wm
3q1n9jnMrKYCSc+faANmJtxQJA/PXdpPLppC5pGtKAyQFy0NV5ckP+XDrrKUlKQd
b9BQ06BZjMoy2p5UYuJZx6/GtZ9F/AdLyxnyorq+W8RBJwA8i9oZiGheLuTBsZ6p
BSqFXDnW1rjz+UGLQ8qehUTc3OmlJXjC8X2gb20UqmMBggvTPYpo078o65V1fS9E
tgq7Pb6JPtLSq2jrgO2ye8r9ZOt3gKypM75qnpOkB9Tx9EsDHj7ussTGLWYzqp9c
sCh1z065rfSM+1s8kUMx1xyi6fMxfc7EztDP76sSYQRGZgzM5jiF2O3Bl8tmhAxm
qVCYqc8DYjAlfrF8DOPowpB0RcErDPoofsWm0s9oxLYGrmwHPWkflmthE9RK83xF
L/9ciFXKBC4hUz2E1Zu2T4KU4qmhEDZJhqkq7uggqLY8EAuaB9y9d+n7UBXJZPw4
V/ksLUk6n8R1qPSNpuNM3sHGRHZtO4DLcVLmjlTY/0WEP0BFjcHspW+nqfdQV/rG
WVFzcjFNSD7Kt4t0Rkqopks4xgTVQ/+B3urGAzXI67HueyHdV/mXFwOBaiocPyM4
y5KR2Wvbn5HRdf2+G/gmmMhv59j7d8GSs+2fipd3O5k9sm7rvR1oKwijH5sTnC7y
deJFcar5JgSsOad6AbLiKzXimpoVxmhm7RR3MeVlJn+/SDgqKl5UId3FaQ/ZjDHm
RwXrkab7b5UkKX4+i+Ogo9udUBY6hN4g9OryGBasf/3EqxZhC8mtYiptizxaRsgX
3vqlQiEvZGq8J4iJD0DF1nxvTTH7/rxQQtyNxvWXpqNxGHUL2WVgw/JvBGPr0Mpq
LMP2D9hHP8Pi7ks/RVIY4rVStj9P5cj+lkkdsVwZnumW52HkNxtDY3xn3RfZ2egB
dFs6g1RETT2FIoB6+wNMghP5DWyiLhr/OO/e5Jm31k5xzFnDdYjrDEIaTJbAt8yi
ZU6QnKHGiXfsML7NriGDnE0Qra5bXb1jRTMrqy6OhwaFU5PESAHaIfxjKUTvNXcY
RohlmL+t0DuehiBqKi4v6gb+Pq03HivSUr7KXitTKtTtY1pDeHwqqQj9plKwdb3X
O/4TGrngs159GIqQwMR8uFfdr8Hq5CAtpIsta9W9Pzv0nfADgI5fjq/cw5kMDM1e
bmtiPX2eVXOOGLTqFzHFY2///O5U1xxjOq+dKT3AZ4kaRfZTQlj0OXVO+quAzk3d
gjurN3JAXSQ9y0vVsTZfjMWZK1GuCoON7c2HAhJbOVb0IdCnc5yqabAcEHKCs7pz
fOQhV07gZN2tlWGsKLuUz851xSaCK8zafTrd+u1KDLNYC9rLnfFrMLbG2NMysc2B
gUT888cxWmkSaguMdB1MbfEDwyYaAsEQvU/+EBuAcA70g0BhiZcc6kOhxWiwunrx
Mj4nE3j5pw5ZV+h3D08fdAllnvOGyOIySmUvD/PbVlXqExzbdIbzEeIs1q/JwqLo
LYBM6QjNwUFtrSlqGDu5s8hB6qT1bbXcevaIBzuzGIQC5CMbhPI3mGOe7rxQmKB7
rPBHt2ZWILeWNKhpw8k6YErauZMamxPn4VGZmGDE9LoK7tA1CzTUvy5g9MXLe0Hq
rB2xVn7gtE8evRIrzJSDH1WN3W1FFx2QTxldEgCMlbSiaQQBF4OFNdw/F92fr4bW
yvzVK25JcbGmcNLBP41AN1xRWh5TMxAbENJZDe5Tyk4OnK62MJ6YE7uIpkdqAYNc
pYbvunldf1G1agpGLMBkHOUkxPw6TmzKBtISFs2FpSfLiRlIDA3iEcBwvf17g+eo
6W5KceebYq1TZohBIw0XiPUUir7hO7gVMxPU3WJ5FChr5B3hLERzLPpavu1Du7+1
nKytQ+mJbXvcDnPTqmoGGFTJ7JWFi+FNjZ7Gp/FuQl3VvvG53oyvBed9y4MmLWet
c2zJvMtdF2u3OjjdfSXRaeyFFRMk8UxYpay1u69n1pwN48FPuUYK6O3TVUkobGH2
tT+q1eFYIv8cU/5OXvwk8Adu4vCRX+O/kdc6k4ZDulIf1VJqW/unqOO1rrPlcZAv
PClSVVeo5gyL/rqulQg7syPYovDPmn4t2WmMc/LrbanEgG7r5IgS0U3DPZLaL99L
uaJnmqPhCIvycBdqN28o5itLSwTRF0sIHcLiUWS43SmjvQLco5WD7j8riHpQDOZE
KJOAUIMLjA4mjpRgCQBh1zr49Fir1SaI3RDq+7puj2n6yE2CkvC9rZ8HDyLEdq9Q
NQnws3cA42IIAq0/vLtQFKshJ4GHMYq0ywhine9Kkcr/Lzk6Rdq7Rh7Z83coLjE5
oOUGXHoePOE4pOXXNe/ZDF/6QKP5YwLJCNerc1je90Z+GMrjQ2NF8GYvnKjkVMEb
wEdH0j177p/p60cQXpehYbiciQFB9vyu4tIrBvucaHWBkWlBMtlh2pPKYpLaILN8
i8M5g9v9x++49XFAetHgobhoFW4eJFNaM4yOQTxt8ga9CPcEgAU+rxTKov/4iR+Y
zUB+Dcrrk/UsktOUpZKWkTCr/yrN4joAMjg29t5wE6LltkumF9P28tXkAIn+CMBg
xRn5Gdo9BQhTQxB+SLyZJuAjsRr3qgvXWlgW/yeU7WHFbYt1LviO9RepfeJQbzz1
fMyTRurbx5i9rjhEbSpnL2SqhOOImOm71tiVl0LDx5gBjkii89HO2/ERcPj38FbM
0vN3u5QRw3QxiihY+fwRqaiSBBD0tlCZnYznULUDGdUtkBIxWQXUEjLamz0t3PsD
mEWElRXFL0jUwhAghkeLANIv/R+F8HuVG6RQaJSvuJTr+xzMN8iB79xvk+e6yVpi
geHXXV9fuMAdhP16TZodfBsKibFSexrqVS4wGHh6RKX7+DpqjWPqovFI7Ur3XXTU
FhfWMoIbvK+y7sbm32dxg7+WZe2JoEtv/I/gVzARAmYtTPMXW+LPUm+lrTrm1QCg
ewrD20zVc2/267JUDJh3TUNyKIzpm//RaZu4IXdihqsHjFTlWepz918QAUmX8WBT
TJ+U22WUbz1WslzNIiTgG9DCbNYQSdkUR200Ar8vw+kMEuCEPnA1VYrHeoIqM+8Q
W9S9oSIa+paDpfD0AGb1mPIbJckPgu8/98qXrRpgUXngqya+fcdiJEzdPKJcimAI
PokRtI2oXN4dO7KjB+7okUM3eQhInqAP8h911CFvqUyeI+aTIp9ZqDOha1JbTQLi
ExkKeMu3F5FXh6ci0rumP7ZGOVbepcjouLVF3STWgPRog8AMfEKI+BFdZrQch835
8DT3QJx9Fjxzoi29CK6ARacuat1G0oSvFvVVBXRB9VOBhLSg9oDFvqjNr2im+TBR
AVB6+243ikPXVfkKNC4klrK+E/utvlqFCEztu2JU2cMuN9lRkzZQJsFg+KA8QJRR
N8ehWGnjge+VZ4lsM+mreSYsxRkrwxOvdFas/ng9n/T/Dc/J3CAojxxnibB8q8F5
fcg6VNVqPwiVpiI4qjZcct/NJfkbifk5BwV67RtGGdDDBbQfaWyGExOysHgr2Ml9
ob9PdxJ9Z6S6ppZO1xcktyp+6dfuznhVEaCsHsQo62mZuZNWtnwqX2qZaByfua5S
3avVeUV2Pp1fxFfL+BKnxYmr1+WbvfbE9CL2RH+uJkYgt72TJS1zfxBpA009MF2a
urFc2CgnYJWKocVzYlY8iKyu8+7lwkjm5yCQKWHDMXTKXVo8aC9NJQ7HnXwFhy6T
Qa6JYnqnngn/gBeMxy0eN1cXb5PKhjoYMGjtXvusdL3hk39EFz/1nezLOfGLz8h2
uN7ZRHgwRr32uhuLSrBfnW0fe0kxzZeZA424B02LQsmk+hSvf9k6YwEFU1ato8ss
eDjwVX7eb1Jd8GvYjaafagj3a5EO1pqCTihGs+XMGUfXdBrmyYupInAx+um36EkE
dJPWwkFQV7qxgG1DztCyjCepzJk4wmmDlKqX1Sj6hp8IDM0UxOlz9DQ4i7UYr/xF
GrfSXYWqvnX7pBkRp+oYUNLfRuBoEyzH3Jlg5YscTvGOu2XnKSQRlt+Y7bxWQHgb
qYe9co4HyRDvyJG4gzQp5Z8aBlM2TxFzSrqSIcl5IrPKx0U4GI0Ws+hqZ2Hxveb5
UaGqNbcruO8t18vXi/BYZYfWn/sl+U5uWG2WoY7O5JF4KnqJSaSlqKbb1uXLVXEI
yKmzLOPmV1wEgveoMosUdmIGI9aF587S/l2cLgrAqL/42eCfazwqys78GU3mvU1A
Wjzt27UqAFf4QEW29IgoW3KRXtRCQOAVNVUiRlRsLV6ITr8WJ7hpMamiXLkkIIj7
+wSKBqwCX/fxLgG6Fjl51GupdFYqvcKKX2EFCiHGbD/1uBoIfWGYATnsKQQ685xo
uhZbooMQpHE235ZC5dYDdhZ+JGe1Ga6qG2S7c/GgJhhKKt0B4C3DJVPgogHywoER
9afIxTd31pJUsFHPbIpvN4pbU9Mgx8NHn6+bkQp68SkNxc4DxAwsyeq93q3yYffB
uJ7QB/yiBt+Lxe7LMp1nnI7ctgwf3i0p9bfLqqbUe31IqkbUdidvj9vYZY0ACLwY
nNqNWnRBUw21tu0jPNR5RxeyVoBYOpQoqhdFONC5rrNK4iyCgUfRuKKL62hmZaOa
tbFfhionb9tNOeEJ/FbRWt0agMVeEs8u/gAhbac6R4f/gQieCQDDvgfBKWhCxUnz
vClBwk+F/mQOEhTGlOa5IePw6e6lYLYgTGhkWTXO4zVK1gjJBUK6HS+ikg4zTGhE
MER0UM04c+yMemd0djO5hB4YdHiig/5mFMb9pJTanTZIyn/ltcwHB4DdJ61xGk0S
bi/13jW2EieMn21tGYQXuinASPK8M55pnNG0+V3c/yC22a9sbwI37bAHsCeYtwF8
2xMxqjagvc8hffuHUBQPmzVgjFF6iznZZYU8bvXWCt8JPKGriJegQgsOfJPqLQg/
loaWoeJANcd0Zt/vS3hdDnUxLl1QIZNEe1zeEzWWs5Fzi1bF1f3PYXtHL8f8P0lg
i1Lio1gQ54bCdIu4o7BeBIUWj3z9//xGA4nh67HJnqPZjIE9pZa/eEiZn0T9pz69
87UXNNPgfm9f6mbivi7tMYqvyoweXs/M2Yl+mSs8jZzuTXi/lOxR5xFqcD5HDyaV
egB+mPG2i6My9FB6xIU9IXypOuJa/oFlNnFuGpfIVpifr5AMcjHuXMXMIxoBuevQ
jH8H6w08+cN3X1nEDRkWpCHcS8Rvga4L8PIMfTl9wJl728WPS42LxCbe4Awl43Zr
sOdpW5fNCf0wUa0ZN0vvF/URKTfodopiPP3rxn3n+mYRAnpodzJHEYF0R8YHYkkr
rRQFT/1Ug6KSlfOporr5c9sTiyZJdmKmfgOOd7tggeVJnfNvd3aFox+S/m40qX9H
PZ+VzdUunQkFAOmJrVqFEtGQBm6ghTv05A0wsLa8GE5qZTVJCrQtNyfj4u1uC1w8
QPyhpm0g1TchR4Bzj+IaDOP+yn9zYIUoN2auVuUSq63YV9LbKdEyBdcstCFkuVKW
o1kxX8QoFxEvlNrKclKtJj0eVFoF0t95PnfQ7VAhPDMeAnlMi9v12fzRjqaBFNNJ
kcLuNVIJehZR5l0qM3eHqtGKQc9k2XsDQddkoJmJrQZRSa8YqeLK+Aos3VgFGQdl
2Y/WC3dSAeJjCFvu0dN3n/N++jszEupYtNp2r6saCpSOrKi415ZbD8AUt0o0opuM
BehIz0QvXIO8jI2Cjgs1mEIHyB7t7+HnrwY7Tp25Ged0OKrur6aKD2WThUyRQXCY
oP9HaKx8ugf8Uj2qgcygcscgLEa9SrbXku0Ktkwu1/KFC/qgTFLSrK3hsm+rAk1K
cFgzWF4N45ePZCG2Kmbci/KnoRyOcO1JnH3iqGwEx3/oyPmnfbFVIrRZzgHH22Gu
ruQ5iREyn9UimZxXLTxSGNFqGzififMB7Cr9ZDsPpTtt44b7ZZUAX9GJBDp/fUyK
SQgynIOg/2DeclYLHEUduLcPv4/BaDi/90Pjz+oG4G2NpsntHbYl3KxhR1YSApF4
PPL0C5zobGj/G5xJQupWTMmM9zjuUG6KbytX9vy7pecxFmvDU0EjpKhCtFqU/IJM
Q/QB2F4keIpK4QfiyQMEoYVwETElWQqYOPuhOJCVY+PNju6lnKIG7utbRnIXibct
2GSZ8OiIRIRq0I8x/ov2p0L1STcI4QAkbaBd5yFo6CmFhG0J8+KOjlLijfgR58fu
7Cws5AWt50mg8I7hdst6YBvI/yHdwyRwNkiD4/HeWZkqCSoOqoPBMWtNCFG2pLti
TK7LM94H80QjBi6x13SrGwGIg0JM2zirj4AeJuAW0HsDQVkbB4JBpSdXjy++RhrA
dsSbwTvA3STJTnH5PxXx3TkOPCkAEVj6nUO/QRdocz3b+bRnT7EU3SM+1MuVMExa
LrptKTIFOq7c8Z9OuUl0IpRAL9y68ZruTLRA1vKxdj7rep8ho+7Bfk2Kx2cXhfCA
tQ7j4g212IoapAeulGB9D/UPK6VzRrg6JbLdomXI5Z7HBjrT0i3BvdwuF8FdBT3S
dL8I2I/P5JIiQ419sHSkECqSxBjs9ftSidwPamYZco+fQkWCi2dQk3ZD32GpTPC0
IPua6C2dIekDI+E0PzKU4Naus6/T0hSZT1WtS5VXKcw3xUgNRr0CyqxIaPlijHXB
VgPxm5Tay/1HeJt1ktyJ5J1wb5sNZ9eFsoN7L8un5DJ67syFEEWcaNSRXvPAorLd
BLlyaaf+rwQ83pRYyQq0BeyRcAeIs/XD2ROC324v/WeDD2+UK/qodgi2OCVPSMc3
SVUS6WwNPQavsvi05EDtD/Kp4Pq8uzAbSy0ZW38Nokf9/bjukLUYAsQP0cjzhijA
NwbmA5t7+lVTeULytUOlf8iwo7CdbgvhntQ9+HUmOiwqOxnd1vkDNjI34Xsop4og
sEInK3HJ/okkdd10jaXpLHrp/Pj0EdQpDQkFBuUfr2j9cXNZJ5zwWVT31JM3v4Qc
d3iWD6Y5Yq0nerFe4+JfH+PS3aRnsI60ouXZ8M4f27txsouWnM5OdoaYTnUz7qgD
AlI8ke7mMYcBX9vXsZI5LQdbIQhYPpkgBQVPLrfOv1f370jooK8rzZkY7gWgsU8A
1v+J4yCaMHb1demiZvALGnBndCop7W3Cqn95v+s6XQF3AMwmqAwDLqwBqCc9T13b
aiYVGSSKZh+L6JEsdCFMEnCMRqRVe7qk7jE9Jj9GPNZx1D1Eg2jdbRmQcg67AUhn
8ITWdnUbcx14ow49mbn2EiU06WM3cvpoYef+F1HzeilMyST7IPv6IS4g2XbTMXK+
kH1RCE70mbTUYxmTQaM/ChV0OG1YjO5CnuR8wt3bSpr20a27i/bjxXgGnZO/ut/E
C1f6PFaXujVcxHjYJ28UQ+WedmixUdMKBGiG+JY9pyZPEgKSoMNc+JttqV9BCBoa
r6fnEvL7JL2l7dDDKSTHYVVJPs9IFS7GakuOK+CJfm147p9mrfufqoteL4O4/tTx
9RK9dqw0QwMojNrNrKK+6RSwgDLwgYty5qlHbqQVe9E9OvGfIhYR+A3+AyuoDXiC
8GNOylfE8/VDFGIuuQviERFQCtWmnX7WfjFNONVdDA9WJx614axW7Qjb8CRGRbR1
cuNqDTFawphGLlOxYa2VUXbIC0d1aEFFhK/lqIQejpULGaVijp5mOqLtFICNXCD0
/8i+CxhQnqr2F98Zp0mPc8735fWdJ9JUlbaJiXod2YKMtXLBJSEVUlvyZEplBWTO
7sLS854Xs2OrJKP2evuQ7MO8lsOMRYKa7ZCo60YAIHLbJjgmXPjFLuXa7vkt2F9g
6S2Fy8MMrw7OuMTpkgvQ4l+L5bbhzmntSX5lcYHBm1o8D6We8H/WQ4sU6c3eEFek
dhNbj0xtphqYNtegKQVRamG6DFd3qKLhZNUS/T6ZOcP8Dh2lelxRiXZ+kaPs0R0i
hUFLjEws7DcU9JeKx8soUsthA+O+vZ4P2pxd5ezZFalUiHFuntBB08P7Q/ZdGwII
u2PMnGs9Li4QZKDmKSPdBdka/A9aRp6h6QKLYgtBF1Tx8VjaJZimU/Uyfw8jVshz
2Q31ZuDSIDRI8CH7ExBJeiGaOYkDDgJeOx69NINvuu6p7Tuu8nCC1xBboua9F8aV
7Oodo9Nu4LxdAXtaZz1ltRZVvYGnDPAJC5dcpbHIKIsrmpQCWOSMY1jxMdXo+bTp
9C65c8i8JEj6bNPZk/JIZk9RYUIMg6a7H36OhecehgEppsrPyRyVC7ELQ/dtKhnj
mBEQlZ8ZdhNb2z6Q2VbXMcjHLww0AbyuQnOLvLC/NiR8duw27/RhJqWnat9o0eM/
jkce4+jRLNvhhm/dskYYZUecAK+pzR6xfXdRjCWe24BGhmIGkGOBz2Bs+57nXzc9
3L5ri5zKpgRmbX/YvVtKfyGKxz/8WB8ADlYaeldUg+l7T78vO3UNcl+ZDFJfTKAI
zz9Jq/TSuEyfEDRK2w8ydlcJMR5e9qTKyGAtvVDJIHFgmM7sdgTgmsQCngfXC7Ij
UfLQbDe/MxsNc+z29VvkaSCNQgjBOJui4GkhxKi4pWXjfKEX8yMpMuEIM/j0PrCb
3aFHMFLlq3Jgq6mbtMLJOg3hkq0JIwL+4zZQsl/jvCAbQA2F9BZpLuim2h9JQVLj
FbFuP7MzvF2bXy9csw3oVdWl5AOHcXYKbLTLAzvAWKVf0wAbi5egzgtp6N9nhaOV
sRvAzRqU0jH5WFjCDe4H5Qt097Ur9WoppWFIStEdWx23opwsbjOg+WtRcMTIbkVk
rxs81VWLa8/uB+nvV7ncpSRUJ4aFJbBzt2uS8AT3fqInXabagdu+Lyxey6ZAb5Xe
LeEnGn7YBMXMyQatT8f3/LWNPD4YYU8bzBgY1bXzx0tB1YfpPbyXZTEYPM9V1hWQ
+dnBDmgMaFiWfol7wkqSKmsgl1DM+ahzvl9OX6WjUlnH3v7fw4SM7WXZXWqorAN0
VjNK68viapHM7aVUsZG6TwVrs55K2r7L5S6XiflrJwaJPR9oPvp+SOcmr6hmu2Jb
QcOT0OOzRtqhzkdi+eAs0iDbYbCYZU/ftb0R2lF28zp0CFDOD/h7wx5I6fEBODJp
IyTGszKRL2evrU0FW/kRd+1O1rTaBn5erIt1hZK/0C2UDK1GlZYxVeITalryEv2L
KITNRF2K9TD6oBdht5xKzerLD0gM36C7tnxwdlJtBrLvT34nR9M2+YKQjXV6Zppe
vqNurrLcncl7GQosqUpd611yymqqKO9FZcYfc+LKxaA01pqKUfbL0okRblJpJ/23
Rd9J16wU/7Efvd0o38QxoOecXFbihbB9ytfpXyxkuLWOKNa14RaozlNVH5pLbOaF
384vck2pgoWdCTNFaV0Xd7cU2ssHYn37JebMlPrqaE3+3wHVN3uIcFHTWkHdrhlS
1d4MyqAUZoWrpM90YHS244wJ6y0DR9Q0aiDolpsbtbxiXzq4CdAWgcOiBe34Rv/C
LUH/0A17yTzvxtc5ig5Hek2dUmTYZw/9yPYBhEu+Rbeb27jvJo1N1Ob4jaudFtG1
h3RD7H/u1p/FgX6m8SaLvMR25/FldqI7RXzbpOOf1QGOO+ix4XhAS7GNyZxHm0Sx
cWJaLz+jDYpUanhBWDe3YQpPm4vre7T3PdX9v3OWgpomc1zyGsyEw97HKNmOoeEP
5cQtB7Rqj2B/G3SVVyGs+TrjmMybOHFK/5PjWZz34AeG2s4D+ohrihgcZz63aiLW
7beaWFzVWbIlfUR1sxTYSaz6iMFKoFSL4j3tChSWNMITAyZ6nvVTMSeDyg+qQviY
Hd+XvVvqP//Je9ORKH7KhP1uC6tHoqNM6dgz/4TVi/yLrmK6I8PXgs0t/NPoaS/S
pjF5+/bhvTOSvm9AGC01ozS+vUEyAPz/Ksv3N1yJfTiCgSMmZVv39rg8M+yH2pmx
I2U+/QznejIB3zkoJrehfvw17D2iNYEyi/953SZcxv90coj5F0jKigIFFAWYziyT
Fx45du9zraokYZLxVKaCHaCq4J7ffPMIxzAbut/XXkVqJjjAqIA9XIWHQcU+q/V1
4Zb3+/q9vz6lBVST41Zu3eVlVs/nw9rMSMw5KKfx0XMmb8Te9JCRl0ama7E6ssA0
u/jD2EkSEgL/cePOcRgb2NnYgdWWyH2pf9CQm2Mbb49MFKsc5fytNv3WzKbvvC+V
Tc4yJtc340FONN8kV7i6chju3MqaNmSqUtYaDtf4zROFUFb1JB7+sFaaHEq5Urje
rxxRM5eB3LPbT9Q2aZ/Xp8Vsq+9K0HOIpQxejZ6IEZGPxWZPqfjzx+y86CpRCQDy
zr9cVp7EZ8TSVvdThEdeVK9yNSOgEn8VeZ2SSrU/HJYfnlve+lM3EKyil0Vx6/GL
x/cRKiVv0ueO/cJHoGkLbeu3njEI90Kyb6c/M7jJnWiHVupUeGke8BQ41t0Isqml
jFaOhvBYdv5JU/MRhwvuQ8vPVBWR7dqyQZM5NU42eA9YMaO9Os22++vz8cukkiin
fE7m4pnqhtjNHphkATYm+MqPyrQjcEjEjFO4zoMix6ONtEwVdDz0FAarFKkFpHF+
OD2PzPKIcLUM6fOQ/lEYDWy/6MeEnwOFmAPjA/QDnG5QtHhcqMX7I8L8OFb3+ZA8
As0GQtvyxJJU6qur7shlB8Wq7fT0f1ZZegg+tEHNUDRe/40VYHY1eEBeENlYUKAt
OdfHQlpYSxq0oJPQ1iTZqslEcGbwDmv0uwNmp3MxEnU0LHVpJWEwnqzrZ4qEUDWD
+t46g91O+afeckSTo6hpd3/tCXaFa/6EDJCV80UA4LdsOjcQtuBWAFGK7V31yfBa
NBlRxiNB0MFg0LYR7wpofxVLZk0DqGAyu2XfHCT8Umw8fjphtf78gvH5h5S8ufAg
5apPaVp87liRsLFn0EDxuaitPtE8jgFZJl+j6pqkdMTI/xugbYf74OSNmOtBgfjy
zgGJBHp5Z2H+iP6mFzXXUCq6d9PpmnHPExIbxlum+XFli9r3gyyjwqDEbhfZ5+OA
oPCyOJ4o+fQlm8IdM84wjiRZvIWorpSI4Bfkus4HO/DXseDtwcVRvH+Pb39BaQO6
iBQIKBI/vtmSG6ql1JVW3yTs7x69Kk+lLCDmwaEpZgTpLbDzcJr30eyRvY2PCvie
IcUMAHJwW61Od+z19T4qGr68nNodZIwhXZp159ROauwO2BQ2jOMCJ/PZ9S9+vGOH
mLR2del8XRCK8qIq6trFJ+OeM2cD+s5v31YuVJSVy2pYc2UmZuu8yMVrRT/mdoVU
F9YZl3j8wSTq+dWHbmXTIazU/bC+ELbxsah5Ao/y+pM8yDRC+SztzZMrOvfylm4e
J9mOhI5muDf/R0ZGIN0WchVT9Fn9LUuut1CnXmYK7i+g3if2g5taADk9HpodSUna
m8fUpoP7PoV7JQ/nlaP6ZXJ5m4pragi4n/Xn4VYso0TqvgPKmc1TyBjyE25DAZIj
wF0qJn4Z8JNuNtKZBKyqdGciZQT4mfa/2GsnCH7CPF+IgAdt5kJ7D9tkZAOpFQgk
PoKUT6Hyh0nJwUeaAS66GdOFKMwdqC5BwFT2gDgZB2WjHPEPBIc8l+5FhtWFWZzc
SABEKY1S+lq8DL4mHuaDWPUn6/3/XE4tjlxErLRbBKfa2v3dpHMEH+KafVPQ+52Q
tF2gW1F8Q0Nk1Vg/axN79/pg76wP2yyC7fHkgF4zsCY93m01zxFpr2N1TxnJnkJv
5yinLabiikMtfnHYCZoMONXmddxl/XgawmvWIU4uyXVaxkrMRwsa9x1CabL0sXog
e7qms/uiWk3Ndm7rDc2i0ccmxBEEwgnfUJlZfBQDSXXZbwbMffsoEIu+yZe6ZZag
cVaH/70ieWXyDyV/cB20PometdN6m23E4RK4WMYf2OYMXkAgF8R2a1wDeQl6YTCn
ikA3f8VAk60cNJ9599GivvQbhxkndnlfN4tjFrnC8aceSG3dlpwlMIlsMyWtkhFF
iasAM7LaqmHPH8HVoBAVOerHXheM1+Nh37EJUN4nffJ4mlv+0LI6Z67smVljHDjI
jga96OBsKN2kMiUw/mWxMIla4VJly31u0eaF7/pm4sMOLqPIVqIbhhQC64YBzgbq
b2j73iX4Ljq+TQa40mpw5k3w/d37jCfuyEnc4BWsFjhoIgc/NwJqvNbTOsHnGXL3
LESAUiQ8sYk6oQsmsSGc0yqVWqJs7VtnNS1qA5xcAp//C4oh9sJ2DGFmG5ozdU1D
Zh9Kd95DBXtgyuajKXX3wP1nXHFSBPeXTgDdgMop1C6Pz+My+LtUGOeDlQeyMjiv
qqmToMvQw1YqZ1BRF2TqN2UQtItq1QvJDoMnfrKa25aXybxvvQmzvjV37W7abscy
BwDQB8jqQaRAS1oLMk+3vbSaT2gSXmpe8W0ARMrkMxK7nvY8EdORpwK9+atEvIvQ
HHOQiDXL/JXIYC4c+xZJj3Imi3zf0Wo8hyIO71H/+1/dO1Hp2kSRuv02R70Y71fJ
SFDtC0DsTI77KstELPbzIovNxVcK9PTDJbP7l/fTX8AEoL3GBfNKl9ey+RyO9z3y
GnceOoebECojCu58Xag6HnLtWMkXYGvvot0NZX2bVP7Evia5IzpgDz9dgd9Wxisk
8E0p45dB3B0buTxWZ3UaTdxJxNd0Ux5K4Xxd9X+HOR8P05RYPvcbadH5+8GmAf0z
G2Y+5uyxaCK/4S1ebpx4SHvuHcN+OXlbMDqzHff2QukOupwLLUAGsBy1Q/tuIoNQ
bNiGLkD01qwH93abwlXlIiqRPwGctgx1zbqNtE1L5pOz2XBH6rDrUy9pJU9S2F5h
Cgrje6n+b7FMTnwxsHOvAFXix2oGBWyp5qgSyAzHWr/wKVULeNhsyi7WyKwqtCv+
5rxQBWmKWXbLR3n+r+xIPztxmYX0KyFXL37na6zm7ZZzIanyYD5ButiLt2uhTQYh
DB/ZdZv+g9k+wGI+6JgaHDU8fBqc+FU6nJsxc4rlA/hawJAYWy7pZ2BxGV3gg8Ix
v/t8wrdWawDTeKmmAcUjjezfUl1LA99KpXFT9HNER/zVuLhEL8rrvmhprmiZ3yzm
KwsyGA9iwAX0Zeh1tse1sTOiQD5q8cU5sveEEZ/CG9073AxruqhiKNB094DpzlZJ
LsjmWC1fZ/7gC7lK01l1TAnXaviToaASV28AY04nGngzOeIM7S6c7qF5A4Ch/JNd
ZorFZBt+qam4RHY0FOotgMRQpmXVSh9qOEfqxj3wAnHivGmczgWz36fPXXBHVGqC
lSEaOgIRnc3mROyU+IyE9fCwYJQ15G4DAOqw52ew3KY1c+LVlpsLrYFA7NVQgu8I
EtKHETBxZ1wQzl/Dgb1/5wJdJOya/sSicx/30ug8LkGjcSt7dxVuI0JdnRH+Pv1r
HqbKaEcCsr+SuMQfwxLn+TfsN/Aj/wfJQOmfaMrvrekpup6+gte7a2yEB0Ik7Nxh
0pDaRtXsEJVQbIm2SuLddityiO6zlSnaJVOgzOWkDGjAPu8laDuXwRpfGAiFTmRu
5ARVXojBrNbZMgdyZuBpzmuyPoYo0+c4Xn8VeWlJLRYoFfmlcNv1ih6Z2HXWm1LP
3p3IjjVDAG4UrAeFuGEKUdyPMxhp9dPIxWlL/5ijqiLqBMUHjA3Nuhpr5GfVst1p
+x+gtLxWA8OEDR8LNcKdSi42H4sy+OC2NvD/69QtBhmjHGeo2ut9qpi6BQQmkh7F
LeD6yci+H0D3CW1l25CpwiLkj/ZO8R9M1S9tQVOpzFpo5B1xgng/2Syl/hSGMDgK
BP/VM/rjpVFGQ9Xnxb0pUGIo16I2In8f2YV1dIQYfI2xqhtHLlCs+nMH4SIfl+Df
DzoOnlqturpFYamRacYxWUefErfbM7ATpFfK8XxSLBpEYo5QufQsNpaat/g9tWJR
svxlEb7D2cAZayxkFfn9G5L63XPyfieBNZlpEN2mBzqsFyL6Te329GzGyh6+Zfpy
+6J1hEOogI5Dte/h/gD6RxuG5KIIH9mgRNjccDCqJLY01Vk8VgZdsnf6RSKyYbNE
CcMwsjS5NgkyB2j+hxBjwTplTDwYvOiADJkoV7G8WTSovmR1KZk0Y9nVUzZbVCkB
NAN1rHAG8JEkVd/LnGKxYqZcuVvvRySerWAQskMkGGFkU2AjQLdKUu1/3dPGd+Xx
sZ/hKhPUG46nam4Wx9mIgB5GMAj3Sfe/Tk8U6tlcquGPj9K8oEBJBhXN+syhWGzd
d4uTPzJdH4Mqo+c2uKUhEWCwcNNgXNUzS4JUz2RMF3xNYsbmveLg41wK4y72kyAF
va0H3488/lISbRZbmwjPga5B7GWcsdbqlkRaGaRdzF8tVI+dGbIlO3dNUYSk7Ez/
R33dy7pJ8CDjNBcswRMy5o1h9XL25r1N3i5bhWgZ2llxKm5aFi9CYlI2+ZIXDK+V
I+uTBgF6+p1O6oMXppdL3y7pHn2xLcKj1KF3Xtd7FkOvOrXSxwFXYl7YGWNCnBXV
rM4/2NyBKiQVdVcpKHlBj81cUJdWzVtnP1BqgOZMhY+JnpsXtGYc5CiY+puibkrp
QVODYv6dBG4F0mGLZzd3Z4VCmqGVRsMYg9zXn5nCPpXpesoKDpZLvHZy8LXt8Zka
Gyk0Fbl8LVKJi0LBpQ/7lgTt3eCaUvTWjekEL+IPTM5YrkSExb/fOkiIaYH95tTL
IfcisIxBAecmQGaw8hn36km+x99rabQWOAJJ/BJxraXrWzyDfjRkEUAYMJKoXLal
0Zode8PxEm8AqE0Q5jmztwX7Sn9q+B8dMbfOtPV01nFosgpYE8NxRYdkrVMmJu+/
PlDQpQNrKd9YPS2Qzi/ry5tQwTp0ttEZKH4H5Ockid0thojLH7ddHiGYEsrt0/wr
yh4HGYIAB6PNsN2+UM/qSJwD0EVbOJqM86ZNudwb7eN1Oi6R0oCW9hHd9u5/BSTg
9yuzuRHRBfaR8Yh52K3MW62CaKmUBUPFbJnb8/5ugrYWzXePix0nz/yZc+aLdgOW
V3i8WB0JTOCyMcnUX3lR9oJLhHOciL4x+NhJmGvcYTP9qn1RyNhO9tP4IRSgDdIT
Bmt1sG3JTxZq/QVrE1jp1DKzPii3jCGDiolaq7w4n1rPjmbwH0PSJh7cRzFS4wIi
r7YG0rVT8EUFHeN/UBRLK7g4dsUz5zGXLNhF0N2/9LDGDR/kStIlBzEX4Elmouly
W4wMiu7xpH4cBVL5otAazd0eF3BtM73VXEde0VWfwuh9zgQ45TMwIOYPJ7NnzT+4
FtI623ZTQLRprrFU1iGH4Q+MSO+IF4kLODfbMxmYQ7i+j7k9BiE0JN0Nr/aHaPbR
2bj6CQOpROzmzkvX+1+ET0ZUjqsKLlkh98IT7vUjAXFdIztqOJk5uCYvOwr8j4L/
86Y2Y+u8y7E/BFEihNj8IQFKkOwxuqB036nAE1h/CFn3tDsuCfkT1dpOd5SdEVuK
x6P0XRz+PxATIem0Qe5EBTa+i8CTA6zqeLx2KMg+S/cINZeR0l7KMOEeCm/lBiDZ
XCOjwzLPbvnoYhRKPwyAhj7mKJIwHxXUgxkKDEynFiLtOtHigpK7yp/NYHMrlTE6
cp+hFdVxPr+4wjhEROOP6DlTotBKCXvheqPBotGVgoSAnk/kHWDm9vKemOFK9rC9
IjVfv8lL8lnTSDsM2qMtTVpjT297Bt2cRe2BXd460Wh0KBJ8SUfe1VsyT/ghnAmb
F8ebgYw2y0jbEj5QSmeSH0r/dbljY77nHUGNHdal680kKJ6CAY/1/5oUxCrZHgA2
Iian0fSerw7Q+PIiOFWcBckgozmP5mSQm7YDHtYXJY6MK0ytMU7zKTr3VneKe/bn
anzggGJSrPjXFPYQmMp1dUN3AE073hd4ZplKdARgnwQV6pS3AGheNcFHbeKO0GRu
89+OgjJE8N2W72kXuzpTihtJw3QRYkjoyv9rTV1Z12+9XAY+Tzv4QiK3TpPs+sYq
CndW4AK4gqa06+7ESrAK38hp0YvGBOgON4FezGrbeVXfybqUxu2otgQyW1XnmOVw
abOzNOGwxrXyiEjaHjxtUBGR7DGf5vILTrE6enpa1KMbNEYLpg13uV1vk6kig4og
CI4v1zHQtEz5TZ7wq5UUMsauYPV9FUFHeVLAJ3w4HRrFLhNg12Ow6E3xonqpA1sS
b1dM6tFGykFnQcpR3Xzp8SspzJq8BD+cBzE7j6kHd/p5SqS2ne8gwau6ni5DgG6Y
bn5B5P/nF06u7MgomcNYpJDCyhMjCwuHpjpAVnpYiiN1JUQYyw+iBuRKIyatUEZL
PMfC8lx6aRYMlSJ3mJiIK0uivM7QWKAjtSL/feVsKocA6AlA0yoycSrYW4XQP3Le
QsYO5PIPbiZFzq8Wv3p/DMNmyD7RbabJxo9ApbtF30vZi1VTntqGaLqO1D5NXbhU
6p9ToPpC/jPQwSMFmlIDcPkUAR+ql0lxM9wzdqtj6iwm8ZZ85wlxICS1bpgKpGoa
SsywjFDVkTzOxsbFzybqwtDwjVBeEsOR2dyq56ka1aIe0X4RaCR/TQMhaDGrI10c
qWTDUSLPPAF6kPN3FyQgGL/37M8TGLkmldYXg/s8EhC0V6sRIT91H90tfWI7AQjk
Libooun++sV8DPCy1z9+DzJiyWaycSgD+7uqGrCrzFuoOgzEQdPjBnvVq+cHVmjx
7M2FjeIGRCIf/63f7JM+M7lPwMZgIyTrTlH6v/up3rM8CnS4ffPaIEzIPOeVMLwW
aVHeP1mE7cpjuJX8ukaNBkK7KL8MUrg2yYQPj5OoMCGhB1FXZ02vKw454XVwPf5t
xOPcuOWFxNSoBmdNpqLzbJM7T2EqTWqeJpBtudF97geNMEhtrxbZdwIZ+5IbJvYu
HhGWpq9hTpleAtcmkCUwMv8jlaW+evYK83AsBT0EgLTJxMD/1oo9xlmZ2z5cKlGp
lJrn3+oWLKsaPnSSXGs1ZIjKjTaD3Wq5FJ7ZGExybWO0nugyoDdNSN66AW91X15i
9snr161Zi7JPn4ipN1hpDiPbV+CnAJok+WuPufDldICEFB2H4fzEKFpM9iJB3PQf
XcDK0OL3Qh2XrrPjKO46FT1V4NNGJySDG4hp7fTesKCl/Ge6sFdv8j3gug1cpvgu
S/Bp0QhjQh+zn1x0KclUNcboPAcyp5yqXFqWNpoe1sI3R3xYwPCt8C4fIhyTXJD4
qSw4Lr7ftpqJJeehkwVORPp/rzj5TKVsqpxvDA7+2+HuA4/tyasXPbaQiP3POumO
6CikgHFZXi/0WAhmQkeKJfsc7HiNSlqNaddOPjTXSWK5be1yIr9yMGm4570SFRbp
PZVVoZ7Nv5aXFh9LJwehWrgc5PMtQ2ClXvTnDwZNZuF9m8P8kOtvcAKKHj/v7Tly
xm4WynTeprmKm+D9Ob3w/RbgzRK/Y8xkr4erWp308SGYzIXQaU4f6+t6Zjs5WMYD
vtyaxoH2+SJ17CYl6McJNfsLt3fizp5BFJ+oOPbdkYcvhwTf/E+4oNS+lV+0iJRZ
p7q6An6FcXbwPax8gQ1LdnYZKFcKlrX4LHKJi5eYJXaogICV9jtsI0IMaKqCDG5v
kFqEJxkVLJE5PWNjtAL5I2nZxikQ5W+SLMIUsVyjqePXmKwo07LWLTaA21ERbhvN
nTatP6smzbm+GXIsQdca8pI+t1/GlSHyDIVBP3/OqNfQJg+zpj8b2vhnwksnO1y3
FMUv9tOLeeVsVFjQmpzF7k/4aogsy+QVh6WyBdmFyo8NWLaBjXMttltNKVP2quUf
2R24vpYnj18O8uyfHrUn+HtE8d+ZiGa5Gnh0QeMcSfIVCFDquRxn+t8nU5OHThHH
eCKoKTeyA8/EL0mD/nXE/Y8Ya4FqYEQqVNwkl9QhE/VSEl/S5NAwW1Bfa59Sffjn
wVBI71ttksh3062hPXaxkPtVs1AvbadYk0qR8Oug2peP35MXBm2Guk0e2a+rLNOA
dexonZW5TLZFuCp1xBA0aqos5lg2HU17FyBswkYlHx6DiEHNOrm62mjtuC6XR4o4
BGuHRL29LgKdIOpy5Sgg3i+my6K5XrHAN5sKFP3Y8XDD5fXsenlefAkM69jJfPQB
97UhUdhyFKqzDdTgBjObKFNslQveybRfzZ1IEBPplWI8M79zyvG4VnEfTTgyWVQr
sLeGynOhaNDehu8RifRVAiFpVvCfgphqgd6KspluVC1eAUk1nJ99hjSlyHgqH1LW
Cfxf2rRnJyblmdwoU0hH0G3VBonb0W/txtVw533XLaVsixKrKWVSFygLCliy1Md+
OJ7dw92+ZkU3gBlbPK8lm4ltr0EAuAhVQWWEMbkf9yHaKSkbX85DH70+94TBkjKl
arssA9y2tfFJ8NcMngwnSFJV9gcwtHbmjzW7vQTogGTI60ROYH8YuPr1DwIu9+/k
2tl4yd/wTKymYXBOOGXIFOMJGeKbPvE2fYTEz6YJuobhoTRsBxjZ8INWYkoX2bHy
6/QzFizHnTjrFqp6LSgWY8HOlqGHd1fePxifg1jiNObqVwzXwlSPdPZ5xXciy5yB
5zeQFTYrIzd5u0kpku0iypJ4GtujGhXhQPEnspGQMjp0FoNhzgt5rrG8ag2jahqc
hQo/t/9BXPh8Ug/7rn4VAKEOK9IyL2hsvf9kad9j1GurshkKdAvMoMTshZGo316b
JryLbFszbkLHypPUlSIQpdrkvBQ0m3ajrXuDavlMnm35vzfnlJVDZK5Yq+U1qCiY
Lvco59N6siEX1ZJJEpKQMZrJQDP5gvqm3kUt9msaidjGv7bDqYzuTysF7xYoJ3Nr
AAjhjnkuq11PwAsAkO0r2gN6G7UPcF1Z1ZISfUZrk4XzlS0vNq8Y8YqGXbz6ymRF
h3L804wEhsGmnBDilUKI+PXbl18+R7w3BdOAI8o2AnL0tdNY0YYWHsQX6WusrA6x
UpbV22nIKJatHFys8hLCv9+EEi/3dR9K91GfKZmUgmwhnR4q7t///i4FdDxQ7Bow
CHMXuF97t1OxPu1NYgJ9djrTOM5MfmvCMsBHZb5PTe9UG7TEfUzo72TA4JzfTyD8
KzieyRDKrCnDXkOFh6FJt9Oqq7IV/4ONSdc9drFNhUgOFED86NFlINGXvhkeat8h
yzCXmmXpTumSqY3HqDvkUqmHcKah7zxzWUMRoRZ2VKrD0vRTxK8jz2vGO+0w4It+
XXku3rQKl6qWIMaDYIabjY3jOqbmMGfsSuNLmKh4oTbn7oG0eCpUKKnxN7PGF1+y
w0eMo8btWs6qxtFueK7wnqZVR/+JZkR0CbjAqC2W4JsdSCCvdrsYLHRu1zlCDa1n
PQB+p0qKUmJCritDBU+NE4WcH7h8rSCNkV3/fT7EMTkWwosGf4Tp9iPuQiiIqLCd
dPoT6r8z31eDtsPbsLDIQLw3UOcAD6hyphgAMO38vsbb8CqZs8yzeqGhTE/kpUnw
DOzwBMBNtvTWpLSvnTf6xE/CJMwmNWe6vlO/cecVojcmB+TGH9WDXq22aWWOUOD7
ojtNOO5TtROCXc7syAUJ63Ep3myBywOJ4W/fI+OCru3qNZReF84GuJZjbqXA5f30
X9TOHCAbx687HIyZUq8TFBS7scfVUE63fKrFl+r1JGwY9lw/sPqV3IF3TmeDynRj
7/5VE7AYWGfFcV9q6/hjaGg5TdCRM1bseIA9rgaUdWflzu98bImwyS4cg4232nbP
3s96OeqzJcz6XP17kpHdmCw13ZzrxMbk1NSeMgRdaE4KBJLxM9wbiD4yvyYLlTXR
isTCAotf6qq6tG4Eo3StWQ0u3veEaxazL2XDxsiXPtDRK/ANLcvSFQn8+d56aFUe
hDNFPlmCaQX/l2mX1YOwwReYbeNmdefdkyosOU/9aVa5XSqX/CjlHOZCvMGQFANY
vVLiDASee73yXcgwtt2VZrDCK0koLOJOaLh6ZskBcNiRvQ7cTWP5MefVWPAw9rlC
YozyEwvqrcDoNHIkVEB8Cdzx7t64T35e5x+4mVQVofh9gMiXMruGYQ0eomLhxMC4
GuSdIWpFrnsrSLbcVSZazgEJ2NETp9Uh+Hy8knW20uhAJ9w6pcKHJUeaJRPZQDC0
wYvjEeUzYM4g7T3FuE0oD7riijyi/nljC8xp9Hy9gIuVDXc5FmfKZ5ckbQo4MTXA
v8S6RKc1jV6wvm8n2glONOGrdclMRjdN+pPXhii0Onif6tmSKnFJ9X9men4RjaoO
Myggv2kNQ1Ncbr/fmQCrW7QA8WZTt4BJcFXxEsqf7D8KI8mSGDRaT01xwTTcvjEt
wxL55SAPbybF9oujPkIGXtS2/F7hxuLnsRHznSaghgER+0bHihEpGGI9QsVbD6PW
mTOyowIqjkxhLlJIsF/qJ4gbLSFov3GrgBBxIk+Pl8dBRx+XXTcPyzZPVMbyu4rD
f+JeXb18hOguO89qql0cLaDNADQ/VtFWHFiOlDMmtevB6r27+gdAwx721jE7f8RE
gjY9rjYS6e7U73R5ugsHE5xac5gD4TqbrSORg4AUMCdznHus8lCZE8wQsfxg7Mtg
+YK3eGHEDbiPGCfKuebou/5BDP81Y8ALVAyDq/lOPujuns2GHnEzZ/EuxibNODXA
Nqd4C2/OCAKlQIxkEjFoJVOGSISQER/y/IutEa9uGVd8iAspWO/qevyNS5PzUTfB
Uxc4zZDHuaGZ0sIuX0jo0mzFM4e6NcZ4lyjPEH978edpSNVJRWPjWz8C75DVnbkc
ruGYxV2d1v7jNz3S6oYajvODgwsLv1zBxBJXk+4jhHRcjocWRk28GFiP6Xb2mz0Y
IJ6HWDIA5dB3QUPWfwyOIwvmQaybAWZf5UP7Aw0aC/wavUjJtSPnmlxSBoEu8QcC
FDfVeEUh1KbIHz8ZvTnk+eeyS97fiDYdhxmKJn5cNS4X0LVEDXEH1yN3gm0q3FMm
rGVhKtMwMPzC1mm7QreHADmQzhg+cIZv8G++ujxcBQY1XbsDrzXcCn2jhMUPCvre
E6ATMYKQQIvtyKm1qWz78BG9BjUQk96Rfo/sPFrLvoR6jUirqEZEzSsR02rV1oJN
NL6hzTwNa/l6kglYPwGj/uo70HH6kNbApsgcaTdLiYydGHYmXQ9tyoq9OD9HnfPD
qFBJCdpisJh6JCVzJvNcHmcnicwcytBVOkPQCK/zuSW6TT7l7WkHNYmqMXCKyUr8
xp+9udU6Rx54Fwc7j1nLso88h5wGRtdpbGoT/bLmbMcCM+ruOAxIhJw3sLiInvlT
mUXB33mHZXDZVbyOlNd5xyW6cpv4e+pD79YBHLGvvoKRD8EXKqV6QAkQKT0RpqTT
ALYiF01hUqvWtUORj2cgcsG7jae5FFRybKwhoOTMA6lZVQ1nCPXj5vxbk76nn2T/
tqYvJoMP6u+jNvdV6HN3sDAWumq0q8ljgrZz5HoQALvbGG06DlCESiFnT25qnYoZ
uCpHQovKYwI+2CVIJdtJLt5WvLgiufESKeRIaFfT09lYmAqZv9g5Z432dW8+HD/b
71hBkasj05rts1pUCaIIDN4l6xYmWOeNK2teye08DUXm6iEDeOLRb4cp8kdgyYNU
6hYlv4lkP/CCosSLzEsol6BsV9pC3S7iOizDzAcxrL+D+c+klJvLrJHM1wlkW9h2
fFxV8Wu7CJ3tzZKcL8EwrHyC7itadKKmjF2pUWnH2ADnfRh8wzJDMusSSUjNhvon
2GyCzWOYhT5q9+3HE7GxywI3afASz+xY00hhq7HLvKJvnyvfytB1o4A29aabj6IP
kn/mvPTGB0iSo2Yo2RCTpFJNGP4XlOoe9br5utqDH1ZLrSh4w/W+KZObQRQHFrcf
2/sO6AA9TQfYYBvh7FxW1UyT5WH3OPSNMAEojWjFx/WMqpTu9CgQfbsI4dpxi9Ua
nYKKTfWrarkMoUxPcpEQsdbr51ccvh+yh9kK/G2L2+Kz1qVlIt2ROtYG//Ew4DlK
sgWEJZFLKOwpCKWaRdMg/0memnq/ojeYlfa/WB2hYzrsIfSURqX8WXM1hyExkgUM
8g4/meLkUyfLQPZ4/aoe+tPVibREodcGEWT1tCEAIo/gHNfvujiBbTy3fruKp8cB
bjwNanDuLubxK182tCYSOgH3N3tBkESlQABEPtes+JKW+MKJA54celUaljbQtYYt
W/3F5jtuKn+zCNUiflio7GOXYBzaQOz/KkOCf8D0y4m6sVsG0749MXQsSxURqgDI
ld0Zq4fLzx+8xfMmndgGdQpAVM7M999tmxFkmC0ZW3pKj6xZDUlakLhrx4Hs9J1e
pBGpWF5j5L4il0dFVVL8CPfyAw/7C9yI9J9PKpMYpP9uCVuYMLpElIYZOFs0+fRs
rOtdf4GbgnwoL8bx6teLCj1+VNxqhVdScFkAtQBiWR2IsP2ydcJFE7Jk2G257vMp
3PcIeF/mx0neQqlCix59Kk068zbAPlOu8sfK25IKVZX1IF5AL4ld5LUr0YtK5w2H
wgFfwnUz9n5MybpjOwkTZoPQsssPPgeRGGzsbcN0bUcUYMPN9m54e0wPpbU30cuw
ecAZ17h59ppuIhUTDjcwMTDX/oDI5sqVDYTkyghqlV1XiP5v4Q52r7+oCJbfU3+9
F9h4P9HSvpNM9h+II1VTeWECiWlMXssupFwebH/QMua5dJp02Wh8++Nn8aLNpqSm
fqwtZHbS+rM59rTLwBUqXtrxii0T01h4zFFVyBpy2VyvWaJn3bTyZvN46Rxuuvox
0DFs7XNe2d9+jV4FadYF5bErzH0OXxU0+ty559fbWXyNhFpVz/Bvx3lx88GUuMZf
7ZWDNip1Iu3LBByfkbL0sobzk31CDhkDM4DZiERYC4dKXCThOJ8QH32Wf/jmNHo0
MqVYLCWyx/+c3osyz75KsM0r9q1tt4/Zx/PCFAkYaGKOqyw3JdpU22x0zOHNNyy8
lFUuASn3QMO2BvPN3COZ3/1mTBWkQubXOioF0N7arVfh5CYHqS74lQCIVbgUqtfQ
Ixo3iiAK/4YXORvqIYnCl/XoN+8dmtzztCDSSgeWchBBMC6nndMlCL+lax+KgB58
SS56k6c/eLjsZgL5G/qRmL3TEewgn0ShSAiwq/xhpGB6Ar6+GLMVz16X0Vbf5tDX
9fhsjureKj6P8YMDhwjrmofUIWPXm/41LPFKYNx3J0yNbpuzArCtSbgjbAoNZ2AF
4krbsbPTbSk4Yapvnx4fREU9wwjki012tMzYcUDdTkKtdpK3WJtFfS/HyBcMYCFT
a7yo9KljFhZuuLIVaDQjOisCJjs9AzuDEOxN0dzFk8wiHOTkL4QlKiEvIfXJ1lj7
f7OLWGhD5YGwDvmqN9dT5pvjftFLXC8UATmg0lM+uZoduZARsWdxH796HK5ROAUm
4F2lqNmvfWDYz55tiCbSCsOwXd3wI8nfMV/vOsVb0RD0tTP2Wu2y7fgU1BdMWhVS
zFYahMcUMm/k92Oe645KchGvxY/5W7Fzt5ZwUZWatPPTIv117LjcfRSXoBTo1tXl
Phj4dALrg0RB6qtrZXNLEGLUSGkFXZgpcV9Ju8/1WaWgfvOCF29Jlj+7hKhjbcco
5IDrsUFykSNdEIg6oAW3F59lrIc9lkBn8bQQyBM6/VqsttEDpacAwrqDb4y9eeVH
rT1YdHsdb3HqB2zG8EsU/nc0WL16OqcGYO0LZszw3zSaBf2HzsLiaunm5l6TkmGC
g83J3nWQnRESJngUG+qKS+iGj4Eyf2WYMNT1zNnXIR36oet5JF9QJGP8BYUm4n8X
cgiMPn7KqmLGMDXXsHZZc+TzF+I9dSj3WeVDxIJCSAzkd9fTWTFe3efJAv/ociR3
bdJjPjOievvINDq8F8Lrb6W3QQx97v7495ZQ81jXSHvFOhkacRXvRmzyEBIxcjik
8BICuDfHcWPZUWCyAsuLWKgH5J8mL0Yn6QQQNSvr+TO+nr+a6/arfuWHNPEHB4qa
OYIn53wTiGg9WLrLviv3Mu5MhMr3QpkA5IvURLMcPccfMMdckF14cclXYuQF6Kro
e+tp3o2GbezEphRc7QdjYwoaQJGCpIU8704ATsXYOORu3kt3D3h/5PWVqlkyER8h
MtU5H3kuPRZp1VoM2hkubrqo7M9v9fkWsr8Cts1aAnbtBPPNhHi7wUkgX6VaQMju
eshDCadCCvtheHzZK0gEeuwVkc78Etj8uDYyPhodTG9OeBqnO4EPAWPuC+XtfnIM
gRTak206T3HQQqdQr90ibpaDsh7/inqzPaVbk7BSD16lcS7bvd2fUtTuAetSaBG+
fAMl9Fy8lyRhtsgMQMzcfHK6mnqCMSiF+y38PJcW7Rb1KorWHAZhAS6jd6pYTXE7
ptkjsHHrWujLwU41mX2i78B0imXPBEZB6pN7IP8IVL8BTueA1HwPkLC9f4X7w8gb
0odinMydbO9PciPZM8fNihaTjpnVn2+hknMQh9zpk7vQzACAatqJ1aqkjnIJokHY
3GEeaW+Y4J1UFr77ru05xnxpbO8vnMgIHFoo+nqH0qZgq+BVfDG5hvm1UMunr1lD
DUYjnYd90mulmZS+ViNyPOntnbPRcejqj8logZASGuSdvgzypwZXTfpbuBaattMq
6Wm0BvqLpOFZLL0xpPUNWhNs8+w7dqo0tD/sBKuKBpzoBWv4gptGZzJfK4usbZ62
NVOQJdXTHR/EtR+Suqeq96cT+rMgg/icWPY7MC6x9jjmqllHW59qmUPM6nAXEw0S
fLhc/yYHsO4NsOa9fDJ8VFGbvBGP79h65IRwUmtTeS4avEg/IClG/Z+RFwkJuSWh
R88BNW5X8RFXrzJg16lm1pj1Q2Z/Ay10md4aIEju/CK+E6JBFKE4H+soS4H9Q7fP
gZoO2z/If6fH18Q7QAmWewyGNv3Y8+IlOZ/CsOkj7//MXYUcvZVZ4ZPdbKzFVFJO
w20t9i4sjwhm73aax4hrAVaDxzPJW0cPH2/Vtz1rUJglNfoV9gjOil04QBIWlO7Z
LW+djgk7HeV629Cy3z69ZQsEqI5tpm+b4B51qdqU4nLyZF0YTDuoXrPhncWLjlBp
lmGcHVdqVF131ryCYXNP9vs8gp7naRtXSakCQzg5xFNsE1Wx8J3iXD77cSSW7mhL
kpclNwaLDbKXVKk7nLN0TlQbx6N9yNVScbZTG2mN++wo3Bu6gHvIrlq1pep/obc0
FjiAjL0Gt6tSarkXa65QaIduJFdVjWlr1TDU8epSTkOChDCdREG/mUroke4NfIsv
JLpu9yqMqQtZRWEDnXwlrp3zY7X5T8WenzWa/iF03zJyJKCxtmSofPpVmWTSL9Y1
1eYKaYl7QmBpNXX3rGu43X/ZLOQbKBoPNCNWP54RmQ1v4mZuMPh/oofOcyzMBF+Y
3HG7juLUxHoTmCA31rW3KW6NjZr6v2JNHKYvfaGPfZulOB8XG3I8cPWHmNrXicrj
C1UEFqDXmHKZeXBk3y7RFkq0Y8FNX5vh48EFbTLqoP5CFL1hz5SI7RvR4fTYBMMM
kC1h6mDYGxvYOXX8pPDi6sCllzKOpcdNHpdirUNWD93ZcsubnNmO+rwtaRf7yxkf
1AWkEMO830VNAmT0R5jrKAEMWdbJktWFKrZlZ2YfGd/k3+mKL9np1ZK7GAcGtYVh
XapHMkeVazNrOLVXLncNt7jxoNfAK/SJSwh3kHfnOIfn6KlsWPsJf6pNmPz/aHoj
+lAmuX1apryoZrpZ9a/4l0bEoBQeIqQTFTa2uuds0kZcLRs/LmRIQ9vybmkM+uqp
otYrhqYECqRPrXMl3rlPX3UhoHNVrnqsu4VFCiz+bh9kdRi3W1Pxt9tUCa1QTSZM
tPA/aWoqmWRW0JVKclp8njxGfkDr83ez0HXn15/RtW+hsMbZn4xMpP0gYM2d+Tux
5QLFLGdq/hVV5qGVDYpoUUAwmQUldDgAukTXHlQOaVC3e4GCFwAr/GLy9pa7ktwJ
fmpaEH3vP4SDS0v08OAJF2znREZxsvZsFAnhrXBAJRW17BQKyb4fTGQiZzDKfhyc
qT2BheqgFbeFq1Wdo0d1xm4oUgC3CxjE+uOuIX7gc8btVKN9qHDMcE7hlDtaExSH
WdpTxps454wbM2Bi7WHXht07OHylqUb0IiCrPUqeq7BTFjoSDAgmg5rP44ZobG9b
GB/riXTQxUwu5QDWJC2dtIzxMZaf7BN7+rqUaq898J4GPiklW4NvRJb3olkE7gRG
KXZBfG/IQEB1HAyRy7MBpOr3c3Mlhd8gRf9hE7XfOAMl01dGW8AcWCw3+3zPPWY4
2UDmDV/nUIBfAqJvII6f2RUVYPDumEJz6rSuxy+kQ998pgt1go6/BKZeapblxOHX
I4aBzhMXJ20x+TuFECiYu32HrDi5vvj2wdS+rlQzxkJM7JpQv1BjVyFaRYyovd7D
0qa50HrIMICxakhTpZEfCPCtwHOsomlXw8fs9w5XZWl1jXicKO5HbxwujmwxcGD+
57jXIEyMpOQS+inFMZ7c2As7KYjy1KVjE70Z4Ggv+y9aeklKkDby+714hrzG9wVG
eFXkwq78TEqCKuFh0P0KccRdyS8Fe1v28kPEYti273i9zlWLwFW60o4D5k/0IQox
FYfoGIcx1aDUrIoAmFkqDYunZly1VD1QpJuIEo3vJ8QDhOrgNn6pnCpg0xjrRSs2
LXzjGtoqeWhe6B1kyz4jagQ9W7aEzTvjRJc+XRWziMK7R/GB3fnR8UH5z4CofuLg
QDgPsxfNp6pPvRePqwVInBA8KrBo40fG78CYWYfvrkdYhHxZIE8gHnncKq9n48uT
wjzTW0/PpNcFMqheLIgGASP12xTWAmKZtr+ROQnnFaY+qWzga+E8kMKPBJ8u/fj/
cgAon2ZVffjkOiPELOhdG3sFrVKswUtLbUieOp6Bxm+d9e0yWpJcHGJrTnrDFEMD
o2WRgdX1Nv5mUPD7z8QSC5dotaQJfcaNgOJwD3jQZeEWbNhq9nb7jvD1ec5MAkP1
sz6l28Z5tPle7UfyYfIMZIeGU8o0/wk7oAfFbTDXG8v5qFkDp7WHzma0Yjn8oIl4
m8w+aW7YXzA0R/7vJiWH/t0h3g+VMFTjFu8iJ+27vM7844GC/U2eAf0Wda0vXmw7
nleBSRHlwQTTzGR7UgSIrBlvbnQADzrBHXVP+EM46w8XW3sbg7cylBQtxAjJFxwC
O+gNP76f+hfz1tFwVsb1hLa7TL02MkbwF43lTppjQ/1RYJHmMTLLe0U3eAEFLwbe
mZWpNGL/1cw9V0Imo4yxqelJ31JXTnRtT6FSowwQvsb4cgrIyfBUQGOZfjKTcvq4
FapIAStkbuG1H++s8mqefC99/5sYK74J25pC+xSuE7UyOBhvt5ssf39Sx2vXDGC/
HSI0iu73t92hq6Ep+6cwlP7vPsWvxCGmcQzWVDVQqvv/H/Xr5GP9SGoKNdnHPcfi
FrZwZNSB5dnQJtu0TngeQ7d6xHBsVogY1Lx42amF7SRU+6+OIg/DZm1nnrDYffv7
vPSwMEX6hJhzVEr6bI1ydPLnU6ugVZ5B27Pr4lDln+ajGtgoyPKDwyiAbEMQgocR
rZxDss7bRiN45sEqfcequY/rqRMK78cDeQn2vZf4QjchBE1fSXnMoDlmcY2WT5ds
V+ecoUOx1wgVHr/PJ1InCUxUyVXLy/xhOj1Umy0NtJQAncQ98mvVBSQZG8G7BlW0
kSqMxc7bx8/JIem5wBwLpfPk29bgr2cXOLGVVhvV1b703vODHnp5eg0v6SBkkJDW
VKbfYRsrsXGt/uFf4lAEMBlUW68hsmpDX5AbZBlXa3mQ/C3HtyTSUcXonORpzUxq
sfCMknVUNxpEcKI20kmk3QYpsxqm9lH+1Oe2+yRM0wYjFUmSOm7jOOrTgyWt2h7m
2tXfFJUI4R2cO/CV7r8vtcERjJJFAQnGpg9X6hbeDNqxrxvVgo3KAqe4jV3MJ5Zq
tkk0oceJJdfH74kewdoJpB36gfK+I0FM5Zg029hEsoRfE9VptL10jBb0ApxM+9US
cFGVcyS0gy5cYgGF+9ogy5EWnE8AjMPWUT/toeznmwaoPUMJsjdY5g1RqicsFZzL
uKEPVLYdaHxO/YU7eTvdvpAxb4mdsRY5ZlL4GuHlSXjZvfYA+xE2F2Nftlb6f9bW
66LpWVKhAgaX+vq6UBRwandXyKPiRLgxyc8xIljsNvAlzgfVmeIhE/jl+/Sv1kNG
CCu9U8hDwU4B4Wld/aRVCAq5L+C29tviQFZmeyP+VU2glfqeOyyv9/gdXYtVC6sq
Tui3CvOsDs7L8/klDLH4GwpK2bBMMOnZyaT3HUmFvw4280NwEffo9idj41IkX/dc
vegMMzyjsk58gMHhhNc68HBAfTtA6sP3Yg3BbNuqRaZY6K73t5Gz/j0tp+6wOPpK
Hyx2UZBoJDBbffDOaWwrhMO3BMckUrZaGDf6gHQsrOuXoV67zsBDYMCwuo+Glm6B
GHnzKQs46yh1o96n8wfMBEYmnaiSeWcDoEEEanKyNVTvXGCQfwiqUMiL2wAQbBZ7
T/bvY7lonvbe4hZcEUoA4mG8AbxKL9eTmbgMU4oDyCL0xz5eNQIm0BtnCPY4tsLU
K1/I6kn60V6HzO+2YQLObBOMx7rtJFEgLQ/pJngTgck7jWldOuRwmGWWiBwgXWjL
8Qw6+xhgYkUJjcJi/guT5IaI7kCLsMjTNxTmzJiCxwH6nquDtjNzA5yQIMJeoo6Q
weV72VGG6P9XhajY1KhYcEtVoH/EURF+xi++Ngud9RR89aY5Wq/GOyR1oyyczmfp
IL+xdj/QsCY2ds6aHTKrhUEhv/DL8Sc/rueW3ywrpa30vQn1fGFg3H5JHgkp+NMv
Cneo3x2yrPLzQ8VEow7xnIDwWpfN11Hv/Wz/dvuP59BGZNBKRyR7Gu8K8hcv4Cey
ha2NncEXyyzRUqzOfg8knzdsWVXsyHOw3SSOuPnoOYtAYdQR/YLhsoA7TkMxzpYW
3yLxnKKO8zddxySfvnVpgIKMaT36iz4SoS8vJ9zTPSlnooZiNx1QxECXTokdPpwu
BYmBxx/NqjXpeXX3eP+Td2BrNHSisK9kLWSQ+hRuhA/U0zVWKYmYQBTfNp/rrv64
cdOi9meVPy3X0CVt4oMRdjSUaBS8EtqT1xf0jf8lxExWF9rxlzC04PkchBO/xv6m
cp2rCT3tU09clPFlZeitDLixCZMWJoozTkeIa9HewXfO+zgEBy3gaQkmA7/xoK0h
N+3XEwrkDS9YhoVHvmWcL+PAnjWy6dspNkmWdcTt10nVJ4l+0SvP/17Q3Or4qZyO
FOFDGyj/ZczOHhD++6POnjUaD08rJfUdift4U0V0RCggCFNJHUv9FPGLMI36rHiw
b4Vs4d1s4habxo/++Cj2apVA55E6R9yM+nIOt6eBbtPsXOCIn8TTwkssigm5l9at
AOXABI2jH3j0o4xgeZtMNBggBGqyNbmJffAIVjpb4yqiKlGdZ53QZ3Q8uWhcKUVa
wxHislq/jTVx20CATDgqWg7UAxiabliDBc28L5EvrdQ5YpHnQ8WJLz4gCyJMBo4q
fVZPxpJOsXofNXgRFPlBeDsP4cgKyoV4DiKlV9qE4vraRsYFVKJ64Zx8My0pACGd
xqfD6VWyV0FGgpgkzH6OPFtZqBnq39d3ZQS7SKjlnk7l8q57B6rXfbuBzZXRxxlu
h09v047rbbhNjQla9TPeUq4jRDc3Ys0PsmJ6M1Aopiw6hNOYZJmm2kp+92JIja6E
W6p5bkHx6qQrNh8T+dawbBznQNMPggsD+O/h2qW7CxXkN9EPt0V7On6hQAD8NOTz
Ljop0YEpPYN8cwX5AtimN8aN1gbpMJLDsfK6Ob/7y0C7X/3h3tIPC+xZCGR2IKf0
NRbhoktM//XpOCzuq/xEtPiAbX/W33hr3dJSGddpLS8HN82Uqz3uerdkyeR9+5jl
sbFPIGDQBBcGYCrZNLr3g8vTVaYgDZwRszAPIVJDVLenYf8qVFxYk2HvXfTw3XpZ
miSGReSg+OiniZl0YGSJIXxYe5z+H30S+sojNiE/y0CNFaPXz5me7lG9sOvSnEnX
u9c7pCOjCjiUyDEHqLetPUOrOIvg2yOlae68P9BmdAyJsXJcggTLk0XK5iyWed+Q
qdVQZiLNUVIizGjQKmEiTCgPiotd0+C7f8hnqzt2oC0LF8ZFi7ZH1IYcjSGYA2o+
sHWMfzZk+FnYWN71r3Lw/qV5KRbd6esHbYz3zH0PYRhsSTJUlQLXsVUkjdoAXylH
lmaT7cGknzzUI4ogQRNnxVKkLbYyR9s/GUi5DDU7ZvK7AkHqGOiy6J5ozBWReHdW
R+KuAwseMTK9jcbPhDpZaj/OvNSqlSjJ/LVIG73wNnwCeLbpU4i8S7cNeW1WRQuh
BHxdQaRoyXb7jpMoRc0oCgL8zHRzdihhK/ZKlnFW8ZyrIXrk55CZJn3C3zjoTJ6H
ZADAP/Q4Ez8ETBxYcPf+AgfMcPaQ8p8f3brBm3+Ef9gjpwGGuHJzoD6fOhxM8tkp
LaKDaMyf4mMbImt2zRoNzdvm1ypFzpQIAziv5f+0uZYyYOMHNUzEz50SDi9XDUtO
UNHYkVCP9FcVh47hHlEZcaYQob0DU0kH4Tb3mqK/ti5O1AQ3/pS5yXg9UXH44ITx
R9jDqSxEXiUCxiae1NP7QIttCb0wE9RXA7MUNTC2XIXfy22rbf4VvjjrivX5XtNf
PVjo56+GupMhybZcWLg201jKfFIuAD09A9GOGBfD9ZfyOT9dCznUj/6ozVq7LsZm
GPVp+VOGf+8eGhF+R+oA1hgjN7knKzcEGjhS/DizltS/tNLzUZhCqrKdkH74dSuQ
RR2eH9us18zix2e30xkxE3HMcTq1X1vysZ2NtzPgp2RL6bs/dLJyjnyjlMpi5Q+N
KzNTSZS30HERjO1X0PYykaLtTmf65oLLqra2zfm5nLHYNw4sCCXFYOV8tCOyUaOQ
BewJY2rt2ep4uT6ZAXTI++bkvSYmp/4RnMMkVPBcaq3ldRL3gjFnlvm8G8B5E9Di
x5jR/KNmflj+OkR4o+QrKJmqY3jmDQT9wsV6fzWjTesI7d4eCCCS1hNKQn8PTdEw
t2SS6gzZI3I66dqKP0xAlYzb1peOLZwXcx2yaf38jXiZOVr4YQoW2iDIBQ1XY2cY
vKv3sCVaFPJNUlSS5sFx36Kd+1pJghep2JKuq1QwN3VH0qXJqKJtLRUso621dIqX
+HRejiMWZm4tbDsIgvud6Sb+v/Avj0JHpEmEEbcvxTULNo4cIjD7ErygwXpf/s8S
c1SqJmuNZ1rWEbjHLLemXMcvGskaemHbhaIjLaAaX+BknAfyOeog09YA1lgrVI06
xs/hSqot3XmTg8eZpIX3b8YK5rIqyyS5XIT2qA35K19F/3D8LF9P5IdY7w6D3xaq
2I8QQuoRFK59+AJr5xyKNTnU9CuryEjsXtVR4Q9em37cXeq7CkCfoc2Nen7/gd3z
jcDp3YliJcDd2znEsgMGmWLsxvhX6iIZ85abRsS/6rA4G2FOafASNqNJftVhT+F+
9KkEkDbRPc6XP/7j4ayjnU7vsdyZG7u5wRgZQlqi842w7XP+rAc6RWTXq8RmkIbD
GyDsCGygiqwHXWyBjEjgR2Iu+s05DGTaSYvziIoD9XzxMMz3jRlJqfIESCu/ZXK7
uYu+7fHL+3eoa35K1lKjgteAHgpnT2Qej2DuEE7XWpWUvojRcYpcWYIrt3uD6z3f
6Tex0Drb3nwOz/ysGHRe9vc9hx7g3SjXXsNRgBC0OfO+2+YVV21CVpBWECnEbilt
soypb4blvxYNjoWbxjySkvrmpKAdB1kGhWPdkSGggfYBN25VP/G7j3GEu7fH1dnq
OqbahiXrofVRHeYt8hHagiorUc5H5GdskfHmNpIu2vQXRugU0m9P20BUK+t8S8fH
iPM8kNHgTcLDTRbzVEm+wK+gPzO8p3yKflVfYmNXqb2Lryqw4NBDeKoDG2hSQfjg
aRYXbnkdgYhR9qfz47JlRJZs6BBvopJYexBb+KH+21N1+CkBVaiNwBiF/fMnezKN
/kLtgijfUKmSmB+/JJajEUCzjqtdwzpukpxy63vlytMU0+yjGFNr0IBWSAPVr90y
vzGumLkMbOj2Neb7N8d2M95BmQ5TeK7HCFjZ5h4jKCgBMqHS1St6256TXLmxkKpr
6LMzfpwvVWVR7hJ3zQpRrtSAXgxzD7vJjDWxOe2sLIL5xQbt8K54FSXAOCSMPBGP
PKSiX4+YSzI+uEhgdaBeOWtESmqQw/NlJh29PwX7cpzmuAEiyo99VQ5ADbM2OLe/
mNsBMNjnpWln680+6v/zJpjUa9WyQ+L/GpbwGuFnxQPyGwUA8WlNFi3T5tdNvA7X
GV0vDUqnxJ/YzJApwdwKXStS1wrulz0m5nwf3AkX7R3Z7uiXPepnv7GEdTD8LAKq
7x5ZrRatoHnCxZHo9/VVqPUA6aE8ZcMg5Gt9yhsl1UJ5axkt8smxBUlnW8P06/Nf
hmapB0NCuBA90MwP1HPp2w348ut+GrPRtqLy4hrkYxMxgQoODmn9iTQsYDXJBcTg
6q/WnHxRQ/oIH6PzcwNbtF+P44qq/X+m75M5cn8vQS2WcLihgh02gXg8nZ7gfbHt
NeLGfhwqnDVhAlb94zOtwKn0Eg+11FRC3Y0HE82f6iFXyHywl13uHESi6rLjGfbz
2/miF4eX3E/aj/MiueS+wgbwBL7Q2FhV1+SsOLvu/aUVdPyfbKAleh0JyLAc+Eoi
sZa663xCkcdWCTMnsBPS9eLLB8UdH3TZC2tUenbs1aRkWV3fAs1Cb84Q2UPCwSPj
hnARcdVL5Zj02XwH/9sJE+mdn5dhR0AFW17B5kwqbeZyoxHqDYH2f2FpVvICoAlX
7XNcS1nJ3Kxs76tQZEJ6QZh1mooFAa//Xyt5bI6SDpJ1FqdBkUDOzilvsCA4ZxL9
aJOU9IXiIRSP/XeC+Eb9FPvBrYqh/yQYROLvwszXn7Vx/fbJoC1Ts8wI92YL6dPs
5iBa5e+WNxVrsLx6TLWo/5YzbS21rUpIpecbRoAXueRI6yvUYXVdlSb5Rc2Nuyma
ujEUHIZU6LgtZr9mJoybrtcflkpmwg+koJpi3SfNTy7UzgD8uNo43/lF2kj3jQ3I
moKZSizWNYVRZ1wfsefm3nApU4gkYL7kWTz55UG96qG6CF1+8x7CMgvaVYy5j/Pk
CdahxpY840SPTMGjCt+iPbe8SRUYqmQ248JkVVrUk6zcnqcbj/w9s2ira7ZpUNKM
SJQTehxeU3a0PsdRLmoGxk5WKAXmIJumLLVYPzKacsuKu8OJOPUULIAQlhzrcJzK
qSU7obPsl8K5WI6SZOJxEZOW9RMejSjnlk1Tt8v3YNmZ98uTHUNVoQVJKzTAZzkO
Dd+GcoQx7fTqMH8nKt5IcSQ8XohDiIysA2NjgOPnb/nQ/CDSsAdQrdZ7m+5bDAAl
h+QJUVgYDV5rl21TDZ4eGr8IFtdty00Ht+s7+MKF530cu7ud1uLvXwcwch7A6rjd
sR5C/H6fNH3zxOaqD1dKbArTbeMCBoO+ktvCzjqF8RrLcJDlO4Gf5IukJ0R9BQTo
8wZo9aCoG3RFLVwIORdrvwYSh29UypjT8rpPRlX36vnyWf/X7gHLaqEYmT+240jI
hljtjlKJpDKw4hGJq++xnUD8UwMyjadE0OMJMyhq3A9PR6/pZ315EaaTHdV/d+I6
bouCKG/1O76vpCTik6M19N/SLsq/57NF9yIKy3/e1mBL3FtES38b5png6usZo+q9
5pEq/I/7gzRUprXQ04LtFNat49RnuanYB6xbh0d297NPfGdm58zhyt2MWqeYyQFz
DC4hk8iu5JZ0dxM/zXYG2zyMFcPvUWA5jF0+pDfCYGtENfIFM1qTQ5PLgvgqz+AW
k3kciH01sqMehKTJ2fYTt79eOSq47tWADXK94v3SkPcZjIrucWdYogjB7smxmvR/
W/CAPOhPl7HyxS6su1Ur6VSZZb0eISM4rJS0KyKTq4URn/NbnoWsl2xKTbqP5deU
syvZu7OSlQxc4400eekmRNZbikwTOaHJScqBtvKQQ8VLEpezJ4EKezuPqTarbfra
j6vnuqeH8pwIJUmoN5bjLQRtD0F4yfHPTALQdDQCoNklgksMCa1MRXNf/cnOKrmW
7hY2R7rWzPJ8VbhXMLlFSqVtMDlqjnIlW7YEVYIuSfdSNa6uzd5O9J627uK7pOlg
kT7+gyodRM7XESvJrFG4fky5096bOxVy+HzRN9JYC4LV80zdU+JWPBpjqWpJlKmZ
9DNll6rHkKb5LYSZ/Oq/rBeakKXRM7gnquPCNETrODDhsyep2idrK5HpMve615pa
pyfSN1/1xpnMBbWYeSDyQ663/cU16D8eF8GQ4QAjlogAOuJN7OC86A/uuFsyPBzg
sCUtHP+AJ29lZfzeGHzidRVKJ1GR+kPrShAYQuOx6qL4qVNXR+13E+ay4m4ex1rF
a1Wm5DLrw3Q+UP+NdR0uk/a6JbURgSW6jv8E42BpA9mH/QpoV2UU+xdccLybl/qp
1i466bB2JRMuWwPWs3hsbahVVPJyGmfwCj1LXq1SPRJwEFWXebX4ZSce/4eeY1xK
NdgZ/wCVGiv7+e/P4BFIck0V9sZxPihWVzSYkLLSnCS36LSXfYFeeM3hjtCp11iE
8OHEcO7qvzY/Tf+pDnAKki5PNaLSLsT7Pf5dIn+TXXm+IrIzrf3hNNdA6tq9wyRd
NoA2DOdKfwG1g6h5iiK1naKMieMXKkCH8vmVsyJU+Z07UijLIkESoVpo6OppYtiX
satJYq6Wn2kYxHAyctet+EGnXh/52syesd8VdAmecnsJTDfZcpsL88AwbpQewfxd
y2PtsnasOhRV0+uvbn7LOgZ5GSs6jM2+0TJLxuh/S+Iszbktk5d/OFQGvcRJYoKi
WtiaXuM1bL84SOQIZF9K7H6EjaRZY49g9BgJXP8Phu2V0CCwUGf54G3zypGSRm+J
t47pZcNX1MZmTORzmC2cDEKl8kwdCE6e8ZjtGl/fzNJQQdHzyRA7X+tHW9OqAzSo
95Sd6lhOFFPsYldrTTbVpvIDV1WMDHT5LhTIMKnMRKU+B43dBmGmG7S62fqGOZDQ
wuBNuxKSyCbiwsnmgkyMOlAAvUpk/wM62vmSIVEyNStWRfnRiTbJxC8wOFcumpCj
XZAkkLKF63YvTaJE36wNzYv7Ge5EtOMs3FXAub4agMypC7cHMoSTIaNUqrOpFjHZ
exazP3PniqEU3MGldCrEgpBO4Q7+3GEi0QYt535mrz+SxYo1T9V8aNhV6rLR9wq6
9vGyY8Ui0Nb7A10GRj23va5XSAZmkbgsL2z4WC9q32tFhgKVp7rL3ZrplFCfFHkY
volg1XPEf6kbOddduDZvXDGpSuE/2xNOa+n2O09UAFhKGNt5E/LWg15zTHzH+iYv
iuxI5xqTzoxxQJLVaq/j3Fxa5LAtsrhy7Pr2/q1F7DdOvEQYVV3vkIF1FY5k131z
O6krOH2kk/V+dgLC5dGz78bvlkVUyg4otqkcoPHgrk/yFTAdKOmCLAWOulmuz9hj
oudhcXwNnFf3fb6vZYs827ZnM09JIVsgqbzlW3mYtW8dtP3fCxeDZJbg2ysbI3Bx
o4hOTVL7J5XyvHeV7NKUv5OYMLbPs0fGYRwxt8FqdHXuFcBl7xpVULyfpwrEpv0y
Qt9g4RzPAG0GnUJjyCtbzO29F5BNgRs+GWRe7OnExzlq2cTOrD29oasMTFhISiHH
c3rZdwgmjbK6AS5CTljlpvGJj2VeLOdFxNgOtzdHNlInvQsjlYlcEL/zr/4xCRf8
pN1Qr4OlZYtB1yGuHpmHtJ0lkqlKO0MaTFm0MLN42TBD76FG9Xij5WFeLYWNyr1b
3DP4U1qhD6v06KeVbPKy6ZC3t9v/DpV0UE8XfeKQURjpW1x3RJjzQZCqSkxSZaJR
hKiXoyNoV97IFysPhy8rvj3B9YQt/eeDlxXdkmkSDlM9yjaMozJVThF5Kfz9KPK3
Smr3Z/oitFiyWNalKgXM5iM2Y/BTWUFtME2VfUac6lu0DiZFqo2jwf3dz0BMlMqa
jzdRUslOHdE09ZnZb3j3fLSC3QObSTiZ+QNQ3OHxzfUnnQhe5PXA45pDhDK/2WwK
6tfeqsODinPADiYDSyAbiS9GDz1hjIJMnpYbKRYu+ZJQkM9Z5/X/KKAhVjcHIBG3
BTbOXrzRMEXVuAMd1hTpnV2sC+kwQ3nnm5EJVZzjEgwOab+Jo5r9GVhTgRIO3gGv
a35MC1DcZoTpu0TCTioMJfPOZcDFT9pID0vVgwjVc4RPP2WjeQSP6/StkNNhJaoz
NxIXI5KjPg9GVZqRGaSt1/UxE5Gm/G5NSfXR5RK1xaC9iZ+xDAmqKPvfSC7hCJcV
qgdNveQSJLNT590lawiD5QkLYaGJ+w0OF7XJC0AUCpTvJVlAjpzlnSaoFkvCWAC+
DhhEN/zYjfSpLxa0tZYWjDPcneda/JdC90l5De0Pqoo22UOTqzTFjoocp9Atgglr
wRlgK2FslCkosU1tRzSFEPCZgJSNF7VJFyVzEiYjZTgnsHoGjOOxhMTuuYIgvxmD
2YPY1ZGySTys0zuAMmXy661lPnA0WXV+Hnb+c/rL8sUOxphL8aXRGDZVdT6mMFjE
iTWKRe0Uk9g43gBxbPDnD+bpG1+DO9fMaSk8DpihP1P/j0wlvQvPt+i2tztP+hlD
hZNufp+7IUD5FDqbGRt249h8/E+n0Z+ninkDHDp+ZLBbQ05ovuK5XnGQ+i3zcZoL
W+KXfiktoLAIgvxJcfERpyQAouIup9O9BnOnNTljp94QBkXMmJlxFaO0+/ldlgTH
QpB+lrKCNJQmQd9k+VZb84FcnQ7ndyUaiL3lDFHAj6JqukNd3JpISHZd71BYQnwI
X2LEU1OzgAIvtJD4TOOgWC06jVgaRc2sOwB8gGekQkalz4pX7UqUjS5SK8X/cEen
fgeqmGABGyt5a9uTZBEiWS2oujlE741rIy0BcXMGOm2Bw4e38ytQdITBoybuNvkA
lmW2xr8V8ZxDcAew6rW0lMzXJl1QPVUxuATE1KmzhlCnOanF25BPyjIKsKbpWLQS
pMJ+vO0zghk4/JCwka4En9F2AhZdbD6FeZRIUW5Eo3hhQP4wiP3PZAFS0P/vU9AF
OxeR8UIn/2iegohKVnIehUZZswe3yurjy5gOQpIMqJaT9fgwb1x72cqJZhGPRTug
OxCALHQWpJFs6nBjM3xhAbLDPvyaPytaFsMpLTcmPUfX2aifH3+9hHPt3CxhZ5n1
+rwDFiSgTqiaYvOc8s1uFJ5lMDFUogijEo1nvL5+4oM0799OxI09/aAssdW3qDcT
BXPJgg/TuBngOFE0Hl7Q2eoSKsr2oBh6pVjKk4AuquEbi4ZsMZm5vLxQ3mqJimQO
8K1ofnjoCbiq19BGXGVXvB6+/WaEpCPIks9kOVXWKuFPWXjxN+I/n8ex0W9qhdvO
U/ox5FWzLwVWGuztvlrjbQXL1XkJOsUbe39BXUrLrFp94xrWP/uEku6aro3GqG/W
dzaYaeEsK/NmFqjiq5dsBBaQI0JzS/Ek4q8lpV/yCIfsgS7C5BG83PC0Pi2QXToN
SIjrvYSOVJ07yY13lRVc7FjHMg2y7sWzBQG7s7BAefBgRaz/QAwIHnZJEvnh16iq
F4PCEtj+ZUeW77N9/FZrAXQS3+0NNaAu9D+sSzrlQurkmSxXwh14htkIZFk0xgfz
aIWVERY0Scl7CJ+zOeBsI7MP+VhQztxK0KhKx6ki4zRGQ8IIUE0J9x1Oa5+zDFGw
wydbQLxbjpNEx23yCDEFNnnojSzb8I+NQ3kXizcnaDr4fYDqhs+A3Tt7noOqVHsc
MGqq0omHsfVWv2q5vIGhDEZ6msT7fFlSCV0jebhp/oe87ska/CbaW67ON1hNc10n
TTRqhf3v1iGV/mV5WiMFQtbnMn7y31sj1xWiRo/qEjX7XR1swAe+KNFMhgp44jIY
f4LH7997mwKHXGMu/z5Jy6Lsg689twUUjyjCHtgT/2n7OCD/tONkGxb3kkBDJnml
ZcCHpc2AWEzUvMLL2vHyWYByyPSZZ+rGxzPnGWUfibayVXvN3ZwT2S+wnsXiQT0q
Mn+/GOh4z7jQu46s536qatvFyu07vESeXiBRf09VGeRPhyqr1Z08Ej71tbBpYsyZ
DFPUn5KAMb3tLFHcjCFZAn1Q5408yocHvUtFQBeoHR5OkgSmxUzDxaeSVnAPaU8k
o3I+xV+89TOfPDDc/c1IOaq7t8cUwNZ7ECAMoLM/1VUx4wSK9qSSZXuzRRVqv3Nj
O7WcV7LqrudAC3+xpD/Zu+6wcDAqdB1qFQwYpymAleyPVLJDtpYk5AeTui9ILLSG
CB9HQP5Su1J3MsN/Tnoeesm1w7jvE45SkF1k95vLHZmQOF6W2/dw1NJBzObutzk7
2+zrOHE24zm84ZbwXNYwMxhxZRbcqUP/WAPNyYf177Lgh6oRXrZG0e+F0TpN5Ya5
E+I+06Ygw5sVbEXdFNV2uWweMl2Fw+tqIje3yKM9jGeV3JwfBSkIVWL2+8kJ9kgY
b909r6b+ZT3WdExGxO4rEEf4hKnK3MeKRlNr1LThtQZiP9An2CYDzfluLM+B6K3+
l0QHV6Wo1sROhfwf2lFmhUrpilzq4YYPiG1ggbk4WjjZW9VJd3arnS/poEmEMtWr
BrJaB7czE6V6DvncHpzpnjxhyGAB3KVC01P/23fpg0lttu46NEslwOoJKADXi2HQ
hvpF+ir4nBk4LkJ1DwYcXG2pr8tn+O17SQNsz0lctNV6R3YVC6W8MBoJapaSOAun
OPVcmyiVjgxuEXTJjJgxDXKU85ZTM9g5dhwlRJ9IOQmRqM5LaFm8g8cY89I7h48w
HoI9BnZbEw9/1Xok/mlmqqPmSQ0Zm85ckoo4OzhztmZAC+O94j+thFtw9mcOq3z5
aRL5eklGtjOlSQjphh+qE3DumYAptFJPRVxujm/JULflUYmWflWOfcCCezWxS+tA
aOeXdj344lYa80SN4F7Vw4pyJvDhG/C6mpTIEqWTDIw12dHwi5Xp9ilsCx0JcvZp
JVj5RAz7xJFA8BjOibFaT8Aux7L+NVKXM3G3N2rG1HEBWuyxPQQjWjuLbNXn1BtM
EGabtHF+jfDUHAArY9PT0oi3rh/aFB7Tk1bMbkDMAj+1B2tO3wLfLX8d2P3oq8mC
EzdnaMkMjZSF+VQaQ5EfjW7oxFLYvKpLY0GTBYyMtxntL9mTfCfJ2M5S+nBwVzR+
1Gg2GGKPvxV4VLsosDOk14ve/XjdgRC7kA1ainRGsHXhL1NMht12JFAGMb+X9l2S
Kn4YacoyjbjWyUd0UTZ+/rRb8l/0yUkVQTVL6zWzQxlmtrndwyh0WSSTNUkM3FN/
r0l8HMcRuAeaN8ixfsSrLFYqgvXMQGWKcdDXuf3LI6sY5QbHTtWjXqsfUO5y0qLm
omfkmlGIy9m8v8A9gdjN9FjS4PKoOf+2duyh0NFKmvPCKdLqtd0D0xoH2z5KuvUx
d5u1yrfhfywioTzirQQbQBbHxoC0OVjCthYIxFrXrqS+3i7OU10MvN5zieihwsk1
Bowika7fsSgAWF0IVtinHXPhqwQx2bN9fTXkFNOxhcTXZSW6mel+kcJ+SBpBrzgO
dEzsYb/R7LaosbywSNpVPtbwzKGAkAW8wNYQAkOkGI62IpPP567QjVeSbtoWgiLi
e0Epe7OociV65gN8vnWewNDmtgdeQ1PjiQ2Tj4nSpUsOAkYhlv70N9L3E0Vck8q2
N+ClJ2P0H0hd0OB1RWmMGJo+KP1tiTgauojZxe15orNTUJxIq9AL4M1mdmqMhmk1
2og214R6QCqbOsePZAecykghNxdchaij61tyoJ/DuOp14PnN++K19D2GR3cBCGj6
wfjIxedSXf96MasUtu28gDNJicY7DnP14r7kCuxXIaTRPv7KudDI3U7R4uBTEO9/
mxoN48peMnS4D+N/qHi+NubTvxzknl+RPRxH467gBYVL14hJHJyXISlh8Zo3Wwmb
cY2IjehVwapeQ5MNHer2o7Q/zLcFSxFUtDebkTPD8VPvDpIZ+i0o1R9Dtw+9oTXW
IEGzC3s/4XMLLNrHFWbjkcuZci2S++WcxeGrIW5+fgxdnNvu0PJ4ogOzqJlYCLFE
DLVJcdSAMjvU9mmLtggfpusKFGoPQZTVJdhCV9l3++GjUe5NQSByqqNfZYLCPOsm
P77rOTbeOkUfHDHugB304EFMeV+kFgdGGU53uZjaxM2e7GWkGPnZuuLstiYXbP1o
IaTHEGyF0suqjtHYGNdJQFmYS8RaXI94OWwCzVc0cGm2PLFcbYzBkPZb0wQCjkeW
yRkDKbrxcYDeCZDfdmq8e41RU/tVtzIOPDfl9Irj6BZ3VhMc/KFqDqkdZKUO9JBW
4Mp2gXwVc6qXUg5JEF3VWIXrkQCK+rPtkeGSf6a+dG270NY4kso05TsFiwyw+nrh
lQTPyIh8h5Td8xvF11o3ALLifCKwB534GROGoJurdQSVV3Ci5h3o7H0wYYLTADim
YV6NmtKhW9pq/ZQh3b1fGvFG45yWZE6RBcLYMX6sWUko/YfQxfRhOcvRsYkwK1i9
Ma9VUwnjDmCpEiZ4diueaoMGs00K97HDJ9W81k5Z23jKiWs2efjGh+ixRgBIiZKk
THpCKoZkFNi9tkRxur91Mjf2g8njx2akRexOrLRaZT13/AXFAtX1IwoyWcjDR4BY
em1br/vAon/VzDffJ6SxOIasZhDb/S02RKEdc03FgasUO2nbdIL+9XIiPierf23z
nyhjicq/lfAzLyv0DpIB2OtiS++mm/OzaePdGaU6WFjlqePnxnjT2whAnCOSSWoV
YUBmygMbVfd6mpEbZVv/1pvIAJxMP/Z1ohqy617osdBRFh4TuAytEcLEEeH7IWUN
7ymsHSwQ4PwPFn7rb+zlCCn1LK1jtzzcusa8nYGnJSAJr9tNmidRUrgPyjM20FdV
y99fuufDhDOY2W8WWFWJnFkyUKHeE4JYktWRVM5XpUHCUNqmiuTU1NIB/k2XxRzI
TDYC0cTRCH2DdN6Nz1KUJZk1elKEgv4vMxVXnKuWzOxz9UbzSUsS/dWBAekIJOLt
CC+CiQk+72Fd3D3054I4T0mZy3inm0oQ3kNfa6OMz4fwQSETugPIVBxIXFtK1nED
8hsjwyrCPJnm/7/MSpUQfxtZMAH41p7wb/wYSirskDvxL+4OchujzdDX7MsM+rke
HlQme/+IsmKw9f8B7jvOTPuW2ZnAVtS6OBT+ZdQmcx61fWX1w9ErvpIkizAWxfgj
0q26b0qDdeq9W1RhbWnOwrIHj1NeQL1pmcBW6AatfwZ8llWNsJ0swuKQkwkY93PR
bAJxHVwpVWIimIa5WahindpOGpWmD5Gb91h20urTJSieSpUUuxJ7tGISuMDqtBxw
R3eRIuK/rGbrmazZ+bNqgCcHDz1xrgR9SDqRGDfQK6FRwMsFSTmpVnBTQusGyWGZ
qk+QLW8MId1hZkIHBYlZlRPWfLYdWm1LQqHYwCfnnDCFjHB4y6LPRnGkBFCAmB2E
Mhe6hfPiaJl73BijJXS+igIYwbkfG0FvWj9/SzlNJOJw7D4/LNZIi98BHPAm8/sB
nW62WfMj6AtGBBZObSH0EZITKICVWrG660CEqA9vNJ/GfmbIC9eZGi7oQuskF5dV
5NStesByF4gf8nR0ItzdTJbE+hw8KSyfHp4r9c0JSx75xwf4FORE3JoWuiITWmG/
nm+bmtY5hn67CHz3Ge/XhuwFy4bZTg7Bw+tujVquH7rl8czUElbhvfwfMJaGPdt2
2tjBgoHMbjCJ9tZcs0pPAiNLPewqfjSRNZgk4i8nIfxsIbxeMng4jpxn0hu+Qpl1
KLXSKs5zJ5CkMQ0M/NpDHbLo5zK7ujarl8SfxRVPRkFu2HGs6aNCVtb8k5mEYsIf
k1rAV9v3O/hEqkoVndLcFqgtHpyIEFl+csAs/cJh4XPZc7F0/UvM8dyYIxe853/+
uM1mTtbEPln+jCajU8HNaMJDHXRREYupRwIWqktyuyHtM8X4tv4FG+FO7EMdguMN
QYK7OLBrpAviTnEs+/bygYD3jXZjG1ssZvaH8tRtKoCN/aUyiEYtjfgjvbjXylQg
mHikOFsY3n0LKh64OCHdVsIcZ082x51OdI3y7gqM+1hwLZQXx+xBMJUgAwlTcbSc
2tf1XP8u4sb2sUvTkgAVIjFxRSIVhaGcDX860RB3PNnAbwuyQO8EQuWoPmNw9ceu
sElWMa2nCWUrNr05vYRnP4zXczvjvJVABZHXoe0OGV6MIHkMioQY+d9Av7W/f0Uf
ptWdTtWfqfQ2364uoK+5OX/Cf0/QOsXYl6Hs3+2m0OAki3dzmLwlF32maavmhV1g
8AYv1u4G+MGbrzUEhQN/rpe0LWVhw6XsL3UD8/6H8Cp55Jurc7P6NvIxjK8tl1IX
aRF5/N40USfOBu+QFz3QRCTi9B80UGLg4OpuepIH00HyUluRvfhvZ70ex3MIMvvg
eid86GvH7SP7x9iGCYARQ5m5AJklD1W7x+rv+74+qyhb1Q6pT3CBhnX6gWryFqkB
YZPHc/XR001EaEmPLYCX7W5obzp3Vp0L1bm2b0tNzsUB138U3rkZinPW4tD4+Dek
QKzEWx2hhmfvd++cPIojfSoGjM2jxuVfe3wZD1V0z9KG6JMkfGpHItgiS5+/DbBY
Ak9/qHIfmMBj0Y/T+Ki3XqwcX7MvlVXtCB73EnfP5abgE0AMOfp0YFaqLlJh9GZC
Yg/EccvSdO1YcB1uQdyy/QL9Wv7lAtLgCawFMbvTJoUNIX1GjfHXuQQHDEtYBv4K
GVmq35xz4jeSzfsGD2UC513VXx2gdm5aZERQnMnO59okHpInApSv/CEHtYtQjWid
1Jyz1rCCZsxXchC7agKI16vA/HPb2F7NtNZQGMzGj6ScCluexjPlvOHJwe/Dx/6q
jYwlyhRCXuuSG7/lRxiUyecYh6tQXmoFPuFBbRKoT5/Hc6cJUZsMf48ICfEwQZ+U
ft/XxXHlj3gynzvng+qpX9/vfmnoL3AW/+bHGXfUCv4lP8JkPMtG4PXD7F73IXqa
dbPdkjMu0Quvz4OD2jTUsE0kozHLU/XevkDRW7BMMvaUcvhGLi2Yv9EVgrNjD3qU
XVMjbvafOsu5N2awmq19mPEU68cFDTNzYNAMBhWxw6T1UMD57HNrs6MK/DIG1Gig
I8QCF8i+n+fEESQ08mMjbPwZlAhaJQ7KJo+MDXyeCC5S0gkmAtmBngrsukyycrmp
GvISpdJ/7AIsgcX2fCefxM1IKjPBsMd31XnQtsIFN5+JZQ4ZRMGQxPnt3lFENuGi
y8BO1mWi3pUXfp3D+BHDExx5OWrHLSOjEtWd2biu0vqlUkT6WIgKeA9m30/4+I3+
hQCZKQUJ25E03pfkdLdor+2VwofSUVTm2i/W4dyHZakH5ArlNQUBC8rZamKQvekJ
/UQxJBainLhMxO4Qc8ObXP+R4Dj+Y5/cA9BqPoeeTYJk0U5R2jkWsHKlVIjdLcha
i36gZZ+3ZtUyYzKt58qup55bqTMsXNO1P/xd/z6G+xaKtyrIjfIvhqaVdMHOYbvY
zsz1BWyZxbO7jGFDHnWMga/wYeSAfcoeT278O//g1pAsD+NrH/9IYHfvRaoSAUru
H/xmUBtNfkslONieFPBFC6rifp4xwJO/8vnihh8q0QGUlQHr8wydSgf+KdOL9wxS
QKy3A77ej7f3bQVAv6VR6yiT5N9dv2tQvbeVopkSZIx5T4GOM18vYc1o0n7q8Hrj
tt9MzOuYOyseeYeaRqOSLaa1pNMJBrrjVyHOAep1I0+wm/6IyByeADqF9Yn3FVQ+
CBvRSpJPs2/F/GbbMVfIK589eMVPb+bjVWkLmTFYAaBYi/qLZGKnKZoRdt1cHpbD
mb4KSTjX+QOJNM6jhmTG1tHdAT9tNcq/cQdnD1XTRE+viDcqhjee0EOKRMRMabGH
sVLNAcMnVqcuzFk0G7F/0BG9/76ESMpab0hYqDPsTaVFqvvCDQYmozm+qjTdKQpE
tO/OPAX2vZtXD/rt58NojlI7uXNzcJHpnt4srLW+sBOiH6kEwLk95chBBx3o3VkJ
O6FD4tDIwBcbLcmfu8IbG1joLWIGxEh6jxQVkDDF1EF1hfpq82pX98voWvkWt7rw
euKTwt8FptQ/vah4mOv3ZW5Enx6yh+fQCeaJVJZFa4kE3S4Cl1fd7w5yflJ117PI
QfXGVm+EQgk45hGhprXYs4+GIlkxt8gc01YftM6Mc6L71qdusLIFr4nFFMCrrBCA
IjpObUlz0N8CArx06yCTmCr2gOXOa4sSX1Ue5tE9KP8PmNgR0GC0gPhynHiy21CJ
dCRkYhjpatNowvGPf1MacUWf2Cn7G7wp0N4sT772oT+sNatGdQvgPkqctSZ0BWha
yv73a7RGsJJTquVu9V4jBvXcxd7pAXcGuOSa1OflblHAxcnksP8rHfVDBxnr8cRR
8g2IYQi+pDBsBqJY1Tc7dwZS1xgZ9mJXRoITedjmqmTMSaHZkmNi+1zcnXbaDI5j
ljcZrz298kwrnlwwoc8NsiQJaTsytgYfs3RFo5xBvLmMhz9ONwzrRk64/gJlN0UV
xn5I1g21nfvntEYekF+28RXiW3Tu744Mz2DqOACi1gPJWta2nEIdzYnPvuCsOMd0
At2KweZSRXEmuPHNTjP1gTrjHU/R/P4F882PyQFxggdkdonj3pOuThaRs6OrhjOp
WKTdY2AUaLsUtW/8rN/poq3UYb/HL+MXGOVdAC30dPo0WXxBCH3+BNFhy7V5+CLJ
Wab6fPDcGOSJ3kST96M7oY5QmBAQX1KIaB9RpTjWHp3d0q8dlUjp489VyaPZgA6l
5u45dZWY1VQAFdydj2qgmBZk2NxIKLoFUYWjkE9WQiEEdvJgVlSrIB9E5acbAb+N
2fJTGM5bYNle7vCw6ShHxlT7WUD2WDIACrSV2nGqFnAV28hkde/uP0ZJuRzBvO46
i3H6pxhmEu2xWm/7MDGbPfrsvNIOyM7LakfJgsr2ncldCZJHeRJk0k/Tosc6Nx/z
PUWYFaUSTb9y55E/v1XufoN7lzKrQ6dvcO03EO4Eo0Yi8zOaTVOlQ3TtpFEp4qbP
v7s0Z/jKx1ieLK5Maw8Jozmaaxlw/bibNXORwYHB8Hy19rjCAiEfsdfEvRaWG+GJ
/Wq7wYyiYUaNxldJ1uV4oxvmfJGb3Tye+xLZbgb8LfyLX4mt67jfFGdU1c2Kc+Hh
K+hO/NRzK+6dCwptFnUvl3MXter4bqVc1vfSv8WSiOett3nb5xJtnaq6ToioiptX
lAaFDlQun950IWJheVJDxWgnySro/6toir8J/sWWSDZ0KdjtsD0dw5xvt98bAPQa
o2hXz+S2WLULJ4mD93bnz/UqfWiQ6pAzr18c8FTxXV17bUqNGAwks3YjkI2wFBkS
EJOiIR9BQVPLd4CwbeSxxWzagGBOPsRWrP7q3z/w3bPCgonvYPP1dFNGACv88EcK
2Q1e8ocL5CPf7bPegRLWTVJq9R+wH9v1JA0ZBwks6oyKsTXHLOqCY8yuQk3MUehK
1VtZ4G+tcNUtrgl+j4/b3oDsGxv5gkaHXTa2Pm2iJnUGxtcRZHyjphMnM9I+N0Ti
OX3YbGX6/wUzXfZ5buwAr8ONsdicsCsWAPoqoLtCkzmKv5FK4q/DIKBVPlfp1zrF
PciUPx8J4BK/VC5ezhmUA2NI9DVKg2qfgfxjFuDbsCxUacT1ARud903VChD36Uve
dGmF0vMokL6WpURq1KiqUBUzXFuhl6YokJ8eW0n1kzBBCoBLnOs74S5nlYkuBsIu
dZ3UeU1WL/lGs9NRNXe4f6Txvxkr8zuc5vadeVGV2Ixz5CLFCxIdcSeBDBzFK+h2
n9Iu7n2I42vlbGHvPEONmZpiLYtuB304+Z09zplScqf5rtXJeRhk+9UP631WaV0Z
IYqRdluN3bI9NfQuIp0EvTfOSbCVehVEHgnzWHYDWnhI+/mlWBV6gOnqEWkEodp8
pyf8iN0b5KP2MUVBqJEz/DTYz1h8TigUC5XDipi29xeozuAW06eOvIxEA/xVPq1Q
qCpSOE7oKhqXJI3jaqZkO64nZOK7LTuNyYbkWSWB5BAGdFBxIuZ9uLyoFu2dAGsf
X9ijeuWP4H1y5J/yGQSoG+81h01B3cT8JxWGoTLt2kE3ofIUJWg7zwveyrYnlSOk
+PBIIWmtIVa4j9OvE6M4ZicqGM/9eIcW5q+Lq/NtSUhZo8l15LabCN/OQrUFGY20
qbytQYjcpD3Z5+dCQyB5m9WgO/B4nxlevI5Ez0O56eXORohSUg5m8IYApQ2D6UMf
FgDUStE0yfXEPJKYrZ6oPCndCC2e7sHng+m1RlTdL5e7OSx8FQ2ZG6o5jGW77Lu0
m1UJvew+MsKiO9BszmtsOqteeitkZ2Aw9ahabzTsWNu+l/xGckRQlYfOZ8cQCSRh
Sl5MGYcrelEGGBG1Y5SAjbx07UtqfGabm7cnFcJgsw5yCgvJMyIlzIYC6O8fXyKL
6QQAyVRDglFfa51KlSKOIabE0YoECp+PZz38CYK510MR7DjHJZWhR1KotSlhtQDK
TnTyAvoYpN99o+ePPYORrCv6+rNEY7hpKEtJcvR5kxxqHpc/on3ScKv/Z8wcw81n
O5X1NoZQgljOVpqnMOe7JQXkwQmdskDhx0wC5bEfw8DCVhinZv5WkefetmtL0HlB
tgDq7pD4t+42Cc1x3AUH4RoP/rUPH3ByXD6VaWfsHe7fsqYMUf5h012Xx2IFGV/s
Ewx+8eIDivpInOUWWUuW+di5PzHmGWWlRSVPnLbdziOWqaWHWk3xhENl/W+r2sGv
85qoHQ83o9arjDHZI0IFq3YoczjBZFDlTcuFCa3Mp4A9tBR54QgsGZ0I8ns+/lGX
mRx/l4suBKfS5a/Vo3BSUqGPxhOpxqijwmYfQMBPXNp5LE11OkIaL7KFe35WNolJ
Q7kNXmSV8pMdki4gZRTxyd00qjg+zt0QKYd+F0+gK9l3st18DTAo0IuJyfMDvq4l
RC6kpa5GE8Zrg2FmtnwCZiXrpWivlaVv8ez4lBUkeavn8Cn9sitktWVgnfoHV4at
hL5dRaHwILlmTfKsmv+LaGspLH2ZK3fau8c2OzXMLNaEmWA53kgjCahYais/QK5M
bcRGFaHS7U4aWQPeRFpaqll7BrttJfFrVuG5Wzk/F2WiVDFx8Yoh2i3gcqdFpRMp
CqZv92uAK1HuxfwUxv1H53NFtP5N6+40JvXHeqzsmcc6LQciBZUeGY24D/8gi2tu
SNq0UQ5tvnpXMd8F/NekZplg5y50JLVavzFaPBjRB42xcTopbOvpFECXZaUjZWjG
G/faFe+0H3H4r5SZZ9iEoh/LCVjyuDl+Jog9dQrWNndB9n+Fzb2+D4V0w2+IjK3v
QMJGOHQIg+dRZaM0Um8EC9jt8esNyYaI6DE87QejKW1AZKRzWPffTmvEu7oxmmZX
mF04ZxDZQ6+n/AvVBgI+jm4poiBHX5436b0yo60SxbH+aBiy5Y2+teuWeZNnz8kL
YZrtkZQylP85CzAIUlGSnySwoUEEUsycJR6T2sdeMSw4YfnF8rWxB0CloT9Oq8gM
jaaMU/AXY+VCquPFzwaKS+yc54PeUUWzz95fMpUxpwgmFTLs8/RMgBvuRBdto/+j
w/lnCLC2DPbTx3MUdLNGZhsLTSx3LBI8kuenokSlOrs6ZqXxSh0qNO7Kh87XcVgM
1OFUyXVAbZJbwXNdRCGmexPK5wZPScv/3jyxj54UyMCODP4T99+M9BI89EDnW/tB
ghxqlORFhwpXgmI3vKYRu3Q97FjLXmJtl4tqeG/KeE+gLZ7J0g6lMPMN5iBJP5hf
HDoOHpVdIcDv4zBMEaF/znY7Vh9Bgnbps/ARK/mWGf/BTCzA7LOsgl3w7deMbCVl
ltLnlZF3dG0Xj6JzTImnl6TlmzWR45T0GV3dO9oyJfdNjTg5x3x1pbky9253ZvYE
f+hvB+IMJWsBOgRwgVfKweQLs19F+Mkz2G0Bhm5CUKpA6+8WYvIGx4CCwyrZcxiy
N95esLAfwwCRbNZF/zGGDFyxrVR6buglGSybuoRCgaKQqfDNh8qcEHTYRD/kQZas
Xafz5t1DYwx2kEwSa3QCo3BBac2ZyA4K3vqmXpE/pheyQpbR11F+hpQ7Y2bnYm9c
0zz7CrkO1mTU/IogDsFJZ8ccHkmFP+oD0p5pi5T8IWnjTmcOYZfrHHjjdcIWNTcZ
TiL/kKVnsGgcpKTMD9E6FlfamQ4CMyL0Oc14cM0rRvpFsduq1sHWawa4mRfqfp6r
1wZYMcumRhZkgjTVyULRaw1ik78+MHWAAVRzWoQSg3WRNMwRiAUfwjAEDBsegnyW
5HUpU/9nR86ILXaVf+UehfDpLwFNX6vFoQvH7BDB9j+jsT1PP0q0w7Nj6CPjkbWM
O1ZazGgNy0lSI8QXM/+9XbV043XQdoLyNrl6JYIG9pWcR4vJNC/zIjjZzXAvqE3G
hj6kBxqojMver9Hgg+tTxU/ElWweWi1HGzQRVZuyOMazQuroJrl7/9JNw75cV0/Z
iOQYJIenFEieOKH/dZY5mj+V7dFNbTvCeO3zJyNWK8COtEKCeB0P4cXCq42e1vvu
u1SUwEVMWq2TqXel3NUnmZtMKUbqS90seX43wdJUAheMeX7YsCO8IuJ6fasw4mbU
Xbo3P7s/qzFB/ryjk/rrxrh0Cym+0fYc14pTJkUVIFsqB68oegoEp0CxwxoeKKgR
B+pYZL+ffoTT4qvOw+6wjq6vC9y8kqOQ9Kb865jRVbvgsA8QikKpturTlZgt3E9N
egTASqHXzXbFE7IfQLyPQssjeH6jxZIC2SSyadjp57RxKqM9lcCL3XN3zxJ1t5Nb
NA+gUTDKxHg8M6m3BOlP+q34zgbzno2fCU2l88RSadA8rY1FHP+IGs2ay1hH0iSW
KqLuanP6hmwW8lWs+y8v5V2QR0czsr31gVqLR1yE8voh2BqBccidMQueVFzBqhJf
gOtAq9vHuo+MXqhskuTGwn7eW8WN9PzYwspmNWTE0dJ6BHIEHe7sTY/VjQmzSMdD
BRoZnXOHR8donS/gbSF9H0OfUhCoeasDi+4GKK6I7usAJI29APziy+dzqXc0t8l3
J/Y8QV2tCeKbjT2zzPrCupVTR7HafNCHbjS62n0/FFI4VLXPKnr9EuH45Yw9wM6t
PESgV423/4A5L1KBEp6/drvjJzUFEy3kUD+2Oou4DFM0ZtKRvQmeZZJPNOGZr1nZ
y9KD7vy++/DxdMzW6ECumH6DJzbUM6OktSAu/VjqIk8bzeRJ5u3FWdFteSLLBYQH
VzuoPlWWo13Z+/sMxgDw/GXtMAu3W3fwj506I1FR6H1c7lC56rzKQ6RY7IwLskM0
k+SbOqPYssc3kkl33vdyjoaK7BJwt743pG0U/VbKrHmCT54HvxlNHpdNzziFb77v
Qaiza/FnBlIE+Q005bBuLH4kbmyI5DiVs/E+ti7qZjKUQ3uAAmRoew3mL9PleFV0
NE/gmdRQlNI2wmzoHVWRISXUUkwYto3279haPL4ScKhJzlWBb806OCc2W6ufRs3v
q7lB5cGL2RVxqvrZ7ogYK5TV/8G6X5JNfxQh9LG9jVasXsFONK0vwpmGCvCQUrJl
EboWmDlwwfblBQYUt5vUdpNBC7KK0HqPGIpSZeGQOFVFlm+fS8j5Oob4sGc8KMst
TE+om19vGGPcMIb8qNiAxejVGG5ltEhkl3Urtsf1+8CedrrAG9lZ3js7DfFL7tNN
vukbgVFuqj68w6LhN6WoceCmjZZ3H7YuM3XT1bZYu4ZpBb7z9g9fVS6m/t+rlUlV
FMOaJB518Cmyb6oVEAzn6IbHtwSfyq1MyQRDu8EQt4vDIykCN1VVoG2Hvm4+RiPa
fQORqZlc0ZfpEVcLKqjPlCtdE8ILO7aUgYz6mUexII+CSSxhsGfT+lOB+I0qnwsy
tdGzNUrSfySwexY8bKFvzrxJt3LlXuiQw0hi1XTvV8yu31e9tfK/gR4BYwBUUQOX
9bSOSH1S2Us+zHrvI9ZQPuvRMSi0fJPr9HG+dFlrzlqOmIoI/7qHsuEl3QFftKNH
LmB30N6rtBgddVAn0Q7t/dpQRf7NvBfzJul6Ujk8bg4QiAmnBfTsGeBJyYLRtZk8
w4uvHyTQCj3t8TEDXTSED64X8xX4qV4nEWdLea1R319um21V7CnENwox8V9hNttj
+xzJFuVrBy5jikLctkKPzE4UYCHRcKkbNJzeuNBTy/TgD0cQt+G2neeEE6BDGOl8
hUBXuYqvWCGl57s6koTIx/VHBsiTaGd/rrPxzYVKuJ8aIKHUH9E3sASPuCXj/yEc
Eih21gSG1RGXUxS/O2F6ITK+tZ0FrUnlANEwzr6Ifd7WVrlOQKOJClUW4Onolhn3
Brap9M2v0Fdrg/EdWPvSdMm7r45jZgScOv7Rmhy1tDn79qvojRfaJgAPC+epCrG9
CXyFz+WKfKEek+0NjbZO4JQ/o0RzLUT5YyNiXkb3yeeNTeLbOcaPafx6RUfBYIv4
gwguLlIpHTNSQ1fLkuiEP6pxAbgSclgd+Wk0wMt+GCkE5uANqFjnDFgEU0n/9VW8
hjwXyWZeDx7/w1HkRvFX/jxVoyjuxZqogk7+ZGXK/HKFUhh8Z3QaxW8Fp3Fub87S
UKXCs4r6t1O9ONa1SAJJLxsvBji9K5Nzx8QDxMuKynJLugYMY2rVePbP4+/27yYV
LWXEMWXAlW0vw7OvNAOKBVSHKu+1mdjHAwoUlDddFRRRXHDqA7nbcsPmjNLnXdqN
p8c2muCKBKooOUcwgU1SgjzLbQGzry9eidFqsTR8WCDx2vzn9PyWX3hRW1QbCP4r
eActsuCBed7lyWoZRQ41Ff2pLOhi5THBFShyJjF7ScbIzoSYHAGYPu9A+GSGW6yV
TB2FRmyy8oxaDYDX5dIsYUfC2hM5XzoDYoWi62bNG1guBKLL+Cx1snyU3WIsjsL6
E9u5r737Wrnv5TrGKzaL4J5VFgLMpkvuiA/hRt2IcSladFE/1xBwBkOUOgryfQV1
2pxbSHjEQtXMU3HtI+jjDp31Ni35BNpM0xd47hJr8tEWErLzkILMoQfE5nr6bCv9
V+TF30IScJUM6YXCmkFHUtGCEM+l1YL+HjOi/q5UfExnBgDSzJWfMdTkg7TaBg8t
dibqurv7CWMG1cdo1e8kCrvi0DLmwgrv3RPynwJGWOrKBK+WqaOSz99j4+4Z/VNm
Pc4tIgO6J9rbNU2aQdJgOijJip0toS+/8TQbzIGDKCZh/y2XktOBsEAIXGB4fys1
PlHdUGsBsI27pJVDSc5nf8LgL1FytK1A6fKGVn9evJNdu3kv3RlFDf3znW6EUx6O
A5IBNKTWyziv2pdWGcqowrxuJFE013y3heHXH7v1Nr56iBgAuf3IAHDEgY8I0iKT
vAFbnA8Qzlb+HZdfGbQKUK1utF8/PEfngRZKHCxtwQ04A7fwvAk9WsHCXt/vdNp5
mcQGXhQekuMWZkp6oM/MVjdh9twUd4tfuEUSF96Y3gt8am+d+/g+FKJy+lqZ0DmQ
4VD7/MdxQRWzsllLR5gqVRzKIL1La+502ZPHoOziKhniEGCRiqyuTz9d5enYgZso
qWqv16corAEswjKEgiU+Y+eZI+7va2b78HACg6F1JNfPp9AS0FSrCAyIfRiL2+MP
Ca90cs3lCqTLSBYdkFQPxiPNxubVj4oOvFWT0VhydXPXYoEn7+MZQ3YoRAaKFneb
HRaYo264UVyKUGv/c0qfxp6XWRhTIGud98u05bYQz00MLqQs5fvx/h1STSl9KNOC
JzHlz70d14GMVIO0DvCOwvq3zplY/ZyMp7Dk+gv5DYMTk/h+GRbvnY++6OuuC+K+
oKuxa8ha2XNrWJhx71MKerl0jponnGOGiJlR2Irm8pKuA3dhvneXxobnl1iw1xE+
5phsNPC2bZL0+tm5heiVQ0AcVtTkiCXaH4c8gxrub+SIzKRVvO+krcjv4/FtudSJ
ddaBNeDKSFLJ+yPfN+n/XZ8XffkCqnOx0Uq2nbkcZI0a9qc1LIbQKa3sVimW/ecy
v9pi+CJ/avWF916llkuOHe6cNiiicHpiZtU4U7OVgMEmGIbZlIgPzHfi8VzlyZPh
PClOHLj/dimS3ND0qaixOza1kp3EYmaDvuDvF8A2943wUkADJedMNDB5VImDa9A9
X45xIBqHWyLvpCtj1cDya5Sunk+nJ/ADL3p1KEiBtKp1tvRiTJCIHVXG8XomfiCS
S9skrlQ+bmcptpjOCYHOIfx5LNCncT4hYEC1qS7SI+5MGqd3ZqoBK6wrUzBLrKHC
qav6HkoglfJ+3Z2XdTz4Gy6i2WUtVODWWWvBpTu6AS7DPxiFpwo28fRVwPXgWcGT
PmSnDcWJfJvRCEl895tVyJEr2YOB76fjlIEL+H0/7zOLpO9yYgON/C0DHDXdT+W+
U2IFThQEXUVeCdxTk0U3xDwfGG4VfO1GrLiDaOxdKiR+hKOhqhAVDQhl+UpibZxF
qK9/rhFWp1sjvsWbqwPd770vVJ15xKzZDAqjfIo4HtEIP2rr6cjKI8SfkFmgRB/2
CxWC6L1GNaYwRj/Z1ZDnHVWSjfwGDPZOLthvLE34aEYyOMPr0TJQ1zhfRC2luXfD
VsQ2Aks6N3+/SiC6TDRR3kOdnsg7GHXZy5N4zhYnXdU6EnajZNOrXuDiNCs24Ym8
jrPnPbNDeaDN+L+RK5daZyMKV30dbDIKhmeoGb7YvEOS74i2R3vvqQuD6wyI6cGA
xQCsEic0Zwno+63zPzhUePPbiamGYJ4++SLwdozsobWcGI02uAAzFG41o7fcsKts
SSCwPUG5ILhMWK++D1l4lpl43OUCNRZmmERDLuCzfIrCDmzUVonWS8Qs/wsnnFmU
lEDhFPXDPkfEqjM4a8z4PCH4TwMmoSMsJLovMcYHMLwFXPoqPxX8+N0WIzrvzunf
+TBkMVpNpyKZYTWu9wRcW7frC46/1AbXibYJZYLaBEVuW6yFm91skz5znFTUr69p
wsYP5htDOxPm3f3vvVoIIhR2OSrsDl2JHwwBJU7enMxFI+nF2VYsojxhZfnvPFfZ
tuiAm/F+a0mxxS6INcQFmWyqulekLRJfSCDkF3RblssdDxOMRDvKlL2Vsh0mir0+
K6ff2NFy6Hj0UP589xInQwQyI6/NiXpW2B1hkCde4JpaVGwmBtPe/8c7eB1N9T4H
doV2YTpcwKOuaI/vmfPbBf4VzQYBQCO6hQppwYUR4JKboPi6pQh4+sMeFDA2jNny
ZZpt5d+iQCS0M1vc6KnIpGBR0d9JeZTf28ptOACC+4bocFofhhtgX7MIvnQsTvkP
GSntnCj0c+g1iBDKPNSfuJDuLAk5jrxMGuHT7cuwsmvk1E3XQK1xi0L949+VVRU1
S6Z/+V3HL+Gw4v0kkHIMh3th6Kz2BHeJB2dDhHVKQKM7qeVuALxb6YgEHOTRBZDn
zB5/XxAkTlZJKbMsrBrN3NwREuzyRvXc/XWyBotR4VxFK4b6xFGVENUqm57jt4w2
CUdMJTsVYQ418m0qHKNk3mOfWNB3S72MF7ZDATfZYush79AygQCMnmGiJNVnD6m8
4/21ks0x9ed/yc3iiSv7jzO4n7NAkIKswLjLfCFFyVA5SvJptuGbt1f+ThmL5iId
X/Kx4LypW5BP/sZLdGhfH3vHl/eHKHRhPkT44JI52ANtktik8xXojz568ximCjJ0
Xt4P2PckyegZCmsV0uwFfKc8h71XV4V3lHi8W4CMOrbpzhoAML/9DHjAO44FIg6a
NdQMVmr2iKWFi5nxePwOVh6z773oDu5aoNwiTiFynHQE4Dcc9UrFhVrb6w2yZ7dT
At9YfP7b6lHIzBp4jygW0khhFpOwjj8lvvM6zBKgKGbNQAS6WdoR9YjOEw5w8TWZ
Wxz2A0h+N0aDRL1xhpBqvpGg+8DsuCXLY3VJjZcQ/tmB8ks06QcdwJiLQYgGmWYg
O+N0nRjdZZaIBaEHH7PcmFttYDskiQSnn7h1ad7y3mU1NF2bb+DQxDD0Cy18iCbM
vWrxcRV9GcwdvgbpXGcLV/8KBBnIpAiMDtjPcvI9mgn+dIlEX5IZODcisXkaOOlD
Ge8sTcArUnSEnv0Lqaex44vr4H8H9x6/x9r2RFkkVNNce1uNb/pBeoLdXFRsDr/Q
MUKF9nJz2L9W7txnjNHkSQxR6VDFDbFk//dfuShw80kw6spc5n2KQFhoDlcdGUEU
4XGcoj3Aty5VATvFGfq/2zN01iDQcezjkrW4xNaPqvViLJJspF+ychfQg/qDpxmC
0Jr9jWYcp/TnW7AsmM3uhzYMd3aY6us4PE9B+mW1L5ixOlnjM+txX7Uh2gGgH7WL
hkGSIEtlIumr1orzxhnwy0mQ30Nzja7mf4P8C3JKSmMeWf7zjYVmi7d29qg6Mr/2
ih5EYuUspn02VG85Al6+dWO2xGg8/KA3c0WaO2F0LGL2p2+5CdJrV27BaJxAmczO
09HE4OMq+/HnVCf3qXDjqMi9TqlLTE6gP7YtoROX9vdHrulTF+gCQt8y7qFYvaNU
iGW2wszbienR+lSx4gP3nfYLRDJRL4Z0p3UtK66ZwqVNszhMYVB6cELJz5qFDrgE
MhRJtl2/wYqBiLCwcaIpYXN2B/2t/muViUwvc/6y1XWC6fXMzsXPMxqH87uekNPG
HAwgzD4KHbV0bG1uAec43PY5wTcHu3K8/PgY+YE2ykkHldXvgFtmIUUleu+LTAq+
91cBkrozJ6hdRhI/satdyY2KxjSo/CLahqrzGH4isDD37mVHRvop7txbwU/WQDEx
3WjhcWInDhWFUvRm7OH7PdDOxIuptDcXpzROwcfd8lFGeYG2/AZDjMShEd4LvBkF
2tTjITNY/N1H0WCajyFpLiAsZISscV1iZ3QW9op0Lu9Jv0MzX/KtQLJ6dEX83Qet
krNyqS+0jG/4n9S7IY5suXYC8WJwnOTGnFAkhzm0MU24GKPjlOf3pzqOQw3L24dk
Rp8jJMVbpFjb6hnBjkMe9kGsM3R1q872WX/6wdE8NUbWVXnqTXi2Rdy0G0LQUvEa
rVRRXNB9cyFB9I2h7+TSGURJutldf4xQt5/Jg0Qybms7dS2Ib/BiPy8LHLyqE2JO
FCiS4DLlnlJcWoQn40vylAE/q4bhn/rDhbR56OFt8m2OVzTrbA1K4xMk95oINZ1d
GxQSKV9uMO9EFPvm0prHJ2tlmPxy5j9pggsmzxp4ejFrdDVMiZ2WYJBo5TYgJEiE
HyxOfaPQGBO4FEUzgxZ9MYqYMWGGdwy+dScmWAdIXmVB4aLdKHzt4O0QpzbyWvW0
7Q3JsYGWVfoB0YFGoSrBE1mxhheL9pSwzghheitOYXgWzCW5nanrYcPA2nJwGDT9
R9Kml3I7u4XYdUIkArg97rq8aLXFsehtDgbH42L7KY336f+mFGouap49cyhJNf/7
3w7UfNxfmBQacjXZ1g9QUnPUfVFC0vQMyv9cI6+7GcemuZSUT0p40PO4qNqQCcRZ
VB0l2KQv5aIXdf2rAIWf5aniy6RZ89wyPGKMDt4NwytE52xr+IN08Q4GFhPDHFQf
LtaCYPhsaDxOsUiHUkbBz8gMf7WtskbGbHtSjKbH/QEyQtyoguIAUU2+/vbgENrj
1zUV00brEnOwQ5eYFGWByEBl8IGarjszZNlOgRmtVDv8+BxhBI76Y2v67lQ2CuTg
W1pfk9HBIEFy4WhVJVNW+NW5NbYY4ZHY4X7HSiF8tyXBPmTECBXfMXmrGT5TrmUg
Gnw6cxEH9GaN1olARBSThKrB+DCw7cgG8ApeB6gnu3A0eLbucF16TBymRnxl0rdK
qdjbBNMvTC6IV/xfFM9IpQjsajR/C5NyD/+hO3JRTKZUbPmcqJrpRZvxnb8mu4DI
FyM7HVSoXK7TMQeg7CN1GlkJbUB5erQfY77XyXbPU5YTAgaLUxrjpn09Pmikf/cr
pA7aBJ2P+mrprYFrWL9d9Uv3H2xnIaJmfZeLSxUbaQ1dRuc9N9/Y4bQThFzyfqkP
craEu/Ogiw0pADb6I/fvcHvPCKIwdkgng/ZUw3ayUXKosiJc+HX8wA5i2AeeDoBH
xNFVWNFGvytYwa5Mk/PSQnzvPMHFsOZCOQm3Y5YctPFvMwPbYbn5xBiNOg3OdfLt
MuADlNCfl2KY0v0V/MAUA7w0B93BUUtSQYXQ5wK5kPJ1iQo6RHuYveOCh0daup7a
elHQMYgeXd1AfEx8Lbg2zYWJ7ndofzMW08b1dpNevFEN4mRsfUM0cSIVji24mq4R
5RcuLjDheE6CkmEoiAGx9uR4xeP7JlTg8I6GTmk1O4au7SWYeN4NJC6NykmVnGAx
hGrIhw3HV5NOrSN1AqXEMgUu5BTmEow9CGZNi60m3XYYRd1Q/cL6TxqW3kWqj1+K
xOl6dhV95STTt3MF5HUOgj69bj1roMEUi1Kbr5t89A1p4O+8KTF0vL89CnuMch0B
oZXDZIqLamUHqhPBk7LfmDoumjhGka9mWnkNN79J6Px4pwyqeYCjPC+bFPEvzp1Y
cu5M+0SvQxyUk8cMNiz499eodn2fNSKmmqZsC7gJVhEiqEmRRy6ZAfEdAEzf2G1x
T+nuXnX0XfC4GPZAM/NP6QOPYy00eOze5TePg3VL+hPBZD3yOhHrBainwrIuiu21
W/xspib5bZC2OL/AgB71nFYI0efEJ/x/ovH/bzyOA4fN81C54SaSKqkUo4r583me
FMbMDi8qGSsJrdJ5SqTCfznbrP1lIINdXSTYCzEQowlR19z50eNRTV6sUxCBQCo/
BhdGZrMg4LSVww4AyZWhpavpu29LQbLlHiwLA5AiZVQyd7Om1xEAD6NZ3g/DGPtG
9U/WB1GtKKMoIeNXb5JIzpYMNqdav+VlfLadstrxjm+SS3tl+Rd0LPe19pWu3VhK
1ztXT4IGrRRIHojPT4mv41L5d2JSXnLgo4feuAqJW84P6s3syEV+lLqfIb9TtsPX
ecdKOGldEZJf7RSLxr+aErfTxQAAWqIc9lg9ildDw0hAg9fzlN4xp1eM6LBbj6zi
AK+OqdmLJv16bdExpNQ/kEpxMf6lywNOhk0YtaOgRILY6kgiRsuvnob64C2UxRkZ
+0m9VuU487qbqI8vcPR/77G49rk76YETacu4CIYG4FciPYwFm8nZ5DaxB1b30z4H
Al0IEyxzPNF81srN/6l2KDxysl7JsXuRRlW8pkyzxLpnULOnJd66Z8SyEE0+EPfO
9M+b24DO3HTA45Oo0dBYUY5ahovyvm2Kfud6HdwkaOkwNg8UGLZeVOYs5JrsLGJA
C97ZzrNn93HlVt5Vx0og8rA9uKXHCYBKa+Hwxp1TQtCO58w8ezroir1R0BUATl9O
+1tUgUTwUJUlBGuA2/sDViHrX+Y/SO4HeXStAvhDHXN2t4cJ6j25EaxxJ7Z/GCJs
IWRxwSyvzURzXNd6+sfTtH7XlfZy8Pi2JOw+oSLfI1fQ50tLrRQ/fSBqdqDr8SVG
N/vDomDspc0qxyQ+uDSaq1V5fyv7xB3w+zDgEYRGTprh0h3SLVjR3m8geiJY//Sr
PzTIEig9g18OIAxb2hmfboy8KRZuTvkgVnCAGZb8BDOi5f9X43nfMM1hETXFfHqv
F8CEsMDyqTEEpugFYDVt7TxmYrwF3dBjm4kqPZu9ojnT91ynOaqoK6hqP/L9SQia
PXrCY3odB2YhLaZb63KrmIHxj0gXWQjAFMpzKKHjoVp9kp3WbDqxMH43S3fpLC6p
L3PuyYvx7LL2iTPJVLS1vQCY/Hcye+p7oziHNNcq+hNSSWHmrKHle6E7oS7rxYlc
D42JXxMeoFfNynBgwaUizMJfehA7eNcYa/Z3ExRgPHSbWLNeXtrWP70107SwJMr1
J0a0XkZY4uhraEi4WWck0jGhJE5mgIQitkR2nv6opYI+qbLK00CBgJLMfnyYB+EO
F4E2Ug4LeMf7i5Y+zY04UewflHofic6CmTh38rCXLI0vEkO0fE68pVQG+IIYnEhE
+KkwlVwFf37Yvb9SlVXRz7o4udslGtCcuMdRBf/H2hSKNLTJQfbgy41UTg8uXq3j
FnpfOGlk8OiqRVC40iOZM7yG4MxkZ/1ElTO+phVcgWt2eAzugSkji1qgCFDVdBsn
xdMJGa17bQ7WGJhhUvMIbu46cZAYE/PDiJxkreu7u0TsxutLmdHcohUkLJFcXx4g
FtUpBZnTMFRRI/wcpu1yXT6f3es0sytJz1Q4MCTqj83GT4mtV39klWB347clTySu
Noos4d5BXYkZzuHqxwL1uxkrW8lNqmF0VRIZ9Kcb5e3JR4RZzJDxcpGxiwkSy6F5
2Km9PP/TkCZQ3ggM3jHeCi7YOZrbo3Ig6mVnu7iUYFZsC00oHBkPAgmYAdG+ODJO
cWADm/DRtFKjMEtlTLfK8uVCiIfsQSfj3ESBYhzgQ5xDD6/ks6rZB6KcjBWs963d
ULAID+KVTBLVHvfpZgEhsNAVSGOQSfl1yB2SLAtWNZQnn/d/ZH4OBD23Vu2vMnsK
pCbGlRnUCVbXW1LPoMsrjn8gRi7eV05/9znL6thom2SmFqFhIBXJzUzqoTB1vhgA
kFzDGoOX6F8xP1Xd6tqCCowEeLu3N0bmi6jyrVHi6Og9G793YJMcTeqo5fRov2xU
Rrby5/bOOTyALVoG2yLRoYAqmSbHJN+OmKJ2/kab8W/Xbw0q5W8w/1nLEghlw7wm
wrc5NLwJUwjm1u7UyO01hdv7aopcKzYxblcVbER2eA6XvQZ0HQiZ6UcFFeZ8LpDL
I0V12i97O83M+Bmd+5QnxlJq8sI7bxhKmv1PSqCDnmkKsKBa8jFERshxy+1AiGdF
YLndbaykybRZzcB+uCR6mReR84p22eNAR2Xk6n1au/wFZ5WHTFG2nEd2J6ilZiNh
GSfB5MiJGM6fUBUa1UzVAZ8rylc5QVmgC+UN9KC0Ucdm4lakaTI8xxtYAVZwXyN1
qRgRCNYCGStZHWEjb78n1CyjrPxkxLXqZRnReg6xGolbcANZADgIcdFVU6M6eAIn
2vwiTWNCK/N9XC1r/iXKMKQS7yuePLjlZYk0H5L/TCFma/3FCcGg+BCjfueVV47M
cbq+U+YpDe5qiM6AQzql8DG1SK+V+Yr99Jkk0Ofvofml4US8MUi4e0NXwWoNaGLn
wfGAa4yVYxQCxPpuOJszGochlhCML/byaLbxZub/qOwrgjRg/o+oDuCmY3qRjuGu
yg/MTo66aaYCAWrl8knbTmt1g9wxDnENJcLoYygV9bqiG6ViKEEWnf4siAylAR7C
XKxF9277SeLpQOuKFjw5w9KaPglXh6WyBCRz1DbzUHLfPX0cogV3rwhOzPn0zpsL
5Yr2/1Jr+tuZsp8jHDtOgduF7dVj+e2ugwkFzBEz+jjNjSQrbGGEBzzovMJ32E+k
rWYhV+YomCRKlUO6aBtntPoaxw3GrLsDA0jsd/hnosiqan7WO6ZKfuRpB/NigU82
n1FB1agLzRl7pKzH1vMWnIVC6OQWiUB6AwHpizRxdmrkEMUsXnoCxLx+OlgpshAX
SufXGDiJ832T5xo81sCLkpJvi2KNtj9hLo/QPt3VPyPwqT6h+dXn97rYqrvKBMsK
SSbMSmPcdMSSLjaLDt9oTWiWBoZQbxz2eW8qeozI+eAxStf/1n7hHKnLlaV9AIRJ
Roi8Paxzb3rMB7oeNUQ5JRJH91Nu9iICURO5zSuoEFLH22FoQmufwyhYMEh1GIpR
2MheTrCwtg6JqvXcChwHT50uwfKUAIs6Ysa8wzaha7XCurIQKXsmT2dV4iKI4kWe
ZOvQs5xegqUQf6DkbFaA+J+RcCCCh0nZyGEATSfptxKureWYUGUac9P7OCf9pXjd
+Zf+zrkbg2xYMTK7o/rDJLZRBEAEVWHChn0Fgv8gHhqZZSNh7OqkfyfhyyMEz6cb
3rJYfQRNOO73dKeFP0LoF4twipz2DYQCLhAQRI5cVYZh3hQ0Cx4lIqhPPQI7wEXk
FlcKedeDYiuw+MngIemK4OSfMihWtphjE8PIQRDJvwIYX1PEbR81jmk3qtKOtcoP
jwJBCNW8YvPpwlXhy4NN6WZyi2i0dLpm10Gxbo9B/vvMInKd0+IzNxcX/EOn1lc8
m6GOMNny4sdy9jWkPv2C1zY5NJ847nw8gDjwFHRDlydHnTaaafemyIxwHfmFWvdT
mp2vbqniCgUQKkkoB2xMMysc5nVm3RIf1VCZRc03bwiLeI2wGTLSJk/cN9diuGqc
POVgqTNfZARNRjr3BKKH3ZUl5Bc1JwVb1LRNE3MfNzxnOBRskRmMM4M/R4uv6MDr
nxXK/LiG6sh+7UO1gF++PK3Myp0hMFYqzCPdgsPyVmYRGClo3xOH2qgX4LaQ7axf
0QOnQVPtcqnLwSpG/f0fqHwx0RxxcGvAL5iWcRURjME/lkWLpDxjUTj76IXPelZt
9JCNDWKsq6F+FY6o76TAoMRO+yqJWgWItHN//E+wZ4mTqVASay6WZT2YQgzXxfN1
i1XJ6hJm3EZDtMxLOr4ICYmRvkJoXivwyKLo/20ZO7JEiXsl4tqqPMGSDKuIM046
6ggm3fVE6Mbj2wLXCjs+eQ+VE1Umi+38aW8djVZbqE8u+0AVLp1TbDnS+vuYL/st
m5IRwTdAQklfr6Oiqx75Us90TcIg3bqq6cTXAcY+F/RLDtOY1H9s7HBFF6o6qfNS
S0ezX1CDflw8Z50Ifn3r5Az5oMYYJMvG+LYQfGkYyEX006hoHlBGyO44wMOWebvN
+jMOwreizKiP0zG2JPaE91ufKiTMDS1ZrJXD6m2/PuuyrPjIzvbbYLNkZ8NmZMWu
PqAZ8IOcV+M2HHxelG+7m4A+73Rfhh+kY+mIIuDISfLxmlvuqp+EH+MNhkxTPegE
NS/x9eT0+Ar29c+0S/4Z86J1HWYrUzr5IsRReDiddOVQ0YinMH3qL3SQpq8w8w6p
mdQ6R6p/oS0yXPj5xYOOf/9KM2gOs+NO9JaJy01BYzWaO9aUhXAfuZjop8tQPjF6
9SI7Z+Re7Fm/I/LwxFmXlmOJILXU7xsvffPlO12+AV8xrM+GjLre0K8LV9ceaXhY
Vp0Ii5zuimGU6vx99SohLZKyPntwJGgxjeXOWR/GOTdnU2joD/35QIDVNLYrjadi
qbbn3/iO2VebySJFS2UnHiYj6JgojyVMPK/aeuudr12Mq9bMXF1Sj8bhfLcNohYb
BPX3NYVRn0UiOXT8IlEkrqq3C9ygxINtgENnn0JD9CUDjbEN59/wOgNxnQq+anl+
gM+eqQBNeltzs6FJPMosziusO8mCqQo1o723NZ6ts3hNz8/yz/015xngF9brsa28
EPCtopEE9ECXHO2AVF+w7rHYGITmoi3NvomjaG3mDK5hxluFv7qDURcea6+eHs/m
dbjXT+y1hul0fHbw4lqlmu119W7HnUFEFCgk1HNw4WRuqgM5UV7wN5fYteifmpX7
RbeouYKKt4rO7+wSi1du+3qetIOSovISlV6TaUkRtlVMqbtPzTB2Exftoe0qBQI8
Ha1TX6FxSc2WDcSWXuKQGosuXd8yKAh4g3xxHAQ7GTSDmFLuYkuRzdSUn5tPfUpt
xdr7YwwP5ptRaOvDw3kl3hYuYhDbGheLmFRovz4bEQaKLcAPIHIH0+1VoJuQjZ4u
0r18IsQRIhemV7K5YD6WYc1JYJ7GJmfPNb+x/e4zOaKiI1k4PAn1NjVSuOeb6gzk
mUjmeRdTTaHsYIrtDZ4sI3h3U+Sr8oYY2qbP3ehabcMXTByUNGrMbCXwy8l8yZxB
vI+zB1HNPufWj9LKlN/Zy3nEm7Rq/t47sKG8nLstbgMofRnKnyq/DvFAczLnq74E
onG10eKxQf5EOAaNL3v/Q/rMIKcqzkLzrgsKTfx30E006zqPNNJsPFqURnvde6Bm
wE7gefGJ/N6EzFqts8L4DmNHu+o+To/g1bJCJR/6uyiHNhf11w2KF8vBUm6zhLNy
Tiijtfd9TKMfGvs3F1LNVwiNEp1/MNSJRZkj2a6AKLiCkhRVeWVFWuIPGxoP3kiH
YIMzfjTJnIufw7DQl+/9Fdt0ueijstW3VE/S9bFAc5z5/a4MULSCdRusN2s5u+sb
dbRM/bH+B2ZezQK7SMTuvOGT+E7BHDAKYxmu//wxx5+ymu+G6tQoZxKhSq8ViYJN
G7ac4iJIjcmviIO/W+OW9K1jV6yHsgWAruLKdRGw3kUPsd0RK82+N9gkxIoY4lw8
t6h6uw78caVExwvspNab4Rq7WWKuw5tIezxFFCxbqBqZG2S9qGQvSPyUpLBTE2Xr
XNxrUW91qW6yll6NO0EZlKvVkMhR6Zlu1wLjzcnmJ0eELEtc2rIVuUfEF28gjV3h
hvKlmn+cXH1cAMBR4CazNPbqpUcPtTkNt4Q4sdH+7XfJLI/Xc6sxqNV5hL12w2IF
/Dh9/clOuGE7e1WtLko7GCwjZqKgiGUAfu65Qkls7TeuyOQHf+yhgLYPnzSDPvqS
/KA7VnMBBXvdy7B+2Tjze2wkTisolHa38etXdgRjTVl74k/4MptT4KpChGyq87bw
cKhEncbVx38vPO2EDa0Q7lamZ/PbVfdmjgzE7PTkEpXbayl8XcP3BwyCxgWBjsu3
dC0ZKOjK+GiDxjyllAR/4UBuwmYBEhfA05hufgnpqmk2Sunp6/ILmlG2575TNj6y
eLtGfyIn6M2qv2vQflIArAlv/p6KcTPAz1ue3a4qj8pc2Z5AR4KSx+GDIHCgR52T
AAcYLreJj9GKTFuwoFAV1zoh5s3u/+5fNw+7xOVGNDWTIc5L0H0xMV8X/nx0rOQm
RetLbjD6A6/BMsh5AX5evd7MSnZypaN9rsimGJi4xri2dQX31OHZFRnDeQtvgFbK
idhhfEZ1rGmErXYejgOYJ/e8WR/Mrk0vNYNOocJb+SxUsAaZa8kowgoWU5iVSopW
5QjZKoY5CKPIfy6wx21sOAkI+Jx1hZsztZRoawIu23Vviw7fKDI8atI0//qJZtTE
o2b8uqEKMHLS5ZzGx/jdPIDRrJePPDdl/Rw1rWDepEAz1Qdy7XzwBoNAFihoaKAE
IQpxpf2qZT6ijf1D3EJolwvyJpNpuJieM1kiFCsREhc2/77hJDrZ5SrRRIE4I8LD
8wlfPlEYU/29bxg3YPLSjRDJ1cbct75o9owH2m8KkmI1d1sHkq0z9SP3jHxkN3FN
XQsHFY4zBPd5hIC3xOrnZG4D1eXwnovezxs8bbJHs/RPO3chRiNvPjWmXh96vSMr
RujckGwI8vTifhM22DygGltTmGZ2Kcobqfk1LOwAO6A78ZgmYpZEsjtXUnPAfaMC
dovzZ2hixKMntzCUtVVk7oQynNjgIfPA3e6FpR4XmOnd8VyMaueMi5q41M5hqUye
anroafzIOY8RTTs7LzvPsPEKWyuHXoP/kd+rfj+NcYXu9rZ9RaVPKb+1DQrk7Lg/
RYJq5enEaFNeocrLV5Zz2m11qsuNPfIpB+AmDchusOM7+6pf0MvISY4wqUWtAz4t
apllJA9rwZR9PzSC6ykqGNktBZhNafCSIgu+6vBXH6QPWizTsDdkB5rDrGJMS9BA
elBmkeS/UCKK1HNi4DmzJofFnXCube2HFWjS0nUwKjY5vR37kuQlXAi29Kn4pYnC
GDbKrzcfzIwaNUYmyIzpcGwajo8wU/O5Dft6FfEGObfj3JI2i0ATqCCPyaVPtsd7
jy2I1T/K+1gXUwJl4u8btGSaXrA5KftmmhXCuO7zl2EFBUPcY5BKlMfdWZiCT2a3
Fx4e2KYVP9/d2xobRGCi0Rei62TUIgmlCsum9sGbiOYd/sUN4zuJBHJRXEkoJx8G
KRxdN34iaj63r+FTc22siWjoTHmiwmHT7fhezhqBdbQFhECEpE56a2GquwWWi7Eq
NM/0ZqmM1yFgQN2iMVm+gV38k0ICyhP/unDApLqb15IuzdRp4n+x3QG9ntbzWLbV
4TnvZcD+kV2FFZ5xjxlHz/fX3YHBE2n43FOi9gbslhWi5o38yy1doZGcGWkE4SO8
o3nqFSaUt/UemxkKW17gD/84aqBduZEeq7EwB5dPt4d5dpGk9rglINkg6buqZmwg
ET58ytP3HrN1mJ+AByGnWX9rlg+hFb0A06J7v/A4/i29SxhQi0odBOsYMJmTpPmR
9O+3+cp8GSLF2NfYqhZd7AL+egvvhvlTtETAlFrdMjmy8pieXyqw/sv9ZeVUmlN5
ffqMcfB8WA9ZoSP/ARi1wIOKUHtC7JpkwhRZq+9Vnpf1DNnu/TdyXU1ti/w704g5
auk75KR3lJnwEDy0Tnjo40v7YG88c2j20BeYtFGqik7RnCAuESe++8cup9xI0FLd
6+Y8GmYlIrqmJgNYAGP4VwZUD1ZBmWldA9K3CkXT9uG61vrxSJn7lZnUGIKKKJY0
F7HgRKOOzb9xvqRiGmWWtYBrpRIroBv2d+rv134qv3MWuL8ihnOlOInWATprJavP
KEyJwsJSnDKYK3un2aJtLWrsQ3EVpOgYD8REb+sncuU6g68IkZXU5ivVWSfVvzlO
EyRCTJGG8rKMjTxuA/v+uwTJUrsBG5nbFR+PVU1gfmuylaXxqNdCJx6BXtaKuCfS
O2BE8wDI/1+tPpDiVinvn26Ho+mUypxws8Bsry0WdGnXyBe2rGkoKdVrhXUSObOr
jQo3b3Tye2o9boDzoOSGQTG+IayRKlFpojKX7z5O0FDDMyoV4Y8aoUPtbPFSQw4Q
j3E5JU+ZrPKxmv5h+cHuqDZ+/MeN6n12YR1ZPuPbWLFkXqnHq4i8wcHa7uXPDqrV
/vcDU4vCOYQfjL2p90gG5PCBpBBl4lVtirga7yqzDUxoF2khv3tJ1Nhs5zDbXVQH
L76mjzAqEmWInyXUudPym5g3MXs0XT6nyXWKbm7rmwuiylFMn8/BWm8NhOtbkRZ4
7XrXn8eqLb/leXTNwPDyN7w/cgssR/jBJI0wsj7e/VRn74CPt8LJho903vir9lXe
m7u5/wyiUPy5pCISozpWomLwf/n8D+gyNN3vQX622Jaxyo7D2/44tOhU0//CupXo
LrW7xQS4OBZv+1X50bUAtfc2yxIQntOKVgk5b4duWBSFmTBsOAAyxX+ASK9CvrX5
if/H0GMjLyDqFbsfz4zZO8gLt300HPdq2/EQqOpeWnOW2by2JCzm0Bphl4VUevui
MJZpadoYqaqZo7Cijqg0ESBBZGSmXuM7Ub7+GTejURSKFoMRag5ttX4jC9IFZnrw
+rmuw5t7hiZtq1IgIV7FIszs7aU3Fj3Bn2xBfhCQPdURjOm1MNzCpXbUXd8QLtc8
eAqZIHLeGJz4ustN9g76DgcIMl0WPRsEA5wdX8FtxhSX2ZfvDgQrRQ2xE4LYaZoj
1f7he11ffVGsz8xa4nuynA7OGs6HF/AifOgCWonJ7YlFYRc1Gd9oBVO3whet5YrV
Bvuio4/LGg+O/hSy2siSel7zKs5QvMGJFfvnuu4rCdak5MdxS6sQ6KIy6cyzws77
qKmSJ16gcE1hGJgkrSBd5WP9JSlKgjcKZIe7CYoKdgPVubojOpsIV4SldG0f1Q/d
CSuL5OmeI39AnYMPu3z5/1WqARebbsS9NrFbHIQngXlxGG6pNbSuhdnWaguoMT2Q
W3SN66aQIAOfG+1wKhceuDitKzk/gUFiDsgKn3YSpXE0t/LUEgHYsNGzzqALL618
qa2A6KNwv8RaIiMiD/8RVzdtGa+CDG0M5YDVXc75JhX8DSBk84M7Nxu3uyV7BmfM
9itkqm7DA6uRR1nSXFp3mBjevvTYAjAqqiTxnc3qVvEC8x6OkylmWaHFyP+d7YFE
pXhexJJ9hIWWCzeKPfjmiMjY349VPHqZslsuxgxjNFF87/5rkAzpZivaXRipYadr
GKev8r6pRz0JdQOJFAzXDzBxXSYs6zWDngeI125+2WJreOrqrh/EtsvZ6fZGwH/e
SDiecRW/i861Gjf2KQvP5pXmrIvWu62EmpoiErQ1qlp3DD9dwo2gl493sA7DABo7
PFVxZsFIqJKb+gu0/US324FlQLz86Z6oGZM7s16yzD4bBUmTyqCHabBD2YP8DCEy
0NzfC4ZuKXgE/QKBUPtPnN9PW+h71sghxAts/jisE1JzYG3PjQIS//ywVvvYZUEx
efKuEcWdEwaJb6r+4g26mYI082YGOi9jtHMmVssSsgsW39sw2huR/7B+0nu+hOko
oltgHKMU1ZLiYlUkonBMsj282vNxu/DvsWDtvUVACYWyuRY58NJm/121Fj7Fc1ov
v66PrnOcVdfBVj+V9ekOS7Jztkb76XCcDk6z+c1whUNGCHdUX128ss/uOsnQZFC5
jLOzjn4cC1JaAczgu88n4ox2sej8yFOh67Rgk26R59xFcdAINpW8wlScAcLV9r5K
nF5VQ8Anxz56ILBGbR4ChtUrS3VDuice0o978eqz98XX7kcVRqBIiWEDR3ZgPP3a
BVCtOVvn/vhbYIIQmBlTdDklToCw5Rz2/8N+/xgLyLboh8qUos6a177TCm1/EQDQ
ZmXcM3r+cjPaCI6ljYkyykso5ZYZOQ++C8QAs5EbFPDhZTfO0aTvZihQaW/VpWcW
M0i7vGJ2p4PzW6OAbJ4EwLUbVkTDNnbSOU1CGC0X+p0AZ/tB/vunNzK7ZA/cG8rO
XCYP34Eym0KfwCjMryqkBvzpftjEo2xhl6gGsRj/XGMWerAVgik6rJTpHJ3oZ0Jb
7fuxc1SRO/eQGyUq0Nycp25Bnpd4DbmNboIQCwskkbuqZeKHwDSepY4XCyYDqjXW
Pxd6lw8AyQ7SVX6dgwYSYx4ZXnYJ7WcxZnDyr5cSNtypUS2q5FKTAbMA9+RSS/lR
eJkefCqNhvvjFOTetZ+hUaaSvHw3+CO7Fx92DEX36/pbsADraFz41jPxJDpXKQHW
avkREsH2BzHlYhJbqEIoLjoE/vdL5VV/4jdxGziBIOKFp2BZ7wiL3hzcvM8z18gm
GoqTzmnGXRsA69zPqAO4PnR5PNz3c/CUNdF/Gnd2C0iN650o65oLLBzbuNL0Wjlk
BVCjAgcpO8ixvSyuzx6LvvansjbpqGTvTneSdx/HeT3Zt6mBEKf7K+1grx8paQOs
yaSBx1qPuA+NMrdOmJwAzCQRoAwoxugcY8eDcEbnBEuTQLxXyz5xMfU/NpKTTO5n
PW0A7RrF+cOiM4dOkHQibcNLGAr7eGdoM6d3Ry+u9GY7B485HPi9fWRaj1pwvmBk
bpnbqukKbmmFwuNp36+gxsic4qOAVFLyU4hilbx7VaBvIW2D+veiEU+mOmu4ybz4
JD1fhqDLBf6ESfvW4DXc+0yZsYW+L2cJFhP43m0fLqS0kquzfPhaoAw1d0wmk0df
xOrwbcjtufrxv3s5ra33AeWYv4Ft2lBp8wsM5whnyXW5+DmkBC3kV/6wbwXTKuNU
1MWzbVfIJ5hZ/PqEkLeLcvmC6wXk65Lyb1lOtTJQVoT9ZDhfjFK5qI/vd+zjXyCl
AXH31NZ43PEy9TVGGUJR32XvW6LS2zd+0IEj/m5TCpEoDF1uBCHFHRbBzICqrPiM
/gYLEMM/MWmipNdOtDSshv+l+zQCepaZyPq7BOIfYumrWZ6A5zqLHa9GCR/QC0e4
uaquWaqaZIKhn3IXijJ8Ftwc7QzmnSJr8JIbw3duqHqYp/C75vTOUYAc9TOsaD0T
+SC2vl1gvCdzqt8KwdVPRICV91biO5CrekaZ7zo7zsJ8DvBSks/glTA6/LLBybFV
x1MQ1UeN/OqVVssClRLvjx6YJ1rXLgKWUsTC87qeyOpx4LuuIRsmHg+AXC1zZ3SS
ditHJRlC4fbpMUt3V7/OZPwrrYTjCTLvIefZBPXkicliP4v+aCbTa/OfcRqbhDI7
B11bGjpxDH5jcUb2tSDenV6TkQFv/HN/xe6LaYbsCbTEJFin3MCV/6lHaUEQxByM
DsOw2mNDL1kYR4dgHLMdQAVlgvMGm1cJkxw5AhAaOw4I4lP7HHEbUwO7ufymoowQ
1rVEzjKLVy7kpu1+Utlix6lA15jSWaKlyKJIQ82UEExP3ZI9eYGG1zSrv2vf2pmv
T7MUNWf6Dd2tP602gnuSi/TRMdU/xC0oRJ+8Zymoh/5YJaSYDAl6beMMaTjowdTX
w0JYYCpQ4Ucl6HYz59gfFI0xDh6GuFvRiAXshNsH0CYkpRtYUn2jfw+UozTUOCfg
i0SLArCJ0Y6HEzDcdh6QxVtrIbMUJVodsgmwyYtpk39bqfzByH3BZHxH6i3fxVbI
IlR27zklMmkGt0jOp772py/+ss6tKL7Ln3vK4NG3LkNwUFjCC3/rt3ZpbpYcJG3m
Nn4geApaAAFrol7mtIkSG+X5fMPrOjG2HujwQrjJxaxDVKq+ur+VbbAXVPR/klNV
82oPENp6kVTGPfIGBdc9YpSfJCJn0sKzXbZAGOJ6+JAnKeXaZMaMayvq4UxfnviI
NNDUutYAtRZGwFEYIa34Ab/8QDxmz5E3HOPC4pC/ufyvNC8DiGWDRUCQ2eK6yK9c
bFX9HTHKi1tAOVdA2ni2iY8m1wp5fUlyJoUgqzvnjRPY///fzEyhnWQ3ZUe34w6T
BcSKfSNA4FbKhAoNqjAfgIxoPbOdmLeWtk84U688T7sMrjVlz21eCoG3sUj7ZJAW
c2B9l5hT/m/cw4INK103yo3I8p4oiFMBC4iC26lfXQYk32XhS+Ae+Ehj0bhSZ8ln
sw9aozJ21dMMJiKLpfwIwDWphX5Fqf0ZcsU219/EvS6o5mc1g5WT9q9J7sdgQOCx
b5DjZ4xD0YIQowZtCd6CGg1mooSNlxWI+oncXCvkFeK581OkD3q01k8Tpfu1BQby
ykuGTe/+0FM4WSrEZ8yESTxjYkrEhUypCU+SCRIN9QRYirl0wMb3kZsjdn5uyc52
unBpkv6bJpeJwLR0TH3j/reZ2x6KsdFcmSQuOQQ1ncmxiHgpJzfQvG/wjiG+a7j5
MR8aUqzG5NaHjBI+vKtUBA+O8tkpZzyuXT3KgUXXzcXZKQ2ivYXSwElL0eqJegkI
CKOsf6yEO7ZhKK602kjdIx/TysKd53nxXzMcR4XxJS0mxhvCYSYhaW/yqRjG/k3N
jko6aM9UGHhhicb11fTqJ5F6V9dK/wcQzfV2wgmRV1peNN3aiOQSopyvx+7RTYf2
7lESH+Jh7I5ChTRi8IBDXFPegj9Q3qOARDXsIuztZhV8uqk1J2g09km+iWjpdBbT
TzFYrCc4/wuACrLSrO6EKdAX7nkOGN+HxMzi3cFUjTPDOwch1S+APDxBkYtrMYFU
xDr8FZJVjbPt9A+49IilXfy/c+HXVtHO9UxzQrk1mPJta9W0GezGexpySKZWh+D0
+3ECXaycSPT4r+abQwbrfsxWNZJ3gYvJbhukNbbZUzRLz+miss70WiYbFFESN+c9
5gcG4obCXtKKMaPNrcotcV4rloFCkPTWwrcnLKqTyqSjmE1Mtx/ItyBx+bdOPJUT
mPaZnXuf2Vc4lwrgLotjWZXV+M+9YNkZX57k3PYKrg8bUzPyDN9DsVHPoAbCmMGV
ebJjfkhnl5T/qc1kxLJNM85gW5N1r5BMWEWwSfqr2nDv19vnEnvOqnADgOtsPIJL
bBuHauoaud1o/A5cIXdLnRkcXO3zK5ug86fSstJwGf12vTLP65z9ZXQ24HLikkh6
Cnawm7u1c+Y0RMYaOy3Th5kUdA1BM6RsztmXM+igD2drK0IQMcO20DmgV14ZV7Fp
JYQ6y2iud61bauPNRdb2Rsw8ueNuhj1SrBomX7HLylLDkxsgd2CQXojFVA5+4NlA
8CIKQ81SZebgfzxOC5LCP2+b7OBdNIWhmJ90qgWmoxadOhmjgZFv2sFRuqm0cbtc
qnkABbJa3ekQVcXC7j+rI1VzBAFe1L9qUI6h3FVLUCYxngSuflnilVB+Npm6Awk8
yE2jrY1y51W+Sxylp/Z8wjLYEcIfpa5ebg0yYtCQvz9q2/0GN5B6uwgmdrFE54Yf
pkkpl5r/d0OzP8izhCOesS0LXjrHQupXu1GSd0rYM/Uoff1jx7jZuyj/jonFLfmd
DsIKydNKCg2zGVswU+cxNNfSmXepTVRUq0dfq+tt1u0taogRIIGg+hhIKaTPIfeS
20iP+UxcNyq23aTX2MFO4tj1GC0QpGhtt8JBT5AStu7RLPbXQKOZd8gHrkLHjmgM
iGga2GZjaPnir6XK3dpYfztlcYZYwO5Fc1mZjOm3OkrgbV2ILMojG/ada7QJ3j7S
0gatoM+lf0cJZxJvyOf+p1QAR6ijYEPmY5eMbPa4bSb2LnXJ8G3nixZ486JjipLt
z7uCVoEfql+OrLMctQ4nE4CCIt+2/F0Zbk+WfNCgORSGL807ofyc9GsUY+VoEzbJ
xzuFcZ38YbC9fm6q8v2cBHgHKtouxAGnjnbifXOUKqRVy4uAL5ElY9DDswzYTFb2
YWCTn0l/YesX8EVn1JWO6+x8aatrUM3Zbt5JpN75rw4bcfGLKGexpsQn9RSo1L+Z
MpT5r1KiOFkMDjkU2yd4G5QahTP9Nzwh1oDm440lpCxrk+LNsrdjmblzRrxq2Br+
17sboU41O1h+QvzsKmnuCBGucRRVfZLO1lTFyHPFsZGbhs2FqWD/jAEmV7DEeddR
+u7pXDCYYjDEkOtdoegTYFhAdiiVttXn60Nu0bT8fjj8HZNoKMnAZJ9NeHNj+rmV
+NYGTROjcrwQE0nSaN6wqbX+bQPoOhDNUtmKgn9rFga9oqRYsjAVe1AzQ0Qt+GTE
yCJ8idyOZm800sclqR0lo2NWVxTR+2mVV3R98/QffpVq/8sWOUd5fP0hEZ20ca3O
z/Vi5dQXF6CPzT5iIry3NVsJFjv9ZHF43x4BljsmoUIOrJkx9/H4DYFB3Pems93I
Abcu3FwUtDX+Ydbtjit9KbJoq1WKIMGzWGNnbI+O9jdFsSxLWAhNaoAFIdHDZuHX
fCF2ln4Nq3BptDh3rW/PnQ9tf+SSJkTC4K7NsZjV62iTG4Vc8OFsxaS27nyWlonc
p4xXiI8h3tGHblnC0ANmc7oNhYanNsk7o1Tac5lTKc6Sq2N9PyMhInZsOEiC6LQs
4yxmXFKCzSR+93tszXtb0M7B+AfWQAb9y+1rnewVG+J41caKxjkhoTphpAWhCFoh
tcA5HkvpmcDVROvfT44Xa1BEALfuE631UyAaQExzTeMmY6rW7CbOnVnxsfL7RZua
YqOfLw9DC1mMWbBL44imS6zwOQJO8R0pFClA7Ph55+Mk+zgBbW6Ika0xFzn7V4YM
sT137O7kDUwr1lrmrGOo69vWuVZNvXi7nxnPk83Ba1AEDSSr7rBXgIF+JHNlaByd
QTeETxZL1AI+nuubK5BvBnMcX0EiARJ/yq4TFhu9CAkC+lloiGct4WmHN1ek2UXR
FAR1CLFv9Pqj0euRJn4AXsQSlt+OXAIBp6jyBVDDY8vIz5nk0YAhVpS25SvTrEyB
MerP0cQ/WiRqVNp1NnfnJmNP/0CYSkSrngS03s9+AQykcgsWEmsrUoMu4v0pQ/2I
TWVRQfCQhS32X9jha4XvVSppuzsckZhvN9kPC2dfrMKybbQU1wQW5hDLV/P+529X
/t55M9l2oC1/hJ0zjf+25ytq6+E4nvSPNV9Kn3VySm7X+BpuJ7ycLORmsggJ0ol3
yn7yjl7FHnKjuiYmFBRzniyylZ7LjniRVHsAK42CrSvzneB4V4H2NcmjqgADzQY+
zZ/l5r3aLNegVO6wxudgUePk1sTEBzJjZYQclNm7yC3wSJYmy1iGMwCZdRbBODxr
MRzNco7sW56O9js1faX5o/Oiv9AkpXgE5a4BY52e8i9usFPPp0NL31z/hLIXaQPi
n1+P2viQs3OcYvB3Z8OxoU3pvKJSeCjs7yG31TlojriHzmQx2PNBX1y93+PVIeWK
VF15eMdF0nxc+AcWRhcoFj/Wj5Ok/m0uS/8+4oo5ULTwDTD87talPib41j1cgukJ
zCCAX2PiSKBgKDVSKCY2i8qq2o10vBDVopOeyn3ChwJQ+CcgCIiN82bncQ3WwKdb
iHsXaduyoOnblijgeHCOcgbu745qULO2U7dJ84wify/f6rJGCv4XX+ltD5AVF7JJ
I2xb8pFaOHRJ9jEtJGm4blBdOwc7e93rmLlFoocCQLVnNaMGudw2cUITEA0WnMJU
jy2tvhkAF2+lRfS8CT4tpLJa0xyngdOLO6NaCCs30mOMoQnKHI0xYgNO3t5Zb6Jl
Lt1FtugX+NDhsHJcuEH4k5A5aZhsSg9FMMDm98gYuG1xmSMiJmSpTEwjpOAbpdjL
ACqpOO4OKmh5E38/V6RZde3QQljaObRNJZFbJ/mXPYGjMigc/BopfPPyQzdZy4r4
tVSn2URc5dWDN3BFUXurH/J/vmJCzRm9Ok9Fz0yZkLuZMDho2xdwbJqZf5OkFvQO
kKYYv6LXu/KJ4XA3k5cxg4uOl5talGUvP1fe9it8KaSXqxAO/ucjfeWcvcgVfcPi
f89O8R8nDYRMVCmFBX1wlVFL+D4H5Oo/6EIVx3Gq05izreyPCQObo/KfTqLaEoxd
YQf7Uw3L7pBBtccCNHNL0Y6OKrPxpwNVd1ogz7Z0xn/v/llN2rWk/ItIXj8xUNmH
AVqREsYnrfAgI/JhHD7WnJ78i0C/miayg8SRl4mtAxUCIaTImPDEVMXGt0aNUEhO
QqP0fDYZUQqmdru24t4Dz9OFBtf6Lt5+rneMO5FeitZXryG1UIh3MknlfvAOAej7
hU+k67kvPRGjebvYDhc2QTTSBXzmnJluOYwh0evjR6fbVnvH5zpkXyKMwdPiVBO6
PC8B1OYsmBYd/ozFdBWIzHeqoo8v9DWo/wgoa9IPXmRvQyVkvNl3NuXmjPT7kZxQ
n4BAu/Lt9OQBovspV6nPzoBO5IfQQQj5qs3HmpPhO0BtRGhLY47M416H7brEqjrs
DxrwtooXMgRusinNnFwJJlIKEAXkNFRUTNegOkmiAD6TmKkaQm1nalDCn4gywFfh
P4OxTapEKWFfk4K25i+D+kld4cFUmgUyl/45CXDHB1twR08yu9NaMcYYZOkxMjoY
XaxYOdbq1DwzjcSy5NWL7nsFMdtxwpqCzIIw9VZ8zR88Jt7wpamfVNWIIeTilokp
nYXuldsMbTFDtWwWPxC19XFC9L1CBh+8ENJ66bDFtqAa/rmYuLJBSHkOwr2yxBTE
8bUb7la4+Z/g8bjUkjroYcl2T5LtuZN5btH4LBPLdc3jFFuHWxnGLoLgMxZJRUZh
S7PitahwHzNsrDf55Lf+geBd8C16rsk2sTZkgfnqrus6ownsS7Xl21sY2Zppb7ZJ
65bE+w7dJejsJyJqig+T89NVRXi7eI8UzfuCkt/gW7VRPX+3BvuskJnJQU1Ferik
TwcvsWyRHFkQg+gRtztN7FImPH8sdAR8V/CGtCqE0wOZmF3EAPSOOfz0WZefLWgk
gmUpPkwUuOw9L9sZR/o9PvcRyYU8aKHaBHs6vpWNk/qAslQDa+H2Q0pBlopqTfgR
QWZWHqnRj9L0AWpqGYFDKFc034d60OKq4Sn6NlOg4J4OS6Ce+qbJ86SvNUpqtqXE
TrLAHrOst5ZP3QaaQ+9nAUQGW/SN2tTnRwyGMqsBKz2ZWH7qYXNVer/64IkZCyr8
oMG3j5Q0GLDcg4BxbZj8VhIEL2/mDTsWy4g7vjEtEOiLN+VfJi4G/czj/EUpQqOl
fPq2D1lYc3ZNi/dumIA5UtFEwuWMkxf0v+HpkdUxoAuxow/3PrHixzIA2bkQjVZM
nrpWEw4reJRi0xIhj4wfzk72CdPjRyLlDasCr75+8BOJ0ezBfREja+5WDrIVCXgl
N04sN78EAlxOqRbnEQzw/Skf0U+dHimpsjdlCaliPcW61DvpxCzR9pDEka77v2+N
2XDwNeU2Q2i70hSulES3wRsDReuLdcgEE7Lq7d8om/njSQjRwwWZoyJb68XIKezx
j7YBhhxZZsq1J9LwTBVck2IzbuO7lg49QwV42cXH0op8VILbDcy6p/S8EZO12Y2r
Yg7cur9gd5HPbzGlYRAAoLvOWrhL0EU5tpDqNs01E2TqRcvsfTF5xT5YnQk4N2a+
MCPyQgeBGCyrj11j1uXXKLpPjkl9g2N3w3f1C9g9Fm1Yb8kO0HLdw6K7OOwqifeT
BwW1vkbxluGGd0ozLhkcwDWJeisVAJzLyn76xDA1EusC1XD07yt0pQLKX4bwKRB2
k4RRfRbLqWc5ZPgDfynqVvZNSlAWqVLngYgA1OFII7X+s+ZV/YNdgAp1bsvxBNa+
T05uWA7PdFo7RkuIxw2ORfu19uyTeaxZS8FCwawK+tFPV/Nd2jwDR9uvEA+GYaeo
Gr5xWYeEoq6I2L215vk0f/pdtBdbD18UycbjoB2Aa7F3gwT6KcVk8xEGfDQDC+pp
6VMdG401Hrnif0RX6tN4tWWIxInCOKuTAQS+vkmC7somrQfwU/BR+N+ysPsgEULm
lER3t3BFnz16tWCkg4XD7fCUanjYKtZDN0jWIRtWcS3DClpaLObT9TAMujV1lAY6
C5KYpOsEARbXBKjrie7Ps52pM+L3ZQtRWo4kwwveL1CS3y6zK36nf08IRz3bafVz
kA7F7aKG1Wl6hDrzQHiQKGorn7FDwoHDQi+n3d+UZnNGUFcBDvLBwg3l9+fm9QF/
ztKV0la15c3xXZ5YdFanj1tFK9bc16seZWbT1tEvaPvazH2v3Dgf2PWzQtRLE7Pj
FuGmacjV+9TpH0pvb4WUXOJEwwZ0DpwCbRe6cIDm/VOvzORhZn1/SFU7qoazzLKr
/nPfAPjvMzzFIIOl+nn4KjQUBsEhCWOVDJk+l02MhG85KbQrtQ4+1kqPgLwpED+4
azA3QHBkFYV8XfZ/WLUlPYPnl/W3X0O0Y9zSc+i9nyYCjCEgwNBTbS2IIb4jHqWy
7GhRAGk1yOphzjF+Euw1TtMLnsNmE/wfHJz1ErvItsSEpMBMX0rsV0GE1ptSjoly
pxKa3Cg2yQqCYBMwx9QIMg8jz3IX9YZwBIoae3Sw7SlAiL0k36Vo5eP1+a7I4DQV
Wgin7P3xFPZgW9eKpU+f6noMj89FdSOwsoCBhjPap6W6XvtfBd7Vko6rFM9SbAfB
OcVqvnDc8mmCprIMsIYAYgY3of6C5Paj0pxQ4uiRFjgXjAk6dQgxba9XsnGEvOIm
DRttLNonwp4eaKv5y20PEsVQy4gO6Wq9flFadu1F9hvPQovUN2l/H91lmjpIuUa2
mPte2vdAWGu7n60gBKLsfm4tnn6Vg4CUzwDW/Rk2Q2kpo0X6xNdj0T42/J+8NRK4
1L7nTI/2Z2qcYNJWX9qxy193zx2vHo4oL9vBoYS/jSsVv1W1VDlS3Au0JJw1ncsJ
ZSFGwlVEETvnnOQwCg0L2p+ddHWjgMQEC3gXr73+nD0S5+eGJb3xTItQoqDXq3MC
fG4Zu9N54GkBgrnOdmum4AtcC4zcfeqJg11V+hsMQ+U=
`protect END_PROTECTED
