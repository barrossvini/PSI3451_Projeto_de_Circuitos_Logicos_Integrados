`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wRGphn+r4lUtMgSmPCITL+qpIel37uioaoymD55yEiKugAf7sFZl4UpZ/vZkqGH/
MG+mK1pqkt3f8bANE23+Vde5WZZ/PXVaTGS0NbBvHTQ7V8w3lEFDuUvzEFZxLmZw
aFkWBBv7IMJxWpxzqy9ZkrwQ4wn7lXEgGLF3ltl65cO/Hzo9obpH2jykFOEgSNnT
RGU/+BFGZ1X+lw4EUQlU2uSI8aDHpFQ0VQskyBg73Kb8tD+XFJ+el+4GGqPSy8Tw
aoIwyK4He6OnRbWi0E6sqoK4qDqjVPuzC2Qc0eTAjwNzvayUS6huwJDJboHZVEUn
bu1sJ8PV6A1Wx9woayhIsuwZeqPZk/ZVADYmmtdvJprQIUwqLB9mXxYD1nR7eTq+
9kpdmt5gvdNLf9sDL31BC7NQJp354qIHH89RajuZ3wqNJah51pGPjPFND0YaNcv7
UeVG7aovmd7vxOD0KkVH+M2KkQOz6C2rn1N5U2XWTQZS1JG1j5Qo+AAsD1b2+L3i
J44Gvjrg67hnwXT9ANjkt9b6w7p2qfDTwdPqeFJKN+CoQVz+bfUhTRdA89VN4n0K
ngTE+L/gOVna2wb4I9HsrW0Q90HiUl1ByWmxDFnGjJdXI+UCmFSWzpwG+zfT6Tyr
c5+dvVFV+2rOUUujmd4ALNnadR30HgkB9VDwZSUvIOaQc0hJOuaSQJjG0EV7WMph
JzOPsiHxm10vM/XHjaC6jlMnDAJrvZHFZ38cFbv2txNdZn0dnzMryatBhZdqZMbH
DK7vbiqwmMlu1JqYGqBBdildS+tXSevv92ssDqnSxu+CePY8YH5JFoW1VT4itrGX
J0wahbcYbn+zxkocCA0Hk2aJUcFWZcO5CuY12g48sVqA5Acy8yy31tn8TR6so0Ia
8+FCI7E974FSkve4ay6/h8bGhCvZcmLaqKs5Ijt5N3FrrUnVQBjxoCM5KChhle2j
FXUSIsHFAKI2NsBK+FE2SNQ6ik6HekCOyP8oQ4FUKl8o495AQWmLf/wIXiA5Zrzk
HlMctfY1/41NQrdnkoAF2wQKG6u09vU5CLGvT5DCu0IcKC4TomxMpV9GjHYtuoQ/
vNbG8tki2KstIyD7gL4/i6lALovhGzPXmgLXNEEeExlrKhs0uTzWwYtc1J/L2ZU9
hrCAhtOo1J08Pj3ofHWNtMDATfwq1tVaiQmYfhM6a0qrjfMaUAwEDMYyoPvr31Mm
`protect END_PROTECTED
