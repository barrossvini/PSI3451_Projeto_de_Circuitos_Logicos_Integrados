`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fmopd3YWPjeeZXQQgIRtILUm7Vv2P0emF1RkLfJ9LcAoQ35qlo8RUABeqhPnJxwx
Xwgl5VD6sEXkUri9+SiWPNJb0qen/n7ZPHAkE2L8OPd2s2eUWqkoyB/ap3xrS7ss
yL56NzWces52QZnCIzN+0N4AwrstqQ8b6D/ZfZiXPBgzSomLxnDFvW0x1lVXStVR
ns1LetUfmdJRx4PJN+83XAFl3BJkTl/w3mEq4lCiSXaEOh7sxHAUfjgnFXI9eLvE
gjGwQ9bugKLSp9bmTlCNk9KZeKecWEBQrnC79XNYiWupbEvzNvaaHjlzLaA/WOk4
ZL1g6qjWfMZTe+J9fw360hFUZX5++X9nq5tqdCK1oFBk1egHRZkx/KQsC/q+59DM
u5boHshcvpSCqifCyc5aPaJ45p0ZcKxqu4dkFSqTztWM9bnRMcgY8YCAH/KAFc9g
1wH7hX74wHrhWvBxswAKjdbssevYSQCPivkedc0cNSOSR0rNNXXSRk5o8o+S5O52
NUmnPNsBm7q9oe6qA2plzgGD9CcyN3rEaZh1bCU8q9bnHNOPutdcxj6+McDzdV0m
ouBVpotZaaHbnubMcnsf9dAxrWW2iG68AvC3tKd3nRB02gn/Rpu5dk6hw3qWUIws
8ceI7H0sArSRuNqzwdMfZnRfUKZPqNyG5bcgB5TDwsQvt6LEqTLvzc6/jwGmIDhW
ObJmxIoHXJLF5crFIf0vvDNAM7pDB55DQGhCWHbRqxtVj3VFwrNw0FjZ592goN1p
NLdoHiowSDZnkbvPRrm2QhRSZItgTFkkt2JnHgvxE4n2oW9baAoh0j7jt6UEoQTO
LaVyNK4KNm70jDSDWi0FHQ4kSGNsVLM44PNXrlAU0J3QVPAun0X89pDfy3ITmMot
6b9K2J9EKja+fofNmbhw4mOPuw360tKuOdQkeG+spyZemfjytoWhIV6do8qR86Ee
ouejl8tJx0sQDGfhwYHvpCRKaGuTdQHdySw9jQa2M8RYE9EpKK6NOaITHqnzuEzL
VGwSH6XW35RIN+D2TpH309UzopJMFtaNvLejagUXAumsHg21t+Mx9DN21CDqkuhp
n+bpSYAlvM/J1Ja8RzrZxrHxEpB6nNxGuUW4LNopHMJ9UQCfzfUadaV5uv2qfmdL
2f00HVJPYgsWYJyh5wExZMnJkd6ASCfHJpoJXLqckplCZdcPmV83DFlNRvsptZuG
ZCr5/OwC+w0OW1stjvKdt75qVNq7frbz8O8zc9Xi2YDCqRkzhbCmOjwvdaH+73+a
+1SLC21e9YKMuH1PAylH9pPq53u1kGt05dfiJkjP3rdyFoYB0AtxjsYo326YOZHG
R1ESH3rx1hvUK3woxOqlWUvWGS5C60BRBvZu/gRz9YZpJCe6s5TcB92XbbZDzojp
NAO8sd0rSZKqEeah0yIooudyzyAsJtf42E5s8r8HWEb9nmZbHuF27rmzi38lhTQ1
Z6MPaur3fJdl9/fvDsT901+oBiId6KJFD4hsOIulCCIfDx7tOJqRrEwwj0sO/jq/
AGVB8PUlTMcNKOzOjOIYDrffsYeJmQzdL3ZCqSUZbvrwheXTibjWhaGW95J3roBO
h1uLrB2UWfA0l9CZjfC0REqJzGq3xyU67isMkk749MvwW/zvECIX5h73takfewME
ycF/Ywk+y4ntt9O4LfmwhSlMwHRSxq9joaJe4mz7EhOTF1wJ4rg6fRxEpFUyHiPj
Ybx6uqZyBIbUtzhG6Vq2jthlb+iiudhpQ9HGHYmmaqNBs4RHS0f5x9G8nSIKP8gc
lQCW489FrPg1Ppb2qgOQY6mI/pNN3giiRGZiVZG42HcAE5tlWtk5lQEq72HjA3gc
fzmbDbRZbkwnIi+7iRRI/0woXVuJmqn3ybpTzhPfWUOv15JqC9Y+nMVGxerlbp9d
P9vzswiJvRXcZGsQVET9hzgBcJTYh9LPHDIjdViXV1X3djAK4P+DkJWoglXtuSNM
D00QkdhG1O0z0ZzRcbHZHonMnJaMMSpad+QpnePI3klF23F/T+sHS1Wur5o7MqYZ
bOvctIasMvd1Cd2RH4jULx1w1+QeT3M1cECb2MPbvvidm1AoOq3qRy0POnaPAajY
SkQO1M8qCmVw9MIai8vChEZCifgB/kspnW1IqquyJV45EHvIJCuIaTUwzY4R6qpl
xZy/P4HyGSUc7dDRIgNbhUPxmejpfTlqKHKEfyZxkSoTsoomRQy0oh2UEPRzh9Et
JnEt0ytoNiWW9gPnJRTPdvAwb4iD8w9ODf0KjfqN2Osn9FWl6poewkD13JvoO8zq
wdJHoiO2lB3kQSBichvTTAMRVXMMRt+6KUXk/a0z+XnT/yWCJkrUqZXbNIYFHzy6
0yz6D6HhcRf71HHsuAvYIOxDXr0zPs8bea/ZnRHlQqHlVdQA7jo+ddSsC+kKYUke
iGv79Jy83DW/pEC3x/7w1J0vGdADLSQjS4+Q2gwML+y3DCE2pNmwX1mXxFsIi5sE
s37rOsIJKCc9I4h14JFozp9smGOOYMhzO1qG40OfzaDJABRTw4T1LzM15o0LVpyq
XusAh1N2y/YY2jT2/C+l8Sotd7utGPWzi+POW3wwidj9DPl4xDuqVlJP5ykvxOla
71+RJw9NVAgTOLQMLeV+wv5D9Vp5cNxeunQQkN8VWHHB8dOkjTXdMYh/EaUsiKGh
SS5eMIzBhAbOFoNhYj+MheABM3mThFWzgIIJfteE0ljABHG2smuaeWESUcMHb3WT
hf+QkYRtryj2df2Ec7H0cm1GuepWKd/c9xERO+c3OlQMzdi/caNuEERv4hj2UHQM
NOYs/wJpP805Zz1aTFD5d0REYr17BHINYRS/5QF+JuxvgvGIsLdHlMh3nJFi0gV0
+QWl4G+1WWaI026kh2Lu+BevoFNrtSMrEcfS3XasTnxaFKA9iCWitsUlu3TV+iAZ
qKBitSv5/H2SVt5GVFWbr0lhIcIWQIQ8dG6D3gaBrwBCp5ZVPM0zXIt65Y68Ky2O
WVPIuXSg+S21uYBCS906sqp3bZcoSXLLpTxRSe06MMZTQe2Z5QiKT/kEH+lms311
QXrH6rdDmKScL+efA04jSALTbUdiAJwPdC8Aubv6ME54UiTIqXGJCSPwneEI8Wss
83hJYE2xzVJe5qH4VkjpfLT2PUTjlU7jNLSbDezFhhOvhLFo2de6rs4DzNNJgkfk
JhVCE+QVQBH5pc4h/b1Yl62wyPIZt+EBsnqa/iaRo8UCB2clQ4wE0dB4AUsz+Kge
Z5VIlnRtTtNr5nElFo8kNd4MhWEzKyq1/AnRuWzlRLjj8qehSUxQI4DUiFhlUGpr
NCWQrzupAFhmsfGrC4ni0sATqseG0+vQPXXNm1Vki6YNJgxbx4KxtWEaxuwINb5m
8nPitromQ0dhgy0CYKz8pBe4KPRFblEZCjhkcQK/xWe/4f1eLQe5BHAWRhfzGGXq
+iW0BYrL5OmnezTXL9tsnO9woE54AVsw6u7pk16DYbplPngigoM2fkCbZoYDBQr8
jqXAezCfH0cVUqZXG8KiyYtA8E4ORYurJT5GF75TYgXlSzIRbYfA6QyCWl3Fuk9l
XmjnPbm36apm+DQ/3s+XVTuXrMyPdr9UYXTNyFd8k5CnQri6D7IYJ+VOfqcYyL55
BJIunN/1nna4kOI84gxOollJsHzGV+OZ3YEttfHGHanAEz5FnPB5QKRJSppDE2aH
IE6rRptKwQgMe0xtJt82YdbR6fH1JSphQVtjVK8mWJSERI+/4sLUtdZ/YClVc3pV
U/iBA8VkUBww4/HnTBWDPOmLR/kf5Ist9uqBPUdEL2f2yjNC/E8HAN3VclD+JGtg
MZakddXXfex7NmzUg6slhoOiPkJBdubOOBmkQnjqhUYAJNWdMJ6nD/k8oVLWSlvX
l4AxO7VkEbxM5OH6XfehyPk6I41il05xKGB2SlO7+stkVLoUp9dRCKt/Q3cWnzdu
Uj6El+oR1b/RnuirGnUhYDN3yD983FB4Ecw2zp8gSQrT1iqkNzRK/I6nNP6qZDwo
DDdR6+ZixPd5fFa+HEr+Pidl30evZBK+W1Sn9LA1l0AiHZBfiAN2RQtPigC7RRI4
oOTW8sCU7uv1F/Lgm/sN/sivDx377teuzwLCVLes3VFrX5WRbtKRt2UUeLq3m1kV
jpfKRBbCim+YHT2OTR4Ys7iHu2x4GVsdVtY+EyMIn+5Io7wNvP6jkgNqZI65BmBM
+Hkrjbx5sqbudje4pYjmVyXR81y1RXHv6tZfoeGvlTq+vh65ChZavWsFUZcZRk8q
1c4Ocwv49Is1MhbTXEzK5bWtJBskZYSOzYADYxQK7PS0hc5Vnk9tCxFXKoRQ6q6i
qbnJUcM2PuIf9jwiHCEhZk12mHl8s1tfqRhyHrTJy9+LoTO9a5Rj2qNEK7l6iAWK
287oU+fCUXb+s5zNfILOtYFsdeomKrRlV2zuEshjVBB328L0Dxhuhedp2tVQf6JT
KSb+lbny/WYL9w/V1m0VkZ0DYEqQHiUgJEHfGFomrpfiJYv4LfullrttbjCClxoP
msb1pn07ztJbEhslKjvV9HBQJW8yuUWXevqwXmzJjfgKhvh0x6wa9JdjqByCeuX3
wCKGusFXjKeexDJywqnaULtwW+04415dyT4X1Zywu3sm8KE9xmicUHevhRD5tcoO
gr/EFuzXzMWKufueHPxyLBNHQbpyWs8K5y2Yb8TLjB3C7KhZ7GLfTYt4Kcbs+jzG
bZUNikV0DeYIaEc1ijnQOdPCyojgd+3xVxzk3x4kskyljaaJ8opXuTvm1sKhyFX+
fboE2wNU9YEY/UGnWwKHodkPHFQ8QwPN2h9E0s1k/ypZFNGD2ZcMSp1ahObDGrUT
VWeBjoP0mJJggY1tePhlxNiiO+JaO5bhSflTNfJ+WVBMspqGuIFJV8I7/jAeCKXZ
9tGphLVpEqMl95X3W1+GdExDQOpiXD9Oy0AnB3tzOYZLXHyFh2VuEnTAzemEXbf7
gbHpr7Qo+sad4hLkKNoQUSRwyloICFswBNcuo2laItgAkn3alTLDzDE+HEPwLoGk
OGwYJzrrKIWO5TitPcTw4RtboH8W0myOYLmjFX2mNyf3ROdGuLCqfkIsU1INTgO9
ee2Z/WlbBBbd1lzeLXoQ0lSGw4FBHGnP5BoMBBdJ2giWXgFgMRm4sA25U0IZVxrr
Rk4h/IMQSMwdzt481S1Y8uvdKUSO4gY+b+mom+a0JU5gjRO4qgAwXdEXe4/d6pej
osiuRPshtFXDeHqSap2FbrvilfLyHRWHW4Di3S9/zIHVcWIwfR0YNCJgnCrrYfOU
pzqxrCF1C2wirKuJYOKtv2RGWYuoi+oShgezyf9L2Harr0PKofp8S2AnCLbrR6/4
3V1upQMQWz/2tDSAM+OVoPjIaRz9CL+sfDYGMRvN8aMN9TeABrerNQ/pM/BkJe97
VKZJz/FmarKYOS7o+gDEiThLVG8MePAqgq3+3XURZndOviLfhv+qeJ7b904IL6kp
LaXnhLCVW9qSY+Ch57uaZ2T84fRHM348dVEBWvYqdMX4p9a69JA2dMVeJLpUHJ0a
K6AYhXhsjtH0TKFjZkHbz2kwLIrHcaW+Bee8uPGcoWxomXYk29222L1/69CT75vb
BxCbJvv8KTfPRreGuhMJf4dMeyhEE8lKMDkGBwjcz42zHh/nl9yHpQp4dSZXkqYI
rVIx5zMVXHWfH27tycrkRyJ+KmMvPgiEQiOt5TbXOYmUV9TirwutIE3w0g3/XAVp
UPjjCD7fklyGCh9qqYHQ2Cco0rezsy/EM7pmpBcK27qNAieZUio5TJDJZxI16fnH
9EoQJBv+mbUK1ZLGx4ih4F76XKI1SfkCvTe/d2202tS/SqnAzpCiIm/di0o2Di6Z
mlsSgOuKfOrEnr+5IkIoUHe1y/HCXMi4JRd6JKfofsg2WpKtlYZolxRlzIIG8nxc
gts3Dg966Xl+QBghsu37JBOdPq8iGlMX1Av9oA/uZZIAiYF+8oG1Ocpk0uEiPqtL
hYy+t5JqSFTjM4BqnTvjktrwY6xpFirJCegdIgQsJZo62dtrpjskJRKKlP3A0a+q
IVQtKoJaHKp2XP9QiLzpD0IsFrdmt3QCLDe+vjMDrCGZdQbkuxPnDRcJ3icnOcAa
vcwBDkwFo9cjymBhYkdkKuIcEcTuvRSZEsNMd5cmXcZ54RhZIYz7weTNudFp9jLi
tACQzB/3+Evw1FlIcgqRNaBKfe6UeX90p2Lf4Dqs74Uh+Z1DgE7LBGj2w1r94WNa
j3IETVigrXVoQ0aHfmbEeC+qv2YTUxn08tRrgQ4mEHfpro6e1xQ+rcUT8Ux97/Wt
9Cy89NcYE1/dG/QcDxUQtJmSEG+XWOO9tgqPyeW+z7ucWtu0Kvglt+0oZ1cQ2LVG
K6S/Rlh+n99GbKAdNWeOPqOfdeTNF1XOefgF5lQ7tUQ3Ci6dBjx42zn5Zj0jMOyV
+gBGK4FG0Adcn0RHxhNYNP6sLga6WgYekVgcsP+64bi/8w25rgeewm/AMyCajRGk
kQM8jx96ufouZYz6MwGKwvYQeRjNY97Ih6b5OGCcoA3Z5DMplmFd60RvqmGKe+3j
KL3DZXjJ3UtVdDWXdDRh0fDli66WC/dtFRzi7ODMF2DN9t0MZCvPYtNswtQykldi
o1WjBS6B4qECUsSf10+wxqXTiXJ61+aYvMxnFh2nIVfL8J+igI4ZtchLNtgIxHQf
tH5zUSP7wmqJqxYHeDASOHBUjowMd0ioJgPw/D1Hm6yaRvUWJhb9IrfGfSwo3Fx3
cBTv4C0PnQQH+9S2fs13SSPz8dZtKFe7LTCHivEp/S6q8Q+iHKjJZ+roKAvpTbFD
iJ4u8EiGZWz7ej/a/21/wclTmgm0BSxLAwR2nf0KJAdTRl7yCFbAsI3pZ5IkqbJq
TsF1iYvQdvQiyjeMeU7gsK/o/3oI2WiKdoGyNjHmiP8bIzTTrlRls5YpUDPGfZrU
Dr2HqzNWV4dQa8o/liduVVpxmoviLCu1qGwaAncIQ+1C0w4Qr5jtLLWTn09SVjPo
W0/tZuDyGq3FJTBYRcEiCeszWUfJHHLw/Zwae5SGc8t8RN/bU/laMaJuA/PQID1Z
zoFxseab2QWyMMYhYmmtM0xnx9VwnCRSYoZ3HmjkvZTyqz5a+2sdt3YORHmApcTy
wHc0mEIoUYNFGXhum8WIt5N4JIsue5EDaz6C3BkpJJrWHUYfuJ13VWxdRkv+kMEl
RvHb8P2kt0AnKTXwI0sJjDGitPjCSKXo3n8rmVIl1QguKYbWmx0FWay41RiIu8f+
vNGLpNOIa2lpEdGwmCVS2urHohTjtgqcHL2f4Dy4QBR8xWC7xxybAwU6gh6UCerw
tsbEa+Onip/RHgYblwlW6V0f+1nQE84QPZ6vsXtEGc1jPajsGm/vYcq3sITM7rRY
jBwU9V2AIGER4wkmunWbs69stFcxw9kYQMm4EUXf6J6p8ZNVIyOxIAHBHnT1ZI7+
xFrI1QMkjAevPPPIVASnzXF+4hp6XohMw1v69njH9Ema0j8daotZGaKgOUCbWfp5
S3YqTJx8LqG5SDUOAd8x9uvMsgEeLgphizxtLo+lzceXqET4F0XVyGe2JdbmhAw3
TxkWy/68nBZYaItsD+GJqDxBtdifW45JEkCbts5CDCO4IsHOj8gdYpcBBA15B0S3
aA1Ryq+qI+MRZdcT6ly50X6LneSnXNhw0A9RWPwQmhx3G3EHL/9ZFqRqbjRQzKkQ
cR/C9zgvpNjMPx7Jn6LWmo+gcV/yAdYwscPlZqmiIYI39Z0ul36WhECIzEaLHm7U
LDClXtYhjIfAbHfSvI9ct+FNQSWn5f/bQE+SFT5npFcjjydEJCCl+ud/lyH8+okh
fuTOQQiwAxGBTOgq0NT0SAjO7PaCPFV7O3I4+scathZdGHtpYKPM7pSdz7x3JzTV
EwcJjWJzTmV3Ec6ycgBZG0K5idKa+8X6Ds4NWDXo5dXyS5CKD1PqSb4fhYmwlalM
K4zGrE4tgLImfiPb6XGiCXDGy0tCaP9gGnLTvnM+UjnbMO3+0uoB62Txwu1kp9mD
uwr1PQ4z5fdpmNBPF5il40lSKgEZGG0w8GC7xWOwa23AY+GEfIG4i3/LtlJILknP
6nHfzn8E0nNXQS/GTL//epOsTZxdSvMjo7PCYWNvzVZK6lS1q6OuDJNfQsBiujR6
g1rjcmYAVHjQmbsg+jymurAtqKNYRqvUKbM/IblfdWgqcqTtJ1NwtKGfofIrg2DE
t3/ODQJRH50YTI1RJFw7hTxENAi6b7fLHJfhuIHutkJltVaHyh93Bfo9eCT4Q3TT
v9ros5jzT/yKh4kBwguIO1mohkiti07pj3RiALwOp8kL+JZg9yI6sz8u+WIG5PXa
b2Yn7i94Xn7/vqN11m2vmDU50U0f6GlemLrrO1uy8tlBhQvLio+61zOuknqCadee
vFnnNjZKcTvW7V63FayKnuvIJ+LRVo8CyYjiauTIMMJ/FH7/wtijhHujgxDcI4To
7rrw1NB1/Ia2fX6Ep3jB/F4+29/qcqswi+C6aaDoB5D5KZIkCWPrhBeh6Rf2xScp
y9u1LHWFFE3ylz4vMm6eckVn25VwQOB2f/BVzF1aUgoorqmZWALzs+0gPZXc8+iO
u/e2azLP+sq4sJfDgOUWGwaU3dr/LFWxpf1QHhddXbVx+14rByUaSr46FMcTSdp/
LFr16iuo1jToXfzqEt4kpVQ9cablo0l78M/EiAxM6C9QmPzblTCKoRHRURPzGmzE
gu7g+XZpTvXjHeO1bZl6gfgX4vKDEpNp3n1msczBwnURSSPoBquvJaw9isGL6GzZ
xczwfooAJTUSbFdZsB+SVP4PMzpzp6n5c5Hs2b1hP6SmCYsXSFIWxnbJ7aODkptG
9eV78FZXDLt64DrnFgUVmpH1WyTifJVzM2EckqkMX1H0ofIDx+NEsfuio4fX1RSC
ZDq+hFHJ0iw1N+XhqhCXQ2QG7bjbwmFU8Kg1rlCBn6zHdp87xdLOhOe9h2nT3ErE
3M5yFvazK4wjXzyxMQGyZze2814+RX4PNN4TtwUM2TvtLsdPxj0PJz2yJTq+FbJT
DpLMkkSoKV5iohNpQ7zP4CCC+VULRb7VqIwcRlp0OlBuu93LHDoGQWe7Vzm4A41A
L+kOsieaHq3e6JmtfmJz7LSv/Z3ORJKdwGMdDtBWB27z+txQVYRXt2Susu4Boc10
relqbQwQvDPMGdEilwB3+XFQUi3utR8w4kBQYmij06lt3RS6BLa0e9RhmeaKsgvy
hqGtQ5S0AYhfCi2T5vxWrqZuDOqrykYSnjEqIVoOutR2iFiZn0/d88roRluxW3o7
XXGI0dKSDKVyK9kbs6sK2lEl7QG45/RWu8gCa7v51O3ZSmpOeVtPxJRg0Nwg/mf5
xcSGLV0aPK6ryB7QPgLITs55rTg27VnoHZv4ryG0UiiCIZ62w10jBgouWtInNltE
C7o1Q8+DIWJu7UDKkvBmeUZgLLZztKdZaFveVgHY8ZOnYj3gxABFbO/EqLGOAUh+
mXIRYLqrVsuL15U6Xd7IbzeNeDFKZ8GpJfIeayQ3aWOSMyQFDV6EWKGSYgJs6+MM
vjPuFp1osVvJP1Dj+eMHuFAhUBfy6khbedTkaUjnThkplwapf5A5VU8z3/UGEUsp
JkrNu2YtlUBszW7djy0Nf4bGQA4zwq1D4J+jxyb7GF3EaScSr8aGJRe5XU5yy9I7
NcXamhgk9Uc/ZrvLkOWAzVlSpoL5bgWkyFjWcdeqXAPUF6qaAdQO4VjoUbeo8fVb
e0rLbT23NSpGQDNfFe1FIztcW7QDV5fjXVB+jnfq8PRmfHkKwHEAynIRYNFsXmg6
GNvOCYQav8lpuM8UV31Bect7nYHsF/lpSDMx4kPtqj518+MNt+WJZbPkFk5SdLJp
BbHUGUNyyig/DM8CrAlsA+xKZV465mCFjTnbJMIzDOI32IjLzBLDPg6uX2YTQQDZ
eJtO0CEeDh5Vd/ditG8vgTUUNrZa0S5PW/b76KM9mEv4Vhx59GhpSp9Gxbzmv56x
ykCzyR92iOo4kRH0m4X03kLTM13dPZiv+EVOBs7SnGltcwmZpG1KfMY7v8qt8gW1
rcqC3zhKusP6HS57Xv0c8lx65qdareDmyUdjg6ChRmxOfjtvHQZGO/YBgdDI4zBf
8S/BJiwQaW04cQRViW1ZzjW9IuEKOUnCNoP5V7d1veJI8wIFg+0yqGzuxsJwb/8s
B4/LQT+ahXHmGdds5UUfIO7yHdgx6wMEvfZN+nUO454gd63X5QsVzW1TxxsxbEJ7
DyMyZgEAgFjx0ZD2dqJRm0NTNo1TdGJ7Sl632P9J/tWv9LR7Aa2nJ8elxZFUQKwT
vXQ7kpL6y0vYFt5AvrI3x1nehsaHKApcDzrJNhkdGZGy/RqltQiK+mHC26MAFsuK
ZGw6/+KK1fMpfzkX5A2OSXmkyO5BPKu3LCcdjuNqOdoXebUVT8OwfOqEr6Nwo8Z+
xWW5EjmdcdQIABfbzQU5E4c2M0bjutV6bqwbxn5nIjb8FneJU48qUWmWekSBwx8Q
A1zwJgfK/Bzc5nILbJ57jIyAzk/CHRGDk+QkjssZiDL2wGCvXptsWQlDOusMGaAM
qJsgkq+Gh3xIqWi2zmF+zS02mh9eZpJF/mj736nfBN2cq/oZPG1O4YpFbxMcXXla
ZkSltGIhTuXdOJsELJWsmtdQ8AvrMO4/2QDctGfAnkzPv74uscwCSI3eufcBiaF4
fHQGYKtJ336ljcaZJXxgY0lrCijlPR1zpFSQJntUhrPc421m16luu+UtJow0FlCr
8m66TE9S83xvTWvkwARbBjCrNnsKSp1b//hYEVi8mnUPF88SiYUxm1+9roZZmUlD
mQKZ94IhuZVlUnR3gszqkEXZXmBLbZDE/X3612LMvn78vO32bU0VdIADw8dPwNR4
hshyVSYOYXQujRJmJ3DL6w1Xy+i3emO7dZ7gvH50D7F+uZkCvx3uamImd+ilz6DG
pyCGvn4oRKBege1EHHGs37ifuy2epUHiBJMJTOYSOxFxYdnrURMFVpYUeo+d4p9I
DxmgN2v6myvT+AcqB2CTlYJ7YgBIjo/uxuYZcTtCHUfcm8ZId/fV/9dBiqYLjABT
5mKOs0jvzMXZGDUoKsiUu4DgbhBvS+f4/RVcAoYtqBgYUUoYqc1QsaakmK46a8W0
OtJmmxXsH7ncZZnbqDyDoRvaKrKTrgVWJghHe153LgWbMY/D0wVmuv/gN42kd6zS
ZKg2wyDY8UOLBOf7vY0etYVEN9UWpRdzMfJtZOCN061HRcEQ6rZ1jyu0xiUw+Pc6
dbtrB6RyYkqgOt3IPNT8RVffiJudr76QNixg0LvdXdzJX7sTVerE0tA9VlDNRSLp
9l+IubLUi4DXRz/FWIqBe9YtA5c/0vRb9BwpA2VR2sfBIfSbxbhJV1j2VjtMOjVx
OkbValbkzwEEH6yT03564CpHSwLXnmfRO9N2WDkGzICYI/HYnXXKvQZUVnTiyH1s
qjiDGci7pKGXoycG0iUEHzyl8tk4qOeT+L5cwgdQgURV/nM6gdrdWuWGc4n8vDgS
o7dRXAss2fcXQamX79qbj3qNvuQ8VPVyH12jxG4n/XKr0xaztKbbs/WHRaolqFLk
DzPZHyZ69tM8kRJz8Spj+uUd6m85iyxI8lyzK/ImVmnHMEkuzfKogOH4hmQk8aT6
EjuzL2F/83HiW/YVX9MIf65oCcykuoWPPMaCJK14tv7YntzTnOyBnnfVtgoo5AJS
FFF2vfOmOnrErxvR+I9oJKb4QWP2GhLLUoemE9Sxxu+Iz8XbOqgORbTB9URSDb//
TCCdsP00fIpoHFCpXND+wJIkDehUsAU9bol31ZKUy0F9Dwf8UbINUIl3O3zaBbns
loMAWfLRg8b3KXn2BSWncjNlqzd5P7/tkq+zW70XcSDVeqt/q9e+Qbztxh8qrWzK
TgL2DYWjcfIJcO7acl+/VlIrbnWMAmOHq+3mPZTm98sQ25Ndl8wkcAUGJ9R6/9i/
DM5ZjR4LPSK09XtNgSeiwtbQ3FABiuMQwwCFEn+8ebn92pIikB4idTFW31TmGhtN
TEPY/QNXRKufDBxIMgPZcro/bo/zCNzX5DLDD3yxmVOfPHz4cI5WwJNuXIFgMYWw
WECalMi65DrWs9ZFsgmCeUL/MiciVC+P3fHYyYx6TvQZl1KYKJ43tORSkWzweTWc
OydZvc/JU3G9lodvviRfe2l7O4u9vfV10OndhTIscZ+0DVs2nS6JQS8jbymx/fVq
gmf1D8NSv+deDCy8E0p/6vTMQfGM+ntWnTYmg9kH+7cY0/EAs0yoK1riHV37RoWq
5gOGptcHQqAFv5ygwOtGcXVZUaoRmc2RxtNdWwh7QHRtUR40mFFoklUtFVHn6VG0
zsjMlpqzvULQKmEN8cDXIi5btzytxWYT2Wpny5WqC/JMMwVgBxj/xNH45VG5lomQ
HbhfaosmPew/Ltl59Z02sLj+LftzrViubqH3GSHKtdiOLx3qRvdUrruoOPnymDKl
mk8PEGKtCdXR2MnZkmosBa6zvifkOqdG0TKn+6p4vypahHzAKdzsnPdW/pfOMopZ
ti3BekBcVqryFn9hwPoo+od5A3utmpt56zFEMEVNY72hcGcc0lyAr/I1Urzfe5z0
syrIEImdm4xK4tHOryb9s07hflFSOEUCi8ci3z22X359kjNPAHQ/DLcsdvowH+lw
qHiAMi5Xj8RhBzNN28kVZOrHTHWI0rea6FO9vdJiMCzeWUnGYEuSCqvtgX1B9cyL
GftrVFtw5jA4wGbEzKU9JNz2Xlwi7vzMkG/NcP17c0OBIBaH5MY3EsKxejJqG5ci
2SvtlJF9kQ2L8iO4AlPcdoqbomjqeKepHjqpps1P913agAryhADH1v+fkJD2qK2f
GHDMrc0e3TApxPKMekUHMJi1Sw9rnV5qTJUv0RwJ0qVZ53SghVGU5qIJ77U3hwiW
9o8nF+uBOlVoNPMTJmBfGWlhxyOgtbDo+yOdypbIF2cQ2Qdp2jzj4f/1to/elnb1
QBF4Qu6uS9jWMsjg13fKNeISa+SsnVmNNiSeCsj9eUbKCRmacroPv44Xj2hwrR/P
5roY+1OgPXx1sZGOCyGFbDno+Tyd+v4+WiMKHWzAQBiQIzSE/qAxu2uB8/F4r9K0
/kYWtF1HJ8d3s7/m7ytqhoQ4fFyU1VVxJRRPN+xpKOTfy3T8T5z2vfunmvBOW17h
/Vh4UBOP/w9ImPfBHFDzgI8Q7AMA+AGqzyQMBIpvJhBcegcpHQ018GW/+Id7tdA0
zT0pVhm5gV6ujYZ0VLWThVEwrCFJUxeRXWotpFkFWe2Zsm+gG2sfME4Pu2CSoGxf
0OLZQfR5uS93ok61w9GHUKQEDQoCkejaNeA7GSTcoTWZgJa5Gd/yJSiwcshQA4SH
t5SO8uo28cWpUP2zkG/auW6YrUKIoM0ZjRV6fGbyFw2eubWmL5URywGdP8+z5QVG
hDx5XVG9FA/5QH/9k77kWURkAH/kT0MppvwYTlFaAtnnQ/gMyDLikhbrzQZJGkEr
owRyEVAfPwV9NvQgzQzqTEB7gQ4CA9N5Jz6CKnQWMOx2rEHsQYq1fkQiz8ZbwCUD
oryQQTKG6s9yj/bWNRHKRFzpL+qg07dQElNL9DGFv+5uE+7GCHL6/3RSYkV13eNY
Q+ENNQQnFNuhBDTYh3eijSTpH8E+btfndLnLKqWys/BpizL9u6+YBK0KqbhCqfF/
1tYHh96hVR29hEkKlPLdZU3BExRcaOF/zghuyHupnRlYiRl7YBkshN0eptfaL5fI
BH8BtqUzAN8n48F94+4RxntryhyrT04oodFgZ2vKATxA/ifc6cs2NDrrBpcOeu6P
kh8N8ov4jGm3HXNkqsg2A1sK7Xfi1lQodL/ptgBncoFL7HEagc3VqH0NbNujIgJ5
Azui31tvgghdSFmPDaT+U2Aby7OBihFU3usKQncTYwBWd1METCT62JPGcJSI04TK
eMM/9g8Z1jIslS1rff90trRtwoe8riyo/wy0Zb2arPQwk70snGLPSr3YLyZqc/ra
knSGnQQuDALBSe8mQGLLs1+SZSFFUyBH1h0WTP2tH7eQSwVPfv3GzGRB3EYMBcSi
80W4SNeGc2UC1ujslPSez7ldtdxxroJiCfAvd9Me4apj0F0qk6eB78rb+aDnWvUr
KNxkJ+QmXSlOWRsFgl8X7UBlJXQTwDyOPMB/7l8vxHqzLb5HDRPH/raBlVobAyYO
Gkngt6+tOP+ZHkNIGCiR+XjZUDCVkp505/ZVNxtNhpLEbYlhowQekNoiTrsZ+1Ff
wwRVawJq5a81A4qXXyHPrVhvnmUdMy9vkBIObaxgCKEG9BdN5/jwLNXZWnUKrIOi
8Eu39CoT3YaooTyUZvjR87R0jmPOuxEbE2sqXz1FCGjZS6Fa/a+ETfUBX5O+Xon6
+iOJZPciTx0fXwhVyJWZHgdl1f2dY/YvDDNC58cU1LY62l79nTm8fFpk19TCL9wC
wHRw3GkPIta7pPEpH3KP3u7yKKKtlTLoxosyKT7liYgBYB3pnbxRrBbk9l3QROEk
cBOhuFyg/yNdmvMzrBjXmQJL0u7oR+C4ej+1ZyX2ZczcYHpwlrM3ljbGYPn5BSVb
66o0oMj8h0AgkjFw6aPNeroCDqzE8RdtPyU/zdRF8RKJXEzgfumP3n6iAjRCfqdi
W3Snh41bQr9lTediDpauLveCOs/JUKFy1Zkjr9B08ySVBi9Yq/bVt9aLUMtNgDTi
XhjRULZhkDgGpNMzNTc9rpVVz9Rza9bLxKRveHg1nKJpuuuowB9AjqK8nF4DoY7f
30BpdHw6iAWhLhkeiDXWGfM/ckIL4tuWJAS6uQXaUxRMGLflOjY3gILbL/EXhyYP
FcaSOKG1UOkTYvMpn43ovPACe4G0XWqVdiJt8Y0ENK/zgEODfqBuI9OcYzYGWkyu
ID2WGTZ++YpqTwBn0c1QPKS1R09zTb+5TGPPHGyrzlBvoml6wfPFbKf4/GAlwxas
bTD7EiOnlmXSGzAu6Kfl3DvSOiTm+vKNG9HM6S07A8WOw+OlpgfsEXYdDgMUsx6P
G8r9yy+3By+yRjcs7NBRA5fiPu7OXWgAmk/fz9azLtAqMX/WtNMbb6vpA5RWF2il
82FYdadtzsU4VZCTFIKJWwn0gfu3JIl9fCqQ/kdRQKBoXWqqf3uLJbadFYkheH/3
jPD5KxhBIVfkIa/Vzu5GA9bmSPoq892Zp96hsTZ39BC+ZbQouoCUUjImS5XYpIZg
Bkc1s7H9BAzOctqjRFoCA0X8R/axXvmikXseW9U3kSM+yKiBkGPCUHUcC3N2nuJz
be37eTfiU3DIDdJJITnqijdFllgsEyEA6kriHVUAEYK/rqa4ZyrhAnTUQVvY2kJy
yDQ1UeNvlRF3JEkQfbXiP4fr9ckNzaH4+8Wz4e6d/r8RjRR7bvL2YKw8c7832/5n
lnGGnC6AOo/pLC5jXNUdF49GMd29UeFntOyuBmzsZzWJdKt0fDXLdalYvbHhQ7rA
gzzE5GNlo7YhIs/mzP+F1cgxiOWf+hzL0vLmIxwX8sRp9cUhZm/HyLFcc1SFSudj
ZZ++VHumu96gJoDBTrJZBjONgkNJYOfC/rYAP5KXhiExta2EohhtMjyaD14FgTwE
rgCtugGiidcqykUrHVNL7h3bGakqSptm+1W1qAoPnAGwKVm0xGbB9ZlIg99QCQAu
piewe5zx7dordxY7hf55TTW7cvW+z9L2b9FRXoGus/wyMBUMY+NCz8DJ8aCjZ/RE
syImVEANq1LEe3/gXpPdeQX1sq3CqDnv6nqj5G42tID1oRx2R3TuIeNuBWVVq/8Y
Az+bZGuPKXDa0y4Q8uD5R5YXBmkZ97PEazUxvPcn/MAl3a4m/++VPLfmAiMox5MW
My5rRFaYJJeBng7jK33NquO+E3LuqTgETbkmimtsti1yDmwIAMPyYnd3aHh11xej
fLgUZEmCGgRBCSP8P5/1zwnOA3utLQ67ThVy9UYGQYSxiEM2hXJEZfFHlPAkzbjT
KMJYHoYdidjC1cU95z11ttEEsBFjwJB/84puhGOZ95dQku4MY0n7aozhdUNjouNB
1QtASWsJqrf25TkjS5sgsVS6L7n8rsOJ+0zgDHbpmyhtO3qQZTTrrW3rcdYV9s+B
D+HbJVAKF8hGUIBJPHTfNoFTB1ae1k6dHvrB35wZakE8ey2/PiNNfKFdino5lWXU
v6s4cc5euk151F7MeKSLs85YDBCjrmQH8P/+m35wtNheajDVbPBp0iEGpZ04js2B
iFcGKD30l6x2GYUKupxrTpAavCxK3UDEMT3e0EgW2Vb4rcxAyWS9D+IRTtkg0/pj
i0//tSpkb9s/JGOpN8k/xi7L0771hFpT/VD6RLRh3P4LthOAvtGVmtDnJgNRgjUQ
Vx3i9BlI1SPC1HnOx1v8btJkXcbTk/qMGHPyMVI+Y3Yx/vd/LjTHvZKi6+EzZjSy
Den+SohEgrPX3+zV1ikZlo1FTsQTS6tZ4UV1zofpIbMGJEEvjdMSqlkMpimOSwCY
6wwTmdIfSE/z4xZxviKsIW1A62tRdCkTtHAv/Zd/CJM5eEGsVH7pYzykkXjQjTWO
AAr++DeDnmKBiuHv0vJdLG8QPVQHVRL+agH4vcZ+ekOD51k8oun2WzFyIyj7f8ga
S9GBmX7mfzWnQAqI64aJ+WoYjhiJTmFl4XphPJan+P7h9V2AGc/VcBLXzJp2AZdz
SFJV8ERifoOXCLQneSCWzwS7Qhhx2SdffZoZXtmFHYy2178TmOlIZ9bwqIXk1DTj
0jWPPaFKMTeCU6BX8kaLetF2ncNFvggV2BSG2BjDj1h0w5FGeldSlmg+kxt+6F8p
3dHE0v9owmF7R9SBj0NLqkKFlxvJa76xcWFoHBq2Tk5nI54tRofFiYOreGQhFth6
TV7zLdglnKFQhIa26cxTZSqrnX46N0pWqap1fAID2IxmRC+W1T+AXXVz/HDX465G
2+VnSOxTICgA1Sw9hZqEHYu8a+suBhXPdAwcmY/0BbXdY8SE+0GcYAPFhVkemPCL
DtgDbyUivh4yxgyd8rLh+eQrkWtZZxHiWSBQvROzgi5uDcaw75aAPBtF/pnUvhvx
/iSnB0YsqNmZeZMBCZPPsBpHcaFjcR/XKxExuQEZDHhgEeqXd+d+zLOM4ubPTw9Z
tu2XcPbSZB8ijfooZsAoA9Tf02GidY/cwXYw3L0k26r9onZGc5LaEqGM2d/smLMT
grssxpc6KgqX6q5ylCDfwqWT85dnnL3ysTSv1PZiWichS4NVidHaeZ0+F9aTktN5
X5B64YGSsiO0fUlMYQzFtIoAzNo+WnOqrQRLASM5xe/L8prAecA4QzosTRQ8XhOv
+xc1VPV696h7/JBTWzI25xFw9/3d+HzdGsVrZwKAYPJ1IxLDEodtZFTkWOzsyVkK
6JKUNRTmwhoslJxONpfwVdgdpjttfQ9aiblTnrYNNpoeOc7ivfncgucd1VWY5YKK
CzN0VCJqBNUs244iBMj5AXruH4ks2UOUlb97LZt35zTOtIpJSSllIboKj3GvwfQE
d0YghWYQ3kCg6W6p5LKp9x/TjybpDGrXSg3+MdizAA7fadoQuHTCylWrhk0AO7Ze
luxD7PM88N2kyBmD8YvJ7KVc6XVNRRkFrTwafbne6Z22tpiyMkxk3yVMlH1RhNFt
PAXHNCjaFkMVAIpm2ViRUXpzDiYDEqtGC2B4RJWePGXfpuUbCHPgxhZFauoKbTVK
AD+SwLNmKkVKIbA91J7cw0jTaHXP5OpHJTfG2oy8PtPkrXOXXXXpbP2Wb0nhskyh
C6/W/EooCCEceB75YdxhxbvqGgDv/2vi0bL4q9uka5N31WQOo8yPZ09Hivu/3IOF
gnOrv/03xC4OQGzTRg2WLq9VmzPviNgPHztDkBcOFGqiHAUvW1+AoajTVzMYw3E1
wOmR/ULW1A4LfAWWNDF/+RbiTZHoLGG6Irs3m2ZjOO1IVevdyKdi9uBlDnt5lUXz
tTQBQSDTJYdOGbQy8h67PWxYjXj7V4Ao0iD4GVVwd9zjwQAYNmGecUd/xLkDwG7g
sh39d1qyLQOrfi9Vxp69/7g1uhI5P1JGQVuVK+xdjEckHwaywyZ/ELMkrW3RokJV
1qeRek3WUzV5yd9cHB6cGYCJ14WEMLDOh8cCmz29SWwbddjSrs6PHtGMk2yCkLCX
BsSHnxzELqe3Hk60nyhFyjXAA40hZjgXKljUECVGsT3YPv96TDo9uHuCnId3Kqta
9LS58dvC9mJUMq47ePVArSCQgg/wnhWZKDW+wnEt7TAT08F2R6wCbrUiSGCwyu5K
hebNeAtxBIImNkwzKaCITsM+toD3X8YteA7DQMOAyao1Ul4T7GW3QBzAF7Af5gbK
PefpWgIH50dC+ywDS556jQ9+Dtd64/UkH4ulD0rPCX2DvxZIFRH0GGjVgJss+E39
CMZFe4g7cI1gdjkb0H9r/43cQdskxdv+/hUBjnKzFSez+GT7oDRb83o798be2Qaj
vaCebfj0+AMSmkedJVOzj7vD2R6mrq5hT65PaJQviBGTGNh0Ghdvwg3snfW/H1QG
nC2cIA3LtBgMNSH+vaBzW615KZcZY8AfrzutrL8JEBtOdWEXRpu/Dnolyaz5rZYL
Z2zfJnUi7oXYybqmBrUD+lkcxxExLwKK38C/BwsV2HPqry3dfKl12tyfC5Mzzk2C
8TmtorbiE2TNRUcxhAFnF8AT6YQdoZHXASLEEfE4LxMBwsJoifL5KJ1N4u6zSm7x
86ioFgsn7aaUhhkWP2XrBJ+8OANwL9pGSDym9Nqw6AYXjEhCYjqkuNat8O76myHU
ITa74K9JOdpedEVMJ6WXVNvrWjoxkJMdcVHiF926bZ4zgjFA/mR/xZpRKomsqPa1
VbkRqRQ3Y9I0lWtqdG+/mgUDQ8KljI6lDp6C+SZOoWuUY39vE8GsiPGY7M1YGEag
AnRqFs8/PFJpnvmhXf3fPP43S6FeVRA/Ylrz0k52BSWOZuNWtEP+nrbltiuezXs3
JO09F+IM2fz4vqkZItrvVnIS2yprPAh3QrhOjAtR0Vomq0DcSAJGHKJyjVMeYk3I
sSELe0+MEKOSiKydkXNjk7P5rlgKxgfHiGgQSOln5Bd7EVAgFVPXCI0t+dbwnh6F
vvE4Ijp42tr7SGz6s/l3xDH345zCLB6TT+0Z2xn7vYE4X5zj+FiKRlCnFr6fETaM
GHIWo0YejTt/eBp6CdmYj3FuTvdbj1f1ccmmS163QOPUA1BQOiouEDjYGr+O4XwB
PNp2lfOR6Bm3RTk8ST6d1zD4HtPmu/Y17IKfUk7wpdw6s/YCUeiWNXcweDrlNnpa
sRAGWydFo/bGIUMxVsdWxQRERG9Fb+pE1XZiTxBxX+qdUoYEqbUF/F/Y45uvgzku
LRLn4GffouQeovCQinH1jDHHNCYuomgfGDbqwvqKsJRo5/yz7UqSJOv7P2jot46n
fe54IlP8Yl72QygNG0d2x/d6ShJIFzi0lrTWx18qfLxWMJjXHOlcmvm4lRJMSCzq
6QHU3QFdU2siACecYx3AkLnQC0jwCERiHTiqrE4Qc8wEmlkNCFqDUuvrDekUDIg7
AklrhbKH2qmn5ISqcjFRKRDzHNg/XU5J1A2tJkgkEziPT+Kv28ucy5HiAt9IGpYb
ylVzW4MBU1T8mh/dOreplb4UEZnQPZyP3kjowcDGm1FBYZNcEKVMjiufQu7meOOZ
rx0a6gguf8JG6kE2BlCdREdbbcPNhReFDy9mT6FM2edOtzdL2B32HVbR/iM0dUJG
+gd+ADeFbCLhP4IQ/KtGcnTSCBNTlkySvkZibXeLIxOPfHYTObUArjCVNfsXEhNp
WFAJ0UI6f/Xf5rIe4JiennbbriKGL+TTqe0haW7ff+adlzp1Dpq39Pi1umtpGhWK
0QZEMzcbfEfo26a3n+eIEilyLOyqinq+9GfldQwaUrstlEYt4ZTWTft/CFeQ2P9k
RH97GmycGicMm9weeI7fzVYu+4BJSQZtszVsBzTsnXhDzps7SoBlCD9bVCzgQf+q
3jWazdLRZjq4vkuB31nT+M/YW4bwzA70UNTUF7yyjnU7ctu8nk4xR+YQIgz650wZ
Iv+b6Wwh5ksCM49OmPSAkx0DBjexst+zYp/RhCQQFZWlxbWfzsN9tG7VL8IITBR7
VX7KIOVZ46vzpHbuB6SuqeOYWr66G1WH6gjcSR6Q02L8QXY6sqkVaSdLcQKAsX2T
ct3rcYPHS8cTiTJmYU6ikNDzjvTw6h6LhA3F0/ayLln90A2zqdA7nOtvYTssvpgc
0RkcXXMQuLuHdg9gPtyWtgkgHuQFSgnQh8EDgNjd/9y9fvW6LqAR7dUd4934zF4U
WJ52dO1fzvbX8lsEBotoTikpNPhcD1UFkqw9b617MECGWteNvAsoQB/MKdt1VJ9b
aCHbkD2nS8BOz/Q7D3nvW/ZZ13XJRTxDN3lLyYNBvTlaa1h/337wU3/XvO1RzLgH
tTrSzU/haWTqU3Jz315zQvVw+A4bO/uk42+9pWYIHxgzrQSgvY8MjS8oo0oe7q4i
B7qszbKimlF4Mk6z6k0sliDs5E0D7/s4GunX2WiMPUE70yeF7nnyN3sYtKq8xySK
v+e9s1gBJaBY3DF0DOogt9+NrdBTmBeFClS2CcxE3Hi7ILAeSvY8UHEUZ9Bg9ABu
sVQupFdOqLHpD71FyvmT7MzoOWWbbSfIa1/UDq6S+D4a3K2FDrddW+xHiH+wV5H8
A5QiTluEJ2q7tgKhpEgVuuhbVLvv+DTyjXxriIAS7+x06UKeh4o0CJ6gFrbolhtH
0NnFDKGjR91G6PM9WEpDzBt/D2mGPsqFESuqLCnZ1LmMXEUGWs8+tSCTcWo2qfiX
IAmoVs5dr06bSFHFK+AnfEa2b4+LwaIhCH5cavV+zxyWPXxp0bVQNgNvQIqeGYAS
d5ESnTLJVGQadEt/NvCL2G6jDheHfWoRZoRMGlI5Rcp3Ytjx3qSwhnLKQLd/5QcJ
IqTajX8ByT1QT0DCM5mLQUi9aakjHq9uVaL1/bdj8AcyX5ae2Z9o+UVlz8qmaBEC
uVoyUxJNXTwAG5hzPjow/ybBEBBflbN1wgXrLGyQSGlM5Ktvn6X8epLIP1LxPeMc
7qU/RpfbvNjCTzUBpoa5BADqFvNP1NF4q7T/E0cbaD5pOvZpOz18cv7YII0DiU85
6mfFP1dMwfKj6BEgiNuooJlrvfeaUibc+tPwiiJF458V2y7YYxvHwQg6bfjOQSeV
TTzloeaZKHxu1wRsYmsbylyHeSYuMZx54MkiEBTIVvTccDvDVTXaW+LBUD9dk/ia
vnHH/jTP1Rke11Tr3QjaFYU6deCVgD+nMSge0/JTUeJ2Js8tffpI6hcnNdZWSRYG
KP6AXLBzO9wvCuOMf/TxqXms3r+TwieXqzDduHHWzIZJfGUWLh5Jv27qYRx+RUnF
ANiXveYNe5kmKe33SBQFhK8olOTLEuZgM4KxMmcqt3PGK5xqZYMf9YzQv4z9/7MX
EVMCGRoMfPpjpMfmuyFwNri56NuJPzHgFq2EpvHNU2W9bChssaL0KQWS/JPOoJLk
6qDl/RY4XlHFJfrrz4X/WpXCE2PbZdaWc/2YHopmicqXSVBeIIAlygHWbtRq7LqI
Uo08ObGRbuPUV1PYxwhy12feKi00Lemc8nzqLwD4a1KTkk8nObui1QKEYgJ1WD82
5IYb329W7/XdiB9sS2WMs5J9HN5lgfNlS/VJ6RSG6EM8zeWkGdwm3VInz/sWIPrC
qSywFkBZayOxbZVEvT1+kXjhmz7uIjbe+0P8xWW/rpU3Up2HOPpiiCBsH8LU2fJR
ZoabhrdYB4s+4gpZOlHpIbnu/n0lXtuJqXhObi2N6B1k39b+H1MTsmriKFvGuBxP
hmsOHO9CYTA9V/+Gb9Bb7+K+5Zve5ymewnfyR//tpZ9HNyIU8u1Yeem2cBt9Rb55
QZJe+TorGzfjSCdezAVkQ2+EqEfCOr6yUqWubY2SdOrbvcvHW/uE9V3RdHaVKg3a
V1rBhy439hIVop7tR5vvnXvnc05EG+EoEjVurgnzghb+YXlef6Y17bI5GzEXBk7O
xzak0lff/vJe7sq8SabiDrCVomRNTPUeiPqbDtw9Sy1UB6LOkx0OogUcIjHz++86
F6XRCx0Ygh+hYoWymwLcsXutKdxKbsFSkw0nFH1Tz0SzcadX1DgisX8CTUQ+uF/r
NTbgKo7TczlyekKv0C4aRWQJWwIr2GyBCzTaibXmuTxI0xOxf1NNs5AVuv2eg1kh
vmmMqWS5gKcOHnadFIK8oLS/k/7Upb0fNJaQws8j5K2b9LQREUfGtRX9kXkOcsTl
vpkUqCTfG4bkSujpwEhZcUtf9kpPK5n2gBtcVlZZTANR+cpiyq+whZDtqkoWGXz8
lHjNRXqtw9adUIQ/KFtrpQ5Wlb/McAWwtMTdM6yw+f0xT4kYP33ivy6hMuIGlXcQ
92laB5xH9u6VLlKXPg/US+0jyvABn8tn2l6H0xAEN2uqX3KkQ1j+Wkd49Kp4xAeO
6QsZe6i/P6CPaGvRuSPR+BzrNwzkFX2qpTkZxPuE2aqo/0uQx8ji/cUI3MU2K2R2
nGPfISJq/gN8Vp7PnHN0Ue8hd7vCEgBOKpBYT7Ruz4P7ui21VGZgoIZcMd2flhQR
KJ7rAN08cG8urwx0eOm+q0oZ2qR2g3XYdsYNVPh00V1mQjYx/9AhSOpNdfYsDoVS
3CKRnoUa9NRh60g994H5xxNdJnpy8h4Eh1F4B3fAsbSvL6Id/bdmOYUVKWtNXdl8
9f4388mCqAIDhJx4/p4e7Q0Whmv86U2LbptjQRkwqIK5hxASOvUruuf28ZsgABHO
SOXw/lZorPeWV6A1A9LoaCQdZMM7/M/yHwYfp08sID5t1zSd8HGjnRwHyMfZYM/0
Wjkdot59+I1+nsLfiRLJgwqs4VzGYRiK5uC3sGxNoLjmrbW3frqfzPC+/GT1Rh0g
WGmeJZpbqZMuufwf0GAIKeNZisQCvwUOytSp/XO2jbfyTy49fyMJoS4U49PaFgSp
fGemKp1YcCuMalKZIHF3KTkZhR9EeOEEWEBSOjtnj3dhclurW3hbpli78b6wWzVj
JEMWIUtFoIzUQDo9FXvaoVaVgg/3IcLqcBR8l/zhh9/5eKzEADPffi4HhpL4I2dp
otVtjsv1qW1stUsOMWK3vkT4vUKmGAGUskDEKucts/Hw9domK/ujosYPYb1KPMPu
R2AcvSk0I9weBEVZWGqTZ90HR3ntHopWPlVznqeNht3bHhrakpaCfW+lYrucbisz
H9fOIBsSJ+HAN4QQ7OOdNCWRDERuoQ8zCy7gPSZYFVqov/I+9mxNRm+4XG06WuN1
WbRWxHI4Ii3I0LxrJ6lautPEWHX5MG4E9TnLKyJMFzOgioRAhEu6M0zvJ+WhUhwj
vV/6Eq5ReOWX3RKfKvOxg9fAxaWHlf5n6BFwqmKQt/LG5N75gOYCE/O2C7IIW510
AbEBQA+M0ZzRfZym9mosGWjAboMGNx4bPRrN2/VFUeeEXTjzAKgqgupQRaOmvzfu
yqQ8CgmZygS9KyFEpcmq2GDW/kcQT35yXArMd9WEZm9wPkgxMzTu2TXJY7N9a674
1awlC8RUyu65mzEeJq/Cm/fv2Gf4fcddzrR3CI4ZscZ2qdKcxjDm51Q2seSCBWnn
HWcUTzIOKxP2+rb5MOHCFlogNI9WiNrdB/6k35qCsGh8kl6qmC7QP6k/ZT8ebgL9
VLbq+BcV9aPgynTAAxaux3B4AGnDdmUedWv+jhI0j+kvoVOfL69wrnb1cmY8FgJV
jK7WElyaxBf6uTsj3smyglyjXyrf4wPjVF+uDhPt+AOlAkoWcKvGs0iDIZ4E4y81
7uyJpNIPdWmWc9znxiiuAHlEXQ11PlQC7erKrKXl3rfUXMvuA3u0nueDbbI1hd3x
Nwgnk9f6emyu0hteGEvJefAw9B+c8dCXk9vFFaEqEkM5uZkpujO1Iws0jAHkeBP6
7NSQsADKR5bnbLHqcF6Zu6K/HzvgAUJIr4hgOH8f+Lq12M2TXNQzltFdB2gkRVHm
9mN9hKZMJGVSGeSMQnnI2EMH5TEg1patV3GgUR/fjaajzPaSchnY2xJMqKO5AuKT
Od71ymZeGDvV6JnexZVhJfxi1k1cJCtocfN7oGIrPdGuGz97LkAN/rbIduWiLsWg
J5RbEatUEgVQ0PjJfPz78YqupEgLmJ4BFNl+YfkGgJ6mz8eEmrlPnznDiOmWF4le
ocFFRCM2zuXMcQeJttALReQI6MHbxfi4nBd9s1GWvexe+eej/jJF6OxZBiRWZOtf
HCiSk7wUre3MP3G4/cR+agamyloDNWcw72S80by3j1D2L6Z72XfgyyIpxfF+ugmg
7Q/dJndpvpAVEqy5QbhvMpyQmU2EV3Re+tXG+f1DdIUvAcmKbf6u0KVqnFSGE07y
ByzIndWkUXAA/4NO0Z9wHb3NQMWfjjh//Qehcd/IfOY=
`protect END_PROTECTED
