`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KwToxW3i4yJMea89gDMrKXLC3c/z8QeiQq0hbTZ8ALqg04Xd/NM7tCTOLUrCbnhN
HX2XHggG45iLAV7WB0O0Qi0Nk0P0kQAYEo/kYYkJy1EkAXOP55GVk2sMODejjJq3
aQU8yjQvRYgtQVZJ6zyNxR7aCjNgmr1PmaKTOqtmmIm31nfH3xy5c+V/vJuxBQ9/
T7SPOfrGgUark0LiSQGOjopoWoUcZz9heHjQvtQYgoeSkIfBWcn2pXU9h/8ABc2k
g3mk/EmG/LPzizCuGi84kp9yb28ys5BLaT+TQxSkuck7JHdKmbgPFusGD7rdj6yR
O1HkZOynwX36RDShskEpgaaIO6g01pjM+3yBgkHpprcbGsQPpEyZl8DBKv6oUrds
i/wTx3tlrr7Bow0/vO7MlwuqTX1EIIkdWt37Y6Pc1OHQKKWQA/UUACEM82EMJX3O
PzlmwQlUrAKSaGJSaYUdIw0aOrH/8toGATJurTC5AtQo5AQkQuqzvEc7bDvHlVec
StkcU/c+ZXOCsvTUHtlx6yjJ5NVNrvdaQTvuzikIiX7/MNcKaCthpogoD4AAXfCM
sHxS6vmzXC8RYWbXTBvkaxK7LLvCoF53rE8XTZYwgPaO4UmQyRngA3tuWOiCbynI
HsPSpSSFcLvfhVRmiFj/eYRUSCw70vIaTI56BPWN/jZcOPo9DdTpLJTzd8HLiX2W
a1wnqQfZJokBrmUzfoXk4M5ok/ZbL5yrtaiBWCnsxQIxiiqt2CLhClmDoFWODWql
2IyZKh3fcDCIYzTwXtY13YjY28SRJpYY1CQhfvvyudzsKyvWIVRbAsRQpHGt5iv2
G5Dy5CB18byVuMvFhJEgTf6C1nXKyeh+zGNLDhrZJPsLCcso5FRZbsc2UltzyLq7
sxhKpcpFrdrbZTAqV9jJphZ9UHjG2y2QoFNwGdz/eXT1UqZxVLCY4ZjQ4aB/b4zA
TTbTTwfzu4CGSw8ZWXgZbOdCpafACjtKcrdaMZOhtsAJGH4LW197BzTlPo6jygL4
QcecksFJcxJHywENYUITyBNw8r99uTFzGttxVTN3x3Q5Bo+iX1wY+e5mPDI2KPaK
W9pjDEOwIeNQgURrqq1tzMgKlzB03kR6TDmH5UaG+2rxS8N5XbuW3xpnfEwel2Xd
0ALd0ttcZnhpW0C7Kf7ttCm0P4PjvX/ULIdXJQchipJoVYOufxY8o2jofWTCuokp
fLPv/DGv79bNf0Vqm4z6FTv4xEXFAVBjFxpijcxmjLg=
`protect END_PROTECTED
