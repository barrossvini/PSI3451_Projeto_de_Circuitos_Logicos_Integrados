`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1ca8c3dRuGEIZHSw4qC6kPWyf8f0ObzrO56J15BqJntr5kf3N8s24fM5V7qe1YQ
gGDmIXXKiapao7QDf/81dskxUvh0m2n9Zg905NP8qzkwWAg+gRPp5V0VgyyAIk99
LxsXFTjfK0y0Ajb1YPkBx+jKAqKE39VEuoyw0GKXaVj4HxkSlIo1r+DeHaa4nA5s
WveQcm7zNKdfIbYSi4fIygFkKiWcjhzWemADEenjXWqaOeMAvVqD9EOcbmoA1zzk
G0zjpe5iInNy0qRtC+qyT2HMjy8l/AvH93wErH2s2eoWHNnODBA6Fy8rmgYlXFWG
ndaACJpzHkjvYRCbqR7brbWK272GgARlUh+8K4AMBl67fHhmhpmwcjp2IgRm+K40
ezsQHrIMbbaP63Pr9ddhZ0xY5oae70ZvtEgEC349EgcvEG95NNPZhEuOu4LUryws
D4FHq8nWeUrbW8aJpJDm70QNXca/LX7+P0OpTcP81fzww2mfH9uAMjBExjwugFDx
TC5hNm1yUKZkiVdDn7XYloTbwUPJ1MoA6IPEsYW5wy/S4aX+h3/Oi88lIZCq+v8h
eXRAttnMn4ABNGrtfcwkZQozw1G0FvyCXZKtO4anSMb9faWTKFTMJkiZcyIsvgOF
JOsome5DrW8y2UrXvtXDO6mAUaxppUA6spZYCPuDOYQFjCT8rdV6SaP7IuQ/KTlx
3cb2DfLsFI9r1LYUTKpOiHWNtXbBQboBstOd1VJf0Us=
`protect END_PROTECTED
