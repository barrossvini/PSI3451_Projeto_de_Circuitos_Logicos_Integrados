`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n4KBL5cCzq3a9g4znC6xbv8A87z9yrfH94INDSEATic6Usz3IAxygw3pHyjERp6N
ZGYOePe9kBgSDApbX9RthkV/Y5FujhBVdRtNhx5uTils9ko0QmD/ERqaMzeCXvnm
2k5qUcR1J6rKT1aClIQkWfw+26iohmQZ1OOUGCR1qOzDUBIw1RSjJKWCr5FsXqWb
7KPzeqmzs6NhfTRvFwqzvbCd9JU0QKEW843o3SKA9MPFzyq4fiz2Mfl+hk4AExCz
Fn7bGUrVDMrutsn/ruMVbG1b7WH0tlPxYYYG2bn5QaytoUBzDjpzBIUPScnFtxNq
MT7nHs0OOHq9PygpTQic9hhD8rswTQH4GHwthHKO7Om3OlvkVG60qfipDHUC64R9
+MVCe2Rre+ArZSoMm6c0nYzrE5euvzXJFYkMzJ135KAqMSJ5DFxzodcUR1byHLJu
rXuA+oFu0Jr4RdB6F/fOA0bblo36fkEFmo6awrIX/ZAS5RkN34wdeZZ6IvryJxyW
69zz9dnMTA9SYW/5EB3uvOIn2/uDEOq75rCnY5hnvAcGPbnsZi7FmvvxvyRiPrKh
YRVzyGr2qp6FVZ9wBcL/qsAM05uFwP4lQkLBflmnJLjiWKRGwOlTpUdQZUCip593
wQBghGquDbF+bOSLtZ9vRtciNnhoYo2gGFuQkNqG7IrICwaN7bA3tDmP8L3hjDbF
`protect END_PROTECTED
