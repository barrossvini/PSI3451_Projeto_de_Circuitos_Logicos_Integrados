`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypyFop9IKxXzeSMIdNLx/AxLqiZzFRYEHhVlZbJqtokFHdXFcp1Qn1k4JAz5t1Wi
HziTN0NOqiU6fz3/Nu6dyHWRVjd/qa8SU3QfY/dEQ3uKw/DFJofBH5/yx0D2dQzR
vyE+UanlGaHMy5JR7BwAcafsYpvQZ3yATFozNdVJN19xFPUq07RGerKYC1sjIIm6
xG9087DbKXo+7Qe6LpT16ndqN6UYZyXzps96fdBu0va4gnvAgpZLnlRiX9Se5On8
CUwGIZb+KNW1pqv1corctayJ6+w4nTDzbi/d1G4xyCgrV8ByvQIWu6d9Tq2ZMuz4
T7gW9isP1O3xexvo+4yj9A==
`protect END_PROTECTED
