`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q9EPAm+jrLvZhimXjR0vBQjDNwZl+ZEAGdPfDr2Jp+/ODXv/t1mR0I+lQjLRkMYp
l9Ib+zAwHLX6fbI8n79QbIdaR3uJj0tunNB9MvzsDOJJfp1CSe+b8uzgoLB1fxgm
9bz66fIW07OovMBzOPPJSNTkGS85vQ6d8a0jkTt1inguhr9C0ubf37RGId6qDVoY
D/3DfUmuq9SrYr0P+bLrN5kv2pvBsOchCOJvWjfiqrMVTHVja2M7zzfunO5BZaLB
A7lMpkzM0P7rqngKeEvAZZSjVmuu6MoZam2VVidB9h2qOukF7KiT+IV0+KlGu7Lm
ssyr1ErWFgiAA2pDyt4pZWE7/EuTEkgeLd01ppU7sY4FcRFPyP2VFlhqNhP5y6a/
mWwI53hhLtJstyce9GtxLa0xPh3vsYPACyDrkug6c4/NpzoWTIlDNJSejf0Zaf9X
krQn5tLRCa/cIaiChOp+2dat5NvSb8XHLygFPljJxt5act1uIYqvZiYJIU6Tjm+4
esz6rWxl7OqKbOXGwHsze97Ga+/U7bZL35U58ltZWhYTQehk4ru4our69NJ/4FH9
swJSytheHeCxJ5SOaCBYDoY3vDmIvrLPWDcR18au+cj17eTuGt4Ww3sj49EG/pu3
DhRwizIQ1umI96jaVBj70FCZDmUnEUdghfkup6Oxtb3WYPXtILo3rB6xDi/aQsO5
ryyQ8SnoWEczQF5GSBLb4iqBBgmqWJNByD01f8JUTD984FuU43k+BrPytsqxPjSz
3QnlC+JWDAyXyXLeKv8b1cHftrv6HYXjFT2+BLJMCzI/Xmfno5Ng+d69UjDRTVDM
giOcioKdCDRguNdarsiRyJf6Uh6ys5Dck+j77WqmB6kffZmap0WPBfgS+MC63X2A
iPCRQEWqHvYNNRDrXB1Dzao8Q9BwiohH/ezoJfMKoymnh1zwCBTpeC10S8C9ehbm
Q7+Hw/1bqbaiUlAPirVHQzT97UCEcj6M11gu5Uhrt3l5ug80xyizviUF9z7Q0S5f
CMH0mZqOA6Z0CY/xCUYywBcn6SFbFyeGS24tXKdCvmdOD1D2kr4W/z3K71lEjDON
7bNzQM1Z3YPbGx7kdEoaTef9+7GEqV7JBorunX34ZHlv/0JjCfjYZxDYIdE6FyGv
rdqKCtPyvkdHQ4RWY3Y4sH1f1TriKnzn5oK/it4nAwubn1CvvB9f07J0inQkYT6S
kDoo3SC2vCI7nHvxqJMLSR3Q8mnW1gKI5zd6soYtsFFWdDghcV0fas3WYItw4Dx4
SyY7lf329YNWtZz+Ektp5I8nvsvX0eoQlKZTlSthcV8ySDMeG0pA2/+uNOIAdDW0
/JvngM30kPqtco85iQ0GN85spu23GVaHyW4HW82h0Vj5VB3CGZWmKRVYE4EKMndr
0tyK1tTho+G+C+jdkmLOmpyC0BjwhMmZngI0uS3SpvXvv6K7OUxnZSefeFLoFPbR
Q+fm+rDOGIyhKSGOCkET5dX31xCPJ2CTqegyyWxXMZaUEupGQKed6zH2wvo0qmyH
jZE6BLUvzbLOmuzbR4TFLXVuDoi3a/b62fHfwZmV6mZRbGwpbeWy4fX5xwQeSTOh
KRvVM8Hs/fr172/0C/BV4rUcSzFGioPl6+XgRKcKR8ay8IyijZwv9sBERL32F+uR
3YtRZCndqhgnYXeWB31WIS2nVyfgNG3xsMfs3ivPtywFOo+ryZHvXeeogiwb9Zfi
DnGfVVMBpTYfgnOKgJargs7zXpttKCU5+90lbs0jlfG0CXrAXtr+CiBeZNfnoqXg
LxOuwTDJ+FXNatjFsim3o4qU+ikCj9w5FWKGkLltzE9k1LobRg56oJfofeKGyisM
pNslc36jYSdAVwK7pcJuRl24uPhLzHS6NyOX7cCiCf3edA7oJiE+sl+E/rlQ8n9D
/UEiesoUqZaIwVLGuZt3c8p8BiA3fjtcV0iGMGYf4eGaEaWzUNL6R2XDF1hJF7uN
T/hYdHgseuMYGT2vZ+RNMGkk/Nq7Xu8dqWjNBGUNE/9MPjStqJEeA5p4zTXT59dY
AWnn9IwRIN7m2wXzMTCVYbfZnuAKl6e6vKB1e5h6pmFRkmovfqtnFkPJL72VCOO8
diIOpgcNVlmcuy05n7f0upxwrQI6duxDPEpBaI9GjaLkexJDaP4GRJ7yhmZR5IHP
llhjQ/l86zV4IlulioRtn2sFRw4L5w+CfQzGjxf5WQZH9GJDoO3nctM50p/mMyRJ
CCU4aVNU3DW/67XlatpiFw==
`protect END_PROTECTED
