`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3FJFLpO4fAAIQ175+TNwmB68BBNVaszmuKohkeeK4HTNGOjrj9cHTscBnLRWKFgI
6KqrrOMA0LSFW21aQehhLpyUrNyYhaaWtAQau5BxCi8HHiPvlCPkGK8Lj6bMB/7q
lkjdApWHEl3vZqKRKIgcA32aS7sg2ee0DDz/yzGInUuVxYjqO9ikYcfT9JUO+PaY
pbCyaK5VQU91cn1RP4B9+NTEMLreahQC70bMYdEbD4O9Pu6azbSEzetL1Ax/psEj
C0ifa+DXPpI7qdoqpcqmre6rL1DRlLFU+e2Y+Xh5r7wThje+eCSHXDadGByFLOj7
YEz9wwZk+iVuW1+9ofg159yUkPdlvA8tu4ruk88eN7bxRLHib2RZfQyLvUbQryQf
deB2O7BaRPbN9IYcEQC1vVzQXMOOMvPi+fiiymNgk+tslqs3hANuPOEonGYy3+7S
BMcu6iAT2phwUTQmvygvZK6rzzmYPrAORmjf4tNZ7s9pmVfkw4eTNjyGGFbFpn++
9Pb/vNZq39T3FZ8iFUUDgIqRbGvbrMHP4yzYWzTClioSneOEwZ5bqy1ahJfCfqNr
i3lTFYmmxz8/CaTs5/GqrWA72q/0vzFxe8mEakvDc+5jGsM4gjT5D2vcFFKvHRBH
94NBUNUPktYAqu2sYTsOJUH6vNk58g+AHsXUJSLhNblwGi0gby4HARLdLEnt7pwO
qDxJHArH5HgDSpxXPFR2b3osvrbncTqYpbwduzvIP6Vf7o0cFbcwS59HYTbJ3zj2
uF0LdtVI1+Q5hRGAWjp5yecsvdrdbe6r/EA2PPWwmOIew3mznEcoTuoxxdEiUqwM
KnBrnF5AihCgSRT/btO5tkMGHQ7hFenwoPzItpEqh5//eABxnrxOydlCWDGq+mBu
lkIK4vJTd8VZskEOpnIJ3FBnBRDIi5btWIdvFyFOCNIn1J4bC847y93q3NUO0fut
aCkhfbj66aPtnQYQ7Ow/b7teVSD8DU9TZssbtEARJy1gJO4pxyR+kcyxCVHfFMEV
ZT/LyzSzoqrINd/QHCc9zJfTNaa9KuJBbwhaaKkOIWiqVFl96oZnpXBpiAWuz9Vk
kbE9ZHGtM+qy1Bl/6K1ADPkhgWnOiB0KLX2hO2dznynVauzcmQlj0Up3hSp55tPg
vcE4h9mI5rk4sB4KhOROhmDfSBgJz9F7eoZ+k4rzVPdMy7bhgdxnfTHhKQuqwqRE
`protect END_PROTECTED
