`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BY/vvLgfqXiKqyR2DEFKLf9vC2hn9gr2LBg2efD5I10dxpxlr+ew/NXXJjIGsyOK
HzsVTdwfArZrvdI8uIfpFK7HpAxH15ssIb+qDE4TUikUubZzvM2+vIaQwRt5hHem
KeoRYHAw/z8Dri9kOxIYYyobqQoKCAtXrq1WxAIp9q9nCTnKyb9hM26Gr85/3O+v
bfPCfoyBro2/nlvVMsAj5HguFsELzEM0/Pl0R+Qt2ei58sXQXsz5IxQOrusrDIQ4
oAYR0825jeGlcY7ot7ZUnGzmzSa03N54aD2O/VDsoyD9AWL8pUdLEewpdBVz1QJl
LbSUlW+qcPjkN5p66eJs5Ndn/63Ci03DLL/hYxkDgV3w4Pbj+9r5ND7aX/ztay3t
kyi5EKwiqj++Z3q3F+FrphiwT6ugV2xYGmYaIKpVUBCf7SplYFFyJ0fA6T4aLJT3
OTHPJkeG3uADxeSM4HQVrjaFYDDg54YjjrtYLXOaKq8xhL8uoFu+Lw6E4j2lJbOl
BaKY5+0foj7CSAe8B0a4R2XkWo+1saMdOiMsS1miKQZuydXrI9Vtb7kioiCsNT2h
UCAlcs/INPjmdHX+wGTQjwxjpUmOo474+ZyMh+rn09qBRZS9p2vw4Z3xuLCIg9ep
kDgBW39V6Bh6BstTuYENhd5a7jDwatO+kMMZrDgrNMS1Ccj91uSaWeV9yOe2DmU0
aWNKrrNLsknDl4faperZ1qGYh4VLwrhQHNrVly9FJplcbdsTpFu6TxtdXiBJ4dcU
vWrL6Spj3k1aL3NQ9O1R/uKD74ksoHFqj6w/71gxLdaEwvy0hLwj+8jc2dlCpLTu
f3L4+Vi5fIwRDJ0hqq+Z47+hnzg0yC/1VDd5Khgks6cqVzCBQKosJh9qniybmO5a
QGZ1RcM5/qDXiAgi0e1XN/gOI/7GO//BcKk8q+7vHGZnjRcqj4YxxOPNCu49I6Et
hYaPx2EZwu7SU9fQ5yT3wcPMWCTQe67RYcYm4/Cs960dVFEQZphnlE9S/4H4hOGq
bpIO3y0cUrCS/H1JfxKawXuin07fzWis45XXZoauyBYilE0a4fwr0decRdIVjWHo
77WHuhfQIIhqkt+TaNl2pBUG2lNJgw9HcLPWqJxKM7DesU1mr9RkYqNToHau2V9z
hl2RH5e0jxdlQce1RdAuTlvGAZwsP8zG70p6pTqt+Zo7JyjMdfqbZcWfIEQ+8OEN
oAvawwCH2Un3iVW8hywqb+6nHZMGzVIYx1o8wzYUcrO1vFrauiVo4tiv3fDko3DU
hIyxDvCcazHdOMlh7Ez6dEX7UdyOUXNkLHz8LgdxqvhOK4j5vI7GKA4MwIGADY/I
VhYCzaGQWGiOtl4wJRAwvr5Z0ci2Ulfmg6mQVSwYyy2tRPGzBSdMj4c0B2ZdEJyO
YR40uc1UYZKWydEsugwbhjp9R6tswCTheSQW0xv4kp2Di+Ufas6mqOpFggWjdEP1
zrFTGLDzFEAilUXBBV+sR3iMk3iFHU5snsOXMp8mkSW4rWME1WQYMVaosaqXfdkM
9QLjLQQU4C+8iPOP3UtcLJqsulA9yvf28uLsjV55DGbQa9CKUaPMSgs6ydaHasuz
HfJ5q4DYIL4k0Lwgeth/+zATE1AHSbQvF50X0eELPA/o+r4RHNSGNZIT0IzZDlic
SZDyK25tZN3P9TvQXiIz6eULq/y6pqZdSjQSmw2d/T4pnIhtQ4Ugve4i8IgHBaF4
YYCHTDWad0xXX0nWheCxLvg6/qaCkrmUbldfKRfDO1c9jsJFIr1BwqhocTtJKGNT
OE/ASOvsOM+1E2WOKw3mxUzn0ZeO55A6+EVzd4krXzTtAbnjgJ0G1pmBxGX7JVWo
+1Z9byXPf1Ww0CzsKp0ke3BS0dUTfGvXv9BiAqy/I2sKaK/wxiLWC0U6iOuWV3Mx
WcHTH1wWRaM7PSCPrlyP6Gnzw9Bn8mMRmqNOTBsRkqcgunfboYBdxBUDLQw6qU2/
nM14egf7IMGB74AhTLV9DWNz2gM8Ga8Of8dNSTnPaw6GF45g2mmO0tRpPw0NQ4dP
8VOrQZR1vqnpUGo3llxBTTwTW37KnKSoEOyQG1ANeuUkWjuILeUrL0s3kCc7GsGY
PF8ArujVQX4VErjeMkp6Vn+eS0i8SpU5eLD2JdNwRxl25Bt55gBvOM8UyahCq22Y
r7hx0B9c/xyna0QX4Ln4ik+IrYExvob5cMSriG0I9jYE2Pq3YRR0z8OXlgrzDqz4
USsBnTepM2F6cyUje8lbKOMKF/VYLs8WuSsTehAk++StYh0gO7VuvpTRJgbKZxNb
xGYe2yDgVXXaprK5InilqLYk0gMYusrASnawqXvK/JsliYHmjt3QNHbRtfR4+BIY
GBjwSjidm8htNTFCDBee6NzVHtC3OYm6wiqhMt0ZEaVVlBKLscVxvlE6l1RojNlJ
8U8m9asjNPnRlh6q2sM/qqg7NdhhgZ9bTaWlriX38JbdRYszXqLXgupQKNo3IYe4
XMdRKwmEDGI+wNmODYPzUqmV9nCNl3b0T0HKbGCoFsUHxPpIYGpzXLZV9kE4BJvf
LRQYgtJ6Occ6Xsah2rjrzMU63bhNBzgaUVCg6xWtK+JCxn5R1mnueJjEVxa5jDUb
GDb5fYewvqUBGwykSb/04B7Wy9jTW5eb1OXTY9E2JFNV3VqOx0k7uK2K9u+WJbMt
xFEqhlz7ze7aTyzrF1ORjblulCVbRlGwgpzfAzI3OimMWXx4X//Ett9urQqzvjd1
HJvUyhWKM8I5sRYoPo+QymnPcO7P1L24euiD1Hi3O99WZKbKqBnMKJTCm0vfaReo
R7xBhTLvX59alIA0kdjvdiQcBTyXUvskIPDoyGrdkeZpKFpXaE6X6JRe+dl/0Nzz
iMBcLJYSELbNHbi9z+uPZmouWqo0CS4Ez5Ob77dPVSwMw33Lez8ogjD8QLOKsl28
FWAApeRTfnNvMUvpJ/ZwQVCyvp4stfUbMNIoeYqR033jPEKJ2fR4ayyadj6QgIvM
rZfcZPOqNG4HO3EHvEb3bdDuwKQXgryACBrKzS1TnLuDvK7FPaHoa8QAE8CUlAZq
g+lJVnhpyZnASdQUE717mB2VEYpTCdRPrkHUCrVK0a41ppuQrIttN7d4NmgCLG1q
7Ky0yTZsp71cvZJfp2xTArmo8iewms6n9lZUnQT18b3joT2RGiG1bWWfjMqZhtB9
vfi+lS6WBcvEKoHMS+xNpEoitmsxgCtHysoyO0wzv85zeVGjqOAEopZt73KReUk7
j0ARuCwfE3YAGkhsuB4H7wMD9vO7JyIn5OQU5AZtdl4ggDnh3b8AS+v3n6Rvnmm1
zohl0Jqa14xpsFVzqDPd8NwtJH7CsmwNDkK0HvEFj5m8Tg0Ho9/83lN8qNNwuOX9
43capfDuqs9Zbr25vhaH8fLSGbCjcpEOJK92FVxKsSFWsIvXoD9x9H09g84/Zc6J
zGmFztypJjJY8DRKTCdHWBeFouNsmNF/9WkXuDnC9/JeOnhZ30ynUleGhS0A//lN
7dFKMmjrMJ/dGsBqR+aOeN5r7EjjeUfEnYaZwQknnXl/fk7+BXRqca+sipSTGiO2
J178vZ2E5lAxx7Pbe4PII9MjATkqagVDfD88+kxhjn7TnL+ZScT7gD4/zTSVpfKq
sx4/hMv5Q7jqrAc4IoYTtnjVrA+7k49Oj/MIqoOLxr6Jmb5UjwmbuQ4jEMhN2AIU
1+gDWRfK4upyK3tSQSKa8n0D2PEt9S6Saa0GcQr5wd17HqbqBAfMmOE7Rki7/et+
TdOfYy0fsB5ZRrWnrjj7Na/EjgWU46594VbOlgu4e+trQmxKvI3v9jF+cH7qKlFI
CTlDydET/M7A7pyzFP020CSpqR9/S7xAzQwoqTjl/Me7F8ZKRpWeEXvX5qjpIziR
4gd0RT64RYgkmazDdLtccptrj+1Cm+0zoWO9lkbC8DNt6qnMThw9hxA1pA8NMpzO
z2/F1y7wC+f1jf0Od15IbggXsaeqHIl8Y3p3Ia4tVDJIF1A8k7uiw5OmJ8QMnxBB
BdT324mLC+Y9sj9nsWXmTRFJ5BNn6ZLNWrtxe4+9OIfj5uTi1/YbxjxNTqE0jFp5
/Bf1fb5nu5r4+1SL+m3cSQgGThctovjPBqFrGgs9daTfaRQYIg75Xo5M+ZLx1la3
WKy5i7AqdCN4saYc2ov7S0AByweI3Zggk3pajeY8sixDt6JWCztWLPlbc6mrqqCk
x2C2LU/2L1M6ofKihwRTF6CB6lnzzt8VxDMZDMf5jMLPIR9IDQmqbAZKppmkLpUA
yQhYzYBQqUvjciblS6wx1ohxPAEpwczQBWkUvt5z6pn87c/pSb07NAR54sQYuari
DD5k/YNSl+r6D3sccPmVJxcd09ZauIUVeCzc3PS7z66N4li4P9bAdwM/4VDYAqxb
Mbp0H6Po9GaJk4qOO2lKfu3kicIbfN8K/Y0AFVGUl3TNJgWCTH7gQRB6KzxpkqD+
uctm1WL3XfXZjEgvw+QDn9VDkzl/6etOYyixFy3+UxsQO9vZKBSbK5NhclyO0P2D
U9SunHt4uh/HQKYWA2Dm9DKqYo+DmUm3tz2/ZIGbepb1AesWKJyLBxV5tiHNpGkd
O91AMEJGSPPM5mrqpbRzbxKWlfs+AVnheQn1K8KPGQVK6NIYldXHceZjgLwb7t2d
R0yTRBa0CN3hQEL6S9eGOgQ0JTl7p8CbFfNyNeBVzIkBBF7CE9SdS/2A9p39fWZf
o3d0Efpdf06wD7kixdpMhf3GrHf5invyqMrszT+V5b6x0xSqUDZDBxNAH1NrUsi1
LSWrQb2HLLJtzyMBLjBfOmz+Em3eokXqidPUfgs7Ga4kuneso2jv0CZsC/Ul7yGc
dznKkYL+yzwXDQSzS0Jow7SpN31rEy1szl8dqsoG/vGItZ64c+XlPj5+rosNuDuT
8ifspBJ1Gw2IiCA82OLMP/NaaNuGXiUo1oouuX5FmYhORiqWFkQBoPu7ypaM+LsR
PAJsdI3ystcXTYi5AtHG4GyKDTL/Ex6l5SJa4BBoI6PrDiOqwT0TN5K6HJT0TGbk
Ms/SMMFNDhJDXSRgBIJ+fWTaeWd0gF/aoka6GN243t3xKkOJeYzSLFmXJmmtkzwx
Wj9R2+WC1oYaQWx3J18Q+OAkFVod7BUpGyfMq9NzxCAqeMx735z65muR8q1S+TMC
SutUPE700PvYlIVmC7cuDQdfY05kn9v+rTh1f3QSiyF/lXtC29qEgcviFywp09gF
kl6Lj4kdVUJd00hiq9+JWQwDP2zbrhOwsDbCH44bFIHaDMYlqEFU6BmRrQTyRmUe
eiUNGUstY6hGSTIJ3zYrzdNB0cK1Ju3gnBcGCzkZCxn7DjRyho2fVZzlOL6Hamne
WmLtbxcv6G2SJDNKBJ/nFlhxi2YBI9YfONChW+3BmVGA1lr7z+8DNAOyBirTlPka
pE73nFFTlxRmSFcriwToe+MqW536+VVKL5SsSEaLCNODP7U7VVrJaF5FIPZJQRGF
LmrkH07a6AEzuQo6bDgtOOp4UE5Jw5RsdKfR+xzS4ZEtOlYDrxQ8GnlZdEEVPHfD
Sl3wjUPQvAuBPmO48h7XKQRYHc0P0ZgVyxkhgHA7ytJP/8tgaIxmN8tznTOqjNRS
I3Dsl5fzxd8wlXF7aCi7bKzUPzEtmhK6q1Eig/FxSejUVmWhKOtZfybyDnYgYyNd
JLQ8sOSBCoNUM/6Ziwta6uEvOy09Stw+Hap0RoLpa/ZGNQCfhK66wOyonmz5vx3R
8k2Ffg+pwD2SMjA4L+Ab0gkV3kqrnK8gfMMoTL8bASn3iFRPApzpl7uaVMNFPZnl
2xsPrmvjMZjOi+KMw10u3AHqfpnrWZTLI9vDaqO+BBfHOrNVCCoevtTT/zVda/v3
QjYexl46hOuBeRRIJ0aAh4gnr2lwo645vjk1isMFGF623P5FIbNBHbTp7cel2KJ+
IE+FdaWFfPwZT/bhWcgrFOADpg1JJAFkluaWhdJaZOH0UVMSjVb1g0BvQjD4mnZy
cC1yV1gLTfEo+EY4l1C3/JfBzXJ9gUjpy9Xcp7OjRIvimo7d8Pk8ipPHT/T+DM1/
yFIOFogM3y8WZJAd6iNdXqIyk8Ex5KsX3i13dNcozDaURYaUNZmziU5D0QOPKZ63
uTcm/AO3R23ohmdhqCXQjYUSFE/zPUQGkJ+N1gxNycyFlJltcJ267+22YaCITITU
t5RAOwjpEWheuM02OTl1j19uiOlrGfCnKHS7epu3TTNJtk6IaqIEp2dgNXZZfBXW
tqlF3xrNE5+5w7UQMT6ZFluCkVySmXOYBiBEqyZl4Zg6Xcfm+j5t7/DWghs5lAdp
ck9spceF/3sjvw8EgVpTgES/doDiyxATU2nfIgkPKn///Hz0BqXnO8lHFU8plTj5
UpZGIpQGTCyDdoxt31iiHAUxOSz8qQicv3wSIE1zIfKK2jBy76FacdusyrYyO9ow
wRJA6Wbzr5lyC4lTNoBIcfYngwA8W/0+4cWmJtWm15CZhR1+X4Cd1fO4lC8199e4
vn9ANkEJ0JiuANbgHYiAvc+y8sPqWP1OSTYF+Y1VrGxLVAt6RaiEZNJ1aRa0lr3b
yMzl28gQSnaNDfAwj95vD6ThlsmrhE42vvW++IBLxTEAq+BKpMMPez+ZfvYGMTfN
+HPwukbI4d9/8iTN/Kivn+iIKfswGAWOaep4X+NOCOLuYlzkOxT06hjTbqCEYCFt
+P9sPVQYDH/8TjIQQuMx650YiwD7uEek8iAK50F1G7pmG/ONMWD30WfMPX6Fy4JO
XHiricvVqtELnsKRnyyGvs4qvPkdk8zkzqdQAGLhhZ9HySf61mrUGQKMNZyN8jg9
/YoOLKTzkcc94hT2gDSF1xN0KxsGdDtrEgAP9UAXINYq6dx61r/iOQ0s8ZrLCR8Z
VAbXbv8noWB3LD0h0awpNeXu95oizaeSm7ua3JxmGPERb1MLNx2hGYw/Dv81+m3r
StC8IpmwyH9IAaawfVHhpS0zphCvGo3S9X7CcajbMn4ARDaUguShFl7azxb8DDEn
49nKdYM7OYIZvgPmAytPdO1fCU7zWHx0kGeNxUyM2YBzAxY2XpAwBWXw4Ihg1ehL
qD/Sb6RHLvICHsyC9ann+FF8GiF8ISMpAwhxQlmTn2+BnxRB7oH7EP1zQXsvrjZr
I+U1A+0hZmJw8igqSZSmCuT0lnmch5fO6FKYHBCAmG9bI6gIbcV/66TwtVCQhWRv
av7mVuMbR/OAPtQtlrtJ5RtaAZWJRRTvt0uJsl5KMfG3xfMtjl5yKbxa3bklccHE
nIHC48OY81aeyca2/lbgZ7jELs9qZmoR6J1YBgrUc0rWKfXHe/VHQ3AkaXwWtl7S
1+kbk8o1mjy56ozwrEO/XF9GP3Yz8+UNO6uAgQa4X/n0djbFG1MeYTV8AWt2VeTG
Bevjs5DBbG3+yMY/j5HID1QTMM21H48txBUdJmd4FopJE1D71l4eZE5vLcdxjFk4
tm/PeE64gJTiPALSxRK8B+JGSrSZIUKqeik9NE1PYrChMV1Ssga5r0Gtvq30oWW1
DK3qNNd4WTl+JLBGMTXj73ss0cpj4dGYHR36AcNbtaXrpgbz8/LggTPYUtewbhyS
Za0EYgywEydy/NKfBwyI6j3AJGG24FqsxhkCLUT1ru3gdr0hIrX+evju/ycZxzQE
xuidY+S892dYu2VdIjtjAfYRRW6IkzMH2Dx929vHagnNKCVO241q6owh+tXznPt+
/lN4UhzLVsXsqdg1niJLA7LumEca69CgRSKJeY/etQ3mve3eWZY7mVyJGkJbGF1y
cr3Tbb5gcxfZomjBcKzwmpe7wOTUt4lmFEm+mW7zycsEbChCa8rc2D9qandcwNQy
oLgeaHXl5jWkXHV7ftm/xzynpqsAYWkfLrm5bQY62JYruGWbIQ9sSrJuTetpoR15
jrI4KKfhO7Exj2bSsasPsZntnzPozUn4ga8Gx7x7RP5sLsbJJaMYu8arz6rQ2+cZ
CAOzUKbfxdXSD6iMd7S/Q8NEx+zXbYWQdhuDCkJFmRLnG1Tu437nur2ZqgmjgiV4
K3KHE7J4VaXtuDU6d/79ZbFLHCV70JjeCz0Z7gBIg/iPhYg9OJ9TuQsN0rQi6IIV
aKfwPzzczJ5SbQXKYsIRYaSbyis+MrtEZVR8VxAL/WGFd5W0RvIwd/CixD+muXzK
H9bnyaI+78vgAcwTQPiq0z4sbvA5hxjvRMgHUu5yaqsr8g2C5n0/VWlpWQzDfVpq
YXDjydRhmuvMxd+KjHuKG6kXFr/QbXHH0RwA5z88Dnbre8l7+JtGvgxCJKT8EM4H
3UW1JEYvRQPbc3F8JFr+uVqM7cJ4fAk+VVO24WxRlKlLn1X5m0hdomi5uePlx0hD
MLN44oGJA86ml/5lOZMsl1YBLLlGf1MdfJ17Ke5nZD4ofcCxuhF5XrOLTOnPboSC
11ao06f0xjKJMb4EE6yXFBu/qOUifi179w/uI+UovRr0qmhrlwsNT9AdSno5JMGb
oDwTAkVrlV8VNmi7bQzdnImWiZi+GtPb/9Uo8L+xdFdWZliAdti7H2/In8twgYlz
QlzhjREggjDZXRKsI5bmJqfpYvbr76EnaP5r1Z5R9/PStxj0/a2LohE0Cvz9X3jV
98iVq7XlLpR3avlQahsN++FoGJcf4DkZAmK3vcuZ/m5jo4U+J4TeCmqRylGF7t3v
jaxF8UWVyVm9fFCJQFScOCPEoIQUmGwFCqQ63dc0oXGTN1jM/q/2GZ0fxQONKP0Z
qWlRAwqyMo9rT+7LWW7Y29RR7l7st1f9dP0/bN75HKYX7z+8iKWbdJTiBBLw3Xcx
SXVYhy6kc4bi0dESjiK9ONBnC41gMO6Rl0wigcTPcgyF9tf4r2ubNzeWBv2ktyNP
hRKKUY5Le1Ty6Oh7Le/4qH9/hPfNL/PvCgEVtTnLtUmw0LrOiJy1HSKkOx7SK6ae
pVpjlo1/PzrBLAZa+XYFetIec2a/8UAoT0pmLYOX0ceABkLCwYnOXgSaU3qpkFsB
8/A72iKQivZb38PGu0bx2i/jXQbppnc9dyCt2wm8aScHxLH9SuH/DZMvUIwQNfc6
aaiE8LUyTRPlQRwKOVXhSx8wctxw8RQ//V8uSPHK4Jez/+sR6x1BU5o1Ml4UVeon
Vb9sX5JlGFhmSr6wbNxu7Ikj1c7hpqG9SpUD4pGMNu66xXkdy9R2UpduPZvuZGkN
oZYSOLV1zDylBKT/iUg3eeBIQVe2NSueiTMv8J4y8KuK4v2Su2rZaOeastjm26n0
JOmtYwocAAhn9DbjdrJdp0nUZksbAN5JOs1FnBJ/USlcT1o8gveWq2/GZPV0XwTr
6JHvFFAgeGAOUQauhNABbroQZiRkQq8Z1yavM0Q5UjOYx0h06xZb4DMK8g51Zbr+
tHA1OJDxc2iqhDUqgaYlsP1pOC7ATfAyCmQzxqdj+x/z+klFPOF3FyZmestTNWPV
FTq8BoV9jWXSMTsXbfFrZy+JYtkR5dsxxwrMhywhncqGo7rcWx9vzEBK+OCNYz3d
BoNuB0VJ5gmnAo/j8LsPXl7ft18Je6MTnYrNeaKxN2sire14WTQYg5aI5hJNDXUE
sWORKnZrO9gaK9YC47H3nuMJdWJN4/ZtEimt9TSfdMWjBDiNn2/c3bdNRhUiqLDt
oaaUpjCwheYOZUwc4PEsLBeC8KnHT+ZK3qNvAFi2uNIwYycxHFH6scLY4KEfJNlY
T5RkbGSG3OUH+VLLkwP+VUSX652af6pP8R2K0JwZppSPF4OjwYEvsgprwLNTXzSl
Ra7eOui/ahCgnKI6faGUiB7HIgWVK3b/yiXNWPFRMPB0jZA4cn9g21ilNTllYL47
RgWx+Eyhb2K72emU0IxhIxH4uYFbmuQFYMfqxxihiVlX3soz7Dzqtw9KacJ45rUi
mN7oW11RvXSHUHDmK3FsOFeje/SeWhHMtNbH4AN87nC6E3SDy24QmKXNBij+tFTa
2uuQLs4vP8bXsrHs8fA2xyKuOXePCsY+DV6ra8AjybFX//gPjU3vyKtXf0LwSZTU
SrRWA6jsTSH4P7VDdNraEKV0a/czt3VkqMfCRkVvH/sd1wRsu2oMbnFUlzN7iq5b
hnXi7/0YTqrWPXwrGK8RoqhmLAnhdL9ZAU0U9nmXJDaFSGnfuyVxOVQitfzRqWLb
eAWM+59gdx7aNNMVGfClVZiTlmsvPkeZYPrplUgNqENSatgotAywinZde5vIvHOI
Ax/vEgrHk01FKoCnTn58mBgNwOzP0p3xW1hcAyqCXr9BN2L9ey/XZUd9c6nltskj
9OGEhpfr+ZEr4AKdIJAlu/TxYflj2rMekJrAh/H1MhntncaDIbcGaRHWfRqXCvid
ANAnUUCmsvUUpefWDzA7tTIaSAhUSCY5XxznGHTl8/UDZAY4gkL3SiQ0l3A/+k4E
Ew3Bb3hw4Z1fxhYKcoKuWmCDK+v20rdnRX6qjl9WpZJo0fgJApz1Qdev7UTp6sdB
p7a9Xhu5kYrlhj9AgshmG4zpreF7kd4E4/rOnT7VGoJvNi4HAyjSEihK/mKBQxs6
9DrwL8ZDnlkp+J/HkWYRxoLaQiSDmXAsuDVsT46aeBhvLymTC28aZh1KveIzm8td
s+X30WMkL7dn9pL/3RYhnXuoTWK5ru2sRnvxEd8gaIDWgW/b/8xejfph4DGGmivL
3pfTv7N9ovpMhyMgszVKrwOMgFDh/cHTElsvuLNIJ352BLpo34XfchSxkDjk95wB
PKlnHOmii6TQC9jFTl5hLJxdChvDWoP18CHCAUxhbKYGeTWm0GhrsPQPmKI6cbAk
pGcvBitZbM7vmg9k5d7zj0eKXxkFJgASvICVCfG6boc92LiSyZLpUppmsqzbsNae
glDylyJKIDVml0KKUB4zXgjHD6BBYvT89qNXKramzu8c5zQx9L2QST+bZuvvE1+T
ly2x8EeWGIJjwc/k5Lbk9C/GHSp89aqmHvPMMtO2HGEjmNeVpl4I1psquRWQ5fw0
4+RuqRoc5qZO8Wq0kTCpPxvPXhS3KPKhCeluHQe5tFxn+nYP2v0Ny+V66bgcgrH5
YB3TC6ZolOQ9FSrsnbCx00/MOLIc2YvC7SF67rkjWwhunWxUVbGOz0Oh6q4DNuOO
Zt06eoZhz+RGAu+dERvgBdycop7ztTygNqX1RBY9l/BdBv53CbIdw+MkRf3Qk528
/d+K7+ZfFI3kheFqNwCkYtvDi/PYkpFp7JWJshhcCQD2zFlz+Snw7bi+DG9R526+
s7N5A7gWzpyfo4KhWeT0rGshiC1pO3bCbflXUVQDDn6fV+fRq3IW7KmzbS9C0SzV
A1qApEHHRZKKGO43WplaCe3tNDGPbU8G+z1TnyyPtb3E3A8WWZycENBAI383YSbl
5OOmrAoG1kTKdLiZvCrDit1XrYG2uqctC+tKV7qK73OUI5HZeADQmP6bN+stYKX+
2pT9hsya+4QwCSpLqykYnE1ie8rPsQInEHBqrU2P0vNn1W29xF7IKRVPNFbs821z
uGvRjiIzzT7u1FHPnGkRQfx7ApWYTrksa9dBBxjcGdwvUvgvS58o3BUMUZiRving
7dusIvhokWbjdzQyIyYLYybtqar7yU7hbA/igayJ06Q2xMsL/P5g+pIKgMbVCLS8
bsJclSLEGTb+uXwbur+CO08jJrZa4utjpQ4nZ3nz4lW9qDEzf7aHGicgwtMvOFhQ
gzyNTH6XM5AbXmTL/XwemwRyjwmLvKQ6yneVBeRHM+zdYG5Wzcf1H+X1jKktYW8+
ZDmw7ZqH+CCL3ZGqbHQ0lhBZuSVaORdFb6wxCZnT1RBk8NcRFTISFIK1qiPc/KGp
ip8mEE3U0lMZPle0Zmt9oRrdYdu6hc0ohuov32jJ55suBOusficfUo4v8GrKPWIF
sCuyW+LPmtB5+Qs7OKRu5N7u6+U6hl5wiCV/R/ek28s12bLo6Epx8OFfz7Pi4pQs
NIeNLSlr+LkuCU/4ZwF/GSKSbQtefvgj4ZfPZF3gpMH6QGGoflwsh+hqGHIdAatE
kw4ecJRJJ0QoY9uk+Bvc/3lVhqpsGRw4fH1Aa2iqhpYhBv8+yW+Zkf0viZQFdPOj
94glam44Xrb7lgVKsXfKbrduRGdDAqHk34aA+Ck/79sF3mJ1PdWpKf5GqEsLl/KH
BAbylt2nj+4Vijo7wSD4rRI2tX/TR76HiZ6AjlRcRGy9J6BhhPsWpjF1jNqaD35I
ZZlmK/nyYI6KZ9YZJqqygnOjQAqocrCQMyUM6zQdIZ0keSP7+vtcZJZObikMg+v8
ZdODva7okVwzmLTk189Q/eTCYcJKkDZqr6AkFk2sfrMp5sbG9Je6YGIcRdUVvHIo
s9RADOSZKqIr2lDS7libgwfYOChNpwY2fIxR/fCFBKRf9/rJGU8e10pkfNCTClje
zn9h8yn5MuFZI/4d8OuPI9apSLZ8qAXYUHWbF1IhcWF0Hv/Fo/mP7co86YPxzMT+
gJp8zK8uhSUEUyGILIJTLBEaWkkVRtXfgouppQX9y/IP3GOQZQEOiiGO+oWlm4dh
DGXVnBIKmkgw0Cp6WcidEIP/LfvNxNYMMyBrwd4SmsseqxfXSgHR7CU+hJ28iHcm
NrFRK3WOnXcOOMaDUNHhESHTpgFJrQPv1947ZLgi9le7M+GQbpeV3e56T/m+1aQ4
LpE1aJEdLgp8ZTpkondMEVtfuCAFumxDsGw2JKCamsQ6gt8PgQcudcVa2DtHrzYY
SgcQ9pEWysE54tJCv8y4rOuOvSGEyDKrYJh3sVt/LvmWX0RU1Q1UepWl9Oa8cfur
7a/ATEOBeLvI3TAFbBSeJ2rq1Av/6xZHA2t2z8UzBa3TU/2TF7ucW0nXFpxuCa1M
2hKJ4mM7wx17GX3j8S0v82T6iVtw4F7vVwztMOzvtzpG6AlOCmHvEi7TPXWfBk2p
8FCc84gMHihCt9NlWlSHs3XTTBhVJjpXWysrGu9EYT0pyAloiwD9psQPa9gvqRgQ
VU3zSOjHTw4StlFhthTk5D2LDRF2OHcSI3CFjVpHE13tUJOwxWvF12ehwBqHiaYc
SlTI+G+yD7RdKg+mh3kTE9r7shN1TmVINHgX738M0jby++hUwbY1RDByTmhe2CFq
+aSCgtbpGp2Q1RieY9pGRJj66qVYgcRwD1PBO6rw4ZZEzjVMejOnQuznBStJv1+U
K3Vk9R0HzbLvxQ4sqYFm3Yu+NmA1dIWJCwrfbBUy+7QIhxqFBGPaEX8A/wSZXxBM
/PfDbz8uwRllJvDZmVuWBBsCHvIUoqaQHhJ9zbbacisZKMPMzOv3zv0xy6vANrDT
wST0G0blpLbT4ObVvZF8TyVBrgyBDQHON7bmCQJWQo3ehpITKNThg2tnRoUTf9hw
nEwEb0Fo0o3Hj974Ip077svnqkAq1jXHF6zJKAq6BWzbsmAfumvlxkbsqTnJuQnv
AL+6H5u7fRAb09orONBh9NjT6UCfmyxoEc4cucd4xZQRawS70AfcU0cDmLefwBMi
GHlrmDNHg5tGs4HFfWlL/Il8UH5xSPkQzDAr32OeMyF/NXTMSek0CK087hOiWBuH
3sxK9cVPaTDQnoIH21wRIEBVqcNp+6PPb9fHDdnqyByQFzmz1YKO84bJMPBoBdMe
1S+80RKz4JoPqhDCN+FJNQxuP/tR4/ZoGZzTBBNQ5v9uuip+h3Ok51MZ153sEYj7
QWUrRt+Mm6AkPTk2CKxsDcuxJoW0Wfc2KyfYOsZ7VKE05BO5K5vAjtpWkCWs8Hbm
QacWp0jHtH0V0bi7kH09PFtRiayuLV3BzxudVFH6XywwkyL+c/6lPT312y4cupvI
zDUq3yMV1Tjl4dMwYKMPrzHryr4rt8z7qhMeSOgWwDZHJWrFOd4s5haxvaphVqRp
/LKTFacJVutuVLDMtjQaDgR/NReWWbo6zkc1WCtjSpLnGj0CHKcdEssjIN+w2HHy
Ye3x/fxacunKa+4YRZbCPczlmC9IJVW71ZaoYo16XNKG4kPMKihn0q/CRCY1bwmO
ofAiN5F4zxiCl+p+qubiGOuIXzXBwhslY3/TGQtS2SjWuvF5SjtE6gYcOlr5htNI
E7do0aVFLya8HIIXfTQN/2CJvdH/on0c/Ag8LMsI8f6ShDW9raATMakq/90bVXYJ
VTub+ba2VpgNh3GCSmjaApTzCjJM7iYIYI4dOIPEVnRI0g0rR6iGeD9Q2U+Waf54
HbOZqfYw9U/ElYN0LNkSI9BlUGVnqIcnwKChl13SKg/3g7vSJ1WZbwBUyS3pwON7
10mkMQPsBASSr8hnHSE2vdPtE2gNIZX6fc+HEnuAaGw6D4sZy/elejZ2Nq5vXceS
mLIkxC68iHPA+u5TQ+1jeiG2cobYILRhKbB3ek6CQZWLbKIqAIC75fAyIsUNynUv
L8tdoZ9pVlTPAxd+9M1EYpEDxPyOFPkzkTE0c2iwHUr+0XSR3UCaU80xGl00Vryu
Ig8qKefNI1KNsCeC80KeLNgTw20cCi+i6HOl9ueskCU/N64C29meGGRpHeH1z2Jl
8W1ZXyC7dxD832waOYA81h6gvPB7yQH7tGDUJKt5pyuw0EMfI4d96zj2XvavLS4q
B0sWyZIHS8Fn39LVQxG2IhM371C3auYYxgIPuj7x7kAZPoJbInlfhlzgSMd1pj+c
fgEwKCYWPL/NtRCPdGd3XzhLgNteAqexGbdBmAIUAnYvYC48W3f+g5D8/MSzHH2U
iiQvhaNHcC3iEHsLRDTGuDMIKcNExyhIM+4SatBr8eO+F1Sx1AkTc5QteYl1ZPql
DuSysK3JImViJnGMGlE7+HSt+QrnxQykvmHjCFYrgvh0oyiXWJtegcOeuvS7TmmX
bqfpxiwqRZoW8SfgM8O2bFpo7XjTcv69p323Yj2XkpWEoyl23/kv2kAV1dflQ4Jy
kdAq+CmuJK3RvrZisH2ip5nGLgo5mdbHrIOIhsV0HFOA1T8kqkXVr1JQ6zGbTP4L
MKaMKg9G1GThThpMiWWzz+ryHKCRyLAHnV+G3W2LSc/BzO+oitzkHGwve0H/VGeB
o//UQW3pqNoX1IrWzHSe8wJlNj/x/uBOG+d5H2wjkBspP4FT6inaQe23cXI+K3SY
CrTAycwBK3Yz8HJUBDI+njiOEdL/lTgr1jk8ZrSilx7ImVkgZxSrF2duhSFrbh0O
kg8UQOmwq1s8x5M0WZHjRI1/BmnMXDcoRRd44izN2SrSurHmm9AMnT8Z82/G1dtK
UBb1ONh2ZVdfPFaPyuShA6zOFR7Ed5IHMe0u0b/EAOsbl8Vy7OLzdWsHgXpGSiaK
Nnz91KeAqX5Xo+OxKASqsf3BesX44DsKV01RrwhL7EnyaWYBuoNsyW9qdKGMj5FJ
bkqzH58nPjDYBYOjeGkcqd79XAWJcCiICPCjvlJMrFcZNeNyCpOPOhHx8WxW8I8X
N0anDkKj/030Okq1cBq7SvfewOFEXuZzOF5Rxyc+dOMIn6waAqurOVyKqhFu1/Vv
hbcBI1/ki52JYxUMTICUU8cx6liZ8OA369jgnLYEQHCgeklmo5KLH1Pq6ynN02zP
/vMjCj80HtaTjubtRthjULlJYlq+7O4Psomrv7kw/vS8F7fXqdc7a7wIUHJpHnFH
+AD3uubCWBcW014grwvp2AplzQHyb9Avzb3J5Om+HxoXixZ6MYxNhwlxW217GGSC
NXPETbnSibs8hdG8gd1Kpnv9sUjIBmZ/JrrGwawbwJ+0b/Q5+AOD2Af7IPKUu8jR
KpXDe/Y2kRNjPRSH+erd3VYoK2KGSFC+Z/cvj7N5zlfiUrWoCjCVbqNlKvCU14Lp
M2fCASzDtSnvTEPQk7xbn+PVVJAuTPLmKL1+FZv3Llv/+54r9R1+hwjPpfORWNJ7
8cxvui50lcZrDdvDkZAWXxV+UjBfmFf5OuT3Phfy0FpVKaD3SD35VvRvL5i05I8T
4rEukDlOurIKLysLKdpo6LUi7YInFtBvY3oPqZvP9tj3y180DFxO2CyOnG0N6WTW
gNZe201v2cWfo1mlQpHh/YLx9Z2DDsfw6Fa4fxUxipzrjBk1mgRS8KBlnAwo06Ig
3YkdQnLfdrgb8PdFRMtIiLhqB2A2Oy3Vlk902Q35aPL0yBxjoxX4wURgM2ROjKlF
BeuNKbfgMN0PshHWI9hNyyuEqj4XHbWmcNjP3s/JD+OJoYbSQFgFxMEM2NA15wW5
JLIow7xcvumwTbOQP07oW0QJFiiFrrydhBbNiuyxKv/U3uUXNZOkQ0QX4f7H/m0B
IGo5PbzjOGTVE+8W9E5Bh6ZrNyTliAxd1OO03Y0COTWBT1CB7MniHLLwE3Ia7HDW
iZK5993lr+uDLLdVmyTl7T0Pvj7HqYvSjm08y2TG0Bm6ch0968cv0btlzzbaN3Bz
JLQPrxZEb4XLRvvnHR23kK/O/BDuFEzDfl6nWlV/PDuQ/zvYEyjaJgpdJOseIVRy
ZsWPg3MQ6XrRBdacMzvQqbd1BPDwixohpkQUpijDyroDYIyJpACp3MmT7nGbW39r
rYq0Jkd2FRVbecdJYEiA2jJU1GO9YKNKJchx7eZUmYm6IURDiZDQMYNWrQDL35tr
HOsZyeWyN/O6MlfHcFK9WeYEh4157VIvjfcMqa4/I+XxW/fynrdeyxG7JYFD+wJw
E5IXUMiWMNh33uv/+iVwjR0CkB8qVk8zd20Z7F1ptAJ+gcHLiNmquj6z+QgTzovx
+54XYKi8MTrs4FslCMFeQgdUiH2T26pyXM6Hp5b11+WEd4DOk59Js0tlhnBKeasS
4CxhljmxAjOGMzsGURflEZYF/osc8N96zSvCUg3WRGGXICP3WuQmfDKbX8C/LwUX
8c+0j92GIn+mn1UlK2ZsaXwee8kyR04vpPW/8SiBM1D/fQGQnHt7/S5tkmXr0w7F
zhuaZ/nCLvYNTG+BRB4RuQUnDlEWEkHJgN5K++QzKIinZ11/bSM2ln8NDre/UC87
Qs2gYrQhY3akyITaSm22M22kn9M72U7LBFSWhXnDsAlCNmcMLdXCejCpGj9TZr5E
hWL293W7gctdq+aCVoDOklmasNLEQy8r/TPVrZIuj74zZk/CDNy2EChQnsopTovQ
tJFKGMJwlD1/nTye/Fm1HhOTz7Y8hr4XF9+rCQi3MGcp5mK/1L15PxhzEQRKwdua
gPb1GwKysot8U6H0chycQ9AquZROfHnrnNDGW0kxIYftpIlyKjrPNCGWkWX3Gkmq
cCcLanwf1ndSMoODCdfWgB3VxUQ59cDsoiPP1OBU05A0r0MGlYZ6UhH7wPqPENOn
fg2HnHewUQnZcuPm+X/CUFIMS4ns53BjaKUNBDRU8l9nvdKpXAv7wfnRQERXABQ6
S1lgvGha3nTk1lDlIAs1QJPq4CQGBaCB3w0eeYgu+4iiomLdJ7GkDVznoxud/Aa8
hE5WnQc7ab2jkWDidaG/1waL0ksslajrOdL5jPuot20uyl9UZYZqKjhTgBN5DM64
9Sh/LMMEHgculTFONYLYdA07jO3JcIMY72s/Ycwieopx6c54NiR4H8js0cc7py9Y
f3d7rBds0bZyxuiYk7q7GISVqWwNwSSbQY09X6VqQJPt77rUt3RddskS3fNUYZaU
vOIDPCMY27aQw1m+KpFwOaoXAYM80hhDTY1eXKSVrCWjSd2ftnETkVRNjE5RdzB8
VBSH2CUdtDXdZPzzDVqJMBYp+fyuRGXoJoGUN2IskopNNjPAwByH/rKp4Rjy19ZS
sNTjJxSn2Qu40QUPO4/+2fIdo6hJnjYSsxEP2Ch+hvHnTfLWPyf0fRfxx9z79Dnh
htvY0cYIY9ZlCgiC3qjVBePxeucYVgyIO4DJU5W8sV6X0uPPoklDFBVQ/sXyRzys
4pZcIcBoBrWvvZaDIEEh/Cq+9Vp2RmTeQLWNA9c+r6DU3ShyGCjRNePVJ6JeFTzC
4JCO9nEDVYXH5WRZdtq3EJ8H5nCwXOPDj9njSyMVhfZoP/Oery6B/oB8D+3ydhWF
n+dI1wqUXSPuwt0pqLzPDAcGZzkXBuHhbRQbdvzRpRFzaZf0UzGJlQEjK2B+pnP5
Sf1fLgSs+EAtFUt5mQ5S/AQcVeFpszLf8FJU84vmYq4Edc+JmupLYEYnol84+WTg
HW/je+GDlzBOeeGJL1S8wj7ej39Hs1IQtD13jNQk8KC26F79wt2kGb++ooHJ8yAa
DHvwL6gDLag+STn/Lze520i7VXojDkBPrNxds2bhQLEbdAtAqYcTpuGhTvOmCiDb
KfuNwANVbZsiS/kiHfcV5wwx4/MxMWfOGCDFxARN48RpcZkp/4KtZERnXTcPkWJ3
k6AmzHrieY6gTrAuOjDqPHwq6gC0vtGhCdKFOETramvF3Oz6yQCq443Qf5Ypd2q+
RJmdcpc3umciLPGzWB3aCJPG057ZWsMKWCmuSiXSRR1ZjyoWWMQ6L+NZh38aoz5Q
pgi442YmeMO6qm/tU/t0u3GRVEUmHAW7VXdv6TJWHTsFvZmDGWeVpfMTcWJkqZlT
F/m4bZVkuvEj37zfAAv7zjaSI1JenxlVRp8mKWpavu0mu9GaEvHXI88rJhP5eMqF
bxwx0sS7bgFSE8wF5WgIzYQfylDjRFNJEppDQpNIfVsBPG8mQMt4SQKert66o4fs
Oc5ereFHF/4k/8XhQ521so461pgVxuzpTGrvvlsnn1QSiWUwWZu1YRL0/+cOi44t
ToLiWq4cicXd8hDeEWNPMNHxZ8evnFlh+kabd1R7gBBj8bq0CC4p2I7RsFx9t7vY
NhN8cfPoKM7/R3DmvEv/mnLFnqk3aSLMfXKMF5v7ZMqhaZWgSB2MbAvnC2BDVBHv
gAZZYsqd4NL3dKV7IbgMEwMGRU4L9JFOr9PqpjxAY1ZalZjUfDNqgQLZc2pnmn5E
c8AueWXibZ6WrZ61pxhow1f5+GuGRKXk/tGV/AWgDN0QIif0h3zqxevmql/NSeIG
y+6wDtCQKy48EJzO9i1EICtUBdS+eohkhwIE3b68KT/SILbaW0ru4keH2hXWizhl
l9cbuVzjHB4sX+3Yiix/WEcHA7lKKlkmqMJBEA22a2f60F75ak8N/vp20vCtE6Pl
0jO8QFuat/E7OD2n0UF1yZi30bDgNkqI6qvMLhCQPo3aqE6h7P+Tog6v/Xx9u7sH
qEfBN4a8DChELXOxaOlfLARDlGXsXqDBeey+fIRK2AJa2D60ttU2ZuoXPNKwwWvh
MbeTsMcK66fTq6pBDmuNSeOa4G2AXE2PNLOORY3b+dvPlIECjkTEVojTgSB9rueT
NRFr6Fu6YA+ham5xTcsOrD9lwZuyULmPz/0RN2ZaRdJm7UKjx6R5dM6r3ETSk7gf
Icmr/whpxjmQySlDtEf/Mohkh9X3O2qsZo8kzegRBgIBO9hDHMOjCp0r4Db1X4LG
lSa01R7RJaUmw63UJEONO4UYPDWN5ajtu/ZEJ/BO7VLXpPLz3GJOxO4LNyWKJHIn
3vr+QPAsyjY/YvYnZqxMwpZ/26LSf6nSPLpkYIrzRKQmlJZCP1iPpDhneOxOWtts
WZpQYT9YzFxpya5AA8QqWhDQD0DEyKO51la/8IJZlVREMvFPcNI6zFv+N9D2A6Tu
iXnBXOWnmUHkApVRfr3ffk/ZcAtf23wj6KSc6ICja0G6nt1d/zqpH55YG9DYca7x
RdeZG4T5iQM06y2LmxwuLLfnmmk6o14bl42zEbnc6ox97x5196t0/Jor2nsHinaZ
F5Qy+bfQp9SxPlQsEYOmc2cyGaeWsfB61ENwl+ksrMyCNx8BMNg2fgFQn8uhhHVP
KJmatFZSZK++PN4d/2BlegmHgD+GjzRoiKQVGbA+k4gkZ0A1wHXG35wWD3tUDjSM
QAGwvJLL+Cfujhkg4mYndqgSd56AjP/WnQaODexqc4vjFFQ6RhW/9GY5nXN38FuO
DjtGAOqY5YF/1zUGGBPDkXWoTKC/QBDIpgLz+z+mxDEq0Totp5gXfmPV3FYVc2no
FkfBZ8+4Oi//irabvuFwOeFylQj7HQzYKqwMte+9IE6tXMd3vIp+exH0ITDHdNn8
ZoXQZ0QkOSrHqE3G7i1g2GabTcjnZj7V0Nu2lZ+7aDOkIM7In8TnfyxcJJAhSGRw
p1Z+uifcbP3k1qiqrdyXFFl7cufaJyr2Do8bQB1xC+pTTJaWwKol8ifqXHOyuT6K
X47cyjjj//TN4VZ8AhGkaJdAeQ3rcf92L6e8sOi92meJo9K+58rgfikH07nZrUH2
dA/lSbP7mYmWF/MHeZmv7oa+TPaoi9GGbPkQC+lpoU4aDHMbbTlmn5EhUieJmPI2
TpYQ4613L73Ksarzfeh0G+M7rPOPHtSsXNWEM6+UMmD6zoTuX9RJsdaB6QzbeswC
x+bcIxr02rk8Om7dj7yawELwdGYXNej8oI5auj9ZAofIY6TXSPSIs9Ua7BEvePvO
P+nlv8rIeZiMb46A3hNUAJ7BSTLsChFxbC2UWU6giRPOEzqgOwswGK2gmE7pqmI7
4OHX0aJ5kCWMxmo+67cMM+b7eaO7neOHhRffJ9edyr8ynbmFbABdGkhlY3jzOpbw
LFS3AAnqHILS4dzDlOlALiaoIn9YX2Gj9UTQMPZ16KQKKIq6NEBoHPORDen0MjhA
21vnQPIjMT3+9VrKjhqsi9p1t0aPxK9uUlVbyLGhOZX/IdO0IcXhSUVU1s5Ksp3c
3xUT556venKlEQZP8sPNGKKwO3kzh/Js596Vi8/ZgFcWVi35xrjzpJJBpfMMNJt0
3WoEg9pqrgNhc/C7bjCbX/1FvRs458cOYISH6c3ZGvrl0zI93mVIzA60MUlh8IdK
eTcPcnUH9SQxVfAm2j3V/sfso4svr6WYQ+7krAyAWU59VNv2/oKHdSZ1YqOQMR/4
l+5Cgoe6DtI2bCldeg3E9WRMDq2FghP4tfEMUyb8+S3/nF9Y8rpRu5e6dJUifUfX
F7XVq+NF7RVOY0Cc/l8oL/ztU2xUeV5GJKVhy71AyP5xmlLffPJKFc5iI9O/9tWw
IdCTWox8uKOU0x4/NUJUjLkcXOxD1M/iRLfEPhPXpFKDufN4rD6iaZovDmfj6iJ1
yj76NJpGYB+v7eSb7qnebluFfAuzbVPHsMLBe02kCr2XvpPXsA6nk63lgrRnqfid
wEGxN1n0Q/vmTZIJE5l+gP3PpJ+u2q/pgnu6Dm7MPo+eEFYYNOgbkr4az46Iga/S
K5J1dECB1PpC+zp9MlZALH3Vo8Dn3allxcEYXp41A73hUvXDun+GPPFRJfghFXIf
9xUGadTQ6G/KJ5feFgPNTpbdAHNrSG6qrnbP5IULW80OhXIj1G4P5Ukx83ExgS5m
6Q6yuAOPytROnlfBE37o0nE3EvdVFNhkUn6OLltZhCH/vg91aEuSQFnoYFM3AIWQ
d4smeQAqeQCjCsrSPrRGzq869gDzGQwNgA5GvRu3qdRVvySvq5X/rL09jZnh+R9q
G3n+8B9dbo3fneVxOuzBTcmn54Ecv2qDhE8beRSwso76D9U6CW5/AZqZcb4/D+bb
jw/A1C3BYYAqqnZj7EV0dwj0TXeo8Q/L/90JPV2aZqw8LqabNlcblg3/WQ0LvcU8
ZsUbPCdjH0r1uSakL/VWPhH8AMhJJODvn/BVVV9Vd2WORM6T9/A1hZaY6Dfi36gV
ImpIo4LwyaEMy5HMW4RGQi8B8JaGDlBO8EkzlnbOzjyEHr4ySLUeYpjAYG5oMjIw
97tLp5Ks0nwuA6Dt86dVregH5e05uWoznFzQAlmn5mU0Mm0RzCCaKj9/qAhoK8BC
cKZiuV/o7BjKMwE6qcSquT23onRMDkPL55rfCx53xfGB7hqiQn8J0W2MbEpRP0A2
OODW9vPVD5qGYfjxFTHEpi6MDvHXtKpjeJFHrhClaldoP5WcLwPgK01hTt4MGMqB
CGfm+9EKeGc5MpFqrPtETcbfDsjn14TCi2MBnagHU2dQfSxOAReTaQVvoPsE58EV
1593vWKgo5tFxgiZb2xVg9/iM9MMffjUYO1Dy/201lIOEe1MBHht8KSNXlFeiES/
glKn32Gm1QrgsaTbLBBK0KtulVirNS1+oGur9X0yAUbiuxe9CANl576o8iZLpnwn
EyzIydEtVYCsKbAqLA0WgNz3WcoaDGPL6Kug01t7VEBTrMatBU0fexAMORGWXozR
DF8wDTaIqz1PghNKT7LFOyk1KumHhHjMQbsFXiAvT/OjumbuS4ag/VUZiqfLXLhn
mUsGzF9QUFtzKk+z14qyd2oNUjRyYqR/49uslyMDYlB4nscPjRcGzyS8ZUiNckXm
ReLkN5qt6Cy2TbRPkwKHVxIjM14t2bKffqJLh6NeLwr+AHpG1QdJRZIbJV3mTLVP
rF7pqCOIOZXVk0qpAh89yVskGuKq2Vw6tBetSXQ8XU6JQlw3DxNmzy6ZhccSCOzD
np1G6iXlaxJGz6ZKLo6Qjs7Of5LBZT4GdnmQ2lBsEWZhzdxgr+IZYArin+RxJUAJ
55dpaToL7TklcE+dxIhrEPD1gpgLNsMUojXzXu6S3MuT0YsYErmVCgzi/ROstlg6
RELY/VnV+C/poZY9S3aLb6ftkCjHFsTfa0TzX/cRQ30YzHmpEPZdsKfwHfAGMudC
YouZ0j4LZQExuy/Sdv6TjYmetdP8wQ5574RL8mmkRjfYJD+i8e9eGDxBxv7oXZFd
Gn+uvOotwn6ODwsaKFGzjvm656dz6CCrgZ280CvzN+T1Sh5V30LJQoQs2DeQnL0i
iuFS5VIQMFXEhFkTp+1Q9W+CAUbGv7PomsTR+v74vPdk4Bhq1XgcR50NAi3FWt1N
SZLIwZ450Q8qX/3xU1Xn69jb0ywwxKLrSk+qO9suOJBOFmN6s13Pu6p+E2F4Zcbv
S6CxuKduZcmorfh2H5e8xou9bUc8U/K9OZfE5Ycj0Rou1IgSzR3Y74aQZwxJNkJw
Xi5IPQ+kbcm116CJKI9J487kz0PKylUhsMKzlibY6MMyUErNYzHMLQFJr+R+HTyR
B1Gx+Y9qBeRMnIWf0yCtNfSffI/LgZcYGt0qTAtvKi+f5iwl0yfexC1Rm3J2TiJn
ZlfDCz0sUs9iksIzPvEGgBsPxQORou+pA8KEP5bouRVCyRHCOfBWuqJLvEuhhHnn
3DjxH4kFw+cUOujZMpMl8XtnsaWIpjPEE+6DaLlGsAHw0LW9dPowohBWxv1akYIV
RapBBpKZS8K8ZiQA2/919fNRSZZatV9bn3HD16sKz0qWw2a/ZOontsPTcHDn6o97
ctRxzsYRqIV9xeFvd545VO9gh3PUdx8HFu1dkntnYJUvGKPqXxt/T5vs8DZDIwCr
+Lk3XA+Rr/8hVSXBB9cDCfpYPUi8J0ieRH8/F0KnApIMeRsmzvCjpEp0LPl40/TP
N7/T0Lqp9ZsnsN7pJ/w7JE91UxppEAQJ2updQqDey6IvqOlz+Ev/YyvfFrvFAvkQ
IRS8dozUTIYBQsNDhMS3XOeFvq6mTYiVQadz4rmcz2cVp0b94Ks/rbXcu0o/8bih
DgSfVjaWME+6GZfnHo8pVCmDKr0n0xYFApnaD2/6jI176NWiLMatrKoZqfHNBi58
WV84Yxn8BF6HSwVesZ02oH0YM/TSkBJB1mKvNkXLTZ9qCvO6u27UMKC2qbROD9H4
pz9cdQZocpv1A8WWlgZ7LxrV8olCgNpQdEix1agZ471rBGSIhuXAy4UBJQhrBHjS
95wZaO4/wNektQcap/aj8YOMNPJAl5NWd58f0Kg1tLwwPrN/MaYm3jUpZaKnXZaW
Xf/cLFsvqZcbk+VUHkND7LMn46zt3VdhGYzwvBj3pjR/5V8+yFOpDU/ZwhaT09YF
oO5USiHqqzl9VqjhCsX7l8+p3ZNQCPog89YQO65IVeSU6NUkRBy9lNU05Jqi2JD4
ItHvNQAA2i7Gb+sx1e0LHFGcIOtRQgBNstn5acG7xy1KwjxiMV0Ag3H7PHqxK7Bp
WhlHc5E0IiwEPa4WZVzanLYMDQEQwLqdH1CMTBno9IhfPlD1ijHEuK7D3FPL9vDl
mdj8COzhH+6S/Z1JKTH/Y/UJkbMYb9M7z2TYATJGCePC8JXqHOPE4NGWj2v5eSmb
o84ZPozJ33HWwVIIw9nkB6/eRACt+1INJOv87QCR4MQeCLOYWpurp5bHWsILpW18
5j/zA1c/mB9jhb/3XAuPT9Cd4u2pCEbSj/It+Pn751acX7gBkGkkXw8BLSrukOWN
k/3e4artPk1EHSVG9GnWzkfBKs880nIMsa1JTEzQeD513BngJuvpqCq8/XTzH9pS
xDnBjpEa17GYQpay2MmgXGiQBrqkIhyHQSFMb5P1NfpW8+pLRLxwdzFNDcERP5Tc
2KZp3sweCKA9K39Efu8gPr1AOze7EwqyGVqMqhozjVy5fa2VWUhRGICTf8hTp3Q5
ieY9D0haMehFxc+PIUwN46A1qEXJxWOBkCewLThMeTbPX+Zo1IO6tMX0u9MbOZGO
c7HayDPTV3UOkI3Bw0zKMcutof0NqoxgVLnBWSsA40gdsTkDPzo8LqIdz98Z9f+9
zX41DgZ2z7wg/tsDe9bZjF5qb7/ErlEePJ2f7mOEsawSWGxDizg/WGrST3wcV8jP
A46hPwlJAaMaPw/fJLDgomipkSHX9R2cY/eZ9WM97hS3OHPAXj+Af2NmaStXsWUa
mgPz3885HaB3joZkD/dzVrlRDSQgMMrFCDmcHNRVeR280H1Ol7HJiTB4lM05N/4w
LPlykJEZyWYBPeUvnq5Xd4+n/tpUJ4BukmgqDN/FR09M+Meftqaby32JmKhdI+Qk
vVErNdApPoaJKuy3kxS0n+XHwR6q3t8DS5U3MjfuPFinzc1Jq7VbhJJtwU7ByGHm
SyjFQ8/e55jMdICiOF4vC+/RaCrCIeNuh1e4Isxkd/0tq+lmdnyY7+5kN1VZ7HX0
ye/o2hH/PsmrwqE3FCxXxmNMrBjXA+uR6Fj5NPFifW8H+20JDp7FCPgq4hM6gCuR
g1dut0IxCS1Y1U9c3uWfCYzvQsbZxoTeQVP+kavl9YMvQX68pPDjQbzhMy2THBQM
zK7/OD03bW0GknHsX4kfhGm2Iwx1z2/R4+PLH9qrm9qvuRncNFjes5Uf3IkZW1j4
bR6asw4yb+WCSIEUSSnT1CScfXBx6erQnxhsmwdN9uDEKFYCatnpQdK7nKyxjv7+
ZSkm3ou4UhU0z+TmMnzxLpO6VugyT7TbMX0uX7/UOMYFkDk3Iwf6S9SvDebO5Yl9
YtlU8UKmNVuw+jsGLsPnCYq/AeRldC5oK1wfUG291e4TzCKlN/K2tUburNTp5TaY
/dj9O4JpCjBMLXtokytlMeOflFo13oTPJAgxs+S9LXX7EveRK/NUnRDUDFEMD+3y
m/8tYDiixPoTOFd7tvTtQu4oCYMwVUCJ64rMNWrBNQbpERBbWitzGforn6wby+42
IQ7uilut+44hUn6gU5kwxs41b7qRY5mpyi01ft+IfNlOoYiokf/3Yj/sAYxfbJ0b
mmnYXk6PD7Liqu0UjRL0xFZNzgGrpuobnP4LKRGtxBDClhl/bC9gAmXhjjP/+jZc
MU6+5SVDkny61+pZKMjZtShvRWgjtHRiybthAIzXu4eFgUzhg0q4LDRv0AQNGGNU
SEIH8yahzJgUSJ9SW9r1a82tGLlDaUg8L5jZSrvrvbF0Giqf6aI1Z3hX6yywi6vq
5oeCPU1eW0mNPQBeSjx1zJwJ6mvyfsnytgmV8dXS3P8Eq4XfVLIGyGn8eYawqB/k
oGbsLu7atEhcjEHvu3zb8dtZAVdvxS67tfuX0UE1AzE0aLfa1bJxDjdLQw71LC3A
xQGh8xrOHunAGgaggFMfQEuRHDVHqeT4twPB/PkqdF+hgPCcDYXK22jb0CUJTwdn
F4fBhc9rytKM0dwYxb+HxLQXEbnQ3OqQx4gH/5g/evx7hXDnbHAmqcEEUwHVAqQ7
8u4myy0sNAyp1PBH/NGNdbsPvI2qIuKxn+zkVr6gsSpJJJy4uauWJ7Z+TXLqNo+S
Vj/433ssyUuyQEHYUVsQ/NsGyqMDTLr3R0TdLni+fS1+pLIFNiusIfcGqz7yt64T
hBhdDDOEj8cfBV7rS0QQEA1Dgu8koI21FXB+ILv00ovWRldCS5Gap9oWW9n86Fbt
xpSSzA4dIzXUixhWUIICQS94KfblSil8WnrLuwu1HIdNKR7JgQxuFvgdaMEn6B/Z
sEp3O6kClZAy4Zjw2akYle9UVViuDHa9i2Qg5jL7NOxt1Nsj+s57U4CPAwa//70R
Fn9WlRR4V8e3h85Th/q4qUhRGwnf3KJsajvOZpgtkD8UU9h3QUXmwplJrCX2XObZ
8Mgamc9bwmcykQZhJ1gqzJm7Wvz/qhMjChniWjkSLn4ibOi+L5HaL9WXdUUHiW+J
eko3meUJcvjRtKDm+uilVy8kdQgTzBuR1l4H10zQI2nbupKSbVAdeDDPj7xmUUD9
RRka+rJP9NqFecVv9q9j4DmZYXdfzJA6IeZBCSeGtuofJ7YrZC+llcfU/jLRn+rl
n1eK5zNK6sAgtDS2B5lq2qfSe4x1z0fLhfMgYhZrKVT0IzgGh/xQra7Pdl6quubm
mXSqVjRKgJtmnvO0hRMVcrF9tCujxFuMJzfCTR8qkYfAI34fWKo5NlVAn0jYpylZ
sctfdpKfPWWs6Ea5vgh59KKKhbGNVhXfsU4ToV6FAiT21sxMbOVt0qSvDqx/vJn3
KNyIZABADOZiIifKWHD7VJ2sMfNZ4NaHJDhps1Z1Jo5A+LMcpX2hWZPsEfrWj4cE
jX/wfObEGYAJdAmc9TvvKU+hdqROQioQET+dQZ9v0oa9TxNJCC+dXpwObaK2fiDZ
PF/KXsPbVfnCzpbbYKyc9rZQKhixsNub7VUS0FRzZkk0srsznn7O2L3ratT4hM3t
+aa7oxTo+wd4PrGt66Pi4IHPDNjQlYzqTTJkaYIPeHllqlLEkjN77hdIPGMMoxAP
LtrpKZmkgnI3PXLi42ICZpFVrrkPHz7wxnZIOcjyXvBrh1E0mphl+V1opHmumPHj
AVVq/RrWMr2WL26yy/ROcURvf8g2Jf8dbWvJkCFdVq+iydTu2aIyRX4rFcbPEi0k
aq/MmHdJuIx4Gf6Z2aQKdNtOHbdrAtZOGY7wwR4CFIcwWzfujKoc3rugUTDuF81A
yK0QEKb17hHmkAlbBVzVipbHI2Evxv+Uxl6Npg64NlUbzVi/Sp2Ig3VRZ3LCZQpU
viayVjrsHqxKhbp9f/48UX3Hi9cnHwvpZ5W8vS9YEvMRtpzNV/3V7bA0DQ7I+JH5
OQyrzXgWMvTi3GEg5GZ/Ppr/MjTkyDqjPwm+eQql7cHGhzlfxTgEUKTHOXAtEZzi
s5wfdYhRrO360d5r85DDXUY7Q/RfNYgLybmAECwDDJN1YtpAtS2DupZkBQboUASX
FXbkW3cCRcNWxVVY4/Vg4GAU+ZgtiaX7I7W4SzF2rneRLAcaKtFPkr4FRApsYMqS
mV7WSJwyZuyWvh1C4o/RCU3GxwGOD81vayiOYdp5E/LRmbDVCLWEYM62LuqTAwEX
R8dOUdxWx2RS22iVyfItyenlDYQAZuUn18gBaC3+3ts/hp3Ra/TLOqLttwdPxXT+
iabiIKtuhpztL98uCqMV0rVepjIYycLOGX4j+dNz0zQLIcI+M/haS3GyaG9lnDf2
vbvgVNnppJd6tiiURuOJkHacBwbupO5kHSqncJumsLTLiVteWAKAI6of7ygfllCl
qSlUPSEQ+RygDqdvbaKzqXcQkcs4kqs/CKJb+tSOpBGddOB7jidA6YtfvkV7vjuO
MtLeI9JxKctY40/INjD0Wawx/qxPsN+0egihodObEwi84xq6Lf6hdLHAAVAbt4V2
ZeEkvdmbpNW4UpHBMLJA8LW4xZwfS9FsSZXifbbCg6lEdJtYcXKVBUO7fX4LU2Wz
6SwNEQ6Nf6h5Vi2PL0xQH8VOzPMtSI87pUIIue1/yAIYAi2p2sxVYB0SxOReIl+0
BAAMReFVmmbsuSUpNY2EO7D1lbhG0ka1SUM+MtihvPpBHwqYstKzMzV5mZ1hGa25
CPoJoQ3Cj7W5nwmntzbZZYanBr7i6WsSxFlQ+c9D/EKysJApNNMLGMPjuUncLcRB
kPL9kNtjueMUesU1aMnm146JLLZGmJN0C9zdsDPR+lGd2pgg/UyDzuek5H9Jn2ht
o33rw1Z1VPPs9dWtezjU2WqPiG9US7eXNijjuENdQqcvp/2ZesmRWESW+zQrH/1X
CBXu9bzXndFTDHQB6l8VAzModn6VSBuUVyXC96aFnHecfTXG4WFHOhObDgV8znpC
/XeSbtKeixBZS2eH0Vk+86GRFMxgPH7WIh/a8z3FXTwc/FmhHcUObqX28xgLF3zz
yEzturoLSeyftpj7sF8S/wM0+z+8RN2eOdhTbgvEYeExi7FHP/nkMGrE/tWHF9Xe
i4M1N7ZQHHjnIIsXK6E2uT+gfzfD4FTn7UmC0fAXB5PSGVe8pkwyv/9xqLA7CZ91
VwaGWzr4DzeN42ZiSxfLBdT2KvDFTELhgmoSnzDQEsac+aD7LruD7mytdqty+SOa
lhzxWF4EG8xAYp6ZFTFGw8ViXyLXj9MoC+T9SEWbfIIAmbUFpU5PPB5fcalyDl3d
6z7+2GIV0DD2M4bgmO3ThutaKgQBxb3gbuafZ3v23d7ZTMUmwdK9I5hidphjBhDz
lI5H69rnJazZIVNPONOs4mFgR1a/MD8UrX0qU2pFoUeLP4kEywTjg28RUHo7eqKk
LpHKXshZh81Ss2JGikKq1hYLoUiWYD7z7Yb74Vj4L1uW1kD+iQycmQkv9HyJQ1AV
b8TPD4Z6e/EyPow6OrC8U09J5SFYRR8gkIUzoGBIJp93CDCZoTZM1Cg0CstbxvW2
lUypHCNDxPdNUEKnAgOScUkBrdRa0MqWOaBCkawgNqQ5UvjxpJ/Ns0Q1n4g1d22V
gB++ATCp8n59aJuOvri2l/X7TK/0r2XLaBR37tK0UZdVwuVG++zYQ2PG/ravkx8d
uV6SWwmTWADE7YcDn3x5mGaGtFK+10h8cJU86U9p6TGHvmoeFXHbVQcYBw5lvoaf
91rc++HZfKHqb7EnlbHGhZgOEkx+GK6Y5Xz0pxFYxU6vm1GHLcuRZ7GytEbqyz1U
yiTlwRocsAVJi5vYtvCX9XJIjiBlLOihS69E/XCiblECM6xwnzVvrHqCwyy51gs2
SSKpXACa+eo0g/W7yT+1n1pi5XsYH6M9KpFg6O3Zen+h9Lc9p/y0+8v6VuoUX+Xo
zEIAzReygQZB+1ngWjoRI6ui7jZspt+Wgiy8rxHyjjfs4apuGsphNuOYhuCq0xla
noNkdqk52eKVhBva4qshA6NPOvKb3+Ca/42jugxOpn2lZHjW4Qi6NPf7C76xqRD7
tL458Ca98ug01tJECO152/aUNjnatE9oa05jMhLC5o//e1WDoZNvSYKKvtLcCa83
p/5iNTA1zYo5l9I19AaDZ8uP2Yvme7oJPM3NkEl9cG+4+DW/sJQw9B/taT7QOKQC
zgKyh7BYuOVVYv+aF847s7QVg5W7hA5TqO9Ys5Tq0SCdqGaVT5muYnjj1UEon9kW
AxThQzsstnVhQyljiSwIftaELkFBozZU/5OJdTlY+ILbup5OBBk6gGAd7SFItuCW
DqUTJegcIORWerf/aEqloIReZSOs29N6EQJ7rtH95TCfZSSsNUHeICDfhC5aVdv1
JXiwZTy8WJx+2pltw3OTu9XebEdYfX7mMIOa3aJ3QqqOf7nYnV1SnQ6i5wF4KcNG
a93/o/j424HZW2uXaFImZ6lHDbrdoSIoamR/ldXPnZIcTRAJunlVhpGa4la42HVq
vCYxza9c3GZgHCMoBk+74lE3rIMh5Y+hcDJ6EgOnwvvZvP8WpNReP3IcjB+/XX5T
gJX4iOsCSG0LZ1vWG9nKAcqKcbeuBn9dpR09JiTLA7dG7nTpAZccN+WpSG12GmU0
4bVGSMtBQHSe+oAF2t+bLcjLKm59s1T05wsjzDkYYmke/b8qhgg2Hco6TlqDs5Xr
WvqUz9FhnZt39Q7vOgbO5Da55/y63dUCH5Z/IFS2KQn6tgXA8mFab1rZj7PtDEOR
hZjbkKw/exNimDsoqQgDq5hhhB6fmdx90SKYxUA0qJ9YEorQ/fr2cjmFIZeu5uJ4
ZbhB0toicGUtvh/vKnprpsMenJfz4aevs6vnrEfPRX/uVQal0HbQz/gkR5aIdqPt
C/jonbL+LpmhJlsUOWOnt5xQ4CeSyZXUnqc69WVAxy5x98ryHRUw1kJJiaWyg95b
PF3F2sPzn9YrdqPhrgtPPskAn5FuUtPyIAzWmAzBIHZJZ9EU8OWojPPF9iif5C2V
4eCqE0R2/6U5DqTwjJrSVKnHeA+68kp/KMKZPw6QE+M4HOv2mailI857eSzFLUDF
kitBHopgAfd0YBKzPtoF7+8ZbC75A6cOb4q4Ka4jHxQh2euTEILM3WILuefHF+Fc
3oGwzIFpuBZlaB4iMOy5flRT/zrMLuGDUiKuIwjyD2wppUKl3bvnhvrg6aVw8Dy6
thhybpmON2kK4x8PnMppqjv0bFry0dxpDFbD4kJ3YWz5ThupYB9iqNwJYHcMnEu5
wSBl4WuqMne9U/Fy9/jMrvZCddE3Hm5IG8fqJG4Bn6vmmSaviOPttIp9yaLGahIS
BviUWiKYeiW/3Rx09u51OAiQ/vsCGQFgx6XP6D5S9gB7oM8YVkPw64Aqp0zywk/f
+/eemptm+hoTMcEovYXGIWXMI3ISmLp6vLebBkYcorgSAcGVBACfNkGcpqOAAmgT
hBCQ15KOAcwx21iKS5k06dxPKR4zxAhEqk8m4GMFoOKqiA+0Ah9j0pBh6Ww4+md+
7GA1/2ljXa8HM8mi6Byd7KZ/7Gci3AJb49sg7GS0fWTExVl+ZfQHN7ECHR3PM0xJ
q+cbBAlUQJVRknWKfevBzINvCMrtqXbWmVuNTRmEAnVtavI/SzjKbgyFJB69huKG
GD4zmQ39LiT4ktU+3sxyDqkf6gJBtw9x5Bhnvfrz9NO+989TsjiSAA+PpjzmBQu7
DhICgvL/zYswzchOulLRWbgtBCP8aU1LYbsowUyQFHgh2k7h9ncPFdwZM2KDck+I
xWMEj6D0XIGfqaeTN1cgiRZidD0JfE53At+NV19jB3masQho++eG4Dw+1DETX3aG
854VF/RPlm4YTbv7IxOwht8pohTGe39NHaP60W0wkke9zcqaWZcXUaiy8OcEEOjn
BttDDcj3EctkkHvqayrK7bJJyD08Ixp9w0asPQAHK04TmwYFt3d1TE3Uc4Yi6QcR
1XsXqKt0PJWue7GY/hbl4amRsG3d71G6zCsSt5H6ElYQOF6i/obwBPf1dOCvkxyD
NZNmGBSixl8kE4n73ZuFpU256obe6n5rNTLDTyvezzWlu9wBjznr8J03CzgOcK4N
Oei6t+LfG6GvjvlyE04Fyh6/863YtwjQkt2zb4x8FXdgRU8aRCCfykoQhgVItHfN
SUI49W+X6/SjtrJnwahEKE6mhK9DOVcpTrJm9+hfIbyrUqXLlAtDBqB2c+Lxlcc9
/Uj3/9pnPgST7iiwZTAgHgY+2Fo5th0X0nTL/kIJOixBstUq/9RvVWXIeVaya1Fm
AK2soIuxTa3dCXpjjhMIHLRQcC7lcieMHS34sk2oUIwimOK70Yab7I5KwTOVmSPX
sPh1NkKrW+YLNS3LLLHp8kkTST0lT8zFZGvqrlgXQO+jE2rpUpPxnITK60dpGJo7
3vxG5obZDrM0+gIqbqp2KMfuNwcOMPSZPvbq1FXkB7fvFl5urRxwR0C6x43qDZ8r
DtviMpvkZOnllxr2tO5dA0Q+Sb84G8ejUBXifeyhxtSh3dSV8tPLp6ThN7dEPp6A
LuwqStSHDTDGMrdI5lnux7Sntv/3inDUd9MAG15QGdmYOSE7fUFJAqVM40Cg/c5K
z6vpan4PZesawJTF+5TXnbiVUaybIvK6jNEXNbxfVXFaWOAFZYOIpBwPW+UunMj6
8IZYv6wZZ6mvdtiqPDNkSYufj77dcJVG7GcFYKYc3exr0y+fley2shOXDOAlZ58c
hhn2fjoZc4qRxldWsk4vnyTyXYBC+r/Mg3rUXi43JspVaqt8QXyS4w5088tGQtSU
ObHsglTPVGZrQ2g+XHOsOO0Tvv6dIQtI0bfwtjFIqjBe7DeyvVmrVc/hp4GqyPsQ
iE0EaKs9X2Hqp/PZX4dTmaC7Lp3WvpAj8/QQ/YbL+nGeNgsyMLH0nvkOH378xvA1
Kazyv1b4hIXrQBgPl893FadygyVSdj81cFrHiAHAMA1ZqDzHsSs3+wte8oRtEEg2
re8z0f1E42VclIZuy0kAO1ECgQe/xUVBqAY661F1YLeCIeOqxWX8PpDVRMsqcHeX
28B/c4PhFCjTPTfaHbQxvEZn8fapL2oC30Yue0icl0Pr6sWJsstK6AFYmzVABmPW
LHA2f4PHHP0dn0XssFrIcz10Sl5JNJIn2hwduA1yM4LSaT++DiYlbzFGV7i1lPBb
ph7F9THCLpsfln05VesnpJcbHhUV7L4QRv1Ns8+WtzyPQ29qSjZQ0RiO5PyrNwbg
wu3XZxy3wjwmc0dKMzSvzgwElLJBpCa2muPLmqEGmULnHbtKF8esWDqMn9a34WyA
r+fC+0MKHLKrED2tbXubTUkkw0ePGj+Fxq7+Sz9SwiDd6h79Lhostqz+y0S8SP0/
eOLVNOQ6EZlctXkp90mHB4OR527su4sP1bO2AmgDpgkLocu/2tgzisCDsWI8Z781
eJ6F1Zf+cIyjuo+VX6exqzfjTIzf2HX2GjUZFZyD2qGBlDiOHrhLrh5ep0vLB/Yl
gJmnqzlyV0IJeD3uMvlWt7QC2j/b6FghvZqWk9zcpdKAySHzEcu5VBiAR84RQzYC
FQ/xdin58T0Mxv/iOANHKA9kcmlwKyE47Kd3jqm/j2DgBRrZYuHYv+ZuvjRmK7Pz
Q9q7Ypx4b77sGYGTUc21bT7cAsyglJBRZOQ59RuTd0g9nm6H6mHTaijNqvID48kV
0Rd7dL/UT5HJn0GfuyvmhZ17RGgHttNJCv6h3i3RuFopQNLo51mfxmJvgmJ3cBPR
BMvdyMcq3HrHgxWbVx5Iea3ieCW90uyozgPwUYotEtxQloj3ZyLoOiDby+s9jCTG
kokge+PIxmJZ35d2C53j1ZhFALUYDHuiCl1VxvFtIwN2bNuK9FyY4oqQ8K6866IH
028cxZUN8O+SXF/g/dXU2frxqepppzFY2O22S2BlL+/65L53DpSh6fQ3i2WLP0sY
fc2jEAkFUNDUZCJJkUovAn+iK6pD4Cgs076nZJSCWoDiphTdhA1qOFg1op5iFvBi
PTaCU6f8pfpKSBXfPTTX86SL+eMT+j2zRw0P2525KK20hvS+tFVRYJ2zOm4msvRh
haEpS3AMxILp1+U9LiIdz84+tF/9NiEorGSYT1KoVqnhtXQYYwY0Gw9KlMhBplnX
J/sGsiI1J9Y/qWd1qtYfJ+B0iNW0OfR+yIc0J4zszJ1qg58Ibj7Jz6flUa2bdg97
9gVC9yhBiVzHbfSTp4z8yb1Pho1q6uVQMrHPQkP+kPci73UA0r+vrdDgU1Ofilve
KO35R61a62hnL5nxOap5E5W8z+yT6ISpTc5fR+S2CvgyY9zkUVfaeq+/sWNGCMNo
AqfH62UaVOZ/QOo4TUj85OrUyWH9CxAtzY2ChSO/rzEhDIi8qaCyJKo7jU2Z8M7K
pAZQ62AAZLgZTO4RLtPo0uB+3eLNdZukHhvOcoZnxnYmIBld65C/FO+AfAfMsYOS
Vv16/pCB0e7U+6NsQjSo9Ektd9BKLhpu3hp3vVSInKhlYkGDe1RG4C5K5O+jTfza
3PlU7wFhWOPtF1XE+ILO1hLcY4v4K5ULY+jLIYeWYjh1LamG3EeX5ryOsnWwoAQd
vFv5uXjekurZMY9fsu+fBsjGVdHtEJUG6fFvuyVcQPdmRN+fphjcE1+opIAcozrh
EC2oJ4Birdjk2da7Z3wKnb8SIocoj1QiRQ4yJrmVZNJF1u4A0luU/708UEc4iK3+
kPFgc+hcWDHpLjwROvtulO7cZfjpNvNPHhxN1544uJLl7cuYp7gDUQBrr60TRkLI
urK2tATLUmlT8tHaqSTUdi7WE/1FgXZQOdN67RVSafyKlBqjcZC3dYeXWVRW2f3q
oCUO/i2wiImHYBHVqjZlr1n28t4ACkQHaM7xf5Ln2pPlMiElzxWgjmsjE4kJtdyV
3znXFoNKMrQUkzkItSdRqFjgJ5FLpSkJav5ehrhLsjSn8k1D22uP6GHwYpOkeVg8
L7JwLK2CjHobZx5u1iru3USUTdDlNEiAaUK2AkPMB19chAXQc2VQXT/z+/hC43LF
9aH+aFKZ4nko81AiCDfP6K+moADF3JIIfiOkY1EqZthJcxxBXw3qyfWTFL7hGgVH
i09VZzj1QAsG0amBGmOtvQlDf75ZIeZG8oVfWAunSWbl50SYecVYrWlnds7dv21E
Hbg0TOprsvLOFjshzyx5TQ93NsnnMKGmODKW45qnkE9aMltwn6+wieZRUmVOAwR+
EuMx9d6AMXs5sZCH+9IuHKohsdn5yFCpYS5quR62+IptP2Mdy83EJxx5hb9jFAf+
KLmBDMteTqCX4A1oYFSMiTonGbYc9Y6zDJPxm2YiYiMh7qv3x1+ZaopkW2hm7I86
guJqnSfDUNgBM3yQDK0fTEpgi2hYsuWRoGzsXClNUQR0YhJrePtGiaXWZMK7Q1TC
29KpNPAVNqIbS8hPgtODHsjamopyDaUh+edfwnR7E37qJTvsVgnx+4jNExH+7xAR
sFgDT/TUnapHMr40tw1Fh2pNjc39KYKx9/7WrHlnyCZa8RLM5pl9kffQ5Ry++VV9
BhvsWnc9wj4ry10adm3ufPsqmGZQ/jjSNcbto44iK7+kcSi3bULfLHDeHoN7228a
b1/4glM/rgDhjOuWXnkPXj5E5THYQsxskkd3D+F6D0mlSgZqC9yKyqVgEeybc9Ti
kVEfyYq8x2+tqYIkklBL7/0Ex+OfT28/XEYB2LgK19wrbpeycItjjrNkXAB52rX5
827Sxjepn/5lAD2uJgMfPOWBsShO7qiSPaP6bfwRSMj+vXzlNoChjOU3F8R4L1VI
i9DBn6/OJUVg+nzDuY570/447bxmIWyXipmF7FOCuwSx/jKYHW32+NUIMjkWu5t5
gx4fQwGrrFfw4lRHHdqQ9AgirxZHdZc5yGwSBiGhKdTAit7B1SKYX6ei0Iy2wIbb
yXp3UGxVrXQpQUy31ToY0bky1NqtTedWXg6IuLS2xUKXccA6D5jn+YJOcL/VG+Xz
zNBgU9D/UoX7CTr4BFCNzU3idt0pEgpw0DVnh3iYpj8PoEhBIu2beFXogT47gCf9
xXOkJAO3xVnnJsily0iulwh9AsRuNHQ05aRc3+TjpRlu4YFi22Z9K41G8PvkuYMO
z/WVoCTrx2FEPbqVEfGKANDsmGgbxa4R+NLzSo1GhzSEgVaJmD9gucyonF0Y+w4B
K3RBdpWTgytR7eBXbSMKjTyrR4jtGfRavyafIdsHMoR0uf47suPd6Sz6ys56aEkx
AkFkQVcWEmpzuV2iIRNzc5fMTgNOL0oLy5xNWcY3pCfDrf5HXjt7LSrk2EHAQNhD
BTbUbJJY7J7E8vfJaYAhie2N7ziGFVlVH+CJcuRI/fF1Mx+m/Xd/6QnbtNYUECHB
lfWpAD5FlOraPhlak/a1/DMSUrzvreS5tlLp/ly1dwb/ZTB+7MezF8oh+rJgD7tY
ychzr5XVy8hsutPQeI/Co+gBQoMSuo8JjMhVHxOiYhNhZ4ksJPOF8/ZEsG/jKQyl
qJ/8BqQyncEMxWIn3WAc68Oeu8KRFd7NqVNIZplyVvsGUkC5sASWJkWDlCLmPFmV
Agapnu4dIhKapKPpZawp6zsdCMnr91su7uc0IN8FRwv1mF3jpB/tUCeizpCeCihx
QVTU13Q02gpfjZmlPQtqysDtmE4SN9v+8ZtLLqdbwfLCyKShyy1NdQVZU0T9cvbZ
OSXHs3chZrJXw+mGZuRo/lTZ053c9yqR9uG9Mo5XbfUzUnzDFcV/eFOdasc/XPpk
RCJPLnx2i72sJrEmrLkq6AyyR3UKiPpFr5K+WTwGng42CRWpuw437JoRoD/ooTGp
j3LOk0lELr8kNp8jD26suEJxEeOVLviI9auRjGD66st29VaW2kg3IplPEHlJTBx1
tHVAXrzggPXymBV5ga7QdAaTo03XNaHtd+J6v6mZaobnXkNj+Oc/68Qtovwc6f/t
SGDkjC+cqsfrL80mIta1HkM7gkapr3P9QoWfoR8BH/TcvLsyEWNpphdFrwTxOrjL
qBL+Ev9Ma3Rm5CQoAMSfXe+NFet6aAiI+W5lfLPZ99NZvmKOfkfujP6t0puROBsK
wjcQyfEnl3q9xsC2wE6xS+SZQOrKvsHy/Pp69joIzWjPAekf3Hh/Im9KnLpUOiKR
eYa7bTyr4CBGhSwSCFjXTosTWPvquZdqpvVh8O/nQ/Zua5JLd7yrVMuw8TY2MkDs
36WFDiTPkZSJkupsErs/qM0Oc54b52ZI3VN/AFPO5YIz7UktdpyOEpMK51rIWn2e
k20QyDriE5M/Xaz642f19I1+4oChDovVwbgA7QP7Ng0JRnZaJEkGt5qv0BqETtRU
GxKBK5Gs7W19quw4HDOQEMLZhIEX4ZVPkkLrJsFnzt3c5hsX0hmsTyqNSGRLUhO5
Fp8zQS8LdZXk8ZO+7TEy9lGz+obUZFTuIgq3DbILHQ1ZzPczDG/E+gQnkpRUKB5Z
O4W5gpVkr/QiCem2zNyUIXUYhISEvwRZT5TqiDbuzpVjdHKRf6/I/4bkWlVJyXog
98qaarbALoj5JGuwhsbraxHlhFFnPee3tmVnSMgOjXpUn+5H+W/IqdVDXRjujWgy
QBlKGU4h0h0gdk0CdSQQ84GAzySwhq8uTbuR5XEbZStn0dyWU3X4XkFgZ9pNPIm/
BhKFoYC6o5z83U7IGeEdVIptNpTUzyHtqSpbEDqAnGrVDpeENkHFYJgTpkgoc+X8
X73dKUlGyPny22c1MtpSO9qKmI4RSsGUY6OL7+PjxjbXGifx/c2+PV7+LlcCTGd4
OF4yIZtIY73qR4cAFCXr1HoAQsCd+e1ab0NKpVb/Ktf8oP6eLp9l9S6lmUJjmcip
HUSiyOKsu0fDm9NNfx8jDh2yVicaVGJZ3c18mXV4n5hUFGwOjYaiBJOj9JvWnIlY
P/FXgE3W7x3RKnFAFL7S62Ivk7UlDkFMnFgCdx50/HQyRp4DpeCDp9c6OIFl1gk3
aUGdmHmjWZRUmh/hiNg5mbietPpQT1HQdk6XeXBZUrm4JoihVCELnnFfN5baMvsE
R1p6jjzbDXaU/y6UXLGeRyfxFb9gtBBIa0waot5fvJUz5s64g8Ikii/GRYluxWXw
j0OhAvoLvLF65cAgWyQuUcvoTFCIT/T8VoIWFNjKW3VeIsmlUH7TCokJIPt94cnR
l7XK2mppa156gPnKhKu/xXtROxCZGhgfKhL0pSRf0wTnpMu8RDwru0uL1k1mFAi4
yM9ROzxQn3kgFLKTLTsixPOGBfVQDal3DoPEZbnkF9eVP19l0VvMvcWAv48n3hu2
aMxPOYvfe1A+F1x8f1naBLJQd2wI9mLx5lNibi4WjDMKJUbwMu14o3lbWN0sSZ5Y
`protect END_PROTECTED
