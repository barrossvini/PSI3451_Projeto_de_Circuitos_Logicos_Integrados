`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7do6SCVnx0pc2Gwh2Ag/Xbkmy0qb0zqceA/WTXtqLvZkyB2Q+HsZaWyyXjfPapvQ
uRB3g8hPZoS5nYd7/tFTcFYCupQWrCTVxiTn313rGDf2oup7vMCVWPamGK1pAa0u
k0R+axRCyfhl5HT1NhizQFhlA2cxseDVZDlhgjvnkqW8x74WdvObufD+M9wILM5x
/LvY5U6PlevTCjvtKDn5EOmr9XoD9DkqR8P0PRUKWL3sA1BEIrA44mq+OYIz0TIe
CFlHHDRdOH1QuJ9A1AAICQDFEXu3KCoErQdFxBkpobQdbe6QBNfxSprTmN+z5lby
MlAm2aHBtcOkgLNbRjXcfdOB9Wo0SoIOoNXSKEBBXRl9G9tv16zddkPRDcqbUFv+
oYMJ/z1PCgilAYy1uZXI9TIuc8jfbSMtjJgK4LdoEd3dQDBpuTFynGVz6GU0o5ne
wK7UrHfBoe1Qkt8CI1HgtXCnF/vCWfOIQlBCL90CUsI3255ze+kU82fQ4Y/vJCRS
cqPrBHmnM8XcuHEg4we3s/AHPeK7WJB8AVskJdsrWjUXAv1JLlWD+pd8sS6XFSiR
tl4xUaB86Eq4jUCjKzUL/5QmxS81thGaEc/5X9tsaGsjh8riksaZkJCzC6klUfCL
/ag0ij7+gA7vVW4jSvSbjBOSszM5A/7+g1O8NyeFbysWiVS93PfbiddpLtkTHN2+
MK8aTjfuIi4IPZ0ez3CwgWVqp777dCOrhawvXT0tzfpu4beG4pQzPf780clKqkHY
kmamJrhdjPoVlLupGGc7/ssXApb8R3O7mPA+yBi06MMuxDF19Us/byq9+cDGQ4G4
tKQXyU2BfudaGOOvyHhXXQ==
`protect END_PROTECTED
