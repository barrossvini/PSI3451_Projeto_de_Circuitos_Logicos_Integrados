`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lozBqehsOAUHVkDcAErbsF1e6k9wSc3GhSjFlCfc2GpXMV3+r26r1K9o3uTh5lrY
CqPFYXa5u8UiFsS2qaCDFbeALz03Mb1sGHuNVm2Kw34nh8OWpsGNxgr1Dis/HwwT
GJaXOEMYVoawcGwIQTcbkVHf5Nj5D7/TmTTBDVB6UriFXrxuXHradjY6Ak6a8j4S
hwjHsLbjrNB1e2fkuD5SsN7Rtqbf5b2MFsOiS4WN+isZ1/9aOCI9addJ08nvpy44
0snuZUk/OXxBm/2CBmm7DQHaaNSXCBEiWmWY449haru4kovEDUWShqFxiKbpVkAK
x5hd87ihy7hjwWq0gA33KoNsKfJ1ABJrO6sfyXZhEieHCFj+1D76Z0rHqPadSQd8
JnRFXa4ODjvgqbo1Vk5V3eNggux579cAYsmPPFoTdUQsIuyg4SB8NzCDdBxPO32r
Rn7R7f3zEfBvjWYY4C2X2DcHck3MUl7Xy/XWbo+Hlqv+TGt1aLHjqCTZMjJa48eN
3ExMQJWvFgLpDEAKFa2hAtKPWS9vU13Uxi/zDImQt0W8PnqyKznlsDTXbFMqTPmr
Tj825jdvkr62XC3DIX9Dz6BbpFC6aK54LRYhMu+7yAZD01sQ5O4FGYituroowUZ6
cTCSK77Rg/AnAjE8W0PSRd/XyX/dwZH9A8N53mMBgogYdKjjfkvAHFFxwB32nJGr
o502jcs+aqgdc95LhduyqXS79D9HqB++xslmZhTShRILRSUMX5IcYm32XqU4VhCR
bCCVLPXz7x2CpyJNeSKaILXUV/pXluTbNkC/I1sZs9y2LZKj6Cq3KAR9BZk8XXvT
BzFuLXPRqCaqLhhOcDHJN2Y2S1DhD+GD9KJotIjwPK4F00Qa7Dt9qz8j9ma5lP7z
c1aIpWqSut55koIftIA/foLNvYPhRZFDDNq0kVj2HTR+jyR3i6Ofl7xcO/z50Z9r
`protect END_PROTECTED
