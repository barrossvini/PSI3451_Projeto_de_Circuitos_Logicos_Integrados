`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EY8QlZnFjMh7p85ZZ7xChrYj8tnaV4vSHfILQIaIoweRUMlz0l/PqKtjbjmcR8fV
/pSBuVQorUedUwC5muE4Nkm3clHpFmp5jBHa+z7BupLnej+HUHDIRndeEEAnGAhP
1sYQmlqHZ36gqgGg2MnT/GaFh8KThQgtrLPT4WLCbN8HDuicqzHfK52RP8jq9VFz
BMmBq2OLuZgmi0BfjbV00VUFgsqwBm1O3ustrI+rwCy0L++Nvz1cLdLg3ChHLGIF
KmWurXunRwmvVl+VDv3ub1qtoLFCJ5hLTsnSPvUo1BoJ0XUJIsHYcvIENy8YAsV7
gzNx0euOa/8rOziHqzWXGq7G7de34yMOBT/P5NvG6RambXyxygknuIHojZF9vGmJ
J8XeGvbkpZLLK00+SFNVurM6h4VXeDbEP2LOum4c3bhArilS/XevfmumAHXUwpJg
DhgVK+iGkNhsorxxn3T+l95EOOWlimANFT0gvo419X71VThxgdPhem3UfjPqYCTx
hh9FS4fYBVA8anhcc3/JW3ZRYVXt4Dr795uryZQOesAXOKq9qFcQbTSeQin+gwZq
ZcVLGaZPYTrMNpt6khFBJ2WAM4jjYC6tlF5ciine5nfjhi22tEwMvpnVzPtjGx+Y
VQTBcpAoF2q4TcQTZameteOxL+vROP+VWAkc47u6YPpNgWC5SXqILddKrX92zFwY
cIHn65c4wtNYd57CdOv4gOxvWwX1knYDDXnEn5LbwZqlQc6MGaMIZS5QWfva1p/T
R6P8Wp/Hcyb1E3Xd5TK7mwf+8FiOcAoy7nILd1zGjkTNQZhRE99PddRnKtqEE+O0
+2bP/AmE+78+JEDr3dlezRE+lmy8ODX2wNFnUDPUpcqyR4Lk4pZ73kLMc0C2Ondb
xWCoAoCqnX264h7EEaQA4kBE5zkZBBoe4hmayWmuYit580RjnhjFxDlfwQW193qU
xDf0UIXiaijz5ipCQQtLjS0plwCMdby8QrwQ23JVXWPXFvjWU9xOgChluDXCMKv0
bEqJgGCDuFetzRlsqVLr0Flc3qydSZnQKBlZ1KCg7n+MqBz0rf9SYHut22iOkSR6
SqyNX3AXn3mLUBIyyBIIeGU/7bM8A9AzuFZMBpkFrtM3HClR/oX0tLTvF1C8qzbZ
fh19Plb4rEqVdiz0GK6jDTrzaOtWmJ7Sw3Tyk5E4oylmutzyVQqtx7cAh2py6pG5
IQRlN+t/EmnbHNBqwRtkEdA1Ry8FPOUsyqCqqb0pno6+TEGdimbqnTRVsud90hIx
KTGFPjKIMZ6ZcP1IDCUV/t72en6k6usTqHwKdpElwA+I6iudedqiio4SjljgNyz0
ZehOLqaWPsIpibTVFyIA0aJUKv+3Ts/jAUnKZqgKQ4ep3WKCtbIkOUJ9ukAaaOOk
bVWkZQVpeWIbMR7qrCg9w2h9to6yEOJwUmXGyU21p21nfZ/QLy6Pzzxlmavr3OdQ
XdMqvMsO92gudNQfVAkT3sfrPPtWmfALR2Zfv63ki5ASbaEOPv/Vz620pHE9YXNY
rBSJRYQeqneQ0geS3R6sXIlyK0y3xQ3EsfJ8/80+00rkf9ryQb9IsuL9h1gJVgJv
B3bU4M+CHV+pw3uRX55uk0748PrH9r3kvYaGgi7LvhOlwWYCOMbJlszk5ZI4IG6C
pFRxXm8JIF+Ojyqjkby0948sUvZWDUtOHghRYiSuP8AcPbBjJ3N2igQ6Z9ovl6cr
B2DlfG6O27LZkcgvENHhJ+7hoaQAI/EzeUQvs2tRzuClOcrfebzRr7mplvM0ccdR
xdeZm4ZFrsDVgoSuxnWmfVxXQeSFnUGKWKYcY0n3O35F9+Z5m5BHTPB0gM9CJPD4
QnHeiJhU5tpHqvZ7ERYICJELyzOR5bAwPXqod9GmFEBP+gF07Iig1DRzBT8UaJLd
xQbs6oBA8UTg3LjBpoQecCcn09+Gpcurasksed8Fd0EY6Yz/LkcyybJYTI5qEzmC
NM5ig65V3ZNuLWKt3WQStuUh8Va4VBYQLoIJU+gnJ8EyHJj4nbofj0BIqyzhaQe9
SiKLB9HV8w8wf+lQFKwYyxrf0VXQuV/95U6AhI5N0zHtqkbtChfG6A0TP4e4oLkG
ihmamsDB8q2M1eUsLZDHMpDmbc0WSaY25MZrguwws5QQlCm2oTDtp9mWI37+uK9g
NqY1Ei8na/psyYm7FajVQuOvwaXfvXwLbe6Yf9ARcHtL3v4qnl+qkhmvB+UFZfXO
XiDP2Ffz15IaRDKll9Fdz6gL69+CpGkiHFUUPMvrh7qbokDOJ0ilQedOfa6VX1+o
T+QCsfcsc+sVg8EcwX/LD/zrUOiFdIfna3dBL5UV/0e2SOqo7Zh79f93bL1PDJTP
hQWXnUi+FDXHwAl9AHmXkHpT2EUTkOJo4ws+gEFzA1MypWN7wmMXm9hncwZKgouS
SD9laQY2UfWavBQLmgZxWTR6qAtDBeY6Vkah4keMI1sC+mnhpVeIGx24CzYbne5Q
XzVJc5RBCGte3IciQsofUHQ1TrjOHBFa8k7LSbxzmvJxejPcP8aQiJ5zjeWH7qy5
`protect END_PROTECTED
