`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PtDNfcR6IPzgMUxyPHR9472onq4LwVD8j+ejW1kI/Sp54xZrAHfSQVPNO0AlisD9
/TMg0QKVIWpkGH5bHhxUZakwrPdn/xVI4K+4LSwPMJcMarukr6dBvCzfnmnEFLcl
e4kkUijuPA1u9iQapCKx+e/XbBjMt3F2Mq1pl4jYGZl09e/9FFHXxSBqeoeo/Bcm
9lhRcpSfKW08UHZtBZEGM6676RoPA8yL8iLEN3sj5M9VwHqJuqmLLZnMnja9fp0P
wPLNlU8sA3zedX2/JAQj7Dp/vVTmmc0M3/Jex8GAnHC76de7DiuEAgOY0dryDtNC
c2bLbq76rRPU++Muta1H3qWhP5Mvt2C05SGKO/tstzyd9X2SOeiYjsVlPu8Z/iUO
Ty/ACGvTFO8HyFT+Vht0NLjvrpHomDQgYJUKlp5w5jEeCwCyYZwzgM6xHlV8976N
Z957hSsFWmVm5iBg7L4Rb5efkGOOE8Q0XWiuUKzbhUn2MjQVR/eSSxeYuRXVacJb
hcEpnGMiT+7h177m+H5l+iwLvLm9cFDead1kWCV5vg11JlzPf6X7HAMCnWtg22vX
eKHar7RF9yX1RiyzuKQOgVVSOh5o4CkfzXqlqFqyK1GiOrb1C1Ih8uq6r1s6xDzI
MzKaWgc8to2rToOBHqknawo4arEY0ue/2X8UP4EeZSakSiRvv0j1Dt44mvgTxe45
DD3JNmuTxBE52gK1qvXq8tZn+L7NUUnwXymUB0Pm2HSJXgFpRfjDqUWd2qG3VSw/
LWifgUO82JBlshOcF4NrR8ifoTqpSvL7zS/ohijrxEt8lmrvp0GPs9ycqRM5/860
LQPMxjJMeOq7c2Q8cvnqz94s9NjLfmYq0yUdN6CK3qnGVbsz63j2e2MzF7oQjb8q
iXwxIaoRmzqRukDuZ0B2uPdYWgQ2Ftsn8uZbqWv3uLoNERy1cBhZAr7h177ICFQ0
AQWCJ96IXzN7ZKVdNRupDoocNiHSeHieR0kubHQgX1q12QEr3imkw93RW+7OELkb
4n7R82EQadzd3/aJpctvz3gg96HXE+n+j2dGarmkVKo8lKuIdwIfTCzUGjbgHQbC
QTxa0+VuiFcqE4Cvc6tfJMOAgsSxwOTo/8ipzdn4GGWU+SMxtVYveA6rgBeITrcF
WaH+Yx1NSw/5dEptD1jnwjmFt2s0NiByl0CofYeSvL3Wg5XY2gRFm0pKm4sIP61c
PreEHEDC13KznAOCLlDWralZH/DChvaCvG4YxDbJg6Zaqt1u7xaIyNtaSrbU88Fu
1oxDPrYWwwKDUDnNxgzu4pLP3wqnthlUr60Ylx1V5TsMMLeWIJUtex6f01f7h8NX
dNhaipFcBXpZqQdgOMQ/Gl+1n3gUd9obIHOh8rB5YWKsy/C12eNxQhlgcDTeosC/
lhyCDcRM5YTKAofq0J6XDWb+lWSjAodOFnMDO/JsMnQCDgBjOGu8YtathvbkKpTL
AhNuhP1nfN1znpk0F+mpQe55PblcIb30ScxKlaZEE1rr9us+HJnrLNdMESIxNy7N
M5xRwxhhN9V+r4fojxzdg96rr/pJ/3zTv2oJrL3mFxct10h2sb4W1xk9uZPzjt+C
U7P2fKc80x+QvZ7sCZhREw5GreCG9/q+QzrQ268RI3/fKce6BY8ie0jgu6HyqVwV
kikzJMFnVxuoMdInk91c6s1bYNUwMqxe0afDl66786FOe0ePOgozQhRtTNwymM8/
PGGuYibss0X5ZOoyKYvJWR5TQPf05uFlH039j0tEImZoPJwFy/jJ+EP8+M9zO0NC
IZQKfYE5lsJ/KAh38UZNpsmFHIJ+j8f3gb4Fmnj684piRW5jOT1mhYES2VD46jjF
WHWc9FuNkXg+3Q2XGbrjSMf2GHjfLHoZjffYUxw2kFqjJ0W7cqjT8/UapdAQeNOx
iBfv70+Gisl5NriL5m3DT3JiLJ1O/Lxqzggl4TfUpizFt2cCBc7903CR5tW/enek
KFjYEPutTQ9triPX71MQyi9CUyZLzv26sS9zHJZlwyeSY7+KMOERB3E2dCO+sHX3
wfrEpHLlpPq6/+HIjQjBFvFd34P6UC0thdLBJR5LMWpqwybIADDxiyYRTkb+dA3e
3xhptgdoyYQMwzrC2CZ/Y5aPDFqYD8HNjOA5obrLKQ5uNpTOCRqk7GY7DSSiAEkQ
UGFfjy3P/S0EBtdtn3o2WFzi0VWTyrSPVDJBgz2ytUIIybpCL3NcRECXDaDrbs1S
sGgQeKhH2lzHe/zlf8YBC4bndH9vp2tP5sHnpL4tVENcyQTA3KKo+1F1aOC6oJe2
1+D14D6LN26+wGI+uWKBBzoTQKqElqjfExFWUxNflHBUONSwhF4CNOAro110DRox
XpwHv/0lIzd1JIUl5JL3G8gWWVlq53/t0bfvjTxNcLEGnlEJ2dFij6SrD8n//fVY
YqzaHd0wqZXaDmoeiAol99LIyCMKyj4cLzXvpCN9lWq+vKBDJKG0JpcCUw189ig/
EqBF07V/7/Xc6pOIslSByNiQszBOMHdP1tNHso/Olh0ThAHJzyaFqc/FT5IAUl0O
O9Q8xuhfeVKxp/fI+Xcnhyu6JnoZ82eUiTDrNLbT3TFALECCTagJFNcKGOduVMa4
x4rpFfK/BwjaYRfnDAfclBbuea9ZDr92DqtBKLB0OxXLla1VnWUi8jn8zw5fYX7J
EEnUkgxOdXWXMJZ18OIrHopvGSE5MvBoRSNZCpX60G37UwD8TmxidBB/A8+H64RA
5Iu9nDjvlOY1ToqBDdbr5OsVof86F+LQsLkrjvOV3D6Z9VTVfdotltydfB3vlvHV
HuEAcsBdQtjdt/aemOovB7c2NlZuaJhKzfscKIT+MQXSLwts7oNf5i8A+hlE2MlT
6PQ8eVRUTne4f2nyZZx5Ahcwa5PZyu2+A2eNmeOK2XVvW7I0g9GXjzEV4RiB9TPy
gQus3SxAm/uzQmLcrBLmUtUhKV8WzKusR8+Mqt37Y3DIbLa0jm6dCcD/8Oq1vqA1
u+qVrGblvTkX7oeTsPvzhu+8QKiNw9q+1YYa7bZjIeuswG4KS3K67Xx0GHjfBvE+
UOQW3L/1WM51poTI/Ev5FQnCA/C7g9ybXb8qSxZQhlAObqCxm+OeICx0+EwF47PQ
LTYls0RFj6Dd5o+mSPl9jviM9RWuLV5+ts0E8JoMJVKvCPVal89WeoJ+/ol+TpA8
jxsL+V35Ya6obj0DRmIWmlJkr8tcQwBRamJhYbANeOr9iNkLyyHjeK02HL4cmRZV
n0+nBVYxTk0+yJu3ps9EWvo8FtOmFqIpXCu2kdqFZhix5zkFX5px9ccF2rXIEqMe
+XCdaO8hvfTigp/3H7rnUqadoqsmB6aSzU4QI7rc6MlBlVBZjx3YfDADdO+IFlva
Ouz4f2nj3gCJjrNucxa9r9wL5ekT3nFNS1qZvy3ZLTzxYG1eqCOlFJzb9Jg4ee61
oX5xr5Q6pr5FwdAZyP8XWIlDtfV+xm6UaeK9/P3qzzt16w4sL1svYy1NTOACT938
g7jQVFXHyMaOa838V92mvqLp7bjOqAN3kFR97cfMURQigw5k61FLfux0UQwuxUMd
o3YCuo7pfltD/6iYhdFiwXDigu5idpKQwEdj/B+7Qo8Etkzx4nMQzs/wIAwedfbv
huVX4wEoWxRBqYfSq99s1eAquy9DKgDdC7eiPoGKtJ3cgMEKovPu/mzfQBOod1DM
2lPS/mwA4OAQHHYCEMX/BmFiUUsVA4iRHSc+qcsltu0lxi8uQ5zTW0C49wNif6lR
XQ5EIl/E5bCI6xgU8a1Zm6WO5VYnJvEglh3aRyYHZ48VUqXAPkM4NP1NeNbeBLjS
kIHS0wT1LicRxcZkd6sr1B4LZiJq5+0VBa6jz13ocAlfvfHIdRIUAwEDNRi0bzEi
1xhqw1vjNqDWa0aRNnH6rMZT2SgdHcDA3aCu4Z010aMHvAQ5pq/QhnBakWZ56sJB
ZmGC36N4OXei25M9XSeWbAsfpRzTNOgpYI18QKa7vsVYrwadEcCpAldkphkPhVZs
TosI2lVdwhwr1a3XZMo9k0FR3/ZIAhxOfAhiKl8Y9pLWJL2x2rg26J2dU5UjBudo
XmhZpubFzkdLPxQIwr9Bn21Ss6iMTLrsH8FNi27Wa0zgoEGn1BCiERnIDvPMASzu
Wdn4zGHOfWYIoA/k4ewL3WZuoKErEG2VlZqUpQFaH1T3hoP0qhyZgGPf7Hz+JLl9
D6C9fJ6yhArMDBFDZ4KP8lXq6Fr4O47cHjucpVevqixfiI6yY3Y6msS4fD+dgTa+
GrhdgJb+JAgrT8CKQHnpxFLd3GGC4EO583r9DEO5xmqrdQqTpSGIsyJA+gGKHKfy
ax1b5rPnoNFw8BP/9+hY67iffma/TK8MJnypr5HHZ6JP0tWgiElmR2ShTH+Iy45F
PUn+o1HeSeEVnYLxnAJP6NNs7/M0MWAPonWBJFUWQ+k/bV1bAP/eA6m+Om8kdcd+
Hjc6xnSyEahOEVGgnDdIxfYTzQHxYjDNSQJGbOuBtUXuKCzMIBGaJs7wqqLGMHDE
UlJVRro+V5t1Nw3a+pqH7FrKQwREc9mSJF2wf3/sbyhqpbQOAcdddElzeNnXP9Jw
L9vgWidEJzkerFxTWhiQxLQiGJr5EsD/A7YEKNxgmKprnGjxQYFJuSd5se1LqHLW
2CnJdfHx5UVqHuz1ec9ETz8Ckvn5jeHw6opTBV3uh9yNWGxgw0q++lsj0bv2hYzO
0fu3CQL6Zer5MAouUp/Kd+4eRilyNlDN7+G6p91iabssroPFYP2EoAWNgeebH0n1
LEt+El+aX/ZMxUIsn2c6bih0uBWtkUV11GVb8ygVPFdtQzOV1ypZrLm5rciOb6f+
1pfODrIkLJq5SwzySF4+u2MrU/2pQkXXX59gqP15H9VG3IgeeQUEICzc/c06KaaJ
NV6WCzk5UigKBMFDQ4VAnifkuZWA8bUKB4WtMJ16cOOhkyC6f6/19Ua38XYF2e0N
/IjEqFll6he+l6hVM7FQuKDOr78xWsEhHFW8qq1UY3MMAjG3mGgwDm8T7MxQeL1V
QpHf171LHplwkfoqrWAs6vZ3uqZugxvqPf99JuxM41Qwo4YQvxVjEI7m9RK0efKt
GlFTqbF6Tt416T3buT3k161gkRS4/apemMnLG3mqM8hJaSfmU+KDTYD691FHCKeU
wNNh9uD71tjfgKbgcukYZp+dXEYWQb4+YuRLPLRBO4QkV2nbOjhZ9XcY9RkqIGpo
CdhEfGOG3scyDwyaeerAzPS/CEOrND5l79v1BSu+dl+ZfLjGrLzZG4gCWhRkEnau
FMVWtCQdOsE0Cnj9Q92fwVJnlcsN4fiwe5Tmb24bloGvHpPSVceNm7mAbda/McSW
XtE9ExC6HnVGmO6d7sn4bSpY3SFBctbpjCKyT8UdZyg7qk+FFawl0eNusdd9PXru
w7P2zjjR3GNUZ9yKwn96+9AKwhHERd93lwSJLUwa5OFeRaeAoimd3SLhjK1z1/Jm
+937wAtrOo22Z3nep9mAECa18Bl1nyRMc8y6nRj3dfMTrXMyPS4hujS/rs3NQOM8
UMSbo1I7Ldj3fjinoQySHpQLNQcDvvXygDZMK+26ZwTh2PJjQi+2odRvkB7sQZzw
hf5CgOyFQQozGa+3Iqna7hxBNIF291T8o7hKzO4FElfNvmjP/XVQyIgVIpnlGAZs
j/9n4CaZpd3/jvV1FnDYFW6MCJPQYcdxz7FT1+DARc8RoUS63BAh0riJC3LUE6hl
DypPJA2K98Xkkx/LNOfHkQ6wC4qiQgqQ6rZ9SzjLvTwUr6YqAq88pMqjoJJM5EFE
g7oJXcpP6OjDRTZyqbHIwnbGQzlxCAhqf72It/WNGw0x4i8fWbaVn55XTmOmJxu7
N5xmjwQDkqKtkSoUgbwdKGPdBqGmiIpSa6fhruMR1P+woNv4/RLofw9rx5XCP/xG
qbEwKYUGlIhCzyqk7SK3Db3ec/tD0vMNwC1p9QT1H0xDJZCkUWpTzeQ+mIxsrCGm
ga8htrSvKfKjzgfPg+iPOy40ucli2hK++eWlrt9lGBDfxP9Q8e6FCp0mUKzuIeZP
K8fuHQ3lFJO3pssTMynUrsXGFrB4S4mvLW4yypf610L8I045mlLMGOR38wsyEDr0
2iZD+yoEUhM20TARWzgB7AJKyEjaR5E1ACQ1P9K6+aWleLy7mV16x5RE1Xn0db3S
DOeTDWBlK0exXu1NyG57jvBhpIzQlli7FvTYxYfPkOGcQqK4Eo3W/mMG5oIl5sPh
hdGmfiOoGqBeNrfXYtykAxBjbEFsd+YhaMcrqfEoHI4tgdLY9jc22aMY0mozvwrn
BR12QT3npQMaI7FIDYxN1qRzprlre6U4w3pPyXR5edSV0IWQYJiUHU3wPxjlE3wM
KNV6BGnNRx3q1ljLSgOiV0Tvrrd9HJjmqLi8pk8bfFFGJBaOawtesL3nU3Xd7W/z
Y1xUrNxlPe1nzWEcuOcQ6yMA1Z6htUHc38AuCz+gj5nS1eOYITDdVuOnSJxQSwqg
5d1fFo6TQEniO1zGHbxkNEjeYoYg1w/SLGOuc9qIiv4wpobGiwiHrHud6Gpdixm1
fK0EaiwkGWHlpX0WVMqsyTjyhslxljc/SmmvMqdQNShYVgtKSvbMFJy45YMg4ov5
5/U9J8BEt/1nkOrNPzyTlUMchPan1UhHTHxn8+35H3LwGCZVztToQAjlfnGR0wQ0
xW4ENWpEjSxVlroeph6rGzQUyt1FPkOREcrZ1xlEdHErxe+Aj0v9zSYN0Nxas/3K
DV1iwIgbimZwK28QfIhc/iHuBvtbEXYZPoQmchsIxtiruN1e/B5bpuY1P3/mPofR
IXtM2WDz6ObuDg3RaLLNySC1vV2lYaqfc+GopSTtzDYCeh7LjAe37KP+5ndakWqH
BemgmA2+oE4tsiS5GwjqB+/gK/rggY/vEJjf5X+/EQiiJqY0dwnxWimfn0kkmXas
j+xrbodq65a78EmJ6i9TZr8Pk42ojKRJsvVYojohR1VFK5YW82HdrHTwMnj1eeej
QZT3NoXp/NW6vNK6XKAU9hjxLem90eXZZ9+WPwIKzy2R32T51qHC6m6du0Q1PFVa
cIZCuHDrkuI2QZjhaHyGN8AgPlROhpwnNwn8hVZnku0ZZp9czLPc4X/osI5O54B+
ED3ReVeWWtgFMzC9v0Nqt83HxZEkrIjRVbw+YCf4ZJBcUv5evYQEZxc/tOb6km8C
7I6n4oiKJVv+HRWAfAThErp3ap6nQk0o39SL7o8QEji2ZBTXUYjHBjKBGQEWZfbG
7Qe7mgDwgZcjD1a2fWmHxIDUx9o7F89ozNUWvBhg4Ph5B8GMFg/r6buQDeq75+Qh
omDKrgtOmMCQLJzM1gjzxSlvrXJzlXHqt5ygT1Uh4Wtyi6p2EjRuS90i1wjJ5sPe
E03lGDx53LM7MiR0f5jGAfK/oGL5sRJaz/OvqST8FIjIHRmoGzEx8PGhasSG7PPz
oG+S6eC9YU0Tcjlo11Xx6Zp7kzg9xXFTaunRRxZjB+H/JRdVBhabvG6ZWOipQzVf
8v5Eis8ueyywoo/KMS/07XF9ATszSIIaSMZqFRNK/TaoADdst4yUUnNPMiTLL83E
F3arSjLc5WyMWBkEJqNI1x83EzmYrbTu7hi6s5PK1QDTXncw79ij4f4BM2HC2sru
XiJSk/HkLNNWPKkNbw4c+1ANEJ+iAfDuYrnurt1UcEiBDpE148BIudY7BLjhgHXG
GZ0BPNLrJ4gln+dTBep7QfJ2Lw7NdnplVNqo/rQ5jAyqetVtytlSpqivzgnRoFxc
0v3/w40UdANNYEwufyQp6lbTtvMn7s3M2bMsWx70qWHbnHb3y8420ELa1KQy4rbe
GuwLti03PdbNLZqS4jkHZHkSkytL/rW71m9Ct22IHBxR115f57GpSlXgbtNr/I5x
4ak8fSTxJ8QdM7+SCMYr8EtBWfMFoHo7ZzR5kBUlAjKYaRJErhJxJEbQdzOshb66
/0xwtTcRWs1rW1EeAFNos9eKlXPWtzb+bf4UpiE9CX23h9Pl9jrMMuVh0VMgOrtj
PyUrTgzEQC5qukjIW+aoRP8MiLOBI8R0mSlp5g2mkR0Nf5lLPwtbF8XRFETH01Ph
gzY5B7ViHefjtVgtfgGe7V7VVEMSm1+vNbzkDIj7eTeRpxVTq2vAzmpKQSEu2zNu
v7LHa36asodSaRYlha/1eRgoKt8f/v64xKaIwqPfPNnkDTB1g5Iew4VM/jDNs2rR
Eaa/5jAqL91nD39RAPgBmTaeQdRh7EjymQu5DL4pFP7fqR3agZrL9ABHiWai+Zu9
gw0dL/+2FXJVO1lusiqbSDFYOSqd8jBJF46IxNDLgaJjSWsjCeF76xBpesMe2GiL
ynM7ejL5ZLTqSxOLwZcv4C76kZVMk49DcuhqlauQV15dZEReqSrcSOlqs/p5fiIo
6aNTyZEJ5sbCTN+A6yjYNgXU8XSXQEDPts9DWvtIy+soRtDWE4HvdKbp7BWA5MML
dHW2TkuCWdcw4FU08f9iJS/1y3uJnYNmxzXrGDkn3E1zTVjpZnzRC5fQkOr+1x8C
UB2rylpZHaxmROIebUKu1T1ZQkh+gnhJn0RzUjoN4xm1BDjstwsZHNPucAJt2V43
E4OXkwyrpGnFaMwb6wuUlB05GiwQgM3aFDShNbng4NyKAcINcf085kdfcU3Nm+oK
QpCQ8mP7BeEKiQydjKKhMxVFiOCNR0dzogFVIize08iMK19iYVHVbxjP67Fpajeb
RRYas+Zo5kZ93PaR6T83/FIdF9St5XUdFBCM9cmY7gZ87gC5zbiMqGGiG6Ex52SJ
IjC24F2OiLtW/iF7ad0pzeAU1oZrlUp/4CiIgQRyP/MoK/wL0TzNitQXWI/i7CKg
uWrWLmDKl89F9wMB+6xVZP6VLgh5M48wWnoKo58gjrMJS6HbgyRyUsIcVuLNyuYB
M0n/KWU13DAeqQQ2SKW3sxfKu9wW1QUZIcb4jA3e79Kfcgc+NRaPtarIQP9MZr/H
LQUpPpAlqHu6rtz8i9oXu2d8GoyspTNXF49P8f/QiXbq5H+mjkWVZk+WC+mCW10x
FYF5aCzL0fGtjt/ACYJiTUdRh7RKCz2rJywXd6QbufvXj/JIlLQQ5aTkXY5JGP4c
GtmjPUQ2ee3me2LzV5xCHJJbixMgOmStMr+q2Qcdb4K6oBf1CiFnqTrM1QMOwJ+p
Wiwrkh5rEOaF6fDU9WH77mm54eR6v82FAEf0ARZhy0gfldEkhRmfx+1oO6pKIhZb
qNL74IvcVPUOIOFiXWCess9JbAJ1IR37kB9dM9wZ3p/ZVyAIu0Obuh3SWEfp/ym+
j/1qtNL7506l7oxtPt47uoOMkAhGmEMtG74QIZodfhKe9lMGvhD8dQmsbVg5Fxce
UghdoSP2fOjkg7O4NYngdGd76qDiC4+tp+IIHrOFAdmabQ/UGIlOE/e/a6YFLOEA
OLnSS3NNwBdtZKDRP5WZZ1rz7adkjX6FkcbgJ1yMDOmFQFtupF0mWuEyNj1bA5yn
OThFEaTTLu2i1ylLzLQGBD2CNzMORosbi9Uc+vFj6cbAAQwK7SyeNLM/AI4+n0JQ
2cI4odcwFo83j2hEuEHr28DdYOmpzkKAzj5kDtxGQQj3kRXz6sARqhKw4BW4nzWO
ExGOUTAat0ntWPYJs3ZuZVhxi8xlobBFowCz/a5ZDmEk9FidiRxl27RqOsW8T2cl
5mYNxh3MwxP/L6AxQ+IdCEEzs0wu3bE9E4xcfW5f/f60ump4ya9aOsIohcBSY6vg
L/0KUDhRBaFZ3osr3IskBrdwZLYAe9uOWolCFE9t0ute0RDIo1HfcljKJD0nc5ko
/g6sNiVWDGNzuR6n2vnJ/6PTyswDwiXm8XBSfbnsLwR7+MZeA0ln7zXGUomNhf6S
GZggJ4VpAvYPjJhAjGwHtQvKEbjpw+k0rvWtxDlRllbSIHHYmVzBmml9k9aj5maE
gYGxm6+KR5xJl0Jbr9K782QFij9gGKTjGgkYdJTICWbZC3CSMw8UFNdg4DleLx0e
gmvAgdYIegwg7vnoIKGWvjaYgBy9Y/3mQpF3hIowbGLnTLEsmIgf7OJa1csVWZF6
43f8kXg29+6Ul4gUZYwWSPUWArZwT1AGeEW01H9j4mo+UkcDJgu/sl7dUKFzTNOp
SS+bERi1O8p7EzL9g12jI8uawC83tK0fZNVfNyF5VavRFzWZl+sN3TkN6iCj8HM2
Lc7eGw+heBf9huypX7UAG2Zyj4y2HZLkiT55yGfSXHWfK+ujIEQvFV2J62MVCa1G
ImwHGOOI7XdXsoH6/aZnbOf/E1rGEsl24KAJ18bawtqBSG3SlO5aOCozaJ/s7GtB
wn/9NP9f7UdN9+KH4GE8Ajr+qv5Lv/iqgPCUchGcG6sLEFQgzAEbhSMDL+2tkyj1
V2WKDGssQ1/ONiZ6KUDPQbxit3IsAQMQk7UXXC/siz1dmbkgxtPDeFSxJjjtgxSm
t9BOl5HM9MROvOoI/60LZWFuI+o3phSsBA/VFrAtm+acP/54sOK4tzokzvTshhnn
AX9plIM42EBofufRiP1I6PX7M09RkHC4ekaROu+tSBDoKk5JC9DbSdT76PgJIO+y
GV9a+vXTcfARArVsaQmPX1euF7J3Z2KCIvS7LSmBw0kb9njx4lWS933cqDhFj3Ry
GRohXxkvj9gAg//+d+Qntq83DgYgWRmj4BvDe0PTb5bGsf1qO7Fnr6blXrGTGvtJ
DaKzqrwpYxvKyEgc9WkpAITe4I+nsPM2N6yFUtag2RSjNU6CKoqvDDiLVERGxBsn
PPUMD4T5t9a5XCSXKBhWUflzp5/QNvMUpivl9+KfERelxNHcg7tEd9B+t5gwuxm1
6JmS9c0pglAxBtadAHKuelFSoNBixKIZzCG8IRpCYbDIcP5wY4dSxHTm+MNMAwat
MUWv3xJu2RzjVoSMKuF7bBjJUbGwAIKcjddRf+sVF9iu1SWPXOKhJNFk+JGzd1bB
mEDpFnJ1TO/elHRrgMbN2lOEUm9AFA29ekJHJSRtiBvYKOi6eOHvHDHVOuafNEdg
P1xEgL/GRDP4hO731XDAcLKYsrDGmZu0fLbmJ3yFAE1VWyMw4762RXnnFbRbkFZI
ku8upfdedkgOXJK4TMPjTyNBGRQCym98OomHIO2a5osqgONrkk16YwompMn6RCuJ
9nMVb8RZU5HacQZE2iDlxzpfyrmUUyE/lLkpm/UG+Ho9ZpzY98LXaZmLlpJu4K9l
LJJGNe1bP9QitQItNyfwqiXJB2wxojixvn/khvPAwtwMgCBmpUPXGlG9sRpYtV22
zOJn7v7epfZhKnMNZWx6MnAg8oANBwjkgKRXTjs2nTp73v86E74BGO9NMwhLkE37
m7C9FmYQMY2FbkY70YsySBUwzMfCC16q1a9AzZFx6T8O5OX4e5VbscpD1MwTqORN
LjduHstdXRDm+29HPZBRmoUz2PGtuCoOyy4+31HoA5q36Oua/wZHQCBiawyZ3C6e
6kIGHzK8Yp3cx4wV47wAcwkUx/WT5Acv7nNloRAdQgtTiZZ1nJhnJFe7mKQsPcCg
aXg5sVU346Z1bXpczz6//e25+rpGXG+nIt/mQIrnpx/IRYHLr/RwDCW9eyWyvIgf
BB3nacwULfoGaTJIJCKEm2VOs7l5D0j2vX4r0XwpkbOmY2zZfFJeoqyi76fIikyw
Sv6pv3SATEeisXpdy5Bs3q7f4r2yi2re8SwW2hoT0aZEWRWGCaSlRBJpUhCiNLE7
bB3LH0VUpjLgxVvJ0UJwWVk7bPNV4EBrVrh1Oxv9v8pzoKaJfD03M+OHt3nnSind
Lz2HgXyKq9gX+95L1E+KO3znGBwDLngfWLuatqs+j99J3AMWRg0Q6ISSnpdna8ng
BlR8EwiThAzvTfwb3lOw40btqU0ySiT4Y2su9CT0g7FectZNm2m+JqRnK+tVKUIS
T3mJt9ANpmUYYrrdKIpqbznBsJgry2L2onrEhlcDzrxprqfIFT9F55SVNYzvxbTn
ENW6rWRTrkZ/AGuBw7hJfQVwbp2smAs2go6KDPMuVIv5T9UnuBCGCwe0tLRSQs8N
Xe9IXa5JNE/62WtM3R/hv2og5myQTJpWZhJXlLYEqvo4VCdeuQ6bCaCKxKqxHDnj
9EEHHMXQWMOzN3I6+Q7V7WtpQJ31yrQOIGu7AMm8d8CZbOkicIb9R1Gsa3SMjSae
ZuPHmFr46kzrx6OTbFbiX4+xgp76qEOXN6J1ah/JT3+s5N+uu9VjymZCBkteBs6b
Ayn9KxmhZJvO5elgZDpvOhdvPqeGCgIaEDTnHcImMiQ2hNUepOxOVlMU0x/dISyG
pB44L/G7OTYTZOqhpyK+q8m5HvGu5c4JiiQxorEVHiY5fUJ4XeDbSZeuqNt6+/lo
+29g+b59ujk6DaCn+4lM64hWQwRpRdrSXwJIfkGSlMMzNvDOO4KmWG1ZzAe1yNBj
2QyVWNQJ43d/8vJFnDohmvupB8nqtlVFL9qvFCoe/WCF/WI2ILLRjucVsRAMwZy/
ZlnOg/fQgWFvaunp+YVNaiav+kkfXtxv6RC7fsXLdEp6bcXfxZInaeIg4xk3FDVV
PuYWkoVXtn2wVidnOZCLAM3/hr5bh5oz8IacA/w9psS7TE7/ZflU0JbsyMCcqLGk
bajoxkkhiZOSeP6bk+2ybg==
`protect END_PROTECTED
