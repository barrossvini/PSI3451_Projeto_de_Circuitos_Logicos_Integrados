`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
noMgSK8Sl0AOyMMp5zvdaY5ShrwECbmiJA7Z5kz8GtSf2VfvqLmxG6qUBIPZEteK
JXWQ/VPm1puXJMpgdgLbZdzr0zclZwlQdGaabnA5jGf56x8jIW0BuHHGzSaNxW2+
AQpLpwUIxdc8+Gwf2vLOF25QSyc6seDjEdMh8W5ePMD+Gikad8/q6i2KmEHhIX+g
ZypXXDprKZcYd6ycDWfDJHylxmk/hN6J4akIC4KBkuvysgC0ojpGy83PJFnjQjPW
WsLUOig1LSjgqIi/hFVHg6dVZrWO1B2pgG46/gO5DyT14v0Us+vVfMc5B3ZaZsol
7ZiFkSxokHNeiWaTAKv3MLQ8bzIWaFeLyBrCAWJrTxJ/Q4nEGPSxmbf0B8WDDko6
qy6cJIuaxIkYsb3XbqUp5fPDDeg33uOqc207woSAZ7YToYj8O6Lb2/01MYgsxR1N
6aK9clIYehmkm5sPd+3o/iHyKgd2vBipR+2F2FbZqZY5JX9ao/rwezU/3c+KLYhs
ADud+sdxHpPGC31tnE0VQvhASnB8wPoRHQqvhCsc1ijIZL+0WuGNRgeyn6NdV3iA
xfABq7nhk642Vu6Iig1BOs5OTd5fGo6c7i5HymW5psHrBvIAll2Mx+nD4oZCgft3
EUgycu6r1mxBqLNoTVPAfM1TDRZiDt+cYbC4fCIi0ftjhqMs731QE7uFVsDrVX7C
1sxiQuZ6t/347hTJV5TIQ8cCh/HvkssLQeZOzjZ+eN43UHlszhOhNDdh3OLkdKZW
dM+1iJbWVyShL7UIEBPuFNDAFCpupXEt4sX8A0ow9dRcL8GcjqGRZg5ai7lE0/3A
s4cDfqPWDnrA/9Zla6uqsg0hbEwbb/VTTALFUtu25mvBJBInQAROjKKCjfPQ/nTb
o0dtDkoaEyueyKVKgOuyaqMYn9PvcukFkz4OdV3vlEdnOvooqc/MspEWKtw1gR6F
6hOs0+McpL0Nwr8lc5h8YI4ArFHDobljtM5I6vS9dHdqme+Zz/+dUzMlhWxLyKCx
pSORHN2wIU3zYqoex9Vs2p23nIcUwDLRL2L2eH3HX2Ssf4hyiSlRXMmudAoOQPu8
1zMBRFGpANPoen28M3uH8GHxghMbJD7Qh79O1Cgkd82lLVPcMDec8TdkRqMomvYm
ODbVrXIMrcdYpNB5Gan05EcQmx7qfZeqth8Ez0Myx3lQ0NKc2ap96qLjLDQvihUQ
+hAaN8Ip/LcoDNKnu7TKUCKpplkTEKleLfDT96MD54F1TdP+4yvo4neqOKVrkucC
ExHu2HurrAXLkQVnz6mc9moSnyJYrXHmKJIUBR+gi7MWE/gcnY0gvDzkB4EaKtJ9
N7ZaYV18wlX0H3/tSSQC2wVQvn8NIQPCrzKX9s3ylhU++QddX73rJVNTpgVbrdQJ
YDA0o18LPrxwBdTy3Piix1hCWlWHG022lcTMA1GZn6nm7ZKmCZPnFt+/pDFKhIaX
cjOIs6pm2kqv1lL31frgoGvhas3O8XYVJVpI2ta52Onw5Sm+uN46jKSK3mlGsvKC
jHy1RbbjYYpSbH+szkJ20jCQSqsyeC7m8Y6P24rNC8bEi6HWMV17EG8QD+whsGnp
dkaT4s3eCLGFlq096SObDu41uC9pGGlcJLr7S0UH+bJ5fZO9P9N6S6m18zj+Emi8
NxR6ajA2FsRvYfANUyj2wiUgAzLR55x7QdCQOd88ENFnRoZgB6HQvR+Fen9hbflL
s002jr+sqEONDrQjZBg/iIxeajuGLe7meLcobb91QXz3AFZiOU9EgolUQDlDumr/
HiJYCnobt0xErvvIzJsm8YJGUkgwWz15LHAyUjTrDL7O+cOj9N2+6zusxHECKw+j
b7gsk1lFsSmJoz9mg1fOZATYBsZ8m1jEM5+a6wsgMvBg0WGZwtG9NPLT6Vs21zwS
3cLwsDnYBpBswvehBDcstrwJa+3r9o2ZKmkdjjo6D2ntyR2nXQIOHRux8dk9kO+e
/hLsUy2u3eLL8s+iwTzW/f/R5myeGHtTXCgj0oSaWpLo5ZGAORkBpku3Nk04JPss
qTS8BkM98lFrGlHqfJBiXwTREztG8XPyIzqcujUJBhIVabE2JN/b3tdxm4squCeq
5ZL41pPNZmw2cBoAXGihDIU/Am4spjKGn5XWsr3rADnr5+FvaYflkOkgnHPW6bJS
KPa6sc3sKzaJha0+qFIijvfRtmOtyY37N5N5ZKc86YtRFXMgL3sPEAlUh5g1GRPY
0SJg/HCn3KWvvutvBvveGhwJ0/MtINzvSn+rv45H8wpmZvnh/vmhi0KaKbEiVD7O
HJ/K97bb6pkMA+Hebh4yxdDwkl8GYNsaQE0OtJA0CoYWV66E5QH0lWihe1q+AIRW
3e5+boSjyVX5DaoVRPeucwZC8b1ouvwce/SZLIT8LowS00nNah7nIpnUDUDfhXw/
YFnvYimvy6OsBZu/yec15yLKIODM9RAi793dvodyt2KOeofd2F8D+v1jDQAmRt/N
4d5DgxVBBVxzSdttL9i3TcPXwpKlbXlURHhcoQ11uMsN0cmBHEDfXYndGTOnso3c
tedaKcMADR2h0FrMqcfPvYQLQNE1I07MhKCHxfihlHu/KjH+4cVIdmBAk+d/shun
afOouTcbUCkN8l34mGL/AN1U/nc3qeBmCtsi9x3xcXl6jlpfRdcxuXtLZaWOp+9E
7ANjiGA6NkJK+CFDzhw8bKvskCg5gT4zOs+KWvTCOh66B1VchMM2PVwo0KX3c/Tf
xSdsVVi3Q0TEK0fo2P7tEcyGX2RkWnSsHfAazbIWBu5XvDkNxC2qppwf1IEcPbTj
V7VlPQTneHXI8BgrGWIuL0i2W2DEORt9ZKMVb22cXDcQzKvCEErgXgOfCommnLgH
sR0uylfgHcPsqgdyVc15w3LBP07+M1o8vK2eTdtnOiDXKixcEmeO7T51PKHkDduT
ACX0pq/H5D76utwvojzuaeEu9ijCa9mwijG0ZdnwOV1hBO8xmD0zuuYBjvQchBNw
Zu/W42zdfaFpTX+CJ4MD/LQ8VUzp5QiT7upVl4olkVF1zp0a4QXfsYeo454Bpkab
rG1Br3EiIJlcn4vva6eUqfO1Yquj3yOWR9eozBeTSQKnudgBun2Om/DGdZOrz4Jz
/Nhx/LnofbehidY3j/R2258dG9B3YRxrLd0BQHO32pYm4mGBlOFAibkzzdTR2xOz
DvxjYlU3UG29n34wgypnVCL4geKf2r+kZSWk0/9XgAG9YgbWTJoDdPBtxq8bKGNl
r0QgP8APTIkdmHEymgsD99et5ARhWhvonVecJPrfL4BuDZ459RHKlx0VbbASlnaF
YoGVCii1utRECSa5sLYvqcqaocaGgmldBUEZBU8avaWdtWYd7a50/msf9bKs/GXt
j39THPqN1J54af1DRglmQpCkog57e1RK5a18xv7WgvktAyLLgS26z116iqe8Wze+
xkhia4vOk8TJVBPk4HD29tEo2pvq6iTXvoANDj8VeF42O84SWNMpWEPRHkOtS/DF
xfYP6b69CbCvnCm9LJjo49adDyEnNxqyTdNVsQ0wdVD9oT+A/cI8gSMCiASZZT+8
WteAf/iVk08kEwVtHm8Hh9DfIEWu1MFVp156AHcmjhCHZyUlCCo4Uk3SYuC4vEhb
3Pn/RYfuUjuxoW0xtnTXlZZnOvGOu9cwoprmpFzdcy/Yc7FhrHjkTK0Kt5cpWGe3
RhJ26naWJDrsq3YBh1phhTGc3/MB49ERjUkbTjC1FWHDYTNNRiAPkCwU+CFW0x6F
FuhPhg/7UUwHLiIViCVoDlpN3vuC2DpOzDgOPoBBB0SqWSz1F0jX7CoeQlGTzocM
Y8IsdHewLF093CZT46PVXjq6u7oV2if9CMWutkMnhFcjlYO600xcH/EPNvNRzrKD
Tept0TfiqUA7BnepCYMvdej7ZH0qpMXNL0X/MrZ40irGOo7m7Whln3oOQe537mBH
Deuiz9IGvCXw5UBTyWQ0s/wzdlYhw7dZfueC1K9VtNx/7YcZs+5vn9wT+pASxhC0
P69Dz8e9hatLIcNQI/tBu/XG4zbLSw0r4JSqhrj3pb9Ku0Dc2G5IPqObQevApS2Y
HH+PfIFkT/w9tUBWoAQsm4q7o8yw0DE+vjoBmVfEPxVk+Kr3HkzZCpYueQcaJW6F
BhpyLXGiXtIKDn5fBPTe9P9Hknr9FH70JZMcWPBIoY8l27Aie8Y8mLCtcVO+qdiG
vaNWn+cI4vH/GrBnel0P560t6iwPRab4ZlzfdQ5veZrAUefck+097pZIrUAojGIL
z+DITXS73hzfvuA0Cv/3r7CpMK7vqR+I8H4RuZtSNTCyrHI9xddoK85kpTP95RfO
heyH5wy9tx+vn+z7dxHVfoD0fGDVrnXIE2ViKUEe2we42UjaJE0gxcEWNpD0ybk7
gN9z5eoX+a0CG8GTlBLZfkxKO2GsL6L29yL9U/25WQbofu2S7aNfEW+LP8KQ6Qz6
9PVsi+OTdhe/OZSGERxZZUkLRevRhesmHsFR4AWilCwu0BX7609WuFrJHjXuLEPq
pLnGsY2cM325SPunD52ASViYrMR0n9dcXuGDF7W5HEgeX8aj/AG7X0pu31/9bb0V
c1d5zJHWIoBO7LHBLkeicXl7VGsfyZk6qkLgvpe312BAxDqAfPAn01eIhRmrH2dU
YjD8PWZwXrXMD4qeXSso0BbfQUKwojwjP2ii/5/T8mP8wRF4VH8BTdvyhQfb/+nW
8YyeVFXMscdv2NAMpIZLC6heelGh2GUfqM0C4mYPa/gvjxhUbegRMYUXRVYdJvUB
GklKkmrsKDrSZQGCkyi/dQI9eE5roHd/bHdUku9j7Pm1nf1F+RmB6kAikPCCIPuL
9rfL/nK4Z4dHLcYxrZQksjxBYvOOAiaM72RMlIt0SZ47Wa6vFzE+R3dscfIqrg63
QhebgeX+kJUN26LFmM8G81ab9OcMxOn4qV/ZMWXH05v4jujLbpRbHVROJp2DpN2s
CJCvtr4wxB3PaHPqEgyo3HwlX2VfJdjDDk9yvj/5sjfrK0M0LoJOgjkr9x9YattN
z8N7UaPOZ6ntoT97Q/8lq+2qS8ulGEPcJQ+y1uiGUGFEiqvLjDETWRDTyTZyswIF
bNKr+worMO81BjGqcupLZ6zu0xq7uPTE+CpuxYEMzTBfOV72lHL/5E72HQ6dvClg
4RnEgRtjUlQBe1K42azVtkLrDEoL+d00YI7iEJIzZvicZgzOs328SfP9WNKU2lix
o75OH5iegvGww1YRdXEOvZ9AnGlORbeDZojuvU6NShMit2sNxa7a32ms9e4GxwIa
f5uskFXCRVk52SGiFENnvWRdO3vY+5LYr4R/Fmr2FN0xTVW/VlLOOY+a04R6RTo2
zQF8x/XmesUStvYQr09/blqGj2fyeEvLkwy+ixKdUuRbfOgKEa2wMEn2bH+hZ4OC
U+NA30P+TexbIM3ouBl6I2obDixwlNx49WMfi1WCFGNMEnAEhVAXKmr9bpPiSjcc
3YaBVB19f+SDworm6R+UAFXa2C8+cX1lz3/XMsZ8cHnjb193WnDwClV4fVUnQfFN
uhb6x/1VE5JKT2tjW0N6cybuRII2te70C29E6TKHEaKes/+RQeCbUbLOscSqk2Yq
++V4L6CnXNew679L6MuG700iccvp4fUs5059C8dsw3WPACR3p+F8OZOOaBldsoY9
E1u9fgipzlDyJZLO0sqpBVZS//hH/wsu2rqCNDj+QnyEJwQbkJJ7SlHzXnQrHWgN
wM2wiASr0apzGTyktubwGr/DN66MiYAKy0e5vbj+eZNMnXf2P4E9gjGUFqcZd1WP
PyKuLkChx85X/AS/j8GrwYS0152r/zuiGunaS2d2pWj5hx13V1vK8sZ9blsHNqsb
Se6bzW6vW2Y/9jGSUJhmD3wkIA+MGCojs6Dp9lCcRv/M2EYLRjUa4FEq4Z9jmRPQ
Y0BIPs6H52xZm/u/Er43VGDq4n2oOgFHd7h3+1Xcmzo71Nd41cfRb8L4qVpcAF2q
k6Wi4Uo7rMpFw0QyVPdfKLcHVwxPZyNlNtVtgNUyedhygiBKLE3v7YjU6l2f2hHk
yTeeb7VKb48Oanilv1mM6sX1J7gc/5AcR7jhiKg+cneOd8e8HtMWj7Qq+75Cy9B4
p/mnPXWsQB0wCP6+6bgnCTlGIBAvpWoDqwXhzTGqIcc/7GmxWEhEwgF23CVFSJuZ
rDLc4HWawPrSoM4sdUoAOavfmWeqz4QqgsJrraU8zqfc1plFkVaUOwBwa5ff/DU5
CZOmu05HdLvYkHANa6giHEyfFoA/s79l+MhBEbpTqk95LC2DJfs9v5HuSaBwru2W
fIgHStGuzFeWLiFLmP1m0J9/mhsSq+Ul2zGCpHOILZHLYkYLuYpeFvgzHGyhPqdW
ruQEMjFYkRCHZkR8PqVff+KijBtHsEC/B3mUNSQxYTiUMfU6lgakl4q3lQ0O4m6Z
yDfLAolPKrfw8+4lsebBdo1W/OzShJAWmTpuhV9N9sTHTdWQ3LKq3SWxM4NG5EWf
p0VAcWJaXpVp5cxZj4/mcFjcYjUTSd5ZUexLot8Be2WZ8qJCYFs1JAnjJSBpeKq9
LjClqyVZmjQR31ooPSyh+QOFkqnG4mnAnDlnIiEJFm3WPEK1xY9VlR4MQJq+g9m1
/2p6GRMuozP7DU4chNl8uq0g5Ov6BgKVXzc//1wJmLjOjdcWa/JLAJLTM/Kn+9YH
w42L+v5eTWvSZ8IfA55NoSltuwsNcCs36NgOBRQiCZiPGaigI/VQwLuY9lCvpwkr
N9i1M1/wOU1gqTlv787yTD3zWirP++Mz3gQtUnipLTmz9aunBNH/3qQPzEjD6rqd
/d16sZIjUU9QEUQNajgmDqDIuClmrvaoDjBvquhPMTfRoYJozl04nlkZpZy07eDV
rsMhAPTHoUqx60KibYPs94Bzpv+DhfueTlFWsOWw38cNvh75PqzgmfOybl6544ml
4t3cKaGPtVwCtonEaoZlwKil+46XIgP+Z2RTohUD+fhbhxPjjc6BbMHOB1CHyhUA
Wx/LJsAre9mHnrZHApGw9cfgVyh6fZr8RbuQr/X359bD8GSsrXF5ybovGeao38jm
51vcDb4Ty0qeaLOpNj+gNEKPyU50DIp95+l3oh3pc9B/Zk+gi7GNdzn1J+XAcnjK
xPrmK1XP9pTaFxFPACuY0XsTGM+owbuTV5szjIfauWpsG/TKvE7Xf+TzCKYgZXbU
xPXm9MysZxFwei/WuPhjIQQTYZ6tz289GlTMSVfaVTJ97kOapf82WBFa/WZkaWtp
oatjafkhGDkUSdv98DEHNZ59WmTIEJW8Vpk8htF0eEKx4pqPdUuDwHLQl4y1xa4K
XMc5D0gN9vBkXJiep4gIXhem7tuNpvs9Et3N5AEE/S3fwY1KGEinXHj6S4sY/Dv+
C7M0IKnkox21xnnkvQ2kTMlsCClnaIP7YfARvff4pY9/9Isy0Sja3MLtbAr00vJM
4q9hgYJDJSF4AEC1IWEvb1EPBAJliy8YIvhb7QB1jxSbGXpQyNgrof7KU/citCjp
KvH12RNfeWV0JleEz6UWoVWSe4yguH/CgXBj4nufOrh53+E+75oEqKKF2goLsTBk
V4YiFtL+Uf+wK+bJXT8RNW58qT7qw8W9lgFMNpM6GQ/v68tIPHvtLBHjlOg5yBq0
vlsthbmboMlq/sA/QIVN3FfyOCwXWJVSeoGmUP/N3qcVoUofqrrfjHTRehdzPBQ9
NJP2j+AogZjLCPDuceQtwP8kYhr+uIQDA2qnN5euovDOdt6O1fM4Vg6tvQnTCsRf
aDnnHyggRb2Efg0J2YQQOQl8RzJyfZmukS7BnDemLuWDK+90r3AHJEQfWKkTQ7fg
BlGujYdEC1ZICD8ETHaHzTollV0fCgLilpQ/gI9P/UGq/oOEPwvDI04IOCwZet89
t2e2FuzGs9WJxZy/VFqj3oF8T7gniVbu8JU1+1uAna8WPUpWbF680qVLTe5E7qes
q5bDKcnrFnsrsWhyZbw8z2RsDa0XLn73JRQBdHwgOlaWYzF4u9F2e9GmvdY+rIQL
rUKomzgGsvBIXbun40tZL8rVGdcb/ZdMuZzJswOcCFYdeQNDxFxSt4wJNaSviAyK
2rpFIdKu3wwY0EpBhv4DbuIwXQqZznUOqbOSZQ++wYfJh+Aru8pFYXwq9evoZI7N
vFwL3l56eNKQ9LCZ1djfcDk2nuXlGGe3yEh9j+vlgzOegF8bitUnK2hphVWzTptm
AJzy2f7r59BKFUNd6GA91zx+LndzJiRijxwBr8l0eCzLkWhHEFInEBhP0/DLH31y
OMC8O0b4mYhtqjcZKIAH/NSjfhQEUTCXgdYuOR+98A9BOCZyZXokF8xYF908RED+
JAvkD04JRrqcqp7XQnns5YYGs869s9gGWS+/MffZ0fYiIgQ7TF3P9jBQq0w1Karc
sMh7rULqFRnu1DFbRgbUb83Vb4D1CproL1vB80vsvNGqR04VHYrFqpzYYMwJRbAw
T+QjAkWj4V+jrRugshycgo22B9S7PzwK3X1qR7ASIJSID9jacg2c4k2Kxvr7DaE6
28O3yN7bUHmZLyMxi5fDl32AWrYLzTDUS9zjPekbd3ZTo80E4t5r59Lw6tfPJIFy
XPnTaIPxMFG2l+29A+7BMLUb2oV+DyfaBLHGf4xONTLutaKHaUrc1Idc9LTl2pvi
bwyo8NeXFQzDUQ4a+DW4W6K5AGTLRw4juZGOYXbDsk/6FZyJkA+FUtQsxzCUzzE/
XD7SQ6hhf+mad2D42t9NunNJGuGHnZ/XY8ybeF8r6T1V3v/rlTP2v6YVN/oaKgjm
UORbs1z59R0vQim+04pFg+UvtWykg8SywUANT6m5Qudc8yvxQ8zdB7UOerpKTH0s
M4BHbNKmOxoj/HTmwvFvVuYCQ6L6zikx2Pfu9oGiLxoAdJtPUT2FYizpbsOjeLvn
EyUzymbpa9xVlDNtJ815Es1aO8Z1ad9S8DeQ1nTqHWFejAHRdIIbgmaompfBACIi
mIJhsNjPzf/pbS68DbDl7cnM+YgfSb14VV8d1+AzD72faGBYV6y/PKD+6xi4AoCd
+1QgWwfjYutwlTwCLXcIwun5WpWCn/iZoNnebcvZc3Gfa5N7ikqY5yKxm+lQMaoT
OXK5jvrYjJTSC3TqJUYriWiFVUTJOJ60XtkvuhNzt71VzthlKfpBZK6uA3nTyDA1
i+UXRgdmapopT4neGmWsRqk45Wl8OtRn9JCnx8dknCHDLoXYNbWq7AK0fTdgNlP6
vQ3HZWfKBtYTzX4iTBRFYnHc0CGzHncigypw+llQzm7lF1h50YuLjXsSrll2lFwu
x7TIPRS8HzB4MfOjJWgC6rW055Av46RQPjzjfSDrK/y1/Xuy1R+G1MkF3fFpcWWQ
Li6OVQ2PmxHvUiyMTXaig+p1+d/KOLkRS5Egr8Z8H0yXtTazfyvVKttBX3b0SaAv
yK5nipZpNvKPPj0RKhYZTKw1EnBXnZIXw0X/rZq4XqtXOq1YJXZLVevPn1yMTf/k
NQ3PFHJlYFGA4mGJMnENQE4yjBLNLxMFTieX/mfHQ5M7oXxzIjF+VqSMKaIkDQ5E
At8FIawzDfGdshh0QQ8NFTcLmZpcPcTW71piNCOzdz2fcvAKDX0VOt6bOohpE6C4
6IK5uAHTNTnXnpOXU+S+qSt/EgTtA9HCotu4EylKo/EhnuQsJC8GMXbWBGUrTM0t
/z9rWconBlrOLkpIyBuLxZWNu17y6BC0Uu+x12rAsvZAA/kO72UNwbIRZX5iOWuU
53BPTBFnsVHeHMjTtqpjRnOf8+FmX75bNx9Ijfpbg1fs0Yo6yM8noGhJnwluK/OD
+4/6D7JE2FiCAnP54kAozMs6uoNZAIj6WJQUdGEN1PWB7owSJzE/eW3jc8edVWIS
dSuS7mkpIkhzhESN5X+/UILZWCQUGAYAqkLusDalGrMzLzlyQag1s+q6kec4HHmU
OuRS7kBACKvsFH0e8IoGwXDmx0B4Po5CimzfKMmdAPbicZ+DBtWl7MYYLIuk0yvo
5QBWvWp6aQkeY4LtKLBYsFG6A23mcPXgn5LdUPpi5GV5n7S9C7MfY4qFSg4lrIiD
epkXHgDH0D9eIy0X83HUKgq7Ze6+hQbl3ej7T+pvE0hSQgjQGPAj4DLxtmn7DQQo
OKOihk7NVa0IoItj5MzH7sAlMXVezqNBUDkOBRwCLWP7anR/Htt3agcS7mn9LGic
t1y5f0qwl0U4yDnfiQEJB7pYYWKmT2DxXsk5I9KD0DOp7iL7mj+jJbLtVBm79GNu
QtQg4H3MH4Mc4zKgsOCf5hEd/ZAZnxw4rj8U6t1haxf+lrFyTr82v3lEKkYhX5sk
pb5PthKBrUe+L6JqWWuTahM44bRgT9skBAE5Z1BWS870G3kYvwN2pIjcCNrYbsv5
ORUpHrc6WxEEiT3YsSohSHTwKSRBKGa5YaCyeiNi0JyhmqXipTW7eHUTImMl7uZv
6UKeczWP5sGE1u952ki6j1aLdNDCJSv10TB1ulvNqaZXy0gGM4LQ01Hlz0XdFlXl
ZTZKdHQvdJkdRzFh5uK7YsQA6fkBtEA8qhp5WZwke0M8ZwtsLuSEc3qUx/KxIr/2
fA1y0R6RVpkcZ25T6UCoKVDMm9WSKgeTltYUJGo8evjqgGYaAuoT3/dbYt7gMXFp
7yC0/dHVoYqXI7hizYoNiewkKkpstiPAa/W49gG086CLYEQP3GQ5bZi9RuKiqzTp
uCJm0N9BNHVh1n/anszrhkrnydAUXg6V7YBxgY5JQcekMnDwCPCk9GH5ghbeEkwY
Lag/1YtV+/nl1nKV5xU+52vwbiWsP12zoobZaMp/pwPyrIWZTiy0JZ50hXSg4fnb
`protect END_PROTECTED
