`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uMpD3KF3C5XZs6Ha03w2Lnf1+np/1ub6t2Gpy3GRMdCny173onBSHutF/dLHdI/L
dc4HJDjddTqgI2f1MClzE30gASM3fDRgv9zascDlD08wnEeh037dr93ZcKxjjii9
4YtejUfE0SV3BFIJ4W+2tz23le4Efbyf7W7uufvuhk2LwGDIpOqgnNYf1/Vrf9DK
1TSbZjXGWR3eMHt45FYv1U9RhpIID6ISperaagxUfN0kthMIjWFBS2Lwt0z5aGEN
6rJsgEV2eahaRADyDvV4WqU24PmOqYCSDkTyGlF2Ua+FXgnD58jhnVGP7F71Ij0t
2ArGWqg64dYIUJjYL1CZRCRywzFsH2GXxzics0wMn7R5nmUUAvCDFC8d9AhqQHB8
I1ZL96N/6UZhq2b0m86Kv9Sg1GzI0rDz9WmUShNx9PWsUewwv0BUu3yKgCfKMaLz
cmFYpNUx8fAfJdXhziYbGiKVA9PbRQ85UFm4knaa4mrgHxPhrT3Yoe4DNy2yYmIq
JjUavH1MVCmM7EVrd/jJzyuAfZiUhx190BMGjDzqgOfZ2XSKgtvq1G7oqY6y+Uma
YSeRzG2YWuD3gbpYVEaHHXRjYN5zf9sOpecjnucTxPkH1iJG537lRHsv8/bXXeVb
DGkUxPp8yTGu+Mx8R4luzdsQyxuq3orCGSqYZuLIytsfgIYo9NpNK1fpqMG8zUiO
xanfWcmVk9AbEagxODnwFoHgKu+VRPRT6ZsL1hMJSyBboJ6xNeZrG+AXLG9SYeD/
5wz08ILC7WbSTwNO8Mvx/GMp3Yi7RDwbe42446dWdSCx6HxLZldkwpat4IlR61Aq
DxoSi2/PZaQDHYIkZQVZ14jW9TkQEhMDepG9bfoz2ZY7wWzP78oVxiWiPDBfanNV
WHUxJk8ald+0oNuVslA0D46vPEfifOFgHntrmuf9RkZHqEGzw2sqyi6LcAehrcVo
OXxqGOEuAYesDU+UHTgEJkiGibjlK+FBmZTounePhFbWdFFz5inYgCIA/rD6LdJh
k2i/hZr3Y0XutLDySk0tjTGguJ+aR1Bhy9+bWkXVhZX6WtZaVOxF57GhYXwziI12
G078/GRAbc2ugmUihAbZe0VcRf5HzqFMt+Ig+WescFQWLzDyEU3paRkOQsKP7tf+
TxoIjJNJmkkvTsG6N16DssQkAzGJEcpsE3VxIcuD41oBsqI8tPpFTYg3DQwwjbX/
EIbx+mk85lDylXbtscUDWvVOCrJHyB+Gyz3ijOB+lqQuoCRXoHvzcTAK+WZmi9kD
mtzBWAMj+Ub5PWe1YnrcMJtW/Lxnah0soY9U5FwsKHGOdCBMsoKIsKFtLAGnp2pM
Gn/80F64SzNMBiAYrEMs26klyfmqTW4FBPjMy/uE50TUpMQGgpbKAZamV7/Ybd99
xUWHOrIS1Ed7Ql7IxeOKrWGsiJHVOR9/VwgCk+9yohdoK1vcXa2xENTWkDkac29I
QEOYL/F8bE+FW2BzJMqqd09VYDNqmyexjqb3xTpaAxihbhXP/7kTEqrknWi42KZW
RqqQz6cyreInIR0mddDMTu2E5zLVlf4ae55L57oqpWGXIAtFw+VjI6qKJI9vKMen
L/ah61bs0dnZ0oVhZLFHBr2g1M7+9IkThKl7g4HJeXjj9xJ4wnTEV1YYeYZnyBEj
Pz6RrtIrTFsnPNOSKWNAC0NG2vXplXuv75N42sBWIMdGZ01WREvQsgzgzP6QWwyw
pylIHOXlnNMOoTQNXRitn9BIwSX494ZgX6+2jBr/x2U+N24DYI81ROSTZOdgEyez
A3tDLffys9PjNPUDiehxe08im0F4YAmb09y/uaFpn5fT+WxiZdlf0huQ35mv2V+k
1SGEk9X96T8+AnhWDJuGR62Y0/rj3bI59jptwEM5nZRNOvvX92eM2ITW8fso343x
JjDmwTaCLPx0/e+7FYXTA7qludqYrnwe8j0jaGdEbLudn0EOYgIPzRpgPX2xTLVW
gJavXhu5mjJiIiaCjeAmXZRPX314R1hGSJgY+PO8IYfkPLrN9/EK8j7WatqSoLHU
DhKd5RfJa7Cq0QoGT5rrHKZ+jMDhyD/3ToCd5/i0gxZO6Ye5Ff8IXu4JYDtmPjBe
abrpF0WXk93nT/Xl//sEY04ZfWZ2cat5vOBO5qj+hwuxzSGudfnFlRnflSmPvoQp
Qg7NEf7qGD7/NFtrhXJA9Mmy7yul7rEljiPzjfu+Dlv1SgjBpssMO3JAYLWiD7Pi
W4RTMoor0MyDv+XQtRhSX1VSEe4LfiSyTJiex8HwAHCNUFEnYP658swNH1Ej+1tJ
HJN3oW2J0/7T6Kp3pBsiy++lMsjMp54O0n9L5WfO3YUejOPso2YffbblONqILq2q
WHPRf6nrvWC9IjYi9yAsq2v3QssCtP693HVPNLUoJ5G1g7gUvIbeK6n1YjMBnFad
4IMxXxLOOAug1L7gvZi16qz3ESvaBM/bfB9wLKtVnCeMFHo6L8rneSB8Kr6VMgO3
ko3eEdei+fAHxs2FM8yNeC1Vav6kbaQFHRkqZsXVGSROfXSin+gmD0Ws1Ytx8NPP
VLDuFeDja75IIZ26Gc3jGXc8OIr8753warODDsk6XNkYtGPxLf8gmDCaMi6Dr1rG
ljZebKr0hEdZGdOI/mg7tUXSzOawnYSgPs0+mZ9RnXDfThydFiXNI6zuQKE8s8Wd
PiAM1Ukhg0uiaBDrlCuRWTK16tPjPP/+ClkfWMJFYhG1ENpz5qLf4+PyA6CM3xd9
I6r4oTrkyVvk1V1EGUMnHU5VpOsmhHmWNFc67UYv2N37AyMe8+aUOEKSHru4ZlWZ
DV8HSs4ARPRjyWMe2mI9Nr1CL6E7+qg3HSr+nvuU8iTGijIsVeVCGsFHi0vjnYVm
X8lvp0kisatvaq/GJooTcP9mwCjHW2cVFlv5wUSQi1d9gaIMWx6zZODFx/PuTFjH
UqqqYCg2aJsjPN/2eVI9O4bgK+2dtYZph8VU9wyVueaE0NIVdMo05RRvYICV0Mqc
W0BENkviLwTS/FvVSTF3D3c35WCt9n6hAZkPOZCh44enoeKmKHeY8+xJtNVg9zbE
sH2SAEbfry36gnWYGzlnSBNPmGgjRPbZBJ3hsD7sbuqBBIr6nY65lawerB9x/gT6
cYJqvubvWSMFfEodAePuhsCo4WiHMNZXDpX0ITI7XVXQeCRCYRQ9ldBZ5kjEmsnA
MeLDj+tCdYy8KCSLdD3HGilBhES8mfOKTKDbovjpnWDAZa8ny3KITJxGdmIzl4CA
6PTkWmPIxS7J25hHDnbGerS910UOTnhL2X+AlmT3TwSZ9uK69d2d9g1/LUh0V8Yn
OslkeH1o1FIURO8jhCI0kGmiVGFP0cTXNJp8MgKgNh49a08zuDosaCIHs5bh5muu
SSS5nwrHtW5mr3JFZ/c9mwqtQSuiB7CIMzW2IDxSB7Z3mKH/LwD8k5I2UmITEJPe
vt03G/t7nywnwqB4jRryxuuIzjmuuWpxso/WUKSvlJj2lIP6RtUXG3TQPazTplQe
dawzB67uuzqz6M176yN6nSAj9oORubKEjJnj4xPokB3UARUfjSdgrx2IP7xSSlJN
dZ9HENqgZD+z5+CG1yfbzEPLi0+lGK0IKP/bCMusD6seTUDre58P8tc+fyNqx9rj
j1VtUwVjCyGY4Fn6v/Tdu38cefXKtQp7PwkTh48DJJJFioj9OVTmqCedEKrI4BiW
FcCeS3ZgKkd19eDOzc33kIoLkECPMl/6FoY+gV/ofkT2EJnBLmiP0hMn97WVn7+9
fp4Lni4WbN9crMxfSu22HZGpNrKTu38R1A6n9UpZyZe8E/I7/8DqYiBmptk9cSPT
QIEVmtZTrn2rN3rrXEUIjR0M5akWjbNmBZ9r2rYwWssO7FEcNeS6FPfedWk7xblE
EaEWoL4tEpBkS31ruwZTkigB8kSYTXPDjl2Fml1D9eFpjGlRRW3vG+Pzae81E/Ud
0aidJxW/7eSdLKDp2Jj+IiJoVAVcPcaO3DFYMQ8qJQjskKjPIHR/42P0NHBLNXzZ
gWU1rf0VpeGafDtAm28K3RBB9Uvh+CqwKVPh0CEWBuAaq0AkhT5PtCVep+XWfjMs
ZilDySYfT/QjCwxtq6eNnA3SXgOAfUCj/me5Mvte/EI7IYQvtpFq2n22pyhCdNNN
5i8DeuxQVQZaVl4DrJLYypwMtROnfJNE2MBSEtBSAWdOuUPgr1/bO7VU7aoe9NOs
oEt6IytXrMCsccZOv0z82zK15lHruugJh0jahQQQKNI76i5dohMcYtsIFiCRqr3W
dv8lq+RQfSORcQVUFP8qUjyqrONUqTRboNG7cehlw8q9hwn3eX+PG85PYGvW4RZs
McNk0n3gmxk2yrzP3/2I757e3xZVn8lyjMGxA8lgYaPu+hZpyMM4SngzSQmFZH5o
eHjYVaJxavSJFtYh1AY8sbjxjB0HNwErQML0+qNM9KIWR7fv5dYVtUGbS3L0XyGO
hpO4izUwGncQHNxwahpKV4ae5wLlA+bYs/xloukdWJGGxuFimWBTXQUMshY4fQSZ
iCM02H5JJVd2ewlzASytgAmnQ1+CFIaU6aup0Z9XYgpC+zbxcx9Nihsva5RIkYMp
7a/VaMJGQwhqkXLsylK6nPCIWNm9Ko4EGghi5eBbrM3CjuTFPRRkRXVsTdAAt9M4
swZMbqb9Sc8yGj5PwSc+AzhsFPjdTeRqwNB132FLlHCfTeqNWMSO9Nv8uNi4CPgs
l80hwtitILEuKtEAvTJkvStSK5dEYkr+zJoTUA8RMLTdEBIrApUoShwU+nsUrfxz
IhhEHn/YNfXBoZWLyliUhlEXIY31Ai2yTkY12jCvK2YuNQxbY9qwTx4ldjRL7c7z
QxSiNzOOCzhnQ7kkU7ibzuq1x9s10oVCyYyboWJm4dE6Dw9zggJp2iVUK+uiXfhY
9EcfiWuIg/QMGV2LUFL63rSEvzag0U0G9Jo6MBDJAMHPNVU6GV7bG86C72kOJB3I
IexThbCb1t1f0CHSYNTNk/gZy8qRWpdTuweD0loBhy8XS1xHSB2k9X35/BE+lsC8
fjetka9hQrW0qn9Kaw6vMFh/I0n9WcofqRL0EXfh/PjfGT3uDhVLE2K1OYmmvyAZ
C7nKw4uQMjMihVH7uqIdDOzcJyHc3xTzmrggS/dPZHtboby4Gyf0j957RU3TN7Jf
Nqn2MA3NtH/hgmBncONy882TA1OLyMNzxe1Rg1iLeoIng3VJerLyy3fC8vBMDOas
Fl8Mg+ltFwhsIhPiUVG6DkzE+fpStgXi3ThvyZEgwePbE8a7SE3XfzSg9lKWaCyr
xyvIaRcE1i111lZtuBsWME3B9UkUBJ+fzY30Vbm3hYXyBcIzUP8qYpKIa3hp6YDT
3NXhXvTMIYTNCNQ++huN/dNI+1Tamj5B33RwY/dVW3hbKKMXAcVB3TJ50w75vMWX
ip0wJQGZGRMOVUDi8M5FybuFX9FQfbpExzlhr9GE7PT5Yj++9GWOPXMoNxozvrRt
Ke2mYYlzagG7LXlyIKJ3Hb97suzpmhS5vzvosHr68HgJftOdjS79Jjt3HUKTDNsm
PQqR70hCYCOkl+1hz3SuYJiPjwyDSbR1Mw1VO5z2zKaR/TJjcds5do35/yCNAnCu
8yFD4tkX0DvNn+LgubTYKg==
`protect END_PROTECTED
