`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/O0ESJqWNTcZpJOjkZRyNd2+JNN6RgO47LgZaqu+KxqPCBwFHhgWpXBmbNicHal
GimC0XD8mzA5LM/btn8xyoVlx2yWgrtBMFcghFZon0fqiM3X7tJB3AuxfQadfoli
zi2/OmWdf3PS2Z62RwQB+ksHJz/ZRyzGqcjuOX+rKWT4Cg61hQEfAnm8OVFz9MFn
iRbjZOyBKM5NgmysIM/B3LSshpOhscjGHrxdHfa2YL4x/ndSMCXTyHibhUEGIZT1
HPICXXTbRcOTsyVnrjEdBZ55KDXdMmBaL1xv7m/NAyO1e6dOFM2UUqjKH1SQNGuc
TEoRijSDd+mtol3KYGZHorxdfiDjY8MYXOPuUkiff7tvCoYiTpUowdBBUMiYizFO
pTtGWzfSBEfjHFH4+uK5mToReXS9fCwgeWDKqns1tHkGEqpCse4dUmzLTyDWAFRg
v5rHxLER1CNYA+aKk+Z8AF9AXkv1FuZ3gk3TMHJwcNoeXxd1+CWmEx0pxsb8+qiU
0UWrKEWghH7yVesZ6DcdLasHzZfmCkKQn3erq/0cbYGb4LHIVKRZgc2oK5PGwefh
lrr1F4SPcIA8ThcQ6gsLNIpwPgSVtJCMyyN0fONHh2w08uohyFLgjgcvjbBNNyGD
CAwUzjEex0WFIU8AKF3GmcfJ1VHUCTEHjmNSTku2LoItn05Mch0rXl9+M7EVDdB7
sTt2A4Bxswibg1W1Sjr2in867XTdyPRRR/x/8FT29deZSRU/kA/4nE3ByvXuZ1f7
z2zF/xhO/GQNBeWJDXPUi5+jdN7NUT/nothn/yn706dh3JHqTGiWQbo9vgYtD/8y
UiP162yyX2bqwlkvsIHwrMWvLCqF1NQoJWiB5CroS0u72Itroq2gHCyaHMpN/TAN
4iON2cwklxayfhycoGYPZGZxJO8f7xrqqr8PCX8hS/fBiqUUX34sMb7q3MdyNeU1
iLPuNr1fCJiqH3KAsDi4RrRe5QYLiQW6bcDHOY0M1YBpv2Gew+cuY01ONm3Od4BR
5JA03/u8vQgdHsNCWXf/F5Sn2L2PfsULwzZDzgFD4hNnprvYFsExQLOdWSsDRZic
1oX6eof948/PdX5mNmjls/0Tx0y4+xrQb0O8RJbR5DG1hzgIpRXLvg9JDEjawAia
r+PZG9si62zM0XSomjzrXhfS8RnLwAXGLf7OkRWbt5LZqqfeIiyxx5DxVgLuj7hT
ht2ttYC6TB5yoIxnknsqX6F/Ajc1NHuxNUVtJtNKqL/KuJRS7Tm6qFM4Avy9AJzX
64SLDW5LO47zz388HyLDGCl+KKpHNy2m20RoTCkflCnOOgZaS0gdLXnrOsXcXFQI
7VoaWBY7TMF5BEsOtNzN+HIPsIY9MacAcLIcEE2E5KS1MEYx5qbvWoIApYMfWEqM
5uiuXG5CxkafbjzM9vhPDY3GLP3HMm8mPG5BPhdZ2ugh6FcJP/jvwSe4LP6m8ufY
TJ5cKwh28cn4hJDl/kyinYl5NA/Lue1DLcD7MF0lfCWCiKXGy2J3VQFn+VcXKK7q
R8fXaaC9kX6TWD5gkkYC6MKI7UTM8XqvL3U0iZlZM+3tQHbR1I0tsDSuQMiF0qRo
AsmeWtjQcBmlMvUnL1qlRf51/enTdCcfRjfGzTCXhIrIeIrSuhvzoReI6esi55m4
TpF5iJ9GrUDigFqxhWwkSD8ZpVGugwoam/eMkbrdrYU9zFnu+cQQVvGGx2nYzZ9R
cSHd2Tn9VAOCwhP2oLeZ8iHBuuBZPiqGIQCK7ihDY28CGuH+Z2X/2raJZ3zyBP0A
9VioKGfTy0eLVXMDKgSFmyyWIAwJ8g3YmlRHnclYSNPgMhz1W78F949lZPyCKGTx
diMzV6p97cM/BgGcLpZe98BPsdpZ6V+/s2fuhvAd5pH1tPHTaNtUWtsmOf7JhALI
x8u9W6Scs3B4Im6VuhRe1iVGRoVHOgm74hEL2whiMa9LCecYYWz6B9pEHegCC4Fn
klZUjxvc5pu1yIP9bStiVKjmpYW7kNiBUnkJ0TU3sT+Ufufo9Zessm/V8dPblP+b
ljbmAQNpHBP3835MNQ8fiz6UTBo5OAVqd8x/nAwXdHXIiycmlbe0cUXoXZgYVJjc
dpE5OiZVTg/rjAfgDYkNMiHGFOKSI+K5MGsn2uLzWoNCHvoQvs9thU+HvAsC5tes
dXs2qm0e8ubCrAjlkPZAkLY3S2nip3dKL3PTdUvhkz3BOfjVc+yRi86dNuU05n1g
5ILucN2APWa7tlqbrXJfpG71FFf84bW4AP8N2XDmiH9IFmj2SA7YA39nOL4Vb92b
a7WvSL9nxiVHMxJ7tKSdzn3/7iZyg/vKAUimWyIZyynx5vROVLPHTmz9DALEiXxq
VIKkwmER4rkfJaUxD+PdcWBXLwkVFircO4GWk9thO7rQ8tUvF21T92Wwua+tbCrc
U32WJ5i/1ivre9jh03BFsYdMqD9kgGVJS5bOsDjwTLIKgau5E3hYVD34H8ZPsSP/
g9YldWGON+ih3XHxuumUPZssQ73pBxZlNIxKe0Dd4DcJCz98qV4ak9IKOgsDQiSI
XdtiJHv0Pae5QejuVo1SvddAo20pvQQFiZ8q3rlGWybRD59d7GyupVhzf/4sFfON
+MGCl99UAQ1M4PDq1ENkfsrY/m3rKVobZ1BsfY57K7I8ISZK7VhCCHadVoyKkgNY
davCr0Nzm19bKZw35ZKU0yf1D8ikBJeJGEod6PAtKgD1OceurOZtmGJhVtYTc3CS
EJvN9mXWpLecqafc1Dq9Ya+7HYNJcTqrXjDP7Kzx2vqRHzyufnAUM49/MP6aAqp8
lr88WjvcOhejLnoW4y6PlAYzX5fHe2EYLhtK3yIOIa4PvKbG5xWXibBgv+DGJkS4
l1rl75DS5tMQrymX9FlIrPOJpnUKz2erRsTCxtNbGws0/MTpMvROcAjfIXqbTjg1
BezL1e0CePDtKZkCQ+Kx7MJZ9SfNX5kXOkxMB4uvQlOM3vrnF9gwoWzQvE5O9fMH
qh3KfSfpYewchsjKhwQ6tzLvH/9OGyRoKXnGsa6qX5XDw0pq0ldKNoaCJVgbQUgI
l4iiLCEQb0RC8+1wEYZLkd52IM9LMfIfjuzmsiZk/+gPY0FfKJt+BeK9HIc6IBL+
Sjwbn5qwta4XJhmdJU9rqfjPjrsEEuuS7Fr7twku45eJ+qBOE7/3d268mClzj48v
1E6pNqFO08ZJbEmXwx/EVAcP3kpvAfagjZRaP7xi3L8MvnJbH2XKSIR2cPH6vnel
4GS3XH80CKK32u0O1kU96O2BWIWoSZU3DOumBGDyfnYvtz8uR1WNHV0Spkz+rrAa
FmWPLCbxfK5h1VrBhiXqg1+5NXZnZbuD4aMuafxPqKysdkEIZOP+seNzYprzTscT
ZW6oVyeHGTkTZkol/choDtO8uGgqpbetNsknFTCqsn9k3ZeDleMuXOW9xZHu7PRg
XuPzqhyZUQUhTHUTcr+4NL4Db2fhK5GDgowZasW+jW42cTxBV/gUwP+OEFQYMAzS
NJUlZwlthQVyvbAIih8e1eS6XTLdFgg96eWypOCFa1r/Y0v0qb2N/K/VXV+HMZP6
uias6ssQgpDaz6S0dmb6cUvo+9So7xXJf6JlP5xfw6coxx79kUWhs3BexRqPNKUA
P0dr/bJS53BlT1pixHoEj91o0rDJpaYZnO56s3iMx+gEpKiq0hpcQnQZ2JUsvFnQ
4LubjiA57dHTYh0mhejK+4gdH9ZXSTTYnfGhrxNeFPxDiytNG0R36i13b+Gs7qgX
ABqPws/pqe/MBNJleKUMFr9g7xrelbvGZ2/lnGYjch3FExYc0odJZIBabSflHmmD
G4wejvg117JnF+hl+njbAyw3WA36QqOoTTEL9WWdz84sT8C8lgtXWpir2v1tCXuR
5wCCtpt0S4kWHBiaAMFX94dlwBRp9BosU05LZLxeJykb9uKcUTAOXMlIDz35g/Af
ECcsaDpGdZjNO8pMC+9++2L+W0H9bP++2Qa5jye4gWthO9nwbxHG2+v3yUWrQkAK
oxOKgIiAcoRoV2PQAqdoYCapcnYm/XQjUZfLNgHSz/lwjbxEkjaNT2ERGGBvw+1i
ECoc59QeYVjW2Z722AyuTPMkkgISq3mQOl/c+kqE2sMRJWDOpItUtomHhXMz971x
//NnF3+6UWVLEq642h/Q35lG0zP8W+WRXQiXvu+/YMcVoFhpsFr43LtjvIcZwMPc
BARIUwPXHuE8dXIaQJR5aWJTGBBnlH0zGY8dsLKz0KY6H0q+Lp1xhxDNx9bni6nw
8EWr3FJ6tEn3yeBkEKG7oWG99PZbR+1pB0sEH0Fl2noDiyywrnAUSuH+HXruoTpw
FbkK5OmrT9GzIcnQohSJtR6+KZqJnN7yGpcqWgC7a3Dh7+z0V7mc28GO8g+QIe1Z
Z01ADQedhlHM9/bzn2COTokJqxoqTpydnt3b+qlOlF8xPPrE3iH2n5tIA7/GIJKz
/rikA3NtZziOXQ4v5JWtiVJKAQF6ViiXxcSRU9ta/Z8UDPjnBFlRFC6prHohEGQj
MRVj9nyRFTthPY1AZaRhpVKVdMGEh3xiy/7h6A839/n1axAj0PTD72B/WRJB6H1y
tA1QNccQsc+emr/Id5dOtmQHoxPcR7sDopHni+f603jEdcDjLPT2oGpfinDOGhS5
gcsZMA210S541X6HnjYIc8PeneTPhotxX+b4P6gwBogNLp1RktPMm543MysUoBTH
dOzqqEA8uPbhMCmYk5rW5tv6xO8aFbfwTTWU8zqc1bevYhO5/n0BQJwtUppvZghv
0+Y4PhSThdJF5Zk1WMCDL2KUhIa4vqoSPp7ypbtn/tUBeIO0JWjNgJNkrAm7CdKz
hlDP9uXZK7aY6vm066dJ5Mo8rp2o4FQC6p3WnFVq05K/2o2Gm4zABCiFj/8ZAcrR
keQAOjW9maJAdHcfb5rZEAPtk+n9dVreLVzww645GNM=
`protect END_PROTECTED
