`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2lS+8LOAvylEdEozFwWJGerV5ebwaKaWgliXxxIz3JK5G0Zc5djTyXq/rrd12lut
09uBcv3Z6X01Ek78gP4E4nxieoVcFdLNVHjQ+nEBw75DGdAX/CORXMQ/l0jPdWba
8pXpvBy1KyqHHIpTv2HbuIkgx5jA/N5zuZcjXTcFIH6GRw8/c3NWkaSoAXIz6AK2
NfY7903MXQLIZQWII+h7GUM3Aif19g54GdwaLtZ+IIBLObm4HkOSOaSRAfLz7mun
onusEP4BVbC2xY3UnbwuDs/n0ZSXtYoQHPYlENX9QACo4jh8mHFQ5FLsPE63Ug/I
Fi2J5kWPkpp+P7lbzGCZsYm6aYNHXL84Fsu9RfpSc3rqdt4w9NYB+2YncBs8MYkN
Z7Ny5JGOH9ZFgT5T5GN0Z8D3FPWWh67cmfW4T8QSx9YooJ4RYbthi17rSBmcQo4z
pf4Jr0IVxc98d9+0BMAFQ5zHOCVnsE9FzE4qxp1l/peFEd97uq45Exuh358EJvTi
kpOy5sm1qKAivEh4GpnaV/iU4kH4eaLtzmlx3NJCWOR42VCahztXo7FJuHZZk/cE
i31G5UG3fuMr/jiXBFyycTY5azZJj5PoQqBZneN8YOkhWS2fKnoUtfLfIDF7r+9W
O8yupjL9Va6AP29SLhwRx4aaZ+reb8u1YM4X4h4DqD9twgUVKOthi6frQ4EkA8k8
pvUkg4geSjg1uuG1Yk/bgcRRtejPQ8wTgS9Jc1k5NZC4v8mCE6ymlz6OR3f/ROTD
hr5Rle5MsxD8LNJLaebiYsYk4nNmocUB/MwOQVpruwvR+ViVVRS+YNvrsU+4221H
p2WLtFuLZM3deACm9e3OPMMSzuxrkpC7fpsbCBoMWX6dKmZQqKYOBGCBwxlV3KK/
SY6ja9LXGl0N8FIKfWg5cPqpGHmv8OKRB3DYaZkhNkLwLCMxlHO77eEobwmovxHW
9311yjWX0AbS6KYBSjCKFueHiaoBFGVp+YKO7dS8+BnVu8D5pJ+17Y4WzwZGCgnU
ziCZkIrxBiiUJsriyB0kOoJKUFSA1DhSvOXEsND4dDBFT1jRfPv2Tfneyy7y3lKb
lDi7lZMG1Y1t2Nb0kL7jcZeukQ0pwDJyt6KYapStiR/RSTmpwWg9mbyKSHhXCthf
+nEYqWCIHBq6zLAXbn7MKc8TLDrGo86yjvDEgZFKELfxsacMsZAwCO1LUS2zqTrN
c361eh4Bp0nu2KSYm/J8vlUH01GFstze60gS2NQRfKb9vwcj+5+Q1NYeSPOwvFm+
YYTk2o7DM17+yWb6AZhOcYrR3zcLfZVXnSUzByKdpkTTQW7TcDy0AH35LrYGX90Y
kIgVVc9pw8hvSSZOoGs0kr7wVpMyC956zyMkeVSNxniNZ7VcDgJXSlI29zqrseYc
3gkVyY/D9ZI/b3KPME46sMjQzNz/Vqhj/juuN9rAund88IJ8zGfTTYVlhk5r/qRn
oVF/QaO1rl/ghXHETDtwSefHf35XQx/xE43vj3NeAkfLVXQbghyow6FFuKYaplZJ
LsILf2DJjFZX13AOlXE9I64QXyaLXxDvV7MvwDoJ+gFzZ8OtksOgQLzuKMljsjIj
90q+5efp4TVoVpsCXjXLuXtyk+OJa5/iWrtSfLxn/QfJMPH/9KPX8iJQHaaalZZx
f9IHVAyUHXBXlcZHrHS0j0sS71gRNfqhJXBjRCRAs4WQ1nWUI1AyuH0l+Nngkg4S
arNpQG/9+COQJLeR6tPVogrOezj1sOJhucvT8ZGdwEt1hpKZF9twnfM7LFKda9EQ
gV/mJhJntc0fvk99w0OmRvZfAKDpEQlVnGUf4NtZl6jTkXWb2mieCYCcHRfB1W0W
aEUoWE9rwGlABbYQF8fnpFb2t0ILHyWkf12jscZln+x7YW23BsjoaCPnMwU82Zj3
79EyEd17tm4AKUkYWUDgfBfTi5iq/lJnHQUESDOE4GPSRXNWu6Z2wikS4ySCq74p
eYvIW4bY7hfMyFJJKDlKRO+k2yom/+xB18aUMbygmrE8elPZhuPbWfWKZUWtPt0I
m9px9vaOdmgHJjk5GIO9fndB2G1gGuV733b37ODnudfjJnHQXuCxewSW64pcHODK
9Yzxw+U6nd5b+/B3PbbCNihISNHO/i6SsoKK3wFQkMG8NT3fqXXmAeR+Cs8zPioA
tgE6edBUSYsi2iD2iAiACiXcaWSPElmCkuXI8lcXEXV9myZMkHWzeXY6BcVFaOD3
XT4l0ADG6DL/vW0NNGKne9qXlJtdeEVUfKfXltm7z1sqmYW9oOBrlKaVKSnGGCUN
9zekzooDImjxgzaRGhxqasGxly0ZeFfEISRjWFLJ//sEfn4efbMnOQ/mQAAnJZzI
NZoUdHH7De7mR7DpSKJtUkJ9oiNfCCw8FYVyU7TU4fEdneLU44DLg4plAJXYNdA5
mM4tedAo8XDiYVSeqfa7xPaihSqH7Nxrh6YFw3dexTh7sGlV/VesnTwMHjvvxMw0
iZ+6cz0Mc+h9aZfkVky95hsjLU7w/Cs0nH7d75O56pXqi2/Qkt+TYjzQHMg40euQ
YThXezxmdM7PHCF3z61AuNjLf3DKRKxJue351mPguvCosYA+7sY4Qr+gLR9YhYK0
4Wkp8J1yOeov7sihO6Na2O0CvbvAmgGJ4aG841tAHDcOb1HJrfEmLv4nLWHSJmCK
rGkCO0fuosZXCFFMSZZyCLIwvcKEWLpRH+bg/6ZTFyd0ZxEBa8NJBg0K1iZP6n6z
qsUwp0mzjltf8yrSyZnNYQ==
`protect END_PROTECTED
