`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VHiZVqaisD3o4McUkHtlAe7aw9bcFJDv3+R5oNRVfcsylfyyM4g46BdIIqsA6kWg
5vwPTmBUNCC4UhSAdhEi5To6Gha9oftaDGFNjiazoCu1Cp+FF/GJ/EH5jL4uQ4UN
Xhs5sJBWGS6N4M5Q9MJV93bY5XipK/wBSMI7avvYxacIV1mNJdnGODB6qb6x/skb
xN/T3TerY3qnIf1R/hhmmXwNEg2rwaGX7JrQncDqZFW9wAD3Wz5etIvs31JYLr+5
tW1F4KiyNo24B+Jj/+b8bto1TpGMUx3Aj5ILULXqtHDpmpBWf7D+pZiaalraj8UJ
hq9Lon/gqmGilZ3jIKzSUeA0n3UKCcUGGUU5rona2sHrzqBNL2ClF+LQBN1vW0J7
vvJHgaTu+vl60194nXpFc4rMs/gjvtjsFlOskvTml/8AzBER0qcjxfhjRr66nk1V
EPCx1ivzst2Ip9mmprffQLqEitD0VLrdcuW4b6F8zQVNSDvdt6ly3JCstctz3svi
DEL0To234HLM3y9B6jBQPx6GRuYJ76R+pUH6t2gR5byNHuWBQUG/+DaiWTTH2IwM
pWugaphrnOEaPpRHS0sqN0VhXFA+h3TdeTMP1oDncdQBrz8wyVpU/69s6Sl3r5TU
qOeu/6kLeQZbIdERHnfPzDBd7LtpjoW2vOBV6ROG5dD6BzTeaEmE5oIbO6bmEpTV
nLevAXQ4NGlBL9cCuDunQklgky2UPkukBtx+puPqEHIOGMhe9C4kVJScacjGRLyA
HdDFZ+a/OEglZ8ghYSoS2ENgdSLijIdGASDZ2aT8LnXQSTu8KCUieR/O3KpATFB8
bmMpmbq3Hg2IiGzYJp92KTPyzedhz1NEzoabvfJCPxXf5nKij1d8crHtzhjtFc7I
FcWhtDUZGNW5tdVADAQzn0W5TynuqD+fs1vhoOABMa8WAdioCMhtDr4JOH7NoZf5
nTr3cYl5f3lKciW63qtt0a5nXSCsuMzCrm+H4T4eIjkNwsvBS7YeuAtSKRTebFxs
TlcZm22k3/qXd/Dxt3VBKWNiwCGS6Z4uK5MqzjLtSuQD9cHl47drPGzkYFyEtFOx
cgvx/mPIPOseA4n+Cf4IUFl7esgvckTgi0PJ+kmAZaXqW2673lnkeL8bWg6Mvif8
4luFsD/RfuiHYJtvbwshYnWFHPmneNmFdCu+kh+JEnJ1Gd1MpfchH6lSSa/wxQuO
eIjrfHj5kTmte7eho999O2POynj0gUkYm4RyZKW39D1thS+aHfxQ8z3ZDiwtLEh9
IVq52jUW5lMFeyD22sqNYcra2tLtQ8tV6dCHvWmOgq9wcSg4bn/2WTNS9i9NYZF+
5IPXDHwxAp7tZ0DQ+LECP82SGLqKj86lQksJFFo5jiYnWBQqY9OkJZzHyE4f4CRM
VtUKUQCYfljdLcCV70dlJHhAuNv1J7RE2njsenvTdwvR/3WCq11DDMFBNxD/OHzh
qaD4vQ9ctEaLte7HHcQ4ZPfO53e2+v4aKehrh+ocBPfNzqkhN/Rolu4c0JOP0RnD
KESePjlxdGwvVc5MdgBG6WinphKtygo9s0MEd9OjOhCpvybz0/UtuYFVig2UGELG
`protect END_PROTECTED
