`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xD6HroDdIY92I87VvZYMsa6fnaR9OkW3gy2I8N3whIOkiqz1GYUmldRjTxUCwR71
AZuntjf7JBjeHXGk/R3oXpEjO4vujBbW/prqDpo0L3bdo0aZ6JfslsJ0cZQnCBg8
oIFmFIvUJ9u8/2LwQ+cTHdD+cd+aY9Q42FbmKqCHZ3CjpkmLxa5W/kUiwWBYb+cN
j904DBd8HjhIlvwu0c6bXkhVkoVvfd8MQI6NUB3B/B3NlaP2LEHhibFETMLc49rn
i3ACyzG7AKEjBGQeyyPfQHX4AjX+UrapvpEL6MYdT5/2d35qIPIK9WcBJ34GUF/j
Oj30iUKqjqYSb25VWFbo0EQ2+e/XRNDv6/69lYkwIzxjx4cf4YACG/RYOR+ZYi2t
kWUHAMlBpZ8FHjJMNFTcIT6qg0w4GKx55cGQSrguk9+ngbEWy+6gdih9DE22daqR
m7cMmFHBp6zzHena7Hi9GuhOvNXHEwDID0ku+aOLyZK46g2kGSWKlyDTOjf5ekB2
wCXp9gdjRluErUOZpRd/7St67gPgCvCVwNEYVYPEoR4fKkCXcEPgIC25DQ/Ug/kG
ijCc97eF3IeO29YzSTPdrw7+QS/Z2E0aYHQ8zzTnYNTHlvnz4DN7GhyJK3yhrvah
dWECqqYqyjeKZASbG2BEtVto479atum8zv8Mv7EiErvk58CvdjchB+840uCaQy1P
UEMx+/KEsqGW2GqthII4eA1ySXD5Waco+WEd+XxOOXFRcmD46VruE2JCy8Fg1YYo
d3KHPqYTJqKogKKu8w3ceLqucgMj9HJW8U5a+r985W9zH1Som9/7HDLqcUaqdrzx
1CnDQTBA9ROQE5YURyDhKmi4vPkAtpN/Nw0ebpDK6P42ZnTGFqi9oMgq74Kx+N+i
`protect END_PROTECTED
