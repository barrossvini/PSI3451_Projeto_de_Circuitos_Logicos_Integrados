`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wadkOrS615LI7MrVleV+gP0ClHI+Z2pDyMs3ndpqAw8JvRa65aXfpgpygnjcXaXu
lvNqW7409fpfDLUscfitIS8NQncIVC3X3CMlIFMVQ13QvhFrULwNM62ojBITjekm
iEjKCkCUhYQ2LSfCnXOWeQ/TrUjdZajeAWsYgHCPpcYaj45Ub22xEHjh+OjvbOjF
XijEmV+081SGzLPaSNQxoz6Cgqvl+SXZQEF4KYTXGN3Z9OD8tg7TDWw8E2P42LUf
olIUJjXTC6n7JDSU6PMQUf3EP6RWgewHLfBQ/ECJ+c35SBthVdCuzfDVkv3KDba9
6bPffN7ZnLIs+TfVudsTTKSTgP20S6Cds9TRqivywqwXxyZzjmbis5Nnm+M1+343
v//0d/oZlmNROSeQtjyDEeMYG5mRCgKyPg4/uR0ZLY6eud+cBL7K3jXmhAubI5Zj
2tSBNdCQiQ0DSbIq3m7hNmKA4oRM3CDC2UG7OSLQtpCUz+zrW3t0sgb7fyBnp2Md
th/JrKzO/D5EWRshKZNjqIahWkd+iR+t3kRZldLypR0ikwJBLR0qUUWawMBZoWJ9
/+CXd0EvM/9LZzD3saOe15mgK1ZzmXngwPZSKTfOkOr6vv39qIBhiU9d7EDoPV5c
rGW3S86kRvqhESnH7uy0EtAqjoDoocMOUJmxD3+h+aXuOa54HPrErxNsQRlZZ4En
lLMZPa5hYfytYZkJJTxKwUndPzg86zP5/zzxs8qXMsNjPFjGwVmibzFezV3oR6cX
ZNX4I+h99USOAatcZlPXD0J2rzuajE/WMTjaZI6iEhOIihdHNeSTp7gqDUYfPO96
`protect END_PROTECTED
