`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M4zXl4g2n117ll92gEA3eneKFhoYIp0QLlAS5i/LVR5QNXV4oCLEs0YARvpp6LM6
lpEq5W7SE8Va2jOnRUr7mjgImAh2ssSePjtFU9Mt42l3k6YJtBUcNhHp5Bk394cD
jfYGOZxUz8gpZ7Eo3/lZlea9JHjlfgGM4wBfUUV2pgzUo1Vpq6/zFQgr727gJjN1
YQuw4cROdWprnAfzDF0RpGluoGywAV3lRaJfOqb2QrcAjPx08hhZlmIfVvS5C/m8
oqYJA+vKBO6Br1Zc77BW+r3nYmdNbGFTD1lio6LbafvDgv8pmq46c53kUx1AaARm
/tljCHM4Kg5zZMaOvIZiDKjQJD1xDOh/XzJ0dPsZimQexnxHJyd7WYrHuUKOHGem
QZVXh6eBzDmSyuX5TOAKh6tY2+wbxd5HYSOrwFr/7FQlVXciR6Ad3HBoYFbBdIiF
4KBehJ+BooBp3bV/wm9ALt6CBCasVSniPHJMsBdX5BYG2YjU/H5MrCkqc2nuy8hC
7LZbxLP9l+CNkLt1u2lAgsY47Ki7ShCo77VrY2k/qLa2PVV/UXInmwS9yk6MeljW
o+5hMG+hAra+iS6OzueyAv9X7xCxVWIGNbK8WUvqUmAzgzXsWEsaay52Mer60y8H
OPecjFlX9NWyftmmGM2cdPADQdxyDGQGeD/horI8Soi24xBYSpXoYtwKoomwekWD
v2Pyx/u0y3Uku25f2qDQ6tV08HcpFJ4mQxW1+uPqh9ryiEya+G8h/7bYQI2zU60R
/Py7OKneDZDb8SwsVW+v18lF69D6tMCJDV3q5rwAkdfffXJ+jiPUYgipJ6xQ6Ph5
fFojw5p0mtxqYRjjykq/zYE/5cJZKabzIUY5gji5bU5WqXOOJaplJNP4N6Gm4Dvu
BS5HFXRV7VAIPkNnKj2fwL43aSNboxifMFC5rg+iYpA=
`protect END_PROTECTED
