`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ze1Tu+AS2xL2HtYwdamedlD39ELvaQMvukeBwYAq9AKaQrxZra8fDRnlHpSw96bS
PZH3osppA+9gx1dTv/T5B/cQuCbojoM5N+UKW1Y3TblRyTeWaxXHSwr2XCEQrY5G
CC4CNEOdRfqkMH+3Wd5LTtzEpcbrR14xcwn1eoGzRjwmdSxk3bSzp4pqJO16XJuP
M1ZMwTIbKU5belxWOgYe4+bHVo9erqv8SIgVrpAO0XdWP1F/Cl8AaycmUqMhqCmm
RLfH/jAPY05pipwwFmGPcwhKepfPxR/iMmgrmIdpPcwWn2jE9J0ndLuSEF7lV94X
dDfGFm3bLp8xroH0GqWA65ulW3y2oDN+Wy7MDfeXzdEpncicPswF56Yp3zboKrUy
2jGc+6C5YSpfF8vKh+kWcPdTCOrupy2fUOtmvYZ+5Q8uzbxEODzffy1+XvlBOT0p
9s4D9Sq6RyBQCwqWS7fU7/Yky5JUGEZfFj1HABdmxcRsqAF/eC1fbW+NjRLu65MB
dOWnAh7YVbpcqS47rIJjYu+PCKDo1c9EKeKWIYS3UjeWacGRAFjUb0Vrq0O54ZLk
O9lMk3YOcs8pXLMKCcCiRI7QYj5C3TkasrzQpHCTczwrAspdZOBoRGGC76f+8PCG
k1pL5yUZm1wlN2wICvnCyECyc4XxvWBomV8xGNLf7LXJ5gCieePZRzGHNLATdsPm
6OxSjf760wSHrjsM5yLV+45LICF00NdL/Wi9/g1r/d6R1opm1nYWKO8RxNzSchlg
FUnOVHaB+qSRzXTGUKw4Pw==
`protect END_PROTECTED
