`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iUhNYa3z7+NTWMyeg5Rqe+TRPMVB0GnPP569iPTmZOTESAb12OBHtozrpopBRWt1
iHKxTNk58IVD3Wnp6/Z3T9x+F4OKWHr2r09KgCoLyI/eURfMNNIZBYYh6PVDgUDY
KKxLaO51cz0zxcTAnZzClQlcGpxiTrDqsuCpkwCHziDIffZV0qwXRuH3BdlaIfTt
9enN4eoU3oXTVYVT62U64poFGBqgSgV5Xo2KvdalksLmACooka+cCayAntLrGBB1
rtiVxlTehxqFpqZfsGyT3+iNitd8mUxJEfIqtxn/cPibw9kPOaJiQalBLkr/q6mW
2C89KD4ZlZmj39upZM4z/rg1Pdwl71dE74WK6mLucfIfKxzlfn8NMY2Q7AL47KTK
oV53+RNfNfqwB9p/oGgFKT9zCgfQIvHSD2NV7okN3m9gA8I0cbrAepNHTd2cvbPP
UnrFoOIfw58ba7RNihan+juhKMd7On7kzfJxvwAJnLPJSXQdTSCzPpVsECEoAg4J
hxCnYAxoqxR/ILplG48m1DZ9p5QyrcQyGNHPoNquIxNC0MRznfAI3rDusNQ3m8hm
4ThPfiU47HSPPTVDlXn6ESOHlknZukER9YrkKodqqOz/2ZAbhXd5k2B3Cq1kZ2O8
qfBckK1RcCnNyJcobxs0yYwSQE5HycKoOQGg6MlLEOmT+4iEZybLAbI2Wzj5SARC
hHK6/7X+2fpJVGe2rKuY30iNAg3tFd0bgLw0lx0g1m4Vh/RH2tOGlvn/Mc+r9x4m
KeZZmA+9GcNLowLt7MozpZWCuT2YmCkhsyo14WQuwQz1GZpSTiHCr8FBeTIJFe8t
92yqe1BZiIUVrVqxDIDJFct8rB8DZVDnsYj91/QHfPvCX3k4B876J3t44XB1a1lP
J+kSAKqRorwqYRzsZMl7qbXpKCVa1/Sj23fZhZjvQt3TbyB/gC86cQ9RJwNTfPk9
kZxtGiYUH1I5uT0Te134DDcbjVMTzHWXzJga31mQa62n5kLSprHAH4jSxOCXvYbo
EoOq8u9M4eWG8ExZHOoUIBTmACxdUkJpISv+ktApvkYtm33yKTS93rDl2DDdniYO
LQR/mvwu+qrvddU/17R2BJ7ZWT+gLwt26cnP6kga98lC7ZPyqrAkLwy9MVWmqnW7
Fc1eXb+UMw7KTkrutr/HwI9jL6zT439sGy4aLK5HWPS44cBq3hxfwZlZ/0dx2Mlo
pdk+5WXBgA4ajicRNf+yYuTSH9Owc2nzZMTPMOXEZyXz+KGkt7p2RhT6U4uZ7xoE
+3j/zC/6q9PKE1grCzq0w5YQgT9oQgxN111Wpq5KKDp1mcpqEZTIZDxgKIXN0q99
7i8vcEesBsoDnOewjRZkOMEYlQyHmiEjBN373JYY1p7DEW6ahCs+V6VCJzwItE+8
MQHkZoKcZoLh53l3PCLRU93+p0G2wqJGIialWvlVJQySQWvbOewVesHqrSYRBGed
K4e05zmyNMZ1XxQeyipfVb/JEySQzYur2bRrY5sAWM9GCJdSxBNiphVeZiKvqpUg
ydw9nMw4j9ZPNaO+kJfXsF2zqzqx5LdFQKo4iL6jX9tVlO+NWmF5kmSmxfHIar9Q
+WcsS6w6Aa0ADnBpi4GudU5SPMD4t2aNXzevREphubXZ2yLUjxAStwbYHWroanTt
/5RDLbAqk21vIQFIYranNPIjsm6LVxfxZS0yFjLRmDaA2y+yQ+OxAcfiPalNSxIM
jDdaaoU+Dcaj1iipDcw5OlIz4ZVB0jsUmYn/2pd+HLT+OmgX+JZv9aVpmaWA8dYC
PjYFoAWtWQBwkAYhC646MiCm4jTJAiw8CbmaiBEBVyFuZoSG8Xqt8H5l/vw7sHhr
V646kw/IwJ5L1LZF+MXt+VXamBeVe4o2tCJCcDD9b6YryfJjDYIoAnc7yAgP/iC3
Z87jJ3wnu5qnlj/2jdjc5cNqlLNp+r1ltS80BV1ahlBIjguMvKb/Tuhv7HaLmIw8
xb7ATN6i8LJ+KwTKYnzZMuDk5wjutRI8DvJVrnnkQPO53ToaG26yWEXv4Pe0iDLA
CJEPgWRQGP8ffkX8qqI6jAa2NBPDxeGeLw8cSK5AZQWd3dT6YJNmy2e4wQNe1801
RYngD+Yqk026+KGuEDVTkhito9AalsQMVZsTgSOX54Ujx2HM3x7W/C2Cq+i/VzKM
Qfk5eAc5vE7oRD/ReDcLn2iSFEV/pnT92AOqaMdV5LGrER1w63+bCdwWrw66ZiI8
RNuRnUtUnscysLbIWPF7F7k92lTuzyg807M1uzd3VQ1Vi2ouNd3aG2m+xSDelm+2
ejlOT9528mg+lAbEvW2+8YkxezyHTQT65SMBICzkq9amds2d0OYJybgvgL8diTXK
J+cRNURDTWAa/rQrhYULrHQ+Inq5l5//y3wZU79fTmJTV+ofHF1hhT1rxvIObTdt
s6kzOfZAZWr/Ha6/E+Byv5NCxKjIOVSA3aBERTdDNOW3dJaiD7l7FrlmcAhP00HL
+AawtU3gYp3d9yY6804Vm2VthqhNJbp/vgLcwrD5gRVTmAkobMBxuw6EI/H4n4lU
nXJV9GNYOPcMFtvN+nVEIj0/oWwLyNTybpIHLy6PQb1cJR4kDTPRsl73BaaxMxq0
bHi6VnFJdYjNkJjl/xa+UbCUUAAhf/NsI4H6jhwKqYdzBD248EgZXKKJtp8zqRlo
kI8Gfz419Im5Ejl5yXXqFfJIv0000vioutPfrpsrcgYeWAPxawejplGBUbMIfAMw
IkTWso0hT3FuAnYIvQlz1fK88DIUZ8ypzuA6uohdUnWMuY5W3sQB2H5RTh5+STXV
R3K8mRcahzBjdp3XntPWhSDW9J0JNbwc3rAuemSkLuoU8SQhx4ohnALTA1cRwc5N
w2InSUdJtoWalRwax6soiHV1oe0NjnPK60Y5XnxkL2tgEi04v5qiS37veQlyMhDV
PVi/aCgQ6/cVUWhvHZeQq39joSn4njCGCzRZTr8XLzu7esBeDmGlknwZKmZD9fyl
fDhd54GbIXLqcqqxkQPw8okItW8wUZdqEEs3uY95AokTqHshb5eXAU9h8SOfz/iI
tWoHTDPthR7Y7tnsiZJtR6u1IWNcgbTfaE/8wbAgHneOc7xKgKblYMQJNHdyTNz5
Gz+Rv7ilDgnbUsZ+qFGmo/RX7VdHRaWds1pGJyUJ7P+lrUkyGXbVUmwNEI16i93c
kHGPCjz/t2tiN5B8BJyAcJCiPGR795L+AdKjzyv5WmxedNtiiy/AbNvgfljPbOJb
ukfUS3SuOky8ACP89eE9NNH3AWJKh4NfWtYJ4sKTOMjOD1co1eg/WicrEiwNxFel
wqdgUbQD9FZWnpgGeGR0CsBz9jkc13uwYivmKJHfcud1BRHVU/+a6D0J7F79wpuo
fgVPKsHiSaJkhM2HvpEWKHxAOh58eqXZgU/Oz0GgemSVUlRKwYNHYe9wiUzh8Sta
GGrP+uukw3iiL5JnrbFEHO7WNTfRUzdpIR4KcHHMTN0C6AkaR2N47KFpBAW4XcgR
2t5lsFQ/gvu0nX3qw72W3K7QzmOInAe0J0wtQX35wYA1CQpWgi14xxyxAHkDYLuc
3IR1W5Czuy+ZYTtLiFSJr/ROJoQxE/XpQc6QqCu7yimDypk9GMHyQihYTMF7T6eu
tcVV/oOvuv/s3VW8wGl5q71wn3PAGAtPxRaMn161238910gcATkdOQtsYA2AFJlH
mL8Bcl6GSMjVsH0H7gMPrMR8aadULakYVBlChM2JutuPcCTJvG5c56oHS1Su0RhK
pVoyTlDQjN+eo4oj1as2gJRL4CwI0WLTDjksDSwmzAdOeYPDBtYLACHn8CZSb+ue
gcq2PBU1dxLA4QpCZxXUg2JwXOHhilPYuhUQ+fGVJOuwMYg6ErxlIFrgST46E8I6
CXrmA9YRg9BtZ2IWmonOXL72vHJHLz5G2vJNcBVRUni7fGKK8tMazPW7fFhh5K3j
q5ZFjg+VT2kWo/FUpkYhuJLKTC5GDsrE6+xeHjF/JYCvCblGLFCkcVc40G1Ibbht
4z/tU+B/cgToISUMiNOWAeykfieILLil8SdnamP5qbQL5rPB99mZ+aX3FsKUFwPu
BWe+FZbMzsA2KOQLby4qTvroGruxoco49Qthtv4mQjF6sACRr4fKE6NEIYocdgMu
nyBEOOhgnyiXH8ERH/oxoNclCDYy2jarTLlN97X1GGRknbr2dhXYKfsDdMx2uMoX
mJpttCKZWOrIFSihj/lMcnCYBs5Z4HsGmpF2I/t+tHZdsIKTU9bY69KqukRFG5Ks
CnvkAcFZhb7fNS9TcvJtWlgFQXxxeIJfd8GdIKCgyvyS2VkoikOXHgpOe0Blz2Xw
3tvRxmEgar8j4nWxtqnqFCgO0DrqJHViLE6P7tFgW0qxpRLqa8i2P7Au1apWnaVC
e41l2AC99IVbic+VUiN5nTN1MhkTi/xuoFyQER9cINcqVKi/CdCZKVck9+zUzlDM
PXFPbjCYgDxPn4Fw6j3RqFGgNJ8UBIpFEv0Mg7cUV/D7TdLMozqh9eQj1M9IzwIv
JuPG/8Y0+kj0ixfmywesSsYruTZ/KjKlVJI28hkAsiFkheTA+/5gbRRfjNN3HPtw
wkC6GZu2pGo+kGbxorIGiYdvAO+63XsNJz65VUJyAMZ9L+qAA4fe/dy6KRFO1Izs
GWsr46lExBPRn9Yc4W4GTK5OAaQtbWXjXduM35kNlhAdZDWqpt3u0L+N9nkBgPRe
8sXN1JPo4O7VNDxk7jd9oHzZYmWyMjSenlZ7awu86VIXzU3QiQ7GAKO3Gcb3eC2c
fQ2cklIQ/H4JC4B8ssB6ERpDDYnZdpnfg0HDEaaoD7P/YXVS93O+UhBb305EUOyo
gNtqVsZj/3aBC8LdvhHCYDmtO6PwF4pqlFI2aA46HbfcpJboKWCqQXtoC6xCCKfA
Fx4/qedRfBjNq7rugUxqCYVOCrfwHYce1QJ+8P+sO254E6GseNgqxlMO9XUkBGfT
kyv2oG6aunrUSvjwKjuFvEWCoHe4MBMYzet47PxILeR4bYhEiMVy4pJEybJ0LHX0
Yjxpyqlvc/ExlxYFY4gNpDU52OftYNZ8ZOFfnlLUzam0+o53sAk5PYevDSSYZ2Rv
EXZ6qd0ctC+FibHsYfuqGP8yxlzwkj8gq/k1zvXblwFY1pG0UmeF+cDterS3pSvj
/wCMxmFQItamVCwsBiKZD9wR7sky0EefQT09ZBxsFbA88ud+KIWr30Ao2+WoK7oa
Wg7IMazinTPB8YL2UGD+tYLRU2wA41L/E08yLIxgiS3B673dtMB5D36a4NylKw+8
YdWj1GykvotJT41BtRsdaBnFGJjHIDh8YH18xNMe1YGujPj+dAN24mtSCPt+7vbN
2/6+g1swROKJdQAtOMhc4CqeA8u4lMbx9QJDWb0MQET1iJgFQXliofTubbKcb5eJ
/AATJhKpAfYUwhCuUtdZ2/4c2vf4/l5FFWxSkBvslYNI3ZtPledqhzgZ3CGiJIMN
wlPv+Cy0vkoCKm5Hm0pAEbdjVKDTgS2f2pEOm7OzupvEvx0CZeQe5hkh9us6gytd
aeyth3gZ+K787k0G+t8uPUyFOblo8K0vbclmZgRPHkj+yq6AjTYFqtPj4atD7q2W
RV5c4ZeMWhxl6ne5LIbr+3nGyCHngHh7xvVFWYPGPQKtfWifL746Wl48VRVRQ53j
1YYw2iByPemLgtT/Esg7nsL9d550GcONeT94yiTeoCGDSI7YD80R1Hf6/SfIAejo
IeRCQ9ObeApLKGmLvrHGBaXeAA2yTp5veLTtv+xgDcpdw7dNE+K+aeuCNmRholTu
mXQvvWSxpJGoyF+yDrscXT8+qejKqnLMmwxo9zI56Y92mtlbnwpBHtakegHoosG2
kmf8RCef8hJjTAH3dgdU+W/6KS38kgyw3H6G4DX6s/0ZgSi/ST2fAvhae3zNk/j6
Rv9EKPsoPahsENAtKfLp8raDG4cB3fHG45+MoFDhbtvZiiwis42ZdYDsSI2QP50B
7tcBAfoUi/3Ngg9Wsz0jlXE/NhSYjipw377+gyxVMEfKW+d08O5T7hTtqEDi13Pq
3OEGHIO/ydvz99NGm1E1wQV2OnoOTC/yKWh5iLEOwM2uDa44tAB/8o3g6yMlqaKO
jK5fzBZSlJQSywPhVue4MJ540FRX/bt5tKt0s8Xn7Rwns9Mkx/jBBQfTbsmftBYf
bm87tyvxhfa6eR/OVJ9N+VAywgR2RK7FfQrLM6cQ2dMV1477Bi6SonialUwGkb00
q0Go8Y7NtrdKiuZ+g6H6GLHkm71KCvpBdlBPubwFkikSDyouFcUPObKVywzrw5DC
HI99mADoL6Q56lKuXosWT5+//jQ+0AWEi8VS6NcSWUKZAD3tdYVM+xvRYCftBgqa
2y11BDrQbjJg6OX7DRIDqjnr5UAztdIfQU+SCdOriacSuLzlKrXDPwfQO0PqpkCq
TwzBYgG0koLaqBVXZ9MOME6WGW7fbIZx3WYmt026ihS7WuW8oKpQY/KezXypg2yC
4ssveKl/FcqYKsvRWVz8dO4PsTIm2dqREWrd+OFyPiTuWTMAkmVVilu5vfIKFzS9
GmxOWEgyWMQH3gCAuWFT8Xd0NyVGN+X4a1YqK8c/2VULtYH/6yaTb/SuDjsWo6GT
U+ceDLk4OGBuTiw9Gk3pK0t+dstwMIAGwdXnWoH9VxsButU5CtITZmngtBgovsvP
OuQmZ7NRBfvx5NVNHxi91w8Kp6QuIloy25n4OfqO9PQ8cGNYIUg+fQHgB3WguZxo
0785Kg/8tQEUVBi9L9pyWUvaqwvwIDOrCUomL0cqLAjdqs1VDSrTuzeZGPiHnbcv
TKlqwExRXYp91lWuqwBFXTihUd+KMx//5tPNCTOdE1RxmSsYTo5xvmqFAJ+3VEwp
cqO9SZrCWhacUBjqmtsIJQna+GaG27yH+IUErvmPQAmcPvqNA9zA8jIv35ACEuty
I0tU92hZQOnYthblUJdPqIp+O9AG1w9wtHw6Pwt+SaL0WqkSavyE1UhtRnCEBqe/
vQT4vUO/POVr9CO+EEeC63dpzu5R0Wn1mKwcFXgQacDlq2E8qpHQsRvXWRmNEDjD
yyHT3Azasi8PcCBOKHnc8wcGR0x6lIGMOeXeEKDt49/63Vo3ztmq7gG0RX/OObfW
dxdfBXle43Bb1OCv0tOQ2Ec3oEY0dGXvilntUWLqBGO5yr+Yit5Eki0ipJbFpw7T
nDrwpokNND0lF+pl3MbhS55RuxRvyrXeYARV3VmGVqQ+bRhSuGND3MchPJu0W0U2
eXxD+7O+z4Utll4v3nQbIqawB5Xs2xAJS83iMkcgcN8cz+M9o4EWpDTlzucYan4H
p2cEXyC3xuyImPjCWkReWXBWfZD/ah9OML+LtXwPsG7JVBL3crDekedzpuAMLVFT
GjD2wKLAhrTHz58Yj0qDaUjHv6uDzf6ygN/nAX209iqj0hgPgx2qm13vPP6RpqzC
kmOG1qlZtRd0RN0iCKA3xjjoU/X1NX7yi/Q/K/t1kbCa86Ea/jEYCZ7uSIrFul9y
tGtwCh1KuTUiDpjn6OXC0gLxId7UvkQuUbhAZ9/Hb+Nf4/Yl1DBs8Scv4uu0scVa
ZkHcexmd6lT4Jhw61w+VwXVL2kTsj9HfSphv4xHzz1X/xp3kR8vX9iZ8GafKSPJN
j8o3Lbdi9H+ks0gps/jbWckZnyuKs3fDL1as/66co1U7I4qHe9JccWFPSrd93UP+
qfgcGnsWThchGs9yTrsmckA/9uf4X84USY/Oc9o/1+0+VGM9mQMfMV0RhWZegYBz
uSHuvPMIlrmmmqgxd5L62N9eNR66MShNQwW2agFkkj+DYGyGzl1OzCai4lG8vEFR
/KyaSnwxxO90TIp+SQ6fUv/AatcEtknDOPZ0v/pN9kDkuNCjss8ugtaAPuzU1sIh
PF6Jqahk47jfxZaLW26WzHDdAus5WX/S3aUiAgoNXmiFjiAFc2RvWUgExdYra5vs
3HRvMqcesKEb3g1XPbvot/TWN4KGYIziFStu7IHOZioTqIseZZbSZjCriFATa54S
dEeomVYqQOZEqcP6roBLpyzv730heJfPngBkE16G6k+pNCUtxG+6faUPsHPk0B5x
nnJbyq3BfvV0z8cdZTFb2T8uDTefusXXaWrh3Yx6aFgyFWuhjSNdasS7rzZHzv5y
x/y5seLddN/Iq6sSonR8S2VhtBTZS5+8+zVMYJqqISEE6cwEpkLaKk6LwR06uk6/
r1Y8Sswhn4gfjeblIGv1SZOwGpsknBFeDNkv7SU4kn/+kh3/luPu34eEpv/Gk4By
2uWc8tPnaJjydtD3k6R0WLIGFw4BaoabGDGrSvev1dgRv7KzXfDhCaXdPuJz8YLL
7hJuwXEnEhAeP9eOkVM6Muwzk+XhrZcKXHQSmimypXGWDa7Yb2JZOjEOk6gyGIHS
I02o29EloSW7xgUiOtRKdbS7wlLJlHIldLojWvUJJMPp6WxGJc9x6nPRp3eV+mNe
WbN5NI5HPsa9qcKpDZ0WUutGl1DPaOSynMWfkTFlE3Df+JXCPXHomoyl8C2qrfEm
fUF+Ea7kj9DWQGZZ6cyzSQ1elcCQG85damHuXDGF2GbtJg672K5uqVHlL28qPT8v
XiA3YqhEIdN6kLycR145Xm1uBsT9cKu2KFdEmnHMfGv0rCGCuS8luZtu+ehK1Mh+
A9FAKvWhbgxRXl5YItDmTTjw669WCzTsP8UleMkDVg/ze6GKyapzm4DlfoWBtbmf
QyNbiv2ZhcQemjmPkKn1CQJc8Dz/U1Kd/Qpdu6CVJkHkeut7Q6WwhLiEZUZacnGm
OEJIxpt/LFtke91l5h13Oll3RrNYOq/VYiT6VEvn1BaX0nTwwOa7l2pr7XaEyvTM
h2aHOMxwTg94zjoZzFkvJpwv+/WQe6I5bX66z98GkxjVBi4MXND/eCGRfqsPskTn
hUKt0/sODb+1WYplX8JKhqpAXNSUXcyfs6aH5as0urxiuK9zHOFR9AU0mSx5/abG
F01K3wILjygEIZc3JtqqwML2Zl97HxFe9L62NOBdhc7F9yTV0a2qMKV68HQrcgXH
yF+FGdKiLJisyqwDX93LGkOrKL0gw5Ie5zbwPTx69dm1aDQuFRi7kKV3iXf48Xxp
muQhV7Zl0CN/hHGArRxWLGU4IhGFqrFPwp48dy/OysD9aR9MJAr+TL6qodqMCB/G
sODhXii6HgdnhzhrTcXbOPHyBJpuCrSmz6vaChisHIu/WMwVgYLJjTrBwe2/wowH
aJUTWpvzH7dRcWa8mKYPpG3wx1eWrEUamsaPstlIFKjuwkX/2Q8uUL5MHVRFO90E
Z3ncQT6MlYB7PLomfHtHVm1raZ8s63hkJdrkVXipyiyIXdq9pfSXnqn2HTb1G9gx
5sG/7NWm61xN0WahmPCreUWSzcjpuuTe6QvgOE5aVGd0PN+Aar3sGgHRjXR8bLNr
pNv2UEWISBof+tgZ1HZ6zENf4YH0/LPaJdg4sdwDtqYqku7HvIRCwDJTVHPRfUa8
2hKkrlq/ae8eymUyJcU+JO1mfzrgGMSxQaEFTAIMFM5AlCumxXb6dgWYz3SV0HHA
af3itDSmdwBCUEeCApMFLJBrABTqEkEehCOO+XgLNWkdMUy6SahZ0JUEffU8gIkk
BZBOOvSzC+CNcVMuYz8rInzzoT2nGvyvMKsDhtqbobhV3K/ce/KQl6FChUbdXwGu
9hpBUvSOZZCtGTU95wfFCxNMr4I106zdCvdXmWgdtF1ENacCSzsS2DHhCPnlhKXq
p6CPbQM5HXykLh4ca0YftBnqa28P8ZtsB7aCRI3OLOSjDPJErOH70cqv3F284sRr
03dBQ2jYmfLOgCCbxqB19pSWNfohytE15RlhUqNHTkdPiKZHAvWremA9uF1gezfq
w5n44s2MdS7sibwCT4Oi5KOH4qKDruLYGoAFRKFRRDE3xje8suHlv4aO8xTFfDcJ
BsV5Bb6sNqHMPDpkBSoozdngOVGyWa/yyXRDW4jVLlbq1VVg9yzrDPUy2d8kiDAF
F8//3ThJsryEB5R8OpmxngjL0YIYSkUlprVd0zO0Xlh95oe1cswOuBtyn49hvB9i
VGY9j2IXmwDwVYJ7kga679sndMmDHMxU+WSCnAm0L2U3xbIQOD/5OIOua8SObxI9
LlezdXz4lNHiClXsdkJyI8vyJe+pz1b/1wpzM5pz5MJhb8DIDnnFy3E725tjfm9M
2SUbWD3uhwtUhok66pTfaae6YX7YobB4rnLjAxOvUo66uhMxtxQkgT8SkHPmd4Ia
j7UfmqA0TdkFV640BmiWdV8miA51XBfsxLtP/HcoE8sd9PYa4k1UcXmTt2eXsaUa
8WiWGiGm2MAe7VHuOLtY7NM3ZMD4xEgeIJgXkU/HM1wbtElviQVcE3oD5NNzt8Pg
GUqvhAAWXAisqLx+a0IGpEoz4emPBAw9acAs7S0y3IhWPNKhPVwQ9dJWUxmSci21
S+NfaLysKHfwdwjDKZ24eSnPuS4h9MvxcA7rFI5ff4r/xErhG+b8h/zimitTUZ15
IoVeJhIEuldTwewI/2xVjlV8++bmOyLPdzKUYYl/4m5B2V3q9LF7b4BaZVhzVA8J
2XbqERxMXo7GymldfP7uhCcv2M6b0bSqDF21zENJfhyky8BfuaYzCS2G7amot9ct
pr7bPddXoGFKJlfhVn7L+lYtCIc8DwZzqOaZ2gh0VZSWDjs3JaMu2IzY1e+taHTN
bAd7MDD0Q0bbizgL0OOrugvYaaMIIbYT3h97gH19bDan6VY86Kux/WSJaRoBf2Pq
wQyz5JVXkuokGdda0oR4p4p/Z43LQ4vkQcWgsUD7HqP0SAhwfBtul63C0iacQBHu
EP48HCCm1S4wgVWfnNazUfeQ6swbj+EISZwkXdnziaRblb6hgAHpGR7Dg/7vzav+
F41GrUnbiZQEjtgF7PORVofa1u7+TSGdNCgCj02w1zq6nILAmRlmYHc+A3UhGfGE
s14lvz1RchbkoYFeli96BJhgDnGGT0OjMIfYpesm+tXWZZ9qNGWz6svk/jfj7Oig
SlgWeOUvcdbE9MEGzaA19RuZMUAq0ciRYxlti+5jYt5JFnc+QiLUajvi5SfIbHt+
ZhLxrQIzSHw5O7WVzxhmMdX9HTTeL7DsMfHSW/2w0yJ4lIqGLgut6lwWMwgffhiY
l9apFQ1hIUoVS4WPi3YKvRJbgNb8IS3fWtQ19zf8u0UnaGLsjaEfrTb53AGujLwL
DMdGxt/8DplPPanr4Fr0rEHcX59aDlhBQgqqIrfxi1dTa1v2yTv+mhgBtuvgdkjq
t9JEbh4h6RzLSPge4o2pjSuCbTXbjGzO0m/lpvC6AThPLMDKo4V1Pb2DNHVBnfBv
qLEAxlmx3fh1p+G2YP0EUDzabU34pUIkKNX3A3f2VLAUX8HmX3CMAGWsgxQc4HJw
FhWy3UGbAhdEeWng8MhoPInkMmTtDadT4lo44YUWfe63yN/NfL3cesh6K/Z+0J25
j79JyHwBPxcb0WNsqVvxmhyb3YDp3MEx0SnGA5IlhCVFVDLrmZK3Yvct1yAXnm8G
cDVLxCviM7uVn2GQnZArmGCaOe1hh7JiYkn+ynFfGhOR0Krd2O1jHbRm6VsToH6K
FaFPtsx3Dhhs+OROzVwMPQF1/nsQRtmDb6SYgcHM5CGr74CCQlOrb2Pk28i7uvk/
kz6c3dOcsMVQRLqSlleenQO3ti5SNA7KK0IyVDpfNpY5+v7vw3Q3zx2kgZyXhReT
cTl1X6mJ02uxVToJqdCf08tIVGA5SZgb9PwK7yhEWMPv+tjjQTDOD7CQ6a9xd+vj
2JhIWLjlsw7lJR4LayjlF8WIYYKby3Y/SfQH82f7eNORxAJ4mJ1TVh20/14mY14Y
yyC70dMvElf+0wDw+ZDUfahx5kW5UnoLDPE71EQwR+lxTQVVQH4S+b0fdXFmoGKN
dI2tM6NYvJfK08gh5gxyKySWUCuDdjItacBz4RDE0O3JjUB2kXIumk99fnrTnCSB
3xsNH/g1Ohg+6UGyPJ0HTyrkinWR6henUEyvrFNgWvsNT2l+5o8j+W0Z3sY23Q0r
uYawcRUrOI8QZYpJTwS1OtukJJ8FrA/Hw1UigM7EPtG9ojHd4moxTmbMGAAfnIhe
YwjrMqVko8JeVRO9KMpH2iJeLfKSqXUXxfIoujeYjPP2NZoWOIhqFMTlCFDarpaz
GUPH5bgUZyrwCIc2m0sORk/yiiqxeu1V/QrIfL2FxWIpzl8kzdxG+iCteWoHQpkq
7euzhfDLlHEItNK5DOSOqxUj2TcaYvvyj9Wjj4/FYn0xId65MgXhMq+gdNb3cxPn
AbL2+2CECEs3t5UsikhEeIocz6AB3j5Vx7qoih/GkioarEqtb4DRXKbymD2X99wQ
KnS2Y29iDgd/TajtSdRYpMIC3ntZGVOrTwy7hOZT1/RtHQ1Cgukg/7MVEAvD1eFd
64w696Ss46ynA8UTyAo4OAe9saae641yZ/HZC1WzrYqRQ8NJRBnIl57QJO8uY0YZ
lLrulWaXOyElInzL/IkpKiV4R6WvCfBbJyINepJ9VjPGmyj+SvsYazVsbwKzK/FQ
0ohHD8Mo4w5yIuTV3iem+NG+3MaDDKPDMK8BX//vdFfn/fV8spg7YY/2qkUNAj/m
VAPTQJisqtNElphNn8wWZncVRYP+Oto6oY+Cf/vztMfoinmihEhO9Jdbond2Hnfy
KlTz05v/wbryk2YPCnXQ0b77vKdh/BJNJvVER/CQG+7TubtRCde46WUyvvkl4nep
Egp/Y47wrGNlVV88IJ3l2GM8oVv52Wu9oWqHBO4Oc0MJytp5pfsTjK8AcKhiGv23
o5eQCKuSSdhVPtzgpAUbd9xFd6xGuezuZgusK4rcCZEu84mELObPki2z4OKGP86h
fPPlwaEzyjmsyxWKruXCIdvOB4jvh05+q8QSQux7+n7Tzo88CbMH1IFmB9VBZYrl
LvBXSgCWT+RxMHqZyWdhOMSAUnMDEaLPmuTexhmrBWGwTnI8m4Q1upejcv776DW+
LfFO+vIOXL6xH6/pMdwbD8jX8gp0qwHPBQa1cx2ayzaD+1xAbvPl57lBmgSzAFXu
BpNSUFxcTTe+X+jHYkHZ/dtMtWrS98rIhnPwcBqfxZVinJc2CDL7VQEB6osCZyYq
LIxs1IABW82BGk0ESigAekCP04x+twdzVWbvgqpP0Jq65MBcGJ3XCPk7D2zkSKqe
MEPW203Q0Yv9wN/hOmcws34NEnvLd74CorIEiQ+kD5frYY0zHEVneGQaf+usYqxB
MCTpGavwzLBWli2AsPc0lviTVsE5YZj4lKOZHwBdXYKAs7n2tZvkPVcWELwHgjzj
9IMsCZ3dD0pb9maZcM7Ugd5eoDt4VgXnGgm1CuG/MmFVTj93fEQ+lp/aK3RvooUZ
VrhKSe6UUSK4r1yGStbOVO648ZvtiJwavjTnii4xiFSsCgqYgWXxInAG1Kn/zc3J
8psY4gA5V5hsVfQczX7XKTTAfz8TAwEBw98ORiKPN0Fm/v/v63am1wP3CZL2E6+w
VZ1Eh5uHQAKlJfMNKGmqx3Zt3GHQ0qrucYGA/oOyWPG7OsztLlnuyvkQ5c+tcPJE
zRH7Tmg9ft8acL78H5XCF1MeDFzhzk2BToNw70Xp2wINO76mlqq6J8Xckgy8CaJ6
35whiL63HyUjPhZ8iqstnr8B/KPeGYvdAlnp1te51Y7D3LR60AuQn3Lf843FzmeS
51URwhM8AuEwKGWvvSBOeAi/jBsEkP5PWzLQBERGYJVKYs2m95tHfzrxO9wFwMbU
YCA4IHPfQf6+a3nfKe84oX0Ntnj/F4oNdRTELwrcjIVW0YyyMRyARMOhWNNFv83m
47gry8wxl+sm08i+0yV8gQSo2R5/KkI5CQAMmNUnuw9BrX9QhbHj8YsH8DTVuSwG
DtpcBSpwQi++9QJ1bJP8CgTafGXcXab2YqKFIE4o3zOWawy8mO5x+8Iny7hWIzXt
PIRn0+uYkbo26Y958/Kdo0RixZaKKpw8AnYAh6Jwik4R0R0k8uYPCXstANbSfUb3
h5mRl8vVtZaBsXRBHV2qxuFSeDyiVzq7UXeoymU3NltLTghlgxW3GkH4ZU5gLEDX
dATU/1Zyf4TYzhAHPu6EeLoik5iyWaGGhKwUKrG1k5yDe0bIjZoUBZB/P8EgXri+
So1nCnVPYiLPRbBogZnk9hz2laLICEjAAmX8UIqFcU7O+4zZiobFsGvp+vSqf7Lj
96YNNlOc8EBGf8GKVcVJQEP3bBu/+Ch2To9HiRUGcR6/fFbexbxTiJd3/yW0ctHY
R/A/ZlE8dyFNEQCO4XP+1pJRvFeIjshIiIPqJBPHE0eaMs8vMSj5UFqeULlmt0W3
TzvLBRGYAubSO8AxzB0ckb2fZnmLwD3VCtWq0g7gLBc42YIsYPGe5BdCHUy4emf+
saTiPeiEs3K3ySoCMjmpZAVGvCDrUrbgvGWrF9wJ5g23PK4VAXi3BlU8wuT3esDu
4Vzl2d8w/cgfGZeeZP1fWqRs8GeGImq47qJFJgGaHPa0XztojavUWTvRkCNLzXGc
6ENvI2hbL3RN42RO3fBMnrKU8iUPG5+WS4Jy5cinCTO/s34crX9FZAQsdZ8GrMuc
1UhjcKO0KYEq7XGvQ7csvPsrXHxHUaud2cHawPZNuJaplQT0+FCe+3eipDSW6eUP
Npcjk7scWym61r529syaJBwhnLHMxLNOVS+w75LV2mK7zU9yZFu/NAdRT9C6AAth
bB8hoOZRcK34L/+C3hrdcTLzUn6VakZDspZX5+vod8sWxl5mHoQIEIL4lQ3mLGNC
GCCORzwQ0VL6W9UlcYsQqcx7VAoSI3X0q1YDSHl0iZt9KZbQEoWSgFkPkX/shz15
DbrIr6VSdh4KvHcsAwzLfFt8XiY7zhJ29V8yWVyblThl1E8G/f7dja8t3qx9phQ7
dDZqhWDHRcF+6PrkOIhNkHhWFswXrAVHbarwTOzXCT6yi53v1l3Sl6EgJKz+lo+S
J+mK93CFJeB27tDGXhCVTo8OY824NiMiQSyu8kG4JzEtmcl+HTES/3E7c8z+P8V/
NwCurayGFIITlhR2XI26UKRFpa5Z/Oz5QY7EnMjBk9l/kb4T15bYTlJI02RIAe2G
Si/+/zqJtwYOuQ4CG57FRfH7T4m6HPXKT0Pcpd/mqgUc/DOErAO/SeXwkVLStHJX
2vgUib0vJPNLz7GnuiA0lsV9X2G08G2evG7pZSE1an8lRO2bn2l6JpMOXofImazB
4UKvBrAmES7Snna1/lX2sXp8GAKDXTAttlstSPPvQVE3H5yQoU+sdMhrjPDUdUJ+
FrbfXeRbJV3a9wKsFFIjMAMOXgcqsT3lerfAkCxkdL1wyxW/h5IALsNk+xeKV0T9
PSKWmuITxbYOycFlQ3Ep87Ce34Bt7SNuDDGYvQ7Lzl9bzWsq4qSzoFjdir8o50vK
jfU0xGpNGBHsxXTNtH70hUhuZak/IL12Z9EyYjs1g56i3xbcTjFjfeYH2EkjAFLo
qp0LewA0TSPAKX/EBAgiWkMo3iXdbWHqMsijzDypV3g47zSh70/EjkMJASFvodBY
2AoTNV7xdDS+qvn4JMagTbZaboQAUW8ieDtfSDrRZOhnJIe1gYEOw6CTg2cdj500
O7/TlpOyQzAPdNRROE21smFh+EmXXzJD5iDwV2649JxAhJN1vMU0ffWUJnsCg97s
+eyzUw7U5kL1l8OEdMugfCFhXzVdSSyAUESG+EqfCxSjKzEnd2k9UvPVqbI1qBQs
jBRmYkMZEDS0ALEwrsgMNewEoqbmPnR04LogM9PkdkOOKVhHMj8E8Rp24m5TT7mR
UA8QoyG83mijRpKMbDAIn8z4UlApPMpoBY9iQu4s9h0pWMsIG9FGBlmAJJmP8uKl
3MfOwSyHp+mUA2XZ2lY/g6LPJ4Jf/g0itoaxIDVA48hW3R/YIat4U6ECaoQ+zPBQ
uW6OBZhBIqTz5eh+6GKxrDmv+ojLqdNrW9Qf3KDer4rGfuyaBBm5gY57xG5eSYcR
IBAQWvR/CNJ71w8ZOPFuiaHSSe1lDEk3F68Mvn8D2QjRlnFoQzIpBevIAehIlA44
lW/G7zdqXRLRJP2JK2eu7XObJZVYa+HE5IKkZXQOtMH8ge8Xyu368NQTYm2BxCRw
/y4uf7e3pW8/fIT0TSyDp+CA+m9OaXgneWC95CX9DXCEfW2RE6VvBXdqKg7CyCAe
C3IC9LfzxKi39mpIl1y8Yg2pZLcA34jdq74Vi/MHFl85HIwJidxbtGalc6neZSWN
eH6vHC4ztlCDjbk1XBAn4aDAJJeV8R3lD1/NGCOYSDvzvLZK9+Wwep8ucHrySu9t
/gd3/FI/C83x5P9yz0IVsq5eiuNrOlDcWxQE0+HhaKLckz7aiXZs7dRlD8jOlTnk
8NEne21IDCn2/oUhFhjWQaHykzD4lv6olBx2AOm15pxCxA8zDQ1Ezg3tKFYaQX9l
UPQzPrNvUPmXljCuyX+zO6RIB0V1g4jo1ESISNWgcAM45MO5wCFqCkR3E8enfg6i
sCdFXc20UeQHaxKVJ9teE/Vwu+utYmKO166h6sDGrlpKDtW3IJM4vEFmYz7g23gw
w+990C1BdjQEvjCPms4pzP0ooekrHY2UgsEE9Lxvg9ai7PrXy47ZienVoTZIllAA
DP72wY/mNs+EzT5YxQWFao+WvC1kaXHniPaSHjcZgbl7kqW+eaKa2C4lLbRZfgkp
LBQNxxmN3YR2BVmgDLhziPr4IVnG6ojSLWfGoij7rfjfW5wEB/y+tE0YCwnFn+7V
Bp9Ypan2+hVyI+VXqAM1Wy1SCuE68d2hX8QFQ0VVFTHt5PkjqJFSZsmhC/aZzkur
HeZHfxrh6OoV8xrtTvlHk25HHygyyQ4b7H6JbnI4nyyrUyjNU0fFQBshqvGQSanL
45c5R07IMuj7gQFRqOZYr2KljIFpTGXb+MDVD65ak2phqX45rkGh3dEWbhgIfkD0
ZyBQ1mKgIsserpaP1PaogbxOeqaJaZK5zg2Hx7wQKHEyuE84AHjVPJSGquKoyz9Q
VytuObB2aJJmtDCXFU7CSVAvPsMHQdpgw8/q9r5qeDzTMP8wyBvtoh/xgl75yJ1M
dbL+oy8y/NzDHqGqg0FMWxastyrKbfcN6cqdZzGWtGv2pwD0jYPTZstoMs09yity
B6b7+2XAfphTqYXBILiUQ2PsHSCJBy57o7xgstKDol4SPZuKUSdbENw+oOoPYy7O
opn6cCLgTmQKFyUzWifzvEYky3xqvqQnCbSaZRkfC3lNziP/C1quZoFh6HozyEfU
8POT6Ew5eF2wBGtV2ujAIuhAJ6rmpcMgRX0iNt5k2a8X9HHcFPVzzwWU0ePLgBah
Cgnj48UFf1c4+LrkqRXR3/1tugt7evD86zib+XEeEi0/kFR13h17M4ln64CIyHGJ
A0Tr8ifCQkzwpau/mddSvgb7e886HB0/P6OgO0lzNHVmsFgFu4iA2IRtw4r+EHZ7
FRUX4PWBy1Hu6wCr+rkJDH8Q7YYUD4/ESdvxy6Z+KT0BQn3FpBU/xbWFVjqRuZrA
Wmb3zOQMWZM0eXRyQnBfULAUzYnZ6ChylOOTwWdDesaO0ZcYH7kuuYfZu3lx6zQ8
QD+uZgjCrZLHuWXYks2iE1NXAbna++KXZwHCPgOYat1CO3b0/j/lkto130vz2TEC
b6mxl3cdD1FePeaRMH17UY36gcD79TgKNxDMZHcARV62xXPqGiRKL2X62mj7hTUg
xuLO6iBqav+tmhPg0jCIUrUiWkr12k1xzsIq2aR9wFmws7ApjW7aieXtUtolcPTv
LBQKoZ7dyjm1QJ4joyCN2M7w1mKoXHOYtPUvKRIn01i7oagiKjsB/r6MBJ6twyD2
8eE9I0L5P9I/NhOUlbJSyWHUmSoRFwFyy8/klrG4ch714B1g7blMpFnsGJZWEHhs
7ly6bgvGRxDYJu8GPNlYTMGO7yAjAGkGh8ReOVfiUC5IzYxYmTXT4s6vB0yGMSM7
XtfRmDD0LeteQeaDKFUEmnJeONz/SFzsJsT4mNOnd5TVhDNXRtKiENJSYHrgXat3
uS/qDoNYqtF62qyrOxeylxLs5WNS9mplSsbuAjClWSVYGqQGG1510RnCxXY7hctO
hBdWuVaOsOzqvKA79qD9izMAw3YfeEDsch3jtzcZG/HRHLUsUvhnvuJS104WAxDB
4RnBQh0br80wbH26cfboFGf7vco1hE81kuu/BjeYL0DtgkYt4KyXvz5v8uCJGapX
bkAAhwZitsEE2OTHmVhNKhkVrH23UAtUUY012wXnfbq7DcLJZYUn7KpFHJ/FcnOm
7S1Yy6okqrLZK0i0h2Yo031DRc4swOtJ/ZhamoNOH+d1nGKB4dsQSzY0ltFAUf/J
xIjZvkUjCoZAEEkEJzoEf7ygH+HEToxdIsF8tdN8qTKSmnayIE7gbjMk9Urnxqqf
UviciwfmwcLEYqrr3fjjsr/G2etSH0m2EsCcSVfp+g2cwUPuz4QnLOfQIrPJIXJS
lfUhW52LdzKYaCkeBvZOdpoge8hYZ09l3/0h37kG4gwaQ1FwkpHPFHxY6b7uuRRn
iAOHkE9VPI6K15cR53Mzll1moSsb3itMsiw3SMV3FZNGj8sld4xstabfqlnUNLx3
qnPAK94A7mqbAUkcmpnbbWR7Efby8mPhHFYA2ChpkT+fLgMEFw8n2vpXbvLBJFlA
txraJtvjmouXhJCatMinUUFRb5YQfzg1Wzqyo7mGEOQ5Y7SoDgSHroVq2Cco0hYA
wD/39HvBCdS2ruNACZ8gfOU8JXPhE5YsBJo2HfoMLbcRYndtPeD34s5TRyFRz005
Q74hZspdt6uj4dyUuAHaYoA0JEXj9Ex+dVQstv3rMzffF4XiJpxuRJUNSG/H9K5U
dbxj3jR0rrW1eiLQAXj30SJYpYmLXAkjd12G/R82Hv33+Lh2qkiCYiZFaPMTJsRH
sdMV+UyOxMapJsMLNv9jZwV335ZIqpLZTJbP7KFFqBmRTZfaZVTmV5B+tmfWfdY0
ShDvaQtGPlPkPM/HBenxL0ypa2pPhYw8A3A/7+TZxe/ANq0XntCcHeNMn7oQf0hS
q3V89uVBVl+R4sqrUeTXCVlF4HCWdJ3HE3h9qx41kFHzlP3Jzz4PR3pcUt1eEA8+
mqyABv1pfihMl0t8T+caCq8Bnr1MWLQ/2uF4qHXEnUbvyRuqyipDvxCbc1ExSnB9
6P7HJmrs8qBxX4FkQR75oosGyXRpL/ahXeR59zQirF/GDubO7UyR3RVUo3ulYlZ9
ajthfg+v+nP++VZD1xlb0qKhKbvNaNwruWsrc4OvEDXFyFspJy58u40elsZYLhgJ
cTNFyI7GBSA2OZ/VdKvJNGKiypjBOWMmZOORe4J8d8TjmqwC8SkgQ3G3adLaMZFK
aFya8XSDriXgzwcHg8qtDLFMGS3nx54N8PZJbROVOjmT/ZuAA15CPjbeT49Qhv/O
ob94zQqF+/0NFu6avC6cez87BB9V8pYOZ31nkorrPH4o7dvIW0819tQ0kB2eYCYd
qy7Nnw1UF3yfeE5geFLoiyVL6iq3OfW2gF4FzFhgfZRfvZqeGePRonkXNJuX9qKS
j0JhsOpbpqp/wmTbatuQ/rgAfS8sTJ0DtokQiE+uUApule6X5zRtqCIjCku0/0r7
Rotdgz+mkeVmsehZqk4S0F4dvlihp9sCinfFrNGkrx3/rqahsGZW/m5Qn8FClnih
wqV6F8DPf/NjYNnzQLd8xvcwnqtvSVpgsBDgY7fnaoeZ3AWbgQKgbZ2Ir/EG+B7T
IiiSrWXb6nMMh80yhwKYynZT6oTNjKwfyrqT37jWoM7q8M3xVPkKaMKV4AwOGKTJ
AXUfQ8Zh2Q0lw7euIxIMkUH1NbboKokExUfJ3BdaDb8EbAhyCuf1py0aV3bGOB6E
qn02NEa8YvQq/dtRMzh7Oo/k6ZQFW0q1BgRlIxm9HJ0EVfY23eK+sGUdS6IvnJil
ElphukgN2cLD9bR0DI2aQ5I91P0RTNg5kH0b6cedXq740CCMhj/r/ixgHZ2qxzYK
NID7p5PUp+Ovx3rGx+CLzqPrcD9x6OGmZB8KoWdzRdYKQYC8h5UExw6jOVukQnVI
2kUBHyqZA2Ye660V5WhjzQx4DGAwFEN3vqgr525W63fXdjZQGAbEcuRIXwgo/Bnc
AFKccrk7/qj8TdsrYbZIct/r6vCJILIgcyyV+1cqsjh1vQQngx2rWe010aAP/5sd
pizcq0Q8p+1jSYI7XARo5lpJ06m/XgzLbZyXkQlphBMXXASJ7W4Np4EZ/eyfTb5I
oBtGSkNQGCMA5OAtIUUMH3G/FiLL3SY6J7a2ty+Jh1cNNssm5XmrgT0c36R3NPlN
is1JE/CvdKhqDJeXhKVWnkWKVzq8tGSIdTayaJz2KgToA+hfhVJt+K1pSHKenV91
K3EcYUBAY0DeeObYrvM2uxwAHe32KpvJkT6ARWwF56arREwNYfKyA4bSzlZUeuyC
9YEyFoXtfH/FrWQujnb7MJcfRCAgDiIHCK43Nh+XRWrzjiOsiR29+2m7ntQ0+hic
IdvHiM3BFU9/2fooZx+g2hJqPp+7OZHA1iGIRb+RMgd41Lb17WP003yaP1HNpW78
wVwYiOVTGVQpum1Qt04BHojZt3atn+PzqBl4ZrmcR4ERQy22Gg+6aJJPsILP5Ee1
Uts00jn1W6n3ff7XWmOvrVoXZWj9z2Qnbx0MfyH8lv8y1SsZMBzRmiXFJuSHni4+
ORKfjC5/Y46eT8tPZZ7Ra9FTXyla/zPFQ0Y/jzR6plC16AJZnucRX7wTH7DTd3bf
pZwpxCUzHdlF71M2f8NnjHp7C6q/JtTpF5ANx5TdbrGwfGfJqQ/KsyXeNEebJ9g4
ATnasa5o/2SpQWTKMfztqgpxRS2UPdpC+NmzyQyPBGXOkIdmtm6P0LW3FNqzc2Ym
Rwbjgr9ATRMZJe5K1nZi2jl2Ob07UX7PY8wVjeNPYEECuv6rtMZ7ZS/GTpkEfH1Z
PCrCl+mgnyPxQu4M2ADeFx0NYcaUSerBVB2/wgUABHFWYsX8JdO7UqEzUwL4AT7Q
G2k7U53753MtaT7WVDMm/tbGLcgkDB4LetF0gODdM0Nq8VrUISCTSPOu70Q/2DYG
qgtvI7fxLBjk9ZQ5Fk+KkY11SZRDl6Vx/mvP82nE2cMTbVRbp7cIf3KpKfnnM+TM
WeMdEhOY2ZF9qxPYgcCxEE7jLg4Q1AqBwaL6hJadGx9kSgXtVymO7Khb8fYirvTD
rUg1zbOcY/GEzJ/vgDAb38N7kuAXu7WmA8Z7tGT07UFbisEDNsC/XIpeXRGFXX/o
4NFrr/XCDK38+NdKMFnCbWEMfb8hpafO9DqZjd3P/8IxpjJFh/9nW69FZLKeSd7H
lhd10SXMXYnP0MQy0QvNYr9YXESZjCnNlHwvpHdjbmt6ayb8PG//kpf8MRy4edzX
RS18ZXoe3Xgyfpa7iSPmp+Cm8M+K6zCK6C16ysZfq7+Fw9lgpljHpXsWjBSnnGrf
jxmuMmUUHIT56i0m9TgLlvAUchN0U++SXKe1iVJxJmor3kMzcp3s3RpiD9yYcmYn
Iy9m/XXVHU2YyaDmeQhWNMcLt6M3Y3cRj/3DuFjHoQzMT8jsA5tmi7G9tGuJ00OS
q9W+Ul5Bsi02CRj0FCQW1cKTE398iyDt54uK0/kKBUJo6UhnkKWlsDe2TEIjrn76
aW7hOEZW/z6xfcMeLsoZuOBJVUcADzO9elazm7MR6P3Wgk8anZoaO1jmDJK/m9o9
HmeRzurhWiiOeDOC+o43orUQLr2mV2Ijq3qiwMvOMH8xtPkiRWCXVl0Xgwg+GNHX
ZRvip2lmid03bmr/KnY5FMTpM5ETKfiqXOXvgIANLjKgrfrNlQRE6a9W+ZEqMjGE
Yasuq/C6DK7LCJnyCMNj79le/QNqB6cembSMAQMfwb7FRP8hjsE102OR5XRBIEbY
C1ywLQDZPBiu/WzUpo6QDntITTiOsq/MwKruFKuIb7vq+90CvCoNZe22EI2YhVo8
lOaUjmfHc67hDiXWzOJe2qf9iqsVfOi4oqvmjy6L882eL0NuMy1uctW8Az4Pq/+K
iFZBaBXoicAsc7N1TjtKhY9LYbS5SmG6kSLpb7vgdh+wA2KgI02ANbnbV/Bcmuuw
LJoEHg6MoIUVLXVJuDzwYqvt61ijgXkSb7mdLNEYq67Mu4UF5njosUsnmpvlrvL8
IdJizo9VnPOh6TqWx6B0P3yIITQ+Im4PLWYLMR/vr0kAfgGy7Ud9XN3Qmdfyeo/j
LEnhtrLKGXMQ2bn0zI1AbkIeE0h8310ISUlMfHSVwWFlO4tdyDQqCtzR8/x+6FuJ
WlxdzEAdTiFzwUjCdgtYQuw20hS+8oljuTsajdBzOx5EORXt4ATb8M8RJ0bE5S7U
5yfQojslP2cyV4NMFm01bi7U7CeLM4WFy4mTx6ov+Tf2X/wzcOm0Z+NKjRZHVzEz
mz1/JD+hbE8BI9fKIs0ZIP8unHYbNZ4LvIt0V72YYWyohHg4sba1RZ7dziM/uqy0
gQOeLgyMlUKJkg13g4G6vXQO5Z0NACNLMTXIv4/kpZMCP3F+ghnZ4M9ojDDTgXTs
atyMSswrw/2Mtu1HEzYB/UkHKa23ceMPxojswmMxTYEMsopr4BCxu9b6R0Lluph0
LOjF96sALIcWtZ/k+w8kl+GMd24XbZuY7sm4cO0PrjWmAuG1S3Ejtypr95emM/VQ
SFNy78u8pzi/f32uwM0zeXjlzPSBFPYTroklZcTZiX9xDZA+/n7pwP1tp2zA0fYG
zwqGDS1eR3EVfz4GeMj2JkUU17E5N8akBW7k4ytKjUhcNRhkFQeybG5FrU+wKXvO
5bczMb6VF3FqhrYGnCf/Kz+ARfiCqpVm2FPD1NT10ay0/IHqJKg08sAg3ETxihNj
ynakQB5l/AzorarCpf23YdQV5Y7Y/uP+kKEBOLYsSHvNWB51Hm0QkzvMO5AiJH8n
qj0BCN5f8P8rr3Op4x1hKC98q9377kM8YAkSiwV6r83mX4ygJtnzPImVE62gC6a7
65E9OBGIUiDc4AhwM28uxtGRUkjUQa6myg3MGgf29OJKAu2kg/i0HJQsNVCc69uJ
0splpk+hJxAnZTemE6mxXU9C8/tZtk2xo1d3r2d7qWbbi/7/N2bH78t/AhJCceZ5
BghdxsCoUmf67Bwc8QzOH/+AtUIIojkD5poEpfm0eDFeFOocp5YGnBYPym4IZZ2s
ggP8b/YcVjKtmA/4RlN2AGwU4A8e4wogJyzyjmY7zVO6jW9+EmWIaQNbLz42ltqf
WwcHo8iIbFFJNRiy27eUmk2ziNLkvwiyX4DSlK9uT3ZryK0CAdQvsvnlLYusviGy
YHNhDEZjLN9zTY16JL0UdMP/SGK8k0dhB0ELT+ZVF2pxIKy0RcOy9agJbAO/OulA
AGD8M1J68PA4D7lTambZx9gv2ZleWS76Jy560OPQselosO95rziVXJ+Xc20ugdqw
RoggD1f7P/TzUjxlhBGSxtgbrLhYXzdOm52l+qP682EnkkO30fKL9qlctI1iRn84
WMsfuB9f67tB5o/H2yex/iisQCvN5wKHDa4Q+Er+6mbk+ozxcXzDyaFX8c1JPEAS
2UJ0lhAQd9CX9bXJnv2DbRI0c5kgFSr9MzQlaQTzePRuuevV2iWk3bvmv//E6uLl
tBl7LRIe5r8uydtnJGJm2hSOQeWBo61lhx3fXJYxDI0Nal33Qi9FG040dNvMyCv8
k6sxqRmzVXUr8ja6Qli8d7lpgO6gRQ+UERHb25ePFs4IBoebP1EnK9PGKcomA8KZ
LRQwPp54riWh9xOIH0srXPzOGzMV7lQ2SdVXcd7wobHLEMDelhuXKjfwMn5CIdML
2t1lSf1BXTaBTIn7XeslxcQvoyVdsCO5jQRg9rC+CMzRXVHzuIOYDKxJAOdvvBcj
iIsU8p+DoOojg9+IH+K7Cw2aha3+gQJDPtAwDL2mQQ97R+JUCJCc1ifDBD0BPsSz
ZaiZOGBc1Mxh/JH9z9NrC9Q8d7HCbZW2f2hiQqcDHVmrpO5mUw22xOFevCU1kJIS
9ZPxTFaX+dlXyBlzxbBuz/U1bQZuoxFM5XhSAF9AYb0ZOOmUfEteRQ2M5zKzWv7T
VoEZmB2Fi81THCOwlIgf52JpevPcTwXtNu/3psT2G3wk9nHhIK1Zj3jWiKf9N1Fd
JdF1dzfy57UdHeNQK6TCegRzulWxax8eitbX+3+IcWnDQedXj0Eg3eLAuFa8rop4
kA0Y4yDCnQA1VfgHB3iPrUAlJXW8sTUmH4Nz/tQuBh4iRQURDnfhjiiBjrCO0OS6
PmW3AK8+zJDgusZrasSMtHj/lyyxkv5narWaNL+RZunxxDg1KRiMJ9+3BVnsJBKH
3ThxqcPE7qhhSJRRDBkk0ixCzz0bb6ZSnj55YIx9mH0zFdGK+6tFxgp6hjZ6Yc9U
mZu4Ep8J9JVKkXJSgo7Bxf1cR0CED2ZVmp1NuNK+e/Riw61o6Uk2gcPrl4hoEMJX
W2a08cOePFPDdDXk4rlPI01yX2rW23Xnbe965yuCGdEbX97BIluCdb4c0qX+Y4M/
HfN4qcEcXvfFWGQ1Fsvbj5mMHMyXTLtfIBEFD3Dstxko8WE0kI4RpynH/YUAbcW9
N0oWNUs+UXv7i7gjoIUyVS9p4rGITXoEjm2INeMD0rzce2mC2O2e12E4n5LdVtOX
bFZk+JbGm2QqBBAdM7+dWGWT+SNaLUiLPAUbeDzRT2V2aKQl6tSI1QX6qiB5wi1E
FqK92Bu32OZlpT7BKj9Lm9uPsrEF7b63zeTtSke136+n9G01bB9gJcLS/ZkXuCvh
3cPlW7/JdKTDJUpdA1akcRzOXZS3FvPcfqLE0x89KuhLN3KEc5qKf94wMWKmC+PW
17OgPHfQi5gxJx8brhLPhMF36NZwn9ypn5AWj1BxMI/giZqUJEWV8834KN9vVJ+D
vK9lNHzElxubsAToGWAbiJ8oxEyqgMkWjmBzpDxNVQdhlgBtT8hEAUD+hH3b3IS2
N9TeQJsMX6DNqdv5O+E/VNrLlRE3J2XPrQbUD7+AQBxsR7jacNBceRs6BidGfknS
44VRREirBRtNqCgPQTTHFzC6oBdWGt1QuEUA+7aqrrhB+CI5PIKd0yKnsHZwKSuB
V/+CiyMv3aTmCoWRjOCBjO3yAz2Ig4P8shZTHuGjb5bqMfNanXbdhSi5LNbvdTTU
nD0BnR8I2Re1gMkizynBW/7ndNyCI6bmCwOvnD9taygAtnZPlnOi3fkc3iYr4wZo
UxRLSA3yx2gyMPZsvGXT6Vs7BFJZHwLtWPZMkCa/uyOKn+vbR+4Xl+7OMrc1Abwd
AupXeteZpMG/fRFdCZ3hFh8K2lgJ/QOfbF7DOxQE8LQd1yzTUyBw5cJj6nendAXU
gqgVdcDAa0cmFDw2si5GRsw4jFycmj8ipq/Bls9M6q8lH32PJnAZz7p46kNMJDmu
jfzwRbk0XR3boU6bGOAleq+ZyfkJwuGL4Xr4M9VgY5lBaNFO/Mi/tTe0KCN7Zj2k
MudKfM1sx7tLA2INBhWLPkgnyZylLHXwWSmzqeYAkZkVNioGyWJKKRGPUPdW44dR
wUokV1/dbbJRMTouyp4mgeDiPRiNk/VuRzC26z1VZJJupN3yeYqrUBR1EPWckNU4
iRVHjSCATYbt/JZAKEnOtmc4dEYa03yELfEvU6lktJcBzPE9SKfRRMdMVLs4lEvk
UKcVHgNbLSYJPiRhytRJGuygm0uLi0fTsEf0GKBeTW57+uWg8ZKd/fXzRjozYrA4
dH8vsLLToOnE19V14cMHdCaitPTlo6WWb//8Kvni/gSbkLgsivJeFbl98SVngecp
dBhzuJ5s6ZBkPIHBnpm1wc7ztXpn+S6kM/r50XQ68CKCrJ/GGJ3yYr5r0pDKO4o5
gUA8lz2/46Xg1MU6179uhmBM12k7wQ+1TDh+LU2jcFu2wxbe6T+faeXdJsPOqgeY
uBxL9sf9gDuvE0/okOWGHycpQ7Ix5cj/YCNuwm54kqBP7OGv82ZmuzNuu59oQldl
3/WaCBOGvyJcLMUplVVs0vFBmcHFEnKC4t+izYEd1Bf33cuS7CfNs76Dwb+i+w64
7ORoqVhINlNPBfc7vZp3ZgJE+uoTTRg993xRH5bKT4EFk6kox/3Yt4T0GiqXF02I
g0Pppw9xHWyuc2P/fPxZzB19e/dSJPGTEGJtrKDdZo1bYbcxnZBjGDbeqdcOA4tr
6rvecQ+ECMznhklso0TfQroB7vA0gBfeOwo5hoKaO3J5iVFWYNXTkOFqRhwk6bT9
efuMva76v4hhoNEkLXvNBmXjXJQnvVpqs7JFLr2N03AeLnSW9JtOpEJMmc3QIEaR
nx7xXEiWaSlB5+T85PWA8y+WnTNGJw5rf6wpTkpQgrazxnrjLRxP6kBVcUU1ef4Y
bMLtYa/w5t6KVlcAqTsGdx3brE4u99S473jfOwrIUvkRHPRoMCOsWpc2fWiw4y33
MQ0XTkqpQ6Pcvo0AJifi6VWDK2leejUpwwutgLgwAVfGQb5r05tc/xt9jkIpH02g
FU9/phPUqB/VhY/QjdMesmqOq59opP0c22fPkjvMKjxFmdXQqfRKTrKxtD8KyOQF
9NPihdlj/CP7A3Yqi9iJjAcpMfLXusNQze2VAIkfkqlsogTFrTjjPN5POa2s5F0Q
KdO2e84K84XcqK/o6hSNWFhkmXCovvN7LBigq5YpRiXQxXF7Zptbk29w2O+TWRFD
Gu3vwp5WqZzFJJsY0eh0dFP2v9YVv3hchIBVOOnsQlIUBKhEj+OBKZ79sp/md4kr
vi2V6me9dAb6F/Q0qE/a0hxV1CvtXQjNh/3k4pjYmlDHio72G9kLWEwtr62kuPyJ
8aXCRrD0pf3FMqlIpT4xgo5MoR5Rmtr+mugThCLbKBiSzvWjM74au4E3JU52Q2gr
bzmIucPuENopdZgxfSVkd88QTzn7jdK0RYTENs9JSxlLcbfr28gedkeTOtLh4RRL
zj8QAEAeDc30Mg36C3j1fLJPe0oa53MvVCkzGW/GyfFOSDqdQPqWlik3DdoW+wv5
T5xAlqe2tawRfbwYYH1Lv+lkWApVQCr+9bk+9Dcq9h4FonhKACrwVhEV9nIMhIeS
HZJSTf/06Ead0gXuslVXHlrJwKXCapE3aA8jufy0kHVFnbR95vQHPPTqIhksl2R0
aQPSkq0MkK8r7aWJAm+IgMqRcZHYIpthuxeuANL62XIiOFxTurkmMxvtn8KhYSVu
Z1Ls7JVxQWmntmOJea5SA34+hz7JpXZM2XanAsIUbOxr05hU00pAocSgj777vmK5
uy3ucmwPIUFTn8ewY/C05/5bebsqGA76MCGLwHmHy3Hy4zhWb9P/YhD8umuuniQj
jIDNnQQCZcOAJmblN3A+RlxmTp49eVteuPyuSOoL08xNlYX5TgymHGETVZCEQOyt
1926R+//YMmorH4Igz2JOYntOjUvTx1R8Ey2yxl6SmfblwydkEcfFsa7VsjJRu6/
H1ETsAzKHfWL/8IJwZaumZGT4aPbBo9i0Z05zCPhz5vOHRVP0IUK2jXZf+UBQ5vt
lCISq5H7EFL1Po73Gcudokq34ZfkHQydK6engBZtTtpeGn4LoKHgJtM80sIkNP4q
Tr/LkbYux4PEGN818gV2j6zrWCruFdPa5Rt5siD6/ODrAHR8SFxzq08rCW7PyRks
SvQtOxSumr7YowsSw2ZeMZWGFTLCSAg9RK8d6Plp15QWK0nt8wPEG6AYHSkwvahx
eq+PqoDlsUhLixXhicd8ijVAVG9T4H3ciEw5CQbAibxuGrp5H7ZGZBU6uvTl/aXF
/lIjvjNlsZgLgnv2tnCdRS73sSV2RCVfBUF0eb6pTNqq2dyu+QKxDgKDQg/y5uj0
gtL4bjSTFSnCYVW5bdYkWvu2oV2qZ4xFXUmltlI14+dwwtjPKEZKEPUvF9OyE0Sv
PvksHKffvy2B0kJqEmfYKwu8DKjT0kcW9wcpX8jou5hbtg5auJ/6veRdr0S5lF5h
watEVVr06NL8XcjPh+pa2L4/1gFYFvJBRBgZ3IAhtAQpmLGVGp0KEep3Qlf0Xod3
aW0zUUOAfFtX2ITX+kSYkCUvPSkhhVjTXfF/SdNYpac+Oyj7x0qKyU7PLiSdGwlg
5djfNef/KN7xi0y4j0N7fen0F4UGQqv9KC+3vZ6vYN/4UO2iHn1nf9DOtlj12SQf
Nt5zG2onqXm9yaXTEAFNZkuJ7O4MVDsgS4SHKCxU5c1lYs6K03I7A1lGz2W4jAfa
K9iA5CYugNbTgqMJB/4PoVvMKCx/S4mKMt9BpafUPmLBpk08rYZSJDwAECe1xthT
0xgPcEFb8ZN64w2O7JtxYWOUIXvtjIJkqYPkzcJZiTcqp+JAl67VCWmpeTwZX4L6
J9UFklbyDx1q3RljIp6bZod9bRgbVJGJm2ybUi/nvZgUc3RgK6VRcBUCBGLu2Gea
wddNar47cOFzy+I78iY86d1YRXNV9nJD97omCxCtt30cuOGV/36Qgqty1LgF5Ns/
UxTxVltJqQ4OCp7l1hV6JBQW3DK1SePuIOwF7DVF61S2qiGWZTvfieZh0Sb1Hu2Y
leQhDRGzpi++ZyEZTYJNwiREbrV0yI20+fi2n/0NYRdc13gWGhzEP0uTtbNCYLYs
9qM2BAPNpwXDmpCZRI/xefPJw0kbycwOCQGNi+5ZlgtaqeIMMCrfcYOmymzfaNZs
Y+zIr7Xe9UMDF+ia1hOWz+2qriSsyglib9fCI7avrgQIf1vrCcylPHKb2kJ5/vA3
Vm04WRdMToC8fcyr85hSHf7xWhlBS3R7Wxgo2gEQJDaZfQe2ShLuy1Ti5i/jyYhL
4j46+8wF7csiwv1ntouefWUs73N83dindLMoWoHZAjIkHVClyw6+zfnxmVybYol4
+2JAKLXLwQErjaqU182kU9zAtOp+N8QaXQ9HFStmVEqVKzMmjXKeEHSC9KMBkWwd
dUllb0DbW4M6O1ZIjBKkom/G3S0wTq6S7W1hdGfxffl/UMHvF1rSaoK67Icm4Oqc
F1FkCLnvysNkxB6zFudso+U+Kf+Buai/oCGanhDDD4P/WWeF8cG7g7CsgsZ1NxVC
lsiE3IvuLZck/Zy3uvuJSs3Rgr3FWSiPgrPb/Tr1zvL/wJ2PH449DnZx63r8K6yH
UatniF+kTzQye9Brvn7R2CYEWEsYROn7OSRDvy8oaAXC+0xXs8h+sgfIGs5ClTH6
s5hBcmoK+nfr/tUQqa6uaoYeamXDuEMgBd4e1XYJFff2k/SVxP+UAAhCyu6+KS1Y
zNlSizaFQSIZoSihz4AXslhZDSxy5tkRyhWlabKnyRTB1S/GhKRlAdBt8ykiTew5
+LGY3tRxt+XSxdImlX5L7gJK2lPi4pR4ExftOUyqQeSk1f7FzX1aH8AMRstsx7Kb
Rdpjtx+PJOdgLvB3yYsUL0thYTahlHG6cavOHk62S0eh9mPvxmCTox0IQ2cS8Pci
eGG6+fhyB3dnRacnO6Ld93TLL379kcitSfUkusKTDLNnqBAFBL6pipeiPjni1Bzx
lPLZauILcxXg/8eBJ9UmAphHWC1MzhKR3TELONS5sP+R0CK9EshOgaZPSk1tIvX/
pk6sptRXfVNBM5Tk4/aJFs7cP1NoPLYiHUhgMbE3RO/xpsIx8HvKudrUTs/t8egx
4Zszvn5SOAlG2Kq5mczwX8cyxjIWCwcjP7xq51/Egfxjzi1wmqCVBRAntPof0LXU
5t8CuheOSX0ZRag0rGgvomkGHsDYW+/iEATHMBVBzwufAZXUbYs+utnWSJPqESX9
suaB5VkHozj/DvWda/nZUXG/2NBvvGIQulskmApM+9E07sKzXxVpzqaNgL5VRyOk
mutn34m8lEB1NJJiD03EYAQnEdabQkj4lPCoa86XN/iSq3iV/1ACR/CnXZK7qHMb
LmZIp6xxZay9ruH922a3QQQMwvXtoXVO9n3irFPmrAxoZQedph8FeLborFC7qewl
EBgzImTTr+WwJBecWy3Mlu96d+RhkT6Q9NclP0Nn4OKZfM6Plpitj+h6ATfdzs8p
Gr6ISm3Qk1GMU9yvvduybCVxWVBGhT0qqGdXkuG0uQxR8h5AzYyYLVHunb4GVjAj
MRi+Imckf3vE83DTffZ86J5cR//R9Fqc21hSTzcaVsoEODeE/S53jrHdaPQYWVY2
wT+TGFBFie6s8KF1XhDyu5g/DnI9nd4oxLobEceHOLK3P6iP7FVGD/c0MZyZnxxU
b92Ox7VCe0fcLgoQNMPS8AG4usYZ9crSY0XAU+7tVAlfwdiBtcc2KZHRY5SG997Y
y4pjohL650oLtQpPkxvYrZFJoLpQT7jO4l4VvFPZEJRCMB5RZKqASI71w5iTLp+1
ZC/OvnLW+9WLaEy/1WoIqw2RUmPTikQs1pDm+sJgV+GnSpD7d1LdGfADT4wnWxQ5
NX0nL2BUOo+KREUEcuephiyGvZLGZhZerrDzInkwIy3qOpq15migZErLwK9TnzRu
fds86EUVhyRLR/GnBe8eIgT2UE2HhRPzTjR7R64lgOdrt2KVpO3tRy5EYC8VG/Kr
jkr+Wlv1PdORC/R79zFDbbw3gcTC2T2TXD8o9vaxXJcSzrgLit0VOTZc/8osXI6A
rRzNzQ98S1E3WfU6TI/jU2dXy9AZERt2RC4O9k3M/XghCLmIesnL+f38f8mc4MHi
bvt+V8JPHndYKBEYgagfQHHXZLgPt6sav2/Z76/4tUQmkLlW9nJMGNkxWonaE1z7
koD7PvkwiMBbJpmFbLR1qsioPUaIFgtMuFgKw0O/NbZoHmLbex8im7N8whkbcBeB
JohTlC3VvfBu/bAkhbTVRH8V27m4rvU176mGD2uZVg9cP+XOomApkKENmHotiFFn
m5euMbnyTouuL9kRX/tnWAskuRBarE9mkVes5YXdwLcBjpKZJni5TgRMOKclyz4i
/mL/H9Un795+yd1Sx61Do9UPLanKoE4mU+dn1AV1feY0AIBocxtgzQ6OjOZxh5t8
1GZAC6osfgCI7JsV4YNXcOVoKDCqlFw5n3HebnLgahhFIL2K58ZOHXD9XvTPRwHo
0AL6hLIPYOr/cOjyEnWAGc/FH7ZmLU1ggXzZ/BTUJ+xrx/nbB44QtwgOFegSwMCG
BxegRppKDJznghOLIhned7/0/n3/g5ksaTMy0GTuHe1PDVdiutvictuswPMC6Whr
1lEUnYePuvS6Z5dXga8XscY9mkkWJy1Z9EzZA5iBFTnaJ7HgtTdVoZtvVT5w51tO
RkEB6extPS6yS4r8AXabvrl70OGLpK5vDvDqinAW662xY4T/9/ouRFppQCHnCByd
r6FN9F+6g5N8S9B+9W1jvd6UZxUJ5fafwARrlqCkU54EUBJXcQ3wBFbA2G/wKNj/
mqcwJ5DwBxyVb08qEQqso5seAz+mcfbn5rKt+3XULlGFjh39Y29wG7zuekI5knNQ
FJe7gjQ+s7gBEppRIytcEbhSAPII5IljV/7ah7V7UlkPGuXZpuLVVndTsNBG4Ugz
s58xpgJeKfb7sv4tfxNAaZWuVf5kEoKGtjECOj4HdDp0Abe9d9nl53BZwDkcOYXw
iTZCTgny8VGryj9jguNjWqLTxG39HZk4OyWaWoP8+p+C2MSskFqClKiknZd9FJ70
ZFqbIUn8/GZUj7ogGpN3k5YF4hNkqAqEgBo8+EsMvXuSxenyVAVRZ2PYOny6VMtP
wOBiTmTjREN6qC7110+AH/Wj9iKTDry43KnnXqNMdrtjSzng995ZH8ooeNZVtfwd
+6wUfqElR8HzPIpZotLERulXyjKAgJzq0pAip/zo+T+++try7phoKHsce44NGrlE
PaAOEJRxh62o7FemIpViiSKowNv6GvOSRYnNHfCpYgX+JiLo8O72up9LFE/NV7D8
SK0VoaE4c2Yl3alUv4wgtKfmkbsoNOiWbRuaYVRkdSJ0hAGpgWmfRITtqPo16G96
RJ5yOX5FS9yr3vAJ59Re48L+nivAu1We8GZp9JZJkHCWK/s7wfzVB558b1MN2n7s
zNO/mFFrkAlaEKwbO0xcXxfUG5cYVh4A57FjbAnigmD6LLzNXAJq61fZTJbSmMqX
CQ/WEb3HSbrziB6xtS1LJwxvXSzBhZDk3dk75Rgi+DB4SAMr/R/lxQhwqkqvq2hZ
AhdapsnJv+VeRNhcP8OwXdUchUGi2HTxy2moPnpqiXowN6/sq2BVeAcwdaFLJp6Z
ODs/PKQU2IK2JnGhm+2Ss2zsjuILAWVsJr+LZX6EzdboyrEILCRkJ/pll6L12mmL
Lga2Hus1Xd7P2uw8ZLNzUmHA769JNx8LEFmXk9XvBNjxxuMsJzAtI15Kzf0q9uKz
VCYW6SSmUSQHtDQr9HLsHpEDXy4tYDJxJZXH8Tekgt0u2ZoI64n4RuZVI8sAvgna
DF+7ouUtAFfu9/8KrPGg+W1HZiKCTCVvGbHM2aJZfBUG1Ix0+HWHeCWvi2HJsc1X
skNN/87XlrCzg3uIJfd8rl1CGWrfxVKTg1vQXlb4F+91FoUtsllPwuMW5ftRmSaX
cyyJyZGERsWHJQj5FiH9o6ubQh4mvUExPB8XzfvApTHCQDMHRzM/5O7ApccE4Mfu
iPNLXH95EjH0jBmHoz9F7Sc3M2X+z9N8aI8GkXc1nxILk47AiMqm6uOKyMSav1n2
8KqyItk3C/qJiG23gaELyLFfOz7MZBlYG8Sww5lpEwfP2tEKomStmTVjmlwuNnZ3
kPbgK9MDxA52Gr03ejcty+uPXO/LRDaeC9nxMwNU6QmwDSbhqXqOITRC29C+eTbR
TcF6wg4bsPjuIXdYZFuavIvF9Skc9KiqmXjjHkveuizCzX0hmp07MXUJPBszc/34
PadFR9Ob5pzv98kGNxcVR4iDl9ZaBZTMvHolU7Zf1nry3XlaVjvBHLGj1IkrYfv2
UQ7yCAT9LCi3KMnS6EfGNqcp/EdYg/zuw7RmIJur4qzqKVbbUhf9f+d7Nqw135Jb
x34wUVC7Dhw1ATEMmZyi+4QzhMhUS8wGb2mgrwKD2XX9jj8zVHK+IW2iUKZ3NObz
TrN4AY47BpRE2eKafCctkwqKGSWBWEtt3/M7mbNFzy6CTooEwrMeChQDodGIFLe3
2HTZhHvpB7+VaDtWqol0JIobTs078WFC9zDbrgD8cj3OQzUk8oN6nKkhsbzCvKNm
EL8ndE6W3n6k9D3vjlhdpfysK+7Uul5jz+yRNwJyIeZM3eNQhWZuz8WA8qv42HjD
qxDHbkriVUEKQGhJAiwUV8xYdx6Wm2Pwd5LUTLkk8TqLNC6/3Rda4NxLU0IpW90P
MlW/X1LzLTdzleB8+gI4CFuox6qja2Y55CseflDyr0r1F76cO1ouIaXRUjGgrEve
bxygpWGZA4Oy0bjTW1Tj97VIH7Y7UFX0IMwNTMf19lp+rVJJ8fjQ1RzkbfNaNUUA
+YGp1TlrgHJzPBQhzQXSgHh49N6vkkd4h90UT3iFDuS/Lunt7NnAm2vJVCt252ae
4DTOOnwb7yS72K5AFdLuqfSc03o+LBsUCqG9ySqGb9LJ4dtPAB2yAh0/ZcZ780j5
npnv3/hI8PHX3m/ENJ7+DLaE8QzP3VsZw+sd/APc/i0lfQAg+Olq48ztFkTAHMwr
3qswLA72GKmU5Mwu1U4D/PcWfqqiTCEERNMPTNUnHUrJKQfCyS+f+IDJP221HwlL
Oz7dOt1WrqmfoHJylTQZjeqSSmRBonhTJCUig2SNYstPky6yTJVnzaol1yFuvfAL
Y/BWGC9zp5/l4OBKw7ZuYVg51BxxbgZrbZRTj7C9xiuJRLBISqI+mIZ/u6h2CmbF
+lSYEkzlCgn13Tl949HJZoqaccOJ/BqzGCnWD3lI7FQvuBYGADPT1mcg7u/sMm81
Yul57ju0Ltc6kk/Z10AK+Y2L1hW6iSN5VS7xHrpjIzePXapAAJCF2/xhk6E2Ki8u
l/TK4QmES/kt64dDnlhoiR1mud/ZHWqFMyCF48kT51QdJ5SIr3zLDxkkzSGHEgF1
qRgZ63blSN0aAhUoJdpV1fK7xSch+JtV9WjEI1m8TSifqq6RccAfW3Yb8MoPjxSM
r9WsKoDZyaWT33ESKtI99nIS/TUY6w9dyTTNMSkQ3TQBGSlgkehCifxcQ5+va5lC
oSKfAbADh3QQ4+Q8ue96TVNX6Jzv6u/E27nwQLThKOE38GEQh01mCT7mnU6r1Vfl
Il7o59pzudypbbYazo4oKlsHdTmKBvQSP6vPZWri3fVI3TYZRavZr7e4N2lkB80j
/0lWnFuLoRcxZ7cZ/Y+Nbah6WPYmZyJeoSOnEPeds2I96xjX84hdIVTGxb1a+ADB
bLosTWB3YMpnOR84QNz7dwj3xxwlih0O4EfCVLNept0WzFfpkurV4JmCPrX65p06
wEwlQUyisXxGJ6S1I+hmnq4mXeysvBrhN5ReNOY+WqKxfmZEVlg9C7fXDlhnd4wT
Vm9ppc9U7EZcdH174T72ivRvuWhcsId25tX4mS8cbKIlDb9bMCK0LyeHMe11vVin
cT0UC+SJz/pKVYOc/51bWlcmNzXwL+LAdOTCiJdl4hmVoemnr4Kx40MZh9YCM/ni
ghSvIBuqZZ+AHc3Og4TFW2YjH+WFQzMl1mKv8+iavtrEJi5Z0/dnuQy5u4BcKS8p
SPVKGT0oUPZaNj9q0u/EGGkP/PGCA6UDstgdgcQPnFiPBLtpVs7XhQqaqgxY6LAs
gJPC0tsGpYZylBB0DY3+hWneIvAmYHlXGmshgU/XU8oaVCPhSnqmeP/rPrbdeFGz
A91ybuZvrto/9mUGodUdBt5nSNKnvEKn5tfBa3okvrbF6rs0v2qEZx+TVftgGQLx
ePuRkZZ3QL64A/yw7I3bpUvsiiP6dO5MSZPOwj8eakAlDnaK6fq1XXVBqEX8F71z
xgmM/VRJVs2mgPIgaoLf8GXmoRDp3DOOcC6FXF2Q0Iu3KaRGF4frOeYO5QaSpgm3
GbJ1wAwQ6QOgTQ8tmM31/qo9dIMaJcG9mClFRfBshjlto+JyqBdjaG7BIH2ZSH8Z
Nn+vBj2Y1OuwH2pVbJYfGkvCSMGqEUxltssINKNCILsRdWebNZlowQ5pN4amxO7s
0JXn5V6V1CfpbeaUKKi9bQVxej2vnltuoq6Jrqml/8X3bedmTxmmBxuZN7H9OcrN
h9hd6YVHIBtTJMjH0AgQOmMlEQ2nNboZBjddsFwvSC3ffs9Nir8CWs/fxtHwtSA+
8bo8oDfU6x2bJubg1EihEY+Zqe90764ggN9XU6NuEjEwBcGtWSJokgv5jpN3Fy/B
yCbT1qWieA5peB60c2e7kNDCMXYbHQCAFOzQbIzkFgO+8Fen2GbV+bUAVdAYfIJA
n0ASvpTBd12VriyFEaW5JIqmBDkJmU/5rUDU9O6MvsN4et8ZiesxthLSP9jqOla1
j5kpXHOUOjPiqjB0xP0u4O3mVF67ijPSn48bUGTHix1hSbt51MzAUX3WlU46nYfR
5EoMgptpZZFHM1IR8sEEcQk3vpskwWxrjtiHkJaQF5XJXSo6UbypecuQogZ+4ibP
4A4CDvFAK08Rbo7W/qzrdvdUm6/A02AWsOXlj+kFvUN4bE1/3JPokuxJx23zwKPf
skraR6crjVLekazj+0sCbYdZ36vIPeeSIU3rv5JVoR/mtYWJozOSYL5JOzgO7Ojt
1zyw64er4Y0vYDT6whnohlCljb6updQcH4J+qfOXpyVopRzz5k19J8Kun8cv2nW4
X8mjFe1bUgXFfcWN+6Y0YTj9mwv/AnotShXOpCEdPnzTbQUAkhTIGuSaNffRROQt
iPdZGRtrqDHYJFnlQWhZP1kA1RMjaNfTUHkIm21JUb1P19zDQ6yHqyMIrS4Os5k8
mdkH/b3F31ClE0KKAUcW/NgAXER3Aj2p0fKxvIt3uqkiymxacgWAPDV+QzR5VMIY
MO2S2dHb1wjzGIenm59EBNBe6a+PxbWncO7Ub2oIfUUF2xYwcZpy+Icj+OXhBfYp
W8YKgUSMrdhmyJpcW0Y1Ww0DsOKf9cpeTEDxDWPRcNCVg/mbr9TIHCWWi2xDP5Iq
mla4iL/kfLc/hmINg0APtsWORzBQlC7cFFRYTQvyEqIjH8CpBcYY3GIvLRgDFhMb
wQrS9X43D1/vghgvf+reP+ARDOtbF3wDf5kc31uNLAEK00ZSisYnvgN5d6rQpb3D
Vk3UL+To/utVzSb+rkAYIUOpigDiCFZ4oixPtPMDMhr5CIY5odHJSmeI+HSsb1/2
BoXejgn50H54Tho7igUGyV1GwDj3P/7rVuEePbW3pvQAxd/NY6PRJCKRU832l4Gp
HRnC+kJFuYOAot3VWiNfyt126zKpbyLNiB1DmwgjsIvewxNic6LIlVR+QQLJsBS2
OPcUNrNGEA7rvKsnQHzOpHxmyItXWKbZRNhLbLNpALNJcVpTr2Hk/ZTVALAeY+/z
z8Dw1S9KstLOY+2DDITFj4OVzZ4iEx18Z/4cxojAIR2S7Go6hDx1kmwW8FpuvNE5
SUHdeTzDfhI+UgGXE8s+aDR9lVa4uSSjFVmcEI6VJ8FWYDtpGzU5sbT08husfaaf
+uWveofMXAKclNhLg/QdHDbm9zgdrGT7X6PB4zaaKhU/O4xnfseWgosh0LimJmtm
eNX5kmlWMHAtnb7vqlqLQ85wlN9vExbVdy0ofEq/De7tmrr0rBOqoVNLo2p/3Z9q
eVnb3+1GkkzA4n0pjq0CPWEKqOnIr8jK2Ow4SEr5XPrijEDkpOTqh4zVhUj8gAM2
8wMOPReynwkDXzOrMbZNhvpnxxzS1Kw9dn9dHDSFaoVf2fnjlPxgYIQ3myk2U2Dp
LPKe9uOevu+9xFFgynDUk2z7umZfcyi/tuy3Xq12rO1p64agjVgTSqjriroocXRX
ezymVB+0JI6ZVP0kLw/e8oscQdXD39qJaLbsy37X4/JL1RPFzBkz0FiXTPlTmrOO
wC61iFsw55Qd5kChW1WAzv1d6SnQgxj/otcCTkvZQugIwGU3kjflA14se4BsYWdr
P4RVEchq9nCqWp2V0NVfPKZ6tRKHlxF2vQ1YcB+IbcG9CkUuJa+BiLmH29Ujjgax
KvNGK0PpKpfsHtyvkBkOSwUhZ8YLDsVYfjDNrQnApmi849YrCLqtF44mIq/3mdBH
KTlQJSgk2dofjuGck+ibgqDEl0l7CjMMr+xVlXtDrCr0sYW1OW57JOwMkIOrvkod
+wPOskJFQls0EeNxvttKtoMKZxZ/ZVq2hDIueWnCxMXbd0I8siZzv8pwpfNsMAE7
OdWgVsFv7FVlfDhqD1RSU9KuXctLy9eZ50SoAw3HmX8Ob9Ck8iv2BRhHCsM3zpRT
MIHD/MDU7zQ3qGf8y2hd9ri6NS6BXaCdKhMjUyXdcXfBlegcPVbj9GCCkfVrYVeK
magGO0kWh4et1WUnTQN0QX/8qcQnUQB3Ol1KHNGXQaGWcZlYUSUa8FiQJrw2JD/B
O8g5mONJOj32H924aZYT9Xne0pAGY9YbqJQTNwp9BYEdoz+EPTDpoUo/bKxM/mOx
SeH/c+MoHdwIdE9E9Gli+csJoA3DI2eN7VQuXuPutoBavXjXrBhZiMSzOpca8mPq
4FMUOyMyluFXI1NiLngsMo2dG7S1hfvgLWMgGPvHuGYI+K1W1oRz/stW+eZI+DP3
yraVwCQbgBieFB8RQcEF7wV+XhmN1PBWfJgWYmtsMYjP1cWemEUp2SkZ7o67KS7W
e9tSFNIj6jJQwEQaitEEXR/sMIJ9InQaPls/aXT+8SVdACFMLNKj9WisndES5Ax/
m4aeMNtmvvHhqbGoUi7utLjnHzrP3gCE0ApoVWlA6K/SrO7zFJ8JeyeFYBabEM7+
cS0K+FeBqfbKqfAzDdMHEouGSUIy5g8n+50wHt5i4wVXQf4YkdeFntJiMRMoU94k
zhUduILiQXsFS1dMDve33RCE5ECbgmVMdo6+ehrdV9vo5CNvstzAnUB3ih7vc66p
yhBCmoD0kkCpnHfVSyoz5zszl+mWuzReBMU8yw1aY9hcxk5qLJKx0YYLAqWf9wnB
6GsC1mhByom0avmpVQFW1U1p+rOLpGuGxq42oYac/NEpz2C+EKqNSkPHL3zBgu8C
pGyL+b8x3EKMd2MEyKaHL8ZyYkqA71cPnhu/UCmsTXZ2Xtlyj71R3grBg7NL+M+h
HtyE8WTzEj8bbe+vgT6VRbI/EYUbSrfieHLj+yTklybZZ4YF3s7pl459MmnUbKY5
UNWw4xlbD40xq/TVt+KtjxX6Usovu4OD6oo+YJxIzJ3V4HFl7ww6l2L6BqXQoDJO
0ROk4NElnyNxW8nVHFr4PrTP9LGaTHhgM4D/+Nc+ewvJ+9iMbQi+nwNY6OlpLEY3
YvCeuX/ARhE1ZMN/8fx1bNVCUkieGnnqKWocRDy7u2okoESDY5KqpZqHHgf5LAGf
xAxL44OblQ7ILFYJ+t/1k7z5PE5a4atxA3YnSOJyqHQz51iRSfwlrsHJKtlGN6Cs
szP+j1jCJvPyppy+nJuXsXXwxNH5Z5/VFLsWdHDujFdD5Jjaz4UQl5i09DyChQ31
L41ODTDNUz7X3e81uTlTp67kmIH2D0tSJjPmZZgt2bGnfCm2gu4dU5nOhz2rYZ5k
7cHfXjkT2Urs8UTN+vRyU6eGNXEmceWGDQc2IKbQD3o/TMWkwnr6lZ8vm3f7zK/z
o/PAPjAv+yfrPsEMGOMp8MGUdi4rF4r6oiOa13QpqQ7PFx81MwR5XLsV781KIcIN
x/0LYDotBdUUrle1s2vsuCQbsU1h4CWZJJdouEiclRN66+DuJAxRm6sJVe/Nvc6w
o7VqxBoiI3WvM8WJgpI/LKIQ8B8ol0CCzixbGjF/RqfixZ792MiEljOqqXCTVyv7
K0yHZHwArAGuCqRfXD3u0X7K0tOcqTki9eob+GkZ062d+yRR+MNGvG7GiMAqXYcl
eNzu0wcZ/j/iWkQJRgSBNtDHWLqiw0mgacuxiDjvqutJQZfS464Dk/Exc0CNLmM9
Luq6c4fMcsX8ucPs8XD5BrRSYUiSr7WrWKiGBH85vHrnWSq0mHGiX5CEXbk9oH5q
ob+OdEDFYf92ZsnN9m3RSuVLXSYKFkpjiJRWmedWoFDex4swTsKe3NvuTrkP6bZa
vn6lNjoaSg7iz54zcL4q0txhduqz9zs8zSBOPmMsufsGoxALB5YNc9kG70RlA9Ec
HSB/Ja8p8pKT+3+CXOWwteGDTMuN4pHB5SWqMxbYbJ2bqqPUL5w3/93qMuj7OtY8
MUQWnI8QHA33mn0AgLDUIIVZOP84/2oVLmi1KNBTJo2WuOSqRWf9ed327U3lJiPl
yiGwSsnw0fvSKmX6asvl8DBdiinasP9lfysNmx3h5GjSK9xJlQIplq0ok3YFI2Y4
D0smkELa0BTx8gGTa7J3LaCFzL9ojL9USgqkcg5GlpSpIdBYXenDZrRzKBuf9TAj
mLFSb1XW+sYFOIidCKG1M5+TXkPgk6hxFDfQ5B0JJdbH7zxe2tOH4lstb073KmGG
vh4Zt1wXYGoziE4UJOAm91XwhHMzZmMtMEL03KaRtXdSAN0w32v5FQogUjlpPSSs
QOWK1brvzVV+YNeSLIxrEHlFZ69CQW+4lxg1jAWiR5nEdzHa/EpMqZjoBqm5FbSD
fFkufDhTxHVhzVqz3DrOW3V9vcdHd1H2vjI4pNp1VOb/F5qfjGNjpec5Kk5nIKMl
x2ax6MQYiLr3eEPeWoJlcGuZvXYO7mY4kKQzk0bjALynbGMOK6we+TX4jnfnjQz5
WFDU3WD+E5ZXg7awsRahXCJVvRUfDyn7UZdo+UFKwXkyQ5djkdhNfU4LqWxZUgTD
cpCt4RWneZGd5EM0ElZ5dHLQUDam0SAHqs3doKkwY7VpUM1wgbE3N1vtcmQ9KpQA
+4zwAu1pTSdRCNG6EJC5djRcKoxr0Gbccr+DqTvNWGvHrDN4Fh87OPrn3qsNOuHD
EuLn6f+MWd0G9jhONW/d3tZhSKrGBM2XXdx/pUcExUKJkHPcIILnv0KwVdPVoyLw
7oIQumXVp85odhCVxVCmEDQ9MU8xDeaMxyU/X1sYgfXXItbFlNF8H1d1V7aJ3YFq
QttayQ0ttNb4npgdmMDoFDmb2/3JAUHiKsF+IXrruoq5SYU542DymHBrZsyhh+pc
NOFHXaVW/sQQGKGisMS8mHbIVOQSwyrEpQFgxnSA3Gpw8bpBcBwFtaWq4msdUejw
SarpqqHtsRmVHTXHIGkBKTHzlE1CNA0kyeJHmB4KNzYn3+uRXlmlNRb9ARyGmr9S
5xFsxxJzQR0+7qB1t2434O9fBUjVk/l9dEhS4lwkBE32WKhf3t5qvHQmiFSUhJ0Y
d0LXia1m5P6wTAfV9AeDc0zvTpOhh65gvuMtnOyo2scPFXRSQwQFaf1DCFAabOhJ
xXnoRSNE8GZvmotSP9TqqJI9d6+wiUFr+1o7sFwWJAF9gqH1+4BG3PnTnBQDvC4E
hL6/oEd6/gR45PVHgwMEDKgYbLgGUB7cUH5nxZ6HB/4pliRLCRdCZhlGXlcKu9QJ
ZPTm9aA2soL/k4ufeY5P4/KjMn9WnFuW3IQ+E498W4fAlL4mbodSr2t194c7v+Um
MzkcIN+G3QiyZ1LMLnuxRiKEaK6steZI/h8716xv7J6tVTHiXyIRlALVrLoqUO/2
VttaBxgXiy40K0RtsOTQsHvq1pqJ5AriH62zy/psqK/+QE3qOpqJCUur2pIYU0kg
dJn91BCkWZtd+0zKXNsGWW8m7hgXBW4wti/nY5E6mt4XPh+Q/bBIjFj2bhfhrJ5k
gEuD5vgcGe1a2jbbIJ0ac00MjbHBRdcSM/krUYUUrmek71N7e8mOJg5n6HxcJLSs
LwBvtQuRw3YU9eyv1DmAVUuIC6HSeLPhNTVdI3LCuwR28SdYYT7I+1s5xM6GWakl
zRPfr/yZaLYp/36n4IkIgDgPG6SXe4UjRmQ8pWPTCjiL3BuxnywE1T1V9rn7sG3N
hYTuCHhNHb1CrXD1bVxax0vjJ7frWFPLAyUpae0Bls6iXNlj8EIkG8rIeD7Kj/Cd
0Jm2v/yN8yfNu01GVa4jbM2Hol6Ux/i1Gziwcy8QQ2zdP2KvCkJxhlCCknCp2n0N
D5siXUC7bHWlYUJHkxh0nfSduYzojbS0zKdRCOjuUkYMY8/9ojeYrgJecR3CGfeF
VyCifDZpOMhsX94Obn6ZThs6XOExzIjHAry+YuzY5M96IkXlNo8LeXEQ94LQRT/G
2iYeDc92vRCDssNYLabW6v7k90PxVkc7q+utOBUzf2DhsElptWZeckr8BHnzsYE9
qLIs12H7sARTE6HLkyIHLPzo7Z/pP1dqmwtshxoaW/+ik4f7rssC7XXQO68yxJ6e
E9mimSut16yY0nV4FbNQZK7I5ckjdvqm9Rv6gNpCOEEWVPBaQjufH8MvJeO4XvJa
+4jEzsvmAnZgCyfh6OULAwzj9QJ6C4tvzMrOTseerlruVmvBw8IlSitpm+KV/D4h
eOmKX1gc+hStTP3wh9yK4bckPk82Kdm1ic7XiHzRQETe9Csx3aHAFWgW4l6DgHu0
RhwCdeAazyxsL382A6T9Q0qnBuGOH313662PscLhGCe7onuKrZn1E0bGLMhOQpK2
Flm5MT+YTtyvMYWTIarD84IwDvzhStQ6PrrvW0rICWXj2EgS31xlrXmiRVVBsxTU
ALjNFzWNqJX5y25Psqm56vVE6mlAjiwZOeTDI4UtjCjIB1gQ8AUckSOcLzgs1KUu
ExziONrEp46OYT+rv/nilsexbCP1Wf/pnVxMXJLHvHMh6vpc+U52ZUo6wnuaC0Qw
tmMefmgnNsJDt5i1OG6Qi7LaL0uc4wsK4zuXRkLkPN91fNXDH5Uer4nF8zqPiI2b
Ay1RzzGSMCvwbKq/dZ09NGbS3xQtCfK21wWYA5A6H8/jP6Ieef9C6dMdOOjtX5PG
uNt6qc2lZ1kaDZzzD8WZg3TSmqElnyJQqiI1lEIElczqAgyMeE+RXYvqAOsABkrC
11aNx4arDMaAGT2b8eyLtFoGkge6KhB9MeIS9/Rvn7tBh5DUgHmsowNfU8Yi3P5g
r3mC/aMdg61JC3uFQfna9RJSgnZ7pCWcI7iiZf6q2AGMlRWDjmKCvdf/O2IDDjDW
haps20Vo8XdNpnnLxjHAv1EBOJN5NiZse5Jwl6/Ch1HRsKHI5y7yU4uNFBsYUdWn
sYsAuYEJ9oC9yp4p5LGu1FQdjcxbbclgmuzVhOZV5jYmqkgDFoE0XZkzDS8hnyIK
gF+xH2mYHRNm9KlKPMosLbOuVKSKV7UkHQsqOQGkTN+za7UQJLGHkhkqNh0IcGz7
y2oQcjho48uhD8qvjPklPfrBQn/0HIjPqlrMXgdDdoKDcdNHCB8NqcBGRRT85iCH
XKLr6LRdeaK6mbHuP8NQQGI+ootDgdjTaER55/tYk4ABHo+8stIGZ8KC4cmR2UHy
gL0C82E3bE9W7vgR0rT/Xn+0I/sAyGtPZ+VqpV4p6Ll1kll3kh8ehDXdmKVtkQBl
68Tw0bGdQ4AxwzYeVZjSAvmCv0Tgp92S1dMCy9DyNgOUsbN21LFYRennXqjrpEWU
9zxp9w02vJCLqVbJidSxNCju4Ks2EECH5bK1UgnLFayp1q9HNiihJUFEsvfNo0Wy
Zr0CTPpESEfDXPP8vKIvCkv+0c4CiDEm+yNrFkS7fHJxnAN1EaAKVt2RDAr4kXDx
qpxFbSJrsX0Pva9QkGQpI3L4ZuNEQ/5EdwC0pLb9XTGymJP+mT6/qMjVIjiXXr9e
fXCW44fH8tlNteA8c4HuGQF+ug0gX/kMEFrjpJJTiscvgqb2nHnvJ2zs/v/ZK/2W
66s3DRtIDtRG20k7NOAkJ/f6y1RZPH01oKPwhH6dSfrm+TodlaXExfDcXwhjwCZW
hJoJjddg6znmBhm5ZKTBYLBwlje4AjpRgnHNREcoUzE9XVHcksxXqxfkh0ViWvJ1
qYfRAN7T3RdG9PQ8pwklYEx/jy9HwPUBYWuDR/spA48zYqtYVfx7HCMV6Jfuenks
uGme3KJYyIyG8fPSlKl2nRC1RJyFObXgQZPNIO3Uk+dKs+0jj4/CBAPstj+xnXwh
935On/nZ6C/UkYukgs2KtusylD/BlZVjxsdf4UAi2aWwdI73wEwk7zFeMsoZkIRK
B3ye3YzfzBIbpXemK5BK0cyfhFo9hw5QUPh4ryrCkNoX9z8ftIkvsAioci/BN94k
f8SfCRnNJvOlXBw3k+DhD7tjsCDBodeWNBsXKOw7777ZCHzQngYrFcozoWvjhOn7
bTXOmcXvOO2RV4qHVMbHB/nSujqxHd5qGN7RuuauMbgFTHaTCKUjC20hjsnQ0KGn
4owG6Pta+9aUdmMN2cEnf6RZuPV25gnc9wdwFi1Nx2M9YY6HRDgUcDc2NTlFqYC6
C4dOT6KLfOBUMsBrkI0dnCvPS/poAWyUKTrCPDzwOQyhLamZ0PlsxzXmHUUfHkxb
iiBdT9Dg01OD+8KyMPb1lEguI/cTCom0RAWM+VPY0sMzHUArIbqO294LNJkGkxuH
ZkWuQvKksYJnrkBt8uO+Zl4p9d7LsXZzSnxNP5ng0EUTKgCHK8GRjp64bu3ESk9J
CTI4bPpPGm84wCWMF3XO3LP8WqDXcjnzbz0hJo8kAgK6/dF8eF3MGrzuZVo48T0V
LX8836h34prKSwW9AHN9zP4VXW/fu/zdiUV2ap/2jIdW3N1VmuEA49KtSPp35qi5
YWzgp+DYZD5V1yd9mLTlhxgD0gasqDSrkOKjZSwOF2rU6b+8F9ESKzf8XxLlHZC3
EQuQoZFwSYlswPOH8ZrzhjK/+1RKxral2fQofHLBA1E6FXuOFR1pkB8qSdJCuVTx
S9zdNbSp75K1HpNTZd47tUIkot5ZcKhtV9W0BF74SUIx2WmoYXKfeBqKkmpwNfcc
fpqGiYlPlpH+tSeOR4vi+d5K5p2mfj5na+DJxKHR4m3KDe70VnkjLdPHeLrMnLMw
rSEeBQb5QI8KAOqjDyfo+fHHIWQ6KpHuqQhxcR+Eq0+rt6W3qTHOzj/swuHJAfmV
T1XRoqlEL4bs7l9zgXGXsOXlyJDqiztq2WgBkDg9fcPOg8Oci2yWvKZVv/x49fh1
+BF4EZzmxis9RVElfFAqBDUqEhPiTHGOUxSPL8Pgk9XhRW9hcmhGpURBhTo0TErj
seQfvRblNK9fssurX56zcHWzJf//yUEwBf35MM46WN9BlpDAK8HNqmIif6/PsgPD
gdj0oETWz76j/Jgj3D3FVg0/u6/9q0b6rOkpnSvluso4q5srJpFGf8+PXVxiCtj1
Hw2lZIGBo7fWLSd9shNZPZKPxXF5S39iS1ROde8so8oTAxNWagJ4s4aURjlNCNNe
O4klYbjPkn0ZM6XS7josCfMIYmgvobLMTpPu6MDV+zX90W7CAC7SUNdu5NEP4C1i
bnFBshV1hI8rbV9l1VHxngopqVfgT7qa9dEucGjmE8NcoPm7iYGg4ZHBhoaHk+iK
4I016HtQBkVAc6HqErSkHfoJgRNapEorlW0DjBxSpggg9Rvuhs2s6j1/A2QNeT++
3W2DMmMK8gnNwBRk9NabYmyt+92c4pxX23nEIHrYDUocFJhH5BDOX26ISZcf0rso
sdUt4opryVH+2o11nBLbWxvp5rY1jXym62wWAvXv45EdEadT1nhse2jE1xU12lIZ
PU3Rm8LxzxlTQl8B0RSuQ/D2x3OFa4TxwzyxN7JQKJGtjQkO0hkhJihchQAqoQbu
J/LyeAlAujPc/+qxJFWRok6c7bRyRz/WwyFKvpXHEwYkllTrAx+DYejWR5O+Wsjt
N8D9RDdnRzYshXe9ctZygDJ3RSqrr8dprjRM3f+Ff9skQdGXXBMQYQUMUA0jXI6c
a1l3pH8Sh7syvmnqb75MROSVTQs2FJ2xYhFfjj1W/nAMV/7vHcGFcsUkW5tbh5Wb
LO+TaxcFLQb2yZ79w830ANQ3lnhPgoXoxHhjF3w7hsLm2PlqWnBl5S8H4t5nr/jJ
2VdGFJW8IxZRLuHEwpkDxfq8zObRhYgtamlGq9tZoOfyXwY43JJIvhCTnrdli64i
YEogD1oHzw1p/WFdqc6bU2s2/kSvuVifL8w2w5JqNSL2ROWyjuwexZmd2LQ1H4Py
o75VE/KDvhbgxA40+TIZUrKUzTSQBel03piHx8cfKAnMdk2ArAixIaq1ycNEl9fy
afNSIQJYEfOzhPQV/9Bl0MA1TE3U80l0bPn2amcetc5gIWP8c2IMrwMFjK5Q/n+6
GIhIT57VZyj3WNxuBRfllashLMqTAPg1ExHuOP05l67ss3lMH8uNa4BWxNfHsjcf
p0VWpCimcHcSoY1JSVEf3C7rKp0KSuRk1FagA3uKkQ+1HW2CccX8u3S9kheRK0HT
Xo68mQy26qmbtnsw098X1wPvLzD0PKZmIs8pcCc1dCfaViNRqmaT4Eu9F4DeUSMg
LwXA77doULzC4DnmWUjaImr+vkWMBv1u89dGpEDOzCBCQre2yDuhrAHHnJ+aRcJV
V9oewHNzhct3fS9qBkFSEPRYZc9m1tQVxGdl/e8sQd2dq7008B3Lv9Nd20JVRNjf
Ke7xEBsqyc3LlpsA0RmCD6OgT5po020ul5UxWj5390FVMGtvLfWtkjQuQ8cGP07C
y3fPW3ecmE+eVwJzdlvvHNDahzNrRaMUdlaN1/IXt5cbDsdGvgDiyY3fNy+IXJC1
yUpKmnFSmVMZgAVZSYtgENrT3O6GirKaHU1lVxm3TVOHAh7hEkrFhKzDmvqklj/6
RdY4huevQgwG6d3jmtRxx8OooVB0wTbfHWmtrAuaYlC3rJ9NcPx0pxHAjrKDVV5b
YPbjWSPLzd1Mx3TwD6cNQrP9G7QlCcRR3nFWWIWNxQI5u+WrG4Lh9d4uYSRLATyY
ozwJHHayhGgOsDZThSkvkA1kFHFFSLlYip5emlP2N7PiT8OwIShsl78Vz1vkJoOM
Hv6SJ9KdDrcrfFpiFnIOVsb/bkzc5FWuh6pv618fmdshy6PM027eBYYxC5JmCYfn
8xWbxmWY1xzCp0tlq0Zj9rlx8YR/7U/02hqi7ntyXqvQPJX5+fI8PsQpjPSHi6ik
9peG0AdOVseMQY+0fD9C33WEQf+ygVwI7Pg29HjodI6yQb017/SNislS8KT7ml1f
YsDCG5htRI75iPCw1L1pHGLGTrSYUTNvjEnGmgk0GMY4T+7qzO831m6xWkWdZ+xf
5lMGj5UUiN9Y+MoVhFJP0+SF29wegFN/Hwk7/D133b8bWrMzyRy/w+4RkFTBqj9W
rLIHwouF6pn2ek09CIr+820jjt1zqkHkamjKOaCCo8NJoP/ZI0g1aA9bk0bM43Sr
eFI0pQyt9FbOL1sGHf4iiIOwkBHBEVX+mLwPdZGdK5QQMn/dRXTtWWeNDq8ilMm3
HracMjrdXffSxpoH4/yALgpSCDZj9u/evdxHRZV4Hfzcl+ouLsOfa3K/lUNrnFaT
9P3xZF8vYUs+4KmpZwXDizuyALDBvYAsptxusofMJJdgfoo6WB8LooDn0lybehbt
0NCLD2tUCDqG9+lBvKmkrF3Flpafho6eRw2/prfd1wPOX+EjLi7jVuuRvrIHWRXQ
9XRhaPAmgoYfC8cpaNWwqRcAjIHkdLytpISVjDF4g4b/OHhc+HDH0nNBrfoIB4zG
bcKfFi6KHVUddAFuSH/LojUb9VZd7QEUOdcM8sV1G3z90BsYkt0TWS+0SNrHrJVj
RpWW8j6rxH963gaGGA86zj24NgAKnyjGuNKer/0hU4q5xJRJyD+mbHCsnEL5VN0A
w+4/0csCrnMLoqvrxyiFhrOX2+l3LVSDZvkyzlEw2Pm6/KPBiDN3amgo9F8/ZCv4
bDJ4yU1XH+7HHVt9QUqBSFd7L5sfqJ1BoL6HRL3vDOUyjjN9mcpJ3zNaf4HrbiY6
USkI6exQiFTGz3R30D9bLeocQ8V31YiekzuKoHZLLHc7TXoQ0w2KXMFqsjd7BiVQ
mi4Swqlg043bp+19YZCnnezab6oCOuzcF94HTVKFx1lenZRKLVJOtz8nWsw1NnPj
SIkMPTp5TPgs9J8mAIUl0kd8W9U26b0zOIH6QRHb/v+Z0XA/gAGhI/rW94rcBgcM
Revs2OkV7dQhlN7PVPUeZMFPhl2U57fk2saT3e8Zbwr76LZN6wa/oFKMdKyDmfG+
AnInJIhlK40XKb2Kofi3Ylq/3Xm3U38ucAmCWsIdYwjgu46PHfy5nCNDXTqG91dk
65mUmvXAD0vKBROYHLRtjgzr9xBbQdfIbVmf1FdJYoVkcp+pm7yX3x/XdTUFTsl6
P/UMVPCOKjujisGLZkQcz1sDVJKxBgDEpPR4ce1SDcbep4Kpm1pj/S8txc9Tpaoz
0B9ZbKjUVEwhkW7Reng7nmfJisV/NBDPL+MVXyY6RLX4O1hduMXeIEV5uebG8yBn
3JreKyR96jUGKscv97VtTjv3fXcnwHEFNkFwqfYgzSV1roYwxYb+USKIYeLSwfGN
4SN/5B6K/OeQH1H1U8gt5AJm3aVzQT1F9rHTJKK2jNQssXnLjH+5Tzy+DRdrXKDb
iTd4+MUu0+/NW1oIQdGEg3Rp2p2x8aBxuIWq0TpLKePSdRCdeMGTTKZSzf5JX8B2
6QAdI8mPAiFeux7lNIuM33kI8cA1F/dq5G6oSLeUA7gQvWfBBhWbxaIBQ/GZYGsH
SDULYKMBgoZVFCBpy8WiZiXslnCuy3hY/xIvA6PLv0qOOebM0EQWAzBjbvaQwzij
BnKuSF6ynHFtaBQ5TKixdHKck2qqBABbOeiZq/hiz0oaUBA0S8p8WIapZag5avwi
yB8KzHBiGvr3w3XDiM7qNAKmykAP6N7Cfvesu8Glz0IkqUD9tQBWG4fkXkFu/6jk
4M4Odo7j6dgfadd+xe9OSctHfpq7FQBpB24rPSsoSzxHPC89XNRn+crTtVaSrp+O
vbf9OmSnrGQNWiqZ5w0qS8OmR8OGoqDWxfGbVHOiBhBPnEqV8BWnmrLnKS+HdiLe
oNHEOimceadxJpLhy3BUoCw9ip0zwU9mQsY26IPoCOX6qvG6ZLqEGtcSYqbRFtNV
j4aSpafRYRGJBLhNHaPW4buacdBYWfCp3k1TGERIvP0qKNpsjwUGYE5a/76m8XrA
K/cfXk8mEp/3M8EVAde/FzyQKEuuuUnJoxdSlm+bkj1gTgOBtv095Ohl8Ae3EhNi
w1wHOXAr9/KLN0wBrvHPLka+pw+REbchWfcP1uWERGkMUckKWcDaXK1n0ST0p2TY
cIIpJvfHZqW23OuAcp7ffOUi9/0jZZFa59f9/+nkQUE421sQyyWxfr3c+bk1xWGH
RR+WGvcgthbtltgfuhRQYcQIZmA1k2Z7GPXyMrfWVz+LzhZNYOWtc4EapuzZ3MC+
7JmCQJpJxU8Zh/qZqrcsYGjJkxmiB0E6MY12cb9uDlVL0KvnIbQgN8WA/5EfUqcm
McHYlR3Yv9EzX4qjqjg2pUTQqer7IZOkyU3M3J+cZfRtH8PJl1ZB3r7CjLF8XBLL
hshA0NooBzENbOvP5gfvhAcD3labSZdtWGjPZMlb95mAfytB2Uu/kb0FdJUXxm7f
8nZeuuE12YVQ6K3ZsoQTd6/iLmXyHb3x4MgiK0ZcKTW4fhO/IHJMFvursYmQ2+8J
avcmsEhxFyM4STeaQvD+RfiI5Fi9ZESsKFiIwQgIkE6bYuWHgUiFe/4ANBGKRHCz
H9I/GmKRTKd7tnlgwlZ99MXQq/2kgd5OfmoKgqdjax0zj92zR66PynKNHermL9iK
tPD8buPmarvCo+4ylYGvi3Rcby+ZFprwYn6zbzDXP2EYpYfmND9Z4aJafDdoXihr
Dy45fzxrHEkMTYr6ihzoowExnsxhRAH2maq25ljhzfdMIUVGf+M+OHR/rG+P1IJ4
lG9fGUhGiBRBVvg8Cb2QGV0ctFdMnkU7YKkalZw98Vs6TVwdxr2TEmjFk5EHNsiU
WP0Oj/PrHL727s99iv4arnXyDt98ZX/UK5DgskPQ1DcrSUmTMvvqtjn9yjPEtnKB
+b1lxd38OEgAO52bdKY8zGHPdM7qhA1W5xjl96JKAI40VhUePt5ira/vVv9l4G6X
W7+CBo6l34ZYrn8z3a7dDVrhDJIxq4klr/tY+niD4IvMIKFXpsh3UFhsVfqKrguK
0hjexKdegA1hjxPbdv0dNEuMl3TB9uAfkd50yeeOEEnt4n3v7KQubP8pqPjrSQXf
gBWAMb9VKPoQlq89a+Mz4enu9F05m4AyAo1I6/50mckA1bSKKksvuCxkOrHa0ZLB
zzNdz7NQypmtsnGAagbfCDXntLDIK+/g3T0+3kHcfDW+txAsIgpkIvaujOyBA3ur
xIcO7r6mv5PXXJej8/cB7mu3Ju8ZWHzfN1c0bfIR9jLs9+VNbGGhHgm1vfa1sROy
p7m+Op+s7MEuvl9+DQSZwHjeFkZxow3T1veqyBEk6gr/lMzliUIkuXCuEyeqNWFJ
3QtfpsVJEsUkHhqBQrutev7tUQQnvY4w7jujsPVmpIAf1zeAEMlKE/IyR8Xr32ZY
X7a6mtGBzBFkx0GrcL2SJ+my6YNZA03vZ0e9NjnXhaaTafo7RrnoyEJX8cppW8LG
HX2xXcIr4kjqbero73D/u2JcfOYjgYdUZbUQW+lBN7sB8ulZ4CoVoZ1KIFe2qvUU
F4z+OksDPhGYS2nUhMsFRzYOyN2ix9FCvkvMrOubzX3sCSs7x+9LwsTdWBpyqXvW
tbswJCW5sPDBnyAfzcD7GflVKzEGZuge13fblekluohO/Q6xAN9mORPpaD6iA/Dm
6NgNvzE63Qa5BpU7+LoB7V3/syt3W6XvgFaOmIwrO3+knDEzjN9rKmI1jigLFiC3
e0NeoMwHx0/WkgoJlidbligKWiBAd/P7eNVKsfUdR9H8/B9e9YwAve+01egvayeS
OIgnJi/+97AJs3x4arDqlAafRtgGySA1+n3nDv11/OLJNTHrAtmoOlguBdt2JuYi
o9zMcsQNw/rUnH73IvO3CvUX9epcAp9yOkXcpOC0Gz4KfHqmaf1BVdNQ+SjqI2Ct
NLtG8AFRJFhZ1pInHHdz3004moaL72hLvmDEsl/TQ86cSngFhrm/MrVgqHzgN8Xr
HXqfJ/j8uJGoHB3YIDz746QqwxxpUmwfEb7lvlTGU4D8OToCFeFF8kzaOZXpiMc9
8FCnes6MBxDI3bBM8CXLu/SBaere+WEeeVC58a4jFFliN1rIxeSfRhhxeS2KqRys
plsOP9yYDiA6lnA5R1p9s8dywlWVS6fHSPGQz2BGFOKJm3rb5MJ6dGyvrTGCeyp8
zNiFzKXwJdw0R0zZzLjJ3NhgTfDaY50W4zBj3Yix9/bndXI/HuHqQJL+ZBTK6FyI
Hw7Fyj10MEYyfwJs+9LS7RxhICOr6EXklxIFLHZCY/zUwYFbXH9+jgbjUdaOwxWz
D/NXLKvxsjauDU3pTI8va5s++NjHNPMsUCMog+Ryh18E+PirKPEdNqRbV9X7Xdah
CarawgL5Akz+shc9pa7pSLR/YJ8yMjWFeFcddSQDODwX4orbCGoHzd0XqDJtY8H8
PqbxF9a6ME9/tTPaYI4t9xoog5f4RDzX4gEyUzEJySA+sN2NcvcfNxy/covVzOau
R5fgl52o36UIj1C2mySrl2wEE4ROWEJAsWYUH/N1jFUHevBWn3c6Q7btSLpZzkJ1
EEGJ5li8V8C5b0XN/5z3E0lwXHtXGXuCjtzy8dOzstRj/oS1QRLdrjhgwzfm/0dX
HO1xJYRViHIMga8KOzbrd6i4sa8vw3go8YLwQyZjNtmNNBkXxz458bVHD/LZmaSi
lyfa78OkqCEW1gRzi+feRLPEXRIC5NxD3fzyTMEiRJ84HhZ4cvnZTet5pn8PGSxN
Hxz2trONB3KnTAkZs7X8DucM4/1QCYI1oIhO5bPIeYoSJM41QjE2a02ubKR6jPnj
Vr2+0WPzPsqogL9mBn4Pd9rkWBlF6xEF49Uj3iuHXOzUBOZEBdAfUk0cVPiwCWeV
Vk0exAml6GkhnYIl1X0YZ9C9qPnjV7hd2VGg/VhUrScNDFek7mLZ2zqp/PMbxPTY
I7K7tljnZ2d0PlqJOStp6ilqmcFQZHkZjtuL0+QNq0nzqRbVxSoUsPERPgpfvaGO
VzMWK4wktSXTAkRWIVlriKjDJ8VTGt7JTMXXBZEterzD5TUaQ9Hu5Smb3BSxRhX/
2L5/vPuzAnTpG4y5CD+GONzu4ccinGyMXIjEIjOzboa3GoZb+FzlGaTAd9aucGME
ig4L1NELTRNAPLbrn3SYLece01EmhFQE5u7Dx91OsxFRyeegYge7z9doQ5qDIbX3
Siahftq690cJ7Pc2Enh94E59DEoiHYnHOq4FYpocOprazSODr2Ln8vWHowX/bog3
T0Fq55J/ZyyLwlHOZORQfno7BNXIIOhWlUB78qXt4ATUbVfUpxLC5oy5stqP0pQM
clMBedBIVUNce1NTRT2Whzt/4Eglo0O7MTWundnMOXmSYHVUK5TxzMXdo6gH6g9R
iOZY6IERsdjND0ESABD1iVNstQ/0uB8hGYJVYZ/cSxOJPtxXfXpsrfqc8j94Xv75
3EihAMZsTK7MrUXzuIEynEiYY23QPzmT2EUZ+tpbehvNgt1PRcU2Ndbbt66rR32s
XpFRVoaQdqG+mMTT1R0P5j5J7G9Er81jbf5ScX6xLRoutdceejyibtRSvuJyMhHa
JUXXH50J2kx9j2Th5riBxFJtp75JJqJCNi1CblvAw1iULp67cZCn/KerChSozHPz
gh2gTzLKjVw5M/0AxzoReSsSFt/AuO3b6bH/5ESu1mKvY+UmGOJd65ZSpA1O6PoV
Dcwi8u5UaLoxCnXZC9M6KQEufUIhrnRwMvd8jnd4ZLrGWWq23xu6ucr3PlP+b2mf
RWBwKdGL4r2l2FJx9VF0L5abcZCm0Icb1eK05hwg0xlz7bKrrHAw22F7Aec1y2tv
jVUm7Qq3DOCDNGalp2bfkBKI0TyaDgmQS457G1L6EGJr41HGLTuv5xRvgzIKq9Ku
YTcFlCr8V15LTxGMKKxmq6gpb6/uKmYBKSuvwIX3SltJSfpBcYKmb1ZuW1buEENk
SUhXcqOD/N2vUBjpXq1R12Tha0myIDL5lyRkPSlZuxaf03QKAEUME81Nt1ZXDlX2
icjISxihirmnvcreh2HZT6RmaEMTcsik0AYSaPQfZx3gBSFGBnfeiPXo5CxYGdEH
BTVSROVpgQf++ERmhh+FDxHjHqjhXgp5VLNGFbXQtk1kFaitC9iiBvwzFBARbdI2
lpxQT9OmIETLxRCwUPFhpBUcP17QXvVqWHp+WpOhCmzJeBFJq9Ck5awoGJMYTJUX
QoLNZnAbtJ31z5KZGOSzpwIW4C+b2v2oAK7J8piOtl33jCtYg/c8ZEVeLztvzScu
jLD+zy1UryYn7mKR/5YbQza9NU/iIBWge1uaHAywcqUsmWrmCUUnNVmH0sVzDYP9
DGdxwejdlTZLaHy/y+6PmZpyOly//4tmHflb5e5o5QfJKopVT6BTmyOuTG0Rh7F6
0rIrYB9U+d4Be9C+9/RvKOP9FuAj+jCYQjSf2QKEMB2NgStJg5NRnwMg31PMjp+O
1VhFTbvQvivwCb2Po0TAObQowiC601AVgjSsDukd5aJzJkWTZ//NACB2CsAaGecn
xq+6v98bbgPmb2N4d8j6HZe/XbSL19hggPxFSa0EBpgvtnVc9jCgQSbzhyfRzegw
Qvf/IDCBn9FgXCKL+dhdvMJgGS94BNrCavxC/16zdajjxQKZAcVShlqQNJqcFIWt
E4vFPFo0RxtPOmcO4FtaS0kKQJsNmfKyFZJHGqbgWIzG17B3r8Y9DkqoCihX7RAE
/SHWDp/vD9XYL7/8yak07yN+cPF5TAXt47aYdrfc4tBk/E6cGbJ+tzQyGHnKRvss
9X5I2/Jl7U88GlZaojNPfhX4pYvk4jnlE/BW2ZAQlmjgYbyI2AKLt5wdxdhdm2pv
09V4ruX0D3tPcr6xAcCO2GJkaoeDIvwpSxwQ3ZGGqgbr18kmilcHS+OD5m9t1wEJ
uEp6bmz6lAb4bYjqyO6O2w8isaF8E2ys1c/P26GA0btnmaLbcsIBPXmh4Bp/pHSA
XraDAe64SgS4uMXLKCkFqEkAodmr2gOGdxk7Hmg6cmTWxtU3U6bc2RAyumrJ8uw7
nxLDurYOGR+iQE88whEu/0AmRBt26KGhwYJiTZ2rDNzy+Ysq1xbXg2SvTih7n6Bq
bo1eI0yeU+JfeQ2oZoA6ybqwiKhE/XDRjP2npGmbBDqOcOll4o5fJLP92/iNpZli
i2ZFspE+B+o9CL0fiSxKDXMAfJ48MspO2z6oGDLxL39hdYpDGd5NJYrbB6hb528r
SGfw905h0bsONI/czaqppyVFH5hPU2nt+/ZswH703WQGycZO6Iw0A7BnD/b2nWuQ
O2vXUvpxSJ7ja+tgxkhH//oaAU9+CF3XT3usiWpXRqKl7MCDhrbODKZKMHVMVqt6
6J9cVVgyecob5lW/NTwAPDOsjuNd3UGneGxV5oaJvdoYb0AbRsCd3gLlQvGMd8Rq
W2BERQzaRQp0c2A8YEqLHHjlSy65UjWmjCMaKDXJsmLupg9xnMR4Oq+qyZwDXo4P
lLaTBOgv+or5q9xeCClIh0WRbG6pOyGtGTDHLQRFKsoQio8qRUVxNclY/G1EIFPL
ImAQWjwRd7242qE2MipcOHcPD/yiXoo38nIDuK5FOEYu7a+Mb8z5OV9zWys9TL0r
JdYD6FzQzHkRio0kqq1Exana+bJM8wXGszEP1Y7YSFQ9BVeieZtjQqE5r1juRx+T
PgcJTYO8PL2cfgVy/wWGJqNHxj8R2akgFaxUegSLYVDDuaHRPJvwgenPQA4OSCrC
e9TAe/lVya/HNVizu0abeMZNvc8GouVAGAhW0Z3fj3VytLVWgU3R2R6/SOEkuxYD
d9nFbVrJDAIbsuF7RaSDSQ1ciho0nIKomMHQCC/kY0JVLykeu9pnhxxoEH3UDeg6
bsR6n7myyH0xivlj5qKZPfUKZHqvPTIdrLiXP+SunRSZNmi5u0EcLFoMOwLq87OC
xDC0icNZVZDXkXlzYpJjbRr/2xZCAbOUQSj5Mhdy7CBfFjdn+zWzwg2CQgk6adcu
P+9tnSuKuQDG+9SLLYbQnMzfaw//+Xa/PWcogPENHm3vS2wHhP7IoHHpfeR90nPx
dpZIP8YdY4u7eUFO/8MEUPqLH63hCyPS6Jyks7VhjwVfZAfN9+BFx5Tj9cuqj5V8
I2lfWsjGVA/+VHvmTkyabSmKtHESGZUXQkYhQD+ddt4MDu/dlMTlprsT1zoDkLcJ
qyeQbw3oPbhfaEZO5WHTcbN5rmUCJoEV9CDLIZkInLVPSL57eEK4wjowXmGeXwtl
nYu9jkM2GlYfB5Z6bm0JihyzoOP8kMJc7/uInwD2+P/ZyCGF0AMQCFT+DZIIOhTa
HtXVGp8efh2n1RGWr+TCbEPP+HUy2sLFrgL4UTT4XIHhMmcb4pGfjmAvcWrT+lI6
BqmF8p2baDaTNkR/b/TWG5Y6vfJ3lf4px4wqHSYmcfHxj3pWIhQ1cuAQk+95M5bA
MJ34TqbOeqY3MgMvBe8PkJu58uMhSAZXrLVfu/+ZQ2oRRMfHzRKOCDkkTzwmYXCw
KcmE9C04TKU5AhRkgvepO81LeZRLy7mugAaWt1Cr7cCQDi+W+yzT9rUzOxiKNaNR
BwehWlFkNTk61LZbxsBOZ2027WW/qTNbk16HCU/CtE+MDAQxi064MfrTL6rUFtni
/ql0jAkrCcPFa/5qdqcYhN6dUmOie7X3wieSUuSDMt21XZcjES8LLbdtyPT+aXie
Kn7mJaJTBxeJ7zVtk3A9Y59W+64gWE/1lALgO/qTeKrFedgvVSRCDc51k4JNxF51
GoDNM0QmMSRXEIcEx0Yr6AP4cHFrx4VBWn63bUC7JN/g3Rn854mXBHEmemBWuBVi
xhM68Q0/WrhS4lq8W1ZyZ3p9ZLAU+kG9siRTUfUuRX+VraF6BkbOohi/gN6GFzJX
Fw00hQ2k7Zjf+Tqcjrj9AfRuEhL57olu+/WG8ciRRLNM0/jda4uKHBdmvsQP8O9k
w76Rlc0ywhqC/f9n7uVrkrFSpka8OQ5laWj6eYVgASu+FDRaJSf4v3LgIg4mYLV8
7JmCd2ZumESp4kFg8YtC/XIQ3Q6F3+owgOyMBmREZ9/+dHE3i5vP9gH19frQT/3N
buqo3iWd3hUBVEdygCoewIr5FmOsqh3injhUcAQxHy5dVrXu5OscbUWooZsJNNxA
A+mo92//n4KkaxH3V1RvJSgRFbQt2oIUfvm4DnTPZ2VM0pn4CleI6610D1ntxzoa
/vt0YXlalaPyYg7wN93xsH1I11omRs2ReWq8icW6Ztv0G1Py8gEmLnlb3u7RryTU
Kp9z5kt/XHZVoQErLB2U+o0NEumNkjhdzv0zvRouCK7jdIsVjuGhtH6GRIAonYbl
PO6R2u9ec5OsM5d/fZndciQSChSG0yXar0V6C7QWjlcOuF4QwLgFoswZXy01Pn2+
RDD1/spHbG952TilzkYVZUfaGSv0M+/T2+xaJXFTnzl8Pqxb0UzM8kX3a/R8wVSV
5T9jTIqoqxqwht+NnS4uIlww7HYm4pOtn6tHsg7PG4lZADbkbgH6PoggP9En61ns
nQfjTj2Nv26nsBOkPIOdIRkrwKQD61oz5opMOApcsx772o6OHwYO2dn4hm7wpaHy
ZBKA4fGQZkxz2VVhWmyhwtQsiJOe1N9XfT5ALIXEGWFQjUDMPGRukIEdIjz6UpOO
Zxgjt9tk8Z3q2oODOuvUkSCfeXHW0lAAneZeiyxcoBMDd2E8i4x2CnFN6U6gYifz
hia8WsWTpnoJADm1YMyZe0Hyz2OrD4qGF9TU6VINHTVCuo1dNOFujBGi/abIspCW
0TekCgW0veIFhYkCZPm4VzM5+Y4V0swBwOqr7Dml3m5LN5iKhIeZSZ35EQBrfo2u
CRkUHMdVeflbbeogMdzJLKTO9AYKGgoDPfRJ7xJTAsmgebaH+claKvBRkFYWPFsB
cBkChxbRmGRIKPoz+CcyunByBsQmDhEjBM7h3Zk6eZtXruqDzoHEbbpw9Tamyk3i
JayLxkgUUfGLBZ0fttPP4tARR2zvmWUE/f6BFsUU2RVRGTE1Yd50wTTJ0rQuHfDE
LysY8JjxKqnkaw44ftX2LRXOYdSFflMeyuHOGDJ4jRQZ5NffV1NR0WZeynhSm6r2
e2sd9vGmnshBIejyzjiU4bK7Qp6vbhpvXVXHM6fkw8/YW+263IaojjtsNi9VwkKf
EOB2KoHszasjG5SoyHWK6EfTB/JHSShEYWjTt9ha/3f6HCrhcm8YXQwLTMCl8ScC
hBNk0rpY7Fo/c5nF+frTnc7atDDAS0I2lO1E4JctzPwmuhl+1Y186BwIGqRyaIy2
j8MGMi/2M9c5Xl3SkBdk4CLRR7o5hiJEw5pJGVQpJ7snE2GDWqr/FEQg6pEz3nHF
eEZP+mk73/Zf0gxcTsAay3mGyqQf0TXBT5+y0CCoye1WSFZaPEmKYLNUDxSgYiFB
IK+OxV0EufZF2QA7wB1XiF/JObee94zznUF04eVVRkQAvWUhyn1M18e9yafKqwCe
cS0Su5nvjuyEi140FI56JM+6eHbuQXfCWVciZs9DFRFopoEZE8da7PYoPH7He2Zu
crr/YfW95gjCL2EZ9f+6YE80MPiQa85bn9fvun9njdmm7QhePospTvhgyU5BOGvn
PaQh1sKl0bRGHvIo00Sq18zpGmTk0dF52P3mSTw5pBWuVHIwKMCG1cQzHmt5AndG
IBFrQceEm58oLwbDgIv57nPNeBAzJjveMtgIwUyBlOaO80nrJl69gZueXqkDNd7a
53MGG1t3jc1g6UtMeoFfT8cjF+72qVnkweUtCN1D18pBqgOLMgVCwhIvU2Hs1ORy
cmYBbs1NwXpCfwHeEKwr8UTFHdpijqNS0/8vjEqowwcIt/ViyTphOctBdPGONkuO
gb54f4AFwBjOFC50nWhEqGvRz5lMU33DXUBtePC0Scgnba+blxbCpt0x6wJSfNqm
/MRdNSGfX4LDILOBTtGaL+3BFa1UL8SDvSixlxuVsrfEY+B1Br4t6y7A7nj0INX+
P62wxd2l+t3DdTGQcm5Rq0yzC22KvQ+E3h19/WoZz8qS4wA5AZgEXZKvIIQbO4zW
t+sV4ge48WRRDt6DvsobXj/RjeAmwU5WjdZvs8CD8p6Juzbp9dA6wm2CRNd1Zex5
WjDBDREpcsVyUi5x/p/EaQrT7nt6qrF2eqAOmh0kr5VvYLk3Tmlwse/ZslZwmkew
1BhtLa3Dv8Rev7NNaaWJ9g/agnJlMxrtcLWfSsmtZXFx/zneqvfcJWbmZ1EyH9NF
hmBWTncPExWmHYf2p/cGju6bAR/C/thyTdby/Ebml9Ks1PwXae6SbsySugUOTMZb
wXWVtVJozHVPeIpXS+/yRZK7MAz6EbUFRXIn5KnVODqvmSJlKDpI9rbsaBz/P7Vi
rmmZbHHlD0UVEaEuWltM5VFS6WOYdVA3gWbgdiseP7pngNONvEx31uXogWlUxGQG
QuSd0vojfut2Ot58jA0JOPlJCGUzjhLYEU6rUzYtIgdB2TARlOHtRG3Mk/hBjajI
9gPQQetLSHRZfEnHyvL0CgebkBDS8R4Ke6h/8bozDRDkh/yLRBH50GxeuSBy1+ZZ
3X/QVKCBv4r1k16UtEm1Gio7UJxwCas7j3l2eBZheFuiUaCCwdw2tzLqO0RwFJYL
gVcSCX4Z4Anzexbi2YEQQM0NzXQMe7N/NaIOOeNdckHLn2LyFBz5Mjy/XbkmBuKS
GP+Cp4xdm2XRenCnTk5g2a2NmR/JbM+vBxHBpvJxXwRDLm01dazDU7tCURsEWgae
txVGY0p26IFypJNxvVYB8b71TVwGKWCcJAlmtIvESvORtK4v4V9ZxMThJGsNAgaH
KRbomnnIgWfcwQgue4r4y7kgX+R5iiVGqC7J4xakwWkMPk2UJYQRx8PaiRTo0ov9
krrZ6q0UOgXQpMslj2UO1QmnZ+3nPrN8zEx7ynhDIUAKfrOAvGXTPvWbvVfo4qzF
0t0/KeDSwKa0BCSJ3ymRWDWnNa3hINwNUkat7EeIS88c5dSHLVmL7LeVqaWWY2hk
zmAQRiICob/tksAodepzvV1FQLzWotliLCUxEXYear9z5ajYXCqpB9YRzhUPFCiQ
Gd7yEtdZVPtJP8VOX4S0o1iw8f7uQQVs1melG3+nnT1ZuLZ1f05ezKB4Q4VyujAE
wJ6599KYj5CSDUBLHIa04QwK/W+hYLBWVrDVfnqTb7Mb/h0qNFUts9/TpcYuJTyA
E0j/bmUnBqV+XODNK9WigIMGubQqvwhrCH0EQccL9WnoSb7dv29fnEbjqNFlQpBX
MkhqscN+8bf4y73aN4ZQY08/5N7azihhQPcY3FKqd7YXArV3QY1QhmMJ41JUX6Rn
04Po0mGbp+idV70fCyu7fK8vwx2lk8iJNRCh6aWQ3//UTGFkmfaZ+6YruzlOQi4j
u30bkvC0GsLQiqiBPF/DpEs6bUZetFG+Tsk+wRNnBFuyZU7XtusIaZtQ+Zko4343
z1pribLM6aDXmBybkMlprXRNEmb+u0vrKESTYWvWbMMel1rOocu+OSw14B3Qr6/j
Mo1ie27PE2UgQceXfmoMQn5BygcB4sTOhq7qRSGzPx379p9p17uOciQ6U1zSWXF+
eFb0u7Mg/RmFoEi2KzNb7knT72gezcsSguL7CNIL6es+YABAIGY5FvcUoj05XmIm
dJHV9v55gWfytEn9zUXti1Fz4zN4yhXXXy4LQVdQKhVfoyk8pTZ6DGOJANcNTdye
Lh7CbCxwnYQBhj37/Tl0l04ILc/UWFakdIXN7Iz+6Qt3TIcV5VhZPz9/oiGgg2Xm
dxiCaIZUCAqGiV/7f7GPQrFq2+j5075BGFH1NJuo6Rs7LBs+27DfIaHM5cBVQEwy
BFckSrV1GbT3b/uHrvlUMWezFDnWHI7wp/XNGmZL9iaqyNL6hx1S27DuorC0yEss
oZWoFOSohdQ/RFVmzkzU2Uf6YIz8jwuzWJtf4sdqv6vCPP1BEQg5nOjpKwMlMiaj
VQ2vPpjJ2wc5onJ8B+3kpIS5Fz+8w3detH+7UNynsGMpFGfm7w2XDJ4WNzTKIYHH
32hnjtcBVz6rGmriHOoY1up2ygNXxGf6n2PcNLXPwy6ZfUfpXEr6pzeDQysBh0h9
4zExH+0k0RAwqtV9w2LmG+bC+/lRdJsZb5XaIZHoeoFTBG0Ll9M/UiY32/SPHWV5
7S2h5zyHfa2bzeVRDrEKXuw1D3JCZIdHdiba90oJy2oewp5pU5c0c+g2qBOaP0A+
DwdICphCQyxi9b62YxXpCRnTX9isQoeZo3snROx2NbUakaq1rPRrBXtcpJthIHTg
81/0OIypwcXaiT53VGuO99ulBYrkUWamDyudbhJTPUgT0VV6hj3lc452fsd0jaKO
QAVNdAFUYC3WZ0h3hBWL9bbxEkDdpYoA0JHNthBy+4Hyf+0/zZbitx6jSp+LsfHE
niCmAHwvOmiTsKcqMj2Qd7stN9/o9cfWRsw+2nTqza+HxG4ihMf7iOgp0up9OrpU
LoCKwNeaC6Ujn2VPy7+S9MmITcVx0R9eTuMnWKmPYQgEfxnxeyuOzr55S16WF4s/
PeyCOEVntd/61+/JhTzo/ORNB/Gc8As6xD31guYxh11yuu+kGNfaihtra96P0gS9
BiJYVuhw140mCwW6pHm98eEGIxXRDVQ1CbX31K3ppLNVOaWvZGkBG1OW946bK+UA
gxYDPi72R4NRINVTWbJX5ePQQ9XE/fYbFKyXPBD2zafNj/ujh6KyPqicXOLYOdwJ
LSmosDQZQEKVLigzKj/8qQKsvIwBiwWH6aTKZ6ngkaxcszTWRwxQ5xOghwWju3Of
taRwvPPT7YvKm+6N7d+ImBwimTc03qJXDEg205I0QaRf8dKN8sTguAvrAEzoxTsT
hJdYyx/+HclDiu5zOL6KsK52JlNbBZ1+fvZ++Vh2EIuNO+wmiK4PynX2NwL+vHrk
R/fSFuN9C7rd0Vfcdl6Tr/TCP0fPqs94gKexF43gLTLCtlW02gl+CcMWwBtxnGxs
VqcsWmyngftf5Ps2vqsZZMhOwTffaX552iBbWPwVLGB1tE1EvwsMpeyOnGv5Teb+
IXRLiWec7+aDXIZpt/jifLb5Z8qTGqH2+zkz+8fKemr4a4v/MWIJSB3vGhdRKrIU
Fo9N/GjGYhQBamcm2Zp1+fnuxCA0vV44Ix+pE6sbEQIEKul2flQr1C3qSFyTTvne
he5J1SB0qEkSCT/wMoaST8RgyVIBkVHcsg8UFTLkffx1tFjIlASW7vtY4sMDwoqw
uqwP/4KPFJottpGdLmy9vPPE2rpVJdavix6/Fy+0569vq0/YDsmxjDQJ/nTEXjGn
K/MXFkKcMKXcKsmuT3Vbn4t0xpEWbd0t5la/CQbXkiuqGncHn0oxO6UhEPLnL6kb
xsmR/OQYsAW9Kny/u3rUXTjroIqohSDQwqmT0bk4tVu0F1W0XOFOC3GM7ZdtQbl6
xhjgjjkBpkEuWIx3r2GpTGFsunxz552XSKY1WtP0LlbNSUt7FjnPrPvhko83VqWZ
9vXOaDgKUw5x2X0P4CApTMUNo3UOejnW63TiukudbncyEtPFXmPzRx7rlwJjFO4c
MGduwzrDzoPPABudrNKdP3a4L8gY0ZgEdRrqQ9sCBB2jnJNKaw8IjDP+j86BN24o
8Y3njNAbUFjzMPx2QoFvV4IzLD6m5hoTBp1Zq7xIlLyaARdAl8gm5OqLck7+qaRC
9smH8utWcmERkZ3fDAH/iuU2DOhMuNuxi7SE2n0bbqj8zXBAn2sJTUyApf9FwDw0
kcDtFMW/gPms5YMuRH64SmABYd9P619Ofc1AVm9qtBRUTrl36BENZxikjI51Iivg
mcqS64ktHLFhbr73WzXMuHi/mJ3PhZ1wstg2PmjhjS9t+tNWQMXRfrxMjb0ZfXxZ
RLA6fjQKgkxye2dYvQvpezM08chMed8csNuaQ/eTucN929ep+UxgIqMTkEnvW1VI
QwGZXnHmwBGCazK4bW0ORflJAhBxp6w510HEIwYaWZRKkMGWtxWpHGREFeJ/XM0G
vIA4ZbGBh3GRc6KP3N+ZBueJOoaUK2A5+lTcdYnHGyUQPk+f8T5YfeqxKf5blrVZ
cCVBya6LHPsnS/dCfzRJVqrLFPYxIuvvAN5E+BJpTv12mOVdWYXk7sJKemRCJQtc
PGcQHK/9skAbTMJJ54Seltb1rZq5iosr3FhrPTYkX7bVnRzU/JJdZcysR1Sbs9J/
pgisvCANqYcc1pQp9WZfyC1YNztPjM/KsgZ/YxAJJ2SnMxeiLyxwXfyC+8wNkHYE
ttd0aCNgsjiBbFA6u1v0obH97d9wynnS3BcTSAVSUOPh1lxzpPPCdnmvWir5nR84
ePrPg9jTfQJWtMept5uYOxrtrVlmGy6eQz3dUrQLRN6aYpqb0drSPlhOraxrKmOf
IpHyXo6D9xVPjE+dF9vlkSLwAUUA4iSz4nQGqR/+R55rpJ76RSpfhlRjUf10TYqX
aEoKwaBN7rOX1XAFgH4IlJ8EjO5G+Eml6w55ozueRQw5GZ1/ipiivQOjNP1rlo/6
iulmPk+DY/c1LCEotIbSxmNFvELwGNvUcVM1wCQm/umbOeNzfXTocGX6qV/gdaBp
swTbbiA4odQdLFd/sLhx4NMWmwvyusECDe/Y+pZTsI3SwmUbaVTKn8oCtAksS2+X
DOpejC98Kwsu3uHejvnguybx2/tvC2+KiG8VfpoNtjX3WY7qUGN8Ec+afMDAVlFU
tLIqA/JmlcS5XvSHWWNDNRMQ6x6Hb2xbOvvFSCszA0n4S5oQ7zvOhFy6geGCPQrA
KkxnyviPAh8fotq3olvdl7zrReCW70ieV254xitzfx2d5zZaIkJlJg0LceKBH1/a
3SgC93mKoQP2S6uR6RBMR+C40vYZnaNlKT7fKp3eGwyU22iQG/k98FJwPRUOLpYO
P0DG9GvWEjlwB8Q+yHo+lvcckUjRYtSlijzQg85HP9KXpyxEfsUvUMH5nJSL64Sh
yrHgL2B7c2bbKthaMalCWoHGjTEUzUKGXSYUutATOV7N0uoOlsijqlGGRtztKTOl
eZzC6xUOMuYB18O1sjZxNPXLcyfO289fIY6lOLnhgI5S00+WQHojqSz7Lwc0lSIU
S7cueGb1WnpWks9WaW/BZb7zyxKCWLRjUJb1nNawTl+yAk1OMkJ3spaeDUJc71VQ
peqQAfnIl+PaI2s0f/HBLpskg32/L4LlmNP9H+XL+DBnVFVFBrsrqVUw8+LefKve
VQnTXUggiX7qBImGA4nwYgvNTEAjV578W+6+Qk6rd7jwbXdCfJW1eF2hzTJY5ZXo
Jnlo8A3GZNmjFvUcZXCwRqHz2o5RAw1TaT3YtheEg9OU882YgkKv5ToENiLNw1+0
cCR2ZpFOuL5NDS1la1z4X1THlqB67bpZCWPrZ5RybwhxAHboE4QwxZWpLC65ToOG
Xy+bpp4QQMJrNecFiQeovs4ZaUI4qsklIYmyfh7MNrwZFuoCZtCeER1VD2npU6Lx
p384ZGB0a7IgMVPBvrzC/nwLuWXvZ9xoeWHtIx4FJTR+kt0Dm7rzDUjWyq6eFmEA
qNWvESYtRpRkEGlLFpA9lyVcC2H3/SRkMbqSPb5RzVmPZ6usGGkyB1qjFykDXVqU
b4qwC9XHWR/Wqokt6ERjn9ShNZ1l1wq/7EWmtVfvhRXCvkFGXkGYekit4iW/w+1T
hZqmUey0CJZGnNra0qKx+I8wPHVRhugWo5GUjW1ACvdtjETjjzaf6oh3vhwYYipe
Pr+yX7dqknybSdnidqLKbAwc4CnJ6ku+/EmBJNC7w8bo8C8doWSsTjmLKTe1CM/2
Z+mSCs8v7nQHUHtghBGeB7FFDKjIyTAS7rgcpsmyDlBsUQvc+ilAWAd+zhCZ2Ype
eldrBU+K+B3rkQQvdeeBuiZt4fhNjyiPUHlFek30xUrmeumeOjcZ+/7FDeK8ysVQ
CngoV/OL9Y4pEFoRHXGlvJmDRR3g2IzIR0hWoTGQkWJUUkPQIxGPV8OCGgYC8UGH
atDbMDCnigPZPXOrm7bFzDZgv70X8caqp3QtkAKKGwpE/4zHr27CKxUL94wT/50P
6hxlRMCzDsCFTdp9Dz8tEb3g3JRdrd/6h6sg4RLN/0uScTcFhGBZ+K7kDRJPoeWy
/RMF3wp9suQHkJvhndh1Y5haEmuwT7W7f9iF5SzESKQVXBx+3ao+AzMWqTE1TRVp
zJaQQdu7n+fU/0zptmupWi2MxbIVOoGumzd3TQLkLaGAuVEB/3eO1eIrChCU/Jx+
PbZAZfHqfvyxqNxq0roHLgyKsRoo66an/OW1rjr7Nbwkd2tveWspqjFjKiST0NbW
3AzMP3ngcxPsFOP1KWsRbCrze9KZBNrBbEAcZmU44xzqEK/QrUBUYtBM7l29Ms2t
Fuev6lcZmmiWNIpOLQQ6VXkMT6DYr6OARbtduM1u6356TSWBZsg3PHJ/Gy6zmcrF
H3ewwbIkXrOyv75elwW5mxcKJHfajzLAbn+ohlkUGKUhTuZAUfGKkrJvU3Vk5SuS
uf5hqm7nSxGwLeGQDaJs39oNHc6ayhTWV3QZnkQbEvu4MaRWrbkSFSzgu12FdCCW
K0wSngQoN/tGmZPhY2dBVUGqEqTg0ZDYiPbirUZSMzIMOjArbhKbJby+erniAyms
FH4JbzDZNsmVeHivsjDUdDoZzvcXExaoA9Ip/ELqJTmKrW1DlP5zA+dH60Z2TgZp
09Z5+tbZyREwwDV5x1N3y1Xo6tqvSLVSurErKAKo59IvluenZ6/Ykw+c2bgSLi3t
ExBz8w5hpohND5aH6vVQ3+hjqZ4dPJcH4M2FrN1rfmNFAfMBUJbIUB6KBHJ85V3G
tD3PcmNeXqoARX95cAwa0dqYvJpGxF53YIqHBy7FIVwb6YzEeatjDKqpCzGwSknT
61VNX7jNI5JD0+7JYFtkXwPr1wUYc0NZJQOjbbXLW2cZ3JC56NOhgXmiXH4zs0h+
mQLXU+Jgjsx7HL0OUDUddWwZdhPQfcjTofwhsPWCkZJR9WWfgBJw6w4m7Gpv1x9j
lIZ+jYSu5ZgSVFxJHP/yh64qgsvCMbGElyxhCF8L0EFJtbR/1A1W53DLLJucNxFG
qXcfh9gfmMoWEYw/T2h33AJ8/yi4jJT6BGzjtunKMF3YA6pM4w9RDs+9f+yEqaFE
GwJJpfBV/si/JavdLzFLLlMHH00Ft1I00M5aqiA1s2Isev4doLEEW4V0GUfGHsUZ
LVK865I7EDBhbRn+FgnXu6QTuzaMXJm4wUbhHXeHa5o4QDxn0tP2lbViTxD2hu8o
YTT64JRzNbn3oqyMKFTQqFwyQ38L13LGQcbqJiEjRBMrFw/WXQT4kQ++hXfIpTtF
eZIjj1g5Ox3LfFxUeUsKVi8lFia1GxV+NTMFHBYLCt/9jjg/BIcwy+p0UuDgbM7a
wL4G5XY1JLnKZeINqw0Jgpe5eBCYFEMKvHdHF7IfKhekvdTJSTApwRAJBrmDXFwa
5Vk4OMLKmIjsuD2e3963DGZb7mOUUvxRoPeYEzAFt/zG2PN8EWozDz0a02zFxHKq
rN2ceYoejgDe8zfsDaXQXMHfyCIJp77iOYVoSNlcpT06hQeORvO50Qzl+Y9PCx4g
jBA6zWv4/npf8ykBlPUoH3mDj2XlFdSPFzuC87VfsWY0I9x+R8Jmyj1Eam/qyud+
rOkYLz19prR8GCxh1XS6bcexLxbB/VpRnaYXVri4ap3T3X47Hoes/W9viyzyDm6T
PJax6bO5kUXPUAfnzozQfp9G2+pCRfNYo72cd6OjHq434weNztdYoCoiS/oz4mMj
Vb6X8wkTNg4z6BIs/KPpZB5EaM3C5SnaOye4X1vZXZn0DpN0JS52q6wdTzoK9KDg
3yxfGrk6/bh9LP1UpeBUXIuXqZeboUrOciYPxq0QOXYQInbZjMCU9cQ/zKIBoPJY
93vFwJQCwoBq86NAJ+hrE0PCTEoCPBpjTp37g8Ygvm60OW+LsrUtbK+a3U7FtSvO
q0qymp0KS71xochcKdyNmoPnRtCok5cXlyf+xnn5i1QG7nA7To4oSWtDpGjj015K
YqYW+ov0vQxmVF1YmQVDS6zmvib80JGKneqQbMhntBAL0SiUjEFKv/TMWYFk8r96
Vzm7i19yh/c6d34cEfuNox1SHHM36fMFVNT66xXdqrXREVaEVIUU69h/611kE4pI
+mp53w00tnRsnyNgp1EFA4nzD8t0KUTdR/EmNe5YAW9kxoAP4vL+q6nXe/zjz/ri
WJ4vG1XxBqL1yuoyfgy/dc72ZbJHYDEpocZSbz/ECX7cDFF0nAGx2TvV/PZzcVyz
r7OWlohLzwIfhgL/Aae3Vg8iM7wJ+dExea/NyheEoRE/YInZ/jqKD35nv4dDYQrO
Mz+4Q2SpQLL7QRuG26q3xK5tJ+z/C5p44dz2cL8Cykg124MS2r8hoZFwJZwZBHRH
V4kqfMpRZrxoXSWrRZvy12nKKZWM1rUCN/xl4RjfiVxFHzKaKiCYaIlXRF3N5HH8
nTv9z3klYothD0tq40jArKdd24JIpKlcEmrw6cXgdwzsf2M8QuUXcY3xeUMZNVq3
weHQxAMbhcFinWbJu/dZBKk60xFr1ZHLAHvYIiGXwROBElvUiaxPsxkHCxisyfVw
DCTAkILSqPnjQgrncrcMDI8BledIdTmaq0TaMyay6J9aT66TFYxRUtiucTVVUoLR
JpJf69WID0TB/Eo5Tp0ZGPdiyy4Mrf2fORqS1a4ASQkc9b4Wt8QDFCDsCQ79LHBJ
hv7IVWYfQxqqKC4vv/Mmc0rZ6AxdJRaFmSfFKT6xOSeG11k2F8naoU+nQy5xWvzF
UAUdR2i306yBdRdl6T8Hhb+erjrmiJq9SsI5irrmpSCePLgAbL7gULf2nViIc8Wg
OKampgJSf0aKDieOhxyHBeMTxcHlpR0x3Frp0DSfPrl+a1TfM/TYuaDQaOprUkwF
KC62KI/WjYxyD3vM8zvmI2eJvS/Y71+xLmJCZdVRP8gQCztyItOKb2rPoyExDXIt
T+skAuJ9gl9lTZVXAPTT1jY0v9d8aOo0epyLZYixB2LNeD23jY7hl6qNsOqQADxl
PWjS54y7bIDFUFu2pNq7eWrSbJ2OKQeZH3sIMf8ljYzqsjr3jClozd2fTG75S5xQ
bSZ8ltUcCx80z8JJqE3a+lvjC47TmK+yZnonJvh77sfI4PlgTV0hdlBcgXMlRdLU
mjPkk4MgRkOFbBYR5vlXaD5pabimLTUIcmKNbTcdt4juZXKaDEM86lxWGKc66u1Z
6gsiqD/FlM1ZMVinbxpb25h9uTbqbqCqDeQrUK2JILktI1N1cwNdkKY8zUrYtGm+
8QKyep+o3Su2xIFnzqZUJ9c53ghEOt2RAOSHmPFwIBG2ioqMskaFBz/44cZu4hXb
Np2mh9AAsbfu+lFHSxyA4c1KFg+ljtgKO7beX8p4JUpNtaOtQGBGXVv2Vc2ekGDd
Hk1aWVvzryOuChKWwdh2U6ZQDIaMYQaQziqYV8WqOgQrW6eRqUQlEVc3RiA5stqC
sNXbbNOtZfSZU5Gc+qUdlgOqOuya+flzqz7mNsRauIGYpHratpyzhEP2Itq83ZsZ
vpDJ/ldTgRJQuR87girCXiYmrHp2nCT3D5iEzaVo0fU+lyKym26nxFxDuYMXKo2g
fXZLSiCNxkWPpNMbX+bGS+DNs6dhpHH2dWJFNtoz0mqJLOHghZuQP41x3qX3FSDm
xYufukce7Wc03x8xuMbZJmeZnvzeV/Er5oj2jxt5KXI6mc6ndoz4ThRHwWBsP/vL
qN7G+Io9q3MbXnjydDedgcciMHx7wUcP/trGOJFdJnO2OB3IUq/T3kXTha+VHfMv
sTmo7l3bkFMTojBUqQ2z+uGHdYrI6KEmslwdy/nc5s/AhNudcx4zVeUu85Hn0780
s2i2cxvlAXm044GDECUYBpYKy+a0EK4Gtm2Ij7QYdpuNr2JngN/eDItGm/XAdamO
ggtEBglsBXtO2amV8zSLsjlB3kzxX0/eziW+/mEDHvjYKFR7tPhdzgFWegv0XeK4
XQmqH+WijRDARiwKUn1EDv7DU59zBNv4E9BI78H5UcjZpytn/ST0ltvA/pOqDbaj
zEjSR2fwWCwckUfZjkFCPi0WxwmwX9DyZjVoneg37gXVwpPm18+rVzi1fb1dMn+4
KtLozeQaOBXtUmPYdy8NJ3QG5vTGiN59BPqjX2KD5xicGziWDVd2ejpR1NdAHkt7
z2QFilc6v1UNeny49jYE2QycELblOuzQMQgitjFrGYyS/bdYZqzsqeoRvJknRPbw
h4WfMwBunkCQZhlxFbvSEwz+jvpZDQC/u84LSZDBIZQ2qVp0uzgQZdapzCssuE7d
VObmkXt0tHPxABe32io2Aw4hiFrNwiRKyxFb91HqDXSdj5BhTK5PRQPwhnzYtJzs
8WWBve1QchM1iHoAWLV85qGq8JnSVPBjnpy3h0zOrJ7M/Ang32xRjsb0TX4uiAQS
tn3/JcYRkwEwCcMZVIhZ7EbvlDgkc4DsX38c45pt4PF+4xcZuQp8cHpZ/3eailb7
FXgGVfoxChEcPM3jhQc49NQjhyMJRDDdTux+J/aDX9Mh8DqKekqkT72cNL5y9ZGW
MV3ZlVPH9u2oGfMzrpXMnHFDU7n3UjBKhCjjM1BCQp3q0r58CGL1xy29h+wuUIvH
59Gz9C5qS1uHcWSIlNT70YQyLTTK+VK6Vq7cWB3j3ilEDaujY0Y9Hc0NmGkl0rYe
HO10o7qdSD9h8kzBebtnKhiEQzcYRdPFLcBqB7DfSHtLYlx3UI8/ZiPpSAM0arav
UBuU9WidVaQyI8TdxIgSJR9F9b/SmweQjPmdLszwxhCYy1kLKwYKBJdUZ2ccKP82
B1+S7wKvv/iDrtHrxEhxztVD11k2SaoLUvHNvFYxnFSgqqVpAUjhB60ytCzKZJA+
ol6Xnj0zvhgJzKFzjU0BiWUhVFr8KACp/b+b3mlmo0D5/9q00Pga1BWOpbIx830I
3ObFVMl8N0slU1P2BZ7l1+N8bEd54dP3x8Rr9Rytxx5t7u407rLGFBT820BBfaG9
FIDLSbZaLOjVDLjwiwHFhGO9AdwUzXNo7bJjgjHUpLvHvPoZQ9QPPLBJp8GsDVsi
uGoCzE6yydA/VHdg7WXlStJV3wogpJ1uNMLYMlajvvaJ0jxden3KqRU0bH5/Cpf5
EKXs3HmvGkU+CaocX+2eypDxnuCP8VxJDwSlqks+SlMM4YS9iAsmWTHXJ7+NZ2Lj
BG8RDOayeYK6kauH2uWoYTvKx1UL+zThc+RuQQvOKCf3sPQkr7vCTN1HFte1Kwki
QUKJxwMYYr9LOgdINZsoAhkIhzoEbPo8Jb2WCP6gHCVbUYDTSduugukiRbYlNIhd
MS7fceU1oqTWy9Vw4PuOy51AaYSAVf9wcLdaHCMVUMQqd9ozxb2SZgNUl8iPXV1o
CquPo8kKtTNV7YmYXkEkkDmPJqWiQa8bzLnutEMGnZ3hwCjpoLo1z4jADp5qi3Bu
vqc/nvAym128xw2sYEKwyx5fy0/qx0EWT+cFTnN8hi8uKcIYQsr56Qcfz6co+yQF
JvFxQ0Duo414dxHNwSVYd/gpwGdt+d5PxebU/u9jC3oC6r/kLviuPz1TbmuWeeS0
0fdQ/s68nDatdGmCGz31gpPxQ5+MHXlvTYAYInheBKwUfrDrCC2qqoYGGrJ4QOdS
jD6gF7A9DqnR9UV4Kxe2UVt5I6hwPV9Z1o+0HAhgPfLDOE0t0p9wf42ef0swdTf6
+k5QAoNuaOoXbnrbIGiAjX+HqX5bxvEIsTAF3Dc7wyQifrhHuGyxMV8bN+uCfE1S
VV0wC9ib3y7aPtQCzSVvEvVroWrLiH4jdBRUEix2kI2x7TofdEwXKa4VKs8nYAJR
+Wx/pZjbnScx5L8W/Q2oeVf2BGKL/lARv34YYv4iZDrEXlcKdSjZIO1cWjU8+9bB
c4dRuK11WSxrjp3+igXH39fe1DvOYFejskR7eGCapViz3BsZ75GOsFkUjfr93RWm
uH1xLERF0kJ+2qXockGUItEVHMizNZtHWgLbfEppVBfSGldP2YyxcrCrq82E0ENV
4nCstKsfo41pY2Kah17KqQHloqBdU5KQ0efk+aoxfTeZVi7vYyJH39IXh1AQPyiB
DFbCncH1ke8eWmTJlTht3dYE18hHvS4TGiX0/sH7ophDjg+LY3noZ+1P/9wyEFnH
6CYFje9QT4M6swFRO/VYwU98w8zvEbrhZyw3M3rlM7PXp1DCyyf+SkBj1uJWQq7d
Hp/33cPhmGyydvjMVm3GVIed1VS3SXek2YM5K5hIjBedgtoKnHCdCJl+wAh5hSdj
3D9qdfm5+0JIIcUzXOTEeDGFw+QbmCUbJRwIebVp6yIDkHTGU9qrp59ZSZJke4RA
47A+BJu0s8G3QKV5PNvd7+ZIbpJu9n3+Hax3l9gmJbqFnl7OqYZxwhRTTMUK6osq
i5d7kZ9rvlx3PzjbQus7sCbb7DXKeINOgXvdfZUHln5cQ4tnpHJ150i3OTfpZfS+
iTHCYcsvvGsZAjwivbZYkcLMWp8rAaCBKIyodQxcDZHUrJGMIUaMAG53EOmSKMlV
rnomcpPzmD9nEtbwjmXSsUNvs5hCC2P31rAmrwO2J0chBC+5IZvX8ycHG3O5FKHm
VOxW6QXoTXJeG7SyW7OxX+3jZ5M1g693UNpCOIucCVdVoWkHiWiCD9Jn/OcbMBv3
leEuoIU9Pm5hsLixvgWYRRT0x5oxVm/7zr+paBzVC8Xokm3ajOgY0ERBPSnPHzzl
xCCGj8kr6Pmb+2wjSEI6vdX2KYLycUI4EtdQqb2SAWLmNCh3d003Z0u6tbcXEmvN
itAzS5mFIa50UOC6Jy7hTrWYEemJd9vBdz0MfAfa1dsd2wJrSEwvDHu23oFfiGbZ
FxuK/jhNuZOfVMTM2Fpa+0mNjE3QQkNRJFfpC1qrorPABtpChAI3o54QexCQq6Ut
s9y4O3mw42ujY7aBjDzYMM7r7l26OLKG4Hw6qjGeyD+ODNe7WPRX7/8OpoglzMsb
7YFJn0Y4hoBqA1QnJ2Rhjd3XARb2EsBCwIgEPUMw0UMKE6q4zHv8Pdzttq4vjqHL
d8Pi9c2PVuhaSDjPu7jJjp5feoRZFSAeSW8wdrfM7gAKt41VNPhuR6fzNapIWkSz
ekL7CWuu4fFowyFR4J+H6pqcyxI07SsciNQPbUwl8HIMz1qKSwXcrunxKmZnkg/C
/4qD+rm9vDz7IvF8tOouEjeAVaB0Pbobl3jQUCJPNXV4ycUMjnv4EiUS9LNiOmH7
6GGoYVrGxplx8z9DpoNEO3kylqBS6rSwlMewdlD8nBM1rMgljcgknBKVPDeA0fla
EwxUbd6+Ev/qiPO1iu75YZ8t32aD6o6cq5kToRuUKRYoMnY6J87TSmSkMC+EZYCC
HbuYU6ff93w+A5wnTz6/Ak+Q0+7Ld7IpozLQWlYQ2Amu6/5DpV06k9ugDeGrQix5
Ik0aIUMNvsLH0IBElbAxe0AX2ERPIB4fRTMW3MOhwMmqNuZ3GibQBvBXZTls1b3o
MwbcsdzJK2bUhoXCtIytg7eykZzSk/4S7jtPEq4ewcPsvO4c4lOw/oNRtUWcpMHK
+dLJ3gYKdhU4eMT69YzGxM02rW3Tz+ouzBorTBAnTKHApZqI9WjS5/NJfLQ86LIr
Lh1+a+/F2mGgoqXVSpnAIioSnMsiSDYpKqmWHPImevydiyfK7FxMEUfav2SPNSAy
h0JzrYuUjwwsffStjSKPz1R5C/2MJpW8IFu5MXpx33e+WuqXBwprgsSq4aL/sdAP
67248NM0yZDdCbLR6i77/if8W1wP72m9TjKzPYKWS6SANve+/MeBvX4OKP9NhINx
YLgDkwf4a6cqhui5Ax9/GdEnLGU0SvCDe578pkoLFWhpwxe/uXxo6fOaUKftCwDf
Ook1KhulQD6clWvOCYI6YEGxhV0CSadC2+Wuerdxev1YjM9Ye2R78u3yZ2Nmjkaq
ApXKDB2+iSJwMTu88z5Y8tVdwVcyWKp8mecvdZUTQ+E5cUoj0L0tyivVuzwFMWDq
0nUScv9Uc1nZ2wL3unUElaBbEYYfJ0d+MpeOVo9Ym6PUa8tfwTmjJV3Shs+qFRul
+FakQNIT8WjKKPXvR90Lq12Wk4gaU1g+Al5PZJk7020c5J5rTRFpnaUJSbRIQ6jZ
S4LZ9KJJzCxPIOiH7bZj6xFCm39g4zuZv022b/yT2h/KTHn6Z8nTuptCwuY+zaWW
ODAepIwYoTSxJ9rAyKEyoRFI84anF+/t3R/SuugpDVpdu4qzlkMZPz9YjSmXhAdM
9U+JLJ2Y4r7SWi3UN7U1bzgMQM05z+KSUlznZ1GGPho7zruTwgZUumlPNGn2ec0x
+OPWPGXDAtuO/sbG5ad5arnP1jtB2oyEAoRNSlGkTm66yxiIOQ0pN29gsCKBcdpj
7uz38bUuuHz7grvpEUbKVtWKoAcQ53J6GJWEtquthO1nzOaanbTktxdlFZuvdBhx
UhNCBqo2zNA+yF3kqFRp/HGCn9EclqFQ4ZzYnuSJsrAOAga8M32WEt16O0RWaQsd
7XJADpBN1AroO+6V7bAetpW7XRfIoopW+Ucq0L39DWGEBVonMRZOkSkl5aj0G8TB
/7UYypQzVkUq5mzZyBdD/O5M02c3IeH5gjWD+0MXx2veN/irZvYQUFt1UTc58t+d
HEh8RO11o89Ih0UnceYWX+F824pB13U1eSgsTPgezBDDH4/OFw24/qiy1gQzc1o0
cdx/ueS/VdHL8E2NUB7cqnD5Es0mgKU6V72pvFm/kqLOQ57SlTW6+3P7dPWZQ7uT
FQcOAjaH5YsJNucjGtVLDShvjedvu88EHN1n3AN5GX+QHjSb12CTckRZpvwdyVJa
7VOsA8Fg+NtPVHq7PEmbWADV0YtlKxZkhy9qvLHqYZD9arviYFxYJDEE/tY7F5Un
NVKKwAYdeIY/thZ98402XWQCEGdxIorW9bO5JLf6+v/rn4jQn9rp5djaDSnhQM7M
8csPaUVXXHV8OVqt+oGtGQiGWfiqOU72pjNh9wavWADXdmHjFB9dGO3nyOhZIySu
Msrv0jftPL41umzzO++kKrv+ebwk7frwCeF+BNLPRNPT7/nXicK6JSZiU7yyQ/3e
pXdxM4hl4o15s9hrM99HCiRy79lVRUj9aRrpV8JdHo+8le3rVX7gRyoxYCARjKPz
qYhP5IqxVOh2SteO+cZ8TSSphVB540/o4aZzQG12oCmEhp8UT7jZRyee3MbOaWgm
bYoTqGFnZLohY4mlRDpSXB4qBqIGKFGndWWp6xDjMo0HkNO+9CoUlCUgqyV8z5Q0
r4nnF0Cb3cd6wpl4GV/ajBSgz19gq5lz+AqiV60ffEtDyX+uze4fhRzop0NaMfYo
y7SpAIdLrtzgm0GmUz8PbRbdMZVOmrDcC31oCsJMO7ToKN8DufJOUIBuqROxUSuv
q6vN1nZYiMf/8MbAUUpTeneypkw1G8dAmrKBpDXLRMA999qa7umTGNMBRzkbT5hC
G38kgK0xZl+t7OfLk+/9hIcOuwZYwcBWAccREOpNu5AHDiyp3aHODDal7viM8CbK
7eHuPNE4Bah6TkXwGO0f3Db3Blkco3rM3xHcll8bS+fveuVazxpvjNQlYFzff0Qn
+3ncMQZWpCz+pNXOpwvpXwyrJ7fzoh69k4YvthkQZ8Qttc4pLk/llQt+rjRiW5Q4
QHUfj+qZMCXWaFsjJng/3SKLr54IysqMkAcdgMyrM3TpFcY4FSV+FC67O57rJMW5
no5drN4wgmksL/wbKAmQYrIWrY1yjiO+ZPSqOQwkubUp/1KwBtN50AQs94QBqWJm
jNQeHPLRKhyMBomwHLYWgAT/8/4WJ5FE2ZqMPSIKMa4s/T6mG/j1z7HSYFuyGQgz
aLv+m9gqSlIEuqAVUaCi8sy8Q8P/Te2ZKMP7Gk+jEPeds8xLlHPvzeiCnv/Mjo9q
4/7dOreqgdZbTBLyp2hdbesIZhblxKSalLtXhBujiRFrNp2zey0j1ENjkAAVUbvZ
VCbi1FMM7uS7EvbEWgl9XHolGlyXfkuhhfOrigFyloUT/WqZIaM0joJBE8HAYCBv
/H6yeTelQiB6diWeQniJYC9ynVtgoI+Zbo22UlX707fE0n5uXU8lTDnxy/faey37
y1zWD8LTmiVug5Qi6NeorSDm82GBTR2zYnbx2+R0e94=
`protect END_PROTECTED
