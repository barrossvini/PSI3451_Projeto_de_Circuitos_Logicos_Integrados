`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oipbT0c1ZK9OmiRHYVBC3PNMZimUyfGo9rKRdJUUZjn5i3PcNEg8PaGx+hNHMMK0
5InTzqJMOS18F8YGvlMZzF0PjUkUX0SpP3gYy+t3ezwuLtVPecABqawMOiicdPNC
ZtbIKKQ4dwSx09kYDORaOpybOzActTxCOc80W8wHlmYtj65b3GNPDGD7RiNfni8H
hWhyNrOBvbWN/qNzX8djDSykqbjVEtHcPMRt2eSmo3D+UxtHydNTqUP0U223ZN+e
yzr6MvOpbTkQfkwArVHQCI109ZgmAJtj7CYtHOh2qVBbLSNEnNmk5Na+/QyVFq2n
uD4eLj4BRY5wuwja39LQDl0qPtKMZdBG/xon93u7m/KwUe/7S3Xsw7JQkAm+UXcu
4O3NBe/A82sJrFJHtwRYhqLQ2bhQ6pVE+NjIYhcam2F/Y7lQnaJNxJLfno6no+Ge
8W3pjPs03EHZ6gydwgLrGnaIBMcD75uddStzBxeToPoeBvSV10sZo8xUJ5AkOXXz
UlNBxMM/u4SHpdEdmbSZtS0q0p/H5lYF3yxSDY6UKIIiOUpW3Vu4SFvSMSacc6cD
RfD5Uwm0Wz0rNxGoS4t5eeaVlVAcENP80seVWb7tN9XUiY8yLnnn/jPI9rwvWMOl
`protect END_PROTECTED
