`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9O/ktf5r0KnAMSNDUCO1eGWdWQuSvI59HIpVnVT1yoWrFwGFobWy6nnlhIcA35Io
JiD7U5LljIpMWhG5BlmRE7UBCNyNNjdp4tE8xR+LbSRZjrr3miCeU31lL8/e6vbK
DWohx7G/90SdN2xR/KeeyD7sUzjgBZy9rBUD9f0narv86ZVZWMF2//Er/G5XT1i0
gJHDvAEKsGIn1E5vN+jTdidxI6JYejH1eu8L+0WJc1gi2mm5ldlkWFRMdlNJjsX6
fC44SbuBuuqV3c9FKJqon6+xjEUtTjbhuN2Y0W6mKKBg1uV85eHK8RuEMRFuT4bA
YbSeOZh+zTyptVtpq0WklZKMbdy+GlxwfkDlX6nm+MI2j9GmM5w0qLd/jhDPBq8F
o6jA+JKlXC2Ltz6hRXN7+ddrAgUyHoI+8ceDu5bz9s+1igL24+Aw+90sZ7WOmLDV
Lyg+xTjD5uTpG2y3P5FbZ6vwoFez/3YYpJdRy1hb8+TTO/HRsMn0SdVCHP5cMnYu
mIqweTMcLHEMEmygJT+n3Q==
`protect END_PROTECTED
