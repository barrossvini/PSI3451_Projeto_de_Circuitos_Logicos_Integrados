`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C6ycaERcdXSf9sGVaIrnB/6Ji/Ik1F5dvMM+zSvpWJ5NxVy/dAUiyxMXKdBsfisY
iMV97U8lO+4HufqLKG0KMY92b/JRJOI8Cc8sZ+ONKJB+y9fqhA804Cc46T7ALSer
9DHiX6Sbc2IPwi9GWFLHZJ+DKGpuKmma5TewCCtrmGn78ACTkvRoQeA9tArt75TY
zBsdtK343dKGoSTbV4plLIf2ZQgjYHgrTHh5JgEEhaQ8AnovWlg9LXC4tILNM2pP
koed7NM1Ew42btCZVi3e5oXeisz9kn9/tglfsYxeweeQ7sFpiaWWGl0hwaoQd6or
FPQWi4xKSOK5hbe1D+gMTkZpxhyeFiRXLpNpzgKNwaNPSacKBWV/bUpVsxu8bRCV
KfDQ20CzpyheQAAVFMFsL31ci2q0WgRnXoi8oj9BPDH/ykOSTJsyWIBQ/SqyZQAW
LaBnfC/pBrtg0iUObWPIidhvvbaX+L0m8T/cy6DbZjxwtIqKSeRl4tY62QX1CNWt
lqNLoU2OiDNUd6ALMF6rfhWcZ6AYbMk1hFYrCdBKJTqGNN+gWLDZX/gnA3lyPuaK
IUcB0fkM+50M5i2EcvKyXB7rrPjR7aMbyxW9Fr8AuaU+Nzj4vaIDb97k6CETFd2y
taP/fwfC72J32IM0V1gA0XrCsVDMlmkMehWFVWZxWUJBQw/N6jWqTsYxQWlpg8KO
c0Bldpus52aWVDwQwPjKK7A4Qppw4S0u5NTRxc/ar/Gl+BeTp9CI4K+oTUfP7AIl
SgC1hmyHP3vUCOLN8aLbqtnZ9YQGuHvSzNK2ifg4z9geTMPiPPu2t8QAyY+F25RY
aFRUthdDl4PZOxcmD5IrvtvHqVe3+DNyl3bvDUvQql5ytFFcPzjFJHySZRf9OHwl
+0LBPP52lzWW5UeMTHXmIm6EfUsUsAUiXbjTQ4X7eGpkHxFqqehJXtnlhiZL12f+
d99h8iDuJqIDjh/yHvQokMBZ4opWqX/2aTEGJGvTfrWId3OlC3hKi9Mv2W4LB+pw
OoX9Grrlx3nBTRhkjN3EeM6D3T/B7yGopKfExGR9MKaqgnYEkAxuFnM8Vz8zTnKN
F114mu0ZnD7XKqKtz0oN008Oz+cxygyuQ7hhIgFP4Eg=
`protect END_PROTECTED
