`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qW/ldRpTJNt1oqIMjpH0WwtozYhGv17WI0Oisv/iYFK9cXlFLXUJLQg4LNKdTPRk
fi7sPWTck0LaWsM7RnDh/2nCHgCtY3AEjXRQsOXa3fauug8BveZ2Z0Q4IB/CyQ/C
fSpIioz0dB0JeRtVbKGXHfolZ0E/dksHvXFazj3J9RJQjSkE8q8LfEhIkMQvjQYP
3CMfdN0PtT2RRP0u13UvrzI7VThov5WpaquMvh2BBmKFb8skxXlkxx9Mw7bDmvXM
q2vyVMhL6dWjOVBfXvR5KiQaqbQy2NFw8J1eqK7qT2/rbEilfN1LEkl5RGAg9m1A
SAHHPwiCL278QOUuNEN/NeVmPtGx/qqn9SbK+E6iAkNi0BLzLuCl9Td6dRtnPeb8
0HhfQVaP842v13Emuj3ZAlxh09v9PIJt7w0iA706Y2avka722B0qpuzDzHAikGvy
/QfVsvxbbSRU3PTBoRrMG62OE5NpOzYBS95Au/4xjmeFIM3YyIHsI/dF3vyFagcz
R1HWhOMK0wy6ZC4GVhIKVtOvlh5yQ2qW9p8hS0E7nj253gQjy/VM2vo0ynl7x6eH
bnEo72MG2sv/iycHmGJyCZ+dQK+dTqJg/FmwsXN9n/P35sI9A5xjbT1DDjhHOAjO
PiqmBFxCT+zLY1iOJQeElT9oK5vUm5xjF54Y3NTSfIoKYCBSOslfDeiCGTP12kux
vzKNdnF4rcT1/pLb/9ADRpBgwzV+ozhLO1q2o8NluUxb9+zlz9jo4n28Q8LFFCf3
/TYUiL9QxwBZh1KzNQR8VyH3Ug0gjs18x+l4cwckqko58geyjVEKTFJoLWrsk02Q
VQAdcmec7VtN6gZIiYdVD+raIjL1Y/5c5aFfpi/MoEGirOQINMNEJrUJomG1TyhK
3HLnkXUgDHOLKX72+ZZSXKqgq4CnBpnPnWw8jTOrldQ9g22L1dJacljnVRfc5hkM
eYEgJnKCBgTRnJa1dDKLrjDXrBiFa3/5JXpx/p7yyZLpVxO+vUid2l3qb7PaNRgi
eB8a6UsYzb/B0lxEBXHQNds3FMolsWK3spCnte6HUgZw5yUiw2KjQL2RGjWeh5tH
eVdtRh8Wq+9zaHBu/G/eQBRVl0stfyYfVb+8FqYovTyU+gR0CyR4kfkU+uSG2fWn
A5ade/Ws9VqY1Xs8CCkPWyPsO7uGGjDlWK4GvgR3U5r6botU3zHmTbdAKUzjzIwn
4TisJyOqw5lCKO6XVHYlrrlWk9X1TDMiVUAYWpXvAWVx9LO2a2iVwUnJjDQIcj+S
0vJd96mKg8kyBmnKUMMOATI+fjCs2zFagEkFEytkIQSaEPdeMManOu2mYUSLlAH9
K4iihaPk2UQ9RsIN+IJnugbnzW0BPl8t6UYUybhCeiD8wuzzpIi2d+lWc9DB8OLw
d9yZ/U1OpGtMX0lBdD/X1wZNIEG+l+godhrv5Uqjy86RtTrQN32QbbHRd0Q/7NDY
O3Kv/U+jpuJbuZLWwndS5mTZbgQKbxZfBFLJAkxL5rQFBGies1LfdYtmNsHZQ0Om
6YgpvTSo7cwW7bAMeoZT0RDL/Oxd+lsazm8oXh3aifVLCnGUGucP2J5RuDFLOJVS
lJ3mInkLDKB60RtnoIzgDzS3A0xsaM82V49YxjryDgYB0Zkn9etViXWXQ0sh5MNo
rBr0ATuGnzA3TuYdVzqEyaKXg+5kysKZvS47Svea7gzHFj/r/k/EouyWEn3N+CgU
PJ/P6KVs5/sE6wxSV0rXUVFhCWG6jos7ERibGjQAH58WNRWir0LN+WoTYV0C/1Wa
inszjlPH1ksnlfxnULlmHuc5qrxBLUymoKo+zu71j8Fg1PXLeLLtLT1ECFo86lBV
O5Dk+oM5DyDpaLOiWIgzPgehNHfad4PVHR8KDG/BHJeQTK3PCdFSIvuQVU9dk6Gf
IZdqc+2Jip0j3khHR1F49wysx6E9/aF6sz8dEaz13uc26tpuuR0HEsAgzK6nSkHt
Da5sFz1atps7ZjKvptZxm01OaDIoW4RA5ccaLWih5JWHE+4cTTkbuRCf2mUm/cpR
6YInYyBAd4hL9PaZbCFuIc6k+5vjbRX+NqDzkG9yYK2T+3e/Vfl0ENvSKdE88PxW
uLZqLYvsh1aJZO1hGBM9al7MdziMHSCWi7G+btW1jVj38V4IA2dRv7ar9OF+Jgql
KoJqsFiDA3YcsIcgbzQI0ot2yws1Nn17TzwN0QL1rw5Tq4fIQK5mG1rASdAGPR8Z
xeYoJeosgpla87otBNmssNdfmZOVgve8B61kBTcpDY/hzijJSpeHLm3rw8nn2cIB
HZ2A2gJ1dVfKH1YKPc5ZDWyblLVagTmVBZgCsosEo2bW4tO+DHjjci1BPXc9ox0h
Mv/oBJgT9F/vZElVymA/nG1htpIj3vPiH/+LZnk7XpvntECVVm+dD9nDjlFXYHoK
TmAoqR9kxwkOPcvSxToGzQ4myNflC3pImNWNc/S9cjH7nc8tcPXlq1LV1lPAmk2D
g3boFIlxosBxCUN7rNKNWTOfAyGDSjz4xEP3SAbx7dzcWsqg4t08HfSqCxLo3p9/
PPxMXRs5XXTD72pPfKPsQM+nO9Llj9E7YASdCnHKAMce21Lh5fX3bgN+DEpND2zu
lJ0y2V4oWatO5TQGeKbS6tV3TlYuTHZjnWbXod/+OUr/raZaPVaTXOq0pDbxbZVs
lmeU+QxDaKFKGxrGszdx21vqA5oqXLTH55BJWf3mT4u3EXEEL7Atc+MUHdB/afeO
0FHHxx3eTyCoYnfaBRpyqnRk/Jbobj4GKagNbzo/HI+tlUV6bU1AjGD+iBBtvZkA
ulZC96KAzhvu3IWdQOdoZiZJFfUff2+5KmQrE+gzP03XLo5RQb242IYwS9NR0soK
bIRxroBajSLACCWfBNfFV+nEEQvQQEXhR46ycfmM+Xi7LxZti1TymZhe0L54uzkh
OB96UuZUxBwy2IGjXvpqT//XvcQn6T/Z6fdR8PgWr84CSuwEcvyakebnezz+Cthc
ndn7orbyIBQYWDj10dvXvGilQ67OZD+a0GSWfWMJKu+BRgO7ZmzxnU6b0LDDveBt
3XIeBroZD9rSfMXmX63/O1gyGW3weY9wRv9mzVFqyxQZrU8J+P5FyJHgcGxUEx2F
LWupIi9Aoen1mkqIhapyC9rTQgbgl6X+3HVFNZUkeB4tHkZXJvV0On6y0TJYXMW7
60vj7x0+9SfW3QzOghcUDbQningrTPVZu638RKc7ncDHzm5STdWq4CCbLyauTfYi
UP9IMnwib5qV13kTMLNT0BgVvSZRH6b9MBgBJreiJsZNRVd2eiiiv5xqJoSRHy2W
U6iud/0b0nZrfFkz21qXY6wNWPyzzLnXx7KEc/prm/yPUsi85FEvuSrw1qnpbaT3
+Hd0F2eRVWSx22H1TXI/yFHe5qLJ1WwvrIkcCTpctWaMoA0MsQactP21zP1BFD3Y
xZZcjaCV+ZaJv7A+JsrHgA==
`protect END_PROTECTED
