`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tc4Qa1yxLwORGhrAcMMRG6yZZaYnGSEwp/rTSJmpojHmXTM/T2MExJu6BcJuOa1W
k/Q1UVJcr0q8f1vAHL4E/x1Pa5K/uB8QkjqZTzcrYDSqEOXPLwvR83CqmaGWWC7B
p4swXyEpHD4H5GAkrbq+UBXb5Tc/fN0fGgPzVIYhTRrh6orurebaZLYx6tQlrM2J
u+UPaYuFkoVxsv2IkLwl7lWJmsswJsq+gBlcTi8Xp/AcvMB0B1xcUQxLPjEXmPy7
CyDKwSO8jdWBIqRe9ypQUJYvmKUiD78TBCunizhDp51s22C4TsKvu41ayN7iuYO8
z96uVURNKFqGm+25XhDx+ylAm9N5i4GSnh9tdY0uPqOd4SkaoQY39lPa5vd0lkR1
c9NnsZvT+tscgybv6IRPgye/Mc1gmbCtClTExUNW64Rcj6WtP2osiJn0WfX+jrLI
bmq98oCAtCgrxpsV3Fr1twWdY3vLTjsEX7h8WbUhMZ4Yhx1s2uWVNuJGZsPCHk2R
cg3HYdBcpNuLU7tLU/XE1OxPjIBL6jh+MA3R8abvVJk+XXpo+b58C0HZxG/uZjzF
Ny/4auICPKZSPwmnwf+11wCuQ8jb2ALLAwldf8pdj4swSSWOY2e8Rlnu6t0kp6LA
G3GybzsEoW5EPASjegQGC0WFApMUXz+FEdrj0YmvR6mfemIsNReVSx2NgI+hf9Hs
qaYJeG7WG7b9z7uZbA8BePyLc58dHez+juSdZOfeWTlBqAgPtzYXqLIevNA0JvQQ
6C5wBZGKcCK7N01/lwHxO9EhULhNPuuKmmOEmlhJ3BGBDGlYuMP/Y1BG2AOFMbV0
34ncn/3LVXCeus0jJz8GlVgZAUvO8IOjU+PyDy6NP7S7/MQ4wKIygXmrf0I1MJ+v
ZZnO6VVprfTSTAx3kWsZ3YLz+5M78CVRVMj+gaG2fsBYJikXqydNN2kwbs5v1Kma
1Z8Rc7bBU71fw5ixtCRhe5XxmjSwrhESMJeH54iCozvUhR2PV+WUxl8TeBvCtbq+
Sp1XGMgYgKRywUTPbQoDKeXp7fjzIon+NVa/MkEXiMniKNYk3Wy6nYXGdWuS/Yl7
cehTdhhhUhVFItcAYZV/d8dX35os71aEfU5nsrlhZDufQQWTZiTUEW1j1p780d4R
ZrsvZ+yD16dAliG+948GFVCXgiJxOo1QRhR0/jZxF4g5bLcNuRuEm3IiBIJByL1m
h6D2pM+FJbWwyWk/1Pc1jA==
`protect END_PROTECTED
