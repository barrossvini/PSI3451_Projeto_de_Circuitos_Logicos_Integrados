`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ElcPgFpm5u1xUVyjnidI+0LlpubshKlilk4/OBczxZ+gM8xVedHF4Q3IqJZjFlgR
aFFb4/rXJD2BOA0hcZBcQzKSo8+mZc2dN9NX3VEmflrHYmvJbzmLTJ4foZbUbf7i
a9cxlYc8dsKEwWvQBe4GZN24+vr6OzFpPj6UfbNyJk01FzXNFvavfl7QLUJ63Oid
0MT7RiFfwcmlPfMQ8czmrtTTxBQfWInAllK0alcUOm+YLb4Nw2oQkjp5T4FfX7MM
wkW4zquLofcXncLhosszR7GUsmUAx+ThRChPN/UTGLptct7s5HiGsTO54Cv7EwFB
eV5BzQDRvk7ZtyE8GSfZuFk5wXXqm7YQN5G6UZZ+VkcG2rOURX3SvnZGbB2tFqZ0
/8yu415dIKkfy8zIP6lmM0T7JQhmsLX1CQtpLb3bE6vFenjITzq94F0ZiXhuQadf
7cvTXFMytA/9LSPwR07B+RoMYYQbSQjFLDXI5S0pbVb/VRvKgYuVdR3feTNW5LtT
yAv5S7xy4fXRmGO+UIGi2zVAPdp2Sd9y1yHcJEpn4XL+gEQsp81cS5kTdJFQbU+j
oS8SIzdGxIRjUs16OjUWBXhXVgfD/0oKoQ/g/tkuLeFBzRzCjneDiCu11JvAEH5H
dq8MaznutUD+f9bg5/MjhNbeRHKbc5PU6FA281T5VDmFh7BOKdDSmtCVEjve54Gs
z9fzpn1AjSVzKV1+rqMwY0pl5yFPdEPBi7WHNNPFpDVx3KPhUgb/hZFfJKma12IZ
zE5rfhCcJF8ZfOmUfvm0ty8QolNO07t8WaNu5NI9yzngpKgiWyAhdjGPJFtJ3jCC
aGMDPvCaiLemweRYys1cOi5gAw8txs9ia3duWIMg+NMDRCzOCoG79YbQvGHUR3WP
7HHHZEfhNtbkic6sUfosoulK4cfbUEPNPeJLzjlayKfoq7On+ijx7SCGrDGIFfpx
kneq36zJ4tpLZfEO7u7HttGy9olUKr32Oe8/CMmcKpfREQcQvyp5p+YF2weaTgJT
tgiL8wwRsqcHKLV4ZJFXxsF4qP0SQX7xc9nkT3Cy7hlF9EUh5HEu3YGLhNCmWDoE
eKeE9SU7oYM+degjVeDz5eCUzbKQWn8AEoHo8qTqCDe+8H1LtFYXugT9iA7QMaJA
C4D/gLLRo5ocuP6wqU/g9TKagJd4YkNatr/TtLwU+OQZWA9vMrlt8KlCknC957ir
7mwF4mRAfTRfg3+k4OOa3y7QiSrMeVjY0y51vpBQ7vOKLrl5+KjGyMHstWlCwiqZ
yuH9slS4YKXtKV/Rs9RfUIJ5XqEnbDvt6XWFCMslL8yNGEHltfPA6P305ELikn7r
ndV926ZpikgvbWRsYdquhZi7LvgT6/jRhrmiICT3yVpJT1AHNFNc0LqAYpl6RahB
qf+1fNMMJKt3PK98tIEQK/Xk2eZGYGJFxy2zGiuTggIiwig3nIKOltNUM14GwAGV
xn9rw89leJco9HDJRzeNB58WOCNdzhZlWyDPnLMntPqzyxdtOIyskbVBINK1XXzX
tKDiHdgm7f75lkR9g0nG+Oi7dx77Q4WkcvhtVk52k/fPoZtC7VW8OsIf7hB6EYRe
sI2FIjwj53pI8k5IdtnaeHrWWyh5NUSMpTGR4Wn5UeUBJ9lEf3kQLzokGs4eXjKE
4baF02kXznwhgjLwi4NkzEfoPjGcJArN7EmaECdCpz/0WYaKOQ0t4tzilft5Uufc
gDJnSl494Dpvn852Bc4Kx3fAVlIZTRSa6kwFgQiVyGM+DVOmiwLSGmXKhbzU+vSA
aXmST0+UqeAuUhnrYWTHe17W0oTrJ9tgaTFKr4egtiXHe2JavL80/p2aEy9SmLa9
GYzkL5ZjvUzUyMIk+iBvE4niYg3Tl16QCvhA8l4g+N60RzwmRt9xzmpGggTvs/Ck
BSloTN92YBmoOUwvn72SIWWtOcu2Ux27ZDrk+2FzGVGNsBDF+1Ug8PrV3o4PMCHA
QxYSoRKF9KYojWxKtpcZE0U2tRkK99iIXDmh5HcmX+ehwVWydJTaNoEfVk1rtZn0
LMpACl2O6XC/iLSodvyQdip5Wz8FftysOUUoZl5eoK1UkDMqhUPz/CJ1FkDbIUCk
mHz9jsXh29QI62aHkIWbU2WbFZwJ4Ng1n5f4+D0dbPzbnBW4lbuc6In78LcX3hlt
dc2ImiZ/LeMP+W82+w34KSVEpha4O/5pmfioOAHnhJiJDfgC8W6VS0vJGGc/LM6V
2G8eP1d1yJv1FNN6w5wrLpdd/1NcW07YahVS3d7Sn+oHYScBNmaLZDXZe6WYnHeX
LBCs+onvEpbq4YGE7zScyylem3M6OXP8F7hKelQigMLNz5SQu7jWtbV2hiZuehgU
IJUqAjv6XFLnGNx7dNd9YpGKY3YOp1uJabVB5qdnmwigflxoYug/KNViQ9xaELUp
pZGx/gvEdf/yqpT4ajFBRHHOnTfWBHuoJQh+WXfom26ASsV6tupbOTkmn5AJWwC/
v80hadfAlZyychMDFy9mTJJ37CZ0Kbllppg/qHRL8jzvV7hHYv8PQ0CeekPkoMkO
v2Jk4pvHw/s5VnozydmnLd6+YarWOC/2gKW1JfUdypa6MuCnNUdXFkd0ESggG1dE
o1sdia0NqiIA+ebUh3yTaHHG7Wkc8Cw8ItPY2HElICbOfVXea+MNOSxG8/QZ1u40
xb8fu2VLp42+yBSCqoXtJGkDD8hLytoQnP5Yh0KDUyS9zDIgY6nlWvmOnxy1772L
o3V/g1lVDwiqf17ljYfpSpVv5JzJ5pH4o2fHqYhK4iX0WWeFMW3XZ2rz9Cyj6hws
9ke4ddB3m5Bzs/Ve4aJu5bmyc2/S7YGEQNBND+94dKgjOq6N1UNuzgzn3cERhyMs
e04m20JBbzb/3F2qKCq5mmxPd8OZKn9VhE8AS7+5vNgSmdZivfJ33WkLSnIReAQX
K7XGHsdQERsHGvIFhmU5LeNU/BTWTen51uQ+HJ2ajdvFwNCx8pNHRLQs0QMGr1CM
yFAOo9Z9r85RqTCFYRD5mBoGSrqFc2PKYxsh0lc2TnPL0XtQi+bMzwQySEURlbx6
Bfj6Bzi1Dl/RWprcvgYIhPQWuFy+XEdIMDaq6scc3C8zrp0Oq2rKiqFeIoDHxxgT
HL8DirauXY9g0xZkJI8eL7J9UR8WYoIlMnLtGxldpL0oXAwf6wjuWRSymmSRB40r
eHouQ84inGNJhMAl5bomvArHySLQHDUI+tIC0Dk0PmNzY/7bkeu5/PSgu3LWzRgP
7nKxJ4cSSOkPiXc88hTSm2MMa0drHPDWmRCqHSAUz+qTPVAvRAlAqpOn6qKop1H1
4Hq/wdTLTPNkU3lM1AwwdYVBn1TYMiTyYd+sgTNYf+ATF9RaAmjlgK4aBrDcJJwE
fH4/xONMx0y+KNmX/02q8cOwJvJ7saQqb6wJ03VjlNNIeNSKq+lgzPDcZsdGHIQU
kkG8wrhcucjW5vbgPyjo5wfxW2UQMqlL8hnvOqZ6eAIHGoKawlO2d1FD7lJoBVqu
Yo+9DYTBVWsM9E1EjpWZZoayJCSRu2fFHEiwEqZdUI0PFdhLNXS6K/2cidc//OR8
RX6FPU4KZTOKbJ2+GI01cuSjJ8VLVcp4JK0cqvD7+fAwJKhnlaXJSpATR6mLi8+O
SlyqakhkeYVh8Ahnf/QcQp2utvDxcMVVDk4Sca5QTgHFhzJEIG/PdZij1ELArJIQ
vq/I939w6Qb6DFULZXD40ZLYJlU3Q8gVHH268Rb2b7knvamApXpnt69QCwK7b3Eq
jYUeQoop1BjGsYWYB0aQZ7bvZ6DdoE2flsMtYfg0F+B2Lkez+xua1eo4uYMmD8e9
9kE/UzweqbfN6WbCvH76wKv+qieNXth0jWyBHoMiJxtCLzQf6ZzY9xMby8vHjIxh
rL9Q+bF1ywUBXIKVLHxiDJcdwCSQPp2cv30Ei52+2NbXZ/N+lyOouW55bJfVvgpz
7aglB3ffeVm122FjVF+mfgrbJbtzxhe8xywEwPndR2dFx2GqcGldG7gCgddXdW+Y
Y5SVxrUI9yGXe1T1fHo8kOfJVw4eByd6dOKPpykb1mzkn9o2mat+uhRxd6NkZLxh
Ck7YSgeNb3u1/xKHrfr7kkCAuI8LBmuzzWXdRrNiG0ym81TKBenYolY0wz7Ax+vB
hf0ZLxS8R9Z88diki8T2nuTZUYG9hoS09OzjPeMxvOgM0jspO1yCJox+FmFuEnq2
4qGJddlOstz1QRxyr07E3MInHrnGtOj83QTXFnkcsyWY33imTAj9icDqfuLKYY6i
UDdu6ZXUeXC4nTOSFca/p0lLR5mkay1MmWMBivzGNzjbcye6VOXj/Am7hA1JE27e
aWpwXy7uZyCNN2WW8yQg9E4RWi7jXHJ1rWkGLWIfjTDnsDrUBspembJbHuzntTlq
bQZa9dmw3tXpcDzHZKhT8ml3t9MXObEWAeBby5LyGdUIcYJ+q30TnW3z9hF6vRUE
KIfb47ndZNx0uT+1VFnF8tznJsjbdvKqKQBcbr99gBTHCvwvIcyU8seKgn2i0j5m
TxIPd/IABuhx4hA1DmJCBuK2I6wKsgJYB3fTyY8l5RyyXm1qh6A5swqwbCfGXxlm
OoljCgKRMMiQzyuM5M2uoJxAkGyult+ypGEP7KdVi/vpI9CN/kUgl2uHuBJBxKE1
Eb3tfGoH67PiNGKSx5feWR//cFAk+yhP+UXaz9JTz5bJUJIcO6c0uknVjP3JPBBx
rHmt45fO7UremimGMCAzfoqz/0z6YcvXg21ILFMbSfZN22bFsZB/mvJMiqSSB/56
oV6usM4ycpHg1CR/EoD3NOTFxDOeKd4ffuJQKmLutrN5vHC5HDKPwZeNGmGo7nJ9
R33KlvT6SxXzLb5KR6eGLLAJsI641XI4nrf6rP+uhIu0sOrZ4b+ak21nnAXgh8xp
s66XWwGOHVkHTVb3fLfa47UNECI3ZmhTuP/ap03CmARH8awHZaOLvxoDy8Edt5r6
YC3NBxDnQ+dhsPm1jpTTY28QERHsKnvVnN8ijTd1f5fL3PvCtiO5blqPa6FjnryN
CJFWD8UKtNJfQWcxbLlRQgkJjVdHeBufQ1+9lZI3yvtWLEbGdAePf9scCQeVedi+
Q966PoWTi1ABoilZb/E4XZfpNQ/uXkPTGXg6iDs1z6Rs1rRe/E0qL1BcCU/+hLQp
kb0/11Mvf1gq/85uBBdW4OJpGDXiHacpPRCChCr3yehPpgBWWRVxVAUu/vvE47xF
oyKNn6acP0rmYAwZRrWws7s2cOOh9aLIdZmnw700PjjTT18augna7ruQlPyBoTRO
VuBdQqMyiXmCTR6If51yOigMhg/5wo0aaeQGBg4deuBaMoFfkptvBftEdEXdd4SR
16ytBv6/lNx3AG+dVyoRMvgMxOQCy/qHc4gVK8JYTk5I87bz0yjAYgO32xFjA1m2
gBqhthrNzRNAhTL9kuRWILwz77wkeREcl7MW5HaN0zEVvkwtpOTLr3Eo4ARmaz76
g8NHGDQcKDSF73b7lqHpmlRX2FckooHZS+NITvePFqoOKYCFvOqH1h4I60aPltpN
Wg3ONKt8w/hX1HMp/yJ3/HyU+hKTXe7ztFPvok1fqUg79CSiiF2QprsBypJpH1bT
IMNIdgCKw2JDfysLpRCxAIcTMPM7VnstbnxsQ5RBHNG4zivha7iJZdSkLQ0DqlY7
OYNb0vjD3HAVhX2wP2T2tTzUOY+InnwvaxTEFL0VcJxCQiK+1DfVEET3iR4JIdJs
dHhIGD3Ycp5bD4WMnt4xe+I4gl/g78BD7tbllFjKqOpeJ1g6VfqMOiNVfcp0+rHs
ypihCQ2XkuRiSik2N0wJxrzApua/KtaAoch3137D3ln1OXqfLP8xdawaKJZljDVc
R1IamJuPr7I9kyGX+k/cTd1FUCo0Bly3vLO9Gorc8nXFYc+CrA/Tf5X08Gklu6JQ
a4QHPMBknR6Bpi4sFgfZD9fsdzz8+pbWu83mgHBwbzBmUmL5IfNZ1QpckPknr+cl
adnC7k0u9cGqpOyKyZgncnUNuhBPFcwEz+esB4ObvNu+y7osZsQ+k1kfRXP8YK8s
mBjbfCGps7xLyJzRrnHeVxa6t9UDSsOPsdbE7qE0g+35XF5Cra8IlC1jfD/HkKjd
J9WafiTbT9gDR0yHxODtSviEZB/zmkArIUzEgOwrjfqH7IwFAPaoRllnj4NIhnT4
a8e/B3MmN0UDlarRAbsnTKz/niUV3Ujd/Zvh4VTdWkFM5BcbOTYvXq5YkNwcNdl9
r1RANCvUe/KehAe33/Mm3CFGm/cF0C0OQKaGVOroKCEyP2TWbB2AFR6nqA7bPIt4
iRJ+mnUgPUJCXfrJ593t+sBE2QkokVsnCPtsm+H9bAGJODh0Kem8+XLmRYT57r/i
fI5t7v2ogRgzopHzVuF8fA7hE+lsir/0/uCuKUYkhE0ed45YzkZQbZJvlFIL0x1r
nzkpKwb+Hf/zMzkASEMfIHL633Qn5aJxXiP3Uo23mUirTRXHMyBhP2OGTv4stxSb
EBMmwSsYlR8bZdQCoDRZxtQeeW5QiPqhNHVRdX4SqQsqa9qQd96AJF0SUM+jqi0U
PlhlOa+csqgRS6eeBZp9OOZDaPZuId/77THGDdz69s8a7sUL6BTQwgOeVrLx/8oX
RPbGstB2og7ak5wgUiceeQsMGZBXmF4cT5KM0iOYBfXH9yMjS3P0v8VVIYgDea36
3uxs1Dsndmv8PrOO7BTHkiWt3Ni8IyMibTzlP/mkChj/4vD5yEOvELkixk81X8il
2OOHp2uwV2ZszHsVMNpWLoBRVO4hrQqz7o3Axmi1TJpl1G/pk6zQ/P25CZbqLUYL
Hwzfs/7DxkUg8gWdcLvGvKGicOQXXW8m7yD2uyGjREIEeAjDUEh9VC1C2LvgsMal
ZI1auqifDWSMEY/EhU6HFkqUVp0ruF9gk63b0Rdij0KlhAJ4iDIbtQTFyJdj7vDH
WkAVOvdEM5lfk6sIipn1/PRl+q+lzwI5O4AXmwtSfC+60feaJ/+sc8+0Y4OKcZit
jOON+ljNz8D5SsI7xli8JEtBR4CYwOAcqJ0aF2snWECHClrbgJda4RmlfV4qt8eF
s/9S0OvEQxM96sTdvRTCJ15rY7Z8B8nU4n3VyHUibOfbTqvalEw958sQkATo2t1u
ysOQb3V8S/NbdzAq1IVtT794LIMaW6GBG9Bk2SeWD4CmbEAQ9l19JnAl/SAw+Bc6
NZOS21SNvUJKiazZrTZW/8rHllOLpH0kOxljSmJz52V0P6fa+x8HlvnziuTgVSLf
PVYnIv5MJy/bnOstpc4PPqHOEbJfkqWV+Ayz31wmipdrEL1JT15KtkCSzV1Gleqr
L7bVMONTcUdhzDlIKlCox0s86mRunDzzB1zHbj7Zs+rSv8AZlGrC9HJKxmUkAK9D
0KmHu2aWl3m3NXHr7g38U1u4h4SGpPzAD/c0fItz3uhpFFzOu7o2SBrngvXtlEMF
0gTXuWPN18nPSzOMPReEDqZFfOVxv7PP/6RvPPLQT8T68EkYDbVHyE4vrwcG9KNa
kA55Mm0Al41wEhAfioi8exj4L2g9baAtGqp/6hmQ+NMvnTXzC3HMn7zySQ16MRR5
N7sHCvc0cZI4UB5C7Yp0pvAF2VIehIu5eAqp6+a8s1+HPqK/DkbLgurMvVm56cbC
ZYpvdlKRijny9vEIvW8vs1GnI+QUjdASB9s968QJzQA0z8J6mMuF5ypGVPmXOy+L
9jhUpyEW1o4kM4b+l2Qn8aPb1wnx8hA1toBDpeI6HmP5mwFVQZMXz8qTwTw8TENj
Yc7kCVL3x1TtDpNrWZ5dJTO55jhiEprRvD/6rbPRWeyz7mfAUOmLPItoKB4iEl5F
qJ+UWm6c2XGSIfMooRJVr9rOTWWzjLQ7knIzLBsg9TmbSdJQVwcEbWB947K+E0Ax
26+TPnZEatYPgaWLRnHo+sriGpiCTyjWlfGxHbaee4J0C7PAQewmoHQ8dWDbjQls
ahhLEsEI1P3G3MHo/cnJg2KwZ+DS/xve9l4is5213eDc+gZ9lnRexr/i+4oY+kVi
DpNKVDDSrCxYMPAIsAef8JqXe8l3XpVctrB6CoSV1El25QbfDhHiNWUy/lmQ44n/
ytiCGPhxJmwcULSPChCVhDvsHuwlum9UC3/2KOdYBlpygbDpQlXut4nEtigfeqaL
uGYBF6q0PTpQlb6Scr/Jb9Z6tCqXR/mzof4QhOIrHBwdB3cRRhirJN22KAar5xN0
Kxgl3mkRuqRbIGGKb10kODHKMh+SBdl+D1ahYCONkviLgdnVZ5mSj0u8avLJngDL
GSgZOHbYSuSAtnc+SLxXOaRa/loruNSYmJtUHIDU4r5mbN5iHiwN+wi4fC7sCeex
OceybHf+EpWV2o6/R91+EE2rEkpH2TmOtR1IknoQT3Aoy9whyZifb+LOhOJuqPu4
OQKuMfDKZGG+4WPjskFuT8KmFC8xlsKk1SBCeywd4WXjrsC2Z/pe3Ub6u2FLK60f
CvqcveL8xpIj8Yq8xStnmRTFVn+9tcBJ0IoPmj0q+VGPwO3U+HLjF5px6JpwRVS7
edyvig4O/DBXr6guiertsyQcCgEUKfxzzKzXlMEkQXW4fG48MZOUF7Arl3k/3UHi
rIaV1SeUOxm4+tQ2W7PcIQcj+whc28zyPXUOfrYPCbGUqKGSzwUOnOdHqkQYQIEf
2qjVTQtO/eTUu2cODlh5EdKB/WZyfTXT84r/7ZGmvBV8EiGt8G/T8Vy5GX59A7wd
ZwIoNTgbsAPUEHSEXY0MyIG4dl5vC1gzgu3tNMnarFWlHk3DcnZIYlS146xVz+59
M2BTkRCQdsJFvS+UY5wN6LNzOiYgN3cePReGvtbUD+FZZqrJPaGpo/RQmeyhN7lL
d18tJXeEbRGjnhWm2uI0yjtBI7O8R4s+gfFN8fytfKKObZhUQn6CFYj5JbBg4EJY
fnZNYfnJ3WS6CN86SH4HrZcZsDAlnnYBcwG8L1eAUVSs3hrrEk8IdDxNqhtKxZLQ
p1LaYAKEDJ5jz9WY4NCpafUk7FJ7+35/ob0kVqhDzPD2ASJgrsUfxmVO9ZrzIZS+
R2Jlr2CEp8zQLWC2SIfxYw+q0lkMC8HtWzhdPLTqHRqoYo5EOPWGtkJPHQSoxWR5
7qqhEMdlN85j8j+oBqAai6LJVuaAkC1H4jI1FBDqBqjHCQSook0+W3nI85Q24/l0
d/AKYPet8q9t6hFJI7rxtcR5sJJbRu1elETb8sn/JB9/A4kGsBXaZybswnFVQnYc
Ce04vTq2PO7eomutM2qO0Dj+5f+WL6/zvsV+jxsXLIyxSyWAoDOicLaWi/Ihc6Ls
TkPbVDW4+hK8+Lfgk8+GtDZRr5DRy/r83y171Vwpuh0rSxvqxulhEIbLK+TD3tgt
/8PZ2rvYHx5P7gQi+fPhppZkj8omuTVeQY2ndKHbGVCgJLYRDmsoqZMRdL+grZV/
uyHN0q0BzHw4zU+X6oHKOcq0KOeWg3TbK99X1TgoC5WAYMQ0FMztfx5Hmex/2SEo
riXKB34n5aLoofewCi3LpMYP1EELFDP29h+qvAI1DgIxDD7oVW7bBXtkvXNKk2jM
x4+eWHzSTaJzsbt7UpNIhkTa4e08KbldjHNaI/KY5IM8TJDe3SmY3cKSFWlUPx5Q
pt8sgsrxmysqMCXkF8yZ59/vjMQGluFRG6qa8RkfvyLI2GiL9mu2b9LuelvJTMWW
MczNgDr36SvTscYVNcPmUIUk61QDNd16JIl0FZqHj8Tljo+busSu9ETvCf6fTRnD
3wB1ICkYbphx6KsWkBcQ5rc7RcyhF8t+iL4iAWl2Pt5wYcemICJE8lL+lKo3n2a5
ccri3ipK/y8ZkuLHEpU7ekIHPY5zvObGjW1sNl3lUP41eqrI2YaQn2zB6YH1Fbg9
sM694WjzvkIEkMTxIcJvMl3sXAokrU0WClgLrG7n8/y8IlAQThsDu9dwJ1xJh8Qt
fGi6guFRCW8ga6ZXem3vIDQst6dMRerHZhrou9+kiovRZ6XimH3AeLjhcjnf8cDZ
nLWXf78kUcglKhPukogq2wm+TYTJbDlVBVBwYktc5rHO+oAyU8ozzCq0MvRr3otM
h6+JLv9noNPzfr4xesJ7owX5J0CDYu+T2Q9P7XjfZx/nkjGUCAjQe3iloDCedED2
fY0/im6+6Ba9xHC0PjFXu+GspbqugsJK52xuWP19VjG4S7di94XOu+GNCbfudG2l
gVuWQFHZb7g2UR3emr5fw66C8clOcMR2TgORCAMCMHwRVoCZ+c1PA6b4v3E6dCfP
aOud5zGBV9xEuNRJSPgpq/CdbdAbwa2AWosikmQkesBkSpsQ4tMUzPF3+vwfmHbY
n8l1LuGSb0BBbPnXAfNYK5YuJ/Kln1xAXyvOMFbsGe6aLzSQk8dMnZHOJrHKbWdL
o1I4UYB4/bzekDs024onm24N5PWlRu+TQEXQOTVxE5eXqnBp9Wju0VAYg90ADjJ7
LVETBc3mIn5b8/RU6GpJ67Mkbt+iqKitEHA4Q3YS4+KHKe3zIX8SnLAZ4eyr7uGb
lnzGoMJ37ESZ8Li3falcN2sXX6AQ5awq7temAuH7fl8hM9eetvCahz1d1shw9EsQ
lpgCP72RKfA+9o0znWIlRMhiflkSk/6/V6vmcwbEMexCShs37YcShvvg4sT+bPjm
KgfgX2yZoGhFMdOick/YlWdAO6ETJsZAfZCbSlf6ItwpIADCBpVFDVrovE2di+5W
YEfeVyf6GIKQXrmB9wdFyg2yItMCLt8DAAvdH/jw1HRjtelcRpbuWem7Q+MJj2dF
tL+68D0M4mfdgU18tMwevgUIKnknZmKwaGMaC7JQL8xCsv+G7vyf/bA3Y4Yel0Gy
oOtP5jlRONwGT5vXPf5ab8HbqXJNGGVLSGhMce0wDcrKzi3MX6Pfm8ZCl6f5ZPN1
ljdt0ZPEalIDdjmhaL/KuCRny5ydSLw+mXhCSpJlQC16VBT92FD6tL+hbUaLHc3R
dt9AAYgwkdO0G6OZheG7sl4aHixXN/Z9HdeszwGatvqUjq/CT/DuwW3z0da3IvsB
Bqy7ga87P0oHcpt9XH9DSOWCztE55h5cB95Kl7EU2O00/W12C4NTlhq+gKT5Zyyt
EVOhpayV1GRE7zozXNIOOhTgTFiiFcNzfj1LAixBODjN8y7WKE/DMibnW2b/cvs8
TNuf3XR7Q8JQotoPtl+uWkHuHKUgEjdJ+e3wITjHX9nB3EFdBbUj+sKzJ7zPrblO
mHM/We+VH/eE/L19jsPFrGbCqb6yHYkAEKdRo+7R45hmM7KYfUpvm2zIQHZXE5P4
gcE/ywECgopmA5M1M6b9oVRusFe+rlDJgDN5KbkzP5AqcGc88FrblLYcGj2F8zzm
2STQLVJ5QqU8X6i2MxnzCcmveyV5jqPlHMlq6Q/1AT4QCmvcZjE8JbvWtWrkn8du
CcupvBKgkdIeN2n7b5fVb/w+C/C4U36N+O2Okg67fyhM+kl9UDsoS8wGy5yetcSr
eTRlu6n/srGvsnz322fFQ5UdTfNIWYhSL+rY0ppJOQ5IXMGGPVNpvvP090EFaV1O
fW+NRX1e+9LP9VITjGaW3E34ad0Cz5MchNhmyJQK5eCSgomujSweVH5nA6tqUmgB
Cp/GfiGT1JlkHTA85uop3b0lcZkCZUIXF6S8lx7ktwap6WfMpwp2qadSCA11XSUk
8IWoGXUIMY9nSMunsdz3XiCmxKz+bcBZFyGaoaSQQRKZmQCNnAqM+atr2utKPd2W
rd5uxtb6rp6PApKYydSbxPhJtOKP74PeNCcqSLhzOhW3xccDT8IUCWfImHuJYzOf
HnyiDUtQUz0j7U8br6Kq1c8v1DqF1ABYR2oERRuCMUnbe9AkF4dONIyd8uynPeVt
gmPfiN+3/zA3tM9Q3uBBZokdqBHd1kvLJMhZxVT8gHOiP/k/xnsjQNW465odTEFR
W/rC7szjTPIzDkqn2WYIyYIPfsV4msGU41vDhjOvEK68AAmQK/13SYeo8LUG9nUu
u0Y7Q58y+1tpgqWrlaB1bVW8nrPZvGlRKxf5DcPyY1vo5fTA21lo+NUoAO/G+sPw
btsTr/XjZn3zWEOrc8WVyqln87tQVy/zfN9f/8PFZpykNm9b4YeuRF6rIQb55muR
MJtbWHNLZi42RSKwdSBifnGQzRqJLqKcetwD+nFOWUAvRHqtb1NHGRXwVkh38GSE
HZpPXQTvrhjLQO5RCVq07d3RnHzM/xoacdZpyOktN6N6nWE1n4Nw3ihyXGg3W9KM
8tyhlDwa4hXs266RYQZ7S6N+Lpsyt3HTDB6vF3pD0Z4zqg0S4/LbqpCMAY/78Jpe
Sc4vHczH6U8Y55LMoyFQc+YhIidmirGyaiI4Kh6QZPkQbdS9G2WtuTDYhhpG0B7N
d3WpO0ZzjnUZNmpqvx5KaMkMxiUqktC4bHHnbChxoZvcXe/Uda6QyarjfF0BkAmu
A24bcp1bFwinTSXqEPf6yyAciBA3bjs+MgitOm/ZF7GMmTwFQib6wLz3Utpb5vhn
w2B4EOvs8IaObDrdwS9H9oykQS1/pvFTyXP2NrjzNN15eVfOSYQenH2LVIZWSO6u
H7OUArNUQHr8jbVSUoxxOSivWm5yeGzeWSiV+dgwadg+B4AAb1Zy0CiMmut3WqhR
BLPNReFU0fnoPn3x2ZshTtNt7oB2xuDUxJDmLsIpw93a2ayAxh+EU9KeGULJAGzf
fAJWZeOYtyK/+CH3NU+Hz0vlaDGgCWHeaK/rveyHKNk3HVF6Cnx1QJlXckI5L/63
+d3yyJYAaDYOzK8S3me7ObH4xeYwOwUSloRDLI+359lqt1hUoMCGIv7hi4rInNM5
xgys6O3qDCvtqGsclFs29ucCVGFOB3R3pAYVpfHjQ1/NHt7OAfgttAkJXKwGiEN2
eV4A+5mo34pu0VIgz/H8chsK4JhNMu1rEpig0Dqdt0fh5HN7IykaIRmzcCz+MTxr
1/ruJGB/t3dWzjAq2BYZdaOW6pVhiy2lAvTQIdy0dnUHQNuWDGLFsBCWr9da6PdW
3ciLrripwWuCrygur//IsLeb4YqkmPVx8omtScYGNoqMAzflLtG/mIDACUWUXqG5
w1UICxpK+2657WBja4lFBs8liqQ6D6hbg1Zr0rpah/P2YzmQZfYtyExqOw/+mDeU
H22HV45I+PV5W3AA/uOGejrzRLy7ltaKZMgd6DqJ8xH/apMxkoiRZSASVSdZOwBS
FZWd0F4Ju20xa0zjawxVdvbnoTuLqZlGFUT5K5VfoLvb4YKjKeAO++RZQqTeTMVF
nU3DWAASEWdguB5J7vdXBHeRT0N3fW1n3SDgQ6kWV25DyMn0jCRRSAF8NhEjkk95
BESemIpg3c5kOD8mvQkXkxd5QSqEKNeFCBhyqLxTJ3duMOqPax+sZ5VAhvLkwz0Z
g8QqSJZoGfQ7ZFkWA5SHWPFfyRwGGuBZeFrdtWenbffkxmATEK9z0DSbctFwFGY8
9FE3qxvosB2d6GFXfVN9tnx6hHcpPOBuUUNRCUKVSPu2Q6O1wv1U0bpj2hhCZycy
mA0hODPJfPPo9mYEfXX3S5XScmvAfGgb5QUzhcz48tcpF0F9LwQsot9HaevdFls6
ikOlPXVWgJ5BMn1p5fcXKaFHpeCXEzmXyjMjatF3/v4TymEpqjTb1ZBkkCW5N53Q
kko/khxdZ62n+gwj6VrXJ6sEcdAmS5XaCU+xVGOQJTVw2nfXdTvxS/AwG03XKbqv
no0rrIgJ0BFDzLnfq5IGIh1nK3P/WNu9N+iDaIeouNVprypXXmpxVARZ2sfQ4/SO
siqlzCYAycBZygFehd5c+vzTO+Xz2vRcvHUZ7TH8awTkp4rWbafNjJb74ym4+HV6
mmwQuFUgleJy0HnobPsYyn6XzJmTmYJTl0iUWa3nGgWvSL0qkw3qepeMUItXCDqN
1ZQA8QiPT71EIUgTPKTRH+3Hot7WlDq5FfMO04UmvUfOBmQ6vvbx5X2BI/KHPvWg
ApXmgDRyWbl9OVcC200vD2ptSbPXUnaYyEO+DmoLVwN4TBw5slisekCISZEp3a5E
fM1aozKdihstDxTb8UxfzH3GDS3x+AV5r3G1/1q3jUZYSJTJgi72L54J9d974uRD
1YM8YSABVtLIlEcUgUendLKLEfN50FoAYkJV4U2+lwvQtTcGnNKdoBnzhKj/ljrN
2+EKYnaghyQE7c315fJ4l/O3IWRjTkrO/+oKjDsS7XBk8oxzS2d69Wucngh2b54i
n5pM/Hd+/pxuTxEqxeM26OHXho690d9Oal8LRQwDIPectq5HTSi31LlCod/asLvP
IaF6isre2eM14UMDgYgLYfsIOsf59bIOBQJsjjHprQT4Hkjb8Mhr79Ck9C56ZW/P
Nu1ALhnFfM814oEEhD0GIJzZVKcuPyMO6JG+3IzcgWuabTjXU4Bc3vDdbheN01+C
LueQBmLRs1gCPvfkly+QuWseHWTgOyH5By0GknBm+SFkgT4YeZ3nryHJHTUty9Nd
bVgah0Xo7BdbWUE3bjxiNrVKIZm/SdCP1emIk+aH0aZb6n8S2/oQZqd9TQ/v69o+
mftvxV38ifz4JeaKp/DbJwoXLDBpf34Ym1AGuPhuWK5ZU4K0bqIeeZcUTfSdmfDY
5TkKe0IJkV/smlaA9EqQnUpfTXymhSKgbT85k/NuIbr00KBQUbi+RdebyUBaAPRK
XSttk+SZHw2cZVEMoqOr055XGg8bah7jMUpGyZFyRdLs0yvrtyBiyZmyGEBYSppN
Z4lRfFDkicS/csoeDdJcuIqlzbrnblG1zXzSlxTKQb9OIWHC42So1J6w2iDuUIaG
WgScGmY8npnieSrdhOdXtAbBUDmhTmvqh6r2olKUogUgEyoH2bwU2I4Qze38kzVN
ltL1d8MUZs23eohFxk9sHpFP9ZxML7VOav/AuXcUpvi2Cao1PhOJUQlqia9UhB6b
+4yw4MVsrEu0IOV5aMbxnnZCTvVQUAvugUU9R8R8HTJktmjyM9viJDwdVnwpWjt8
0deXv1d03rec1Ry3Fziyo8ztQ44shYAesV+A+FVqJzgC055AX7szAe4557oEBTlz
bdZJA03gSWClBj0ERrSvMk9yVY/Wx67DWx62AYlx4CzM7EFPXdIouemOUvUsUbyw
RmirZOB70le1pAEdAHnkBqOLSJbe6bsLjfObT84Kith2joZElFOwHDXm0gsQlj3A
Oeoca2GmuC6zwu37nXCAg3/GNFvEm734u44Ef4oIN4n7VwE2ZizTxl5hWH15uClh
1l3pyh8GkY6BKdNgYhRGRswf7DeSrRbBSLPkXc6ik2PfH1poMJE6LdgZQPxkH8PI
ip7mRVXCwKrV5lKk0r9rllR0e2cMIME2Dn5NTwChpB71r9KxUNBj2pnH9gBD0ypu
EKYi/h66MJv+bO11/QBf97iO30wiqF24UdXyeSLQOa1krts9J18+D2w2/5FO0V4U
v+Novpc4IarWxbsZQoVbmy+NTbvSNQtQPSL0cHt1jbXOjTXCm8GZ+NpFAYpNSUWc
2FnVD1gneMT7SCzqiqzULyPvyB2GpF5/B4Yobb7WBvKQagMEVl7kmVDUFBLuVook
ItBFWJ99BDykuPjNVXaz0gVzdpomgs/74Qk1CiwMJR/RBxbnIamjw4ngEBVMh0If
R/aIL4wgjtsriB1P4XKsnEegVz3knZD7lIFfUGpLw8bm66VqnTnC42vw7kMspMcn
H/ZK7uZUmoTInlVH1XVyO2My78KYGIWDMBkqf50zQJrAXejj6HGRKE5LyvTRuD8U
QRcrVSCE2bpHvY11ZUvotDcfDYOhEjwWN9NTJO1+hnZUeGCfiuCQQIXXYhdxh/s8
dIeGvSc8J5DNaEqSUIMtbhKqStugwM4axOWGuPk2Hl3fXcSnikLaX+2tQUs6C3lW
g+wNR0PTkO2i9Ow7qGdINN0DjiYpNH8yHVc2DJsIhCP9b5vUctqJSAxMDupkOPWH
v78tvGGA4grdhj/sj7gQRh8Nrb2nttmH+M5PZnSEimdIZIYAL+99uPk/DEJR6ymi
lR8Qq+RC1aMUQhz/ePfBZkT324UvMTmTZLq6wqa1fAAPfKaHzsYNw3+qzSf6jFki
E2f8g2mfppDu+5dKcIgjG7mrLlRnq+NvfyufbQlOhOBNji8IR7JT5hs26+Fbe07a
uuxj+DLJfVbwyggrbivLQduuy+tSx4ASzBCUXnwXlX3+iH8ooOvywthcRWwH+Ywv
li69dPXysk7jwtzzsBJBjtUTZzDDt7oZKcTzKnZUK3Q2FeMxO9hQec7m3vWRM9Wu
hztUKICU4NOJnmF/hFwCZNK21nqRT7WZ2jqpLt1DqiqKPjXtqAKebXsa2xROvE2w
on1CDtewVa85YG5xOaFwT3u50HpJoAcPXymvFknmPj5Dg2m0yNQ/9ri3D8TIAPT+
r0b5pnq1HLjHSxyQ0TduIc6CisgKSrggxXhPXAq6slScXF8YPgc1WqzXn4wjKvSq
WEnnwA+sO72gUdxCxzBntT4I0+YxGei6iDLhduZ4IQdB+V1B4VuYoNsxc1BbWGPN
FAjm9/P3fx2DFH+97inf+4Sa/ig+XOkw5JT1CdGNLvrO7aB/bpa6/9RqmcJOGSG5
5zgEj6YltS6HNe6qdGJLCH0NiAWQC09tzjSTJvAnwlTMbqORRjmfbQT0sb1vkNm6
q5BRpf13Uats2aWGEXBYN4TbX1adQ7MxziVec+p1TmgVIQcTBIY8jCQEutIxAKPQ
ht87o6eWGo4HuO7Tt5AVBUs06RFfqMn/Qc8SavKmPEsAni/cQJIkk+scsh3YjUXo
2kffdm5IXLYkQydCv5g08rwHh+zY7C0bdUhH6ChSvmSp7sqp5EXI5RCh6HsyUbTn
BwdKJ3GJsfo90Ye3GkVoW2MYCBW2qMTeJ1iel1sOXlYrrV6nl8eTgGsecWMbZma4
4vn4QIJCEaZYm2+qV3a+4WJHv0hHOPEGZ6/F0iTWTJc/m4SLE7D5l0q9Qxo7Si5j
n9Gb5Zf92jH9SuWyTeDlMZBUW25mIUEfCcKUUrxsEWV+KvzVgzlfsMPW0s5TSZji
4hwlEoeUew7aEKiiV9ZS11sv0jrMMLzImG83L1IeWoqCKj45Ur1md2Pe1j2kUdqr
5pOOmnYEiICzbDDEzTBy3lB6tV2r6Y4fT6f3CAtsca+XtnWqoNeBmT8agna1ftzo
lh3Pil3FPRHy2HBwPzJ8oQb4txM1ezjrslJyjNBDo/qcPAFd83T6Ic9/SAkMHp8U
tTG3W/2PQD8XWX8wGWV3gHTNufCsHBKAsTBTBSMHgdXXJ3NUrrkv5WbPgwrrqim0
Q7mBxOPL0mJp/JdQ420ajpR++Pyi4KQFcKwVQqOKU4bfJneVa6yEp4BQuu6PHeTh
mvf9RfSkA0LgDLY58VyzRq/g+OtyTRJX9/qPGCuUFUcsMKu3c4yNTKfFKS7TISPn
dNHVXPF1+UH765A27osa8vwRLTqCKLgdcwJpAR62IG4Lq7ZKyX6nI2sGmxhhVKw0
WyxBK/isW2FwnE0Awy4s9P932MPaRd19b2pSGDvOZzGcU29VQyFk4JGYvSTI9YkS
FGAPsA8wZQfrSndbD9ebkAFaKlKn54EuI93A86ftl6z03IhxONDLQv7Am/6Zfmlg
Hdq3fKbrP6hzhq8YQrQRQnpW5Z5RoHuTF0KrQjDWnQTGgVWlGwpBM8OqLTKWtIY2
SjUOKPFmMmMwsPIXzSvhnnyWUAM84Xit/2VEwa6rTZZM5Nu1wwcv9K9enRJGaewJ
yKElyxpU/WHDBkLBcbIDxI+50VP4T67jk1y4tdTIqRYFP+i71MguhGPCPgcsDUPA
rS89t5oviJc56sbAzWr7lZrhhn5BuCQrZk0ZkOQrm+0eV79ThDneQmE1UC9B092f
WiNjYXGp0r5+kHNoe/7WXfPZO9B7nTX772graKMKghD+BwfcQqr8byKMXhSLknUy
CNm/oJoPUVaB55lyt7zYVkWe+JT4eJifZskYUkNFWHhjT/dRAtKVcpxulujHpLD6
uG6OcmWmWi8GiqEtUBhH6SCVVy2G7rz0BMDamamYcJUoqQw42I4jX0ns7h4RaqKC
9M3MEYRx2G+iLTiPNBslwQwiW6087xoJjOsZwWeMtJuM88RPijFxhgipDW/KgBgo
+sjMTwN5tMt7qZF6Q2rP2WJUZaai7oSp8T0rp4f9sS3zm4CnOTR/wavcfFC49wGr
/KsbK/IOe+hgh0FeOPC0OlFmujFr4ulSdqktGMD4u4SbFmkooiJTEPA/if2LTFLD
9qOgY/r4KNoxeJ6iKuHz0Yxfh7QIECduRkn3Z4SH/MQjOO0972oxLel0eMTLAN4d
3IZQvicOehP7yJVbTOv4KTSOxD4Vo6XBMpbp3bnmHN9rhTR3oiDxic2Y5St9NlDB
46AqAbrtRnH5BW9baLKxYoViVWqORfuWbbtAwUzaYDzrcguaG/C2BGc7ZSgNs6KF
BUbHYARgwyZva7rLeW6hx0OUURMf/vip6MkOx7tjVmPUpgJMNDX8m7P2qF6RY835
9GA4Q9S+oB9ZSG5JbXQQ8P1A0K+d/adBiRspkXGmkK3vbNIlVMH5bxmZ7e1rJih7
wy8UaCfha0nCSZOF1QN2Ir5nwgurXrPkIuL6vSeBLDFHKm1nCyWA/X1SimkbCs3S
9LyYqRoVLl09jff/dV5vBkiYtrW0xIRu7oXV2e8NQASqOEoavHWW1ACzo0TY4beH
Dcn0Jd3NoclgwlacZilqawEJHKqpKS1DJ2FvCGt87g7u7TqXLfRcIBVNabYIoWTw
7MA7OS3LzPIRtoWdUDhNwDUaOTIhXMLZxhBD7Z9tF/5LNz1afeCW75w+CFoYF9AW
/TF4wrzTBfveqfPcn/7EP0kHt5RVVBCinLbA4yNMoQaTwPyJFbVi6dCxWm3X9aIt
aQ1f1XDmF6Hv7pnWR/8dcvySWmor0WuoJ9DgcggHuaO4Vvibf5NomCpEzpizgvsc
KbUlJMew7bpAMw1y5MDdWQ1jZPs8gqPv4qEx/6aIJZZ9FrSNNLJLI3rGwd3ThP/c
xJ3mc3q0n6H0tt/1z4pn8kGzUIPaCj6TvscJddTdxJPESlKKr7HoCFk4Oqh3z66a
tdGHN2BYHwyawCkbRHn3+FNU4L5NkvgTjitm4m8294exznCWhpWcASa6axUOrW6Q
eXnhZd13acbqPrcL7rC37MgtcNK2WAZNWq7eAVhcsvu5iOo25vz4juShJdbTJaHz
3omA92gdkFWMyZm3wcWj/4BuP77hWRdrMt+H9RzfFKhjUoNRUMRhLNrMZAIumaNq
nwuMPLyS4jtNMEhGfgBXbHrBX1F5JL3GSYdonICaE7ENR8j68Fa0DKci2Gtlvq9u
BFPgDBj7pIc/LDHBjTKNu7r5Hj/heufuWutVRko5fyfGFFTA+j6VvqS7q0v3LIMQ
AHFgmAl5kjy3uvxT7PXj6e3rYkaZwlbdbrwkoHv+P3Gp7a0oJQTMUGzvge5Xeir5
NOXk54jf1I+iQx4hC2PXaNapmfZvupDS6m5wbY8CKkh+a5QfH1V2fN7V0E7LCK7I
QljzdBHR8zvP9bQIKrvfkHU8lL60a5PXZU+q+2IlVq32JoJi7/up34RkrGBPDkMG
7/6Vhqci0pSq+pmUdxS5Hrq21IPUuYrqmgy9JoCs6hC9rIxiIi06yv28QU/bYRwa
cXuJvIJLQpfjwDrwwN0NxClojW+Njpwfj0OnYTwahQ8z2SPv6/Yy7KZxlHV+R8kt
AgMZiHMs6pJk0sApmiupwKdqfP2ZXcnnUVXTgl9zhAeSROReXisNAg32+LpVWREu
C80q5i6xeWiBciZN14eldoHNiXJnoeyz8pmt1VQ0GFK/cUYTFBw6bf9Z9VBlzjd+
rJEZuXsiwkd/P8i5fAWpOMWdap462GMlzqH93cbiDkQbR5rPUQF3mx9/E3uRMH/Y
pA0gydUHZCVelGyETii7bMLYK/DTYRRrsBNMqUeyhsFLFSA6oLOnDtgGxanWIpiZ
GwcPKfoKOYufmY329GkqqGH+oAhHww5m2U4ZtFbaGGZpCdXGUf9B5kzIzSp4n6Is
bmw8M5RrTPAp/FFm5PzjopVb+ok5esBJBBUbQPlUPb68y8TeC5mXwWmfY015rNd4
rLRHy4pb9XWodUrJ6/htdLfcUgo/HxNxyNMYBGnRcbHXc6oZWMDdvbLT7UMhXzNr
/RUmlrghuhKsiY62VYGyES7w4k1q2jV12nA0pYI+A70UD5jKqjuHR9M5lJUQ4elE
Pv1TyW7H2fulcBBn6hadbiWkR69dIILOwtrjhmBAs5TmsJBIOlWn/xYKTY/C83Rz
bwuu9qfbLFt4KmBRfa76cqTskXzbFCtHOz7nJUcj2IMqqFK18ZIGcKEGhxA4kdRe
y1l1WUlgqPEYGYR5SQlfv1TCLMHG2mSksFAhNqX0St0enSwDKF3xVxTiMjhoN3yJ
R7afQ+p4tGe7oefISCO9N3iNZo3dSikmTQElfR40VDnYkaFvgtQCybzFmBZWLjgd
Pvrk/MiS28CrrrblUpeS8CDNIEB87KzmPhEZXhtzMYOVGlSFDqOJaJaTQuiuR800
12txR5ISGxtDvVVD3OYJc5PeL3mCaO26BQWZPEs7tIFLYre1mPokoZfVk4o/oBm0
KIdQ5qj4Lg9sTyewQTeg61/rsG7BAjYUdz/lPZjfvjukN9/m20GrGA7Eu0y+bVi7
7DVRX4eAIt/vAdh1ARuj99mnboEVfy9enjdznALHGIdQa4FuP3WSncv10PCec+iv
bcyj1Ctr4xo+xtPlPaOHVIMX5YKam6Mc/126uF+QgmHZFfgD40K2PF9MutLS/TFC
qZHjY4eBrSqISfW89chpDLTVKGix+DF4RMMWZsIVn2XlsPwcEyDXh5weETxv5Xvt
ks6xSTVmdMfnF/cPiLEIKVCWL8qJ4+gu5jwikcOArj0SHwlxu9rSq+7DUKjBbOld
Xp2bFA6fE+OiuJkjNlr0x5qssVpmfWN9GEThp0RcNXVQ0Uz6c9Gv+QGakFyoxIMp
kYmakO5XAkyEmam229yPIEj0MljfDg99EsSnsDCFrQqfJnA1+JcMJ9HjtE0RmXjD
OGoKqbe1x8YRS8SRm9FzR/INvbk+lAvrxHrVZ+5zUJe76BkpTnP9++/zfbke/9dd
b724jh+ofjxzjzRvCk4HfmvUBl/ZvIyxIR23oPhgqbOL7jrPbyyGFfXdfaiVDYYH
an1PG84yVZ/D1W8VKydJzoVqf0uoauEvWj02/B9mSzK6/l+G8E8Mnbz3mKfgSmkR
+VFvvgit3mGY915jXUBeQ9XI9zXlBzj4oILMj2mbi9bATTcxXtJj4vaJhuLIzovw
mgMoMJ5jB7qsY1Sed6JW36m1TPsQizzxB5/pNl0RTx+FIJaTx6UpKt+FreiNqyBf
8NWomjRw9qo3tYuI52M8+GLfAZDR2RXxiJiFbROAosJXemhF5UWqgYv9vHgei4Ob
XV8tbGPy2DCy1DoNaSsem6ZWO7ClVl5GYCMeVhd8vZO+2rU9+T7kJyDGeIymahvZ
IA71zWVBw6QFGkFGEHCEHtxhm3UCGf+b476MVr3iClI+jEZ+nuqmYC2RSl//PnOb
nqTsrVpwyOClTq1/D6lm94rC4CX9VKwv2LIQgfYNhZtrn2ja2wyhoE1GZpyJzB2a
1n+r1SyKh7G32tlmWH0k7WS3PR3eP8MYT1ViDGwVY1S4pZ3qT2vjwW3zCtyEHoHI
U5j5cQ6ed+x+3mX8trbeI4xhYGc0cQUnMBEYsuO+qISyXh5QVVJCQgz8rM4V5+Gi
9URDHog5gmSY7CDspxS9A8Oillpl/w1ffkb+74JFHXgh2h1o2RzVBpOORGfsOdiO
JVxjdJRe2uQ2vX8V/yt+8w9LNB+uNprM/wVYe/bVUX8nSxlUoetaUqEVZvcvatS4
5lLbPes5D637qmh+GKpFFPyJ5/xFxxWubaKRRxQJ38yOs73P/FxVefcrD2Zp/2Mz
GwerlK5LnX3AnR5RSauiYfkaPc6apNuYEd+6fUiUjs+t+9sp0JDvcL9+cnndgqRl
vIMjzoR2VH5ZSUAhqPPPPVYc7Cbm46jnfoBNgdvafHoDYXMo17PUv7xN6oKSYHjw
lwDELYF8eu05+SJ2YNs7YB5A9FV1stKyK3qolZGkY1m4I+1EMcGb3r+HHfOFIAjq
ufY2Jjlx5WtFxeUWVNlzNIqxwTik16GN+/hm0lfOtEEkU61oUdkWMV3s19SCzoRi
dKdUoogSqa1fgQsIirE+sZGfyOBZptaFq30UQ6MphRcCqn/ZMiNvn/WrWeGHby4j
9TTpby2IGxUj0weI4qUBg3Mq773ngOmhRdthqH4cp3T5yZFybwq4qSG9IsFrx96G
+zgP3CWy7PUhKOd+wIBeXeITgFBHCDUyGpQfBsML7FhZzb0CiIGsqI0d0avoaE4G
QF1IaOGYVBH0cQVma5977keeGKecOcauZWjkUibkztm1B/J27+ku+8rJLa7A/91+
2NddRNsdJZIvs/I3dWSkcqRWfj/+CNoGVRYRy3ftMpfImlgSV9pOPqQdcVr7kZJd
SzO+CJbO6UdjqHEbptO6DTOtyZp66oq4oBU0ifDIcKQLcYZi8v+uamPPc+RCVIEF
e+QGRXuwHGiqS03Ch2+mviW0mIxkeVB1Gu1Yg5KVt4ikIumu14taEX0uHvvPc+UT
DYNGJaWkw19xA2ubhqrIi+Z9ousYokWfVSdJohe36l2j/c11d47NR+YTiTIOY2qJ
uUvXJXTOijl2u0I+FavTLwjGIH2kmEWfCAfua18ziXHSIPLrfVbrWbS+JKxu9j0s
ym9K8M6troD50oE+3HA+pmIIahaft3qUZRaquOe/ddv+qmT199z1CX9xcEptPDTh
7RazfE2Q+rY4OsDu4FewqVCEAgRSC87jzV1Rk+55ic7AoMYPR+mVsXAwofi3Wa2r
a1WLorWh0It7oirua2DDrPGxqUEGfl8hJcL1A+WsnqA1AkMAJ/ust1W1FBDbD5QV
Pd+lt8XnFuWpoX99G3Mm3iVDlLXnuX1K0Q8FmZF+AT6QWaF9/LuPV1W1njSCwB+d
x16HkLs2xVQd7XbBIDIE7O3VKlyE6r+Pay7U++OQZAC/2bstdcDu2/J7eHmxiRnT
KseJ2u8lffeLRWLRpw93PCATj/w6v/KHYExC8KOjFb/NYoLTie9Slg8GGOKoWqPD
R2Smzg92sYQ35gGEtlmXwUy1SOpEV9Rn5rlUxj3Khaagl0RTvHDcwCQwolRcJQIi
zKYTLYNlaypz7zk3OQ4Qhf4fl8eZ3YldzbyGgxBTfT9aF+ZOQzo1/AKZS8RQNujj
L7msXUJnWkXu0cTaUyR1qzXwhfAxyg4dv/4mBreIKAVSc3Latb/rSCDez7jK9MoP
EXP+Pb2qPmD2Fyhtz2OvqyBcuur3nBSBvwX/bv+k5bLUmu7VhnWlTjdDuCGfXyC9
6jbU4/I0VumuvtEiJeqoViok/umx+fvb5d7PxEk9O3fZwtx576Pf1u/Or4o9hBPs
1ZS0dF7Kw9FgKKljvIFR5MesrE11Y2XFSnIFQpslhGteqbxmpHn1KmmXFRQX+7Pq
bzb7t0IjohX1KO2+UYP4dhztjspkmV1WHI5tn/9qxDFC9eooT8tO13gnjXg3DsPx
j2JoiGmt++r9dTyKW6cuDGDjhBq8D9ztT35NXVQbwpLGmwyFdJsM5oYd8NMaxmxB
T6UR12lgaVQKd3jSzJiW6FS9+M4HjPIyxkkvnCbst3eM6DwS9L5sy2BN9zCtIaM1
1kjS5LzkF+hFnoPBe9fELDHxFNpDcVGzvQ97g5FDfpRwAc7vRIKA4cmnOngzDluw
5GCrgN9NAgmmYaoJwHDhjFM4HrcZTCPmRXE56HU7wHbeGBDdSRkzaB0IgsJgW8x2
ZfvnW+obHWNJbtJ/zgtOCsRXR4G050KJxC7eXUbr82mm5QUJyu87aGcaqboMXOJu
KwKfKosGsK+7vhJz1v9r9ANmMKGOqggRAXjoh5AX4pqcIbfa5/b7whsPWjhVtFQU
QeJFZ6LbTvhQs6JGhZik5wqVT69/za/r6orqMcrg8kzDjRBZkfb9uSQmuSmNyRez
8oAdUpsUHRBzUu6ie8cp89HFYZoLMP2tPOdJz/saTDoyxzISN7/60MEtzog+vdzI
7z6sMh2NGtFSDPFgdzUCkSf2dVd4W5u7sOvMsjIhaihsZ0tJlWRs0wIICnOrKGhT
zEXPHG9fKyD6ZZlHCSckaufuFaT9eA6H2S+hpuM/xb8ATRGqmG0y8QiKjNv9eOw4
UX0ctxRxETu/vcezCE0JoP6GSI2NwPZpFsaQOFmY7UR5o0FhkvNq55vqGeO7tb1E
9ftmmCGHQCGDbhNH9oy8MOOWey+xk2VAsKVPP6crUGy/PCPjSy7muscBzcg1390g
fa6N+RILtWPkvCotFqdray8pZsuTIccz6eE/hHZe3mVHXa2Wn933TLVn3EEINmB6
gtdDYbh4vheQhRd0hNE9psP5PjFNx4h/hjabPuM4apo=
`protect END_PROTECTED
