`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8eVmJShVulAPcGEiUwNAuWow9Y3DWA9mzqpLUq1S4pkgmrpDyvgYnQWub7ZluamI
ZBhlf8aFIrzHxR8+e6DLaRH8YfEBZY3qtsCYo6jM1FtTmVu36EbGi88AgBCt+L67
dl0S/OO2IPJoqJ8+WqIGL3CjxUMz6pp5/BNip6JJ3gwXJFDl/KELn7WHZ8pZttjw
6VKFV0Djf5g/Zi44GhVxoAtp6uVFVaySNjNfj+ldc2ytqf1ICy/iqnGIeERrJujl
x/mknrGlsjS8Ouuh2obEJhGCCGlDtIgg/sJTMzQF8GlLfuWRcY4LYmsMNUN/dc+m
gHbBIJKlA9ZTj0UvxKEnTFMp8NkB97bsGHFG4rpAHD/RXktojz2HJSGAHnetOUnL
1MWRhvSDqyB1pkyXmVBkk/je/z1f8SXWSYrgSXEa3L9KjNzxYOTTVGsFfPvs2fQH
/w7K7qjR3SJA45eSRFqIUAIqHyAfEeztFD7UePeQzvHeuURlmPXV3TCm0TunSA5n
11DIFBIpgflxZdHQG2uc6yCp0jmJdsjRMxnJkgKDcxRm/HZcGsCr+Grq/MK1cBcW
Md6ybNpA5EsXKcyfDN9QupCZ8AEiwujLlHhD4nbv3RliV/kVI1+bXaTQ+30mSit0
kgsa+HrxMrZf9xUHKfvJIbpWpvg+zk+O+T0desLr6C4G3vHzklsBk5hRo3Sx71fz
l6hJmwsHovs1xkZ5jE/kTbemzhzfn83i0yoO808TgWYwfIAihnAalTfIg7FOHmpU
IlouyMGpe4nmtSicbTc91tWo73dwY8IG1I++lOj4WEfMovMrc5aKGoavy/ZmBIrx
JsdeEYxSFOc0gPWxC9CQQT4uwgXic38/lJDvyfk/qiPzi9OdnRSPbMAJEjaTtloL
816j7OaML/tk84fvVBjvtrbbB2A/mcxKrlXb+zi9sY0axIRFe/SZ8WMJykOTA+Tl
lpX5fUSy5OjzNhhEjFoNh3AF9R3T0KJN+2yagCvb+F7nRnVFoKQbUKK0b2WLrmMy
nvUJxQHR7uzc+QOka6IDOm5tZ0J47lzRX74w1+/6sIIbhBDF3D5YnSmxgKxnxL+Y
aQ927LLcvCKGu2AmFXgzoyWvLBY7v0/Y/toRBywUN+BzjJDvzzZokkduniU2Y6ao
BBLEjAEvMi5g9txZi4Brng==
`protect END_PROTECTED
