`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
idDZVl5aLU66tHJRcwlS1NsQ9Gwx0cOv5bDp+NAThZoJ4x0Jae8mfRFrx+Bv6xYp
5QZ5Zgr6GQ4oEjCiKV5npmt+T1o2tnaoEb1TfjMB88AHk5d2SVZpw+6iFVzX9K0I
8rFyK0TSPm0Sci1rmvZXyKs0xk3hd5pRmW+SvYa+GcYADThFBZcLG9rlXfy+7Ohw
jBo3fFs8vTGSpIDbEB4/P0qBSHXRNl35L4+i5fZRLz6ZiX1uuRtmJljIqSGZC8ue
cm549GDdSTMH4QfLaf6V5PACg9WuI84GPNGJXTTeQOUBY2/coLP/qtehdYZDWuLO
fa587sdj4/TpmWkbIqtNk3sydNJSw8ge2zcBw6sB9ByHeiYAiPOP+fh/DuTqxtpE
EEp8USWCF66NUb1B4GeL1Z+GTW/qqJOzU3W1mywSpqfgv8OnnDxLqvAe/QbWGE75
aEqBwmzblR4fgdhrL8s7WEhEdNCSb58j+1WwLRlTmPQ3v0ilTSWB2eCWYdkAdbbs
8ytlJbzWw/yYN1i4Q4gmn/xsDqRuTJVaDXSC+EnlhotYgt7PIeBBcSkxCDjQ7+ix
w4g4qXIduNjwcuJ04u2+RhSBvhiQLRZoU5D9Bw0D836H1tcophJlh4811QmJwXF/
TEpKnRvCWBaFUn9m4IXzsYVUGF4HwRZn2zPo9otWVLPfaSxqYFMuTdTEoQ4+YtN+
jXTZrGrWPgFUbR4x323Gn+rU2Pua3mbTUyap05koVdLkvFRYsuzTkvTI/NMo/L1y
LGitFrO5uMatPXt4dS4wVBZ/pKIWa/R6SqHB/timRke7haUvS89QoCDTFrPcnpci
`protect END_PROTECTED
