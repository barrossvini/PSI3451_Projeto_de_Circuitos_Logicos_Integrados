`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2zcoIzcSfrtKZqY48JTQa4s1ib8jmz+wKWg6mCfEdN9W/Bwh1wOs1z6/9bjpPsjk
ge//vYX0V8XMHMPKcBWSny6jrx6f0Q2Q9SiMHRnxebRUOl99FK8cSBlTv2RgvIhp
Nw9naV2Nw+snlpKGRMZy4z5ffKB9dMAr2I9Hd19XlgHlz3JVYTxN6XbqFb0S13pw
GQaW8xxesnzuB6ZX0zCQvW5p86PsA7E3M/d9cN3co0iN8luG8KFyW1DOFiAnMIRJ
cn0gLNmmR1ij5ZWvMeBukdRSu9JZwXni7Hdk/Hcj6I1dAk7hCMZfD6+EA6TPxecK
0kU+j8WZy65r8r2uflC8DvGW6HjWM41+HEFNjby3oXpvQYqHjuD9rdnS8dr5igFR
`protect END_PROTECTED
