`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
guHgl9C2UhnlYQINnoOPDjpOncjcTPeJF7kkgMufnctdB+3As5Z4bh09iiEXd0u9
hBty/amuF4k3Z0oALL8oaoWVMLJy7746KjjCBD6KZcX6RW7PvJZyQaOsLpMX5V5w
tWyFEHP+V6WrYUa6w4n5KvFH9rzd1TawaCerI9MIC4uX8OA3F/KjoOMYhXXoskRP
dKRtcPQ6MGmJnT4g8QWvaDbL64H3m3MnXU3wBDuoqFE7XqbleJHLPkAxbkyTZZQi
u3yx21YLkWlV1MzaULqMSX0Mo717xYhlku3OXl+R/errCDQA9cgImfSJ+Qh2hb5t
azbQGqOLEt1szq1aY52zjeYZuDXAvh/3sI288O4yKbmN+ONDAeqkrUj2hcfbls78
CgujuOJ1usKqPxcd1JaUIwPwciEpovn7gmLRMUiaCaAfXZLx+0KnwB0coAXmI/yK
UGnFpyIOpzmOnecAlMvQUikYCw9rrglcekzEaCumCyyYx1SF8E2vBQ3MIxc+kawh
zPBiqe1WB5JCBEKIZKH6IL4jOtTyuqLG25JW+lfusV+D5yaXzbfo06yTRN+pxusy
HCsDpBugY5YOI7iHKWiLxbHU9WiImDHvmC6A1hfjVfTL04lKqTwf0Pe84TF4QrJ/
pN5ohrR7997FU8jPcvGAT6xQygMRY5rHEaLrQqSUizq8WUo4QNviwzkHlJcdLKve
`protect END_PROTECTED
