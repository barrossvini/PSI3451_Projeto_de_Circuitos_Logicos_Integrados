`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8kJycCHspzgZAxLKg4uO8Ci/Jg6s9K5e7sIfynEvG+Sbt8CjEKuxBBsAAIygxpIW
wf4QOPB8RFKUBoDkSLS/5UIgOm1j5qmKXwf868VBoR9iNQWdb+/vn+Csmdiqy4Be
ssOxK9j4ScEJz8y9eMUZiKky5/g6W0z/jwLJaXmEawyCN3PVO1Y+qQ+HcWQ5XENx
24iujHyZwHbuVJCf1EdtbXNvW3ZesLC1bd74/BTYucnuj6977MA1Q+h91O5Gh+lX
B7XF6b0mh23/6QPv84yQm9I87ySBjd/qigV+1z+h+Kj5eR8Q/nAX9XSeBInTZFeg
79dJC+yljW0AWK356bDYJ2T7zUOM3kTQOU03Fp3mjFsRyBp0MBjiq1TipvZls/pw
JBEInrzqVaGrH+VXzVUeqGpo2KY3J2DnCFKlP2un9kErnr43qTC8mn+SMX/JVIVK
OdJWRn8rJe5Dru6cAImNS0eaTkH5zU8Ni3hbTl+8cMPj7NVamdRSiXeHfmM4cQQN
0Z8Pi7Ea7SKIDpe6f5k/0Uvsnzqy56nlGsCayLGfOmVaOgvY4XSHUPXtfWa3jidW
nqe/E70bNwxhSEH8Fq5HjQdK3ljJy3kIcKVvH1oecM9pPmmzX1Q88bNKUQoMiU4a
iGJJTOqOsNZ+FYy9DZnyDYnCMk6cbeNq6lLtIYRjKjVUw2DzGU6rJSZ7wQGMGLpa
T6JSZzAUpFPilRkiOE8eRP5iLw1PVRIJXP4TnFEHHPwJo5yDUGk7z2Mr3irdv5iE
c+QbaSZaGNZfx9jkaDpcWMhhBgXdDgwU9ZD014sMweHnM9XP7HINZen+QXZcwrHK
`protect END_PROTECTED
