`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cMZnRMQ49JvAN9Geo/au99KdvaZqqhq0HEp+9Vh7PNtxWQlJ6jl7GD06hycpQFjb
KYEL3RZa3wlKeye2bMJBr5usisnq5RRfxUCI4FwZ60j+1x1N9D7wFpyA9Ut1MRSG
CW8yw4lBrDdXElxslZ0oQovVRRzR8xtn3qgbrk2FfGRMVTTTBvID25k3/WQ34Rx2
7NA/RkOJ8OAQiyGijfzuEKwe/2VqkfDWEEnE7tW0PZmg1lPuLkCRw+hA2nEMqeMR
IxtyCUHfT4NAH0pk1dK69tTqCSCTr0ZMxBUwWOFhV7SskT5HLaTb3dJ5HSHWrOXT
IV3uRjvyXym3tRA94obJCCJ7GjwJbVG7F6RBBVhLpCJa2qGuoomW0boHyhBqqO1P
BxLZ1v6qlAGIF53djDoEKb2zAts78wJAjB4cdDcZyI4TbTjrM3KwoJ20AU+U6Tr7
xjgiS3+M6s5Iq+6Tc7038C1J7fIZOdtYCPJOSqnaB9olCdVvmDgXO3KCVeJrF8S5
oV61lp/3ETyVv0pV/NI9gfpplf9osyqoCn8NZ83Z+5f/YigSrbsN/Bt1o/Jn6nQ7
RNDex84EFWSi5SLQs8p5Soli7r7bjJV1CbOcpEvpCCNNHxcPaqY3QP4lu7RYoxmn
E91PZV2xB1014yMyBEiXf+fEny58oeqSg0x6WSqqbRahepVXwEhUi8uzRD5XnDQM
PFnePhSJoUVOrBkJV4SQ5FUV2GSimNqgFNapxWcrzMA=
`protect END_PROTECTED
