`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0jDsr12Y+7DqC3CJONKMFdmFvJQCjxt39STOugX9w8JtTbujmXqcuSt37iLmERS
IrV831GSiPKcAX3Lah4kgUMJNcdWPqazpgrWVHYp9g3Pr8thZoN+/4frH3HHfj75
WagDRA/2HeLjijO5xxbYkwqeLClgdrVt3iFHSbfdb3DEgGDhUqODlHqTQrIIIgx6
jZF53ZbCif29bRE7Bj7e9X/IqUDVkmlQtkriw2pLE4mJe0185Zt3u4pd4FyKcsDr
DOibKUtq8mEsNOscowMNKOgxDw1yLnlNPnoVrXhynoqsN4PjHcXBZVQ4QtWJaYWm
WcSei8mSTkQYhtQejCNgbRCObq1UAnTjEIku4qmTKIdaRFRLUSAii9lVk4j/YYyo
CiqnVyYOyHJRRkJ3fOfqCvCYah85PelM72v+13xXdo5WRvsCUk99wkCCg8cDZik1
b/SBrAUtwxeeDPcHoC2HbGY3DyZzmyxPWFB83NFh6TKrRQVLaG5H9XUotGUcuavT
yLWMJfjILTiwU7c97TgIeKpxSEQwMHp2Vx5Amp3M+8BYrIQ1MsFUPfrYgWDFXAUD
XnGMva2eaWlBkfU5/lhdhwimsAnC8uGQYRSkkQ6vqi4VbPrHCRL/BRPLTjyu9DnC
0w8uuoOI5f75y617rTocsH9iDELgWke1DBNoWYqrZa4AWpsOXzvHIms06FK5FsBa
YxB3b4DyjVjrLM7hk2jxebvIGlmPkbA27S/08FzRanHZzGG9uQ3o54WX1HjYm/y9
5HmjGBViPKtjzzkZqi1elcErnFz3pzf/5a6TIZGJ8mNUYyUnTpwXOJWYnEoBGn4s
3rr6a5eotexXyRANqTUcWrKUwYz71TcBMz4s4xtcMZdqvZbw6qttZyvGJ24O1ITS
uq2pa1wqI/uN5pNrWFPh9R4FAJZ51TFYHFOBjJU+1yRoaHWGJvj2jOW6wZ140rx6
YMbiAvALVbnz9/Cg8MR2PLnV5G+IjguL1FwfnclARfTp19Xb7H3pFj4yLw1Hxp8v
3v76fN3ZwJmZTeGE37A4SyFbHAytKFasrLrN9oVIhwu+UWzRxMo9Jhv6tD4S30FD
AgXlmd5TV6Lzyl8DhxNIubwuvmdDN95+WkgAC7bftZ8iToal3eS68CRun63Xd8yi
G5a1YYAKfRiyhDdsnP73At8OEuOR7X+/Hs6Gn/mYl6XE+5vrEL/tKY9Y0eCAN5c2
n38zxZsQ1K6fBCCC0n81wg==
`protect END_PROTECTED
