`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7uqsa2t9q6Nz8XXUg6h5NJkwSqVpdxXrGwZP4YNeta4qjXeGHP0te3YxNPobNdJV
Vab2t/kMJ16ogjnOCv05PScZ0wFayDQ6xrbRq5bzp5veq93EohWMQDJfEqdTn3VY
4HNs/F55RkNBNg0Q8ckSDIZnr6QHryJEosBIEa+h4VpwPZIjRQGRH/tRIQFbycuG
tRSOuulHaHHiYKwrDwlhihWdVYe/r4oB/kLUr+OlmpBZm/fcXX0mqs8OYOI2EUSG
93hhgb45cPQh5lPw29ghW8CrBLfes0xYszHtXvacBmCOtBZUkrGjnSSBO0lw179X
bevHXC/JXblgpGihPHDEBvlY9nxj9GbblaFd05N/WIC41iEuHHEHTGqUGVfbvsL2
Y7JQHcfSJ+TaGEvAzbl7UJjc78iX1uF6SyoVROIDuJ1EHAYF5RfduXK3wZIy5h9E
SfseP9cjN2x/sd+6z8k7V8Nt9Q3IdvIcGZUg3URRSYzjVVKUGpThIbQaXcfhJwNW
kp2MISg13rJuNJPSUVhEmfAw+5lv230vuZPJc4oVpHRFBZLCELD2IkR/jURa52WO
g5G+49AqVK2j7NKByPKl4CbcVSzJf2Mvxq3NXDlmExLvfEsZC1ZIh88GWsQnwPNA
/CN+R8/P9g6jnCLS52sGNtmipB047KNdQXSxFpCfZ3Smexb+UQxUXFZBCBrNlcdM
w3+85br/TEV6mw/aPDb121P/MRRuCiUZM9gHwV0e7Ov33u6bjDNxwXkNp0mgCKg9
3eyyVXMAqB7asPra1pAM8etwJnAzLHMIrsrI4nAGqHicezP/l+v6C/KWwyBqOaFC
TAoJOOs081ErGJBeICKlpEw7aiqZMKRzfIaq3/M09atiUuqTIVpdVzWsbe+Ki+PO
KWUJG6msFB7jadhRf0scve7B95oiDkXJ1svtPC/nVP7FkwehGzuCDJvMBywC53dd
SK3KBMUFK979f+UsfdLOBSMJH2kIzjjXeK6xnohHHjiNsj0AU4olKAm6X6Z99tPm
/W7EkTJpgF2zJrXy5eoQhbpXbgSA6CifndDJsSgtUZHGs0pQNsTUEF1uOovUea4U
JYQoWxI+jVx8cJ2bSHb7LvvUEpDDQ9P1DBye9OKtzLKC5dboYvwkPAhV2ONbMpoK
kXzda73mcVo6bWI/iCciXp1yN/OyYzl+gneZXVjHnj4dSessBunImyEcV2R22+SS
lSYSqQ5Vn5u1+M7sYWKRyGXdVo/pZ+ttA0mlmG1asKt2SMp4aHw8LrJZ+MJLC/Jx
Vb2I6aFkEszlYXPDUwgay+YlFPLTygKUWQjp82baMZQ2zbLc4qX/oYLHaGogdYeO
4hKD6vdPwQcVwmBSBxCedh/H0n2CDPS03pWDLPCVUK2f9drsj/jjMMizGJZHuBNh
E62rvYeMpHoblGlSnBT+WxJrH1ZndtKC1Qw9pgvsphf5llz1RnUMsSVTDNyflRUk
4Xqqn0D5BD1fOv5qQvGwtxUHtviR/tFF3xU0gRpZEOIPFl6ZmJBT7gwUPY/RUrxP
KkVsBL4FPz8EgAmoWamOXy5L7gxQkIoFQ0VApZRqa+s6MvfLMDKgRBfGgfequ4ya
2FJ44mNzgwnbrBDcS4enqg==
`protect END_PROTECTED
