`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hq2YcfkGTUZqlnPh3kZjtWgXuxD927YxCDPYEkmxjY5n6pzK2KPY2CGKu0bzIB9h
+KN6Tc4rmcdytSkKLjjsS7blExHMbjoe2TeECbkHX2lbzh0Yy1G8xgKaA+tH/K92
O8ey7upGm4qAIaljHxUhJFKk5J6je03FTKan7zWtu0f3kHGSu3dw6rufZPkG4fwa
/O79HV1irKGlLK6JbCxBYEahRtcbwxjdSM9lCnpTDGtUtq9EW7jR6xvz9w6nMJ09
cUPqkFG3hsVeqNwhtz2xvf2sgf+bbXkfkdDWPtMpHhHc+5Imkq7IskzfFB3qIm0y
4McQlkauT0It3XbYXosDXkIrcO4ZcCIyXwje41Y3gy/3kzewTtzzlSk6XkZDnojV
Oqct3exGnpKvAUBlBcRVsosgkBM8aLJAgT6Lg3je8gLOWYoFSz6B2zx//bOv0qwP
JmJ1wSsLxvU/sE/L65trH8kUV13NxX+aMF6f+zhOsa/2GH+ugQ8oFOowI5ozSzDN
+b0kMyJeLTHnxq2eVxOJMdn2nOaWPtXcbgb/8FeeC/mOY4l/ECQxoFlryxFkAPdi
hIMm3qTwufRPHXMu4RvNeOMkQME+kMhcpXNWvnjran/xgIb43fuB7SLOF+1A+TY/
IUuKgoj+Q86MR4cejblmbHCJBFjdixG4GKnfstxMS83EhNo39FHjT1gZJ7hjJrrJ
dzLbjCOUdmta9BYGtwWftA==
`protect END_PROTECTED
