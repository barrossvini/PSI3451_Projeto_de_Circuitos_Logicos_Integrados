`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GipNDJtYIlr9x+FNhwh2FyOhRk1HHkd0l7dDVGl1MZ/28+wvvAbeEFRIxybRNXCU
K7TDwIYOWOlPhcByVtupMDyZy5xBGwpfdtv7HryIlMjLGMLW5Ae+vW2ATyxW/smD
TpZYmuCg9JImU7572N97MfiTsSqrM/6zpA9VHJxLbGZlWvkgyAMe/aixaFj4aGbJ
VeFxkJSdS9JZ58/AvZSxst7yySWKWIiu7VlgtEjirAUHmpWOj6c+MFDS7j38zA69
aoz81jg9axJP8ea7gStXTkcapGkKaK4Q50ijHc1Al2D8h0Mtu1h0TcAoZ2Lc5m2K
mEnZBBO2OKMaZ9d8pqNSvcsoiJ1eYrnNOevL+twE+IJwpxO0REajpmg0PbGqnuZp
5kXWfY2DoBALAGcmtNQustkE/IhVGVZeEIJ7u3BwaIrIUcmg3gKtxuO4zGyw6V37
ctO5Iaz/XGtbaqdWVdmZWgNQg4bcZ4vuxzF1NeD5bCad9TFoCPKxlZXl5xBrE4i8
nlOiP3+t9+vcC2yxGOouq+/pvuVSCvNTEVw6ClghcUMHEwVFCYl1FXk4oGJyDh2K
E0HTLj3JgzuQqSDlEBo4s3E3Ypy8kPE4RX5kcpPxNeeuLGUk5gjptWY6eFpTjX6S
oT0bNJgb0m0T3r2k8FMcKNtllh8w2d0dMcU8cO8fuMZSBFIkPyikBwJ/nza8Gbkj
XHO/fP7pTKLQpnuOdQvzl1fTaYst/VHay4QaRzGqbjl7U3vVVKwaxWPhkx13yhZc
gcJANSDrpFD27TIjc6DucXm5I/HIcMwBU6mvLDP5UILQr4CkLH8J3f7KUP08K4Iz
FDy1ojEMT763RbozPLIu7oQqV09xjEsKYULeNGCEPkVuLxK2FEUepOg+ehhy3arh
lIMC9vr/l9OCHuU1MWdj2jUfm8z5rZbDqFgD6j6y3IVz2JFbBPHYYUBHRBB3TkRt
rROKH3R/nqoJumBwfPYpkm8hnq4yiwDFQRhisi/DvO5ik6dYYbdKqigkZIobtqST
szUF4rXFAOs5ZFI8c3G8DJlQMQTu+QgvU1A3Z62vA5jR8gNlBYfI6YV0GxjRelq0
1iqqLS1WkMPhnvXYCCHBYPRX8PGxD0vJuAFWkIch/ao5q91LA4XGopeQqDNUqFX3
1ga5zai5C71IFcbIl+vSXHugkQIf1A3IWzpOnmA5JnitX1S7jlP4nz+s/m4A3pTH
e14IWTGQiAL2EjbYVpwqUDw8mRcq8aFxLgIPDIFowgeasXwlgGfr3DHBMRCZyrcT
ENNObYvgMpfvBJjRG217SaE3tUXuKoB5xoD7wjNHfGEJSu1DAbIOd59UJSsWOyQl
0A+KKu11N5pxwdjusD0nxGok/2gUmCXAv36Ah11aiM4a2/Zwc6OcbKVK0CbX4nTp
13n3tIN/lSIrHoKfrIsFyhX1ElsjfAIIIVtVIH11es56kdivn7aStTmYmZIpjdlV
vMGoc36iYJhWmT037johUcGiqi7qlffWxK8yq9/2d1Aw4Vc7zQi6fT1BVyziu2sT
GumXEftTqZoCRIDOt9TvUih2eIGHf9dH8Ol3nX5MT16tcZuwwKUAFLTBRS7EOHrP
Imba5B2abtecjHLt5vO0IoOYk+B7dxYPXoJnWE6L1eBM0HPn19tnXech/sCJ3ucu
KKpj+9lDo9TruvUYXekL5LFE1xl9w08JQ/HlQqXDZUnc8LC8E+ph09bKiy8xeJJk
bxuLTTw4rDoqO5dWOgolq2fwZwDFdgFIwtcYhVRU2enjuSSytX+JESgzcopUVBs7
r5t3ZUELXBHML5EKr0ChkkgLkkPSw24QNb3qkjhIVrlLvseCuraS+kd33fKuXY43
gf+6Xa/KvYiuu1dpveDFeNtcUKqzeVJqSy2r+6QhY8jDKRA25ZtTGRKlNZZ+3kpW
iFLnTxBCf9Eb2D6sD/b+3j0WCPw3pMTw/JPepkBdBNMSDEtEqRYWaqLHbCx+8qz3
JBN+co1+e/6OBlHsq8IqM9rAjQficLrU9+i1pcJmqsNFiLudHQplYnYDkj4VI3Gs
CLYuJmS53hmifSCMYNcpjoTe2dRrNPUCODlIw89iBlJEINtHcs5ejGx2X+J2zdk6
3zsCtu/6Y5YFcgUeqDui10NBenlmFGVyQwEMxbJrlhbLujmmn85lc0Nj6U1BIP9F
0vLkGS8xbOevK94ZxihLfEOUDox3Jh8AdWPI520yyL0eu415U4MZjx5jbdiTZrKC
fLBRLhN8mO7giqcSA/oKhQOwW7l5sG85wcfotBnRm0ZT4rpIU3L3loRuSRNsxwVY
bVh34ASJlRqDlHHTNkHJJga+xa0FZ3+tMyNhIjwzISmpmmqN+IMMPIZiskv7ANeM
NSuqvgwH1VGsyvTNUwyo5gFxQzo4GF0bguoG6uYkAERgZh561Z4tqS0Fn/SVedF1
dC6DTDRtE1w8MDw4eNXOLP1O4jb3rp6O2OTWkPmRZ2yR7jYBFUWF0Vb8deluykwQ
kYXxIvQU60HMe9NauX/6PYToImfBainhDlSxw4S1nts9zgdhaCct49zK2op1tAp4
sBJdOUyJsELE7P7NULEvvihB7MqthKjTzCYCQQSNm+pXjq99RQ/Gf3g4xJZvYXQK
luoO6mkYixytb/REtMCcR8Y5w0OZv8O6o6eJsqx0ziYP6ncskAkUBI6tJvMJfGq1
4vn1VkED6hZyqfIbLO+w2t7kqm5tNuGKlxSJA9x9fDTuL/zCsdXY5VP0h5PSvL99
tfNZp7pEpvGSQmMMYkSGIFlhTXTl6dpnGU8XwM9/OS9BS7O1vqnp5Y8jNMMbkI7C
c+F6JZuRQLI9uCj4a1GER7wVFW0AO5MkHgNSiZnthed+ItE7CAB+mgfEM2+kI4kG
JxMmhVohhDtW7kmjxNjN34s2OqFSBKjrhhkrKKLcthzYp29krNSAgeIfg+0P5jjT
zbRaN62i0KoTVYNbst36i05nr58T2yXK7FrXF5tfHiOqV4GDzke5upHychRZ84k8
tCwTMyplkujvKBYN+BbFzPASsPLk0V3UPtrTkQs/cy4JSFe1qXBc3oTWJHLrdfhT
cVDxyaWuaEBLL9/FgKDL+8Bl6q2cNyPp0HmGAU98qBZJBra0AF8c6UIiGlYmay7d
b8KHFYrPegl7mCrnI2fxqEn5nLMH8xS+qTyOd5ypyTi2Ptzhxbv+Mf/s8ldXS/+7
zF/aFLDnyHPFStz7O+PYWuNYuH/HnSad+T2HwIGjbMNmGxnr2o09uj/3+NIpn1JB
DyMcX6cEpGRDwu/MNe4QXTjOMYNoybl7bMqN5IJ+1O6FnNYW2nEmZu3L9FvWZoek
Zx7kZ3/0aIiI+zqNEaCfl/N9xfKVsCHtJmRDH9wLuSFhIgKDJLzuXsXAY0wyoXsA
uUFgcnkv9JqDl+JXb2C1MEzx8H4vLwBSNqFF50PEfsW/F8rKCCfo2y1jR1BoDqOg
Qz+LwEBl8D/z+D3BMxeh7DDErTQRLHhHpjExVgkvcScbZeP55xhztj52iJerwx0R
/9FbIbdLUIEuYs0ye6Jp09g0/CtMtWpGGFXy9bSztsUVp4qeJr1c2vBV7cw1NaSn
RvnNBa5nqhiPDGXG1u/dWGjadkiUYY4IxpO2qUAC1l4woamE4oMEdc5zuesIW7jj
L/4G5Lal6k9EE5ZDFmM9jqTaA5oWUiuFcGM9aC+RC5ra0Q9dHoqrU0fF/PcIjhSW
0nLKoDN67uS5thV8DeFp9PFmoveWVVXbS0bwI2ZpJnHS/VO9yU5f6sUtKDQrbefj
+NrGDIIB5APW3CG7qTPP2VAStarE+VFkOwbSDHOu6YsHTet/GNAqoJFWrR6jHK9B
dJXqAQswLvSyWbfX348eP7TrY+bH2ia7sjVZpMnQg0L14tT5Nfl+IfWFy3sttM4N
zYiryu9765wVmvgXXa92TyUhZCweNMfK3Kf2PQcwElPhQKWb9gbgE/Q2VyoIMz1g
bFsmFu/+SdA3yTSWOc1PNIEJvVazn4TKxzOJQgQovp7qCaLPZTITMireAsBpHlmg
nNdGgFQCA3hwFj9pYyAlK2q7UncF6LGm8QKMmtDh2M0kgVOF5e3AUqTf49yxLjjq
n6Z0wZYV+8lIr107IsWnoyf6GakyJC+uN6sG19oW5Lo1ReEd9nm151rYInbJv+sO
0QkoCh8iRPLOU25ZjeJtKcKVJ+eooz8H70G2VKzTdm81oEr66HFPYrEqoAbb1T49
w6Z43Aqrz5aLXIsrNq6dgk3MQFWXjImn5+VmydzWWEGY1dGo7ng2HKI+DEo29q79
e4rLB5CW4iXDj3ZfbTyY3jc9n0hXVUbEWmm7lUUrL9T9NT7zVeGZ4dfMtZgF1Kts
i+c+qj5ry3NmMMV33zJrdRxhlXmrZHqPADze2LTaSvJn/54Sal7W5CV4xAn+xqvZ
B7g8ueT5budxVSp4l35A4dUpWfpRYDfU8spUdczt8CwHCtFKPJMBpSoNVOXOMrEx
yFG2NprxuVD4a1nPqogaJv/gqfUKLxPOqsmLi93yxEsitJvqWU7fi9vXWO0z0f9Q
fjLS5fbH2HIYVSZLrsZj04Wg+1dz0Rr5r6oTJNMJhd5dQcVJy4nIJMpFpDv91dDj
NbyF6Gy3rZgR3etnpubHpsSrpFXJZOmICZUR+IAaUKpiLEqvKyAnPYKPOpdi1o5S
7JvVxDq7nbC41+BMQU0oqvodySf+9wS/g2p36DXAh/a+ucRGfxndfWruW1R5Xe8U
BTAbX5dda+1T3kTzN8QoaLGZM1ZssENf0v2vH0sdVI+wx8y2y/4iBPyXnU/mBhoh
38Y5DKIlQUUCoCZ2Ly7HIF3/VlTVqzhLfCeFA+yeAhoyuG1bu8cYImRGqWABzuCn
JpSfR4PcCXDebeXKhctOwAV2RpGVVkCwv8vzU/3jRpVHxlMYTtvAYbEPuCvt4PaL
9Ly7k7uWoHwbBvn76PuPRwk6HNVX8emEinPlY9UR5GuQlTbqwUHeB4IotrsRSEvg
Xo3RLnjUB50KQ5Sceskcz8nFbdJMbIz1kqhw6S4RFj7mjs7tB8ZeLzBSsqjWq3w1
7ZPxQPs5mRg5sVqMwY0Q317jF+Ze3J2JbOeBAmiARb0b/hszz8a4AOOE/jqT/0yX
NEzyOv+blzkc5Cod8LH7gQuodNJVEdVW8LG5K/gjdxkKZOWsXcQorNEMN9jjR+4Y
xwJ9IyZegE2I/0bx8BjCGqqVtKjFTM6B/Do2xlGiLbsJa5E8Cd8Gn/p+79Z5xTsy
ZHVN4I5T/C3uoKgQkKOL5iHAFYrlRv+r5zBMehYB1noQhI5KW9K0skw8X5Mq+D0a
08kb73Jb2x2J567H5yAKPR1gw9Gyog4K2zxruLCRwltENBFCkZeNSWUp2DTsEfFl
/kUwoSRIazb3eDShenzzkreCbD/w6rLlUOqkI+TVnmiH5ytw7ydqb/4sTQ2DYgYm
zOIQRCMOAZSRCiubA4ZcBYc38+HbwkDLYogVmws9cx6mwXkqctXSzAUPvgOZeRDU
nj0WylJfaTm4NdgKXJUYOWMgGLiWL7TQvmL+Pf6SbdAwt7OEdcA6I2xv8wDHY2+m
BfTeGtexssxuFV2myHFImWreKtvIIX7NOM+TSE5cyZnKVcTUDgoaWGlpo3A0yxE6
2yR5EvAgXBCqkKTTzO7WCEzRqZYVPyRIQnjHFOXvp36WiuiLqr1s1ZI2gh6Awq3c
r3L+83F334x0RuR3ACh6m1Vh45IitgkLNAZJ9KdP0xb5YZADv2jeTnHOPde6DRra
TKgA5xH+/O8+ki2XmFIyspFiSLybMLyNw1gW8lWc8Mq06Kw7amldgx/QC8g68cWe
9y4xz+YevcnwjbSnJ76pag8lvVqJIVp9m0YGbAQ/Zgdb/+78ouJBiU/E9pldtmaE
KrNyx8a4l+JFHMHH4LV4f/ekBYJvTticH8FFpWdYu9DAfTr0MYa86yTFVE9mv0kh
2IKe6E5SWZXxrVl982r/IHjcoydGWHv6fsoTgr3ccZX49uSV0kPXj0Y0ew8GwDck
IpjVjYfYMPVBo3Ede9SpIo3PjYn3fvhlRmiw9FyMNDmAddPYV4ukPdKFYouJLfuE
44EC0zcwPs4aF/pNk5kmMtJRD4Xfo4APXEPDMkMCuJ+aj8rGy2+hg8dXIYVlCQKD
0ryjHgCyaCcs9qBuwG78HUfHf3J1/JXpodnNPFz67M3sRJlOiNQMD6hpJyjHFd2G
zg2e0ycciwDKevAUyVdgoYoDw2CEApzhCNFzhY2tqqkb1NO7oMTKjihui8b3O1B1
anJBDNXsqSstVV7tnkhbaGjrIEN/QoOfeQxcMJ9qKz4bEAFAMw/UJ1UxN0jeFOvC
Z8GCr8A94WhqYuNlhN4hjD0ScIV4/BVnIAZtE7ACg/f9HFMKzdGCQL+0NfvpLQPq
YCVOULj3ygLsGyuT87yQTmpdHfuhByFSuqpOmb7FyIlWpb1YrOuP+v4hEZi7aX/x
+k8AKcAiMJcH6ysX3/VVUAKuJpurwQXarH4618vsuhv5ucPyw913PINiOuioFelC
oJT8PZmx8QF9+j8pIvUXi8ysywBtBo7GpyXSVeUqkvoPOrnI19tNpI1Bv7Xfmlzf
CGG1KAaYktLLO/ajDFqv6dXqOlHe4C2wpaC1M5DLLHRi7FJK+GvwWav8OhLQWdE4
VJznFfPKOAIEmjvbn75ZipCgbCBOhAIjeAJMv+9E1hsXLSfjQ7b0VTg5aO7ACZKF
P8OOKySWJg2Dkfdo/3IdEACEZLsizMh0CZuzlJBM5sh8tQ+bvo9tBQXoEqyHMRnq
PsxpMklCJlKeOO8b6HQwd+3ZlWUeK2/iOK+8plOqU8JGKt5Gbfbh/unLS9G0PUgi
MfsF3NB7XQ9r4zAMz0Z1fjfODHLaCgWw2xxQRTC1FjqgQVn58g5YZH9p3I5ElYQa
SKLRLvboVkPOjcmV3BvSaC6Sx8ky9dldZrtKs4axBsNQqA1io8dhzSDd+SpRvhkT
qR+0urpoZUnKOWx6MY833cLeZmlPuyabTJl0ALKSBzwi6s33/83EorYTHrSU8w+u
ao6SJL6MlUFXnTvAVRK6vE9ChCS0O8ljP3cS2qpE0Er0DBPd60z9A/N6yTFC5Ajg
WwEaFIvYohfvGOU4X9aNYuMOshJg+eUZafwDXbAQUVvoN47sNsEWNPEZKL2iBORw
vttMOhr02YWM+x/kWeGofGXoI0N70UD06gNNO51DuZ5C2306nPvlPyxFrhT8Q9/q
uh+6YxpEMN0P86A7wuMOU8x0ej0urFCmD/6ScCsAxabsATtwvgWxr2US+fOm2jm+
c0S2BIQhVkeNNpQVfxm8i0fSvAguqLOZ6uavGj+0Cm6nYx085edE6lvD+IObjQgw
jdm5c86lXgy7nAHQVFayai/Rl93dvnkzS070RPrIpQg63E36rRsM+jIQJqnRMluC
rzEFJEyh2tGbh/30r2gbl07q2B8gp8/HUNg6ji1+xCpmtreLL+MNSaYyH1AqfISm
oJAdaZj9FtqJJLcQOjawZ7T0ZahMoVJ5/28eW8JJlEvBx1Jdr6bJpVzK1a2Nhs28
wQrhev/ruf9273wE8hkfG+yG+bVT5LzB09itwRrL6PTV6lFeqz3YeLJm2SNX1dtO
E2g+Z80Iz/1usV73wJ8QMMpTphLGgL+UrV4+Eer1ozCrnejRIHBwC5vhCdRyDNcM
xHWXmBmRhFqpAaVQs+54zfR9054+qpNorR/xggJ95tWgQ4iniyN88dhHkJ+dbaLV
eVjn8G4tUw+8e4s1z0ASe6hxWYim63vzfcNehcAXyj4k7QWmZF3eNBsc+/iQ3DFF
pPHUmdHMfs6fHBjExKOov5DyZeT4fA+6cZRRE4y5xi7iTkLpgXy9QXK89oHjqbuc
PXM6M3ZbTQb09Q1ziv+n2QTMYwBZW4KSrQor1FCCUvod9GpZZfF0QOUxh/dpwVNo
nlfS1QrG0xI3RLzX2GHvIWws/RlMwOd98kVtLBczl9kMNYq2JNZbO9WNlRgO6+84
EbqrwCyIpEYUb8jfgdNp3zxesNvzfc93WQO9duMoT2JsRiSQvOA2Jqaq3JL2oi8Y
CdDz8QGCBASRhj3g+vzuQCYK+E9IhRiLIuUch2SFxmpiWSOKZZKQJEu8MQPGi3fs
2Fv8uBnWMw2q45hMsenj9xqIET/3Ejz57dj1o4uRFK350H88aYyfGp8PQJV+cWUE
d5cc35u/Lezv1mnG7cFxYEehNgISlusgA6gbbvaAtbiKv4MGYAuiXMecspl2Ochu
SKLHlDNx1siR8hkbaQPuNGjo9YSmzS4MBF/7tX6XoFEXW0YysJZ9dvnpvVbOOXWb
WEzt8ZdMkbdi2NhZs53xwiR7XEXbZfizcWmzYljeUb8AyGk0IgJZCKY03JtWUZQP
8iCf+7RmekloJ0PrXtn7tI6u3nwLKNwqx34t5vMu+8dwXDKTpd2+CuKCLn3OpUmb
gw+lbKqdVZduvYjsNeBZlDPN77T+ZEL2rAC+U4b3LDKYmYllm39Yo/BlqQwwIpFj
AwkXnsvuy9LmxF1+Cm2hRS7fNJ+4anU2XUqKVHMB8tEPqF0ovqDJpd0qej9sKqEr
s96JxU9ekNtvuhQ0BfsNpMVUXhUBBLTm3tXCbztlRIK9lSVMyQrXFzuZMnTSePJH
WXXvZISM1FLIrXcJ9YLEKX79W4/a/zBv0qn2CKPFgjqrjuq6Qgv6YeTSBOcmEFds
1tiOoYgn0Khw68pVg2A6c9mFbLuSc7Vdfe3k6Ync9h8VaWBBFxK6+DVNKi0+KWOC
qweiOCPnHiZk0qEf9IUjZjBxch8+Lf0GQ+aSNjJbOPvvSo/uAc/LiXZXIfqeFVVQ
ebxUd8gKFGGe/KqIzF1GzuVa546mF0LBNCAeZUJCxdcGQcN9A2b/61seHbdGFSde
bzMIdHCL++IxkaPKNdU3b/72SXS7IyP1NVgQiM9n8FkFEVrznYRKzwILMa6aVz/y
2Dszb8vpLj5YwTytUjX37BgWuIrqtxh9WH69w9UQcT7vGlbQrRZq3LrddY0mpV2c
eSsd24JzsYvRjL9J5RAuTnwr3RMt1jgcrJUziYMr0AXDfdWx6VM1mQu89Tfk0HHT
d2z5lhXqjCDiP7/lL5X5ivacKOfGGScidwsjzkpKKQ5zmS7NXaIvUUYNoRFtdq47
kEq4CGFekmapfSa3vuPRzVDTeFvEo/Z1B6BuGN0QAKPgSUKV+3JjjEFwl2aYnGTz
dwb/naw16opuIG5TeMfLz/MoHmKDWE/hV9xrB6tYUQClpTcaKe175j8FDs6ea+9g
ulWSjHk37Yv502ntaHpi4C3jgINnCgHBeKKbusTVk3svxjlXUjLdesoNAiBXz4uj
ZnZC91N9x3NcSbK45rqgGoh91T8EYZw104hwMJytH43ZLjC71jp1ZJcPuXQPjzHZ
RKsbtNSIg4HsCy4H2CU+6JXwjK9NXiuPFCAqhS/CRC4Yp58iYLD0b/tDNSk5UI7Q
PuvgYBKblzS5L35Ew7kJHIyzgVaYLC5KpCLyZ2AG+M/S21sM9ozI9DHSe7MOTUc0
XP7h+lKL6oadaPHE7evRh3dCDM+YSaip4xRJbj6A9k/ahUOVIo80aohlHFA18XM6
EAqMrfxc6HB287jxUJcWoP/FG1GmbxpvadiIQsxzvOE6oZ1kpEnWYXYoE6C0MjUn
tLu3/qRzTi/RIYKdu3eQ70TvYHQ+y78UpfqJcAZyo905qm1JNSGL4r870YomtBpU
YQ9Zm/zkek1+UmLNaFZkib1vH1RwVc+BBgS3ewuC/z8Sy15Y599ZyGxHxFjC3xdS
w3+41cCeuozzT34ekHvQ32TLQ5r2schqrWUCb0DkGUoIYpJZ+n6B9aHtbajGqnp9
0fsLoG3DhUW3+2TpjuZ1vzhfcWnRR219BbAE2iAtalAgHMWeC7kEWOKAFuyU1PUr
IKI7rNBShvrr56FoTq+DXQXQMUpun+xy5pQLztQ/Adl5duZBkbwoGv6mH6dT4NS6
aq3TRPSZpN8T3EVws8FoJhKDOiG24wSR0oW4D/lWcQV1hxqvsNfumu7TleZHfjHp
LpD5EMEtq/epNn69xo6/44cjDOIPFv1K3w8TDSdMi+gQrPaKqjai81RGN6wNbIbf
TzxDsZvxihbRgb3BjlsR5K/IX+IDateZ4rLyfUPQ6eVrxnnwUCnhc2XOnoZ/eOcs
AyFSMyE0HXDuFzp6cU5rXHwvNM+MoH2NCa/QJZOY9K3DsqIbwGTv4pQzayQS3da2
qgpgNMLLgry4kvNP0UgKDhuQsyUCjJQoOc6zSZhyE/axvMMaKkcgmNZXTtOaPgGG
/LMWhj4ZA0OzIYpIJ52CeCgV5o5QPAJOaUT0O8CTMeVc/Zt3WiWwCEkPn/tD9axj
O42k+NdNWBzbUBfJhXKkGDh9L966wqGllVhRvBDFB9aXfeVAtsJv1VXUS1ZN2WPa
GnXVjkH3SzkVBV7G6FVSsAujd5/L5skMV06Co5M/l4fZCYF0T6kOzJ56jB/4WMVt
aHkrwhhta70li96QHx4or9NNqq+qdQRv4knRul0UNxapCoM+RPZBH7OTAPzVWLfc
zAWZDKAIQbJ9aZ2Z/A2saDoS9pCTN1ZJewrc9pWi2w/K0ad2C9ST+5PGKuMIKxt+
Ez8AuK0FAiKPIKaowKkQDDW+fxUf+1mRP//SCcHO8M3toLbF4fiV31kNwdcmV4H7
lzamJZ20XkqJfVHh0H/vpyQ0779DZjHSuUgC4bMsit+L+XiiRm2lPR2PkFCy9ZHa
PhK8sv8ViaqbV6Lh8kYf8my5Wr4431fbDJrXZAWX40DoYfdl+9/vyVFoOIpzdd77
umwW/rH+udeezioOwpNJex2/y7H55nQkGPATtxIAOyWsP8kwN2+u+cKiEsgmLK2s
BAnM+Oy0ULNokVvnuLATp3mXMQLCK7Z0lwiFZo8d+6x13hGaGptBotnhBBPmpxkS
5pvPCTteUX2Gd6jvbc4buqvkmMJ3nKayrgkR7xSPosc7H3A6ZkE+SEDMhI/+9Oj8
LMiR7swsu4g64sLGZTggB3dJWtWWnb5bLfMBS1ZdKAHG2JPKU+Behcvh1q3QULOa
IG3aWQQ4eLRLPTlSvJBWcHN4iXYt1kOxVcXOCqORrAXSQaOfHHUStDNeEmIxHtky
WcRM3YpdX1Snpuz2p6tBebenCR+4+yGiZ8oddeCK1COpLDqzWU3sNroXvVglPdLc
Ez9fFXUhpz78yKPGX0MJk8rX6ef4Eu/ZcuOBG5wSGIuicWsCBwWUiT8uljpHcReo
QuTXyMndFd33VOJj74gIjv1Ce2cNSr6Qlm6n41KpN9HD0ZbYcPiKTzSRLdUusH5y
58aHXEmRMO2TSYE/KfZfpq4eoYmytm/THTgq5mUfW6D39FVNd2Z+JiHFAzoGjyUX
+IqAoj6whTMuBO/YaTyiN+auJ8O3oJ4v+ZFpN1KRjVu8iCU7gnLV6f0ADfGLJItC
lIyYXJsqOHu1CuzwRzFiFq5cismyPEpsIU4u16z3cO5c2U0oeqfYSVC/PYc7dBl6
Dg7zNFXoR9FukuXOwg6U0ljE/r3T39i3eAD715Tun+sbmhe1XgwpkNXzzmwUAiBN
oKjX01BLkpLS/pKYGII8Qfhs88MB+offNmhGZNYpwZ/9eqdXVkWTUiqpb/tdgUHx
AvAqki52bxwBpbtwS0LC9gk+NtLMFbwo+/LxvEWDJ/pmYQY3yfEuAnyE6wSAh2Zn
FfE9+vZbP9lZy03/VY9IOLRHrlIoXs++LNVGmTav1uv2KBdHtGGSwnucCMCyZPwp
Wvw9OHQFtFP5fGag6br4DAWJNISP0U536FZKdWX6OoDC/UcKLIPYLnUGBrrPL1X3
/vVtrfYk2qZL0JiT3CgLhkWdUHspKRkat/uJUe0c9ScPiArOHXwJzUsq5bdW5Sa6
RntmNldVYFhqim97OjdveBXkYcPMwfaNMe5297G0WKQE0TmSORGJYRMXD0ncGMLK
D67HePx5E+bBAbf/M40sSljxKf4UeW93xHkedQ1SMYtLv59Y0f9idkUodjTtyPB8
MeY7sZQ9EuDIHQz88GX+EGnzaHe49YBNAKrK4OMSHrAvH4EMkI677BvcuqPzwF0Z
lDWkR/6+IsFcM6ICrCUshkyV+PDiPYAiGadtve/nZwEFFhv2IyP5k6cmZxwWLva7
0t06hCkzGpAizVy8hv5xvQBfvaWujKd3SnEqxb4oWjo5TDCMyYxJjD+ajbeN5eXX
7W06BJD72FYQ6K8tUbixLq7ZRpmlFS22DRg4pXiTUpQBKaXmFBZZ2saxcWnwSAyz
jxkm39e8PCjjqgsKHOeeueF2csfWQCTj/AAvsRnCL3RpVJKI1nlM/KxrcL6O8Zag
GXkKgqfL8mABRXrltkQX9846n/An+XXGswwDCR7bHzJMjv2I7oUs217C1OXevHLJ
aoH9pv19hRpzQnfCwjp3NNFwRaxQws4esiWkrxQPOxlnhV4anoc6QMkMyrWupBcR
5o7nU9+tluNHMFEbk0e8O2YOg0mzKVQbt4dsiOEtGGQLGOSHJZuq7n1eC12AKfVY
LxoWNX94FK2Ws+9/w0XPbZtbY7wiSu59FiX11REEGP8uiSuIITINQWhX1YJayb1j
0/3YLFCCU6VLLf7Ey9hmcgZtdN+eI+HSwlBNg1HZh83DJT7ryqfvZerT+cZxOHka
Y6c+2Avu/GB2PG2FlytCeU3ZlbNyUKj6Mn5WykBlRr8qNuVOydpUqIoV1EdCF13b
Ft7wYRuXRMWnypDF+8sWgYcs9+1bol7Gqt2dykFhdTUZZOBhIVynY8jK6JKoxvWF
QcZRhw7xblgHXyVohEfjo6UsjuJGfQVuENiR7oJ4ZFe4nyqLTjgjnmi5PUsl4YGe
+2da/vv0InOgcfGJ5rS+/PNg+OS17Xb80ukIliyGTYMrqKJ4e1zjm3Sr4Nnq9B4h
0/axZbsnL95xCkz3o7OjSrv4MS926U92Fz0rhuTnfE1sobCEp7c7PyabtL//pFRY
W2JwLy3tq7nnVGUFH7gy+zwD2CKY8bvjohAGJxcE4+uML2JFr5yxVQHnbwbtvJbm
d0M3ClUUECL6bNJgGxe6KP8l/1jhlo/m0hQ+izwmNPbmUPChgb1trkE/S0jqsUIB
8Bryn+7lBZ+VoSn0aKIpJPNEphpdmVlluBy+uKwlDr42GGTjzQOfa6kM3/efdCYq
t+hxBhU/sLTaorr7gfBzPk6yqMfUrtRor+Bip+P5B1AEK1Roir/H/IFKDL9GW2Im
t39c437JhvlakemX9VFgxnwxvVrMoT5I0PVrnMyRh6yVRWK8nfwfUJXR/avIDt3d
M4DZur0A8WV8uxBvFXpQ1UbruWhpMBc1vpL3nHTSOvWfCOvapkXnXmrHPhstNzUm
c1Uxh61T2AVsa9Z6EFsGB/LvAC/3lWrPYxrF03nnSDCPSbyNL+DmW0LrB2ywhUjd
a7Atri4llHUQCN1FEnUp9Kdt9npWlGXbRmJRR4rCkUTpYSBAPlXFdqD6LwR9Mvk7
yhsZUNwcMC2mGAjdP1Hdl3TDN00nCY4b90exIAttt5j9n8TEj99M7geowJx/HaJb
Bwhow2Kjri8SylQRPsiDNW+Z4qcu3TZT7yRir3nhBIvbePxheSNiVcW3zQ0E30Bz
XVs3eL0AZvSVaYRUhYTjAAVmSXh9+WeJdAFYQCODwh+SP+JjBKmsgseGSyDSn4Fr
aksCZ4s3ldsj0IKZ+dq8uKXSTcA1o2bwIKb/AODNn/Rg3do2xFVJ1+IiMozP1v5B
CPGAQKd7jrL/mxq3uaEJlk5xLCZrVLd/hXMfX7Pllyqo7uXBtGkBZW3++yFRtBq0
O7a3GN6DJSr5m2jYSz1/h6x/rbdHyWWEOURABICcIeggNwYYUl8CDp2QGWUB/B7f
MB+jo3W7L7b/tfCCzYLP+40TvJOBGIzlDn9YSPhAtOS6BFQiglXY1K7ZD08T7+5J
NaRXS966/sC4QzQ/LP/mmFnR0hH/71Qj1wOjB6piON5t6XTl/t7AZo/zzJJ1kCMs
d2K3ffDo1wZzMSwYuS5xihSL5FZ/kMVlAf4/Gw9Z7Z9Zg4R+2WiVPsphCTgB7kLL
NELCDaImE0BiIYyMan0/ZxJ8LaGGSC1sEkgsIzJrCe/Ixs8iZH2sOrfDte9yFHhW
KfVzYTB9EmCbz2rqQxMfJC3RBish1uLx7G7SxA8VglkHu14VygDYBYbmHxR2w38K
yH0M7ftSNLgT1tPyVHcqphuTZw/HmV0s/9C6UayJByHcVAESOwngw2rEehp1gzoW
QyKuvA5l4cu9299U9ofTm4mRIKh45gQbMqlbhKR3+09GipUKAwJY3fatWJIdnlx1
ZlHOodWV0cTkWfgCaHR7Ddo/Y0oJVcIpIpHVOS8ssNO07W9CuQz24uKi+feXao3O
JpE0+MY/RQ0wW8iznRofnj/PbROToEZqYNVIuQcqvIj9iOM1NCviLifJArbF/isI
gGgvL7PuXj6UGrO42VOw95DMR1DKb7wmXV2tUlp4FH5w+2xqbFfQ6Hy0igLeQLlS
3IXKHT+quI8Px/sfLL2j97igKyB3++I7z9dVWr1e+zjc/IfM1BW7ssZMBazAvYMb
tBduVCWB5qwPT+tl0tjC4TjJ0+AzbfNVoMxwU0vsl/yRbJ9aFi9pVGILc2LTvRZi
JkYIqKv1e0ZwNUmxi+WAs9bmmuh2BwFGu2VEMdhYmXtr+93N1uH++U1asR4j8izw
P+3Kzz31n8LLJEwQ0fheOyZV0Ms2SSuvUkAHFU7GR2450AaC3chPt0Gj1iRpzaoE
74kgh/pIGb+8g2zhdtXsJIxBDIIFA7DeWz5UjJ44D5ziChixRqIexIsrwoh1oWoe
AH63LuODrIuLgp/Mq6fKatwDT4rimUk4je+NxoVjMNXt6x4FQ8KpvxWyHGXzo9ub
ntvSVFNylo+TM08JWPjY5UBbfVuiT/IgQ0juHNAdz8FmLGw+R60BomKc8z2/V85h
wmGtDh6SYmMen24SwCvtyY/gpZRNI8/hLUgUQKHAvOr4PFu72IBqAoik4IIritmG
6Bi3nZN1PWS6tgisIz2/tqsn/cZPKW5C07SkeXp/Ul7HI7vjqdVjZOQHbZGXHF3O
5DiDdZp+BZbIitUWoM5htgGNeQCC/P+sjIhYQNb9tIq+QglE9Ep3ZptRMpc4N+gc
HU5tYy1bS0uYyPJImw0EFpprjHEF1XJ2b0SlGLsfaznrewFns+6u+nTWG7QyDO1D
gqGsIsUDsxQei4LkDvBvkqDCU+Th9CeGX8Y9yMsWvMwCAALL8FkF2Vy10P9TIAuu
Ms245QTcQ5Z2c7tFqX6torrIb+Wn/N0JJTRvLWdgicwxxhMyPfxeo/HO+I1F56y3
wbhXj6PkafHepqXIYZBorhPCqD8ZM9JtKBJaWGXbheIa79sn89D52zayy8rJowKW
lBEN58bSjvpLrVKlBWiJD4pbR/6y1RAGUjU58SI0vkuxO2qR9aO9Js6Q0jqwKKSo
ZgTGd1LeoNZ62xlgMbR0hDYdd+04RsodkBQmNSjRhjNgSEvrZJpMr0VDqOOhf1bO
V3DoNmnkXvjv4zbuOmlYSzSDqXatht3KUdMavllYPFj6yXF97loE/GflvTHNhqdT
hBvVeOQjNuI4t1LCWtLR9uNPK+6Wfgm11MgYxiGyaevvIxUOOngVNz4d1USdiFxM
IARzLY8RagJK3CG/6f13XTP7Ab0Gjf3X6syHf2pot5+JT7qZoaTiLQW2x/fusWnh
GRrElN+w5o25uYWE4MzUw5IvF/3eRlMMlL9nzTyYn/yZJ9shIU+s94FiyBfk/ReY
4VwxrkpsQL5pQLZZwTT34WXWvXxDjsxL49oUzrg6TPykXcpLf0RjAvD2RiFFWiJ9
SvrG+lNxKGUNPPx2i4M7Q6uyMcACad1W5y9CDwjuTmKfKJ88KWPIopSZccnRWoxa
VqKWQPPmavS19lEzg1ieLtsWnDf4KLI6RrwlvQlPr4gB32bHdEYGamrPUpBzQHG6
zB5GglEC1H61OT2fyftPHPNfiMj4DJBlrOa+m1/JwdQBOhkC5rJyK3p2Q5H+5e5c
xOUrYj9KZbo8NaVpNxZG1VoqcMk9FX8XHhz4GOs+woV9riiCITv34x03/uJPvyHg
CiPW5NxyY6R9Bj9f7tOmpCg7QFqM7dVLiuCLS5MYiOtrwP6i/DLAM6DxRYVbo5EX
8p8XCz2ZTLeKryi0b1b7LmI1VoUNiocmseApvoPn+6SmP5/CVfPvpYeeidYu0mXM
aimZD8fUTXXP9LUx2sUi7UdaRo2nw2XLv3Abgng4T+K67AQiliTbzvBZn+gdZ6wo
oWQg8EniCThWKenn/JeJe43m5b0ldpuFBj0syPCbCEvvjVAThrthW55LuSwEvk+V
++gzoNQQ0aaZvP65byqPLcOqLpK3L0Z77KrFn6LPohH0P4nj7x8stMMl1zzJ6a/U
ekLkF+H2nHBrEbynOPrfbVecvxf0k1ArxOGVmnTnf+0nRQAC1iwNrXp/xSPXhM1O
+snL5WO/1SPzlAuVvKbOMdKbO0eLuDobgd7oK+SV/f+QqSK/mt7VGuWKxO4zKLsx
4JGnQ8JSz6y4d2c+Cs6W24/yoBZFVcu7eb9Fai88inepc77rhJ5E5s3xta8y55mc
o/iE6M1OFIybzmdWiXM2lGYXVXFPq34q2w4puJ3Ho7ZI9PQQtHOwieqWqYhN/BRn
v2vDvwWjXyKgU1CsyMxgA4ncc7BlG5cQzdzVxRYTBO+iQHaNQt9LSt9+KIHy0Tma
B9nS9w1l6hsNz8u+Wd/GySfuK9K/KylpNI0yf/T2fIBkuKI+3lA8NlcI6Wb3+hmy
lzgiqgnozOywUdR6LJtI0gJA4Y5zhzXvpU3k9LqsUD+d4QGdrsO89B3DFYXbiBkn
qHuhwirnX8PrbfxcJcNQZcBx69WXVcslsUY/BEEbmNQXOL8JL5Ld0akDa5+aPbG9
FUxPUM0n38uT2KlLUS9ngoowLwrysgJ1pI4l86hyawN3MObIJIJ31Rc+FKQYC67B
44kbpyruI6EwOqB54ib4QyEz07pmJcmBsNNYaJ9PdPVOdBgxz6v2lA0kKiQQZkDx
ICuwx3bsjbSgqEBG1koyosVxbugZzPveo33Gpd+itwftm/EPaKT9bdgzJ+ibA51+
nKmwl+hYjoSxKfCoKqfaNdLzKYCC/XCyU1bFzRQ1b8dCVQVv2aQYyRw1qsKqyf84
ETOCNb9lnbAj0ej4XsbKYcfFE4qwnqqpiR3JO4oqdiKpk2kSj9jTi88pUQ1ivLRz
53YGIERwUb46lExM+UuAswzJdq/31f3+ho9Yj29pKyEdjMEn1I4L1PPqynw0XwDo
ZhwiBrWyfoVy1q9yhdeIBfodAr+FaGsQScISohvC10aulYDhId06d4IskPYCHw/t
VBFu6eoDHYWYzfUtqmJviD0n7DiWsODg+RXYqRdrErHshmyerYa3NbB6BDgAyCRC
8o71l3NylJBt9TWUvffexyzZV3kjAw6bgBQO1AAG0QPpzT87qHv0cIp6nPrUCzPU
LvxPVnA+RDDUaye1McLOOlLYnpoksrv2jRP7hRjPwRXQ/YSi30cfuwaw+vHe7+uB
+E+UphF5Zd8Ssdu3Hn/idcklzY6Y4ECDz7v1X8EKxBdr35CNtRM2wQgnAPzjSMxH
Aac6ZTFrwhJKCg/l7me2sMDC733a3MB5GKSXHYxyfXI1ckxRgMyTNkclCoeY0uy5
GJeLffNdNrr6NK2V9+U3ml686ILFd8bDLqHfC+0lOJ95y7PYIUjr63PVfpt2ghRw
7Y/hJLvuj10D8DyYqMqgooNLwvSDqCS/CXW1FELVtZ2WaGO6WwHZHB1i1x0wc8bo
j+7dTtyjd8neodsd1US9uWL/BKkDS5lmEuS523Sa5/TfHYlPLiABqFX6Vdjq//7r
kFhhRRO5BSVGrz0Scj7GkljmzQvasioxDnnmJ6KbwFvJ9VEb9VRlNG/E6ovjYLE/
A2d0qJsrUYd/aDTk6Ovk4tbKSTqMcWZ1+K6Ql2Kp8NumVOMwwm7oM0ma4dI/hYz2
k7keNPlCdvBC9L5eSzHC9xOCtJ5D2/Ek/fValE4O5e+3l5GWGCfvRRHdjf0KnANG
dLnek4K3j61Ac1KzGbOBd7VT8WXUSPXqpHc7ARvAwylurmzQ6gy5ozJJ4ynS5vxU
JmxFY/w+dquAUoVJNvjBSidd9ZqSpFeW4O7yfNE+Il+yjAtXfqr90ZGHUozMdeZ0
skUAHG2Xvji7Z+a+6kTfcp+XSGoKaFmn30LHrVyuFl+eLGb09QAl+qPcOPZh3P88
F2R7kPvIDKYpc8CRd4W6YRXEUilj4MCTMEech56DQlUw/O+v4vRBuxoOQTitYwUf
yAYGQFZfRdEHA776ZgKyifQodRtaX/SBYCvUvXDzGKubduyRwT2IeolICisBn8yr
OfuMiDwPuqCeJ7JIk2hnUf2DrHon4E0FIsxuP3uKOmleMGdC9F1SvuhYfOEWg9qi
pss6PHiGp4NO/dfGbrw4PZDU0WqXU6CzQvvkOjzYNzjP50vvYosJxiCS5CEq+bJ5
KZnYCxeQSzmFmzDL2KttkxuDlnclvdMz1QMGC1PcazybZLwtGboTeDrCbe7dgI5A
/lhsxO0LjONnwicBN/ptVA/kSds9vLaiOqAr2tGQ6tqTe14YFZRu0VsWrZgOPpni
p3kMbKpX4x9g1NXyHCB9Bg11Y/2oij23JOsFdC/ZVoqG8JUjJtzcWtV5/fZjmGaR
0d2Ewro6afotM8xehl7dj+qZ+i1ehZw/2AwzWLWnj4mi6zl6vw2H6U36QrcBC3XB
/UuX2OqZsCmQAcpy298rBs/9lJJREdtVmLTXqNLVP5Ad5Qv9EO6gemREH4HfWz6U
tYIB4eDE+mFAHGDhsO7TUqcfu+2IOHUAs2NkWR0Cac/xB8jHKPDlss6P6ooxbZ9u
oqqeCPf9Q6eR5QDzFUODm7NuyvpF7YZ/uPKJ/ao75eEgqY5wJZWRrI8gBSaiBVjs
g5lRUvLhbN6lkQh63idV5BTdqrZQmhMPhoCyFVU6NOidR9IsrefSrFGiUZdlHpH+
uRLBeDtihROeAtThLrNz4ElWvfDsquhHXaU2LWwbGht9Ph2abjNJONbRYSdaI4a9
lxpFCyhGBp67VOWkeTwdHDUaOdDUa0cFLY7uFlvfDeqsUGPqC0c9NyoUtr7Vvnbc
frSUl9q1Jrtd6FMzpY2YBmLS13PRF7XhhPl2tenDBTCd5amNtejmDFBL8jv61mu9
kyPYBNzn7Fxpq9omIRaqsBFxrD57wXJGKEjRkeeZeUGsMc7ZNwJDydaE7ILdbtDn
rARv4sfOknvNVhzzunikjIXuQXgzmfC7ZwcD5LSPzh1TLNDQUs7IkvfGSNk9enmL
kdC28PwB9sDiP07kT4EMdxZZOhYDdKTKO0lmU8gyF+aN5zJnmB80Mr25INSFHpGN
v3Yktlvmje9NVWG+wWQty7uKOzT57V4dSFHqcZOWXJbz+uhv9d9EiS6u06PUG9Ha
tDhlaxQe1tFakOSd8FRPLNbx5zBsOBzxJyYr2Rr2ZYlRy+GFmrFO2gKoV6wQ8ZqB
GDgzyJ7JGMFpVXOdgtn6DTPPAWfdDZj0ZwpVZ8I9b9JndyuQPzhDnFj5iVfoCjtP
IdvRlTvfLYj4fbjjMmF2aPtQjbbYWbjlMLHAol1aeJxQiOKBnmr6wZtbrUCVkXc4
YLO7s3gjZX860pqlhai4NF01ADit3m2Ww9huI2KNU5R9FKp8a83FY09lk7N0rbrS
G2psM9KyWKGAqMbL47reLKMYUHXW6hf3uKM8eiGjZqh1EddqQx43XgRX+iImXK4L
MN1vdL9VOZNIVg4Cu+goAAVFx4mGJYIaihm5fk4L7vHOn0MLm/tVKvBqOWulKBn5
vTk7sTOpG764ATlubvYh8TL1CNIeFCIQHHCbn4u46ecrkr8SYHtQ6bT2CUh1UX1N
uRfToaE8wLUrHWwpHuB6DCsi7gD9vjiEzKxfQrFUMBJMr4NLKcjUaDVJqKVVG6Fl
ZowzlssxGh57KeVBwvVJ0IXECK1cYgBl56F2EmvzSqwJIzqH/tlqtzQCHZSOMlxs
3GS90VWgamj4POPTjSBmp7ok+vxKA6lX2EyiWI+4bemnZzBxqUaiXXLHC/g/y8pR
nYRW0OKwMWXENLK+IXweVhV1kqf57R7T5Mew+I1aWEz8Os/0/fFWfwMAI0uMyLSC
0a46PCWWKKTb9D0zn5Uw6dKndx6Qy2BmJ9AldKL77tqemzX5BIjFl7YIwUqk4LRf
+g7e8LMYBBf0zFdG1Q5RKQiFkDHLoNLRR40RBQcscLH3ZMGD/IFWsr7QmKownwIs
/WikxrPIcTx3U+6idcfh8iQQYJqfH7TC0foAw5/dIbdXAKQdsun41vYcv86+KWP3
6surmDQ/PMSyinVt12hSoD5wEk39EiNgMuRE96HlOGuzsGtTpWdcBUJQj0Cb3q6H
IbNGdWAhy7Txg3JtHvHZl+uwxGRmUWKWFagQ9zny0d7P60zt59spNfPMBrLPj1Np
i+c6xZIqBarb5rg7+/VDGG+nCMNWTDx268faTyAJnV9Rvq3zzx+JxZjD+cAfoU9B
I9ecwVKUsMWmMR2LCbuysixGEWpqnPi0YLGiO7BlfAThGriqNv5aOJsbvVjlz/2Q
VIAuBVcjOyIThKnWJZrX/k5pvdkHNyR7tRn3pxQeV2d9KJ+mpcareGrCKlP5G1xK
Y3LdC4Yq3PB05syUX8eQDWArJ+7T24SSwQDrVOREj26QJV5wlJlvQqvBQWNAtF68
1oKz9NSuqgcuFIg7OYVg9GMpkYQq0KfAlfvkGU256gJhbC2letm8sEQ7pghMvk03
1hB4C/Q/2Z9FryQTLDAc5+ww35r7iXBvFWacMtlqz+Xwd9RWHfMn5Fvkoo6IoU/J
VMV6WFaB5WusBAuiZwVcbM4y0sIKrrJ5+QruG6fJqJpOIlLSGNjZiFReEuIncTMi
WnBJhEcRoMOZA9nu1ofxFzJeOJBaFwgdat5BXJQZfCWHqkTdjGGGttrdEwlL1AZ/
ZrZTAxdPvIjjFZ4AAwDqqk1Z5CdnCGBHAQs1SM0tyMJffqRLHjvIO6lAWaTa4EqT
GtLwYGmzTeAmpgJGD+0JxbSC+VLYVqiFVzOYMal73b55hpZn2gkkx1NSSFGNUPc1
BpK9BKDsI84qq092cxkQP1bmjzxah1vTvhTQEfEk/etv/NvGRJis9QLv/BUik4Pf
nR+hs6DNAb3wbWweWNU67j3CWANlW9erEpkdg7s3RrYkyfSoLEpFr2arfjXozd7S
FGRt/fnA2FW0dbXQxXTI4OwjNaZwTsZGre1HsatU8RIgUXF0WFLVEy9yTw1rgXJm
BeRguXCG8Vdi9dPtfqQo2K7dgEKkNgZ9ArVwZeAsvSSZB+MkUjNpjyHegdvP26YV
p46HFDOfOsNdmlUueNCe3Jk+D3wRSnHp/22LzorvCZ54Cf5QFn2N6+ZNpteTDTXM
yXmQC0Iy5nG8/YVqXhz4uQQIz6lV7j+QQcS9YpPCyP6qyxJ6rJ+q3py/rzUbOwrv
FS9kbcPUalf7Czm9Q7mppqTl5NVsqw/i+eBKHfSnf2HkiYnog+ozqaB3skzqNDYA
L2M3GKwOfURba+eEM1lneMxjrWQFzayG8kkDt29ys7MykQm3bBxmcyBixndcSTS6
6U9T5lLRrwNO1EqyK50QicLBF3b+NT7qFzakNF8dbUy2xklskjN8D94A7+FpdKDg
Kz5XsvYlSg8JmsUXP2gJu9nvG1DuJIapWQd/mX3nNsuMd2tu/IIne6bBVJyqU1iF
wWF9Lh3eiC1D1ZvJYvFWojCFQZQOcT1Kyv59/dNIxuz0zM6sBvBcxukGeiMwc5aD
L7eux2gcAI/GRzsFtkWlpUTyVfHJld1C4SoAbrugnII5UdRXND6J90e/S/D9Na9g
fDCDhL11c8WsXsfLbHjfR60TQux4WvNpgSFDRm+tF/4zUsb7LXtsTdNHC3xPii36
QpuuR63qGndZvePCBu1SzqcVk2fMJW9uXI2GqDHxcZlrP4X93an9nexJulpwSPw5
dRm32xF3U/QwxUp8QneQ3/8rp77w+PCBOH0i0F0Pn2gcObIa19k9W08tvNZSW/66
uT4wSrmmbFaUaNp9xllCa/SWqbi9UDMK5gm6TvTzWb8e0nqCUnmuV1gbDBdl2cef
qcLlEcYdV6HylTOtG4dhoFkSStWQlUPfKSiiSV2elIsUFqg8XL7slOU3teIfKpi7
kTJsgzfyX8EXRkLr1XRlqa/5g/HDnvWKf+1oNeVk0Hsnx2d2YYTMS949g+y6ZMym
CsCf1I23eMzptDY9B24eM/RkdsjKciIkzCk8ZzYzzxzW78T/WnUN2lUF0p1SHh2o
FMPtb8wplTEMU7PLkp+7MBM11TxurL8lJRpbPBrLcVIPFCNOuYuSbnnIkhlDx3TX
/7JmLa/j6m2dpKXKhV1dQekSV/y2py3lPz7GOQk3nTTffjKaP4uTas2GDJaWt7JD
x/kOaAtpBnpFWYRCLbciawVVGj43G0D7IwA4Gf6Vzg6bPF5ap9jyFqTqIn4qU5Ez
iSCHrmmX8Q+SmyB0NlWluno14RItq7pw2NLvYI6UEvzFMYH6TDtE/imj1bYgCmpt
xumpcYzyx3ZKmq1Eb2KeXOtOr/i+3Zwfka6LQVgKWYi6l/UZcUstgd7Z38IKzYsj
VZ2TtTUqeM67HFBeNEY6by++lBNOOgy84hTos1VtwuGrJRSB8RJKhZKMDPYBbZNp
hZpeo5tbl6g0CEZ8BF7BYhTq1kzgA4euWZkiCg7q0YPGcjIqKBMsadg7gsktD+3J
RkXv3n1m1EMLiHM+67sPOsV8wr4huDFseidJkddU7Gij9DUYUAA2Zp9yDzoO1dMF
4I77yskPsetC0qFHRRdPW3WycfphjSiMRQGTu7Lc7YAfU83/TdJXRX+cOPHQ4j15
5HlovDD+5F0MxZX3MC3Y3xLqMha73eMHx2BSA0VMf6OrspxzMtuMLn21JlRYWNtk
ur2+okmhgtImzzHlp0n38i5xQ4A272XxBWuMtl5EB4dh6j4m5j5dz0WjJUcy5ESz
lBihkAVyjaTR91heT7MbrkiPayp8b+WPvRuoVyU6BxdpAR29BqAJ54/3BufSEpnH
oNSCva3nxxo8tTMJXfSisfwLeFFUEC3e8t6h0JxP+TPteZ64X2BJlV1D/8EnOsZj
yqt8PejLMtC6X6bIsmjfJM7ib7dp/hr9RwE8uQ7pzacg9hlg/BiEwhHj+KfHCKk+
OlbTVOeSwYUwBT/fDONCTufoMny0swRALpOsPnzCeztnKxjQe7T1xpnQgk98p9TY
EkNdzrMYdo3vHESzEnRMlIDEAZ9S+z52GJB9/hqtmLqTvsiqQanNWhe7ymPxZhk6
uKf72SX4PkWXhnLEDTdy+wsTdgaQiizk7c/hY52H67ewAtDVA/JkeBG0MGiHe14p
21sufxB9jo57w/WMeRTb1eDnsU5HRaCxY8vPZ8ovHuMvF+w0YtuvF5e7evcxn0ZC
+EvreyVu3pIOeEbW9jaUGY/V1KAonOCy0eRP6LNVyMoHERDTSaB5U2Q5EQEW+zKT
g+mi/+6lpBqBCjyKfJw49yufr8MNJuD6KEVZFIyMvLFg8HSskSLc72nM9TgMbPTn
3kHryEqPiWCdaWlWYwdBjNPK9V7Ddo9iC7Rpbo8OX+I6F0jsNNCSe1QJ+sduSIhe
WH3y2ZT25UPzq03YGF2D7ls797BCq/8sK/593cOprpDyTPRCrbUnjgZePutCBQ/W
4yRRJ3NkigREHBS128LrlQDEzg1aSjHJ1ISS6YFHWsisQaqcGgHHUoAffe2pVZV+
3TqTbt1bcutF4wmlEI0fk8CGQu0eTvYrB8k1GrtENdR92G4KzWx6RgxwTeadAKL8
v+3fiz/mz5izNaMfQF9mqkdmw3UeralM2zP6QqoVRAtVOJO5hKanVOlLeYSCQiMa
sA40q/vtpPgmfGblF9LRgwDfCqiwF6Z2zfvgSx9ZrwTBC7f7vGswfG+ETTh9t/zc
U1CL8NPiFEhIAYOKKaSqPc/9t05C44+AS7DqusPq/BSjd44qrfAzsOn11+m+XNgM
2w10JmGAJjcHyJS5/GwAohXAiHXzT6BbqRgZQJYsGbv8XNG7F3ForFmQtL3IH+Hg
spfrUyfu26HbvOWBw13WT0z/2ItfjB/wzZK0Uxm2eCG9Z8gq3gltYVcStkRzUmBE
9X6S4UDGmUOPkg/d0ZibiA5y8S5fHfcp2P2cJiKTcJYN2D5MwUYP8Tx7qFWIQQ9g
zdg3XHVKzNPJEeJJNVXXwIgCiA6nleocSxkVcucG3EmcVKVlLYn2otbW6sI9mccQ
TEkQuaGeHDxeHsfNwES7GaToK7HL4K4lTBJ1hHueIhw2xqkeeF/hYLuXyxpubgD3
UXlK3IylEyksFoX9NCWHAinO678MvDtW+uNy2BUWCCjd8BHWPTEciYhyABtstzLQ
b3W0ARwiVWbug4RmToMP5QpUt2fSgSuUxmYmjytD41deNVpcrb14hBYa6iIKwK6o
K5BkxERZQLhEkKPR8+6Ro+zgwNnhzm//kRHEWOGiytQ+EkAWTOQH1+r1im3Gr7Ml
QLe85gPTptll31O+1+hvvg6r+SXcyLoYZn2u+DtVZcbzRIlOOqyw4Q0YwSNvH/Ts
zWwA7KxihJNKVHWS68p2nUgAAdIAqXVve3Wujo70w4ce8wmx7bQj5pKTJVZ4bC4d
4HNhiXRjbVAYQfYdj2Q95r73uif0FhtbbFwN/OF+lRJREH4/lfp9NNjgs6bUlFnC
/O13dH/aDF0s58S1tXv39feChAg1hL9NoLQoBOM+mhBnD04qb06ARlNFsdOasM8g
ZmBi070AxJlUbQxD8utoKXhzU/DBFtbp9ppbByLaQ6KQaXeTEXrwa2VAieRl+Jio
luou1wKf2jiw1KbIToAD95266uQhTzSjVWUk3iJ30H5EFz7KZhz9HnCJ+iPZBTEH
p1qF6GC1ssScPItAFVBlxWnUyE83IsAQznPEAjzfgtTCLbXX+QcUh7/yShLyl2yc
0QZf7+2NCWgaBmiBHK1U7KRM283z7d9eutsnQJVpo5XKG65jwlemUhi7L1cbm5gD
Mod9oz3xZC26iZnQLkqTCrHh5z9efEksCbY/OXDyhoFNSsFCVNhHCrvstnEjP7y8
o+KYBNptq5MrYLf335I/UbQlzna5VWIVkfRqQjaeFCc1V2SGVsANJd8Uf+efa/rD
qklaMzPJhDJGDpxARbq5L03AWhAARYX3OROMWynkTZxYyFezPkEBFCo2LArm4OuW
E9efuAAxoruOhB5kT4qh/LnAaweGZGHjktK4vy4Nn06Jkg+KNjK78rfi7YsCdBUk
q3Tu2daLLiK2nRF5MLhVqF4lmTCtW4NmD0/VD2UDx6cfRX2Rn/idJh2/k4Vy1klu
+NLJ6yfR3HJwamR/6ZBpPvKUFtM21lfG8p31p548879IbgSxdCPho+cQil6GV9QQ
sHZDUoHoJp8OJpiL5KZTpL+VvM4bsU0GrfOBxIRywXuhSFWecPP5d0kYJmEHgTH7
yMwxMKUfei4OXzTodyRf++C1Euf5okWetYVgXozLKk5lbWpLZynT0gAhiZBqC2uN
mOADVvNzsFqLOx8x0RUBf2iLdGkcz/OrrqXNjgNJhj250R4JwL8XbTuiz1np81eD
ssxQFIRdMbFOGspWHFkP5+5mlkKwLshNAYlhxdAkCkHOk8jrP0ym0G1Zb+8N8Me6
9XZSdpVRGXYsLDIJHas4IGgYQnLaV5UWBIMoOWnKu6JsgrvCN60qe6assDL4gPyq
iEjjGQYcde15loqZqeI3bt4O/a+ZdVgdyzH/0aoOHxCJrwrw9kysOn/F7mISJsxW
KEAHT9IJgZvBRmhTtBaUDkc2HtfFt/0yxVmW30GTk4NkVSRpkgLcXC21Rdh+lfTL
Cc2U5sLti9I9ST7PA3NO7L21Q+nJC7IudAU06tpM+PvS8CTdtvnBGnZi1gKO/8u/
WSQA3AjiIJA2XZCA7iPtMTWNLsFREVAVvJRAiPCikZf+IuEk0qXt4SyRvhmDEw2C
3HczYc3wxskiD7YTs0acZ9zGqwsz4qV3I7ZGJ4GbI1pF99hoC2PjPBQKQpzNRV91
ubBTzz9EE97AsKChy+2lcH/1AKthqwsuQWDtPMD+Q9fPHZKpLq2V3PUeu3NBXplL
ox9cuymZV6m7hkl9tXKu/LD7IlHQwPqvQ7b5EXR13EgeFbxpuD5Jab4Rw3pfOqms
v6hNPwogWEasV+pNKecTwNz7kA7LHraaCi4vph1QZjTEam6oGF1bsvcnjCmJaF86
dCTN429vnmI8Wofgql2AnDb3gSv99JLrRPn04s9V1ZW72d2PyjAt2ONRE+emqbot
8WiwsQ5SP61b14jDPlAnZQVIWPZRkgK9FUqBuIb/waya3csHjmNC1QbRZ17VDFoJ
ZgGvAJxleAUKHMucK396iSgv+YRMvIWXFXyZF7eIf7LpUt8b1f6f7iyWHzTfe4xa
T+cG9YvybMjoKQ4bLn41Vka0TrGPYRL4PhUZdnc/O66ZR7o/XsEDrrUNHNsmdf1D
KYxDTGj9QlxcSnMZZ1TmEA==
`protect END_PROTECTED
