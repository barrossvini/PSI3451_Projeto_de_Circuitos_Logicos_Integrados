`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CWPQORBWQ3T06zPfgq5VLvM64UQwEm/lnmPST1ubURUtOYGCaGSIKiNndwZgS8c8
S9AvxhAHPgh122jao6f7578NXswUMzRgIHOICQa/J/xzU/2cMUL52LjKs7a6SSAE
cd3KVsbuZ3yNIn7TalobSgWavUj0GYfrMSgwhBLBdx1B6Ghl1OKz6LjvGI3Oxm/i
u8ErJliErI8ecl9aKM4QdFFPmSthUjNs6Nv0LNPvzU9lVhOPn+2HR2OLPGwdskba
EWe/sFgPlQfxERl0wRPRSB+w0mzX48XCz9uUbaioHnIIp0ox3jQcCiU0asFv77/3
cfI9g9Hw69Fv8jyedfytFAE3iVGexCw8m0LbQ9mUAd5Erc2A2pj9cUOirkwgNabc
Tp/WdkPP8KNauHXgwBMZrfZHyy6pmwf8Rz+xcafJTzWhXUcv03m9FEEnenX65JoI
8ux8Fbsr/and7Gh/kgBkdsLtwqyiw6CR4o5kAMpELmT8GNNadGy5TB8SIAzsAR4O
A64xBEwB7D2bpgvSMXDXgyQo6jRcI02YbN4xfXOhkmTplkx2VBzFXx4LBZ+YU6qr
How/OkXKFImBTxoIh7IqKDkfmoTWCK9QZZkLKz7WgLerw8yLBfuA2dsvJdFY5vtn
Oo5ZkMQwiovUBJu4YmnxkeKhJuXm4L1EHKt6oELnz8R9LplLD0QlGRiUUqYvXZ2j
kGYTQpYx/ikFGfBHO5qHGZYmiWUOFCSpdur/mN+60HJIvuvtdW/i3OoIAtO3sSD4
XPTde4MhZ6KDTQEd7Ko9rcKect8AJUOSAwi9fToD5ZoOB9UlMH2rWvFJBl1BBEnm
PZ+jkT7Re+aRw9guUlFwd/Lh9uG+GFAFJmJvEfsXxxpp+6Z2vx2ANDPpuBmXEYfB
lT+y2IHdZJ+T31/LFOt97kevUGLmNl4zfjSwzLuXCL4LAkS/RPgknkJe1eXGCZo2
kMa9Bz6Mc5oM3FYkVnt6J8GmNG9w5p4DxYDHMFrFxw34NXTbLLb0ONrUjUJb3N/I
LkEseJvwqk6heU9xevOIjxRO0DIxrKkydSt3jEOE1hOTrOrd11jMAclUB2beoklg
X9tFnwIoUU574WyWWsAvg3lQCECSsZkx0wASRL7tKX8cl9M3HHjKNWL6BevyP8vT
8UO4mRTn+ehV23qNfqy99WYdW/6w9DbsxyxHQZ3GoFPHTk0ssV+KLTePBd6UhZpk
50ovlF+Ygxn0fYCxrPNZXYonLQnx0p3fUBPXdwzd0Bl46Ra8/cgwukmmkqx76fEB
dMi1pnPeNx2/+Q2hhEFkEszVj8G69uD+OO51stvWz61dlM1EszEk1ShldMjVewGz
ZO7WbzsTvj7+B5PG3lET8umjb/YaaYwoyNDvdA7MFmfem0L2KtkiJosQxq2C0Eee
xrie4GOd4P0X4lxEX/uV1Q==
`protect END_PROTECTED
