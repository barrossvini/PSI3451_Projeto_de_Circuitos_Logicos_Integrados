`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Fsvz2GOJtkm2yLAZaLG0M4MWzZrMT9botzuX5aLZADkzxV7hu+pHxAkcO0r6W9u
Z4eyXi91KYOze+5DCDcRfJIf4HURf5tuIP6X7LxFxzB135mVbiLG5VEelMNn/nPp
bw6J6d7Glrg07Otv29g3tmayYx184t+yjYxWDahY1q0lyEg0zgXN5/avQgDBc6vR
el35FLW2AzMhtxNhINeZgHQ+HFVhpCj4lA3FLM+MyheFyuG1h6A7zyrhlMIVLb/V
FgL8PHKTTdYirMLwVAFbIPJm2pkv5SA1r3g/tAU9OYpfUgOFF+SFY9utvXBpiweT
W7YvqJovldKQ+o0pAeZaviRMJbyEv5HBeKf85dxNkkVxGi0O0PppcvwL4Jeqau6f
MWgPh4E7ov7rnM3znwYa+XmU1CnI9+4lSal8tD+B/x8dp+EjMEkXz9xtaYSLvW55
juH9qgBpwPY5CW6QZX57kpZO/pw6la8i4CGYaPEwGBY=
`protect END_PROTECTED
