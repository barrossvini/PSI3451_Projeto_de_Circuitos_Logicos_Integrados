`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
augUOF7HpEHfZ6oGG70AHMNwOJ+HZ5qQ2kY6TllIRx1cfy6AC1+QKYXnLvo/8hDd
0TeoBvnCc2u8SlW//kW/Q6fjs2yEPTZDabVT1FxjWakBnbyEHqPzERr2rSJABuda
qCZRLrQwQEAllEM+oteToeFXlITCsvDHQGboOdHI+Jo2Ky315A//XIcLt7xD3Vce
ZDqUmyxI4H8Bg4dkeeAttpy8IOnmYP5PANsgsGi08GdI2kXvpHYyXlVE4uSjovw3
QKuA9hsgtOMDyZZ9Zo68AXCKuWf7V/B87HTADaMusM1BX25HlNjaZV6MC9h/zOQB
bHIj3zSQJJPlMulv5gLVh5B1xHas0ufnQJncLsKuXlUu/zQ95d/rhBMrNYmA3Le7
X9X+otGdQOxq1ZuBe4Y7T9yaYD1lZ9fBHTjtwnAAVDoXEChs2GutSSIJgfkHEw07
I4A8RMCVUN4/6pTPZ8aDb2mrrAZpA1GTmJ4x48sc8NtMGV1ORJZICNPckCIxpSt/
xBapkCy70dpBStYQ7zl2OtOLIk9YEVOg3VwMJgZZyylMrW1q8rdixHxTyRRmZbW1
AHF9afQ7oOc46RX86MEB/6wiBjWs1usKoRy4GwmU+CRFlWx6Pwx+T8MuyAePrxMR
r2MUioBo4ntz2PtSUa12hL6TbrwUhqjaHb4TfGLqjpg3OUX/6jnDCqY38VFZJwfx
47GsLCZuHpw29cTb7tm3NqFtc++QHZHFHE5ms0NG6WqrUVimJuBV6wxOTZvCjGCs
7k53/LN6WCn5ccDpKLTy1nv+RCqz80sXj0Iq3ItD3FONLDM7RhqPQ+eX4evCBSm8
TWpnimRd4j0e8KcCXDK7TuFTTESBp89hnvuve5CxK8b+zLIIS1eYrF3l4hEVR+1G
c+2NZEscLmQCyd5+Gb3XdyL8sNJRAaaW8HCRF8qZ4ORhGI3OeVq888vIg36WJpCQ
f/+Mqbd+FYgAVsgvEkxxJhoM6BEQNP4XNd2uByasBGTyiHlRMounYTwylMtx0DyD
Ow2Wlyj6XyyWxAO5RgLhZkCGhNGGfQpI7rsvYicLKk/ABfCpkvZ2v7uxVLnkOkw9
fP+bG0Ciaq5+3d+s9C7hSGoVEoTi6T5gbrPQwDEVBHtS5wP8jfINizAoBOIin8RH
0cxBO5MiqFud/gC73xRQIdTP7EZ1NLRJM/f8fNc6dJzVDIZcIc0LQ1sedo9OdWD1
ir+xDex5e+/G8Xc+4gmjiwKmm5X/Tw5xrXutKNBGAXn2UKwGk1UdU1S5hTycCcwE
W7/NJfXM00mqUUG4P5o2D+m6Goh+qSYalm1pREsNABGqjJWSalpUGJlrx6QTEBpQ
cWKsZDM7adxrRhdVMjQb5wAbOigdkamFiZ45bY9toyvHIvS5gqZlfBR30ySUAP2i
e8TLSxWUgUPGlnmiDjpcVC7gGrEQdETv+sHQ+oeYbVmF/RcW16KwqtMEnLlU598g
ojQA18tQ/ekhEAQhVyZmJGjsSkU8MRvTCBqgT1rXjrgZz60BoVIXNQtyOYWzAfeH
Qg1PzJJ0CGSjYPNO7Lw2qZh1928sVyyEg8zkEKWsQqOkRwYocqyr9AigFOAvf/HI
p0OIZvW+iPlt5RDPLw456czM4uYNbG5LuHfkMw5MVZg+Q5tR7qHgE0o5WNjhJtyT
zYhH6AogRpNp8ysoVCQIaTjT/+CQUk7NWx/z02dE+SZtcBsvV0M2rDX0hcNTY2OZ
vAKWLy9UUU1agk6p7FUiXKQPFLM41OIzyLkrwHjNetK0EE9nQYoP76PzFO3Pjkxl
w7fo3KEoHXGjWoUOevSeDYkKk1Uttkk0mYaSR5Ha9JHVgjvoFImTM/3kdufxHZxs
xJMGnAsRvfKxY16p1lrrs6KnqULr5rYRcNivMhjnYEo0ZMuzjnDJLMrM6KBFjmfC
XN6sRauyFH1GEIhsPbsJGYrqn5fS8NSultbgFYzGqAjEHhvVR3/UH/0b6udaXMwO
+wrlNqffvidPwuybaRZ4I8qJ325qILVujphAAChgmDBCsUGiWkqo3D/vphSz8zvh
E3LvLkcEKMWNhNfSi8fYg9knNfEMp8ZTkVydym7MroQuY6w3F9oQg3niqsKWjyPi
hWBGvAaO1K5Amwpxkp1MxewY8+YQfbgAPH03MVkRW5g+d9CIvYFvAuQSZL2Zrdp3
WTJmOC8qiso1UCT2W69Xk1NYK/4yRjxAq192FrKfHjvnCIINioidw9LKs7Xp10ug
4dHgClVa/wxftRp85Ls76Ozq8ypBByVYXfA/wPmIOnAUP7sJCDy3zHYQpcnbQfHv
6qEWfYLi/ekr9dObnkHE//GMMNuhT9YJEuump+kTedV7ER+LLPE6VR0fnhFmuhDD
l1kJ8j0enoSTeAGCY9abLe4pqrpQHCh+bhRZSgxF36ru1L0Iyvp1hjzS5wVtZP3p
nFxHuXeXHHplX1s5afDl9doZ5zjcV5LQIYsx1BkS1t99/dA2Z8M0o5KKiGJDXNCW
FrPzwrN7yXtpXckEIZLoNYWDstb2m5YfK8z2g0A51lPscel3iht8eVShJiCP/x9L
/dnf+rOoZq1BOulKqgCkospMAl8Np+NXKtppWLMFQxtSrvuoaLgA52cOWm+hHw+s
kp9+/sU5ou6EO6LtxuDtFH7hJo3Vk0F37FHUKJv/UM4F1U1feJPuUUcy8nw7V9wZ
cy1KsZRd/jPKQrh7kuHCIVTJ8vHQKhU0d2tDc3b4Rzat5YPkjIn+DpDK2D+ZK/Rf
Ugn2ELAca8foKNhoHWtWvphmZhc5F2Vu7gBkueVgYfxqtCCM6Ep4fhJyrhAAnErU
oc/7aWwI2VS5rmGzA1twcQs+I3d+NFwqfYqpr2QeqqQ8vd6Vpjp7QN1ZjJqrTCBd
aPll4dXPc69D6XfeXY73Mt/HjTldoRPjigOOa9oo4C2xKe199EQpj8TJZoDer/m2
K8nAdfb79MQpVKs3rabGVkwbUZxwuiFUwSmztiWcl6xnhUbg1t2xD8fcSOWQ3XHj
8y7yun9NklQ/Wtayp6wMJ3+45rFvFCU/gDYw6R7S6jpT7vuYfx9Z/W5m0HLGDq+Q
ibZ+N+fO1PJ3xnE7uHaGAuJVrUCvVlBjDNgIfeRL6z8aAZHCvYHiAER+PznWHilH
gIDpdPJIBY9cDa2bjneZX415OuZ1XrvKLuWjcvM/IzOqfin5P5Mck11vvP2prqI9
8CXRVF/CpnBShKS8MPnN2TA4AIbH9zXduQk0Bdyf6afdpl9t5yEp92gpNc4FXmeI
0/t/I1GijS8fA/z+00KuGOBv86OnwyVPuOSWHg3SjDYHY45DWNRrsN0BAJ3Ulrk/
CjY7H+uWlGYyVPaUBAVZWsZtFFxuqFx5+f1QuqCXxHN0BGVKFb536CuXB0hOfkpN
X4h0m37OsmBhiA1uOzbNl+ntxB/XlEEPzyCjB5nVrvoGxG/x2abSX71+Ow6QHnVM
7PYnI/ZvjQE2jtGUZ3OIJlNUPoIdT04/Pn29WnegQADvGtHDdgQZJxtn8ZvmJg5Q
Ful9uUw8hgyaqJd8OowBCvjl7tgLbP/cMn4e1rOOmjJ4qpJWVsGNKyGN2CgoLMWj
fyv/vFKOhrvvSTikqs8JvPUzO7dKPwNuIcl26kBY97gE7zeMjDqOXWv40dvRfgCZ
NRehNtc6eCISCol/xbZ8poqYp3zCe6vtgqZcrn+b81U4meUtU8Faq3oty+QnBOSp
KowX0SPUOYav1PXOGa977zSfQsAdTLBVmLQoddcEZQxglIryKIgI/vnJOBYQCvBi
7uZUNpD/0Y8Bqh4peb1S7rjFSqQHUk+yaAiajXeR+wP7E8J+ZHYpBre8w38baX91
xwhutjNJISGoZ/L9DUzLPYaaEktfjIl/7wuIzfvclMv7jEWXdzmLTBQWeJB6PpDP
DsAVXF2Y75I0uviH4P7JPhdxexRZHn3HbLQDMPG5XIcK++1a0PZaVZFh7XOvhRGn
RRd79qUpVqMMfIxp9SKXqTgBYr+CCfTIaQ2qrc1NK6zjT2q2wu+ZECmjbhBE+VTi
cUMcgohJCF1FaCBrGjS3m4I7GtQ3ZwcIIBqf+6tvyr7L8MSy0DYedBjOJQ0QRr4/
XNnfLw5AoVDovdn8haQX+TJDOIB8ZRERQ8vg0yHYepq/WN5dfeCtibRJAU10FsIy
y4Ibv9a6OwiWUlcCCuAlGxnLwkWl7hhgF26zFI/XGKGzck7bSTPquPF2rV18t252
F6h41hMUDPuLZNMUNY4mOJgKnozTQivx6s2JhL+L1JNwBrAnAqzI0u5k8oxl0qj9
7LbFZckduRjrM+kvElFK65FhDcR4anT27J+BxH9JL1kM+wennAEY7zgl5vjIuaMJ
tJ/jXKMKYxiWiQd+khdXSA0OgA5Ioa+zA8jEBEyXkho=
`protect END_PROTECTED
