`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yOUtFG+AIlbBk2TN+SIGFr1BeTs96QbOTf+0z4CzI07vjTVjnBi0PEnxGABxCn/v
WwZgKwUXnpKYoK1cYVEh3pvIIanAyp6xNdce1kbrw8HO1cXXB4dfJJHuP3mjIJ2W
9rxD45njckMkCzuJ/ypZRV+9tqQc5CSvp/qqhiVdyR2iNKp561aM0e09/g0enitD
/iGggFNhkuyBukhl+UOwIaDjmlnTPTZPvSeHAiwI8rJY8LVe/Em9fWwj0NtVQ4xy
0svmYZQc6BcWRWgBhCyOVT1OPoHAvdC6N2c4e+xAey0Xdd6Zvjyx35k/0CdEGRtx
9cgycSSxJ66SQYD2sRWEqghsr/U39AfkXMYcVhF7xH76XoeYx5rIVhB02d+MogTx
1TG4Msms6tIPKVHc+g8stpGDQLPuUB8ECwCdkumErhEH4YCvl+lzsCzkfo/z36BR
4jQjvAwDjSKVS2e4UPGWna5hxIObZZkWxmVNi3lCFhkvg+ycuBxj/uvkurWhDELe
2ZQIY4/lJer+mAa+qrqX904PlExnQLujJHI7IltyA2ttfMFjrsmVaIJcoCQOF5NC
Tu9eXj5/qYObqf9JxY2GzlEFMx7EY8e1YvLaIYnrKhLJr2Lc7EVLQLDnZuS0YDbs
S9M/nyR6ZfxDWP7IgNcW6kC6MMOoFAekosfW5aoKUcLjmhCTjdl358Wv5i4yn1mh
ssf9BXsJb3Kt5qpEITiO8q4cEXrIEuHtSATxr7t8+NIvp8U5thb+8kpUrobcFFBn
0jQ7xxruc2gY++/+1+GVUGx646pTZy1A8KhDJzapxjkdW9EWYTF7M0DBu+7Lxq2U
aqz3L9xcGqhuhQK/EHIzONMKm8auQspnIUPPY1IfPTXhmGuf9KEKWovPLejeT5hu
2GJ2D+pFHkBwEOglhk69fVmnb1D11MhAr6wzc7clUP8zd9ooDYFNK7WFy+Y2K1Uh
gtVg7+PF9r+DUTPX1t4F7qyAgW7yRwkPcAwkyiMapcqRspQ8uErLZtY0ARN0GENc
F/11BadFTa0iRBAFosu3RYd4t1sFtypVSppqa5PIjNaGpa0kdPb3+QsvkzXzKx10
aShUSS/HIAFoZlsyb4yXYgDnXBo3UJyZ56kNKkDmSeeLpG0x7SoHTDN8d+NdBlCF
lH9VLDEixsvwp4aKBCwnLGrBNOU1dCg86+zvZ3GSY8kkO0tJoV22dPn6x0cQxaYw
rTIxGtyb2vs1CBGJzBtDeAv4M5bb71pk56/ap2EK4HKX73X9HeocKXsIAcjGRNUR
eW1kbSLva3sK7MRz//Cu8u6szQ5gumcPoUhOZhsQM1R+OMyNkeGFdBFUSWCUXgvq
tkuMBngnjy+yfCdRVl4jTadVyo1s5rbIL62w5VFV29EcynUqKILFqCq8Gq4IrNha
bEX7JruoDm/2/NhNyGl3bnF7CmCB1GbQ+HpJTmSxUtCmIg5DrijGsNd4FxGZJfyp
killWquv7ALdwl8X4zqSsCI/+nsPtClLy8VXpw/G/jcH/gjMIYvGcvsmhOk+5ZTh
p7DGuqH4cqrnwUGOdKo30xkAc0jTwLztLeak0a3vbfO0X2y9zBK2QRd9GydSZMmi
bWpYFVJ7wSfsYp7pS2VwsW0wIub5bxPG4FVUNICoUo4ydvmMYgJETugTnSDMIT6v
aiiw6nU2nKIBrkEfdHo1PAr320yZORZm2G1CvDO8lNnda/6zmwARDNAF1vfF59Zz
QTIsDNmpLIlPExqqnhQKbIlj7yktrGRqxCUWI8U+is9lD3eOM1bc1Waa9JZuzxKM
gOyqojkFRgJV4S8ChQW8QQ==
`protect END_PROTECTED
