`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6kVkfWGfrpNEkqqoLsIJLrfBtluHYC0hbhGj3f8G2ZeR7fGYjrT8qaKg2rBd2PJL
a34qIjtGZM1xNQgzKcrPKh8tNLy54vYrWRVvo/qYV3eSS03vV6D0+bqEWOHfjsms
H1k59wHgQYjbpeqvAwifIvGthmkZexaU875S3kBYjLZTXs3VpK1lJDPXpvtRSNRt
82wPEvdY4mhdNwpt/OsN8HZ7M4lw02mlw3B+QFDw20sWUzECJij/lmgkjDxA9Tp4
lZo5/f4DHF4Y12Ti1qx3zcRk5B1usOV5tLTjCjtwKbLWkH8/N5qnNGay+Fk+s76o
hc4bVfXdycCu/rgALCxodOst/kiCCQZndlVVSWriAj5F3svpiP4vU0uYG+xoCK1V
bJEnNzKCBjaiaZywplMIJVvc3cUrNF6qvMtzaHdoIMBL/ZCAjJ0bt5/uEdm3GJ5i
tbHuhjJRt9nXreg4ldEK3Dq2ASqsvlL4n3byR30JaAdKO7X9vwM1+28TQn7tOppR
atn0oIH6Osj64yqINkVPfzFKEgZk+atP3lDqJZjqHCzUZRT6HxMc//ES5lQjPEkK
rDN4YTLWAq2Ms6dr1D7ZFrwUx4R80L7Qqovc9uXk3OZCHtd49/hi84wQk9fjEKLx
OOWCz5ORh7AtP/L1SQ/C5I5TqSM6Pym/JL3b9WFo40zkQ21txwBSFSrr45FvTz1q
q0N4NsiqrJvQLlMhPiPPmMuIIf9Rb3cAoht97BS5xs43T22NTXfL6e651HtAH1Hu
u5h9fAscL3YdJyfZLZAoOTV6RWtDpiCJNYjcMaDlO/qHTvqso0HrnKhYwrzdwsXm
d0VlvXIUquBceE8sPR9bL9QE1QrJ3fNibEWQmGdVtVpSHS7c8T+ynXgTDIHW5wXc
LBj5hoGjx1NSTGiUjf5n266E8hvlYwnWZCI3QTMyKgPsObDYWBe14Ybi+4EMdMk8
l5xJZk6vGKjY3Jtfp+VYIzGk1UkOrRmgVRXBP1DBM1RP4AASY3ekAUqxbhq3ZJFa
Dqb/ieAwC+ic7sLXeoJqSEw+L+biMCuwH0xZXAGNxoqSvXL3uWr6dfn54CiRtlFg
TiTs1232Ol0LvKl/5RYPkZWRPTT2Yk3SH0UECtLmqA/vWuhyaErQy5aWyHdsn1Gy
jlC++FnOJ57ld9QnYjV5U4Q5eGou/VOZ8xjGbMHvsvzgLzuZDeTDyFy3Oe4Q4ngQ
/XwOrZJ/gAdutQxrNFrphOmeHxaBoQ6BGr08j5U7yRM=
`protect END_PROTECTED
