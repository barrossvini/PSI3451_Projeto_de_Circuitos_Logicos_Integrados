`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
taksoeciu9nsd5hySOIghXGTVkk7kQY4m0QcZ8NlIH7M8rce7AULV50WvEkZxUbn
5VVz2XJ34o8IjD1474pSpCHXLQPRqF9lNxSivZ6bIoZTSe8GVg9OXxXkkz8fQ02p
/njCkNlQ3JF5H81s2b8jzwyP39cKHoBFwGqkAe2BaDPQuo+xIZu+vh6jnqrsUU6B
8oLAc5kh+eeWeEScFuWfDiASCRL/QFwDwFoC4GaRXjkzoSmXYtBuMVT4vbQi1TvR
6ci51L8YO/ZBZYOJdzkCgqYtZhHaUMGECmg8y7ae3K8YRpAX/2M8pPRqLzdWX2rd
G93cb0y2gByAqqeM23lDuUM1hQsqtDbqLgMM60hrqdcDVMa1NIFkujcN12lHmXM/
wNRPOkl7cmjEvZFzq0c+cTdOVySnfUj5k1D4CRWyDitlAudBOGfqFnMG8xyNvmyi
WdAOJFIP0BVaBQ6lFCCNLai+q3q8w7VckHPMHKr8iNVsxMOIOmV5qOgXlC/sl5R9
WzC13eNE6tToAtQjRfU9wuZEVDIZh9h9mS5k0YINuAzzHbHxTGoyFUmsXY6Hs2Rb
sTggcEb4gSBGsktBJKHKxy31vYGSVLdCmPCM036XB9/bKKSG48ZjrrTHjAQ+Onr3
TxdQFsZKjaNPCvipExSibUlhBTA+9vFtwWxLx20WSZCkayLA0tevkDvfsVWvpKC9
1owBantfXPwwNNsB22vucL8ew8PFQ7egv/ZTBwbdX5brgD66VpWdWGd/yriSbNdU
6PE+lyYYc46BqJ8gcMNh4l2B3MVmfmoptRrtLJkC1vLkJQI5rg0/9bzd3cvxMvUW
zsvZa7CkfuHput+QFFIFMx7l0Xq1t/BBAIV2hrlbvMq1i0jONDh0PYW4K9yxAdq+
d7mR6m8k836Am09tbrO/RjKFk7SfroE4y3FvG93pQLU=
`protect END_PROTECTED
