`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bnsjivyytK2TwwJXssCIf3BIXb5Mbrob+++xwceIsXP9L7rmugVFyJ+ZlfoloMUF
aTc1zeknqolGVLq3Nest6OIOUqA9YMSVhzZh7y+m6/wDomJy+UqxsCVcBWJ8ccIb
hUHOinSoGv2HbrjBzkvtNJe6zCGcFEtxPAJVOpkMyLVgP/wo6MO9lXc647f/Vief
p7eDAf7AEco+dnl1UKdQa2x1ZhMR30URIS2U9kAWXAIwio1j6rKvshu/R+psxbSZ
VGigBYvbCEcy3tD5VZhSRdyIrnGECTk7ZqOw6WsZIibNxhwoHr/Ez12TaZZSseS9
Et+z+LpvBpaMzpHpQbZ0SwU5HRyxBntA/1Rj5ys/gfq5WfXEq9quz5BGFXWJYH8H
6oy3oYUlG5M+T4Ysp+13Vtn8R2S/8w4TEK+WDmr+0dhqyRkigSyNjvRfHh094LIV
jmV2VqKpDRE6CsnZJz32+Mb2a08fL0sCvQfODqmRMqoPvfTg9UOjNyZ1ZBdUXEwR
a0bbUONkJ08c7D4BCBzwxndPTjV9/J9nOL9hhFmUc8+J/l886BrU7E5sSctK2HXz
kndW8KPjtueocVrZbx5GbRTN5cAeTDtZ0qcRB87AeJ/+lX+zVtRz7hOUkj+TUfw0
`protect END_PROTECTED
