`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GqwGu2kWCmqZkc8PvPV5GtFCNSvUS4cENg/AFOnATaXw5uJP0Pz2wouWC3ejJVxq
YsWJBUnQ0k1ZdY0YNaVl/z1znKDZlh5jtvBmfGUy9BmO9v6voAuSyzE6Iz8sYV3x
Ea7Vmp19/QX2bVT27qjEPo6DJ2QrdORsXl3Owpt5EPZdN5v+ZexL9DbCo4DtPVZi
uD1Rd6K/ya+tKVwhjSUyW9St+r7eRTaedmLHyH0y9U9YUC8ckOb8lb+8kOdztnlm
/ovAPX7DWgp617X8oYmmIahbbTSk26JrmlgLx+n/1+B3Lj8nA9SCUxSlk2GgR9dr
gTXZZwneivaa8ptF5q1Cj/YWEfekKGYqvR9i7jABGVg9zJs06dpRWpEmamyi2Zwz
+DvPEKO56k6+ei+uUKO/qcC2aFuVvmR70pcV6C30k3jPvqbSKbGB+mYEDYY5R2IE
dQ1h71mnU9FJ2Wt1mf0soxpROxIUlXGuEurgPcfygYO5l5EMHFEOm42+bH74ouZ5
GfhUtWBEnLEtmVSKG3POh/eFA4dCHx0MQWjT7MQQ55xpWj/wjE5840ndkSAfSwey
Uk8igqXwZiDZBgBo0xCX7kL5W9jQvzixAb3SZfxhzTBNQ+zQGhUJcEd4/t9OW+Wy
Buw0Jn8T4aUxWG2p1MepX88fAoGnG1etml4julDYGBbpnkp4Jpj6D13ir1kK6EDU
uhTzv9NsC1lS0SQYwtCiKHsQlJegEU+S3/q9QGI3ENHzALk7DQcgObF+aKijPuny
wY7C7qHG45apVAbrtNaRWQ53slQK6XhJ5PtBtpNQjlIiqqEa/MfrMRWaUgZRUgsd
g75f/0cMlCDpW8Hr6YNIkGRQZWDDSbqVHjZPOTbn47NeXw0ZiD61z0dOORgdf04S
OwGJYkbqwlJY+lplVGFcHyvADU6K1vHyjqGPm8HDd9nyr6DS6ehZe9q5pwxJoBhA
AeJsbtPWw5tyB8jYtGyhQ+p46ollyB97BbIsLMHYP45gavf1mZfDyut7WZ5OAOO9
RfOtmPFiCHyhXV1QECibDLgSyJOK4L+FThz0U82Qi0wDfcc018/RuboZVX7yf0N5
ZywyGORRfXJJ54pMTS0uzhLKLdoK7RTXH1UAOXICTeS5oS0BrQwiVu64gX5t1uN/
TLCV0jMx5gGiv46zFVTSuhhZRTMahY/q10CaqBJpG0JKF3KEZdEtrGTJVTHqmVcZ
Ao9mzKsQq8tbR1gxfWlvqJvMGImncjf3WdKaJYCH8BTaGfVNa+O7aXJEbUfsQoMf
DQECfxWXd/09gXSrjyiHIyMnf0oafNlHaMX0tyzfZ1BG6+FBCtGiM4BVbwElZacL
6JzqzEQJEZsxGuG66JeogUJkFaG/D6EmC3wckGHhU1W405OcQD3gOKWM/85x5/Y9
XVert9xaTHWbWrXCFn1u1tiMZ+nLqVAd7ylQlgcfNoo8lu+ft8lqR55Nwoghy8yL
ZLK2Zw1E8hIbdppljXyc+XlUPu0mTQHis1NEg3ccl4flh4TdykktlZ3B/mk8CP2H
s97CQt3DybEd4J2R3jt/iMfyYCLyITFjMsuQ+RmVfzmw6G8GZgq2oUPpt6emf/VA
NYr2eQEkOB03CuPtBGxKtqQp2Te2W9OZsz3hPYoL1ng26qNdxlQ7xfhb9wXq0orS
`protect END_PROTECTED
