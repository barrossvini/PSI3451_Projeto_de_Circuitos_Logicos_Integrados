`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JsfI1wJuX4Puftj9YMAR0lAccp0fM5sOkEdhar9gfkS/eYj95PtAa8+X+HvpEkFv
JVZbooYieu/pTkdTvWjC90QqKkDqFHkCea8Xr9rdxUWiGgg+ZMLr/goB/6IZRFsX
HAcsohywXxWPszyQYBce06u/9msS5BVoxAL5ZUanHMOFxH7jy4mZXTxlqYsWGsED
9VB8WGlfG0BfodCHHE80RpHAmXvDtKt2HucJfmqlP0JaFUqwGq2palO7lRtZZKXV
ervG9zbia2QkE6BO2CQBnWEE/Jvp1IfoNiPROoyj9JPJzGNou5eltTUie0Cy1Gni
hbuKlTCG5bDZJyJcmGCpmq8aRNpiT7gzmC4NXvkhQFuoG28ziIPn/j74EJTcCwih
Uwrehp7z8XRs0RLIpnMNmwlZz0f/5+PXIggq0wEGMhV3ilnufVWM3vCYfJKB9A4L
cEuFk+jHL1wJCm8HFCdkCUMeWQSCskWmOnuf4nwqlqvAPNwpjuwRTgNsM/fsawMz
P+R4Wti1RBEK4D+dgNM5JtRbdpIvdyLdbazsUBRaM/UJulULHO1DWXTErR7YQFfX
DJGWFwV3vVr2AuNzyn8Y9tDYt3tilDChPtiDAUUyJZCFb5TKr3QEXAnjuC5h9Tm0
iDpLfkYEYv/FYkjx7GelP6cnWle+WVbFUc3ZsgFrbsQXkJHGVNjCTclZu2LAuRDs
APCDp3HWKKToVyH8b0iSNSb5csVEVG4tklkgzvUqLUieGYtUnJOkIMVPvnk6wa4E
9oHWjBuKSqKMFoScUKzqcBu9EooK7rPGMLDQSkCFZkuOdDg9YNBs3k4TDbFgJrVR
RGWd+CK1HtOrrUsGFiJ4ttRgkeq2mjOCxjxUQ8l0JNvxOCZ8KYf7yd4CfUtnUpUT
u4tyNunVoItyMLM7Nj0W4RNuD5ZR7AYjCfBIePGRlI31/+Ge2HaO8OmTHyUHAZ+V
MGrbZcrnSQfGzmVt9b/z+4UNlt8qOF5dR8sIKidDK4OvjrJDfcKOmi9Eat7mkY0d
KfJi5jWc4tAsGstACGcruiG7lVAFxGBX3Vpt5ItAppXROuuKhVSUMrwOCpR1Gzea
ls/fy5jOEIcilGrBPVl3HQ1C++ueIHkNGUolZol9FxFK6kOjSzWC9KK4xmwuoDdM
bNZeP0w/qhv38mhBvhYA6iAarIZSJ5vHHCk5P7XWnowxRznA8tWjIp7ClPxLuc/Z
z62LrA7khiZbz0o9XX/TAZzgFMNw9vyRyVPDYt22YUweD9ZuW4y/ShjK7A2fS6fg
hdPxgMIa8MixEtO0w1sYMG4aPNynMQU7wlNUn9GIibNb8nCnPs1fkyhuBcOzH+oK
1ialyGJjMtoQ4hIJR5P7re2Vw2QRt1mIsabfcGQQ+6+Pj/Zq1CIi+7/hdar7xRNA
CdUde3zW7E3kK+JVC5UEUmFTsw8f30ymJFY0ZQQ1h9+RVjScJIhi0HH4VdRiPNwx
jSrDh/MiWU3QB52NFnovCQ==
`protect END_PROTECTED
