`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dkuaSJnG8+MEauSPGHsvR/VregW1/xUs7mNASnPLghiMfhDhcbQX3X9KM835SMVj
b4qoCJpN4YXZOK9KaL5iXaT+8XwxToiV9Cm6ahEkP8cRzUMSTM1S6H66E2HwTQg5
07ej6WJHHneRagbX07/3GS8W9AUXBnNzj0FcKXe6KZCRz9CyNcDJlMnfH1H2mdf+
9QkVPVDzuxhjEmZreoGw5RAHOJPd/NA31VgwMXwQ7bw+3Rthpvb0o0rGt0AHGBSV
AuodGQO+/TasKgMAUVS18A9y9g5wdspB8PAuodxXxZzH81omN+3UCwfCCaVEO7wU
6MaZCtFuuPKMdZGi9AhtKsnmw6VzcTnJhHMSxECzynt0hPt0G1+aO0hZ3OEduOad
AOOJd+B729KJvT/cy8u1HrGgeC+mFEIW4IEocbcAMbiWO99k3a7n63gmOmnsv0Cj
+NPT9/xCmE8g5yEI54FBHLz/Lo1XAsZyHwlGmR0WEec7c4ReXdtaVn+IEf/GGGhS
Ext0PSXeu5nws2a2XHdTBd7azBw0eGVwgWlNDruDa4kvHSp8CBi0z1FuOvwJTBdY
EooIeSGfTls662MM5mG6FD3S9gdiW8qRuse+gjj+33X0M6XJI40TOfc8e5NhsU1A
zx2nwe0MCGf8oQK+9FfdHIMK2N/8LudX0XQoJyvYfb61zXTU1II8bUsXMFXYkszj
VfsNRERa+Q2N+GelwB3uuYCGqboG6MnZU56XxsayAS5KxTBNzpzb5tIiXbu5ts+G
`protect END_PROTECTED
