`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tl/K8bYh47QRroHJqMWGUKiX72jUwl+Q0wG8LBXxk27JIMWvNscFfn5lD/XG+Kav
IC6xvmS7VGFA1pUoehCovqqJ1gl9fcNjZLs4GYPvEqL1eLQl/Yfhw7drfHhH87xh
p4tnPw/5//4xkx4IfCZ4uTx2Umu5Rni1rDbbQVtsuSfu9jqlM2AiswzuOVehwCKT
a7tEjRm3iG4f07+dSbRt6EnUU8ha0D6K383OkNzVJkjroYBI4bMnakYAsRtksxl4
b1Tapnfzt4uaX3rbEII6wvJzbub8gXaUKP2kxiHN2GJnhrv8BxcmMwdeyWId2B9t
o6piNkwbBNWrnWGgnvwGNi4VbP6B5sKC3fmDD10CN6f3gJUYDuQZ2wkKPTKtiZ8h
CprWGKZ31mDnyccn4s4OxCk1Wc5EE+Cw+qqC4CwLDMZrHGVcyXj57TR8VSAoww/b
JM1FlGoJ4Vh3OqZlsB2og5j1Ozyo8kgVVgjPDM9NwERJXNuzFzq51jMPQpB0W0MX
oRy7lCbTj5b4ahp0qUZKu5CzWAz35huPnOvaXOq5bwTFDI7RtRnJf10VtQ75NWUj
t31BFlED3VC0gnRbe+LBORPHoy6mBV/y6VPoCcM7wOyOYtMxEOh+ff2ysaz1/OWs
OvdQ5SZrc1BOMNtImzMW2a34h7KxW37Wy5TVWgkHyL5qo3FKpxf2RTJNacvgk2Nl
Zl3FdRThNX1TBxwJdzaHCCG2s1UEyNa/VrkxoJLx6qrrjGB/gBy5HLkUYs+6+l0H
IUUD34UUBccw334Bz3v9raBKBWeEqvNlBHAEkXkpzqwBqM5gTH/96ZlwgVe0xFt2
QrNAyrj5SdC0kd4FlP6kmcTEGn4OEbudRHuqpjArvVV9ITbFFV4CrXlHDmbiK+7u
52PIDcuj4FpvHqjwjtGrs66BN3IVNeAYdwaIOk+D1CviF7TGvGKSV/6H+CVdYIBM
np1o+jM3rSaR3soEnFF78jyABm2kw0yh1Y0Q7P+03rddHEMrYiiXX268nW9Kau4t
BZyh8n6+s0igsRupq2UlrDR7xKQECLYeJ+oP48S/2ZTx1G/4F59ki55qnSMbHBuR
`protect END_PROTECTED
