`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nTlk8f8X+xzDMAemrRkqrRn0cPTn9nARgOcWuf8f28vEwcvcF7WCC0mrLevAYsOY
DVTplusxiWHXaXtQIrLM7g35QOjYNZXpNhIjBkfyLo1r5Dta5ld4DRlNd3ik7ZJT
6PT+2JRsmGNO6uHQvNExQsCbM9yHMoQkltH85uwHBhTx76jnu35muQu9AjgvA7Kv
9n5JcAd5IMsVCaubyfJeC0COPBNI4+QheOb0MOluZVtLMYYpH0YDReN2svDW/d7D
MTlApJhEAcNk288evqzQq7AGPPBoC2UztMyd9VZna7pdAVdpq5oO2noyl0UuTiL0
2gs5/2H2DOiplloY5Djgt2k3zzYGwGVLzBUQlSyP/9vAfkw5H2kc8ppX+wCTJDad
dMzZSqyC/9KlZZb6BjlKN6g1LZn2CddrfLV8Ko5K9tGpv9mnkcSV08n9UbVC7B3O
GwYgJwS1ny/Z9tk5H+3wFO75M+68LeSjcvVl9AJ9V1a7eAs9+zr23QC2iL0kZH6R
18FJtvCRCj5uONrq4MSa18G+5LyfsQohZuCxExCUPsc02Nj2QKG61bUNz2/r3N4H
6hJC8Ohhss3ZfVpTD7RLLkYrPIzYhToLYQnfDDY/jNBYGPf2inXQYJKWfytAtYmX
2eVJd9pzUpTc/ZISU5WfKA==
`protect END_PROTECTED
