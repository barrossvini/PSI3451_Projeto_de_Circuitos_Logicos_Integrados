`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/BY/Hf/2wqE0qu3bvyo0qCxWreXxnJxcfsci8mSgFS0v8ZPRfLPGJtmp11qUI3bu
UiRksqbrjS4OoP+ignLjlrcW6PzIvNs7Vn3+cupZcss04JjsS7+nbrXuRMzIClBx
7q300M9jq7ACUGZTtG2f61KutLjmoqq95/jRjByP+zNQ0l0xoQL9gHGKSdubXI9Y
T8YXcfuIpKpzfXH6N9owoDiqqwo916rnQWMdNUjVk3/A+n7wq6xZhcuaAaHQ3VF4
VaUXMNzH4RVdz+q6kTXiR+d9hKwJ2L+JKh6YXjSl4J9lCcEUeSRyGee5p/2+Lzr+
3lBmPkoh1PKOxPSKgbwkgKIxMaI5hVJ3PIZ7nCuRXP4517nTlyMZ99kBICEjANYD
YIH+FbXEtYtHIsTB+MUFxQ==
`protect END_PROTECTED
