`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H6fzWrrg1VEbOLFDNs90QMma93T98EIirrpD6uZKLWnvR0SDskmK0AIbJjUZwieJ
mXAsiOn3eds5IpDOz3GNN9mMce3oMGxH96Y7N+HZNJvHXufGam5Dw6hVLY1d0YNs
31SNnTQrxLxPZcri1kI3V9foqE3vvt/Ku15dzDRJunjRSeB8jJnvoqkqBo4Q9jUX
pHe1CTvNzT62GDITU653DOhF03EpysqmYpk/bsxLWr+yMpAreOx6Fde6u8N9F2sR
0YUQNg501eFBPYsx+shB/CZ8bvcittWOJEcY9NOOX/RLTjDZuUpYBLmk2VCmPvGk
niI3M/8jzVaoz5Wk4kwn/HVksOnf5pNiCGQHtFLz5dJHyL4RchGlmO8LzIYj/ja3
I6TI+3zgQ0R4TrhENyzxqQyUWzqyxvA+m/gVvpb4gfP79JPsYiUaChmV58ZDHPw1
DgmUnMHafqUrH36Lal2giF1uTI9pNaOJGfdkMdfX8kBFrZLSwpVS0BObHTLl8feC
Shbwkhef8Fb8f2LivW5fTlod5qfT64j1j1VoocCj8JTPfnhghg/ghMuVvKU2iEPg
BdV8xFjzc8POJ7UUwDj86oVhWEJ18pYll+kGdMTZYT63WuXTIttuC+yJZXYBAeLc
g84xN+E2+2PReD9X3vxNVW1L/otwYQafm8Wa7V+NheXFiN3PuF2wkW3wUHE/ePIR
fMeW5/ui6JtBuCn1FpgmJpdO1Wh72BejIWrtXtouUQaV9GSc8PKvswVxLxkB5+U4
R/po48zFa0VoMeaLJCPkJtk5AezaNcsNBt0IOXzB8OnsXrElcY9y9204i3e7QmOm
MZ16dDBbxlpsMxr6EP4RCjCPEOpPwlOaxZIi95KT81tERhQgS3/d0l9qE1gYXGbl
/3tZQdwKNhF/FtLWI7VHqVWfydAN8w8iqgeM4O4WzYvvsS6FqoOhFeCymShoAt4s
Qh8gNJ/MJjT1SaV6uhac6lGhJCRzRT2dXaHvz34WHdQgUY5lZmiFUVnFZVJK2tIK
zdQePm+WexXiqDkvakGpuc6c0qP3y35i0qnFulvp6jr8Qk6MM4IbPuHDxgT32odl
jxwy2dt4oIINvvpm7m4pn8feDIlzZ1+IsrkniXnr3yfQxd9EdDqFL+S80I4rZo9a
nDwaKMy1R77YXIMJF9y+HO5+Sbf4sX9SU2FTdZfgA7WdoDT/7dZtQPSxVUjfyVYb
vLDThqwIYK5Zq7elGYJEMgoXRrU/2lux58aWez3hUQ9SAMypTya28jWtvvDJB4oW
0TDLOmNXjbqPa9WKYFwJMn/tkXNNVAcZ7/kV9s3r1DRmRpUuIQ8jXNrQVkR+7LU6
OTc5cKYkqy00BneiYsCUflMh2wBboQizCGI12RD9cJArYYObnteGsqS916u0WjAh
dLLZSSBTAB7WZOQwbrZ48VPIXfPChWexEtd1uMUT+Ir8qf60NHmD2REplpaxeGXd
aey8WuQQm2xgm6YbL442yundvUtLKzitqWvjAqQHIvQ0miYKqLjgim4FX7CRnA5W
ey7awmUSx1oJ20CF1OaPd6HFeZivBmNgf/2FanPjn6VJXdpSy8PCpjgJl+kPDihX
8dY1+JqhCqo87LWpzYulvVmgUtIBBi02Hrh5dRVuVvpZ/b+gyY9jYdTMfo3tsP5d
4AEnDK11eS5bp7AjSQYgP02rOcmHsPZLzbnnfJGh9TEXdb2DbH3mo/HhjI6DvZQ7
0QIpCjbpG/oMq+Zjic8CVYYqZ32vxNm5tMFNVuavSgUla9WzZfIVTjzfSziV7/ad
8IRWwuhQJeCw+vnZ//ny60a0r5p+24/5H3JXRvABhYYSgey2f1Zkn1uMfukgfDds
YUnAp87M2nLyUJfqXntFb5IHAOkfzVa0M1j9rY+m/tx+c6gJYGJiWcs88LLaeihJ
uGj/EBcJ6UzFFF6M2k5DkkzdEp/2Nvuf5TKJwxeCv41xmhx8lCNGnuKZh7q7B7h8
RyZrVjknzQciSem30Z6nIM8CKJs5mlc6zgc3T/1tXE83QGEJ3JfiWDyQt+2JWA+G
vzKgDLJoiAtCwVDgEXHP5i/u10iEmhnjQGUayNnZWPuFHAP07tic3ZrkKvLkUv2J
46gvByJF60Q+/lsuBGOJ43Zd5otra3QkTNtsCUIJT6vi1XlEM9s8GHiRFy3UImjn
yzIsAFD2WvmVvw+Up7A64jedwYtyTjGN2oDictzcRdeH1wFi5VBcjdmy3y1ujyRk
NQEbSNfpmQ8hHSKNEx6IGmevHXbbhfRZ/4Waw1ayJr3bkq2whMKghSYbFS8YqPvc
BGrV9QS7KnOYiZHmCWeSl5P/DnXqBjNiW1C4C/VgRv4XXo9pNR3vg+g4Uqj5F/S7
cAwBySY4tjFSvMJMBjl1DY18G+2aViI6i98lJjQifgTp6ecCiKvlYQvxTd8ID0/m
Fq9X7pUQq5P5VRDzGnNl1/1wJxPTXQPeL0QNIU5ijQRjbqHnuuc+qU55g3X8WnVS
yM1xCGY/nhybejECmUXDaeDInKHcKkj/gbAqvH1d14eWoqosnEJ+o5LP/k490ph3
unoQ8RnbbK/BMgPbXamfVnVFb3Vk66Y7+dh6YXS3d3acnaegAAejGH8ogS8KmLNW
8xKEWTde5SLR5DdA2FE+LbzkrY8r33G00SfvIgMpWRv9gLv9RYMLk4P6XgCrEP+G
bME0Zn2NBh3EroLvVSH9k46CB1u2BjvArTywTptxcZF9fmCowU6U4pdHc3ll3C1k
6SoqxhLfQOe9HsQx6k3bNag6ta3QOpzKp/dplNG7/04z0I7WJ1PDKzmJkk2uwEw8
r4YPXI5Fu7OLbE0xmfU0IFlPKWELj+8jxBV/lJ7vO8GIEFF8CzX8AdRum3SjXw12
mjmC57DaWoGK5WkBUE6qd6f1arSFzAbEgioo/m6CRFu1+L4ZN3FM4y/hFXGAzwKc
+v30f0e51pCq+N1dfXk1+9lg9jamlELWdLMj7j0cUGw7c9pP8GfSLCPoLyCYgZ4A
yUUBiTWFIM7M25XLmmjlQdt3YVqgXCK+rMkPzoXJeK9/SwaY3DTz2p/7Ovo2zAzZ
lZcFouL9ZfNaEx6fFB+0wOJOy7k4bDLn0LrJKERZo7nUH0UWKl1PG8e09IMUkiV/
lYYzkA2CJ95+myUEOSVb+2EsD9ON8xrUxbKcLsQE2IOePXVeDXNknpNBemHwgRYP
PCfwIVQtuicMCh6jwdT/t6lXvt8fsXX+5CU/kbmGtHW5xqRlpCA94TsL3Vfl3Isd
BkpCianIlS80A7Q2DDr0HQRM1fqylHex83nFGTOZxPIpquAVFithrePm3G8wde2e
aeA1mc9YWwic6Mp160MA8KnD+qeeQh/Bgf1Qr1de+JUWtRSvGWXuvQO6wuHhmwsI
kBZNvLeZm8bNTDau6pUVHUZEojw9VmEN7EqGVKNecGndLX7pBEO5GDtl3B/HgMiX
o+w5mtg1oZFOunULCyF3QnebFpH5EGnOx/C7AvKAOqvYPvz1OcfuvxTbKGgMUeYg
vSC10WDB4NLUaXKaDTt84hUK+Rjy1a7Ot3hYhB3Q/f3FLysMKetE9PxH7x4GLgW7
YTyhuTBHHUSJlbAkIaQwM4/ZJd1tsWHihyOkE/tLP9G4AC2Lo6etWYD2b5TVtKza
oNSd8D6oV+M0Ao0Adhks44b4YG5fk/sIH8ZHoILiyx/x2CTJvPVgnA5YCw+O2htJ
GlESRCqjm6l1wHTLwxOw8u6rx06Ig5tuysvUYAZDz0LXMuOaQ5Hyl/zvdp+VbVE/
PsKsq4yyO5F2fTwaCCTE34k/32JjV/j/Oz31k11Fx54cubJDSnYjLO/jYlLgz+E+
blcPB0Tp/w0cIxKfBCUq1u2zrMrZgbpNr6WtT5Z2XsxBB3IHHl0yvyGlDwr/kEgA
Z+p2NdpFj4uM5v2ygvDKL2WNcjMn/2C5U9Rtlqc6jYArRg7rdo8oEVMHQ33rlRp8
hMqE/MhYuSwnqaDmqdx+h3aXsUiRKiKrsCD/c9pjByUAQ+M1JQbWUt6GBKXFF3S4
ofFDdJmKYKut10XV9KDqLr6SVYkg6lOSwbVVvuWt8MkF09uovej4gfKhjf6FgNQE
ur91hioZFgnuRvKXb7FRk2BCv3UKvJvVQih4Kf3P0YpsYABokS2yMb4T3jvLhNqT
wuwtio/GSQ/lKKOaA/9dO95zv6V+E9zC91jDctJQ9JyVLFWl475CoSVpBKrJsJXq
VTyShgZdk/dO/lYtrWW6rXkzWgXZbdr7cyjZ3eeNBiKuzft9oYuZVRw6+PXF+z3K
wHHKdrod2bQSPWCVZ8IGiG24RCnAF1qdlRfhU/gqxpmtTRD3NA4KKqZ8TI6glx02
/syshCulIfaZIESfhiOM/FaAVj4hJ6TC8MUPDLL8GJPL5/I2KcJVolsJAjManDkk
idVhs5uM2UM3bMiyGnQKpm2+JbG4w4O43HFGGnyuBUT7q4qF2JVmvPsK4liAHXAb
s0ZILgbupbOZGNdVhydGeIJpZBzxqblx8Yl1np0FzcALFmQrvgQGgIEA436w9ls1
imf3o29LwBl92hFq5Zz95ud+NNcCMZFw1MG+aN27MdPAz/hLv4dtYj5KnV89+M6R
b50GdwctQYfWEWYaWs8yQuc9RUlWCQbgrxpezb+YxmbIm8OcG9XGeHeHGqfcv/Uu
k51IAmSGPHFTzgZ9R2A/WbF/Yq6oa00dd6GDgHOy9D8hOSeiwGkGESs+X545KjcH
NUvUgscnNknxkmiy3ZSUD0hp+Qrn6bnFpCkDbQ2avNW/wGWJdPu//3n+Jh2LYHct
LldS0SFIW+4ypUJ+ehfZX4pb2v0ldbCBcbXTfLWbAA8OTT2DWbgJep94B/FgOhiX
KDoRRYQrSixuhm4kpOywHSteYdBpTvLDD8rnF3iwf+nl7sXt7UOmNs4xZZunaI97
MoKYXTeq559apl4l/EAghc8usVK6QT5D2wP5tCquNWjMi8hMF5tO5mNhrtMtYULX
ZCu/FA5N1Xu8MOmt2P4I7fmgQ/qsUrTovIhg9z1FYRV2309e6/HjK6kydqg6u1kC
7wWhqHLCZ3PYB4IFmjzGnQE1bBnLSGeczwdjqRgUBKZbtow9RurG+ujyvxn6J8gS
A9QlhkrbLJwSk9vWiU/l9iRGrzZUP0+DFjMsHamzXqAotgnUsX4N+XN78E0ryof2
lfOizTYhefhOjUPUQmIa9uP7sMx/FXZy1KafvPWRN5XcL186msVJucm5hYlQRC6q
NqKU4CypVBw+DY9Z6ITh+12ctG89ZOlu+N9vCZO0iNxdzTl2k7vU/j6Aq9liwoXa
P6VoC+weX9qHMSxVErNhtkRFXE9CG3kgyeEZbOrjX2Z/GVPh0rsJ1zIJ82ZifmJG
mefIHFFUnU4FJAfbT6QZl13Ntcs7QTD+DYYbmAqDStTgFXh4pPwRtfjZsxtGJNQQ
RaZxIVNh67cEb8caA1H9M5qqnaMSMW5Zm/EjZDBQB4aJsoLYafOvvgGk5e6aCPwN
ZQwl81PoD/mKjeBbkh6YOhyNbcm4uP/2CrXf/qlI/jQGcE99E2eLI/Znhf2HJOrk
6uYaCrijqVnj5ClITTuO93eONxow4SgPhpuhH3DI6BuCTDHXk/sNQx90Zjc9ivZy
RoS0JVvNfW6T5Pg5SA1SfCbj5d9CtPKEcQ7IR7/Qq+ydWWNC44lxR0rqgMzTu7T8
yNzyUWI2decCXFYY9Pje/yMQo9LhJMZWBJvOKE9nV8yYS/Trc8jigwC6KynobpZg
m1qZZEom0k8Zf5zSpiAQSJw/FBFhbQdssktLk9LBHqoWLYXT+ve33rV6Wqt4c7vR
Vb5AjLNyjDz8nvxyAmJUQsUrZPSxhqXxAE+5SCwnJYt9COwzSu8E63wzvrTS6ZT4
/6v6tAvhdXuhfctFcQ82ar6wI2hKyLBNYLlzGCbw02s3opEPZ7nd4KahfAl52r0c
6B45aEORbxBOUFyyA3/WAEa5M4weOZW6kgM8m8V2KajdfHCCpi7z9tKxUBtAjYdq
Uaf99FbKiA330sJ2Estc5gwnXjq6T+w+f8y3/uDEd/8iyfkWKaVIvlJxeP93q/NN
jcmWtKiPKt7DOyo2ggiosnyQyEynA8e9hkRLPEOi8b68lgMweto+TmGXeUjU3SRY
cZlbfySLqBKsVLSrAX2S6zJ7GTAOhmm97lMaEtL28nVenNaFwdtFaEII2URxwKZW
kGSDDO6dY2dNpRJc4imv1SDdgqObk8k1iTpFboOaHrJZZv+wrI0a+bOYSQd03wIZ
QVqOFMku+p2913ettPouL0FMf59iNU8LJeNN6yc1ToOT395XyvYoHCyFYy8aY7jz
kgdfzssa3l2cd5Jqk4c+Ym2BehjSAHOgdMGRQSEtJT6VaU+PCD1eP5fxZIQazL1K
ad9c4TkTnXUy7INIYVnavdO2QSmxMOcLvfIIqSLCPVhO2s9tjBxrZZADgmrL4HtR
Xrs7tQJ+xSCEVltPsSxcExwlQSzbTc3pttlnWwV8EqH/cnZobdH4ORwcugNLMEUK
135/BNCyTnmYYSDvrU7EtjRDJPsIB11fjk+PmjdoclrWO9xUqb8gvWaLriRMcsIm
MUH0fogmeyXp4Ia47pz1/LzFAKn3junFudhs2Y3mAcwkxvH6kA0vcGKfZnnUtF1J
awSX62KH23eMP8zkmBOpFy3b043rWflomOABMscm+K7xiIEF66zKhUK0QODqV0bk
WE8rW49mOr+fGso390VRb9Xybhu5PSoUjgGdPQy7nIY3MplJGkTsxf++NG9BnJcW
n+Y8PvkK+Qf9gTckhFkUuwGKHKvjEgGLXjtUbd/b/LeyLLI/NhwtQ1f6nQujNGSl
LgOEv4PwjanYjJzNNW35KxArCltTDazpSiHZOtpNZQ7dhB6QZfb7YepNZJZ+8kgr
Jl2Ninwbf8k1IJybmNI98IR9DoxuXmZt7md7HsHeu8XDZ358oO0+rFvhdYv5czWF
zIyzg9pavl6mzAAf3Dnm+AXjzCamJwEwSZgJAm15gO9m0PcPqhi2fh+uqxREukhH
nMiTYoSB8Y4NcUL2mBhAYRtG3XvCObzz1UyndRD5rgfyN8DHc11GTzm8WG6zdieU
CfiDoY8jyftcr3CO1rkxmH3apSh/n+U7Vf+kPCOeQaDqermOvQu+YJePXuRbuJqT
bk6y28PJN7mGMQPLNXDZrFKk1wHxECiXUIoljuPUCXByzJH0x5eCS2mMGEu1v4cZ
Y4etisRHYpEE41HcuWUZfA3GV4pqklAVJ8Aa1074L/+IVEaQPCA1sOVKUNeCtf4n
PHWruND/R+ozjLdmo9uYlydaamC8nKze/CeQwtfmVOn5iyL2LGq9fk4PSAIG43C2
rwK8uLdBwY+3bj5sa9HK9cOlS1CteIxpmakrGz0sFJoPwdRAvdoDLq+KFM2JU3px
LtZceZ06meCvOXueoRHJ+6zgWbsZMmxvO8Npt4bH35mK2oMsf/0OZqAB4EARbjC6
HvG3J+25fVSQnzHxQdxgMS64OyVb6O7uwBAC5px8eFjySzOXM8MSsXt+mLXAietL
OLJc1o5LQvCqxf2jW++jvJxgfn35P+IxA7TjKcQXaANHpNWQPnGOrU/aAWFn9BSw
C/CX4LMd0of+lSliOxq+74O8ZOKJbHv+qT/pTHXkIgh2pwNhs5/KLVri0m3h9LTP
azSZzPPbPPiao+dvlkGnJjujmVvA1Rb57H4fBsh5lVnNX9nS4vRTZQMwA+ir7qZL
Pq9Yichd37/3czMuBnF4/sGsgTCvjt+LmnNjMp5tPnkkDVONnjMhGphRg8zYS0Em
HsJEkCZCjFH8reZr6p6fco8Uoc7Wgv6tccJ9t4ZeWTN40PtUsXs2o40Pz9QyMhCf
j5HNJTvliSrhSNQWLirSwaorIfdHX0TF0S1ExjdS++yBtyC6BDFI2Ma23EJhj+BD
w9D7+ae/stnf/FylP6iP0242xCY0IsE9WndwoZ1zvFgrgizOt3BhPx0yb1kC7bJN
AtuP7FnNEko9Ro4/yYxNoEFfOSd9mM9BLvb+4SjjYLlXG2b9AIoZLaQx5qclGPMT
vCvnd1C/5BeMqWjxhiw732M9c56aoTkJqh1m1bkxW/oGEHh1wXXGSIRQguq7/V00
aMjH/IzqMo7YIq1h43pWYYXoaPtGaCppOJcy7RzgOgvy6I7dy5Rr4YkJhP+Jxv/j
jD9PdmUM3rNuwNwZnb60UvveOKFcx2rbzaMRRAGz7EZxcMIP+aX9WEX81dLZ+K+m
lQ27Nr7kKNALjXEh1oZdjA15xBY164mFAIyA+JJn+B0e3I5HSrCV4o9oaFNdvc3f
G4zhRNMKlRCUutfmYNBex4dolcXA+oDZnsoU23nsqpA/MiF9XMUQEo9NzfvGFHJM
1o3WbkHuKGc6/M/TjAQsMGfIv/iNbYqlVugxr6otiMaFEzIccKI2zshjM/KSzgRY
j+h7wGOS/L8U29dM93l+3HnR2e62d8EFEFvpwgB62H41zDGU124wDhORGqNPbZW2
VqvpOhqNAFYnDLteRq+qGugO2s3X8ut46N1+jCwOjxERG6UvHq6g+Lq/n6AgrpjZ
PY+mSSIBsvOOxd5MIycsoSkmpQU2Gx7MWlsDzHOGWNolLuztnRZKe0cd8WvSQA0s
rUnZPFp0z25LLeJLl4atnxUPI3O3h/QDZ5c4E5Lr6fzYpM4zhg0ltkVQxOae1czG
ZSxUyspwwxRE4R/ahYI8EtE3DWlXQNuOs2wKulVzNl37IcfvpzbYYQSN6oxfE6CX
OMQRQWUiu0EXW5aKdIInm72BaliGfjx87eGv4+YyEYvDvhsxdj6Vck4+TTBVvHs9
0rm98dK7D2CzD+GxE92G0gp1XY+FRMjWzgv4ru94p3Ls1xrX4vAEPH4JvyiEO2MY
haKwcqKhStT+OF4CRom+WqaoLjodKhvzGr9MQSIqwMFTmibqh2fBQqh3I0yyP16m
ChbOmWuac9iJNWf2Cn7gMyZEQsNqB+fnTkNR3IGPtDx+VzFmbMe23e86C0b5TWdG
ez08Thou+ktjkbYvlOdNH7sJdnwTvu2NPY8HUsHCc70x4VsZE6ESqQp/M7PgDpib
m18FKSajHa0HfW7NyWMya7nM+xyY2robsxa7nWMqUX4Cz5KNBR8vIGtKO0B5eP2r
m8gFZitT6FDT12hWFCau/VnhM2TTEQH5w9eBLQyGeC0xIpOA1RAXnxxt34kyycY3
JmTEqPaZNjBnf67zyNSWFLX//HrMIL3Dgm+u8mNskHWq7nc4kN7apY9aNcJ9LOYJ
ev8J7xiVktA72/TTJzzMlUxkBZ3yjdK1QgwnpgT01cg/i2gxXC39YuoOyhS2/bpQ
Ld7XTO0Uz15LSXWdJ0f1aBJh1+zj2ImO/2V82DrHsFStn2QB46nZFXwAszroOCGr
QE0OvLYzGFYmNDU5Wvh47LT9YlNMvtuYpWFdT5L1JGL2BmhZrOZNUKd6T93bpgNi
H6crJokP0ymIIWLKs8ODQ63GzSAJuYGD4As7nF3/gLWhbZVRKNp4dJ1uipbc1Iuk
kLIyEc2Yr75D+7BK1JhLhHWRWHToKPlp9DZ7l02h48J3R1JaW/kr/S0QX5teQxFN
llOKmqq5AOLQvKdbzJgWfhV8MxrKdPRD4giC7i5RQkM/Le68YyZfwsrLIhchtA7x
H8k16ajp2dMLsMHfL6sJ9mZJwFo4nqDvsYcih0OwIcs4zFMgp7tyBTRRiJe/3faz
JRjKN28J7VRvwj5yPUVIinUO+eRjKDcdcroFscc7f75LftxZRZWB7024SKQBuRjw
Ou2A0qg1cGY36nnf7LqaTKanvmGQAvcF5PwNWKElEzCX5OqflkQ8iUzjTDdl3Px8
syuBrNk1sa1UTLg1OgLRnQfcK+AeArm2NDiOGdA8WPkZjyh051Xjde+GSkHzzyTK
9BV5u/yMKfXHbkQDmqiwpWIVoQr1MTzY7/qNlSSG2N4j55DcW6GdoupHuwLr7TuW
CQYyMnTofDQvwZL0dMC3i+KCzKoSSJtcRoq68aTltBjV3DhpbqfuJa9Zw3SrnuSp
IPcNBXnXxo3n4RaVMatwGkKD7zAiHEuh6dNXiEBK1D3dhe3PtAU22ab3wTwZh7p3
9C+7cre7hKANyhWl048Q+gMIYN0NwPOgIAfii3MkLAR1iCdUHpCygrB/WWwR5fUD
76tQ9v0v4zXH/OeJeAuTSTrhTHwoFKJDiYgIIcW91GURdRGAZezGN7Dd1bIWtWHa
mofnuLhqjKs+gb4WzRMZxCQUj4M1lTOmQNPpbSkhMq+pDnZz+WEvppIsl0A2og1u
C41d11adlRZlIbaYKsX0or9pvhRbTGEj7tgP8zVeGLVKU2aDRS/s2qW1nTkchcZp
+85EHNE9hSZL75T8dtO5g/leAXCn6jjII3UVAIz9vJsq6Z/eGOQPk1gVn70erF6p
BHKD88YjO6SehGvysqzU4j7aHdn1uT/I4VIyQrTrzBAWwJDGVPJpjclt5QO5SlQf
DYt4D/QuSGAAwfBLIepM9PXSlSAH66jLGV1EdGukAg02twtXIp1Dpb+jBQAFcQqH
YUr7EkU4VrH01WGdw2ubgnS4dj63xVx9D575UONlbA2Si1JTKN/SfyEQs0FewvZE
Nxkv8Pe3vmBuFne4DHkUwGpQTn/KFg0UsxGaAP492oBBrwImJPNB03Oq43WfzvKk
nhKk11r8Ze/odiR3vfggxr/hAvazjffl0i7l6MHR4gBzbTxtSvuK/hVPzAi6udeM
ODfzxr2+UwawvNYJj/kdgPhC9LAjKFQCokQ9eHycfcUGJ1uNgutBiVoQKXevlTdh
NWW2li/8JcN95e5LZukEFOSofKv2096F5LHcrcWAyHD2qLN06xmTlyWG8Ra+vWxE
SjN4K8kMROwfdtvVXG4XKw1tswgn8/krckShRL3lJbTQAjv7OI+F9+z1fnESsV02
8Ido/EkfenrzOnmCNCca6NqD4R8aYh1GhYtSm2HAJJVdPFZOBYKTxvL5gE7BssGp
61Jvvd94al3iy/TT1Hsq3Ae33Y7I3d+C+oyU3aoJPP+SnQsZDM9lJBfGRrSgVVi7
9U7ULJWO5lQxNVTGOFwbekjpZMLzRVoj427C1ajCwNGIk75c+5pUBgDeVWCaerMi
RFSTDJzix55BiNufu3yE4irZWIt+sK6wNK0+DbH6vRc8NDmtNQryUL/DYDVUcVnp
VAzvdY9JDXp4cXY+g3XoAEIoxMybtBiY/FriWAjaFnGGQTDynOIeaFx5BW6RPzNw
UBrJmC10Bmw6i2k6TM4KSx7MfPD52b3dqQ2Aj72cm5/JqcfsXSnUTejOJCiD0nq0
sk81nQnw45jlCvGIMsOzDVT948FKdQjTHTanCTxX5R9w8saTjps7VUOSSUgpzVSH
ctVTxIcjagQPT1lcZwh81ir3Vz15U5bccINAIyHfRz0ZfukmiAU5UDKwBdysXPts
xMDmJ5sg8yNY6St6c7Fh8mAfssyEmxcBwANXhLxpS0b3yI1VuYyX6YaVSzSw/rn/
PMm5Na05ZRjWOLUGB6DrIYcsPWU4aUV+nS4r0YeK2/XjN8yS5G/LJwwHD5+rkRpK
sSmqEggH5yI/BA/rmuz1feI+svDck5ErZ3yHv/fsEwZib70HQzpKTjgTz9gMFm8X
1SSNO1rPmTFmx8Yxae+yo3UtAW+PQZx6bcf6Hs8uKed8GIWT696Y1/DIa6E43aMl
eZwLY/89U6fR73BEw2PfZLlaap2dSO/IgDXaYv0xU6x+sUpPKJ8Gri4LiDnxO8gD
mXE/GDyetX555hLvhCvt6AJA7lF/iOyHbHlbjtvffXYoyA/k7XKMD4MbO3RkNge9
6abeoAqpxE9NCdtBlLBv2ZNbB4KB8GHVFS/T2kYvfqltbp/Hr259H9Nut3cSZpc0
kKKq/YszC56X+DEop1qjU7+1WyZbel7KfAzZOFKJLBsUNVv9FrTJiVDjwe86WXh7
g7zPisTNoNyt4dm8b4N4gW0b97pRCv0EfHYsS4WBUVpFEUF3Ev1HRcCI+0vWISGE
bnpDOWhSLLoIRoc7jRAarArK1ZnpReBKoY6Rod8RQ3uY0/D9lmSjBpetNk2DazhL
o83j4YzjIIqCCh2R9OVKrpUIPgaO6ofmw5HpP5VUptLMIjsm69j0GHOPbpj/lOrn
ukSJ3rnVli52tefirR4rd+WJPG7o7HToMTPT9rsCnZ7Bu5wmQLoX7dOLsT6zeQnv
4EH71aqK3UUMl7Vv7NljBaO0hjadIAKvAt+DEIKxuKoxLD+HEEfnQ+Y3akS+u7E1
O/tBLgZvea6h4lcwkGgXwie/wQ7laeh+knVMnKNXPpCPg5SjYgsBf2hRY/V4RY6f
ary7H8HMigx+fPsgZwiNds6pzYuQm8K/PrOOgR7TZ1ixqzR3R3jhwyAZ1wyok412
ixMYGBC9B3QO1ycoX2r0KL8JLyZy7OCq5/TN2TFRulYG3LOoSi8j1aL2bnxgozge
zTjiREoF+suFvRzXaIDNySEftmB73DuoBJMx+xOHgt6rrIMhbDdOpnj3op8Kdq2Q
u+J5bAhXtWctxNdDZAYqrVC33qw+BDd0GYdhUI+Z1zCb8hAfV5Q+xOHCy4k3toF2
3iuOoIpQwB88YAKlDGjHV2DQIk9kujXtyc/WuTtdvzlEuYQy4z4Sxjs8uw/o5dii
tE0/XMC6ImujhTFGFoUCE04IUvugtHXhyE1OUQzYs7teaDt1g67KsGtzAW/fDgzf
R2ayYEto3UfrR1jEjZ7MCmzvmFGupw8TAgJCaRWYX7Fyqb8aUqXDu6Mk4iLaEKeA
YSurrdRw+3mpBEaJy8UAsFFUDqmefwrlRnMQ8gpAJSRG5fx1X1dJVNOrcPJ2g5sn
fMxNRwbKf7OmFTKzkYcYihSrz/EA/q7ZW5oKTDt0d4dB9jb9Oy7jJ8TgqULPoVgC
4oKSMchq0TlyDyLzMLkmqgKBk62EESKI3BHgzo6FYnFHKQ44tXjAV5a9ZfQ2KRV9
Cwx+27kndBhbQrJ/86n4vRbT6ifJMEQ4kgyjwjp+sC+o3xWCx6YZXisCJduhwjgV
IFflBPa45Tjjj+tVYpdoMwU1YTxorvOfu5prV0qXanOuzPhX/Y+RH5YG/3ItGule
D9uCbDz0awQdGgamehMYWlaz67PJHa3Q0spdV1pxGZmfvD/Vzi4sjk+FDmlXbBxg
Lx4a4bC7jT5RnCWJb2+YLxg206uvlor9KadmAASd8UXLpxJ+aYcxpGJoxs/ndMmn
7XcsEiIJUeOB/o3Un2OckwXUUsP34px+BK9vTicova0sxkY3mXBxEFtFPRsHAfik
VgxA6oMczcE7FF3TJDSGKZprmGl1L7cL41D6dv/turuF4eihrt7BeFHs1O7SfZTO
v4nDZ9tT4Or3Gz5soPGEM/XwfaF8EegENviLHEssm7eNzSIMY45EySZbS6gjWhkc
dRhnKzJMM85pBYGDbk6I11TwYalCqAKvB7sI/A33fE3P6qgPSlpLOXWsVl950d90
UN1pYvRuPfAV6gc6WhuUN6v/9FUHK7fZaxDKdDUQ5y6H9iIbhXe/OAxJr1m8C+FN
jn2JASFLw2fy/Gq9pyH/tiinsSj/8EtvWI4RXXayGKezH79ilQjdp5EuLeIR9C1G
l2XhNWhUtLzTYdiG2+lrE4ctqkVYaE5Bay0X3vOjMzE2K78KflUy7UAlNCZ7YGCj
thHMXv7Q9vyLfZ9GSONBlijDIUGfm54ptrGI4giQanNeLmvfIPTelRx/WmiFMlYN
iW7evcbVTDxi9e/m4gGT9I/SFJaEYrMUY+OoVmoBcTj3zxjcMdBMsfM6kKTlm71y
FC86+6Pc83QBHMeIqDnPS0DIlmHQ5WhSzMqrOzmtO6nGgwYDMKBITiLgoic5zip6
v/s7UD19qw/jf3KCZ/j4i+wtIjmV6rvDjiJ7WSxk76iXoDVwLWosEAzUe/BXjo2D
/qau6iMuMVX0eZmZJtjVrychfcFjK52gDtjonjV2MIXl+GON5AUZ7ZYMurnu+P0u
MwoIg7pvc3YTgJS73ZqgNCWjMhWNUWjOo7rj+jSRAGB3LChavF/s1gy5qHZzGNW/
FXkiQVh1o14eg7DoFm6Cqjb/t8XwQ+Nrxzy1ybkQ/bq3VAYsd0ue2PsmZpdqupiM
7ryFxuGRtac9Z98Bj0aBx11Vo/MPQZPFpFOA/VAioNsiv60R630YaIqqhDGC6LHg
EPdibOyV0XQpLI6k4YY1xeEizvUOXPPtnRBshosTTjE6qL6ytt+/+SD+G/HFqLxb
nfyzxyWYNPh07Rb2MUapBtmWqCk+G+C/PcVYLcf0CcZ2kbqxG+ldpu+I3Nr3eQ37
YNdEPVih73a2Kt37UYW/Rh/dJW159BQuNfuIts4BJGFG4J/BwF2RGV8gjKg+C6uz
ZaFwDWY1Rrs1sPedfv8mAN9+zvACOS6NiPpkBgJAeP/Rkc0xRmifazg/1yLGFcdv
AC33sd+9iGO/tNkJnNE71ilu7I3ln/yPiqCHvj2ICKy01ueLYT5nGDxaXTZKf8Mk
hqxGogH8K4Ajj3muyys0n8FkwGkZhKtgwFDOTbGOTZLL1o2AmNBkE4bqK2ofq4jS
/x058mRKhQwDZuxEkrB7/zc287CqdOBNf7H6UjndHQN/8UoK+0TnD8n6XFEoU6Dd
3MRKzQtjdMvdZIo/5i/grbVBSbKBwmj6yNd5pU2GAlKEIstJQ6pIMs0VAjirW8KH
T5C3L7pDLG7gp+1H7v1zBsi3hDavLOjlXTu6xEejYB9fPZi9dU9u5TZhlPSqbSrB
lVMYTfb1ZgM6Q6pChVIyuO02Oo+NCxXmRbmhdFcNMXatG8tcmHWDEsBYcro6niDH
74QoeqiCFF+ymYgGfm+OAGcsRqIEisYfS9CBGtW/ILHglFLDGem5LEOzBDvZaqh6
H3LHcxbbCGAKNpXUtfGCWF1v8VU/rbLJhQBSYjyWUl6WE5ylD/g9S8RmEf1ykjHB
a1UQTciS3y72/iAtVhS8qSpY/fQ8yPG3jP8zIFaV/dyTJDKTy5Yv85CRsI7aldhd
Bu8le+MfZRopBUgP+BO+fRQZpPGipScqHzguRoN7mLmhQP/CAuuCDniCPCvSYq4j
UvvsFGYIWTL8VQ9DMLTo25NhhQoQFfO81IS1k2CIHWW3wZ062hrSMnbIriknrfTJ
GJ64MBvOLd94WV4rb72vVIu9VMNNugRunuuMHWCZcyjZORVjQUirirEw69UVNKrO
pwav9d1ijs8EOglFXcLVX/1BnMQ1AyC7bOLs26s4UCMQqTQS5F4ZddzDcz1BXYsd
AuKN+0ACSe03AvVENqeV7fI6gLPG6mrX0BPqJXAndV/FZIzsghrJIWq+WhFOQC+E
c+MsEHk25mTeB47FMEyLOANfVLxeUABhNhB4MFfq47I3ycJ9ZExWPy+28uh5Xbu7
FFCvCnunBHKDM7mqV5QUhO28+RPmo9r4rkFgKZG+QlGLODurSwFZ9Yqa2+gQSZjR
oBEA1ndL7sDFtvkpfHtBZ67EMj0THGBmls4PzBnSxBU7a7Kns++3dEe4q4H4JvzZ
Z7UL5h75qeIpMvcbiaIcAHj2js33dYwJ9HgIvR5fECPrpBrNDb6AJAjnqjCsNalH
jDjPS+Gw01VHiR+4jkJ8BAUdELBZaaSyJ/Dzzz1TBir/DYKPmuAI1Fb2cC5dhxZa
V2Fw5DAlf52XS3WG+yKpox6tlXkACBtgPqLipvdx8uk42wPXfLfCQNOAl0sd3Rew
oHhQ/fJE6cmVXdfYB8DyySp31y0ZnbenkjmV/Q6uhqsx6P8k04PjAilLEGgAw3Ag
QF5ktMuLpSubtG85ut/uaZhELKd+Q8zHqpfen0ErBuIfc1vGrS6Xln3+mp5I6eFK
KJAhw/qdXPdRdNzH9bKZqvORcl/K+u8pOMb/swdQuP00F8bLD+ASmzOwOcWANEIR
e7/K8aRF3zsD5nnwSoQwfOIqEc83+PKEBJgti76Y4CyMiT8aFDLgpyrgmZVaO4nE
QJJpGdmP6uu28tEbohVV8JS45YEjU96KRPaKa/l6+SBbPSkArP/3+6eG1I8XqA3T
1TKk7Sf0buhKGJxt2aVw7KzmWObzj/op4E2etyFxACbvk3ZXWninFwjOgDwG3tQj
GoOuzel6IniTqdqWWx1GNCPwTKSND3BguZxm3MYX/2lOadvtNZWK5AnFPKKHQQx7
j203smeDpIgqJrw6li4AyRTHfC7B4cPgwtPEsKbjWN+dmbUIT/aGpVwawToe7kAN
h+sGgOT4WvBxPTWc10We3JddExABN7H2dkTjqbE3L+FuWVi1UvQtvKICPbDAw0G1
z46MJp9O5mOoMgtAHj9DrgnBTX+q+AzoRgjWtjoGkC3hYd1+By1WNgTegfUAShGo
w7dD3LOp2v5cb4eNiEx3GfKQ/tPT2MnaeOtHuAyWARWvGlf8rWXmV5aRumnimAO3
Q7kHdXcjIQDmFa4ltjO+3YpRAclPEwL52fag5hT7NVRjh/VuXVqR+bpk9kfeaomU
PPn2DTRGGM4e+D6MRo00cKU6c0sRLZ9XcND/sW560l/rTC8m+wyUMOIcLL8Rl8fH
1vu5mHjNZboUwu3WbEVFHhNBRrtEL4kExmr90YHqBjBEm1C/bHVGh8H+i9cKM6HP
AuHY+pXQTCFkFE1XgxS6SNvl+zftg/3z1eBzFCpP3Rx+JYaegFVbrhiyDXgdV5wL
il6tSpZlfe42nh1Bkb9XC2SiaTg1d0hNF8Dh+JGXy9h010nMGGuusirsr6/sh3cV
BtcEz8a51ImAYvDWlFEVmLHQF1m34GPIJ05HId8kL0zl+vv2Pos/Q2Zg4HB9Z7gP
i/EEQlNn9tjHawd2NFpd9wIGeyqmDmPYMARdaQKiYWumYeR4h6F2wNggrRPGOMob
IF3DGC6K3aSClWMrIkeEHTzhDi7x2kJQjicK/Hjn75oASgYWgzkV6gWZZ+9+4yve
4B7azrWQbJkB8RXjk+6Bb8p63XFhMbnMSv2S5jNV/LSPXQMrZZoOKaNmI58QCmiJ
1vYNWBjNKbIFbttigZoKreGScI7IWQYKXfTaMwVtbPERJFMZ5g9L4ey03uT5Zv8V
F16nU3YluN3Cal0ippuFRAt7JdsxFlw//aFM5mW8FtA4k6SONOZ90o1lAGp60BeH
e2peaD81wr7cprYwjoKoDJZdbDR4Ag3rlR+h7sobnEfpJjuFFHtI5kzFxzod5LMv
snFV6V5n845UQS0+a/q7LAqVvR9HR5r6j/OECCznFE/0e2rT/C7Pj6QoNPznROtk
Mbf9MwNNxw3IG9ofVE0skXT97vOYppvomGAQxWk/l2/0cGgXHHMpnNOqjAe1Qv+B
hu+QGvCpV9b087xVhpJGCJurGKaRv8RQy7g/S1B8aUXmIAJ5pqoNMmtgtIHX5LjW
gAOnxKcNx30qmGQsIL/FNJCuwa+C4VdDE3KYh34YpdCSgLTHdL5eN4hjbutlDK8e
9mOABBOAKFX7CoTlWTGI6kWV6krd4WY3WsQPqD5N04AwEHNQdnDw+GxTIaiba9vV
IlBtc+vgFIY7Txd1+KInRO1QmFsURMNgWBBXc5r77ZlznjoCSPUtOM6GBcsD2OQW
H5Ir6jZO/nmFnUd23x+tTs52tdjmzt47EWT6i0PDzqwLEBU9UqEh+0HXiM9mOhBw
VPiRGbDNTU0Pr0U6buea7NiXRi0Ve70VcjqVj+ZVuEk46ShF89Y7MQp+Jbr28Vio
din8IoAnXlIyUKArhSS8Ak0Tz5HIEme7oAaPft2u7MG9gz6l1BFGXfHHM1tCIf/J
JjdCjl3Ar+CmloBN1paOFwouacI+Etew1WvwrzsJxSxaVabpTDcgy6CWyM+YacTl
r82BgOBlJ5WV1jHTUGXc7uTf9PWS5JSRx2VoLvDk1zORD2Hv8aM52QUvSa+0k1rl
lzWeZgenKT2uEDgKb1+f5RiUMRLsGELibHZeZh8BIXVkfe0pvuvNHfK0u1KtJCQy
rjsuZiuepwn0KtHXV0wCD/N+M/m6vG48GcxCUuDuu6oGhi2vYPCkour61ZtrRI+J
JTaUeHKgkT4LgMZ7qKjbNZpLSoXBB99Tvjkual8K4gGhaABY2X2qigFEG/fhq2OV
9HoOfgWISfQe9LlsCJYFrdNaeCv2wMWx9trd8GVGvNcckkxMbYoylTFu1tCZ6tb3
QXg/+GI1QfQGBLE+JQV04vp/1LFJf/29M/jGrxkrwkbmKBtFTC0Lal+Fe74o9rHD
WMI7yF6o/T1iZ3ubzkYhAwXoOQOs60wVJvvUX3XYRvQ1Y8v6Kzx1X7PWdqEjySfv
P/FhdKlpE8qQOoJvsBvmY5lyZHzf4hjh7sGgf5ZQTzSflyc92RJn9FS3PUCA8zwX
0cNVkCiXTABat5Kpt5t+qqufX6NxZNpZqSqjNECy81K+9R4IWvu7zuLOY4pyDgz4
BOHPLTDO32A5ct4U+7SwsoFkpvzV0eJpIgJj1ayu7h6ZE4h7cZr+lKViL9Y8d/n2
GUyxjmXHk1Q3TemDTS5xWV4iQ7DSFcRvI7JhoOUgxcQn03C3RLYV7k9zOTAABCGd
Jm1afK4dqkgxLpj35zFyF83YG9N/nZjtoeqZ7AmtepI1fMKRDkKS5c/lFtEsTxSj
1CvqJ/EWOpPhF6H8awMHMh4wwe4k4f3uybSze/ZzYsN2m6cvG4j8zHJDnUbKOUGQ
BlAIuopAfu7wmkI3l1GwtziN78E3wH5I4NoNYq7+kK1En3G0Tex9x4WF2ETCUTa8
UVhbIhBZXoIaWmTQ69NuJXi/YbXQfYEnQpvhKY5R2mDq8EDk/PaFQdzMvolNEexU
3GMgnE0RQp847ga0Elz7S7tYmhWgC3tmuLHd+r9ats1JlIfHByT7wcNYblWE5BUE
Irb1V4Er4nczALSD4lUXq3tPKZPyvSV0mkNbM95Kd4WqwUSta71kReFscfflabrH
ZjhWkjtBjaGxK8mnJznsWEBvFU76BlG0/i4D8eEqtEc8n8kdEdKoNiETui4pIQ3B
WYaHrO1a4JLBFgAm8tJ1bO+lno3lVLy4nPihL+7c78FaRsUJvF+6aBfW+EbVMRoP
VYFuYDsZUKcMcQSiaSHHuLEKJ6VQ20vqlOPD1Upm7Rn6le26C1Ytxn73jJ1TTMRu
qHrigZ4kJeCor1r1FOB83P1xTywrotnjq7cZ0qIGI8DCSSeBPv8ywgvjONeiISxL
4DpJgxf4i9/pK58ICMSlxD0PenMKBwisnIzrbQPCUTgR/P2VwdHx40+q4Lc3Zo5M
4Sn0E8oFaf6P4kN6Umm6Hv1R1IfW9E9Bp1BA3Bk0sPK+bkmVRRf+SbQx9Z94DEJg
73nY4RsWSV7JftiyVizyGdiepMlaNPIP7O0Nh3urPZAyTnBO+XDTT6FmeoUO3uUL
PtRnrmEjVxeWEodAqYnizFoTW2kXvKiK05cZMKG4NgEJhmDhMLogUt/74fSznfjC
EuBFBd8FR9eDyyr1T2qsls2ZT2JUL/gDPwuVYVdEF7id6Mz53iMAKK/c8qf9Uxqs
gWqA6DN2zq+OS+A6Qa12XTB673oUd1h7e9wAEVJtNp+J02QNWnwsOLdFISedLrR9
gpfV+P6AvqAEX0/Mrxwg/IFJxjsiBrzl0ieL0Yp7KOIRgTbqFJO5cVKKHfEAub9x
XenRI8941Z0jZCNdewUkxqDjjHxxXPDUlK6SYdNc4SpCnhnB6sDwaAqXp1sIaOi8
3TXev+mMBz9biYkJOITfV09VQK2rX8Z1rRale7u1pwsPGTgHrsdtPFuU3TVcwR5R
CfueODqUWLG8OPHJ9xatci5oZs61oKzWX6mFySvP/VYyzpCRuGfZ+jG/DV861iXV
yf3PgXAeMuNiX7bPXk3y0bF3uu+lUwOgB5yt1maXwuKIbLk6S4+UCSGi/uZvP8PF
WLnLAV7w60A1iiVp5M49wd01mLpszvJ0UHlGpXGRUd+u6f3qGmEXOdGMLjKIew2g
5GSmTuVwPZpnhGRg0YWN/7WjqoVNzGLTFEaVTSR6AW5zzqMgEMYDvWZv5WisRTBi
WZ80dCtca+VzKYmOcOVedgF3GDYkB6n6xiFKFFG6Ol2TDOwglDPXaCF4Y1xN/wYt
B8TCe8WZK3eQne9aQxm6HVl3pmCB8WJPVBHHBEAJ6HHmXY1TaGLXU1q5Z4HJIQ3o
GnOMs1RlnVqyKFKw/1pWHQse7t2kxYtG/HlpUFnakQWkA6OPmYn4b5SHaAdv/WOy
sGZ0u56p8k3b39bHeQHlDYoYVINTJ0poPzYEiGSeIU8qvy1LJy8mztAdqfS6a+Yw
cD7BXdNFQ2Qu9H3a0AQnjzxHGW/nGT6NEF8u2Q5sBzlSuvnRHcqUapKHGqkOn3lS
Qz+tZC3fuYpKuQypn4Xafn4kkPnGiONJwQRqJt5ho38aks6RgniCNI6YCYR9Qr5t
45Ren6+bw3c4r6YX7m5qN+f41HvViF26GGM6Ssm4Y0bajVuIIT5QD/lzbGndDG9N
3D49oRY67cVl8IqB/OopkoQ8o5rZEukMVwWYjhQBSwyqfbz9OPHu7lmlaVFdlNJu
2V0+w/S4iZdXYOLatKlreKqJ0spCZg6lD0WjlR/n3/77YiGadMC/UIXK1uk60iG7
Ahrj1JDNzfgfgq+Ovm9RG7Upnl9/NnonZecc3MIbzeIvetQ5N3HsNxh6OD3iEa8d
vpIMYdRG27q5ZhosBha+CUIn7/Roredr0CY89cvbTSPlHaqCTyeB9uzPprF4bqqn
13nVS/lg1kyZeikWz8WOBainyn3kza10fjGq4riN2lhWu2/+kub/Zge07qsXw+47
nWJxi7crU87t8/nRD0oZkrZTAXQuYGTTV957qItng6d8ThznSpYZEFuXKomfvQI0
WjmHoHxM5jb7KXDDMIN5Hmi95HzyvepUVmX2gsH6xBpc9URnxXWPDjh9URkpHVd5
p4yJ26x4nJuLu3bb0EX2HDRDSPmWel9vUv6gprS5CinldXDPlrB3vj/Iev8VmU/d
fLK1ZweZqK7ugEsHdEpxNONu/x9Yx913sHrFcYlECuiYWmrk/4cPSg4cO6w2ajoK
+fBTnj/VLWO0YPJeFOtpHy/rojGrRawDUfbYf6QKpqMe1ZDCikLGNT7XOnrSD+Go
Nrr/XmcYwxrweOf2nSIR1WcBHwWofsZotFOv/u/wIIRDtrMUTko2d06C/shO6omf
Vfl1hBW3Su15J8DrV7E9cnM0FvDqoTzYLlrm8Gk4HjIYplSHHlkOhifhqY45alxI
wv3m06jiEtHUq4T3zH7d/dQav2sAK7OmBKUjtMzeXK8e6COhM+ui3wNSWlqkYp59
BlgrpDDXKHXk2Sz6tMBplbmT9xRQnSN1AbJamneVZVWChZut0LkMbDrGHGd1bOXa
TH2PoxBjmUagYbWq22uQk5UWIRgtH2AjDUNoqnmhw8Vsnr3E04Iq05wDjrl5wBS4
l75qnFzkC5CWkptkEol+fzqcEIqhqDgTg5YMzdhgAQKhGtPTWXrsgrlHRUCd68na
srLcdy1RSKROoUefOoIkoeuOZouqPQIdBIujIHOG333DTxCChmQ5dd2vo8V29053
O8+uhFPdscuL57Lgf830xEzZJU0a3F7Rq/kgMOm+gyjcXQItBSAg5WjmZhxT83Jz
/vDAENTubUm/BR1jIpo632CkHPzH5zRwzb00s/ZUU5fjAZJ7Q2PoroCCAHBJmbd6
N0ns/5/JaHKqmvoQnwJ9X0kvH0YKhJmmJYLo/QPw4fVoNNloJW/rg25jIHeqzBdt
of8hjcQsJluuZY9nyQKocBi/Ox2DmigI8QWtehooR729DaLOBdHb/zUlJMKMsucS
o6yihQzKUfu59UaQQ/jIOvI4XDv6y0cQUzegkgXrbuLW3pp3a/bOJkghT4VyXLrY
dcEj6V7ZJZaG5GroD5FrFclDeum9kxb6rLOdklAKmcfXVY4hBlb37c50NoM2LG9O
JJqbwGbom21QFLzJ4WbtLH+dyL3cz9ACup/JzyIDnu8ttUSql5icfxxzjVS/RQOW
uNcU29o+0C9x2S/ZdkzxiKdwIzlNmOtk2U5pSSltboYH8vh504Lugh8kpzXClpUh
74Ar1IDChcSJoZ4I5bkzR3yDxUHUy5MyQLJ7A4pbx0PQ2vrUZrm6nzcRtXVha91H
hE/skKZtjXqB+tjlgUfagUtvF6i+dXAXMZkz/55y6dKJU98CbhpH8LoE+qExyp1U
QERnsk80G0GjX5I6mG1DHAHYBQnT85oUeQOsB8b2u0uoHBsVdj95LvQQCwFIc+29
SROx1gvyT++bCkg402kOLXDzgP+0FbJAzG9YzNWphWPQl0y4RrBC2Hi+5RuAwgEF
fJoedNhR2DemliOtUDakXBfuSQPHLs3HS12CKsMRc+0yIm2fNWCxIUjKZhZYYABk
9xJthRl50D3Fs0LHL4SdcERxB+N/4s07s07Vr0ja8g23WRfyoZvORJOqYwPWJwNq
Svdd6MqgzzdUdC0ZusiF25K8XFwyI1EeoXPLKC5eNbQzDUcKJtuNAGXka2iQoGZP
PjHtCKkQbQ8llKVK1IAgESjkyDz2+ry1MN+yON0g0fOKuooZrlA4ZdN+0xN3xF+M
h6fQASMy+rTGVcvJXDTU78fmqseJEjTwhJKLmcsoJIoQAEh4oZT1eZ7CZOuKDaSh
AF2xGds47pFrNxEgmj+myGpvRqy1G3EGrd8/vNFJSFb69nwm32eBW0RM4MipyH/n
SE0kIkO4rdMt0gkGJnajvKqbkURTC9h2/XT+K8cs6e0oefpBi+h6h4j7P+Q2JN4R
c3LRYLcQ4ZvgdRTiegv2j6TzC7KuOHRQ4HbflO97+Z9YlZufGpvogSdbap15ZiIS
MiWyUxEIsjgUX89NWP5tY5msTP0B6sMCJdbemUf4kYEg6vPz/9yt8uMlggqhL9Dg
pLoQ7OGGvj0icxvyFLT8Noca4Bn1In6gswXJjX/6NwKdi7VGRLfybh4a1NQ0a1r5
gFL0vHHKDI3GQW/j936AIcI7GPTGla9OSK9zd4xOB1ZdwlMH/Fug7eRgbIzGdv1n
4uBl8PnPEf2WR9oi7+ZVwoN9DoLC2w0ri8cQ+Ak+ZWk984OZASX/OTWLPPoQeni9
iv8xs1F1+1f+VSQCdV+SOWVJURUNjbAguFlVMnGx6zhw2diKVt6ddrDP3Kyrk0F6
Pj/HI+3s8us50nvUhsiU4PR61lPWREdd7IN2Kc/hLRY/nwzVY8Cox7A/QTDiIfgh
alA3BkgnpdIeiAxoOiHs5bs5ILcI3iIrS12fto6E4pZi2UwLer4QfBsr+gS7eW4I
Y3blxvN7LsNfCVdfYEZcYQZxl7X8t/l+axk36IJiEyq7wqZmpMcBpVNwpTaJ5qL2
ta/v6B+fF5PSjVL3UVs3T69zQ2G0q1B+lXUmGzG2BQz0PLryyG8ZomH9GPB8DG16
xI3rh7MZ22VEvM0QiikOgDZO7tTMRV9kwxsbUW0A04ObZeiVXAbakhkFFdxEFYZu
yJiqRFcwVUJ0zMSW6wNhd8ZqbHVOmSNV0tq5qrCM5o9wIA4A3mLf/V0myaxR3L18
JN0/n/piX6xA9WPetLFczzPuFbFYcyqcqewpxThH2ag8lC5ZdciTL+yG/t7g4fVv
J+KRaXtIOM1tVUtQ8mqrJmop5c0dPGV1/YOoxbyk6X2cQpOyirNU/te8FTkFDPjt
sXvqdxBdXsnP+YI4ZVaMl1TuDF1z8KIv6lHvJPfYdCDQi/oVhFkbj4bBDe9wyA4Q
B9yYfWxvhQ5VMJTtSv+60vLhlpYTOA9dlG1hqfuV8FgMg6OHLnfqvHoxuawiJ8F6
Q1oa2/5eXitjQIi7Zcw2PcxZaLEZXkVBrurBKH/NsOlVf5qvQEexooUok2RztZmV
J7RyJeaBTuDGAnHGeNtWkJtAILlus0l2K3qkK/UG3iTx/h4u0jJX0qJJSxfAQk8e
1uKYMg+h4EKDdQB/TmJ/kbAXOX+Rr0bkjPA5fUBOu4//cdV4euwr+3oATGI0tL2u
XUTW9FlqZNcBPQRr1idw28eZdMtdkwz/sa/Ps3v/H3Gof8rQRxrdO637Gxu5DT68
/RUsMRcFl3Vd8P73lepmoVUJ1f4juzBdt69XdxKnau0Duv7OCiLTfecy2GNj0L8f
9q79JHZzUlFE0fRSoIq6v7El6kl3oG+lqaU5I8r/u0gJ8z9vGifLFBA0zDSgOB3m
YktTxzxoVJGvIOvU2T5eD6KDWV0jhhZP3My6WI64FUIYVGMY/pYLhlt/uBzvNkXw
vCYbNxTiVdYJMuERDS792gTC91+iHun5gwXiAt8atNlY3b+CKG+TVaIlrFjI2ZeA
31DxMn+I8TzxcKNOVcdV9UjoLoCQ54jDjFHIHULtOZOK6LfFO4RYxfRuDUnWvCR2
fMZmRfbJEg58DbHfRVMAvf5ElTRynVgJ1Qo/mCCgG1qk7QiCuB6RSfRCLooNeyiO
Ih/DjRnhDvkwwnxtT+SmL6f6gdD8y56rQT6kWfEBmMrKhDk2XFxoIHH1zdeEMgSb
BDmg2PoDmHkImStdeS0YQ9PL0N7fEE0LECkiqxoXv9A+RcOnPCK+yuKcKzXBEdZ8
sf4IpDvWrdwGBDYTiWTQnkfwoIt/D0+N8QAmO5e0TV6J1weIgEmJnb6RfglbfigR
0tDpXQ3Fsq0PIwzsjJR/SSlTtWEroEG2mCEuyEyqnZNchSREOUL6slAYsBzKggox
83s34Knr9Z7UtsXilibuEWNJ5Phk7s7Ac9G22pEYY7gd0MHOuCRb6fpzyzjyC+VP
wUzHPOM1vJRAKt43emCvdYF1MaVu2c+spZ5IaAxCWxYo3S51pIU8WMQ32rCu3HtO
xaqV1svd9XgAjfmzHcD0og9tdcjQq3xRSUfyKOlH6VxWYgxSYLHi4lvac85foJhA
fhCEcOGodb43wojpRD2V+rHqHAW3ylFHbliHK3TuJc+OssZattAoAeTVuRYTh8RX
F5KereAH/PArWcEDTrW4aIX9L8PDrb85pdNlj2XNB6KJtGCz+s8Q77PHvMe/6uqB
Q0AfHrhVyWH1ZbULRKU86eaurxf/37EeBFSH5M4aYIs7BxJH7Ziaejvt6XNi5Xwz
qm8FaBDu3HPC1lSKUrd6gry8qMdt8eD5GOMqxBJpkJej65CN49ZllaFTBt7B7UFo
IqmBCAVbV9B4C4ashMYjbtNb2UtRZV+RdIWOkjDWyTmZNhQO5aiNkJkYdQKT9fS4
T1BtuDnGN91QFcv13DdzjDfGBY1uBhvKJPqc41RtJw8IQPzLSdIeApVVwvuTzxkQ
25KoQ2dTvxENxHao0qWWYc8LX/oRI22h8WmVVMTU6mhRuTyqd9ExwEcm05QMrTb3
/ttzPVtG0+VneRJUCtDww22ncktvM5KBoUO47c+6IR7GLDOUxm+ETNalCxRwFg5p
Q0LlzvnryJ9TugjAE8d7/lMBT8EOCzIS5x9A0QU+tZxOf3vJin+nk0AxhkrcQnnZ
xD8e1APQjDzaxMuPwLD9+GJNkc7Ef6z+s4UgG8zVVJpGCcJglUfeGfXeIKutN1Um
ND4NES0XYptcjYR5us2n8Zss76pUEoQGEST8XueJ8ZpppA5Mjt5i5ylyfAsve87E
TtB/CbdNtKSWBYIjgDU4+CDqIUpGuZlEf+1leTXdLziMm0kczcD8HePNSrvkRhn1
DDB9meTRvJc/6iCj18GEyyvpEclQlxuYQhHnASoW1UUYZhUYAb83XRCB0Uq/UGZc
zbTTlgS+VNBwEentRt+UyyaurjMdzT4cEfHl1C6rXCwMgB83XW/rAi7R6zST35AO
/EEulHvJqZKFOyOuS6jbVUzzrhEOHPxzVcETCratRXy7XPdHEFxNkV0Yjka4POgE
cvM8ApoMMjH/iNDL4lQLi87C0G8o3V07hUsWXjQT7QzvDYMJJeBRzlio6uUb4ohP
KZz5jzsXq+dJ8gaClxQEYfa0nQB1WKggW+yOIJ+FEd8P258NTHk8KbMgcrmLSvSc
ZhW9M0hSWiKTCqqWKNSZv0znmn4EmKJNoJccwlpj25/5V+DuXMwG0chOKSdyNqZ8
mgX5sU+e+efjYgMo0meOYl8TGE4qP1gVXTNbmjQ+LhxEQB84jXmfGWg94xT1b4gF
kcU0W2arNH2ND11J073I76FWC2Hz6f7YUJPwH33O8r1zVAcreZOLeFMMiZ2uFLls
wZjHY6Piyy3M4U+o0m67X064bv2RuUNB37Pwoot/lM0n6SIs5UrVM+mhYsJRvTkA
VwwiS7JDHSYSJlE+u/Z1xVT6DYmR0MxqtJG/JIAZ9O2av67bFc/QsK1ehptQx8oN
fb01tE3Vdvu4wLk1LeRpmmXPTX4YBTgh35EelDRBr76gpDHSYdp/K4/ZSJ0XJGIr
npqB1lUUZxtBGiUZu1P2J+XitVJPYrxOgiG9QZnivI7kbcxGjPWdn+khZ+g002ip
CFUrp/hDbIu9nCOZQ9BrTgEcXrkTnL9jRk0dWo4Ljrrtb/CivuQoYkPRase4BhJq
3uwr3nt/+IYWDulVOQjNGPLH09OgCPfUL8P/Q/gIMHtEbtqwXqfd6b3mq5JVoewu
Iyr4MxiCcQCb5QEbqrxFtik0FJUbjPJn7l7SXcu+nplaYUvubrDE9THvusQHK4mU
xIpxNfuI1UJThMMwlxSegFQ62k9cHlDDTXizwTvijQV6AulbJMJTkL8ygIhjAAeI
nrZBOZRGdVllVN1yODD/iaVeWlePjh5oaRnwsnzhYftW5icNEOIwdYSHKdD2FoN2
vDzGs+qe3A495jkkPSHY/WC8D9REGUWrrevpP3ZcfgQBwnPYvxff6BjzCk5ldjAS
wE7GuvM/5NRD92qo2CFqwS9qW9LC8SPJTbWXT/+w9V1WPa+W2hPa4EPbvjTuEX3s
T+j+ZCC6+i2BSNMEDvEToO73ToUseHzo654CIsimIosTnqFO4ak7cp/C8wgE2JrL
D/JjYRQ5khlbeNH+MBpMgupwElsSwyrrjaway8OVcPCgtsmLME/3LLTnBz6uMcfe
7h60f89CGYKj0Ef1YheUyRrJuDdivpOzyFmKCAn16pA/7lljpf8ulNicIsl03+C1
cscmGpm3a/FZ/ig6MTpGmRD3iL8a0NQYdZ+yVVDppARicjMcDq9WpasmktA70NVL
eQmBV4zJW2d8WsacxU8CrVGOdQPoc7PGI/mgJdBQmcmrsxSJLZHxAW1GgYklc+Hc
gfpnGvFrcmrdqKzx767aGy94tptKxYpIXjgvzYryf57fOyggq2u7vgC7qvxYsDXt
XW9TOn4a20w4/lvZSVVccEzfZXoD8xtd9kH4D0d108UpUJZUcmDEUg6nnnBa5hdk
Som4hB5+9lzWGq8/Cy9rHvyRxd9Ew6mkarym1VAsxZLg/npvCvnDzHahMiwnsAny
cnSG+qcqeNlJ885Lyy0FJn1GUWZgt9hu2jWrfd2nuGTQppahOpYTRXYtF8dLlKKd
2WVAABbz++ZNPd3hNZtzeU6yjMR/GaTGRYJat+l2VqZ2yxf9ysuzCmxEGO9HIvw9
6Xl9a7NyIjwawInTKqqfpEm3Gv8W/Ly15BAawsES/RAo1prkMSr6/1WIkIaKHt7g
BenZs2EYiDhR0DSsb80LoCpvlP3/R0DZY+hFyw4ywoIfKsZRt/z9mZZ5kQSf0MgS
PsTbJGOHyxORu/2Y/0EwptafjmCAXJxzitrfDdRBs/6cnf4ddbJBamaoUyVlRGQX
sxb91tWOJR5SU8PBzWO6UR3aGGROaeclQAVV3zSH9U9cQWhJXjiel/Axn5UjS8KP
AT7cgmPVI0NQE5i4IEQsrQKMVA1g3cv2T9GoyciaEK4CeWigqXsbbi2AZDlN4Snk
HTCY0DyclWpcaEAQpXg13N8Nn4Y1EdOxP4YWLTVTv/T1HZ/uJyRo3NVk5d31ssio
zTvHrhYfQAdH82RUZHB7wP0vWt1wFnrAguXhFWx+zcJLMUnkZZ3+m1vZioeXbNQ/
DvR9VPomBYprdCRqyt3Y6HotUv3YUu6hwQJbO0Ysck0+yxm/ogrAXLeP15WpPjbz
qg6U26ZvylBWIlIerYIoiLDTAv4MzBi1jEdLOngcWn7fp+BVsGXGMhcf4ILIRPQj
Io9qKg0OVbkxpJjDR4IeTVKs9o/qjgFTCKogScUFCybMvQyaDNVKEAy97viaMkUJ
E2eaSHgrESRJ+kephv7peOnW+DgqwYWVc/ewWPhjMWQgK9AkC4q0nOhjAR3fiOGG
2BgAI7zxbkeOLYS4BcIkXTj9nKGF3OyO1suusmZgRfEDwusqkkfUb2X9z/JF/FeJ
HOfr/SHq1rq4hWNgVtSeHVJQbBCl4TyUgkaDFbbPTGuh/R/U3Xbgy6r0JlYTbbs1
eKLsd7SfrgVL8SllcYA4+V+iBQ2nlOoiBRYChHtFTgAEPm5tJHdB0wANYppHEaxz
QxurRKZBlGOwEuyX/H9GGYVWXUxb5g7ucJxk8RAgm4yAE1jTplANqM20MNwmeJTp
4MncOsk4k9U8dCqrRQsoheJgCPqMLpTrc79WGkqYHShiHTNdjxU004GaIinAUC+r
pVvR3oiHxiwMeI2DutoIgNUqdaXmEeqqmPoE39ZryDaXUwXjqF5Oq4g0rqHKKmVk
xp236Ohh8hMn3XwoG7aHk2GsrzJ/5KW9ewDRaA6JyFvHC7F3POQLuY/T3q9U/SE4
hocUp4uQMLsy5BDdoXdDz1pzNdaY8QFZdX6Z3amNne80b+iI41SVutRs+3K7kdzw
JOKmo16NcIJ9MMWfMc2bUffq1l0kHZzeucvmp/qx2q4OjBahI3cd2RdVknHM+oD8
Qok0U05EWgM1kgj+r6lCTVyAFRDeUmFi8m4MJyjC+3ptQ+HVriJJvd/IJjyNSCh2
iU1xadqMTzhDKsxWE32xLHPaaG0ygzzb7kyfRKHIpJfI4I/G+AGt3ZC7ZTkjHxXf
W4AUpq3O4PHVFztadXoO6aHcir1GYNtO5xujb+fcVTtQyo4P55nf4Ts/fdCN61Pp
QhzcaJHxcsIHu5xQDZKKCwCVvhxOnn7WkNHYynz/JWSPkOUFmaW37L2hegG1Cvtl
xExZtUm2W/iArZZfBPd15hDffFDmi3aQItkxiNXVtGygyH9CeX1V7vxFPVXOUm+i
QwKl5hQBnV2qjLS47X9h8T4m/yJ6exnAHMTeKs8mRuWrjooFq8RlTE4ep5roGSBj
nNkJCnlTsQjTjou24ak19MOeXIfzD2OhgU3uk9npqLL+DrksSv1fusgpvRif/cSp
QaptjygQZO8SWThmcQpgzzfOmFVyaq4zo58vOlYYO7sHXHtg5LwmDJxgisSsbC4I
a69jFrkqEcyUAAsTiUEKlmwjquNXvyLg+glrA+6MbAzf3txSI0Im+GPCbjxWoHyD
Few7P0HD574/9tr+VmOQgH+Ml2NeHl+ku5ZkOAyCbWUJN3vRvmHegvTOcIrRiOgl
1VfRXzaQsN4nVcLCK1S26QKSA7nUxmKdMoyoHyt9qzt8oW5mRsadAaVuXD7P1F9P
KrIXaREsdjr16+xU4QgMFcptXQ/NNmgphkEAOrdVYYOd+8dFVJzgDsJ98ymiv7ft
nPIScbtvSzQ0C+zmRlo5vmUppKhy69A5FsUoU4wNNNRZLDr6e9Rhfi9X8hLP4VvC
lAnXNGMOyWW0h4x1SvNq4+A7TBbb/n+r+zURmTZc+6+L2ZPwAwgRPAmN7AYhzCNi
ARtItnmPxH7s1/GWCOnIMCR2M7xkAx+pC+8GKnLqXCbwbLlp9SFWFKPffqa+4Ndq
PX/oX7TnttbQebwgV1HjczTxLfluxLLuVUHrcT70F2lF3YyjdezapwljFDVvadH7
vlzBY8FWgPrC4X/KF6nwITYnLXcGYLaXuSd74T5IyAq2iW/6iN8HutTSckP7F5gr
KiMeCqsref3KwME21X0k7nu2xilfBxPh8Fp0DkljNoCoN6uhrmdy8nkLdUJN/o1e
WaJDp8L0fi9aGL3vmi20Xllx2FJpHRXwsHNJp9lVMqmG94EhGgqM04z+ew7jzx/Y
iOPuwMxf3dMwDQe9W2jALHKX2BEDOzz4Es4Mj/AgR4GMuDrTcNbIP/syXdwBfbDz
z42VucKqib4CibmglBDEnGCmBIwgEk8py1bRCJDWqQFw6FTJnlVt3rrqTW2pJ29Q
2jkld0fdv2UE42+xH258JKErtOaeGr/nhYN0FyBwUxSRIkHG+eIAxe6Q85eN06kP
umrrDaV4t3Ixs4e+b6uFqJL01lmE/lKDCORUdzEUGS6ICjf523TCQROdMWLGOHzf
A4yxYyMvIDmuMnLa6BxfVwxKrIy2VgNcOLWk9av6CiP8bk6J0SBDvjmC4RR9FFqQ
LNicxCh2YV8mYn6SAMUiFybbPOay0svluTEM1zFwOy10X/RZSX0ZrvgxNauT6fxu
nN+pH5fC9+cOf6RJjaSsVJd2e9xB+hIWd7/MFxqgiuzOsBM94QXrVpgn7/+6Rd0p
/hnDKl1WAvnpLLRGyUsTl4rARPg6CEpe/kUxBv7rUq9YdaLONMcUhTmodmHui4ZJ
OVnzhExGIy+JzS2YLnxhxhivHFLfd44fCWcbGOaQ2gwveMK0a74Q+H4dlxD4pz+i
uiDEjVlknxQBw2uqw7ZiO0DY6qWDQ50JW9bDo+1kPWyYQveJX2syUoL+DXuA3AGu
FYeu0CMRE7xsNZ4mcIaj+4jUoue0P9juDsDzTwsfisyQYD/kii5XqdXYvATb55Ed
mfH7BZLi2V1LQaq73D67myTvxgcpUYg2DLtU+phUJ70Rcw7fmroMvjSfUxFCx92J
fpvT9Vsz/7IdFoT3lK52qHTllSAFhIz/oDzejcNukXpPBBWAaYcmcOtylOIX60wL
FWYxfzpStWjYX3XU2TylYBETGRqprwQOinoMdH5USXMJcCKyxKo6xKg5uNUi6PjU
tqYw8srbJa5j+r0TgIcg5dT3+X793uSW5TTy5At841Ux3zo9Hkc8rtvzx62aNxHE
ya/ixn34a1nqtdYo5CU0PJ7khm4G1CyQ3CMGyMpVvB577F3xl9eh0R2K1xtZ9+9y
qUsqXDR6CD5BwPtWXtoVFTKGzCHAADTcwMN04amdeVbo8TEu8jCE6mwBEw6j6DTK
PYXjFuimBr8j1oive1ZU8LnxlrZ4sUchhz+mIrcWAkIJMZNYOWdU2imC45iF755t
GkEiqpYdFG4x1Gfvq1Kx8ahY3cs/qoz8pGkcNn8t7pjVCBH+yzvCS90ITph2lb51
c7cbEXi3fTp5jujhoZ/IPfGYniPNkoBBlUKom92p9VVjnGL4vtu2/9dn9X5WvYFr
iA46j2Vo5UhJBMo1f++OU9sd2EQ7jjGTziIUN22e+nqfviy2DxnogDUz0SPE0Tpz
PiSIyVdd9mTMk6KCD0G4oP1d8jTG0XlbkgjYsCKpIlCwNpYdNKQ6odm9wXWqpndw
oCpW4Gx905/EF2O2+NkKRDJMGq4Q5rDdko0tada6epyhzUCdXuAa9gKP90FtoB6W
JhPE1GCp7Zq+g1a1oTlKLUY4oa0qbF2nfQ8HhjmpZIoeeZ5YQyzJcCvupb3XHONw
aQC5EvDPwwqyNvBeApYs+2fxehDkA0XWw44DbdSPgxDi7yayno6gFeQ7wtRw13qW
XCjOnkAfTAZg5zLuPwKmAnn/B2sndUPTvaAvNwdME9U7gv6hPqR8jqRcoX9J6+Rv
J8IA0jJv0XmV9X2aK3NsmztdK2eIO7g8bOiCz44TYFZtir+jRmMkODw4vT1A4j8/
G3hv5anHzL8GBABREv0ejucBN+LB5NMMuNK7Kx/DN6Zh4ZvOAg+QV0d50iAjg3d7
LEoovkhwJsU9+xBcgAPiK66ETzsOoeSuuveMLp+0sOQokAHgTuEKi7OB8FOb3KY4
+CCFnJvRwR70cWkp3NeUSu6tX3gHR5m4W9IInJMLYg4DO1VE50QJYxlgkuKHv7xz
soQRilQMSio2e63ex/bDJGm1vWpRCsTiL6uFg4AOPeSVIHO+DWopiMGB1Isvk+Cf
sCX4PeIaWM5ZuJuuQNjitV59jdvJyr1XBFpsHL0tqVo4xbx588jer/ov782309Pt
mGBsTLxsFoPqS65wdhCfpdCv7E5shDe02EHwaRRtGRJOKQNn3c4fP4w8F1uFVok7
6suAeMc7bR26cp7+f6XYR6JtiFEZzHz2Mfuw4rqOhT8AE91uRIAvyqtSlSxKqTPG
e9FR2S72kLNl9JlLVoEpa7CSEI1v84xdzQcUP/0qAZEOZOE3DDjA/K1ZgcJUf708
ogMgCIFLJydlldpJ+ZGquPibOp8D7yMmdyrKL0R6s0/lPt2V4XJo3KjfXC0fY8/f
eGV4BlkOTiclRzXWhNK1Q5LDmTmsg96UF3Ty6fnSIYIwSkv5MgJeMkejFIL+iQhS
74Hmbb1ROfrs+9MWye1RI2OtPC/LqJXzga75FAtYwSYG88yFewYdTfPnCID2Whca
ZZqjPl3uLJ+FZZxBZMlvulfIxDLqtXkwSNOntV5UBx9SBQjMtnCfpLL2lRR35amL
+ooBcqNGco/iXkDiV2WqzFtqnVl0KgIDtazZro43px/s6xPKuBurPr80UMzYpKz5
h4yVy4I5d7p2YQlfgxmPXmx6Hzj/2/X5OgNyETMojoIQT1DDMBsFFubudYUQ61iH
Dhr2p+CaatLudrOqQs38vaWW8I2Cb0e1uBkLp4rQofi2gDCkqJCX4P4PhlzionhA
lisW5Akzdl7DAaRwGwfZNCUGcdmGEYNP0L66gb5DnST/L5O+ugR1EKnjv4gaANUg
/ICQMTzcGiU6KZhZoyT07koSDkhbaz1mExhEsybE4O7IEqBYczfxwgV3z/ZQfUgs
BpsolkcbHMK8saBth6kXKuzFcfPbFvphgWiUxf5cLXLYPgI2BbPGbnSkvr8Q0dK7
xnPX53g0uNcNuM7Kyq6FfipYMqh8Ahg0KyDXkSEAjFhDRJICSAa9WbcbYt9nmEJE
cGgSkuDhyVQXOTRWYnRCogwHl+RxKEATyjRc/jsIJ35U4FrTlEX3gI4wAnpfrIgp
mdBs+m1cm+t5QqVCaV9F3wubRXLbLoPfUyhXYkBsUsETOuV1h5i3Ic/W008QK7ZE
RvRb/W55ydcpYNKAuYDXxFbI9AO+bWuhBGxav0IvD11qLXGcNGQCSzm8qjnZIox5
u9WdiT1Hj1w2mK+JnUqSOP6YK5CrsaUCXm3I83FUT13n9wPc9ztDpwH1kG2FR3Ir
KOXESffzyogs84FDUTcJuhx7XYHkXUoC2vu4SU+9Qm4Ne5D1nzYN8GCOtaZg2GWt
abN16hlbhQ2gRj3WKAI14kgVySGyGaUHbX/fCPB6Fys6eNfrzdcgxnzD0tFopJiL
BXyasWO2xrVGN8SC8RfAupggBnqw6pqxjXH7aA7aS7hlsFoSG1tZRWA7zjaz380f
tIXed4SsjGMZ1t2wQtWrrkSfYP2HShr67lMPNAj/4Cv9j2KOBdbhaxVo5vvocxvR
nthA9+LPV4LHwp4mPo0jRqsdjRHEI/ZE5fNt1r6awNZqtJ2T5IT6HV2TARbuHdqZ
oR7xzp6Prxu9/jGCo9AEUyDJtwhiKnd9hG82q4cK5YzxbXd7fNhDm1VLOFv/0K57
fDrDFcZuVsnlnWbwp1eYCi31ICRL1PaQIrsJ445+goX46VrNn+gqHc4N41oK00s/
6SafuT3pARu99UbS585UPtiGr/EyH4e99aV8xpB+SVt3jxmAxZsngVZE1MiFqPkg
f9r/z7KQZNrcieWsKme0m3DASdIglpJHvGCgm8YbsqtvX1MJSkCknG+on9PLk2qw
3TRqg39Xs8lxs/xhiLF/fygB61PenIVHZZeOnWzvZeKsj5+tZ5dCVoqh5FNx3vgx
h4qKbKo8XSXLWE/Aw1031Ij5SZE96AAC27ZkfigeAQ0W4SiqPWbUt5I7A+dI4UFT
aO14FcHcXTC0eMocpEy4iL4YuvRwLtTX49wogHcaenZv+vkPLbNyAgLi8QxNCfK/
QCEw+VRYVv6NWGQsFlrIUdCW1njM2KH6ME3uk2N93OwUeZPLXmOSkjcy1gNocIl4
dJ4u9Q5DURn7eM0HPmXDwpl/Awt1L38tuliQVIO+t1dixx7ejcrslYaR3kbYlTIj
hK9UkqTJ7KDzOKf+SD3h+fmifs4oklYRk8f2WygmqEX+O87jiG4pzdRXBpxoM7zd
F5/+CduA9RvKeVIGPWDRDVsUy+1ePoIfxUjllIO4sNZ6UYuKIKHkQJhaH9B0p5bN
ch+rsQLuxSAegld/+GquXDH2c0jJACwFQ8zDOluCPle/xwml+q53V4jpzgWwB0xM
RGhXHysU4q3UN67fpkH4VpaHTZ6bwnekx1iOud8JocnrSTzYIb/8VLnkAcD/6HlO
Rg62hesd3qL/nkRGpCp0+ZOZkfu/weBqiIEQzNKWoavbQvErrXJ2CpmNXZVBlG6w
/UiHYnRxXJVGCsyxQ11wC9rkBcIb9X2TcMSc1XplAuVOsMkWrLdRA6F6rCtgJkmD
hw1fMQD9XsL1kXGkLViQCvTZBx/y8PTTRnBjtXC0euDUkUj/6CnyGyPJLCES8vMV
sptkKpMzS63rOXTmGycWdB3O9HqcPPb8NhZxyVzmCcgLwdYiM959t80o5RQRPLUE
HyGqhV+BeNWzt+mvbImV6Cxqk+9tadBb0qUmwsdg3PcIIecXU7UdGh8AQujGTJr7
f0fj4Lm6SKQ42+/5mnUipq9mPsOrjNqw/yBwE88vbgS/wympijqh5+TDgIBSb8jn
4rKaP5J96rG93nwoJ0iy7UIrfbpup6H3A1wA0xwDB1Y7oKJlumNiXWMT4DEfdcV2
PlTKCzakL5dUqJBKWaqRuC6bqPQ23EFh9gZhd++BCv046AmXdRAPnN25vquXGcBI
C9HDPdb9Ov2gd8W+KHZPROAZUVuUVDhF/3DlWd7gByIf8UIQqMyjCfaeyNuHH3rv
Y4JjrBf2TG4MIpEOUasaoUu43YcuYYFd9IiQc9IXv+zDZqJN5oMkZs/5Z0S+ev+I
iKKARwtHucpybIRPezuaaghcWu2mD+nHuuZkvNP1zWCXL5mHX/lM9oTdDTEpA6lG
G+/Lo8K9nEAKyIZrzvkWNxh7PJFM9JiH65VYjKCYKAiF0HuADt/dAT/GX/tW+znb
oS+t3Nxyq+tY+l/fLCtkNJDwy40TwWfiWlBON8jrBt7stbOlOXgx8a4Yx+Y6Ez8k
7bTMdmHYIn/ALjc4tS93E5S/7twJeshAy1xe4SVd0DEYc84cGRBGFV8SNevlvjQ3
YvcSBgNc7409c9qze3fzJLAYVbslnlQkrDPyriUxxnHKCPpEmLeiy9Zs13IaQucR
1UrPnHIskbet6QSR9CmZQ3buJlVrB2Eq8t7Wkp03kp3NPExlvfwdabkHUAXf8YIF
V/v9cgzaVNXuFyuQxTZsnBzQRp+NzC5bRk8HKohYmYI5A++NutYmqNONAUdEHaPg
o+YK8BWEp176ndVVu/51gv/eNNW22yVhFOadqUV8Iov8nZ0EEbaHc4PBpGccyBVf
qY3WT2JCkbDefHRk/xPl6la5c2NfJjXCO9KvhhfSV0kUoaaJMN/c8suApQS8O922
zjanBDBW40y4CN2lqv7O8qR39IPxQxObnu/9cabatakm1NftuxvEJ360yyDS/UUw
LXwidIrgYbm42FNsdBzcc4EL4IJG2zyyTNVv7Bpg67pCAPWeeZqEYVFT66iHzMYu
Nh6x8CO02SkKBalE+RuT8P6m74KxCzS9YywEPRkUcE3VpQY/fXUIG9YKzDJuE/VH
WRcNqT5bNNO4tA8ummAw3yfKHXle4m6VYk38erV/ZzFAvlKvgPEUdgV+bP6Wt7E8
SIFd04qYUprSWMO3QgNDmnx68xKraG57RUUqjnmOOAJyFGTKY+ipHcOVrRWDW6b1
gHGMIEZRuk/ceTlyTjq1cO7a6dBoDaLcRpogZwF9rsJ4AS1l4AICDCT9fu8hXV1c
rRN2wSdMqOFsWkPB8Sg2FJp1e7sVtdtfH7lxLyHy+W4FcZ6xALiGWw9OZIWUbL1u
X+zMd7SUX8A6R4YA/GI8+OkE/POm1qlx5ARfWgxj4EYZL9zbW289TnaUDZVwoPSx
SlW5xtyAD+jv79y/wS3RFUJ+jyCoqybM2vwJev/OXr3F2fShucgcnTz6X2eYzEVl
3BelceECB2EbrIAtSOVWtz13dcu7NLTZocTtS4/NboEPn8j4/nEdk9N+DhQtnvQa
HVGVrvDhc9zgf3WMtwf3PFWZ1oxWtHpJlYV2g45hdb10kHOi+Mc+maFppZphksYE
o1DxFz/NuQfDb4XyfDcXKpQT1SNbrIh8fJoujaMK04jgnalCF7hYIkLW7EEHDCj+
9CeHh8NYUzJextXdpYtSKjDiY0mqy3x3kR1WoytcaS1Dg3mya/vU+r1grk8MUlnG
A2b0W/lmkZ1XNc3HeOL48qZGVG+OjbPDdLyf39aSDXi9Pn9k6KKNXMtz9T6fjVYc
H9Dbe3fWwxvIx5j08Who5eoHMPDR4BeAs1yaekEQnrY9Jo9I9h4Es+Ez3sFWB104
xpdoAoIJwSGv8D4Cncp/T4+iVT25NTCSQtAqSv7wFCzlgccJHx5bzZCuTHTYMYnD
chuRKfTs+76fYS9I1Kphw0YQFmrERtgN2r634uM06TOq4LHkrdj8vzKr7JgCdDG0
fP6UzCweymz7jV2x4R9hR2hA3fcfnEVfMxNsLBGi9V9i3eTLOuF7ypuB8vehVP2u
szHFGRiXAbZ91ZxOCGOY+GFVGFAL1hQcKAoli27FOOu8xmCPwiXMAKjMJn/dH0a6
LQgzpT42RY/BN6PjuAilYTsf+Bzyad2R5HJim6Rvtz55/ZJ4QwuD74EJF7lES5xa
NUrSS18Pc1q+DIg23l6YpdzAulRb3lqVhUQ0Qym+x9FQPXvdvJB/RY01xmWywcNr
7y8MrwujEsET3gf1Y13wUCM1aLuhwEtNU2KRZG6aptfQuizX5vc5BhwpDqAmCjxT
o+79/9/AJSiyX/Kab/MhdYsN+cEoeYDh2lHHTgspfxUcdg3p3RVPCB+uqI3czsh+
t2Oa22mpn5tvL83zOTv431gKxbij/gD3OKNN6y+P88bYNMxd5Dg5AKfBlmfhernM
C5iJTIBAnyUqJhZ8ybcaBkbPrLStQsvyX3UHqONn/ICjdL3er7B46nInjOD7cKOy
3oFC/74ljdQ+Uk0B5vAIv0yQuSVeWsxcA7q52tRo9+rh3ApauK3dUgIoR0IJgRYD
htqmWCk6guALy0juKXnYTdMOgVOVg6k1t/k0UsXzyXug5sHs2/PpQjKhDVjxqDK1
1DooNo9VtxStxAGHLjvEzJs9TIxY3QR5YozXYJwDduHexlv3RJbTTRjb23fM6Z2O
1uaW1LILbLHWHibrZ/V6BYTgsOM7+c32YkGA1twuY+jTTevp+ncj2BJqWCl4bjej
wmuBguvojRNNTzFyUa5nrM/TqhToKYx9FFxAKtDcq7HJhzhCGCAFH7ITmWI4ARIi
+Wv1kDtu8SG/wC7MZV+e6hUSmb7bY144f4HH9W0Ckbk0ND0snurSgn2HpF5R1AKy
ODVtqtcrra3PeLQ7SOA4lSNb4q3EdIs4fCsSbJl3tEa4/63GP5q+WX4wsmImfFDt
e1IdIF+X1MhCx0Tdjw8dtzagNihP+zwmrDcuNSpfWjP+RI6sC2ruOX50ha3f8+Ks
`protect END_PROTECTED
