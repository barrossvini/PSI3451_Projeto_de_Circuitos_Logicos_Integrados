`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iIO7cSZj7y3EFxHGk7RcHPGwOzLfMiGj3nf321WcunCmU3qcXEaxxtB7KOqZ65zY
oscmGlbuL3TNyKwmioxbLPN6h8VZZW8rfZZcBhITkWB5ZieD+LL4aPhSmlCBPNVi
F+kWw4JTdgdxIRNHo7UFYlx9SjbwtNMMJ8VHILK5iTiCI7Crcw/tuIViB2SjM27s
3EtgQkY0YwJlAwctFUl6k+NUX+qY3ay5LuRjWu9ouI65nXxB4vB9VRGriCLDi6qj
NsJj65tObv1J/h53YtD2M1MqglXBRYAddMlQ0J3clPKvO0OpK4p6pCIkxY6+ND8c
wgtC4Xs16h2xwZYhbklOp4289Xe8sQO3sVfU8n4oaRGWaHYdS4ccTCerbG8v0RiZ
RoDY9LFijG3Qkic2hedGa7hSmaSocVTLeAe/GGm0c7BbMwO2WxDTPxETySz19MZG
tAH27cEt5lea4QJUgQyz0wdW+z3iLLR9oUZZMG1xz2lnFmiqlmKvl0MVrdw6J0Et
9mODRwMV8Ex0BKzKgPrzleToUA+iRLW+ij6T2XKSEbEtdkGU8B/MgBvbR2tejeNd
8OpF0X1Gsi22UYa9O22E/V4eUueAdAEvwfU/RCH/iT8xjr2mKH7zcGAsw0jPmDae
7TYfzb8FCSgPCsTGY/Bq7M8cfGy3SKSyekf0t8TR40HkS5tcYEgfmEDT2UDNjfhz
zff8YT+7rTQN3jAShnEKfYhdOZaJjOVgr30XYyt4KP3pExvYHoOQJ6+YTBlrkKmC
8+S18i9cHs5M5Xa0XojBsMDZemzPVMQySRguPI1/A3u81+wzRpQLxw2rZ4xIIMMT
o/IhloC/jeuwk+h5fN/2VqyKcCw7fypdrNxWK7GVRilP/t/L/SGD5AZDb2LwvLbw
6DKYsC5JUQHXvYWUlDS70T//TRLrplwr0i4L6yv+cQazwe8L89W+J33SqUH1ItrA
f7zAPHVAcDY9cMJzCAshU83yjxahSChw1XmBZttsONA9LLz6VK5R3MT524mn02XZ
bUjW0s7F64OIHahZH+hxLbZoAhaCYMY1+/iBioIPceR29CPI8XNB5sA/Ki106LX5
okwIGHHP1mz6X5Ewj6MABb16eA7rWmMW9Hf6hjp6+CZfelHKSd4zRw2PxvSNRwYv
U10m2z+i6lg5iZbKBXEoChvhElK9I1p9h/ACje33gTAwAAqyJKb3QYop9+ZQRVqX
CoLQwu1R0B6hbZlkjFLlPIn9/DJsfY/Hux7SKcyqZ+k=
`protect END_PROTECTED
