`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9WPbc0IIdPXhFKKzVZgBwfV8qC1E+wBinHTH5dGdKR5m4+F3aCAbwiaeLhphTY2
DjuH/vXtfWf6ggw8lCPQ6Lyiz6WWLQ4Le0k5YmUAB3aWG3SUDxiiAohQkGO8dO89
buNS7nWEKwI8Q5Z4s3yAw/C7jXTASD6Rt3t0npke6X94kajGZWODwNoyxkyQ+cRB
nvYWimt4vvzmlWhGt8sMjRwjFK7DrPL4C4H2jgjQgg13vKqBRLhWo9EK3btepHNk
DLf0w2c3s/0S7qDLRK8vILv0986NGMKLl2E3qjZgRrUdAs3MxISsHAWn2RGQ944Y
cyszWUTtJYwAKm0Ls3+73SXpnmY4M/bucEJIC/oP5MZjsJzUE+lk1Ys1lAo/RUE7
b/KGELxU5n83iGjXVwXdlDCiHJZ0gRm8ux1QzKVhEyPdYSiFLe/LpWltwa90EDdp
j5Uy8IJs3rdN7kPQ0b5GTXkyNRb5WfAB4WL3aL4/VE8jGmVtBDrr5QnbjYNRQzNV
QjtuJQQPQy5663DYNML3EDhmf/A4jS51+13FoNowhP2hb/p4I20/yunOzVKpmfiC
QefoCtToDGBHSmZHVtvu0u5uVL8XSjVvQ1YX7LwE5YnJxWbz3bZkKbPuXgHE++sM
Qd+RuhSIvJb8fDgKiRtShClr3OZXHSTYdL1YSUmqwaiVEH8WdqoSxsNtM10Pw66w
ADnVV9eG97rKoloNdCvNFJGj5zUSwOdO4ZCZKa/3D0ixwaogUpv1Q0HPPyiFeDaE
tnNWYJYwTeVMaK/4mMtBHhbW+D2T1sfNXO01Sm/LsfnrsKnR3yjVux8+AyeoYc3i
Fb4CKZMNsTzOJRvRiw+H6A+IXAlmrwVOM73OMqWbJWVOPVXD0+4Dx/MckWi7s65+
rGctwaEUpYzjcdyzd92Kql1cvRuuKOL2XKf3X0MrwlUtLNJk6IuOg/W9BoR7L7sl
xDv1Isq+Z0xu/b1MZVK8HmbtEudy7aZC9WGgHwXfpsBwgfHjgtwIvJSyEEYzrCMH
Uoor4yJiYE3d/wUOuB3PI0h1oHrOmoDxIR5mszRf3k1JPjl0zBu6DcSAeeiehWY/
ho4rNs8vmryFcR+jBnfROFTUIUipSfv8jz1bFULNsjNL9n9o/4ZwUBBfz/oArWfh
J0X0y/NPlXDDlKLXinJQaDOnvdAZ6xzu9y08+NLDPUlDNgiKLJSwZgOdQNpm7pBZ
p03eIRjLsY/PdWgjAATa9V5lbI8OaWZveVR0u3r/dKstsgm+QDw4EOVhcOgwUCI+
`protect END_PROTECTED
