`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AN3FCHmVToHe4UxsYG/ImW2TciRkT4XJbHUkqaw7mq7Jk7wR+SZg4EZY8eZtclsJ
Rcb8FOF0nlnFiyU65OFabok1E9koq3g9ZzfR0Kf/vVriYBzlloNmwDnAn+IZmVnt
Rztcv0VmTiGOXqPrvdIAdYFIQfayufmusFxntKhO9aurq79xO2S+nXwMP36yr4FL
H7uLPUlGfecjliu+MMhfSj8sX2o0Emuxhsoam9/8bv49Vd1TNBydKBYOhbeWIhjF
j1+nyA7HHaQbZtb57yye3nXpTDowcg9mmj4q8t4gNFHXxrVCobx9LjS9AAMHEgL5
2xm0es/QIMzj/1lzq38VNWovgSBnihbWZXhwVpCmzcz6TMD3PlsbiMhuU+8KOYR7
O49zsRDD9NaY1Gwg27pfNbuwhw76w7bn5m9SdBOq8axMzHeo8rI9IokhLqMZxsJ+
yoPA56qsdqLR6oOWBkMA4AbKWbSVR2pLM43H3NSMYnO1VfBc0bAHNCtvUudaLNUs
wWZCD7BJGIkhR7Nixs+oz6n35It4pCoCIGZI6HmuDaUPrGfM+Xj1uj1OKOep4YPE
MKwG3CLDbGwKvItyJ2ch7txP/fdHh/2Ve0OHR3SauTdQ9B7n1j1hjz9zuS+Ogout
jidiFRoY4X4gKo/kXCj0+567y6coiP2ud1vWDIn27H8=
`protect END_PROTECTED
