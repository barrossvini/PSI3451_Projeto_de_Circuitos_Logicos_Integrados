`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
57mdH7itggvp/P8smHw4lYTjpGMk4ccMiXbDO3Nui6s3ARuju5URla6krQymEFia
Jeyrsq3N7piheDVQdr6X29Ed4wFeGjSQHvDq3Ze4fW4l+Cug+QaSg8AUo4i9gIGd
J/yRjQGs8PKkyCdGZFMVzQChz2moMoEZv63wkZXaBFSfJOeHngLfUpncws7+KGgY
0nINBfWmSpwAPXeyp9da43rFLCThcrZ77sMew8rmy0W+aTdWHNwxAj47IKyj+eTv
0GLnlXzzAf3oXTZDuNSbchWSmRUd+g7PcQ1eCP9311Xh2+9fvWsUQTnJuCph4rlg
uKDcgz7oSe8uUiRwfcuKB9VlBRRgudzAs/rDEkR+Bpaer27R3enI2EbXVQ+uhq0i
oKuRG3ZhWrJJN0zz5rrpK8ogH3TfiDLg1GYN+3rKdRd+YFuzR7WHEytC7JscFugX
Vf9jZrIZDsH7lN1z/9XZj7NElWao1GyC1CjL8gc73enQT7kkS4EpT83Pk/EGyR4c
5nKzkvr8XgTGjwY5Sf1P8HuWsMVGc1PuljV2xHKEiJVJcrnFrLaPgGI1hpiznegJ
ZVU3EoY+6iTpmzzR5zH6UwV8xgNWCH03nq1POMKq7lYIT6A/xlCFWqStzu2j6JyD
hWbh71H+t/eXwGpYjJRN2JNtOLdyl9D0SpMqvSrkQ/Vz64QXkdhJzhco4gkcw9fs
pK4Kngc5CK/cPyJtipQ5+zl6vo6fD3kj7/n0mE7i7zdDk/s5uO3uaWNX0eRUEgKa
OLLiQYH3KFdSYfLj76j81+sYarJ2uHxoymlnf6JuKsp/sTV5s+LVM+qg3ndvYNi7
J+Kbtp5jsJfHqPurs67SOKCOudDtBVruiOBgT1jJVJf7JpEtH30qmsk2QipTAzK9
BkgpwdlH9aXgwIa0utlWZ0jxIn0bMd4GrHJ2O9tGGlsPGP5s3Bs7jZC7Mkb4yAtV
gOJNNz+GwuoD0OzSKPyKgkhyXeS8abD7ZL3wYiwVZCA9NYY3xTSP1FLZowCZnd/v
XxK+mkMjgcTAuJuBnwATPra/yUAnZxEkbyvd555avYPoOoZPffC/3ZHkr1UV+sFl
qy2QnvnJos7sDgnSPijOaYl1e63peL9b3KsfqIULwAWNinloNi3EuDXlf4c3nbsx
cDf/xfJU2UaTsBWgLSFRW5UJ7nWXBiv+TkqJXAMt8Eg7PgVNlB2g/sWE5uKtubiV
bXgRIvMlABoOwRUfnsaWy2nF2MOjG35QfHu3O+rscn1i02OI78U3QOLLp/QobJul
JbrXkcSIBlnQFP++cXEm8cOmtmn2IUgEYP6vrxwNjP/ypjorVEuiWmk10Mb5zbCp
htjYIxuRq5O8EGo2uMgCwxBPClDIx523+3pB63AVNRJNHqY6OPbKPovMUmgWINuw
pvFU4s4CjwiTZ7bi/5apu1mqx7B4nn5vvIrCvnQJ2Yhyw9U+MD3155wdJg13xOeH
`protect END_PROTECTED
