`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1qR7JvWRgRua3/Uh8ORoG7mIeSq9CQdJQQWR5tMnZv7dxZ7sLDLNfIZricCK+G8f
aKqhtKfBTiQOiJHzFBHoxy9xRjestXV8PfmwP52oo9PDml3r8cv2C8HbiFHSxttr
qHLbmu/74VEOPOi+J8qSn/Ep+3p5di45TUEBZ5uYfIhQP9rKY7CipBcKhqLzelkN
A40yOdTr3SRQdQLphYgI9xlKM8bTlsMf8OVzuHDncfVspWSHBGZZ9hi1zlIs2owT
ReQmREowSlUxAvzsGe+CfknzqvsyM5/Gf4J27YAcV72KqvSzvtXqYSdXYLIT4SA0
775zuKGQ0W1+fwECwyv4RoImjm6ZzfsNa0JAYLyu44R/Xy9b1CFY55jdqwKwmNL8
XWX2ttWeqcEiv5ioGiq6ETh5KmJ8GsweSpTQ5ao3bsnxwHtUCUW+aLXmlQmHDcdW
pMnmclNjDdSO5mVbsuWDTUqlqk5UIlpB18WiZrfRe3PNlRKXaymYAfKPBuJ3luqP
/nZoO5BwU/biuzFaMsIdT4/as1KdbL65rZEuB7V8nvx3ugho1SBvMClgMxGrSxfX
F7EUDfrAppz4RS25N5ApYpIcjbTBlcjh1FWr3OpveCN1pGYzIP8CFGdUMhBtyvE0
3vkwB61DYOCZfWxdFT9w+1M/oM65y5f4ZAVT/jqr4MsaiUTLcjpsMInL/OnS1FQZ
PtyvkW6wBWc2sDp4CCD07TrZnH8ZztdO648u3TCJ3+1Q1pXkUQhVoi7QR41X2dWq
YWW8ja+wo7sGvVxrR0BEUifZHRV95NjYmgf86k49FlXq6LzSXN5lEPmoDkZhqHSx
HP9lGs+2CXq7ylgpR65tyGvkj8nuw+MDP8s2hUXNO9l2+ynX1SLy+wNSbHWhv812
sdyWmKO8tR+KD72lCdvwColbrb9UCk6A1BBfKfWWWz8=
`protect END_PROTECTED
