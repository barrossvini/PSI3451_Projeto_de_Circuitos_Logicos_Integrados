`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ATR4qBTdC2bvst2r392OYZL19QXR8EfIYjkD1Vdq4uT9zY/XVllmskTCxEHdvP93
NbzOPwaAQjUEHaWhE3GNZu+3TbnflffiAKNuAdgc0QYwJmh7MAqgOmCzJdlPWjPe
MViiQe/e7dSry26b8bbepw5S09A5zLoc4gBpedJr1K4jYgbu5Cpmv13E2qqIWTA1
mKn6jNnqQz0JfQOX4lcmmBdS6H969KlwoBK/4qnmZlN4SYnwrQDRy33WPEWl44ME
TNRVs9eNQgPcZT9oIcLNtqvTmuUE4gHjc85sML+zi+ow+2k13IlsNW9oy4h0pIYW
DjMrDH8tTAUlURQr4h8vZalFJuE2xf57yXU9luOlgpkzsJgDWJlivimLG+nLLbYl
en0it2fIdMBvIcCG3UwvzL4a0zbQFmxRC6/K6DhiIOVpvjZQklsCGzN00A/HcZN0
dsvIr+rQ6LbGM4n2nAVYRbRLvS9qKF4G6Afs2g5GV2ZGeINN45Euf5PJXkvQj/nz
p8IMJVS9KQkG0FivScet08bRSTRkaZHc/zpqwQrdZQJd8XI1+CJ0YH0CxH/ZK2P2
5WHDlDLd1Aa4ba/5jtzoKClhVWAStcJYQkItkC5/9seoMiSe+eYyppPjbQGD1IPU
AHdR7YjhiVp+Ktjb4pMVSS9nHrPi/5t4BkHoUPabgSt0p5x0D9Kpf23d4BVOrm7e
CBvqgRXBmTUSssW3FlLBH2YZMOYpjKd3ohJzqqpgRyE5xUwT1iON9quOf81qaKH5
b81eyYB6Ue2/sSsdXhno8ct9vyYOTmj+7dfJEL+J/3OZHiFVlXust+M/MBolF/Ua
Iemxmq+YmPH4L7Ny7hVOCmV2LzgmuWcLZikua7VSDv5cQBV8AOORxdBO5hEDuo/u
0IXAjnwbvZ0qfk8YBpaq40cegjZWjbNsQRevfDfrhUmG3GeZsPcxyogqMlwpc6sn
J0Tt442AKum3YnCFFWSe5kchbtswcOitXSb/IUqNOccLAXqyCoDrwQz13LuQnqxm
`protect END_PROTECTED
