`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UPafSlxrC6xeILqyBJ4KjGwUfXgVOIFkSROdEjOTP8YGQQE235mUYP7rhswdWH/7
gNRVzPU7AWCn4rKllPS3yNAQ3BNJOfV+bnSVQf5K1sm57FXTacoIzCu5BsF5VcsJ
cx7pONoCXrQftwo8l5dFjrpsQo74VfEBtuAdVfOkI0aAfxbOYnK0McCu4/2877xB
xUUFvOejX1iksm7Er+Aqo/EcDSQ9NjcvBXX9ySTzKp2DGu8sA7E0IZkfe2uozLhq
Hl4VAw3ilcvUbWbCdFBvB6cyi2Es65vSX4duC3X/C/fAaPTr6z5gVEBFXNOgCnnw
SkPxmSN7GdNuxYD9vslDkc8g4V6KFdpkwKrkmKJ74wUTi2HUsJID0tNyyVdn1E1x
zqIaEy50usb7IdVxkrm+UguKr6LNHEmwTDE03XrHu8zMlQeY6okvqljzGoX8VigO
c3UEMLiaSUJ4C8ube+k9gnvdvZK8JWAncCjwUExh0bJjNxZ3LPHRAVW0DlqNlNAH
eeS+VEIoBG2l31KM1dGe3BhqagHs9BdehdM48LvG/rww0+xQxkvry/nwRl5M+Iku
zN9O3GX/dfD66Z6bRHK4mWzPdW0Z+8+B2TKcYPTZow65QbcyOSfDo7f8dM9nMTlD
4XRXXoU0iQvonjMtpiMmNj8ClDQStDL+LUa9JVVC9K7n1w/dGjGiASnYZoN7xsZM
`protect END_PROTECTED
