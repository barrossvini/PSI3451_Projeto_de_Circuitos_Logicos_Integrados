`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NICwx/OdPKU/2qcqCrzLozb0mKAFwU5dqfPyJkzK3mh2rasvnuMLcjcTougKpHE2
u3a6TKA5wSk0rr9PPQC//ZqXV7RBGEkipJASg9QtN7aZFpANTrNfMmLLPb1DSIQ5
WZhookpytrygIeh8KnP0S62rMsZVd/CHnRWQCVc4QP28k8UJyjLhxvJTvMTZ07wz
QsYKjSBVQwrtYZXFI4j0PppMwrPsukQPEig4crgE0Ym6VVBY+FGwEFuc5Z6Asj3Z
kNEePmCXOlvo98UqDZowh3WhCgPS1S+aHf7VbKYfkLmcn12/7wVJ84O4IaksrBM7
yqPLZxMDXRcykChXcwevBhc/HXgJSeH+45kYKFeahBHIUAXOOUGovG92G1puloef
Em/Q9LlTe3mYG4elh//SY1toIvIWHdKNkNJgJBNhY3aDvkmfUJya3Pa273+mgT4r
bTMkR8+laXL1P3lgfI1SKDulRRWi7edS702TID5kwuulSuvDWuofvKWR+/ELWpFB
FYP6Fjg/sSPVPW31hApCH3UQwoCvSSxCRXKUpezZTZA=
`protect END_PROTECTED
