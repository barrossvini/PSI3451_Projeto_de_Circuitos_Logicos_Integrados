`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mklrXhUfqnKA0NnhvyDDig1I31XCqIagDviWJrbgraBsF+MgtfADDMSsfk9lVJmH
rpS//BDtGcRQCzw7WRKCAHI0Aam1zuvRx787xN5LfQiOLe4bdv4As7+wKKrx3Il+
2NauQGR022davZ5Zg4z7UglnnRejuaRiyGnzaF83sfdoag0cjzuqjcfSUul9XCGt
fdVcVQbkXztDt9dfazPh9AEZ0fw4nsyJ5q+TCfrlPBqyQNmmX15Rm+Nqya0vNb3V
ft+YrybyzZ0x3LDDOC797495IPlZ8lmxNtJlUqtdrOxzV5uozrG/tRHwniLWYmke
n5vm/r5PTHZR+lj0yitWs5o+yu/kGbMb4421RWzvW7FEAGjBK2cvolW8OYN95d5Q
bc83P1/Cce5Qc7YIhpUSRpdzkS/YrbfGh0rp/tuixvTeDBptA5z7Id4kvVJpdBcE
FqBmtfO8H2DXxSd8IwTOa3mU4BzoCevPBbjvDnmTsu1UEzKb4Im65kgW3J5a687+
9+xj+0zTHO9UjoYkB8o//s0J2C647enlzuvsIGRkc4U=
`protect END_PROTECTED
