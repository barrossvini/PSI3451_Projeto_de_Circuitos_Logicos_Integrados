`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSx/0SSea7CWN0mjXUDv4UVxnLbEiUcSZyxhry4ZjULUC0SQ1EqOGhnHIJ0Df00Y
SDjvaqt6EG0nKexSsuUC74W8Jm0liDTDmtTpP+3voK3Ys1Dv5hUpYI0FTDmVVxQt
Xd71e6TvjEIBYVPBXsS1JQpX6a1T4LORgZNP1YrP1fpd1ReM3HRnhuiixsbFSOMa
ztnoUxGMaUiqDGpBj6Wj/rMdpWjrCVW1rds07L3hXQEbA/8bCOcyPtJKFc9l542N
WPsUpVB4fBYK/yI2OfGtfxIutFYkb3k0fOrBZVj6/eK/uSSndyL3l7AJWVPr1YeY
YpgFtr8YBDN36dOWyx9RjKyNL/FoKTtvtvGaAnbsqNCsKPDB/U8UeQWTosmghwLE
RDZtcjTAbglNDqk2zhrVO3EkfL8jRcHRRADr+1Xuj2nTFCmy+DA/0qaU3vTBxtuU
CQA8UJo47niReOd4Q4NXnk9zSXmQdzZ3JjohXB4P4CTJE9Ml40/D3LZtN2SIkziI
kDQMmrXy0JGyldgeIgqTqU4GpFgPVkxbio7MPiU7L7zsiPFUkAnZTEiO9EnfXStS
N0P1/Z3kEozsoNgYaJeQ1LbC5LGK3P6hPdr1lvPxtoUf6Xc8ENhZUM6K2wYfwN/M
nhL2dghWSxO7OaEgwEtwxP7fWCRtG8Njf7fn/4V7ko3fa0VcGMISw6IVZDjmYuN5
zDZRfqFHLL+ZyfO8TmPS4J6XRLu2Vyp5HtCaMCG+/Tk2UeXXzHEzAXQQY/hL6jCb
k9WEzxrEQ+xTygliZgLaseeE1q+EEguLFg6wayCI5pDYyhbflcN3IhHVvUlm8j47
dr/JPhahyRSK90QuBNHcXyCYKJp0SwqOeEBzptYAse/i+EtZcqTwPvMxrxHUGtKX
pW/clkP7i5xPdCCNdvkgjAzy9iINIG2geEoN4ZkMKDeJgFV9xHBh5wdJt1wt5DNh
znxujzD9Q1eAz9mxJAteVzzQnndp44G1csTZriprlbcs+LYUMvzHEAlAxSvQZwFw
2hElv4lsEC4NVz2GC6RfQVBpIfiHUBCLm2fRnzcsMmetBPPtUv79sl6i+UhGUonS
20ondEfOWXwFsB50yQSgPITySbSTyE26YUlOSFahJydMNmrs8DLIMGncrgshEAyo
o2Dt/hgXPRuJEI627S9oSFTAfrCtQarVCWtv2bYgO4BJ7qavffHsOmU8jkLXMd2g
bvVJLXGmXDL7X/9eOLEXyRgAUj85lNDLqsVdM1SXSB7cq3JMfdMrHbVvFQyUUfwA
u4kJ0OSjRZOZgAW/vKsJnfLtAFyv6HCjRSDBGtZhcFcD3NKAyAAhr3A0p1mT8tpf
5RVSERH1ej7pNHdAybHpFkZHp3CKZFWsF/UFz6KDjVVJrZx7vsmtzVVTWH0SQPNg
Dvd6AcmbAkNkVj8n6t7IKazKaDmqU9fVtrnH49Mwhy4zB9/nC2IRRolpG+Cv1L2O
t9HjxYbeYFwDzQVu9BaxJ3vlNB5d2EP7RmqU+hXiOr5YsO99MmQfZdtu1BJXad0e
kVeatq1falmaJLtRdkKCjNg1MmN5PZZBA4LU6DjA8mRRCgdSac3ANWYBedHeTAk5
7/euBiUSk8LBKT/IrOlo4rMhe6HRh4pLCSiG8rITFEQdBoD4aPWoSZldA4lAtbUB
tCrjKY7AlGEeHpurD+tTA7KdB5SEBXJG98ogiOaOJISdE5UtjkvycVNKL0jCvkrg
bZpFw7GwyXiK8BKsQqbWOznUJ2nKdHJA8i6iNkV3eHDwaKzeHgP4rnQ4ebepfg6y
FhtOVvCsOiCjo6y0vtB4huMuwbiEot7lUaY1s259HiNicuZAn9nZKt67vmpGHA/e
+YYgb+6LP7NE0GaxctN9DHIVZYy1Knc9PZ4xhv6OaBZKFVgdBsBCngHii1izcJgZ
14YP/TYyKS5YLFbTMv/fM1kVjwwliqMCYKsUIIJDY+PTG7pwHtO+onAksH2Argr8
9/Zn3RKR00FMUY7GD8SzOQDmeVKf4nB+xWLpG6E+U8Mj/RcD7P0QIfNt9ilap0R7
t0pugfQsvPpVarNDznmhvc3cUxmAsc5X94CQUY3G20rCY6ru9cdf70XHU7AnBPs3
MAWWT/jpcKdmQ1TpoO3yut0zbL7KDp60kQdsQ9GmZqrrXMlWfIUnJF82wXYorQhu
aADTtyY6A0SfgDsXqMmtB1XbFo5pFdNvaqSpY3N4NRLYrB9YHG7JpQ0uXV7mFB8V
/mC9/+bL2XQLqTJ0kq6ewahsOwIjtlOrT0b06nTTNzo1HHjFemv11HRLtExpW9Yp
+aNFBgCxIwhioHy1JlcbYuX2AHoa6kTk5fR+bVKh5qqbkjqOtfflxvzUmpLMZHkJ
eUDbewysyEmVVbMPY7GhI0WrNY2A6Syh0JscxiduK3thJUvQKNmciW+kr6zDnYgY
4oYBgOaLvza//+R4pt6aKBdUXT+7YTCjsHEzEuMWEF+nyQfXHbW7Xi2xODtEDZUY
ghK+4C5UH8zEVvR54DzGd02KNCEB4pIFBsO+/PE3t3kvTSn/ff1qePPICKdxIiNW
qLfPoeiXcxmpN4pXlljeydncrAS14ni5xscCFE5ufI+piiI3nb9V3uEYeCxL3hd/
eZJcqqNSqNzvRwulDGUpVdkda485V4ym3VCsME0suY/Pfzn1UiBFeA0PlhZHvGJ3
/fBoq1ASshXw6tuO2l0fDfkZSpGFzy23ssn/mHMG7P1AIQh9qYesNh/wkefAKDmP
822QzPDmtCSy25ahNOS8gYwRI3qQoPD4l1SMO0ZgVQL14zgyIPZm7oH4wJcv0DgA
bqiQ6GQT0uOqBEizqyW8fw5HJQm16lVjUrTUZY+maPReauYnC6NluZj6xcOHDya7
rKCbcuAgA4lkJPUtTLesaoDx+1Loh6jbzMYrt0k/x2RzbcOZgev4/UjnGyfQxEkS
cT6+LwpucnhnObJEYk/F47WdDtMwpXiisAxqpwxKfmm2CphmT6WDxoB/fCEBxHbF
aP+F1CXzNQ/5A76FsD+VeNpgD3DM8V13hKnBZCS3am31xR8kPNk+5N4Rl/RdwO2b
/ckRQqFvSQ/CZ+4ASIv0vWkxyRcQ6nS5W32YflY5Fj5aAVD1nfuLUaP+o6YJ8z6M
QbXw3adYH55JWYOHx7f+yRlbphQSOARHhup0OUX8faKY7qif8hTQnVU+WoEW7qb5
lDQSbtAQSJ9T8GImckz6pNAPb8O0t+WmHsDd2QeqYTnAZrWMKyanl5svw1iaNghO
/TnCNMXFkfwKvljKaSUDYag9lTqvwFnEbKTPgwA3uJ/26a5OQ+621iuYGHzVW29D
Pjh9SrzbGxU+oIFwAfEj6rIntfxmoLfUTPwH8zMDF8wv9mc47b6o9Jc1cfehNXvR
6ki2QVtP112TDUaK37iYzmDdjIvz/MkmGHc/7da9d4tKhGSfyaZ+5nAEw3/wJA/c
dYfLgqW3MByNbQurNP4ze6M5YbKlr156VfXSs5gbQVxH5hJuT9ICEUAsONcU4RdW
s+8X8FqomZRFeySrt2wjD4iHrxX0yTbZ8xSPazJMSTr+waqgnu8MnVyWZhlpIzIG
ANJkaYcifdOufR9Z8rmXeFPrU7T4T2TdWAZQUrAH56VT3G4EVUm2Mw2BmLQSbwVA
vn/Oz/drzgdX/LpqKLvGfquF3qhoSolVxj7r6CGVYQL0kdjSnqzo+6mvSRHp8bYL
DcE75w7Vy+TKoanNMkYb95UgltD0khXVDhpuCix1akxSPaemBiMu3w6e4bhCL8IC
Hol7qaEMC4SixOMEdEwkXSgic27c0PQUmCc45nAcgzbTW0CHpKlN5U9/Q0JXso10
tMTdFCMPCDs9jbmfhDD1hX6FZxl7gMJxeGAF8uND9UHOBI1Dk+miZTvegD59pUI5
93N04P2crxyfaGFe+01SW2C4tbAxEf475lqGA4jPocBNlH0rukYkQfLFKeEvop3b
htkjfh7AMRrX5s8zw8pVecoYHDX98gwKfo6mvxeTpBzsOj9ANgsf4mUMcFndIYkZ
FytMEMUTsv2pVTG6FgPyGI5Txc8BT5mLgFiOoxVzlO7nCQvHk2hsLrtewv3YoJTv
AnMcL4gonwZdho9zgcvkky4gNMeINtkJ/mEuWYcSktOHE2ZLVm+/li54w+YdERgd
VqyCJNBRPQ/1I0z+Veo9mrhCCWFZMRlG3ZMAoJrMZLUz5kEkEHHUD70ZzKX/k+Sw
I5/JhA4sW0XaJDKkmh+w6XM0LJnzjh8nbhh+UMavxdosovl8z72hXzd0Z15v2C3k
6Y0dmo0yonYjQXfhODbLqrh/x3b5SQJgRhf/dvo+shfhWsAJ1Vn9HNd+v25sQTrg
Jq2Ee0MfRzd/KabgjJdQApDFNEmhaJ3OnitqbzxQNzXVblLie3efgl9Q41EeF9RP
JIw6FeKshDumoPHRXUG0Fg1nxMFy9lX+u4TsEnenIN7zczjon4EGm6+yF28KV0fo
Oc9UobzbMVeAaBzc6LVvrdtxhF1I6V+lSgHiToW+1inNPS/L5q29UjjARfmx6r2S
fb7BV4UKdIWJ3AZRVe5K3HUxIoeoethqliJuj3TCKnoevsjUN9VRtuEalU4cuo1E
rD94bJDDB838unrgPEINOndiG1sdhqmnzQxV1XAidUwc9//1aAnVjqdBUqyqsNFR
DnlmQ6O6S2dnZB9Xejll6D/6G2arjGS/AH4n0x1N8AsJWNQ+0X70Alg6Fd5jhG4Q
0nbEapDGlz2eYfBTDiB7TNo8BemmGFbMbaXMY+KzIO+VUnG7Np7YYXkh/qiVOGXp
iVZPru0pyFf5ZuUK4b/78bnvIx0sjDThgxVGzWA3AO1Bf0bEbxZt3FvLnWrnPSOt
UknWcyNFbcjCwDS6auw7wmGfuoNUHuVws9x6c/GlGSetA++rFx2O98B+iChs7ZiJ
46yJXRdgkpnhZfoUA8rAm0fuV3QyXipSP5Q9BW3GpGMbzn2YSHBCCs50WVmFwia5
be8SgcF/ExQhPJd1iuvfE0iyOwdqxKeBtInysPED84S19oLrB8+wlugMc/gWQ4La
CJJePknaCSdExOmTbD8OCObInCLBgTasI8UQ75++UFUdCLfgRry99ENBSMS75i8B
DAm5JcK8YcyhMWUdlGM6PruNqbseGPqyqntMFSFZbeVBvtAecVAtf4/pyVIO4gUC
GJhrNb8bm1VZqT5MUuvn62Fwa6bY9SSFsUvRQmTKfNJvwXbwpwWRDLPHR+bwq0a+
sBAaMO57Dtn+0yAhAc8Eq8p2PtZnV8gnWcuJZ/zwUr+EZ51TwMBSNZZlSGbL1wsF
2MljHNEZwxDRTH7eR1O/kPWvBei+DosDyyozeJmgmPIj37y3B2IICbaIcessG7jJ
zv3yBGM5ojeiKPkMRSiBgkwimHoyKN/YaWZ1rEKPHaE3Z1v6xQGG1Yhn7TumPMam
v4wYtfQoa6087KkyR7Jm3gHZ8RpGkWAIyXGx1BjD9eN7MuK/MMtJMuLyHw+AlsjB
mE0Ewe9xt2D4xHIDZxFAgWMOoCQQ/2wox/CmsPEVNz8lMIkB08vK1prCPOhnTeyd
raP17A/bkHGrNL4Lm9iFasU5+tkhFbFCOVzka6+/HIerP9kQowloAoJYWEU/v8nK
I9XX9lNGkdDx3XvObIXrLFlgK8veYCAJTyt5vQw4pUsXQvCcV6lbglrNWiQXJifC
PIkdwA1kp42h25ROdpH9vRN4xX6ULa0oyBTtuG0V+yDB3AYCv1n3EFZiA54/J7NO
kV/J456AkTxX4PfDvTCFechfMvTV4eI3zp3R63ndVv0L4wHsnK+RGvhCyQ2L8s17
CZmSKM+oxcX6rObhEsrPttgbyEfaVfdZ6rQCMqRS2qL55yQGxRn8zp1Pax4EDWT/
q0+ejRAnVGAM2TtK2PjbIIcj6QQRTd6hEt+DzHmYA/JcxrByTsPyhM9txuVJL1rZ
sg5UFQdsHyuPXjwr1mC0mvrzrEhCIqF4aZWO+Oi02W61rXRb6SiU5NEf2a5WZ23P
Sc0dC4KIPNhby/W8t5vvjuCwEw0jcqAgcDa69brIvtG5f3JQ2BaBHe24Xm7pJa6E
IgDJ6JkF9bYUDTJOp4q++1Ae8o8VyrGU/My8AGGk9i4/FBi4XZNTKm8gundtphSt
Q4o0qB2xbRASftBD/THEdLAJ4yql8s3TFtV+PhhBuiVm3nJ5ejI9ec+prXK51RTH
NOn/qb6tqI4ETaSNHcGHKgkFHg50HCWSbqKT0b/WbjAj3Oimx0S6UzmUOkIyZx6e
/bvFUmsX1yVm15gqQfKBc+l5ArC8m/j+J8YGB3s2eCJisAkX6Xf6ly99ehEX0CXZ
KLT7fXDI/EHvaNY3Xy3WFJo+RZHvWwePBLQbcX/mmzVKZZI1pijw1yHTVau66K+S
QHjS+GNpFng4UhEBcJUVUDsrnlPWyRNg8/iMH138nxNbZ2rsboEU5qk/AYPb2rM7
Ujl4YR8mmbuYm427tgsiFXpz3iciKq9khVI65yHOSSB6C0JLDGoI5l+yqXc0DjLE
rjvRIC5TjiWd5tppuc/AkSrciI/qKgw3img0WmLASyFsUikKHOaSfQVbKJxEhdNy
ninUmlvjW13qZbD9dTbHRPnX3zhFzNyp559CPGFKAK1c/oPi7JCfUo6clNX0+Ykq
ZDEpTfEmeq5U+wWCDEETmAGso9davFHVzir3VxvkJubpt6TtDh+Zt0rAFO937q5x
/2Dkx5Z9PfIdXQp5AHF/D8VQTFnzWJdlA9BtWnXywzjIUM+543ctW9T7f0euamyw
nCF1jOOa1TAIlShk4WL8TCqK4Lqt4fUGFM4u4fwWUeCHFH+5eSDl0ofrfAn+lUfA
RVtAH1GkB5qjm+K+BSmh3hwYMv13pYj07YBWWUNi79hYEiIwpOVyMQe3r7DpoHta
34yuDOiDWFWlsxl9ur1EwMlgWukNhs6KMg2NDuQf/bENeJOrZznpSIyS3awFNLWR
cga1fkCgqMHFpqcUSkVI5TNz7awF/pZUi44DKVv3of4gGL50GXSTuM+qnoZQLUry
Kh7UKlURbDLQxYQwk4VXSimqS56SIYAFdEWsVz4zDE9XTx8o+m1eeiav+PilOEB/
9gmCJXfDiLhDJGQNF4ibGoHda/DtXqbh8tIrov5CoySX8FJEctJzVdvu0MvUHCZr
U3/5wXWFg4abiq78tDmy8bPawpx+KdcKzz74lCTYuT/pRBWfCeZZpCXRea/Y6qaZ
gyCK/DlyRBREpATkgFP6Ur3DVTjbqometn56j6yVWiasjzEw2OUIfnqsTMnsI8gU
bn8z8PHuRvJ3/3PNPTGeM4IpkLwrz0bjZizVfWwGC3fPzXXetjSiHAKsuQNsPczQ
LMvFg5+0B3UWdmdyOcxdWjF7E7ToRRXMBjVWp6BQfSPYPYsa2Wo6AgaBjwcmWRpY
PATvJIK5WQh+dUO9GIXGrbBttIfx/L07EbZZqrxzx5FZvo7woTHEM20r0K5COBZw
rhKh4Sm5kl2SXAloSgY0g4ilw859CevNwci6Mg2nxoiQ9Rb1nj1mopE6JbT+oTYF
msAv/VuFHTq08xMXttsUUh8WvJZS8lq/ut/MiJFzEs3AcRiXiTF0BTqh4rQ9YCy7
jVeU6dQpTwlb3FWJyXNla0JpSeItuHAdUCKlKwtBZxwnDlPRWSoQ+97ReXPWK7qx
Cn+tQ53QWxikMQ6T9pCKfvJteXnFBsxGhQRMQ/X/BaBvj9JbezgiDB+5kBnK0ZTI
E2LY7VoZxwT5K9LJeNYzMAi/T+9uiKMb586xGI1aRTgC7ae6D9qf1F4eO1sKIp+S
qeMFFV/oHmbqbADMSL6wXNIJ82YLM9EmjF9tH96J79mAERE/6AP4BsG7jgyFhTEY
y0SrllbQh2D9OXaEl9NzqkSawQ4W+Mk+VcbLdjzArWTsFrItC7otrosNBhG6yE2H
RHno0GHJ+Q5ut7TuhMtXrZJlXLju/UN50aZte/+ka1KH85Q0kDAanKZs9VEFVBKb
1OfehHzVvvqBmPT4tHsgUBSr1uAb0SaOXvlNuoptHreWfd/Opl7QgOmwG3JOrMjk
D6Ps8P654jwCcCxXjZA/EhvIcJSlq33a4KkbUkIHmMEnLmk8GltTcIqv360ySvMM
Ye4RYXsGIv6zZZFnXVXKEqlONdvf5gbMM0a3xmPoYSC6GmCu67at6hVvxtFo8Nst
Azj3K5G6hquzlODmqfyPb0kWuRQqW/j0A8ssciJ3tLjQfOpWR9PWEoh5YSl8khhT
asOKykBVdnfBwYXtN4tkzNV7C1ebCkuYrID2FfhWjSiJSKBj2px8/PrFvq9MIdyu
Xv9+0t590C7S0gHdgkF0htlOFQpRo+ilHa051dbpZ75NmlGNPJX9PhdpVxrhnq1f
4C1F34GDfXHGVl9nguXjAiKHRkBdtj6Zm6KuS4UNtaKRTpP3dL34gh9mDxI6DUo3
7BAA6wFNvXMADyawBPIz+fby1tuR93BWFBZj2hzQiRHUfFmsI9bODtHDgf9EYzgU
R6sVkAXK/1hxlQSVOk8ioL7gq+enNk56LTd7rWznzrRfGCSZV8d2+vasaLGygQ5s
3XRyorzDikIbPF6JGYg7VCJQ/B54/sUhMWVvmvIXKcQNPVTUemuXymgwgHDfVeGe
5FTiUS8sKdBn3Hdo+8AufmHDXNcVdSLZkAsZQkgm186tdtY/qajYACWkhlvOw1iU
OObDIcfePi5YdaTlHRocHIuib1/ecNLEJKBIowl9hBGrY0p1XHwcegW0dLurpzXW
iQNdtbZ9JGxW/uTNVR5WzgZ7fUIEqAbMWozMVKJMRwL1EWbtx2rFIJCCPBUlwXRq
t2xVWnTK1lEva43FGbIYS3kGxqJf4XGP5Dm5L9hJZdT6lH+al3KMpvnAmj5+RP2c
w9dmgAGIo4vU23fD4REC+f10MthpJN70ebhUE2L6tE9TerZYTpiZmnIyb0VP7Rlu
TJwsfzgAbxZhUJwyIzSNdl+QAcitcG3JxmBwsWubywB1cbUS6iZ/ly6m7QnsaZYc
M2QmXCjz1JI+gzI0xMAcNxcVvWiw8ImoVUlu5oNKFyEce7sGcri3/NS5XKG6R3kp
LoiltE87MudGVKoypUtWpv1JqMt/x3ghgxWvLx7IBNHJSzkeiNV4hqeRLUh1/Dtc
xtPYjtZzztbh95X+WiJJVegrzH0gCL3B6ASCqULY+bZy+0yZLKDmkqO0Gxa7UHjQ
ocxmjIqEgMhKokAV/z675kX0yBUNNtz+m/Kdu9GtRzO+pGV0wSnLMG6QztyeSvQU
OaeOQyBeu3VpAKCxXb4BtBSNokdC4E+13FPNiW9r7vdMwE5Uzyi9aTEV1opJnChb
sdYdW4lJHOvmtXVNXmgMGmGHnS3WoZb/qNsZlIopG7Smnh2krXssrOHJmEmmKtAh
0UO/UMz0kEjn64Ncixu9mVIff5cY/39vXgAtADyx/AvnrY10g7cIJZrRM1fENenX
NltdD+ObFgIIT5nIRB9NM/LMJ2OXxSuNHgN6zS5LyaVq66ZkmfLdR3sTVztKc3u9
/EnHf2zp4yI9GNk6poh4reTkocG5V4A8SRZdWSrhqqO2ZTwbycvNEr2SJUF7qTSA
Kzf+UCAI69FqRZQx9mL7eLrTdNAap2Fq9fKeaaI1fqxiDtElfyb2d35SJmdE+Rq8
XavMnV13iR7GD0VD1F4zAMXUq6MPvaX+xThLnhG9PEUYbjH5qMwoXGDI278UvWSE
j72Lo6bhcN43MUHm7vYFhNZ7rQDX7ELnOfd5uAv6jwj9WkDBQTYE0cVeJTo+m7lu
grQGE0VrkkMSUpLYUPtNQ1+wvLR9QzRXES4oAA39tbPipTPaVgLQfXvEmdG6mmSI
jGvQxi3v0qKeuMCfVDa1V03CszQ+gEMQJaJVnAtKkkQEzaQSX7AcxBHID8pf3SBE
EzduO1Ej4h4ta2byDDDzcS9hznCNXQWTxozMZ4qGmFtaxV8UDONqefFU3uRyLUDy
kzWGgnVBUdciXDpTCg1HwAIf2BYb+nfnQbiZXMsoY9PCGpixabxl5PQSzE1FoSw4
qlnbcp1Am39UDL4rzZfNOS3Xko9xGQo8eJOdPSGNAzRFHG6/1stxJNJbTWoYBbFO
LhuNofDIkWaM+h7greZkYurt3t0Y+/O53C3Abyspzrr1rdN7v0OpMGjbiuxbm+ER
7CvqXiM2fiZJ07zDChsSbG1vo1vdMTTbMSPJJk6Wfom+dS5svPdFwHuEW34PKbYE
/lxRXQ9n+Uw5LNsRCQshWfefDa8rvwKS1aE0WdBLPizTTo8UC0JzpN2uOElzg89D
OEROdDfcKj8F2oNWM4q1XLmtxbIaIDN6ntDwjTZDF4Ng5ds5pcyz7CrjGMSF+MSc
KiC7+RZ+tsfkMRXxcKvYOWJkrYPF2a9Z7HF9IKPZht95Xokj0zEGw4HqotV/k/As
7g0RA+sUg1rQd6P0qhqT1XvxDtik961/bzoYk0qi2NHlUUP91HkXxrjN8EziaFQr
UDk/1hNVYBou9EO9mxHK1eWpy3UuE+wSRqvFD/4L1WbDJP0ZVdgetbVUPglM7oha
zw1uReKYopd7ISSm8TZUHzGxuEFXnL0dUy69u4IaiEZfpNs1YcP03A1AygwSdGlJ
aWQB2yVQvTbCYFlfeNLLhzriVz6kdNF0mqC/YFeQahhx+/w10pQA00gnLFetYva2
AuUHgRkXkl2uDL1d9+0IPZTCJAzFBxP8BH4E8kuDiqoHOPMzT2TGTx3WNX8jzH8C
rpDmotThpQ/RbNk38+Q5MgDkbxcwOd4YsT6SD0OnTedhWXOpbNfkjBr9HU+ThtN0
PklahZLtOOGn3o2WgzmTR+wEI49cQ2cFU+vQp6kIIeKai8axRGctddSKTjyiYdHj
1h0r1lLQXq4Nh+StDA6w8ubjLodXV8lkpMCG4epHPlVVV30Z6iD9r+ljW5McT4j4
bn2EaCaWRn8+aM7Nw+owIBcrUcRn6ubd8g1VK7jnqX6CSQbIEekAaYop+OQ7RMuH
30rJidc7tAgHKd26t+CrTG16SinQDavIW38zkR3maB0YCaR+tLHWPKin1Ni0oYek
6KFUvXSyMpOo76bOT5o2McHF/06XxaJ6JOdOGBKYQT1luTrxlJv64oy87eW9D4Ul
fr0AIsLV0U7bqdo8sKmMWv5MWEA1BT/POsMLgv82urZk2F9DVFSbRtEI8Hyeq1BX
R7b6K9mRpZxHnHeRBre9vqPEYh2fQs97OR4getUb9y7cRrMboczWQUEgSd1qmFGi
pXEepn/6Z3i5sX2KTnK6PWHwM9Usan25Rt/jUE1hcyg2b2AX7RyZBBRknx9r6cTG
hJeFupRD714vgl3O87wcIKsb1I9Wv93hv9ZqkdoyN+GPUVru+NMiLRPMfUFundC5
CpdrZ7xTJZsXf9eaRMJvB3446hofoVH3EsufES8986u9S+o3CNgpHg6MTNrgo8wZ
cpm5/h4oyr5ns2qIS6iX+PDa3AxTQdIAeCZJgljt+zw6bJOE+VEUtFeX6LYPlMy8
r+p9rVUKDy8gSeptw19JB/JC8GRwT+Y1Woe+oLp49ex22ud7pDX1M1tMegDlEKSE
26RI7LhCRPYGykYNga3FCxbfuUrko1gpNT++9gYBl+H1UpUYPxI16Mbv9kn46hz+
MjQX5ivTSu0zMywPFtBQ+y1M2ZnbRPzWV/zInGvvqusqe9PF/zn9eqGECp5ect0M
juRc1TQIF3KMqAoFgVneq2+qpjmqcrG+kyJPVSQ84gGpxkOfnVnU0nLjqVY9qCwX
FI6BBoeqBUU2ojcrG8Xy9OZvc/xsfSjocCeFIvvttnLrC2Cg211iSBWVDk1ms0Eu
Fkh8KPmDHgJuIAHmBcd7423LtHan3LF/cg5g9XePyVBIBLOCnWDv1Z7fWT8w7lBK
VzYm2f+iaih2MynZL17qK8tNHAcO4PAuOob8c28Pf7zwQQDwknT4P8S1ja12CYiK
86yKKW/erBmSg3qFUqWK1nAs7W/r6RbhbT2gUUB+qBP+ik5NY0nmDa8StthPRumN
1WMtn2T2feZFT8GUMVv0qWKWY/Vwonj+PjeX6TArsIvwFSmUsksbx/FUvDFXnAG8
8+Vbe4QATA8UNwBPcaXxAl7ekAS/mRCb52trRFBV/fNNBjdbyK3e56y5MhwGo13K
MZvQCr3Uhpb5wrLD0hOp5S4XapiKuDXuaV3rvFOzsW9ruZ2Xqem2JcMwX24aKrbz
9ej0zjUL1X0bdBtSAPYJ9k97MZNqJhIZFNCoahRws8UiK/kdRGhFZ917KY+7NOah
kXiFVI2dS2pl6XrX3xn+BTa1L9uFA8WrlrAsA8MYVvkag0ShbOGGF3q+R5XzpvMr
r/RsnjhYP+c4WI3mkZBv1vrJcrfYEfU99CJ8RO9H8vguGL1fOM7QQaOo1Vw8a54T
m4RNm47U2G34yeOM3HWBCsyRTjHTAN8k0XzH4vQ5c0YzK65ZVfjhWzqjOaCPuqB+
ybI3m06Az3dJfV8leiY6qswb4qqYcrxpeIUcyrfvu8W/WjLfmikuWywJEEynY/J9
kYKHyPYpdLyE4e9VUmpdcD8vQwf+u+XV44GGEJeXk6CmDvRA6o93XX9V39GF+Gvw
lN4HFL3+OGCqMJaCGS/MEbWeC6Q+eu79C5jFgGhD+ki5hO/PqWmrU+JUF9wE9R16
MMcAKFeGImJCjQZYrNi9kr7Vz1wsDUYw/bsHxpCrdqxzWM4IL9leL/fKpArzn3kd
p2qQulRotvyJSFRlPPuxYgon8I27XqMyekQq33/sONgMMAP5LMKDKpWWUpJj+3N6
QjzOikYQaCHxm7Ost2hCd2Dn8L1xIaTtJpDBuL0XqwlDaFiMps7g1FVUn6zHUBDx
W/ursMa35XdyuSFnFOSe91rmP3hZb62bVehOoAMeAdX/g/fPGLf+BqKq58e20o30
FL0LogrBDCUBwupzhlejnwyeMeByJ2+SdTR0bbkB/3V0XvnrSrutjTK/5RsIB0GH
ZgAOYWgLk8yhgv7R9oMTUEGNlXjpzScDifxkvvJzYdxYrF26+2DkqK/QRZJCibd9
2Dnw/5F43xUpz41cwqMGYHPYiuxFkF4TreyCUvpDHE5zirVgABXBlSQ/TLcl4pAz
LehGCpJ1qzgDljewrm7LXtQayJS7+0IrSva4LD5tNOIEg5Qix0Aw6zWGK/4olrtt
atdTh2s0JSg+/0w3SB4++wBpRUm5nHl/mluDuOsuoyQCNnsXgvVQ2y0S6mmNVbow
BHDxaTiZgRCeEjiM51vt3//NdeTWgs7ReDTYmW7zmCYYj47w0CR4PeC+5M+nZxsn
JHjocKgUtXyDBvMkx8uqlBNN+ReLOBxZ4ZlJ1wkLEqNWv+T26DE0+58Jp66VvLtq
u5uZTdg+ri1AOJ7IYN7Q5IMJexGB8zW63R8PhG9yBjSAualk7GziCdYzWt8/otoz
0OpLWGZEa/Dn+lji3fNrbK/ra4iwls1E12SRjeySJdb8lRwszw8jgEbecH99+lkH
BlyhYpGmVd5mI67/fueVrV1y2yBD2GH2D0iqVSn9ZRAN/rR7lWRBzN9gNJIZN2M1
qW42UOqxDNyh6y+zzLplnGPUVxmy+fJLqQwzmRN/i0D/9lj97znQcC6JYj7mre3+
iy9iej//DdkLRsE6JuThN5EFnAAtsXE1oPs/c1zhcoUFSgDEZxiq64ZjQuW+tEdA
RtKRP2Xx9a+2bPceS7Ld3sbH6vVLXCjtAkB2Mcc6CmaxHRkmxWmrbyrOMESyMfmr
sqtYM8DYIcvQN9E/fC4MZlX62P3M+zRhfYgUtwdt8tsp6NmGikV+IZi56YMBndAu
PAavNRmV5U+tEZ1QxmRM0yC8r3EgiSTyL0EBsqDXk7wo6sA7bHuuIaf/f9y45U1V
SlE5rPOgg1jn7aNRU73g7PSwapPx2TwS6Lc08dB/Owy+759/kN+p6ZCcWA91zNr4
L5GWJ3WwgI5MoKVHdFcHN0oxhQys0eDod4KfDmcIi90hoVrFv8z1YQnM3CilxhMh
MmAG2UQfRFKpopAxEIvVdLj+4K5S3jTmxWly99wV5P2MnoMOT5OtWy+mnQTydoHV
Ityxo+A9hISWr0LrRoH3Vg7rItQigy4JJ5j+MCev5ZZANc4RJ72FloHZ2LMvl082
u9SDvq18Qh7I+41oPNVXcih6dtc+ZRVeUskCzaFned7BNkGIaqwXrWW1gI/JRIbv
bQ1jptIuKsvP7H2fu/Aia2D2+/LkLsCXWvhn3SFMqKQ5AThZxeTe1E7JhK+10FqL
dcjiIHnMZwzkdnOYrnpMYhSKmbbvZe1c7EfGZs9oRR1fvX2H6F0izIy52iLAvYSR
+7Eu0MouCLGmmmMZ+7hwOhp7pHsjtB535HrcREsvUhwoNn7KGTYMowuj0m9XtrZP
bX14YqUR/QCmHJ8LfP/qI6sU2qBRky4n3nbX3BBrqqiPKJeAoIBW4NAfbSqfowiJ
INR6v5eHHXkl73iX7zYB1/4ArYXwveKE8KbOg1k1hManTHmiudTxmLuqp2X6vqRd
nzXvc696eZakns6JZ2VBLgBqImXAhZb4p7wLJrOWMr6rVFHgY6/9P3+iiiXOkYcH
xPlIlDmBO1wZDyemPl4gops7hGi0vAL+sd1lGnP6DlhzakfTAUFyRmbwo3qODyI9
nA2XTirUGrgA+i1MC9eELC5FSRd1RhWZNHIpQo7/yMuzbmzz76ny1xggI/tU/wL7
RcFbTwpDS/ZJfBlFYAvv0G5PTSMrT1b/FPtl94xXfoH6Cu1bcyfTIL1VXgSp9EdS
Xp0Ph3WfgrnsdRa/JeiEPxNoGp+qusXLLHo8y3hM6xfxHdGyjmqDMgXzD9wuIt/N
/DRNhyP7VKUxTbhpeQbwL/AWL5Upqo5qKoCZnVB620fLuvyuhUFgTLNul0ACir3T
Ly6xGLqmcaRY7JGioiO8HGjYfc704IEcK9tCSpXLjjOOo9WaL6iGM9wkfdzlGeeo
TMnxLZ/u5f7E8pPmvCbrNRkR5cDshmNB7pl0O3CeMe6sVe1+yV2qalvSlhjcufAA
fUy2hSfejZGqptkOdGP6JqtvT5yIicowXEvTqvmlE2j/aD91hw81uR/m8qN+kFrv
PGTNlr0QNgZhk2CrTIQ8J359rfrh9Th7ttEI+EUKOcmKcs1/ZGOsgCA5Kk9aB9X0
vbuHiINCXCJCUDOQ3tEnp3k+d7LlzK9zFvana6QLQQc9K5ijBdSMcLFLrRxS6lRt
M7ZQZWyitOJW+/ixKYSsAUVofqew0yX84gRQ4yMJ3pi3jlQElhoLUnGYevEl4wsl
H2EccvLchgy5LZv2XVZV8jaVVy2f0Fzmb9AjshMf1WFmgoh2MZLjjVQz7F15GFcx
Y8+c4gVew2uOIFo9ZiHDlLZ2uAbVAXlxXxbjJxiFi98tbRGI+GQ2dwkmAm+KPTfV
XqMR6BGbO9cntFgONwx6zw327ChkFnSYTYbVKp5oiE8prRH6t7o0gOIf+AVkXkBh
D4GGMP7K6x9YvjLrZoTnnTZcLFGRycTbIAuQt+CzhtJ5Izvjy0x6GlaZwRp6xh0l
l1fM5MuDEDpNGmcIGyYJO9TpF+AavR0mzQQQO2BSci+AwEtURpNE+qCqFc5ppJKR
wu0xfsB1WW6wCxMM3+wQNuD5Tt09MCONJ0C1Zua1qgzuLV66koSnYt81GlsnuOlF
vZus6lwVYVaiRomGs6EO9ODpZkUyYFoGtLsyqNGe8rCTi0r4g88rIXUJCBpJ3kGy
6Wo2tJDpq8RObVPTNwciG9tZHB7PI4TGUmGcVo1G6hdH4yniR8EoX7BRQl6fixOM
W0ZfbObDPl31hQsnS5/aKbaffpXIdVFpuiBsk982He4NQe8ub58THJ1dKBjfkn7K
QZVe/pUfmMVUH8MWaD3V7Cv1sV8TmEacensp36/MWQ2eorgfaHUQl2IvRTqEuttz
mZ3gBk/o1TBrCwYPZKhb/WqmeiP4b46+fyzdSlqOK7zupMsztKSRFrNvwh0ktPsq
I0pr/BbhDnH3N6Kaf/O6ZV5SS7ZqRX6KW3VRaNp/93Y2kdPobH+dB7/8jQWrv/k3
8rv3PrUa5CUIIiQCk1citd2eTpLss6NmnuGgCR8W7INFe7iXBxVx6gCslmt1t7GE
HZLUcggXpdFIqboaMCHk4cM9/hlR5HSJYyUAeG+yJh3JPe58QI8Mvjars3ocNzf+
v4i+kzCOJOz9rOmHgYcgMa5d9YpkL1V8UBj+HQe34U2v2hLZ0O4AFHXx07zOXEYw
ETwSGDNDWfThhZ3KKyIvJA1X5aQJc/fjiNmfbHDd2xdUJrZTGO7gYWzbLFkTg3tZ
YZhgQ/WhokhmuK86INgtZaO+gRPwFHKGJDZZk+7cgKnh43ZmQVGsCRNGFXXou7uO
fZLqtbqAKFe604XweRDLYUAiBJYwOxG2EZ8pHELMKum8veV5osByuYIa2Ft0FmDd
CkQyUpizZRQAVnOW2c7xNIyTg3hKrB/xufP/VTolInGZzRzX/dBUT6BE1bzgl+3D
fqn5bq2SAptnAxHDjsOLRzJHMIJfYjE8+/tkxa3O1SzgFYmxd10WV/Mj0bnpTQfE
Oonb43MZVhSPRrtXKDlR2SCHrqx9AmzZprU7r2PgICxfKikPOhW3HV29gtgTwbK6
cvNfyst1lGI5VjAdGXe1ebCXnClIeuWVi0ZOWlTYriNtDhWeuxYoFo6T8gTPuox1
mwB1mURbZRWgphKfdIMZjJbJUdf7KIsYPcmc6u7fD1ta5wq+pj6rmsPl7zAX5rHD
p0Z2rgozebrjeFvPaz4Ubohdr+vjMryN0Ex/MKCYWh9X6DSKX+9YdXf+vY/a6hsx
oEMmXeZ2OdZvRHV87EuGPeYTc/pCLioYczJn3fK0tWJqo8fqjFOe/azObsF2/DE0
jbH970s4oOVlNWPhkpm91CEwfxCyVKQOCQ5siBFw1cVP8z2L13YuHmFiUs4y8rak
o37dpfo39XIBQWkYmjC+Z582J23wjMoF1JVSYZB8YpCHsBnXDBxZcct5vFkx4XrZ
9z4matnDezAGXJzjuqmXBByAaC+YCuVes6S+Ar16VDClHr20RFI4wZNzPdUdx1dm
AirmjkdVlDhDqDJ1kjEOaov3i5zrCDeh0ziE7K6eJBnVHkJ3mSVPLkJLuU3XGIpt
5Zz9DTliI3xTm+gZp3CTAv3PphFxWqptRd5O3uo9aO0xQHcE0ERJLTpoKsHAKSiD
HSKiFEGZdRXdNwM2s9R+B9f0F38vI44+99cN00wesPgxqYVK+1pLZfyTRsAtJupk
gOgFqTK6QbhdLKYhQC/xlwyEorG8o9p7xYb9GdZZ5V9oCCGF7hBwEdvFZytFCDfD
M1KzJ3b9cFJ7bmuPn/YOZtqIKbrnlrweH5t62RXoyPg3FjaxfclDkX2zsHOaC9vd
y3pbXIYjUiEm1iD6mogNnddJb7TopJC2iKpctsAWduKYaJ2ctpsSMcajVPUie3z8
2/AwdNrgqRFD55UW14SX4xnRzyZ8aK8gT/JwuwaKIOMwq5aoD3FhP97fQ/MUk7f4
e2dSNgmAcX8tXziLGEAPTscLwv3Xd4E1xjBNxf5CgcTx4hDqhxxQQGx8uiwYY03y
b/AzZjV06gL3y4+U15iL1+UF3/QrqVnW+wz9R8sqp2PqgxWl2XngOVSxM1Kq3kla
FIpijieB+YvWxgxZZ3V9YKByHYrU7pYzbjUls9aTS0lZBBOax516D0bQWRTuY0Q9
iqamvwFaSDk7gQ8bj/OSDPm8eOudlzVhJ2JfT52+yqBLAUGrwFwfQDAWHaBst66E
AQKQg9k357HYeLjIJKx806AjW2BKvjXK5AtUAaTeBl3putvN3Y/bMPHKj8yGgBxY
SXFEAPFGoyJZVrs1eb/bxrcEJBT59rRKme8Q4F8RxISy4rtJJdmoDh+EMeJVA8Fj
6nDKleyp6YZ/Ci9ZlbBQBGJ48CS7LC9XyCQ5L9IETYcsoI7GjY4mdndjJVduvxet
b3EZuFnThUCefwTPDv0zDBMrHW5CPoGdWAF8bRilkt1/F18Hehv/FIddpco9gHi6
SlxLwXQyvCP+vTFFXt0kn4t6hlXMnwUzh2KFw4t4lQq8ui6vwieVCwgjgFnM+KfE
NARnndZW8JceE7NHnpeGrRRY52gaCJPL9Vrmxl7JaiosyKV/jliX5PJu9jUwJfoR
DioWrqD/D5DT+/VVN9L2ZdSi8ptQQDZ4XZrhu1/IkU9wRlX3XPnzTVe2q8Q2VNBF
jQkWO6lY7UHrmeZ0UTE6vLaUm5+59XP67LYaPwlf99OBtIolm9/gPUnpeDx8pQmt
1mfio0Cz0X4Tb8GP/WNfP+MYHiHH60ovPPsFCkLf2wKqFmUyxebyk8IDKmWgOTJs
z+auPss4jpHOVxnGvHKacHBfcybMwFl3/HeERNjnkTJdgNgqCAsiScW6WKqSlOdN
hLGqH2KVoUurXzZ3o0ikTDiKh0DoNpN7q8pFNuzADgeuEoIPh0Q2wMs6rnTSKL7S
KMzDsm1RmWZDJxUAb1u3uKyU5ZyV7mhTgNjiaQImL7tWSyU0kn1N6KEtqsGEEV/F
4jIG9n7U+U2JKUEqcw64VBlAH6NkxjzykiXSTb669x2B2rzeqPios8Xw9J8b5dOH
oYxfd7rfF46cpqQnwD4pgZ8jpBx0GUtn7EnQ69YYKJGCNN/GCR/mFzTe1g04ltdQ
dRVzQ3MAYufjY85Oy0kHOn+YEGTNT1fw3YoH1CvJTihAfduGyo0RHrRGMw1k99M/
A0qf63a02GgzdDpEDvLYw7BSA8M9rpDw/GoFq8bRWkq8D5Vyw2xNykZDx6R0S8OS
OFA/DOwBFaldb033JVoKGRoF70HMHEwDDQ5dX1EsfnGsSVUtuBsgRMuNhk8Uv9bG
Zzu4KYalMB1sRYesMzH7JPmg7ER7tj3hywLkwk3W3ReNpVY96hpkzPO3beEGxf/U
0UwzgYhnEONsd0rEZwOOHFkU2rqlXnEnuJeZu3K4Oky2DDVhH8/xmql4dFIDwA/n
GD4gGcOUO+DbYx9Q8OQhQjzUA7Cn0GtjkwNoNnPxbrJyE/PQR3OQ2ELPEy1VrCkS
ytVD2KpxrYPF8NbLRzMJnwozWbipfBmbjhcwS4cgDNKBsakTj6pXCC3pGg8TF0Y9
KD6WnGj6h4k/csLBuOGzG0jOtr/P9EsKnU7rGShljigrkY8WCKkAx5lhVIuYpdBI
wBjyDvCn+chrmKLXioI6xeFta1SVOHgP1Zo2AeFg9m1IsWTDVPUtRsQCCNEQPzmi
9YbVpoxI5Wh59XH6GeZrwLoDbFhmHI1yQVhM28fGDgfd9ey8uMhXz0qEzkCZj9a9
1BS/M2qPEmOosCNxmffBX0ceKVaE712LBLGUhoF4Tr950GS+KV6Ku/xueR5qD/Sy
SQW1bWiS7IAyfgOikGPg079zBP1jt+jvhc9Tb/hd7Ejzi0jD79U/y/HNCMZi7P1U
SsFXbB2sBCX/HPlG+xZ8vxeiaAR/dpJ9Rs5+4UvCMa8zXwwmUkrdt0yDYC8r/tDl
fSjLMGar8tuJ8oI0vU2NmpRLxFa4dR8cgz01Thy7MmDNoTiV3DMAC/S7NkWOJ1kO
jKP7YgFHmQ0NtY5RsNagXfT9sPrc67BQ3tae956cimBUTGNh32tWpLr3bsyApoh6
tVlvOq1VY4CqYVDBxB8YMjbD0c3dzL3pGOka9fD0j/qZyxuaqu7pC9IKzrmtwjfG
UZ/RX2YWkOtJv/EL/yKGbgrhXQEKxA0KSxlgdGiqIkr2nIB520iEoM2P9Un3nOAU
+kgklEYoOlAqGKC2nLWU2sryE3tbU2mKHoCmEmN2psaGiVpryUzltWV6LyeWHMkx
DjmSJSc2o6nZ/6o9aB4QDXZxR8bH0La0Frwo6cNvqG6L0cmgx1EnsJJHG4fqtpHR
G8DvApRtSVHNkGxFu5ztuT/JqZMyHOn+Szcu0R60lMuDijVMzb/gOTa74KW5b/XF
fPxSNLvVS89wP8TLWfFz3LnPO40ZUe/XRKbr1Dl7TGyHdEJVOaAml+R29t3EsFiw
OfZ2e5KrVp5Kb0wzBczAev7LGE3wOxOVLgGY8q778ENKoouwg1fLd65fsahl1DvT
ZVH0GsA72uf+kwuQ6VJerTjIBB64OzDf143GqBPK6hFHvVYTfaa5/5t2Zvm0yKXh
3L07Ke0RegCtsgwny238gdW0D1zBfhjtPXHupFA8mYdO16R/gi5wxtW6MOTvJ/Tn
pQehHFm2cVzKMDZxTJ757mKuOzCmrFBVtXSUbAu/pX64J1x20HkYtosk8dgJ9M6d
IPhF4FAvxv/PVJKWh1lHB+wIoq2YcDetp1hOl5EnX1j0epAabKtfejrifwA1OuVu
wtjccAVdSZ05pTkrsrTzAYG6hd257qcdlGXd1CUbKETtW0V1oIDa5+6k87+/Azsn
W7c2xksv7fco414mQeNNeQ6OSWHpMrTx4tAyWWeZtJsz8OKhoVhQ0LFDn0FDrFT3
z+nHe4WeVdRh8useCLHlEQIaanztHu3SHBLimV0+1ZW6WjIpvgqTiqjCGn9Nw9L7
2x9OtdB6/EuGRveT0QXm1wtkZCpIOVDm3p/jzSLdzLNcte56AJzJQeGUK0/JcObK
WZJWfVH3jymFahn8PiM5DH9PJ+yoItytFQeBGxKRdblzTbM4btY0BVblOyFDgXiK
3rfy1L3G8rwKsMULEpnRLLWMcMqk5KAdczXpzuWCbn6x3b8QqR/TwM0hChDTl+KE
6BJ8zsFENyn9agRVi3H23+D7b0w3qamAmE1x49yXBtvi7Ywmz6w+1jNhOTbqs+y9
+JYvxYR/zr35wij7KjV/mXo7Pv1QOQHPpRD7kxps3+x7wuegBXom9wFD8Wq9l4nb
3yymGdXPZdKauW+t02dgJZQmOpxV7nI7t2fP0uW5phnPEYPBUAgWbBLC9VnlVVFL
OxrZY42F7FDRZmisG5Bjj8rMFvPxeDQNI1l3qGaR/t/5YrjHPWDrGAVJDPBq8wgl
1EDVMczvX4ZzstuXNjc6/05WYjDtLtTE035PwvLv4Pm1LRuPm6px2UxtP4eca1pG
1KBPKZ13Nb+OZcDkPsmcNAoH+e+ymmCZ6P3u0Q8X/zr1ExO5xHrpngavsRhId258
OF6lcyrQt5pxN87SeRorrhZwrteUB/8y1+NoKU8xjKuHseL4zxJtZy2a2Vyyk2qR
RXrKffPENyOxqNASZYjTrflYHXm6ytF89dzw7Btantm2DzJBf/4LbhEo8fr45+8C
exUwYGoCZNUisdwhHqpLCXsr4sLUxSpv4Ui46SWmwB0sLpeovt9B+PJxc4Wb8RlO
ql/mvIU0wf2+2bHI3wgXsPl/+h4/ekNZ4wBGwrTmNcoHiD+r7l9EhYHLLihrZDG8
EcmC/zeDcs690FoNiOUb7xkzk0wHIYLltBvWbRkuX/qMnoxfHZAzKZ43IV2wn+Jw
8SUV5Wfi7/iCnu4s0apj61K/cJVm4TZ3mu87d4D0brxRsBuH3VcnT+JgOfmDuM0W
z8j0cGDoOGrD4ZU1cTY0qzkTO9flke+Q9DJv2Girzs6wizdqH8VlpVQ9GaSO405M
L7e/OooWd6euQZhf+ZS0KBIes2xSydUj1pgnXhMlh34ft+a77xE82cMxlHW9cBrc
sbzWJ+XXaexjV1RI41eu7i+D25cXCRSxa8ZHS/6OvNs1I+Y5NyvT4Cs+/N6DEGoW
XJ4ryEeNPYaPaIOSmbIqy4JLyCgyKHgNoDPVWcjXA8HBd5PpXAcGhdjzAa/I/POg
OzpbGKhu2wNpvBMlrZl3opm0P8+djBbg7fYOzzlfUMtfLUIG8HcXNEA/vBu5D/G/
PXdVl/R1gFYJGxUzzl3zcho+KuRWEtYBoLWtvkRq5jQY65PJjFiU3re9hJPoAvIQ
a8fGuQjt2HeNlPriDRxPrq380Ut3b3a3CiBK/ryoLByLiipDLr+x2qlkHx6G4UL2
wDvXLN4eqlB0ijWykI1/B9NVwlLkNc/IiTTcn8TukPWs3jg24cgqs1z66hiWcKh2
/6gYBkn6jp+Lz8pcFxeU42C+9ucFpBGKy7zZMisSSsSvvGjEq5XmjV0lPbqZPKi6
JD63VgCyAPagsLwTEvVpdnQxL8df69EBQmTjW6B+l7PRs1oqGojWwrKyhLs9DOj4
Xzoeio0XUkBC9dNUQTinLp0bOKowQhyitcjydEsSkuZl1l8LBETGv/N5Z0aewG0G
e6DPmE4nWllvk9mob9iW9meN4H5dkGcPYVKhluTUCKJ5Q+SA3QPzqWhsLh30Q0AR
9t8k+IsXqGDAekxcJxwXjBi6qZLLIal+gBzkiBdV7plSNN27a45SoBl1JjQnwQ0Q
H382Tk71IBTFdo8ub0tnCMFr/RzwbWWmJiQEauaahHzQ7ZDNWBbt1NmwJcLpwx9A
+ypZDInkfHYub/L41/lN4FaQYbrSfexxCmtYO+811AaA1C1cvk2TA1VGlWT9nZxy
UmdHVOaGeElstmcMAFo2bGTes3mSQ/IMbhipSW9a/GgLJ6GpFPTTjiILewAL1WWN
gmaiJfgOtn/xaXoogodBxKEwexCnWeOo5Bzjgm2c4HQRb/nRAwB1YxHASv3boZH4
NIvgalRTRg1do0YYd6mCbSBvHWTW3ymozEUMAASdAzXRtHcrhtS+Nnri6Lp8F5vA
IZUZpoGND0+YBRPrXrF1aHTEGJC3BsLM7+tHzuVhVuws5peigc8weTakCAxQLWKn
Rq/kcZTKvZtJTjIC+ogeAuluzzLH67uGmEVawA0gZJfMWM5bl7JoPIZnofyEX3N6
nlAtqotETRZ4pAL0RbNdCreS7ysKXnnj18fPPvQTOZ11L1fk1vt2PkE6E25blOLy
Cbl9Nm5EoZZ6m6XlNiMnsfxMCfcMbNq3QKh9cgCRa7RHp9jnf8uPilQjoGTZL9Cp
pBdw91TnH1wSHoNJlfTuk5EtkbzuwbTPzqW067l18COQLTx2TIM3jhhyHQwbsnPW
oYSe/vVjqyO/jQMfKlT1s3lFfwKklinDGqQQJoEpz7vgO2ILxCN3C9umPgXzoua5
LsDepfEKLu1YO6lfW0fadxw40d4lWvRsgpeqcUWSuf+MANHM/xUEhq+W5yjsZ7+M
MRSpnwlo4Mv+ooI7G2f648inBuRSkpKSr/zA3d/po2Fg3rBjctJj+a8n3QTcqm0L
h5hmuPXWT73G7RmMEbf2GNkEcd5RJILqq0NXgKfbVTJD9A/ptADcflH/aV6FDbgb
b8wLujAKEP1Bp+KATdcEX9WaLOyAk+8NMA5jEDs+LrJ7HH1o+5kbbUu7gk6Zo7t5
mdkjoSuRfKpiF4UY0vYnRSZWOIrvhhsfonLbMBRwMUmlbrVuFj1tOUjBz3n+q1Lq
3wS+t9zKNk2E2VtwOkECNTkNW3wUEH+xK887UjjWA7xuvX9dRz9qAe3wewzJVmSj
I4sSYTn8fOyO1A6OXNgv+CjTQpnCxN0ELJFnxR58qozVrVxPZ12ofE+qk+gqhMBe
tmk1AFkkx4qGlDHlls4G+6ttx0+tLvU6OfGTdv/yEpCfsMpC+r8j/5VtH7LX1USg
PZiwz5NUv/xLPOj/t2tphiO1b2hn9ygv/sOeJ+sElcVMPbbdgrVo+1iSxomcjktz
iM11EuIGjdDhNgg61hPHJ1ocvnvGVUL47rLTjcfw/005j2omi36NXEgMboj3VUgV
m1TjE8rVdMeu5GROHxmGoITEo60wD0x3eF0zURlTTIX+oVWiX78M9RlWxKJssAFb
1BSWpI5HqeerbMqxEYBezqL8881ns94pH3pBDrDnUzsq67H4GH64CqLiSFxBtHOa
YJlo7/MErTkb48kAI3OzOkzLYDyKUbRF8qJzVd2hStpuV/AxVesZGJnNzVeL19do
EOpJoE3fKDtnJufMAInw4Gd1/dHUHG+uJwb8KrSD22mxc27HS+CvrmOmHzMEodGU
0s8I8vUY/1mKIYe/v6ujrhwlQRaPeQfv1d3dW9TW0lP64WsVYom9YWWzNN+5gwl5
jUQOgq4j+G1sbLE6OYOF2shkp82YjzNeyebxT98m8o6RJGVy20OnZ1jJD6q/AXkp
FN1tzc0Hi48YbS0VSjhwPV7DLwDD2ZiplfofcaIOTi+AqT3SWZWNeV4Bp9KKtBCt
teBkqxP+g6/g5by/Ik03lp4HCncPDaKRoekOqqWcwVRPIodSLIEGw8TiOOeHuy7E
x342MSExSOrQfW+NYSKIiXm+a7cMRR2IATCwBNaigOX9SRphOLpnSc7bPebQ6cu5
OUnsQ1mnSmUk8o8YZBqWPE+XpPd2p+gefeO2lk9L1zJ6SUbpJroImvHpbWfNClRF
mpDyvffQ66kIBKZzKAlw4JMuSvqhLwlzHEloN5k8bFVIWPM/0+qSkQvIZj/978/k
mzLzKWPkshZ6oXk94Kbk28OoewM+TFJ7lJ9tAwnSqg9tdRKkA7TQENyYirP4jBHP
igtoCXwIJhERq+YC4xqXsahPsOUApo+I8CknROpwGWGnBsR5A3lxWWt2guPk2TsP
h+X7VihaLBiBsNjehpARIpngmmPfkl5A+oL7mywadp/hsga4ZULlpwOwXuN9hePi
6YTea/K6EknEEKYhyvvLAU6upg4Ym+np/bpN0F7l3l2k9QHePQBNrZkgRb/rNW5M
p7bbU4WhWVLkfvW8iPiN+xb5QIbo2PIsTAP7rbrRUPO3YNMEzDF/qvtDpnvnl7vn
p/HufDt7s9ZE8z2jDwjdgp5yq+KxN5FfN/F337DEUp7sU0dZVutBSeU0pv5XYpZM
rNRDN4oJUZLOAEP7iL/ct3hY3q7NWnIytEbvtRgi5yxkotNrlIdM2OX1MMVZ2B/C
ldm0WpSCA9qRGgzBg1UHApp4FILVYY+Sw/1h7F36hbEHYmPJUPkAlPg843knDH3G
1euQVitXPWv318yvMiHo5BbQShEUA0ZTCrHwjn2cL224m4FkHT2GHJkEKkYmFf4G
BznkBfdte02VIly3VCNsehFHE9HoDWnWIX9i7hUAg2Xye7RM/8BRd5vMmQtfF1Rg
W+5etWLeGKCByAOP6fqhRKWo4rw5q4Ud44k3uT34T8kPFgoYnOCJUXpZ+9WIoK89
WXw0yfAp5BAkCY+UG+f8erd/1zvTZLI7mlcqQUuv/947RvK4zVTjrGDlrs9uwEnZ
55HAnGy3sHA3XnSLRrZhdJd/RO83g8Y5njTQ1LppCNd+rMvyTBZ6NniB3QZnO/2A
1yC5inFO+Bq8fibBlPwFIR1CirptWduMZs8yOBACu989b10Lp5f7L9JCZdbajv0z
Jyi7eK3FfNNYaz1Fn/9pqMmbBqOHFg30Vjq0T17odddum6+uoLzcBiKAYfr3duKi
+THcXJOCj4SSvCIP+R2Ik0z3cLt4c+a9RD22xAnP/mDvR8UejaZCBnSP3FpxlR43
cj/Nip9egzDocIIn+wepnkRKeuoGP70ut7UdgcI/EbKnt/dSu8Jph/sNeMiSubFS
sWxavtsC1tub1MAW1L457otbUzf+yAAHfn+EPYDk+NhP35gwDoUZUs17x80E6zMF
On3x9vQAKv9V59u76VbTOxnxAqrl4cNi/VJCHTsvozrm7TyNxAxegScMHLgLJQOB
KkPlvRIt+idRMQ6YXIVOQ5c4Kkk0GQDeIRSOQIzSuXrbaFGkqxB97/mXRNKY+Rjm
BwPy+EluHNpcu1+ydjSKyX61d9TJyzyGwqyk9AzTSim3KvzKBDeh17L3jZw3z4ka
65frEu6pN2Y0fT+e1CqRMX2w8YPGB570gzHlbRloqx/IRXguxstpZm0uIaMeeZwR
3Cfuwt8EB9f3XBZYRZfTACum2GMiPxOuDlEzl7K418JoWaliW92LyHSCrEgcpWb7
d/8jEerhLslZRPWbvY8ECYGebfVIFGXTfjKQEfn9Nb4K1/PoJCNrM/ZQFiW0auDP
RG6Qw3him/umalU+0ipGxSJ5gHXayxhwLz5fvkY/7jB5eWdqjOqIATaf145Fnupa
4gyz3+rhMh9s8hPTWA0U1iyPA+bBatEE4yEvyBo4XM2R2b6wRFwmWBhUAUzCQcBH
CKG18qdNoxg5HJvZHglX4hQovVQfHnIhFWkXv4FEQpR4ljoGM/t194DboHGGKkJA
OqPrkanQBKrBrVtu2Wh8Wik3kcF/BlwzYOVuf1CSROohfrEySrVItQlA3LtFNQZg
It/1Ssfb9ozT+F2Gh6AIjOIsZ/q9CjK7yPysyylsNHI09Hbwwop/p21veojyk/b/
RMdp6xI0IEZGrd2SXgTm9YeMfpJ6fa13QzvzcJb+OgnhJ1zfwbF4giyyFgVo+qS1
p8G4t49AC4AOMTVbB1wV1fdxDRM3XNMQpQrb/qPcZoTxkb5jidAxu9XyyBmgkbxR
ASwp2ds0CA1ENSm8v6onniL+GYUYXaPnEVSK3rISdxZZRAb1HI+JzU16prXVBELZ
MEiHZ2wDoMQaI5l1KGq1VldDparkWjX4oxff3EXI0YW80QGVMd9MsF1/TQ85NF+m
2axKhzsdo3xxBehFdNu0ATmp67wthP04N3oUmrgrUprGIpv0cmKgkmL6khM6vfDW
yvkdoY/i61o3mxlanRkmU1ohazSqMAus6IAKo5ZDxd3iXVj4W8g8jdFTHZijGzE+
jrCE5dQ/Z9WtRdlWijg3/8DR6YORO9OssH4pihU7QVcszvhfXcseVCqkzZD8iMVu
mcrGgfn81nzHx0SuosGmJnkkm+MJqhtZaGrlMw7eIVuTyuqlvzzTvhfkviUubh9G
rbR0clLKQVPp1CcH3iAlZi7L+ZKhm+iEjg0/rt9V6tIeC3n9imRcIPgZXXRXMer1
A87G+3hdU178RQ/oi4MS6LrqK9KM5PYfd9D1OXUlEle1FnO1CZXuwrQP2DiEh/9W
NImoat6VWUWFkIgcYWaGPUfIfkeLuRZ+TTnPbk59+SE1mP1XSYFwti/nRitfsiWs
Wu5X9sWrVj8wVBaaZI2VO09lAwO+LRf1JoxCpGlcVUcEfizcvvH+KdIZoajjL01+
j9pGCeGS5c3yPfy3EjZHjN6KutvAfIMcx3Zjix0kTgK6dHGm78rUmR7wRD7K7us8
ns1AIgmkzIx0wgJ8Gvi5utbAB2vMPvn/HNYsHrolxGSC9fYgaOTF2ZV4CCSPfXTA
99lFtGxFVgJn8DR7Xm6wUt923PfkgPER2FThCUPdrf2PVklzW9G2RRdx7BZuUBfe
aczY1CcZXQrj39eOg+3YmfbbJh0NgYV7OQPrmSnZrzIUtx5k34RJMRR9w5mwdyyR
aRVEsjCku41HiRPxLKF3iD2PFq5cUSjfl0Rj6xUW+G5Ka75Nq3fyE1IHEQdxaOJr
vI1a4Cwo6SZDQ1Q7KXUDqYG3kX6h2GX8IUxPzMoEJEZ+/V4jpEsoYYQZa8Jxpci1
FIhG3PRbO3m8pEr7gjy1z4QBqvwhvPt+l/vQ3/eZWUgC1A+aYkqMa7qRbG9X73Sq
hiQSPXWZy1x0bFavLDR6WrLFK1+nQam4/m9ltzr1I1TDOFoi1SLPrWGmo7NoV2T3
SYNIZqdTrMZlvlmM4nCS5wWIXVnf5586m8ppV2WwqxWnY4kD3YNablEw0iHw8YMX
E0Sdwjgkz9fitpsca0tJBlhph/6zQvbpSETxs5Q4ed6hmispFEl1B6mh6GgQbxgl
pknSoD91C9q+52gPTS7gGfJ/bxK8QJF4cc5iIo3QXWzEYJ8pNZ7P/ZW8DQXpl8D/
RSa7rSieZrO4OyPdGtESTvmxCgA7lFCiViR5ehgVMWTCbbkSiEPHWV8JkwMtd5Io
LuBVRZtE3pVy38rwUWW8qYKSRwCdZ/FNrJ14nPegkUkMqqjeJx1N6KDk8MXuctE6
eEevIyzuZxpTs+nvFUy7QhW6xHY82WRiC0xKIPKr7oPmNBJiVgW2DIFMBu/XQcJb
gA1rGQtYRJgNuzVJ7vaLUKR0uAODAnGiBPjVShUhKqTWt1Iih7wFlI7GVeiTJfz4
Y3f1kCM1DXsUqjV/KbHv0HCkbEpPZO1IbP0RU9Tp9DJf+6FTQ1miUJgfOugUkGOb
lkf5uRTnSSX92C36RwkrL8Qb5HEU4fL1CiP5OVvLHOJZvM5kiwSpL+ypWwGOehxe
7FQkzTxtlun3/8DWNDWO5yoocHpLQ5H5muw+97vu8enje6y6x2CVCerM+KDYysoX
RmrrsyP2XzQnMNgTc5kY1Wj81xTAzUHbooDoR2TiQD+uF4B0YTcM7DpAJWi4cv4z
zyjSrdXtRksI+mg8uWF8a5LH78KfL0mSJNz8M3NU/fzdYac2PRWkwQUD4KQEja/A
1naj+9kKulBxUzC3XFb+Vicuqnbb5p0uhQ2esObo9woiAxK2r8+qljCac/gNQZ/1
TK96dIMI/aki/gvewFefAIEWZ+B7XlWLYm9kPN14saKpPPs/RGa8qaMyToHAdZBh
+v/jcBe9fQ8M2Z68jmYveZAKXbNb9DqPmdj8jEItrfaHVE+y7yZYHh5lkfStI9ld
mA4u3vSS+qPWTsCV7juZitFQnLzhFuNOTtKDASripNREzxjqex055Uy2Ol+H8b8T
W7a+YBaM2vK7mJHiBTCwQfAKnag/wr5K5l9ynAvKmNJ3kGP/IL4HQ1KcwfpT3Bw5
XBaFytDA8PRT8v1tvSkR/PqNRBMgWJIZbGTPVmoeupWXrSFWZ0KmuXmjNf8pVKp6
vdIpL7PtLqRiSxTc9LEXR2mTX7K7F5iR0VLt4lLBYeTf6N7hHO1D8CNGtnTIs0VZ
J2SY1Jqfu+fO6kGuKfv6uqGTFofLqrfYG1zvOiWRSEvj01wf0SZxnSbkD3RAx8sx
phM/ymno0GVKsdYICnSQfwgReqK0i+UbUVyscdA9+xkNf+jVBcDTrl/RzaOUT2sG
JQE1dEZnbvk/Q3WH8UY7XjYfzAdJPNA6es661RbjdHcaFxtjdE566Q6Utiv1c41D
AQhx5xx9dWqkCaHEsiHzzr26ap/ijwKtli9aMDA02bNv1NMSFErRDGRvpRJfJmAt
gmMbjj68R3rOPXsV1JYETL2Jckm8kwV8yPyaiJvDW6c7Y9aGW3nA4GAG4no3W7qq
CbHQFenyI3zbRv0IUxGT4DGVPsiClrHr1qnvvLDbKIb3DRwmBlfqxotuyhCjxVDj
nR44s/Hl+iYcjhdemU3gKv2edGwgCs9DXN4WjuVGESGfKblji646ylXEctFSndNU
Xoi6XUwJzrLveS6iF4zEE8Fy9FcWHia4K9H6ASncE0ILMbHi+mNl+OJCarWwj1+d
oHnmJB1vBOwMdS433ietJHKexMowsG4szuCvZJH7vz6VUK4JavQ1GhzjFDp/uurD
6jhokeMJZuW6vrp2GS+t+hCkoSfvBWY9YkSCH4LDoCQEI50cHB7OU6VfaSqh7ZoR
Bb6bdMBMfdCaEU7GrIqORTR2Ocooe6c6t8q3bzZ+CoSKmQp7e6JydnapZBix2B/K
carr3zk+c3Gad+Qz43QywTXbxDj+wW0SwMrNhrcUjFP4C+1+tFKaWmm+OTlWBtgg
8TtiznKk54r5eXD0Y1AWS8QLjXyKQsohQbDWFQ5j/f8wKOpqhnifrMRlqnDrGVEd
dkxM+4XWLC0gMVDF3+rvDrDgQldeQscTEkUjEjCkTEn7PxO0L/dCj73UFD0aFbIc
N/gbOl6D6iwYW2w1Cj/bip38lKeOk4oJkuVus4GeZ8olR9MKARuImMRxJ++VhjCp
lfdVt7TVaCNTB7RrfcuihYAEOm1ejCZyxze7wGZDkmvfjsY9OuoexscTDPXOYypF
WQW2WBCWl3YH/4MFijNTFxKkb+2z0DrPCirZBbyUQutQEI+xvHH6hS77v7Hnibhh
0z53WpIIPnbR6VsjBIXuFSVEHu4GyEBgNJqRPMZbz7zqeist5YiPsxuxe7+898Y0
duFNuuRr/gsSo0W7g/mUoXhKoXjqofasQrWUGcsdMiR+x4aBCOJ0U/Ax/B/rI6CX
ADd8L6SnxPOv5K7yzQCp2F7QXQntQWWLLQ8Tk3h006Ekdtw7RD1A1b4wlsiMmrgH
HEwRd264N3oJwGbWb2Qt2UhfGawqbAVLgx1E/zkEY22OkdpNJgZ6wF90nOYzJiVT
FAcgTPR6ysQhP1iSEYUV1KUmwU2gTwsawwM6vJ4Cqr7tmv4g9Q8xrWWZjE/vB6zB
Nj9DcAXJ+mnWC10NsDa3EtPzne+3xthVJZWiOBP98gqJequcgXwTwbmKin5EG7vj
zKFkvebMBoWbhnm3AIsVE5KXbPJjUmmILFIracPvnZIiJDBlSSAJGdOzWUCm+zin
UohLhEcxiovA1Su9+iqfmELGfcJFVuuZHuUb7xltZzlFm4xeEdapz0vG5jzo9rAs
5kNZ4U3SnmIR2m0o8XJfJhv639SGk9Il2saozWhzKmwx6gQID9IQ4jjoQ1XxpSpI
KRVgEZewU+PTJ5PgwLIwbw4j7T+KGB0DA2R/5WBJ+Xkki1YbrBniqOo5owGNeBaq
Cc2eBIfBwhqzuUT83oflv8gEhMDp66ttMYPgHHidVH2n9zX/L1l6v7KQqLnOZGyP
J8cCoE4d4ljquZdP45zpBQxtxNX7ktiXSVOHro3MEgogkPTVpu4iPPclV4giAG/L
z9Vf75T9tVbv2OE+/UXqkSCW8t5sr43JrmhCTqDY7sDXkLSxjQIIz8iT2gPjinZ1
5qz1TDNccfLEaKx8NjXmJpTDNyHnlPn1WWt4OQW28lEWPngY6zgEUUc5GaqLnHSf
JJfkfx/FKdXWUV18QofPiZsslmX6Ts4mOQSkwpbcKk69mVEanC6IdRT7+UeyZ9Qv
jTL363RhUR1e+h/H3RiTQDom2TOexFnIWirXYc2xwN+9G2f+1LWRD+j84doVSsnb
JfrvUhpSqp0r2SSxTzQHBKTzgzrBk5BPny0XF5BId/Rxf6Js4UMsK38bpNyKmMNn
5OegqP7B2wzumZ6BEYwnmeXlAfNWVoDrqYUButJUGN6HOufmg90AbER1ENAI2nVq
AurwOm5Nuy48RajmeeGD9yRlr18uFAYylqWM4bvO4ggdif+EGHrvs4jWp2pX0418
J3iDvxkg/5i3b206E5nw9HJifKpg+cnFHWW8jcalHv5qTNJqzLAazt4LCADanirX
DiaY2NA0QgIr/6VjhgGsjDz74VuSzL9qwrm+RUhLwTWEcR2eKHxzhRD09n5MyMES
v4lFdNfaj+wcf0IZLC2oojzxFE9O3sbEZQkvyyTLDKcB9bNlNu5DC3GnxICgRbxp
0ZHM93mD7JZO/UAaF59VBwJDvnFQ2nbqMxh2KNwFpQXtlniezkGKX63bIKU4dm7U
dwhG7/XodRt1nBYLgOvVcNJcUcX/+9cX8gUB7kE3Fn7Dhg6czrSMoNMy/LvWUm0k
3Pte5I50yiEeID4CoT5cZ4cuQd/5d1Ne6isN/xDCnSxUgxK94EszGZn0r9pVsDV1
4tVXn7UrLDjDgYt8m+UKmWjjrN4es836ny6G3+h5Uje1XTgbwoTHTXfsl8BxU+V3
buZQAQLFyqjBPZ0M0A9usPXemv+oux0NBUlVnyt5IV1JIyseQjlPKW2K3pSMZ6ec
F8D72LHHXrovOfxwY3gFw4KoMwM4JkF6HGqEx4pgn42igyp3fejnrv2bHvavfEIA
OelA+ZEZCWZz4+vkFkDdexqpiSAkZkRwBvJdKUpM3ESp4IoXfX+xDQaJAeFNHAlf
wgEL6AoubVnkjhJnIHkvQAMYIPELTjNfrNt7gAI2WChRvHg6ubbPo6oQfMHIJCoG
TRTBypqnxVPzAgPnhRAgaq9T7YS8+pLV/MSAhwnI3yPSoRSxIcGh3TryncWfbcRU
VfuSLUPdc3rtYStrnxSSurFxBM0Xo1jdiD/2BWgs0D9EGg5t+OddRJUPSW7TMXBg
D1fsw1A/f2xCNzIXfrZ/KOlR8wlpbTfQyw2uH223qX2eThxZ7tAwCjmsETaC9TGb
oBiQ6x/zE/wg+nIsEq2WKhFYABvSsjDYFPArHS0+ejz++b7K0xb5dpNbvLGeG7Kj
pBHKyjgth/AUJe23nvqRuqTY9a14Gq3h9TOnRpSjh5STtCOgKRMsQ9XiUkTa/gYS
WqC4sA3GB8RtRMKqnKAE6wbOPCS5GBOmP20xUIGvNHVg4J72d7hn+ZVzuQH8CuRp
lab0AhXP+hMP2pV5uKzATODr8zJD7/z1owabAz75jTTY+tIaRyvz6OSX3SnpE1o8
tZVVpKC535pn/36Ct4QMy2XldwSPwNvLXWrttDEMZHuDwJFCHOVMSv2H2QQs/Lj0
A7L7swFum+1wW6OGXJhuceqLyPQLkZUwU6M5VfcMwjAUO0hOxbxg+wxH2PO3Fqil
taUrkjOo4kJgAjfavEQjSOWemxbEiJCmZhzXcGdrXMRFKybvA55CZmvcnA4Frgre
GFsRf6SncapRe5H/VB65WnNo9pAYg6MwnB+R8DzPnXtWFZ3aVmlhI7AhGdiFX/uU
bsgLKqiaBj2ZhiXGZKZsrWSngDA/GuH3aLQVy+hDVPQAp9V80U3QotfQTByXGN7b
2ByvC1K+Uf4lRmo+/TrIzQ9NvkU8yZxDpcAxNBCT9unL9N31dWrEKZBtbZXEzpIt
Va4Gcng50KBrm74NsSGcboG23Wao/BEM9VcJkgJoPh9B82kET604w1c+CQ397Gwf
PRIqA/gYNP5kQIjrknRL6JMHA6oP9Q1lAW16VLROte+eQ10t5C4vR3g+VPdhnBhB
FZr1xPtJf1FMalImjbgWwTYJgZ+bSzYf8AKFZBJmMINzUDSiPzQ72wGCMY5mXlZO
R66+VmCo8uJCCxxvzpZY97yDq5fBl7dEQjDqBoV8U08JQFlrU9k2j2qXzorJVuMr
Ep9EEl5v5njiCJKhWgXJ1PZjC8I4TU5/1sxh/Es2sgi7zINWopaWonDW8nal8Yr2
rFNF+Vr7fcGZgYsoDHs+nESCzFn9c9ldcrS3088iMgQJ9R7dSm2mRPpN/iidhS3P
rriPsZ2WLT8qXq1R875MlU62IuaqhoP8epbawoB0X3+PUZo9UJL0WSTHwNhEMbwm
6Y2QRvRlN1QUBWwqUghj/N+wPghQpGJHy1ASpHsjppMMKBVeVU89F03NgVXiI/93
5DhJfUTESilMPLh3d86URVg5cFsstF6KT/TGPESeeFdouXxjMTeF0io7ejvLSr6n
dyjeTIf4GuyCxesbM1T8MiqMje8F599bbndnjJ9n5eBoYPtTjbENqkAr9gbRNYvk
P++/pLhkxcEG2P8vAXwnwFTKbo8Abv4bT96+27ut9FrpAVGgXsuGdUnWAH+pQnnW
TFsOSY6kzoVJN75xZCuFahVzDQG1+m+z6kdRGh7lWFj/aGUwhcL4rPDkLkivTWu0
iDcepGQK6LR1LEIvAIAylw+zsDtTkDwkyOAju/tX9V/0XCBzI/w3WbVT7OXQaw+l
ktvTHlTpgrwgvl56/E2SWYoVJNnF3U2wSMxod3jGFfo8K+zqtprKWCRq8f0NY7JH
BgxiwCfP0PzfdGxc8ZsLYpn2wZKbQv/Eigeg13zHEb7DleGIdAJ8mTHvh67cxaby
jLa0NjKVGXD3pDVkRcQ3TszbJWigRvKq0VD2sMb5hxe0D2YAFqE+410EFO3bKtYI
Gdzk0PaK4UIUh25FYlQepKcCLOq/Yv9XC+NYE5MZVX5wEDUZAgZXSsv0dzlpjZ6r
buuXpVmQEQ0VnnocKbnWIncoHxbTxaN03Fd570rUFcUx9Y80vtNpFYfsx31otZj5
yg3i7pUGldund8/KfJQ7p1c0c1sATGM6YiOdr+gQYrqyckaDa+0m1WxtymBFyH3h
QsQYytwrc21Rtn1RWJzkDUJfIdtUSL1oQ9I4NnPMcKXNZIVWsRvpWuIBMVdZk3DG
drAEq4VBK3EHaAvgHvv7OneGR2r2A0mGyvludqRVp84VftWKryEliEtt6qpMcC70
8LpHxFK2mhxuhHAuBn8fouUw8tMsSHo0wxblFbpG2HsIJd8PHQow+HB3L1PTPlM/
DxlGyx8v8Qr3f9CodbIeyoXXAbUf0q0RZZ4lQuOYg7U52qLiHAGAphzAH4Di6gAs
3V1Z94zEOyKqbxNpLDSsSeZzEdELoC5D5+lbWmkY3Xfw6jzL6sktllLMaoKzoSrj
HSUGN3jEDIfG3zBmrbwn1l8ig84IIIgtGfnW+uaicriLY7evOd6Ea+Pwt4xFCybl
q1qJY4To50CY/1me6xnnB9hbgADSjfYuW/fjKCowznxrFSZvkrXm/CQZvWy6ZKk2
jv47HzgvHU/gndf9BFQP0Qd4Gjl/PMkIhX7rfLA3kAXon6s2ZF2mZTHPmPZrZugO
g81LTT+WNGYUUOG6/SY4gqNHGtbnBEj4UZs+4UQgUF12TvkC6qWvOtlQfd7AK6oo
4oTH0QfcSDjMjmKlITkB9dRN3bgS/mJ6oaKbBm4UNlxnQApmzqaVbOyRRWfSQzOU
Kz1lxs2EZDejPhI3sHYx4WtuH0/TpyJvegThu/q9AWVtMwMgjGi23E9bZVFEtbtv
AC1Az0QJlRf3HSbe9/K8TefGd+hJ0v+kNbmzzFUqGSSseMBF33N5APFyueyRi8a/
eRjN9v5K7F8uHBSJ7Abh3ULLFVeuUkTOGduXUM3I6XRwIg+8dxf4mgc9j+M19TE3
EUc4DDZ2iZtxyuZ/3HfUDPhTVFxBiUkPvxbI9CI3NqjZ+AQEui74yN7SZdwuZa50
bDGj6dqL6rKSXSfcJIogChH+JWx4eZAR4jtDiyIFP2kbQXo2Vhbsp9V7R7FIDsAJ
s7xKcUoobuyiwZ2GZQXklzXZ6kmBxf2q+MQtAGS5p4i1wTDJAdhc7uM30YBpfBjB
gAIrlrInDidKdPE4eOjI9b6Lokz/CP2+AaU5KGdbgzMCz9obC9Ybk83wBH6dwR7t
PJeqoZ0obWb1lGroVRUumx6tbddXDfWXpO8TK44vMtSFA4PeiFXjk7SbKhCXRn+o
+AjUEi5qODIXp1deovOtWX7xtrzC0NJfbzqiC6c+5lRXJXvagmbtaL6gjl3AGreF
VVyt/SGQepJ7SAkljbjAVvlZpLFcE4XKDoymvm/0G8gss9g1qch4PJGWOY9qc2tS
9fvGSRE5ZIaflw+7W7NeE1zO7XOExH+HnYOh6OBUMM13VnsEcsA52/7Y/qV4j8pj
PF31+sXZeBEchsi8l/7nub7rHMqkBvfwb7rrao9FkRVaRlwxPpKCIJdNtKOyHtoW
cdBD6Kr7XSZ5xH0WqkLKFKV45aBtpapcBDevFxDMO3h+GHDu4ne0pOq2Ea1cF0HZ
rTlgt9eQJCqNBdR3CiDPv4qMzvazJwk7x4N0gf9SSifsR+gVb91jljMDsqjgazLB
zPrcgVxYGZKclO9wOe12VKjyn7tlaxLdI2kqrhfczl/9YZhOdomm9LwtXFtDlbyd
BQ1rCY/vS0IjINb9OT/fQsQg63kvgEDmYyXFMsIGrmxwGcYzUZ3LeG/K50vaY6P7
IaW2w95Sd+8Q5sK939jc9MOl0VGqAhhyQoEouifbSfaIGbv3bn2eQFWm07LfjVX1
Ou4RawZRCya7LovmdeZc2cz1Wwemqhqc0+OdgnMieakG0LHAfAKo3uCqIGOn2BqS
hns0M9DCkBSV9iAdSsyTolN7FfgHABivtck991/uO+ABlLc3m5N3RE0UEzm/SUHT
5IYgeiSFWu2eTxyhpQiDPr+6LgYGhP+t243kvXdKx0d28cjfwRYv3xQwlyLxzjEQ
8f0g4U84d3ts3LzcvQvmi7uev7V8sPAYukXbJzsDAY17HUj5A3hOriGSCMHQZNM3
wELbFvqNjrd5fKCV3yBgUBgHw1obz2i7F6JNc2zoOSaqsdz0SimmqtTlmWCWneIR
UUtuxtsLz3pYTY3ZJkfPd4ATdp80ZUmNYoaERdNjOxuAqMe+qR5c4yIjMZ1SzBn6
KKX/R8+eqYicafsYD+jra1DOoReDYVr8J7Fhqmoys+iERSJ+bp/v4EubYsej/Vg2
m2Cjw7s4QFg5uKuZW4vI6tb5Pd2sMMuYE6NoQtmyQ6RxU+QXn85bY683gCjQRN8o
4rs5Lpnl8uPKa2FVM6Jd5RTrbKFHn386wUaz3MBtlo/b3ZPhAiY/K6kzMcBESBo0
J3JtnHKwcD4eeEpC6MV2PS4uiZZze5SwHD/Wy3p0uHvgsEp8lAOVyOadOkg7CHxV
f6mkaev5HRXB99o9QxpfJ14bXZ/3ndqMMBDbrLHIbV3IiKe+MYtxHkeyuvcqXIhW
pZUzBbOTEq99tEhnyOcEsBAkp11s7LTC/KzDvvQcc37+UVRmN/f+cFBSwFB7Pxcz
EWQlXIV+2JwICBoD6kqEpyK+I4Q4rU39wJ6DmM6mLgGmibsajvdSwsjoF36ahslA
GxEzVx49jKt4xasWESuK8O104aQtntx93iwdPKIA/bpLbt3DP5doar9eJyxDnSVX
TC82rKrSsXVtBiRpF4vrIideNoq5dx7ttWffQNPIux7uYttbplx1PxKB6XPdVbGR
T9Kp7upUMV55N+VIB/gIgx3Bt7Jo79SY3FQCmdD6/ghhmmsqk1cItp0S48TNSjMF
R0d0TU5WbkUB2myXZj3fcl1kkjHAZ47QZ4EdQf7n+FUxwnIfqjKto0OQ8epT4aMb
telcICKBOiTMtinCrKIyfSb6185XUQs5KsqBQrrfn4ufcOHnYs5dOnEBYDwlKKs6
sx05WJLHeb2jMD6cMHaY0qUhdmD6aN9jPwai42wY0JXTUHnqPYN0YMXmfTNa+aF1
jsWXpMidSBjMN3Omby5nZIh45PNCBwhz1hy8m+aVB95llEoQ2XPa7rpfxhB7tUbB
ZOJmsnlV4NIOuzrmN81aVJP3hHUUcg6Hf357VlUg8qzQdm3xw2JKmQewtlhaJZ7l
GImTfVPKbRYggTyBIrhcHAtN5NS7751u6I/NaLcVQZFQ+omcHeKbWwgcLpuQqEwF
qj7H45e2btnIncW4P3j9aJozfk8jkeGq+HHtzzHdVX2G6oObN+u27BE/4+dDsBmA
ndpNkD7MVlhAyobwdbUT3jL39XuENFBN9zcd+7YgMM05HjvcdZ0dnmYVW+KcW4kj
ykfMSCmJU4xN4isuvoJNDojDXf2wDpiwQNaSQuQL+PaSyT40H1ZPGRiZN2fQsAwi
K+b33M57FocbM5oO7ynmhB7w2l2Bh5vbOCltEzVVF5e3xk0gkAOK0glhZPnOFkBo
2P9M6PxIJK8fJiG8tzlku1fvWqbpyejZNTXzt8dDvNSQs6Y+X/82l+J0MbDsE5Wp
1/pbz/sjIZ+NVrYEM6Ai8Kb24Yd9BC33+eURd0kkCEr0XzWCQjDebGajGfmpbhDp
+/wpUHOFSAOfgosQbEpOC4JaoOTqqntcd9zerYvVa5kTrrMJu4EhdRS4uApi5QKh
nqGS7QzafoihYn4ubi6ja5Gt657tKCmjraZbx8onCcBElQYwuNF3xhEUh3r7AHEt
/Dq7n1Ya66m5hw13TYvlzod2TiO80NB60mpvTusgvwrQFHRDbQ9epwNtAKR8eo+9
zx8lreiPtpDaWv6NlFjjSZTSXz8DtbSZRlmvphg5y/Kg6GTPqis2YXQJAQ8gChDS
q6KHFFuFuSml0bmZNHMAwPFYG0n17j+bvCPuMrPGmDqdOUuUJL/EJSlXS0QwXfrQ
39T+WyxxtHj5eBpEXox36cuSXd53ehQp1w9Ev81kQhY/X6YBIigS6vTZtnj7vfLn
`protect END_PROTECTED
