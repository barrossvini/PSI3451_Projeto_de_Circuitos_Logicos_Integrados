`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qzMq70P5VSmsvElXzRaz0PJ9i2cAzndBrpXjiZVfwj9HaYt8tZ58kfGoT7GFlCei
NI9MLdlUIvdY7dVCHWqkgPYwv2wVDn/1eT5MYlBl+uLJpjGJfh4IPsCLvzvVo9TU
i150FopDOPhYRic5YYCtcNvWdWz8Qby+ZHSDCHjWXXHCP7ChvNbl5Nes5VVZJBXv
LxIFF0iNaKcfBfy/He8pJ8Suuanv0aHs26yxX23D4A7HErqmXgbdf2gkHg4hecnm
5RsmGLU/0gyTYPrD6Rs5xFO1B18CdIe2tACeWp2j19n02X3GDVarglLIJmGYDptA
Wmz19EsMy/AuT2pjyc8823OayKkMjvEfNEi5QdSj9qEKYzC4KnlFXhsfrXJ3qLPt
ZG8cI69WPM4tQUR9Ekk07+tQwEaAfaFy566Y/GA/4I6GXBevZyn1g/f3LeFmyvQi
cvJRHIaPYynI85Gw7YMztwwHmp8Y51gk0TTPg/iclB/e9ZpN7InYKUlmIAqMgK8v
`protect END_PROTECTED
