`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tvfQRSmR3osgFQTDnuAn9v7i4O/7mqntzruSpcsQ3J2YwrYK7zgAlmtye6DPGdUV
lQOujR3YREIGyTBffp9N+9iz/mHsAGHq5R9/9gqsIFvsImkm5WHdQ9g6xXu/kJLb
Cc7kPUYFpo/1iHtzBQuEMqrZCvZ7hahfs15B4nMvHVagEo38oCIiRkFc9tVhnT38
A1P8QCtS0m8FWZaeTUfO28JliPBOPUd1diUG2rnL0lfaNJVB8Ze6J/P13mUYfNmc
GlX4qImPkMSCu6JfViaoYLI8OIkiVsaf49Rjm1iNNreO9igjWhzMrqvF9SoEh5NA
DfySNdViN/Omu+3zJ6VmKg==
`protect END_PROTECTED
