`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9vkzFKu/2fFvJL7CVM3CtNoVc3pufHrsN2eYa/JcPG8U0LR6v+1pY/BUPtvmCFWh
oE/EWQ40FCkh90FQcfrpDCwwmXcufEUiuHLOMxsQtGWlPpB9CKmdLrdLTNPKwIlU
vldq0PHdm6sLn7SLzVJE+9kU2ks8sM7uFtUt2KIetBgOBnl3mv8xjBEVVTdVp/te
RlRH3BSSAN3g54J/6vXBtp11RyyFsmGqXBltEjg0QQZvmfWdBuXCaUmNfy5fu//z
hgu87bd1gnXSfnP4NWgdb4vkq0RTtafp/Qd2/9LeV+m/rFabaRm2JK/CeFOuGKNU
K5+5Yi7g65J1tnmq3XIJfBsr9jjccrvv75PxV+SlpiePYjUJq93jysac+KFSSrzv
2dfZYOojCxSBT3/kIcwlTPRgSswuBZMPcjQYv9pUmYHIZG1llnciCgE48Pp2hf2A
UOR4Cg52YrGDCQoNWDSeECeGA/5/fsckgITLtnZYv/a7dRWaS9PxwQyalHPobErn
JVRnaH9lNesDHJXCCYeyhcx6qc7r//X1jhEpCdX3ZO5oNW3W/f8u+JvFHpUS7FDU
20jibCXVJWqEpzYqOwXgx0UvMRrqo2WhFuY3oZ5aO+OVdZtYcTAlygzmAHokOIQo
AH6EusWyxix5+JFhi0Y9ePgmptzhlNHGUOgmDlv37m3ufwksp00iOPj1B5MmNP9J
7/ThwusP6F05Fd4Li0KXS4uh6HIZw0HFfpH/ExFxfSApQH+QdNvH2JS8GdfiW7Vs
QLuP24JV1Y+t8IWldkql6/x3BuYDnWQKg8zv0Qt3HC6XtvyfKpaBXvvRMgW9DCQS
baku1YFHO1WsI8FW+/7lqS3SUVntU/YhbSfJfSbir+wbdyxmovN7GW9T/vTd2UlR
a86SPdU1PHr4Da27EHesrv2n375goXKS/XriL5+Qs5sdYgrztjgjTAg/vGFu5Us9
bvc8YCBhRJWxuzaA+MNL3RTGNMXGP2pioznRv9hJD9et9e5TRZt6Yd8EEk4iL3Tm
/omrlzvjleW4kmamct0O4f/tsGauVhNQjAe7F4jE70SPE3E0BcMJSFsKxKLrE8SH
CUxPHYoHqssvG8WrU7Bj+/ID2obfEjOXlfSo7zhJy8OAjAndMNQF3MkmtJSBQ6Z5
RSQgF+jO4FVlbxsixlf0OHnbHRl6lOgl2/R4FkIGS2wMmcb3piOt0TKcFWk7N/xE
DcrPCwpwPbbNx6M5VCPBaZqCHOttMxHPK7y8/BtdDfm+pPWxsyCDRKscWQmRsdLb
tT5oORE3swlcwuHoM3RSOk1AIcQzd7W6JQY/R+zsqecCSBGUvSAdCSuF2UblP96a
sL8+DCXyDBZUkCW2UmJ/RM2OqbkeZQi8kwsPKXnYe1E3vWsPAxbpO1BT4/P3GHvy
VFOpp8X8LdYCJ/ME+aj8jJJVzJyTq55r387L1sCk9AfYF8KPk7bvwaeh1j0T2UoU
/yARaxAl+F/hBSeddG2yBXwxMqAsoT6e9M2x1PEmnYg/Sbc7znW/Vp+z7QUID5NE
NG38zXXqe/gpYuU+K5H2yS3u2gEGigYQoTl/NZUlUF7JNV4Hq5VPVzxwjc+5CDuD
7+FGL5OnYX8CRzcVVD2UhDHBnnm7ufK01z+tnbG23ROG+6bjyQWFkvakBH1ocUN9
EKfmM7iK07q1SFDsnmXVArFTmaCK2sJuUVT4R7t/zYf1Vx6QYp2uq0TXV4lEpgMl
zvlozUDXRNRGixtS+8yCLEFHy4/O7OSqJrIfqxBavG8/uod7s/nlHVvi38m9Sjri
+NRHEp61bR6m3YmapySWL8bMphPmk4vueObptYqM3Ruk1Hf/3hAwxiepjFM/W3lC
KTOmCbk/KWlUAcl38meJzxCcENoYz1V6Ol57GffGFzJYoqfBQczHvFrn12uhO4nq
jeru/Qv938CObapCnpqbf0fNqnIFmF8tiMhn8Yo/6ydMdkZ/ISYt4TlYlBXHmkWZ
qYrHjO+YscgHA4nCVIuHvMqtR8snXQlkUR7av+VkBTXf198ZyYTGsAFrgG7G0Yma
D5JTeqdVkHhjVoIUB/SvpoYXlWcs1v7zqei4Biw27yCI7XFByJRJB+RmH77x/sy+
VI2wEwtTCWQ6arIlr09TvhpliuG9qutm0srdFrcndl2F55qqUspTURkqYRPqDXvU
OdZXVYhOs9XJHzSXrR//xyTbdG2xz8kweocv5gIl2jc3HlB4P3VWgGpQGjq5GaGg
8GPzRFJO3cN5Uez1AjpMRkdcYLL+b4e6QyD0tscCLMK5AimOsW7vLj3Z9eeDDuTh
me2gONpkJuwkyuKwa9VoqVPA5GtwXsLRO/34A2t8ozrIHSe3KsTA07p7yCBTsbzN
VRiIJyDYAd0Qk/aWh+gjmLtuTWrs3WaLPo7D9XQ1ao5J8QIB9NpPnfrSolsG+gPX
mEhtIt3xzlXS+4dnhEx0480nbEQyVKxxLqB4WiNDdTVRer6n0QbPHLU9cPikIikj
TDaw3REBOIVr6hbBXY/pKn2EczzqgSSs0tkCoNuXUTkRqe80UWkCKEe/CIfnrvm5
yUucTrMkhIkBX68bb5UKFD9XR/72ZU8IQyREPlt1pexD3tH/lNZdlllpq8BY/hMC
xa1UIsFaeQyBsgJXNdWJ219GQ5d9VRvePOF/O9HI236s4lcvbjHYxmAuSE9/SlCk
FI9Xm1IQX3lTJYyWyxyoQBl9xxAz2cqmK+NUbYeksNqRQnAwOey/gXQH0Re5L28h
SR55EQKodUTzPpjvRGJWpD0B1d/lLIBSQgpgVfFqDBISelcNWhWQyPrl5KjgptSk
hQgURl7WHIgP4d0rucYBw0XTBykjwmm4k6o9DqJEDgTZLgowLeSQYO3N7c+By2ks
fR7XqqhvbiQYnDPf5WdGJmnKWmjYaxTWnmYwg7W8x8tySCdMmROpUikIiFeDiTlp
R54dsK9Szwc8KD8xybp0gLRNZyKx7D6uLN9tUYDJAaUwd7DENnjkdojDbSP/Z5yk
N2OunNqKxhXyuiIVgOe0SOpkGqFb51b2R4oNg8KyeiWjhNq1Lr1AYgGnu31WiM+E
kJi11TLNzkED4v9n2qqj7cQG5ukHpGvrZyDOFOFDrrVNcwQFrRYO4ErpaJ9MM88z
qeNgZbOpnUtvQ3GqQ3xQA2wZy60V6OIbI9OY6OCi5NWYAK5gi3x33F+pmuh30B8P
ewM3hoRWGVw+N1nVfH6D+tD+WtxUQA86qe41krhPJlHHkUzAz/qsZkeb4c8QUgoB
1PEr6ZZVpVejoFWiakluikfqS8Yma/g3Xbmm3zPW7J5XRjBqTt74uOMNCjO7B+6u
K6bTPnHQapoGSXT/9U+lgJAULFWYEMhyOKCuR9aT/Kkz2tM5dGw3Z8o6C0D9JRDK
bj2BkSxiMQUXJmNa8brDi+ryI5/xabDtyzLW4/UgtVaZhzVa8NwiaUFfpcSdCjjx
9bW4SpLrm0fKdLNG2nQ/bu4yUvg2oomQ+mq8AKAl6Bo5jivSBJtspWm9UeYXazhS
fVmyfyJ6mYVxCYAUYyc6dwGpEB3gXctL6DWIq/WUKJePYf0dMqChYUmQCtnBqYEE
mG4EKIkC/lFtDSovRHBwzyLPeJ18yY61rssR8YOedzmPkdkjrqsgcUQEKsXZU9Nj
KykwJ4tfSxheIpkD5uzofWtmYpe39y5WmEhdjMUoJmkK4+n6szeK1QMPm3mQLUgO
AeHEuRJotvhiQkXnlCXmB2/w1DqUNRbvHOROkddgFkjQKeAYysfHc4nd/HN1k0Hi
/B0S3cDDZeenTbtt5lP+3naP5xZx+wtNTnMXs0ws94a6Ky0bj4oJ8vBqwPqEP6Nt
XvZXxf+24vNmn8fLsyISBWzn2RI80Ymehd4SXiWUyVD1vQhsCdEgODWdiNrqsnV3
w32NDl00Y4pWSF1ViMT9Tpf8SzgUuaRtti62T23fye1ZDlRLGlyyLEh5nC0VCKvx
Tr1zM53UxaX5fYHEJAiLBLZy8SqK+9UlRgu0aaDibv6GbpXEv5L9DWtG3n0qZORq
N6tbsRoZ4k6FRBtQVNG5ziVHHnbNm5Lsvwr4RmjgoajL1ww63+duM1O/ofUkkPoK
UNW6+GMlroLz6Tj/s6ioId3DhHqVdA/99/DL3cum/ZKuR9nyNZlej91ijwXXG81J
UpK93ZeunpNo08kOTedZFmP5vkWk4FUR5yZhMx5uUDxf9Zon+ddhhdP/cRkpydjF
MQEik8YR7rgMrbxM7tN1fx20oTchJ2UThoNg59OwZDJY2lgr4PxPR4NDKWQirkK+
XDXmnAMxaVAO3AItUjl+F0xuYA66citbfEHkoFZM0dWzEEevg9Ch3zo4OlC7XseF
kjn0wVebMC3/6dCpbYzhAfOcBWLNIS0QdN5JOeHoNQrG9h52hkH4xC7ZIeLRUy9S
EQWI3gZQdJpOtpWUmS2JVc9i/se6iJquGEkMXTeRCvFXWPGr5SVxZWIKFZvVLGLd
nX7jbvH2fJzr7Gf7czLhKB6ItW+KcdSxCggrdGjZqUaHprtgIqE8nZ/beF7FrMcq
RJYIiNNTUecUNPeRRv/kJRZIromTfVjYNvjGYxSg/TmHUXLFyGj+YMuBYiBbOt3J
uvlSsvpvMKqwd7QNSS/ccDrvXCC8xiiodzS6E1Aq3bGbd5lcQhGPMJ4uzgPlU2jz
5fdb0knjzs6x4romJwjbYcb6zBT3KgAGhGaML7W1LozUZQoSSx2kbgHf1P2PYmHB
qq36M/GdJ9sxVu7vVfX/Ovtyhf9r0GQFMy6F5H7sPiihlR2rFyWa4Dbfmali+zIY
59rvLi4TOlgNJOVVNi/NHtNkomQHZiMZvIxwQlO+8u3TVWo3OUkJ2B50SQ+3G06C
lweTM51mdsPiw1dxLvTOkmXVhEE5D/drlL5X0k+Yws+ZZAMhKh8UHIhkEbz459c8
w7Q7b2DvVMMJMaxDRyOp+C4OmTt04RNGsBwHVGK3iyrFIOUjP1T8AnJ3zDYiu7kH
DpCrzPpLvivLY5Puh5SmrzsffLN95B6tzIFjWi4KQDHPv2PVLz9qRkWAzrv6Vyy+
u6fvn/gEYSejSBoCuR4I8Hdb5fCMOarVNYlwTAPBq1vGARP/bBzboPqipRWf3v6T
3z/mDNvBAioy+JvQZYkeFR1gS4o3Wprhp9OOxW2a8na72OpfJ0xEi3/4ABSavgfx
Qyymv/jcMmErKMmtMD6flM8d6PlWWjdDs/FW5+hrjEnfDsJYqjAnfAtDNrzZvA/j
M5O0xs1/LEgvDDT1BtxFD6k4hLz6E3kRQ4wfC6EoFXOEvOEm4Eu0N4nkp34f8pJx
1mEuppuP3KlVQB63jah/r3Ye4SbzKg+Ls9suARpRASoyJa/g3g0sFP0MIZN27X7X
J+GbKl7VC8K4jfU/0oKj9t55idc4wkwJp3PWcvucwm+KwPRcNvZTOBTFQIvYWjH2
iUbnx2qHpT4qENbyNn8g8EIUFNwtSAAQZJJcXixS5TX4AZTW5r48BdKekJrclIZs
2eivz1LvKgN1hQzaRabIqvwXiomqf1mgq8j3OdsgL4nij+z96Y5kPilRT4JuUDaH
Erhs1Hscjws/PPv5+PaMJws/ZaTF02zWRMZPTiG5LGTLdCuzFu1dQ0l7jTJp40jx
JqD8TwJWUJz6okzbdJXj420usVbEaDbNTV8GelvLWEsjKRwcJOVoBfsTfVzmmRXh
EvifOQEEniUBG8hZPfQXOO0ynr9YSb+ymIh+FxI4BwqkxQG+P8tlDkbK7OpLz0ot
14xIa6XUwXAwKwiAW+mt75ebIvRXXXbRO0DI4PweVD0fsC8aeIR+m356ER9d93Do
KnFqTrOpiYh4CDC5SyEYdYoz4qY5lGPxbfGxeHbj+YRQ1221t+l1H4AiCLWGpJ1W
vdppIZUJVN/AeZTfgYUZUzUVLLbmXyTXrWRrbQpmhvJYM7FSH1AfEnxlkrzAJeR/
XpoHOy2XmbYn1A0OYdGqAKZG4WkXpxpa9j2mEZPWVeiIn2Lwy4LsNhJV/dWXfk6+
0umSrD1V7w0dBfXqxojV1gpFyKOdithO8wS1tzQ3C9Hew21g2NwyLl0dbmq1lMrQ
XnRYQbPSFmKGO9bSL5AXNbdr6ZkLeJaDsn/9DC1NjWTF4G94JVwdlxYHbCu7nKVf
mh3fy3A7UifUKBdKaK3lY5jvwACTfZWO42eLbsktRok7KhddluZuot0AFELcg9qH
1NXK4/sFwbEqfA5AYwVMf/oKdLmyHD44QFQH/WnZBP2s4r3D7oc9r2pjLS0iEDxw
PV9SGyq6TVVOkcU7jzEycpz/A2558Ll2dBeoJgRZ2eKRjBiqsKSn+0zsJZRVg09H
5OYNHNQQ8la/nBEH/6qIR4UuUqhVoWLBtTCz88i5Nmp913tFY/tSPiboMbRAuRtY
mGwsCbmkkbZWh709lAjBK9d7D92zv9aALoh9qf9WI/EbVslE+PE0gqiOgbJp4Kly
iTxTI7aUSXqDDtLlQCix2qdhjbQG8VcbepjcMheyG2MYg/vB6kEFXnjihlSNcg40
jZGHEuuuxH6cV2IkXlbjr08/O65ZR6zRyCF43dwSUs8THfwRF4XjC6KlUkOJ8Get
sXq7vwur0/VA88XdrUi8f+WVG0EoQQUvia5td0Oczk0q/orHbNQkJRIZVTvSzNTw
9AboXCZgtgTz1GcWS7EdBvexZS2/qsRc8oZvmc/qkKDLsgfUVXldlcUNiMRhHsGd
fEi1s7bofKEm+BATmN9ulUGaNCtWOhOslyWOouVUCEsrJkZMplpAbV7HfbN0rNFO
hQDEqtkF7LbQHGqp3OkNqJZMtr3JpRS6yrjyHrI1TGHCkeuFCLc/bu7N75cUc9jC
eoOTmhUqdSqlfB5kKMvgHyZ8ouASAyn7TCdz7rvWMoX9ySHcSznyZJlMWm9MdUS/
26KrdY73XZCGpT3Re4UM9L6JvXBCOQuXMtwkLVV99MN+JYMEHoc1IWdDCrywHuUy
eW9cLQhRWWWkLX63HBy5PVndnI89x7fnf7/elU7VUX8ftG5WHtQu4ILzIufsFT+N
yU3VuKnCP6PyhkcXe2s45sCO2u8OHRmBscDRQMWFjia7h92jiOw9m0NXhA8QnBwG
vqymZtM/bQwU0Pxyg1XKPgTdogiQ1l1QKO0zz0mQCTdXxqdJEQURLUcAt2mEiARD
fRHWTMftrK4Uqf0Ia14DNVh2XzSWxYVttg14Gwi/stwTUzQZakh7TT0AFLa5aFrz
nLjE1GqTMokUUP9bk2SyKpGmzYSi1QVX3/d2/IzQOu2JfdMUoPKLGTPPiD0ShYBN
JqRxm2KJ4srX2T/wmInekNNLHehdFqqo+i8abfHB5fB/4qEpkgH9zAyD4Q+GTkJC
K4OnXD/Lr5rKsQm48ArIaIZ4ZGIxk4+qmLrS01Eyupc2pfN6ys6UqMAKfz3OSH2F
1GVbaUYQMKxiVrcgIR6bDsaCZlkGHjpdUdzW/pkSRie3Jw/QbfvnRx3KMhOy0TXc
6f3RdoUTsGyF9XlaVtaIE0uGd9BF6mUCdf60MOkaG9Afe/ouqturAf60WSTrgv+u
ArFBdZGocmnlATcvdD2XkGTWTuTMAQsg2Pm4d6Gzl1k7C4uKzGbiXQ/8TOSdtwOu
CNpcCtDPUHN/Gxb0RARAaSNKVZfLQvM8QwZOuwddyKpzpo3L9hYEq35A+P1a+9wA
PurF6wlEvV/jcw6GC59klJrLOLohH17FAh983NXClanZdoWdox+R5gS5WiOVHFPC
I2u0NxVWSLpcju/1xnDBwf2exoNbeMUjKTBQnHk6O0c9rjfN6mq1oMxNngvThKHT
1qz4WtqdzonGjTjli7zgQ1/Nfjl69LXubWKNPNd4vCfQMc+A4NgqybZ6JTlBgkCv
KbWMnHTvD7aCWFM4BN/fmgkHKmsI+mzxTPckCqfE94VKUiHazyuRrIytttu050x7
XXvd8KfvVb4vGa5cBqmLdIOqTmjsSXsBB5vEHbTrTguzkyHKcjWIY3Staz1yaF9l
PaKATBEwufB9K3Hp6L2vH5jio4Ff9RNjwEkxTJUxf73bEDj4y70DttKu+Ro14N1D
VCug0jYLT/ANkkhJtEamXFDB2O7Vjg1LhCYb6MJjgLjD2XI4joZCHon548oR9z5w
ploXvBgO3dUNNoczlv6QclD09Dl64SHoryf0sHT8hcWg0ONGLjSfps2DkTxxw5Ol
M9i1Qhy+yHQ+b5Bmsln02b4GuTtqBkt/1PfNUhxHetEBUOojW/f4TFtw7fq0mtmt
p/DcQWnT90WFz7lLKzVd8WKimuKnBYNKPwJkNKqfWnAfOoSBHDgT0M4TZ7KwY1lw
EbvVGA1zjNo0+1yjwIensIORL2OsG/FT9D8nazjMmGqDya7I4m2uVgTqJOXCFJbO
i807uWibasARzwtkY3tCjMxKt16BbcBGvJ2zWRnxSX+C0E43QePgqlMV3sosJNSp
ETRmw84Cj05p4Wm0GxFLUZi8pG+69xgy/D0oh89UdiI+VH0OHqEl6wlylIi/KRdg
hXpYoOv+V1+RKj1NZirmMs+np+qIYuNIL4kCuMPuD/fFBCZ5/n6sx4tpm0iHdWWV
hT0ETHRSW1mVjsEWeeumGR5S/26PB5aR4WJUsIgk2YMNIIAjbGoayRWx4oowZzQu
kimC2/sWNDUAJBpjPhDeowWMtPRhwHjpMhhhx+q5N8ub85fy6/9SOH8lceV473RJ
IzWfbrGCI70to8wZHXP7WDOLiGKZMBTGPedx2eFTUIgpjzqhWcGuQa98bcY3Dvcl
K5kI/0Jmn6IdHCGNvwQUJzxDtSZu2kpfgULSe/UP0+0uCwcOfQ1YlNfOs4Z1ekK/
o5APk5bdU/wSEynDeunTOpauWoYDwdgPdgphoXV0RNdN+9VvtytnV4TQXc6tvhVs
NPd/E0UBivlclSj46DXSqtDj2bqEBTc96aM54FmaL7KcfyTxY5zamKJwNc1B21bK
jbGNNvwtKOXovzPlMRsKSdkRKfHn6qQYJfsp77cKHb9vi5203Ao5V7XLiBsmXNTC
8kTUM0CMKZs3rq5Guwegw2wmWHQYzyybqS9knDSe1yNR56tor29rlcShBKC5UAtc
yO/B1MUHUXH/Y0v+nVu/T7M8DK6dz1ZoVUOX5OCKlsnCwy23KYMgigBX3PTCcuhi
0gfXRF87tiiq5HQtFStlfO/kC8HTQLPxMReIyFQwiG9stY8YR12D+qsmcria30o1
XLoMUKp8n7JPZF8ooJsw7HOUVirAtnrvjae4Pb7E2maYFV970OGwF729IDVPAAjo
Chqikip8LZmaHEs9DgNpqmpCgqFL0iOEcU/9XIBi4vxva/eCVSwiLTQzNWAiPEWb
ujRqeoAOU3U/M6TfJs7Nyr3ko+/N33U4fbaPaDvXryyRNqNzSVtjHMmXn4utiSqD
8jHo56zMDPOTHnYGm7aNqOc14LaD73DGKDf3vSIJsR8WkRQ7xJe7eYqd07WqB26O
/MKWsiX1WwAc9P7sD0t3h442D+aTWBUyCerD0NgbqwmYKj2gknkKa16h2DATtRHh
qaQQT2k+nCqEMwz4/MGlAnoBw5kfcZ7VKTpQDfMyDTv9uaD5x6twKCSX23dd5feY
9MTlvtf33SuWKmO3Y21d3oidaXTqQyLMcKKrnst8VRbu1iYIuYAS/iq67RccgY+H
9TT7lwerRHEWo7/bmCGpV8rP/Er/no88vRqsYOdMPU5c03AYJRAzdB2eyE5tKuj5
TJESA/WUrt7PXOye/33w1D6fI3gtUz4B/wwYc7kjwqWpRNV72aBooTxgVh/P/wDm
h/w9RrNEd5nieEYfHfEPn1hd5As4hjeA9mgTgK8zl/19WG02zHPYn70bmn4vyARc
mQRug4WpiFjepI6EheLT1FsqIE7UkUbYjE2UopCoB01MfneHG90g+1xvT98clImk
R7CtX99cxCQGcE9C8xM+mhOp9AHH1ZqwvxO2bH8c/LCbOHMUzlLW6jT2jId7wbkU
l73Qrodix9XwXzLsOyXn9T7YmJMemGHagVd1+3Ueu5rJCyzDyqCQAXK1hs1TkFDv
cNJOLnNquCrgu0jXOvk3Xl+m01tU2mrP92uDgTCmLG0SnO049uoLbaAqShkNFLT1
G0eMfY4foUxB61rxRq5V2REML+rO7gP5RJKvfdXuqSByrodayw9RbsHHNxV2ALhe
aqRVduz19tbvjpGo4uU30s1um3I9mIJYTra5ywxstnDScXClsmPUB/uSaHzhyn4F
eHNCRtB4MUSgPNqFaVX1LYnTYiOqYWGVngAkBM4xQkGG2hZSJXYciKJqOnolYM87
2a/0S0UND4W05EPxRRJO2NiNhSc2EFFKBrmxVv5/Zyd6tgc/29dPniHff03FeERR
boWYgxSf96phbDEJKLvxrw9yOT3sKMuz9z/zlApQ8i+R9uO7fIyCy1hvLj/DpWCi
RGx5hxxm84P9VaMPYnnEJ5uY8ZXdXICQ2pfIuJWdsXPl64TJRAUgTAe+WtgP+Igu
t/KO3Li/nwNNpHEB/Ad2hHTPRKBMDYxZj/LHyLadAavGk98VjO0esUwlMinUylFH
keomUl9eYHCRF6swfFTTGlw8ktwov6b5a9y/rgRLOUceVGz8/q3fEzqEU5ChInHq
Cq9yJbTcwWlY/6eZi1C2ry+PiL5GzyiAHBkYIxByD6Yj/WNxJaLktI+gXH0q65xl
wSS2OQBpn02YtIA4FtU1ePYbDaVqa96ej4NQM5eyuej+ekiGLKBiJx7lwFd9Xy9a
QqFs3/nUyJardnDTilieYaOZhXHF9YT52YjwyVKjCfu5JYhj+DXvn3abePOfgNmN
fkzkPrEinNoRRUPAWUBvpUzH9c+gdgxpcKbxClU5UnNLoTMxfBU0uPv3oop21zZl
XjEa4+/3yvhUwTFwd0wzZV4zZ2bmK9ReXGHh2Gc8HVLqBsAtVHrTq76bGwHYQ1Fq
5fAbF82qJDIGCWIdjDMt+xeFAoeRq6cLmitPz0OUb/uxpaDW0xw9UIiAlV7nugAo
v1cVF9QJj/NR5Trn/8C+wExFZSrIdRNSIT1tvyqaSeuqPUvQWCtJstpKcxTIwduw
lnHI6qwkqhu7ujuOJjdKXJ/Majrr+OHB8YF2McpC2tDYxaA528/j4Re4+oSSSOHs
mgfi8Speb0pvEaWxfGtaQ4YXcwoC5TIHqyOhnHsEbSL3JPn0oI/OeaH+khB5Oo8R
fHFclxh2swEwa35qeWEKyeybZvGWjY1WoU2QumZqa3knv/9CUR59iymG6Mqqe+L0
jiWUriFu2asPAMmzcPWqXiD/GSwd2WdK2Z9IbsGlEijOFgINm7ybswWQ2EiD5/YQ
SR0iy8PurlQRp65rdi/6xZBrU7+I8vrmhWrTj747Nj9umN7AylWCHKrPYiNzlIqk
UkLFi97SMMFnxPPqkY7SbO6CvpA6GuFuLvClIwHGL5NISWrZwpQj+wmvhDAIl15/
jKCln6UcmlzomG9cz8M1QPSQjwAz9vbiH3thPRudMBQP6+qwhRY1cFXzyTr0YS6a
ZOjurrPWFB9eriWUIekuHg46j27JB8T4cqhu42+wAFfDsKZlAs/gefv9dArLK9dS
Po/RSDrQWol1Lp87TvX+R/NWlKEKfQXyb7wPpJ/Ollo2wB776KtAn/VIWV2dsL/7
5tc4siI6KcjKoTn8TmDU/wbALgOisdOaboG3o+9G1+SfffbUUrnW5uMhgWsa92pR
hWtbsnf+OJX2T++F1UXzAyD9R1+OfctVfiA114cCS1shQ7WQGanfG/bfDYARfmlq
vlgH1IHqR0v5flu0udOa9ETNBxAsSUX1gZVmNMaHaxcCwsYiuf7XswHmPmEU5vbQ
LeV0yrx+4tfukrAwtwea+0NTgz0dI67BUjxZqqnqSIfImPPdctxCY0dPxnmAWrY0
H7CU0lks2r8N8U/Qm+NGAo9JSe1cqlWaZYJGbKoTIF/8iorVzgmpFzKSzLumHCjB
9TEnj3QpE5qkGDZaGTHsccRco7p1x3VrpqI1N8+ZkHuQ0OZB6B0FzYvJkV7mMm/6
8l0CASN5pcxpy9r9ntLlw7zHeeRT/qNlon9GDEawUA8aWN5f8UeL9t0T4nEhzAy5
HUqhEPDiYddUscB9r+EI1jJbBIN/8iWAVMX8MzS0EIFNFg2SfUh5XpNjNUAcD8W1
eDvQzB4rOBmpI/a3P9GoFYUn9ZoffU96eBE5kl039hSILSz8IOyLCtSXHyNHBtTr
nRq9ml8uQH0fwxxX8hTDReGcrJOFx1qvfVvgiFaKhfwrQGNPpHRaP0IhKUJg7/LN
vsj3MgppOpnR/nzTvK7jCSGCQc3JX5Y48euHVmCw9yt5iwY8rxtdLXixxBMOGcZW
LlLW3Fu65RPqT3gvMD+ePvR0XTOH3Wbe20rbEdh7acWpqkedeDqMGrrSf19WLZfe
xLe8XYlOIQZdqrCZHcW3zdYrTPu+ecaG6Xu+E6AMPm4kxNgv1n0pjRhNaxLfF/DK
At7a1L/eRv7P4nXS38feW0QpbLPGxCCKPiBchHFboWpJYIqgNvar8UVhTSvCvpvS
J97h15zA6Lx0QA4Pkfgbs49DOOxPBAyWFYbaa7ysrTisIxTcpZ9vEt3nJmLcYaW/
ZUqhba4FUCO1y4b95viNbmGBCVOo97NEmEH80u0WKlyB7aXgaIf9Jgg6ASHkczo5
UQaRZNUFUXgFmSLRQkYNsyDERL39WvFK1eqmRP/mMjHh+uHLuUUGneATbiVitSzs
vNkgc+6Zb74/t4YmjhTpCX3Ul2otpn9/FaLp8ilKxWcmke0e2k0yxX8xobDwddmd
/Hxt+vmvY1rgvJJiPMXliL7y9ygtpNl2ThfnJ7oJl0MaYIOutYqPmk+amf7VVUEm
RrY5nOtd/QjQ/2cw3NIO3H8ReULRFNm3WqgBPVFmRh92NOkmOKVBWPt/v0eYmjC0
Y27FoEb6+HlqerGl1NIHq3M7CXH0QIoyN3HwT6RzM5SykGs/HN3lF494Syn99/gA
b1cYkODofoyp+ghortpcJ7RkxFljVMBsfvwQjUum+WflwCiccLkyYtlk7tldumTu
5e0Xt8bp+cI2yBwBCuiQi8dMcLAvYP5pQSoMzsLORcqHICT9C2vXmtUQpY47Up+7
P8VMeRP2VCm64agaXYLCRC9SBAges2JW1g1GSgxByjFidjNDjCL38a+GE0rIYavJ
y5gvlbeXGyuHz61u9SPnQZwv+DQ66SBUNaw+cD/08Qm8nmJ/6R71diqFWpsiCnO/
1ky0/6oHfzNVfIj7hH3EafMiJfWFfWDqq4++w/1lu6iTo3tKG9Q2TQ8ojHu3sWZ9
vAOMPZQbZ2totFxjL+Isb84vXsbbX2MZvmcUYp/5yLBAFq95qbYJ9xN1yn+o823S
xYY2nWPzsJVDemKAtLhQp3RBbHrw8Zkn8nMDkUVdY5AjMuf/x3OAQi8UdaK2B1Ps
fh5Vv9R9rEk2om/zHmbDlSyG4zhWgjlSRF9sMLNiIi4iuPD+ILuBGFnnVf8p+T44
Gu0yduRDkcaWkqOQGnEsxcWM1b2pNoIYs0QbbEbYO+UeV0nljCuJ9jz+VgZ56wd8
7xRaY770AIY5OlWRK86eY9TBIq9GhkGJTPVUDcsw1xoHPEXlEOtgIAi9u6NBRh6O
wySTKl6rckWTnkBollOwF7EJoHE/Gn6nYxhVWfMfWY0yWPleaoRb3stx74tzc9Pf
5dv1PFzH9RyiedNk6sAQhIwHrHVlsaLNDkUxv6cEzU8elQwkrNl3ug210/5F0VJH
bLOOb0tielTEkrglx4rbBZixAGMmskYrrBc6cHI3zdnURuDU5MXzym5oH25wa1qv
kC4iZLGi3jxn+S9B3G3naY9oCpu6tYYRO+SX0tBLIV09USmOnbQ5L1W6XIzYtM5U
ze/fwDz2p9tvH138DN9qwxO70RZzYbVVIojlst3Egva21dCcT1EmPgwo1TT76uu5
dggIvGgHUEHv5pX6NY5jGI0wvH4gNUSr0JTMLYE+AOu0ykd4FtCw5vB26q8Wu0eN
06vuPxzeH4OxJ5pw5YWH9e/MzKsfNMSSmpkjyfBA8DXw830fkjy5CwYCWa+f/Pvf
RvX11SIVVJ2cvzoQN4dayEXmZAGdexD5OQlcV4ZZdwJ+2ngxZ5Kfu+fpdzYCXOsU
vIH3c3jdqbFjJdIoFNqm2jP6+9GjCnTHoxZeA7GtQPa4O+4iRlLyeaoGWaeAQMz8
thGT86AjvwOYS+Ja+j1pQo4EVhPcVFnRgzWQY92/fM2s0E3nXDebMHAmlL5BNEdL
iZPiitZ+tBi3FB4mAJd7XXnczOUsrGWoBUjDvZP4B5PcNNngu6u5Qnw5cnpPEZpD
fE71ZX0xAbIET6NO3nmSpI4QKG58IUSwZI8xz0F9P97q3LLLS1gK16A74H91efHo
SIBL8iAFNbrAWlattpm0tq0pqt4qqzTeMGHmV2ktAmye2F91cTlC6U1NlQG7Ak94
+Y0GcUj4IKCHU9YBS68++/DaHC8rfdPZN27Z5JWPyIroHzGGG4ikSztA5Jcdf/Xl
3iRYCxSqRIUrXtmL+OlQSK7uHaNMwNSLObxbdJ7FnVaVbgVjXySTAu5praukb7Rs
E9qcbBQeBoUEBVZN4xqYWTh7ZoAxlSUO+IkeClriiApScZsqIQ8rA0ru9Qi/JaA6
6V3sjHUFo7vOQ9sF9uLfo+emLEhL6xFpZ6RLYZwZqc7yWSzD67NdjSKKrIQmQYud
GyJ3FmalY4Y/WIlhHUoBf1XXo6UkRPCQ8q7vpvsGVHuUcypZfa6ZAqYKA6vttNrV
9GNZdqlfK2Vc9qIn3warLjTosh06lSyCMD7G4M6HzBTMdC+LF6pON6NSbzEbUQPC
XrdlScfKm/s0fiQ0+2AgWzxg+8DmllaU+AXgJo6YIaC71E2WwH7Gmbl5VGUMDWdU
mE60anj6rkF3QNYCbbnfcHcjrgbgAhX/8Fl4VkHHZ/CmYkqSrGdg4FSOaOP1FCvo
kgs+R9ifRy48qOX6AY4ZO2tx5UU54NQPL09i7fE1veI11qMXiSuNsp/ZuBscj27q
WYJZXDTdcfQnbYW1uC8Cen67iFrqcU7UahRd7fvA4ZMSeYYZsDd5V4469Fq7bGXM
UZHnaNDk2DdOSBuq0oTSX+xyIvz+U+rvQ53ySJul/YYn1H3CQnwlnsR+Jxoei6FS
hu3eFjKZw8/lxPC9HSpyGjBhOt38pxm2ObFeRoCD7RQ5YSghNdE7m9+rjhmgILOo
BPrqaisPeNEaEgjJdgWKWZtA4/M3EDmLgt/vloq6Q66wca0YomGGfEtbp64fAHeo
f78t0I33doT6sCNQ27RunCzYXZQqwSF9eveii2/z+h7Z/xLcDebAUkKazqkGxXDd
2GNQEkufZFukyel8CBgOWdjZdSyKVYm2Aqj87WIpEsSs+sLgqz644rIZbMuOK0FC
loTnBg3JMJo1o6odgENoxI0ipYqJt0RW8iWFDsJIv17CnTfCp1kXmESSEb6l4Goh
fHMzudq+cP0PZYsvTekb/+zD+puScxrVGRvVMHKKLIfD7TexFNCIf1micfxR11TC
TxcGp0qh8Hc2gzhn5VEi9iDy/sDFK+P+fE17lyQ2qzj2ywqeWXpBj//HzCWZ0rBD
6Rs7Aoi7MagYmgXKqGqWyl+sIyE4Haa5npoyedJ6+/pLqCRzyYfO5znIut6XvPSs
iwE8fJwlUCb6/DILYw3clhB5lkJp75m9JN7fhj0oLwu1yUX5BB8GjHSd58VEwmUv
DtPD2uLOREIAci7ANN07aEB8ugElRrJJXnIv+a+o8g2yaqNQPupRzEGNEYHIuT9s
2V80CbYZ99ItNWFPVo1q+JCdGanz72ZlsTaLvf5e2T65HdEDpkZ2/dOoVl5+WsVd
yj26OxSlcS2NAFrVFUO4Tn/ch5rGpmyAARFbZ4dAofv8CUCT+8T2Z+aYL3PWltO6
P0zPmJo3+LVGf/3c1QyHFMt8ZVDiNlsqfReyQ3hVjLS6008YQJfWz/ABpS3D8TiO
di3SXldLOD+DQrh9Eg8+S3/Q39/TzUJJyAoTWlrMQALDeCjnRmf/jqUXReXsFtlZ
3ACfqjtpViiFOalA/boYZNjbWy7WJSEyebFpLDrQ6Lke73u6Tnm1yAyW3YVbHF0g
yWwR+/EfLD855J7PwVtNKPaWFAB1W+br5Rz1S1eXafWfSKSFX0tHcuYCtNiXBtoF
5UxzMjP4M80JTomcMgY+qZK7UydQ58BOgjoOScx4s29ZjC+0FuqwzxbUAOuHVa6j
0miYfC+kEYP6nBVZPoeDytHwQLzXQ+o0NjUfuWMpUtwLTJv9OAYzVzEPv31Z/heZ
q8JD2y6Bd3YETrTQ6IiwRDKZBYgIaf1+MNHtSHkN3FiZxdTjLfDEol5xC/dbJVP4
WkhxpPduXgIxYM8tUUPQU0UhNincnOK3S/3I2LUQvIqGtTQa1ny8WK+Iu+Ah6tb1
llbqNa+Rp6p2VEPHsh7Bko1pYn1ECn3djO4W7YG1c7RdbihvUGsdD1D5oR6TN66i
4X91qQpeRqKF4Mewt5wQj6IATuSSt85HNrHIN1maemM3eWABTOxj8iLcwy3fmDKh
N/UMYbqiP0MaIimVhsFN9d7V1m6tyAzg00CvZe3eYGbALAkkdpK4i71qYRW0+bpz
InkvM2sMm3H+Ay0ueiFzsbJNwFdBd27oN9r3cW3mDfPLeny2CFABdvuxoxw+4LFG
JBwlIqp+mDr1N05fkOHMCR2SQA+DKOnOZU6iIYpgjla8flRno28cE86kJaJKJkuo
6VvlHQrFsJAGTliYQs/lhUhiGvBkqgEHrW6P4609TQqIJEXk9Rud5wtuHNtPfkZu
D79qpD1qR2dh/PfxvzQ7Ig+dN/l4D36hju4evhlPiV60+02Pjt4ph6zdCci28ZGF
7EGjxCy2AcN3ZC6Vtzbu7ZAnOwncjFiAySnpEBv7HC1J+yfmzQPQuNAkkKD2EVJ8
+RXzzxI23zf9wLhvJ+EQownWj6MC848qD5y+csdbkaJfcTM74YgP7LoFgtS1Focv
pub9dVX3eXOiUQKVsXPillFqeb1mzn+wUIIEQ+8hRmmmPi0/h6CW0eDXN2Uf1ghZ
WZiSJAUEkQmsdh+Vp8qFDOcBlYTsGsUONfwyyWR6HM8ikOtWx5Ci2aPDJRSLiP6W
JJ2CkzJlJspCZECJx6apPr7ZQdZ06uSrrflU9Cj2O3lwXsrSHUuwRnc+azYijk64
EKS1rrF75dBt1zxs8aUDjsqO08bDjdDaBiyDEZBIruB+4KsL+FDj8allgel1ulnp
q8dWsgogTSBv6bfrLdQb3qZ0paAujCNgMURuKsGPi7DnmamyPa9j8V2Yw88O3WZO
g0DyHgX4Wpw2J5e8rmg5HSsGzjJm82+UmCQ2Ye8cOOTdVyrZmqJX+CWvWLPONuTX
tn/QucmnPXvldu9PGnhwWEiPgnEOdT791aK2vXOEDigFiacZaiHJbx0eLRUmI40/
hTKEuId8kmtXg+YQQDC6alPk5QeymcnSquUAZa/vXmvrtVQMns+pAJST9qp7OILI
M3GPC3Q2EdlnF2CBroScjXGM+eZaOfMX32kYODyvXuvF+0Es199b9VZFQFuENYz9
yvkGftA2lQ3mPBTIG9QxqyYIQBf4lVy+qV2Bttjd1qVvIqZo1uw8nNkSc/QSexgQ
8Xp7QJq6iUDhFJQKNKOpExjaWPQMnsIMjV0ajeku3YSukrodjBkX3TgCFyCEW3pH
mYtjOx6PfauLQbY1m3GzGwbLlJlJSCT19ieMj4JLgVZ9RZXBJGIXSQ25SSr/05mw
lJ13pULhzeG87HD/qTJLilnOxHb/2nmKTeeQgbafq6RfgJ8oBJQPrwjad2bwU5aW
/G1ieXwYaMbwcKOlWIDjMTd1/EEdgEJl6vBMK5J/j5wzeOsUg4thoxjanXS2tseD
ZoeENWTQZuUKI85sn1+EmEXTVNCAhizf1tZdqVEOZt8fsurMy5ajWOTZLVRwvsEV
tVuXPMgNzsywaJrlH/mcl6HSYz5ODTutIA9oDAPlh7Re5Lz+PCrmNFUzNux8hmoQ
DoLsuA/SDKwcw55ZAv2L4keP1XnO02qD89DfCeroKiOCfVETP99BCfHzrF4gnXix
Zc4awp1BuLjJuok8mW1/lXfpsq5vhRHQujAVpw6RBDhUvHPU3IhMhLY8DE2/HdZm
4GyVDY3mPLEHi/qXDRGCN1wGlCp+V7LTk8H0TEP0/Ak+AmWETNSWeZ1kLqa4ss8J
poslym+lTl2KnxIFr3DM2g3qaJtLTilVtbSkawDpWWxsNW64jx+OCAWr1b+2kc7I
WqciSAtn4zMLLGv9F5/OeUvr2c55aKcThfFQWyYwB+mWTRghcvFBI/2J/njs1kXm
BNJArozOX2DllQxwGS9ZI/6PgUKttO3pgp6pj9QvqvAyFDENQhQk3VI67OPtg9Oj
2F7y8LIndjl5cgWrIK4Mj4r8Ql3ZmU+IhgqEAi/rxzqMuC8XaeCEGdM9+HjQF6fL
q7qVw+686rcKxmofhp6wnS3HR/RuNwySdp1aaFQSgrDBFiHh2dWMHA/R/lzS7+SO
e2C7RFYH4sMdv2nRgXfvrNCHM6JhlbQc5GjZTY0hk0st2vEfnxRXOyXkGP1vqkaz
A/2m5e2yBpxMieFdZ2jtxQiUqqIYsq1mLpKqTqAssCeTaO3mcX5PZiLHV/FtyGSs
1CcRQg3snnaAbpWFglM8w8qF+EQUT56IvtO2cYqtL6TbOLgPcXNpkWObd1BTcx1w
amI28ATc6koJK2p/3KT3sYzmofT0swMtMPzyPdVTMAoIQmfq+lFEP+o+ObrbXxRm
IkmoE6cP5ajJaozNnT6kzHwg1JwrsmO1y0IEusH7rtP2qxENgajhpHTNBgNqGrop
EYZsr2Xs3GZp87uPZiqbw7B5xl95szVp1TZAy21FrAH3O8zBuGFDfaZ8h+X2SwR8
xNkIBGyfph6SejXtWJYPRmNlu7qRCv9+0eznO6J7bK+NYKwS9WCA3h2V0Flpt83y
vkq6wvzT+d8JKPSRb50ga6wSgTnH89ZU/CCxUqBjWedl79AZMHeL0GlgLZkBkFmU
MhhUrU70VYgKflZ8r5dQD1luwi1yFPh2++e12QWBLY/LagKYjSe13D/VOp1zFmqT
gX1aLSB8kO2p5s5JS+AL0YwAk1p41w9gzNkEV17gI92t3C4dc+g/QiV2Z6xeyfsQ
dtJ/yUK4zlT4XLHmgiOsUBzYsMBHIxiQ8L5zL01RhDfADqHDj9rsII37z3lP3PGL
fbAlgwf+e53AWeP7bcJfVpAhz1ThfODrbuLC8QJPjq8ku+VZHnIs/gWxG1HddTcb
YiKLtPdh1swZ4xNY6lsQkhqK25U4FkAFhkGOyaGilaE2kwmmjfLoH5Ww2qD/ZbWW
773Mw9RMHNNYOAqi52JonUfOOSLROq11Vn2QDh0ssbrmjAYurVolHN5s7L17ltLT
+frJgDgDdS8M4slBf8Ij0DY6wR9h0beorfpFFV7dhuibVqw9f1eCTvKnomBKTRnM
DY0Sv7XXjLHjnOFoB9mGGmxoQt2oz4cAc7LH8jJ3u1tbwqTjpqCog21sUXXkRhY2
lofi1cYDIKcoR2EiVOs3ATDbp3HoPgEVs5AzmjtHsc6JrtZuG7i7np2UnMfO0Q+s
lHv7MpNRaNwOTWlEthKvrH1Yv/LL8Z1yBj1w1sTGplbfSIW9F/lg4dkCENQZUb2/
Pvs3eeEIa/tC1rL1fbHA1JhTCtzWeasFLHIgyDHBC3xHk0doNlbg59H5wFUDFwQ5
DNjYwILYxzEfa25bjqjvl+l9smMtaWF+sCXxyHdXKPhcI1feGfJDWvoFT0k90Ucv
yoISF+Y789HLJrEAuMOvcADe2bnfb2mH3V/q8dz2VJmVFmIGUKdeo8o+IW8JFlYB
Rij1iJKHH+ENQd1UqkaFrnksGIYuYxpRxWoqXdQnLGWqJDWec/COOwHi3fpcXF7u
w+ywggIrj5l29rJH0cqVLLfU3jqxKI1nAMMwt1bMHhwAsg9EQikjHtLvlW+Gqw/Z
NgSdLIbubYwHI5X1lW7yil8EQqSa6vQFoki3msYluweIBUAu32JGvoOvesUVCgLV
FM34UQAKJ5+lF3N8851jHLmYYPmUANCkRQv58pSEQHdvgvNDnqryGcSDCJyfE0cc
oU4VRLVO32mL8RcymC85ezzmP1lusab7/l0e9dzERTIVFnxuRyMNJxWoRvx0YdJc
pppL+4JQoTOyQaRrz1Jw73qJws4iJHe9vIuz7wlcei8lM2vhhLbtptMyXG48dsLO
+OBH9X8aNNLWC471xvwALUs/FgFOvUjeiexuqJoS9ELeyPCHgIX1IzQUO5EcZEzu
N/tJvSBEONMxGMwP/ZP+5oa4w7fRD2dBHNgoWDPtv7af9glbH+LpiwzzBMlWz/sw
6rLpucdI6QuIJeVdaHe7GQWm0yC8RvbyAFKUzyp4CoH/NTFCNc5CTRi7u4Apn19x
K1Cjn97Eh6ZTu6RsmFFoOT2mbbA0Dq8SxYzTX63f9NUqdw6fq8hnOgRVK6oQjwT4
5F2gkkjFOTTqLhaVISz3BMs6NAYMjCZLQIA1wUX3OGU4BNXydJbYpBcmkd/KWWzo
u4BixIZ8jDQ+e4b1T3+fG+QdFw3n6VOme4V4MY+6GD1+xOjsRvxYLTlkD5k/3hUS
mZkU21frVOMU4OxWLp5vZOjef7jtdpTeRt9DGN6H7cm1lGPOPw1fAIpPv0dj03pk
NfaLscDP9AzRwYUfhy1piEfwrNUauQMJdK57TL+BieHFlCUrWxzSuhrK9uUvTtFZ
19GR0kE1qKCy6JVbWO12On597wQ6funWxY/PYjHfhfeP/5h0VEhGqsLgzyspcHvx
fx7KttQ5pxdcgNuysYGa6WXh0yJ1Uxr/EBXzJM3S3AyTXD++1omQkPLmjDjIc/bA
SeJnZFa7xE8koGUz8oEsb61v2GsWiMkyA4y2XvcVKXXmRwOrFALIdges/ST4XZCs
VUfNNGIQiZDJvdiwb2SR0XuPuFgrWHyV4I37iWhRRGMZxU5o5MymLlKQ3nZQChq8
ex1zgwSzmxl9yR1KVg1vKxyAH+x7IdLxbjhdpLDbsfH8V6GS9ISJdWfc+E+qQ/v6
o8FwpqPD6KAWz5yBLwSIn76S0h8nrHuG0mOinVIJ1jb/sp8oQWIUG7+HqVfsEzGs
E3Wo5m/QQ0EFsqOcbu+hF4x0oE2dTdzQaTCE/PwxV+/YysDC1O5IZeD+EcEpHrd4
oAjeREZw2uz++77thjtvnMyEcv8se/BhZPmVX2K6t1xyIDmRhgKL7ywZ37DyIYnZ
Rp8c3Wd87pTPUlW08mshS0y6/6qZhOOVnCBbbDqvfmIYWmtt+WF179PCi8zopvRh
9Mw0p3vT/6ddYU/yW5rHDGKk/VBrTgTuPhZWqiT3xrGmNjHPgP3HbdDF9UmPAf5W
71YPVSu8QbbhZ+chAvIcDUZNI0NboMe7WWXwcM3FbaBPuBAuXwFwePhUF5XZPHLJ
MtcWt1iHjX/uSeFSON2mnCcBnEeqpw8gRHkPrFmNlLTG5UqSwnw3vMBMapCqpuNe
wvCmgRPofws8TrXRbsddFgVkZiYqm/moU+Nf1BKxFz8ejswrI0OURRinHctiyQPs
rCX0okzChWuCMKTtPZE2vfAYIsIlvNU5og5zlGXXwOe7FXi/L6fAM7KzoKUj7CUA
AkHyKYHks+k1C3aAM6BbWLqVKLdml6xkNevHWE/M1ZY1bR/Wm9pFV5DM1kjEKdQX
FpbJ7CeYSAArie0MQgMhJQnfRPNoXqJ1QsJRPSgwVcm7cOb2mFrn0LF9iHFZOmJK
OmpAHZ7VwE7CmDpOLMUYicuyabsroQXpeQY9KzLGRuvI7mS0pAKs9IGQXHpDsFMO
E+zzX22j03qUf3vgkEJtEwNpOjVAym8vaTWEbnC3xbb3/Jhjz6JvPQAWFZ7yWC93
MzZb63QCK6qcYchuvKOTSgekoZrLt+z7qO/GTIjaiikntX3tLEAyp+UdlhKdJYge
teBleVV4dDL9E+iQQYH1zX0KuOWxuIDFsEBLJ5s5Np/pKc6JfBe104o2KUhSx/0Z
bKGqfOpUzgwy/0d80sxlsoZkWSDav26IsS+Y5fGGCkvRV+OxwR3nh42b5iDpYyRe
eU9sWpflukfhqzB0+xqPIRQWC1bGt2JT+DFP1q/25rdMhIKRUxJloXHxLpwdv3EH
1oZ+UTPlD09Y0zQdh05k2JmeaRwefworQgGXigFXjXoNi4OpbgDZPJB7d5cqwEs2
PCF+gcfMPaMifcp70j9fZlgZ3s+IAuNeeI2z3+X5kLUnEbCtn0y0aZXgKrMxbxzk
/NPFZcLfwoNlbvpWQF5D/m3a7lxB1Aax0CFWQMD4AJZrmDAMLaasVCoGte5j3vpP
NEwMgdA9mayq+X1toENFrB7Rtj2sXgqem/5gu9DZH7pbWTc1fPsZpomGTHOsoaGU
H/2yPrUq2qR/rSJiJ8SrjotFvu/KY97W1P5kHyNOqo8nyfyb5JuohG0dnCEsEpbW
lzsGySJPSa96kv/Xk8yAyN/MG7GLWPR1FYp6XoNGQlVFXfXzhKk+aE8EhOXUnUUU
0okEp+C8Xo3uI20XnDEINbVKZnSyNYoaBYQXgZi6pbgumrkBUOdFMMOcQ5g+tr9K
sviTAOoCIQR1cX/QJb2KbZSJ6rF561BRLzNOV2/Ik81+ndYJDBEKCPamwfUt96hb
wdE3mt7BsckKXwyUxu8Xyk5sPHtJYbcNCPlKYUT4Gp9TJm7jho+hhjcwuoGfymWn
2I0vWfccSRXEenUALXR8xMvmHKBwU4o15RVRxJdQSfhq3mGLc1iAw/kLV29WdP+A
hHezBAnUuhYhSaxuIhG2Rx7dmDX60dHxhR0szSRPeTzpqwwGBzEEs3wnthWvPxHq
oG6FtloCbqXBAPDPm+cS69kTrYtTM4OqDH6hIpifCb2+JXAiYT1oqLUOQ0aZxT+G
8FKJ02cqCqSR2+7K6IEfcECwT3ZDBueQBjFb4mpUwOzyz5Cqfv2yW55MKYzdXRAN
ooL1BD1hNtg898qEwEAzDeSbpKTW96qPle+4DqvlZTggaKyUefudzilNnB0Q6mOK
iER+o5OJOhIdtBw36z/azibe6681KR4b38rx0a3tGW9UyLNXvzJiBpLEdSCZPzWC
2ubNaSndskA19UN72wEYb7oL6EZV1BUg0eFAmCkwrI5KcxaNm89ea7ZUUJcDao1U
PUxKJDpOn6JtCUPY3eLsdN3B7B9THtDeHLI5iBnCHBuD956ivOjH2w+yUMUXcHJx
rKF4ylW9DdB+9igmH1b0N+Wd+qvYnZFnP2aamAwU5eM6ApcDLHEJbYM1Gqc7P9ig
HW11WQwmhwWZfjYaXpXCGsiCtslayKzOjSGemCrVYHF4I4u0Tn0knYvpwzUHemwd
4jVh5LQcLc4L5uiw7y06U5Ic/1vFwprHmzlignCqCw92Y3yR+bzG7TTbeTb++abv
aR7IdvCJWQ+oxjdgcP/0CW4ehOddSb74uizUQv+aGkn0wz3CRAZJY9mJmu9voRB9
2ufO2vekkSMTHdZPDJ/UmOu7n1cDPaTtGZVFxkt0k50CV3TYP3lysCVcdZ/I52ns
3Qke6YBNVssvffI3MMKcKlIHfOvsHPPrEzC235JDpuy9Nj89/O6raqOJ5+8Etb4z
4EelN0WHUr2DPchIpaj81owEGLF9QSVqYBAHD6kUbhw6LL5KSVDhJCJdWYr+GAdm
Qztu8YgDSfSxtT4Vrm0x8NR6hRoRS05iTllVkLHBK75Dt/TBocSkpeKpSjhVU86i
vltJMj4fnxuKyCAmHetufjb302gSc/N5hxtCwxjpX+6WfVKSmtuSm+SGYWlCaIig
gJB+R3K88bGHB6Xj8m2I0p4Wsb/JgUyO4I2iQ9fCoqRvnlnF4/SXJlHogGOcSOYR
m4/iL6/UKvU9xfcDVu54jGfhHodJYrXPmU2e9Xm/XrtTx3jOJ6HlqC5Ruk7U5ZAo
C+sNPKplUAL1JQMYTZKHxFXQ8eh/01Ho03ZsAlVfHkqLoBnX6nEys1tviFM1Z8lD
F1YIawvcYbyfslw5w98JpnnFwXqqZTTTmHgm9jls9dKj38Ri3tzyMIswq8Ishar5
YKa5IgNh9qor5TlAdcRbCHx0pc+8tEcsUjTgcidRNa8QkwgRMx74gl32WyrfvVtJ
4LsIhY0qkhvWTpknu8mB338k+9B6DgIMe4RGSUbEk4YjnUKCHg3WiIQy4YBunLwc
wyjS+GRthHsAjdRp7WFJRCmORyJVptWbkM0yRpSDpDML+nIP5vQXT0oXDrU0ucFt
fcIUYot917fnlNiGXoGWVGL08QAV2bxS23/yBwjv+w+QPn+tfIpKePlSqcx54w1l
yRkWy5pVc323jXRSykYqgsIVkJmAiHHdMdksMOu0HaDV4EpZMbcaqMol701U8vUh
X0B1NGnPXpVXhzv3OCoZFkZitY5WwEnMtnV15VjkKp5Rx/fSNCwjDmAm7Bka/GUF
MSAneOWXw2Go1njNdcs27I+c8tsIl6hgK2mmuRWZLYMJ/g7GYoJGzyCa7VzqC1Uq
Zy09AvaAEp8RZ+mSkCvgJATW0rpqCqMXiWcATq2/6P+mT7bnlkSEGIBBJ8YZ1Xq5
k4yh08iz6X6BOAwYW9hmlgC8V45ck9UTEBXbxXvaXqQfV/obaD4c2gGFUvCCOu48
PosNvTB5RqW1rLCHLfeOoChnHasMu7HzcxVDvdzks5K9rH/cQObiBsoHv6BWv2XN
j4x3DXA0wGer1O95y7gTEdb76D84svhxb/n4oKT/LRJLGMT96bV3ArFvHJQu5XwY
to632wtXw8XYdsMg8QhkLI52i18szealFbno4WgmGP+CKWzKSfgAELRWd6eq/MzH
pNjqMyjkKEEYF3RnhOusne6RSkiFroH1kBYbQWqfeJ3gpQ3UeSiLOIPMTx8sLHaK
qI5fr0AEmHy/qckF1rQlw6UfYHNtWbIiSt1/Hb/g0cjUKgtbdTTFReSnhFoGo6h2
JhEE0DZdlxpuSaEXHzpNFAEbvjpSLY9J6DO7av0vyu60nvSaMwre1/A3lSedNu8w
dxrc85EhcPpCm4yRhPQM0q5+Hs5QJBJ/wOb5VU72HW44fvV8gjyQXWLVjSKTB9V7
Cn3ltYJkFaWd85takX0M1ZV6VAvlWtywGv8rWIwy/7DqJoDuM3waa1PdBOwe/1Ul
ZZFUzjvAuj/VZ58fb4ETfeM1Uz3GuN9+dVOXEw9k8OxAUVXWUAww90XTX7/vP+RT
7eBTqe8oubyifo2798ereLR+l/xEHQPPPFlOafs27Grme9r4/Rf0dziOg2Toxkg3
2wAy/ZBjBnu0v2TY3yYrtywiesu9azL7iUS6ISYdjNPvs8+d1cmslR0Q+bN9u3Fs
d/GH2nsQzQ50B3urNzRQb1HSNU0D6SafnqQQO/JNIjxlqmgMbKtNRVm1UNL8MuQQ
BkdLAZnJ+6apev/eelc8jhXGdOR8Ar8r+r2ZyXlX8ylpDG4270PJm3mVWkrhRzLM
ygS4VGCfnSjfVa6X6Tk7A53b4qP7IuEy6pvfYZzH/a411ZW+TCqb0aSBMW6M8pnW
xgdmYuvZ19UpuI+peNESskOoKFVRd7Y3Hdj4DdDG1kBgmx155BV8NafKzZY4fCg8
UfrfsTNjoYSXbBm4ly1/ZRdwt1ao6Qi6XlNV3tMBmYZyxdaDYpoQIHwZRi413TC9
/iwwno+Fu6QKQ9xOa3GxOiX8sSCAfwa4+PZ0VXCqNsBnUu2ySYTSlMYVFrclCuz+
BIwb9QH+q7OpHG5ewNokecHf45y8wLJ5xrq7VFxU+YQY5Ap4V0mKN9uQOotFnkJk
/gNq+y+ZwFc0yTOTwqVC87cApfiYgGx5+UGi2RPPi1dsl+ec4H6TpGOS2rHaAohE
tZsq4Ju6At5JHyRS60WF+ZQkpfbQx0o+O5EaY276P6h24boG3DxhwlliTATyN7r+
vKXFOztD50G1jQjIef6ltLF3Qh9ZPNCpP2+IjClfv8UnEksJWbRFwCyLF9URzM95
oHEKEGMgvY99jJRWpVobfkrabEMpun4NSzhs3n38AGsIh4hhLDPr6IZEbwICbTH9
dx9Mr2igGW3i92EL8JXJmyIcj8luJi7BvCEeOlAclyqc+jGauV29WxpBt+DNRUGy
6P7ZnwZgxWuRCqUWo9pdQtwv4Sa5Mb+dzXIC8HJGCxAxJ2Vp1CT+DOawFYJPfmJe
HIMFFiVKdt2i6Uh1hAT6mgOzAqpEPqn5w+4zgJn9cGsfmDbeYAkFSs6uNNzxSafV
IlZKBvlRIp5QvhsBDj8y684rkB9TzU+iWkYPL+A+6nVYOlQ3CaL0S8oFjPMlUml1
GJ+6Wr4mK8Ptcn1TKhIJOZu4Inxsju9ZrDZyLO3CaKrzKZW+XHFBpi7kVRQkh33X
fJjq1mI+vFZw7NGsfE5Zv4/SeIF0N64HkSLn6q/TuSf3fWP2vaCWb4vEjvI9atyR
w0NhHvMJyqC5ZNwcvHm81BBsqxyKmW0Uj1D1aiSD5f9cUdzozyaRHMQFdIsT8M1Y
3l+IBLsih2yeCVxCb9GJOgUTrGVf16AMQEIPuJMhfmb2rAs06Z4yoaFW922bkK5W
CDceNGpq8pl8Sfpp0VwPPrErGX3EybM2w73WUwW8HriTYIGya0YXGrvabr5bBwW9
pOfxV0qzditk40dYtfulURhOvz/l1Uf9FyDWDl5tJp7MmO/0Buzwigu+C7OFuXE+
1bgzPswwjnE0wBXlQbQ8oexwgt6F5A/IVaM19lzHDLv7cFTpHoKE8UW0Qr2Q+Gzk
tLOHNXMciA/vBlM3WoeLbt68jdC+aUNUCrfptVHdG+9UmfhqGn+72KIHAz3KB7gR
x7q/HEZjz1fk6ET3IzudykXIQIO0usiEKyBzgt9X+RFEf1bvvATMnAA4DqKWGqs4
zmklApzFKeCfaLeV6tRwCMFYcmtHzyEcoEAg74IpWdIyJR2wDYwMk1Y1ZKHbcr0L
0EKhoe+s2wzoDOLDRigDKKqQMwrpAEvUqen7hAenAeCFVuURFwBEdaQse0yjH/ke
5IfvXXAUJHRPK4b1eQmjxeB6tIjDG9zjq2FAwDY1CBCYplpAbrdNyMJ714xD577S
W0Bb6F+LqM2RTdMqDn8Bs3uR9QeTbfU8Jo3HaTO/SmFUe5qFW6nX+PKz/k2UkxSl
P87wTfLvZxHg9zHEqUCFdnCSp0A7ibrH2O4dna4+NvVCkRUr3U6lSTVZZaL+jbBl
4UDNR0QD1D8s6IN1NjB9yyy4yzSu0ba4xuoxe2YYKztgUPW8axKJfJvywVvPulX0
gdDX8f72xporND5Nh4VTV5mvtO1Iv2S1kWTzQt9aeXvA5K1Ya1gXKksO55rtHqBr
dQmfFdIGrHyRk+XPSS4dbdFrTv94eW4yK89boQel8J7Grm1vX+sepbbOQduwlNAt
WusVNDEMr280WQjSN+yEEHVzAKKvhb3kepGl2LYlP1DhUR/yruWBGFbXigPoA3Wo
F7hod9n/qawit5BlRTFwfycwF1KktoEj16hLcIZWd3QC7//p5EUn9bvSVaNhuWx5
5T/cRkiQ6XrbNM+pWj3Ji4QgggarLjOrNUSUKL5kb0Omnm45fXgIefAqEX3cAWdw
dS7C+2qwI2IZAOrq4EZOMCIga5gVaDFM8+I2Sw9TSnpNILP+Vy/sUJJ3FlWOX3YE
8ifLrdzQB4B/EoorWm9475kqQlU3sYSTTMjzCb1Uhhk+joW4jrsp9HDnFUp1Pl36
h15SMJ5nryYu4eWxTsEtfqwbZs7LLIB5r56eWuQL/yKpcj+Ek8Y6ySkOCeu0U8pi
WBaFCmsCwyLFUaxMHW2rza6goGvh/C0EWYC0/Hx52Vq0KnR2x7C865X1bhhSFg+j
3QuPZGig2al9b2FPArm7oTOvGi6jV9JefqLZpGynye9heC4vlnYc2JGpigOBrAhX
7Jtj7/F/I37dX1vCMb2NkZNwsteW58bjghamMHgSuexe+QC9fBcADUTXd5e4rL0J
6C8D+w0P1L2WsW0rnBT5DosRtCstdLuLw75qoBoeiGDHMdKYVGqHl7Ibxm1yXWrj
4u6CjQ3EYAyjA0Ty/FJhnBQ5BRWqh/I61z7XhdaqDCZ9eBswIDR0lmOJfsq/n55r
lvpBKSLUuPNwkzu9cd4pcG/rQachHkzGGN0yfBU0yOTW2klA6mMOINdLLt4Afy+b
rmBeabXJ0KZ/EPpDeIphDUJU3BBmqC5OwvrC4+ZbPDM4UOYkAiQdSoNNNcFJ3wvO
JgkmF/X7J3BIOC04MHCg3UayOaUtbECztyWwZHP1J1bQCMaKAZkec1O2L112vGde
PIPcj2iEWt9bHYN75y/ZgN6FuAdat4DSer3DCCVOszFNuG/4mQGki+vi5ICzuYBX
tcJCbQINfNESv4z4coNBgLpCZaHhpTBq8pQvJZhHqTJCDDOzQIvcsJZDtK2UJkI1
OZKv5KioVJ/QRyN38e5xKuNzPYq0po1wwPqs8J5aPmzuruM7PVknFpdNN8U7zwwq
d5SZEGqTlQWuoLKypNx7O/02dBa2c1Zlgz48pmf5fl2o6kmtCtutM9uPHxZLeG6L
U69XGhRqo7boEG5wNN+7Imsd6xkaEYzSeC/62HY7iJa2q3jdDKaaplls0L81I2z9
VCqIQTTlEFoQXQIiUWhQFBqSQArsO3boa/yaaIQ2b+svsKV7YI9te7v/aoQjn22V
WevkZ2qBI7/l0ZAawtIIxUU1vaygardGlB5dnthR6oJmH6s9cZPLiGdaq1+iBzFO
a5W01jccJA/jXNwuZaPZEYy+Ua4BUpelyd3vxwGkL0Tgf6UCY19bo+T95dlKIK6J
1iqT2ti6xnRx2hTrKf8k8BPc8sE/VrWtHKYKo55YRYOeXbnZp0PhcFMZ5+tUqTAD
JJfJIjhpH0uJYD5N+slqyRqpKt2h8M0vE49GmFPqfJv0qjZ53IWlCQSn7lu0PyWA
8t2r7PZHGzaH7gCX4ZGn/OT1vnzc11weN5GqH0tqEkhENKZJ0JpTW2v9FwPVAgUv
38u0FjLP1tvvozNEgjRY3PtCDVExsLqLPo6BREI40LX/YIrGxbj33Rw80pgmSsDD
WWR4pK/lLw2z/7QEtRjMvLuti5PuvjbkMtjoi+MxR3Gkte5A6XVCZVxMfHJV0J2/
aFkqFpmZpAbPBIk6M843GPi0UgTOD/K48ZQY60zISp8FZPiAXMaZBvar8i3rlqCm
Bhs1vXBK1ufvadwwg2mlTf6ShD1BKor6migJsuTdMV/9VBK1zlpmAduICi0UlJhH
gXtgsBeWaDZAwyiQWSOiWbFemd3YUrOnBxiBBAINb7jzKO593ETengT/SDefs7MH
BQyhELByirR25X3szoGj2lDRFazYrs+tdwKiFI6AmdyFZcQFeRrIPRdUinK9k3Vx
cSz16cIXXif7sv4/Yk+kSbdYb6N4MTsTVcaPQwJPkfMWV1PND8pHv+lSd5zAKKYv
a5ygVFBsObc79vxDGGNwvOw5d9z/qeFicyoz4YbxoQtKRGqglQURx2Y6gL1GenjD
IBf2LENoHP2FCNEChvCs1yG6c03LhJ/M/N4aeX6Y9WX/+2ZlN1WecJmlKfK3X1uU
ifEHKly7W3vKGRlhwUDHTi8mCiax8m/9F0kQrHPdZA1g1524vD7MHG8zm7ncgKi0
DRhi07A06tBodE1S/0M1AE4FTbBsW1/GYPAOc4wEgfBFlAY+4ZZe+E/Z/gRhTwUA
ksMpEoAR6UyZG7nuhpWxteE5oS/Eso5b2TowC2u1SyXq94QGALHKlwYl8sFUzQI4
SnnHN3I9jYORXLIKtQQIEwdTEBlET3tFwpwTnJfwAFooODkkIDFJzOJGRoN3f+6p
7hXuaMvUgjOpiFASRBrsOHW1MIQ1zUHyDxykEraZ6WGt+8UL5YbCvyeeLgHn8kVL
eVo94kM1aLGrzwUkEHiBTmvWjlnRNtgCE3qa6ewa9nhQHkGwDZSUgC1FlAzLrgUQ
D15soxZnAOlIf5JxB4owFcRbaHSHNXZH4uSxSkcvDcGx2Gyea16+DzJfhWwT1VAX
hmzyQGvA7FWFjHbsttwVRlXrrxj6MJqhsaoJi0BWf4DyBRP+6zGrBgpgjPmIiT0Q
T3VJ2deoDUHEjAqxVrlpkMYqBn1eOi6RoDIgVhBb8QOU/4DdrFkw/RxBaSEm3AOz
/fRNJGzgZuikFiQ6/o8j50VZo1stxtHLBmPAWrhkiMppxxQbU3/4g1kXm9641akt
SMH//lpbLRWovOjaB2C0ig0bYM69w1qNC9OlcXnrX3lbYeVjrT+CqD3mi0qzehWh
r9y1CDEtjaE0faIJ6o+41keTJYlu3wPDdFmj8ul/9TG+vpsQ9eVw4cr4EGkl+qT+
uzuUzZ7MOLgPd+fH5FEb4bxlSa7tPbCucG/+oU5M0amO1Cf4SLp7Csq6Ouysz/1B
kwTilLmrCEXYptawyrYYeJfXABI8nQgjFSvHyeaXGM7UeaAuzWjTT1TXMxOj+E/9
B8Du+9Z15ozbcC8YQQkxZ9+Ok1NIMjFSQkT672HF61cnxW/FDydVFpa9JPF0eaTH
UANCtkZWH111ec6FH4ZZ2b2k/nKO9g+nc3w3nPY246JOzVzK6gVoOIC87v5H4GeC
wGx2PAUV320PMKSuibOxPVru1+dOu56C7JmvTzCLKdblhpEL5j4gdj3r0N36jKKI
MVMHRvsyp4J7sE9NZpMU/1wRvwatxYxUbT3lBQLegn52VEeycLnKKyqvObV1QDhy
xcvK1dJXOSALm6xyNvZdSRWAimnoil1NkR/pYphbFDxwPisZhXhB7x5nB1I/2xRK
IiFE7kOA5Ejn11GtivGr88A3x544T4HVSNH55TGng1tBPsCgZ+NtD5Hv9A2ssHM9
ahT+d8SWGZ/I+H4QKEkrrgNmU5Fxu8Ah8dKwmdjda/AhGOZPE06BoC4cs2L+eXfU
knQ1n1tuzUEVTRyMnTqhdB2aBqMSM/ITW38K+w3bO3KOZSe65CgoVlgR3duRmHRg
wah8tLPyMcpLoxDV84ylQ/lDqJ0uwLgP0oCkfE2jtiauo6Vd+Dt232Xf2Qi19At+
VIdi1HW/YP3b27F1V9WYz4OryUSfbaDP5mi3vMGh3BegG5NqdSKRNopjZLP2ODxR
J1zzWkeDrzLfbyl4nYSslLg3T1P4WCHq2V4PZZd732et2y5spUjCP2TtQhJi0Rsd
mrh45crkROESGAwZxT9cI79/j5Dxm7qyRZB+qjfsJZxWDDGMYzEGtDdLAMgIMJiL
v8404xs7oy1Ukg7DYCBETBaBJowTivLozdr48vhuJKFg0s59E64JHguwSh7xDA+s
nb9KO6MElZv5ZKjbHAK0ZhRAuQiqpdoL9aU/cAmaNx6mlkYiKjqV9OgbrnhE9mwk
QAocGdTXHml9nRCwnRLipBuRuJwS0HD/krUPHAASsXS7kEc3yKxFMUDmsMqFzq2e
f+R4plEOa2rM1dRgXTHpbgbCjb7UfWaKGJXEWGwG/LWBj1nNjwFTUuGs9GPmEsoT
qF/lE8laD4/BKIC63T09ckpRa8nl4ACvZK0Ss6qyjR0grjsE1Elb+fA37I1uoVvk
bFOW0Bp04OsgvCdPVXCR/gN2vVh7igHkAm4qYQosHGus1bQrPriMgFG3GkMNg0xB
pvL6F1xHeFJtpWzLcshxwoT/i2VP6hcA1whB6n5jmSl2lfCAeECz7717sG0u4NoS
fVJJsrPR5Nw0NVxMYhqfAoGTIr2pdABOyftkn9rghmUkAqBSWNp0VRlqNyU6zdUy
mAjQaBOvTDfLmbb9xtVLBIeb0tT1WUn4F+EKjakUmgAWCWSZG4pzQuqpMItsoYFF
rGOe2+oP7pki3SQNDbVFz0/+ykPgJ/7P2mv6bke95sgeAk+EhbikHGFuVjHbqNm3
GHGDUKDJiN5uWvd2Y8d5bEzxjqFzzblfjbf+xYi6ZHVqw+Gh3nW03NMn/32sqkvA
bz1extpOLsCeBBJL46JhxfjfR4Sf2THwHmy3rOvWFtpRAkMFRtZma2Cz2GdZWwtr
dUUQpy9QnjdVhkanodiEiwAiwAfUPghs+ADQVT4uMtwHV7LEBlSfXLOXVPzMkr+h
v//we7P/iL/NDf7g2BD4Q3cbTjS4OY+5IFwzd2g1nP7x/UeoX93AWdPGoLOcL7Pf
sRZ9CzMBnfWhHgdnjKeXUXYbwB96WLqPYaPYclTYwizQimsGvCDeHwQwh9Lu5Y3x
cBP3Iuzgy0+nawYfe3EbCB4SZnLRXjmRH17m/JiS/rXqMYKfIU4TyLVTje9Q3YEB
M1PrRSKgCtMfcgvZ5lzyH7vlijfRXtOjbUSEjXSGvcQByKu1A7Kn+AfXoSWqJSGU
uLf9qM3ryZtkNBkQOxwA1GCVRDK3gBRumqRKWC184l5R5aG/FhVQOjxFp2f6dPoB
4b2UxQYh5bzUzolbXpPzLuyI13eeoXhIaE1qvRxxW3dtIPFVPqlY9NgyTntAtDrW
rO2doayXN3j7475H6QFKi4dnS+VR7fVOm8BZ3GmMktEsmpbcnj3kfpQ6nZE5ySeT
3krZXLnEoguNydjo46sFCGlxu+bjSrWj9fO4NtEy1vPdlfSKPeTPcc5Unv8Fi5qc
mj5nQSpwTMRviXEIZGTfJ40ocf5LZz4rNXbqj6RwrvKPW4fubHymyPe33PJEj3mU
fWXU8Ne6k44ZYyUj/2a8dpvoC6uMzF4O7GqkApaMz1e7JfevrEomfllJl5p61oby
Rvuopxu+RI7v/tld9KuqteUvjoOHQdLy+JxKptbonRh19z6zAFI+W42BlkoQU0Mb
KA7FzauDb+dU3Owq3XKbNL8usMdSaY10VlNoOSYB+NhQi9vm5TOqPucvFBUM8JTC
Qc+zLTCXU7m7miK3LmLRDPLJFEPnbh5UhQRwUKvdwUzb5yO9Zr56Zz6FeWSUPRWR
Y7l8NCTtJP5aLhO/fJvNxtUGfUpZfXpV6KmFK5wJ7XLsA13cB5Ga880HE9tYn4U/
IElCWjC6RMLRIlFqLIs593SHUY5Z2/h1nEN8Uhoi2JAkBHEHlTgYQSQyWTZItHQm
r8TfgNXXmiIR8dyRvWrTf/s9I5ToFWxpqPQrhzZ2QPZwjFpFrGtOVThi0MWVpHLk
IDhhNcv2Z0Szfw+AA9I9/WfkxMMbpLrlcgaVIw5QzjVQry12MpeAf9QES9CAAMy0
cPZjGFaPt6b/xeOUWEWi+s3iV7pi4HGl0vBmXkSk6TOkOiQV1DXKA9pt6c4RWUP7
bNpBtdSALlgunjplFoGP15uvZBTia/z5qQc25DOZELKm1GUCKUu+s6vnolE4oABV
ZOmkGZj6URNc6xW85yzKVt/jdxPInoRhwox66djNPFYoVJO0lX/vADURs2YBMj8L
LVMXSZdxTSGU0Kxo7w/bBK9RfxSn9hZpAQC8GGd8cf4VOlGSowkx0ir3EHuVY+rX
uDxQkkLKvSxQzcqZgbgHHfb0x376kBFIC+3DXRw6wKCr4G0j234bVYDXMDXJnno9
6JGlLW5ekcjCC4jfCsd5V1ddowP7yCF6g/2a9lw0URLdxBcNZjvmw2oG+JsWd8R0
nJqJrOOOir5iZQRRJ+jOnXwziBkrATArmjEZSu19SDNjG9UJlOP/pJGSi3PjryzF
yvwS0rLaACslQLAftvIK5Iwf6LvcEWKeR+wHVrDWL0o+Nuj1e788U5od1KBfGxY3
b4UNI5reFd9EAMq8nE4SciwpnReA/pzEIw8pnhilVzN4PQOlPaObqPJw7xAJ9ALW
4Or5XOrduTYCvFmP15lzvsnRImdRJ+mGHnRaUrurAcXpo6REB7c7S7JGq5/W9qKd
svr2KR1awQE4UZSlwoZTFJ720GNvv8t6tvTA4EYz4lh5jlY0FtycnTPr8fMuQXHo
hYCPY6CUqLkQWtk6I5azvWNzD4rT3ZMDg+dFxB4zi6CuGiQgXk5aOVMvvI+YlzFs
gkLzm73J4N7ezDXPEKwPRKjFGUFm4Cq5BqT6ZFhIvCWsE4dywHSbOctr6HPI3RKs
oY4GzGCz4fkN2R0cKCDPCQzcoJgGvJbxw25b1MvFZZs4nUSzvMIcfml5uEDqKA1U
U8NYS6c62R6RJlvODcHhTNXsjdrF1Bk5YvJyGSzs+CHw2sThRIlR3kiVRhZ8lsSJ
RSRaftANlgMo5gNcYGq7O1CkI2tQv/s04Z/bMbcZ0Tek6DxT23xb+FHPP702aYr2
3J20dud5Wl0U3h6swmUDu2dDrbgcKZ0C9IoUk4yRB7xDexTfIDmcUnhaIptMvpma
py9uixIbyb9Y3gBPlQD5996dsb2E0MzjpVJ3GGY/SXS7gmod5DKZdR8tppG06g5G
rtOdUzjya7tJT8gwpX0kfTUTg4D5tHRcp0WjLIaMKoDWiSV8ev9ITTknQNYZvQum
Pi1iA29N92LSvr+c0LXDsGLXD1rONkz/pN41iY2Lx9mXP8Y1NEIbTtwwzd6dwvvg
/Cl/LVOjQehF90elg92hEELgKcZCH1PTcth9IIBNIbed55dfZLtVc0ooUyxa2pSM
CTjrzPVQ4DnrqQMnG9VkSKf29cyr+wTjgxR3ZWsighLXYxSLG/VVrAImTIsAvtDN
V9nqqROR386IZACGBYkY96pe/KNqyQdEISxQdshySUheHS2ZpJCb6omX8/he8rNP
vrXe73JOVszzlWYSUrcyHFCHQnPaYJOJPsiMUQdwQXK5KwE4SWKGoxe8/kP+LoIu
8gJOa12J0V9REUDGArPGdDi/ZvB4/OL5nV5XpGpQjsFvjB9PN/lB2gDXUQOmaLm9
orhmgwa54s8kUEgqtFvXfVFKnzdsju9Fcn1KkOiz9BOm8g32Z8CitQ4b1KcX8ACy
V2X5UpImNEeooYDzJ+FqGIT6f7zb/L/FssN5gZJxWl50S2qrLLx9c9S2G3c7uGFN
whyyhNOY4ibFMjOpKgHmnpXdwShmhSgfbQe1R9SyDvuvHO6q6Yl7qHNwo0F1VGJi
7SOrRWzNXuXQm3tXGu0IS9UI0swYMqc4H22OXzVZFGf54f8qLBOJIk1ItsDr3LvG
u2m2ORFAFwzcgBB/XjRdbmop/UJVuhoQ2nhj8bNzHZriR3JxOn7ZOKew5kwRJJko
sDFzprHxkrEXl0T1GKQhYaYVLlD2GiUB4ONGGK4kF01XQY64yY4R13A0weJSkMl5
SLFiAUM9hSh0PjZmpC5wXN8EjwS77inlBfn72QWLYSgiIZXgsMZMycNupvgoMVk7
CA1syRRX97lx7UjcChTRKsV97u0dm/rRfmusoruo8vj5e0lSdEhIMUQ1/D5B/J4o
fWZYUEABCiJqR0uE988d8ExgrmUhx60pA5HZGSpB5S0Xk/jhijgrObM3Yl8XU8Af
deSOAncqKGkd92/pdBSM1WVKsH/P6ASxx59yrderKQYWEeAKFmU2cbjv2n43r4YY
JPohru2N8WwINJ+u6ANr8pHtOGZq5NcP4EJ9nj7gABvcvgHB34EgeW0AzJIyTRXY
ncuXVLp2f6yhnlxAbijBgeRHCvUARFErvIM96rXpDHYQCNYUkrg5NIU9e3UOARjB
0YY0I2Fi5ZDGU7BZLTYSOKyVnj/tSK1+bA0O0NVUU/GMiJazjc1lKfAEnxWRhcQL
HTvY8J71hyIGcc+QasVONzfTKnItOEuqwPNkeIvMZBl6He6XjldZzBaWulEakCbp
uBWhI+7sWW6aOC04vdv6NRkpxE/v1hG+1ybTIBbwJA/n97BLMr8YuReZW7m1xKdu
AE5vV0gXw9kTEPsGz4Rr6iGOqCm0ycv0VdrcLclblzui0VY9KLejpiBM4I/nr2uN
4MKRywUYzkRqIBn7aL0/QvYLBpNCXq9jl4evqlbAFgXm+Chb6IsscPxQiHWd2AN/
hhqHaAhx7KFIzMDE2lTQX48zIGwsIa4rCFa/rL43T2dC68DsgFZkOiLgHiGd7igs
ya50hxH0GNThDxFXkHvK8dFs5dSYOp0QZngss+nbL6WluTRUPZT7PkAs2iE2Bp/M
huZUt5DkNvprhHNuZLdpIcAhBGugxtX2v5/mA6SI2Xa+p2qsNvtMeR85YIOb+8uj
VESSAhKgIXOcxTbd8a0+gLa7SGtasilaZ2ILSmbztC/0Mayhd/xNcovB0Bl2X1Mr
FLzKFfx7KAxk4vDNT2xFqEyrfLSSzE/obSmZuaBl1LWbZw1hMErA5ip5GyKgyTsU
VrXvIKDWeGSsuEofP459XwcvAWZ9vyAOWUaGa/q3sVu+YqkDHwBDdwxJ9ptLjFJM
BSuK4oMjQ5RTZ1ai0TREWrkmwsJHjOZ5o5ANaxpxGcRc5VG3HrHuIUPaUnsPVuaK
C38pIFky6n/epbKul9WDvPx0RRzDtgL/YMk4yLZmYTK4Kk2QXkqxpqDG/hCP6anj
OfFUrDfIe6Pbo/f81GiZiKp8Q7u4E+one3Xz1+mDPGKMma9vgx7KF5OuueJ8dP1m
GnJ2DSTfFNMgo9lJs96SCc9XACQc4RVGuZIOb6uBeB+6v2T0amoQVLxTs3pY5CCT
MxcyQWFnpdXnyr1W4AbYedYAHd94voTQn8PzgGmN1DelK2Zh1v1zQFFMp1/huCuI
zXdf055t70ZKMD5gHdDPrHVInp8Za1qhyTD+7VX4WVr+2wlGuDSOvzTQqbBOOJ9c
VP0KBf+4460WBaArlVMXewsLCT6MB2TRmfmwTe9Cd842yOfFBOsLSGv8HN4zGS/X
65Y4XwrRNAh1BpkodV7KUhysTEXkde+gDhEhaBXKrEFH8Hb0Bm+MSHQxjnQE4jwE
PDFrfAjhsM6ryX415fvOpX6nEoQ+N+wHjdMtXZHNPPJO0E1x5blQmdK4dhVkYC1r
AIlp7DhdGPFGNxv56TAod/lf3E4PgOhR9n2C/mNxAivTyesqXlCAtwaG0osJD7P1
PCB2C3VyaRAesKdlGSY4DEtxKC9gBuFLwCCYJnsFCNjL4sv9Gn9Gd6WV9MxCMoH6
LwERNIslM6uRRwLKgLf/lIC3Ulgk3hgmRtKKjB7zvtPzd7zDZPOncbJ4q24t02e3
58ZgoFv6BgZVTJoG4mKJBAzcBxLnqJltEWUSppNUPZAm06L0cUiu3r1pn0PaIxB2
W3qTbxdfvi52eBwlIgxtxPqPqJmgacq3wv36kvtSkJnDkXzjxp1qEINvzKtRMP2j
Y3EOPeFrR1l3C0VnezlnCSEqWbz7Rv6yrw99Sjaj4UosLdcNxP/+vF5slepe44wy
fxCI/kOdx8meNk6HhO6ScjbmXEX0OBr0eb5n14wl9ymzEYg8MhIXfBfzaRJpjr+d
FlcppNy9cS6qzQEBzgx2gbnco+OepV71MJvgEiDJukfw9saVWI16/bU4JI23cJxJ
lk0WLRLkVzD5tUeTQscMvTsGRVgjDmW61Mhkw7ujg1FkcpyEjqtMPr40U/cWZMxc
RRpDEafVAYUszqKWu6jtjcLe+D6pRz1QNDCF8hRZl4nvJURbGj9rpwnzHiXnyIRm
XF2XB1pF21W5lPHCtaVgtp+/FTMIyyA901ZB3yJRpkfsSz8bj7PmCjJ7jaxff7IA
aB4/pHiWGDD5EXoR0P3DSmcewh36PsHE5109Cc7Y0nWVB62SXmD8VB8Odj8IEYvd
9QPUeZuX/nA6n0c++XbK8hSZ9bOOegqVF0PuEVEBmoB+aXIrBLhdvHyrZYMk1KGB
6+Wpj6BSgeUzd9soHgdM8RD7SiPNqPYEaTMS6xDAbs4wvnpsxga+NPp8RFlaHOJh
qXxuPhgKUfKExM5nveVzZv5gROjHXMVHM+2Aq50P8Ebo0g+knG4BSlmG+VKGbJm2
rYs+ElpK40ZTgDjDsdl//xz/IxXHkQF/UfOaVVhy7Do3JibepEHETng2jqF15gob
W2aSzY/Ky2fNRtvD21AwyHyGXu1jAn08wQo8fgPk1SmTXbNqiq6cyhLDRxDvmVM9
p7HelbdaGLQbcxct6QkNVNw04UUJjSd4pYHBQy98CDfOWPIinyfEwT6JJZceoqex
ALLOnGdtarH6coiOriQqbx+gk7APWSUjg8xiXGQHC2rTBOV1gpgZsBkWrZGYvwUa
uuUuLzaEu9GsqDR6Dssx93oToPFR0KToSOePLDH0Op7y0joxCrU1matlaPL9dlig
wypxu3nV90100rvqywaMGqM04nZkrutEz5dvayN+FCS7oOc7A/4OIYVDnfIA9ZkR
kWeHM/3TBggZ52CwiqQxTGyl/neeKQ8HNVoidLtywEMD46aQKNLSwQSqMasSXnnb
xn6tLIxES9/MbHR/ujLqQ9vrQeL1RjyqFIsEanhnM+ejQwX5Sw0t6/UNZ3i59VUQ
hiWlP7iobfqNT3wS+JDuNNxBHCqmMkGbxkS94x/Nt2hlL4uOV5iz9BW/wOy0m1oG
+RJOJymfBBHQ2EkyVsqIkSH0NQWRQzDUBXkz7/nsl3qV/EsHUIx5Z1Xrmirknnl2
8oRl1379aNH+yofjN3pywu+upFdnYThz8j+7mjtD1BCm2r46T5ONudgEXXWgJAxM
ami0tiSX8f0/P0s5HX1oBvgu0bDacwgqkIQ6S3K7iI+kwcPdspxJpaXX8sVN8O3Z
ZfLRrUqP+sQP2EvZl8bzj9f+x7Kq8Y3GLodiOpjwzVb/BwzvuzV3yFe61+Fpk8ji
QyTOGetOglzDHjTruU7YUchVa0cRdChqUjfuNWHNVXLC8pNBAvQg5QPII5n37SVb
CNXCgTrJ9zIeHzENJzd9hyFSDXX000l3xzowAAIvlPcPXdn6ekgJTMJzfeHFSEIr
TZRMkUqg44nh5cXwJTejE+FugguGZES2vYG28mSWlrQlrJWzx506ML1zdnfr5J43
Vujp7WJ03ITgiVb2e980FPzIGyDRJXK4AzL1jy3G4liRelilG9aAPEXbZsuBMIxq
+VBuCRznTce/myRxrOBsflNpZ/MPaT5MmTdgWxByRKcsBb7ZbCwbURSD2n83WdXP
/xEzLMDuPUlTFTOfkyS1XxzIyUNUuF8h5cFFHiSro3wRFtJOxCc6/PYPtW86Ogdu
gUgP5fjVyC79gN6DV4VKF1JVUGC4F9KPU8E/fJdUNSnYTUO6gHukKRNdxLebXk8T
G8hg81evRGAGcDG+YdHns6ocpcAu9Exzp24KYoWISb0aBxj/ruczTZuqjgfEiSEH
CcmUp2N4gcqZ7C1vu2qZcMYr5BtJ4d4GMGffRw/B3WyDWXBAwi5+vzkzHVucohvc
l3gx1NszRj3hohMRnto2/VCzE+Lw+vJrlqAqXVlpGQlFb444TFBWCvz860iKgiPY
85xHJxWbzVrdoQkn52o741SqO8oUcudKMtKlLf/OtGiaLlbqxwg2qFejv96kDbtH
2gwSILIIHTvBZHzqgX32aghkX6B6SmY0kleo8oY4olqL4+4BBxiPlZWSwRGnSlVt
fbvW5bG3cTFYn2DSXu4lV/vSHVV9xoenxEXHzY25YylPo3LhFKIFJIxvrq4VM+EN
37hF1LlBFZ3U42hgp/9Rncmvker/n7Xkb3ogYPUQ15LGOvfnNbDF9iJVgx965bQX
knOOTiNLwqs2HQ5TScyGicMxQSlUrnUs51D8K65EpfT5DmrwxksNSISZ/tSr27Sg
fbO7VnnIcZkzhMFepO2nXmEzWvCZs2pv30g4lPHJwbIMdtO12AfQnaMeKgFn5xDY
mAFmIZqMdDRUCT4jgvMe+Ii6hL5aNjWxeE1nYVWeeQds1MqP/AAGkOX4RW3To8tK
Q51Dj1wP2fcZPd4JAzyEy/AgQ5dTTVi+HCxpFzPRBOdWXaC/rikzX2RL4/DhXxPV
xxK69OkOqFMrtwLYl+HhqwZFv3KqNa04Ej8VPbaNYyzq9A2cveHm5LAtyY/NbLVb
tNTZp1X8ztUkG3rMkWTTGPxM4z/WoeZsjRIwQqUY498IJYRglRIqGWH218/8nevZ
Zz6spviTk880qkG3FXROn3YQLQD/QGtXTWOgCMgUQExhyMeMEU1xmGdVGks3uAp7
hIKT9s/JSmvDg4iEAXV1q7sEBcSJoEry53ti6yYu2cBxf+A4AMVSGc/teucNzBYl
moTm7BFiD1To83oKLErcwKt7cW86R+UNUsVDq1Vx9oCjQcyneMjaxruYzYZQJ+a6
j4MnoqhZveVEeJc58nsPFWtaRp7/EQK6kUO4hubeNoMXHZOdGoKEC3siD6dVqjmu
J4STx3FEjyZESNibVK58Ij03LF0zL4uLw2LYJZTCIVir+hPnjYZ0VK+upYcouZFS
L8kU1j2LCU1vTJ/wV1aQDPHr4eLk8BLwj536WdvoHr6iHnO+pbeEvf5BysYbyff2
vPnZFEOpdgE59sigJSIwbbQqS40LoYthS6JxBpyTbWnNKCpk+YgFyw0tUTnxpD/r
RzuSY8Z2tIRNbodx9QIziZDh2UGhtk98XLt3QeYbkIa6YI4x+D+GMVbXm81YZ+L2
o5CkhBcsC1bJ7+cwqDAEpw3gHaA8blf+W5UrjrKcddvjpZUlGB540ZFv5eHnDg5P
O2eP8Cy9xsRJ6OqC7uhCVTeSX89+J6rSR7wgIE9XE6IkeS0YuZDUjqjAvyf+BKI5
3Fyn16r/ryMWLNZR2INeytWgyg6FR9qUOicFACdqzmOPQYp1hOA2KDIh3l+ciKkJ
HAvTD5Rj/5uZc6SoPoBsu9CCvo/MIO9Ph9ZVcbjhm/RnD6NwVCtO3gqAwV7G8D5H
ZERjvTRhHiy2vcnKDW2gcMSvq/YzO2mhuPP2TZP5pw/EiM2WRf61GQuKPvJoUK1T
QEjtXAsQZeNri9hODGskGb2CZlLhp6eOW9bHWuLeIQmiJ11uEU2upif41qMGWRNr
Yrw11xyrju/nR1jgT8tghn5kX4pSmamu1Wy7Qyb/kXeqXMptUapwKmK8dKydBnj1
bLYcXzwCpFO4HKialRxkmvGc86EJEV6qkHUqBYYaLttWFZhlEZkPRJFJG7Rw1/fq
Pth//FCtKFf4cDNYR/Zpvt58zq/Zen/nL5+vAhl/cMEmR2DT1iOevIH5c8lutxZX
wYpcgxV5g6hJlm4hAyvuHZ0HRl1yQzKlua/B4RHUGCl3ybRszQC7El+sfCFxybaA
igEz9r4P3zq1qJ0LCjvaUo6jjKJFBHlSx3oFW+Z1CaHvRzi6mq2QhK6Ssd9sQD+3
ITgvcx7TIoSIfS6MzAn2m2CrDLh9V5c+UMAcuC7WvHHViZ9c/nWuFXdoqA4QZFt5
9og1xV0KSw1DT4O+8CUH8ZwG7bMwWjIvUInsc0M2r8UCaKZgfjb11m24ugMnCvpz
rMuBdnYcD6adRw/RORHy48Fj3ushCA+UiH71f6vTD3h1v4UayK1F4MqILzjLFBxy
UokUPpVelCJsgNTTm0kq6QT6RHExWvQ15yY5B8EpFYkigkBxrxYSCUDGPAZo+3Ar
wvPEVngKI+nA6RZybG8WDIBEzYeaXBY3hJUKhtV8vpQUKiqsCOPmy6jFTwcAPSDA
qOmJR0k86IePWr/0RcV0vMHb9VNgj2NW9XSnVJ1IIhW9MMIvQGFIKZQEDz5vA3zn
Gd4RbbxR5SHKxlbsRxE4ys07jhVGMiG9J4MGmosOMK4lHhw03g51ix1HX7rm3EVy
n/PDW/iqkG4b3hg6jmAi52ofZ8gjXZits+Ku+K5D40gFskhe2yGka8PhA6WHXwX6
SCPdxuyIBEDmmqsRVXUCtS1Vx0BsupyGCtYQzLn4H3lfaweaaLeeTuodHbbk410V
Zp5KB0rX0hOjgPurZESBv9MixV6qpi41071M0XyjFL4UiGBgMVg9i09hhzuujlz2
L2g6xaZoG3A+UlP2AR+j+ZXCLuLDUTRHZmqT1oH6GHb1UaqAACFrPFy44zxmRwuX
AvbmFP4GFXGCit+nAjPi8D+whErvhINhvBYTUeiUT90Zyusap6l0smvqdWkm6+Kw
pcbYWDMi2Rnrk7X/qQ2oDOk4LJDwFXrYwTxxxmTcZuaT/q8kEu6f7wm+zKFTnvvn
1w1qH4vHA1lciJCJ/mVJoFoVo10iJRWWX3txpd7zmekqPy/eRLE5aaw1br6HRyh6
SHcFLiH8IOaiMeuvN0YGJwoEBNRCuwC6N8jndT0nUbgM9/SAJj/QR7Ewm0o9q3vg
nd3S1HXVwM1pkkR2KNQN6mTTdx84EK4pzBurs1i4wL1NDfcJLd/8PFSYKaiY6BDW
99Gie2Z9d76qE95n9TqqbExV08Y0FOgxsazjwa4aTBHs6Zlt0t5EZSV6m8lYfqOp
LluOQYZII+kMX00PXyrNlaEecM5h8J3yqddzV53AMOLVBjp3O+m6xgFgXBK5IQn8
LSKpChxNRKOT13Hc6ahhWcG7mIDpE0o/6BNWDS4dpE/NXJk/68ofbU13xlxNYNPd
9lncq1u1MrYoHxxVDw4DpZKvEiNGVa9EH3eiihJgwKlJ0AJKgkTsmztInJB+Qap1
iBvfBCDVCNXXroVb7Gc9jp3fflDAhcIa1L/Q6EsrW3CWxccB8YT+8v+423MgkPYj
VjPW3+u7Xw/NAqUx8Qgb4ImP+B/aWWTHcRZCSswwA9Lq4kISy6X8YSPe6Q5PVBOG
6lD3mgKH/6syF12OhNDtAUjt+JRIVzBkurYQgop17fIW6j1k13N755/S/GGZhYQf
W0sIQL6e7DdXne1Ng2196QmfS3j600IMFxivuW5TQw0EsbfvKv83YCczZvWkzSyB
2r4gRX0FaNneY9v2EyajEBo1J2iDM5alvzuzB2KeWQmMWxdgjFXuTCJ34Q8jmal9
crSQgKmweR6TDu5OfcGYu3ZoCMRYSCGDBtI66JAnoUwZX9ofTRG0VDpIEyq4t29S
BG32BvbnN4bQy/oyrQQqb03CSMIx03P1W5GKpcna2cak6E7u9TtAB+H+a4XTh4l1
a3mgh/6nd1vrASFQX2VPabAMP82OLFuq+LD/1mnZRut/bthe09brdL0ip79R54Ia
+yRI/D0ADd6pw4pl6wX7UeEROpDpfzYWgiltZruWwD9rq2W3DNfUDyQT8Cji9NeS
rvQCmIQtibrkAskuivK16bg0hZmaCEQYxyhdDSO3x3ZOSOLgzMixRJmiRLKe0mfp
PYsYLwZXGeb9HGNu6pOPSOfIE+22B2lSlwPx2lK72/H4T6x6nhTbfjavBoz2BUQy
2xjXzdHka5k/Lr1F0C80xP32w2+f4FTlcJ4qRzSwGQ2a05HfOMkDnzo0ZouLcrjU
GZ85JosNGfX+LPk0ZDPo2qojL1wYCF4+/beN7vzjgUgiHbRKyWVzy3m4PfxB1qji
KgYMkVWdQhWkHuJ8PIdGRpMzr4GbI2LjULpQl+fdqi5nmzbUa1s0SwZUjrWlAWAC
67AZ0CTvD+pknyym4mOo/iSYtu7tSRfxeZabU9YRTRfo82zBjrkS7XYDuQsqdKCY
KqWoJ1AWiJn2bTXj+JbIBbVge6Pj4BbDjd+wDuBVsfg1kqVtghcxARGuvEuHwomt
BsKmWqkc9Y5UUclB3KVjvxfo0hXb+w5WKMmx+ruy9dllfTmVrCewKvgZalyRwc2b
3NGrrE//2zViLpZRYK9PgcjvvWSKK83Fk/1ZA7vPPPCxdtFBUVfMDsLB9abn47f+
5Hxb7o3PTYElkjWDCdO74bCnqcl43/XHrxEva+3Zjo7ADcjUQ8ab2Xkhnnbncf/P
+D7wuThv4thcXBC5gsQRkhoa2l91vUTfoXEy1Hpi+OLWPmMOtZLlSkJmxae/ztgb
YUEKO8oRzxx18F7adYloS87Ye3b6P7Dj1zV6KVBpyp3dbk3K1Ad35Gu48cI9uUI/
h9zHgZYrZhx+rv6UCsL8VerKVmUKcNldHDCkSgZZ4Sllrh0sCWq5l9qu/DKVqIFW
ZIlA8NIJQ5FjyBSohxjpiHKes+7gFRwuXoE13KWxbsPupnlsVIz7lukxt45dZRQX
4HxYSU2J0j6oPzzMyiflu4z7KwN/86BcQFu/NPv47O1iP2HhuCnYMQjc3FPpEUO3
SXLVFY8kOm5Yj67rUGpAqYgovK+oYLnlNYbD+lc4DZoMJX6LofnDYcOKfnUOePvs
s9D9JNBA+Y7glIbvzFXo2P7x9FwE9gVBNl3CWYHYADvmTa2tMucag7+V0TnYmkgo
qejmRGID67cHoMUmRwOJCt/ln+WTRK3GMVwxqmu3YvSj0UM/GOmX49XEFxMfCeI+
Ahzd6TEAwHIvMa8EIPuJodux6v32D+fu4lWJzVGkaBdz9wHPzEIe7BfhAhYkC+DG
kdCiOrwmLgrYNDIIFz6m8G7rGavum6Cwke8kEsK0gsWxSWMfdbI8xDIMvVrWDNxL
g4ZZrHA2VFtZq3ayRHwauFBlBTXpqJVcMjDogmHLoL36UWCBYZsu4l/2S8ej93XT
lUHx0b9ZHxvb7TOZVqdNTnumx3VKd8eXyaMLe3T3kWWqS0FumRGOmCZ6ULqWNNDt
GsuNpHaG4mqTCkyIroXlCJ+C/wwKxulb9UPOYv2IgkBm1L83yu8m0BHesIX6BQGk
G1Jj+NhM7aoc5OTXfRbgI2LCpAC8/IcsD2ZEeRLrEAgSLxQ1oU+OTALiJSfL5Ypg
sxhuLrzcTmMdAXJjSbnejR0OBBQWUPfhDqLfEN+uzPz4PIkhyARUcgZNm9MEtloz
MBb91L2nksKEHiVZwybyFCaumXG35/EBfyDh+iTRxftgz2TxVc69tl+nllMTr93n
Up3sR2FUfIx24iWEotCKc3q6SGCwiNz414vP/ikvyjQEpLQMtssS/hj6hDJ9yWCf
vkfuRH8BbwuWwoZKES0rFL3lXEXAficvHidlU22m4S9Pc4CwEFZdVIl5AtmUJJCz
FEtTMGnbWLdpDqFsIYb70IeZrTBh5mZsNegKVXhBQ4oi5pZXL075hOgvJwDxpX5b
RPLtxcVGfkchZLygT3Hlcp0d+LZe1Wyh8bTzdZQcM1u7AqWc/Zia9TSoCPUJ4dZ2
UxM8ycAt+9vgCrQMfIN6zkNyL+7RDo6fT1NIRLqELB0UZOv9hv2KlfUAA5B4EbYb
naoxYImHfhun/ik7YdGKZ+/ZaqlaRpFeN+yQHRlSnww1u/wfuhFitCZDdY/nNrji
uhJRb9NH7X/wpOJVOj/FQH04OArO+tqGoEO2ekYG8MalxAxHdD5X2A1Yy06Z1Io+
j52hzphrzFfdXMhAu+ow8qgqx33oh/8Kew25ZCsEQmSSxiDgGJez/UVd7KopkFjp
W1u594qp7PeqDLenDuUlhjpsuch3kXHNXErDzCOZ4YhD85m3mhnK6g2NC6AiF39X
JAGKjKlbz610U6C5anzkbfDhliOIBvxt/NZOCzvgpNa+i30xQnAVG/CGEHgasyi5
aEqbOH+oWkGQQMwneBBYqTFQJG+x8sTZsLlT1jYQmoQX6JuLZz/9ZbmHHA/KDX8O
buwrIY3b8iZjrRBFzJuMEfb05NLn/eOsF0/NfXaLr1899WjZTPXcaKT3HRn8lvpy
NnpCp+qxPGTWhoEN0UJqk9hz0aot676NdKE06DhgLRpY4PbBmeV+ToKfBPW9hptS
246Y8cmaZ6KhfdvvaC07GXV0PDmoUg5owkOpxbjdzIjhtDlPsG7rdldHjyeh0ngu
Fgrau+jdDzwbc8vpEBD3S9tkuI3JUCbIqs3GyMhOMVZGvxJzv2KhzQ0Rn5uUYp7s
oPKzTvAR+K8DQ5ul87YUU4DqSVOFoYiBg26j6szuQUxM0/D1iXA02FnbdFr+F4ww
MJp9/j2N6abyPbD2IxchgLFY8yF4Ban19z12KvUqyuF6bTFIsIhYFWNqrekWk1HL
0WBa42ZpjUailb5e1WAe/tP/gSVZhHpjdc1Pxszgg2N4b8zi0Xyu+T7orLLqj/gE
DZmy6R/o4YxdmVRaFTbsaWkR7pY89tVEKOxxedNc7ZqbwlYyWFmlgawRtq3STVlV
2HIyc+hKUdD6cs2HhWmHt6bffK+wzoYlTkBPg3tugtC2TECiozO0uHIJ98H4Qokl
2zdEnFeUOjG6pbGn3fexesCczmLrBzO5RJqyD6pObMUsaNGJ3cncnhNN/cUpjL4r
wLpLHAYlIe6ZzWu2bdsleXjgO+8AJqC6tP7sGSfHrj5Q9pnpRpsCoVHFmomhkLP1
lOD4L6xxuQtlJ/uFODlJRGCakHPpnrHFipgbloAnMcAA+K3667QoWprje4IseUfC
OqEfCh9lgNJeiqRx3igjKeBVrtk+IGIfZdA2ukqbkZP68K176zCyh+9GTqb1o1M9
HIBRphgQkbNeKd2Ht/dncHMN/aonttmLBqRG6PjqHdY2e3mUzN78pBZLRne10JX4
3b4JaZ/qR5rw+cxFyiqv5rrYvmeM3vDzad8r4eLhwy0gY0TAqv4cBlvJY0ZgBcfC
XmzDQkjMQ74YHMJQoiRZYcKW9MLXHSb/NWO2N5iTsSdKrUeVg6xL1lvv44HPiXvA
Nnd2InMM2RN6ALhZpqWiRIze5r2X5oR5+hXk0iC8J9AH1yRmHpZt3aoNeM1M04Jc
G5TM1OWKoJpP00fBdoIxZ7EUk2S2jiqxIJiR4sS+169e7X2GyF01yZQs6pfzEluC
zPtlhPUTOH2jBpD0M+qTQZfwZDySNdsYV8ey86DGQOerPUI3J/H4pMIEaIPIF4WX
leaiUrsHcE94U7W3ZUG9OZq0CGyOU/hTM1YZaS7t0pq9yePr1IC+S90U/prUeuGd
4uvjWkcpz6KfGHlT1ePLTbZp22woTKbVZa9l1WVQBshrZK/lj4YUJSsyu0t80MIc
2QjLbg1adzJPyOP1OII6eL8cj0gGya+VsNn23OhhPVIEkEMDJMMWCiTFhkOf92qa
cUdXivmJZBEDNmqs9slO+2MVVkYIrG7PIUqHsj0tH8OYgJ+53DPsC3eczJCBRkjx
2tGEbExdkr8O4U8Etdw4dBIAbZPPQsssXgY9Z0jrMEUz5geQrSorCnQjNVKesS8K
zA+K6sYRK5nB56U6BWX8zSkM7CnuX+ehit7ASstxB4JTI3zqoN62ZnWmR80hcaS0
0M83RfF2sKLTJz2PcSVd6Z4VxzyYVUfx8XLysy3/YvMBvYlrYeMpPPStMeR6BKsc
p94AaAmtbLsyaD/me3+SLmtsYj2U2gJIrUNSgeX6CE996tPeboVJq+K2EDRLRJlk
kbuVtyCVkOql/HaZndbdUtVYFGt+mPOGLQ0Bj18K+fJjjdz7FTZPpRJzOZscaCio
g2g9TbTTHFRwNPjO/9CQr0QPDLT+iuJ1JMk1vsk7SnUQ9oB99YyiGXlLoWWLici0
8czjHdy0jLIcpASJ9X60wLYfg9QfuOxaLQSBM3VZJVSB/0nQ5o1FlTFMoPB4ZixH
ClEEIV8fjazfx2Q9RTvU2ZMSUMG8Hjt8ojlIg7tSP5aQhzdZ+zkUYYCsFSKxFJq3
KUgCirz//LkRAh4zNQr8kJXIvGN0iZWzmPvSRX8PDh8QC0CIGZfXylWoSzVXciJu
dzUpDXJjM6dX6SMNRphNjpBnPbXKnX0XCSFMBgzHD2bmK7ftpnNZYkomvt3Q6X2x
QayQeaAQFnNKG9uZg7k3rQcybiIle4842fahRAeVjZm5qWRohfehCTV/fvN/YaDs
HvqWnd4JqV/O0jMYN01GH2YPUqbK3pCheXM+8+VNkfM7bbeisQC8C75Vk1SX5EdL
B1GYRUuGzOuho8rITUwm9iMdZbOFXuIgkOGHtuQK/3zTknqgTItR5gRboOGL49Px
Sl9cHtKuoYBqcLThs1f44f5TTiLzYp7GaWyfbiXMd9vIfZUZ5q0VwCAggUpic5iw
dqzNeleaaCWP1SEvtfYYpJ7qte0T0Q60K3wmEMlNTAuY0n7UZf7ThPKmgw3a/qQA
0TQxMHPcRxN+0SBq9nZWZTsir0CwItjCiK1RW9KPIbKhFo+c0Sf5ZIku6DpQF4/A
5onPq9D8Qqg+Q1SIVaZZiJQl7FOFdVM/r8dYjIxDX/D4MvNOulR1TPoC5PL9Q28z
+WxzqJsyJ1s7SQOi4BG2leRbq1fe5+66cyE07z/Ors0DJ8dIeoxtwVn0GRp1Mjae
xJdsbkXh6/NLjTok7W7od6YTIVtvLHVlqPIXb5pyvLfxYs2btiHKFMPdRZiH+hR7
V47Q71eXYa6w0LVCBmAkn5R2xnl8g7VZ3BqUp+r2ZP+/gsC0hq4Di5ogx6n81XVA
SzYMw4g1xy1FMmfeK6XBKoDN8wah1hp/YZGqrr4wD7kx0xFaSazgS9SbqIdd/RNl
FOuciW1BxA07MsZWIjF4Kvg1466xjx1WNglopJ4Gc8TnvBOsyp5I6QtSVniAnFPW
3bAuQRDElfIuDONrX9E9L+GcWmnfibKurj52luD3SIDqc/goW5947S3gFwosy+9l
zjkBXXa19EVMATRHzJXnbMh3fz8mx3t1mJUDjoqfjXNb4fK+WfHxiKdVw7c4Pov1
9yDpwxM0HIc9yrCd8OpdJkv1RVT5iZTRJLZmqvhn878jy4DCyPLYjRS2nrjxWRFn
c70kDYNnWd1UhwNDR+8MIyiACIWAOBU5Us9/8HF3xlfyArIanaO2Ou7t9uljMwdH
2edtlD40MXi3+ydQCeZdOjcXNXt1QoHgyTzOalUzlx3bXgbPwjgGrU7U+f51Cz0s
1ickn08IozXiLiMg8eRGgQ9rV+xkgnIgrvMAjE8vz3DhXH+FUE5MHxkBlCVBeFCZ
j8YKMkqItuaJ9CPltrNxh0lr/VMfssPf+15Ae16wAfoYOlivWdPoy9BzJdQSJUb5
O4eSqFjzLUVT040PZ3ZkMTKvNZOLV9tqhKQxEoh4bOaTijpu14AHvjMBpPHqkVdy
a2t2NFr41DzVEVfH6Ti0QsfOSldENAmssTJ5X3Fg2Hy0EBeMVPjtaYApjH10Jp8s
TbBMhkwNbUlWzNTIMCWr4wWGO4tEQRPyZxu+Kh8s6Op+BbX0wyv2sYUWdA+H+JNC
SesFThc0zo25KPhNsM0PMnocEyUC/+3iHGu5DKJKDuAs7drifDu3WWZvncnBwIPc
Te7p0/yRgqkrjTTag1Quxzy0o8cu4to3jT2Cir8sDxMtHLQNkwytzqNtLh/wSutu
pFVylRLuHeP8wYUZjn70fMGsy1G8PJPeRRkrgrxUkf2KhE0+0FCKqIaj6NtuUQJv
kg91x6pN5wMKqYnyKhYh+mq3CK8A9/EQCxxBhVY45cLIi9cmZRIZzv1+k50Zjtn9
JUubnD/F7ju9bf+rXZfjgj3rovvwP9u2yXozhb3UZia9HJCbMoaLyOWfx3CT04QU
QMHHwqzSOJOR7JIp87SBBVzsCFHpP0dcambDwTMX2OZbati8u/NozZjv5zPIBqbD
TdbFTu8aE8FGO3EqtJAUlX5R3uUuJwmnsXaDfs2c4ANe217wey8JyiIaxzn3Vqsg
hoFyjKl609LNfySjRlf/vw/tElEhkZik0YrxvZMFoWrP9p+jAj2wMaLrXW2jd+cE
c9ieGGtMv6oYuBM4Jf8i58kAKhxwy2GJNoHxAYMTmtUvylRj7BCmqPfeyjF+KnvH
bsypR9qW9zENtmHQPMTJS/a3wPjLSIq1rWQK0FVhLTVtRY3FcN35JGUXvfpI4odp
XW3Vd2gYL+vinXtWZX3Qojbw5N2DuURBjf62Xjidq16K15JvCtKAJn7ZjIoVycLu
gWQf/QJHqS//qBtvKRI+PNmrkC7MA7cWRmRXj+vjD9aiIR4sweg0wPTO+eY1Cafd
vLdRChgW06UnjyOl8sHOV2hmwDWNhzm/4bLx2o9ILFAdVApNl0EUXJDt9WPjg63d
8LUk9/gkQwGi0JcmGlEGhrBX8tZ8erAs7kYZUY1iCYxBTr8hxliQW7EPaC4HhmNP
FSfc6/zSFFXPQQi9efFIVEYUczHXYXHQAZ6oKukUBaqDxymat2y8CjgpFeqLDde1
JjBH6neDHsRX/BhHV0liIF1d7tf5iQU4jlLMPOxEFU6gsIc+rBlSP2wDsiPqZdYe
8osD4si0cRASST+i39l+TuHVal0FLR5HIHzbs/B4rvsgvm3iZ8LgXCC2CwnIYwtn
/r+aTRbovb3/dkEdPO9iX1HiWR2SMFLw6fIuD0q2+6XqNektLFtIPJlilXjVQDuv
8oAyN5WoQc83CTceIJMxbcpwY5AGab0pJgx7RI7QCMOg6PEvB6t7rpW1XJKogKBT
4O+1lM7/9gFAyjsqJt0tQv69S0Q1cvtoVzMOy4jlILcMJ04Ig75Q8WrBvf+8+aP2
YQpHJt4ehJ+xbOIIg8KmH5dXJXiCcKl9Azsj3/744xcXGvSvis6El4s/u2DI0616
RArG2rBP0v4Jwuj2h+RRoKPIZF72+yVQTSCN5wxTwHVD1QmsuL+FyI0K2v5sKpQS
yt5Cn4ocIjsjat8qKTlVOTCR9MG4MCzGsVWUJLWxG144tz2BHe92RnMSgRLMQMwI
0J4noR8gcEaTS0Z4UW2sXy5aQaX8rD7Vvwwaz8HbndF006x7fD6KY7rwXOIJ8W1i
/mOrV4rk4iJ1m7PbRTb4ajQk875EtmXA8Ca8aA4Pu9OJS9ovFHh1w+PVPONXza9j
1wiwfoKWc7mG8LkT3LPiKQKIMdm8rO1hLjOB3dezkttvfeonlyZuE523c1G2BCMl
mClCmXSju6oS0FDjigghZmMGdQ0Ye0wN5Rr5oh19bbtz5QMeP4a2nbeQd03cPo0X
DJbksx9SKJ5Fq2ZzOheepcWyP3g2jus7XptViw0D1lrYLbI5YTSGan93JWgmkjxM
Z1sVD5WkfTZeyajdvhujgEtK5k8jOk1UrYCfGwQGLAytbXgtkdrxM+hE0Pwlld57
MOeqv+gYZmwzut8bPWtKzGGIbupjrkDApRzG/HsULEhUB0UZsongLU7SIGmlyG5g
pvUDI7wwXjLGahneWzvq3P+De2/NNSUe80mnnvmUSLkyp1g3JUYVs/D6DsE4c0R8
wKsI7yTpdl6pLYwp4wK3XzpHNfaYzhliWhuhOhs2DwTcNiP7OtGiTLkog13U9Yob
upRfXh6xtrMeGLeFkxbYRZnXfQq6/2vZ3hZKD5KILvnb3nNkjUrmspF+rBB2Ylax
40+3BVqOarEl0nU3KDSg8dFs/QLUfCdqhhMzQYTI3u7QBmc3yGIWlc9YAZIrvf12
4wS2oY5ftaLFfrRJt4KrqimIDadZ9SJEnZekfXpyE9/3QfF2W7Xrm5iFpmAiRceV
pkxlsi5UG67G6skL7IfuLGnb/MDWvmZv8OxGkh8lRvldNgY7HK3Xk1uen3XVFjHC
9z+NNMUBgsV5w9KWnpE3lN+BbTPqmrK/xR0D1GhKhBMqrrR3xE/xkss6Bajfae/9
PnIG5PDERS7UaCwWcN30Jo5ZpMSDZaM6iEF2JIKhhM7c+mQQ9kjxZKturvH4zpB9
ESoRUH5siiUcmGRc6mEjieU8RaojVoxr/3rK7zBxTRGLdVrYb8UnTeSQ7RIL1rYa
f7fwen3tn1QC5owLdF2VitMlwmIvO1SZ/Xttc6cvNxBPAlOFBpc0JeZNMxP79RsW
2ZJw75TzybZFaQq9i3cI6XhIH0uzBhWBaQoBQw+pTe6eWDCHjZDoqcIXR1CZQiE/
XXxfR7KteXuWZdrXSpuXkBbZXc++YChfNHgf/pYZRqgJsd3AlJIXgOyMkL8d5/pO
LpEgEpekcBZvTmva7ssRx5JpqQQR1rLRr/0lMzBBV0P5za4KjBfDePvYJ/WQDIQa
I4//pEojEluyWSFCGv3mmUNwDQgmqAqenLwOjmnL5DoVJ98eIhBwKmAEnRuAstu5
svI0bjXqBmYb/558lTn89OqfZ/MRa33Cej67GvZyTMUcDKK+a027tG0RfCcsU/rt
WQUv5uycl6tEHikvi6TGbRofEJbasgxDOfO4+3usEDy0vK2xKSNKLddc8YjTZQ/b
iCc/YjNTVN15NRPssL6GLS9OxXxFzrsl0lC9cQEL5ARh4A402n0HzEcHmk1p4w1X
IMD5HUg4o8/kJAGbvA0ylX5CDpR1M8DG/VwJ6M/EIy0nEdK5nmJCo04qPC1zYn7t
U0kpkTF++HhH6uEUd/HlX7UXgIy8qCxxD668oiFjaNpLEjb/6gZwYr6kr5gKw++t
bYqKLfXD7N9UcFB96nxoXc8Xx9QoYu7S2b3yw+EbF+aYSxAs4QFeZMECFenYc9LF
7Kg+iY5hu/a11n1BweSuemLtL5bAhP26P22yMnMFNmnp/Wtkcur9xKIm/N6rO1bF
jwFntTAuxiNsDUZDa1WySDlenGkqPHQljguR1DQIUCir0ZdT0dQuqdqHPZOfv/eX
33mG9x/IS5THd6I3lYxXcs9sNPkjxeyJFp8gbn8Alz2YR8BvXThe6wlBk8Fc+lPE
GpcPIiEfV1fZNkrR2/wol8hqSrwMAxjv80pju1RIuTVf5JieDxpBNn4vBXLqERGH
lrpgUQ8VOldkG3ptnXV2lpGK3hvp0q9NeHJG8AlNVTkbqVAnq6yY2P1qmBL71MWd
UN+B8IhClSVoUZjqqAl2K4234EA05RIV5GPp2iP77vYNBXSbxYWvapImFivUfprc
/g9tm00EtCOUDWUI2dLINPhSdzqE8h+vxyfNKwFZOawmGtTruJsl/kHsauT5JiYF
+fb2DUGmsSpJXCxg4XGlz/CgkuqsiS0OyKSTP4YyvL2IJSQTe9jGORyT2GvYV5s2
FQRJdpK/ajbZ6VeSjohRR6fkpC1Dl63RdYsQ2FxJmYsmSjqUddIbZLZAdZ5jbpjU
XtTfzugbQQZEnr/RWHS0RRK6TJcR7jEy4jzefDxLGYzUeu+uLgquY0H6JdzRbVbx
jMFrdNBiianJtQo+mAFUooKi24rzBAiyVFWw7Nr2k4i+nscm27+y6ropcl9sVVH2
2A4uRE8V49/VGANhQwcoVzFleBG0oBFSpXzwxqc2BQGImQKDtafybG9ers79mPmg
qA5L5InGWCQUtadMtVslhthnGZD9CncSnZVYJk4oZ9ywmpA+bAVQrJbNJ+EwZh8o
rT78QdSWHJim9C/kKBtl1g202qLgGMOnqwUYWurI5IjLCRRQW8060XmxlRXnZec+
5uekdOkBnDMHaq7SWaqpv+SF86iEe0wOFDUk5EXTcBvyFH2nl8bI3/52UGilG9PE
D82I21LPspJcJ6JM6shQk2nzTL3RNcTgJC5/w3R+koPTLsxle8YWjQwSeQdbJ14h
JkHEx+Ha6K6+TD/tml6rNMtcywGRZkLc25yIJqD1FY84Tns/svhQ6R9HDAyYbyMj
cYe/TGJWnAesWkShtM+Wgl4BZA0Yz/6RpJcvx0UduwfCNF0122VkjLDJu1RqP32X
2Lkd4H2ZYjyPwKekDwlfTjFKOsUmSK5bmzNGKF0QTG1/Sudq+puLrx5s9xzYuGIo
cUHQp+LxkILf1epBctC6MGgyp2XyZtzriwBORTAoWXhBn9rnf3LqttOTXRzvW0LZ
UfpOOh1EeC802qmz0SHcly4L59lR6yJ4KTUVSYzEZrhgqQ61qoyt4MPAGqs07YzU
vKY0eXicSNzyGsJX0jKbQpaE8+i14csyRVVUv1GfVVA4ZlXRp0su7xtszdZy8sjN
kCiTE1hv39TYMwshSKNXT6/35aNCSV5pJOFaiGajDoaHAE7s4kU/ijviUHepiYon
Cldsa+Z4UyRM8ytvJeHGXYlnu8lHQnym6jwgB7McuLjDY6KQsgy7r/z2G2hFsgOM
BuCwk6gIvrALbJ8E6YYDlLNb41AYgtVRW2mL8PnsPfITv9wJL1ld1kc30Vh4Ilbl
XnPaKFSKZyhkHeWaqP1TJX+W1ZWFZ92jhXZvTfPXIU+2G1fjEqe/n4b33z5ajxbs
B5E7SwEifYhdnGzyYRTK0n8L7OU+Hl2P08EQX2VDS6prFBExxB9I8jx9Gov7ozy5
w6jk1scAKwvfOoFCino3qSrmG6Sj9aX8CJB7IpYWu18f5n7RJjzodcCRATsLOJz6
GMPZ2jOWNht7LjWW8QQ3yomdkPx0pcxlOPk2wlbnAD9+9SV21N4Dzmas/aspy34q
J/4LljZA7lN+fEVtT6YKB6qNxrbEYSUA0ICeU/OgoCNsFEpblShLd7zwoUBBsC6R
EroErhRr1LPOagwfQq24qaQF5kSFCEDGPuZZPUL49MXq7PjmJGYK9DqJC+zZV7ER
8qpFn4jdqofx3MLF6zs4kZCWOlo0leUJVN5SEMng4UICJWWm+Bsp/+CGoC5hnU/e
2Xs5QymOcGORN9O5jygNxZ8yTcIq7nI+LKKd6NuoN21rNtkFW3g4tUMThtop1HKJ
dCpTulfPNTcWeyrrmAMq07o6iGZDzohMb2VHII9Qko9CtC/CxjBetdl1o+oONySw
ACNmWKPM2wtQSFGUQcRIiBXq93b2cUDJ5gled0peg5gHDJ9yncL+Wzf7W8B1BE4j
NAf9RnJxlXHJRh8e8FW4Dr619oWlBfcqVXBGnnQhsxkr2GCtQKSW4FZXjkNesYEB
Aer0kzKb2YL4bdHi8bAKoeCmzl/DP0eflFbbTSqtf+LYVYe5oqJ4HPY86lIFTjk8
dYvCfFN9yQ9WDCPP6fAhMIIruIlorcYP76oRO3PTKJZ1iYmmZjmPL6X5AWksu6I3
SN3yiHU/uyM2UBfDFRjrBZ++0x1iHSrss3p1YQv3aPZwZveDbOSwYNk4crFEv8uJ
5hBvAsawdYvvo9ZtKjaXfayvmeWjtEnVhVqltaJp2B9FcG3v3DMxFy5lztf5CiwC
FmpWtJXXIaF3K6CJtTe+ikeVhi6fomEpPKGMT3eNrC/GgfuH3/sGE85sh6Gh8EE6
eWAz23CkaaUhx6EMiDCf4Hjpycu7LP8Eil6m/h+1zwobe55e7M9TnpNczNNNAmPH
wRdwfKC98J5NyzIj8jgTv5DdmabG8pI/lzAyACtJxYaw5aSc7a/xh7tHuDi/j3Pe
TsvJcfsZFLNMTowccH3/+qXMp3QfKoMe3WLyvJ5sv3xqORaWElAxViscwlJCkFez
+glqJ4xFCzycMtFEF5lyslUfsUjRDpCmg9rNuOz5YEO0nQdI/uuub/r9Ml5hW44f
3HS8LNTP/R6/29L1Sj1zPhrlPpfqU/ynOJN74HcpVfig3PEvLjnxXGowQf5Pruzj
ot8LAZr6DY84LB/5/wjZWmEuqfmva8+xJVzk9EQJGMNE5h7xwgABKXr6E/7y3ZvU
6ZBXeU3H7KqeZQdSa96W4ja5wGPBKo0e8mzhVGbqdwAqQflsogaIfvVmT5RU8Ohc
Q9Pvd9S91/VdsNkLdAtt6DCige9zsq2fGF+NO6SfJXulmi9QGYGRUHi/OlaCsndq
RIVyWqZdFEpA/0GA16iYtqIzjIRbWfs2yAFqUOXFLGpZSgRtDZG3UQ0hOnpnFCve
4g7jWlGoSkjUPjHytoxkRRhUqLzDhBxaGZwUh0zNigN5R5EwQAZ/B1PcZXFKL4iD
/ce7uwkI4ZwOB6a7S03U0iw04Drnr8dUUdn07MZSuCUD6E+25vvgagRRBYYZSInP
aQtE5ZaWLP5sbXxgQDxKSXWEXgW8R2ezDpYITj1Pkfu8K6hk8m8TdQ0BobzZfXq1
uP9+izkli7xoTOzSaNLOoTM5lVmrUVDMM6tLiDrc3DUColz/cV3h5gDC+yWsaUhh
61OtDAOpqmj+zDUq0RKYDanYGHX2Odjs/N3+ew3/9WtMd3NRD3M1fK4E5NwnzU1y
cUKog7fAtYxskOM4XJFGhm/f2oG+fjH1msCzVAZeYPVBU3la758iE7zV+KKOjDUg
Vzuz4Qg6RUrNYaDby2ymPfWZVAgl24nY9l2XGEnaCdAI8xM3PaP5ShGSlf8vj2yw
hxI1YSIhswNoSWPw7JdSvpuO1rQZNt5xIm0Dde2nJHvFqdi2Nv2xi7rVYb/K8Ort
FcHTOhdcGQ0jeYeFbxbjNp8xxXUyc/wmhZ3ThuTWMGic9NIDm0JUS+hxSapXzXou
fy11/rDL7a5jHQHSu9U5eQB1HCBLI2Pk0Tz9vdPRnsasFRQnnGQwXCN/v8DvlxUT
EuWjCCbUIKX6Y9M7CGmuLQEDJFXB9p+DnSXqDiuNO9/L0AvRupeGibItF+3NUiv2
+eLStVFa9kKsfcLHwEvE/QMwj5+weZvwxh8jbEmyeUbVyn5Qrr7VI+LmzVbJOp7Z
uRdIRceFVWFKHrJjR4m7eQPqbF+ySgsxPPXsUXJi1dyn0QjiSOclcusP/CjnZNnF
SVAYiUsSmdgEJatvD/fz9ah4zHzWc8D+fl8t60MjdeNDdapeb+Fli1enEFYATkSi
mChsPdLxgETuDLpVnuogVAbUhjjv84b3dqO4Y8ha5qxs1BMZx0rFcw7XHH51Kj65
6wE+tIDh2PwB4iC6B/+8PJf290uBcOsfw1lgJQFt2WyHJ3KoGxoaywKNjSlZv+ui
NY8OH6Y/RoaEFVd73TToMhGsbaIwP92Eq4NpZEDbNlajBPijI2VCthcv7/1iBfQ5
Yin63r+A+wIQZOtugBZlVaK3lBasB1Ib6MPUFk4w3vUeJWCeFKEgJXlBukqXDA9t
Hp5eQ5BaSmJgtD/rjnFEU75wUQFF5ZP/yHTjHP4cYjGtqLsjoSmrkZZvhRs1rlub
FiQIeNEHOYT/jwqrLlNJyMs2jVPasfJJKb9uy4ectfI3tgaybgXY1OPyh8zSM3XF
5//Q+gwR06XKpkVy+FvqsKL6ObgloPk4KX+8HeXxSRVC1RLMMY+fsK78C2eEhTRU
IWdzRxZ16aeJ/FTVRyM08QqLYffem9HH8IN/Z+zs5hk/Zaaxrr85XbROm8lR5EDy
CAeDj21PdW3/fHQ9acfT/RdnYQucgHVskUBcIUsugjNISGoPeGgWqib5f2bMCmlx
uv7+H4/OdY97Wt68wwtbIdzu70MkAz3OQRxLbAaOoMWuD/GVEasjo2E7cj5IisIF
iJ6KQft7T9LYqxz8oaHjv3eqMmrE7J5R0ZI2bV1N7/uY55WmC2RxA7p1VcfZ6hll
r4RV+Jakjz8B2zVdJXa6uYGhzGPjLe6OTiXxY9wpDIOOeVaNG4J8eptJK/ZIgEAI
e6D0EjXEy2iLQu90CbtPE6g3bZaar135xgnhB27Nk7z/Ikjk/gbWd70YIN66BVmq
+EdqKSK1lH9ZCy1dSqBAaEDVb7dKIccJCV0meOwM0H3Wi0ojjKgr2TWXy3n5q7ju
C2FuyTuGk6Ubtce6xUWUdDytHZ0JGiAXxdoVROSmDRj1yg4lchh8I3gJMh/GNju9
xDOclcCRpwpYTvARxXzMx4U0VsDb45KCoq2D79D28/PuV5pD7OWUkvx5/dXK6u8+
YhfdolkLk6DLgqJEs5oVlW0Yau2o03lvHrOgeOJBedRN+wKf7+CDfzdIHzQnZ1yE
Co3J2LwhBZGEoNH7L9VlVOYHeCUCgrxkouy9ExPHEaW2naGrlWyGMCl0cs22nt6r
3k2leM/fq+Km8l9Dg7WvpYDyVd7Opg8ytWPuc4B8EFCqMHTPk7h5BnDF7vQekwGB
b/ZHZw3W1uINoLDj7ET+4ItqmqKyh0RhewVEv5SORj+q1TCkoDtFHaOYIJNX3Tx2
EQTxKgp5QI21uCm5UFMhwBGfzhkNe+MMyorjq66p8V/uAKyaJnKfYUZS9l5foUl7
E3zLWtj5tRtPmDc/NUBy9kT+FwfMFPWh3YpFSoWTonWegpPmHQfYWvpO8D5PhGO+
U1ovNkHNWoxIfrWc+wiFI9XEnNn1TjSou+JxhRDc1uojkjwfeD3l7TJxf0VPKgFd
hlaBQm2fJNZVUtQQKOEG99kXI2VwlPctlGwsMdHIw/3zBChYlLQA/anbsyRfw55B
7zbGkql854LrscsddvFqlN1mqrc+GrBA/fN+Vcl3RQyNMQbUmzYNgLaaummHmfla
s7qwV8+M44XJoU7KbNOjhEn+wSmjKtn9t9z28ab9o528cepcazNiw+UMTeA+Oy2l
DDFL0IXQMlvKhdBqe+a9nrurPoRqL0K9yOd62CPC5YhfrdDcIeCo2oNjUCFTxKk3
Y17uzDDSzakMHnOccR6YZsvIUS26ngzUqL5zs2Yg7zVmhcXX7CX7z4iVqicpG81W
8V51iQ9bp2xGf+WLvjwubElrLRKMd2eOdLl8WPAZcN1lVg5gQy79wgSFRI1kYqeJ
nsoJmzubBmzd3RzteylTtxLN/WJRLqIgeDDFHG69foWcQYlUWN/fXLDFf7tTSynu
ZqkPb3HLqtrit8loN5g2/Lf0TFWrPW7hVc6vvqp5+8w6o/GRrAxHicJA9mLobUyy
Ya2l4RLO+6U1vMfDwpTakb6FJw6vWjlAj7JLKj3xDuaJveJNFJlMsisOJel0SaP/
g5Z9TsuqMnJsO5yNJF3U2CmlGSDZJMQGC+hvltv7x90DEe+MVmcbxheymRYe4Bv2
btP22NpJLhw/4g9tOC0j0ZvjuXeAv9z/CpDXlcpA6PSkUQQGuDQLO6vJonOQGA/f
loJIyIVaXa2BQAC1Hf3TseMWyJD8oDffDGz+S2snRMno52D0fH9WRF3i2rl54iEy
+rwKpmSQ10AEceoWn5oU6JmreGZBdzDCKYq+wMnL5diRQTLjEez4TMwT1dtOtDS7
Vfc7kXsY8BJJ5zRIeD8FSPP0hqJ6bJuhHbzn0bEydArCR9/3p94tZ52ouyaZo3+J
lD6FhJ16bwQfB51Q8H1Q9a29okmGAQHH3dcIY4V52fXlFhhrhe2ORSoenaBZoKZY
6586dsU+XXzalq3u1tnuAsaKPkaRqD3ERyRuNd2yEIq8Xe32kygm5J88Mg4XQvYO
CLcyv8eSUVIc/IgrWwZsqRsOfM6bcRn7Chxx6FEQjQH66sk7DfzmWXd2L+t9soyV
yU9xcT9u5HzWLm7lknCQparpxGVQ2enxY11Hipt7hOYotl1/fiaP3Syw5z3Ot0qH
7kXZWyP3t6sdJ42rYfESFVSy55qnBlr4hA6rkSOmBKmMwlXkhTd+q77pd47P+QYt
aBT3WjLqFNBHGLp7EXjZeSaGKVS5S0CbUYGHktTFlEz6BZnbh/ofA8sPPk9bueKY
cBor1DyjWlefk4SWSmnS6XghbOFNnSDhBeBEofG2X6tl2EmQuaTUOvn4dRazIefn
ofboVm3TA7CCDS4Oq2RRvuNcxnKwS1yrlRriGdH9CDKsPLcPfkFyLpYP6BuUj+Sn
Xsr3oFUBD5ktBby7A1UVEediRin58MttTrHuPy9aLZCrkCwMXiOa+qTfZ13Nl3QG
3PXLY39K7DfN+SKw1eQm8Bn20gy+I9S/mqjjcLYlqqsqlYyihBnvEbTWDEb5yLG9
O//tlyFk6Z8RrSIc0Y18T5ulUVvgXfrZFZWmjJMdzkOfEAK9OJ5qZL/c6Vpt0uEB
N5DeM0hnKAucqKTZosSiqjfpp9Q6rsUo3CKTYhoXUoO+LDDo8dHF41CH01FImWDZ
HfQWhKp/LnOJ/Td2snGkW+546jboGLRhRkv/+XLlZkUIWdXEy1mwkbIEDB8zBL0L
FVhX4aYYGJGWe9HU1KuWT84JfqKNOB8MhWPVoiSMR6FGfS9RrkClhIDrLyy1gSKh
A+pO7UM19Vg15Y3ANCTp+dZzONRON/Ppe78G2r58baSak8Nv3/8EaquImVcE1ow8
rn34ev8Y0WYUgZsELZm+Ldd1gGoh4SabU1ApfL4Knt9GztWXSHb2Ug2CPen9f4dU
/JOZNKGInU/lzjjTCiSZ7uAGBTX+TXQYYf1j/M+EavlA5wqG3xEYeCm+W35qsNyI
4tHesmkIXNZOkR5TzoLRtba1us5an02OmjmWmjrLm9uXFBNCvhtrdIgYvzXd4esb
yIdjnLtLQiTozU33KrWTCPIwxzah/rLaWWEifekA+cXEgefXu3rR77pHz2IqwaqY
IWm2PsSRp3BNHBPd7XDTIa3uSUwC3FxIOqY3JujcO4wYuN9khLndmO1QiziDZZqi
u9NrrB3gI6jeF0xtysbQGS8J5SpzCIPhTHfv+YNlRd2Yq/ipIZyKhth5YavMErKH
/6n+Yy9z8noZPE59+DKgzhjhFI1FQRYGDVgHH32zQU6SFEaCyP+8dEFjhud/k8MX
A3Vv1yMhIX9xRNUHMDmjxO+gT2aN5dbGBV+Rf0dE8RJcKXTIwHI0QLoGzf9Y3UPz
Ydfo4xKgIe0XpG3zz+4bjoZ7dsenGGONJtA/sLzsKMWCUSh4ET/bCNVkoK3s19bf
DGbI3hWKY4eBd+9HB7H1MuHlQdwKKHO7xiyYtjIs3uNGqskMi7LplNtnm5fDokpi
SxJavMbNd+BBvJVEqMPB42cHCii1zgg9r0L6mpg3Ywdzm0hQSNb7mRIwP170gyBS
YUgrrwEJAAervzFVwjJIXXXDdl6/SlmFI7aRkX4kljSlE+Hp7j2o9odK9x2QDUf6
QYYrh9Nl7T7PMT/pF7/Hx1i7xUaR5aO3S7iJwFwsw17GS36wAR9SguLV3vmGaIBj
9PMLR46es2B6/sgcuGl0GkjyIb4UpXaz9/3enL3uOiJz44s4Y1+B9OMbbaIPug4K
RqhsO9dg6ZAnN+iNjjz2kQCeKvo1E68Hcl2KI8NSflNU6VSJ/nbypTtF4/oP33QZ
8MZ8W2/nLIBvU+F80VLvzKOlLujsUmeTjMjp8TQ3nYyLILSeMjqU0AhrloFHCpMy
8QMMB8icS6PCWlWPAJntwekK9Y9gXddVtq4AqSpuI1A7VOBp6ysCJmyOpalEN0M5
At36pvjQTMCVSgwrp8fX0KZwRt7XQPFPYAvCEHhK5YwxR4JZrPCsxO1sWItbRKS1
VNk50BHIxtQN/afGlUbaT3ZzEtNwR3pnGYpmp6aiAtSZjZGpfTcB2PbJlxo3r5SK
v/uEofza5dbGpmhRmzw1wVz7xMMN+6W0k1ufAzKe9fMvmogVPj9xWxYhy4/ltvjB
+r0YFzSICvROwPrg6/qlJ7Pg6jQaQPFNUU9Gnji+jO8uJ4dXstvPMWVIa0r63VXY
qBg264Fvyvd3DhxMLx4tX0BhqXoVhFIXRZdMzmXcAB5Af01IKVEKidDaoKkA8zK1
gLzSGLuDphv/9Uxu5PPliKuSNwmlSyLfsr7sPpcSbKl3fYJGSmdDjIY4yWwXBWg+
kxgNQ3l+z4l7G6McJ1EC2N17yCYWbkwjfs5INz/i0R876bQx7IsD7kgZSUMSZFg3
CUkX99xG8wEtq78YyETu+QKeihT3t2oigDalgTqduLWwpdt4ncLzO8Eix4YAsWjw
/SdR/bhL8d37gTkxneiz5oEKRnDpXrMf8CjdWc6JcNt4U53m7gnun7N/TOImav/p
xdpJaMPBXAGzjMMJUF+6SRo9kmG/t1CsTz401YudJt6o5dRVJe/GKb43//4/iTXM
D0ymvpDISlSnSMz7wGC5+t/aDT3W2xJivBzcptUd/cLDJeDoYPDFefRxofytVqLn
EnkGzr/VTPU+HMIJhBC1vk5gFx2fsgCLpGDN8o3RW1uzYcfXn3q9jhpU/W0q8UUm
X5MJiZHgUvuJtUTr61Fxwj6H9hf3eG9dr4qO/y5oIGuBHA+HvhAtis4QYI1IIVsP
tb2Q3Y/i6XFIP3+EPvSsA6r/CsY3+WY/RyMFKf8wUDyVt7NnELh7HbHMcLfJhqNf
psE2LefKO+ILiYdJ27xX3erA/ydfiVPH/EcPkPVPV4EX9HiHJ0Zg89nPXsg3IQNa
KQyva1iJSs5NTBWakMYv5oErfLOAhAiUENydQip8REMubViRksSUqS19gNlmeZYu
sggPEXOJ6NE0+tPZvbREAMpdgSz4CDS1BAojtmNIqAMDrHwDWJF+Vl5Xu7WpWIWj
x6d8c/xplGbSL3n7soxS7rqhZx8gk/SEXLNrh3WEe3o/2YsSNl/utUSoN7v4wUKM
tvhO8cashGtmKwHIVCNLLo0pz8DoWhrT6wcpvOUk9pEiYapPeoJF7QR60Jw5OPZr
VQEwQUMryFJ18L5rkbMZwxhHMOJPdJZ1JMOdI+UNKny4nu6MFkGiP7aUHAxeXF1X
JDGfF/8hSOiaDlj9r4/dzIDZisacm3ZJ5C8I2QhcUhQ1hXtBKfiFUrshfK/lCi93
UFL7ms9NZgFzQQHwQy3yDokJB4Y1dbqJB0dxa8a9kpmGAf2DQcJFdLde61t0ncMG
/+3wePS5Jz06Yq1eZF6bZxSLr4y0wiRyYMtKcXplv5nMnMsZlL5KnLdEydHoQqyD
Is9zHlcRdkiPIcJXdW8o9s4f6RYXrV3RC0+WUZPYxhY9d80n1Nt0h4mdB0rCChaa
YIX2OjkXaN84cjm5EBSbcFmOy4zvW152LdJlfT8SBptREBWrSmjA3FzB1ZLuET+m
bWhX4/UJWQ7b7p/DFfuULiMN/pn1TvfYc3F3zg8QHWajMZKsO+brFriQpRYaZhr7
IKG2l7tyszj1V5bTrdk8ntOwB9a7dOYweDPa+vGoa6I1iigWOrkUepacB//R0Oan
0Bq2YzuIXauhvXfBnBAq/atCMrc7ZrMGwWxd0/5ERnfAPFOtdctWSKPfuSGmjGR3
zAZndK6oLv94sBwKTjmHxVZpbR9vkBmpCtYpXqOAbRh/VBkDfxsabpH+Agrv64B4
z4cYHNYRfW07ujQ1T0q82pVwhgoiqUMwf6PsjyBPVhdt6hpaLVFSOQ8Qf+uJrjuc
XMvmXpNCwQmP4/zDcr3SYNZ7a00ZtRrLdtfsViLbbJKaDAzMBkHCmZ3teLgXfdfe
vKlPbos08FBAAyQjadqypyN0U/qPFnvJE6nBO5imt6kl8STbv1eV4uq7NBCP2aLj
OlPaVndveI1AgxOliY8vmV4W9hiMSnOnktK3ekPeGAOgIB3kXJIxPUhUP7wIZB4e
7vkrEyrUg8ODuPtNB5qB1hOTmb3Nbz/8n5j0aOwc/x3XS8X9vrvKtIGZL7lkMX0e
vgPDqfQq9IhaWL0Rn1lfyk8QOFWC1Z1bxJKGo+k0Xxkq9NCefPeN7f9N6LwtzOft
42DY0/nrGzA+zywRDJspia8RkH76m3OZbL2m4EQrNjbb2+bqNDkS78K0XDxhf1SR
EJrKsmynk/UAWZEiLCLNqbJsD/9gVRwG0z114GKFP/YIWKyQQM3jMZcORud+Dnjn
RN0Y9ewhR1nldDG1pCdcA1ITSvhPPwCnVmLjBm/v26crkvE2GdS00mz3CICnVxdF
mALUkmEwmDmM4RiGwdtDUpGIRbY6BXzvAWCLB89lrO/3qWINWAEMCyIhZ8J8WrIz
zACvCine1cfnWcx6g8UPgP9iZYb+afyX93pZ4VSrVclo8oKlKS7rkCcpA2ZUW22c
rdE2/M+NRQw61UadAHkEwJFRX9ps+RwnyzZGUKZXKkyjQ0uvS4YBawH3LAgGvpBz
6vd+z12E1t9Qe6mKegZrJi8+Rf33F2QquQEM43sFQVU3phQPwc4ulFUESDpJsEa2
n4KdZgSPkxVR1VVEcRZyhDJ9z/LDUolaqzEC/qeqA2ThaKJBV2kCMSvvrF9y+UHd
/TkR/o6sS6REJAWuhJ8m7ID+kNrE3s6jQ7OqzMLVuNPyRqax2V85B4UpCXmxGzCp
BO3YGpI35Rf2emuyxfmchojqmYxClbSijMwQlJteKMNrF024DXYy9wrMUispduOU
7nQc1nnRmXaopLYhWTXMj4tMxTLcd11hMkCWQTmzTTeKV9dvJICu7rVARH2DgbWG
zLPqIArfNOU6VxqmtjYfJ9QNzeXcRE1XHbJIo9/8e5nXePBImI4dMKCkRmIEVNwh
zLu6w2ON71Gx3f0C9chU+shl7Vi55G0etg7ZYtppQJ8WCUvgXtnzJfE+dd3nvhuE
fmK9svH3Z0mxdFd4Jg6a8mJ58lx8z1MNdAyjTtKl/1IlzQuNH27rGZMVT7tb0KJP
d0ExIQwFN08imxIIPNEtgc5PkHlD2BI3GGgDbOftLMv8Qd/vHhbgnklODPF59YY1
ym6l6S+M/zRy/DQLgECNcTniClu2LRMZ9nmatOx18vr4TiGnTjcN5hoCVvFOOEst
r60/CykuET9qx+pPSK8kRqPpy/qca8wyRVCXbO7Uo1ZbMx7oU6jo8ZmEZsFQEhnX
7SYhMuZnoccejtA8bJhyGk5BEwN6nSGyqn90P/W24xbhpl8S5I/CnHgqHOzIfUKS
A7BIIIj+dH1WR7hiB36GV+qjG+ZJqKHGS+hYqQboosdCfujiXoj4JGvL48vDpKPq
KiyilPYnQ+dVrcqPmlZD5fy2YaB0mtDQ49PvGQELqOpZkLogjJWfhu/MfF2oCD3P
qHSlOztWa4RxYIKsi6AZHu4FSg1NSZWAH06OmgkJmWAzQc9nT9Ts6+YeQ3GOFFgI
MB7ISaD2lI2ht10EbzGOQQq5G0PL8acCn7+iBqRcdS2/WPj8HIpd2uN2RSowTnm6
MM1yTFk68vHocweEdecPSEYuiWIoOMhoTnS+sX/obzcq6WRPPudD5BLIQnrvVPGb
0K0jhy6DuYWbnblnsYBiW3CBcT6F0D4477tEiUl3597/AGXpkuh2XNnqVBgy2amY
u8KDP7iy7gmj/KilETflXf0EmvB+lBLvbxq0QHw1cDgkcZK4g4aj3LmDPJY7zsRM
eGYuaI3g2Ns0+5H6LPT9t2wdqcV/ydyx6/p6tSXtElLkdrgdHgiETj7ZJRoOxFm0
W8I1tfNuAWYkX2H5vDffHOmPvaHQa1Fb4yOl/b8rQOiJCRHd0fOwkTfaTEfoye2G
10wZZJadvyY0rcgacflZ1XARmZxWpmH5xvanNgljB3yLVfj3gs3vkavXl/PBfN0b
FW23F/+z/2xBajCuMeh8kP+HMMk4xGl84GYgJ1b0sDgP/bpQU/XJZjq+7HFRmoCz
SdIE1JUeg0SlhEZ0iw/lxvWT3Ojl9YDBBcK7Fj1kVZMwSvEKbh4KHpDqoNesT5VL
o3LsfBtx2OdEWGye6Nu1GbdNxt35cC4NCg9ENVhHJvgR32nacvENpyAG7idcYaG7
ad9B3Vqdjjwqqgae8MXjijNKLm71B7RtGLXOItLqxk23d06nKiAySPo9p5/NAaC7
hPerBWWPqqr5qVIPpxVbhft1pIgjfz5WMyNinrd1FXVj20NVTzFO5b0zlmIfcA2J
JHxPnGaV5CS9gOjP6FFgvlRhOPGv4Dmr6F13Lg/JY7brzUE14Iheqm24Va6Lqq4A
L761RtJohBgmQEbQrq7wCOB11bicgHoSMSvWj/FiY0Cq+RrmcYRDqCxoqjygPVxi
xEWADzGLeFuCf9UbFCig+08dnwnGJWbKvDhfYc+gLItslDvLoefJ/yromv73v42I
x8QWf43bISuNzNZxzQrvzKtUoSl0rAsPd0MistxHGfj3MedrbbdPV1XJgIuEZ5Xf
dtulX5nn/8vIrWwTCzy4MY+mb25yEIVdH/MzrzWRFc6MEBSFY4oclGYjzJjB4Cs9
n6ubKfjajS09Fd1lYK68qJWHRFcMl075jiJ0YozXxDGqs7IFJ/Dc1Nl9UWpc15nR
Q4CBeSl+Ar4OkAkWYzmwSs0NMkbEyIrB54FijgMGx0jsR+qjc83szRYg8uBRDMBn
me8fVucv6CCHmOb5VtzG4jf+lmNwi0EwPqsHh+0lFP4Ll/R5GObNWVdIXmOCscol
W3qAMEadg9NRfs1/sqdzCZBL3vz+G3WGp8ZrmFir/J7gxL+sZ6YmebKTIyQspgtl
RMHarRmJK/+8h3AWEotbsZEfqt6147F1dN/Mk6ixP49omgKManLLF0m+E0QZooIe
eS2vdMPYhDxIQeeac7og2cHRrxhUXepdVR2JZ8pMlix19f7d2PJnDH/M+0wZiZUB
MBRr4VWuNF067z7cKULBty/hBPuPfhelEQ54lPiBGXfkv6iqNmjIc9xMUJ2q8GdF
Ab5YXrF8JsUNEKXCbS5erQCddVYZFoYfOO/v8b/dsSNvSVd9pzuPPhyZJp2DWZLM
CBcbs3AC0ovTvujgkB+VgzLezSO4skNyfYPzTCNtktcK8nB3jInP8LmOxFaSRdjS
Y85MsW0WU3WKnCv2FXcmtqr9yNekswm4HynMDf0U1shnh16XNBnX/XmMrcHaPbAJ
4FRdnF6J/sas3/ohCbXdR8pMJzgEPIsu9voBz42zb90yq5k2Q+YvWj0wxG1vSoTp
D8ZofHdBcTD1U+RM6T0ozwjlp/5XMSd6ceGL5e0fzHnqYbhMqHaDmZUL88GaVtL7
aHRYR6YsLOsus8nxuVyW59Yw/jGn5fCqd+00dII5QmUDl8uWG7uFQ9IdBe6sLYg3
lnYJ52AwkI2o3sUG8jcstsXYvqXVCq/1o+RXdufYoyX3psVlBfxbhVXjCr3yLCv8
F5mkoiEWHGz79UdtK8lR/DJV28mP1NtRQrlSXvAMpYdIqguqXbkaZ76n6aLzpjOH
z3wOB2ZkWUJ3vW3Bu4Bm1VM3wANLhd1lTokTpLigKKR6QnByQ9kWlF69wPy7V5wO
8w7YN495XPxtaJB5bPGbtuzLUtbXqramDJo7TlBMGePZt5e3vDQG4ENLB+hk3o62
yLD1xMsAJ8GMa/9IvABKBgwGYWEMbvrc5fJFCC7gSLLoh7g/4Cvnuqc1NcM+PkKH
vpp4fzZzmxs1TU6oBqJxZQYz/QW4yoRcrFUocn7xOo/MesrdwBXCehmGMhnA0sbV
ttMqd4dETE5KEBcCLfpn8kSmXC4KvD8/Xu/2R/Jago/CnIGKQjMhK77JhH5jwJnm
5jNGetwyRPM0JoxlG8xJZii4u3hKbKF8gSVMK15CzPUW3iSIFeGmMAUjnqJ1U5wf
M0HAygH/nEdf4j5ZGD2iEli8Z8epG5kHBe8fStkZYZC+cziC+yRQmS+ZzjQetdkP
gMZunLKO+kb8ve0VptFe1ALncfXKPhRZfnPqxOaGs5BI8x1RQ4b3oe+4XIcYXtbs
9QZAESF6wMBMT3vEUUS8eDON0fWeWAviNZp5hsGoN3hBfhNf1V6fmDaUhJDEXlFK
sWyUt7AOhMIdLN5aLfKDtMeUC64LF+QGFxU/scLBn4gFujt6jbcPM6MGIT5J7wSJ
glLPmCly4QmvcB2GdEJg//0i1gX8w1SGBNvEtwYJdUn10XmVXGnf5s4aV5z+Xyr6
+gCy22btgkU/47Kh9XXFZ5IKywn41aL/sw5A7nCXl7VQwteq5Tf0rXdt7utEiP1E
g/T2BE7/a0jk998WY5OPKVtznbjdMnya35oKCGEtjs1dCmaBrLpm5/vjvbzbYGab
GVD4DuLVRgaZbVXOmR2rihCYEsKheo1U2LuYFrCr4ZrPHi3UGgzH+9PV3pijMoXs
+Js+l+HI5ssZw4rRjt0NFLe++ag379SQW1LImliXRrdQJN+i4jVO6ckUUWiuxNqT
InYbPdJ89WmU98MfmkWls3RqVB9W3IcQwg17KFpGxITy8ynZH2X9cvXKmrC41+fo
rWoRFCH6509ATaa5NIWa1AYJ4Ns6MUKN7Ttx0Dm8IZt1IxpgClJQjw1SozVuyCvI
Jsj/5vZfvFSCdlboyp5yXkUcbcVpFxmMMBy2YTyM7WU3QRSYu1YeXDyfcFl05COj
7N7d5Q7QWvemeC1fGOTok3jOrdh17RHbbFNsA1eT2di1wgN7JFNPMv8wTY40NHRo
hiAkIpGi7EIjLrWzRVzzMO9Q+OM1CmEMy4OiL9tQ3YEoaUuB4P07d09OsnA1zWyL
dXhi6ngvAwAajpsWEdUtup7aNw+4LOQdGbZlxROJI9RlPt4CdBjGHsFqNUy17+cP
oSeQhcCLtq1A2h7F6eEAtzs6bH9KSTiUz07oqoRH6Fcq3/3jKZdUvQ3HGygAHG/i
IYXWEDpAtGWVhYWWMbvsP5Q42e+A/w2D6gtlCmcLbXaxsBzORK1nmg7R3vWIJEfu
B1Doxr7RK+EDTiNvj5vZJmG4qnqQVm0AuTs1NNdW14kmVORePX2yAUaxW2BrzhIZ
ioZbLoeTgtJS9XGjOKiWP/l63kPm/6u/FTONYWMSgDIXktlgzq3IQFPPiBPfPlq9
BFY1DtBSl8LIfr8Gj1E5gyIqPmvDgPzmYvnpnOaYf+ieUnWFe3rOXnkjZ+vltkue
21dRnGXd0H9zG9V3XMn1HgoXabPLmCR/twdcPZPBz7vO7QWlQlosaUuPgKESVl6G
t5ytbV5LLBn/1yiSBoVbq6S1I5BjbrAR7yvqyMQrxRzpbJxBOQ9qpaPrtBH5jZ/o
OwbOSLcKvThpdis94Q0TdcFt/g0Njgv60TUuLxJMHaYNkOfC/Nnp7XhbwY6gOmlr
QTV88zDMUoCxhsOEPII4L2lElyEirDFJ47yEC+GSeXEObAl8mmQv5/bMn+v3p+by
PDQ10PBlFbKyHpKDue2CrNPgwbw6XW5a1W5CxFvnvOw9EkNL8/nLIRb3osIgtBML
CxDyvjiGoH4VJDDru29FhWCNqihmWKYxREPikbJwLWumd4bNLcEJ+4QKu30uIgMG
B4yY06PftXAZkOiXA+P+6yg3cRpYjjBs5JMqlyc42Qs64Nqiel3D0rZTeVt3HmNR
GqLx9GFXOiVUuCWJxQmtkU+Fcdc4JYye47HVhCjWo93HCJvUn7IeJ6qO/lhXuMBq
95VsvFJj9XFAbZN3p2gKp8f39vrjvn0Azdx+jRFKMjLteHXDIyh7IDPvwYULyjO+
anJ+lY470L6ioutKyWOev1Ls4wZ9NPEYp0d7srEbYZwv7DTifKI+ow0knp4stpxf
ZXuOn4pZMzZUDsRxUw1CY247M0porgyFmyd5zGBTKRYUtFgyG0W6lfWmjbbDSgpk
Wv1QoM5C31uJXeB6urT+ScgNhvMpWfQ0M4CqDGE6DjmUz36n8AtNQ3VDvjUgVzY8
ZyxdY798JlXy+GXv2nNJMiyr9iJeNfPGalya5CIIs9UdDoP+HlSW5SFFsJmth5Lu
zehQTHDp1pfwMHLnlx4Rj6SjAO+UJ8+ztS+r34Jxao2WVkkBiY0Z4yT47b0WhaCq
/1ZJCsE05Ejk44OBMjshxL5OvoJoiUmwfdkwwFZCRuw5mTE2urITg0YviOns447L
jPbi0TK5zZSGqKZATMSxhb/2tjaCLMJp8WHQ20e5PFheyoGF2YZjZAsphQAPNdg3
P0oRB1aHPLja06lkXTK+kUFNiF20BiZNEYaotrQn0ZfbMoh1gh8EOREEgiWRGfms
4+PLqrM/kRE39yoja0E8YYVbH+RyrLEdy/KBGGn81GWoFj8BAIH9B252JrI5dCNO
X1cWOj1HYqFDV6fJGvXxed8zYjXFcrn73rH2jyIqQHZnYv0pm6V7RjYCw0iAmQAk
Y6+hiJ1OG4MVzeDrpdW/s168GuqrkaMo0AX65bd4HXbzYl4NOTG3Q6TY42SEjITw
z/XFxn2I4eBeq994rP9as7SJ6LNBCRqzHyhdKV9hLtbx3ONuZPPTF44foQh0+Ev4
6Q3/2WslYMzreBK4ivvx2mon3dqBsYs1/NngyCS96xSF/abfBct+B7ssTS0XbIEF
wPXwBCrl/8nTpO5h+VzqKWG2FVfeoez1bBSqzh+FDjHdj9Em2XP8MClVJVRwmXU/
D+bcyZUPydIbd4Rmw0y3YbBvh3EUKC0lJ90Dq7oSxbH5FLbELsEFi4aa3K74T6d4
El9eZaxlwJ1kVsrBm5Czr2hQaQWC3Aezjtr5jh+gGE4DWdK/0lIIueLGot/+8Auo
F6pQnQibM4E6UWSteoywLktQYsa8hwDH/zC0u1rNGLXAoApD0N2lvFLZARExd7FN
IcfASleltn542AiX/COzvcF5h+dqWS5D/EsOx8g+i3YN8X874DT1Ghnkd/5BuHT5
4wPxQMTZezxtxUjt/Yvjrei8e65w2f946TCrC90ivtOXfuA69aDfj7qFK9SD8O4W
PAyL+3xYT2q5u8EEc3Bs1SYo2ONuHNkwrYVTyyhKbOI44B43mVNkxR49u6G36ToC
4J4Ejoy09TM5lqSsV6B/d2gAZ6f+UDQrIZKiZ7vsGdtu/wWGLyvelgiyi3jz17VP
mM12YZaqpSlVGH4MKvYR02FQIehhJfR/jl9odb2tQxerNVNYqB4fTlz1xzSSS1hA
jR78eth51QoVv+bhv4Vavz1f6TmBEgQEtIBZZeciaoa0wdHKOA7EW8kmxrdkIKk3
LvyyW0zFctOTMjZm0MZ77NFXP95l1Idm4JMjvPxVd72Qwz/ZMfAKJSPPMvoQ4YU0
4nJCwtiJx+puv1953a9WTJ/c7TxGh8Bm5C07/65QjJdqqqnhHjJXgI/fUyyhZhgY
slETg56UdqOvR4ueZ42AVAwbqlXiGGtyX68eA0xJgvtQEvuEvvyI2JFvsUp9zapO
PmwrDynUsIf43JhGR/dymrTFMRVRNUTEdKOvxmuomACpLEKklORJRBEfvFehZcLI
9AZJp8EF8ZP4thxKmbb29+6jndPtrJD/WNUHYR3E+GcxDqa2unoA9xb9sOkf4ZLo
BN9fw7gPjd9NfQf/00YQIwtLPL0+b5qKSJltZ1ybghdvaxw6h1+PPbPFFfrPK4m8
Lqh+AlOVAdU9AaaRw+O9hzWPon4gPZq3eeG9wDZfI77H+tN010gdtYdEjKlDJKYS
tKU2DcmM+bbINidnI3duenRMUYEzExLqoZ3Qv9PhJ79Kwh4Rcrko2nhDt5SZwPIb
UOldphxxzvMr6p0qbU8ZKLVeEoFSRAkT9ty9aEhZliFWF1lsa+Fzgch0nRA41t9u
/qseM51odAVBf7OcWLf0rhCLzQzbOm3mZnGj6+7lpA6CJVRH1g8MY1V4sEtS66nm
L6NWykIkWYw9A9m/yhK+rf41rLno7dyEOD4Rl1wS3vzc+TGeiy2rsXKc59tm+1eq
5bh7jvrQwBEVoC7VwgUsvGJqUyIiF2WpDPD3O5ZoRP4cmMrOpkffdR1BHz8VXPhn
8rYY2ZcC9PUyX73qpmogjuytHBygszm0sGPyTmXfsbHMK85TWr/ffukIPxNMJck7
gXHOsRB88TFMTMPXG19RJRoXX8g44lJ4jNyEkTTNbkyH3KJ/l5anrAaXCWekQj01
gpf2sMMZGX122xM548yNvZs8xQ8n13nDEnTdy5U2/MFSjnu7NKbov8R75aUc3L+u
EqrXm6Rffu7xgemNkBEw6/qXF2CeEVJZhHiOV9FHwolRAqZ/Wcv1CgvWH2Ya1qu0
WGp28Eg4uwN2KuHZe3mwAwfXdrKmd0ailTZJLqeijRshETcGMdtSkcXyyrJ43CuN
/WepBbYGTCafZtqVBSLuMXm/iN5yMnVo8be9BTKVGzclhhzIiv+u4HxnNFwI2KwA
/K6/lJ6av37++uqZRoUVc1lF9tH4gDy6Zrl2UqB0jGeOEmd7kQ0keMWrCh250Kxi
n8/c03b9FTNKD7plL99nlBA1N7TBOH8DJNjH3NWlfAWTRamCq4kWBtzLHR9bFf9j
7CtizeSTORueYbsaNjsCuBCIBFWh5y2dCWr8nakykfdkpBiX31iH/hgQ+yrYjIrF
iAyJrd6z8q6yCjvZehdcrkRUWxP1vrwbW1O/g8NWGTHNNNaldm1dMRLZv1Kn4aPS
3g0SQq2bcDA5SxWHeufHT/57lcCIA4C5ASKNBKL9x9weoP1qr74a1sxSOKK30gue
dGXlpgHhIRGlASl0LeqdQyEMSqeqX0RBG4u/33JzyACuJiBXRQQiAehm+twUp7Vc
7+0oKEl6AOswqPy0vTRxAfo0xTNRwNU76zXF9UaeV8fu1z9m5hcQ+q0SDzzKbhnq
LL0CljrS+ATLapbb2w/PNcsmapQ9p5ejOtg1TwNopqZZEbJIZguSSqXtZsTgw0yt
qzuo3fmpDWppcTaIUJXP2exsGFGZ7Og4zn4FYxc/zN6mcU7v8dXltGWvN392e1Vo
q2kR2j64MToUbDnvQmeuSowOfUrhIbFGJXGHET17FiyFfEeifKHfA5+78Td12tYm
xE+ZWAot3KYOUxGDQC9pUqLg/0QiEOWL8ONJAXypfEm5w2wpVO1iOvzsyH7LUW9j
Csu6UmuumeacVlqwjZlDAa1RNn5E06gZ6VCJGONL8Ed6WF9MlOY2iAhIq+3Ww3s3
95uOqt6AIj8jGePb+QDqby7JBBFuvtYcDpkqS2uHOYcfClDgUBMvEobeRmNiNjn8
TERmHRx7Dxsx6OWd4/FsOUoECtiKAw5MOvOx63fCp9VvXJYbsxJdfkXCgakzLkvO
5lMj1lDq1LmuPrk2FlJD3Ek10YifUTHN3wyWX+i/L9pXQk6vz7mI/vs/Q7TMEzcw
RbwtyoiEsw2UJnQOV3k4swBEc8OAsqrYXioJ1Re6FREFi2CS4z62lPuaiX7acEmZ
m6l8droIFkizfH5YyU4AWg7cmJAH5CQOWfzYYbvFB7CGmJbfIl6aGS4Z6jP32YWI
duPkJf1XsjqiB7TZneczxQAQeGgGT6Py8FqWddz4W0rZF/OPiZmYEKaqFhXHEHZq
sBeTeGimgakNjtUFe8oCRBWnqr/BJaLKaUVXq9ur5sLc1UQS7Rgk3Bbj1UQzjJXw
AQdXlfmbG5BFLO1Ptq8zgGPU/f1XFDlMjAaJodcqcjuL2wI6uWK/IVoSdXZtpqGB
gmoOk8oXuTGv8z4IVElrO6vrjpEhp0TLSVXQa8AJvFLu2EDX6U+Ww541ghrzX2c2
Y4CziqhN1D3v5XlEbp2D7l3OtYzKmkb+ahgO572M1GJWWhpfjtg74SuKJpKHnW9/
sLwchkIlivJJ+JYZoD30laMywokhw4u9h+DHAIrEOkZcONjdTt0mI2fDdxV5927O
xxyfkSaRb7cv8m01oHEUttt6XXXBYHGQ28lACYVe9LclmV0g0VvBVg25fpAwTHRM
MOnvX9J2ImVKzSjku5v2Xzs6JrJ0LupnMxBzuxz6+G8tEfeq8BRcez4SXsvr26Wy
IGQL0Ez7lOmWwa4Lmnd9PUQsfH9XQiwxXYTag7cHDzr6FbTuOSOdH/jGS201eiMz
nz2HppjHjPj9uwsctXRKWhUF1UQ0rsAdlZ0Ta05ojdqwrYWeD4ofAFlIkAnh1bPK
8aWtspFpSysfoMZf3yVpUmxZ0Yk35SN4oNosuH97UZMiyChuhRnXk5yDY9lI5lg3
t6XA49Y+uRaLZsvz9M+lUsQJyMhzGSvcB03xBNVKhZZKUNe1NVYYIIrCPRKewTOc
MJ8SCtZt5nOzz25YWc3ipnfdxAlWPkqQ1qnhpmb7AQ5CRLKCUB1AEVgqVU7ALEqY
TQAH4m2KqeATsJMCxuyJmZZWjv5RQRkQE+tdV1YHYPpaPYPxCsoak1WB/a2QqVGR
pv30egkO4SuWCa+T42EPXhQE+Z6kd84Ng7AQjJYAaFfJiScGpY9VJZBrNkuKz9ql
+KdSgL4Z1Y22Oe6vp7fGR866MYE9gIqml1ndYkbgKeuC+3i8U2L22DWQZoYwZdIp
ocAsfnMoPp3gLxE7+kgbru+VuIXJ/zGhI1a8MRIhGehpiEkTM3j0TxlxwLosjkuL
J+T33ep0lZUMASctflh51LFJ65Y/nx/8YPJvP3prW37IUuHS3suBjn78rG4WXfQB
uUK5rZvwjl/WJnWJnvDxm8Z1wCrvQQd2dcX5mkBXKTUejvfXH9Tn5KYDdKiMcaSO
wponRFSehfqtB43I6cEDXWcPSG9VWWUveP873LzfsJdpYlJzcQrTjoPFBVu2hpKY
E8xMVoxulfpRm2KD2HqOg6h7cgDR2N4Jz2AE2km75dSDTxmHYP6dcktR03mkZSIP
tAqarlUPcyytbQWfrCTO3urDTMAluxmaN3svWlySXFiMd4HFJJ2rNSPeNamujM/l
iC4uGQLU69TnefSnM2x5XE3R28AtGaN7NxvagKWEw77UTORxqEJ9emCpRxhaZLEz
kXM9j7vVKYcMIuRHXD1ZrwIdxcN0LBhcK8nJ/djn9HVLS/Y8yWiw5AVk9yW6xkO6
ee3T4Sjx5T5P0Mu+tU7pHMlcEAYOXUi+bLoaSn055Brb56GVPt73UfTFRkMnXEh/
aKZsesRpfIXiFogd2OihRZ0DWaz2eLHOgiwSZKhLvFGSMAsknGKhpTR26lhC/7n+
jvMHWVrcYK6L9+GK+/60Kt50HxUsliJWypptRWT+MXQsidyXryIrjBpaZiU88Fvb
MW4Q4IvbebEGe06mDIM4HMrHb1OMODmHrjgxzi1cKibgKhFDO/IY9iuUWCh1A8Xx
WA7+JWLaqjbXrWhPMAtuo2zjjs+Ly5QhK2NuQGULovbcC0TysgnBbqOECtlZAd79
gMy2W5hgaXlduNhnbDuDtiXvjOdrteVsTwtBf945AQ7OeLWk5xxxACJaLgMcpmQ4
yBSck1G6di+PsicF5FpOA3mOmHGscANtm3fGBTXSGiUr8+bCYbw6U4CPwkeafXtg
TtZF048K76YSeOEGJeu07wzhcLICetBiiMtPs9FDr5MPTQikdgjjBd4eibK4BwUn
yQi75zdynNP9PM3PP9iMbI+Pqs/o2FoKZf0xGg1j3hV9G6ydA3G7w70ZWY6h76jK
ADdeAAyHZuFtQ+c0an1+RLJodJS//20MyOAOrY/pxHgO4wI4r82XlK8JK/61YO/Y
M11YXm8kI3HDF5GfIHVlzYYS76w/HatnG9EqpwMxmcWFx0JfyM5Q5jf7Mxs6eDOv
/d4o/CoD4GsJgk5LeZSqqATZkkq+geu2XmwbXkLO8xk/jFlw3C30+B9LL96rtUFB
tHQIAIhce8vqmbbvh4tbzIV+/z9l6E6iSeOOoQ9QZzxeW/yRs6K7CanIdaBL2Xw8
xs+x3GKEctt+zhkueT1I73FnbWHXoanz5YjVS2klzS2RLtQ20vt9XobiUjfQIAns
pbLSsx9zjpVky8qOO326zD7ue8/mXnDRA7j6COF3/13dKqpzca2jUEqVnnXKXAsT
Usls2Gl8cuF4NqNBdzmASeYyWS/GpJctzeMX1yDgatYx4vFsXkAka2I0uDzxT62K
lXXDvB0AuHnVDe3FGSgCJ2vOv+Wrup4d9RtMrjxOtMmzIYb3L1ezbjODyvt4aRBU
QCo6PUSQS4Wowj09nYelK4w7F2iyHvW+kGkYs7HCPcsPUl3upsuYo6ZYurY/ctAS
lvzvFazBdjSyfiaW2rYbXW1eqALiMobh45JYOky4hk8ULzensBrz75uaXR4QbUvF
7da39kGCA8YB8tOEbROlQEK4+2h5IEkG5g0zzu+wjjbZjbJue5ExpbkPFiOAc87r
On/yOOP+7L2SmpER4TORi1WLPWGYqhK0i9doeOGOD79H9oklJAoy4Nj5Hlv03WG1
ocyTqGGSQHcGQk0OTror7aphqH6uzoDq7u68LTzciiTSM63dNnsyEOv0CaZE+4QS
QnpsOOLh25uRTmQgmj4FmTJODfdR9Dl5/McikB6LfdZzVzF00urh48+8sFU3vfj6
g9lxJSfIQmSJe3bgLBCIeImlcfBtj+VXw96U9WeqkgXvXCPuHI3T+gHr0KlG+w+e
wzSBYW5GcFQn+ub6yf9dMiHH4LpPqR4eLZUxwcrtF3t4z5K65XWZrEjG9ovE1a8H
9ZEtOdRtwAl6nnDCerobXo3Z2WoysNUs5KlMMgakOwBJvx8nLBEyNh4kRaG65nf2
ls8+PU4rBoDo7aIewqg7L16l/qYqaNKseYgNw0qIs2HZzzJxkJzCE+ZBvbkTmrsd
d/ddy6SoUZCsR/rRXSZKiTI5qriVn8lLA+ip+jMm4R3kAuT0nx5W79nbL+6nwSgP
zul0RTRvrXYtHQcApYS2q3mZLVf9WgTdsYWDNdV0pvinXpujtQq362ym8jRKklp4
LJSKjyNe9vxvd9zdIDVzE5ishoGks2mH5+L10K0ko1+DiZBEq0nnXZqGrmrcjqyy
niWA0sDn7jGWOMhb72MVr9AO6iVLMPcopP2Mwly7JYa7KDXCvUWMUcEpkV1Lagct
gw9GINlGwLn9HeJXIMdsF3Ojv7eBix2drc/YUI9VKOXNeIs1nCW2hm4nNKwp8/Hg
YPoq30h+hziboNliJUPOV/Q+h/o6h9pEdHFID2uVLk5s3p3h8//vUnEMdMnB96yA
f/H4BZzu/PaN2i22D+0qjBgAMt97Eb873J8pLLlRDmHFSCfxFVppz1KKrk7ecEFY
pP6W3TeQM2hk4z2dQoi4aU5HJVue9Xu+uU5s0iPJ1ZN2YXNp6ktB9BvVBYZte1Yf
Mv9VwHBRFKF1r0Vx2cmEkeBNEkrcdx0y/sE78SdF21/MENx/V6unJx2o4DyvkxTT
nB8b3me5Me9DX8JdF1+zNkboJxd2JuTO+Zgj1+TMi9OHRodLpcqtL42qyhvNXhef
HqEiOCOAJOGplY5+ulMmYqkhmkP4En2H34wsA9hlNReYdZ9vxHcdstlOOdQIJnFg
mgEGSkgB17vkiVWSH04i96ZmYJ7pt0l5/tgJW7opiQSWaoyUbANXjXdfVHT4yvY3
r4gMmHwid0IqN9zk+4ApuhrbZxoquj2FiO3sNKTdqbV6wn5HqDa5DJMJFz6TpA2R
iC8MzEE9azZNX8B4jMUobB4dcPBGTPUGr9z3Bu3+NzdeG5VnEceNRUPjiWHHKj15
XqA7FHIpqhyuSMReGcEfSoegXUbOSyb0K+uiHyjReBCh1kyXmPrGKamKY65+nrA+
QncwGvSGE15ogfR3oplnLEL2DXqc2cFGuQ4EY70QcQQ=
`protect END_PROTECTED
