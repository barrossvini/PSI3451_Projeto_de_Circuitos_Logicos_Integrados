`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C9GXhf6K4rPlq55cVdOKNNmPWn0T3UoUaZqGHMkJyQJraSIkwNYrn61McT014wjE
3/bAWnfNAYnQZco3Kr4f2EAEy/oJDt2/JeTxVDawrIUP1TPf5KVWCnLbrP/KBLDg
D3VAM2vKlJF1Mvdq4xV0+XMMYpfPs1R2BcowUnAxDqy3dgtTK5/yLEdd8H4mrp5c
gmaSwlpN1WnfrF7Uyd8rVDLB/rAEAQtgnBEXfL4c03leh0EvILs//5nnscy0+Jc0
l8B9iW2ATZ0DD6xHwB9U+1U/NeCaL9sE+YYQWUt19HT/FZ1hPDtYf7bKWhZaDrrH
zX4YX2E34a2OVfwGg7NIggvwb7Gwa1EhUisuhWLc46KYIWIiV7TboOKt36yrWl92
tj0ZRmXtURsjpPqB4idYAn6YYItWfvPSiQ3mTnfdvAVbwNdVxXXieCakpDuTibPt
vSQ8YnQJc79pioYeWfRwyBMXOWHqKTpCWRFPtcgtJEupeJcgDGZyjVjfBM0PkWy2
aDSYyHcpHXoJfd6kG8RtMerHKi4HYi8/7rKnaUDM0wkN0nJ7+sbvqdX9FjbR6f3j
CEaXampMeBVc+udGExew91POsEAKwKjGiha3nIwec4k6Y1E4QHvqhbEFm0K3l1kb
5w9xxv99VD7zyKCqNFFNo5Hf+pPdbdSSm7Sajg/fPGE5BRXdPzYoQjUx4kvhfkzM
/of0mtCSyCUS5z9dSwFqawP56e3SFic0opbktsiPd5rDrHWCsh0zhPTXOjXUtxzK
QYhzu29KD3tPCc9m7g4vjr0mtxS9MBGtfrU8KdXoifxufCmcw68pDHxJTBMOjjci
9E0HwT3yIVgnguoAtGlAFO/ezRvlv0vwJy82Ha/Tghz6LNuo4Z911JAtFPDTNccY
fNi8rrrhyM6MqJBrAkWPRaRO+25ufTAHoyfVV/SDi7q47PreatO9mFHBw1tT57t+
b0JMSFOpfL+jqoHuEAQl9rgseNazqSB083Cu3k5QDnhRJN0S5DiwoYuEi7GUYr4V
lpYNTxNOsQ2N5AY5IeqfYeOyjrCuHyd0iHDv9GxsA1CfkoZHHMbzwN8XfaSR5qJ8
`protect END_PROTECTED
