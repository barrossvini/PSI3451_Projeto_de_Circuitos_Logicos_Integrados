`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMX7r0HnVD+EyU4UddLD/Zowzr/VbcsvRoQ/5D2nK+fqwKyw/A2PCqAYZZEqHdeh
1idZqp9l7fygmVMuWJunHfeZ6NUM/0E+qkE6M60w3m5We2IW0JRQf7Hl87tetnkv
lpltEj9tiH1RKRif9INY6aNuTl08GSuoJWPX7HnyjqxH1ULqhmI/4Yvsy/fOFLn8
27FlYsX+O3cTHck9BBtr67wRObvOsL8ciY7vnD0SVbZgq6Oe8b4OJpboUebBsbNN
0saJm/mLpEqv577i+ifX+T+C21a6SIN21thRZk4KKASfcGSmD6NSH0erqpXNwrb3
MzCKfQrxjYhcWK9omXnS72wEfGNIZ2c+hDj42NL/aSJmczzTzOkCX1PDMPXylKfl
T1PitpnZBbLerGrHRcqpv8sXgTOQQjXp08me4gw0wdQ2tfKGJvBUgW6yTo/t/zfM
jUHkx6CBRZcX/nwtXJp/YMfzFJIDWDjSqBC1xJPmugDocgZxd7RZto0dJTdrcae0
JEWHwLC2KLvn5lbXb/PlDoldWeA19aIXg+c/3uoYUlv0k/hv5N5MGDZ7t3guVfGl
eh0WI9t3r3BMAeIZUbNj8A9k/xIL9ltVJWPzIbO3dhPHHPEh3XrmiFGKPYQoG+wN
bOWwQyU/FW9wzmQhmWDo5oAGa1FM+glRomrt9Ipk94Dc/0ufZuOhy63bJKHBFmVg
pnbe0IzEkMeDO4zU0Ku5UNbCAwODnxXy0xllk6lTuraQDAmVGdu2cKqoPLPScBOq
pMdw755GSYyLh80hofpIiTXaGvG8Zih9lX0Wa0o/1OdSyv+Q7ovquRGMfp1iRuox
xDUXE6UGI0hec2Lw82HD++t5pohc1JgnjMR8x64N4ORwUOqAldN4d8aVK8G3DFmE
5uk8mFQPLX885IElABRdFahkYu2Z5UHhk5lAw6IyKL3YzvmTh1CIwgK9b4utwswv
S99ZIX0jqog5U3KsYphV7Fte+T1+VP37GkMpMevbcJLZrxBSIXpJ/rZ2sYOBsqUQ
6lGbZImtYxfcoPn63CwHebTpvrCpfEmYi4lJ0nNYcyY=
`protect END_PROTECTED
