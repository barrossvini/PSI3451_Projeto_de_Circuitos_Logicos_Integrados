`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PE7ptJri/zebyk2WSHt2wDrbx6ISYrslOQRc2VMGxChU0O0/KnPY3EVQvVb2oT8v
4byW1qRfhTeTEMKwdSvQCIe8raWaUu2UEnLgcenR6rtR7ml0Ca+QTOq7iW680onp
7mx66/bDTj/Oy7PQVbzA+cyf/hcN9Yz1jMIXl5yIGDrdlKBiiFFUCPx3BA4/Rj8U
LwunA5+g5fZabBqBHeB5hhDRk8Kq3sJhNsiuY/2NErxbwL4rmA3eXEsIFEP+Z2ix
GhB/Ar3KkhwSljwNT5nefZVuC84jGK+RV/Lbq9mHvqWOuDiZGSxgbxh7APe1+H64
jdWHuLKaALf3OTHVHgbjSRccr6tGJcNdsJmwT/Hyz42XKoA4IuZlKIrGVH/3L2CZ
ioPhtA9WgSqA0vbw9CMN68NrXBwrjlLC5XVRMNsDq+4JaD/++7O0Hsx+E5xjrBpp
YuxxxZYK/AI1NYi+H0KC77ihZoWpmrfQ+ElpevKOwp4W6d34yLV5IVhWBd8zFmA/
CJmt1eNbVW0XtfbryPVnBt1GSE8gpjUsPX9dRTgDiKeU3nFJju6fKuczSlZRao4z
hXj2/w3NmfLlpQAp1XHYVgEV7/zhTZbeOpIkD4anJzflOwf0iWqtH4Q9lDDERZj/
qukEESYgheaC4eRTsKIX/enDRzboRDmtqCVUClwDkKS2p+QtgAjE3VloyMKlwPoc
8hDGq6+6TLelEzjo4iaYj8mB0nkYpWXW90YLQWDkjKalKw6Y8xM3h25vzYZQ7Da6
S5DAhaXbw/TGJThbuaNqiXfKON0Zr6A+PEFuzRZfr2dT3s7roqgaoAubUAkeli1P
9uqn3NFmrP8kwe1sLXJstB6xkVPv7Xdgngnmg35q3xGA2g8O/3cw4/oQY5o0wut/
Micf9CeN7I62J1Br8FQz+UxSL8bM1ddDszbkWTvT7f2h9iB1zkecQ13YlrFMatS7
uJPPt2H+szZrH16vAXg1cYyCMB5XvOcIVRgeFG3oiFUxJcmfFkHMYSATVdBOahfl
LBqpOUaDzVU1dgLrkI1l/ebvUOAql7DAb+TSAMvUUZLrKKi+apq7wR1AI8c7snwW
z5HgBLhmomWwKl5sD3AeFEGBvFrYi3ZRNP8d/1/Fo4afELvTVo1yA4erxK3nAkfu
UYDI0PVPzKafpVVgypcM7gOaHJ6BaHFsHwyBamCq72txq3glWPtpfus/YoDxah/t
UjDkSGdPUDXpd2nu1po51LmP+76rlQbQO4iKuLVSsnRqCt+asfCJFABGKX7lZ6Ld
1QSjsf2TGspbs986dnrxpTNjKkx3FaJ3ciRaDZRKGcKQE6kHlcawmWnACArZPjuh
SnwGiffJCfWU+o9G3waffyEK/GH5hudSzV70kro7D0T9blIH4i/NBQ1sSwjF8r9T
EuRbwv//kdXyb/4sKKzXrlHZU6SjbBD9nDOWkKQdafpwoARlB1Dfv6FLqZd/Lmbf
RV5S3+zTjI8gdqOb7dRF8pdqkMRZw/q6A5rpK3zw843BV86Qyxmxh1+jyHgxZtYF
tCl/PxVOH7TI+XtWZ+pF79wVYcLPWDviIrx09UFYJORHpzV3qP8fp6JjUlPRXX9e
J/MUTJCuCb1xjJwGX6B4/M03YLUor9nTkQ8WA5PDF2A=
`protect END_PROTECTED
