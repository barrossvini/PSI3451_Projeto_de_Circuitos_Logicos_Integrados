`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5xDPPYSYSatJ2bjKxWbbTPOezjLyUlIPcVv1FSv0ELOiYVxPyo0J+fSMNaGmoQfe
0V/rJO8ymVqklxRsQ45UolL+exahsuoEzvhjFjfMNcA0FLA4+hC1Ypb+P/Fn6Y4T
Z1AnBkbHqFH9whTAlX54uavmze5t8lmHK4dXx+YcLzrTCmFnYgDcK9Fz+HQCYucd
23B93oSYnwrZcQ77VGJ+OEcSBqI4JdBfh8pPpMTIozMc74A4c2CKPyo3OlE6PS8p
v3bgdMDOOPeS3faryIOmDX/w+uaTBkGCpigvl7qGk6cl3hHai9HNQfpR1jIbiU03
HPgI6N36ZtLSAPJBf6uX4+aqFkdYdmKqy0IiQMJZX7/SyUnakcoaB83MpjrUSOf5
mxJV+jRrfi8WYvVbxK03c4G0NY5Drg83ecWmONKXl5CfALcswgTnrcOfKRfXQgjc
HOnkUs0fYkx3rCuTy8Scd6BPiwTdTRn0toPIcNtf/CkzyqAOF0h5JKt+hyAyp+T+
i3BZzdQwZTZv+uX4OduXpcMs9iTLkEC/NRgjj2ordFMdVE0FlowORkMVMNFFTyto
wXjCWZQkz64Jkv7brXTcWr3QvuZkOwK43jQ/q4e+6W5YfhirRwQ3b2hkppolzY8g
93no/hSqi/hfgkLIVI3ei0Uf3Q681wWyBR/syAkSiQnVwKJh1amVbMe1Ip+Jep/l
G2gZd2WN7bUQHgd125asNBNhuNcEmLmN3w3Ym4qHhgOzC/BlkTsyCkusSmIUJNty
M3nrnJQL/L6jbGHSbqlYLhoptYO51I93ZGbVIY9rz5Wh7VYxhEvRMoKdlVrufoYN
tjnacmK15L5WykeO+PsUk/eeCjWZbX47HzNkZwTjFgOePOSVaYfLSF0C8g5mC9Ie
gNJQyqjVvcnoY0DVtUV7BKD73tksrTFoAzXrRoWzroRL8RdgfzsqmoO148u+6jn7
epWCnK/bq3cYJ1Nhqlukt8fAT7ThyWBzHC8i2XRWGRchpgft2jpAeck0PEwinHvC
NImGxLNR9g0VtASQUx2SiOWwWSnG8bo2yqYSZ97Aqo63VYyc3y4U1OeA9OVZdAt2
mwnH09ODZTBY6ew71BaYo4EXHjxtQthIyAzBJz/AqdGxRUmQdWWhTzZaZASN7r+e
HTHyWtVcrGfllCEJJCLGBzUSQtqAHnjmpStxjolOdbBCwxmmEGv6rWQePDGm1nVa
39yeHQKsIMQAWg841328gZ3II0gFzzaDBqPFHWkg0zbtPOip2UQuSmQTueTAmon8
krTdDuG3DJfjLaWis2WQbeHhSQkbTw+g10Hn/V7W2jkd2heqhqrshDrgdezYIXs0
dDWB9rBRRKB0WwgMQSTpD9wBUWwGBq3PWsc0NwE23QXmI8bic82MotLQYnXKERqr
mnB8kW4wG9d3PkcMLJd8S3GXTWFB6ciwn5Lm2HIsGlVLVCqEK9JPifoo39cmRqvX
yg24fWmFvl7mbj9HABXyBZPs53iI0BVc/jIVwp29ap5H46dXFzoxArp7cNGFKIZg
6f38n3msi/z81qs2MBVTTDNTpigDcYVaPbqP31axhNf0iN6r2TUkjWXKGRMEE33U
CoctJDS5jVCEs0eiUcP54M2NyGd0RoRmOptrq+dD/4plze88s+pq1nxqwUB2mfVO
mcsS0qCcUiSsgufS9dmXBiaocNIyESvDrXguCkyM6nKgLPLzrufHTmBCedh3z5SQ
4fcEBJE4GuArerMjNcw9R2j4ebUZfxVYKmQYN7Mi3reIxF5wggT8O9wVVIS7/I1M
ho8TAhMVRHr0qPJ0c1qaebeetQXTV9YOqO9qw94MbTROqryxULSMmPjarWdCEqUP
yUvpaLOW3kNyox2Q0kf9FaL3Irgyg9AjzvSzSisU61fiiFg78sk3dl30TD+k660+
2MgnzK6OPQK3xQRQLDTxlNWe0/BpFCgOKJcmRJV0uFVwszIoHcUtel5UL5/1G6IC
ncRpWKe5sGafkFunpRztLhj5Br5swDTNFNCe1iUtE8+IVSk3wnr94RJS6UaNWB8g
3ZE20hjiTt9PisA9bB0DNxT8dHErYRNvmU3aG0GsiYyeg0rSVVh8pu9EHMqeLDAu
rUBGRWqWoeVLZD0IaFLszz24W2u9zKsfYe5kc7PpN4gptaPabPfayMINyXy9kKzf
ovNRo6BQXbTM78ZY8ehAFKJZF6ow5uZZb7BlZwE1MLLn+1bEOvr8JFZdeq6dlR5l
4dMZ4dswyQ3wpBWr4GmU+pFjhsBWV5fUAmfRzM8E9jPTbJ+R7dVF6m9/+8V3HlKj
Dxc9fWQqfTgZgpNcZkOjPsGQP/bwoFnFImgc48Pf24X2zzbxptzPyIlcPO3GuF+I
IieLygONceVV6ibOHX6Rueb7sPi0t7DY4T6/rxOmavyCdMhwW4HMFdhsQtF0Bfsj
k7ULm+3cKed+KBD7x2/0u0lNH+cQzrcbdXhg1qz0uml3DarDtZO0UVa4yX1lbnh3
NN5lbGHFUeYaFlfb0jZACO6npEXQVzn8rXJJSHsAVPx1l4RiY6G9fY0PLhCBArJo
6As8Z8q71DFJCekGquaHEKp+NYjflVUwoVnBaniumYBag0VOxzXgBkR6gABi9XWo
fC+hqnajlQSB/+oyVsJEuUrFvVTwudjATkKy2AfYA2IQE3GO+M6kljuZ0hrTRt1S
aUgfjgVseY/rmnfQjT5AcNIoTc/VegvIiMSc6c7bz6oIFH0cTMWeGOhJjNMRX+W9
J3d7J1SxNYOH7njEAE3sdX++/akSvetFED0MaL6evvzj+lwyxVG96gLyn8Il2ow+
pObsCvwcjD2Wp1yUQTmVOJIUVe0c9wEnzr15D1aSQCt5KQ/u6F4zXVyUVk65Ys8K
aqYQ5Fxxp1S8FKuaa7IlemxpBXx547p4HxWTuJUOuMYlxdZxaHUvvPIiCiwTLTnE
heD1qoA30cfqFJn2MLDK6ndtEMmmkQpHFv5XXyyMh7r1DyQ+OEOEWmUDRooIXK3D
sQC2LR02UTPIvzVGZYnG/lZBNcx/aZWB1hoEsizy+FMxX5sNCP56xj3m9DurnsC4
JEsNSAudDtN1tTMGU8PKNV+dR0EiXKU7epRivRGOGvmFJDgzpZc0b0Hva5Ca3DS9
dLJXeqL44Ia6YdRW/t1z8PJMUqfojYElbsO5Rmfp0dECXblriZ+HjWiY2GpA9fFL
/IExT7vCb7BakvbecX3oY5lwqfERU6k7eFWQzbm5f8wuWaDLeTrdCTzeAa7Qf/3N
jdfp6OLIBU0ljw6FH5A/0P8SiF01ZAhhTONyn/twRUhPGS1pyvGWYTtA9IvPRdqA
v0igZAqyKzEW88tRq6CF0TtLJaFaHBHsfF+lFIryNs1Bub/V7cT++O6yc2EOfuB1
WcXYffBLExZQ73rdWTK+IxWSyDLKupgUulTFcQ5vaK3FKtgIsyIVkzIKv922SORp
zkp0pQFSqs5JD2yEd+0ecwBMU+1Rm5hQZbyPki4h2QscEGzT+QxGFb1rU4RCVZRo
pexjkEio3NU/w+GjdyddisuN7t57IJDBgkGw9v6YzNAxx/pCK3amPzdcBSgdEcX/
Ehld9BCUt4C+gC9fiXTZtxM55+8PtnIAG20X2ax7LCI1ok2SvzxbDO5XC2cgDr3c
ju6jNLwL2aiS3fQpY4YWtfkODU3Rh3EsyUeUnXfFodf907diTFftTDEJkf+pNVf9
e2TsUfqI07y00/r7hEEAzTMsiRt9nXUYni05rc0DFxyncS59XnBOi7U40+Y4b5Iz
WGZSWS3KW4/jaZzp3eJYcDkxqpAreGvWqIrQql9Fue9J5N2nKXc+QQEifPGlXT9M
bMkNfJhR6bUqjMEPdBkNRvzWzgmtuJedArhT8TMEuJ3kyO+6/6R3V/PN/g5JG7d3
3WSuqdMV5fbMAGdrfqkqPeFKCCUZrZIDPyNcVs1JnkCsMIB2a/6Ljdg6vMQMnvUI
bDFXjeQTTDD2OBbxYqnbtLziYMyUugWUa8NzefiZyD4bQXXnky5/y9BvPbaR1BQn
t7ZKX1kvHGT8KM+w+yv5+67ZIfYCh1QsesLqlVVbpmnkQ996NroJ0E7J+RGejScS
FfwJHWO/cwMp80pE1sckw4JFOv5SMw/FdMxOEax21HKNxmi+f+dwa4vhSBcvwvQa
x1Fl6PoM4G7m1c+TFhluKd06oBU9q7A4zTZNA3crK5XQUtV9xMedMT8J/1r42s8B
pEFgQiGwYD9svNBor+FxYlz53OOv1xQjso3TCxqWs+Dv9JuhaaYEpWrxFh3sHyOK
vTPh2E71vUQE4ZmFH48etvqCjIyqTjIbwJtEoi5OKjvnJGdKRW3clv3/cIvn/mJP
D9lrwuqYvQuVzyeqwr3vAFq4/CHXXcFwZtzThmhf7vY=
`protect END_PROTECTED
