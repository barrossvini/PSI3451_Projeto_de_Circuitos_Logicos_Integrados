`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EDAfYYOP1z97Hr6L2BjwellUzpBOUsSpuCjdjz76fTql0KEkCLhVCnPT7sByqEYb
KqgmoI50dEVAjbmA+ZdhdpCQ3S40jTAFiyXI+4J92GbxZwC5zgT4j3J8ZskBtY/C
pjO3T6XxZRuLCGZ2CxOn1tlcUW7bcZhFLXFsQKhqJrdFwX2s6Y6hxkZgbDqgsCHV
4lVwcF9Zmm5XcjM3h7Yz9cQLRFmhk15ByuukmPgYOJDL34SKMxVRPvnjopzVFgV2
D5MQaKaS5WhTT0AtwIXtQ7hj4Vy1l3hnlk6Zg0KQGzNjfmpo/IoE3qM5utk5PxVL
/P4lARLfnAl/iLN2d31alIYYowSObJfgBtJlKB6zCuPUfdNU3GRvEP+aXN0quqZv
nu24iafhZ0W5dbBI5G4AaVdqOvX29tAKGxPQEFV9vt8sCKmGQHbNBh8WpeIuWzlT
Ac3CSj78B8GnfAaJKLODbjhfQKk+7zLI6Ovh1nGFtiR+jAG84oX/ueqxv6CLa9KA
n5N4l6/uHt86v3RDhg4ZZDhxgjFjG1YVN4evD9CKR+QO7ycKafDYUcoIpQubl6j9
akb1RPUsoNuqF7ieCBH3+uh0RB9E2igPmt6SAkK+JSA/zZbgPzU6/wwOm/NrykBW
sXFqK1I8t5xBbAVxEo1EeEI9DI9waSshvpPdacfR9uLi2/KfcWnosF5gok8O6RxT
WkaBKpVFvYTTXaFocrVQpr2Sv9xn+N7evT4QPa6VboXFbDWGsZOzxlM9vFU/nD9/
Of0L8xjDoc/8/nV2TiZIvFOvbtS550vBTiN6MjQA1m932QQNRhGjP7NKxsWns1Al
cynLmQNHrwTWD2Q8mYC/x0wiF/ImJ8dvldf3RYPNaD9Up5Ev045z7vcgZnx8uP5u
RyyKyvCum/Sg/I/2Zomwd5jTKt9ZcElAwMK9zK81r8uz7wxVQFYvXqKebXELFBha
+gkp+TYwAcaHymrFG3d5pBBhc59M02OAtM83/3MJCeACVeHqRWWj+u4d2znEqhO2
K+CX1uHPVfVlC7Y2a2J4I5m13yjvHqlvoHZSyXBo0gDlk+ssjsPBu4SYQzYQlISw
M8muDqbqtZy8VHzD71se8sJYd9kCrU/aVFWqQeNrO8wYhzfrpHkj1pBxK61CXSPg
xQH9Id99V07IXhBfm8UHlLdTYkoHUk/ix9zaq9uvDNIUc3vZYUSBLDfK1UDKM11h
T1uOKs0lOxXeV7d6g7U4ms0Tm87uudoP9BEy2FvKyDIevk5qk4Pky1ZLeBS5ZjXJ
C7TWiHZ8hTYUoH+f9KnbEj/RbVafgvAURDxmoU/KskxoCEvh+MwevGaFND0jTl9I
7hGZaiWLwm4Pf8JtMUAtRSNTBNLB+vWW4H7mY+d4Y+Y+/gAEmeiPmvVI62dFq9s9
VaEb8wR7H975UOqg60lKE77DLtkpkygfUwjYYqH/VVm7KrJj5vzDGHnKP1JkL4I9
vs5GdLZNT5VK795NP23WE/zMaYlWknTfwsCeBPPSRPdV7oSKkWpGij7bScQI/vNh
XeZwlKlakX47uB0SeZzUkQ9iUtdwz3aXdEjTtrui+4TRchzoo9AJW8S/Yb97rs0e
WwLE3iZU3Fm9MI1nB1iWmPrf+UI4zQgPhCfvWbfwevi20NApNAFTGSV81k4O5De1
0lU66W5bo3/W6Rfy6VD9UHGdDc6735icRc6pzi0GhhXxdaor1Nn5WKIp4YnPqApT
CcEOiFjsUMVhNWAdoy8VeruLom/v/+dUoyeh56NZRLMO+CJZrbfxmNx/vATPHRrC
DBFbRJDSiZmV4Dq09kr1QRdkju4L4TvmIZ+ugdw8IkBE8UN/HtnJ0Nj8kgsbtgUd
Wn5SeEmvlY1f6Fj7eNSzjxSyNO2hjrzQG9xF/+ve/79G96/e+DJBd3DybS2T9816
geteCBlIO6PxD8Z7nbl5OUslXwGwKrZTxDiwHLVRoH8t2ri7k9tfGcXqRxF7vKEX
xkoR8EqZpwShfFQd3QBcUY7M+CVT/qKqiaSx8+0NKUNu2GHqzFBcJVU61JUYvp3Y
mZJqYCp1zKpepKm7ZhiSQo3awMZopbv5P9+8EC1eaGgB3+wa1o85lVTrk0KuXJTE
dBTpU+DEOX1NPchc9v9Ti+utxfkIOr16lK/7A0MX9BBHgIt2Q927ReT72y76a7kB
PJX2/aSbsbwmAzKGCiKcdeM6sTK4bjdqr1pDuRiEailTTVcbhorQCbqpyfart+4m
8PcuKFny3LdwqqJIXRtiwSyM+FYNlfQGUlyr282+XND1bpPvllwwCim6bldpIIrR
g+YIWbG3qZZbo2Kb3rnXLg==
`protect END_PROTECTED
