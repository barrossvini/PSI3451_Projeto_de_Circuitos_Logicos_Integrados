`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rz5fLNFxLtvE6fGpOLovU+SrZ3jws9Uj5WoE8speZkw88Jcz3xf+esanSsMTYucM
vZXNppw5s3FbE/4q+H9ZhhY8Cbsu5mTF0AB3rVSRogsXrkEThgr2++9nw0MV4pac
Qzu5KEynqjWH1cz/BgYtL3VpIhNSQyRhstNK8k65kHQjFPjcfbIydl+wHY9IMHBM
4WgFYVxDb+bCMHp+nTWbz6BQeWHWepTdZNyuMCFA0i1/5EtGsIjUFpwPoDCixq6+
sZLtcPTdWjEqcWbqFJj1LRq95DKy+fNDN50QUKkgy1KaNhWXvLHPkCV5c3Z2rbcO
h4C4OT8p5jSSe9a/LzXvkUKcmKTUkNtHl451Hx9vW2SEuF+HROqFQHMS7eGV2jBj
oboOKr1EVQZIlZpBZVliQHsW0Vo7JBhfdeaKisv9d7X2HcRTYYvr/IVWIgPXwv8Y
mTSwE/07a7EigCIosDDK3a1LASHInfGU5rU7SJh1hOnQK3yESU2PLOZ1HMM8LmR+
rq7u9zG0p2b1tnvgXujwf34rFblU4L0byKW4DahYGVsUx7K7AMDBFFc3BM9kly3v
NOPX+nP82hAARErw8w54No6jHnzILauLPFSut4MLUgwDE0NxQiyYfJNKOErYpFs/
GAdwYnCwFGihJ6cwwwWdV70rLRLQa9JBRdKwSHyBealjQ53/azqXf2CphEjspvRX
y+WHI2w5JG1PDyscico/tDuVBzsvwzOs14q8SQJXdMVl848hZUdZy0MJu7HlLMDB
C9SpXmeh3WO0UYhxTdioFFiQfI8vA8DUAw7TN6UnqIEIeG4HBBN9Fy4AuUtpoqUd
LfZpSm7SW3sQOVWrugP4fiR9A04yebkxi6n027PspJ4=
`protect END_PROTECTED
