`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zsadiYz6dHLx5pJdLJioafwY7mHFgqUCwPAAoGzcgQERYCx7jWCrVQFRCsUwkWRX
JOjaN5MRefYQP3Mn2ppC8YAdN3x/L7STHYRFE2EWZWQlACabU0JEROKPZx3Dm0Lg
+PAUOZht68RrGsOvrlGa+7Z/VnHtHuR98Scn64CXSw8a54Oi6LpXtxzUjiE8/16t
1suit3pUjTH8ywIaQxqMS2ycgpGepBnXVfPnlqTzRsdXOQPOqEzoXgNqMu4qRk3x
IeMdAWME5LkjCXAQDL3ZlH1oE53nCqoE0bBQ0Qh4Zymi5x88FB46J/T0VSn8w+87
WOUDKv2rbHSMtSvNJZNTkconG5oPE5G9DowVsG9yi/qP4o5KkSZgV3SwRkwNv22F
Ez5vVKSFyauxmHglW/GX+rGN7rk0YHc6eBaHjTNAlbd+TxqcpeLo+69As1f3hqiQ
3Fn+TyEzIbZx/t9lGNRItV572A/fXthHuUMtynxxoNGlVgFZCanp87/4Cdgp7mBo
jwNQS4XLLKyAElWuJNjt5Xs3BdkPDUCSw+1JRdpTn1eSJoHLUBO+LB5PXPM8771q
3B83Rtaki9ssDVIVLw20TDk0+IxBADS9Z/gDZaitjKVNGiVLCFM4e5L9M/Xh2D2W
doJQGlfVhCag74toPtYhH3Y/pbSID+5gcPFRtGKQQoSp7YxCFbxEvLtz3bUTCqAd
E2dN5eIy2s4tdrR1sauKgjc/6ZajSVuUbJqSuFC0Ub52umNGafPYaOpVAKRl7SN4
4UvMqccwnzg5FGSjineC6CAQFfS2lfNy1CrCMmN+YMXvz+hNP/qC//raHuquxUDQ
SCFyPyulcoPTy97xN4dVKw==
`protect END_PROTECTED
