`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRoe1+v9sdv6+hqbVzv5sCI7RKr3dx77rhHvOmhNNaM+z29Pwa8ESF1SE4+6d6iy
+J4qx1dAAZvKD2/X8YCwu+oNFVFDtcjJlh/1RxJqOaie9sIrJO+H/GxIgOjhsDpE
EVfNuC7kq0TRdl6FGrYhNv0kdyJKsS72jg23r8Yyf6FKxw1L9bSKVIOWTuoQTlB9
TWt9awJib+F86rRPmiSyFMykXaTx+Ce6KJrkyWNKUxVevvcojKbWmWQXlzPDeRbe
fcEdfYGd6+aqlTbDhgF6BnHT1jcctR3qKxXbfAitW2qxZp/9Uva2nMSIS2gaW02Y
l0GMjlj6MwZa87kZKqw4Gzt7yWoxgkkDCjrm/+q4ErH67LUAWJrUVYjXurvx5Nlf
ZGWOWBf7G7lrVYLn3Sd7YTOMC3aOuhB3MJS3tpDaSXL1QF9NP3+OQ+Ocz6BmJ1pL
DdRqdffVdXumUNFGkitFJ5JOiaZ7Jf+gKFUPNP+pVg+vAE7BQv9oV1gbHl2Bv/VS
UU7eHYctTLHUjfT8zTiF0BCrBD110IpRvZlopVNTNXSrE4Abj5mfc8pkDxyZ2Vcq
bvZz4Mn5jyRyRAfQmK+yjteEUgiBvJzNTag9zwcfAOPBmDPrVjsgFzL04j+2sxcj
G+ZwYk5xOx2UCoZVWGFXtZEWR6Vwel2E7U6ENKtgvJ9gLcJZu7Bqta+zX8UKxKsV
`protect END_PROTECTED
