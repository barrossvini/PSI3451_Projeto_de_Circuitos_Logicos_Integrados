`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fC0PhGQ4gqYM7NUhBEM/JvWjeOvfXH47sjN/vb7G4Bj8BjC5vOATyLP8E5tcxCB6
7+/BzZKAIRVdbV/zDMQ/Gc71Kxvy45Ryt5ZsO3jeNalnQO2PnSloGJsdlW474tb+
q0jdXvUAUCglECaW4uiBYykr+e/8CNC3/IugPWIrT4ZPV6WSCrRdV4QeBVJ9FQIv
zJzYPGieXc54pE9OM4NmkdixPJ+bGXqyB8chpKs5MslVoFMPTT3pTwv3MycJjDFW
bOvCdyuR3sTaKEaua9oiROYLNl5gv/UJ6TbxQR+/nra2ijIbCJ4T96jkW7fRyJHI
8J8wxk4t18Ob31+YipMvgTHYmEN4/mgdKoeNDnnvKDWK8CPgNW2ORJ0sMAd6cn2H
ICndtsP6ZtySkkdSsyYJ5dJae68P1UOVkrZ/qjfYNJhH669AYNNJ3NRdWRRzZdVP
eYNQVsfdOUqc/aH5vCV/d2G4L3Q4SS2LgWJV+qRp1MDERL5cz25fsfZQdncqFcnT
ilDukmLadFt1VXr5K9sQzCK39P0A2H+kBondfQJIR9/JPXsi4DWY+vs+PVjkN5dD
arcUwHSvIjidYhP4DvbSAJOGNH4vLDEGxTj54i7uKxu+hW/gDLCQQD43EowJ4qkn
FhhDmwP1y12bn3g9RU9dAxln34oHV2lsrnigUF15Y+h4qed/7wjALepwVrsPzmlF
Po0ov1Rt43TqCNwR7Q+ebllUJjfIfOdbClTFSeCtSugkuWeDtaDLj13oD3kcqnYd
YMNCGXIHqXTU/ulcOs8Mp9cY5M7qda7c5pcCIcsAHo+HemPbJtYJviU9HKFvbeOa
PfOHI4Yi696I3EUuyNCm8uH37pSNJrWh5yHJfi2BNpEQkS2oXYNR32RydQPTkMWz
oUfe//7nTbHRNir6Hr2XygE6yMt2oPUidT3uSbjRpX/g7oVAZhfKCGLUdjkMI3JM
0DLKK81voeD2Khh4Bblc8R8c083m1dLphFeRUy1Fp0gMrdGpXLvKJgXT+dwhVwHs
1178LdK/T379UlaQdxfXEXaOd+4eb0yfsYLKKcEUHZmMfWIPIyKOMfmBko3QH2y+
um7WEFUm+ncCYzeQ4+AqSly0MRsYKda0Lhe1FV5MC9J18bhfzWHpmo4u+olpPUhj
DYtlwh7+hpVTydxAanTwSigCxutXVMvoiETbj4hhNnjg+Fg7CelA7gF1TyIpmaoI
wRk625rvtsgQeUHddjOuss3iy9PmsZEdIHes419YgAL6C6wipdpZbsEGkNlp2gwM
lBUBYXCfOcY9hL10cka6i2UzHrnM2vxvMupZutxcICsjeLP2Zv6+iriPdrNRXv18
ECncozvKCoQ5UaX04TLqncJ3Pqvj0yiIjIJJD+54g2Z5YU4ymO7dris7WbgDP9N1
Spv/hDVdORF9aZnNcIhhecKJvVW8WMuWdpok4kBdeBReeiCki7Qdg32XqTSs+iE+
ZiaQdgMDbeA8S932vklNDLSz8wbEC8eCC67UiyV5cN9fZs3ugkzGYTZIXNA8HPph
pRe6Eg98W02V9iA1RAXZzmzjJek+s9HBnV60Z06i7oOP3VlXEi9TkFxSeydCm/HS
L4z+XNIF3QXopHG2khruO0jDdW5EZP/SHxv+nhYII2iW2C8fuyNZc6mvlRMSFsPW
h8LBYEMdNzHnyw7nS1rE3VanzGj7o0F6eT/CykHOAydnoDYtWAtwsnhafzD5gJcp
V2bcANTqk1iyziH3paZwupeWjqIrkV4UtSvIKJ4PWiN4d2LvT5ssbXXWxCnd+san
MKjYbRlqDlRmXPxsJ2EKRONSky2v1gUA+JQ/YG5m0WmRYKl3Cj/sGfwcx9N54umq
Zacaf5IApElRhNR9kkAsa4WxzRhs625hUqUfLTDnEpMVEwVaQRoSGXgglAC2KCUi
UxoSw+N2Q8bLXUH79X7FjPcBuOCbf92fiuJ6xZ2kosAYoDlNMGPmxlqy+wgSClHd
3dF3mob724Jygl/BXtkoEjKW4NUtl+YJKzeqmGjAvrsq3ClkMERuV6fCygvvmyQu
nQVWitR6eth0zBzHTWBxsiBexrPu8uTyMooYwhUr1yCVvTEAGg6uWocY6JhXe0fs
yTlxQrQbopG8gerNhiVnbEclY6dZ+KKOLxM5AhLpnPe/ZpQsLrzv1dUniKQDpqoo
974hjo3E9rlcj32sEtR/3DimrzScBNhoCjnXXhUZWNYX+4zIp0OTc448jNuTd1HT
wzKGJw05DOXtIhG8ICMmaB3esp24PvppPlalmA6B1t657NxkR9/2eHOzZrsP1QBk
JXShZ579zBgA3mLlyMvMnbVGK9F+p/tU3I4pu8dbd7bkRq/2tk+I6Uem51S6mUrv
smnikz9y+7R0ofMeNaTzYZmM7Du/vuBCyZ+TKbct9Ovx1K3hBo2OVeEg27wlCo+Z
/keKNP6z783TZ4T4navEaIO+pxIvqIYOHL2fH8A18djTaefFP2czLr4Xi3CKNIlL
f8TyvFvjp6Qgmfyf/r6dJjjLh9/J3vAfIL7qBUj5EKSCBxdY2q5c/5CdqsgtBtb9
dV431vuklSLfdE+PvTq/CyP6aQCjGYRwur833dzjSmooDrKMs06RZKEwH3hyPPEs
KJtLOocrnIwiUCPURPqEMz7jldZ/+QmXxnAuYKZ6xjlZxYkgNI4awzI97iMsUQqv
HmJTl6bjSZoKSrltW7gsqmZwmEG/U1gTwR+113YVSST9nTzc2pSs411ku36BlJKx
NRx3ifvsfcqffZhtAorrr2BTfAYfrHuT50/s6R+Aj4lcCVmHrbyJNbjzq733FjTE
mSCe8DekdEBxCyWoOjZrttTQqvxVB5otqe+D+3RWZklUWMyPFBuL0w8NZ5Djt3UQ
sHPm74KT+7SFZd5w+jPo83RSujVXaF2dYOKTmBasmjtz/qu1tryusqUb3Sq82cQ2
HwgUr6niEXr0ptJJTxmhIsEZOI+Kt1JbJIXBxYvuNuGT3AZ8KofkBirHmfVwKR+z
KRGxLiEBStXitZ7pbsYafghPLJEs9wWjrL4gY49h/lVK5EkSuYQG6/2/JxenyR0T
KGMaj4CYCCT9yQ8c0ATqThULOL8V/WZeeJG53fbVSZzRN/AqRlkVCTZk6QSqisbz
LmHjeWwm+gvbqRSj37ydUjWPBcjWybimFmuXwuwgaUC8ksqUPMfZVRxEHhxJfxFL
K7W8uQ9wALCUIUop2mOUL9dUZYBPl5UsZ5n99joUuKl6obKy65JgjbeuERhu9Ev8
tJIdeDLp54gSRXyn7AGCg1Xm8xLu6mV7i9+nSKN0t3L9OHhcr6HJXxY3rwdT4Vta
HEm3vSjIBskXUuGUhcmeeN1CbU1eUPNfU/v8n/tTbFwQ3Z8urkdGON5GqHieHWnW
7YhDhiNctElR8rdh5a6rwy4G4+9jjT9ZvdeNpBRzglpKdxxi14yGdgYEwry+1VRv
OcdARFdh8GfvG8mUWW2IvbvMFsk4Ve4PJr5p8YyyuqTpq2iTzypbkbeDsWIo0noR
gC3rK+JjUq1tyBmGgMc2RhlI4CuX2AU8j4MIUz0kVtMjFFV/2CeCc/1oWrPW+647
dItRgxbJWaxZ7xaPVc/1Av7Az4mu2A01Vd+i5ajxmLQV43GF3zDofhjjxCS5W8C3
8LTa80xVoLEjPf4jarnvyHNJDXkKkYJQ8l5kIvVfdj2aM84Bl2qt0uDJgUhhGKrG
+1NCUONm/YrllvRM1pj19A==
`protect END_PROTECTED
