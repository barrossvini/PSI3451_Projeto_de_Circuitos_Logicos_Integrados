`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N8VB3tJ9f8dYphsWmFpF3lyKFDuuddim/Rx1xAzQThiQB1RHOucXDnvWp0EDjekh
xWpXbCrWqkWhcdTBAEMWFvP81FHcgkvkHfHEE3VwFVU1nNJD3N2aLsKpknMuYQNp
bicY22OgiFIgASHBEzGtcdHUEZq1WGR8HIULj6Y1LmVlOAbhz/M9bPUkg801kw9F
CRmNeW9znvIA0nEqqcou4WunEPJbOfUS5EUcTYhMguNAq6hBKyPurvXt1aIhLXx9
qeAx3ep9KAkOAPuABAlwziV1PeZ19LjhJ0jXiHdNTdAZ2c/quO2BIrQ1l7qOIJIw
BBQzpKhMCC5HA+/YDMH8zTmfnEwRUtSwV6AVHnJUgUMNXCKJWRtWrrVQt18Z6fkP
3Ovw4sXw5fp/BIJDa/goXIooT8BjJUAetQSVgWIRYJ9Z1U3dtqcXJGOJnQvgDrky
lrw5ffRreBTLbeXQxVASn/nGi1bVY0DrWz5C/n99q6KGnEv8oThcBSpARPwMiCk1
xsL1BIw3SOy75XOyFTvncgvewIoUfpPBI1iGdJnFmmrnWJdfFK/b/ouwqIQRf5fp
3W9iVdKl32hXMPiezkctZjN8nWTrwKRufV33TPBjVwGvEd56BpMcDODvo+w9K4ub
bdq6f6MFbsNkYN4nTtSuJVAN7hgOIGb4fg2piR9dbw384FD+ixMGh6EicM/MuPpy
hTTivlI5uaDJ7fDHmsbHbGPP+skSWzOAO79Fn7qSubbdVp2WJX2+frg5Fwk41ZSp
LRgOqCjYFOvhAtoX/lqWZC/rm0aYtjqU/an2oYm7EQT6bqVh+/TnNHyPZKzMbxuV
FVWN8X/NfF0zeoaab/sUVqIdUsaQUoLo9Fc3dR6hPJNiT/j9OS70ZpQi+zqww+dU
UfIOQJDVkbSuSGgPS6rDtTRgGd9Lu7mp07lyLhmIiem+1y321OpbU+2cNonxEj04
heUpaHzitvj+PjRXMLK2Ml1tEyE2/budJgDrtNapRFFiV7bMRTTG5M1UxjJVoBA6
FHazf6puAppWlPh6jMa5rsleAsHY9eaJGW3zszgnbk3gBhq5EGs4Vj3Rc5XJbp6p
dgKNd/At/TNTWOfYoCfehnwgNT+udzsmp0Mr7oogrpKLyrHwF2OqbrZO0pggTzQm
t0evj5jUcbd0c85j8x7TS/RYu+liA/ut6dxgACSO6KFk50grxwoiaa5GbZojBDeg
jO2K0QMKHdwqvqDFay/j4EEdA9okuNtyswS8B+NQzuw2GV603BcqW0dRGdDj8Y6/
oKHa/0FbCafmBI2hm24GevLDbbuCSOyFtnRBW20qsTjQ2p6tNAC0CnndUQxIxJAy
wir/tTE8I5WO4bAgxWNYparPMAZeHK96dPHM9sYtRdiNHi+nA3aaz5/Bg0HWhrrv
PEJv0Z2nh7oqTNzrhkJrVlLSAV6saQP89MnyTZ1/66yy5ZQppZuanUrVXJVhrsXX
Z6vPyf/tNV+d4AYR9cEK5FNXnP9bMSlUrHPOm3oh98/oictRfyONWtkENJMlzBQd
BDlbly33cgtC4BDD6Y+ZsQ==
`protect END_PROTECTED
