`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TMfukzsOL7F1YGgKdoBlDsxteFA/m8YFy2Qg4Cqh87ehcmGuR68OzWgB8+LtPFLS
UtfLA8thX9kJLvwwIhEAgX7KxiCdCwvAX2Oy9VaMjlpJuOT7WjM06AqoIfdpKz6V
92TMs5GzcfiJXADkx+tQLnidOYZWiH6gb7aYU10CkuENu5I4vX0QLzpexss3ShrB
OEW+JoeEsLmV57oi56A6nydcFtgNFEepJwnYsQJJ64PNgQHzn7hw3l35F6s/mQCQ
xUybBjuglEgoC2IWZE3iYWG8k+f3BbXsSOPENQwQTndOEbEmhe2ZOZWtszk9GstU
xzyPug0A1otIEuk2jpPQes9/Xe05P78S3NzTDYcczuMWl0mFhbbGNzj79gVggIxU
qRfI26CS+Z+p6QIxrPj874jys3NBBC/hMahU3YeL74sqrQPXkzevLLnvYXfLvKIP
kfnm/n0RHnxGjoXTweIRZSbMias2gNKz+SQgyuTAq29H59eg9Eb4ZqjwECDlFmjb
m6qPuwemhaWygIHEoRBdn6XK7jeoyXUVyW4Vba6OS8fM5I4cmYmqwGa8XTD+og2F
1lvyzxOmxkU9qnLCdujMfJOgCGiVh+297LI31P1Np8/mcXwKylEfIOIshOfVy6Oy
NlL4iiEI0y8WZ1If3N34B0J8zJBTmaLzn9flJ1Ny71m1nb2YFF49jrNwxcQLSIv0
kBA6jh2U+ClRhVlK6nqPSX6Uiajb5QzgmLHJrLgUufuBxWiD2h6A5h3Hs6K2Fexb
zU9e4EfVBkEKxhBACgZ9SqUmGZSDUQX2F1q+cjfImwVMoeQF7+zichp2VHdcuhgu
z2H22RgL7E7xZlZfnu7SLLo72dzqb6l0LSGgBA0xcVxPzrV8pD275yMlUSUnntcy
j9eV1JzoBc7Qkp13xCHzIhN88+bOjWktdYutmlG2C2OTl1ddctCmsnzrl7hGx/b1
9Nbj9bSKi77CKeNbufumWAYTzYatHHZBMXmru5GoR/3URGAEGS1tziI49NzV267k
umiHIomisxPKF1HrXOhj9we06n/u4xBHYxUcxNAN1rHFRmrg/nTnwh/gbO+JAkwI
PCyRfqu2SkEm04n92X4Hd3Aj3wY0SrFdx+uTi2SKOjWhwPbKl8F9syIc3zsUEHh4
88tbPmdk6EWn6JGpOufR/9wM+lLxmZ788oqubzEstuCkef2dOlKlMnzXZ8puqKvm
1+gig0R/Gz5nUbkNS+2JWmT3UzZ7dIPD501zGVwDXfWqQnak4S2NtNlqD42Q9oj8
s4T6FlxhiOJRumc7QAXc9sW5Z0O28QpMcTGhgcWbQKgxGGqcdDguf9Owur2M4bdO
WAdSuNYvS+dRzOTOI+Fdgbtx0govdbrUH/euT3+bJDVnl61LYrDVYeWLzQWTkVlY
vjQvl9vPrKHC5a7skdtZcJtl06tpj2Gk8T8U4kPwFmY=
`protect END_PROTECTED
