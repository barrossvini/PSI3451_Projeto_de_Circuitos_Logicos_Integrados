`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1TRxljxU0/uSm0vfT9M9xQtJmcQGX6tWbRwYIxGjWIQAkymySdKLRRfrdYwPsJHS
HNVRJR/AmFRmShZjKWI87pC5SVCYbvhSw6zUaXGK6l3BsDAenexpcjv+LgQR5BkB
Xlrazm0HG6qtRvWHmArl2TtHCmjurHJ/JisXYN9T7rhy7kLvjBp2uOOGavETo3LK
udErjE6u/oqY9aFz0AiG4h5lQh5LHKBEUDQ+FeWiic96l9z12WQ5xvDtv3Y4BP+k
IQ/4xQx6JCtshia1zSbP3oNODoo+A486jYPk2xFycrACbOJ/O1bZKzLG9QIX5wWI
BNnJZLKzANS6asEs75zT+3jXCSOJlaxkPNDjV7ihyyfGmoaYwGejZuiB8NrDWfzG
nJmfRpIFDY0fVX96j/wKwCR3vxIxmnFXCUaodbeScfUY0wK9VpiZWEqIag4F12Y0
PrFa7x0+MV6XAF2fQAFavuUNkYUtt9phJsJbDEEhgG4lcBlqtPc/sG68IjKtqTGs
GIHkzuSg5o6/C6FVCh7Gi2v/PmKUK2TtP/sxumOPCMrx58l1uFg2ICOlfybJEoTx
IpzGCWnOqHjvHTEFgyYuheGlOjS17Pggk/IMcNfeLsYT0P3NWAdpjhrMnL1A0Uz3
SPTJmaJmKM7IRN3kmK6HcWJHy+OBBhfAtkjvxQPKW1wmAuUBJRepibVy1qwn4LPj
hw4Nq8M427h6sN4jIW40bLYLM6yGYehAg28ZgCmbplsxgcxmeajdddQGhfUs2vDo
62f0AaCbe7LtnbEAO4PmZkIiosKTcyfKwpMKJgjmim3GAdichm3X7I5/NGhoN32o
8vhCPhi5WEa5vcBh2oasJsFWKjE7L/+8wOoLQ0UX1mchi2U1xAQhfx6I6Gkypub+
vcTaSXYAi+vYCZQgiDDTljPZj+jxlcu9rRxJaZyZgdJatZnFs3CvTKLnq03Nh7Y2
CKB2HLBrIegC1Jn8czRvRq0VyjxoznmOlT8SgA1gqpHIumu8Uf05qk/d7Hkk2DAp
N/4HGEphylmXkkrEA+Xz5rbMCO1JPOpA1OBOq5xJ4b91IjUyqhNhTLjabMvEM4uN
pA6G3+G1+iEZyIKu6dZAYYuEJxLrYPmY90hwrP12Uaba6mNqPC6DCpH9P6cTdlOn
q1eKA/eC6V5GVPXZHnh38Y/Sj4UYN5abRBbtoN+m0QLia6HGqie6IIiNtE2ZqvBR
qISzv6AgQO6M4WKLH2Klb2667lA7KcDk/pVem5J2ML1mW8VARn61++TpDgdQ6t3o
C1niSHfLJktCjifOzQE5fBt3OKS19Ez+8X+wUo67XEHcHlW3Nl7PjbCjGx8dDaf4
CELwAyCLqPJ9lUMz9CNsjSAYWMBHpTqwDyiLXDFGx2nAcJynCUIj41K4+ykJEL8x
L+ldBB5XY78a52OWE4y43jY9/d2wfgCT+3fGfn8tvQFsFlPLWqRtRjOfVKja3XxY
vwdDcjRijswCxEvfI0efR4lbHf9+gOKP8Kus+v5oKfc7AO8TRMXk1eVZi38Kw8uj
e9TAw0ctoswXD/yOtze5jCyKww3G6KZ7Ui0j3l8ry2e4vgnnfBo7rt0bZlNLudxX
k421R5ujuTS8DOAOmWx1ljFenjmmf7yfSEEUE8v6FnVfzpLY7fn0DCQjM2R5XbX+
cvAEIO0cQDT/XU3m4D/IkB1OK7r2kzNW15gOVddy5Tb3kPc4QC5jwrP/TVAI+tth
l20Hu2bxLpm5c8jrH8er1ZHpktNc0AWI75/FhM/hFvvH0cvknt0gOrS8bNQwJR9n
sHBYlNvPVkHi4O/NzCP1PVRbanjCEWdRLvrJJGLs63Y6fRZp6McS0uBu3/BjOQSP
rsKMufhBK2gnUeEnRUEbBGfVoA64ZJrOrrN5XhJP/ehZIov4/4qBIgjx9lCmgS8j
r3CxurQqFOIUsAtUh0FXNM8pw7xIhmQeRWdprxa3eWuv9LA7GYl77XbDCagM62ou
keRAWHaCsirqPfEGYYDfd5rbfI99TMz0wuT4btD+/raUJHPp9VGmyWwUwGEibbAo
5COWsfxbo2eezo+5GnzvQ0m5Z9J/y9ZTjkXt6Lhqa2sTJTwTOtB0UnfXecggpvhV
I+T6LKr5uZNwQmWwgyiRzL799Are4lPnqS6s9A+riJelwuWWklabs91GYZb+GFsK
om7qXVaPCKejZZ8B1eJEan+BUvOcsz/HtPvpJAaoYldShKLMBKYliyGAVf11tUso
Vv8lOUfdlSMGVGqpXriV6E7aKi06UI8aK0/XD+wztucKV55L/c+ovGN/Y0mI+USk
bGR0KUGiTue9nYXzWASr+jGC0qIYDX0nhHwXDR5iWocHCz+byKyROAoBehQj6Efa
HNbBAL9S8NAKTIWK+2tXcx1vo+cdIqfgsABFi+8aalaFnLPtG5MRlvRy+ufT3e4r
EXi4LrR2LelSlgWBoeM3jON9VmEAdRA6smv4IdMd0XqNNjdoXOlr3kOvsU1Jyov6
4/idRL8bsarlfJuOOZQta48of+qiKOS5WmL9JC+l1A2pGYZWN4OmvMcfgGzMTn7j
yA2c2lwMO+F6CzZW54gC4sL5PVXXdNEeVrxCc86zgvzkvVq4p84pj4TGEdgydYOd
BDZuCDggWcmqouOK/dmgzeOnd/DV9NyOYJ1KwvywdS9CdJUnXCTItSp8CLhdsjL9
YeRGY2Bm5dr7bnL+ZcqWvWdEJ6urd46DM+xDiYh5Sow8rO2JZaeAIK3LKWtaopEm
joyVWF51g1P3b082hB9gUXn68tmkYunbJIMbsJi779SD/I/FoM6L9fc6R4NQQrxK
WvqBl8cmAnAxTm5zM7kJud2XQPAehGwAE0XJbkyN328zTGdDBa5v6Nzsfy4cpdDI
rPRg40KVrXRjeIHMVFn+cawQ/eb3TBZIEeJPyt4F/DInar5zyVU2PDgouuUEUoqa
82o0WwDemfglez4qbYmgiznRZFnES+m7lcNI94dFhpW0hWDJM6G5nQCuHlMi0Qwe
RhhKagl82g7XovRoXfpNd7Gl7YLt0/Qt6ovaSL74WVMJgQTyN89CC0a6wG9+EpnD
TGLb66GyfTkJqNu8UkirywbRbn4uJ4cOAoIEPNkCH1Ekj330KDQVPMr0xSTDRjHi
nrZL19L11ypdwmR/sBXHK/O2CMBWGySqzXKlPQwf38V27rLcR9JtUb4/goTRXyUS
XYnWhDIEYutoTTg7gduTFUIE2B5xbuqVFbR8zzrdyReE3zILzMK2Jse6h0lR15ub
ZCouTg5I4PpD1UbypRbCa/NnwAP6rWq2om6rh4gUnbgBgksJT7bhk45IJfLiluPd
orfKuqFgBQG6E/BA43pGqywYDrS9FKrRpUlBtY9ZaM6IbV7Ki+LG4BKCwM+Cirny
gmyv1zbpgMFBgSKpLr3rhwKYH7b+4/0kfoZur5zvgJnHfhOWViq9nFtwpnHgkKR2
1xreflhoDQF4j5G423Q7Qeb01AqrO4mK1MGAkmXwW99hluvRK1oQMsIuYEIsZ0O3
X5niUf2d8PWyGTnVN6/UWCErAfli+4UVKzy4HJNyCLS9ByuaqIgVNyXJ60Oj7SiG
W8Vb1aqEHCx5VVnpVDD4fA8seocpt+/vLusoBT3oZvdXO+nVYe9R0lddCJJzbqih
AvTFtles0yRO8hnxGjWMKWL+La54A9xvQ2BguOshaHooKgPtrcU0FPYrtBQmhK3I
rpyivSUam2kKotrpIm3G93tGvEYPYr7dwo5yTp1XEyEsLIDDSyR3QJUXoYZj/GQu
ydja5p1/JnnsLKupgz3nRlK4zax2t2Aw/w8edFQ33hnI/t8I7WLKWcw4pgZTJbt/
VNiVZ8zEFok/Tp022+AbRcxepiQ4gWeSElsEChVnGJCDJcmdu84MtgKx1S5NxFGP
F/DaAHKINBAde1cmPb1YUPM262F6iz43iAr6ooe2Td6QXvi7epcTqgPmpgjng2QN
TYHtM8tPEbvO+1nT5AJevIE5GrSb4aGYhU6SJfZDJ3EpUMzQnOTSuk3kWNoe1bi3
vplSOIqOZFNhxi+71Sm58fMnVhMIlIodH8IfkiylH5IvwLjHI+EjUQ+G8y0vuCHL
fBFRte5KD9yQ5AsUP5rvdSJZ29RiIKda88MYse3K1e36fRXYm1/QVmeXvyk9+gNZ
Lag1f2UZDn9avYUKjKiBvtVqNUnA15uxGdyAjm98mMiVXIadX9vim3HFvJaN4Ve6
Gbe8iPqz3hCyhCWbIoLiy7KcfbcNC3daEzG21vgLrFJVjzRo9bJIdit3JKY0DbYQ
CKFmA1bdrNwmj/+xxy7QFW5s9L39+SXMPjx6ybLST5kbxecHOXhE0Y41k7GG495I
9HpEZF62oDY0gFPMoLATskIdG+VbQXDQH3pLZduKGyFBy7r0pOs0fBQWHyALNfWC
r88Jj4mJ6JmyR3sCz0YtIujmz17PGu8u4NWLFutBKKk4BQRyIgBhHIb9s8ZrVbDQ
BWzoLXrrmnQHLztqb8MFnYui6QIk5mHDQ1fRhvfpx3iom4YYOvDMc9t5VbRmOHJs
7QWXjlBsT6fSgmeA5dSDDsoDKsC5cmv1ByJP+o5LyRve/idEXHXgV9y1CZcYeR7B
daPQLmUB+pg5TYfOFpkyUUindvntc4hLbpfenQ0IMh3udmC+mtMmgbOFd2L348P5
/zx1ARNgJfOz0iTzk1a/IHT5TGDZsiAHJlWzpz/eQ2VnYRc6d8yB653HOG7RsOBc
gqFkYoOIoPPOaDZfQxuSF7kE4CyPoTiEyQMaGIEbDZQV8nn6/Z/lX+YcN7oyA0GN
mn/rKjYzz4Mq9slU1ng/odxuqCrVjXYC2ReZFZeiK7hsLlfnhlQHKah4mT/LSQqD
yPlYixTjqDvb+HnMoTSBcnYEtv0FAJBIhb7o1N+oKIBy9W/Igq6p+o5GcnjGTYFC
pQZHpLvYfKj/I0p7bgyu9BgVGumGfIgrNT7b8YS7Di0cCkgJgJ4++VCQ/FF9Pryt
AYL+DXkww4cnXyiCaXcrba8b1Dv3EBiEWwyfVJiTl6G0vJxyhbTPsIqgIKaRo0JM
HSaZGiKD1xxW9uWbCVM5AfBiKP79Uy0NodvGxRcyOrbFwA21wyVLYHPDL0xIgSzH
MioLYVN1ugeV9RsBhEIq2PlLSk3Nc7Lp2Tn+eM5SJ0iikE9gl1/2DTPbD9KlzY+k
B2WoqIURxE0eDi/k84E/lFmTLsbt0UDLD6MZSMYXdpbzSM5hXM7dORgLxQE5WTny
HggkIzUCWDLx1Y2qvUQ3yhwnpU5jAkiFUj9Nmd/TO/TGjfCCSpOhgcTJ4fAyS6Fn
`protect END_PROTECTED
