`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ufkUWohWQV3rI/vR6YbgxsI4HMDhcOJlaPA05fkCjnyhdTm+hVSLbiD8+chmwppO
4F8q6DYZMrU//8m+qdO8HvCDjIR4kIHWiMgNDAI6AnAmDBPgJ2XTLXWARuOZHf7J
1Pgv7EuwO/tPUXboWGWiOTDGVde14BE+uY5M/YFnks7zZK0lZBW4kp0p5KfVegTR
LPsnEJyoyM5WLhv9FlfL6gF4jBQ+m3LQGa5SjYJq6S0T3mBulr7qlkwo65DThXJv
Hx7rxQy8MIAn6zPjpY/qkI+3NuRyLXN+rlIfskIFXzkqysDvsVPoKrNZ3UZogxzd
h2sFU8kfrG+kG/z4cTMTaFLdqXcXPo0AxUZDU+XAX9TaQwqmmgJiEYo7dOIKhlLJ
7afnRlFyYa2VmXoMgRJgD5R5BtqjwZOyhwlmR5I0cPNj12xsg/A2PuaeRrH9Wv23
Ig9uwRBj2vgVmFQr4mwUytvtOMScsc3ZodoyaGog4QKePbwpyaAQ7r4pzXSWu/gN
tfTTuPd60ac+JHtxXuSsPx9VWvXKBUwaHv2Lz/xw7vtKfDTx6cnSUtBpI1Q2L5gg
EiLX335GdJ2gGI+XNUJ21QX8aJFPu1mwFNG1v51W6+H20PiutbqmxnfJVlFY8YHN
4QBCCYKMOrreOI3fDk2ejNmQS2BR5nnW58RuC3n/qx/nOokfOJeRqwlPzK0zUodE
UwYVdOn93b4jmfjhbGE8BNP9Kh98UEqxcdXbcugMq4wZEJUIYt8kUtjGKSIbIQDo
Mvi7urw5KD/M/+GwHHAo3UoQ6pcCEIFuVznM0denI4zx86rHl7bLkzpJImOJGH93
BXWXYacQviTdTGqBNqKFAwTXg1BUn1m1qgYXgNAbcaGI0gel7vCtnO1BxpkcJJsE
QQW2M68ubcDl7xWor7mA5WCKtvJjOvDOf/gRazLco05+raMw1EdzDozyFaznd/OC
mZTcjqhQtlVxriv5AtRe98YkmKP5IsvMSo5Y9oLl/f+X0ick/g4LEUw9VBEWd8Qg
ke/H4eCm9GbTnxW6GOTYLUqoteXdp/LSJYj06wUjQoGYofHxa7x929t1zpT9sgrd
jKIsMJbGcsVEPZqlPuyThmKrMMXwhd65C1UlCMHmIjV2+Srg/KLOpnwFbwv7rOm1
EEu7TV/ahpyqH5lWF4Z3NpCARSf+3OiRRpvaJzZ0AThwqVfmMvgXby6D/VS2VE6m
/gm+49wKbpuE7AUvvLa96E7ajNWS96YMqcJxtn3RCGyBXD53B13mcC3wSxPd+kcx
YDREEy/xEofkCg6G4GKrlR7X6ALKnG5pXeHIGyBnFIfWu70mL7r9NevhiwKACyaW
hENfTxOuLDo1MeF5jtga3gH+SHdsjrNFQRW3ySSZvs48hn1DTAM+ISrKmS0eu6+z
5VKLoZQOxs/ofAFj5UKs3mIcIOUSbnUAaEvWHBfE7eCjx2ZP1yFK71nhcMW/a7mf
+7KLqmjtpWKtEqnvLwjurrmXvwgmc730EeAwRg+dINnPthJZSu3VETlFHMyxicBC
XgDYrE1i+xz+SRz14Qc7vpuTie0JiUJ0H8wRCuITy9KbE9qa9UJRK6WxlTmlwYXH
5iROxtAwifB6PnLJDJsCYXXY9lAmV6H0zyAm/1eAPWYxhsqQtDp8SXnpRxuBBuYV
/A5RFnaoFDahFdbgU19dJRYA5OpwqOVnviR5ZZqkDmrGQZZG3tS8mOp/5LQkbvTC
vs0dCxCjx6A8tz6nyIoofm28ldjKahhSzP6oficeJM19UjP3BzF+IgHcXo8rDZ7u
`protect END_PROTECTED
