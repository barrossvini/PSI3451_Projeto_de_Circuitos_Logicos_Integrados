`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qSNtjv+Va6SYiFI7EnJfegst57om2ijJyfE2nTUprZfHQdqsJh5PDg8YxvX/qhrD
Msrv38oo/Srk6r0k2tVNqy7fOfjXdItISqWhASrPFyjrfr8C/+NwaciO0O12Z7Zc
flV8AlSqcI9g39TWrjtLXKDDhfiRYXuyFYKSqiBqJOYEi/373v5XSJ625f3T7UsS
n1qOTgc0LGfmVRy6NTh3YVGK12y0zCn8UrM8qfrywjDnvCWB7wxXGC8w5otp7sil
sJv5VODAH1lgI/5MNsNTsRJGUqi3vRZsWaUQwVsgY0UPZYOzRfWbZNDRpWjlcyyv
MkUC54JRO0BSwalWg49wpxIOcSqtspDE6qd9lZB+JlLNSOcbsg4lZS92Ml9X5Gvj
0mcoEHEQ/y+jW7o9EtJf1bFZHx1ln1NUrJa1eH2nXzro/fgz3YYxMWecB97lw+z7
0qVWszwy2PkUp98LcYGPBbfFNvratqE4LaO0kdKueSB8/67jHS4/swyd2SrZUAEV
UO0na7pITDq9mF74L2z14xMy1ScfjjaKkGW1nkir/9cAfCmr8Y2PDPmW5gof/hZ3
Ee8Vn+QR829f92SU953ZGx61X9yJYa27Y63QWMZhnnGa/7zFfGxiMB5KEB0ALrY3
3FyEvxiI2cXEYMiT1lPrsyUGNHdyfAQ1oDFwm4eCGyt/5x1dKwMZBupA1dbO3FF8
tJOMo/DnhDPdutZ5GDIPapQhDIsocevs6ycUkXIm/b3XCc2ZL9que7UFi+Mqwylm
s1cTz5nx5tqfFhiXpO3rc31cs75ut/ex9RTpVSCaMqxsgJ9O/tE0PvG51JrfSo8m
91c+3Eg6AH8OQ6f4avI7bByBSSKgi9e9vo1PWFPZUF0SWw9hpf67AgRzocWCpZsD
ErDwZZWMPfxVQnaBVXYC32mSH+0aQ+70WpBD3rPEl6Q=
`protect END_PROTECTED
