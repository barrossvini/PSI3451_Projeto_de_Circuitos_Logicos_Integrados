`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nb+2+ZIf3/d7POK4UjOdnNse2w4UsK0ygRYvc5EWlhaymSnnp1HIosjkzKcIeElw
GW6AOACgrfFLbqDSsYQZHTxeb/DI9IeTAAgQvo+hDJ959RNEUZ0GSN3suH2R9DKm
5wFnKguWL/UDoR/RJljQL+fLMihbBICWT35FJReQGeUnlu823hovb5q7uSbjeIOC
AdghTDRwppBR8TDWC3jYRpxFNZZI+WflXCyOT5tR0UtHZfw/JJ4lO6s3/3JwfyBi
e8hBEfWOnivwlbti4iDjpxxOmWZQOguvQD71JrhgrdK+WFVoX49beJKmqfwiKigr
RCiFSJMCcMumjtsIL4iUnoB7s4dvQRkK0Ca1HBACN8S1d8Eaf9U7KnE631RDpnBH
Sgqk3kMt6XsMQb+dncPf3K0IUzVCRMd5ZZQhhcTfN05WnNPgy/CgSXjIBMK8Qxmf
ND3BQ4zrU4Hj3EJyjSsD/VBSs4+qxa4KqTQxlZklmnb8bj3+6KUBWY0M+sxonA4U
Mp6b3eRXQB15iD0cc7ZoR3FvVQlZIKqWJPs2/ePkjiFFKFC800lpqmjyCNUu7Nc1
uO+iwwuqTUIVlEk/OWufpOp9Qy6pxF9wSaDxyd26HT7niEbhBN7zVHrGQjGRQrqm
tpkpCymqgeK4zO379x/gXEKcPkUR+agv9HymbV6C03trXO5QY9ybxaYEoRFGdKQZ
Jqj1E6PZqza8P5VP0T7OPKXFJ+wnMeViZohrpNcBouWS982homdv2yzxr9JsBvTn
sajuMi0AsytdqEnTECGty6u5M3Bc4f9wQXDsqdFp4Oh44TMbN6x/QMfZnuH0Qcua
AYJ0IYhMfiN5cQI9AzGeZMMRH7lKVISQ+CjG7hSByfnGqINN31F5n92GrQz9yUIx
noNNjO3Kh2g4DDQl6/hc/zYys1OzcPSeNoV5StlrhC7AoHq1WTOE8JzfPoAbcK6h
BxyECZp/mykdumTZetAFoem5vTom3qMy2sS8vYH0wjDrBKS76DPDljozZQeACG5q
VVxVBJ3N5M5g20diKY2QEyNJmY6IUT4SzIinjJkT7JXZB6YEsM1eAA2CUS8+eBjb
0mDWDziCeIKxqGVurjhLHIoGjIlKVWIz5cQTmZxdf+INtMEnEEwGy81mnKUlVr/t
S2E+4G4djHMZQxOeknif7ejdVHHfwv8B+jrORBth5wHspVCCcMh/k4wPa1u0yHP3
nqD/O9bHYsK4wWSkHYfJUvm6RdgMbD6kNdM2y6aZE3BJMwZ/XIEpo5MQO0sn32Z7
Y/C+5kEXtU1PAe+CRviI89Qem3CgBJ14E2FKYBhXiKGTh80p0xAmpyV8eBBgXzzx
jQwvzeDPOaR+8OpbZhcYx3uZIAnn+97S3Q32ufXtnYPJA5CytpRnHXpWwamLFbxw
krfJlyGFREODqLOS7132P1G5xqpU9OBZDvc9YSK/GBAzxi9A4k61P4r64d3jcKqN
lT4lRu51j/TETeZre09nHNVrQyT91l6EqVo9glMTd51VDhvuJkV/dpnQGUqfye2C
lb2LvYRRt8vuCu3hFACv+A==
`protect END_PROTECTED
