`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5M6lmIMkHSepr2EYPm1ccAoP+WCyucCqel7I9spehumi6WmwHMpYTHI3Z5C6Cnar
UVapMHbKliORXhdMbOgfmhGXJyl+ebZakKLFnefHiWByZsy6VlUKoth1EzpQ2raX
5aZCxQ0l2mZQnya/lpm3rvrkZPoEs8965nfCeUfDgJaO94QPri6djUdkC0QuqrNj
w9e/AKMrimjfvvuVEayfHDuwBnbxLdM85c8vMJYwg/QogoToGcJIUE4Gsm9nn/H4
In3RSyM0xgUAeqImNZQ+kX+qJnt5m5G7J+zwYkVS0mIZF+A/YWocqAHYnuuNqn6p
uU/y54HAA/VD9qjVzsE3M8wT9dvl2FnMY5A+jogpMNT8vjgq41x8W12FuI4h407e
IlCiWLGlMI+kSNsYzU3ZKhuyvhd2GAz4VdSreEhrZ4YLh1d74y7IEGkqP+TACxxD
Gu6AUpk4NiavscltXr2yTtSrS7sR29LuYq/NRu1yHD/nvDjn8S0y+GYoDU801rKZ
FtO+ISEsnYkbuM65XgrkMJsHH6IEWUEUn4jvJAxjy9C4EFs/aZApTslHddPyUbFf
KNw7uA2Iexru94sYvTA4xFfZlEC8UauOvK1/WfygyGd62oOX41xD7otHtADxJBb/
Bn3l9BQc9QNWhXsnh9VLtLfxuu6gthIze5VybevjK8uhf3sCplUwbmMGEgnjkCgS
QKYLHEnl+g1R5EVNvLeUzbAdgyDQeHTWyx0ITDswM0hhJsvb+qkSJlS/CUkZoOUC
qsspdXfQMBdo4peTtIyTTL5sDp0luxIcso0bHmtLmn84nRzRDKZXHebUY1r6hkEb
JiVMoJLHFVXj3qw+b2Ojp0rryWwi8kDN8e1/iSlOFf0+E6AAPFBTgE/a7vjlB6Ru
WVg+4zNzWBxAgGM0c8YX9JLxvLVyd4U4SZd4yli1Gd6bH243WrXg8MiBPFlafm/l
A1yxjvuG2ls0a6qVPEAiCeA/sQUUF+f4Vrt4dZnJPCujjUUEcf85L4Zx/opsCvvC
n0PCKjCxL+4qPMo0Rxwwchbgm9weA+yjhtZR8LjvII6fyWwKASNtqB9raJvfiDlN
C+rIwWtVbaommKPTFk7M4OxsqHBGuOXcJEo80OR+ZwuwtCS+pkJ03tWsXYYZ5jyK
7CQImbD7wRAFMyeBKrkJakE2yx6UXj1/j0NdoRNWNI6QqzhECvWwY8yoGayZ0UP/
Fe+unvZcyWEwimq4wKCEcYdeAXUGl0NMq+Hne2U1RO5POjv12RBEDAW1rpB0ZOkE
K6md8rfMUFYvvO05rdoWPJtEfgYjNRzXzEQbBzr4WeoXD8MP0SWBk4HZ87Qao1o3
25CXIJzeFqKyfNa04xMh5SYS3ziy6/lrGtC33Wj0xHJjT+pFjY1EcbSVqrSrgiJW
0UmAhusQdOVfPHygjn0DwhK60N4u+t77WP5pZlXH7XilNJ2KqYjgM6Dp5djNvJaI
q5413DAx8Ge72to59gdvBcGwyDHuDWqtusH1pGalm00ymya6CddUkR1R0EpyenBT
8AV+Ke17auSxktGErf65DtlWwq1OWLYsCW96310cDzLwLGGeKkGszWuPW/4GbfUi
AjbmYhoK+2LE3Wsn0SLe3ajU1BNkG010ysWdD59ofVt5vDvj5121x+arh3vu7JGI
RKTh4UFh99tvrgsmcipzH3aVwsxAvxQ+lbE/0lOm4LnxCp+njGk5qI+hx1Hv9YMB
0/RJA8LbiIY6/fYDevfcgxcI4hqzKvvdyuZwDmKLSH7SmADicYIi0Sksybm2pvaF
l+MHveCHwNsXVsFdyqu3pJ4l4wiqhJyIIDJz9xMK82NO7z/ctv2AF46UW88GkzCm
y32OEZvIG9i0sm9dFHsR2QTMl2Qb5f6Gv4XwopPi1GK5RHFCrza+gQl2ot3quEb1
fLtDeN5pzuZIqOOeeEPhOi8kmMAEX07tCHQbANg8hz8b2anSBgZIVXHjbDRYB45+
WSclMuX3jGCQWPlMdADDW20/HFPTi3I0fOj876Hfkd3eqz5IdkYDUxYG27vCw9MI
kslss2yHvsebuuT3yF/nErgStuY1uaxpQGBmwCKDL3oY1Dbc50WrALvgkNfYW+4Z
eBFV4V6V0dACYP3/FdsskIq8vMecxQSKMt4e7wiQU2exxmFuEy47/NcVFkM2sY4Y
qwZQZdfSWEIiE+/bFe6gXwi3YwWfrnymT6etRi5tHLmG3qO4V43ML4CirovzAyYk
gwQlUdIj7akJJBCExNT7C5HeRCxoOX8S11V+yqk0s/X9T0WZNuTjWVmlKB7MGaLH
kjrdAbdY6nchZpkFgCqf76VwtB3+GMXjb4TFFOL3lBCNsNLqgxGqGn5DOmlG9URa
Mk5TUTLiA0r4Fw+GhagsmESD2sEWb1mGlrffXlaFD41vHfAueo2/joOGVLTlMvoB
lgGy12kzdU4LS3cunCksCU/RicRJ+ZU/ar3iKJcair9Vj4QveqdJS1ySKSRyy6EJ
seT2otQHrMXSRyWs7S8EflefiX3CAYZFZFby0rSsP2kTwqVyHz7SJf5TKgnBAnji
xO6p596Q7Di/xEdbRQCK1cWYE5aT4MsYjWuRn4Yh0Z3qmHCKz1bZAIHw3TBtTYth
+QpeapooI050MyBqh5XVdl9UH1huRiEHNv57mkeotdvyCBNUn91H4IVsZ2RJp6Fe
vC2N9DweVGq7u1ETCJ2lB1YfWzEACc9Rxarf85KXwKCj9eSVuaTNdIJF5Yw778zT
DJ1pAqMMgheoVJH3aRpc5w1KcTz0sAEXSZTYfGItjIl6XVP7CopGzenfhZbMCKdD
Diyxr3YC3/Ku3UaMU8JyJL+zSqaEV3s6hCJWewSvzEM=
`protect END_PROTECTED
