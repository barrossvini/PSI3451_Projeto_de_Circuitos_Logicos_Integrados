`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
29AgIdDm2IPetPK6sSIui54jzq9KsnKzl2PkGq/z10dea7m6io6Cx0g2T0MDj+Kp
Fg9Fma9NGiwIudXKRvATe3v0OWI/3FIVygVN6LNdiCgCE8ajddnzrromqLxiBfWy
6kn1+RQUbXZbTpZKUhJpw9uDmkTqlrdTQEJBQADoRny4TkzwiENYh4Vr5VNKcJba
r0dpYB6UPUhqovQFiZX2+1GeM5NZFID+teE3H+JjdhnNswT3JPoWEG20jIIQtExH
3mapSoh/OPKrjzqgbAUvEy6AAdw9k+GJSbkMwQGQR7Jih886xTo/wsjBCYl16WuT
IIv22H8YYoPYfa2fnMaJIGRViLJk1F/Yt8MGJsCi1Umm4cZ0hV784Gshmz6xwRUM
8oDzMgewMf8Tw/up8F+FgwlD3VFMQuAYIUFDfW8Q/gnPsWB9w7cAzPTc6ZZZ+MQz
LF9iAcpjnV1OVxJ4jQFQBUX8gM0wMGUPlMuGBChloWnS1KV530886sLp6H79jDg6
Lm8AXUkZhVspTFuhE0tAd7vjK1r/CGWcgJctfcpaeXGDQbCeU3twoZnbCkzBBPUH
LG+Na6bK+b89Ld8vcFIsNItlEH7k9nkUAcmr6Sn0iHhDd0ogRjwIsmvTReJhKbwR
OsVsRwMMcFlBPSmXRpF8jF6nUW+ksBqEEPKM6X3HNI+RvefvIu0qD1SRIgNv65KX
GL2zawe47J4SPKR2m+9mKBEF131PhzQUZQgW0SegSP0rDOdbx1WkRXut7WWZjI3Y
8FSnUbra2b3E1PIXf6eq/a+OLjT5CAF0cBqDNvNCyCtNIXj7ypguthyRn5gBnDMT
cxMkELrCX6hNtdcR2LkPnCEMk5ogWaLE1MkCAw+AsIVUv6L6IkcOGas6N7wbMy7f
Du6E8etuGq0qMAgtatkqachBuZ+pnI+myD9Kv/5ZKaIiuuKDixreDwfilIjV4qQb
0DKeT+X8V5Q6cQr/DzBVXl+3ppx/J10iaD/aVTxbqojm/fLr69XKUkeqfYDYmydQ
z7cTTQtLDU1VUC52qd6CDGTLA6DSqhTZrWKQ2EpiZUOwhdftcthbOuZdAeCLillF
CyPKFijZpNp12Pa5ogTN/E2sAPDhCRnzcyxfw/spj5rgkN+Cs/uhNj++BKJKdZQ2
hpUsjWd6uiaJ4nekQY0m9+EkHY9du5+abB1JeeC2ZKesUlhmf4SYzvSAIMAeFrE3
qLhWjTRk34b14Cfcks8nk4yt7Hm5x+AhgzQ2K77XC5dydzCmW51dCwRU628RmlSl
zy8PzQXJDX6o6GyjCZrzyf3UdmP0BXGmaMZx4Sx1lTO+IATFO58LdBjgbSpADbRe
hxnQ/7eGgAmnMy06tAz9veDyzR5K+GK0oauHC8kAMepruIiXyIrkL4SREbllYtqQ
b3W4ZgGrh26xNyBkLEIYnCa9+eaEBg7+7ZIVNndn3H2FSmNCIGug+txXAUeP0QWd
UMdTc2Y7QZUipTffE8c8PfStCH1MoTvFjbRBgHJhX/Znwbrf0PwWEAzyDqzC+qEa
`protect END_PROTECTED
