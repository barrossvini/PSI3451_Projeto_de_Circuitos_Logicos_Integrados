`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5oESTkZKcoOADyaKyey4zZzBU1SqbKsEThH/QID71Es+IMYbOnN01Ifs9fTaV5sv
r2Y/eWidLZ6QlNRfnpuEebUHIuCEKjij1CXCV0Yvgu1CnbjWUB+0JDw2aitYBx0N
/UDXckndkE9P/82MeX5moMwqEqQlOvQw22MZ22Ntxf7NRh2vlINnG5XfIE4yc1BS
LfmRDtWgYiNskgi4cdrr7ZEF1pliWuKfkjA5sBydOmscXqIZ0TaD0zDIYOfsL+dy
qeYRd4zfFyEe/iLiDgZOgov54sWD0jrIgHluWH68r1EtbhxfYPsz02q6o+T3fTmP
Q+iJ+wpbbZmReJUim55Vxdp63Sa821b8VDjnQ9iV/3FKDaoGAxIoQ2GMswNpa+Cj
00WK8Cpln6jJewziRmyfyDC9DILDhZ7TNKRqxcKmMi0kxtgPPhJJ3xygCnr5Vx87
MtXSDs+C4GrIOgafndo+gg==
`protect END_PROTECTED
