`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8FupD5uibe+QR4W/eKAqTeim/qysz/hzuxlw0rhh69PIi0A1gpsprrqtEkpn87go
MPAi+g3zj+ne3yWpiZgeyoEDXg/QkkrmcTORNrUgycKp5L0nUVtFGipJXS6+SWZz
rFhs4WCuqWkQ60PJfg/PSXRTFnbV1NQvMNNtsYDMAGrSRoAZKvGQ0oYZivRwC21M
9YzUxqIZiY1ihdK8t4qjVV8tS/YO2XMdndlCUGwaEnD0CMEmx0+AmCtbdqBvDhyi
tMxJq2kr8BESU57U7yqBGdeVwbqhfID4++9s7Vi4RqEy7cITpsdFDHCts6EroUWK
wvkQroncpdrBfKLI/86KYWGDjS46LKpz4+o59zpEIdZp3JA3Lqi20lSqGOmukFT9
+nJZvzGjLNUf7dl14Wx4oo6Gbf1jNMRGQLsjG89nKsAgjJQiwuLV8j19ZMkHbf59
gmh+RlxKwIP8x2bAo/8EyUuIqUHE/ZOni1MO5yZKuvWr9Xw8Lpni0VTqX18okpBA
ftaEtyLkIavA0e60U5RO/SyiZUgbs4KME8BIu5vmg7Bai/Ildhs05L/7xwA4Mnae
SR42HamdUihhYkcIa25fW+wuteb7RY4vWV5HMN5RYVE4dgSDtJl9mKJGPJ/36C0K
xi7YSILZCRjT9AoTZIJW/mAK+3dDZdx7jMzqOIYvnF8pw3hUDGaAmqnrnUbm+vFI
F7zBhx800DTwCRxnwmoONJFJulGXd4VnjQXt2NAuNFzcabgbcRVJgJO6MqAfd6GY
kYQXkwMHalkxyEZmOE9xd6pL1qTQGTM8YMADlioCdEjaEmnHEJlUb+8SYLe2PONG
n7xn62Cd1Dz6ccUc4nneDAEDzdnBlsxFYM6KXadut1NdhO1toR+hwLyHSure6u+O
h1JNWFnJlDW2t8qD1Pj35r8By3/Gm3c8/MbuQotWt54pkxKU3Iiak7OLVtB6iXtN
XTYjvDoElBOCPqXisNRuzn2aW+KRLls7/PUkMUlqTIF483oarkW25BZCwlDwEalZ
rzDOayqH5pSwXRrtARJUg6iCyIyOCq0gfRfQ9U+zhXxi7C8M0zrc7iUMf6/8Qsk1
E5kr9XT7389g84mGdIyqWsALX1rTpAwaMUddE10Jd7H4hxZq4Bbk2Lmea3JqTBOa
InC1DdnQLkTAQ5fC3KYIfuxGtvtkdzSv4/joBtcqyWzG2qg4lZjMdtHjXU3q/aV5
6O1rcso3qsI2v7+Ql5xyXO1gIsWN9ZK6BGp8oPTFQnhw2YNPY94g75tNQbLT5plV
HFFJWu/Htixs8Bz5jd8N3TqPhN+yarYV/zYSvoFo2S2rvFUfQr2d6GhzKz0Zg544
fwqXSYhX+Jl40SeeZE74pcbpPRGiRkCoP84xS0d4IXzDu3NmCXzySj2yRjuj8DWx
kqNss0kMHe8EJsMHOEquXY5JjRwBVqaC1PmYnokwh/FGMOa0+28qWrnsgHem+GtJ
kK6yWnNSjEVTKMytaNS4HQHthGkoY+fcw6e6KtT/dmMFy4HlI2rIQEdz8e0hRkka
w8c+cnaHUdoBcBit3VLKsQztwt+NxnlPpRCkrdu2YflqKFwI+V1BX2JdZPFrrVip
nJxzb4D/6Gcjuq+FeqvvjskB3bR6cKbP7tWTeObyxiq+9e6L3AWVq2/NVWyeMPx+
dn4lOAcdd77RaP7kwqkGusFUnXDjayu6Lw5zGESKYtpU5UIfVjxgQGOAI6GVg1MY
VDFwS16/EhmfWKuChMJxcW2YrDlgjAmjm2MBPswDEIX7WrVBB3p3LH0msGq9b0Vr
Vbc23FzywWrnVukgV11xG/dBQFXvMV7O3g+bMrl5yeC3fuGw1bJsNNwsSZaL4Dfb
CxftD3mN0VZPuGvR1dQdyArjh7c23jZqwzM6XOP9sl5QYAu5Nw4W+SKVbyXjeOZy
C1lszmTYnZf8UzmgkaqA6fhsGOiRxXvc76CV5YNbzIj85O+I1Psgyan3vDoEDLuq
SRgJ7/rSy1FLBHgMs3AvksUVyflURF+34lxHdTqYjXzmWVolGBNHd6/JY2GC0/7N
bGK2+SrhRiidmkzJ/9oQtVtbRofq6nzCIvApn0dl25qEQgRu6LH59tR8QcD81XEC
LJcFQj1tCPcusyaE2kAgk1zY90OoY3JF0BPhvz4bEgC+NuUbJ9lQIAh2lZs3HIdj
bnWyJxKD+NbKnMhFL76Vi2lfSF415xwSGBkfdzIC9OCrYyyhx43kGQFu+o5wnV8J
tXcbjHDssTEPi2VP1guKgdxnFrC2asxNRr9OSYG6ygzitaUPiofWK6ulxOBWBs93
F+zEqGZHKEmkQ/16Aq4Umq9Uab/JESauPWD2SEH33IRrJrYDsgSTwZ7ph9YMZc2x
XEkjXfKL5Hsr001QkBtV/InTUOi0l+EtNDjylRTY3347a8kEYtZA80f94q6dR2An
IhFykKMpb3tthAkDNOjmrKRSFfgUJocO7VLWn52NjuW1mkl/ZicCKvTHzlUGki9W
qVXauhya+bxvRhJtN7igv3QmdqRQUAODYye363JEgGG92B+CccV3/53D47pcaYbf
SRohXRsAh9yx2wx+YGQrk9tAR3R5HuswLCsWYwtAlntUTyxFONgywSYvJbFy496+
1ehqtPnUieaEGne8K3ZAKzUxuJ/0FBmpkswuqnzpFguC7QyaBOfbA9lqIFUtdBtw
7V6OiIri9O1g37sA7J+mj0ym1bQywkosxvdxumdtwWdX2MmCFUSLXovdpd7UnZaT
g/tXdgehXx+3oEt9UOlYNxEg8U2VTpWL3+I6mvhVEais38Ubcw+LjcvfQF06PmuD
VSVH8vpvYbKLNzLirqwleq6pofJPLtSXYOyDtVCvE/6AqZOR8kGskG2VHmaEisVD
yyZnBc1s1ZNVAkah63Y+L4phjEdMQltaEAV83tRuX1I9LmXcumknv+PUDpDig1q3
ym7iv0B2Sps/jDIKTmZZ1dil2YQP9/Dmz9KRoZ/+8fY8dLvz3kxVAVwbJzvIr/xM
uqhJRmnGV4m3laDHUVFPg+qexXDHWiVQi7GOgBxeL/5MuHjOZxsYynm9pRseQKP9
KshdC8Om4DI6hhrEQ1kJJ575007i6HmWesOjSo47vPKMqouKXXueKms882ysCtal
KUjhm/sTdkXcK4zBfVmVZPnYR+iVR5O5jJh55Vbo9MlCUqE9EbKazkL46r+0NasQ
+EaatZPgrxrOvuEvfqpvI/ZVYldTOrh83BbJPkkKC6effaCbaUcpSxVuSkm3tzvx
qnfuGQ+WeOmOkAagPY0YfLzglA0vXvPmPJr0OcGXmXTnBenLr3nhQKZYd/Fk6GWB
Kj+jYmsdegZIs98CPkCmkf81k2rLRvTkdpOgcS67AMiXTcCOyOHX0y0+bXl02xVa
1Gp5qC9lzuYhtf4yWKs344bJtIGrpCD1QsX0FpSxD7eAcuY2Wn/yboqFqyiNxGNM
I5T7uepu/PLdCxBSejDpnBUqpUaXPTWsm/h+zzGBIcwai0+U655sCXh7gy7kxVXp
2wB72w+kyLudJ7WBEa85omLJSaG35fCqmdJ/CBJKSUZfFN3elOaQIeSdxsQMecxW
lhGTqwOxpV8jHrg+Ol3+Xb5Ie1UNXXbHD1svZgk/9Mx2+M+ap/Hmbol6zOC4aKQA
u0YCdDG6gop8eV4FSwrvZ1kbOp8uEK9+5bUKxabK2lyEzTOjF2YOiLDcek1yYdzc
BVpt9t5z8s/gXTiDCRPCUQZK1Y7/9SkVMKvsYeeIWyPstiv6Q8LZFTGNJ5WJ7YBo
WIs04/hKR5BxOT0TJZo7SDYE2iBEERgGfMP23COOLvFKMQc4e8dGZE9rR8vXZjy0
0YaQA9CxJMHFpnpLO1u2/7yDSjh6wAVGOLUHUQNXhzn9kJQ5d9dDUDWdtsAunQ8k
iFHnCDhe+3lUEQcAXU2K2BY4bjYmxBEZtfV2kBnaWC49otk63jby9SLXqeAakrRP
9O9datzhU6WLwTJ55HfG8JEtpGpKXAbc5Y+YIMYH+U0y++jJl63MompBtIjtg/5e
SMqgUHcvmg7sG+F7GDT7nzHaaLhYZ3kJBVw/BEhCYe1I9VwThBnakPQg0p8VoYT3
Cnwo7tI8KOAwemh312Fgyy2THPq3U6npuArSvsFKQ8aDApCjW005Av+VjwTQaXma
UL8iUQ4UH3AGwsz7zqmKqSTSpNOLmuYDNNsQKzNp5u2ztYP6DunTubrWPYly6snh
AWQvb6LHAKcjbc/iB50ljgBE0kKykd0zXfyVgAAaJ4CfpInsx9hGqB2AewZsntHP
sGCFnRHLh2PL/+HSbbE6j/AnwDPR/WG/+g1EYsYR0FZm2WDbzUMfDv6HA3l1Vx2x
wzh9QjgellETAmfXJJggCRKtU14X9tnL06eIjmlyz7W0wT+40ihEinoOLA71FSs9
youzmy6dE/7TaA32NhkJLQspc0jsrrMK2Jd4XXKHZ2Fqq4nInX9hGYmXxU755JM3
M1Vue5ywb3wHW7OAE5WQ/aBMkCiIKrfMcpqBPa9f0FU8xwTMcxoSdGQy9N9u1A4r
/qhUakZbaPr6nrhTD5hZOHDfhozh6u9jiow3O7p8yN47LV6szIr4eznfyHc8Bxui
Gu2VkoC0n6Ryej/sgKsvkPFrwd1jNqJRhIN8UQpkMfELe5RgDq1F8d7JOzK65tjn
/nQhMASrrY/Rst2OtHI7aFfGnnixHOvsM/+/GlvXotOMyyUu8Zhrjz/JjHgRZnbs
i4BS0rOdcC+xj5y8suRjwFfddwSqC46XPySrMrcsNgiKEUzy0AlHe6MMb6byTn2e
3SHzZqVvt7pGcPHzyXJ3lSZwbQtEJ9lguvzsZ16EpL5998QV182gs2yJnyPWsYMX
HYx8BfLsy/KzrrrHsXjIng636JT9ihVBvdWX0mnb2APvIfuXkA/KrMAvwkFGQ8lF
GHKFC+yH6SoKYEIhsPR4eNYUlCcNVBQcD1luKKb2c0GJVDOZqUd0NT6BVSOUzC3x
0zE2062TPM/B05vGfiUUpYwQHmkBBdaAD0ldwd+VMFjbhF5VtcO21D+O4Z52/ObF
EdtUHboYsfQFK6i23O/dY8JnDdTngxqX+SRSPnPi/fd5Cw6AypY/CTmA9TnlmtWY
b8MBUKtL8q6GYRphTQBPrtunPIV/3DcI6caoCBGRShPSnIydY/voMEjcz/VPqPBq
lCixpMDpq1VpsFj8sj3WYmncx0F6ZCIA7GjJTep9cPN3v4nhp/lpIF4lN21C6ZeD
PD7tC4y37Nf0Dth0yvtHqVWuNxfHhTG54wWKwRUeMbkQ+oAKnGqHcB14B0NyZK37
DQbrEWJfgedLDhMhq6fWnIypINv0E74T2H9naCsHKL68MjgkCeEbe2eW/wbmPCys
v07YwHEwfq/IOD0dhQb5qRDytXnmihpEEDGf7aXz0dCI9CdyAbTGwpqTlkzKzF5i
dY27XFRsL0tqsZjSwucKA+zwWXhDsxjHjpcftA2AaaJFiJxQ7E8yxpnOw16OqARW
KMiXZKpRdr6CiB2RJB2C+QkRNaAWOAGtWTsD27kj0L2klBtJdRDZVsDuFApV1Dh2
vEv7s680uVmDrHG8lP9wQQ4R63MAkUCfPNHOPdPOybjKTBh1SX7l0UUiaosrKtLM
9O+tYoKpAPuqHQVR0q/qIRhMBbkBM6xAPOCCIf0G9ww7lxWQi4WiE31+II9ynvm+
ksy6Tg81j+8Ikuql5FNU+fhtBsZkcksJNDyFuqMFLaKCFPC6hbGQqK2vqWtg8sUi
BYE0BQNwpGcxZJnih9yCDBB7nBXsWDuRjFPj2QIznQcc0iQ6aCpRS9bgsfC0fgIS
+s5DNrxhHDKOJPy66vSWTgzHqVXOKs5hDkSANDvwWhkhuNlmPaId/zgwiuLWJY5h
YyAZ5QlPj0pDg75Hg13cdnvMS9LsT6S4SeKliYlStpUhhcuzogBHusj/kAJ5/87O
sOMl2bkIabe1ZHO0q/C7re5lkDkjpp0oj4JmkvBV0FpB9w7b25TVzb/zXvJDl1om
fds5iTP0sg+7PXLRDOGUJzmQQzRjn51NKzIgufw59DbqjSpJk/08eiVMPOHRhS/4
l8iHmE7xy7sI9tXf6ULetjPdQAAwDhyrQR58IwEOALb0UH3TlfDlLWy5uPq2ObAk
GP4WJMiiwn9Vt7obvK+vc1Y4Mzij/NXZYOCRVsQ/eKAG7Li0Nu043EUDCFxc/gQv
NKGD5nmxXejiNj06rjQVkom4lKXKb0yYbwxbAhgFPer/1Rw1bYVwlcgh1k7ZmbuH
jUdXnUxGcBXdph8zRR9Q9y1AfeXKGd4U6W36+k6nlDgucGNnWt/FHB3ZBCBrlzfc
ry1J1ZJtuXYitiwa22LO6wWyLtf1w1vkGlAi6MkP6fzqMMuWL9R/EWG6Kdk0u4+s
j77KKSNKd/PFdDYSdWfuLwNxK/PfXb2WjN7vdN4U6MoI5EIL91qlw2fsWeKgT8M1
SfPGXX+lnAAjBVHX8Yac4jXV0Ic4AJc3eq4w3eOzhF0CqFroKV01ATrtcIoVehEF
2qatRq/PVC3ZXntA8ESO4WfO0TArvWyPhV0A1GGkVx41Hdyfz4mmnz+QRjYKDUPr
aTvIm7uA+BryOACoNgQ345QNA5V4/RY4QBBQTo1gTPSbMTTP2BXlvR/XclWli+GF
y0ICkbJ9jT/d5FuEaHgkPF5m9UUPYKg4aeiybC6n2P7PtvHNecbStFYcoes+8FBn
wRYTFZ6HRGHB+R5w3/yqt/1eQudzVZkjQx9LuvQjM8gD7qLupNe/FNXIbbykg8Jn
lhLVJldWCOgQ5ekKZG/Aru7dp6bt7wiJD7V7Y1pzHZZeoS4FC1kj2kMeZVgH8hD9
m6aRUuZv7x14TG6n2/DnUEk+88ukYQha9KJtIvidKcUWmzzkxSkDru4P5TvDn9qK
CdAePPXPHdtZNUx4HSwiXOkD2C+TpKwRGqWKdV/RYYkpi+pZAdpQLIix7YHZ8BS7
7vLez/pYTvZe8/Ixor5lSNfvLElgVAAfeY3kxsNz+88IM7+OMdU+f6rwcbJyl706
1KBv0+ovxNx7eZKScJFF3KHFAbbRMCdjhJEZbIc4spdbw6eE3Kxon5UzqZ0LYTvu
MyltRgt1/xRLuoACAP0Si6mnntL5S0+U/tRq3/QTdt0GHxkOxiawmP64N/uXmESq
3pQ/cYwvQYIA69dBfjjgt6JPsJJo28mMf85CrAzRYERLbGfybf3AXYv4+KCi8UJZ
kQ+rMqpqxi4vrwMtF4zGPVEYO9npuLgguZSBvqbzPzFC2g6T3g5aW6QkkKMma0Jx
rbJkjjhGczjaVzFziklMf/nvL6BJnUZ1pPWtOW+MexhYxf48oybmUl/FiNwfxpNw
dgMUw8W77V1hkcXjkz/WcacTN+SlRPatl65+0vXGqwcNCkcxjYuXrahds5JHbNLK
CDoQy35+Q+XW63jCTF98nxJ05h69dewL5kyR+z1ASodLjp+fTG5cShOdt98Fo9EI
9Lr1k/Nc7UeEknvJAV3KfR3WQone28gUQkg6rPXwvcHeoagjEy4PtCPgZD2cIUxj
XuuQIIYRtd7P7N66oM0BBh4vYyCAMm/A9+UVru5H0IW18IwaTANMsWihiPWWCAnL
vUW87GgU35tozbCBz2yCnZKCVC/yCQR70ILk18qdQX98Xzdtv5kcwlF1GI8lnGxw
GAONrzIYsNM806Xs6x72A+NypM5xTmaiCvoNm9FgAE+e2s6BZih0Rr1FQ08uCSFQ
cNpAI4fWZHazEPy5leZf0GwWVZT3BZj7HWkSZi9x33bZCxDoapJ9zhH6bVlA83R9
lCaZ6zYB48KV/z6VwkzOAitsvMsxbkoL6TrzSOk3eT3lPK0RPqL2TT1clmA3RkY8
ZwaRdOAT/JERDGD9XKIUKhJhxBLGsxyzcgwhVB51R29Pv7i8JJCa9HgloWgW6Er2
on5n89Ghvl5mRsdqRh3W8Ef6ZO0Mzy1ho6ZEW8joNsXgArFP++Y1EkzX3I5elTMV
a5AAgsW2IBbdw6rXAe0E2oqg6jUO9Flzkn1h8F/b0dG0r9rMfdfZdM1BQK13djhu
iPkKjDzCiLIP+OomiMaWVq9QJhnjOcBtgTUE1tquebMtlR9ZR6qb25gRlZUqsQay
9XbReCfGV9cSHQN1AvJsGTTJ8a9aGSnQP6/f2Ac3iKlnimTcYvGGU2133Y0KNrGd
7Zqj1I5E8rwr9Jl/ixt9udxRW/az2Q8M3OvnnchGIUDh6QNXQdA2HH8uRmUkEZDS
91mmr/4eorknK/iqKeLrh2EcPws9u2jZcnNzT/+h7MWQ0oPX6lQFkOtkU0MM3Doo
y4h6Z6UKlxohNmIs6TXWs03CvUlOdsIiu2hApR8fHIEk+n5ABZElJHUhTVf38zyo
q2DApqAvad1jRH+hH+7nfa9U9BhqQcVXuLF61wfzFADhet+7eR+lq0nT1VKqQZ8e
YqVyllrmiAIkmQydU7d62MfnW4cuBVJ9UjBy/lBEGTzFcJTH0f+ki/dcY7TtMlQg
9HPe78llsjuLElD8xMwWjLWZEDrpgSRIKGGPsO3KvoesUuTcuIQB/F9xl12HyDnz
xkq32EfImJ4ZzZ2O8RKtDRRbDjTj3WsonO1BtaLx6MDEnTJyhF9fNnd8Tn2axHYL
LhVXe+qbbUpXCwR56sYokt7E25yUyugTj2tW8MaVPtJuOoDS4BSFVDBXAIjo+V/V
CB7k7HHOdXX1US4LcaPMXkLkI04yWoDDCE/pAd9bzdTcbPVeqBNogiyYDhlES9yB
JPAcdBNUbRD5WHW835Qz9H9ydC7ZOgfjEMRZIy+/Eyy1hnL2h0FVh4eK5QnGJcOV
FIa4W5AspeK/qJDk7GdH1ObTCO2/0Fd5XnrBKVIZZowpQeb8GV1C6ML8pnTSGR9T
322cqyvNkypaP9UzRsBD4J4OWtitU8UC2bJN9e6HjhwmLYD0W2KW1KqzXZBLnAFw
YsJijAGo3+m0kZqYFSsqSXIA/QVMEDk6I9xIw/44m2mUSPX0mry584xgE9U97Gqt
ncUYiL1H0/6qdwNiK7N7QAy3OBypFCr9W5jt1R08zjsXjKpuqxzCrizJK2aqmhVI
6S4yjKqk4VJNUkv2qq9ta2PGSPKTN44IRPlzlpNu3DwV5Dt3U9rsdA4AjU+lY+E7
B2Wxk/jGLiRf1BLUVVXO2/zvnatDc2ATTWaR15F6om9kqF7azUOZVWZIkvDiYZnI
PBo1lzATpNTlcXyre3yKbBud72Y5Hp+bYpaPJFEw9Nkal3wl+4/xiLLoL2BmlJvw
l3NYW5vWlkRqET2PAZLp0MNHai/H2lqZruULWM5A8T/dJBgBwusE2LprC8W1CXg6
MdwaOlPi78yhTbzEJ2D7fXfEtxmHYrfXuAE+yY/eUy7gTv6/13820C2Er0dhz9ud
tqUm64r7kMIPPdWBB2GAz7XY5zx5LeKnWRDaNevFHpwOMWGDb53Ei6XOmrHxbODl
/3j8fvkahl919Oi6hrv2GGtstNnhgJHRnib9BPCrqTeQbnZcC4bX2uC/JkK95AGp
BPsd0HW9B02EyZplPMgTcysrZA2zfEyUmXOsQUHH/FApzyHOIg9UDYolgZO266KO
frkrhHQ0USUyeFUXmKFNQQy9fj1aWAgY/PkttWrGwlUVjEYUfgnri+2Gax+DPuoT
1K9yL1/oix8jToNyh9niNksYbO0sE2hBF/PDMXkZPh58OHKXkTnaYwRi78s3PpJj
DK1FW1HjKqBEFncgJbkn/ErkOijvkgRGdQhl/HpjRcI3wIUCxz6oz/KZxe33NFsG
Nepq85byohshfEzOgeQ6ZDmZnKnuc8Gxkmr2AHDkda/HshI68qX+yhMN9VIWYkp6
xuGgy+SVe8VsWFcvyk7TCcsRdiwBQyi8PR5/NdboxG55KE91cfuyoq2jR/YTttYa
XJCX9hE9lU1QrR6m4VN/CUiLsMX/qFvUNzesQN+8K5tg04jF3Q2WNT8PWD5DOFDe
0p9DO6NLzkuECuG14/GVrEQQ+QFI2BhfGgIg73wg5EqyrBrourtDRiWO7B1DE7UV
WbqhN3k8GobUkQ13F5kNNHDh5x3bsfiLefoY1EQjInNIVSDtTWNKuDMpJy7LQe+x
fGNqFTshbd14zf0K8hgNm8EUafAwm5sa4doGOily+YTjv2SUfS63ISO8019EPg+r
BzBseYKdSbOWP+nt+nkD0HR/EsyZ1YstoLZESNb1iX+PZaGhd0LyWrssWqTQ+ij8
LPK+Sx+t86jQ6c4iSKAm6ZbC/OEGiSSQtVs57cVMrUCCgXRpbbyjC7Y69PyWQPLN
gwjqbtAbaFSAEA3vePhkQkuKdN6ho2shTCXUnhT95SNJAOPfj/VsSUyUGPBZqFkO
6MPdQgKjXKcnyBjJjDaGUnfjP0j36ZTcOvZApGzhPkiKT66BIA+UIG0SNNsa00Eb
hHBmma8G/M1nKOJxXPVgi/9qJFFJHFiBX4jKQP2yWHrRN/Gp1D396ZkbO15LON1r
rYd3nYuInGxGa7NouoDsweVq9+O64ld72RBvyxdgz8ntiD129KHbZiFHtFQsv7c1
7iYjB1yLGUS3tBP6STddBCoy2a7AN0FUtKJbd2WvbyFTwq1Dwrmjg/tTEhN1CIPu
b4WDUB+WhF7Rh7kcx8rQxYz7JI+1SsBDT4XrWCsCIJHVNIeNC4Iy5+uFS/r7Xcvz
A6qGmXFv4kbJIepu59DviUZk67HlMvYWMp0/aCNlZqRx0er2uHVm2OdLz0wdnpPA
cP+ZWMrA0jCDLohSgfRU69+BZzS2DU4Crr+84JXWYm8IMJEwDcspdLPSnGCSbCqz
561+UJEy0ty2x71IIuWva7z5lG1hcOQu6wAfhwbT+FYOAMVUXY6Kb9dHx0TTXuY4
38O3pIScgwuIzWe9mk573q3fOFt2aITZIOiCirDLITDP67kIIDdWfBTdiMWbhQII
5EWyXOLIElYw8Pj196PfADdXKbFbZvmBrNpw1LkFA0RxhV8d5Gx4mY0qz/DFlFgH
HxR/GxC9hLb/xgR4gHWofHmxR92akuT07gHrZQAD2oRWqoHPX/nZ5qSHTKhdOW/E
FnOdsJtsooUyTVNpzgBLeGypetiFLJnegPlI0wFmw3ouKH9/W4ZlSC6DeAlJyVNI
FzuSuDjVodfqNPUIiW3eAWu9Cyh87ymHcNs1wKHL1sputLxSug93JjM2I23zZCOT
l5RtHV6n0M4yhB6RL2S1WRZu9iusxM2G+q2zXRqYq1f4FDDWCT4dAMC1AvhMg6Fo
4hCWIWubgFs8iFCBdE/Up0tm8XXvDh2FL0OVo+2nekrQEjDOp7kLqkLcEUODpsOx
IHewBjGKsOBLoEWwD+abLsn1O4iq5FbZVtajtGbQ/MD4hxMgZ8Bot8r4l6E3eLXr
xrXgMedMa5f+KfheGCwl0c9hmZ2CEMxuz+pmpBFYWgMSyXysAV1/UZnItu9m/iuG
R4KKsgLIkIvjJPIeGFpx54FN9NvWmV/TAQ9mHD7DzXDlxL0BrCVT7goha/qcdNzf
sh/Yuo8icqPczxNGnBW6EGo4wZU3pzarfObLaldrqDwQ0jjNvKm+FU1rkk8GaEfO
dd1hggigXv8tM+a9FnN6pPaZ8dcrODl4Tj17e3WUHTtShWBYNVATNb4+ZtcZjuQu
mhEUdLwvmClN99/+usH95BvPLR26wrjiEe0t8REnCO/LcDw4WCPtUUk/Udx7/IeZ
MqN7G312OUsR4jGhVlFdPRARibMhRPTKI3HtG5F9/DPvkVJ4x0podRq0hoNhyQ12
yMiZZhEmr5UyTyNbnDxU8QrqbxDXUpxd0cvDpNyaxIrJsD4Th0tnicRrHaxsg2w5
AooqamgRbZ9PycjoLuVAi3aee8QUt3x7vmwzJfycv4s+QDLJyXF5cK6tjp499vAC
6QctTdAmEZcqhEDDpSnL3a/NTxYOMTLaffxNpZf8o0lC+Vz/oTyZEfY21ZxvD1Cc
xHx9NvEhJGrA6U95kxrdY/R5xoZz3nsxyanxbAe3vV2Sk5/Tp6CRqux7+bm6Hlr/
QBasY7UGcnRwAInYLS7TM6FP/P5FiSVRjromQCQ+7R8QP8okgz3c2JbePgUIprwN
1e+g5qJEBPXvEZBupTpSQh1uYXEDRZf+i76NA8Se/HKGcVlqoj0UPjw794a3xXFZ
Y1M+Nq+DVHnYmKpGsSWI3Q5Q4KaCfWlKWGvmmGmJuESpaq2Wy6qtojfHgt8pjKmO
4/b1WEU/mrbaMOYdGBvxMn/GLGeokR/m1HATkzDZfg9kDS9avOvgZ47j/6hUO0y5
QUjc2X3nKUBOGgmkBRkEHn4vdJK6wGhp70Rlz2s7WPV8AbWh02mLVg39dYHi+o/3
xxJJp2pUeawAFoVJ1HlVOl58F2z9Z++YVKOjViSWgJkwh+hY80FuxbVmISioq4YS
bqOi+/A6ioF4ofCSmhcXpLWEPrsA4W1CpE5V2NhRZNMV3nb+INOenRIZsXS9wJ2R
LGEKhdX1qFTv43MIvmpwvWoP2JFQUW+261603M6V25P7kU92q7fhuh7oAzAVdYe3
WW2st80TxpeSh2nM5llce7pG/SbzjnrAdcFogFg9jv2ZY/3GT8I0BdnBlU5TSID3
v9aiQEY+N/sPLnAIYfgb4FRSOmxgoIixol3614WsqpykQO9GKQFavtPFJHOrPyPb
Yj+yRi9tNQCkN6dPua/dObEpRtOYJSFWbwkjgOmbA0P3atpn3KriKQYBHFTqBwmj
mtkmHBKKGMTSGeiuH1cbA2h+JsdcGUyeOvXvqSzFuuEJJCC+ZF7kFFpzxigAnyXM
9kbIpZtJS685cCtQdEz01CjP9xwiUDckn9N+j8g9cPUVakbxSDUGByB4i2G2baR8
PneA/pKx8yUXMRcipT0D0s1Z9M3SGVFLpZ0OBOfWL0DG7xM8mUi9YboEx+wWr8YU
U9l3zEthB8x6zU/tfvDZbQXXUzVCR6LOJLM61l6U2Y+03WKL273oB3gdNZmwpwZO
o3VFPDLwKrk3FF6SFFrGatLlae7nMnqs41DtTDXtKvgCyLRoJzpqrV3TOLNfvLEJ
1o0HDdP/UulN4/rWzyMoqy4q6+LiM4mCFe9gI5tcGV1iUpf02/3AbbhsfqoiW8X5
AREAbBGGMz03iUTOhtlMu6PwJzJw7kqGhnAA7FWzXvawnIAmzXi4c7ZVcbyCsp9x
6x/H5PNQ28mYRYmevc6h4Nvvp2B9yhHHzzzuy7kauV4aCwLrMQVRvSwLCXWQqYpv
0ofey2RcMVIwLq1nBp9DmpFFYdzOAqFH7YBe/moR9sdQsFKXfJGnuh12nzvXAOPR
5XVsPrAN0q0S8eu2uikHoVSJGwkAkArDk09rSkO4fgMBVZEu2EzCFk2UnQZZGIZM
WL94SA37+MKN/osrMjYK93MUN8ehSxMtO7Ipli6JnknYWYI4P68DANmDR7s3YdFE
dBHDubkWIX8dT3QFF1gP28qkEEuTPXruB1CzNxnKaWdDXvmeKhOJ6EtWLv1o/8VA
aYGxCpp4xRUi3wgHQuYybjOE4heDQZemWoP81Cpswl8b4kwqa1uBKvy/wizA5WW7
TAuoQTu2P/BizkUhn2Z19M0/6CBXY2cvAxTMt2zFyh4ONlG2OAQ5mva9o/fGf3qg
45YUli9WqWjY89MfpFICt37Mu1yQ+1S61BP6e7JE9Nr0XUPV3Y95LzhgkXMlQDEU
E/VrgjOBu5uf44l9f6nCbn7FtV6PDeQeM6qMOTZqRalXMXEDygy4eovDCRs+HJsQ
LzFkGTgqeoOrMahQXqvgPob2bQVWRG+M5ZoxB5Z5cZBdo6+EWSq7mh5EWqsAWj1d
8cnlyVXULGCCRR0aTG/sa5tGLmFuwj581wUFlkbN96xnE1RxsyjepBCX/jkicFaJ
mz16H3ypFvHKRtTNvWEn4+jp00tyCQ2FHrzg+O02X3NiEZF0yhkqW5rvkduGu5lk
fSqNDEsXNHA0EA4jADg5Br6cKODlvpW4Ek4+Z4sXx3zB0iYNNuDiea7RPJekWOhM
s0yZRNJjsKdgqzSp0YlK9rDhOeRiiqXpkOADtWxTm8xnw2kSjnRgke5UiXzbINJG
3CUffcAwYgJW4z6tBs7052BKxiDZUjyHYvJnYUZ16jcmuSMXkEe69lIOjisIUEOi
DzQgedy/9b0Fd/wnScKESfGerG1QnngFu4SLzdXN2XLlS727GAC3gNEEKkL3waRt
tTyBFrhv3K20NFTnONByHbM7IfbdHQnDwgH0z/GZEZGhUiz2lkmOHl0zDz+6wS5K
S4CS7PxE+Sm29fjnA3qv7O+cAxwZ8RfOXW0h6Ze8i1RmzT3rX43ZeGN28QlsQHrw
OE5pLSr0f9XPVWW0C9AkYoN07Ay0CcmchSJJuPnHlyjhIhK5GU7PrXjy1aaBtwsD
1IQSVy9v5jDlZI49nHd8cLSVDNpSTDg7w1TxU9PWaW/rY+ET+/ymginSgzUSvGXo
c6girU0YY/eAPfo7a7fs+ZNikck2Km/ISlefW+BMqJaHbCSmVHSANM1fdS6EQJq7
hlpKBlVczt6lajp/liSCHJMHYUcm+5O3xCO+1s8jmTEIHkXhOg6xrce4PzHgUcPH
z3gSLbuFLzMEsWooUD94V42sLH5nDlsGrNW0qSb9dg1qxkp3NAKEd27K+UCXAo2K
9j+DusYEp423e5L9QErB5en2b+YoxQxXP13zEueePiS4rrgao4e8xgSiefIKxqWd
+UqyB29pTLTC/PHgD+Spt8zeUXCDsNFGfABJ+9cnVUxUuYkaGD8JvuWGu4vZJYO7
ubt1jsPmKQvLSg4KzZQawiOWBY9beDk6ZNp3mHXcnkQcwfTBHnm0oVxoWoOfd0tl
EE+n0WgsehBhACKeH3Px+91dg+21UZcj/0lmwYTfELr18FAV9Svlv2JwvrzzQ0lb
HnlyTVRtCEk2bFvPIVrqxI1oajd6CGg/p9EL4111JIU7mepKchRgK3n8/I8dUbSY
VmPiMEZ7c5Dp4EcE9rGl8CQ3SuaNoVGiyydHyHj0wB8nDzWt+1T4BafCOXWaNAKE
3BdLu8TuaAwtqx1XAftoR/XRjSU/RMKHebAl34sUMOIdqNCwaYwfWDGHropWSEWF
PEXTrPMg4s1zDOYh/lmG3EbsdGuBZkYaD3JyU3tzPzYLPh93ifXmXF3KJJ7Yi926
WdNpa4/MD6xm+LheySwQ2hBikLiXVZuUMOIzcbgkxo6NNJSZvgeJV7oR8xsCfjns
fwimvdcbE0XUBRLGK8oKi3up5e82RoT7FCifQxmKS6cyKG4do7THYjSAtbmKK86k
Q4iwtS3gwZRCpx06oPt5y3HjhwmizhJdcnemQ1E0vFS3/j7/mLVXMFIOMhJDsZUg
rV9dbEGEesrGSjML9/WwXPrR9TjzRlsOmMP69ofgwOanMpe0JrilwvdkIrmU1BbE
PjGoSVxh6uBDfmdMSw142j6Kc8hghnGO42XTvHnthJz7O/vllLVwA+bk07rPlk6k
aVlujkC7BYGh1+Wjwo4Sy6Oj9Y2UONhcGmKE/Z/8P6P3vpChwHnMeaAZzIx6W556
+DsnuPk3opRt+Zdd8x7zoxz09BsIt5sY/3mCXVIZaPwcCJcIethUQi+PleSD/4cc
UZoQ85f6zcVlxE9De7g8gvjb1dKq9qv8gsiKcxPf/BWyi7EY7K/Wx8YNLt/xaoyX
51jeZ3aTjiqkbwfUMF1DmRYhuOuueEgobcN40e4qAYQrFQNtYHJs/XQP7DLom0KN
SNjubtfLOidyn46wBxIYqwIHBLOb7RWtEFWIhyey+PxkXNZYtMfKPuKBBzfL6a9k
VhJ8q9uvnpAacr3rcJDKIc+MBCGMrzrMBpjQuK9GvWcbaS8jdPXWVFeG4VC4ppJq
4pOC39uO9C/2/qHTUxQY1SLjiLrugwsM3hI6gK5DTEmejsWubFPh/fxxTXmVNSn4
MrW8Rad8en09yQa6YZqKpkFIA6aUAd+t8hPdYOPmpPPIa9EAUnb024aG7Yvd7Q0/
v5wfOP8T6D+mB3aV3nd6lYD9LGQ/0FgLrdtx1zD1dns8Ow9j1EKQLfoR/kQ4VYFg
xoNNapPxmunybqrF0bj8MaQmHE4I72qJSUy8l7v9gOUutikJ5mkA6qC3C1paeTmP
CbXxaClZHxiE1lN9AXrpINQuBLTXh6i57vSE5y+lAtuBY85r0Wb83G34qdiuOrQa
xXUS+rOS2C4Oon2ZoVWgqKfhTbpjchTblJ0vJraZTMvObBYbK5RqkuTloZyklLEG
XJDvi361Hdf8F2j4cUiOycH4O78/BeLZtHE92oUgB4S1NufLKJH/bQYN73iL354l
FK6VZeTW+tPKmwEo17VuqU4shXxTnOYN7KMbNSWdEbz7sWJYNJ3ztFdenHDmVh9t
4LslF0D1zhV/F/V9Ei6/UU0HjX3J/GxMgv0QtMN0NOjmJUm4VipzMIwVKY3yUt+t
4dpOLj83Oc1tkltqfYZE/vtWCb+lyy+c1AoJbn8i1Ny1G+j6TYZbDnsSctITP6lb
+WVZgtsBqXNfvzX8fABDSDyh9q6Uyt/bd2WbILJVcxFf4q0jOphm0dWGTIA/LHsO
jVGR/kRM3N5OPWLFeqxfcWFmwhH1As+ZXxeCe1q9A4U9ULftX7UnkRcCLmhdqmTL
JJLqyOMlJCRR1c4VfhO9rdDgDA3lkdD/1gxEMX/aTRv1TlrEOFZVfGbdC0MXXZZD
2uw4EtQFSsfP5Yw/QtCJiGSe809JLLs3wQUCCrfb+KnzaaX11wKyo2Kh0bu0Y5BK
/j7m5WM8w//8Yxzua6HwJVkfLmjZihob7bskfD7tClXKoL0xxBIFTihGfDMMPI3/
zS/9evZAJzRLEPak2iZUi6iNaL886jpNJ5AxAUOAYlvZOndF2FSwvGHIFZZkoPmp
Bzu4ExBGzyYG8K+f0gGU3f91NkWO2PGRCFHZ5dBP8onHMAWUJKjmgKGf51EG+UYY
iSr62qVzY0Dukw9wdb45yDar0IRyvw8TVpTKyV2T67EuE4m9yw0UJqqxtXvO8TFy
x+wwXyDSEswfCkhoaOkKTL0MMcC6Qu3/MtrD6YAx+NY0QI1cGgscZsmCr/s9TW9u
EdDqdZkPnpxv3fk9tJxy3XjneiTU+pyOP1sQE62VK+gVIhC43YzCBbGWWpBDuj4F
4k1/VFnOQJeAGi8JGEar39i9TvzsOzGNOrKglgfgyll7uCtFq3bxLHCtlU2W2R52
R2oyrEZxNjKYT49JMA0qJB4IJ4pkb83IWPpGFHbC4UOxzOndp8gqa2ntlvy+vF7m
NsFwck5K5zSvgDNNUjBGQbE1325AhXSgKHWuh9zocN5bk1TLTYoLDeJYjM0t0+JH
Y5FfuENHk6P7geqJ6KOVr2FvTpLF39TH5zuGNGYxvrv81Tpexl001Ig74CBHzCN6
cH6L15QV8JfBqBm1xY6giRf0j7X4OViGNPX3S6JsUfgtzud/8ig+Zm4iiGZUIKSQ
h+ZEmNswlg3a/c5AQUx4pBoiR/nbSVvy7bmpPBcmEJCnvF2oaOSoLBd9UzOvPy6P
qbbkjG7EZ6gSMxPoaS9qcrwvdx3Ll+qqfFAZPzeRNUS62EhvYS81ACdsv0rOF77S
4c/f0L3VS14IkDI9w3DLlK0U+gTe396ofiJOyvPSSYug6uxTLBheOZfxrmesUBxu
iBfqZuLTwH4C8++r57+V+eU/O8HS/CYLSfGNeDE5ejSwY5GiRAWvZg9uEcId2ftm
UPcA5cVWPoR+eYm/pKIHnXH2XjI/swgKQ1b5UqUL3bDLexdvzy1mGC3uJJ++Lgre
VA/PgkjZYUuFN8cwAbubf3DUIa814vRzE2Jcps4Wq+BAna0SnCLJ8/MqJ6A2L0JK
h2lqF4D92u/qCgdTf4HxyWdSsW3rhefuGs0m9C7JCwzJ2ocghiwhifRra9ByKxmc
AQ2f0GYziwpqqQjbUEK7SAKC3JQiOzhiIknSt0IUVBRE+9vVSeNh6upPnGzviRwF
nawqG0wcBFTPwj9NFuKpm4n6FAKeEBeafipVRYapw/erEUf7KloYPYKVAQU79RMV
To8wZoT6LrZm7leigOQulHclFDLXDNeL6RMEHoZCaGJbKRZMVXc1tXzwcOCTJKOU
I4f9c+uWxZMNLoprDBnNdfyq+1YkRe3mDSL5hCSquiihfncjI5fE2dHnUIMlTuPO
PC/2Aa8wApDK3LZPUsxDl6sQ3AJ9EnvX4Q8mdABXhRRqNkjigJ1IHV+x+LZY9Zp2
RZ1SeZsOE+dw3ba7uGZbtJLVvW0+UxQPinqz/0o+hPZHSIU2SWxnYjOlHolURotH
4Cwsm4zr/6mhqflwgxSKs3uGaOcUE0NdQShPet4qXOdl9vMhnnShoHNSGXiFIKir
3GuHPnEyRqcTeVzVI7Xy8Y0r7RgrEe02SqNN+wuCmt8PIXlxnQtyISEthR2HSOMf
HJk5DssQzU7GDWl3Vgiu4W9ghxF3JcD+ohtMmYWCtvOKolCzKpNMEmJPAlDO4aGz
YENRWZUbnIqX4k7ce/113JTwNzENzdz2K1H5KShYsE7yvFTl3A5mbCL5Vzwn9zE7
ZXBr5LerUfmw9hDRfeMNsw8n/QqQo0cRrCOE9aJhpARIkZWrFKW+M+nMELqAFg3k
rL2Qs0XFub9DTfkxp3VJkHYZqs0dn9kUSshYL7sAhTyikfXjY9IjikrIFkjshTPS
oxZsL+qhBoRePBYMREuY+s1MZJOxxSKlSn1w5VUpmzesaM3IagU/e3hTWttWnEIq
bgcKM3TIiVdo/ztSWzUHIa0E9SXBmf3JtAILy5KxwbIvT/vKsnCAxcRkD4bckzEL
NWywwm9JewNW9D7lfb3zDMMltDmkdqHds+h+ceembAyu1LbDbSMpNj2mQhzsQKSX
jCWtrMB7eQPbXf+1cKmW862WsUTNrGc526qsyjfA4I5Wo+DW9Xhh4swqP5uWUN/p
tbl2Qu7lhPhJu71Qn2B45t5W4FAaZKwtiiwHuRI6lxAjT0za/ZFyPD6DWJYBQwpD
P4AOPBuNFqweVDmGa00K9AU2a4mEb7cZsyNhpVexDtlZZtNU92Va2aQZnshVDzih
434L9MCC7tkOPpGyCmOGr6QD6cP1y9fYeOAbipfy8z0/2Fk0kcEc6wpkO4nhkAUj
tOCGeqHiIPOFGi/P2EYyWAY9syTZuang0X8uG6m7/R3pkvO2EmpSwGiiZ+vHz38l
X0Kjs9NV9/frGjNeht6aYoWVfdQyXVytJH8o59jj2P+LR1bnAEQbNUalSWK/1sw8
qbIN+qyMZGH7IHiTedegA8UDc7EZU5xa9u9uFkiBFMwgYs9ztv4RPWlXdTHUqhrM
caA8O9BvHhZdKFLOUZ0vF5BS62jexz+BBeMlqXsCcrYLLMH4+G4jzkAVC9V0ksju
2ZsERvB8HnIIQY/WMezjx5d0eYbqj6gAgDpWdU1PUIHXMlvhsjHw2sEd5QWPkv41
RORLhnN/xC0WpZeo09R0YuYKEmPyi95PXlnqz4S+8v/nBt6G4+4HFnAF1mqPHG5e
pCKW+vGxFNbWGNEznduNKQkOOSHggnxcyvTWcfwH4u/M+Y1ljGf9ak4oOeSExUrQ
aoiohmZ3qZYCh42XmnSEkpaa02mDYoM2X1TKgjCt1zxf0f8Bl3eEIXS2wUgnVkxo
74Wqto/jh2CFWMuSlMyAZa03GFHjoI8kyrXx7V+fdZs2t4wLw2FJg17gur4slQ0e
SIJQy6wCe/fFqwcSamdgLk6BYibuRAJLteJuJyp06BUJal97XzhTSVavkhqwwcUG
/dHbjUcdJy06+lBNV1d9RFgQHNhvLHToPhak41ZqgmMqUniULVsNruX+qt6jG6g3
U/O61ubn1aSlLUhZHI536VlNtolZykPe0TE8OZYz5C/I6MpO1l8NPMXDrHdgE92Z
pWn1C5RNoJa6J9lQlmwrg2VOq/7XcupL1OEe3fNrn7OzOqjA4jODQK+iDtT10JT4
e6l9kp2h8828A6DHKLnFxgaiMwxNaDwaaczwuxFnKFQK/JMqDEG5TTcie4VJ+usz
po7J/eWPbVMo+FbaJD5AalGOSazRw/EE1i72WeEwDa+xO7UW/az149ZaWMrozvgc
rvTQoMRhn+TkX23W3xIpS4zmqPJi2Ny4eDMEIouwr5WzucCxT8JvMQOb2eTpyK4R
WUarVkKObYznLdIlX+YL+9KBKt/BTzH9FICIPJlZndxQeVUCTCPkrMIVIldcEki5
G0jzy2Yw6Vzs6s6EgBsmunhneDShIGW5UzTYuAMqiDXf5k+xtpvhKp8SWNOm8JcZ
OXeY2u0VzX6ehqtBKWKJX0Whoi3nvm60g/NTDn125+lIX9l2d49zhcchwyO14Yjy
/9bVNEHj6RhIZmunSB9wfwcLOeMTWiCEPyYRpQU4hyRv1C9CKfYO52Ix7/h4lyGs
ftDyjdvbY9qcj11xK0EAKeXz2dcJ23Ho7kEkvHyMf3WC2OEDmQuZTYSo8R1GzoG3
Oxmhbzh/xcmyXgeZiYgaEbq4iKBUxzldhmtZPZKrq3+xn6COj1zjXsjYpqO6h+pr
mSuhB50sdnWAJBf/d86rJpdk4L51BRZSPp5XX4Pekth48OP0LvGEzUyx0O/J6Kog
Hu3y+AiqmXPyYB68kCUNmjY6bpVzq9EVdzsBVLnK2X7X53/Ae/koNnGBSD801i6O
4/dBOGgxTfxbGJzw/wwZVEImOzBP07vK47LBr3nhbSnBeX2zaJt1+gk/e3U+Vo9V
d5i26q7L+8telDL+VytPj7IhxALoqGSj8Uccyz4Zhzq9OOMLdZoc2CFAcyeqLos2
P3zvezGrxMWRhYjVG2Cbo4DcypcKY+hKSBZ9kISIFGAK+80oSx8589iwCqtX86ui
Di0vLfjfhBQslicnqCHPjvIUo0JWAiOGlP6v4Yt/pmBmmxkGnyD4kFniiTxka0KM
2Syfcvpeg9/MZn6lKsgppKQmURN70Kpt4Wn5uwM56b95InH4EKGpr2Lu3P5ZVYE9
Bkxr5rm1YtSDapYD/mot0IMd8/jzy5IzsiO8FXzWaSMDkjAIs1Mdx6N6YcSI+f+X
xtt73vwa28Qd6BvOcUJLySnRlKv910VinkO4n+8BoSZR73uaui/QOb36iwHohNFB
r3kfefI1udT0HvFMYkByBlLpyWAfXPlSs3kyXwDxXtfoMEEOcpOpzegp2bgDDNn1
GVswfnomU8m7NUPI8mRGxCi2+Rz5/VRZP00Nh5kWCFLwR5wvLJoydN96hsjCWrsM
YqaxGz2vkFwX85d5F/aDo5OZljwtdMmUUvjYfvX/j7krf9Y9hkW3Ee2zXLdPDcgd
zviP3vpS1TxVGEUKH8l6z8Oby5x/Y2HJ8XZ3SBEuJrWNjeB3lvuM9i4AaGMm9/fE
R1DBM871EjZjAao8COu72/N1QKYHnsDJ6ltCuX2IIYu46RwLHFbB5fe4ETZSfS1K
J9UTrBy/0UJzxZB/VBJynQU2yhUjlMBSNXeWjj3MuD/q7ZoazML9ejwucVqKmQGr
TPcQKqV/YryqInV0TLAwWc9DZlkG218yjNOpq3MLSTokR8UaMjP4ZWSSeUTDcOG5
3SeG7++vFf8xz/gHxyRrJUFD4Y9HeOpJF+RRRD1rIFQyVP1dQYXQYFqpYH8KNonC
lZlCgXeu7w4b+skTtNu/FlyIBRXG/ZYZba6yiYODjqBP4Lte2ORd49nSFKSMDeHf
aRD55IuXdf/0ruZfE1c5H+Zgw7N15cWz/gfXZQUg0NeS67R79TztoTGWiQQGdSaG
97qZvLAy1XBQfb6b0eENhAL1N4roxkuEakqUAqozMqYo6vULScnKpOS2FxUoXlTl
oXxJSNMTcEosukS8EcMnGOhS8Jgoy7FkzahxvstEJOX0YKSO5+LDnVMxEdJOOfNI
QdXTAbcTXGWqFHqi0a9VbafCzPPfQEFRDg1y4A6lMwVWRo0rqtlRkpl9PsqLND+n
CzH6NaAxmdH7KGTDX3HYHljwuhtnIpHVYn8R5O0n6FsYzwdUIgyV3EsVYgYWgY0B
lN7dn6q5Tt+uQjYMBGQeotDu7z/2LqiKYkGi8/hRACsvh9l72MnTZtLb6GjdDnKx
X2l90va0suw+/5jsZLnDMENphGSQO/eIjslW64ABuHMB0HC8gS1OpHNgoEYSpcXq
FWfq0g4vTVi+xFKIIZIH9ZP1vZj5fsD7SS9xksqwdMnZRTZbz56yII62gMmgVZu3
Djj9JBBl7etbgneI2gm2TDme/sj3C/Gf0fsAcoxw2N+mwpiLr2GC6DzvaWYBKslU
4/le7nUKZhP0A47pr1iQrhIkXlTbXIJ+HMfGkuL6nSfEK3u2rBolsYOwj2y/wgQX
5MfrP4hfypOmutVVuZ2t4kREdue5n1l6Ki5xPbDAmC3xTh0cxqCffaUdLJfM90fc
EURFfRQWc2A0y8cfAi32GWkwmUoiu/aM+gybwn/+KuIvXZh9V96sKRVgrEsOnHq2
Ssvg6rSDbem6kBI6jVzytENudMeFsJAWFtgPKG/KEd9KRfK+h1dhiz0+hSEC4Ddl
Z8lYlRWCfWh7hZ2/I0h+MtTP9J2uEzzGVj+48/d36pT+7Hlo31kICOpVsOWezIGM
ceLLxzNYQYuIAt770pfOELMxJUrWL6Tzj5jykxgRdve/Ulqpcyg7AGH5WwYBG9fm
1LYs0joUV7znqu8rZqX5i3VfxPq7o2aYgYwZ6U0EIOz0ElorzAA9aUfldSvLT102
Y3mUbL1WN1TSm0ody1rAPRbHWItvtuoyB724vXQMwjdVOQSohGftLoYORffAFaId
NAcJ+Udz2cvg9FxPTDeyD8Grt1sUJuxAQ7sPvJLb/EGmNrYK2fYf6X+6RNYoLUbK
I0rcVh6a2QAnbV+zos1BoJcRmH10/5Lf0ykjpK/bvtlCRR6DXSbQHtSXcjNns+7U
GQVAVaDYHsecu7saqyPUTsw8FPieQoZwBwxjIQLveJBagksIquQew6Dt2T3TOpJl
4UPjDeh8NQzqP2rR8JMS5ysuYg22ynHbBMFNb608kMPFuiY+jXaH76VJkTKHQmQH
oTgAKMoNqfyp1wmWixBOzOjwRxFjr0G8YiXyPNwSsgrHYg9GAC0cy4U2xUtyMS8e
cLhdjWwU+mTPQJCL4ndZXM1zQOE1yEHweoOBpwvtyRj1URbLVrt+zrYsNdS9CeKa
A+0Ft1msQMXmqdtZuQhWP7rdMGaxU95iq2LYXlCdnhitVEbr9hyrTiAfMxGiaKPQ
b5pEO3/19eTbNDx6vdm3NI0fblW7Ssad5n0LcFuS4CMKg7ZbMUAInOd8eLQZ286w
oO7Z7FaYxung+KpIJcAIfO592QJFx8JIfUya/0InW/OgFVZVp0kmkgjFFIxoQNTU
L8UNzj2ENa3KTbXH01NvfPHW9GMf+cRBp7HeLhTalvs/BqdYWdhAMEI+QHFAn1Ye
TC7lROXU08j1nICq2kTWHktGzpiNXrsaIB35UzeVc9itz1Yw/+581XOUtq7bvy+X
bjd7yit4xWfOFFLGjW7b0Je1Uwv/AVx6T7a1yoWIem8eyq1X+rXjzzo612IydEcN
IQUXtemSUlyzrGIoSix4osCq19As1KDiw3Fs3Ad2Jr7F3JfDnBA4tjs6bbaEze+9
OfYu20n22chdSWzwk8EyflbkjCtXlinD9IrvvWIY8W1EabR3CJ3mmfdi1LcP3BwX
cNCCKWq8zjdaHy0bwpgF43v/JInq2or6EQEpAOtQBpA2Adm19pixhi+WyVeGtqg/
zv0EoE3wEDQerGhkYICqK7XD1p6iKE29SJocBLz+NJRdIkEqXIRovsvGucRpEc8/
9auAie5jzXJqfClLiDnmNd/sncT4hHborZ55lWLctn6Q7ZhyP9oPtpSt2RjQo22k
8UbFV9iW/Mmo72MEZIPDYTlgeiCUw0xZjvJglNP5lhEhP660ePlzCNW9/EwJ/Ksq
WMaLIz6yIeucfYShESr9lpn0SALj+UVq83PxfRmrf6yGj9lySOPjbeZUzTYGdZaU
6DAeY82q3Jvmzj17YXK14Zpgyu3UO8B4iazIK/MXRgdbBwy+L9X6GXgX12gMXEjS
nXqR0wpLRqHdhY66dQpINwcYqtlM3AzwYI5aY0ACyZv3Xp2qfMfsvACuK9xRNW3j
r1s9boeF2g7rRn+xlBekS/UJO19z3mEkHg42s7RyEVHTjQ+gq0sAP6CbxF2aoxfe
vy1qZCdLd7943ENhag5iscaXdWKadUYAzsCclPejnLl39087VZr4vFpfVHTzBiXi
mKNOY76ZiUJ6bHUuthUR3Kjvk31JZ7K5a9KjnMeMuEAzJ7KYIxHiyE2nrI/OJw8+
vLKwNCz529llb8HhoinJg90M5Nvgspq/PRRM8ntPIF0doBPOnNF4+4sx9g1+Bm+0
pTZqIxjGxvHFCcFZSF++7hjjGcJ4TE/J6ql7slqc6XYeMWw9GNnTF3bB3PRkgkk6
ycaLT/xi20wGh7Spz9RAW2/zuEEbzkbNkkNiatB680/ZrwnAGTZXGyFGPuEfb0QW
Z/8wXKIbBd0wZQviIrY7OU6PFNu+PuezsfSD4gA9mvnlRuVj2i3Oonv6oOGbOzx8
kIBYm7P30CXiNaEGH9+XbTY7gyD+f5KYjoVaoCg3pf8hIzTP/ej+/mXJtc3Awuh4
pmYoFmsq5pcYdYYH8QmZkhjI1nEaznsDrO89K6ZxXUjsOyV10H0d7XuNQTMmbpxM
IDRwKPNJYzbvBIQHecMUbFQ5LT1AjXONvt++I0GMCRyWXKPxJeqNMMp7EQzZKaIO
Cd3MgMrw62aQJpS6IWjqvrIOOzwOZDV5EuM/2EoZogVJ3M9ouybMY/3vg8hR9UNt
R4YZydw+NzqORN3Z2x/LqnQy13uDAX6rpHghZeR/Zra4PjcyvtyNzFfFUqON5QJt
pt4dcoBJkrPWHf2xdFLPTW+Hhb5HOhtow/S8Wot14LNzwUF32ErbQvBSZFRpSi0V
Yt5Ms4lqDHt/h6rB0PHYu45R2pbhtTd/9yO9pAPzdgK5NmCrNSVmCS8bUj78D3IR
uX4sYBrWM6jYcfwJl4+FT/aBc/XQNxYiHFAiqO9YRIisqlSrQkmzt4jyJ+1Eyz1k
nYIqvYPETv+U2Im9rto1fJ21hzPBOSfdaMD+2J51N6UBq/otNya0ScInlaxCqRDN
K/vPmBrsgmxFhyo5LcQh3/mx8SmJSCYFiCbWYfTgk9GCE3Yg9tXOsN49k6f/RpdU
eF4Qtc+9yrR0U/wre/PILT56iwU6tu7cB9kME/RqMVXLZag4+eEclZLUGmkpEZfA
r4Ppblg9C5Xht4zHpz0ahTmde3SMapGYSIqJwK5yCWLqKImlDDeN5TLxNWQH8Yif
dn+AHWdkMxCw3yDmV2zbnaNH4u7wXmWSCekb055EF6an7KjrRGpsJ+KqTIp4CJb6
WMzAr7QjuY4nXAbPCmAYrzLWKyk5gOyMoVTBfi2rWnPLCFErwHcWbIsz86/l/8p1
4w8lGi3VW3RF6xXfhOBg7BZwCzGiVrZOcRpId4iqZmfYB1+PfHnQMbtCQafHl0Ly
IaTv7g6V339P9SWiBmPpApl9TkDq3ayeZcIfgYTsU+j1fTMn5XcXTQ+VRupfyBNj
TX2jBSePjdXvKrsmrbWvNemhr1IDNJsZgI/c9Zm9G0krBMd0+oAiRkVuY5f/8JTd
HImSF+yuVbS2HqflpuLkg91FtpoiV9YELieIzwO+0a5HfQh+WgbsyTIv0LpsTDkb
EQ4G/OW5ehrcqzqYXbEl7ktZtUQfwXdqhsyaaC17USbLnyzYjHF7wJO7aKLvro9R
sHegM7X7bG/D5ke6buB5Lp78VU9Vr74SZDfnllhMCQmjebX35FNon2/9ccRuE+Qs
lofxbTMjp/T5fwCsnT8KR1wpAzHGxELMMqhiT8KXtP6sBAJq63RzSNcbX0lXtQtR
zdUy91SfQUmiujrJj4Y584ueBJKL5uayP4DVzZyslwfErbA/c4Y9jnANln/KoGHz
tNXHt2U79u/jifq+WzfYcx78BqCXMvQ8ngxoOPBTMwCNMVSInrldg8XX1kK1frcQ
Yk8uC954g9+q2N2WkCYqtHzmvwQEv+jBCw5fLaUdrml9r0RSyUfcPVyEgJm/hcA7
vgQdVfAks1+aTCzKrfjCKyexpdtDxEM+4da5LOs45eHaNz+TKWnJGbkzv/SaNLRZ
Gf2QfK2rVJSWvPRHAl4n/k+NdixKhaLfT5HP7V4vbee95I9nhdOI9U1LllONY0ZD
lYuUF3HRFseCrEl9BTWqeMA8XjlTcoQge3gfjRwBqvKAN+1meOK0MX81QAzp7jzB
icQETOTVNqmLAhxzAl64M6ntFbZuB5B8BfD7zx3mxVQF3OhUifxCYWTVmuK67uRV
P2hz1ypWoTD8Ru1PAXI8QProCz+2z1k0VAF57XK+S7Iy6DfLbZf4wH06c8hac5LW
+6YzNgnC90qUPSt+qJs2SMrLRceIWaWwGXh190Zw+2uPYxD3vhw79CffIzNGqUND
6vwAwe0WzC8f8azM2iWG1WEkzCTm1VYzs9mHG6YagpGy3bpffAZ4T8sPvVEHSEHm
ql7hkGkuAJPCD00xgP/210ftGdV/fSXYgHnWQnbBbcS1dJ/5FQtOD9jCHuRMx6ZC
zVv08hpj1m9f3/dObcE32ejx3rWoywvdLA2nlpkeSfapckY00rB+6aADqYp3+afh
PMTjX6qN9TQw1UK4u0FtFvx/WR6v80Kts8V88CGuetPGT2S9O68YjtED1/NRUk7u
mSqj9bMW7q8oOxvE9gFkSbRrx7agrHU+j7b8E25Is1kCXy+ts8XFmi5MvUZJpgS+
h+mO3V2dZ3B2HSNF5SStmUVvp67s5J9Jhuy/+xX9DAOcz4HlVpvnwzAFNWLVd4wr
N4WZ8gk5CZonYXfVGt8fX2nhM/gZD/jHw7d7B5AUbFs9uKNEq68IXL04BVAzLbCB
TBFSlGsWeyI2+4DK5zFp1nmbe3mTggytL6jlNaSXoDhUX8jQYsUfeWAC/vsJyD6K
TOuFK3QbM8eqrdfJbPVTaGK1W2q0peSttdoeM1vutCjxYx3X+4ZtwPsagQ7WKAO1
Pi26KfJcMSx0DpS8K8GqhBEQcSkqFAR2Rydx9lTRxGBYh1hRNdYPr57PzynTmUsK
hjxjCL/1lRzCLvs/yJUdUCgmCz+zISJUsgRCspGaHc1/BvBP2QhnDqL1Oq03JYCD
UwS7MRYhCCZzh7m6Ai+u1fZhbLMnKfMjM9KPRtaA8zuSOUh3i3+RBJ2IfR+TdBoH
wuTUc8hspH1eck1jRfDZvgQuSnqC5Ds6bzYyBe6NGUUSJx6k2oANHq0GPgGm2/fd
DHcJQdPLnzedGzYlQ9pC5W4VIkU0H5KooaEwY/iBnZxP3Nx8W8q1PjZm/0qXQazV
wZf+64eJBdZKrUan4W7uqix6lR1Bj8xUFzGKl9e/PeoQUJEpFmxs85cgIi9+QWkI
mmas/UagluQ4AbYJ0TuLv7c912/IfUZqbFQfCL3zaXookGdn2JWhspbgTQBZveyr
zxwSTR363j3oZ87G+kkq3QfU31d4oSSjKVCALRoq+a71jwHM3COxmomxWBs6jVRt
QQe4fImelPCaDkZN2620qLB1VqfHbH0t55iTeG+/oBfUUMl33sVzSDMHjDxZRyns
jS+of0XyBL9iuTvltFE7V3qjbYynnrjXjZlwOzHc+in3nKoypi8mUFh1l1SPtzLN
fyVrrjbN4RFEf0BbWmbAT+JnbPm52e22orVxd//vGMNmWZ088adwEz/vUSRKH0O3
YRC81A5SgxPEUTJGSKMjhjokW6axURnSW6iC5shBNKJO2/M5a6JDwv+EP/q+sIK8
X2JEm8Rygv6QMA5401lL0KrMx6GIU566D8PqCG5wuNKhvAF0aWqfw4UzPfbKl5Dj
awPboC7vSwqc3P0ARejd7knR572NDp8GIgOjn83rEtxP/2Mfzm7ohUtd0fT19Jqd
yH64nRFKGRv4yJIlHLSkfg+bNqEnPE/JLeU9zwC0FPpMsTXsmB7lc1O7h3+gGNcj
3WPv/R4pYzW4lNZoqLuCpwtAvS4OVodXA3WJlS+ETgu39jsYQcNTDKIxqbYAriE+
ZcsykMKlAU1VUh4+KKEKpp2THLjJSBAgtbJrvXLdnTGlQrKcqlR2225HUYAZ05P4
5IVTaCqYAoxHnoTUslvVtmDybj6XG6nvoOS5HsHYJTzPqLDqVEhwZ1qsurlh0f2m
/I9oASbYtkxoUM9QQPm9vcx1IW4KliPpuDqPhXcDtC9irj2iWBswMjViN7Z0F1bD
BRrtxmooR2B9u0mF3RtZ8KweBMKJ0lwhGdJ+H8q1ULtKE7TFmtskXtfAV6uxqBZQ
SgCIJpPzbWloSk++oUhxoZcwn9SUZ0j5gfRQJRcs3eQPRGZ33ctZZxgk3shmZYrA
u6EyyTXyS4OaQ67sGJLdxTBNJSZ7xrtXrtNVD6X5Q2QeFyp6D7QIPlcyVX0xRJ7c
+gnJgVwRFJzoU145X8FMfeaEqYgiva3WWnNg0TEHbiTawJSYOjS6yTQcKNzSAJ4m
W02Vc75HgVBWcV40pb7mTOnEAsbAbc0MBHV56oSlZH9g4tSgVvMMIOUNW22WZLql
pU7OsPlJQMFA1uspfQH1fvRSKccbS7g/ey2YmJvBkUMYIlGwZgBPHaCxjn6TtGmR
60KzEWtzXRbEvGPTbPbt44oR1wCiwMpcHtMAcJ+emG7fb4Pg/RD43DkrxzGaRuFE
MT2lc974CwEJGGUolAiAxUsvKrYKmvmHxLuX97dbdoPVJJEms1aFB0MrCD+SaUG3
QvTRaZLSgM+1jz1teUUr9k8/16GjRdGshIYDkrL/Da71FYOunT9TyJiUNjopDag7
yxwhx2gzFeXFxG5yM0bN9oOgiFuFJjIdCUsyi84i23ZlDKNNWusvVkUNUJOeU/xL
udhL1nLWkwypa2qgzg7HazZyfbjQa2DMiaLrJjyD59SqgY5OJ1Ms+xjwxm8HkiW9
xnRBHbBNrvt21AT2PGM5cyyk5fwcwj3WlEIrN29noUEEokfquFT04vruMzD/I9ie
ccLH8uD9T4N9WD98G89sHAHoQGW1iEOhaBfPptdzBGfwlXJYxKMRqSNBe+0lT/kt
CkcDYWOqjbb5JJNajzZUpqlujj/1hQ9Dz9SwjBG9M+X6mF3ALO9FmZSNemCKam8Q
LC5NFIb6e1PVjF5R4YtGczysq6EOs70tQH9m4KDls9vbSoQfdLr34/SQy0jzTm+Y
X6AS/1HNMd7xO/Eu5NlBouBBjCmGk480LRX5rmbE8JGDJG7y/KqGuu8nJVFRDq6D
kBCIPuU//5qOpbMppj6O0T/FDBT70HWtIOpnEHd/wMyMNN69sEkOiztHlXbm9LQ6
K2/L7k0vyqtnfAJ0ZFUc3Og/kRVaP0+aWkHQiPiUxi1qu2nd35kEf19ppQAiBm75
eCQWyf1s2JhMuk0s4UlfQ9RVH2OyFGPUa3pS8Q7uY5C1rqa4Rp0TX9/fpPaBdbyk
otOp0q8aJn6waSISV5OQDRtUqcF8s5uZJ0cL4ZYhH0bDTWoQrk+ky23jZsiKYPIm
bIqIVvhFXZweu2tZl9uVfMnzpX7oAlKtt4YdbcmaxlilbLGNl7yZsX6IQiXtYgX1
l6BYRsLyLlqfN1jVx6kzlg7YNEBN2EH0z1P63cBGuHJRVitd3QsFhCvO0kPL9fqP
S0lLyfA75vMsA20qL2VL/39XRo2+no69nt4sYxQaeB4QxGnbLxNzDjNfBX4qOwsK
7rwJN4w94d2ueHCZpC/sX61N8OkFDmpULm01IAg4NvJIAuzsltKQWJeGsvJW9ZW8
AuIBE1K0sXsUkxzao6U9QCE9+RTs0nV3i2SkmE5kmB5RAhV3cbfIoIX54QbiJqY/
ILAB3hA5Pi4/f4R1WXcJ/YHGkN8eAGZmH5NNRvo/8CfJ3lIQepts+jSX2ZSGnLNO
/hLQfKcXyvL+NydwNMjSUG79GGY3UBr89StNTndkZNSPxyW2nO3Rfid9nsyMNv5I
f4SYvSKYXVOFdg0OvdTa04tT9RxFkfpoaj7JVMt0TPM5V50tncD5cPthpchw1cw0
MZN55AC5Ia5FGtZfhTummZvolH06/9v6JNvLhYfb9TrUvbwBPLAmmjW1A/gdE0nQ
ltLdbo5yKAtv5Tst2QypsjaNnPrylM7GQH/ztam4ROSWJGNI38Jas9DwvR2I2Dnp
XrBPE29eAuIOr7mibgsCJhMXqdDmsDWqaXTzHvxHFtl1/Ce71IeZtNQXl64I4XJG
bLdom9OFAE456nWDJaeCFKQmPQsszfdKeJXQJcNHNpGykO53WCbDt4MRAnkwGinz
T5UFnUCo/lGjXAWq/NWtLt91MRG7pr5WYwgF+lIFK3o7sNq11+8c4k/fzLLmTJLt
3FaW5XDKISWRqFdz3OT2mmoeXRW3EJOuBPMocrMYNyjj1H6RyAPCyUGKS0cHi7Nx
IC8TPUkGz+Hzv0sidTf82d+95lUhm/bh8WcdNkN4JnOa9xvJj3xoiIN+ks59doEZ
cBAGEtJ85aBWeJDAufl+U6YPe3sfxgZv2MXmJuRj+i3hwe2nwIVHkccIm5bgFVMH
Cg39yZQiorVPfd5k4qc0PunCNzCHWjGnJ49oPCGh7G5da0ij5uOwoxvSqMcz+QUZ
ANBsd+KpsSZ5TPTBwvGzcBquJ7qBFrzQGxC68n2fwA7inhXrsuEWE+ppzhna7PIV
PtrYF0BW8rX9pZrKU2+438dQMGWVWWztX6CgkhjRDCNwk9d9ApPZqd0FDf2RTAf7
cgHv9Oj79yHa6iANPmuOJ3aSomdvn3IYZc+uPL8gNgHlSoHtatpLx4H+m5igu4RS
YtBJifbAKIjkomVFy35S8LokwFzHXCZeJtjGH8JxS1kk4LgVB9+SlC72C8gVEksC
msUTDEiZmhkoTJhyedIGWnJ3TWrKyhX0F09RyKG4nUPF5iRC6w+6IuqJI/BzhoUE
Hubw2OKv/J2CoCb1P7lAXwh1Hv5cR0tBsZ0bPmtipXyDoBlxWjxaKPY8fMpH0V/W
upRSHqjY88sjbtKRCVvzXJB9NVr94liDDNnEM2fEqbNDLhFlIa1+Jxe15mIq0arV
x5nftK7JrhWr3H/HGmTuwMMeMeVxVYL5icGeThsgx1fEN1+vslFuZKNtBDhosRcz
qZ1IlaQ8jPlIJIwk4gkYrY3iZPd7Ch3/nHMPsfsf+S8pvdx1SmAaS/qTFcBA9+Dp
wWqoU3eoas6z9ZLEELFrwtT3Ggp4Q62UubUVIUfvwMWzS2FcVbOsbn4dcS6EEqIm
cKIAa6ff9FdSHrwS0Rho6x/NeC9aK7li+nGf+C10Qt6Twtg2vUXzOfHOnCS2DpEg
3hwtOVPne/4gB6Ppwc4dy5x3AIgLvTT0ui1lIXlRhLyy2M/ViK345XKXn0CefdEY
6PBWzCh7JbAW/FVMYLTyKCbkTma8vG1PKvy7iR1QF24xiVePcrnk3nGrll2gqQ62
hHlr7iZR7cyst7ojCVj/3UUQDLD/3sOT/NnOJbthbd+Fxffqh+xSoLYpR5td7yXx
6JMHl2jJfOTMigGfLGBCkuZTQTsHZO4XF0Fy7ztNJpgoDOzE89DDU6r4Wfkkun/g
XDlOvEJZdXkDjuLx1/9ccOa/flVQ+MqurKrUwOvgm7L3LfsAnXSt6zIj53A00qwl
IeiTPgAW8Ah50/CBw7/fQ0NktukSYO5kd//Bi1ITLMPgdTIY0UvGrW/W9083Jo9s
EAQGm3dIHWKTyIOKmSizBtTeOFmy1Z+yWfyEwd2V9Pnhj7ABUwYmzux8pMH3goK7
XTkAjW7VTU/zptRrsg1/Qsl0KFV+C9Zh19Hhz3uPZSz2HoIsPh3d46+RzINDXDLp
0GTe9yEPNq2Fdq/duzssJaU6OdjQQoSVUR/iMrwzXVQXkt/eqJyVifyAgnL7Am2J
OUb9nX6RwWdUSKLMItr+KjrgMpbO+Kp6ep/xTFkNxneG2un1Cnwb7h+RqmfGzK2U
Pmo4swgJFdJ9Ye9r78AVrVXYjm2+xFvMedy9AngvGuLuvmNKRXMz8ODRYVqxjkDz
05963/g94c9ko7HyCBFX6Evb1C/06NKGp/JT/p+eldFet+VziYiFZlYlZ6lt+zN7
7yqUGz1yOT14pH7sXY+9/aD9FS0n57t7NpaE/rUn3eqVNGe/pv26r2OnqPjtnkAE
hnBx1qkIIIwihMT3RNtVVyslSUGKX6Br6dDobQo/KHhComOr6PQb1MmjcQhnJnKj
rOBEYpfnSGGGsEnzmwO67Q+zBLtZRjGJ+5rGoNiuQ5N3097M1MGVx+xiAels/klt
R+JwRXG/gIAVJ5iuROp+KKGot/rt/V591UTfuO1PnwTpX1xOaGysQ2x89G7DyRKT
8lJ7gTB+Cr5d1eDpLltAZwz+U3hgy3pU/5EDKy+ULODs+z0cd+/p6ay/IpDX9F0w
krjSUzQuAV/pkuVa1MniNw7gca/YA573IbEJJnZ7Cf3Lvg97ARX9lGGG58rWAlRD
Vr2RfZv/jZt4ZpNrI5lTeubMmU8emfQS2GqDJtKj0TOQL5ZZwSRz9zkMf817H/iE
ocrey/DYi4OlcLV2jVWAZN4grY6YSGw7FzYA2xAG8hojSAhiq3RFukNCEOVkDgjZ
e3V2pAxjM1pzOEr1VG9CF2uXc2gs36h22/548B4C1u0HEMatyMHhek9Tot7853ce
gqOXkCUw8sV3N6aGIlPK+W84w17WwDunKbaW5K0fCArWo1Yui5DjsbKPUdLy2ODa
0n6DSknLI80uRuGNyiZZ2F7jD2CI1sTM4CPzlHsZYj0ioFLNz/v/pHTTG2SQ5OMk
uB/zcyY1tv8KaXRvmLhNEUbEQavV+QIUevqx/T/Ab6T6+m827dBPeSitK6VGbw/b
yLZq4bV30nqniMNjz2gKHaFfuNNMEiq+p6Jkw252mf2nphmTKCUQjnP/DBV04fzy
PZ25cKuusn4YTa76ZE7Ho8ZwuyqotFMpPmNaP+CrOVCBb1oJuOJe+fJEEBBlBHue
nAev65ndnZT8JsRvf8YXFUm9O++zl5g98M1S86FMKkun5slttdIhtP2F2AvIMy5/
GgMP0AYz6vxXckpJKWYz42HuPGIIRDfCCnghKylg40/k0phjQQUl2O+DSJejghSh
fF0+Qy/z+4hustzo1miHxggfdNZr1st6HBDk7dL1kEKYHnxQJASUndDTnkbJvGwI
i7l7voA4yvMG27vbIeOTM1bK7ehJq2IH86WT9SxmBTW+rQnfWlkZI+etsz7NZJqS
/WohFs1YwZvtimGNLoGPgdgcwJf0QcOO09QloDe62nlVlPU0dBvnrnpPy/0Ug/xj
dFsWAevyPAqhLJHUrZHemqJItC1Qnts7oWiZdU9a5nlF3LPwv33MW3VqI3l8Xro1
N4axoQci9GoSUMQyaDsVfDicvDgwdLZpZS1tW5fwh7pWsuk4hDOPyrtXZ5JFgrE3
QLz6paGoAYtj0emo8YkdwFFb2FfyUi14K7VA8WC4XNQ9LmsCVdGgAgPDvdGpE5ox
nGl8VaZH+fknOVH17i4swRVP7DDrDhN8UepmxWy6gHVn2x9ItbosnreMEIDyBiAX
ongDCFQl9w94b4rWiVovfXuv7ErX0ZGT77JFeTOMLpK1MxCVAWWA0Whr1i4so37k
0l/IYUqUSIDW9Qv0p90h6JucrHbJM01gPoqnigSoD0dBltLzbtKrZh9CaBvivsoW
M4p4PWBKcu+N7zTVS0vgokcS8xMZ3Ub3u68OTfJU+dHk06kyxBKmJqDR0Ht+0wtv
gpZaVp3UIrEXg4A8AH2v4B7Fhsr9SfT4kXYH0Rni8Z3XLw2vEzUoqyjhdzWxlcSo
RsUSBGbHFgHAWwL+yehofwgPM6S2VCX6gzRhRHHsColVTXyaIPtUBe6fJz688mM5
4CrbgOsfls0yneKuwpmMBdFekn8lzK/FliDh4bQ215nEh7wJLPSuBDKaXiKgHLg1
8k5wkF/MbkqsRCRzljvxoXOOZjE4pDTnF2WMF8yyD6021t/vFT09X2YxAc9js+uA
pEHaED5W+T5CqMew4yAZxKaCj/H4sTUhkPCyuCrB/CplTSNim0jPpQbs9uaj3zDp
vraFU+5SaonmFjckiL95UR+6TlUUndiEti5A7BHhK5SOPeh7atyc3cbvpa4wCzEc
BjqHOwtH7V0pqg9eNpoMPcaBYXyHdWesW6sP+cpH1ic2Scpv+X4A9ML6R4NniH43
ZFdWayGS2dRYyS6uN4CDU6x2ksE00Gf/MIMJb3DPINCAqbLEJujsuUP3pMuHEgE/
f7Zv+F6hwocCF9oRLXlYGjj9ac6KOLdaHEKc750nB/dj7xPWENxa8bl4RSEmE4KC
lCqF8BNGpcZhfZOtJqhgS9ZP0F/isnV/BlW0364fnkBcUkwgFe5asq13RdHzqjtN
xJkcDgGPDIY8nfxgxDTaDyS4Y4GKKt/w577HQeyktnKHP9o7fPEFCZFwgF6HQ0Nm
AyHHWLh8BoHwXVR1ndE/rRFszFiCbw/T0NUluYpwgosgumK/3bolajMrwghYbqeB
V/iT+GKmOcvkGREnbhX77aRpWhvJ9Pe1qlXQoFGgXitnW8hQCCm6rdISNLofu1XU
AWCbCno9/MZ1r2TzrzZ13Swnw56tO91nAwdz6nX7sWACKFqiSUccCM1HRK5NSqh+
vkV7V5BQ+f7Qy5vW1Y9a6o4M0d8XpYEyHBCwxRLsWHViJPxg49kBjl+c1uM+0gIx
MtQ4pWHtHxPPm3HJbpLtjPg8c3x4v4pF5o3uVEZ4qcVxm4ubMJ5GdUe8BDjOw6Zl
CoB/k6dnXb+zC0RL5yFhKJabRKlsM6Uo4kOJ1pahrzjeYuars1LnhNrr10sCQqsc
6UkZ65OQ00D8onAq2WLT2Zie/zezw/08l9hHwXX12pCSVkM8Ytjd8KJIUvz8GzQw
01l9IdiQdQVEYbzAFwZjULkMuuXfN7qZUL2qFyBtgS6NTrPt7M2TGkeLw/HBuD/f
OjGqSrP1n5bDxnG3GsIsTE6/57A+rcV/mtZDt5WlExPFOJHgftyCH1yOuhuEEV9H
82jmtjDuzBdKrifuQ+3UC07egVvghWvDGTe/VSW8C1weanL8QhGWBIyX65igEQzB
jFRkpruGkF1HcMtIT+w2sJKh6MzMR5AZIMdj78UenRTVNTtwUwOFedJa8rKTPDuc
G1Ab1tu3pWh6PgP2nGiMSWTl3Wom0jHH2d+TSdphj71vgCH3j2wwI/ZILbVPoaCK
i3YHcERFsr95ertl50a0KlDiFsmpl6t3alSS/E99RrF4ipujxDak5u/gebF21ziK
e69huyibw/Ngt1ZmlzsJy3mgmFitzE4AiRepTH4vivKr5WOUs+c5kIymoh4xYb/W
jiiuYrjMPNRoCitOF/lSieyPLQYorU1FVhku3rv+Md4lktoPwaPkNB52Hs6nB+Qd
u4UrhZ4ZGROaO1w2cOI8dNUARP4voThRIzC172v56fa69QTAm3ZGR2aBXH9+rvto
F/WePDniO3VF5sT0DwYIhjUjISBkm+xl8bl4mq5Hu2pNxcNeNwmeVUnigJmLeLOj
fUZqGPbvV9nzd9BTvJyz2I66D1sU0RAvk+wy4ZKUmZ+JKsTFZ2PP8bFtBSvk+iQw
J3VTQ/jBYkqSiOa2yMH35PYiuK2Ji6sTdS2Ji8c1BFm4y2haTs5m+arrFzZmgBiW
QpoqzFvQJJEfO7yFwYj78YRsbiwCyHVJ5WDMXHdLnFPW8TV3dZLeBq4HP524UxL9
RBrV+qrvtnhkcPu6oy1bLxM1cfgyG3u0LpeiUhDR0zD+5SMyjfunra4tfdzsLr8v
Olu5j1ZpJDTKRNtyMtGSeR2OkMgDxdluRbEEyHn7EPxqti5Nbmi1G8uIFmavZz8e
qs8Jm6GNPKccdqtUtuUQuVkItB6o/VyHNwIG9jWEKaerCF5UchvFesPHLfrBA4XT
Xp+n+xQ8KN7y8Ea3sUb/qyyr91NeevdgVZFTFvK2kUevwPpuxd7bGOlXuVgMt2eg
uTMfriI5+v3l95PQAC0jeC4Y2IdmHnriDS+4KRYT3N5925mK9AUGmGjUn2c9gK8I
OXb+KJQXk9oR+RwQc8+V+IZ47yIpMOeyeIhVvtIp2c9Q3YUpM0ZdFCV2XACKS0GY
kvu9p2+1Pj11K5M1dSoRh0K28MeRLtDJ7UJdAjBOTJRdPgmUm2O8dmXxVspcfC1x
mUoRoBbF+cD0lc+G2FN6arO+m/aYOWS4GnjIDLMH7hHYXO0F4bhsxwYQrGsAbmLT
oopZliSwMQwu19tPo8Moy1zXAv84pfVkB4SAHWNKn+B8ubSlXTWOy8IkbHYcVFsL
F/Ppz5dYSoQSJpltQJLdlfaL4Lljat6dGNpwIDNbgfWelxyD5k1ZMfw6FPXhisy1
nrdVhOlQYQJQA9dxEoQ2vvyJY60Oaps2RA/S8VSCxSm5C4A6yFqe5UVycAawo0Yq
EWETbHJFjKCU5273trD2MEX+jih2ZJ6n6taiWXfaoetgmlZe+UriEsLTnv7AbGSO
JVPQ75NHoY2bBkPCFDw4HL3aFRLf+qknhNIvnGbuBpDgMGq1Q1wjyD0r2f05eRc9
kHEL9xNv0XFGusTg8bm8dFBeZRuPVEiNJO8BAUMxL2ylArQZJN0lPh9KgMNZsOv6
Ts5rKehvqbelMkG1PuuJuvpuiuYGRVvDU2M9kIyTNouoArZFgNInhUaY/TZSK6JA
fI+6lzToqobqFNdU3AlahqOWE8x7FgKnQBqOdS/k2kO/EOiL22fGyyS6DP/rWj2W
gjDnT/5iCSfhDrGmdnLRscvM9jIelOq6kSYm0iDUt9zbXpyIcGf4Ao2FrQ+ev/eb
t7gK0yzohCoaoaAtRdV41PHBenXUjs6+qpI/YtBqnfF6qXVWADvrUaQBzhkFwHyA
RhM5LX/As9LZFKVYNcRXd6g9qsOJtjtvY+zyvQM210jEfpuYurHoIrpJyX76VQIY
cE+kyT3YkMsCRmmIR8sBwX6KqrlZzKTLOd+AfeA++z7QnxbkHX3Ox5E4GXYVC2ur
iATstX4HaJuVxWcO/rfOJBXP/cTxPpX9b2TdHhZiwIqBCsR3/+YOSmaP7BQtjUvi
LWNGvU6K0DWMlP3YkcMLnLQymZ1Pj59THnGfhFzb5eYBPXi8KnNw5YGREq6hIFip
aq+0D/QzRVDVewrK3cbdEdQK0IaC8ngN2RYaN6rK4JRxwFwh5NllQOsIne2AT3Dc
ALMsUlbiI0TmgdyCAKAzX8sRmuJhcfI/iTsLLYFVDvT0Pb7UZylbKefJS0nUHRGY
Rtln6HHM1IK4jGhi3s4BcJ6zaT5rdW3D84/rKf+U3sbzh46g5qwxnOqqeutqrUxb
gs6PnHzkZDjuoXlDPJk9+nTeJCs8XFls7fnCyPDdeb4P9nJssta7bStxrVcseSng
leoCm0KWh4AJbrsIg/pZBnshhtMinfmozGE+1LUwfDGxN+7dCtA7+d421T7tdly/
XMxytuaB1FN1tHeVhE4t6/PlTMQEyOCVWX1MsYxj3kls/FQDwJOVzm92MCXrxBso
qONW6DvUXWdBS6CG57/hUnCkQmFtb3aWwMX3//psNslEY1wnLOUDRvgbJIXKwySD
lLLc/JnePFciPfB9uSlxyWOKePQ+Agy5U+Rns+RTAVmEYbLLHazjaU2g4fJ2GGDu
+eOECTvbzifl3aun1BWzaf3bS9yBG1sNEo6K1FcWpV2BBOaeo5jNRbAx5Oz9Y8MF
BsV3fYIfzEkuL/8+RG/tnMR26CAcH6vsFs5gV2KgyZ8WkygLXGg0WIjdmGpGCxFV
wqg0IqGjrNWxV/V4MRnqwbCyYnXP3fCnbAXS8QWFk3dwIJvivhite+W3FgT+BNBh
Va77Zumi0MuHa4V2OiD+5HBjKvRwI/MxsqSBdvINagJn8itVyJlKrmC6pn7HTQbG
qPHhwAzoO577nMgEbJc2FQcyQan3hZlQ3mtkC2z/Ysac61uTfkXtI9+2rxZLgcu7
soBN4FpRDdbKpHdGK4unpqo+eYB5Dh1jb4WuVZaJUb2pHL+ZVSDGbv9ZfBlGkThN
gCcJrcMudc0HttRmKmJPkgHTDMNMwi5XFh43ccTnsAXuZ/ao3mG1G+WjuTMlm075
3KdYliGlFeW2paJeHVS15mMXkuvxsr7DR8VxzIBNMaJWgUNViFFCx9+v9cWZOzjX
KaQo3Q5wXAQ5IAy4lcmJYzhEwvwArHAd6DL/kmjdt21LlNL3NhIFR+HWcMBmYu45
7XWBRyeRe1DV2xfyUTnPbxpX3dmbjidF4obxjrvpb+HSa1rxEWT3D+v5JcEjsL8b
dejnONEJcC7UzpE5S0ueIl3dQDyzLdKw8BXZ+W1BLKgmmt1oG+0O8IsYSU972DnP
fBsXt+mQpUAOYqkWlc6rrnfqIJtPu6ZtdeFOQ5OSSuJmq49PIVcH41Am9y3nEh4D
viMeVZsesyE9dV+m206uQEU2qb+jgIgcc1CsBGXr9Rwb2oHy6+HXrdoItBazrWnF
Ig0aoCdgpL0d1wDjmvCMOXxxwKCQK8IaogBxIRJl3i00SxHSq8Av4fSJTD4TshkE
kVr3xInY5hLCmim57vMmYNeUKNwI3VZfQJ8luZkgdD0eHHMurHZaKSMm4v+aBkPP
X7xcTz6K/6JbEiWiGJ1GZjdBXtNwyrYs4rZIJixMxwPen/6WToWpe4bsvvx/6s6d
3iq9EMs1btJWfXEBqFk6oJYM79JgvQ/G/RXP7IMi3gkIeOFO5iV7kylvkMXzA69t
n6IezHR3m+vxp7hni8Qi5oKQKTxiIUOXZKb3KHi1G14YeWFjEpMLQIhnTJomxOOy
De2T1InSRGToQT4gsF/HKUqkt8ePXKvgVPdu05haFMsg44X4E+lgmd7Gv2lHIN+y
6HVO3rW8YAxevDxgqkntaMl0HVERf5GcN08HFekD05lF3O+WG7iA/NONpqwkjOpx
E6XwLpaPI1+xKQG7YrZ0c+dvrJHFI94lGdY/hTte2SfxLOzJjH5Yk0yzT40x9nXh
CMuHt9Hs9dDsvGVwcnCfepgixrVeJRRC+t4MIHPd/Oy6oeO5OfXoc4y8xBbZezM6
WkZ/L0QWRPclNrwtaRGqrOLuG2B5V7nSGbcnql1+dzNaD33zDNfyFvTE8wHX+R8+
fDWi/YyiXCrf3yy/rOCPr3WBhPjPlAsnNejrgy6r9wK1ZGmj3/2Ar78e+rORWqAL
b7LhIf4Ql+GYdHzr3EhRKfcaj2fPQanEI/73M5lQrtUIxBIp9b7b9gXxd1BWbj0n
VdHaOJuW2Sa/fRycZdgSvJ1/41ZBF2KU2y2HIheyuGQQHQRF/ebPtxnzN7XsXG7i
Xp20BLGxbug+xGLRw2kt9RN+dQDN+B3mMdMRk27CFN1WeycDTy0UmV8qs+l9o5SY
Z72fsIOJa+Va2uIJHb/WcnX7tvV9uSZ26EBhi8ZnjXfF05tZRLJ/1ltS5UHmxt/E
qFzyyl11BFw3bf6V90UNJPZivXaltAD5LqKwMYt+9aubBYcpfE3WR6oZBB7iUmXz
NX0APe0mt/IxBnCljvMnBiu2ZpX18tNZXjTmjMNA1JQRA9DdR5aoOyU1i2DTZuRn
Ary72nxda2guRD+FwBubb37P9tpWyGIu3HEaorYyCKHN/fk5xYd8ie0fXdCXM2in
OM89EBL+OiTnJnsbqJ5f5UZL4U1fhfXVfHwnMTo0envL6oqJohudzHRma+b3640y
vUgA5Nx7cxtpSQ+1Q6/sFq0D0XMgdYIFqFRrw/hT0k5E5iOTH8A+FdR3G24Leq1Y
slgX6cLNqq2K+UTGEWJRFEBUVII36NeRKCb9Nx9+5CL17H4USE02uaxxq3I99Sif
LaDDXLfnV9mIqCNMj7V+BmoPeCkpgcFqDHrQa73WftpDiSwzTKsGgkclbokIv/pS
poBqhGyCgJ/mX069OKjUIE/GdIEzpgWToZ7vZjwoVo1sjY2YWY/aZsSB2Iy3Mjx1
an+SBDozNrcAXwa7kAxBsG1cvTdyom93kSQpSxjS+IxiNeHvcr1LCeC/q2tyg8pZ
k05Hu9gtloLUUTnvRGZ7djWzuna6j15f/8FiC8dN4IJCqp4ZUMnk+IcQGFcb4tqC
MQddjfLsnKJ2G0RtHmkht0GLwNgFV59Uw5FX1GMQusYsaVblWVmbxsrT6KxLhox5
qokFjupltOmMX+Dq986qxnKaqMb8T3sEfqEwfUi7UhMxhZRWbUPbQvnUK99HovYu
BnnqTR7slz+CthArsHFeK/Xlldp/kGb44q28gfYZzNiHnGquI1la1JV6+LLorY39
ih32+zaYWrSjhGAU8TGct58ZCc3dLWtw9ojmEIBpFCAkEDZPeyI1LtZQgs4/X+1x
XUKhoLaDX5KBmQHZfczf+nLf4t/9FmCUbOAvqjypUVpNIveAhpHjYgA4sTmFapcK
ctlq5pYsbF3qenHrthd8ShEKRHQfj8FdYIYJ1yHoP4KHD8WT3yxcW5bsrDJZDU67
fP/oMUDpIifjH34nMad8abt27rQGG3nCBlrGSW0ULFq9E0IDR5SrBHcqcj5jLjzD
lHGw0HZfA1yBDa6pW/EBvkt/nG5SAjouykvWLkNQE/jDv6kq4GRVdiHw2xJJhGQe
nbVKAoDCaXP2OAEc8LuieJ0YI9FHrHINtU+Is7vxsMdK4oy1Ae5Tprpr81GjClji
VBfkNh92vQYE10faNBSSZ56kzTukGGXTEugplVGi2ivbdGdhyHn8MsAl4oBeUsVb
POcnUJ8/pxrow1Rp8XmBGUHB79KLeBPGsJAq7KzdaNrlrc/FFOnrGxRjWtDMLA4z
PWl7MU/wP0onKgzXxLyb6lrvfZarQ7ZTgIYlZwOSqTcHbSIEUimb4mYrfv52Dgg7
uZxqH8NtFud5tEWbFBFAWOAaZF5dnFpQjqZK+MEH/E8PMo6TNh+A1mPM70ABz2r1
xV6sG+fwUMVv5ZzalMFQF5VYvcvhCNN6pIuywkCsTyvVirkcZDedsx2W3jvKdL5G
iuokAzLEV829W2vJZkXpjzmu8TXFXO/FCAS2XQcekz4ykaAeywCDd3KIWXNbz9l9
cCADcLpdJUnT1WDCsVaL690QJb/12AdK55LvxR8AYGWacGx5MzapyBxnr8veLrmt
vqoaSYcsDZEw8dFXkeP/1Qe1DF7hGliEXz7vquBh6lsSYQ5WI+QtlEsV8xI8KzDm
admR2lYpmrBP0On7T4EemMep8s3Ipy1nybcgz5ynFNk5zxuwM88KkTiD8ZT8gZR0
1n8r1f5809G6uLTDlyjaWwYEh3uKfO9W2YrVtlxTBU2mp8ULioJf2BDFETELepOx
C1ksZ8Be9f58mHJ/OFWUred2QCZaWQNerajiSl56SUd/YtkrPSzFYJRF/s0nQcNi
s8IDtcPfKiZdjuk6H1f68f7/NUwpetx4wXf9X3d9rtf9FYVWT9yDJPFuOZaNsuMn
7cTazxq5WApYAAtR27N6VA/L8KRnVCaxvcmCt+D6Z422x2asMe8IwRCUY26r7Mrf
HMP5mnMtvOQAw5sK/CpQXvgEHi/vEq9IjCTJSSfCKGCra0iPCQ62SoDOw2XUQqwp
WkDhIYO03tyzapnyRHPv5jssNZQwaHedTKo07tMeAY0CRBsEP810TrJBMjPN+DoV
+wY02K67TLzfm/Ld8j5nkjClIXYQ0pJSEnB3zyTubaTUGdwAP47zgrwTKDzJmc/w
YdZUzTGdp6t7ppCl9gi4yUUvYW0cmlQoRSqx3Xa6mhEQNHS2uJGDGYQB+aWPzjCA
0hP+MkoteYgnvq48bL5wN+uz3i8SBUqRyzkpz7+dPFuBtQrxCR9nstKVprFYXaBP
fJyc6XO9AYTavm9/Q+5jyv8EswC7qtNnaw6cdboKX5BGiOpfyd4lwEsQR591UFOp
vwYW7nQ3/uGeKdl4F0kZwLIpgql1Y3UVzZVPcwDbjYT1v+ZUGYJrTGAQz5zOUJPC
eFW+ecOvxwqI4FAjC8Hb7LmyKTVAXu0Rz7G2Q74cuZnJ2IC9rqq1/za5XSl8j5NV
mNbPNhNN/5WZc5LMMkcFd0U1quKlW7mre8zHVlZWeJJaxE0hgAQVD3Xh6Km1dX1v
DIuefvcLgXUBm8b09lZtZX7/fR8QxtU/bAqFt4jSRMyIXmu9cAAQFgaNf6Src9fZ
5fQojGryEOtHpQrubhIkZSU2p+L72fzPGIugIbfPK1nUIqfxAsS/20qs9hm5TVUh
ngznJI+O39PldsVD81DU8ywOg6vJTE5dE495fdCC3GxxPyxhTOFSLQV9iaCyWJEP
ZaGr+HMEtX2iHxZJm+sCUqF+FGNy+I8En4FQQQKfIS7GAnRqzVFXjJGqoYex6WxZ
8Cb6fCvXyTBgnaR8AiNVvDgr8MSOtSFCAPsk0Q6cBDscoxaFwspnZ21CGcO9FdTK
W8+3ETprHoaOcAcg7VK9uf8GAlAZ03dTNMAY7KJY/8bAwh4AL316C0Q1qMOnGzSV
2fQQO+Rczwv0FP9gBuzhxdO9reyXtOIlE8yX2pz+amQsFXVRAnmYWBsnp7GCdwXa
4fabZHv9xejh41AmVq2EnCLuqovcUcKozqrdoq3noJ15N9NflewjntVD2p8V15BP
UBrB6Pn20+1F3A93jGrqsxb5lEjZW8T3nHu/5qXlI45wJ6XBirbblIhj/vc3G+4G
zTzomtweX5DiYBcFYRpenuPduG2r1oWzLkcUCznJibWmKQ0zOEEg6n8fUBQ7DdzR
BA8NFPsFWP6G8S6uRNLeHVRaAbE0pqt6wGBz0XJtq1ihhbzCNIU8P9bGncYcaTeJ
yvfvwAS9nwVSEbrgx3RQXqvlBGfKltrglmLRhqXLeNA5Y210ZVqs8IhDwHaEPEfS
jpDfwqxs1prx70AE85NcHrHh6ZtP7xfyeLbUh5nvxM3wrRxunAvoX3Ko+i9pwrDg
gPtJVkT8utKhJL0n/qC4dM55UVQg4sE3hnSOOW2v8YunR7fyGWUWC+Z5knBE7Deh
L76lwPkWTqCcFlHXMBqytS8KzhY7W3vlWrGdrC4psUuaKQjprFwX6BlfG3CZqUXi
xnFr/oViO1xXJpSmtmwAxQftjiza8G8tpOWDJtGiGku5wdxBb596xXuX1sk/s8Qo
O6JOPSeLo5JwvzhytxckB72dSQ7VVJNjm1JC9MfE16CeisqEYar0AxJH4JioVaW1
xz9n+Of54SUNdTUDCRT1hWACT5fWulBFzsQmwE6ggkNQfZSoZ3GuAk953CDACoPa
X8o2thIym99p/NbXi8q54A9Qwz4LgRmf+tLfibOih6VnTtnOm6rokMmrQKpq78px
P4txw0ilziy6soOYvVXdp7oDvkfUyDGQtK5mv16LtasP+Pnd1AoRkRiwFtJtxt1o
Zgwiex6iGiungpvxTaxIog3aIGQeJFm38SyLZ9l3aYFE7vRyxpfHvV+i902tAnlU
Ah1aOJG8w2vRv0UJCPLTP2u3g/otbh5eR3njz6hAOBDpmyFGMQS2P8rSWXUqQV+J
fdrOT6xxYRANMQKWD1PA9zmzEYrOuZcgVus/pOxLLrUGQIXNx28DMdER564TldU0
Wpw44cxE1tVnlDEIadk2rQFYL/esK0PgRL5stIY1lTx8H2kz2kzXSNTQT3BjA2Io
kQVaPTr7pbDVX2VWHNCLgPhtCWjOrUdFsiOIuZcXz+QmNkXhOQthwCwBSG7I9DhD
d4fSZFNFr1ku3/aF8RnjdUd4mJCP2ymWkY3s4UK1/xvfFa+TDgnD0Pvyljxf9bj4
U2vvKAUJ8gVf+F4e0IA1fINprPUrn0LE3k66CNtAem/PrrTYtg65SXIseykvRIeb
jkIPRdX1E6pOx6UeJFKlj3FDVfztALigBWOIYHMjyJzCiIeFydw7KxEvFO06TKda
KFatJxiw2NF+DhcDUCbDrVe96WCia0laeD7wrr8NuEtA0frF9RCZcQJsiN99lHk4
vNn1tUeKNFeuQpvv+RcBzMkNrc2e6mCtITB474Ls1ASEqGsOIdCfh4X/bvuI5Oxt
MJQ+9R2D7qamxE2oxaF+vVN/ZQMr5YRL1BxrGOEcXveCEjK44qLGkUSTbrAGxsNy
NDQIBs1yDCHb6oc7SbhXZS5y/q/HnoWZTgUuNejeLrBdiAhnUOVuOGE9pf7h9I00
2wepHSkOwazzUid3ks4pcg==
`protect END_PROTECTED
