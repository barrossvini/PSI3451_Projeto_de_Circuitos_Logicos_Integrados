`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aJlMtloUZxmaMGNWnTEA/SHPrLW8PrQceWHiH3GnmlOMgSVeg4oF2dvpVcvFhk5+
OlHUKyWysVep7a7dhFXfB8d1jT5aRMrWOCxe46jO5qgdimUhs30xPweBFTZQ/f80
p5p9GEKPYH4q1lWTydSU/+lZKIpsrMHPwm/F/dhLshvCXmPj6IS8lm496v4O4KOU
jnLWh5CFhKL2MBpbsyKKoM+mXis9d2SMmTmejLrUN2Jgu7Wuuy3nYHRjYZyYGQlw
yv1r7/+xqVqW0S4jo29l230DGkRrDJlIFrNNHyTElJjR/g8MmvH76fSLQvgm9iS+
ECxNHN7rcE/GCPA9g04hyBBRvLIhcI0/tavWxehGpsaKKgghpBLu/lSFkIvB1ZM8
wMEQ7jJeIlvx5NQQSs8V1YjXbvjk6G3pjfkXgU9u56zc7qyrXkEXwI0D91Y5vhTp
IN9D+tgNtRy7yTJz0cXd4VrDdoFShiLqSUzS+RsGi5t80ZPbHfNGysjI2Vvk9tcD
XuAET22R7Al1n10HB1QgiefbHxGaLZZXdaxGjGPCUUE7vihnisOtIB8Z/0mqS/EB
nm71wu+Nb4NR/rP7AvFv9zaTz+nf0mdTiBrKq6HKzgkT+lec3PB1Hl7YNIo4ExVQ
6D6sgnofiWgueuCQsoj8VsOWLy1E0mT04WsiTF/iB9aJ44ioej4kD+uZMOGxSaYb
`protect END_PROTECTED
