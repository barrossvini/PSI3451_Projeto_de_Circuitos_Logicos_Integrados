`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WDKbg1Nq1me54d0iiuEO1ZYfSbjpZ1W71ARb8LxQJK5551BszD/wQUonHzWhFFet
jyHU5K7EvE0MNQACWpfXG7o6IiOObV0DHa9tL1WMNJsZLXUEq/Ml5AUrOT2IqsNv
22yGbxlzhzCXwic21ysRKC35vlVzfKcF+6QIxYJqfpWUqVuSQ8Hacbuc2ELP2M2l
qbZ7PmVA6iBy8ifdCJnmNF+oXYD511z9x/MoRnFXccKX/R2EocsuO+wDp35bTxe8
iJzHuxYp7vBAl9gYzkS0+27LcarB7u7XFcMlx6VTyRIjMG3ET+nGzmzTC1+MaUEz
DKUQNgZvMGKmVAVRhZRusOXjdAXx1IwNDP6b/LkkH+eX96PDTD3Fg0tGXLMwJ9Xh
ZJ1HKxCq9DQBbhGZ/Ntc03IMrsibTnVTsjkudZvR61yJNh2vhgdjydP7CLncP3Wh
scNDI6HyTABzlVPkxmz1VU2Hm43wNCXkU8ugJFFJGt0q7y0/23u8klZ/181bpe1r
cjfYknskzQGWWlqD8AgyMYZEu49FTyjMQeHRbuppdsczJLZmB0FaJebP+68RK2TW
OjnQVJOC2KB8Cp9ql6ry4SmxqZDFWgITBC14SmO/1EkwH0muooHKB2SW1WtMCC1n
qvSWuXHYmrPrpN5rPbMYlYO9Imvutgp7o9dJbr4eUx85t7wWnVNuREVe/6btvgtH
43dG20o0VCCFoBCbImE1tIhkJ2A3OeBNzO3oLvtapwLpqs3d8wqhKEBi7qGtRQia
mdy7nxKcsztMtvjsEItAgw5Pc88eRMziU4j/efwcnIZ93OiLrhsAcOm0j1pd9byR
x0jk6m2bJfdH++p74p+4PjG2TyttLuNB/ivyvauHtHs=
`protect END_PROTECTED
