`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+SpplH5YcVf1tyNWXta+2x7OjORnZkkA3//sUHagtk4N2O3j/WeD6AK2OMYhXS4
RCVPHNhuwXPNTa6R/x3O1Klzn4GdLEJGLXnVlNdZkTHMfLffBoE9yaBsJxvfmHiB
vwxM5cxht4/2W95ofSrsI0NhNvJ0tDOrc4uQ/YpwmTz5DjgThy8NftcLihZzH8cq
pVcMXzgpikc9V2g3A7mD/Cj0V1lK50wf/esbYng9Kr7UjRDFTIE9NMI8fZcnnHzp
p/Xmvy3piv82eIFB7ZALxtmNy6MJ0FuyXMul5lllPsnkfjKAXJQNu23IkRHGWN1V
8V5dSu/ANkbjdzpEG7/D28tJ48SAigvgjSRzLgaZzhUZUrkDTXGK3uWk7ILgdklg
x1CkP0MmwIFcnuDabPBgeQSgAKou7nfH6t+l1xBGe7wIpwvQerrqtgkvUKdQIAvO
aI1vrnLnpItD4Y7ewm+QMCKQrLiPYGuIAlUtvdPgPAmwDmYUD4lPbfDOn/6Z17Vp
+h8m2WzcoPao5g5ko+s0mMozkS0sgpsjtKutlA2zuFNOzJqDHh6j8c/sGSIPdNkQ
pCUkvVDtAd9RgfpTJNgtG0e5LKCgHL9NOd85e36nOUZmFqXr5W/KGRrCs+hL3Qy4
az/EcdUuA8Iu/nZsv0r16P5j0wQPRpFlKXneApWGQ+wy+YtnLOu1nim+4sVbmOn8
M13BvbCWu/udSnHkU7+aN7VEXQ1MyNIj0L5yw1W0KJYTh6P56MbAQO8ML1xAUimS
fAhQJncsds+DXTyxkmD5UNsyXOP/CMlzm4AmZzn9bVsPf4Eb2fQoQmAK0vcXkcnP
v9ICHSN6rLvnXD13GXNb1LA/C9WHixQi2YZ8D9N7poxMKLSDxG8rF83UbdJ21VD3
lEO/PpWQgvR+FXJ4eeBtyNXQKe51litkfx2ZWghBf+H4uW63yDPd2WEbRqebkXtl
9//rPP5cJkuxbxHy+M8S0eNVV2roVT6CZEWNcboBSDPZAFWKapPc6SHAFOSBR88S
Yb2fV9goNcx4pZtgG0GpuykNcYug540XVyBoE1/zL+tIlaAOtOMaYZBEuk7KIgE8
1uEHUKH2jt6W32V4Jsza/g==
`protect END_PROTECTED
