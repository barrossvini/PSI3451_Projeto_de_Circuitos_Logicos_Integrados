`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rmh0ntsnlgPYAsV3fGZAhvxatwWcEh09+YzbWMolL0nuZ66wU1/gXZjkGq5Q0ss
NfQg/+3ZLwxlnDN5923zc2I0szKjSIyeiyRJvYVx73IfGER8dIfNHrZ6kYuIp5SJ
2hQbRjrzwLGWzhZQwxgCiPME/XzFs5klM7BS8smZ9EKLcT5by/UmtLH66cFmlzJy
WRQg6YglscwkvYqKP8YvOpgypxzRadPua1bgEdqBgDhMEvI6D7hKx/fRARDjartW
XVwFpiuLzR2sn8mg2OgflfImybchBNNTFUwN4s6612iNpzw3C/UvBbhUfRzA5QdI
pEpurgmCAnAmuaQMqu8vSJeM5l0KWrXADCzPz7ZPD9ofqp3E1669dfAybdmfK7hD
2gArD7bJTXpxLpStI86UAfp4BRJuqOZlsRZPh8jePFtR3FN6ZXyQ2eBII6VQtzwT
z1WqGHgGqz25b1kWHOYRX8HKHpk0L3I5I2L+72WDt/jXSgJFMiyV+sPmdShX35ju
xMjsYPh5SzswJwEd6M2cdfiqj7Vf1LwgDmBFVLxt6DnLahNuG4DHP6CvmrItpQiN
NI2PsRZbZ1nezhDnPDxQHCQl43tjJBp0+J3knWfoEF3eYIx20wpFZd21eW/3AjBn
R7BFQ7m8tKmgrXkl3R6sB0BABQ/rynn1MdbxOz2hmwRDIfpUgwV9rsu6Dc9Al5Ne
OPdvVonbQjqF3Ukh5FmLbV87rQBczdfP2UUp+6+9ArAdqLylvmtf/bMb31CvSzNL
/R9mEdCDwjNz4zZg0pK5g6Wl1XOmv6LSXVXhlgA41/c3kzcLxT+56gK1hPhVnUnM
Z4oY9wcs4mQlKw77eF2anecFaxMK1hwFgSUamXjTZdp1bTQBnXwW4l47Nd/5EukU
jGIWhB/nuObPtb6mLsnmEvduc2TjWKjNFM5+X4luC0c=
`protect END_PROTECTED
