`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WT32OoaP7MZaiAR0wsjxOnlXZv9O6IlgZfRPRUMfUbcFSFJ4fORldfB7tI9DccLT
jvpYY94llzFVr4GnPU5UttlRNUQLqg9GC1H3917UBEYXhRDEK4Z0SYcQnJHRuC0t
rBP3egsNNVBgYvOJypjfsinzZ2iYHbv68GK5XkE+GfNpcUmhj3NNvT8E3A6/EUMR
fBOU7dcFSmEyFwwpuS/ELM+Ce0LSkxlmeegNJoj08q74UTmXaSJ/Kbbp0/1RGQ4k
cdcwJYJ4N9PF1zgYDnNptV97dlSFxnAh/Ii89tQpWC0LBGb5L2ROd7unvf9ZXFvS
GrF6TVL0/+8Eqt6UQVkk7LoDkz4gb3JanYBLlIOKoJz5zS9+MxomcYbbMrWEyyMC
`protect END_PROTECTED
