`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OGXic5ljdJNoivRNsvtxcI80PGdm8ZhpCl6QVLtWrBzWJWfuLtiE67A6ZJOaU+6B
v5zbQvFhM4SSnh12D+46ZkpBrFNsRE72TGdNWLPFjz9J92UEJi+F9UIWnOkpK1kA
cw2hMQfk/fT8ZeBy665AKH7lT3YHjNbBHz6fXGJk+z8K1pDtoo8TgpedEUAO8NQp
B4kF29bGcpjQIQBCnmmLt589nqQSOJMRcEr8nzD0RdhsS63F63zGyd7xDvn8Zn7H
+xCyBg0FBiWwQ21mF0HUX0CJrI5xNKmwz/YLxnjI1f2cZlTHNSjUT3GcGSlIj21N
MC5qG0x82/LTHsKlmA6x/cTidrh/PsoKVLvzHS8qpzsiTt8FwX9b3zO74P/H+Y3D
IBBp7PLA+nFowOOw5mL01L+kuz8ReAIyODkMS5AHhbE0u0qBMvtJ9MnWu03QHqLJ
82aDsqDGgnpXBsiVxlkrR+s8obONZww+2veHI/JxD1UpQfdDaNjN7UhKGMF+E/nD
qL8Pg3Z1McajaKVLKNjPcz4lWFFz1Mxvc3BsdD2+NbAX2cjp8XHnbJvBHAeCkLWa
IPwVRcg/KeKBYKcR3vU+VdoEZSEC6SJ2RU0kv1myfFD4X3QmWICDpcKyQDqNx7uD
XECdNqrR42NjnimrypJQVm6Z3THZPZAinwbHjfbp/dMYmwvACtI//WeBiSzXz5i2
SUxxUHqmGxcVajeGCZlw5St0y904EAMF6Anf5e9UbMfMp0CEvdROs6+pMF97pMAj
CJruCo3ILqC3I8F5rt+LSY7nAhHYZZOkjLs1Fhz6Qc4d3lff1kzQs8CGKTO51wY4
iNnsIbo+Fr3IJv55KxGgNTY6nAymdQYc0yFn5eZkHpGuSEqlhSDJOOWPIqlcSgv7
BrQgbSh03wsqDYuzDmG1XOplc+GIKZSm7AOKlpq7x0DmBvp8eS2hGo2swuQb2j6C
0M74ujgVlxtxSEGdVu+Lb9g3JGNJhA5U0ms4a3M9sVkkRDKTKzBXJkd8SCb/eawl
F4AvDro0gzJce0wFiwDHJVvKd4Fpe3pC4ra13yD6ShJ2n7Y+tdn+wQ0J/AuZRYZ1
9161AbVBrKq5cCGZo7890uS+SvLx8QEYnlV4RBwSLcX1UKRv7R1lA5CNNzcJgw9i
dAfhGNocBmbqym5uPW87DI983RTikYsWC5nZbsNbxKgPIkV7b0biXVBzWkDXhntw
EYHhv6qcCR/Uol7XoVWaqeaNqGnqAlDmnp+a/fWaOXd1/fox45pTdpmtI5jxB8q0
GCeR6BmWPf1LGawvraXFFFqYoYu4fASwSyTpOIWZFh8+Wch/38oFhYOBWvFhdIFY
6MWM0CoGDOx5/GWR+ucrmc/B1e+lMt/mA/DY5yVeZ357y6Cm8qGgf7AUVPUy218U
GyI7mWWdtRRK9Fje7HWN7s/KNKOnEFT7oJHXIAabdsHnV1yJXFGQJk6+lJkKjWE5
QZnbrrrTjoymq10fC/XmFXQQvDV8rWLxLulWDagSKs/bpOk0+FnHKNbv6wt31omr
Sqt+fu+OWrtYsYAX/0E2hw75BodbJ7fKKBc0F5b2/MgcpO2CvfpQaOhbUzwUrxGe
EedtOXqdK94qCmCx5MwBJ12zKnbcilgVRIqFYlId3qRLpX4LmZEGNItyXyxpTYd4
CsBzD6z72+w+x665J7DvJ2IgI9TTZvQHxD4Rcl7U0qv9PIyoGsM2fX5F2qMDBbMu
9NtwBc8z0wsPL20ix8SOQ9hGp42fz2owEJbceGVvEqaqrdvRa2/ptunVGHrqYiQa
`protect END_PROTECTED
