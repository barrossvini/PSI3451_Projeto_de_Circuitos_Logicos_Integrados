`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTR9pyu2+aJdMoVcLXQQvTBa2Jzuo6xqmFYBeHN1wGEmxuVFKHnxasqmEKRpMRtx
epP0EUf8c0+FUa5nl1hSQjvPwSTGHHKlxx3a/IfHpl87OXE6xCrTyeAH1K68Pv0l
E9JGVrMlgS18i1wdMM6oBFj0Lh03qcxE/bc3vHSqzz3TIo0XtL4b3wQnxXaVSCvE
vS63kf5gSQT+FsJdgD9DkHSEDmq1MovJ9QVNNrAKKnoyZ0b9BCMeg+FtE/akeUMq
S2LFVCY4giITW+aeUFF6MDTJ1HcPyb9KxONikOBdSTEZlbLLtoAG4/5ZS1WmSC4n
tirnPYv4Vph/qp3lVVZpqr7WKOVkc4iC8Dar8N4QF3EeQU9sGVD8GHTdOb2xaNPZ
gELlyze95sYrUi/zYj14C/TSc/vwMgrL83vei0W/033+oco+dumUIcQMGbCib5YU
HOSZivLw6GMA8wQmcmkxTEvhjwfQDmS0q9wFWaDXh1YsO030pu6pwk4mCGiTB6aN
eT4WSEXM3kKYT2DbHHFzbmy34v+rzQ86qkSCqooHaZwFqwADEALY1m7ewxByPWk0
`protect END_PROTECTED
