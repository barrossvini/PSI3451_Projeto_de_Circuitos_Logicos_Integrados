`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zanQH9XOO4UGDwH+rqYXxgU+vL5u+HDT4J8D9i0pSAOrsUSNSJ7vkQfSNhcVGMSg
cK9VYy68JFazKVR4bWg/31WE71jfo+rcWfOzX42Q0mTVAH1syV4iT6beVSrS6eAI
vvYDRFN/uN5ysX7ujzIU9Um+KHGMOMtqUmAvuBw7z3IEW7/+lmglS0ztvRJCRBt2
0Kiw3D3JdnzpjOFK/T6n6xA3WpuelmCHK5LSqcZ8drjgrQF4deHhRrBU6vpIdKqs
jPgY8PwyQUZa7Jf36Q5ZSqgCuN4KnbUXpSHxc3Arg9xwa/i0m0l5O8uMyGTKlaql
QYWTIk7Bh7xYvjOeuav3Sd1YYcBF/5Tu6yJN95eOS/1dy9n+XiH2ixEMhsVTE91s
IDrvcAyGUQQsdFXp+sv0Ew8Zq+YDMGYzxID0tgUuBGjyChuAIK+3w7QwzVfczbCJ
N9bryRe7a3r1HGnCoOftyfPY6kF/KhPY5Hz1R6XGOfJwRLLp+UpbGgFCqV/ZZqYV
Xsnu3Qh6Z2AdGvrRnY72ZFEYISzel6TTWDoCV+Kfo8a6fR1wpUYxWcCtAaKIyOwY
psHcB7rYawVF8smD9Nf4P343NBErp5Ho3ungg5rwbcdhOJWs+w4Rf01y4TozN4HX
HFhbEp0s9OTbAiHthanKU/5fgt+4sRmJwsCQ8HQl2nzMR6M7S1iqThRQaPp8Bttn
Bz7CMCDe7uamBhuLjUNXXQjP1u1BsaWTPlEI3FoR8DPDr3Y79mCzOGZBcx2hmp1I
tqKAQfNW0x/F/0xoaBJAVzzj221M5BzGKyRWYoFRRiIhO/OYnRigVIhMiCG5CxMS
Jmaf6wKtukFWSCLIYo1QluqZ01sBTIPZL2cJ1mTHtLNjT0cy6gyQQtyQ2xiOKB4O
1oVUfO5jmEw1BJlERZDoI7mRWoYjPNt5vDsdoAK+//fbIY3VjoPqkaD6xjP/FE1x
fmtq+vHkXtGA/Y3/CpYA/+udZT/m0yIezR006iv2tS0bSPZHfHAR4xmwI4cow/N8
CE6Rh+P7ijSS5oxYhKrrHc447My2El69MLpL5s+Qge/fnpP6O11ajgRst/gdoVQj
qVIvCf2USe446alIuvc384x90bfXUBCITeDFNOTbX67CLAynkVIKtYeLxocO652x
FjJ8+rQFS6PrVQd6DHz/aWbtOSQ9UKpyIr+AEvGjQr9PZezpSEj7lf3wcy+FfC9D
4YtQq7dCbboIcHoLANP58LsvgPQFeJqCzPXunvI9QaRJzhS4oRZEpa4LF51Xg8bJ
nuoy6BqOOE0xTwcy3a+C1K3oWkIzin0WbUOv6UpsVfjQdOhDPdgKjKHPaB2oYrl5
DdsmdMJIJXo+btZ97A1LLv+/VcbsEG2yxYkohTDd1bV6Tbsg4EPbkJcWIMEsnUJv
voa1kWyBtKJqoK38v1Dz/MMWpy9V7OIDNG3K8IdLLFE0vA18OktywCjm456Hlymh
TO/LQDYvdFKvGV3rLZWzlP42AvOw57Td811haXztJE9mAYj+DfAHaSxHhlEGrenq
lh9HPur9g9LP7LZVCiJWmw==
`protect END_PROTECTED
