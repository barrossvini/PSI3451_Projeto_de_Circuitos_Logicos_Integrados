`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nfEqvLXyq3GYkGqPwL/R8BxhL5Q43rV7edRJ901BpMerHzZUChRlQt6DV7/F95I8
6+67nRYsIXPJuxS5Ct5I9DIj4f6gNDIvfvE+1GaIF0zSEsyo0h5ANElZpG4PbHii
wcaxrdRt3L5RFcmldR/5gStpm+gC1qbrKbMCmxdEKKAO8wtVlI6+yTu65Q47qJgR
1+JpHnAmTvB3IuRM6iUCaPXr093aO9cDYk0J7/Tmf1L7YxGe4Uo0wpv8hNeoonmi
NHN82rj5eLkGo9sdnRz2fCvF2skiq1846JlfEbyPsz/o91ywQkBfRUuu7zhsXPqE
ohd5qStSVM4shknug+rT/mJ+RgZM3aUH6t4+utvmEJVJLLr38rz+/jsejcSPY1gD
sj3t3Hd5M/BmAgA70s40Xapq3DdBEJ3uc12HFMKWMMkWXH3MgmKL+TubZqqt5Rqe
vUlcbpXUPFpMJt+pa8eYy04+6W03zOr8H/srZFZLAAJxgaEC9XUnxgJQZf4O/puh
x71frkB0G2njYHL/ksXFhf+j8EHeO/keT+A71skm4XAKt7rxSd5JP9ym/DX7noDQ
Iiy2g26ETiOPhMWJcKrvTplEEIvT1hbdpn5em+ctpZGxAXcW9cJ0M6+spAXsT3br
4NDaQ8H2c/wRA6PoAVyTpvfCDtMsPdtaSqmHOegRXH2Q+/MkN49ccLQ+9XHr5ty/
Ai7rzAK68AuU5bPStjTm1Af/MfjWWlXDfWKnVIMsKWWT9U2zaP8vdTNvpfqQbxMA
iojCQj8BQz4puBFq+2kvq9X1YwZ6MtNsXHMjurEI9IUJLIycNd6vyfCZ7L61gP3v
TYKDUtPzbPYipAkSSrALfv7+p2W4ANWPsU7ME+ed3p8U+hXj0tvB7LqPN691KWw5
44oLv/Pp+Niot4F6GIY8fZoKtBwsWa5Tmpd/lWZcp9P3Z856KwK7iRuAN3C+XU6+
BJXFzmuAIaafrxkLpXCvILx8Y9RTWPecc4AC6G/G+mSmCG0A5ceSmF7Zvqz04ohS
W9731OAtS5pRxX0GIcaWUGqEXuZ49l2xrbh8xQIx8p1SPGyNteyxQ9s6YsZAbpx2
Qlc9aZ4moiFoqwiNA70i5O7z3qBL9u5OW71akX7KIOGDe8feIk5FeEZAgNap7SQr
QTN5i053lbrcrDtIVZFAIGcKZTy/0RhqvxrGirLVv3mIilOWxeAxMpZKJIu93gtT
lUdhgkPnAlN6llO03qfSc70de0G92WX4Z+/PIaTp62t6+ZMXHh6w0ENi7L2nuRJh
xH9wHqXxDegfTV10cFYxy6V4UtMBwtAG3+Sf9hlqLQ4b3UZoN1zksrhaxb4SW74r
6VfMs8e1mAaVnWJsHpZnAMsiyBXSeXYQUzk+RexGyQtw8G403mzFGV22kCjpXZLH
XIQrW7A65pMxY3hnxRK2es0tWIiLI/x2cRhgeb+tFcLA2OWrXDSa0q/QCCcUCwJJ
hZ7l7FRAyF56fzhs9PzXkFq9ff4CRo9jMWrKZ/MrKh/+bqiCfqRqoAjBy88flPpt
/3O1gQY/AdTq3r5xjtIJOacWFjGWCTySO3hCFk4mAiGmN2Ai+Pz95mMm0oqFTHq6
BmexUEgDn776AUr+0wR1DInIXyruwJwyvVOc2s+HuBuA2e05i/UV4QyKPdPGixn0
/HguLwxXQIDBW4RGntB7VWxsGWjT7IeIWlEfbitk6Cl6nCBrHTqjgJyToxp4fL+T
hPdsq5bTlTTUp5y2py6i2uAEshOthYAFzyqaBKetpvuprk+bqHJFRbjGMQw+2qkr
5bzuZ65rv+wGNTv0yJV2BCxRcSJhgkOUqpOI7mBa39wUTcukMlP4736Ph54Axv0k
Hk9NJ7pmEhGzR11dCpaG60OgwoP9m2AOJWwlRmtKRD9J2CLUzTOAbtkvFtEBk+5M
4sx2/DjrkKtW+yrBiP1Ysb0z8QbQLX5v94XC8bEvfpPwY5KrACm1ATD/wXrEvLqo
yeDWo4Kvt67hfxsUrHq4UA72LXkwx/BGI1YQsP6rnvHJXpuIjoAWAAyhfFFYL1Qw
vil85h2FlqloAAEqOUGdg0eaWaAz7Z7Wroxa7EKp/oyv5xXPRppealRMTU8iikKE
sP3JvrFv77WQnz0GCnyNR2xQVTWoDZRhfBRPW68kuJDtCeB/Bjaae/vQQ5sVVNTO
vTp0exe+WOHplkDKk7MblvjWyUzGERLmCZcJ+eVSYxWPo6zd0QHxvBJaNw8Ollqd
WSEiB0ZveiiP87aVWiH1cM6waV3FJkxTLmmOiV5h6uUENHFeZEnWKU2mMH86oLCp
qL2gSbKdOZPI/o7YLSJyRnmxZAxZxJL1T/CWzBzOhkV7Hrq7YHoJXLb0bBPtZ+SF
36DNeIfUjxB5PH3HmUqrhJxXeV50jQy9Fc3yxjXyoHFgcNHQL+BxvDbwrlffPJnO
1MGLPp3X/MKpYQeUjd+uX3/wY4NyWXOYa9NEr/8Gxc/X1qAjfI+7MyIjvaXFEHyK
CHZmrYc6xdaZB96cVPHqQocnCTLlrF1i16E/EEgiTDPVV9idWV86xZxIj/0Xv+YJ
L+LWBNXbo/bBkI5F8MJW2nHH+tjP1i0SoXIP3me69B6Kw5nHlggCc57ijuhn/0fY
otmAXX79lhIEKy3EFVUfGxz6gi50LgXhKNbbxJOoUfXlkAv7ikHHZdqmdSV/XLw3
Z2kDoskI+L2nduYYbLvhEHFEDvqXxTnymgDmFCiHEqj93aQI+pNvEQTFofzhmuPj
G3m8J/iUXi+uBD2s1fmwrj9Gu59HXjIrxzzOsdFYh+kaJfpAHBTtlAq/qc4a9H4t
4dSJuwh7F6JP3ao8PB0PUVhPn0qZ/TTsk9fL6ifVLSyKqxgEgrVMGqyWZlEE/1MO
vtRhV3D217sMJZKfb6I9FI2UroE6/e8HC2Ofsq2QbNVV8MhaXobjfNrluA6Pf6OO
JawXrYxd9hoxg1QmX8rLVobA0AbnCmzwRlTtkP9kA4qutRQRsgdvCbKNLUIG+kTt
Hp/clYPwXrpxHXOQTN6aeLxmgYuOvtoDTB3zohWFbdVt4PpURi6S4+01//F0W/Jz
0uQl/ECJPFNr/HiYq8W7CT7vsf8n9a/iH3WtHRF2Fr8Ho6IH545lMi88nh3gg1D4
4rfQutXdzZD9DTgngsTCIPRIxNB5m9syufLXYBzPTv+ZOiqZJZdijZZtv2BJExdo
y61n4nAzSKiseM9nIlPbRvgTDgPziEHcTqiOCzOEOoyBz4+vlXRRrGOr2+DiPPvZ
Uftn6wx3d7bePh/UJRx7BvKcEKMj/rPLzGJpbHo3YMo0OgLUmuuRicb6n8ZcymhB
cz2WELmvzFGx8OMtDZGXmQNeXExNJhxeaa6ChIsljlYe9N+T9LJ8xBTUy/HFjnDR
giw+rvV747dIqBJZMYyI0teqCN0rJ7aCq5IJ+O4u/KzTONbL+tihrzQVJ7aePjGe
juo6TthpLkO7GU+v6xeyW67oWjF0NrG4cYdnxy5jZ38CCD5KVvFWhDgNgGcLVAw7
SiN8OBd9Nxk3qJtXfVQ/a5jw811oit9iBTZVgszzNRtHNuetTi+QeH/Ltj0wA37F
UYbW+RrZVyIL+JuyMY+ygwPo4rkZROPBUqNIzs8JG+CpN3+LcbrwV/4jPNWyL7s0
TZj5ew3jJtkY4LIzeQepBmVFXzNGw5KtbdnveLKnWmx0PWx28AV4m9YUmMC2Upk8
XTfQsbFSihcSIbtQDk7+O3z3WdatK0p1mI7ID3geeBhIlBfYk0ZDELKKg70J/OIi
EIKVzclwTIb8d07UBnCVromQJiSwbG9ab3TMYPc+KRp/rWPTcaUXVfMXgoyVs+fY
MaS26pQQ9Erh2Plt5MoQswi95az1jjty7QDlNeYyHhfjH+GWAvFP/VUV5+3bwgA5
19ypG+Nw5nP9rvTUtALRpmEhgtXoQ06XUOsoSbU+8J0oQgsQUK7vxq72zmdAin7c
bZMj0pBVCWPF65yiQFdByruC7YkZNv+kuHRZZ0iDbMVOJgJbxBOIA+T8D4JOUXOh
TDgAqOcfb0ro7wZ0ixitdqyvzEZKr2xgAOdJZqb7yH73YbmkZz24L2kuJVVb5Pa1
vSvjUXAF5AZS7wOCqo2+7tY05fjxW/4gPTckYunjoH4p5yupDr4V8iFpFq9o5pQZ
z0Sc5zIACsgXwNhDWo8ZXDaMn9bGayRcWikpHCw3R09e78qw9R+d8/PDwPNCVWpf
Kvk24NitcmnhOi2yE9ACp88i3vucNHcxPhbNXEoxjNnkik6c8PFlzpL1Qt01rc3W
YCELKU2oxnrzrs0mOonIdkcIegl49LjxPuAVlDKOIpBQtMF1CuSE3UxxLacUOt0R
26bCdozwz89ql87JqF4Htsv71VCW2HOCebrI6Praonk2ee5aab6ecykM3s+DLFAy
BRjATPutrp7aTn8hhEDTeQmiFW/kIraU7FSp08Cx9s8c9l/miWHe/EV1eLBAxTUx
zphZ1weRNSu6ZQhMJ+7MoKIZpmeG06nkZ1cGRQrvP+xh1dKRj4RdYzZOyNxEtZZu
jH8jDPwY8SbSaYRSn2VKgRuDTd9kqxh+VylRm0Q1AxxTcKbmsNspIdIiEXMvrOX4
AO1bHd39lD1wbOhKdVXlHp2QFmF+KUcFGVoEtJUeNpkF6N7KHCgnLazOAaON3Xi7
yni/Q0CvQoI2EMw6dgON9ZeoMyqZIkQIG9rhzUnhr0Ud7a+PuxfS+g3qqkKWVlPZ
24yNzArLkeSs/j3ud+cjb2PdzkqTIuRMvW8uRuzy2+76ZYBUs2U3/ebJ6bOEFh9e
pg6jaJp5hEV/Gcmf+fP+RBd1N0tX9z4yIoKpm8imol3R/aDQzYtCXFzw1O5LaNkE
j7edOzifmFTr9TKNldaKMEys4bsurOyujUu1GK2CxveLN/jwiSNYqNKufBs8LIvj
8rpoVjMMUFJfA/rmReLB2RcW5IQeBaS4RKmLeR9CLM/U2JAZM6XMjxbDjuhB7qlx
/3d3mznNVw2cq4/KwhQfzvwrP1ad3pVJcwpD9JQ3V7ch6sk4an/b43/j1FyHgiXM
o5qwcxReHdhYlMO2XPs/hQ2F0D/KpbRpPnV5t+hOWHn20ShggljGnoaKGjzpZXIV
Dwx/cpRefxZOzNhhcBMC3004S1VvfyyUi7YS4ukraLxpRZSuiqyV0PY2/UIj6bxP
21aEMGh7o6gBb4VI10kvjcBZdlXGQGUAEAHe6ES1u3gwW8aBpSXHtXEpA+3ry5RW
g2slsIE4kz2Dznvmqp8a+g==
`protect END_PROTECTED
