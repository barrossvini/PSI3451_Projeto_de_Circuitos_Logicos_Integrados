`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CyyuicMJVDtRVY9IXUT9pi0RyPAFUSWyeVF3ZPZ8BBUSSAnmakwQ4NnmBy0ge/2m
mzZ2fPyqOa/KDZhUkuiY80T2+hjSpaRa+zlr/gQ8SLrC+g9NJ+nvjSHDFUMOHx2f
Xdq7EegUp+ho68rArJUWY+E9OZvld9TsLY1JOAPc34PCJQPOh5+J6+Sif5ptiVk2
Gh0wc79xX6xya504J4MEXsomR6MTF0ZTv0iJXhTZ29gfWz+03SS3WVCxM2BqnUwQ
5K6GSZfzUEkjhaX1JxlnJC+HoOn3EFmnesfM2YkKLFlQfHZ58TcR/jFwta1sUUvY
HHJijvYO99HHBidfVyVXHAQLcYd1djPlsNi91XvYjH/dJRhudcGxCGb1Eg+YDU1f
7ETV6WCP9FC/r6Ah3FXMFIKIU9/BqBFHW28An3p9W5hUD52qyVvvxj7gSNpZoejI
szBBqFoiyVXmbXW8JKQr33y2ZZ39hynR8lBj3FOMG2g3ZCjV7fAO0luL+EBY37Tl
`protect END_PROTECTED
