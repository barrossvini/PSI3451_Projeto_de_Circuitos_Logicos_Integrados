`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Lz6RjDMMy+nG5FCrbFhQRk8kEvgLFHJOfNw0PkqPMlGdqAAfZ0Xdg9y8hqTcATk
tdlPVDTaCmSnLxX+b9o857sY8uoZfDYfIIkUA7NLecZ2tCQzDqNmHSX0d5VY47Py
5DD+105TWRKCsmTL39LADUgHwWqfNVeHi3DgLgNDZZmhTj9pQ7o09ydabNZtaDFN
f6KC954GeHk1NQkKZArNkCUpAH8P+lAwmzSSCxsbbinj9keB9zFiqvvyy538/A6M
NN2rCTmhNDumt5u5ly5hYU7gemCyfnBYqgliPrJAKdpHp1eiz4oqOP9VY0eJpfE9
pb820Sjq5V9AAzhUg6AxoOPCS+lCrSX1FCfy2jhY8HJPhU28jubkNZ+D5phmXPAy
jK1eQUXy4wfaCY67ayPw5jsY+aOYdlH6kkCyzizaYnajexDu459ERgPSVilKvPDl
olWsur9hQYCASnHcJYLeei0rrSzICYRW7g1Wx27EbHiy3ftMP7SfM5VA3dWBo6wq
CUASYqPfWA3UwMZ1XS74GxjV4vEzTXX0H0Q6FglRPUaT8GEtNGjNTQBhYqRs3AVi
ITX/wZIfRKWFM3VNapiFDIydTwzGpFlf368gpXJRfdrAg2D9UYYkczNsVDmutRqy
Z147jhM+LXHix8jpooOxmW8SZBGwCdZfiFEl/NClTv1ZOlMFqQljbm48OUP4kr14
sa4tSr+bM6X0byPsWdvoxPJMD+jucy+gojZ3NpEY28TzBDVc0tmkA5iaBYhGwFkj
vmDqcng5KAhMa4ce5Iqcv7r4yJUT30gnHNzWwBzH2gZcR06dj0DQvlRJ4AZXUDlg
rAaMj7PtYPPllEkTtfxIumiy0I4oQrm32dSQsvRlXbCMavU26QFd34/uXN4FveFO
ATPfREdqMh1rGWrYCKjfVznQaeAOyi1CzCBoBuuWhpFg0H7iEg20IbB+ivIqYMjN
W17QZYdnvhIM3sXJn97Phon4PLEaREfHa2+ksEZvEgz2uGtgbdMn7SuzvxYs+iMN
Y6XW8+mTmi0kozYOcupTpbuWjG/F74wMYjFgqD5VO1TljzKEZCSBdFblKt7bW9Gh
ceyJmTuv+mnXvW+pyBUp/s5sLoMXxujtaQw5FJtH4p3zDs/3/WGNURkJRAsLkZcQ
oDW8gFM6GMnQ6aurKBttrUa/E4CHIvR1TPh4KGlF679AXZjO8SXIkzO3Y3z1ws+1
P6BVWqRdYuNbURDSDfUZUKK48nSnh0I+Cvoy5mRO7mfnJb9iTLBVDRGW4rHcAecf
ByN7ChMjQX4BvRgaqDChv54dlCWQffWxAkQm5JOThlip0cTSMEdSrme9kNFnw1VT
6m64aNPNUVn7vi/WiM3NGKN2awhsSYb3h/NbnITs4w7zOu6LKbjIcY25Ru9Q/X+Z
gnaamsJwrTWmzttUI3ubGT/fUXSIxac32NOgb+0B7enLYUjtUPv1GUNR2gCj4r2r
BvZpdegrmCYqefTHSw2TYLWtLAyGYaMFHROCK5ovTzR4WKpZkUvguYPq5ZZJU0nU
kbAaDtbkYdiERI0GWdqjKfbzRJM5RB+shW6Ba1nyPggs3XPdRs8s43tlL14JhgZW
kIdWoYfGq7VRWoSlc2Z1qshEFkQZHNDCvXra42QIKk5tgg7tgVCxOof4NWrZ2HDL
j6v5spP2Std6WO4Qa9uF2UkmgANtwwPtgumM0918Lmkioc8u5MH2V93lfxabH5Mc
pDIR6IGZ1o7Ig90cwWmforMm4MBGQfE7Kw+5Nkhz2YtQVkmfnZxvb0vXhaDqk93d
I4qvPVjKYfZ/dBCXcJUjB4k3YdCdvmW1of+I4VA/6oywlq8m3nwvqEmNclqGFqlY
FXTVUlFYlc+oSYMbDrFAJrSjP76uZA5UK6X1OLQ4PMgk+X7vdLhn0/Fp7N4RVpwa
sTj0FVevCwbTC89portW+HayqSF2vbG6myVIObNocFfoOE49ZhEfxvEOm3LYgmFB
YsVWbiXqHpQzaFmTYC5ndPVWfKmlXdGa4asHRn2t98A/rQQbapzYt5pUqm2MPIDE
ps5gvt9IEUNYtjF9GZqIG1SKtV8L2hnuNOttiALyn5LPSaWca46j0/sjcxHoNZs2
ymXuxMr7amI4hEruJ6A8rE3mEOhcp/3JNWuV1wUPFasdulTBOFfWqhLJrAWQVaiI
bb4cSTM5puvt2u+qtiP8GXdMN5W2gXNxCVXcSwAZ3sGLB0dpmjdTnRAp26jkivFw
YYxwF0KV3gTHGICe9KGI1vN7lD0zgiZLsqVvPcesANigdxXuAomdkxcV4NpD6OuC
1IIuWZ2W8o0Z2lK/Xi5BUQ6z8c8Z2aqbH/UBqB3JgHyE/SaGhq626g8d9qVXToFm
0w+lRidX2ZiRlxveC+XcwFQujIDXs3TZ0hP2+Quo/8HOJwb8XdPmbjw7dm9qLsQW
Tq6eyq7gii9p0G7GroqfmAKSYCo3p8AXP2hJi57HSPIHzdeufbpjtzGQOGNXJEB0
l67xjwhcfo5aez83CP0THFTdJwmShraTH61yUHL1//De7WCdidowWgnbQoHTjvi0
P1rLXPnWl67s2SSkWqz4xORZEkCaafghfFmlX+lvBDSvh3wlOUnUqyRaPor6YdK2
l6Nyp0hDRLlsuCsA3Wc9hcNdGCQjNM454LehkbfNWddR3fdIXNsb0Ozd7aHcZR+5
xVQ4KcPyk6NxHcratSPjHof0fDqdylZUWBBSz7V5b5qDl+XeXDS2USpmANGMFKdX
5qOUgkFpwi28KJRx5fdYNuHkOrgCJ2b7qTGE4GHHVglvPM8xPM0hKCXZDzga+BaP
rzWaKjJiPP4onzQtOa5lY93myZB6mH7ixJoQ+o+JUrU+RZrJK8JfuR/saPtXo8F4
34bOjnMhsptCVXfduHGeN1CJKS7EdlHOYrQ7Yiex7KyujZUMB9NpjQcf9j6jbShE
kzUhy+paWBaouwC128RsZDhSKEIez4MIBeqAIU8oXX2t319UJ+gD3SLlHaJWQ1Lt
lBT0ZmfBsU30GepHxvDKAbczGu2ELpRapVekZR6zoidv8LAAhRTvlKOClbLR34/B
sYP7mactSvHc+R4MFmEVsejVvprDpywH9k5/O01x2ZsrdI2Qb8I84bz6nxD6cWZE
PUVUZMKlAqMzn3jejP7bziYcXW+x+XbhSFbxM3HzcERlkFcV7ao3togqc/HgXktS
d4EOnS5FGXwMcgmju8BdXx3r0B00CtipYDPtb0jWr9kIb4t9oqBfGIntPBpg9Mtg
XhLmapHRLJsy7+NCQk1MCi3kKlnxtXXyseLBjxJTBfCcWvRdKHb71Dpozzs7UjHT
JuZZCnF2yUQlDst8wFjmZbIodhrEFbFnGmdn0z0q8IcWdORzDWPHLgYxgo1JooQM
qREUwpVEJhan4egTOYHyVT8m6rzPbixyJ1k2MxQh6fklqfaJNxvGjqfph/Sd17c+
yF+/iZ0n8HH27J9WmPJZ9E9pD02RtF6fHTxxOvhs5rnqiEIIwJIGz/VwLXXPBkQk
0CSvUvK1pzHf+POG2y0XcS/gf3uH410PGxBWdBTptyoI0FRyvNt/FRU3Ab65uMcU
WgJRfPNkzFFENPKAdKGgE74Y+blbT27tMtaxwKdkPKi2NN7CSGoegWHi/iNOGtcp
F3UJMm6AChF8pXdtwRoiGf78aWeG7p2oaheo1Q0CIKQpxmw4fBSBBbtM6IbYU7Dm
G9GVaGG83FZiCOHSatH54ivyAufoRy7H65gMqAkx0S0WvVGIOX3q77jO86ID1/Qc
+O546cHlON9lb+tPkdPJ/ea31A02Gp5zNSvupzVUv383BIb/VLAOhwMkjMP1y+IE
RCIyruKy2tt1D6Vn6ArGB/tQCKOYErIcObH/dAJ4Skjmp35ycoOs1CbzoIHn9SuN
8aT1dpkuC7bj4PFzcZ67I0aJqOtOREjNvho7XfjxtTdAnJZKuhUaz3+Mp+idwsjx
BsoL5iFSzlVOxNd/Ovgf0m48o+p2B6bodUw6NeI+JWrOinEZOysXMystWqPB7ULR
pPgk4P+1ULP+AAN2n+I4+0LxJruYAnHOT9LrgVdFyfN9GhHjwL1mSaqnV0Al1vlX
FJUPrf5cBc7gSc+c5HRjehJokEhvxescbUIJ8CB+3toFPiUQI1+oWaJcqfxwSNH6
TbJm0sYmhEUBHIczYfHSFH8lzQvZ3qnMLggoP0GmCsVJX8epUXUUk53WJSIq3EIo
vmeAe7OusK29eXSdua45bjcig0BTbruXsu892lkpfjiQ8XqgOAJ9gqwpciuGkYca
KniafCW2p4IfL2peKQg8/4/wwux1qlXk1a4CDoECPAIs4WqAwfAmbz5ORTBf+D1R
D5ctk5LZZz/Jw8Y1Fwp+rtzzjkNxCBmFmXCyXzyz+TNQok35YaNxGXJZUq8bbcxm
GlgXuCp7qfvBezVryDy5CWKXD/Jeb+pRvVnPoF0Bhc9WijxSR3fdx654ANPKtv1N
zgCfxXDxWCCYHh3HtnvW1Ijj2ANwlBUpvRsUpTL6/Ffo3Ks8T1nttRHUgnquSE2B
nQ8dUGls0/NXoA4rlwPunez1Ppq2SXneovvfOY9nykHI7FnMkTeG9+vlGjvpbSUa
xxSYg2AISR+jbK3I6RgCOSYOYjio2z1RPCT+YpNFZEkx/26gXYwFKDwkhPWdDxlJ
G7eY83L/TPdrCY7dR2t8mdpOZwtiJHNh1ytEKkF8ad+rLwpUxkOWM8xwbe24eCge
lGPbD+Awu8k1m64D0XhTwSRbPFIkpzTLLHdSNnnyzqGqId22uoqIeYcEsxUTEg3P
vNXuXrnFeft+pVz60vcPKelOIbpJQRIiPBofzw9eSXky4yKK/A0Sk99X21te8mvn
h3mySRzsfYG1Z4z24IUt3y7SbBRneS8+x0OXebqQX82+7vPAVKhRIETJdNeOyjP0
UYcr1ZUetfuRZ3r8mY0PrwYm/dA1ZrkMFAH5Me+674X1FBIAA2OcUUXlhzr3F//b
sCj4hs2SoR8DhxO1tdTJrlyOu3DaXYgNEJG6YcKacE5CEe7Iu7jvl1IlFe42GCwD
PAFyeFlD7Q+XLGDnL1t5WM5RTHVXux1u+4zYK9xt9UjzzbDifZg6rNB2KiOdCaIA
l0y8hhPQ7SNX0pANf9HaOhdC2xOphkzFUssCOeTcBWt1LaKvf61ynvmq+dipjs1x
UC6Cx51+HIU02t2n135aA10Y4ZA1vahk9sa2jo4XImKDzsUXsZPeSjBN4qFPyGfN
rj1w7fmvsdsHDAFyZ18g+9Ehq8khd40cKbkwZJxX3iUKWmPgnO+a6Uu83jLIsW9+
irEbVMns4YuZ499KF7HOuX0SyiLOpat++hhyXHjyh9+VtIKqASn8WTgeTR8Jc1Ni
w5213alRiIBaoPqxQy4daPcinR3zYO1JnErwfi3EhAzWZuysenvl1QngphyNk2wC
73XOEKN8yGJwz+tqpbunA3TpoYgAGhKmdkOgV5R+L+Gc8oy/YwCBYwEW/ss7iL9r
Lz0Q7JwlLX3zzBJ6Q/QWdRwwqpatmNo5cD1s6PoasiEJHJC0Bw7oTJt3AiJ3GTBc
x1HDzYCRrtj8ybnWXfNWNHzAZLCDiiOEZpSahpqpbAaJ3jctxYJ12j+U+KRyITIn
1ZTLXkMkZht492QUT9Lbdn2SlCfAWNpN+R49L7ViQOLfa0Uq0wXnF+VRIW5aiNx8
dRrP7NxGKCBf+j1q+1ZJ1xWx8pIkOjKg2fvLk6vFUyifnSD639mQos6ammzjaKvo
lEHg8AolCwT8L+08+hc4+9j55V4MNtZ0LGe1VAmIWU1H6JvFg7vN5eNGra6InuaJ
lO+wTLm32/jz4cj9n7fF8v6w/QraBNgUJWRRKblrkeTZpOATt5ufvJLgz9r7ypXE
MXUnryFqtnpj6LmFqSqCottU1m46OWf1/Bzs+5Ee4Q3PZ3uPD4yrYMctQCRZs9bf
FhsiJgJSBVPqei4HwEsb8w7ZlEw2dvgU8KGAkRPMbex+CngWLImh+Uv2X36go3k8
9nWrNhdA6DPFcvHmyLC8XvF8R/hwLb6uSNp5jZlbo+E2tD6TrM/nKsjq/vS1uIEC
boFiPGoBDQG1xUhJpgl+eE6OlFgP/VeQkcaKYV9/tgZNoP3r9pAWEHgILq++Hphx
WjDHoc8OS1yP7d9WOoJxoA5wPih2vdWYlYhiJmm7+sPJnX6EKEXHb2ibye0JyPFB
CJ+vROvYMDnN/F6t+0k1+tihqwZATZ/OKt6vueDRHuEeP9GhCkaspI1upgOtqTq4
/fei2GOex2XMgwkGmHNyN0i/RGC5LvOpRmKsXn8MiQ31mDiV4yxgFigGJ10PoTWM
55f3eJmGZnC4y7B0/i+ayUy9WX1KdFWqHud37RF7zmbsZ7EdQzv7frj87/YGKHBN
IddNWSyLXZ6WU0xoa+XxnvCPv2fo9mwPh+feEVTCcgkGUfqIojVeQ18G2bzCnuhQ
QvvpZ1ccDkZ3DKvTcE00Uej+2RnF1HYOoP1OWZIn2v2NRRKneoOHi/HJt4Fz0/qN
zVdG/QmX916mxbEjpWR0fWXAc0UGmSmHnlErkjMCq1p8a57G5bqdZCQkdvUGF0Mt
tLA7+jquYOl4maG8X+i6BBMMk8M+ZOhg6OI8SCofRfYoNnFBDs5hz0BnMdaz0SYj
uWE5OktYAhY1+AkYgoZtwJSL2HYQJXUqwOsFHaaf1GSxWjRo2XBvjSpIPIMAQJy/
f+4MKsP8Mwfez5qh0EW/KL47gF5t/EaudJh4cFoUX7wNpF+jTLIZVc14Lrqwg8mf
ugm5lZuqWm569r6SrgxnLER8jzfPFJnCyEh4mNDs3POMwjKa2hExfekT9KaEYJvr
nNsn3a2kEKeZ8BWEKTIklX6c1+4Hfqg/FLCASvwui2H/2JTken3yo7+Gjgz/EvwY
oD/nGDiujN3ykfx5KMwcCNs+97PiKVt9z3DgYjDp7yplBVw9badDbUfct8pe+5UP
ID5vZnn1BnikGVSUocetyrckZfhCMRcYpBl5pwTxZ0xfeYZ3OmS/HWYtnr1L3DbD
UnS6EYFlz7eOH9JOERvXohqHY6+XoZ6Z29jzVRIAx8qSUNyYQxo1/4ErKVO9Otgc
OkMDce/XVR1pm+M2jcvarmAQxqA30N9RAAyr3RXGlJY1SkTIUBJxSrzxItjE3FgX
ZZ/NcIpdbFgIa6o0Iqzw4cv/QvdRQC+q+ZsTZUPfF5Kfj9TKKXmxfSkG27/FVyk1
EW2mND5+Ugdp9Yn00rvyB9Opi6KfBSovz26X/Dvh57Lt4lb+gKDKVBwfd9i1mzma
bvB5TJcFIznCIprva5yWp3zWsbMaqqaUmms4xh7Y8ZaQ51LNhFdbiZCHb9g2B3cE
xJMza2yqK4v8d8muo2afoekN+0zGXyz6HcxbzBFQG1Gl/eFKm2THjRko0674Y/OB
27CpSwZ6O+HCxdHpAPwmuSNrWj3kRHwvpRyrE4DBYJUp1VZfyRHaoHnDbZOdp84z
o8e+8lOT8xxox4IBDeG6JIHkiioFUypgZlP1SVFvYRp4HIuZCkQlIx2gNt/TcfG7
EbgCYS/gxE0IGtFoNuSmLgc3GnU/AKdJUL9zSlWIMGgoYpQYRtIf+Id8F8/k7Q67
vuIUzeKZi9aR7IKbZ0219abkU5TRsUo3GO3EQevyLbh2Lvp5OGt3xFrL55ACXFeF
lZMCdHYYd+sLb+Ctn2Thm2xvHsj+FNLtMAgNQNPOGN5oJFvuCuhEi1Tlbk/g67kD
dAN5MOLtFLf0d5QZvfQCFnygPao943xSBt4cH9Ma9r2WMQKrZ4BgJDPhzJWDkIdZ
teFuG0xrmuIqayqnQ4od/tGzpwb7Zrh8a2DUtH3lttU+cAYkDzuMAzVk3JMfCHqa
8BDzvOz6WZb7bm7c2xVPLU+PynNrga6fYGzmtwNTs5wwkt/2G7WW7NqnD2lwKpoX
EgZ8yOWydaIrJPsamsK9pNTLXyH0XazUCI6whCM0nvMhr7SVHHiAZp8vRCjdRPem
DBi3uike24QMB/JbffK3KB6uhwPNg+nkRaw+wEiZkcA2KwpeoOehAWuqwCBZ9Uye
CqiiMll9YslzICeOr8ZhRiNK0FJp2dF5XgWQ+08wAwyCx9KSUI33SIZbElBaI5xD
IA9F+gs1qpIkZKBP23vP59adifg1HEChJ/s21DHG9DJ5geFf54O4crwndMx4fckq
iuew7Sl7wdWTxaGPA341/adK8r5xVCOGOVn6SqDq9mkAltRQzlDyA3qZ91AM+4uA
iN98VHPAu9zLxopFxzU5BCz18LUN6iIplqI8ijYQopKIb3pWjFcCyMfaowPEEUlP
q9SsDk20Qwobk0rnvKHPMBZPj3yDNGQU2EPUPOuqx2FLSmzd8GzNUd6tEEucJ38Y
zoMO/JqcQjY+PF9TF7UlxQKz+x9iQRUe3KtUsR0mzrvCGcERobnMvxIycyVsMZFK
nAIyqMTBIBJ7/MIPM1J4wI9941EQbwbOmRJ6xmpxspKPNoQRP7ByFwIW5lbMaHdM
I3c51J48wD5IeJ1Wmu8DryGN36fUPfuUJ3FcJbAqbtnltiXRZ3/y/1TrKDE2xhL3
3iCYr9rRhTZFnDwHDq9krJHwlXEKF6NDmM2Q9Gg8KE6R/O+lbaLPBgf6V0pyrcLW
kkZReZOlIXeQHJtsRaMKDbheYokruKLCvtY4Yw2KhXWQD75aY4FHQ9Gh4Q/3b//H
2jTh8SBwgTNo3tmrQmigo0UKE5+rAwX4+NRG0RQzBnjX6q0dYbMvynD32iFqac6+
DavnM/FVfnyYwVAS8bthHEUeBeV1/ipCAR90XtEuT849BW9FxrII52zB3Hc607Py
ABgMSnZ749aMvFxJMi5PTH2mTBA7SJrj/GZcCS4xS+cSPj7U/VPRgsbbkCdU1CVG
BqArDekQEo04veKssLfKyhyta/tleqozwYAWjMCxuh0yY1Hv/g5MZSyBz8+GQo1y
NpgCVz11tkhgvgL7/1Kdu1i7XccFh/KWWIdH4KBA/TTgdJ5tYR+u0MWK4PwhvAGt
R9CErEyDYJ7K/vBBEy0bnGgj2qZUT82e3bpr6pC9c65QFzT9liPiFsXsyITcX2nf
lwmgBhvorqM94yzWQtDD8Z4kiet1OsZXC17WJVYg7Rzu29G+HBrudDlco4iNkn+7
V9o1DAbH1uRjsAczhdjvfkAp2itc0ykwvF8ESos/C6+VyvGht6qiY7L8WNFyDB2P
T+87mt2XDiluUTJc1TkR/kWiKWW9mQraX2gRTlM6UTaBwr+5EFs+RzWAS3hI+N4W
2rbLAudsAKDbU7rKs6chBxyTZzTxWeMnMWQH48rJ+2nQo5zB2ucT62Bad1KPbLmo
Tsi1zUcQIJfJACgk40APyheoIOMfNh8Wj9w2LA+t3QniJxkzMqJ/GNfb4aAeOBR+
dRDnc+htfFjZWJQPhxYhOwSz+TZEaqzQVrP+lOCg4HCY0UUTsqgc/iQyMFdWBmx3
dx4kUThjScdhdJjG1K47apE1dhbSRt23mGv0lk2SwuMHfB4oth++zy6jDfEJSexF
lqFKNtnFfQvArHbFGj5LmBHM7unKEhJw3xCUnQAeBkzUkEOfmJylEXKiP+CZ8pu7
GAabStC9jOV/W9++C1f/RpX4upfjzrJdaupAGbD8Tc9sXSwfCMxr+SfXCJKcqveU
LVHWQydE9oUyuPEhdw9HxwJbojzKZk7eE17n2PIpCXCGA3gvS4PTFj/1NYETTEkL
q2KD5KIUQ7MJ3I2i0lfkQeXFYPfiFBjWuAXKqU1v4eTyhwZJSjfkqXr/mixi9n8g
JAZxkmiREsDbdzHLkMpu0OZFuBeBMmAoKswiHpZerZOC9Trkz6syn9pAg/T31NI5
86KOLOw8slGb8ChDCcLJ8sELuBWP/0ZC1caDAxcUh4tWdhu6ONKVrp/fSAuEeWh5
8b7a0PNB8AvU65S3Sy1RxDEsvGNgdg+8iKxKEXkn62fWFlo9y+rKFweeMn3upH5V
PZrgrICAuwt2zH5iGDXwcSNXTLD7RYVYRzGtvIuPsjVzhoRLJJscmI0yOLZwq+00
8q/hxyT3k2tixL3WglmI4efVQ0QV9O43PBOdNFseuWd/+NUgrGDJwz67QQvTiiD2
vCknnakUIKS1IkRLdZIRHvF9Vm4vGZ7NEZOYVbXmztawtcaZwA9W053Vbxi2liLS
0PrPiylDtvvQmpjGuhpjgnW0rRII6wMH6paroBbKMOSpt9jMt9fBZTWxfwLSkMEs
PexYecuGF1soBgl8yEOWvYWKjyOKLhVyjwoNkVrRilja5zRGphk5O1lcfhpV+ZIs
4pEdDm++GgaXUqvLhhmYyvLtvyiWqsLLNJqhYeQ35CWanHaPTag6l8LF+3FmxtBn
N6U0/iFURYb4pycBlF2KOwyN45cJsWq++iGXxbGjFuuWziT/DvKYkMo+1GfxZmpB
rNH+zkXyVhqu4gMfnQl0bBVqmTlt/YKdh4e6Qcqj0JZuuG1iJmBPuuQMRmwZ2cwT
YIqn3F+JcubdYL+JyhxBxKVlCgwbI+95CKcbYVC61qCxYwzJcl0dHGdHJpJyKOQo
KFUblkLKA/bd2XAFJsQCGQFalJxbdLTp6ERsaKuRYLV6Nc7hwasvfhrfj5VD5p9G
mXOR3uZzAc31+geePgdNn4PsQ3S00qlCAAs6jtzP5MG5MC80Up9LjuBgpWwGFT8w
GqHBXw8oqZy9FcRoi5sohGICm/BlOdTMEj92f4Qdb6ISFN2tRYgHoRHOdFNCEB52
zwHloRb2579fRQGA0FzvNG6XJQm1LQiRkm5/7vz6zO6epA5ZsQEaG9AcB9unKINU
BvWlyerNk2n0yD2jS5pfv7aMZNXP4Tb/8BkT35WuzKvUxn3sbJxyF+UWxkBEe2zk
XM+hm9mKrLFG7UPdo/E7VTCAajgseLyBL9Wy3a/fKGHCE3BlINwvKE1FpBNMCWZz
h89EXhJ5X7ES2UuXNQ95978Gmt9debY+2lsoWb2CspcqUoNSLv7YHiV+i68tjntx
QOloqj2KoYzr9FMfK2vTUDdUrR1FdXcavrtcpW8ALy/fnPD8h4nc7GDA5qV2+iT+
regKE7B3IlmH2nGj+qk72BuTxjUTH1j+Z3k4eedHYDU1OLVSe8L22G8/bVnDH9tg
iSvVtGs7Jz+MAr1mVbGslywu4FmTIcdJJeJzfXqRoLQR9M5prWbVI2iOncGjeB51
A9CV26FXHPdDemExBwt/VLf9tyiGZV3i4aSz3PCaN++OXV9Nd+wJAW11U/XAXhPL
9Q2BK/zCcpbaSSbFapBm4gbQkqvat1QQ8BeQYBqpMh0LX77VKTw8SEuTyc0tJmdi
OJbyWBRb1Teqj4aMTmrRQwbMy1nx/JVpre2k0yJfIs+A+AC+4+0qa7XAzCjs0+qC
0ECAUSPi9/0uUdJxjSkwW+0w/piFYdRGEmhFN/+TN/hZ6MgxmJCOtth6ysKOcl8B
wvl7ozfLP+UC7ShPy9D3pDM+QF48t4WBeYbH3JxU4riwCt31I+DmMXHy57bHV6bB
ZfeLuAfyZXw/rvyU8sjjj5+05i5adY1q+kch+6H+JZ6+5dqxhuGw9TQj9vkBkBdw
44sliJINR7SX4DIJ+aN+542hU4lkaK04hK5a/+fmbfe9jow+2vCW6iYB6l5TSjiy
/BqA1cyW0JBa6d6OXpI7y/FrSkD9zu/CnSdwVXwYuwvTmq7xmSPDt134ZHPrGq6N
dLtCbpyEtGN8J3KO352F+iugAkWGhzWG0+j/7Qm1+DKLBsJfZZdDpxfDcBAr8X1Q
GwdqjptR4Z0zN0AFaP+bMvAciZVYfTL1t78MSQ6TKdCsD85gZuejxW4SSCfzX2RC
BtqJrSjahmuKXuNZueZwzusta6LvjKn68k5rrQNm1ddFr5Xva4EzkhUS2xzW63DP
z79qL76ppJEoSMhcliP6A5OsxmS8wD3uHrEW+BQUp72Hy8jrftMq5jiiVKdhuosZ
Udh309CwryquUQbRj1aTxa3HH0O6jWWNdkE0rUxQNBX7wpSyjVTotDwPlyQg7Mom
ylKREplrtZ1g+3Ci5rYyEBMx55jCE8GdYWRhlHBgwHA0Ji71JlmR+8XFSP9eu9v6
8ildNyVi+RWVD2qv7imbz48SnVlWAXpwLObuY6windI8rIeNd49QGxHe9IrSX9K7
pCXvicN4rlgZL3p876JHCOoVz90IP+wRppIVIxpd0FQD1eKlmFySlyvrKQ0hcj8x
CKm8isX63/2tQVJ023rA3YrgQeh4irKSAQk+lYRe5+aTpAakficpq3iIitYmorMf
ETeXWIZrfwtt8gfM0jG2whL4RX1n+kFj3efYgQgzsYwexVuPoQom+gwQjdadp1Zk
8JvHTmQvpivMvdSxnFFPJ7ZeiLm3LSSgS5rFUW9oItiGUGjOvLCPsWmWIvum1k/x
VUIHfuWgQhgdjE+53rkQFGA9dXuvR7Aq1y740vAl8Na7t981YFm4nha/wovAZ8Wv
hCnL42htEefmaD472vUjta1CgSI1gvSaviwbIQ0gdhLvkENWhmXdFM1TWUSFNUjw
+E8gHF8kYjYRDkrfkWM+T2J0G6r6T1DWk0nDqPSLfsj11T8ZnwYpuGpUHc74G48L
7RD5ODR/xU7MoVGHpn1FJwJuAn0eZET+xp5PkXp33h/3jXkPIU8ovr/RYZFYz0Uy
y2HNvrxwLgfuC0I0yxuDuB2fIMxz446OZICcYv3OR24j7WtSw5UpBRU1jYQ3w1Z1
4CBu4jwFZ+XPY4+g9nyuHJqg5RrNqL3otRdA0ZMYxfDpvkOp5/dv6MBZQ/kmf+Pl
uwTe3M6GEVkDc0CzwFqCl0X1aDmDz2PUAyEdoV4H7uQ2pkT8wyK4Yu/MFrzvXbBf
OnwDjhWqahj8FVSYqeKRJcztlHCQ0IdvOdodmy6bcPL6WnGZRi/DmgNLaofgiusp
neVVlQcvUav9yL7XGgUYlOlgX/edM6RC8yvDqOuChnh8mA2Z2sBWHgNo/rUw31ra
A2U0vX6ysHCMlJQ4Z6uHRgrf6n7ywDqRRDyVzRNarp7zEYD07edzRM7wo62vjdCF
eZnaEv4CrE1YZZK4M8QA1tL8rN03DNPQF0foLSqqfeh5UNKbwvTb7zXWuAts++QQ
oh4696XvA+/NQ6QA6BMNmCp8exJd7bp8R1NrGb+HcRaOnY33Byjr4jb0CUADGiI8
ecSc6c7WPHlfRWhww3bS5ftsVR475lm/m5ztYgPic5RMza+JX8JlKxv5kcvD+VdK
UUrMPqAmSeKD87YXisI6aGJMOQWF56A0qJbXwtD/Kwxra9KdLooxvNhflMj2ZjTg
/6sIZMUC3zl3kbXmiGprAgLKFdQ9RLynFUteVyTVY9R1wMHJKyDz0AxVEOj9cllp
hJnuGCVb0+NpBMz3IY1wHdQEv1YLPdCyuHnj16VwiDVjTdp3XdDtk5DPuZr14MRW
MwCfnrwff3dJf8lQMnrKayyyj3ztI9uUNKBYMEMSTsNUJ0BqGdatSOxtNPomsbNU
S+v5Z9rqXEuor8Ndsgb2xaKuEa9I0nSFwxsJNUQ2wY6Flnvecyeuheicox6lAvV/
staZUOtTG+gz3pkYd8+U8lneRSUmImLwOLKZG54u6GUxAuB2rSW9qfa5PBbO6zSj
41e6AqLuwE/k5v4aIuVUdKSeU6ICqj1aNW3542JtgbUxP4z1BLst1JEAzrs96ll1
Q0q/GYYXWlJi5CMtY39XpOOQyvOIKcm6CbJ9SthNHG8WFFikNDCOXcp5gupLiGXp
e5fZW/nTBFygjKp6IXWAOdFa2P+xI+UqseKMGHM0tZHFX6PR7lNvmIO7BoZp4vzi
/mnwjiqMX8j40UR9BSBQUljQfwX1rYJkHtk94Zs1fISNVeIjxuiqlCzYFV32wXIf
nRhDfkFzXXqHeoSgBUxzPXPQvmnlDNG+C5rBxr7WtgSjDcq4Q7Fd+hE7EOQjMYau
cVJaZhc7Hs2ftIUsLq+c88NeOdDA5cd0DpKBzZRFOvQWfYIeBeiKIMYHr6OfCPe2
m37jafqETpZ13n9tMS6chf064OpG8x/DwT1RTNPV68PhzsqWndsEKdsG5xTq5tHL
WKT0Q8dVYZqzyNqfTUOYElK8RXtR0wu9V+CXOw4Zlqe5eazkzC9JMOcCmmxy1IkB
g6mfgFAmqxQ/WjvQ4rYyg4CHFE0dcX4Pbh2JvPccc8FHjAYj5TEG/oEb0XmaV1yX
yalVHmPBZ7R0+i4wkA4Z3feSoD3ISLaAv5yuiQxEA++49ctaS7pxLYEAX88Lb9al
DQzpi0nlPaF26uyNbImA8NoA1Y7rtStYw5HDGmzHpeIadkxGCFEWny8Kg6sPfYJl
R4B4mGPbcHVY/6jWrsUPY/cVKNU3Q57jVuSWqumH/lY394Dc2v4fitLGiZr/tSm2
NAPpzEupopdAX7zEQA/bMqFx4Bnd8ybIPq67IhAhvO8Mq6MbtxO7VIX/5HAQB5He
KsozCSbogVL0VjcJZJ8OGdN1dB2ucwFfaHcH5Y7IZDSMPdt7LGzfISmOV3b7mKx+
nmrD12XSUjIppfYioa/oEw0hXDJ8ttzRostgx6PtuLV5DuE3S5TPu/iURmqJ0MBE
xbjAShjLGEPhvdErpS60SjCk8+LSWcGqjtY1zqus6ekYph1exFAauJmI0ZvaMOFV
ZiafxpmgadPDn9Q/2tj92Nu88TSVkMzprcI2Oi7taApRrcz9lDroUHnYapXb4cK9
/+f0orIsky+M1X77d5c4uVDPYraAkdJprpfK/I0AoaDIuFbOqDHuWf5gnY/tgRqP
ZENya6ddjkYz5h929cpVgr8Kr6a4ma//VDsiCqsgaSm8QXVeweX0r3mD/is+1/dD
cfInNYKf/SZg/qYnpp+ykcpHuzypZ372z9jgfrXyT4Z6mulveCbXzlMz8hBLPTSB
i/fY9bo/b/T3I9r7ATqA/BHxKUYgWwR3eXmuI4ihXJU3eRnxmDwmSmwrH/y5a8ss
T8sSTtUa6jb3VPRJupLnSOXfEngPerk4jaXS01tZA6zb3OUMpLHjjzDzpEpEZAf7
YvJvcl+QeFng8SKeUp6ELEJBsnQafhexk5Fj+6jb30qC5tZWfNGTuYDId+D9YiHB
eBcxrplxMqqzZpcgY07Gc/f0RIzyBx66DZenOkDZuY9uQAgvbhclCryP+IONR9iw
rDpu/jt7CNA6sgaPC2VRw7cxo52KtYjlgopf2Or+X35Lld19Ku6UoFKc3W4njCMN
ATDWc35k3bQsQtLKV+XzicWAZbMkRSVPbZ/QzzgQ4CKEg+oEH2fPfeHJB0k2SvSX
RaH/9HDV0f8ZUaaidWNWt34XAZ4eAUPjI4n1y0FmhIe1dfltQgfmhYtIp9WcIn16
DiZ7UCmellzLoJujlAWFOyNnMnBfh3kvjSchCAiZSip9zdNFbJO1W1MNgtutkaKr
HjARSvUyMEWZDkuQnUg+rykBN+cHecJIx+O/d9x3Xb/TMHBLREJQiwCVg6jWzh7h
v7ul3tf9dAybJ6Of9/GPh4C+ve26t6mu1j28PhHIqM8hv+ttVSSUxWp9ZDkhb+MB
0Ow+BZpLF3cF51qhm8AmkhJTrAY4heMVdpwIwOUtZRtH8k/1sj2iBPDJChadKTfF
zTlGkJbEz054jZfBC2Lvcnls/DUNsQ5yay8v15dXCNJK+syLeaLPSvAq/4EANSC8
TAFmsHgGRw7E9O/f9O3WH+fTLJzpfDknS9+ypHOHb2Au/5RYV1XnTNOt3gmX8rfo
pRjDe4Za+I28AFsk6PwKYUrykIes1y4OjzsGA+g1OtH5OuHnYHmRPyLyOVgwhn7r
QIixd8JWCT0VJxSQVT8RL3MwJl/QwqOKP+VLRrgPrPAv1N413vNxoGN2jvwl9887
D8WwZUaJoGHgOYT1I9KZzoRHY8ZjZRH4K5V6mjLSocEPFUsBa6/oa0ZpnRgsaywS
hwA+mX3jO0/vSdYr9lGC3LONzbJrggd9Llblhku8auXrvNOIXJHQAH2ZcfDaKIxd
IS63aGXzg14Hrm8f6P1VtZiLBugv5N6Dgs/Zvu930B1qyNjSR8yxI2z2Ie9MBtVa
XOEj9pCboM8j5XweoM7BktNtG+GAGLQ8sDwFRX/TqeuVfCUaxz0iu2+kpaIP+dIx
xuPiL5zoK4HTaH9fMjsHqeQnF83xQB/8HeYZ9fIMt6McxYgWRwcfMusIZworGA37
V/mBZZk1gTifOvkyZtbpgwMMhC58J5YjiAXECNCy+DLqEOmKbwub0Ei3Nw08im1Z
9lK/jvUOF1LgA/4zfrDSV8IxB7UQJp24F36b1fHRfp9zOnL7v7mfHazzksz9I8af
lwI2f1FMONeJc7vFaWnHsLBefugpDimsA8Wtg0EdLtX2vWCG3vWRTeAOThLjdCqY
mwxziW/AeQs+X0dZYuFlXOpLtu4Qg0GSezL86G8/j5sedtFIpeOz5dpI1P5AMRV0
sYP4RY9XPfLWhx8oxWDgsad5poSOOV9GryUkpXggyjtV27qDq+NeWBSuG0KM/CU5
uSpczWPkvMSIffym2sctDtdyaVXhOsKyhLEaftRvJpaUZq5xiYO1uGBoKJsktXfh
/z6f1UIFrmEZFsEsCalxn4q1vWb6Z0JdQx6IAX5w8JL4LQbGMQRNovocYeHudDTS
VMEG3f4ApWwAAKfGDS2/l3OQuaN1SemlSBYf9jGEkb3NHLbC7WXlcE955VqkG0mw
LDXft0q+ZyczuP8Amn7eAWFgFhGkIrSg7Gs+V5NNri4zgSvt5VuBEjyt/u2hpmFI
bsJ80cYM6fF4SF3Oo/b35/rriSJFe4zEcQHBDbJ4q3T48varF2tkE2Xgu3ZAhM23
UVg/nUvH2jScyojCpzHmC4BTKgeYodpVhaLdlipmxlYt/CMw+45CjW6wAhWnd0Pe
JjkqkGpcXO2kjO4Ykw0/FCZsViLQyr61rKEYexhxV8QmfY8d8YzgP9LsQe7Sw+Vr
xpABZDZKpN23Vuev1i13OwA0nTgfLtaiaWi+kHAeupquGm2r9UgYqDuQMTbHEI7x
mslPlMa7rKBge6AQoMa5swGL8ApLOFbIAhSimOr0W+T2Fx5rnzgnedZrj81Iepks
p+7KRcG2Qv6eX/83FHCGS69sNX91BpLcsKEKTbNtAtlaTDMDDIyowo6+GnkZTK51
N2ilAYiXGDCw+dSSlx7uyjnqAoH7+qn4iTqgvmYLxeG/yXiDVp90hPcTl9enRVdC
2voRLaBXFpKVsTlW4bUMUbjM5onl2GXUnCUN25ZZZTpwc9t0rcd/3f0YAplT8tQ2
4wtmIgYLna+GIYNv6imY9um6TKuyNJPX6KaDINhB8tA/9CC/2Mp309EAtEj3bZOp
WbuwY3iAOuFG3iwd3NEyS/qk6uZYTTzMS+Z57RrIDgrPJrPk44L8lLuLKZKbjeKD
Od9vl9FpS4GaVO8aXVfsAXrmhAIE2XpH7FZzotC0RvnC+y+MsdVjP5wgDsLUODVC
QLrqTJDAOfgtpr2M+mqm7eSq3BJBf1E96scYBC8M8rptxwFQQjVVwgmSo4ljNdS3
R9J/rAdR+rQdVeongIOL6Xs3T7FBYz082v2C+SUtUFXn3wW00w/05N/4sVnOE8lS
M4TGJxqHEL4ViiolEHJV2sJS9HxfoVP0QEPaRNJrnpJdR1Y7TAuPgV4H//rNyir1
fFm3EBOmpFuEvDXPoToxh8FVue8G637MT5BF4K0OpO9aEfrM4QzKq/l/81ye+MoI
o43wdAIh/NR1/AVhS2SPGA4H+FiLeDWVXu6U2R+zX5RhAO9m96F97pdtgY5Wol6p
Y0sP5uT9pMLib4o1biqw90VLoq/082nJ7KZk28VZwN27LMl8q5Ysc8bEkvcnyDvl
My5cSn2JlyrtH2Yt7ST+2u1fdu3lMsewyemb5KREZ0ke9I445UdaUJd8Yii2je0z
604U6bJQJP/oK466klF1oaALE4gy+ImsfSW7G4prtyal8ZXttpQTrvVr2mmz26wV
lTvxD8RoeZzkzwrKGG28dBGyDt6GzcrqowXoy0g7Yhn7kO5etekTIforehCV5gYm
aWs51f5KTtp9en3zV8ph3WNxlPeLn3efTJjU5YdrR/4mxVaEUN/NrTmnz/cgbYab
iNFsJ8nnfl5HtsKb3ysV0PLuK0u2p2Ai2A2/AdIBQzeZj2bIc/4eNXCOkmpPymFf
LRRvb6e9P638BnGyf7aQgWqAuhHxcYi3wuOxyrKCUw2NntEQ+TVcw5FvyyRJ0AsA
wD4VaxvvM0ei5jbG5ibHzWDLiJkyUTkIEbHBtUrMOlosIJqzs3M24vCYjXiYyIE9
CwS9vpobOr//4uXjDsbA4LuCMCPz8sbjvFzroySYWKcY9rCDzPyXYQXpqtDGjtdk
XDDHFoAtfm3qZQ9vCzsR44LbfhpHmhJJW9pwxJqoGIly9Wv9ytUmVg0N6CS45U21
HJUlGuTqfQJdda3wldXmFydyUUD+9YxMxD88KZDo21j3bbVA76C852eAERksBQlX
2jDXAuBvKEVFCwVBBKXdKLtnZSfJkBgAt5+rhAHSsHpn7bm2LX2ByJzj5NWPLnY2
s4ljdWu839+BhReI9WvPJq3iy3QFpZKmNXHB/sZCpuFOj07hRmtz9Wk+wwOj0VT0
nz06zADso+lA9Yzml13eMTl+1bMVz2T/Klj9gPnjMB3KLvKa7SNek4gqZ4dCZfzG
kqhx9keaCvdqAmKkOp06dlxh4DUCC6/uTa2DK2c9T5tYZ2DsUdlC6mq2A5fkWXIB
sRq8s01q2GwPkVALEHyC8tIjxAMXaMHTzbURvbk3R6AnKBnnvNx5C1b9QG/oKe0j
lWK7Bk8DfCXMbbLvz1FnYa9dMNvNJ16D03IbZVNgyzKtxV+4igP5CRx3YS05ux9g
+XZcNTizxgQE/cKhn18y08wuNyO0O1gi/ixiZ7nVvjDGphpo4QeEYG+Qe+GYC8vw
LJiD+UhxapjylCyxkDa6vCqWo+D9084NnnbUbiA1/AwJIbsSgGKRyJJ0fityxUDK
8/M+ZHAsCArkh9YaxtSx4mlwDhqfdF1fjf+ZOc5a615xF02H8terpu74UDWqAm8W
COFlsWF6OxRfi42RPpKe0G4++CmvoJCpmPZhhu52E3wVlBXQfvzvMpqbjqVPkYHo
VgdQ+nP0293AFu1YgxuDw0fmy0raBLgYgBgMF7ahS4W5zdjNdQbAAKEyqGMNAbiJ
tTvdO8zm62bTyveuUbxQG1ZRKcqgfPpSzVzqs2ZRgBoY8YKD0zMDIfKKjN7HZaT0
lcLBazBKjm/UKudXKMhjZOwDfW4NNzlnDmaTgutxdfzf/isCxdmA3zxC+5VIDG9d
FU6mDctT/QO16ZxTByge+wJlouupmCjSFiKRb8RGvY/2/Z3ml9Ujj1lwsWczxjRG
CSrI9jLn1hH540li/8HSC11MXUOCldRsoPf6VvIrXDVyCuOjZ4Yyb2oxJw5QOXEP
ERg5mNSwuo2lElewl2QPdZVCU7zt1XTJKfdnVZWTc9TiIEPeZokVDbbQPLq4PtYy
DAtLizlPrS5/m6eID5SUZqpSqTjkMKoLveB36YK87Xg9nf4Sc+Gq70TwEsURG1Aa
zj7C27Yxc+F47OSIZ+Gq8sF7v15OdyKc7BGRPTarhNX8FbKxjL7yJ1qWPeV8ziKr
WrAFIIvSw/am0/ZxPvrVEz2ZRvdRgibvTXwBceI7rlMciaFzzb9DJ4Le9l8x1DCA
3uhk2sP25MyLSBO4u7o+YPdXkTsvcFFcWIRR9z+GSRZ1zpxYpT3H0yIPmSRzA0bp
Bi5nXgL+s7lNJx5rLQmjhZT+5TwlnwcbuXmUpDSCRxpctG+V8kCOSzbmIU8Po6H6
5Saj3L4EJUDZ0ZVHnbPtGQePsdUpS/R7Z+CQdug7AzKtvFdqtuhFgg1H5uYuHdtj
XYU6GpVqnRh8nNY3q1qhsdPy8bJAODQmIpaGASDtAeAZtDNGM50zWO31P4JLQ/C+
w6/1eflSQBoIlnc/6Oq7HZnkKSXhsQVZWFiqVHBw6LDDBxY3n5p8Wc+yxQ26H6zV
Jw7V0LW37pqvU03ha4vURXQLhl5f8473sUQjomKR9DVD5VMFSmWQ2svEIL0BUFJB
5VG6eCyEjs7pnqotrSYqXkgWRtHwwBc/AyzxWWMJzYsp0c4T6s0Dxran2HtZ6pBk
Id4qZ0ufPaEHhCPbvNg/fs/62wUrxs6Qvk9oV1Vscb/YW1Vb2nfNU908Dhf1c8wm
3vibVdOBO3wP10giTOVdjMcbAFN5GUyZoP0dtmmSSCDg5+cFRYZHDnQRpfcKBUIv
o4cSsyOKhNn1tnAfRp6Gid3wGAIOSfCHnrK1NwL4ZueurVK3feHi49GEOUh2Irjv
QpIItbF8kj6XZNEI1V3lGXCRg5P9iU30/qw7XHMbBOeNEUrcSz1HxlXwXnNH7/3Z
+97d/0h/NsmJcjj0cMLpYMyMSJ/8Pqsp8RnSKRUOUg1bv6Xv181pGB8EwEdEsXlB
I2IFIacx1o+vaVXkVXo4MI0Xj7uHZ0/Bt3z3PO17udReI5xifQ035uWgvhTawqcQ
OCqgVPQjFbrfVyppbpqyQOlRS6cR8Uat8k3T7epbOcgBp1cQIKZXyjtcvTfny5b7
kpBxBqJrmL/qG4Xz89dSPHimVBzMWkZHh0iuriKPJd4u9O9liN61MCCZ74ctPmyq
SyxJ2+Sj3fbH/+xChMgm985F1447Q/kqS8VxY2WZMYSuMQjrJSIP5qZ6GpV2rLaI
MKn2tAPEp0uHRG3xYI5JjbFkVolyfl8OjrcsU8dPEuGyzFk/6c4rt27nLLJ71TDj
HYjQQwk4avUy0FilRuiWIcCg9DCsTTmF2bb0eAWgS7R6X+0OmlTI+ejUtdb5MmIb
XZWd4osXunCCYP7rX7wdyeg3d/Yhk0kfq4vWYiVzZ0aVVRZTILTTPWb1HNxox6Mv
lcc33WaCt6VnORxodKCPBOk5fXmSXd6d4lJv5Q314o7J4u9R0y0S2hxAs8Ai5sXL
gwilHzspXsgdYG9Ed+1BwZN7kOLppf7XPEHR7qG41jASE7CW6Hy8hVdWpf0nBNbb
I6Kkj7Q9q9VY/fHrwJ+48WmFrMiik1zkARXZvgNU9iJzSkWTwQZ64Kc+Lg3VdM+Q
3+rdkPemJ3PX3EDdIJqaS1k3yMk0rqpvlMLbfYAU4Udnfyg98fqA+/hXoBkw+7Nf
S8ii3aAcVS/8aYT8dbi34F9aR+5ziKy3CWQWqqm7F+vp+Ch5uNZjFDRla6a8xpsZ
A6eU0iTPeT6vPRL1Lm5BU0Nqo+9SP5JlnXpphccdxznNcsULWmfYlSB+RvgXCv5d
LvhChVbYJ8FiJnkc0DuRrA0BPOh8rZbylTPmqt+e1EQTNIK7o6QUsJ8qGSLfl+mo
tVyTlFPZZrrRqJTVkVmAwaEt+5uX7mqkJC9RX0SBiUTWNk/jMK5W9NByWE1PzyOs
QmtlsusGgbGdu5aYvI9ZXAILwg7DRyzeqmzZSzJ/btLZ64JaU1vGgd/mRry87Kc9
6Lc5MdfmHNWJWGhQXT1bMlfynowPdfSWX9QylL8Y1z2cqwzrE81nqUx6Xr+mckGk
D+RTWNai4S81o/cxA4rDVzrnP4lAttj4gGoaqu/4p+AFLPjyiLO4fuYKG7eeVm6N
u5l0OS+7i6JvMM5lucL16++qdIEV82XWtU96lFZ1PVaes1PRsRkPO98S3jzqHxKu
+lARtd98eGCncqXkwMdWLE5eMiPn88waol62dsrjSNAXmkEJgmv48CwZTalngGGZ
0k7mtf5n0bi6kfGOlFGZ1dRPVWhZUeMPBh/BIpya1vlsa7eNH6smofINbEhyF4yP
UzIUSope4DQkF4a8CXHdeSWrxKnfSxXnPykORCyaDK2eqByvO784qfK3VF93oFw3
tpcuTlesQWY67EffpArA5rvpCSNMWWy7S406EY6zKWh2zQraSWkYjpC9ngSB4QgA
6J40iLjXrwPNSlwczSAIaVANCGkrKWLCV8Nb+BwElZhp9SoVtxYy1HYmEv5m1WDx
NgEKVvm3Z6a2CGQ1b+fL0NC25xqmjnTxGkPCT8RYTGGnCO/ZeTCv6yftpbF4QvXC
bmKeXbLnenCfKkiiBGfCBxOhOpXxjxIcgBxXZgZitGMhM3h5P7zc0sXBsVPEW/0r
lNqazVj9H3kckLVfElQppHtHBquXx2TY8vApkYf2exE4I957iFAkSGqljS21FqsG
gH1GsiGOnWtkQWcHl1M0JybLmcYDQk0gKMCPjvHHaKjITozEt692yemgktKWw38y
D/jo5PG6X/tcJqPKKp026titwXHlM/4XZfCHeqr93SMF6+iQ5URXsPXOVU1ApeUd
qmhpQ5tXoX59WlCAZqxGDilV+uwSix+cuupTzfoSg/YGumarQcR59sx2DfixZDbz
PSYzu4cnUaG8nYCYIK5czjMo3hDYBoZug1uqw37HKtsJi0jh2D3I6L0vEHLONzDk
vMG2Dfy6ns5/v2DMxyNtl8HDRTtk02ABRIAbVAAVQzJYRZcfiHx83JVvj6BxZTzg
8Rq2/zQe0rDNgoezp/4YelLw2fpCWpwWIkZ1cBJklv7T2mTuNAwz5O1z3FWscB7M
CSrmnpJxcG09tHrrwIz86xCJw57No+ovsHQA5Nii1re9A54q4mdMYxbRH5zOwWgH
maMjti91jgICJsuezOCeXbXO0yfgin5M8fnkkiJDqdcRT/OY6udi8MKtrwPxT5CY
5fq/Di4wMwK7R2RQiHlWL8gn/+HhJ/G3PmLvtHkvtssc5oSa831rmKnFWbHvEl6a
Md7MmWQJkyCQkbE3EyeY3Dme8E5muS7De7sCfXnGujv45XiAjMTTzRyN3bADOdn9
9tESov5za6aYvbOJewcDx/072Ey7el7KF8lNgSs7fPVMwXQwEXQn+HAL0nXYDwGg
fbUsYlPpfc7VNVLj1Djh1SaJcpy5mkaeOcb7TJhQu0/ZxvPmv/9fJllKTQqakJcd
fujcvRYsebNBQ7cQr9RKZOFShsANZnhaKIYkPY7SzjAKQD9HhIlW2c3ytPY3OLjJ
wX3M6LsbljfJNRGSBoqwmS7SgTeok825uxT8o3s0fDrL0sa4TNCozPCPZ+i8g8cu
cTZwevv8jMn2sZmImEYU/3/b/FRrnjmpUKQPdP2ff9NM/BWHv+0LuVmrCfQvHSL0
cnlSh+dA/y3bvpnaFvkRcPHLFixS1mRTdcYEycAj0/OZF7GI1ZW802IR2ZO7coQS
XGCp74puKXIIc0UiqON2tHG8kAzLvTZ8bl4qqYB2dR06UvXT23TDFLPpI4RK+qF2
eR1zAO/ZwZpKYfe73CQxGMTHn0Nt/9ex02+bZw/u9WFdY7hh8zqksU3p8buIoNjc
b9z+5q4REUJB5fHOmhFd6TPeApq1XmIv2yDmCsgKgwzMEBkC4V/rbC26+SE8G+TY
9TN2YnTg6bA/OT+Ak5ZIh9sSCXdFxw9EZ9P1+XSum0EiEtM65piYnMeFRVEb2YvF
Tk3oD3R/uedhIZAscal7817fx2LTJSA5fAKx3AoaS+pWvTIm4/0NNunDoJhudE1B
4R4HAfp1K0hnb/Que25aK1zy0aoWyE1tw+C8oimJ9KNmiuLqpuy3BWQ2aIDGUkWr
mLU5oLV1IY0TB5OXwCk6svDE8jCqhfCzqKQfM7mXgdpYASIKLgpHo3uxlrxMZz4D
9DX2rzvfw6F1FzhMWHKcThuoaumHeuDXRV+Dinv6yW7c2YFWv/srMPVbEak2dzyU
Q3B+R/zgdmd7ANafnDlL1PFflEoNiutoFGvU5WRGTvbiyWPw9YM04ARpIKEGgV9/
giiFbKaG4HHGjS1LdvQvkJ+wgYMBgk3a0rQ04HPfcj9ft5x4JR3pumDIXGsWqry2
5t0dmmfinH5bJ9TJYstlXTmfXLeTMEtN1OCTEwiYxtyrcPkzV64LbeyPeMX37wTd
FB+VP4uDFkP5cpnRyV3cOOjLtnxC823KAey60r9VP9dxTkT0PU168YbIFk7TFNjg
VrktZ49patM3WcM1aUcsMR8hgI4pj9yDPQCsbih0XwUFfw3JwZWT4S4d3MMHZwLZ
cxSTezERCGkvsGqGwAmPPxota2JY61dRhRKBhwTwUvCWtKGa+DgZTEsDswR7gi3L
MyRCPSj+51bZSxTLd8AjkCPRA0W1zSy2tiJsl7YvPlzS8zdx89AIjHlm6p8dGW0f
kKCnAGmeLLPdZfZ+smIZX3sXQ/E1mXEajZXLt0zZfxqY+sE9vL8QT8PrXxqv5qxS
8KbCeMdIkfeWW6vOxGY167onmLEl75F7ndM3MafsByML2QJ0Ed2o1p7R99VeetQ6
bJPdLg9VOZEv/qykIZpssNr8vX1IgOanchChVrEcmqpLu5rZIzSbY0/37CMsNugi
Jp6N5RPWat5jWDrkNkNaX6QkOcJ/lpjcHLIQzukvGPqE1akiMjio4HWb0I/b2c7F
xrp9N0xnQyZlvAuCaqmUdfbKSjALkA9P9QoVR7f9C44SEc6Mjw0LBqH56l2M55+f
+rcNxdv9p+NQfUtaBO7/qISi09Fdwq8DdkzYXlXFBTsNu7ZPLNxaLB38wWNQwrNo
KCykluuPXo4NeSBDmdNBcAaMJIdOfgHnXgN8pWwH8GhIuKsdRSktzIJNcdSCU9T4
A9Ty0cw/DAR9gRlw9uzidzsvREKV8fIa3zMkDbAvYwuvjsQpju5fK6ehi3wPn7CX
GS64mzXEe4nhaubz2Z6Jsgx1RDP6BDZ19Ybh4Pk1mjKLuVUAmvJ1NS7ZH+ipNXEO
qQ0G0Of2M1ZCD0YlvHtfXvNWa6K5xdMThWcmOVi723WgZZexgBcXDM6nqeyvuRXs
cJ4TJYof8OD6x8qS4EXh1xcQMt6zvgP3Ub62BnnLKmptsQALcQsvErazY2byMhoC
VQ15WNDkHGrfDvXmfVXhJ4zxo9n+2nqYQunuJ3ocAwsmYS37Z3MwW7dFZ1McW1XI
WAmkoc3JyTGq7gvSP4/NDApaJqE6EmjiDr/RBJK2Q/GdotTGm2OHg5bplnaPlQ4X
GVq22MEcwKspQD8JzXBw2dMHs2z9tuq1wvxYm2hI4lPjHhVBJnzl3pGtTq1CyTSJ
0RFGb85Sn+44l+L6wqsqc04QTKws8hGosXnT/O9nr56ZokdZ7inAbO0d7vE5+1zj
xBrDQWJpVVGuNmBt/pkydkD6IRRei8WwysRpTbF0sTaZ8IC2kdA33FO4GQQGPjq6
sJSioxjnVOsj7sZhaqQ/+i/bFyIK6OTUXF0+5VR+HAO+L15Ew7kpWyfGwUii7Gss
CYaKVcXRPlZHAp4TgVvEvMQJCGaSRN14Y4JQFGCeyI9WvztuO3IhSSKSqG9d8+mG
nWeFcAU3ODYoSH+e5jEucHoSLapR+W/FpspgbroZgDNHW+/ZsnXWMLtfFCmiwNBE
tmN/J1CcqDAQtNL9FUb0VetNUrBQgerw/Ly+CjxwEPCk6FEjFYYEz7cF88bEceYx
/TizkocRBawSOav5OOAkeXSxysV6TMjJPX9xr02AhP9UGJW6myVeG0Ovz17g+ML6
SB8zXqyVjxmspDzAweENKA4xg/yeO/uQZAK/8PxQH/56aEKIboASnLSHa/iO+GkV
384vX1HpBdXOl/F9be374A7v7292ygoFzcWZ5JyL08+QpzDWV9gEFvZGPvmCEsky
X0DlOFfN1aKRPEMgd+4a+VTedyP4zvk4XwEhbMDt1dgUmVBR4/ET7mby3ziIFhOv
6kJBxhtEXuiQvSUfl/47qGhJjG6Fhxl1k6FDFGziaNm4XFAAf3oz0H3yNi8XBFh7
psLeMl2/4fLfIR/gnXHtGNwn1EO4sas0JnoIy5XY65LCHMHHAS92wnz1OtO95cLZ
6OkfOhdZYMbOju5jz5yNHF+3tGWLHUIXJziJp7L6fdc6MCWbJKzfqYsnhtK9hDF8
LnHiOQzY61qOt93yl2z0l6JsLN2OEdNuol2ola8EaxYUqLDW2v/5+fKIJAxz94wo
JOmp27r9Upwld3WsDpDHyvfBJYfMvnVbtgwWqt9A38XdJarFo3i+uJ/lyfBiHZkQ
iNSW3m7mGjqFztqfCDriSsUhnjPCxR+t8X32lZs2gogsI1xm2VZkiuvwj6EC36WX
EEGAxxmdqeyJKVomdAIMb0Tpu9YfNIqP70yDQQKl4tqpQLGSMRe6gep07QYUOz/K
wr97UAXYKi78r9bfASzHUjaUvylT2AgV3kodQIxlmh1xu+P04w+QcyXAe6gJzhoL
cudiRNV1vljrbsYgEC0SQ6zWfe5IvaDEpkEC/NNmM88VvJhdgdOmj0C0Rle6lseA
AvV2LmCF9Lv5Yke9fC2XrbA/b0dPnHCAdO9fMOo/FTpQ/aCo/W3uV3EIY8HJDoVj
yPIbRzdcfTQiUNKirXanExKCOAoquXeakgt43lV3dJXgU7+ZWNTDbpPNMSXXpoZQ
fWQS86d0LjPzjT6kbh5iiQsJCizGBFkuUa9+3uan5vdWN9YmTXH9JGuPgVab3pQv
LUC0NmV0BEA2J9E/xD1/P6NsUhZ/23Y7TVhEWk6ko1HVQ3Rrjdp33uvO+k646Lus
pDyygKVdtdPC6m/JUZEXELN6ogJqXCHgyz8J4xhbASCQjbSiRW4pJko3tzAUZimO
MrpMpM5UGc20EBn7rFW5iN6S2Ds3QHdvGgvowIMkE/SOkgZ7Cf1O5FBdiYtvJOw+
osWI5UuB0hdGoC+PIyzRwIzkCXXm+R8zR4f8ci5lb7OzZL24nHlQjBeiMnRB1xdx
oxi+lsB7EmSvc8802P1ZKzI5cgSFyntRszLLymBDAqvFK3/XllWmjMsC6DYMGq0j
OjvLyB4I9+iM888n2Vl6Aeu1W1tdim5Ub2CKRI4d1wTgfSGOVcjFvV06HBSmh1DN
WDVRjy3fJPnsXfqL0d7iRvIh0PsLMi/Nn3/CPTKNqjJy6A1xxhfRNHkZ+j1O0qj8
igyWe/7N4jFPL8EYxrNPO2gewXtuUBDAjMDtsnGTVYpP1/jryoRUCLAhsYR/HlRO
tar9OKQL9yyFzeWwLpf+Qve4aUWlUaeoP6ZfdDYIsQWm/iJIWdA6JQ8sA8B7yGDm
0e7LGH9pOm/MSHWgAevxrQu2u/jQnABNHqtShP7nm75nPl9zB+5DDSzt0XCttSLq
IMCgRizTjXkTaCxcKWWgRFmzfxyTh2PdW9LlEVh30SXGXUPErxWF7nkntdg41RjD
GjD5cGkjyNE62L0L7FRKwSm/gto/ANIgM4s9fx+WOnhqZhIA1uTsnzPXygPzC5Xs
M/HgiyYNjybkWor+43Iun+HwJ312beAy4Fp/xfVo7Rgpte9Dvo+TZ9gnQbaRp+k1
L5x9Ug7EB9qDc0/2TL5UiyhwtRtFvWhFUeFHiKlg1JdR7Jw0HiU4ZIGXh/53mop1
7mr3qckoXIFvvswcIelCRcIPaulbcrQ61hbeSR9fXeCvIvqcTPnOEnGliqsS5+rh
3hJ8DM86ShgyIWWGTpHefmPYZdCvIMAnmNUYtujcL1WZSIjXtEoHh90QksLKocgw
6qGMBRvk37nLWCHswNhn+dxRenM9jdtBg71Zl4iXSQkhjiLSRlhl6/XjW4Q3NHkR
eQPcqoAHFB13FveBdI9xSV2g66oEdQJnHVnJBDMPFims9h1zwFEA67qeXYN7B9Vh
T6L3JDXfyDqH+3D0Gsjpue0ReKpSQxk/JgreDDfjmA7WuAzzlZrjL+AhaHrCBHJc
7v5Jp8tGgZdCiFFDbg+h/XxQJh7HZ8Jqwqw/G8XfeJ5V90/Xv1VUZg35I5tJDoI1
4s4+WV2to204+55WjetLKILmaoyls79Nld1nppBoWkqBh55X0AiHyE+8e9jld3UN
ayzSyu0OwEk1mHD5fOq7MUjDGJZ2G68GJbYCN13GbvALpgYyZxVmAs/1z+9g819i
HG9vVjUaq89EobYvcjo3/Ww0lH4kuFARdEQgkcFO9XUljg1OOFG+UInm4viQDoay
C2nCJ+Y8WS+o2Kn2E+7lKrhtJtClBDOuTGUwV6DYDdjQk2/GuKK2vq+RmUD75O3V
UDlCqFKdatFLlbv/DbhLNQ9yEFSaOUakh0bfdhsGSReHxT19c0vLEgWZk6MUFcJ8
iIk4OyQFa4qwDhfA/tz+el78isWUu1qnwNUFhcorjBrtfUd6fwkrno37WkKB23b4
xMZJSBwbKO3t1xLx8yx9rtb796L2VlkY7XExi2avVnC4ubFWQuw/crMBozigxG/e
JDB/aIeEgJQUlJKPFTVcVL7ITetsifbIaXvIo31Ka2FenX//jbotwEPvogljBuzH
1hPtezrYNGvXt0gagIN5hraqi95jFJWwafq5yGSsiYhikiPO8xLFAvmKgQ3j/Tpo
OVxHSJYRcHlN2mFNtBGu/dQYpn1rBFjcBM7+voaiSB8S7+u2mRzla8MypgQwGTdj
2Z5vxtw+vf185i9xps/2VK3FixmHJyEgsBe7vP94YNdWrNdoBYw7Hx7BCghg09sY
tGWYOa53RK0vyLuiqWZhfOWvXfBCIUyJ+mi8pVwM355bkj8bAqx/piOWwTxyP54V
KupmILAS5ZHFsa0Pgz0J0A4p8gCNtYyq8GkYoNAtLcpX9RF2rHH67IcYIkB6LCIo
lKpzJXPf4qfpJyY9tjNfgCYv+bG39jxBBluYa7vDH3loERd9GGm9R0xkCx8RQ9E9
xhgiWiSstybqXhkFbbcmcyzPYM+RZ9rTEfgJZZQG5+Kg7dmht4P5zWGd5LN4bJrl
TaOVzVm1wTec0oDO4NP8JyBpAIBx14fU5ZvW0mnVBZ7Ev8TtwcRu7k7TmuzbkXGx
bOqpl8czamAeQy6ld2ol0hDPhDnTiWAeauAg5bIa5gmCYDgMPfMs42fqm73KD3R2
3Ll69IUPh3dKWbLH+8cGZgk3GbFvb/mmWx5Ls+Oz98/JYNMGe1HF1lI8+3e6RCAE
viMjCfaPmPn9rmep4P5th8bfjbKRV/tRir6Q2lyF9feMXD+muTsMG6eE2olCNp7y
3nILxMXSr0e7lSeskYYWIDe0bwuqKZY9SfTAd9fjFZtXHiohV4BdwmP8FVZu5+bc
s08S4e9Kg3mf0do/UpMIMEqSu2QYKyzcmEl+w9l2CyPFC1A+g3Dw4+NyIgm50hJB
QZszbrLNtbC/QyJjm+vYVFLfCCjxEbifOHRvEgvryjr39H+F8U2z/9+wipGujuCX
dsfoxyhwf1y8mdk2Hl8N8DVXTjySNeRwFB060oN9GNkbfshZb6FYb4LXFePkhlMc
1zVD9KXgd6KlRJkf5eL8cehKKmnZoJNX43FoDh88Y+2IFeGoFkZ2dvUFnApO5SBW
oy7KKxNML1F56MWB6D3ApFpe7C1ppWSMKBQ96lWxGkcmNfTvPabWOZZfNrArGfLy
Jx6ixrCUatNH5UVvvR9xyclVM1ZgePdMUYhJqpOk1/WyDOuYKcCW9r4BdbJLU3AJ
t4VnNb6YPWvGco3DgAfTP9kwq7+rNAutCcQSz36FD9QLJkouPblmapkpskaCaEkq
wtbjDnj/mkWAV3aVLoWDNl8NhvHUC+l36z5VjGJOwscOoeFhF8fSKEZRuzraHbUT
Wjh64yLNeN9TR+fhCHGG35c5qFaJIhpTcEVQm3NoNfxLdZr+fthn6vn3o1owPKuL
kvI4segzGaEmy2Vt6ZUAgTN8VBN5CanqKBsyYfpz/JBzL5dCDYAOb9nnjP+Glty2
jNk+PYSYkrcXwd7tY4aesfUksqMhvzu8FMJtAZouGnxmMV5cBtYUKWFnrIGoCjru
yUsF/fsfDqy6ZqjrvcOM62Acfx3bEwI/3BJDERMh3RsByVNUf9PnrdoL0+40aPbO
t85zvZV/ajukc5pqzgKuci32dmSju+M/LDgUcTzSJ3Mz3DI2iX7VJTp4MECPL+Gf
t1/E0445eZtzrevz9+Xfbv1PQyg3H0uclR8jqU5OGo3m4GTlQVulJXQFDlh07R0k
x9Koj4aQ5sFAL0cNlUvsJCh8GByk6n5LCfto9bit40bDgzpZ1TvOPHciBPHbcE8v
xtiBfKYO6h3GovNz06NLaeNNyXGgk/KeVQocjUAAz5Qx7bbwaqZiNGVUr3iRrmFa
mKofFyIwBOtHIfN9eO0sCV37gZn9rRaUvUc8WRO7vFC3wez0kqZsp7d61dEAyVWZ
o1Jd1R0XhbaVfPMMf87o1Uh0Y/O3EiwXZ1AmTk2zB5jyHm9GnfZh06HUXL2InLkW
egAXk8U5L8Ql5TBaw2W1ZO/bCjYD+kotiNXIxThlpLjACqhdzslG1qeXMu41zwOp
ByyuXz6mDjCzdF/Uxb3+wKjqcmrwIdfl97DH2cC+lUXD8Urs/P46F99KZKWJZjnw
sA4wxhGrUTDZHVvHGYG/Hhsz2cJUZNr6g2Sg+I1lp+PIfFMvYZiL6BFE9l66bgJ0
4/z1RJdpn5QUqo+xgHfL09iZNQrpW6WKprZ/D/FnhJuERhTiK6g2ef2O7ZKM8mEN
E0EJOtRylKHiiL/uVcQ1eviNaHyk1H2pK/eUY8gV80iRFEfTV/Q1gkuoHzWn2sZN
JoSJ0+WZIDGbnwy+ZpW18gaHKDcLwb2yfRWZyupvH6SqHYcTkmG6f3AdlV0r4eKn
u4HxiU3khWdNLnPIHa3imYy0rMfGPRqjt4jm2Iq8/P4D0cr6dxN+gQLgoWbfCZmY
WIZ/0pIwhaVLgv3etU0FSk/4ue0P6vLQTAx0BDZsSgyrcAWDkVB4+Lsd7n4JRuj1
62VGuEq+xpb2eTT8lRiiiE3Mjy9fzVHMm8IJ9hu7IpMKyGAIPdMimC7aNGRAGJth
pnfhpNfxAHibMAoYet9WmuHAtmxKJaoPKYuLwhF3oiKbf/dhPCIAJ9xuZA4Mdt0C
FVoEJfvvYcnmqC01WJDC4S1wkmjHK1f1pM/nKs3ihizeQXEWyrdQkDIHfo68NjVN
H+JfKWALqISgbnI00ieWc8nO8eHyM555uMKro1nrjHGUABb1sGRbrKN8jylkfryZ
gG4OQJBXqdQE4MWpM0cWAimLuiokvOhRuqiwINrz4ZGV6ZI9aLQ4rdU8GDf8km8U
NOK7g7JtMJCPiDmC5nzhEENQbDyq+OLAN90Ime5rKBn8VLcVBEfXj7LlzYkLWH5q
zMBCGQU3PMk4d5KKonAyx8PjrGBcW3Bu7OFQ+fG6EGeqpdnV+n0BwOQh31iZrOPY
8X4Ets0pUnV+wMZRGMiMBGHW3yAdtF+Q0bJb54inQyZo1Vrwaua/bZbnN9Jo5Wl+
79+a0gsaNkcCZoFVcgGPyEuMZANXZkEJhkYi3Br5aJhhLHQG3hFEpG8sjZT2/Qqe
V4tYfzlQtXUHu1e1vc9groK9qjZFG17pbfpwTbFtM1o9h0l7yy0RAyi01yaIS4nu
eHntvBbQyvCB+G28ZYMiAOCpzRr568eseea8HlWGWcEsn20orQuvaD18twOxXy2l
0KInuUYaTjrqFKLUgNAr0f58G76V97t0HhGvCeeggPQuWaSnJwQYDB1/Z1ugCrJf
4dVTx0oI+2H/INb+0gzfjFTj8DMwxXFOmts7lK0/4OJFak7DNyZzhhYdWOKraxWk
QnQpzAkw020R/8d4T7yesO3MiY4dJnyhmsxyFlVbTf40ckOZQGWXGL3y4Z81c0y4
6QXCkrpzh+IQZyryiecYtHLCtWzoxdipHICdm3y+qXlUpREcL8iOyFWipkxuzZcS
VEp3BiO1ab4y4yWMdEINQYvE5DQLOIP1rc5YQRmzlfmOEghRDRV7+tI++8/LLBH5
f+h0pUvhJ7DGdaRXlmKRW9dy/fUKNEc8KwOzqgeAOcriglZrF3yWf0gWOgR6RjCC
r1I/7mloqmiBKIRI1c1jrP+C77X/wcAjiUqL1Xy6zuGYvkSKemDiEp9AkLN7QFDy
oNJna4prZL5jpB8TNaD3IqOnS91wTh7EeV60v/KO4Fkc0SSzRFZSVPm24iMcsZYI
QbMmeff6YACE8aOa8iom28K7w1n61b9j9OOXsu2c1pnY57euHmbf3meH8P7xPwcM
zKMnYBPRkR6oCRojuziFcFWlpJkIjS+kKjYRqlUnXLw9O3wgzBgQeRCLyfsQDFoj
vQ5TML/nR/gpFN0OUOtCaROiv6fINSKAT7oOw11f8qLQoBRsh+VXYb3RNE9SHYjr
UdbCTKMN/vqfjiGQ9+DtkATmfeDHQH4XfhF6pS4aeIKJxm/AuY5MTXMaKwELEvja
fMQ88IyOYRhKd1wg3HJy1CGC+CNF1U8M/+BwtxHS8arXLi6BQ/JbhOsuy/afIiH2
womy5/L0ggn0K5fC7u6ihqWtwrTD1sKywMS16zuEsLIhLAYiV0cBieTSMG+JQR8T
uwASoGUHmVqJQ/xBScnfnv70rP4Kmf5pQ6edmlWNJ9MnbhpLl+C7I2A0GRjR5rRO
03BcViVV49rlztv1KcUhsEnPZzMKk+M8gnWATOYyT0HR2nk2CTKi2xvwjJkrp5ed
88F9SrOjY7TYSgfnpcvPoL+z9kQj9TP/td8lRBdzK1WDWC+A0QuPp5yKTBlnUCyK
SNeaDjPyTvsAltnWTKSew50z+2DvLDqdgJJ2pmyYhI9CiTfTLkKnAMSKg56GGVqJ
hhfdpl8gMBtjJ2daJXoYlU8E0Hb7C10JzTYqYM4kvN69FJrD9Sz5+KJDmQokkJB2
ze9Vj+qYvS1Ej0CrVBlFAB0/Wr4bLL1od9a9vKgnJn0LCBXYRytWMzug4UilikwL
WJN2Tw9nI4k7elZOSqVoLnvq0ZZtanswHnWYolmW6BDJplUgDHm/okNnwvr2BkXT
5akDEoQLq1iZEqOZn/TOlAe6CEbKXdeVaV1BD31sNQSGdSdM2WVE43niZk8Rn35C
YIlRanGeoO1OjXnRu52QwWfh1Sga9WOTzMk7rsPZ99p2XfFDJlZEgl3u0QCpcQ71
iatiXg6YxSeO07MYpnV43F4aI58fnhn+jxrEiXtPAhvk9s4N/LRSJl5zppwLmkEm
/8pOfbk7cxdUb4linUGp6hYeyufqxxHatXQ2b2syhxPkYuJnK/vg/V7jTWsZKUsa
wbGVstenEKwmsmy2+RoxfJFqwqT760sZuNCArGOKGub8c7hCuu+MOK734gbRgW2W
RGZStaWO6jd8a27RFbxfeXNp7IamyjG4a21tJ7MJr7Rk2CY/3Ei1W05fMSXbjnj9
BKvoIdhfrDUSOiVqN3o7OsKXCgd9bT34dso1oWo8RgaBIi26HT96NUbIp6MLH5e0
frArA+Ulh2ArMJqUE+VwKV79XwIO3vtcEw6d3lITvomJYxpYXVLS0q2rR/jh26Yh
q/GkfvNdBuXEzYXL6R/to9p/1PMiC01J2QmgEe2kY4vSZjZsQe84JlJvQUJFvIBA
BXZsQ4JSHUIeeY0otdzpmWSaq6aJmj+1sG7QO5fWN79MetS1SbEVderoti+D1Nrz
j078vp78v/mujGHz6tEwCS4OM/vbi64kuikS0JxjmmdSAdsrTtQBUm2KwfV6eUe1
PLqvzWmR0zAbluOFilAlCw2s62j9fgfwp8jttqnCsaGDgwZRhTiq9WAagG7KDTfQ
CqyXg7lkO977sz3yGCa9cOzT28KJVk6yqd5FguE5/FGqS9thJCGsfj7WM2rABqa4
qvgWOQ9z/leTiMlYd9NMPDXtXwb4ObQkXC6QEWIx80+hzQbJg+KwbVgqGZzoRb7J
INzvmzxPxJKxPMBBD6ACgDSUlR2B4gYG+o9XQCt+YNN1GSt8EPKbCWz8/IGBl+Gu
pd4+YfattpXtjo/tR1wGTAndI9/QlB2LaiVo0fGuQbydLeGB4CwAQiDnAFqTcphi
66zmEu7Z+iBtEaNBsdiHU1ROxL+UR4FKPja5hMaD8zTetlM1rcvkJ2ri9dBB/Ske
NCbpuMzYL5wWv8sczNV5cDIImGSic1d+wduP0A+cmzoPfPZfJaUj93U2N6EFAhO1
vaIjl1EtgxFAhf8jo/lI+4E1Kw7CF6L+LIj5S+mi0vhgCBVXlyrTSMLY+JxzMkw9
jl4zwimWtg3jSChNsWEzHcmFOLl1pNBP8Xaa5woyLBCvn33vXqwDmULCCMXaGWQu
ryjx+Px5i2ZvC/L4jh/82jhA8GQGid65tp6GDziNulQMTNT2reqkwkKOAmPEJaV3
oBLtREPqYUvNpnRDdzXhCp8E8LePbRyzD4bmMeyfxUU0IFchg88Zn9ZMwg2Wcp4B
VtloESWe52Pu6HAPVSZDTxfvw3JdDGNrkf2a24XSmgp7y1ELPIieubhFUlKM9IZC
9uzR0NA5dVBOKqHNbpj48GnJLDNeE9Zihd3aWcMtKgnOhsVt7MV0PZi4ZpHlC+GK
9D/upw9xWpad51PKkeCNWdSUSOf8Kn/h6WYWB82UIz28xKxI5Ausc201/8514kI9
VdtaUdRewbSJeWHBxHWg2djcb6XrPdxDOolwcT1FQL0322Bg4cQdnP9CsfQYy881
wDeYIX0FSC3mhca0OldliT/YzEcOma4c/ruWt4G5A1vibY60gTdNQ8RG1w6QOWGt
kdeBE7T7VY/e1oOTv3ND/Z5GGS5DB7BGJw4Zc8bzoFuHLUXhL56xWa+IwuU1h15j
3xdVbmeQhNpUJ55hpr+1ISntS/XqVU1vntHXvpEY3Lf6J+7jwqI6iEiTTZzVxau5
AAOjRO4/wZlEdAoUS9CO1DVqUt9nLnTpYXeOD/OYkKy9sprT6he0D5FuLQuo7TPN
rQn2TtXQ4xD5HC1M5E2lA+sy0UuGgoYQBfCpzCp2nDW1UU8FVlrSAZ6jxx430wwM
eqLd3NAiYwx/3mrFCkmGsYILt1KTqOU3PFI5o3IMrOx3f/ux+1+QvHfnRZMrqbks
2E1kDb6RiVqCY1A0TnuAbw6jT5t58TZI/fopG0Pfy2qSL1BPjUQUdRIBGh9ujTIK
DBsWUi6o5I7JALZQhaw/RA0wwKKt/dc6eUdHtNYAr14h9O6XlhXPtWu6OfbsUUdc
/s7LLz9iXTEOUDQPsSPxp1QThJJipg47AnzYRtVJ3upH5UnUpiJAPXht+KmF6nXY
l9dGCSNE9DPDmqhXJVHlw6wjC0Z0qEZ08tKn9O9dmSvUnG7fv02/0EZ37UykViva
k9lE3dPdzVNCCno0XnqJN79IORTVfh+AQclG2tMfRiFrN/GuZRrS6rXGRR162M3b
SjIc9BLsxcdPyEn8hVKChuqYJdBjUeY2mnZDwTyBbsWt+8ayTkU7pYjTAEF7FttC
FNx0yxB5aujqgUwlWvL6DsGMC/LiLL540Y/sVe+/PdqH/GWRAN8d1pYzHOUnNv8o
DnYSBtrU9B39wO58PanThuVvjg42Dl9duN9HK55JTZsTKTIVnMQosUeEkygcqHwH
45+X1u6ZmNLp4VX6P385MGQBhisHiqyxoaecdtPCiOqLGix3W4deeVGPNdJur7/O
hltx7/SmeMcdRd/VD5OXPlZ9GfBpnunuTYP4LIARoz0jERvkdXNwym8nOpZYYHoG
DWJ8/Alw02/e+ToeWrw3qy+C+j12YiIeAHhxAe1Sp0i5yNIQLVrxBkO7m2GC722a
Akyq3sTXaNsl9MrnhzTrPYrO72cJ3+13D4kM51npIgWC0KtvRsZysZanhhS6rPqf
30JnYroEyv/wAbe66tuJEClbkejQEqdV8VMT3Oj8oemn4PKxhRZRt6nwW6vl77TM
P0qZcz6aBtrFWNObMHoX46D4f693e9nIvNF0OZiiob/uHPTmrBT1P9PfcJdJcVdz
nLpY6E0f36kKxEag7d/PdKxcA6FCtLcQAG+CRACclo2Bc7nHqtTl02DKYJxkETMr
nvs2fd0QSXPBTJjpeaQWIxwgTU6875G4HwfXsWC2l3R5xhRjFge5sIiMzZNJPIMx
b5XyeTNreQs5ZlaFJuqb7EggUKX6zG85JUs98LkKMlwm/8RzkWck9z1Xk8HCC6OD
59vrfu4ig2cseSsFHVnMqX3YHWKexE8rYsu6X62wLdywK2KRa82EwVoIiDkXyBeI
tIJXTOC8GRz1dYPPvEGKBf1QlYTjoA8MTSUKjpDbZklR54yvqZFNwn1cvbeSLKJ6
dNlZjs5wLoWgfDvROLZRTp38a236wXlXebOjQ90aZuO/d7cWiDrA5xkgHhsvJf/r
XuQJAlnY0EuAnTcF6h+e/9ePfo1l5+BhfrI8YUyttydfWHa5v8N5gFOWJqUZvi9Z
XCxt58yrEiNBxtImfWcT90bMS6X4kMwKkS59/chRvGpLQQ5VYTFWQHQVZGlOesrE
3uGSE1vAZ9FHy2VyI1DItoRuWAoRfzshJenCOrP8fyVPqUsbN/RC3FZDPZFjZSd0
W8hyyh+S5cgBhWHSHvEdkRFoWcRtmcDGCkawMMvXfKwhExi6OwAmGm7JzMva9UdI
BiC0JnA274z3eht1l9rMK8eL46YijI9GOfrOR6ba3qQoKVV7fUMh5azSTcknHpDJ
Ql3E7xUwMDmo38C6veRafClHzS+1p4d96apsITUUGs6ie4QMdbQ/u4JT5kzAibrE
slBRxfrVFFMKXuXgULvHEERciPmKTmYt6FKuQNw9J57XDRTiyr8Q2urHehAuKMZs
eigHiUatE76F29ed1WiR6l77ent5rexV4ABMERNJoHbZZMsTd1HJHMg5iAWCAQiJ
1ZCim+4s4Kw2+siILESHSQAak0RLaViRqU+RWB7kNyBujnCyo/i4PbgLM61Zxj35
ooC7bDukvoG8YuTcljbRzIf5IOPGg4jW9u8rvCUkD0SKONCY6bjnnDatdKSZy2ly
lhfYq6oIHiaD9E5dyrHS2hgRB1duEgCp1uAsaTiW9w82DDATYHymdGqG6IVwgMuw
nlPUmWZHuIs85RTKoLXf9QRCfrqAdgpQm6ivsrV6T02VawYClHgOF+xRCuARf1xj
K6Au4ItZWfxpalY6B5cIX95JaoJ1+oTL4W9oZ57nz2AIcANVGzd1d2psF1tcl+bn
3p3V34xS1XZeDMF5vNGRc6z9Wdx2Buad6c+/gswbpF5TJXYl2NRFG6mQGtNFUW0v
oGIKH0APhz1BVyjXCLu85zeeoCiGG1z1O49WD7eeStEFP1D5eX58uSAI+vn6/JSd
a8RH6B1R03rTYRc7bXqd0fpuaJnXun9NXI7Du4jwovAaXEvuU7IqudgigPKtx4Fk
ZeXNBZeJH1YDl4EXyuk11JxUZgSN9VTg3Kf+zkCTInCOLR6lGaom5L2YOjqB6k8P
21OjTaoDbMOkwA1/TpDZwHpqZMa8B+36mGhVgKUHtjn88SYzo72ul1e1LvvX2u/h
d9qo3xnzTUqECgn5p/VUd5q5EEtBEq8l+TU8CRnpvGn3b6Tk6htn+QT6FVvttDZC
BXXPo7xEpjIluaiQX2hAsyGhu0C4YnuMoF19w70k659YDldLQ7DAZhPuOOkicn1z
Fvh696ddXEimY7SGyCixrJzQh+1IQ/AtLZL++Tm5GJus093kRyh2fP7kp331JxpS
tGIiWxdTpdw9ohgLQb8ng/L6bFNZyFQ+1agiLIHGnE+nBx6wgfh62qAxsY6dm4Ja
Oal3pX/sV4e9n/sK+yl7xbd+MOUrOnTn/Geq0h5Vn+/+2EN4N1s48uwAqfJFEeIm
RW6WdeCXL9Ea4K0D6Y/hyZMTic7S3z+LniPwt8iEnMNDYciW9N3iPX4bL+CAGmaX
OFCC3InYCEzzWtibw5h7AVTBLV8W2sLOlrOPrPSPaFSa6WL56fqVL1fMQBzU8dhL
CzFI2O2BqcTMgLhC+/mJC28SgN54JybSqt8TkByR52clM2V4ml+9LL8jmesuEdme
IcOWE2ltMp+RoPNyq0qSsich0HtzKXBygnzmIRfszUEim+NZHVfpba3a14ZWa5rl
G2Ve3YcKM75Z/9ZtNlM8+q1v8sLm3cKxLsaqZt3PG1ZUbz4aKUt/L+6NHrQ4hdcM
6yunSkcfvrsmSZk0j09zxdfDYFRDZcITGWkz87Q5+lZgTHwZnTRMt3nxXZQoC6hB
R1HG6+O7fgsQN+/rq/CPvj71bBiOA/jLGsIepibZnZp7e08G0wRo4JX6V0F9aB1m
0DjonzAoMcYpr9jFy86+Ytd8UXF++nR1j9bfB6Q4bgpvxibGtLpJhuU2OdZ/auyo
XgpxTWTB6QHVC9Ma2fahPQqoH4qQYgAAHjVIg3fPsh4q4cD7Oau3SWM3uaOa6wp4
nqGPz3vYZzKDnDIxo52CBehvqmvOhdvd7gt43T54541StfCKFEBO0fYc1QGxNn/y
bI+GZIrVdQXx/AGojRDFwIYuyq67u86IRV86V78AuQzcGnzy3S9mqlESVvoxHhYb
+Ys6yuOpZiyE7qFnEKqBNeckgDxxLXhyDgaVwYFq3ZGIkWjJuy0bH0yyvJqxJDzb
SWbpaAzU0LvAtUkC1nIzbTdXNZl4iWg/WJdoc5Ykx6vJlt5EokpTDMGfLDgP2Nz9
YIY8y+D1HxN6E5JC/+8DpUOzflM3JltbUfzlGCndAtFWaWm60R0a2iizfSqM/eKz
Ympzc4Ob3viHIWoGvz57Lp4K2IAu+2tuVSFWGhw0PXDQFaVo9jzlJfMV3/uWjO1a
asbsfZJ1chAoqIqPF0H8lWctsDnwPXI/Y2h1yx9GmfFawBZOIVhVHN1iyX2Qy4n2
eKjHAcg/zZH9i4tyXoGhgTwtKBPelrt9fVTw2BA6Gqb3985ty0L+Cb04wSQKeGHS
pllbSvWQ/XsyMzua9eqoEZ5qUUudXWsEHb+fzF8MZALDXSYKRcV1Kd64K32QMB60
ipYX1osZxsQpYD5Ie0lfN0DMy4ODVso8A8EyCXCRf3HUXoZ0+fIYylr9hlzmSJY5
qnt921XputdVsy+Evn349Nx9i1nOW2C7frmuIAKHGdIw6ZB4SfONHvC2+EF24yYX
nXc6/2RqGTsTKuwHQwSlOiPPQ6yo/TtUH+u5F7IMbPObYvU76TWZt4m/KICMbJ5S
5ySqFBzUU4MaAEvVgnpOsBYRm7QLChjL4aq09iSCNuTaU6U9a+FkoGymY4OtyfJ7
xrD/hMtBtxj7Hr5DCXn1HlzQQ1W7pji604w+XD7NomJ2RkWh9cCrzEMINj+VXIPh
SgFIOUejSTF8aqymc01fdoMBJs8/8q1q+kbgApUvSME/mUnkbSwen/bF+odiyPuJ
CBwwdwLndJJfKvnh1cOwxhE0EEq5KlDpSJXF2EiL7A4o20PpJjKrrL7gqZl4x47A
Js9oix4TAEQO9vzSuGacj8njBBqzbgH+1FWRRDD2/7hXHv7kV//iFm1HvZw8OZWN
ST/vkw5t6vKHkUahj8YCvXkGmM4/H0SCmGxWtMcIWN1ge71KZKAAoJZSEq1wByVY
SzLSRC/LvLRujiakaiwuDyiucryhdDRx6O8b3fOgHzQZDYyG/NunaWqD1XgxjZgR
OH5AB+7RfvQkSq9ShAsxRKPB3KUm+ySZQ2KJSNbFX9WmXqxw7/xg7luCYsjeuB2E
IWmPH1/Aa8m3+pdSN5JlWZXtSP+bFVowqmTQd0a2gfsUJDr15qUwmZh1xjrzw1vM
7SQcHd28t5jlHTjEnA96p0ybgYd0pzYdxi5w8wp0h4IgeC81G3DUeqMmOUVAqb63
FqN43eOQdE7QRDkgucHwazISXct2x3UgpUt3xQhlc2kzJAMEgDRD1vIij6HRkOGp
aMbnxp0mYhf8jisEmKqaSo1O7OpeGVs02MPOodjJ4UaXcdArz/rOhsfyTuayxLDb
gAr/8y8SP+GKCfJ3e7pMWgMOCD26xggyNjIatK46q5apkKo4QktQaM7Q1OzRdlrk
fALNiRsxcXHwSrHqCqAqOMLXWdq5N1JQNtTm7mPxJoWqEMCbWI5/GUhdaFgHIhtY
xNIOGCbr6r3KmXKrUBBUNJcicyRjUWGDlzoMoDLPiBvq4cplP4STSUmPWSpV6MMb
BQyPmMjS9r2dNvdG9dXjR8uDVKt4qIYneNBcWRkBZNUXQHjdLH8oDfcHQMsgoHaO
uzY6i5IXxHCYRZXZWu2WtJHde1to9s3vwYPQmGaca3PImgupDd0UH2Glc/wXm4hJ
CWmPUQegi46Aqd+eucKWj/Mp7WNNtCBKEg49/kVq8GY2Fz6g9sSJHfxVmhOH4gk4
gN7wSJtHX0B6mv8/CT8x18w+SH39nSWk30N245HGHXJ8v5/ACjxAf7+kJ5xPsaYn
5qtat3Veo65rb30Z7haigIszHrBLMITbF/JKrrT/inYvr+JemdysdjcVrwWylmDX
Mdq/dyCKhy8gJuEpmem4DfLPYyuuexahiGNUt+hUOGYrrIyrCmEA8LVmo0+gVXPE
2KXyvcG6ZDhybMbCjoe5VyzaiiZnfoOqf/FVUUm5YAueTPvHCdTgGjS5ZMJ5mm5N
XYwzGSaKsLnrnoCGVSjvqTP5SiWaLHOM3ALgDmMV/gb6kqfKizPPg25moI67+hU8
1lHoaweyRR0IWWimS/5sc7j5PxI5urmPgsgyfHRXd3XfDZ482eGcCm1IjdXKvJ6Y
SR/XSsB5pk5eZZ6Otbb7kizJrKu2hIkly7g/jTCjFLpmDnFh+dh0Jf8oMZbGQa8b
abx8qmzL8XU03ahnyNAVMydsPshzWt9Q7KWFodjiICpmAUoGWin9Ep/9Fw/L5gbD
Bnhy52yF1kD0ZYyVjtI56JM8LiWEgFkC5xWFSMgM+UMKVbzffVZ362+zs4I/4C1B
PMDA6J7xxj1FWXGnz0kLTmsIY0mxwOrVKuWp/S4Dgj0nuAepMWWZJzWrKF41sQpK
SrbxrzUATXXve+ZxHaISBfHj4nB3bf9P8lR9Xq5invrV6Ddu8VnkJsEhz5RF4GYH
Q2oL6AS0/JNjMJMeEFcxOIsVMWdWNZhYO9wAbQ+MBBcGR7jihYryFGj5ZFiN5ytt
thNLqsumZqtLW7KQJaJyMFbP9SVlZMBoRKdrG9FrApMsognxHaBD0hWDmky8KL8V
oSnPLRl88p/oo6PKbgfWM2BtPRfXuN1IlhB2cfR2J8XHmfLNHLXnyIW4hqZxxDp4
aIgpmcEU4od/7NmecPEhVBzBZi6k2PTVWT3rCLvBq74WA6YVgFsJ50RY68MpFMoj
FiGvQFwZjQzxBkiL7uEsYoezgBD2YATYrNk7b2w6ZrcnWylse3hFHP0DKHyVmdGR
zmQj7zQNkQvshLwZ4gnsS2AjexlR24bpG7iXZCQsnw7QHixDradq0y/ZCF/hYsR1
MHXo69aAvU1u1qo/Rk9iCQ+VBQLjSYP3EEzz17WMynnj0BV2WJtZjO6XdegQltMR
GXBZdEPUj4je0qQph8qdeUN4855XQFVKfp8STuhryKNDYFl0WPUtI+bvbSFCMAWQ
jgVr3Vdg1HEXxuu+sypOf0yNLBiBa7VfsL8nMhoHr0KC71wmKlXZVt4Wt5c3TbOz
Q3ROOYG0zjMd/9999zWxfKtdTU2F5FanP5SnqdmyDIvm7OWKB9jzf5Ej/nCwD1NN
lhL/cFNYFC9Kd71FELRgoJUR+m18iWZ/mUpj3ib8U3+ZDDsXToPIfppdUKEcicfX
NFK9NoKMy84WnjXZDVcwwZXIU8reSYod0EEzE5Pg3po6SyQ+YsyyErha8ShknXAe
zq4EII6gM4gERptP8I9UO2DVIWSTf8etnZG/cffI3vBnf/okkhqes7v/1QDlzC0l
Q0Nei4pblCmA0yhYLA1jnApLXNuBYCcPY9K7FxIBiCuRADWwHlv57bsyZtI5aZe1
QLtAAIxiOh6OTKbp+yeLKVMMXWhq50/gRII+EVNLwKWJL9aZUS0Dk7frLhdQ421f
XW+MIufKcsuaBvjtP9dkFtlbEfLO9mHC2Q4oiN7YOfE0d94yw2CwJQd0irefjIlZ
noWE69Z3FUIc8V0sJx0WYEWc8cBYzwZZtSh7qeRS+aM2gxrULXjdxQBWdSD0huiB
QobZdQU82+n8BQhUXqItEvwOp3L1VfJsGwrRyWQCIi7RnOB2NSbSv5MEDibRJfGz
xp/kpYxcIKDUbQ6fj0jBt95UOTvOzPiOu2zK2wWM58f6/aXGxSdqD5agsKqL3G76
Lh3c0OW2XRnOOY6Tlbs8nSsVi+pu6DfO+jC7h5L4j6wDWROxTcq08oLfa+g3ZoKE
AnEEpLWVvBZrqVc4nKgcUi/imGa1TrLM1hKIlPzlcF1jdI+HjebeDld8ZZbDzN4F
/sPyaWiOVvhPX87MqbYpj7/KcS4RFP+zEoODicXX2uE/1ghlHq42O2CgNDLsVSlp
vWLFYquIdUSXEir4DdE+Fz2kzrPXpKxi21KeE0O4K77+iFTc5pkN9wUW1qrM7dSl
mALSsELoDSHkMxV2gcfpLE5KNUvasDmJKvEM6X8DuNA1hiDtU2NG5k6eJOHzCDbl
/rJkAnvQGCIPcBhV6RUWqGuqV5rNMdc3YKQhJwBBUc3TjB63Aa1KRYKB7niHXs3F
GqacsPZD5QN0sgkk+6fHQdLa44KVtvw9RnvkIrJPsR8Jb435N0rqIjDlk/AkMUil
K2VPzGR/xTsLB9CsdAwl7rT3MX1xdU/92NQBhuH5sa8h5oMC7+wcBk/Gt1OAc8+j
kL5iY6ZiM/q+lBZAPCbRIrnTT6LJZGo/+jcqAJBcS75TXE9S0f18c/ifAfSqgxc0
yb3xPJyADwxpLGipfHF3LP5AtxjB59r2xu208nKMEp8IAekprRiWuFnar9R7TsV8
H2xxw1TZ3JOVbJvo4jTPGl9jugUXvvD+Q/bHDDAfZwO1D3TiPDYg2xOQe0PI1QPF
eSXToJdOpPwPh6gh9SLDM8rxZPON3QwMX3eRbL/+Y3/ctuLSnpO1sDrtXyZRhyzs
T3tg3kjL9VUaGrnlEgk9EkE+7v1p+5bhsR0bdSAinjvGAca4kw5nXEk4cRwGbSor
Jf3CM6DekmfzeI1Kpm0JFzQNWhiYZEx2L15IT3R02esAyGnBAoYPEGs7atUh6BwE
GNYLD67GrSt/AiUpIIzzdIZZqOGzUiv4cA8TbfY4USs/59vvP3XJXN1RtHw+ihcQ
eTdHg+gVXY/NeMPFSQV+FqpNc6Ae08KDSN1pUOIx6R0P6/kE/2IVVZ4P+5WGqhgT
uN0pRFJiHmJdr++aD6q/Q6OKvWUV6Kb5qvSSmzlDAy3e5dvojKuqcObzPlelyzN+
lyILt+pUPPlK7cD3R34FIsoB9Bxo8j5WJucwBav7lGQSL0QWqgjKJfyfwECSQa6J
TiLnzDY3c+oyNwqkoW6brq54EPvU7y1esMK0jwodyqVBsmdfjM9nWhZYIVkvRnYu
2xYBucyMLcMZRsM6w2ZW68avr5B1GygIDH0vF4PXdZdcYy3N4xEbdxJeJtIDl/xO
QuBrJ5Rz+tOLIS7B+VFVFEXCWggXclda8aO3OquMKNnTfabGWjS3NzcAezRcl0TV
FqekN32W0/ZO8LQ9RI80wPbQjmpdFASXni2LnPt7t2KqeijkF9eHfbSEE4h+zKYS
KSqQF/ranrXPGSdehOqAT2YzupRYiztAVGR9WBj5NmTFb4N7iZ8q1qyIZV12mVb6
y2YpAF1toRLzSwu1X1dkDBdDTI6gs5goqjNBygiJLrp6Xn4vAW/m9ZJkZs9YdemS
/3t9H3l+6Mwb6oPtmfaHj6Not3BIt9sfQ94x/MP64U/V4vhZXL4NXeFgswgfuyLY
fnVk647iOMjgM+XQsXZOc2czP52BFE8Q/ty6+ifull8h2HvmFyparqFSi32IjoM2
4bh83c/w1p6Nv93jDl1O5NLxKKmnyBbXBHI8YSp4C693LRHWW0Z6yWitCE3gbW4i
B6wVKa9fucQ+c0mSaWECGgX0iRjmOqvjxMk3piJnuEAUMZiLPh4yjY98cGzPDXh2
12EF2KAbuUCd8vUj5w4OfVllYlNCTbbUy56nVjAx6KuSxW3nWewY66cFqSaJRdb3
iOV3hpWC6xpnZcZ3ujV6y4VuVTiv0ab2Fj3XP90UbVlBT7QqFHAXjkcq/YcMgLfT
OMUUXmyIZpB0NW/S4IEd66OGCJhiaurvZUH4cQY0cVHm9MY+HYIENPiUnxDbksAF
Ll4BYRh4eRZXT0QXKiPcZNA5jMj0SxQxBlP/gMzlyCfkXPfzUI9pQ5flA+/UT5eF
XP521SOM6KhfsqtWHA1oUdcO8/wsagMErXrF+Zki+oNGt/KhsE5wGYfj8em1lpp7
Q7aKRGBIYEKDVEAoylncqhinVfonzUVpu6Wlw5UJCje4KEj7MvQJ6tt6tlpyqjYu
E2LjM7wxMvTNJOBnpR32VPVPW4yEh7Yh2dZTxeymo2OTS7EWXNVzCw4UJUJW0WU2
y4OxRscQgZejq1v4RI70Ag7zNrVrqdOYUrDKcxji8BCwJZCnJmzJCvBr3Op++/YH
YD6bY3AQTr87CaqF2OGNTKFhp/lQtaoRjT/ZCGxwNERfWjWBvsF+QU+oH1VDle9n
pDcAa+p1qfPmKMBtOru1OmnRhYAub8ZOR9i92ue7b0BWrhWZYX44MUGPBL8W6ydv
6SQJIZBU9MZ29pUVSyURbZao+f0avV7otdEX3mh27YSBS9HMb061mYx0Hlw8flrP
x4ETr8tw8MFfNPc0tJz+G7Mq9ISK7m1lLGRc7DVs2JStITKVwu+u55dRZGJgo6Pa
W7yVcpQhraI0TYR+n1ih6j6YUygcJZnHwrleb7An3j9Sz2eJywimYnTAf/VBJdHJ
K/c0DpYd2hdMHbMWBV0zf+t1Akj4g7sqXsS/xVDqSOTQDgVryIJYCaWPftAvgWaG
YV58r3nsOZJ+7Ohkdm2VgEzvTCK0Fjz9ZUMBTnmiBxqfnEG7dhFc8OHskUwJI4+U
4FuJTR2Nr5EK5/n1If1aZtiDK017tn70jsvg7EvsXi+C6/pk6Lrhf/Cp1l5nVnTX
NeTRJp4ekFybha6U5DYdO/ZM3Xlm+67yxs2X/2joTBI8SFfUCYb5jS5Q7A5IQEib
rTwCdbzhbKanHwqiWq83xp+Cvgfhba3CZHXCOz0kYkfue1tLB0iTAvyvs+brVmwA
82QlcwtQ73TmDRFTJJo9GabQ3QVoDZGcyecgfCu+sLe79HbGR3QHFP+NwaPVCv5t
oJh7mP+eWztkuLKM+L8rx5ZUBybFqCykwSqMFoInkKd6S/vLTRZm16KXhAIhPqKZ
SK6prxMLlBivDnTGrHuMMER54aTjJ30O/IPFRLxvkoOhAPSESbE28E7FFbwlGxac
Ev67LSmDQpwAfy220I1uwdNqm/bcNrqwDDyVc5Tnm/NJTOLfm/sMEaFDp4aQy8lC
KbTmTPLz98/yrDSeCt0Xbrw+j8ZLdSPCbe8Pe4nVsKoA+jrwRpbu4yse/QpDggL1
AXgmWLm1bAMU9FAWsxIZcn9Dfw5pqoEKjB1jRA1U3OQOvL7/NvX4uNVVY7oOU1v8
ScGhIneatmZM9VI+H5UYfT5sfo4Sh4oVU9deOCz/nlTlOxpPP/btGDbeWr138uMe
fBPNrni2jOO38GszRSjakWKmRBeYOYett9sxwdglKg/wlu/BXO7EyWos2ZOlMKuP
YIQ9VbsarVtYlOoZGbbAEPC8EZKO+nxsCmPJuJkXaqTCSDEc9CJNCMEbhsvuKmq8
/fp3g53hPd4vT3qlwsxg4YtvLJY/5hKxoqg7mcaN0YDIzIv5t1apx5w1xIimecu6
0W+9zoAdtAQqI9Er8bJDSEIt8e78xESAKhmSHlajE3IYVgE+nIPDAPk5AljHHYEP
ydDP1to1IPyx2MqJx8/2pUOjk125oNxQRAyzsufeCMqvfTONzJG98mCqwOS6NTfZ
UqQh+Ui6BoopHt4OD1oWOpViCnhY86jCQU1DC/1pCH7KKReLIzk0N7CkIiFhTNRB
uLSpY+KKHDLOMcT3z8envTdrigy2/SMtZDstxl+Y7RyQohInyfWeHxglvoWraRB7
Co5z5wOGcxyG8NpaJ/vRThUmqoSty9alyK1GFiPHjrb5KeAAtDgY63+U5Jiio1c+
iSvN6Wc6xhjhP8t6M6XbEoU1/VuzkEhd8mzTLS4u4MIjvI1+YGmI5PP6LOljb812
wYzFVlK15faasHejIFiNZma51glHUDkhmDIIs3oa6zNZ+4uQ6Kb4mjF61PBkiAw8
JTlonrgdP5u4kBImhiDGK8mqqQh6tcBLj8NHi66TPn7bl0IQvh3tg2BSOmVcL+TA
bJ3DdaZhLWbUoEPgWjgXIr1USDHbj2A9f++lBUUysDTAEboYrIDx+IS6ZiHRqM2n
/hhd4sDJ5tdyOIkKAl1lpLdcHbvsIWcLaIt7TkbGS7KVd1JKiiX+CIrOpmaGHq0S
v5sOS6T3vgxapFWWgCz0jZyteatjpZkgJN+dkoHmNkTeUWBb8JCIAVWCau08Ko+x
5w9JLEVFi0/Z8/gqn+lnxk+f1N4YXxa73li2CzSFQo2sEFitGn+IoR/48pWVI0ow
t5R/5ul3cjcJDJouogCAO9uyVjj1aeQhCTRIQNYUBjqnN4AfjxYag91SZlD8tV5V
VQJf/8wJ4zBAWs/VSTgsuVrnOYhklKkpstRKDgHTFgs+u0DNF4Wm6iJllBIrimrV
mVQ9yTwUJrSTYkFtnddfXTX7tQ9Fl369HDqYNifoRZ2Ri4GSH+EWkuqrvUBFzTcw
nwuBFc3mYsRc0FHXoTnKHyCIraom/F4DSLiKpuUKii0OU8e9O4+S+uBHnl9KcZVU
P505sGMrrKkiH7wbajixreiXL3QH4KxUUaLFD3GbLNHffWGnHuO5+D7EmbrpcSHS
K5c81piX8XF0fUqpPzjrnxO2jSLTh+HWLgKW5T8CrgYMe+Q9E1Ua5GN0Zhvxwahv
zlgPeGxDdlGg9T6L7nuaiyFHoM6f3pdXh62SE0sQEC/r87prcaOSD059rs7AWHVR
FJPmWch/KyEcAl/GEwTPH4tJPLICt+ivwIjz7GD43kNgVx/WvZ7cjGAJqzNbYPxW
x9a07SfUhAm7zuRmb5UQZSQc+yd+0LvMe0mAM6uHxxFwH5FLNRahN7yHnEw915rx
i4Lwknl79ChniWQ0zma+61HbYGyhuD/z8aEBlprIk98yezz1HeUALVL2T6DmVAW1
bt97Js74bIhmDE+/VfQp6gFFS/w8c0YMQ76DoCifVgLZRzkt/lHBz49As22tWAo4
8rTIAwwFMKVApRv+WkWS+djoO3NhhQsyUEYy00vc5bKf4S84iW8J0PEAA/SS6M9u
2aHz2hXDHlfUcl0kE40kFNkrA92fXIyy0boYCWrb6ZjtHuuN9FzU3Js5zsVI15Lq
oLohGubhIt90YmykzaEdTS4G8oPDNKyMIF0EPjRsQi5O8orx7J7R5kcg+nj4FIs4
K7sLJVI1e+9K0PnO9csQVlqE7O5/pr4cGQrEqbwU8NGaiVkdLth4lWsk8kHKGtSm
vjkiKCADzblafHeC0A82bRquu1CMhz1EMHUd/BQBTncraLZtXgsrmiRhISzmAFdC
JWy51uuSa5NYLQbradosZwk0+/vtJw+OtfVhfeNTNmfv/vcxZ+KGHpMKYXZaS3lF
rjkfEtJqJHdFL5MeXHutzJ0LSYUC9RcrDbE8kh9HeY6rEicISzRj6dMh5RWptkxx
NE6wM9bX+Op0qXT4Uif5A37yOwpsVDChyqfMwcD6gykYD6f2mMwISe/bCs/1ytJ3
wkRaNWt4ZLNg44CbDsk1hEsxDhdUvVdWfPx+uJOXoEtuTcnUu2k6GsYyd0O4o+OM
NuB6ZxWYQ0v3FjszlQCb0XPs5IbRehE1jFATL2nReUJzxVlXRsZKZIJ03OJwS2G0
nWysaOG/VaVhUwb9qOx0/yxAV+lVkErm22XuiZuQibF0/FdgcqqgICH4NKuYM6Eu
Xr871kD3iVPitNDCy2bhi5oLfYaOLssdmzjClb9fXxSiCVtG8gmVBLU+MHJLB4dX
uamwYcflQ07QZa1eD9mzRXd/3ZKHQCU6hfEJhDzaDkMa/iwQHbt1JViDOLNX7pF/
Vstu0dfPdaKtnRW6wiBCuZZ+ndDVOFGdn4VI9tYhUis5o9aamcbCU6IaFVCwT6yE
Il8mL+XCgaaT145d9FvjK3QQwwTaK6VoduqC7xT2gFwZNuRE6T/nQKsVGKWD0cxD
akm4yVNl7cfUmdbjnekWFCvPnGLaRQi3pBl2Vby8GI/E1p0WlnohGsrPwRFP034P
revzBi9qFxyGmpPyNvx1jhmDbwniUu5utYh/carSGT/cCmEUEoiNWh7ALHIw01uM
X8tEUjIrHYuTYbURRt9bg74HEyGNqZzILII5lOTinKt0bsdwPNUptCTixvcHkx4A
CT9+1KRDLssRQchUronvNv+5fLaPADRvrShQywt+L4JkOS1HU5QqIkIoSggSqZyI
FREalm4IO7lLvH0LEp+g16vf69WHagLQ3fXkcB2MI+7nr4oY1zyp3cEATfbVTRmG
kB7h9bEVtIKpjHpQq9VujqXqC/bvwxV6nedMbq+tPaQ7TBXi2BUG7+40ElqBfUHj
rDw/JEYXVdMR1FZ3UxVvEkVCUvG7P6lntHtIoTwOEVQH9KjLdDYW5bAi2/dogQaV
WwYg4fXcxBwGTN6dCSiuPWV1kherH+irWB2yXbK1CwrmeCbnMi4q0TfVB0Mi76wI
GrNnVzS+4tXYPoqebNlXMJf4pB/+DJNFj3xgoB90Kg4+FDEXV61UhK5qSo6y07uo
/eDqAcHLH1zI6EWZTPZlSyby3KQO85HmsU8dOC8Z7vm4fkJy5f4P8rLdo8dzZFpt
YqJ1rEfPaUCdrnqHJa5Q/vQgWDE8e3krKW9/QuPFEMDlCCXiNaBiP0G0WjRJ9sZx
azptjbwvjKPu98Cos/SdcWApXXFmQZjLSPuHR07g1uqsQgZGqnMie97fU6U2+nd2
oW33oP2Aj0z2K/csLXSMHKipAymIEOy+e96fcvZi8FEJA8BW19kFplqid4PBMHSG
zbvEMgrhOElsOfVM5kpioIVn+G8nqIvNXMJEzkoCnWQrTzmpHCouG13Y+ChtVlTJ
CRLqDNkqJXEJ7Mc0i5sbjauHjjSKiVO/OdT0Hoih8tvAv3n5Qq2eF58EdwoCMeSV
rfGYgrWP0GlaqCG6CL+JoDHl6+s+11c4+kdB+yjSXZ1HyZAzl0Vmi9+0z5LIDdPF
LhDa8eTLtmr9jFLqb5M93zZuhJkxTxfCMBctiPCN5eqrQzVI1VAUcYC0cb7t8tgW
fs+hn3BJwupty4XW1MY23smQzVwZl/96fBQjb1msD/w9/MlPjQlkWxEDRNEAZ7e1
WOckjGeJbf5/IXYbJvawpo16fJun4C+s26oTRghcAyuiLmDoLItZ055tEiZsnHW8
SBpjxzGTTSsjjtjqJqFKdiYA0UkEjblVjMc3E4A8aZFChU/obDsGowoVcxLHeRpM
OPmOsONFZkmipyyDS8JTBoKVMh4UHLbjGy9OeYlOtvKLcDJfezJfvR1mPuJz14wr
eRwW5TRuNSQ7GHFQuZyCl8cgqNYeJ9o4byVFoZHNK8gqqZOP/DUMMf91Gy3A4wFl
0UrTCeNZC69XGlFeYDEz4eDMW4veRUvDFAheVBgOFPHcOAKIiAyRdXLE0zYz7h+w
3rp4V/J/q+3/zHv4//elLKGy42zflkr4XOGTun6/rZY+CwMVOCvB/DbReJ11MepP
5ZhTnh4yPRF8M14ZU2o6HqDadCfcWAcAEsWtSiMLzOtcIH9ETXXl9N60SXYgxHet
t0A8jGMqKq5yDY2AF8cA+7kL9m2GWkSNmuX7wO2BDnLhnV9e9AJWvJMn+YPYkJnC
OJnx9LiXHh6UEEukdO073Pdgj4Zc0QmYHax9oPZcEW71dWd5R18eEyoPof97dHfo
0cIzxOq4no4WdAZ01OQLj/uHMCSza7plI6lN27FgXXJ1LGbLwMUHYu6GBlWeeqCL
PnbWOI6r0+sX/uDkPl9qMSHxlEU4ux+6GbFf69Cd71BB8NTjQdt+1kD0crt/j5mu
twznmPuaFfe3TbPiVLmuRUYpF/Nlxn3dH28pH29tHGVXE5vV4i++y6v+JxeXdZb9
sikAl8ofCgLfSAk2tV9FpNV/euQW0I98Dh//z5uO4IqHpcm4ZV2CvRTlt1zlptYd
a3RhZyWBsp8fkhHp5d13rsZpqs7WfbNygiFg2gdBpPalDw7pYr3So9H+QsWS+aQJ
NNV/sv8kEpRVN5H1o4Bgcf9LgZrUdOigzo3eHdPLXlcgCuSSRrMD6KIXq00mdZgT
N+rd6zGE0VS/SRBTPb4QAsdNdGEbt3Kq5e0+IbUuXt4ECI3guNuiEfMyuuKtt+cq
Ow4tBHJUJGNa8vC+pwEMAmJ2HFyMECLvcqKMXzRyjHo+2qaD/vhtCNQHwTLsFhUF
UCz9kA4MR3+/YlJh1EF6s/rdW0rM26YCuRZPg4MZcBfrtmDVcCAi+LL5kEeAmfd2
`protect END_PROTECTED
