`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WcgaXCjkQ1z/yfXH5bKkJMmDHWofFRFKA/YSFQRPMIxINUrvZZff5U0YEW46vAcs
52IEi0SnksW+4Paun5IC5VA3AxOzJsdGP+0S6vAbLMczXyNWBfDOpeewKECpnEeV
oqrvErS4r7l49jp1rf/XB29bL0AFcvilpihFB3bUd3eiE+rweu4/ErzHDfCpG9Tx
Gu9WLA0aVbw9xaryO7Id5IpEnS3zUPFkI5cKJVjFmefkJk9lBlglweQnvdNNDe25
fty1wCU+sD83HyKc/uVKLUjxfi8oFfs6VXI/30qZTIBZVMFyW6xJt9MeqrZC0rtn
oOyVrVpv2v6uEpG0qQgu+VyIztP07ka8NX8Fhc6fBSC6L5kqfuDx47tkRl7VgBup
xj3kY/HoZs0u4l4VSCzY+XJYlwAeTqb94/pvOHOc9cWbadnFsSRAvav24yz/jfT3
VzFKjT699YP6hZaDrJL4PPzfdpootEK7g0rvvBy7DJPM1CcndrXtMsv+kSXf5W10
deGcWNQ5/LbALgDJbcEcihX/+iPBxMi9qWhIyVjELp7QUHJrD/Ff32YCiFasPSjG
bGFETa53/LgGwL5lFE282RkdQ43l51e25ruDaEzw5LeDCECN7VNhDkzlPLZkalKc
wPLVvHQejwD4A82Xapj1D9VYKqhI2hGYcYuZFGP+OjXUbel0FL5SWBDgjGRFLGbM
aDYCQbxhOtHIVQbNy8FW4TWK+/hTjFi0OHBW2oYdF85ZEDTmH/aHC9UJWREM36F+
Zo+V1kRLfqoGf9TtXdygt0jL3SJF2oCy1vGFHN+KWz+i0Nl2GloQkOX1qE663Jke
D1NqFL4XdGj5FbSxkE2NVtu3tAPy0z1ERKWoOqhC8SDX7uNItVzP+c+Ya+CDTG18
G/E7Ar1F4FHcl4yxuGpyYgRujr398Tr2izkXXFAkI1dsFS+A/JRfXBPHEtWMuUg+
HQ/5irNMgCtVF3xOf9K6uka3+28DcrMu0pvMB/leEgwjTCJnjQudkjbPd+3O/3Qb
uADxvoLjK0nv3Iqpyc3RUVh33/Fcron/QueHFX9ruMsPIyX7LNiZ8n81C0uv3Ps9
5CXZ7sQhjryn8XJMyJ77iu7DdbgTIUj0iQH778+aF/9I2TexcoF8zocJtjQ8Use+
okhuQV4YOs5Kcuoy0hyzd5s+GZ4F6ln2tMoQ38PGUKBSidRDmMnrizUX+PiHJ7Iu
8j65T799LPnC2K+qQNG/Cx4Fd6sPy1QMGzD7I5B7h7JHFHYdLpanRtb0AGAr7qiy
BX3ZytW/8GD/FVzJjMtzSRHdeJpg8f0IU1VMhHqJQMCb9drBcgzV/2xWmn/aUL20
SywIAK1DNm9WSV3rT9SXeSBR69JWRNpqT98NBzlFiJeEo8ji/+RJYcha0QNk5KvE
o0as8PjR2ytX5bNzdbjQs1xhtdrEGj7GJNZoMTUDlMUYfXxwHhTnKbtLQkfphGSe
mLPDEUm1S749CrW3e2tPyJG+HbObRFWvYrIxew4nzYz70oPvBxXpMqyVFhX9uEi6
u35bEgGoXFdE3AoLXHjfkcDplTYpXv7KZ31LMJd503P3zKY3MMu0JT82nbtNOPra
avc0ec9Fy2qXw6HmPNuFdmEAOLuEncP7KneQdn/aeD8IGztBEyDaD9P8DZsZqx93
Uplwc/lFmAYcvJ20k3kDsP1jEZMObopB5y+lWvofV/VtUJCTCDBU7Wanhd3jw6y/
LagkPw7auehwZq3CruV/T2iJ+d6KcO43K09olBzq38s9bo0EdT8b70cSQGERvdYd
5hRuvQMqaisfuSwMuV4LriCLi2E1o2FrbVpKUPKy3XNLltFQzG4W/kvSSQCaqMMj
BL6QyogJQViY2X2EaqYScB60Ek6bMRHlLWFeu+iwcrc0Ow7K7j439cut7IiKvFeE
VBTkKx0s8wYCumXDmFkpLgNq2iVYwFH4ZHYGTud9MhM2wY3NmbGkzzc7OED2Cs55
L/zoxDWwQQu3BhQHtzn0Nes39idtD940kR0MA8W6hF4U7KrAB2r6okrg6mzitaQq
vyfoiwibMl+JI/AX7rnrOi5gjk4DjetfXjjrnWLNLFNsBSW3D48+wWmweopesNK5
REgKPKgx36JGFrR+sD/T/di8La2/f9NMBj7i/hLfXT+XF1IAJ5gNMrHRNIKuO1i3
8oHwfI7OlkSKW5X5bo+qJHojn9MQv3lXIls/COZi2afHmzvZOOeWeIlCerU6X2Hs
T1lti9Cf/HtOWM/75qMX2rBmn4oiR/xJWnityzNmZPq60cJZenEm4uwRfS8o9Gxb
bSPd+FGKNTJ79ebc4hakVIKq7EUISogIZp6tJpU2xVCuLBh+YvDqr9WE1dWgBzVy
SGeSHknJ4sJrQ8GNaoAwDE3pq9xd0W9ZCqSZ0WciWfMAvj/nzwO3JlYRVWj/QKZW
/9gtSWxS9+Dz8E+3VDvcVLD5r80V+4Py1QFG5WEYKmxUVflIuyA9qhRQBzaQ5Bq1
y5b+DQI7HcIXKdwyC+Dh+kNa7iolDo0dpzuxHMRE+tIsi3GrdlIYvfPYGwluvKo+
P5jZvqRX6Sv2iP+3qceq7WwFAbVAsc8YlbjJskH0P9FUzMSh1uRL2IgP0AKgme0Q
DaTqjAKspCpiwz/RJ5OJQagsduZcFmA/wS3/TgPFkWMPqiEP6eGrwXEq2xlt7PkQ
mkjNz9ylGMdHWHD77sqnDwkzqvsCz1I1ODMvdtEHfB3Yj+vX3XROLB1/5Evr2Xwr
kZGbc50tIcfPbUOM3WSCFTORkC8sK07Als45YBsckc9R4s1K72MJEELJcoEx4/3u
yevTIotc2xxJhEOkVkeFFPCJCNgJDGSGjbZx7ldy1Kka9zzKHKtbKjTiTfOq+/a4
MDUgA9FD11GxR58J24WwamM5KiOyZf6LgQyYFiaW2QvpJZdTeRJridCfMVLsZwAG
VlDzaWzv2YHwrEdI4aGyI5/W40avnmdGHTrE8D4QeW4YfOTwHOgV4KN9R54YDWgx
cVVJkIXIZGiTbAyWABNCIf1GGxcruRGyrbiMTmzfKIJixJ/ffpFvIs6F5vSsYNHT
ODEVm1uJxnGlsYReo17VkYTX0pEhIrQWzWBZho2PA9Hz4nZ1T3eij1Vpnv7PjTgM
JRpB45MiyQXq1iMaugITBvjF1GCKX5r2Eji1TIlRl39LIhnySvodUTl22CmgThlU
4TTMTkkb91fHHXbTw7RXYSV3OsPe88sdPTQxSuySOQj76fe/i8ZeOhYrdlmmvEaK
J4FMD3mYhkrmffM6ujloN7gxxQeBLcjf7FWEkTTZhrl/2Z93PfrscK/mA+r8SEeP
trj8uZaiH71Luw42mLFMgLEv+llqj264KbZdXvldwvgQpwiG2IFEsJE+E7kQ4D5C
jbv+wTd1o24Lt0pOCagQ1Sf9bJfsOKcI9vwQNnXHQf8mcMj8U1qqNjPi5MULPLtg
FbH1Aaxt/aeF0A9/rfheMNlrctq8fyCnIGGc2iOnZ+L89YMJKzkOM3mnux2Sez06
Sf1jesP6V7N4CinGO7Nncoh7UKy9xUjIMywOv5ZIhrF0yaTUXCG9NZsbzWy54xCE
Yr4avxNqH1dusz4abfJTEswv8qgbBpFFZgllcUFx460ls1T5Jeizv+c73HWIESzD
Xz+6Mw0OBafeUD8RhwVX0j8lmettLEb8HX5cQqqHdbPLR6fRxwBUw/xSmCLqJ87U
yPI2cH3kMPcn/sCP+xsA9OVd3JYSbDcSQpzvDKKGDWyeSOZiqVVXToZGb+iZLV4q
9D1356cJm3NEXMKOKbFMvUx5LzZYXMFFN3K0D4PSt+/Mf2MSi7inwlZsnw4pRuc/
CJelcFpPjs+ff4lg0s8FNce17Lb51gRF5jaFo4NdaEemk7qxpXn1JHJfF9h48L0e
w2EUQta/MGEtO0qjEESg6ybyMb0H/V/MI1EFJfI1WuoASYtF3RDXmEn9zKPvWKoQ
UyHM2vuYdNTYJ0s/KdLYybZFTEBEEFbLBRyOL3JCCd3cA/OnuCp8k6A+5jDGeRtf
ay/bKfwDD0WZz2n9C8+Lw1igpA9aKEXAaBcTJ+BGayb5oYCiT2MQ9glI1gYeIxol
UM+6l1u5rKwmOX7YHIlPBCtc6nOFpNCO5JeWxDMGZ6xX21jnFDGGNPFvHbN2FUuL
2JdAevoOPDiV5Ik6lZ9vvbQQkMkPkE9S93/9ljgYIn/FtXTu83mJD7rqBjORLEhR
nGRLUiMSsCmNWUp8LJ+qUptdNX4gFtoLeaLLrRl2GBdAmhYb4ha9zYp4kHrZ3Mrj
RvmoSYfLoDt9EyohR5J6wPsO+xozK4zskDPAnVGMwEJlgVCHwLnOxfWgkKJrTy3Q
ixWLV5ZCsVDOFaHEjjQw/TC/W0e9loTIiQzMe8lVGT5L/+BVFUIaQ647LzK3W+mw
t9hAine3GUVeuH+iOEfBe93FKcVxiOaL/b9p4vKriN3SmDCLnMmZ3jS6/F9D7n2e
18GMlh99Irfyq7mhAts71geG16ifbj/L3UgFkTabMGJ2Fy+NDhQ02uI3TUoZnybl
va4F/tTacqeWaY9CYyuHHC/d8RcZGs9db7QM0uyymjSGEshrLxJt86Gn6BVlH60o
qevAPeR+tfDFQy5jUE0dsJ4XXLge2wYyGmcFvJK9vX2UCR8DiTldmqYJHFkXVo0t
fFJRFIcvD5LZ9OERRk4YAHpNBWgHya/0qPL4F78LalHyoTegMMy9ebVpuuucGlaM
WavDjWbymuOTXOfxmw1B+jsdHrCQ8OsAspZpDag7uo8UhR9VP5PiQM+dXgnhEpVC
XhcaQips2U6BuUobTf8mJrA69PX9Bqa09OHF4B1LPkjvpLc0TY9pByHJZjFzrnzq
a6g44catE9VAPIvvT4LVFjAt7nEZcl6bdwJWiqtZp34RUQG2WK6NU5HKly9ViN+0
VFwy/hTzX3qKH1eIxtVvQ0d2c37ph1IdBokKR1tcexcOa8dd8FV6/u7V5OV7YjbB
QV94vWVE/d0H1v+FLOKiYaFD5G+551Tn+fdPrjNyqulGw/5QkGLiIIjV2zKmQEvA
MNdnbTldeUvdx6ybw3FiigxPu5tT1ojJHUOJ1NpQPY/aeaGcp8501NPbuNv7+HzW
DgWkBspOv5IHxpIhw4PbpOUXbg4jt3vnbZU2WR5ygOPXAEbddgB1+FFVrIE6w3aR
kBaxnETeILp9EUd9p9PiAPSyApttnWtHgXzzS05mtg+8zGAD1NI/kO1ts1bNTIoa
XDwqck0TMxBoOhww7nZKYpRA/6opd66NvfSzj3b8SUpc75xc/eKsBguMSHTHexKC
4pgGGPcxODHQfYGoiN3JINwlO/BypfvnfnI/s5ls4kkOPo+RSaE8uitngeNnt7lF
VeRkwMxpo2CYS4g7EcMEIxqDH9Akz8pNQv9Tk/YURuR5Gx8vxkpSvgYl1mev9D/P
FC1w0cZfP33y1ogL9vxtguVjZ3wAqfsukmuxeJi+ht8VzdxRI3Tvd7YScKkhMHfN
1mrpcOjk4QtZpN/f0nW37H4q4knkdfMrf4A2QpjRCuhZlJXZST7+XOFBaLxGlSkH
0S3WWcnpW1+loy+vtBACQrnlSkJsuGeDAuo0WLS2D63tLk7dYfCLZ8ScQX/xAPHe
IbisKuezt318JyZkzqap+dZbxRBDoCbKdTaeOhH49oiQkMrHcLh8IPn9dS9D5GRU
AadKTpbUM3jg2aPBVAB8m3R6YwDa3FttfMKb8AQVebFuNNfGpeGxBtAtIdqIbBAp
+cQ1TXl/klXI/4ycLhMwC8MG2bQZxxfCV1mWAgK4NStUWqdA3/vd25aIIiVhH/6b
cN2M7zDYH8rp8dTxsgkrC/zpnIRmC8uyB7a6mnQbk9KhqvRbvNq30yiPcUEN1dNl
LX9BCUgi07Y6lgfjmeDxqxGrXQnqFXlQ41U0s2I2C7Cw1rJemGEQHYasllnswmVg
qzKiYx9XndPmZo6fNjeVgxKTuVNjRbrANCjh+cBg0GT72Og+hJZcHaNSN9igimVw
Ms1vyDWKiWlKv9pt8d7UMcOLbZdVgJqo3qAkSpWIelrI7BY64hug+SB9eEM6uIcH
pQzVRTRTmu/YxgdgoXwkGpAkGDFn96tNQ461TxBIURbJOdbbxzDtIWUyQfItmbAR
yOYVkBHfjWGLGkMH8GM8n/FNwuZymKlnl8QjfMX/dVRCe1rmm//bf7TFZOb4wSZj
0t4eNfPnarvjAEN1HGaebInLWxQ2c4P4QMPCpFtYDiW1EaQAxHEjSC/G5XJG7ux7
g/qU4aSJNF7QmxWYOLfc++RNgzm/fzCDEz21ESlWebsz5FBJaiMChgKKJZGdfHPz
And+cwo3GLSKNRoLfigBraQfspWOaA1rVoI/AcaEmy1sdk6xpi04OZdANkizl/Dl
79dMA6kDWv8oIGo+N+JR+23XNY8Zq3x31YP1MPgRM6zgI0fMtY2GFI3AjUBZa1Im
n6xp9HFdDHEE9RcyxIPfLc692SaaBn4tQ9hMSnKgTQTRxLqX0m+40kv3V56QgyKd
/iU4hksxleBFOlkAhP2vxPU7F4nhz6IZhKmUR28NQj1mPOGSyzaUDgu/eTkpjqZ8
028ahHYPQWWmJRCS51eA8G5bBNFcaG1gAcNPMKq05vGY6G+PlDpI6HjV15net/rI
2k8AuxFZfoXJkSikv23jfzzl/TXxOKolqMdI7hS2bjDJhdvqqhz+6rEZITaz6jiK
S6zXfbed8yKfybgkXXxoSzBdGc42I3+aySBPnJmG35HW6uHDMhKoGsnKLHlXRV47
QiACfhlcHFMSYrLSE94K3xrChQgSR5hOtqGD31y+K6dLyxHToOnWcjnZjt0krlFG
db/qJwRkZW8aCVpvKY3HOyxnIFKnP2bySdzjGNEpI3YblOZBtzBxhCaQ7D4lwOnL
VlkL51ZUdzxbkIrPFUvf+GuE559FJrM7GW+kfDPhFRvlHlmfX+rYIw1/9L6eFiG+
OBvYMJHbch+HM9fZdRv4FHP/NbocH79ZGIWT33awQARu+gO3MnLbU9YypKSGAMkZ
1SqZyaoULTpF9rzPnmklJ5yN5US0KoHy1S8XOBHpCeAaSwc9hIIlmj8mvyn7E6I8
NwhqVOb4qHPj/0VHcVycqUNPZSLEDaDvCmMYnQHWDvit9va9FqAAd28SmBh42IPM
JO0A+wKH8l9HnJmOfJ+uvc+OMqa48j4QOg1W9u2qbumODAd73Arsxf1lFY7WXUJV
wsIPK1Ko8TxwyUhM257cvQxMMNSbGUCHMcPCOLq7HjOjoxS8ng2jCgQ0wgAIed7I
/+agHClIfZ5g0SsugWQ6tJO8BGxarakhZZxx7kZMj0vB0aQAwMAJNXONXdq7QRy4
W4JF6pkIzs/B1jatdcohVUwxPc9Aoyp/bwTY7p8iuPLZsGbbJ4ZjKrgal+7eJGhZ
7wLKnWCBoPL2fEatt2i3nlApmFDmSyzZlGp0e68tXtkNbb94hOuwpZknf1l8IlGm
iGkVWnWeP934zsEPiJGUIWXQZ93lvvZyjmwLuRCuRa73LJq+PqvdudWmV9AgH1Z4
QCq6mM9irZWoNoO/w6zUJbUcfLPk+90HUyFAXtKUJ6lgEh9D1OCXStVWf0SNlHLk
6xcTREmLbzXgJwG4ocopy9fOy4RSXaAU+4jKpZumkjV0EgUEDq/Xwsm7+pNYOiwN
Wpd9YBU9m8izj22GVmNU7OC+RuuUKhyBC1hheyyteLVdbWztv2UN89a7CgSaBYq2
lga2pLBY1SIU5HQnVSDyNkqoFxYoBagTZTxXkYyZ+5PSAFtXFRFUsIsSKMd2bgfz
WMN4tQHoYLZHVtmWsN3cKbAhT1xirRAaR5+re7Wt+83pvy2irtlGg1LkigGSP8i+
twwB9X74pT+DNzlAu4nquulNprfPKyTRpUnFkdiYp/q1lL2khpPnVrtdtZCLe7Ow
DJx91C1Dnkuks9srcipFoOwy5hB9pji6c3ud11obiOUomFnCAaVcgGqeFeSBpvXW
utmw1/zdu+JFic4wnaHIrGxl3fDEicp3Fr1jdYANds5FvuAwgYta11JiO6Ua7l6F
hgfAOyUtGKrD0qpVzi9eT1g5r7EvP78yQAEHq/31PbflWAkcS8jNb/OyMOsYVTFE
y4KqR1tMj7l9uvCTzkCZD50F9xBESr+rlw5GGm//V1n+u8pgnYLsGQ9lEbX0/nqp
qV4PZgwBuH26zc8KE0jGB1WLajJ/hpxe9OqZry9GNnP/ZDCc73SzKS0d9ywARhMI
+fWEse7qZ2MCdJxtQyKRdHczGqhXYYQWM/6n3Fhl7x75yhIcVPjbd3SUIb5DTKMi
ftRGCFL+WfIvyKYfyMaE1a+GHoJJQaHyff3tVpuTUdsTj8ajFTz2ZmaSVkLbF8rf
9iiB6NxlV8Lp8AjcVOY2ZdosVPEySyU2w03lgTfMfbUJNPK4L8Y1MA/QoxM7TRNd
CjGBOQCQPCeJNfckyn5fypkfZE2mII03JMXZpEt6TDj2pDGreSjr/tk/FX/MthVl
TSLW3hF29AKSuVxAot6i+rD+dWu6+Y2lsuh+VCRcoGXuTfsMAIxSc8uKIxcBTwxn
ogNijiaT+El5z9mmFb+xcp+fmg4XSNUqzA+WCDFPOmFIRWLKW6glaCo+SZz8+ggX
dhZuQpOj2qvr/j0y8yLQhkTl7HLBUXXv+WMnaiAM73RJVHKxg4MBSTrpDlBJaBz8
dedm860kc6qON8O1gUeS9m9GmUYEnUB4iYiHZTFlNJYQRMiNHvLtI++9Ksgzz3tY
B63BfZGU6xYg0yXN9fJGq20bfBjRjd0SzJvo/I4QPb7/EXWuYjbMFu6wUD5X/EuL
eC1St4VWV/+q37x8Fe9hk3CEXU57dWvAFetLIDSF25eai3Iv0gBFbZrVgg8LakkQ
ASqNHpfYqGLd2pQ6OqvjZlcvKHanJ6P+x6cjWr77VWgq+lEptrRJTLLrZpDhqVF4
M9oSrfaVlphQ3Vqmy2NVtKaNi4ndvdgDISYlEmi96DyUKgmlQj+bWWxZ8L3LiGLn
jL8q3B6bLJrOnPPWm0hWLJ2fcWjTNfOyVgkbwmaxH5R8SbbFHEz7i5+Oxa8nI598
21UXwUpauo0o46RN8zo+Ju1CB/kCA5se1nzyZyKaoMxklWplVwwIPDIbPHbR8mbP
KuEoDE3b3IIa17drQgNJM6U2nWp6yXMljvz73kHtfFxn9mVhZq+onSzx9niQ3KmL
glrQhtPNNqxIUj0ft0U78fULM/TddvI9koVAlMRFr0Gfrjg02+SZc7RBIht+NaL4
C242ni6JDqomkSVBJ4j9wrnlUY9tQFOgIpPAsAu9C5WSCg3q4u66FUswTSg/BvXy
dWCWkVOyqDutwuzfAplaVjJ8iL6GS+fyrgGt1kRjgaUix6+riNOlcr15xgttI2AN
hMKG8x920hRzVs2wJyUp/TwUq7N3Jtb5n0iJmGi0ToxEz6YT1TnaO21eaJdqXlsG
hLha5qZMU5gaNreJUGF+Gto1dN68oVAyoZiJE/64w0SypWpJkx4ZAd6RpwaNRqL9
kh+vthcwAoVvIXZFlO7vhxTJQ1SXI+nYIDhtL5iFTFiJH4gaQ8ClqztkB7MrO6L9
TW7zu+MemKWWpRh+bG2GCAgWJkZ9Ei6c+qmCkYBg0MLka+EdQTZm92/BjxRsVqTe
TyAf6VNRsrqqe67gk3lmgaIbg28ySZYxxPMtevrBoD+nA/9lcVWznUleJ6UyRwZe
4if+x/FPRPJ96NDEhpEKqbvRI78Zm9Xb4y9lyruKd+/G98Vnf7ecTyom4aiF3m5w
IS5mPH00kc7Y1aiDlgvbCn59aSBLQ6HW+Q8YFHeokCJWqiulb1AKSltLT3rtdlvE
EJU2qICCe/CXWnZ7x+Qh9YXs/h+KOGGpldP6UwlI5MQ5ob2Awvv87O9ibeCxC9QZ
SjIWbwThfGW5gcNFnC2Z6rZTQ+/vbk6mPCftQJ7sR/VXlsZbNGOA8dZIUqpORTxH
jaSIgVq26/W2DGDpGH6mEQLxQYHWkst2EKXDZnq3QuFykITG+r0i76iu27xWCdxH
oZ2MMpw34wDLj3JLfNZQaFXR1uObBWGloe9qrITMAC3pOAL92c7QrcFsEbIz8Mqa
j2kxAPXn9PUen9ZM7S3VuVkV3SDzZ1d0+h2mUmxKIRyz1Ly3ydMODKm4PJ/CiRwF
t4o4QCzAM4qnydTdh8bvfR9NjA4F5LjmeiHMy7kuuB0Y9GuQ7SF1ZDTjm/9PSSD/
iRxcQ0YFu22KzLEWi9gKVb4XfKYuFVbQPgGNkyoi2BfT0iWosqo1UgJSrJW88SiH
NN+ZG8QbiC1coya/+RS91LOo24rqfj9fbetYjIEEBDT8BhAFq5uJ9mEV8EhPFigN
epPc1uWwvp8uXzhEzDyHinJQpQl4moydppFKiDX2iPAjiuVFU1wHpEMVqnyOsw6V
9lR0oV1sYHwWj68CfltLu9LWzpSWMWmWjqi3toSD3N+TD9Ynp0Vtueu0v1dr9JN5
WvvSTCv4zPzL7PFYyyXO2hACbmaIPIP7CtVtbLO21wEDHWN92hNa0LKmlLEaeeuv
D8ypUFp2M0Sed65BbgN435CFXobxtvat3Q7RhC45cBUCGl+qGUFNy+q4ZqKznRpJ
2Nmaz8LCnBu306ZpP/HQYebesTLk77pBKX6Ps85G21LoDMiwup1T861BTBZMXJNM
VWiUlHxn2oeJcWdtg48TNxcnXqucCb8CfFjdv1hGvGzOHSyz7mc8NSDIU3H+dzzg
Gllf7n15koWCQHk+ROUTKkY2ajAJ35ex56dmGTrcrDTpswlNoY1ikJ2Byq7nXKJ+
//0e4Amu+uYx5h8rPVKp2/RrhJHZnbaIhcSZqeMuHPpaDBUR7YCF4/ofOP1RlwW8
YDng3WNTvQD9xeA+hbZqHmmzvfbFkI7JNVBVJAdRYPIBNamMTIALDHwUaJQWjZLH
bKLQbZwSIJtkgaRmC9k2OVi08daDb4Kx4bjgMi8Q1A1WMY7JP8y2gMQcnKbcCv1J
0un7VklCYg6fEkzKhdFDQBUHtGwfEGbwcDwyLlA7bA0Y1BGj1BuKgy5rlLFSeXQs
J7mE2X31GNevyyh139yHdtzkxMyCc9FtkKXokv9v1XymXKM5mkHpmUX/EV6p9fqM
RBS/xeNcqPhRA/SJ2uoBZI0u3iRPWM8oNL/gcpuKLOPAIaAs7R6eZgAevXPkJ0cj
f057wGRR1aGrEwXyFgEhVILLvQTxfrVRwZVi4Mga9flJypJeOyzYzSvjSp6SDua+
fBdxcOtQ/ohCLYNzDXzV5AmXmSlK2oPbUFUA7RgqLtgQtrL8RZrlLajtc6+2Cuiq
9FGFDIL5yLr7VjnAEWOY1JE7UmjqRCP2e4sbBS1cU0GmnfnyXmKAuOV+8VfAnuCs
CcN8gv4iwSr/uIQeo3TKAnl/msp8ZpQYSwBQr1SPG8m7ogUnaRwPpwsPondvkx1P
WmJPQSdototw+JS0xS6L/O/gKM7B4DocSl+SQ4iTIfY87bj9xLwAczEdNeiQSw8k
Tqu2jlCkQ5lw8ymoy7o5DaWSJw3Pmt5ojNu6oFn5gfic5C4qQJkD64ZSWpdmMo7R
0fBH8FUoqpYDWvgUUTD794BJ8NrCk5aLR4qzR7x4l9gSS5Usbn1RFTzwzMYIKFds
kt7nBJxXyFbS/s+NDAKojkv03voc/RssDI8wOgdheTF6Dz/385eeBIk11LmOmp2k
alE/e8Lxi4tb1yfGczkrb0HsPwkMDj0x9TkE6ktKUDPs3KVDSz39e4tesnwSlIyY
DmTfA8pAq2ciX6agZJVBZryOlPRi9K//HrTJ0Vzk8HOmM+WxpkK4k4Td3IF3osCM
ZzP3BxHK2M7oYMH54mLr2LTJFwtgLCWCI5IOCrlwjiucq1ycBX7ged9BTEQDlmhq
1eVzpyNSS3wob5sXiCNewlU5eUD+X77elIwIR9Jaan8MjGz3u5eplKhSkJqZQT52
4D7G9iyXXEdzvKO1hwzp+V6fyKXSuThzPLmyhM0gCskbWw6ji6fKl+mMHFH+RKvi
RoXllaAY4CSmuRY1rbaVvfyvl8ozfO8NpDlBl3vNHjEW62ec61WWpxjG7tNGHPrL
QJUzOvpwdUSeg2Z6vNEMxSlj5m9K/MeFgGEetJudLaXmMknJDnfigbaPDsRGlTMW
bryW6icwRRrFJdhjSovgJ0xvIohiszdK9StX2nzVSyuVNXT1RYIwucQJVdOre9Ep
teyjWE+Caiw631Q0ZvkEbnfb3AjjGoDFJu3m0EhpSmsasakBufT+0slyL3vajkj3
jjFa6DXL9m8dhdWNDqCYC0AraE1SJ+iBeGWVnKGBSTKKB62OnQTDO3EowhzgwwfG
Y9ccd5peWnzbJy4l+YHIrYnN6P8XZsu/mDO1C+d5ZbowqwBRLrbS7N2s/AK8sDw1
U6dPqSrG8G1I8bfmzpetTQDGt4Q1R8yG1OtpZCaR2tysRGgUTOWPE53Fu4WkM8Wk
F6PX6VZKzG78GDEazNoKOEgZzC+CboPdh8g5hSQ22dqfg3aXTffSVGMYDp6r4j+l
D4SlnvGLd89F92ZgwPOmH98e3K753IfhkTBSYWkuUNCrXNEqxNS5fQRBfojb5gE2
CdoGa2iBBWosaDguREidW4VOv8ZGGDj+TDaOjfYXJXhCUwOzJZ5LXzbYiUyCYFRM
evq3U3+s7X+k+eo6W/YPF+suQETtfRf+F3Rhs+HdiRxeJGaXAVaWALX+aWn/ttfX
PON7REGboVg+4fgPByKNl9aBnxKCl1/Jmur/nFKpRrHdYKZ6cVueLgf9s9tZpNCQ
AMete3B8whDYu0yeWip6DWkGEz07rcvswhcVpd8FyYPUbx7SrP2n9CvYh5NYqqAL
NLcuhDj7ytMlwHjqs+y5pd6A3jilXBCIv4X0/oh9xQLBrKVLQLcD+yROe3jt2LXR
UAExyrtU4PVVwcDYJieoGY542lJwDq5Xf4Ddc2ieF//zggjbklDwVAO+QwjjzLua
jaFyhjxDsayJW974bmCeesxvf+58HdHHL+Gqm0SuoKqCOQC6WAcT8BSr63SmyGzw
9f8Z8iRHXsCXuCCLgg7irhlIFyu8YY94AgvCOswIXSYK3R5A/+0gn0wssIiOObh0
oUt7sf3SC7+jkk4G/O13SpLHUz8gvFdscSboGn5tWehNTfKCOTTLN2wiWCgbHd7r
jh6tFZxRweg4Nn+bqsvWPazHjkCt72StQwUHVHl30HPUub/QgmKFNDVa4ks+pkAs
vIYnUlBI+pnFsNJTfKDT/CJ94rbmSx2XqKFRhr+BJqeP7Kh3+Izpmo1x82HGRjj7
vHmqQRDC0F9IayK+F9E27NaLSvfpKR73hvK3kHmIzLwL91wb3b8LUgXOABvOxCc9
Xevp9wgk7TQAaIjfLjqn/ucNubgyT3CvhThesM6ty4I3ME+Cqdi2J527ILhvrg2P
qkgyWslkLUlVWzwBmxkwFRE2GLbll3Ar+Tj/mkmiRuATPau8iw1dXSyuMeg41uZl
bvPvIlnq8kekZd8eYwinfOEHCbJVISzDVoKIJlovMwgQXwOLbyJ1dcPmv57h/nwV
nt8gwRazBAtgeo2+Jdb0Gfolnk8MTGEKz1TdCygCcq1i/5K72w1GHIz3HU0/4tQ+
UNUgdmc/t6WxRTQ3uCRAroGb1OpXndopQHtegVdWDH0W5JaGw/bf+DM8YXKN97Yc
jBraDnQeqFxM6PJq6mPZUXLcNcz9HlzRkVEmnGb5KuboHeg5rrDK4T5L8q6HjR9r
rsYqkW5237krQKc+djvrjoHWNx/kCA0f8/nH0WhYHqKsckJM6BsU4pJ9OsfDFjXJ
E8/pQYDJLJ2YlJSmEFCA7i3oJwQvzkEBnd3tKHFtyrCimE2qkcafkSWaKWJDt+cz
woRgoHwK4vlZdqhpIL3xGaJdixVQ5/KbAUbVUTsDiS3BMPcgZ0QM5jRp81sm7IrP
aAwhMvAl3/4iC4xBbdFzmkdiXcdkw1OcBFicNgFG398Vxn4eneQtiC+uqcacXI5Z
gldPA3evJ6yuV10oNKsfO8X4YH7SwjG9X2TmvNik4xcP9oH+K471zYkOaV0D9a17
b0u0bVI3k2ySDJIHAMMNevCmVhZsU84eVkH6H2Mf6doVip2L1UUFTd9hDmJCLcXf
Q4eT9boxZq5/TjRwqKD9+XxcjRvaEcUlYO0Lgf28jd3KfbVwGIFxUsEO9Ga/lfG9
0laQoMlzFevwUjaqqQHnMYdxv9VRc/ntMRuoK0O8UGEbkfxfuEy/e5vkIcLvA2Ob
tfkcT3gngZnn+kYDb6lS/vDUuqHna6/6+qZTya4CvGD/3GA4gtiiE1mAe05bt2tu
TFETGFdN5MkhP+EzPJMq9wrfs/FNyRSrhZQwNe/nxI7oB9WQFBsvmq9sRdUPdPbU
MH66ztoGewPAeZXrm0c69z48aw97+xI2str0qErhMoMtD/7pOm89oBomSbuN3Zue
tiKkHvZxpoeWEjqgTvNcDbTHd+QctjI9kcj0dwnMo3dFfudIFR6BVAnAxEAW/MkX
slYakRbob+zwjjY6P88gdEEc8vfx3VKm3STW9cvOuvtinmIavWFUnW2BIHakH5bb
91oF2DskqCIfQA1ufk++PjJbd3Q4CI6cBVA+KH8AYqkKc1J5KQd+TiTpHzdbd/2c
I4E7pAD1tB/GziFy7nCDK0BjDtOxMrMtreOn4r54u/QO6sDJWxReLlMaP7qzN/XL
6F+1ywEWChsya4y8F+sLLmnDmrkLHEcrtpQqRpe+a+iUpz0OyrL33kBnb7kScnRu
81qpx4zvMKmeMH3p2ryOl3vgayZsb16m8qHwy/5Qkr5eEmcdUfNyglwCgqTeqHok
z2hGWRh10cw8fiMh6iea10z/p9HqJoR52oOSaLle1hAn9MjbZ0qdQHo4geEevueL
smGMC+7tCZuzD4epjaJJln/OOkBVsrlnydkLulRSm85T268OGoomyEH0tRklEAlr
gtuHiKhwl5Z6YB6UmBVEpkTNHiuu0fuIMFlWdaA7DgV2yB/ga3VQEdawDHlB7rw7
uSqKvWHnVPJmu4xVDik8WM30MVvK34bMqysZRUwM23efrxsqbPdV7jwxyELHcjFR
64JW7dJ/sKsg8pT5pE7wFNH4pHnx+81oLpCbw/88HzKKVCeXO0zFoNhl2TgHSfuC
0AlmQycdgxHe2trKiA285DVe+gocTkiTRO+BoIXw7im+rz84G8+wfrorpyrWi3hw
Tqr5SakSljE4Qnq+xohw8wajBsB5jCccLG3GgFiX+MUIvPTcZzvg6SyCDucGPSBE
GcEeWgF2Bz8drXCC+TxQTqnFctZHPTK/sHfcysenxyfcMZjwC0gqtHta6JL/cSoK
Vim1NSdTAePW7Ms58KA3hUlwGCtAgLx0UiVZo5CIXNP6YKYZ4bUBXVBBRo6+vh6l
YVPq3CCJ9lnbgx0YP/sfICSnXTyUQE0mddQvWgNJD1Y7bBQrO/LgUiswQ37TsCZI
v7j15b19p8MgdWu6yt2TRKrs8W0PIIC9+5s5sfY34Y33HAs9rasMUx+u7WGTDhko
H+G5uoSKOmbbpAzfI9MGiCdz6ZSreTkOoAAncxhMcZvfLteF6VhcbQSnM6NEgqiD
ZAGsoWl10zcwAOX5JxJoyLcQA3wF8/Rle2M/+NzbWKlNscjPtzfzXRyPA7l2ohjI
sjzBKYQkRhng3Q/cv2HTPaWb9puBqVmOuOL56dC2uYgQrpvVqc/4thx0G33oGHG0
BO36SY+jpj2hnZVtKCt2bp0u41WZzbqNq1L76KVh0XKGCjmZIH22BwaJfLujaBHf
NErn6RXkyd4t8J62xkmyQMJo9g8g8Wqidyfh+UR9Xl9PYhVpoTpUJCWYPsn3hmIL
LZq/A2z29JBuuTjuy6xiB4P2ZkDngz+A/SvA/h00aczxvch3v8NVmOZDqR6N087R
mviPJBWkgXJ/DkTzCTSwdKfdo/UZ/BOXRUX2F9mLGyCr1L6Q3btvh133vY9fKaSr
3zVn+SMscSUzqR7k/BADeFBVdtaD0hieHhXSgABi+2JC4XYkY+h5kiocykm6hFbb
0mEn6rbwcEGYd6hjQ5SkdtoFKJRIz8wEzlDDv0gIUX4dytX7I4p+S8VAv8YS4DT3
2NCcw+aeR/tLhLwQkQmt8hRnVrgbsHqsi3+tBw/3lCrvSDtRH9oe2jtZfpGZSNxl
oDesXQIfn4TS1HRPy+HOWxHc04Z9XxK6nfBFKn/3Q0faiLpAbNqshOzDB8IKG4DF
nObsdPz+QEjZ601+4k/rKagJyO5OYVnjhG2SQmZTkBNox8iS45czlyLIcqVYznaT
h98uLq3RIMdqFghgiF+VmzbYR8HFG69doNJBfm4GSAG305+X52p3rXmgAYgckLx7
XBvFsq6bdjxXo7JnLp8/5dTjc++xya5lIT5MynIqLEJPkVZydFsrLssYkvXF/F9s
N0ygvRj3zLl2enxVbiPeIJDMoR3Da5abnaYHS2gWrFSPpDhzDpFuQ3dwx7Vbdx6e
q/pUeoBZ7KRMeAg1xMTvY3r7iDnpayEp4uANnHNT1mKjsuQ1zWODZzZarsKi8+Dk
1ibLyFCTs5CR3nF9IfT5IUShwBoxObNmxv/49aCat4GZizChZ/7hMt+KnDpUkYN3
U6HAtuNO9Lfuyhiq6AMOPLEUtBDQqLAmcgg1elvx+A2zGMTFWXUwYKCIkaMevVOI
MN6LjpvirAIV3a8+AX+1a1cIBLOZEGIfC60cZ8Dc0/jy2KmNPuIED/MsuPxmfoJl
pvLfQCKzIAm/IDTbukColy/3Xuc9J3cozT6rNgO4TkfL2bfho8tereEFDcoZoVNR
s+Z+rpxjPNR8Sr4Dmud3me7QnZi6U91o67rFfCdsK96Ixd4IS8WkEKif6eXluZQJ
eEP+hyL07qeyqmul8r9XbEbFDmD31cEj/56LJCnoeVK1zuvVhqEhdRndIC8tBMan
vM5Tu5nsypjm7PBDdzklfzl9pLBHqPAcsBQmvHoM1et4ejyBwDDFGGwQuU04oybR
lLT9beQCtY+On5g7gNhZhuKcakSYCO3ef36UPIF9oYcmYlqjseNwW/ro/j1oSOM+
0DWZZF74T/gJHJqUEd3nQck60IEaLCai5N82viiyCDPHX7mOgUa/74DOzGs6mvL4
1FcR6UAmaVsjkBtIu2NmrWz81TRo0SjhB1ZqvcGRrBUA/PfBa0PxcmB/ZHaQO/Zh
meFC2uRfbgpfE4mC+pMi0MGGMQ2eJgUU6kHc8czN9qL5ninUEYSFKeQEx1cTVmZt
Oz/f/zwNT9iRpGdCMC3oa5nOWun+eyGyVyskQY19V4eRebz8yBzSYgt6OCI8tpU2
Gj2HtgoUDBF9x+7gfa1SCRSJv8FsHeHPXNGnFuFxoWjdKoa549BnSX5umkDQ31Fk
EcCuVa8c7CkN3USq2a1uOoG2iiWrku/kJ5aFGi/ULaQN+ABGM5ksAMGHrZgnFF0p
V9PrPwC+U8Qepl8sXA4ecxeDIn6ay5nuiszf0Gek2sTmOKGm1RH17MRMCVrvvbly
34giJ6QDah/6DKI9OIN+Jhtrnb74JqwrgvdO0V9OMUFb0lrIqCDfXro+x7jlR5tk
09I3lYcm5ht/+fdxE6hE5pH5dTGDwO4cwGpWzdhH2EJWPZS4XN1hsuw96+3wNB6A
mfNTGAAbQNXhy4lZeS3segZrGOjhxozjqQMtZ1+a38eWuZpGRiFqAQLRQKbMMrps
8SA9I4eReXTBJ6ANTZNefjrwEaCxkrMRw2KckOHQi6MyqkEX9/byetMsspYNXyDt
hemLl9BPDkH9jOwMeXwuzb5bz7ohF1kcD5NC8XYBXGGNMZfarHIZK/JydF4Rbjye
MAIT7Hvf+0EWrAY2Nzmq735020+mOzjrA3hWeOQD9xMrX5ZuLHLYHzWLBuc9ndD2
E7W7Ryf29cO/RuWfsINzN1E3+zOOc1EvY1owo85jUm24Fn42xuUeV1ywGD8oHqW3
e9ZOKMR0jvEU956c8kGQezCUV4zcqlCmt/CsRu+YiEcTcLPIZIJ82bngQbO86bKI
o0vvou+FxWFVpSJ84Wn/CpF5BhYT7IDTzuGjeP5ZOxtrcG9fD2raj5o7g4K1Air6
Bjf2vVKizM3mS7V6GvKg1ltXloCOTAj5rKaLBpWoI8Pbx41YvAmHX3yP7KKSNxHZ
bkZXW0w9OuNneL3jaTyrhcmOTD05TDj3nNtGdBq2tkqi8810qXnxhUT58IsLCcXU
tfiItZr1PjtzVKWgWU7ZlCCeqa1LONN0B/O8EnHN20KJ+MYTaqGR+IHluP0XLQI3
aGF6e432j7Sn8ZCudYYqobAr0GGmkto3nuX+I6srKxfiL0TTjqkefXE9yz0PQmKG
q9sp8YmjuUlrX3/BW4TjS3AQAr4ufX7qSqIJnsu/CxF224KNIuzZnrIcFJpo0hly
F7paVx3Y5rGALshmc0fsMAgSNoX3awDlypscww+GaJ36asW6Xj+Dqz67lR474iHa
YYFMJgpVvmU3YDJDOVgj5DO6TZVIkvJhbo+0IRYMlsVdHUFayxiRJOIWwL76yKbt
O/vVDmCDaQECLrJFGZZytJUW581d3XmwumihcCu+DjNtrzxNGX/Q1PuFmFgrE7jA
1O9ewNTS7SUlTFIjy6ZjI2WOZwfJMjavofQtYRCGW2Kk3l07c9zKuvykzviCGJVP
N+OAK+zeDpCPxionF3xIWhjTGiyNL5uSE7XE+c67e9LfHfTe1qHQvqcOLe12DYET
bAqrGNZrb/GlG8YflyrdyE4FfiTM2G/gryfjDWA446/02+5/yJFub+5Y39GkZeEQ
HwVWIsRDphPmtwNsLhrNKhT9Ltjn9JLBT+QwVaOigUeSm5jr2E0Gyr5quoGEvloL
Le7dYy1GExIeFhInAx7uj/HYr4cS1PrsZnUoSLDP1nIqYiFaNzr91KNlGSeo0yql
89PJAHSmV2GO0g2yAZYzt0qgt44SsM7tx0ILrV0Sw0lXUH9IdGj1rPd7Yd+ak2kY
G7n+CfGDfkmc8+Rbs65slKPqnpXAA2zG53oWwXr7+W62g2V9MmsO2Aa5qe5+pO+5
faVXpoxP6X4lS2v9CR5kb/ueFIf0Uj8CsPCYM61g9wWGloYCkRzuzb/n2/dRKorj
Hhw9WQZ7AkNMJfLPBEqpYv0kcTaY7CCPq7Jm4pP5m0nEj7uMmsw5bclI5USSYabg
6j5hEkZdttc92bHgUe5U/+K6ix7ngXwXWjSV/SgMdtdJovPpb/7pktBGgpBeuRtG
l7Qi9knuo8j2HIZFjTXZVmfAIie8KY4Np48HgyE+kusv1qX9+WXr8RmBU7H5QEhF
GBdzGCzL+tyE/My2uQq88YpG9kbAkxL8IWeay39RmeDjv8oP+zNIIBzZzYHGX6ML
7KNegQn7PiojFn57yuNQx7bvSJqZj8jX/zMa2slLhd7qb85w5D2njfjZTm3nXhes
iZhWFXvq9VQDAR2zgJXZbzE9YThbfg7+klOweM6q8fdY8v+O4iznfYEbr4o0+T/E
73SkBC4U2JJlZExOYDPj1YsTzSEWpKek7LxorWiiC7agNT1RrfYVd/ZbMMgV745c
fE5fra6QFZVblV0krIbyFyx0K9j5Sx+AGk4JWfFoX4ij4Y5jy2e+/zjtT4er09G5
h64aJItWtrMglbF9DqFKuFaSlkpvANfDllWpr+kpGQBbKofp75wOGLa3WrzCYkNq
NkDnLPAZTi1CTsIbtrJhgdXnqvS3HkdnAHWN1EppHkdU/OZUkThidYi5NokO0Uyo
E5LmSEU5j9i/M/xf0c7lxsLKDgQqrVyrIM5onerOBb82eVtC6VG6DLESj3i0EO6J
4heWUvnmfmw2vkS3G93CIX/2q3vpbcrdJpdvwE6wwKlSagM5tjp7cMXmkRQj7Ftv
HWZdxz+BGlJco9MG3qJISh5qUndS2BuvA1cFMevqurd0P9rra1Js14TGG0kDZ6po
jKwJ+bmIE9SzxsSU7YuY065hO6bRAB9BBG9QCfMX/NJVrez2vdjfY7r58OMZwmzb
M3n1I/WpoNcfTa7Fd733hi289cbNHxiZtI78koUa3iqTJdNQATLuh84w/ZvuFwLP
aeMgC4oFcU+6JprYJyrwF0c+yo3ogG5gYGXiHXz9lI+4cdoBr9Ep/PiXzdAf/frP
O2BhSz9CnzYXHqR+ICLvre2WtgY/FRxyqcz7MfxkFLIyeNh8nuvDsktBuZ6tznro
OiqFDbvD3Vm3EyQwpHwbjypGD7t/yOyT8oLrm05WFpv7/rsxQ41XclIadXK/UBf5
XkBjj8oBpszqQO4FeHO/h54YtarpNs7SPvmii6xFladTzHxvghBJkcUBvTGMQp/l
VzPHa7mPfRTyHDvd0tU869VVb8S+z/6wbxiV7HCSEEILpKiVZeWtUj/yAh5CWBEs
o3zIzaggwXw1J2VYHlExkq3EMMQS5UaV5FL6OGHvrrPxeav+YVbDZex/8lYrNhy3
Wt5fNFbH7PfMR7mEET4/bCWvBgEfAE0VzMR45hTqrKqSHB2HylRvF3ParmiGwJGt
0beCJSQwUhERy9k/0E/H6/Hwl8k7/6aRBgwbVaewA0iS6+gWjIyTIfTK2lhtmwXw
q7A8XwwkpiiGkFWwgKxjU3VvUtm23hyAa5poxncmJ86bXCjzp5/YIB/UHk4OGGkI
GmziTWC8RbDSssdt3+1DDm8ldu0sOyXB2+Hk32lY19weu2jNmauSW/orWC1fFkd6
iBEhORFXc0TAM5qLSdn+eimVd5bQwkUZDTc2erME7+FVghnU3zpuagqgstsRQXpU
NUimwKAoSv9WJW/LAC7f5BNl5SuOw1XHGhZctkqUYEtGvPaXjM/Jic1XTfub7bab
CmAZIhigJiaRKVrhG3ch1zWqlX5UM8BFCuIeqb8KIj33Dj39nMqUkt04sUMfDtU9
Sfw7A0mqWXnzl2an4GDH0e98Xazu2hiKfd0rX6+BT07JV9EM9oorzcuCyuDEh1Sc
UXZPaAE5pE2JLRClgEfcrmT8dYHjwsMSY0nsbNB50gLtHnfwiVUlNquLUngBRAnJ
ESjDzjRkA5PiHWqvcHhC5VeXt06kzb/koP3eRc4GZRHIlTSbZMDsvZx0/X9wpV4Y
3TydS+IdlIatgcvXMcufX/O5DDUmduyXOim3NhgutPZvoxBudTPkqMFM4O0oy+AN
551Tnwi6qT/2WkW7uBeoB4DrVR1Mf0pqGSDtCLpzMWYKCNfhwuzgcRvytYrYINvA
TrrFEf2EavL+ZBsHm/ctQiVBiRoVW69v8bc6M5qNUYhvp7RoZCgsVjdtCXeCLLL3
ettp7k4I1zbHLGHD5m6Rway93WVRj+xzEji5VdEACYOfCWonUd4FotlRrWWxtKm4
ig1BFFru72Mr/f2lcYWZfm74CePIm8WPsQzoJuMgK1VMFv8ohjyBPBlwxRHadcNB
+3gPfsrt3Mmj3c5gp4C6axXeNzIXMsYDCXa9h/J07JAbyLwOsFnuX5T8l1zKkCmN
HlS7HVdljQ7nEoam+6e9NlhH+rQsUMbKLLy2vS2hyJzVV1J4lc/DyMUfR6XQQdis
bDWLqSx9bDOhS/MCOqHcZeXj/SeGwgkXm/AwqCw/ndtRFTgjhGFRzmU33S0/8xXr
lO8hdsiWsMB7LxfTlhSbEtLH6h4PpXqXJz089yAmV6vl4KUoSVwfAMaXzxNVC6/3
eunsdioe8u+zQ2d3jI3DR+g86xoIG1CvtpE6dDuOkmpcvfChSkXIVh+PR4uWQEoj
fyxc1qXNJ6LX+dpsENgJwMgJLIjqFJR2nQdS0NW4e3OayH438ZkT3pB6lH4SsOBH
I4usIifB+QLVtc67t2at8Da2oN7GXa4wmTWX6UmFl3uGsCkJG1MV4WeOM8SqZV+T
ZF1vZh6ipTS0brI4lC26kiNbw6yXI+Hv4qmcwCs5F0/NoaLpATvl+x4AYsycAtT2
SgvBJe0Ndy6aH+pveTu5RrbIlq2marykK2H5AYuI6uRUyGpyXHlqxKeGlwp0u/vc
MbC2yq8LrBp0NztdxaI3a83qGIWfKnjNnmzmaDCEg1J+nsksTMtEPDc+g83h8rRm
w90PBugoE/Ixwr9uH+SNbIXMHiKr6Y8jL4rLBBSwTIIi9TJmteRGrd2ohzZ06w3n
x2IRSdX4ljRnGOH5CjN/xaD7nCBg3PZO+oVxo3N7upiqiXg/gMn8MkYdvIqPp9td
2oP1Gp5tqzUqLWxkYzHxAOK34uDsxZxc27qAIUq/s/nX0WMKQCPJCi6Uf4+1V5bt
Aujx3gmot6MN9hqBDo6mMQhiHAgOKaeV6klKvCDTjFLQdZNRyGJjYbpOxPoJNjRU
GZIjip1RLfG5+sAKWA0qy/hpxN0uFl+RwyCjgVhNVDnf6XhrvDeVRoA9+4uDFRJ2
OWYynuOCdIAbFdID856lKkEKPTRLwk10CaZagPxD3vErpdHxrmMN9hVhdHbNLaO9
Yz0sXemD1Z2NCod2oY7UXAKC6tSg93D2Eu7+tcif5yMoofkk+phb6bLjYAuTupVA
fX2lTpvsZdMf3YT27+dC+3NHMLvsfyxIjojXhWMtxeDg0lGVe0YKZJsvlZtW9TOz
TI1Yp2lkz3T8/zav76kC5CE6d++Uh5JTVf4FIDfNMJZ96D7iRsGGfHEffJTHdiS7
w+y0ZULy2s8wU4waOG+2tdl87Kpi7OxTM2Ul6t5/l1pmwFUdL+lE5AGUDQuDej4h
Qp0llSxv518MJ2lRpAumkvucbYQ+6yTbqpw7XTeumWkaIV94ezYCvc3/yt8Uj2Iy
nbzdrA48kXOsBlZxQJ3uLNBvkcgdtQLAFKaPdjH0JrgxNbI3sOrNoSTn/OddrEvi
vpNeGtHcAzYZeR01Ro0rCHzR+NQrrtdwMX2+5uWLqqdp2PE8VHApgilSU2leholJ
DnAYkXP/5h7JI310bc7OcfCVYcja8HaBr6NVR2djjj9ZWvk8+fcN+DKzr7hB0DZH
9C0M95A38sIr3hCsmQrLuAMaeYSmljjDnF4bNiir/goRR3avKR34M7p3xiwzZtqP
vN2Hah9WDbKo1gNK8CeETF628uBM1tdTNXLXEyK91sMBEbYdqQW93wI6YC++jkBn
NixBK0qFrZDn7RW/eTXk7kJRy5nnWsC2wSf7JPZ3zNYj92m5UGQRsKZ5szQ3fPdz
OkhyzQjQ0xN8sfj301ye+bPwaiwqatCx4NYAO/2Eb5Re8XMXECh3IXZar+UKLjTC
T93O6bAd3sjR5dwcC/GvzAghr4mE4sd/GamxS6jriW47irY1daSPBdyU/8vereuy
JqlKvawrbkGIg68gSBEzldEq2+B6nz/fj0tahDCjxmmGtvp8A7CUNRN88SAxeZkz
n4aAyZ3TJLegLayeK1KOAPZoHJP/oN/gIOpzSOY+Sjud1zuClQKyb4TE8UChLO2J
dxW88TqoaLZW+IqpZ3yLnlGTotVmVXzll3P32oOrW5g+fWm2K6hZJaPRntLE792J
RetIx0JJXKDPAigegC6gV5bOGK8bdDY+3Ym7+gbTBRv/lXnGQOIIVzyg6wlZW6nj
Q0NMcuCaZY/7wwIbGdb3VDu3dS5qEFp0tXOOKkr9M+SnvQHH5b/fEpJfybVQ598l
4CbcWjrMzJacU7Dn/17ZiwUWmjmfKuDLCQxZEHqnbp8LtzRH3j7QGxi3e3p7M8Hi
WWlJm+Srolg1CQUjB+5VyKqwpgjpcxHx49PMJFdv4ehYCnp2RlxOIQf4RS9Z5KSF
LwzqnJ5gcHUuScfvqZeYQoj++izboKrAOC3iYZwO446Sz3DMJnNC54tzudfB5Dhi
tSLuZeyG50qgGvFHS+B4oKYzSOKzjRxBb6rEWAXwOU/WRIH0SQ2vawG0zmq2WxBb
mjFEASKYutYyDyp2Ml4Jzdrlrq8SW2NKTjoM0OkMTm5JbojLgZlmFsxnKMvkyrw0
BB6CzAsUeHR/20W6xQDdO8GJLJrNstXpzes5Pp+TjRdwL4Krcy9EyKc/sriFEgVy
SfiR05GnCj9FRGOIn5LtmPBmTEzXQY/aIZPQt+R1xKDKA6UvOBVKijNeQyfAX6WG
inbSLRNPL3TDAeF1vSlSWdoyYGMtQrn7vReReWyrWfojdU+P22QqAQLBckvJboln
+2Z8jU97TisGQRleBhzC4noekAbBi44l/zFyDgo2kNkTIr1P4ln/8/mPsTgfU0Ac
17pFP0ldWeMR04HMk66rgyAyYu2I7BjeJ5rUjksnQtM8eUJVNRoj09SXHqOqWrxB
8KNCGKkJTjS7kcvdm0/HTOT/urpiCQ8xp8/EbyjOagM9Tc1lwryR001BVp+ltJqG
HGsKeSLyCB88SEOjoEHeoN55vZOFO8ciFncmLY0VV+dW/D1EcxqQKXrBEQdztRS0
qRJ2m53pGaSEB6i/zGhUYQ5SDDSmfDCphhV7jQnF6THl/RkqWCDN+Aau+Vho8/mJ
oblovk4N+GetJ9MNMPsXfNclhbc44sthqpED010W0lFihJXf4Lyfsa8N6tc5JTEf
lsdGsTlfhjNzsrR3FmstVGwwtqJuyG5glnYvcw4nPg8PI6nxgx9j7faKLo0BdIJl
IOIW2Fr4r2Ffnla7x/M7YsiX1q73/i606U6iteVfJUQ5u7W5I1ZR8sRdfK51348x
SGxtZae3dpsfhc0VVc3/6jtJcsOdo8g8PyAJUhN/qDNpw8ni9/PgP8ubwuh191IV
eyFMLOkyKIOxwyrSkMYkqN9lvwGGd0qMLJJt7HfPr2Y5LLrdbOnWvrGolPOyHGg3
8PmvSLZkqkiN34JXu0hykq98nHzVLAI7aN7x1pVP3R3JlL2FiyJhWwZkIG0+gLYu
g4DIkViTRLjp0IdLaauKLlv2iY990qFqgiEulSpquPBW/kdHOPksruEryD15Lvso
gxG0FN47oVRj8G1pvb3pWkM4SZ3h/FBK8KXLhLB7nRY6p2Gs26/cFo6gtwTXb7xA
jp6zJPVupuqWxpFohrSUNZXSXJ/BMnhBGgxfg7+qvCVDDdV9ITFy5r+HCNREO8Yi
dsiBmCE+L75XO/iS9nwUJZjR6vNh5ARNg0TnKc237iXowvuqG81OnYz+W5eZcS3O
5kj7nFOmGLqfNjZTGu+zig/AQchSGpewHWIDSWw8DHzff69qtl79gc2YNO+D325F
8YllPcxUEFnCEcnTQBIz9qUiyny4tcoSTl+1IVDhfUi72o/QSQMDTctP2yelxftx
bfiWhNOKt3EYwF86laADsZKYu0saXpd6lQbciPUPFiiq7FpGR0HM+1iAx7SliKw7
GoeIUGNhWMDyF6ECsWyGm74l2sg+e5Ni/U/U8n+skJqrmjSJjp8iKDk9LyAb2xoe
S7paZbj0IqzO8OA8oUxXkSTB/1OmCbyEzsF7X6oHO+agctvE/+itdZCcJxckyYl8
zhQpu2HeAdHPqLNnrmg0YqbpPKmmrj0lvYHDLuVnmm8MfB+sZQLyC8BxeJp6NJnr
Le5tCjfu406gBnVYynYVQJvFnLtkPKbEgVcbaxbbVk15akIcmLB9pCVKn6C+1d4A
64RFV//HOtTAHI1nUNa4O2yef23BKT4wkcRJ5uCJa0/IfJvYhS3Mg1kyVPhNVpJp
ABUIsDFCV5x4BRM1B2sQSIBtmtCPNNwfit+RbAzZmQQMEpiUGSPq5p2hNjKEeDUX
SXJjeAv/8O9LNsy+oS4sKKACBP3ZyOhV24XxmeRsod6ENq1ZhWvdUEwTR0TXyI17
MVuEuSkAWJ/cPH5gVDV3RDEq8vkpk9JDOvxFYF0U74gVIigJcrc5IWye10vxYB3D
s6DudUh7MIz0C7ksgvhgmmYoOmyVx/VsBe2vBfzlTJmFdqHBEUu5FuXwFeYhT0Hp
m42f7U5yb/GYhXJ6/3IfJxE+Wm2u59FnnKHS47hjDbKU/w/x2/5CCV+B63vjLZd6
PrZ3/Jj1nNPgHYBGufWBC7O7Jo7uRLGCygo9lF1LSkL2l9z7vtj9O05z7xb4Ds7V
AD+73pZTYKxpcuKb1bm8dh0FS/ohBVoQUeKhzWDRW75Kl6TMKG/tU/ndXHv2JHRN
YOaymc3b+4jCrtoQ9v0KsieoWDSIOjAID+btOroelaw2ZarcZRzBh690kdL5OJ9P
R+YPnYeQCJtNScWMBmScu4ff8Wch28sfKUH+qObGADL3/CqzGxGmGfEfOpyZR+uZ
7Mep4n0235YDwtLGflBU6M3iIDt0ZghqCn1lKsHDQ/eisTOlxZMhVxXwPTW3WIMz
yEUkxVKwdu2CFas9hsuyaOHiCtj2q1oP/nmUVE1jKSdZnWzXk4g46GHQKZxcO9gv
g0gIugiIusvmpkCg6URiJhxNtdKHvgJNAlyLiiSmrV5U3RYaUIZmPgfQ659l8nnj
JMn7Wickw7DRGx/WS8jiBY5jircVQbAoLdXGvETuHoz3qve0LZU+mXDxO/neHOkM
Q3Hv98oLJVWZ9upnJfQnRfdrbK4XSRrtftUrNCBBUaTB+tpneK9K2nJ9BNWnFME/
0sFaVy7KYeFEjtSbwISaM8EfYAqfezTx0QqkgcVwPaceEna16b7ksU0N2/vsDy3/
W2Zmxpqa5pf1azYvbASiQT29Z4E4CffzSAy9xkT42NVW7GeXiT/NDY3A8NOMnAbi
LXZ2jh5N7LnT8lzZPRNKalojQO8VzTqbrCXFby/H4eeGcgqP49iRYTwwygoBSS9A
nw15dvbaHoVvG9mesx1BuXUA8ZBa7VWjCvvU4faGgcpy2FyURi5nqCTcMWen0uLA
f/Ulz7IcvYeGFU58pe+4CLLIjZeY9fgnqg56vcDbp7YbEUnE65Dj1EnncLUL3fVE
KDEKMg3sgCL3FL28VtmuNfNdg1/D2aE107m7cWjQ1p105rMUXEM0Nr1SPAgevjWU
rx2yMIgxZ3QvuT69VVDXo9Q5SkCspH9wz07EyxgvH8MGR0Q0caxZXAcQqIq0CaDD
U7XWPsXSnuvVnIEEnsO7H2mjy5zrDPR8tkI6EealbYVYttPwRht51vQsKK2zFt5R
tF1mWGAQqXU0448onUYf7L45k9HBSX3/29B4m0rpuYtxBFxP45/5y0aNfCwlgLZe
3YRchHSf3j3P2WM6BlTy63c2HLjQW+SLbYHTDb7PbRTfgxsPTsxWVtU2DGWqvAsV
BekGk5vOq0ZVZiG7Z6KaAyKjhnK728aSSk5KJUB2Cpe92V/8BGM5Il2ASPgp+Xid
P2qKhGnJYGxcUUX2ahVrTCvsL3PIrdKnJ+dhFqCBP5kbkV1jPFYlDSWmRSMEwi2b
hg5GMwK11AbdGZZI3xDaKrmpTxdV+tx7RG9Zj5DOetc9+keg4m1FMtl+yNxumExX
MXsknBWd3Ayt1hwwK+m6s6LbDLfePS1CJnsuVK6NjQOWkoEE2V6TSQRP/UUcTe7i
MZ/DBwRKYTsnoDP7erUpCjftkliWVXs5LqIReN9S2bnyhIDFzfTGDQ2MVLasZTR1
CBLGmAwTRPuC1f7SXAZF92HUE9/+vz48G5VQC/YXqJHXF0f2n8EBoR9+Sk5q/Osm
BVuiVXCtYFgEdWBNSRcPwWyh8+Xa2Rrhx4Ck6+j5+DeY7cyLvN3Mq2qQmv/EcTWk
lc2bM4tW5REiIV4P2s4QeCGjVIdnUmkkA/8Lq7SYtAtyO7Ws42UgV2dkPc1W4Wdm
/e86Wn3XVKhT2SVY4WkqvmGdonv0jzTqZby3Un2lc6H4vCiK89TIMx0M3qfNd5XJ
osPgthpqxyD8P2g+Xv9fSBRheXs3FpMP+0AqPwrVFXo9t29ADWFRGW5sxz+OCNHo
+0RRuGHsR9oG0y7znI1Q6LpcaRsk15aDSzWKL2IpjM+V3IRHA2TGJpKSeLIjJ0S0
hovJdhtrN8h9Wut+h5jP8lVLMbGMbjcwor/tl1QdEz9LAx5kDfrkmGvyCO+SzYiw
S0z/tbR4OVHi0FpQfurNusSzB12YasDeo1esvVlNlIholB12BGEdc7uSh1+Tx7Fo
efb6tuZ6rBAi9XLpYFLYo//tr1GlLdmyQOfsHTPi4e1bJpKPXnfhtIdE7EWGljIH
413p6WniEbo2obnFYehrEb2eCOvs8Jg+nvJ/0uDuhDjA6QVN7aBLGQG61/gba4dI
sErHdM5idTyhG633He4NofAfc4qIAcRusoW7Cmy4PQz3rYuHYgvaNJDzy2mAV02P
9iXucC5WxBQJU+lS/dwCenCI1KJswiDAGoIGditbg8NM0CE7Qg0edVhTK1TERoq6
HYFAIoUH3gP1gGCuHQftrVFY1LTyJyoHcUfilsw9L0mP0D1QBGrbB+EAI1t0g/sJ
iLkNNRAyQy/X2k2YuLa3MPf1zdooFI07mizPWrf/9ZWMxGMR+orplW8LH/y6BVcl
QMrNtENGMPNky+U6CfHANsi4pKC5jDct/pA1LJUOyeGUPhndQfHoTwGZnR0w5ul2
hHgam4d1xHZCmH/6vuXEfQCyP+5AdL+l4+41Z7yF2L6M3RbJhgmCGuOsPcKQzUQE
Ref0NrHYaGq5WpWrHVWqWhpUPTbYqWYXT2KFGGyUHT6HNRC6bxm6/NDA67Qtjblt
x5LjZx0NQJhdEuMZSgId+g4UQ215LFcpcO2qilzPqx+hPHW1C7iyYWAuRllEdxMV
BJDT7njB1QfaqvQ/dweeRdN8gitniN6XdBhtXKqGE91ikC5S1jJBvyW2GZ7oPfXO
TFmfkf5Dg1FJmnSHtdJewl6YgPpONMrjMUyVYRSFad8eP5IG2HubHxiV64aiVHe5
ZGT3eD6bRRSiw5q373pCrO1EDtXj1r8gCGfwspZPEmiDuLWrClyDU8qMBApzYWJL
xTQTnsIDzdtDiB46tcPBA6Y+sO4AB8tZ4brOlwyzcJnEA3ip3pEzT1Srt5ixOnQX
jE2GlEGG5HHtyYhcgShG7fBy1nj1SveCvPsnMpAnm+xBHoOzIl+mPlroPkwdFPZu
6eighOwyPMB6EsKbuZyYncoz4B+kQcaBWlPUUKk5XJfTSbSzm4s4hcxe8Lga6TFg
Ysh1Wf7D27xF9rtP2Op/588hY/cuTRltHQ5cZcphwAWWU9W9pA650oRtbCNvAWU0
LBPNdDwt3RGmYBMEIMcrawt1rWwXV53kNas5HUdXL0ecXzq/m3rb4YZ5iPZbw8Js
LkEb8JP/JTh/hYNqFOD7fFfV2BrXmEzk4pfjmsXAa7ynX9SbqfGdwuCesk2RsPPT
f1uED56vYrEmtctQGbrWukVAopc5GdU1DUH4srWbdCJjobx53SHxTONVaDrtuGjl
i88ZH37cKD82XkNjxO+qwkG/s+91/CYOlliIaw6MpWdHuYH7IdkM3/18u8SnThWk
rgqNJQJrFnN9uiiH8nGUINhAT77JU5xEhi07gNy2JyTlhASIU5Fhm06859h+U/w8
WQPbo5+8Wdw5j6pVXl8lErulwvTThGX1vDcE7Ky73Bom5c6/O4GykbCDaSzdKuiO
+bW4mwJd5vgycvL9FO/VNK9yL34dR0TwE4EjD6zFqc3D4FG1WrP6kLzx81kxTHAd
JYbCV22wn0/kZ+MmVGkwe1TMs1mRzcuAB1e0cSQU0/8fHl4gwTgvvkD+ECcF2aVh
zWSWKMk5U3q/8pmIOBGdxMQe5uplbCW4fGmARg2XkkX0LQbMmnvrhcsn/y27hMbi
GnZJY8wJJyRyFsXn+21FoNlqS1RBAexz26VWnefHN3MQINgO8fUdpT1sJvJ8r14B
dy8/MpqTu6c5In7CyH1VSVpleUfdv/ctiy3MFGnjVc8UnqksU9oXO9akoM+USbLT
MSn8Mz7xqM58Nc8EXB7mojVlPnWhdKJKSSfqxgRIcYttRp5vhbc58KFSZAWahQPL
9x6LdmcQz1BEpZIFld8ZJQBoOXNcsOaocy1G1kN4Hx44bqvfOIee6cJxK0FpOR8f
/4ZomTwIVa7jfvzopW7G1Z6PZhDHUZIiQKtE6nU8S7JrU8pXzL/BRgqgVsR+2uS7
ceGoEd7xyZUOvgRJFfcbxjB2hl8TMX/Pw9C7WdLiFPNC7v4jkMn0QBxyRJ5PKyaw
6+WkkBp0S0fXA+gA9QTlkY6L90BNLpzmaPyiS7SmWmvE3tOFpcNg07z0ZDQF43/J
WcrDlchqwchhA4cL8Z9RK6UoVcpqFDzlRpEcEAluyjoVntq90kIXGqALfoFN32g2
nugOasYmXDcH5j9j0CvDFBt8gilJI3KNMspo6YnTsRIhNQ+u82OM77BFDcMwe32/
VUdbyJL2rxMi6lcA+YkhyrgAE8y0lEUa8o4o4lDgj1yJdeuRNhc80SQS7KCOjIeJ
+iK/YBIGYIC4M1JCsegnIeZMCuG82Mlpvabx4+RgF/i9k+9J7LR5Kcq+cKuPs7jE
bQ+8g6rdASCDk2O5LiGFU32tXhF6JLdnxfzvo7lulwtFAQz6EK4YTNssNvmWd5na
z1HjOcP+h0FZqj93mF5Dz6OusctYWA/qNpcqY21b8fNIk7E+oBz+PiJUwAyqOCPW
Rax8L162HkmIBnvjCqh1R7ut1DAnCq6zQ7Fef+m4YAFhDLlkzI9p5BQLcSxe8g35
jeK8Cw4OgNvdk/zyT+zQgiyp6Lpv8hK+WGd4FLJzXPNWQ9JMQj/OJh2FAkoYRc2o
LXdgON0M0ki2hWHGE7B53E7D8qig1NUcKiZKkFx+iiULIyWIUqbHazkoA7AmSQYm
QPB5VsPhm75RUag5PQgWAFECXFBk72zN7Wdfkgj+P0VLbPcgOCUzRQOUiGcwhV3F
YlPw8syRA0462gfCCAIH35E4vR3pNs+Z2CY/958pf2MU4SODRWrk6Jaxhn6onfP+
kwqR/1WxJC1XYi7ZSSL560AcUDYPhGj/EgrCgjYNvytz/Wm27QFRoDMWCpbcEAi2
MZyA3pitPmvUoSK+PiEQubPvFYBs4tbCuk7igGTLyrDi5nlBOvL0CciEVILSC36n
rQgJQDGwYBwxtBj69ccGVUbwIqxp+XdWQOj6yVXWxnW/KD7UMmapKg1IASoNrmEj
bKFcrBXy4cyAyPqm0AA22PQLIx2DD7tH8AFdScRRVal9mRTkhwzSI2m+RQuu5yYJ
DSa/Mr7hh1D6Tt30nv9P4FASw3sPrEsmFz3hrYy7BlgKa7+0etDkVSVe+hbeVBfm
Gb9r4bxGhzp+C2OqBpaEoxD9QddNd4CME/kgtcIhpdkRuSu1k6lOFGcpfN743mUp
J4sJ6TFJfUNK6ih9iwLgvun6X9vU9mkcuvcbIjXmZcFDI4cMG4zQ7aW4KVBpc/kp
iDa10r6VJv+/T1cMkJJLF8bZ/4YT4a7SPsFgn/457MzLk0Cyx35QwUMojnVReMRK
LuIjsg5UvzCRiMV27Wlf887s2H0W8nFiEn2i7LF0+y8JRnVApPa1xUh+YDoYsgAv
nQdM/P/PiR3dFDjxueCcRkQRzzdQUpR7YF7VYHuiq0JuJzMXt7uXZuJ9K3nSGjrL
MBi/RMU4aWUy23M69WZlp3Ga+jJiEwj9jfyAjl1oByCMNPv72mo+hGvL1/7OxTgP
uC9WG2QfvFz/cMfHOIJ0uqLYNg50rInydQXKbPeVY3d895KOU8Et11qsUQFnC21Z
0UQp7cdJ/5G9zDRDGJwhoHwxJEN4/ks1EHHqAh0es/biTIQXEcRx7jbiEqGtbvIt
PKZWlqKHQOW7E87alB4C9lzFvq6UMjTHAJrEE/dxv58fDPxbmIfdcIdjMhPp/DyQ
wsfIfvROZdTdmX0asAeZnHV1YG3wvo9lc+wrUHWgsVkC4O6JIbvgc+9VVOhJNral
gGTlydh33o3ztEpeBaPg77OkLG2JUIm1wbSMdq0X4AOZRJrvD99ukKT7aT9P/U7+
B7cvu1z+1t6Q6/Gbak/EnR7MMM7eN28cpXxpX+Is7ck5ovTvos4NwcaHMOsAb/TP
I5cdMA8NiMyfkVRAi0TVj2Q7v4kEiS/6dxDZqX/CMNnq9TASs+k0VuT0xU9HEjJ2
Fw3v4qZoP8w1Qx9tNS7pQPYKxeWm19aR/0x+TuX7Aac7WElsfp56izQ8nyjqAY8B
l0rvLVQY41Bn0vHusFmX+W3zJkW9GzA22iEPWo+4fw3qE4nI//sLI41oK/5QuyXi
9CLXMop04aTP5THTLsrItN+/eBgEIx8ZS7fS7SG2/BvW9hUge0W/dWOpLNcV3md8
74DOxiQa3ecdIKtTtauwpJHotzhsyiSl53rJ7289iG2m7yqjayCaxPQ1quWJEdyP
I9FnsBatCjC5ztn11SJgB2PKZS3/N1LW8iQd27dFEc91LjH0fW7WusnrHhkSsWF0
cpXYoXTalOg6iFgXWYqGURF0AB+PMV7qmrkvbWgWjMS9kLIiqIh/UMKONHO8ohAn
vsT9a0QL49Rz0eb03Yj6iqRf2vYwWUGAA6o06CLcKSSvSc/V2PB7kpjtGcu2qgPW
i786fo5sZpuuKJ8l0iZ+z1INKedtOo5mCpsuaB65r1/GNpgdiyQVszMLw3XZTkOL
eC3pnHOwnp3nykwZPBnBgk4Q3xkY1j83Xui66HzgAuGB58KiwuhM5/p9ZGTdKfSx
AstunAqWORPI0fRXzqitTQrXCgMvkPSeStRIq5TshFvhvnIe0E/apy+mVtHtaGf+
dzxOzP6etlNWcY37MH/G3DFn9LBNoVl4Znn48YB8L3jECxp29A24AWENqvBz9xuA
piO4kyU1H6qSa9YgWJV6AkwuigMgJn+ohQaiq+07ZZw5uBwKhmRTw/WngBsRa4+4
knlGnlM3NG11sWNiWAECw8QxqhpS8uWb2MIAqe5su0G/Yr50KlZHHXrqRFGUkcIL
XGF61oc1PmDwDYKqg8y2HeiBGeMtZGyDAKnsnmJD+yZhLGTn/uwxnInL5Nxkfxuo
/q5HnvsLWvyPla0E1CCWRLxyLQXUw36ZjpDpgi17OL8M3IxVUmp90QCu6OQEnAlS
yuLNowCZxq1AyOYfkM9jXTO70unzSfhGkQcsBrTMUzoxNisZ7xkeN+N06wotmJnJ
IKup+ZI2eblbDrprGZbB5C9c1gIdSdfSFedy6r5lEjKGFm9g7Fd7l1KQus4EaKVX
B6QaxMXZjBCqjk7PW6t7xM8gQx5EqrL1ZKJG3ESCVjfslLHS/HOR/laOgteQ7+Zh
MbCw/g33VKnId/46Deqat83J9ykK2o7ob0c+ck+mdxIQLKQIn18TQzZ/tyYoEPFI
33lRDPg0ZYfuPoKF0RZc83dQPO2BfJTU/XgbcEML65oG1OSOWHNI295WiLdR/eAj
kGiE0iSI5/WYEvLO2KURvlpPZhCwDV4JFjZ4/fnECBRAuCr+AMgubfrx34OiZDIt
4tFdr8NIWaOnRPy6QX0FOBbQMRqM95+xWHY1PunAajhB9goA8v5bHzJ6lcxZpbIM
cTiXtOuYPD/YR7WENn6MAmans0kJkf/4B044Epnq2/6EVavdF178HHdLKMCMrHdr
N/auABfFUkO0ViqUsagGO+D1qH2QfnVtGipvO2NAcGY3Kgn+Fbc1ZinO9R31+8Qq
LY3ryuruAFrLWklw7pRPbdsSFf1Ly75Mcu5Y8RMf6xfzrkXjNiF7wPjK8xkz7WSP
LGj9sdgG/5zPrdx+xF2KdbKVC2rMa1DSiyo1J/x9e2X/SQR2Ub2OzJPSMaWaZDnS
bEN3KfSsR9kbnfXFsFLvu1pFB/x/0P9kCMdqFsy9s2H2jJ+hfwv5XslHWJfC2DNQ
66jNMs4O5lucDY9TA94Rb1dUbLAGwcqDIQ12VEv2pFk2JpKtm3+LF7ifBhNgFQYr
yziAQYPKGN2LESDWpU8GhT90pRq2pcEzONvJBBRVtvXhRcAVioBfcD0I8ccizj3M
my9rNKHy9QDkn7TrjDd7rT8tvQN3lHDKQrlQ2sMfQ4xREV62+0HuxViteqZqSb4w
PA4PCvbIT3vw5H0AZstwgsO/IA2P1HNI2TMt872/s0XHc5QSSD5/mLIFTkZrJPBQ
meZSiWe/FyxdmAOF2CDctkXgWjwNuAIzvJyLNHTddTQI/QlSL5Ilx0nYB29BQhkK
ki/KVMg2LBtCU7fBNMVMsrY6WJbgNput4cPr0tv9VIiLdpgCMsdAGI25WqYs9qr7
VSa5cY3IhbF2gx41mbvTQJb0udYAmH+7BHrwHDh4P5NSOXYQmowLcQhYJ7Gz9LqU
+SdU9b8KpW/GDzkSTBM38V3SU3vl3NDf5LhG9qsy8eh2/TKCcu7aKPTlaFmPavSP
8/Vcb3EUXTQ9mITOSGSEI4ZVL4Z+/Msv1LxQl9o0/Tmhg6V45RtukcJaV5fu69E3
E+O0sknei7QUeIdIIWOloKJgTZ1sB/LP5TeQqrTdEBI8CXi67mUT0yt8ncy6odit
jm3piGb8h9ajHYco4W/9OwE1g3merNljQWAqzqpDVY35Qguu7Ka7Qcju0Mo0CLWt
+9aAmv6bqcgHZO1iiKFxB3v8b5Ho4Jrtz1OYZSk+Pbj14ro+7Lhcby4PYJth1k+c
kZq4oJlX4UiKq1Sd56SjHoMwoVmn8B7J41TBSmWaqlX5ALPzGHB1yhFauCzKB3YS
hEeoW0cPAZuwTFOU/1BJ4R4cTo2rm1K5AD9nBRUdVeQEzCFTodXmOXutyXjCDmLu
DmGvBQ8FnDEqCDBbUTcrJDviVkD1gwYWc1Ey+cdLkoXUT/2Qe5WKaITaJKn7n30W
PjFtruXny+zNJl/g+JhLGb9D8BsDhWR9VcZNyAOqltgNr4PdbIpsr9SCzsnjxHK/
iy8XD1LwXWhGWLYx3wCZ0gJ2nGcR6Vpj/rvGgZWkBQYBY1kBHGKYAcI/P2MOO5fn
+P7SLWpyLMohVG0Tlzltbs4slGAV0kmpRioNV4y0HM9ZJ7itn53OEYUFXYy8hu6+
ssSNR6J6Th+b2yl5Q9qiyrbbxtHEY2oM8Yi0+h2dnv6xGc5v7I5WDPhgl3A7KCZo
Tn01oqPx9WFfccK3B1ZLJBMd4yvNq0kuC9LkfDIAv8LJXwBd+jiZAIG4z7qN+VfU
2dyH4S8UdwK9wFE2RNjUkWkEN438XdwHua6vvgkj25pU2TvCsRU5FncasgQZdshk
m17sqM4z5qT37fl1UMXvid8pHGolMj0Ycp5nVcS6V/IOxnLRGr/aE5SEvuAz4ylJ
T0F+vr1IlheDbryW+cJGCO+N5IngeLqk3KZbHl2iNER8X3E3pGQlrK3nzg456oIH
XbS1yBD1kkEFEylsWe+2oTor6EcLG27IGAAUM0TkzD2axLw4MNAoDjeJMidB/Ru/
Lzu6pt0W1lbd1eLiTWia07L5VBoluE/Gv6QMKZwLh8SsOPP+W/luaiIXNh7iBQF1
+Si1U9EOoXJrvancT4ELS5eZlekJzj3ELHoVJO1NesWTwPWkoMJL2KN7reK11pD0
ObPOGsl7St3LVRjORqvH+wbR9BTvyGlyznjdkDXTjspgamdNSBzl8fXMDdKB0BT3
/oLJ25P96XFYPH+BiMYl85Y8DPybSKzcSRe+GQB85DlvoRsi2Tsx31k1t/Xs3b5U
Y4j/55VYbduS46zsCZdKMTyuC4Wx2h5ch2QAryFHTTJdRyZ9PLiWLSlqYB8FyaMI
IprJQ77sr3+C9SwSpOg1wiSog+T5FKCkI13b1SZ5IG3GW7wgoqo+MZ5FpuIhLlVV
/EoccbR1VXt8LvExzX9N5Vi6LvPlEDbQYkMYyh3qJ/IA9z46ylBeLnacafwwL1SZ
nWqaK2pVebRBV921sClcT4g0iliSznLxa/xkFH4E6yJaLyyGzdOBRc5kRT4tyMcz
+9rJOrbE1ToV1SGJbMAQCmiPsB1h4X+wLEURe93+3HLLbvqGs+qqEUZoKepYumQ0
OuW6GRSp0/t1uEYa9NUV4Dw9B7ybaV8JEWE2suLv8e+y959WWbo2LskzrQPTBVNf
XlRL6h4hjP2U8L+l71w73NQpS8fKzzjbZze4SElAZ30VXKVTjjAyAJRt5yrwR7ho
hi4SyzL1PJAi+MLZu/uHm9BubSsw1AwxI6EKbtzVs4+FngSSTt9f4tJ56DfHRykQ
WxTeLWxPnfOhP+vdvApP6gFH6Xv5t4MkHWViZ8X8fP4IwvTAuXECZ2X+8TW9zjQf
Q6iU6lwGHTxZWERPRuQN66qekgpZWBPjS/x1hI+EX0A5OYvZCgRCH6PDBqZkhg95
sSDaYvuZFxX8qATtc2r2AJ00zGfciUgVxPcv+0xktPUH8qFLDxE8rHVmJtSjfnPZ
uOpWw7G0bXk0kKl60omLgMlABQAehu2NZFL0XxgjDlizi1ufDWSgcoxWPQYxYT6s
2qla+0HVZKQuxfghHuIsU3TsuR6DPG8lHSC7RdSHsWYAbqVri97N9iQYSjw4LWaD
XaE7rcgT5My0yUsRm/QVzIpv6C2/mJVkiJy2u/miuQ4dmmuhI3+GnHYjLNaCT/Jk
MbPgL3UmSdBgRWMSBlHaTjzOqDnz2nyLoX+R8z08umahvMaxBUDp6xfSsXFcQDc/
bKkhheDNH6u5KECFyAUPaAMcEthcjfyp76FzTfhzgHwB1vr029aD0FlQHquqabsE
B3Fwbdc5THDn/8Jhox04XPqmOC1rreWPMh6dcyn9oZOAN0y6QlW4QnvRgOxS0MHX
hw+XgdJpIwwKX5x1PMxUO8VlP7AVIhTKgEtrPkhVkcy1NCtIB6J74UnqJFjHc3HJ
f+Bv2oJIthbU+u/iWKbpvBKtHfegBaUuBSx0XNQ05vsmL95NGZWpoW8Y7vlglaHU
FbnFoTJJNxZz0m70awH0MpafrzlHgqkQCcI1yO6xH92yNtg9Vb9lI0tG4DpHaYlP
9fjP/R65EVWEfm6cOkxUpP3hGJ1Nc3CF9ss49TINRFTgxormMnPn6cCGKCsMMYoL
2KzlkQ/BY3DE92pGV2MUyWfxWELr4/s63hokDf8Yq7+F2Dv0dP36YKbqhAUWuSpj
QvxeJdswPtLDUUuFftAGwJHi4Kja12u4e+jSwfuhWUX/5R06/A7lLrILzjJUkn72
utI/JPcKz3eX9HZNbmoHm41co4QejC/8qX7uJHU5hg1iGwd45ox5WprEVvujuZ+S
t71RXE0isZiqiZ0ksr1OXvSudeLGryVa77onyar2/TcH/c/CO88JCQhpsXErG5ij
eV3cO/yZqAKMcOSRpsC5ov5tiCB8Kcqg+jgRl7C4vfi7WG3vBaYuwQjA8TisYux6
KcdzR543uEGf4BVjCBy7BvW8vv0ID8v8h4HpI+zk2qQzxDQrzCdODY3QCGRvWeS+
FXuVMhc0CwVNmtSkjGQNdfT/zomBft5pzoipjRpqkcyKIjvgZyXhGx4Z6bzH9g8h
81BwvpUe9JHTvChA2O44nEMkgX76MvO18aBVGSm/Kxpx8OuHF73Kpj9ldzbvnwkQ
zx8MzxVWja4p2SvQCEDEK4CEgeoFDS90GUBNBCnDBdibGQF53jzIGwFxycA2G5QQ
P6zKHGSrDkoaBIwP9R9dk2KZz7CrDk+RifhwVUIj8GTDq4kEfhM7EIOrVOCrzsN+
W89cham/8QfaZOmpM9eQVwt+PkaoXAIYAe8nEYkVxdEaixjsM62cAvtuMD3ZfSUr
ZwP21z758BiugJ8zikLLhbsWoEWthv5M5uaasuePMVHeNYb9Viw3ibv5Dzj0mHfp
Mur6BqLgbEtikZd7rG/XqP69/BQHY2Kw/CfpCBKpY41GF3RCV52PuRSoVeYwTyAS
AW6JPEa1k6ej29pXEbEt/1Q9qOqWSbqlS+Eu2tIlF0o83HGkzr9BFeK8WC09xmjF
TjKabl8eqAqp8/wy/AazE27T4DLlz9oEy4lPkRe+D48lX6pVL4vRAHHcbtEE27nD
EVK1B40WfBnICa3fY+Ovj8Ur4+rDGj3sTO3bJ2bujNcj66yFr95b8l4o+zE00uhi
Al69mDd/3eeeWZiVqQ8UsLv5A4mTb0SIcgh3mFL2kyxgT0d+LhDHteGRmDdx6l0H
YK4kv+iSvcpeY2qtC7mL5xWIA3QE4AwWrz6QYIxSmw2/cTD7t26PKOiO0BfUB8OZ
IFNE2lLncNCyBQVjCDRPrVlITnLJFkJAgZI9qc/YAqGtRYT9sfVfDO9WQH6s4YWw
xZUN+qT049FUTJWrSifgi3snno2q1jxsh0vo+gFdtzPCHFXHvdUih/FwSs0mte3c
SCYB+8OBXUJrSux67ZvSsPDZImSlF0He60R4dkojYx/5rQLUb1p+OdpWtXA3WStc
0yn+FgRYVrp0q8l1yTTpwdjO0HwEoVGu+T/ydiihwyUaECZLHDl+g4hgZQQ390nV
7Ok9HXjHENMihXu6DP9Vm/adGiQ7PKrZ+3So+oHeeQnJteVH3Kn+QjjTFrnkvLP8
U5TcviInaDoMX994NbojFTmldGHsMUgh9V5rYQoE4+oIVe5EwBj6bThqDPiMJoc7
zIeImLf+GxqZXLeyTkLFfkAxzhaGvAK4MXQH07yOY6uUOBdAkhJWi3OamJS4qp1q
KEBOaSveVOvu21EMJHxL9HhASnK+1G2iE+WiyYz9IwvE4L622TWG2mnGE/hTDg29
MlEU6+RHBtnGRmd23zwI5gDpByGvpLnSwWJf2wSGxtOGWBoMGlaTnT5/cecfuYID
quxKhMZ7ItEcMXszD2ngf5VcqWDlbE9+Aw7ADmMh3vbDFnHIhN94IR7FckugT6cn
pHAa2h9krEkNk6VmkV/lK9nr+81mcSVEczyIX8h/0cS+OtkFyenlBTlpestm4NNf
iC3Gg/OMSWwhSZzcS2vOGuOUXo8PSeO4jAlYxfe0qsuoij1R/pPlJhzHy9lPEB4S
oZNty4oxju3XbReQE1i5tVZ/S/W/GWclvYrkG6V/G2mYCiYXKd0HE0xjxFWlIg/6
fPYvOu/B0PE/6iEIaBQbuLEMw3P9VRkD8qrEMhxGy57Jh5vHDU2sET2PGr6gnOr5
0y3ipJYjIdOwoGg5byzLaSDEr8wPD+1PLmZvk6OcXlOyGqUtlLRdKwkdS6WF3TYn
9P5bapDbDNRf2vnMhzpMnxdFm8JphezsktQgd51SwQsxUDqN+XZ6RdahvoaqGHI0
LCF0JGM5n3cMx0ECwLYSLQKLXObmejf2C/DH66rAndJeqEOxPpR+SlmGP6olhDe1
KRmP7caGahAkpM+E+/zCQH4d+Y2JeTcy4eekHoJyUM5a/gDmJk9lOnojVh8yaH8i
sbTnVfcGIlxl19PDsJisnOwo86+XC34gysxEBieBs2vPsV/OiUhz2eid1Fh784Lx
xaI/CMqav9nmwYRA777Q/LLTTdr8W4IdcThln0ruUg1/ge94vNO6+J4tZIgFrxOA
a7wIdJjmMWq+1B/OIryXCpOPwsOcUwAs5dthrKWG0A3vRc0mAomKFENiLEcPTGuJ
kS+6bDrnPGxOTAnKPTwqLYGDyCqUIvOLvoZ+PyKc1Diuo2O5rDuAO2mKpMF0QEHj
gt2UYd3CzWL+FsJ+5ti6zHOl0vgRBN7dOc6FJY0l74FD7ngk1Lk7jYYJ8k7Nf4a0
N1HF/AlcvGUoy6ZeusWrW3NLeUH63kHkrHykpvr0V0VCzjAOUlu/N1tqhoQJWVdW
YA9sQ6TObAdwQaDkbailmIQRvTun09vL7A50KwweJN6xf/5UbsDHbPXYwOjK2l/u
MelpU7DYle/4HGvkkZX87uO0wuD/lVEeosfJlAJChTkj8pB6UwvSli9Kd1WJVOR7
RjWDVsuDYzdDefxvU/bmZx+QGC7UPYm2m1NsrXMI80n7BNad5VDVgvQJ+4AcEgnA
gfe4PSTuLOmy3RYUtDuNg8/xrz4TaQoMnu4xohHnQabgvNA88mG0gBau0vV6Yvg7
TURgo1MLQLVR0JOax1Bvm1y+CwEzgP/2xxOvtg0Mh1nYRe3McsoqWrTn7t8whPpJ
XTuneQek2SoRfSAPlyH5cmYYWWrJk7oICatCBxKAXjFkqWtvcfryjq4oODsKkifW
Er+EmZ7BI4PI1YvTksvxkZ2GwuRNeDM/DjGgzGRTZAcIzoLQ7A8NdI2brWY4KbZg
PmX0N2y5i8tb5ame+6BBbt17h7GvGPGtmhzVVHBnhCIWXGsJD3ZW7Ibp3aL9tVXH
K0gFEb165gVD992i38oqPix2EJiwn/9FPL43EGutWMXoVVnjGQ381OVibcGy2Egu
B65Y+6xrlwmaNwXvUStCb7aAMrMeNLvH71ay+MFmdQ5XtPa6yWlNUd/Rrev7EGGR
SSk7umwLBLzobB4FaUwxtqP4ALe6srC6BGHoMQX0nmnrkLaZPa74iES6SGh97Y+0
E+K0WaEBbBwseHNFvXAq8Ojw6coSp9QaZ8yhqHhndWFWy26flGk5vFcE5tjhR39u
HnQ5z9BdzP24VB7MQANqWcW28bgLmlMSj7kCe8dGabnIvX5zKJCHgY8u+owKlwy+
/T/ZC4kMZKyPFPTt8tpANnKMUbu3Qnmr3Eb3c79aStLPsLIU8c/25VQTq8Qfj6Ef
lxEMUfJUowRaONWtHLRLicI+uvnu/C1YsL3sptfznBPOc4QCXlNFytYb79WYXS9e
OjxaZ5DLkW/ihfLhBxz1c7EtbbEaUeL6DKRpB3WhtM2umDo9uEoK9W42OcMLOMS1
G9kZ4UMr06XFS2IST955QTSJlCGCWRkpVleAFiQRYSxEmM+zuyokxRgGcnfWhUSY
sL12pquSC7XeONHzdZxGeEVIBK7ZEglW5DWf69yGCxR8/r3l57LYoC6g2gg2af+M
rqTPySKkEO5Ks8sOMey5kc7sLNgnO8DxvCQV5HnQjqAethNbPo0VbECKeL7LdlbF
nfyI/lNKtU522A2kx/Is/LRM0TQHPAQbBVEv7syMN8/g3aU8SGi/zmqcAb1pnNgh
+v3OHJNd/PJUL0/tMBpy8UB5HsmZkzJBdBZu8BgRn6gFGVhOlKUh0Zz56Yosj2ae
4JUlXwNJu8SfG5n+WK2ASjqDDbgQRaINJo7eKhpzN27339AfBfN6Q89DupOm3gzs
vvLZdU0gab2gdopo7Yad7Za+f1xMUxReTYSJjG6VTRlIVc+bMVgXD9nqrDkkGY2S
qKIAaCu6YbEbzw3drnh6ZHYvj6Z239bXpruGkIgZD5Yu7K/V8vC+vdY42whtOSEZ
nnQJxSn7HbBjE5suFWuecsjX8XYzV2CHoVOcPJSkYS8FPmJvFW/PxXvvPQZ+po4j
H0DrjskdN19XfzXjRomsu5Mv3d7G0qTUI/uZwJWRwSf43bw/HkP9If53zkFprkJD
JDMTiLMLmPuQSo1wlparDhdF5diNE/cHIUo2JSlw9hYkRI9E1XiUljOTH3WNtSYp
BNUzg03ffDATgPDRhMozJGnprmx/wm4uzndPvV6z6rH4wM3mrlZH7/YhkJVCYOLp
W39YZvPyGZaD7H/A/Qa6cDJc5G1lnucLOHGjc38lSMFo5SyUOWzpPTYX0qGBCigj
dFlfiNcrwYv03LxuEfXRJzoobBr1ydZ5aXIKkacWDQAJcRxEWwUZTjeh9v6yfUdH
X7qwWs+YLM5aVUMkl7Fnsa5MoVrTtVGMyqzZHMXewYroEbj3RIMGU3KvsgG33m0Q
7LizDlkyBolBcDOSQ0uV5NjXeKHEa4AQbcFVFdes+wWErAHzdf3HMnArmSA3b+GA
NQd3Iwvp4NE0r3YtJ6LQRySf6hHvnltdLRLbHCkwzv34eTzifnJnOF6arhow/aJx
8oOXTUfaWMAo/98j690p6NnP4SN6ZxJhPJLMuIDEjX51Nrk+wdTC9s/tH6ZGRrgI
UFIZQ+K/yeKW54Kup6+0OjsW7zULh+dPzQA+awU1WC7iGvhsZK9izJ54s/C7ckp1
HilqZRUN2hqqgSnUZSVjewfBr8EWVcuJ8uuffu7Vgkyc5FwG1A9+grXSEvKhv8D7
81Fqyq5dpnjV8JMNX9jkrNdcEvYyroYz7ZSfUB97WPPGH44/xZP2pQ+BYAVetHw+
6+qoryr4hbhLYKYqaDl+ZCsKjgP0NV1IBZErBqNDAXKPOjX3YaVNIkx9kzo3AGqC
eWzRAqh/HJeMDPDIpTVRVLGA3OdNfiLuC0+WWdSbuNvtctOeSdYLiKkDUWUjg4dk
LlTLyXiZqWS+rEdJ2NDyLu9gB7/+Mzq4O0cJ2jbwMWDfcBJspVmzNCJFbBQ8gpBP
4iIMlkP+B5LlGua0AXmCrQ0lstbt1l0IpeYOH/RbFVZ2+Yf1d0q41FqRDS06fLYG
PNrT7zwKxTJSbZ0SeqOpeOxsITEjAkN7dxJWnyji5ucftRsdfziJNKZFKqyjeWr7
nZCcBLiOwdAotNx4cRTi6lXqfbZmaFC6xwbYm/tSBhgT6cRu3bQZ0u6CTAfYHlYK
ZhUpRoX0HIBq7AkWavH2pW1EnCxDyYCWWSdWHaOO9/0gFgYRQn2ezf6iH3gofNAz
47oRh6M0slCGKaItJoz85OOMMUn5YQf4nx91V3oyznW+WjVaO/harksuaLM0W+eB
ek0BcUWY02sNWh3+8s6MKx02gFVSJYp3ICXgodAI434w7Wt7zAh6eC9lnUI/d0Fv
L1W9/nq1c0AEtVRk6daz3e77U3nDZRqTwQwg7Y3571IjBCFumcBuLLDUnkB7PIlZ
Bw8jT7UGkKlZh++gWYll3fW+kHysU6VK2IEwz3KueDoCTgYj3X9u0mpp7uyOJxpR
e3gJFL2Rjo9zH1mUN6lCLv2Ld2khYO+8XqMSg7eAvPzb0Hlz5aiDCJkIzL2xymif
5Ls3Ql5WIjpvt931cfoqFJY8zgInyT8XqdnzPGRBORPPTjot3hvB9MPBuisFrb9j
Lsl9eO1iqRxkHRLFwf6aIgRRHS1921bQf1TpDezUHrjGPTsUxIQ0h0uj2TckLNZj
ovSuBYacRE/j1sfCkxmoztyNQXuFOhHQ9Y2kKYf/dtrnKsqhreCjH+98bgORaScn
gF+jooDWrUvfX+heYPW2lW/GHO8uv+Bjy5b73q1uxcLb88rV0QacXMwtr1BwzatN
mxWLwOyP0ziFADK/hxEN8Owt7VprBs8RSAgcFIlVj4cScgE8pN9BZMcHloZgOn3k
hee8nPLNaevscbLNrqEI/Mb4nQ4E/4tn3rgScvQLuocKaIbSqw21NkRPLSN+JY4G
0knVM48kOC9RBJgNu20j3cySvOccSauglCw2MuFB/snoSovcWBrKUK1r0/dihGre
81drGY9CWXRr4zGZJmuKcGpKuXMPYBT563UGPM04wmnjFt+FgfvrE1NzzdOAGx4w
1wjX8QZel/PZUfBkRAF+k4yh1Hawo0zIENPULhUymPxLIYFwR40Tf4v+EvmGW292
5AH8sNIPbHmSEWzDyvsOAPuyw0uhydPnThOCebJ5Ddep/hEPVP+x4h17imAGi+Dd
tkKqQuyUm6VDSz7zJHLirj8zg4DCrUw9suL4qILc3/X6OCZyZ83wVqWsF2wASXra
w9TChkyKm090M1PZZ8jD5NAstmzgWKfFYrmocViPqBV1gFKh/+PW7ndDI9ItGWWe
RObhPJ5w7DSvD2balofJqBbTM/O5e7NI0DMQEqszkIXveQgW0lmNqC4ZNuVd5tnC
KE6blY0nCe9hkOe/xE+iJWo5bOtR4U4YJ085pdD5D2ywKZGTtQmZot91SmkVbg0L
AjnvR+n9O4GeUmqi/SvZWqn73vcbfSmpZ/Ov9ykCTYlo1enyRRAw4PGrCWGkM9UD
i+gfS7l2SIoDqwUaWfMKZQ7Vp6TGeAv83Q5JQzm/iIE8ZKkx58ouIpCRLQ5PjlGx
Mp5eGEHLQBTULJ9gUnI41bNzGzciBP9l15jzLFxIUxN7oDDovw7LjoIU8O+rYfJH
Y75yR3i8j9v/sZ20ALguieGc6Gh9XMLOM9SCFXL4aUSDrApdDHn+6JGRK4ud/qTb
64CP6R4MPEXWF2PrcPpJMhsVFC24LrfGloEXwjsyBhvBsSbCSJoIiK+K747DHWBV
WYnjcPTyNiZkCDjgkH+XboWaz8jbJrbtOsip/3WvkQXJUrJdkj97ZUQQm/tNKJ49
9OzYxp0CWuE1dGFBVmFLORJvYCIT564x4NMXqDNz+Auz/mTrqdSpi/vUBXglAxGk
s2PiwNPwqIvVL3+asCL4ittiOeYEIbxwgGRdgXnCuwdmXNyJktf8niwSvlMxuvZ8
IF7kUyqS+0bD/nS+jazB+an0bsmC/W4pvgaNku4PRMzUoQsezLBm8vqFGjLGdWNE
p2cSSgEgiy/L89cKCukwdO/T2yhbVYAT5IuZj9TSQxiQhRaTWAJX5RFrxUVIImEv
nv/DAZBoovSFTrl9mS/ipuN2LqEqA/tnvbCWF8QoU9SAvERpD59PYFdhid7zLzTq
e9dMTj7KOQfJ8y8gRybMpKrMt6y6dECo7DaIQxmof3BVCw9opKwm3OPdfg9Y+KLN
TubsOKzt7ljo7u31LJ8c2DtR444HIXaUmKV5kengR57fgm46bJmlMI3NQ8ikO+qE
Y6jPd7qSmcNSte3TsciXFECoQ0obArS1r9Lmz+ylifb1ekI6NXpCABvyQ2qq134L
snVNjUHiPnjJ2WrjrXIcfI6oxIZTO/3410DPmHP4XxSKyGMTwdHwelu55rxBTzct
Xis1vTmz2LXpYO8NEeT2dREUdY3OBoade3Pvs9oH/Np96cnPDbscQoNB8ENiWsev
uasNEBV7ZPy2wBbHSzNH8Ic3+1Hii62HReTAFMlDM86UuRDRNR97AZ16oiYFKc5V
UHU2Hsg4blTBb3B9L+l6B2UlwymvGU/QgtF66lwj3A2PIOhSJRB7Tfg5lHRhE9be
doVUN647aTW8nSEcujCTayEjAd/OmNVdcIMaJZVS7hXzJCqHlZahbyYD4xtlwcbR
kfOOS//rnT87ai0j1b+62VlbT6xQF9hD0hpSQ8ANYgADBsGjMmzXGyLtv4h/me9k
ZsbWhEkEnpmtN5DCOUbECkj4Wm/RAjsRasAuW4XzfPh/hU1BwZId/O8McMoDEqRu
qG6I8ON+e0syzydkf8X4GOZ6kcF+ek/v445oCWjTbJ6hWdYOirXCKgjr8r8X81IA
BdJRUQgkeedhR6bbKX7h02rDPh1fh9iykNLMedOxB0yBr9UiDA0qM7QORRU5wgUz
q49H1yeqSKuERzDvTKtqLFHFqlKIYEzH/QVpReOZeEMWdd1uE0vUtobb+3Gl6y7Q
j5KEvBw9PXIJqL0N2HW2kvqo1M37DkEJd3zBaeB471SjFWGOGJApJ8+IZ5xnb1xh
a5k31B7GZXX+Y/rp64c+rtsaSmiEBzZlBvrPnUpvpjYJIDtKJEmgmX2sv7mJB71B
ZFCF+dTHDknhr4xF8q35ChM/5xpy3bcki7EhF9vVkfriP5+dmIWM22vbbbMrGaRi
0jGZut1/DpLR4p5Pn/yonifO8MlQwJ/7HaXjRSRm9FnYF6XqPe4A2sLxPEdacZmz
y2f5o9j+r6eVV9nIAtjC0YAgDEQuj1KtUXXfpCTqnTOQpiVYV2IFVfL9RagzwOJe
go+lfRlUwbxltghkxmSjVZ0+K/TfWMOF/tqz5MVM4RzjVhf7vY/FakRySYQg+0QA
IPEfC4rxBQXTCJw4lCJL/l0MxvbrVbVOHUCpCQnaFUI4tqQ54sxcOb1uEXiPleuv
qr7ryg3/nPuHdfE260jj1K4LLMorg4f4d3jmgywFNS7+1ezbVIcPA7qrKNXJSMuG
7wKA0JpvMLeF79fXlMg8SoW+9YvaR7+rVcWNJAVKOaHXTxTxUfMwt0DCYcwoJXB0
E+c0kACZiTyqasuEqg07cT6jsg+Bze/XbHgA4scYKo834WHkiSC4tnvNJXnSlBtk
bEFiFTHImZEEzguAPaIUWz2unBswdSgnHmmIUKF/PbRuMs9b3dPGAExDZ+fhqLo+
dzs2fvjCzgck3FDAZ4lLNmXy5bNOFc5tPCVr5nYAm2AL4aX8pm4xKrm3G/UG5aHm
fYMAncuq/xI6CaxyaVvpYbpErssd0d5ycKnwGNqkOrlYUKgMH7U4GkErAnHMhwDR
LgegZM/5vp5DLzPKq4SoEtCdxZ/rrSOmKJEqVX6oUoT/eWuKpnN/hhPdp+qk4aXI
Z5oZO59T/DRfmbfbHeJEUXlK24/WRAj4hf+C7iv67JaV+ZvI+KjExwwajYSwpnmV
VQAIpBwymRQq5J5BiklMmMJ3/humyGvG5nSZrIJJFxlc5W6jjweCw5TEIHbr9j6c
T+dGzQyb1q1WuYfsWdlub6wvWkp2R3OxhWYg0saDxCBLdOjoSODTIwR1BaCswc/c
sHHRBVw7hZv84SZiGMHE/CVE/9/SuJ76CwRNhE2ub5qVntnhTGf5KXTJyWRic6Qr
h6bmRaM68f2i0Jd4PYRyjmxfteSznfao7LTSSgMjcP+CF6w3R/frqgfY8K0kyylV
dVCUTy5POB6gYmVVewxaP3EnkHjAlQGou791MFuSNPb1a1d5+z66WBGgPpgEgQiN
h12pkPysw0240OKcgm8M5k2tZJlPVbvjmMOY3heLhHmmrOKhWv/7NNGX9wsKw5WX
hcxSJjN796YiS8bJEnYN2zKu8CaYTdp/JoE0WjVXOxaFwRFBTpPcV47RnX4kNGHE
mzCLurnKfAeZ2FlBlwpPDs1+f6WKx3tRMNvzi+Z8bA7kQ4hDct2CvJXT8eLHYZE6
Z2pvez30t72SN031V+Fzhlkj3g6Y9FzHKV7re/Jwc4NVGvMr1ks3ybRcjbj65cN8
qG2zTPUXikCQBOZYvesKVN1sgpHEhm0AjJ+GVADlT1qUUjJ5bGckZEc2Z1wSZqic
+V1NWLjqXz0m5kZ/jRjHhYTfFBPAqBPSYCDDA8rK51Vjz3GROl+hwAPQl+3a2AOB
GKpXC8Cb7eAa+fQhduX4PTnxarUR925rYOZbgW9l1c1fbZZ0L91aLIHniA9xu+ks
5D8Ed/SRqKvQM17jZ0mKjJPtss0icJMlAXl/4Jta7ayuXvgQHenXN+ZfAPw17ZRH
zv7ihZhlT6m6ImwxT+riGSkbXeLmey4xWF9fUU/PPFBJpI66AK7AfBFJzXE6Hb46
ZrrVHyBTBc9IV+Bqjq2PtBuRZCgkREBKxSemxAdmc9p292N1r/tYoWL3x5qMHSwH
ZZKMFBTxn4rCfvmIt4y76FzFDC/fIjFQr9BN2JaoqIcQnx3T28/NyBoPabLy9N5Q
VVEHoZn6vD+WzCgHxmq1gNZoEzViANsHcCC/mUef+RuhyKPfaRT1Bj2FvR9aGTtP
R8DCq7E76hMjThvKF14DdZuBJlKEG+JEAS/9sti1ZpfY2/M0P/B+lmFTTgiNaWlM
fASq2vfrDAM2FyMSE9taiKuEVizkKsffP8aCSNahPTf76XbJSppXWYmfEZyqKCdd
NnfBcjU6KUZaUhz90isQh2sLYhTJaIsVGCvLcZX/zYtnOnoHkVZxBu+BtEYgXSLP
Mm5TWsmbtL2uwPMpAsaJhtDeSYhjwrU/egzC6znZfw5+yEjYs7TvX7Z2ggUvkIQV
zTQDhmYQCv6KufnQlnD6f5fDKNDc6UVASxX8GmLnmB7pxVCBjCb0ECD+RLX18aBP
hUWilh3+NFOveb3ElhKRI8+v8xpTK1hF7cqyk1TUmXIBZFHxfm4fbrOv7qdxCl6H
Rid5tFoWeUzP1pAjSOdCYCJWtihArfGhRSqHQorsPN0ZMKvS2n+CEgVkU0K4rkJ0
2XAqGxKCtECFkxojedi/KUOlgacj8PC7PqJ+AvoDzLiEdE7tCEumOSNLWspZhBPF
3GYHDeVyIbtvzSywPZhYX5F3IreJARvT64cU8jh4SvWyYhNpIou65WInGeZjqzDP
r9KTwOa8q+zw2IPXp3r22XGKnmpFMNIrqDWiTZTe9MVTKqJMWZI8Mh3V0AdTWkLU
oUZhMmc1U2SpEHy2y+XZRyheIJEK4qxutOTzkxfuLWUj8yrg+0sG2/Vl2UKokxOE
Avl83VmQ7k2QP2EzIyZBpwEfaYMGqkK31x8FYI0kgZ6bBGYz3Xi7vfC6WAMNDWmF
tK0iK+TmQ+Nb+2H45oSs1VuS3eRBPBpWtsL4hkJ9BRFswpZ/wV5rUTtHJOjzjnZg
kStmL34cFArOKwMPC+sxIDIFd9yuQLRydJwtyU+q54QngIw3f7KP2pZWfSSBuduy
IksEoan7smk+YCiF0NlSN2+AcN+X0CBTbgPlak3sFyPH5eMQ8DNnCrJJ7BJRY93X
KNfQCSLC+N8uINPU7I3ixfh2Z1RBnyaGj52RwZ32+GYSyIY0rQRBFth54BRZCf+m
ev6Vd63ucWTv64EQbpYqXfVPUUB+HVKi9Mb/8bBtxTEhlRSgaoITzwsm1EQuqbk2
zF9haZyjmcqpm4IH1Edt+XV6MUnrEliVUTwvviXYhYb6sA5Y93WmTrS3M4nQheOF
gxojEC7LI+YXnDMW2KOyy/lI4VZlqazTeU7F3WDP2REVqdtIGalw4vgjuQYMBFgA
RWb8UHRaoe6oC9peDbQqRPXtBsUxtQ0st+9SL5NiaWgyUkD3IKc11KDdNec7J6od
H1LnP6F2w7CqVLBZ2ZfG92aAIkBpbhG2osif0YFB2aR0D5m1d8qtntYcUNWcDVju
T/jOsHpmScE5rk2Gh6osiV72/hUe0C6IxrlNjtH5BuW4zoAmn/Bb7egqxOUZHrqB
7T3P4RRZmgY43tuTZYvq0lbysPBUzaz0kczzoOGARlXLIP0qjipqYGjEJ+S+EH0U
XeZolHPndK2J3RdZ9SttX/5vd9lVsKb/QHUVKNOUPY2W5lvwnTiM1AJPC1tnshyR
ZyMKQxKj+e0iA0n67OW71pbsZIuahkJrCpx2fkVM2Amz+DVOp6a518ZZ5j3Gi+pe
6UJ0KRxsdA+Ebda3dW+URniIaourBKu/WW2vu7xAfvx+u2+QLNAfvPdVd+bf0lnM
zDab5p2vQCLRmaI9EvFWq16A2zoggsll1cM0B/BuD5UZ8zVkvaVHXbTId4McwYzg
M78bucJY3WgJ2PRoqsjNCSe5d7/yVR/qRYBFMjxHF8VbqV9ydFYtJj4yq9hHSr0q
UX6pkg8Kd64Br0xOvO/WMjfRPpX1FVbbBgnhjBMWT2pN0ppP5pz+sxtyWoF1K6eK
lSE4goVriQh6K5c6jr9OcnG4pXXABcnaaYfC0bi40GG+KrXA+X4CwE598lYNQfvt
keEy1FDEciQyDVYcdYI33W7WEBIwboNWvUKRodwdLzDSzYYXTmA9vzjwdhQ0KwA4
1Rl+73WkkUz7RVfo0i21AklCnfo+QdBdxtOf9ay8p3uyp0SKDdxTUXxi/ryTgYok
b26hXwyKvTOhAsqloyVbmhZY5D/mwDIkNVYeZJVNamYkgQxUhIcs8m2MoA5uRXIh
nYXVo7UcxStCvAEnUdv5f/WYm2XomudZXK6KC3JBG1KkCwLjMd6SbLFHC4MXqbkj
NOGwMpnLAJhSSGCZoEBlpDEO8TXEbsGFwlCkgz0wkOlUgJqWWeoVpM9QqYR6KqKc
ZzZ7eDgiLRHI6OBE6GI01KtFqi61/aU7A3ym4CNw5r7Pjst+cZ5/lx4mFl8nT8YK
5NSMV8z/6LF7SKV+srsaJ36NTfpBIckoAPqzEbdsXzdyjtwJsYlIlMXrOk0IyZHq
Sc6axS4vziTCP/ywyciskxJXaMXLz0LUaAL8+SkBjLMh6M8HuV4ZIBegoAa2Z1eC
djDKrrdCg42I+9gSlvPgiMnAnGi7McLTKOcvt4IEh/+S41yEkUWQt9f8cke2VHkI
vdmG2M8Y8w2Amux4G8ogCgTv/9puRfrQgm4GQKpEAQM0pyPuT1Z5KMapTQwqF42Z
m1kn2Gcm6kZaTpr2VnYS84Al4cs1e+mjpnTiR6L3b2XjjEPYW+m7pbeefjmtTZUx
1F2Fivy/PHZJrd+3qDnESj/WC6iF6Dftqx2WledhUAQLD3h0P8jSXJ1WbGDj8Z/2
oh7ENDwpWA/nC/FswTfwUK02Ft0a0D6MuE/2sFLRTqWZd5QPleEpy6hqVNe36UHy
TFteeORpjFRvpbNe4WHdz8prxRAYSrODJnH9eb66lqpxSFrcK5ujBrA4fGNABto/
1mkd8Hq0HOOe4NSbc/nwXu5I24Nx7P9yUAOPbQjy+NA87kL/hsW0nnQz5NMXmIHh
bLgwQhXET9SApyOpZRN8nmRGHgwMrQ7iqXWO14KkMNpP9ncwTMvUfkynhWiYp6oD
Cgh2kGYJaaa2hm349dUOzrUiBosCoXC4UDt2r0xZw1kQpkhIotmVa6zNiUSgvYl2
OOi4+Oc18sfoP1UHaHKtDclgbL+jckIC/xhXG4XG0ciQQAntL7UAXJA9tvdJBGat
GglategNdbaZ9wkXcUdVxDUE8KzhcPkN2eKjxvNGb4pYU4qgZfmdPB/JO9d4DzUP
zuApt2QalJbrMYWep6vI2YPkqM0XUGnkmCtw75w/Fd9q3UgooFg3+0YRgB4onCy8
5ZQNaxePWzuoJUaifmVwHDrgZjdsLV8v3gGLSRcqOC1Mu/QzuzRKVaEs4uVDHydT
rlA6uggoF8FoIhaSPxTobyXaa/JQ5NAeqjgdUgk76+0TWWuoSZY5vLU+cPlZWK32
JFaFr9nVIuGID8mmY2cVx7RSLMJ91iMeL5Q8yUfG/0+ULOsGf8UDQJHEAYe6eaj7
aqnacqmOu+afZi4+Sef/ftfmvH1te3LpkyCzQVHG6cG7iU3WenxpUK1dLKmIFZfm
B3pM801MqcTw8Ysbiphom91epdfPvn5dxf84Y7rYCd8V8CyeMduuz6dOXU8/AYBr
5BRdGltmBSH+2jlDJVTt07cUOIh8jvl/X+R0yhEvqQEJuK2zB2hszFodMNpVLdmC
Dy7OzwsSTuWMJw/p0YSZ2EUIT2UmSNFU+6UxnUmeWfe0hOMUmOldgV3ST+GLL8O8
GOSgCUzCs7c++ATYywBG3neJK7nBJIH4Gf3bbQak5dQOgalcy9ZwBYOeUEsxOlMD
Npw/J+/Qt23IZHWEa/SoSxS62wRQBInxYIRFTQqQSHeSQdV2wR9kSH7hiJ37a+/V
ome4OVDzOXZQR/7SnUU1FPh7RvWW7cyFvse4OnPzEw3b4zSXrFJ1x18EDRtq8Asc
4TRvhl6U+Cuw7Iip51OpSkQa7xdx/uUrsKMDpnBnX0AfsxaacAb/tCmrlcafBSjA
30GHaQGxok0r6vXL8uZmsaQUzbaiXqu2fa28QjNnSRcTGG2yi9NL8AXR9Mqj6rEN
rKMWRUTw2PpnLa29Tu5FmgCh9ssHrZtB5dBchPT/x8beI4vAkwfPrZiAUSrHZytd
5kvvZBQ+AHc+VWoHkazZR4dlQArHuEvzkuSGDsS+6bgjL67MhdKSd0geGzkeFN4x
40DxrflWjRsX/K7s3jFzgo7zfk1QFlFFJHM8PuRCq8+P1qPw+snEUA3byTvxpSyY
E9NgB30+kEqilPfxeiOSgOU3y0dyRrYEl6EX2g1Rt4j8DlP8wvHXoQBJAzH3JMEb
/Ci0JbswzBwTsTCPeNWylk0bqUMoAB/wdY9x7bpYQgGYd4OD+q/vap772/NodG0v
uKGLb175N8MGoSo1r3O0BOGMF17tTU0E6pXT68AovSZ/mjX9ywa+hdQGY4WFFPGv
S0sqYZ3rFz4mqKbDVAdPZBwOa8xar9rmf2+lerYhN12bZtFS7o9btqCns8ULDSN6
m4dH/sw+8g6V5/3nZbfJ5PHAUGRugJNbM/fSPATbH9WugWxNrWOvh1Ew1FxwCSjK
1DTzoXmMApX02tY12S2FwWSOL6cdIQ2qQfjOIga6rlgMIcKfxDb/oVVL+9r+mzkn
i+ON9/KJT3BalNw4X0Iml5mhm0w+FqQ92sIwnoOOekXqUZiLAx5rayDXIUT93ka2
c7NhBZqIQaSAI9bMbHInIFnCgWpXm5ckuHtqsed7f7ip0cinFtvoPiJFP1aGDCvR
AEGDDClYlg/qI94ic3hCFtahWqxgwDUoC1LpZVTHHdwP94YXgBwXj5D2KJAq7hXq
btScraE8uVQRDnWUKfZamYZt0hkZ5+Y/y7MAMQt23Fo5iUdXKrnF2s12pzwiWm7X
eiHpkmn13/NRclu7d9g4j0z/U9fxfbcwUCDHLtSLjgNe5RoVpYF5dFWeQZP+gQWA
Ltpp+Z15CL2Qqi0Jq3np0pnQ2tjj6v7olbRPZRCOq1BRqxVtbW3S1uuCQsJhgwZo
aquhiZP66NvFeGIdLLrwE7jC/WjjXIna+UE/NA+ZffAXTcdnapUiAAyMGhkg+73I
d6a88Bmy28FP9zfKcG60ye9Y9Z8U0DzUFgrr684tM7Ko+jLF9/pItE94nP0goeQp
7HPZxivNazpl39jj7fgu+3SGddyqUPNjAK67D5IWUWTSnlpbzWPoO9fPkhTU7Sgt
NJl64ZcSf6B1n920aycXXPuZIfPeuE46bdCr91hIvrMsHzu9CXH1QS7XP/Z9n0og
BzQ0I84t6eMv8K1bPXV0ZB0KONMl+HWdCAPjiRlKflkXD30b9yzF1j+5svp1+79P
PH9VCSyoo/4M2Y9DsM9sS4g8WtOsGM1C3f7ZureUn4WHw0dAY7blX4Lq0SHc7URl
YrrbL/fDEHh6bq8jwbdBkO9/M3OLA0yOOmslnhoDl4vHiajSXjnnD1L8OmUG/Czc
lVULjH6lWm0tBoctgbQR7JOJeNYz/RuwDiTSkuDPKHxDKvkwrg5MomzPCcaR5Ims
g6iwq6iZJxpMe55EedU1xFtnzqRM4HfcTDX+8yKbK6YrmPt8tPxd9FSyIlpKq01n
ne6tiLmr0H/uK8wVqF8o2OBrA1IbKUlo25Sb8sRse880cgzzL8pYSwneWhom3Pr3
9J66aAJdJ8hFa8/rd/E3P/dWIrHNFHeUsUglnGVIsUcUxCjGPQI3UJCMUdWE/2RD
ZerxBn7Vixs3+Rouc9BC53yOgtbl9caC6Z0AdW/MdW8j/gVbJQX62Utz4spIJexz
qScd/QLqEFU/1J1S/+3FpMOtirRRoKvlrVfaEHo5dk6+mpueGjsStUjY473L8/FG
ZIbbVy7TJZrhwdWJT0xktb7/DiDfqOTd89KToBMsnjuJ81Ej70t2FR64MAwgqXlX
cYKtd8rEiOUruedUPxg0Rb0r9GqnnpSUgAXagOC7E/+ruX77Oc/qCXZjqTM9Hrk4
stKjspzIaDZLzkrNz/cWgldxkPX3hF5fVAyHYHh6xqdpEuqBRTLhhtMiyXI7lenR
sToASlITzy0cDqe7XTuB1gfNhTuYobmtVicBY7YG7enyg43WvUgpZyjvQFNjUHUA
efofHph5KLEiPPhB2bh+E12IGW3XjqcKR0skZDRuRvFMMlL64ziIcdBOHG2peRnv
x8mSrNWV6pibAFADJ4aa2oeIv5IgMzWJxf52h3VFczvUW45SeKjEm9spmc92YxSQ
aiaDzhEeTqRffWWRN3sl5Ptfk+AERV7b6HEJ5GQUNjsMe9oj+gSLNVDpmUo6eRyq
3e4uJRFmh7CzxtQ818ZAa6W4UeNUqhJTE49vYyoVDdJnC7BMlMTyp4NCWPjP38r4
ngKBsheXCm7UYJebeYmeax5w5qattLzRpESRhBpIq9FQyGbu6T2Y9HJjiG7bOYXG
gwv5JuuVwrmyhdxcUc4q2DdKQ/YqeEL7C/TUtb5X81ZzXZKNhS46xKkJXYqNBK5k
ErIdFXmJgSc4jWUg+sHMPWSJgB31wXi9tSKg/ZCHNu5PHxEtckwQZ7qImWOQ5tpj
P7544Lz2i8Sjr9E0omeFxAnjxcGqr/1zmBcowisKLkDgvGGTiiEywXAGjeBvvoaI
Kv1OJCmmfJ+GMpjVM/7pHT1aytNMPGWaeEnY+6pve4mbsS8j4l3NnmYqmcAxkz0Q
Nl5VQpYKwF3S0AUlAdq3O6TnSx3f89J3SJYLlOh9fYXtsqzdxBtVoBJ4AA3LmTjL
XAq1hMeF05r+VsxkT3rqYA49Z4a4GpzFRIuzVkGA3MVjAwJnAiT82lu/YMBh6zXJ
J3//D8TQl7NM606hlg53LrntkfGjmccGpCisc6iI31rfB7rQqHZAQxz3t2+AugiG
yZXjqb+s7Pihib9LaFle5cWGRkwCgzxGSCNZ8vgW6ZJgCITlikH/waUixzOzK1yi
9BvljCHdroAKnTvyPv1ZbcAIzRTV7/qbinrnCxwYSNwjTcBas6dTQLWTg80xUfsa
wDUTf18oIh8NARglkyx+1JhaoGqdgWqgGU8UwWlPFl/NnGIAilWimrH7LfLgladx
+3zIcRyH27RMi2hJIYPVJqBTJA8j7bte2CMPEPVgg2oa0fhTcWGvIDcvIH0IxxdK
NxYmBrdnGNOJuyufejCOjB38zD+DRDJJhZFofIkIeV9Xu6AQzu4EbfFKvHgWmxIy
GGNJAgGjk91tNuJJuog6kjMGXcQbzcc8oftAFno2t4XB185V+8kFbEWegyZ1QSLn
0Pb8wAiPerR+FSLGtCyXjz9tq9JvLY3eD5qqPcHRcC5PGvSvLlozCf7RDmX875h5
`protect END_PROTECTED
