`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xPFWYsX7N17d0BvyZE1eSUZWVP3DVS06XWff6bQrvSP5bWX1765vtiSTLJ+nWpP1
Jrdh77XWTSZr+kJkTTKOLEwbmxnua59PHe6ldabkllCGS3YxJFIYjPzQhx6QiFKi
e0QZ9jgiKAygIWwhCkUE/zQmfJxdyZ58RfyEbgwzGAWxfEE2cIfJBh/ksVu2LHdG
FQhoP8o4QJ6Agx/u79vNt2rVTZIZrcIX4++LkQHl1HrqpXxrIIp+P0Kpe3dkKkiX
XoZBPzi4+hiFsjJINlIVWfhaqAXYwix8KtQFKTv7wP8sMKlwxxu9KtBg3H0g/LyM
faD51zIWbYDD/Sf4iSFrmixnyVEnKVMaDb5EMEcsuFhUYQWtdbeLuWtXxhC5XMic
54iHyAARNdHNgYK0cc2tC5RQ4r1SkvdD+/8w2u/yVozikKC5KhZMmAVBcOuJRqyG
prXQknU8njt1nqHCipqV+2+PcR4eb5QupWeraj3hJg5zY4GCcO1UsbcIymA5CXQ8
ABTSvz9D62ofm4Px0i1nnrwrgFkaAG2lQqtDMFgyfqRq4ylySY7JWfY7SRsAmwdh
ArjtUOX53nLVjraVu6+FlMk3pOgi/DZ2oyDZzjZwVgvJBx7uD5DDPwXKoFWKVY2I
jEjCezH52VgGIc6GksEwdIshy1F/KetWjJPWLozn2W9zNNPmqr95/Hk4KMOgo/79
n6nZT/dInYcI0ddYs30Z+77FQNFeps4qSGn75N7kk0YtwMYDFRqHx2EOLlY+xehW
JnFV7qfiWjX/kgVWZa1HLhjkqSNif8mspN6RF+fuILrKnV1VxTpwjsJR+Yr2q/ym
vAfYzyuS7vnR5tZZLOmb7/HRg6uK2RHvVN1qccqW7u5NMMkvDC3LlTBIzxRxFHsX
w3MYHs8EuUO/UXVcwWQB99tvRcgtcXb8VlqsjldmYwJGXzhDqtS32CaDNFz6PKP+
b5yEzWT1KkUUND/8bsm5xeVFLVlbYersvRMwpuorUSG21uFq56hD/nTkHifmcDot
8LFyd3FX8Z9BUWzBpsmqu29zzpzsjlAeJ3BpfLyyzOEKmfXxvjpWAaai0uWh3Nlu
nlyz8zkN3ClfqVXLOX1TzA==
`protect END_PROTECTED
