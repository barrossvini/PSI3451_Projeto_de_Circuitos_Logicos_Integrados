`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dGjTECwGBtSopwWRHzI7ix2b6+FSybJgnmEFT4L3fgduOawWQiDhpHTRz2atpqvF
uNPF2382lSghe0T+8OEpNJ2ADFzfLQ+wvLyJ5L5TdeF663Pr8kFprZv7dJlHYOFm
azWS+8DRPwrXKmuOxcNY/wzAS8RAB999w45XGWYb0ax9h4eo+r8f7JWiD2pbZePg
/wiqm0A7fg5b57Tx5KlxexsIsd/45swTtMaIlpels5iQyg01qEZqHeGaYecaNo1F
TaVmo2Fcobm7ZvhSfuqxa6MZQSu6CeAcFgLfo1ilGqJ1RPr3dpOoHW8hO8QwcpIe
kjItiz8Wu5nAriXje8yZo0nT0lg9KCdzEuT9fxIL0xq97lFJZjjpLdN4RRaDoPrl
4QknZiCq/ErNL/MlB+MYjBAXEwxJi50xsBcAqjX0WEmHH8WUyrX1JY0SBkrg+CZE
f1vOGNn+l4fGIvcvdrL98rTTx+I0gtMwo9L8xG39tk684pY3aOjAcJrErFEFI7DU
ftF8+tY5X/YWrp4nYJVcGTaqJhEiEi4LcJPswV47oHJDKenlI2MOLLR3KWBL5+fY
A7Ur1YB1hWYjkpUS0a9nl2RShVy9MsWHikrpbTG6hSuBGOfttuIBrX50QMLyPlrN
YDiMyNnNgrbLNWI54LVe7ogT6Fn5ofrZqpl7157+K9eNhKz2Ks9MR8BWZ3nrBGpI
OOvqOJForXeUIVmEpdptiNLVz2lgD9XWdfG6wPnNjy1eS9p1dH8OkWv5xUvYEvfh
MC4Cn5gveQqmZDwy5sh6zk4QFutR+79iFfBE9iSepAz+feyMkzfN61zyBhhJLiU1
YmVtliXGaiSFZyue3ynoynXumfvCxG/iVGeudJ7TATBckUikGGhmVL8daLC3g433
hppbb0Yceih8/5ZIbne/y8Rsdy9sb3vlbWIoMWFHMimTlv7DJhucHLRouRPDkzQM
bY5SKR/i7Khn+/HFEDH3RXXtMRY8392G56K6Z7YM9aui5PyTPOMmCQM4j9CJsw+w
2art7/ERtdXIo/U6O8dSfh4SRK5x3Kxq+1QppFUKQVJgt10SaXllkXp+wVgFERIh
bHC1G4OtVT07PuPJu7lmsCsmnR9rdcyDCfM+qfjhzVqlCY3koXaL3Xnf5RnQcNnW
nmTsggGye0hG8I6FsEUV47ozdj7yaeezTDOyv6QnMVC1p7H7BBpJkEeb+yfgPZYR
tlDsFKzCUen8wBHwkiIT8Qr7GkTuPmADOboqDKyZkMKNJvlc9zvxqymKgTMKhTWu
hhJh4XA6V5Uqyo9Xt001kFzsNlyzkyhWZ88A297vOwALAvaxG/zFkPy8GWopAN6S
Si4CWnqLOxTSwgyermZQYbshf42LVwBupE9KJEmBLJf4IJ9I8AmtZTruZaRXyL6n
ODWNttAVCIOqLQ8E9BXoR+bAw9+i+uM32cKLbtvybALZn2C91ym6dBKfI8RfOzo6
loh/FvPSABg2xoo7YavkVVUkZxgFd52VMrSl34khrKT82yoh/hpsqFJ3Fd301tGg
lkuhm4ei5BTwjFU4iH7URXnmE8WlY1APLwQQL6GZ1TG0gKijNHfY+SGol6e/vk6I
l/AMQkzpX7o1NBAqmFwPp7Y28Fa2f4ag35hwgJpuFYtaqGUajyz/ar4JAYGmhXFQ
4Rgue2MFvHjzV6/rDjt/dXzOnCxODXUGoATnd14vYDstlvlLDoUIh7Pfru4iCCXf
CwyuOwtMya0EezliB2ZLYC5B2tk7WSoK1ux1yTL5p7LrtM3GjFk6HKxR74DBCDKq
XPW5JGdhtXrhFDfXCcK4mvy2Pk9zDVgw76yBKNm1bISrv2OH77Kb+x206VTuoQpr
25M5vmZE+wavIe2maSmz6xcOtfjliLumW3dQWbnga21K7OZOhXa517wJigTSty8N
ykU16jHlXtUJ0oZ2fzPwpXLZfJwr4G5FzV043cw1do5ql9VrNtx1/aTgkUxKovbs
5W6xAxIT7XFi9WVQWIOHJnAvA3SJ4L0d5HcKc4Oq6SbxsqN/zcsfW0d4iYAO9tdU
wv3kzLdZmWZD3aJMQZRRXCQ6hOprZgkOe4l7OxQETyQYVBISdW/I930TuuiF4+LN
kXEbgX/MP2b0L/qNDnDeokhOyV8+4LiIFnfuQs60efM4N3urttX22Z3E/eI/8Rg1
VKwMgydSmzLi73YH1ar5c1+XOv+rgv0PNJX8RjN4TyVvXX+uTNTPeUC9ODZwHH2x
70Ab8NOI9jKbxP5fR1kQWKC2MnlRR1s63XBPrH1Ata8YcRTqP2UXxfxdyD77kdH8
Ma0uzP7OHJDHpcChuom4J0kU0wIjj8ahrlwDfkGuZy4qaNI5UdMB2+0/5Y/H1c2z
`protect END_PROTECTED
