`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XFSlIesUDyRgYQDNITUifmgy8i8N4xp9RwdmzPKXxIVBefrTjZr2DgvsG7yRfley
bYyvqGp7Y8kZiguB/hvBOIegeaMDCn/Ct9qi5ZW0idEOQI3d9uy33T6WqYBfskJN
M3sK8PZXepvibH7OjgBnj80835qnYADnj15OF0dfT3Paj4aInIvKOLElNzurZUcy
Sq2RY/b4VLbZ6tq1DhMpdbwLv93Mx9wTrAhlqp3KUcXufzp0k5ovhbHyMtD9hAbJ
V5r4PL3ui+dHeMumzj3jTdLe6XmtvhpwUcSpF4jF9NmFeLkUFHhJxnPJZ12DAnni
XT1TgyW/8vv0GxIA4hdWPXf6076eVOqBEki2a2p8LheNohBdCqk26cCi7ngydv0f
W84nWHWnTybis76BW2cvPPluKnXa1AnxLIw5U3PN7fWKJc4J/H08yW3r3miZXV/1
9kNcDo2XMNZJ6IY3P6dfTAcG+X0P9izz9rp8BhbClvzZidGqbT5tCXKjR8/i8JMm
R07BkjWVOSN/XDKdJxySj4oDLCICrjATMHIQGyuEa1aHtjXmPmYJ6240fI7o9Gqh
mAv62/tBMIf1IOxQYC1nkS+EhOv7gA5qrAvTmryTmh18fMmql2x9tW7x3waI8SKI
3LBFErZtrU1eMKl4T7sPUspUwilegmLZyNl6D18q9HmIrq3IT/qF1KSoa+SpMtpX
PtvlvOMAs3+2W3nVAguTNJElvj9WDb26OCTPjm6l6eEizotqEBOm8WDTjXkyarNv
DMk20UQLEuXLvCw/njX9h51YKok94x3ZyeaVvb+XckL9TC0nuWiJRuOTA/y+J4UT
8sYyZ0SfHutyVi3hHcjPoT5RE91qxlJntifqcoFojGlU8s/Q+ZzdkP+SLpcigqzK
laXUPhTht0Ky/nrYC0sWS5Fy3yDV1lFmtamzAkjWIZcOv+6ai4MK1gHzkPemPNwn
1Av+gbNmFmVHCeZxrLJVlquwWJ9ac/auanjA9YX71Ec5WpXKlHj25+cz+GvSj/60
vERWkpOfMkUJ9FmDeGDzIeOyMAgqevYRIejJMCtDfspeIKKAlGunSTcjbzu7Ve3O
G5s1dL3nmlbUqtTlppDsjfn8ZVSrRqzwHR4zeKmkPj7npWgShA8ORqwAMsvKGsMz
`protect END_PROTECTED
