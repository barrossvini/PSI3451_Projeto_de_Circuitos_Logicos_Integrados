`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GwedXJO2UOY4vOE1UkoszjS/bcx9PvspDKvr+ifdI7gn5nA5DUF6usTAq9P1pA2S
PZRgDH0vqCJqZXQsgDePxOBWU10NjQt9M1n+8ZTWadH22Pb7qwQby/uvn5QT3H5N
q/oQtFCv/rCLYDgGz+5YP9LkDgFwx+DNQ+8QZWgN4kkKXlY7h4MdiuztYiP9ovE5
iYtkbeekRN/0HJa4hime6fOWywEZllqcNiEUCWPjOYcXvz4LVn+6XbdjuU/Crntf
PZLI5zFCn7G8yuL1lf3UGyG9ifI8UhhHV7/eAmZiB+YiezQYmxHgBCorfippfdxK
iFYL7aW9aEtp+8iI+Dx81NwaDNEjkcq3Gvw3XAxWByohG6Kugcw6vCGR1iaSy72D
0fTCXp7+DNLNsHJQhWR40vGV+FC5bN2A9i6x4UTUrqqzjgMAqV7ZpiMza5jJieMr
ZRBRIlkgrNkg0rtsKScOKynjTv187s/3T/JX/6eLuIylTqMQXwlSoGJ7uWIrg66w
H01TXoKN5MXSz6TfHRP3W+H7ybLmKSN3FXp03oiLloj+xeLBBm26sBl71RA0td2V
XXIAUiC78koA4NH1BztjUWldtW09z6SpbxhGdFQ2dz00zk4oV4+6dEQAp79diQg2
gajhPMzwIErC1gMqVpND+KD3BxEZC6YeuiVWiV2t/Kqqu/BLF6vSmDAQGQ+5uuNU
mHNj0TQNpFesrf+iBU3P+h1Y0oRegMG9ZOpMp3bHGFpW/n7Pk83IAAisrSabHPbm
xnUikDJH6HMh2f4Zrt1YqEyNjFUJFjzz456yl7/bwW2PHF/H2wyPgeNTl0Z2E+Qf
qWRXLRqRyXCVEmJrreReEvWFaA24hb56TphxOLFFGecHBhJSxw6iogtkrOqvYRo+
EvsAG4WktFGxvbA0wLUv006Ijm2O0AOBIJtBxOjn6gs73ylpHaUJmwfTm7EcEq8G
Vwf2SuY/2kgOIS/2MZH0vuFMFYYmLsCasZuG32yjGWkNNlCaxT4tjbU5djnTMwDN
8ACsBoCZMTFeZddHGK/apv47G3x2fE81fUW8iLZby2zh2UGnE2RcthWGJf9ie7Je
qRcuJq2Rucg6Jmym7kZ7do1NrjyIZ2XQ/LxDOG8fGtxJtFojhUO0A8xca4YRC6JI
lbHLMGI5VUJQIY/273l96P6nkf8ib1gvIXmG2VNl71yFO0swjpIQdWxz8jMgOist
fEqhWEjiINKMdKTHbVNd13logjlfbKbePMC1QZOYC/I4aYU27i1dDStak3YapjdJ
NeUFhjTSJIqc83pAtE3pRfMCq4SPjgiOx0W4KYLQH5gn76ram3oSomUJqYlxE3Zc
3iZeh/U3Uqc0BHm1x4F8lTzNJupQvF7VrcoQfoVQVIefLtC3fZPm44egWrLtsM/V
y1l2KYJYUic3UAFXiBjdY5/GdFjDdhXz87NFrKJvB6CXlIeqMRgKEzmmXgK1AWn/
vCgyKAw26v4aAFVSb37uCOZCaytAQVHJGAqiMBt1hSnk1FSpl77+E8KImIWOJxLG
wfcFBFr9fyfDwwDYG8F5nioMG1vOvlaTADGGp0g5iU1WElv+3U4QbZUwwC+h1u46
mRkjnk8R38P1p9EoZ9P60s0FJtBO45/5O8RRLbMS1Apzs/5IZ97IjEytLkTpFpvU
EK2U5hrjkv4RTF3VZzD6NvaHy3cJiGt3JmqEOdXEbHKeFBi4+wnWIaaysJm/c8/o
inXMrH9WyTkmdyGm6kVgV5LU27vUzZygjkFyXyTVkGf3o5Z96WafJl4tuP1oOQqZ
B0youMnEMjAkEGjaxABelC8GZnFnCZnH57JJYL6z+yGhC+adAkMB4AhN4L8w8Gd8
m2hij5hWeSTu2iCOU9Kcm8REv6dQIokY5czJxuUiaatogrMBu1D6GF/7RQg/4KSD
zlWmcd5Bv/3e5IZkw7GJXO3EupgJdWWptGRHdki2uh3EBt2mh6bNvUncpKYNDcwy
TdNW/WSskkEul6U3dTuTXmqP0SwHbxkcoHSLKjtZ3bHYbPyYbxu/b0XT2OYfqMzL
RujIcaEmZ/MXKsYi9mA6x9o5LZxcjo9PNtYiYaAOfzuQCw3CZ3qPdjNPAOm4ZuV4
IX2d7iJafGVmUe7fF7x4ZnmEq49Zf6HbzqfWuPbX4uzdoBBLtFoeETiS2NCzzmbq
Tgn8F8kns6ucFGFU6+xigCuCV3JrLsp4IK6ZVJq5MOMxVW/U1ulebNAAhbGNA2/J
Kj3gKbkGAUVjIRotpZSQTPOa7seGl6hK5RMYNaewMURWZXSe+nTNRIvQ634cZBbc
gqdWM7KfMPGmWfJ9/R2YAyHV31gbkH6MDsbUrwaBEvVHFKdAUYUn2TsTQ4WFJloc
WCDeze7sYFWuq99BLYkk9Q3s+G+3nvRGDXngPbKa/XyCeY3G8p0ykVJrCODpI2O4
ClfTtIyphv3wAzAZkKO5zIHyV/81El8Kg/4q3T0B7CSI0uhATl1G3KtzEQNV6zqA
kEMYCTg0j63WYJOD5cupn88CyWKR3n05yfCWPuK6V9GPZZCydkuyIo0DRAHKEc8a
Pm4qIaNfdgGVuHkGOiEaXhMcW2PGb5LDMKWnHO8Vfhke/HCoihwKFDEKCc299OYC
Ww0BCehI4rVVD1ByQ8B5nQ==
`protect END_PROTECTED
