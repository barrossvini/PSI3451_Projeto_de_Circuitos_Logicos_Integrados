`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Emugw0nRLP+f29ectrGlcpktUHuV8KgwWlfgXYW0RRyVnECC+B1umwt0pMoUcrMW
8QH4LevvHF29HD+RbBYODr9ds60OiM/8fDNpdhBQIv3JuOypmQCa2ECF6aUeKlqt
aqyHXlGE0+/82ybsIi9ksp3qkQwBO4G3sGrtUQ+HulQRmBOr8kH8IDG11ou7WGzN
TsRgoXw7gg1Rsqs77CIJsF08kUz79xbXQ2Saa4BXM7YyD8/wlYuUPwCpRWrIcMzC
BKJicqUjwX6WY5WkB9Jd1EwFJikpngryIYC3zVEzzo5bdI1GhmaGvKCqbpMNpZQk
dFZjQQFyTDlbFSyCIIjxPR4WNja0W0BBsvbt1d3GdzS4ZoRJR4kILQAE76Bj3rhr
UaT4TDKnYSBeoM6EfJWq2l/Po3Vb48R+qARBPUIOexD5UGid7eqJoExaHO9zPX1N
9MB/UuafjHJjdaFtgva97+DJq5Y47bQDJrLvhQkuMRkOWJ6Zge4OpPiM2e0Yxu8M
fnkiXjRRNonamKK5DqqG+izCvOmLJo0OB3CaVX+RIqI2PL22nvkFebfHBmn8xuLy
vETpprBlSOaRYxLHR8msFVm39GPMO2jgPxKLuvMO7OG2WcuKp//SRCNqCQo3KMUL
lz2gvQSGXlC60aZ8f7Xiq7/9WAHCl3BS4E9FSR3UYC72jRkpWKOrAsxCsE7rAnNq
osDB3Zm1CeVQBiIWHylmoOhVGQZknDYuD2jmK+FIz9/WByJwbX05lbEwlTvcs6Mr
skZuUH4EiBkP1oztUmtncwtbwikJYp0YcPd80M8reJC9hmm0uGKa14YUWz49KqlI
g0X62k7907NKh2CofXgc9w+pLWQtuOa3wyMAcw4ibXMydbDHHo4OF2XiKbSqvLGB
OFCYWIov+78pWkEL5sVdDbTCYR5PSOy8hL05KI/3XfcI6UEnN2HXh/aqmeocYlfL
WXwArKshAG41kmdl0UT76o98846mRYsMiZaEoiATL8TJK9IQio7XrDdk3KewpWBO
l8JFa60Bao6KfSNDrmNvsYCNftSdGImH9LnOLVtZHUdJm22vPO2B0nFj1Uhob4+r
pWTFTZj0xwigPDXkmu6BK9LSZ/xjqYhwRuHFQuWoPXPYoib/cUhxrQ07fhRvJKGa
gm9X8RQvLvxFo4l+R1LKIg03ckkem8l80izUNw0Ldwvo582JDtqa/Zt0V2AD1g7r
2xvSj3ar/SpSIocMEQSnoH9j7v96EWYb3hdYz36v9/GA2RTWe8vVMoW9hkvuq9rX
LT6jtphLtN895s4C49nOxHd84Ci1PHhf2ePEk1xAu9vZyrjLi0b6fJkw4hPZwxkh
HS9j3ma32S3g8eSfrsVPGTKkh6HUDszJGVn+3QQp/JwJt/Avm3ePsxDk3RpVHb32
XMFY4d4fr46ilyB0wCBXcMmbibv8QhaHExX+MQfa9XzuM2Laqw9o7Sn3LXXHSa7k
J8i6mKMDpMecOmpJY+Osoi4YxEtm2l5+L0sqNfwUrnT6wT1x5jOSzroNa6EU+xy+
+VF44+tMxaDPmPzsKjsRvMq4HajERQMJ4hz3FsvuoWBz3+GMI/akErMvhaP+GS72
pXK7l1zOn1bOgMb/F2DkF0e6FmKHnW10EPhY/zaNyavyyvRauEBBIvyuTczbh5ar
Av3vFItTfk8KIHxWOb/WoRldwYboWEFRr2Y12pYgsvVR0OBSJjyy9i4+CSUp3HWF
tsCmGxhrYNKHGP3wpkXREvzceRi1y7j4q/wjZ7WxOZTED7Vo7IVPq+RbxRMt2L//
6+xuG/vQfyzn74eumzKhQddkslyjov0jfmkCUFzY46ncvwIxB6YwGduTq+eTiKA5
nwae7JDIZMt6fpXS/2w9a7oBl0OoaaoWJmcMdnDLeESCFHW+lGRX4cv81i5LIn3v
SVeTXCWXxa1Z1lW+CAzRkqdpfR/IEDBX8rHUDy7uNRlyfFeF2e+6pk32Hb6WPidd
oaMe6nkl67KSS1jFa0twQr8hlT+CPD/oxuHs73jQpUuL2pBBDf7AlubXZ+09YkC0
2JuZsLQgy3CGyNWzxg44vz4/P61JKDtqcyhDtdUfzVQLZHQopeJ7ZlhmJkGrVQN3
AmacEIdWufjtW/K/7ggURyiSU2h4NaQAvxacE8wcxDERMkhwAY/PmhU/iBgoph55
5V98TohJnOVdvXLy6uoQqimJSVQfMrOIanrekN26Tmm/hCifrz3zhRLjFbwtTTbL
hPsSJ7LDiymh3SMXT1S4tglsL4PmB+odCC+tfnMiRem+y/GWx/nz0mXY0NlWiHbe
/z6A1NZnZ1rPbehVFhU8YOpicoqY/p+pmoVQpeeNzS4M/StpvTeOrZ/lVhus7FZr
DJgpJUBBdV5jAR4fbiaE6v51VtwWd1JDex2+lwCOg1pnSOMRrRir/AF87IIQ17Zj
udMKLTjWw3vASmrLw6AzhpUsqNWxPNxCZG7HUxmDz4Fr1jX4NomkBEb5TOZWBAqI
oLvbqUMXzMaC9zWx7KhFDWwKwDlKtD+HYg6xuucp0YiciPVVRChMRgQSg5mqhVuT
MFDpoPmtoO4tO9HZaL/BJBqgZxKAjUm5DLc2HZoLOQsBR6BeJ4lrmyAja+I2aQRU
NDfCeBAfiyCQmTntl+FSZQ==
`protect END_PROTECTED
