`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8mrx5Cz3KzdMptUip2lY0fUgliCAB+RpiP/42qLI11ONjX5CA9BUinL2ETz1e3g/
5UcBNPd/X9TdhmtxYjWybHORBQw9bQ8BquDd7gewxRRHcBH6UqlfKbndkPcpFC1z
cIdhfBya9qFbSi3RMNgowDvTJ4E42u8+TQ6S/OrW0ujobywcuyaz5BjsT6kXacpL
/rh5oY5yv7/BrOUUToRBQyFTJibq3vgPwTIG8guZtjhSB1NzEnGkpADzHWqKheQP
P6lDREcenkLChdZuDHkg1tytKaEA7PU1eBzVyMVF1fnvT/zGHLCcjBJ94zgGXUEN
q8t/2ZRKJc25etYI2NHxvX9KZkSNRo9M3/mKS2cYMOnIIwGhE9QRxpQLEUobrm70
hyM/v+pm7Uef/31tqvHD2YQmq0RsM+UhrKpldRyZ8xEWYNyjyq0/4Rt19F7S1Nb5
6FP9KvPZAwbifPXZMrZUYP3I3YEtan2QqUYOOrhqISDQe8pwNU4UWDfgv5WQpjZ+
7qJIIYhDGxjPIaQrBQN/Nx+zo/mACAzaU4f4sb0tyUw7uZShe8qju6wNVSuIlku1
jrPEfpsHulIhTinDzp+VMOTbS9HDNixg9pyy9aTeQueA5l7LuW/sFx+iA8SvSaGH
3HXpgNMmrGC1ohx/OCNRPozmiyfl8vCy1ryAoNfS8+Y1FxL2E+7V2CTVyICFUa/R
s3maFeqIiLOQjaHuXIAxHh1sn7bsEL7m/eKHqnnnoDwnHPu7FXnVSDJ4UQ34lq17
x15FKVcINIUgU0iHz8ry4Dpu97Gj3wq890NzLV7v1ELBJQflV/DQnCgv5FJ7PvMh
vzSzn8DY3FzUadgLXdgHWcZG2YpDU3AkTQcUVLZgw9N41hWXHnurBRLdQws+vQQJ
/6UoPbzmkddngYoR9Y1jq5sT0bwzEx0DVUCEcaBpa2lFzFCPTU7BOLA5Wldc2lSP
odcMgSFfjYZw/q+GUQbmxdR/+rwphCFIscI0r9LvgJDzm39nZi5j5lmIntBsPalG
v0o3K+Jmd6wt50ypd57G6bdvr40J7g6nYCAXTOdcbQRAmevIlzJYJUyvtA9lITM9
PNR9G05kCGAEtktGEXubMgRx/aIv+6HCQX50LHmOQdufQY2GyJgJeUrJE0eX9a2j
6N+VL+nSuXNJ7Vb0zSfhBTU4HzXaE849/vR43i7/NNdbUgvZPUXQXCfJ3jaZfCPK
xle5FEw34rvuiho/tD7knCGm8sXRh8Q8jyx7SP8nWgxPZ6JD/tQ6SjDyXptBUBl8
qHZtr+lyUlgdAo1O8rmBasVMDDh33UywHhxgzCaBphNXUgGbw9Mklrgg3CwDh5EE
qNrgQxkog9Ip3UJX/GNKkZuynA/uLvK/ynxwCF0crw+7xevlj4o8IWrRUCelAQyg
viI9jExRlaySTmJdpqMiYJVqbHeVwEGEfwYvQ7nbAADdbQSQKgwfWxdzL7E/y0/a
QbGACnVTCz9zPs6Unai06KcGBgVduYa+cHmCLHjlldGSXpfm4D6zaCRPqtPIogQT
ssh61CTA7NEe8F/lgsnKlyPMkE9SrDGcdSzCRG+kE2gz7l9mT98tfchbyUlpzp9x
5DOxJXS5h87f0UjavzNjlaKtNZo9hTzo+x8T+LKP0e9X0yNlLtkMnhrnVMw4Ft25
gosLyDuM89XTPgUgIla2RVS0Ph93JxGkTQvEptxR6zmzX3QQCRriHiqHZ4GjLYQ+
ShEe/MBOeDHAomCNZHe7hvgoOIT4AZ34dXQ9ra6//91XdTRTQjBZWdu3ZPaDmGBd
fnGn6PXSuIw0p7LVjLh5loG1f+JWgoiEF6AtzDJZcOzGVUuN7Jq31cqUlbzPW7WI
B+uCHkrQcOiWG2SzrSKpCdA4YsYR1tCcY6oTRhGc+tS14cnJE6O6YlpiufKWPzr5
gglykz2hEVz47Q65tMwp0sPXaFeQFynknJdungjiljeiLBiexa5LrYz5WK7+adrJ
cdhP6DS8NvLQqC7jSx6T8Q0wKzyV5N8bpdQrCFqTxeQ1fVRr9ceXQTDRkKn2Z+CM
9LxQzOpjvkbrKdIxhO3+DMgVD7F00noO3x9E2CaJDjmeqeMK6CFFHZjHI4rWCyGH
piljkWT7QAdT2qLo01TQdhgX6fLVxHYB7s5ciGbN7zopRmQFiCjr6gX7UhV7KFRc
BqJoOzrDZzL2RW37TmSjvPHlD2eWIaAM3nwowKfZLzdPeejaefV9aO8Qm4Xw/Of6
nHkLqlinJkZs2bU+sfyxkEGSyjWlN3dgJHVOglFUuzq5PgmgqkjUBIi31Go+K7jn
BbYHSAlMTWZ/N/TP8vvZY31BbNAr0YO/Ol+MUadT5BYk8AQ/pmpM9UjhEWDbed0V
mau//GNqcRfLVI660HMA+HUCm1F22Wn33n+dCdbaPXc/BxdisZY35O8S6bq01gOe
KMtrhQQ99+s7BNs95DLZ060WRzyghSM6BodaI+JTdzDT4+SbYDHUn52BKQb6mWOM
bns4FUhtp410HfnTEiqmuldPeV/HnjYfmXksucnLmGoQGl2BN2rQYt8WBYrvBMg8
YhIK8F/R/i/wAIEOTyZerAAMJBZWUs3go3WyBJFmh2herwkWKX60qPJ5Vheubsnp
QsgQX2Mffkeo3D2a5weu1WELmDsUfQcIoyXT8TVaw4jKwR+D+6Mg71s1d1W5rvI6
cum3PVnI4pnYAtWV6XGjEqDJfOtQ7R67yrx4PI+3QkX3kjpGSKDLViWAZQRsLQ4u
8nKqJx/7rxdCqsdxtE5NG3dhU9ZBQ0jQBoh1sGXXEqTS/VkyYegNpcnD5LyXrzm7
rH8szctTKoXvhwKzC1Zep6kPywp5fOCJuLxE/a8uRxBTKRSS1x5V6ZUsdreqzGc9
XWdp+ISQB607MPWOpaggSUFGpIPAzIxdOqXreOnj6Nf1Oexcv8qe9EIaYTTtVwUp
U+thP0V3eL0HsPw8v+lu5EtxAn1Py8PCvXQz/diLNQv9V40M4SAAPg1wowlUEss+
18Z+PRZVIB8B5b9mOvWYySwIbodY9WY9QlW/l3ia3WhFLbC/aEnWNgqIuMMvb2Mv
Y6VxCJRUdwJCQGKa8b8+BbDKMkafb8VU43nQ8I2Ze6YrdCEDE/vIbfz/0nfYZp4R
5nJ8C39qTvNBOFk9l9+BRSpMBQZG6tCLUNKR43GkGdujQ2CfCm7jkvkt3F414xCt
uCEJ6qef+i3bsqiXTV7kvLM9/ghBD6OssrH/7vXbaUJKpJsM3/yxlosDOISliewN
uzpFHvTJzHqsXnkbD9lX+w2xAC9hQyuBqfj2/+WcnhAu0g9/lD8G4AxLqyhJXDAa
Ca+AR6o+i4PhGK+wFfBe1lc3B579SxaO5SXSULur3UONfwGc/8YaB107cIOaG7t7
nqJBbt1r3xlybGis1BC4an9gAOG67nOGj6d3pwEcpgxMUWY/8/3uabMOUnSWyi17
9jV/v6xcedQtjdvOx3Owj3IQLRfVbR1iAv/PHW4SV1LeuZgMbcsZ5Q7SkgiJycqp
Vpk2qJr+m9CnW7NpkrZPDdmEOcpS4jIBQoRFYwrgnIu0fxisVcqvHEPmXsbnvAzr
YmgxP70rOg2rI9ssZpxEwMLzd2ACzyfugpD1q7PP2HA5SZrqGZR3c2r+vh/PC8e2
k8Osf7rA3NZw05odAj+h9a8MM7mQr5UklXQxF92ME1UTpDOPwceeRgNrWGNYgWZY
Q7cINjPeURq2yHyWGgA2djJW2UwYIQRlMBj6rVYk/Oz1dgVjOU6t1mO4pNwB4az0
UWCRs9J3PL33FpVuM2ODqpudK26Ar7hlorjMV8Z3YoSgQStExJxti+rU/MenfEfv
hukELseg8kJ0frN2HvAfq9WiBucp7fsLvdE2dAUZKr97xGnnIpsRrx077kPeasqC
L0jfmh4b7KxUmjQBdN2z84CCzL8RgoB9fvNwSWS9Uk20UEfZ1m/H19+IPv0/rsdS
Ld2gHC8lvA/Jimy+vlJEpC1vi3Ni2BhxDyoJ1eL+UVJOI5zMwzjsRjG/j+283xeG
g6RvPW4qoWrhJl5Bjl+Upaxq8n53tVsGJyHTncQfJFkD/XwO9qYmny70FOnq5Mdp
HmXIpxhLVb3E2y5kjIjcOBMHXZSVY+d6ZqJ6ssUVPRVoHZF5QmWwyhyEMn5UOLyu
W+AD0RtKdE5SYi6Jw2/oPkt9HCNNyyQzVmCcCC18mh9GTleJpfxN+WArRT0p6nU5
QOFqLBCoMrEPQZYK5gBu32Kw77QgOX9LaBgng3cP2Npin/j2zRaWNBVJBEiVz+B0
UCovYF09Rokw9h7Qb8s25DDt4Ni6F47lKYlYJ+NC4cvj90/cdf7eMKcriVvFzKWg
YmQdsNRaw6Li9ORsZQ4jX6Pod+OmmRuJX47AFyZxy9w=
`protect END_PROTECTED
