`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gFAqTRrLkLwA+c3cufT3gH33xlsx74zNL1hkQxggPyU3mxZdYwlaexIk1RXt5Ori
iJgLU05yFkiKh1kfkx5RXMNHS7PYuP2PK1Aw+mZlCH1csYNJt5BD4eJMblix2WJg
aiTJ7X9qd8LWzlPJBmgS0h9Yubi41AH8wZt9r6ictKyDLn3s5nWEQrGKBGibguRH
BAWPD3/ZlBtrBcigcbmZ8YKsBXCL988dVKbRJTsQ1TV9mtPtOzRghFYYNa/WbKJo
0wkzcPdZ/on8lGX5nQr89vUQPTKWAehlOAB2uCPdPoJKALAFbo8fvP/wjJjqamcC
qyJ8ZzyyLw3eiBmN+yfMxClBU/LqN8AesJyGIhqzKI40XqqVScZOV0DvwGjaEFw2
Cmn7GuHiZz0zQOjz78UExrRuDXSElsRceaZ1BmjTiQzlG7XHfBZJB8AvKX/MSP33
sMlObauD1YbuYhb0mkI2Ug==
`protect END_PROTECTED
