`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NPXDhuyQckqv5Gy/cOqrqLkWiYWKgie4eYqz6laSzd40nJBCup+jB/VgBYvoGvMo
95krIEyub1mUwmSOEjNdQQQYyBNFVEZ4MgIcnZaFFTTzUwbIoikvwfX1WhaY3D7Q
9a+B1Fd73Asv8MzGGcaPwHnsQa6ruQyiJK9XoLMazymIEFkrIkt1US0HPklcOyAO
up45h7OuTc26cBinQ3XV1R4EPj4MohffkgDmGM6YefvY4O8q6T2za+6k1P9nzTUa
YpYcuFid4LVtAFdHFTfHLTuc1LAshmYnt121T9t8S+SAl7AbDPpC3xH5EJ/kwByx
DyKrs0tsHIU2Hdw3qSEZfGurWGs3U9kHZtz+ICSdLWOdt9Xhl5ufp5PlX3Z4D/Q8
d2m0R53QDz29AGN8dkDcy1j92hPZ9fLRLNiKFXhGD1aAxKmsDchu7IKhtvUEHLDv
zLTy6d1oyXO4sXEHvWRhZvdKb76x01ueGJ/6QZtCAn7lWv6LofG//qWYnph3ft0y
g0knRHeXVVqmoueq/aCNPrCq51NmkpCKo7JehHSSn32+6cjhpZZ9L3xOZntnFilR
D0SXNpRusivQLhha2iZeeEVqontCMFUcP6ZvDKwgS6Uu1JeCywraHBUm/sLu83Zj
0R1cpUISiu4XRGn2LNjIzydgU/jsp6v7av6p88qXFE/T+ruI9h6j6hwDkQHs1xtk
e8a1QjfGhJg6eUSIdCu92tnJxO0PIcpW6t9wzHn5a3g7MFLJdbmfxBfVgLNenPQ5
QuMk3VP0C//yr6hf2pnJ8xxmnpeeiJH0uBJHSdeXQTVny82kxINbuZ3aUSI4hRua
m8lBLIWzlNnc7VFqLnMOWXEqxcODQMFpqt/uuKb8/4XbBPpBmvUrM9K1KpjtNYDp
w8NOmR/kFjs0DDdvzEXa3V1dRLKdBJyA4LD8veBuepDm8gHWsADceFLUfFjLXaZF
qrlsbpMqxgmv3JIXEL/WVSJPKtIpCyX9VQX0vMCQxAh5UAASA30xbCpYxXlM3U3I
WA3i43mVNnFs7iOatQI17+nAj6e934BVE5KBRgDXOln2Bb0WmtO1fgVlfJD1EGvP
Cxs8emoFXylvR1HuM7EKJocE6zl22N5VlrlX0ffEno/SKQR3SsTE02qUyzzMyn57
t++HBtJLIq6k5FAN74/xPx6NT3RguL7fQSKCr0byj+hSBgM/sSx1rdxrYhtMNc6g
YnWVV1DPkWWoG0ko7wTVh9rD82ZVJ0puDCalYyFZ8pS1koacEQBWsPkeLwSiH6S2
momLpZbAgktQEretpq9Hbe6AgGG1HPHQQQE9urv4P7EkpESE7V2p68ORtNNDLTHX
uJDiml4OpijeNaxsGamufkEIDe/FdAyq2Mi2ty0MPN6X0cZur4pJ/vuKnCQEVf/Z
ds5PSK910RpZ+BkcPP9ExNZGNcEKf4Kns7K0P86hrOWwHczPV8v7a+X/pkt15T0w
2Tafkhi+KnxWMxCJQdvN+vYdmsUWKzMCxZ/nFgXLUA1PNPR3qyf3RTD7VXLExZ1x
RjKjOJ9Xp/OEJyQyoee3VerP0G0X/72Byk8yS7mTdxO0fWQgYWVckE7sLT2g81um
8imcrmrLJ6VtU/7nXiNTKkbYCXE0p3OMWXrr5uSKmKT05izx5K/GTbBARWIWSa07
3oEPjc7I8RNjmnPJ6R5Eb4uu6xxj6s2fF23u5b+Mpdx8o0wd8fzp+It0H9/tza4K
rJ7fozeAwLbYs/bq2skNlSZ/2Ec9hCsBcs1n37a2PV8GsnG8W1CchqA018FxrydQ
biL45lBGpmbNoslNmPhcmQNotCz6Za+M6cZZHebmi/G+Sma8Wlj3gIaI3cvsdX0k
/K6i6zDcW84uTyJWSwhTgw==
`protect END_PROTECTED
