`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vxW0vd6zTATndDGU5ruDd2Z2c5aDWGu5TdxOmZxjfCFiCsxn8qpgC98t7HqF48sS
L6xDBa8C/37Q1oVgONGgbpDEwbHYT+KuBvv2M5V/sw+C8MEYTUhULbOOMpjY6M7Q
4ptfkSYpWN5KkHmTAKX1kJWyDAEP//kPINn8dowprsyCFmHhS1k6hypRokBYdtWx
5AlXPuGaILDqAJggXZD1yTw8w9psUCKpR50DLwQ0aTik8FgLRCH3VZHOFWT2MPPz
rIas1l2blna0ZILEA4OBo/j+cPFUryHdJW6wCumhaQfiPIa3ROgDHHb4ZIwaIGRh
WgRYHd4TIrEZJhjhMQrZYKsEjvYRg1nDAMPc2/qYnTr5JY+ieem7isCyrTi/zJGu
gQhJRXjkfTKRb7N7zLREPk8PURytOuU2AhHjhTo7D4h/nQNer+WdfW96D2NLSt8s
1Pm/kg44UDGoXKF/8Xf8dMme1WUAn6letiKG1lDw0XqBkr4eksIf5r7qd2tqNmSn
6k/nLvOniA8uJBOE02PGlkZnCmm2N1p1+3ZLK8qQEtki/+KxhX2K4FAo8LNwOTLS
ccQTZEIGfCCgEwZzYiDm9aN7HAuD1l+AfOtzSK4uBCack/ZJlgCtgxNKe2gB0F3M
QvIcM7WpS5UWgyyhReOu0YOg9zHx0LIp3wJwc118oYT3ipBXJ0Et8PYtgOdFXkSu
/RY4kSVsY30N8Z6TioHeKfLM1UIbgTEBB20yeodcpAwiibTsPc1oV6RLD6NYbvGC
GHhdY+V85YF7f/Its4chkIEPYgq9/ji9sB1mejCge9iLgJR4cg0YWkUFkndXmHg5
qE0GREPfXyGHZkncM4mJVq5DHtfhja4lAiXubbkGZIqxyartEceBLcf4WhPgvxVB
Clw4LZe+2QYk4/I0RjdBMi3GISIx4zqdRsq/eqQJYkkRxHRVPUfeTRYzvNfREyIh
7I0iLSdG5ynOmDlqdu8AGQJLfRO+rweoQvChm5f7MIOziWOxewUVXcnMEcam1jPv
nKl/BdyT3kHdVW4KL4euSYOi1drnLo9nE/uExc9AxBKg5MvPW+oWeS1MjZn6lOHh
EIdXM0CFgu0wmtXd5aCHehnDFdmJxq/0IXQUhootsqaTqZd3AvnhbaRV6Nyl1hRa
OMDrWo4bV2x5SWfdYlWAlWWg2wIMzXPSRw7DpWxVy5Y9ApTcONFNcv6JQeYkTFtf
o72dHXrPWHOlZaH5lalwqooCjnXqDBL0NUXfPnbRtHhU6X4ZXt1XqS8IERh1RLCw
iV8ykY3hrCqbDV5lMZuyyjgf++z2koNS79SiQj3w9D3wvZT/K++PY0iNhZ7/4Ist
Q5PfTGjyuV4Z/IrR0bYnzvurFNxBU5U3hhWH78WeDP+6VGNcLiKyrTM7VTorWpGs
yYFvkWCQ0/gLCbZtlxGHUw==
`protect END_PROTECTED
