`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/GM5Jv9QbQtolnxzT/LsXOOPGu44z+z8PySRj18VT9mMGvDO7zRFtDZgWkag+hut
2UnG0EZsTMYeEoZ4Dj9z46Pt6LifSmZbBg1Z8U3Tv5k/FOIPlCm5gUXekfWotzS0
yE6tXGn1PulS5yL1cJq9jJLSYJTsWuR/e5Dtnid/DazoHncKmICKy5H5xgYYF2vZ
O8Saef2vs7twvjxbMRpPA0XELRJeDL+3sdzHeFLpHXf0v/2L0j8fUbNad/1zr+LT
YuyMveM1X7eUHTrJTGBGXi2eKOZ2qmhfattx3tu+xPo/zF/OwQ0NwiNzsd9+jEek
hGFYEvyj7eoXm4HChsJ++acPURik+vI+E4dUpDULu+PnrieERsfHHxhuqDYrcH/i
5prS8maMAhR9eEirntHx8+msSOZ7UIJH52elxKQnypBa062vCrbvypkZPldDE4gS
7ZdcmqcpwomY+vMYO2GCYuLCwsKod0qbVVLdp/wgrAsPxtdD5np39QqtxPHQftiz
eBIlWlxVGUGaUjTaUMLvlE6F3gyPptXA2oELkupOPMa5D5MQRbwS/Wxf51bUyZ4S
996QkcORbAitWkeRA+XuZwrFYPojY62Dg+ivFZrK9W8ddNaw7gc7op6smwHO0m/h
BdjeB7plmzpeN/l0OXio6sd5NztUyNaXrqnVczqw+iHa0baVSXeL4uAuiiRZPP3T
aNzeOkbjQoKZfdu4rCnhDA5KKHFY3/A0IZ0ONDrowpDNZm1PXw6ZOJUQwwrachBT
PFiDIbI7PYIhgbNFd3RgkEXzcZo/QSzjy7jyexd4jdGq/v9B1FNXvv52E1fhYYgR
Xp8whj3BCfBtxKqzE0BsIOZIX/yjnSxIqwtv+/twon7zyR3cSE79IV925GOmlBrR
iMyoJRe2zrV5FqeDnRvBTHQ2zRqomXnrGjA9C6kios0xIfbqKydKgeU/yqVjw/Tf
chSGHlWyKIlClrW9Dqz3AMndY9BbtDQ6aISYT/BN5/Z+7vbjKfkieGBkduERwEOs
wkakLWyfLzpnUmEcHXKB6YhUZ4snEAAFALFF2lCTKYy9eBux+zundHRXIAzM5zJC
lwMNpJb78BXKDo70k6y9+eNi0JD3o6O6gWFkrM8Pj66Bd9oKAECWsC898tagm5v3
n1aRu1nHIvLlhEclGy1kW4xETvF2plhrko70RwrJdecwKK3eg8VBhJdloIplQfIi
ek0MJ/cdS7wBPyu1BdnRcmfUyXXT+lp0Agc/IO0w20ZIu9/tYlr4pS2dnTjd/CQD
+tUTwTrBf0i54fRzIWK8IS6SUopevZrz5GkW18bHoWtDV/n7MTxwPJtwXVWoCnuw
wB+plUYF0T9qnBXEoHx+W6iE0dpNe+SeYiN1TfbjHWHJqp4hG3waSs/1ovv43myd
ivNecmcTHa6yWEKRo13P9w//+R2B2o4q0HOSMUCABXnPn+wrO3dMX5FoujNQ+ROs
YFor9QgzUg8bvGzZ4d/SnONYwJRrzoME7TUlNmuHXh4oZcWWG6oscG1yZnpOt0Yg
qApArzHayCdao++KGrIALcqw3E5hH+z/MmCILTVyyNoLkEPCZosRzU1wDNWK1lxQ
b0fzYLmJGVQmNWyUvyYTmA==
`protect END_PROTECTED
