`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MONHIKzxGR2AsspZPlBjyhjwZn8Qp8QjM/Hto4NlJuaYPaZ6YrThW1FGoG9QZNtM
6CICAvtIhR13arQmrpWaJX99oRwy+5McWJAOYwItL8IMX6REEB12nnsPn+S+B/VD
wScyv2XvdRDoBSlz/bP7wGuVRSDCet4kiWVnbn3VryKaUm062MBK/06haroSBM/j
z3lr4XkzVW/bbMEnXQINdVsQPjPfIvvyu2uMN6bfQaoqNo3UNqUoJTRXJhYf7qpC
YHlfkyAK/wGNm8sVf++RRybu6vGQLPOaRrFvvQsWhGiZ1Bk0j7e8bCj01kP9Au+e
MdbaBD9ATyH7D9R+3bopllRgt76NVJgQtCp0OG2heYaoxC9fBSi91g1Nzgct84DA
AqozCVK56C38lT4M3QYpLyt+PAid3HpG+SQ9qTpm2LXw7FWbC3GusNU1lK1HeQSU
S3FqpRor8fw4RvIxPGiX3sCFZSXZWKhvBs+hlxHtROj6u6653ohs3dFwB+TGwpNr
Q1/QQ1cpdemlkto/dKfxl0U42eHA9eR/Mngs3lQNYnlNXO2bVZ9AHfd44sXfrXjX
WwjM7EpUYdkwf7+84PwQmnYMnWOwqDiJa2dnR/EsPnmlasKI2Nfwmz+WNS+++T9D
ZgyKcI5a3aKksMVl3YZuDDy93728NePuLmjHDVCtyCdRJYufZIRLCq3Xxs8V4ME1
74La3Yax9cdn68jlcUhk8q7WBDMGbuP3fDY8fKAHD0xnlyY1+MHLY+s0dauV7lHs
0tH2vPkFNfU17mj7bH9YuQdA62VhbrtVY5CpgJkPaTh2UclHvtkeldAHF9CF6xFY
P3RNnsRR8PL7qhOW52IK5gWMavivsVXDElHLQfSFlQyLxlUWv2WgMGaxmjxEpfMH
0UWW6Al6syYVM+UNdW1oQJ38QhGnLUzgQePGtjrfWIhjyS5lI0wQnwt86VM4RY3j
RBEdTMMSlJRnkG744c3xMgXiO3tiI1RqYzwMzfanoDoF3I9WG+SgQszh6hXG6X9S
P7dXwOhctQQWIUb5Iact9XHQbtwPyqflk3MDZo866wZ2jy83TE0t5OUUM9lygZBG
CFn6Azf1Xvagl0r7w1gDXirEAr9SHd5VLJcx23swNnE7muCyjrzm//Vy7IV0L94t
0AY9JUbFFk5v684vMop32IVhPm4K6JerAQkbiYDGoN21SnJ1FQDeIavmhIrkfsBe
HVZdkDy/7kbCDz50qo6KIn/VQ8qz2qfV+cfGqskEIw1U+9DOxIpBv3HTz9WRDV3y
60TvjvGljBZWCETeu3cUW5xubRwMCAD/mvn+2h1LOp/8Xk4gP8eer3ZsM5u7uRNH
uA8oZJgveGFzhRUhDqrNyk/ZxPwZVtakpFcYgaNqDgZY/J/Hge/CY6dqUrXpnWo5
/LKHTPRBAH5U/lLT9qA0uJKzwjs5aLIO5fyYNWshZbDUHqM71uTPT96jK0o5Ah/z
An9I4wJXBW45ErAV3q1EtyDxim6OMzDZhxrJ22CwCp/zl1FB+u3i14bETIGvW6US
rX3EdJq95GAj1Kok8N3pGYJEfxbB4AorZmjymqp73LIifJu6rsxGXJ7MKCLSE9hc
X8iWil4QEs9nHKs9Nzm89K0ZCUOxVBdLByftCc/aHk6k71iTJH6dNgk0vqfUMv7z
7oPRoKPurFeaUTrdhEVCRVkNOPNFGj3z/c5I4e00fJr6pfrZPNJCFyWvyXzxToGU
UCQS48B9PX/TALbPmyUVUiGNzJT74mygY7V0L++TIVQE6jRFkHH5CIvqaLQhtail
4nIOQOxAI1y7w7brm5yMuRLcBouXOKghUXKgoRfFQ0/hea4fBYVdj4jkXIoqkE65
uoDszQXxjIWsrRha6XmBBvDqewUqLPxKYam0n/cZODD13fJlCFCa3s1gn0qwogHi
p6lhYtT8QE9sCMoEf/DBoHX8sK9+6r1n0kfA8IxTghIxScWfbUUZb8k6hPQ7C9Nw
ZBJDwioaUxyspPvuXfYA9xtZSz6B1nPwPfaY+xkox0ohw3n5vSSL7TjFFpF8cuXu
JCH53P4hbGeS63SB132Yf1ob6whha4kPVjw+E2zBG7iBNjQOMobMLhUKI2mzKXLl
W8YGqtaDKgxsdb+BKo0h5RLRECVYjVaVu93R6zdMNx98ZfyJfxKEONSp9eHix4h2
3bigqLLtHOfR0KKEVm8iIYrTdkhptUYOgkhljAbUMDYfCgWkH/7c2TqMkFOl18yT
MVghNNWVBDe2H0hkOY17fWXVwzmqB1aWSLyNfGVgmlUX54A+sTO9CfImJwuYmo7F
5HdKURhlGAmwfRz+jFAmRKja8xuaBFUWjYKjPP4XotGDQfy4FX802Lgjr9sSW6Zx
ShKma8xp4i7oJxwvxWfojimKw9+0bTgVZjbsDFWqi/fZL2KqGLvWb5SZEzdteCcY
EnZdiLxu9A/XGBc0dZ9x7zdmkE7fCV8K+UiPlFfuxYTvRCCPfE+kWEwPSV/i1s91
mKtVolmgHCEJPR6Uxz2IzAZ1bsx3TanLIlYd7YtyXDv7pku9tEL/UJu13T25M+xz
gv7RDZGvbnYkRkFznCka+WCppi0uttU4QxF+9jJw5mzWnMQgUkjuxEmLKrdJqsKR
i4qaBFsBB+WtTQ+AmPYlxT71hWX+qNnkv6HxobHtr/gppzQi4T7xFq5HL941Rt8e
v0YRrrkBGueBl38cL/6Vx302JpIo+2kS+9/NIItrutw91M6yF+iHpOj6ov7SffXH
S0sfKnIkCrDi+wNfo0V1JPmtchhxOgW1EZ9qsEqBJwfKZzuh+AVOCvVyNhCuM1zH
kw3vlfcDeCDaAWAGbAE57ygisku5JGtEb5mIn5L7NKG2bdTwR+sdmp7tS4kEdoRJ
D1rQjLjA6X7YemIhc8W4Gde6eqqmkcLTN2cH0pn4MuF+64rur3L2miKketryaMAG
4Xrdj6Mp41Dq+xN2jxRaa+J9yBm1TgWG8vwwfGCR8yiWcSIrewilTlzThHyQND8d
lIlVS2jZ0glXR4NDSguZhUYJVQT5ien9OfK42wtLyTdq2UDQiw9lB+qUnAhhVjC9
r8806xV0nyV4XKpsVQvL1uV7JMGbKZ4+xORB2TmvGEr8i6Lza2mp6TUwWVadwPbV
Scr85HCLEItxR5LQ4l74JPuiWkbDnn3jZOyT6WPAa3ORcUAf9Vw6IOfJP5+mvHkf
B+kHxKuNttQ7rspGwmJiCwiNinHbvc/FEnLXyfzD68ChU1yyIEvBIVxmSBo/d2g4
Zj3ixDG18T/LvaIz78siaDe+AmapqbbOJ6nTfJHFMWZRszqDDv+NI3n1bNbx+q0O
Fkvpc5ckEfUO9hYZ92jNAEO9HyP8lCzc40jyWhtM5Sazd8NnfV2ntqqzwkpH7No1
JcgkUiOnTb5FoGidaYq15h3CeHGajuDvNYIfeVJOHAvNt2bDBhnhHdHEUr2ooe3r
Zs7qITRyICR2TsP/kTUJayW3puz9z7t/wk+kCE39Folg4O572xz63y0FjTtOjd9Y
00p5ZSz+qWJhW69JpOkZay/znDmyPkrBRoIub/Prz0cE87uodcF2WeULGcRVHPAl
dgqJbl2KjZGVjsavZtt/P1rEFTfOVOInWp0fbXvM4GnoXIk5zVC9nVBShmrAFEBX
GiDe6f43OfUHl9QxHgeZz6RabNFPKhvK/vEwg4q4rSsSELMuELzOL0zPxI+X0t6G
BYINRdQvCCJv8eFJsVJnDMFFV/dcZgx+5OG8n6VG78Twsl9uBSXUPACmiursu7Te
1ruKtEUc999zYg7lqNK0i5cJ3Uw8w3LGYlFJ16NPID5AsWxkVIbrdlZNCpi7OUTg
vNnUzB5cOMliszh0kgxwnuqYDqRNVyCWuPJFpCQRSYAknBYStmNhmAgWJm96yPrJ
C2eqI/EoFppGZinJ5Af1E9Q0bcfzP9i8aDFJMxGv1zzDmWPlGNNo/JhwrJKOjOJE
lLz95QXakZxiVtHQjN+gchbTcwZVoZxK5vDe5j/ewplnpIinQqixf7Z+w5ClTSyt
C9TUyy+mbCdOcm2MVR4wCDAN/Y1eNyj6o3SJOWi4SjTdlobOj+qjGJ6cLzcveKEU
5hUWqvyrRUU1x9fR0umbUO3j3aYpEZNGpUUnjC95c18a7vJ93BHz9KWMMqVp2O/j
ra3UqdlhOqwB3En/0JVN+m+24QvmWT9Ix7qgiv4HgwzB1NQWlGTVt1Z8p3aPYZ8n
DI3fBf6Jf/s9neiAU/42inbbYPE1mPlUISWnQtmbz6iR2nMGK7kMokesj2slMJim
QgdfygLCl2Q17B8i0QJJKvXgTsbxcTs42PxqAEDFoxWLNWhHPbjIp1kp9Dx1AIK0
mxMACmtepI0biKtA31zyE5WbCMmvielLNEvU1kGnYOYWI18Snb5DJM8FpU1VLNYr
j73WxbumY70/9ZiAPPB6ec5mFrdc2BdjjYf6cb75Q/5eWVxPaRZmsfkNs3pn9mLy
pPNdsP+YQATBpN9oUJFXsYKi1txopN2YTugBRSVLkVyCg/2pxVtp+oX/UxMHNVbs
umD0FNtU4bjFp5U4zHnzhSE1QqG8z2w0ZiVUvYUP8wAkNYCARNvZ6Sh3IksfIkiK
GNbeWCDHRO1E07DaGbzdz4/ItSscxLIa/4lrqavgdOEC/IS+4YxSSiZF2X2JNMmb
4EDpqNyrpn+B6t35DrmH2c4achX67InAjTBrX4HpVv+7Pi5ex2SA9Vm3jaIxWKOO
PE6uSdLpLbo1qxsaci7ye5Ykivi0GOc5CpxyTzA6lNhB3t/7MMNWP+/aTZFMQqXy
/JQ+/v1sp78jrxZCuFC+WhZ9qYGsVaaxRO1GeivgtA+fnvy1QHBRdz7sQEHS1P9e
NRbZb5QeZTpNZCSw5dNMgpXCOaUn49NqmrnUCnuS4TQ8vRXxLF3Zqzku09T5Vb1O
j6ZYI6XTxTFxAdFKyAE3nctOQM9RZrXdK+bZ5I938AiKrtQ7gfYF1/3ECEJPzP+E
b89ibkfYfSHzADxFaViUW7vazlN+nUoSAoctfPxQT9hoX+gG9XpfV38BcPYFy5a6
FyG09/l2m6QX/V0LeKR/XVMz/KMabzKkw68DS/mM+Iq0WoVpuy4zmyKaJ4ScWH7a
GMuFsrTyDVAi8KZfCU+koCdZaVXJnB58wuBoh1xpPfCBqqj0oS/GeSxGywl4WwXy
assilKiYMA9SdFlrTU9fowRLQ8AL3VxVjsrAFuKDk0dtdgxVvQ8h2ycx6wcv1UJu
CPji6RWylpeTj4rf4hg6qiUD2Ot0flLDZDvpuRshkjF/xaE9MMhzSrm011BTHhia
S6qt/pkwMtS66yLM3I9k17uK/KsM149H02VW4cZUQWiycQdO9CZnJpo6qpI5ewD0
Ukpkhj3xTVLimEVsE6hVy5ItkDUtOTaEAxWGSZ8Q9CErKUTaZ7jkRB9K6jDRQMvw
GH5YZ1B4RH/ehh9ifZN/mLY7I1iNoeua3kXN0pqYQcaFHT49YBi423/cVFjdwaVr
1HfKnfHiRDxpxjvtJEclFtYI3S8+8bVuh8YK16IbjxZ7EDoA8iIQv43wY407zYh6
JneGathGAZFf6J8o7ubXqTSGyLMyRASpASimB54wHalYx2eYcv1xjFmRrcIgqde9
Lcnpb9eQVsBnIiZSaYLCcVPPt0JWrzPdxXPFogptomvUQbLEXf8FEg3ZOg/vozUp
18YgLD6joNRHxUOWr/cyDy3mXzeLzln6wBLGyG7ITi1keYUNEczF0Q0hy/INWywf
vAruHMZIy0ti55GMyYJouKc0MYilGQrMommGolNOGDamzBf3ByY5aTYVEExGfvgC
pbpDtElCy9iNn6gPQtII52iEoeaQVVmxxDsEzgdyomnFrXi6s7p3XfuEc1Qy71FQ
EgHOJXVYbsIkgy3JSQed2pG/IgOru6ROofK7heeBzJ17V1jTpPwZ9Ze6XwUhEBp3
8R0QHaaAphbex+hTR66HW9OXS+cFNLRKKHgNEjxQcSjPPXjt3FUUBwC1jG9r3g6E
e3gVmwzTD7vH2/j0v4flhOeBSplA95qoEhvmVkcUDFbFTidm3wHaqChe2YE+LAG4
7yeo9BCA9BU+c9RUOSGvnxG1Hv+HYfU/l+TZ40N/H1b+2yk2T2H1q1GfTpEjcEfq
j6N/Qt1NC4Q/ZVOr+o0JNUuloibFyB+rdepAqzS44ji7j6af9iC/W6fT/MCJYNPM
wxlDmzU2DanKbtZxOX6G4YQm/bh8ELuCnfPQ2xT493JxoO8nX9UrjhFD2jcasI+Q
GH8u7HGaRUEQ0EYmj3ahYM6c3nwfV31ZX2Y24VnRJb6svAFpztYogWXgczYmKjnh
0eP9or17oHG8MeFG2z4YotWIUW8jz6VfgfVU77WFyV9SaNN/V86VEpK7onCVYg2y
VMIB/9PFyk8CD6ScoDtJOrhlmsOhC8OGD52slcShN87lQC+HqVSw/G+eVGpNlr2P
QmyVjE6y25J1NZ04CwkV5zQkn0pB2o8Flu2nWtC7ni8tc4EHJgbo8cQ2IAJpyJtR
eoq/6a1yDp2ACdQFoaCcsPLFBkPgbPhEArfe6p7Y45XKlHlHONmQDZp2Jl/WkQmP
SOvgR7j2QD6nwWwBtuOuWO7pTTPwWnkWvvYRUm7V4iRocvOWnWtqf1TCVUnOidsQ
3B/cGl2k1SCc/7KaKPUZvFH7DEoW6Ag4A2oZ+0dhSIL4jRZNHv2Uxn5psHfnJAsP
WjGU1YBrhu/ty5L/w3FPBScl9k2F0d0cW5lQaZV3XLbGGLcr33H7khkI2szyC+VO
A7LTm7X3yNqbmDKcQ8OQAbOHlPYIQQrAOCRxGMirxyWErjLGi6DnUx3PsK8uWLA/
drrJ4G8VdDlY5uOSbWDjmSNP3h8pc7hKHlg/V/qRZCcqxTd9VIvCaPebTXNCq20/
L0dKAPpbwcFVrF+XedmqAAm50Vv7tJPX41fDQLxURHmYJpNUrTCDuL46m2rR605R
NwQaVE5JuvM4P3yl4rEp8d4xafGuZpNFHGJzK4xLmrnCReYDInDfXi1id58x8tiT
YnY/Dnhy2RPMbCoSIzMbRWrA0UGikXD1/ih6eCZW69EELnGxkCpOTBYDgMT7uorN
JAEbH5xQF4OSDz5Lor6lf8C7Sy79LlKsqzO9Wxd+pXsY1/WCpmaPgJIirTz9RMbO
gWgJqY3/R5qKvzB+aSCJs2xL3HTo7Iq1VcVZBhTYAp86qaFMgwQ2uOydX49YV5r2
QINPUtvlPzB8hg0ENOUwta2rcB5cnyoPOX8B+F2OqBhJDGoUuiAjWHydjs/Ra9kg
NdTJKDZgp1+/bjGsH0vy3sbGXGOa0i6ShxkD16VeeKk7ITfRN2JE5nalTyg8Elyi
aKKAIxiBzvoTTagW4nf2AwQVo3ccfJO7Rzxj0swSAHR7tYQowbjV/We//AWB9QCh
S9s5l+2FlUaRKfGFu2P/fhlKylRoUHgZtFN+k+Jx11zcNLmuJpnHQVo5mSyGrEn0
xYV0EP9YhVVzPhX5pNnvzr1ocK9W7t1JYP/ZF7GFfn5U6xPLracw2RO/qmvVI5uT
+uTGLdHkwMffvBNquCU5TeQgwzDTvTifU8QioxEh2J3Xx8iPhJo6dT3pZR2H5EvI
UvKXB7GOuDakqpy6zjAAuj8hbudywW5iaU8tzloCUWf2PT+S6Fq8vzRP7Bf0vr3x
tE4AUM5V8nPQpiCX3aCyu9j1uH05FVkkOa+Dnz9lCl8JMeYMAVjS/fuN0Q0WHFtB
ZdSKcTLaxG1FtrMtu48RJv07hlU7mIp1UN7bwKu7JLIap/EC5WyeylKnTW+JMD6L
cGG6hVGx6s6nQTOAlRaFMmsQP5mCvXRBkPrKJGeI8aE0JRZoUHgRzjsI7tz4aOTW
Sxq+VWyy4q6rk6NFUqztl6BOnrqAZNCF6XbU2OosSPFlQCa7nQ73zXhdGGn9UHYP
1QStixixrzamayd+f31NHqMvR8I8eJTpYamK1B4O61cA0aSJjs+u33o2qqsIHCUt
3m/u48N1o+gZuvbgWRZkfw66o8XFLpc6S1mFsAvl29SsIyJ7AdKehmlYTcDA3W3N
uLNr+W/8wlo0QJg6NDvbPu9qTubOFSM6WcOKVFjiptQYcftqmyUlHOGaqTLAVRYz
3TsL3Jtp+upBOZqQL0OCBn6Zc8MIzRfm84mt667/whCSW/HzdwCu0PCBY/wpdDw6
kue2B4b8QY1zucOjDNJtCAUxYvZCfBrRp3QAg2M4n2vIbJPWQKtD6Wgpyl8dMB4h
poF6lKtXFWWhWJZ77U3uRtFjvshLANtHMFQwyvJ3/70byiZ05bYruFMqLTXpJSw8
BovLZNFLYIdBnMrthdlo/km2f3m3bvIBzgFLJRPLNm9UxD8tIQnymT94Nj2hhbVT
OQbQWWrsak9TUsHGnQPTQSlwXp6KrQFhNj6S5Ya3ST08NjFcFKit5xqRDf75mBri
f1ze/mVP91Ws3+gFgkRAOYQLRhrxAvHhpqPcVymXcLhPaDXOpqS7U0dHCdPh7vYo
VY3OaATkQ6NzZYSQc9EwNKe5kUndBPil8nvjNU3R1GLrwJ5P5KLieegNUehQvpPu
5x5OKZPHYqulJkhWrZaQIwYmSXzwy+CwW/+i7gZTolzyKPNraebQaaFhU0hBOqss
IM5hMdWhow3gULhgCwUlfF0+R/8kvD9xpeeTIJnGiRb4k+d2Gh/mUTc3J0DdjtuS
Kj0WIjSoUyWAjDw8DrTLsmCx9gToyVsRx/AF0+GbL/83z3q3BmBvVhABmz81MjJ/
Ghq85B+JCbpmY8L5Y7N2Xel0lxI3rhW46J8Aj8IfxIc4lZ86j8KO+N2yKgKaGA7r
6Z3IXRUQRMGiW5KxpZMTUMSdTVdMbynxQvPKqk8w0pw6yh3N345rZZU5ozmRB2F3
eOHzlMnt2Ll9X+2soLQ3b5DIqPMLvgVJiSaAvy/QfAdccrK+8v1KGWJno6ZsryQ6
ig+52sHQfVAcXBejg3cX0fKS8e9RYuJGn+3qy7VtsjeXJK6zrfONBre5qbjGVf/l
vZiPkWW/7YzKE4Y/H4Vs7MP43mJvQ3/bZEUh9oPpaD+66PefZkVxCMS/oBe6BaP9
zFjBAacg6dF7tNSz7jug/EKoslta4wpXbanosKq0O4f5Wa0g8oriSg+TUDeOvbFg
cC9eMEGwaieICETtz/vISuAuumdiQp8Mkec3aAjsfgsRgMLWePHnYuWS4STrQCZo
0vmeP2n/Y7r32wy+XM7TQwc2AYRPNVTC2AxDT/krZLBD+4oL2KeXc3nEp02Kd0YZ
Q9MfZ5wViEpuE9mHYfBovdf0cpX4BXgr6JvZwHIYoKpqMKnZK7ixux78zaa/xjet
bXFfBMXF1mki4iNB0CwnUthkq+fiClyjwtqhLfuOf0/sUzvDBSgkCKK9xU+YFZbe
IsLD+zDOwsTdXAOOUfLnnwIXwEFZPndlgjDe0/Hl5hAR7RronFNNMVus806ULWeF
wK/vuqsQoLSyNIpiINOrhiekcDRDybfAjwQymdmr35U/y+tePgRJDoqHXAmPVgW8
5eR9lmmVccbp7xYaIvurFoHVZykrxBgFmpKXE9C8sHuU7g2T2/tWjsR5pEBDRkdq
A+rpzhoRHfYWzMATvm/G95qAAkZ+cWxIJ3floZDXlxVn9pvzr7wtLqZzQO7vq9BJ
SFmoDJJc8hHXPzBPDqBMdARDsM0BfLuL1W9hRUlOcrZTO/h5qJdPhDZDYrXAzLnH
oeCxir9Boy+w4oGICgT+aJ/gTis0V8OqQqihFotjBxo3If6v/ttGxcVo1hupVCYT
rZi+wD1L5lCuLAGCJv3ijC1chqz6lgdkGtxHWbohl7wR4kpxNqf4qm1ZLOOdZjMc
7b6QnN5svugXgWd0SOymt3cLhnsV/TqCA4Q4yKzpyZgAm+xuhp1C08qUbc/Wkgxp
LswtWMVNiOqh3K8Bh/JZ6akgid0C1mat/94IiW0RIjrTvW4n8zpkbnUdzhpLw/y1
xKnxhszwune7C5R+tL6v/nAesY9ppxGZbhrtvmSycEW4FPm98x+Jw1UDShyyiwDe
jbg+JlzWPHUYD83RpUB28jgpFlKUukJ+ciK6tnDlT/x9V0l6ZzZn2nlMTPw4yeGs
Wd8f9YPQTZ9lA6LJt4GT1rWrWJPeYFbCYN6odm884Kwu1IdsNQ4LjbKP8RhnwtIz
HQoExYF0zZ34y+iib8NzoO8ZNzmEvw9S6rY9fEgF/yCJtpDt6D/qpG/xNmv6AlTp
mZ1ZYDl3YXvGG3Xz5FWE6/KnsgxPwZxbZbeXFhuRVj3LeosRoQ6Yt26F1Ma3SK5L
uRGAloeD2ppMGPiM404FvVBMZH/uQtcsxCb6drxZipI28Q6GguTnBf96QOzXp8x0
YCq9w3I0oZtWgoVXR5jQGs7dyrQabP7KUQFnoKdKaJV9zzZaLnry4DNNyAFSPKto
0zazkSZnlNcr6lOvx6qGndUW0ZhGuw6YTXJGU2TNHpILF2O1Q8FHdsckcqZD5ain
Gdz9PAaIZSOHKsxx5HxHmezFlm5coqL5ssiFkEYTZpseNWGL4cWesISFGPKg/H0M
hWe6W046meB0FmsXgQ8cPVuZ/r2o+566q4CjipUweC34J3Yn8GWJ1h39Q29J11Bc
ZRgFfy6zWWH9zKmL9sXtsnEO4DInangh+HFiU41iWAvnW/YnrpNrPcV3vMLxTHGb
fNMkjEbUk0rPoyzB7elHeMl+IrFY3i3kg1or9UNxTBV4KFcO4zfSuAtk4A/rE14I
It+VEtu5eGd0veuAbpNCQRs8omP+3VVzHZqsImipCaGjdAPu+esFUbiL9r1N3Jvu
CxQ2KbP4GuVxkapt8N1nRQZi8lpkEn1FV5UOo9CqNp0kMAADeEbKK/iva9m3a2D3
NTbCyn+myNidQUMVTlkcjlF5NJ0QKCCHCJFmY8qGoP1P2yB00Vt4Z9/sRZEpRCE7
qan3H96jQ9fJSsm9UeZbDGSVAWkfq957LjbftkURENagRJZ+MD/GFoQyQXVAOTt7
gdg3D8GR7JbBSeswYXcQzGgQg5nQp/ri5LFojy94ky307NfSHNJ1iadrNW8rwPR+
VLljrXNC0GR+HwOA+HiAFuxGCuMrKZ+onOJOMunoq+2zkc5f+7QKrGzQq1zkTENn
cDRsZFQW5H1LFGQx1l+vu3YcI8n1RdQDYU3WQB/FnRuyQYzrSSboQ8eGwwzFXU6f
Ut16m4Km4HNiXi7Ly4l4wnon2jR+tsPPibM5ci9mio7bXVGeKMwIrj8Hqyar+vmk
YBD9LWh7BUGW4R9qIcyTPwlWfE5PjA641KBiVC3yjoeeibg7N4xB0XvKLzY/d9gv
dVgDVuZZ2HilUkFEYi+8Y4xPyJavcLHGyDJ+PWyC1aCVAa5tQvQCumpXbiH0MO/e
NdWKod+v7oL4rHtWIVxV8WvlFJcDQg/D9hKQ1Ihw//XplwBVYONXwpTU/O0+kJ5F
VV6krAJb1BlhzNV4241Da7pEc47ab/Yw1hZ+Vr2N+jqY2QZTMYIEbu0PyvhnAsPp
uB6vyFJGE0qshELnDCSY5YycgFbTj2FHKpPNCGAoXu63WAGn2lpuDx91tEwHtQY+
mB/s8QWht2Vucc3jklw2+XAkQz5MZHWAQGNh6Nm5STqUOwV1IOV270DljPB3eJ8R
TrZ4b0MAqF2z7Pcx75FJRLv3DOF6skDxD/L6uygMeYoM92MzyVvEqo1ikoMLpyGA
HfbaXdpMA9b7AYE+fSNmopyyaze3qca7VpbjVFCliYYO0s0/QoWI+/i9PIOnslqz
acNm+na7jWZq3ePVi0QO/qatmbtBBBEADqfLv1sdEYsckuS9mtcjTt4wX9WLiYAS
P8pJdIda6HyUqGg1j0RCJtnICwwUP4bYighJaOR2TFjJnVWcL2ELPo7FFo0gOl8+
ykBSfMcREleH7wK4adQR/KDvB9IRptfyYKokSjAWmJgj5vbJ+S63gUa8Xz8AacPC
930nZ3exR3nejHuK6CFjsuevIun4UibXcWoHmjtXxNWWYWcHGz2cuMpvJo5wDvcg
0pPsWDs+ohdUm00IoIc9LHnnRgYlAPtSUwVF332aUCF3KcFCNaRamdsVNdm+MeyU
YTsKTdt82wpus/RyvZqasHdXy8rzGR2avPXSxw066/qo133Uvm2ezfM1tV8yh7aj
Wv3Ij361YGyxe4HzwpJFpnvFyXAvFo1M2UEE5LeLs0LcaMq6DDtsvCpXi00GIOPg
q2/ruRRXjcwTEskkbz0slK9CLuY0WniKuGLQNABwZRidv++5xDC9VxorL2o4nXBi
qS5+3SZMHpJ8mE+2EdtHoVWxYssFwiQl62Aa19OPN5ZqVHS3neRKQBr6qNq7EVUn
5RufwjY1RTod10t+vPFGOby65bgxSh+3v9Z3ErCVlUWqhbx9II9giW56yzD4+VWI
Tt4SWBZScxgKI1yp3f5lx9lWhdbyMoZxmNJIk/6qPiFDI/GCjb3UuK5F0wjIqwgI
jdA4r9T7wvfTPK/U/3+oB6BK69NuuDRHo1MC8aiaLqzoUpRhznErhIiE8MpOrD+p
Y4x5MVFoKQlR3o6v64QTc79V6oWqCdMNvC4+OSskEYJE+VwTXHbZWBeSCDMEf951
Lj+W/uEh+mqWve9dQz4acWYxLD/MDojGmKr/PAS4p4Ss1eROqiFMqO1OUo+chnCl
NkiVbz5VgoUKMvhNDRaxN1DWnZWroMAdAlB9D9f7BFqYe5605MlozJ7SaJQK5PFe
wecOJ+WefCRbAbaZ0nkCoyk4zSSNYDNeXhm0ctWAdfxWCFqkjaxcVcdsugri05VW
FSqhLm9iRJf5Kp8VkqqH0718mBmTTzPqkRfNAZlZjgpdeqEj/AQVWyT7nfEP/Iy5
YWhx07AMZjWrbU5UL1i4vLoL2CqqB8/E23AjQwahkTzhEKx+2x2PH6MyTlHxmx0S
sLdUC+CmhpKI0pbdzNAXKcOm3AG7g24kZobSGeymqHmFMfD5NsPZ5NJeg3kz0TcO
rDVabZ0pwz/7fD2Vrr+RlEdYzOCetXp4Fx8wUzjF6robyPK3aw6n+lXfkrjnh9KK
F4PrL3zN3keAUEfRhuUUbmA7VQL2b+fEU0JqDCyBb7ZV0946fu5B5K1gE0u41sab
Oq62KxgYaq4z1cV9iwfdxJ33JyzNasCTaqemfeszROghGh3qLVgwcjmAyfckIOcP
NBOVd7WRae3WytmKmGqRJNbSWqPhVlV7SAWFJg+QwLJtE34JoJOUldcY+e963XH0
wLrDn/l53Zftl2KCgHU+ftd9PWBSxEues4ALyj7QUNft3x++U9A/6iw/lydbDwtn
ypFi+FbFcP2P2S34+U+TiSfuX9jv4B+GrexbAvu/t3SMiEx6fojhmoFde4cvGqKI
oDLgAd1trDl9yanOrpPZzVFlblEo6XiRsyvgKwiOFG/YwT9LnMIxdMwNgowAnu1f
bQis0CtbcMIRP9BuJy858Zc2QCmqPMW0ciPOPzIYVRpEKS8oD4tvLHduW0RHcIey
6KQNthPV353pZ1v7x2siBPdTBiL3W98Hu9HNfJbDE791r4OCAODlxhMyh18EkQNf
nEEH4Va22vTOO0TjAhSmUUACuGbKcoScqyo6Mco0saXxtO9UCLnWXh86bkn1BX1y
w/bPYHaYar8Is4CxAcHlu11UqJUJVxEeNWXVngsUTzOmmzbpi86vaP1a9ZW2XrK4
MDWsOiN2n1viJjYfRcWT2Qrdg1qJucx51vBcgqOwe6EcEvClk6rn9MxKzTEoRvOd
ujXQ2Z4sM9tSAroavRSm9sZUYpzLFQrGMWSa8/Zu6VT5p+4ikILuyN3bbRy+Cnl7
zr+C1mwcIMe5H+2p/hMTj6YnOBHOIop+vvUwe5uZRXbNxWxgH9Wed6CzZz54WZKZ
pYOWjzmuqyJPRqsOzHj2a0Ie57HGJrRtk08SylA67uak9QCxUfdIcywjJVKaL1gW
RjEuGX6PEUOo4GYt8RMAdE5Mu3R45amsWUKDHpoLCenqnKO8XAX7v6OMmG8pYCln
ao52xyI14GEWPLEnHglISXSbevSsIGg97q03jT6oe7F7DixY52heY6UGmDlrgzrN
lsknIZJYUjsTgTs909hN9MMz1liW5IyxSguT017yp+sbrw7qSAm0pEYMgABB+Sgm
Pp6T6PfuZTT/9SL/Q9ue9e05QB4t6guXy6tk1LkAfSC3D7oPjIeQyMitGQ6Sa6DM
dFB/DjfHl98uTUXplzP1XxltooMjlZocf/nHekDgEFB4JSjdI8fOqa/MKmESfRGq
7x/O2c0wmkwTxXa0JoBYo98p14xJ0g+A2GKvWDNMzeNFZ4aYrAskMfGf5fjgfUtb
p8yUpcWWYEP5WjFv12WJgDAtV/VAsVTGCERljeKhTE/fGFjG185Nze6zEWTCzEA3
3Am/sx0R2EVNl84WBvV7240hgoHLE6k6R96RxJH9CofcpHYBAr8qvLWaR5dTQI6n
QMyjLIHyAfi0LdIBuUvgR/O/RliKWZBC1BS1U4q6O6XRImNNWup9AeNnyusi3x39
qeiKyVOZeRTo8h5FvlaKIDxjjSpApUvVWeK8ibJ26gaULVJD5GHyBpTmLCzWGMMM
K8WkvtoVOIDN0F9x2yCG37a88DYjnIopEfVtNJBqL983JwXXkGYj5dvisWe6a+BF
XDvwgWgZYrJHJA9WCk3nQhjwwS7zjth7fe0oNSJBbux/X8nZRxQDbHPSkvGNqIZx
KD8b9pjCwZCXwsQGB4jSVaJ/FbCeyJ7DawvXhEqnH52T4WfC2zSd597yZxJggNMS
FnivmA2FbWtJVQjBnhJEGwKIe1uQ6Djw8kMDkYmhOIlt7kmdnvb73q7DIEMH4gfn
ThfW1HZlvbCMMB4XkDb62VVKkjVg4AeqtN33bAVRwjnupNATT1OdgX7CQ1UKJWB/
68h0uWW4R3QrnUSE43dCpzHkBlrf3narQva7qHh/zwIf9rJEdt21Xcn7VC5CA5S+
PkXFnqKo7SA/XT/XpFn0+Om8WW6aVAuO0RbAolJEp8CItHGwm7enGWHLX9CWg+sT
r20ZrRcVACHwdplzHi50/4SJS+CH3pz/KPxx1YpH2Wkf/pUyq/kKoTjJ5xsnDaTb
ZLcZXwdLpXbfiw+YMBbsc9zhWA0Jw7ti++MKshFyxXngxui8xLjPy3lfkxrWESF/
VS7MEXbC1WY+9ZoQfCtls1ex6D3SWVG5yQAJWfiRNJ4QBEh9yuwfFI3RCzg5G9my
juR1NkrFdRClBc6kpCOxRwESYIoFe0XDJA9t+dfG6bFnPoxad5ndQkQXAwFSiCR/
ls7hA0794u+O1zGWuicJqlUmAZQPDfjG6WId7DUpuxQKwBHMdP8w3micoRmtURhF
uBNX/o3HQg/lRg98CiZse3LeZz42mrovPgLORa5V3s0TvQZqf26+DlA5+WEtZhLu
yTEvmZsuoHMLZBQ58I3lyUnq1C84CqZXvJjQszSAasoRRYtdlvD3dDUvh4ezzkfS
7ft5GokAV2HoABQHYvsA1osymgsQ7hV69q3HwQG4s4iI+Q0FKpP/0W2za5DrcKEM
OAV11iWJYZv7KfYB8ghGPe8baDGBFVMFlrHbLWAe1ta8r20wHjbeZfNIww+1OWR/
IY5GcrsBnPRbwb3EjTRPqvnFvxiGV7c0Uth2pR7YHQDD0+ERiqmB5NMqyOw2Z0Tm
F5kvowEaSjHqKu2blPzJbZ5Ltx5vjRFy7xXJIR5RdtNZbEVi9eUr0epAK2N0Qlix
Tg+exfgNsDtdPxHoUGwv2Br3ANAopzy14vrq+m16AgamwOCu0nbVJiZ7wm1BLQPw
XZDN45FOA4jR/TV+mexjF9c48Lc+s2Ii1nq9qVFKDVpS631IMMS3CCw4y1Swhnd4
GKvWoLMQ5K16OCkmHkHndVa+j5EUw7q9x7E4uJ7sEbXU24XQt+BdH8/nl5tKweV2
Vn9/EM4MW3LuI3Sa8miSPibB9bcXeKOa1/LGFZ8QyWpV0D3XILDjXnqdl8Op54IX
xYXWQFxNKKs2MydlsB60cSKUbTjqMhhmVvuVOTKij8gH6UM2nUxpoheYA1vO4PNB
WRJlQDi+s9+wHiKvdUj3OVPfhQLiLAUoWktHLUqCZUMj8zE4C55lTawyZf2oAGE7
vcDu6Hu/S9hhf6qMhIg3hKKo+8v+5gp0zWyIBwfEmtG17JaUNn5PEegRCYgVuZMT
Xm2P5NLerZByEocQyf5klWPHdFzdJSmAo3VdH1UNHvpSDFoTUb2+Yts8aT49qKFq
rzYlzYSFUEh3uQ6KjPJVms5tX6hCiCQ0hbyYSl0IZ9/GP+I6yT7bIX9ExjkuOKN1
MxQazppCXgUf04axE8kcG5yCdoD6tkU9ZQe+tJFjXA3oPZn/sfqN6JDIknTqVn1G
BPnv3MELnnoaLQRJ22ToqxK4XlJ+bSKjhBwzW3a70zRp+t+ydG05HiXHe/1ynPAp
4AbB/oEK36ZbDbk1+axyyvYnWzND2/q2yi4qGbhg2MoR42SicZnsP10vs2r7DQr+
h2KYhCNjjoh2YQl9x5DVUY1k2zlga+E9qzEBtB62iGS+p8C2ICBTlAHdZCRxPfbN
+4rzWgqFE+WWBWQYIBf/3E/otgcg8d47PyklE04XeD1bihsdv/nZbmYE/sUvdLU1
uGQrRkT3mMRS7Acei6eD1Au31FhxojfbmMoO9cVQB54GgLfc9iI5LK76nmsNkgYq
c+AuF47IG+DOlHtHuhpgYtqOiFwhKUkxYnU8oho5xW8QLo/lXNGga5tYmpxSSxqz
N8/gzIK63++F5wt0Rr0z98GQwVemlMovDiIrHiBjfgh0WxolSOq30c9WHPaFEn8V
WyvU6fsxE0Lq2MHtLKEHUTwLO0gJuvM3tHXJuRng2q2osNrgIv66vWy7sgr04aqX
kobEo6SieeYVrRAbi59GGg4jMfvb38HWaBAVsPq0w6LjieIzB8ZsVcTqPKp7VVak
yLqE8txpkbqXP/pU5jFu5P8JgFlxmY0CwzEg4W6v0ov99QMTVBNYLNp9e0KikEPC
Kqi5MxuSKjbEsUBKryYRsVRk4Sxf/BLC35Ck4m/TY/bHDJ2ZL1QgB+vxGkq+cCzl
r3tt+MQME/UiL8G7TGDaucK61MaRFyyNGPTqNogCCxPydJkKqqVj7LzTzSr/pylt
stC3lv9t9Uak6KcX+ObnQPjK3C5N1tPBaB978gr2hksanu1VU3I37ILIB9fV6CKm
bahcV27FxE32BVum8lXGKP8otjL+oyf5yPIFzTV8k3K18SlnTlsrhA5KP4P2H7Yz
yNTjdCUzcf7rXdBhDLDUGEI777njS/4clTCntd50axhoTO8tpzBFc/r6AC2H1B2u
pZzBSWmYyBE0tWEvRXIWfcAz7J1VL84LbeQe/1khDYLUgXBqkbqZnsYumf9LkmeS
NiVBwgoDZb6RL/W7ytLMI2V1IsoYUlPlwlfIBopRhsC8t1jB45VP9uU2EmZvc4I7
TJfkWOgLtevZzdV3EgP/wGw+Xj75VtAixXPqICrhd+VwdChOn921uCHAqHbN5EyS
2f1Ehik1/TeC2N5j3x1r1pJG+Z4g3z9sY/HAAv2H1UjVx89etAOX5g3HYNQuaUMe
rnzTspa2j+SoFUM3guP+h+3Q8UeVAbTRqsLKH+cqU7lOQnQN91EVe3e4dVwEOTG2
Ns0OM2d3Ly5tynEZcH/V+rB9xekwIJDRQDPBHU6UyB9SPmyN4nv3uZXt0e3BiAk9
3Rk2PTyNI8LDx1SdSqmK9cEPLRQu/NgJrvYCtcC33zGt3sUTVsMZk3vcUUiAPvio
Q9Gns/gh0XX/cYZE7hHNji6WPML6OjaaIKIiHWaJnG1b1OGdJqnKKP4pW9oD+jJy
+5jBj9EvXN+f8WRw7dpBkWqreCxkMVuduWEn9aS4/nQFwZi4l4Bo6Nwo9j6GgxxF
918MVs+2/r7G7TFqyp0cUb7TlzugYMFyMzaNbNskNcF87wEMMUxnhC7/ncqYUDHn
UyFs3Ka/knWlZHHuGXfJeMLpYS854mb1HT3LvzNUCZd1CM4a64aDC+GKuzWFHg43
2BPkkkzMmByczmwGSTKhEz79fh0QfUONZggIpI349T+Wxd/DqLMoC7eJLdS/Gugf
+kGrw+i3C+qDIXc///tGuwd/0uUHxhSgsYMHHLyWSALMFGWoJebw7EQugcv9DsXt
YEQ/RRAHA7KbmMk4X7ElDh/Ke0HlYPN1TYMDsnAgFzuN/+nr1DE88zWlitks6sLc
1XBcDyBhWDtq2Mmi91CoEkLddGXi042bvxtLhe5aopHjDbT62mhfl4x2zwdorORw
U79wqjcs5sNzqBzgUZA9w1UTCWWPMnii4s1LHK4ncHE6jNsMTF4sK2jpr9Yk3Ci0
OBAbGJUJDUg7rM5sEufp9alb5/86hnXAlkH+aHWPKChnynETuPo+6xk4OHeQEiyz
FIVpENYlLorjoP+dZL931sHJAVaqSAlbhZjmd5aW0utUabr848l+i8Z2FPK+Whjh
Zq2ITKuySocUAf/fb3XTN+8tZ0Wj+b/xj52TNy2tn+Ci1W8OxIxfaD/MtZseZG3e
C2OTs9FTKCL4zHcb0/YUkRnsFYZYQkDPksq6MrFGRvtWw7ibSt1qmXMx8rRdkzQ5
0ezMQCB46nx7FlwXnfOA655ZRmiVksMI+0jXk55yxryYwL29RMDAJgBTaXoG1yT/
GZ1yWDAUrdYzla8adv6u+0ADN/2gEN3qshJqvaN873BwSn41C24nOQe6dsLw6OPm
u2uHRCpvZ1y0aJr4OI+svHOXUUOEbeYuCbbjYWgEpJ+NU8/JYcP6Xt8NYgInEjv1
4Xk7p4lPinOZCoq1AWZhJeXMbFZYI2O4nQJIiIizXf9oftw2sabsuK8qMxqpFi4Z
jnH1ZEDMIvIfKLquBmPrDvmwitqPwU1jvBK8ulZ0sknTRIWQtU4GiDow8l15/lcT
R6o9WA97h/HV4qQv6k4U7yqKWwo8TfYvXtjeiryKgXELkwbqCuWjvNQKcZwfMBar
hM2U4gEsgNtFovBVMio6aHggHyS29yL8YHfPGa67+nVpYFKby2//mv/4mNDxvwOp
GmXDjCKgKYFwR2buF3ihOiTjSf2P4gVp37mTdu6EQSyiARA1QyBj4Le5a4pJj8pN
BU3wZ2MI6GQHPJsq2avk8Ux6MrlvIUrWT7AigxUJBkOLDm3hMmjwrIRngJdtz8Yt
xhTSXjbdfIBcIiLYGwa0kLj1lK5N9u1BGsAPDrxlNgkJFIv6rBrpJlo7mGZ6L6lc
uVk6BsJ2HzY8NSSFb4jodoshUpkPoOFaL6yREb9m5r6VJdRWPrzOoFMEQg0fxSb+
GtZSShP12JC1KUi3qXUBPLLwKxqas12mJozx0mzkll3sHzLpQeh+jXe5jKsaeMMH
9SBKc4T7YeL5oCgB5gUZVQeRtesZKrqq7E3QsLErYnxBQjJXbkcUeluRETNbfbLJ
XGw4McZxJV7JTwAlgk2WZB3n5TaJE1yIVoYMoCgUoI7ALvSKlYsm6ifNlaWsG2WI
CFzMa0B3M2cCR9YCbJNmkszplQhg5oRYiAfXz0Mh/Ymbjn9I57DHi4FpV+5DmrxV
qDSSVABdnOTX4xfq+ZgiALXyuTngziNfIFXhbSNKh4P2P1iALcH4FYa+LbI1FNov
uU8ICo6HqyB/oJtZfqvzNDkuoBW7HIqT+xY1Qzdr0NGEFagVQmZqDUUxH0M9vEcO
Igkq71WtmQE774hURMUEiq0L9fl4MiHMZPvbUK2apA4BmTlOI37ghrbHFRD+itB5
AF7WyfRogjZD/8N63RKO9YlTrFaG84ilE/kxN/wixicSYVxrbZ/MVjnWq8X1jKE3
JHYoKa1pbuDhGGRjsFEiv+jva94Gz7YROWYoiDeRE4YGSwt7OlbGsULtQf05HCKD
bJMlPaE+lV3HtJEsbXTj4KX1J+lB9Nr/HcoKPxDfHpNWiqPspLWmv7DSl3PcemC8
HHksCdse4UjdWEz1oS3wohj6yqa4kIk5VjkkNo+d8pXVRtK97ZxT+oq2l2sCSiLy
FKYchf7H5M6M+rSTGEiQtse3QaLZhmiQzb8aF8hKZALsG/pTkQ1wd3nWlqPvHUFP
b8tkpRtnMcaV4ahz73kHJ3dJXMtm3lPcuk5ktih4hUa2Qxgc2rzDKr4sutKBrEi8
OUdXjYLyVGBMm5ic3pmgau8xeS4UivlrEjMnPy3bHsg/oJlxuHpvu37lCTe3GnBv
Ol8NVswqKC8FxukLCSO2bQHgXFfzueCNCFf2HvNqG4TWvPflq5gSNZjfqWEh9k1L
Y6ZVTNxabk761/Wb/sApfAdaCIX+Th7v/YIknDV3q4zZv9C30a3WeJ87s68rMSI2
9loQvOGAOUPY3sIL2GIZ+HPRDCyRxhBFS+jbQyaZlCd8WDVMQXEheM+AnWFJKBiD
3x174mPC+Gj0YXoNldtF45O1u5pCgOe188rZCbDGX+pnSzxfzbFst1Tch+Ld4lI0
OnRqjUZx6bhy3hZQD3rGGgaQM7dGYEvkhjbHtgGajAmB7TmsvJIIQa7xm0b0M2pF
BWzCIen1eoWRmY4yH3XLotyJ24exwgJXW88p0ai55RekXh7QXT7WmyHsFM6fbLxl
lkFbv9prrvzQngC8XdWkK0U2401pVJwAMvKutNiUh3P9vxNJrs51LG4Z8dA2wiT3
ECvhvjRDNyeMtiV+tuljLDtva2KJFpQznLsJ+IwQMZSZ0ij7lBW1PMFV/6TWHG/c
fq4ySrGJiDiNViIKZ99TRaNVlSkpVlp7qcS8UdUKvD4R79Z1hDINlUt7cdPXPNM8
yLEyJmP1K7b8vJxQJTIVLAdhSHSH/wGtirTv1X9PpWq0QbSRZl4t+QfcKa37l/F0
Adudixz/zQW6l8ry0Qel+JqomU5r4OFAWcHQnwMHY7vtRQIJwcB7awQF+8NkPpGj
e67SGkM12G3v+T2WTT5BZ8tZ4qkGJs8BjVxBTDGUXIpcraZbW7w1uiCcsMuNCR2y
Lia7u1sm1cA+fyWxYbA1xdnLgL3vuOJkPzubPTOamCco+4b0ZViGKEh+VEcllMjN
9J+YiaGub0/A57nGRlVIB/BIbvXFHqqpflK6fmg0i3vh7LeQLUaVjU7dbF5piiao
9ozKDwFJPu5tmnohV1f7eeRSiV1IacG2aWOwCaaR/Q/laf+Qhx+zv/SfqDfxQE5t
LxOu+GZBfoV81b80BYES4FCc7ahrbplLcNAuZ1fPgA/STZ7GUaop089bNn4D5NlA
MHLR9t1N8yN9e/TieUeEdxCkiwSkVSlECGGUP51aQSJOMwvyT3YMbR8PVS7U5sr+
UNjVtati+LWkQiMiUHSNyw/W+7qbMuoUxhyKihw3xWxlvZGY2BDFlBJACROtrXb9
uE1OeszRWQOZFmiJ1FUnCiT5omChQ2NJQwgo76C+m724qj7x3zLkLDXs6EBELw+R
AR/N4uGsalCtWB1hkcHsbc+IBllC0hUrEU6TYjV3d2+5rVnofKErPbfEywvFh+h0
l7n9K01MbaYtcl9x+w7mtOBUnF7YKNGcEoWQFWwIl54OanCogRl7P1+3HDLkyo/u
kC1k8Db0Px4KMp0Ft4XUDXrrw1xWkQ/VzkN9BKpAfphf5Zviuojdoq2XqTZLg+U3
598ER/hMtC+KUS80C/+WrcOiMLo0+oMu6s/lYSyCrpx5TZc+b0/j70EyLhtFxOV4
pscs28Gc/ePU+VFGvYgchsZhibhVSan1p9InffigK+vVAqoXB97kdo6dLAhg2MMF
WfLUgiPfWXwPrNj8zO/st4MZFJUWLbiH4d/k+1GEsJzpz8nH6C507zcjjEZgWpQp
rotb7C7BbpPiizvu8reLwU4km63/I/9Upy7m5bMEXODcPvt2mpDAzcP5a1NCxqCC
ZdTARU0qksaFG+9A1jzXa7+3Ybo/hlSLUu5M/dOHg3ln7+gwoGV8XjymNiCLlm1k
CQIUZor0CazvKGToBr5r4KTP7nPuBgn0fOHjMgNy58qTJi10Wui9pRIZ73oxcwzF
PglMHT4wWEe3NCOsYOQ9phFI1b/AEDXr5p3bNiVEaq5WUPEyvmum4C3V8U9ZAfRe
woQoqiAf7lXp4v4AtSAOzCVOtpDxahkRr05l+6IzLgf7CVRgLm+mGT4wYHWZUsdI
VsXD2vnOeUC4oCIYM2mq9fy2Gx5I7suFdJRse/ho3es3Ym28+shiCXMs225ODek+
ru/U853tsMa5uGZ7z5hnYwsKMdi+wHpcH/lujhYFDnAGeNWkNSDROZtj9a/P+60Y
6SMrjM2WJw/ExhdsJZZlPjHzDJlcnP4WfqKlFfbka33njPRQvHCwf9Ev1/UjNfgc
UpjulLtUDNekvs7zCoPw7IgB+HnBnuYvS9LwvZYcUkKqWQ7TGbOHmI7wcfsxXN9L
luxV++/40x325JjiFqPy8KgTk5gEO2NiT/bvy9bPbVUShwpMHKkFWjQQpqGCpoEk
IlyOc5a/jsySKRsJ5NjQUAixdRHrbmKxOLwwhdzW8mvn/G98Wh5yVY09v9gxdmwz
UpN0GaqXCiYtIp+eVMkLZ91zXhHIINl7EgYFxs23bGvzfKcAHWveVbhQNqVnRRhY
TGyu/1GMxQCnIXbibzH7vb67X/KGWdnsF0Hqke8HErz3nL9UmiUEQpcMppNg87LZ
xGoEpV57FAs8RvnqLccZtu7JKoLxoB7u8LSc3NOdzUQATgObodhzAw43puKOmkub
EjMZG4gSA1t4WxbRMsZHPa/Tsdxx3RahQe4M1c4egumOzPrZLODXHMRs6Z+FNs1v
w3W4snKDz9ongxMaeEqIvKw3QDuHRqJgwumRI0oOZlrB+mUEB16PxexcODsG+KT0
zWMZKg9YNNQ19+L91S+aE8oB1EzmBBm6mLxRCrGZNmi0g+pO9BvZ+4tJqzMu46ko
DMKqViG18qgpAF30zb9DiSA+Jfou5ogbd/SRl90/kpXgOxIqWwO5S2yzLssoebuz
hTJR9heiv0haO1a5zDhFeMpmvwYlC0yjIDcJEsGLsrRoEohfzBCsGI5w8MeVP5HU
9UU9MJfKW3Y834I/YFvdr7SdugN23fVpx4z4HaIYi6wvI3ioUL43bM50MesdzKhz
4ZIOenLxea8Zmqwdm8QXG5khcVUbZzzpY/ycvgJ2YQklJDF377HDD0tV/RR3GAqp
CWfZ5rqEEEnwUmLF7Hq6Ebop+O2mi5X+/vUZQrkptjRR6u3JqcRPSbjrCGQZ7VRy
vwFKq1dIKdKBREVIsXjDu/G76OKsdNfk4bGpV5cuQBA8uTsIyZ/eYFLhz3TYnmdM
fJsIl9kl0y9i4gEvu45zz398pGJdL2Mef9VhAZYCb4uyaM4aRVR/pn+3sC/y9gwi
vDvLNkBwenbTFgfFukKa7VreRrexnEMGjjUWY35pJyOdjH8NvwlKBTYxrWiBsK77
4x6/hXrcTkyU/ftR6UyewcPJCg96Yr2kLIF9Cz0OWZIre8K6y17u+tWkeOyPMM2r
37w+CW9lGDoRVcBuZs6x7oXMpZhrxRn4QgajaNc8BQIeJrc/LiDg0lurWMdTq8Ox
Ded8d5qoQupKRczIFl6BRSXqGAftSQhP2pygYAheDuWVmndsiqL0oVXl1YQau7sk
QWDrKg3sAfSmWVj6Yycdd+ck+rbv9KFzBncUjjqDt3Z+hsFyZOoZKCdD7o7rSwMR
EEm5xlKsHvk3tYzE29xUZtLzM1RY6Qg5/hIBqq8jmi917Z76cZQfyxxXiiNbU3xq
an+q5nqpQps7RjwfQrnKbAXm6zadF5W4bqxEpXpvyjyWAhhr/QSo98Hda7QdhL+A
+UfB13EkC+zL4LOHaG76sbnAHhDUE1VPLeB7zxJdE4Op48TRowrru8Jti4t3p4Si
zxjD29dQlMhhJ4bFiffL58ozKDsknP67OfocCxkWoUy7aM+EVzdBJBLpCfK2g7U9
Ku6Rcgx23QXVA0BJcDUATPvUWAQ32mZNUflP2vCwMHbMlCCSJGWHPHAXORJh0DC8
MgEvuho55MePhpwMP3pCBSJdE+LzmqKi74JMPcQVeAeVKRuCLqzH6EtLTfYm1DTG
pZEBR2tVvuJf3SAMoAkNmPC7wZYCfQPAF6lG7rTttRAan4BzZ7svFkSGMmMhMZkG
TgspGWJNYUxd1s4loowwzC2NJQw22tUhgtq8zEG1qN6v+0MbgtiImDj5bO7J7W0v
QgPCg6kU1G6PhyDkYDYN/H2eUX3APQBrmAwiWKOfR2GIu2cinh7TWX6VG59YR81h
eGi2BD4QOBQQDvVxgiqvOB3DH4mRoQBZUCO+9TUXRzyMUM+eOCFwTojkb277DFSr
b0A+Z1S/+LrxnNLO+Oxt+1YDscuAge2Iew6gV4e/VbgN+NegQ5ZcigHmeRWymP5s
/zLnPp9e9oTqIquh+CcQTXFSy3MYN06Rtz2YCxsyZeGQuFZC/wptHvLQJxvodVo9
CIrSE5Lm4Ru4LEWaQ7dD2owzGHgsMvMzemC1MQ3hIOwQp3L1QNOex342lpMou47p
IwAJcpPn1ez2gH3RcTTdod/elkGthBSxehYkP7Q8JHNCaTADTyybE3XENaw2n4Tp
SK8Z3IOEdaxYurw39DO4bdNdOsfx7HOsDbnGbmWRjX5kRLaL+R4nONfyrnD/5eoC
+XR2zQKbWoE1yCcJS7qezHgH8y+nbwAxeixprf6eXHJdvGbvVvUaKpd6TrFLAOwX
FTfWVkSCwsSQ1HEvC3Oc0J79QTz5THksA1KB9TDUsSnc9iR1nazpAEq8nycrLfLn
XqqYHf+ex/y2UXfSy5tCe5jPci9sai1YgAFUIl3xPEI+MdrZ897dieiXCHo1Qsuj
35L9WURNwC1itJ9HvR3eVvZn6gP8J/M/O2gu0SKYz5qnDhHnu3IBseIQloB3HrI6
uTYwaGO67YWNYse6goKwBvYMKgK/4OME3W9FWJJ5IeCN/N37dkCXMCejtQFL2Jdw
M4MAx9Vr8phlsn4xShYFtqLxZb2UYdFr7c8De2HcHVsC5Ib49OOjOsuJ51OU8NiU
UiySfy/3e7m8YMSPoyR34ZzGL4ocVEGNxGmOCwUOAk/MURXQJwOf4IkqIV+X6bYN
8B66faDKQFPRtXk6WZEFZIi/iiKnyaOkQES7W/Z3UK0HltEfN+S03HFRme3vFDnW
LWffgNVbANAkf9MDljrBAHrtLcMrRdUG/GAakYh1omKrSW4OidY6HT5LfLyjI1bT
OIcbZZjG2q9WaYCqlwEj+RwaOzHTBjDrfGu6NHPThkPzDhN7rH7nYDMxUlatNsoO
KUx4lmp8nR0ZA9aHFfAOfp9+MHjHoZ2HLAnrh5EHpZPqX6fTVg1vugRC7/xQhMXQ
KDyBeUFBFBiqHPUtWhsXoNOa8/m6qJlEQd9zmVXkbJMEYTIWyiNGbu6UQOKEJlWx
ptF0k62azAGtFynlx+A3+6Kzf1p5LnIjHGqpKAZuF0CuVxZX39YTYk9CHETo4qtM
E+NS0V7GtUmb5euWXoacTlwSH2/6nAwZLd5EUI425pWTPxt+L9tVjf109Dtsow9h
JwNSf6eTiLyEa81i9IeVk9eoRklJrzP972FVO1xJ4nqP6oyP8iZVHRbScfxDR7Gx
1tW78FxguTY920eBDkdBdixjpVUQ5nSx0pkudw5KzrTCCczQnCl0AzV3UGPEEpsc
qAUrFsFVwBMm7eprMknY7AUF3/BLGaRm90VaxENu2WPCJefsWYNz8aLQEo5efF6Q
mxO4QA8p83TDz570kRen1UoCcGSai3jhrwvRrkBjZ3BaVo9GyuP7J5Q1SXLeyTqx
PhZpeDBxJZ+j0NxivQ08JkZvBYhF/OlyvZyMHRVBoYbaN0uuAhEsKJjgE9e/ulZG
pS8u9nEGOt0s5LWRP716ZHIRTYlqLmFJeBGZ7/T6c8HPiDDJuUOiBB2/adBlfi7K
sqg0AXhcRWVft3ww0gZdoEswqRkYrZVydxaO5YPZCKkPNCr33AvhcDhHe4G6zK5l
uEZeV/gLFWEkCENrMhgUwcYIl94Do/TFsjAeMR2IPlzhAtfVU+KUqpSYyFSk4Mev
6b/9W0xBhofHjlWEbdioWec/dPMydzBHbj3C68/mNb1jJOrfVpTHX/3fLfICb/0F
2qEEXOOCU1mRgkmbHyO6ZcPWCLRhbCa3G2p9uMWtGdp1uMg0/aG/nJlbodgPaQ5k
jfi53pkWuYp1VsR5VVoMRWqGrlatFtoS2mxT/CM5RzoMLYBFNfOI6cmWK9YQ2uXO
wRi/HYJfu6PYkI7miW98W5n7Y2LqksLGincU9HqZ1kNPPCEuxmVyAp0SAx0MTjUn
w4qBHsDeGvpwoHgCa3tcZErfK7D3pnip0wzIsW+6NzXoaOcjQq0XHsdoRgqTPlb7
geArjjMbV7EQS7zdtkp6ZGzjMC9vjnyLkxBt39Wx0K7CtFX2EGlnPW3tagcDRYiJ
B4USQXtMU30MYqAOJhGYWP9dAzzz4F4oBFOUNYCNazjLv1sNARaQu3MlujpDbiIy
hFc60kU3yCcXoEDvuMHzh6iIRUnNsODYTGDTku+cHJx0yUCOMle8riFF6VQxNIPu
7e7hQKOXay6E8JhYzrpqCH7uql3gZ4LlHdN9cuKXcBH4vlb5lhO/RMk8VZdf7tnO
zinbgHe5hldjUH5vu47birAuYnkyzUHrT65RqU5LNIWlffDC9S6TA9SKHsYDJad1
gtgIsWmLLuX2etj7UMfs2yNE/VuXeszTgJH9ThR84eDnBmuDJ/BD5//OJ29LKm5o
LVK/l5Sjgg1xxbBDeWRFRnre1bysYKAQu8EGJZBNBZ10FQ1xVMKodckAe+hGW5Lk
oytB9CQpNoPMkRycrjA5uFEsdDeNxi+YslDtGpv4h4HnyVaqU9EF8BBftTOX6mvE
0SAbaRBO/1QK+kn1ZPREQs+Jyt0W5bWu1Qs57jvnyUqSj1dZPELsoM2eqQlfA6ci
eVyMFH65JK9cj/lpHq4YhjtRVukZJmRdh/lRstkOQWJWgc0LIQWn4sI53uqRw0v7
nl5Uutahy1gjq/3FGsUIHkSol44GphIBbKMcbWeVagKhEDUEwKascF62NrpQAj0f
5+86a2Zx/sg2dPjI1zk4D18/d+JHt2q0etCE7pqyHBUyrAteoDLQfSyzKD7TWWzJ
tAF/EingWkJX3jHs/GGPhuPl0zi/wjwguHAQ7S95nQ++ytMN8elwrhkWzoXh2WQP
Wn05TyGSTdaqDZvK+ycE97pNFZuq/qX/rr5V3DKAER1/ItKtcpAcOzKilUrnVuZT
/Kly3zvZi3xIoZ31kjsdYk+VEQdfMBRpkdHpRtjd6tULLr9TgMA6jur6+QqANIBc
/koS9b4yog6j9oSgObUHufp5xSccLhXShAwbKxN1LO+M1ut0o/DtTOHEWuCIQQDa
52WzaxsMGlFb7LpDex0KHi/IkpRuhMANKK9lUGbOSTUo8Cx3b8yaNOSsygPDEh9r
QBVd2KbMmLH6Ywqbvg901L+tAHaKn8oO+lWjVgVZRFRp1yBNYIEsEl9rsIS7iep6
PDsA8RL7Nzx0UaTUHtChMB71red+T7zmc++g8V8Xb1k3RdRZ1YpFcopcPD99g5ko
qats7JTW5QbKN4M7XPYtST2VdjGmtpcc3V9cFxX/OCKhrgGxuUVf9rb0wVDrj9kT
u99XhiX34FBYQF6dic/4tWjwa2EOETf9XUcsxuVuU9D2yKW7p9/Wwu5xvidZnZIj
PaooaL4sy3Bp6VKjT/7JUcgaY0/LIlsPoHTRr83uCV29ZHErvxvUCi53n+z10b5g
zS16xVZZRzHY6R2ycFmcrRzf1nqUF4yhoNNVCxtHyQDcPkdyoQxPkmQufvX3R9c6
u4OLAQIE2w+fRUeq+dEX+nfZU9qPUZY6edd4/yvMIiJkFBxx+kvpyPBUlghzv6IG
yRv6QbPsXq6ARWq2G2Qn4g7vhQ2eVcQ8cHAW//8w20VCrCt89qBIEVan4VQ3SIFV
j+Kbegw+suJvy7Tl7JNAAtWoy1ESUWRbygvfpm38AKdSD1yu5SVYpj7hCrjImmdq
hIylQ+FJQ2vXq7T5x+TljlO7froUhNFpRbVsll19u0EAfb/6Hs6SnIJKg7DVgdhz
XgWNtSfW532nJBur3Q4/VQme24qxAakUy/cYoiGfkUZ61AfOpLKCUbgHJD9GOHTm
k6lqeU8Au5q2B0SV/hxbNchzCDcNx2YQES+RibXTk3tF5d5B/umF5+fT84qpiXSx
sYfaU9f1lkWeyZB80LHpONRnJXrMWKEhyvlfxUF27NJzEVU0spVmvYEVpcT3KnEs
FGh8yzj/I5oRMoZoenFXxSRE8i4kJVuqXYlX9j+i6EV5DiYi6MhB9LxbXHLcREBV
ON3Wd1JXjda2Tne9GgKEIevOV1p5VXKwkh0UhUAWt1E4or3KyHQNVCIvnVdfO0HG
36qnhEypkUtmJcmlpJD0WvfSDjQhaZMbsHcCG3qq25E0ByCb/N6MzCzrDv03YS49
J/wSK0KYGYp7klP8EKcslqrCLI5ieu9QY9K8pS7SMJYwDrE1nb7g9Srd5PVwyKQv
3ruW8H28vVGUksmJOHWhWDFhVSyFbyDHQ7q4sAyIIFc1hmA9f7fC/e0F4FpjQU8j
d8Pm23wYQgzfkPNhEY6yDMVHjdAfH8FdZNFg3aGYeKGk+iX+9tIy6s/64NXc/R2i
Epgd26T8mocbqa6Mg3L0Zx6nuaKz8w3TLgGC26/DbWIJz8Ajy7XiyI3lJ4EAYwrS
K0BBEaDA5pAGwrMMkPW/0wckn7/aCRfTqOZiuxnuGnCBLfOgVMTR1fjodw/OooNR
nd7d/YGJh+rQLYLm84XKsV/IoGutjQLhKbN1w1TbbiDjIP+Se0D++YMFORtmD00G
Y049+grJyTQ9MFvogjAzkM0jWgEku/5ZQnxuttjWdMJ1LUSPuPrvERZ7Mc1OnV2r
uASZpFtIfmd+Rujl8yqK6dDcRbqC3l7jDoMbm9PenCHUFibFxYgGB8wS5dRTUktv
pe99v2iu6JsIoLeM3cAweoObeoujxyRINDnkSYTztDV4tvwAYcM7ktErE2jfyd95
oMrwqvyTr2Cym/alJShQe3GpOyKO+llh807fiAHCRfi63xdpSiGfjstTmvAwKYM/
U+1sj+6DtD970G1bxSZ3mKrdBEfC7Ome9XMDh+vgO44cQ7gNp1EPbbVcEguMLWth
YzoCkSygTp0oc7+onWzZarjthfXcxPtz1FMBf9QT1Ds+adsHx1pumxH31x80RpdP
hVDXXN6CgMKAwo/K52wt8lOoyUMPL29LkKtot0Gcpg3btSlh6lQP8PhYQ9+S5ciT
hafr4jQ8sjCsiXq7zA6oXrZe8LpJdYg//rMJvN2GEQFZaBckBKDJ/n4GrouUlvel
eZnWXtbaOp9H00p78zfzkkwtA261HXO+8ZL64PiS0nrwPDyMbrRG8LRdJjaZFo/O
U/wob88/O68lYT0/LlKXTaEVfLRkCKWsNRZagQCwQHTPshXwfxFYH52n9flbTLgl
ztBtH4E4KXaACVRRqNQM1tVQYomp7p8E12cVLKYkL7zFlJiKz803wNKBKO020tGh
IRusDHWa3wp6idVFiJjP3cwGa+G1BOn4i545nYdDi3dcEDDScKf9n37KF94vwVjL
oF0bFH8ZrJC3h5nzKXowsUjb78qMndA5xIPGQSp/8cxrb4dCE59Gbj3x90M3MUKo
TzFMlOXciafSvmiybdJOZCDIs6HhDbhpaZBNk60UjiAHx+gSHdeaat0mpjXd4ivV
uu1rkn/eQHdcUv30xt31f/KWEGZQDW+eOLRerjTMs7gK2Qr3qro+1HpWUpRkC0f/
IT3TJcmMf58nvlR66OxZgH3CjHzx4xtEPJ09XxZSBHQoJg5x0TZKYsPJVangNI+a
x9cGejzPTEokqhYrGbLh99iaLucvCnVGQMpNnzr1zyj8Op30ZTomyjCzXNTAdIef
LrsPXUHUn5W7r0QL6FvJzvUlS1tEjD8GYKqUXGzkxe274oHQcQK7Iu/ljLp+CU/W
p0er1gwPtFAOAcXrs1Ef+QdGQ0vWhwsKgUcu5zuR3b3nOFUUIzcpPM7Mf5fIorye
WJQAQTFQI0OCxLvPu6zPHkB2Z3IEH7vzesAC8uzPcvJ2vlbF71pJ69yndohzz8yg
wf+/erdw+3gm/YpiS93otMe8vchhZD2WLzeCSyCSfKiMxun3pXXnlVGRGrEkqqPK
KutRWuamZJF7t9HI2AwR+GURxRxL7g6ItRyto37astgIDPfkt3Lg3uR+li3EKw7i
dCpycjSQ7wd9gfA9SbXITssswMARtf/bSiUFiD88ExHazsDyMTboxVn8MARc1bLT
aB1cS/5bmAYPYy7sDllLOwPEMPqCmsdiT3Q2hAqkcx90Zr2aFEk4lDlDjQUfBnny
6/4UtFAUyzSJtbtFghcdIpxPRa7UB6hfOTKWHwprU7DUy8Dk83DD3Nt0HFAHZesB
VACpECkr/xGaPZaCGLX91bR4BPPtCOWUji5M7B4TYQDmli9CO63uOSlBLQ4KiVUx
vJpkhqVfm9DVpkOxo7Tc9KysmcUAD/XEtDKvC22AqHQrg+J1b5BVcTP5PSKjOmAt
BdWdPxaeKUUYYMmDMNi1x5QCkjYWhU2Hb4GvBGUTb15uB+vM3WSt9gJGFnrrJcgJ
vw+R2YJwh2qnqHFzhE5uBz8gc/2JKKqrFy3o97FE69xitaZ5zcnrPCxWviFq75gj
Xsfm5N/eKaYpuKXz/Yrre4d8fiXTXmU6D3eJEfhuXZ8ruEqQoSZx7a1H5b3DGfDa
2OOzEQqm14w65zw+2SuxCdl8oBv0rGzTQ24uTkd7eUqCZZTokvyc01KMsG/yqoUA
n0/BziGdxGwEYD/6TiW8SyWhf3b6tkuIsXE5Fp0IC228ts/SmpD/995wZlCNcyks
itkDup95f8lz+kiHyycvXd005RxUnsvRlH6KFyP9mWy744WhzNii8nAMPXEeugsU
sq1Ere9UNoWAuheaqDB5V5RHLpgROAyy9EZ9IseWTo466i5YuaXAjwNKqfITW856
lM7UsGlVEO4Wk6ehtx8xqXSvAkPE8Mke9zqhYh0WiP12Ci+UXSpbZ+cfk5YtCgei
N2vO8XcpJGqIZKhKu4AhVfABwJry0uDmkSNXPlq1xZcu2vkBc/50CnixRZZuBCsl
IU3QEPniyJwe6BpIjyfOVjUkn6gzmWYqs28Ignma4gkQSxKkTExvQT0AX1KZPuKt
m6pMd7Wl6YoFpJTtmg78c0unIF50tWcjro/puHyaj5iamNz8M9+DC8gzgEzcrAoy
VdKIeCpT3soQqibd4kyEAsXk36OebhnkcTv1Ph/iJ2q2aciksl091ZYOjyhb26oc
j5u5Rc3iIhBQPWU4/6Ro718pq6nizxm4LrshdJ3pX66BK6p4MA7p8iEAwe09WxPG
h72gYN1EDQVqIPtTzeMNWhZGKiONW7VXE5XiBl8436ofwdioWiwV6iwlfQ39URgX
TCUdESbsyFmnJJ2OH5IeeLWQ8xIK3AqY4rp4OV2FI6bq9fpxthJxxFlPNhih9w61
GhyyOEztwvojhEt2+hH0+M7AqNFUzslGnOKDK3RK9X56xEFVGejdWi4jJiXskGm2
oDeBHFZAg6Jpl9Q9bvmN/BA2zROofHwrZsD2Nxqyl0d1UNM4AQqEIlT4lsDsw6E6
NcfiqiZiPU10FBlIwIDIkoqHiBQg/b4PmXBlVPi3IA/644xiBJyX2HOuvDp9GWQ6
WlHvk0ViCeq0F7nytO5VaqbrGmDSUx0fdLX4izJAbhVetOs5scADqYklvT5+K/j5
OY6gwk1/6cecibLEfnXDyspCUdILl35TptNbEuv+DEOfjTdHchZBiYli+t30Fsna
arp595Od9YpS+WeGdAUOxER1VwuuDs8/i4POBIpiTB8aX4wI4tYe6yjjHA5pu7K4
s9Bg5nndjqpjv5uziaTqy0DLeYGbd5FPkQ9up1u9yNzSggTC1XU9qYvbW3XSpNCS
Ku+wfrd4gDUZwfJcCvilpCg5tDgXsbZcyf0xFGe0fOSUL/6BDvHKsnIN1wMxkB5h
8mkMM69brsmeSLKxEnlIxY3KTzVa2fjMnwb+Wjks6g3gMmrpY7qHwZz43ROvh28o
+moUDQOR8+Hq3wUzz2ANcUQ7fngBtb5jSVV+pNPW81AnlNR/XvcRuC+YJbNbGzzQ
0/ZS+0Xk/PumRSQvZ/RImcjXZeg0BQ/wg1mQrFVwgB1fhO4ba4E2HOmGWmYnZrR/
bGaHW/fiIMemM4RIwKuqR5H/stbR46eYZCXT4Mhp14Cdjj9Hd6dw3AXSfBwlws0d
zx77DdUx0VopUVnmiH6Xdn5mOdqx4FhwvOe3xHVaDF6Sbw9ZPQPJIUkOHjfU3s1O
yeOkURtcZUteFx3BrpEukvWxS+h3XaY3Zvm1svQ+KFPDOcvAeOKecQeolweinmf2
T2kgtogPgW+AfBk3v6jCHvA61fP3NpWWcCbgHkuohfUpCYnbAK6TRDgRd4W6ZAUM
qrRieQk8h2tnwC+UdOvmP1ZhlBzQI+6nVO0Ia2v8yy9cBo/Qf4B00cIPXdSVGCmT
7asu14TCWFQeF9Rysv3nNhQdH3enrompoumApGlMqRLpOdiKnUINCnJa/u7aEIAc
KAp4xKsyaYsKjmAbCAuktAvLT4VuhdGa7NBYIT3PSJbunuVyM4ihbs0+Gsnmf43+
9ogtWzbp5CwsTSeT/pGlNvpuXoGR9o0srWc0w/8qYg+ylJkVlBmZkosv4HK5WiAJ
QTIzZR01+5KhrqvJv3foFSYK/X4mxacMg5dJONCzx81/WNOeLkCvPXat70AMDPUl
MHXicxfHSgiTgmfAArhtF3u2rhD5D3Uikr9Xwwryi2E+Gr2PeLLNIK/IGz0rps64
ZrhhEBy0/XzLGTnsMgzkUwc04B40YxP3auQGqwyUIliHD/EXQ2raQLU37DY5NfJS
Mn+nDjSpBYuFPU4HgQSHmHHC7iLma1ve8n5eIfyMWt2yNbom8QhnmJc+drrMTfv8
nK+P3GPUHXOBVGwpWXEZLoIfK7lMM1sjfbruLGdKI0f041hjfP51gUdiRB+Nol2r
vR3BFpZMUgLsp4lgc62tg3QoKCXbJG18aWmA3CrlWT6TsZaGGdMeGwmARYCK5g5y
2HBLwvU1zxl9/yHzMR+QedYDBKYlGEKXOjxegByLF4b23ehF6gOrqDGvrhKkx7fm
d4VZNzeIpXU1ZfNOOUIZMh+c47O5d5klB0l6PS6S0qcgXFj16SY0XlO1IcMb3L5M
KGikt7OaSVeuGZn9J4iMCBcyX9BKMBitCLHzxz6FV/50jMbpUXVpENMvcE6j7mwS
jQIry2kBu3J2Fp00aknUdoM6YMk+QHJlqVscjDO1nwbDyNhLotsTehgbP06zZQFe
buVdfLslJXl8N7EdjQHWnSS12j/ucfDF74goqmhm/HfXpURJ9FvXrF0WWlCZqP3y
WqN2spJn4NjdttuoP0t/v+l2X5T4Bsk80I94b/iybnYMXAFk7k3vI+bxF9m22kiL
AMnk405Grqc5TXdYerJW43BuaUNBhH6d/DebOuLCNboCtdMhS73YK4j/Xwj5zw1/
vO89XiAQT6GbW6bwt3NNhLimvr4MJlWHeQbPgrOIhOEbJ9Mp27hqeNBor0uSeuGn
3ROYKMoOpUHne6arD2RSLmXsHK7w9x2Iz5zsYkNU9pwIBeG1wGDPbwkvl9uBcJvJ
VQpl4tAYn4KRr7fi0ySyJyWMqSS4Rfh4ZDn6oikRavE7BK8gnVOT/dGszHkcawyf
JGbOh+WS8GnQpG82sQzImWIk87VfKKnu8wnPxnkhAMnqWUKrNb6Hyk4PqTfJt6h2
hquBvwCIHB3E0MA8W5wkydeCAaXj1uOnzuM6vfzkMYB3vYUsw/7bz2voB+Tm4YFH
3RJ6JQV+sbw+gox5TVXMCNd9+bH2ff9GxD7nZG07J7L7Ujiyh/E3qF+KgOldCxbT
CETCmNdVhcUVsjiK1r3UYaWUPrSFw/OkRF0IXAWPvRplrs2q3UV3DdrNHaAdrdl+
B8degjW1tdpy7kgJcq65Ay0jiO/r3mbNEzHqaQK2arZzVOsQC9vWqmtVdZX5VnyS
mcL5Lemv9pnd4fki2fRcpciBTU6m+SCbdAV+lTVj8Uk74vR0BQf+ZbkenVGQ0TKB
ub9FfOPySL0Ik+fWNPI6oICGb097v4AwVUQrtMYel4ozKz+3Vt4+fzStE1Y2X6fx
8ssL6/mPGEUiMBpLO0+H/xE5chqXi7wTItk80/yWvXc5Zo3xsYbBdI4AkraM++Fn
aX/o66pW9dib5/M+LsVUKXA1Y0xoEbbdJqY8/HJ6ovkZINd0AwCCVC/RTkF41d4k
BL4+YzjtntJd+O4iq1U9HWW/7t6Ypj/xBCOTfavXhJsRYptOVnrTBpqVXaatKsoF
IVsw0Am0q65EOb1uVivp+VIJX/JGSoy/9AveBGbO2R/HSvA1AF3f7Ono+KNLkjTc
qFzjBi1u4nT94EObzQ8/pQAs6z8/wU6hxcXHD2a2KdeM2+IlGS4XC2dXmDz9enUN
uyK49tIZ4/E1vMwjgEmzpq7urY8I1fUxvHO2s+xH4IBiG8PzkxNC7Cw4IK6kLXzU
lNfiQftkpiy6C0vNvlNTYFOIQSsj3YlSqrutPs7MJ8YTglA+NiiDCrAoFIR8HhK5
8pym/StnuRMwbrayV+PJ38QuGD5rA9S/M8UM2g+epH4K1GX/zmm5jVTYmg5LNi7I
hniXqkb5vG7kuuM6D03e38MnkerZ7sbcdjIS54wdcxJkoITdbDgT035/k+61a+39
t+12PuyB/n+hc27ofsIg6cXdSGkQXK4w4GEpHok9ar6+UVFSqcPAsAsWwC6uuQG4
6/2clNRHiQagrSMVcfHj5B65Y+DeYq7UnBG6rq9TpizSmF25xfrcDzWFm8eprqqF
r1FdGP2Ao1StWfAgEv3rktwQkngwCLWi8e+dt7PI9Sj74SVjOOmS394YunEO1HUg
rPV37f7+NgJAi0kabsVi+VFhCH94Rf0TdbVoeahl/i0CnRgMPADE5SOy2QjuOIIo
4E7tZ6lP3g8C8AvNe4EOZ+F7a7eub4nhxsieEZt3K+f/UOoS3f1g3cGI8887qP6Z
lBQz1LvUbpEopCkeEm94MJ/cop+FaILnbLc+pvuwVSBf0xPpxBXO1NVOyRz2U6J0
+XeIxpT23mth/J+4TK+wpg/48tUwXq0qL/RtUR8Gi0UqVBJJXovVDyuZgBo+9xgx
w8BZTN10ML9cqUbT9XRmY40OJ2AI3XoblIlqdHi4PR127rUtX6DYJu6LKCHgi4uM
1CFghgBiRIocy5x9Iy35AJtZ6e0XdIdmQSDgigudfuwfx9kT1IuMWvzEcib8XBuI
cZv42fnXBIWHN9ZGQoNFWuUoC8O+WOq9YyZG983FYfCT1u53KTDCldPXlDoGhwtn
tXmmATYzeHV1EGV97Cg6XPpucx7sfZZwdBQJEdXHQJOagsnKdWLYCzrT8lm87Tmp
tnUf8amKiAABLzPSWrp5XI3yrp0cravCwXCon/4LnMwFi4X34LZ5hPBMcO62SnhY
6hMq+wauMwoLY7ZhsPnmblPYL9F1T2M35kA+IvDppexK2Zh/1aGjhd4VxdZUpWex
9YzlNi6DjGI5MroK2uFdbE3P/urVLQ2fJrY0mHEQWdXldpf/rHezDKIkYpOZ8zMh
CF7/LjMuJaSYIrEoQmFd4BtOBb/4VrnhywSzA9iMNEVW0R9jGH1aKWdXbLTr4KR3
FVw7reB9iabIsd3CVG3VUrQoEk0oADxMIn/+U8bT4o+VTS+1mHbOUvLohnQZsGzs
icZMztsaVwQlhZwZsPHxSeVIcgxVvAe7BZDtrgWvkaWVmNsSj1jE61ma1KpbhDci
EC7o3dNzvbY6qs7odE4Kw9Q5A4WRCC3GY+7M1IgfZDmL/L/PHxZyjzJMIYMjGixm
ADlWBEk23GeK45xHBmpghD61D+Q6eWR/OaUIj/j7wl+3VhduojYG4tzvZLh7mo48
d43CdcoI1qHeHK9kbKWVE376vbc5MdG+zXVR1XkibKbZGB/DuTFdk5jzNEZ0B75B
WDxurk+92KyRnEFxxbQsq0NenQCok2EejzyR2va1zrVMLWpjStgfbGgM0e0SzGR8
OmNqs3dNWQ3iHB2tWzmQP3IGMNb/gPoaQTQxV3DEr4RcQikrOp2fYKoaXdP4qcp6
Lm1EjPz8BAfYQpXCgdeQETjzchNQRZTiTP/Tj1L3IgF5xV9qVcbl+vDrDlXq1HD5
WMXzCUXv6RXZwPlXgivJCJlXnXqsKmPedsQYIj4yz3xZH2hEWWMYRN6efy/HnXtz
oBDF5kIIyKfKs5+4oLyGV8Ynuz31VoBtF0AjJh6DezbUzvdP48Rr1ncbb31L3J1o
aKKzV2qmt7Cp14rndacpNqumdZkckQ219jUO9urkk4+t25BMOko5i2ye0hRi8z61
uRJgGoAGSiJhMeiCM9VoDg8v96voXW3fY1bZFl5adolfDWM3GgvdmVz3wr18QVOo
2rhN59Mk9iN2RZxi2EuHrIsoF7k52ivHMezZG8DXnQkUrvVPvH+OYeQcfK6WtE40
ePhZbkEIzEQzY1dpdVAIQt+Cm0lK3BHU346Va5+bWp++vlY1Igd7tzf9jJXMFIaQ
IEQYF4nWdr9I2oFPL5PrmbpVUbbOj4EZwpgZ3JkfksCaxp0oDiS/KwEHMEGzp0xn
7sBOa+zuemoZAJYKCWApwUSdX7iQMYlVBGAeImTADiEeMui038WiTI9shctTz8jw
KgbKAugSOb3Kt5A6VVIdr0nGGYZ1o8JM+XxfDkuwIjhXG5UgrTjmlSFrLb8Dn3Wv
s+5MwHlbzniwQPnOi6VtszkkuDLP7azjzsQF2hG0GrnkI8aGayHFJ2DVzJhucqsq
HF/ZxUbXpXMYyfc3dD4lFuarX2I52gzrFgFO611OTusjSmc1en/lqamGpoRSruzi
ApGEYhR7snOyo6Um2a02A8Y/5avYEEM1odd9QiHQUii194C3udeOxmIiG3Sefmqg
1leYQ94q6go0QapkorMcA59KbqpfiOTbox3hCKqN2HU918ElAzGf/Jrf6jM3KFe/
MFuj+hzHF+87HfjK3HqL/YzHXlpM3QX+2uZbGl6BzFKUAW0cROoFg/RcnpEcq7FW
7tTORz6oodg9wpNxnMkbru4b2gF3QT87P8IvvDp1kuM6FgX9843KTDBto2I1fbiP
rXTY+q1RbdHpI9tjbL9KOyXlJY2udAwPKcFeok9Yv4i+9/SX1Y/9ZhDrhH7Tpp41
dwiOW4MwOmVDPrkKQP08XzoiiMWHU/yzqQXx9MBqmWve42/JQWdKD/GVcBikF9Bj
Ru9FKct8sa/BE15XCYGeR21sq1hyXFP3W9GnHf54MGOrTcAtHbmD+jFvbbPc33ch
Blt7nYMpvyUhxgIG6J5kZ8S8J0ucCxvNdDzPsS2rrE4f0aRYly5JRNN1q0XjAz4H
I5KRfJf+tzMydvKlQ3ODqC4i7OanRCKVmLYQZYTY7bvSNQuz0oMncZk0EBe3yYsM
5wSmCzwgTEKkSwHH2Nquj4r2oGGDj5CSCuvdk5obhtmYj4m6gFUIrsuh9DgAXJsF
jDmJ50Oi++5Xg/FzUWy/tc6oNKxdphVt2nHMbQgqXPNT08Z26J9xHxmhVu5GB8AR
Kq8HDGAyV/QUoNgAmUlaEIfrVo7ZOxgQ/Sing+YQXEF0SapCtuplQVs+hCAyRF2t
E1r7vncYwhzdYgZOOzEAxdjJrkpMZr567c8X8FnK7hbGI0jn01GIx+OSQEDo8kar
CTNRc+pwlib7m5663Cs9T7vWyMp/4MJ0gX6Y/9xOEc6+0UOimmuI1Ph6V2PyxUGW
imC4mCzH0R14EiRVMt+QcGVULvp86Kxq6uu7Dzyc5jN3cntoVLvWnwHm+uJvWazo
T4IKO939ja6BJjYEpp+ecxTf6EWCNxKJhIufkVVAsAKfaqauDNhoJDUrqUv7HP1r
z3XYoK5sOkL+G/7hoCbnBKBCFw1XbwndQG5sdHzIWWoOThm2e/lPTq0CTr4KMSd+
B1JS0Zdvxfhie7C67DKEJBOrgN4AexWnuSvkkMvOntELGMcarb+ovDWKHHTQz09W
TI5EeAgdITzGQXHkYB66pq6fxjf36qlrolgVnxIZkjXlxigYkNVsLlBTSenzH+AM
g2PET1sorku/7xbB6J0BoHQ2zMaoz9rj3/9k6cgQs3yxV3TFap+FFqd8wvJLU8eM
K/TMkJv4eGxPgOuowGaIVgcbL4GPDhSCEEJvyD09aYW5hj1MmYKuUx/fw33U9O3T
UhNu8+34PZOCdbM7Up7LQbqPIMR0GVGvjivAq+2Ha+L14ZX/o6mypC3RbIhlMC8y
TrNoIBaQWLCkPrs81hMJXLr5yfR6VSEEXgal/jhugzC8KTk5IM4Kt/yzQdgfHYCk
Xnz81iYomBuVivykMMTaDWCOtwgoj2jmNS3OMcc0VXVSiAqnK1BGZkEYm/AzPGti
z86mDgWn9+M3tHq4NPjA5fDJ1wHkza/II2w1LucYWen+VAKh5vc4R6R6ILUG0lps
s0IZO6GCSKU6gfXSJB5I12WcE3q0k0UWFLwH9nMcD9Gh4MOYyBUswHj0vkPL49Xc
2IhSEWzTDonO9HB2Yp5C/UeSYe18C5+nmn/Mi9yGAocn2CthHp/3LQ6+KpZGGpxN
Hw4Rw+v79Tm/e4uUqaRZymUWSilpHRPmzJXdwxEFQgibXQCeAkv77JLrbWHmKyHs
0EA4rtBV26HHJvf++EhqLwCHon94gFJwbyeHVaEBDkzDM7TMetyVueHHYvgPx9dt
eZzHv7A0kL5qiVpRgGUAZpIxyPysJNz7mhXgJXGIce+Caow9Yn02nxgfq6A7KgJJ
e622uJaQ+CpCqmyGB9P32OuwPYco+1Zy4cl2NPLn3FwWCtf9ctJJKXauBUZSepEm
u2LVUvT/1JObDuAHvZmk2+wobj9TeOR6meNatujSu20iFwpEv/dREX3vkoV44qnW
YzqJg5/sZwWCk+270895MWQuoVkU/AU45bqL7fJ77IOJfYW39TIU6jPUtAsJkbJa
ef/jBDacRjS9yeY0zB/sg5cbdXFE0SRZD19XyZLdg4PPcoRzFh0e83SvV/2Z+GVk
iR5uMvJLQuK46wusN1i/kQqQcVfuGAtIHtZ+Xvs3/Y1wUXM6MzEjAmkF6hqDuuy1
aM8l8301C/f2stE24RR8Ge3pDVtjeEmTnczVszj53wEa95g704dP0IrB0ofimNQ9
iyNa8FdZoWK8D7BF5/zhGg/QUb8n5Zgv+yY0fkmwVfABHXNSoTQqX2OwZyQAIjo/
nOokUkMQHUuOyh60Zg7vY2XqAc1GASezfinnhZNFEpE55psaNvCJ+H3KIGEyEiy6
XulWNgiEQCj/Ar/RFZa68v3BF/VLRadToSNPFjMyizxOGSBzyT07EXG+hI1lkWlu
W3edSRiy/72qFszp6uiAvukCzpYDlQ9UMpT1sfh+11AdajgzianouupfDkHDZMv5
oGbAqJlk+iOyiw73pimXi2P1x0r0htouTBLEUs8JGrKFbNkZbUNWLscCYT/xNHqG
pAxh4EbcvZAkLpFEWOGB6EWaeIgXd8/61XqGDs1yfU4kyTHLk0iqeOmA+oIIElUO
itOPpxE0I3SmmEkXsvQ5tftfDSfKJIQbtdH+UHR1f2IFhKb88pdZSeoHDAW/wu/d
1DVCMPz5POE0anUaeacfe5wCdagJjYXjh1rvZOzM1BIXE//i9RX8XQUWG2dbu0tO
r/JlFz3/GHws3lAmYyZLXaPjNdtv+NayeOXllvox4hxYX+XhdBBhTEsxa6qwdpHT
5gn9OfC1GPDgZ2isIdRBjiG+M4L/EVRM5SWt7spPD6ktCd7/aR217MfcZbqWfn1S
dSX72nmJWmjhGjiKu8thr6qTyAeWrMRmecPos11K5k2wjWfUv4K0W1pZZQBiVASi
pme47f3bFIG54+46eDlXohsetQ+K+rCzbwXWKDfTaLR6yBWhIIzT0jfC62YL0Kl3
7nUrQ+shh54rypTTq7MpcZ+tsSH4df9zliWM2xmC+r6lWR92olDVspI0PhIntfVm
DMofMc7LdShMsYT1fRehoI7prRDJOd+F2F0mhisKvLkijRhRBAvfFZDPN5D436hV
JbrMaWs9IMdAYLsR1F71tDtHhuNSQGArpF5gdlokz0s1P0qwEF13j3G2NrkukXGi
idVLFfUlbxAc5xD+Cb8so+zO+KPo2vxfvscvp6Wwe7l2lnmp7STqljv4st0URMsc
HqUwBar/UiRcrIRlfnrbPRRKNBkNMUiJWQkLeqVfmZLYroc2PZGqtFC2GBYS21sv
G4JuKYNvlb2PVCv0+ueJFO0Lf6GRkIsKObClE7SwXra0X66RazYWicQ9Qu9BSmba
TQmtN5fupd7IrZSuSp2zsz7mmFHXocpXEN9MbKelRWVmHDZWESM9Zroa5xK+Yt37
+tMfs7RVwdLKJogN98rINYN6rZpV646zum+EHL1uxDeihQWQSGmRcRuBsCyaXOJy
a80TGbMQn0WXRILmbvZ6UVL9IET+/139v0n/qBQINVGqvMf0K1N1wEY/6Ixx4Aca
44+uMvByNWGmLYcn4+w7d1Un1S17vnSYDzyX9CUVVf+vh/EUjJuy4QVzg0ZC6gtZ
lp8nyScBzVQzNwP0FzXqK68m2/gc5Kx6AuMT8FZtdtpSKXf6ACOdQVDshr1krfPs
6uLaf/4AzhKvngGSBAQIF+A6a8q+tJYtj3sKOKlerm+8/k7E8B4doa++fnGfDK67
H0tEG9vilIIBI5jOpg+j4pWLx7Lrcny+keJChDiySbEv8oOp8FeiHxsO5g8x8mwm
S4ZyBYX1XwfNPg7I8fEzr2sRnk7TnZ0cf0q/a2xRzsArPLJV3zC3saNrrKztOxFI
MNFRtWQcId5my9MO5slcjVFB4kBA6V9Q1IyvAwcwVe0meXqIG5tdhQR2qyK+wjUR
8rVQbvQBtY9tDio4s9E5zHOTs/XhwhK0CGNNwb47qPu7JxJrQunHMcQUm2xS0Ugn
WtrnC5+krQ1bJbDLq96uWYznFbkf/2CdMmPtmjsZu5RQt4d9CB9q8GOuu2IlqUKW
hIKm3vVtQYsmDLrUftnFqnMmpuyYw692nKu0WHlNAN0+Kb3NVHdN6B74YlFUUVM6
Dq0r1gzaNdPcGmZapUibPuOFdhVsegR+uCffQOicYtWSMXJcOkSg7XBpfNqs/lny
ltPWVwhz45AUPj/eMez61FJmVRflV9cFGD5f+v0X4tSau6WvULKx5V+y5gQCm1uD
4kXBTE0JoHxch5qh2w/3cccmAOKjE5XsS51NgFRmHCOEaSgupN8Ked+83ICMOHgX
6PXwViDt6WxYpILEeht89d8xIFbiKmKMByYyCvF993YzuANE+87bP6UVwf3iWlr1
E7vWxsQxZuZ6zwIESedY26Yi+DuJ381sZC4sSrnOZcWgbGOYIlJ532FUZwdcXCm/
/Ui6Vuq2GGD4ZjHpz1h8fdGGlkec65bTp4WhvIXYed5WkK3b4hR7UyjshsVTUKdS
xer0ybRNySf8OzYBLMLQIS+Wo6PjN5VmnBAyGXNPOQcu88GNpT8peF6UDhnXkTYp
rAjFl8hKAiDcAtLHGfkvj7JrGG6ub8u0zURT5VoHaqRIZZWByOtd9RmwnidKDiVi
Ab0CiHhsfLQX3ePI4DodtT48vtkL56FXS1cLcDVpB2dNX9CHD6GaxKJnkPocSlPO
057cdrMRYu/HekQOM/exOYBOhtErbW+DeRIkSSNNvuaoQzoQaPOQS5tOKjJS4lzr
WOGcyyUZGZGis5BHXCC5RvyfuoxNnTcCkdUWUXOrZygADMqYGlwxS5EPKoS9cWfE
L7oeEpvEKQ/XulqhudVGndWtujgjf0VYtWR5XHkOMtCaREDl3Qk4RiJfh9vjNqbP
R5QuLOPCyisqmR9AMWKroUoIkE56690vBaYZZYafGzJf2B7BvPLmqkpe7f98JWNt
V0UbiCk7XvwFS5acytiMLpwHaQwzWcP3aYU+HN9ew7qkBc+bCJsRdldut/X45Rtk
SKFGpB+nJeJSZe9MA4G1FJ1UyBXYRP98nXLQxmR2qH3D2unIRP21+gcQWNzErp3M
iWokA4h5f5RK2nQbZIHhPpjrhj/wJqfE4OWkNGtmnaE7AYXz2Gf9YBzFgyTDWb88
hfh3GfXa1fDFvVQfOxw1WiMopgJnJWom8PbofmjGbdOMqJ20nusxYzewj+dt/YaB
YVNmXRePPRSM+aiDUlc9nqdt1nawdtmv+VRP5W0T481h04neLtu0wuZSO0AzBpc6
yNVZ9P1IIFPLMxVzBcLlJ5/LFzsaFUb3xXJFD51qES96OiSRMQldMx6Ql1ZTF2Hp
8HsHPg7JWDqF09Xrptdg1/SqRf+AETN+LAiFp1x8DJCzEpYagdYjGLpaF/cEBjQh
BAMQ8bL/jhTtDi/EKz1Zpm8NU9zvKG7kG0DoFpf4AjAwLV2t4gAl/kc+pmIPyVJ/
QnhQiRHBDWtgjjUk58DI8E6NJfvbh4cfIZ8EdQDtqQFmPh1Wbpz0mTiVgFSFAY4w
Q099qqWCHk3gsrtZ8UHn3E4Z3WX84jLZDjGJ+t3okhB3ftJm9oMmU9JClKUtXoLC
uBoELLVR2aKQylcZA6JUM9/usQz6UL4/Yl0EZO2Qqf4B7WKSjs0SFQAM9U2AeiJ9
GQ4StVAWnDdgeCOnwlhfaS+BAUN34dLoQ0xv0C9KRHvlkL3iRyGr73ofvD5gORkV
WluYB2Bs95gLKu4nDUgfS94xpcG/LKMJBzGsZ5knErc0Y544CwFxjXrR8W5ifU1Y
w4ogupRrTN3qXdzZRb+XJYDsJvpjaw9nT27yx2Pbkb4vpb2fMH1mbxH5WdHADwRs
HV3kSsGVi7i6FIf5JETvxiSKWmbv89+p2+1GeRd0QxIW3pShayPOqeu6vGxAdmws
k5MoM+Ktk9ooEuVs5/u2QLTVSkhw9LyRYxIqm0S0W1yBPHWz9sQbOWYlI1J4aDSk
xy9BaUPGx9YsYWYJ8ddVpwwqyQ5UbxTrKIi42YTk8M7yoD2joiFNkqRICW05hrUr
ldRk+Q7hpkQq2NkMo5Gjc+dgnQpcY8MeGWld1aHQMcNqPhSq2jicPGO6FkMPB4WG
fza15AzaL/TPORn/TH4VOOhabJBwJodfbE7sYNkmiCEV9KirEcPfH9m6gc2yO6GV
LAoyvHq+S578IYIRWEf0iJhjJk3GqDPQrOAqPLxi2YT1VWysMJIkQOK1JayP7FkP
Dxfp+cdXnbnmXJeqAt0qty7K58XffwLCtYEBdhwDNSkwOTeEdMtkE0QbuAVgvyqO
tPszDfmf5pAd8pNafCmdx/TEAfpu3rpj9AGHSeobQdqv9cDalGAOM8oTPlApgAVS
Eyezt8QLsPB8RMtzDTMc/o2E7EJOrvRGigCSDTPiWe0Ey1xLOu1K3xDvg7qg9bye
we28NIoBnrc+VJf8uYupGde0N5Tm39dg0ObtzmrjHK3B4X+HL5SPrmxt4gz0GNoN
vJGQlmttBn4zIoMe8ydVswMELpUQXD/cihzDc/g2lJ4XoTCsTrBvHwO2H+xLfPQy
e+8s7g6Xrp4TqI4RCzhDVgCoYBDfSwgaZVu6UhOwwMYtGhRCJuCftAtb4PoqhoZY
1URNgP+I/egnKl7GgAmGmD6+uXssv6RIo4VCz8uzUKIwHcB76xgqnlPw0x8b9Sni
YIXQ1jWMWzvlUlzVlaxnL5fKARkj32Z1hbk0uRMTCZvhx1jB6pmBzcqa6o1Wq1pG
+WwGwg2m8a+dlI0OOeCWaNTFyb4wuJCjvV0J94BCsa//vOFFWKtiVuDRsGB04MUZ
cDVp+dpq93c2ls4k+dW1sFiRHtc1F2Su7HA8Q1piW/QPUyyTM2C1e9yzFHJ3xPF0
G1xTJm+dmJPwvL2Tq8mBzvWAECXaqlvzdMy5fTZ4xabXvfho5fT6hPAMRm6Nd76l
jHy3cyIbMsrLwc8ZGDPhhYU6eP7wTZ2CId1ccxnM4XwPOQs5BJ++K63uhmjTx+b4
LSZSFJTZYaMX7TfO22YDg6V5izFRdFNv6PU+E2TcZ+W2gQOnMkx5B03wrIMd3d74
UZvo7ub6Dc0Kty59DERIXFE45Adm4v6aakKruBvCLID/tlRUEQNIopPVstxd+VHQ
okfbqGNd2r18tj2/DHYAjGUxiNgIC+5eTbhYVAj747YzQKXirAnE2GbOpJenCUUr
NmsdkjdA1E/xitO5P+CCEkTPezUzr26+6kcFoDMLGU+mTop/YmYKWBGAYIC6k4nR
8kYY6ZQbW7xhfdt3BZ0eQ9WCVMn804gkszjv83fCMjNN5QU1HIzkI+fSggfHxPdh
JUewPAD/KqNaljeEzLmDUQNNbxcClw8BRV1cSRCgTdDZVZ9fj95Uk7UZ9zitBsh1
199pbtLvC4ATqsKo5x+5uwoghqFwOPip9YKsywX5pdUXtRNZPIKGQ+3+8Kl4gf0L
gFBCE5gkcMzxhxsotMvMepsO6xwqKSycj5zBdBfrNoxk50jSXmmLtTmiFC26ZdPG
NQXn6sqhJBNA8/F7LatONXUTiCuxs3ECsSU1hN3K9nzVcFwgovKfO0Dm8KkHyKOs
PG5Z3XbawGg7a/Oeb43WQmGsCa5qw8oaWJoy7fp6zkf9Ofszi9gzru9ttbHo787P
S9K+CG3Uut+P73zKjdTqRjOLLTPpwpV//Gn6NURyhnq1tvOG3csrfdFLG+/jPmR5
ThdO0Z8Ggem12keV/IcIYhf+Qe+A13WWGn3V9aQRkG/z3Jxne6XWEN9fcLUnNN2n
Cxfr7wkl92QrJgH/kGi7OJk97CHQNah5HW17RITGa5xExlydWtFuF2saWg87daxi
PP6OPjAEx4V/wincKb/U5Grec4Nrq1iNxsD5by24Os1FFcHrGlqcJ/qp4bpuAtiQ
e3k+lU0yBontXhy7awaaYGUpB8gX850XKY6QZRJbu76PV2wsCIHWc3XoayFtnyHy
HvlMSJBU4D4o0MpzWNMjf/uEdSq2GYNMsTVzA9hLsUohypDnhq9sOHn6WocJw9wI
PdJJDP0eujRrH2sSsT3LN0du1wX1Hs5ORTO2q3tZEFml4lLkmaSDXt+7WbH9U8Nu
dsUTrkQxilhtFK8NQzsISTUh7qyerDd8JZSs9iIGp+Pd14YVfL0tai+a+uY2UOHY
c/Yg0sNoSa2hGRkrTrNTzYqwpNv0TJxzsnGBHCCVX2X1LVAPzBpSdE+84pxQScMx
YJcUZHzzoDaPnPbys5yB+BTevLy/KNi1kh5sO3iKyu+8J89NlZYsFizAJgw/Nc9N
LPGABqqTsgTFOH7n8swsLg4x++4Tnibh/P8YUXZK7/N9cLSatDMKlt4BSia86AP7
TiQ+baJOU4lc1TtP7yCMl0H8411QAgUgH5Ac4FpdAdzqokBYYInNaoWWLCSSYroW
7BBLa/ttQFvOwCVjGB4yBxFw3RTJjnwxg4nj3er5qBXYAKkyJtrR6S4W33h+Mj/e
4k02gQvKa+r43pGbZ81Hjwm45cJCYwYtgEAP9UnL4R5V4gdMownc1k0A6S8LQMac
KljSA2v0XwqTL8oOgbfgTX78CTF4inWjFuJjsTFp4bHl7VUXXMcHZyAL33PxhVmC
VkqHmtQhkRe4/8QuetIVajas0zMsuhH4IRyz7XNtPdhlYlhcu0i82WqRpdS7fvEy
e0LXlvC/oHxDlKAC+S9++n+KOAYyj/3TcouZvNQOPFGc9OYZOi1YODGjfbYULUhP
dKEBaL35QVoaa19I907IQuSsFhOyDqBPu7OnfTvWSsgXqUl0CxKfjhmGo+pyaHkV
nhkRAcLv2bGhKLg7LKNzn4Cqym33+oUnDFBEtHOfTb3YSxwX0duqprOmroPI8pKh
Jc3bYAkbC0oVmdFF2pXNRku0Ael8lmc30yS25PaCntMbOodjaejDCQwgU92dL9en
2pfSIw656eT4bjjJpBsg5tdiIHD6OGstqMxhF8/TYEhn8fTzfZXDmPlPctcvr+/t
hv6GsqxKsqsJW0LFuz9ExpyD1NKNvvM0PjLM9NErSv0ERRpG4azqOJE9NO3HcE/X
O1iBiiXJBDZS1XUTiVR29RVKd7NbHq6Eh39FWmzmLz5ZncPeTbQrY0jTgSrdIxyd
3hPKdQbthdkjJ24uDjz9NtrWo8mScsS2nAXXHNNMcE+e2EX9LkUh/uBhlYOeOmWO
YMDeQ+j+x98+PTUTGoRZ4QHPgepRAuLTN+fxfruP2YAUyMX9MiX0D5/X51O/zjdM
KGfVcZNBnbto7HNksKkuNcZG0sK9KaE4BQY4/BEu89cKBwpxf3AJk3ULn2CYm1an
yzVsQaMtmi7jmqRHW75JmjjtoMsNXzx96BN3tSVD+1sdOH/hbSA9kwXLXUAODitD
KrGaNBm4jtD2afK2h96n5GogD4E/8NAHGHctHb/RmKh1Sra7cenIv/K6XSIpzvtq
1bhdRXcKiZcvzIMscGof5eaq1zczo1ae3OtMR1xbrXKjNh2ZxmFUQn3ypHzdES4i
fGwtjAZdD6rq05rcDed7A59r/PlKi71yal4lj/LtQZS6CRG9fh92ySYTAO5zh1oX
cperTwdTLZ5lH3yNsiFxDMQNugGXHVpiWWMpgnz4I2T+ZrTEHvI1cv4yeKJuqc9O
33eWTZCC6Bk9jTfgq7lCm1JtVgdajXt27YDsthHRTc49UrTFNSiHQf4kEHNvL2za
UCVfy4WAtE8FjLTCIIbpqo9R12EmgKDEfhjm1AcBwjTtEp2zcslS5dFPvX3ASUYp
4DUczj3M6loM9U3UgnMSnGptJsqI8XRuGlZEASJ7RGOrBDcIRNnUepKk4JtoOHLg
vyXmPfxxhwmXv8VDVRPliDV6G3g+Bxvx4AwbBczweDue4gdu4H78RXcQH6JADS52
0paRgKP0OZAVyX5wQh/gU0+z3cTbanYxmAm8H4tWDeJzEoo4hP3Jhbp6E6hx6kbN
FVMB+eu3gmDAAN3fRillypSNIs3eUvZYarvpFBwtFiJzTJzwmgYVWuww4UFKWjQr
74Lcgm14jn7mo9N0ISx2jTURWhCgHN8kRcb0bwH6LoVcLD+4OHCG98Cdb2fBAhG5
jDuyhZx7k9alYrUfIz8KDfowlYQCijpkVgrwT+pgtwbcjI5BYDh342DOgD8ROjm8
//xHp5qA4sXXoXSrsZX1A6pG86+cQ39+g6hSG8n7sjXS0O6Xiq0OJB/SYGp112A2
lZozmEBsfI8I/lhdwyR+nD9q7rVNQ2LV52S3NGzAZyfaTo+a5E5WRPI35Cyh8Jgf
eHtWOQFlnDCe/WQaV1vB1vU0G/XhCMFJc2RR78AOIeYyfVrHFDwM/qjRD6E/TfBW
vDNq0+fdJE3EUPkp/hr5cb0l688G89kQm2lXkdkNHmgQmeDJpTfeQU+co14e1AlK
N9/D+AHe0NLaFFk0HJZgdnmK5Q/wG+g9VCltJiuInz/3PjNl2/4boVyEd2fXCDul
HEsb1CCA8ON1fZzuxqTHBn4BRJJoj75egUzAxNEVxl3FpV5u9sYZ2dd4xBogqK65
6brBeArShfY8x74S9jAZha9gwkBtRRugaET0bBv+FnieXI5h/Mrtxg6Wf3nhZ7Q8
D9CQkCUHns3e3jnjXH3wyBmNvwhSLpnodOXwaSRyZ3dpwHd8SQeG2PxlM/5cS88U
LoX4vXkATHSXcc5sRLFkEp4cWthu2exEUoj+eVg4HOY1ndykSSlfIVeSjBjlr6or
ksww0xInbevEY9GbMTdCCl3DQ4Bm0TzU/K2+FORLq7hItEKKFOluKdqnb0OImABJ
xn8ZMm6Sv3++H8t5EaaP0ZN+xr+ZaTFvGv8XSKZ9fgBOcYGTsA2+RJfLYARTyoT5
H9cKVdkhsoLaO+NF+pyR2eUYVX3+QxMZUkA3Ka7yVAw06uXtagt9rjTKjlsu0XMw
HH9Ef0putRt8jdw8JBACKyZMLTLT+FHMLaNsYbmDz+uI8gXQClc5QNNsxMOGf/OB
7vpnY5r7a6jP1kH5eYNwkFKfEViMEMYTSy6rLAwFMfOrufomxV/l4lskhvUgI/NM
M6X5C8nHBqUaew075m6U+V6k4SbiIALNP8Zo+/vMJkVgpPknyr6yVo7+PCOJZvF5
GHExduVInrX7FkZT7QIj82XlSCuFzxbPc9An+brgVv5hL7vW73vhnUUV12wLr1jQ
g1bCIB+bLoBHocB6GNL03cZqTn7Zbb4QuVq60iN0oXpaoS8MNUKxeuZae2SXG5yI
p67eOaL5o8WEFQ7DZMzf5/kWPNXSRyVEYbF1LpXV6Fqv3rgPrlALRYp9LQfJljVI
BQnA6RAa1ho1SEUbltZdx5o8qyDEp0R8csTrJ1Y2Hc9BukdQjJYcZQ6Q4eg0QkpG
jNM/pUMqa6s3yK1NJuujfIuYrU2zANQ+wLcijd3Ap37FP5j4fY7j9cVVPQ3HViPu
KIjpUA0nsiKrY3ie9WXxOFOYwyHwisDbZR49KkigkCajQdcYTjkbJjv1kzhn1z35
rVPXEaqPMPX8UesLCfRgaTk/5YaCQHS3E7VyPR6TrjpFhRJmxXHBkyEBOKeb81XH
ggfpiXAhi7SSUBsejEWxe1UsNWkc63IuaayY6DTjPxZxUAmmBMp4GFoSkmpAjsRW
UjCeh2YxIfkYMP3zPGLvshmn3zDD5B5dyMFJut7wSgYDvIq1VL6Pd/A11i1rtmcG
Zstq/luXVtoVF0uSbu2ppSVbR5552WOM1CcmtXn7wOluOyvvAeYAvIx3xtM6T7Jv
h2Ue3MeOup92MuiAJiZCanps9cfEcR94bNmkXmSzpXZIrxBy/Bl5w8z8UxhQL1dy
lfXGotdMX9Iz4E9jVsozTrxqOqXYBDmqDPmEakZMQL23H7lv10L5MXRsGc/RWbVw
r+OqKZJWRB2YVy7Ff21fYptMADjtbBz93DYXkgUtFeOzv8Kf2DS8jSS3Lp1IXTLO
uQ6QPHQv+9tNMgI8HkZvQ6+5cAbCudJAs72FCMlYb3vhCNFqfCsMe3cI+AXbBfGY
mle85MN2aXAmG2iPYBBFNNef7Oss9osjwBtN19L+7AhOqjJ0b9viAnBOMzCqLaxa
IkLLxv6zSHTpKzPb2rKK0D6CddFv/318+voHiAJrOvf2TQLTJbfxgn6z18kjXQFD
Zbbggbr6zrmb5P6Lq69imiARBl3zyP24zj/jZ/ugSj0kIwTC9wlT88UGHwabT45b
6uhSpe7B4b6gtiGH3oozGTbnmIDVp3jYpgOCfxjQkbFs0RdNtbZMhNHZA2ZzxbjC
gw7PpbADYo6KApw6ygNsNCmKVafYpI4Z0618LeVg4mljPjHGKr+ySphimT8KlFdD
XxAmmxaYdk1Hv/r6EB0rRSMGTv4jksZZGQwOWIJkOLg8DfuiE1Dgae1JVasZBbMG
K1loYwy2F395N+krE7sfDzc/HNVRobokOtHGQha/m0YEuAWlZFShUikXLIxhK4uw
INHdO7hbxV/0xyXMs3lhZIsvZBZ69AgMapTnIy8YmLM0+JS9sY/UL9RM7OXL1XLl
ETNV1kmwhIwOICm8Vmy12sw1a5kbsuSD9A5ooylTvTtVS7bk7HFSiBfHVi+Qgq1q
9TWxlCGl/Qj128JbftzcbqYR1YJK7UuhVp6T0DZw7390fdC4Jdezgcs5MMaBEHnt
DkMllTiD1fapRtQwLMShGWWcciXlT5n8CGIb6bcd3XGzViJKgp1PSnIUutGmotR5
T4B7kNwm7hLnHNamDMcPbwojVZyiNoPWjIYEQbngVFnBPmThlzg6HO73oxATEZ34
534ymrckMr9H5hIetaeRvl1UBAUM9sEauqaZdrMCL/tRYQaqQYjz1QtQ5jAF4tsJ
rpoFNOr0712bw1V8c/biZBUN3U+6ZzYYFqz0LimCYWpWOEekzFovui7qW4vwUed7
RFbCL330/aDZm41l9ZevOamgwKxKwE7/ZPRI194EueJ5b2iF+xiMEPDAUtAvm0dy
VS+He5YfuFJGReDPSl8bitZanrq5YOq83bnoSA0VEhbvZtoZSEjdwnXy1NY5NKmA
HSs2u67eL+DBu1arATuJ2sx5sTyFnFrlx5gE/eqAoD3c53imBVbFMGI9A5qpWE+n
usm5roEARFfZKrdyesjXzL7eUA2MAg+E9O2dbwf/kBZ/EpmTgXlcr5m1g47InA71
hwOCFM0L17VH4YW/WUOB26whA26OrY80sBawb4c0h4kHGWq5ifSnrwKSpodY/LOF
HgbFvwhM39gFYHUohuIGtaZRJGi1yd8+PyongPL8RpG4xN4P3MFFdt99+GU1b/0y
JKVrffrEshx/g+Oz8R0zs5mhWX5BNCeAAcLWSPkzuOoNOCC4EivMu7PbMS8de7T+
w9zsAnFi/Gu+/GqI4f3iQTA8KRKkQ/uAtmrHHD18xEdIpn3sllnWq5VHn4emER6d
TXyKf1SfYvwrT84uXdefJGGX1qhOXipU/ZNRhPaNCDrV+NnV7JGX0F84K+P+6Qq0
k2qEFgt7Jbdd03dbXlgISdl+1c8s9jpQd+fj51H1T6An7nIC1P9+Cgh7koEGnxcy
YVNe8YXmy39JXGlcvVh9ntWnLCSp+N+RkepNgif2samCw1B1VUCkFJnhhF8A/IL9
f9x8JKascSTeVEnBdy/hxaECiJdBD8gIsyt85c+xoLmOoNEmStkKziAyL0BIQZ9L
++yE8A7oBDcVp+KMUrsFgW0nhy896LothbACjx91Ovno5Ys3af8DgCwNg43Or2zZ
l/uWOEISAvwNNLXxBJD0BXuxuNdyxOe434EWStzA3RoDo9m/VwI5VzSB8+CDXN7T
PIdfBc+F8e3cFkm8nxQvwN/j4F4ocNSNTj+YjHtcuwkvlZUkD46Gi1s8sc7whQGp
31vFud+uR5kLelcYowI0QVLqtuBN2wOWelcUhdJj172Lc7HF7DGry0tA+d1gnraP
JqqGyB9lcCqTSj4WFGnFpYbkwrXbDzHYCVYSkPrcN4LcWcwyiRdPERJEY3zaEIUE
GxGoeUi8uVd4A0o883k7+UqUS6ZS/JhlojgEtJsYKumZfgsJDsiEg7ZAaSCS7Ob4
xPDjpiqkYYFSgPXy+JqsREQRT1HQEbqJfhfyd0nmXNBFEfFjP9Psv9cfPNNbGEnd
6TRgC0+3y8mkEdEQ0XL1cV3NKgwJzvGOE0Pmqn7VhPPQxpFgd74CphFLQpiC4WZl
SJqXhJWrBfq23BlJg+yR5F+Qe23A90nl+QTcWrNP4pSgwskOzFHG0SHXhNIdUAZt
mO5HohftvANO1T2PeVtmiFVSizU71cP7JIwCBiTqYzXWvFbNENhQ9Kde7LaXhP3Q
giF9IVqkdR+KTOrtCeX+vUdQdlbfkDXpMPCK13XY7Z8Q1ecmwnXytfr+CtIqhEEM
DsTMipPCktuyTjHBMqTL90I2/P1w1fJruJnOuE57izzNSul74LXhWxbTgx+fsBpx
BplDz2ka7VgCk1q/X5BUGtIixCZzMrK6sV6peCvJXLEZ/KqWBjaY4np+qEPlcNuV
XsKs4jLzAvm0cMO2h30HXDiHNyQZKOVdP2GeVMZeXRMYoi9JwSTj9BlO5jVoxfQJ
jIxzvdCyfibpzJr45+nGPqdLPkFf/K9PP9vy0ENPf+pKa/EfMDagB8fy/Of6r9XO
L5GR730HHm9CzLZSTW1OCDZ/ph9mMwCeDNohw7moVc4SZBE9g5jPlgI5qSaXCHMw
jDyuL7/UwlQPENCCOEj4YT0GlHI5eL3JyfMyUhq+wO95wCm7eQhPhWJyW7/sj7Zl
MSSilpUfNAUbyGOf72xSu9+oR47KpdlrqiB5wxMDwwAu2kL9Pf/IgESClsMSz/QO
+r0fC61Q67OPnzDEBT7LrHAhrOxLgGJ2K+hh+kjkoIeIyyobR2BpJ9Pb+ip1g17e
tPrQgnK9t+ILfIcnr8wRRxcFj3XdUhOcZw/D0ZKWHLtFyZ4ST6oVjbd8leQiwi9u
J72enp9zYuFLECAQjK6MeMNAW5LwHkvEVWKPRS2jzJ/11d1J1zggO0LL9MXroKzo
4FKC5v3TeJ26TzGJc8WTd84VIb1IimfciKFbSKNqEH0FQYu2Q074hpneCRryOMaz
1FG9Uon9AsXjGjmEXnUtd0lEETJcCZlpEUN8lcfzboY1Equ1NnDfFKQJvZFwhEXB
yntCqjw/osDsol+OYaS36tzWHNrpR9MrEUVpHU3y9SXHCzHdNjHentlYiS/h7Z52
xxe0rzyC1OWKmEfqVt3jkevNrveiTmN9aum/qMyG5xUEbvDORN4QLwXM25dGE1lP
7EiKGVSafK2sooBf6IxpgQR9ErGmmeZo3FIwmENVPpyOzjpIEbRpGVZvlrK3eVV5
dze4L8E1OQ6/WKOAww8RBsqCxmMSrAzZ40vT7zCMHNCp6U8c+ecn9izkO/2e/Y9b
g8SXXsKkVcQYPsgdyW+9XhfITIgJlLo9sMbf1A4NvAwWxyKS6dP+ICgJ51I1z/rl
yzJrDLpAhANbjR0NT06M9sVCr2EDCV16ViZ1qznp+0STuIkC1NFHOGIWPxTdNKAK
BnUKVz1htHFTgBVQk5iJ5IMWoAHzcz3DBYchWgTHFjQ4rKPHteA9koFz0tIwxWr2
dSHHRsL6EIboae1DVL0hXoFDt2n063LpjnmkhT3YrAxUw9WjNNdfKjfU4UlWz6SB
TKOd8ZeaD1X1lNsGyEvZ4s9CF/CdYtl9biJURRT5uOhIF0PSusiIc5BUXiOevKq+
QRkTf/YUqySY1pim8fYsVXLy6Mmz5MM0pxeAthdgUBG543632Ee+h0lsLbw53pyl
rkXuxYTQwOyt5amKfxMoTzLve6Gx/sbMyyru8xAv3X0tnvylU5j9ypKUzNFFPabB
V2Lk3PHCLN6kjyADpd9o2OLZsxTFLxTHdccYv7lRTYa8zwlq4U2w3mmKJujz1qdD
OYsx/rgoZS+faO1Zn3pUB6TTFmjRNV9I+BfVZD0CJaxcZxd8LIXf9N53zqyp3OrH
XXKVWdH3K2UALO7rRa6T+KORvnnSAKYel8/lBCLNYaroZxS/Gl4BO9KSErITWPXh
BDe5A/kfNeBaKSB6Bz50UbS3YUszF+VhU9ieRZpd8+QmH7eL/9WDxFAJxkx0Uqzf
ixuCcaIPdPsR9JDu3OxzhcV180bV6aNpHNmbWNViUnmmgAhlbrb71wyTDx/hF6n7
MAnZuivNsvP9IgbcxWxUAS6s09q9sSRZ0PDooUjpvzxe/Nk7H70+ZrQr6lyE//0n
oQ2rHMxmHknUCynQ/FeUSKnWUqIgo/De/yZhDDPeOGUcdk5M437OMKRkLpGr6a14
bt5mqDGPWPDCOsDGWxUiL4vUWUhrr25vTNfUHzeJ618wa0XoZpu1nxBRKVuZFL/7
Xi9fAb+/1GAtz9G4kMG6vmSfmPNCpUTwsBJ9dMVcqBQyMEG7nTkWB3FkwTz7j8tD
Qxx6yRiooTQQbdWTQN13Jz0o4MtMmlBb6E6AwPchYjsiapcgrFmSQ5duEas6PDx3
uTahvqQVkqcnXmeAQ29BKu8N+2mce325JvnZ8yhNsZx25o38rqqNxaZsonc52zxn
C7KX4qULz4SEzkyCqlRZc5lFswFKgOr5fvXjioiry8pBOMwBum7NelmBVPVOs+4w
2tfnA05Zei4oX2Lpfs6o9NC/DMQsIJ9SSLzNfhUMeTzlN6JHm1h6ATbRIfnrzQIk
iUfnI99wDvNVpwyVybtuFWqjjzvZoLNy8Oy2EcwmhBFHeH4OcoAbM5BHpbBzZXwe
yjQW6SRfnMIIuoCvLYQLgxbzn4+Ko1bS/lIOT9gQ7prI40H5XSCsfyaslmR+Qo8h
ufvjYgGMShaGwdPLv1cSYOlWNxupD24qhpUG1Q6/iiVjiMeU/p50wBSc5XeMe/4z
Oz64UGhrCldfl44ZCJljKAs7QkeJ/FQI0yy8nzoU9Vur46tZJrVoy5cNXZpjNfY0
eTHgsHNlQMxOX8u3PzQ3UXJ0xZazYwGwT2/ICJ7ID13NaL13NlNw0ePNehiAmJlM
csSoQkqZMUQc661lh1wukxL6FYkhJaXq+8za1ndbstoyGaGxZf1QbXiBNinoDmCU
B6p2SG1KuxkgMVGJmkPrvHwRfRa110TgQ4q/f7KihfvWM8cLPFhWMoEhNVdISYDe
O0sH5IjnmA19D7nb2QGf/rL/1s1llx9c5QTH6Yb+NpWocRNc8Tl46fQUzAcYoTwc
+AOsKbXQR2e16E/yxhZleQEF8nr8ZdeFoxH4pVUKruXbimKGFa0gJiDzwalzV9cF
N1F2dAF1EdE2gw50pZYypRtQu8buzYCWonb8VgmEutuDFFUXzYSQKbirrjWPPNHV
lrHS6NJKn//0klXvJHSYELzN9aGNH+mlxdc0MgT/SFxmQJ03Rrz3XcWdJNEsVev2
ZPqCQdZuCJbqgtNmpJiDzYUv1Rr9+hZeEq7wZHOHonNaEaYTNX+tYua1Q6B1IyVX
henDw0HSIz8q7FzbA2KLmjiREqhGmF8FaFQxg0GP9D71A3SmSx20sIpzMQhyCRIM
HGzDef321mGgcJsQpwE6yYHH4xcvMu8GJIHvzbFFlathaEo0vTGcebPVL3iY+9m5
14S8aQSTGTLs+UktF8dYQ3Vkn/Ez1Y8VSpOQR94n7V4CBeFypQVSGvrGfl0u8GOO
Kkmhq8xcSJyOSUOE2PzAZMfpqvwKSBrb36o77xgAmqAoq3vNPR/UtEL1wgfglHic
GSVTsDltLSCYa0KKWt/9SF9iXeZ5Y1OgN/eqp2rkAB4wjJpGPxDHFsG3OGBQCVLn
CmZP+rRNp0UGOO13/i8/mBxpGzvafXGiA2f/XjUg4GjOJcZ96+03D4MEv0e0Hczj
94kmS7vkEwngD2uu/yrlpYgcItgV+ry1LNVHj2w2RJbL6cQtDQkxMnaoUOz+KI8Z
2RPfyHK9W/srGiv7+E5rY+ySLGg6NpDqiVKy5WFZOFU2cV+6GZZiGWO+rlU2UwTQ
02je1DZMButxzfI1iU7fYcpq7Z8SZ/utB3Z/ae684stXj6VtsRIUUAQ4HF/IGECj
qFU5o2cPlc2RjKHYL5tWhDRRFKT2NMAY0w8cN5dBGlk9OaNhcJBZzz3s3q1GnriZ
DXycUgs5lWXfOoxfY3Fu+rR/0bGHJMGEW1Jdgz7OoQSS1GX9V9Gitt0Zdn41iv9P
s8n04x84uloSNFWnm+qn9Z1hXKYuS/5dSYxOe4oz2mO1gVdyCkN0km1c5v1ZX7iD
qqcK3UswL1lkfGjQSpoSmIwocc70OoLZqY6obtxznTMEcrsnNVqbdWeMtpL1ekxb
8PWAH3aYVa9oWRdZJRpx9UT2MD2Twmz2Q7fI6N6fe4ceXoSvB9VbARa8Wg/mShvz
JA09bhwz0S3Yhi27EmaSduR+nKfnesEEOAvSWMnfT67+s0ERjdzbfwhjfMe1KzbS
is9rAl94Vm0OjE5cyXIGEjS6lJU3IjGQbrTkOi9iiZJoCIHfxfqc1zMQmZGq7CcM
czpDeLbFwMEb3Lk31RQuFBKcBhKecgg0yf1Ui/oxp2baoChyBr5tjdKYslFzoqjH
Cj3zK4U+Id09dBAJ0mlYDWTbJRGkGpF4xvnXfF1JQZF+D3xMrv/MhfhRJ+VTGYUs
0VkYwedIcde+g6uu5WhRHm9B/6GLOIIgeM7R8cgL3biPV7DEoBXW057Eb4RgSJWy
y1v+2F0GWtUhCOH57lRWZf5ag8bDkaf7w6JLPMBxd/L/p46B8XDzK/1V8L1CgVe5
NM7bsq0WQA4DIIA2mWFdG/WOtyBC9lNv9cdkJUpRR4423X5QYOLTHp+Cl9Zcve7D
2p/y+Tv4+3kL1PDY2LR68HGkAqNr2Y/osLB/Q3MyyWCp6o7HasWuzbluDqbOpaHc
x78LkqC+Gyk6G8pFAStSkNFpUUC3g8ncYksDbmcS37mmlcFNDaUyw/A6d0uunf4U
MdVqlqf9L+4rGV2CdkmyxpbBcywbTVlDsIFG7WOuoDv3OcPlOJKks3s4EUopPy+T
HJRJuJylgaWL9KDHBTuGxAG5P1Kh5vppt33fM2uzj1ecU+P9lHmk7avATk42Z03l
ZRq7ab4UCdnQ4gFTE+T8FRo7ouKW5czNIxUcNPXm3WwuNRv1KmJNgVjgnjUoCkB1
/olt9CgyweziWlmGupimfs4T1kzlGMiHb1l7/KhUkOQrX4tTTz+4zHTAaUqMkTMX
mf+e7+fyaN/GuvPt3Py9SKpPgCMQUTYuDy5MDWEdneML0kCfhoIyMUmg3umF67WZ
8P6liWdm8iWd+Kmt6m26J4shtda7Rx/DsutdxaK0ftIII/lLoq3xHAccp+ZloT1V
1LJydZYMmVjFxcYINgA5MG2gA5OAXoR7tjrDSk4lduzbSxadHyUaHwrGe3bA1mnZ
VWgRMWpFmNyaXG09r38EAhmdPdKVb4X0MQxkTt5OUuw1usJ0jQw2kvlKzINO8cfw
eVLCi2eXkU5leEyihVmsBupb4vb6v8zCSs6qs+6Mrjw+UZisK9CKmRC77Ppm+UMX
vys80ItJg8HpxWUx3djmI0lt5qvDgBfySMoB0UIVn3eY3w49RRpNm1TyinjOKw2q
RgzjHFlaFeuMxEk2LJ9Tve5KSzYKfXlmGoNn/NNAi+D6IkMOxPWkG6CNgjhkkDwL
+gNHxDPNafTT/tkvCr/BCqA+Amda1CrqPdx1Z9YzId8yPABqaD1zWFG6sWdjloAw
sv2W3hBCB845Sfwvah02f4eR7eO98I92u2Zs469W1Bw1I+TZ6jpdF2HNSEf1FnQx
w0ElhPxu4Vq36B1ojVnQziLYerTqMR9fUnMLpLI1J7cqCFclcShp0IY/RmhLh+Bp
VLvw8lJmN9JG6O/2bHHYDtHjqauAkyiaKVK/L9DxUqirkEPl9CWBFbh3uXIHnHwD
Az2yE2kzLcAlxzO3Qx058WskLcbrmA/nmxWFmPepnDi70PJdXtjCArwjHH1km9Nj
7m2jNT3LyD7/p0bqjrIdLl4v4w0nSJ0YYPVZ0CQW2CQ9+0cWfpMQ/UKliNzJpU87
Qory8gWXwaiQO5BKtEzZXv95/3RyDXBM6ukaJv8PntFNQCUxQEACjwKS/tviYJYW
HvRKCLYzoRY4j6tapiJNiez5doPtBPFotHSu3urnM2O2cPebFb7zZ3vqJty8wptu
juULtWZfSPkAEBVsvbp2eRbtuIRxWkpo38xQlc7myBSpZykyoQH3/UwV3VCnL5h0
FexyhFguu15Cbu62+M89oyzsy8ymPnxTGFrZRIxzKXZnN2MI9TTYqwAnwdzVC460
it+Zb2lFYLYSasoUD5wBzxEwgqkNapSpCqNBlbbfX2KRCW09+8dSesFl+Uj5hW3a
r4rNaMkCuA4Q3pSRCteqY10PzU2m7LC+g10QhuwJhU+aRWqm9p8r1gHxVmUmTFN4
OPIs7qRQhjxVAwrUa+cpaW2NCNCuXxcKShPK/uQn78NbPqIzsEEPYAxIVhk1eL0y
jg2kkWzbbUbI3o6XtFQEoLbSSqn6vBZawxXDeX/c3GFkL+u7s1AmXJL5Z/puq/NS
HGcqsqh+qXVWh3JQXkeFhrYk0QzSofX0nZ/jo+UToFCWdQ/jlV8z5y8zhrk3/Kr/
lrwCP72lUQpUMsMuoHJsaasBwQj/5hy+dnQ0UISeAJe6zvvZ/6dGDWAc5AbRZN47
TiX/yXVTrt8eekaFUkMx7ds5tlzg9uUPwtJDVjamW2hb6L31EaIwmjUbcvNTDref
KHSzj7VxzytAnQzhsw5X+b9t5GZSdBWjuIAWUlXSc1DFi5sEzuQfdcjm0Gcrxqr4
C15wu6fY6NpDksoT+uwJ2Qu3TrWBLDrGFYq4yE2TWjCTemlorE3rtcGPFWNBKh0W
w3uQauiaYDx2XRXaKPFtA8aFa4oKKfJqVEgwDh6AwWNxNSnQRL83kJOQSd11hqvD
WmCBxtpgmDhInai67H+0ynpRmbv4pAd5Jkf64r5WsqtWfR2F8XlkxiZxXo4vGVrp
At1Y/69If4QrAkajXVLlz+UMjSNYVlGPrLuZjasMXkPWNTkqLB7r98ek7CnzuZKm
N5WJbZLa9fju3b847eKJuzNp1IC7fKedwzzPPn71D4AIi0px1RGIMcTsFCM+Ow1O
Ww9efxBm3GSPIF+1wR31Y0mWGk+ZUbUW1xHxkyJ3zc6o4tUtSdX4wiALwCaem43c
/TAaCd//NQNLZMzZeI6G06GEqLt5NMGCcasXdejt7tfRKcSHiPaosoqTaGgb4K1s
M9uH3cpo06HsO3M/khLEicKfDOMYZ/4UVEpvE76MqITOgKWiUqjJZH/6wG9v8p1b
r3rPdojboPRu4AphrrC+wjXmOyV/Eaa9+o1MXYZat6tUKpAlrxYauJNEkclcW5mO
UpVHcm6oWCDckdrkAeMwaN5gn5bLx9IB4y7PBHZoQ+UGhH8vwKLc0MRIvv/lrBlR
TLSpfNd+mkmcXSRfGoKw1RPeOIaIQAO4kgOpgJh/jZHpNNrzovADJUDfTH3sRq2n
uC2g3TCozupzNBLvw7tz4WugmZ5w36Y+KrGxsZq+H3v63Pj2beJivI33HKNcfilh
qU71T89nns93K52UAFr+XgiER059hnXZO7ZUiP2b3r7dfCPHYCzhN8l8buvFlpBh
/9S9LinsSGcer9vESNeecZdzUhodbuSW41zCYVHnJmBZ1Wuv7/jzy/3d4Wkxzjbk
ZtSAtY/cbI7iaxO5si/VGZdDOo/gljjfSRArrEvZs8DDnYbfoxiI5Q/pfn6lfp5k
rhV3V6dD1oaveX0zZYBqy+aJZROztCcQF3+QF5MdjwNJ3vR3eJkhTekVyMImhU0y
54fd7U4t+KE2ZfNzghB30K92Xn/r9NGeo8Zvmd5N+aP++WwuFF2qLW011Rlx0l2u
pRKMAEQEOKITqwkcRfGacsr6fJEtiQjL3RX2+D/nCSF1/dAyIoaA0n0I9pUsXADE
e39lT6HOmGgDz0IPUKnE6ly8uGrcIwqzAN2JdjtuFin3xVQLIhbDXPl9nVwfShFp
WeFJfWvMOmB4QQuw8BX9ip5SmDvatyBNCKT9GajI4RDtTl1kVCMueoDBWyDIQqN9
6W5/lfV6N81RtO/Il+ua0QTJodsBseUlZZWq4oG5dkPQuxKAJT7VG6WRYLz2aU+t
Y0SXdzqJZOOwVcLAK1f17yd2NInuQXWzvAX3Ay10TxPLSyTkGcu3H4tDtL+CS4VG
wkDyautY+0/ImFKKjgA6yCKl4DZz+W11GjP0rbT4yxBYGMGSZQEj2dIFlpf6qirl
+Q4QufkyRyRTV9+fW2fytv81Z/bZdPtK18R5fHjEvXwhKJZ2cNf6ZCETzvA04Qj+
L3JF6tnwULh2oJPWfyLAQRLwDC8XwDpQVMV3Fno49e8irh+IuT9akdGNpAWzRRfk
mCyFcD2vB0uf3hthrp4DceY61I91JgmSxkVUD5Vbr6Gab///dD0B7N6/FkFlfC7q
C20Ty2JBTStb16HLVtfMiRJTuHlPEEN0GYdgYU6PRMEPMIbi3jSRpFN/5CIr/0vZ
mdJVWsNPE3Na0oIwMsTuB6BGUrqYVw9kG1993wIrhx0OEetV0XHC1bAKPz3u3vz2
zogEqzMt4GkKTtYMpeMhnAc/UPfAHaoEHwFsiCBmJGtV8KEv4ZI9j44AgffT1owO
V/l09pdxOUVtOJ4vkH14NCCPdz9cq/DEnevpbIncf+5tu4YryLWFOKgr/KxyngXg
Y65rBKJAtgEhErLQbXqIaJKTYJ4cPOTYYPqrPouPSta6hwxQz4m21odnAMhHBi8O
NkzLDu9UKmVme3O7Mn9s4qGKpT5MbSQ5hAxyLfeps1SgVij1dftycKRMYeqPm2w5
qU0wnxAT2faNpKz1KBKHoykKI+JWCM2qTc+usElik02TSzSs0z9IRooCN62RF8yX
zf3W07XYPAu185Vo2LDVUqvm5qAWdkjTeD8tuAencaYItjQ5mZzZzEYq7ZA+GHIQ
f8e5Ri0gOflsu1CCE5sw8Ld72TT4v5yiwW80DLHiMKG02nNCS/Frmw1T/rHW8fk6
Jh1KWFRRhy7/6dab/olSPGluD6sNKBBiK3PoNyDAD9u+FOUrdSpZB3nLPWQaM03t
eQIWNmiAnyZ/pC98Q/b/roVsvzRnjU79pnnGj0UJIDgxKDb1URstu2zSobgwwfaP
qPX9iPl57ZGkT8cpRsFUe8JfBwAZgm7BU6FNdk7wYtrHobAdHiW5fMCY13aDGCrj
WqMwgH69slKrNrQuS0dHUANt8ikbSb36nUFmN4LweMs+/NT7kwXseZ5QkRteMJ/r
8Gh9zD6yPt0ytJSHLQ9pBBVnBQcc4CmeX/z5pz/n7h15uSuXwqDjjPXXOrvZNSwo
8Kx81V6M0yYhgqgj1mfxm/srbOxSL+N9Tnt/mRUOeA7Ou3q7M7lvrcb2RnQ5FHuB
pWaGEcQLe0+YI0xyDlQZsmhazk21GFIDZSMnZ6LupIyaenyp6QO+s+qt1ywyiCO3
8X7pynxWo1DP0ICSZDMgoug5KZQm9BWTk1fQVEIO+lFWuXuv041TbCe11Ttmk3WV
8vlhskzQBFQ1H+VZbT8rhJx41yJWwpNOdD3sDppArPEnYcOWJVy3doC7Va+wZrzH
8fYwmW8tqQY6jImQC3BqXrIZ7LZwJ+I8V0UoY0NWUt8iV/2/pEsA4LVwRMRH7673
k8VzHaDFiRh5oUkh6f771eI31r4nas1T2BEJM/SBHS6BuZqINguS47EbR9gvOXij
0X949zRjKdA8A+EK65Q1i1Sg3s3MexHhh5g0HowgZb4KApOF0fwEsNifPWMiYVVM
RNjU9kcnbXSf20oVpRoBNJZ3W1EQWXj/3bmP7u0xW3gwslrzQxgXYH7+58gORQ8v
CCz9hbneH5vlARuzH3x73P29e+jt/Da1tYoqiSnte1Mhv6ywxRwqRNYM/gFDex3M
oXXryCL4ORS98AzMdjsReqE18ndLkOdJHFwuIGIHTxBuKN0orwc3g3AmdAgdFmPS
g7dscou9HCw7T/4a301mdVU2F+rZFOC0lOXqW8SOXQKhEzygJH8RpQrPvqS1leNs
Ilmb6rocERT9L1gQZK8+fQJKaixuSz7cruJJVQWqeJmwyBtYtDQuVIekaI4mwXGL
wL0MzHF5IRmMWUFZSrw9ErJ+k0G9P/2Wl1wiiGqzlelZSIkJ7rU1PIssR/hJojMz
xnFiTimG95hGHPYNYtT9miMwqlZMZI9x8KRCP7D4JUNYvUg30mUOSogW1ZAeo7lP
aWbcPEPzZQoNj/HdcfHAQnr19/WNtHBm+uhnxjncvIM9iSJz11OdiyJYAenqcx88
qLJik2n80hoWf90qyZRs6GKCNFXFeV2F03mVccEFmYNwAV+0z1ycTQxloqb3hBD1
NV3xe2a2B/QxAklGBDN22lCjrOJ1Czkx08+daJthrSm1zMjDsAGsX/Q2r9Tlg4Z8
vAeBKO0m4fIDSlQEmuSLr9DtH9WJAz8s6WV1+2Me/QQg3ZOA1K3LiwIOsbl6h7jN
YtvPAgDhErlsw+Pa+zJajlsJqZvTNFnnvUV8+ZP0b2Q3JaH51OrPisYebR95viwi
uC0Pof5FBv3N2UVCNPLxsJA/gHYVOf//dV2fuEjeCW3xN862kNYEInY9oTlGL+u3
wuj2TxYNVGS7M7nKqED9l4zAxb0sQUTA3E3HPh8nqMfkcM6EQUXfVDFDohJcgDN5
A86os3l+yOEkZZG2kwXgJKIUAogbkSQcrmvLyuUeIJyzGzRfYW9WWjfKLlCZUBXY
Lo276Iws2CQeky26+YULNJgyQ1TTJedr21VtHoXKSJC+WnXdjLc22GI9gnvJNTva
rYQIwEHtyToqs0kRgZ9sV2t53JtYo94b1zJ0CSeoKq8bqHU+HBpNPKfxvk62+0mT
5U1cCXWseP/OykC7fCrgROwjYf7dSOCYo/SA/4U3AmUa5/9NSRQD7LUxTcZATSvY
hk0mRwhB3dBoFSQgrtqIFh5ampworMC4T0lEqg3MK8zixiuYmGam2/uovUeqwBK4
qs6J80uB87DZHIpbY/mxh88AOBJDathYKXx15YNmaBDmlZzYgmA7AaDKarhrzCKm
kWl8065aOwKTEdVFMlmNPlxn9ggmBAyIy9t0DnT76pIXd7SPzt9+EDDD4AhXrNvL
glvSlvheDv4CvJKdkjcniWsq+Irulb+50UvoaQGW4UW4kR3Is5lz9EQfk/Xnl3an
04m5w9wNVJkDA+nrzGEpD3gpE+nZbGUTLMP5n0kOXEoanqUYQ69V1N5LNmNxVnN9
f4ONV5ZFP9Q6oaMPkwbRkolVAk8v3XZzBpoZ+lFLK1wkPQl5cqDtY05vRsDJzHua
AzEgZD4ExsRa+Byii6kfBtd0kbXzwIqy7vinPKPbkn9uC9Zl7bzOL4bMJSLPj5nG
hFqbvPWokeR6uHvSX9AWHauNFEjeufNYb3P/S/1C80gcimm6AL85OqzaczRFoyyE
b+TmIG7n9VD5YWZKlF5N6v0kM+IEeyAfmUDpo/8KQbRSjff0X/uB6xTEHijE0gtT
NW7fICemsXK4qZIYmYYyyJnFDVVbyCVWH1vlSwcFNgY970AlC46k9mgpkEpUjarl
QgyWVs6jWmBVRULf532FhZ0ngJZyc2jmmjmS0tWAXRA0o2a4U8mP2NRBy1u1ln9x
2Uxx55tuT1P0JnKIx6oE45u33TF55W8qdJ2tNthZy/D8GQqAgKUqQmlH7HixeuFX
Wd/GUc7cgIOEwbBVix9uSNzEwNPUtaGeY5I3gSOr8E4Uhpn/CC01X8VJRZs/AJ33
NeJCd6hH7beclkR6lXkYjDrsUmxnfWZr9Nd6ZUZJxbj1hMJFvkJwDK1L4igwy1nP
YAFMe3/sCDd+MCxDnZJoQ8oaWQqO/d9s8fTBAMHBQ8rvO32vtoNwpRJLPAM+vh7r
wFCEu/d+++gcr0aHBc57F/ywvLcywBMyHydryxc4koQN2EtNPVoslk+6DETAfH0y
/9tnXzswpEaKfSX0f692ZZPsM4a1aWi4RaVDp4UPllWEEkAgZq4x3R+xK9w9DIgK
QC3fUi9/+y6C4O8MBUVM5rg5xfBctwuauQQ3DvzlkpRku7JJJzxPVV/4u+WG4AM0
klwmAUXhkF4vkopV6SHqP1O03Iidp5NpqEi9Ci+rTuuFrHhmblTYjWLz5miZGWse
qfJrstieHVms7J7Ex6f1WPmqObX1N9Zkkzr4pWczMJVnIgDhFAWv4wTBdTzAI0JA
JYtc4m0seVnoIZazYxJ4x79IC3afjr60T4HLRZ8gweguQlV1gbrzWQXlws7MtL/B
EBy8sg2vr+S9ykfNP2rz80JL2ScrKS1TiDIFvVJWxhH+C5BoOmZ1iY5GnnynGUiC
aqOKdgzafUgUtejsC1SYqPrXyj0D83lbCmxWDFdnPW+YIJfsDiWKfijAKL2KUAVd
XdxdbeRiXIHcO/UTna2ws7M2yzNABkLLg/ib+aBPHFsHySSCX7EjcDDMocZnczhX
mw5M6uplENKaqHa4r7RIvtxUy3Cs5QnFrWn1iD8THNtn7Kotmuhc1cCRX1gpEEnP
iufP/r0NtvcSznpbDStnS5RJnWHPv2l2nGLnNoWTgKeCgTZLuRwx+t95UHISIUpG
18xVtLB0LdcdKuWBrs2LJBOxDNc4U17zxWNmuNt4LLpAxrmM8Y1dswbesznysGz9
rkggTm4HqFFot0l6NiEHXF3oL9+sqVMwigZ6vkjKx5nLWH5+T2XVAvLNDailg7fN
DCm4SlU4CYBySNU8FvxgE/Y/gzl/qy0aQSPvL4L77w9T5jem1gqL3Pzju9f+w5ya
szX6FXHdEGXeOe8IVXpZQXQ/Rq9U9Y/PnKOwUExIwTz9ZOQj8Vu/vwi7FY6Cau0Q
QcbBMBhGvehQJzSg1faSbLUblp2gW3L5us3HMNdThB0wuPcuS2IYNVoR+9T30Rg2
BBXK3H+4S6M09vMtbRCcz5IiJhRrGbxvY9L5iSwH4BpJl6aHOIcXnIlNr1/sWTmK
s5ktDmGXFIuHYOib1JoO1sQTfRXCfvnlS7q/AELWkxheDE5IT0x2UTVhetzpd0ct
GFDKFpOxp9uAxHqvaAylspVKtn1bYriMIwUnT4BRmHjKlJmgpFDAVp2Vd11gLNPf
pDkHVJNxXHcCX0o7/QsTiVL7bqN+2hsGFFcAo6WBtPhUeGiH7o2P4L09Khy4YVOw
ro2XlxJz/atKC6wcD/UBHJt80xSkDYdKcT2j1I6EVjoX+idOOaGSxZmFaGJv32VN
x7gyWngllCFkbMDm9QBO4Cx3wcHnRiga5V+yIefUnAaiJFCb2zurzrP2h8ktnHzi
G6px/2Qlu7XlbR5v/0PAJ5hFqVKntGIBEW3UgvdaBEcE9Gi+KxLek1SmnAxRFu1I
5cTaRiG6IVaS26x94LL+lZ8l0CYW1OxZ492WyG1RLWF/VzthtOkJ0Wy6O9TEbgx7
xQPsyjsvaapSF6IGJDvmuRy+89YqUz2jvD1wWWoTzWoajyRZbNo1h6Rest1LTMXN
/dgB/wexy1wXhLRGY01ZCiZT96sii1GV8kx69d/wgEVWA7v29xKNG4k5ZQHSXxZU
pfjIgCUZFURHEPpeB6AuM1wC6R3z4Cd6Waw7n8NllLOOsd+YrJRFq74BZxQUap/B
4T/X6T5nP2AnzG8yTEPIvOfZWG2uC3wQQbqgiHyrBObZwB//dskm5b9vRq9raUlw
CMis+83WYYGLVEfhgnpdY/EidHWSAEe8+L6L2Nak7rE4ljCVsSnyh4vHuVvKeSbl
4/y89mQ1WlQ34rXblOavRKlebZlDxJ0GgsuxW7bcS+j5DvhdbcrSogqmMGBbnyyN
mPQKHDDgsMyHLCmAqp0s533lYpn/6KvK86PdsPkDE28vr/3Zpg22YowU6o0eIPdV
tIhd5Y5YnOnL259bNSQkN2mi0hOh9X925u67JeJrPVceH6uanqzgD26jOsN+v9DE
j67HMJXIzBkye7htAYjt1rbscyHRJqKD65Vip2bWPvIe5ghwzQFcH/hKzZYqCDCY
p9YdYPF8ApzGOXk9hMqFhXGfhpTT18twzKn5f5xRwie9usKzSCwDxyTatQFfNmrF
p+MJ45CzlZM6QJeCy289Aan9Uuvw9rZFx2Nqj45dOP5+Kmm+5R//7d3yJUY73vxk
aN4Y14v7SGpVEnSQj3gFXqVZ64pTe56ZiED3HXOzQ9BADMkmXsh2LJjZZZ7uboQc
n5iK7/iQ7aIKcg8YB1f0hd4iDEYOrxcF+pDCKT3yMcU7lxtiMsa9Ca2slsWBDoom
np/RJ+9UlfzJcpIF833p6KFlXdNnzSxeFsAc+C44c+0N1VSqch6tyJ8yHmJIVSuS
BdwCrkAMuhAxNE1EU0ZZzvHd+bXD1GCFCeHpHn8XX9GFFgeuh2TIkoY3zS7n3dPG
R3EIZXjLypCslPBT7SeZed+mU7QHCL19m/7I6ld23Fv6fxCyERGsFbQjeCYeC7cf
vGaYpP0T2e5YpoDcb3UZXQUcrGKLCB4aQC6h0SeKXkQSPg83aFSbCcJH1csAjpQk
w0gSGhQncaBo0yfrxfxyGdh9agsQEyWc3+gF4ZSwmZEOTOn8PIzVaQ4XK0B6ugcr
AaneNtw+B6L9gf+S3TxJvJydW5kqk5Kr6wPSn4RSfUyveSn0lkrMhBV5ivyjR1oR
iJOdLdBSsldS2N1pGDNFI7LkKd8WpMS+ZVqDuujrDnB7ZSgTO/Xntm2owtW7vYVE
/JoT4aO5df8eLaCVibJ82TqF6TDqAeyP3ciTbFCCzN25foJ7bNAnEvuqFrNipaGz
LsFQafLROgssgpgWmmUEkXjC+3bRoIrT3NHIl8L/oXiMV+SwVmtf6dHCjE2iNiyD
DM9L8c4GLxHS5oNVmzE4o3vSZHwxYDoedGi7bLoGMPPNs9qH2jkd17ZNhLjtjBq6
fayEw8d7zrf9i4HlhR+PBkgbOSaQlSjO9IrKDW29YKr/RTmuazn3DuZ/ZpPWUOlH
jqQmFCG3XkY+vmiGu64J1P/h03QgkclzD4DaJwIehwQSBgJdSqgivwNujRhsL6dE
fs5vDLcO/iDiGSkyIGgM7a8s/cl7st6QM4T9M43AzHU3WCOVKPlCMwTlcx1JaMAL
hVqjZxNQP10wlwKwLDSsvQMsOBi4Zoa0O32RPkHHjXU1Aw2bRjy4Li79wA35+bV7
fm9SnEe3ZZh+c1RC8+fRq9RVwXY3md5YnzDq/GJdcR+PVUzzWUEPyQdD7Lit2nZZ
lh/S9NUFZOKctaRH8nVRVBxUgy/GQhcrNsh2/mTTBtoU5RoUQE7UNTK7EJ9ht5Zi
PmueRZTogIbRPmH/iOzy6Q0QDWBJ3kwI3Z1C3SdiweyQHkzVLRAwB6794DIM2Qq5
zgR+AnTkMNF4DtSED3zK+qxxdPcrCdl1YvBOaD/ejgGTk2lTyZK/E8JbeqflJY1h
wGI8kx48tLnt7Cmnbn3HcJxXJXibPuaJSyT3J1aHHcyf2fbL795loAabxT+36RoP
VIo/U6nbPGY6kwW6beR7Ffa6y168INN49kKVkVAijcBeD9DzGtfz6FliPPPRbdW3
UfwoQCdMpk9n41iLUo5y035XHQt3n/5tN7LuI8nodMi9Ot2ZDhFfZD2REdXNN1lS
7ZJTlWYx9Mo9FBsBpHx+KOrg8zvtwd/E3MNuxmSkHYRbJJcL48LEMXxrSnk7HR4i
CJu27Ze1LbBg8XEYOaMRfUXV+4bLQX6T1lGc47Q7FP6K4ScrdLudhtah3SpDtiEC
/LqlXxwbHntYVN1FsA/EebfCzQpnvFiTPIATdslUVHnRszHPQFMvg/ZI2SSIZVpL
mQCMe8rwTMbubc+jz7+CGcb8AXCZz4535iPN/EOy8O28bTWaphoEXOnIten9hD7v
xa/QGVH4sndfQiqgebtvesyeKZivIjQ5yvynTSWKEdQzok3CPiOQFVCGkp1I8PAp
fBliKtWo0isYe1AsKxQDPGcwXkx2UySDs+8lNY1tah6OK2SRjbuzKruw05SRc3p2
MrNqfs32V0o7VjMlf8UJHto+lYsO2PrZ9xQ5vWiesywtVNQzu52FGn4/FoHT8Hy/
LQXlRDTl9k7RBbUMVHtFLUhmFSqfM5sNZ4klZuW2q1243qqnRjeIVnmtijQKkJ7U
mVb3a+DzH1fetbwSQ2QDbNoxq6Js/5YAtV5CR/QX/mQXWSOQobbxWmod9dk7RP8z
EYdg7OFLELaI+Z4r33LO9FJyHhGvS+CJjfF1wjB+VdBToFhgOicS9GtwBKmQj0WB
sBN+4Eah5tcmXn2iL9+pQfenNLkoq6xX4VWk+gAqmPRA/eVjklNLgAcSsKh8/h3m
m4hvir1xdhT+dsKOc+HmLhlxhLEGTcrFrSCkHPmPvXx8ZftYzwVfQ2kEITQyiEfS
SRZnj/ZwjUxom2hRxxBq+D7imkhbsuFXlT1ZQxRxTh2jX+8ai9V9B4Oji3BMNYoX
NONHv65p1K7iTOqsrqoBacC/ymsNPD5WlSVsUuisSrtqHpDo424D5ycMSn1DWvSK
PVgVS8OLLq9lLyu6FaAdvdWICb/3h2VEDZ/oOi0QOIqujQ678ATjA1Nxm2bLJp0h
KH/sy+z6JnGGPk9oc5gc6V4ucOfaLIPeC+g/gaLQvIX233l/MC+0lskGb2sPwrd1
hCBErj11PLtV2+XRffArpOiFICxIu5zBxMPk8UKdKaQGj7dMhU0qBmA+2cmMSf9z
1MTcnoKiBC/rWiJoxbLSkoyapM8kWr8XQBCslWcxKAUxNCMyEgarLwvP6ufmd1Fy
mw/jf1QHALRNtSmwDsV1P0be/YtOYNCfuQAcWnn6hqr2rwBi8PzvZsRIc1cUqY2P
OrWlGxhhmPm28gK6/R2ACHXkVO+jNLpR7avbjb+qvw9gr/pRhgzC3B26U5hVoEZ+
dMuIYlWHh5qpjz+VIfbLV0deqVBMf9RZf943CmjBxlF3efsFPtq+n3L4qeR+Cuv8
tVZ+aFI8QNuNDlxRuGupZUZR0KBNT3OeFNvTOM6ZxPOLgmF4e1lCr60KNlBUxr9e
7dRhutqfmfr9sshiGrFoiTJdmNIe7i67PfSpbakLHBdOp4JHdIvthkZarDQkmXtI
VX1LQBAUQUIgexWwuIa8MO0LXl/BA0Wn5AxL83IJey8k14pe7tncLHl/72Sxsq2g
PtLlRJNcjh3v/MA1N9dKYqLl+gq3y/DYZ8hKh0J60vvSe0Rb5VNAOG7+pkq0qXM1
4k6JvxQKtbQJCYr3ukjlfuFWaSht1d2+TfZ+1OWPHxz7MLoMdFvNqbrXZLq2laWO
6OLvucnqLovTDIX1KAGDa9PZ+wFob/ruC49iW3PimX2G2/Z6Drsdrkdo3K1gbK5h
KxTV7uWCGM4cI2hVOs3jzFaXNl+xiZG9F/bpGIe9HAQAHk7VnwT4bRPZbI3GqBMm
rzBvgauKtL5O1oyVDlP+tqo6gRkbjFjPErLNqLboOQoMez2Ok9Yir9sqNnXrOIr4
1uxMZ1eovRbBxHEAx9LuHkbHfKpgG7iFxfR7jRXg5eqfiTC39nRQAOAfoZi7DG51
YUTCkFBtuc/m8HJcA2YV9UEHRLkrTEj64l+z5y4L+zGb5k6wZjUSi1L1sI66/nbf
xBZlbR8djc0p8FJZnr/mpa7ts7f53yomS6UhsHBBA1WyrKOfoAyttBCgCp2yJWSu
qcRciMltd4Co2UwocufT59z8d2AGVCKaUGXO+J/fD82bFPxMjvEmSn2USlbNsMzS
zByhC6EpIcg7ek43SX50mfAn6PsLBDTVk9OuSJr3S/ohA5vvBp5kM8J6wrBbT6U1
0sDIYWelNLp2xIalDDrBlhEMf/RARcWjHRnRXJCWBpSuQrWvMtzkv8YlBCt3pHGA
4Ilh09dsWMgsvqrcv4hXAvvcSxZD0Vk1LkIzRoG9bm+YQCNBA28SqsoYwGlS/rRn
rmCU1o6ivncCf+wZmgcY4eiBzApR538mTPYtL2DOBmeP2GJHydBAxDQTwLEdWI/D
wEC7qc2wqB0LHdvz77yC0D138xjAK6NcU8JSjEeyW2W3f9ba74qdDiY8fZNxGgkd
vIVsEsTGYAx+F/O7llWwyHclQA1rEXiA+1ZbBCaxSZIqNIznEHZ5mAkVT43Nf0+E
n9RjGlyjz1uV6/yQ3TEsLZy3daHI5GXAlbKhzEj1R1SwN6pWi1fy4Ghox0ZVtPp6
evufRWBDpyOTvJvL2jELlEos/t5ExrOGtReolEVDedMKDQPboVOWDZlxdKeKIrDa
lJxICUFUoJGB5TynRT0YV6B7f2qoPrnry/jrYyBmx7k91FMcyJVM3I0i5b6Cx4+l
3xnP0TpUyqPdiDE4l9dWQI27wogSqokbQI+cCq188zjAygCRENv9TfCnzGAUkxFE
dhA0n54J5XDnIeiA5AN+F5NCSdQq8LfiFiZ92X5xLp3qHtRw9bvJ+GT7iqq+mZO1
DytBtZC7oGNp7jO2gZj/PPnvaOuJRQWkQI+trY6IzcPhHkkvDAb0MPcNS/LqGp6+
Hmi+FNeRfRmxQXMReAOMAEreZb0AU4LHSqcfuEveEWbfGF103tNv14mSOX0zSqKq
7m1R+sVTfIM+cjrybJHyzurUu37mq06fMW+1341HvxecqTtUef/ET9XOAWbVvw+Y
itm/istQ60z75U3ifCguBjgGSPsWOXVtUgXNJP+Sbv1GqbHnk/MrtTbI2ZKoRHqQ
mdBeIJs4YPKyVd/uV63Bw2FUhKd/4E+N9REByZzqi5x3ZPXvSJluVM6FnxD7nCJh
ODUMvtlNyziK1BPJ/rVisO7TSMyxbvIgFaXN+X98gCrq3lagkaQedMIB3connWuT
+96tfTFY7WC6M7OG47bE9GM5Tu5Ia+x/XYz1z9olWUPxIX0Pc6rHwpH7/yXgCGbB
eX+ZZu7gsXuvAcwGCG5mIWbvxsvoRIhn204ajGpglRmlDmARG66XmA+5kUcjkyZX
s2ryuWfhpDyysDQDu4cyKHMuSX29Hxzor7+EFBg8A9Zcvazrfq42qlBHooDeRUiO
0oZPVTW08B4xc2CJfSeLJI5f6uRijBqMhf3x+4H4pQkQqgKsRfcKcaeZafV7WYpY
MLVOwFBYUV1KBG3hJO/ohPNtaBBTaLfnh1fMkOuCj1heFbmdM4bEwysFEdGfA+ge
6ddhSYt65ZZnhKW+KJz5Eet4Sy9E4+KW3R3tRMgFoT+R2U2yH36RKjfaWHuHZc/P
ZnxdXZk/yIg3rUSskdmTiVC0Pg9my4rlqt8WALAxdxWWktYkyHv5eUfvfsCsjXgc
h8VWCrDCU1ReYrjVIPklzLWhQf8RVM5XHW7WNA9xpKgT657+5ZVGjXk6HSDSUT3L
NR9zWYSRPoylCM47G8aXxzFtrKqlnpsneZ56LyiMGmMgx9ucLWLinNVf/cHSEL+d
Lsz9NhYEad3I2XRT4l47kuM/Eca305NubdTA1HiBJHggyP3Ocmw8k2/sm4doUZxb
cOkBAcGBMlS3xs5YcHr8Lm46ho71uwkrUazB5TfEh5t7Pa/1uN/hORu69BNrOkGH
JFud4/9vURcrwEbi5UK04Wq/Dx51Idagq6T+LrEaeUr/tb7lr+dQMZr3CmV+Lm1p
gZQK43ie4hqxngf8TRy5xnO1pkZErqayLjhJsFuXHX8K7RYJTb3/RzTOI0jgHuca
2EQ1uZkO11h9hag9e6uy7TU7CoshsAMSN0g93BXL2H3bw03slYTx7/E7KzCNDeJ+
CQnt0Zvm8E6T2Tdy3oAA8VTbBHrCdGiyvbCCTqYJYzaat45V+GxmBwSus6VQ/AzP
Eb5E5wEC1dPS9c8PRKSEy0Gqsb+VDuGmg/9rjh2EE9h5g65BXuurM5mJlV66VU9c
PI719BExKZ90/X2sqsEd/mYhCkv7lZ7+pnLZUbNz2hoqY+brwhsxOXbMdNbxvwqg
a3/zJa8lHERTnmz2movsvqaw3F4hAP30A+Dm3eBVhba0twjkdRi9eDB4X9nhBqDq
c2jdicBuC3+kAZlvzfVRdVWa4f5mqOo2FbidJxFKP4i3kJrlDIEJtTOfAQo5mcCb
0g8GpA2uhvUByMshPKLUKJG/LzfQoDA9ZpcNvlxnglzpSP26LUwwFOOaAwxll7c2
fESgRcqBnha9qyGvDVDxfbERqnNxc8jI8ALcvw2Juzy/9fFQW+aRA6OLQJeUFiGi
44rfLsxlUKO7OmOvWxxYOs5szAq2MlwsRGsNBlbuv9oeEu/oOOn+CVwspSOrYrfI
ccoCjwJiSRvHCM5IxVP+s92YQ3fycsB0J9b9k5UsjlPV2YxGv+Qe6ONWy3E7tzoN
e9vo4dhkWYeYjYvfWS81mU6NBWZH9kFX/udrdYcqJ2qAmAZ+tXhu81C/puebiabl
F1Jj3B4QqLZpq/8J7C3ZW02Cnz/LUS5JQhCvgenJHveq0IK2xQHPm+mwyans80Pi
og2SgmMWpIIo6FATeFNbCBE+4kJdttNc8iMhR2wm08Ka4E1e0egCAadlZYCdHTvX
hjI0d+D31M+lMb5QpHfrzNS5VQnkpiOUhvFE60H2j+f7uJWbu25AMcoQr15/bfVb
T9duk5F/VntxjGWAdLQ+BRFBjuf4e9Mv/N+Ap3eFsBZCqQP9KQXNJPgTPfD+aTv0
1PraOhv4jT/9/UJ3NDPWlo/cB2Ux8xC+VyUGlSKRP2jjPwaBhjMIVuCPJwmbdXa1
z2l0Oqc32fuCPWep4NXEQFNVpoq10HoczEKq7ne6Zuv/6tqJWeCErc/0WLt/rajg
pQrZ7wHnel3im2wv6XfgLr9sbEqNUi29wGcKOoAPZ/SseHVV8XSG5CZrEUU/3Bcr
k3j13Ki4j1315CqV4YexRMnKbLk1Mwc29LUhFEqfRKZnTNmYXmR+osuqTqRaOMWt
3gWd9LVi/byNMljSG1ebezAeTV1DrNa/xSieBHi3jsvnbjTKy6oYab9ztb2MDlHr
giwMURe5iYW/0SPltgMkdVHdT/C/RKK+nvSK7FMtZ8pfLmJm4VhEtxLmuPsfEQow
AY/7/Flc3lwu3JWc/eyHVCBbL8d6moRQ+evp5bqd2KBNphTp5cHj7UTH1711rEUS
ZimggnAGhiLxgEfRuWFzs6qWE4Z4WZqcLoCZlhBwmoVpzh7tDD9wmDBHQdLtQFHN
I1lsSg47BkunEdqVNiZloxRLNB9DSRDHzHYPY91kaygLK7ZCvAf215VWj+IeKYlD
QxWB/2uHDD53zx5OOiWbDltProkZBTwV7o/9dNTTJkDwDSuSj2ERyVrrvxqeqrNv
UCZnGgqfwmCWToBdshA0IqBdZB9tDxvrgmb2jtQvN6cMkCxi8PmGz3Ec2JKHdGkT
6TL5Wcqe9HqNZbCfy8mR1VJfuJHbch0yWpiG4pHiZt1CMFt4F2SQdT25r+jky58i
iiuswHekH438g1n52bSSRIBmdgtezsajV8nDL/fd3qZ8besBAJsx6AiU/l+DHqgg
Fuk95MKt1142p7UHbyWbqHAQAzbRoGKrc9d6DAOOlpiubROEoxLjEN/DMVhaC2Am
d+UDm/JwcsFZzqR38/Pxr38Q4o8gJLde2UUg0XNNmcCpMpcj+Ynviu3JeOBQJQNH
/JYfOZwBav9uZeKLv8dGAnj6mRvoybz6EtwcKOcuoq3JEPCe/2mz9AnZFVMpGyba
k+F2n79DIKvbMzPt4Le7CnT7R8nxjpoaUjuRXxojxrxwYjHQq5A31HCHGamDiOXC
T9Zh8tzReDsQpcWzYZFhrQPjypWjLmAQ6ZwNa24f5FNVi/JLhQPZIOQkE6cTueF3
Cx7U+Gcr8FLwcyv0GYOGGALl+Pd+9NK4Kh8YiqBLn5+QlWs9eaeXtP0lw0o/h/Cj
u3mdjPPMF60AdFeVBU2j+KiugQaNY6ojCSb00lV3ol75AujmhMndwcZ6oyMbPayc
fI6oLN5p6Cm+TPyGrhaid0/h6D6ZyjBD45AKiR4xg54aHuhGAzaW25HlRefpT6AM
vX5EuE472mlFMxsDliaBTEH2Q/6EQQYMwWN3y/AKhCie38ha4sWL0GfSuiIWSrvP
XHqwo8MpcgAYvP0YUz5Vm0m9+3jiPWrjCfowr1tfeK16lsaPJYf2Mcw686vmREs+
cncJwHvZRN9Vx2+NZKWd1RnDMzCG6nPBnNc1qVHOuYXW1aRoXzekGgJzdWPEve95
gGhQHbqJCOmC5MLZBoFNWMPuhVpTt5fIhAJaUT90nTRbZSu6kQtFEeHCUdXrTJe4
bzYjOIaITtYEJMPI3ngfXxp1IaUZ7kzJywZ85eIBmQ60dlU/8mcHrzpUobzWDCpd
ZiCSMERZIQNAngpIM5cdIVEKT7ty8jvSiTdEDmUytQ3glgoNihhTvkHl8V4vX6Rv
zclnCUM7FK03hroLL2ksZ0CGz23nE7+FZEB8nd4btDQMoWPFScvwGXA4w7Ipml5l
3/aVkZdmd+A/0IQ6s8gkY9ae0sNfQNcs+aaAMMSOhbuEidjjtJNgABXE9liEB6/g
Nv3Z993TS/K1NDs6dfD8jtzmMb9x3Iah7sIsabiEtZr8cv3JMXTHeEFom3izHO5G
rWxGlfPJghphNWcPm1Im95WfkP/dOOG0LMwi+3xmC6HBYfVVBM1JKTfLXnAvKkLs
zIIoV7sZ/0GBHZpSkIXz4KcfvoFEV32oq9NOPlHS8OV9lw83Nqqgw78aAnmMIkFt
HeXCfLFaf95twnpLR0AM4DTZrIcDIZjfgVCJkVoNIwhmE+f7nU8gQiWC1yEpmRJy
2BFTwrRsj0ELCg/dAlKJRu/Vdwy04FLBeZJljJp1B0oCjSModNrH3IuP9ukv2bxF
J+3Tik7pv5EaqF1oEw5P82uqooDfMAjnxkCLS5d0RevTaXqpEQLNRryiKxMOFzNP
umEc0lefzJzCm5G5iNnDv6H9JjLZQ2Z7JPihiip6tuRF/qt1fmcWzdUWeqiAHkzs
Uz2QddcXFpLGVE1vXQCKtrH33WmZGHaWX9u005M4908B6z5dNjDpat2XkIdjNXOl
ffISmz/VECmBHKN9Ty8LDvl97QamGZLkDr77SxYPldhAyzddNpy/kHJqyPHZDtaI
WlOSfO53p/ehOCFBqegpyMjVVgrMspsvB1aeoxG8K/+JHZ0BFzSU8GQ/E8P4Rl3Y
BDzjutXxrDV6AFdfHlvOX4YvQQJw2iMqOhhRTQmsYw0/f7LmSr2RG6LpZWJZyUh0
EAx0Pwnm5RBzURS4/DZVwGGZGDZN2PNtBI7NErV8lbuUV/NABoF8b4WBnUR3/4QI
E7vZ+/ArrLkdcHFP4R+WF5QaoE5jFcoLWNTMIVH+WLBcsIV67iaPCKYGuOoF3uat
1qGd/SDEgn8Eu3UYn4LRmEXYM0h3xPxtVbl2azNQHqdhyOfC4n/LoYUcJpYwDHdR
oihvYQ7K7MDNW65hDcKD3SqK4Btyu0f8xvFxtoDjUsCQhe9J6729piL/iLb46XDD
9UnwN+OrMfEp56Sm6UfYBLcMLchtNB43aAqOQH0m9UEJWxc2afxCEZ1SXfxIgHhq
7PojzTLvc78dR7GODtxo8dWDphrtc0Ou6/siKfIcUP8oZssHDmzGixNeryhwzyTa
Zi/L/5erNpd3zz+BWxWsDvzi1mDf2eshlfCqeCDss2rpWM0C/wxSweqvZiFhvirK
qaVWehb4Ho5BZoWKKmDU0vTAA6j084k9t7jNlF6UmbtYtoYSPjtJyCtm1fILbYXn
icnO4PFpDWfyV9XuBrTk2glwu9AjwgVmWgryqapnlSK/TmEbrnljQ/JMDNHtbEov
gybsY6g7IBP4dsQTpTOYCkSb6/8ZCWML++VziD/QcL6tfAXDYcCCfaRvzBQqf5/Z
oxydrUVC45h8wc84MOZ7vqJYIjhuNotOtebcvJB+fpQ6NX9RDlkCamkSB/St+gXm
sNOo7adL7ARw7Dsa0RY+UFLdJlVnqPLTX7j/AIqSzX12CIx5qZcXnJzs3ksO4ZyE
wjJEnqmn85jqqptz/dcenTt+6UNlPGnG6kbQpEhn/P21/JfatiK4ziaOsZ5t2hv1
RZeSo2baeWj0LXA15LYVNHDuKUf144ivVAflMOxs0kDpqKYLnyjjwRty5p0/F0Ko
ba3Vy8XJm1ODigcJ7FALQmcr+9BwbGJCmCIc3CRlGrrdCsKRcFba4juR4KU6e4wK
aNzMcWUvGXVpcnSjhACTPV5IBxI4X+vFWLx5QChpuVc2Rh9z8hstC298Kaj4Bvse
VNF0ofsnL0om9CkrK6xES92KRcbcwWhe+JBa/f19P8jsqWnjTegm7x5lK7S17xpD
8LgqiBhXH+qkJVZHE8q5wLAIm+LIqoByJsKd58Qhik7IsqZa9ES1ZQ8rTZOGoShs
QwmJEHzHpI6sm2frTp1l26gVChQW5TQAfttgrptc2R/pXWWKNiEctKaIgQi7Mzkv
SbG712B5ABaxhy/pkzodTt78VbJmvBtCquwKNvmHaMCCXJwNXCW5bIR+32ouUox7
CHEanRUZXQDhz1PeMdNdxormnWX4KdVgtThqdZcmPdRTDGPAA95HnremlxkWmli8
hN1FtR++SQSue/OtSjuLl1ulnJZQIKwqA5aaPMBkUR6w1E/7r9SkuOtDtqmnoqGW
TboDVD9bECWoake7B6FTUweQS/TZJhWhJ57XXTgAlj9tGG3BVMbkCPaMZbLBVHWh
5UlxDFU1KtgtrOzN8Q9f345fQ2eNhpeOr+OTErGugPuPvMPMQMV/weVDHFisvtfg
UA47wPu7ubLnFtiDbcZN76kSf0LAg22vfwS6r69wrM8TycRGO3eKC0C4NO9ZDnLm
FTvwyKwXSZ/FzmQ/uSy0rK7RZGNqMmVRfCkkLNuJabnfC7cvn8w0Agorfvu4bZ5H
H0PrQrF4TuwhS3K6lGRrUzY+oPeuglnZdiQMq/fxH6/L/e4wjbyow0cXHBUdqtuU
gNPiqzz2xaZoRIGHZ/Pa6ecXMSaSobPD+kiDdMCcuwI9yyMqx3om4vusbj3uzV3V
rvY4wQClw26ENmoPgvqNmrRxIEvl28QADOQlC1XDmI3TRkU5tPUr3UJerKmCYIqj
iOjvLP68xccGL7+LqzKJkueGLq4nvUleqUQPrG3Bm+eGWrWRvTTGGEv+JwAEfOlH
md6ETp6gwPdmIgKXc2joAbyCpsZPPipYZgvqRyN3VuiEf9Dp6d6n0BP4NIZyg/Z/
CtCWOlbnmZICxqmjrBccphrRL+oDvr9aR114SDyOHxgBl7RTMRT8RnROJh8kRmoR
GQ/4Sx6j5SYi/zDoh8nh0PqBVPPkIKY2cyFRnJB0O1XpkyDXFovWfLYNxykvz0Wz
qlvYyxlC2EV2/iNQp73MsyWxwxDaPF3F2YaBbAw/2h7jc4Fqif6gBX2kNy0w0gdV
TDF5IzVgO2Uc0RuzQ2addqOpHQrF7IJxxacGcvEkcL9aBw5/66BNBph1lA5PabrJ
cYmiQAsVQ6X4NYUcOQKq1PdV53dUQ0sgvIIXIA4A5lanutLlHtJZ1VPCN8ucOB2c
Gm003EX6zsHN/hf8Y8X2MZbWMhILBjQkws7xAn3yl/esb/Nm5eWDWmHkwk0T5BZM
LF8lf4HYpbZXFITUZOPsydnS0QPXrN3crdbCgdZsln7AOe6AUt7+tzVkou8wQE0f
DtoTBmg1vtjUN14CdzfRI1Rk0RPEoUO8bNPVrPJ6Wz5PNtU/+Y3OFlauT4egMjGc
HILqwopSYA2NFSEvw5vbvbqeslI1dKoutXI6Yqj3yHP6ZtlxpDXTS3+u0cwbVT8g
7W6zde0RBTH9rPKH2DR6Q0X2Aqw5z7R1yJfu2xjE6APlztwURZBiXEKlVqnZpHgB
kvtM/xy1nvan/JnEnptPsjYcgss1w9KNDf/v1+BgppxSuy9BzQa07UhKC9qXkkRD
SVjEVEB3nyxJXKLFmpigHgASuuBwZG7uARHDmWtXMLDxwn35uMQmcwuepF6dlDRL
sw/O/DD7HZff1mkXmLaM9alsqe/nYFZ1q00wiTqFkX8/2dZvE6iFqEI/YI3KO/UJ
9qy99MOlPrKlVeqMn9J+RqXvRa0AR2aRjAlLimv7drnHG/JHIBsAxuuhT0r9jDzU
1hmh3cF1eJzrtM7qxyK2UikIG2QVSQ9EHexIVw8/yOKxcZYoa+zQ+3OIhSF5dcsx
lYtzKaKCtd9/1kYPhJWrCcjtyasRclHCyayvyamHGI6O77jRSco9aIrFBXcV4V+h
aMoSu8Gu6KRcCFXXpUg9xxYIs5lMW2Fd+Xfnb6EQ/hS1/Erl9eFahfHt6LDtJLIc
7vvRSuwKlCWGE39WkFArtirX2s5Vadr1EROnr371BtIp509N/gr7MSDdj8eZE42v
RyKWboIPnxtQdtfP+EI7fgEVuXrBC3y1l+eeFo8FjveTWr/E5ShI274Z8MILq2eW
Swb5b0RMndX5Kb7IoJg1MQQT89a66Lr+jBu1ssvOimT3tXe6fPxZqidJZzXLzMOf
v4+wXc2XTqU4SZz488TbNuGU+xWMrUIKY541LaE/DhrVyj9/u7wX+YAepwleZ+eZ
uPXdFhXGUEpd/wgn6kaUVQndP1UiTfoUERtcbp21eLcH/WRwvj1XgvWC4skGO1Wy
B1/haODsDGsHIkzOxBRstW8V6oM6FNwT16FIhM5T46DdjzA7zoCDxfVG8x7XyMos
TVg7lRxk4Mjl7lIq8Yc3Fkj6NVN8f/8mEuPwGN1v3ztPDtY3GRq8tKV35Idnqn55
Ce8CDLKgCBHbSnhZnxmO3uMV0JKy0diIpilrfNTgksB1JqS3gSKmNrEr54n1Y1Jk
ayTwy0/oGu8HhqZWBQAHNLvnzACK0exJST8X+EubjA28Vi0MxfLGjmCBsratiC2C
rqN4zHUl8TPmlnE/b3cGv2BhOYCCZoIUG9Kqpw69Ivkko6j+CmOOxMvlQTJ/+Gn3
cx1oin7Gc8iuFQ8ic5i+apL0j6/aud5+0C1T7mv3+IwqJ68TXOnOmUN/TtfolysT
J1BlGh87VO8B7l8pYOz7DSaEUigpo4nJJOBxIpjQemfHCPCEvFeKYeBI2lppppd9
aPu9OiJzi6HNlWG0+jzgz/LAN2quhKKnj8kzwm4Z0QF5VeXG5d14/dXRBChNREdA
Z65lp/v8zgxSAgqvFR+RaG3Rpn9YA8tEY9DTgaCCsqtyf0ALq90y1hbTLvUlrLNR
1f/cR8quXQzQc3KIudxcgrCacrpbCy/S6VmZPZ1fkPS25FbeNfLzaHe8+7dor8L6
OwUxvHTG9VMDcQnoYOLVcrajKhwiYdeFu7OhJ2U1QcyD2lKrrf5QYB1aijt84lZ/
bCIIPP6ypIOxt83vyIa9n1BXCvWt3kWk29lTX2HhrkAgUoEKcAT6s6G8ssmCKBEn
BIiYz1nFr9VnyS1FRdSOXCZHujur/w6FvpwroSMQdpHzO7MYo+fXWxGeOWREA5C7
QXKDecBFnNlCge9AJwGIE0bSOcC864NEVkuZ9fi3VICR4VJOrDTHoPaYiODIv3HD
L4Mn1CWyqrCOyRv6GUVYTS1rxyL+pDc76Ll4cmkuMYzcCqYrnXZs4MbV4Rc1FEYd
u3hS7V9YypFdcdxxALkDm96FSjigbQkTVrHrpp2iZufZi7UBrxUYP55sq7MAl8BB
CFX4BZ78PUeSQfHi8Dv1NdTE05shYVnWREEkkxbb3EhLkF59Wp8saZWALq6Fq91D
yv2qPVLCk+PWVjFG/aw9DcEv/g8mZGf5JIJb+55PsKi6fJIeg2r749Xsb35pWYjS
BRtJemgCq/u6f5dffQ+wBDbTD6gOvCDSPnp2R2nKNA3qAcyTOApYvd8OKvAwTL3W
lCOOdgFf5QKH12QlAdHLT/ZBJcagV9ofdGax/b0R2uBUQrY/4ODv3eT9Fo7B7hhy
U3AqpwqG39QBdgGg3S43f5MN1iiC/kqybQTSBh8zJcBuQVu+MComPIov+5iC17ac
ybB5Xzqowx/ov7ZTDrdMsjGFJ1Y7/c5pJP66s/0sORxGoMhc02rbx2UEVxBjA9Hu
DJvazh6SMjvJRFhlCDxlLTnoHAzPK3gJ5qwEgfRPJxHAwwAfBMUhi3ty7imXE7yz
gyrpwPeQxyFxYF6A/9eqIfM8ekQcRWZesUMiO4xY0XJGPkPrxYO91pflhIJTsaHs
tompSoJ8JzoXweBbTCPetpX7mKaAAH9vU+xkiXpOX8XrvrCweek9MtUM4z/McRVr
ap+AVlFAGCdb45oi1ajDyCCA1FaMWIiLtBKXVQmYwzXgg62LqUes6ga+RmrajiAL
rJ/0LoCGgneZzKIku5OLl3He3GyVvoYiYb9QX8DfGLPIioU+tINH445taqn0A4Fx
LQSua2q7Nf/6WfzJeVrnpI7x118LkKgw5/gFoSOXz8QW8iQSG7WB/LAoR8QrN82f
KWdCZD8tgBlDsLSBFAAoe/BUfZuBevCUv4llZ5C2HkBe/evc5LVSPyX5WGe0Ab+F
QUnPtXsdXrqK8eYBIdTGLHRp9P3TcPw81i9h4GdGAADuU5Nym0t96E/Ath/UYlqs
z8ImQJmB/5NZABWLw15jSkjbX+h9T4g2oAOguHzPxla+bEJ4umWA7eKc6FpddX3W
ZFwiF/55Ky4TqSSkvXskweb3HUuWjt00l6I5dUI5lCBdVkg9G5qGlRzV4nLIxUzl
NDlEmZ7sqQIrsD7ozK7cdG3hZT0DjudyHJ73qGAVk/UBkVBTpWtf5soM+3eO1l7r
9zGBfWt3jVtGG5USweVGtJo6MQdDv6/76heQVFuq1zWx7qI4YJa800bz3DW+akLu
c1EWX5EjLml7ct5pud6V0a/Jx2OFZo/cEPvRW7Gpypj65Vc5DkvZ4pWf0dB1Xxld
RLK1kkmVgXjMpnewF2dO94wDm28oY8tJDCCtWWeNwskg6jS5Zt2mAd7z0YwO9b3B
whd800dd7KmWTzcwcObsFaD/NOOV4BVeIDsJiIJCTn5LtLzzPZP74eeJJkic68fn
vt9iUvRlBuGaiU7EH3Q82fiP7nMBeXzmaWdWfTzZA97Xf7KFQCb23By8X4/dH8nh
lRdFzf8WMJcks7lkZLoQVzQ5DMp22J94yIEU98Sf86Pc46vlgRbgUywJmJAOQgFp
Nz3MEMfGC2aMsSdUPnrFp6KiNxuSYweejMG+oU5fws17DspjZ6JHkP6xPTBHP17X
ty052D5nO9+h/DbT/V6eQ1R/+Vcje6pB3oMjaON6UbTkjIh3JZAprH1CvYP4SvdX
SoYHaf3xNzDA1GnbAhEBgWRGXXc9mJoC3kPBQxUeetuFPB4Gg12O9EYyKjXJ9mRk
cI86RCiHRYg1/Cm7pvnYon/ktWSxPmTtOtxXHVcs5qQ9YF2uiawUNDPgLba0JXJ3
Ke5ma1RmXzcBLxSRyzdLtyD0RH+qSv7FlxWX592vWnazp6309DXyj8ti4qyFCHv3
KcNDLSDnfpFNSN68dDx3vO87cixd6i0RDGE6e/N7pUPExNkJc9PyhD9lf5FS/IQL
Ih8QZCcF99GOG4JNOZ7w7WNAuqkgEGgqkWoe0Nv0GooCjz1sDLq/cNUAg8/YDAHQ
9sbYnz8yRCbBKRudT+P6ckCHOZaCr1lIiSs7bfjnpI632QCWmS8M0VP19Oh7A484
CqrrlsaKZV11ysedCFRhNI8IjvNEfUCx6nHTugp51fbqwp5DE9WOoohoFGQiGqQD
9m3zRlIYhUo0ubAXjTmh43ifsckwBuRES9GCFx3E820XgonIPWxrRWBukAMWvaBf
nFWLI/Mk+2MIJwCvZh+Dn0ycdkus7E4Y2Sdxo3RrgbmyBFGphdIW85OOrJYXqIq7
hW2Y4AT7u+dSj/Xb4u5WiR8DxIGvfiWZ/1kns1wk5P+KjD7pKYYDTmXNDxIV3msz
OwWosdmJTt+bMQhC2CMad6AqeJdre/8yYOdipp0FS9vdlMrBkwztrQu49WQFpBSK
nOAFR1sXL27m6SMTb7sGg3wAeLnrRRbupuKNX6FIQjUWjO6fOZPUNeB4UlIecMoQ
jtZ6nA0TSc3duwp3XC2VX1JQ8K23uPimfj4/ERlRK9EHCJOvAI/gqMHCUS6ChOQq
v/NSsSKR1zafFHVexfBoCQ9CnLn3uVTXdB5Ho66XkWOBOm3NgoS9mqMtuVYfUfH/
DwXdebMZTy0R8S6YHZqDd80LGnmsRHjM6zAaN1yl05QNOPkP2aP4VgET1D/rER11
oxkmv7Wrzp5UtLTL7CiQb+fEqv+exuX0J1sOFUrUI+z3Au4DjZzcx0LaYTh+9aqk
8/FtEdiZyTUgMMEIMTt9HA/JC9Vc6or4cWZgQPg5DBshXBxgq1ikcVa2SNmAIsie
pgc9XQQWiZT5RW1jKhJk38p1YI+Px5Y4SG1VOXwQIfogfztrSZ6XLl90ynV+4NIZ
0QlxV/i3RuIiau7P3A4UrDFUoqwBMP4nzUg3Ba7OnfMl6+j0FXd1Yw3mQiHJRDgB
BnLsVyeoPj5WReObCd36ush6TOlPdNvXwoZKXzexeBZQ0Br9FRBgeq4ohC89yKlq
GuQEQFERVrfJEd7IPaSTUd1+91SEhK691M6ywWnEGRbG/ykJHrBrr1MCLjOrB7v9
PnrHplp6CTZT+38KKMDG8/4X26WeiE9nuZTEUqlVUPDfcGrxKFQWWbn+IDA1foOC
kKLhutEeqNOZELGceH32tAy8i7I6OQ4bOSAbKPpMUnhKkdxdTS5b9u92K6ujI8HZ
n0CxgcKh5AQBPK5DDvFjGPNG86IA3KkNs4y58cyocuCGAxEJpDSp3N3caA+CvbP7
D/EfkT0MovQtYSYyxi4vK3mUY09hBabsww7Vja1PYzjgCmqZeoeer8UqxlhGqouL
38WhTc3OS8eYPIv1feTVWoO+pZczb8LDbLeY1QoKQEHQ6Y8iGhVBk89k7ceco25j
XBJHWfmzOVfhIqFWwKjk2KSMHCIp7A6DttZCXCZfCsfjqcvtY9at6nEx1z6/766k
HJiJ0BtNjL4wq/pP0ByDO1nGLuJU+ogafa9Y7zKJ85zbGQDKCXXQM//cHM6sPk1v
N8Ginz+XxBV1rCxn7qDldJNrAkLVXjFKdm6/uFCp721VMc3MuoNUarnjajIuCZXf
iH5mu3BXTXpmh5LbOf8JguOyQJvO6Gp3yYTpFIF+PjE37DNJEGfNod7q1ESyZnyg
RuDxP3vRZhiawrXsqGfO13CPXYdEQjC28ObCD7KUVSw7fSozOxkM0rSfghey5UY1
ZkUcAHqMN7+2+dN7AD02/zH4dBsTGwKVVXaDevZsfhaRq1bZQCiQxdAS73rqE5o1
u+PFaVlf+FsNxTF0h22zAbGJAAtWEdOEIoT3h6oRUltmcNhFKJwmKzNM+hggMS0x
XTE9S55gDtNlY7nnpe8gWOdy64XVOn1HaDCQWdpViWboDLmrTDRXX7LbVbvoZoKH
UesAnVlqjHuvm5p0Ez7Ec/ZB/DSUxyX7C/gPPLYyhzigIUp+bldXorLz9ddRfZ6p
g2z9TUtkyx1VQ741KAbrHAl9/HQ5k1mWzXQwTwlU9lBJUNCAAW7exoia5YHcLDkJ
z6Xg2c607rUUC+zooFc/X11myxTVqRhnWImwS6OQKHyWTdl5ypjKhywUs+a9SgB2
loj1YBNxT+TaFz+k3eSggW7BJFj0vK8air86Nx71Lem4wuW7StaU+l9Jo1ElvJBZ
q6nmllgsuyBN1iNkAH8avUOJ80w/qyWzWarEksk29phGfNc1tPyb2FGPOjEwb2fh
7kXy5dVkfd9uArztT+quq7c9f0eY3zAMwO8cZlahRXukuHHVa8vF57ArUku/1Rfw
/EhwWQcwl4/ogv4A/ns5Va7+R3MmZpxqWN6GhiA/EI/1vBTZGs3eth7hIWV2rRYU
3ReVn/ql1mytMSSzs5xXOv6iJRFwbGvwkZ6A68TrFuUf7/BvlzduSfbIdMK5v/j+
m9jLPjrWy5PLDfOmoXwNqEkvt6DdTw0o+ciMtJS75HxHbC+Pu37BnzboJnpjikDh
Zjy4s/bZU6lrpWk6YZemBut8bcfaflWLfaHx2hggMHOYRDPahkbHW8BvqIHpkn5Q
1svVZvwqvFdKF18eRbYfm/hyRaTrPyhb1XpO0dKEewjEBe9EUgemBo19UdNoTWQQ
uc02tQIUOF2MDyPybfIK0p8paY0pR7cj+za2vu1I1Z3yL9Pi6GM5EchJ8POoLQ7M
gjzeu0PKiNQVmtdUSg9sH8l5ZJjxHZQ/tD1yObTPJ/ksdePPoIdr6eT3mE9ofmQV
I4KQ85l5Un9UOlnaKQRyETywrb/ea12hsZLQj+VEbxlDg3e+h3nfs7fJG1cr9iRU
jheUmms3wgQpIl4diSJKjvfBgqN+wg0hXHlwkHYS7EJycYCDoGAH5t3wiPkqrLeM
OKvlhKYq6USNrbg5ZP3S/wA7BbSQAfqk91Qloa7sSuFYsN4/PkGnFP0Qothrh5X5
0BRHHgx3/6ZCZVL1bZ1KltS3F2XFi4mcGETwnRo5znCJ2owgFEDLJm6sF2HGp3Ek
xGdKqE/3l1buor9ezg3B+dbS8PcoUrA39Qx/b9PVKOAxmcE0eQqcg3q5YzQOsAxn
YUx6P4nvZsvcaXMyP4AdQ+LgeuHyEsNkEZkeUThySEBwB5+R7aF1M18qK1sTJYks
g4g1ix/keSBSBZOWfkqJsSMAyYGh5D+2K2o//TVLg/PqvgryhFseWWh6xJ8vzvnb
7gcD5dCSBXir1W++j+rfa9PQvQIVTPECtvesguJEJrtl+Y7KdUM/4ktjZGnIgvfb
HXNQO/rpt6FZzjLHahFPnYcUtqutCC82FsuhpgzoDnX1DZcMYL4mDOoneuhYrLJ7
Eoq7976XlX/+AhmpGS7c9Y8ebPS7ub9NZaCwhlA69H+pyGTIaLoxeqppqIR2m16D
JbB0ZK4rCnfurf1hABO94fUmIeSMKCcTarnxuOkQU9TAQPrEypgzWw7vOp0r6IgS
hHues2rSGwDh1rOinyj4aDsgu5OXFW/AKwq2i7jij7y4X72tatoAmmP0dgwz3lSP
6PUNaMzw2IwITggS1Z8u6tXVEIXZdDWPzpXlK7D5ctwKmzjFjiWUHCeKiMHrhlIw
QCHTvH13cU2nqusJujpnUG3FrrqS9/Y12qwsP5wUrSpmSIJiul1EPOpQBE6Jokpv
pB6n8IbwteBCCfxJDhhHB2XdJnuODnmWggZxTENHmm7dxwj0+uh35gMv3O0x8wC5
W8IMo4CBKl9ybl6GfikkA3yWrPALODjjXbrh44mvJzccYZcRFA4cjricvXJLtWyy
F3qN9J4XHuEhi30HYyY+004o14f9zEozilnwuK4ohOhSq2Vl0I/Ib2ns3JXHGlOz
SWH9eNjy7w0uTZm9yDvtj/1x+43vh4AJ+eOQs4+7plzRwn3Ns9v8vvYRhDrU/SjW
rgzvQDTSKLrdFcbTg8sZEXGFEIrizu+OOcldqM2mrxlrnjYcJbAqm/fOI9qgFaq0
6rbokj6XLZYoPWtZLlvUdZDV5zpeVWexTe8D0c6V9EbzenUYPumpFCkloijkmlEA
FI1nenvrqhh50qC7fd9/XY63GLCL9VGnB/HFuuJZB6N+WeJFOV7tHgzuhGpomIaA
DtjbxDYxAlw9NDNL7yV5A4ekExngqbP+1ZIlSzD89WPWV7ZRF92suyhbtF2vNW55
qCLikm6JvWLRvwywbeq+u9UMczksvLOVG1+OtTYkGUMrUa+jqnJqzLB6Fi9d+Sth
bC0A9Sj9IH6rtnkMPFMv/VDAlBXwpZh0BJ7YyH/Otq0kLRd0WJmjuTHHLvhxEues
Zh9R4javQIA9nUTCf1YGOaYkHBaV8gTGj9ktW6W2h0oralpoI89aWGme3QtkvtZg
iv3DJNUadXpISAKcPSTHSe/CaHFq4H3UqWgyTfFof0rQ8cBaPnOeXVGx6+Q9neXi
5w8gQMOPUgwsMW1+/uVt26UmzQ/f7VZM+3t5RRbg3dFTITQUr0v9lF8QvvhXXuGb
Vml+3omRxA3mQzqE2BaG/SB8cyjjiog464KgJrXhTA/lqGPyzNwlTA+XjbIUzYlT
/EIrD/P/yNt+JENZpcJe00xK+1JSjzMUyFPFoociGNQiSRzzNVtTfALOPL2dwqTz
uMXZj0azSnNuqE1frZKtMrYeQmthQR40383HbeUI6Nbt1dJvNSv80kD91dPFs+z+
InlW9+Gx/nK3YeADXkNMT7StytWAXxxQsytFNOjt1b82uv1MH9ewN5M04XcxgPfF
TWs85h0tWyXpoV5uXYsrsJHNknM2CgpesX57mYP6cdPhtnJVHoshsEd3Xlm4Jnq6
JTFTOGF6OTWYAGA+ADaqPyaZjYqM6p7P5CimO7bor9L90OUBUi8j8yESYpYeoqEd
A1lVhx6XJtd6sZnfXHgkhi9UiRnctC2jSvVMLZJx/GWppT8EzgmkheZpReFXE1y9
jaEPx47jBOvdDPt2MkcQmngCicsjlEQYDS2oDx9dGi0h+IKyYWWBTqLxwPWrcQhz
eTcqaIe9o54o2iOgoQvcv92+nMsRJ+kEWUXqbxEvSKolxWx1L0gYcAbALxZ4zrWU
lZRhIhuvK0BtsjVqeE8ZY5t+sPneRPvxk9bmT9Z/ZovwD1p/U3XUVzUHdmpdSFxJ
O1BXeVt+4ezOo7y12ACReM6KAe4Ryz80f9d8WCRQer5ZHNrVe48cv3zpT0HmW75x
75nXyzRRytuwPUTR2Nwe5q34DfzJTrBBBoWqoifYeHomMskJZ25ZkW17cm+Z+qF9
csdhh702o7jcvz5Ap7PMYAfkfq+t3jbywBaV9GGxpB4EtM554i30W4QqmtaJSWB2
i2UqEiw61nYF425kTOafXxZa1hUxFBGxcOkmVoYJqf1RnfJaFQJRej2NeAa0dyZD
bq/N6oeXKcF5P9SJl9CPoQ2nozlGQIlMIOE651+4l2EGWXOf+vyel4Ov1LyE+3xU
Z4ICv+e9gfWH+p4Tblo3A721aUaB6VQcJAS5DMjV3otNuVOGTuBP7BY9swzGGs6x
D/Hyzg9V5EtVrVUrDlL47B1M3/h1URX70UOhj5HL3DIdqPxUp8oAT0VCcM9UOnlT
ycfKAxnXALxg+mPvzUdG5zQI0Yv1k5oDcaZ0TXe+AXAwcbR0X4Q38HUB72+JDVmD
wPy5+PeGehPUimiESDB0ImKTwfz+Sj/WpV1BysTGyywt4hZBIlGPgRRQ1r9wWqCc
DHTRKCuK1LAScugwngM4zBdDF3/lBtP/adtmWnrYHtgl+dNdRV6fyJ3y3lUpP007
syYyB9SnHWsFz5+im2wtm7eFxrG4Nk+YcfHn4EN/wFb4QE4SywPiXn8rwQDm5zOX
M43yQhP9CPOlZi5WdL4ju1tQqd4V2q8I1pB+gWYvdWVpwu1b6O2n6gvGiR0vbz0p
KnIt2UaG9c+pWuIvNHkqsn8HkrW7F8OA3mIK4dbdND3b5p5cgmd4Cj9kofpErEL6
/g9/V5GKWCH0wwkKu7J7ZtZveGAj9tylap5l0kabXMSp/nlOlEfxq2zcVJektRWM
2NlfhHraR3P+L2qOM1/xxt3sdbSYBXrWapvPmnntKLBY5zTQoJIfsZX+rchH7I9Q
B/tbhqbqfwbZ11lQKE9F42XViTKGeHk+b+/3HPHi1w77Rb1M7DHcWED+eRnSKffA
9s/1GIbWGkv173cowOpdzXNX0SoSQrGZCu8o0Sety6SWmRxYqN5UoZGTnIhA8Fx6
Fltasybh7fTAZcAHuH4ePbjvHBy39RVwePlIPYYvUq/6nxnH2b5LiHCv2YbMLhC0
Am3+nIMlnNYGY4sjZj7iRlPjUyrlI36BNBaeAPVhC71gxVokXfpD8/+Cyvv4x6+S
s2jS1NEGk3Zn72+jr7MJGwATd1J10pKZ8dpnstHIkhtoWHrwGjCvYj5qlR27pi+o
KU8tyBR97KSjQO2kfKX+ZX1A0CbHNWpSA7akuQm7JLbnNCALBeMrBp3mQxk+KTqt
Hznus60Mw/aolHnbMr+jRBFpBXGONArstPeZKO12pWHNHx5+i7iRW38Qr9Q2O9bo
3FRsN+ARCEVeHS7+7Py/4Wa1nfylDOl+Vrrw6rH0gqyc1eVTxNEos9kto+pgoZGU
7+M8A1mlg8LzsNkTLp2PdF+SXQpMa1wxt9OrZtX1xVH34S1CBAroS8aOaOVjKZMW
rQgmue6wlS7OuiswduyJ7huSlsziIof35jhkFucxr4iMRjsOejG4L7YimKoYvJNS
gh7HujZH3PBrJNwMEHU4R9YpTp/m6BmLMbHV/dFLpcoDhm+PiNzBx4GbaAa0ZuH6
5whZsEwia+gDX/X0eVL+HeRx5oFNHv44Hl0O90OnU1Tuzchd71Mn+cWQHvS7rSPz
l6Igy/Y+7P1D9YxWn/4z2WDC+Wt/Q8KeRF/Ikdf1JpCl2x2iNG82aZe8L/6cMssi
U6tQix1Zx04Qkw2bWYq96PNw8X+ybUNeatw5xPS9yu26YtJwtoxFQhG0UgyUKGSH
/3znpCRJMKWnFAHV5/AJQcen8b1eIOcDZYcp0TsWCCr5DxgFZ2gv6keHdimcfVz5
RoCY3IRw1QBiSBYyQnla78OnewvefYU7J/kPIyqAN9+0OwGF/nEYvuaDVI5/u31y
vDk2z8ViqPorqi0qxX5l8PezNgNPXBWybq59A/zcqbaPj4hFjPCscTBN6JMSbb6D
VyRp6NfPT005mpMEPuaM73SDM3bcnJj3JEN6gYSlJH6kOSxnskyZGxZME+zBHnGW
VaHxFs0PlvwdJcfkuRo3tTe3xW7hx974n5ipeUjvmzaQSHclpM/rpIJYMelTZPNL
5FhtBIz9azqEVIf7AXx+Nt+9ljuT0FhXj2LAFV88pOxuyn6lsYA1cXu5BI2Ra9UP
+7lZiqOBlqGik9eIbJSHRQosM//m01pVFFlrSghRk1b+a7j7g9rzGBTJ8K3x3xAw
KzgGxDYNBDmykHrKiJrLmEmZRVTQKYkgjODFLJ8SvDitFQtyjucGwWuJilnN0VeK
UPqRvd+6CjfBqVK86pHToLZICmEsjbwNYbBexrIdeDJy/d8EZEeHP/z1NZ4XTuZi
38UK7HH8EGs661NTxuZKGK8J7zMLIqFVerDBZXeMUbM20+8YUUqR3LgvuBqM9dRf
T0xBgHpzscjaTlzohLACY6iTDzFxTPupIYE7sVZO0iuYuiBtJLwvpt39ieV9STxx
W8OfO/x1J1pRwuytqHDTI9CwxcnQ/soEot/jiC8KajnZUD0o/TpLJ1GBwdKX4x23
LHUO7s2mGTsd2k4dyjqcKHBA90XCLInTfyaHcWjgn7Bn1BzfxX/KAsdWb06PJRC9
hkjj34gt/fjkZ0ePg0RM+fTMW0fSVfUlKC6IRZq6bzeVxRbfYMVxmWI8b7Tx04yP
f/q67Z6o3Uc6qadBzeSrct0bAL9q5ZoOxQdXAp/++Z51kZz5WQhpVYRFkhf6PHOS
u2rDLTZ02lB3mHv/sRdmzL2JAH7wt72KclgrXscTIr5+Hru6ikEbRcXH3SbjKxkD
gc15FDB1rrauxMw+cr4yiTrxESFK/lKOLMIoX90TC5mWdf5tON7QKoLByQkCb75u
IINL/z7pdIHU+H18wtiYirP5pjnZ/BrzUhwFaO9qXGHF8yU79T74wxd0C5tHGe0q
YyGqdxZcLr/H9fi0eEUm52x4+rhtboEQeNT4zD+4QTYCCfyvOjUt+yxsAD0nj0Gx
IpM3qFmmjja9AZrLAcoUY5VFXevoD+KrOPQd7dIeI/h+o2hbz1M6TaYtiHCjBBCu
vnc4IWFQrT9mEe21ZlAeujmqsAWoUMX0pquOeyCaUq+nf2sT5DgT/709HE2hNwhH
ImbhvePDlSdCj2cm12LevAuLW5eDXiUMZxBbBZp1LLCfWv6eH8rvE85tZWws6cRq
QR4XlAWSaYwmLHAGhPl17htu+mAW63gCh7eqTUF5aMQj14h6bJlMH1gvqc/jaNMr
da9vXelbiDx1XgIrPYGzkr67r3ikFDWvDZQ0rn2Jfyyo93HmNVmm/36WwqE+ltZF
5M5Zu+72jNB4NG+CZnA76xIN7zDN8uUaUf+NTei9miW4KZjA5lYzNlzxaXFS5oaF
9pCsBuTBIu5cP6Oiy0nSxxRDF2rRwm9IAoFefW7S+Hq/+FgZjMnBFHVGUBvJbCn/
pd17E7dUwmSI5FOUle5QpY2PRqBiaZ4AoKurFCcMuv3Fy9hU6b1Bfb46IcjxUSTT
sObmO6UilIDEBmi19xtKrr0MQ4NlxfEdYenQyIfSLe6Hdh5MBiTeDUJ9w9UBpAUl
bGz1wf0Zqmxwh0sLNm1dwKNWQAW2xpxMcAhntnL+R9lqT39D60JLCFqrZHdKFLdi
SZ6NHD3zmJ/X7hRKfYMgXkNs4BRmb+dNzo588PvYuzv7WAjDbsvVJIii30cQgl4o
c043rVjvlekyLsernoA9YpayKTJSf8yhREwAlaPG6p1v4etAvnNXCp3toby/EjNb
hSrBwY2uPa3EZzx1XxDe/XpRD0GwVCXiTwkh9QGjqD184ii9NEVM7KEVZCAtghHC
r8hsEEhTbSSRwVpQnNhc+hifvOLJRNUQBizKAtR9zSiSK/BKp8OABvnQYFNC1APv
QrOQIF69f8z+DoPNhxhDW7Lre1TSZjbCT9l5SIXZkJTeuSx3o71xvJduFjHIvbCl
AGzL+h53mSEaR1GN+72gK7TLajjCIELx0wqtJqoxRO2eITGVJ9ISLDJ9sv3CJeeg
tpH/t3SRMVWLI40ccyGlpyevZXdfYKQeyPK05Q1WkwPisUUjzHHbcaKtwYshcPag
2EmWNgIGqIALLetUmj9FrR/U5/rzfw8qbT+KHCoojQL3zPtU4Mbe0zNHyQZODquU
qI3WECwtEHq8rZdgTBsPVAyPDA5PNiu/IesIsj/ARF0yr9LyzseE09I4b8B1IYjC
ry+GYOAcfLRy6pyP8GREAqKv4ikCJRf2VZtxDY1Du//Mw0iiQh0heP9n2kzkgdc7
1Kub0uZmZO2LOXRbGwL5egFo9oUcNp0ZmYzxnJHTxsVx/njfqP+cwFLkMG1X2vUM
TPHBIZ4HS5V26DocHTfWrfGYXeO5on5BQ+zxg3AEBOZ/8clWGyJJV2NmWVDBCTAi
XMkXCYd9bt1QQ9LUxM+iUB83ULELYduGiX9GWzrUx9GIIKnRu+ZjrXuGEZxvz6lb
LRjrpLl1e6rOr9FZvWlGfq1eYbW+1TbmF71oYB3Mm95appgH2Z/KKackpkugoR9x
k/wtd0qYUR9QcAwH2sbTmKecf+hk9eIroO9CubNrmAjyYs2kWRYBThYoTHFF/XZM
wUoFUTa0zlsyw7T/SaR1ARP+Tvd0rwyQrDAxX2ZZJdWUDUrg5hwDaI4y9raelDEu
tmf4Aj7MguKOYJBwL9XnLO8CdMYAgSD3WZ27gVCjsiZB/+MZHHIF0USxLnu313yB
hGH+1PEePUzxgaLbWNklT+pX1h3HJ87e9zcx/FiNQs1Q1kpZIXPo6/nIHNze8Qwo
ouYnfPsDuPOI/jav7swOq2GQmrgb5PypGPWGozKw6KI2z+Iy/WIdFfX4+AEqJpwb
sSQHFHILxhDYguBlvTDWkAU2m7Gazqjh7VGfWeroqp7V/Nidz6a4viQbM9W5fYa1
9z2ioHBgwooyxZVDbENgATBD7TmxEqJl9+/YSc5AJEF3N2AiUHwuXW8qGBysPpAF
6/9REDgQPYcj0tloNU7wbdgGDxSTrD5L0/CaXrjFejLR0Ijydf2UgEPFUxILUjVV
0569Wbdq/X5bgm8F8sVfcupqeUSjJO1moZgyNaiPfQJdyaqV63gAuE7Ykp355Px5
/9RD3oxmIFexFBV1SxEPl9VFHwU9CnqIjbNzhndzTGRy2rPVamnP2f9DTrMwEmNT
YPGx4VqLWcgzM9/FUa8lUDAIhhbAT/Zjqkuun3BHbBHjRH8770uRHANiEgN88CA9
C7318hNgXYBPvhY/n57a+eUVl9ZzbO98E/fJLuufQTenu/Et+kaDxQ8VZQNKb9aI
v+xhSGV74GdvKppIy87A96zA20A85KnigYfTSCwRwxO79E1XheZXVmk70BImSeG2
vulLZnq0rAM9/Mwu5JR9Dmwa/e+/X9Hy34zwvjFzD0b5rt0A+/h3BjYAtfTzJ15W
xaoluVv1B5r1Cs0yuXJW4mxPUFoBXn/lkB8Gl5XqLkfg+BD3ZprZuT8eI70DYZdd
PViI8wQbQuD/HkHIQakg6K7yUfaf+fqgvzioMLnQlp0loMWOfMwOdj/7eYoQ7D5U
kz5FYhEUEe26dphsHrFmIHliFEYO6+fPuRhLUYLH3ihwFfkJq/HdAJNlLDBNd5YT
YIlLlNXzrqnstX5XvGVv56YynI6TWH5BEWIJCBr09mbqimLiQIaCrGkdWDEHgxY9
3kPpKOVku4ASJz+AiyQgb7/wfcNLOIYZdK5fvAKolRHvdxGLTuk9vFnw3zu53HrI
3kmRw8NrNWl5rBhSmzzmgkMCMLZd8SCD8t1ENAJFQVeBgfjKuwvA/Samno3nB4mb
yL9PiVYSa/Bjl8RSrBz6xyW2BkN7uLGrVUS5B7m2xoHNYBkHBH9w9XCbCBGwyMd4
nDAY79eDLt0tbaAJ2saPcQ22SX2KUaKpkuXX0kS0BXtv5D8ixqxJJX9xPd9HnHoZ
8Z6k/2xQn+5i+gY9VF0dmpW3tmOFreeGomsl+4i7tZqMNYlOfGNShvPIhla9L1m3
q1w4zXTR+wHDtHNgpDsC0aGNpWpeRaWOtDLzuuVPWd1P3M36Cc+Ft1rl7DaczvGC
rZMrtUQGIc48ceBXWFUKN0r0aZOMKqvRMT/jVtLjhti6U0SlRtQbYcCNQGTr1T7M
qu6BnT50XTprryFdjz8nLCffxmgLOUauoWEpHLRLAHgQP76Sg04auksrrW64SUXh
AOKVWFSe8s3UQ4c1/M6CXYjr5s4z6Zhrr1TlA5ekmspNrNPj8UXEStmMG9xmJc+c
Nt8yRK/TTjDhd3SZnP4UOZWsMctEEzQn/eSvrZ2ASgPUdSUGJL6MAQL/K6Vv/EeG
Az99imF5TzpiXS+2YjVNpBvWaMJRzVJYRqhfkiaXke8DN7PmBBvAsP6p4c9rSIXM
r0dmH66TerqUOJtzBFj1aa22hDu+VhabSGoxNz5prQO2f4kMSKc7xWECRCT8n54M
k34+oDUuYx/waNCJtL6Fs4d0gzRUSPX5017Z1WF2H8fji3NpbT5IteZrmLxxIq5+
ha0XK9bAEa3uiHjXaBSAXwf1UpTIzhmi2QmpN8kZaiyPjKdzvCeyZSDu+rQquzhB
LUq7hqxRx3tEp7S+EhxifXjy+sSMwo25HDuUjBrc8QJoC2sOGFwdfnGQPr50mqyv
OXnOsN7859TK6SCKNNHBE8SDnT/v0sBSSxKzU3GLjFAjJ2WQ1S9oiBrbHFJg1GV4
Tois8jQFGIUrp2TIh8o6tkkskb8OYrSCpkwdful7udRvbfPIJXYnl9tAM6zyP5DH
hjkm81huZ8pqQchzAu+C+4x02bTPdSTAPDAa+rK+7wYr8h6ayAlZLobLVBL2ruzs
5uSdiBEWSfPUvkkdSxElcqG5kvyU+m4l2r9iyG2dHtjZ0ZVjC4i6E94WnWnuAY4t
xbOw1wnn1pxobiD1tA8E0TXCsMBaEerPg4NgKvAenEGI9plRm3uzC0vw68twkavS
xRGYhHM0+TsMSCTBinMLJJqW0Aidt2DQGC4LHPGkf1tHtxXB8DJOV2f+/PdKq7Ng
ozjtkKMtG26BiJVqss0CacrzNt8DjIw+ZX1hSL52l/TDFurp3feWI3dfxKNI1BZz
lgqXownEG3G8pw8R8TrxkYz+dQo6D6bZXbub/MJfWJkrPVFvmblA63hUUMrQjXRz
8wJYYScRnomS+m/GVxjOn7tah3kZMMsWQXXeWQJrCIVQ7rjxVlTX6webDwOTlTqC
FRX3PmhFDzd2eqCd+yCfMgDMI7wHFC21eHh8FRsguSj3Dm1X+lFDEne/RGFJxxM3
nHo8sEB1kv4jgnGyTeLv8JpRHGM/wxfihtkt5OKgHxy8aU9vSHlm/+lTqXdRVFLn
XaFRYF6qqwpImUDD9UclLWEdGczsUHJ+GDF1JVXXYahDP+V4R2F5K/Jcw+7RK4kP
egmhLBZORU1rs1YKYU9bH0gYAVdAyVzxRNV0yg/YYBCwlxDVCoKU9Lm25z3/yykK
uYssOc8yC6Sv7mHEIXR8cmkd1PjGmz1mNhjEzlbwBZeKf0PcSEF/8Fz30Mx43GcM
2oJEAoV8yfb1mWp/o9BILw9BTxTnrwbaoCmOnAOyMHDyg0jbvK6HATD1fG/mROLF
xVQ6z283c7wKUXFP9YB7OsgEC5JfqL6ZeX1LU8DAteTZNCW46ab9IeApxAf/Rz1g
4RqzcMXCoM0pxivnhFd9TEgS/MPDKQlVbZB68sttqxvq19tKHkykaQzRmKPGbFPb
FD3W3gRN6zuhQBlbP04GLs5yt1/3Cnf2BIekb5BsFx8g9ZsltLVmrGyBMMlbj7Gx
aaTBmfJxTMWiQqnWyFXLv6U9FFaz7+W8rsFh1DVpeyXZF3pSv9fhlVTB6CwnHD6z
HGbqF2cd502pd9Q2x5C+TIMZw4PT0KvqiJAs8e05A2SyLIFiNjEW4EWiM7AlmMGc
3mTbOUbLk1/D6k6kmTR0v4crayj1+NxoeM32Ujub5Fji3FKcBaxhetqoVlNCSgMG
qfbtoLW1KrJZmALMwPoqWxd/jahBcBoj+Ikjk3vpRQ62y94bVu9fq4vCFThu6EqA
FSlYhGIELENvX/oAl3b6H0Smg9+HmZAWXONmBLHdiPErSA3MbadAQAEAqGZe4eC3
Ypt4u495bQMBYXIeIE+YLD1gSZp5QUMzNLZk0KK2ZRkKWd2QFsM0ZpUjQKbzwZUp
J9lWpLwI3CN7zwwvoBr9xJm0abAeTauinVa3vVggKopW7a7zBr7IdUD/azChiqz3
wsAiNc6qZzeaZ9tyss0vJPXWjQHI7pTObPmwbiSScy9mVr+ziItpXrQcdGzBI/7M
9MpzM4qsobpE1xULXQRIyWKuIpBmcJ3ddmDYymj9k5G3cUM2ApTd0YJ/wKqOXdXz
aNeCgqNj7NzlhTZILWbLFiCZpWjYsTwNzNndyWL886lnYpzyHc1QWLXFqHfnppuf
4biYFmAffaS6LEihMjlCYvRUiD+ya1goeKmNLKnovSKKk9n/q1sPvxxuQ5oluFp7
Sfc7tmGnE7T/M+p4gd7BTni2jXEvjIrRNz7DXGnRwP3DLm56W4Rr6r1VpZExnhA6
Brp+Hp2UnuskYWEB5OZHSH88NKyTjg854IHB147fhfGnHMkBMm8AxSsaEFS7kvEc
JnicNWJ7721w/pfeBXeTZ66fmyojPZ9sVm9HAfvBBFkR/2YzyTyTj7NcT3dJQ1+S
Tux2O1K3cJEBCdohKQBuYvqnurwgfZnhbaMaXhEJFQAAugGIjUus8IXc5c6SfzBX
y/5Or1yT5SUkFKxQN2LE+7l/8jUXGGA4Xr2t3vm+/5vDAg1sr1JDXq20pFhkTUjv
e1fR1E6zu87QTkS11CljZqKM21kcT2jWvmilpawgWbaVMQTdJr3NbYhajLH7Pb9E
Sbdr34aV67Big2xjXRzNh1L26TjTxVyAkSRFJtgLmlYa80NP6bfe5Rzj2Hy/TZRZ
zxb75jGK9obzq+K/3bAyoItpWrafVQc/CoSJRRAo46mF+HQ3cVxcS5HBYri9X+p2
J2iy5BL7lmfGe9is26HwC7nyAA9N9VLmUxhL093z9GJm736IEXOiTkZQO/uXN1e7
XwDyxk96hWDhciXXiX1LZNS3ZNRyuWj1UA9oQhTSBVc+jSzlgmQxPHa3fandFp47
7hvveKJ8WUG7EuNt6enBhsHZv2OcYhZL6SQ3YC93GUcQsoBYe/ITLEaAGpKMJOis
0oBdHYvFeP7gW87vKdev9xefKe43GwO2pHhcqfXlyRb2t+GS8ZkcRKIwma7FOVF7
OJz/xxpp3RLVLzsWWDwAQMfQpe0SbDHu7/9OHXywEx9uxy0YvwhYzMB+7HjsPR/Q
VuL4VqfCXHOax5ADgUid1srXB15wIfF5kzbCaqfxoJ5IP4QMGBWiPy0JSyCX2ska
u2WOQKGs9gassh2+K30Ib8LIWmQ5ekLz6qiFBK8LBQkLnPgXrLs6SiI5ixw4K96Z
Sv9OeLa2hjFBmUGOyS0ge534PRuTFVIPdSlmjy8ut8+UHKyoU6LR7KtUtGV00JFn
YlVqgdS7UvnIPn6EVrtKyizkGOoyoqM1H2z/pLCvVqe41OyMpOhwX36HxuiKsf2P
pk4LIYtLRsLfAI5W76V8M96ZEacuQBAfxhNuaKctNITgaXbraFOBU5p8SKSBxtR3
FKcJvjb7DRUPmKbKXwSSTLwMOWKvOSJ0dzMe6J+5JJhv0Lvx1nxUtnt48RPuRozh
lqCMKwI339ys/q9rDzUevr5xOes45gDr5AhWo+KxwvveorEaT0GprdE7HG4tHL04
pAS+1Zk2P3ieWIfKo+dP1OiiNKbn70dCIMX25QM/xm8NMlABYKGxJA7kS3DjaIt5
hZ3H4yT2b00oztvQJEejIiIW3krnzxdlGD5s7+Q7oqujg/GgaDwn+Pec/g4FPyc8
0MHK8eOGHAH8iRZeNbs60tAftllMZeQ7L/6HaWpwlfUEgBl3RKfv4GTUc4kg7XPk
457P57O4VBxyIxH7YdABEFFGs3SAlwMFcwyAoZOYpplX0bm/XMiiTO7qEU4uSt1U
gxAW477pUz7ELi66Trakfr0qgun1gg+2wRKLbeJwJnmRHEfOuHveE0eRSmVj5kdt
tgAXpojQ3Fmb/O6mDXXqAyAH7tkyNSMwsqB1tVNICwpGENqF2DDO8LzpUBPMbQ1z
pnOkDEaS7tKch27qhirtONnRXghXlciismfxDLBRU5bAglcmxEHR5SsxBcjZu43q
KoaUlo8xYzcsKK0DwoGvPP0HkXCGpB4MYx+AvoBBLooEpGkYTx5XawJN1LXx27PL
W/GKYofPz2kNpSs7mI3b3GE3xbUMJu4KkXmZQP9pcf3H9YOn3x17jTh1BRoM9RNQ
zhSqY12g0PCPr4oHk/tDSYiE6eV/Xy6iytmmhTJ3NfGfIaTT45xDlBgKVD7WemmZ
2VyM5hwCnTq5L+7kTU4daxpFz1IXQt5m5oV4/8BXpJbsUNjZqSpFCi3/EdAl2mlB
NxLMk13Qy+yl/+n0o9NzBzyzEvUxJgd5mw/1pYlk5eUTG1mn/t7FpMRKB1THIInW
VJBpethN9O8T5/Xm8XomX3XUWW0PGqJ6xM0G+8GWutT8i64izRyaF+nS+Jw7t5km
j2TivRp+5+qP/TOK9EJZ0kdMEtPIQCjXvBypWYHy6Zc5XAVIYCBMa17NPURqho0f
Iy9HusnFcgVTRJZ30GyDAfIPMVuoRkt3hVSv23dTWKKaI4wijuJFjtu/6q96EEOs
ARIfjAQIg4t5svSx7aH7boi6GaCGJwNM4kSWUozmuX5C3mwJjzRdPssrv4Y5DMGg
27XSbQcZ6VkKwBoqWUEVzTlvMkPX9TzJaVw7/oM4OWdTlnnisAmatHz1zA19602r
EZos3Eiv2xW9TE8LLf3uT9PnGn70qbMF5kpOdCSdqDWG2Ar0yE1ZPeM7HqZPZiA1
NwC4HkwBbb7qlaIELgpj+r9R33CxunJyZmrlMUQh+wKF6EbM92Ft3gkXTJAAGfy7
eyxBKtF29EuEmpSEv2eCn0cYJdEBWrQJ38cT0yd/nDYdCaMyKIoTFZW2Q+34iLXt
J4ZhmXVpR9Tp2tMElCY572J6zlwC55e4c7x4vsKy4OLpjxJ0wLvlQixZ4sFRRAuj
7+7PdI0Oof3ZBuEF5Xup2+UwiFXLSKeJyHfWrM8wfmA4itqTUDlhZD+qg91MPdpC
jJ7jfRo1llsp+JFvIZDkGAV5wBP/vllfzqATxn2acZ6b+LAHDP5JetwvThKhDuva
peluu0DiDRVQ7vtUcsvtTYYJ1AxiWvdDRZPrS5LWmbaRtZhhy1PogHTTyb0jOXz1
2o3g3EBKZHLriQSvKMGjq5fln1APiE/Hf77dO1mAIVFEW13+s7cQoe9SEzqPJ2IZ
kXm9PmKu1iXKZ6oaGE5imOOqufGPNRw64IwOSpC5mYO/n0XQCvUxryriP3sQrpEA
fB87xAwyQJbNk9JTcv0Uwi5P7bLwgRFHmHTZLlfjaeZ4Jg9kdFhHg7Tw2by/ndRD
0/eipjNZtQc0T8RMfUtBkoRHwXcEpHnNoEI821WALTYxwSXTWPqc8cj5mfYVNGCz
L0e4kuR14oHv8uTFtAX8OYQnoMLHxTOeBZtMK/TOeGuc82YoCRyF6hlBvzFUU6iZ
dwtaBDQQjLpX9zIvv5YDK4BTiNdJMEwxMGMOCrAzuQKq7az8sRtkcNNWqPgtcruk
vHK79//zCu7zgV63snypiLMOAOhH7Ux3kLT/CJW4L9+r2ootoTmnXlFIVPtCt5dQ
cm1eJ1y5k3BsbqTwrrb+V/HYRCg1fasXmqby190gt0lkiMOZRE9rp4u4MrWOZpRT
A6D02eVGggdT+0uz6ukfdbfv1be8Bm277oRc1aQk4AKJ8gciIBNj1FyCRa5k2NWP
GI7nccPajWsumXlvu3Nj5WVUviJrTnjoBO7WQOsk92heXx68wpaTOKH6ifTOX37L
XcYCVIMDFAR2Mt4T7okvbM+J8LzY1dz1U+6K+dj8LiX2q1eMuSlZuoU7nJjKnwpa
5K4Gr2kz23hmmeEV/t1oq4t8TWBO65lI0D3nsCXa8bk5+8ke8chMi6YQCiA6u65X
V8yQ39q9h785cDq8wIekkX+Qat0hG8lkRDZFW6AF0Ve5lxBBdUu3iTnKbm7IuCdo
d0nHIoCP0ZcYPz621Qa9runQlRPq5F7hC0lODusqqWi0B1Wd6l91HkJCyeJh4sVL
0PeVrC+x3ECNWH/F62Ivd0NwWQ5rG6zduW/AgFT8VMrPErYpEjp5IAWcpYCD8pW5
y/JX6+EQH7Ic52es1FABBPLCnNMjhi+IaeHUyl1Vjvr1SaFaVJR7WX5wHCC5s6i6
ZgdHZUka+vXUjigzhmHNHxCfnODZk3MlYOt6sgMnMKSo0QARr9V9phyS6i9NTGLk
qNHzOxBHrWRPXu3g9huVENEuQ4dubK62T33T1MrQlF1wMrM5X229ycVUe1jRqv0J
i2KDc6VUqMf0C8BOWj6Skln8IW9+MCNqjgi+fEngxGEycXE2DqBfxpey6+kM8VVC
LU3zCM7stI6zBDf7o7Q5BP47+6/ua0IXRNd6g10tcMbRVUPfIIxPFJ+vN05W5APv
VsvRYIp/kYqmTy+G+2QiWFOdIYIcHPHo4Mn7lC/Axi2hT6ud+2ZQNR6qavmRB3Sg
YV6poUMqws+7kyCM8fm7sRdMHI2M5V7lmGKwr37pA5EgyJuO903wqUes6AChZOZI
7/NhVX7iGbau+jdVuHhh+GXpntDKg0G8y6yFt/VHdJZnmcupntBNEB10ZOWN6aIF
XqM+q8noywT6vwRW2tXXPa10ZdT8+eqz70rlraW6WC7FtGAT9gCtWeyAOfHywtLV
FDmDCvKmLp/YvAYZTajNcS0eel+2yUDklJiiZdrXA0JceNyze+RpQk8iHReEtk/I
HEInFHrldT69X6bGywBoyyifgydF6Jfqcl4x7yJzYyZxdcF5S8Vdr9ZlVU1Ep83N
Sf0CYx8eaBsf5gOS4Y6wJLRzZFgPQ0mY8ZCVRB3lRlQQZxIO2uBuvmzh76YwLjwp
Fresf5x4nXFsXJDF/Ts+d4Btdl9fRxCXbkO2gCUvAMBqDzQR4HnO/0uyTZ4osE55
nHX67Mij/1Q/PQKq01FGM4QJKmOdgAuZc3xoTOuhqx/bHUgF4RqUH0el7YJV4e9u
5EcMhhD2QcjGzyuUSXe0zirTnJKoFPqtKf3bRrzxOdyzBzFwdMPJZxaVCL7LhXw6
pYn0Z5gBBA1dEZA3Wj0bpjE7irMhRgRg45+TpnQvtzX7AEiTn6rSQWKnvkXVbSL7
T8rT2Nmx6OSwApIfjqSno/Zsv29G8v3A1zxvAx6eDtSscPA84MPzUDm+LObQfeDX
usXXKK+6P4Yatd8+zDA7cub8+gtZc+DvaOLa/K2THg1D6bfNstOJUkni8K6uORTe
ygT7rjni66ChpVZsfqD4Y/gmvX4QXb1cNmL/shkJOqKt/1Ry5pNdt7U5NP6HN5LB
RyKXUagbXKf1OyTw/tS9F0/MOpvhUv5MbCXpUqxSPGA89SwQKSzDqb3c48/A4KPz
k4MuuOFlCYM+sRRDJ7abMObRcwjfE6Dq2DBLsPiaK2P2O6AdyCwwsFYSzFs1Hwrm
Wpp41Tq6Pn8Z0wBjFe0zTy6uYk5n903+LiS1weo4YGGG+xNUDhnpURfjx19L1EHX
F9RDnHeADsanx/UJJPYePCXgSDmiKH3HfHKE8NknSBHreABUBV5DeZfR/K8azlTX
wY3T2m/V9uwOwX75B6lyf8uAT9EYYiHuPIxcxtfxr4ic4DGn7drE7TUYqvkvPkn4
ALByOl+kXHGcmZ4bLxh3jnRf+4sqdODcIL/qg9aWgPjE4qe6avw0eAX1FUNVt2na
lfqGrLzT8/cFA9uoS0r9ZtF1C13ZJavvLPLGNRRX0loM1eUI6I2RXGfXq9kTx/nB
OUI+DvXq0SID2kzPP/E33tyt60vAh+MMk16KizgVrDLD0bSgllWHE6//jrkFxDBo
hBfR4dpYZEgN9bQSEijcgiP/0IAhyHrKr8qyNVsHdEZGUw9jUHQLRqDNIwfHbgCe
nPxSjVuA/g9gF64hpnHcp917zrFWNTEWfYfjcQFqvT8hEYTDDPjZsy7vHhPiouQi
VH4JWQVfbsx2hSHw+hEYTOTFXAu4a4M0D4bFHMuTQbYZDytkhK8iF3UdM+CFAAVF
lg6JVx+jhLVUe/nDcjtQ/0c2amO6CRVzaPFRVn0k99qkBUn2p3teDEJppwOVxnBw
sDsoWy/nBaH+8+TcqYOsemh/jBTtRL1CpL6z1PLVkeGlSYnKcQkylm5zd7fT8CFP
qGFCIZ7a2xlMuwhNXwKNmSeFSGGeNf0IKYu6nwJBBDja5AL/15mg7D5PAzMScOr9
sBZq3EYtfP36nm0S1D7KBo3x0gE8dQ/aY+XmwoCIn8nSg8FyHxia8pmh4UP385T2
hN+shtf8Bv/6s7PzwfNhWSEfAi8UQWgBXXoKVaZkGeWsF4eoN+8NqJSC3K4zfhXl
b+a/Mm8UkbXJknP+enf1pH06LcSk/6JWX1WynFFu3KuVPIgeAlqahJEifhsMhBHZ
GQT25HAgl/8jeWjYWdeq2FkdDt5pRw5tWEnkt3Dy87S+lLbJpCfU3pVHwvoBVhjI
hkwLIZu6CMf2/cRQreCJXj7Em3bjyfssCSXYXsvERmY4Opk8j98yXZcTjTvEK3M3
3QaoYrf3ttE3lC6Ow2QyoYj6QMOiXSzTwdkDzd90esf+yPK+QiCiIb9vyXqCNAre
QL8PtRcW/dQt2RovrHiQ1HEjxWccgV8s42r8P6+ESsOjo7xvHdyyiKjJWrRV45+v
Fq8Wd5wS2qxKbts03cjeZi9aH7kFIWPOy2Ns4YT8pqh0loAVCEJTIKu3Pd6t6gin
T0foSkPvjWs2bfqzaSy+k5wEvLJ3hF1mLE+kydDZGtYUenHw4/WId+qEOlvbKnQQ
qVtC6nsNMA4OXqy6xTQ8ytS/HydubZSN6YGV1z7Ip05MJ3Ab3nlEuXQSn2YzwzDC
wPN7DTrBQZvNRmFebHHN4POx/1Znz84R1WywBakbaYMU6LOVrrt2a4pth6h6afZP
lH363kNBmkAyz+oMmeKf/sGqHg16baK2d027EJBkkAWvR8iWR0gwTSh4p1tJ6MKV
VQM1TiscvNgDf7FJ2R7pJwsSSqWncYYACE3iDv0vbEUp81zC6thNFCB54cF9kO17
DYkgEwt6MnUpA9CgXh5wzL/uxRad72uvGBK5erPlEmpKAU8AZAuaCxIjlZ3HS1sj
EFXhQrJ+iqXguGYceUsCQlWCFHMF8+qhIJaaMe3b9WzJSTl4QcBLHHcEhM9dZOlO
EnT02c2Rg96QZUR8MmuVUsZkjCFXxMs380Apv+YrJMUogRGB4IafKvJpi/qTF1Qb
ZAOLjYZW6744DFUk+vfjvcwsJPaoh6D3+aN4OiOURHLPSxigQLS7AYO2UOULK68n
6paHLHS+aOe4dEj+8MWgmoYiDNCuUNqblQkLiZqha8Zn9dt2fLMf7LXlK2qr86SD
WFISPR7hJ8OScfN/dXs3HdTSkXvmkefZ9CfC+fHKLut4V9zXFD89xqZ1P5fxsLWz
IAxT9orX77JQ/I4FLH0i+hTQdu+3/2LoWHLM1hF+YFOQglTXxPm0RRWOw6Cv9Zn4
baZ9nUKUpQ4krhojOtT97ClmYFPpcz2o9WAiQjhWa+tX8AK8dRbgyqpg1kaVJU2Q
VtD2DTY9Oe4hqBpDohHgS4SSfJNvuTzPOGLYBvd1Hs34Ljae8Zf9MSa44jYZrZ0B
zweGk1GQToLi8xo1/FmIfvKD9n+hXQxio5rrPfCd8fI+3ohj2i1dnCZLBCd4B9WM
aV8/YgOmUgkjLI1utQhACscWnbAt06728wAAi7QGpGVoFkedSTiXb850ZUsRB1dq
3DTG7Eyuzw8XrGNDDcw/gt/Bjn8z4BqcqpvrLArWHMJjXQ5DeBpq7Ax99KX6yUVM
Dq45PEQmSW0tlVu1R/JVvMaavaz2aLIEbrpgftrogmtKZahoIWsNwJkOcw1XbCP7
92XCr2SCWtWEATtOw/HhBICX4Af9Yf6SrQX1voYEhNEiLwlZic2JYbxFVE8imqHM
KVUo5aBBpncp8/YyEdVdkEabUWFjwGrT4t4iVpBKHJdOQN/xD1gqNNPyG8NqkCdM
cpkyHbJXP8fiuJRb7qvU19cpwHYe0dndw+Npw1fev94hAz2t4C8o+49gDgAKKFpO
SiQxvILhKJmOoCCx+iJkG5c5GvtQHw1EhCR9inwI89me6TQeJKPdBz1kYvQKpp71
43e69aF1Owp4iSl3qMocpKct+3NUjbbO4xWledNBFhL1TBW8f6hECloUHW9El/cn
lNSLTOcHbWIowxxZHmByIOXbzVQYL/EPbynmkmn/TGePsL515yXr+xBcL8gyEd/z
HfBbtvgx8FKgTGz/KFMCw7DvLytj5LpGNJSNioFR0cLCjwQRFamy0YoZc381CGaD
FBOw4SCg/uivSsS4+XQHi9D/8YMfvd651LFYPPT/z3rbQcdUW0muZwMxoWBoXYpv
KcK+PeG2Jxtu4YrYVuAnN4G+bKTVRTHaND1JQRpjB26rIbZa0yMw1iGDqigk72Fm
Yi3f05XHA/M1xb9PEC2yiWk7ppGoUcJgCnj5C/uBpdi6+dQ/GeYel4Z8C3LBwwvy
nEE6U3pLbR0REip9MaZWuSvhzCkDKS//jP1WIXhIZvZKpfJiXxSoaOEy0av8bfGc
v3dNA2N81pfuMpz36ehect6CtrkEDMhWp7khRlOjITvTNWvBvMhQl3eG9+8BcYFe
QppQsC68bxRIRV8lADnMdsQ9lVmq5e9jnNNSLFVc+AxOuasL+nS7ZSt1ZVB66JI8
tf6+FdxxXylP582weEQAve49tfIOOE7oXk9x7fermxJgig/FSy+qgYX/CYMGV7Qv
cL1wu/mQfeLNnVL8lV8eeGYXx6POWyPYyPFH3keun6SV8rZeOgtKSbAkE63rlmty
zTZFRbnMeANtXDm9YeBZacysFN2o2y8+H9eZn56QzKE4qcjcFedJ3913LOlN2twL
xXg8JPpVefukz/a/dr/6ORqoX19oO+50GfQK96HkDk9n4Acs70FTaXfUOtrTZ+Bq
SDun/t9W5fSEoiI1uFSidqalX51dRxmcePyhXnUNz94Cjj1XqOm6LGt9zrppw36o
aF8IwW48AgmR7rv9Ysj1oxYHEgxJPQAV9OaMDm7LQlknA7z7CEzxskMinLitbnI7
L5d1qD53BCzB6m2qRhvtEs7pIiqRg7DVWSMbIWu4MwPktxQZRcJN+4dFkSrUtTRP
O5nAwh3fvLoTRjmd/jrm3Du8zMFIjZwkb2qNBHtgyKulzvJyUmKF9qsDx/iaB5XA
oY1sTAsa3750URsRX2zQqZKyE4h4K45wbs+JgjEeAkP7z8soJjNQNo8WRIC9AOA1
rMmEjCVvU9n9yRnCVm/kh84orFdApqOlnmB+RLapj1cizoQxe98OCr+5/h1ZacZe
CfaQ3vDGAGL9NIa5c4hdFqeRYIybg56n7xPIO8udCFX6QNUK2oRu4hsW546DvQeW
XarIX/Es5/qx/UgIJR5ss+eQsoE0pbJUNzeMnH+VmgfbCL2lgbuD5CNZD/GPkwTE
/KiT+7/tlkE32Z1OXBfhYDS0x0l8spKrFmkKHMlJSvm265S+fMagz7cS+4zxuNmS
QLBFMxEstNzUq8uKo8syZbHxkzeVRZtAbsaZPgrrhQnS8XIkp6Orh7dyOMzUUcUH
5e6rQ+ovgoD4l1N4+XUO2EYRfrGQMaMAicq04m8HsdnKtb5wdwr1aOKFcT40QZB9
RnKpOVlEkVstUq2z7gPPY37SU+q60cvV1M6lQTa+sXUZw/LajwYhETE2VyN4p32M
wSHp3YmQRjxkm/VZS3xWKU8PGjOkde9L3tXM4DM0C8IGD2X0OcMnO1BEYPcSDEKV
JR7pOfEFthEa3F95aDnB0pd98yWR6r4eiXWtnFywtxz0O4mzEcsBY9wx+A1Pgb2M
jc2g/wEJ1+2CYW2XlKXJuYanN6ed8qv4lJYhxLZe/1bOVOaz6WAxGB1c74yfeopJ
U5CRm8laljT1lJIJnPUo1qRYH9a6N/5jC9zqYC2SnSfG1/zPzXO/hwiIK3QxgDiq
VUoOBbXsGhl1SxAHgKri2V4GrjMCxQqxlBUiwNHpW9zWG1reEwj5a4CYREeJVEHk
ByMf3RFjDu7IAZ9r0SPcyxt0UPRFKtLo1Z+oQAN9pnGbNWvif++0dpELWmoCT6HN
WRwBvOxTdNgJQOqyQ8cwA/7u4kOP3AYITSkXvebz067QBqif3qNz90r9SEuZpJl6
xpumaeudkN0hvGFRYeai3DzVjHJTRT1474FK0YGSYwhXjRjktHFhTzIdLVF52Drw
YdhvWnqHxosxGIkrUw3rQbcKk1uCKU1o2JHvCERGx4WCfSs8nGKV+KlxVinEuDNz
/XrhwLQ67F/HwPsxYzo3cTo9dRUnGe92ins6grRejT3jXGU6rvZGwvcOUbvcKPBS
bX1qCEHYqYcLERKTQhpgVoR6scZDBQ2eeXhcV/Xruxvnzlawbzsscp0OV3wvIubl
DyWegcE9BQfeKhZbh4tFhvommX+qWn62ivGEns7vys0Njgx9VHEmxWF9RQ748zD6
w71p1CrqTs5QD3iNpnUm2BwWT9/ysKH+8vdOXsOIHwGQlel7WcOg8iuCYcc1JP6H
r0gRVHD7A5yS8hEV0bO/xcy9Ha7bQUOygMyK96JC2S3hQnQ+iXqn+KI+juGzaxzh
n7J4lI4+Rj3XCdqMIUOCPpdo/GVTPjnVgyo2Q4HBIO2fR6chM7Zurs5t2dTIfgwX
j3OSpXxZc3KlnZPI6VlUplotqlrGiL0xlPyr0BPXHcw1S7g5QHzRHj4P+Iwj1hGV
UIQR2s4tqN38mZfbJyPP9X2j+meFhgPZ/KUmlzGOcdmA2Jx6ZUfAP+07SyKzIXFV
q6IidIsi9ex9oab0reJ8YxLswh+oosF0jKFn9+kx89wSjlevinBR4+JM32lwyv/N
/5F/9QPZ9pIxFrespd74Emfme1zgCF0QHJC+Y9xMc8KHVgCs7XDp75PUQ/pljAhY
KEYcDatKUK5FxZMpk+yWCLxwhL85NJUqrETbLTafHRenLCe3pv3AEBtWBrncpq/P
XLUlnA/haOlurS6adSIeXO2Rnul4giPVcj/pOYcYAHNzDCSydkUBj3XMOdDtGULs
LyaZ/FkrG64veTcPsT4Ln+asnZxHlQsya3sGRh/wmqhq1rgYA3LgrG3CU9nY+1I5
nhMBUZw2drG4jbmf9LZclDjdsGrR5RbRr4U2WRBjYu06WGAGZdcN2e7zUuZkvCoz
wB7hbgFTbbbj2s3RAdVrWWod8AyTGodiCWHxgx9woonzcuAE+UdPiNTT0VHn3N+G
fU9kQPP8whQ3dzH6WdqRCUS3D8ScFX/4tgCr5sYB4IHKC069geLX28vsoaRUKvvV
lArH7gaPygXgznsecpL2owA4M2DCS685/juYOkiOMHnldoZtnL0x3Ntfs69TribR
W/3qHHCcdYxKn4rhnQJ15pCA+k5jN60Eb6JBtwyezz/pwahgGgNq5wkW0DBfpOzK
be9+meUylJ3DzGANpUJIrAic7QFJv0IoGf3kBqShX5YP1JwIUqcBKUa+DlJ62bsZ
IQiCBkokoRlhB7n4GZ4J0EiLdQlof0znFb4gHBNwDo9X+LBNscta8ERBnmpwyIZn
66F0dlddIW3lA2L1nO4UzfK8VP4+TYCdXUsgWhJZgrkTwH0TCl2dDiMaBX494cMk
U3hvUte5WPbXjQLI7v5QiQ+/2eAKQ2LUfG7tQ/rkig5I6to6Qv9mTQMlEFifwLLG
gxW5ZEmvqTPo5/OqLKGdkJehRXlRcXunFpv+VpmE50dzLFVxI672rFpRfT2BVoTT
uR+5H1TZlymRw2aL5/775+0/zV1a4MflTjoR9wZ/Se9hy82UewlrzkjWSp0QEXxe
eqUfN+eEqzrE21J9gCAZbdEg3gVunEBSegg1QV2sPzjrHcWoBoss7O/XoBB3O6u0
VBsUx7xAv0OE06QEnYbEyoVjIyqo87p5yxOAbliKru2+XH/xQybRteN1HirkqVrK
KrhZJQr8Vx7vF/9pApv3Zce/Sk/3WlJyJEMwHJQUyZi2F4t2bMVJrsW0IuX+zlds
ld6H6MWoL0qtxjE/SvIMuD+ym2/rmZrwH1AUWo9Vj3fjBpdxjPZQvdcOnSQf3mq6
q0DpRSHmUcs8UrJXVVJS7JHb9k8rsEUNuEpy8ZvE0Ol5LLGPiFCyRkHBB6P7EpCS
PZ4MIs39ipj4teCuV6SUp1wzMkna/cagV50qj9OuwAlOdGE0Oq85zKC0UW+ajc6M
dQZctED+7mqqRBztdbDLEX3xSdFrHpwMvdUZ6aSFMpEFHcc9uJBj4IpvK34xV2vq
GXIjeJI/fMqi/YvjDJ83SPpcBtJ/Wd0/6PBYbLrrz3zirVyP1dvFgWTTaHsasb59
shr9nDsq4Xix2kb4Pfi/WUY3iWT2nMpYifoZ0N9tF5+54kZZTyDV1YLOqsui8lQ+
OrGM3ztM+XhoQh57BMCXi2h1LtvSsxZPNeLNCRWu2ygTVFafczpH8g5YHyF4CeL8
d6i2bWSqXahjZRCYHxFlY7Rk5ld/uouc9FpLS9xssv+Pw43D/S0B0aUe7CMdUER1
+/LRUSguLEV2ujz+bbpiKnfaDFQBUtMNUOlCqqt7Kbcfp5lu24atS9p/qRyekTq1
c1HhYnR9/DVqlaER4e9u8AF76xdlcfR5x010T8GWogGQqBHEiNprguLgJnN4ZTp/
1VpTreDxjn6s74ntvrdhHfhNCWW9bQ8J1Bv/CuFC0m+oYELtmuoexuUa15OtSbKQ
nTJ6FCS6okjdXie67bbv0hz/iqnIc3BTLcGi8TrN+bjziSpcaKDzCtny215kPqXF
fkgTUiVnnG3uj+u6XGZQIXFB6C3QGXqq0mNdGcxhr4KG36eiZz7sMcG65gSG0QQb
yohgo3IYmBpQocP1IZJgp3W3xHNcK3UOkX8OMRVk4yRAgRJIr8jZ2zkxAKgZHH9+
K34RPG+qTrutCAJUvNWjHxnDvQy7Rn9S/ymVZYf9LoPENFECnU/WKa6AAk/PCwrK
+IVgg3WNY5PF3TteMYlGMc1AvDFZwT9LRvuygjrFVyQnx+G5GYVh2CJo6dgbh9vZ
MAdgvOjotieniGdWQ4U4oQax6OtV6PNJmH8deLK2H86KAZKQVR2CEDG2i6ScmoMW
SrwdZ2ZviXNiU/NfXMgBQwh/yIumdGKfqWG+Qb/98KIoG/PXB0Df2TB81q2rNBl3
716wVRTUnfQCmYdsQgTa3QkjhpphnTY57m6zGHBRWT4IPh9AunHjm8kUfaRKgcgQ
auwLSa3oEXmk2ai8N7C41wk1Ne7t2g8kVkmWhopH6IlK+gJZ6AAU8k4OdxfvVPzl
TgLEnx2aQYbqQXS0bZtwzOYSdPo/deoII/tXRDvGZf0KH21JLT7JSit2iWWckL/E
SnSH1IP1aUP8xnS/GPItkowvLSx4hoa5JNxoqHjacdgcu4v+ev8Rs5ADGpOSBv3a
0+oGm3B4XZl8qYQb9I+y9IhE0OEpFmsH2+IJilanrFRlURq+jRV5U2lJ4DDOO1rr
4Vhu5ZHz0g6T2PxUknQV7GywWv2kPAp42NYSq4aUyiMDM5L2MjNw8xVk9b6Ka188
5crb7CXEhFbe5E+3WRyOLLHayuKPpOTF7GjohMAwHu/3a/6z11s5VtKos1quB/t+
fon49CVZiBR8CSrOXpfU/E2KCtAJ1wFQ9utLooswGb2Bkd0wbjIQcRqkMadGMuKV
PCpX6Y12RSbCCEbWOTcQ92cyfqhgOoJ1EJ3nz9hXAD7LHklbNUcMD6Bs7CeKFz6G
EbeAZOYvpQIGVn58Lk0VKKta+Iv/iH2zyozMO/AYUSrRj/r/tE0oTFEbTV6THcu8
G4+GC6BlMl0iyCHWZCsbtSc2xeBS4Ll90cN/x1lnj/8JvSfWsiU5dfYIbFJxFmIH
hhmi3gmLDnPC/1kKkFk6y659SdeakqHvTjA01Qt0PT1Ir3xQVZ0WbrxmYZFcff4O
Ej3i6jrokgMIURIY0X3Pq6Vi9jvz5iEgpyNqwgiWqCwKmWR7uKiKcYPFPx55QgYB
dew7YgLEygbnZO8GoGUdqXFN5wZWJbLZTAIiu8OQeLSn0E2MEh0B8N+z1i7PybOT
wuwn0sGEpAfMnkwaQ4d1mksIEPe3BhmFyScOoH6vRkHeMpuvVRSIUBaJv2geNzcC
H1k8Lu8S4Cz3ydVWUwFeZxMFVQ+Fa/mZ6BD3Mtgp/5h6PofXWTGFT8JV725lR9R5
wd2d5OPFeQiOOxv9ffGQuDKMXWzpzeHxDshhuaIj/Q5AZgVGtqWG9XDePIyCRWWT
0hUQDfO72A85dBU5ZupiAXiWUPva5nexXjDCEUFbMSX7z26EvfB2pERNxU54lzxQ
l+XbI09nWBHw6dZbweA9txrEWiRKwJch7jxJPtm/YQPdXpgmzqgzcAucsmFFZmLh
rItCbxX1uzykVCZBndtw1cSQKrPb0kJZGo6lqZOuNSDvSUmaAHbuPZyi6RFWu481
S25jMW8NPmXLnpkUwjM4TCV5OxDitsAJI0orHTqepY+tYQ/2HTmfhCRhEDlSy1QU
CkEh7QKbqa54i2droFuCMuWM/m5oryyw3934aBXVaypLj5cHEF9Cd/uK70qO08S7
8FZ4SmtKkElOJ7r+yryEX3FKO9reYGtbtATulMdAECOV+VblsRAlWKY5i9MerGOg
6jVdTec0V1e1+R9JhmSIfzskr95HqFHZi1T665N9H1EPvjbDvEhtN3aGqRVl8kgH
9qKI79OL4yE3KCCXt0o4nHLb23W+hcHFp+h3Q9TTEdGPlvGrSCgv/vTF12ZQEjYi
Oy0O6pLcYZisTPJCKRPEOpJUOdEstAIMyxcB7YaTb2nzF7O0rNNRLEX7GZvEkiCb
g8r6tmWuun+Goc3NkHyxX/VBqe4WkyUwfXiVU6QFOwzqkq1YpS+our7ZKgSgRoGv
WKOftI03qnVVmHK6yvcVgDbat78uTXftpxE3DdWpA3pPwGpn8TOPHm3xW+wVbhsv
8cofidAZedZLT9g22nBtXwx8IZg0G53lJihKL/8V1oa8L5DuEqhvdyh1xjH90sGo
rMh5lp2ON2/q1FND9ssKHzEysqnqvvrm41fHE6/ZUjNQ6WKe9LEFhmxpTAhiaw4e
KeH1MntXyrxyc1liI+b3Jt3nsPqGJJ1VBwfvUBZ60FwJRSlreitGeKivY+NVtM3W
zVesupRW/eif7FQVzGJpA8OI1NqirU5tflsF993GpNy1hTykV3G/r8JgFpzwk3/b
+9b4Wa92yWWcMVdA083HwJXx++zn4cNWyD/zD83jNRd+GiTtLQG/ehSlgjctUW7B
EWiDEG2P0XtoFd40hfaDJYTMataed3z1V2QXTyjRaE3DXiatvmJJHFHQ+PQqUwHI
ukWZlvFYdzbRsR7rXVUCRLD1H0eiLwxcioq11tEHRILPq/Wbs+78IN0MvtGQwyWw
LcIPYG0zf5hwdlgSs4kV1UnAfsirgybTYt9H5Z0U85m6vUsVme6xrJbVbJvwpCNB
Afz8HeDtjevS70sWL22Oq9iVM5ffM0Is0I+XoMVPvaqveBb8FWFXD1TIFnhyz9Nn
vx8tfxTOU+61ww6g+0hkE1OoKpU+DmNIknFqReZz9oItKSEgZT6o376aCHxZ2RKf
v5tC6k9kS8NqJx1RjfRUCEtoBl5PfxCg0LaE9PmDf6z0mwhTNul/mk/KtF7EYEAz
4vi5+hDFrlNR+tfNAeJZ+Dw3BRliFpuKdkzbSGY/j4WzW2k7x8+XVLd+D4b3XThu
duKE9Iv4hRwAGDVnUryiZ6oUy946grnhdTXkifbop/uFhlBum8VdDs9pH/YZCB94
dE++BRNUwiolEyd/H0DTS5vR13RMNfW618iLPulNIA+Zjf3Xha8X0EMjxkSXPJa6
sujEmWWv+8Hjflh9DT/ZINXsVBHv8ucYJN2mBmI9rTD+CLAgSxD10KCj14jW802g
Ju086Dbb5DZ9XYYIL7SXGTU1PBjJ5NbhyMIQcm/fD2DFqZnCelJ6LFtyKGkUgMeN
y/YSR7XlcW/lEAfguEBtWCO5AJUx7yFFhpJrJkRdrywSIuz5qPHiJabDt6yF9oId
1eu/qL9Ho/BKzT2K7zwQmbKOOu3Ml4D+82/5y69BiYmvxRRJfyqRsHl36h7PqzC0
SXXLZuehNnQjchzllTSMPhnd7kMea9zS6TQWD5IVZq2aIBwfAfl84YTXcHFVVG35
QRvwKX5vBuV2UGRV40RkBSmnHR410PT/+w28vL9Dpv0XrW0FUB+1hRhNZFjmrU3B
dQ2a9ptn5QFm/D9fPBzDefc9K8mTDgxNuS/V9j1Pn3Bwanpn+ursFW6z9J4NlANZ
paElbROOi7PFBuAtgGMai0tebn8JC4bYsCqTyVmk7s6wd1ptUKN5MKbuCnlc6rNe
S9zIl9mazS/G7NXPG+9uraG6vFzjEoe0ysE47St9zc9nmjoREx+F/l43XP3cqrYv
6h+eb0msocTu68jfESv6d2xbxQR7gxVC4QTE9qsjd09o6J8xKaM0sVVs2VywRGja
rTAPM95BU4XSA2Tic+8o5TnEwKHwRD/41CjrUUXJStRCYhQqrONJbnYaeZcSqfu9
zQhz8LefJv4/S3y9vCVI7vpGjH6CYqtgn/ZLw+y6mzaftkoj0k98TD0m1/nLukLi
m7VwlE4Ma3bdtgc0AmCOjqizCEWaDJG5pxU9aCpru8p/VigxHKicpOIM1nXWIGoV
jHpQHS5qBxqD2i5003P1XS51+rGjxYsCjbNMPBGQfEuEAAkeAknRgn+Z6R8vLQwJ
sSupC10Moo8MQfYgr0JyEs48yuznFfQffmaySlYC/kSL9pzWn5Beu1oUdg4KL87O
9m+9Wj+RybIBsjinDvJpbNidg6nXEmdyrbBqTn2+XfmZJyR7GyB7sq3+1rGdZTAi
SVAnNvl8NbZZBthi0Lrxh/bPzZUMGT4MwHhN+6LbuANRrwxAF0T+DJAi1cfiSZEu
O1j0IXdgraEg+rCfHVzUei+KwoA1gYbnrPkRR8ux0u1v8m5/3y15OyH1H6JboiRv
eohLD1mrs5YfgaifxJ2qehBC7FMB9eZt2vH259ZPaCoytCtarM6wSeKRfHziXrL8
Es4JzB76TBucrfhV0L7n4j3I9R3EuiPo3OVqtXEYkgJWszxE6yjcPxifs1v8DIX2
gTk6hEQt6dDFCSSNITBNitC1R2lMCpLdlAjxUaNe0178zf3Muk18Ub+vk9Pss+v+
T7ZtLOyQZ5sULR3RATDC4Hn0/XbnWRGcRpdg7Rszw4wFfl9hHJodJEVhd+b9cSJP
B1BM3GrQi26ypeb5PwXVpCA6A7DOx5YVGyGYZtcONXNyODS3hCG7p20r+G94WSpl
oif9w/Y2tsOV9IJj7vVjI39NYBABdWcwNOK+yp5/JVFNxLZpRkLTBndanUDlhspE
Sm1dtYvroPdhPrGX3s5OROzMX1up8mj4M99Yq/ea9hrwrbW9cAbOX+SmjCmdYcfu
ENoKJO2A6oTZmBDZSe+6FEvT74neorA/Yf3VtyQFyMva7VHHSq5kHBeT7lWwzo8d
wYjqOMZ+TbY+meNwUlqjgX+tykmhtyXQuO+eFOjwwHQOrgYiHDGa9Tt/mzl1lZ4U
5t2LHqxa3CK6F/RdoUdr9K08PiHgFYbym7e2ONj5J7dFsX8MboHPXnf3Z0HL+iV7
7IIcjCVAhlcRkdWgBTpamHK7feq3Dr2lUMvaq3oJ1IvaemxEARmNxXq+iMgcYsgK
uzAZTi9Nsge2bCWEKt1DOjWceVT3DtSWOyuT7wfiFPf80FWpCKSJ3TyHI6kloaiz
PpUL/VDsWJMmDmaU9wDESYkoTbG6QowCe1yMPmGVKyFNw9MLZEYYjwm2YsToUMt1
1/nKr/dEshsy6PAXZYOIclT9M+XVkDmW/vifgxNkcE1FTF+VTq8+V/mLVVmPQqcf
WJgsIyVU2+BtAzxZz3IoPIdkraJeB0eiDXkm+QlFAATP3lTZWH2j1n3FGJ4vqa4C
eGXDo9hum8qbiJW71f62s/4lT6x5aBLJMy3Y6a75hP+hYft1WsVZzVCys2446xBD
RAnVXn8wpHlWozPbkyfWl1cc1GCvGxfpKVqjoJBI082CafDLrBue7C8MzOh91ykQ
FK9FQpnlLalVtFtmqj7y99K9mWwacMgeCdW2lmy8bRFo1Lj2NDG2J3UxmEu9gikt
il8HwXAXIcyxZ1OoM55UHtrc14wsSmhnhTR3eIKJj3D3JesOUcpNyoEWy2HMBwkO
iGyMPDf6rlDekOPgdedid7ifd+oRTHIGwxVzAJQqsNRNTOUT3FpIJB5X0g3iL4be
ovLUVuk2dqZcdXWyscQy91arm+Btsj8cp87ci4LCtZev1v+jm3LGrQKrs7MOtPjL
Vk537uj9HB1me741PxCSsdsiRnheNxHa/XVMM72HUBRFndMFU3phkhR3Lp+TQotO
lCmONw/O9i/NehmcqcWT2X1BWwCgi6yg4rm9w7V2dIKQch9Qfc54CakBUaiyRiq0
l9tdfVVrWgb7Jle3f+r3HZoBkZUxKmuo04z6iyGEd2nUWW9oBgKKDmDbaLJx8T1s
lpRf9vsX0w5Ram3O1KBl8n3wTBIV0izHXmTmRQGAqXV8euxJbSYW/KnGglraH2X+
T+4qEDWTivlqbT9ZJwYrOaY/g9ZSTHLD93xcz1BaqWOt5aL0lU4pVM6trkN8bDb+
bHKfYITIiR7xMm9LoAmD65UsKzj8fai0W0yDRX3VJHLhXoYTCHWsRxFGiPuumyOI
QJMvoWmCUVZ1pP8Ti+yFvnGAgZsyQ+wuOJ8udzOIddAYZrkbHnw/3J9OSmtIdnfd
LJsZlKCXNtroA3IqDs4Wo92JEcWy4wq0iSZqbv6eV5sdJF1h9xAPif9JDEckX7eG
xMGhPXRbxjzQnpHLVkpPGd9UmpT4kdbtG7KDNDRMkT8WheU20mXOCgdohG/kGWhR
AN+TEjRg5Y8u6H8e6R281B7w4km9xWEZRBM6iy25VmvVGdPJZeXycfW7lZdeuSXB
DRsmjrl0n4C+efHAHa5xwNtsMsrlkg+oKI0gbo5lno3VthD3T5vKK0m86WnQgk3H
K7Ip+plj7LqxGjTKJNajmDBocKXHzU4QFWev+nxxhc9j3Fd6B8/1Dqbp12G6/mqx
/APVjnPVA8b7TLZCLwRzyMe7UAMdjleY3JL03GYWWjko+AkpfFnfeWshPM9mDjqs
SrvWhuhjcZTR1zaEjjkAuJM3Z3erEco9ugN8K4RtVoHQyQrII6SZf1878oFYnejP
X8ZhsMMhiaNS5tJmyHju9BP+CgdoK7O+rzljyXaNjo9H1Jc5UR/VdORpv2rtp584
vlRYxSc909PJ0tuapNl8vjVT3/nCDtqHZi9gIKnoVwXkdU4fJwvy7yXbD31UWv7w
KPaf2g/NvLBM0g+igftFPT6h5ZnWnb/qqTJiuSv1aZYN5XljQRUYmLmrFnY/ICmP
bKYUww5CT8eIPUWl10WzzqH1ukqcBE9MRWRYxg+ZWCPwBXlaxBF/6BHxEY5VCXeP
DC2zEGBkuqgX/Gp+h5Y1MpVzDAWIPKVgcVJYCz6J6tuRljqqPIT+ioqasM+diYmG
a7+TDpO9AJgIhPTn4mrcCzSsemNk6KMF7YsRP57YrQ2m8XoBEHpH56ZJechg5IyL
ll9p3kg7oc//aR8w+s2Fa1X4UaHir9enc43Cr15/2zAuC+O4Kg6V85tA1sXhfFaQ
xy5TwEaWCbNn+Mi2IBDyG0pj2JPBcipi+JfzqC0GP95Tj+j5GWRIL5lUZTwaCfm6
n1Uw9aySzJFTkJXROypmGFLp8Wy4iWADOd+8C++pVUBB/MBpoBjs3looLhFO2Q9c
aOVdwfhYT2ecU6wjyIQIWHn4PCHVyoOz30zr4DqL8Jgoq22UmRTC+o3HJL2xXvHx
hWJuMvh2BLeNyzlHqJHqZirv9A1i38woSGQI5++wysV056LVBn664sjNf8pIqWF1
9WKDAnvZ6FbeKu07lfW8697DML7Y9V2FSad58TT3nugLw0Arp/69l4nT5LxZx0M4
pfmkUGycOgO7Rvdge5Kq014uiONGah+6jg7JZPPVf5RGDA+IBc5FP40jJ3IirSnP
AxGgNKMiowqz+p+L9E00Bt67a3UUjotBdJQoKlw/nE0pgSfHhLWND7r59DHBwzy5
5VPiqOTuobbSmi7PNImtP8eRrGt3Zs6SFMLzd+nRS3hrCbAn1kazH7yGjNGcBks+
2S7kQHH+OIRuLSd2fzcygg+KH1O3dYgKWnoyUKyMXr1e5/BVSaU5soQ7Bw1zZrTP
6GWljBPKS4fTWvHksOEeeV+xbVfvnorLvlcbb5Z/LwjfGvF29MiyyqJgIME4xPZ6
eMkxpCbLt7seCe5Sw1YXPBF8GsI7UJbX4lbsz4W2k4lkk6CVQF0U7y0ejNbiEMU7
wwYB+e87SfB/Yz0QzPMavbGgbuGs9jSyFIB5CJG785ixKsUt10yGmNZxcCQ4KbBu
iCODW000jOOd5ONdCY3wlc50ExNHnjJI5G0qO9Snw8QWDYkMpHt2boG1HRe0zq13
P1SyG+TvS2OZ3xrjF6ufck04N89DusjlIcdzV9aMB05cHrTWaGXw1512b0SPQdNT
gZg0mf3Ereqeq1odGhYM63mPnCpjzQ1HHNyQRVr7deQAjnsRYivPw+h7iQPEg4tO
wks2WLw8wb/ns65Wj7khIKokhGEah+Bs+bRvThbyh+/8KbNKMnpsHPHlUc9AiWXz
/yHwZe0EdA0TIcL0+k63E2T6NumUClYzXBlSji3hGxDBPCJZJ7mjVDnXCAOE1W+8
9vG2MXlb7IlRVDAe3ydlXesDj31u1waJvOnCEQAB2+iD8WdAgEsZSEL20LFFqaBT
zlGWrXbe/DavTnAIxPrv+mGnorCgKmQjaIyZ/OSzL9JbD3PaMIPCcz++cVQ7TC7A
DPi0G9G6kvPQwlVCfOjhs1KnlYXkGcCmGzUz5Afsex0LIAn8MWPgVtgfMQe+120y
/HRwf0uy4kvbjCxrayWlmJQ1mU6N7QYTpiT5RuANM8v6HX0QGOwbSsY4deGazah6
aNNMYuccy4PZ45HN5O5lVHlV4Hdin/g1BJR9ZHb1u6d8URSd7B6IZR1VUc8f6fyv
Ekkjq/R9OWT0REawjAabJfGKZ1nKE36u/3SGGtA8GQ1thoxJAVPCobegIkJhBCmf
+jbs4rzY5ERrInTen5jsyz6i1DlA+2ezI/5yifg8t63LSyH/uYyo7IfzFB7H21y0
QKgvBhOSFu9Ay7i0kB/QiF8q+jG16f4jau4hdoeVVPgra7N0KdU1csLpVbmEQ7Dh
bjY2l65ngFsAtIGDpiI1KbzPaxOzPf6e4YNBJCYA5B6gx6EYZ4cHQUKC1jxxPJs3
Nf97SkJgWkU1bgOaM113cgolOv6ooMcFT8qHaK9EKefR1r7kQBWltX/L8xa5uqxa
RQBvVRfPr/SRjujmsNr0OQYj1zLa3jwLdYxP6nbyVAR74DebVsuH2onxfAaWW4zM
V1PYlbE9TNJOkx1kus3c7jC3To5f+jZ3ifwaTxlGiVpM05+EBh6JzVAkNz3BYiHe
B0u9fIkMmjX7A00FQvgzwPhx7VB4k316+Pj9x8MLLqLv6qcA/QbZLYL3WveAkExR
eOtGgtaFhRFkyyj2lRUrQLrP3WdrexocgovL+QuINHnc53qdx1JWjljV+i4NCIR1
fwK90KS3UVdRm3je9dMbvnV0CANTg+uW4iDCpeHD4JQqgBt4RHOZLuagScUz4cy2
52q82lqWG5dL7z9meO0YYlsLgnI2fhh46+O+4+UCy9WZ9uhVMy04C3bvxypLgMWt
wyRJsGHQyn0enRr2g0nR+vFfkFdv9K4EQ48l3fxrnPBu6dPIsUO9/SAdj6PTCYUo
9OGMLpbfclEdN73A/heDnvp3mL/M7++bp5Qr7Vhzh+MzAurhK4f1v57uSeO8QllT
Auvgh/EesbY7fROD8rlm1+It/ZEqOdvds0jp7Yhel0zo6GIf/dJBcVD/hYp1iLlt
YR6Hs22qPWUnSog4gLcdKC2XFS3aenjfGA6pF6fSGtD08+ybUl7G1kpmhVj+i+Z5
jQ8OvcTwmPy6SS0YQCGH8dPws/mrAyfMS4wSCdbPrliK9QFW1XjEjCEnax7g3Jrp
o4pkTRN1T6/H6cRDru3IfGIuokDWCJKP2gOUKI0XrUb1fQL/mZnkZPm5mqB84Eb1
eCR6g4+FynGxlVv0TYwXUuSrBd7LbbqNYSoirzxgHXlM47KBrRH3SBXbiPqCGM8Z
qm6UcTVLwddg/k7eiBPQfuG69RCFqvBSXdS015gTVNzDdFf29tx0ft+7MhHMjNcv
XtPPiCXWKFMXLNGvcTtn4Dp/ZOxy2oWbPrPuvOJa9cz4peuIaICEJyD3ODffgJFm
GZ8OvRos8umcuuaQ6rCZPA9pOxAb+jUkwKpFumCumPkP18lmEn6uDoEUt+9/QQ/E
wwf5fBCftJ1gY4PB5WfzBF9WROFbFYF2AIoRrvNT4grXZ+JX1/RPUsGr0Z9XqqJR
3Zqbb+GDJgsTNgYqFK1hE3d6cWvduhViToo2M5ZbRjVzHW8Falk1eD8MaZEy1BTJ
vRsPnVdcxSDHr8BwteUPfBkq7o7e6Yf5O9/NcCPeFj5GS3CKREtG4gAkIwpVnqhm
py4Q+d3UN3KSEXGd1O0guXu9G3VaYEsDgC1NSH/1so8chS+XI+mzXnKKjNhjNJcZ
fJmS7GcQE+PkFTs6PVhpoAwrcgQPpd28bFk6Xr/XL7ihuXCIyTbbJ7JeCI7g+HZA
hbycZvUuOHCUvwvOnOaR7zVqHo3HCSQMSldTrUixbkpjYZoJ0GkDJVzR4heBLoa7
iwpE7mnMQCFwvjwaD5rlRyQ8ESQhOjpyRIFh4plAO4cFTmN20BvMM/WaUUNXCW2L
0ndmaK463McQmo1EsB7phTTksyvj6fcFUMHwB+RTY9AgXNh2/NDS4DxEv3C6JYEi
uaZSUUKkMz6vC8XLg/TLLbIcpCpZPOubTDh8iYKKUumHtPOuuO98rcdh2+GDDxN4
DlJXp1Ll8EPzCHS+xl191WHOJFasrkWbw+u7G+rwHEkmoB0CIUgQp4liryqaA/PW
JNs1Gjy3tt7a0NF40IxXnHsKjbgmUUpo/LWX5iuvl2d9P3wKvRJwEDR99aosGIEH
Q9W2YXP/ibuHGH4b3PdPIBXfV5pBlFHE2pZipYSyrQ5oOIulnxewxoxL1vKPHhuU
paxHO5yyJ/h5pCFTbzw9IYQUZUJu7Dwqmcte0QRitSU1ssEunvJP8rpkxPmOtedv
MW+lWg9q6ggbpOOkZ2/7Sgb/1wakvHaC+uwNTZjHI14wNFkf2jCFWkS1wSwpJZMn
RMxjhTOJRJoJjQFThiD3dvRSlTj7AR/29BIzSW0wqbrjXSKf8pt/0bYpxJdrbxU3
p8hUV/8zgmUtu0JU7bk8KvOyTB4XC4GOI8wbGs8if/crNG2qDlQ18vME4ag/irEH
fVM6fYm+jKfO9Du9mW4atsc2n2rZ+hEoqqXSIEoxhl4YRKfNp+KO0q/6uFzakdoR
IFBvCw4/bdNqftvLUh2ixvrAozujn128nwrHjr6jd/xUOaEMuhNXHHGj5MFxmtwI
3bCBdNYWU2FbNnEWyfx31djATSNU/EQDoThLy0yHSwcrDiwZu1pUFo/Cz9oG6K9b
32AfiylzUExbtNOxg6uCl50htR7D8UcXNcnwr1+i6o17V8ES3mzQwGUaQyGmZi7M
vCQe9vVVHtT02zQj/lSroG4V4lVseScW7+nTT2CBpvLrtUN/OSXlxxMAJgeUcLJ4
xQaAy03p+pGWKNn3sKqHX4uXqlfySFej5xbaJO2vhC+hPh3IYcp864U32GI77qh/
ktdL53cPtJ85k8b4drATcM8Cfxo+a+FJQh+fz+K5pUsSHe9/i8/HArZg0ZhWs4iq
hnL5NnWh7G2vO36ai3C7A89vkkJVCZXEeOLIbYiuCSRrNcQ7AMYULYN5UuCo6tEu
K1b6C6aCxMsa+6iFOdmUpVadDD4ly4oV+Iv04nLIFsyDqgNkWtZOlPp1Kpmui7VG
nYF8LzQk0pYa/uT82a5yQMBCGmethbDI7zH4VNhaw1Hh3tUFkjzT8TrGXgFy3Aj9
RC6YJMmdN1gFIm8hg63Q62ABGBs8aJUmFEEpbf8a9VM/gBH2YtMq0C1NhyarxPzG
70NtNVUSQmZn0z0PwErprhZutRgoQ/paUgwzu09YsAD3jUcxPQl7Oh+wzWV+ekpN
nIeNz4GhTjLGVKvifyDgy8ughNOJ9yzVBgFtFBzlzZCecszMQOrCEoTmXciINEVX
Scn5fu6UTm/U1aIKJDiTBI/RmFYO9E2uBygQgRPfHco2d7/HNaqSKJQwumQtjxep
lbIlmFSnRALYSmQyDUkCWA8ZwuZxpqZz2kC/W9N0RTUNeoVWr1p0EYAU085t/S24
J0Uc2QtHV+x6OWXOToEE7ovSpkvu05TmctLJbC6fsMg2bBAHLDWpEePeAdjc2/gF
l2YT9ccv58nQWygXQcwmi3JzpzOczklcRP4GYLNrHZj85lyWeUEIKbSwPnmhbF37
0j64NpbEf5kmk3hzssTp+QtCOsC9ptJt257eTSaAVNb0tvWAk90vsSAZtp4nYOLZ
1n6KUoN1eYjEEg5+2jDkhlhUR8WTzMxYJBtb9uZFMJkc08nWmhLFjGZYL8GRyN1U
DLXyFAPbIdnrI+LfaoqJauE7qPfu2oTK+1aUEw1LVYzSIMqe9CmmNNG7YecGHKUI
vTxsos7LR3pGxcJmcuduaz4R0TgHUiVAPMMO6f4uVt+8wUw03ddtWQjItkV2oXFP
W5b8zKdM4jSenlQlLcXafaKnJtRPlV2MPxpFgWXo+dcQRfW0oUyhSW8jEX6OGnLa
GlKV66RhEBPz9WqoBRM1Kbhb9KWeRpJqushU20J4FN6QZjc3USlBpqKKGqGZunKQ
+X1IKilmpaXVsFH+lnEvXZcnskQVcpUdlenjewPQUE7HY7zXsIOnA2ZQ8WxjpB4k
3wr1B9WncrpXpVoQyEONadI73tyW5cxgl5V+v5bJHereuHEtFjJzIbCwYaWl/nrs
GZ5baxcxrBq9eznT1QzXLYv4YYlYmeaZruDq+97wJJEPcrG6rke7/icQJNnDANuM
3ahtb5N/agaFhKGqR8tIj7zE7wafm+TpI2Su2FvUOaVJJu6NH3BB12NLdzHhAkqb
0lKxsp0+3qHUEdySXZ/HPTBbO5hkRCa2bV73Gp/0JSbUT3foyJuysLKwSByzShwV
d0v6NCfnrFsKs+TV2NTf0yUqMksFA+8Z6FRfObd6xew8FFGabDgidJrJl0fmSd5S
onN/ZbgtCqMEBLRSzcnqDz5k6oaRtyMP+H/nqSNOGt887vTPWA6A7AgqkUwvehi3
v6FiMINbeGYzTm10nV2JarpKLCz2QNLD9xhel4G8Mdhj+wv7/bLRYTw9ngTHFJhU
nzDNZBL6ORd+lMTxT0aQ3TCY/OhSaJqXuYLprkcpgrZ9/9Pq8rUsxo9v06ooap7F
uhIDmBCE8E08WO+/cxHwTxyUCyQZZSiPycqLM/gw1WUhgfviduH1WLcMF6yzrzbl
bDpEvOm3GYuXRgYZTmmUqZWmr0wmQjpOYr6HxFgrWweoCoRXtSRy3UD0D4wNzGVR
K0fWal2rLCLvVNKQWHmB5U8LsFoWJx4lQlMSBFg5O5hJvsssjqGDtHT0tTjmUJ+7
xs4sAlD0XHP4imX69C7FLKz1i//m2AoKrC55W2nDlJTqB6CcSq+x02xnxrEhEIQE
CfkUB5DR3W96DLcUtM5aThkAeqCT3DD+Cdoo82ByuE3GPT4sUeV3AcQjJB5hYQt9
8rgtK0fkXl2iGM8/Wel7ErsItAnOfPNjyO6VuSXZJgLdXxqKTy4UEXZK8+2qVk7n
/TCfMaoclzQqbaKkMBUaf18xh/0AZjf0ydjtmWJXxiMN74f2kV7lFH9wSW7qKenL
wn9GOhmMaObjgX0aAIsJIfm1ZevAcCnZjGkaRC+pzfYqfYcEh5Yd8Dkx9hVhnaB8
zEoJjcuyu2iJsjvXOGe0KxbZELPFHuaK0w2L1Tg8MlRarOSpB0FaePCBFSzFyX2t
+G1rv6qu+2pfDhsyvfyDtA+uMmP9bZOv91k3xQh8ITFeW8LuX5MB6VW+zJf1vyk9
sve8cKZBLuASajkK9BvH7jpNQlNfNf7P5gWtJAfelcZDDj6CC7kPjyDpJkovnmi2
ipGZfvZGBufl1/bFBdw1ptGKp5bWMEaPTETe9TRSSBVeQm5gZxI+kUn5cn7QET4k
Nxz2PzLtMWisLKWFtfmEhhlg86y+Q5rXVWgwKpz37iuzY9UTeIfFeuXiB+3Nm8Zw
OAOWUlSEHqYuL3107tkprfkFVlTt162gli9CflArbBDGqMHF4ueseHvR31mS00eG
dPL0EhAvhZEni+gJeS1PAqC5Ch5Nmz4c7MIZt35OpowlDDo12sC5iBN8E/g6CUdv
6DIsZYDslnoZM5tfB+MSv+Wa9cBHJLxg+h+aix7v21QT+ZgPf6JnB6o4UD6MAb+y
gJYqIfJfeXi6/yLm4BoJVoPSqXt73Xb2VgKQEhcTIx9+EnMvwgt73Ix07LmsJquB
YHQqzUgqmIIPdtS4N7yx4dlGpCffqIb2Nct3u1buXrm1mPVlN6VWItM53NtP4Pys
KRaIMHEhDzqxZY5PHD9CAzIlKfD3ticVOsWlZmNYmRIIRvOaDe2X7nMjgui/8Sqg
EJXwkhYNeCyEvGSij1BES8i0EqGuExz8oOMeFGpryNEoPiuk+l89HUAy5brpKFAU
8D8i6eNAR6lSZa1qsphc1nIe5ySGr5ojnc6VRtcvFx7Kjh5DdnEwkxy3sf+hERs/
oc4MEvQLoR/VZhiudRckqgGX7N2LRS8lDbyInKjppMaToV9rbCTq6KQ0WMoDECZS
9x2PYVW02MOkPrZo+MCrgcjKmHbp+iA4oyGfKff8NAieBtggKhDllBa4wdQiXrG1
MgwE07uZcSxGNuu4zQ6FQ6dDChXVc21+UQZUsNlRTGQhWhi633vlsbfHpZcUySMN
MGiIA/djd0ttFEYHMaR2Oj+WVc92hgPq6c/uyFP5fS1kFwZTfbynLjGEVDrMFIO3
nlhYrskpceEggApa/AYOGH2H78wVvkLTHLSA1WYsSpHiMrFDXtWtTlQIkNCzbKu9
falOVtX4iY8WmfJu+U/gJxe28bs1MCm46T++WApV/7RQB/+HtzIFzHcgbRSByuSr
UF/f9wNS1ducSnX5XWq70zA4potmWEWdLDvnzOMoIsKJDyLcQwLJ/1kAqJztQHvU
i5FuajK3N7Tn5uAJ0Wy3qh4mwzJ3DDhRyPy7GvbTJAvR+ipklV7pw8tWBAS2we9/
P0I2k5JuMprcOwBwWasrSnhh0XwwgBkrFh2IozN3l9UhN9n2UvRQwEPkOZoH1c3w
jo6Xn+qHF19kHBY2hyDvOmnKQ0gYXajh0WoZr03aVtDLLzvoHtqsblnRtPvNXu9+
XNbtu7Zp5jHBduj02q8klprbufmfEV1ajr4JVrcy/KE2VohvjStQPH2sP2qABkgK
+CXp+SJ/Op0FFe4coUqNjdVq7Q/Fdj+NF6GbytXrW5mCvtNgC1QVteiCZrV9wK3K
SmJUnC8lqOu5CVhc8IUDRGDOWGfNI7pJfjkYjzhLLANpxLMXE6DeQ5deNNCGNLKD
AZuuhJ9BzXBpCmWUSnlOWBT05xrt6Wen4mFuz1RS35per6Uv3oxmiL9EIJOlfC3O
+jCDwTdmWGhK4lyT5/HBJOei/pChIqFI9g78JpBV61yDBmmoU6UtdcJ3sAs2JrES
FJhx8zaSlYqe+w3vWJ0qnQvuG6kNGxTPHOynQJRUP48cEVzXJf7LhR631+KAx4M7
Pn+oO+R+k704tYen9mDuWlcZUmN5LXY6kz/JUB1b080RITXnucZrBJ9ZoDNMfsQ2
WVc6hLF6ZqrJUTnDof1PWjeWk+pptwcV3k0w7CMUDmxYOcAoCkm8r6zBaQdxq0XN
2I7XoZwHn6n6VfU2ZTmAm4+LwahUFKQk90XGunMzqe0ONnG9IeoOl72YCWnJ5Aar
xKFo1N1nwiYvWfjP9qdjCQplbAU+moLdg1ejQu4PJmKVZgXCOOG01xx2IEePS8sW
Gp2ZyvMlWhN2HeFBlTvVM5ws9fQw3xdhAU3usb6BC4GqFVUnBLDC4w7Q8ilMcxNQ
BzRv6WlXsN9eWM3TYyysc9EUznH4FQXBWwVUyiCC0Yerzuoti40CimZzX/ok5dQa
heiHHtt72Zt5isVsrmdqJb6YILURz/4Hu7NNKgQ6Rk8aCc7I6rrh1pQOjRsrSUn2
P+c+06gejg3TiB3hED0f3uVwvPgEXdajBH3MdtuDr/F6mL5So0DhpaTpi4DsBEoH
6NrvWfFNDvo97qA3USDNWW/O02yy896A1DtbhMRLrsoZHxXB8/jt6alWxjZakAo5
NzERxivQxHYZjuxd0ZeYqzq5ZTv9bhTmfaao+2EtJw7rSKy+rnpBchaIdumhdt+y
duh3mW8Rds3n59lYaXhdkF+RIbqHLfPH7cb9nkE7sBdb+5eZNKPx9tFcn3slwL7O
rq0bYqKEH23WVVIzisFyaAEGP/UGT46y+VatBO/AdvmNtq+33ejNfdgS7g7gPxFU
YSoSAWI13+NAajKHBr/LggHF/RoxaJ1STzKCkeiGIcZ+Z4Ww7oUh96T9iqG59OAt
87DrolVk9ngUE90GMr5xGDriyZNWpKZbXhmJMjKZq1NwS+wXRIU+4PT1sCzj4q+k
AxBjM5lSdnjk5V/nBzbAxmPzM5ZLNFbbwampHuo9QbFL/ZR/uH7wStSgQXeNKqOY
l+Edm3r1tQ2oVK6XsCfbfE9wPcNpaM3OX7LYgSe1aXYyUt/t0sLO7Iojd273k0tX
ESPIXj78iCvtHt12X3CS64SURq3d6nCcTzDmSQaMxJWNNxInAX81VBT0eu5Srukb
LvdlaaEWowswKBsFHLFItK4vlt51+PimXOix5H/g31JDXF1xcWTZQL3t4vWzhLyz
IHH/CTchxpSMUYObY5Gg0OQRAzWEH7XOqvKgs67btngDEKOwSWqKvqJ5gMm0R1tN
AeJSnStv4TK5CY23iiE4kjOqfnJKHHQtChmkWNJguxWJzqwWqg+AtfI2o2uiE88Y
TJyYekbsTUzMKF21I6KLO6+46o8MtyQsQq99MlT5h71rTabjiZnSoGsSUzOuisqA
PAJItC2E0hvY22e/mvS7lafK0sLboYuzg0czioHjixvuZ4wUvFfKdHPULt9+z1rC
1KCYdOxApuTfNWi25i/ceK0b5t7viZ/YEQ82nDNOj8RkcRn617lrrvsHAR7xQgAE
E7lCmBIp6GBPKOUO6PcONzSW0ppu8/26EGT6ui5RpWVgpLZARmE+qjX8FW2q+qIK
FL39knPVJxtiBV2ujP2e9ALAULpn+6SMteoUz6PXDqV/but12+xBmUbanxX3hWTK
F1BOaRNzYrI6rAmqsXjJ1OwsgQJ+bH384vrIcZMiDVAmR2XmL47mBp9eXmaTWdAl
xu1XTPOoxEU2Cy/AzBnNuQwgUaafn3DVeZ+GBrYhGkZvHByV5jfQE/Hnh3FCOZso
Xkwjg+X0EJ6b54QF4Ea72C9aGFGKl6LYMiHBsdYdstk+yFX18zYshriblfg5d4lb
NOQ5F/wPqjQx6BaMQHgUCEJSpglVIZLvRFABk2XjRkYnmGOjPMtXJACykSd5P/Cw
F9/LIZiCzdsOlU4LHzaY8mX3P3IiN3IS+fegXVJxNwRvMHYIw2Ok9ptkCuVLpDuA
GUy1ObzwXemwNfaiaInWHLRsEJo91BqnD2n5cd/SOvvx2x02zs0EzfITkUMC6zFF
G7b7IC9PHJom5HWgAg+Qcu2iX57ItWJYpxThwdKehPVhoNGxkEuxSWhY+YcZg1hv
u9gI00zcxzJWNMmSSpUwzNn0UH2RqjpMlj5vv9Nx+LfLdxciEtqQsLB+OCOlcpl/
ZaulZJmbeEQFNrWHCHvAcEQvbpJxiAsC1lVK7qDRfLuOKIzuCg4/mVS6k5jbVd/l
XztXHc401xXrz5B8XIpZZ+wBzOjGxZk9iIduIg4X3zSPgWX6XVxgF2Krt5TAdfKn
1BRwaYDrM+5OCa2xh9VIfzUqCXYlBL/cROfZ8JQNtjSBpGzFAzr1ZVsrRImE127x
E7n4KqN/p4ufFZbiNFf0TPFUXlV+Olknei4rpfWHsuD1v2Em3NoHzUVR0eNZR8Qw
KUMgfofH1OJh3Z/+Shc6tjthKWbDR9AzEO3+k+uHnRGs3t1Fx4iyM+w6YnkbWIb2
Lp32G867gBuQQgv5wL0MCc0faL9UcIhL73+xjM3tTttZlSUNTje5Yj6t40LVvQXq
uQ3lTdS5b1unkj6351Rh9N9dwOzhl7JWvbKOpot92KyXR9c+gIPVpevmuBrjfNVG
p/C/r+FGdTtf9kFF4tlkAI5WQPAH1CK79oOl20v0CKlDJfrczYA4hWzGjgpVepfv
tl22o6SBcEb1MmbFF8DQ1NIG+QPM/EH0a29SqI0J7a9eHOGRMhrPK2j7J2Df9YtV
w7iCd12OhQlXh9dXnpEcNdDzE3ryp+h8gr+0VhGgHJC9KcjUGPEklncQFc8J3aaL
td2/aK79sh0dOJZnSNRAQzRHW+KtPkgYU56S30Fg9yy9UGOUI+lIcBwzqDwKFMQB
DiQdJIVfZe/TaMx3U+16fez2HhGviu5plOe6smhAbb6m9zm6EXTC03BbCMTmMDdB
NSCm2Httpp+AEZ1bdgAyMRqjuCtqoXNq/NwWHcdEv3Zg0D0t1EIlR+zBGD+JcuAc
TXqp4PWYk4rJLNuKs3OxSd/W8bNfaGvoEBeZUWMdNXv3MKmOF6hvMOr8DXDkmeIR
uIibONHpp+3IK7LEgn6f6SzPiosSkQvT/j1j34tj9Y2Fdb6KTtPGsAgob4I7vLAq
68G6DOxExMg++xK6sDcSLeeHeLb4LAFC4icmkWTpM1lsTc4V8EZFdg+Dq0VXr8WR
QOz7TiRUkO9sVHeIxvoQrZLKg3O5e3LhIBpIc7aAHrwVOk0ZmViAnh4dKiiWyuFu
ZMhOPeW/td2/Fnrndnh8vld4BoiXNkaOPOQsGJUBtpAyD236XeeRHzvv/U0qop+v
Z+vxEtLWSgERpW3NXMizjIfHA8mFg3Lz4SYx9TcGTttKWprjvzfxjLepN8xgZ19F
aEa7WwHlZ7W59KcZNSfOZGuhBXv1VM06dwSSltEY9lMkv5mSaU1vvoxcq/e79h9T
ewdT0VHxNlbBYPWZT4lOLi9GwcTRXMBpvHdCBtf93mqhBoDxImtxUHWxHZptGp1A
qimRu+ZJM8Lj3vTqZVwoMRK2FWsk1VCNhYOmb8/Hdi3B42cBp/LdJBO9YIELYYLf
m1a9vgaoMAj8qXyvTIvddet4+7c7P9B+d5S+3uJEn0AR4j1PsZg6zf/cUJWDOT6I
TYbMUT+MlBWypGpQdUjYLpzzt/kEPvTECvay1vFp1yU5XDytzvRJz0VAuwcYWQJN
jOAiItzX18yAkI6yRoouADcGIJGkY5G8klVoJDjU21Hb+LMZczAKdJedM7rph5Hs
KB0EltJ0/RJ2lpdWgewokSPBRQAt+b5WrjPcrCkrsqfVjVwPCQRQpUVu9iju5kK4
2o8ZA99uI6Hy+RyYgCXjivuFgpOG2hNZu4l/Fzw/ILfDRKZySg0/iA5MoJ/XxRzQ
7B2ym4/9s//5nh3ThZMr5XVlo2LcijFmp2P1TotMg91NSpk5VLCbRRdoZ53m6fQd
8mpOx4cZw0Cg4LosSqxWoOHbm9645+OziEnwsqpCe8fZQvqwWJOpJGXmmvWszRoo
qfHe+2RUPEEEEf4MKLiX+meVgdeHKRuWj1wSwOelwTtEM5Atuns9C4rpWj9gzZ6g
AZ7qwDlEk5Mcl9Ea6Qk65md3XwafKb+pq4DZaMi8OCLFurohAl0DbV9GBeJ6baXs
noqikx7JdReQWbO5wlOQLE3o722dcsYMOlCceAefVP5eKogfJwPxmA1skuvvBFme
0Z16xrZNJ5bXrQPqT/88+xmQ/tEL1DLFM07zW6HcY+rpQxjKyJg8hXSq8aefa8VY
I8BP59KNDla2l/uCCHmUXyy22o4wM06gcgQE8qZP0jbs+wjXKVg3CzRRR7Nxmx7j
wyGbG/tzCb/EOP8Fc/PjLF/1XsVIcdSHBo2BAAXOy7G14/xLuG1G1imDWPQ8Muod
h62BeaGx+9/bSHQZZHS2uWuJpCSRbRKWDyFVqz3L61C8hrc+KWLmF3otATcLI7+A
KEbdzcNAsRSLNlSFL6xLmVJjIM2/xZRSHTyLwxw0A4TM+m+KyFhfHlB9WEnl6CBr
79gCN8yyzAQkxTXppFKqIu8wcgQ9be8BSJ6kiiN6L+kzMa0JvyclGemJ3i7Zt0xZ
su+gRO9Zw+wdpOsiPK8q7yREq3+cQ/VcF8cc7vpwbZdgvLDycyAOOxWijwsvH1/v
Kzc7eNqChayuQbAyKSHwkaInMnNtQrS92fl9fxWH+rcvoFs3pYrloHtFrIVKbWC7
JhK24K4DrJGTw8w5aoDXyEFoSnVc367kMVy4YvvOrDoGrVxbJLhWcXxlqdKN54ED
CUFoQHJd8PRI6+Bd7aEU4sjLKlnoHQDug5TVpQHJwTQep+K8xBMGTGBBvWG/SoO9
HEifZLb9alZ71r1edbaAIDQkAZkmJfN/tg//V8jOQOQE6QLDqX++BUMeQs0qVjEg
kP05lyeR5RakqVRgaz5KnWPCH4xnM0JBt3Fel01TLYpm2QYUgqSVWosHWONF9o3l
rbOG1ovm1qb6I4o01ZNiVkdRGoNh2mllwdkSE3AKTUwvSAZ9FhZWDgds4zQIQmD0
wO5Fu9xH6UvxNu+x9PhvG00CdwP5xzY/s3ukz/JH7wjl2MYzt5O4tALGbftE49QX
rIC7WB24Xs81RWGWiJIi29kbKFuXsURYBm9Gr2awvGh/EadmOhDRHgiZTgr0X9nI
42XxQMvco3RDG3ipf8CTUyKuLU76vp/tjZrBz4+l0quO/BiNQIDB2rMjqFPiLVQB
F0H4vHM7vzylwvvTb6B6G/M2tRlRYyNdBBFLG+RS/b0W0dyhnlvAH0tF/P/TK1qT
UjBSTQu3s8YOk5X2C2BqQTDRKczr/9x69UDmLLye3R3gTIzUERS9LYaf2n48ywVx
IcfJLdFtfWQNwslAQQAjh8oNk7Bks7xZuiJX4MzMFPm88kt4SGJ5nT5YAG5yvPPU
BMQeAPI+6W6tZLmSZn11OU9n8vHa9GRU974o7kwLpuiKiQhdIxLsOiwvusXeRPF5
f++RjwN2Hgslq8TSCfLYzcDvQ6V8UZ9Uz8HWkQZqBx3Mu4S1T1qtmd937A5Ut30s
tZSVWPrReB+26J8gDL7VH5lbqdcclIArox3eKqqcWBKZdPqL5ptgq3G7m3593NW9
/mn1OUuHGX3pPzfeQXowt22gm7r8U/a6YiBtGy/hBTLdkM4XdNxSqXPuA1otwlGe
zM+mEvRhMaWImtBgrcLfzbQoTja8jRWbFgEn7NuT4UvDBuQpKKFfqnOgOZi8qcNK
0XDbrTnxFtR0M05D6TEiiY5Fu8fI3xr2it2rdpnM+Z24EQ1ZisWSbt0VdBEGdunG
DQXGt9zoP5cYb20JfrCoH1nk+a5OuXZDJ/Ozxq81DAMMWGSLcs2FeU39k0wLlsHD
QFuumZwgbRnlEx4s8dB6IRqC8HUpaVjaXsM0SGUC4BkTn3249nf6U9pBJa/PKIP1
EgIxOSg38fiX2+wD33Ae0/VQ+oHnBxd7iPxwTBcnJFlIR9fbhvEdQgwL0gh977Os
6ReIIueF91iA7gAhxH+Wd1A+lQJlJapLmP6CrwmlAJEQSwU3s1AG04xbbT8XxXRr
2dwJlp+6Uy1p+a/wj///f9rYxIheceU47A5zWeOwXiF9JA8GRu4m081qE6EDTEhi
t2qwe07TKCWj8CZ/T+SjEG79LT0zW2PYC6C+/5ApA8Rs2EfmBq6PWHykuWeHC16D
TZtbwo8RXAt2EDCkIayZK41cobueIAgGv5Q8/ka1c5/D6kVgZMaccAgfwTZxuEIs
d8Mln0GOFSr3TC0fyswsXX0f6FY9Lh7SeE7ouy2SCunVpE5hWn4QmEi7QHKOwlzO
7+NFmGQkot1rKoUzW1s/62+M6AvzI8S532m4QymV2BFzBJeXE+amNr40/3klxVQY
AygQCxdhl8afhHGS9P/w64xljrYX8ao3ponbDVZatFqECP5lGGDGb/n94AGxxF+h
a0x6HiM860PeEpx5SG4iYVjjGp7eqWFmOA1M5E25rZZWR+AgZT7s0FyccbiXHMHc
R/F7H2ihxVE1cBab26JNgIcv/J4qyCKhmPCcgJEjTD5Ea2IfN7kh4VQAYXsKQi26
FD6Vs414owv2FixXkXBP7HYNRQ0zYr9x12mY9eltbFRvzGCWRtoVhKsmHxQHpa1P
pmbcr2xjrPj5kS6axSkhvrFYB8lK/X38OYAqkDKBamT4aeSyJSTmraATG5b/WQpC
eWKg5amLz/hF+TTmbMUjpFTvRtfEja41B/qc9CRYc4sgidw1NlU3IFJUqS8U6+1A
fhtkqDafpT1mkCYAPkdeWn9WP6V9RB3hGuWP9eJbzDHxqTIEw/CvjyuYQ0DYd/4c
rxQ3dU19AaNEpl1Cy1vb/1hK3tX4iX9tcMPFka5QEyHOB5+441oXjmQFe3YclBkV
62vYQvTaAjnnS04pQkjWDE5YAFdMlR/2OzRtW30zthhRFijuQucPzidRnGPfOzLb
sWFYCIDTP8Gf4+sHeuLdIHM/+0cSQfe11+h83fMkc0hThJ8fWfIMYPYsvqrFZr7b
gWA655X/HZUBKCxa9MmeFMftLB/BHFVz8eHmLcSLublhRod7bjLp/3Hz5B19dTux
0BTiAovFNiFUT7TN8E1dVNf8FoFnOqni1ULKjk82naST4pWekLA+MDgZYaA/0jK8
yesxuytfElS8zbIlYJ14vn/UeumoO6AxzygN/x93qjFgMvXBspRkmeqeRgSQ2Jel
aeqbojrmd4qWz88E9D5fApkTewzno9s6VpZC1YJ5RhZgcMMYCybVNEBZPmQrVRsz
FxRHyi6uPWGevIOhYQJ37sbWkX2Ha6cckThICj1Bm5O6OxmFCaxAcfcjp3uqBlG4
O5h/1G2clbUTM/TTqE7ZfBaj+4o9Jq2JWJFVd/hZaMpGQoKwrVyeVcyFYBXaB1ST
cMLhZDAl+D+4Y14BAjsxt5f8uuTiIxMPXmq34jQ+z4mwM64ZoLp6BtXH6wIngO9o
6Hr+qDjM6HRYc4voteRadnlsgMccjCa+VwyslvqXkL+FtXmU6w4QR3AgvNnyCPZJ
FLbM1uQALkluuG3okpo/rdmbKhmFzOvgSnlCljfjTQZmmNFdDislJNbDJ6BJsbT+
8cQfuKDMhgHu9GW3od/MT0KWYxd0otbH2QStPnCve42HhmFM3ZCmANVwRewj6uy0
+wZIzhQY5kqJXMV3kmLz0IyZkEeCX9ytMC+KAoQe7IZlwxScjQaqu6bjmNco1atz
N8/DvQ7Dt23EaLn9DOx54P1mLMEKyJGPYHI5p/3WGjQX3C8nOsd7vU08U9qp7EXl
QkepjuxADZvVrRuosSdHmdGDAtRdxqQ2S9LC0NwPIDa3G8PKUb+J717FH12F3lP5
xCSEt8UAFelZxA5g87VPj6dYbQ/JzFbkM8cCbkmlPc/YU+gUCFd2dNClu9/trH9o
AhFECFAmpEmGRMXJn9uaFE0XAoHitDAcbSUH6UURPooiigvqbPAxgw3VSyaa0CGK
drjsh6Xvc66fdHqDhI2Kf6WAk9wASWwvflwkK7GHfIrs4GLqgE5ReOVubvKSuR1o
fadGvXJLYhtnD116ZV56j/Vfmy+fulXXGlczOgE6cIFPzBxErPQbmLArqubUXWq8
B2VV6WXp1IAiPEEGpu78bJABKEpjWotlCmzha0UyKhXufjqhWXLDIij6WijszqI5
XK6/NismPxVvGPIx3mIWxFTZaNmWAGt3rnsV+2KbNNqbgiJeaqBnORHHOzaY2yb4
gfVxOSbOya7AjrFyAA2i6NQ+5DiyuqQ+Xarq7E4zisV+g5fR7cSYH/gvurMACKi1
eq7fIZpz2NmOkilTy/3N9lry0G8Cps22F+f9m7C2c3ZucAOTlRGKqhqlwhb8sgj+
wZlc2pmL73WevVYAC8baPkQwv7He15Hxx6Xp9D2XDqr+IEWF2syRYw7omLhnF/yS
+3jrfFnFcVDvl0aXgUhq7IcsEi1UJwdWPwTY3pniAP2WqneGfJeXgUm1282GNWdb
Xj5Hfel9BdtZYEyB8KQ3h6sj4gAaVqVEF3jJtc6F/wgWJl0VQN2eG6ioHZiuJ6h0
x6WWj55uJhhvnraiiavY1kXwshK+t6Oyu5XlxmR586JKMpUVIhGLpO0nBv7tT0Yx
P/KZkplVbxDjYgl5iF5c5s866t3iJuwNoyzpxB/4l3PMwz6Mu8amx2nwuWwPXB79
dKWQ8gmENEnbYYXzxmzBuEN5b40OT6djdXZMVqNVrTTal2l1Sy8SW5RHc5QV9AWt
7JAgKqOCgmtwArsir7sScRh8L0fqLmw8oL5eGiM5JMDBBOf5CDH1SAhqs/mlgyA6
pL22wrZ8cWwgiIMHPXxkgU4dRPERBoh+8rLyKLiLB/xMr2zHGHDh4ib/hr0x2oKY
wDReG1xbN32k2FrAFhVKWx7HcS9OeCdxPXjd2tGlggZwRclVY2Ffinm32ubZeEke
zSdwOIkGVJw7atxsFfVLaPsAq0M7rhnG2g0fMmHvDCucnaiVTtJwWWzmpxrXAYpm
NbgYOv80WslcUPQVu2opQoUczq2DOCUc8HqHPiHYrucfValkVecdzbQ8PZPuLdIq
E4rGNyj7rX7Rm84IW02hyxBznYOmIVOXM4jIwqc5SMtcjbnvodiUR2lr5yCj+JWm
rzIkKpUOq11ISdIdbuRSukjj2cEAhIUDXTDfQHOmPw5bAQcv83qlgVspmq0iR+wu
pw4N3RiXFUQGNyWxFOmBJJqdo4kxQQQaGzJWCXoDlkeJxwopGMzfts9TU40u58x8
fUhOoYENJ9B+oNbL2Dd4nQDnBshVLmUr2hz2n4UU7DXJpszyz2Rb+afVhtk8Ztqq
tX159lgeW5xa7lBATDyRbBK1IPWsxyeiOQVbNl2f2FTfJZdF/WH5cyyalwKPicwo
BlbEHEH/9iW8/Ir/tqRGpR3p3fpHveYAX2ibEc75k4Qy0UzpDuuwTN3d9ghIRILl
Nql89m4JHpDwLgiG1QBj8BGx7aNy64cfn5DuADwR4khtZCmVstPv6X51YjqyERD+
51ODC0toMUpjPWaofoTBRZ99IqkBS3MOtKKr0VIa2e/TGlMWwHancAGax/PWd9dg
fXUhc5Ixw1X6GeZ5ubefdudCec/4cL/5gC2QcRGk/XRzG5NtonA6RSi+alWkeOG8
vdugg6BEo52urGWMsMgaDiZyunRsZUffFLdAiZNdxUwwUPlsUyOIEAjDxq7mmO8S
RHJVMWZ5nYvM8u/Kq5IjyF0LIMNoeUkDA0pMEuKUjjiykKtrDStDIfaQrhT6Pt4t
1UoV4UhWZbr7C9FOUBXPrW+osT20mo0Rjc/PQH4Mgvae0JXajbgSMRSRKZGBoSv0
Nr9BwZCcr5mYIg6+xfKyBqjMxPJDt84Bmc7fozW4A6Cj7UjBEBTG+M2llQCJzM7t
5IAoU2nzh9ivQkgKTyxrTWz4Z4mQhCbqaH0rHCLaSPhOoAo2iskT/7My8qrVVfpt
hAFvpSn/ISSty9ltee+AvM0uoD03+HbbDE+p+V3S6BIecDrj6dgMt55R9oFDgG/Q
XeOjn86rvcpyHzzWFmO9f5o0bCfuZs2UL6ytO/Vo0fm/nNoLd3Wb/v9Hdr6gh08E
1H1vcCwlzi1VV9zNA9xeCD14pqzP1uNmt3otvrsFoOiyzVW1n9xFnpYTymMthfLM
W+mvJcLeznx+qpsO3t7IhjUTvtQ2cqp7ulOiwb0r1gTGYkwlNcYMlhsfdCzUlcX8
lgPGKMQfyqt5wd4V/O3eQIejszYfvwlCnyslGF7kwVJP1rlGBBQxVMaNk7NOSLM+
qokGzi4+KI8NoIkNsz5IBn8E9WehFz4hbKX5/c1hUvEZfoA+EWi6SPdTYrY+0cKo
N8j/UABVo7mJhB3qD5SqIYzCqqhKhuUEM3vFneOKsE+JmU5MuwY/rvej4R2zTkFW
fh+Q0JOyYcbljEOYM5UR9GIGu18MmmRLcLi88Mx1rYvAMpdz9EjRXw/SYuNo59/p
CtkCDktDfMSBFM3iI3PmQoPa2uZy/vPGUq2FmgRQOC+3dbSf2erg9/IqtYNpjnTW
DXeqoRwGR7oScKQP8G+Q5+Kq8d1DQPeGpHHUHqCEH0tVLP9HKzDtwbEGF+XRI1Ee
HcR1vEgpx73MaMP7VoJsveehMoK/5d6XbHhoowQxLQs0PajE7TPipY5ODmSQfyxA
9rJtp9QouqtQ/t6Ygmc1HOEj9rYz5/Oip4FEmHJlqkVpZUerQQNrMDIHvGI1wpXg
LE7J94Tg5pcUoZ3irXg6BsR1SdF4XCWfNNBeuM3KSNFYydu1Kqo0PUWlRZ2OpV2j
k6rMgjd/Wvj9/JGfslE8KINS9isE4wAYdQvxCfS/u7Ky1InVJExvpuT1rZT8OSST
i1Bo4TmLs8O0uOz3SkSYpbvScXNeJdDuQTlkiPfSLhEAbaWLGE7BJ8OvcoDmUhr8
4Ew3L0TUylspSppyv7PFfCqhYodB9b9SfOqJc2BuLsU1s0C8rHf79PXyFmuD6YuT
CSaaQi8lBfLEUN2C0SrJNVrqgYzIRVYJImTjFY/Kd7T4LN7hbeXFK+jHTjjtkpXK
qt/j4nU2bHNKGWRWQ7Em6lfK0r7789UdF4WqLX87EQjJqFkXK0A/RKu2gM0V42m+
qYg9NJtlDladaCQKGORH3Q5DVAy6lEryUf3FLgJSMyRt0x26Q9HFJwVq/dx6Dvmq
HXQFH4Z0ik7IEIxvSRx0dJtOyrNJDAsifipn8+yGfqJgaDskLdj0UH0p8aqxkEUX
x9g5Fi58pFveZk3B/qUuXPa3Dcggvazg+acfPpmqbi7UK1rIQcmVj3nR6e/ZzCHS
g6O1BxusNdHhaXdirFSo/xijNbquuj7Z+Gbh+691WCqr/6ujzZa8m60iFTZtd6N1
XatcSav9q6f4KJsGof4eskXq0egShqTMaRKptWGO88gJKy/1QmDl4JmU/jAYJGfG
BAM/ljoC1HsWTFuafNn2PmUUQH6lJ56m5+Sr9IvN8tGyd+XldLejfWQ+PfzcUJLs
va/Di1E0kCnk41v50Q5QU3AMPXInCEEiP28a37pTDuFZP4DxbBwFoysiVxLcO3YM
UKiZVL2AAbHGH6pADY0K/GU5Kmvw8Fvc+QXlidWwsDytzlE7cXQOI+umXYdDWDkQ
FVvlF4M/WO5LAF4Yet/KXOBmBad8T8cad+oFzP+jz79YGkNjd0krszZOJdNW22mb
9cHxvkyL65NmxNZBG8zqWU3hdb2dXDlZs+GxVZNWS2seDaVjN2yX8a27rCg2HYDA
6Zy9wGXKA4r4rR6bwW93VgkLMRaHeZh56ciSzp8weIzbBABgGEMG2tKL7+p4rPrE
9fO5JnRIGMAFJikQ3t7DQr5fu3W4rGoH1of7ITtCnMPDp1Ect7ViRhH8FQVxA2Ft
UwSBjb7SYRDk/+rY4puJyNsNQ+0tkXAzPJwx/rdzixlgy+GBhQdTuPVvnSteZJyN
m6KvTho+4L8D4NGTJP7S0Gig68UboO+qqNd1Mzr6JY5xVa8g1pvCo98HEo+sN1lp
NnKGdBTkgeyDSt9faY2WQrIol6szZ2ZVfKHHUY9Q+mX4IaFTPLgmXWGkayZTCo72
v8IOhaUqVUTNG2agCvDTBt6sM1sbbe+oF/3C7etmj0CzTcQXB1HM+ou+cHOetDGC
g4tyNKBFdfUsA8P46ggOeB+e0lhHs+GsrIikts/V47ZLcYAx3eHh3Vfe61X3lCmE
xqiY0+zyp7e0VCtF+UImxIbMmsj8Z0lh7XoOWcUZ4gkbznxneCd3NQPIyAwtK/FB
6gWlQ2nnMDf03+YyW4qL5MtEJmKfNLqCip/xGabpaNPGFhcC6lumo+dbJycAPU9x
3CBTQVNmwhkVw14YLGPA9hI4HIXKLQjzFfdsTCHwkUFTfog1bw4Lgg8ms2g0FdSz
EGZx5xBqd39frjmWDwyFo41yxOlrwP2yE8fFR02wXqFcWtn3pF14doxK3f7oIvkc
TDym0mGWSLjQRLYmn2AwyLOhmuCV/D31owQsn6FHt9RYP317hLtoxxQWpVteKWTW
UGhE0P/RN/VgBRbMLuciBXRhcpZPre7pMYsI/FleKNzSYWEBJZuJoh8ubwXE8lwU
c9XwnbGIwGAXEvVM9yFXoICE1eifYVeACzPl7rcpgzv6tRmDnnilFGiTuniJkGAz
0xIS3LhHLAThaXe3F1hDjvT/CmQHXfIr/xfDrpV4gFoMt1wq7snJ53nFhC4TCAz3
EPchXddkHEKW6LnjV575hNXd2Q40wAFDu0Rr0FQ64m+CdRW8b9dyogF/Yi1c3e1p
I6KS608f3KBudzQwdrpnspUUeBWRoV0uRYRC5zXci4ElB4wmEkJv8PfIiT9Q4SYK
vfWmTffqK9Kg+gxRhmXSEOdJdtM9XoAWySnnzJW6zt33qH5RAtNHv64DYRbMkqY3
HA4H53xwncKpO4kOI/7rNdymVyvPDEw8Z7Ex3eHA6GdkSkHIZsjw56Cvy7otdXUP
BUb6op6wUV61vW8OnrYF7MEWwGsjFGfymj+WcoEglBaX5ucL0mDGJ7fv8MGxS0SP
DeoTOUtKVvjSRGs0klLllDgfrTM03ycN5zalGbsAXJFBNvdMC8OaPvPIppTr+RYL
Tdv/Fpi3vDtz2LJMDDRNgVZJp62codr59vQS69WlNuX4hhkcSh9SLPfhESsePEyw
pHvo/4GnINA22GvVoMQlFVH74yEiEZ+f94X37uzYVd774Il+oi45iJ7Itf81M8zB
oK6yqnl6i5zQjllzisnMJRyZzAgcEmthGzGT9H1AeXWobWWb9CH7akveE2uOH8e+
hfGAIZ4KnAIGxYZujIqH//Z6L/Wh1rpxv8AoqO7hnHs0iwgPVrVFW+m9R953g+C3
7xemcqYHNoNVsR31C99Dwkse1W6eQNcF60IxDKmDaiES6FSlkg+BNR0Fw+ApqoGq
AWEuQ/6+/vMYrviOvOn1L95/sSG7YTqqMXmr6mFSl87blJ8BfE1SdhlCNEO0fWcV
2csIGUh6DrS4EpjwAR7muxnJMJF6am9Ooi7gebf2EF7tAjjSIfLZ7TzxYbjKdjp6
8RmAwhrBbIwxMYK/a5nodMV5OZxi9Oa0p/I18VwLmf5D4YqImfSsu8C60sdTR8T3
5xrBu1R7EEXIr3vH3iLPTSsQ83/PzIXtIpWKMhaa8EjvMVqcR2i1b0Eb6OFkBmpR
AXM2Tn1900v8g/nFbFxmzuyCLJFISIhxE0itQ8IbSOh46Ul7quzfe8jlYuVSmmDb
ssKGjqFO+nEsHgvjSFp7VOTGTbkucmHGKdRcxPvJELFBUFphgGalz19gNGCqE9r3
kLmkdxlw1pNHmWb/2bSQwwEIGdIjkxW2L/leWoSWhM7Ge3tRiwLuMIjPIz3iVDUS
c+yIXBdkfuCX8q7nyOdtXeZOf1UWIPRMgJ40HM+02FClbIDm1ETyV77MEWKb8EJP
+pW3ua2+oWHsmRNPMl8gs60yj0jfHwPLhsNnv+8UkjBFuvljCJn1/i485Xqa0Msy
HoWqt5Ucq+KpMfLhRKB7cJ1yaFHb3HP0wmF5myb5jFdRFWVgtdaRtETxak7MpA+u
aR2KFpnHCyBSmq9juKq24C1F3Uqd/M1ywTgRLgRnu/yAMbI3rXbD4DKLtaTJ/Vfk
HyP/moVv/GXUShmR3pzan4FwERZLvkWxAXBkq6YvryRTAlFnuZaMveTdXi4j5WwV
QPlPCKUJjv+SgpMGRSymWtwKmBLpPow1seGEE/Z4hChOCJ9yXiwLnZzb1leqlGhD
5ynO6s1lhm3EAtZrFjwNduBRBkmNyr7d215ZLDyDkkt4Yk4A2AeOeS2dnXgj0bqn
3wQszBp5P91wX1WGz+fYN329c8t4DDIFlIf0BOYkVmUDystq2sPfIDqnCthNGjer
Ja97il4oRaa1xzsZPzjKh7IdMCGK8LgTz5YpuOsi2eYqsdhrInDN9miiFzKsfxlz
1+iTeP3vozP/HeNwsGCTZJgGUqkDWkJk2u02eKDKZmt3eU4B+SFm0DfeEXGrAQtS
hZMCfdtWKbSMvSwI4CM2argBy/o88GpYvFqMUbuRb/YkvNjhYfT/ce8EMaAaTrWz
bISYRV+NCdb6bGE6csbAyFb4xDBJqU764rRTsJHnBxbpbXE3Is44yf8zETqIK2KG
/wkh8627itZ9gATTy1vy0FPVb4F706GmwteXVP7jubUp4YBp0vU60pnBzljAi1Cu
j9EnjIBcG+XumtmSc2a4o9NUgC2p+fWMGfSBcYO9RqiNZXL/nvXNOnovFOGqR6pd
1lzJ7Y+NW0X+BUkF6pLKGWKPGqe8gjF2iwt5qBhyimTdR6qQBLU4SRwGi0RyrxA4
9NdtzVThqyJr05Z5A+/alLbDPy/qxlqsH1Q5qLyPwZ4Uf1/tCZ5eVNLHuGwzle2Q
+lrz+wdH0BbmNLdp0uUfTHNWMh7W+LPjvjBGNCYBYoz5FuUNX0HaJjKYrXlmcxQ1
tBx364a/mBhDiJAh/beXKEmbCfXKljWzCKMUDf44dw7gnt14IGPe049RKYTNf1TN
pUgTc8xk40+N1fVXOXnPguZBYb4QSd/lr2/50EZvEVocmOxrGLt4IKaH/Dj1kuLe
Uew0Xomv4fccYgLrP0HpfWyIt92Am9Ryope7gWnzsO+z4quhOkvY4EjcncC5FBo4
KxgFTuYWvYPBad9eUm1j8rU4JoJy62i8M21Kl5dNI3gG8uVd9dTnGE5hrNfbsQO3
pVvrLeJBHEyYA71r2HDX/T7dLBEIrtlZA5ZJVhu4KLldhaM7hWF24/m531/vMcQm
Bh0f2JuI3bXiPwOF+xTae6VX7YFDxx6Z1aP/U+gWv2qncPVDixs5dQ9St1eT5Oo/
p/CaRz7tLwJtUn6Nq5hsxjqfctDjQVMEdm4IKtm2+DDEs5l92XcNryNdIwYfwC7M
+d9mRSsqkcjjHFZYONHm0KlsJe0fHcL6f8XBqRyvfLy5W7hoG5ByU4PcWHgh+p5A
A0cBZ0RqxBh1w6Dw2HgBxUcxcOw8Gx0js8UYftZCD0Pbqy87OofDXifvHwS5l0lm
cmBcTSFleBkbmMOXwvgnmR3DW6ndp+QU0Q6u+5bVTyZTgM4YxDSWOlTImbIWkdEq
h+vcmKSCrnQTDOe+87cddzb8I046VdJ2JaGUKeNobdFJIfjl/fHgkQe7yrj34Yvn
GUqEutjplYyGWO7ErA5ApInzxuqwlPBPYtg1xpuwicIeOCvYY9GTaNB49H3OabM/
3CkWz5WUdG4zviudFo2OhKdN0RJnjm8UcEBD10BGhIR+fg7rOwu+adKshjmvOwig
ul3lMHfraV7qb5R76j4laGE1UMIICybaEDhrbVFVFQUdtvzZgHm3niY0Go0CUqpM
RBb+rrjgGvTMy8cT7Pt7TJ8r5IzgNaTQwiSlUri1SseS0iPtNIKEVFS96qgHkrof
G22ebWFVDmZx4Wvw7/GS3InPMMgjllTEtIjN2Cb8jAevbi3gR3Vqj6ESXfp6OBHN
nojBDglGUWlJKw4rH6fg3Rf5aqMaP5Dq6GdNcFssFg0zWc1bCA2xnf5SfkufwFtc
R3q2EuYCqsKeyR7Uxooyf7ebvAf5bxPnbvDDp3Ai3Pc458SIXBHvaXAlQoJYd6l7
zpXOFiFXUmjq712Gn1YiMKIGYsCnE++d+wA9RpD5cbxSoWNnO43dOQxpvJx+4Fsp
gMyvfLToGh/yDTg4YX1NsEegDun1oz4tvZBUHSJzw5g3ePW8zgyAHK0/kckCc151
D2nowudF1mdd5ucmawTQ/M4Pk1rSLibcjPGiRsHCNT9/2bCfEpeE5Gogt2eIN4al
FBH3Big7+dxHFehj/lOvoFx1F+McN20FAURWziIRv6FuuQNX2OmYWl7lAgBx1e2m
LQcHQy200eK/E+9FnsO4neyuzieruQKlRpsDlKd3fawL7TckwIeX6wUbEYRl1qkE
0V76NMQN9xvCzPqvD52U2bXUlahGOtZUssuvD3VsstSGp166MKxvzcifooqQddJX
l4VdDp9M+smfJ7/6k4LYQgHtgluHTf3HF3/94r4LOBzrkDdwXrRpEK/EcluM+v/l
IIps3ck8a4SQ3oKsaTOBXGHLV8stbOfCElLVE7hM0PDY6rLrutjqwNI1EtVrBGkF
2pi2D1TReLY7JpTW5NxWw51HFOmbi3d8z+EpE7oGoGpUAganxhbj8CeTNSMHO0RK
ZNiGRNwmQ+qLG8tpPrzkxeWWPSmlK4um9FCagpgbOd7s/+OxPooP+EHd8YrGpXmP
+vrPSBgKHHDFDWKlGNwX2OzvCMvjTHpGHcQJXJn93DzLUK7i9txcyLjYG/h7DHcK
HEx+Pg48/bkhX6jKzoaFrLKpiExFSiu9FLbgepxVQrTAQwmRU17HEdPvPgI/dclB
LTeW8zRPAL+WP4TCPR0eUbQtFOqCu+QFpPGyBl8l/dYCfMUgSlzyKTGoGuZRGmXk
Q8rlUDyDXEXR8lNzjhzCuNpFKzINbwFAYoETWjkTyF9+AfZpydDqWbSd5gGpKmYV
E5T1/vP9ErGTEpz6wPQ42zTHsi6nT4jmeD2Nsics7nlIv8f9gglZeq1lxmn6XwzA
sxJ3sFqeQQtlKN03lXQKB/I9iqinGbrJcQknL0fSWc43ZdlNwCHTSKsqQ6wuoxLZ
XyQSFa9V6nTRNcxeVcj2z4MqFkbJY3Y+G4bQ8zHrRc+Mt2T3x5BFsJhZue4mbkwC
Cc3ifl3AijV1pa9gr96wD+Kn89cr6ND6ztMgR4TSaIaiZWAcT3kGxb2DyXEtL5mc
+MTKgxo0wOIrNar0szzRyPo0y9nKr57lZhkwENCnZU7vn7AcpBv4QF5fUKetuxCX
IKPyn5g6Hgzl6udP37UwaiTaqVZPAW/L00Wh9zjJameNaIqlN7Z3AijtFSnTU9Em
rFIOJBJDekNcaUNmufOae0xXbwt4eyokJ/NGlq6Ftm7ZrAfkM0RV4YhG8lMaT3E5
3AmZ3F0bkPujlMMkX0II6UIb/f6rh/aiud4mLlQ5e/1CaJ3bB9q5bpQ5RMy7qEoY
BRea7o0hDR3CjEmHf1P0eVLjxpjwG1IvxpeSdkEID8vqRccUhnDxlNuRbHglcgMC
+CLwI0ELaJbDfbsX1TkX0aYMSRcT7wOVB4H9ZUg+kqk7iXklmGCsGNMGpK7jO5Vi
cl5qy2qBgnGGQkf6elhntFfEjel5ds3tobel0Yol0KttKb9mtgC/ifMJuz+43Dwj
Om9IX97S5FYe7IsB0km2zohJ6H3lqbFprj1CFTaT3tRFIdWZ7E2Xt6vnxg0qSHCW
D5TYzCPu53zKicvXFNnagjVGHmp0WixCs1Hs+ncHOzMrzl1iccHv68EijEdwfMIz
Lynlsz18+E7gIQ6ZPcvyOlR2CLbrgLFNDkfF61dntcyRYzhsAtCs7RF5o/utByV3
S37E0/W2NXb1dH4kzs5GrOEWMA8+7l3c36iqaQv72qKG/hrcz9xVZAjYvweZf9+G
7S8jl992rkQrFZodyvWYbvuwk1XnYp4H2l7JdzBsjU5ANVFl0b+M0w07nF80VtSf
r4NpwsyMkSzrrReXRXuIkdbCZxwx+2UOEBLgOpV+nUMoGHGVfpbmXtaDOxf3ZY+5
/n+I7eUbq0CPg7VlN/ch7WaZ7VihO5w1U+cUMpnp2lyizbK06T6E0Jmej/QV50wl
jseN+arAIVOlMtmls/lS0fXXGFyH8T76PaD2rJMVQbH3BcsJ9dQUd9HQl70IL6O2
xIXSOZjKSD6wtsPErowbrNBCojcusojS5v7Q9x0bezDWB/ZSzUwg7TTtm8Ku8pDb
qhM5RkEsuOD27EvBeVkApfix03iWGGMy8zNlmLvVC2jw4REoCgpdnDTEFsITmVNv
KsByTD5n4deKqFQNsNR1WI4NM38Ke0hQMiJTD6veziCLL/aUi6lROdKbXIpuZBSz
RwbKx2F3daDioDQHs44ovcCbmZspaTiosCVLSx0JcnaxDLl0PYM7NkEpndF/75Zd
vupmbLMo+AiOBn/rV+LD3W6B+KamJ/sdh50g0NS1CIwFmlVU8QVBHeC4pWzxd1DO
8nMjXQLgzIzUozmkiZ3DUuCba9gFvXsTr7uXDWD1PWu/cQDWv/JN6NwOkwGaty6H
pIT8znnmah/QYYoNZYyDQV5ZTVygQiTzaxJsiHGEdYCyKQaHNAC1xL1bu3YFEmk3
mepwiPDOPTnKXLD0pAHQMT6lT/TFq6kOOt3RqeEOz3FcYY3GFlsXCrxa5kaV2VLf
QAHvOE+f1FW13T9Dpuj3pKTE3RrmDU6Fcq3UU0vFJTrTbovavSLA4I0+aWwjFH8x
88xacp3+nuV6KcTK3QuqyPzil12/XDRQId4W7evbglWxT3d13cdBvK3qBsl4JXaJ
uUQCAw+NFywC0aLnqjd99FQJEWz6N1z8L7q/dOnk+zlZ9gVWBKoR2FH4xnN3bfC0
WxZFRgsTnZt6r3XDaD7C1TH06AYVkfCApoLDt/lf30yf/Y3QNcfJtURQRIznz67E
LbfWuX44iwzvEFtiwA8Sd7bVtJ+DW8x4R9puqn7URrguPl67HrD5xehwSVLZ6lKO
BEoy3vFzRjvVD9wf5H59kPLwfR2V1aWS34zgGkoqRg6pjb1d7Q64U3+a/3k3a7jv
R/mGVbEeVbrXpcV1JKsLya5ImDPlEfH0ReJymieAU69rz7DNyu0u5pdp+YBqqgNw
VHGkXCqqCyuN+EBxoLHmDlmidYvbGu/Mz7qD9EHpao0NZ4pnE6yBXLo8SqKE12gY
L1G77ftpe6hMMcp8ptF8w4saXS1evnCEnuwlPnDyxDzeHSQTyF/AzWStBJINcZ49
ulq9fZtact80LP2jZrFQmrR06WNizgL4VOtjyZ5U9BsGcs58t+vKfI42rrWIbXvr
d9l6XkRaBW552J043v72/QPgEGIgO8tIIgStEoNYE1hspu6Q4j/0GYOQmWXm7pAn
OwBuTJaxiqoJciMjOLI4ihht5QYjnqhlhLfqLRV0+VC+O5dDGx7zA6ibBshWwB+Y
TtT4jl7dAU1rrvCI2Lh8B0mVcPjUSRxBrWYzYKs+xyTbgLXTxXjVO0WGEeMpj4eG
NBdsXOcAaWFyyN5KlpfIfod9gBh1HB4rZ86qETlDPjSArkGR2TfJNz4HsEhWkdcg
Nztb1PkJDS8JFYmzHJIzB3rhURxqwWZLpU4XyAGFKrC0AKF7lMR5W2H6Zmx1RjX2
/Tw4b0ikjCs2y1bdYG4LlXUwcVLCf7sPlD/ysdzXnoFVrNY1HQiPQOEwh9MbDRNe
srgboScYHTVEA8o6ECWJ8C1Xt2CcWCihZnnW7VcLCIZ0pVP7qRQGButD0DnN6sOt
YskcX6ThP7oFujhyxu0zy6mhqnpx70VF5Wk6T9UsX0aDrjkHgmXYTx+0jFo6pwZQ
1BlDp+qYI9is8eVemjvrELBkl008+UCyF7bgOFKSaz8oGMiPmi59MbK+N4hARJas
BPCulriTDrb+6WFE1hX4w1xlL4ZhAkqMzqCKkFiszk4X/q2tpsI6Pwq3+BzAdwbA
doTQBiAd9sWkMO+HRLuHMxLTsZsON+Yj+0E2UzTx8wfs4LJXEtG71yqyAp8xyO5i
cmReok4I6GlI9kfj9tb+TlMMLq1IDVeXPpAHGmwbFQaO+0SLNhbvOekJWlbn1P6z
JX9DMlN4okNfaI3uHKi+ZxhoEEaa2WIJNC4mFbQvMdGSizoQNV3VuGppoXK6F3BX
dHj5uriwCDuHu0LD6xCYxpMoUe98hquYoD3O1Ai0XZ0tgZxPjWSN8LOARY2bAO7H
9B0U2/h8RtV7I7SFNQ7pzDxKSFetE39JWq7KofBzt6VWIlXw5BcH0hnLlhjXRVrE
Bo7W9L37frHUug52F+gKDzeyQWpcrf94DxOVuB7ifB99XWpnQqKOUHXkPY4xolMh
K7pCkxtttLdJZwDBO0DnzO4odyYPlSwHS2hwT3yzjjtWoo+2pyFwjoXaKktp7Nw/
hT9EE4bZgg71r1YOkLLVAcPjPtb7qckyrDIIweR8mNYLffKdfJYbIiq9ZDKzJpCD
KYqPHyyDx/9zHfSmX8O5nmAkrCxZS0pyclf0dmafcieL0ih6+l1ovpK9pSojHlic
E92rPFX3wQMeFWN/dz7FimSXHXAFzboLXMs3d/dPYtD8fyJ/4LvvOq3DOK3ErsKH
R9v3Z2qEJ17BEfaTV6i+raQ4dfRwCr1argyjXoxvKXFzfQLl9kRWl9vwW15BBL7l
/3cdJJAhMvI2K24xD1Wy7JE9iHVViJmJ8n46mcvy/EoCPi8STJfAes03D5M/Xaol
7PVotA7ZNkCE/JULG9OtqUj7ncsUc49zfr/66uLuoxaaJuUFUKrqCXdriElHtxoA
MfpcP7fRDXl6jT+lUSpYSa5uXqj41Oj7LNrPPW2E15PIMyoj8q9bKRj+4UycoBP/
ib0ljQjz1UTuZ7+5XsHvwVz3rSNkMMxHT9OhKpvWBzUXOSFHEt86pnBB74UcAUlv
7XJJXPGIr+jKV+CcDtSA78CwnPyzRhbuA6WdLGPfXUDorPf6MHbvaT8TD0Gt3Zgf
OGr+m5jSNEg77Qenmv1niZ8phJC5cLt1wSUSRXAX66jbH1NX0Acf+20Intwcv/w5
uB0IdvUbFkgQSQSLb8fCgAQtTqFeDkILZPr7ztGVMT2VTTgHMAx6+4xzna0mQYEC
iZaC11/Gxr3cT+2VzDomFZsflFLRGTctanp7yJh6xkEYAvchvU9aBWJrePefZgB6
uwtsd0xiVYZLsg9AdAsclJkoTxjLISDrEfPqOhdeJ/q96woxIVfXsdGk5uodUG1l
I91ZvuE03SsNYcplU6hHECVrRHotD3q9JHfAk871ccR2d7WuLzblR/6GAMIhZIzE
UzML5oUA4JQ35e+j2fJMwnLmEHQLUe2Sg3cngDl/GHWIadfHyo0pG/A55QgtXuNS
4H5Y2DsNRlyCvP4lgMIBosK1PZ7WcdGAC3NOpTF2bAgWzS5giOJIddR1qR3+l+Iq
CVt8vgL4dBW5obXB2NQ/oan6Sw9cNlU0kEXIGM2TceEbn4JgXMAUG38Q8zvVp2gi
Zl1NhLajx6wfSrf6LRMQCdXIbxIVyo6U0ZWCwbrsR4hSJWWjAfD3TA9twcyUY7UQ
MILIUYsb8DK4Q6Jftk034cfD7WG0H2Cs/REficlw2TlHl2qePABJInsrTIlSzoqx
Gy4FViprNW6YPc2GCUWM0kjqxtn/GLV3o9z7nZ9TbGd/Mo8JLxH+5sCakWLkNq6l
3HuEf+ACtNQjbPunQepG+jEgtRVyH7kxJyEzLaeiPSefNHX00MXgJ8OLe6WLT54o
m+NXr7wylKJXWZ1/qn5gCF3lut0e210J3OLvVNtyaq1gqcs87gluWsQZinzwmBN1
n1ak4rqg/ePpcsY4CE+ze7JhBus44vGJszKHfP82AAWrPUm67eIsgRvr/DcUchQx
kzONx35xyZgaK3a5VX86y0U639OD180S6fz2BOpk6Y75l3ZkdMEFUv9wIs/iFgX1
IGGYYCdUOU3AR1lBSm7FFnApOY5g2f6KsmrKsov5EN6NKeeb1pkUZxWFieEsNzO0
IdSU5E6D2vIA6GWGcmgDufSdxeXdLc322GQwK4dqldoRf2JO/2yvN89aPJqyhpet
Tk2BRZxoTLsRcEaFb0j0eZZmXjOy635bHkYFAtPQfB9aSMpsJ1ZVgbPQbr4qdRPm
4PTGXn1rKaN1ux8qoPQSEGZhzW2b6SQwhytQiOv+HyVOFO47nE7AFhXGDN43Fw2G
kKiRdpUdHUc6Fe2reGNs/+ZimxyL/czw2t8Vjz131+VMk4/DGQnRzukJhMc9rCzl
wklRklKHjidT2TXTFld9Daz4Dq/ppLJcMrMeN+hc6gmH3y1urFp4e5m58JL6Q4Kk
2NO2MOElPM+Q24K0cX+B/gyIPug6RH4GIsydp3n+Rax6FlJQtzc80M671Nqur6XY
FX/WTDZ3fA6f5e/8eQDFi8clPRZbuhv0jORqj5U7yNrEz4TSy1DNHTaz5vy6R/ri
vh5X737ZZTzd9praQVNQRRXK8ZEVcL7u9ogkbRN1cUTlxTUyAcwPKOPhe+3pEnI0
7OxnH/9ZohXZqBw5nNBj6WqARoiiUhK0zTjV00OUEZZaprNJN8xHnyMg4aV41Rom
bqPORMtA7q4aEYJGp1GxHefo3WoSDiKtT663twaNHs1zvbmZh6COncXDDC8kKosK
v626eIn9oq2jLXWbcxUDUaDL0kfnaUmU387Yqbsonuifu0RNnyHjMo/tZbI4fzc0
Y/HohGH6CCQpiw1T/88CDhxRMPbk+gY7aUJqge4fdFaW70FEkH2Xs6LhmtyFWKv5
Lnj6zwSiOGNbLJtR3JlnqmsbiQw2jYQ13AYl2lE9VLUR/N1x1x+ZxC3etFS0SER0
0BDmbmOnzK2nZLHmL/HLcrtoP6FnA/riPH59DmuHrbScYw51E5aUzJmNitt7xM6w
fjJDQQ/MGRMTgKvNuXbe1qzMmNyazzI8o1mpBchPFdKTVy16HvhyGAkH6ns4/eVd
M3wQ5FEherJAAMuYpttIdbUQ0A6nc+D09bQ90UZoRktSxzloCsRN/G9SybfYldwV
xM218suBgVazivO58ARiT/XIy1C0xYZuPrRxYZ/MVujdlqGXccaHt2uFoofGloeR
gNNCqJCbbq1aFJcglDPnvPpVFhrRfrDxUc9N9yASxDGk0DzmQ1HZy1fZhgzvqsCi
TsnCqWCuQa5S5sqYr4cjWkE83WZGy8i/SeBMGSjQUTSkSwNE64vHMXfBy+1YnUdn
kYyyb4VuFFgzaIYbnQOOtQMkrjHYl6zWfXJPO5axc6Gru3Ny0uCeuPp+6TR0CBdi
oZVqeN+bvQJ86dAESpluZGp9BZl0X9aFeWYavf5zL5Mg5bNANud1a/Gydwze9J5b
JA50jRa4vAZ1vbL+HsV5tIcl2ecVsM6wy/GaLNmwwrepyksevqz99C89D7LnMUke
ymWfDNx6FDB7NyRfwRa2pNsLpNJ8tSAk3mxxJcfQxipVh5Pxva/kESN9CrZLoKoh
dhEBikSQrW3CGvxlMyIb4XIZ+cPQjAEnbJCiWEBCnoAd1leol2FiNQFS6IbdyF8p
opXr1ZxP2TlrwaDWGDgGfBoH8X232L6+tydlr0gZ3hR5s703sGCltKVB2aUJU73k
D0//xuLfmmut7Pqr4b+A+L3j8HEKcfkjUuXtr7OII16D0ar+r3YlMx0tyna6Sf7N
naAzC0YZTVyv1vUODjicraLMxQUXJFIzKVfDzkvSsm7tGXMhpTaeyXWltwjF80Tf
r9RbKGOnha0+800UkbqBqUAD8EVCv+G8xqiS9/7OhtY2EwgkM2pyuKxcrpmTdEfb
fhx5cXDJSo0k+zsHM322izQkknQRz5qTCjsa0S9+HdCxEeoo4E+aqRjer0S+OXWF
q583V8dbcKrW4srwR+yu+0k+Ylaz9q2LiajHQ8wVtMxQfel3VUcmiMbeSPJCenVt
k11zog0lgFEbr1heBaMeWdX/TTMjMRR2qZa/oUJDL8m7dqb9yMS8mJBIf0BBOLGx
/bGEHBS4Z2AdIBLkOVqYweuL1fSb9nUN1pfUIAr6bRIBB9MKwvI23LYs+MChMWBg
12I0OaAC+YWSuYoyXot1eY+LtQVc4ndAz2k7+RHmypRVwRJNwcfPSrY7DQuJOtzO
kVAm+KG+Scey9IVRNLoRb/I/8li1B+rrhyldAja3XI3paiifoZhM3sPKULWFWcR5
NJ4NEWCIaS1wPvjCA3/f2aIkAyHcCBabSHYCwIIYYwnaJzrHiS7kAMDcPbfHraH4
18GlKTWFyCNXUt6YJDUD6/RZvHGBytzuHr2Wa1hBm5ikm89muJLrkFfX2MkKGqKu
TtM1hGaDAcirwGXJWmRopU9a14k3+pVSCFIRj86RhBC1f4/p5oFCrHnWKyELce1s
eJU0dgnMHr6wUHXNrrpzcthsWx52mh/hbIbFDt2/0/7DOMJJO8QJtBWK3FM9uCzy
DWFag0b+au8j/v68xYSJkmrwGPaXpIw1BiTeLZCMcDcc1zWlwL6WtoR6OkwBldOs
NUGNvB+ZS6WVYKd/LXSDrnyPmIstW5QT/bOVhjUHWM02BPZvqu+430Mm/cVWXDm+
1jY56TDXfnSIOnWGkW8BV/PSpIaNP0MyncjTbHO5RHFouTaAOoYERUdIhB629+YE
SBP1+8I/GUWmSSxZza6DkZZhP2vyGHlpLGs5rVrpPOxUAMz2LMEWjwnsyy1LdX5D
ly7IOyifryTi/jg4TVi97ex8xRDfHYv/tSVkzrBeaGr6U1/ukKmLui5JkLyr+G3u
L+babupbC0eUO9ZEVVG+H2gFc0KvwBD2FukTD6KrEdyr8s1cFmx8zQYQGx9BbRkG
+bAhept030ffGSB5lRuv4hsB3k6VRDdbYj6zX2AWDU3jVXpgmP3BXmgo75klCNuR
XNh+shJUzRyEc6iie25kLpuqRleN6e7zg+RemLLBZmLF1O0RC81duXvzrgMMlDOp
0s0/3hSO7OeWC0cgugF74g2AKFBA/15wMqmFte9yvvqPDCIhJX1YVffMXDLOJf+T
KfYnDMYRFgmuIO4nHeNwGPOGVWDf3VMkXiKubJYB2XWTdfIdYao2D67sFAZLgi3n
RSlJUz5uWECxcVmE8JuHQP9OdZ7u6MR9qAk3XMYCBgO4IMutSWc06SqaqM3plZpr
x5Fd/W9eMx8I8Fj8QFznB29HPoomKzDZUuCOHwfdkVIGKmfeCkc8aVtibCB8uN6C
KFKKXQN/wIL32nMWqspjrjTmfZyaE3rxeVbeYv7FjboUznSA+KgBA1dFRnthwFPe
3kgeugo7s3Mv81oggzsFVHrzWV+rpFFoCWxCIhJcU/hfNrnmKZf+R21Kg2XpPfms
EcEKaNileThDPdrN2YhbWrPiKgiXhUYQ3tlYFbV55rapdNYCnmdU2+Hi3UOwdwTi
c4GpinNNyNYvwbRgLjJANHFdSX1dFnR4OaWuTYJoUV/gkjnuEmJ6NEO7EiK7Z80n
HUEf+bL5MDt52ha9iPuvFr1Ua19u5H4LxO1JSjV6IAL1QwexcmaJp0TLXGEj/BZg
3sVSvb+fic7Ft+RUcjq+348BxgdQI+w44oNcb940KASlqVCPwrbVq98b9qoJj+1z
r36xAcTBOMcgHlYOZamVldEnqKDX87lubS5pYuq+4a5bu5Z+4D2SD1AsSMrRG6NB
7PQutLzyillnhy9Uu3sUtjp4jGM+0xaRXfQT3fB27fie6f34re1MxsHnGkp42SpN
EtkJiiZtYXubW1dlkIP/jtVQW3WGDh+Ehnafz8f07X1AkgE2R7rFIAot77Zo8Obm
FaRx+r7Yjy91dTgv3Xcu8ozfhsxscLtIuRTiYd1jBBOd8bYEqSnXOGO+QfPOb3TG
N72739y3sjx630oP+eMacPMjrJNMmm/tzXIaemJ/0F16K95H/q/RCW25ru67KWo+
hyEgSmrw79jPL59CdCm20ExVRqycKQb4SngNGJhmfPWpsd0GGZMeKxX3x5mUIhAU
kd3r6Yx+iVPtm503Sj49Hrffap6SSFe/M/cDfqqZ6nZbpwXKLnVHg/oXWAaKKSl3
+eU+k6lD/igWdRthCi6+xaaLo/vVHE7JlINShcfp+4CIfrD9o5j2EmpNbzMZgDLn
penU38gDMuPgpDmq9hcNUbPA/T/u2JCsYiqYIAcxfa0M44UT05bwfuvZaPpROnHA
PHt2+rdk7nRazbdYJXTcUAGSbDdfkqGjtIlqloCulNUMxigZ+EYsz6LtqlUA8oD4
vqtfvtWoky8jZPXpixWdrb0FBIFTHJWlMmxry5Dc0Y2ajj0ZemNymDDRD+bMmn91
wSjeQ7RNHsqteECajjr92dN6Y6OlLrV8VuFGZf02tUmFlaSb1S0zvx4kb0LkoFg7
9aE/8vV8TInjyZEApcCZgZFlfwnPL8YxaFWaiqzv6ikS6laad3fDuVZxgIn/6WyW
yu5o2WOhNIjakb5ehpysgwaH/yuqhrBBynTKwvNjI1iWGsyjMNsdIpu2DVUl9we7
ki3y/X9TyPhTd2bK3mPFd/P5PURaUUnOiQj/vwoqHAFmwFpY7RO3Kpvrfxn0/bwc
2IO7/UlsfwkGSHm5lBNA/vPy52Lnh6hDb/igyAHdPmiNC9BzZYOSzeyJyS8hGDwb
R5daY0YTvgIKgfh6CThUaWHVjHixQ0NLpDjB2+aL6Vwj7N2E9dYhUhuk2Tx7HUo4
IcQmICvXb+XCXtqbmo2Q+x1bZluA6ALSGlcHNL8wLRrBMW8oqJTAKlhRq+oPy0Zx
ZpqmIXXGXw08x/USU+0M1jPAV43iy1jJBGyfBUjIgNskQCIsCTZx/uhvnuiRAktG
X0B3cW4M5oU+C9vLdDRZqm/AieVvvkQWdHLY8v0lDL//e4kvQDYtrPuLuNWhpsWK
viC4rW3YsqtEI09/T8o7oMMIqDu/JCYQrMNA8OKCE8Mzfhv4IWa7Dh3hYd+5RLw9
36T1TqYiCAMVSw809YI9MZBfnXALR+QObzGKhQckAFmASqnSOriCf2TeY8MLSb4I
vJDaj6CrjsCKJkE1S5d4mM2yPm30taJQlAXNQ5yAiZtWMTjzEdcnwqaYGW5Gyaxy
ikhjOwg04j1kY/vQdPCwG+nzWDLHqEv+ZtW6g7y7uRCundFfig00XwZUQC5mbK2m
nYRw4ae/sD2Pozt+bI6D5+DaqXwm3crCGi8YSuj/X4xHtJl4FhrrI9LvoEsz5VQb
V+KTFrTkU/41gv+I+v3HvioSgYJx4U81zgS4hLsL4s7/lRt/+Ox3udzuBzPwoG2C
dcptIrdU/e60JyMmtLRx6eML/b+1QuJJ/xi+Ki4IAMScJsAAbuL/jivwe5RI3liW
1RPJ7hOYuMQyzq0Pill1v66Y9yGPWvX6TxY7KosSiqwExZXt3RW43bOlCYUDdQ5S
r7Ie7fchXwCl1yrQdLtae/O8c+uJtRnttInbJJJHwwqIDqDcdlPYbhQTr135H6qW
uohbZMWMnREq61osjemKIRhJQDP7OBXynaL9ezWhP4CiLNs12u14BOB4wPUytCEa
IdjgmTxP4mXbofRZKIswz8wOWZPtoP8Knmdihb1mM5RbR0bwCp04DEe92O97CZ3s
Hpam2PL8Klf52b1ZWWesGatIN+wN3HtXAoZtavffMly+VN4Xa9NrVp+L4JQw5QpZ
PlOjR1d1RGkFNm5RfTb9lh1oH89Dy1lmnmCYJ/Pso6Uys/bWNGsGlOcVMgUMuIdP
tdyVCIGadKA6kJNii52X8wYlyNMXQ4963883QcT3cJKqHHfxJ7P6wfCNLGJp64ez
3DTwwFY66IUjE23GjrAiDD0QxXtwrFhhj7ePGSME2Sl1D0iPaRBVSkwXfIwNugTY
4vuq9zOjdZhFatGOdN77Gala6TQLbmQMTcgpjomqqmOqy2uyQ2XZmy18/i0YPvg0
423D0Ay1Hjk3wyJJDgYergw2O5NtcQZJVojukB7GILWDqwy2EsNSAeRqMF3ZmBI3
u/3OtT4E7ehSV/9Abh6Zx1DWxBF5Z8AAO8Qoa1Tx2Bm5jvVmu8OKko25fB1b0+rP
69F9Sju7c09Gh4FO9d7YOhtVAepeK4Zbhl0r6HJmBofJsecBb5+XMfV7XWw6oEyR
iNBU7KDzK9rirZAxOyP5ylhU9OjG5PldjQJJdkfSZuhDKJH0NulW70eAk3UL5Alq
zgELNmbn3kB0eCKnJU9zQ/liDRu0oqkZBWLekOpq19V6iaU8L9ls82QUfQiTQBQI
sN07Ygk/b0a7/nqi7Tql614JwQCYInEH+mU+QXVrCANOFZHoHj4y5P75UHymldrK
8wYl6R/M5Tq2LVXLZrGg/fRpxtQHV8fx6tYZckEtXcgz8ART7srYR/l2SdpUK5oR
lrCeyGYd9YR9bVbiXxgo59r75g+up+KWfyOicGbmRas2Kv6yax82JztjNWL8vvVg
Ftch6xXeRb1+pvYERdxBNaIxB0jLKln9dJOwcolpDnIvxWS/c3wfDy2zL1RhC955
dJv+DOToqwGUEPZX5kqSxsxHZOVRAR08erd0WoLLBekNITIyCQefXGL95WRCnP9F
oddEGYNXWxQXAVbOYns4Mv30hZx0C8A7uzXD4dY9OyqrloMSjSRrcRvbk1ZRtirt
xFovaooBG82+zrEov9SgNA89uS/ALRwt9lzU/etMyzQXELo36d34TDi/pMROkHPg
jPZ5kRUhQHDGxP62dIEcaRjeEB+Opny/b4s1Jhml/2OC9LAgMf5O6mLX/EQL5S9L
rWAZjaQKpBZ681MGqnDlhMUqmxM7aADpXRHvBq14kKpxMX07STuLPm/qZquPtGJV
BWneKaBRyc1T/svFV/aZzq7VM62dxW1IxogF7gqiXtn7pJVd5rxvmqgHWstss6V0
qrys4CgPg5Pv78OWUp0kmSFkX6ntrKveEE+kGFV9ffKpAZtpCc6WJ1OMIHNSzl6W
Aw4qMo2OVDXuRF7YJey0REBqf2w7dtWRa5C96zjzbGoBuZAcAYxVbAe92TeWtvWn
shsnm1pQVJkrzpYtQWYbMoXvzd85t9Ev3icqcszKjpGjwVDVtQWuz8iXSEdpIklX
KdykfB2OjOyzZVe1VwoA5BwoQs7LU7R3S5MBXESFKrxK2f3M1spzv4cvzSFpMANC
RpkOwtg0ueoTRUb7o8Y0Lc/OZxz/s9sp9rFP62EP5pvyt3HNTvxROf2EDsgg/wOY
bc0pp1BnShsyp7aAHBKaMkiSw7b5UPFdYHi09zynvalbEQMVtDSRVmg76h7IaXmS
6VngyYlWsHBBpbc2tjOUwKx2R2ZxV3eKhJa/hXG4kFGLWnVvierg5QO41ROprgNY
vXMFT+MJZbNF6cAs1zaW3a6K5cgHC8XoffP/gdNZsb1q+eHavyklX80k7mC005rI
duZjZRx5/S1yUF20sHP9CU+ewnPDaAHt6SxvTVDQTWjnKDJooGHK3Lvh5HcqfbkO
TRrVsxgAvwwZ2oO5AhTMJKF7m15HGdH+OglPoJ7fltgIKSk/P9jK5pxwTLtlwQZW
da3HtjyZwDOIAvN1+mGINZRwxHUqQCcdaGvRgVGRCgrIRgwm9nUUTn2+qDYulgO5
kxjuSBCktI67J5MLaBX4mkvB5izOF7xWggujuOBnzR5fwXiMrwqvw+y0dHhlx7r7
KoMMeGcNSQyD1oPdnHFdBGDIgkeHqF6K52s717NAjqfsnNiQ3uVs3sd6xpP5q8iw
pu+pVz5Tnr2iGwNsRc5c7Qe1NxopG2Zx+0bo+zobYd45s6+qV6zthNC8Q2xZ/GUv
5cQBnaIKzZjxYBESuSz/M16gI2bXi/kHmwk4s2+o6WyyPu7aps9PGGbHR6nh2+Kf
faeX17cJH/29HAHSGYkgHMhUqn3df+GA32CcY9v9BqNs6fNf+Gm4p/Uo5IGuUWtv
bLGaCeqaLM3mAzBfZuqyK2dDpvJLTgbXaFxwmXsUnJ4LkyhTgGDOTFFgnOYIjClI
xSvk/0baXahpcPHTC90L6Opi+3AJiDf3kxGkVt384mQxXPb7gXmKADSX7W/auibk
0inqRd5hTEQVJuroL7eGm6ql180gZhyGUepRm8F5CMmMFsr8mvjfRZmKqHkKoSzj
aVD8kEwAcEEAdnddW413ea+Wi2hoMxUjeXocS58dlrxK3GUHbXKQivp0XWdL/wOD
edrrNWV7q0mcjtxWUiVA7tJNCojEYkeaxmNOarACKQUkRCJgRpy4mZqmnsDf3hV/
Ib7g0flFe6Y8HGvcz4yh8Rvij7rLpKMOohQqtg/wtj2MzIuPRGj7XDMKZOMpliOc
67QCULQ6ZzXc1/51gwJ6BzNBjt/cF1xOXLytx1IKodE2ridPMRd6DBJlIkYKaT55
oZlI7RuTSTrlx+4zFT97DRiysaFKN0kg8QtDt0eMS4guCd79c8x6CodZFwv30mkA
pKIk995MTiTERLYTPdWEjcnGzvs6soxGFUS3aSdve/LZlouEKRbqN9ZR1aZ2Gs1s
LH/VUhs3trThBJLRZM5Bcu4m8aGMmOTMvPLYmmRBXxZs3NJn4ZmglfcER5UnZ81b
q97O6QaSkMeWXgxhJo6bzYYmEmEpHdESMUq/x5RKC/UoIWjUPGF/ry/Gsjv4lEa8
O+op4VfOnhLUF/WQ0zJJMPV22adyhY+D5hbyQD2lC+bC+QWGuCIdutiIqqSBncJI
LFpbNnoKxxpqvXzYcFv7qvFIRaFYW+EqrTJW6Oo3R934UJaMTdnMhfbnY5S9+fKz
BcHQnpkwV1BB846G5CoAa9qfyrfiLeSi129dkyDsW0IMRe2bkFqZ2m8vp06wdsJT
8/3Mm+eTNMzNtqg7ZfTnOd9eEarggF2q57HrsA0JMLi02fSXNLpXjZ19Xd3TGvqp
06qVRfZM+dc6Fno5xmp3cmvErmgPSKKObo143N1ZHKAfQVDKoo4QcoKfmxCAwLhG
0QqbkWZa83e+RDNmYvQZRMkDtF/queAIqh/S3ltzzeg8UE78kkhk8oh+VhusOWQW
YSGBon6persEO1iZN9GCvg1BqboHhBQlhV62qFczpRWRuKO8xEnoW9nqSLuIDOnZ
UO4kE9O1cHwc4HXAi6kgbuHQXHVjXIdEIhXHtE3yHOj4G4l2/48h31wNwSVBzcDs
RKBi5iL/Uaye33fF4IBqzoS7+mLwETW3CK2MwCEejPRD4cYbBIg9A07+XLZvxbe4
6nTwbZkX/gHOMSxYjo8sLzIE5by0kUnqSYEoLRWPzhhl+WejSlOF8JmIxw0oh0Kk
1D0ea2I5Ms/H5KaWW0A089069c+4s+VBU1nH0DwwN8zKEHShg1x2lpgsOkqYm6Al
UK9t67n3+fVJvzy5exmD7W7BThkg3bQe6D7hwOU4D2kxcXQanZ0nAccIFJF5P0sL
NC9itr3yW0VH5rWGzck4eDseO0TLvV5qOz5jNJ1mUOQ/BknaeJGrZv9q2f1B26p3
3XToLA4hMUFWnzW5Xs9vg+dfG3JaAJ8O2BsCV6fT7zABW67pGh6R0qINZPS92jQI
qT0RMAKUDesTTl9OLzA/ir+BOILW+vWTgIg0ovEf8xgF7V2Hxxo72DYz84mI1Yw7
08hllpVGPiVROpe+4/Y2cyZdwwZCJcILOVuC24ibW+E3y+6zyy9L+idBBYPnqR8N
ODRUjYVr+a33ElbD+uwK2Y3d3cVseCdNTAyYN64NMa4hLuzkm6CoueZ4VNjf3S76
kHR4VL/nyucY/Si0hRF6jt1eHILLDvT/DndIsUywuk3dWUelz/VOKQz4ZBeu8KkK
VEy5QZCayLbLUadauAKbLLikEIDuTJ7UrTsK9loN88v+wm0syL5aeaDC5muXR20e
z8q4tTfET5MQQDEhhbQC5JgR44CHAKh8dO9MPWrpVswk2oG269E78e6DGKrD2Zxk
9Ey37yxbrrpw8q/lHFY06oVu6ICyPYdeWO5Cy1P6/pRvJJLJ0EyBS+hg9MFw8AZI
IbQu4SQ3tOVPIb4SWDGd79zC9yVdZZX2A3hLRXUCTSZ+fIYj87jNcuZqt89Cii1E
5aXzCsKDewrLwRdOPy1CeeaG5duJnkzFyzkVvmGdeDWViDZr61ppD4PZy9/GEPPc
MvM+glh3oz7NF9xk9MNWrsnkt+QApUrlXzLs65mLF6U/Pf+XvAo8QQXiJ1n5/fwC
2f6n5bcjy+soE3qP57m4DUaSz4uyqjjGO/jaWKxJvNA=
`protect END_PROTECTED
