`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CrdVQ7FHT7LdCXAxnsn1pO17MCct2QcRhqif7JDH/cEyIW4qg0Vhrzw8PcVWLbUi
2jPMYb+DbvpIF32jOw8r6RCvxZpyRCCPCb8uVnHqr0UMdBPKjanx40coADcLZ1p9
IRJDkPna3lsw8+86lOUb/hvQI5kiywl+fgVEXirk9cledl7cxoU5wnnrS5jx3w0j
JPfJtOawVrLAk8TNGTc8ig450bEnkB0QyIy5v6iGG2LsG/YF6E8b+6hivs1JiROk
sKK08TqOqegsdC2UcDQQ5NAd8W3q9Z0B3vk1Y2ihn7bOrvxmCIVUBDnlChMgMw4g
eoL6pdlaRu5QrSwyvK36phMEoo8SMTjZ9DtRx9+V7P3Wcvx0TRx7JDkW4RDLwats
dYxFQI1u6Pt2yeOJhZRPXzA+fV/WJK59yJyDiksKM1VrXluE4C8R/wMpZ2uuNP+j
KaeI98CYDr+o1gy3awSj0oqS96yTl8kNgIzMtdW2BEVOytWjbGgVNVWGgSEsJiXQ
syyEZcWpKqn+eGq9SToVJ6at+02OsgMq3SqCBMCX8XVf06u7urxoKNbvAuZZnzDU
/n7A+OuPxpLVmlSdhjleYZGR5HgnuIqsSCrgY1DGT7AgXEehzp8nxPba19bB152z
L0AqWl+KqAoZ2r+f5SMt2yimDgkheoAteGhnLAqEHUvijTwLmnCsgAIoeLsbuAwr
rsmHqoSliVLlseLLh6DpO64cJ1dvyDkT8a6uM8z07ZXRYBqzlJbiL3sd6VBmtWFR
SUqjCBLutc9TV6NubqCTv/fVZ5NnNb+WyZDcLFoaMwrNX0S0M6JBnti73CtviZrK
9BoiG6AEATecfeGJzP+2wKWZ6YwyQQ/ch3o1LhHkj3bUBvPKUR7ROUm36+nwWXL7
nItuC505NchkVCY9RLpQDhroXXe5m8ivO6ynCIFxoGUhmvULV6xMX3QcRguzXxx0
vdkMpCTv3AvqHyolFj4fCmmNHXTvhdzU2Huqw606WO3jGkyBjvTcjmuF87VX7B+U
Ut0myHJ79HvXSACLhl/KuE1KQFT6AeSCjZ5S7mKionrya12JcGjr7kxNSCAB5Il3
fhp37aRzWdzABhn/b0chPk+N08/lEiX3cuuSRHGMoO7YzaWyZS35bcyCRrNb4sbY
QkXwzSbY682h2oJeodWNrYmG8KFgOixOHATXinP4snSSYlenPfz2gjitCx+v3KgL
bfrjJwUgNxrosnpSXHczQUezYDP6cVKrVJPFTyj6pAf0WSx/LVI9oTsHbLLP7WkP
ZQrxfX49jCARqeOlirVp1SKOwmwSIGNuYFDwx6nVhlZLbFUzRpDXky9f6iCDMhoC
ft70wumzD4Yg9YPOj9+54r7BR3/ten3KHFWkyDbc02V37H0frL0Io+rCqzNnOayZ
K+2CJ9xqae9OihnvBs3penX4DlwpmCot3IOiS9wgw+S/2EhqRCp/A09RGcShgHzR
h5ZTmcN0Q6YMetCaMUJVKgReLPw3CWfJ3qH8UrPpRGQ0mdxDrcXn2+bD5SQ1eF6I
3HpCFM6Tt3qSXTiaQPS+nsga672qv6vAHJYQCXRRh+otx5OtQd+sScHFc025o+7r
vIaiyZYHjuxK4oRlY9R7nNPY4VGlSfXGR9XSdM3GYr3SLXMr7DGNex1vlCqiyT4t
sWZf2YhFO3mj65HoTAazE/cwm2mqGWbHZumi471cXOUjcLm4FwB2dpx8UGLQrYLS
6ObrWnWeS4jkchPShMg5D6gTHFAmeKsGgSK2qcI/XmfQP/BPYsWflnzOexrvD0TV
xQTaQ0t5pMkJ7XHEJ7NcMwQhsNbT8ZgZh4St942kqBI+8B7kL0UeRdjERNlTt5F2
wpKxAGB6Unt1jMNUifOc9Jl2iKgc/KQByN9h4C73FNkC6xL2HXg/qm8Kq1ZNFtnj
F/EFR7zBZlqyyGl3WFNByfSTQjtKOYIlfLI37qNWvwIxV53N/dNvwVdWdHRbgFKB
+orpFO3U5oYhpLvyB2EDXKHiwKfIHSdNRtfSkmeJc7wm4JXdrAoeM3EHR9O2mnUT
vCx7sbI478ufsYwbGiGk4Ix7CGrliDb+lX21s4pznrFpsd8RptajlUcltnXtJKmS
qWtE+4XPusj1DvvMcE0zGGTxAnJ1Dq8mVTXRd5VxZq++aCGbnsQ3HJEDvhNSl0Qb
zV7NJkJffJlV5n0M5kD9vk2bF/O3XNrR+AhDQqe6a1CC/nGFRPdH1dLYx+wib1pn
o468kSDChxsRvxti1kkV63BRSkeBgvUa5JsbJRTpsnO+ekXTHnbyxb5Ds0EgDvol
YvpOgYBvRXI1ySpfYQWKt61Sctuqnvtg2U86kRrYpWROwH4N2qIkkQFep+IBYxjn
1OkPBsEYDPycS2jLWf+bUeyQGqaSZ0vAz3W+yLiPQ+Sc6PV+/7IPDFoeqP6R5Etn
Ss+RMa4zoiXjL9pRfh0zCEBQX4m/c3V4WUh1RS173XWXV5ImAuzwpOIIaWgYLHUZ
hlS1tD0dYkeYFWrqSxPh28PYg4QQ0uHM7xK+uSOE0z25dN1XVp0y3qEXRkOLnbHb
zFdGtbvrQ9MQMX/ZpCNaFRI2SzK/eyE4JOxgB0oFVoEu86O87WZI+dtdI/gz4pDd
cCdhLf8i7TobvWwyNVnpC1CyfVFL5mRbMrDyfUAQtOFw1yXRDwHJbNNCVcXgJdsU
CZi9vLdodteQ+G4QEdprOF9Aec4LNaSVtA2tuZK7fm/hBOuugJ54CVABByFvXSfG
bZvJbMrVnkr5kf6zqMaX2rGaJ6odkOoH5PnPntHLw9hwE8Pas8TkXUKD1Z5qigdp
1xjll5/UVBtTQ6tSRGlE2UDheXHtqz0UE2RFeNS4gWRzSWSSggf3L+SCe/ZeIB3c
PRKSjrKk9ynDAHymWuEnwyS8TGNg2M/B4vr8ZRDR/6WUq+6quUSaMq7aGiRCBamJ
iEIcToYAEJgrfJ83gKuqOTjhzC+9aKv4jyNEYIFpvH8U+Jw4U0CjiBIzGjrRs3J4
zMw0gXlLYxOLLAYm1aZ6xvf5ZzVK5WD23iFX3JtFn4Ya/Lf89Mc52yH0EE9fnhlT
gjq9NsA6Mpeo5cnWKr9sc/Pm1aNAv9MEFomguf45/eE3P2J76TSaV6CQCSqRvgoP
xriEzYFSUk8Fxx/eVwtK5l2ku0BbDisIp1HzgefEn7KhpQ+Yd8yXQiSVMaNH6xVl
MeuZL5TMSHA9+uymfuuFGSBUGDN8Ca7OCLiyesR4zti9ounE687tm5zTI/V973LB
1oj7cNqxbVB1XBiZ5ATTf+AgwWH+HFvpeTD04IEXg2j/rQssvKBh7bwz3OB7WVJ7
Hiw2gUg6U9Vio8t+IhouL11+10PgpniWZJLJrjQ/DRRd8UYSdlDm1k3dmCg9u85x
jcwn3qj+yBUkwTVtLiKqcRCkeC9z9pX/pyX2fsQcGdsOqK438S4g2CH+XMQlAGcX
O/iQJCOgBYsnEULBLCkeh2yMJvvszE7acP4hXdLuQ6cdg0IlAey35WrGoKAvQhjF
NC3aatyyajH5OM3/b2XWzR3CSH2iHGobKm95knMbYjKTsn4CXv7DWgcK+uAY9ev7
7/9G/Y0zQ07I7aI9g7dX4FxVBcF9ERnOo/U92OhXuwbe3XNa6w3kGE2VhkWeRHHw
0eaxFFAlJQa7xFKfFmjCZYBTlVAzvGrnvfIrVCwRBMV5WnXsJeSNh8K4ygViqAdO
Sx/0fbVfO86ra3O/hlqXuY1W9Rob8SKy23J17ZV+WeRIrve00KZWwtRsN8kK5UFC
PxNSYT7pS5jNCWT0Y0QIlSdqI/DyjmN8GkqLYhyAj1YAAPHLJW8EEomwvM020NvZ
v5ZyvkTDqn9lfh13n0n8+esVj9DLTAxMupx2Y2hbiBklr/o7JW+JN31/V7iU2FGt
zFLedGtDl4XIFrfLmLhZCsIfrKh+oDAQsxwNbjLalmAA0cV+pz93pe3I/pDwJ/wY
oNG99xncTZOTRV7fuc0ezSi+mgKGS2FZ2JssfosRkCvd+7uvBtVPjGP/GH2j0Ufd
PuW6/tP1HnACfiEdVhSSizljYMBVhKunpBtqgcKpp7xj/Slq9+QOjPuX4MePcRpR
x2KMb3nZ0UiebnI7PjGfy1GVO17MNB8Ezb9Kpd+GPTXVFi/inpm4oYANLVkKWQun
te15PpQJKUosewiEwMKUAvdN33etmz5ZQWx62zcieCRaQ7+pF7TEtq32tpTakPSi
cnTheAihbIMZwf0z4+cGKhA3rmFiSXeANgEQ18a0fJf3tSaG4U18EV92NHidJTl7
q+dsSfWS0uGfx+Cp/zCHeCOL1fF2x+NiA5W3hMux+Ay6rrR0oT0LWhtDrkeQeiBt
Bwp5odF+Qr4BkNJWOGcSyc3pYIsbUhiazbBZjPHZkxB/8awmSsplSxJtj7Qzk8dT
IiZBy+u2ojttypSQOhn7+Uuy5OZJml/3iSypgKM/0Nd8OtNQOyW7jkwlSLiWOveJ
cRpL/I0X5u9rKY3Cp8X3n32XQ1trCxzuEwmV0eFz477zPM8pSZZ2fH4A6CQga9pC
3fZ7R9dZqxrNTO6iKJa454+o36mB8AqGEpvzxLQ69HhrJkQtZti7EunlZiMGGHO6
K/W2emTcH/SMMQraXdRO69sncS9xBnqqL1yU36aZqb1LJdq4Yg+YVL0HY4aW1ceB
40NpE9eks1kh38w94M+4aM+NaxyBPrsP7TYixbtYJow4fmlOacQhdcqd8F7AJ5Eo
Pjl2p8w7dhaOgyFa+dM6kX/Ye10MxcXjIW6SHKY59caG3TVcanmYdotrJLHr07ES
t54nsSPE3keQNk9jM1JTTCXvRZVYvmisSI/eRG4kv+l2tRHF5ws+51E3/agYWpu/
u2WlQR6pNF4qxXP1ibPOHmpR16grwppsn4zYIG/2Ag4BRDsIwDNIZUSWLTDrP60N
vx8m5dw4DDm7yGNl4vSVFHb5UVDR8jJiIVUZZ373MMVQ7+kwsyznXDNDSELQmLli
5kNHixe442GgHOFy14XuayVsimfMPKu5ANq7q4Ww5B2bKLMJXkyYl2Vdbh7V10oM
poKzfUKioCW9X/eVCe924emiPtL/tCGsIcLGR6CczuVgBqcVxX+TXGzR9hyTfaJw
hhaZfKD5epQ83H9Q0iWL165mjpa62+/NYWibeWgirsfNDuoh9RbYfBjzJ0CHxD2b
mpLkaUik8AkoQyykUf6NiXORFbH6yZAS+y2yFuRbBzsLCxTLkdUesjlbh7dYXNns
+Th0C2+VPYVM1egCqVdqnDsV9w6Edxqp2nXVKtflooGVWSnFSh0FxtXrQM1nCFLC
8ODGztTuZn50zGN2kd8i4KiJJADAR9UZXIZOhd+GrQ7X94j+HpT2dhYP1n6EBdRU
LPvCEWh8FMiDWeH+6LThZgItUkNezvm3dHJFSG4FCb0B1liB2kaZvK80BIWtekuc
T9aZXpu3jdM/A/y65RfKRhiOSvpmNd5rPhnsvXH9x/qWm17Ft8XmOMs/Om3d9V2T
WeAq3kv7mEvA+m/+1rqTKlqorpk9+5Mrl017OIkQLB3bvR/hZlPNn3geKD456bYg
iO8VAohohb9aDZ0q6RADOPXFBefA9dtJ+ilLR9xQsNTA5ybICnzhZNzMtojipeN4
12HoaTQQVgRYjDUfRH8Z9KX1dwFonGTb5KR3CUttFuDnC9uxZ2UWP3pdsA79IUAy
Ux49OkfU4o9T5GX2zlNed45HREAcqRG7Cd2DYOkqSe20FehxtxMLD8VC4Q4AGUq4
NpGrFXJAOsOG1U8aZrrCEdZnP/JYX9G/8oGU4CPl9FgccLi5liAFrpeR5rCZybow
kLGu5w7/y5F+NQRsRxs3nR3+oXKLmYULwj5chdjFTCqSKz/q6Nzjls9Erw7pgsu9
cQofxRbwHK+B9jFFTQ10qQYEXa5fDNRgR2Ff3GikQO6JA51W9uCCeG4RZ4sMeNUw
u4GMksMsmMBT+sv2dntE5a1YJpKaUREUgsbJVQJo0I3xTls2mlNLPCX2eKfetMpR
1Aj6G5ZjPj8ZGnR02Wwz82VL70mluttIg7ywhO8WyZdgW8k+siDkJlHTK2ONxNv9
4RFsxn3l+HzVpsQISDaf3mfVfUmuaJNBwdsuyKjb+PewUFdhuCBNAAkHPCoiaJpc
y6rLx2jN+4TUwYuQIiY9Sigu7jAB7+f8ycdrYnqeZVCws2Oe0nYTEv2MJgRRrqkT
iS0pm33gLheF65pCj8+0emmhc2ydq/eHE734yxpuU4ZuLoWbz7XJjNC6HRQVh5oI
Jk7/URl8SfRGj4SzarhUXHwC9p5qFe0f+sR2hqqL7NyOVx3b5pA6miabKSf1iICb
aQE2x3ClPddM8mTRCTGgtSQ6oKCBAn/IlU6YdFl6cnX6RRenUJGgcRAkP6aYPu1v
qAWl0wfP5uLaksin+1nMSu123UhzA/BOQWnzCpz6gAiHQR9Ln2JW1z9rwLngtMB1
3zu8DX3ZYP0WNF9SsnU4nPzU029xnLIeuk1Frhw0pRIPoVE208r5taDl+pswGPR+
1esQxB7lN+0lbmb2JnYBunnOqWV9YxPx46ZJCOAyfYcWbS+kkCnl+8SnJgt/v92l
XqoksoT91btq9xzqeimaOpWeqCq4PIDp9h7Adt5TUpttohA92R9Er5VGfhuPXk3v
Xv6YWfpaN2d0SRFE5j8qRyuZFVl4RaUm/f4qmHv8KBL6tparq16UFDvMGzaNklus
qXCjcdTgy/t4F0McjN6OpF4VDRH5M01MCaI09+XSLZcJ5elL3j8/I2cr2RjBPzG9
D3PCD5MGuVHRgsY9Fvfm6/HcNzjBk+aiup7mhx6rFDQVFZtmIDrCX84gbGVBnAQT
U8vh75un0tqZLZnEkSgtMlUOHKYPpY8I5H5o5k1Ow3SZERxC6fp8r8ynWH8+R+vi
8Ntf0gi2ahyMMT9uY5kwaj4dbyqJ7ykkBntLt6gSwB0heXZjxQ3w9VzH6gLriJJw
z9uqm9su0CEYbJVnt0Gf068YZLNODx4GgihgGlUINasXYxDwO48Nw5jqnanCRGG2
EIKGCiEGaMQOZjSMI/xfuMgCJNZ/laAPSuler/MhweFcnARUkPjtBTf9gZS75v/Y
1MgaJ3BZcHkFHt5/O8ci9YE32QTKmmBre+bR2dGIEbgnneCZ///u4j+o88wjkrU3
esdWj4g380WKb3zTfXUzTK1OPAeYgfJl7OyxuEmrfajT/wcu/pvqZf2Yekr3rxOU
4GT45frXAQHyELKCtE+pf+u6MIiE45GXZQMfSIySh9JfCo28Fyq4s2dM1l7nLccq
TY5aDT7pRJflkbgihZWQjBVoBj5QveWOVuK6EsdQx0/qmPEsZv6hnpMElqxOtd5+
eV8cXK9BUbilsJlMcakCo+soaPQ1QjJjSMgFItIVnkNDZR/rADJIxW9OO7c72IB5
IZHvni4TcLxNPYj0IU7tGQHbm38t85N7w+eaovW+iHo+Gf30eGkOVBu5VEx4/Ja0
tkXgTYfLB9jbDiqndonFCE3B/1RlIaXZEC9VBkTdjywLS3TYJ4AMpwTLR5PkBvZw
FCpYRoqyN8tTVAIxIbDHlMnFGFmnQy1HNtX3c1jth6OqWrikt+3MWeCmPq2UKKNv
EunYfhda7u7r5AMYTob42Z/XM8uD0kuUxZvWoDsdKT/LLuJc/2NNLPUSRhTNZ5Do
VL0aTeq5Kk+FWt34fPwB07Rpqz053vrkRs5oOnTbzAYmMVDxKDPs+CsZeuQ8QF6V
p9VQ8XG+5GNJzpG8UdcdNKXD5/CNdmnE8qmLBcFWn1FCzD1IXnq9AnnJgeLc5qr6
7ZLOldndYNU0MTC3c1vPxmOVTcOWXWELCQZ4h1nVjWnHTPvhsdaashOEb/afiWfR
aEbWc6BLpZ03jq92RcStxqEl3PPmq6yL9p7h5wsUMuD+4jq4kKWbvOFUUynMvlTk
J4NHcl7uNcJw6KO8oMSR9W+09tChg4ukMSNci9rvXA98Ep1TUzWDCfOdTJvPNYYS
TELl+w5r58GH6+WL27kibG166/2Ym65qyV2XOkU7otNWgGa18BZPR1BR7r88kKQa
sjPtbQYmry9qfeyd9SdcAS9VXrKt4QdaHwl5W2svqLkU7gxFwGPV4eRRLgXcdvEH
pOrjpsvcyyIDXkCuhZgds2EfWkGzB8rFBneb3mBDvpOKeQP7EHxlJkcHfiBZ+iHU
S4pQF7M4/sQwMXIeRte0aFDE6YQpOQdFTKsVrB62k7uvwYN++3qzGKrJphTmU02F
5dOkf8Fe2ia+6KXd96b49ksDDqhgpCnAUbGYB+Z2OHJCs8tDjbThwRgzd4U4fqA8
kc3Rnyocg1iS2IzjI+38UyiYM7KVLLcEfVk8cLsIoa8nsxrrepsQ8IrRNu9/T5wf
Z8Ojci41wK9Ntor6cN1iH61R6SZQ04PG0wNoaDqEIktvhdKJzFJLhLDXM2ECMai0
YpH8KAwpsOBeu7t3PO1ZfhRSi4RJM5ez7LDtKE49hlY3q75AYuVaVNXmVf94LNEn
ibdmn+zpY5W/mH8wtX1/hiGkThDVcQpADsxpt8tfY7UV3rXQcOtaEAyi3+WrZQ5A
Z+4fwgGCKQdrwLyYlSiRg/mL6qGd0HU9H/2ayXqTDUM4rd1/T6JHzpA6E7U5YEnB
/+aCboVFUbo+VuLoWA2KacAURsAr+yQS1b7VtSk0AsTpPjIvGabjw+8AW5L3B8DM
91B8PTAobi6Yf5s+ggTmlxjSvc3IdLJa18mv6e6UrtEIqqYHm0H2itH/opH/O2Bt
LUIIO9F5MBNWAlAATC4LQMC+GPGQC1y2mILQ/jjnKTNRm1hcEqmK084MYWZKgmGl
HodSkrruEDW0lISKxS0B3q0IeDNYHBzUljG3DWuyXiX/7HBKUdk3UGYmvOxzF3QF
54jjzVldUqttGTkZjvK9Vd4+Pd6ogq7KWEuxAXPhAHRjAAcPkKBLn4CtqhLU4Z48
QhZxtdYIfrY5r46Ot4g2HzoVYZXpwUkm9Kh5wpEMC4FP2Yi0Vwq8ZOgIy54W5EHi
2spSzaCcQoyggJrkDHrrIceYkHjJkMELHquikeu1v9qdnKWwhJa/9nFtr4bToovA
QbGfQWZoKcN/DTh9z8YHniBKzSs/mhzRdC/I9Asc0/H3DARzIHn/lNp1tP4RkJII
I2Y8BCf09SXLAGSea43SKmX2wLpgoyqSM1g9aC9FgWCeHnX7ofJo648eC6ofI203
kqx2zvhTGc04lH3bcTw+BmTyzbiIPbmKM8qQSNewa4CRRCY6uJOYPrivGddZz60L
SPTQysb2bpqOhdB2raw8mrv0xcNhWdhudcBdF78n9T/DRhBa16ka9wqTo/58bYoy
pVNH8sppcMfXkhV16A8H0Ku20quQhY1xNrCDJEI3JEZfCniFGbfq8gKcJRTqrfin
CIXN9DUPELLf7BD8rQD5TLAsxvhFtqMuy9jZ+2dxY6b6YvD6UVYYSjXJAGq2qFYR
b0LtW12V37yyohL18P6l09SN+bat0zYcByBrmUplDhOs94yH2Cm8r1It46o2f9So
+zJIbt7HUbmGwfRfUVhrtlz7sRhOlWKRHnZN1re3UDEmXH7HTyKNeyZfaVkFJ1n0
0Vf1E7boBYVvyUT8ETEeczW9yz8ZQXgSxLwfDeghrypUEI1sEjZOWg74Zdi1FkeR
bPCCX6KLQ/LOvzQOu6F+OFpYpOQ0s+5jpkkJ+NX1UOtptPtw2YBrcRPCLur/idd0
zNV674boVQUpg7BqiIrwNKXA00StT8zNOICGIF8deYo48NWFsRqASJYnldRCAHRV
ShGTtuWY3Jc6FCgk8YVGf+WRjuLA0/M8oxo7tarOwlQ3Xrs963WfPpdLjUf5JIPg
40LtWTorT9Dx/LIX5Nc5ZSz/779AU3kSiz9ekFQAGXsrhkvBle2FnbeIquEaIKY1
cceK3UYkU2L+gPsjhe4XhHLw660Q8iwLKvYTFwHefDouiELLVXz8M8zBt7+CQkI0
bpHWofzZPBEPwpnSuRo14M2J6BnnDh2FSrkPMftOBvJlzNI20BZE9O96FvQZDMcS
PPgvug/jkUvKIB8Y2WapxnH84gMpsYhKFFFA3AOpCzCEsvh9b+EJwbLYLuFlpVmw
KLEt6u16VKgTbsyOEVjheEHV6mTmQzATR8VLSGs6gJZwWeXGzstC6cdOW58lIHD/
dG6o0ZBhbzQ8GoD4Y3YnoM+iOfu9O98csCC6Z+RyVmO8BZEKK4mM4nA1FkM6WHcQ
t9XBeiQJfFumDKo7ijs9wXMEcvabHkoOzy9HYKz0KyFsDc6Jkelif4eHrQSuxHpd
1Ddn66uU1Kfc+Gf2oMfVKEHaXlTwWwXPoOFJaKL61D97fkj7jAa36abwLH04GcLs
EKTZTRx3nKQP80ryU4ZGEEtpwKEHnW0OfeYoXP1Uzr/HqxObEGMWgnroQg3nAqiM
flYfeY9taISkvkLX+xB7PD2iHipgBaE+gj1S2fEPCjwsdd//X+ndqKA0WT76gg8U
JhWpK/Ji7vq1Nlph6/30s6J9qw2JAmQYEWYFQ/rGrjuht3TObjvnPVpeJC/0OqFc
Vy4lWdVXyVjDyW45KuN+DQdXVDHlYBvjCtVVjZtvy4iiWaSFN358HVf7dbD8sMTp
KTaSB8xcL76ufsE5rJ+PLJ9+fZF9eo9QMd/7faARVASigwWT+TmEFfedL103UpKU
I54gc76Ym9VE1fWmNOLsGRIPY/WqtWHl9WcRrS+YF5w9djFg9cX1ygVVE8SuwIsQ
IEzkcmrW6ibPI3kqeTRgzBjVRYqj0V8prOxWnkX/GaAIsTms6xJD2InZeM7vqcD+
6gK15/iguZ7Svc4t4R7Qp5iPpL58xqo5vkS6cpSXenBcIF/euvhR22e2XgCx4CF+
+Xby+ae0STHn2JqzqsNFRhoF/j0wsR5wmosOnJnwVejK9m2lH0UUv8kMWrP3fbBs
ocYOjGQil7Olf+TC5raaL7mks9oeC0uuu4bpVYBJpe6F5EeDqGqmH3TYtGInMSwe
oi/WGcWrrvjBycp3SoU833eqn/yEdLdx5oKC8Rti7bGqXRA8LcRhMqzHHjaYA/7k
+k9rkLKc+XSB64v/f/RnMaqkyLqTEvlwbBQ4MDuVKVEnNkseoBq4FoIrrBx0rzqc
5Vq3XYtrnZe/A4rbQKQjDKgpLnnC9bMscCvqUDzBmMeHrjAgQMH8+E/qIfEGrPaP
gM1/mXXk2dAz7BuhJPz99p6mDcBKr5CHD9jwTB3cBpzfu1FUeFFSXiQyEbDOq3JG
S6VXFyWqeoZ3OUJnpknwEf2doV6Qg9yUoATGQXMuoPceNDKoNXLoQUE/2TPUPyEH
BGEC6cQr95ujp2FMaR/Plz+W+biIj1JRpZ/qWHmWBlrpwD3Wm3gay+jHH5FvnE+r
Gzn2g0kw75h/hil+2IpQ2rOPG8J0MKkzmZ3yDIvpkd22X4Q45qkH7iiQvGGAPnmA
/TKj1hKgXr0BuWOkZT96z1JQ/BIn4YKBqxtmM657HYomcmCQK7NbaRoWQYY5ldJz
wR5U2vMNr5bKKhyVIRhRS2W9tlw97RAgBEzN6uFSHGFm9lKyOY8NsCn+FzvHTk44
QIvwcK5HqpoLJTPGQAvTRog4NOPO761eyOnEWqNwtEAOSIcRnARYztyXryA+5WVi
hsLAPt69LPLXybIHcJgzis52MKK5sVjpyLGVhdcuKNe2TE+yJ6awW/AI1zbHF94+
kthAlPGaj5W34BhAI00KATx6qRFFW6E+nCXa0qHnzLWaTxNhM+ZkRk347c+Emksj
ujfiTXnWOoRH6Xne9oLGhvxWEyR0cNFUK0grw/nLurRZ1ky3dfKdm5e6egsr381A
jtC8q382U9deVW6141rnhU3+lZsPK4jcl0l8M2ghgB7m1WXY8v1uK/4b8X3fxL1E
1vErhB8dtQoMe+w7hPBDnEKRYdbkzQLyzcsLAFQB+HhiTX3FLTzhhNxeyTydmz8l
tXfS4d/syOkgA5UBilmZ5UkpVE5VYHO4AUPAYKK8Lu+aKRRioA0LxMHhxBtGmsuH
F3WEqdDHDSDv+gppEAhpC34en49zBdNVElIb3sW86eydKXwqYNIslHKITDSCOIu/
k394jCrMwg35FRlOthAL44PCrho0H293KkDLVbMpWWnTJJZlhCvpj9j35peVMAJ7
Nk4+ycFmd+c8a8ACoYfuGf5iHMdsPqh+DmCC/wSwHNDLYdF/F8rW+SC5bZ/91Rkz
6FbAnoI77x6SpQB9zLleZcLdmmWve4RTo0kEN8QVVPKqJ/Mwwe+ypScGvZXXT1EH
GGeVm0EB3AKGBWj7pPGk/hHPnm8BKuNfetABNFs7u+6FkvU7ErGkAUJeTbd04oes
DmxyJAH9bAoFhZCejhymyvxQ1dESdkNkwqPM+cPGZDcD6RpMpqgY5shAY+u/8SFc
xqDZsHiNR42I0XHs9+aQTRMaKptPWE5uTNtAYxiaCHQzOq1RGUYys7OQ3a6J4TIZ
tHr+fbZ6jEm+kwkvGCoIaP6PIyhDlgASVGvys3q+Ko8qEe05YmJ8QXtuXbJessxd
WS4Zx5jrPhdjvLUJqgGqFGPJOUWHdB6I+2X7ZOtBjN2ArmXlP0SjoWj3svtjoesV
FOvUeZBxrFqVU052YuNYI6eXlHQ2Bfi8HvAn1JQ5ZHwUxoVcfk6eM6i4w/FD2sHD
0TB+MlUQ8bG+AiNVYicJEnnHQ1FPJlxnbbZjLmU4KVoZCmMEqhyN1wC6ZHSklOIg
htSM3272Idhxt2GMwR1UvMdpqOLCXfzAVAJRX+66PdeKTd5LFENghA5N3ezGZNKs
JyEFQ6zsfuhKFplv1KydtRZHPqYHjoefgDO1SCVyXydqx1DbNXegazJyWNSRIL6J
rSTUxvmMTdlnCho192GuI7w+5HaS7BMPObtpXYvtgzJu8IhSSYHAozfOOzLh4ZG6
zUWTVrd0axSjqSoTKZT38OVIoSZ9/iBXFIh1D8OeJuSi7DP9xUYKfA5FwNMmSi2o
nrOgLbJ0Dx88lEC+g2/9XHn9ubiNET/E9lXOTV7yAIm/JjK+EDfgFdh1abYMnNVD
ge5Z59INKNEK8I8xor9s5L2dvlesHuoSbEjvSq2ZaAOsGochjHqnA3Y0OoyNAyIJ
7QRWM37M2B16MQwW0c6y/RR/E/J4SQsmMdYUXUE0b6PTGOSUcIn9sPQJAaowjqv9
OGj4mY0OiXuEk2hIfqCXplW5aPqXkr7cdJ02UBeMQu7sdNDT+clLwO2MdLwkbOte
IUMWiGSoEIMPSJ2bXFsHsHnahHBsjKpZLsOWFDOaLNOicXVAW24FxkWtn+45mRcq
He5hmkTJ794hFvnm1azZtGFUb39zyG8bgfb0CUSKAtKzcwKSwaUHr6Kv4XrY0w2u
cx/VAVwZoL7rDwBZwng+HAn/5Wztn6o3GasVaZafD3uGeWiCwxOA94pLP4QV2gKa
1BDYQPb/n1vl1GymJpzNXohGF+XCrFlQHvsHFAIV9RW8/0KbmmDQubjWOHlSCwGS
q8YUh/UQ+FJNX1nDdkELRuCXxm6i09agXgQZBASuvtkHFDtTHIWQyhaoQD/Gp17T
wJYOazu4D/blb1lz8M5nw8Hfs8Msc/CNm0UUP8kNiWP2/fY3X5SkguX2mYMN4wNb
D9WLhLsMbJuvS79qCo5Xde+/u6+yuu5xUoQ2/ufMeU46ZHVybtbUXrHTgn1HTVQX
0HW5UfLSurmPsdJfPquezdsM36JUJhm5cYWBMi1I4qDPsv5Mmk9ZCM5wuWzCYBXI
rotd6Dga/w0HpAUb2k9YIIzymWi0zU/lLzAEIGzqFlw4iZRL/r/5jcaQ5wVPDvIs
FdbT0KjIZs/UMDe15h7fZ1jRqC0JzZ/o17W3tiwGdWNsY3rGfi5+fMwWnoDS1TEJ
j/mCCRs2cgW+dn8Wf15hV0vB/lKzfhG59y+U0g4CkKtjMAQo6fSAnnw91YUcWuzy
OKtzJaxiRR0iTICbxPEclKYkgGL+ler89/QNC004Bi9Zhoonhmz6v1GcqgunVOig
vuRIRGuk81xxtFpUjrcMmS0ltAuz0uvmjBvxw6NHugOyq2CFg3WH0Ryc7zts4UMY
TCbR9iXLVACRyluDbrYLcnxVkhPwQ2BqgeDDvmfjXcYXSl3NungnzjvF2Rwq3oGQ
bQxEb8o1TzCBb0QJh39Hf0q/hQPsLtQeme5D8fOEu5Ee1eO5XElPPDCmczwQB6GU
LyQDZXabDueonusdU2F6NVO6T2YW53jqFFZamExEG05ltO+ezxT3MehyWvDahXAD
jhuT2C5/kTYaM6jAlxFuFMBU+jxRuZ4rP9We4c0SLaJmNigDn2rbvjXJPKMN5c3U
J1uV2FNB6/ZG9dRJb46IsqXI6ZD+ubNm7Ws4P2GIHYkljzopZTjZfqI1iMx8Qn6r
EArgeJrugPEjb/3dvZDjym+0ZMk0nHHWx2tFD2o3jhBqn1mNd75T80QfusOpIpEg
wZbNnA6JPIjCkJBeoXuKn2+gKkh3eGVM1r8HrgWLYjluVtY7R63FUZdIMwxwggJw
vYSDM4UUPJIxGN1f/MH3EEC8abh0hH3udTWfm+Tmm4xSh3RASMM2SmPDJUbnOfc8
a5Kj6/7Rz9xiaakYMoC0071cL6qQAbfabTN/xzCC4hM0d+Af39fyHorZKJs3HhG8
Ansi2gwnuLKI4NfHf7sdjSTQCyyGxEyABmxb6fZe/fhbWqrF49Flm5RaS7MVtL5y
R3w5xkCz1tumDzyOAfZD54drV4ALR28tWslO0TRakg5O/Ib6R5VszRIdPWWsSdBe
6U3U9djb7LKlXTksbIpuntlNYIEftRJrp/fRVioSRl3Bu3wnVA0ZdsiwZE46MTl8
06CyRvB9IIQEvhjvfHV9Twzg5ltel2fWOVoh9boVr3iic54Ztts+xQOOK/26kVSn
FgImuSv9LsCXXJQrQ9aHk7LSPdMP++Mf3wqb49qw3VWcxQW8BRJ9pco6+0LawgA3
wxoN+Bt3EEzN/U1istCnrIt8HhYADHZZ2yo60E6miRcWRUl6ACodNkU4YP02o1jt
Wxuj+V+z96KgIdd1NVYPbdysd2vDyqpkfj9n4JHj/XjOSVoa7cZdAbcMyO9dCVqM
qjMskRJRTWp5gurIclQ5qBeUwfaO7yAHyqQn4r6gXNtz9NnEBi9QBHNtfIwakURu
TCt0UsMY1JFhr5uKg8iVj4fFhcd/BZ2/7lChciIJC1tjHUlaaNZqJotK/3hBrfdQ
4a6wubga3N3c6qj2JmnA+x1spSAwi+Jr1Y/CHDLUC5o0cqQlw9FnB4oQ+4X6UKrL
ZvdF+z9oCWvRbcZEquXmB/7cMiox9eKYpF2s9qqSWBR0voh/sN89o/whtgLVD1F8
PqUgdgOUNX3ZlP6xCqXXu7zHwRIFiYUBxLH0IGKiFr5bbCzvvD+Yc3As34ZV43O3
hZEM3x0iIZEl70xef+OW7vjz5RwikWFogbKbnYqzQtglCPpjIwqnB0PfqmcjBcut
r2uCykllcvIYXa4nJ30nb7y428cQyB3pDjsdqAaqmQ60r687U4StIbEKo4e0Ubi+
vgfBcYw+dSzqqQicjtgp5G4P9h71aezTxdzvMn0rWESsMFENWqxEf2Z+FZgjcXxx
cvCqpvaOHtp7WzxV7nF5XewEEJKHl2hFYYnUFWwRKGYZw5Yw4q31fYQzzRFxkQq5
jQXZF2UVUmPWL8YXnhWfogvfjCyqe+Svh/on8BLOrMd5qzGKNQ12wVBZJtx3zL7M
VZXQEqDHRXuPe3q244NijDayOxmvtf1EYSD85Wp3nGv1vAQEljZMk+w0n/9fAOaP
fnzFngLKgn+Dc9ZoKWkaOKGE5nDv3K7XlOGO2/8+2s2iJtQkEng6QPB1Ixdn26sk
dQeX8070dGbdsLqadio29/y4G8jRiS6rMTN3UYEbHvuZcC1mmULJJ3og7fWXQx7Y
afoESG+tStED86BcSLVYb9TfJgCPrlbyMCXCKRIh2tIt5HDkIDbQ02NoRVp9Z4Je
8TwThI+Ky/K5cW+jd1wxA8Om34oMrWHAmv4MDd2zVkmPNIkqwvyvUY5x+ajz2rbn
jCJZw8ZwWcoQgUxwNrVHfBllBGMShmFtXp/v+RzexTOflLKTT4b+LjhoFTzqexaC
D/07dR71Lcwn6VUdRdu5SIxLU8HNTegyG4gZ8cq1VJtN3Q5Np6pdCHgnJWuM0ulJ
Y8w2DxyZjJXEMooNgTK7jauWuZ3lJBgwKchrM/aUH50z+ZVpRb14+si4Kh7aiDW/
iA4YAIlG5kYeSpSW8KX3arAVzqRUu1SmEcDlgcnMj9e0YA3CL5E/ShdLMOGgxx8a
FCx6AyxR1iZRLySFobb/+mh1gmSLi+pzGIIJhEl9cC4+2OxQfTbvbvU4lAG1smky
OAtAKVnUcuNw0rdTq2Ub8lTabitc6iMq9Yd6GBnNAGMGKdkRSq3nsd3dSlgHgki3
SrnrFNYPzidCilR2TN7ZRnZ4v6aS6GHJsHEM2oljrZDJTD5pRFpHr63GOySdaNWU
WqvbX1FEB04R67MFUtiBd+f/2dzXMUTUjdiO8iwPWt9HgNoQwa+w6/Day9U6m9Zo
UCZyREOHW8BxaArzJHEvwvRwp45ij4N9EInynI7nED0++VbXbFYx1jikrwL4GUTI
d/ynTEfmi1m4lI0kH+dWNIMoqltslcNvhOhQ0DhkiIf3FMLy/W/duNFYDACAi4yG
pjT1hfbR3b04uGrjcG/9avFUV1iVQ+gFhobgb3xp3byXJN2jK4b/ddIL5owiZ7vu
cGCumVZ/scK/RoMuak5yA0gp5HZjH+NUas8R+EQbdX/7cMVgPYcRdHdBxM4azlTG
V0lPhm8D5m8KUWoqL7+xGLAvNqJYyWquE5IZwrxfSHnfWKG5OGmy+OiRUtP7OTbV
mEyIsNe8CVxFLZW3LU9Qee7S5EdT1KIl5wEEjVaYYzbT7PjlQmkPUr+y5ObzjlNl
0BSOzliZknnFqBP7ywcbsnB6XSP9iNB1aI5f2NXKPEhKiVd5A71WIdlwVFGPR+f+
vygGl7LhmRcMmByf1lCjwiJXW5V3zujUHTm3fEgKBMFVKqNReTFo+GtOdG0QpY3p
0qOBDEUY65MBoIrIbJ7m1R6A+sCcQEwqtaJ+xkqUOwGxYzxKU8RKfk/JlMqjSSIJ
p6hBkGQgy8+mXK1TQkHRtssBPMTrgCVxke9w3yJGy7ULHw4j5CbLsEZK2cH+8rdA
kRjaB/fznhv6ufWRy/s7tx0Yt1v7OzEpZz6L0YQsWY7UDUMGUXpqWo4t78fh9Q+K
r/puNCrhvwucSNyLp+LTfBTu9vj84z3kU1I3Xe6eiV96NCMRfJDllqoKS60TPK1D
tE7IezJVl68u8PjpK7LAJ7V0LQdZit3Y7OI5gR3o7JDmILfbJWfGEFYNFQ57/xgV
R6fFJlrJ7rjSLY3/Prd4z/cNDfcsM4ziiG+NrBVtXMi1Gpfb/CUCxvlNRIBwSuRz
bO/UHaYWovPLlTLRR0lglG/MZsfMn9xdPs106lwWlVwjQv/pfwo5X4eCG84p7n40
FRqfUa8MGhYEaORKNmMF5jcqCMzND9cC1RJfmSTZ8sZWK7ARApRnyNpUvhT5LVgX
VyB+bZHKFEA1uGsMucOlEqIJN2Acxiu5ytM5vg9LILCuEAeA50k3D+0LxvZKPGrO
R8cl7bzvwbFSdlxkrkIiHAdKiCe83Cix+ALP4V+TLZcPCSjJJeKvX1l9mQV1/f6x
ZS/M5brC2i3izphhjvrR9vsO69egxz0KvnYg9bzHrmbYse66dfqILnAUFYlkbza1
YnHAXAoGubJNRAOdw1bKhA9a28j6fgRwGiTS0fBzQCVlyaapQ6o8elDmgSSuSPZ6
IwLHA6loTzHics9DsJzgIchDHVyCs+MNafTW9S5pYyOqRiGCEc0k8qMphzA6UUiR
PbkLEHqsYnhcu6X9OOkjF14yxMVKWXL3d8iCo5X7TNOdTUD/XLWWDMqBPBHB/Rsz
B2Av65GbFLcNJ+PY+HdlWbyOTlxKQxvbkZWtX8KNi2Nb1zNkkhECcknZLu34m8oO
hhLiV2gg6OFsjPW2jN4E7buq3v2OklQQLj8rOy8woqu221wgeRdgj9XJulFaMaaC
Pab41AlkW8TnTWPBz8FZa71uxQRkwI1UcJ6rxuYevFu86yypLmPc/Z5z6wrNuSMQ
20EE6f/vEUUrJpG4DgQ1+4xxn6VNseiRkkzfF085gm7QFBzkrgWikRuo0tS/uEt4
Gc/l30/3IW8lnRe0MrR5FfgCSOLQfIw4R+Y/8VrJ9JfQ9kZTbvkEi+uZwqRkywRY
+BouRTihNnYFrmj6tVYVyU4ljWSbk1e3Ap7/Q5M1cC91qKJt6/Hu9PzauXNdor1A
deK4Hla6blg7T+Qn/BaZ6mUmq8l2/4utoZd/ezJ0qz4NeBcQTJkX57CPMvnTrnms
TTl3fje1zyIA84r/sHWzUALRPQajCSSBi/AVfKOmxQ/vUVDfqagosAFQmEl47Kdv
8bov3+dNcGplg6WY3uiOHMBp+XqMeZ6pZhZ+lMGMc7OhTeJ8KaTM0rQRtzXEwe+W
Yn5wZESpnWP3ikAa4ljm4HdSagRufo4cBdm/Ix0/fGuDnGhtmzdWw+AEjAyJ+6aj
ui8q0uHPt0s0dSisVL5bbKBIYQNPNEvGRY3q90rc9eQwUR86/1RWNfwzvViKogVg
Z4m4m2ewW123Jues8vw6SWvAGa1HwVXzODcArxee/02dAVlZ5RH7h33V0dc/d5vu
QLOAJyd+V62c03XABV5dYAwKCHx/Ybd6HZwQa6e7sHY0gTDvOsiwSr0NZUegFffs
0jzwBy1kT8gm3WGxGv1nEewllPlRhPG/i+fQXbES8bSHElNWuZ722kqx/oMEuHId
KYUED6qnPzWLglNkMerLO9I15Qnh206/avTPt/9/OiaVXHVINBJ47Onvt4lRPAja
B68VZK42x0/rA9Fbn+rRTa0fWR/6HkQ111npHj3zAAvApO7fA6QnxApKxExdt46N
cr+Lb//wGIIb+ibCBeg5OBKqQKO44co/IHkxmp9dZC51DTC7ry96gRJSn6yZMo5A
Hz2vja5jGONk89Dd2BI7teaw/fDuflSTOeF4pFrWzN6vI8YVXmv5Gui7z80XUkgf
8Y8OSLHuf3rkf0z23T/tvAVxUoETjqrn59xLxFeYQMUT5Ja3GC1GNQLDK6uhDhST
08qERAy66xqMwPkUA1ksNjyYBVjZYPwuAr6shPeVQgPfy//AZOKWtyIcmT3OfOjX
7lq9EXjQNRV6R6+4RBOp7C+G+p4kU9QzW+2z4LA+c062nOg09bs8Z/QdBpgPIqjO
tC7PkTkyPmbysInPVKupOEsj2XeWk+5OFRfgFEu611nFxSZoJkDeawXvGk5bzHEQ
eBLMducz++hI+mZMstOl4S0waIR3De2WqNsKFuScMxJ3dQIPd+58U6h+qEWNd7Pn
GPhXVOni1O9YIpS8myGCdAGnFo6oen0YzxBJdeJFm/UJyJ9Rah/qM6aw4ePnpIvp
LMEMhwckQEHELMTxYSIaD98pHsSqp/isgLiRbGYOREMQLJlQx0669sPcq5nrf0Zj
xICNWoBwl5oTaKouxtK9K3OzEP6/ihPsfkr1dmQ/z2DclbXAgPFWsqSajpi+vEgN
PlbKCKHtWmVwYpvbWSc/NZYm2oNLufSEQ8gtuMJ3lXuaxrrALMmTHCe7P6JFLZhG
cWqdjFa56YH9u4+mKiFRveOtVyJhuQDc2kfWNJrZKPAdcU1rbAeFsrV9qKnkAmO7
zZfWNoPsxcpRQ1VfPcSed1mgTztaHBKcTJ5UP+ALGChfDIVnIyEiP7oXdgBqIr+G
vmFfGIEior9iMIdWJYcmKm/EGqijlPu3bqy8G72nAPQ6mlwiOG+WLJydtwAlqrMe
evtOOm6CF6mDWB6oLKHGOP6IdQVlNUjNpYgTw1hLTvE/1FLOwYz89oQO/jjRdqd4
pIb1b2eFdhYTNdVfRHxYBL77WCBvYLF39cmMjWxgmQONQWBImekrbWGGp4aYyybx
0lEub0j8KAiJvsJBCAeYbmicn/4IP0CnaOygDDoBDUIc0LUPRCuo4u6y4grfDY3U
zy7RzqhAwQybXlY9Qw3cG5XpnbKEpUtmdlgFVpvfU90zwWgR57G6+zcmGfvL9QnK
YxkfK/5sHrXMk4rrQs1G/Dt0fsFHSSg5WIUXFSB636gsEMBDHBtknfpYM0PyTz9U
wARRzg8fbxu+85AP79uMjIfaEOqUIQ1cegmLdlIxpGgrXERIc8qJHx6iiy9ZrgNP
9KGfhGLsFx+jDBoZARZG2Tbu/XvOx+FWvAn12nSxY5nJtgjoovl8NCDA6VidPO/p
TQkas3XzZlKyVER16Y3ZNrCEb42VJChLrM/v4esCTg8j1EPV04zLZgzKPeEuBnbv
GQYXGYNTg2CP7oDw+Qy5tIFm5aU73Ntq4HOs/sRLbBOIVA0WyR9NGc5Z7wB1SqBJ
g1p+cMhnxImF5Sco73oxDsb6GmsvjVCSn1HaQCG0pOQwWgYm7IJ4TfR5WPTei2KE
6VxipcFhlpIoKGdtyvwEwhxbGkFVlFavdcwsWHwIdngFA/FhUqDpoLVwksZh+a1X
cmwlUL+V7lt6atR5GNtpfoKrGqEDXgy5+kMgn84GqCxVSdQemqt/y86woIrQg00l
HdAgUncfmFIOJj8gfraaVrZi1vEzeB+VZ/qpGtkN3PkB+E4dTHthrC1Cwa1SpLcz
SPztWP/62q+ckiKDQluQJYjJBA2g34HAQ8zLfeA1TKBA22Qyj0ymD0KI9QXvGmKP
n874pkRNg3SXNhfIEvrkIEfu3SnIDOqWIXuhUvPUfQW2UyQz7YOhjZxtuVQE+xvk
Ree9Tzo5u0xrC95ff6oQb4ZC01RdZ3Cxup5HUUvPZeVOHB0yGGfSjBk7xa6q50TO
oW1rQlJ0v59qzOTGRdbMQCWuqw3G1I8TVmmT+WuKhcZkhZpY16dbTOuYxNSUA6yf
HL+t+FjKFwegrwA22/hcJBPYLMyAEMHHaaIdWZtdsMdOEWjM8ib+/Ji51YKYZaJr
TQyfFsesO7LYNViKoSAuFssq42ArqMpI+LcsQljEQ9OJ19enL0kMVdIgQTJ9GGkT
0jx9H3NoJjdLJIljqf8JsAsjRLFE8j1K3BKxguJUaE7Dd483A/xjWseIkvy91jE5
eBTq6K5gE10Ytot0xeGQHCNjTjj9lyI7Gs2YpwrqbC/f//UBg4/Oqn7eQtEfMlFq
r2dmpaOD3XT1ao15YuiIZULW/3icuWq6C0zSNRrCCueOG05a/+Fx0HwU6wa9NpdW
4sGy1UkItD98oHXiOeK3oh3TP3krV1n9jahreY0wTwCttmjHIXbPDtUjQU2N3t0Q
fFlrKPEf0oZ6H2WlgbAGjjH7+/6Xt00mCWScfaTUlroSBTcHnB1yeMOlPG7DqERI
7ZvUmfW5XoSV98wJyQ+L3jr+445ADqV4/nANuU6zEoSKNusss10NAosOeMhSz1hY
dgl/VN6XUyUcOVgeTOiif7TORPUArkZz0r/vJMwjCc2hVHXbYgEVuvX0zqohnSzy
WhsGiXQZL4bJTaomLDjtMYvd/l4ctJGjjb58qZHYtQBjNxoJW56X34x891Z0B2m2
mvie1Pvw8FLvwS7HQQsWa3KUyxih8x9joCpOOqAejE+ZXhXhCSK9ouuHJDpN37SJ
MCoszIwJE86WXjNmMJSg/Tn6GQ/48xx76dMCJYBi2IUN9q2ch+zLf/OMYGkufFw6
yVO35Iqu8W/q8/eu8ksr4kZ62tuESpjSSzHHbNJaaQPOVMkLQw4clcnU37ChQlhG
Kr1vlmGjc9YCqznHCDSsvz/8qYZijOK6U2/BJmghVWsIJFmJVbFw1eJ9cOzTHmH8
CefeD/eFlAiu3vGTJlEpOE9FKKCbIlzVGo11HaeJwiP+wMCLV9Evesf5jX4hzsN5
ne/uuBFqmTTehSral2aQuN3EYQKs7w1i0LRhTxZENB0f8F3hD9Y86eqGwFnqewz/
a6m7Hm/M5vPpzsjYHORaOMaTqH4yCVV3YLmXL6hkHBHpaCvgh/KKn/rooRokwKZQ
Sx8JQTYA4iDbznIBgOaEovw8arsrwxKGLoKDDZwiNG1NcZPIZKQOkJBp5/KNtMGr
QG21OCHFkLWCww4fMS38cuPk+SNfKohFp5ij564Nx1IwvJMxbD6gdhLIAz4Rz9T7
Fj1xXIOWBSuggWpJ2EBn1x+2en6ywcvVG5ycrivv7z36X9AiMrXqWKgRYmjoAZzq
J/CN0SSONukBOYNLUeI5VDE0DSFNR9MMe7/nih2x9jw8Mm2sx/cewNh9yBy4+4i/
yPyKJFxv9m2eRV+KCdIhw6GgXJNihKS2dE3h2PfFaZNgiwSaLduijnFXGb36oXIa
sszEkSW1OxfOhhcIrl+canBRbd6kKLwKEiuEot1WJ8tJWJoRV36TZZfIsoA/dMjT
z1wQ0XCiYIlOh78/fJ0b3xP8uf9WhY6CC5ezGzUZfYuj/OTqG9LZT/lktUtMt1A4
DouKAbnOOv+iMIyTMI3QmA7AAqbeSpsYLtZXmZs0h97xEZbdH+iDo7R22ZxHz/+I
A442l4sZV52fyKN3KJsjxzbHtfIxqG7tgxuYw77Q1Rgn6xzoVKr+/cEnCoi4vzY1
e3a2LlhCCV4Kv3SJvc3balUl9kDKm1WLUOAfZyF3R/X1BLJiihIN058nBKiwYZwr
4LMQdeyenLKZoh/HiHM+MB/l28+GVmTTFeEallIEF7VunxAJ89C8ZBc8IGgPpNqR
LRtj4+WdlvYvTpcvDKVXhPuuOJ6Gvrc4/OEvz3LCOrSKPz6UxaHtqXE0wpftUk97
H7Sl0CkXvvq6WUa7Gp9eWeC3+C/a8gnT9TDb/If0iri+ZmnNRD3GRinVeYn2c50x
zI3aCudraa+mhqDdFYEqBS7QbB4/Vj5TOfqt6beVleh8IKH7Hhylmq4qtbpC7vj7
BKcNbYBtjrM+84u2swiZMvFcCIPxj1dGHSEj4MDrwJd3Iy4ocL6TMfmry7vaXqC8
amufbEeuai/hdMaJRddo3KagthuKALeijYgE0CkMBCDIixSYD59Si8UEXnR3mIA2
om1efwOvHwnPlr1y3mld5Tp5qQh548hFbtNQTBjxx9Ei6w63seNSpOsNkSszhqBp
6kUfN9T/P8yTt6Fr+4Tg5piqUYiKAl5f0z4s5f2HPxjr3rYpzPF/u2Sr/Pu5RZ2T
hE9R7cEuP/WzmC4FXZYTiSpfrDw21OnKCPJ8yxXVg8Vt1hZe4su6A2e4nrmytVoz
cVTOpHgVagPRfM7infKezuzQjorwxvWCmh1+ygSLH/KfG71awE5ReWguBPzgZDca
g17IXdp94EeW6RaIe8uM7uJumF2oCLPlbjuNqmft3I1ri0ZOoTEPqWd+7KgdZBtt
wkyJrYuozbtAksTXqK18TklMVUSHCiKe+hvNX3fprqgPeQBP+ePFi6YIf8cTeFD/
uAqjLG7zPetzy8txHuebcHuJLqxu9ov7UM4gBOmYbrRrPq0A9cQcUuM+D4VgomNt
LcAuaktTrlt8ZnC4UvxMWUErcyWG03kZ632VEqmGZuJnv+P202WZY6wEAc9R7xLW
S/QZ9BWC7qlFlqm2g0kLB14gt5Qyr0Wi1PshpA9vfxOFF/ZinILWZRZz99FMwWIP
6LGl7lgqYt7hTIzrB75yetTNg+xR8L8eB5IM/aYgomxj+czDNTPwkaS+33G4G7X0
6IoH8nVkVIkYdCEEu+C4oTcWrFBajWY5vcLnP0QVSsIf3ed/XDEKU4mMFOwzv16u
2iXWt854ekjdSjkiF0Yz+MJ+wvrvqGK+7Jo/36agQEmjxy9EQ52bn5YYEx6kZjod
8PBwu7cruzyJgbn/y7tUtk2WmvV72BjvZ0OgcxFnAgSZYsAFt6ewiiGGjH2mtpqs
/FEltzm9YKde1kINWQ71Pc0vkl41OD1wdEcMNtpSwpeWBtDX2e4yPyNJaIecMtgG
RFBwSEZ3XlQ5jKuPUQjxHPzBLbDwse3WTovhspFyAFI=
`protect END_PROTECTED
