`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgQ3fNl4QDVzBA89ziZhb8ZBaRxI4YOWEQ9e4luWWSBOSBKN0Q3Z9uoNGzOwifen
kps7d7Yf0HkGgIe4BQEAh+cW8OiYvHjduw0kZO4Cc0xF1YMXqhjmMyKET3xpvQGl
oSASaBv2jRwkf/UvAxjLULPwZxi56alS6UKq1EtA5ydnRMOUxKx6pETV2muxpf/G
AHwlnUaP0DzsGMprpgO7Rtr1iOMIM04o475bzSly+5lsptqTISW0MmLccbiNNtLw
/cta5tZ7sQyT1J3Rs4Po2vCJofUxzmKRCFX4z1d9evgzTEfWqHkSH9MZJxxyzBmE
r2K2CwzzOmcxZhzm1gxB7/q+PtGS6qeisL31o5JgBw+pIsIf+Xu47Ggf0+ySXWm7
BuNF7jRBa0QBg91UnRcpY8wQzSBwlKk+42Kyb/AV+4iYcQLbANquO6SxAndTV4Kn
gSv3L4HmDD2c4vMGSz3qQw==
`protect END_PROTECTED
