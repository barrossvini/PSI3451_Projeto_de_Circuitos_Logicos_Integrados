`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cvnGi5+hOp1kytl6jp6xnG+JFdRwpiyNFrmdI5/uRQa8X3GzS+uTCkxee3BGnRn9
J1fLwsUZC3SD7aqnJOVE+jc9p+s96fdOS9NJ64ALFys2pmFcB1XLWQ3wMQEDhmgT
M+b+/FiVveTTAlG2FPjVAG09uprQr5Kfii242Q8AChbOCoxl3UeOj+uli4/I5UoO
nGX25BzSRd6TZPyQkI0EVHYiiP/JCkjElZIAzTvmVCCGMThT+WFyUR8NfPy7/I3u
1S65544eM6bG25uH5EOqfq4ZAB5nMFZIHY6HmybM1J46xeJyWyL+FygaRvVdNVo7
O/VT7EfROd6qen0AGJiL/5A4o1fq6AaIge7/+qOwjI/UO9cj+piGzOir/20pw16E
5Lp4gPnAVrvIJtGj9RpqajPx7ahuHij5r/9iL9aD0d5h3BERNMVj4ZZcbjbywafD
poyIH3VQX1qU1zu2kznDHvZ4liaj3m4PRW3l5et6B8ewWS6B2gi4TxQjIMvBiKbE
e4vpwXV1sGBkb9I2tucgLbRcNN+ayq8jN2YIgflmN/iF+/gQ2FVMwAYTNKwKkDkc
xfNS+mHQnW9f015Xkn42W2TcrhgsaOThytDQRo2O5gPA0n6RJ3a3UNqzLMdb34Ip
YIkK8ukRNr6HTEuW69aMbkJqgENLo738Fx/SFqG3UytT3spk9GeMMHKJvPkj5Fw2
s/vZuKXbGmPpC/wA71tz2KrtIQceB74n/neEgPsnqlnYPRSQVGjXK9uh9tjDk9tl
rFmvRowf9IYbW358F3Sx+MsUl6twLlRippf6FaAdi46Oa58012ViuVM7+uBFRQr2
GLlmhgemPj0hANtwKK38qMItBaWS7PkUGt9jVvd8kjD/DjY8FnuT3TMqL7Nd7yeg
1QiI8X2P71QaHQhh8VnQHHCsq9obn3zs7md16XPvtkR2gl8t8z6yLI1AYJmUKJh1
jU3zrtIFGJWOuMNoVV/telPjxRxUl0mpcUqU2xfkRQ08VOC7rDs5Ms1fV8RtwN2H
qR3aiBXDPCPd/y7a83Wpe4CJxdj8dOJqO1ncxmtSwFdmdbrYSXOvv86r2kTE+opZ
69RZq5uAvNOznzQUAydEuWT61N1jn0R8NOcdgiJzEskPJAOI++T0OdPmK9xpC6uc
+YX2wU+sACHeoHoSqn2EEhK3KcgXiXHCjcHEXCoc9bf7bH46nTgBsIHCQnkzg1bS
4TsP7Vs7gxwE7Qc6mVNJgtZSJIvJuvkEJxXkog7q58XPat63Xvl3rmlijDyb1uki
nRVvkpG5vl1WdK0ghI2Y5avyJBOZKgtmK0eBqIv6qaEOFQLC+Ti3GMpLKeg+Z0xO
LtsEjBofiH3zUXIgrhb0PvXl7LQPCpOkpHjifwNw4z9xQi0PbnMY2OUWY8Nd00OG
kM1mDL0G0dHRxy5gV/UTi15//FLRKAzmnk0NjC5lGklP0RhHVM1mIF73yLzA9Zev
o8DdnCzSzf4BI2hFYJHEsRcD/WBuPChVWJH3m7/6yGojR0xOfJvCq7Y+bruhwhkm
Zo+iEQVF2kwFs1F0rhlJv8UXow5YWq9n++77KEB18a1//NSMJrjas6QKACNzwcPj
okBlozMa+frHfmGOYAnFsyzFqCa1KtCKMWikVLkp4QqiKNdDTALc+M1mqdugXLKv
xurevmnRrfA9Sr+L9ALqVNggZ3HICpcrysMuw/ypeOH2WLSOaJhJQE2fT8GB05XN
uI9FKno18KyqniHDpeaelsA4KpuMQq5CT/qAZVDSOa1VSIRnAQXEbncnf+eAlDry
UCNkHLswDnP7j9zE04WbfsRJiBHDPx4YqEAzAH5Bp0YkhvlJn4LA43GDg506mObN
MpGOvESOSw/SQ1esM85QgJucvtM+C0ylWjtCS3egiz1IwuqFVRz/odC+rq04iukC
+0086sqO+DSo+zraNw4VRCWNipWP8JGeuARWeMX75FR8i3IdjDrhaNXmAv7fRPz+
zBJsSvuAwWPvHkKSCY39dJEe9dcRc75qpXYAa5U7ALx0pMG6ATGwiIdD1Gu4hRPn
KhHBkf9zzcXDJOwgAXDgGxGDVmbIF4XpUE2rHt/7k3WcHqO3LLw61UEHicUz8LDN
5YQlGudpk5QP82HE/vGhT2IUGZCu3J1TPsETa3IZjE6vq/hK9R+NrdTPEEDzRoRq
mKmC31Il+1q4rQA4bFPc9/b2GECpzmthwc+rTGAJd8zLpQBBNmZeDKtAyzzRuThu
85feKVGjF0IEBgTm1AiXMmpTcypv0oFoamqDMEgLaT9DJ9DKF/rRbBM7THwggJ+d
S/qaFv5fpn07bDnAVsdadtHZYw4W0yP1eIH2AbWJ0MEAEn5c1WBxiQ58ZjtTdUVv
hZ7z1OG43gL7tbtN+X56WtaWD+HUkMpVlxNHKAt2dADJk/K4dOUQrkSpIab4WTbd
hdHwBfB3tSs2fEuqfYDdaPTUcWEriLwhqN8E3sZWF6IVYfnUkIF3GRmYo73gGa/K
PpKFeMf0B141QcUWCaMlUMqMCIX/70Opsb54cHcppbFdiUQD8icvmbohg5BP3W+D
fLdtjIy0uduq8bVjLMikCDsNQFVS2X+z8eFuoYt9g5KeQS4FLfJmGyJkhkUrT4DO
sT1W0MrCo9+3kK4y3O1UAcemQvMSTftwqdQAvcfFkNeyzMRr7r4otnS6O387UuoD
p7vp2PB/fMNQBUwq9w5/oUhZ70x7qi68Y4XLKsxjla7YJI498BBimyZ1L7hS3Hx2
V8Yxfuiwpi5e5Q/uEmsi6111JxaW2RLPS+YV0qZxIivjSIQ+3ZIR7q5ea4ByPzHH
eyqfMdZw7JWA6JuFXGNnvOCizFwJAXJGygpRfw1MRUeMszcrRzuX4urwrGAK4hNt
eyvYXFNFj6gw+so/atuvyQLwbYNhkX07CvVYdTJisiVIQQpDlO1Q2kghnfYKasIb
D52hlwqXQSJaEWQZIiS1Z5W1Fn1Yb1UuD8PaFXiruJk+8m4km/fkvB81FLi0ppUF
CWKKHSG+VKvVP1+OSO8y50l5LnHffYsR+wltUh7+m66igp67CSH/TFZvVLBSfqCP
Vj4kiHF3sPXh+k9TI31eaVMqNj5J53i1uwIGJztRS4KPQORCZWBjYFUsxHINKvpf
ooP+h+BfSy9YoeUlMrldmq6DgSv+bZlrKCbl0QiXwmfWlJ7edGtZ4KL1fBOO2GQ6
gd2kHFCBq7nbKAnGBpFiEcZvAAMktu9KKdEVuvUJCsKLI20gaxWzQF0zeQ08Hg2y
uRLyjhFUCGlrqT5GC4Slar2E+p0D3BbdPYOEue+OEpDA0yuJRt5ZVYVrer8D85FD
6aipD0dKjhtkKLjTCMI+v3VqiJv7OEMo7wsy/zOzmcnExUfA0YGYXEq63SmGupJB
OvqJ2RaPLvouIUggmcmdxkSuH+RtRL1YYxT3M07zl91P+3/Ywuz/x1pDt6aVCvAg
s/kJsLPWZfdEEZvuV6kZ1EtUdfqmSLYd9i3QeL1lcrnO+NkRQDhrwCMjpLh7btR4
RL5srpsHWk9nNjinaOM2+TyjouN7x2GeqeqRvlg3isEcY0iNP0YuePIV+d/Nz7nW
CLDubQCMRv1aAfdFAVTZUF1RUS7mfb+E5IcfIgVi/DYSPKzjYb88+G0nJ6rEohW8
`protect END_PROTECTED
