`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
juyXuqqEKHNK67eQn8tR/Yv6TdIHHr8Mm68BAebTCRm8xqfSE3pfq9e17dHmS7Zn
7ZKh/aOWNBfmYCJIZvLjoKg1rGTObXPo9hHNcAPYtuHNpEpD6CTcvZ1YOaC964N1
qKezOcpda2wi7t3S5G+vyJdFwYzCO4ZNQvpyCHnbfeEXvi8t9KNaGEMA/YrKLeTR
Ff6tj8INgNmw8LAf1HN3H3UMBFtmn1cRdsu20fqP61dlwj7eLTsDtzpbV8gu95nn
A7SVID8vgJ4pCzqSYOnOFGqDGcAbwiTu/lhsvNPybGiw24aK1xg+yQcbhpwE9/1W
VsJgnywtqGtoRZFBltZyf0vdfWxiMVWVwy+Pn2YIDb815BezvgUbPgkcblfAjwcW
GlQAabRdJMYar9latjiQ+PcJ5V8vvxh1frZEYG2bQTLXn76L14HWaec6IiHQpWc4
eQH0E9ar9PHmQzxFtjlZwCbESnnPZxI++8uXo10Ar4m5d6w0XuebYU4OrQnbmRsl
6dSZmSiNyv5zGnfG/ZpvBICZ4rpit1Mzv4GqwAhGATloQdKO1kBXPjradRtvD7OB
Ze+PYQSJAesMdM8Z6AfekPQVytGj5kDN1cX41IiNwSK9a00+kNrDPAEkX6FQwz8q
6D20J4L0euvFfWZnQuRInYXDG7BucWJvtm+x46UmJqBarKAQDCFAlN0PqrDKh9Et
hyTfc/3e9rIjiOhJD72iaRqFaCHgsTAsssM3cH+SalyaBZ+50UYB9o9EYCRakfK/
25ISMU0DX2T8WEZ75T6sw2+kqA+dCv79RR/NtmTdHoE3vBxGLUYjM1MoiMvMsvOY
lNRenbPJd5JCOFchmRnmgGsBm3jpjEw1M88g0noI/+7UIRYbJ5bRrRSCebF2xn85
EgKpRCpNA/kBrsPLXgV20n0hR/jLhGR97wcHsMdaWz2qGrlpRfdufUIR9oaAJC+q
mzPZwhXNZBNRqedeLpRCwnOEfNJbCUP9A0+iMru+RLXRu5VnBRUEIvlCeJaTEBiM
718yOc4PqkZNpwyT0+mBdt5+BqSQPZSpQ84vs5lRIivRE2DxwMLFDiLIvhgt1uDi
oqxICnhGWY/hb9ckICHaMg0zf6h1XAANP9dKUflHrP5owa1BdL1L4QhFqZzFB/VA
aq68GIex0ZDd2Zg5xLUNzibIzDztyNJCHEjNceRATbD+UKkzav1CJxXY0qC0BB5f
Ms9qjNX2128BXcI7my0IcRec0+d2URX8Q7TD6siwdQAaSHGEgWcRgFxQxaLvDtGw
NujIIiiw922+obPCAFVGNRn91kpDQyHrFf8wojE7EBaKlLAcekGH4XfVwvZiyGvU
8DHKpyqMloW+QfALAbNROulJLUlhMIpW6bmCDxXr1mycp3qQmFqMsz3KXVjg9Vz/
wB9R6h1GnT3aX6s7+3G4RJ1PM1YBEKSxGebp1MqKKaxVu8GMrPXEA9W+KV5Enp7n
9dY68aTm/y2TCDo09LVFLNLqM1BoQEKMoyMLc2xPyWnVarClWthdzrw7gknsY77f
jvU9LHlixtVGKj0OBw/fICiHHK0oAFySaGut66GFBV9T7fItpdtidWogyqcEVrs9
4tzKq//9+4zxl6d3QVMUWsWLumiIKwIiZ+d0ZQM2LtovDbkprKAVcVuYkFpGmdnS
R9hTaW1g5Qr5VUOPWkiw6dEmzC+BKH7uLbUoa1c5jakJr5pXwZHTdA7oQZ97tCRM
73ZZr7UAC02PCZ4WJiR15a7tqDcn+o4XEbrX3puMAa2o4kLgM1NQqslKHAyt0ANz
YE9njPMXFxusErwetGIE9nLN+KinoYnyOUZoJFkV2U9OSzdqF9WG0iaRShOvEjCT
tymG3ZrmacMW60jkV1/nHjh1hVpY0XQjbvKsackrzL5jA9nT4ULiwiVXAFcl7O8D
mIjRQtNfjmZpt3mbngBPtCCopC6exJdObO8ia/9C5OrbzzC5V5GyITsILZLYC5Ao
9GUwl3QKvlGsjVgoTnGyWVVMfOt32M4N8SAEvJu0tol8XmRqmUAUvuMDZncjOUT0
WwZPj2e74epVWUSC1DRry3R7IJUzWFlgyvDHErhezjdtWR5JaWRwaOqhhBCXMNEb
8v3c237dv/rCY2r8+YD5aobfAEfzb5S9CsN/bgKfsnL0darbFz2T8mltzok7Mntv
tTJU69zAQjuojmTK7sTLI7C0HNLvPf0Q0jN11cgq+DZgxLgDKb1EdZ5464oZ3bsL
JS+xjrcC5wfQiYbZpl+TGtAlaABngeACYl8izAH5Gju8g1GOqObEH69JEhPGj56L
XqAL4dl1X5wC+zvq5JKBqHV1nOHS0CUp47rhuh6U7qgsblw/DqiuJKSvuMwtVNBK
nuzSS8N1XFGwl2UJBIDoW1KO881iU9Q3vG0ktusfp9kIsc1DikljErv5V/fscofG
YAWBIiC5e6dhgisDjAMfhy6tji1U2xihSjAG5uz8Q5HTfzLi8hyMrwJaJTT6hoHN
jX0SZVB7UKJA8RpZt48cDMePiLPLr8OYeSBPQv1el+8hJF5qB6GkWAfoW6a2IgJ6
hPBu6csV+DzWPpjEDxR/B2YXoBL5QQ2mYwY/h9GGSQd0oUmsjFt5MLPvGkjJHLPB
HiZyYoS0/KnJqLxKHh8BxbgEjTG+fQ+g9sMXcxlmH9k03uNjv7zjPrk6mI5sQmVw
+RtuZu+P62HrZYRT2ldHhNprGOULH6478xYK393fzVumVH6vT46S29K6muXz6v1C
SppWxJaFDA55WtlyComc9gwaJCD7QtfYl8KFhEs/z77Zw+yLBxMV7b0ZsmZbIAT5
Xm3kgmoPeG9vkTsei3bsuSuyUZBBZSqPWTlzjCGamWZBtCyzHSCWjynhEr9FysRz
S7liqlQBCpCVJDiXmDzZ7fWCS4tHLEqGGm4nS+CTJNcE8xMI/OlipxTSWC+b54ZU
YR4tTuVj5qOG4M03Y7NPXCAdIAwMx1MHpo/8C00yawth4s3y6XlosFnSxD04n+tg
fDtbKfBWCgFPfe07b3LFMq3r6pRrd7zWqjjlfn31X9y2lXWOtukXIwIrtrxojqt1
vz1tEC6XhnzL12AUvFGtLF+CuVKDF6INwPHQnk1gFlWTnuzp/yvZ5KJej2Mn0KOK
JIafX7ZKatrU/mS5CLbYfqLKVVt1vR5Qv2tUY/tnFSA4Env5izRISKMVKvfugRZH
NAzj+WonP/Evxy77AetwsIx2zZQHdfvuyEIg9QcJY5zhah0NiIgAlBP3FoTo8vla
CAvy3f167AAaFZSvt8SmyCE1aRoUeRUl7YqbW4eBg4qBPienkqpbz9172KbJeLu8
zAI23tf8fqdklgySO2OozINYUHK5AMHDN4yDjEW+1APL/N3eoUY6Xb2GJi16VHG8
NTIHxidnciAT4meUsodq+45AR3QIuADMMuliGJS1N9J8dx55fXFusf9azV47fS0D
+1cHmMbCv7HVIL2FE0fjdP8CNuyhs6+smH+4LuVAeF1PuUYR4TyWB7MykUZIYbEA
0LWSgUHewnTT/O2CIKZvx5OlE/fxfSCo4Ix77HTvhYR/hf90XeAlIVm1IrfKAJJd
PzGJr/LmYJyTlF8LrfIwzmLChlwvkYbKmHXinToY+Rq+t8yFG3QEfWdpyAoQ6mqm
bZ6w6b7JP6haWhqlyQ8KhXgNYy/A3h1TiMNrYdy0bU8WWR7z3C6datvq8mwpcA9W
rzVwJv664i6NkAAezrJOZweZP0i9DddIaayUCJZ5zIZXnttVI2akg4EZL16Xg1Dl
lCxNY9hf3LQo9DacRu51wpJOfCrGIUEf/me2smmAnwRRQ9+HwolguuJUgeVRROQA
FTGtecO0BHjLoQ2+e5YtSthm4kUj4LFXrIAGXhdbA6maCmiZseKOCfeaT6EyAJqR
0SoXCmGk9YJvjfmOQCdhVY2KyPvO7DCJ/+LzT/OJznPm+9ycPSpIk4YzPD3ZzkfD
YWVcaJ7z6WramsSk2QuHdZtl5kJFyx7RnH2mailbrEYCZDX8eqhy9iE42cyXLVAQ
T4nLEWvx+V+n7eh/1i/pbgefoAUEXyqqWHNtFy5TJDGq+stob/JqOCPTqx34d+LL
dhu3EhgGQBfuaQDfqNhXIlFU/Po/9dUWmLtdDqaZrUhe+bM5di0gYMMebDUlwTlI
5+iqJaOmZFn9dE7jC1hBjqW3zR5+mloTuGpulNIn24v7BRQztO0bt1kGVj0sVCBC
bQikcs/W5RK97sRnpjF6y1wUlHRwABLEK7EHOnNrssAGIDM1AKuTx8q2B2O01BPN
n47zUXEH/3hwTq/xozZJG1MOGAecDoSLY/mizo24U+jvYAhfbFqHQrkpPq0rul2K
t/nngf2EAUrlSBynvXqUQq4L62UhpR98mCHrptcnQGxiAccvz4QHH7QtI+HwpFwY
73FlYB/LKqQa39qY5TZjFnFKV43yH1Wtw3mbYFj3UJyXT3YeT+d4RqJIdyNY7Hgh
pbTYXQRwefr0dwyIsQKXXC2h9uIDE/KadFnev9KYD701JZOJL6RF87bltfK0wBVG
RKGIFsk9PWoIOa2OAn4ZjcUCfa1//bZCG5O+MVaCLM3dmK7BFEFFEZlH8WCRrQ45
Pebph9pLhmMtRY4HerVPKHqADAjhd8K8oRNCwtXzk/icDyn3NElHT3F2PuF9xxV8
G8HMxL0+/QZV5DrY+G07SiXfZ0FeofW7ar3KflwPB//sK2B2rftCQSHT9SMUHSYn
IgHreM4aVUFY2bSONNz5jMsrGMOW6erw7hasOXlUZnk7XtoyqxAkLKArb1sTjC/P
K4HQ7M2drGjdjQ4YLbhfacn1upUBRUWFx4YbU7snKXTs7KwMlQfk6lPtLNTwbCcP
5X7LDRIAEV3OGKge/m87cMOi9KTLKCFrYo0ToZN55ORy0EqM5HuERMS0RKlMr6u5
q9fk9YnmIQBPSNtrQr+xxzvj/1ePO3cQNYM/fXZy0N08nDdW11tFABc/gVroCiZc
u90oYA9TPRETZtBG5zHAkkG6+Y4fxLXT6qXWjGiMFOVXlzvv8DgbFkNpuP9zmbED
m6qU/pplpbntz+T0CssBFcQyKNf5zEOTA9xjBbqpMaHmAemRR/xjdJVM3wUrrVYG
7RQzqmqAN3zKzXbAOnFzkSRIO4Yw55Xeyo7bARuzEufI3jTsylOoykwUpxWnhLJK
BA7tJPgiGWrBVRUtiOTeuVo29mGmkba2VaTWU8hwVXzfn/Jx080r4OfxFI7VYa3I
wqCX9Fc5rrQ5m8q9zDX29GG3ytIk4ILf3rvCNt2JAuOWKc/YNRpRhJQhP3yegun0
WJtMXcCVDVGcbm9TIdV8yMWsoEbM4n3nwKjBuW+3ellycDgXoNiYsm4H2byzd495
1go8zzX9RSZcUSpvIDHA5o4T/iLdeDkDxwiRA7cAoO83KGw6Ut939PK11riCUwr3
38sSNLc8qRC81MWU4dhfqu3uYbABdyh9j3HQqfX7nAaNAHeRXEhQFyaDFuI2LLWD
2lcfzdLAOsKoemSpiKJZ/hE96VM9TicEIWLz7ktnGk8qt1k8vwNBBcNG4hW61Ie+
Z9Z2rwo93qqXShzBeyF/fnkQJfcaKWui/m66Exw1TnzTvlUzPrdrNjb9PAiy9fe+
/2fLYx5TXlytasPtK0pb8F4Y+Ws5OSFXWyKVrd04bqTyoTfZkkJLcSguyoiic1ug
x2ZFtTzz/ZMaGvoecCGAQ1P/TIjp6LYkaH1b3PiyEM0iIlNOa+96Rznu3yFIDsCb
KLvwzy9QBR98hpUpP0czd8YNJarUSN1lOjNAcPHkokHMTu6hEBo7nq7AcO8D6jpK
0U7KX5b6XmwqOXZydm/kmbEDOo3epiHCC7zqN3pYVqacaVWDBShCxMo+eIlhO4ch
53bDyXR7sgeAwiZVktUl9SH3e6c64IonZRTzz1++nSOJD2EBAlYzicYU3NrkgWEo
3j01l5qJ5vYbRvH+VjqUOR+Smwt0V6VvGvgA9SkUjUjMbzY5wmkFLjBVo8N0u5y+
mFYMkmBT3/kVT6Ce4mQCDUb2UzFuoMFw0OBkfWUeMf0DN28zS92NfPt7JwknlzLp
J3P0BI4kcADzGnRBuXTv6jMiC+JU4BWIjKhmSWOkJGijUnxReWxhtaFCLFe97hrm
io9kvHZmmVkZTIN4IORnWCynMYYwa2DX/Tb+Mp5cdV54vBwoE+d/ytOExCRAiBE9
vcGMKeMQsA5B48MNrXxAS0XtghEGXf3iJTd5If2ytFDwcCpiGmUMHHzM3Y4pzLHr
KRx7zotvwc3UovYUjSY3lSAZcqZL7W9xRJMBOA0eqrQt2UuppdKS04TDiDkgtXQz
bbEuSH0p/yr7+VY0nJixh1FxfI+gVI97RIQcx43aTLmHaJCQKABMwIasA3WNtoMJ
8dOeNaqlOHH5YhedjGDtyxYBwumEH6yxq4iScp64LfTn9kozRMiOFlSOP8Tp4ZMC
FyE58nx81o8f4PxiJQXVTcNbFQxyqAJnNZn1tumbSZyIfLCbQnCZGNga7SSWS5aj
VJiBSHRJh6ZCEJg74LpY9vtzdIN/ZcKBLufscgCICUEO5eCMEpIabRkMoZu4ET98
6Ayu5SYZxpQhwz6plHEwmaUg+/CR7Q48hGeoeoPUSBURvRJx8lszIM+2F6ohp8x6
TuoSjdr7ywOA6LB/ptxRknzp3uiWyU/Rx6DI2S63lzjrbhFb2YetqvJqGY9PRzRU
s2fPPKcogXKpk+n0TBI019vx/dQYtuBUr0IJ5SQkkv3MMZPakGMo2vZNRLK6ToLG
2SwINhUdUFvrotZ22ypLzhEFaz5QkUKR4yKo1g2Rts4kBNd+q+VJZqu+6CGXzmyB
p5bahyzZlfcFA2PqJ/Qjwx1kzeKrD9fbBAnZpDc99K82qU2a95AvYQYRNmp4ALQp
Pp4mI87+7fHupZa44rQtaUivGG+PJ+Nu0B2+pRs6HSNS0g6Z0rfk5r+QIQSvOPtH
dg3MiffTNSSnvpmhB3KjI2sV6RPHjyFHtksD0wYNcjEURYste0PpPbGU7OxGgXOp
lFRuW3tall2AcsaXkrtsrjG1qil7g9AkjvVDgoXiMahCWzycyPpaeb1fwyZCGdQM
E5dGmHeIgJ4oaWQB+W3+xRVQN6juXFuLbjeZgspzA6gvNYlbmPDs3y0TiAYRseiX
ew88FKUosRLuVdXMExeQVzgdYB/UW++68SG8DXicSiz3MJGVVyE9W8ZQ3/4ndISn
yjeNTrVv/p1czCVEhYm1a1NNL2UPDMTmOUopMhHNOdvAdg7wt9RU+LN3fnuz4iiy
Quhpo83cOjasovCKOYMra5mCmMpVXuSq1/L/ai6/No80rOae93rknH1KP+gxa5Ln
qV2dTvCGwkagYmD4cIM/kBOOx/5ZdpotgRp6T9zpmWqsDcJD/gDsluvKrj4YiRqT
Mi7ophLOJQHYYfbpUk9f01F3/S5/ku0RoilIbje/SKdCI8d2zKBCxOCFBeAovbX2
aWvpyk8GhAqwSlt9iC0Q/6J+1OV1vYcVyMxfx/ixMNd5nXe8HUGwNT5y+vKUos2n
UQFg+X1oz/hvVcy5TFJFzg6d0fUjv17/BT53pQYVuS2bynHvDVz4E4qG6FOE3nCX
hrVt88nAZi5xdU9TEwvmOs1mTLjkcq84GO9raWIfATQuHWmiAe3FtQHx4OHln0xE
JkpcpM0/M2PvUWlFAC+t/Yl9iOc4sO8NyTjyj15Q+faDQ+vsHe71uxesauPs+J7u
v9aF/X6/iElDNQcN/yw20aGzvDJRmyKOfIAhB6muuhS/h9A4u5dBxxm1RmjAb3YQ
7ajjCtb5VgZQQH8fd3vH6glGoe1GAhtyKEfZU+FTqclV3iZ+AyTe4RCc0HIvyJvt
dkJHbxUEN+al9m+A6GBU20HFJJj38zHimlfMezfJNGtMyiKQUPQbzsyQ4HLwRgNj
IN2pjGp3mg0W6ENsHSOfMv6oGjYgFqlv2xN3PUX98D31IyCYdeixBZEPScvLcSyp
xXxO+BGGitINR7/crI22+CWfO51ahA2rdcLeQYuOdfbsMLu28AomJ2ZjTiMXffYB
IKdIdpWGZDfJM0dQETeU98jHj/KcxIkgffhWIfoCaN0mkVzYrRbNgc+YP1U5V+la
bciDTbzeHE8//4PO+Zys8z2tF6jJ7lyJ2XSKbYk8RBivu3h5ms2c8bhTot4t4Icm
Rm5Fl3olwHvavnRM8G4UC6pEjIilWkVRzs+3f6BPEaOZDlzfQVDwiIpm+jJiJm/p
6iWPD8r5L18ipqSDM4CmV0n5Xbtk/faGoLoTtjr/TnhCCLvNpuOKzxtXR0Zo65vQ
/pytVTRWTxSBabtoq+5lTMJktVyLIBpwqUEG1UKwfE0wC5uc4iLKusptdk0nci2i
+CfRoXnOaWQxH+OdMQZPRR4xVkL6d7aL/ZqayQvRQ84NfPx/e+zRUEEz8/xiR2m5
FMq8Sc7MY3FBF9viaUpGS2/s5guicY0b11Ra3dR7txNvuISJN0+I25UWlyc2r2x5
4ZrOXJG4+P21OQi9BLt2iX4C/TRwZ//rz3kDAfDP0W3JO1xM92qAMRjJKHlMWh9F
txUOiUxtVppxlvv1nSllVYSHJ/6vm0kIV1Yeztmvnuhv4eatcgDgU2FWiSdFv7vF
kUrvCfCSfsGv2bRCl45oUYRQ+LI+4Bevh0hqhCr7K7KBMkEdsIHGDSdqAlf7FXCh
YlNjneF0ImikMkOWkpzSs2ysF4p+ySR2hr+++pdVQSBN0+WCJ53ygHIFe4Uox6jC
kK6Y87phfpDaWDKSCCj+ga+SfZFSQRQuLCg6F4LNmtGKEkaONEvIHpusePnbW/jU
/EOgSjiW2EpD7EihDHWGPBXz130RMlcQ3zW9XNfmpyk1gb/aSMCL0mM5HwhEQYqK
6IG9vI5S5jW4Q0gKRO5CzUuEasYku75Y9uBE5AwOtlNRoelvviXXF1W8xLflXagp
yoNTqMwAHeVRI0U48+i72htek5HnRLRyHZQumvHjRpITFeZPFWwUbDwfHkJRJR22
Mm8W9TKg3wwjdGS5WKeo0ujLke1T5ToXaa4F2ic1GT5YzKMxYI1Jt0NA74XpYF2E
3vIbMuCo7HpYw7IatfVj0T9HXbQOugcuU5gOB4/8MZ8azj0EOvswwGrAAyNwjvk2
WjO2LMMYZigzG2Zz6nXJDGRosrZQGeT3ClhjU6e7gT35VmLvNK2KnH0yKRs1q+CB
Y6oI/Zlaw9J0QGl8y/etECqBXkk8wKx+sq0Dw+kvGGA8wX4ohBY3X+Np07fS13Wu
Xal9eBFGxg1XKbli43Tb9+KyImXiD/se94grjwHWuvxqU6rS6siZh19i+dcOIe9a
Pkuci50RysYy6IRzOOadYvwgwpIsrr8g8c9ONfWo1SnO5oDeFfB81kjnh4sBK0/x
zpYOFcKSIwLB5Hv7uj/Qsih1RRTsUVXMxccWCPz0Rma2fr2twjQilyqvi4gILfPJ
F6q7j6htBhh8NlEOY5g1IddCGGvH11bLNClJQWRgtshzPdYVkmod6kwBrLoOl3EC
+iB26EuMwmjgPMjfHbY1yYUoaJ2/BN37604VabTVKaB/CNNcX9+laRkq8bNnwJtr
8E5V07HKyBwaf14GQKRteG+ZxUpijJFFue9xaG8ro79Ovi0/ZDG6reiCkR8XO4Xd
LIGirSSjmGbD3zFXlBem5wn8Zxv3YxN0Xoh0Nt9G0sUhrB9PV+Cbza/xtewYAiAV
HU5iibPMdq5c3UmoTx7fktHKojZ9Q4pkU+T5xLj/Oij91U1KNWp6/D1m83uMR/0N
nDrzNp0RmCsYgueEwcveVL7+bzXUcCJ8R6b+wC4TtyeUqADu+4fpwZI9HCz3a2DC
YcZbqEN3GA9Yod9EPPsQOkSSGZhuEs0xhDZY1oRlmHPl1D8MUraFIazE9K6hOhxQ
jijkijGb8AHi0EfcCRY+KEC4htkH9hGG4rfchYfViUWO+XIZo1YsG97F+0yv9wHm
tRq6Lxjqbcz2MhcFuT+m5ksf5BDLIvOOkbJuGaYcQMXOn9Z3xwc0OYs+yGXkl+rf
zEcfwcDLd6AOLcIPe2vLvt0uHMeGSE597Y+E+XoOcyEuBr8b4iJXMm7AXN9VL0LK
sIs2+eUcbjNCGUns67rdJC8TtjxuDCmzxkTBG/7r5LBLIGT4k4CtPPweriqF5fbw
Ix8u+EXqqEDhUi871yxughGG7XcBNCEkH7y5RcWaKnAQzTpq+og/On2gArYB9VY0
py41ZDTFhLaBpNm7abCYmdjxI3SeY8pk03gMbA3F8uQDqLDCy/8s8FbDVbHGWbYO
v6WgPyV8kEhBPgnXZu8rmReyyxSG9Ku7cOTyp5TSh+kNKcR7GCPbN6VQGwf0XEVb
FMObnv4ZpaoLNPZAI8PqCl5HJbqN+WZRirgfy3UEWOePnwr9Nua6/OOlKb8AuqYc
ton2dzrA1W6+X3fk4DEyjvM7EHKOb6w6Nau/QfnmP1wtkEXnGT4eb2fnL126gV+P
kElmfCdDcktbFNJilVUEsoCc8WppQAhAJgaqTckLn/Re/O0QSFpIe8WS1KCLJ4i7
iJEtpeEMbHUX5jISHgmAr76aRZUFucMCG8C+VL9Eg4LGhk8fESBraeo9sFb9eiw0
DBS94yaeRmltTyofNAfttQuO9f+/jQSpx/i4+fqfYW60bVOQzpBLy0Z82AUWsA+E
H85C2fNkrFsOoFpiwuEepDpUnSh6uYuh+goddAyr3stnpRCKGpN+hDKMwIGlZBs2
F6nwAjntgBy5ZQ8c76snqN4mfU8Cm00aij5FN8wd/0C+YpLOgwW0kZoODPUrsYAD
z96H9u9qDnzxFhuIkNPRMbXo8DnwbfFo9G6IVgPK6mPrPwvzAm4cNkIig/4vchMq
zbe5tefHwVETbvMoZFhZfgFSPPz2h1PoF1pkOMwjGd/+iaP5hkmDJuq/95qSdeRi
6sqzSPVn+ltAcaGhtjKPxjnTSAUDJ4LTZqq93w2kEPsht9liJI17PXzui30mAm/t
hvsJEgr3gkS18DVOY8Fuj0jdRmiyWxyyzTimId17arofQSrQuEpspcbTlOktql0m
SYdZqwwtfZYT3oWtiCkoCZ1nst9N/VTcNY+ytknum97ytdID30/nWkMCrkK468xI
56v+HSHak6xoiDot1Jq4esOAMwsqlc8jUUzKIJ7CEApxqWEjDv1pyIF2Gctoxid9
nHyPBa4/Bnu7VL5Gs6XNnL9EVxOOS+QUQwVHNlopvDtWvE5BEhINz79BFKIY6pLc
qURRgF0ZyEnUdvoIHLq7V6vvkH3KUqkOjQgoAogM5K/aNVio5sRf9q0GGcGfXTEs
JYQ+c3ZITyUkcHqae7zI0gNtETaUWhOd9IA/MbpfXmsMIXB8897U5PWoRk14Em/N
fvJf6TX8R4PBjfiPO6XKK5lJkd7HngAEVZBv0Evhzfajz7rv/BQN9+beCQsDtdU9
zvkL4SLH59lHczITnjI5LV8Bh5/ePx+ex0X7eRy7xL4Y6DYkYhBuPnAGiow1U+X6
JkdjCicQAIKRDKyNs9sV0x569vLU9J7tOjUckmiAubwyRId6vNsDjVPaZxQ/NE+c
txJv7iXE0ooFw7w2vtjEY2aD+Lf6KrTAsW0aFrlvfmv6fe6B6lIi7zBkWFFSZVbB
I3qKWr8iBdmmF/yCHkuZXJB2g0SBLTCbBMKnpO76vAp5Wy09r9cUo/Cf/KTI8EBe
6+XKXl8X1pCA296xjWAaEcR9V3/wTISlK0cdsHHd0fJsUolgI9B5ULugrjSnBxrH
Es7fqF9usXDtA0qODulYB8Mx/7S19+cO1M4mBgCdS0n96+E0wwGtqqlEvGBfbg2l
T9mFgFRxGry57pLSFLfZikHFR6k5lRSJVmIjlN3tlF2vov2rnM/R4qs2UFAsNPj8
SYr51Nq9XxXsxlgm1/LHCTEyqAe8Ps+YIBf7k+/FK5IHPmb6/COPaYQ6nEssCow3
khTm20367eJ7jNCbV5cY/Ooe9tiGBGFXtQFJfBJ2PrPjDsF3GAFxlyS4uzIQs3nU
s+QLqC/s3qcmWeKA3OXdyVhUKg0lTwTZtoLqr1oPhTqrRixOuDSu1Bo264Wkj41z
GBNv2WZeabBe8WajKiYzEPXnEUP/lSmjV+oprXHFaQrTQ7fz9XkY/1Poxy4w0mTq
iAxOyzRISaOKid1RrfSkqUauXvrufydfzTf4Z7QaDhrA7IFX9FDCrPY5gboknE1I
No2b0XyZ+aQP5kB9Wu2Yzg7W1qywcemL7rZqElEnhoKIbIkt6N1JvS55V6jv+3m3
FpQddUjXuAkpeMVBoVoxlgOj9iVtjGjkpwVLlTDRIvQQ2FCXNdQFeqCBYMogNdG7
5S1kEZc+3VHGBMyh6PDXGoI1peNqxn2oi0ngnqFVovk35NM1L6neyl6A8EyUza4T
8GSOOs7ChnzyCHb15uxdUq9q+6gAudkJs94I2nJiFcqEQBf4HQxMSJfaFDjS05Op
dcQPYfqU5pTdFUdUCvBRecvpiMzUlcY9DTPmFzlKsne6u5SSmZboScnHw9nIpM8P
wj8r23t3CELPF41qEYeVOvPquTqLX/+tLZFgZopYZ2hG84XP/NXWdMVmyXKKb4xd
BKG2Pq41fz7KskNXcn2qXI90d8kqsRgc0Gn+1ZZLfZdHbtI6th8H6Vu9biBRBA7f
llb/kGS3MEy8hTSNWtVc/eUFcusf1mdjKPHL23rYzip5yB4n5UJj3Weg0Kp8HSzA
rzTdri92JDsG/FQcNV8Y8nOU8Ji8TTOnoYVCJb+LMRo5eSLmUuydPs1B3JCgzPiE
98RRvKCIrJ9Z5OuTKbB1SSoZJT9QjuewMnTFv/Pr+1Oqa0sGIUZ1QmbRf0Dn/ruU
vvpMKre/vpxsximMX+87K/bdLf0R4kUp76dyRnVo0uek7KFlxL6yWmI/VWqn2/5n
xgAbcn8dvEK0zt/Zb81+/Fkc6ayp8vI1JjsLyxfbq4Gqacr/mSi6VVge6UhdLGA2
JZ3fN5KEzcjfmBZDyYN9eCGe53iwIe9PWKD3rBuGedHTywuYAdy0dFGtKRq6pxf0
MCtzyzm4UaDNx0zrp9fpx6uZinzynnxrXBcZmvC6Ve1vCOgAhNdqhd8qRqCZ2MLz
4WTXpJ3Ios0W0PoLoIEYb/P/HB7KruRxhZDhodGlCrpndp7qgJflA/2M8GMMyzq7
BmM8FFPhh/kGbTu55EtWlB2HFEOZJRt4WEgO4kMi6dRQI1ghkqkFhMl/4+3HvUla
Rg1yXi35mTD4ohwO89oZwVKLyadGBbiEWdq9aCcqWjFEtOEIAfnOw8VkwOTKaQyK
qudXHfWurqtdziipoLNoCWV08g/Mff5TyI/mpBP2MfK+SC40I1keAEjkvL7rKTr6
D4WiD74pE1x4Mm5hxlRnETBR6guFpNGZ/F5F0UGeI65ImIHHBhM2u3na0wpQAMoF
WxkiECl7ft9oD5cP3NFRqI2Bg/nr8KcFYj2rcB9zSYn3cbX7jIxJ7NC3LufnWpwR
2ifRluyrvyECG9mEXHu+auJ1ff6jVec8TYdo8PL2xlg2FbnUmkrxqhUzIn+sqigE
i3KIzCyt7OuPhYCDNf5NagJFlvC+Q74+LWZyPw0w3dNinKbTApLHbHLUSItTEqEU
hat1GPiWAC56HBuQ7J7eiv/BsJhgPoLEAYh7O0ESSGAs/wEfyw+rWwPHHmrU4gP0
hh0YSLjSt7wBLbhKgavIT9EppJ4bIKV84VFdEyPKe454AsnIsX+PWax+IGs9mYCA
qLuFkQKIl3s0or6JMslBKfYjImgqLogEki0z+TgRi8RjJYnfUZc07BLS62+N+AY1
u513TyD5mJj25CcaJv94B6XnpqJXazNzzC6Vb3iXL4dcBb9esJm/MP2827f2XFnz
DDjoxL52dGzSFHd1yTJ5VOkzFywKmvJSmx+/Ag76V8klqXo3yfuRRZ+jpx24CSTc
QE/O0NdQOVl49FP/e7PpcoaBkXaY065ifar11Kew02uK9Y/qCHck4Cdz24y61Okd
fy5nMG55kG/si3P8hTp4OtmNbGFBAtZTUFNju8jgaZQuTkb4HSvzeRu4w06n+CWZ
p+kOEJT4/2w+6nfe5qr7FFlwm2dBSRQHsB1uiB99/kC8THFoG7szVphmUL8UsNpt
BA5UrSAApD1TTfa6rh4mmSabmzN3rPtjALZZSDqDNQVMl0IGZ7hKT6yGqh+8xFfZ
M/B3X8eIfzraibhrFShfZTf9M4MpEXHEbHH8nXD3FxUCtGbC6enHpFuANbG4Yneg
9m/QH3+80AKOwNwaZOYWBuFR/5CgerSWuVQerBf/PaC1P37VM9GYazQuBW49CUs7
gIJEsdj/cDd0aB+wGv201/K83iedSAYqCBY6/GcNuHdaSfsE/TqtCikWYBaNOGdP
/99bPp13kpUNeHjuJ3fFt089SPQEPmg85H9AJU9lMZJaI0dvOzFymsS09ylsGb0w
IOnAj6hcjUMaMjMKLa6IqrC38TyhNs1GxbvdFPcF+4tyAKZI4mYySOyVW2A58P0I
tJxAgtrn+JGQzdbwfqf9SSGS186s40Ch/329gy2D4+xu/RayBwwq0mUpck5qeOoB
xia1OifIx6kXYuvWDfuNX6PDnvOKxnJT8et6O15qumSvaJQYIRmAWj+Fd33o9ue9
xZcszgypHx0S2/RYQOEFiAH2PhASQ3K2+dHkHvhjztS/vUm3m5j4UPXnTDDFUY0V
jdH5uGNYKQbze8RdasL7G050g76ijJU+IM5leStDM8/9DptAvs3xXhf+URwE/n3W
PK3T5I40xTVZqkx/KBZilFiPbrLX9PKKCGVygkSkkqQDgoJBG+uxS+uRVqlCJ53h
4zE0nPfYIEdaMJSYAkgzMDC5F+mqfMldYsAsQRkkxATpixkTQvakB9EYSoG5nP2I
SfD0Bkt4u7XSZOzjKWfhlC3/cFi+XytBLYvbea8f8GHrCO08dzavZQsQW1H1+kaP
l0G36xefrgts9DR9isR+k4Y3eiQn4G0uwWl1d8BwFHtuv9Gybsnl807ZZu2+XSgI
bC8lc3s/kzdzWgDH020U6hzNwbQuGB3egUJa2g2rBO/t8/4RY5flHTMX/zceZWuA
SdZA6kV5y4Tv9mPULv41F4po+14BpvUnlcYjq0jx3TkhSxCh4LxgPIyEy8cTC2EE
ZLG028nKOF4ewqLshFsn3wB06L//Ut41rmSRV98Ud/66dxKVb1QaH7B6Iab495Ti
RopTMZlg909OWEYwlqNa/0sCbAXvIDKHrIb0igDCSgIIjG9xnUJk5Od/GLB6qsrq
fhV1WtvfUukhQUjI+FnjWyZ5SHf0b5B0e3IUVd5p14RQZOj5OxQVbLCN38Dp3GPC
Ty4b7pDLkrkm1hu9u24FjEmEAR47nXH6L0Sf/6rOui42bu6CL5jpnAr82ydeC3+U
RSXC3yhK/r2OxLF+dKtdy92rLTDuETxiu/LCAHihRHmr7EdCET6gGgLZhgMkPWkv
58joP0UjOFYccZvJHGLIEtQ7g8IjCKuQgRdg0AKV8Aeua3OtvMHTUg+NuTZcnt5o
sSuEQ70t3Rlg/2CEwiV7+cbJYB3vYifeGbycias5Vu71r5FrREImcPCWMn1z+GRg
CE/iuTUTFpEBX4BK9Smk/Dowkp9oVSMq77p2zowF02CR1oQ+D9fq7NwBS/jpCpRG
jVLijo+B6yoYxf2pJkgrMlZ0kwd9jxDl8C+Y9MZoyM/9rNI0Els0gr6874IgxxlY
ZkCiX/U1jGdvxeJ1AgSyPXTCT6NzpKPjD76wjjuGJo0hM4XkXqYC7Sx7cIJXCQhg
BR//vMI3U1pt9Sq8LOaXBDmjTuSCfLFrCAuT10taHwCwyso+YpW05a7jjuQS8fef
DWlq00bPmUCFY3leWNZGBH3pOTyhNnxU+ALUTpMmF5geHM7o4bfpUDmdR96A2W24
+hpwTufJc7kp0HgfMnYwoj24wRNo6IJuGW2yhGwbM3+WKsnAaJEJvLV1sBHcHGmN
a+GHs06fVgyQmjCAGLo8ioDZOTPFuH2JWGM+9fInYJVScn0Fg69i0V60A3BqJwxr
95RBJ3zLZNlNJz0D8CG7kRXj27wMkKGscmty5bL1z8iNJlY+D9J6WJRPBByVSm7S
QvA5IgbXKeOTvppN8tgmDLKVAK6ndSMjfmrT6c9r1sk8jQzZJrO727YuFI9ee2iq
BgT9VER9ytP7fvlE2DZrxAqbkP1a/ZQZpTHcgMXSLvbvzJU2GgkdlKUZO89ueWGa
aicL7aQnKvofdu2pKdDGvUpGLpeq//Vn7OFqJ4jSX0XcL8ZyNfzyBUSLp4vwJFGf
B4HGGXKpXoOCzVENg6Hu7Ms62bc/qml9VaZARIFM/Geb+b6tWLU0tjshcU5MB/Aq
ncGovqOgkAiGiHQ6pjkq+AhQQudEVl8Z7vGI0kZQ5pza0pg14zS0jXkMmz/eBiMt
LKNn/sOOBIJ2WMH6PZZIkX+OYwly/H1HCa0dczA2mItzsTwQqs5UshwFHMvIJVkn
hvQZL5MemDPbfiS/GxLOAt3+J+SqIfeYJdNfm9ThubCQNePR/peZhECcVFy+ONGu
tjqcfnD2WW7WJt7go7zjGLyWELdEAyyVFQovLOfPgAUFm1kvn+U2EL0PttRpZcy2
e5qW8srQPPq2iU00Io/rkA0S/z5T9dzoFhBT9Rhv+u+YtsZRlnxDIt7KvmigM8nO
BPbc4u+pjVgO1Wt+WBiY52EH6fj4O7N2u58/4RT7NcBYM9330e5wKPpgULekdtgN
XLhh0dyQzqtoGLN+apZ7OtQRSOAYbEfDXjGmEMqZ07+kCILmKxl72Ac48Cq0/+EY
hsBBYHCgn/A1YPdavUtXpWPQMSpIOwVI7T/voMRj0lrEnMhgJEKIoQ8PhCezLBmj
GzmZF3V/hY1yWhGgIHqpfmx5mXR5utPWcEwmfFv+82EMB1OXcxJBSRWxDquLRkLg
rrUMulbsDkNNnvm+e/29SX0z9BAVaRtR5uu9K4FkGGnn645Y1NMb/Ugy9Bne78LW
ROJ1FCFnU2wadc+d5Ikje1DSTsTPy84B3pdVt8jWmNXOUvawtqKQ7cdpPVqol0FS
a4wO/CIHOsnIM1HFR3eJBZd3bE1NSpD960CcTvEwkSW22k1yGiHfTuu/O6O4HQTo
yPtKfjRCIvx59GHPa72UT0TompszcJlbTVdO05k81fvihqsFHgR8MKLrudKKW7hj
Ep1HKq/m9p8728C9gY3KB5g5yXHbXlO/jJ9BqF+WXdNOrPjP8L9rprwg/lfpRTkU
FZQusvIopqhVOs4gqjpBmFrF2qLT2wdnHyNadoV7f3PXUSoUYc1vYhb2WUDgFKZh
7I0LbzMHVqUaYq6urOzcYrC+Vmq9IQr8CQk/FdApACtZHUHm2FIug8QeD4KWU9Xp
cF/KNAH59MKujSJVncAAHjjV3dEamcqSzK5NkdbOYKULOw9q/D/Maw4hoFdLe2ip
oGGt1Rx3hIu8CTuSRJlpmi+GQHl7Wxm8ft5AB3Eik3TSKIYrOHP2VrgA9flrJLPW
GFf6tu3nbrNEVA7EyJE/09LxUXrb7xdUWrP62eUI1wW/BvSPABFraCErWet0HzAH
X4AAppr0kEXbfusO7DsTQwXaWFnfapw0E7TXXCl04FkA9AquLI+wgdQJxsJXkPTA
wS7FAWOD9Lp+kwIaYZgM3tUKmycb/wBiYUHjtJrnmF+B2S1T1c8Mw2mo5Jyu/C2I
FB1196F3J7v4rnTwUWbcX7IzeYFX26k2SQCoRBwspjNzomkKKT/27VzRFOaQL/JK
zmdvBOH9O/6mQP3Kjcj4QlJuAzncXLBPryosFRapXL+hu20wsfMMc94LKKUQ7mh/
BLTgldRnFooX7IJ0dV/LxSnYOYio//my32vMvO/QOtbF4qjIutNWxZVYTwLIhosf
0VPkbJAX8yOp6zsXFsofQv1yd0oA8+yYXMhGgRAIyf67i1GibChRCsl4+YJjMqYN
DKKmbnwXVQ53R5SM+tXrKXhJsQFano9jDbQQZnDVrNlZMcU2eLVx9Epni791gyGg
qkX71K58WN1G49vkGifcEzGpQKycaKpnicoKs3uMgU4iYrTIW4hm+ygK6Acg0aQI
ke5RkGDJZXP0pX++oZ1q+qKU7MIr/udluvkquOdfMBQZGgK2I5R9GWD9uq87UKDS
QxX1g87GV5wwfJRqSwIqHf/tWxYMe5zmCpZGmzAMC6mN+HQwGgIUz8QDA+g6En4d
ex0XPBsP95kfT7ENlropSRc03pXl1q/7V+zLZtEAkV6X8Ns5org42htJSWGAlOmd
M8Uhws3KsLFKp3xbQgzAaSI2e/AfTORXdR0YYDiD3ZnZRH6PbPy3VEAWGiCTRqSf
uBWu6fiIWnOkVxni1f8aPGAwstyfI84kVPEgjp6nmuwHyssbIUCf8zUmbdLhu44C
oCF43TOxniz5khiQ4CkOpIwqBveRoKxgR1IYyjjzO1cUVmp5/V6rSQ54lpQLzpr2
SKSlfQLUgQhqXlZPGbOnqot6tAvBb8fl5onCl0YQp7d1cDSqrpKoWnvJ9w7UC4Bg
Dr7xtnDI6OXGIpGa5tSHbTaGnBhhfMJQyxMXR0ODNeKITP0NALv1nH7pabPgU0Ad
EqxeAiG9CfDsBlwIvOK0YAbF2F8jXq1Nn6fhzaEwoolYG9a8OgnTgS9LqWczeJ9S
SEAdhTlchJeyOjF5MBG1arrIBwmj63t1gDRzOPRnCJTAMc6OrQnm3bGkHhr8mH5B
PVMcrYt5PVYI8GK/3RCiFvZ/DxZpEWeaSwdeozMdqs2R9Zz5pZV3p6WXTpZ9FbR9
9QEdSbcdMfCubPcLViyWy1eewMq74cn5piuH60JRQ6VoYmusVJD/QAiJl2HN4SRk
DMM3ikNAaFd0OqNLikGsRO0Qd187aiKQK/jdHsFeTTWOH5LW16WTWQxPwD2JerOj
dw4ZQuMTn5GYgJQX5xgONdv+Szc1IhvyfSZA8lcFnsuXOb8y6VmWqBeKkoAX2sLU
9DU+N+WnUqxuuIX+Ddo6plf3e2v/1gP0cDpeCsTf0pcp681rcSj+a3lUn7EJNVwH
x0YJdA1tUxEUciETCKb9f9Nk/+8Ls2nDKZnR9OohC80Hlvti/hEKgPzSKW/6CQDf
51CDN18kgggH5dYZaLiRXA29ThxZVniyAWLj6QDIkPsI46BePbJRzILSEWMjnk3Y
4j2+6UedZIzaj6RhxjtVWuBPblQ1VI0U7PcOeXdzEkpMllKpf4HrpbWcxdTEsEVW
MKgyHnUXLcdGDhl7bOY78WZiAOjdzGD7wiSHV3WAfHlTQTcwSsfjTKm+htIuFXJj
v4kgdDJkm+XCPnGXyr5B87XCjHQq4H2QPEPSX8qTBrDuCXTup54dWKRm5Cn86EJC
fD+Y0/P8PZuQ3NCp/Qz9IGYP2ZKmXWAdk9BwTSmz32WKd4BjIvknI5/fkzZx/dDR
Gmq3K9YX1H5e30RT8MhclVRX00kzMh84GAdiebZgiWsaNBkMTvfi4+rvyMHjaoBD
b5lduGHuTKricj7YN/cXiVuWgp8ohUIiwY4KD7dax/dOad6LdL+KS/L2E3C5j5an
bJa53NXgW4zmuKNUYgV4oSdwZQT/+o4v2XZesAdL32QQc60Ey+sbkUxBP3F9LkB3
kZPOcsJsAn8Pq6bUzUptLngkvqw8ZfqynQDyNoumUlGhsffeibklQff5TY4uIcBV
O7VcSWKrJy+CEzx+kaSiPnJYoORqZ1tOdJdPPr8xEhPqh4CQOz+Lc8CQ5pekH1Pd
B6oDoQF0r5/WiyuxY1yHfzvuJqXHJ1r1egWJCdoCk8okxBKRMXJKI9lpkyzXnsV3
RY3pcZbOpK0n4nCBO8ZLeFj/u9XpllF9jtiIhzf/mi0XxDhcXtt5duU5wpV5woM6
GwIH8daBR5ypPKiMkEY0kkbKJUkMLN0F96Ki11dVDEQkt3QGqaoKnY2JZCGI+lX4
UrBgTkYFxuVaKVz2I1nQT0TWU9kHFYP0GggefWkz5K0SY6xXXwRQfS0j9Ky4WIru
ZlbW2ct8GQWxOUI8zkZUOTZ41rTFBCh2le0w1J7z/bAHRldtDkkPhe9ObU+XfiFS
D1HWYnHl0k1ScHbaR2ipkjWO2E3BUuPgOOoLmY27Gdfr4HBz37ydKtW0f3wH+naT
E3shMAyPhtQQNpYJ4J0CJhdDSJfxce/QOyjpbGINQ7vlIkFh07upHP6cJ5d12XG5
hCAmKTU2LClIMObE6ipjE7BSVOsBf4apt//yQ+tEBcwsmQhRq8EO5G0G+6cN7IT8
ZojtXyyZjU0yJluBZgN14MRR4pCc5uuO9eMVHMoW6kTgwWGuO8aEJ+WTU6/Sk/B6
Jlu+Vu+yKLP6uBr6kraawGskxbOst56iq6z+T7u8Jf7rMyEPBfDrpRUT8CIDH+RD
EPMaYlIw8uiYM/dQcGlFm+SuDv/zOgLAUl3vKpFeWnIGOKqC+vQArE5uKFxaPq0O
qxZIgCta17CJer+Sjo0V4rZfWAjvl/VDxXgSsF6JKY8ays+3z513RyiHJYGtp4R0
4T5gz19JCPIKrNlx8SUBpYGSQOPlRiwezF7vXEOToSdEm6e0BTt3rL89FC7uIJAO
OLTn/48Zp0sslsTt8Sg+goqf3LvRVfkLwrhH6qDWrVdnwUGXppy5pu27MSQ52bEw
4Jnz1ziFPldjRxHDBlCVXwwfQ5T4P/zjqbiRq43tHZinctx2sEGE/uNwVBNFa9c+
bdhr1xxcx8hIj4NGdSO0e19GELnwVhvVpVlJzsqVLof7dxSkcluP+10S7DBGLmtn
QKC6WQX4vueMoYxj1XXd0o9IyfT0AyPbcpaIrQMvISNg0bcuygoJQYeG08lFekwk
caSV6lx2xtY44A/04CkOWaOFT/pBtw66FUDiTz+50eXqz5OOyv3E1ksdZViknfi8
MNZS31TVJAll9CaldYgnwZ2l5xqBkNbX0lJOOBLDFv0jhB3fGLq00EW8KI2MQZYn
+s1uIfEtzpAb6/QPRQ43R+r96jiDsXvHSxL1uuuGGyHXxvJ2L2NnhwO90DfAJY8y
UuU/A3BTSVmVBf52e5qz0Pe4V2o+EX0XlWt9lb3UNu/ohOUKuFzx0DjaeeY0AIbL
OfCD0wtlhyWI6ErjhGQSGIyxglU8g5785DFuDQfXYkPqyQF5iTXoc5iT/1WiGZVc
lTmHXobMh58SAO3ms+ramJ+NqH+doxj8DAM1Bnq1DRu3m71EngWrNQ2URtVqOG7R
kMQ8WbwejiR1aIB/0uZjHg+GN9S1dOvPdwKjmaXMVZFVAyohNX0UapKHp/t8M7/h
0KQKEu3MFnM/kgGeJJnb/plAs787RvxO/yUEVHyKZMdgIKZ8qDQXD7+VSoVfH8xg
htS6XR21p9f2NO0dokxQqU19vHAhL9rhLBHzIinH1JMEUYqYAmo83ON8o6mUzslT
T5dLgbdAlCJx5sUL8X1eXfHDvimL6fEj2gNtCEYU0CY12yWlykRSbAed1tIKT1YD
y63sQttVqy3o1UN0W8cHQpd4HdaBhMVe5hIqcorl6DUYaoEFlZK9YmyxCKBOi138
rYZ1bVUYzcXg2Lt7WMDlSy/Ll8yZAiThpxR9YL/4gMG+i/GP9yhA+lJV5ol/SfaW
+nMJXPh+h/w3M9BXgGnvLfZzaQGBSDmpD8siqDd7sP62c9efubzwgrrt7r/Zmv8l
F66VKGp/W/g4MjDGkm3xS/XJE7rfjCrZM+FdPb9SP/vISllezPcZF8bEvKeFa6UX
IPmIRyab7+oCohLCXksSdp02twGMzvyoLYRxr9PE1gsCGMQPRLlybdPqLUjYzwDe
hRlaRByjQW61haG2jcBwNXOL9xiqaSSi3YKzE0XojXKHBjLpr0oOTbjoR1eERwWI
sJZBlNnV3nwGuEPZZlXpz4LDiIXxMoyneuhedhcsjQ5QbfFmqmA1X7Nl4q4I2S1Y
ROiPFABEZK20KPOOuiL+3dpu4Wu7FefzUVW4VWiSZh7tMLr6IvLKxbthhcCLUlEL
J28O/uU+43s/yhZReLV/PPGi1GxyIHmsPMvSLWjHrBHUVeod0VoW8rQ1HHt5Drrd
Uk1rHBtDkNM7WdKYWsvTpm57wCXalGOZXUbqvvwT1gd504cIMtkGes1Lc3FMEwyS
tk1brfbyiIM28kt6lvMGB+AW7xlTftN+i+AFEhniPl34EaCXP62Cx4TQkjgo6FQU
jA7wrZnzbJRHN7kM+XMONQe9tPTWrUl93BQE06rOKDCi50lXyU+12BMfeX736Dx9
ihPaxEDn8kH+LRSrUU7+18Phgje+2v0CDPK2JN6uKNzkpSdUlH/gCWDQc8SDbVbn
rXUB55MFOEAMxmt9Qr2V9iyJAiNdshLbn6lA0+wjFSyNMP+utUecjBhr34eeL326
8ZMCLEyAbfxpG1Z8bkIHwPy40api7HodF+dc68jw1mdBaHrib91YMalBQ1p2qqZX
TFLtnthPWuiHaTDJND00ybtfs2WMCxkRz2ijZowtoFuFBsZ6C7AjT4wS+ZMMvox5
WUKWWToaVkXZsA3qnFG9YQA9YYQJQjsTvF0fSQFX43q0Aw2tbbeUdKVoiYKQ4v/h
EE/xMpjk6HO0pH+5bB/Oq00izlQEvMf/BwMvSnxd2kcz0s1aNpnNcRYop1KrbXml
QA0ktTODrn45fZ6Dk23AI+4EuDL4n3GJLXGCL35nB2R7X/NWjb3MXDwwuDjSZsP2
z/DYI62chr6C/6B/8lyIjKpkkWtTbFOo/ysyFazpREGnyZuMtNZCiOBvEM0cPqCx
xZjNCHCztRKxcfN0OTlCFJivorr64F6Lo28pOQ4GuQD+geIiUt3aag3KeEhAskqy
ppdRT2HeyMrpkdPmdEgsy+BVBz+y7f8vNTqtOpaTb2V5Q0am5xebhxRRS7PFjcau
abLPyeJD5t8fcEF3VYyv999u64RxI1jPlHKAt/ZFRnGv/MK9F8dWGQ9lNOMIhnyv
E9wkZ8E0R7r0vUzRWMo3ZXLVf++gqDV7jVIu42EqCodwqkqeNWwIciN3inplUmRx
D+m0WsYB3nWUoBqGCaBn0Xybzl1brXfhveQ3gVBTrNhK2iOE9Go0tl7WVI86j1F2
+dswUEkPkZ5RRLR5AVF9ztk8z8Awg9zZr4EXdaNmKdYd8HvCqZ5dq5Jn0d4U18Z5
ObHBGyLjpN1d83X+twQ2QPKkqXwg8sYrbPq6r/gfzGPyeAVw9TGHunzlCxDhNRSH
e671QyHzvRV1V64cSYRyAEv7nf6L8MxoQLyxM5ZDH8BHYtHG0Q67BctI6BJ4h0ZN
QjGskD0qz0XEtLINEpfg+Ch1JknunQeoa42DHwfAXHeIJEn+fNQbIv3B7H4JaPOr
Clh0YDZqDmnDmtmclFLi8gXBl9SmwPndhGZZIA8dXgUge6xmzvAHufXPc+o+F/ZV
bJHaqA4pS3iZ+v90ISIjxOyVJpyxX935Twc5zVm+jksxENa7jFyV9ANfRzUwB4RM
Q982mw7WoYldPc4NhKUs5hcjcMe7gkrvSL7OOP90yr2wp0g/CdrM9U9rzDaeES7K
vlgZPN7RLdIpnTAVf6rIkavuq6T5LydDy8k/uwr0lYcs43DRvkTUd9mSqCSVQdMo
MxbgHO/gvgCZhj8IEUfaY8gDAsyFZ+XbJfZYIY04PjyjQKHdhd9/DRn6HA0eRo5Y
uO1q5cxI1FFoXtQ+EYjHKFsgHJOVJ5Ww8KZLRi+ZFH3O0mnodVGQ8hYupxgs7kOA
VstHzm8Sf4UCJL7WCWtgJMwnh9c48HQSZ2gatgPchuZC5+mw0qVfh/nDPP1++rQV
z2NfLMz9GCRElkXOyBAc5QrqlSv+b98s1QL7pPbNkEE4QfyxuMha1kgrHElKh9Ge
+vUx0hbNQXoVmn4c+eCXQDYc0jW5bGY5se/AuA5DVqkwL5Fonwi/iRSGdbOtHPS7
tozwv3vrW2JJSS2+FtyIWULtRPUk5OZSGKcAnm4f1MO1v3HpOE40pIVFxOvjZDe/
KDbiz7CsJHKZUM9DIAEA8M1YUDc7QevVRcXnTKCb+Qk=
`protect END_PROTECTED
