`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VFDi5+xMTU8ucTmzAAWnEDlzjPXnttDI1h8uwJDkIc8wi77pQtHppCxOyXetV6mQ
ktPQrd0wR/WbPaDYEqIJWqwDzAu+GRrEuF2j6b0yZUBbOVLPfyeOVoo+X5877qgu
XQYwPYuSRFoNuE+VJ5WsvtfHhJ1hsdnGiaP7jcJm/dzdMU5i/CDroLJJeQGOmM6V
K6rnHDbD7/GZctAPnPByFAio3lIDXvw20yLh7i34ng4BO3gMD30hKwnnU85v9Z/b
neYqYd389Sg0FraczSmw5D6YMHojLWbrJ3aNrR88QUIksYcw+rN0FlMUwATaAYs9
T8EAdf9YsPBuHuuKy+pvro2JMT68hHVGHQfeVkr3Hsejp1fxaxo9f8qOENurgWAt
BJ8mzmufGlxch3A3OeDlMDKLJ+l+OI3a4vJ//juPvrmqAYisUVSpQJ7PgNB8PnE0
CA2KwIqweXzcr6AoyffQXx8DLjo1G5365x/iCBKAIZfvo6mU66iO0GwdfhBljtIL
fX10JQI+/gWOtswGjh25oyZrVuJ4kewbGkyFZ5GuGCsWbAeuTe1taA/HSEgS8z75
6cKtbZk04z6K8UrqiH4NDu7bX0TSpnhS6ZSlOF3T2YpF2D+jkMK/jhLAXeaF87/0
eGGvYYfOZl5C99O/+V8zewUpGSo7u0A0Tra6/K9HzGkMVir+Ehy1hkgEoiUVr45o
6aVl0kbxBNMYXAb1SjEpOvyXhBwG0wpz5siDlDSM6ap1mF5odM5huIlKzuHs8q0n
NxfEJS9qNMLTyFsUlo7l40T69tieZku3B306JLp64Z/bdTA0qTYsx2CVxJ3ElQXR
hfFbIxiuNUd34DJl1akSRPoQsPo/jxVvcPQYdTJpCbI0RTlkBV2anrlWCLeV0hN4
4EnTAcVVrop5SsvhepuPQQ==
`protect END_PROTECTED
