`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N58ZeNVJwWuKTVIqNvinFp1kn+CEfx6hgAHuHK9TDXEnLTmWSOJZNEjQ9tfiqA6Z
TWjnH/8r6ySL2fjFDNwwFNEXPgyRchK7d9sTXdIB3rnw7FJQkIte14TQmLN91knb
95idb4A/r2s+g+FJc7eDAPSecdDLnvbjut58L614LRJze8KneZ0UzLZY67+BFQru
1Cjb6jf6nF/+OTE5RnGByf+khBRLH2SwbQy+wZj17ker6WPHDVQdx4GB32l3LwkK
kYFr4jT5XeOX3z3PtP3hucZ9b14v+V2vQPXSZhAwQtGo6Jr7tdNci8NhH4aoBuj7
WsPbXpI99UnDTeVL9EHqThZa0h3IvOoL6TTVGqW8OqUe9N5zgbtPO/gOFXhduooW
uYzVf7UEG6tQcHwHk/Iv04fakotUDVgodYpnWZLKBPZIzsNb5Qa5WIsdt35iENw0
w5BzXmpyGSxZsaG8PgYpLQDIOVmF1ku42yh/58lRoCsICSKLYD7lTneRRXIxAON8
r7i6tzA44+RAVAUJ4CpQ2Iuq/3N/omfBzIlRZSbpshU2mhtNtcGK95lyqq0tpKQi
I6B5t5mWRk3/l3R/x2RV3MNn6R8giSRsnOY91/y1eyRD6N17F5zJ/qVfx316rEzB
jj8I/FRdFQE3ziGfVWa9m4mInkX2IrS37En1w193EN6SBjLD7THlmeIM/aq4fFX0
aCgutI/s7fmJOSllkk//j1BCYSjaClraB36xrZPvU3PZbhZVIyu38NyJ5Zf/x4oc
hxBphddY7sEC0c1QW9VvSlg3lEBh/4QOSHKBQ7x07MNzSsTNZ2jX88gFmXDAhF4v
bcXoimzO4ixvf7jiGVusUapSOs+UN6waA1UhA0HUbfJ5+aX5Pyh7brmh67eLkBwF
S/1tSzdO8DvSFVitljxZqr32clcElHAaDUEhJNnW25uEstHtKoS71IM1SyUksApO
y3O0aGR5hRd2RHYUqd+zopZ/2x6mDgv8u8YgyR+p+xWCA2ossEDrXn/fJ3MQX9U8
EnpnxjtSnKrW1CE7ro3FmTRbyVCf6jqzf4rwWDIMLmqbhu23mGw1FRk2tyAMRcXN
SaJ2g18+fAsERKN6PQrrfdCAoxDT+39oYcTuHizJCNWV5yrDm1NNafbGnTXQiaOV
OHvZMyW1YK7RYeRjkKs5/d0VpBpOm73XnChhAhb6NNuRIOKlZ1enSz0RV7M9akn8
lsH18C8g2MW9xUM6ydwawssGE9syinLP4xnro37TLHbra6wkQxkrZmUDZyMloLCr
39IH+0cjaJh4YEkqZji0w6Q+b65kXtPMwYTZuFdAykraxgUQhXzHwm8ybrXhO7P0
dFNVoAPCeSDucT+3fwGsGRb1I62gBR1VHcyVdHR64mna7MhOMUt6oYf13aNLplSt
p+cqFbMGRLW4VQquCAxzazc++OXmXLCgBGabIRdwrjHtDbk/5RdFNyziH67+kqiY
IeeTpmSTr1h7P/v7FJ/H7+3UdUeykI8siG/APq4TbyGfUAUqxD3LIZtrGbdRprXP
8UNjXF0HUhL3KgRLr1FoS2oxerru2NuYX2dNlLiQw5MogMtzvayFkLePZt6RBpXI
DO5WzeJuB2wURKVtt0PVE34HKGN9Z1BVuUtM2gg0qjjbeEVPcpGV/2rEC1HS3RI9
MYCz1G3aNqTSZqmmV4N0AYtvyGQFRbEb2l31632rTroT3ESXaZO/PYewA9zzk3Br
wvNBiseexPtJ6osikBJdS2rtu+QJf9hgKQKKt16BzdI4uOIfalZLPkLJ/yxM5idg
GhLcLH0F+M6r9Am75ObMLaA/0U5C1Y6E9IyUdFEIkbP/wlaa/+j1/w0grsYuvWSv
QCZgEWnba4PTnnCJ+CCT6eyO7wB/pY66XlFoLn2uOubIY6AqfYwHEP3frgCRJzfx
7zfUU7QQAZu/NMkRRPp9/4s7xKUnTUH9NDBYGSCjWfgSmq4cOiY2Yz+P+IVpF1e0
3raAzzOgERDQoGGnX5dCg6KNCyV8h9XjEY8sMJ0TZslNdMxlxl3T/+hq8Ofx+Nrv
gfyuHW+Tk3F75Tv96vBbQn9cjV9hFEB6ZkJJ0bpwA5ja2JYtLTx6bcXcgRQrPQrk
ogG2vQbC1DAYoksfrwrAWtANUszTzs040RKWuHiUiqgKZvoGed1bG859wbeTQcPy
xp0icIZjd+1jHhYvuIpL4kOvwss+BuZiSpDwRXB6NPDr445s6xFQBxOAtjvsGiFQ
KZNoGD9m5rWlJKEwWyKyidh9r7CFox8CR+oJ8xXKrayqqmzscpLH5YCfRziZfmtk
wVu2txZ5H1StaLQ8DAo6jIT9umEBZ7jUJLmCRFJ6lU3EVYc+zB4Sk4d41SA4rXxz
PsaCudmJWLP6ki5Y9UNrjerJ4VUd1ny7dRLEzDdY5VQrIF0wYYWPRY0W0U6LVdBO
/OwcphUbVVGWhaNaoJWf/VfQLHAsyU1Y2yUcOiLTUmMcYqR4XW6ZchsuW9IBtwQl
pQp6r8N5/RGfsArxF0xr+QpxLFkjaXqRlEihq0ptfMFMSmxE6mmJ9GRGo9tTenFo
kHoj5FESzgE7HN7Zt1veXnrTMaBqR7nJK7LMOWbYrJvpCltaH5Lfx4QSoTcPX112
9miXVDCqAdlpy6QOzA2q7V288S0wr4F9OMiCVd2dZBCQbDhVfUVOz/GO/ryEwSan
Cozy1157TJqmX2mAj6iVfdf7j9O7I7cZRQ010v66bORyjh1C1fTD1xffLWZtti82
oYx4iQB9SH2lFZcmZBBAEKQsCx8GC+ljIFprebK1haB4ipxg92VkmiuQXVVk8RcZ
iKUOEaQ9fUpKUzyGMD+T2BNU0S6txjdpYgH3XFXwsvNPxjBpYChG+TedAsZct728
mnObD2EyOOgpMN7TnGnVXzopqPIID2Lj9sglzsJ9IQ7ANVMa4KG9D12GFpcDi4rd
tbYVfbf26I/kPRKmC0voKcyxJ0eEI6OrKcNUhj2OEiFY7OgsQfY6uqUhMEcL/B3X
8FAQFEPt/JUInpGZoXcpzZyZyk/fUiO1UI9AR3E6cArrROFzR1Vt6310Ehiccc4R
CpM6HSUV9wOMj2hdG6uHlKv49TYrCkdNsEnIfoNnPS33ZED79UrWLCb7lg9+HE+x
RJvY3CuitXuCSX07vFyoYU+3W8m/f4Nq3Dk2qHISfoAKkLefQI69kU4sh/Jgo0+6
yP0GdZYlfjnCDWLJzOgz6PtE2KCVoRe2NpZA+oL6aEUpJV+ceK5aXJo1uwORnvMC
3CWrwRvmd+AHI5artBJyXFjnyaRw0SmU17jtK0yy+hp1Th3WOVIbP+YJ0zW6qozp
0fulQreQuSaQaEYkH44LaAbnmg3iKBXfL6AxQmuzmvR2201cSvo6SksKtNbk5pdG
yUCAmpyUWhLs8Ddn/wU654B2lPttAKQgxhYMw+eMf8aumWXsd9UBuhdLFD5uWF+3
oFHdXzoS/uYTNV55aXgPPCc68fJiPQwedYIY/30XuvJ/f/TUgGOkKPaCisIBxjPv
bj4mBmUTGAMX4FChsHQjVbMYHasmL3OqGfEncxTCQCI9miMcDbthvuIcWbN0+TdW
8FXpFa0kWk0YluqXTznQ4Jed/JeGoG72VApprIFXnGdV6ZNTHixJR+hWrz4fNarK
NSziZ+jFeCFseczyYb+00qjZ5rwVSwrJuSQXOw2L41A2suyxpMDmGs8a+mR66bmx
vk1iQ95aKcKKfQ4Nid3OTDVl7r0xiOl4rseoEOzSABrCVyvRfZ3jUA1RYduw6sgY
mV8+b/jFshlvDJiClmzYKOkjavzplsIo4R2T/Q2BLTHjP71OB/5mQS481gOmc6tp
n3ug7s5Tr7rpwsRVPxg20te+SD1Fg8ElrawK27lIB8dY3WOupH/NodIbpq8VR8sW
pL96MJ93/g9+cQeYqjvVDjfJPIC4zsQoDJJ63CbchxBtAbg5BU67ZAXvbImrGrcu
dxvp3AH9GOGayEvbdWCGl431IROkFitC6QipICAGJNtUkCFb5CgEP8jOvLpCkwHj
82UQWQCw8IcPpL6JS4ZdbK9c9PGb9nWktxy8yIR0O0gx2h8/c4H7jhTvrnuLpSwz
MrsichFPyrOz++Q5EuromY9j+qCE29jokdm8R0QCYiuvXTtWMRQHi0BzKsJDwWEc
7EpvRXS3Uya4IIq6FuqbCeaRx5UWm+GZKQK/3rtm49EUjesjQH3PUYE7of/4+CzV
YGLtUG6pjGau0YaEp2BWTYZhnkSIGmkeoY8x5KCh/VfCrV+D6M+96FfuROM+PHf7
WfHH1EJCY3hiLPrwofVcGVwp+yK6Z/Yl2UDQgj5QKJdZKWch+F7jjoW9EKZoz9s6
Pm//213gZjdZ7F2SdInqpjtQjpN7nSKF3oeZBMZTg7tWAf30nGFbWKnAeaovN7M6
NCm1emLWEBQlQ2tV/sZIcr/vhoekR5vmnByagHKA3Su0XGRiWXhMgeAZWmyi+76m
dJksa2G0T6vmggUyE4kQ3NWlFwxy4y3GfFEsvlhF4TLNq14MzMsVgmTVtNq+TZZj
NZDkEkfUvPe+2aDAYTDM0USHSSCMyaQB8XXLag63j+bO4x76Qru7ovJ7EH9sE+Tr
YMnnejlKetoVDrv5Kt+549Cw2hoorOoSlVz6ByaNEL7+CSQ5TesJfKhBn+96SqnR
OdsxY9efmNdLJurET30NgKLinGuS5ozKK9I9m8lSW26Np8eB16xl7HBOCOELJHvd
ODf8glugUhIpu8jtTbujn2UC+gF/e8QZn+UWsebdFzhyngN8urwh47eQd2dXp1KY
W4REsEhjbU7v8lozLHTDjpm9icYp+XaO/24cBZ4dUQ27Eco2oOJI1CROxHM98hUw
iDCNR2ypbAicNl4347hEQI2emDZHJJDxZUbFpYuq3YS+Pt6KFEKcFF302DiLm8Ih
PcBSEX6nMNCSlHXy/XHQx7fv7jzmHKMiOnPjsCJCKEYEyUtyYTMng1W9x4zBI62z
i6mZJy5FUgRyj/TaIDeweJdtZKIinyV1AkkyIID4ZL8tEg5gIDt7gbzC96W3Mf6b
F3RWJjgtDyqIozdMzFtOOH1YgvvLEbGWbAJPJWMgoZ3w2mtW53xkhG9Jt4KZbvcW
g3sIZNTaJIg78QwCwwIsDpWqj48PqyBKnnNE3JSSxvxG1QXdzhNJhCSTF0EuVWwe
AYqk8E96yoQNq+J0bDK5zTk32z6fT69DD0xc5HTLmY/7UAyf3s7QmOfg/7n4Z6BH
4rTD5Oc5O0XW0M7z/txXvbVy+1JyqW9ZK/+2hicLAV8S5pvr+1G+3sTVDwoWNPlL
1ZibePJ2Px44Hyo86Edyg0UMFeaCRmG3N4hVFWP/GXJB6et7UVfz4MevHKxgpbqz
s+9W6W5fqKNnyRkP0q2id1ELctPZdfCj8KS/gr4OYBXMpIM0WGX5RU/BBcnpCw9E
dss2YsLfxCZznqHLc4+RqqZSgNdqDf+5dz/40u06M+j91eoIC+5P+ABguukvOMyD
5vdDJ/PF8u/pUo9EmKq4Nypt+5PQ06S62Okp/Blo3nfO+7q3oj848xbMHSLbprPa
KjjxfLOT27uIY6XsFH+KSw/Eho/mF7R/3QsWXQ3MquzFoSjgHPHMkqsBDHRwYgdB
hGhMMxfoMcLIy2hktzpZ2oWPOC+K/JjNHmAEbIQF7Og5FNdsphAfo6zsvWweeyWa
DKYfVVPlB94HT7C6Iu8gcxqecjQ4derEbzO3mpfpQ/IZpkRS07ytY5YjaMlWUCn8
ZljhlzHl06UEhPnCqTWTzXK7kebbrJmfNBLoMYxcBCd+aqgB+YMv+/uwX0Hsj1P/
YdIc2nefI2RVE0k1JsFajjM5CeMXZ5XTNI1icmz5Gp7cfye0uadU5jHTt7oaJE6+
eXWvqv+3Sh51P+LCECem2ufGvOtl4ZdNBM9RQ0VXqAuZIHkWz3l2DZScw4RUhEz8
GSm4IvixMI1AQGFiDlVfcs+x8d7BId9WONg39UQQbjzIESFt6kL+bNL1NCqMC1r/
kBvQmJOqy+tbnDfhIzGs3q1Dv6Zu2xGsGYfqVgT7zTNSeSzww1Ln30FeBKNW27RO
pugfrigOZ2tmV82SGxX+UIGoEMzycUz63SWWqQFKNUgjTOZByl6bWZRGD20neFhh
pysRjGKdQrrOvTeOkAyTU1HJKeGYXTcTsoUqFvqH+TryGqaOJT+jkzbLczBXtthq
UtXSnq8Q0+WC7fABVILCweUWtKSxEeIRMbOtCJH5LAVjDiHfkTpLXXF/ROoLopx7
8u2I/xpEdumh70xl3wrVXk5ZnuSnR4c3ueI/O8/6kKv+tu8mYo5dUvzFW9W0iGS/
y035n8GDTRrCd8fJhsjC2THW2JGMrZ59oHp4rirztgru6aURQ6lcMyFYVH4k4Pus
o65KP7aHzN4hZFCAZ/lJFBEpeWfKkySojjyb4DnSi/iXPCbia91FH+OV1Di9WJTc
YL/QQ21PiuQ6HQZRCQmxwVOhdlDdtKjdsb0o0DSmqUT89ovPyN2v3OAtDGjWA/w6
SqfwPaeNcvTGgXD1HjHq7dpLy1/oI7MdY2ZA5U6e58hQxgo78KxDiaLYxh/l/lmg
akmh0v0YitLTnII1lN5V2GKI9dv4BTHW8VdjKCtmsJDjijnWI0mH9oS9kVMOdscW
3nFTLP8covOErntnK70zYfQebheJ7PEy4cPVe2M+55X1s0hs5Ksq/JYzS1FRtwgp
9fM914nwOcPbNmY0uxBsfY9a1eXnvrNtUaHc7BTg2nm8YgOFIE+O0+sYxSUhDX78
D3GNV0Noi+SE1TeDWBP4rN9dL5z3oLGO9HnAWfdu+H/uRoPQqjqplUmpjcWYU3E0
SSyXSV+mDKRDhL71u22UjC20oS3iHGnfgNgfqe7NztARGvffd2nZ757PXHMpZod4
VcGzPRgV8SPnf3xbdzPyyUJQVJrtI3Cv9xqeV/XYLHXsrO8oGsiuM/cKEbBZ21RC
9gffUCOQIyTIi8pEDjfVPZWulTxVBaqhvwGIETfZ96TSOgZKN3AiIVyEI7XJTWCY
7+1zbfXN7wH3BoEKpXt/Njyo03IZnQ7ezH0mngl+NO3LwWIy4HsN/p31zlClCbPt
zn0fB6eNw0lZ8BMXzA20m0KAwZHXaOQmlgg4EGeF1NSxXaIx7IFsO64haCNw2XOq
yPbFa1VlbXlg9HZB2Xz1NxnEFOliiJWcSszBJtAHw92n5q4Q6tTs20SmQfcNJu1S
lIlcXceRRL7lE1BjXAXUALW5aNmRMApCrPDZizHh/Zd0rZwgCgcKJAti81ZPCi13
No0niL23OopPD3cZWdJ3T8zirPECQ8xm6oat+VXhi2uv7LiWJgBPaaYKix+B4od6
Xs2LTh2bMTd505mZD5BqgWtYriv42j5tRHXjhFS/76SSAUUa22iLesxD5nGoCH5Y
/cmMQ3qYuhw1y+V96NrWbiddikFkKshh0nwJXxIoSVgfwe97DoDzNcuEFWkHLv6R
jkRVKbDb4Xqk9ZqrukciNuUY727r2qDr+p1A+gmt2UitF850GYXHOSlZBUx2oob0
+ZF/iPT25z47aQKP1I2S5hu4O+ApfFLeLH0RBsulpxxkA8wnWBT14B70/UsNlzZm
hvHlG7ngkwoaAddc9UjoedzLpZMxoiOnIPNPqpb5t4WVywFDRMjBe6vP8ICXsp1Q
gjbQloF/d2SiRQawC2rX/vN7g9kqkVTNXBMLRR0k7I6s5rSMbc8JW3iphZPJSbEd
0i6HF9+82Qg2Tt4kZQrjCiAeePG5JT+AXV7Yu01SgC/qN/Je67G5B1/WnipDYcqG
Jc4JfDu0kZV9DKsN6IkgwdWSyh809iZX4MJggrrJccTdlH4mo1ABWazFQ4xbfx2+
wX795G8bFdDi4ICmMe7pRQKxDpCL1NJ8RawY41FP2u3TuAzNqGjiJShR8wjQzmeu
9G2kcyuueWFhRipTeFgFLQrBxn+8I7i19s8v8lLBp32Ck+A3BmJQ1CXYy2fBWE1N
+7FlgXmaKTYg7Q2CeHp1aHsDvQXiOr0VF+EyQvhIyfAjz4fp3W3F3hcdKiqaxLEB
KXWK3zynAj7EN6gXazTSUS5O0PiKXTgbiouqGLZN2iEUblo7aQvpJP9/icneA9No
MLa/Pa95cPNWXa2PC4bWQama56XLaBrgsmbTznaTJS/u9Amod/mQQHNjFYOskskC
d3wPVWk7erR3yfsDVkJuuwifsMK10qSUocVf18egcCH6TzFss+iuokUfWHdoOMDv
4ceVcpTR1DgKB9w0PkNyfSds3mpZyq6PP/dFhJuuC1ltTS5uRP9REPQ3Kv1eyWl0
1/yX4BrgUM8M7k/W6piUtW5a316Iwli3HiirA/pGLvNzlQUqySqyAeKrb9DNIwRf
I2Vdohn8840GmqkgiA/11Kr7p6kFoAOD7S0Rz8XBnyUF5a8yDSHoqV8//xGfLS6a
xvXFW6xwLvYGN4nsAp2eaoSMko8JRGWdxTOYfs7O+FxTcuVy8Hjzb5SCXRQUy3C+
W4Qmz/0NSwtKtYJq1pFjHeYergoyqloaXCEMDCdnE5unxOQrUNtAPjal6BIBTVkG
Yj6Cbxcjilay4FO5R+o/2RbqmBNtNksFZfRdWxiR01k3EY2HDzCcHM6vH7uDxbqy
L1D9nFYBjKRloV0m0g3L9oB5Gx0tlNBBNl0m4UeqMQkZa+wBeFmK0kI9fKt/5zrZ
MYCmkF2cKBcZQaBv3rh+Zm/LM8ej2aNNjQatMi3/p2bgRxBot7PNxF/uqV04yETu
+aJRHtbfCfpT+87ekJRggaejoJZlNbcijZvX80nGJbRPbxDJ9vIXQssMLcmJoRSp
Cv5FQ644zLbDZInukF3pS7RColJTgZ4pgXQoYx73uYwD216RMGWhfTOAFMbEJrCu
59ZdNgSaEFzErg+5Kl948PYjzfoZwpnL0LvJqpGV2mJ6/AYaTObUkT69VhBY0Dq4
N+WU9/wP9SjXM+FTairhXhWJXNqknPxF3P8KQZuH/TJkhchz4RYVMCqba2X8CuAf
eXzN3NKaIUq6Qonu5yD65oQ2o0ETLkvkcQ/wFRVDWhYIGvaZR69FxlETKwArqs2S
tKvVdsVcd4VEvss4AI+IuDiXff/O85Nc0KYJcfAJWcx560ocsYFYCW2N5sWgMKYd
W+eDl+fMU8Vptgt1V92jnGpu1/TqhDyOTN65gv+XlmnEB9BmvJbMXlCGP/kyd2ey
wigGeiHYjuQfyVXF6ap2O+rC7F5awHqpPHNK04q1MnGZg3sZbae36rBSZ/Qz1cIy
4jlE8ENME5twLqobFGAed3E66uyoW9f2fyF2F9NG5gBOmYWaQT0HucadkBmn1B9L
lQoz0Qm9u2GBOpx9p+l/+qHpXEe7PqgXoWZUFLxhFRNJ5hDwn+6d7jPRfBOjx1Py
T/L2BodEf8hkReeLGUdc1IXkFq6HM+WoNv7RsVDtHJemcyVZZnVNW+PuiufppYW1
FilvCOItd2bskxCn9gpe1+hFN6teGWGP0qHZdR7eTzIb0u12C9NQa2iHUEnAFCbf
fct4ntICMjsuG8FC81r4uBF9KZQ+UpvxAVJgioOgz6//WYJOGC1crKMdXDmJbh8t
hCEhJYwkAfbzQPp1OVj1mfJqhXIB1vD2E6HrM6VahE1AkaX5mvY40ReruEdzhOff
fVRdbM53pgaUGnW1hK/OAuZ1lWLjg0h3eN3Rp+s7/9aSVSRJk0cY0NPadRF5XYhq
x0fJ3ImDb+CXT2BuE5Sw5zEg2mpEBJ6wI0SsrGW3pxW7pQjWny5pDfOWHnfX9a3A
L/4Ju4cQwsMhaEh6CG+lDOnX7F0Txw06QSSdLDqP0wXU7GHol29DlA+LtCR04WUG
1pv+B/2wA8HZG+EP6q0kw/WMFQn/JahV1hR5oj8ZsYTMQqNe4TIc1pNWfFQk4DcU
gCNEurmg1P3Cao+sZ1wUTAeP0m3N4iRfXMKySTFVJJcApLXZuel4UeMrBi+gGmMK
NX4yE+KXZCHGb/vgMug/kIl/QtxlcPD4ZASzsZ5RGGKcerX8aslSB4ltXuoshkyg
29/fegnniDJMwxOJ7jaqTgV/HM6honU13GLFCQX6ZqXQpo5Me8kS4DOQ19Cd+IGb
X3N00CAiUCaFgNdexjeYlfFLNcBrjEOUEf8D60P3kVAQxh2NPWIF4+y/pspj3ELE
tZTNBa+N3WYL9P1uAFA2FqMOXl1VgGuP7S+gYpJ2wwTUpqKEZ5DvN8vq+02RubTq
Bk2JLXNKx9GWYnmKq1KyOj9H4N6wJHpzbu235A7SUVc17E2eOHGjjlH9tUMMAplq
JSMutYRD7TRZruoR0DjoELAwL21YwVHWOz9T3pLcW0ec5/7BT73Kr/BrFyyIBBxi
RwGRc8SqpQY6ZX57OhljbRus57aqCvsF2WZ/2go1LHRWErH8m3dzPUwLeDFr0djX
1/xE4D+P6N8iHxoYaVpzp+lHiyTqMf6I1xWGhzVlhZrkXRc3L/24+8N202DqJI5K
NJbxSgQU16TsbgttsIx59ETdilmgAYtsDBARUsJ71eE5sKnj1Pvp1hdWvJ9zxbUY
LzIZCoyq64DGgGuo5rvcE2wGSGgxgUoyZNL2BSjM404UujaBYEF+t7vEuAcFVovw
8xlxe3vfSzbRj3DtMa9QcDxk0fh8e/p89dplzU3F0AO5iPuU9txgvbiveKRFYDza
wUDYKsRyuG0DyrFE+bn/NdMptLn3fWjb7f0L61fDuXD1gfaZ4oFIe8cnHEa3aQw1
yO9Ha2ScU1uFI6ryxmJD3luye4vR8HFqgQarZQhdOvU2PT8kqVThjPd7dTIKACns
txaFcTOJIq/JwChaQGQweazs0ANEFDksDYBorg0k1I9azdcrbzqQvdNq11PgriT7
wooRrjtxQULccw1UYWjmNhg/Ia3ltGFwByexckUdOJPFBzV3EU5fmZ34627jYtMW
7BwIzKwbVBaPoxldlPOs35ZNmeZ2UNHjGAFCA4n2OmlLjWsqdFgn2ZLlMZMCz1Ob
YzW0UpYzWNTlJq/JyBFGUig38Xkf+r7fqVLuyPqqZvbUdTT7uvfgeKnEDrJAOOS5
P6Ge9hlPhVULVNlEw1E4AgnfpbTkd/l2y1/aovMS36jF7lgtACNQc8nxIdhuJ2uw
3pKXeH3uN/mAfoM6XPzMU+R3UnALItksaX52wuuZRGD2uc2OJL1qI9A25hMrb4/W
LUOgwnFzV5csl3TLWnNkJS+Y2wDkWFg6EJNAoKmyDlmPniJtA4EdA8SjtWS9aIMb
hWgp+65D7GZXuHjM7XaT8l1lsmqsHjKKeuAG561wL4vAMavnj2oAR0WXMML/xWrf
AgDKsx1gX4rNqkYqnXftT+oK5VXM5x8eVpKa+5qujpfGMVDyqcOkjs6ri7Tb+Z1D
SCzoHI9ssha6z4ZcpySp+rt0Vf5o13M8XWFS3cWfNNhmUxytytjjHYPkefQOK0/G
JnZ+ajvBzaXwsgCRz3qY1JKMY1/iSNwO7bK6E9rRXB5vOVVNEa9wbusgta3eqpKa
/sYKkZpU+HM7c4tmWFulb4TS2LVuNiEA2WqIPHKUSGG6g1g9jIrj5TFkrp2vlBGm
sXyDVdtRmHlacY3u/bpEVCET6vlsoBEVgIdlC2TFZYAt0I38YaeO3rf2Xx7qEUh1
mrE8icUxx9Q8HQJ2DilYaVhSV36POKlxi+Ar14Ktg2/BYF5Z/nzHWkpQGHmma3rx
2U257LcJy18CAmENRQ0vhDW9jAPwQChiJ8Rjk67d1wsP5NPQ+sx1IPP7pwwt0f2v
8NP48Kf1yv+N61k+43OtobvFJDFbAS6fRgMV5Ou/Hs/BjMleiVxswjgADZ5BdSk9
T3RdSIWtW6eJpKvtwDCeUXrQFpy8kgaXfhWj6G/Aj8woPCeEMYh2mxgwhttlTEHA
PfzBgphA+XzL7sN3m2hJKqGpIm5YI+CcYmBHrMWkDRjN1Vv4rkiTAYdzmFkrks3e
07P+nC9ncB9OUCXFHNSGtz431IK/aPcyxBKuEaNqcQ1pAIEqn8F3KLJhDin0+nBn
/vg9KE2UrCqoC4/j7rWAMZHqZOMejCtUKfJw5HslK5Hu+9wssjzxfL2efZbb6cBs
wJS4pGYouFFPA503ipZfhFLwiZcjBt/5RDzARJfhAA4KeXordX1CTXxDIfyZiY4K
JxYaIipnVirHLkbUGNnQdPmdWAY0lLCCX0MWh1Qmy6M0tSC73RpIdexW1uFwdYUH
GURRMLCjTF4mLZz70rQpp7JomCzuZisqwgN56UVV9bb0PV2FB8TlitM3cZU7gd/s
wNk+AvzFI+OOf6hMLNqcM35CrfZftkh0gYU6RBaBFoO58BeP1LkIiz3Sx5QGDLc1
+4ZenIcnNcQB2EO1BP4/FNDQyJuEkQIcbolEAJEgq8VKjwZLGPXWmTyRB01R/Eqc
PnkpSyjHoWpD62NhpW6DkTuM3QJ+6Ki4x47jByP+UUBO2kB+wO/gOZSFGGKV2sDg
3WAWUdeYDO4QQfmBx5b6R5F/ZCGL6WVt4ZBK1eDF7bGjQ+wvOd/Ns08x5SjV+3q1
3rU4bvDHff+Ec/qzDowBZnfvTcdF60GycrHIO8YMi73vmGSdHHvjk4OpCT/s/Ms6
4TyxmxbRU+daD5K82t1VyGB3XPlszxy8ytV/WHKmG5E+qWrzyslYtMy2MBJpH0Vr
UC26/fHSok69IRcQEmrWDLYNFveX34lmBvdAGg0GHiCLXlfSBrUlVlbJTifef7s/
UC7XJYcjWYhMogEfKn8R4Mm9WMNBsB5kb+kjcdo14kN4gDAWQX5j8ljVx1oeBKSq
PRgaAcXzB97alnFpVycLcujg9C1BPjMZTK/AZog8YfQ99BJ1IySU8JWv5hpcYMjw
jMgQklRIMR8gNloCzqua5IDK+nYX9LTMc/0XzecJ35kEGMw29bnVWfbTGoAMo9eu
KhxkyJktLFwremq8KVkDc6HX5RXwUxZKMiGWTJmD9PSC/jyV3mD8qtc4YcOFfiWn
zOnvB89EvTXShkbCUO6oO1ktH49pRlfiwE+GwyHwDMNwKQ4/ip14whmAGBZA5NnD
/BFksn03VuBCH3V/EXzP/EP33csQS1IYueOSxOF6xcQreppz2KLIs9QJDJTh8qZR
WQLQSPkjcnotokTw9e/MntfccTyVrxc3YJoh6ruPzns5ItbKX3jQ2/VeAyMnhl9a
X3cZKo0r0x7nw8HbIzWCK6wyEWrgxufDFeXzNst04EOh6CUaqRPT9m/wes2nyXmu
HjadU//e/l6lSaE17uVpUQvTkdG7flOr3x1pQgPZY6RuPprjQpTbloxnbYqPsmW9
kf2KNwBroSwOzZdlIr/xpP/B9HbsFcuC0ujemubIOK1D5fHJMgtswJT8Oycre8r/
CpQjzr67G17jUptKE4wCd7kZuEitNdHei5aLCPH/KY7T+zu1gdXZD5XX6XOFVdi1
f3c69PUiRmQxKzBTw8Qx44WsNJSe29LfJvXvujPC7kGvf5i6GmuUR0DwGkprcvMi
I1cHcGmZqgSlryNpklJuwTqj5ed7cbtWfkzX6oUrfCgLZ0xKHbYHSH+Dj/8akViL
HPa3RNdiw9Luu4ATB5/Nfz1LC4QGnTeBrssuhR/XKGLyzXqG/K+Sr6Ufsr+Bsnm8
aI0/lBGtTYI5pBUou0hsU3vcrUU7xCI5Z9yx5l50+oHYWWey0281ir64YLoHvUzb
V+14BIdrlX6nJN0xBZ+jkIQFJwSbAPw4UBeRRtlzysVe8WOVZ+88XjYtqd+OW9Ma
hWqlTdJ3VzkQx7vk/TEinsEjiQue0zcGZ+CQIHT0Jle7RqLHmgdVbbIgGhv6Wnzn
VIf81Ns8AlHJCdbo3m+xTrF1V3MFDzSf0y4f9WUymLVw3PoKpJtGtM7Iaga9tN+K
dOP3Vhl+C2UdNd8UBg/zVkX0N5bYhJf/n58v25Se1vxjV4+O+N7gDg1YJTSwcocF
mehecQI3nbygHFwrLQSBYOQ+AksC3yIqDY3gOJ1/3Dpxkj+AYIuQXmOporpJTR0n
5nkP4fuOdvjQhKxpdROBRKw5jvCoFoHx/RZXrXI5j15GSoQ+njDDCcxqyL4B2ejJ
W/ehHDVSK8SstmYNO2JG5lrgpe6EkiiTPGvnMK9u0Nj577nw5tCPbmYcIrfmX97D
jpERlzbT8uJ4bzxHy8yENJRawu2KVnIlq3Eh1Ui4G0so+M2e1tI01Iwc7nlURUAD
/UiV21Nsv9Q/orx/jDFgVwqehFTZfbkFCYDgHdyMktXqlLHiy7V8l+rjcDrBsyiG
CULxYTetMMuLsRHw+vI2C3b473Qkp7cZFWsQdEV+UU+jMvVPRPSg5Cigm6HfX9Ki
iNcN6s+OBMy9rSAQ+6qXq6ofNYW+i/ognd4rVcTr0wdQWWcSayTmc5q7obtpSK1x
tt/T6rtdvfEroCYyV6D26UNkWGTVgkvnNJnxL6gr+2uVSl3MBJy5o29Vr2QkAZK3
wv716LFE5u5XxO5G5l+pjR1zZ5C628JPW34n1R9B+nVrqWAjsNispYmECVz+WBKw
cQiIfD9oFhPJ8hLZCXDugCR1QHh0EGklT/ZBcE/YN1V3W7d5OHDpElcP61fsuc3p
CxXpWfYErth1pmCXyKZHiAMT6lmkUKYh2rdGyQRUqWqqsrWQHkgVd4ZHZAp8ZAw8
GJBbyZoMecZ0aQ3GhMkOy+KneD14uhQicyB18/0mILOHB7IvNR+EzMpDzPcDpJ8v
3XpnVfvNkACAOfIRtow2KwGCJXMHWXmzKtSMsvqtchv7VVx3t/3Hz8XMA8SrbY78
uWIVaPUQlSysEp2+Crsp4D2k+dwOeA8oOTNFvlnFHVnkDm5U/ASwo8teAPRjUNpa
k16WVyRuHMnSiCOp91KhWSG+g2Y1Ew9uBkBSFq1bTohVID1grgg9I5cpi43Mg1F0
B33B1Ml5j1IGzZl9rgQAWZ2goLLBFb4nr47pDiYC34Gqy8Jhw4KLKyVZoJWQdHPY
XIPfejELZpcVcK/6Kdnm3NEOaBx+jpAs/jFC6BPXxhUG+Zqqs2VhhmCzf1SOdCyX
g9JwLZDn7x4YrZEIA8rgtRgKGSYb7/bhgGOWOpdMXlBipsr2TFxj7dsvIRBRukZH
0mk4+iSplYBiZHKEWf6yoeXq/V1kwoEwvU8XVBGxThsEmjApzn8eoYs8qEXusvKE
QddwTHjdM3z27HWc1/3sHbPDgrseQin3EdRL6gd7WCuOBo8eUchIcFAtKrciQpqM
Hl4ryCLB8V39BZxLBJAMUaeXroWiZO0k3yk7lnfS41XKPLEDDDiSM1xq0Gj1wWik
Akh37dwUD5CFKMM/l0D1YmA+9QSykFd47DHqPFIqlSK223adwpRGJgWJr1nOnc8P
0BmhAsrJV/3IQKEc/PRxed51Z3kwy1pS93l9xhVCHsCFWASxRUloPoi5E2Mgby36
2/Z81uitYxztNPpvS2Fdzc7WNHtQbrYVfToj+jzKmiJN2hEFjRWYyuomHyANlpgr
uBMc17ZLAwfyVZzFSchV8DV3w5/lVfOA7lG6yO31Anol1mmnPcVPwXYZnVcPjPgS
q3vxzmhCjOIsslT/GWc484CR/vnXterv+A3zC5lMY+vW5fIslfTXkgKOe2W6PMZM
PxOpc+po90hcdtlWfGLhR6wFHM8Cy7P3HWfR/Bxatw7Soe/42bodrZVbr7PsWf3m
LtganLPDtbdEQLvd/Ses2Kah3sHWoqqaAe5vB6su4H4=
`protect END_PROTECTED
