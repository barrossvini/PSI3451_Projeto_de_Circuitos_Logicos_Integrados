`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GrKFSgkgrRP2Pb96kIlfImxssCHPMsUzIsVfVo60XjWDDBbR1uLaF4qoS0OUqBtV
/rJY1u2e6K5lbOsjpDe35HudrwpJMvWPAvP5qQo4ciXJqYh6zF+R+HX9OJloQCr3
1PkCJp6agi5du569KudtLlnn5fIoVrpyEBlECOxIBSUIXeR1nyIFRaGVvTMLQbXH
AMBj+ZEZBSQbN8MS/aV8lXchYAsMSrPEmYeZj0u4+5wLjroCR+eqVMpnm7/2VM6D
GBF132LBnJdVg5s7ZdJxkbUN5zhlUjYWefG4O90wLsaKgAnd3ZCJ6M8tFgkkCXKI
MMp04Fbm1pKYDsjGCgo5cQsdYlTBMzYAujLoK1ld0pl+PL2+V14uni6okHXOMLYc
tU2zDCHYDz0O/70tMMe5/jQI+ejnp2U8zz7w7IIPIgCDOw4mXM2+pYLgUDlVWI0A
A79kIlMeFmAlq7AxlfEll7OceTXkMnmwPa+1iac+mbsnJHZElxjj/bCUK+wzcTZH
AeLK3UVluCAJsg6k+kOpuXg8c8OGjUcBXGgrmo8n4O4WrCwahlGIA1XC42t1a/MB
6E+CWwwjYE4FhYN3q/0tYc24dIRsVdY6sDH6H1zwBK4U+8IwYeLmBJnQNR7mGn9D
Mp5gNY+p0Zh94CCfal+MMnu8a4I2Vjr2hu2U2a1gChw658aNq+1DxGvczxTuBHXq
WIuJTlRlHchBg/nCzUFAz0WijDHtEPNJb2Kex2p+W+OfmVUJ0W65T7H3HxSyExeh
1CR9g/FURriOx3bwpWsnRapiRcnoyx679Ax4lhYn2N5I6l32OzwNO25CyBYQ3wa2
NBuuU9NrrtIU7E9DPwRs58p2Ocd379zm7aLWUQ+YTJN5UWZRwpLKAheEinqHIenL
woitzPpNpKLlYoSPU8iN3m4/hdZJRMt4Uo/bwL7yE1oPDjgATAEK1veQQXMJFwNq
SDds5tAZJ6vSMHYhUkIfQ0GLl9nTiiEHU1ux2X1UJII9WrCxfA88FhgYqJpK47lr
bPRClaJLsP7H0lh0knlW5pbCg7C9FiezA+X6Tti9qDNuAiwp7d8nA+6EzrSEkjBj
gtIRloQxW7P2l9EILD59oBIJblk1sY7SV+T9tJfA2P7lKDHGas4TXiIFH5roxPsW
Xw5EeJZ2Sa+vHu0IhvvQDI96dHlr/4BzXhvTDYLH0XEvvC526Z3zErPBp+IFYj4+
EmeNjgs7Dh7lX4x+Jvz/ZXSt7wnEDJStpLiaN+vlvRU6nT/E55C66OZV54en//eh
DomdU1DBBivF9W6wbDfcQSBWw/3IDlxcPpgBgloRepCQM8Tld+YjGZJaT3zFUXOO
hOcibsNSYIDu/FrLJmYM29hW3+hvi/AVAlI94iflUUfcruKT/Hyn6thRU1JW4Aye
Cfak2eOq/ayxEqLOQCE3b+/4AeSKZMWPD16H14N4ajKa0LT6eHTPDiX/C4edaBa3
MIRoAqiCD4ywtYx2gjuNtRwj9kWOvbIqmVJ3e6yUm5uJqBiGUNwgl/kahqnzICCN
IO5DY3FemlhNaum7QmyxetxpuhpmXHgaqd23z869ojY+eQp6tV+5vtvwvezvFw+a
jcHQO7n5npafYeyh/5Y8IpLu4W8VUU0ce94lQFa45QsPBxAwCF7ORxG5hEnkpJAI
QrKKAEillMYo4QRS+BlphyGNVuhJbH3936+jgjYJdsXn+Qe7S45mLvKiuIgJlzii
ZeTehhPHtwOXd+cTHLJCSef2HODZMdmussB4wI7Zk2QTk4GH1Nm1VxhCs8n3Khrn
9WuMi4BIGnbYwD+1QCilifGhlzX/o5wetJQ2fWtryi3rIadYLKdNOPH9Qr27RPpy
pZum4iA+Fy/BLVqPt/+4BvIjYsL9BT9NgMmG1Psus8glD2CRl53w4pcYvKDN894F
cBsVmUG5GT/KUGlws9pLyVrqy295g/Pgj63Yx6m2MaXLAd8Td0msjKJmJsPiOGkD
Mkg9f4g4tepzjAjv5Hldhp5g4NYVNuRL6L6yal7aPYFj0neosfvWIVZs7639n7Lo
pWsAVK8wMu+1hxHY/GSX57HfWml1FCy5Qmz8hMlX2fe05jLQ67m02D9LyDM+tI0V
xjnJZw6Wlgl8B900RYub4+tMwFkSHWRP3WrsxeO5gjuDxOmlrbOzOhAbbs24zgeP
qjX6DUi8hEYJGQHrGLQqrVuTLNS/hso+l7wBBF+RTKYrCi/yu+ocoAyt2rD9M5Uy
Q1hi1EIOM9qzhvl7TjDcUxkG01s8BtddDPS/NUARPHcVkznXbuZvCIdxqFQLBoEl
TO1T/EScIU6V8ZIClfLbc9+V1kL0DTLTsYcK9bdoqm0xK++sBeJPa+lKic9AhErI
hCVr4F4DpZt1+AJ9wQKnPRYNCCwRXbzBY5GpdzpKJ00Q1A7MQBzonLA42JxW8q6b
gif4vXs5Se71eF5T+OI6m330HcB9obSDDcZxUIt51tXAzK0pLXB6/fzK7Pg8KB/D
1+W3xbtFycmeidNV6ndb55UKLgSCAWD1IH3rhJZ2hvrEh+ojwOrJZtujI+4cm5PY
FwuUEYJv2AkkZfcM37G90+JMM+G/lGg5f3QqccQCoraHbDSkWcLLlV1dHlJ/+bPk
TVtKWykriGfLCZXtLIxFXFr94Q3/cIg/IK+8Cx70mErgtLGPss5EBcTso4Wjq6Ko
E8whFOzX1KrUh9gE2cQHP2iVUJUy/325taT8hJNHysUs8JIecUIVpHsokNoWvacZ
YQIGgoZ9haKSdOQMrNZzpctCNRIjuHgxg/VVW2q6RzdbFxLi5RCuVJ0/FOibwx3M
Zj5RD6Lj/pgK8oLlRnPr1Jj4NYjszZIaceswal4aATnfZX2a4nyFrQJWepNMkszQ
A73iYKRIMO/NcPlgCmbLhMU1qNEWtunGBIf4uIYJZoLt3Dr1llNTdWtaZScVS1mc
Gh13EpK5Hd2/41JjkbCSd+5xJOMxIabeq/fQLjI/0tSgAO7PHumj8QIQq7lefkJp
BYghQmKYQskM4BHCVNMjTCGMjrzDhNcHsOh/OD5t7Qjy67tWr0eIiXCG2sGIAh7V
Rtk9ITZABpTpRDpRl2vrzI66fqOt7r/ZcXYbhPzyoQYiIMzXvODtYiqzB1OLwYAc
PQODYbacERoLtOJwoeMwTlQ12aQoDOefIBtAIXgW5GHBJNe6RBON3FZSvs4xMZ+j
XbleTjq/NpgRyYnoyByo7uDknLpvgkeJyNNf8NmID7i/6DU2LuJk1j3u+uj/diwR
1vHhlZZ065WilbhEzmKQGoTYZaEk6GrExZ7Z8aPoe5sWPJv/Ef9OdqLAiDk6XxLc
TfHLB2L9S3Ioz9ATyxSOQ8Lsl3nTvgjYq61GrE5mdVzN6GiRskvV6tXjPRENym/o
Fbs9z7Hb1JZQsJt5VW1b5Yas1IUWt+VJ9Nhk5uRR1G/xKWIwg/b87yZCjVtQTMxB
7F3ZjVvJ25UvaggtOGxRTQy0+DOCK/iKwlUx2L5XggInsUHexaytaj8CFVVIzHay
/BGi1rihS0R+alULGPOAZdyqD6YZYxTZnRguGj6NtBvwYku8X1oxq5OOrWCb4G6I
teasIfGe45RRstIAEkMOZYqxhZhxFyi4BBbdCdG0mAiIgekjbLqQuUpvInidvkxs
3fck9Rs+n34gAzhWOCE6HQs+MtncKbVAawAAwnhemjbtadppYdprla/O/y21bvmB
SlGbkZFAAYFfYBZ7jI290btqdbcYc2hMnw8Z2mPq9Yi8PN2OwxFaWncfY3dYCcN/
S+Z4J0JCHyX9JFzxTCWDU1m9zmDHKAfS9DdGXl9oif6Ia3cxQktYD0LaqJW61PKw
u2lpKv8tZsxmKZVj7GgnlZekSsE+9yGC7AkYi/3u0FChVqVjxk2/TzwV57cMx4x8
u6eaGUulNWL2PmI7y3C0RrTdJ/KVIqzOCPfQAV/vYF7BuxOXVhkfmfNlvFRd0RhB
7KEKmNhLgizgl1uwKCjD0qZKrZ7LPc0kXLSqYgF8eTIXBtOIzpdkt5Ydy/NpJzH+
XRCA4xcOYGzBve2ypP1M6lxLmavEFCFSqzdziag46q6L0dX9C9RJpbTpmojRoo9F
XOabsbL80fgSdYezWlm/qDvDdFRGe3fmuKShhV1OQN/RLUU5YoN8Wir/7rU3eRjW
e+jPJCLnYZvvjW5H0wT0sA08QiK2NYUJ7cm4/CSGxba4Upy/2hgsKjpN9rgVC+e2
PfIbKrPv9TH3aSMTlFLEoVoPP1Td0XY8D1thqRrc/vWvZkOiKujUxUHxlNgxs+QH
0W6zciFmlTSqhXioofKdXfZacSjG7/VAAI+ZxrPKqIrqZjnYt0/sA+8skB9s4EQ/
7Hemp9O2OZoDfkvceGnPSObV442Vf7BbHRkuYj0DMJiVbj2K75orhlVOJHaFwAfl
o6VoW1596pEWwdDFRBQYKvU8G3qO88UPw4QMvB2GV6MBMJuw7hBEX7EIEBcNZbDp
8X8zyUmhhbNZFortuOxIDI4tF7l1w/WTYMOF79b0so/F6KmXNy1AfIPuilZ4rU+j
UD14W/FHndduzWroXSIFj5D85Nt/pZa/zmlpNggrVZaU2vw/vJ73QI7DqdMETUDi
NjTLzPSRBZ0Ev6mJqdiGSJHsUAdC6b7TVfqR609WFgdJ0XoU+OcUAmlF+FzpesrP
jkg1nMtLdGd/RY22N8kwJkxMYGbFfPZQlMothGhJ2rqbEBrQr0mQdXldi8XGQQ78
9MT/KRsBDn3lVdvDAiKrRAlb5MZ/nd2Ux9kQjyR1jIj2SWjPO51SFWqeZIMMf110
e5bhgdPbeirnAygNfxqsOD40a7SmwZnuSP20zh/zPhq9lJhN6LUEHhMceEajrowC
6mFJOrOBFIezSaO30HI9Ux0tdDevb3RHrSBijlD/dRyQyCs2891KLWJLaWTqExhy
groLgg+sO1mrX2Nu5R9Ca/LDUHLk+7MdLtvKORSPWRGEBAiUmJzKneAjAcjgfaL2
LrsdGYhTMJXGSLcgRpHafPcXU0v+cewiiSF8o+cRTstAK5lu77TpG4jhr7niPXYf
mOi4o0a4Q25d0lLUy0uOedQZo3nQbJ0XrxFcnzWxSfWU9ByuEvY4hJtAPjhIA8zS
BBDiSWs79Kk4FRll/kU+ClWUNaW2VF6N3fu2+zY8iD+7RI+M5tIUZxBJ8bmRHIjy
zz3Z+WCaNHNpbfAAz3GmWfJyOXD3iZTB9gajciP/3K1E/hBZzWXqk3R7pfjRCwAL
/3cghTdl82kiK/EUHaJjDXsk8xEIKJZOrhqCEv7ZGMQSnXhd6c4GgnHGAyeDk5RW
qzotXEzlvotDIkDGuqlHy3ZCM1+Dgm9T431wd6OCOnMUC+2cnwGLdVIpBsOt2TnV
xH0NsJhh3rEZg+Puxv83VtL5Cn6niGd8jrqZrLEjApM9EwiwMhQRD8OGTqEHSdL7
cVWjTyyh3+OG0dfeAz9niQkE1bAWZbSLztSJoCv4JMmDHAO+2WNmLLzn3a2ARq2J
uGcErtMGBtMLS1eo29FVeCsYPrjxlWbPsS+fl4EKcnQo87IS/Dr6s1wBNETSqf5i
6k5X70n6F8o8dq9/D/+aGhoiNobtuhqzx9/5K0W4IeyWc1Pa3QWpfBWe2f/JZzCU
OyYEMCLEOzbcgCC/MqKg6mWQAs7gn6dRfPngUfXiW4i02a2P2jEWwub8fS2vLYzp
X0nFOTu9kV9mHdJUklMnH1Zv26zm3II42A3Tbttb/fmZ/HmXca8Yr5GVwiZJJKMz
btLBRpR6DjDIzSV6aM8uUKmbjZe7uYl66vzupB26uXIifPNfzB00Qs+WNQ/nihtL
vu66hTKvqweDl9Xa/sK7Ml7v+84bXIyxRiw6rRXDiayPqmYlDVmdswGBS/TLukUd
sEQ+H5NJAYAW/wU0tWJaXPqvizD1g5FpJ9pKOmp9T4653/LbKFlgR7hwIwNyRJAM
2QQDfT54RwemVreLjszdH0beO5pTWoDjLhyIJ+j87j+xIinhu6s61CaK8aJhAP71
1GZDyXXSJ9aUTs/8Z4HFQxfs1+xCeAJ8fN/mk6LCEORRR0+E99thgqQOrXHfsK6d
n87Ww5YTVRl9a92XwsLCkOvhdkX1P7PRlDWHWkRXMP7kUii//REC6kVKrcouXSTu
qzcAG9zvzjBzJh92D3bqPx5CdW7rxNqUMIAelny7mG2M7vW7ZZWe8fqgbASA/aOV
b+ViUQtmJFDSkcccykmeQcyjZf9JaDTKCiC+wi0PgvDOR+MrRvhyZc8I7MtGOU5/
6G7gl/+IsglgVT8z93jHxpHlRyE3ZEpmpCMu6PTkUsW0taTNT+pBgp3KOvpaf/Op
l72Pobyfxmqlj6sn8xrIL+MwtK8exe2+CGhS392nwH/87XjmM8ku8A5zTKCiIkar
PzSze/MZcBj9YXlM4BvOCTfoEMATz9j2Snm8kXBu/vOCyKNDGBs+dr85mcRBuD0K
C+dzRMCvFhoibkzqqsBwqOyF7K57FOkMFaVHwhhcU5A0se+KTQ+cBSpLZmlfXETR
XeMCrlaRsmMa1K/CsQOsO9VsTcBGUL52kkwRm5VeB4jy8UM4vu+BDzBXblHrZncy
plr/OekBJqUX/HGD67dCYrbiN1s6WR44TJhzcpvuT04OkeGpHGAfRwZGLhUXsi8e
9jvlB6JHQEnRQ9JSPtJdaQ9p/N2QlCH1P4HTRTIXn/2U3CDTP8DqDi/FPuaN3fSa
/C+F476/8PwCHl9n2sw5+yP6b/nvOOKvyDsT7E6UV5q4JOpCirHjqx1d7IRPGFdc
M1pPUmWsa4UijtMmQ3+c1Qo2ypncRGZcsfmDP38ZfGuwvUut9ljJUScli/0gEwOe
YLDS+Gdsesey+ubaK0HLH/58837/NFvQw+RBYd+3S9XYPyM5D11exPr3TmwrPret
+KFJbVO91TRXMhQbth0+DUxY/YWMUJ8NzKwKXSoBw60WDpbAjbKCr+XVKSn0j3ep
0yTVsZDUdhV5Fz/KdZE4w7V4tQ4daWFb52GbMfuAEOAm8n+C2jcuwnnf7jdFmACr
FcSf20zjLuS1yH8elBr+RUJ6+TX+81NByGc16jKnGCshCsXAHoO+nRu8p/82tGt8
JlSRKqjKqsv3m8DpP2brE8zSH9QGUGdsb11Z6k2bPGX2+3LUHnqkVROImfWYfIT2
ULb1sMLSLdJY2L65Q10vugErBnH6hZhH8EH3Q4RVCiS9KS0KcGh9YYIfLaLm8puK
CIpTm0eQBjSXHZTcBemjXxNk7xhZGslscDlbfu4G4mUBgLQwIuPsPLfvzbqwgn0O
p5Dd6ERfo9qIIMqBU+Ag8pL6wnWCoV2PTuM1WECi43GMTc7bnYnqdSdrNGCvX89F
K1EA5sOMtnkfkzNM6GYg+vhyQ5B3O6ZC9/IWHEM9uw9fQELu7Ue8A2OcEMEyht2K
7lwV9BXxbUxepEUy2rC4sSRNYdPzGp5L/0NDQiaKKbWOddoxOtciZFW9hM1NFfU8
lojFJoTpeh+ERyZZAM/pfw36VjGDCRU6oLClz2C09VXxrYg331efsa3z6I7kOes5
dHuDAdpawxH05oyJz2BXp6hdS1hCH3JgjcjHwoR9AH4wf2Il9Bz+npjFkiTzxzPk
9drMgBrNxjBzuz03Rh+sY5UEoTkCP7yjcx6pxpoj4fGu1zgGt+ZeuVSBfzlh2zPE
ujC22OgKJfJUTSMhJqFKP3YEmwEmZ+azxs4PLse6xu5KDA34Zdmr2xSWPGq8ZJGH
aLxjuov6Rj3IzOn+KvUOKkZc92WIDS1wDM5eHT5I2dMaZBI2YF0sJF31qjia6U7l
YpyYGJkJc+68n1GSxWyy0rfie9MY3j1zLSbvm8DTblN+phIyBF5TJT8L71buNTWe
JwtT3Tzu9PAcMjEsDWfUw/lNvlEnzXDUPpDQOSLvgis4mhQrw184NKiuhkBzJjZt
seZKoyayyG7YD03oUDCdClu4mdJPQRK3itq9P+qDX+SeEI4IRFHX3KAH6PHdaXam
mTpV4cko90NQzmtNqnRnMPN50vvBsoKXAy09MVYUZbNH2k4aBGrmaMZZjSlZ8oxa
lEyxudY/Q+ZjTE9X7oV2+u+EIqs1ifYyz9SI6ceiJOw5/GTak+gRDTodmMPmCpbU
yb/VPPnuyxMlYVRv5p4jzzb3p90UPDjG9jy5CyPJe/bLsg+ey1aJWuiOtQo5vF1A
hLwBrcVTTqV7CMIv9ZXgLCy9R43O6nHNGHErr4DhzoQVcs4OamKgnekQGCQJJYjr
tdfMI5QuSu9EONueAQ4uTecwocJgooBjCqFks2Hs7LBusSvZXBrmeVe6ahNgJbjq
vJHkm3yO6lZvtjyrXs2pVBun0/IjzP4ANQjq7Y1Lff5YMWZC2WB/Wz/oaJrDM/q5
OQInlWudjW83O3G3ODkRwxokuY8R9XtOuZc/hT44DZd1z9lFKQ6scOcCpFJmUIAN
eK5ife2UAR8Od6tVsYBRJw33J9qGfD4ZF05KCxJ+CptlSkiFxkeqTOwEfu2/e47T
d1qZpFMJE5RFVuc+uayvPF0MQcIMnf6Bt7xOYiIbYbhVwDyjRkj3sk0FOaNDlMsb
51Ccc9HXiDlV+NUmKPrTU5LLp0Ix0ijkwG+9stUzDteONP/0xPD1do70iJGEwYAA
UI+kva6+vU8r2R0Ur1upyHQ/0JNgzRHffLNFGB+k2CkhDaWznyyJjFID9sz7Qo8g
N4CiviZFT1G299uZS6buqxAEepEvJskiI97mljmleO25s1p3mslcgxmtGpUrpqIo
gWs+jsy9DJmxyUOY6e08/XcCHm2iUwnA5w4rEwgZtfu08SzvZRtIgrnk67L1it3O
TlQvsgQUG1uYCJkwJWFyTEVcLNRarLdXBcqXP1Lsjjf1htw6x6vdaMnm9xYmeFAi
DRURt0abOLqVeH1OA08NPfn/rW3USAEqJ9p3B9Di9bpA7HqKtGIzufABto1+srRo
oPBd1TSuW2V09NLhD8xFQiQiVTvfzV1VpRD+oDEx4nKBW1IWFvOIMLksvdZDbD51
NEiEYIslQv7TZhjbbdsWPf4/oxB2fWz1RSe+n7bDV89EvYzDlYzh9uXCd4UlqDhz
Ud45sl2z2oouttpkmb/4KV/UhX1g2Y6pWbUxaaEGyASP2PoBkW1FYFtujIq3GYhV
5ZrHIzfoj47iHMZgiL3wbEnBJ92UBo8PB7E5u2cffpyH/9c8LpNJ4DCKK+9Aagrx
30VVPE1LcptEl2pMaU+roZP+G3Iw4umoYjl8NuMEHtevIo/yfnPGtv741gNhcfTY
Z249kmyxES+erOTtDziQ3nQ+4sXQ7r76n6Gs8Etb0Ncq5SBGO306didV8Y+5Viln
Y7IiH8yBL7xfAYJkXHtXJdLof3Y+XqnuQZL2q9JIPC/aZjESprVWE4wVqirdhu/M
qN5a4/7J02GD7FIzh1jvEEwoVwKvmk+ujCkxgY3GaBD9gfhCQ/aMktMbggu0hJ/B
WTFCBiW+i8d9tPWekpgq7gD6F4BO354o8sptRinKCSa74Na1G2Ycu9ChO9i0BORc
YjUdSHzOCCkX/SpTPN9w19pGx0mGuMTQB5mZKkaydWS3wPfZH9ugbKP2s6MByIp7
VdK1TGCYzmrPNcdAayaDfmA2pKhd2sBR4jczv/IjtWmxxb7b9NEErGUlmm0QXFvn
wEBgbCYx/tHFMlPVULtwg4JgysYTjDa9p7YigD2VsSmQpGsaeUij/3f12Sl/CoiQ
pNy02LDz4Epz4o39uKbxTDzp9T+PuW4fJc16GyPXTW7uFocxyOdSKXzqMI0EH1OM
OdmEEqnULgQg2Gs6Kx7WBE/fQX39+jqEamFwH35/rTP/KaB4ihfkelJddl/kGZFt
LYNqzI3TGQNQ7yunHScuW2ot7HLuk61eFzUfK8FChJckitMpjV7w+SoVdKp1ABDf
fl1Dg/qxeItV+6kl330A3HdcgwtDkFZdGVY5/a4loTeOY43icr3FynRprVlsumoe
9ey27dsZUnBisw3DvXyZoQHSpHewRVrkuU5bq6emiQMEPCym5C9lp52kLYC3S9sk
/HhDSu7/IGVCTpoy7JhSVUTtooT/mJ1loumxskKcgF/iBEZurp36VUnv8F1MYYEt
J6n35kFbuRBy9XlMMi4NU8h2XaPWEMQ7iZsQAuiuTpVTJgYWmwnxE1GJyRH1zBPC
MwTggLGP8C0HKZEMfzIrbtRYlvLeFp9IP4TL0bhlduV8cJ8wVgaofWLxy9ljBo+X
nNjopUkzqcL6m93ynbsBiGNw0X/IOzrHgVYPn+S/EqMwTAdY1S9coz+jEYuVT9me
ywnEULHXcz6HZZNZcUcp//WmqJ4gNX35QD5KG28/zbbo27gadeosOtJW/HODI9+W
wv6KxujwXD26PW8vnxdIUXknIb98Bvsmn1z6Pb6+Ic2te/YTLIScq0RcPSeGOtsH
CmfpBE6KbTTpENjNvafWlqpPYBVuhnRVwu8KhDTf1sl5WBYZrS8WBB7fiD4iVu6v
3QdFVw5zUvQIudvJI5Uylo96+z6nANr2w6r/bpI6nJnvP1u7Q+cSfiiGocw6bxWh
G+jTm8iKP0VHYQfHBbg0tDPpGY4S7QmCZMEa1P+HyLvaKYqRuU9ofMRAtCquyWIz
VZFM5Rfwj7uiizRXMF0xyV5mOjUcBXA5Hx3er5Yf8cYlF0NpsKWmAt420V1JgZ+v
I34+TBb178rozKJvtLwannkOPtn5hTIoyA0uKur7crtaf9c5Ew5wJt8weMAdCy4v
NJI1NUWDufDF6vtIw6cpRbNrx0WeStLHI2eknAZrNUzmAuSDuXDk6MjjXdC3Z+C6
HtBBaX0hdgTkKdWHxvff0yLQAfbL2fQBq0LbGbLILI5WSLx0bmj8NBe53jXKWbnd
+tKujH2u9OMu+QDTaixVFyVgiZfCqDvfTdJFJctnKOqqOdXSC0v0Q8RUZugScfQh
zI1DItdMbNK6lckfeutokDq/sdN9AWA7MWAiVwP7WC0oatrTCmiRV/XzEYWadCoV
pOICetxp/IG4Y6HvxBEadL9bMNnm4E9ENTpkR7/3nriHpEgc80Cfuq79nospjRan
fZ48E7JwXlgYYK/ficwERL5goj00dl8MbXPW4DQrFAmC7IehYcV/MwFBwiSDTnE4
i+GdLVLsr/mdCqWvwdHzg5Pn6APhdZwa9qrGPkWzpp17VM2uA/JvJiXgb7AA+rAm
jb5WYSfb7V80FyY3JrKn4vVJKXhX0jRO9CuoxqDdB0Lv977OqB7fFb/7VnXAd5gW
daTQDbUFsvVOMSZMlab1VWpj5ILH7GQQpk++0lN06n8BEzLwtmi+Dz3Of2I/5Zaa
UK/w5/rquaOG8PEk/E/6u+7hLiD2gmLipkxnyV/ktJxuT8ut8EHA2dkSM/CLJkpR
UHUW42luboGbrPDmil4Rf7DpAv11x42QA/SRTZMt0iBrijgpV8df1Nfe1Tqoqvwe
IE2D30yeC+w4INnPTx7Fpb9XD+LetKGGw71jzPU5gMQcGjYym3tp48ERKnmZkbGQ
aS9n85d2Xq8RQ+iDXOUHn63M+mnSWdi9Ji5npvNQfh9H/Ig/4058T2ae+EiQ9BDy
xZpxFiwSLnxYLi+KUNe177+EjggdMv1RLkDyFl+RuCR8Ib/Lz1rc1XzGlaBt18wi
1nqXTfCnYn2R3QySGgk2dJbCMimoMUlSknrno0f+HA67EBQGoGVwaLZiE71vJtkL
2r3nKC3jzhlvjOQKsejU6O6MZ0+uIW6lKuX7D5C21h7ZFSS1IiGZvEX8GXq/ocRv
ZyxgntvuEP6YiaF0SdWfpVcISoJiiMgjjpUAvqI70Ab6+RDzScJ0gV/HukAx++33
43Xsv2WpaR0LKevqhq/6y/J607Si7re9u67ouOKEtxXxxipWl3xhwCpMUOHZYOAi
jyslQDXdoB7uJzNyGlfMYgZHOFWUqtSvgTENS3DYrHPtN5F9vQY/OKHIRnaUgI/x
j2mqDbxsbUenOziHT51emeocRdUek4DNbkkZeGAz9naN5exZk9e4uMj55hxwMyUT
HiT8ZfHxXAxDfm3ie88d+pJ6wRGCMKWodjKS1xiVFSg+4laH/1BLF88XeRByD9PT
8LhIB9A15ADd2OawxnUq99wqbRwqfTHC1tXUZlrM5/kME285HQ4Tvf8kYZvErcCN
V0znfhUW0j8ho1dPIngeNUL3LVvvVCjy/clMAmqZAM2sHr5mhr6YaPMWIrnzdI93
qQzv7jli0H41CHCZrHYxls62tudNx89i9IeOngAI+84uuVD7/F0xI6yho9zquOI5
BE9BukMXpzCLKD0XA+2iOJAsMfGO9MxaKNFhZ+hIwKA37d7W+O1Pd0CEG09ohhwR
UzA2clFZL7wEdVMciflMKsUyDUx/XUi9/+XLm7/yAt1qZAaoW8JTqNC+c1u7xu0g
JaqH08sBCJxKThCTpGRlAf1LQb23cXOyoEJywcBMyeP9hWNydhoAI+PoRSOS08lU
iSzz+7ijvjtwcuK3BfgKIjeJxr4YIrVQedXpuodLPq8OTC+bJMA9LZXZyjyRia5f
2cHotWWAgnWCbwoAnHDA4XzItZ+IGfZywz7wUh3Y0r6QRv8t0exrfcACTmxRNFAG
L/CLqa50gpFCAKXDJgwa38dDTgNdDt42DebFXdjBk0loSlntlSwMICgZIqj7xsT5
y1HrGyvEoicFqy5PZb0s4YiOzLSCC8wxNE1OopWdy5FYVOwHAJcommojfFunkDqS
uykWVvp4j/1AXMqiUKdgzQyY6SjliLyqQJy30xJX06/YLznH1iuhxuCvL2PecjD2
dOiHnYP1isWad78MKqVurVOQSzmGu5WFKGMbhIoyGbcpKRYhPNkwMj7KjyEyWaWd
dDP/uCcYoXybZiRYVfXHWMBkmr2ZWk5foDWLao1P1xSfHo2DqNQZI7JoI6WU1LVu
moe4oNlTISwfSldrzBcKkm04R2Tv83VxRxlMBxVEBemvfiuLUqJn0diptt7PA0JG
zugP1C9sJR+KeVFjSuqESLO+9tR0cltQdORNWuHr9MS58YRq2/i0MozHCDGm1zXZ
DeCHruvQSFxoB87busSgCrNBgkK3ay760LICjRc0vIrOjBo6Uj3zz0gMQOLxB3Vz
wpZ+94xL/9cpLwOpOOd5b08kV3YZ0f6TEAPhbTlsKPYrcy8ZmBztbrIa1pZ/ptWv
njSw9f3pzMzp4muMBDBk3Qnt8jJ2z8P9NElYO9M4dOZTDc/ogrXVTMpS+0x6Wb4f
cIkOYcaYplJcG/QhRhfYWsKVrMdl6C95GBS7wbeoWDFAtCIYAYjU8pDXk6xScDoi
mv+gaH0gwoZwkLmwRoi9oNnWF67oR6dI2Jh3O+yKnN/0iSwjX3dnbdGCYhiDnkAg
jiLd7yMKS3P6HX2vOdPp3I+zAOgIIZRF1hjyCwpGPkA/ph3Bj/Kp0RI0fVTKAxic
PSxxbuG6jxeH6951FUrJTsmLy83ll1Xs7BXUjrAuoUVzqlrcRpVrqpXz6iCa8R2W
eS7yKTwArSYDto6UrjyVY12SoqRc+wDg2SL61V+u4cHuVkp8Cl3MmNO0Xfefs/PO
zkfj62I7SmJybNKhteUmlUxWLfX8BdHTPsU4pqnsUg2KDgtYPYicnXWHRbN0WyKS
87oICsXlEnBFlBtSFVWD2rHyjjTgz/n6A4jnC90kEae/xoNq5BLEmDJDiAgknZco
ukzY3v/0L5Htn6bUgdqq20Z3QRrotBCOvAzHgrJfRP6vcAPeSyk1BQZToKYhRvjZ
8CMEnfrO44hwfoz1LJp7SLbPeVXw3MA+lFkp7Jfu7Gr4/jjRoQ64icjG1PZe+YbD
6DgKqq2Nu1mTI7UEXzIu8cExKFzwYJJeEbd6fX236YF4tNixu2YxV+ydjNDmvokF
Dz0Zvs9Y/tO1JPN07CRkebScSn9e4wg2TkQQTNBSeLohR7zC7Bjn0/v9rSoNsehS
/B1PzEqYcK1Mk/gBlLHoO7Qe9l/LjDl5alhLs/6YhYftrzKryirgCQMRZsX/35wJ
SstI5dLVmlvOtAkz0sjopoRw2Mq/W9nmLB+2wgOwWysZLNUVxLmouhRAE6wzT85Z
fuorLv6UI/BTlKE5kgiJP6FKUFA5wqEUjotlxuQxvcgkdL7jB7QwBvbgapR+gzXW
lMpS+2I768kdYVKF9CAu9w6OWXWfWU2RyXCRPm/Ij03e9PVgvRNNynwPfL4oFkyd
H8dAbfg26iBnRta//lrGSvbLpTqmpbZhCo0ukJpqoEYDvtu7d0yM0vcV1cJlqBKZ
bxGtjw6Yk4SMCNEzcG16SfAnQhWZVjaKK92Ft0768Rm+odu1Rp42jqzBapgwG1wx
zONecnr2BWweMqzcd7R8ETTzCutQfEb/+XBKaBFcKm2NkDbLhicmwtOplxUBYcnC
PP8yjoDD4YAe+9dnuxkUsQmHJplRtBOlUx2n7iRazHQjiR102ghvWbxE+dj9sHg2
GXYEcT1U8SAfdje2AfPeFin//eYU50KezdLKgqgVCVqmQe3J3744tL6LIDbRD5hX
8cKrvpxcKo5hbDfV5toqoeRtnzTdmtX1kE6wdow/XAvBxpQIoSk2uPDqKlu2blO6
o5ERXEmARcQNOIov8Vtx0miYFZZtY3BgP55vg0g9OLtUfYY6PNTlfnXddjCXWVFn
tyPSRZnTft4wMc90canyGJWLREV5PK3/8kQgmhLsWYBsq34wZuvUwmRa6t4aY32a
18hvwIusqqKee8oVENnf7/TVRLKWEpdwMVRgOp/kEQ9KovqLsSdsaKrPWaume5or
t394oyA71F+EtE5BfpGdI3qrgUwy+5A72BhQiBuNAVjMAf4J+/yhCNJ4VRHyhdOk
mitlrLlbEcoY7BgYWNSny80jcEQThJKSWSZusXxSMi/eKUuCMttiJ9zSdqwowEO0
y2sr+Elmf8eGQWMxcYQ0IeK4n4AnMBhgbg6AVMm/Oatt7MTJQ2/bsmu5hNN0xFI8
Wt7wXiYwQEWC5HoHqH8dc3kJlPTn4FSPH+Xn/YIhK4SmvaAjKXQhsNX5ooEJkWZe
52J17jGDEsbHbJSQ/3T836SegjbrhFl8Lx7qfrbBTi4mFihDTh+iMKoR9tLhJInQ
fGfnbXEtc8xh6gN4CWKdPCj8fc3UluIQ41PLkIL0X4bPTsBaT64qDmmQRw/5KT/G
U5nqmYEZVcrBv3FcpsuQLntGUMgDbd3M0PRsdqENzl3Neiaw3050IzG9ik8XKmvs
peuS5lkZNl5d+hlq/nETuHyfqaZNByKA5FPVH8rkJVtG+cKbSq+Zzrtk7z2PlGZj
wkP+4Y8nUDm4QZnT5oLo1cVXSOMX9vwyM/RqDt+KUbS1FhuY2MTqPmIoKQx/5xGh
Q48afP1c9vADqBiTzEgrVbL58TkGiMVSs6YUYGF+4vnG/X79c2ujC9n+xACdEmjp
doWyidwbgzpn1+ChPE7JZ9cxkMrBOYWocxepZxs9Cq/gwD2cDyOE5/8h+GOXGYs5
rEEBp8svXCf6sl6Lh4sZX1h/Tb86fgh2yjhyH1hi+a1KUgLVKsKMjwMFP1aCaZAt
PPZkP+cfvMlwe++P3CjrJlNlkevHy/ZuboO3lhpQ5Dhb+xtejMvTFn9xK9/HuuaJ
5fbEP/AboD3gwai4zo+VdrEt92W0Wd27MAtGXt1Y1eeT6v+5/r7kfF+eg7zmW9N1
cLi+fKD2CHFSKsyATSpRRmzKtbhbo9xGTFG/a4FBu3vnIU6KkL0vE5hJFdSzfobE
eQwPx9Xnuar/6PWy44y+VOdI3fHui0DHT9AkTCg9Ol29CDXYKl8yVlaTUKCnyLS2
dl7H+WrcTN4iajQkevP3mnTmyutDGTG7o135qIF2i8LrUbH5Igd89rTqr9GNR5+s
8VYVGPGStzZ9ABA8c2Ln+i30OzRXJ9ckhzuFGrcLZ71TB40TsjkJqDknmVfOL983
yW+0ziMmWBRxi6ysnUgLIaEe1RPzDEhHa/JTkzsRhYoZCT0BobAFlAUxsgmwZdyq
oN55vqg+mb9TgK99cC89QlBnka0Kb/Y1eyv5rgpPeLS4acncvSnL5Gjw//8GdlSy
gsJAMKluetN9VpsIOepkkBCgwLjkcxztOucAo8NJOGFfwNFeQ3GCtCvPE7fTKTrk
EtgwuWded1PtxCg0QS5ZV6mrnF8jufM6BfJ3oyORpWE5yxkqGHu8L78D4Ium7/WQ
nuEFjHE9YhNllxD3Ug6kENZj8ijLx5uD4q99hAl3wlc33fWqc86mcKIEtGykMgde
qXZwDimfjMykoQtBTcdXtfdIzjNYI4BQsPlWbl/Re1udoqUb0arVqM9VXLXMneDd
mI++yCFnn2b2mKeFT4yVdY7qY5t0h/6USW6zZ9gGJtYu1RSZYehOgTxhW4Lko/iU
82u9Orii+kaqXQaI4gjkhRshwFns2+oYEPOxuCHmVujQyeYELnC1wgnBhmMuFek5
ItFIPZUitgm+rzgRrOXC6iGey7amxaMPLqE+siORb4WAXGWLgDqTi3eTcOYGA9t1
UcbPNT0G7SxAhkkBizm/1fV6I8y6JgcKw5iTu+52ONVbh2rOSqO7VMBu0xsUDXOB
F46NvErKnAikEyB5ALZVxuhA0lMj12YATCnNEKcu2pBTmcRlSiFiCx0v5AB2gF5G
GcCTtZ3WDqeKecRGsv/3Tp8NMr62sLTpa+P+WAo9OCriRM+VxECmxF4Ju5VuEueX
YZ564fKMO9s+ScNnV3HesnYhLitB/PAPRTxRocIuUt8+7sH9ha0yJ6OEtdsSZ4Kp
69Vyqkch2fKlGTP9td2YFN/61c+WANBxG3HPDpYdyhwHGi3RCTYWSn5dDjIXBLsC
C8OG4OGY9VThSj+3lYXxgQQ3dlhMPhMdphmVMGe4SAbWC9eCZ8z2xAJ0RZDR7GoR
6KCgWMWbSWs+YAiH5S44QVFpSfQI1tZnNVfvA7YsYwlzdNP/0t69XHPv8SUIjkM/
FOVmcogijuDpYkM0oFbcxPtyNoSAcRH3DLLF/3fgo0wDsa72nOUPlup86lbZtsMH
z55txlvHSqQZysFZPCoEvowSQpMxyZ3o+TI6L6vMuI6thSMAe/7Z+zBiTKx+sZvr
MThAS/F5KUYubRLR+YO/ADo0tLRGH/L8OlgUP53xZ6FegX3ErkgiWI82ip8fjzXO
cWwXBYsAWB8+Xgtgj4OTV6D9BqBXa6HAOKBGWG7guCtbAO+2WFlUX9jlEXYJOdDk
IGaugaJNXhqO5JrvZX8bOTUvY5Mk8+Omi0ax9mPOZFn7EwDJ8qphHAhtrImfEqQq
bUBj2Jlccjr2fMWB4tkw9sAZAAbxqmFrPzKtqg6qsYSbXAPMcuXTg3ruRU2rCfMH
u7o6VuorGAjHT/f7ht8v06asdrA0Gb/Ifv9jbSm6ct4IDCg/qJINpyp4O+DAg6aN
5VmDJH55EZ3I/BhHRgPSzLo7VbrOg/aiJJCZZ0C93bChaYNsCapEzQNfJ8NGkq8C
frOoXRp7O21OpX0N/dkYX+W6aW3BwgijgL860uIoMbVtm3owAs5L1lcO97J2f8Tb
OKHdNjlcvui2n2VgWu1SU33zpkDrlPe969MeRsng/q0mlvQYtGSrRQixn1T0hqUi
P/+tQL8a4e0DbfSxdwKx5/LuE3ytglC0qK6rEEvX/FfOUajx9HDzZ8IED9oRROt1
qit5EDs5nltRP5zzByHS1e/H4vynncfvxOOLMLQZal2raU9wuk7aYreQBvn1FiNc
/6f4o8uXVcZm+DXvt7bVtMgrk7sFqkqPA4CsjdentDK2+2hwI7EbKYWnS+lkVDS8
O6KEPTdIggriqlDm62KQ7q1u9BQ5X5A7x2YaDPX/Q5ZZIJs7CKsrAN2f2cax7P2D
ayii4/14LRkOAHFLhLi949jiU0KmyeyXNoshdIW83bx9WJKk/gXEDl7fTLZpdE5X
S6LcsQ3a6D5HfogwB8PStLesx2BkwxgJ3MJrpeFQxRu1TkExMpmr8UohH81DYeym
tnmUAmBiENSn+S9XTc/60Hd4Vq48PjnVA/znjuPTsUZF2LiM6olv3+Whm1cxQON8
pSKTeo8VAdOBO6JIuohaE47P6Aqsf30oKevoJcHB4KztGLUZwjHRvKNr41RBkehI
ljocm0OmGxdXmmjr7UmNeGsyXGFuouScOdvuJmd10PPQaF1EM/6He2/trabO9Yjz
7GUMq1dF0+uRM1MxsOVWSekQAAZN+qTLvrQcyrSRHp3/q1rFvgTb+JKmYfMgSpDb
2HZSQfND8LytVHJDkVEvHgZbv4TcWR7hlTgugPdTyLlmtpka9PMPQRwgnNzM+Php
8ldQBv1DfiVgq0QOrq+hQAtaHuToNFHkxDv3C/aEVOehBJhjgUkAj34km8loEvHV
3SxxSiryX7isNhknV5u4dGecoMV/VHOAlf8gbM944iJM9h1JqNrLAaxS35IRr0yR
ZMvsT4LjcqIuObRxHHwUOmJEF3z6RfqvXSSzVK30dFnzKrlG+0459TMeuwVeodTw
1mZ7QefsKtaBxUAZ3MQwJFvU9c+UOzYo7SaInYLT6Ce3tdMb9Qcc0E35P63Up13y
sC80TdT4HQE6WVVO4GaJr4EthHLGbMfYEnILPU/5UD+A1oFN2Owqj5msoSEysrP8
jO4thm1/4T4k/o+4kopZuzULVMExiBTWkaTSlguATcmfRx3sxQ8rZeAQUWfD2Wir
tlDeXy45tfqejzXFx+ZK17L05q08yNdXC3CWAgocys7foGpJWahjEqQqyK12D61N
FZZJzbfxjD+L2AbfaqSF13odUNwfF93ZBSzSHqGbFBkPrXr8OACEmyEAs4Vaq8oH
zaHrGzsNw8LpfmFi/wMuTwSMc1qTYiIblUyQbiHT+2LzQYQ2pM8O7dd5TX/eY9mz
yKKSqRbK7SFCp/nv43NgjasCVliyxPQJ9FC0dj++KvCd2cU2PNe6G2ktTWk1lxlz
UpKtyl0wnL7K/uJzfKkiME2PVGUfm+lFh1qHB624hWQ18r/xLs30TYsGvoh2iqN5
p9gAUIUc/Z4VEyfGUhV8iIFXRyyNf2L1sv4hEhO7UPgCKwvs9iCEhD5sDdalDakg
kG4fdH5qsgn3NqFHf5ObAxTCILYJUpfgrvVPhbXxfqP7SgnfcACEbKZl/nxw42hE
W6BHf2IEvEhhutI5u3nSigRjWNRhejtrZ4qyW/dYUYxVE7Rq6X8z5aFgJViab9rC
a7oBdYcy9MQpO9pXoPLz8AQ6P25MIYJrobaNo/pklTPbglYDLKlstcQFRquQ77Ra
gviT9o/xT49WRoGX3+DnryfTHm9jaNfcUO6wiIbO5xX4CaMbNFPTA29oyJxf2+Zi
YbWtsBKZAfRea1UjQAfqYiqGm0flQlwbhKXfciwSr2WCtod21/abhZNX3wZ5sWaF
WR795iD99uPL9W6ZYEpWcZ/sdU5dH+IP/g1uNutYtiOXUhDNMYBpPg+gVbGRD7Ka
vrWD6ILmoahVeBT7NrZXNlmVeFaJslLaQLg229RFvWJGERxHrPHN//7vUDvGM5lk
saDu6nArfrCYTC1EwJNm1B855ZLzSGx8y2PKKlgp3bo+U9kYDDYB2Yn3UOK20est
PF36wzjm5KTOaM4q6gWm47IUXXW0j7mMOfW7XMhZTSpZI9QNfMpzAd+ZwJiTa7j0
1RmnY788LDdm+dzKTztiHVKsmB5tfIq4es0Jp+JgoOJHtTV7pnBPm9GsXonFFc1P
qqaQ6DqWk9ThKqY6kPSGvj7fUOyHeSpQls1WClwDoFBpsCyD47rA9wJrB+T9txJp
ZYgdPEcvkVoqAL+sBOYlSSpBMC/SLBsJpGLt4Hrzd8UzZ8j8TAtZSYOIh75Pp86k
zK0IqgiLTi3Ym5FMCPXnMeCfdN750qZlqPbIqRHTw7uFBDZU8rLqyjmMoyu+vhUh
/JQbU+VJXzRN4a7C3GKI0mjO2BeRnzot4ud9w7UVuRuedk5pW5popts85LZdq+r3
NIU2vWfAFcNYQRihjmGADIVJFOTBHu3GzAUYnY0kyIE0p0fUYF6vBsccjs0LfbK0
qXFJ5snbd8Zie+q6rWyMlEd41WSMZo9T9oqG5S83STVrpdFg80F+KOB445xrrq9v
K/VuCkvM/2MfMdUC0sdnTQ/NzFO9z2rii/ExRp3um4uiFxvbUKEhSA9wqI7ZiY7h
5cYOO6XhYuJFFFjnxsxzTp2tBgKoN9OW/t6lygUun9o/ljTlfUSZhyYC7nsuew4k
bzh7r3J+a13Mdx6L0XlxVOJ4pJoE3OUjIHBUYxS2nrMTbHywo+/EBB/KhtBim/e/
Mo85A7OWiatC/QD3GxR5wCTxi8G/8sLznOtmnYZplfuyevzFqHGr1CmqRdsRPDVO
hb//+N4K9MpazIm87tJKCQljV8z5cEykwm9LINTfKgi32zTXljDkxLdhtiBl5bnp
W+Y3CT/QCdZBypS0KKx2o/pugWeAZN7JeFDVvncnkhKerBKxZ6bHkw/h1TTwcYdF
50UxD9R/dW4hYwYpU7CIuU7p/uJw8QJvrHcChGxs+lnAGfVurz2/6UGTYXy1Gc7r
K/ihbRqd2yE77WWf5mRTktMI8FSn1AKxs5b0k7j3FiZ6vICJG14IIC8ihg0xZWKr
xDTor1QbmuQnXMCcwhKHzplz+hpmhD7iNToJCfn1iq4LAXnEQ5ghhmzXfvmAZZWQ
qmhsYeBqobRE/6xb0wQSikWFqlwN60uDrXnPauKTb3fd55MxLK38bDoHLRGwKKiN
YqCUIY5o4EGIIKe13xL6X7PanyJ4xyyMChS3xVFEKXOYxbsBwov+rzhdvyhpSFHX
MLPC4215Tzx+d8F9mv/EsPAVhPm0A9CUCwoBPK+QwVqeRYL8Yo8jd/1E7GbURKk1
3IH3m8uso2TnzeEA1hsxy4yejRwPwPMLaPe3sRX7pkEdjV5pdblUXFDNgoRgvvyY
JJC9CJLVDyrnPGO3guMaNh8SMxQtGTh/tR796z9vBf7FTgRHSzoPk2Yctz4wwmCR
hHvl/+KXqpsoPJ82IKfXrU5h5N7nGoroWcMknwhbRRLWuxVwan6kh6XylcUWc3My
G2uQf8cfAMojdg87XoXG/fmUcRWtosKScrXeR2VEQ92bc4yKNV8frgzjMXkkvP+l
RP16bXX6+NjebuMUWu/MAA6vtHlAvsWrag6Gmf4Nbyq3t8p/opl6LXiJ+D2LpugT
NVeLajORlfyY3IJ7sf8l2s+/870t24YIIaw88ZDzRjKAyivELGPi5o/fMNz1c/NL
cKbOhBguv4w8nxSR7jRDO2WlyXxmgoDjHTM/xM67tjpeXUKzmHS+GFHPOaWKTy4W
jXvU4CGE5HyKs5SL9s5+ADPsgzCbWVa3rdjM6wIwhBFLOu9BWTgEA+gMq4ssmymK
K9DMH/T/kUukz3LjzSNFSxHBt+UNhlyf2nrdIDjJ8tjOlNtZREh6prfNfqKsdGIH
jko8nrAddvPo7RO1b85YTUpk7TpUtFugrYQm64mQboPPH3+67kuZlQ/fqhKbir3o
53XeI3KrCT0aaAdesx19e0rGrFbKVXDeXBpwS3HCjt4Uqta836r7AWCM4aB5lxvf
TVFLJmL7aXrpU5Hb9fXVGUNNfrEJ/PHK/OMpq49fN8lZKk0ANwBzN80MjkrqBgh6
oezlslfDNgMtsvzdrRZsZn1OphAKB0b8GUH0uRASomdLI27kCZL9mmuYhIxIDIRc
0xFjnaMpp3w1p7AM8X+osDRg1cgy2arfHkeFfW81ahK5TCzT4L+WMHmcgtJTQHQ/
WI4Z5OmgHPR53/alMqRqFllaeQMboYC6u9zvF+mquU5Zxe0pWRfPtiG8ezxcZ3jn
9g7/eU0S/ejWAk/6fzS34PaXGkrty697Gjx8NFOpFOkiQCaw+/43TVe5cCuwl5XC
Qhiof8/HS7Mw8C1sqMoGU1gm0iXWMeufJGmmyIlsBrXbuRle+MCmlB6brwmbOekC
N0kJclicNtde/FKhSnbFGZvg24mxpWF97KaQfgIypyyp+3Wd2x/RO7qLyUlB1k9s
ha7S/z0j1EysMnklibvNre9fZNHEBock0k6/Wx/Q9wnOCYkKLSoGS07nRkmwk9EM
Fl3hRO94YAsc9YnHo9le5AHmReJ7TPsiTHOJ2/9jW2OWxb0vUBvW8d7piW3pIjO4
aE0/K8nwlP8PtrT2mFJyFJKQ5cedzk8MCWq9IedIESEZmvSFfZnCxVVfPhHBgV/F
l/n/T+zpGdW4WlqWwshdlLyVxgKkrHVc6NQaJLtWEf67xSX9hBwoiPxojTdASQ+Z
TiCr0fP2P/iLvCoAF9XnUzVy9u7kTGJap8IX5F/ScKjZgf8H2E2UAq9lirZRxHv4
I0rWP5O0dF8Y599t3I8H3mK7WkTJJAY0aoNwDRrDoKua+2iZO1H8KmuwXB849gpb
uTwnz0GFpE/uhOxqPHegER747/R54+/VCcSn2+gW27j+0OnEkeWjBGbhm4U5aHAQ
z0yft+8dIgWbk4NwdxdA5sk2kxM1LbhTcd+18TddFXXT0WMwd/EdLohi+U78R2lm
mHZU0gLV7+bCkTs7MaOR91sVYDh2tXwjdwF8fNvkSlEuQtV2SwC8BbP0mFGd9AAD
C2iG47SgfrwZS4Mn40xnzgx9+ORC1Wyfkuslknk7qh+nZ/BeJwN1xgb7NqHtIEu3
GU7LKCQsjINrpA9yus6R7ulmQMyhDSLb5rK8eWxFK2uOWxmotWNp6inwBCBJ6jVD
GwpL5c8GJoe44ZIIi1ctqb+lcWm/pmiaJaZv3ScIR2PyPO3fdbUemBY/FadNfNj+
/E5Ac9dNxOpGfpiunEeX1pgD/7k8Nvess3skPMzZtgPaclcds6/uq+v/GRwG5+Wt
GQMGDKgSPlCGy2bQ/0jZbSRLnaUwlJC59EB/+DPwH/rk52Tl/yu/sHZHrBcbtd96
wFhee/CiXOOjmToK9/mYE2oRXBeISGcLiBYySQXhAr2m8ZczwenG+C2GKR3wE1GN
h9oXFe/OuCBxYyHDuuVlDBckHBa4mF09T6o2JCeOnM/VJdgQsfWa9gGcOsoUdFYf
g21vdtSvz0bxIdsyzqL9mK7OY/azdWJMToVtxTgereZGAoya6elt/87i8C6+ewpb
S93Ns4Gwj+Re5zT0EraMuzDNbSAgob+xf7/OD8Wav/xZBsP3MofDmE8TzQz50OKO
9Pno3CrjriZSjkgfPzTqPi7iJOn4Tg6aIpdv6DrirOEkCFcoNDcd/bNYTJMFCEDH
mgJYg6/Bq3Fb3MOGHXZVt9Q5VajYt/cDkr7WPVGOci/R/6Esbi0XGHqHpSoI0dap
EEkm1x801Na6z0hoDOzfr8mbCalvU35WFGa2DM86gm9kTo4UbtniPdv/D+UpAb8M
GhKqZnxbhcb0hWSpuJdZVUU/DHg8YFG8QXWJ6EkioPmyXJ7jJ1jFCPPckNDFRI0T
EfxGvvynrndzorHnmfvzRzPqPJRkc0zb0ybJjwFDY0wsDFQxA937qaGliNRM5VL+
17Movi3He8ntyeqdGsAlOVen2UEfClVkqrQ8cab/rcj/nx5pUU69I4tCUppxX24L
TC9i8d2rACruTiCpWg3MWNEFnBwOqP/3dP/pfkegfqLpvMtlpOQtdFBI1NNPjaId
odsj2LVKs5ctHr8RsrbyuCyCeUP8URXixq+BdB7OVZQ8nQaJPVIqFHol4KmCi8yc
/t/hhyokKVP7BVuUAQAwEP+80YRon0Z3g4owsYQefhxz3KJ7ky9pt/zc6C7mbtT0
lq6gJm1rF/urGy9XaFwFM6yhftq0VoZ5fnRUQ4Lsb4BxQF9GYoaEiPf4fBf1vk95
SGUbAqXgI7JKEbK88DsasGWQEs8r2ctxpqK0TuPZPqar0D86fIZfznIoGRML/LMj
9K5rv4C+2p42AMrieTaO2HYJiDwKXI+scRBLskiF/Yb0XE6TCmrP4AudvQijOQv3
/AIjtMFB7cXtqF7YMG7OgVI/Fbijxge4qtiUQacIpllafVVJsOGwOxbF68CDb/Qm
ehtCnYBviOCvzk05VRE8bBy+zSO9DQqs6m+pipS3eL3ddxNMG9fP0VJFHWCxOH1a
R3b6b7FNe+FZ5EECXGXMN4OW9s0PjibxGj4AB6jEDWeY87MvlVyDbGnWtnIvcQ1g
aK189VHU4EZ7OhLgHYO6lvvQhlnqqjwhLLaYj0XLLXjOMK6s0O5dCkdKRtZfixcs
OcXeCAvipt4UBKBJn9030WYgDMo46Z2iTykVc9uFrAF+sqsmscKV2ZD6siYB1BaN
BU6GXJsabzP93mbEfmlyvewg8AmAekYK9+pvFLuYF3kuFBXp5+TbIA6K6RobB4I8
DR7DbkKls+n8u9Hf0LqL1Yirk4ijXEbrV2MJZnwkA/qNtzbx7FvzTfEHcjLYIWDs
ySNVxWM0sDyR+DH4iFNL75wdqwFyz/cj25qID2x7kKacl+Vz4csOFBTpmoWztTO6
Vi8tXM8HEkVGynBCPcqGRxjJ8tqfpl5IcerWG/wiD3waRIGvpwi8YHwUCyx+Cf/B
T+R0rz5HCnkmHGxiVaSB/GWSUGQFom7BBvi9wk1EM0AOdGmyseR2Q2miO8+qlRzn
p7eYDpjzRUQjuEcseZJ3rnjCF/8ra/avjtbKe5Tpn4Qm2omkSIT9JL+VuQIyLudk
tNahmkBLrupFBTJD8wPR0m75Xn9n63Xza/Y8Ns9DcSJcpSN8uZPWqzCYpxlj1L4F
0ViTRt2unAnSfX6qjJWSmIG5TFNKsQZ3EHah3j2TSx8Xn7Kw147M5FOPRdpGR8wJ
q9DQXAtjmdFaCLbi5cRXIqXtOw2WlXf2/Peo/2liNPULgCa2qG5U9U8e50uy+8lL
hhkg+/5B1pgGWxJVdp+lp4uTKK/H/RchPJtqVRX1t7hPr6xnaWxKEZfh5NdacifQ
GtC//hrMbLFe8UFPiTj9a6Gmu3x8m3O4KMCpdmSnCHYZrv0gWwRi8rKDI66PRxgW
Cufr5E2F8HU85mw82/Z2qEHBxfTzIJYXDGtQ/BpxR0KT95TNczlkcZxRbQmfAry+
/c61tuJikvgOSkKhLXQTb7vaRxmNUeSQyUBVVeQsGxoDbBi9DbWs3BTbsnGvNkxm
7exkwTCcTRr8XSnKG6wc9TapOzCg+rHYpUnqdNxfEOJK3M1PJz7bINYOL9xH0+rI
l3SpyVP4eJlaN5D6lmWvA/qer1/lxi2CZD5ARZr5eOu+wcgw/jnoI1mqXt3dyple
WsN8kOQjxlHhWv3gKUL0vV1S7el1i7OsHG3kxcp/eCX19hpQ0naMRxAg/+bOc2po
FU1A18kOkPKxDTmyotMMOEaFgKSDt3atX5025dXnYyhXq7wcM506P9n3Gh85GMzE
Z4CmaARajbovz2KL8FKqxv5+2EPA3crYnk95ZVYUl9+vLOZbzHT433xhswLf3cHi
lQYQUYC1fVBZLDdmLhIM2BWqBPOnSLK4Mi090DeZ4RuZ2WOWo/AmFeAflf2Th/Gz
TvFHMoow4h32/a9bcjO9t0YSgusoL59X1wmNv3vHO8HFB9tMOK7jvNvRvVdDQDGH
iLQLbifCMcEhJRT0A8Zx/t4v79sipS/XDPbjB0PJjrQpJ/c5lxmY6qLfC/u+j5z8
9EE1KoJXp9gxyTN3N1aWa6tQVKCEdQTbNVxvVgwGlUhsXPJnBghPPQux4g42IaSz
SIFkKVyLMH3a25YdSRcKjxBzqJA6WzxO0y0PsKUDpVL0qlM5YK1IUw8AbbeJnsCZ
XVIXCvpOqFGjEeK4HHCU0NSxHlv79HvZd15yfddysvhr+CZkwL0WzM3GEHz7Vz13
/97Pake9vr2bmbH+eqbKIoSwxkSr3uqh1O/Qc6rIrF+spl7hiVj/v18m6tYFb/6L
EjPE9hDH4lfpItqB01TR6jojd3Jk+ZM72Pwm3QDIYp9ASEov6nl4HA+wTPMOit/k
g+glKllvEnsjy+XNxKcmiUbsNsY12uab6inNd9L3mxarBCEN0NB/ud8b5VPYbIEn
2S78QfdGELUSLbT4uXKf/+DNowI/rbrnHu5Kb8JL0AuRHwJVNLG4O1/CUlb3MdKu
xkIgMEJglAL36Xn2vnMoeFuW49AWs07R5GfZGXke1N2pAk/IT+81S0wLPvEQTmIB
gPd+HO9gPY+q4vTDa9bfy8Bw5D0dVX7djzHaR3ztqubUnAvLClw0gUUPT0vvEyn1
/PLps/xmYH9ZNu6wcnGKtlRmijoFe6knXZboP8ZNjE4l3xgRIgQMGO7iCsjJWIIs
vfMkm1ZY9fS1rLSQKpHXysjCRA/V9kr6kkKijLpK78hodtr/kmluxoquZxbDHx1O
FJw6SnVgd++C5/I2QnWm9ahS/U6kWiTS+KpzfHudU+8iCWNepKeGrTKUps4HkyYg
WOJGfe+d5QwfWdkxUTd6Qca1+6tihgBRmxGK2GphrfqGG19IYaoC1gSy3Z7OCTrk
EBK37X3rlvbuCPOa0ew/xdH3qQLYKHOlpNgmDug4ZZ/AXmsJFcRn4IC75Vn8HJ5v
wu9v5d0YnmiqC33DovhEdWAFUfWQD2pxRIAemroUs0wWd+cFLFgsKCzf2SepBRQz
ri546XWRdO0pDkXR5n4yaVEUkXvH/lesmqb6V513Kv52o3JLjGHpHBJlhjlJSjt1
/g2QesVch5QVdeNzgz1RgQCwbUbTTsYKkNiR5iEH9Ycecsz9DbVin/2Lsrf980Qn
kCKdPD5HpUZHGXVx9JRqXIHZWZTwlk6428HXrgnHi4CsWg5dx6H3h3jMQM3fE8qW
VUCvIs4JurL3r04ujqVzCFL1sCFIP2IfUTCXd01/0WO6nURSrxGe2j/v4SgTfSQQ
nOKyiBx/MW4AuETBzKGw0TNw77f4YCfsfWJf5cLqBaU+qgvW6HZWQD51bwlZAX8T
HVqOAztf7aKrXL1ZTFbXwyrngVZC6hrLQSpObwRYg1ABpo63B0AyuWi6leSNvTrq
XAoJU3mFo359WI5cMoOcxHhsE6FZDM/xf2aONnG1m7cjElPQTWW2eOl+V9pznFcL
Op/zjWwmvKEhibRYgMpyew+VeJtV24FnkmkpB7iXBqsDb8vcb1fwpV39kq6QPVoV
XvzC15BefgG+fVGTywXFrFhxRBaBxjTYUQDD6HlNTRjiDseMK7uAgL71tY378zTT
Ri1B4P5Cy6pV4ZmCMv2WgFe4qsWrsRO/agO9iPvlvi8kfIkPjUJzCXnnX1GKL5zs
zPew64hgCg2IcHYTM6yBIDwWFlvJDffnMuQ0u4dkZyUhW93hvW3UdgfpnlV1mwN7
DNKfo/kSHykQdvqcJw7aei+OkarrvxQfSdJU9IAt1hfU+DSsk7gYdCp2vbrMG3W3
sJcKeYwP+m5Ogk0ycxeO0C7QSxWvO0zu9i3+i+yinwTuhCBXazyZUoCUYPQUjChI
rpL95x2MUr1ECz5Z9jV/oYnLw6iOWGqRtanAoOaCKOR+4AuDxtVmCguzfrHNneKg
+povofAUf4xj6cNw/rzh2y0WYw6Fn0ZLtZ2uLLAQSbaELWpHDjqNKhq/9O0M+mRi
HXSwS0mzLDGuD9yd580n6VgsFBcwOlhBmQ3llO8XuXUIYVAgVV9nlQq1vCtKSc4/
Fy+HO+oh/n2RJTzWXsL3Ha/3MNxSl7fqyXH7HZC4fLTOZh0N3PFARo/oaI2R/tCe
rE2F8p2upurTu8lOFrBtG0wYzEwU6cLyEyx6neyGxrvOokgrIQYbW8kDmmBnMhWg
mm1OvgTyUM9tYaunevcbwxer8MIiT6Ok8j75aqG83RrR9XRZQW3kkAh/SF8Dk4bX
6qfP2HZPXHJlboXzxKmZFrqvkXj6ZFVkLRfQy3PC6ik3SGRlYfoQSnpjOm4ozsfa
UkDwpXvmDVK6ZL1SXSZazBWq0mfK4AP77745jVuVRgP2VVefTQecaKacGAQkW9gI
KBMJRjyVJE6ux5sXgqhmAJkdRSr43lEj/bpLLS3msir+soXm1/sPHLPVeNZMzJMF
r3tUo6O98cdsud8NyCwDwd4iPIUjojbn/SIp/cFHq2XCtUkmlB8NLHRAJtgnaQ2o
DSYQ34U2Rzbl2GfOUbuwVHhGcKnReriXw33pWZ0TlBlpzawAeHhKTrgMa/jA6nA5
+0l/8pJYq4UHCE0c1BzUq9yCiSc2pgZdJGq6TZigAQSG1AuOgP8u9fKrd6gBlstA
VlrSUASC/cs5D8gTq39C/v2RH+1n2qAp/teUkmceqjAB9Zzgf/qAhjgyex2ENMuw
ivkTnidBZvbsZD2Imv1DLgPehDxsfLXTt62iKjI5CH9hYvPNUhA3Kyl+0rSGf/k/
SGuWSiO09fdqC8uuAeAK0x6FVtD5cLzS9UN+vX/KwXFmpYR+DAHdgXXaf8dqBxtB
utrFDtuMAZtLM+mjYcpmG2W5mE5Wj4E0cAfn4dFtQc30ZlFYq5F4v43rwEZProst
gTXvq2xBNwuL4oOeWEe5WasyR1Y0GkW4dY7Nj78CwFDQYfoDLQQFZlBx/P0qKZAx
jz3CzjgTZCLTMbcjQ41ZOJj+s7gQevUeNCSttI+hPZGwkE+gUMbIFyT2pSRha088
5jqO/1BaEfVzu2onthnuarIjdwkTQlAdrz0cRNaREEzEI9FLVHVEbZbncp96NuB9
XTsUqQDq77gxaxOi/zBL4oNixj63SXjC9REKtuI38zFYlvLprKp+7yRSahbJ40rk
JHOG4HvKu01HJDwjOtnC9ktJnYC5n2L2F4te8fqjN3LKPWxWQx+FHxntaBz8qhb1
Qj14PnCtWyZ9wuUaX7JRH2Y8GNyaIeNBV8nAlUm3yT30NKVYjw8seO6W0R35PjjB
YKJPiIFryFL0j5lNV0pu130xxERb06vaONic7rcVikiX9fDtrJ5yP69ywWOjHz3u
myn54E+uHmc+gUs/qUExmY4XYsZOs0KcYRhoDsuG7hQ70N43mVntCsRhLz5wcqWu
ZwILZijEO7D99k+NeYoorEvQzRJx44EdImD9Lsbo1eaSRxUnnbQK2/8q2NdqnZGc
L8gQhCCukSyNQxGbRWr9UYQ6/ZoPu8w9OsmhCBXL1EUkL4MIGBWGs3TiznmmxiGc
XpDZQqynWabtTuwCN7l5P6WoBnxLBS76nauM1H5LZjpZWBFmnLJhTy4oXVLm5QEP
0griUDbxHsbniAGPaZQws3Eyh4PzCDkhkJyq+AdWZaIAeP9aOmS+6TQ8CtQgCJSn
wJty/WsP5cTtsph/7VPSl6CMYWWC0yJNHtNdmbEbt6UyMhe1dENNEgolxMrnrdUk
d/7vNORaiXL3/FMUGG6Pter0FfT9EkCFR4FUV2OWOJlfqLEepMMLmrGRE1qjzfRn
xebWavvRoTg/uMxfCJxjirCXGb66S0AfMwIvjdkPhjdHt9YraVT8gTj5vb2SEh1L
1bl8EGk8tiJoh8ZwI4dTp+bYDcsfGqBM6t6RGNKsEbpAqD1e7pkVvVBcBhxX+CFN
mil5WaC6p+Ii06qs/Pok1Svs2ajACGwJ7yA61NYQiUPhy60eop6IFcf+ldN+ugnO
r4ebykNpxgfKebdcug8I9bAAIGTGOOCgpKteWR9ILtHSh4qzwgafL+bIgDPAOZAD
w1S7IgpEPFHy5dRytTH2JRLPv3cnl/v5eUandRU5B9Nm2Di2oo5b9GP163x85AuN
3OKx+8Er1oeZljMueBM/phPvpo3yaTeZ8cBqGcLVn6GR5FmnhsG6aAeLKm0o+9WP
x8WmLVhpYGVAR4QKLQVpw0/y0BT3nbJZPyYErUdhRkfVlXnd5jhm5NO41wnuPxhX
wQNkM2+5cOCDAKVhohyE18dm/EhKbPfqO2rkgMgK0nEJqgp8A8QV7Kk/2E5hvcnI
faukteAg6I+ipUcuMs7QxVon9YUD7R2xQb1mttOSP+RMmcxwh4or3b84lAmg+JBW
SnoDhKK4fnkRKN0kX+7udcAqE8wapH1b1rXfBatJExU4RkjvIDC7DBKL4Q5LvL9X
oe7Tg1BsdEb5vCUYYoxTdgvFgPkBtYPXhHyGaLXAHZl7JHuJvMNlXgNrKfDvd4gg
QVEXEp3paAXfvakB/rItFBSE5n2RbS+h87xgcC0VQ2I2cKC4/CPsQL+Jrswap6Vx
RMlzk9RlNiu8cnFTGVNp+PZKMLIUFfDZIN6pkjsdYw8lIxpxJ9eQiXA82NUwB386
KhlvV6ld7HTwTDSmz9XCJd9oGJYubVPsXTOYk5cyHaP3xPHRsHcAbjj2cyEz+7rD
49Y0vo4rn8vrkh1qi9aiPjJ8e6uAMeo1hrGPyhbMuwNSdyO2O5OJ89Zm1oZhbjCW
luSJM3a6p8ZmtLB981zRADtO22hJPRPV3F+5rfaeMjXEPl4dawK7taRCRcJRac2f
5Wkh7rF3K0/gck+hl2NThgph5QtV4YY4gCJCIIxvmOvmnV2eAVElPrzmXhW+RZ5/
/VoZF4Zbb84/o1E1ZwXjg55XrWaA0nXXAqAuBJtEvHpu31kZ58dsYMTEKP74A8Q/
yQ6klmaEE25olRROX+pXIWbJeIzA4dBVzUdfec8kftefrm++Jrw+n2bcpr5t3YFc
jSqp+yFgp90tzOZEDYq1uiJ4iPJHrkDWBn++l1SRRpsgw4ER4pbwHOYKzxsQ4mfq
NTXgaNFwJOo6LvVng+2ylf5eZekGCt3LOBOvdsCjSEyqBRl+x3FxeNBectcDvjHt
2yW/b4XoatgPqUaWGr+46TUgYzNrfqvkIovuCZHziKAMgy1dWWnJzgvH8oSM9jh/
Tfn02I3f5vUZKJeN2Ibu81IMkB6+zQr6vfJ8ktnSvcDkMoBvx4xq+F9Za0WM1oiZ
vK9mdFhjDbSYlZMLhOBe02fBrcOCGHLNrApnEf30b1rnfMhx95b/iHn1lT2PMBht
y+7ky76e8WMC8w9518Mx2ZBrngOcwua1QkqdvjquqOlGSLrdNMpR7IMZHzO7WKKL
HvnHCkjJ/H6XXfPfBfhNIx7BwERPROhIskGQj1LhJsaiOh4XWZm/5mxQalkRDZ2w
/a6qZa4G9Q0rg1VM4hNhlEiubDcg816/bKiRzI5U4Nt7+ADy1cbP/TDEM+TCSnqn
uDE8YAk6mdcLLdDjQw/aAr/e+TNwEIAqVnD5KQKvdg/HY5PPOwo1DH3uMnyoKVn7
uFR9ZjAynJvRM9pR1Ncufmb8h3J+Q5zqqeTv+hjIjikalEmbMA7dVkcmHWLJZjkU
zD2OqKWTBaVK13wZDDL4YofmhVo5IT9UgB/YOkoUtjJigNTWrUKDBR6ZyYJnQf98
hyZpnkie9yk3qNNfOO85Y63ph4lf7KkpdpXU6HXbrreSTXKm27xQhmgXD5b9Ng+B
s2U1nhheumxf3GY7t2u1GvTuQgWPsaGUU2l4h9douELWvQ0A2ilRnfw+8XuQQBhc
BpWuUT369FZJu1nxbZDj2tag5H+QAguBuhlCdX3spSTqgKbVnoS3MaA2p8F7nJtQ
QJkoXqH1nFCr5nrVl3OyDkggwWX3rZfmLUpwRiEewcrDkmKZHl00obAg4SfK700M
0kNZ8aTpIQs2zRWir3lGK9NBI0JY4rnW3LHzoJ/xPeijIqsQ7GElU2XQYRFEzj98
XUsxWy+BVkOR3FTwxW1GytvIBXURIaUH/feEAa1l36dVGa0n3UhslOfvuPC+dpSn
kLAmGX7DN2Cmsup2iniqibI8RUmMBjFOoFXkbsnC/eKe1MskXEwwQ4vNUIrB58jo
eamlVKNr0+dxkV7E+BeZLhytE0TrKZb4BDBSx718r9kqJLIKyInnZOmjAsmP2S/C
rjiB4chtMWkS9QC+RgkRQcmPAZhWdDz6HsLjAbvEmB9gJy8h7y58F+oP8RwUi9JX
xk/HFcvnhyiIS9T03Q5l4fIBr0vtUq2C+XvouDjn3D7L6pzahlO4F7wrysKciWkG
B0jqpGcip4BkjHgEiCWsdeJDYZZfWL31A2MS5/0tZPvueXhCDrY4dEGnv491/9C0
8cFTQLLhBFYI9tbZWySI0PV6ecivs79njOyxB7bIOUeztwsivguyNGmqk1Y7Jbpc
uRe0Z1JmDRcuuMuhtfSyHdXezvnIUAtE4F7EOVANtivhR0s3923nU/6F2IJdjByT
u7GyXtQ2zMiECNWV4CFwCun/mlUMU96uVLfqQfpiyjrgP9Cx/6PRgJj3kA4MR72y
sSaYFVLvZ3TjhVSrIZ0iy3IhFvTwICSKY2AzaVF33BVX4+vCr0NXZyK2DdD8XWiD
xP9mgBEhnjlib2yaLm9hBJbcxzmf2PT4xyruHuVKNBXhMNamW4wm9/UTzQgBhae7
tQFW3XaZCwOXXkj3iffHyVIB8tUAfMxMO+SBpL4yXPHQv9YHkEIppnYx6bfNVQkX
CuzzAf2brad6XQZW57ArpW7TEJZYo/vXQAFxC1VuN0JELIW0XG1Ks9reU/yEHldw
xJTDYvWxmRz65lEn4scMTTRnA1S+fvot86wqgItBsUWT66puQDMHCCb6g37qQmWx
ozCM/MTfu6so8aYRtaByjrN/ZetfbEyoy6epz9OJfXqePkuom9EveoCejeyqmFau
UdMha9RpEKexx+BR5EqDCE6Zbfkg6QOWqmYqF6OR1HSNUqcLoDWLYJ66glo8p2Qh
0h45BB1V48PXrbfO19H6BCHRYyJAxH/lNP1l+FDUQemsDaxGFjIWQcjYu6bTYzgm
YyyjU5sI3GViBrw8zcLf0t2BkRTdnm9/o2Ip+G70ONVocqNoBUpmmvpihfXwRKyC
7TmYXC/KdqRVBEH9XPOS4Mw4Ne/3JoS3g0jEv88K21RxA1G97yf926aaJQSQdyoJ
0gm1t6mTxBUc6Xpi/UefOLQ7MKKnjsIJXXDJ0PnicvMgJAQo92Cskj1rxaFyY6sZ
Bz+NMcR0OlhpPZrXVbCxhShahOjnfNpUpfBNPwxP/65WZ4Owkz/+Fe98L4kLWkQG
ZYQa20ks8HFqlAfZkM7enk/QHYofJWVdMS4wfQ1S+rSuvame83Pk6i9UhCl5XVUT
ZCI7Z8FLDQ8kIDQZv68mpiBmXPesjBVSbxKxEhViPc+JZDTQJcDEd5KVSezqKZN5
IPOjEwIzgB3j6otvt1UW30buEEZa+xOLNs/U0Gk5ue+EZKeMuYaeEA9O6oq41PTb
8h0UmOj2BcTMv8H0gMHsjrbRB84nKz2W3K18oURiG49vNiLfo0hdriowWVC9MfIB
5gZPcsjFuCU9PWYPRscLwhtUmXNYKSgjZg9beEjtTNUX4rwbhIvHeD7OnetNhmox
JuqSmLJAPShbmSkevXZekGEiPDPt1eE/Pr9qnuzPIYkkkzWqKd+x5bMN8RACvnE1
n0tg8h8mK7IfZ1qu8ikJG2I5uxkZbd4twFtPgCkf6Wpi8/+jrGd5a3BF05OJiRk1
3cCPLf0qxv9pNO0EPmnMGnFVlvcuVyKQDBFvAR00ptbH6aBIOTNZ8DDIKKvAmJST
yjipvhhETxs/RNfuu/kdxk2JxOEY0bHkx2+mkP97e8gfD/3beqMR5KIPV3FM3G9L
hO8EjTM6EpLb5tq5K1st5ZjwMpghhdW+/9fBEGCRvd1HOaf4iQiIlt+4pOAsjPDG
cGYDeINJb2qfSlSC347efgJVoPex9STxB7LBiUMOXgsUUqhj65d+mckT2z/qv8sb
dhLAMwtklK4P53gNaAqvHMDa7QioJZpcxhhYzHUAi0Vt4lm7n1Efi89Xdei3Nvg0
9ePk7VKj5qRtXeUofo0ggxYhOJK4Bby90qFaOEQSTixJRIJXH4uyt7egjBAbkENM
a5K2qK13P4YylH0Q2ESsywUBLaE6iK0OahMJWLiJcPRVUu3280jFMsVDSmhWMpOl
Ka8frBGt0cuU+E7CsdwRRRr4LEJrfrdn2jrGGGdf+JtdkciukL42KitSFuE+FNYB
3FnRbxWDGqkTFtrtmh9DG6UO1Xvl7lCBZA9b9I/3I2WeQei7Wa7aD9Ivtp+xwyJE
KC4vgkk/BQ6NCDvUsq0r3p/XOw+FjANI7VgRDsNscxxyt9LfgiPOwiR1xZnIdDEQ
y2dLdcm7VYMhpTVPd0Ox4xN0y+O5NdSYR3I3yb1L8sYdMJ80YGeHO2GoNkEcpf/G
tKC0tOuhC27fZsfDJL6sBPVSXRshW0s+EWVmmEuHfH4iWEPVqFjmstniUls9R8nu
U3XbQciIndzI6nDGRre0tyXGPV3Z0pfniNLkl0Fls6HC5dNslpV+U/AN/jHb52AW
n1N5gxPFKnglnzZU6uga+gFJkznQsCI375fXDUBtPVOS1n8YdFVhQy1SHosZkDBr
VSfM3npnsoIOOBx4qC3aag8ih6PuFue3ZSNjEd800ILSTy0dYVZidI0OXoFIbU5T
eGSngaTmxloVZLerlGfZGaOSrO1GV7ol9aCnPLrHNI4lGZLHZT9raFnCbwl9KlOo
HfI45QUsFgjSYSPdgL1Nff2fnrs0imy3UkXiZ9rPYuYYEph9PHf+AT/sRUcdFJhA
Rwe8QA5kZ5LP64ujCUwQ03Dyq7ui/Ky6uO9fWgDmCugxj0BtnjSc/rYc+Fj+dtJw
5rv5hX8fidUsjpNsYDJFLHnUBD3Qr0mueT1noCDmIY897R5tc3dHOC7BIuEHY6/l
FoFID8O59J3mCNA7h5KPJ8e/97P7uPrdqUFvpfEYFY6K0+If3+TEm930J+1HLWf0
bNhQkV/4onnmn3VYxOfVn0qij6ZZUzbcdgRwtmQ9ZTPhKmFPlC8vNzeEr0RTIfRd
BJJZVhNhXq+JSb6xn0tf0WDNsbyrnfWQmgFTkXMUKMjcXt0hbhEfX2Pn6NEt+9M1
FeXpH+VN/OcZ4yo7QNeUln67/qjKOExCzMCFlBsE4zLq/PozxPkY97Ed1bC7Oa+0
Zqyn3qYr1u6f5TsnZxvQy24U832ZlMD7cfLsVK2pOjF0vd0nrZ2TZ+JjjvP0a0YT
SKQJXTtJ0iKJzAxd3afupqPK01s02uCvnOaR8PXD6b6V2JPbYMWLpENKLlFHgFR+
9rLyIfAhXPIAIkph8IDJYwsT/XZ/56HU6e68r2S3B6kHQpb9+awteuBRMJZHA47Z
66lyeRdl5Jsag6obebTSNH8nUAwiukD78slWWZ3wQ2OJdeTakzIK4H6FuvZIYtCJ
sj5eNNB/VDg8O6iKdO7ma8ihoKh95etbnykDscnSMXLHO6y/kX7Ocyx0/2/UlDEN
vmROW2q4442T1BxhrMOtOQQ1j28X+YQTlDzK+B++CNPtheuXBmjAzOV3bhkhSudd
Fx8CAsc+FFE4NXWJ+Pib2/p+iS7CyHQndkeYXAM9lpmNSDCW+xmIsg5tlmIzvZnH
9E63FwfPtMnnATrWn/B280HyYjni+DFbht/oZfH7yA/UBLlNnYPr67JGSp8tkgMN
2s94qJA8PyBQox14Ry+807z1nqQhbB2xxso6GDeokhP6NQKO3M4cHZ020MRKNy9W
6oUOLfFJXMfN34sc+LOb24jgwoVgf4WPtYsb0gIzf7A5UgVMs2up1hz/+M2hI6YF
L6S/lHnSLTRr6YRC/pb62vm3LxX1UzFPrw1bmHFEXMCjPZe5U77mAwbGkYbrqlIl
zQ/F4gA+JmNrgCDX1M3OvhgzO5S6le4uvjYLDAPztc3btNK3S4ioo6h5UoDRyykD
fNwF3jGJ2dcg237H7pb9sBQilW7eUcBNGVH8O9bXUNV9OgVT5/7zBSVVDWxe4HQa
rpzGva9CgMn4IGG2FdObz2Meq/ugdukZvdo++nBgx6i1JjUaiyYRreTWiv2qvHcZ
O+rpMj2hroj4anIqwPdpDi8jCi7oAB8u0ldOW6NWeSzszbSKF3cFxzBomoLcCX89
uScP96h+wkhQKx9q1+yTGmq+BEpCltVIVaE1Qq1KnQTnTkMuYUjGK5z+uBrtjDBK
R4Uc7CgW1scB0kRCDLcEZyHt7tGWzR3d7kZNHLUixfLRt4c9RBpFdFX109SEZu0q
LicDCyDKx0wRwaSW4GK8fxRmoWcGFQNCsyK0YnoeKhxYAWoNl0I+AHmmqG+E5LEy
rJmB6BD8STkfBVfaIwsY7bUSH5aQ/PgOhQq1LelDoIpUAStKZGRhzFH9grUg4dDk
Ojhdqe2JmJ9u2ChLJotvgbWNrB1IpubfXetIJwi7WSvqEi0QKXa3zkovAbH2Uub1
jfjuOXNrrk5ACFj+pw4ilhNh9R8kmthVELm8qE1AhcJkJOQycqC2afY/FdC2Cnbi
VSJv09MjRnxJRRt+xNInonjTzIcNMvuYN11ja7byuxug4eMQ1vyEGxb3FUd3vZbv
dQgeewjxuMN1dJbfgbcvpPLoy/OvihwKRMafWbYWEWtIMlowXzzokL/EZY9xKDeI
G1H9x1IoL//VhQRvW0y1Qj8Zmny4ZxBOYrbYlpy/3wc6nR5qd2DZvfPJZEKfcQC7
k2a1Hb22pocrKft6Zk/7DvQZsg4nO+ING3SrgOQC1lW+qjJwf16Y7dfKPnuJ4pFN
s2SX2HK8zJsVpdwZyKr6LGiijDMijoYc87vyTyYgsImnS3VNhFHLro0UYC6MsJka
gaFFa2aBk/LzGCXSscifrS7m7IqbJxrHWwND8ptO4Cf+YY9aQST9HLBV3hvnvuAz
F2bppAcYdl8YvZRaSaHjDH9ItyAmN5E9uSuJvmbdrsw0Bbuspa2dbSzUKg03bc7z
gJzqgMBZTdbl5wd+MIYnFoD/rWU8ltfoKRUqn7mTs/pn/lUWkunzYA4ja0AASX55
e466ZMEbCruysSF8FCB5RwKu/p9ZFgExlCPIJRqam81Jmp30iF/izbrlCO7I2dqp
EaZt9kE3CvZZxZWIA+5itf3So8NSiVL2PyD0rsS4NoMfTBh7Js+ITMY2cvblc1LI
f6R0FMekZZdFVpuRpiZE/latNZqXYuV6bRE2/uX0Gtnwxrb5YJOPaZpOtdK3W4cn
NwCu4C8NSB4M7gEyA21eIoTWhtPzlPMSI/ovQITA1+2vzNSa3mjo2307oXknYSzu
2tmtebHq5Oa8ZnF0H3bN3BETqx3XOHSdNM18t9zEvAA4Oh8Fq2xsHvI2Zqjn2ol1
b53V+BTY5KzVGmMNHc5ioPaxxfthKPIQstVdbO93BzokpG8x94d7IzEpyw3q8eiE
wCdFNW9yaHQ4zeH+PDlOejW6JoYOfh4k4zvs7m7qq1jVgmY7ET31pFNziA4H66tw
9qFiXOoBdzjBXZoD6FNQVHbsffjavtHKEtEDupo7rTvIqATQb4k3wfjOMZiNhQyQ
eq/HAdG1vQaqlhSTsiU5Sn02fLwaTuqpkRqi7hQXcsY8Yckt4kQRW6+DHvCTFVG8
P1yU8B/Fp5e6MDVzQVlHZhOdsBB3eYorvDgjbwic+0sYYPk2nYIMT1jgxUTqMlVT
egTNey0zX6p1m0AVYAcOG4KZwBc2mUAZebQjyUcFjuzuyJ/Z3v5prf9AtAKGzK+A
FzMSGmuqDTS89Cy2ULJVL3QtMyqPmaGJGf8jNkz9F4ox5GMtzeocV+lGmN79pJny
SNEMgz8C1ukwVIPfTxOMT6pE6Llrfr6bcKcR3TnGUUx+KeS5UBmUXZsGrhCIPYNd
2x0kUNtn68kX//PCF+IsafyClsFZ1i3ZuhstuxejoD7aoWHLwvF0fpKquBEpUXDr
mEicckNtC/Xkopeu8+vZB+lcRf7Evj2AS/NMOU1yT79HuwElZr0OIShwZa58JlC0
9/+KnFzi1arGW5OScwB+MlzsGcPnl5mzDGlAbeujK1T3eF8sUcA5O4EMvblYZniE
rSNpK+sp7c8xRz9CYfPaQGIINlSp1dBIjyf/vBRttETzfkCDAeElq2Bajd++WcDZ
yiOM9T4bpD/hUm5fKVm2anxiJ0AYZrMFAYGah4Br88SLM8EYE4J3ftNxZOPUNalB
S2+usAEu37QrtFNk+FBM8ZbNlcyrCuYUWaSPr+kIJXXn4DNO26lDk+HxGshRk4tX
SC8+oFbBggaFu2L8lPzXozSUcbrQf0TtSzRmt8sSBQKC+3hqwPxMNm9FUzSYI56m
6/Qwp2S8Bn/yF+LPaLT6k+otNvG5UetFKKrxhiCcBOb+3wBqVPSGWMSHrh3W5p99
+iViIjWgPD8diz+UcFAtG/3zj1f234t5+hU8IZTJThKEWeUrPgwxeYcEGQ46N0m3
bdNeXXTt4esOxfP/Tth168eqZUYmPYfxVwqhlKmr8M9JZY9muN2rkl3wW/1bF+9y
ii1n+DaQ/uYefi9qd/xHEJcNY90ffW3CynSBV4kq135q1OBUyE+K9lS1qDyOKInm
plu75kDzN0e9x8JObisp/WYy4mLc9QpOLyzaGK1TgXEfZF/CVjyjcc0GbYx/84A9
nMyn7ht2jr8K42jsEFNMfi0IWd1NhvHICcJ1Iow2OtlylaJBEkmW+FmYvXCB7yA+
W3qegILIcJY4+keyGUHCy8PgCbJRIziEmr1YCYiF+0NvM/kidXevJ5xPtPXP5Suw
Izl/Og3Ih1RezTcf3h0gMxZlahGSzi4PLW8iB0eV/ZpOxa03W7hY+Q9ucG2qgXTo
1eK/J+WviyfhuyghSZ5yaaqPqKdBEGQYEoYFYKuEedpwKlzJ8nnHD+6LJ4YdOoXG
bT8aR5dScB/KRmDYaDKqpAATlOpT7CnOngUbjkwF6iKEXKSy88c3tFFPsyWUgUYH
T8mhFcUyxFJKIY8KJWaLft4m0uL+Wuzc9J/7mTEjSedM2xrYCm6J/VEwqONkZNyB
CAuwLnS7PuZtSLpNBV64+71qfgZBgy2HkxOK6IJtgm9S3PqDHQAPK0TOE8DPg3Md
aHRG2tx5NCUeL1YllP6UeoLhOibb+xvTW9Vx72TQw21Ege0kYTK0m9ZaXYwmb92I
yR3nrMuahg2aHMTqdFf5xqKlRLposWU6MOinro8G5iJVQcJF9pwE3Z7HYB9V0MJW
jZCExMYC31oaNCOjXI/9OpRq0mF3L1PEZOAufST97rRnxHyR7OA11Acr8fntJ4Vx
SCLO2lUjof1QYj0gPiE194Mff0nFKNtIr5Nv3utdqA1kBsuYOB9cqQzO62qYske5
sGe5ft9buw7SoOV9nOUomb60lbGWqeSgPBe0v6n5jdVehSSJib2q20if8XN9dB3n
leEjMjR1i6Tl/SUZLvfYHOUTF/SYAbToMzYWHq9xrsi9vwdr8gO4DAl5zfOfdymf
I5Ri8RpQWnGViBgQ3f4RNUDFK1ED0Z2BPVZ1YmBxe6DP00I31MBURGeGdvtA4Giy
zZTZIXlJ8bgs/yQze+6zQv7xKmRrXsZjhtK8ftjRRQVj8inpy5b9NlLXdPTah+UM
3D5+SdCOO0Zy+X9ZmKTKtCjthmsPNO0wpd5Wb0NbDarx7tMJs7KQTlWqd7s6ztTu
aFanksPA5ivw5XhQcdn+PdQlKjim+N178DZ62B06rfSAOHbYkO5VqyUFpNXcfAM0
KnmqO+6/0ZvufL+84t6H/VLR1QfW3OImg5jJHWDPdMTkTDbKZR8giFdr2aq7EG5A
CX+IdxJG/Ltid495C/OeMSCeEJdgC4KjuLRDi0J28c7BWulhwtXNhC4x24YjrWhB
`protect END_PROTECTED
