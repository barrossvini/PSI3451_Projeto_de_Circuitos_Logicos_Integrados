`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6x+HoRxTuHTF5SdO1MKkMuY+mO2dn8QIqa4NvzOga8eqpAqyos0AuHGmsg+lHf3b
mi86TgrJGyeX0eTV6NIAWWYl/xgnMtXUxrB/jk6JfRsiLX1dCJou8Wi2utgrVo9P
/N8abLiOXUwyA+7+l+tTp3b8YGhOilzlVi9SxY/JxQSh2gDOsp5+B0nceXzP8Esd
UhAGsKKUD+JUfBJQTgL6IP1COpikNsCexR8H1ug0mVbPITbRFPiQ+/yHgIrmAT+V
QVsSCufv8U5Y3DPQ6ku5cY6mySyW9yINfhHH4qTM2EyYDTch6L8Z/ki3EL1mEoAu
iIxO9Hl45txezt68kHSfnnJFHnjLz56wj2RRSOT97RvpdMohgDgOJFIW1cNn8h99
6iaicjv5ofYHUkh2mdck9OhbPU31jxgNlP2p8NBUhuMovo4XbDVj9UL3/z6djt5P
PVbM/2WMSNLhaXb0c75cOfvs8W53KBH1269ZgQhpDqrTi1hUBIBJuffxP1XogF6C
T/SsobMcfaGdhyXqnYI9SaL77oG3m2lxbOmrycOKNH2doveGpTxv+t0xBiCvOEVH
ISGVyYqEIZqGv2y3C6WoRyNQoOjyAVLGFYGXw4E5CwNFskuKcrzBJfoQ8q5yIVjq
Seax0KyMq8EyiNZb/yKv8pazIYS1djktSqGadnFFJURjo3WVFvRaM0cJJ6yAHRYs
DgE9CwQQH6ScXf6OVcprWKRSSIgbTysrXh8vZKhuTQRd5No79AJzGKMTMRu/O+vx
YVQQwXpfyFa0eIut4jIOeI4G8nS1X+PHI8g1wDWEbORA52o6Cy29nuMDXyjNKIUW
GIOULBcHrBQ/0MpyN1d4F2f+Z7tBx4i7EZxW7YGUDP6Ho3eGjXWqLnQJR74Gy5Jp
IvWWqmFnbi0j3T3Gx7bfy0aN44VQRstRJIW9m6jRbeKyT8c7QAk/Yzdc25jFt+LA
q0qfC7BBI7AamZjFcz5tIhpBZyMLSGFI4R0Mm+jk/JGgqE8cDXCkTZXEbS8l5Hks
dDmhh1VtP4/LG36rcNw7q+we5jD4oGrhl/oKx8Z5wrtFyYvmXCZkVaDs8oAsF2i+
KFJmTMAlZZU8Kc7VSNA9jRDfRmxDrwByIQR5X3m6+AVYBRYzENBC3TtjyMGmPd+G
hQNAw9AFf3Rh8HHS6kXy7kLsvvx9dU4Lt+Gqqyaq3vKpFCWoMARBmoT3GYduncIq
EbBDZ5lKpReoip0bxfzmqLuhUI68BdNk4wn45SkqwSuyffPbRdL9ze1UVYEciOPp
fKmuKlajBBFWHNvg+BoyRHnYR4umyWuXDT4C++L9R9QT92OB7a/xYKc39oD8qRXc
CWk7nvezrnQAw3kvoiG1e5eDcuCA+v25DA+CgrlwM7Xya8Uzchi4EawlnDLLGg/s
FQ3Sdkjs0AvBtWK18e9Duhb0BiVUV7we9hdWi9/LWH5bgjjERZl6iYIvt+0ZWwqV
neMsUR/AYrLE6KURvCODn5ZRuVTpoU6ao9BFDaow3JiclV28iqE+Pw0Nq9TX1paU
bwZ+Gboo1mQsqiyjckjcurMqSvubIaT1InauLlpL4gIvbibuQEyP33d3BRZ6pu0r
ebKVeaEjnR4jSWqMVoVPy3MjFP4LugFyn6j5A+SZtO2M1YySyUCeMQpXOhu9iVU3
Cnt1viZcJhXf4K6ukTDzjE5C7RdS0wb5zSDA9O3KcQpztV8FNK1a55Qquq3zX1q5
lSmD0bdeo0r63KP8c2cuomBZbG47DyVWk+DSaDnYPdmzPgrryGgWtIxlgwVvH45Q
Zh/AjNFg5TiDgfz8D1xlXepY4U5bAz9zsbxOMq/Fzy2r4/W0iKjLHGovQkdg7vxl
fhmAP8wuH2hI+ZbxH+PKhx5MJzngBpFlGbxjwAhHRegjfpCOnqDelfEON0H3eEX1
u+5r0XxfgkGRN5+zvJ3PP4lH9dNqYK3LgWc8wMiyCH3pSRyFVxKXhjGa5I1j/OEw
8prRQ0oAKx/QmETve/TyJeOKhHnAPLT6+UJWl933bY6VuBktQtdEgzbWQL2Rjtq0
l9ut/cSHNZSmW30T6GeODO3UGBKHbBaiMIILthHzl/9UrphladfZGvg1HkOLvQ6w
fgD8YBLCkXtcaC0hQJh0R6M88lGA6ds3mpp6IG5ErhtAl4f9wWPAgSJV1MfvhrU1
0EI3zdrZ5Mh5vamUjXG5XdlyUvN7JGqR8vCFj+1CxV93Ybv335SOzVgDq2X9Hb3b
dWbairo6DRQqcaW/A73bHNWmQ9MUb4ecEtGBhuJLz/EKirQ+gfYNJOcLt8258Omj
VWgzb1TUh2NfjpZV5Z7C9D6UiRqpWZPzm7iJpOtU4KGCEXOGK1hEeNPeQMxvN/97
5yXU/KFjMAYvDfjdpS5ZU4SMRqg82SELBIzGteGVfJxeAPjmHhd6RISDn5uGpgk5
nOvNkOOLyXoA9BOQcTJhC0RpnNBoLqU/N4tMHwuRG1FcbZfbEjqBuN8ACFAwvkFh
5dhfhxnIRPgmeeRm3k3pE1ZFMdEWt3oe1xPLSTeY6LblZ2hsM4gLGxOVYy+5X0lT
Lg3HvhbWuLhLCfJ1NaQ1AnEsiccRn/Rt4n80z6drvfesqnxCqvmlwVwwDABBr6aF
39YRjqWO+GXPhb6qu+opeYtt6aIrFWBmNsBWG/lu616HJMIzb+2+h74cgRoN5WBJ
wryfa6WmLYDcDagxLdTzgr4Y3Q4nZBNJSF9IuMKODsYDK4RY3Vbbbq2faDNUqd3j
BWK+4jrtn3yoxrjOn5h09/7vG4kM13wukGN61lCJUpRh0wg6m59fSNwXlXhmojqb
mzTy1djGnwDZufxSadVyJE4Fn4zv2g2n1bF3P83buzO/sLljW0Cs9idjOcj2G3wo
WuPRTz+OxDDuMWAYOVqjOYhcay5PtzZu4bbum1T2jyMdOOUGUH1J+6eAuqvDNRnd
iCe1sCN2dKqSQIpsOcP3r4rT9jpdb10FpJ47qQ71OAHhjEeN5s0HbD1Yk6tC1yRR
vwrqXljorMW1DzgLVt5uO2Tj8lq1Agpw2gqpvHK9WkYkOKeQjYGzCOfIej4Z9/5q
5txO7xHSXYWQF8GY7hUJVI0tKjCKRSucz0Gk6c237QYWXPgrT6E3Qd9sDb0lUtTg
/4/1Pyw2NiUkTf8pORlgwNoaXvt+zae1ScUb+LylVPDmiMa+0HFd2DMrApDk8Qy9
V8roQLNG2PTHRbcbwJl6y+6wwC7CklvELDoN2Qkgg0qeOtWtMcPQbXPx/Vy5zRLz
ZCFQ9zR61nQHKy/V+nQiQ9Zu+oaGab7qsg9VEsV/xOFBuraY63R8DVrjW//7MNcH
A2BjgJbX3he/5HAGOxSCApDN+CVFyIcJQdayNqQZfmpu2uq1JX22S+fb2/vSMLm2
01zKdfsE/nwHJ48/r33ttsvZlLMqtEUoXQc8kJAqEBlRfa1wP8P6cKIRXe7X4YFt
GE8Hph42UfTq4JGEV+scm5u9hFxYJ6LSdNLxB7B2CUatBzxLo7hNzONmpc3XHKXv
SWzwHawF4PILJ/JdJeR62Ns06fpYdYFm3NBmhHDTZBVvLGYp9KhMulcwVb2cAw4y
ljbowk+cISVXqhMSQzc1oAd8hTfZJdgtPaKUHXut2sfTicSjy8i+GNm7+IqstZV+
cmz6qpBcZpSHxpNy4rNjrChGDCsbVpn9nEB+Z00zPHw6WYPda2ZIptSoMxeQurAd
KjsVzjTc20eNmr7/ms74zAxvypy0+EQTu7MpQhbLh7JHA+E0wkj0yumpJxsN9/wg
2j9jhQlJ+ndVMtEmtODmcctJWX+kyZI8eZY8JnXY3OCJajChDWZvTmgxTrtno/iN
ilUUrIvzb7itIkmkvoIJ+P6aLsvP+V/g7o1ahCB+K0h4jt5djdw1RA6XB4b+I9VR
ZA0lwbSCTHeoSg2TI1N91BLFjinExgRbgKAEJ+gZFsc5ppVwP890YgsPWewA/4kw
BZyUjQ4p1J5ViDl1toDrRmr0WLIBxRYwiYM84n3+oiw8zwgQg+6QK8U5fROhhnLW
DfWjVr0uUMNQIao2lCQ4NSqfg3SZln/zYJesHdsyC2+mFdETNc6PbTkfoYl6qX5R
Lx5jYPmx/YFMesQSGAqDR5OsZDY1aDys0fGIqcs49XkQmVBX88BZ+ClcrVjEYYaT
WIr80fg07MrFTCRHyXVD/mKHP/ZAZEaamVE35lxgiAVtkrgzYIJZvyshUxrB1kaE
ujsC3r0SurHQh55ICrhbkS8hujMIR+tE1Yz5D8f8gb3gS6y2hTu4XbYNwp6iM84n
x8gb1ySFwRjSbEvpsc9EVUvF1apNP0dk6BjYBkOaWAweP6bNh0KgJHoukpVXaN2+
0VYj2GCv5AsjC+eDoBIyEKlJirh7zrIxdbmk0WG6PcvMCY70tcagKtSioS1bFYQf
qgYRb9op8KXzE/bqRkjaUzO7JRqTQkJiOD0m5g1Hzgc0f2c4Pv/pwDmWm+awmcaE
wtMp0zcpZZO1v9xVi08VcFgnuEIK5vKrsmur9tgdGKt9AnhnNMETJgnYrGFn+0En
2CBpChHQvoma9MVw5dqz/uvb77Ny3OW8K+26q8k7X+ATD44nLoodhizwuSeNcMqv
DXsABrJc/Swz5F/qJWTLju/zR8HGDw07XmOwkTz0/YiFgGa6/5ItekUeGc23CnGY
ZIL0gsahRALmJ/+juAFJs17wFH7A3l7wqLhMVOzZV1Zo/t1YB4PlpeIF6TXlcjoV
6XA8lSdo93ziGV1r+zbnU3wRHAxgArew1FWDmouRCYmEkEm/XvDEXPd1hHX7In9Q
ll8cuYHiJpzTT/FmMs6Do+H981SgD5pYAaAZCGNqFWTSUycTx/jpWmUUZNjXY+uG
odX/o7khzhxEf9Y/o2KKP1ipikgeOYI8xbvnHzPnzOwETp6MFOTTJ6MKsrIKUZTp
dS0WdBXVbas3lLETxyEfuMfftl9i4Xj/VapDYuRFnw59ZQQPszaAdHxk66Dxv5u9
l6UHksGThGWZoKYG50e6ip5LemfhnHqoib/YLMImYvbH5PHVxDWCtbs2pw5qGos/
H6wUnvkLTBzsbZFcnMbmTAnUxOGzGuJVAl4vKn9LCqhqAjYT9ti/wtcEtCQkjb/f
4mqEhvdkeuJs66gYHk34mHNZodhVgNcBuKbz5DJ2VYTVdJelezjee1znTm/sfING
ATldCua9HsYwcy+H4L0idqg5z7TdSayZbijleLAgI8iQIfLUYnZQkkLBu6qs3TIj
fc0dAOAyKlLJ7MzHeetRwjFYRlSvP6JFztniV5RpIgMCXBfpKDyD9/GZ2trWWgbS
2zJB/f8ATHKGl4iBJ2C9ZXEogFWkCIztgVk1DY+b9GbrgEBPxB178zCUPWP3rkFH
8mwlvebi6+2wdHufA2GPgIx2LAN33YFTt5GE6E0Kcyr7c7fsyfQ6EEAfJ4iRy0Yy
2COMOp2J/03J/jV5vETVESsKAm9M18+CYFulYNaAh54ZFcdx/PEXJhGdq9ag5JqF
/3eCNV/OvszNzH9oEcLG/5czD6PjM5gKA0q2RobA4YgeVdfVnsFmrxlKfcpaZKyx
rm0/xYAoWSrws2HYj+mfqKajTB2X6KFNcO2XOSm5blz8OPLK2u510FHRZwKuj0zo
LyWND4DsYtsOZTOPY3jeuiAz82SGj+ZJAqRGsOaG42oLk+vEJ01aGqh1423i/xFc
4ekYyWewsmdpTraxF8Zh5erRl7lTA4XsaH8teQ1FDuTBhK/NllwsqITgUIGwjoHI
Y6xFHYLzAXM84k4pXpFjoRuOVQ7kiELchCzQUaTb4SpgsEThlk/qt/QwlKSb1dqR
tr0WPUH1a65ILwmzah3ODxQW5bgKlfE2BPDB6byUjc48wtiKNW+MW1t4CIPtk2fq
bhKWtDxKwgUX0wJzdfQeZOd/OPayLh2NdZhZoFIT7QQsnor6AygtCp39sChoW6ny
u5rYUxtjvwSEJE8qA8CylUd3eq3qS+VnSmYWV3i2mzw+J2N+GrSpFq1DOKWQUMG5
cAOZSaZ8+gHHoyA/Faq/LfZd0u1PvY7n2/5q/0vx0s0U2LyVatpo3/oy/o5gSCBB
qzSCcEQzaApOniF9Y45ue+VIBGbHYWMFrtOpE7u2ttt2Pjw5FmtnsHZHFh0HpT+w
f7qN1e2y00UjNRwERWptHdbRVD9Rpj1LzNWRGm06lmGurcWwcunQpBSCrP93+e9n
2BtSUQDir09q6cwt6XMv+aGpe4Yl94gy0tAsPwV7RgEF8/7jQmBV3S4TuL6asTVe
cijR6RZdiw4vqsqIS9WVqQw4oC7awskZBK5oMHKlrm3pQqfg8LPwn0u74I7gWwA4
supNfD8qbk67HqthTGKgco5aCHJDc46DoSqVfOPvcGPTm4J+MPIGm5RPa/O1i00V
rCMTr5J7/wVbU1TwNtIdJ3NSyUC2i6T6/BcSePVUEAPxTHTFRnDKtRax0/VN/fiN
CTavgCCVK/nGYZHcQC/TLjHtbfdgWGpfEYzjolkjjvJZAhAcc5p9yL/NPJz7MtYp
a5wGSYuQVAElTHUuuHZ3iiZABM7ELWxFeAR6DK43JdeYK0A5P/4dwJhipOYaIcZL
oo1VGSwnaj2sRCHax1pmyiYdpgzGYOFz6z8kE2p59KkxRmxK/PYs3XDRd8sFwWG/
1271GwyeGgDk2Gn3lmzcHgG/cY4QBEfVFJOwR1U39NhPTjGdyzPygNHySamD0QC3
A9e2HoKMjj8fUZ50PTLUOnv33w1wdgVe++ZLqjVunx6GlY1fTsDXARk7efXhvNf4
rofuYJH11oQ70Yv2kaub2zKlOT2hMZr9HykDHMQIaZ8qS0HAfaOZLqtFZ3rCmKR1
IZizYPQ9B9M/t9cVsMZQOJcnKZEXu1wLXRJ/IZwAKW3U6miMvghZhm03tCLZhzYq
qNIJ5rDkMpm9/a3nISVEB+yafBOPczSXydUATta+P4dJuIgZxeqUB86XOz1ad0BX
6jZGTA0zqPfHM/MZrS6tpEXiG1EkjmWqaSgrMydR8mKoY3/VqFvsEnYhIV3trZwO
fr4UUMM08+3gLlckwU6uXScWGR/8nHDHSP3h0mVtozhDNa/rJIHtfmpjMYUwMwes
G6wtzvBmRfH3n0+ar/Tk4ziEnXpaPrStDbtBFJpDEg0DXDzIhzcGBX8m//Y4TkGs
w0VjO8eye+nhIcSYKbjZVdjkzGASv1eONc8WlD2BfKYg7GAhZwG0Y/EdH9no4PVy
3eZtTkKox1eRfXh/97Fh8nWy9n7CBVvR90VYfavTcB71xx2tlWJudJRnuf0GI5QF
Qda++NsW/r3ASgR23lWizA==
`protect END_PROTECTED
