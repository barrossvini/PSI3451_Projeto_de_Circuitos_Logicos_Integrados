`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jao1UJPFZDAbZhp7ukOM+bNQS/TMrzs6XBYu+/RNdHZZei39WOKtAokmSsf+12wh
gUMangSDEOV4LzktzIZFGR+uZmt/wBnEWsfDZQ38fM22H0Gb+EAufxw66Gc8OOq2
x/5RSytvg+WKep4CQvMLT1ySpM9Dga0Zo8s5xKPPsi+m7C6peUDUwEbZ1m9jUGJg
/nbkOvXcFOHdVgEH5y9LFzshvPmEMW80EwyreE7sWMZgxd3u3JKmvCXTYOvZ7wJk
VtcDSuQ9Q7CB9oEfdGQ374EBaQStwSXrm6Zo5QD/dFAZimMca5LTwITft3ETzuGx
mChrD212OUjSnoL89KLqOOj+cIWoFa64Lw5X9fdU+mmr96EWsKQ1bOoUO0Yp9Xeu
CuiduI4/YqKVR5H5MQR0tbmsHzJ69uBxoH8jb7Ta5Zegh67pipgTMddvzyu69+dc
K/EqaLURE0fM2ccoTVYrFqn6IwkiqQqUH3dGsEq7p+G2JEZzXO1Qlf2u9V7cMMYe
C0TyLiUFRDmTAiMAuN6AQzH8pQ/wx6llNSP6M/1ssG7Aja9XY+sYUY8nlUXiR2od
zOWvSTYnSXSFF2DzWJFRT67k3R+Qxw1aOMjMU7fKCsft7YacgrgWzAsgeLxpiVbg
8wp6rCNLielqIsnVxJ4sEBOludj0u45TIComeJRRIYNqndx98X34G6w/zeqh+h7k
/PaX9GPHaOdktgLm30mKE6OHRvnxiffSJkW95406T2ShDNJy+wyVlyrO0pUcGuhr
vGS+/e/1UB6nzUGnB70AfxR3DdsOVOqITpHRzRirO0TfUtdM2cx40ootUfw75EDt
ckFx/DbpSZjkTVcCY/EP8Q==
`protect END_PROTECTED
