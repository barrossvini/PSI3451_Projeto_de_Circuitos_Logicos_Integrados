`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+x2yKZbbI+7SN/InqAdzfjZ8BIg/BpxlYSI8ZC5DSalMOVJHfopCW3Ir+kjLIKVX
4PkQHVisiw+vTMNe6TgXB621yREnDSrLEXi9pk8iXfybLc7uZmar4XvILlnFXcrl
pMDuhJpbcCHs/r8L2xWBQl6Hst8IEyafeZWCKSjsMxjgA5c9kOCe+1TJCwqRvh4l
xbAgWz4VTDivENCxM4issv2p6jNXM4bZklJ4o9viiNzZiwdc8msqouQHvXP5axy4
TLgkh71eNg+fsRzM6feBx2JJj8eIYB62VUV5043Ird67jR/UxUYZn6wYx4kXWH6g
kknDGZsJ1DgicdGLv/Bfw4A5YWDPg2nQQnpcVM8LLPWxJukuCNxFHUR+8dgrSW5K
RoQBYS+op993LX1aehIHV90xUL9egM4eIKDI15gtDjsVa6L1GvIh1DgldTi2gfXs
LUZ/ghzEGVmbn3TXQS3o2QAg0/G+tF/Nb/1uHs05gSez7XSUSW7Xq4bLAbxuXM1K
DNnCFR8rO2jtM1t+JeRx4JRNHup1EvT7KolT6uqAP9WbYe4zdooiKOoWUu1xwKcn
H8ENziI3IMNncnx6bZqWXD1TcFjw/pgBATjtzOc6EnwwsFnbFD3X5dCQuDPnzrjW
Ijnr5I3ngzfB5uBaBdBTIzc9Zsp7WUXiZSpuuUc2ZWqviDj5bl0tjGNX6etVlc9X
NJq2MyX+mGVTDPyKWxwKUD4InQx1l0ZFeG0ipCqDEQ/ILdmHaQcLgsdBA+/yHO5+
imgPjkbnuosg6Qvljix7HVkEJ2r+f8/pW2B7SxEoL1/b/6mU7ud/Ad2Q+jLYbuRc
cg4qANEEF0xlHlISyhbkeXozC6oRDrAVv0Rv8p26lRMEeZFyDFMIitaiF1MvOO6g
P1PLI9e30L4xEQqd11yJbsGjeL9ZHpws4jZzON5xVUsspO+1ExmFHPVxuGUSL/7L
UmOqSElHf24AbzDHzMmFd6OnM8MQhEposFheFYUSZoYl4WmUyE1bQ2i4DCIhGnHF
yPt63DxEMUTz7wLyKyDiC5pnKjJZrSEeqmSRtuAue9otC+HoyWBq+YuRYQk0x842
UcYvYwGtxk754VxTKIzEe+eahdxqRoTt4jLynOQTQJjV3EiLospQftvXRUq7THHM
am3+0pZzX1Sed219Srj4RXCHnj30jcXut2xOufdOZWrjkAvPHtW7z/6a/HhK2l9B
ITHJUNRdjrFUxn+6cqtRifB/O40d8WgfnVHZc2DTZFz8KbuI5B3Gvp7meEL2oZzg
ZyM2tJ/A91SYBRfRbMKLBbpBfDI5GH0KmSFyA1sZhzJ6z1wdffUXlG5wGSoMPty3
H03ZA9ThcztEDWbexXhmSil71DqofU+2IAOh38hgdg+uaEu3ZSp8Q2drU/HV5tTD
yxiAoJuuYjfaK8gbIC8bx4yFWD/4JLnnxcBxvvBuFHwYOa2HrgPzKvCNrNtpgT+y
4JREmNZIeaObbOGXq4SzETHJ/TNB6ujVN1+EeFwt53wJBl/qXhE7fnWrcKBgZmdC
YQ2CRfiMyIPb8pvWOGzw+xBjng0N03NqQMVIfPc8dJLjv3UIl8flxA5i0V/Dkmm3
5dtexG0OfSe7epAFpMfoxPbmn17K3n3Tw7WAMJRhbWQXbP/DVPZZrWuCMTcMlz92
iti1pZnedvFjL4PthAeZkfjjD6lvlc9VXAba+85oUSrXbF+EPg6N7MD6uioYj5Sk
PipDN7DR9KBzmY9zVBUATspfHRZodFT88cZc2U+MYz7XcQ5my09aVwH8XnYdYKq8
lj9HW9M3DOVe6i8uf5EwbkyD7RLO8MUsNGj0sE4wwQfAQeCZIXXVRjMql7+mXjNM
Nd38SUasfMsbA0fkKZUZ9eDas5T9hAg1LVmkmPcAACwVxTz6HX+wgLHCYo0gbB7W
ZUD3VUdSKDiwPugpzQhLsAeetlTn/CLsif40ost3HyPpx06DhYFH5PlvTbKvNl7k
luhiq0QBEwMzUNpKAfW0t50GTuSpMp1H+MKkV4oOBHcGluITboKE7VmoEVblfQMH
DWOaDikhBZnD5neCoQHzGCq1mzxxskGqo5o/8KQfdjC5RlQ8CLFdRDRWyHugw3Fc
VpleAR5jfaMd6o/woH/aLiNgPbqCr9C62AH9nanOYpyCjOgy2qCk9xwngKpLFt4j
FIEH9dzz4EiS/kBVcYx5jrdN4ycTBzWzCsGXtmRYTYN22hE0Dj5kqUdgx88VJ7HL
4FKoZUreBIqbLKDrJFnAFURgYEW9MCMSkUuDXMTgDqlr8W+Ba0q+NblWlupFP10j
xazRV3GL83b4OXjkXA9nf+GRdz0Rhhr+RopY99GyXIycrkguogyuaTA0wYx7LSbN
UxmJw1jWpOBSAfA55hM2ru+3+o+KxJtWuKyiibsnk3s9CKYMn75yxEny50xYsXAe
+fMdlLZSywfgwvRnSKof9siQde9q7fpqvR+yfMGn5h3B9zxzl4BqeRNtlC98bVxd
k83Po/nSyfAAAiZt/574ERqSJktsNaqOp5bYeFsVo18XrVG4lcUsqIoouLCPuCf7
DzTTlgY1YIZLzVJ/QdnMp/ierbSCWY5wl4JbZKnfpSzr1eE1fWvYKOWRefGNpgFW
KOQ6vQwIoRPI3hraOrF/wM/+dG1HOi34xs75hpP3Q2JWSlrq7u49v+KEkeUCyDZO
F2GmC4jieI+qzBmUj9Mt/blB8kp2SBU8w1hk2+W73yVmonsFzHA36hpCj2u/3W73
eFxbSfjxXMm2blULUQvuwpvnLUQVvfoMLfZhVRZibJfV544DHDWiRivxvL5YqaAK
GUAj8SDmxiN+vUK/lozTuUpmys7XlhqmRi+nEFSWnHo9J9rG81U1c0jrBfPMVllY
5JKwePOYHtoRnPPdLbImNJ41yqB38betxhiYrwPhDoOw0V1xqU4peyXLNS167QGe
fFTU/fTqLYJZkkuZYJAyxI1lIejMaFRfpRWLR666R4bCexum7l+zdRggs/+hb+jz
D3FTFOZJOkb2RBKNjsFOxUbDGbES1+uEe4YBju0gjwZNyeEOCBf2JkZk8CL9mJy1
Z8V0woFmbtn+Z3ruyvWpyl2KHgxMc9BjiJ9/i0WLcaqZ6YZR6NMVWkw2EJk3tn92
5DGr4yFpGgLdkFIQbUNcoKwqlhe5sZCdIyRoDbovEYyv1uIiClquqRPo9Hhe7ZBi
kEmjKl2WgGLXx+V9phA+YsOi8XDGpDfiC1Ps76I05CTMpnQsPQapzYxZrmYjGGZd
J8aHLn21NCbSAYO47iSdck1FsVg/z3RZGTMksVYrF49lWROCy4rW9PAGl4Jxx7+N
p2ZakBqBgV1Ui36QhWMjZma5acA7oXJBC2CV2ctjijA9gqzEl1AkTcGHE2n7XZYF
cZIc5Th03ah5Y5cwM43ATitYCpODCs/oW/ONFJGhVnJwR7tqThBup7tcabT3eZ6t
F8YcuKHBmEOl1SwS/EJtOXZqrOnBx/QmfVjFEJpU9FKyLBdKpMpLl3LGBvlMHgPU
Ul0Zp93IFici/e9V383LClWggtUB+Xr+BF/mHOeiKWx9xK1XBeXWkFDujhenzVJl
cOhL1Q5pqFac2lwXDwEwzSl7sd9d4n3w4gWICd7N8TMHEjHylq7lUF4qlN2nVZWZ
S41IO/ndQDiDM8LkHOdot02UrdSXuBZD2aDkunn2Xd9WJ/M1rlPZPbudPQ+Hl/Zw
mi3Mf30Rfw5FGZ1LLUfbHncJ6sO9E2DlbsF5bSjNdZNRko3ZvcKfs0osFPH/Qn/l
lidhQLTIIgnvJVcQR9JYY087nRIOYpkyclY1cAtETtvBVKCJ4EGsqIl3tsRo2FHC
brInW+u9nbUajrXRAHr9BvqgdhB6neEp2gtwq71+CG4ULfWVBIB1dXDZMB5uisbZ
zjZiBiZ4LxXxr73zWKzbu6gm93M17bk88EGxSlG+y+q/cNCriIaVJNLB8LlG2aHx
xiDtOXerFgxLJ8Y+tiqSMs1LCnHZYgqVoseHQyZDj0mOBAiKThP+D/qvJ5JXNQ6l
SZ89HpzoIYzJJ7sOzj+8tjsO6JWQuoZVO+Wvj5RRpADFTOG6T5WInPeWlOhRJNPP
LslKTIuINo1oJmzniRlQlTnk0OqS0CnN3xMQzyiJ/tAbHXHE57cY65/4o+9ilA+Y
sSKX5O5uDGNK9Rh9ceM0q1EDWFPFzgwHXGmKj0zeLs7tqWq2aiflJXGO4v5atVFQ
9ILz8TX5ZqvMSlNE0d1VAD9KsJa74EYOQoRoqXN3/8iFHzZ4LylaRr4I8C6mi7PI
dPDKaCpyQJJBX787/VA2YtUrG8lOFQLZbhQCJBwIapkk+58ZksvlL4olc38mgY3z
v2Qg3i0hKaIzxBcxT3Z1QYeceGX4xDNACP6N8WI64xmtyWNHC2j4cImKWcmDLVg0
Yr1BO5M4HJBHvI8cbfUNFTTrGVom9PJm8vKFEN3rJzBWrvGp4Sy0/x1o9agioeGF
68eiSWnLs0adfR48Zd1wqb6RdstNpBTLpssPcGNodPk+cVku+HkLrr7/HMelp+S1
Dd798voj5pmQXaUS0xM/xsoIUOgHDDo125Saa8NVu422hrEO12L+ssljt1GXSBsM
gTRTgQT3eRjdJuNuOiEAJGEtkSyRcU8vlHEOCyJ2+rBD/c6iCN9QHjEd3ORlBtYT
O94X6hS0uB3im/4jQAL1h5FTvVUk0ORl4rU1HXTau6sQpLqlH9MlSYl33Deb0nwk
XJ6Fu/6C1xwIOlVUft0L4w7biPu9QGRzF+LiPFl2+0zND18E4ryqSptw8lR85R4W
XSD9AIHGn+yNDblsdnuY7f/X9EjjdhN0k4TNDhbzSPR85NEvGmkoKs+hQV4QdQfP
CuAHyekFccPd6m1hmF0XwiGwZlfC7yiSSHmODJtau1M/3qQ1ePB2fsPm55D1WM+t
tw6U45XHV7H5uINL3v7eoxMKwKRrLlwNjO4OR3wXQrAzEpBG5b6a4a2ovpEpzYhy
fjuiJWpOKn8bMXbRrYgQ7tiKib1iJHda3NeL+7epWVJyUtK/2Df5OozU1r8IbIIh
POnFMUPJxY+yiP9sL4O+2UJYsppKo/K75uVIc1E7YhrbgUNpUTrhYI5IQWNNNOCC
BOSwO/jGBjOo5zx+kM545SYXMD1vP6XT/aXANJ8TR2XCxPFJBDgtGTu7gS+tLNfY
YXXr8KviU/qbi09jhUD9BZCb4cae9/7yXrAefvv/EidH8rF2Oblx1JuBStHW2JFm
sBs845SWWfiWDuwlEet4WvVzjVYplSvDBv/UxDXaN3PcTvW0BalhuLqC02X0q9hn
0m9pKuN0vsU38I4MZzpJGN6DlnPQ2rcySG1j5GFRMOP+DO3+uftl/yEKQQKEYtJN
rnizE5zNBaeG56niFK3/Nt1P0UGCWLKB9eRzAPo93V2W18Ca4AH2P1iUey4mjzx8
7C40zYo5R8HN+sCGUxn3M6bkYnfacWPTb9zREqStG0wQowvcd7rR7T0hUjZal8S6
6iVPZC4XdMV+iWtLolMf2iY1ONFw+1dCDD1jyBjvk9APURL5Bg7zLS+m0v9zTxUl
bTPfiP1jUj7m6aCLjZ32+eXssLWisnr0/BY3CtgqEdcD2FSLXl+C0QzLfcGiOQZ8
u7KlHsZtWNz08P0sLCnOYwGjH+nPL7cxNlqyrgp82HmBMG6Y+xdsQqjOi/ng8PYZ
x/y6YkyBB1DxM/Tf/jq7lFudWLXhm+H0v2OBA/RnVXnx9mhlmfyjRVl/LFHXKkv+
7j4fBij1uNLOIPg6+WS1h6+eURtQmF982VtPf8m+ANuK9jCgezEw9koWWWg5gL3+
wZZfdXFYpXI0MmtauN2DqqX93BIFf7PtOq/X7RAAR8C3r20P7InL6Nq6JlRB/1DF
990DbAyhhCJ4jXNEEjioPhIgzIwPo7WabSMYcwE1s7ejI9a3L3b0fTyfhaqM/aQ8
bupODGLsXxFht75zO9SVPgsh6hM0L2wFMHxehWAPdlQ6oVFa/zbtVaQdyG7iD+Oo
7/3Ot6tmK2mC+5E5TzuD3oeM6ppgvvTbs2TncI4QQ409+n+36hLUjrkGstze5iDb
axNuAVvD8wbH3cKRC3b6YUjJ4mWMTbB9xt9JFSCCNT2QYKE00+9cmFWVWTxpfxdr
mQ5UrlbVe9B1vsFfFEg150WIO00FFY3fUTeush3HuPMRKVXp5Gypyx754M1CGD2n
84MQKIoFlAtBQde7cwKWCUIGxaq4DqtNZQbpP4zVFv4U1dcyKOWXmg10+/7JLvEP
4AjrMJYjB1HKPFIzKQUvW6d7X9Ui9I5IrddApg5HSXINRiZWKIq0j6BYF9tCsNmf
tZuqhlgTRlmf2un69M7qvoAtDtt4ycCqakI5Fbbz+oR7m8SZ7poozpodk383nSWh
Tu2qEOurdclOTAmV4Mb+D97Pn4DaCtL5sC+6hfuxfmK9BqvIKuYDDlwmX0zPp07l
z2sPKpNtmPVvqd8jIQK/CRpurJq8eRoymPb2daZj6lyCoLZHB4RkOndCRyQFA1ep
hTBf5gK7pT7R81jw4fbdL7zrt3bOrVF3lgZNED4tLrjywFnNxdn4SjGF+4b96MXq
ekxaOOSkYa5TlcEaeIlSLhzs3N7Y4sxIFBVQK7ovtkA1mAhwboeps0ZDbQ8mZThm
Z8TURWZlmFbCiOd4IQ+YTyZOENclu2+wr7yI6ukN7d0OIPS7/LyxExeG/BV6iMNX
zHjCtfPntRwby1OV1tK0gtl2P+6JvmjX4NzVaOIWivS8N7GMGpAvcbddpTvuE13N
lX5sD2h5dh+Uk3gn5n6l/ZyabJh3NljDsiFQsyQ8r3+9secflTGstQceoEYd1HJF
+7YV9MitPNQiMkFmT9wdUKzWaU0pVEbxSeFwnl5LClWdDxVntf/MFLDeD8XnmDNL
STdg56vydLMhF2nbOqptcxu+pc+0tyvP4J3v/FPwkYubIIPfG/4FRe+IP01iGwei
FDZEFsQIfRCmq6QtZ8xNzMThAfscWKX0G+YxSClOXjeLkQzxWeQpnxj6EqFEqXYX
tBThK+jIAd2T033859OFQYP5IdKl9EFoYJSMv1ASmA30LVuwlogoY58qWu6/bga3
6r2t7cAHjkYm4ke7I3vB+jJ9h5A6OMP1sCLBbxG+/4tIF3Ni/uTbxh3em4ozg+vX
Uiyd7N27ZDQK888qd3/yH2vmr+R0hJGR1cgS1Drum7mOKRXX2aH6brODgMF6iW5O
SyHKGaHBD+ALhROW1UCtQEfTtTTgasz9NlUquCD+Pj8UMTc9AXrlVxkU/xlecFRq
zGGnJu4ArxTskUziaXM+/aFNA4u3nlgfw7TvJGqjoRifzGAYmbp0sxIf8SynXQLy
YZqnMEc30Ms1auc8aJtAYReugSeki3aLDi77U1FQOkCS4DGzlbGZVO1k/mWr9yIn
aldbYqS3ONdCM/e44xODIpz5BXlO+9nBrFYUQq6mIRKgTXWZ1yVWThYcOndyCTrr
4uKySOcCfhiPjf+7HwRPCYhz5VhFyuDSdNfY8tXaKjf0wkd7hDwJTxfFfszZRhlI
MvZpSpSzyQJh7eiXIkmEv/+1oJAKXO+aEnMkzz+SodOxwI/LlbVz361xYWVH/Lot
LLifUuEmBwZV0j3htyr/yBAs2g7OfqsQagANI4eDm4pkUtX80NoC2Ci0BECjfyrW
gMOoXsIuT9e9D0Vst9dX/b1kWHlb15a5Op5pTla9n+oxNBSsokukTWn/ClbQodNU
em/yeW9CVJHS8uyemFSXAtaGyoilVezhlxsgr/v3CQTei1OzjmUC0BJUZDd+gNJQ
3Hra3fp4p+TmUpWyFPhf1E59oe/XXrrKiCVEMr7RD9TCi1u5EUh1UVX/MzCh54v4
favxywc9pmfL8vBwRimVgHu5lR1aYt6LvC/R+Ogm2MXMIxRgdeadk2KEpAHdJFJp
N1ejznOORGt8DmHXQYlQB0qosmhIXYmAxiuC09MddtmL3mVqRUd4THM7pjVW3vbV
LIoq09EQyf9HY369ujUExDa2Bi/l/xTnZuyAh2CcxbKf/JTfsKTmAXJdXMaL2Fso
wkfSvcNJ5MI8ewekdhyq5e05sI/W+V4xHXUY9cA+SVlIVxQpew3pCwK9Vx+kEwN+
EjV+RnTMsHMYz4Yrqnlx4eYv4/uBpKAby0REviZT43D6FTBW6uuBy2toTQvN5Pu3
nRW90XlAHZmI+5QAtzjF6cMWhi/4JP+ZEti8vbOPLnbc+zELbTJW08JSoJ6rDQ0Z
ILqC7+m2CcSOLjeeSkwZk86+cy1X+mU83qY/YfmRu/Nr28RG9PwuXhlYtnomc0V5
2gvGpcHTgj34kqrFRoUI5Ew+aPNyp2qAIgHMnELp29qTW5fAgx1OBqsdm3D6HJf+
uo9qokl6K8jRKYZtTMMvp0fgL+mXEDTj+pNk5echKWB5T/VvPpvP4lyXeUhIQeM+
lhrnaWh9+KLZLVj7f40dCxvJRjOr9M7DuqCjEuBepjMkjblbe9+4P2sPCRkgr7o1
EWh/qhsxij15tXrmD1Jx3orBitsICWpk7Bcockxeusd73A9mSlLHMSwy4UyXNd8g
tSd6cu7dI1IM3+Z6SIgmGDKGxsvuLAqR+uj+1COPMjj/Z+VM7P8vRPw9cQ1KbAAo
QyVxM8uwbh0suUeF6AOBngGG9xl6ajB8UxYzd3dxZLWyEDh7/bi5PQ8cwD3cPO6o
VulxqZKigzjoAq5dtY/N4I3eypAFaIEu83SaG3XsfULOfVTEFaNulKdv/IF8tfnO
RUiXRJL+9qO5bCdmqyTPgtaEpggExY0RYVQ7KKPLsgf6OtnuDsk4jTw1uFkRq2dl
R9und47H8sGRSKAoboMUcM8LJLInoHvbx9ndF+NmbMMvcwKJ+1fHqAQ6IOjp05hu
pURxK2Kmu9HSEYv+65SxENZDTlUJENfv57uJNsdVBg3OKf0UX+r7F7FxpzushCPP
MVFXDK5RcwIuSn/7p5uJ1WiPebtWvu+nbaLQ5UpMHN2e7AZw2hrkm/hdpuZuJeTT
Zl0t0FbIpuLSyfmIiebE5yD3XCaq9UjqLMWq8aaBsOiOPk9g4jn4YgJT//5diUsZ
3C8n/aSvodGAJu7gD1i1yiOMnKHYozEpvhtPUlszjuuXP5CID0WoPOBsDOEhKqYx
xlge+p1woC/CW/gZ8bs7NqlbIprt1HFmtsVsHDfjMgX9VjOvpyiDlMLbBUxdp7wq
YFqb0Ersd2mdr3LZA09rfLOKJUv0ozVHBxt0m4dSonQeBgPi7sIiMtqdnQv9xcwi
XMufOglqN8G/7OL6Bs25kTD0epBJssEVrW6xuAps2SgbhNmjZ/IlVpISapTnx4Kz
xVYYkzsjRgGwT/iSHIjRGjEGUx5WH+BUO09eq0Fgp9i5tg6OBQzGTY2nMPNSFW8o
WGjyjZvhcF3kfI1zfx0cdZyhAG1APksfZy8Hd6n30pImnv5uSIu2NohSMcR4FNJH
YYKEuX0OjrnxnDFNo2y/7bAeFrX0K5V9sYOIirhv/853ZERNa7yfhcZtopBz78Hg
70X1FDQFa02lckTNeTJrC3ifxne48ULr9TvgqdAQeBtgYM2qp2MwKuViFUWM7Rx+
odkUU6FRVjr1nn/teBsxCfOaV9pe+VG5lK9kvNtqssQjknzHLeq0RwaFyRZl9ZGQ
JCUP3el7TSOB+UJBtKSttZTam62IukjAXploRudg8NIsEzMCasbPcXTK0f3P7UqP
kEabnJ6pHzT73LZVdvp9MUpuUf2BrG0VFYKBbGEWnhhqkmsmXY3a/nZcKP0d+7jx
EqChxSXBt7QSyn0/Y5X7KHWo8QHM4xDknQXieVIVgmUXzDUY22nVoH5hfvbsR2lH
RMTLoZGZvyf+dEB8mP86DUBsxLVMaMAJedtXclCv7FbPO8Gs27qPjoMWDBt/slFZ
v1MuS4i7KOAaWmr0p+JpEb5BiO2/ASqVZaBlhz1pQel1Hu+tT0MkPesubK/5IjGv
lR1jbPyNNBIetDvh113HF8RBMyJ7VLItWTnY/bmA/jdqr7TNlNiZ5QhJY+mx0Bzq
D8dyLHTk4mCT4owSBExXwyz7ZA1zp7jK8z7r9Td2BozZbXUvNNj84KYNBL0muG+M
SSv/t6WMjBneTnWwqzrDmsIz03k01DBgCKMrnWaBQbIj7sd+6+tXXKOWYq7cIkm8
C7LunXFjvOGsi683vqFaE70Hha3Lc7VjKobRlQ86A70z54QA42Le1F0bMvRYLb0M
tjcolyPLvuAFfPjf//A5j64cmmmlQgtYhw6PeDojHpmYzhyOkYReFiR6bJD60Hm5
qiQv4oEdR7YipyirNnf6VxAwx6q6UrT/WU/J0XxsTVMX77SOtEDo75qU+XmFjf3u
q2rjPgAL7dQnRL1jqUzls7OTkryH2BPOWxMlz2QTYqSqzyKh5+naiC/8GXbBmJzH
FbfI6u05vJAxYrLa71tmJecp9RCwZUbsWC+S1wVfDoB9uMLtyXqVqCiCBWeoWu1Y
Hfc2NF2xU4QHoqoueBpBMmbJnGBN+qrze2JFStwf2KFAVZikn2VNFvcZB+1kdWH5
r0OyQaaAYeDi28zWpV+gJFRjSPN+k9cvcQwBsfcOrw+PO+wOGDi0kZuSMVPc5x0Z
V6aYS++ud7AnseJWYHwEQTx4qBJBV0B2yceWZX4ACHxGzRomUKCsK1MKDVyl6KAY
umJtG2yGMVdQqmZ7cXSLIDHrW/jA1GgZL0u3TYEmYjhRtG0Lj/edS9KcWAmnS8s0
BOdI3XFH36FQjA/ltcc6D6OEDXclMtntJra1EaHVSuoi2rxrbXV0k1TiTW4akfUH
r2/RnEZClgOgNvPoKGsKqbg4SitnGDV+xVnQvgs6tQgDKpj9TMWm2EBliCJmvDan
MNxZb4S0SG0CL901/tFvx+r/2khYuMXs2PeT7osD4zbBYFkWJwLS3g2FrA5slS18
PjnFF8ghy6KNGLtx93BYxwxNMwIlrTDgwKQtDwKXUNMrtMgtd5XSGPDSfYL8XJmK
m85PVHwC/Pmr8IgsU35KK3eEhTbhfTdZbIlCnxpubaE3bBBQNzMnYiZX/opuQegU
MSZlLnGfCMO3oAYDonpgPPB0lVuTleduz5vx1+baX5rpTckaTo+K+MYRq4BUH5g9
Aj87n5wP656xhFdGpt+0R3HGJYIGJC6d9w9wwZBl460pxyZTiSTPRFLdMO5lQ1qE
225KKTUxnidKKIt8uO87KoglPr2Zr6D7Re2ZL3PAHdfTC5/uTMm2biFPPYErzq0q
FRsZwXeF9phFsitFmK+UyHg6yBwNWlohOkxqw+BE+uQKH76B52Ov3VxfOV0EvhkK
lUFxPlyKxgPpNCxixMGINIqqesyjlKemqW6sqpqjPx8AxjJpIhF1u77Q66Q523ky
hj6B84NaxuKslaW8HIKh19lWN25tq0WSpRt/zQudVINBii2n3RSU1h8+LJzCsWxn
j6U3LjCsJv6b7e4hna8SWvZEt7imci+cGbOUHZ6L6PWY3wSZBIt3ov8MUwsCnYXS
Vx9V/u/rHLKkYWi+T54nq7NQ0Z0Hame4ZZh+eFmJkI+OqrFH6bG+yU5scTmr6/ET
JAZ+XNaPnyy0aDCJ0nRgIgybcibm4QMScgLVEKavK9gvGLI1gSXxj/iiLniNJOW+
X126osqM2B2uZ6WbZM1W/6rymkcutll0a2Mp9rCHXmxECLnj8HnQETSgc7ydXYJR
PC3Zfjmpwk6+OiJl66hZkDAs1wDqi7/v8R0C9uKpj/qLuSv80Nc656tyChaXA2vY
mnmyCHgEaTgzrCvin58Vvsl0+Z03PoAIgpUqW65IQ8gVxwaQNQ1ccL4qNBKtHCxH
f6wLzh5yERBklub0+VWOdcVBQ14NPh2+KFGyO1fcZ4oKyhueNms2lsqLmQe4MRLZ
EPmld90UmDS4+WeS6it0UxrrJC/KeKo4oOxDFFzjNR5/8OKwCNZf8a+RlgoJjD1w
KHWCckMzvwOKN/GGfBLxhIvct3nxMVgaeLVJl4a70f6fSPrEfl4dKqTn0cUu/r+s
tSBQFRbiE6zuO5VDOXWUM5Lgeieph4BsAbsRe+DIrwu72mhawbXPKMuwNyT4Gs0T
FJCr94Ip7QwEspdpXwPetAbUsYj6x07Ex8metigypPUczV60KD1yimVG+cC9N3h/
d+3Qi480Ngkk9EMMw2aQuZIcAQhsvYzw7yAWiPggqDty1bOz9YIbzA7o0eKVS09M
2N51JT+kyshUHX2P1Gk7fE6aWqKbJDRglqNnKglDRJ0/vXxsvAGP4Ptcvk+B73vs
lSE5ae+ctCf/AENyfoZ6+MfdSGvEKrlkzR0JO76YwuZep1zq2JGywc/xHWaOECSu
jQ2aKy72oawbLwWphTR6O3pyVfj9oTCz03C4AgFwFUgHkGumpNiwoHtTdQv+9v2E
wnVwhP525e3jIv6LnFCSCe0kY0r6PVTYvDvQ85nkTXBLlQIv2mNAZb4Yom1sAP81
TIVl/DjWbcEdNTUz8YWUDaSASNeSpx/oV6Q5xT0xi2Ga4oeIQpjqG5zGCjuMkmqc
X8TfiZF8wJRRhW2SNcvv4vq7cn4jXrzSkXStm3fsoucPjhcPMWfGPUMAGJgXAzmZ
UW4ywn1WPjUqLF3X96Z/pUa2BljVIWYqub/fWY47DVT1VxdaOMJZxLgonO7QUv/d
nI0x1owP5Y1s9E0cQxefr00ymbdkHie6vnLhQ95ai0KgNmj6qQZjfhxNv+pC6G/5
XWdbolEMgqsyxv9xBtn17BLPqDcoXFIEv57zP0TYUxsJBlWaw7jRlTo1/oOIBheZ
1gaqjEL/wVQK+i6/qRulX3d3FRjK+TysDJhBVxSrg74q6uPbFVwpCbfD7cu2PRZl
q/CDkgEevSRXYawueZKtxkq3xWNcLv+E5pjknliNK8zFBdHXD4I4uToRzGqiCLl4
lXWmUsn9mvGF/N1QxAe8/kzZ/wQXTMZa5VCz9AP8Lp2A2ErTVho1/CzxnpQ1ESvQ
jjw4zJYQbiSeCstXM1CQMeSLe1fhOgC4IblVjzdlmwJxE0WZY29kdSxu9fSG4rFt
1upGI4TkxKXkvYe6TG3um6/Hw3jgY+O2yc5bDnvD3fGvw7ZAiF0rQOTz5HPttleZ
zJsn88kzpobEIFjmp0l+GAo9ynhk7i+rQzfAhwC4lbUatqw+0ZnYg+WnFoLuaYWH
FoaGiTbOszBHUxVOJJood3z8SP3QqnNiYowIG8qimxc=
`protect END_PROTECTED
