`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9foBeoZB0YjXN4XpxI86d33TpUOxPXSUd/mK8tMl8IsZxWeMRRebB8HWI7uyvi4F
fYaDTIHVQNStzdXdjXw5CcIF6wU+r7PMNH2sgEnfrwwgcyU4CJTMczKMLyQpGgxe
xzpzY6QrrsLaThvKDbH2qGaUGvFNZbj2G1hAy2dejRGZnPkgSktY0v8+9X+ExEcM
2sgdiNyK6bmo40ZDGpBvuc8Hjj3IsGIEX9mTUONXfkd7HSiddBqUf5muP0P6swin
n05hwlM8bFqokjr2OOHqufQxWFg8qQcE2HxvdMVr6rp1ToBsCV2Jn5tyEdCS/pFv
HBnbIO5NY1KfkFPMWe3UeRTjmNYI6W6ozBtS0X1UUOMIrpf7cRShTv/Y5+uBA5CS
KjmEoWzOSSKl8tcajb9i1LNuiWuTKr5uM9Fryv/sMMsMmpEF0pIpZMnLbJSMNWod
nf2tZb2/qGBrUyYiwECrhil7I4FSR5bTRfgAF5Lq7wF/niNYi5kekzRP3syM9UGJ
TIYk15uAgiqslzZcmMb46KZ0aiC0L8Xzc+XFooL4JYn+UlokhqWc9D0x2Runn6F8
YmKSq3zXhhu6BS4j1Dtn4TLE2taGK5VA84IB+CYCajZ7iQbqvYYjarU4vveOodmb
tAUnOxEV+4Ve7MFPAmcgoq0fQUWVJ6IFYa2c1ED/UsTSPIVDrslncaPVT7a6bPqD
yShVbwHwQJlTJnz4XoA6rIphp3VYeEd2ZYFcgtyqUHVITySXtKODBAPSEIuVqi4o
oqFYPtFebWe4+TIvcvMftk+KhONTwZ20oBz8yRoMiPT1NiGC55wqnDuzvKuGniJs
qKxT8sbXUS7RvKwOEl0MB4Skg7LBhBTLLqXbLQkI8JEYwY416cxstXAeFZpYj40X
SWVQ3Z8D0FyySsTTQhrYDwoBl3pB7gvzwLuPQZt8RRuqh246p0xWAdsHp64v9fFZ
AxSYM+wNZUCkNhRGjN0VOzmlek5TpGKVzrJGhUWmXdZRoXJOxAI+zWqiYgrug1lZ
TX2c4+r+BdSKsNXMj6SRJRogClqn7nAYuc1jujXIwHijhuEE9gLMScAQJOsWiB0n
VqJO8lX1QG7L+9RHoCWnSKoHNgGntzSQiXqFDh+i21TqEb+UWYX3m8i5+nkrVFNG
apny5FPOAlYU2O515oESjH/tW6eXlbTaqv5J7JOqKljCSNb9BZi8ifTOr5u/88rR
Lj745dOsve5lDqw+tPw1R6YutP97pPN3Qo2KXtEKfGUf59ltPhSN8810DyiDrPMT
MlO4EeoQ+jv1WsrAveUVIhcLF2uxBYcjvh0U9tTYWhbA665GnRB9KjTu9S2TUoYR
H5Bob7CmUruaInAYg+nOsBtcdoDVPFHJQeBOnHgKi5FhrhoFgGwaLDidlMqfx4bL
Kmuqk44aAzXnTHUWhgvl2hsauN4D7NFEb+nD+/JNAzU9H/fT0v+GDFV/KwKDw6nf
4p5RATJXYvMN1v29MswvJtAFUM4uylYNjSUew3yVwYVRJ7UjZQhpeVoxIRepzWT0
bfUp1VzieRN4ugmtReh3lOk7qDKa72kVk6MJM6taLXkAf1zD6fFQneojDWHnAdku
Sep9kBsRlGq9iO/VPb0Ya9Kx/m4qdF7yJl3Y66zFKZ6ciW9QVSdbR+3FWfdzAcE3
VFF+XHMksRXAmKdLDAxAYk7ZmB2pyjVaCumYXiA3fWdjkgU6xB7sYzDVK0xraKoA
lN6WfzF6a5vqzUFu1zuuCctSYyAvw2TorF04/NCW8/QhSCPisAuCrETq6q7PPIKc
`protect END_PROTECTED
