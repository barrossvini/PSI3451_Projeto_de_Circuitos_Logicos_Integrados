`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3rqpCJG7p4ddDYq2Wq2HeWOX3rwIstRVrPYrhKZlwuZIU71N+ihJ1TCvkEg7t0A
ot8WLCJYyU2/m6O7lCKhczts436c+43HSqJX0GOwiR0Kjc0jiGAAImLJFL8PjM0o
Rt18rsOpujFgWWuVEKTv++02Zsdkn7FuiCCKnhJOtjTgBNH6aTqiXjVrXLj2/GUq
51MWvmRs0th0I1rkhFFfa9H6hqTHo/U5VU/FEJT6LpUHNCGH8OuDi0VjNQFDuXkc
nAxPaLe7av8PkjxI83q3Fovnw/9Rrwdgk77vQLD3iMd4/ofDg99i4xIg5cxax5K6
TNV7eUIURgb7UwtE2lN3AqA6twlzo9bD9KlVpoO4cgZ7iaaBEN5PK5cBia4gl9Ub
WMAJ6h+25Az6wGkOT2OVwtGvAupT3sA4uiAsvcoK8rBuBH15Aw7iveZG1gN+u/E0
TMH8AsKq7dmK0KBzPbj9vZVekQh6PThPclHkTpFmmH5FdWdleUMj1c56DeESDXap
ChwKShrUJfAvYurG4GcGrQWXZc/RNCP3LbovS3eKO6OqUvc/WcOmhg1eeOKlJ76A
7mRlRfwL9AIs0xDj32TyZ1o6mNxA62pBg90EEqK3TWaFVfdOiWovvYKWIr+w++o8
ORfbDKemgY/4skkgNdHkLroyhtBwaqSLQmqqbleeXSTxilu+3uwH+JJ1hJyeBKae
`protect END_PROTECTED
