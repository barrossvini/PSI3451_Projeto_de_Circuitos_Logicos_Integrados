`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bSQTfTzYQ+5DJtOEXSrWKtUG3f9zEsYrLp34ceH0h+3ppc5Ql+yWsCkv4UHCaCsk
kyXsm9SbTpYP5xGgg1puL41zVTPlaKSFQq+L9HtqsP9Lq51VO+tSf65n9hQaNIDe
B8VFXdCY3e9r7KjLUOjdLnHSJHwQsWtCv6/1+YVo/BOkTvvbQVGwo+rWKAAJMf60
xl9yiK8hGBX5yvnsSGyCvgsGGnRyKr39e/hSpdAh8Ov9dxbVjLKvdcTvEYBYcYDX
9/6v3Hir1AApKNZoXRDMEVgQXrqMBxcwvm+fr0LskoXIVkXo/14o04WXcWh83xVQ
PeuxaozXOOA4VHUhswLKKhxJ7eGZYBW+Cvalbndrz4NbOn3vDOEu+fOXR4NavLRP
iWBi7NVGrvCpMiVt2yncZ0HwdeQhgL8gXnBOTmAFLmuf8Q/9om67KfEl/ts+RimM
NxEUOdVm6gV18gU5WIR68YsY8rxwTVa1pncowuq/MBNyQ9amcfY8LZJ8Jl/QJmq+
cRhS+19kvDmyz0kam7XIoFr2N9I07wYrtUOT+Emjcixd4y9SA+V2zcLFxRAtaShT
FxN89UXBYRM8T5p3d50v4WUCxkpo0xhzmsKPXfXCjkQAuWYRjvy9fYTIg/3JmVw2
RZTi/nPJNjMsLO9v1a5pR8eixpRVsE+yPRJsDHSzS5XGOj2sUv6lKupnWIev7Hwa
hni2DKhzw45ngygYlBoTQLaiRkhRzDwvD4b9ZylXtShMLjj4aLR8SBxKnxa7hFPU
Gv55rfabZN9KWBYX+w2PUa4YCGFxJyWoWeT0+6j8QLs4s7K8SG1fBqL5+dqixGGJ
dR5sT2qOvExA0uVVjo8H/vM+2mg2/oRYHm0VMyL4LnwSiQyRnTJ9h3fjvrJYWkdK
sS7oRguw4fzt7awAkZ+giaaEt5N+GbvnM68v7K9FHkRnagTTpyav0HZP1XVSkM6S
+kObHpb80+ub0H/BsY0eXCDKDsPQ8EpOoHRT7sRfNQZ/RryDfplQVLQZZM9DJs4g
UeQ0kjVnpDIBEs6mSdorKFT98f5JTSKsBY9eMrO/Y+yGVyUgkZQZUdFzIeJodqsA
a6zz0Taz/oUhZtZovlfGXNu81kJJuSkDu3jaDypaqta5Vr8dgGcPlFRYknVsz6Vq
FE17SuyFXQMkphJpENFQ0wULQEyMEh4en7snLcUAHJ/VdXnHp38X3uLu/gI2Hodf
Jr+mDJJJ808fieCWTW164tDi1FiKLLJuRIYkmiWGHUHFQEvG5y0y5SH0sS29T4ZU
YMFj3DsFk4el62r++SMVNPJYRrvLv/yb0rOW7dMYay/5kGsBaUkeg7KlUEpH8b0F
2UkLNOUgu88PksoKEehgYs3qzqGx/SrXWC3bJD+UmpZRJh0P4JltlMGMMz7e0wgU
qCaxZfh8bxRVsdQ0e67U0nSZ6KOAFjBTH0KEpcLGDI/PCfpq+kmTPC1iRA1NtWCD
gjdvKIi6mVz4/zm7DCtSH+M7CVmWehZ2knpHa1Il1pbw4rJgq+/z05sv0XXtV2gm
yf+esGC5isevI9ThYSe9V1oCV3kkZcpGJxgLudHtlubZQ1ifr9lkf+KBo6tx8yEV
2WPxNWn7NIFDgqlOctqUP1FJaLavcpjKBfgIAVSIKkE0epr+FOv9PaIA6wsv2J6t
FRCxefwh5t+s1EmNaPIGTdgYsgnCM1+/TMNFplnKj4BJqZoc92Mu/Fk2S7Ed0vp+
9K1ZOMEN2Tjt7/z5Qfn3hp4RfZoGb9bCMxxJOnL4d+MuwvrEZD24FshSbIulzmC2
jx4PNipOQxe5OEAjn+1DGvBptVKiEJIIExn6fxeFKKx+AFMFBhANoovNjbDmYB7w
4D6aMdPAKrzfEaQ6YlRrnF/PjN+xoI0NLZkis3gA9gVz77uOgA2FZzQy2BjYm2xD
Z8KwsJ801UVmVnX1arJeFWhP6JsvjVRaxw5pSEMcMfvAFBReVIhmHBPjCfdyIgkJ
Sc0mZSIJ4FdVM9PA5e+zy08J9bKj7Fy7ZY0+YLJBGFtUt5oZmItWrILgj2JsG8fB
CHT5K0T4BNT4kqiqDOG73AHm6uh12illD6OvKxAQeXSoHCmTJuFsVFns5kVu9+7m
G0lekNh0JHD3nD6orTIptDKpeOQBuGVRu16ZZgw+OHrTHqCfUDN1mo+b5gQ69s53
NjMU60kUeRoOuDOWyRWtNSLUZFDQnzU07DKO/qZCy0DDuVYC+BsRtHPIdTAvjYrq
Uh8PPAeCLQQELCraF0tZMNqay4JTnwNO2Ni4aq2GExCChY247QAPHFG56UIcea+s
Ed7JVj2OQ3z2z6NQI45ebEaKZTYYVMI9KTnVerFNTA9oIjU4jVmPVf5aLUtXpEnP
KTq2EPDvgebFW1RAQLCEDDbPxlTQAgz2xXnze8uDF3v1sfKIOyWkHWHI9S2nf1IH
+pOh6rJbOorBdRhIF2YIodNqgoP6lmRXENgCaad1GEWFfvuUXRV80YbpsTMbsOL5
wPm4EL07Ip3YW6aOSWVSGQ==
`protect END_PROTECTED
