`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NHwZ+99wN6Wa9oyJLXbHeLCeDe3N+FV/U/wX14GnjNsvoL5DTN3U/aJP63WELRwT
Bh3vc6QrUK47lFQF5yvv1WNVpy6ojZqYntFvHgG17186US3OoFGfOVPKWxgrENCh
lOEA4wNt50ykq3nW8DeD3HT5OdlrA+NLpgGCGe+RlDwA45+rJNYmtPIxzV+tN4FE
Fau54DEoqI7bzfIZcoT5A1IcKnRxvr3x5LtNKFvEIRHWJ37R45WXI8fpefhIQHuF
oLZUhIahQLLOsNZBp3RQX3KwB7R+iOGx/pGhyIivvuKiNXrcvgQzVDsXipoxbMAv
vVi22qqc14WPq1iINJcCu6pwkwpNWbsbNl2LBjk2BQWR5f3o0AHRjXE6ddu5KT7e
9L+h9YJMb+o3qUhcD8/YFaWAFiBVD/bUOueYlRoHKMS7yFof+qE+q34VpkTYkPaU
kTDQI3soGY57zO6FfMZUZg==
`protect END_PROTECTED
