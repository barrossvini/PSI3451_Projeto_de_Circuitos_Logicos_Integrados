`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W6wG4RYBwnE39CKY8EO43x+KtMjuKv6TFgIeke3uILtXhwYtQ/axn6sB2UbAbkFX
McYlBYmqs5vT5P0jdJVr7t/4vXBcwfwyMN2ZXwntP9TLxqPKGPDP5gVcIpV0Pi6g
MDmLt/SbGVoWv5TOzXiFUuUnKl2eS8j948/xOu42ss+vutC9d+t+76Lsyw+NaSOs
rOiXzxU7ddH/vmKN0FrMuUvGWligw4+rCG2ExUNyIeqIBRnqhuUh9aEAt0lRJt7v
I3QD+9VyejdLfE3mEFLy0bjL2NxulEvd/wZqOGbbLogebOSovJdkZLNqTOkfgF4U
b8qgQedfeb4d/WYKThLQsiptiCtXZ2uhWmWcQCzgSdkIO/SqAPhSO8utodEmyB2h
tosAiuWT3NKBNBEtPKOp/1fRYGVMLVF+89+/WKI2X051nykmlFqPtm29lYpWauWb
cFKN/5HAJc1IcrLcU3UELtFzrG7k0Metnv+sEGXFyx2ty12Y0WIQxbg2BPr82muF
7qdZzgBDo2xHso3hE4mkdNdKkCOrFlRaD88+LQQeJUYmZtwI3pIrp9INF97bUclE
ULmnGIBG4KpPzNWv9kh5YUJGooVWJOE31SHuUQ7AZlq0/PT0Sb/bEd82t3evyFtB
cLc0x24jo7wzpnanO0uCGdumzBJUWrHLVeeWJZ8xvAlJlqekOeC9dk/gmV3Xm1uP
b5toFiSc2DAqcRJ8u11IJkBSudNyTV+wHpF+3B3lFjMNGPNLFx0U4TO5ZZPpmdkj
5zVWwZPkZd7TgDJJD1wDAw==
`protect END_PROTECTED
