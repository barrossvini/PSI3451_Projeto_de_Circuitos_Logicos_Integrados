`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fY4sMQHzaDQpONsQ0WHYhPgEa+E6txjt9Rr0tSrGlmHW7DsOZKpmvakYCfbD2Gsi
1FlMnjYZhy20vFeI1HAz7CoIfwFwopx7mmv2cPvNVIsLcE9hKRrOeGZtdGnMQXH0
xEbm5R4r4zC26A1w8W/4QIBLBQ395DHIq6719gBKlEasvA0+DXQVy6blykTo7lMT
24LCCyPdpLN0mWmErim8nn8C81oUI1RAAc4Yhk3o09CV+wWMqS5QKkgth5oV0ilN
nYoXGUUibgTH7qefqBQ7//40ZtV6155T68mhyHH72n+Ye57Kxax1Rx6+UR2yqn13
ApwMz9viQoeaqSFLfaM0mBaw6GOBX5VChYJFMNGGrGT/4NHGj2l/6YsDCaeVlp9N
8MTYQC9YVujvQ85+3zvJO2mywuKozbuznj/wFDUWAC7IiHGZXoDs5+BDoQzxi1HT
TLN8HtXBbWaBZXazCwRWPGCErLDaWijqoQ0LjCa2V+U6O+4IZrJaXLqrJUTlgvNe
GKSVt3bjF1tKvvwdIIHEcBMHVd8cclWaAojBhVKGiMtoXiTBmpTUz1U/W4vPHJno
6ICeKoU5/z64qDKOVrS99Z3KXSd5BSl+BEGsMhJu0i476F/zkyyYDctKgU8HkI+C
un3nrvAxGlb8zksY9mkyvc3nXuqRmq3W9fJjTTIds/gix44MuPcfKo/5B9rFqbv8
kOP9NwilkN6N6oU0c1PLQOEpP/uIfMnMJXn/mtENXCRE/jA0XloRqoH7gcERQ591
61rsqteYvw5LORJeJwoaeqz8knTc5UNuaTp2VGkDvQtCjpEz3zLSaE0tYKhaeVEw
EE6nOKUlxkZ0Ypf4cPJCf9qoJsJaLJSUW5AWYT76/U6L2LuxxH0SmgmL0aQXF+S5
vGgiiLKf0q14a4YOw+GnJ19P6YHB0Zc8dFpkQZd6epZKeXlvmj7IByjgZ16zMTgj
rpHb/vTLkm3kquS7Y531TGrHh46DbT2eqKRgqLm45f5kiqRK/GIgR6VllNxrIq0k
5KNPLteVTaQW9D5Z7wIdnH2Y1h+j0oiyHVLu2V11BT/X7WFaqEKaY8Yaal7cvgvH
BcHK4Y0zHmcaLRg4eTPbpi8PZjNvar6OUwiWWHCkuWvRr9swY95rLiq9wKVNHCvP
LPkjbwGgzzgyTR6i+VzkIzRqW4B55I+dPo6HD+XpzkgO/O3G0iS4MFqUkCvkhxJI
YlVCcW3I5nCTZ/OubP5OXkMSJ98rg1bRnKKyrR3WXvpKbGM54SksHl1SKhXrXako
qanhTGLKU69OODqDUaMn3UdPZZXnQuaoUkjZvRUbsiqAOUTopokDWU6ExOQdtnJf
z0kaaNRnxipXcQXYHMGl7WDP4sn/PV/cbsrDk9wlbp3oGSYG/t1Vp69fAo9yvG1X
ihT2J5DK/gespKJv0kzjXY6NsE99CasEZ2cpnmPvFqDdFFaKAs27FbUo5RBFy8cf
0O0PxR61fd89PzFnEaYX6G7qQW1HSbqz6/WColteDpGC5bd8tY9BKOkjOFf2rpbg
k8oYVsBOSQxD6CLFo6RpDgtByYbiHQ+MymLHcSvSxY/2J4Zh2aGVYg/xexZhcHw0
QNosvbDWNSR6i/Lf8RdUd6xGESMNAqV3yh8pdtEdH9JVeEMJs+tYFHMcHBFzsVTk
9lOgFIVD6+a6jH1vnQYdZD+/QaIy5bNXUHAc1ebWfcxCfL03Gl8BVIJWVeNVcIZh
L98rdm9P4CeYkvydRnAVQRMv//9gFQ4MhrPsDTaXwl5dzRiyhMg9zqqYuLeMdCmJ
kk6KC4+1dF1vO5WG0iPatk6pOvzNaaXI1yEu2JalPMMP5THvXAPwWMdU+mGt1ikA
rwyL4oD75LSU9lknOB1IoDk7/8T8fRJ3JOYfr5DW++es3FsgBpbZxjHH26gcQoaB
+s00i65nSBFwUFXrkW10/29NA7Plh9oANGjC26ZPv3ZHrbIqGCpbQzBRyouZolw8
wsagm8ElTHPTQjyr86WLW62ZUcQEtWevN1MjbbPXCQSIz+DREilWOg2jkCNIgXhR
cd26IpXHhv3LAbDQVdvl45uohbqwxAgoMo/ugmOBjACCGrAlDTwpho3EIAM0EZ4u
uyHGwTY0By/hTan6jzRIdplwTRdXcZfjjfJHUBF98wovaQ1SnefF/h+dMl+HCUC3
hJDnvXvPxzZaPAPbfuaDHtjc+67FjYv/7cLvoTaJftxprHbilRemR8iwJQdmlXty
zBToVTQz3BMLUNLNhFvIJw3Fq0pO1WjGM5a1C95snGrSiaZW3tQGBz9s7mb/otcJ
dxBowpiPj7Nk5VWU1RfFFyS05wF/jMEgfSRxWyq2QxGWf2OR4b3h27p40er2Uomn
2xWE/YGr24FqT6dMihjcpj2MZBQQ/zNtG5zHdEuvDtKXuxcgq4gYeC/bEjMOEStd
YL3qflkhy16qPe+xkoIsuWSI2TIjzoMofciWYySg+UTinW5DAyQlQ+cJNSkc3qMu
cEFG1A2T/0HX9jBk0RpsknRhK7bAiJoEGY7T5jmSwoMl7Pxis9ZOvLIfokkjTL/u
5doYv49KbnGj2yHdHEhyKl+dnNYkQIUXf7qyJ6bs99jmHPdQ2cT33WAFV2E0EVXj
ENLoTf20ogBohEGuVc2jdeeyioGPhwavnDjQiE59gRCVtuCb2BDTWXVmhMu3l4kw
ZWOpXwKZaArJFDGOoF8ZMGojRTVKE3S0z1ZKtfCWIarXNQHGldw6MBrhW7qshDkO
bGBwLrODs0ZK2dT67cLGow+24tns+L/36QYe9k9qpmmfT5vrQLkenLMaD1zaceep
41J/0HQHN6ZEJ5sUQScKkbQHtweifGvJnIAZfvjJsDJPdmqZ/Kf+88Rz5s/q6a7f
6oPUg0TU8XvMYWGtrX8HfiTYx3RZjmuEvKDXj+/1rEF2DhQY+J5Wk7Bn2LvXWmi1
vsM6kMNKSDEYfxZV9fe5g2CSvRFMDAj2t+dZS47R9tz78+6oENeol72cmba8doIh
06kh7Vbj9zFsxd2+urLrLvdT/FQ6Gkmu5BoGuz5oI0poXz0dyJj33+uzgFzWOv3j
IN3awDR8lwu3y/R7YFpSnKFcWzs0utWiC4HOQzuFheA2TQHIOnW/fvlrC31ogPHe
aviNjt+IfGmuG6+1aZNok9sj4de3sYXmSL6hRj6sNx9X1ZpY6doUgipjQKMNNlg4
fVCsBE2h0VcLgdQrElbOl3+pBc4zCoSR5FvRvqM8CNewIr4MtY5hPjxycIUE98a9
lcchVvFZ29zHq/ZTQSZDum95HOoVAjaaEUrVy9g97AiPPmTEHAF70/+yI4SLvrYX
OEVxMKiwoFBG1DhoR92pmg==
`protect END_PROTECTED
