`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WcC91ySA2DzBWDoQHUPhqVwkYwCnCV+SPC9Ci5WVHwKoIBBqFvJJG6k0i8zGJFIV
4MkILl1iMuyv4Dk4YmMch3hrnMv5fCa56rjZJ/aG0kNMnfYDmRGWhBlMkiTff2OM
oPpRsF1pvPxOygyr00SfyGZD8CxVFa7iiKru6vGMdG0dMIsoHpFh1l6KSgbiDSGz
UgDyQj0eN9uumC1HrwKMoYsa7jasszQcSY0lonoinI8it2hSPqh8q2xyZJCGKoT8
NSdESEdTwB11W+OQ2jiwOF37iIJXC/4Abatmcx7IKeImdoQH0cUO34rLlCd59dHB
rYiPWkBDk5htKnry8mRZKpVbA/viNBAL4iCESta1iahxwC2iNHGBW1+mX/Pp0dCX
0SPxsYivyAyqnWn7RvZMprezWSHfHonU7iiAX41hZ8zGfu88dJhfQzh5+49ihQD9
VEYAUgX4V/atchbqEGoM0AQJRBfeyRWOXY0460I7tnDe5YMGg2xMunKgUHLsJduU
xRs3+nNnfUeifm9zHbwaxHSKPxcK+UVHOruybdB5ykns6nWBSoWomcJ2lLbrVgTS
l1Z8ON4LoQgYp9Jb8R/Z20YuynYLheKAZN1QKOGI5G9me5aHvnIeumZYhWoZAJB1
XbO1PZlK52KjezWqz4WsYKkX6YzgRhMR/f0ceryanOS0Unm740rbxNvS8vumwVoS
cIguU+j5ClpDhEiwED/4sipm/w/uH8u0KOAQYckX7BvaqY1KWKAg9+IC81PI3kyE
5VKMv+7I3f4eoTjzbpi5qOpFoMuJIDx5MLRICRMwJ+FKtFhRpbU7yl3um/tnXsCx
+tXzgXJ9PtQrSIlN8HR2T5qzCn9jWmKYcv95w3jcMiCv7SKhkUE1fhRKfOl10wg4
lt4AWHc+ElB2tcc/7AbmeJ5jEjqR1ZVCtpx6MkX90I4=
`protect END_PROTECTED
