`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6N1RHUYAvWc5zxyzZRpATF1lps/4ilnwG26664z8TW8ndXVUZUFZQk/N5Vztk/AG
/u/3lu6cPjicCSJKu2/yCJB1AmGFNlMpaay0uN6OQ7wtGWbbhDTKaGICHPz9toFI
V8IjqH2E6usM3DUBLkQZCvVBRqHdujv8p3dU7u+vjjHRNTiz+VEGWAL/FndlRCkW
sD/XM34XG+L1Eu1uJgPdoOhUZjjs06CwGKCUcSMDA5w914sXHiECPszQxFALrxpg
vKqzeL1pZ6D8VYmdM5zZ03/GYTaGE1xSDtm/0KV9YIZvc8UxBTwTgrmCyyTrB7Sy
Wj23LEYYK3tL4//tt3sNMMEbLzpW2wzfYU3ciGshyWxlVY+FKF+EvRY4MiumzjTV
ESQbWDcItE5vaUCMzFfkvdIwZQMdeCOoNjUx10+fuqNdWZ6VgTBw8c3uHv9osKV7
OMfwJbZRcW4rWgQ2Wd00zRq5D4r7seVMW+zsYphA6fOGJZp+jqvi2VcT3OD/0WjF
TOw3jzRyy0EDVeujaM1dO5K9Co9faABwA+SZ9CUB9+o=
`protect END_PROTECTED
