`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5bu7v6H5TKSXekyD1zIAJg9kJXTrrIsV3omMkR8MnMspUxdvk9WHkNhLTgAPWNV
DYRlq1VhTFiT1Yzkm6+0K6utFRaIZ3gde2mieAmnk94YeJpSliLYHwzUSav45sOn
q0YB0/j/TPweXi9x+IdpB0TgvYUyx9uEgwEhraU6A4/Eoq1KkaRDKRx0h7LFPy59
kIz3iGDZ/n3t7gv63H97VGKKydv4P2PucGk2FkM4d226OKBl/vw/440xhYpXvkKs
9cGhV3i0khfVDjKmoHHFepBE5t6/DSlwRrtEar+2ejarvVmkbe+o/B+WIRtwnTYA
kkGdYF2k9c4PWpAVbMIAUAkcaJ1ODHa21bU5V4iQx37V2dtt7+cclIIv6DU7vgGZ
LiUCe3T4bq8Lx3v9TEdpTUjfxPIHUI8breXr8YYhL29HIitmPGWN79uLQ43Mu1Xm
EgyoFdUTSaQPj0QispwQfcfsPq6tivRok/V6rXgqfUXQkQzq8uEvxD95bcbAU4Me
lpszs5Oao8EzvauM/xpRsU70Xmmkyu5wjEEkfYnOwJOpVCi1WD9vClYgVPYLt4IK
hBP8jVcFiDvYM+omGOkmN/uRCc1ctqzSDqYeMgRzAzbkTpeUJSNGGna/AqdFQsBJ
zt4PRIS8zeQiAzXWOVJDkhM3ZHkxDDNrQzqhmWzyrxRpHwIJ4SJyYGXaxWamQ3Xj
hkG9GeFddn7yokCQi/mrdGu4kEiQ06v6f+GHWeq8585dksZCyyMl9XNkIXfx9I9H
oQhEaCJsqnv6E1UT8xUGI8tUKLoi4HLmuz0ubpLnajtkVWj6irmsN69usQE2ZVHF
fujyBIsrfwXPjSZSd8QAxYhdcZ7ui2w1FfRdKN+you2fjEjOp5LIizPQviTFVLnv
QvQWf8bgIBzc/5Gsc/0ozBR9aS6MTwhog5FTpkLdJQWty2RpDKFwortagSFECAbv
Nb/YuoSyBPMfkq1f/f3fNf6kSw2igciRshYHvsbxwplA2yzVC8ZI97NICAU554Go
zJd5Kg6oWLgfD8kN/8WjOJBc1XbIg8aYaEhvWY8lWOt1brPBWZ4SxrIdsRjNtYxh
8AKSfFvcHG3ljxWuldur3C8xFKpt/VbiLETg6qz2fV27Xl7KbdMUG7okkqNy8PVC
+mNMWD4beWYlqqjnmrfnPdwzBr73IQfaK5Pspkbs7VNf2bF5+0Gso0YSm0eQlwPe
YV8pP+aIiQVpxrmWapGRo4OKZOg/KQZvQk/h7cW9Y1Dl23rwnAl9YDrSvWzClyXJ
/huocAZBo01PySjV24bvuJDQkz2Jv8jb83Yz/9wv8QB0evl31OVZgYSrAj4bsU0t
UuQvx8Oqu2hNfewVXnMF1CWevpBpRtQAQ0aH3i0l6Px8H//za9ZgKKYMubc7fjE3
fvFHpiuqHgANiEUZkxzQQpI6kGNtFSL03WyArKdv3AZ9h6E8aXjEkE6BsybRZItv
5qV7F/4qcLG1l/1LNuFyd3KCS9KL4gd5YSyJza53y7MvPn7aJvV+Hp2F08y5d7RX
c+bZrYrrEx80xLWo3rqwSHXrqJ/lac3w2k+f7hWHuiS/nnRdXU6KKrz9CKT9Okwy
0BtvoKvc1qUe+rvMnLjG80d1i52yBOOGPftmalUtCcqL9TC7wDzTeyrf3SvzPTgw
NDx1fJ81V6plnF0MtmFSE7NY8LxCD5OEtHxFY4bFEE3wdiiWS/QW9YM63++ynYgY
TCKXN3jPL62Mx2BhOAt4LT6pBxoBLUiG+0rTbWejNeLTByCN8dyP9TiAWYOdpjwT
tbX8uDMrTBVZa2z/L7pZ8YD1yV3bY+m0cUxMdI5GIxn8FsJJMuYLN8Kn6q6S+H5q
ebUKl7USwtQoJHlvjc5NIOB9IPaQo2kzSGbdK5fK63Hn28F+7ARTqiW4Sel46HaF
BUj7yz3u3hrBtBCC22PEZ7klWziRo/NJPhY5aXJX9ORguZescNT6LwHH8czUVgxb
U5JTz+ChFKLYl9sAeV+vWYo7/5CwqjffruFuZ2x9NrzQxIPmuwd0mTb/FnALmtJZ
b69FfLKSvEB0vFNUfZ/lXq1+i/Yx+pFXlFo8+ggbYgA3q2REIeETeaBhYtuSFB/C
+gFNOekv8D/PmQTenCvCcfuNBE/arLDwwS5+V8OoPXV90jDYXP9sHg9fsbs4oDQw
CsX9tu/0h21B0fsHB1A+zZPJbOqpwlzU+JbQwqcAk9NgJn3lYfOYvgI9pcko4p7S
kekcGwkaR/GUSGhlj7tUn7Jd30OyUgyvV5FwvJBhKHPiFZXbNGHWoo7bVAHQYdTx
Enux4Zx+o5r5vQFQHzC7NODxHHBlAsNknQs7sNCWlV63antrGoqmNs9APUASrIWR
X7X8dxsWLuXNljIXCtZ3VDwDAa4ZhqgIn67AeKn9wPHn9rLTnukyjSAdOGU9Py3k
j/Rf2rN6K3tjBWU07F6HbLekUAlqR0EHAoxTgQTsa4IOBZXppOyWajXzEEPErNcQ
m62xr5LfaJJElwTHyC2U8vdNJDDfagVL7wYTP5qObi644Cbv2uey/ROHpAzImVXF
`protect END_PROTECTED
