`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LlnwZ2AQH/ggNteL4Fr9Giw4jHkL0dPNL+spH5jHVg5Bd6NCS513+d6qvyE+73ue
cwgYvxHIU4raK3ViRxBUDjPjDk2ewIh/e2SigawkO6am2Prw0AuD7z6En/ra0Mv8
7UQg8LZZPRWbHyvMbxerWk6lCtjk+uvDfVGQ23vdah3KWLGf5uTOBySV2Tcc7IIu
6rXcCBmYfNPkAI+Y72d1jZB+ahw2nHnpys5wAes0rI63Wt0LTKzR75i8Tvn5CIy/
qhC932xk8iwdTPxxG3UEus2HvST2wYRm8rjTBy0dmRQ+WQy27viY1DkT+HrmMG8E
Ig+DvONl+Mr81Tj3mhGw/cPYt62UfXqB7NP9OKFOqmm3eBaQXo0FgbbHADgOiPvz
GEss2xKT7AWsHyJlBPl79Am//8XltI0DV/J7FwdxKPZLJey4rZ026BTPrcXnEugf
D5XEn/RMmIrKv/5Uc5dzPggT/W/3ywRFe7oD6ABUBPVAV+i0sdBPKZ84gj5vWL4x
biorUpGRugqgYfr1Qh8F4l9WPBfRV2OZ+ydjnp7RojZWMeI+h1fZyikZ133gK2mi
28yRqFI3H2Tx/M4hNjmtWHaUUd4kALR2mEEvEwQPUh+gSMsFq8g5qX3mYMDORUk3
obPhx9yi6FsVft/jaVkcbtM09uArUxdfOMFlvomX/Qz6kYLSGQxxDrFCMdrTR9uE
VvQQcYX2UDxlGUKLP+f53JDYt9BdRM5k43CJ7EOa9ndTaw10PXtGx39js8YI6Pkz
5ZWpV95I2rSxdk1I5vH18SnI77KdC/TOXmwSe6N38AehxUDEk6FI2aU4idBYYkXP
jfLw0v1o7Uh2Y1FxnLVXQ1D7Qt5TNFjXybWkqFV5TCqNzwpj77P83vuG99o++zN2
uV3Q5dx86mSbN2w5yP7N39dgz9zHucCuNmZfP4iiUpGnVrFl8D75a8rRnC3usOd3
yCwkoylCnjTJ0m+h/wJOimZ9K2w7HHXTnLtZrvTKKFf38unjmrk4pke/NWUvY0R6
wIAay/N3Hxe5U1DN+99ARpq15BaynK0yaBTL/QQwFi2MYYBOlkWM7PCjzXMFE7zn
MltJhTJ7nQXG6/Hw3LQ7psTb8oFkYPs/i6okme1Rw2i+8dGSvfRxEePNrQgt5P51
1ED8+NPFVBFTAMTFaRUr0wBd+i9wKvbnsNtSMVY6n1223XVxeNYYvdr9HBbllYKm
gKiAdChIfmDFIJrry/gH/SPzPSFxYiCIl/Rjh6writzugTGMLw9DzfU+Bdqm2A8W
`protect END_PROTECTED
