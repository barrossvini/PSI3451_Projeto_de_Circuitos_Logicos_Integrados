`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qGsGhkJlGYmtCoQRvDY4zNatd9Hy/7ROZ0YatDQGne20ITMma9ObMqlmWijwgL1C
OOjFzpmMPzAlPcR94Dk9p6V0rwdPXT9WBQCTFWTRkOZygrFurPxAksYB1yAaJYN8
Nt9fywhpSoDHkGefLLMMgoQJkC7x2rxKlF41XvtUK0QF1i3PSszprpDFCpq1VVyh
97S2ZsUZuGZUyP5JcWtWyHB15mDMZ/7fiVh7qkKqaO3TVh5+dPWEjwxKuGwMUvQ5
Ishvw7dPiYwK2Ta9fh/4EQZC4tdFMIgPqf+ofaMh2SKQhOtUTsRpjJdOuIgA/UCs
YjH+NF8abQSpYDZ6nYOgY7tMa0rbQIFnxBmMIfxzFURGhOCfxHSZoSVxxshMMKln
WUI2xSXWZzfedMpEgI0Rg7gd/kIVIPZYt/jzReUK6AqhQTQ9Mr8WoRwmAl75NfrC
H4HalzuZaIQN8M9oqXU4R4lIU5SC/slg8N4EMlYlUXoEwkMG3pB5uip8ETr/C2bB
Nuewy58yc9xYu1b/s0EapexGFwKDgdKO6E3vgwc4bxykwKK/lZyISBIv6Hu/YrHl
wNSUfPJWpx1SmSGjBeMj228on/Czfcx+Om0jyK5tJaaj13md4S+vFsru1+8zA0sX
+ztxwAl0i773WgvQvnhQ4khxYO8koAJELShIGaLNamj51vepZnLwL1+MqmLvnOec
LOWuxv6gyGEbe13o4rqpogWlVeEL/wZUmgMdDXmqHj7Y1rxDf+MOVbKJF4Q8Nz5x
hqcdd2hbmMk0QKxwJ7c0VA==
`protect END_PROTECTED
