`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sWClt2NqOzPSsXs7EMdt6pzD19qtDijzrEqB/hEban2BIXSPCKoe/RkBZD2x9YH5
5ic74j1wALu0GmzlSaQtCziSnDS4xjM65cCx/Rx4k4X31zgjylvmxlXsLOFwP1SW
AMslogBADm4TKekhx9rmfplfgldV70V/jKKSrRKt4iFtylk+CcIXHsyqKYDuzfuY
HAmZPh9Krmfbtcrm/xifD76bbFpKYxwbqkaO4lJ0LkmzKnw5cJyh0tfTT4Fy/c4p
D1ulq46eYhV8zActGqxvWT/4CTb2/WXhfnh9UdOAzE51wjKlHYFKnthMn9lw4XC+
37IYh3G702LRPoobq/4G5Bxt7lCW06wCj8MZdJuLK2eToC8P9itumxujByU8e45b
wyWUG1wHzhyMedvvKPTwtJZtSiHAvEmkUqnPdmINKJnbzltgXcfnLrTfCOX2qafF
e7to0da4f3tmtraHyqyRn9gda2nNSxT2qtnGukYv7Lr13sG7A7FE9IqI/YDZUfQ+
uOdHYFs6x4w46h3mK6yNll/GByeJCKdROr/F/Ww3Yigz+enmtEvxuApxgCe2525C
DPggJAef5mUGG4uA8zQFW/vsv3q6zk6Xa0VNGQK6R4rw6EkVgmn+juio4JudKSsL
/8Ukd2R+a5fi9qie2oyPqE1Zyy6d1ksmQotFDR/HIvXtyiab0sfu9Z3p01Jod+Q2
9PQgY/5O1X/Cm2jRpvV6MBDyRYWhYXw0vVeHH+4im4e5+nSG3cMSpUwbwDudrfyz
gUxjTCVmCGQu/N0PpMYrT+Capk9ahHZ2FgDiBy0XTtUJPoYfuPaJiQaLEWk0ST1+
J5d+ahtbXFLqRW3YpdPWTDYejYpT4GaVtSrzB/FMbK+K8bk7axOD7vOg3HVjYs+3
n627rbvSM6uDYJb1zocR9K5tKDyIIXqLloVvbo2DD+aAkFDGiHHpqo5UaU0jFPU7
2N2vYcZfah1ncnC3hOkf+hRlH1IMm5nCVTOowGMtvZCKQfMnU1jIG6jdB5elp1HC
zTseyysmoPWUPM/69p+O4ZwyFwu/GjNzVCuy/dcUqv1OUElMSi9OlPSPPpPztdOm
T90hRmfF6wcBlULpYtj76sErrfNF7w8/zMGBI/bULW5naIvK0m824JcHM0i1aT51
b6aNliEWaxiLNxkm0+s+gty+B5/UkidfUwhuDN0LaZ72dqeGi3I2KAt/IL0UNKwe
Rfy7e/5ZYRaWEube8GdlldsEXLlw20Eya6g2/NdXbyBgN2DtiuITVu+PNvi/5OuL
kpL+q5EjAt0iIxn8VYhurk0tkwQgSRaWG6CpuGp9G0eXPP8DGG8fivGfNJfSP1tq
ULB+Qr0kZ4a9APynm2iwvdpqBM4viNC2kH42ZMEWo2iUVph29jypEoIJS4Q5amGr
6Wveo0tfzDcENIm4Bw6AmAQVkDJ+sd4lAg4l+A0Og644OjjbnoL7T2T3938vC4vu
e+vLKRr5+8AOSRQV4ZBAvn0QRKGhVVpXRXrSVxyZnxCrEI3uXDqpLmcCggPWTu6p
U7qkjTPhxhYrsmY7jO2zb+duUJ2sG/X9gmO647TsgRCmS/2vFqlnhIpzPmDfTCdH
tNzEcYI+H046XwNykfoNS1ByUbdCxAisWqMbIpijBWtsyOGAqWO1G/1K6fNOmc77
LXNmCD2UcWIvkbSFtTnHv6AMeuriqlZ1QPqBFbrLum09PKtStAlfK8fYtlSU31ib
hYHgXRO3J06EhGeMbY3Zs1Tx4qAYavXdvR45QZbRPezi2uLI8OLeXkZQEoIoRRWj
2os81HMDHqeZa3/di8v3OggmERhpnoDEmfl/btOrRej8pNyPojzy5yYb9+49Fr2t
pzo02beP4zJfg1g4ND0LfA8He52GPrOmutYVtrwd3X1FkiS1d4nyR41AkXBm0EC2
6QH8fcona01V6MqB7LvshY8gRnnFko7hP9fFFez1kwRKRVo44YCauZd4eTGiPPsg
3BBXRWsUBFqpqhujalN36LKtJU23i2mjyta1+D2BxTq81q0llTr9qhfS8LWU+2tC
BOPUwwa1xxNIJWn1sLEuAnEUb6DkY6cTX1xfR1eZip3shj5Fl76X0GJWHZJzKAxv
N1H/EWGsYORUrFPK7YVollNSIQnZTEZzfl6vpFvZa+B6K+xkLmWFfvBvPwQHWTHI
/sBpzjGMrREa8mtUWJm7mHA7npiBNzAEOatu88V39pt6KGVlYJPjpJATxfp5Pu4w
Ww9c/J7v/CfTV+QOP/OjUMV9dTuRkdf4O5bUbLJ9TGdp7rsKyFJkMayfhYzp1ikS
1giu7i8aT8f8rPupGIAdEo//p1DFrjSl1pUxkttaOUisDb4SlNzDkGAZmvFhehSP
BLbsfhPSrw4rq3h04rVbMW93DbVWamg4Y+7U1cKA3qFyCLxJqs2KDxOoBKprBKga
DXF0SARTyUYYf8pbKd4H22jEZ60dxbL9OofoXiRX4wB+Dy0aKczebQtfQEWveRDv
PnHAPRhhYurBctN5tN2w3GzQYTV5260h+KzH3HIU1ms6DSJrlZWtaZKl859jrb14
DCKuZVjonwjgkW9Z21df0GUWtKudjF2pCxkprqouXgEQ1CqV1eBOI2rftKKolhsc
GtDK72HM/UAtNBbR5WfoeEDntsgbxHZAHioB+Hno3i15O5Z7nSkhNspqUtY5jXjp
t0NJEtAk3iqyADzn35xReRDw8C2EtBTLE53dggg+pyMk5bMoaeFXZeCbQl3R/sNL
Q2nQ9/TyEEN+hy5YDV8WayNlD5/Lsk6K8tJtojaLQ8iezAIx3XnJ31Ggp7B/hve7
aj4lySm+0hkAFqCuBJODTmmTjc5RdOGJMnuZA/0043XfudvJzih9EpbYnhZxfrRN
xSYrg4LAx9z2uxIxOjz9qwmf63jzUBhAV1AaNU22+MIHiSSmKRtYITXN0NyZz2Jp
W6oLJ7VZLuMH4+WZZrnEVTRsDkAdthSnJp1eFEBEUSo9HaKV0Cavy6ik0RdP22mQ
FHP08U3Xpf5fxXydGVNTtJ7Z+HiF2/QmEaB+NBB0d4muyRW9BCT6/4fZ+VHZOhNM
O7KW5OdaYaJllPn7lGjKhXZ35BmpqIB0lplHS/ej5TT3JLZ/JPzfClgd7TQE2fCI
PZZtBU1Ixj33tTRpL+YGvx0MSX+qg36PZxOr/GfGs/lB1OOsxRGlmeNxSGuu21Qk
KsHETF8o3f18pQhft8N98AvIwazxzXk4S3folZq3WNJ2z3XYsSztPnv7Yeo8kjJF
sNGZOz4n5AmWwGluGlizfF0AU2pM4kU5g6KPU/2J4RVO6E8pDuElIaaI/O4hERlp
bej3q5ltbpjELKcIQlx2hctRB6cn/JGRWoEAkfLSF5mp0WTbN4Tsm+HxXoodyvRG
x5hXk3b2Ed4a3ZcjAEp0CNSTDTRL/7tTxr+I6qB+7snQL1d+pjCpdnEtAMAV95KJ
JMRzJ53rqsbsqyCRBdvA7gGJgVxRuOk4UJ7wKD2OeB38y9Xjb8h39rMgi0S2GC8X
YjD0XfBSfCQIF5ziDk0S6zaDMEnbJ05QgPhBUycK9EcQ/1X1BM9U+5ISqRoXCOIo
KssRVyKyFuC5RM0iuk7jzdkOpygHJMQdftyZX81srxY=
`protect END_PROTECTED
