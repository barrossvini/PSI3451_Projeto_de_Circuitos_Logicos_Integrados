`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8LWVlb84mObUrKoS/eud6yQ23TwaWvbkzCdo9RXjytrgW5oc9Fry+E/Jb1Gxkfl
1yzs8UhddCp6UrQ9ZsfTEHPpn3N+/dohk8u5kupxRUrYYqufevQzl2s/2RDbo/5P
DEVudYLd6xU/KcL5+ezAZAHqXiixui7CqGV02EUq1a80aNgnzte/xIaZ/HjO5lVU
Usf7wCHOGKNk76QmFVjZ3pWFrw5HTeiSvtuzFmeYZKkY48GX3AQC9NgwcSzyi9ax
In+dxvApURnst08l7vYFPsfTcEe25X3Kf/qELgCDGKAW+3UcMmieAIQ2qTjgQojL
bXToYfjOpDhC+hZZo9RM+fNkIFkFpwiPqXan3dGQGVJd42QpLaMJyGc5K66IBnpe
8L9Jfdb3nPpryXR191gKTedpcaGms4OOp3KTjpckOzM=
`protect END_PROTECTED
