`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8faW0M6Zi8vM4l9VkqHxgDjZjtxmVhjRps3l3DS+ZNkfTOnQopCDEEjvWtsLOdkF
YxaU3garGOXM3WVHenhxRzKaULtH0WRXxUkILosTsfc7dWPIxPgSyd4SDwkVsBSj
y8qSBAVpp/ksIeZEuABvIjeiK+DKyR/VpcYAd24kjv5GgUKgkSpstincY9C7JXmu
PM0KJHm8tV0kCFvzYn9CoQ4yOOIbmu0VDW0+VkSpKiRciySeIBh1uXhb/qj33CeH
FwLgCaJfbj2U56lhBXucc5qsW4rCuhJ3dKfw4Ig95BtfDseal/Zd1tub00wV6gbB
UjzBD/48Pjl3xFZK28V0hohqCgP7ZoDQuyjF/gGdhMlpeCL3lPHgpgqgf9E5tjU2
0+awb2Nw+e8HLVFrrKYRR0hqMnTkrROhvWWpQUXoRZxR9Krot49aSvSQ8rEnJMiG
WEK3YZ8QFKCcqXf6EnS9NzoZj/G+ewldr/TEihsZHszrKRSjHXdX4y0VpAzlyY3/
uHzaiyreXHifgHXU31lYffYtSOAo2UyCb7KVPqnjKO06JP7UTZ4Y2ulZMPh+TnSa
cIji9yxdKOVn+tNX109uW7y9vdMazumBjrBrtMbYFgdjxFvUFPhgm0pDrPRpq21q
S+Qv3ooCFeYSoqcRuE40YxVCSZXN9nS5TMbfCqIeuI+8yg9BNczR4tcJnbufPSbX
e3+2b/N5hKyK6iElpSZtwCADrXCGkicTVEBe8j6GlfImReE2Tj36Ir06Ba/FpBi5
QVYD3qUMgtgd/VdskDIYidOFM878v7kMMzQstENEr65u02Owu53+hDIiZcyxlwbx
cCc0Pz9Kw1YuF8ff1D8wmCkk4PpiiaDG2/yHaP9E4cIpgUVzZG6xuGwSNGZdNRbO
hXRFyEQH34IomS0sIyRVz/nYNbHT21X7Fa81+4LsSNsmEnaTTxuitEhFn1tUMM9+
`protect END_PROTECTED
