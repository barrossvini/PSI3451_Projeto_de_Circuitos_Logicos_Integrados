`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OpId9V4vLWhyYa1PD03+O9Bo09f4boo7osYHymsjGy+bLinl16tlSS7394Ybc+mX
AWVtwBlQU+W8Dz/1XT9bQjV48Xu7Sdce/G8Tk4zqW2GOFuZn4qvSd6j36uo2Z0Ww
0NvMCPpgNUdvSvAqtFz0diQJVuXDqGSNFDPP/88YcPBxwIzhmL5GCmhAGNxorWUp
ytuIdtHS4TQbCZtdLOnsQfoagaMlviwOej1d30Unhrj6OYpvH1gSFl+W+4yxUnV2
1Rj+dCwilvaNURRGnZnaRDEswj5xWYvlh3qLj+kRt5kdVARhR9nVMctOB7358gQ6
eunyc3oSnjJ5XZrnVtMaO/Lxb6tuFQBIdmONNTtrgeRYcAg05BbV29ANsyjQpHNV
vyFIXwmb3MXBESDb+8PHGc3Y2ecqZCNKca80iQYERLqlknM8+n3rti90+kxjC3hq
GSGnaDc3b2txGfWfVoVpR/OCF1vo2E8OiIdKNhN7tWTr/b8dfshYMFBaXvC2aLqV
Jwc81nKV0P74XPA1cY7TlDCog+6nIxaPEIi9vKjLHdoKOOLxpEgUrEb+PYejgIPY
y6xyz0047lyU+4hDadyQEAifWOVmzE1vwUSKj56l9f32rWHKzbDSc8XIZt9r8Thd
gP8uLhWSLIh6KdCw1MjVhhAC2OVI9wSIz7D4WjpB2DgTjRrghsBZ3O/S4p/bYgL7
BmQV8sKseBmcL7RuffIu5clWb0DEAWg/Ez9arf9gas66lYLSxNbYSMssLBFxwFpP
0mRF5dpGzgg6PDLne1ebqqj9dM7cejtMy6QY2Rs9bihjhiVBr9RhntbZ4Gu1uHhj
e2SzsHJ60+Lg0plt2qEJE32BbKTZ7QYzjjoisU290We+vfcs5WSLFHM+sY8B3ZCv
ZV+JBsI8eUCdUZo3Wl9q1H9hOragmCl1oC7mdcYBfF7rCIEz5G0hZAczC4O2iLLx
n+lLjcB/LsNC3tmhWFMPE6WVsXO1GREkSf3w7swgIArMPiZ7XR3vGN4ypvwis3US
cwPjcRrIIZeOb9PgNlJnwnAo9hPHfDQwI1He7BFI1OkJMTK1FMM0acHJWXj9AX9a
JBkaoz/7v1pGmPdCGKZcsx7LfEClzBhwVva1EBfnnaJOrMKZjKyK0aop3FFKXmCk
t7H1J8i7MUwuUTKPniOSE0R2aW2CXbiEdC80Ndk4+G84gL+lDiWDJC9w2xe+JuC8
uu0NJWYPs0ckOy9BAGuNp5mZdxXpc93LtSHEcbXexfORl44aKqmMe0c6ZYldyTbC
UrVF29DdRxtxqCOQys6R97YFQMl0sCNtuKx/4q//SAoTGaA2Ueewfng0n+z+D8Y4
0aP+tZ0RDCqverUqM2Q3/HoDp7/f36Yg71TuZxKpeVCW9kHwKBCGYEotyrl8Wu63
9djniUJlnENdwO1cjn5Fsp8IdGhE0qMSzowz0R4/O624LGjG7J+TZ/knN3C7voBY
RQcl/H3KfPNZRVY/6kUok+8okJylq7YrjS4N3hriv8s7x6lI9PMZBDWMpYCX8q0f
sSHr1jrDJPdDchKka4V8ISFRowx+0JCKtnPnSLGrA6klL8PTm3LVv5hpur3tNa/G
Oqzt9Bjexmo8itivbXRrIvQ9z522h3sk9A+Skq6DX0/N19i6U7zY0BroiZi01cJ4
qPIs5xTvyt9OdoFOiz0iIQEz6qP/qn/IIxml8xtWnmir6F2qzSVUTsGvsj/61mwO
heR0/kcu+Y8zHU023HrksP/IiDxurq0Y+zg/ppOBxDYqGFTEWEsNO56KsSrTzLGY
7EYQ8td2BjSoipWTOEshRQXKAqmrDKKzbpfEE8TP8VGoogsdgVD2a+Yol70BxXBQ
6xU93lLe1XiTiio4H2yAo7wKRA1hcSS63tK7TsZVST3D2UiV29PCQTJyO4iKfDUj
v6Zm5pKMR5i4x4CUOfAhsBi8ls2DSk+r5wBxK9Ak8EQ=
`protect END_PROTECTED
