`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8E44bKbIjoMEHLXRhY0uk8hi/NBXwkaRvv4ucBuE9iVarfVD3tb6ExDKtw3kHunI
PBq8JujkJOwb1v9zpOUmNvjxsXnzvk0As75lrASn098nhx5DgF5v4YaHjCCXK/ji
GQPq8Rzbzp+qp8L0dvSaUfHbOpsl/IMcIVJFUhE+zyyS2lVW9SfAbBSF5cvbjwo4
L7zyJqsWd6I9Xwu4TyDlGT1Y6ETCLcBbpomiXgY6xHJH60hlNwhQgNCcRXhsODb7
XSVFOSrB/SkkPFDy72r5rEYeU6SU6IqKqgXlvpyHFxX710D2QqX/dH/LxbTaSR77
VNfQxYlINiHXxy5f3gQdLeClbSqkXcsFJhagXs7N1e6SYpjGTU1YgUbYnm7vUIpc
kPU5mAvqlQE9DGb+4Y+fuaqruj9Ie1Qxe7JRBU5EBcKarsin9v+RbJbm28o79Ydv
xnzSvTNyENM+lDgHfDyy7uoolWQa0uQGuQVCpqAlvSvk6SikPMrlnADFBoHFTeFp
qpwaV1Q77P6UkyEa5QyeLWh7gL3K0B15KyqpX883lY70LsP3sMYYgxQtgQMpFtDu
w9ibiJNm/FAx4s8YonNwjTq6MyJQWVixjKI9N96bfGB3OXajxRupG/7YspZWv4qr
fvPassDlghuyNOibjIvMckzCNUC/wckqyHJUvvpjLPG1ExybyWBjckl51d+efwEv
shLebrG4VySKqPTB2XKN3KMMjmUhcFhNvS9yt8Q9V793YyFJuOmIpRZxWQ3UwNxR
ShAxAa2bMxU4Fmgp5JA99RpOuh6Kp8HyYL6i0avaNTtR47yqnq029O/cl/USVtcw
ocfLM+EnS1/g8eoiHlJptj75wwo3yayM4qNeAtrF7kp1BL2oFRsOEKulYkpHjF/x
J0RF+ORHWg5nQdNktWfGNFgJPwtkO/Lp0bPnvQDUqWUd/pLnAPll+tWtuW5CXJe9
eNcTLj1mUjZrFTI+uD+SAjzJygguEfq/sq7DPBpeiOOCJxNrKInJyWa1yc5mR9R8
9Ql8QXaFWOoRV7PuyCPIyzhZuxPhRYU5Tep4/uYSpuHR8WMNxUQBYvqOZVtRJ2GQ
EoSmpyRhvCMBgzCFbU9AH0NtHEq2aQQLqgpyo7K4FXCN86ZExiH18xDFXCc0wPKH
KHNOjhnL2RAVTSyS9JBi5OFiSBhQrb02gsabG1pclRszRU6rA1w5PgLnur3EsENr
7wy+z9o8UmHGxGRpFmvcHWU3tg2SdviJ0X1B6XiIS1SNPliyD7K8BX30UhsK7hGu
x96cZ5UKvHsZlMDp12S4YGrXhpqKFHC2XKy7V9JNn/OMRzLZaqSjUNHWTyyOEVsu
HV4otrrjrVdPfFJznxvl8KZ0ACTZe+Hf4P605laYB7esQM/wzOoy03WH3vfzidw6
4V6a2uk9ZoFP/Jo3OYWvFXE13YtpgAO5XMDc+LwQgbkjau/JymD5Hn7vD3C0x+P/
Yd9mv2+/ZUnHzOv86nln6iBfB3jV2HlINE+MubBmBbxRUgzFS1QlIJ3KkSDu/cKq
2m92o9hbRP0C9g176iwSl5eVe36CWzQeLGWuL1Imv1SPN1Vn+Ml8LeohEY6DY88y
v5IPYv6SKDAWBjgpR/Wgu1k2Cw9NlbEm1Ri1dGnPQsObZ4tzrn46sYq67BkQmv7L
N8dxif3ZQbZrCZ6QWlxL940WJzxnLpernLmvFIoIjSsr6pOyTIfzHYWSKaiq6/Qk
++iGaJQjcCm1HE1JIP473iFTxLCLYrKq/zK3aFWegXwvlYtJwCBTNEYhKdTuJHoK
zSSeiOOSMpJDkrzkfc/wcA==
`protect END_PROTECTED
