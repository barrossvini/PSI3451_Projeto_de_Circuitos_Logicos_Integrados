`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
15i8pNmp9iqfqFMp2U4fDaldKkGg2KjGTdHZN1vkHY4tSh6iFz8di90CEsXfhVo9
saQbXXjVGNTv2BmXXcAH0m/hk0mpjonaMBrqf1cr/W1vhJsiHDKvAB4kvxvVHer9
9f5biy5K9lPgDaNnprJH634A/8MAw2m9SlXqi23V3vuzQcaSmSkfBHoBsAkyRaa9
d9J1LJUNyER2Fe6hA5hxQX46VSCAmUvXP7mR2pxeuH0rvZhsj3aeJEYQcvLG53K2
xVWdmDZsG5fP4c3txKui9P4VSeKmp8DFMSjNPAekQhaE8sCSliG239CCZSoMXwSg
sWD3HoxN0aF57wr7EgPO99jF5FLvUzXVJWEy8gtbYLqiYEhPzcEnqB60z0thNQbm
R0x5Yg2SOtpK5ObGbZaAV1yzSA5g5AU7FY3zkEk2O52jZqpAcbAdB7uCUumQQOda
glfQfwQc4+jOX0WcaOXWjhdysOTzGAzOxGZal8AisaNoQw1aw6OVvRLHINyrOKxg
7PiiGusAuDUogFFZ0b3eg7Shm/YdqeKKZ4LAlGxNAHqojd31lqjwMXvaB84kGC10
b2qB66PQILF/vR2oSUsqUU77LtWvBjBWvmniftUfVB51fJJ9BPG1uGFnUj6EoyAM
rNZykQpliXdqvu39nk4uxgiUyx2mMr1I+etQJAuOD/BB12Ry3SSFJPmqvmmPVLaX
Tu6c9SuAm1v/spcirmMGVBO+Pt3locuqRNdwsPb8asMkiFVkaou9B7ErTPBdBO7z
xLkfbbZRoQvV06CnS8UEO9z+MKq7UUa9LGU5MFSmYcIwQ8DLrVm0Af2RP8tbGzei
UMoFW6koq/+6DozZop3dotT7QCF9ecYwT+z85sl51AL7GOWqAUyPxa3doxwby/0A
t5qgAqiz8PiNFTK4/cpfXmDcWPJy6ltmSntgzkHk3mLpixYcII3pVMMc/mab4KpO
aetfvbFR8eCTqaxmhO0gVgU90gj3d6aE1hAI5f57ZIP/WDfiwJEGVyNM+c7Bgc3E
jz0IMcy3O92r4LbyvGOCnnP4I1hRyTMmGnN0YpWoFVKAtFmAqojO/wfQ5iwffCLy
Ezk3sjRZ4OybJ5VtgCX2MUhku+FNF+DLFMI0ZXEBEdQxqUc8YtIZb1pwF3hU16Jl
0WtpiMGASQ1lUmeaHZkXMS1EOYrC+SXIz/9pBlFPZ2lGUkEgjRPIAs2zdSiD4UxZ
jfop2jLT6UPNyJz0TWcmNdgEoxI891k0DkVC4GtdJ43iRpFA7iI0KJzNY6ubRgGP
VU3qVHx/Le2wcKy3Mg++37XKHGSgOjheVUWzzYtyybHN3SivMhV+rLcaFPUGXZ1l
Wdkz8hXWZs1wRFzCwF2zUlcxHvnz/7gRrbdnHh196GaM6mxMwUpuqUMJVmpAI/Ot
uOXKR62vWS/hivCAxKJK+P9BoliMD+hf6f6IpeF/clhaD1YTpCxDsdMC+AzECEj7
rtaH/Nexg7Seelctpk23Zpe+EooV9wANbIa8SQYIuLEZkvHid5aGbC/aUVmOdmKr
yGXA4rnJfYok3iMXeHmN910yKQub0512mkJMmGvhXJUSFx8+EKINZBWfMqVbDqRp
Got3bCdY5IXUobuHiEIQqFZofAEbGuxuZ8ID3ee48NoYFFaxz6v2cNjCuFRUvuiM
kN9O3fH/p7sydTGpn56rx+LQulWxevQvKPypMQnBzPoUyGYlbfoNvGAa2Zh/NHya
hUTPIYDfauH6e1/qgF+6uQwBNVOnWEvZ1AUliEvYftSWxotoiD/jvDm7HwqrBPVM
z2F3vALT60AHPXiZsxfQCec37FiFcGLRqs2tWWhDnGHts936rrLwuNYigTmZF9Fe
tAHFJvatw2WpLnRM8xZzGNoMZCUY+eqld2+QyHWSGA8Pe/frUE80zURaEMj2i70W
lRjnfCDUD4iOC+0iqcnjXr4VhmjK/h1KMaerSi+6tCKyj2fXzTkzIcdnMdyJTJyi
KTEPbQXksopT6ERfJ5rifVuJ9Z/5vOgHEsEyHkX5Oep4XM9+wOW7KoR5LIzZsK9u
d4pj+MkeWBo8FRy1RkTgEDl7ovXTcyWlEmR/Ze3g1vTNn9CewNHSuPTgbsbr0PnU
NFepoIFVTXn2xfW6gyHSTNb9gsK7XxYUTHAlhSN0CMRxgQ8QHGorOH8N8kqcGTS8
FbWYj2RSLuxoIy7aP1nTzgFHhi4mKuz2YaQYFzTJSzhRvOr+CBcwuQzg7ibWBKAi
IrkwIcLcMSy+dSeHBQJjA0f1iOz826/V/fqDDUekzDMVtxUdeSDQHxUd9Ys4gJq9
0e7QhP4aka9u4WVoxmICcg6tXqHQa2U8yJnlCXRd69cx0wHvNcnoNqR0zKCKQRp9
/NbsIOLYI9JvkTCHysLB9evffmCMYmYarviOdmfRrrmFuODJzF+Q09hvn4s1OyZh
qZYg/WDTfrkBDMNska+MGGafkf8ztq4I0BAXjp6V5XcXtCjT/Wj7dtwc034dXyAg
xJP8pnZRRhgSbUoZKCVG7ghvZ66KLtLfHJJdIcMgpHqAu0yjaWROVclFSu1OT3z4
I3l0l5HGkbTfS6fbT7Nr7SDgeepE95sXQ2o0p4IrnQ7l3sno3h/bmEEQQUHELDzv
RFs4GKtnDU/jyv7J3hvOXtfMi9OEGfMp3l21tBHHDGpeDZA6rExoqrN2ieRxrKis
R7mYaT/T1CiLxWmUhyiEWlIKOjdrIDDAV77MQl6WmTPWB7GFz1vNA/8geB/TNBOa
AS2a3PVs28eKe2i/OtDeyyYtNGwcvwncxk5DS24CR6zOa/X8qob5ohExY8JB1R4f
SaeyHySsVbsn1Z63rJ5SfWnMaXDBJaN8eKEl6zw2P+auMCnjRIMvTBbNBQzUh7gc
XBY/Pi9p+yNxfbxEDqlvs0EnuXl9HdkKjWkMkoeeZHJTMdPYHfI0u2fpXtXpFjAC
R4jLiMMUJY9mQlw4t2HKiZfCDmdWedyazZ8kQJG6xDIwNthVIskxSbl2Gbo/OlFa
T1tPBK3ynv1gEKnsGkvB/9/8xml1ANy7vqzxC4EpADcVwhdTq/End/5WTYh0aM5C
scOnuAeNQqBlI4/+JD/qe2TuT7V9FLy2/6rZbyKBeBnCEgKqCjrr22pChn5/VIw4
F4gUXWA4ZUVDvh/xMhfpivpgJ5mDMtuLl1L6SOKhKhuR7FXealDV3kfV65tQJy40
SQUEPbWWtFO8/3fXKXY2GD2J0rxBfdwtxqaNccvr7EnSqHrHl2j2kgTYUDaVNdp1
e9JlG64TPZuMLL7VF8JvOmwmiqAFLT/YA68EHGY5pmyT9ZMQAobyi/xf5PeixnwW
hwDlRaImkaTG11omoVLCX4DOEmwnKevH1VRnX7Ilu3n+gJ3zFnj+7ys5WZ8ThleS
zTsU70Om947+Ov7LjnAwMj0/c6FYE3dg4F0OEDHzWgDXR9kNz6GwFZCh0IP8YAXV
Xb2O1tz64754Lrsfq93SMRIHfh7HMa/hAqILAajpSQazS0R9TJDZxqd5g5fFHzgj
lBSkzyyMBs1O6xqgVmGMW8ZfVpLjZvQImYlE19yXKLz/PpyMCZTY3g4tKUCYUxRn
Bz9/RJIjvvzwziO8y9xAOxVg3zlM0W5Y2jaqaTWfrz0HQr/ROrPZLCgRZiQ6vIE+
b/6USAiOhYEIekVx5zk7EH6NxPUbiXWS+SIYgm3jXUiyQZLor7110/h2y9ys14GJ
oN5MKajfemL5pzq0IldFtQgtCTzx20Xekmo7kvnXaZotccjQbe9zm5sBy77AgIY3
H4nAXX42YkOfw4N9bzHLSjqZw4IUK42oeYQthECrVB3JTmpeL4MFpNv8oc5xn78d
v/wgNFpOJpjGwvGXr9BcV5qZTW6TGXrv64gE0vqUqRcBuiVWB5oRUrg5wBbZYXcU
5I9I+h7+Ps1hKS0RW8UClYUSwNbwNwGKosRPu1b/U1mRCKsBR1w/HUROM72LG72F
gAd6dG0NvDHm4+No753cjS9ttLQO478nWJ/eqORXPweAUwgsdv61M/F7WXxwo/oF
7sE9ZGM9MG4VkEvq3BGr4aWgo8aUXqZXdreR3wUG7WrigLW6C/CK2P5wGezZELmm
93SfXeZTXRXBDst2+Pj640pV/olfuuAuOP7FxH0M9075hhxB621+4gZWAixoUN2D
S4N7QYMKCF+7syaOdqaaTKnnlc/pJp5phyfb6viUI+yaiEe+3/ZUmTPzYAgqaI7v
nIg6in1lgJkJmlJboJZpOYBUi12+nKQ1lsgxbuzVKe2HkUveFy23EsBemHSqDL70
9EeehG/AzGJT5XVjXtcQ4oiTolhIvLm4nAsWQIdLx0JiB4wy7aV5E+d+GV+n8+XZ
9CPq5Uun9dYSMvCcbx9/8oHWRCSc7IaxCPJbk2pf8vXwK7w39Q+TaAz5Z80oWaSy
Om2o+VrFDLawAPS/qUzYb/mGxpDEeYJrZeTht0Gz5iy0xquYQ1GnH/ESKH8HCVAK
UaKtaeuCRRuaSNYI7SI5N0SfYh6E3sD5caxfAwlRDXC8dN+7UPl7KqGCsA698RcD
PP7zKRZ+31IZdzGc0MVkQwYaq65fdbvv7O4wZcU0HoJIyCoiTqp8M5NLLlda3Nql
cntwt/N9r5mwxpjeAtKM623HH3n82srtmaFpxHfcTXiqj0gzkADqeLSliKVrqHNO
Sp4dxfWrfREEZIvPsdQij6yOMss4EhEAMn67ElZ9gfVwb7Hd5D4u9Kfbp9oWPCeL
wkys8i+cf7scNs5Ui2ic19bVVotGiGIAcHNxFQY9BrDj9NMzVfSmHEw1slX4P1nY
kIeyJjEW9l2JyE5FQ8Fipr4nCE9N08eskN5qOH+OpArhwD7I+xdK5nrdVuA2ro16
Vt7vIpI57PdOqEWz7kyL3ognRexHk71Ed1L8zkFPjE/8KggOSOIsXqsbaGV0qkev
3KuwGf2qeJEq7nBa0yEj/N4/TpIAn1DzJiGZf/VwhOaY+IAsSb8fdNT+4OyrFrs5
+5Lx7LWqYSUgKT1tlXNpZh6uoW/08ESjeSndGF3GOPzMb2Fl4bTOhnG4tVv2DaAB
6q+UvrqWrwAOqDmctYwnqpk8/xYIsb/K2jTPTuSTlP5zr36YbaPj9mrJnyX/HdtF
JDOpRqD6eXmiEmZxqsdxfpg4W2dPK5zZbLlePshEc+HY4gPkII8iEqyLKLZb+QkH
y9Sz8yojN9ttmHifZNN/iR+wMwRqe5WqOOU76xnWXjVkLlqNJvaeEijsBbCIlpLu
vOvvmmROrwc1lCCkxwp3766/I8z0soVpkv6G4kyjDYgseO+7bohI7qJMjNZ3fcFz
IadEl9KW70FiCMmdD4CGucdSJcJ8J0KLPIjK34HwVmkQ5aj/NTvwWwgPaqs8X5Gw
1Sskd0AXKKybBgTLiG9gdAzbDH+3jTII0jnDFEnbEWSW0ywob7zjQAQYFYalp0U0
LUu7tA/2vFddXxe+HamnstcwxlUf4lo4OnlUrSr4ON+/DF5uSmFhZ3la+JWagZsX
zSgwyBeFFXj9dsuU3uVk1XvAtkRVON92xZWjnNLn9nShQ54N7Cmn1ykGI0jO7WW3
Gp4MvRTstW6NKvbKUflXoB3I4Exb1N7J0080ZZLYD1mvDqEotENOaTxHwJcfYRrh
edi6kgfFMeb7Ic1SaIQ3Ws30OyvZ1pCwl34LjcOZWGoBdcj8vCyv+jeaC8Tiedx2
fCPQnMqnpkyagpEoir4gyl4iPLgpbfr7YI2oIKqBd/na0WWFkbTdTCpEVmYG80o5
pB1OnwgABM0pamcDokZW3VXjIz1jkwaN6dfOwb8VoYX86XCHhkgub6Pukae+2tKq
NY/Jyn9Ty4CNp68++z3Qf7S0vEtyi2sFHBxSvi/488EemcNn7URu1HMehtR0hFKf
IkKX1b0/0keY3Y/K5XQPn7+bPGnJK2/i+Dj0XZxap4y+nVbGSn9ipdvZg9Qsh5wn
+3+bEaYB4etudLkqvQA4bEIbht0RSysEbrynqxJeHlcRqe3pIlNKzprTUhQ14Ox+
GcGMCtc6ZLdF3Hc6aiXCDjFLC7EXAcCzCOUzz63wthkAR+PMk8oqc+N28JTBi3OI
Z/BgatYJBU9pSMeQY2TXPIYAzgmjyCBXV/o7HQL1xLQ5Z9oYN09EhnR3TW6/gkIX
/ekmVGDvO70DThcJO8E7Gg==
`protect END_PROTECTED
