`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NlogoxG0NGGRlsJGKSJkz3nTOjs9rTHIOQkvtYhu49UfJhjLtcUOEy/JARYyX1n7
0hFSTuRV1OoeHhw2tp12nB/2kC0dE3n9qcegbORaDvjKh4S0LKEOAb7b5aP5m4G8
iwoDlWU3aJiDhOFFS79Zo0FT5kYIeCnYIlbL7rgd8ClXMH7voBD7cQo61F6q4IIn
EY58MVglBmq85bHi2HJ2u/txsrvK6onUn0X7iAFA4OSXNj7fOu3Uo9MzG/hxAkWK
pOtChO5UbWjeKdG7SO7qVdS2VyFud/mgVkur7x4RbmzJl4MfUKe8mfcBZLOhRRzj
rxf4U5scKc+uMimgEymnbdQ2xovbitnGrFNAlGveAWMIwFdFIBtdG/ozDxQwmlaN
IpRJgwXG/SCXOJ0ch2N+1ZC4QSQxv0rV2ji3GgXz+KKx0BVdo/+003a5wHnvEDG1
eOIRz1zeMNNQQz/Fa6x9i4i+8qujDjTVZ+XR2IqJj0GKKs7m7vB61Pm/UVJM7ci3
lZnpGAfgyhyJudqxGH/ReKnz0KxgRpX7NJeNpS+cdlho31uKC8IxDrPnmNONP49/
1AeYUpt194I3u2fUrSXN+88O9NlJXaAtN3Brf4tbpja0Y7T0SQHdM71bHj1WYUBh
c1B0Yxrxru9IJxIt/qbKmPxJmoZtH1za8qnn/qxf3tsuIPj8y0LT1eg7mUvh64Tg
w9tTpVh28XOWLITpDJAwkDufGmKl7/z1DZON7sXCwCjq/gmvGhLNEydin2/wSr5/
HO2UudZOAQSJzimupCp/Hc5Fb9U7uA5nSnERRsaq1fx7BIto4ysAGSd47fT+CHzh
0vCG9dMhZl3a33TULXAXsp9wpfhy4MISF5sFzHc0RF06AO5lv+uFZyPErVWfD098
0uEINUqcRfoXeb2Yk2NToDODUPw11B6qQgvXuj1XO27GDPqAKEc2UgUC+vvfMGoD
TFylzRcHjdgMgHGw/Y87yFQGu+GQsHqtdXz8SeSacFYYgR2HQcf/XfAHMCROoZWF
LMj2NpWh1FPX6EVhCtv7jPRTEcO2haDX5eMLG3bFuqFUx3fx3qB7KT0kvpuGUPov
tRSBukJX9fKX2nRDdSmS4RphOrcRVQkNVIX4jXaunrtua6aXwI3n1UrMR/pz0eB9
1StTZhcIfATZzUUolQOnzNR06c9A4nWi/kr/BqTNRaGWP0YQTI++dM3Z25KRa/Tm
W2jGTVTwlR5uRSLxeZamabqce/MymZdHzQaArkVBinUWn4+Cske7aXVmZeg78HYH
eTI7wVTXDSxJ5wkaLeuzuBRucfYRUSQTBtSnLXxl07qb3E0Sd0XfZ/efi12yIncw
R7aHpmdFLD3Mx2J0cExj8/KM7pcS+5N8C9433axyafh5aGYZndGZ0fUFVCD2nWw8
ccJUbkr0Do3TmRHTE2dxYi66e8+GYfl2CWeXLHGekfsJXg580v/z3lJjHSkcVpct
DRxfXxAtBo8g9YnjREQM/S44fCMEZe8gWHz3f6oNEdourCH1RecNuaoZu10tezjf
RclZGoEsfR6hMcjWhJFlWO6nWAP/9G0zKyPGj9VF/xyRV4oV2TeRWBD3AkiNJvDw
MvYB9GvhRjuGXKm5hacwy2rLMNKKrwHysqC0//bcaQLkj2R2H7SWkjSkbtlCHl4e
yxfsbkBzsHjJAW7zeaJgcufR0nYXezoAcEx/kNay4ENK16ehgEnssU1Xm3hDfqwG
v/HC2b8R3jBHt/78tSM1nkggKZa9lz+/Jdh+7BbMLNqS9c336TulhHn33TdpJD2F
3wQxY6l0AwX28JdqwVQGsYLgBynvAWYohHUB5QnKMO7Ea5/Fjt4A5xct1hVDGAzU
CdFMc4DudKcGBUEUXtBNkW3y11niwK/9u6ow4pAugPTdCnMUHmkgwHFUk3fcSBhP
ONhCDhQQ/yPuOX06FIekODlRXk+hfK6qFvT9gT+OsbvMhKlbuw0uksQm50y2NpH5
UAUuvYoUJrQbYBaG95TGMODw9AG79Xi9u60tj7BXcIXsyP4gp+W8A/y4zAvr0gxL
Vn/2REDFWK0ZYDVZKsQU5+z9xozwcFbnbU8GMGMYqhYkVmJWGOgfcRDE4SmgTp/0
ZSarWlby25a4G8BSZIN41d15gbCC6caRoIwpSIkRsxs+y/Pk7MVJV7zA2idIWOpr
+x1ejxtSUf9DfqrCSnzKRbNarZaahF15rCaRn75yl8RzJb3k+Eo+IIpoW/jJwY9s
htaJYSQSmpOyuVIGWfkOWoizBvEIZHzMrNKsOQZjj1rpeJ1SPAElKuJailDDwD9H
Q+UN9FCLxuZvttqlvAEi1CK5W0Xt2Uq56Hz2vigD03SoDFsHzJ0rfa0B1cOXNHuB
ciMkGEoUVnKNChGhaXTpRMw2kgCgwzHePXuQnPoHBYlzZObERvcs5e+1fKpOHGdu
7pU80FrKE8DH4XZ69rD1M+CwJgi6O9LFw8T+B/RSYIiM86SUZeoiQfFhZ1Y1FCVu
US92uEug7UzzOnrucQAJzgdHs8Q0jMbVzRFdfZP4RKwptjK1aSxa/8yxpW6Z/nth
Prh2+sgwvU1ykFax7khNeRQc3SQTrcYW7PqKRu0ceFPYM7Ivbl9JSJI5EklbDiMR
dHA62b9aXSX2Puis0yUMBSSpPyrAzV/FqmKjRDa+fzij7Ag1/bN0h5mKuSoJPjuh
pMuNjGqBtWqlDwwInDj6eUjdw9JiNnB8ulErPV6b4Fr8MCgMcsTmOUoknJ9wW2Qi
eVrmjJdy11sfIDGj12vZmN8QLQ9d55CY7jiCdghbIutUdIS/97kl1PdV3yizGySb
WjEFCZSE26GOV3B6tse+l+pz+ycg8YL/I2WexJkCh8jS+neiUUfQUXI26fpsEyV2
v77pheLa/iJxPr5h1vuQPAJvv3sG6wFsOzk6JcFLLExzSP5hkITldEK3PvGH3vAa
7PlVQzM35LhYuTMtZcE3d/lRW+vSxSy/DVKOreOlEMtpLR7HB8h00NIprlNzKqvM
Cblre1YfSEGY3iUO0MgN7JucAkosr+nASbRCNJCtBDa5xaO1U7SBTrYy8p3iXPUp
/Wv1PvV584Fij+PhfsCsyZ42gsmjwgjEVjiohCIPxa+w+yroMAV3g/ksULUfFpR6
LOjL4jRZbk58xLhpAiyvD3sgYn7y7tEYnX6G3IhrQuDJffND+OMv2OgvC+KZzeb0
iJ8ec2zXMnz6M3ewB4A7u6TOtGnbJ9AckD4W8biH9gks01gmC9OKjMmbyP6PsWKj
BndyHArl5r3kjJOhlMXArYMGH/7wZI0fiOMkZGC0ErgD3B2FcsB0yMsVlJ1DzMhw
CpD+/RC6XLIALmR9tljoLCLHsGSe5px0fxa5zbBShp5EsfAfByo/AvkmUPxLpcYS
FXVn12V1zHjM56pOg974VlGjPO8PAKL5Y3Ce/RPYnYUU1SbBdHTzoLISqPGk3O4K
2Jw43P/6YIU8r9UuXTPVDOyl2S6qjC0ZNgOXi+DUqymFrJHjrnoTatAZ2Rq9Zz9e
JTtelnzdp/rsgfirutdnqdi8pIaIqtJGma0lrUdcKurPjwNsPjJRKUr6CWY3+fAH
6+maNY1srsSudTApfL3w2CrTzRK7rWzj4VptvIbSk5KnRfDRHeTPyBD+iBZiT3/w
9E3qF1lsla2yJRKjcnVNa1xkMTiuy5WmTP09buN7TnMvF6/5p7S5q+F4qMNdeGl8
5jTFfM8ieaYrL/B3YqtFm/i6FH+bxNrS6m/RP5zj7A5lcXJ45XwUE7Vzkk/2zIwZ
bhFzYrf+YOBeKpaSfkS8BVBjQi0+ylMf3BTZKVKCGPC5AfUU5pXcyB0Kq+K2jNJ/
7gD8Un3mL8/9yk1bapuejgHb+6zzAsDe+FpOmQjuszZJy9FhWR5tJOpXmhsYeyrb
yImzBG4vHELkp5y7h8VnpZ5Y1yXocLAmXpRPG9RuwSNOdT0d56lFdI2E7FP2oA7N
n7emEu04X3IaxtQfiAndF0ohq0K0Ff9xjnbzZxHPFMZXZQ+WBjihj31UuRd0wcua
OQqwYgm9iO/KPWob3DXm+5W73ZUZKH+7SJVeZ9csg9q+K/s+3SO8flziRyxOevi+
OyX76fcYsbgKbbnCzVWgMrRyfau3tl+MvSOaoKRa9V/yhrsvZs0jGca3XQuycFzW
rtPkMG44p8mSYpHPaI+D269cxUzlcy2TWk1MgMRhOw2Qai3YyO7Klxej8lscWZFn
w/NnJDztpNuKn1sXncvb4AkW1MMckMNCinxpb3xFTQQbpmk8H6cMS3SO352TsomF
uG1j8WVquoUM94KIqY9KOYWwqZtKLoh+ERPViue7E9wtNU4ZMHaCgGjOrdQnBRIe
DFSkAmTBod0O7t7FQUGenmqMzbDWjMgRt0wchu7SisDFIl0eR8fIGf1muAr9h8bU
uRfsHrc+VfE6pMuMZP3e7Becicnka56G2jvyFcOeLzZeEGYdobj1gdm5D0kyoi6X
UW+1yCJtN83TofRnE2MHhL+iFR4DIBYvSbxbWO0lGsH49WwH/Fi0iFGFgh4OsW1f
wFw1UO450dGiFrE7bbRzjFwcde8C1Ay1BqV28Q5aoG//bSZEAVhaH8Qedm3nismX
UBdotzQ63PjD8WaGucXmcQft9j50Kd4xXwBfPm2VH8VVOlplK4D8/l1GrmTHBxJV
lblTIQoiFhDatEaMxfC7I6sT3kBcj6Qy2KOzncOwOEU6eQJnEuhjvF8DDg2NsAUO
79Sdev8moVbBoSbC7EBY2BxPJ7xqb+fBOnR82bAO5s6O94qVtdBHMu6kALeNM4OP
rkDD7i4BlWBFx95OVTP5jGjFUDedw9WsIVcyR1swjdD2IftZy87qUu9Ia24wRdlS
KLyQ9XX+udZanMJWo1AmjBp5EXttkaiJu+Fv/SaYMiDJuHbek+s5kI8pgMKHm+Xf
8uhPT7sFaxwo9a7VdvyBaZBIX05DUmjc4zmvcggVO2ulQ+Nf+4BuiA2NndPhQzlY
JPm+L2UVxO9ksunFQZqMkCd5kgW/WTaf0ljz9nfsqc/Yb0YgUReLmNVUovbeEcUC
rTKYX8n3KiE1VT5Q9eHzYYUMUoTGmKCHLqqnBPVcphhpAXubZHM/dpZlzC898pab
tlkY9f27FHqyZu8Ma7TeCkVtlcP/hjW4SoM6PBYVR2Y56kxAArNGNwQi83e28a8c
DxXVcrZZTgNf9dFV47fVcB5vNkcRvPduWCQuSbxghJL+DK+7IO3ETJM2pNlIPe7A
RatTj/MXC2QQDR5K2hUxyGMW5n6ZOd0ArhMoJNOTAFXwMaKXYB88OD0jypz92jRx
4Pg5LgYhhMZR0Rv78QyW4/QAmjavK2XcMwU9koImm8ogJK0E1pqWvpFWeutOM/Uu
ED+U7urwkka6OjooMVuhdLRSaq1hoWTAI5b00LqopfWDJlG6h9nDNeF/zatlmjeO
ICPTWz5ACb7JM8qZU+pvQ1malFrVRFXk5dTLm6xJv+m4oQQaBLqc3MdIFBLT5NPu
1XbNgo16niAEjDZrCYiK33U9O4nxWn7oMj4gKqFYCy7N89Bj/YlHlY8a4QvSD6XY
ijj+v4Gw4hSqblldWV5KQOx/zmEqyfX3s/b5VzC7dKWQqTNfIQzK+dVGY9Lh1z93
Gk7c+a6Qcf6TPpQJM5Y6WgVpv/W7AJXp1Z5usvVnAsQlRGMkBofmBNYT6iSuNilx
n9wsdj+5fh6RrfKrSPL6ic4UpqNGZcM5rXDKSY9DsEiYwrGsGGP3BVPFh9+rCccm
Yi1Ixqd3zN+Kl2UrjrMT8dVo9z+KzzexcTXvMMeh/9SmapuXs3hcUurqrWUvoTGp
hvbPYJD+HiRumK5vzXCGs1Bx7fIt8Kkm/AWmEhAwlF8=
`protect END_PROTECTED
