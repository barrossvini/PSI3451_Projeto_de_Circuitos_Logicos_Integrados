`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
acpu7C1fYf8M7j5efd7JbBGCQMMpCO248SQAS9WOcldUZJYs04639tCol7qEnlUh
rz6v7OPpKoflQu8oWstNwprbdBTciDqRqC/WVjRByXD3OCwpfcaAvFl5WKizPgTp
PfIv9D2xVlHS3kRDxWlqxTx5yiRiZKnmeYTF1RpjZaCun+ZxkAxVC5dutFUxmQMQ
prg1+pn/4pP+8ELhGlFB7pC/18F11Zl4B3CmzWkk7V265pRo8o6Ae43F7RGGgXIZ
VA3tkNGPrptYxtbjPiCS09VAHrXN+izH3n/xwHIWp7MLhUq9FB2nTZJvyPmQsWUq
qDkgV4ps2TYl/VBVJsk594AsHvgmM2RiTwjioU0doexebakSxlu+z1sprR8J4MgI
Cf1gMANd7nIG2TjgTMJNzbP6RM9RdZnzzo0QO+x7Q8a16dU4lKErK1PJOt0aY4yW
y+BmaPwySkEDx+BDS4q4HqW0DnOE/yKhibDwITS5KifnabOFQproM/7N4GL2rfSF
xqpi83OLgH1vq7yJt/lLv6Nbdmkgp2gn/4ImGT32gV5awoQS7xgkhppP63s32Fab
l9s9Jb3IkCsD+FgyadAE6wURVy+ZoPm11DPnEztxnvZoiMA0CCk3ddX9ERbbBoqG
SNTiR25XCoYqsIcWRTDWMD0C3tNG58WUDChK3x0k3u71g2yVCkfGO01gItfWLbD/
TkNFHjrpxPKTf/R0dIqCe6rSXXCjgfZnZIvZlbZh8AJ/qdI13y8jrPuoWHM9NAsS
0cjtNyS3EA29umnuhMu73R/zpjhv4ZBD3ighe3wGRJhlLznBN1MNHWm6WPgKGxqG
ANfuAmg9BDOrTibEbrZj5U1WSoAN6LXBzIFBz3z+X0N5PhRBiIU29w4NhVKovF5c
/4GYv46a/pP81KBShZ5FlcHBHLKkphfiA8l8JBzQDoskDtOIOSNyRrFdOR6RqbYc
wMq3EywSBvS/rL6ws5Fck/2x4EqTqixytEkdbZqvOL38Xw3ooszSZTqyoirm7SIV
1Y1vyZqnU46wBB2c9OfJ2ho13UUVT5QURciqWLRUHtCdbw07470xPrjPQdIr5QML
Q7lpnsv5F9/sTWQqcbvyagKAArXHAqM4jPbO1uee1wVNhVoPzApA5QkFYW/f2nM+
s4tyhuLHVlsncn35f2DGg+I0C0tQT2O98ds5xBQ/a51V5Wwxcw9amXZHc0T/Xej1
y9uEzALxID/W/SvYDT0M7NJdnRAG17w/xq546z+5BOZf8gHcYgIVBBt/IbV5WpGu
S15kUxxy9ny2hyQYQCCPhbrdaouP2serh+b4fuwkrtGJ+oDIt6JZSaJguGz2J7Lk
4T8P62ypRHhUhZdbEWxe+ptfZ5M6GeSz1Yd8/NDLnl++F3u8exO+z2OTlk6ZQh/i
eqIsg9ZSL15nSh1F/6qIOK94juIJxQNWOHlEeA7Kd9ZSdsP/rmj46eESpNabFJfK
RaEbIf7llRWBoUUULIPMsjB3R4+cvACb8ncFliA6KQSragxr4dYtpi2x2f4CLGlK
z/vz158Rce/GvIntZ3Iq3PFAztsb810bep/3+oB3fNzUwGyde1sq8FH1SAiNzU85
bL6A2vSOcDbJ++1Mr7P7q1qHpAT+lfhnG+mOS5yJRiIy7bQTis/rX7+qahkl3An/
10U4/LRA9BTKkfXEuWgAwoYTp479XYAEAz8i8xkoe6+QNN8E8XnePiToHDzXksSx
f+Ghsck6BNXLjwnt2YVbGh5Ihax+zjFsWVBFz6FSY7DOKWO55HzuzEYzOBDUv5Gw
sgnmwp6C7r2QSpRaUCx0OpAfSRBIR3nP3tfqLARQxAyajmLOac+N+/7ZsOScNXJ6
s4ltahpuRIkboHVsP5pRsdbVuB2uEnewNexjcXLLax9wTDhZVuUFD909PnxtkLkz
aGCIhACV3PH6bZVXcZZtDQdCmuEzPIczSDP6ea2eygvMPnKRsgKBFWmIo4FYyFwh
DKBgYwf17YK/NWDooplcplycy39DkpP98wWOhISFvOsN9oNvvwaKE01WstlbNjE1
AOMiXfYhVocoT8+iFQt2n+ywM0DhNyE/WBmpmCXt0MyaZPdqHKf0Yw2ePL+DgcgM
iRGdHAJD7Pl74O2W/wjCxh6/KI8vW6EkdHSkrLJURxr0NYaeWBSHuCvXeAvatdP1
YSpZOl5WkQc7ceDWKjYzFh2PcM53icdr9zbrig8DshOd3FxzZh35mwnf8v5bn6cT
wL74Y5CiQzUYR2MYLrvnbv2do6upDdsxkJBDRZsAPwaPtrD89yre46lI2dyaiVX2
+wcKdaOknOqMwPHXLYUizlKgkbYFT2zHDyMsG8GHhG1S4HlDRWAXIrh4f6gGD97q
CLyor7MHgV8wrDZvu11DeK9FFGM0DO6Ed8uLjo7hf+519fKNm8NVfHVyeE9fimsz
BiXdXoCvyqM6YXLOsf2r2sLotUOXsoKCuZ5/tAQpNhRCYnDM3iu7EstagW5B7eWn
s8aq55g2rH54vjnLMFD2bfM/UYQXh47uzlQpGdETj3XfoBd3khQt75dvFuLsZY14
sfw+VGDgO5VPWZtGS4+rlDMZ94HW8DSlSPATCqIn4tXe6wK/pMZtagqEKBr7qCR7
KjeLuKNtMOnByDiG7tqiDPcHCF6ZnTwMe930hhUan+0B+H0RMemRP+MnzAxPEXUb
1CXVCNpJjDqQM0l44wtwes84pO5r7C6La5HOcybAotsqdjk7sS8WxPEKoyIwhXde
JaePVxyrRlaFzb75lCbT+A==
`protect END_PROTECTED
