`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IR5J9KtlkqrW4mZlQELu6aKC/0+ekgPaZV3edJDngRA5Fkg9iBL5Xbrtyj7/cr+1
xQSeF/K0kVqiT8YMffGgokdUj7Sjwo4yfydkxlymW/hNSEMrI6vvOPA20ShNE/9e
7NJ65r7wALgvhbp/EDAwKTAdEGvnm1oVrSYPrASSUVIkQTnWHAHCm5j1O9erGaTO
`protect END_PROTECTED
