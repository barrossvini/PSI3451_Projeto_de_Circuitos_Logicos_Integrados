`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eoaDduoTrPyT44PJFr9n+nVY1WyRMDeIhq48OSbzZi77IancKR1oefQi3FE7ZndH
0E5zCZLj+wlCrUyBTEj1UWm+md7iLIGLAhB2AOzI4gbqA+xFPYJfM2z6Hzyw5bAR
uoGf9G8ARdMGBApXSW7njyr2LHtqnj5XAYrf14e9oBE5yvilJjQb3TbVSzV+TkNO
sgjxE02FJ+lGAX8kVT5iV/Tf1jkVdYgWi+FIPhrZY0UvFcW8wLB3coeH+LH5JgTP
UC5HQcYIo71IUi96CnCILizaLfNr0W6orq8CUqYe/tFh36F+0sHgZ67Mp/m22jvT
IdRUfeXmyyq9zPoVm7sxXd7CbvmDsPxDZTOKxvBa06wTPfbEyykfVoFFrG3aPRZl
r+i/nYYOqJouwUUwyz0oxG2Fn4rw//IXPYwa1YLGyA3ju8CHNupk+L1vTxfjqROJ
+7QEsqdKWzYwiYuTgyvaGUzUDIdvRgFCiEKT8VSkeEejT4N3yM2nHHXi79xZbHRd
3WHe4/WOU5EeTBFA6fXTZ+Eq7K8CerwrRk+e+915xcqN1ZjDdI/Lde6S5WUGVwAD
lMoeNtLRwxf54+pGmD9kyrGanlcPbmIRjWQY2K6V10VB4YJgv1wcaeRYLnlTvVnS
iKUR28sFSNtGBdpVIbnUgmvSNdzerDl+Xfg9/SEjQ+IPfEiVtBDx1jFdfwCvSeRJ
JUN1CWQ9xb5fSYOMRy2Fa9oEyyykUvpD3oQ+F0TgAd51v0Rjyy8Yg3mTERk5IZcN
2uw5Af2FG9OnIaC9TeCcIEg4f3lLU7BG8DQZ3gLyqg1V5HcfKXGHaJIfbSdAujwi
h7zwTOApMfIrn15tiDCbylwl2jYDnY9f+Y1T0LTcOvxgCjJD/GqF53VFFpR7jYxK
lABXOBn7HaDutbfTrLYvdI21vI+uThAyQ9WX52a7KeGaBHhh3fLHYyVPDZYdVgbq
x34JKj9FcH+v2f1FKJp1vy2WDmBaNw+SaxZ0iAaPH4ySGHf/bOUvJmpXpvVUEIXJ
gBWDblhlbxvYpOAIEgF18FR+oX4SNTSw8yhFA5qLHgjdakDoLaAzTaJpxY8m6KH1
j4ifRL05YqtskqfRe983gJehJf+k4GfEOWQNmMzlQVv5ZEuGSQunubrbH8QtC1bT
BYBSbn90seklMkcw8PJyWhEIomDkw5kdGrT8k4XiRRHCK39gqpIY6d9RcyV1l2mt
C3XNxOhZEw4ln7PTkVjgSxAG8jxsOWMBPUGdloBdsdqcGC9HaZhZ0TxmsZ24FRyt
1hQ2+0YuAfg8/00GnBMO7OYQeMknvZ02PWiPnRbGSH3pshejUntTA4emgHwNc/VJ
ajiUVMRR1XwTdKoUHQf3RWs9MRJx1sj2MV4v8zCaKKnFBHIokJc5F0GeR8+wlxK2
mL7A+AostSdUhk8aJpqJK4hDn7ZLMt3Hkogvgc/jOVuyYUxo/2xbi/7K+STXIT65
7wmZy2Ngr0tOXHFUDq+wi8xJSUEj1/UrSFewf9+o826p137qe03wsDQEc1hb9mc1
zcYSLnD+cuVx1eMlBXQgyKSdFiBEJI66mO3WZ+aGfAzuSUds9or47VOJ8wsS4kt3
ddFjXUQyVMt0aaQ73vKO5vkZVP5VT5KAB8+i2ktsKg3BdVc1Hni6NMXZZcGF8vKF
trwNMsV58DVw+/5Id2+rORfkkvAyha2vW48eFIeUtuMUHadP37fjlUrw6zZ/Zm9E
AkeQWX4WMiQGZUXPXMTVMz5KqR9CAGepL3ftM/VRY9RMk7TBnDGGt1J87VVi8WcW
r+BII9HlTEH+l2jSYM2kkA==
`protect END_PROTECTED
