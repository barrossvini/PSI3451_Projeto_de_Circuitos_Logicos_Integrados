`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uyWHm2LYMCie0daWfLNcsikEFmtqRWtBS2Dp3ocOToX7DRwCrN2kxPezLIm++TcH
rlP9gtStsiVruGSrQVvin+dHvLcKpapKUdyq6kdFlu7ysbzg6tuYWae39KEnRhnn
xchjmO4XlyYSMPMTWFDI//SmPqUYe5fFyd3sYf+tHJu3ZuLM+/O7pNIlEe7Jb3Wt
C2MKli0N06yeppBKYWZ2WigjkyKZSQaUMQRM8GHM2cVHc1yvlSP4h/2tnlrj7o6D
QYV6KIDdhoLb92jIGs2tZnJVtGxTX+u3iP5HDYLEQsZ50TJnsOdWjcia6pMoUXUA
ESGGPdvAgVTNlenmCysowOwFoYnak38rEcyvoVSm6Jai58bBPp/FMkzCvUF0aeTz
`protect END_PROTECTED
