`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vN/JJxr5dkEivjpQTw1XOXYHQQQ4chHb5KhPbudx/IZgEEequ77rNAixqtHvzYHL
BVlG9xim8W9A0cOLE5e++jya5Q+dsn8H+HloygvAiky+7qIbQnlEZ1+Ij+X9mqwe
kkQG0ZXuDyWfnRRtC4nW8ZgSv+T8GFkaYjy64MdjeeSyOddLoqdMLvl/1siatu6W
cw8iVkAcC8lujnoU4i68R51RzyyrNxJ6PQYw+O5Ttmx2jekROUFMAAqdiqn5r3cZ
Y5+UZGCeInFHlgwZqXBqfORCx6c/4kphS6QWoI/orZkR8bDmJEq0iuJAJSJOr75x
8OwCsfhrystSudRojoOPeMImvPMy+hiksDqWQBHO1x3ItXVj7TT+etfXjtQOZ8O9
PbPmcTrIF8QuKEONV9+mO8FKbaVMgGnm4LmgfbhHN0i32eDFT5uwHwd9fdOOYOuZ
KSjIMwAv2ZUj7s3OZ5ttaIme/qoFG4bGDKE2/YG5qGxXZYmcsQbxzW+4564n62T6
z3/K3lCddzfR30ZK27qLPi/FrCyyMYQooSF4EXwNuu93Wu2x1OykuEu0dsC/uxYG
FyeRP5fDz1lH0CrFHhZ0c4tDIt+4lgx25A9NDi+t2D3frk2dSmqUc0bhyUtEV6Rx
nf/Ha7hDb5HPhcUcweCUJYugfH82CTGixyWbgRPcxab0HUAkzdd9UzzTmPv+bByh
8F363hmpv78J/OZLRxGUy5d2c3zt+UCF3askxz8g5Ylh/3ma18oSbfFciXQb/u17
1sTb0jBq/dbA4gDYk40rW+LpMkKnP46GDZcdkCOnlabo5eJueFo99Fg0J3NCVOEG
Nkz2+Vi7pnLHAFzpAtaNnTBrM296il1I0ql8qIXZHgmr0bb8zjYvoZitDPNXgK+0
YyV4AkQeDA1AlyelJVqD4Ts89V6CYhFpcXpCHDHeef6NLRig2bxwpB2wXn43RDUE
SrS/etYZMTSHmBqcNhblqZOQdqQHk5p7W55eVfdMPwucBerrYCVUi837Uhk9cIdz
RtFNJflnRjeONtmCCdvoCwroAggxABlg4cUKxtnzkVmv/ND3Qioc8HnUrKMs0nEs
Sx3Abrv3cEuQq/Tuyu92cvDBen9oLwlSRxL8ZnpAEvA=
`protect END_PROTECTED
