`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tRjh1ajY1kRJXDJprc23+btApsmwsULY6MEBpZTXEL4r7M0hHGGVabNXXhkI76vf
1Ps4xNhUrUFshUiBpiSUn5i2gO/TQSXoXzxlLzfXlLtRckUAza6OWyfhCvjtCifA
NjzCZ2moyjORm8cV9r8rIOkDn+BC9RW7RWaiwP1TJZUjAZIAmnN9Ppkz35Gp699w
onb1UBQV71gLYIZxduL+sEcrtVyELhWu22uuTaP87vIEJ4WR/qt7E0zvrAoid77i
YxSvQPB2kJ02+/CaMtztSAetL70Sg+MfNx6p/CZxi2ueg1FQpvrIhbbiHXTTBpIk
Z4sGMTy6oUgqk5lWK/CL7CMe33x7sBwtbtlTFrMWpyTlHIcaia8odCaehJTAgDmQ
eT1armRcWOkIjZbJF7wUm8FjoYw0VmG77PxtMCmJO0mJX8GsJdS841R4FX51rRss
mAl8v7iAULXIG7ampW4dBAZlEwLdylWfqTvB18s5MqWTDFvMHT4Ne1AUPdweSGbN
8auFQiwc/EzaQuTUZvRGB3YXw/m/vTm1k8mb7SjfFnNPOIY21/Q+S4IAhyWV93el
IK8qXUWkydMTwRibZvkt623wduP3uPw9EHHuLedoeJpCyY/jr/KFiMQscWsIrqBD
MtmPXUIstN8pctp45qRlv7zaJKdIazzS4GNO1gOJKJXevzvf9d4D//JOllk4qiO7
iVyU8NVwA2EtUbLSdFol/c8Hxqvwk5GGKZj/IVyK0qWNN0d6ePqa7LDT0ISBYb+0
r8/EdNddkZIN28ReCbLX1EMC4qCCq4hTLYyCF+t8OH40pjxbmxE+Oo3/rcZTT3ii
pSQ6PUMj/zMebf35nplrY49rfbRFfx0T7MZkNsDz3maQXeLZHawhJxnwvDnEUxUL
lrorPu1UglGSew8wBbtHa8m3tAXsn17WEyzmp4Mfm853tCWsushEtg140tHizQhK
gAf1dwBVySVxYw6VMAlRPQqyLw3AW6C+VS+0gyIopqqr7dz+1/MbJNFqMsZNphv1
jx/T99lkjxAsQOpkCiFpKf+Xck1R/zQqXfvK7ahvsw4kR15DA5RifBwUb74dmnnB
0GzQRbsmgmWb+HJb+OncWpzD/flFB4paO7tbepinshB0oLIKhmfirXc6jWZtR1hv
amFgmvQyQGYw+4uLspSEoPGOusaXe03Dtle1QzvAk01n3TAmE+2wRMeHvrBvMRGh
J915LTmJ8jbSChfpuZDVcxYIH98Lue1DphOAtKccK+Tjb6TYJk6yuEYHk6aJj5A3
MnIDUG6WPaAT4MBYYeRyHCnVp2Hm2nUsta4aU32/Fb0/uP4cmVp0YjFzD6uJqNCR
EOIUo8jHwoCRZkA4rYMRFv44rmmh0EMe183HsaeF6MCvEH+I+WbwuChy1bpUuz4A
4QxmUbzrPX5awc59e06wPyLNXR4Pf2+2drCtT4VcviTaGn71IyWgb0cS0luDhNzY
voIzETJUBS4QqpX9Aao55P90I3qHkkhYeeggiMsmM6UyHW7NrsF6jnFxGWOgDC6V
CebszuQsDUWkrLomSh9SadVUcpE7IYNrW9pjpkpjFv9TnlOZ07As/IDlmtjaC6nd
VSyx38Og3VYXOE4MpFq3BjrjNRWcqbqriHn5D3t+gxIt8Akn6x1e7pSIHntTMBi3
XPtkzRAa+qnao3+92s+esmHypRRdJNg2NkgNT8BCT5QkghSPOrevR2XNJL/1g5/p
My1UabzQS6kEn5fZFnqciO7R7JJoqWrKndyjA5E9kWXPLvTDVEOu2usyYZ6PSsiX
tfjx959AywfGeNHqIw4K3cApjcOj04OxEK9K4lfXKOVxvQ2om4ZRetoN2wpGw+1B
BYw/sjHSPcPnomr6YdJ2UkqKWxJXRo4OZWrcHp1xwp5RWCqULzb/IMu56DeWhE18
kplAL5Dpc5r22/+h5TIa/4Ag2+x66JC4maetSgKZB/dqMK/lQ6Id0AaWJZva5TSw
nVGR7AT0SPaLmd9p5W39gL+rIUTWJB1RRy0punvoCjnagp0zH6VrztLKmFSBmFsx
6mblTUg0Y62cQ8kDJ5lgHJz2eg9Fa8WbKo+N+zGa+1OdThVRC0jd2MZfjsIt1lnU
YSt+By4RYiDdO2kCSehxFKPcgIHvyZbNmjNBJ8vgbtWMIM0rfuZexZSUK482g45a
CZN5yxVnJk4A2167lKNKQfkgPFQ+S6yV8s37W+O7s+ow0oSQwOrLpkPdAgihVkqF
D6DetqpCWISdItmFqQG0HXCQs3ONFTZI3GaEcCea5pQiTlXRnGGtLLR3SVSikDEm
Dwz6/FrOFLRQYbtZegqvi2Fo47q4eTLa9b/T0M6fLq4FpUvPlLqPsSVdXAgpL4zq
HwneoXQADQq6veRrFjx4pj9qZ9uG+FJW7p3Rv+p0Jm9u3rFLoGQEM9/aRVKwXyis
5Vl57iXbRUJAAnp1rZLtSUzCxeweuiXpYEi0qO+mICmUjN6U9beTxBnzbbhrc/kK
64FVr+j0VHqREAkQdq0MHAO73ffLOSwvJzFru9Us52EsUa6PRpv1p94sXapQVpMT
VWg9SivW9S8Xipfg07goGfS1Sdzj34PXKFpa3cYWl/MFKRICuMN8r/lfHXqJmh0R
hlJZ57/zXYwHW/YEKUp9zMHihi6voyangEe2KIUM8HItdAjKYUhs1KhS4BY0lma+
vlhvdOyvym1K18IpxT89hxgQyodabXOpc+rLGZ7OutWIkrf6Y/gotvgCF16mgW0G
XznBfpJWEgDTqFgYk2gTncxIB3hb3q6dm+r9UMv4BPOgSF9byaL2b+vcKmU7Wlcr
9goJdOt6ipA5DS316y5DnWMGW5STd2bh0fB5RR/FHxQHQTCGf0R5KZNpliSY3WC0
6J9tu6K8rDhKJQH8Mr8XGIhc0lNmDOHEAHw3SBcFHQN/TvNamUhqJMu+b/Y0dSO/
j0NgqoUTe6rkR4B9VRYrIBLmdM6XDAWsMJbdxgWwXjjoNHvyZX2d+rFm9HTXc7ee
zo70tPpmSF/AQ2Eh8ibnChHQrua+PRtdg0FEo8WlBi2ul+TqGF3E28I5hySZNzGR
N9zHCq966cDD/ats9Bihr+h+MG2qJORYmsKQnSfwp9sWsKKSjjr8roOpSXx+bJRI
PJLQz7zbRcOHdzuTFLO06aUX61qdLiy/X8hqtb0aaFajvuDvguVJtmMfTpEjsbF4
yl9J0Y1OeMD0wWyDwHRvRcmMo9vEw61V2VndbVggXKWXOqKPK2m+d0nRFh/9jtkZ
xj4czW9Zjs7dabdDUBEmWUrzGk6I5ywTwQ7sYjosYu3TuRaQu2+Q+zS5xeksJik1
nfj5f6TJNXQ3m2AIS8JltU6/mtEV0w7aUUbk5gMnrCg0AW/hh+RmXMnk9dna30yb
KBDXENht2qotfsCnzwQnXPcnoPjOLY6aOfQqYv/LQzI+/2n3a+bVKKvAkyOBsKZk
kCaCUOIt0x4oueep/S35fevxD0cA98pLJ87kWnA3Gp2q1DD+OBFwEn+t+QPB8Gq/
EHTGWkLNFG8Z2CvLXnIOJ2ybZW3vbN6BS4EUaeA2P5wj/FeUlhe/lqGhI5190BKd
hd2d7rg6DykDa5yAHzIyphMeoxyl89fkUiToJTjzo+dbaPvkfytkSXlCkyzQV88Y
JVmbzSazktaDddGCvfW2EIqdZJMaN+SBp4xdkZ4PCv6sTUdi/nsIIGL/f41ed3zM
bBR8oFY6q5DQb8eNyCpAtQ/yUpT+YcGuVC3bLgmAkt6c9xUNxbe8gnCOTnsURHca
BbwBX5cX9gyVvK3mdUXlbuzoqgsC4L7njonF7/xVGoiKNgKAEavU3bO+54Phdriw
DOpvcCzsW8T9jaUnqo7HCaKvUYZhxeF1TJOR3MxaHbNjk5P+Az5wa4r/SfBxYuRU
3e3U89+62evm720+Rq91X276q3/xawCT13Ge90VZ1Yl2Opb3353Y8NMQtDnsFoqc
MOcQ1SWVkrA7EyuY8bBe99lnY06vQz69Plsju/zXuJcIYefuV9VsiH3y35D6n2OW
TMy9O8Y/5xYaBCnEntTeRL9bC1+dzNCv5DXsvhUq303ABkEhs1xv316sRkiZ/Z+1
6mEhLukQlJmiVwzvHgeqJQsfDIatmWJFgTICyysOf/mkbMOKMLbHheKRUwQjo0MK
4BncFOTt3a7OF60cBP5GaHkFLeWNw90c0KD40qQXRh3eEqMjPbsMbLyWWdYQj27t
uSgxcn+B+Al5Ecg+0j/r6KNO7lwI5d2FGDhKW5ZM1Q49HqA75jG/2DB6fc7Nq384
3aDfBlXw6yoF59dAuUcm265J253bRofy2BnX0bBkLaRj+sd3kq7bba2jxTNbkSi0
30irUsxt/8GQ+flKDr2a4ic1dd6vez3RLnakRjjqsuqnQRNMFNRf541Shm6L91dK
iOkCyvHc50VHQDDm7zLIY3tgfRVOru41eDUrcNksIyJpgJvS5x8MrZprdMDXcP5g
L1F0qo19DxQ5XNatl7hT4ApaG0RL3EDCP1m38kpYm5WTStwQYqiygg1+Yj9ykKnP
ZbfTTMxqUuFce4NK7VQhigqUdFafM5Pw9nRxjibigI8z/xc8WXAMC6m4+NK1qHQ2
N5VLWH0ZnVkpnMLRuetI0SUn+ZW1EWwZODAZY2cGzPJvvzEvoMNtvxEt7hxrkTan
ZeNHK+KnLSmTai/49TSl3gijnxJiWnYip1rSguX9vc1Igh1wdzon2dQ+Xp4DYBEo
EJ6S14g2QpmhiskpOXGTH1+BGhEF2PPXmXdW0JiP9zJjLdOZTMIDxRjbLeakQ+dx
UVVxPlBbeoHIA6ivlBotFpyxmLrOA2sQssqGAaWgI2+rQfsO+O9fkrlmaBpOUNNC
+nMI+OyJwzQQuv0jPTvPOLJxt0BfDBtwPtF48JAfIvCwQbp1IbrIqYUGCgxkIg2b
WFp+EDdesHxzTIo7oXdFZTa6qPA+qW1BlClt43YXgCJbuBwYd+dBYpU42CAbFZbl
DrudjYfP+4pKVH3IPJXqmWSl3k7aa37l8Vdwg4LMlHxCrrRRrCTQ/Mt+p94cvf0k
xc+E655bFRe1MnBZnUJjLQ==
`protect END_PROTECTED
