`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XCJGTgAGEjXtGQo01NQOL65TRTieFlJyg2NdGY9BHE5Zb5ZKYSlrd2u5MYr53zzy
sQU6BuLVXKudnT/5fIHhGAtcbfRfq5OlnIZAtwXAiaHcOC9O2RMXC1zR+QSb6Xp5
QmkTYNXF6GB6T5oJsasPeFyKIomH9tGQnBZ5APsA3JYWEZxzP6arl6A24MLUstlg
MQ67FXbGDnXFpWnCjiJeM2GtZUwtcattIhaVb4HTI0g9/UWtIpdONFrqqFL+zVRF
vOOyGKsd6ldbRUfid0Y4i27SH9kMo3bq1MH6XRf0vrrNCZ+GPY9ORooKWxV8WULI
pS5aOQJRvf0XoKuEWxxpuDs/L3EahOPstJuigP/j20Zunim052fSFjrmVQlDPbhg
dSSaHJkEWBWDQepakECGo2G/4Bv4MCYZnMVvo9tpmUP4ROE86YWUcZqrE6QPcCC9
cfx4UEbjDqsf1q2Hz2/gTQ==
`protect END_PROTECTED
