`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IDjt4QYJs/hZCMKppurHB1ulprpFUTgNJ/D6RMnuGxyRPdc7h33EmAbQ1m+P6TVA
fJ3DJWzQs92/tJOFzySFs786FywsZSR+bBN/5VZYxi7aLffjnrDbLy1HMLM7NbHv
P2dX9OZoeXerKnA0sUJkXZ0HnFotAlH17eDnRP/OUoNUEIAsfpCHw9I0JeaZ1ISr
Hh4nj5XJBjLGMZDsyre943jvF7oxpRrW5gswTEr8p7MPLqIN4VAzmnmv929VMSC2
kHnvEKC+ewLOGAweVrLZUA/yBHSDdzJvuF0Y5Rvhcw4STxjeu4acJiLwzW3raYuV
QciO6W40Dongdmh5KHVM7m3AqLd+yOV2EBNqDvJQm63CBz5UvwuAIE4R7fjtTq/5
Kno4g+5/eHh//1doM4gKIw==
`protect END_PROTECTED
