`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kSlodoZpdOa2+HlXugV7DtsWAUZftKWzOpv+lwWty5Ec0t0PaAF4zCRVwE0lg0EX
hz1s1fvpFQbeM7Md6GW0iHgHo/O9grcLf9hIMfiVqq5muWT96+VNW9wNPYTsOu07
RXOCD3CxINtpMBXL19+haPyvtUdj64nMFzRXJgHTMQHfIQzpGl+0itD6fE92xQB9
Ey4DhlQUAt0rQIDWZ8pgToIPXJhx7M7N0OkDNJZ4toOn8Wc0flCBu9guxBShpkk9
jhE6xdUBDU1XMUp8O2KNkVhA3WF30HNrkDsdzB0iZbitNSajSwg0+hZGrh9inDMQ
HzYBNPh2fPclgnWNyTXxYiNJx4Wxl5U7LkKJdvLLKII/dn+A4IiUYqpndBg0ejn9
th+QF2eTr0/bx9ectugjtZ4Im+gTjb+kfLzDhILnos0O7VVBTXSViDnM9bWPXnK9
a6ioryq0TAf+mLEUDAAns9KdKPND2cx1F3tk+UlWsqmqb+CX7d24rY6zr4BUcXH3
coB/vpVHyuoOH7c7nxHACFnuoklw0fn9irCRdRMTX0cQgpqvHvX9mcwhOk+fBDDZ
c1LA4G3gK6NYpLew8gXTNv/Azq9XRvMLsvBpFdMPYqbzHRlcx4voZSyg7cOCFB2x
qC7Nt53v7wA4jNeOp7Aj3nJEfczGysO9RQP0US6n4nXJ1uMRCKq7bLDjjYX804f2
zDKfHIXb7pxWsuJmfm3bFprfM+8PMvoMpyoit4fnnGMP2Z8Y7OLa4ZZLeC9yXqcq
T1lw/DYG1hjNA4+OTk5s0S8vT9HKJy8b7AaZO2oiYoBAZKKM4eHpT2sAtraemcku
9iZ2weoLpejNskfkFW0P5u9BZOuwvpu/kZoYGBsKTEbf4sEbr0X/G8mlRQrMKMEy
JZ6KyibkWOMWOvvYZl4JLjsPcyWCKaXiy3Vp7YL5rr8EY2ti50Bm55qHo+WV1T6x
mFsoP5IoqBP9BNJRZhYlQRT9zc9i7Z+nhHFxSoI2IX8Qoc6usRs+XTAdd0IN5NZK
UjFda3b8da3FxFJPatHFOT6akwwnGHqZHZPRQWWO05Syw4b/6uYZ2qwlYdlbo3QH
+h/wEYDKsJAMMHGXeyoIvPrktjwiNkFMEPC+8ugESD9B0ix7AEvEhL6yN4c/lsLi
qVg02Ik2okJyLsPdvg5/fg+1XSSCchyvjiDNMXpJDqA3QPCytHf5Bw69MRSIEb+g
IM8ISA9YA9jfNrYC1NnwuJzZURtUDYqCgxb3p7sO9SIq67vdNp72KocBvC3+YGRv
Z7eXH0gz3emJ63suQBmQJ6nCw2NJ2D7JqrCbzoDv8hzkoKlNPKxrPzL4IrkqXfkP
sx5aWIE85GDAFUzSU6WWqOpUc6c4evlwzSCDb9owQGwBmTz+tcb4zddPUvsgE07H
MGJbYzWi4jzny6uEAzTqJ5PARpwXDLg52m6g9gh33oUUuzbiROGdBIA03uG4yVkd
bdxTUH9zAMWoaQXUpum1P6RjO+T3Ome33vcwKvCUZ/cOEugkrPg4EGVb286Dkovv
GVN3WvR92o8NurPQ86tsmEG3Nci1MZI76SkY/pqaxEl5r5T7mOw6Z9bqcTm3Y8vH
tc+1A6/I4/CNBwktIq1gJ4igoRsGtTtyRsmruI4WzjSkhYigu1k9YrMS8HwM7cDu
4+NTY6T5mhFBzPmIznl1REn7FLW7+tLINCprh0+xoHhIkbVduMa6Vqe8n4cCPqbX
kOS0KhtTFOpC2cR7yAacLK9syiQUbUsZccPejoBvq0rafhRvvl3eUvrxrbAYqMGV
Tq/k3TLng2mCIb9vizEjNOgZB9NrAxd7IRSARWoagVdnHpHBiFB4jEvCQ1f4FZYh
CXzsQGDL4mOtv94//cVjWAnpDYodlw7O+kXGRJwtmipbRbSAb2FzReDi414WGDkV
uxrL1BffMRMt9wui+oAGw97rBbeLtOICu/eR1yDS/bpiMe7dqMpWEN0PWcbdwS6r
C1PqtxznFrA3DYbuaSmqKH99CMZyebxBydPsJPSgYWQmcPAg9qLiwRE4x76I9zTE
BfmvJ0ItcRyKMHY/HZNPhccjj8pgMAg+c1l3jgRkwHHDOauss666Wy2kJvEKm9vh
zJXoDvpT/mxqNNV+gH7E+n6JCJpijrMA4uEOWL6PHkoqmGmtkksFZJwmYU1Ue0+Y
+OTbK7oqqf25u9esv55ynI4VV2ixpXhokwZjSdEDjgHan4hbF80pzazIyEh7HuU3
1l84LfhmlIYQ7E5xHWzHQ0m+C1NRwF4WgbCsR1985rFSwH/sOtIdiD0CV5Jd6KMY
3QwfykqaWf0Dg4UzYZsM61wvS3Jth7m75ir8nwLKNn8zPsa7YpWv4rcBz5LpGgxD
c4UvGj8aBOQlXdr0TcytgRhgzzKz+ykr7zksgaRGHmpJCSxetwIOMhRFS5/7J9Vl
7oIKmFz0B/uQbLxRkNX3uJCigbiCmc1Kq96JWgjN6LTKPomGt3c7mY8W2CZ3pUpT
rXLzOT7YolNXmbn0pcWp550sIsg4e9UeBFF4O97Hc/CselgJCBOVYWVpjJEenEVs
oOSay54VQ9bbYRj9+81w6jzMk5UP5eJV9yVSt0zhCn9Fh90/fmcH6iBUmNSpDxQ5
6iLYmFwGpdwKGQojBvv3Tvkhyjo/diG/cn4wZFg7pOKxxZZlsDHLNOx0hvym1BYa
l2usDjyIo9u6RfB9UmlgbobpwCiL4wPcuTUoZ2ywU17vda9FXXLa4pFqxNZ9+PEL
oBUwRKevbNwvDikCjLjPckmXdeN5WihQjjmiUqVuXiktnt3khHS8wYP3USGEESjT
w0PsWXmbyDoCtut2flQNAZp/H66TZcWcpUUNQyM4XLIdmrWsqf5SbpZvnQT/V9yI
GtZSBmkiqmLC1Z8qf0660zN4Eqw+88OUq6XBmQxlHywYLce3ZsDDtZqMiv8xgcAA
5RE72t9VAvAr0jaJArexFM61WU+0fRkYYENxXXObLcPDrIbVWoi6JhtrV6Zi3Kb1
wm8UgVXu+3BySA/1fxj34cVJZxzH5S+hXLER8YVv5E5aVB9laWeP3Rex8riR0OaG
I0CmSy99v+qKOx6pZCgRw+U8HfnCzw1zc3Vh+S/gEeKbKjBnmK3fS1FvKRgHukaP
JW2pU9YbZiSIHctpuzzu2w2cYKypyDlfyQNwyHbV4EQPHFjtXEfZwpj5wLyj9yKe
rYh6x6t/IgHqBeRY6KTSUrh31XipEFtkV17t/kuAhdsqLUmjBIais4WbxFr7nD5r
+ulSCjoTpAX7QGDUqN899NszGiSrsaa6ry7/lo52v/iik3qrzWzbQUX8kDc7a9Ta
bqnRNK7jBWZsDzl2PUkzEc4QkZCqtuMuPeApV8ZwlRq57KcfO6AnZcb7OT/C5p4m
tSXDSyevrITCBMafkHCDTTDjPoNfljsfBzoG6PhT76KRjpY8KbDjxi74Tj3sapJD
XA2Frl0lRJB0I6mxLTOULATOxLJMd9Uf1Y8LbNR+4Q45QkkdYZgORSWsV+qIuTyu
i/7X9pq81Lqo+Y1jKUnGNBCV+RRDtunlP6Mm7sJy2SfxQC+F4NYvrdEGR2au79yC
LvE5AtBCc43TABk5RRidYvYZajjIZRP8/cDOU4Bd4sSIchVT+QW+Id5vqnPeEKS5
iCMUTu2G08TWI6PxcTzlrrWOnJflJeokrw3QirkXAQwTjsKv1lAjE3JyMEcVGqQ6
rEFnkSt25h8B+3j1M4Z0Sg9sWgZxwW4rMj3goXBdirj119IU0ryoUi8LPZG+ddly
XAmKheg+0c/IqOt72M0lpjvKiSCxsef22UCrbRF4OaNDO+uJ9V3kTJrMBhAhKDOt
81rdb5/3HP9bdhYlZDtjz5JLX1BgCBw/PMrZa1hVHZpG0SSdN66wO9QiSVkCAiLh
WBiu7xsbzFaLpqk6l4SQ59WNLKkfiGkvgDrSg6WmhhQtE7BT56kxR+Xot+PoLtHS
4aGOrf6TUFtk4yGeUax2q7HDsgW2nqjmheRqM9xVP6tlG5nHjYf5W/6JF39I5T5H
OsGj1uvaBzt+kdMiSnvhH7QO0daqGZa7fy463y3/hKPNKomEhuCJi7tS7T45a5eu
CjbYQRwGz3AgROij+7OS9/Z2THHeWSieHifQAeWrus0R48XeFvIrerxAY+aE7VwA
WGnRgwF0pm0qwY2yn2UNxWUp1tXftOxKIG4j3C4L/mOco3DsYcLOUJRg9SwSLk1O
zsYy9SnLOcTOeFFQVKgHsS4I2vBWnacyL3Be2paaF6/uwTowX1Mmd/xz9Wq8vrb/
668LGJl/AaVntKvs6CYNFbsV6OxOXdlxXJ+KLbqAGMzj8r0mBoqL03VKfwsep/iL
oul+9glmlxpn69HAcnTuaXO5yowBGzF27DIAVADcc/XmmljhrmTgnvYjljkTQANX
ZBYo5/qv/lMed5oXe/hN+QspDzEJBNDV8PwNuCuYUIDevPNRFlfx9hdrIEsnKGGW
3U4DqH//W1NRl7ohdxE4AOhPcPcCYqFQPO71GlRo4dcXQXIEab5tSvsQnaEZxTPQ
74u4boYFBkhaTOl+Egi28eBmKkWiRDzoLxfmLJWnxFHWpILaGkAjYjfO5wTB9qHC
aD+JZ/o3wW9lJk+MviaIBcyzjTh7DuODYbB/M+CAxb7fq47wW2N2oBlFZtXd+6qy
s3zITzcLxfUE81obUoLU1TWHgM2OHspsyBFDXtgPOEBuTvrgUW7m4+agV4yXeEUh
jhlgBfjIBjlg65QSqsvE20UXvL3I7nK1PI6d7FFsWdnU0biUNWLqcCw9FeduATkj
gHf5+ApdoMOAJVJMj/mOFUJ7/gH/YtzWzbeCG3ymKDjQRpMgAHmhu1egkjD0C2nZ
YO1RldphpGMm1IkM9JHETdxjranQIVnUTsMW0B47zYKXewwGcxKCcx45L+28PRUa
eUjOKcrPeEnjTGp10JVzt7Q169yKcIZvAy/bJUL0Da7PRGgk9PPe6YwYqJpsoNVN
CXFIFYg1jgf0hhr3RrHClqmrf8nDtbtXudIMeWbX4E7867J/jDc6X/Wrch7Oqurj
NlddHPGYzbsKiel4uwjvOjRhy5iz4Rj/RsrQnIh+LmbVMQRkbhc7cN5GDHAMOakq
7UJ6rJH2l0voQx2HULPcKyd9f6sbqbIFZfHFTc1ldIYxJmgtYMCikNphnBGqTBdF
FsJZZxj+ItngG2L4a+pjiIB3M2Yml36k6e1C9zY1ixJuGf5mRKuHFYrX/wdXBjQd
JSt5QbLiQzJU+N0KoB/+kM+rl2Uzx60XADN8WheX4glqOs4awWO3NdU3x6F6t7rb
qA557qzZ9FmR+P2Cm3TwIpvaPvcwAbIAPReXij6WG5WsiuDeEjqaOd5vtvd+7jC3
QtNEq/kiAjfSnmrmyF3es6YBOZFAo2Ep7NzmhJdOGcivxD6i1SBAbVBICofu64hI
U5EssVeDY1+a3UgWMwLEztZI6whM6fOYe0mf+QSkw+UcTDncNVsGPkuAlanC0eYC
RG+pCYl0NtPJdmoW6Wg4glLKUCxCC1DwjG2JUITiyVDV0L6AJAWh2rOXybM7GAAu
m799Xezd9W3VhgDu/r2WSqyt9cUmdxmEByQkaKKympLyDh6MWT0XYNLY5ZljtVHT
OtPFoQTFZ+YY+1NPa4MsEa+8fl5ac3zc/fiuZlTc5eTDHVbvQDQeENcTltNEsjWN
HMPNQ88P2J9VoNim/VaOG6NoHexsNvMMIUACJso1N0PyJW5+8Fx4gDPwx1w0O9Gy
Nv/bty+sZ4obdpTJZAtcyUGWrctExwVwkAtIUmtxpoa9sxhBWlevtml1t2m+kUjE
A01jFcMIK1sQhunSfocL5L8QA60j74RM3iuY90Gp/8+IKaFCxiaEjjhHuGw4Eg3e
/n6Zu2ktoeMUMT3T1bieYZQCngJpHAFMKoU6yOOdn0CBj1uyIZsLUGLPmAiBc0e/
XwhVIuYU0VtO8ClPEEWgcbuerP87guDlPaTPXmrG6mT2fnyRlatySCWlyJJ0iocc
kj/2kETiztqb/S99ESrQmW0kNEHYpHdPHAGodHM8gfkPinnp/25+NhwK5yI0X/h3
VD4UPQdcNnfl08/I3g6HbtcpW6YojUiWf9vRBXDyuMfvE1uJ3EElLC0BSwqrorHk
zcQK5box5dvQ4dMErdWnDfA3qIg+uHrfizUQruXSDjVHZvXqWMkCuhzYoePUVakb
GK5tI0Uxi55lt54V6KCAXQTGnrY9PfTo4zg/hILt4a8SGsAfHwYl/qtqvWx2Fqvn
r9OaJdzNjzKaWF6lq5fqMTq3sycU+dhwuffx+21lA0bUmiMJ2m0lZjAS0rIqJ90t
8oS34fRmfzCEHTY4w50vvlCszq3K9+TlZDD9+WLELyEqYXja+BH+9+9ta3Jd/YEW
KcesCP5NQTH+AvzqO4pMq+qJHyfC9cn0LoTMwLpvVCNzVHZa4NfXWpu9VrZ6mOu8
m0qfr9K8b3yUYNdkBBff4Y2LytQrk6ZnuNkoK3vq7HqioAGRAMHOYOj8sKZp5axm
CH8DJb45Yr3yXnYjnkke1NozxRNbQy4B9+9iWC9eSGio2UnBErNq09p8rduOXRbi
ts8SQdKcmWiUPg4Z5lhKCJ3DysEItFI5VUuEM/0C3tidMCvHLk1D/C/rgHAG+6xj
KeApPFgHxYckEK7BCX+9pO1Bm+B6bjAD2zjafQikdjQsODiVJ/4GZEUMrDp31HtY
oqHCLnvidKFXTzlpyOBgyRZPqQPlsKQOSAOnifqZpfMlmPFAxV8TUse5KOd5ORWR
UzHM1tRl9g/4dzVPVUrFvrnNwlw7UITGzvtbqy3uS+16upwvQdQFOlS3QP+KU+MX
KATxqQ7/tyHkxj+I0hHsy0/zGCC/8v9H1K4UOxc5TitwEpjkjQs3WWTRMKQ8bxF4
zxkDDGTDMcjR/Fgxn0XuEsHty4xr5NXE4qIwrw8CYXFKoEyIW6utcO/CfJHuQR5/
FJl2+/40YwmUmHzpQWKd4ovMZy0I5ZM0utjnDQMBFCeXwspJ269v/hf6Vghpmw8k
efLsMr6U7P4l/p2tkx7o5plIsRBRwBsq4RoDNSpdvSZsrWwAfNLgKX/k+kbBnTGn
xKuFOljqxfDhOU35ici/g70FNjh+bQobxDKVEJNV9uP47vTELmh54NvnDU26trw8
wrtSn+q24cbmaSgVYua+4XuMZTDWLM6abgeBImEN1e7M3N5ajdAU8XL9PZa7ViQA
o6XTmrGG5/J+1plRf6KJwFniS4ELMgBiURvEJdmgifxFWoS6d7nYEb3lSqs4tvpP
WPguyMs5NKKWh4wDWP4k9mbn06t1z4t8bU04zcLBWm3XaB56U9sUzDVj2mxyG9QU
RXBAev5HLjNIOsxzarnNq5nV3xTgtndWPAnePIjpQPWqWb8cxPAODlmyJrpK+iGp
rV3pHydg/SC0t4meQSVj59gfo6d3Q4KN1ydGHoReEBdUyyCdoFwVESdglACxJcOB
Okf8/IXjq9Tc2BgCM1knDUZQvOETrVfJmFY7iM5tIdRM0brOQZYKY8k6gb+msW6g
U2hL2oWLzo88v7MkwXtvs39vZIrAX1apFnVa+uozWNuOMXoVDNVCdvV34jCBxFYh
rEGITnnZcS65JR1Z2N5McuMgpPnKpfO26dnCRUFViSr9Tc6fHIhBllgwYA3RXGgM
6W717kgqOjozxiyxyFqKqrj7iHzKweXBCgA68UveJw8N/8Il72dqfamt8UKx5LSX
yDKcou5N2SSPeXIa7Kh/X84JBxro/FHCTi6LuqVWgQ6Bu3Qwfu/vU/Zu0lhXL53B
ZHq7CkDd5+F+rYIBbJ/usG48JG6AoVk/QYcLlHfl5AJqYtKFujo2f8LVM3PgOG7X
GoK18idgbvntD94k13P17waCIMu0WklU/0lTUDCYAEOFt4UPHTjT3E2RaxLjA0en
Iu0SYWaZn6VlMdUNTs8FvAag3cWj4PVJnls/jSPsHtKRgwiWc4QG4SmY+656m9Z4
frt7/T//51cpxCeBtFSeEH/EG05Lw0dbYMHRZgb4AeOeR8uF17y7xzZ/7mEnDYr9
yutt+tS91TPGtpRwNQ7sXyAmmml1FnnD4RNuGdYvtSU7rwUG6l5exjb3YuF2CpRL
0bwcI+2jUKSv5fOdFEV3ezmP54f+eFVdXIuOTHwVaMITW8rNlk7yxwgicIb0Ocfp
2WMb8Rf+6R8PH32Fq4iEuVZ9TRMPFrAX0XexB8NiCtgFNrLcDQhQnP9mxXZWSwjU
FzUinMR42dLS1EX2xeVFsBxCNS5i73tDAUpMv1+OXhGg6jOfWODuL4NIeroCgjzO
E/FoMkcZRcLbWGnlCFB4hnvHhZH6BeGYpbzQ1hV2i+0pRLGTIcWm66534j8AQA1X
tNSMy4TvtPOzifOunPZfO3ZWSpgeJ0tee3tkMqJDwmD33jJlYNNJUrffbRI1BW2N
NS8n0whvGa09lUzN0M2yuP1f/5ypXQUnvKMz7WSo2inF3UXtr6BaWkERKuQvDaQl
qP/aHgMdRsF8X63KKAnB8GVz6+OFo1rP7xvLZVF2e+/4m7LUJcNhCMlfz7drvGvD
C6PtizFXdETY8t2YwyF6FZettitfrG0iXI6FnD1xKb7i0XXl1hS4vQvUn3HSYtve
46X9KdzJxTeBJ17lj2W9ZzsyOvJyJa4CHjQ473iuP7OEtHPzDqCWK7juPWmXa3VD
5qj11OaXowQ+lmxEMAHVfKLMawPWwLV8ST4YLWdW1rREZhETbDgqSaazhM3AvgfK
3IIoxpY9Yq4Zyx8/Yo8gI/8m++w8gP67VlTNLtfF8OXd/QULACWJMDS0E3D7iXky
WY1+eh5n3NdV3y8shBxNryLZ5Wp15wTSYp9/+HHFdeg40ml4xCNlMruSHTZ114X5
Disg+pKJ26URWI7pinq23RhV5cc+xDr70rYjA5T1hX+hcZv8i55GyckzMUTDszmZ
rcyZbzLMRCwGyazoKxomj7ryLZHnTd6sgGIT/IVS7pql3M6mJ5sHd3jgV5aA+BR3
5RlEBptzkLPyGKMrGpEpPEOOehdwq4Uq6R3SFB11SIZykD7FGicAWY2uyCjD+JEU
Mis3dkPkR2oaPgdv62TId7USGTDCklC+Q3aHR4vsX/zXDK5V6dxZi49GicV+dQyy
cTiP1JhH+2r8z+n2YYkzPqHL8PRo+5VYB5I9Vrf+iA853Dw37v13TiNDMa3SRRH6
GVPOMwnQ4FjzaOPYvagNHHyoy8O9qFjlhYRK1YLvlboqN8385ErBRjQF5qTqfrM+
9HOlZBNN5VnwLr45iELaYb9C2dw6yUBvzgZBZQaNkt8Rb0rzAjcAeFQ7l0ugePNf
f2JjVvT3a2jwz3hd7XVyXsjNSGRpu/O+JjI1Powf2qXjTCxsECFju75QM/tvxEqZ
4ub8C9nMxWnfGPfyfi+81oSdizB488e+vri/G9y+ZTQ71kn6HIGHHVC1iq3rLbEB
SwcOgkR0lwyi2UKBuxU8Hy0d4KFLCqITdDpk39GmJcRSB7JJnxIaCAEbXiMLOkyd
sw2GJx7mc3tq0uTJfWuw5hPO68MNtBAS3w+ZIxwT0l1N0W/U/4vtAHs/Kg8vlAom
L3Iih/DAlJ0CAd0zmyIZPSKPAUVC+BTncWzE2dcyETvH9Eje/IDQjx9NqEf1gVqU
/ZSqSrpr3xccODxmx8OUzA9d1nlffSfVRvRq8kRHTgypQr5vb27R4jkdYyD4PiYb
eU8GzNsGc9lzajSJFRtSmXDp0wFZmx0rBqWLgnnSxsmENTOhFCmvJPg2PnsUJd2f
GBn1WyspE/1mT8txSr61dzf4NSssG2wvsUuU1twIxrppk1CZf/FG1Ake8jSJu9aA
+nvB0lFacMBlORRw4b3Jqe4qM/iMW6xLuOJ1hu93dArck3LBX1xcOncVEmMK8oSw
LJI185o/MxdyLVaqOPC8m729lNinSQG/KcnZqQUTsTGCptD76TAJtB3591hv/QAq
VJ+Vzg0YLS8jsWP5baF8E4zsHYB8tSNxKU/i8tJP9bB0ji1v8C0un3bUyh/B/PZT
ks8SMEpO+TDn412m4VGbM/DCBu9CC7ZoYZSosIPfsekRkbCd3GqRfb1mWKrjT2QL
4iIRRS2Wr9GPtCEf8Ui/+yyLTpAz45enoq1YtUnXYhu+BM2lA72ljDPhV8YnI7Tm
1kR0TEJVmn5sFkrpAkn4kO0YdVs5fYvW6hZaowcd1Ps4x77a/t+GsIK/LH91jhMg
ZP0qmc+tvyiu3NfecwFIR/tWuGfVnMedNdUdO45b/X+C0s798XYXxpaodBCUM0MB
7FxjwGthYkAKhujVF2L5lHnFOXHYHqvrZcuOyUdxH2rAMl2F2xszu9APuePVIVJY
WNpMz6s1j0XEmqtAqxZjLYo2ug+681Ng+UMLZZGlEIQ98y+/V4o/a0tRiIaVMcoR
0FqOQIkV3JL2cBC4vqCItc14Umyb8o+4KI3TRtp/T+kFIEBLjG6sIbhYqIGGOUxy
RQUinZbVaCWVl6jVrkR21FkdXs61jMWZFY4dM5gAiOKtoXKx5yA7kAG/0ouTAA5G
zOIqsp6izda9Y5kk8LUOP75cjo49WIkmX4IAIu5cZOz36RwNBJXWxloOunk4OmVB
1GLBx8njExmfaxZurooGjDIFsdJS0hDghR9Oxzq9CifgNTXtd4DnxdqXlWgPBPkX
caqKLb0Wd5BcDGBwaHcWfBr0VeVkVCozQ9lJmJvkf85igx6tZkgFuy/batAPTe9T
kRc52vgQ22BcGkdZbe1f/1DDtEUkmUJBKYqOeeUTNXCLJ5BSSLC4dD3B8Eene81H
YZ97zwIRX+enQPqBShgJWRuNfkhsImyFOwnozSZtFJNAOU6At/19Kf2x3rlYI5XW
qQLjxRUjUBnBv1QJY6H9z6ENTS3yxvjwe6S0+PM4TaBOXeRlrM8dh3NrEEJ25p0z
MLuNYPXsIrvIoiS9LyjITZkPo5x6oP/uByAS1rsrPF+JiTLOa6AjA2rV9ktKZdah
j0p+l1b8jBOJXkIHrQ5/Y2R0NpqDt8wVtM2VRpr0zlbo3LP/6CNuoSmQQviij0hh
7uYxn1Tuc4IKpBxIr9QyYgXXlekliioDLwAmEE4CMeKKJY1bhCqLg0uitG4LxUSj
SanQgZISawZTmmqP3N2lmkT6KIBAMPJkwaKb+30m1wSc73gTDY4Rj1IG16DqYIPQ
QlC2w9TJOlYajUdIrlvU6nKvumJhyrogoMlGyp+zHroVC+Gu2qvKBgUEvK9IutNn
w3+p/P7STQFiP+0gloyVUv6DyaAK7TbGsty58IHFYtpHGQeB1wXPMnWX7zCX/zme
UM1E7ValHpEtlBa5oETHq4lNFPOk1FS09UDM9ylhN0eINMIOosr7R+NVn9NVaP3I
82rmLPokCq0Y9f+sVTy5kbYiSUeRlCbnBXj9evmLktBLo9ofN91tCvezhLQeYF4T
oUeqO/QTyDxP01PYxa507vPbc1ZjOHiUsor3L5jRj3mtVZYdeE+lathE3Sz0krsn
6JC57wI7BoJqW80c3zi6KV0TkG9xv3LrlzNf+HRuwTdelYBkOti+U37M8+H5MWfu
Cpg96m4Zkk7pZGwWnY/ly4c/dcGUEFnZqN2EZwwjYJqX/cFp1hO5c1+b/elTWtpp
qhs2ZDmiePvlLphUQ/hla9PuZ5SdIuViH+mm91A8hUQZa8VHmYrcLLLy5/HbEhOD
dYOnmID4L59LLlL9ndpHTRlL+MazRBT4KM4jFyPwpaIJXhXMi1/3Hx7yJYhTdjjZ
9SPdsx8tGOLgGmZ0Jsi2japH7/eQSbU3rtXMLv8LE+NOMnTKYGW5jH2za1LTUi6Y
4MmKzUstVLeuOOl1U4BNR4Gqw1aa/RlmCwnAMIfpsGZfAH9BiyRWrX3sTCX3tYH1
Zi9xL4j3AqnSuophH1d4TtausS00Wa1nrYpwDalAhIh75Uq4vnCjWpsQppHtbl3c
rA4UwSUlFOWizIoKVVOyc1vwDkqtOKNoZMWqpi2nfFV3ES0Rh/2TtjF6/7WiMnoi
e2nrdT/ipGdMuPiCSX6kDkIuDwM4hsrfaTj6H4HABY0vM6pdXnFrDParxmtj8OSS
nI1RFjjSvLt2JJk11Vd+vXeuQ6HELQ4yi71YHOSSATefUB2bYFo/6SnekOcIEwUR
zg7AzbAxmiLSUwSEHp6tYSE1PqYA1+y12uRCrczYowPEzGUWRlVZ4QvpHTtpLzl3
VjCe4W6Ix3HgfPD+r98wgtfj9hBFXCAi8t4fodz5mVRixtsNmENT+IMqM7ppFRHQ
1pERvyMSipCfLyglXyfCpeog3j5Nb7+iJqD9dw4PDCsN5Sm1ibMHRk7odt85oFCK
lkX+P2kR8p83Wa9x/+4+ah2oqB4GogJICskqUYDI/NBU5ROuLr2QOl5yqPf0M3NY
F7GhZty6KhnHd2ofaWbtCn1ppbGGNYbsF18UAOKKL7YSPau0giNqNT2dbfp2sQg7
JY7DyhqRinTJUo2tDrPohrbKSzWo22sNGHHUekXzop2c51idrkyVC2hR1/wpw7LP
sK9aOfL+/3BfuC8tnp+lJxYDp7a3/S+u0tqcsfwCCDfW8SnMJQFZlZmEZsH6rLTF
fM22dunIDnNmUfMqRHXPg0S+YCoaT+L2KBOafW9SEBlAI1/o87EAccjYPmx5IzG0
UQrc2nzrE8NUT80f+N2eDw==
`protect END_PROTECTED
