`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yb24yPh7M45hjw+2b0xyUj3xzCLiCWqZk7+0lc0WBgz1c0YbM4p+XnqIssRzi7XL
flVq21fV/zYHVTzBHUQ/6Rjcg0DuA81eyagvP5m6LtqsOR4p8wfTeMqwdgRD4qeJ
voVPuad5u/19vY8OxT7HN5HyJ+I+1MO6TvfhNhQxuhDTFCYbgeM/6+3iRbNY/R7v
pnR3Kye+SDX2DmtgGNrPii8TSpgCly3C89jr5fKe8HvyZe6U425l6R2W1Gj3/HkE
ajJkLLRlfgIt00rt7IV6shWImZUsWnY+TKSuhFiPh1R0uFeJEhbYag3T50VAOmNq
9CDe8pCCKnKDX23nLdrzX3/2OpSPCymiARjOlJaM4yAkJVT6OcIKXVI+kvBVkNuc
OIhFkNB3dxUF81P9ZXVLqWPlxmv7ZLBIguvc3+2lMFprmekdH8T7EVLhAICzjPC/
lXBfssLD6JpjVZKsZJbRmshD1dmuWvilRE+tWB2fOsHToy5+7YcZFGBFnBSivxB3
9O+zmmMxIU8xxCBt/gdAdQ2ebQogBMK5ZbyyV2ucJcNHcjMvHv1brhR4TEJxNW1t
euyORoEbMxSh7puE6AAV/VFRN03mO34ifXId+avCapYrsA14q492J194tfg283Gl
Zf0NY27G3sxCyOHXeDdryqmMLVBTwAx9b2+7q4j/6+0=
`protect END_PROTECTED
