`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RBlFaONlvuG7Kaz7vIHmjzqWAArrqikCOgIZiK1qW21jMLopCtZq5eL1cDV3MM5T
gewsKxNPtofURvMTQxXeqYD0xQ4LkB/OAvXwer1JPsqiH3EZLrEPUKlZl3J+//cH
qABlluA0ov6C4IJDwAFZf2LOCaukZ9UpC78HcF12hTHF+YkZhTIaEyPWwS1GVFc6
colCjergfSTLJyj2ZJkdPICN4msMQOwLNWxoxLnilt/jNOioZIfekiwbFpwoc1wA
ZP10osdT7UG/VVR0b4M5YcfhOuWYxtJxzqsADYka0/5fWq/wvvCehka/ZqCvfXHv
I02cBv3IxPEmSPb86wuWK200VHDLoFVnTid0sed3H1MYGDX1MHz6lU4eHZXI+5Lo
E60pEgdFmIRetzUceM35w1bQfCPHFDHuqen+8biHl1QQjo1KVQfYRcEZT+J3BD5z
jjaaX0HurUvqmFLn6uqIQWt3+ZhPLJi+eVAJVmNrNpv9nJanfphKavx6eWNoOZuI
4SouOjbb11OJm0DdVJY2s538fiTspafvDl9KrXCY3qjG6SOeeRr/3M+JiC1N4Ge+
CrDxZcQgIBT7+vecrkMCvIX0o4P7zJZoNt7kwPdma4xMbxWGDbwGzyfFvkkuIy/C
p8X4BZq1Kn+b+c3pVgd9bkaTpwQ8rCxCPefmp82uGKtDHNCtnnAN35iycReSfHLs
UNILlFwCsm4dKch6Q7gUHoD4HwGKPBfVUNweyt70D80q2rqk0Hnd6E8d/gmgVABE
UeDnBgOhCYPImC5RrGIZK1j9WecRyNeAMcTaRp4ZaY8I7joteUW/0wA9YEP+Xi9o
KKNCvAxwevVV6xOgXJOOg+dvDV/MZwnzhjOkYAulAte42Io3uuCtAlaEbX9I6a8x
zjIvxMDGL+gHWRTzKZDocjzW0jQiNELXOBD2YTuqZZEAK+QYFtUU/LZfQbzHM1/z
oxkEKIOC9s8A4HurJmxP+tN4s0TJwVFCRa7xZ3UTBFGJ1s70O06vJALKlBJ+vwV2
X6Nn++0awZCfKvxwtEvnEC+9hpQMzns8M7mqr7toL/IQkbdyP5QTLSmJ9ZlLwC+r
lIRt31CQJVrWSVLSLAJu0AUvUOcrHNnarAFS1k6cScYuQnM+wKdgCU+3F62mRb66
jAAGKgy+WdORg8t00ZavVyuhsA3UVsrnVpJsPxr0yR/kk+VwFIrM+14HNlSoriCk
xdtXLRhBdnrFAIk5KLF9JfAwTkVyXWYpBrG1in2YoHcJaBsEYWbGTRkymKL0av8D
Xa2/yvXA93T1UnOt9f9OEX+ZDIPaZ0QNFKcYybEtAiEf0aSQMIVduhfPMHcDImkh
SgB4bBg3NnOT/Ms0mVlEuP89cnXQ56cSKwZpTpVBl/kwNkfL5/BtOWgjp1O/Z5pY
FsjgcxcH7nlUPYCLruW76j6hd2Qasp3v0DyUWX88je1SnFtb/pQMQY5MBn4Fix2T
gPwDqW2pZq92upsbo/WwsK/TeKuptABb3kF7FU/6fo3LpwfUaoHXiCLzED85jmbv
1xtYwtf3/o2jP9J5H6v+Qx/LH1xeI6EfA5Wc3fLQBXgmmIEZz8xLs8U58P9E35ib
3ZnomsICNUbV1dZ73hjuLe+gnu1gwWIqz8iohCNZb12WiNz4WochW9s0BT/ofmft
5wXb4r4Unknhs8DP6VXUk/xtyot0ruyuxYRhh5BmP+6zvqkeyK5InOVU2mnZLf4D
J9sbyRuJFO92HW+9/hqCO/ucobF/2sv/uEn1EmHlzBqk+MI2TLyHP4kTWYoq0oLF
`protect END_PROTECTED
