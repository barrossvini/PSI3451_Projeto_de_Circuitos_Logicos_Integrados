`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DdRB1JC9xaH0PHtdAmsiTTpdbxAjhBdloHb1IxbmVk7VdAnqqtSBZXHc+oHl4Ut6
kVUvQRVE+5lT5A/005dWA7rHlqbI7w1rC5F19tWcD44uIq1GwSVVjmFxfRR3B9Tw
TZ40hE0ItQJU3SbDRX1v8RXqy/uRaXQTz+iOBsWUs0+VUy/224NnpawgY+PMq5xd
UVCK0XB+V7YQFUsDRuZM6+GYVd9JVtZYUcERmrmMFVsIeB5J8VSNeHb3QlV2A3TS
re7+c5Cs3gJIYc13ShqBGHd252gkBy+FQxwhE1YJAOBG+UsXidAHbGaLyLLr0VyM
I3zRikyykXCMLOnO5ZOTqZnlw5ZiS5fa1sqvQ7mgPQjq6y8e5hhqfiDiQ1FiW3sK
+vS1fxlWpKPWO/cRkJpYs270g5iJzte9e3k0Py29v5U3FDP8uISGtrhL53RKk/fi
U87ImI6EJ1Ax/e5uhy45V+5zK7wfA/FTop81Z0wk2/RHXv06aKKXV+IiARiS0Gl9
mutvbt/r2HhwANqc0Fc0QfhtQHZS04+UmVq4Ob4MTjsDfu4mJbOMoa/01CrLenWf
oeMEojkzWRqBfiHG4630pEIbzOog+v+GRL4RXSb6tZKSZnNhIn4VwxIN3CqI1pab
2HJaHYZy555iCBGSDWw3WgipisIo+9CzwUX+5LKt1ZRGd0eqZjza/DTvUuJIRxdD
Fjn9PW7R0XdlrlvGOTboUT1005lQcFbVn0+kMlS/lhO7ullNCO5QelHpR9Hvg327
eof9SJtw7BrKX+Zk6kdIC1R7gE5QDfBkxOXNXcs0tEuGJxvWM6CUU8e272RxF4mp
1Vk73+W0H669V2qedd42ymMCe4A0tRql7S548ml7yjEws2p5g+omWrsiWnzSv/US
hVKQL/CzChGXEaIn94WueGbQgL/fL1pLSJpR/oblPlw8LnWneRjODeySAZozOYV6
IcR1LIlS66uPiFXGDao8pyq0pZColSEvshZeHtbH6iK0fKWpYeix/oCtRQt6sCG+
Xc2QVnODJVdK8/Yykg6rugvwTRAVzC8vqaB7iut3oL8+Gh8kfq88jBH3nxS50+B/
EGlL6fabLzbofAFhTVgXn3rOyYNwztxO08GMTOBYGuypYc06WPR8SfC4JDC7HC3L
uwPQq3ULQO7pPVM/+wqMkvp+t1CG0jHmLdNpAiuagL0vJADy4iU+n2lXK5KLBL69
FjJtEkwmnRhL1WBveLIzNA3qRanp50/2YXWD0Z09+M+n9cV8efPNIc4y8l/5Vi5a
PXnxmm+usAiOR+3FC6nyM/ysAr/ZFUpU67gIxK20cga9LPHXgf1Vmv6NOkZ43Khc
RBrXu95oKmWG9Eh5JZh14C7TETIj96h/piDtO3YBaxYdT4HGzy777+VwSkz3JBmq
Qfp63JCcMZNHjFgwcaOCh24bGUDf7wQvP7Cc+eM6gzpTM8cF6kynFKYMh3b83grK
0K0MIvcKRalv3Ssdz9nQtBD1n11S9lkd//wKnWiG9RtFnbWnL1QRC2FhDnEPVZko
okKyg0zVX+Jshszk25eI3LVkI8KkavPts+9PJKJF1PsVwFjWCCp3EawfTQsZDE2r
OhZV5h2EnjaRRax7BkH60qQ6Zav65g2Sb0gGKv7r79pRKGwEJtlokjL6YKw4ce4r
s9rqLvAITsCPvgDKGuRxj7oH4a6dVpmXDVd/9oUInlnFgwk9ppd8Y22VR1moqpYN
HvkC2X3bvP5haYhsZiPVbCdG95i7+35TKwGFO/4z8hedkClzLevut+u+Fu4kab3I
O+AZN97f1Fnc2pOwvQc/wC34q9grOMtZv+Dg3N6+Td6nGokxyvtUVWQQ+COzaWhr
fWgtXmfXe0KT3BvHnequCCZYq5fpXYswxY5uf64y2SIHKxTLft7/+Le4EJKTiYwb
yd/hDHNDIuUQF8TlQXCulWiKuzpPLjztXT4LOZa4CkaDxa5b2I6gzE3/x+jTO+Cs
naWAWzhw2/JbEIITpB6srO6Y2Jb11SVb98a0oQvvCFQewKjMGEDU7N9vjPlnBjcu
Q3UFd3lr3CPFH80JJkFX9gkJhZzhu2eOiR9t+iP+biuYBTEDsBJLPvkzaJTxeynq
V1C2G2LbLrds4FXxQG+wa7QFGs6i1ykWJYK7vtmhfTRelNMb+5fZ0j5bKQZ2bjLU
jfPU6NfnZ91W7eN6GJug2XJLXFCF+9E01CqqUwYrWyFScFVqn3HGZQXMBWlq0Pkt
ebBQx/hHHJuQ+meGsVLdIpOUShWCaJmJPupE0KizAWijWgrMKVHKbxNltAtZrT2j
FYL1tT19RdW/n1VYBOPZZHjUQQy+24dPmVAKI00bXk8zFpKamoQiafNoJF2kxASw
DP+eSq2W26pYlnvMT1FgPrvPWQ1T/nuqhTTwuJBb4+s0QVJxVmdnDJ9SCUYMvXol
4EiUwfWyuoWBB21k6CX7nBUg13Bs2KSJykdg1YN7slEJe+/hNYXodMmVMMuLIpTc
SfmRqyT/LL+VHJ5MGkTSg8GxIc8Ea99O2PtISdtuvEisWSuvp9Mz5OaYPIFO7aQO
EvSd6vzWD+4f+yVCwsfdePywewx1pMmqaiuVM1WkRmBBPYBbHdXA04FUoIPU2Fb5
Kw1e7AuMf3tbUmQN+f+Fg/h0hBIxMEwk5vy5H8DzbuH9vJE7c1K6gQ9bnxq5mzCi
Ea6kc3peK4gag9nx3X6n7R23XRq4wKUNa2mIlzfVtQFRH7sDbV7h5sAN0mDJdYd9
jcxQd5ISXjuPprQPecK4lp33ZW6GP7/0B0ha98h5PAEMpl+nqcxAChOZbuiz9pZr
a6Q1HS6QKNhEcKPiFS+Pizwu7+OAX7qR8M8JDRBBaTWpzZTTbTe8NbEdWf+t3Itk
8WyqFTfMa7N3Zp2EDGfiKl7TTmLnXpbiP8Du6w/VmS/MrdiuJZc7XdDy2M4w0Ssx
HqXYnkVqmBbs62k3tMYDLc7cKa2DgKHX3k40oodBDCHLxLw1TiaaF09PEEE9TBHd
4TfVkSm8lSexTiE2NreiRkRSKc6D8qpx4fRhK2ZpvJplS7d4Cop3bNbK1eN02XgN
o31UfL+Xb4Y8E/e0wTFWqlX2jZs5y30B03yXBqDwgoTU04oeKXmkS4cwaDV64Xul
9H4Uzx39060U/lVt/VBIDiI+aB44U55q5l6H36xafp2FEGKjmzujSFIw+GMHZZFP
M3Axi1d4Pszxe/3191CWBPpbGJeom6MHNW+MCWTNTA8AqK3mBnD4tflq4SNQwWMT
EVAuT4ZiHhbUnp5zBqL3EjeBI6y+C7fnZNOisAAZ48XTFay3QWGSTY4Z/nghj8ZF
yIqcXPd+NUfge78SxlrLKduoB6Yxb0ivbm2kNLXG14imY+T2f3sg0XT7unn6wSho
FXAgt57kCLNcBkZ20VsFsJLI8dcT7c7HQHf7EzzyNJK73aDyZTlfarM6SLulJL7a
fqe9yzXLZT/oB4UiJ7I4MKHUUzZOxD+CqPCkd8FtgBOUy0hbWfoFIbmy1I9PtHiB
h2niS/DImpqRVUyOWWrc1RVfqY4aqHmstlhpALJT8qa4ADjrwlBHllEkBuFCxSjn
fXKwyje6X3bIC6q3IxAb1LQ3SGn7WJoag/LG2biBxc5YHlM9DmHp7fshC3OLAErS
rCFlbfgphlDyHuJu06RV1zkDRQECJoA7IqlqV+58E1Me7dW4AW89WTv0AxwWYJev
z1kLwNq1TG0rQWTwU6T+lXawHSABKAVO1WzRKgzU1VP5Y0tk08kMkIYX7Rx5w6y4
Yy4clH5/DdNzFx7jjJESqY0BkVTWLNaJaHanfWfKMWqS8SQR3Vso/q8ulLDAfp99
FnZ0pqfpbBIcLbW/3wU3BOSpi82M9jXwT9LrLHhXuJbnVovXMtBcvDeCz07/Qyhy
MjuX9s9wiLng8u6aXPc3JyiCJNhH9TXlWFKVXbB/cl/66jfD0nTMfxIrd/DzCh7I
SUhQF0Wg1O8Gm5BQhLZeBbwCcyNtg2uTA0KQ4JS/XHCgcndW9sbO5Ck/nvayU0ry
nSZi+5GLSiwPEhOp57VAgMzwRRECWGtq+vqzjqk44gvLZTBdaBR+2uiuY/oz7QqV
7BAb3BNgQ9z/0ETPQOVnVzaVPft9jprelHSHzjuPSv8pgIacfwDN1K1Au1c0rLxM
3Z8t7guBl7kEiGVCk04LkTLfzJqs4Y9Hboub258n31ddLFWr3gP26+BjSCffPRPM
B/rrWN1JJ/RKGXrWvDwnhixghUEzFjJD2D01i7oUwvNkRw6wlSvu/dAlZqwNaEik
9ilywNyPLSTO3fT6RgzmDaYxYGmfwOPEI4sNeTRBFHqrGPQFplwYrFjmr2VMek3y
87vexmMUpY4YzmOpeoQ2apf/135I5LA20EPFAVncG9br1oqdEeM6msstUezKef6T
pEx1/MolU0/4Co8sQDJUwNgTPSVLpCdb5JCn/l0xJB8hCv7Opow5oZOfhoE6wwrS
Pe5emR4Nfum5AtEDDUh/DEjl2hxTgH8XFEQsDIP831b67X2bTLXakRLrsR9DkUEN
H25ulkQG4n+S0mkGBNPXHuNnE/Wy3kH01R0OfckBm5dFi2ERpMRf47CeJeRaUOd0
+Jutga+k9F6bsTzhOwQpD1gqnqYhwabzpfYDJc5NEvuriwY3tupNkfI4uaaRf4YI
OxZKoQV7Q5QIiM3goZvDGiKUt8hIUDD75ue0UctrxWIshocDoohJwoMqEL/Oznyv
Bz5r/QtW16JltW3s0hXqRojZLLwgVgV+2yBurcA2XTVs8UFdkmojoPNd63h0307V
Dyfb62x1ZBn1nRR2L/+Ul+uyTV7IOoHtPWPqOYXqqzV0ke7nG3fX4Z5mAQzpcFu2
ZSUTr33V42AefiNkXMtu6/9w6wg+rUqQqv6yJp/4H6ba7LqXdz/CvQCh/j8YWyKG
b/gOHacoWV/nQxxLOzOzfJFgYQyg8u4i8Kf0BQF8oSVBmkmuwrPkMri/nsk2+gFU
mS5aTwuAEfZ7bZ5NrJn8mOSSOuZc1hf7Mx89WsHGyTelyeRSIHzxKQtyLse7DJzS
vn7zoNstr6t6BUMv7yv+94FyHrLZoJ/P3zvPj9KlN8qittAbunA6IPCKVWqADOOe
d0VwTDvUBLU811CG9DJtMrQIDTTOil7f/62QydgZyzAvTf9KNEcFOVOVhJSIJ37k
72BNWr2IlpSDN/vjJM+sbmxz3IWPAVgR/nIsSZql/ZnHrk1+pzYDo36FupRy0ppg
ixWAXV+IDJd/305tukyzpUIsG5qzb39M/BYYSiQUglykZwMWITg0YIollSE4gWJ/
xUUOYvgvuIK/J+X+pTbe733yMsdSZBpQjJ66AJTZN37Qh9Ga7VjyRyNwstzroNjI
z4PAOn2Bi2xJUNlxFO3OHY4QVg1oSdp5JVC8YAc4GNJJqXt/lTmHaYPo1TO1uFs3
CMaSHCiSi0uNSeL4p4f/zsvf7aKQQr7CuBszagUdB70cEX3/qnIxrHDBxXjg9IkV
8S4UuXn2pqzGIDejgxxz6s9pe8rTxfQe9JZR2o8o9iNx+TQt61HvIehhNN1csIXO
goPLiSFq9WyDhai6mW9EPkZwRbrZ3mPtfLR00O7HOOvPJfqzDaUcxJT8N/1YjflE
fHN1sgx/+KSY5wzapG3fcCY8swFAhd6P3Lq1es1GYoquXs+ZspF2HCBhsmHqWUpr
fRM5IAOKRpO/gD4xRG+vy8OpRX2IaR0v1drF0hDr/l+fQIWOi2uPXmKWYMbk+P0b
KVRMYLyUqT7y2cmcSAdfxmzei/EnRnU1lLpBoHSbkm5daBCPfUWHgKgHqOuodRYD
Z0DIrN2WCOXDCa9f/ZhyZJCX0mgXoxuiy84yvlVl4AMWbKgeNfGf3S2k6IYJGTu1
M7kbdX6st6eOJ7B0wn59jsDN7J0lNV53XzIXpNhMbA58QMipSHQma1oaT15Upd/R
6G65l6AgIt1sbB7hEFKGWEx2bXuy8FEmIco+D7//qcElr4kEbbHqbdmxWPMMosEl
5qefyjyx2f8o2v/UYnBVbqaL3BfPt9dxbSRED7hHUF8L5k9bXASWk1JDDSlmoeax
4oyD6oartPadTXgOuriO8i6yyLVDzBAzmXha0qxzhEJU/NbZzm/8MUaqN48VLDf+
vOhFmfkA1y2vgHdOWKp1Ao0NPxozIFPziPbhZDMoXv+zXyJG7UiOhbdSm3yGyoD1
2kLSmKC4u4KcvEzF4BIISFtwPNt5SF6CMonQEFCweblH5ufC5p9JcvUCvlbiDWsZ
FF9g3xj/rCgZHnmu5coH8oEtCTNDKFaT2FkYe9txkVrG9k6s0rADbBsb16bEGenL
XfLEvUI1Q4gVVl6dMapQXqKbPyCTD2jM8IvICMAWAi8Y1F8LyYKNsXNcVunxnJ94
DfuqHPh1wtOE/6maFxWci7PaU5qenH84IG4Bvr4ZjN3vJRarj+2kRuwgFLWvj+il
AY7LL2D9WKiU2g0j7gq8pBEt+m1myQHpvnDf7c2vww3WqtET78GvbYaRSXvgq7f5
aZxB0UuPFYSUPo+uO1G4bsBeMIdSJyXwZnBSR9SYr04EcyKHkQ2V+Q7438/7y0r1
lw/CbEQ7/+V3MhB+BHxQGEpgV1j6rRgw7iF7D0wWKLNED74tZibWBjB829CDQIsM
Kih3R3weYMyZp4cC1X0g3gW47RWMXuLCcfobi55vHvPEwv0FEKS816VIbKhrsKMr
O2NMB1G7bIZQMqqFGTvkPRXeHJ9qqaJ0G1w5rpPQhLUw1ojZ53WfcTGgBIyRnu8d
L0uEvffiWISXvQlHtru/ox/0HgVYwx3iYvJqVO0XkSrHmFl6Y0/8dLM4gYj4qUeR
AiiP1U4E0M/HmkDYvAxFrHzwSTCDgw7y9r7gkGhlKFC7OfPseK8lPi2bzsLAyLJc
6vvnvOuaCXhVahwCyEB26L+wScO32gzscuaPQSNnSMUH1p9uj3BWosD+ZGV2/Hy5
Arz9al3MCzkzP8eB/1hWId54FbcTGb6yXJ91LwHkTObKy5k6jEsh8dKUERCUE+Z5
+cTCnNg8JPHirpi6OHlPJzfhzoaQ8YKrBR3odloRJtEr6VHkaN66JP0+acd4NtCp
RKYTxo4ed0n5JYNACFpNLhJwUFxW4dlcJ6Op2DKCLsZdY9wtXROUHpuWLTZKKdGx
X7ciI+0xsUaQ2GyA7IxdpaAvw7pHmUz8UpGGTMK6GAFRwe15NR9fAirEQpcnmTqG
/vQ8zWJ8DBv9NrDOWt62AFXx/SEg9toejFCvwl55/+NeqThAtLAhNxuMDPhuKdLh
v/cU4D4iqboZ4zXW8bLyZA4yYmcQ7pTY6jZkmdWtnKactj6cYAISF74R+Cr0RLUe
Gw5+q65Y2RCvTRK12DIdCSBKj1JUS63XfsjqtEpCZsrcSq2vAk89whICCOZuDsfP
z72FVq1Isvp683jgYFswW4Wb3onGzTB803BBW09/DrTj4XQZtoywlbGT54Z+XFFe
tKXdpLXPbxoowj2KT032HOC6RK/2cb0UVroBdIC9NE8bZwdNPo+4bjI70MQ50vtZ
C5q83jE1d1hR15TQVbxvvePHI1pZrbJrQ+wsGr6W34h/xKB41vLBcpxW0tVvH8U7
3nge+nrUKWYm55Yjrs2xGAyG04L0id3ZPHoiZSHFqRSHcwgwjR8TclB9OAbJz9W1
Nx6kkRMSFbGl7foUmaVOjvklJIZCky+yQv3QwVbkT2AXfJkKKSvmesAoi1nGBPcQ
F7PY7wAPEhfWHhsKjlAaMcyRb1AAeleaZ8I2R9C/6puXYDzr/or0J49WQdiGgU6k
BIMZxMdgWaMiUjtN3x/IlbspFpVPIGVPZovTLWGgmxBY9UVI71afwmJq4Kv1UE4N
s9kv/jkIirmVvxJVbJSAxyZaO8WsP8jlAMvnNfK4DMH5X0ckNdTFfBJpCKUZfYh2
q4AsWKmiFB88JP1lFPxDiEPbWiXHwoLo/9XO0mcmBFU6Z4Mp6ffnFIV60ZMWFwQv
DqaGQ6kBs03daXRPI3XhKY2kvf2N/7lf4FIgrRdhq1ZJ08yq+phK9Es5bndIWwqp
3NkT//vCBhlxf+6jS7vftx088CWlOUJxRH9rmB6f2b5/OR7bXWCeqkjSO5nFNRE2
lqGMB4NKfgaiEPPiGAhYjm1ANgCwSWiYmKtmrmy6tDp2bCXkcqwlDjphN5AOURhx
gG2iizdHWwLORjHbZ4otvL+MmgprDsg0VOzDnOfIWvoN27JkN9hbpC7OIKOpuvFg
nnjWe4r6kwqQIOcHiRuuIBZCgulxxUWRYtkDZG1n6ha/6MdzmMt2FOoztl48fbjn
bCYEdz1k5i/7lvVr9qltjY/7V1SL+KW0UheFFH3Euk+FKd0HKOvPLM9Wxurp0azH
ZpqnTcgWEfQ0O2P7T8MUZOI7vPery3VE/ryMHJCAI77RKV5qTFkHS0Jni6Ojswg6
3xVED5+IJ7GizESEnr8XWC2JWn/NJBK7C20mYWSJbZod5LtLqUjARQ2fG2vZWIdK
Qf7PVcLBwGHem8thfVOYGXrPRDn11JwoH21M7QNgQGgxqpzHe/Jo/9/96bJ5mXvW
bIbK+Bbh6MMD8LhBC5XDAT0L87p5t++FsysW0wLppqL4KVH5mZOhObYprdHvtE3V
jZAGwlOgK1HeDK8+bhYflXEu0vaky0HQwq9F3ui7x0jsFkK4udjMtMj6QM896VdQ
MWlbH/QnoF7pXN9KQpNeGgKbbdOCBvPeUocmCm+4kps8+GXDqV1dEQ86v/b+wWMO
chCcy9bhs5qkTIfXGNZdTQ5jugiOhA+m0/Mt/P4fREmGuyalpScZLEZlLFQBuAyg
55H7yPf4b/Hoh3sw9tnbrn5+ZXVy6Ls/C0DwNm2117otxyJtgaWIogkOV6xk9uxk
WNNXZXxnfgIABaQPO6yWEAvi7UYw1thKcagQlCpd+jtD6t3lHg9Ydnj6gEG82Ntz
yhUZUcQpu+FeNXh84aYeZ2dNcYahR08ofjk9yvdYq6QFQA7NFUFeQ3HlrdVJSYrj
+iB+dM7K/lDSejBlxt8HszY1Bt0s1UGtkeq3gNmE3/1s5oErAHjDV666E4B16cHt
+mQJMPjnB4KIRdd6CE7v5tQrrqPad3ugZj+xifYXygc1xREadAIoD7ErX0PRz9P9
DP6cl21jZlhoV5VUNXdKas52AnEMSE36ViCMiR/oQ7p1Blchf3yOre2r12D5M1Il
1fHOUyk3+i3itzHwyknLgLjcBgzdq02haoNI3UzfyKZiauoWhUQ2rknWEsCqbTyt
SwL3hBsayPTPa/j4cWzonRx6vdrUr38BTnR+IiudnTBgaNM7L7mj2hBthJ+O9eD7
+aejwdwfwF+feuP2o9/LpBsb8q5+8rkm1NJkATVVfAMYhdVUDa+l8iHwus0MzRzb
RI1nY++r1bTGsp/YxGt0MjqL1X5RNbdcoPQL8y1U7USxoVJhyqRCtAdZFUXW//e3
HVZhOCJx/adJm8lF46LDdWRYllA7LccON8EdvRjnvPqCUpF0SOCHycyd8nihfuXR
djyE2CYihC0DzQ0rzM8bUC6dftlTtMboCUQ4169sHL+iiU27OjuNnPadaSkNf6wS
oQIzPv6HNSFn056yLGavuZzwDnt573DyYUtvFzurRxOWO4D60Hpox6mt27kPNAbF
G86rK8YaGk36dLd3yWN6F2rbFZAdYPk3Dz8UEq9yD7ba5DsCG6z13T9RcQ0p5AtM
6UyxMN5B/2emwlsp5deKiqmKcIknya3MoCt5Bq6cuN6aRYQ0oRTukLer6wQnWq7a
rwFlha+t1FXwb64AYQ1ThOH8j80B/AOpOPzXx2k/WQ2+/+4qon2s261Ca/ytN9fT
+NePqZ7P7sCaA3E4oIGIvPPUCS3D8H3pE1wVVx0jFnstbblqtjF6s+C62clwfcij
kn6kO70g2ZMI+08txNPJVLS7Or6W/RmqG9QlrzlBshilbUgh/aXM/hPYP1+I12/k
8SnjjwGZEain3TbPnElFT3dc2Xd10c+a+dsBOhGv8OvzUtW78LsVD96N0DeQ/Amh
4UBxsA9KmRdk4M9xrureRA12PtkAIZeHCRFGOTyfW7Do6aBnbzcIZAR4GjrEzpp/
zbpIO7xLPB55W0C7J9mhU5AR7e7EgUtYZYlT6JPrjT9pbNVqHWHDnsYYLY0gP2Uo
k53jmJVBviMCBgWu4ooUZGwcbVpTSy2bswLJ4DAsF57yD13Quv/3p+cyn8OX7Gpg
QFq+YlgZq6pOVPrW2PE7O81u9D9CY38iukrrWtcdVvzbYEHiGgJ45qyqFdPudIbi
6bVwUIYjJ+QnwKVqylc4EEou1FwfNMMSAYkMmDbz0EppOjfJFdRjrmOZYxwONqZ3
GExIgOxtprR+V8ZV1MaMXfeK/L+q2S35C3FosIAcYvHPzNFm663I2foaKgNyLCP3
WtZ72+NTKbK6qQWfq3R1RUtcAR14jQ0DIJjeSENlEAF7wO/BVj1wdefImA2hfkeb
9U90dvkGxl9QsZUo37wpk35vy9aIfSCGP9ZYx31UubnHirSrCG+pBlkzeg1334A5
Cvqlmr+b2PCsjJ5eYbc4ysaG/j5wU6MRKXQ6JiUNPG9nOWYARBIn/DXhrT5ceTtk
a6wZWHf0VDfPeD4ZGAr6iy/vbBurJlneFCbo1HazEI9dnFjp4zgLAWqLpN91PdAg
wduRa+p2pEba4bcF1u4fw/vSkzCfDocd/tedwpNBe3WjePjiXe0J9/J6MqMJUEaX
Kg9zwEXqagKwVGG2bdRhkduOAAoQUoyjIby0ao+KADiuC8UYMaUre8J1yG+mi0MM
aY0YkNu816Ce00K6vTU5X1Mm+PYDK3PFSrf+M8Yy574=
`protect END_PROTECTED
