`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Ou2uXxdCEYFQMUy+pBD84zK64oGihLR4Hxszqad/pIAuIP9uA1Y3NwhdcTOorrb
1/OmbGqoNQmnvSU79XnmpDtaKrE6Lft0kM8YhbNo3EXkyXctGbq165nl32MxFGzr
UaP/QRy+LPwTFziyhjYaPSuEhu4nGdKkuLZF9+QvuYLZr6Pf9i6vIn5Sk6MT1o9V
JNSPce1+zAUd9ddFxixskMs1WgQIxxwJLyhNLD/JC0DTA4G+bty9swg2U3RiuqQt
TYnHqckyj359+i5PlcY5s9SqJJg8M2d0gv48TH3islz8VkOMnb1hXhhNokA+CUyK
N+QzFGoByK7J/9nfhZgx7RobypTxAJ/eGJui/A5SXhsMJ2JC/PaynwHMF/86KG0j
qpSlTCDD7VusVR9lQgojHoaYLuKnx7gDy3jO61sxIJwOLmUamJKIMLJNRbbSzN4s
C3l+36hCsgh/0IFl/nT3zD9TPqRuM97KBjQ/oYtvwyZ4kJtrWhzQ9iQbpCZunKAd
KAZQAcaDXsa9B+tLmbOmapjtj8O4hcDPPuBesIUbo+q5AsYM6AuptnU2zQt8hUXV
Tp4YLEkTiRVxdxMEy4H0Eh7KpZPOywBlV1O8XIugVhd2D+vRuD5sOp/230VtSoXf
skIDYt6FjxwaU4CBzZ/jp/UH5qSa41BiN0e4p7j4HPb8KR0WLUiVwE9VZNMw5Ss4
iFYovhTM1GWnTdqA8NmSoJubaGQbk/7Uua4OOz0bYpo=
`protect END_PROTECTED
