`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
loBJq5qSZCWAtM283lvg6OArH407ohMD5mmnRMs8q+J/HUfnq/V+rKmdwiBggxqW
kcIEP/VEU+PAlU+OxlgS/YFjeR9m9jvnb4I/BWe5aH2FNjSQsJigR1N6k6vcQw2H
+HX7Bx6dITrE2RwmkxjE25qIQm+TilqmK3InLt0eJg1NTGfVL4ozIi2BRMGMgTNw
QWrn8gJzF53wIB236IYSsAsz/kSExUCk8t/eiNY9DnhX5B+FZBFx0P3ime+JjFTw
Xfjxdt+gGq0d1wU5R7Ug1MCskyJ0VmpKAm0bKXHtgrWr+CGdKunPwkUaM+U5CiWS
hmcqXb/bywDsBR+ZLYt2lx5wcrx05iobEwevtUCuURSmLehms+i4NR9h1u3IWQMJ
PjSTwWxhXeXT0Mq5L4T0BsGoJykyRwhWPwWoiGVgEfCWpiKzPsDpcHDwwzIwGwO0
hoCDDu3ptEeReKnJyGudefWWW0s2pESngAnBYqrDFA/H7iOKNePeEbC+PBPa5TR/
iC1jXNNIh1ZtPBBbxn/wp5lJ1an4UBAA6tj74SSWBqoR5HL294C9yPC9CW++xasl
LklMPyKXoQOH6NaaODZdESiVwo1K/F+dJfaz99ljZ6e0R7Qj6ygd2wAkOAWvDe5j
aDtD8IYNnlgIU6q7qUygsB01qUZhLP8sUmY+BrtVoSOKGj386kt5YLHBlPeOwCTz
smyUI+20IS8ckbP92HPHg3AmaAVZdySdmc2yF4xQyxOWNsmHc0ieJrQq8nolG+cs
JdNTqRV1dmwUDm4BvNvDk3OzrNgiiXiv3Kngpuj/T65nPCbMmUW9zz+nHUcFj4pM
Lg/02ysIQ3k6NW/gHuGknm2EzBxHF7kmbJp4NZyKsr/r82nyDy/NZMTpXkAaX1oH
wQHFaWccJpneS4dQfpIpASBTOiDqsUDKZOnjpHlByBi1YFfq5AHf/O5kFAjwV3Cm
GsCUzKeibVgQqj1s86/2yQ7I6jB2rx5UGoB1TPEcaqCIoiKbMRFMUVtS6N7w5vVU
X0WwiPV853rWpTkzEAr7pjtGV3xR6z/IQq9obUEmmPx2RmN+Ln54lTqc5UP99jJP
N7TaN9hN2blnivWrPtWwi0CNhPoIt5bGRg1oimIHLjbk+rpbs6RVlrJkghUCqXXD
MtbGclzTr1LQKMZJXjMuC0zUqnmlT8EUbse9FG4AzSIjpgZZAk8nrb1N6+tfMBUo
xPVwAvH/BMixFQHcYpWYsw==
`protect END_PROTECTED
