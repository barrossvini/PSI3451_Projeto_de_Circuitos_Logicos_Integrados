`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VkPVrdBI9V0Mxy7yajBDikn1DlIH2pFcZG0uSvzXu4W0MF6LkE1zLFAriwpZu+Ki
QUNQeCaycurC8Mc5JPfukjGlHASLwqsXd/cjLIAYdKQuy7+0qcTjC7OX4TUnMN7j
LTkVydIeQ5hHOi+SDQqa4Vyy8asbLh7cQT5i4zkiy2tx9+iJFh8Tr8DwTa5+vTJZ
e4jVK9bPJiX0uYbw9MpucSiHiap5Jjk3dZqLAGvaWpkvQaola94CahQs95vu2rMe
tQY/v697156+bKDyFykrtYfOkIzoXwJyS4GMTLbBj2h3za1FU8jmz1atxQlNwmON
0aom6tZo/QXRgdC+4PIh/3JoxADcUcLHoKKwWJwnsKeDb7BfRgefAz6bAkZTBOnF
ODLzHXgFlfIk+rjPcPG0WJrfJag5olRsmGGXmVBlU/bHpS9K4bVg9PeUU7cRvVJn
N2bjfgZwUFQzYAFFymDg/g==
`protect END_PROTECTED
