`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2X7mLlknacGZ4eWlbVx/oiSe3XAC7CB2M+otWDCB6H8HVgeOaji/R5nhckTzonhT
9XSDOlUTzGKUH5j3J+vSlK3haXkV66bfEg9w/IOuLk3IS67a1EucT81j4HhTtkzn
rf3u6mZOFh8vfpLDKzYQugrts5hkPYlJYBTpF0+AMXKChGaP6R6x/0uaMXhk1g7r
R/GbqPULjitEMmqKoDRm4tnsKKSRlb/30jddSfIlvFT5CIDl5wl7YgfaaeXClFKU
sOmX3L+QgQ82gvK8Grh2QGfULm0HdMhGPwjNk/Xbga4IrZc3oj+uU1HzX0nfToWB
0RRZt4oorRWXgWwNfDtdl4tLTi40W+JWBTqCyK6r5BaacKTvStauJWquOsifauIP
u9cyUWE09v2YyColY2Pp3Ak5JvLwS5QOVNG16QQpcZVVMwFYOY8/gQaDAFdRNFe9
/UyF5T3kqJvYcePjWj4zVdrVMAXZotyurqCcdpaeYD0r5x4u5YzOvfuPgwvVWhfc
sDQL3KA4XTcVA7ULWIBycZ9wyzaEYW50SLqm0/jZ1UGcXPe4yVQHVmQCOBkvSKb8
00DMlBOE9DHBGLLv48+dBABbZdvlnNkSKEmLH5tFki/9s3E8cbcX6iEzxiDmeDT8
4V//uPHnHqsn5bUqV3FvnkLhZGoGEGHj9Xcf8YmDjV+I53nUCtZlYywMgH3IxijJ
fdLPKpU6ZBFQRzvu7HKWzqPkV5LIsIU5eao4KK4O+DovDzunXt2XMhvKdacLZLlL
bv2JdeWqhhFvhY7V9UepTBncZcUBStpM7FPfQBMMsYa/naUllGBtDBdsY9kP9O7k
YXOeIDntrLRT8hMMG4w2czL5syCzSALn/JFB5Qag/+9hFut3FhZwUSDE6GntqVec
+mmUzSs3sdHyCiqHQ23IBywxir7vRZ6VUD0v4CMmLG+BTcmM8LCoUkkDPXw4bnUU
zsA7BXtD7zk/00gW2YkGfFut5N8KbqLkOFxQbEn0JlKm7GVsvu9pQQk6c1Gc5vQH
jl8s3kHA3LGHRwvdEDLVEnY/Lh5T6pPG0SY0YAYmwo/Rf7FJDZBxtPomRLk0etIc
OKNs0fCvvSa1vMUg6VqtmXrjRbE+31W2QBnpb7lljCz8jPSlr+Q0qd07fhtfwsDe
BLv2h/MQM5MwdQKDL61Ac/go27k4PgNAN6dJ1XFYHFTkbGhLBpcvt0mNSDkJAxV4
CfVL7YAR2nvjzuUxvVPQSRcYYtTBYrA0jHYa42TtaIdVBDlqKuldYvKag4sJ67NB
cuKgXH0CD7KCQ/lUMoydwCy+LN66vYazC6M9wBiRTQHIKiyRZ5Y+fX4ogXYS+i4y
87rPr5oAx9Ud0rElHQzDBNoP16cKNANsTCVn8J3n0u9ZBsTRDOiEuBRjPrPr4WLJ
d2/pZ0nOqs/pJZLb1shVlOSGj/CBUmiX/5jYPfB4rJX41ccNSz7hcG0+g4qHvujc
tE8ZnP3dROGZvknSeBSMQcx/5lzKZcGjXvAc2PablelwXrcGryM5WusVQOVQpiH1
8D8cP7QBAi0zsipRR2M7lPPX0/v5iSA74xdT7xmpl7kWoVS4v72MjTdHik//5NA6
eMehztgMBSMcEqHWxGjdEPIqUbjA45rLG+EcXVPcdMNVhB30qoTyb67XmJLz20wJ
nYwdgXjBPtAwsuR18izbkPbVyRH/imeLYcs729m53AmjXqPsmUtUSNY/PqDEFdSL
+cPWCdOc1hadjBJNriNfTmm5tRNTOd76u+qTiomjZlAjZLptjoO6BEa/I0zLhm1V
ozIkfYvAQ3BAbKIaLrY6+eDPxcYLK21R9bWKFjdFsMplDgz1W1OvfxwUDKX0t3te
P3zSVIKxeVOtsUljVu1lFPz7Jjj92Pc9eXEREU4aAiE4aHl6QsiqHCh4lFjfH55K
/wzofzzSogVqVuJWTvDT10wKbydplvPbWom0ceZ/nyJR6EBrRYZxdv66sf98+yfJ
QJKv0lyH1NStXR9gh28XABTSxMJFNjTIGAG4Tm/G6Yo3qm2KvHeJzV72TfoE1WjJ
ZyapLk9MJC/ZpAWR3cToz3bciQQnsceYoT+d7U/6XPdrov5TbITP191kCFqPEEQ3
eEUlHda4QXbI85mBA8rwIM61MedLJfyTodrcPsYg0D0OuXsl0YZ7HUZLqGXlxvqo
N3yu7aStuXSBdHc5+5BVi7GCS8/6+CuHYo25LYJcjVSKT7hbMsmfCnjkLkaeA40i
GK4ExJ5XngbUibdxE+0KTG1TQeP2STtNqVAh4vXC7CmSzOzp2zSeqm/IxRxyrrPV
aalFJ0YJQGuwd6+HMNH6KjVxrYdhTMkYMxA6httomOxZ313K+JwNgkLQV8LVkYBw
DmJ/WddkRcSu1NFBlh/hnvUOqRN3ETSzyDbsYFXIJW7Jqz8zPZWqNYj3lSE4e8oR
2Dv9cDnl1PcTc5XEO5bLyxJyLpV6CVT5d1rny06NsIZdb83Gg4xWjDXOJELq0HrG
OLcY+xXSQRP1SfQt6OUotiNYHXb6GIGWzEKjcy8Un71f8kK+9aHxVnV4iP8cc40E
`protect END_PROTECTED
