`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hIPIlDyR7NTTou/QoyjHzljdX9UbVu65PzQqAu7rAYWLnaV3owi92lRsqDjj8Xuj
ZA9JMhsO/ud4QCMu/4yE5+BlPOpqgkujXCq8gk/+uLbgauEVZ5vBii/jCj3Jw9WU
+2rYgyxxf/Cv9qxRWa4OsBPjhFTuYMZuV3Q3/EKAUzxBPEgBe8k0sQD6aso/mXKs
9E3+bOPdR+TEuke3Bg7nWq5qQWix0JaoWdVb/1HMghEDL+Jb0b8nb8mwuOZ/49Wg
Kjcq3+CRFC/c7ueKVvSPtq4O5h0SdMPGX3UG59URwhLIVbQyEH6gIt0xv78e81b+
O2StedpENGExvfcreZEjS+HiXKWhy2j3DEakI3jvGKA9CGPxnndCkHTjHWZsGuaE
tNFK8syslzLKQiHHlif0kQ==
`protect END_PROTECTED
