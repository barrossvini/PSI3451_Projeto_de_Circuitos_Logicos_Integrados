`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eiu9c+L+X91QmDK9/TepnR2DzHxN8WsCh2n5WE+a0PkmMpLfAk+b9NkGxJTaHvBg
RmMCtK9Bq1x66ssejtjEwtLBb9GVZfbccssd9OE9sqP9F4BWIF137VKGPFW2kPIl
1kfMyI7YpE5DB9Bj9GVs2V3Cit3GbjJuW5Nxmfy1EAGBoxg6SMaf7w54dAP4o5tG
myYymydJqRZ4LQeer4PjwiAVe7Sw0kP7KNB1IwhgublNURGmrcryC69Etz6nN1c0
8z46Dy2q1SCSkDsXxH/cd27T6VZWT57lOk828I1merYrfIvElrwxslSq0tgcj/i6
W61tJTuDXttGmArHusxm1OaVaTEzx27qzuRBh/4J4Mlo4EGGYLTj7sr0VP36JAGI
J6VFUa1p969udL1jG2ARsuCQ41dlDzKIJlnI/VF6INMMgK6siisd84V2o9Jd6c6c
402VlqLmsrX2HVmyzMdE25l0gUq0N8GIbnG1eJVM5hWxmwYvi+y5gbdAG7oyVTud
nPtrW7VIfPDMTKbeQDuQCZj1JNkT6+n4xojBq5rGH5hQRXWk2Hpf4sQQjxv3FFUV
4xNOEvzpJKqvm5yHhg9cbQiH7TwHvRM6VKDFsHCD5hvtrS/Z+mLOxwN/frNqI+RT
djnK+/Sv3qdxZ6iNnFBXQtzRWsKOV1WUhIAtgVCaL8o+QaPU9w7pjc0Kl38qk4aY
QiNuI97M9TH/dRd8Uwyl8iMIZDiAohBHHds51ElW1ju6I7O5JdRgK4NNvFL68IN0
5GrgIrBaNhuijCN56PCqrzvr/QBsdQElkQjEpy8Y5J81+tvdyk4RgbfX6aHlmQgF
xnjHI5WyFlRcCvnSJ1v2n/JsI3BsrjUDAy0bYXxy8TmF/cgRq+MYrbJGKJv7mjTu
XmGXAKeFPqkg24jxj/8D2AA9J2/5IMKJztOiVWHZY3em8nOabWTmo37X56xLivhL
nOu+i8ef3uuDOjJVppLO3FIpVSI3kcDnoOwBjbGX9bTL5warou3T1/4gGCx8IAoT
1jDMbzDJNO4SueyiWazscqdvOye+lDyUjFXkzNWB2Xj8t4wM49JbchXTb5bRn2eF
twEhQPpokyVlBFcpvdIHW45HZHeLW6u24RAGC5pLGquSL4OvStvFJTonBiBd4Q6i
idwTCGx1fdpy88lkKdTq0UwW1ekDca/VGlEorffIsnRszFI4Qy7ZGfYj+DcxrhuC
FcdqzJT4tn0YnawAyi2rWdd+OQvHaIT3xiD/P6elO7bKlZ1tZqicGe2afUFZm5pl
2/ECgsMCatV6jnI8uJQIgKSgtu7WRFDQj/8A8tRU+M3Zqqt905oXPoWUNyRhrV3D
PlI7Rd3CkpgLvlHwVUr5dH3CTuq3aU8rF66Ro+iad0La3QrRFJ1HQbMipviDVohN
LCvHHjnfVy1tnVqAqDmuAZkQxWzYAbLDMYZnDhPoPnBn4b2BWN9uz8M6yF++Jb+R
Oysi3hRP2Kyj6cfIgZUSLXYt8vU0fsF1KliDcRwBGuUgBfNaG5m7yq+ReLH/lYTC
sUd5LgaUNJO91p9CA93D3Jj0mL0nMFUs5c3SJ0TYAZuTZCelGD9PdAw6lL+52lqT
j8nH9pV2C+0vCVdNphbh0+jy+CyWDWESHss2TX7E/swTCL1z/JWsogG+jOp5TL/x
TewTHk+c0JitGiVhQuzLne1qgl5CFRA9C7YZVH2IuWOQWBuB/xxgYGF4gC9iB9im
W+Pwq6IeuiDBiQEqqUGraQQv6eJ9o7LVps8lxg6JnVFNGBsKgJa3wU8z23YxaYn6
ZF746VRtiXXfZAwTvOuP8upAP1zqCL/R2lz/v/EQ7/R+bHOcGU0IeAN1TUi09DIG
VRUyMCRGkb0GbhZ5IKckHvC7PCSX6iQn+atv4hceW9DjvfOAgL5CbpdlmBIBKkOP
AF1Z9Xu7kZa9vFH5VAvtQLxtnJOM0+wGRTLQR2ydIax9Jce40wApSjoqiJ3jskK1
i+/lGB+gvTZTAOz1w+ObLXMowwoUGeUmlofmg1oQVy396izEez5xg/zb3IqQxDgd
nE5YkVRUyoC4pjn0AT6zXv8dytW68dFRIcXuwe8Wg7CA7Zo/FOxkwabJ6VbEUb/P
ZBUiPE0lYe1QMNo7J7hqw+ZyndghwxTPK31AAYBDpz7pUmNxt6Z8g539nc4t92Y1
F4tj3dlRpHZ8kFCG32AGwTSGylSwwLhWUpWp3d/T2trXHELSSCX32jd7pm/M79L/
ErrrcigCM7gToQT35yM1rPSHJsslPVvD3tWl2ywFgh2rfmtxczeKaXJOKE31YYup
ajVsiiSECOYsS+CvsVYY3H9LWXDPZAIz5TN80oz/zYJv7B+kENpYZ0J9ai3Eizx5
mb0f+InV3ggkmsIQvejG+pK9FZl5X8eN7wqdAS/mHuXWrvYGG3wEdd/aAf05G2Kf
wDPgrmxdzchg2vLqDTPsD9DqeF8JVwVToqUY863vnfD1A68/PIRukZqmLh7CdHF1
/9iXwKHmyB7FrnKcOCmy5AyF1fRzKNEwZMtab1Ii2vK0y0kts1G/hKu11ts+rdzS
ZE6JlfHj7f13IRPtnGuV94BQdXD8MefY1lzW2XZOnnVlbG+nY1wYwJOrbEu8f2cQ
wVba3c4HmseFGrvUiYa4FfeX0iKCBd7cz3IoZ7MAucUzQK4cApPEXyrta6Tr4MP4
pmjufnHj0DBVgzmg/q9cx/b2FdJznqSn4cGNWbUMncFWn9WGpvzNS8HQrJIZYVXl
ij3cTndKrlL4EJXRh5f7K+ZRYJMUJvOHxw5WPqXXXfpCZs/27aQoqplL5KMNNhzr
bGNltapBnEGxo1XbltfsRfO95ava//yL42fWrhI41IVUg3E78t0vWfIZkieqSeOs
y1pA1bEnNZOABdE3OuW6BnfHjwPeDrsle8Qc2/yF/OQCfi3ZT0RmDZwNldzj/aGd
qnH89HObi9HLASchnu1CYZiDPg+wnYIer67pimxIQI3pE1f9EFZ8uc3y9j7nXoHf
QAkk8/rtg7oK3RcA2+uS/i57pRcPEUCStRO+p9kjmX8byCgci9PmR6EYZeLx88cB
IyZviO/Hp4zlugpFWM/AHBHKA58XLrRjaYMJCboYE4uzZhX19Dz7HMFJadfozEgp
qJDTQs6SeYTPR/ZQJJbmuLZzqiXml3S4lO97ZcwNlW4HvwiOQHWIQbskABDSa5r6
HLQ9pSJiexKx1GjBvtmxtm+I9DVo0sFRBfLflD5i79PAHL3W3lBOars+6R3zYkcD
ceCabYl7QhPVV7VMGQTWlFfmH6WkcqgA3vLvOxYxpIFUT+mqsyWf3q+LM28xHc1J
00UGJaulIkbhoc8hcfDyWXeLRTeukub8kP3cDfP2EHvQueEezHXZ6vZ5rF71p0Fz
zgC4Repoc2Z7ch6Ib7cwg2ZZ6dRb6cxWtgvF9kkXKsEH3PKWIR5RGIxuxWDdfrMs
BzluKN0UnDM1QUY9Db2/gCbQ68VSHyHr+RgTh5yH2zuIgtp1/OQvVLGo+R2PQq3h
y+zU+qQ7qBJ92PHpuQcsGwCytzcg2oYtQXQL/Ra5jTJ+01BHiCeNHkJ7cPinq9PE
Pho3yHr3vEV4+ifEwMfEhdd1vii+TQKC8kVmU1jHQ2gLQF6924q9tuqjluUoWWxH
jhsk/N65+JCeFmR8/zv9MJopaJEZWq6F8kRMGN4YUnM6SHd6+11kdJxjp/pysFHc
98Qhp0r0v1uRF9og/GR3WyT/S+ZuQQIisUnArp/QLhKBRXGbNMW+FmkJBcW921dr
p5E2D6e/3S7z34PpLgRs0s8ptsy74I8ObKgWA764dqb70jAVTjShs3gFvB437/4F
AsvYjqOg9grpic/UVNI+9i4ctvh1AlNOLZYY1FNlIflnMDhOKDZbHuCziwHvHUeQ
ri0WULE6HteFphDaIlFDfO9v6AYNSgWf9L3IMWrbyt9k0j8MgO1b6zyaZ/KxIaOh
9PjwcrJa3KbOL+evaSkiWB3ufcdDwnp/0wdKAKJyweF0BmKeayjtkcE7QSDz+BOg
BQMx5lDe7aYapEA5yzaaVAYu5FheCuSIQ3pd9uTFfETD6YNe1c/uJjVa4/ik3AC3
48ONbDKtHyAHIAmXFQ/cKbmH6EYUATck8sZBSfotdLm58Vj68JH4Z+GSxUl5mAqs
+NC4sucAQI/+d51O2HOhfSD8S8ObQ0zkK5zn63qv3A0M4iyToAoHRthvUHhfOdbV
VXTuLK5v8KmwiCnrO4bYn91eyFDN5GJduTvx2EbrLUZpgs6q/ta6WZdmggOo4hCr
tuEUsMpbBUChcR2akidpNMM0yH8OYVaHAYJzjbii3WU1NBOImaS2HmKXgXpnSMbW
idCX06RCFZkOgyxMB6jDOfT3RFz/cyymhYgoMoRHkSu55n+o13ttQI+9lsNCHcTj
RkU5tzQfcAquDtELigrb4YOkqTGdlBBMpIM2Lc7xKnKjzn+jAvazxPwMz19nmjbe
Xcb3o5BsDWWWMXK+AEeUz9yQMcN/qMw/WOq4hTY4VqxGpNWQWGVPvmrOHNd7RtEN
PWhhfniV2huPsqTAfHx66CgwBcj28vCRtNK0xEY5UEZ46Jdp6Vu03/R1CQ43jgEI
IJ1p0MgeRy47RIS6bfRFVg==
`protect END_PROTECTED
