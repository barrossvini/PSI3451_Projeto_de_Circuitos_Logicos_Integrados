`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HOrDSroBQABqmTVx/krGh9BilfKQW/S1Xo7MrWPflrwVnz+DBT2GURe7b9xIM2Xn
BlGkkeNdEEozl/LJMPsdB8LT388eLqc87uZRBfZaNqPu3r/nTrcJFvqmUmrX14H1
S7IrBKym9QyVifbjFUkKd+k+E7acWpSLcgKAkB7ms6PEBgwaAdwQJyXgtAeaNVEd
EnHuH7YfbIXytnPlw1ij+rPCdi5e5GsSt5izLR7DuNLsOKu8aOF6i8YMSluSzr6K
itZlH5+A+11GPKlcu8rAiSV5m5aG0Gw4omm/5bRdDxtU2t0Vv/dKEvZeyMlZPHvr
fsUHgZTbTSLiguhVhM3zlDriciSFaRuvkavJF/hKESK37IaG6NNEiTSDUuf1dAa5
Cl6BrM2uJuIWd5hpyRlTcIGNJYPIc0xrdEqIRKkPNS9cDN+JrnQg12H9pytZ5FQV
JR8uHLTkizpZebJOXbxd3xgsWFyNd++8+rEdlqgufY3k1m2A7PF+kwYvWHSfqjui
ZvAdT8Ud8uE87R3UdPBeVaC0o4r1gM3Q2KrRxpjzuxUdwnhnceGONAQdqhqyedC0
E8mA4XUTQuie++tZuL3Xb2Vq35sJRffyvlfVoKOQC91WQm4puNYnhmQ81I64y+iM
j1q6fgcGnuAg9z6MmvXpKfHY264fjvhO6A4x5dlCSH40t17m5Wc2+qX0jTc1wTAB
rM5QTqlWA1VzfwK6qQplYSey6/wXvwZRHdzf8nV0fen21j3Hacou86MGVHxxInKv
OPQx+WYVP17rAEKF6HD1KvVVXlNGF+u2InGrQjhA9zZ9fGBzXdgXYZdzcfu9Ke29
eTw3mYB1gfJpWdXvRLuf9ufXlzzMD+HQFWZdMVj8NGVL2hbeI1SLlNa/RrtdrFH9
MaBlwLPGullZhKuXLpTX/qliXkT/o66LSI87axA0cUqdO8cVdTLz5WtAdmjhwoVT
LN7xBJHR3o0GYBhGeSp8e5fH9I6vbGBDphzpd0RK5hwVtUBNyEcDtX5ldAdz6Ovr
h/4XjC8/86W5HfGerZ9hPi37LAue4z9xwGpUXoQR1nWQ4wJGhDY6XZmPu65AJXHN
/D2pj9y4R6cUs/mAFuybsc4usLmsfPpkfdJTQxrJbaX5NXB9jn19Pgk4NW+xL97G
BZiBBuF3j3Ep308nHabxsKygKXxkfvo8U+jIaXJSgmZ590O/+42l86i//4LTY0nF
lkBGNHfEemfwR9cfgVgwtQckTxXOLLxa2n5JmAVQQTxPwMboXKWJAQ+AD7qd7Xev
vYpmgJC1EsRFvIZ5F7mNphic2z/LUUQxjTQuLZ7rOJufLAf7W06hC0c5LQF5evs6
DP0NiANY5GMRwUyzjPSii7VKdDnwBQfkbfENSXCgZ4ZsllP+kooXiNMiSyE1qg9h
HC5YXkOMo2Y0VjzOW6z9W9IXTw404rAPla5z86gg7tJPNLYEQixTv/w05gPe9Vj/
bRilv7jYCFtY9Wnhii9y2vvUnZps9I6BjKfzkWN2PCOMt1AzED6uteRVvdhB8x3h
vY6JqCV1NyeZesiektP76t6LaXEJxLG9TcSsJSXsiCCevRyFT+J5tPyMZOwX3NWs
AhiSYEpqvKNOhCPJZnY5dy+zWkqzvJOibi68WPt3Xr0rtF5zBDP7D8YB3+iw6GWn
66a7JiLIw0f6M3vr2yrFXZsxpn2OnX5JsT4z59fQ/ivd9hKMD4xgsvTIvUDMVLvT
2GKAfa54+XomIFF/A7AiO9amJswRq6SGpx1zURJI7MXbGNxKZZZwZUs3tEKPy5fF
tSBYvDNG8gJiK1FRHSxOk2RWhrA1LVKWFtV14F9qIojC8oJ0tGAAgib9rJy5K975
ygIwvokC+mE3X8uWgwDyRX4pyAe/RAornCZsbZsyzncpwrZizStH05khqvl+NLtH
YJgpGjSdG1zOdJBxHigWqen0yG0t2cNxg6EqpvPiN/gJbv+AcaFaLh/yk9h6nnzS
8/kLnrQwSsaEhQse5MXMT/MO4sKvmgVF+7/gLP/aLmMpDfhRQHuIoh0K7oFSBxW/
Hipa2FJH6tIU12swWvPAfiSK1gKuNryWQ6wOx/ExO8rWHlFk1wWzQGvbF3ZaAc5o
b//9KKGzAV9BfwH5wpUjFXEJBMbclMyb/fJX4aL0n4nwvoP/6b5Q2d9L1ZbKZOQU
qJ33irGEJxNOCBb8NaK/EWsL5WUTweDGBI7bd/wN21XYwqweM739GWBjonNr11yW
4aYt2AnehPSiRtOa+IaNOX9xyjvITC4hBdnCmK+OdOxKx+csmnua+d19OKzsY1we
vWnFGQEiAD0jNOm292rQNqT6fESOD9BhHpz2nvNoB5ltJ/bcYaItyDENcZU/KAom
NwvoaGD1JfYlBl97f9r4+mK6mNvnemi21S2TsIHimiUDPPHFGrF0jSml/X9eN8OJ
k7CFdeccpt7Bpoa0cyfVSCLnlKVBddBASZ32qwnJLt19qor/K7cvuA9oy6kaXVBp
FqYSrmEbjCpEYbtZ4U2J0ILCo+bB1sDnlXcMMWo8wuSFuv6iwMNioaNKh7d3394I
SZiqxjmV27UOYDQBZPjRiIy1fF5315Pk8a6S++bGltcRHoYigwjS00niweVw9CrI
xu70H0cuyBgBVwkO8JU64ZO/yfllkU4oqIj1iGccUdwAXKnNHVxQ9PrU6K6C6yaJ
GWCSsApp1m9e09Ic00dnlLk8aOEfJOb9jzKcSQG426rrYli4QfbBSNCdymD80iup
rgYtpBww8JaVnInW00v95iTgqfqp8wdRwizt/b5LjI9qztuuD89bLmxKpSsM43e4
OzgsxUMpMBwv4a8hSRQHmpwryOAKqmDk+Pnw42XQD/JZjLTOIXKA9ltvGPeXnZh/
TvIYMpri1XXzHC2fqVT6Inf16HGd/srtymbdRth3kPJP4fZPstX4IsFzb5UZtOS5
R+UeK3S+Y366VwMWEjMIlwrgAtK9WvhJTpvOEc0spATyigq3rB7gxij+3vvlRTYS
MuvNYvhpjNIsLKTdwFvhN4Oy/Rix6vOvMdw0B9kuRrQdnCX3UVPNX3OlAgmDvRkZ
MWcdV92C1uMsybNG2OQBum+a3swWUAsynOXholpc/wZGbvBF8KFD7CLC3BLWTQSF
fTtdkGxR5cvfeWFOo3JTujVPJkIdMgDYZhT0JIZdO9Gn7bTa9aSO1agJYvzLwcxA
zb5m8jlh3Z9Mh+OsvIjramOPLqjPTtVy/Kbcrf6IntkRMefS6r3PTxUF4czk+onT
mPK2eV6qC4sx+VKuVu1Qk90up031S4SOrFyb18yS4iz/RwhA6NfquYqI8lV32/K4
OJu07+qOSgS6cSWyM+C5AvjVPNH/MiOOoUzVjyaKwqrYQI87Kh6labA5bJflnAoj
9Mta76ZRA5BTDig+GC5pqTj3yht/u4kD0iCepkl0LOJ3HSk1C42UhtTpcb7YyUEs
f0PVgQGyEO3FoNglKETTA+1NLWrlcXkMwgd1z6z7yXS8QhsejPQteQ4x0bidANc7
hIOFanFe6TL/Iqychl0dSae6cVasvv1IRvvWn2vvE/aMXNA+eq+wPzvd1+W4ae1u
H7JPqvniM50xXhWX0bA/OINQeffkhDQY45ULkEpfN+dAoiM/7LVL1DYLA87qe5y3
UZ6JEglZ2OuO7lWjdkh+xw==
`protect END_PROTECTED
