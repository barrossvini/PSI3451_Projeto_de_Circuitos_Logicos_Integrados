`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Fc3wqfk5x8XFHaEa92IuyU9xYB+AtBusBLufbubidP4E5B2Zr7cVeDa0gV1JMQJ
QpbNs9ebFP5V3y6fdW+5IUuwnA1gKDZlUFxiq/NhhREiFNWkmcGdiFtlNKwtuSST
hA9QFvYsalaQBZVHR/E2uZ0Se0GqkRlWk423dWHEqPb6dqmCblmWNdTmGHYh/7dS
48jtZGQ2A3FtxIgGyNM/m3KXazdUC6cLx9Fc3if8aj4Bs1FQp1iG2a6CTPhLCqyw
7f53APoYvwxGFs3KstVWMCmj8EiD/aRgVLjyQWXEBp2iD7luL14Y7YfUx6Qd37NT
oa16TlS4ybddVk+k6rFHYpPY1s2XmT9qSRlUSSjdAQMfWzr+nKdCfeZqOOC/BMoL
YfloPWmL4hw4BpCkl+ytgNApX/K1B1ix/JEWo6OCuQbdzadEGFXiZHhz5T6OQdLQ
gJVsho/HF7AT2asPhtfhNHpJBvRWhp96deh3E1U4RnAEb1aNIUJs/OV8mCXFiEvE
yJrsOxa+i/COtYUcLHbIiF61I1w9kaWk2h1ZuaB0D1AfnrXv41VNbP91v/u1j1W7
kU5m34s8sPL4b9Mwg4BPmbalt8R6BMifxgLBXzQesjB9nOv6c7srKGt4iSL1JcTz
MphlbKv50Hxk9AtwYxkQ5YuTTDgcgZmYfX+qe2ympjjy7rsqwi3Flns+Sqi1b/dW
T8HmIORtUX2IHhXNfb0NRZswjasL30o4uyZafLJ8cF7T3C4YSNfAF3gDTwHRkWM0
uZhCXA+4+IzHkM3qS/N2dGnW0he5JQzc6E3S2MgfnATrXACiNtyRYe8ln8ZgwZ14
qYwwb/Z0dnTVtmMUi6jaMTJz8Wo3TtPOkOQy1bcm3do=
`protect END_PROTECTED
