`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z4Je/wN9Gm/QsSlz/7/5FDVX4YwU5JbX8keGJq9qTAfLkjcQpGJC3Rx5YCcAIPRI
xT0pAFFNbb0BN+N4AOfF5vLjOta40bwfJyQYPcZprkX/ASC8Mg3Fm7e+RDDwcEMF
+Uhpn1gN5AbyLTRP/lZyoZOd36YcfF3AaMHeLmq1Qt790Y2ZgJUCgPXMfhMJR8IA
6UapOkRWxn4gYn5dM60dPGSyZGzL4CG8u1+EhN7HIket1elpIiobO2ZkYTX4YRR9
4WzGcJv2SJKljrBG6PtuPOeWrW4mE4ZsjU7H2I5nYXUbvL2h83DPW+ZT1Pf8yojx
tl6qSr2tKZQx4i8l/6mt5+8/wv8UD+3MKMWt7Awx7359p6OR52Hmv2vv+08hEcUR
Cxl+LUltU776KKXumSf94Qy4mx3sLq1ov6o9UidFWWj5qxXOaKmn1KM5HreSXoh+
pIi91De+JkX4yaLSUO9bcFRemXtpajOiopNssroLq2p/7nU2pBUSLEfeyrQsMvlt
J33HKZxUYY8ZfwsKziZHQPtGYubRswFaDYgPHYwXxl5gJvBWGxK7nR5TAmH4Kqzk
nQF8adZSwti8HU6RRYqH2diaxu1oWoNLVQghB2IpioT9i1RAav5BblrU+oIJfn9/
llLbf25tRyYDsJTFBZJ0PxbfrJu7ma7GEikyGyFkkUU3cYVJsswgcbe//t3Is63A
SC1PS/CNRt4ssM0y38cXPH2L533sO0h6REqQaEH1FTRyUTvCBCwWf2Foyvma+FCc
B1JOJcYD53UqC5GqAFyebdi2rWOGaDIzHJTCgZ+2ZdCLpBr7HVsD5a53/tdja+Yz
4w1IXTtXmaWDpXexXjLfaFj65+5NvT1wAL3ePdaBgqDtUQDxj95BBjemMXJ2UwxG
lenOGB8BLiI8XZ06JmDqAj/AQq6v448HIphTIquRAhavg5CxSu/zAjamoO+/v5ay
XNPmNfglXJbUUDfxuNGGzmFCa2KFtWYAM5jxuSz52Q4Uec+C0VxZBsb7tKfGKq2V
DSf58YxhPKxLUnJdOQ5eRkhtPVjmmhO7IfksMlKiEiiERBylQzhHSNHBiIbRgRr6
wSzusO4726jCkJLpPhX0SMfDXcGEoItyoqyEc4e9AL/rw4qSJHMkVMdbjkV2O6Ma
AzPqP5fEbP0gH9fauhBemmDkFBpdPTRoS6/Qv6nV7pXBaJJXV4viAkBCNaI18CG+
9VjrhiH3sSqnAuPtNAewRstfzOHI3f7DblMt9uN3u3zS/STQlXj5QH+SfHXUbiXl
VbzyDg+gKma2V86wx5SQ1/RkFmbkcBOa/2vDfmwrL4rpsC1QMSCnmyCwzcREaZfq
1O141coPR7nPwNZ1txec/zmSoEgI1+3lnWnGEgNAoXWxWhc7LpTFFA7oUUqijQPK
jFg56y544TU92OD40k5puxKbpg83bz+PMWK4H9XbNlUKE4EbtOCmPKFUIEJMQJqu
v0WeGQyQ3qddomBiwXL2QAp2pk0LSdaxvG1lBEES0clwGNZni3k0tpN++q2eLVAR
sEgm/f4/pLBinVio0Oqfig83LV/lzVtZEoH4S39+OaeKn7J53qTYnsSoz7mRdk0c
voo00WuSTftZJUbr47WBmdVF2O2vLqY5+uZng5QcydswGNm8M/NMT9YzDmOm0n3Y
elfk/tXM+I1EVcCas6NvQitT0kzBCaic4MSYT8v3SLwPmZGnLZD5FHT9rDGJk/6x
UQRMVnVNaabWGUme0dpk69GjO1wjqcdOZcLZLZUl+jvh2Mw12e4wvAqFv6Bm1grT
mCeC8j9HCA1+O+YaL0Kk6YMjDQlkw6WJjVVPs59iV50Cjv98ixZbe6nj3QdzF536
EWpUYp8tsVXNNiqOAuvLMVXkEcVh0GIDiRK5wTyLsvbVEBmdldyMuI7pkPBA16nP
fxtPclVxA//gKoRQPB/W222c0znfbJc/h+9FBu8RG1oJ6XOvvaEb3xNzNPbehX+0
Vb7bXIVOtxi92Tuwg6z48j4GkUPA/m5FQbSTgo3nokwe9nln0ldow2Runeu8dC6b
VW1jFTKgt/9Gwaakbh3C7TC93Q4YozisEZZixoDuHA0+6tz7xel9fN9sGahm8/aj
d5r/QAJC+2gHSOTeYiguA78pWwVMTru6uBUC4uQ/dPy/us0mzhqSdvP2lpa9PlIH
KVvR7suPLSwdAkeslMzRhT6Gh4bEjsWNoiMoh4S4V6i0MKon1uvHAFQqSkqivfyw
dI3AnGmgEPwLriRsZW+AhqqIf3jF+mOuImUvw4GpXtzJj9WbA8ST8cYnb2tNdOdO
yyZz0D/5MiFMx15KuuOP6vQTT53LaWT4v2xFeHyUZJ3OF8BvHZnEBcMrSYWZHXUF
/dCBADHJ3yGnZ8UDX0BGYtyjSzEaO7k2BbjMdqOgxGoeHRHh44R3P884fJMEC7tc
IiyvyLgyB2tbUBSLQtX8oTaY6mnmQCbEKr51EbBTgZsOrdzZP85kMFLIaTZ9FP4K
Vj5UnLS7Ta6KLqydRTJyEetj/cr4K1EkeTnkGrPfchlJkq2FJlGDjNomalFb8DhR
sCl9F3lv42X/I1OZpS419gJvVp49yJcTllQHKGzB3ghNJVM+u09AZnN2GxB6CswT
fjPCC+QUPfXM00p6ZguDjRf2klM9/zvIpmi6hhzoh4Yg4TCJ+STNCOnbSGitspMa
Rk34aMqK7JAL9JSaTTNQsiGrzkVdKnMQI79g4zPmAP71MRzdjnI+yA+L+VE/lPAF
0+h24RzT0uVWknWi+JRoPe2qc3kUEIVwhth48Wsnh6A/1bB7HTJQWs07OLVmktYR
w899QanDqSz69ztAJhTuGuJsTXCINcvRZfA226ue9XKkT8VdstF4R9vudOGRawpP
LHjBh0J9M6Tp1fYVfRTVdMsOOhOM3LUdOYAs8kp0HImd+lQNahtKu0EgqWAHJW2d
GfTSYGWk99mKQjlgPJuttRjnpBR74GAbPeUYy4Kafs5rHHzV6qKCAh6QjuAO3xVC
zAKay3y9snJBuXcKw051E42JTRRJknZz+2wtjr1h22WSHU4zdZIaUbpaLsYhDCHN
HTnarR4Zzb9aKOXd8TAAjt2uuhoN4Vi1LfNvVL+Rqi48xrV1WVxwvSRX6uZOOnqv
DvEY59NrUG0XPOeYYIEjZpYny7NHew3tQfWq3DV15o2y659IffV02CkxI6Fn2W/B
EtTVJfQBiQISOpwGZp6UipeaFbMtRGnFDLSV7qMfFgeMvENYgFoumI5TjnswEWmW
1FL9dF582kEv629+z6bho+P0pzQugbEi3cGCX2ODkJ2ri5t2GwmEMgf9QqHZe8ty
fQg4M+7sVfkWvBmxu7CqkwVWPx0Hbjd4eufb6fwvTu7FZIemT2p4ebrOLw468pM7
EJnNsQWHEv05bf7DTqmvEMIrOuIVcoFSmv+pmc+6du7OldL77Adz9gZHy2CXox7n
R454jCx9CWzT2YyQodfYZskLysMQtjDsrJ853IaCqcimYAfjOSWGI6xHP5liW067
OvvYRChtHjxxrYJXGN5A5QXM3ual22xyODvTO6yWgJpqpXAs4uY1bfUp+KiYQsbZ
YLKvGQfpa/sSPYV+N0lYHujh0gSFTCk7c9La3RVj+DAi7mOJ+eac4BAd4nGBwU20
CAz9n+7n6l7t4KU+zRyEjyG2RkMZdFTv25dYdDkU5l6E3yihuP9U3QVH0IgSQT9R
xXnb9gGghNKCmpijBFEh5FWz5dlboRUJd/olq9EGBXPQhS35TACw7xmnEadbhxIk
xfH5VTileS501f0O7W159Wa/yVpp1Y+AP5/wABGWJZXP9TW9f007QsUNVN0WVHBw
G0qTZvDKBuTMhrJmyFy2nr9EBsv161DBA7BroHxyiON2QY23DrKReVTRGeLswnEA
Kz0Pgx3pAEOQwVjtXH93vzrWYUds1H1wBSKo8QlDIEZwdTljri0G+165l12pp48u
oXGyfm01PF70iWTpuJLbMeDHK/e0RnKYHcGpWJPHc3ruK70rkEB2B7cAQsQBZAvN
9E5Q3y+en1D5Z2mUzguDmi4C/9GT51Y0UGu6+0ULfhMESDxsnYZLjoUZCksELcWj
S7occALK6boX4XO7+4DTOJl9UPM0x8k/Y6f7Yae8amFn2zJjhx+ggBZvMl8Ihe1p
8+BwVQ7DTbnwE7zH95ATxOMx4NlLiug1iMIJrmsR3O74Q5efFRabaD9HdaGXxYCA
pzMib2YIZ5Pvbh0cfnkDCM8w1q+vdfODyRMtTYyB+HTpwCy1Mie/ydTH+/rwkSZw
+INPS5eOkuVILoBnl04mcii/ZUNLdaU40nhQnfXOwwxeyShMsZTCA5NhEeF6pjTj
obk4SUH5rvppsfZvwPVy9a/dZtPQaoREdW0LOPFmXhVKa8M2CaRkH6QQZKHHWPyi
eI6xUNe6WSQL3BWoikouYUxwHQMeMvkCFvOjlkwyqHOBdrNYfPxAKpOTf3vpRMPv
ESjLrAVb0Xg5loZ/h/G0dKyUIgxWs64pf389qf03gNakHg7Z73To1bMVGNejhdSC
0M90OO3AzWLhfeX68C/L1jSKe6hInetj3wZRMTscUmeuGvI+Vvwj/ZCZXgEYKzJN
2F85vtyJX/cweOo9yVeew8wFaYQb6INB+yp7u3yolwq1L95fobwGgJvYsie6hvzi
JFL6u2/Vhu6oKQsjadWxKoJ9v8nDncmV02lvMxpMQ1pvpKza510OyQNlOgWpcUZX
8RaKzapGPdZJ0/qB/Zfw/IJXrGLxy+qZIFVeioB8AcE7fWZ0Qm2W3GHjb3u9mXqY
VbxaZSzel6OwWbUnPj4tTqDaJDtYVO/koT6K9OsC0oTxibNGLoNexQGYonsECuae
c9cQUOChKOOKZgfLfUCJupnerKaLjM4vPqMGwtgkjO94HmzCB7wLCklPW1BWsXaH
l6dNKrnoAqP60+jQqqlKShYZLzivlGy2OnL65xN3LSLP215Vc8PxbTPpo/PSDLbN
2t7Kl1wXFH5GnyYyjxYNXXvvVa0vvrieHMolCLTrNBLOQFXBkKw6LptS3Ovv/+P+
xmBUAJtWE9j/6I5ztgrjmSUfR2F60uvN2ancH680TWmCZB8v9NzwE0BVZpwK7m0U
Tyq512VsnEwGug9DtOJd5Bg/7Lapw2yWDnZufmxooceYGhbUM2JS6w/MY68IKukG
3cOlrNTmiQlCr8meEO1JDsYYlqEbR/Y60Xn+mUcR6hjvMzJ4qn83Sot35dOA2x2o
sO9lWSEiIYFiC/RvjdmUV28vx6NS1ML3t5To+FM6M4FgLlTW+v14UCduChFlquZ4
qhZWw5eHShVrchZoefN7l0dCfWDfnb6ubwetHC03VTdFfdUAMNwglSvYiFcVLDb7
PAoR8D4xZmxWTuS0ZoiAjmkQNrm9Y+KNCuoapXtMFvmaEvOevePEyjxk7I4aTdrV
i6rmBkhup6W6AW/NI40Zbb66Qi+SHsNIGcQd9AFTeytM9OPt2xCs3vxaKj49Ougx
Dya8RA8wfiZxgdnBvCHk59XsghcmPCmSJqzJoez6Hi1Pm+yBBoUMHJwcFXbxpNgX
fk0KMJ3fZsKsfPUDUNQy7sl5VYtJpTP8zcjYcRFwtxgPpIWSP98GEoiglcy05JIQ
qD7dxuaxv0SDjGB8yUqhQ7/HJU3wJ2RpktdaA+WA/mcz/mpHcrSc5rKrxyymYy5J
Rjp5b8UO/MX+FY7HmOhWkQuqcmiBtvk30Db8ENqNJL9hsxUdDcK55huZS1Nq32YQ
d2Hlpm0X/QoOutwBwjLEw9AZZuGc898/gl+RaHe8Tz5a/bXJaBnnzYJXRfXxciMg
DjWMvEAGqR+abDs9bFlH1CGl9dO3xpnYl/hMCOf/gnO4+5Wf1jD/sNGvgJNfhYJh
d8RRhv1AxwdofTGv6Wx7Wpoy7QdBVblMjlTKlhWi5LteC4e8F0p4O6gOqbPKsQBR
LVztuQutP3K8zgrnSxbMIvL+95PqrkCLfRigJejyrQg+czhh24Cwjg0N4Od3bw/o
nmuVsk8vixnIJw66R4ZVKDMHAnz9EXwwsFk0AuxwkFjskhaEIVi0VZAJvf48Ucdl
3xgt0PwnZnC4pvNlFz33sKiAxaHDypLACJw+DyBerBzoIStwkuYJY22P1C0X17si
49ZE59vFEMkvTgCbMqvYI4nbaTCYC9DsIgqnXcdVOipWwJh7oym0qdz+F/1qzIqH
NjxFV3KQIidxVHCOR+8FO/xsA8fwhakuoDrrxMi0sjtGCrRwN8vWqtIRvgsCxxsT
m7W916FaRB/kdnMjrH7rSybrUkPt9B/KZDVh4uS9jWggpd9tkkvzFgbOyASfDtHW
ApGNGYkQMQR+rBwO4cMA4M1WvOuDU2Xfo3NrX5jlxLS1Ld9UcZoTSNdJFmUdqivB
mBojkBhLuZYNAJfgWL74lUEF4KLsifDwVJwNcRLyVXvAbm1Eas2NReXw79MXEuX+
PYvJF0M1rN0nf9oopP14F4kvoxRol0ely65WzF+ON5erU+FfBYe3BxhmGb5UEOIz
dAD+NPnSQfADTlcpm1//qVcP/7fHRADKfb5NDrY3UwTkiThRSrsz5zjizNxnY/Qb
w/RdSUIv+i/RjHvNHqTUbf5GZ347DgChOKOBbdBJpJGGsfImu7KKCFtg82BvHhTC
StsGzaJPswwhtUnTegWV5/O5w3QG8dOA+pnGHDykLuDmnbPjfZjcBjMoF4mpPImd
GPQN0ZMRdNXQel6a+P13tJxya1E6gX8sJflUzS0HxPlF7qvw6/ZqJlhzaNYIKrfp
o3/UWAkGBZRq1ICX2v8cwyHUIhtMmxd/6/UXV5b5hlekjL1UGEP4QUOUv6pxY98q
h7r3uqX8sxi8v3pLsYuIckJ7H+UxYslRjs5Hky8oDYWxjY4HjcfTkkHqGlpaGqeH
0xO8f3Pc2iIJUm0Tkf0Qm4zWhPTzsPOOutUW7afEtE27ulMtlBi5rMVD0uedzSzk
ZxK5/rHdb8wBJGIcK3k1KE5wfSJWTJkOghs5vybYG+oylc18j8Dd4GiGo8UnIM2T
AlZhydIu7nC26mxD2P9S6vIdJbyB1/Bd/2rebZSKAY5tSGl5Np2CckD/i9+I3jH6
/rpY8np5AwhoXMJdwVWJQs0Zcg3lhS4i51VeqJ/RotwbV+ZYOnrxiPx/dSIlkQ7I
rP1tSm2owibBq5e12d900R0esk6edsF80Fvcz4C8D1Yg3XZf1GAIuBlzYrPXNjMA
MHhSf2NV8ZSE/heAn2/FXNTVRhl8KFonBHZ9ymjgNeX06LC9CNj6U2NvtPcTSKA/
Orsj3yTZRauXmhTS0YrpWO4+6Ncb9UrA/vLxPkA2j+SnhJEb/Z/0ALpLR1yO0wTY
GH/ZpF04z5b+ZnH6Hxn8NZWOv6Nl1bGSFEiv/1VmQT9HfoLm6SX+xzP2c9rNaz07
PRFBMUGOg+Urtt/QDvDMke4y6jPgEC228+wOHq8j4yi6u1FulrdpBLEvMJsdzwEB
dNvdDOtJXs7H1KULTqwZf4YtvI7bp2uw0jHeRw7x/Hu/gljfIcB/bK6D5IN2GDCY
IIZo2+VMuOq/abmLbWo3Jm3VWtgI9qlt8CjOpLNYaZVcewboZhhwBuxpNqpBHIv1
Bu3Roxippwyie8PtOF1WXKXkCe95TOPl5O8e2ly6/5+u86Igbb69hS3rFrOKRp0R
gXyLc8bWQwEekiS8LQTjtF4ThPaiuySZylZkc38GWcIunMLh0NcmsfpNhrs/FkDu
pQaTytJOjmwqqtEtug0XCBif+pj4ertonG8Jt/7iy9+jPbEszlQ5gLkU8fYogArr
kBi8BIc4q49PWhR5vKeRjDNVpnSOrFkKt/vfm2KNU92vgB8ed6OiHJZ9/uTHG6lh
DYiV3BdEN/ly07HCcsYkNZTd/6Yh4Dk4Uzv3yqE4yVr+wi7ROOLmm7qKhnCTSfLm
1e6TqIr76NKIW4J1tJa823ovzDo4WLYNrGcXzRhqidZeSgVkFO6X8Oiusj5Ggwji
udlKpjTZq0GIjC6SytbeCQtLSPPhOOGXpt8NbwDWtWNneM6AJ4C/rqPQBLmAixD+
LMpPj1JH9uYoxvZ680CCdIocLDHP3HBxp+eWaCNVqXVazz/zTaJEokrrG2tJ6f1F
/7nb0pnddwpw32zHvPNSRAjPjegNKNAK01XX3tneTG5zf0d0IKL4giGbrO+jWPrj
e4T7Yae5kUrI+o4hZLFt4U5eTmiybG6lVoTzJVNi5vFvfe1DopuVj7C1TbmS1O2m
u2Qxprokwj6Ctfxu07P5lBhP8xb84vt/fmMuwgFUN2WBn4DYvcbzD3sv3PguRf50
IASgyq2WXn+O60fKdtCb3PoJT2raM/KSA3PAHk1RzmQm+o6Na8VhCZKNCU66FE62
JW7Jg+vAcjG7KlORQr7YzMOlUWSGQrlBkVLMlmpM+g+bd7/yEgtUPCRzESvfT6FQ
IhRu9LEzUsg3spYXbbHny81wMMKoa2vmoINEIhQ+y60t6n2yjThYkEWP2tvX7n+d
esCyesX1HK6r9J8KcrzGQ+eEu1rUf20uOimTLOS6FBFkJUyIk7t+XzvE1el6YTt7
YfAihzu1LM3d/fAcnSkiU8ZLthEISywKJ8en8ZxiUOqvnPM1zRCbMkIMe+NYCHKX
uDxkcFMdMGzZdJyMpvb700hffpiM1avLi2JF8um9eksaS9LAKa7B/UpKQ0MQfqDZ
wY6ZPwkokAl2iyJgQRJjfDOEYuBATmi/92rhD9mCcQ+qim4jBTglhlWZlyjb5MO3
xWikZ38dXdKD2iE4bOoQdfQB08PYsqNW1QuhjdthDqsb3h5lC/zsNe0UURrvhQjw
grnMUERC5VW1Q6w82F9TZvQ6K9CcX+6gWird1sGLV9NI4TNF0Y8OjDBwsiMBL3Hu
xPtHW+DUJu/3AW0K2Dybi7G77y+WZkJUFC1hD73RLoKN081lI0Rnx3/iCq4DCrOT
mvGACmYyJ1iWPV8CDFosG9DLsf0lKDixmUpSgh/73fM4zP4pWIjAxCBneuvCe6+r
7IMq6+wwtU7oyCOkFj6n0b+ACSrYey+9pMPb69YddUla9oyoKrRWIBT1lTLyFWWm
lfXbh9qw5xnBqDt8Uw4D1ptMwDAfANXyHwepRZhcj8H2KRmWxM9o2kn3pqQDRrWw
gHIohM29e/BwS2mHpl4nbeL0OQBQqStSPa7hm1eLyMqmmpEFrVeFiA41Lyj/u/sj
CKcCP0MWCo29QyizsRMJ+u9MU6xX0cMt+C2aOG0GRRTsdVVw+c8HnZKmz1ngkZoz
RJ04UPP3qtMXHA7B9MdzmXCqAfTYLN5OsotC6xl1pQ4OodKaL3jIPk4PdISvTN6u
RRT/zxRDbTFDCFmDHC6Iz09BXAagVVSNvVw5/aeirq8HJSBuD8ol7ESRR6h5g94V
OiR5XVPeFHsxpj1896NkyFWwppTPlzKmwnGj6Kt+bcsN4rnQ8A1hVDOJCTCz3G7M
wRWF/M+05mjr+Mfif0qAn/YqOh1NbHzDG1tC+yIg3USHExE/u2cU7EylMO5/B2Oo
mkH9T6BGxntZJoov5v9kDN+prTRnRgNalQCuMSojmtlsH/zHmxYFXCUCxfqkLCuh
1stxkaFelXhj6aQLgpBYqiZM/Kz+L+r5eBce5cbO1vnfbSQ5H6K9wa5GKPTLIC5A
a3k3RoKudojBqpIliAEPT/349CUOx+iKAZ6CBYlZMgbdazP0iHX2XJHDvWGVyspl
Wqpql/v2I4NfYxlt9jROp0H5nu8u2CdN34K+zOh/d3oxF80dses2xKvTUiu4x044
eD3OFJHVLA++WGL6MXEQ7f9vEWsHe5SC1Yt88+PsO1GokTKNngNDkrTO9UlfSdS7
AFuRwupS++WJpqd/tbPsU8wJIRnV6m60Pe8KCdiTHewYuidJrS56WbBXJe6SD/BI
Cv1RRyvs4Q86YinMdCPmG67DVqairncFnyMU4oBR+GER9yn0uX1utVHU5Vr2tCVS
gJwTaK8mCmDmJRiInC2mfq3v2PWIiJBJE/Vpyd5m8qsg6Z+i7Ne/6zSZSpNNWKJQ
27f5aPGE3HVQ0dDRo5wwI3blW5VQ051TxUy5jIp6KxgtI4hIPmbwt0HoAGuklBeo
K+gSiZ2KXUCO76b/PfNFK379v9p+4iCY42tkQsaIJ0NzWuFwUqZ1HsJeib8jddiN
2/anrNb6Kp1sclgnB6BNOT1dAm2VhkFE+6CkCxzW8Qnu5MEr7NkFVPzPk7ChIF56
1UCH4dsNHS2rveNSQpFqHfXf0CWwGn8C7aosSQGdlbKgA0WCf/cGx766Y4/WaTdm
2TJVrzuiUzSAMO0Hop/1FXZu/IY8q0s2auHf4LZfG3bzf9qXZpsC61q4eR/DKvEv
4JLW+8ozEeGkxMKMWmbu1jRgucK11tCSjQqtO4hAODhuk/iSrWqKojsUIxLWvlyx
nmTWUKxivBSXS3MRqiWfOI43R7RP6VqKFfI5cm3lHsVJz2YPAzd608nSPGo66qrg
BO5aAZkIhvLLGgaLfN3ze7bHLqGYDQncdGLDzKyR363DdwxePg4F2LlkEhYRK88j
On9/8ipaHhXD2w0aXz/GlyVv6U14ygS6p3D81+hnjN1ZK0WYfqdr6mnfJlqJH7BV
32+iRA75060NeNtIE/15Lm3Wex7YAkSwZDycsmIGh0lDjU5HAOBnMURzCyTAAmJi
Pjf1PH02V2w2T+dzEJu3BDm6jW0IhIIk4ZI7/7kdUhOPVE1LBkM9LPKRBKbW1Fmu
0Ya+viqdET+SYwaxG2jscRJ7nDiolCfxiQXa+wmwmIcCBBxWBRX2o6oLnBi3r7Ba
GE25bUbjuZefi2VrZDDcZwQGj4cvsrjIy1M68l60tspnuj4G2vRh6VxrGXU4jo5T
wjiAgJvQFYnwYVA7pFuafgzQaI0QxW9a4bb8p1BNMwdXBoc07Zyx49aDh1Vazu9f
Z4QyjbvR+xaWSRUQ3RB+ygvN51NB0Lwra7oSj22ykdbK1RD4OvNKPVPDlRX2X8Sm
NXN+2lR9uvSbwuGkWjmp9RzaAoc9cc8423h4mBNANPEbofnB8Z4lAWsbAwcIGSIj
TIFJuf4lyNOfZJeI0Qd7kzc/xAL3odbfdBQOnv0bleHpkzegoynMRC6XVzF0UWct
rEQ0o+4UV4GFDEG6ar1FhGAck/ti2+G4iV51IqaThh7Dfizq9Jz/EFmt2/FzfPKD
PCvoD/k18fVpoggPM4k0/IddVzWd6B1Zjj5X6je2dSP4uSsSOkA+HspMJHouR0Ee
qjn/6MF56+WwNNFZzJmKmfYSLT3RNuxIvcc5DnOmM3V/DpioZ9WSo7OC/bX84XhB
HKPWt8buVl9zyRxhOBBNbNSAcOM5geIdxcySEke3P1R+SJfPtKpA6iyJKkqhk2UI
vagDYoRDFhEQkbkDIYrrEPjtP12DlPzkxlsgjucqZOEH/Jtw9bDPVaNoOBM87EiO
TRXckasjfly4y22U2QHFkY5Zwwj73OP0LCAF/f1KlgyKj2ULK+E0RHGJ2DSEnqBj
RFiDVA0sup0aBuC+ozqIuSK3g1gkbQ9dyJZUuEi0wZWI8TIcY3ibTgxiZcmIPv+Y
3doaeSqwK1t4QnL/p49BvDlolGJYrmBAg29H7TKBP59ZJAk0aExRsL6qB7H8vvSK
4Hwn3vClD7vF6UHdiaR0C15OcGBDgLUoyOwVQzRYKDTguJE6qqhE0uXA2W7ymDSg
rfwXijr+qOkXMw5TCDWy7RKO0hXT7fD3w99EjCTG6f0DXqtBajoiYDONKvrl02/k
t9r9kMNgYUHkn/Sts2ErEhvJ7M89pGDR40hHojXIaa1oK8QKAhF59t8TNQ5NEPfJ
jU8Rt4REw0hK5zFINqdOmYfu0Dr9HPCPNQQGxV+nQcRJS3n6QxDstOTWemF+8PI4
0fcwDPsw+1KqLS3PIT7VwgJI/XLQBNGuuH8Gfhvzht4BDpW6HacKKjrcBJy2KnLN
v1vt/kzct4NK5p+kEXbckV+KsJQvhPHQ//fF43HyKtW9d5nbgs+C1fI5ZdXF6zl6
qK+MibGqrNV4qro6EFbxyRdWMKa3C2a4YumG2/5A4s0B5LNUPitZbiPFnNwzLwqm
r+hprgT3iZs5nUqoJe9l5Zcr6UnBLPClDn2fRRRncZ2zxDoifzL+S/BYtDsT6lK4
Yg51XUSKXHTaAGQitg2hzFRNKq0Wp5WaHJriUwJBCO6yStlwzl0WMktbCwipUe8z
WZWnw3JBVfPuHdMmW8LQ2tmI4peQnrwdRrR8Zxx32PcfJuTudW2UouWSwIswPlDu
Ml4enaxPSVwuFc86jlVjSHg3y2sgfCQsiHsiOLMoI0OcVBUQgLNzZFxeo+gPmyXh
FTZY8J2G9qAghIQwT9L82JwB7BHXjJ8dLZj3rLy/uOq8IbVS5ZTrUGhiOKj4KGHh
u9piO6sM6zuCFNDNvTE1mshQYt7jwfz/lMlrjl1tNBOqilOZa6iqMSS70ywdEve2
4CC3dTFhooEH+JDwkDudihKUca/65bAoVPmgLUqGfn/mU/0B8dq9mLL/UvIAZ050
/cgk2Mp2wJuJKuPM0VLtcL06CwSAmjfJyrVQdHOB4o6BBSfqbNBB41i0mtFjza0e
9fX8P9eqJ2Z2SObib0ijHWyiOMDgoIuoMizVH1hRbN4mwF8LVDbiY292eRWNnMGU
i+06AWnbP1pE0pBX9pxm3w==
`protect END_PROTECTED
