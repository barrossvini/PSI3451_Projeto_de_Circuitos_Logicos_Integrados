`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KLJh6tA/BxBythVq1QsE1Y5fiJUI5Wp5d5pH8dNOq6Qi7SdM6EOBPzht6HuOMQ86
TjPktbWmCPkKeAjJbiogXpaqOh2uo2jnKgvj2+7UevdUq0/RX1DHqxNdQ59TxG3p
OB8hdOoZtSsA/1R6k8vlHuvv4Me9MwQaeKENQ/LCPGK5B7xTm3ZZ48YaiAfgbirX
uSlASuIsQU/cplX7rvqcxaAxIHd1LM9Tjp9QdVrw9e2ctekYdyc/eKmQaT8ZB5vx
+mXpPJRtje8IF9OvYuYgOp0xQ2UvgpqPGHhAh0/zzFQZDE4YyUrMagava76bBV6E
1tgNXuDYXDTejfD9P0zC51Sz/JTMV6dBoZcvYeq/Xltk+w7oM0EsQLS5+lYOqzQg
VekEa9NCAnuF0qfEF4pIIVKOdDN6ohFHxKTzqQkNRthtBM035qcttT80+d55VwtJ
0rQwhg/rU+4vwnAPXxd5yUcEDzSYDNfjpL7oTHzOX2YGv+tBoy0+RCRTiwYNt+8r
XgXpAWY6Z50oYrXBSbal+d5cAxES43d89WEnhVKrlD8BWBQN+xYesU7rr4TQpBF3
uARzVTzqys7R6+Iv6W2HCf1my6lXCbrA5mUfkbX9vycHK5NtnRjp6M70nFLJJXix
81NzMxXaLemywykqRiALPvqveFR+aX5kYqInEhUE4MKZk3qBMhl1uE7AzxbnC/w1
SwtaRvMVziwgASpHtAMgT0C3f/KwLrC0P+0kxlLn6TcnEYQaCMQcZkecWDoma2Dy
3laM6fn9iSwVNWnT0YHCEzYkcywS8AgFekoyyNxiDaxHC1vuqhI5K45ooF7pFd1J
aFBTvHao3kIOjw+gg5o8A0Axah/8DzSqDKXh+OmpmauGJyUYrZXgacbNWOGfcuZu
JtHmqhjU4BFdLhsrMLei8WkrTai9r09JuvN5n2jbXJ7g2Q90HpZgxmey9aoJDRZa
PwIDVOq6DtD2BG3+YYhp4Mm9hZTnrhOBd2X+t1lw2Cs4HlVYU/BX1EmrIbosxCo3
HUI+5rDmRmL1MVxSAqVfQtPhfZhSy/tfWQKwQHex7Og3QATuMrpQcZQBY2FKs4f2
t6HMk0IF1cUAUgaNmHszA2qtxgQe2AHdLk/I5YsD1/ZWRume6zXZpywfOkh96O8j
Xly05959YycbTXdvklSBafq9mFfsXjWzJ1WvVNdyXGoYeufBn2qTv7RNcraK8Mr0
Mi1AP8/8WlugFV456LrPxTTsEXYEBMVkRaY89fup/WECPm1Z/CxGcvkIVjKBMbxq
qC2Qn3aayV6dWD4Eib3TIuif7/Bo2l8RXbkcCI1+WKucjWo6qA7I203YRIVGxUzE
Rww/CEP/suaKoIdgPAheV1VrRHFfYEExk0MfrQVuniqV49+h9mPv9IfsDc+FGzMe
C1Fo4y2dmtI419VaS8JtoFeuraKzNiZVHxUIUe8lRIhYF8b5yowQF/2hn94yk3QL
OuaEeWaHcAbs0+dYuYfjXm0T1XRRxmABEMW3fVjwRP3dyuBSPiFEis6yoe6Ll74i
5iV+hr/ch2k+Hzs/wYwvFiTfLLpSBLHE8OaP1oL8bU33k4/0u2p7V2L3nVicbFUZ
babdBc84a3CPX9akU6FStUc5XulnPAOyBsddjpi+Fh3KWoCCMWOGX08+mCs0/gCA
2V/sm1GmdVJq5tYd3feWvfRPGtlqSfn6MLjqi8UwSqeU2v0+SJgLM3vxjbzh9oiu
PL2ofdGkq8DWUYCgjbrC56M5KukOmLkJ7G0t15NlQlsq+LwoeqBFLNUlm9HOmSYd
yeNZ31mnuz5m5ynb2YeEY4rkWmiOE+3Jlnsgecl13GRiEXM/vrgWbOa/lsfNHu/q
tOUpGAhoWD7VsdPrvwAU0rQwhqVcnE2Zldl+U4n74sHdALajw+X2GRdJ4mgC+qsb
1fGK4qfS0FA5VxV2QvC1nGRrg3KnBbAWgxH4qUBaKpazlAGtYO5qstLOTqGnoQJJ
C50GyKc4bUT/8mvu+KLNtvbov2MKw7aYsrsfH2gIACwez9IlDTlTBFLlQICT6uZn
mN9UR4vhxgzrJjZWHaKcnRGUgBGt6iK0Jt3RVKF8c5CRCL1BgocfZ9aMr3GEs4gN
G2n3PkPLRMnTynysO3Npu9Bi5qFd4BYHVuMgK6sjhcOVgC/7VDTN+1dKc2Y/HUJ5
G3JWDqAybFRZ6OcooZda6kXumBrBVBJ/Zl9zIbiHFHi0xfyf0i0o4orha3G5tB3k
MGE7HB6MSH5BWC7pr9qKyrALe4Y2N7oHGDbec9dTKBTA1/Mota+dtLtNcgg/DSMb
N0r+NQVUJr0a8tZ+qPqhFoEIcxsciXyt+bbo7n2LY37gn2yuyxvudrJcmJDgrIVZ
RCj+jyFbnPO3bB3iLim+NUqALiZ8DEmHLJplRNbvkJ4zU1E3vZsatRmAlQXVedOR
NwaYT1eCPId6pVRLKZ3pK/t8HqKv18TUkXhz7xGhLVJfkIRR4a6Al2MUl3tvDSGI
Ihzc3X6awT1PdJU9nhde5+3KEZislIpvXu8ReEeW4GDrsgm8WhXmUvcVurVyeqvm
DhwLGGuZizDkZS4kgRPbO3P6TIN2CYTpZUSNvehYAxpSMNW/tcLnVY+bbEG/KEiR
cqO8MrJT/oFiAKh6tn+4d2O3b668iub44lrql0D16AZusDuvV3o5BNVxr/gQ1j4B
vCw2uk1rAdz+VgdrZYTLVFKC2CjC9dDEwW/LS9YrcD0IlN6NrDP5UBiMCb40WLS1
droLV0vVoe0ieaxD8hrmKY1KVOa2qYjZ1pVqhyJPA2NI0L9qrlIqzk7dGV02a1cq
gG2f5hOhthorLLYr+SMBc9K6tueDmpjHT/AMwzMV577Kj031j4srNovyxp9bTiTV
+6Tx1toxIN6iV4B9gTzIh3UxUj9VxEKkysolgaUrdwGqmQ1o+CJF0z4bq4qscQ1k
F4mbK0v5OUUGoThsXIev1Fx1zIT69DJxrdY792SonMJu+vELts2rw/qHBiK4R1BL
UnHAKaxT2aYqjbHWOU3NT0jxrg9KvrYNqqhtMPzeDTd+PLNiIWop+rrkjPXDeX0/
3IomQTvV0p6IcJwvofPsOu6ENSQhm+D/8j/p3tETgxFA0ZHwI7sqO05CcyT3O0TP
ImRGPjXyjb54yXo5eF1cCct4z4sgaRnSuStOKB5Z7Al1tCgIAFi2BDCRpR7K0WNc
IOJkQr93qUnHZrIZbh4PHovCHY7hKYrmz8VnrzQS+Ti4k1u+1reEHNW5fGUtpY6F
4j0joFLS3AaEOnweqLcqddnURn7jN6/ppbcgpVKYO2UppcvdLMwmnmgdPZe/Gte3
WcUwApPPMzc14O+zQKgACWP5H0n9eeoYzgNzH6oLl8rTYSK/MkFCEz25YP3gj8lT
o/s0cDOttAgIwxRP6RsSMK+GCDqEB1CKdIXWl3coqpcXpwcfleXYFhl0Dnigpdmn
bYRoz66NBrk/pKOOjd24r60S/1KbcaFvPRaHiVMc75+CQJqDq3OeCNzhyZSNMqTT
J8ztHb7L6d78I6caGPvRtLr9BjhpgLmVtPLj+bSJ8aTxSDuwaGYWQBB6Fjx3dbS/
R4CULr2eGxgwbFJ31122mI7tEyH7TTbnsZYgXIxXOAv5b9Jh0Df5xF+HZ7k24fzX
Kn8xEWJUFBiyaCtb3waIsursZ+RASLwBKu5XMYUPk7qRJjvfGWOwyS63IeoekVvw
SY73eoi9+wffKGY76iuMOgLhZL993i0BC3mvbpgyPPEC+eO3hPs9eN3nDAgv70rr
hyJ8jOoAAaPayW2ADW/UUwAHDo30hWslVJeBvvte8KZfrQZQJiK0IXPBucDLxX68
VF46ESG6sg91d6jQISDj/Nx5/te7cmkaNd+aAzXRzivWUAxfsgT/f6pOomKzHwVU
MforYdb+XgCiG7MYZ++d88GnelgljCmTiDFHn3xAvxeyLpKAKkOPcN0TzgapvYC9
d43pTjiHKj8GsRuON+cNj4nWSG43dSvfmTaILu3eTGNTHrPGAdn6GGWpoBsigFcZ
4X68reqP5Jilw1Y5bAXPqv2N9gt4OcNGvdryFj6TAIR+ODJwXSPlt/p/2fbScyan
ijEg8S+jYkbbBoTsonGA5l8ifRg1lvlIgbfFCOJgQPMgGZP66Gpk8QhWdJU/C2Az
jIkKXoz2pp5iDH/WaqlhSrUQ2XxgK+ssJUOqMqEAjJlQM0lBlyfhdLxEkIhWLiPY
7D+V22NJwpyBcMCg62Jqw/QhTNdMG82KtiKtCYvxPCVjY9mJm1V0zuPf85HyCoCG
z2avA4CDXF2Ai4bdgaQYp5CiP4W9fKtGHK5A3wd9oKXlFNJe9oDjoZa8yZTe0iJL
Ueqihb1cxRM2FA+QEtl8SazGwCiTCJnoYw3AzC/bm67IcOAxv8GXOKAQvcA8B7Xc
t/QXL7KIWi7mlsFYy56BDlt7eH3FCD2l6OMEjlnCO/fcRnmBulxorwzsZFO/d4b4
plcUnAql6lELXUCWa0HxmCPmAi/QX0xkbi0IQhT+am7mlcxf5mBpjmuUIeCO870G
xl5E2aXEE2xiV7JLN+nk1KzaZOy0TtDU2Ax72KHl3BFV0ubl5M+zp0SrIyrjNV1M
7KapNoIsm2TVhhi76oBGsBzqVZhEmjNqV9aoArOCQY8jGOWp+Q77GE51VGHEWyg0
7i4G4q2iv1sFEk4gIC6DQKI5EVish/zMMzbdRg1AHbhV5W3VjL0Z2qcQwIQrr0oe
HqQYjTGj/hecRqwG0S7HfpSLW8I0fI7qjgq9PtOvd/huB3cB5g7T8eiKvCoskkDb
0x2H3ebljOBcnrbpNofU/ydAl2HNWWHYaiV9HPugCMwndLKewgIm3pIpVG8WgdY0
KgfzGAPwX1b75ufgecMYR9IMia209zcWNCoMLoKd8QatTPZKmoioRR7DKJw1jobY
Wfk+OG893FrEk6iG0XNSHLdrleiLiTcGSR17dz4Vs2eqIr3/xHMNsIcyvebiJjs4
FK719UMXX4wQGrzMRLDBy0y88X5WOskArNLI/4cFHzfLUVVKzaWiIHJgAx6ZBaoQ
+Efj88Du7e44G7n0wq4S1ACIGtGkdNs1x333o3jgYD4uNAKRLmF61csuf311RySC
BP1wTiJHv5af7Q2XMP2rhM3JHH/P7XQ8Rw87kPW481hVXGa9C2qspEo6loEown0r
dm99lnm0VFcivYOJmRHqIvnRdfyggbk0hT4R2CrIa3iouCUHe/ibiunt1gFYVYbQ
epGO/BuQ+WPD5DKvYXiqjkN4nHK+Shfkc3ioqGd4AJypt+mcxkt71wxYV4LWPdwg
/uI22w5VITo4+9s7d+XNsAFL14coAg0HyYeK+ozN9WG25E1rLHRi8FQqJQEainzS
61EHqMNUYMoMARS0cjyMtYjEpEKVvBUhaISldFUwcudr+2leDS43ERR3N42VIvJf
iaq8ZhbC9dREj7DqRmkEjCNXiqSaqO4+bVdnCE8Uhx0OSMlB/oHHOe8lSKEiVfBl
CG33NvrSlSP/mnfukVWfYchhvrzkb7aJdk6JE2FSJx3gyEg/sPESQFSYtV1hn5m2
MIdaQxv+stQWQfcXFHj6EiVPjnTCYn3CxWnO6Xx/ZNM2nqvQmKRbHdZRU2cKz/PB
cq/OSveF0PetRhNQRJCSX1oL1/8YjtjzqRdNA4W2y03EVeemJQ02VXTgl+eJi5l2
PnKAyZ8LRypn4hA43SXjKUk+5BnyjjpPRGq+8lF+NcJnp0vklWIKO9VcY+mlVItT
GtgsP6ICK6ZEInh6r6RrQHhKBXEqSH5nQH3e0ON/069FFSv3+5AkZ4Gv0IDwOlXN
L/IgjSa3xp8DoFRND0lNiQwIESbyEqEjAlKkS2TlmyVFlBScDRG2lDtDU6II/bv0
GH5OtQMG3mlLVerS7V0Z1NywlV2cnU4O/PFH2TkbsV5n1d+uZAPd5hSlsTa+Q0jD
TZZhmYE6f0ZMsdPsMGMhx6v30R7DEaWUG73t1DkYrVr+aOGRPtkCtfOYSjFBzLb8
elFLKHt/+GYHrFwBHnvEtMClKRQ885IDiBPuWCjY97DRFqx1zALUKhviAvS9sqeN
TvKQC26WmNRFURo+aZv3tmruuGzNHNds+vIlrORXwhUDA6KDTk6MyXEGdQ1W/FBt
PZfGW0UOrL0V4LI2dgz/XPc3CmXFgGy3KybUwVy4NFsFJxqeoDT5xIDFQXIZpNyD
fzEvcC8PXbmfXFmGk93PD/i1D4ox2aK6Vt84h2Sp8Nc/qkvzodX1BOqXw0rQgKXf
AOTeM8eQkHyKy6pqz1rLdV0Yfr7b3DgyESZueNy/aKNFMgvyHW4oxW//eC4AQNoQ
3BgCjEmx/l8keMKcQc1947IOC2PPp8ZxBcIrn8+c9xItYPB8mtpUs/Jy1nOkM3DT
qBIxDDD65a51vFdQZLWx0UaeBd6ztKj2k1yy/S1g7274jjkS5JlV+KCx2p0+nmmY
+F+PplMPgSg5yEKya15wuiUuRe7SK/SwZ12ybnrvFpsn3z1AsQrIMFiJbnU26lYi
n9zAkIuQP5Va2n35pivW45WmxQuTwLGULvPiMhpMEZw1WCY19vp7G8PQ0Ise6n3G
2Stt5CtW1wpY1WvYh+1NyUYq/ttVT7nMPrmrkNMrjX0sfwc/+XbSDEzmFrdXtqEa
Fb+mKH0gP0CadG0faRS50c6nrowkhFtOsi1gAqac459L/WaAVlhVmOqphSVM2uks
PIyoIBIMgvulYq4pfpOzT4tDQr0EqJvGbjjLVsDdSZgcg3q+Mn9Qoc6L+SQk6g84
aAyfcv1quqTiobMzK6H3e8wGZ/BWfWrBiZnyCIwRDklBCywlnlI/xx6fsOL6t2Ff
IFjwuE0ITGg2hdhBJ6OQ+hnMW2ACJY122z66W9epVPzBaLJrNOaKQUy5BBpQMV7Y
ySdJY7XdljAis1RSyfT/OwuyYp9uIVvw2FzVXxVYctybGWqF9mOCaqBQTUHXC8on
yIxMuYZPBVKwQ376zaHZlqUIe0PWGnHkZ8Jelp9m6T953oHDLYoB3+/9xlfhWyvk
JxpHAvW18Y5Gr/jXg6fh++LFA3IVAE/n/NGgXzHEQfd7+WBYur/RrHyPf6HU4dn/
19/k9lfb6a8QFhdv7Z4/Wn9CbZrd/Ic9CsycwHgoB1nOujOe8HWdUKHSohg/M6ln
A8a5nCLb63VN2G0NeA+sTiNMyIwiU2HOh2V9yLVPoyIxWqErQk39+VO7Tm8nqtDc
DynQvcSitZ6xrYmOSa4hD1KI0q6OZhKriLPCYKlujcTs/DToGTiAVt8eAAcvW/NQ
cZXj9TN752+jrNDK0BOcARau51WN45AB2T6wRE9w4fR7jwDAHgTWHIuP8/czeyna
8JZyJL9Im4F05T3RIr2PaPGuafDE5lYXcgvlw5BfxKtwCp0ij5eRRpoq3NaSqveq
5bqNv5Mf6W41rOHvYqybndtiCS2+hLUJ3TKhIkBqp2GmsgoljIpm1eI6ZqFJqjMJ
Uqx7ZvoT+gncvOGxqGZvhGTrzxJsUFO9nvbRd7sSJ61OBj2284NUWWzO67cAGLQ3
DrYcqa68JmTPMALqBd8qVUHTltDjFbBESzpzNnPa2x88B15agUcNviyvDS4rqu+T
pImi8t4GLClQ0sY5URdwgmM+r2FLR6PluSvlZ4YupxXCclDJRQFw2zpkprwjsk91
2pPJ65pxJR+cOdOgC5WF3HNrgtwDHbFP3YlM2PqAxr+XMqRJTgAwtzDUmb9ltNzU
YfYinSA9qmVgsbr9kH0DyBoUR2Xc4pjpyxdF1QesVaD3IDmQaIDq2n1GzoGEqkek
P7TcNwGzcM75BCXP/pbbsaQpuackG/cy/qgyyBUfuuEm9vH0Cgdfp7+areweun/Z
ekADLdMuJbVudNWzS3fRKEJWr2airef3xIzthZVpUUTTe5ThvNNAWo+c6k3j/7lw
n8jOKQedVDzXQeY0dofjt1D5cNOy5saU8bMUYJDb27PA+vmqcN1Lz9MCI12YuH8e
k9ZCpHXCnyKvPcKYiVrIyOxVgX5Snk6uhKTzmi8ucO0MuuUAnNYYizpcdIORzACz
+RMlLbbo+4+TJ3vcD7xWpipXJ1A6724y8tztN/TSMTU0/L0JqQu4glm+VlUQGlzD
SB2xEznjkKlJnrk+Obqng+XlCPjG3KhVqCWoRjhNb4+7VrtIBISYuaLfevfWbw1Q
ZboQLyAP4DyP6VnGXl9uHK5YLpr7QVKE0U9neNvJyx90ERltCHX+jO2YLnjfzSqP
y5zICkRoHj3AoB5027OaJ1IapEWUZQ8UCvXf9IrYi6cmReeFmi2nVvBbZNHV+lND
3UgoG9PC0J+yyvmehRZSKLZx3/Yh8ZnMgtL11+B2NE2+u2G/JrbdfbxCpNgPrt0D
X2aJxMnmuze0hgXj4I18ristkinEZd2rlEQ4iMbKS0FJAC+S67V9Jhjgy5Q2JHbX
oyGNakBi4VwyUdrjdgiZqEtDG7IiWwzOmixSFvzN8FnD+2GU5xXTGQDIm28xzNBp
E/uqZo7WZslXzK36Rv/ILVOaVcI6xJV41uZHqpor81avj/Rpqw6tlhcaXecZ59zn
716oFC+2ypK9FjZbAUNBfqQqGs0cTawM2jDwoiqVDOkJzXfnAvMM/wRK8ihQFoYV
Czw6XRz1/qpQaGehp/X4XQYX90KY2yAye1P/k5zG3rvqKJ5cM5ljZdNGBqFulLru
1pHKOPUSo1pZSuZxQH48nkX6fenney8+4WJ8yVMx2V5GtPEbr6cP0qCTeoKGKLDz
U/U76kAoTiIdhPorTk4Bn23OK/g9CRNVBzNra3GXVXHKAbzEcrlbw6BNSxVOiXfH
7A9tcbJ6KEkeGyyxBzBPPgkuUYbYbYiKhKhrvTgmt4PNcrUxy+ufkthwPRnw3G/F
Xy7bvBwh1YSseNV4aM13kc/IIUOtIQRCxM1xoY8xEHPTjX7Uo5/0UlIQT54LaUe1
mYAiTOHoGJfdutedsXtLQyElgVvUCCWigAi0v5CiLUfvgFxAxbABtfn8In9ydiPG
eeGCJ38wyjn1DSnARMDEdi3hZCZk3L9fZc70/5wuiuqNPGHB6If9jiyuuXroWSgI
QSAS/EX1Ao2a4IAe1gHfphDt3e5Nt/iKtUwovTTltHJ4K5YYgERYcCtC1W0KPbC6
e70SfLBnW9BJyC3p5rLUbH+sIrSh8TLc+fDeugamsV2vA04IyPrwqn3Q2R5T9x6Y
wHxUSDa6W+grmxqRWWEtnMGgQWZhUHDu4SixTWy67kP+5XEkjGI8oFduVHvcphIg
SdF3mjzbEVCeY9Z02B4ChYJCQIRKnp8jqzt0+5rlNgnXyzEOI9AEk66Dmab3uYmJ
e4KSnX8fwEdh+Vqn1bO+yPSh6/SH7AB6mFPwHeL8lWk6jcq14WnkcyRs4F+movyQ
iWJNGp6glfYtVHfP0vRxRDByuizm2ut+H5kY0g/iBeToejRlj6ZeYUaYII6ccR2H
qRGJ/+hmEaj69+sZU4zYuBW4wQjZNBf15GKtiXTq6GMg6Oo+//sNmnAe87gjhmQa
nXIxybZsCVAriFP3zff4xPubL+xNO49HscLa0Namn2zhxYUDsvXQ6oL8+Nlui0U6
orT0b5p81v106UOmC0oAYU/k5mQLeK/TAiaCBxmfeVGeFVIaolTJzPkGjqZQqOdv
Fq7JDrhyHhio/Bh36sfVN/hg1/FtMhLKm+qdQNwrl6G+bdxIT2SqbWuhc2WooW0U
CIZrWYJkG//HXZRFO8rfJqO/cIjcc+NLoPPlCOc3qOilm/kSR9oBw6sZ6bSJnlXl
dbGlQE6H8TvEXixFM0LNxxVoYbD9Px0fwFmhDGVy0HmPJz8NWxA7obYethhiFMf4
sjZkX1foDbzHCR6N9KkQiV51B8866OaDNGLNzZAs6kMzNuwqOyB8Lu4JZIKJllDR
oTyUdictbEXvkxvtJvNuW7XYEpHj0ZecHf/XQMugQ9k2pBVSxnp4WoLXNPSPkOdy
adXE7RMoqQx+YZnb+LlHs+JprkieKaWgQXAs/pper85+lv+Czr9k7+Ux+OiCLUip
S5dC5amGPJ4KI32P+pWjK01G2BkugVdoLls3JJTJgPOh9xEIaXrpGvO64AXFacxd
CVLrrs3ZMjXBYVAF7I/c1xEDIZ/WxRaD/F58cfNYWlt9jgCli7XayW6/ez2SY/RI
4xgR73sl68g8FdiYwgPvtkKwmY4U4eS6oNAdyzf3iMNf5on/1NEHaWXNu3b8HXWw
kud1QKnLPoCOXwLLXJNPF7XwrjUMHvLvBnxO81ff95jq8syNsXuzyr4jByLzNadT
kTRoDTVxihTU2ChWF6WNwbeQEDaS4LooLXB44gHEtQF6cqVL9Tpxg32i9qME65C3
z4xibNdc/WHP2yX4s5gl+ijW2KE6ddUvRvvDwCV+A7Jf1Q0vfIKlGEtpxiTHdLdi
v93z0I6p1wptytxK6MhcjipxKTaLiDYDwB6FUDg7tYjteExwPOtGeIuYUGL1Z+lY
iYYiV4ALQ+JZCI25nMpfuXJXSpN/ZVVJ9iXoIv0kLmqGMrpRr0hZXXDnzNJv0jnl
QSOmjDWeJ8e6b2GgYi/46XxymxP1ll9XAP2DZjY5IVnR+hdWvbRoNLDl8LHPVpVg
mVChQBESSlNjGoGufPDCt3usjkUWFyuKq+UedNWByRzT23kmGU2jb4vR8pSA7hY+
64IooSVaI6NtsTrbxnd3oX8uzRs5CAdr3GB37C8/PkzLTm/1GjN1u4/JubRlCSwS
xZ1NWFzAIGDJ2r6tqlgjYLJy+yGtEen6Xm3+b1PHpa29unjnhUmItH7U0r6aBqcd
ztpX8bOYpzIqQZUTB3S4ernCac+8UlXdM38Iggtn23kuBat637HYG5sVHJBN022A
`protect END_PROTECTED
