`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZlRVvq1FYr7LGSJHcWHkuFxjgpHg9rnCHvKFnJXAjYmIvVYlLxBz+F7LIDbrtX10
WuEe5cJ36twzCnwCUEP7+lGT/e2mO/WjJ83j6JAMvCnm2ggiUmO4tRCtLi+wnpDB
XvCJaashRk4Rp1stb7N6OmWoZQJB3euZDR27DpXDKN/4u+3aXeXHsM+GkY67vdkC
8zzWD6hkH/wkO06O3F/ciHuLy8605dbMjQ56cENTM2jKsddJd4CX2pq++8RFgQ+p
v4P95AvSUHxts5GwhH7z82E+Tvbx8bNCGr0qs/BT9J/MmqO99uN3t8613MyknKsA
9IrimL0Ogs8ikffrKeddJazPxyqIbeNR6sKtGy7WchIrD+Q1hdmHtfoG76k3C16D
BLXQZH325RcbPiSISKyjouf+kLXahlp0japDCqPAuC2WBSzyfnYYNpFqcs5FDKu5
qz9Tb4aj8Ha+hn+vomNdB9nADh8BxvPcZ19KrlAgDw/NlSYxkI6/LGUyeVNr4UCf
basIxOnU0bEsqOQVNoXxj6GOjl8PPbhSgMwsX+QnGurrc68rMPn80I9n98rMmrQU
zv6zjsEM2Kp1f8VdtcvN9oe2eivc1Hm65SsuYScP7ssIisS0lqJJ9C9vMQSSx7SH
zcykzHJn9vWKQNWEFOS90sUgvaObmbVkn4zvS5+sn6LcoPbWrc8dwWbaIzIV4d1L
2/nCU7yOzoP09G0Q/F59uOX1zB+UjNs0ko31uWrO/Oep5ZscsQ7J6C53dH+ge/PH
UAcp2gY66Dmd+bPihihAY/SSUybZvE4COz5X7hlOm6dfMRKFQEsYHUWpABEVs6dM
bsiS+jxJjrYGCeBmL1IeDMsE/lAirZgxq1Oau1NLTFvDZP+Pn3VcYxf9Ej10F4Ge
13gWWqX4Ok6XR7mvCR63zPqMAUo3jIydzj0l+ysJjzBc8oQHIxJzndy6b8GCn2PR
WIcV+fVsheQGGzIF3kQChx30p2xh/aLvgMWPDoaO1MKfVkZvVKhijZX+d2C/qfND
bH1BZBjwo9+rMo1yUW+dGh68PY9q1li0fPYbu5Kveu4ykQePBf6L8HtD8mRI5W6a
wDxbcHTrldj14flZ/4BicRXTbk0bUMl1FMgyZQrsziQdRG0OZREyaC/SERCP2n45
XcbLOJGDaNIXfLTr0m2hWSXVQNAf4BFQs6fsGfaduk9KyTuK0sJUFeNR8wAxXPq0
opTiuwSa0Mr6IWCDLY/2v6i+C+73WvbIuSuvOzynte2j5C1/tpWA2CKUpg4G3b37
W8eK7PPcLxJJi6pKTuC4/ZsHhs3W43Wtaf1YRvsOAzFRgvYp2Lu9fOQfuZLrtq97
UKrMGg8tBlZYECmYXbENkzw+aToVDkgZBf0gUB/ehJVu6fT9uSUR13nDLCAjRATc
N3+d4PR45SHzYNbWJPN53A/7jTFla09xx1ddR/XnXNwg7tLgP+z0rFFxGFk6IS+a
POXDyT1R2JGww3Xr3tk7vXveUJrhnudNFSeZnwy3JvSc9YjoGuY/7+5YFqf+VCeY
ZKhVJQJ+IuPCkDX8REtNqEvMGbJvXBv13w6s1dfyZjM6uf2Ssv88vB4IWe/fq1nX
atkZEZhI3oIVHFAbHIaQNzZ+Fof73NGhkRFnIMYH0u3TdeEeb4+jJvnCOjdU/qIc
Nb09tUSjUSvBgAWfiSXC62XSPWYZX4T/lqAzFP0hu6pOKXKlUycJuZIjBJiK6g5I
ZY5NZNViJOnchYCxFC2hB1DV87yuxxln3e4NzBqZZSpVQYLoKGmHqFj6oJ8nkGvE
v31LqhD7DASXJzrZ9mD0VTQ4nJA7tt9jrJq1MWfhaZklCEGyf9CfquWV6w+5TjyH
l7PrHACIzk1USe//F3zptU4jnKkFMd9woLxVt4GxQ0hTHq+I3Ka3mkg6a3er6H5M
kDvqUQOoyA6nRMu1e4pyyD6oWg1X4xBs9XUN+N1s04dKRWlrImJliZsAyEFzXzqz
yK4afhGPt4an8vTR8t9jQu5X2/Gp667w8/VkT3Gn//k8maQYPVTqBAuesA5Eh6re
hFuk+cG9FZafWVH1Eq/mVFzsbhArr1mAmld1kKacU3+vpwTtwcIq3y+37ifa01h1
lZiH4SbH3mw0lu/Uff0qFqS8hNLE1waOOrWXF2GZ8k4XBxCskFOcfhXFTk02XJ0k
efjifbNeiMe2CeWToBnF4iwMJl7oCv6pENXgWG0f1N5ncPqSroDb02iYpZE6waYC
Svi4XHfnUMLmWwLr6J8UzPfxvxlnfp1fAR0x7Lzn537q4PVaQSwrhbd6UrOyrFyZ
XEz+UeXez0hxo+VMyAlTnTVkWUi3EBrTRHVMG2WpM93ixUmIkbFO23iF3XK7ncp4
1JTXtLDPTAzlborH6OVC8CqEdzzsF7+/BzsPfE67IUsBSv3SBhHu3O6n4dMqLnUm
uRijGqsNAGtf7KXcUkQZqUVC9EE9w8y07hw6iDDNbCAN94e0dc/9DwQSZQ1ZbbSl
edOEZ6sX03u/QD2nHsaq+DQGo0JGuQoKVPfGHnpiNsTTwDWCdHQ04jcLYB4cnnnD
05ko0KIFBh+UTHyWBPIz1QS8tqRq8wg+oZ71ch6+kRW3wlvU0LCAkG69waUBH5lF
6cIeZgbwQTc7DnuAF0F7+QuJ3Y0yhym2uW2WY7uPyiPiHYNt/88GtP1PkzPAaFC2
qk+u44zQyEBiFoJBjfXKnO520w+y5UCNrQj5V6DPA4sDnS4m1XpfTF0zQwE+IzBq
1k/+rh60JXhGdmg3QMc1bp5FfeZ0ox37YCGEaIjI9wJN/OIII7l8cDPFkJNiM3Ww
R+R8e1Fw+114Qt+c2TaQA1gC8AhKyUkbRzlHNMbvzDCEQw9UfVReqadzyVG3Gt5c
pkqymRGG0ZpJd6SR7wQoqTf3Cni7Cg9/VbCN6qVbFQLcFKBjA+6nyecoHCJpROPm
91oSq6ftF7hfN4T3jjtwZ9NjtcAF8VKzNg3oo434MqKWNPt5hpaZi3lmyk3NLdGk
T+zzQLNv+VCDx6jwupnwRzDyfAFfbNLuQeTzv+kqG8c/gwsnbZw2E9e+qXFUDuvw
I0jV5EKl9EiZAoQ37tnO+Vfv1N57alaOPjO7/2HQt8sce2mZjsnpyd6rkIVZ+Lrx
1cHxBBdP2y0tokuQp/dkVcMFIZqnkNQGad/XRdDzfow0uD29L6T43sViB+bBNLvk
FkXhDuAyOneIG2tZ2oZeSSLEIZ7E4NrEFQFCBp4APXl4jYE2ZuP6mKUXf+XTgQ3J
u6PZP5uhZ5lpQdKLovTXbNPT9tmX940SVsjw5OMfOj+rQZKvFpZI7g/rTBMI3kQA
6BzxrRvJZkSMXZOHrADqN4VLpa/z0dfOoGJHRg/2jZntEqi5l8+0tXeWt/lJv19C
Egegc6OW+zlNhgzI61h2oc9BJzPy/hzdt2SYLQMRzvoqAQWHSmz3JzfOaYxK2vBE
Vd1eZdBrC+Ojw2ID5OBGMdfRr+RM/JPzf+WOM4yAplA=
`protect END_PROTECTED
