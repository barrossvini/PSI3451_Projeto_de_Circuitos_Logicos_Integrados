`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rILjP3RWg2xI608XFwr0eRB7Iy6U+bhlvXhqPRPnu8iP+5VdyWk9mF07ELkFoSE1
+1AKqXjxIBRo9iJeHMddThbAQHllalke+GmWZS+zmssb4bziHC2kadgASWkjvVTt
N36UIzyZDrXhB0s6UpJElrj3UGc9UAy+6Lu1kjUXAyYnudzrS7wQMaZnthAzDvSi
OzqxSkcOm3xQCDIlV7uzzg==
`protect END_PROTECTED
