`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/KaDO9k3BvGzJQc8zBI1IYfWy3oyx4ZbyZcbRJrnec+DL1cnboDS2AY3JwpT3GU
H1XlsxCMbYPhTYgwe0LKBJA5DEELOBVpldZxmyBi2d0Er42DyrUITyYpc3qSaRvZ
51qAzOjH+cF6Q0g2Hl6IQuw3pvIL+NYQcxJ/eSl5CgdWZudKVM+gEVQVYMfpzLgC
MuDYAJiv5QwvnG33kQ5GkVTJVsx/cUcRcxdPGprb5E6+KnfgoJboHrdSzUzcP386
WDwbCUloUsEDWbNEPqPEzG3Bz8jkRk/aNhs2fwXeNERsP0yAXyBvEe1FHKKxVx3K
xcfoHS1v847Qb/tHi0YpCrdpRJ0rDmEIvkiHyYjXcH6wCZsL20KmKy9kQn61jdL+
ZYLMt0FlBU5HVvhBvEzMcjKBFRpuu1a05Hd9XCMc3qx54jnm4yiKJrc2KcYPEC9a
uoH3ku8Rox9O0VtmJx1dKJJ/dCjG6PaDQVn1VzzDJrbxMe1/VBdTre74/9Xa6Hfq
SycXB1p0y6NWq7Hr1rs1vlm6GiwiF7sAIn5w/asSqJRdc0JD3X0E99Yr0+0lFl5A
WZoDaHwUN4uETNyaCecYlGI3d4RX0ZdkaZ/Sq8Sfs/2caEj6vvZZsXtnagznO4Cb
OwqcxGtc1YYkbjhYzi6CamYizsvnkrJgdiixsjxkDe8THhvpYA4h6RJZ3l5UGLx+
4nnXcfUXKxBPzM3hdQIqTd43pFEatKf6HOPKQJJRLcg+8H0fC/BmBS/QovXFoBDM
UJItlDTsCSw5nNcuF7SpxuB/liNkotneYImI00Q38BiANxV/t1T77GLUfxZJwJxM
q4/iyTRSGq4zz9U5eiPZitfpvbwA6MTE4upGCxEqmfXOwIC6tkfKNQazhGdu7Qwa
MXvIKxtt8Y/Xm5beFKpeoNO5HaSYJRH4SSullllnU8z04prg+tLuvQFPmPfqh3iL
kkbpMLYPh5ASD14tR1gNmQu3l5A9UhixuU97U4fWd+0jCwEY9+5I/54fUiKJ07fN
FvGJQNKeFTYT7NCcezevGIB8H+olhQSpGyKW6p30iow+92V7GqCdRHqfFfsbu3OF
sBTJVriQ9pmY7lH//8YYK4x/a27hrZ2YeWbk7jSzl6VHO8xitL6gHO4cKfAL2Oy4
YKdJUa3OBCfktqSHdNVsXstWKrIxEGX1JlYVFYqfgqps1P29RwoPdXVSHYqdGxqw
cWBN5hLrZ9Pp16q0mmAfvEeHdXOl5ngdiCZoR20ZU3gVBrihqsm3XZpF6PzMlYdr
6Zn6LUYiWGgK/cbhoK/knz9Z8grAlWrjYLAZevBGC9hPBdNwqleQzkuyn1dWNkkr
s+66SsQl/IFyH/Dg5WPWnenQEPTZdStR5Wa926OE7M91tKkaORZk/ViHHogfJnl8
WPLFwHkkiu5mlN9AOzK6c94NKR5LBPl2XaeemjUkBVgS20AvzmRm0XRtaqA788Dy
bMr2Dl/q/dwAT+0f/OSgheEOsRJZhpxPaIdD1Lxc4n/DU0J8WlIWuXw1W4A96hxr
4dnnbvCsOjH/SeJjut+lPe5vU/wbXqBDNHnIGU97G6JufFm8QkrRd/Z7TDUCV0tV
lMBNpbxvjvEJOUs+jYnoQomKGeFQSA3hJDjYXtKWT/XtIQ2CzG6EoRrLz/oYurRi
3tkz53Ob7xQQl/I1M4WsstvUjCm7iaWs9VBjbRMaBOgT7sc899thWXDKH2dT5Qtz
c3DEC9yPmDiSCEGiZXyarkCaWkXuaayL/Lx8xFF3IzJIJ+JSyUtWPi1sOOxFT1sk
maz57nXQtiLnzeKgI3/xaKmHLJTAZ94KnqVEgZcvGsj1KAPWZ13XMbYxSnD3+x3m
a2Ldsss7lnL8c/hpSZ4QhLopI2dlNacQcU96cBJ4SPPu36qKj2pokl1rkyOalpWv
YZGWQM5pfbsfdbeUL/B2AuR0f6LL9YC2uFjaL4NpJwbLVO60LaLIPiQQVP1HiMK8
qrChcptnYGgaJhbSbt5Kn0/Gm2gpJ41xkwZXe9LM3pBHfIpfbLJ5KtCUYk0ILChO
LO9pOKv/HSjSXc2lWZtLCbA9ZX5wQ3Q57pWWZLDVwIkEqbQk83VY/6tkVwWeH+kU
1Tyz7BeXYcN1kcZyzvF3u66lj2+t+VJ2SptAU68Mdi0lH5peyerMMdWDrMcmW+VK
jreg/yu8k5VnX922qVd9geh2fmivmZzV2w5FqLLUKOouHMHEKvh/0BI0ciPmEKog
AQnAbiwmvdh4KgLvQrRFW6SOos26F6QLsfScw6wraH2+uJfPl+XEp3GKLxS8XIA2
YNPcCU4vhB6yK6b32nMGG/uLXO5YRhn8oEOTqXnGtsx2g4hxQuZ7BN/bRvNwi0Y2
ktyi4b3vOGwFnf+/igPp6ykRDAlUJIl9/154Vfn5S7GZIWgwYEs6ecpcEGuMmrgI
X7YS0+Wy2sHz3x/u674PhSwrDXNr3It/kAUQe6lHfrJTB5qXQDrOk+KyHCK6sg75
mZHK2Ar90GyaxOEW5R5jFBiqsO/BD03ig6wByxUys6YCUNfPgtM2VF/WylF9Rw3l
wWWLRVGpIoL1NNFAX6GUM/k1wfjrcLFxMT3IWz3TgqGSgIDfA8IY0n/2hSEyiP6d
/uGMK3DHQkxNIPmkIRviTv1snJR/WyHvrD51MF/CsrS4b2FAdXIUmVoaUGd79qRs
AxS/cSrqwjvGO5TuQM+9VTvbOSS8ViIAoHT/sJDXkG1aTkY1LB74GGMJdkKmaHCj
cV5x3S7OaPUc8p+MrdDVCofXSZDZMzVTx8K9pGmeCiG16N07wYhp+vIZAVpVRQJZ
VIGL6pyPS1be+PgAT9F5P1wC2yxZ33fvuvnDXqkVmie2KMFocH20MgyZKlrEhbJV
Ou6EQBAZP8gfi22w30vwmsbmLMOPqez7oeDz5kvNSs6AMMWuqhQIwKung/jCFsXS
m9e0rJXszXbDVWUprurh94vA7t395OYiDqFGTEFga+w7DYY2K6sngwQysW3aNbgi
Hzgl5JODVU9RoKNCEQ7nqwVG0jmuW6ZteAXoERQ9t9OSLIz3uqWZLa6HDuSKeEPW
nr6hu/2hjtaehcGcbIy6JgpY3kiPmYX+2I4n1MJXhP9OX175BjBBEuS3RBBFeQPc
FpH7zNmsz2SyblPabMDyVh7ZDfQ0Rl/vMVvliR5n250cdpx6oA9mWBv8XbLoMiBc
eUF2e1V6LBC45ynFWhVtbd68XbMuWMD8037k9+MMmseGBLf9ABE4oE1ZyACNLcMB
mBXviGyQxaABgqZFzXVdu15QRIWviiYIzSpHiSGsXwzoGLr2Vj2oFnu9fk8TXsmS
MpKajPXpGp3Soq7zpeFD7ysVwHTjlNs10LmYY5PMrdihxeQNFB/xUxKHLOZLCxfD
21F7GXoG075qwMcimifUsaA98l85hjdDtfudtFfWyoiihtwQuh16ahrPmn4XPd3O
myWB0TEH8/CsMi5USrgGJPgsZrd9buXcF7T3Mj9GtFrz8ayAdwWrtzhpYJU1Ufrb
KSvV5EuhacFJ1kthH1BYJF8SpA+ZxD0hHmlFhuR9dtrun7D/cPc3Yh2t1xCdaP2e
AZDF6XoIZFDmh3Htmma0uv/n/maKwCWw2SNrEdxf+gUAaRcksY8VIv+chalWdkH/
Ec3+u4ShWxKrldeh1PL3f/+1jdXDodhiRpsHT52SlaO75w9GK/WbvtSoCMPFckJn
aqNuCKRdCcO+XlE3u7LEDq3TT3wcGbKGob6Iw+PibxAHSZV+G4JkkYiA/x1+mjmJ
LSAsuupRMxVP30ulp7cdeuZVS/6YlYRa39ECc+f71R/gQE8tWPI5IVx9rHP68nER
mLml7hUr4OmC1aaBKjg6JjQnKM4g2xXVzHQhpQqFSewiuHguUBQvYzRGgtkm0z3S
9nIgEDGnnJAkMvp9x/LeYUSBR+RXk1xInI7QSoysq3RnA4OrQVCpZZ7xrgBySaH7
CEKJyPcfqLOG1EX//xOXPu7irkX3t6w87nCZk1HeRhWhJpsH4Byy6Spy4IAATx8Z
KOYYezmU9Fayrjf0ZnEwpL/rcS8VhMtyRRu9dd0K7pzodVZ3jB5XbK9ytMMRCB9g
HdPdounD2IyljW+a2Ll0H2BTHYg2CYZc5W6HJimegiYuRKD42imleRIeV7bTtWld
uQsgW2rzdYLTDOG0ut5gIBFU8QioNnJuyUAMLNQXQ2StYL1PWJaHw4m6lTtjItR7
a4eU5++wAgAJvCNWTbmXjBxbnvl6SuOSvoOiWxJsoQPMOscl2SXVvV89D52Q0+3S
2WUDerp5AQlvIBGO9jQnBrLzXN5+N/4xNQpa1hsnilJWEzxffdwC8Sgd+zUcAOWY
FZfDk50Mdlixtf406JD8wD9cg8dj7OyWkQB23bekz9gruyD7f75vNGdfdVrU2r8D
gRzXBbuDFU9VnKBJfex1m+BmXf00sm+h8Zja15sAUl17RL/rt3sdMt5dpcijtn0P
VCAOPau3nFy5Xw0HOgz98l6gNkZxBAfIT7cCdGVE5lFQIkKp5UKHtlUQRQRnfZNg
5BW0FihvmWvUyi1Tk5jw5O0WpXlnBSMQ0VU+kCVhDd/zAtc8XU8OVjxt6mtlBvlY
rR6AAolLBv9CfylU+1dD1wSNTJay4gmqlOsVFYyFgWdNRiczTZbW53Ir4FKW/of+
p6Nbnfj6ruV2WmOLLnDF2//61AwXonlB7jeWCGKJcj9Om+iuNFxyLxPLDGqC47OU
YM0YiybiJGHRzQdSMsDAyNP5vtJSpSb2KLi2KBR4iOs5mzrIgcGJrBf1J+PVZBbW
daE7DxXvCnYy2AJuTiad9n2ZvYYQAcqxR04Vq8xbYwMjNTj+UoanwMn21UGFr4hI
tNV06PKHcR/tU092n/NFwyjcYDYL/McGck3fTsJkkvLH9GETwlwt0Aee3t3HQ5e7
ErDpcvl40wJj3MtkhV1qg/Eo/tpBd7jHrtYPRoecZ/KjJxQTIe4QRezdXgZ6Tu13
snMm2nY+MQCKrfKstlUePfXOkmt8pTJnHtLpWOBrjipWQjPwfs8VtZWk0SbRCzEz
ml7tlomTmdDkAe4SNsqODDGPYXPdCCF6ANDs8OYkmu0KMGDaEsfJFw8e8pcjllhb
AkhGb2WZj/Vx9I6XaGs2PttMnV4eF8aDPo885hybGATI60TqDdNmtKYFku/ztm1k
zmq65vfTH7WAbLljfVlIop7T2qyJUVzwVUBvF4o6jL7MXZSQLphOyw79Yrmg0uwY
5zsjf8AsqYayRRkHFvTzTu023BIjz4aLzb3TBvTMqcFOXXTur1jHtXnN9DLfRowH
p+RUMqKb7AfSCJkrzHgnfnjP7anG9uWSxsnnuyv0HXfEa3IoPr3krctKibeWc5Y/
eEy8/6FKGYI5JgHuf60ft2kC17Up6ZSAphPHiFibxdpXUibZPOl6HVtJEdoQ493g
FAx4cQZWe6q9Q5JaAfJbowzkuLEkGPfOHwmh0UVpIZKkgDcvLCn0RmmsGwp57l7b
Og3iIu5JV+pLbJbhQI9jKZ5IkYan8dmRVWDMsEXs6GuJk36aLRdExY2xGbw1cMw4
s0zUaDf0KYj8bDp4La+qu1kPTKVh4NBy7z9ihWjxIcBIzF7sIFaJnc3z/ucsNRN4
XdYvfibS6YvT28PwpAwEaHe3zHkvR+iabRhWWLkYlex0Ic2I2Jw/7WIhrtT1VXGx
89DuwzH+dm2sWEFPjFbt68iSfprJ4UbqaLlDN1tffNoYv6/EMaHZu/U9Soq4BwOS
XzAMQq4vE3xR/bQqeZULEO99MPFzuB3jUTeOglDRVlBql1ifjMliXIQXG9n88xKB
msD5/JUkVqilDnuzKJL834ondZ7WrB5GgxMroSCPKUo8VYVj4M+XDOWzComogM3O
jIaCASFeCqfSg9+yVqCKGsS//4HHAsdSLjApNn3V+SWOcBe6LehzYJ1Z4z0V6uj+
JLPY42v0mJdzzMTQljBV3wt38640iYtkvt+G+yfMJ7nqWHqih5nVZB0K3SMsjSv/
ksGnd+RMvIErxy3SK/kInTK185OxTSRHLG6xRIYOAbJS4AxsW3gNGjz0EICls9jS
i6v9o8p92OoRJTEzlTgCYv+AX6k+8vxxLnf7xAjVpSNMWHnDlODUfnBwdNDVuAQR
YgyLAqOn3jl6lrvCLCHKb5Nkg1QQ8G8iZhaD6CqkjFw9ourkPr7XzWA4Rz/Dw2EV
0Z1vLslwXYUwfStjs1u1yNEhzHW+i541vIpq7Zo748DRPxEhl6Tm+9nv2/bxA56h
FQx4M9aIDK9cpEX5VHphGgqdIdcH0X64j8GDvdryN9oD4RdlMMDiRd7HSMm5pDt0
mdMFmo/C1d2x34bxP8FXNMQFK/Ia/cKPZEbzzdwLZ1TW45bvrLgVQV2jFKzUWrsu
xqKBk4zJ96ClMiTlyAiUw6/kBYhRSXrj+hwW+WSTgnGpdALH70cY78oRha9X3sD2
UalWYHKCxDfSqhiLOiSlHMVY6i9JcEalE3P3TCcggP1nG9JsUde2A3HfmTLEl4z8
I6cPMDFHovtZp4DzVKlNq/JBetFGqLAcNgxLLQeGv/UUcTbr1xKjRBMB6TqmmYJo
PhmFFvGGQ2q1Kh+jdigUQ60HmPEUOcHvDejSiD7x+TLtjOEGR9Wx9nXxB9WGGQHp
fs2elR0ui/qE/hXFjTnEvVzVw9O9OrHRLVvHZeBl3hEcCae0uHcgP1jfC9rgdcAr
lmWc1mC0tk0aaeXoabh2+HA0oYFUUD0m2YqreIdgr4PwyphmDgnpPL7mkOwMYs0d
5uTgGvkFLYpNMq+E5Vd/Yt6f4U2vRPoTsrO2IyIvfjax8dVTK4B+/86EThXqPIc/
QreknuR53QukZ8tUNVJgeZbHY9QCjeICO4hhSw1afTJfiX7SVzx2zpgqNp+DUv6k
bM+9rdHlvJDSSyttyElk1jTxmc+1DM5ppaeRFIRH6fgBMGq0RfeOUfkOylpMSj7x
TtOHjrTsPWtXzDrWwZXfwqsjES7ThdxSCUrPIORPV0h8q0QCvhvalC5olHaMoMIa
baux4Z7ro72NmMMpAdZt2ab3BF/mDYyYSL9MwOQKJQ6xYdgpNvWXFIGEVobNMMk7
Pzq7YPNwvZA4piZwMXij8JhwIlkAChJk6+3Ghsq5BvYdsI8x3Xwp87QH1ZG6Cmf1
JOOw1d0i1m+Vn/9XVevlzhcxBKgzRY7SwdWQ6vj44xLtrlLRnDiFvzTP+zeAlFkQ
ETzYHahmCDTMHXZYTb9X1QUaCfBZjMIBf9XWcQmVOmd/WheANTbKdTf9v8RsAlEU
8c5Wh76cklCOoIEJ5LkxQs+h4kH0eMC1M83gv1QBf7AcSe8bs/YhbYek6au9MrKL
1orBUwmlNm1tTSy0P7ehBlL+KCz/VEk7peJnjXhfG75H6uEvde3cWmqqBleb7sy6
BSBeDNZW6U500bPLFNJ+63yCM2oGuYKKt6I3dYlhsBfuYDJyjEvvvsp9G9kkzK3Z
V31s03IUsAglk1pmOLpV+HUDOsLFpPCwa43oebrphSsSyLT+LzImkDWaJBL6WxV1
1khF3s2Cpa1SbsJLYo/Vbx9EBaha/G3uRkRhIGES5AAeSqazkxz0ipAW1byxo93Q
eS7hHNlTl+rfUEFNtjCMrdLx+6az6MsmL8bFaFiH1i+bufyAzyfZ/t+7fc1O6/5u
LVbAh06jCfYXZzUZnczfBrRLfZDhEVY7njWG6uay4KBtljeeLLb5XJyjyXewSsAB
icMUHWf7wjSbrJpHAZjdpjLg2MqNslyvhNqGPTHAcH6lxK83OuKAsZ9zZjdS/0j0
5G8Jz+D1aOkwEJV6soJga/ycmOMSfecRgSXb3HDKEHiVOcgdd4O4p1k8VW9724aP
kX1yqjeuMMXCWuJB7u6A0Yz1vlnWHTz6iZGPhLouYRuQojvldohv31S8rsa/Ixxc
AHXQ7rnfP682gGyjNy72mxC+MNxldMRQ+PqjyH3//gKe7KB9eG9okciRY6whd16e
FBFuz5iih5j8a+//QwW72pM+o283rt2SfZWUGHlxDuy2vO10fdv2Tat+A1Npz1dE
N4g/Nde0jYDMSTNR6BS1y0qLKgEBKvmlDVXyN4jPwQ0ShtjLwt4OmVV4Aqphe33g
iDZYKhnVLVRK5hEwHnpQwCu0pv3mf12Mf52Hek1T9haSiguHlhgUMxcQhlQbSdkb
lLrU7bRBAHqs++sTcFrvccJcnH9EKCMe1heNq99mtl07lCNXPLSdMzXMNoHcnMIt
cjPBDS/2uahnyKYpIOfBg2VuaWNLlnfQM6OwLn9kyBbqav1GZUtj3OeotyGhV1X3
Ihw9nuz83zXjNy94jXrVRSC5YTcT7bKRipYn+rpMvPBeYYAOSo+5rfK26sVc9j34
bVNeK0XJDkVbeovTpy+/7s8E/LnGW7UY0p1sLuM1If7c1jQJ0iqu1QzsF9+g4Cip
YMautHVcFEPFslMpX8XcOmNLWrHwmlMwlZIpm2OhHDrb7OkOxYn/uC5gtbYpPKl8
8R17mOBNVLHVHfqyELSApQJ6CI/t9K4zybUKn3gNtX1nbxVKCmUorsLsIyJ3sk1O
0arbCGftoJF1lsEBKeYo9w8FNt6VbAwLtuX25k4uWBpF4h6+sZW/ZwVLSW73tKeR
pf4CXY4gtwNeU5zrXuchlUm1mIYw+NmWrnBzVNm4SIwT9wyv1iuEjyKsGS62TYv4
1Qd5orj7XWkiRW9F0vLb9E1GCSRjRqP/DrNIRpmiYjflA6Pq2rWpdF5snaTSsXC/
0dS094ADgFfxhNhSSXkMTMkirnwPsLVaZtDAMX4Hzrlb0nZjUklLoJn+JiuJ2Bz0
4luvAVv2MB/lWwM7t9LuU+eL1yVrvVZNCy701cj4H8TI5jgbZy+ui19kHRxE61NV
zwMyxdITlUfpdy9jYYUQqqx3cl1Zay8eUIg1JimBng/xlXfl7Uf08xYfDe0QpRf7
Uz1aO/cBwW5WRSSZUtxoPZOb5IK09iTBiYhLApESIRE6x1lcydj2dxjb/x/QKd0g
eCh14CjbTe/fwsPKX2itX3lPk711CBYal1SPasU2Z52E6NlNEwwtlxIvNg01fSJc
B8EoLsMtdrumKbodMVzMJPF2nMlbi43br7+DJS2GDaA+QSfqE5ocuWZbQquXqlfJ
hGaB/fhMqlrXH+hxepAXSyLEinQee0FWE7QM7kMjn5G5SM6Z1yUy9aGSKj7vJvdx
utxiLCQZ75px/6y16wOiHs/lfSHfJCmjn/Id8u/OFdJ1ya8lkf5wQZVpAOHvbXJO
QOaYD4S6mhv/ZxPvh7bexu4BAn3ME8oLMvCJCGdWVhOXf4cvkLTSSPbNhZ/VOgEv
ongQ2FrVAkZ8MchCQjIHJYpiChwWA8nF0Ilifhvzcq/7YAHRXVoHvTUMGBmqVu87
Dzlxqd6J4XxuXz1e+kZjzaLpmNIT1yKkWvi51ILI5rG2A0LveWmdr2XLq4RUjEx4
Mo55XrvA2BAvx7N84O9znx/pWTtx8qbc+MlEPvenpBaJSxiuQqKV3/JAdpdTZMMK
7bhrfMgDG30I6WBcoOCCMY9lkN77LY1+5ghEaud3jZE8ocLwv8dSC5XT9jTX2Xso
8diSI+qJJX3sTzkZqM+1ScsT8PZSBOljZl6RMGog8v/RXNcIlgdBjfoIOe94fYha
tPBC4y6QY+QCMIUnnCxYMDqlQlAAJKmoVPKRdMueJgl6TbYKBDemU/FfzDHlsx+3
zmWxXfyHdNg41TQ7UDAiBdtB36jfasYVPKWy06BWvgGvSoaBFCbr42/zdYNKUHqJ
HLb3amCZqdsrtQBG+SIBkKbBNeWH0NrgvrHGBPe1jvcNojv4Kh4sJlbNbbMTlYwM
huzJPx6hHkpWVYgknVLeDZIbnn85uMNCp12FWv8ZQaD+KKgOHCpkSqnjLv7cJjaI
Qufkl+zsL6F6qnahm5pGzb+y3k4lR6cH9xV5dLIGLnwZb0LK/2s1W3q46GMkkgcC
dLfnHn8Jqf0D3Mq2+rsqSxOmZEPuWDuZKhfaFiWyj+WSYR0fVrAnQsWRT1ijw9yS
Ckqw3lQ6qdxc30xfA9cYRQqoXqEByyKiiwwDuV8Lfv/zRLFNPyKd8XBMHX5I9G3Z
UTOWnU+DZmTC6BC+7WYr6dt0SUBfNDs1MWQU70pewcsWGuaKfJbylIYeWB+25Vwk
NAKLIpt8aLWKubh9Pqpsk6wH5h0jhLZqSprXx4PmFX+PWFpaz6nyqsfaXnNpB9A8
m6RYX6k6lq6+ifhzR9yXUEHwyKMZbC9qCztOx6OJOuuRHNdhPP3KssEnm6u/j8lg
LhVk8RdjA/ABQEwAFRqaVSupLOuPGDmcEQLO1YUi4JBlhHSSxm9z/hB2rzEdNscO
YKR9+ONnRT5snI/owuKRwHlET4TzFndXLmp79DJQKOndMYjf9xTYi8jKq3vTyFcT
6l08xIepGq6MRdk9WvqXG381UucwUHQc3Lolqjy+gR/ZXO/C1Ld6tLFSWtqwhhAL
vTrUY5Veo8iQHqHM30F5IhvdNqx7eJvFyhkxH0KvTJcaADZHSlpcEuRU7RY/Y6HR
9xNHgP64hwN434YWieRtsv3Pk3mIUJ9O4mVwCzakC/b5k4IqB8qzD/8kbN6M3whc
3WKahVWN8qU/It3pJsBA3KJoYPLoKX1BWm9v6KZYc2sVxuiUEVUIV8LuSyxoCcii
fgKmVJI5SX3NEGS3gxwY/XEfRYUwa5fAhC5oss5U1fanr/EQVVnnOKkwD0pmINdH
Nyira9gvonqE7OllvtlplVBshEzQD3hxndMezH12ALhO5JW6rhStUYZlWr2pH8+7
fAkLkz0ZQ8OQDeYfcVeCxOA/TEHfIrTgs0jYIKJhzwgmFBNsFwEUHjKu+X8tGWNr
27w2AZ6IA39quY43EQ/SPw3+guFZ++PQM4NJp/vCJGXdDsZCbytX3rcC1nQ8Pjjm
HjFIuqXPcLcZM4Mw0KuC8aVFev7+2ptmdcHiVniXQFGPuKSHR8jR5NntUn0BDtOg
sxPIkAgNt5tY3Wc8MkYWHf70wjxFchsqGrfaTCMUwleq+Dr/UEYO82ep7+x/yZYh
FOUV2H7IdmM0ogcZ5L2hCxKkYQgcd7G2hf6hvBN8LpsGD/XPiy1+SBtPqDfGwfH+
nfbwpNWNmdqRk3MnZP1TuQVJs4WZYysKLrlgMwLOzDWyTbcV31guUGCHA7OYuR15
1f12t7iKdK9nlDeo8c9nXhgzZOYYYPGe87gvByPRMwb3kKGg7iaYF6z0SgMyMpp+
VQJb7HzheyUQLClUXf4P8ohJvI3y8mrDuj6wrnF9ClmDFxIwVBURs9Tev8ux9623
m9wbN58SvpSpjXhLS2RQJprcx4ilsUfTp9IV0cZSzIUoVUk4GiVGpBRJdqCGmEPI
osfM6OvPPJ9BSXx7sAXrZd+7xTFpzyWftE63ydlNgVJZ69y6rK6EU8WDP9ZBGIte
VAOeYX5DFPgUqIPKitiFaMpixZB0TVJO5OnMabahxL/oXTNC9RfoR+jWV6DmWSXq
IcrZkdBq63iLPuu3lxSEgk/R1YBaImz0oeF+6xrSIaM1AOp8FYWanJTzMCmlrms4
QM0XiaG9TBCfIR6ZpUHv3NSn3JTVcqAGdRShD4xjljMVGvCFTYhXx30mqm8tE/Bc
S1D9cLib73onjk0iqC3g0vQQU68L6Zu8zR5m71MzOEWlC52WESSd5fy/03fx5DVN
r7rHt+Mx719r5jVgecphcyZMVkKYb79VeV2WuPzaBsRpSjAMCfq6w4BPbsY7y3Qx
smhdtkErox/vM6c8CYkFcMDzseRZoErmcNKkBMKM26gG1XdzccyZ3cK0959Et9fc
GdbmftSJ3uG4i+BhcQjZV0OdkrrcvjfZ+IAvzTA1CAdx/SCBP8kWJy3oRacQtSIL
Z2Qw4Odss10o3q7mL27j2CuOa5M/xy1B/B/LB1yCqxn5zyfEB+Y+qDNWXjv/K4oF
rYijHwpwx+Qf0vRAx1nEtsAUJ4LCQairtpBWg46K7N/t+OUYUkYDQolnbeN9FiSP
iPA7QcOmFmhmS67Jaka2HmVbfQ6h+EuJn6n7UeMOO3m8mmvZ9LYyz6FarGEXNq+3
8Mx9gP/4W/o4sobMlixwqi+tktp1W9e72LVQHkILmsae9XDVExTU8SATNLJjhgxr
SKK65/PLY9aI7INkeV409GkNoZo+O+Cv7HtZgbeXv+CrovvnCdbmApPTw2IToNIn
VqXxRVBuy3zErz9Bzdq60IevePANC0uxfty03WC9gbiVNEaN3lNaBcDondUz0urE
lMrSCGCz9+7WGLPuBzOU76HiRYC8/PNYqAxSCOPFBz/NALEMpCZ99V6v6vBDDYeL
Yzs+0OWjrub2I6tdw5MfG9dwO4XXFUeIuc2ag7qkvRiwVLC7GA8xdPZi3qWZCetl
4XRNiN/x2YKjRg2HmfQsYTlcNkKV6Z30kw7b7QGULrGhzu74lB+sg9JcccTM4Sj3
NWP84MR45NLiJhSZz7OGUG9rQnqvliTeY/vWb6fa7G8ERAuJcv1juKB9pDGmQm28
ySl8avGzmbJlXUKOEqOIJbCpj9+WSHy1ZpwcgUvnDPk+evgKJzsgL/GSWoNI4g9g
RK4VtCfeS1lWTPil+VVUuBt650PkXp1ma/GHnCylP24jaGHiq0YPfuXxCxjzDTAL
R/A6UAR9K2HGIvNzuvNIdsyAA9hIGXGZjhNb2z72WedDb0vjiSrDVp9NWEJP4fud
HQYamZfegZe2oB4PCYXVC/LDniI8ctIxlzMWYiSVYZ4VYGgwNVym9riAwhoTuGR2
Jn3AEpFInSw3tpoAY4RLQcE60zurLbCYkDYDNXlIIWhS7Ju04UwHOPaeA3rAJta8
vlf5UkFodvn1whaLFL2jjAvWHRw7LbKzJmD7pXYG2YSp8oqZHAWUhLmgqqzTGs1C
r8WrQxBDftlO+rqy3lgd4G7toA4YTnIXAHwcNom10i4pHrqXqYVYdI9TzoJ5Umzz
BHNfL2CEJHg+H7GoSIEKGMxOuYXg4oVT+s7ldgchKX6/hk9Ph8q5Huh2Xz/OUyQd
yIxnNu25wdrD/HfDU1l4+5IPBIbZaRbWBIrbQKN1qk0JYBjNeCZFB8HX+6w3KmQ3
m5ShUAj/o+S4AQXYmR9LDG8HRr5QnyTWl37UKMTC45kx38AjLJNmFp4vefiANWTw
CwMWKQkuAUW16GiVJzAdqzkrKcHulVFW5Ty7wFDO+JPacPm20K/bFp+4Y2m9DxRa
23VgU+3uSJ4BnoIHiRyk9bkhBDarcZ78mK3whqiHmqcQ6Q0wfEzEHWQzXll+f3sd
+DBj22iqzLqPo5yJmLzHeN56mmQsNwhBlMBeZkXE0nt2gZPW2WTaOf/rUmiRbzOe
gfl8T3KukDyAe6CcPfuv/FWweaTL10LDnHbVDbG+oTp341E+uTCbKk0MotbSgA8c
rmvQBZUaFE4Aw8d05sJRby4Q7t+0+jTyY8bvgA+VKeerqkZEnvkey0ogsEM7Ds7u
WD5XqZFHxErtYrB9VfTEu2u875G03HkYOJPxlnpkxSvFA1RSficzEhnzwzGJBd+t
9nWZT664ZLWQa7KIsF/58mYwPeXjSGxR2XCy4ckbqQsZAZpFYwYKQAEYy+TxKAlK
cIizw4rRgnIaX/J0f1+Uf/bZmL1DNRWiU0uf5uXWW2sfxmxTo2rNJIEfVIVYV/45
mSfW6LKuDtv88SNEX/fmsYu+ao0kDRt+aszcn1iBIzf/Pi0A0fUC1+07aopIi2Wn
tdN8C3iZCyo9rsE9npr5vt40oPW7ecw4WsYUP1k7IgdZm/gySsmSYmMlZbB8I5FL
+VaAuMYRSt46B3NPxQSgErO+jFyyNZ1AaXxZ2orMjvL308o5NB9PKvrsd9D9z8cI
M265X7xOsT0ESzpTwk7dsIr2sMfARYE1+SvcvmHSQy/206coG8/UsbVkNn+1tkwS
rLYsIBXWbN+y9W5nsqFBasf190cN4OWxyyvFq5LkBXCnErqr7N/+Foe7z0DGHNt8
1XNcioZjQ7QcVJbloYZdyXthCDQWzAiIP/K3zmnA8Vk1HZdsGJhZACFSLnfIgrka
YbKpNgRccUHCp7J1KjY16Q5vZhwk530dMZVpo4jGJbdawIk87pt/f6mU5q3QU0YL
i4rAgXN0nyVVUQs6WybXJ75uwSN+3kOEFn5AL23VBdq8iqjxK9Rpy2qrfEQMwMK3
PuTsDfvXx8gsCtgc90rXYIAE71NgKHjQn2MZGWl35ROCGZ0gI2YbComkNRyo04kZ
Ok5gwTLHrveMcxqGS3p98p8YbavxbyHXNNHmT+YaLVBzIAW7OYjpLaTXVJXYBt0r
PaLQYU9mk/c1Ql0ZkM2WD9jTw8iMcbym+zEcvB7nAm4KRnWvtURuSoEl+hAQaHWg
AaZX1iCi/F3fO+qh8+yMlszULCgaL29+szQACVvBCuvYN0bXI6mzqA6M5hlr6dv/
UZvLJshGJH2K/MXd9oeEK9xPtHhYoXkg/TcpYswoKzYHV7ddpWhxo+WKqJ9iNoje
2CwQ8s1T+pzaNiBAJCGWJEoqxXNuYYLhid76amMSLvPwjr9H/XM3cETkUFzcumLU
+I1DuWq5Up6kStALChw5+aeOs8NS7n4PpSUGFvLEVlOYEGL3zPwbXdNEMwqT2H8C
IMF3vjzXfUc+DTwrryoE2+uf1WBJjKZGu/BKwEogbYIV2Dtb22F/LAMiOWElZEUZ
ug5aTb6Gesyd1M72QgUKiDtP5PHa4Ha8rfNmqqKhH4G2cbgkImYmufm98lwthDR/
0b09Utn5K7ilp/xEKIkTJg==
`protect END_PROTECTED
