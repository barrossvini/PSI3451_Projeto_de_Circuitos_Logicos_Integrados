`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
liBpPNpMmMuAD98r9OMPZoFTRp5p6JVhBeXml6YUiK8BbO8rZxAKv10dcN4CJx6o
ToDYacfmeDiFAnB83YNiP+YvPwJhRUkncJC1HzGZI5+0jLXeDM7N7ljd3tddgB9o
ZwABA+1Ij4rdlltXI7VVIh8TDwELgy9Kr3GX4kDMOZQX90u2eheKACZnXPZkamdz
rX0SCirPWnM2Ogs8Wm3uomR0RqhLLP2CCN806I9IYYygJCwPkVUZetuik3ZsamI1
NB0IXJpVPQRkCkNTMfMERWobSzDpZ+fqD9pNXUHh4mG89uNvN8NA1Wwtgq6OxYUH
eldqTpznVFaI8wdgWhJtxRvXvnvuwBh/EI5Bkyb1d0M2KMFfo2sTcqNALttENetN
ch/TA2b7rNIyOPApt0Hq6wc50zu2aNdQ07SI0/GZyhpIDejxozWbW9JAFF8GBpEu
pqVtnYSzZqInI5qMjuI5GS520qv/iVCf0KuWOsSCgMrU6dTkLtOkKCe6Y+FBTAYb
nOxbCWWCnHpKospTYPQrYXZrI7CKdwz4939UE6ccJSrq6Q2OleFjbc6EIL0rCHRl
ayEXutEty5TYSiAbwaXLuZi9GLMfDmeevHKFwyv2bT7fB84ZCGt1IL+g2Wff4jpL
z7F/IHRhEfPKcOX95CqT9BZINQ+xCRKjJflPDlYjclPZn89TDHIg3BENtL0g/d1j
AFIP/m6Ud6T1bX7nGKHGgDc6NQ1F8gWGO/wijJRat4l0PleoGUVfZoFw/WwXVdeP
Tq+VSf2udQDq380263O3WLQ4wS4j5h1gUoNB9SyyxWV8mYeiI/NZnjEmws68w8/5
muiF5YrwZhC15mKn5Q9pRTyRKTnwAz5DPNfo8NXeO5l3o/ogyPErURhll4pLTFc5
m8AZJ3FYvnOp22kh7Jc2ybAeZb49RiBx4CejUiWHY86qdUtwqRRTnVWt+yG4Oe0a
Zol8JPtLSy4MV4apHObcWK4blSHB1l21RNdeYX6VU4s4lACSdoEsQJKsWHlWZbZr
jXG4pT5nXlvDeUc7LQihrGo0DACLiU3jQrVyOndxWa0al2ErUj4DaLJnR1nF6Bhw
HaqvZ4gBG1UZ1/OKZUnSw1CdpKHUvaL/JHPm5MxYyWal6hYU8pvDYFjEufSuV7d5
LOJLWUm+rnVhd3so7Rges7P61BqxC6w/sRkhopDVEWNC91uYxqQ6P1JZjXAQNSAj
30F7akInYrm6iIb4pNSwicusZXsua28wL9ebYW/bHJ/W1z8Hpb0xqNqENmLxkrmd
ek0ERkNmaIl6QR9i6bEiyGaJ02cu640E9AJY6OLsGINAlZfTSUiwKfINLbUUFcWW
vnk5DHvS9Ble7hbuJOt5TwDhZPZkiz0Z46K/+isntFvGG2Q67xsgapl7+4ADGibB
19VsgInu9/VSsDxOvfavCHp+wRM2pbeyFi2YvCCZ89wjwgseJBjaioiedbvXJ0ar
KSU3IUj9Nr4DtiA4AFjWi/ARnSrPe6cvDz7o0aJIKfu5U4P+7ABOtEtPrKWOLMb7
Svw/aeLzedwfNDk1QrNDWCV1EHyqRp4rU6RrEVxiEVmDFB9soLMWUwqRTj4HsDZj
p2Xyk+jquYGnUop2X7QX8U0eae2FzPidzc4OiU9YbpAAuU29Yef+8qSyArZ43WfO
e9DR9X2yCPtYkzXsGdOOn0oaClR+fBfhfuOYmtw/JqjooCyIsRwxMvGOL5VPfadr
/V+FnAkTGE3iPNFgX5LM3YC26qN0RWjs99gT64GJBsTZJuCWl2B17lB7STWiZbso
ssA8L7DOJCmSIzxS1UIdfyifR5DdP/yyCCQUehWgANW+hwZrOrOk1O07TrsZuNYB
29aoSymCFc22N86BRPZfyRhuilnQH0pkEJUstgM/L0IuC3pJykreekg2KjPI9sC1
GyYcpuuhIxjdt981KQ+i3HnotcguH1Dd4kJxtUfxn/kN92wj6rIYk1LQxrIud0eu
qd+CROa/5hyVnrB19u1FercMAT8zAZg2lGmvvUqFglNsfC4SRQGxesli3dw+1q/8
Hw6hq0W+OOzJMnokRLqDS03x4umClmSJ8cWtb3jyAD+t3wzU3sgzTBT3TN5tVG1R
xxk3e5HeLM8VgtM+s1rk37xYaYRBUjy3QzoXluzCMRDhd2G0TqnIh9qz3YezM/BG
hd2meZuLn1wLJoKVC+KizdEwYMUHsQwHaQgPo/xe0nY0ozS0Z2bAqJaq3k8RUZVx
pAhxcXORY6lKfj7sAX2VqNSY5qCt8vsugh2G3z2KhU04iJTjYXfMTuYLozEcBRIs
I4D3g0l+VD0pyrnKx/V6sgzT1k4JxPo3Y/0DZMXjRMqiNGRt4Bpl7a50qTDxhEch
k9P8bO5ft23byMefZ8wi6/ToUPq68mBgWtqiW7/x+lN+ZhoqIeGdeRvMrtaZLgif
3Pl0ElW4MU/aQnYfps338FPsioUjx9ecEvNokcL6r9QT8mPBgUvFhWgdwA8hTjnD
SkYG1ABson2hvDvmOkjKq8+xjsj6EAxJsuyB3ODy+CaSHgmsl1znY9ULxETnSb3/
U2hIq4uEsmM46hDn34isih58Xz33zM5CH3dRpmeTDmLe9BDw8KkdjLAY4X3muxHB
W62244smYoHZ2TcQQZogxLAPg/5o7oPlDZV4NlCXSDPOkLqOviHLbcfwrXQOt1QM
RsErhYp6b0McXsalkNWZ97GuvsNnVX0tFD7bVQDsdz34kyKsE7Nn1vEKjezV/YWH
S/rQXu2uq/6X9NnKHZnJEMTwaQzonrHDc4e2/0yYRkpqaP0UOVERYBdn7WV+rHyz
ztgZyuKJy9sPp2MnyfdCa66+W4yQauOJ6XjRZautJaPAs4l9HXAQ2emkhH1ZS8gx
d0aXJMqsBvkxC8EdjW+3DVDIuo7aqNHJdZWgw3dNmAgwTxRcHeQy0iq/Q2a46m7N
1tvmxN6uO1tVGpTLN0qZOpce13ZAl1xWgEjVKqvUvmGF6RoFu6TyJYDmlf2LlJKv
nI9Y4EBNVOyIcbGAGJYDP+LC1+wf8MXTgDVswwr4WIxIiA6LfWfY5zMZp8B5TThQ
cqQqmhozejVw4960xq3taX6do0qP9yHreW4TGGzrRRAJs3JlMmOnz5xQ0sc5z/+8
ub6G0r/jz9ERRLiI09f7Ks3Lw/wj7KXb8FodzQ0veD26C+HtB9dAhwYyaksAy8AB
xsKgmQelCUMW5R7ctBJcpsz2T2hxG0TgNBa0y6Pyt2aa5LAoEp4V+1xrGw7eBMu1
yn3oug6eDi0AT2wqjP5ed6IyVNwraBelY1JTmQpXVYzVurTp5G4Lvtgiw+4RGraH
vvbKXh2WUp9USR2jLh/ArypWM8h93bj4+Tj3EWSwl4uQh9Jvk2T42Ha5qFFhJ5QE
S5RkWi3zNHqqHOGiuHExO96yaOOukC0lB6jZg6kSRDIjHMMYUVRKLTQ9KKqXV59w
fPKqSQZZHXc9y59qLvnvtn2TTV0ngCohfcZNEuB+C/nmXrPkttT2v+If1PjOQHkE
thtCdKYNhICg6ipCe3lTGMoMQdMLkrNan2U5w4SbBYPAK+6eTNO7uZEraT2O0aK9
ZsHYknkVga9NFQh2Fl++Fm9adGnZbOOgVX4ci3TgFo5hJTXI1U9m0TgTVzDgQN+k
GMV/5C4Mg77aLO1gJe37F15JphCCkCQiRUb/lf8YF4MhJSqr1wSqTspauzsXwIaF
C6yC1wFl2BMhM2niJPw0yu7Q3h0Rmz8FPUnK4hm7w4RfHJn4F2skMxgZa7VeC8Bi
Q/IdUHDclhElh+P8CzMLC2AgyM8qPpcfdfjULdKxTXeHHMjdCz5bPbgSWBpEIujJ
hIUT0jzrbF78E3Kw3jlBDDY56ssTxQvWXGZM3NleKoDzKXmI4Pg8P12qDZc3S/SM
iK6ZnHrXomYVHaQulRAl7TXmex9AAItj1tC/hZPLWXgvXY2Z3zp+60wErjbLuWiG
IqGSnZFVOHzVgjQBP7Qrs1bBw1ggUOso+a4l0KlqGzhRw9kUSvMoewd3+ELrwIIZ
iUbcT02cqT0TZl+LmYcXd/XvMJTWhHcezDU238HluxJq/vPlSq8vmBquIeDd6bKa
5+Fr/gMlaQaFes0WtgQpFE1/GRdgIh3M0wz+NVY/vHQOGaBoXelaqfBa3sObiMmN
e9o7+G+S8/W5mXaj+Wz7vw3iCVphi9ZmNYo0tj/7vly0Ja1MjttCZPOjPE1jv9o3
eLt2kX5FlXz9aJDmYsdQTkiWHcqMp++ygJh+zAXpJUczMig/wduMgGT8JksLHNux
jp9rHbk8u175dJdplkajWYnT/EcQmH/w6WbRhWsCwN0pnWLwZR/D+J6RZlIQuc+F
EHn9YyVS1YIHxcO5noxhBIU+FWI6S0BBt5qujgfMOwvNfC6hhEXad3nIroM6RmRx
WmLIejbzBt882GgnG7H5iZQwJwYLFxrevO6lJQtnn3S+v7xSV8NnKZgL9pGz0/oy
qPwzPSv+iavdsUiaj3s2p2KBlIYTKqk3Sz+MkUwlmwN8vMWHxBCqe0ENzV1qhVPB
hsaZmSdHyCjLMk/c3RLfkF6CPk/+LgFif8IJs4zVmWWE/5EtBoxvCSbMKH0sm+Tx
MwFple303b3YHY33wkmGMVqfwWhYiLSMDnlmlQSrVZ9D/+pBiTyrMAjGPox6kb6J
xUbRTJoIGdTaLhavH/s5WV+S1+ndzSdCo78id/ouyodAVPdEJ6jiRdJsiUId4801
VzA5fPY0+AlHk0IkYiHiKPnzixPHUSM+Eg3Kg/6BwwOiTKFCdnXP+BXL64Pi886D
IKG/xJd/8T4osWaOI8pVWPdm/3Zg5Y4A3j32IUSkm36mkNpKC77f13fXu4UJElqa
pg3e4TkPjGe1xyco6ha+aRRe3/AaXujak/xvruYZee30uSgu1txIDE6NzWm9TjB8
jlIvSI3EgNE2d6b8GaII4CTbtbGbXEis+L++EcUYqRNcrCafSXsW/qd6l50UlroQ
sNTQ9W5uUhPzSZqZ/yYkOU09Ocxur8dGgh5qU8xudltlhYxhVmA0aYSsTpwld3NV
Kf0j65rWe/w9OJm6X7Kewsnfttw8Vyn79HluXmwmBMhmarS7de5JIIGf9XZjMngV
L5kwaBL5IswswTR0IRnuSKSjFgLpzXlZzah6p8UTvu4c8XFs5VYtjGxBibsxWpgV
pnV1G0plBXIXM+E7MNe+hhyt+3Kq4A5wFX7daTdVP268LN3rnI/Hiy0+hTk3g7Ud
2R/o7z+FSwAaJDuEPtbDTsQ3akrqowceokS+4FNm07HdP5uMuViYEKKZyoE+kJGQ
6fg9k3UC72pgTsjL/nHJUAugCr1Nbsva08V2yMzzPXz2Whss0HXb6UUiIWNfEqn0
HnFkHD5UWty3xr+jirbrtxaEuMqFRShFUxn9LB2BzNc9bfdPwdff6U+5KiUYettn
cZM108hp+gBJB/E1eDrt940/6ohj9nqUytqUf/Q4rdaKFv5BI4EAfzkpmzPMyInD
hoKHj1Qwvc7PFjhJg0NXlvLoFkZK7Tub+ML1A/tqRkD+oOQa6zgXF99eInIzCn6s
6bTmSpOiOxuioeV0YjGCRVRZFHNNtYj3XFlKDsz+og7uncanj3CZePCpkuf9V8MZ
NglKsJCLavucEAHerxNWUGm7kRvTXYDXXyGSOtvyxDsd27PS54AfRGsIoXBL6x3N
ouZJ2OIBebRekLr9eS8RxH6aBVZxAectreVb4nK1xuZKTsvvHZ7tYLLGYq5D4k2/
AxGrFX6ZYXxQO02IiEAbcBMJMINhNGQ5st9y1NSaZlWfQlvswdiilkRhSXmriO5L
uqZiWoSiDy/p2ZyuXya/PnCgzs+4YuMwQLvvHCzIQOmH2XuxlslGvhUrCgsS2PFH
/Np01vZDAwxzFjiCx0mErY4OICh/V2/GQFwultRHrKA33Qx82j6cPU2BhrwAOmtc
EdTjTf68ziiTSH0z/eDS2XsGqpip81uez+b55njLZIVEQN/C1kFtsEwR418F+7n/
rhJIfujIozyxosahrBQnEihBA9E3dYGSVsU0v6L8vEqo98NCVAE5Io7KMelZe4Zn
enROXKaGW2XUFukJFqS+nlL/nvq8ZTDwjc3zLy3vQAWl1pPt3taMOSfwL2mDvXkX
ostwucvkDwaLQdbxAv+2/uM1ohunvMkNgB87EIOTOnosRoURQgPDu1OWUF5RxggL
I6V14KcjGxqKU/0k47Q5b6snzX8H40y7thgMk9EKrRvAgv5xIH8tmETLsYXMrdHm
p4VHcbfLieSc0QY8ZIWhRPtOATEjrqvw8lIdMx4+BY/dWgV61YC+GMxHarXav3NN
3K2Xet5HCk6WvRYb2ZdqcTqjPIsYe3QTc0TKa+GpYAl8C0iBJ+BMiR0lc6VWVPOR
hGlyMiy31seDYjrH6PkZ1GQ/iOOW6lXpa/5htROtq4H2H0W04rFo5stVI1sQRrs2
6SLj5DTtYKwROfIA9QoI2ENFiPpc+nccQ9cQNHiLSBNnxGb0EmjvAe+ulrExfXOQ
/LnPMbDnuM2mhqQICcy/CyLUlWDKe2YVG3Ofwm9JgygHyc3ezfDOVlTMq9NRMbwE
jznMNpV5b2om/+vqdCJNu2B/UQpHRxNv4R1EpKedWd3hyYe54Jy1eydm6BYKtbH1
2doNweWC/hdUl8MVueva5vJIicT8E5cIVqToYLgARq4LGPsHK/jdRbGWo2mi+mRR
/lpbdiKxM2ulesGKZkY5hnM+fUhKy1FZPRFGbs41yUB7pZMb6Z+ePtc2Hcd8tz6J
ft8bnA52oloqFo3TB7w73hy3dunVhbfjxM+tm3HgtPrn2JxGdmWJPyNt/XYo9jKF
TcZttdM9Pb4rYL16D1imk7rz9e5FG/9FKvjgmUTUoHB4O11c6A+q0BqeI2EwfhG3
3nBnBhKEVUbu3GDp+o0oU9i7LvcJoIhyqsGRJHbciHgFKwUdtGFSRio8XZAzZNEo
wpwzUEQazuf//Vi8XmPkImvr1ezahlI7Flq498J1IVzmqcmDBhhrerkekecoud7T
JRiSJTLjfrr0tncQ/24Z1z2O47kYDxiq1i51kN+O0hMcGABwHGftQ4+VMG9ArL4I
t7GYBPsyHHXCbuhctst+luHTI2cm6DVUrQFOSt/z4gWKo/D2KQVQBx3NIC50OyoI
s6aAL8sS3jdPHhGslsVQCrijqA+HWQOI38+jdBmO16wHJR0MK1ra+A0dNwn4jjbS
6GSjNI5hh/Omz5LcogViAQPDyEe+3t02OkUd4xOh2EJEZlXpEIQFvf/lw7JxnmQK
/xl+kd1JQTVd30IYHWRkgfmXqZhg/lj+Yjjs6fK1pSlqX0JRWYnR0exTktz1h/FS
5q2Sy5Lwo7ijgsGDscHyxjnbKiD6xVkVOHhwAmnPxDK+RdL4h57K5Bq/Kl/RnYbJ
8yXeiRtH5pWO/sSnoLwSuwipnlfY4QqZ5oDKaqwhJzpeGKdKN1EoBibK8UiLWK+r
Svbdacba6qgjezEKpylXKOT7DIi3KCbFtc0Lk68whZ3iEKkOybJKKfyh8ZJ01jck
UwfoVm3JLe+RxiAIu4IT+C0dXft61Us+ZxcUlqXZ3pLqjzrbzhYHp1kNjE3TrA3O
qMlrgdbTZLnJR023Lg9m1VxPSEbYpeMUrPzk2gffeNMf4GE5LmKwyI4XT9zYFyVD
3NFFcLHOl0JstYprzSITPUrOFQQefmIK+OscmDPUCTTqO2PpfOfTenBVDo5w9LRJ
lroHhdXmbqoPIO2JXbE1Lyc5yVyMAZZrsBtpIIYipp36i+C2tLZ4fFN487arwNwG
4h/yoAUCCKGdSTjZSk2W89gJ9vvvk2E17yOK4FoVUlin5Q5F+TMFP132fN6Lz3F4
d4nafEzhI3883/KxQmKHAK8YSjQo+pXpLBY+apsJ6vfsgBojwfZCnofkgZuxONUU
yAQDUhrhDUtcFr2nTelTtQjO7HPKEBLDvpYTagl/fV4sDMKvqboEzency5DHr63I
wuBMP/qMSvppNFix50ZF6nWTan3XX7PD/tzR3ez+7dK8u9BEUSna/p3xIgYGfblM
2xoPxx05Gz0E4wZNfolLHAq2PXeReH5hrm3g8f0KBcel+5CkbZqa3/pVSBppl1ls
zFmOEgdebKKmxD/BfJtFdKlQGEsSa6mygxzIOjvnID64fSOYQbydNW9rtGlN6PTl
4ln2ZSzyAtleRbJpsD34c9agag9uFD8OjHCm91Jh2mnVlW5g5Bdl3Qvsjp67oA0o
aUnGTsZR118aqoAvEW48z+G5NJH00npEKeMzaxAl4VUFIsEpbVFn6v7fG0VaMEsH
VH5WQmx6RXKRNEPQ44RivIzvH7SgVivOZ+QQLGWP+2gudCEofctpK2XcaDV0tpLq
m7BdX97jo2/RrqRvi7di2jVJjXuce4ocO6Td40vBVLef5BrwT4u1QRecysydnVpA
z5PGOne6J/hXqZ1+N3t/1qF7JjYImcJANXKUMRBAoaD2OiGXVdZzW3UC8ug2oCdb
DA0UfesFOShJbgZjRT2neCVIoCRAxeoiXzQGezg+VgCqPPDU5fN8KvLb4uK87lC+
Csi6dKBv04fJjcQVwZD+kiyJMcb5MeC+tnBv5gUOD5QlbNMVtSYTHWG0YWIrA590
4ZvX0sI2Wwjqmk/VbJGRz73JtD9vyBM2LID0IkPttifPYNIU2du0gdZm0ZcHLa7e
RCTuBdJFwomBmar6a8ljPWkF0YgIbPcxYLzVhARWWG1LhaqEiSMXuRz0aQzRa31n
D5LtqUpVlf53MUSWqRSUVYRUxRpNjIga5Hnbo9otYv0g8ES2nj0QZ1Z8DTpPJGVo
VjkOBHnzjhttuCBNp3HUCo9iowN2GAppQ/Pz4ARPR3pF65ODNDUhOdBZbEIFaD9J
AZjW10MTnaU2jpTxl/ZSKLg6BN7QITqFOO0gpwUDF7LiaEKGDIvbffSNeWivxVXM
25zilIs4NA+Ll7AKxBblcwsYiQOsDA8WP4VbR/uVgA9LtNdgvKGKkvYvBzNHqKT0
x/CXpciUAdFhfweBRmQM1B6aYgXoTxP3CW2WQvRSds9iYn0HZOICsVvwHNtEo9en
NpH6EIDSJHcdbUblU9VWRzhPtJGP/KjP7YTkU1mC/XIvkgBf4u5Cg2YXNaoD2qb1
Dmd5jNitR7a1O8YaEvH25ueYjphDnxpjRDgYfgWUyBy14dej4oc6RICujzDB5Zu5
NwrZhljBohyL6INuZPLG4zCof10oHiq5gjRUflUBelVD4F2w2R77lPRkR2Ot9L2R
4bOmK29dVrudNt5U8D/vCpoJB0c27Z0+Qiw74xWbynDK8MNYJpoJtgYVz4tqR2aZ
nyk/owDdJETcF8rX3NsaYI9WOCKeLvoEelS/MDQkj9LUo3rXkvMZJr5FL/K/v69Y
kgrb3LsTA6RKRETqEHjf505RdGxO3YDOVmBVxEI1+hWEAhPpkOexcZcDG5nqEmIp
zXcwOUfuLyvrlD/4ysXFyr3ckNKV9wAq/RMThMFFt6OTeUW4EX7FqatC4EJdbxpM
dJIjEaaCqwpu9/3LwmPUn0fdlU2KjeGIYwvSYVkgc/qgtAcDMjoepMthjUJ/psH5
pPKhrgSmfou/OBiDMlrDp8W+Zw7ZAdxG0zUWGabyGYm+LqrjnRIWhZ7iqjcUZtEH
S+4UmF7cwJ0KtEWvNWcg1Mtp8WqKtj6cMH6Y1zV7ebmYOQqgFWlROA2ZV/qXQDed
5k8Lyf5E3KJdlyMREziG1pn9y4oye0AX4ndzPZp82b6qwNkUT4zBVEFqBiQBaRBv
Aa3Ib/ar2qr6xpMMpBEgj1gJQNIeayXWJnakkLpjmQ+tp/r7fc02c71JiRxQxq3E
65V34w3QUdEeHwE/84vQdypVADFJiGSwxHeaAy33iGeA7bum9WfP2VnZVl8QXJyS
WguBS1dJVXnqUQqNf/DorehkdzSVaXsCgck7s27/A3mbn7cw8lDK9zzOAid4cwG2
gOlZodzz98fGP0SCrlurz6roHmg7oaoJv/iwMzo/G9KaZRpQeSBABK28Q2yGHwaV
VmJpIcZo5GfYucuDZeDDuv3A2VycsAMegJdrDJKtV/UGJAdoaswSWmRRcZbrqjca
Z1fqUGNPI+DcovsuTHmmu2oL7Lm1McPPzOojOoMTvx8cxSlYTIBTFltZNG0eVd+L
hW8FY3wTf0NGpDeNAicKOxAvANQ+JcDF8+Pu/rIWYmYNokbL5dvB6Xc7PBbPHKl2
t49h0BOKmAvy3oIKXC7OxVkdxmVfpvVlQFtXrqg3mD+r0HlAWp5eCMXKeqjUjfOR
rAVgxhXOIN6XWYrBBPqljgjn8wYR4nI306zM3pzItpAcnUXwcM8slPxFvvt1ez/p
NFGkWl9sAcUPq+tp3OiETTcA0ke7MCaRZfu/BKTS+4HzKam/AYj/JtJmYkZ9rkZW
G5YWz4JL4aAsIZXhfmZth2VY14qnhswIPRbApzp1l7bmR5FZcbmcYCAOslBBuZsN
QMSEbr1/LQre/tjLy1qJ2GrOLULw+O7XsDNBFhcYVz6Mq7BdArsbf4SLLE9W6jQv
KCpbh2HdEyJSF4IRGbmzaf4oIjTcxOonvbSu2MrkFy5Jp/LnOI10qu2er9vcbNN6
C9/JHud5ejSn/zvld03NuO8y7S3PdBhpca8e+XmABdg7Xw6//aCughKGGosx8NhF
JfSlwZhHUGNpGnkRb3RYAZtTuKCu/9tZ4jQNQCnlvXp8Y/ZyxsEUwK5CDwCFf7iF
TyrALMSvQA3kPFnPtOFBrV5BtukmSji7lwGdlN8/tqL8WcTGyjOMtnOp6seq+i9a
v9YgAG7upQa11RSPbJzIRxRjnSYPTrYUsm+kKnYtfew=
`protect END_PROTECTED
