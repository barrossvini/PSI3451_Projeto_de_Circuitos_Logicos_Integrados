`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a5t8IUDEWrNead/v1gHrsuB8VU22y/my6elK5YaqHFJjrkywP21gx1zoXK2ffsJw
NgvyYwfO0e6k4CIYQoS+qhLou0IpICyiNjmna9IWanF+3IYDcusUzV468Lr8QaMw
OLsrp4kcBQ89gQrBXz4ePU1vwVLDNhrfYe+ahXDmX02xSQd+F9TI7no68QCd6Ynk
VsCIbNdhPVoNj2qp369OgP88uU05Tp8rPgx/62IyHZiAdPshHwyx0lRJhRWSCCYs
nkA+0UEJp58Yptj9Vjhno06mDHXWx51Az+ArZp1xBlQARpnV+gw0nMhM/6L0g6cy
OfF58F6ApFcTKvAWVpSmvmM2cUwupZ+I8Nn2RgAGBuWiHI7Z3IfwHzcZ+1/54sHQ
i4FFzRrNM3G0Nx8lfCKMLt1HOKMnKn/3b+GAXyv4lNnD8YShHgASej/hWAOfp9t3
a8Mm3Y/PYJcgNg34zLA+auCYw+o2ysqfN/tjgyODdqYOH1pBuxBZAjcfyOIe4MiB
G3N05H1IVo41EtsxdFtRiiT9YQX6MHjULdcdBiZjBsl0xY0T6QfSpSWZ2cIU3SfE
aWgh+iJvl8jW+pKFPhguZ+H3Oq+uJvZQCTAxnMC8jE/QgB6Jet4EjpwzPXyQ6Vbl
zhGcaNm9DRGdgP8/2j5DSr5wzUtMPsCr8xY83sVEEebTV4SlMhZ4jOJBpreBmAWq
IS/OB+KeP6W1G9rkh+Gz5N+Z5AuZgb4EICs0tRihmoFurb0U/HWj9mKXyiSeX625
NlPupTQG3Phy1FOkZg/5b20jw0SEfeAydeuUSxnUKpHcs1pxNShr7Cf2X3hyqbbe
nK4OB7ZIpIxHyw51beMStWoy6urvYkNfoJh8lfdUTwejm2VrdgypEP7mA3R7trm4
NZyM/F1EGC2hVCUKsfvB7gNvBmDLHBXWT9W4VAeKW/TBmbzS2OPEE8bGKKpJmgjj
4K+fwrF+un+erT9L/8mUHDgqE/eVUDLh0VtMgxQQorKyplHmEKQAzYKwz12lrKTl
rBZ9bHyttMmJEqOqHTTf30bkmvW//136IhqIwsaR++KIvH2CLU/yqkG/0Ntwigpo
`protect END_PROTECTED
