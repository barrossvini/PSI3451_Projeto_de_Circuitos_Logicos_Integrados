`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tOc8vt38P+ORKRQqSkHkjDQ/qSD/2ZxGMrroV7duRbmEwN058zgtVnD5JPKN8n5s
Mg00GBiFVcmYl2sBxVpeUlqoX0HNtZuxkwp8kKb/XJjBVLOlB6QkOYGXpVTGhpsi
Dm5OzioOQ3DOvslIy79IWvSKkq+JHVAE0Lf3NUbi0/Y3+kmFQGumT6KVlyIlzQED
V2K3QAvkk6UGiXxTLhHMxiYDJa3s7b/kZae7p5MbiLVX9V60/aULw9yrP+1vxN7C
00Y6PV6fGECjm8T91dscwv99BakI9o+TCucPX4nfWTqM092KrCabOkgNkbv6OG/m
ReDTcPEOvL5KBei2ao10/PMvxksdblXTFxUybWvO6FeiyGSPqhMrLabdboMJGZau
xQGBSGhJ764EuQ1CjQlOxqi7HuwLvuguq7kV4uEsF7I272Ig6IwcwRRxWzJKka9+
CuJvgj0cTpCOC1pVEHcY+IfaZkfcqhh5QM1padhjgtklAlQ2dBwY4gS/Eb/0X9Zt
mC0+oEWLYVZwxgfergefp5aL/S8ytNwwxfsTz51DafF6E+dSbL3GGlj/vYS1Wjwe
Bnuw2DMnxW0TOO4L5CR/9AdAGp3ifnbYo74z2KiDjGJNRcSrIM5mqgf+MeSXk+OP
7IsEi1dauP53l6qeKiRJ7G6OpISyIugwYo+kK32Nja5ji5tQWSG/K44BROL5fO/I
5X5M93sZkTxczUseJ9kjmEvGqTDyNZDNfmuj6TUjS/0AuPi1P2iwjhVcgcEymbgR
Z/+aSrk0+qtzcegz0c9xevcFCX7FajWB5vND9QoIuGRrYEynIyOEsR0B6nYsXDwQ
iycOaa+bk8rUS/WovJpuRwsej4vsMAxgRBgESufN2lG0DHblx/yQhksATTgbFEJz
osz4xfbh/IcjaMen/Zmy7L6k8bE66wuTtt6iQgrzyG85QkoKJWGDUU0FXCLffzLH
3ispXi2qtcxg2Uh+sYHdIZ+z2p9NdLwUSTtHjGYLNC6YkgJQZe11GsaWrZo23fiq
S7isAUwskDQPgcG4WieLTx7qN38iff/JHcMRCG/8HSuNIo9N0ny3Mwddk9BVF0QP
OprQooCjhtOtkUVa+KW9M3Z6X2iMEq5/beK7xFKhID8MzxiF21zJD+dQICXC5VbM
SvT2Z+jvTug+YzC0S/SpKelzendqj10+DgL7uIG5/0yjRJwaXD7/h+SPIIWQHckj
druYkUKZch9YjhMk2MB3+mPyJwhU75uHEQLzGDPmG71VRgI/zaFitjW3aX1ktGJk
IO3nWmxF6Rp+nHoNeyKLlH+UeV1gjSsRVf7GEzJQCTgIRwIHnPxsqnwivPP5Dj4C
HSlxq4LPVr0kZnhfmdlvNBadKOoOBf6UN0ukewetkvYn5qSCBFCRnpKJbgIuZFv9
Q9DPU8kdVcOLveIVE1/Mk5NgjT9yzZOZHdhXwWlna4REKWP4DZ/T6rUEc0EbAM9X
nnQHGU6r8gW+2u3f0pw6jupfhXd8YSlNo2d7iZAAUJIs36HfD2sxStG0rW+ZUPqC
QdF9qUnUNfZH1/INsenwRZwdOFPft13iogu1YC9E7A5kGiwkAzAoBwlo76NvTpTH
1soVZp5ihrX3UgtaX6Hl+Kbd3f4ttZbnyrl4yUVv2qGOkzigM1ksYt2lTnmo/WCy
`protect END_PROTECTED
