`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vCMyDULOziuL+dQk1Sa1gAMQ3G4NcVplmzVeTC3k2E4BIZ90fNX3BVEYiO2hsJli
xa3q7PcIeV/UxS/afglrgz+lT2aLEI0EdQCpU6QAf1GgP++u+0JYGuvIBU/AMjqe
JfxyV6RkDzawC2c8QvwhLBm/nx8WTOAPbupkLDPHJjcXeyt2enZgAfadRvaoZLoD
zu8mtpo4xUvZCPaFVXcRDqQLQYINGbGPz1AGIs+FGmEi/iCRtf5j84qRVCD9bgE6
lwsvJedIiTOCmaDebBXASiP2KsIwkxfw78siUPT4qfNIC87ttuTqKi4RXkO9Tguw
IsED1ijnLfIAvnuVkmn7J+legZb+Rsr4+d2AVbzPWTSfpYKwmdO5sfzwwBfcQvT7
YgjT4V6gg5Okw8P1LCClLxLhS1SqjVxzRWgW/2ivtnHkXf9qcQ0r+j3xMbJQpN4k
MYCTu8hF67z3s7eVco7qCz3JOOUfSrALr34ZiUfgZVEYSwluzuGz4ypj7SctkiiB
pJO5/M0vIh5EobKGDYvZTj2HC9g6eVr/hHaMkzRMtmOu5HXFu98fz9UBRUbVPux3
ltwrwQ9r9YZMazwS+y3Zm0NJUrlAwqypl12pfcfzmx7oVHTPIYr+dp+2C1hAkq7i
PeOK6falwMbS18hsDIkD/gAjf0Ku42PeOWaKdkpgu5tCzFGPdZDvtT/NcLrXjD6r
YXY396UgM6toV8Lbd2sm9OTHVTXcWofhNpQbiD5sPcdNbpnouAKKJyxks8F61+Z/
lA+n0rua6cnx0a6+9ItReMY1YKeZuAo1KXMWmP3iqpjyBNmMfl6i3lkuc9ABqctY
3kMWNepi51vUvpczM7+HgMtYuti3W4TsbZDq6MeHx1A+znrr1qb1d1WLIphvdfHP
oKZDBGDXOTXmW0R2HvQu4NrR0d8Sr3W6deK1p3WgUaI=
`protect END_PROTECTED
