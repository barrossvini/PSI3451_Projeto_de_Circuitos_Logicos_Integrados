`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6yHow570hohFkuQ87DHN951QJi554j+6ZLf+7oD1PJs9leraURw6l9sEc5AQkp18
gGyxRl7opdE5VCSwdf4LpxsyZDwxuKR1DeF/ESY271sOrN8cqhzzZ0wbhkLOuHDB
DtATb4IwBM6otvqF2JZzAoKetb1t2OFgykxEHWkW/isGW6HsTh6YaoKB/DMKfooq
4tQlFY9kzvMlKW+KxWBVnCNwM49SyJo1VyKkEPZ5POiE2aiBc+PVlsu3Pnc0Lxzu
2+h1rtmSq131ME0BikcXSs3BHts7uw9myrt8po606XPUlFnrnEVwrleMU/LX2nmI
SXrTmTW5UCscjY7lGUVEuwKXI2ulO1FeCPBO901XfTAQKS/3/lg965ZRWR4z2C4u
NOs7iQHdg8VxVffr+kbbBol9oKrGCThk1wLWuswPH+stTXT1/ZhO6BZD8vx80ZyZ
ZQyGgTq5TYRzNrZIdK79K7tdQoNnVKEJVsxxIhjMr+Aa71Z9vpmxwgmAGfUcvTJA
36luX8E+pOvTd4D7f7N3CDwX5NfKS+mMhETGnRzmj5c91TG42XXwg+fbYayp6pJR
TVJawG9ImVLGzXNRLUJ4qKEWdZU68hGZWYXjo69csF+emL1qspNdT3Jyl9C5oEV+
HJ8GZWVbv69L+gDT6E92qs+2TWN+mwdTmAwjkE7w/JAzG1s0rfTkjUjJurze9SNM
MCktLNSqX2KnPusfB5sMAtbjOJ9Fmz8QppeIoiX04SNle4/ay6iPKjr/cEhWy146
yX30ibKC3bC5IlHMZDWBduR4DlKDfK4bNBFb+O0jRotqZ3+gtgAKX1o59SEUkSJr
vdsU/qpeMy4pcBmau67LZ453dw7YUE28cJUBVxywHOxMvsrax3Gk0rfi8O0cKPK0
nH1M2+9gFJvvtTkdPCm4Zo0CCUjirwwINAdarD24u9Xae+9q/5cxgwoJ6Kc2Ro8g
3Ql8UYKSA5FDKh4Yp8qfRFghCQPCV1L3QyehWEIbzeOi30MszkBTpcEt8msMveLI
cEG+3f1049GYKrzUTMasgsRQKqBQ34f15JhQeXQV9zvejgUp/ojtIBBC0NrxobSo
MvaL5aXhU2x9AxNCaW7fFW+Nn6RlT2sjV0mh9cWuYpd4GUy/RpXs8Bw6a3h041E6
u2xVRBVJMtYw6xB5EX5Sk3BeufZRQtnKIdBHL1hQN1hcz3X+Dy+U6AZpwljagCWV
y8vQD9tgSNVc+iS1JVsTJvU02522EDVt35Uo2GjFOhSyYsmShhvleKWEqC1XZ48k
CxuuQLyD/4kdE3Mz7dG/gwkMLow422JVka2elEhwWk8hV/TKlxHT3n84p/3IXSx4
5gXdyyvuiBl6jCrYGO66ijwHYLrs48YtfDRjkg/nbZevkcYNVuZgdWC+eV2MhfRS
ApLBuaItetxbFOqTMcSy0W5dzMjEH6Csf1zDLA4fAuW/jY9hjRlI4/UOsemZEDwX
itBLm9QvFY3+3Oc/Bn2TvnWWOU6kXWqV1Ewkc797Zr/CtJvFV7t7z4AkdMVQpKfM
uvcs9GJNzyXjQCQGEICXQOf0lem/7lgjOc9XMUoiQI2R/bV5EDSsgmENjUfnQ249
tgC0roS1bxT/yPl02FRcZw==
`protect END_PROTECTED
