`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSQzXl0A/+1IjQ5goeJCCJKhBtWtUNQiu2NpEAt1n8pW9Nw3wEnM1JJ9p+NHHKpS
tp9RprV0tH8qGMl60ZWtycg28ojV2mFQSX4UdJmw0vTPlNdgqdeulLxy0TfuEL67
k14B5tar1Aha1SRKGq1h2XQfep89xkI3xC54g6HibGXC2uMa6FHH1virrBfyzCnk
T0we3VYlJED/5zYj2qvljEOng7tgoGSkEabWzBNSSkrpBS3ET6ItdxH8FU3csg3S
xYJDOvlqZbhA91jrSkZ+Up2rNSwmAaEAuQHGL12c2nA7uDHv3T1XL+FMEfGP885V
zWbIbqc2KH41CDgV9XB1FimnpEosvRTFUkU/FLdqd2UhU+GFR5GV45eRIjEXKjBL
PM228AYeiRzspXBC4fdzKO55chpxDfGCQwe3RutY14nUqt9iO9kbtSLSa902fNPF
U0i8YB0r+CyUxFNq4/sfwgwfODMdzP5La40n5UCc92TgnD8X4mYUYd+Rq75Ke4eY
PSJ3cl0x/rzJj4EwyeKWTX/aXXikmewcSgO7t2f4GBXG7p/5jyU90uY5qXCzc933
`protect END_PROTECTED
