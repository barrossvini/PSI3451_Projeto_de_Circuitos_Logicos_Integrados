`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cvj9xR8xxY9P6cre/ZxQFEN5sADOKwENANCB0i9JxuNYAFwHRitbJOyc1CKYcpru
W9l8N1AWmw5CkcBp7LvuXixcfVH0SbL6K5iiY3jJLmQLYUIWxNcGXQJt6P8pMfgp
660C5AbORXZXnvn6kn3UEHxqR5TclCuqCqRfyOU/1QPIYoWH0LoNbC2c8xc+GZnq
oi4LVuSVZJFPk3Gl5uwT5iUxjDVE6U/uPF1LNomjFhSNwv6Kai3TBUAg2D0SkpPg
7B7inOOQW2eUg2lqcwwEsfOD6eQpJqXOUpJzM6JIRT1HUoZu3kLmNa4ETzHcNcNI
w+rN8FnbUA48zhCxhipyFPy19E9QUD//SnLuKOs25md3CJ9O9uNWoizBFATmBHOo
ZWZLNe8lY6ejdyS9RJkRBW+Ta+YTrz8sf2GD4nT26P4ucfydsQMze6Sj207hW5aT
qOiRF8NaoGv7NnDHxqItGnuJiY4PNaNvIQ2FSXDTPAT/s3DfV6lP+PJn1P4373YU
Va/aSi2xjl1lKGnyvU9H0Gp5qeycMtkt4uioByKt48DH3yxkpGKBoNwGFDv0HjOI
I69zhhb9RRgUQkw12JqBLLhCKVVi3ixXThacSFyJmslhsQlZErmcHoyWvc1dmgPZ
XLylTv0K9jcJ2ob7EE3bit9d2dNxmMVrJVPiRDhGfr0IxFY42W8sbAXR1s1xPfsq
LaaLvvoOf5JlENyMSeywqAdmq/WbpmMaRU5foFes9bcWGTUpiuSITMUENrTXFICg
QOVKLIB5qBA0/xgvW+OGn2jKzgIukhEzFAcCwzxsJmnb65d4oZ8vCiMgPx+d8NBO
zaPiEAjr7tqAouH9RpAL0OsNUkOkg5f8IvmJl++CFR9EfBKEowD5BEdLf1AGKMZP
+ePS4sWX1qf0N/z5oM3qeAOr+LNerKXyZaWfhkyI+n6EREhTU6aCmfWU0RmCACZw
sJtmWmkQZsTcXZZdK78FCVgzGJ5oxxOmUx7Wl5BmnPSalHc66+yklsslR9o1h2Q+
2halhk4mko9NdvCh4c8GNJ+yp1gDF8i7crthUaKvSvtPcq9LX3yVtWNRsrR+udFe
VWpa5AnHGOrhIgSZIE/LFIN991j7d1lEm+cENycZNqZIesY9+1+lUpz6EuQyuZSO
krwwAlb6H+G99OFks16ISm5KCFmZnAka8AHx8I9o1a4V17vbApb0TK9/Ut0WNfWB
qYGtiLOMcHv9gXwkmHbc7g/kIpCd7KyyePBdbwyQkAItc6IyrqzqKdqma46uwsEM
01xJwausbdWy9ExXDkpuWygjGH+IDY+t1PxoE5t9qNElv2+HXmTtLdcFVX5XkQ41
eFdK76Ss4DTA+4JIg9We5CsmgnYD5Fcrky8SfUP6WZ+jro8y5ZjO2NkF21StPvZ7
1H1OhMNto5bt4twc9YBPMCR45eyLob344TyFBda5g+V8ErldZu8pZ3jwZNS3GnSg
ebGSSVYno6Qes4mnnXgLCwamQ4Uq0OhreXetmNbUQbge7Yf0CwugExWNiTjN+fsf
HRPiFHSUELMyZSujeBhzb5eD5Qy216stY/4uqwnlipiHwOLddB8vJRLRVfYcLVLR
DyLakVEmwKXMUNPij9lygEQyHH4ZY8jslviESSwjqIkFajV93oI5pLtsVDCOoo+V
cXYWgSy3B+ORGIQA7u8J4FG7zqCiWtryZn6K+Uq8eDLPwwEUzkn1GrXcVcSyxqIS
pz12l66Gyf2ah8GS0hRQOdJj05bLxSN5KIEoYRJLONaYPY5o/K64wS0bDWjXc6Om
6hiVPygcZKAkN6LAAZ4jyrqefkTtrue2K0DnaceTUpRXiNJdt4+Q56SpxaeBhdiV
7cNPOPkFX1Zkpmo2qHbChW5dKZxoBfTIpFDAWEWbhJ1pkrQ7CkWvKvr7qgkZiZX2
CZcaO03u12hxAxmkyJp1YXvksoTynwIsraMmaDnfJPAVFjTJSQy0QI+pfkqwtDfP
I6tgowTAZlsNFd2ycxfpIl2s3z5GKU2f4Gcrddp6eTpgnLjCTgPj7FAqF7lgn5hr
3cf9hxnk8dbahDlGY9WZvJy5/3/w3oRKbMnbbnKSSAp97Hca4Y9FkktTTwPiBvxO
00/DZz2ozl6q6njdZ+qAZQAMCyow9KZr8vjiTKB4OeLYLilxi5C28oLql9GoEdUB
ZJIZiJ8T7E8U5PSEspZODs/dOwE+HiWlr/SzOPTr04mATSJsn4EBa1m1YPDYBybs
U7ro61PuZ7qwn8Y2yl6fBdnzomQws1BLT8pqtpuisJ2z/CBm2VnIUZb3dowDKb5X
U1HbvZGrh0SRVxrRRRDAMW1vcqwnrQPUy+XKJI4HiEKUMiaJlHyQO7m3bv/+c56w
GRJJt0SWkYgRv4ja8YKejeD+Fu7UQuPoBdupepwrrv44piCbo0GYVXLwofUpIKXt
+xkmeaG9nfjZI+21e8SY+yGV4p+VfSr1+vFJdLbJ8wVK0HM3XCGfplbueBO3pXBx
ucvaQzRQVsp3Q0864r++PAWe57+GiN2dvhSMMKyJZw2oyLXtvQHHNgsZLDg0Kq4e
stMH1UsQVvp7WyERN/F0VOhUXF7cdZdJCwmsqL3oOY/8EZ5LVLBXkiNrEc+8i1xm
QkBpTv3tjHYQ6g75uAnzrr6TFbvM1WNcZ1MjdN06mwxzIW4LsN3tsnn8bZg5V4lm
9UGX/5UxfFSEpOCHhDM0OHyeaSnIvyFFzxBgg3QkijZlDG/y4BlbaZ9bHw0cgPjg
GyD50VJ1Hz3MxjBDzUMyBQR9SLjmSQwuwgI3jbh5DNdlADU4uy4zB7lPKNEXRgW7
B9Z9SGgowOfbXMY7GiohPQZxDiQncGhiv9dlQhvF37G6rJTGgKUOpXkXnZdOfbTC
ESGN5h98tPOYhEM7Va/gRcufYmsbPt85OV1SabuKbXPBFEy1DSuINsOQEiwQ7zDw
iFA6BKsMWzo1a+N5jl0Om+UPu5SUREzY+61kc+I4FmqLmlPsCcq48XyomHajnXlB
ZD70nVlX4bvlpj7qKZltVpW0nnDkJVo1FlomqRXWxIEhwOhN/T5sjPq/WDRtkXrM
nVdRkDaAKjuA1Hcv3jYbPFIwxiaDxJ4gbnxTRqo0MIGsDbKge5wOs8obOiRerhQB
J/bPkExnRvvVvKensazYAsVGap6opyRpT0uB33JR8+EbaC8VKaviJEFvZLMwzOJ1
6kUdvq+TWgoryK0hQI6It852yeuD1Bc5UY8IkTi14rEyFD5sOxNQlI1GHpkzNvTM
9EyFsghDd9o13sqU/lbgfxyXcKQG416xjgZTspm+k6IvU7Z+3yrS3FKQHAnb//4t
fwiQW2pp55PQeG8gOO7GPvfjlQ7Wfhnrdoj1ThIVFr7BzlQX590tHspgif3WFzOy
lEnKYNk8o49uQmJStn1sghoI0dl8I8z7DqDUix9z6G03WdU/qgNK2EYr0BTSIkLu
SohNUpF+nfjDMT++QYOo2gHgkUjPAOFENZJfyw9kH8xkKgPklYUIrcMj8nR3wbw+
//98BUw1kGVweH7pilvlsIpyHdxFhKrrn9iWmTZPKUC9lcB6u2qMl/EeRXLxIjJN
WCE74HsQSWkPbhHNXROQpxTq6cU3DXeempOSwF9LBGrfUdihJ/vgi2h1MCqG/DIe
/UEwLdGo12/PJ9QEPA2OmttFtBXSMkD7WWnJnr4mKtrY+j5xcAV29uiKr4TJaIav
+40YgYWeIicLAK4MO6OsTTTmLTtcT+gRDSF4Q+hTsVjoH34IbkuRZZkwJ3WfN41/
2FBfxvvfghvnGrVrxLswMiikqHgAYk4IrHHVKMlIthRR0JW32lg3S+hFubKLIp28
0BDAUBoKEMRo9anyqRr9JJyPgZ4V1oWhcjFODcM2oNDNRyV/c3Pu0YMaWcqV7Zo9
VxFhN+VOp54aLWY8bbqkqlmb8giYpJc/mYBtTq4p7X1d7/eL+MP04U/GnyhibmWL
zncC0K74zD1uk7104K80wGIc3QfP0lix5na1A4eXeB47Ug/uNBMFKqrebJqhcptR
XKSwgLTvTCteeTVrMAqm68nyqNVVfust+ZdVBw0GKnNv3zJSXVp8ESxSDKcRX6ek
ox7V1ouwu4/19FuLqQ4cJHdVaQug6/D7j7+3eV9IS1SkS5cNAeW8me9fetuWqCck
CiYH8I6XdrtIHFPdBtedVVYAORShpabiBokzJEn4kgFlAHf/BFCkM+JkW3OvhKPh
+Bc9d3nvD2aXp6LhSCn3oR2SkLvONkFzuZltyUXH9KKMDYxax+LUabt9vBWI3Vcf
Y2TvuoqynrnuDULHzTqdDwyIuzMrCKUCokjXq+y256Zpx3Bmc4OlN+sxKRRmxItR
H5J6tk5qGRqPOpaOHimyTtrZUiLhIz9ZsoppLkazjUVjfCLzFIBwQyxgE1ORMZ5D
VbLF8jx6cIgc3OyvsT2tmGyS0vIc1eT/McijneU92gPYxnLk69RjKGergfSRZZ8W
NGpRBkXEbIPBi1wEsnosu987HndPS1GEhlXkx/S/Tohu7Q/ODCb9O1nAesF/eGZC
DCOLf30MXNVro3yB+bk3LOdtEfAw6EUtQN/OzcmceljGrF4+dp7E6qYFNnWd9UH7
YP8+gLZfYs/TAF97owm1UteMHTxfxDOY3lZ0eTKVdnPpW2SJ5ByUrxAlzFpe2sfb
9I/+6LTniGitUorz6gI7pptlAiOZ+zy/6GRrpNuS9qCnDxkY6l0I4qdNidX5icEn
tsgR8PVkcvCBpG4Q4Kkqxu/WOHm3TdTs0Hegetl1VzpOGPPTbEA9+Con6WXqNsvw
`protect END_PROTECTED
