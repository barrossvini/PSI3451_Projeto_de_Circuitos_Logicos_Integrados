`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iTWzhS5UmyB1W3jEZwVb5xCDUSkW9SmoOAJi6Y6e1QOCLeo1CgnKMCTstO5Sma+s
Y/wOOnJUKvEh3YAAdDAUDYbRdniI7uaYCqo50DkEFjuEiAZCZmIYJTrupSE6C4zE
mAJwSDnn1RGnacG19Pl+ls0E2qIY0vBI5nr1o38uuIQupMJc8Oq+cTd2en6CD2WO
lp5QbCMEVSncw/48+MUjKRobiBWULSI4B0D9B1453iRCIKPJOLGqDmV8676QjHiS
yVUyaTt/tI+Bqxe9TMxZTIXO+SpxhSRFQhCsedYmf6bJbtsh3myg5JQJtCnO8ozJ
ttiLh4QvVIzi/GKmRcwrXF+/sIJ6asqoNwX5osaIMWlz+U7JfaW/f0TwHjh6maKv
UO+jqjvjPMw8alYKZwdk7R3cvQPNe7q0qEFk4ynpPDpD/q5BtXkdEMbxlDBapyqv
6vuKkkvH1IkGXeKhnCMiYknGi5eyXmNH4NmuqDgsitOFw4XV+RGy/BKccHZWo4BI
+BdUtqbWpn+90Ej4F9C2opnKigZiSWhxc1CV585f6wNw+1147kU/j31z4CiJvlI/
m5Pdbiz04DRNajvm2ynZqDrWnTDeUleAtqtoK+0wPgLqzeMkkAAvtlIdTEsG6Nnv
eBR6vAXie59PCCtDh8hH/MZzRUI9xfUsMTms0IW7vxupshWymc2l0z865yGF5cuR
IST5GvSh6gkdlJldoHafOZ7tPq6X6BKv63dvn3NT0t/Zl0s3UEm16PhUySdH0b9w
BXVyoBB1IU8f8Ty+Q4De2UusU4EBeQD1m/ZUgLyWyDb5D9mZKpveLVqNBBpqattG
vIA6wYGWMS+HiqI7c9PB4KR0hZueJsMZzpXKbK17PyQSfzJrGPijvEeb/hIbnweM
19BAQPbcUuOXQF+jfdSTy7G6RWUWu3IFplh+DfpHOXp0GyVEyAwYEh9D/i5oJnaX
49cZE73QABI2tHBvV1S37tIO329g5P8Kvh9hrbT+IC6RQscUJiEKAqbKqrKUZcA/
ITlc0jzsms0Zt9/GkK+j/fSKgc1JCligbfL+iYym7zqSOeuw5EXsfkIsYVv4UPsP
t48eHekRLjdYJbpeeX5COrd1ppTJ7Q/f4sT4ZLZaWnIOr0jOxqb4T+PEsV9Emm5O
ElGrg7NqZcWetV5SifceAfHlMY0vANIgo6zUcQDrMEQUaB2N2T731b00voYYAphl
q9Hqnen8k67tmvTtcpVYVlE7FBwGeur8srsYNNqgUeX3p6B4mCNrsp6VXyzGcDAv
UWGm2/O115xGEc4xWcjND2T1OACd+bsE6Fgw1PnIVyVQ3USXnFDJ4jbIqQiriics
SHzVvnFDMKqHsPys7JmfrRDLrILfDMcm1s2LZpLKqFUyh9cG8HmDksumbW6TY5Th
E6/EQVGzrA94+DFwMdXw8Nl3295R0Sar1WIgBI+RQ/AYYtFkbhp9s/2W/US21ees
+h7Y9aSVop1dzR2mi0BGIUWveQtuCbZxQyQAx5xCdkhDMZXFSZUYLiRNVIZlHiAV
5hBn7LsSwoHrSYS/WEuxk+Bpbw+mjdWH4KZD3ekzk4ANKPtdbltXUzAcEV0V8A52
t0jihH0ms1qm+k3P6YXO4ZThDQUgj+coWfqQP1thd+bXpTB3wGzQhXw+2tq61vP1
XZ5Akblu46Z0LKvcsfxPirGbWTIZImW6DT6R1PK8NzQcvc2qmmSLlW7E/qn4X8Vm
xNhO83UHL4FJ+Cr7Cw7jOW4SADID22wLeZd6ISqy+1qod4w72D2sIIfnFM64ThT/
fP4jeW5bN7IVSCg8F5eO9ag8+WBoOCVgbPqc9jmjU54yKVcB3uNsP2XZQWAPrNa3
Ov6EdP+nYlk9djlJ6D5jVueY3ObLuedCh3pouijMpeGH0dtRqJoWN56qqpW/RnRG
C7UTH0hP3C+HsnhS7HuADTBdJKZQ3j3Wv+V128YcK7ZhOkpMYRgVPlapEU7O0k2d
05tuD7dGCRK31p6bp3YsEt07Jzddq2158eZspZmQOYWH1HHxbx/PSo9IifQgKqZJ
6CSFVVU8vx/qN5uf5/R9iqK22E9b4Iaqc3Vh9XdmCRbGmBxUeXvlkAMqj6UoCeDY
f3b3c7x65MLjsBJz+u8QLBzLDkzeY75YKPX9azwC3+/uodOHiASeSqSjqgHuZQyG
OQ1Mki2wwHuIrUGYrsH515fhj/S0k8IthM1VWWmc5fMxPyFmyS3cliQHjxLnY6oW
I7/cMofoNp6xeXGrneWtsp9065V2qMSLzy/K3ShioKByl4+IIaVYWDQc0DVJcF7f
rdaMwIRmGcwVJUjJJrK8wSRuzNHE3sz81Dk5Ya7rlqZ6aMPHYP2tMLQdpKi1t1X5
rLFwJSC70rItwK3xRyJkyfOS/8W1Hvdy1zWeD6jrKGu026tqp7tYAogWzXB48wJp
d5bK35tC1c3tUcAb2IW7Z2EuC7oFLsL7bhjfy1JQWAdy+E86h7Ida0ql1OZBaoqn
UOaU48LvIY88vNN8cEukf7oriPnMf7gjb7/nP0sebpGLPv0JdOX4MSEYjDdwd3q5
wrAJQVsm3xQUCX8oqQaY7rO0P8L/+JrN5fUBW2Xvtcod7krSuiViuKxPtfTFnBaD
JRBOLnhB2z1aXfwDvLRrZMlzXXaDzOBGOV6xlpIJb6yXgJEWkbxiQMG87sY0APSg
VgsdTsnC8wK4R8uaRrCuPE042Z7ZlmsODwERqEDBSg0mTgOTpCXATzuc2dahkshW
ge0valQsS0r/2wtyMh2kaqmATbnZLzpP6GudkuhSe1yP9ja+jUaCUlOgBM9T96qs
WGfxk+VSuz73Y0qRhlChJaWHNhiFGkXnppXrw3Zu08zZ6I9tPBl+UIx9P0Gpr8ak
MlF1CUCqz4mfHKy8+rOWi3YiMfvewG7FKvF0KvHnHr+LLttRv4EU+BXsuSq5Nysv
VIm4LCLnqruiXEydMV/ziSRIrFQYC7bxX56moEN3QALJuYQQwfXWGGYZ52OnY3+C
dWx0f4VM2o0PTohHLnZMGGYKhsGXc++OxiwTNg407inVOciA5aocN8TB6fHvzFYy
KK6RAE52uWAs2/8/xRLUxmSiBDhyLmaG8oA7YAP1q3vUf23Etx1Vx7S4RHzqUElQ
2ho4fNsHkcCfdzpjXVyhJXGcJbgycKFiNnvGPESHjbU392/I3VnxU7Z0RoRvo3Rw
cJZlvEg/jfV77ois+6fqdgczVH1EIvmqENw/+cdOfs5rZUiiF0/mvd8js99en5qh
0vlWSn35yE1B3wCJyNUZzvrUg+e43rDd4FfljxVzg/rAUwK3kKUUy8uFDaQZxaUF
x9fvZwFreJQ59S6V8LSa5iTvdDRrHLEw1O1j6hDdqMza664i6qezuqM3wMV79QxN
fuvRC995OCyzr2soZsaIaRpLarKSBTAibFGQh/4B7vstNlXfzzlu5bkAjNbAiTAu
9s3ArBBs9mx2VczvaRb2c4hlQlzNe7fi4cxhTSiC7bAQtsUfFByC3FDwHenllMgn
N3ZDGRKl0nS95ZPbu/nBafcOOBAg5w3H+GNJdMa6z7pcGxSwZcGARk9CtHGv8KmX
s/s+hN2KMEW1/yjODHkyDhGk5fnp+24imO5BcVjFW/YHLLFsNlwoNhwmkVG3Jww0
tHpjUKEPMt1A+CV9B5l+T9sDbbHYl3IR/ixs5GAB4Ce4Ga0wm+UIVWOvA5DJOhdT
9EQaoSLLgcceb7eSSsloouseo+MbXRpNoV4k7TYSjpP/1AZzuzgi1oBAQxdDHnmc
GH/4bKTAGeBY1Y7RajUg4qSJaG48AxtqG6+EpLh/AumfnFgy3UzPbTaM2a+WVp4z
As7HGml0vZQ7Apt02jfpdP0EoHz/luZb8focKdDEwS/Ygfmqm0srvMZIzW+F2OBB
VjwCZD7W+BENjGRVWs/IKVei6/o+5r3pm1n0OCk7UgxfK/v7t0xBDYbH8ttVEl+n
vJ36AYzTVcRebHB0LxXRQ2uxb6CzLpAPG6GqfCIHWqjDngvr4r+8hsjkKC8qSDwI
mAR5bIfETizqHa727Fy2C+ZErjGFF3wBTt9wWzrTUdLZCyKuzAJ9OpuXLzhJv/Fd
LD6G5NMaJsosp4ISX9BegyZ9d07hHhCeyBYn2yLEly+lA9ZFZ2AswKRo+COxKIsk
92ZErY+DXG+utEqaJQcdoe0GYZB1w5I3gjjZeUB3CZZaGlQurVrIeIzC9/pwd3hn
e3NiOu8kKoth7mmxTxBHC86O/pLUWYnjn5koS+RzYofd/yxdgDY1gLUV+fvidiW6
maqTzvlCy3qx2EcOrh+QDMFBoY7PodcCXuLiuDGQXhKWp6DEqfalnEbYv7ZYzvz4
8wRH0qcY6dxwgdtq493VJHADi6OpXTbabYL8kFSU/nNLhKexSqAsvzn/3MV11NNV
eD1lJqv+vjKAKscLesjEUwmAUGC3FavR0yh0uNhLh2mexrWDJuxVROgkSH39BxnN
oD3sgaqfPQzDoOZgYRWC7kZKK4KGZK0MezftSrX4DpCtcE58O46HmW9JRlehqM1z
xMjpSZm/NN3ruULRN9Wp3uNZ64Buv0T/1HhZb2iQIoyGOAYKEzBt0GReWA19KIdU
`protect END_PROTECTED
