`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H4D6BplG37NaQNSLt5Ef3abT7AIIC9cNbGGaD7/iI8rC/siSMmwEiZzz88EQudqg
m8WtQpxq+Tvs+IfGdzIwdvWcSL1CoNszw1tlw4KLAFCI8NGtOWP4l/zF7Qq7JmIx
EpOt1iMvjRUru+cLLRHJgNHudmYiLW/JzLtZzzT3lQi4um9kDvx7BkiJ/PaKMno5
zyof2a5P/oR4cv7JJDRZ4xMp/nJopIo75iMGbW0VZ75kDFSc81bT8pK4GfoqU2uU
yXWciX4VjzN4fPHuYoDTOH5UHfex70E8XqPd9NMw/W6K/se4Ah9UY1/Hrts8D/r9
TwB11ADJWCwaaTPHZzmPuL5f/lXxTmoh/9Qol7iwp93iHO1lvjspUWTwSVE3Ucu4
0kpYHdiAv88r33skNpmQ0hWGzUIWCgbfoi+fC7+LAT/twT4aC2Jltb0U5CW7UOGp
SfEn8YSJmDEknv6RH3ZOyF+UO2aYCOYHa3/ZO3HGDthkIHw53auMnfrht8bF/eeu
SCEyC0PhunS21m97P9RWKBhY7Y0JHmICDyhtpdrUXAHCR+0NoXjaxtJUywaOHCTO
H9M0GCSUN4eaG1pYgpnekTVbQj5EQPBr161ZPLkX6a+jnj1IoB6EwasclPL2Lllv
XVcZCvoEAu74RvtMpVTxC7QJY2X0reIhydEF/6PItoNVL/Q5bLETHOmGk9opGIrj
J8WHfdnHvnmRtoVW7QivQniLRZgMKzNYfR5t808etCFWBKp0M+Rw1TAVAmMKFfj7
TsYMXspygqELZ6M3GVFBvJUZKSBU9ttxsikA3ZHKPKNTfsiMVsVWl4Ljdd12kCx5
32I1uQzAhjDokyMeqhTa06FFpMpEuHRNBXOxHODkAnVyHLuAN5S7YjPkYd4hBh5c
wL+cC0lY1MlfFTvz+itLso9mw8/3hHObpcn8BKRHskkeGboUQIRruLDwwFxe62mD
DOZ8B/bNoMdRci9c+Q/76xgRTGb9LNjtRLvrh5xalxeaozlXaRjNC1/Y5btIlt0K
2Cdh6wd9g76WlEqdHPNaTWHzr6ueVsQGJMYgvilflGR4QTXY4jwEoHZyUqqlV+v1
qM6Yp1LYHIaOOhFIVglLXITp4nsWqRbE4djE2Pq4BbH6CwkoUMkYYWhJ8BCLpMt8
sMlxj4wpWyjx3Ju0jnFu6YF2aZ2n4UlkdzYCXvn1G1HWNZ3dYg4EKnAnQGF9ie5m
2GfIx7QMX4zsi2m76P1aAeozNapsdX+L9PiCkofmAy0=
`protect END_PROTECTED
