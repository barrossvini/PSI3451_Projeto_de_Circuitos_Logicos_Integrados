`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UK/QMtGOco66/cE6bre0bgCNbP2r7fOSu5hnJePeV3eIUrBiN2Ywxykzd+xZ4wm/
CuKUZAvPpYLEdktV0vq8kOklpSymAZTDVZ3kQ6ZCX6KN2mPLpaHakBWhK3R+X22+
DACrsmZ+Y3x2wM5xoGMsmmREfGqYygWpPD5iofVsBtHmD6uxfZsx7q2HlsgG7/43
Vb8z1LYuiPjCMYYl7V2uTNSyMDqK9dlC9nv++AZnp3qqy3xbJCe2ioNyyfmWZ1oP
2kX7qUyV29HKRJ498mcwX37ztgNqBP5V/tGk2gmO7vrgbSnmd6NgqZZmFTZ1nZMk
y7Z94LIRPHaV2OairMH8iaAxSBI07SxWcQZmdAftnBDbR2lSPJlw51J0rYHaVwoE
WsXEjBvMYNrCmpNWBQiBBZGJABeYWX3INKUeIdik8hT9sUepOIZFqi03KtJ8WOup
yBw/H5NLaXSULjdOGXwfB1XFAzg8qzWVpYSBt8VKd7uuTRdPXWewyxxwau2Eyir5
C749DNZleFc7zYfdrVNRjJyolyuYSaCNlMGPZE64oni1gELj+CCvNuex/OB6XYl7
+Zi+IJp1BTh4MCcLtcJyAe3sZqRNVWn07F3AYEqIOiN0+oH6Gg6rjK2uOCStONWi
cySlqNsK0dR5ZSCAMkSl5e2SqimBcq7wwjqGZjdGE6mOxsRCvmr46xuP0PsVK2rK
kYhajpdbpEUZmAjYgKnXeCnmTvtnTZ/AtgJ94ChMU/ocuJT6N8myOvO1B4SA0o6S
FFVELnq4I3W6zuMo0Xz8xM83mCcLG28y0dYGxNKH36aMTMUHmq/Tyt5NhGT7xkaH
4UkVvPc8upYbwPM4YYk8c/ISGPskjLNcZ4kO6ibSpYqXS+7QfnR2/WPd1zeTYOuP
yLKYoBQJUJRJuXp40DLP4kYE8Beu5ITNoihlzRW6G/TRV5/qysgWQHu8C1DZUK/W
aFrss09/AJxXSWU5Z7cHZ7L/uTzbcIJehyBf15CC7ukoqEXnL2K6PaSBmaAUBFfy
BBZMtKa4KcBBNIAUWDtCGO0O6OT9a97Bdzz3rFPWm02h5nyr3hbsxhirAmrx73sl
8qpxyjTMbW9s9aMCbDJk99Tp6GTSd0BTLHC6VOkXCgQ26EOhoKxx9ejO50J3TG8T
nQoWfXLkbHgBBolAUbkC9AF3CsCV/R++nIY6qS4aZ9qdkTESDRSu6+vbiC3ctY/Y
0ulaF5iMRCD6+VsjR5Y0gvmaqZfMwYt1Q9seXfM1R+8=
`protect END_PROTECTED
