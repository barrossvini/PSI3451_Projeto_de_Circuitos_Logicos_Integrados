`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmwBgi7nE80lqCJXkoL+2ITTMOBfPS68F5v59nJv1PbKsLl90lfMF9vuQgjbo3cQ
6PGi92TJKBFi/reYIe0iWEvTdIUqlHs1q+SZb7ih3q+9rYMJ9rKu5eSgU8q+Af+l
acbqTnW08OtPZ8kBjgIZZhzFTtRrq/siS5bi5RawDhDqHYod1l0vdpmXCkeNg2u2
/q8hv9iVEeasnZDlOxReewKquFxPZlk/5/m3y89pX+ow8WGh4e4BaxD7wn/kdi2w
4m5Z+gumg4V24cjlmji6/zLeitj+LBCGgtL72fVG5N6F2sTsed6CduEc5gC/CRFF
pqzy+jC40nwQ/odiHILWvm8s86FGwCad1ptw0kZXMYOV6LYLWmq9lEZhMnDMaXc0
o/ahRbMlEV8mCPngzNPH7iEyXxFNMsjTir9PGOV6vZhawS6ZVQlKV7K2biI6jqSi
X8iPl3//HMualggbH/N4duXylIyKq3ETGTKWktqviRgoqS2ZN42+G96BXg0G4WOF
F5YDuDJYHucXHOs27/+wevk99fqQy/V6WR3MbNioL3kjY8NeJpcXnqXkcb4PHRa/
OFna/uvpZvGaVJpOYxhFEUTcXWfpP922I3QJYFmAXhlLz4Dpi4LRKLPyjLBuXSNL
/0fK2QWLmOwjd7yGQ1/1JjBAL1Tj8VLhL9LnjmEs5E26jYUiusCxqLPv7i1mXY40
zB3umVDzUZbRkNcrW4l5V+3I/HmuSSJ1fejTBhEZbyJZ8bur8w8gtIr73ckpT8TF
ctWxg+ertyogYmOLxkOfJ94Y1F6+keMofZ5aDc4uDK9uyKVxh0aqius+rjqLCWjF
bpCIK6EaeeZpuRf3JAtzv9+zlGFJTF+QeiZPhhnJnuVcsJayWwDqOws2fh5OVUaL
`protect END_PROTECTED
