`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kI8koarrzYRYQku3EiYQvnf0moXlO4eUvDr1nvCQd65Mgl/t4OZbEm+aRwvECibR
LcnHJyi6SDr9vaZFWMyLg3WO80s4sPPhpvIMpIPRh/XehjawscVqqiZZbLMGIsP1
C2XJWyAs50/QKg/96AQUP/ag/2oQjaINNyedMqPxtkXh0ppi8MvtaWCVvWs7G1hZ
f2RVXanibCG2sXiD9l9IBcc+m9u6XK4eEc46x4bcqk5IBuKmTFY6XwwVM2X/HDOb
atIRyxOXqxyI2oMVA8G+gOEQ9EJujk/fDdLyrchLH0oW1e01y7npEvWA53u4I2nz
tmrxPJiSNYB/ppNXu9WlC1P8vNOwrR8Iu+yCb/XJO96nxHyeWsvNr4doLPOFBgIY
2V4qBfs2lZ4JlR4NDG8v9/pcXYqXzCglF14eKsWNdVs45PYde1+Axr6xEc4dcznY
TW6PdRA5lve4YcJZPX5mrlWY+ZzStKvILDIKSMIBvJ2CKuK0erXnb0UajFw93nuR
irkgyYDWGHhsadseJ3tPh82UX47Dh2rHw2Nrxh+MLcrlQiJx2276UcUr5FF4nFX3
rrUxbQnPE2+qRxdiDLaLMWANk9uhEnR82uSPTS5L3kkid91xvNfVi7OkLIi29dvw
kKHM0te3c/cSq8ANDdLh6yZMUnf8eaAvk+0cLyYUfC1nhwnQPpPMzhn5FspXO6GM
Gt1KrV+imN7a0gwqfTTDcrUK7V0wGSOk9zNChehnkPjncVe88ZHo79GQB5w6vH3p
t42vxRYhchNTLWkorNNSh2TUOKsbT4729+OvYHuaW7xNgU9g16IbWBTGCfB9dlUI
qs+XunczbKvZst8k7C33fAnX9+btbbH3aekeWeg1iBjy3WctU4ZE5GqqZPy3qBbq
kTjF61FRsj5ZNAraa+6O2dzRmg8p7X06T9fXfD85OvhkC7ZcUxu30nRVgrlFFgRh
l50MAGEf/xFDBxjxBsk9VXgD3vpf/WPqisxggkKfat5nYKjnPlFtQCgpAMzFIbP+
z9rI3EgMXT7YYytn+iN1mdjq1cPVX7c41nq6xgKqpQhOLcki875xgISuyTtcI6sC
SkaAbiCEoVNON780t01Z2ytJ/ehXj1SncjzECTQBb3vpJkWgPcVXwE3K7/rquGQn
QNBYIlLtNcAb9REVvENR6V53LSTTMH6pf6fHu0/aALY4wtroPVJh1L+SpFiB7Sqd
egSN1sl7kwRUtStpTZQTUUaD2WetHmkE9g56OP0ebk5WlGvdQ5Wt4crK23Qtp/rU
Quq5THamYGPkLY8/kZMeoZ/sosAVNAbwDWHbOtDbz+tMpyPad/3UdIXsHPlTK3Qz
QuShjOPX/5lD7+YEhdKAeQy2gGmVASLmXFl1uS3UJp+eyXyD07DGLNOLUrSM/Z+E
ZpJdF3uh9eKmOb1qlXf/bE1718fd3NgRupifEnkjlioIm+1BzuLgcXNtX+0wjTTh
ylYspnVLPYusuceowpcI+7iswMHwG5OEvsGTXrTtsv7jWaQdTrwi4YawFkCZnQJn
RKSsw7ULbgCMGklcrEu0X0xGjblm5hqW2II4wpveNk4nxb5nRqlanMqDXtpeInpt
nHoeaV7WN9XlIpGZhd3QcQvnTFaOvCTTHXy/EX1YfTIh8QE7pMGltdjrOUIkrfnN
U0ZXEH0U/VixAgD47Xt2xcsmiFqdeLMP2CnTQu1QUTECm1+wxcl86oVqfNanQT2R
idjl0Nh9z5higQNTqM2uqamTSfALcYzsJPiHrnpd7gZ4bn/Avjra9SnBw2G2ngqb
bvCOGhb5Q8FlFsduJioi1JLp27Gvusgu2dgzxC6ZU943Oc135HOq3yDxSCRuBX2e
OrzLy37rbiqq8SOSJ469B6lIiaaGRXtWtATqtbKhRU0CVAuMUKqK+3ubwTzEaL6o
sGZmlkLBpn6QUNcKa1nBLg==
`protect END_PROTECTED
