`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1mzIeFy5lUBPr83bFBZ9EBGs4OkdMW3q9u9+56BO8vPsBAhXG3+dynSAiZTPaC70
mlAtBUqojyWzUDmRADkKw2g+lVzIsfJXYCSYweHYISjQ98BZovyek3nQh5hGTW+o
rStVQ35UTaHQgcg7v88DhbD1v0u/n6GVkoS0MF5zM1tKuivEH+H+6Wc7R1uQZYe5
y1KmMi44MBKyCXLd4GXI/bNDVVu1dVj1evyzPCEyfKaaVQW9w+9Bjn8fbRZJLu5R
JggEmjCZ/lvIOIMKbsRZMEzImhadc4Tl6DrawPsHQ+4drzPt/RTMWaW1o7OgejIO
aWtBrgHq2+2rTD1V/ZKf0R1CsHo3gcf2kk7SXdgcCnFY+UL48M6njXZOlvVBEnIU
ZkO4aN5vBkfDtgqPLIyU0laCh1zqlPgv7bJOVEEq33rcKJPItWhgagT0bvIuWFp8
fM6xLO86CFrvxtMnSk0oGbk5k9eHN9TDV4iJxxxFHa8X6DUtKeQO698p30vv7tAy
ZZAwNnE0SiIycdFToCi4Pc9AAe0ksGCenAruKna4bVkfnvc2hk+sGl3LFt0ZkqQB
FR47Y0r9Xuf3xtqQZYiEiDKbJg1I1EumgLAdGcPE3lmZvveelPheaArgrmHg/2e0
ReWk8B25TjZi/dn7A0rF6XVSA/2WfVd3HjDvIoBbjLjskWtNCtoq6OdlZXrSxbma
7TYlHIjsiPWXYTEHjDL48MMJvV2rcyRtMk5tniPNiQbPNuxDp1ZqFNR5/TMfgngW
lRJSX9hvRex2b3PYTsyihMPpAEpyJN7t9QfCvFqzT93SvmfqvXy9tTZ6rVWauBUV
GNHJ23pM8pEOgc5zDT77bF1FNKRBPEPGVU9HbeB94uv7P+dy10LQ1Ew894pDkQRa
d4B8xuvQ+mVeudDXMHfU+RSXMlJZ0wyUdjtCG082BCzQokyJo01xDkMTfhDHuZb9
vKCIhKAmHjVHDbJ8M+0vSDqn5xaanmRu3TZtok5Yznxk2pBfsr+xwNe09aKMzINm
1EjzfyKguSRgX8a0WPFeRqHDw2H58qe2GS8YGX3oq6w9FnvKJE4uplYo0l36esS6
VRPHTBHyBSW8ZqAnKulGQfLgYtEAs1+c/KSBwpS8TjLZSMkvPCsrfdwUaslCw3xz
nOj8wOip65qRqPCJjygmv78bp46ytztFyP1ITLzo3nrFSVU7d/qqZUilb5OFz22O
QyNnAiCsVQxMOoayf27fFSTbqQpVapWKhSrBVP0Y9Dshvc59GYOsXRAcACldXfsp
Vx34N8P3navQEa7+0ePU8d9bYzxUsizHb3yd3Pzx919JtZlyoY0+2k8nIdWvPbaQ
qhjLPuDK1DvqKg30BBfnebilCtBVakZkrQQ4PlzYdwI2B1TDSP6rVqfunrtcmmW9
iEKDec6Unqz8jeFj6MuAPAQbtM/kRGKMkPCsJOX9lLx81nj37SSosPgPNnEhtMRA
GWYEV6LjMK0LGKWGkJpY2Ba6zJWokJB5HNEkXGDGtGRWkMYlRyb/d96Kh4YoVDoe
42MajO2P4N8obqNoZn03c9zT3WjZjAq0+I1toSl/b/Bo3e+DJRG1pA4TjyTKmhN5
sdPRhXnBgv2ZYevJ9jaaOnNzwupjX5h1RY7BQOfWcPTzyCuHho5+HC5bWis8spnr
Lw/RNooWjmb6VDQa2atKhO9DoCicnotX+LEJhnDhfrBTQ4pkyzMgEqUPLrA0Xqb1
8KDQC+8p9LB+mI7apm3KRkZuh0VC4/vxZq/5qBu5ATUulxkVR/PpNT9V9Ik03TpW
hxSVbNTlFRR32gh2rc2ObNMBSASvCRGD5haHHGz10Jg=
`protect END_PROTECTED
