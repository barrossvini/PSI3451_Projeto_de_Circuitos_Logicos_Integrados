`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gx36CVJpK4L5vIVxFmepTqzNzMLs1/jFtmczwsIBrQtTYL1ODtFOzfog2qtqo4yT
dlxXAtoHpIb0OEqBW8PddY1Z5Q/QjVfQojLEvAzZT0qjHHY/W7nf6c6lMnDz49d+
/0yUl8zAzOqJMhgFvgkwE8fxOYUmlQmVvPvG7GdttxCH0kS5Db0HI+6EhLHT95bZ
atR/p+dJH3YM4gDfQylUSF0GhxwQIFaCyaE2TriVJH/1e5hidiRwgkM/ymh9iTkT
YWkt4cMqMLocIBI0QD9s8zAOzUUyGrTGU0mB1Xlt1yL8z/x+T/Dqev9dgljBxBnz
XqBDkdljEhtvsoEA0jXqJ5oQy0SefrXjHMSw7O5fgP/8m0EB6udCg2fCNgS03Mnk
LqJm7mmbVtfFXR/72hlA987UIEsIiX6hzYblYmdK1gvdrTrJW9avci2L12Wg3dnQ
Qjcx0m3T/rzGjzgFYh3kYxmQeLOl3RyYIQ/kw/PpV7OyDTCn+37JtgGp7R4UNzTD
R41t89gRDZLgjk7sqKJ2V1hI5stbfqh6EjrtX2sNXQLloN+5sgB7CnI3EvkSH+Jk
x7OirDDtJh6YHGHQpjBZAQUnGlgQTqQayMmJhv4n9nEcqSBZMJc2WnEJR0cMEggJ
WWzhxU/D6Mtx2ELs43MBeu1r4npRIIVgcblBKJQXAQewNV3KBAXxPhfTkUGfqaV0
IJ5WzJo6RvS0uNju6l1QU9k0e61csHy56gLMH+ut75/yQdkeSmTI2O55NH3giHBd
bZte9/Zfkuvf4bGhtUwbZnVnxLqC97PqfFMVBpFofGVzYymPC35fnO9PsWcRb9OQ
4dPEZtQhvF/2tr1HtBzdTI/0Po/zWfl8Z90O7pM5nN7zP+Wp9D16alA/j0obcxDP
Y/+idlfP0ssVq/gD+pIW0/QoDDUCaHVxBNecRI2uBj+ODmjrwbxqnBTmbNsYB1j9
FTV0PnYhKvz/FhmAXoqmUlPI2xUrGBWwv3Tt36UQ2Nj8B3sL+GVKU7C6wGPHZ8aM
bEssPL/ZTbuKxQoXKVy1+TJ1/qvjuCDYLJHLLVuu6c6Ri5Ju5KOop/9Nfa7kePhN
i6NO0rBJDu4cktiy7RNL5kUahBLImg56sgKxqOHBR8Js9H2D50X+BDPg3Mcjo/ss
uDPKFNOJVBlyG0IklRfiAA==
`protect END_PROTECTED
