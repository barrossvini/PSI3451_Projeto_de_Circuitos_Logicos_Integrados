`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7S2qyAWdu4uQvGSnADz2Qo9yDHz4ACY0hXjaLDk8sBGm5r1N5Fjcp+k56dIwbQNE
9n7u4U+Xe/HFYxN8WH92e8EI3CRDxS1IECNFXynqyNABKDse9FGcETvVHFAkT7FM
15D4vk77P7QOwZTkocPlhp3go5pHdE4YsKzmnnw95W2/Wj6XoJJ/zatXdID9+oQv
DdMBMTK8xcj7cldIt1B5lZUZ0KRg9Eyihlhtl6vYsdT/r20LJ5VDAEJR6Vn8PBd0
NERFLW3vSgKUJ8CE+jNEqEVpr8JbAJKQCQezT0kdkeUIhe5Y+Qqzg+e5xdubL0X9
RY+Adp8OPR0L5QlSafefCyIJi6OlBGxLzCtjSE5NSeb0tV0ksJUfBgAK45g+X7w6
bMQ+QfNuTxuZdZwUE+uB3lhxSeRUPQseKlEF08ha9FefdgNbwX3D6O+QEP/tqIgy
ayu8XHXXpHlBttZy6unndJG/NfDALfgbMcACshBP1XCC0LMWqyXhC85SyT/UoOBW
HLuI3VeZWthUlfw9O7Tl3LjQnD1r6i2vFBawq/nkmVrVOeugZ83ww2hKlbNvVqdy
3eS4DqnOEyxgycLztC0it1Fs9Fo2r/E19RD43ZYuuZOCVj2iVGiVJYwxd4rDG1x3
+qJIEWWHUO8RP7HQ+wWKUZp7gn0A8/e9YBepA59+6XXXFUVvhlUtlj/jZE4x9uPS
Fk2Blxp/x8fDpty5xlVKPCFRS1LummtS3HFdddgwxIeP1IFYI4hVAOW7nCzZ4q8p
LJYCCZl5bUFLzQmX8M8SAuKzBUbX4j/YhzeNjWWuXI/CNRcrFb07q7PL28t0umsF
jtvgmSOvrzGAbusSOXQFeq9Fb+ui9+9+9jkWNXXSZaNy78l4eaUZ0mM52g9lDESR
Lpn9CtsUYw54i4AKb0UPLNvf6CBf04ha11UvQuBiANbB0UPaGKWgZyNPCnpBLuEK
coUYyF/aYrdD4dLAfMd0tr8i/9ONHBH+xSbKHCQ43CtfHcYCexrHzfDalHGQn55I
ArYzffbJlqWlF4qEZdw+uWZquPu0wYIPFxm2+PIj0iXmZlJ/fwuYnqOC0ULzDTJu
aZLrgb77lWKhmcDdhNZB7HkbcARDEpxWPnHguWEXZU09+nhK5G8cNcYiuwf9ozuu
Bsu8fal2P0tcXPFFVI+qzE8OTpJnlSRY94ETvOcbzOyTp20JSkaHiIO48ATu0aYt
No3Lz7k9OtTxVtWUij0QH8mENQTkmizzwqF+k+JDWTs=
`protect END_PROTECTED
