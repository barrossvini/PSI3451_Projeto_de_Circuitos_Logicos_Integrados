`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QGwFMW/Xjbh9WFkeyksI68KZZ2a8x/+ZpjkdlpiiA2qlrJWIG/6mq4AvXFgm3/UG
5udHRwuqerk888e4NWZBQYt+h+Y4kC5pbRMXVQGTPn9Ckzy2V42aEfmu8vuBsj4O
KFQ33NBxtYiotm2k50bAUUYMZ+e4zGruGjPL7ji18oa4gfYrVnGMPxw+zRef50A0
kPIlgzvsFZz309DUwdp9Ucn503H7oBc+g9sGXz9jtU1wRhbFEWc0raS3Bt67/Gbe
cJumMpxj4uGjQ7RLQR6QxH5+QlRbHqvNN9y8jA/ljKpk8I1gcrT5+mbO8D+/tmWB
/zPYU5Tw4+2aNIuOph384QMxoOhS8a0J5kpFjJlP9gKa3A+KsHwjR5Uf8vF0Ysjm
VnD/mclJFcAI1/pGLouEQeCkzQhJOeeaob9JKKtuDsXT1bbIO44aA27RDwbxW2a1
cSe2FH15PBsQn3JmZeEFpYoJ4CcK+ynynLLGtVDI4Y/E8wsN9f0mOHqEZ6PAsP/A
7sbXMU3ebRPtjHD6XQOQwexymEYNFCi0ivdHmgUkeIxB7V5Zo/kBtyFUW6Dr2UWE
KyTITBAWndOX1VYMKEd+XtC/RDrYCWROzR35FVFxNpvmtJPJaNHASEphiFmVZY4J
ECoOqN+L5rR5vT7B10kU17PvdFjl1criERQfDkveHgXDlhQEclDtHMxfqSKnulpW
chnkE6iF44UFBMCgDoVd23UO/PSzzSom6at24ncdEk8n20dOTy6+UaSorIH+2K4W
DEQ4d/sqM9gHl9E14JkUIUeVXTcAFV+MtpYmhtsesWiIMsFe5NZ9XPkjRAkJ7VgS
c+c69JKL6QH0ll5xAej7JGMEG0z6Dp44yWEhJaZ3NpfV+IIa0F6Uiv58+p2yBF1p
c4ovaL0BTO/wA067ju0GqrwM0a2xou4CyPRiQQ8lYiBHpmQC9JCMrzJukvVSucOm
ybG40uUgWUQWoZ4NYdIkHqYLXa7v53LNEKODIDVEB50ZKZmVif7bOwbTri54QQbF
8UUuidQqLcf+sx8W5m1qSm6J7oMm8/EiFNwCEVGJDh0=
`protect END_PROTECTED
