`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vK0LUwjoCBxdmW6UPFevsgdb51YJ78aNjYZNVTmMjwBvVS5dxMyJLL2rnwAyeViG
ljJsqeljteqAMSWLFyveoayaS93OP4KW/inIIwG1Dt9JWLVqpSu/cBP2peuGCj4k
0+tMJupuJdbGYoqs+1e2KQpMLtdfwAWBcdRpBxwDYo8B7jZ/lwiH/rHC6K7OSFQf
sctuWsYuoHOTBAavjv2PR6C5JajGocafTLCYFkHDdUJTv8lz4/h4PPaqPjIIo+gJ
6RuynRY4bFd9Ek8VeiknmZ1UGJWBZ7v/0D81PIVI0tWaf2J5pDiN4nujTGAcfLO6
jgsgk52ZJEkZElbm06mP94s6BffSTZocoo2/zO3y0VVCFPjWFYnjok0/1C5YLw8x
KvxHZs1kh0n1cDfc5Km7NJEoAvcTHcVbw5U+SHh7darol1/F2wmpUhhs3XHL030S
NRFsw673AEnhOzTw3+Y107/0QHazHCeo0Be5GfRibjaAuc3yl4SyjiXBd9IyHj/p
jfV8VZ5jTMM7TpBcslLFz1jY/kUW8oFeNt9i4iRKG/vvW2/BsKi9tSgx6TK0GW3o
udtE0SiqcXls4KtRtyU9hbLYTRQCEPxboMq4HRmll8GfYbzeFoOQAbRtQtyKCnW9
TauSh6GtXTO3Ra6I7+16PKbFrSus5NpCvq0F+dae5MtNBz37kDkqGwbPyrAQrKSf
0mJ9bx5LFEUuoY2j2nrFepblFTox0k7153BB7pYbMoPtKhwLXnZtk9MlebPmev5u
p+R7Av4M9itYxRW03vLXjEpty7A4cAmtfRNOe89Tr7X/K+kBnXEfDorqDXqsF3ku
HsjPuKOmQsBZuoxkxy971NfddpYKj6W1T+at4QWqrwJNSCVUjNxY0w7ZzcFgp1MS
3yzKplSP0DgSW1RvC0xUD5UUyWVhDijvjWlVln/uBO6qjMraKt0cKLfcCtG95M7m
smHOT87dled51UBsON7JxgXETkkDoE88DGDsdgXSU12U54qXBbuPJ3EUjHh5PErs
LCgGm9nEN17wmZVfhepVzpHHfHBO0VRLjDWqTEUur8W4mhM2k3T56ZTou78MvDGP
cxaKyEHv9lY3xPXv/IofFdoOkGeF5jBzKABreIML+4QRu2omI9wG4HJ3GutPDERR
`protect END_PROTECTED
