`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O/iK/YNiekTO+Nat/i5/09A4A/ezS3TeYx4+08kVS/LCBZaux5mQGwK2nwuFEpsS
MmjBv9LhEwxNFmoq7r8ve/vURrFYDNcKPmR+jY/UMiKNkxEb2ynf+CgJ9QuQd4GG
gjnEB+qovE5n/AHk2wOVj1SrEFOBw6WLwyJRnMWccd8A3nfUxz4SilfGlLiEPTum
isZjnEyMPbI3O3zx1JGZKHG1qLFdCRLV2ePO/HoFQHRe6b9JAFALtGLdAvURah2G
b1kiZVGRurxHIV7YHECd08lHPnsPonTuAvfqNsZqiK/NBaUmTC5dRe/6HYOAFLwG
oFVGaATrjrK/A5rBTHhFK1S4ruqOO1c6GhBHYRD8NNnJk/BQN5FhGv4JpmPaFzNC
WjDl/pdz25zPuQPaNtnrYvFih8li81EtWtfiOMpJrsS+BlYPF/Tr8OIvgo+9vGK1
VAYAQwiexWIOuImNHOHb4xIbEnu8kbJksSuzSbtf5x9/XPUmk/u1KRJdv+ou5mxD
oyBskj2cHX/PYnWsf5WoT1QE4T9Lsj/GMcltRvXoTLgdZfBKFu+9Y/ioRMfARO+4
no/pB2/Cq0k+m5tC1HX8S/3uSYPMlO7DnrryQsqipQngdlLVjx8sGM8htkVfFYH4
fccJhwCEUkb8gXB681TqZEreE8VqtKDeOeYH7ftZOuBshwSzdMRA4m85Gvw7sAM9
UQjOioj/v5FCiR2cnuroOtm/Z+eNif+fcVDznF2msyZmZYKk4fBGXxDZVNL8cSdz
vUyHCT3Om+I9aO48Wpsj+ilsxFLkSnI/hjjYo8PzqTPGToYHjBU+WqPG2GpWyA51
tQawtxszHs7ILCJQopIuiw60Q1OUmpxqLCGr1fxKN+kT9ztRgkBXYqSS31QJpINT
yv2YtyP+EDYj9C8BfGPRuA==
`protect END_PROTECTED
