-- megafunction wizard: %RAM: 2-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: mem.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 350 03/24/2010 SP 2 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;


ENTITY mem_quartus IS
	PORT
	(
		address_a		: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		address_b		: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		clock			: IN STD_LOGIC  := '1';
		data_a			: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data_b			: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		wren_a			: IN STD_LOGIC  := '0';
		wren_b			: IN STD_LOGIC  := '0';
		q_a				: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		q_b				: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END mem_quartus;

architecture rtl of mem_quartus is
	
	-- Build a 2-D array type for the RAM
	subtype word_t is std_logic_vector(7 downto 0);
	type memory_t is array(63 downto 0) of word_t;
	signal q_a_s, q_b_s		: STD_LOGIC;
	
	-- Declare the RAM
	shared variable ram : memory_t;

begin

	-- Port A
	process(clock)
	begin
		if(rising_edge(clock)) then 
			if(wren_a = '1') then
				ram(to_integer(unsigned(address_a))) := data_a;
			end if;
--			q_a <= ram(to_integer(unsigned(address_a)));
		end if;
	end process;
	
	process(address_a)
	begin
			q_a <= ram(to_integer(unsigned(address_a)));
	end process;
	
	-- Port B
	process(clock)
	begin
		if(rising_edge(clock)) then
			if(wren_b = '1') then
				ram(to_integer(unsigned(address_b))) := data_b;
			end if;
--			q_b <= ram(to_integer(unsigned(address_b)));
		end if;
	end process;
	
	process(address_b)
	begin
			q_b <= ram(to_integer(unsigned(address_b)));
	end process;
	
end rtl;
