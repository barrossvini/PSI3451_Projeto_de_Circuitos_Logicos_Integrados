`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WdNHyQAqx0L8khlNppmfRqZ37WK6ecxHBgydhKH2AGim8X3JC8wJuAJ84wDyCUZR
+IxKfTAgfForxGXgH4wXKwIcK3GDCbyq1594xDD0T7SBW/r7IUC8xRbOT7giSLy9
KV0k+yrLfBTjR5ecSMKLJ84NQde4W0jmnycMcFxNrgXp5egXJFbuY7fK6nuF3K2K
vyUUtrGjt/U+fsALROopZlLx6NKUHvMn2YvZXlreItIybIIHyHcrmCK8kNXSBnYV
JtViz/IWjQ+kTjm66+cYNplUE3I/J6mcMnokx2jAkhANxVYbq1Fv2IA5DAo2octE
S2I4NLJXIqPCBkzCFDPLnG38pja+7A4JQTjwjU4kNntMYlsaVmNU13mYzP5mRL6C
TsXhFUy44slaOB2UxCRBG/f7jQarl+WWqbmjxE0NVa6XqQa2dxmobHQDBDXnB8vz
y/egADUqqQophp/KjBIPfg==
`protect END_PROTECTED
