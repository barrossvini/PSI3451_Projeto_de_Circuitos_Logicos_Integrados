`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W7YsqQnWKvPjCgZylxicTq+HQpcfs/EF5W9Rm4z4/NE7T+bMviqqXJjvnd+0TayJ
EfnddSBi7imIy0A+Aydh/T24LoaDk7Ymh+aQcbDPTzxYA8SbMsduINTUGXTh4kkW
6aQGLy2xcfkQnd9HriPcRu9lTLqAhMiEsxP6ykiYE/qrQ2NpuoVch0fRUXH42lhK
+z6XKb1ZxBmwHll+bx0ccxcES6JNdpcTAJOadjHuXnHzbIOzYMGKQJcD/hN1EgUU
ojUwLQNPFKjkhI8GW7vQ71N3X2C7H0syXpjQiCCtu7WM+2ss39q/rHDV6D4qksas
V9SNC/o3HPke43tml2v7wrQESWJW1yA12JS1EwDxBL8Yg13VFmFvJuRU7YeWeuLK
RlYCxTn9lmX7dc5ZrOQByLfvDA/EPUpmKlPknbSfwaAq5Jbuwh9LwGtDXjvdUjUG
GTVdu+QIhTKeXRPNcpvTY6RSt0LyRgdj2Em00f3xwXpbmrGM4v3nkSMA9oAbM0uT
M5FUsGNRcq1eFdIRUZoNDpQg65hpzxl/tpf94GgFPcuScr7dtKSMuNtFr7ZwxI2Q
yi9U8lT9zQcrOSxmVy86nzeSQNLpbH24U10SWN1rfBim2s4/ZCNMPxdQdSE3bkaG
`protect END_PROTECTED
