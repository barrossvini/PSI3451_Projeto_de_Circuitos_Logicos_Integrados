`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PIe83pmhrVkJqZiKmC1xcnMrCnfncTF34+yQ9WYAWVaV/5ampG93bpJBqw3/EQ9q
1PolxF8DZMavzLVcBCjSmADtvPxSKQdJf2p2eTL4vBF8QBEefE4BdCuq8Ylj6kTj
y7oo1FmV+DQB+cVF1uLnpnVBc7oy6Vfc6M5YREXSps/lRfQnoQqv/KVj90hGyhGj
`protect END_PROTECTED
