`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gc8eamzMCZVaUmw+dRvvcKlKfjOifJZBAkBMqNoGmC3BxeuLUJC+uipPBiOvNp0n
MNoLR0qyTyhcnCR9HKKuCEnFZIi58lra1NRzzVc1plsgwQLnMFetNUPyzezdGnA4
ssbcoawqpC8OpqVcS1yv6OkQT6Qy5lMZP5BNWCoC4gSeBCf5h5BzMRHjr3Es8S7V
5rE3Xpv6qbQrfxeNqXiLidnZ07jJq19dGDPlg627MO24DYtdvgedqk+HYVFIx4Gh
dvnRjbQ5fBB27n3xxcV7/prCGdqnx+xjTwi3IIXsPmQzRi1juHuv3+sVVChIKwGv
IOS29i0M2hbVAcSwgo3cTBYcRDIezJVESWE73QrGS/uAJkb0Avx5zZMUBXPpJWBN
7N/pOnITjzVUiWov/10OIfsLSuR1pkTV2zDXXTGwPyvDO9RJ6UxfvbQCkWhX8wkN
A8Cs6shMoIe9h5wG5Yw5yNUcumd/G6RP3VYixK6BSzVesk6w6dzE4Chij2Y/vLEr
/4xzQFdgX/qz7gf3loD23cilo0P9gjYo0n8ozo9e9/4si5XKcZcZmxQaRtf4C8iJ
4ao0Y9QisNwEDJPvTG+4297V/60E+2E+bfKxJ/86uDNdixCl2NMf710A73XSQZu0
b5PkLh10QWpaWfkaX2Sp1PJ5kez4jEMhe1IpaMCaSEQQX0m1xYCdWilP5h8WFvMB
to24GVhyZSgEkVXRkhbvd620GDGDbQrACbdYgArGNNRpSOjbQ80xF6fLjbBI1UCP
SNjW0I6fzr+M1y1WzFWgjUds519tmZ0dbo+Y+2Ff7W9eof+J86OyeJRBTr5sL2pN
SPW/miBITJEWRAGYRb3J+MSj47PVeL/U5g4FWVmfctX6NqwifeF8Rklh1QgLXQpo
emFgto+xiVYqcvwYMimTNNnIbprHWnDfxQw4FMuXyM9R5rTe0FoF5ZRHcj5WkCIL
F5gbTVssB1TtPkZI0KLLrKP5Onu9UtqxstOzJyyFsLS2UJebPbc4tuTl0XTTUTpS
PJvWyg2TBiNoHPsMq/UEaKJ05fX3C1pFATzFBrnSFNuVyUcWKo6gY2h6qB9Hdm1i
11uxng0Bzuv6vCKbzUHiE1qzZ5Mpl7WNhEb3vISW1zQHFYsBfYwUG54i0hfNk2L2
l3vEcaXEeR5I+jppZ538yrp1bor+yEKgW/LQWPMjFtceN3qQZFiaFEGij+6QROny
c4UrNpqJGlNE3Vkz++rdALNcELLJYgp+SzfAvlSzDOLS+B914HpI0l14v/OTSoNG
IjH5zAU3r3O3nDdd0WjgJwFuxOqeUg85RxjJmAtBLVawsH/ehVXBlbsXzhHOD6lL
ao7UmhU9a4wHvjJ6N3ylOz4mjPJed9dcbL/a475wI0235xj6lGiLDkyUkYmW3Rr5
8xkKqCbwIRIJ/dBzHS/uoMTYhfm5DokXo86HQG0YH8D1FdJUZyg36/sL6yzvovAA
dMQcEzAXzkGmHQ1f/2/tNq6Bjmh3JJeOtdxLSz431Io6H9+wiv3umbn4Qjiwuiqe
ynnPDDxkjNLtGecVP8JBrobj/1q7FiiaoCsozrfcZ0sGFrpc7STPTxSjTrpuKBPt
lHno5MBS5lv79meDEBrjran7i6GuQU99Wi6q3+gmNakfoUIYimZl43YIdsxRGeVw
AhjS60iZNueDt35vwj+nQ3vljtONaLfs0padRMqMF2YYTPzZuCLzOoTevkCkjbje
MrntEJ+uP8rxSL4/XZDE3Q==
`protect END_PROTECTED
