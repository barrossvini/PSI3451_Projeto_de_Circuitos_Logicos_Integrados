`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
103Eo+khoxuKO+bEjiVzZWnRD0uLK3Ky2tppUSUHHkCem6IlBbtyZAPU1MFXReQZ
pRLOfEEV/kiIvCLZlxdBsrK4zzmXWl5+Ok+gIRVOO98BzrDxGNWkmkBogEdYJ7ut
fBOFoHrKTAt7YvAxpiufncu2LL2VfCYRkDLHinVA7Kh4p8HcUI4xTRWJ7T/2qUNM
Fs2H2X5VbK2xmS5AbO9RBBc1Ia32SI5wcorr6CsDqCduNr3bausA86kYi1urvRGV
AER8pudSMAnJ8nSlrUaKPF2Stqk/Qnpmrw9lycKoydSIGSyLGAXs+STi/41AjTYS
EBfITWlR4avYYI8ft8D/4FajOqmglW+Z9Sgky1VT62W/BU07NXw2jEhgjZg8pArR
zSmsGqvpNi0O5b41HqdDMcb+N2EJBfimOQfHaIris5vd2sBUa3RCrqvHh7H2Dh0B
F6bYPtszbJmDr4UtTCxkfz0COP/GpDdnwSPDVtiAefzUUw10duWWB9IWNqJTaulF
MO9FxyNuKhwdaaQnlyf1YSflwmb9mNQFVoAxkbPhPa5cHoIKJ8jscKAJF0r/QwXb
/QyhL3jOgaLJql3mzO+eGCv0UsEWaFcJ7OYEjvptnduikR9U4gPdU1/DH0JKfuqP
o7rx9PseRinGubkAV9uYCwwk8rINvSMVkaRMWYKQm0ViM6eLgDIInHphea5bOS21
T/EMEBkKB6oJIEEmWoZN3HCQh1bo8A128DLPlTwjL6wxvZXpOxmloTbA9ZYjccXo
J7fBsVtInrS9V+z0yc92hKt9wOYLYs/MgGjLHQ3/DoXnLRRqLHpZhVYSlhNbORIU
bzd9vwhAnoLehVIoe9dcsoM3YqcgCx6F3salHj691BTJbmoGl4ns7DhxUNE4WFVJ
eyEokL5OpBDrTguQWYl0WUFXzSreuLz55kRINQh0fXYRfHtmPLIxWbRo8K+N41Zs
zaqVUSq8qX9z9RAGZ2AWpAZ8wzhQ2qlRM0dkKZNbkaRBFuUkx1b8Mr0hk58XqiyX
cIJc/zyByRyQ8wMzAb/DZHJR8QiXIJBgKcSANR9rnYyHWk0Urbtspx2LgF2Fhdke
aG9S86HpmiQZYOsbP+cHwHL+2+PGFpvhKCJETCD0EQ1rVxghUZYMfadJaf+5jjTC
LytzcYGiWcdLLZ+T/CAPOKT/kY5nNoy4LH5trIWvVzfDjBPAnZlhJq3j9pXyvXSM
qbHaWGCiR6obDvt6s7m4YAHFiPQhz7oteogMhVevdzaCX60P61qJOtPxKWU50jqV
sHCWmx+GnNZiG1ftcru1JwICg8JYI5hKJySnkfHzu63hOL0labxnh12WvMq3LxOH
7Brt+BXShDcdHth84cdK91WSN1Ut5QeARa24iTz87WOq+zRRzPREAtSEkjlK89yY
KBtoIHONRqc3FTBbvPKM1yLV4ZcOczGUM+F0kNIOZjru1Psff90CYXcYYpIZ1KNV
WJjtZR5EYO9jEZUPI8kS17a6F7DF6ZO2pAbcxhX2iLlaAQDueJxugFAMrjP3uoYF
jAuf4/CnLzW2/8QumM3Lc0L1n65lY17YcmxGf1mg6KbJ+FE+SzSm5tIWerpHt4zB
JQYkxFTBnAFr8lXFsgj3gaFJjjsW3IFyRm+tUuFzFu+sHz2XSRHoSDuQjGRjZmEB
9jAzIAy1xMHnTfaDD/n8xTFhU4guxf59f4uUd4xBFAIsSD+3Kvl5fHU5K3PQM6U1
nyLiSX2oHwkgzRIlnCkSeEEpfvO4cI6RG8GGnsGVHIeCl0ljZ40qMhUIzyu1yPNC
+MuGcRblG4vd8dc7a3n+MufzVP+PP33uY8O6J9qpdKhUcFElL5OR+CQpBYKyvJOw
iMjWfTeLMWk+lJ6vyXVV0ls8JcQJbemhfjmdI3Hhk4Jf/EuCsN30B0dBt/qwZzKp
ZrgkSpbD5n237zVblsBYxuulkDvicw+dx5V47kkSExS4IKsP9B/qsiH2w1kS3iw2
Fp/rd2ldBsthMjf1ITgt+d3Pt8irP10aOOkuITd3hufoRIQ1D8u/F8cBr5THtSbw
bmSH5O5Scyqd9A7gyT4zZ51BVUVI0PiKE7dBCw3JdQcWXz8kfO8gWX+Q6wjy8Kzr
fwoont3ZWRAuBSfAF7VR6FMubVV+hRXb2px9AAwrZ0ni4ErcMuL1rguAmDqV61SK
x8MlporAoZawO2uhUiGcAdDlWFkssPBFIrTNAvrMPQflnhoeDJBU2gv6cYwGYoS7
8zgOUwBiuoUXPEy239kAOS0WSQbSbKqvDQiih5+vxVZVjiOcREMKjz5EDx8xj40g
zAteMuzGR5KJfJ3o1/zl8AyKDda5sxvPrrrWhZPt+kM0vKyfUNOCdmSOj14OLrdQ
1MUicxrDHgoklZ1TMd6/ltyoXp7WMa/kchWQNH2WzmDsLxOQR2u1C1yPSOlqam4P
lriNgF+deDI1XI8cM8KDQPE8maew1GJYyUOp6qRLZo8HWNUv8ef9UuaYuBN6RnpR
j7ITSTgxMh8AhWRilxXG+iH8wxm1Nv0+IMXHbVtkXJfF3Z6WJIsiRDBafOHmDamK
UoPoB3mUM/ahmUKOznEq6x1j1X9UZPwROuTC3Hkj5EvI1Q8BYp8joW1HbxOAm9BV
CAaQwECoSYYatoWVsy38UQ==
`protect END_PROTECTED
