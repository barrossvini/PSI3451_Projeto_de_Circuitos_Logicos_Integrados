`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7fEF/qGnN1mtgGryO6p2S2By0iyTK0T03YmM4y23R/XkE0CKcnPu+k4IPsIn3y3s
Bhy0K/KQkjNH42qDPMY79rhVS3lnnvhKP34Gue95kwsG3W7Z5wm5Hg66kLIX1teV
ODDcTxHozeRKhjOcKcpgPEHbKIPc4R71WVt25PMeJkWnZVT5t8gLdK+yBQGrQunP
wUNoopiLC4K+OszoHGjLCl5XzJZwbBlV2tT4FLhNXy3bJOZ9C/SGwIYksi5pqU0v
ZApewwFKUSkYHXzcVK003FGw3+J68cTuB3oPShmv9XN7mp05b9YdJTYpZSXrz2aq
jvm2/4Y0T7hrYjUfJoMNvqFpUh5kpt8LI+MBcPd/KIJBTHA92m1FwlbCMg2zmKQq
h2I6kTZDSAb4RXEI7/dedFSZ7JsRDm0BfgYaSlXG426G7Hzf9ltEkmsuHl6K/H+h
Um4NYXB9ZwLgeAIlEifBAINje8EHA5JMnWMCf+j/UoOqM0KLLJw6LVfNd23XjMh1
qTupbH5JWdkbJikT0Y+WJQFVX1JZaj7fC6jBDnkFZ+HV0BF+MDyd8AcYOQnY5CKc
KYIYV43qDo6RG8s8pSFPg1h2ig0GQ0DweQOLqUANG8OupzkhMGNpk8mhnpm78Aj4
jOjsVF0BpuFrChG5MlHDE9sVW6djckkmU3KXnToJRICQ4h1X5/7mGyAtimInWOnB
uywX3j9LLxR+8GjiCKsGYCvaMTnyTCWi2ZZgHjvW4Nm+wW2teqprNo1qTQLokaiZ
XSoG+FkudwQx7WyQkHDDyrAadGIvXT0KSjXFxG/xqId8PXkx0M9QNCf3pzGLOX12
WTn2fqj4j6mnN4kV4+66Htv7dkRhbr1oMB8WsCerjmv5bfcRKnD0XpcWlCqqPNfF
kAoucLSeM84MIkydO7Lro3+I8rJVf5Cbyg2wod6MQ7uCCo9b69o9FsD7K7p03smU
2/RIARBpE7gId9UkqSiPb+njstkaAPd2WeXnktpXuFB2ZNjxXrVfLSm+/zLHwc4/
UdpQ8ApmUXF+Zu+E3pdLBcmn7LWcGrFVlwJlNgmscrXf2yhzhF2stUAaNpEaoExT
8opifAoF/5vWYEry3DzAFdQgl94HRRoaMR0LQMdCgFWjV20vQMyJi8PZiWHjn6AW
m1F8Dxul2sczrIuolD+1qP+fthjfLUQO1SX6s4/NvpU3vWn2CK1ay5hlL0KPzRwL
4OEthh8Y/W+B2g5d7IxTE3w3ZaXTKjZxVQRiI3S/il5VzJeTwfwv3SGEdq7illVM
kJrk1+84k3GAVaZ0M7IbblJKclF73ujtB4faG8L18Qy1qwB3HbVvJovc30d3lATu
xO7Pb7Z3Vy87IYSDUg6VGDP5v+8aBgAYHp9ZBzCvhnjU+IybDSF8AbqcouqfHcal
XyDy2lCNTZyYcmNWmD9CFcZJGtxWf6rjG24JNDZbmTdevAJDi0251YS+EDu2aQdi
PuMXYC+sxRMT3LLlbExDJILxvhxtxJwtXV6Fv9+CqJkWHyHcX5B6cUdbfSR4wnBK
KyvHce18jGyT/9j4JUBl3AYEOQzA6I68Sk95lH9bU3CbTfIeQgkxeGaRKA+/qogL
Z5GAhOy/uUzfmWh+Ae65D0X2+dVdQ+i3blyBi6MFbKSExcnNr3y1mGaHT2tVz5n8
mYWYGD3nmarBfiNhoQCOwatolIdNJtuP/JIBZxtySsyyscN/uho1jwhrbKVd2H/7
RVLvT0Eqly9mLnzZ0ayaAym9umpQ6y1jC40AQdWcIx53CrGh9IH/FjkclUjPPjxc
nTinwI8OTHR+grnKevYI+bAyA9o0We66j2PbOPbU4q+KBBLFdjckdQXgQbFavig5
OfKT2zi2oQcgkzW1bZu3icYXSebyTk3ucMB1hYmHrkUOi5DfUqsKAi1pNAnjM6J6
`protect END_PROTECTED
