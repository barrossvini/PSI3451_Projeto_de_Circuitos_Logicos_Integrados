`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SomPwT08rNtrZN3LbIeKfAI2yHTvTtXa/6fR4vCxQq/Ur2Creu2S/GYG4Mwmx5MQ
r3WBC40Yp3BqMVVigaONMwr7jFG1DGa0sW/tx48/HJ87piJEWb9nNLs7Bhw6GjWh
3sSriG+2uFFuQq+KhmBBjwXtrOmZfKSh6BQFg0AI2id6y+sAxE51yu227CIJmeHw
FLvYFNdm4Eeiw9o8RixIjyhkNkWyTEl5q69ujj+RmKdc28xqptU7d52uCce2jErN
DWNz+JlHLgvFixmWeWo8qmKzRV2s5hvanlTwfGv5pQbGzA9JX20ZerU1VCC/WW05
FtSmDbhTQaRzuoQiGK6TeDtscYaypS38f4b6N4quyJVggTWBnxvURdslt63ba8GA
8/Dkz2aMcGOcT6EW7y9nWW2CWYeuyev+i84pCpyv08L25Qmg9e+FE6LQdXwTAvQL
coc7u7xILFiRZK+cEa2O/ipquVyhAOZMWwEp3SdBGmSovktOEvfVJQZBi53bIXa8
eHdtmrnpxDTB5zs63CYmFmuR/T2cEA/bukEswb4nJDt7B5dUa0LS8oPkoZnFbyJA
rHu/YP+AJJkFucPLBsNy9C74ws9PNaSSVsvp0Gizd/hYNT7phqAaMOU/a3ghcyj5
nIxmtTf8NRUE6kLlUV/TU1z93nhxXTHXNIienfcwAs+Sw6tT1/fay/gn2Il4cS2G
cX/rkm1keuTe2ZAJuTvd4eMduL471A+V6fK338chvpRoyr1PWBW16XwTXaExnfn3
6haapEoSWceP4fvgqB1LcJd0lXhby3DFWT5skyvWtQtzWH7B3kfKBnrWkWhrxmQs
u0NNNlgYZsZ2aP06/v69bxyFhCax42RzYjtRyI0junmPnLpJtw/UzLh2vY0YRDl3
6TyzWxa8qY+6OimGBFhzeryP2ID6ic+dGXd88yl5UESG/UAgLD2DVgRDp4fKJInL
gMVnCjp+LkbYX4HOt31hkqb8SCL0xGmR/AeIgA2MNSKJCLsdMQx/9w6DyLZeHQOr
FnhoWe3FxtIP6R8iYdwFBEygVrcYN+fvnAe8v16zLtEVcEr7P11CpmszAaZLZTUJ
40cRnuX6MZgOPuVGfhp229k18p9p8dpRwLp+IjA0S7S2a22VC9iQIHmK7adaRrLJ
crL1icLMh7ydfRNyf/C1+s3m/3vjOqt1f6NmXA89gLWi3A2iE/6X+M48QbZDjZ3N
cNBADLO3NaJd3JRzw8bj9f/7X6IvXdY7baYDH1JNS0mBcxnK2zG6ikEfVsPpkI9O
9bFTF235hgzq43tG+WMeI7KguJF60zx0eKUlXRZyjbGxD8G3Ly9DqIX8xOik+hRW
BhGwsf3SSjMDcFFQZ1Ay8/v+QKTckKHeba7OOyeUmZzR8cpxk2BXG+QcArclb5Pi
SnSKudaTE0Ohcm3Gk1H4jxtxYh/q/LiX8svSlBqgZeSLXl3TKV0DvGpWktnG4ioZ
`protect END_PROTECTED
