`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3WV3RxISenYYsEmO+tttAGfXJzN3LEB+Q+piSl6TETGin6D+GKY67SuZ7V7GWCUD
hg7Q4QheIakCic66Zl6MEdVXuaifcxKDb81o1vTKu7kwAeeTIGR3Pp1UelfZlfin
mavwh1Mf9FHuu7klTvocIYydOiszbAmWE8MdTq7QoGy3pvm79aPuSoq7mvFbdqtb
bSSiCFL3VzjduXkrYeXD+bqb0wKAUUgEkNc6Z+h7bv6wsnr2LOI+rAOmvL3Xy3WW
euOBLxSmnl2uEOovHPKW1GN5VyHYzTS0yiRD7LHNFbGFR8hmZqo+xCR7u/sttHf7
dGkeP+q0JvNSDYLRfYB8tnVRv4LpIN+hvWx8m+WyG8qwuUqa7oXRwK9Fksi6TqG1
Sqg3dydJqKLU5yZGv7EJ3Dh4v+A0S6TsHwNJs3+SPr9pIOuR9XL4jS11kXrhwSbg
NRM5xK1LRFELjGVUCdlHj3lPvid/6qir+q4dKbjtI37B/YW/ZyxKKc6uruljWo4a
QgaMX7hBrCrcx7E1yQ/RGRiKbLMBbQiHvO0+Osj8fZkAdc2+xdr7/bixAoXHIit3
p3cunmLsBwlLRuj1vlgTkTJNBI+Skj0kmanDnUKHCB0a4StncHnSwWzQjgWx5rGq
hV50M8I5dZebTLAoLprVAYgqTh1tAQL15AifcUB4naIypw+AXc3v+6NYET0739nA
5Cj+eQawzFfFTZonXl2+Qc25WHB6BjHVekjZmDmyLWRLzh+uAdLrCtRQzrGaO/3M
hP2RHcnowE7+ikiMm/HYirZ8V25elxpbjSz4SmdrLol7QRcK3TOb8AFiGGZVw38U
gWwpSuDia4X9bIYIXZPSTU+NCx9hYRAUz3fj5SyamgK0AnvwmbcEQ9Bvr7Ygt8R6
IoFvcHOtr03WkAbzXoywOVL21rGT+7rjBn67LTF3w6K1j1gcwzXKS3UvoohAC+Er
Jsreb68SCvpogFJV936ksXGQ7PU5T2zr9DfBBe0tSR3ZeoWnN94lAEwJNE/E432K
DqdtV/K/FYQpSmWnV8c4Vd8CVGmF09SJeGaTLIqFSkHk08VOK6EuD8ocC1kxBGsL
9j5pYhVqYJmJHkcwy7wDMbsCwyh+hLGICKzOOG2/mVjXd9NCkfRC2KKg0IrtHZ/u
AIFNmVmQbiZAY2aZiHHu77XO79WBpDzuAC4ojBR8nSOGmsfzAAZ4/t4eJUFw3Yi6
Ppkth1G4fCVLmMITfoJpyIw1ifezw8fd7PvOYbjdMth4UQ2Eocnn9PWwHgQQXkUN
97r4IvXPGoe4iFdW26hodbP4piCV8BMRm+mqa72fZ+CcqiozzudVpFUbjvUhmUYi
q9sJ6GvBBe99abEjoQt9L0nFbUiVzXiQm4FoTKipt4Hy4DmnP2mmfT9XHbE9gP7R
UIyXsuYzIAB3urvCN61DDBqUCemE2nDHYWDmEv0RVxdZSESK1WA5AWpwvcUHmMMT
RXF6Ng79s6CIlvlY78Kt+mdOTh/e5CwdnZVwn/fw/BmX+NSyF/NQYQ3AaLbEGu0j
Uv4gmUvaQ6CQRv2HfJdSF/q+9SajU50Q+kJa35z7GVRIgg+LUQorBVcp7tYhNeLl
n/goJN6LpAKF63nkPJuaXYHALi2AIJKgswSS/OezybKJRe+Ny86j2o9d155xgAUB
OBNG6/m0Yim940ZxvhJsaRsCazTEQYvo2DNy0Uee7k0vlPlyu+K3zq4bcQxqfrzk
t5dcpxOzvY05X2NRmffeV3n33sk3fiVLFEiwFWPr8BSzahL5lBcDWD/vieW7Cnun
lDRHiStSbjHU15PoJBbi1Q75w3s5LN3HpcXZiLO9ihAgE+Tuk//gNtWjQqbHNswJ
0A6tykRg4wTMcsQ+Uevqc69H3TUrrAyXh2mFCJkerqINDU/tcePBAWaWiF+8/Gt7
tYppLGLJ4VfvlCpuJuZZ3ZiC6RxnYyVXSk5BCUu/A7Fg8ToYiZu0Sa8pT9iAXc6z
ePVKeI1fOc90azfx64hiUFkYZY3H0IGIySN9c/4Kg2235aJB7Xl9NZnvqJGjSfIH
Jza1QMZVDJYlAOTgpJwQ5rsjdtqt1nFSEASWLoQHOtP434hgq5OYUOnGXyfMI44N
97wIkQHDzbO8oBW8OwekhjfHPeU1SiMmdnxKwcgk8o/XK1t2zxGdaahxZhQtOkAo
iO1CaUGrOLVHqmQE7ZHuCrtZO213OPesbylzU8Zp94wvoN1cVLTuLSMSGBF2y/y/
xkWVZLVeiBKxH/aTTdIh7HdTco3ExB7rg4UMN2Cnfz8UkVJuvZF2ZxhfHEOrJ1oq
+haffsGoZCC9lJNNlmmWgZn64C/j7hjgqWNoyi9l7R9atUZmIl2IFWxY41F15/Ff
eNo8jJqJp4reb+I/Y+pg9kEIYxo1amQ2z7zaQpxOPUJB5GM6fBuxlxsf/btigfsH
R+eDcqNk4WFK+Q34p8VUjNk4jsU9wzq8MupdvzfpukJT8XQ7w5r5MEABWApJ1K5E
6TsFUi2yeEz5JLXOcy1zCW8+wh/eXWUbAq/XXJdKxitYTv+kV62SMKl03KYv9Ly1
Fgh1vLQ5FTbL4X1XB6bpCX9mErUIISnVWZxbuCuKPdVdn5TaqhbPAJmmzH5lJXWX
syZl22wU2rCRaPUcgGxN60nx4BigNHMBG+qcqkTgIqWaFKFcflRImgtldHBucolz
ucEMi88Mqsw43hkdguTKC85W+Ut50lY5dhAMetmYhS7BhmR1VvI58W9Yk/nUc2JI
X74oVB6J/9UVND53HYzTurhvzR2o+HdNQdjEGeLIRjF34/NI+T9ddMtsOse9FgPV
XiCdjAyUrm4Pq/yHpNKxtkds3QiwoFQnKBejBKSbZnHzhYMFBd76tnEJToBICjY+
pg3xQ7Xb4rOee4Zn5fyGa7KS/GzJ3J2d3Z1NPVy06pYizVgYdadrrMnxZLHP7LMF
gigrr2uCBSlbCOd9WiDpb1OYz9fBArX9vtZ8ungYhT6WDos6JzHUcdEA0UPpKeZK
XHGpq9RLAooSMo5SSb2VJgKHi58edmIkfmbHsLc+Y8npm7H27DJBf8OkICds50JK
iEK4l0Z1Fjl6MzwlGk3wxYOii7yIc5gYAK/GaBCyjRnhKinnB4IeabMzuMof7o5C
y+iggWiG9VzHIz2+qb5Yijz9jkyZxP6HRemi38RRPrJfl7+9JnfnCUd4d+s2TzPQ
FVjAwJsazSw4V/x7hc+FIddoMbFS2tU0bl6W6UJDKQeXYQOUHJHORXNvSDOvzPbW
EFIFsTbhTwmhzsV1DWwO+WI0UjhmSXnZJFa0h0QZUabT3vlMBJXR/+3sxjeB9Txl
iv9jarfj4M+uIWfsbRv9OE4clk2CXkG7FfYjWbazRtO6HNF7cWsju/6U55V21sJU
GOOcw7qUO88gYSm62AGcnc3DASwyVI7XfXGGpTtVqP2lkzVfF1lFIs3/6cIxANTY
Xu951U3DdHPKel8zGC0bfXYf80jZq4FAEmUsELp28ozBXqIuSkSgjfVgMhhFLFJ7
vnZW8m4zB4xRPYUdrAT00BEAjvoEjN+58cUUvHM1J8eUCwMkLwSr8lqHcj4GaY8y
HQegWvSTNjDe+e6/YsHYYrDYK8Tqk5jnDTWS5O3JNmYw5byQqb9pOJUrFGmp/xQV
LoreDPPOwUTyBu00g3JLHOWjDnrXSrOs8L5wp8icvHTAELUKMN1LGcxRiHLdebep
e/s7tHXjwRCeofSZ5/UnY/oyTQVXFJqusiITOM0jZg52sBaxzy+lmv8GXensT4bk
c04PEV22p1eq72t4x/9d2AYPdiW3Mq+464wrMEQXea8Er8Y7S3HmXdZMkdqafB7k
BBOPttYWNjpwqIRyETN/Wkv41mGICe+rmM4KuHf0mOyRS2Iz9tV46heu6ZP2V3Lo
Heg6lOzKdizXBW8IbeUyGA/f4kCLzHc5e6zzMHwesBuVXCblla1gK7lM+ESirKNt
bUeCHhH87ntGSo4lHocYFThQV0KVirKd48nvEjTOFNukEmyPhjHcsWlMWPwUaIcf
Oa1UjTJuR9a1WK+GqkEhHcYM4GzjisRn4XEdlTs5IZqWvpw0tj+u8KR91AT8NOFb
NnKr+X3ATo3E2vH91Woe+e3AzfQRFK4XH7xvRQj4ERR8uImmn2iVqV8gNJNFMAW7
NRpwyHqQBJfFs/HgGmYXaIAFyS42zfKrkBN/aWcz0eCPfpUxE8jVQvOl/CHLpxWH
qeNhumSio2TFFitQQRgx6V48z6WabQ7ytI5kVRqlHxIqMDf89/y0qJw/RBcNxiCS
e/tISjZRvl+S19VnRbUjjxOaN73n1TcjUUjoRw3ibY5qJSImC+IuBT0VPnqy8jwq
FTjLGVgHdXGJN0YMCVPuahCVwz4uY64WKf8TZC6LfNR6A2zHepBQ3TJLPirkRYY1
2IeVjk3wB0+m5Lw7oJJoYG6rXBefXiSSQ8pTUAYSpwRI5GHdtV/M3BDamuR8CjsS
+WwnpuQadHOyJLH6NlXEFK6kSL0lobThtfTUGWZOXofEGOM3o3hmzGmlfHkSE6IR
99kvZeupOqvQE5Ln7MYO7sl6u7BZikx76wMqsxnttMDFe2E3jeOYHlj7qabhGNOa
Lk7eyHD7QLK4+o7HCgobCo8FzPPf/70hhv3oRxwl4AccPsLBGrxJYbLtZjQ9QXR6
FRFcKVpgso0vbVNfqo44AzDEv5CpZ0VgpkWu/kLtR61AD9KnUX5Vy6mi/E5nync5
CwphRDx9LN2BYisqg08l7v9Km9DBwrY3q+NferHeXCmYLycC9QVA/Yto62SO/Pt+
UEQKVoL8PUwX5coM9Qe4h8FeC82xkwo1Z0/04yH/bVgzYred6zs5EMNKBKjhi6Wr
wua/U8VMurBgO4ukU0g3sgJ4u+4Zj6wTUkpEpCcqbrjkxVo/j40vUmC3a/saCjTC
qoe4RXqLeZ4HzIkH+3fNKw0zFjo2OtSVcTtKGi0j/+pzURtux4m9Kf0i+0+TWiIE
715HjazHOz496rbd50D1W7hAnDBJUz4IeClQS0PJVYCz7LSV8sg/HftAwaQVJngU
CN/EtdeLVIqc1+NsXSQ5y+jjXympe1ewWFogJ9WawJXAqFzKv6SxUkLkBrwlX1rL
hKmRRBJcn4hnCEI4qmMPNbQ/ZFhG8EgcjrdeRbTfTwuDzW3w61Cun/KXz6LBdbHh
RgZ8Qv7+XOxSw1hp1SZfeK4SlACF+OS4rA9039F1Qz+Us3tRIBB1TKQ+g8oa/+wd
OMEFSb2V0qBc/s4z+DQbb5TUE8/F9iihzJvuwpH/XeXwv2IqXkn1dEI1Vj1DIwHC
6CeNmTwNu8iHAI9339b/1ACKInwqo/JejYxbVgHS/ZiQur+qgbkEIOBtsJWc3AUN
uxQajJGmXv0xLRUNFJ+IcxgAs+SSHVsWcf/yI59zlLoAY0U2F+ripoM/VnNdCnGa
lzG217MPR0MFwk8LsMBNxhZsaq2ljL3UbTxcA/l2tKI13xV9ekvsY5nROWU3OGbf
+pnDwkaaPTWQ7SVTR/nWDev3ZVf2BefnwPRTuuVVNDr5+HonRikfhKaTg2KZHYE7
ki3qDUUVzlaqxQzvxHJI78o65SGjQf7QYzHfLizi3yVr/tto2bQlb4FLlbtKfsGn
DSfF/V8emQVMOO2XY5lWBFOPueLMkqDMnbx8Wcd9JAeA7CLIjafCASyYv9T7QEu1
LcKi5n2ODmfz8gMjrEVZsJLRrqyLe1L02WfNVLtObTu3j+98Bxy76Qp7d8knS/rT
tP8mqQrpYT0pc8RwCvxXsBpwcLtwxGO6aJdMm7ceEm6VTv36UdWKvFIEjczHxgd5
diHJ6kMlnn+Dk1dJByH6DHs1edDgVkLfHVzZSdzl6yBYB9McWIJf2G4AtwktT4Ow
Jh4Tj1MHeEY3qrY58W3nET2g6BYdzQSXMNi3YzclqA2choulNrFvMug2TMf5cIYU
cTR+XezriHoHxfzTmVg9wPngiXIfyG+z4lIzSylTZhM+7mLfYeSadU4llXWj/AJr
0+u6qMWUCDpkMDii3s2OS5j4jfLbQnNoQNV7aO3mwZSD4J42yuMBIyb65xGwTCSm
APQ7FnRh0rmPjXE751+x7cfUQ8wiAOgqANogFaeEjozfdBRqGeylotCO4iuL1D1y
LS7hHaOubJzftKLM8Lmrj5CaZ38sk4qhsC20nPwS4084+OvMz/rDq2uvFcL3/r72
zMU35CI1AWWsw4qShemXno/MxVoKxtki0L+eNdbZ5dthBvA3/lZWBJkhQRkGZdIe
AEdpSteSKlGkDXf8f3uEZ7e8E0BUxN13ZDdOKyLsLSAB/ytxO/XoKj9PYPUa6sYv
8pNv5N1zKZakYDSu/9lu2eM4g3+UZXL8kgxwPckcJL0QiSkKlTBf8dM0qRnS+T5x
UJTFBqqkPedHusqI2wKvpJjYKARPKs9IIKLHEOMrTeCqmvyfTKG88zDi4WRaT1Fz
WiTH6kAUY7CkYQIcqm81XtFQFdDpQv3rVZfrnO+Ay8+uUaywWPAktx7AAAyBQG3K
PmkI+D2KhrRRNBzQOvtEqau1S8oa++Wj1IoQv/736WjeUMuXaOG/A4dxlEAayJgq
3RlMFsygvaOPtcGBA/KXV8Y0PyGiNkqjqFKzVO+HfBcmaza7w/mFErfOTrtonkkF
wnUsndCfbf6r4elXRMfIJpkVrnxiWFukZ50XjKM9iW9EmUgWON94GMPhU0qKRfAb
lhN7xTZ7si4q+Fy2AVuvzyxsGEDZTMEuN33S2aahg84Nx8yOJHT3ErbcGBBgeyRW
wm8//WVsp1dBkm/rGnPJoXIoaKiesMtN6PJ6ZNza1QC2xmtu4ddxiov/kcG4I1Z2
wKrlXWQr+U0Ip8GOjGm2XHn7cUVJCr1vYXcCENfAL+mPucBjzOBrydpRZOUFoRVO
RDOdHwYdP6Vjc7tqT6Nb96oDxnPA9UUdg9hChAewH6aIfuBvYIAkpO6wA2ruGRb+
38/rTrAX/F7xKpvyihJmqTrlpBumFlAjGZP32TbFVLrnjMK4Wzl+/fNNA3iPEC/M
38nGX9wLPvG5Qkm0ySo9Fsx8HvslVuWLXTRazrykKK1K+k/hz8+2rYrbQ6gFmfaM
sbxwN/UDK1mLo06KGwTSzgj2jGZ9jUSUAOfpZ5zuRJ23Auwk/iPKmuids0MjSopD
iGdkJ3/jFq/m7P9Z4H49tRQBcla1Lxwm+4uiq5++QdmyLu83p1ArzZ4KRVc3oW39
w+SgZurgpkeUNShlq6qe52a50SBw34afU/ZbyLYZgtFAYAxqgieclCh9+oFGUEy2
VniE3NIkkdhbxkSAhjnKYeCahnLzcIu3jF4uaNaLwV2OOaKV4WbY+jzs8yISvV6E
OQCa96c9rjXEStdr48SUvxm6Xukzs0VLT65W9jdOmkhlRKn6Ji6gqPx0qhhqZTmL
wbuDCmulM/f9gm8hXOeB9zkrsW9GjIpneimzStZaARKJb2sLWbPy1QEmx0m3gZUi
Mck76+KzLDpQGp0wbqPWyUSrEPHtgRZRWPJWfxwiBuv4JDQdZZXc6UVfEJkGdLRn
0mwZkRXgtdJChR8LEsMlNqF/UVvoVkZVJS8btzDNwbFv0ZcwekIgMz51+r8AW1Bj
DehZmRwcegNP88n3iVIwCrvzp+0QdpfhLme3m9QZg5H3ptg413oISmMEIN5ObW5j
g3K5X2Y5uTOocDmXLeTA0f0i3H0E4fciT5R3Dv33EmG3LstRbc63KtI8yhlIPwc7
UTfQbFxUj35i8+CUcuD2kbAfeGIFuHZASIPljq4l91AF9SMBecC/mCaTE3buQl6a
99LhUxLCWoBQJ3WiS2MwC7ef4s4QryS5aNsHIywr5XyjW/iwx5k7vwvNqLLCK3Cg
pPxuZdnauMoz/B3VgT4jvTUaqvueq/+HpMczbeR8JHyB1l+YIuljApfuN9bKv9YN
pG65nvtnFUKqe/2OVMZha8/SyJGNTb7ErlzZUk99Yf/HIuaU14XKv5gFj9J+WuF6
+KQLd9BGI8CcoBX38fKy85ZLK9XkGPD+wTO+4tr0KdIoTHrgk97bjNX6/nf1zR2C
FJKlZzHTLQuuDKRu6PzO7KhQD9kTSUl++KKZHFYExlmudanE1vUck4fI78Rj+yMf
1vUu4OqP6OKeTnDV5W76sMoNrMTEtIlvQecJnv0v9iqWnPC9LaWkaaVFeRpAUraY
CVAUIlrg/vG56w9bQwLDdzSifPtVF1ZhSaerceqlVPBn6zl4LI0EjuamxXy/iFJ0
4dRLpDSZj+aVsLExfYvBVQxzciuexRIEB58n3d3e2v4wXRpXRXHR2zES9axf61Hp
Hkk4JpzAz9l6U1FaWl9GYx44wVOeWDq3MUpkMAKzR9bmkoas/+WamYmZfQTG98Ko
UGAwjeGLYKhfiIvv4VzCDjgJn9+3Gx4HgABWfYNHYiBfRLyFcYBZAZSMyLM0GEwi
TphelwKFfJB6T1qtBFbE7HX/79ExNSs9szvZo3dTHAxtAkRPBK6p6ivD7buA4yjn
TjMwYZVS1KQPz6+m1VbKc7vbyyv1dmo33T2iM2SqGAZQjGCfqcjKYlmr4yG8zHED
/Morypu24awkbWbVKoyZpPlJM1kGtqjcQAsFhv9gxSfMCDJUjDUbOczbh2r3IzNy
yQRbFOmvg1VBeYjf4CgWMMG7gS0OPfFfsr8mWHB+9vKjufyOEmwb0WJNonv0IW3e
spqgSRnlKzgEP+0XASvxqEw3FkdouzBkD+sSnnAw55S9amVoRJ8Bk5Ds3kZj/v/G
sF9xujbUTHckU9DGk2POZMCY73kiPR/sRmsKju9/tw9kKHL7jZC5vVWDkfZIQ8MM
7HlvHYixZmY1l57gME6l0m3yD4Unj9lXL6QGN4c/eFCkkGQGyNwa6niwbH7bwypk
8GxmmQOpwymOeMWyNMpbqLLEaTK2euCecxH5EAnBr2cDfNfb5x8Seup+ywsKZ731
7HSRw7p3EczRzUm824AgpvP57t6CVagjFGBVPbeecbrhk40ZfEbB6XHDf1GgasO2
A4wyOW5wRmgPkwMsT53kUUbHuuKXfEbXroj9sg9eHB+WKiMOn9VONt57TjngdPA4
yunnQEYecAsSc6fCXmfsp5S3mUEuGsev1QuEblxlBNoyHwOQbsFZk62NrIpBkNsj
q0dS/sQT/FGH/ri22G5Ri/mM7naNGgGbFBYYKQ4m7GUWjRbISQfyoyjUit5ALqFJ
y/8kM4R1SLv3w6P7faDwmbzJe/BEhNs7Ych27uIzoHRlzmofqIq5uGVs0Ui/Ts7z
DNaywS9lWDXFlDBoAogz6Z69n9MPvfPo5CqN7QhT4nwCD5crBQ2rYsJCtixJSFUe
xQVdib5S6ny8/kSgtFy337EzfCYHPRUmXGwHV3mpKsLE66fVBKnYPOZyArdUHfwu
NaKXxOx7dk1CFCGQMLPSEq+t3FV3F94M57zdnfiJVRQkGqlG+rwrz6jWrQob/UGZ
XzKTrT0CQMWkdrPYQBCU/9i9Ul70ZXTC25pfh2OaZiyXZX9u4PopUVXOj0Ft0oSs
GI9mNXrGY6ELfEq7ygpqgPUJRx42DY1xX2JAMyqQ1YGXBmRI4jlBNc5B3o7cGHPi
FLAfDWHiMW4ajHT4HW0oSL77GXgCK5c3EmeO3VZFtHwaqWrR8DssrFw1OOKECezc
lpZJ2pedYd4ovBnMamYmMOdzTDK3yUgZxOT96o9eIHJKXBvHYfiVpQftpJ1eQV2V
P61s5nQ29tqulSgrdDFVtJQ7D0lCrMzWS0SCNn3qrITGjkagB7Sg4JmQd3ZA+/cO
pIDa02LadOz/dG5u4NLasdjvMUZcQDeRo9XiIm8IGLSN5aziSQlt0x/gmJlZwHdh
iRXqROBuBkUTu9rK1QLYglLvi/cUwQONnkiItxFxRGuHmYOJLN0xyvSRdfBBX5d6
b6HZKU/0dMfGAYgvISPpA+ejweQFTy00mP+ZkEu7eAKnBwOatyyavHqitcW9vJwc
lTQq9ByM8NFLTUPtHf4CEMGHOyBXhe7BscMFzSvmo8VLN6V/A+OgY5BqgsQJ29J8
3CPinsBGK2uPnI6dp6/bB5UMsoWqc3J71A9sFD90/ymiyyDDf2kk3X4b6ichBziW
/TjcC+85F5efheh4akcew5RkRPtki2KFjdNqHWMr76p2KwQbYtu9131m4qGTLb5Y
tN+VpN5QoektNqhvBJwBMX3m9BP21tjpuKOaxxSI8jkxMktkE/ID2C7rbmQ+Tfp7
tptR8Z0NVRG18/7axmn/NHvypMmf4Rr314KgzRyKmh+S9zxYqmsv1dwDkBtKhKFq
SOYLzeCSh6zeg62GSECuyI+dLlV/dQCadyViZv9v66XAGZ2yg7mpz7Q4h64f7Eet
9Wu4GiAJ97XqJYuMbhDUkkgknYLxgdXK64wlfdm+/V9l/5qizV6/YNbqMolEBPD0
0z5zH4DV6ptMlkXALzew8nia3/TAqHNzDLJasVdec5Romkv+tOXpuxRXsZwnFJZ7
HB7sXM0S518TZSzpDi03yb/ss0tNQ2UYVfpNsgKVUN5yDKThx6CiO1FTlddmUfxB
9NdKo7MhxZmXicG+d8WjUeQ1ALHdEV7LcbbtlkHOp43p4joguQLTR56GDD4fiOZ3
OeC7zy7jatGej4KPmB0B4Js7eUx3v+SbuCZYUHB970gpTvSnDZW7WCD2gXGd51mt
G4vlcD8xf/4Y+vs8h8BNIDXNwI1CSbq5yjitUqMvW0zRx+itDiXBJPBqQB6dJBaZ
Od//uE2RrEelovV2l+OsYRRdv/6PgjaSHiLMLWToh63QuXQ8p+rPXO8eyTdBFP9s
BZIS2ifpMnZunN201p6UqG1bFKxrDQmmvsE7LNU31Oc/lp627gjVFVODg28hhGXI
QkVTrEgy6sHmJXfg0lSOhfRr3Yu0+eL+L7Yy2ejqu0q6duSCsOrwTB6XfQf88Nis
L20xhZlmyk0JXNWDwmjaQ6rBDF3ZKp2OkgEKbxQ3FytI7fvOEU5iOCMjyYyzZbeU
dGr7WqIcZoe983ZIol2vrFfcMgDjyHeTrbeD8esFbx9W1Kv7JeLTHdYTXz6mL22B
c2s2QRqQYKZEY2+Z0G6OX5V/lhWax7sIluqPcm8nSGstejfI4G1zpcpv+z6NXNRv
UANBHjh2UiLKwbhjEtglnDsAcOT9otFAy05P+UJGEVRyD4j0pjrt+MvgUCTwtU8k
tEaPB8XuNqTh6u0H60CHeGz+7SPJy7NVzjwyzbcM18+4Ca/twdcgH8y/uo29L16a
FQWXJOErZ2AbPpQ9tw4ITtpTmNadQAOZ3mzm0fX1QRGODDiUdXoUVzyWScRqJxYF
zeduv9Rxw0KPcIcDWD9ifOvlYt95kPjqsfY5PiGElwWg/oNgq6YKLkZihLRvXoMs
E2PvvC9XY2DErUC5w2vpUPXWBtrsJsMw4eEurJIjYs3jwgitC1t187Z//+IpeWy5
2rSVgw8ztYK3lPuPC713X11/yNbM6kq5OZJpqxT0FuqvN8W60c/87kGebyqEXiX7
MAREpxnWfvdvI7FXsTv1gCN654tocgEooBAV8AIxQ7JUrF6DYCSR+moItn4j/J9Q
pUII1rgBqNaerV1cdzqD0JeD1dYooNXPkp/nbPgCx2PRhqoe5kLfni2zYSWSdfWB
i0SdL7wFHZep9rKsQyWj2H5Q3AAOEpJSgVc+BvLypPiWzClSw1AaZNESLpiB/GzT
4DYInT5xFnTPt/EWMLA4q6eYtTP5pQz8pd2oXPS6o0D5y8k07Ebtr1/CIY/dhiB6
TaYKC4ViH4VBxW/68RgVeKZO/mBQw6t/aA5VMAvp1PA8dxzrsS7bWgpaER6jNcjX
DbqDssf0Y++CqEPkEz2A6oK5jORn07lgK6RTGpNgqPEwXUztsa3BWgW5SzWufhDZ
os5uIoV672IsC6c/ZcODCt+j6Am5Xj1chnjb3AGTTiifxfu+hqy0MhQqD4m8YjQ0
RUIpIf/mHBhgv9Ci7UcfHULuMaW1dr3BwpMukIMDE07XYr8uatMCAzkOqvkUafOz
3EIEFmKzRk44BJLR2dM9nY/KzopcTSonv80wOS90kyc3uElVN9aJrN/KmhP54eGP
7VdJbYvC3Ht/ZReqeRs8qP5u9t4ZoL5NDuOJheq36mjMaVZDQz9TK0VgHP7Bv5qZ
q5kcF4VfRzuwR+1dtX77offG4e134GZ+MBHyzzAD9hQtmw5J0SWYfT3LwK+JlE0O
zuIadBywUJhQdcCNDqc5M1hxPknvzhGiu4t9b2sSd3JI/dTsYcmXsdoGPy7ycXDT
icj83VfRuUobcdLHsMpqou48W0sDMy8spdTT44Ba8E66MEyN19XYha1DcAto2Z3v
+yIVaL77Pjs2sgjWwfq3AL+4GrgZDQ1M2bF2fGeIGmR1hwp6mLhMEoAqYJOorHJw
OMv5aPpOl1xpgoovBnH9UwR/jcqcPhICydQw8VYpfPauK3VeoAQ/22HnXNlAq+bn
fYppt4+oH981sNN1XYQPsRoVAIwloRQuZ0nQOyocLjHq3e8KHLVetuyi6OKqKe4m
4TVbRt1IKk6FoRas31oxps53uACaXgefi2Xhc2v9LgTUSLef3ihFtNLwKF1iCgXH
b+AUoMilbSrlg5eh0MoHMJigjmBY8XXqXZVXyI/LULEb/2xBF0/PSbZgK/S3+UKx
QmF3B4WdubMtof+PjL1F06fb+hSdMUtLN9LM/NSApKP2oOK9ydGaU5YSyQEwJKxg
sPkfzDOpwGxC0D+WQ3bRal3f1DX6YUZHm9TtsZn2stb9qUy2UBU6N+Y8BoVA9XG6
6goZzN0LAFT2LkvXQqxqt8WL9+GUg9cEnWzH3Ahg3G5zBJwDqQEAfvrJDjbHOgEN
T6mhLUwtIcCvkH699zKccKWCXbZHy2LJ/Xr2+4JbNJiWQNLp7VFFIqMb1H8jb9Ub
DU1M5zhulQDxSWMjq6t7NxVFnUQkCpRfdb/s+ONjTnLygGn9pI3EGiTLF5yDa3sG
Aa2YDyAb6xYpL1oBpF3xBNQuhqqBNrMyiU3fpP9VlwFXNpWK+veTZ4l+H7F4wlXO
mKKC7mJ8e/Qr5IOlTdwCwbnqR522ipP8WB+zwOyVwO6IiGrb/T6c9wHdr0pduZt6
pbd2p1A8Ja0U3W1ZLboBf2jIFw96m/P7WFQRLRWtneM3IKPUysYFTCrjjdNvIyb/
jK1uwfb42u+dzCP68o65l0qAQhUO1LTR3vIO7JiD1Su42Eo1VSRvxm1+IY/etWyW
OsVr2y8FGRSlPJGeVeO7K8vhidBsYXGHada/lvDPmwF+Ka75l/96fthhFEEH+aHE
O078C3wV8S5pApfgzR4lTSNTFbcPg4/WmwoZTDrKWgYAnOqk87Ne5VYKL6CSI9AB
uSvQw3VPIkrqWS2JIMxpBngT4KW2eRw0nSXvJ6Vk9gMexfNUqYfSQ7tzADF7F/D5
agG+HDxxmUGnABomHUEqj6C5k8XCvMP5h7cao/8+APvJP5j/8lwMnj6p8++FRp4x
3Imn3PXHWanTpbQ4MyW3aFLGZwaX/ZQ4QNg3oluJBKQd+v5R1Vlif1znQcTBagWk
wcVmQyN7EgNMpnjGkGcoxupcPpAo3KvwYZ2YD4J/9HHQnUH1FgQA+g4Q/bDI7JQK
ufHPk1SmUis+bjvC43r7PFDv1Z5sGJlGh0iyXyh85D8e2I3zPOwjzvCahHda0QQo
EEAMZDXbx10znz5C0B5hZ9P7gyVwP+ylvjgyVpqcVimyhJTLaF4rgOSBzukn6UB+
STeu79gtcMZ0NStSwnBnvFo/uJ5+KyEqtLlUAbf3zxpfH3EA4w8qPOTBZE6JFMqC
wPUvC29appckNo0tN/punBS4Mz6KIXG139sz81x62jTgUPeF5VFLNHdgqq+zb4yg
5bzGBVZi2sQuaJyqZPcbymEOQU7JYFzCBfbwLSM3pdtE1q7uwp2RQrXdGFnc8trP
lxifK35NMjdORxhPjdlKTR3gZvkKTxAUDmn8lZM1fSy0hY8dETMNxrnd5eDKkYqc
tXE5IJWlwF6zQ8ugQ4t4CwEch+GZAZFL2tEmhuKI5rjpPD4PXgqWxR/uStug+gfz
lcRhj9GQydDsXoPBpqWzd6dOvikUw0X6VeR9SktT/vGx8i16duOSsuZQuZr5Sz2n
JH5OVGzhfVUAGGl1GEnVqY2SmSasv4ANj3/zuVDMT9/bSUEksqrLaqrzVNXQrqVs
ooNgjDIwzlib6MmG26OofL8netsn72hKek0B9RcWiyYHCrNaZp7tgby8RuefdD0s
fds5qbfA53d29wvuhMZwUnMjz/dUc/onAxkg75Bj1WFZrytRWHJHgHAZEHKnG2TU
GpSNUYPz+qrVK1r3bufSfaBFUaangfbfr3LUhuoSesdYxJ+UEiKmBMjtE4PbCPGZ
YQ+UXBHrFDMI094N6ulJhUlwT30k4W+jzfoNf+if7CGGouk5+kjTVJ6ym+Mj7JN0
16nTcHwHn9dm71I4cRxgsBN96WDya5p9y+/shpH918BYI3YztU9XcrCRx1CIQ42i
2oTqmwuR6L1rxZ+79rxmp6ZI9G1de2BP0qqCXj2QamCQR6kvn8gGth8sRWr1fUf7
2Kc+mrQikkSYlZ6j4p4vrO9NW1d0H75o3aeblh8YAbZtHPXsImW+ExfgMWP6NTzm
NFc/tOnmaJir0OsN7eeJEWQrnzYyC69WXwxeuBxHwQl7F1oDNc5SOc+kqbCO+EbA
h0HLl6ZEpOpt9rtRNGkJK6wEP+/nRCa4XN8NMivbVCxLKaylIpzWIcVIW3Tv8Xrh
eQ7Jf5thwqCiI9A7aECV0kvMdXWEfiYXEqROyDPhqf46sOGT57WL2+cXs+8/vRqt
+Gj/OjJeJglDL6V0m5+jD8yDTHeZSUS/vrVu0OOLpoXUW3ztPKSuioZQvoKxh3t7
YCG9a2rmf8DWSJzJIx6B6uAgTAEC56SZp+ftNQZzz1RQnfgczNPQ/ydD9WqPdbXt
b5FkTCT9JpOGtBTj52pRYUSW2mC4ErUW8YLOmYPWHqO3KzXZKb7G7cL8hR3//syU
3IHZsUU2es9H3W4lR4GE1SSkbtSLjBpzHUM3hxLQ6At3uB9U8a4JVGm3MncZKrDL
FkpbtgrOgw68AO3Cqh5JhlIBKgLdoh+5ojZ5ecPA3TX6FUtLu1eH9NbEDsug2bBe
LDx5R2cA5U2JRjF4VuUiQnkYIn+LjZ8SzRPKJnnl5ehO/jYd+1pVgPyHL+NLCw6W
PixBrpXZ8/UhRfQwFL+GjlEC693OAn51rAhhTmCfU87+YwZRd6v9Ph1RDl/h/03K
negEWwgd1K8waECkW6uMVAyLkRSoebLbf6RRKGcHQFRX2Z/br39YuPqL0XbdYFGu
SHLzgMM/RU5viIZgZL/Q/mWrg7dmOXoLOQUM30cUhHKkgqwnO2lSe9pHAGQ7m+G3
OF45Jo3ou7KfRL1yhmF5GgeMe4msNzkCTxdQAMnUVphloNBxQqs+1f7AdWDEvNMN
OFmPErUvOKc7JSBxNYl8vIH7903vRX4VrVTfGrZDtkc=
`protect END_PROTECTED
