`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5pKp8UCBNB9LGCOUbE5atADV2KpylWaM6ihKuxUHr0fUy/tzSf4bW69wFKCSQVu0
efajTej3JJi8a8LVFyBFC4lraPOp4Desrw575Dj+820s9ypp9z1TvrLXa62mITup
SLyKpfANrgPLlrneMHpOKheo/gnv7fmmoUos6u7VelesK+xsp4PrkAzqpPY3EPbf
13jcBZidJX2S7My1BOcR59VLGUm1iFhazCeTMadmqjMbq6iCicIW/BJW0eHV+MOt
g/PEeV5MhvxGVX5mfAHQ9RQChgs45ICLi22QdXi3hrOiap+AqBFW+FwqbVdXPds2
MNws1aKeERjuWPPJWNPuGr8c/HfjcWuMoAMtOuwVNwwvWZMRzJQXuAwxaT3AF01Q
wpiHZiA5CBKpUNUljRCv+aChQBF5mQPNUzyRIkNKsr72MC6bk/e9fun3XbGW/qhs
IbI38lwt82iEmUgWYT5tGnST+uHYAzflV6Zvd1QHN/+DR8O3/Ak1KcM6S7KdoMDa
U1kI4GjVWdin//crK/1Omja9bEjYkPxXbT6xH3WjoqenYuR1m9ecwvNeg/LQs3zs
BSeFR9AlRr9dIMTTKUfdafyyO8z336dMjlZxY4PtH4rB2An+/UkYtg6xz+Gpftno
k8Zfo5xFgmZGq/kXYlUhjIvAjcPKYRBqpUzLG9V34TBIN1e5PFPT3UyYAqEjEaFy
`protect END_PROTECTED
