`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frJhpnoQDkmDFzFD6X1iappNwCJmhD2bA55TaqlG7jj5xjUWd8xwTQ7I4MDfT2Qy
pRHWexOSVx6VZETpMsBCSuKbW8N3ilPXK5I1t+qxNcja1tB6aHjMwVKWrBa2qeRy
CydlPpXrfAyhH0o/VXjN+9hxbLeKrVw3OP/qs6bVP/15Zw+OMGj2DqrwqfhnLfZW
/KSdr3Ei4wQmb+LyJyXgbm48+kQaKphrdPjSTSrusU2yUx0HkCKAQKgi0p1F6ZDb
lqDph6WSetuj+3ECTXuduMZkt6Q2lQocHyTOr5MLbdcRzQWMtzaQGRKLqKEJk8np
vQFQCjil8mz3rW0PDFa2fl2Hm6VXKD7T4nkDPaxl503FhtHpP36zm096r7XHsI/V
pzgY3CI+uSGI6aJPna3ShxwE7s6UzYKBmZuKzM0Hfxr+Cm3leJami/bV4+1lNG8Q
RE7czdAiuuQLabXsLehoYhXeeYUmF7i2flFrCHcOV4sVSBctWs7l/TIT1lOCVa0k
R4xqClxIBwDwkH43wd9+3hNVPNcUmoRmz+4rgDSg3pjk0rTGryInEB+show+Nzuh
J/HtZarrP9zrcNGLe1U755wGo/8OMIjnAzo/iYCoIVLOP6Y2NDBFwqgaR853sIcu
ryjOxhYcqsWLhzOIj0IYgvPcSUAmS7Vajd+HHc4affW8hoBUPm1zevU/uOTUiiDk
VStEUkOSgw2w0MbxmcmvFFCiOU/zDj7yD64rRf4siSyxknDr02X67y0jFTPpalRl
1O/t8FOvzkwd5hYEB1eTPhG7IgMfT7+roe3fQIUran+/7ROz/tUbgf3TEE0L8BiT
kBpix+RRWlwltuTNobJrxGdUh6miQ6ZRPrcXqTZP39qWo9g5s+2ne8AvnVVYE1HJ
Ek6WHOYE7cmNnb6JfpXLGt7ZpWE0knvQOPqERgCYg94eFHhnA2rcBKdDSbF5O/+s
ED63cEgZJ/TQ3wPTZ6llHAlczmusUxlRKWjzmpPXVy2rgxoUmKwOvj4YstGh2wUL
3AE5qbZHYd39rxnnouwijtm7O51BO/DeSKshvGaDQyFVRvNcBiWEg3RYKTlGAtxZ
L/34/b5H0BePpS9k2FiU17otPX1R8As4YGV45dEkHODtqXOiv8M6bKUg+QhtM3WJ
0V7jU35dVeDwvTh6f/TskVHY7r4/wQnX/xXu+ZzRUepMV4Hm49q3rPGa8otDoaw9
yMLE4O3dxKEXEMMYdj4sTiltNDRYiA+zSUsQQ4BiWXIpN1DNOSF/Ws0zjT0tjkgR
ZpkEXdwv0wMW9655C31CAGxpMNkC2HPls6aF5mb2OzTOZo8cvHnlTLn+Ggu3oIe5
NAbaysJf/FRtgLgWchHkxZBCrORk839G/COwxjZIVezeJQ+HQrTFxKdoy/864ciC
RvqaMG3w5ifAx1LMIn/AnscZCy0stu9l6PYyEudDPbay1lD/NQf6LGV2fLYXdwbj
K2EerVxLywfPy4XugVKama1kHahIWjZho7uPo5HU6XtjkAVpHLACHwc4hQQWxYxI
2sg+SQmDnUpQVr7lWW0bE1Rfe6CtAjpWU8VDOpnRGa/qiB5zqmEOyX8uXloIJQWu
D7izziWLlbHcTJxY8H2K2NkTn2k9HG6Svea47ItVgHF1UqspumZpOHF4a/HTEXGP
b/vzamCv6G8hJq7jbvtU/Q==
`protect END_PROTECTED
