`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A3k1YEQ35+T9xOAbXLhdLAR/olJwqhGQool9PfaiJV7b2GHRPhwJP1iCo2JRpvI/
NrPAO4spWUKio4oLuuwaPdmgzc49LDSTrt2h9fXs7kQp/MVeF9kK+wOhqswfrtQR
H6zewBKOEHfha+eyzDnigp42L2MASxIDTEeLVN+8TEjEbUobfSUKlE+uEdkydeHi
b1L/Mr2RHSOaubHTvoL47BRxYUs62+Q4vTgZZ3yXDGZyy7ShNY9a+GtVS6vluopk
05+FuozDVhNf3aKudQCSw/URu/gaWxyUDCxHVApFgDYrAc0gJCYv8Gv+g1/95ny2
RKhzSJgHne1VRGyd5CPRiS752uZMMkVDzeuDzKLvyED0H4i7oJk+Pn2wjJ2HJHS3
6dhnZViHyGVjd1qmVyOUBkNNehKaIsyF/OIKwLcVTtqr23DiD4W1vsvyy1S6WBTq
U5GHG2zI5hkR5nQiYoaxDn8oMUyhcfwynLa+5Df/O2VrX0BHlLjd6yiu7oNLKJlF
L1eFgMWBKxN1qgY1Ozr/oIVm1gIB7WXr+n4uzwlTYH/tALnsq1L9kAhDPH06dKbT
6rSGjb/c/7v8aFkdCXMSyO6R2bRv+kQIk1ZTPPbc3CISAzuccDx+iC4tnOSUb/80
wxrCKA812qvyLvKlTYKnl5k+qzNlvas/qWC3W/JmWvamx2Wz8tXBBlQz4PaJTaKx
C1bPh0HRryGCYPgRp959kvK2n7pFlF9Wd+56lS/Q5F1QXDgeYpN+jk1iDJctZ0xE
Mf85Xd3qYxMmh+v7dVQH+eFPLDX//iP4TIlMIl7tCd7rSSIprsOOSiOOD7QaZsac
/NM2ZNWOEREZPeDFp/1wHLfo9jZ6yjrQavz2Nu/arxjLe5IsbxGVcyk0fS+9+BPy
lY28q1nmABRBRmmHepeCnObjh1Vs+HBTVPQzEB8ZM+rbes4T6swQzQ4915rvnNp+
Ifb5/x1oLjNdQiDsRJYB+pfa3HC97MWjiawiaXeumYpHjTE5COusdCEXWAvco8wW
bGig6daRaXt3YOZ9i0dAsE8mSOnTlMH6zmHSaNpJ7QieU+bYpUbXmbJPd9og2Xh6
O7ArI67Ns//fOUklK9URX5CTEzvGwHEPA7Qiu36fHKv2VAiM6nqCauX5MT+QnvaS
ZyK/ejFZBFCbvswsupm8lbCpswM1Ofm5W2QSu62kPx4rBoEG2MM4in/keq/plqdu
pMc/Or21WC63fZdqL2xH7Fxg/Vg+iaSqveV3vimGrZDPYEMFL/LuzqArRnBkM7F3
`protect END_PROTECTED
