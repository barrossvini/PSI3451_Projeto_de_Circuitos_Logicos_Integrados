`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CX3835OVchiKJbU7dVbrL/6vskIlm+nmZTz71l5+0gC8tvAqOAUmLVR3nVg92jNx
ZgnBRTypjwJXZql6C9AzJkVSj/KH+d/mN5/nultd1iUIkoq6HXRMh+YjhsFEGSGM
DVIyOy6N/1vDovyyEFLPikaJ4BHTVl1HlSbVbZ+hcJEASJGSAj7XECHFREchRVnl
NEWE5h6xa6Rn4o20APvpei8ChOJpJaXeSRkWt1YgqWxY7arUkZe1K1DkKBHJqhVQ
Nj5Z+csGTwDhsf5qOTd5ADvVeeh4L9UndiV/i/cFDHLz/shDjtKQJ7CIitQm8hQ2
jdT12HLxbv6/Va3WbR+bjV3oV/i+kbE8Evi+wfDQJaeB59QD2KjkTJBndKQ6KhpP
3ZuZ13fVQ54UDlmE0+9B2Wg/ByeLj9t00CWzZx6yNQri89XwzBVu3air2G1gNzUU
xJBWQDKn2YgGH6FTug43QW9yKPs6jEPYCHXiq8uTPfu7mjvr7y7qmC/PE8AU2A6A
DiVs6xyOk6q+nR6RU6lyagYgepDIRt2t7pgjzUyrSvs=
`protect END_PROTECTED
