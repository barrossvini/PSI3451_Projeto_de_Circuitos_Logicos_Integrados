`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RnumeCSVLaCWx0wSB9GAYnjLsF/1+7EOXAM5pNW/FIygaG+k2hCeNGIDI99WqGtl
QprDIpxwk2vO1YlYxczMCbIk3hSM3Xto7Y8zCaRj/VVFmpmOxz1qDL+3dDoZA0MZ
M9TiO/ZazBCRAPISmlR6qBMqOdrz/FwNNk8w2U1Y1bcyANUCAqVwbJ6W68zZ8y1Z
DeDJIhP7jIIXhclZpmoYHIowH9g/EEGDUMEfXvX6h36rjJWeq6abpqMG16OwgUUz
B8Et8ceSdEjcNSIyZcv/W4o8agNlWZBUkFmVFIus3gr3mpm+B8d5m5gVyqEqLHKk
82KWN7Kkhke7VEL8qgZVkwTd7InX5PR/bDc0onO9K5F8mxSL7yoewIQiej4e+zt+
MbtSVbY/uhhivGqiuSWXNN79jaJq/TbUVsLAJIaAFIYx/xiHecE26qrgFSV4WowP
ZC5mrkkeehN86cfMOHEbGAaUgn7bAOBwKNWLyI//1wv00ZMItJpdweYxCuFDWhDc
+iAdbEK3qR6Z4HbUGcXREDB4lOVtflv48Jrtj1rEFRE/5u8zvgXWr/mSqIBWmMae
g+DyfQ7OHaSiJopRx8WJRd1Dp5i21Zlph2pkeHNZNjkltch8eW/X1ZbX4QUriYEm
+oVabHLrE18ykY9lVujO4XtaL0R3+0Z4yexjJh2c+0AbgMyaDwZO10NWQvRH69PG
5wqoo19VHDd/AvovqSpocd45LXw8HrDFEoq2whRrupHHbJQ7o3SAUPql+pOgbViS
GkUtJA9nV3qm0WRsvxSwh3AawTGGCFtda3WATUoP+p/IbIcloMI+MnDI+aj59QGP
e0Z7yH/cpFRF549h/zDwRnq5CsbHga6AZGsmZZgQbvSDO/WDVThOLw84P7b/wI2t
GZKvFcuLUMCAysOAh+22fqVydk+YZHgIfuZpqEZPrSmROQeCGNEyXVQnDlisiCK4
YvX+T3vs+tISUJVsWum9fny3KBpDGC4DGGOXp3pjypvH6B9kkDPD9jGGtd50m/lp
83/v6N92H7Ar7iIJXiNoPPEqxla4SXdSugeQh5YjQttV+pPRFc0hZpAq9N6bEqJI
ngIjfrrWjeiOgJx/YCYysM0t/dX3pyV9qzm9FUxxmJhAlRdproY8LI7ye98TqQ2v
55MXt9N4a565SVGfK68UjMg5dtCQpIwTFpHnYuYIsD9RWiAi5skUZ22fPVmQP7vv
irVqpdLSKmWuX+k1Bo8r0P0NIWoKZND78RFv2cSo86GV50RRS/WD1YXA4t4I3S0D
XonbskWnwIAE0yErljMzVE6ZE1yUrqUCt6n7J0+tZb0dln5zSvXgUsk9oi3hlWZ4
EYAAeNPrN7iioauRQlQ4dEHM2VKSgoGALLo4hNzBCcnmnCr4UDVTTqi3iMowvi3e
SK5UCXWKpnSBhOi17T2CIXh6y2ICwa4pEgP5l7IhOaEkGodU7Eo9+s320rQjJiSN
mEZvkwvQfSPdL25j3FUGC82Vv0oqZfKOnD8lpOCa9GOZQSJrqZRoTdGfHDaobcpc
K/c3kVWSy9SL+z83UOKpzB2t4YfEy+oNNdP/LatV0CBWtZcp9XYZJhyG7ska2gAm
KdYqo/f0DCBLrjot6B0M8J9afcB2ph92Nux3lcYKrrzIuQmJ0rhGCR8SL6TYpVij
n3Aq/maN0kXj288Y2X8zi06PbindO8sNwUj3us6oVjOzr9ETcscHzUa43x4+YhOc
32t5wKFeSitDjRq3qMPToM4+7pSXtRxEAiLaWm9pnTT9RjjsJsBRK0IGBxSzqwGk
`protect END_PROTECTED
