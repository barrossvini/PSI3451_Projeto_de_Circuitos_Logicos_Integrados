`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ghoIJuaFMJmqn/FDd2Ez3PmYoZ1+BLJsPbXYWzt44rkXy14SURsqw75Ud1Myb5UU
ARBV2KucCP4M6JNo1ViTwhdkNniyrFFtNGd3ecK4/wpw2Hhzn2YTOHaV504CCgtG
KmItmEIqE8DD4qwTZZ5Dvw8JwdhcewRxXsYpEl5lg+cm3IX32QDNZJQx+EsmUZkV
H0LzMwNBw7k29ga7X432Ye7HKBy+vXz9jXYRuziphpVtm9IZxYfWDQ1lpDYgVfUf
P0qBvojeBbqkw2/YiZMx2K7iZ/E7nFNY+vExlQgOjUADA1FR2IA7/s7CyBy1ZC7q
U/HZqtDFokQUKeUxftyotK20ahGEFtAYu9bqSmBj2kgo0WVf5T0IyW+lPNE4Dkwq
3YMqADxk1Gjou51lSpg26pe/UdG4ihJ0E0D/tHIkFToJlqVmf929yWleKIRihlk0
QWnLqMFb4XE4hbgeouToE3PjG0mr19ax7Awp6s4UCbZnyxpVtqR5NwU4JO7+Iz6y
FNP8S7hkQBcfeEgUn3UmKOj4c+bQ28NKh6bEUXKLPcI5Fi0PtQ3gHy3NuVdQKFN6
P5bg7W0kf53hEXhhuc6sTq8rwxQoiWHnVOkGoiPz+j4+hpiU1X3IITSPRcbWNJdp
CrsvCcWsE6+C2wXb5MFIALBk/dHtGAdffnQ7lNp+7w6fdQgwHrnFvt/rs3YSpADI
+MW9hGSd6bTM5lIYIrD74NaA7/vcSDeQaIl6Q1v9cO+Xi0ooduTI3mwOJCW46NI2
894hRn70IZOHt1tzWPBg0bRu8e8LkhAVtz3qa+aiKF1+dmxM0HT+jrRlSRNk0d2I
PKR1fwpmJW6qFnsvZbcox3kH8gJ4bhms9lvHJzcLsdL5Isd5O50ewjCnkPqGL32w
SEtGKN28DLCNZyhpuDpOH2g3AkBn4mIPUyZT+nS1mcM4+UsHKPCfeOWO3tDxSgKP
IgcYFHsFOUqMVPC81DIVoFnmLux5zGkX6bKoSsL6tpoFhnBQgqDGjAylNm26uSJD
qMG11dYYrvAsSNJZF/B3mbzh2j+3/OwN8K0EFRfcAstVMUk3pLOCQe6SuA3gl8wt
N4djmD9TLwa1j8UOyF+9W+ig4ImTrQHQK5bV9BJMUhFYiE7Ffm5pZ/nFm0BO/+Jp
`protect END_PROTECTED
