`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zb33Gv/+g2gmJ3+JsgWGAYOoS8Mh2WnWb++UfQaQC1kf0qgLIHWNt2zH8kVX2cTj
f3jKoEU1rfcd2AxwXT6AoxFZ2rentYx/+10zi+aqNTQk0x95fPFr39OR4qW0Ha14
GYY+pdbUHbPd2nA+ahdP8TChmKNbvktb7mB6X/g8vXVD1jODoG2c4r1nraiWx0xm
nbC2gy8YQfFGGZ1cbg8lfurn37tfCrbcsD+8t10giZ6evKWMf1qH+wN12Td2vxrp
dmn3ssQRPiMYOY1sg7Ri5Xn5lINgpiCiPoztnm+nCMFYQg1wXVtwG8RtDYGsQrBe
C5pG0SmUVoK3bx2L4cgJWH6/ZU7zayfYgfDvGvTfMP7vdi6vvrEJ4yCD/oiPGzKp
6qNQUk1ZG72vBqMrqOEGK00eA4h0/lkZMMjxpvtfbWUX7oBRv6jTyApbw3j4MQHk
ZxxVCIilQUxmsm7zg/KfYRmK5ffVVoo9oAJoguFbUROR1PuzRBfrqP4CfbYA3se2
EHW+DsLc8Rg0NgnL+9KtRBejDMD8UaaeFNSeZ0b9UDmXVvJkcp9jaWHgc80Qlf8b
wMDnd+Utk4cYKzDZLiJTV3o0Dan1zcqeHezkBKHrGGQm9beCIk89OST1MAycB2/e
K+5CuONIq2JrQwBsFODCjSoC3pVdPIgpRBAJP6fLOsUFA3QruqV5eMqxBzDTb60K
ogUOkK93WOTuLUFmcGN7+yCMNWeVaz6e5gGIdi05JriQEQkbrIWDEA6x1JlKrUKN
LqXY9bWz9LJK2AbyKaOmtB/x3l2QD3nYnlGYKDNOmmjTMuTT0PgefwEYGX1GRbLI
4K8+1Q4sKTxfLHKpBh6wq2dktcKsk+K4aG8RYZh2py+cdyMBycrPwHtfNs9C3BeK
qmjCVNghjYNtFfMnO+QYcyhp/fW8dQiOYEWUOaf4DUOCA1ugeeLxUFPa23t7rBem
OFKOx0gnVxOSRjuor+gZpAWC8/xA3Ap71OK99c4K10L76KMVjDxxbNOpb1sFb22J
cO/ZqNiXcY3k8BClJJDfnl6w4jlRIBg+4RNSHwnbix4rBCdjauBJlNGEQajWcuuT
TYtLbI9QzsYFDyqSzBxVyNFTqFEl/GTGumNID8MuAGbASAQQAotHTtNmQN9CdB3r
VmeDtVv/+rjnlJw2e81GjRFA6QLEu37S7nJ0u65yCizPPK9rRfd7SZR/Bbi8GsSa
g2KcHAKdI7Q8nxOq71MiBIglql8tpVQ8bSuPynCRFmc=
`protect END_PROTECTED
