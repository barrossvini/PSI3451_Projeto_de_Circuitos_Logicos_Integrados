`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fjPHcRfuEHdbv5I0QaIjN6zunUVw0EuNiLiYHDkRTf3CbroxmlJ7Ne9A0CBzRt0u
991RnWLVpJ4plxmAt+ZppQJKIlqpxW1QUsw3ss/jARlrCHNxFtRnJCpg/oUAUKYl
L5FrKW3AkH589hXDqgUFm+g/V7+ewKUPp8fb9NYi7txcH5+6uVpqyax85EpFoc8H
gAg7OGoaw5zbGXVZo0y1fapmC730slj6OK0sDVBeGO9AGOhYenWDheUOI98D3Nce
MrU+EuAum1oXDrzh/DpuEXK7YWxImg/uLuqgCXY0IAuUzyFYyYql4lofZAsPuzMa
DKAGestXPkY4P6q2oXrsb0WWhJGeo5VFEqJtmlKWqQtBLbyFoAO0TKgZYAt8Q8Me
pCNw2Q/7TtYyO7ZVx/cva7cLWbNBonSWUR7HbYCKdsCza4D1EF3KcFqjp9tsR1Bi
NGPb6hrZkKuPSIZRkZm08KGxHUNqZQj0tWw0ePm8BiFUQ7Ycg+rLeXEhyXLWzNnU
WfhtQzIPuVeTg/ijLmYPq76F3qqoIVPdgP++UR0f+zRqrRGECkbBaYIuhdZlZAKj
1H6eCziPwxc6gGOsJiIN0IwqDWTw/DAkFiH9sQ73e4YlaHhBlmxx1BCLhEWOYPXE
n0n32klTb9BPZfJWVK5oPoJ34tNOqZlvJ9t24AkiYFH2iS504oVs0gmxVPbJn3Zg
`protect END_PROTECTED
