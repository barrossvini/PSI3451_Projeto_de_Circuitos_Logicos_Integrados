`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mx+mbfuN5omZhqguYF1X3XM8EFOn7W3PPk561uZD8AKH6kcMr7mSw1lGa48LVGEc
fLD6BIQ2AagS65dVq8K8lCSgxYOR16gGBXMSkSDlfjab98MfQCoLqSUSnA5reByA
gzmakB4e8BQK3HrscdqxgNhfS7rOl31oabA2xW4D3ADxbLBXgXg5BcqSXw08kd7x
GIkNJV66kQ9D4ohwqPZAyL7bXK4p/XSioqgwMbkRLFjWBhQ7IaxqyiIIAnXUT+Oz
WAaflhDrzxusFiMfmvDB86szA1pEPJBcV5YI9VsUpuwNTFZ2Nk0mgXogX04UgLSa
spi26fAymibnh6zB57rsd7EvvtZ8keTCSYbTQU2MlnNXLz5Dvdut3+RI86mre2U4
LBrj4vCSJZlO+Z4Hm+lp553vLvzATVATgXg51uuphw7bvturqeKkJMLPShhZQHqK
mS2HmoqeTpUkYA80xAIjySA8hWWPj07YTh9x7rrfA3SC58X0mrSH4EVlhUXpbzKD
nfda3t9nKHOM4uAxdt26yQuSuOJVPCDrCIxtj06sRB4PYIkixj51397mi6Lq4nBx
QNvj1FsIGliS0Y5eBwmkXSAX2uPIObs+mOnsIS5HXhmbgMOac/lFqHxxn1pT4hdW
0GKyi2tSc9/ZgzUmVDkW1MRAnAiTS9rmWGzyBjSLuVCFMlZvfs8BcIxZxfkodvRT
tOtWDBIvvZORaqypy3ed6kChbMB7+wKUL5zmQrgy2xsS+3IsSTEBfbEZTnaXCSF+
nAhCSOagtr04BgbSEUjaMv2kPzVmkdjUDkBydlWR0A7vmqXS6aEpqCRJbsXO10yr
Fff6wseD3XJg6BfwQ2NpsXaXifA6WZ8OFuUJG6bjxo0gID9jCgSi14gz/Db4Mz9/
9eirAeV5jVDMbvvY/kZcL2Nt4p/68DaxV6gnHbC2RK4=
`protect END_PROTECTED
