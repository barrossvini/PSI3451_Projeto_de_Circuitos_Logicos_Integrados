`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZWrl4T5pCK8gM+LWgrRuXB9SuR6dNYM4WmNWAkJ0h6VroTyYmDDVfWIcV4Y7ybyh
aHnhratRhkJUxDrp+eZCGDQUbXxVuHG+ngVbx079zmSCvHhndbDhZI7Ac1jkZnm3
aEB8Gvh2z2zXvx9/OaUv9UpcVavCtYkBm+IRNImP3EtQx2ye5fh0XyleaueJuqEN
FUY85+yCUg6pyplNntLdVBZ0q1f1uM2xSs+l9cs2m89mNnUof2lKyxaDsEEOzJxb
CpxwntrRlzYvJLgB0xooIpDtsUa+3EEQThQKuaTQGxT+KqVHY27OOQBWYP1ohW/O
8I2vl8r61273Z9gf3s4hVJrgsXbqjrPWS4tlomaIdteQeZxGNWthpEr9V6g5eimP
VrhlAjarj3g+b1NVa+v40TJknZ9eCrpAo3g7X8bnd42aMCXh3JWT1WKDMz1FJOVF
SPn5wby7PbBbx1C3EZYnL/v9XAa/yzJ9gMOKUJygI/Q=
`protect END_PROTECTED
