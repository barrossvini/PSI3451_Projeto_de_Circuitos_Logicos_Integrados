`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/DhS9rcVt7g97DWIOWkEjkcXFDiPz7dNtit8lJPhN4lEnMcoRDXlMwMH2DDRXUbK
kv/uNJzTd/js53supUbacbCrfOmtNcMBvHov/9ZYfxy6B37hs9PEq5AuoJad9r1f
i2mkuQP7Uge5gEnU6GSTStyyjlKsCViyM/yu+BmQBn6hFnQyJ/Y7YMZgsRZyH+Et
VdovSJ1TmMc6B+71bHmYjsBplRAXCG6UHLN2hNyYKab2UGB5EoD4ddW+sniZzzYG
vPH+siQFDY5v4grbuWgIUDp8iPwzVvmsXeefZZiTgjMJeTqBHTdbk40niQxrypbe
NFHtyc1tVcObeIt63gcsI4V4tDEqVTSRt4GobNqtTKiRBsuVFJGsAhD7781ebq3G
FybeVqTF/1ot9syL7RBwULDBzDyuAJRxFFhtyiZdYe3SAmprfeUnGT5F596lsRBG
VesxmUqqpsIK7rQC7mi5ATaQeWQnbfkRtH9Bz2HiqjFfj4z9FgK+sYb2YZvqQfMO
c/I5WvfNh03jINEyyPaIYXDpjq/LImUmhYBvuZ3alpEr4qdk7P8LTq0nZFKTIOUi
Ua3WkpWxPGTIbTwS5rrybzX+KSDhB7e9RtEdSsRyJg87cNEdmj6ScahLmKOY2UPj
oZgPjFWxPy7trx3ErMoe3b96+ejaERzWM35fV3UAZbc1sYvngveVOlKR8wJqxB4u
wOL1v1i4k9PkxkjUMbXX29jIGIL0/eb4EKUgDMJoDxZ7Mnb4t0PcHtpw/IH5usu+
xO1nH75oqYRlSZWVdziEd9wVNBzqFF+YH/nzYW+bzb/lIWXgwXJQhCugJucRTjDo
i8U55Qjt5wMAEqSBomemX8pYYZ/ye2UO86vmBH+N2kAndZ7xtroMxUPMvgv5rcOo
RGyESgFyvOlIKih9MRA8OWb7f0dGNR3Ki5mV6ek4WKM0LmRpafNsBmbqSYy/5yOY
mwdmHgVHBhJ9YVfcFLyDAIEGXnMpgoVMnbGUQxi7XFEOGrdRqruOxPHg3xjIixBk
bEg62UqQQtTvv9zccwDHD3eP+ukPbmzOUJwmpBIMj2T281LHRZxhZHYtLkDE3gA/
QF7LKXorawa0ZAbYIXuepFwFnLjMOsAp+34ZPxKV64s0z2f4s+n7S4GJE3B6VAp+
TsaNNxIFHfERqfcKzf4h7jP6iUag0x0tOiFaDyOQsIU1HZZUYXPLZdoBOcEKPAwX
FpBljw5HIXl3UMH8uY6jJkDpImGkaB7l//pimnUMyvjOw3YvQCgOXFhyUYf8T3Dp
0aA0BZGiMENFlqXMtE88PYjhQ3PPE0KgsE4G+8uW7ravWN0im6OKwuGMr60hD+OU
21eKgKJvnFzy3lSBCNqml5SqoBW/QIU19shz+pkb/3SHPUOpdK5JBh7pq60JjDMW
nofm/Y0qudZlgisAqSzjqs3ZfAze/I89+SSjyVFGDr7Ojp1Dp0KuPYnQMR/y2BFi
K0nfKCiU/0AXFJtR/qLhAra0g54XnI+xiJyRtITuzpJDhWhNVFblcLMeuHUfJD1N
HJjB/w7cLsHW0c3lW5EMKAts2WDoidIv/dt8qg5+UdfTJkIHk/UVCgV0PO9LzVRs
oTcLjX1wEfKV/jz9a9cNlOvEzuDH4eLWYV5yjvEAD2AZ2UgRd2vLr+DsnZRmZkes
HOhlWHAChXQXtZE2qjo0JxqvR1f7TT1e0zKSNqvkzHBDzoqudj7Wud81ffLuUcI+
8J7alwi3EHgFM4G8gD8wMQEdjbioDkbR5cLSPYUo7NnCnpIjEfXKU3v4s+5zpcoT
9fgdsEgM8aKw9G/4YvH7N7XF78DqVwXkc21B3QWNMCcBPSE4ji29DID0jXGOJnwO
tXq2ElPuuSZSf6EjLQnprp/ZFYHBL9oFdp2+L1hUIfAMYiiGsYZXC4LqjzE90kNh
u2X2bR7XHb4GAA5N/d3+PTeWJBnm3bZeNw4291nch98OFZV2tjJoek2QHcMh7Y4n
8GI1av+Z4O4ukrDz145j9cL7i8isuiHET3y1ZxtRV/YVfk7g6crtVPvbwc4bSeFs
OpRMmPoDRg7UAjI4KGWlQB86bK90tn+r7G+QD2Ef6rYINIgcoDBsTsrF178851OZ
hsndHMH0M++bCPlzqYs+mj1c8sRqNbgZLEbPCDoQ7zgsTS/QbiGsAD/jt41oGBeA
QiaQojFYSzLcecHpHUn7vZp4I6xG5ldntqa1oOUYsVoOZZ+ZxeyRCYeTnEgDc33G
rCUora0QfnMaFFvpQPZaHclxnxIaRd+b5MJBtEgTI7l3Of2KJlOGHNoX7wtRWG7O
cBmXGriffhdLpPqnduRqfGolANywWT2Qm0f9laSt5a4jKfdNAduXlhxz4xSPAIRg
EsKIDeCbJKIWFthP2lGDLN9AeQHsI8kgKJ2N+drDdU1YvyzP0thF6LbdgsRA+/pV
/K5DpkskaUuGUe63cnFKmICMDNMj1Ke9AYR8HXVxGMUPng/YkQn1CZjt6bRnvgB/
rmRXXsT7dyUU4k7TDu9W/87ZrZ9ncYNLg4ZZ58Zg/FG4Q9ojuSyXUpPUul/044Ag
eW5eeaZTv5ZJ+6q4PIe2z7dCSXC1aGnAFkP5LrrFIgNAHA3srPp6vSelU200fKEH
iQFoJ3Xfbp2ZoFgWFvNFy7o6d+PyGz3KPONxftIsE+Hnymhypq1yt1QwDhBWxLRB
TWAYSHSyFUqhLedWzFbgmpuj3NnOTNwNLhZVh9XSUpl2GPvSEnKgohG0nXQiS/eY
6j7CKZRqXA6WnzqUaf7rNd2kSGDDV8GMYMHEPDwO8fY8TWc+nK9XUwT9e0S8IZ+B
BN7Bh2A5AF5YH2zHdVsW0156Ipekr3XZv0k94WjPzzhHjFJCGIpCUfzSlTxQSGTx
LvaLB5sHggDjBp95GSuexokLVNAk+z+c72YRcdBYDyVgFcR/JO6pw7zT7RoPRx3u
7dhf9p8qL9pekapypoaFxV+A3vJjqj92dl+8IZZn6u513GHxYGhRpuPEtmGURBj3
mU7i0Af6qrsz+BtV1Oq5Begiyi75w5ZqMdUpwttD238ZDFTwZ5V2UU6cTNW0wide
EWSHBFSphgznKPutxHzSBhRDz8xZKhDIgXR/ypKFD52fTTdvMQFx6f/S2Ls3qAZP
bI3CDiddeaBnbF7DA8NQUDX5AH9GJwqSV5evEzpysaTJmnIau1LVaOZQjM8teDZ0
784TfEYRBg/iIqlpwo7kHKeGCfYnLg81g+be0xsmJmp85oLOHzBWhezgQ8DKKZCP
WRvcKI6ig0j6k4P84L9C1WvQrUyiHFsvOaZer/ZvHhMOjB7H7hKw31IMYypB/qJb
888AIQ5lOTVhRY5BzfVFQSE+3WRWrnft9scmDfnxlnTxqqr/7kxGg0cz9g6BBooj
aG6xlpeX9wBQvF9f04/Yt+vdF7gyLNL9NeHLlE73zZ58vr4CLYZAgAjJ7YspMp/U
6vCFWUIzlblJQgBbkI134SddDYqYZQO8ouhuLihMuElmEazuzH+YBkK7DGwCMIaW
uuVmggL+FiIjgmQWkClDBhNEn1iAQwqwJdNHPDZAYsZRJgdg/fRVB7O8hpJYJzkV
Pmeh46FNH0M9IFkpnJ96FMdYFQVNfJ6CJOkiFxdORF8Nht0pvelO8Caun+gax2Ox
6FkEVjjc98bSo8QHwnFhHy6WgHW0vXhD7+izJv1QDV4T3UZaaKGwZFcXZ6m0ZatA
Rg0NYPHKWsT0T339Nk577bRw5Y1Q/S+e74sDf/hWWqsoyFjuzE21/V6ge/ZpaN04
sZsVmTzR5+9bPbC1cBWUA7S+nrncONu+QqB3MkecfvH5R/FAE8HApNGKeVSa5ot6
KbyuBwq+iuCYguuzQCm09l3+v7mAMAb25U/VluImaE0p/6dzhtx2TRVQblkdSIh9
t7p5cY3AQpbDG/zKoGJXI0raAmAmdwBMFY8tm3TE6c4i24T0VbhoB9fGpNyy9GfY
kgHTEZVm/e1zLUn6rsi1dZxW2pG8Wn8Xjr19Jkzb+llrq/Pp4Rs7XS2OrJCzaQTV
8+Gox7Ggo7DojGCdwWBTH75UzlGoOwmo4vDpNtug2QInovwbO5UntF39hnlVPguj
Vi7NbqL6gutartlIXpiL77Ls1EWQXAi0NL18xTZDTULVfScIRQOGgxrGQLKlLelP
boqZrP5qPoBcN5mTMtQiDNCr9GDdoHGuVwoEJNz491Zd6Z2+OBzH0hI27/Evm5bX
ZyqPOOlUJ+3TCO2oNFuEKEEPWLE/rI14xc0a77dfeFZk0N9HjOeP4VNNuNNKSgcL
sig9pottgIKAjZaO8sKM7Ga+y7LBXeK6PVNQ3EW6J5EXH3JPO0f4ttp8auXPX2ep
t792iIkhTwf+CuthXE1U/9xkeclVDJYTnoPNjqR76ytKt1yOeU2ucDg3K2EM6xhx
wiUK10uWTV9Owz3L9Gs0Qwrys6TObGs+5u9VA8ZMVGbBBm0qHB6VeRvJNt6ITWqP
vML4OrBrNS7BCpCKz4IILMBBALN6a1Q/Zd95p4zA5VNB/JteFBc8IhBTQEddmDuw
MFOqEWepDOiwHTCcjUiEbWydpBFAxaZYWEZjn/+ppj/CF8z9e9q6ckxOIFRIwzVx
`protect END_PROTECTED
