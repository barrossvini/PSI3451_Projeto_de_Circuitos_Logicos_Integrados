`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tV+9X0la4tl47mvGw8bnIQRvUnOW+UW6P9krCgtury0DIoUECqBfkzg7engyxr1a
gWxq0m2XZGoZ+EjtA9LEXpAkSXxOoWgvbvMOiyTJUzG00LIF/39+OGBxfK+4z6nZ
a8Rw5FmK3Y9M3taucEkJG6gTkgnq2M/vDwtSPcKQ895fOVXRw+HSzwzkMvc4LL8Z
KFEoLHETNpMWH+vLvt/fABTFNA/8OSEPc6nx0fwNhs5YUfYRX8R2cD/k90doZ4NT
WNjLLtrMSjQWqwQ4Eki3DdVpY9ski+xH24TXa7zWh62elMuwmWhFyyX4FQ33MJqK
G4G30X5/S6hpV8S2LsTZIE7mVLnhe5G24iSf8o3z9tVp15BjYB0BQxbm7e0p9mmP
VVAmjlU5P3uHpuCZ8yFxmk+KBFDZAxNzDyloZ6Ey4Mw=
`protect END_PROTECTED
