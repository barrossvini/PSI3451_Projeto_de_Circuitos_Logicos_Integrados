`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bEJ1tKPoa+DwOhx/2ZgysM5fxc+EnWkn82RFJ4WbD+8qBpmc3GauzZi3YUuso7yQ
WnKhXlSrB68f32sr4A15crCFvGgVlRslu7/um76IKxFj963meSwLhNHw0PH3iFel
uxcEka/aD9b2DaQBHMprwtSlSNl8tQA7Mrq5NnC6hgeVs41oyQ4UxFaQ2gNjOP3P
I1AuW2yC3I88LsC5aLu13YGwVfg0Iy+ji6/mFIpZYLwblJKk7ohuzgac0U17q9FT
rDgmdmf2sLnMd56w5Zv0DJ6oUTGduFY3ZXFUSKht+TH62u4cuQ0lzT9CIp/pb/0s
+UUoljlgNgeHp3WvWbBInihDGeRi9HKGZE8TUeE4DMLSf4/wFkioitEL03OgxB7u
NFm4tCHxRA3sXUTffUS/tmGv+zLjzrbINOmHHh7BO6j8P8J6/JhwryG8bBV4mQjz
voqWFWg6dVT3aClTUTUFYY4x/HGzgsnDVyYM5n7W8cZDNRdj7G9tMPT3OjibrQeq
P1YehCgFPTuGJxRbLEppCSz+lnrktAhkgXneOmsDvOEyLvkeYhpZbmI80jo5tqN9
xVD6rgONnrCw+MDp/7KUhUhml7HLt2lyjgNEiWSUEaISUirWHoqSS/Z2TRQSnZ9A
QDHtsoMo1/fbY3ZwKvpvY5T3udez2QcctAwImX8uwgxtGwm4Wi6WIKPLhUd48yJi
zKFMweMXXTD7EdUcIbh82Pce0sHMztsiag3picS7kzN3CwvV6aI271Ff+f1VrbJ9
BXMwSH/I35r4iu5XjVkj9He5WsFDKocnmm29edglIIKMqmKYgDmg+qQMaGMAq9bW
HrIvVKk55j82e3+bEl5wABatLMx7s2QpUzdtYZ8n0i1tSYBjK4Cu0JvGoy+s1Go5
AAjgoUGI76a4EmYAzyoGu87dwW5fB132EL22w5ZvcoUNO6gPjzrpj3NYw61lkLPT
fc7m/mD9R4lU4GwtTVviPG8VdJMoq2unAthQPeb5a463Ek22UZ+8eqxcc+RzGt5e
k4whqO/YjxOVGDGTu80dmFwYabo+vScUUp8W9vjoiZdGSMYgNYpp9nkrtXNcPNeC
pfxbHGCGju+qZLhni8ryUGX4ZviB1VfTtfpdN7UsLf8UXXDTbKMXX1XJQVENVbOk
W6kO54MPeDAcS+QEP/LqZ1dQrJatDd1qe1ytwvAY01SjX+TfIgPpXl7/M8ygionn
ySzFuhuRHNvx0NGWGaVNcauIJMsNruYML1jSKKXt/UvQvugT8ViwzyCyOGp66Wfg
d3Uxmwua3WJcER/zKuaqUSc3lelVmepaobL9G10Ai1vFuv7dDeQmAr6ArD4VfD+K
iBcCeACRHDhsjKQF2ZC579mvuz+EsLklv1LXB2rIVW9k9cYocn46+bVvNx0Q9XFG
sZpT7XGf7Z0QzacXMEac2STZhbYAmD5pFimDG4EuZ6t5X7ireQh6ZS8LUibfQayJ
G7rr/whetuzb3c28e1nJD61qxXkwr2If1l8Wb1RjkTqKgn222yiVlH+dqCUBvBEa
WlQTf0sO87YQmOrVWb8trzFIdQS8uNoa4dQMkl4UcqgLwOtJkWGIY1UqW02KZU4d
UKIWETr2djpyiHj6UH1mTHdGnauXsZfdbpz6aa4uR/pftcPvB98A7DXdeW3C13nK
aOQ9peiiEtiZ+30iYBp5PQthwYvg+ztCY9g4bDcqlUOJEJTK/2Ud87MzoQ2bDAS3
oQbBWbTx9YayuHRDTjme8WDWGUBz1w87m4Dwn8Ked2fog92zMQ8Wz6WKudYV4wGR
fAG8dkZB5sAgCNJRhs2IkuH+9TR1ksASwjjRuXVpqmwrtA3JrN/KB/DmuiE7XeQD
xH3yimmIE7vEIH4w4mz8Zuvxl+LON8L3Q/gt1PQSYV9JD3c5IBF9zXWQo584Lut/
itYmL/WNnbL8wvESMLabcWG2TcsaEfwPZMW43OrnSlzjowmM995NOK5qbUdq+DR3
vGWfvuNzhRZwq+lci9IT4hJaCW+ilTb+1CfrJjF2hXJjvk8LeB0FICmqHrR8WDCz
VVydlPdALuLmwoQIoVJA7/uOqL5UCwKceFumLYvMm6qWOO33VDtviIUe/whF18ye
RuD1ziNI755k1Di+SJE9oc+q9RHr/EEISzNR30SAG1fy+NssBudN9yxdMt1Ef1Oy
meMvyVNlCifXAF3MnGgLlJw85u43DaNGfThG2gUJZWqvNrtd6kkaLMg2k31PMSPc
O9eumJV5JCdpF0D/BAZw5FxmdGLLANTam48VtRATl3cxMMOKl3uawLn95fdNODGm
yUdJs5ROmA+62cZv8eKGuG8QosU0dY4TxFhR4wtQpqrl6WZMuTak2YctrQn6ogGI
39JkdHkIqX9sytiGzYdDSz7rvSzRUhrhMKT8/cQmi9QUX7jPKWtuI2gxPQeEECbz
T1eS+99FUYmVxhbSDrtplNylD6BLWGe3+vL7WGyCF+eMJeao1KTSIYjrsCeA7fmT
sQ/BGwBAAVCKz1wctZTd7kn+Yi9qRqY5s2qUY/DksTSQoh6LLV0+zSmIgnoM+oE0
Qq8t4UcesKJgktIiNuSmDFZGPn1RboqTILmQul9Vb3VQp0fHy1c8OZ6zzYPrmrZO
pRDKPwdtWu048ONisT00M8XEneia2OJMmG6RGGDu8udBhXxSZGZlIE/DOjacGJjb
MFRcG5gIWfCzXZjBFW5x8T/rzqzjcuxewu6Y8KY7L+n4Qvn7obOuJ8T7hLi8q4jm
xmxgE/5onrTWGua2bxtW2WzjEFjKPT7uCDv9+E0zRbDmZSF8zXpqhJiaxh/YDKdp
umKEKVB9en6gBfC3/GB7SE11WHnK0GaHiGjg/VeY9mvEGu7+h2EcxM/euiF3T8yD
sXlKjtqJEBEhZSO8HJYrM8CRx6N4Jubk8V0q2MzgdI+QqgU4IAllR2ouWJ6Smpvi
kaxmXVU56Evx7AI5WiJxO901ED1XjO02GWX94N87W+Qo53aWZRwLFXfDfOOckzfW
VBx7b6F//igUKy/bTf3oZJJb6prrCUtWe8+SbS0TFWZ1gcmyrTZIDh5vUMBL9mjL
IeZfl2cF12Dr8aeN4ZJ4ChD7D2G4xGfBsQOP49kZJ111HZ2CP8O9q8a3ZMrGV/ub
Fe3oIfG2izFzwUiHOUeR8MYZrjHtNFKFevIfclekuO70cFRBElUoF9m8fCzjbKTy
0A5IL3e4eK5oT3rfgp1xkMFSsaraeyM2XoWinyG6G/9XVGFG9ySzLTtgmIg/ZgOf
Fy8xdZmXgL4Zx2q00ge3BC6r4Ir1aI9EIWglp3rCWsWW9sGzZXStBxVnUAyiMewu
wDfpIW3rg1cRFaBq3gsHeLqMLGkXwoZkKm99ofrJgv1GjZjOI3SQhw7bAvW3/4AN
/AIm+rA7pxo6tAgMP5PU7DidQeEFEsJlOl8RaqpJGjt27xVZROd5KnGPBStIjRYJ
/L5Yy5qoOLtUkcsvHqPvteeU1wdx/nYNroAzJhJ1ZNJHg50+CRa3V8nRIj1oLok6
DhbHc+Nz8aRhdpJLUJO1WI6U3Qg2TrJ6S0qpjvvXPh1mIwwG5qGaZb49Dj5KXpNn
AydR3zOFgX3gnzva7QkOV4Wuk29zv1seGmjs2AhNLVQVl8aR9jvwNQsVOu1fl0Ok
KqBp7dmLpXhozcy23+z3JxQQ0/C4WYixEnKPZJBWbCQBFhuucxZVuYQxv3LyO65r
a1pi84ouIrc10oX1ic2PWG+IIZZkZxRQjXw9uQA9YWjmnjdQ9KkemlfsBESew1a3
c+v+ViLc4ivilQkQ5INSSMw3yq2snZ/9mlOiFQobJktiu8VIdKJx/8aliHBOhXU1
99WLF1pp1Oqgv4JgfRPIGIzd2ubow4wBtO5c9XZWUGMhbKEqRO3p/0Lkn6tnKhg1
HyeKKDsS+g6QrHSIK0MYF4H2+SBBsrfB6g5VjT6QXz4gqNmH7lauD2mMrgNa/lfx
kvTqWEI8PNcBA3x2KMQSE78fEnY3ZJ8c+iKdR/00qvKnzrqDp0YzkEfXHnJqHlWe
FaLwDMqV9FcWEMZPp/J6KLOJD6MG2OdSR+5hOMHjD8yfrGzjYJZsXW7XW1JPGjD0
h086snUp+XcpOxG4Ou5sPj9Is+Bxe2W0eTHXaAi08Fk8/l/y/sy74amPlcDOQbxr
IbPha5or4hV/vWFPpKS0IpsdzHIBUaAkZBVAYMxoJC9vaSE9pmLRrgaOjBWs+TaM
8JtEv1fCao1fTCw6vhp8SSgiqHJii329wBonFrx9yTXdGH2cBhWzoxbBLpK+DO/l
G2JzZD3v9K2/MT4flNRHw2Idir8O9kAQHMeNydAtHoDqVd64+RvmuYPegRQWr7z2
F89IBXmFmwgXbgsOnInVp5JVE8E03cdvDNq9C2U0jSEm0JnVU+QQWuOwUVQvXdkD
LmiNBxjWDNs/6FVBUaDXd3fFytSKeVA1e6Km3+T2J98EfsDYZSGJRGBUU7vyt7V7
vl21KWdEt8xxH7aYNAnosp7ip6/SCd1d78UoaDOnf0WYK932xb30DNSSWmqYwn4j
WGF7SCNzLXyoS4zGhkvJ8xznog/yrql+ApttRpv/U1a6d0LHng1idVk2ppAyfi/J
72qmFziBCHp61AwiHrBi7qqo0kRPRTwB+3sP+Ln+TL7R4ACj0I9Kt8s7+UQJtqHe
Zd7UjU5kMsA2CBjDk9WXp79XYig2HlA2pl4L12oz4JofxOsuzfle5c5aAHfD6qlJ
sTZG0xs8sVD9efRYKpE9GNE50NZ3l7lJsMqKb7xhS/7gVabNA6bhcZjRDZpdWcbN
Xe/4G7+rODGxfhLpVG/ALJ2jO9tIdKRBkFLPeoNZ+BYNb0uFz90Y/xWf4aIIjuB5
8g2SqZX2QBLTlicVHgUn/hl0a+V0YoVqUZ66AyvtbeePYSbqS1DnZcanJnX+6ai4
peoAnofL92LH2eb4T9RBdHJPLEO1WV4XyDhfj0jG6C4sqvnH9jlkUHeoU/MgJ9EY
fd+fBgpwK7w+nsujiPUGS6c37Q2K4BMZxZ0ZiCFYgU2R497GgK4svUi9BbU3FyaH
Su57V5zun9jzl3pu/EyACSAeWFTwO0jFJGLzX9px5v5/BR8U2eB7teObfh8F+lZ2
/OR2mJZ01Nto/+HWdn9Xe4vV91qnsDKEfQMTrY7a0OQ+ZK7stg+xJYjqmlCzlOLz
8s6UuHAJ/52AHm3rcFHnM7nkXLJ4HZT/nnMy4BIxroRjR0zQxudterw+9fsWZyW7
axdvQaIxIv4biKOVavbE9Q==
`protect END_PROTECTED
