`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K54/CZ58WpVaZAXHyZSKE1GJHiz8iasqCx4iqjOklYUxn6Frzx7a3r5MhCJJufkg
a9zGgen7ZBHm/+pTyKszNi8tOJ5Q6/bO6xSZDbD3nALE8Rce8VvUSd7LITOT02vo
FEudqEenHaPfiZI7RnAk8Vfy89wSrGjgCbGAjlDAa0bi/7XeQwoNKoVwBaKxRZGS
rtaTtB2LiRSGPhiI8GQSC7W+xTuftXuX5WXkXnWm+st3BWmlw7iyJQDyZ+4FU4Ew
FSK9m1bGO1F9ySLuOm06Dr3kENhoJxt9HDPyYeMxo77v/knKlcDfuBf5Ov4dGOVj
mdTxh1OrdX8C/KgZSvyURlbPveWa+BVLkQ7L6a7wJ0JQJurgXon4pMj7KEuhTVv6
iNkmm1wsYfZE9P7VIQG7ph2eLb7poI7QniZ51qyxlQ+dhCEcy9kcTZEj+FVmIYUL
P+D1nElwjC6MJUy2wNWTJYq/IxE5ClFBuveQOYGcMr0JEoK0bdIkpQaY74imnI34
+wheZFnjsc8vN/M6L1tLfRzQiXwQI1vnn8nAGtu0Zz3KrdfCvnnNCcWx+s1lMAkt
HFeWmdzXh/eWfUd93skXgfvxP/HDlQpATkXWXGpPkvjrClp7/MO29JHyYdPbchtH
JuxAD3JBoQjGPDHW6wxjcyK8yCfr4VhpDWPPtbMKNhZOjAu+miJMTcEyRGzIGe+7
DeTajqOJIyRlJFU8HxxFZO5TQJV6Hml2s4WRp1VsEQev8LLGrTPCt4bBTXRy1C1T
7+4YeB/boG1ezNq9jOyuah/lwvqXnAvJZu2SCZxnJlphm34LkxrLpwke+pns1NQ4
YDclFPDSzPom7LsZ8EoYBd4h5G2YRcj5yJUiUwPXM/2lr+EbcwYnlza4UlXRaWkP
VMOFPBo9WwCYiINpAkSV/IO2ia8IbM1LSXj5FU8NojF9osS4x2E9oPHhL6cmtChy
qtkIBGbjA6Z1rUw0HcjWipM4tfLJY7ZQoGZlC/kxsbto8D4rAIQyEN+NAZLLVHgb
BeRIaZjhXrFZMpW5+oFuDmquCvSsWsB0cVexKuMhypKQ11UnWfuVJXxVDlnnqk1M
TiM0ZGZsrid2E9sTrFlFdyrQCGpwjyfH5W2Cady+7EX3kX05uMux+qVLz8Plqb2z
jFv3sD9uNDxIFR7XWRCbhmemrK3bY0yjaUhKkoSyJETWXzNiJBdkqknDgzuhtoWh
lUZSCxGPLQASJMiBong52wOXWlNjofO8MCa3/ePA/HYU1dgDcCUR6IIB3tN3Y63h
rihw+vSeSPM6BtB8awLBSy9SgfiZFD3TpyDn7b1qkq9WWJMuHHBLnFA2cgHTppU2
2Fi279i14JX3AAo+Xa94gbe6XyW7ccV12FuTu4GauLStH7EKPlW15g5puoRzghc2
v1t/Jt/lOFh+7JSe+5nh/WQJn1ED54LdoaBCmKcZAY8KC9YWbIHdzRnNgvrBp859
ZmyrG+z6B3kyraB4JJaW2ulpOiOilqptMU8hEx+01p41qFY++v/7XKJ64YW0vAyc
kiQAegXR2Sa6kyDDbQpdtTaKVTp0XP1xefAgkisZfBDfODLtxag78NAbnRW8XY5e
9Noz8Ru0ZuyeeRNej724fHOtky+W3cz7cWpFST3P7X6nsnnhGPeVNpOu75O+tmsP
+UIYQitNJmD+BoMwOyuFng==
`protect END_PROTECTED
