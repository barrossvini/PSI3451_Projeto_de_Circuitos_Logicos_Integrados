`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SHIuv8JRlv/wj+bJYytGXU/KSR8gGxAoVM9/SfsREBuZx6ZGqR6kEjC6MlKcusyY
UhWly4pmsPZyIouZU8JaLH8wztejKon1PDY591UO71r7JgTx5H9JqVIcIsuVFH10
TNsshYw35l7s9N6A3sI6D2uZSlWNb40OzDcjwu1gcbXALK+0ArPELlmHvh3e6onq
BkpZpe9ftljAuY4dJEId3sC/LjXgHp3o4sj73G6qnfR9SH2s35TvxFuoClE1VuRy
2QM4TpwELslXGRwFBOpPqX7/ZRnJtMG8h4XBH3OtL1MOtm9w4vhtlwUUo3B5yqyd
SXQhzt+H5LwYVzh13OIohS7sQTsTfjzosWYmxq5y0FERY7HE4xFJuIqxz3gphsff
jIdospBtCYZX2rJVFYHVL1fyXWM072diD89yavnAuu88P0nUOj3+gK3CMrle/EJo
C52QBZY44VNlxP7ClclEdrzb7mKq3C7GQ+iPGKHxAA2f0couLWSLCgHxFHMzJ2L+
ehDERD5QP2T67Hed7Hi+vWo5rKEh6/5y3rapUmFzhKVF8G4P7gXN7uLyqZ/3CyZg
lue3ogOMXbiJBjK9DYzpg4DylnMhOgYLz/NDheEHwQ+N4Ew+6sVlviIYauXJZilb
1pETYIB9AMnl1Eo0edokL7N3sneWaUETo4e5a5eArto/mfWVNA35GYBly9oA3m+B
NRbR0i+D8AelvED1WnucUZN/WqnCA6QHCT/xrs0RkD+ESXkM6w9t0eWTY/Yp1xlq
32NQIqA1iWUGZj3lkz4ALGmsIG3fi+Tpf9fInW/mgZHDPWO3RDAjLLgs/mJxViqU
H5O0m0dpHFoKL80letBUO0MXO6hMcPI5Jfr/eOlSWvgnwJC3tpQdD4SQfw6QJ88l
onybqs/Lmem8EH01SLWmFIUUb8OTVhEw3ZF5muxdQ3qUG5Q7iCpCYMweWm6U5kak
5iqbXIybzz0xgp38E/wbpSgd7I9kSLCsVxUoFN2Nr9Mmq1XSbESnx+Oo6Fax+6Ml
iDFHWWMOvfvJywOmAN4yQzplwPzM8rTNLu7TTWxlfCkOVe2vpomboBdr7CGXxg7V
aHRt07OM1zQ8278O2b3ObsxdTd1c62A2tMxf5g38KMxcLoHwxQV1Mc9ubgDzbsMS
0SS3gNN2Ypurho0wcm79jsC/iEzdoB6T+hnNkIGH6X+wSTuzKtJZJMAxRyFNHrDO
ncKIl/0qhfAZFQiPBLd59Xnqjw2gZEjEShvdkPKOU6Y=
`protect END_PROTECTED
