`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BOJuTLTE4u3a8fZfRjfRK3eABbVpqcVWZ16WrsvfnrQmAQDLnqn10yoMDebeTJ6H
keVYQTAhwe4jUqatNbJAjBo5qnX9uiEnxaUEd5VlyPar3eUwYNnPfIfK9TT69zsB
ML0gkIQO6wtY94X8ljfIh2AYubqlgS6xZ24UtUz/zREzy1kYYKNC3n1jJkCDNnp6
l6jvk4GV8oSKNFP/j/DUraEXGcJE/Sez5ULcIX/PnYa6oqmsMW4iLGx0vUdyrC8Y
5ZQgFsmla3rMYHQm1tdiMZXLhaXZRYw7EwB9SatVSe5zqhjcusSAJX+ghHDfHFzg
8IPZQZT5ZZRYGDcs/JtnxpcXIO/8FhbYxkJWx7m5SXvpXKZIpQm2djb4gY5x4Ain
pDesSS5duV0kbWJZt5q0y3HfglNxZ3soN5Ttc1WIW/tWnQ70b5ErBHBbA9/xq7dn
RaDE+b/4o1xd3kGab2fRG50bZYxaYeH/S6WKiD7akMP/o/L+WkuOata4n399fROJ
Pf/vnKHi9HNOOEyu2q6bzRpkFfazAgfwYee5/y5VZmlil+GWrFRt/xi3215AfR7A
vWdpnoWPqTsINBbe8sOTTDftuJl1IRC6JHFo32PTmldP3YY84DXcRABs9S0yaV5h
3pF0hqnSnCgiy3kHVwua3n85Qo4dBi620eyGwpX+AdLhfaxVkpBxPwX5nXttP8dx
MgZ92BYTfqoZ6ShY4/ZMEuIWrxZpTS/zkJsTDi6lSoXVvfNUmW8aJm0y0Ico48ME
N91inBmEmiEL18Ijujh0lNhJYXJ4JmhyiX++a1b7IlWREtQZoCA/ZUI6vC+7z65E
STt/lUej0zXDGPEk3F9V4XOdFPKBkdxVkGNAs292Rixi1vCtTUqfcvOX3UtlYiLh
eBUpNQG+gUPi9rcYyiZ02wJly3SVk0Ud+QhRfoD4cDP6Ja6ftrjk3ww1Y1xoC/aT
tUqvOSRBLVsYsuIB7soASi3eu1EOHQmXEF9lNw2Thd9W4EU9C1bZWaa06zxABzC+
uGwEWJvoSrI+NTqQWCNpwiqfuoIU1cEKeAioJftztvSwrMbdJiGmrcbb7SCoL1mW
Sr94UxRcc8huzol7k4THN837Sox+vWDAMnpT7K9HB6p8tZ9e35HUzFHt2XEhJ9ly
wjRxWYDCIQnBSw4sTXbZ2snFJ4dksd1jQ8Q4aSJ0fo7RJgyTtbz9ItWG09rII64o
bCL0pbMVsuUuPoSyODO2N9HXHk1C0j20KACf1WfhI/hvoC26FlVvcdpeh3NgoDKQ
N/Kg8Z+sPp8E0JBJlfVOHT8Q4u7FE5ToDHI7cs7GcE6VOTMIoPXZ3xet8z9xfXch
Kz7OfKsyGc85aMvacSAu072/Fic5uX7zEl1XzmU6Mu2mpfuZAdeGYEojNhxY9AVp
laJvYOhBFqy46jLHVtaE+GXXEIrMq+03KRtnbuke5qU=
`protect END_PROTECTED
