`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vM9Vb/doLncbnLkvSRTGGKESXkWq+oouaBjScKFWpkKs4KMh76KytiAuM8vtBW9A
/ZB9vdMCpcWgbsSl0GGGh/eglYG1AlhD3A7cb2fI/oPPQhuxBIFN2x0NB7yktGiD
kAiRPCOLC7m+bQYOkH1H5sLI26KDzv2tUt9H6rMrLwR9dE/NE9au4XQ+9XOG/XOe
YZwUViHExRiH7kR25DHKgapMMfmR1eNUIOP1ZLhVpR2MLKHXOrDBP0YRfXUgG+Di
tovlVtrStISEAwZNGWJ1cqQifvbVI13cOAr2MhSZEAiKy/bd87vz6sDbaE14EyPn
D+9n9B4al3dgEx/VE3rc3+1MGDROQpS083ViwR4xEwsDNEUPniO2V08TqMdYymWf
8s0ihDIBD7TbILSyEa8Ww4ywsaM84VFtmzCIvF+MvBeVzPVYFDEIwMM6EDFSXkmk
6ip4SU8NbibEVkT0B2J/ymx9u/ulGDfB2IaOfcAvy6PkVt5h5jeokDz9ZG7fskrS
RkDrlunaaVPqbOGAEMjWv3tAZznrpQLiTcgmv4UcHbYoI47PTI0acwAsK8YBhVrM
PzCZREz1pmz8w+/2EaYoMeo3Sj0GLkHhNCjtPxIK95rc7tzwDxOUjaykuoazgyCK
gqPBFbtxw1Gul8rdGBiulLtpwSE6JpA/9R66wPFPXYsrfKCu5aCgTjifEySU9+mn
wUK/odkjeKK+/c1h5GOPkhQBR8jHCLYfz1UlJaXjdK8cT/aNQFepcI3mLd4oKlL9
/OajlV+YjCC/bl2amkLdaq1Jy2uew0uN3CIYdBnHoVB5GmmsA/7Tosi8/q2IsHg4
EbnDHAXI71Nl/a9/Gbbbi8RVnpu1hipdelX5q46xGyU3fo3QKg4esP+7fEDIToTZ
PDz3OHCyyKlfokSPZrqR/OZfD1XRZSST6G5DjiDGYf0RLZSeqzotA7SxTfywyO92
B7Jc8LOifn5k1ThbldesvcTClY/gvOqKci4TK3+uBlAIq1ShxMDBaWp2MQHAItW+
onc6F0bcP1Nw2AU5omnIs+dTTv8N2d3rHKP3JQisMQ1whkK4Wxt75qum3TjlOlDU
KIunci844F7EmjeHxdTyW66chadcNWkF1FnXr0cb4SYHg7/VVleW/wofO5T2zSGt
/YxqyUcXA0L84Yc2YCE3BzfCJgqgYQmzslBEsYfN/qGT9qzi1+eEXHB87U+p3e7C
gSg5CNNj5lxBYMmyNTw0jVzsQwwagiyyl6hrQCwtxsLMRvrO2CSolCaN+Tf8BJRq
vM8ar7qX8/UFgWLpo3djuptqST46iQ7hMgRbRT52HqgOQID+Cf/vpX/Lp+Cw7nDU
lSuY+1ADW8iVGf3pgL1ZEZwtajeRKWIIpayZc6xvb3ruIOA60VzWELr0EdnDv7xu
AxRXn8ecKmiCBomx77Im5M5sNvEosbhOCaKBWfRGo00G2kNROZ2s7nfpsAZ/vYUf
4dLAbHQBlACO0L+v1knhMGbmpVSHz1VMztMDDVtyI9y3Fw518UloprEUcGMDbXPI
3+/rcytxH5kN6uvc/sEk4sL5VU4wUwLkYB7nUVSR+TyF/kBazy0fl0IZa7FYk1P9
BduIAtmeJzVM83Mk1YTHG7z0SAE/HiCQu2v+T9tspuU66wg1pzY3iMES592ILUdx
nuHGyEE8Fp0WQRqy0TCKpJ/hkaH+BFMMfVOi3a5UT3UmRHhcfVGwoin47IayT3Od
enNACOzS8oyL9CVxCyxhL7s2dEkHf0Gg2tOl1fYNj2e40GuNDJYNjs3YPUplIkwZ
g9bS8iYDWfkaBWOV8d7s0rGqxztI805q2gj0MrlgKZxybGc7z2FDFMid5TpUFPZB
dOJynjgkQNfm7GuFNG/8WNZAlywYycEanXIUNKoXFKRHJvkV2emJEtNqR3jbH3Wy
olqWl4cjAnYZeYuW0kNVd+QTULgxCvdX1oJJ11rTfla9yTV5Ksdhn2ZOHzutChWp
yUVmkV5v9TWM64ud+ea53uECYfhcred86uLk1dkH4yZRQBNpmH0YirDbfKma0rJR
03z3iaQlpMflPVIe9BqB/Ahz1HB9dyP10YV1S9xJZd8K5duG0siy47220dEARDeP
HzVAIsjvGdnpjWSxh0karaisU7ZQikUuwLPtgwAqF9n2je8oW3RDXMUR6CUUdnEd
D9NnPwX0rkBuLCqTfYG8KNluEcJwI22+00vv6hHRWDBCoxcwDVnPRqApP9nm1mzg
8y2An6bt/JgUUYb8KOR/3jZh68jPYA0CtHobcz5mG0Zdz+uWJDhqeJyfNnmMQ22S
32WrclIoyq5gRat0sl1tYfCY+kLrjfZ8aBclL8wpNiiQ/IOseYZ4FhL0Li+fVBsR
g2CujSb4Zp+V8Wxk7wwKaYHM9WsvM5qaSB08Kr7TPQaV8INIbmFHDsdTHsZ/NEkV
YjZlolnaKXZXvvy+RFrEQMGcqnXkbA57aFQQuHmPzXhITNS2J3ze90NLC2eThLVx
ihV3mu6UfYi4wF1DK/MiaONgyjpnA+vW6O1Xm3FHf/8wtNYgORJWO4ZkeBLShMyK
j5aUUc8K1f4DxHMxYDb1jH1feuixWgpHWBugFs3Jy+yKza6Mt3O5stXZ/vEH8bQH
WOpd9eSo0+2PFX19s2sfilR7qVv0br7GLwQAAYcBq42IcDhyFD9ckJAK6qdxXFqI
70PVefRyEVo9siMrFZNXiAMFmvWAIdpwfHoK8PEej/LRGMg3AjOhjrYooe3v021G
wpTDjlZpVwc8GNwheV5bDBur+YoFhO4+iXULmXOnkZsojghYAb5vaPueGXSNlrVM
SlWzXxzBb8Rqvf40/SF9aHmz0gyjSA/cY4kxtfMMVFnyM8JT24QPtqsnE4IsbXUk
vovmEbjPZDjRPxqXpTDO7iL8+EEvFAgjBHiZx2Fw72s7DQtOOWQnJInM0Iuqxe+6
TR3HVqP4WNqDTcLN6VgwJg5UVOXEqbuBq1gI125h9iEpyPQL9Hx1yzgzESjsuD1G
fxW/PZAFk1V9Z9ICY5G1M5SInB4BprhC8YbFdKTHr+ZtGzaHui7jE4IQExRqR/oE
BEFAtfDTpDTVS9C6vtWhgIZtCfTb7z+yZoVNz9WVg84I+nroLhEuGXAz7KP6vO/j
Tf8lhBnLbCLvyYJImIl5SMZE1OvLyx2livc4XEYq9LGKNDOQSEkwC5lzrTk89+g0
vFj3Hr888YMK3xPpJSqAeOT2T2f+iEu2Uwok0AbSqVe63wItF+2RhWJaG4Im/UW2
M3xB8RUpSrOyhfavjChFfyo+hXcWhGSL/O8sIJqabBM/Ha2BPPqenmNoUyNHOmUH
OJVMf9BXDQ9wLFRM++5rQCZwGxYS/3N/QQUxcnrqVTBBSQFvbtbWvSWhe4bNJHyC
KTUZqsEzHJccgwQDV9MFCRdW6dSct4VBK3/56NhdqolbHphMqNaZGtw0qz7Iv8cj
Cz9UmoobaDReH7v/aI77yUd4tNQ4betlBZ/WwLH7Ya+ByZ2ME3yJfevrUugFaHwc
IZYgJHVkL5/bxd5RrMObLg3hnvcY7O5JhFuiy60KHuGCR64p0BYznpu1lQt9DRgp
NwlHew8fiybfvso1Wwex8XC1YS0d003ygn51/8paUk8M9jaV4o3yFc0Nj2a4z3cP
hXgYuVT7qa2skZQP6DoUg7f0bSXLiHvnzoiMabTMr9k2IIoOz2hr3tSGaQNpOyjx
WiKBOb7oWdhSik3ii52jZwMdQTe5NnHVfMlCeX+W8s2HOFKpVjfT2PgZNYxki4yB
Y5LYnqwrcv2uv4TuPYdVv7F4FT4rxPRE2Fb0qiiTO0cLJOCr4QhjtyB6gcIt2sDc
yeAryizuS7HJR/49fbkUivvbEnchRHEy0wKBlprV5qyQfLufUzscWpVVVVlQZ3Fl
3PuMHfb7DhlerUWNACisXQWgQh106YwkOl7esxR9+9fza4YSt72uJrjoSdaU1Xy6
pSilebOpf1N9GBfuHu9KijM6EKWHtqovd6oPQ8sIUXSYIgegMB/2SDnaItjfdGAv
LG3gXt4oor8AK3fkZGcNfT6wUgjznNReAFBSUseEp1c4GcsV2547gi8ZmWZYZLZL
g9VAHl8IFrJFcnktOFhaLnuvU4fUU7TU+Vw3ndMd20bdduoNxyXaHx2GEtXFPUa8
5mPkiYP3udaErzms6wxtJXdNf4mwp3Yp6WyA4bwWcaz1lnJPMYLLaaYaKQIsZiMx
csnxV1wwYrKw5sI+b85DDA731kUqRQUE25ASxfrF2EhB4YNRUdcKi2vpJkEK2tlE
a1i2TckusUfD4h4uXtd6FRS4kIWS67LUEe9gfYypEg/O7hKlkFeyUlA2YhaSN4PD
iBUkO+h6AzM9FJIeDiHu7O96PYbTlHBtlDN0LC3DCh80ytBuFlFFqaXjFd+zZ68B
qwx1+mwLRQg3HzahBn8RRxyj2bpHyEz1lB4PRVAAjuZCqrX9wkyjs7/ipFNSEmQ5
/zyyKGvNJOoVOfxZyOClV8GB/niZK7hk+vAW6q71Rx+YUz/kRrkO+4T+tkQ3SXVx
KB8Ls7cH7TyPONeBfr5+DZNdA2meSeGLQKziH9KKa6dnmnXhRelFTQOgAMaHv0lY
0CyUv6u5m32roWSMJ1gJiuk3ENor2E+gLI4v7xKxJKFkpHBT+NRz+wvmhjyL1sgp
01tYaVuP7rTZczAGEWF6Qv7UQHsUhRNdhQ4IJAoyEDQ5fDCBlekwihiHAtNz9HfD
7hpG5eyEivbo5Y+wJAC4GlvsIMrYK1GtigmtCGgIqgDEfdToM4V7551hn6XO/EwY
EhRmZeDNjRC3f6MHciRehoxQYsOB3ns6Oks91PtVgRF3hNWly6BmU5aFkzDCJevu
ZbBeEhGPrTOyNiALh+3Jg3CjLRvYHXpCLu7RCfH7G15wM4vttuFchBJqGan2RjEc
kZ7uLIL2k2KXjRzyxlE5TkCGXP8kOacUi8bEBq0SH7dZnEis08xSnSh+qLgtv/Et
x7wzO4yQRwlw+R72sF2q1jlAupqm45DmndDWqpvx9eau25LMyfsnYMa38cVIx1AX
4taggGNm6LW7VH8d1Ulck1JiJC7kHLbYQZq7LnAPJe5FYlSh8hNujcvL47SNHdMF
5w6j+j9qP1oXJhfvWzWSgzfW6O6GyUh1XPqmZKFYVPzW/SkbRUGGzVnCi/8XOCnh
fQPCRjzxBTTtUwO4AyffY8YAcRm+zW9OB2gxbbGw4eNo9VH9pHbfDMCcaUBaC89/
NX8P4WUCerM04Al/URRd/miqjHtYoVyxTHiRPpDBEqSgpkzmU6fb3lPWv11AH6PI
axBNpvN8hphZn/H7VsMDwlQznw9X+FeIQNXEOdgX6e1OfMNMBxzX3BlYS11w0BxN
jwk46TOibThmGYXiAfqD/G7hQ60sRomtC3a1f+ksgfUK6Xbg3/5zT41lI6aorSwn
QM1lz5e/GxeGJLX5Y5BkTIpHXIZAa5xchJh45fWNNwpxCgEqiiRAXZ5ZbV24R/pN
9QRX3dG6H6zRJVsgls97OcIuao+9AfaueIpzewarATW3RvTxhkC3YR0tzU9tTcAa
jS7rbOrQueCAb5DuiRMoo9SPzrFEYvhT/CJ4l3IxGwSnUTlTcsPXti9vV1Mk7nkC
7SRWDcNOQZ3BrjIVODmDywBMh6CtLh7f+SDcL+B6hkBlvG/zaNOSCAaNTTk26psX
+uPwHEKzPpXhbgOf6aajz9YjV/gJ7Oti/DtKtCUo/Cdvh3H0lLGGgCTOTuyg3Qi8
+d5MLAS0r35vBeI1eAuSU7quUdXvzyS96LtDmRGxFijZXLCW/O/GzKNSZZTn6p69
eJ5l5tgOAZNeO6QZaEzVpJjpAC4e+ixlM2/Kbego7k50JriEjqmwMrl9DJ9q+HYk
QOl5zoVwZJRip373I22dHDh7rtIVI9DbJZ2ekYHL4qTzuzS6JBRwWXpQuNBtJvd6
uzU6DTWGEsprhqUUFZ+N4sOm5VKyCFNGlb39WX+6t7S39As7MM6V9E+K48iZAMsi
yQiXMdakJrBvja8SRuvu73/Sb3oC4BHA4h5DUNZFV6hoqnIVpoYk73vnB+ayMsFS
IZI2Bdny7kKVK1geZ8Vkgcf2SCOUxZnsTz5wCFokJiMI+iJChCp/WfWvmD7V5svX
01s104bue/kLXt/F9RT0CQA+MWY68jklTEMOKNHvarYQZPqLt3wxkteCdMmDKCSs
BQ2yV6q/sx9OFD8xf+bDpzvMaW+/iaFi3OTz9DIQL6Uo0JQgf6KEyIFrzgqnDPs4
krjFNfhZ4tnVbgbABqzen/PNUwQ5JJjN4khxZkOft5mkvj/ZF9mndMpPoklCxQ1E
kQAwBBFAkA+cV4cwRDP8NWzy6OfcXcKoHHEagvRElq7KE5a6SMAaVx0YmtrtuRab
bs8vG+g4h1e5x+QHdWDpA3rJdmuCeZmATpZxEi8n6aX7Oa4dQq0PTd5YMzzj/dhv
KzSfmipJrDFgdbmBgOoS/TjM+WVTzdzv9gyZxbeanwcK3u93eSMJXrXuF8zGqVuQ
X0vYMHRJ0OdwVubQkzuGZEBEGDfP0P2XzgsROM0f/AnBCqjf09wf1OtOReIRMIT2
deJ1kIRKhJ/JAILaoyCP+XDQ5k4Six9bSB390oytHRWt+rkBR1YvxKq3VF8KUlE/
ZDe6eUwcSz80LCKfxjmx8R3ck/KyDA2G2DvlQ0oytgglYnHXTg0Y1ob8R4e4iIeH
JoM14gUF/H7fYngYrUuRJqlOQtwCnHC6yErSHwBlr657kAxa8sb6dEtzMfm/ArbK
iH5PeiezA1h96s15W921BLAfvrHAgHBngReUsMAxh9rmbuPj9sqwRvxqobDqYD79
YfL70vo6e3akyT4y1IkpVPNQ9F3Yb6d+646GAQTilmfOXKGmlStF4K4ibs+bfUnz
VZ6fmyH7PQJLfRIVxJJuGLWd6dM667adwuEqYwt/SB9m9fCg+CkQ3LmyLV7NRUtl
h6AQhbm9010yi3bSoDHcoLr+6vB6Uo5m+RdizIbBc8x1favy6H1trkf39bYAT0J5
xaQmsyyW5wUDx3dNoXinzjOOnkiLwKIjQXe5YS1aHJcBhNI4FhIT+Ith9LpXGcg7
sMpYgeHf210Ta11gKkYh7G2OTcDoQI7Ovo8uGWKuUqHn9UKMHI/awtEMci7s7bc7
8tjQ56922J97kieQAaU+SVysbC6h5FJAqBVfjpPB4uRVMoyihYRk2IHAkyuumMf5
lSr8xBFIQVRxXht+R1YxvZU6cybTLykfVWBF2hmkDTs=
`protect END_PROTECTED
