`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s9lkQOsCiiDnxUCcWS937geefqeLBIYu/5LhB8sSYhlwTKqM9271RNMnH3Hv8Y96
YFtxjsKlEMiIu8vHZ1e+ho3XEfRFrxlXDpmZdqqw0uYoc2QbwEtL4dxtMCHtuNQc
X9B+7Eyi51L66qOMYqIOh0aYTHswIrB8QIZEPgbdauu+Q6J+zObxqT/B7IR28424
36v3SkczhVG2QD5tlhclLhpT7U9D32Wyf0DW6YqfkePzG9U1WJjLYu1lkDZNRaMf
BBMb5lqian8gNem6DoQd52Cyaj2+puc7DMa2HbKBsdMefRd0HoIk8YWbFhUbZ2mM
t2yYJGEn5anmEaIlh4kgVx01/omhRxPcRE08FTkToFk9fJ8uzJ5iAYAwGCyz52/J
nDFU6ct8ogCT7pi7BkvUMHKwQ1Ajrt7Hqst8C27JVRFANjbPwHSYuvonl4Gd3+ck
p06iqqxcRdu4W4Nsn0tMTjVSKC8cAyK+hTjgPfwupadEcUpCyjzDzNiKqYfm2BRP
`protect END_PROTECTED
