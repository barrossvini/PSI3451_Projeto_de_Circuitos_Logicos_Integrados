`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mXg16ZO9Eyy/wElEQkhJcmoRobDw/Po++nVNbIA6wlnPACRcdySQqIKGZuFLRPEj
fVBIDqk6EGgMyd3Umh3p1HiriUVfJ//NCzCVxkKsNzojw8kBw7Qe/ZqEvEvb/Vpc
7+SOH9C0+jm0Ap5ko2y8A4Y3B0t4MncdScYvgSjlceZZCzdwZOpKMrPH6mpFDG9H
sylRaLjpHsaugQ/6/C4XSykMJTGl/oL6QDAOT8aXNd4T3GM7HsaA4DzlZfw8NY4x
+6J2usP2SYtD7b6roeDK7gTUVb6GA9GUZVMUCq3JiuZKyxVCnMhd2k2dt+o7FqqP
huUsY8Fx5xcz/PmrVOyADaHB2MGM0Qq4QNZRMz0YjGwqnN+nqBKsEbvkNbpDz6bi
SP+xTqrmkWfwtc+7+Vn3v3ZybWePOFd2EPkhzGG9uxI/OtUOElFV19SWpv72AHrd
UUsRYWbqY+H+My0VeBO0YvonamjV3ZrH7QKKwVES5AwJsqf1+DyDggR9id34MxnL
CUjvqsgLOiUErR0ehSYNz3h1Rt/xbj6fKS8PaDDj9L/Op1v0LK0959/UEShGKSZM
JfkAYl1vcZtYncDxJz6jcFbRww7aL26h0NZA3boAUhsa7uJNFuwqxcYffe405LIM
VlOmWz00aYF1fJDuski8HZzhzQiM53xhhbgTzR5tHgY=
`protect END_PROTECTED
