`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C1D4zxN0Fnb9x4vuHgL1mBvM0eahhQFrMGpn7e0UjyXuxhxw2Nl5LbjO/UrKeufX
AREzFNtvo4QgMQyeOQZGyED1SIag7P7EEBLiDIwRmOJ8Z5VbHWHvrSNht7PE5tqW
r5l6q2u8T953BVe++r72jL7kvSZqR5SpM8rtMECBIuzgMBvf+nmYYeswkf9nocUj
YALSrZUolWi7AGRtLdOrY9zxGnLh034GB221OjscE2Vz8YYaj4f/S7Yczh18x8N/
bPtP0nfrNLVcd/7DCuKQwuexBXRxdE74/MYxszuOm6FxQcGZwiqEFn6/HI3j++uk
BoLaZlGoL0be3xNYu+4it69juMy8fSEndXK9KKoocJW7mKrSA7+pmv7miGd4Isu/
YOXWMvp7SvAQ+ZQwbOmXXx5DnZ0L0U/zvuyNn7Kp6e2hePnVtYhDOMS41cmNaFym
nynNjIrIfzUC5/zgVSVplWsfyktkFA9gLhxTJF3CA2Mv1m0zan8+jCwheUaNuOU+
Lqz/bkiIs6Ojtjpxkqbv26/KD8yTd03DxemF9JgJGK4yS9SUMOdzeyW0bcifHZIL
W6FtY/vEk1RFl4xH0H0VePxeQ7E7OJ36dpNp9ErhusJTzwxwHwsRRt23yRmziMK7
NH02lLq9tzSOekTrglttXKs3mRjq3G0XbkcB2smQOg5yiPrS0zzcJWm+kDsW2Xzd
S/i8EicRvb01JWyWtPrvlBpfxgNe2lkGF29C2SrSCsl9jp/KomifXD0lpRig8A+9
+7twsXOfVkBtTIcdWYNSk60u8YsKCvxnsw3Xha2UuTy7eWXa0Kl87I+RmDuRjGwO
QY71XHYUSx6tZbY3O8ZUjSpMFP9JzBAN5xcVrkCB2oS+HyuZ6/NMJqiV1O7AygKp
kjgt2HmyBi+5Y+VfRvJ5A0tOfI05KlPwqVVJiKGUW2MUWnToU14oXGS/CAKg4Z3i
OUcaAbDaNyomIFLZmu3eCwHy69gSyCdJSTXcvtTueOehdlV1JESC74R2x9ZGQ30h
gWJfQGa4H3qCuuuJcyVn43n+8SnHxw0VJDx/8qTHwFckg1VDvQ7Gpz63YhAi7AwY
8Pe5Mt7ChQdrMPZxlaW6Wje7Dn/OnXcPgaWR0jtrbs/jz/+ygoX3o6L++2KtzEp0
oH077Y2M26AaWbAP7PaimY8ffq9MiqgdurSr1lzwTt5cb8pEosAGEfZxtQnnOIYq
YaDQ5m1ytrX009CoUaZvp/S+q1ZwrYbEBtT6E8JRA0vrWy8O59ScPrcBHARDIHRo
me0nyaVO2FLiH+/fdCtGbBmINfWK+OALTZVoPUa9fgnMhGaO+5W1rlIB1+AkxQSc
cugwxnItwgqB8y3eE1hP2X2pjq+BeefER+1BddHQyGjO8D406imKihzMrdwoVUEk
uFBP9KfwpC30Q3ba0ElQHH412BXmMJeFwgDaSI5g6z/BtGdtO4plq4SV5ZZyo8rm
pfsgFRCqgUwL6r8df15+zuZhmVGXNOyhhPoNjpjWvoKlstO9h7qArPCwZXtXKv/n
But1kD108X3Ol4M/W5huU4JPFRHw056mhEPvzb6dr6rm8nUKIvCbMozh9Kf5I9pR
0EzaGzxbOr2niJ4k/c0yijWmZiGnfy9CxkDcQU6haQc=
`protect END_PROTECTED
