`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UrixA3g0sCYsWWHyH6QP1ExBzUqMEI2Y+rhS/LvH8HVDh1Zgq6gMOBsFKcpw87G+
z03I0W/IG5DLZyXJVX7yhbHQIXWYgCwwi8iG1HuEoRkkSIivkcjGsXvOeofdJHTL
3bMZSy3rRGwWxHfw4egt+m9uE4bBbu5mk9CrkuxPmZeTh+/dwMyg0OmD3R+ve9L7
HVyTTJSP996jIPOKkYbdG9uFXWtOoRIH+hBvC9tOsijQeT8+bMgx+cdUII+NEb43
hYzM883MUuQO1zdCt9ANXPPECWpbZ8yZdUTQYsfxWpcGrWCu2s3fuLs/d8O46txg
mAm8bQFM9qKi2/BjckmydvdDQLWvk5I/IcJzVBWKVAVp/otPsFnHz5B62whuJQTW
Wsb0SxFJelG5iMyijaPwHoQAqJ88Qa7qJA1yZa0Xhj3404eCVXkEPZq/2m1XxJOH
lglnenq2crKbqxk/G3rC70OIWx9xFeNVEmk5LRly9ur//lQDMYyRPNMvEK+EkQvO
pYWjcWkj8fNP3fWIit6cRvDvN8IgJiLkLoHXemNeIU22B1/NlX8YRD7TWb1b8649
lF4sNeXDHXZ04bUXt25vW29JoLFwK2Zwqs4he07JAmnPNDLhkH0bSNk7AnqyNB+u
NiOq/s2Af/m/6ke2gsAaTXniWnoGeaijmmICjNUnrq86ixfWH5L6Ne82PGNRPBhF
wmCA/Mc3VCWWjwwrZ9dBpU8yLduW/RzDh7peOeEwdwkX5gGQkaS8JTXZ+PglZhit
Ppc68Eov9FZqf9fooyerxMhgv1BZ8p1ud5UnyCNM47kP+KMVCFN/7xYBtbVv8TFa
HvD8+mo54fHACO6hPyi8jOw6Zgg7D5/n1LuPT6T3At8t52udV395A/G4sSVxOc3S
YEv6qJVXRD+94pajimdn/ZC2eRpK/6y8k1o7WusEYuRVN4U16Pzq8g6mgWO9bNm0
ZCB+w4bhrBVL2BSWVWqWRFXjSmWVoCP+4sW06gNYhfvwkpNRHqhMf2TF0VmmMi5d
DJLZk0hj3j1y9RiZ63ByQbFrjRirKk5qkCJfWzIa4Xd4GlXlJU8mS4ZNVTPpT8tc
QolCSVgA4AISaU3WoKrJVPR2DpodiO9hZXgds0fJKA627Iqevv3NgsAqa1VUCCY1
pL7fwywLrA8Jp1E3xVSHXsDg8qQfCOYP65xDHdRen9vRdOd6KhDXJ3xzMUp3pzDx
Wrh2jeDeE4WChSdKnGW7eNvxaTSvQgdMubQBedPJ/E6XmabtK27WyV1HCMeG0jBm
I5TmaOt2HCPoE9JbX7VcDhtHUu3Lx9oLGU1plTCan4KEf0nSWPZbVdHe5G4KNm8I
2GeBqxMe2JSq9/hIyX4VkW/mMN6jsl//fSAPbG8QTwQG1kBUHfH7KOl4lquGuvYN
h5tLPnLVpx6iAndPW/23GXKSEk4ApxzepayH+ZINAWsfV/yE+mDea/V9IxC9aBuF
hcjIwYPkd/oZnoTpECv/u3Y4blhJDy11gm4Bj86ayG/A+oXz1GZqziuLCbEaeWrc
zLa4jqh/LZDcVnwId/NLb0Fgvo/Ad6+OYvY56pSELce+HLjkXmErFznhkO3bUyB/
6HM4KXgNu7HIN4EaBhxChnuYM+I60ozRuDPuC7ygIKh5ZVzu8/a4aktwL4jIS2rD
wDL5F+SqzMhX9qSv7xJwoWjNGnNviq7XHX7fkfGG6NJNLfeos1+4WCT7Ax9sahl2
NM7w2buTZ98tcGRrXv71GlWBrgMhx74lAapBv9NK5OuxOJfTl6hzHJ9F/pD77aRi
yHGBB86KSt/gDPwpzuRpY25r1nHUmzjssp2iaEhLEImcRYDd+MjpAgaeVUFxDMx6
TItJ/OQX1oN9Wq5b2RwEts1A3ZALkninLO7lFhlqxT/rO73Af6TdCnxtbhcaIJk8
PGkq5S63rXCrTWXbOM8J4GjMHbrywGsq9g/K3UwQQOj4pRBYa35gdPllZdjfNAnK
Kk424uUes9iJMwxaeBljY19hzurOna4j4Aj+VSzb2zg6qT4+eb0AG9XWQEsn6RT+
MV4KeZMc14UR3kNT7Uuyoj2o6BvwNzq6I7H1aCAgPsEywt+/67tdO8cnoIzY6uEN
bq9mZY0sS3wec2O73LOsTgWt8BUeqUtN9Fce8m1mw2hzcQXf97Az97CRGEvPsE6w
wQ1ZISTgSVmV6nt86RWRHflQvSLkHghRcRYfXUDwi0B5IA1a+QK9FemQ2S3bqwdI
m6pY5+c8cV34Ma5aiTCE0c7xMIemwyQVd5/kVmLi+8aVvQQZ2564qE5hIch4fnb1
eHpLCOMePQQF917+o0zETzv94Cf7873gbOl35c6F68Me3uUYdg6GuzLAjj9i9xGP
p78NcWbB9z/x9y5bEleBpHq71mAPmLtmOpVyWcGWM5YmBN6ewddyyfy4nAd7GMJ3
e3CzIn/ahtJ/kroDT5aiC+O9S3/WZzEEOE6eUAEQQ5vHn6vg8OzNjHY0dKIYOi/m
YHhOCoeavhEUnK07Igb5WIrEpQ1TQQ4Nz+gGc+74MIzOtcQGrHZDChiTzwAD5m4P
jEutyTdlxfy7D4Wl0JAJcpOT52bVsdaZEvDXE1pOgj/uFrNS4+fCzqUZpAd4alJw
YAo7QT+KghHRzxpRkHgHv2/IIVw+sEPkrceq4kE8yfzva5yBdjTgmRKnVP4RyI5+
UpLEgyezF7rx4cx29KhbVI+A9nAH7mQAIM9EIEPjHDXCkey7YpjBGwnotaDB1pvM
BGUxBURcW3ycMw7vTGJTrzuakvzLNhIaQS/zzXqUgXmJEoA+LF0PPUslKHJq2Ac+
3yVNGWmTFMMZm5Yd/uHZjRTyjGzdicS51oin8js3PcZIYVaJ57/OR7Y8JhIZftPk
C0Wjn3lHmhMP2TGQBuH0d1Xp8NR5MVAVIE5Uadg0nsuKaF6a9t61F8d20m+xjeaS
GGfuWH4+b60Hyu8Sbr2GYd4fG9eUQWqEosD4luSlyrZqk8Kike2pNKjMCsE2TgIV
fiVirUPEqNY/V6aDO5ZlPF5AQg7oUKTTK3bLJE5nUSHIz+xJateUtQTssM3k0sUy
drDlMdz+ZC8XPZlrKL3OCtpLozV05Caef0seHWF6rchhB39o6enlZvu+VOWlO1fi
YpYbxJGGbAPIQLxjpERtTN6ti3P4GydU1wOcJaNIqQl3mmNzxkHNw7p0Eh6/D2PO
6XzZ7bUb0KabRHqjkSZy0PPivg8IB+YowB2O9IrboZY7DKoJ244+GqbzCllzbzE6
APTT8b2uosLoMIr2CBNpRTg/uQtqXyR0YUUDB8srFGzq8nMab1Ngt4IaBWOKhctT
SBoTW0qSgtTrlXLvvZgtbBE9qTbjUs84BORgH/qHbO9mSq4cxyOjPO2eR1AlMoIe
eefE60kecVqnYlIT9OzGpFacRuoq2SpukEGkTHZYJAqD9ZW+hWqDScEYZihi2nAM
Y+MgZvX3aCEZZRqhlDa9UinZayZjxJnasR+gdVIeWAyT64Ds0l8TG5Ywjgio3JW1
Z2enPbs9liOveQvYe2/uuFrpLGRjU9XD4ActavXl+4buq825v6wvQGaZdib42DAn
J3ItD4bwKooBJq4kj7gar137UYYZ8aQJYSy1uVzgDMDsrKNyY0lL5dN0pXYptf/u
PmMMB09T6hhmF++GQ9w4tjGwTYSMA1nqw/Ykc4jgiDJ9La2Baaeqax6ImvhAtSnW
TrL/jdj3FFJTXj/zIONlRRrITDJX+OZ/iIuBzzn4uFMsYNrlyff93lbCTjKGeR+t
8T/u3cUymP3+uEtCiffvETSUiihaQqbMnD8PeE2HiqacVxFlyeVi3Wlxe14G9Ymv
uivgroGNStAP6EGipBsr/rdrpO//9Gb31QgE83awScEDlvCRHmkN0OVntlwalpX2
JA/uuTx9XYNrjb1PVfCDZwuQSY4IboAXaJpQCrSn1cseTdcTPRAC81l9jBwogABP
UWP7pX/oGx3p5jjXEIlBDVqo74Y2YOan3ndRz44e44xIzWFOgt3uIvVS9mFWwJKW
XYcX61xuZPzdDnE3gW5coj7xMcGcH8IcQl/OPqhwkzyMG30wIF9hW+DBr4146/nt
tTDq6xcv+LFEt/FR6TvUk6OFNyXsg6sFNFp1sA0scDWpGANnBSFNz2zjWa8hobWA
RV1lWDoU6jsfIbRtB7H2XaTM0xKThbuVQ9dDVwdWIJxhY4IB7m4mRxY9a8qDTUyc
c6xTcLAGVTnxFyfs/fA++lyQr8mDmVmVfVk/LFG33HnBck5tYvcTZVLX1BqNQ0nr
QXxp8cKc5BT9Oe6RNrVRjue28iX3Wo7DuC4QnpVAOpXUZt4PUGgdJdK7cqwZ9T8w
Aq+2aV+OpPbvJcIahb02VjPuIauXTfaOMNhq7z8TT9Rtu6f2dJFtvI9AVXqGfahY
PRtxN1bh8gaLPlBY5YASvOdYnjSg6857RtuVpi9kEZZMNrgNSI8QTbvKwoQZ9smn
mJ7e0YLSHfM9ZirSOlO8E642lmZq4l1/L76OlhFAz+ZlrPBtnskoZa9p4nI+TVEW
WEjqz69QmqaGMKX2mxJwje8Jsxzr/UoBJ77J/gHIQilrbjLFyRAwKkIA/jgOtUNU
Zl+uuwTR9RqHokYGMQvr8lOi+kOS6Jipf7Jvyv+M32jf8e99q24jMk9ynMgXV1o8
Plnx21O/HYQcwpvadFVv2NimhhAAO9+aaFqJx+nimYVtmVaQXG2/5REhiNl2SUbO
iJLt+PyYFtALr1b2xjX8/4KjKU4rTIkmfbiVXKbwzJtWdzzdpWmXzrBIeIsYd8fq
6+YlMIMkOgnTDfgKyRW8KdP4M/S1tHxwy6UmhHJJGvtpJyLf2dx/sqrMPMZB+Efd
2Boi2ODUsLzX7WpeL25McNkoXCHttLtl7nR1SbAqnCZ1tuXuEABHJJhouM8YFX1j
aU2SJ1WLKUI8tCa5UsKwdjXW/bifEMfLDzeeGtyr/9tj5t7/dumWRjeDa8NQnphF
iSpESgyJ8A3Qt2CNtpHLQiPkwvrdeUFqJ/u9UpGpQmxz6r16f7dN92FIUKzKwRXN
cnRYM4/bgB5Zya/7Xme1bF1kCMfkp67o/hVJDzcQhhP49pcAdeS70KLhSAHYoEZv
VOy8XKvxOqtvymz864dkJzjFDzp4SA7FPPtCk16F762dx+znEDQfbFgSqYkuphk5
J29hp7umti0D2o75IlkNu99HUtBVZd9fnjffm9B1/7YZeXebVShW/2vTvGRBtGlu
uZmHXAkkSz4hVQxzj7moJqjoCopKJPWjEErk7WGXd9/G5psFoWNRu16Tj2e+wKHi
J7IyQWDUk5uCECRNKge+l8QI0/F/DzDVgC0we7GAFRqfYRyVhfgqkgd7pJF7XZlD
bEdd6FEYnON4B+DRpYtdT8ClmQ/PCLSFLeNJWd4rhVbz8gYMJ1Q28cHc7Mz5vlpV
4ZGvXIG9Y4xusci0Zb6vMMstZzQlg1AlE+ZFDHsSdXu3lpbqfN5a77WpeCBuJ6tb
PTvdkgxmgiDfLuhrlYFWf/fovnoJJvZmam2Eryu6BAiY7179Wie1pqt7Kbw7ski/
zGq7NH3/5wrg4rYRbVJ39aIuMlcRoWSviYZ6l9/PpcT6liAfBFm7ZRELZYXkxmRI
MEzHwq+JWcAeULI4hsQj2E3LlqpIyvnglCoWroH2l2oXj9RKFo4Iu3EXnhkySHEq
0tF374hzbZnGCFeE49tup3kO889zcOhXRzHRVfDvAMCw7mfypScUl0GivOPqTdZZ
yPz+jpxmxYaK2K0X/W345TLlL8If9/+lT0TcyhFMlglBdYBCLEtfbRS+/CBO/pOY
Ux5DW4FhLPdPKod8cQ8MUx6mv2T2vg/QUnm8nhZjPx2SmNXBj9ztSx4b6Nr8oEZM
opZFOCYWg7NPMkWwQ2SIy9YJNDIddkQhWmsxrQLDtenE0hfGKtyW6dj29z6HXZKB
sJnqLOkfPQFVPAq7UC0t0Wm9zrbqLAZ61dhu5pSheY/t7vOpLcAnglmOaE+ni4Ee
qSiLnwGAKUxXAh35DYJ2x9gtiN2ordl2gJ+Dnpt/9mXCMOBw+sBatzfLrgBE1kmC
YOpGJzh7cS1UlmvVBTjh28R5U96F2N32/PTzwR4/QpgxAqPINDVfJEExXbRfDD7u
W3G25lNNt326HVh5L7BtWlX0bLqxLX207Q6djXI8rl/O9pJQlYNPZ1BABELCh/4D
ILs3gav1xiq1lDxUyA9cvptX4kVdmGVDQYf7tYX/tU1DBI9DQZQ8bVvlTAKEMott
AjZwDwivW7eIAdVRc98mMxnS7RMkLA5gsUrbpORdL7AEbVXxDKjCQ30NuJY/C/3F
2+/O0V9e4F0Zos5RcLlP+yemeur1Qzm4iXTTvXmLKM9sX59GeWKJHu/BjHFAS3sZ
9zKI2VF/t+lvFxkP4CaY6ZSSzQ0CGwzLICRqiBmmmY462HxmlsgVfMgQDJHqOkoU
/kQ76yZfsqffVV01cxLbP3vhzQfchjC14QuhgX7aGxYyU4DVwfZ423Jh7+cBsj/D
ODMOBXhSG9mF28wXxd2udZI1SS7XQazbvM06yhaDZtWx5V+odQc0BwolT/9ho7AE
/yOMcEnGFCGu9PvqyzgPW7rgAmp5JX/Nw8Ut/MJ3qltYhR2anhed2NtpjCyalJBl
oacJN6L+S4wqtOyJtSDL2D6e+5WCwOHdXnIV/1b6pf12KJrNzEyXejFijUW359up
TlgdpO7ztXXj4++MFDQznDtYr4bIDEn/sS3cKirHJ+MIRRODeuYN8189y3T0SDf5
X9tiQJHKehgPCFWJJOI1C3/2PyqG1N+0inJyg3QkgSo6j/Sov8mh5RjSUbf26LpR
1mEytANtnIWPh2uND2NqXrM8WMtTIAmEqHr+ob15afBMLaQRqbGG7rmL23uQz4Jh
E6dV+4vhDyeB5vX0AO/QXAg2PD/EUz6BDLFyQwE9QW31y0zGfe2S1KY4cGt5wjBj
PZcCImikXR2Nk2KSnJgkC6+O86ss4n/wOYysJ8srmwuIs7XKkF4zN/AaYtGaYy8Z
HQQywD2ct2TW9kmZptaiDfOCKejAGISpWWKoESsnTO6IZ46yfpvqlzNVU6XaO4cZ
gjrCPKPVgk70VLig7GygJVZ91ykkWF5rkDfjz0PdLlc8sR2X5TRGM9IuuaQAsjXp
GU/xkBs4CBHVMebSysPx+IAkecEgLU+G9M/YkGxsgqiBT/LbJXW3X3EQy7oaHDA3
RfVQ4XZXzGcY9dv4iXDFWnjyYTDN33TbX5SWgCDtDbDoApDckp6cr62FBh6GXSC+
uNWXlL54gNDyYzFKUjmYghtOf5s5zSyeDmVLnRDGxxNt06XdD9nLlBiamWVcb1be
t3oUBFX8tuktZ3dLj3+UL/SMUFcfBPq6cIIWnBqx1Xlbw/oydL29vyHhChrULc53
GE/C+UrmtssSKmCVnu0NYiWc1yqf2hg4tjGjSorpkjotc5f774pGS8nt7/Q3qj4b
fzXDQmQxvz441vv3W42EZAiFaZz8WAiVG14k7qrHyFTO8Qh/vS6JwYpDchU/+WS/
cYf4EtsaqAdpz8qkyEeYOpM4ibaSmQORsC/7n5qJvBP+EG990Rw+JphjTMJ885i1
/+bc2rgm6uRVkkhEG/l8nsAedKGFuN/5uhb1IaPMeJ54G8N6zhwwYWNboEA1F+2V
tbDsuFF+497fqXdFlagLc9fBqQiVDgqbUGjGI6T9APW4dAZkEqwJLW+OVGX0ZqgM
1iICs6TSFwFHpri3C7s/tTwUBrAUs8aHzDcAQ3YabxyNiUxaH0JNWfsGBpyVR/rE
cuDWjS4E8I3nQglH+T+DoEbau5egJL0hEG7Za5szbWcijqgmeAVbMFBwwoa8Ycjd
zaynaUUiKEy7HVJpYgmre1lvWMseHBbzNlOAGsN7DKviqZHbAO+pXDBt8gWT8tmH
CzzB9WwCGaMUbJk5j6QJU/0ThAYwKHaEWKWubXsVZVl5bK6WcYq5hUtco2B2DhOI
wSgOsZRCysLKsLm1NxE9EOt2yy/ypeqlrJT86QNIrTezREASCORrtGLabgqn28TX
9lZHK1F+O59lW7JfR5UA+RqaWL95Jlkqw0Dx+ypgEFV536/U2Q28gnV5Pd67yQwm
GbzDNoPtBLOK3rNU6KEHfmNwzJRURjzVQ7kJBP7Bxqw7vjJpw5ZuwAg18ims/noa
d+txQOiHw4iwzEZIUxe2zxyMh2hjDurMwmTg69VGHZPuJ2di1Zwl4MOGkG9i2OJT
CW1r0j4j+jCu6z6W9x4ovPHauQfGjYmXkiykfTQDKu7l7Yi0G7bBveUFNIxD1FX8
CXzwrO2vrZh1WusJMLZcH3lFt9nnUnFMFiwgHPlIhcknp5JlNPMKIXFuVMSJI28U
hJIxrvGiYUnIRkHVxhmKLNnCk4BvFa1/s4WQvUaISfNjW7CCuYgBgPd1GG2/Uwi+
6JRXStWVrA73BlbYW4bOvsd1Y1+2DPaI3Bn5H3ZiuJ8tsXQbly+HH2YTEiz3PQQL
aOM96AYqCc2k9D919PgYbwL5nWd9UcJeuRmta8lKnU99UYQn12IzffGQkCMbakK/
A33pDrNFQeyFpYmWo2+eensC5beekAJ0O7DFgx07xm9hKuLWPvcpKWWfQJAKXUKJ
KRvjNWy04JJjw9gJFpCN+lFJ3a8k/PRrG6H9G9JAku0h07Gc377JDh0w6379xnBA
d+X+QeSAh4bC0KiNBkTEwTA46SNl62KuYo5TvT9FSEqA71JC1S/xkvdOcpD+TZdA
rkGKQFysOzceyCVDgPUswXF++LuZ4ivL9vTbfbDiV6Aem9onKeUuj7Bxt8DG/9r4
Cno9pPTaVJr0WzPFOkRbcyymWqD/hFLga9JmsTmmJks2ezLNzawg76bSssGBTR1U
yZ9EU6PBgZ4zKB0wuwxK/gVwSeHCK/B4vmdSIqO3qQrNj6tHP04CVTOU2RQ/AvmR
2GcgfIaLzvLtHjY6sRv/wzEFAFpOprtHEZfGA32rlKz/sNJ0MfvFIgFsgOrSx/jP
PUsQc6twl/UQhoJEdO1tw5q04/c8y6141Ldcpd9bnNRm8kJaeNXri7KV6iLtJPHp
mXZR0Qn9L9NYyXcLOEIziK8ijezl4tkeDwuXBduIan78JPsnkpUDzAY63u4jfXhe
jqIRYUxJ6doDUDNlf0pWzPkrZCANe6hyknRrqSuEVKm7VpeFXLNOsG/nhoirpHEh
cif+f+D1G67UmcpHg6JOsbsypoRqnwBeYNi7p2jDmQETe5aHp5bt+81ZK91zdtQo
Gd2q0vauq+Wv8ljjtz/HlIH0L78+Pbf/cT3hTqdVzqt0ECyg5Fw4u1KkgPjSGJ7n
DWvJAmeQxkeMpvDvvXhh9Jou0w1Rpe1qdkV7D30FZioWRga3964HdSVgdE2uZgwf
5FCA/PTS71mC3EhfOqUH1/lUZxxQErJcjU9u2QPYWmB49tbEQDKIAfiYPaQLVaGj
oxeF4UNG7d2ZBYOJB1mEK94Mu9QFi0CUQgiBOmYKatWtYmPJU1KH5DIG+hRVJhQS
Cm9mf7nwVGUPRTPnUhfc6px/IOSfT1Rr8Bafd4P5+hZkn4a4wNdu2haQTdBlpmet
6kprCD+bGz53ijoJtui0S8LFjiqaJNfyjo4WWN7WAGuxG7Rap8XRg+GAeq0yb9nf
Iddp8kpD2rQeg7g5TGaz8ROlSdqie5eFNyKEr/wQ3vCg+TZaYtpAsClVgpBLrvJA
IbPYaHwRSEvtTfjqtmcEIRmH0PVlfSJf62oeWcOxJsio2FG65Xemk/sWCVyhlTsR
YKlNvcYCeQ0iAt7E7Eyw9u2kRQDOPO3jBrwLote2ejN0ENYxwpVTQlcDcr/NBElH
gUeObIE7l6QTlANtkoIfmxdAt+I5kefwaC0ds5Db2OzHk2Gb/neK5ybVo9ksmcJt
5MIwmqUARhS3Q+qdPivkcMkSWlSRIweiLwO4NEhB2e+d1iH1Y8nbQbgBTgu2Whgy
qzwMHx5FbOkkFB6XSoR4wFqLsSfztmuPTnaXQzl26Ir8Gw0ys5Wh/OlETXJ9MJO9
2kEg3EMEGfi4BOWDmlBNinU4xKqLt0YTmC8FvEKndVJNlQYo7aCUfceu/aGqboRx
52/iiCpKNz10LI4a59QYrnAIK3duCQSqV9hOauWm611eTKPV9cmdI83cobAk40B9
FXmDGoqS95OG9fafHusnhtWVKXmIY9fiEy9CqEXvbm2AGhSUYiY06TXDb+C1dn2K
ih7rFjrShCkHhbk7yTUAVHs7jK/HexvHCbFrKbtjtg+zBjLt2PpJETxRtilJTLg2
GE2jGnwvOwKh5rJa6IFzpl+OPZnt/++bfBjuoE5oXWmu2aLXILy3VBfjFapbioRX
H6BYHzz1KeqU76w6e3bzN3wUnDNJ5pcZKgaP8hjXvQDU9/l+WN6Jd5JPuxD82krn
QCwvyhGzbYHrEkPrAG7Ynfm+q9G+axfWYFJHt9OUbCU4rcu8orN4psEJlOi06QXZ
RXY41fIpZROUA9yz2SeSD4PMginOSUqygc5Q/M2/zpV0G6pZExalxOLh5DPpEwlw
9SKPLqBsdVGQYw7bkZ/zUrzlprAUJxM+BBQHyMhYmhJB2X401pMINwqSbUh9QTUK
O1DxF8B5R5nsi0J5FieSmmAtyrcGyTYJHJMZU8qmR0MZ1oOP5N8hRWWRd3Omy0wt
kL/7aw6dCKe/pLYi5VZpzHEqZUD4bKrCuI5pm2pRK1KiHpgrtsHyrUiU4vGfyZPj
bdvF9gsHLDGE0/fQ935CuqsDOSCCqJCRoBFnJ/mjqYb7OfzfxQj6gzDs0bbEZFfb
DgschwnZ+LvBZupxEi+Z24nZEBGdzjWplXXe9h+VRDBv0LCMGZwMHHlIfrURw7FD
yeScsk0vXIqAZ+a72LQKle/fbHZSpB091cMRp3tjdSQ=
`protect END_PROTECTED
