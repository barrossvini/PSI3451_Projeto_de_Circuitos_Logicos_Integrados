`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bnZVN+xCnNpjPXqkSySQ3XMV74YDgp7SSZgqIuHe88gejg1NF28XLhpqGBy9qCK6
YI+dPDy5b5vdwklCFI9We5aWhKYSQj2CEoCYHc9JAQjAGL1JXGGjQULGyIO8w+xa
dRYwNfUthasmpheSFMGlokDhVYwIz+lPw/e2memcdXN2/fwP8PmD6+M3vRGv7B7n
VevLAeJchnsdbBlSuCGIT1JLyJZ4zgoH4ScAG83xn3J1YpkTxZ2WB1ljH1QP+4hy
ZsapvFyvSXrgsu5iSUt4RsYAtynEzfkOHD+O0BMpPm8Kna61yeUUrRjCL1ctvb/h
cqE0ddQ3SnW6+REvwOl/cyd0amgPpiOW53PZ3lSQzCpA+kAIgzIXw49JKhP8Vwto
LzFhI3TSdRRF9rXOvT1IR3ZDnE9S3e68T9HnI1gXZuxiRqbZi/UuuYV47iVx53c2
ZH2ROBXpfn9zcLCi+fym8VzjGxiFgGaI0/PHsX1utPJnbD763FXZPG21J8gn+QzI
GJwSGgMs1JTPW5ffOWznKoqTdMksVxTVLDmAPsqiIi4+iD92Q56M+2yPQR+hK7OR
u0j4RS6wFp0/ktrYIKYnUGZscWeZPwlWZirmRw8JegwZ5ILAj78bP6fZUA+Btyud
FaQou9P287sihXm4kys8itgqZzz/SzhYPTzp7eRIx4yY4klmR43NfDohlclIoSO4
LyEKPRi3tdEbOvkWP7onTBX0CdcuwwkuuwDS9bHdwkqkDN/Y7qbgP1ZrH69JqVaN
BOsMzDF9hOfuJ6Yb20fhQftPpuZHtkxrP3IswOioITVnxzsHuxKvaeqr7wsFdw/W
w3UjFwSgqAkdlIQIiKUdbcC5Z1504t3qhoV5zfbmUYIzLLR+hSpM++PyWAJuX/1j
sd4W4J9GIXq1tPVoZP/lOPTGi2HvYtg4cNLqLwgwlVk77COaHRrt2c+jv4Gi79hL
bEzLD7wH4zyvRV16wuUY20zobOlNaRV8kN9/95XFiA5W2DBWrsF3p/7gD0s4eSv/
s6sRrNYugh0hNjo8ndfJdG8aQPpWEHAR3xOfxV0Qzc1c54HYLiY+6EQsrgAKQATU
RajhWRyC1znE31SwDlibGr8V/6KYgMU8v7A0Al+3IL0T7OBrC0w22thFeop/91ij
isli4TiVjUsf0sz2oeCLyPbk6nE5sERvTFZ2FRKTA+lr7U64wdVl94gj+Ktt3kOe
uBC2EB8zsm9132RI5z7mW2myVbBl1HC/2cnpxKFeTlZzjP9O7x/Mnjesjurv/g2r
nAcAtN+S2TmW8+oRqBuS4LgCqDWbt2b4/nm8FnAD+qhgqrN7VrUttSvWsJSLX5Wz
a7MWsk6811rTsLyNQhnxvjOwbq6M2GX1BW12hd+RIg+WJoSd0cd4dSQLeHkBJGbX
eoSy6FEWN8UMYHrJMM0UtgndEkV2PQyxa/zlhxCeIGHQLwVmc/BiLyc069yFqsmr
booAU4UJlSdQ9Lu1J4XSDY/5xoU1RRmvWrn14qDJ9fpOlCoy9dqYP3CWGJGiYokY
zojT4kIcjpgdL0P+RUPBeZmW+Jx2pxNZ9Mp8VQs3glabkrN2/JPUfuDCwQO0L8wi
sq+DSZ5X5sYWjNFBn5ZYI4x5MLcPjYQzoUPZFz6opSoS+Jf6Y0Rnplm6Io2HNQ8d
Zt1AxjmPl7Lpp3hv36uDALDOxY+AZk7RZW+n6K83hsDfPDnfaAnJVL6fkTDWbs7w
WcyNWTP7zql+1oV/0nyF7rTiN6ZsQiQEugSkBsFUOEkxFO4nmUuNqQFI1iiYUbru
`protect END_PROTECTED
