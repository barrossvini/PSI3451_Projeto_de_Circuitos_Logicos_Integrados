`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NNt17k2Z8NHFBy/LdvjWHYhg6kxPC54TDaI2qV3ytCTe/QW/ik+lAMYPa5Q/fphf
gl5a6KxWuC7LYfRQRLHNRmJMQie3vzEGVdb6doVLftjgEN8cjHDLtMkCUF+OSZ0Z
AttePx0/LFuX9s2oU/UtoIpzViZP10+tMNZtQKfdWQ18oDAaDdSCzY5y762W1DHo
qjUb9UlzOobT1qnhu6xL+OGvzvd/UOkXooEb0k/AaMMNXsVmVk0V/3jJ6UAS+LvS
490tMyUp0acHnFV9f8srI5DGz0kUTie4+U8Q1Ob25r+N1acU2KgONsnp3pWQ3Rjn
o4fkShbNvLKUJKkbrsQSgIoYHLYqM+WZOIf9G7eGZOmVm8NkiM26S2rHoPha7M0Y
0IBFWY0lx64hR7Ef65G9xcQQK4W6TSKzteenioXES9qGS/7FiWv+U+KQpxt+5G0n
wT9LiYwPMjRFossgr7qo2DlSeVDzAKdw1+QNn1Yr2Piag5IIJ0vTWbthgLg2pB/1
JcyKqKmwkO8sQ/y+Y8GSmPbNvMW+Sxfvyq3BYWB0/W9ukPK9+vpIhtclnqRzfxEM
3Re8W6IfYRsV6/zHMfqXOif4Kj0ggfbby2YPOa6K4xZwSRShbjonmMS1Ndi3pFEC
0m/P8HLQ40e1/f9kqb3lmfs/zZ+VY+R4DWWC/+CcrOG1k4IcwMniR4fQHnw4cfTC
hJSin+H4iQVQv91pmjL1hnF+np8EWbSGBRAp9QDK+OGTGNx0hBtF82OzgP2dn1yh
BFStRPg82Y1+C/dP8WrG2t+2gPEmxAX+EKPzS6YVe8uwxMeFp6z+8bCLbld9S8lU
8HT3YsOMWUxs1HCmSIdO7+qsQe1fSR9sGNt5flrvjR2kZpvG7gEYxrQ9mtK6raHc
6fNb7td8HO8LviPKnG0hDGoobP+M2oCb8xp31n2DJWVOTeDhq93YZJ+BNkFjeYl7
ImJXqUCf8nmmQBc0nlfEtWTV/ddcvOOl4SY181/O8x//+qAUqJRwi4/MMCYToF0R
zoWo2IS2sPgAwtW5XXq7n/+KrXy1UTAGmifvSNMUFvHp4om7DPObZKt4jcdy51bw
GFW2K5YLENpb4oJ36Vy4+W05OlmxRwi9L+WPHRM2jsy2iLmMCb5beuQvhFv2Vleh
kuxo/KBImqLRe01vergX9zTIkoncY70SmFbhWGix2554/3h+rEebGaKnd+ZEu4eV
5Op7L39IrwgpPVMmmdk2CR2IBLnbtO5BPFbPvgN4Z61D1qPPr4tvhaoqm8LGi7Bn
`protect END_PROTECTED
