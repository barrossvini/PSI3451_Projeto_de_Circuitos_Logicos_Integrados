`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GiVnjM2WK2Dq/IAmdl8cRRhwSxabxaH/Z+7apl67dhhK9Lk5zBPgvR8Nn1sYgByT
eMgYDZfETK27kfd2+/Okja5xYRSLXd9w7P8y6oaHJ1z8/dsD/U6gVg4abjCcMWx5
8yA7qfVKZj30m9PyIZBpQk29z5bft8r86frCkFbtYzd5zbILqpYT9WKcrCjc6+l8
5064x0bTUEVkSecAByF41v3AcDdaaBA/4vUKtRbH0BXJhSEgb9PQcTlKtXAgiVLn
Uuug81U3ua/cILc0bNEqhzdxO5HDP1t6f7+KEt8YUCp8RjGk90syf5vcPHZjdM3e
Lt1A7NzugiMgmQhL+mahwQ==
`protect END_PROTECTED
