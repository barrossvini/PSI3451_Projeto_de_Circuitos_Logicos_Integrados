`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AhOLunBZiWl0CG1k/isQpMF2o/gTujCHz3QHiZV1/h0A9pBDCv2wMmP0r8MoeM6O
9uWQsmfUbbM/2fPDaQ6Ly5+JnW1em+bpUaJD4KR+nBvV1Wr9e8ZkFk+sCkLAaIA/
fkRjclCmnEgx2RgVJrs/O6WtW17vpJP4ET7obVV2chhC1qagp/SXi9vgIX9H9W0p
+adxwIQ0kH7Qif5HUF7qcvOINmhDHId+DqIKXM3Ft/6yZQrCYvFQNmRGxHNgHoYB
zPtofNDbgslT7GrVgsc8d31Dpke31SSSLbZDejDVCIPgdtFCIjsjXcpIvdzcdg4a
lOM6f37oMSqUBBFYAjAOZfOUc0SA06sqI0QVCSjfKqeW+GcTfzjHaUOyssKh+TXW
laB68NsDKJhvfeFCCqPBY93L4MbgmJDk/+hv+318h2s3AGH67wmar6CsgPEs7ueq
WmDc42ZE0iROUdepxDzG4w==
`protect END_PROTECTED
