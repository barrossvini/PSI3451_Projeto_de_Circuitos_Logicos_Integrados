`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9vSYCKTds1c/3eq2Ovvf81G0iuzVS1mHPrIanGc/p3AtzbQJ+3+GTVpIgAifrurE
0HKEQ+1f6jDN3rdgETzOx4YgEQw4lUFhh/o7IeszyryYtXlqfUewg39eBRJPePhB
mGTJ3SK2Jsc0hrtgVaCbjq15QRRmPAk4I0XbsJQN+nGm7FbZ9XSmUSaoGOmYdvE9
hZ29CwxMKpP+qDsY5vv5JeLaK9wvNS+xxboDpX8c7qCLUleP3mId86V8whsiQQo+
D/jx6bRSmd3Je/96oNAz24efvE1e2cRHFNH/A7uKktGu6O5DmkhUtxeaU/nzQwQv
B0Q295NnU4r1c4WxhoI8ukGVTz6fr61avgbpApfzLc8FxuH22wLelGnfFHYsZ7gR
aYcq4pFjo6pbuP/7Sr9+Lz2oogOhHXdljShW1qMVNAncyvcqzjkuIHcv3/YMdQmP
8sE0/FOGNgFgQ1SFA8MIY0/KpgkgFoJeADBGdq1HovAkiIqCJQ0Uid6vyAsGhlo2
cXtte86MlApCw57ryTmuQAN6DO8tuZ/oOnAj7a8KAWjPAmKvJ0BVLyxunj+K3d6d
q7oSOzFDFU9d6ex5mY+flF8d02o6ObX9JqkDhQTdp8i85Gy4YOxHU+7syrUbAyGJ
UpA7faWPEz1P601eCHTcjqdesjeHT+t4I+tQzkP1kRyZfY4AWApce9nRJPcN/P5W
EHFDXd0dcrpJQuFukplfhr55yTf7UGc0nP2hSuBXWxuatyeveBpoa9r2YXHT7hNk
MqzkiLhACrvIbMB2N2Hp/EaNqG3nQtE2nv2JR8SOmycX7Z6gM3OVMMIfLoWG6w8n
UGM5Psxr2uTa7+niWxSc+7/5CAb58PcWy5kQ1S1xk65T9kh+THVlm3dik2OkwAmT
5IWkEE6epsWAPROOIA8LDQ==
`protect END_PROTECTED
