`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VCvLP28F1FUiPbm9zfEuxC6jxjRE0eTUn6PXkCUqFI8TXhhrW9BUnMkZu4xTOv2b
EBoSjqKqRwBK/NEIebkRxSqzrHb2ub2EBRt6vyYGpuxBDgF1HRfxO+GCGiqzjbZt
Hsmw6Chkx26lkLRUiQGLN74C3vqngnLZY6I2NYDKATl+tAz9ZhKr7imxpEECqtOu
7JSjvgYMcylqNqjeBwm9pISDZFHC0fR3CuWIfwu60vDUBaBzvUMzzPjOWJoI1Rtf
7piUFCzPZpVGE+vbfqmfruzbR6RUFG8whgs2aAoZ9S3fTZELvnzoKkOlDEAWr8sc
v5yPw3N/nk7AO6tt3oZg5FtV4maUIP8SWuapvNgBgI5jYf7OFVp+uTDXoWhknff5
ohyQyctI7m+SpC0ZAD3+NrmGRdHxnlflLx/X76ZbLHTyC0NQuCo3/xWSZmXPbIwm
h/jSG5w8yUc8i0N7YG9fmqrNLeCcoGM1fuKhuUXY+GO7tLk5CO6eabtw+jAsauG0
Uim22GJtC2hUiJChaT8q1SQewDnuSdRaLJJJSIfBTMh9Q9j3Z0vhJz618GcKmnAd
omY4WfTU624AtMt04jsK6+6BOvgdh7BHxaZZhXV+XOBxseXmAovuDgwRpyOT4i1+
zRLqxH6B3XIf5nAKKoeBek/f7kVu8ZlzYXbIH0153EQKRTy8xFu1Ze+VX7Z/PwDq
sYAwBBeffFu769BPMM66cKdBpkcKfxCRPmfqTulY7arPnpdcLwvPKUFruxTUNK51
gXQoHz/RvlFYLS7UH0vEzaujvOw6o0wcbXTg4JgXsVRz/Cu7JiOmD/KqHbcdxYc4
zriAFBqGhgxDhYshWM0JCQ==
`protect END_PROTECTED
