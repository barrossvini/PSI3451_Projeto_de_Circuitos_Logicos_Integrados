`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mdJiNI2/eL8uBgSSO8szlZ3gfKt/hpLRS5ZDR6oqt0Tfzky3hayH5rc+icI8VioB
Ijg/cznUbU2uOpTv+6AW77J37gz0afMXKI/DUKsPcAAf0MqUr6mx8ko1RfxF2S5V
otPs4xAcvxAXlQlaPvYChYwKInlDZtYz/0805giQ1C2wN9DxIYIMBytApDqg2ziT
caCUK65sQGLxCRYkHGaNOhF0CIp814RCh8B25jowfVp/IvV96pqfh59IkA1vI/Fo
C6f9EQRJmHl5f/rXUbd5C8z9gb2HNmlmSCrDdnAnVbPjLy+bCQDkQOIsNjLjMkyd
U9saDNMOUu/4uyfEPuG0R7lZj+RJVtOcJCJvhNO59rMjSWThYiSqCgeMnkomBTOD
NFxSfouka0xtHfozj4CPYgEu86rgSq+49jt9kO0wkw08tF8iv2SstYQnIGEWlzC1
g+xS2loPWDIUGeg0DO2o0rAEs9DzH3CvN2xKxld6D6Gt74Fo3ZE4QVGIzrqyllEw
MzRyLq1H7S4QOK+Y6QNi/U1w23EUKDsoEHz6gk+UJeOby7xORfYlJwQvid13b7B/
H+Dj7vEN5rdlJoodQHNEspKAzfBg3ClWiOoMg+GvBqrZn5jUfkvAIWDsRb+AOpVu
DQwFVvBEHoE8ff8hTHpZtPFDXsbpTnnFhvk4CFHg2sL5DrA7NJO00j+0sm8JHBpJ
q1oHa1eZZ7Iki+a0K611DGz8E2P0BR+HSpwUtmgTweS6xUXbGgBp96hJ9kjFOHFP
qTuSdiTVYjVSGNEr02zkWNXDNUpNfgIA//a7LLi6apFfSJlUd9AnfiTqjH40cckn
4bt2xpwQ9ALOlHGp6WVVXIAOzL/f73/DZmerYZEavTKfXReEHbK3zlEGHYISUnn3
s2o9GULYDhbUJAgbdHZDxeabuGf9AXYfDeefABJ22rX3+OTtom3FNCtGJeC/r64R
sw4RDgtmXBjxQoAWxFYvbCNgIx7nvHx2ShmJM9Kj4t+jZ6yYx+U3Q2Jz+w0sY4v6
GM9uu9ZNU4XNjK10Is9Xm1CJpv8rp3ish+4B8Kc8cvfpYrbAlQzQ7NhtET0U/cg7
r7/WEH3xD5e6zJGEmOyYoZQNxKgKFAc7ojNSuYxgX00edYMaHjuEhJH6VLggj0cG
YNCsP1M2nuJR9KpjndiglJL3BzWFvhrEYJenokEs7zpAcusxOokPm7EZNnZM2igc
YtQBgFJx1qIE25ubNDf5V4DfJ8ldxlNuDFJyJX+dNnchOFeW+fSmQCzK8mcA6uBj
Hy2j/qeGfB53BBP6GnMoEgB/VjR8AgKzZ7oPdvgin/8D07heuaPVh4ydICsGBnHO
YlETWsKUcjBhNVyqHFc+Qo/Hg7eeMoxU6QAXrNJHGf9VRPp5O90HUiJ4PUIfUM+4
t0c4n7c+LC7JU54AB8HYbpfR2C+PwEELcHj3uXTeD0Biw8/F6+tvOxQEedC3Zmp9
xbGGpPFV2UIAsAV3K3mRyXkxJuaxYh9X0AuXlpZji+qeZFhtcLqi3wS4PyuxksCy
0kovDngv63guslY//LZ/gJ5qoFi4py0BKnfoy74Aq040raWk8RAS+OlSWT1hw5FN
mJK3NinIWyBTaqmgtR4UTXtuReNaIfBR20tSuF+wP82FqjZ85xFIn9jEObi19vdu
drd/zqpr9/jIhKjVuVvb0US1wdqvJLUwdhXHep9fHpM3+chUDOTwDiSJ2NAve3/4
7wmwuoLnpTF7e1fqiPhEmK+R0zeD+yp4ru7poB8Kn/wWLaYOukHnmBYqVFK0dSgX
awEKaLV3qeUUfwfIzTONv7Kfqy6mk4nBiSNUeNAfgDKxEeucf2VFo7s+vlV3pbmb
hZAIuiqxJjS2W2bvRzZkIEgkiy/RoP/kYhSDDQk6VZwO/1TmP6L3piLnrwfrJSFf
q5meqpkRPdSicnwzjXmyQMrdS0MdujmRRazFmxRp2lQXl+ruPaakNJB7UumY7+53
HMfXd3HXjmWi+ZZ1dmVe/RGdBGmdIjpoh7Oi2PbYJKYgJcHFuIV0TBxUFOK+CEXd
3J2zdTA7QlwW5J1GT77EN9vdpQ6rJe7mENs3o8wz9gzQH/5NiPrm99TGCNZUqXky
WYJ85kX9aQ/VwpFJesuqptw6O4J0tUoZaCc+A1o8kbb6UzDIexwQLaGLF/mTwg47
KwnSnOXmSighBw+c810dava26SbLQX3lWCFnFObKZjri5eoZeib5n1L2tdcncscj
wL5AzawGvnEG/3jy7lRjxyB586EDrsWzQCz9hrZmohHGB9MJYsQ4VloXEXG8BRtg
K52hxeq8YZVGaXZNN5NTb5tW9sAmDdMiEGSNkPwx/5a5f60Xyc6uHlb3E2NFegIZ
FLrAuII4uL2NvDGSMdBrAiFGxyg/iaqp9UTD3fAuR8VDZpyY1BpqDVNA/5bVhiqo
UQ9VX6In4YoIEl5U/vwINuK6hypcPgEWmIPXFqhxqjoM+dfvBBxigqAGOoeuqK2J
V7gvlz9RLD8nb48P3qjdAA6KTaksiXY7ZgohfkZivyXpsTcxDqd5FTg1V8LTaepy
u92kXTZLNnfQF8/jggoRIUa5LNVAfoNzzAtsppwVq2nFgLxUmi7qir6JnmDS1Uii
RS9Gt7iEtv1/yhsej8FgzsqQToY0uUzYkm311PO6g4VRUwyv63eaFGIuVp4JmcP4
MHi963zOE8EFeAehYGI2ZRR4mmqpCNyO7w1yvPxeoubKC46/qQ0DGSmVoRoyQLVj
xUpgu2WPAvA767nElfXBSas2iT2cS38DWp78sJq/qf/zNerC1ZQSQsMRXK+BztoR
mL+v6kuRqlIfu0qg6G3avj/QLxZBvuaSpR++7yc4Z9OV+QM7KRU/JUVJhB/B7HBF
FE35RQiTToYPDKEj0fr+8uZhPQRO8tPzttI/Scl+eNW7/xOS5++bQV/dsKZ3miI6
xpGcU/oo9p5mwW/xGKbbWk2hS2QqECf0AI23qcKMTuqriNONZvAswHqbt68TkHJE
r2qL74mcVvC8wkztplMvvHvhs3gwrwuQG1ZT05/rzuuCJwRJY5UhlPnEzoR1isfJ
KnB8mdu3cUI2FWQymy3dD3hNLUalQXk0Me2rvLST9J/CFYm20WIKI3x1I1Z1zacx
LrCV/vRIm1x9EilCXyW4GhMSMFU5N3iSN8f/sWAzzEeTBWlMwV6GVLNTcfBm9ACN
P2Vnb7dwL1Sjpj3Ywj6k8lGYl3jacm4CFPi4Be7in8SOek1pXtnM+YoYz8EuNEJ6
Q4m6SiNeJ1KCO2YyZW0NDjCl+zFkgbqQVo8TyJIsgybksfkouNVRUB/e1TyJVuoZ
GcdceE8kd04XytP7gWjzEQ67Dmb99+dZZulFiCkOt5mgJwLehGx/xneJeivsVSKq
m1Aa2wqSzheX007TFVatH9PjPSLt7MfUwKdZ4GCu7vy4NSdGddl5zFoPLqQiG6MV
VrqxzfFvhNBsU4pXhpC1VdRRjrzCEJ3QzHFyH6ERXZtd1VKKOb9ZDYdKQtx1el1F
gU11U5s/1nFZIF58tkRQqRbfL2No3pqrFV+uMvKNBtrCwaUYf1tRhwQ77c4tkQAp
r34YmkJJkcduKvW7E/RVRrmlkgMGcgwMq/GdBbQ8N+SmtvenRmxLtwB870vl677K
sDW7y4cHnrCoQv6gW0I97xRpgC7L5u95jJTnwGZ/0ezEUrWXfH2LGvmEwbuLFwvT
AxgSEFXXcdKAf5Wl9Luyfhl33LfiSiN04arwehZPjmtCd70Bppl5kAmN0la9pI7m
MQTrM540HtnVRvfkAnx6PuwVeI/Pfgk68WNnZosUSnCMnJnJcxvY/nQiOQMJUwuL
VIEBdX8TUi02L1yOTzNRI/KZkyFijvycJVnzbL7OxcdwueBmZjTU8iAVXtHS33r/
20uB1GdTR4rKk/l4u1RrpOFFuijFi54R3HtxwyC26+Yxc+Wle6OhgxfEhBb5FCn4
7gdlHXgp1ehiuP7DtDcGC2NkPeD4GDgdiJ5NYY19iI32dycp5v3CvQ1a7oMo8EAG
EE1WD784XKZzItccFT3RB5yRY4ow3/0G4PdWtjQpgaRbJrzdorMAGsak+SiRqmcu
eAb6nblHOwiB9xeJS6R8l676oVGw2+HrvHoyiEus0WBUC4hKrhT/NTDf5iepPBY3
QJX3jRxfgUNN/e0MGNUGXa2rFmiwMMTBNqECGSCk7x39etsbk4cOsalJrI4gOys4
pcrc5otIbhXb4l50qxrngAZafbuZIBzmTpPF8AmrKm5jUofdM5XyaI45vHTiGRiM
WfGHggzNuSSGDHUcFuVzewDq3ACUecngMYvrAcs/L5XfiOQqts4PlbgOIL9Pa4hx
r7ETaPeKoT6xImYa+5l36aSvyKtuuyEZItHfRSAvJLeYmw3d+Kiw6F/OlpD+8M7H
s8vUAJwmAd/MctStAxJHoSb1SY1y8GoRP3xdciC5qPZSMz8jEdOf4gE8R8en6a88
5Nz+jpIWx62bMJFKV1xGwLhwYMz20l0dmVNAjgc+aAaKJULpZp/7HJ9QrO8nwWyw
NihKFlAAbRCW3WjyOA3GopxeQzLen17q7rP8LzpdwOmGmp6jfuwBn5EXNaPFNGCU
nPCgZ9WPj7Wg5xWhNYZIjKsu7oyZcaeOrp/nV8CvzisV6NwscgvXHXtNBJ94PiKM
4z7oSsP1jxVbaH+DFNi8BxdgF5mEmnyvocHcvJViTO5jx4Libv197WhVvcRzAQWW
l1rDcuZDrEkeGrq49T86hQXU8Gofzj7StauopKUCJ5w60/hRJ+r7V6A7os8t4oWm
B4N+QGOBDeUn3MaslRmoraxYK99d6kxPTQ4/XiM4xEVlGKeouq2Cpdca6wNDB1a4
bk9WlFnShwAo2S2g2rVn395I1oDqIC872A6IEnRG5AIkqAze+/thZWgfNB0jCijx
AKX3yM2vn19bO4UCCm13zKEvLGjbWwuX59/NpqgVqV+f60Q21MWWvHYHlhOStVJi
qrqnM26TmqBPmMdKWumAApdUakNflL0ezNMiikJPsmg5jiZct9owc2T2cXg56aDr
VHcW2GfXP2fhgq/eml9qpUL+JlVFdHb0RMRnXQIfE/lSiQFxowiDkj1kqX9EBG4x
58R5/3jPwKoBat9jZnq0wDKLvABgklRN7wBs10icWsUZ5JMp21Ja5Xh066gZjk/s
bXVRLBmAvh4MsiFw1eUhLLCG9/kk/tRe4AZIm2S93kRTGiAfHUEgV3oIZt2AMXW5
PS20oW9fGLYdiKIPfMW0LIeGKZSwl7VKCvqbHFkIxkNUPGsmJbaFCy5UrqFpxIYl
7QEvzDoUgvxqe0g5bPhQUX4I/g8ORd6p+jXv6wm1mhoIxQrPSCXbW3d7y07g7BLz
W2aAznjA7cd2MdKXRNhwCVgT/RSC09aL8Ae+86D2x/RTbDDEoRlVg1AvyFONaIa8
qNp599fEsgdlBSChJaEM9zhUuOgp3o+2wU7gzyC9aM3A1ome7ARxtLJ539fhJaGq
e+M4XVoDnl+1ZivRUor/KzOdNt8tAOmQ6nbQT0K5pCdfQOxUsSqQcrn928hPcoor
xYSN/8Zcj9xrJ5odwwKHdvh4Q21p2RLpOLIzzxA/nzObzHYCKHaeeOJbxbkhd4WF
p2Fx6wPEwdWMjnvL3e71JgSq3epAD+ggxkQbrpuxg7XxRTY0RVdeH+blhI2PQ36i
iXTf1DKFSBL6WzrS2sDdtmQNfeb8DQVojJSw9CFTZiac4R/bdTAArmI8VSTezM93
HsTodSpj1npjViPM3l/xdWi7MDUcb1RG+jppRhaW2fiAr7/qEDCHITpvBzwR4TwN
e+CvVpY6qq+FRG9ZnKqEtVemAfa2PJu7zZt1Z7JuINiSDaSYyQ4ulutHudHoXfmN
JcgoO5w+TuI4ocKLMSdS/7cG1rOBtNss1OfWWS7eRreLdlm3TgDxKC6bNID+8p3v
pVm/Z3hS786ZEOSdtsniAt8OUln3X7mMp6teDJLBAKHj3dHYcRIxSscCCh7Dn+WE
zSJ1pkrS95AGEL5dSRRCyoUiciClYiSBqbxGr6cxots+x0wMKKU6q6PU5vJdBci7
ZKxGzt8I+aSqci30aqTPSvYF2GBYpgIjMi9Ckn40hgKBnWij2/wgtTyAC+CwzrxD
GctmRraqY9WybR4T5oaFqWgzbET1l8Hlt+QrlazBisPxYA31+fD/KXM+hGi67JjR
w7h/YdIiCW71TIDlxfAw9/07G5INCrWLL26HeCWyDF3qDGg2DpLXOpG+euvpffs9
iioWzGjkaQSC+4Zn/HAh1kth/S/CZOl1y+7IzknZ0w+JAZCk+9P2kEobZ1sMNFut
7PytADl4KzERP5r1d/O8k6cPoMcGnE/HU5ZBqHngb20JDBPPvM/BDuux+FiGOo3T
Rkbm9V3wvzX6EbNyPhgMOVViLfCQvn8/YdRrKtnlRIQy0hCbqYxPRcKmOlchEpvj
MLJ0lnkEyGPNw42snohmYeBGUQAAq4EW5ATWlP9PHrMd7k+nmuJIRvDsIy0SzvLs
VLD4G24dp/oNa58sXNdBWJQWHYAb7Qd5Uyys+cPNM7mNW03yiD6z1UNJtHEHOs68
fLPLf3XHlcZDUM/5jRyVVfCWK5KFp31g7QfW2ci4xFb/APDq4IYteo+T6oaCl2IS
AvT67mhYdLviBbGXmUNK5BfXO7TFeV+p5Q7uRysCHt6Dg3qk9zyFFOaUL47Jh495
79/8Ywpwk2JRGvFJvHlQWEPVnTmkMIzfKaPIzgvl3Uh48Mu9+SXJmrdaHE86BnYc
DU5nXiwcOahmDvmdiXPX0Qc5mQUYhLEnXzCkqU+z470QG8V1qGAY5rfV1daP/5Ho
0F/xFeCAsTYTdOV7r/Zq58Wn35D7lN0vAeZ+EXxoq9+CvR6sWmMlbfKPIdQXAJwP
tdkb3P93/bpj6bGtdcIGu5GqnfgD41riYxvnv7g0DGt31pdFxn08IOtKieZmYxfA
fv0IOEwiEK9PCmW/TV4zeDkKUULq99rKx4r+na/unjRh6F0k9vhfZShLj7RP2tpR
/T7I+PhG51lySmzNPEtfnZU2suNuH7rNRLQW35lBsPbWW9Y37ITmn3EnDmGru0aB
dw5DX33Vw3xK1rEFfMkdSoxKqqdTYLT2Q7s6whdpYv6unFnQWzSqwNzQirsI6BN2
uU3cL+lcmDhxA8/8z9cAGIjdryJR7OyyoelbXh7Nqu50BahrnL7lR/BusVrTUSUh
xnaLIxw/utl74VVWJITB82bA27w7DrmkUZkl+N78FzKFNWQsVO6c4iVFPSoReXBB
ur01ElyF87D+j1Gb9q3LnIWQ1Ps+itdwxsV0V6GDLLj5WKG2860yXYeXBoxHRlFz
K9FBYwKZImhk2KDOSTwU5yJ1uf99oXPMU5em53cvPXOKS7UficiE1o4qUonhboxK
H2LLadjWbc5cK7O4IxmTiHzLc0ihnHwcf8Nx6x//OGhzIZj5gFQdg8atDqnYWzpa
hOkVBwHmMAZnIzSsCfLrYzUW/V7a5ci70x+Au120jmoVj2VWepdwHT0R7Way5sLZ
bAvBCyP5zszhPIEnqYx3PLQ76gxyJ5GHJrPfB78prmVN/ui/eiyNbmuMPAw1QSr1
x+Vbq/aJHB0PMa/XqGlPDlGPf0ftDOCQTCxFKSWdeCiiRsqDbWXddCrS9Xp6RGso
LPaVVTlWvLlJ0Bg0+74YVxAwTn7NFzp/xTKq/gGh/OyjvW/+wrO43Q6F/rFDSJii
KnUqrjdBcG3nb3+83DgAuFFbkcwyXCsrYXn3wwuWcZipaT/Awje+cEZRnuPqIJia
hZRgbrDRi4HIeAp9AK/im3ukwH5YnkYh91zzY9NHYmlU1egtWeS8I9jc8B4/8VZ4
PehptABGWIlxORgrDa7m9SBGRlNCyovJnzrE2cJ5JiSnXgE68k39C4K3NftpxKZx
sX9ok1h5ZAD/E4sgUMSqDLIFXzp/EeSkzCpCc7aRTAv5n/YUzbqpPDJHPy5phzJ7
nAbvwTA8BRYL03nFMtsiq2t5VJoeNpCzlTV4TwqTePeO1YV0vieS60TjmD8pupy6
TZvRpvnG/zXm3IlHFmmNdPC1AAv56doMc4aKxgRO65ykgGfAbXAMgk0pHxfsMEjf
KsBIxE6LacCtAC7FW1hgbPM6Nh7hA2HERKJOjYZYlRKXyf2SwOW2nsVQ31d8CUZB
zS+TJ6nEpU9mg4pMniqUNdND3A0hOzZlShXYfuQMwU1RYafolsZ0epzbo3ZLwsey
G//upeWO3tAMVGEAhER40vXl0Gs6Z34IhTu3fBqQmL3govYbnyVQvjp8TbabeJFW
nZ0ht8WD5AF/ix6RNkySA4y8LgDPIGFMrRVdIJmWLFJ+/x5EnFvIZCf9HBfBaU4b
DaOy2/jRRklIXwtsqSU/IrP7YJR6WEh9TH7VZkE3R0dxKo1SGN28irDrbwrRlGWC
5PA0spHo2dpn0TJR5/cv0YDlURKQTTUeWz96X6EjNyBlnd6Fyq/W6ktg5wBCcqD7
+yCJeOMJr1vom+OUYX3zyHF+h3AdRTJzNi+56xP+WP9VUqjQGtdN+D0dGoqB71qS
h/3telfjvcwlFA9hCkXufKWiu/lIkGd4+q3da8spKV8TYZM4ArgavQOcHdl5Nfvp
u5CIwBvUrRLOtpNTd/DaS6+hY7p24iz+EdVRsZL7oIySRbSCjud+nhJOvmQQNWGM
isyp/g9RJp/V3CUH0UkU5Gg8OG6feuQpFuYOGoTHJsiF+nW8Dc3apHJAlMqRxXec
YihcqsNgA1+HZuXAU9Gf1X5AV82C5MA5jhkEAekdOd7iE1vPwhwMOSIriklJO+PT
dwqvNMgP8ftt7+oF+eygSq/a/R+ZYviSTC3MWKwGQ5qupUJeCrX4Ptj5Kd6AeKwl
WhcJqm19j4fzgHjgaq2DJ8L/wXxM1PkdGu7dFIW2lNsctbtcaJF7fISW2i9yMrpV
8Z5p9lGT2FDPUFZN6wFkRID/V8QEVhR2lJt1UOBWCKSIR1H/s5wfe5gko+IWD+dQ
V/+kOhyF1IQzbIGL0SMW52z4CeyULBg/lm6F8hnmAS+Xu8BB+BdEhyCV0Ca+/dKp
1ezZnKAYVNwl/QJgS3U970NpgS4LQxeDyLLN+aIoAcFZwAaPKrdMT1s7Lu1zmkbS
t8T7dw8iq0FUALjKJFJ9ZppCeMsTr59qHqXBcOAf+n60PO6zPWcoPN68v4o172ML
8hrQ1DkJyXM6HxDLi3GXOw7F7iBmJW+yx7M8sVBop+nUJB11AMa4BuPxsqjGILpe
h4476dt325sL5j/0BC3Ls6qxCk3FcQuPO9STSMELZvSzHzV3H3jbIOKaSqgqmplc
Ck7tn4jdrdrO3/bPfOoSPN5Zb2vqrEUnNRYAq59gm6dgQVFaNQxTW35lc3jwUQIk
2Pqh/cxH45CQqaHQMafh1ielSi/8VDvSI4S9SZS+Oo9iv/JXavwAdcf6uWwFGJPp
H+jfOs56If4lDYGp4wijB9XrVT7pIiZYxdb3gEtY0NVv7i+wnYZAEpdUGlVdjeAj
zYph0DZ9qgsSN3aTfGsfVhN23qfyJ+SDw5Nx5NfH4PXS1iFoFoFOPV+aylEfrEEr
3h4T4JUd5CYXbLBq5uiCCaCDQXDyJqrjyTNd0nnM9prFBjsC3Rkj4f40KO9jDHlc
UJQlPTRGc7Twky7iPF2ts/hvfyaBUQS6Jgoe3U55iELgBJbp1ovzknvGxJQ6CPWV
iJzcxbTG/fXvqB7TxRVEIktG5z3LnMyuKf4gW1GcsWEgqbP5XiysMZM8+q9GrUJb
IkboJJwdlgNxVgWcKKrft4XdcwDsSQmX4pfFpUS4slaZ5i5nZNitZHvespGtHMXq
yPb4mvJXx34SLZQhKLzLRfpGBDk5hLijm0w5qdlYkNZNHunuqUNXYNWw4yB7ZsHv
0hyJnwtdw/PyQAioDZP/xhxC8tmqI2vLuO1Wu5CLK47pcpGzBfLo7seSiffI6APj
8Jf6n6vN0XJrby9v9lkRuEVfY7uXwqxJsMb/4ODRP/YrPt2chFN0Aj4HAxsYa2W2
Fgl+mQaDfcBm3odYxYyJF8edSzOu1pmpxHcDCWLxzG6R353ZZlW/du1T86ntU6JZ
Wdc2yBnNqIPX3HRC4568NwCBevO2LgiFidLuzA8sfekv2OvGMh22lE8NodHQxrZ+
yzmky74GiAJSaNz/eSs2WGF+s/PnEPjm2GeRYKhkD4YkGcrzTghXe/3aTnlf3xbB
mHfDzIO9bIGjLsyPgcWNUlt3B22lpyFzfr7pIc40wS3is+lpdAYc2yYy3QDa5mLF
0Y9Ovq5nVEl0oWSg/GjapEDAah4p9rAXSkXYC+bFr8PwWrATPxLfPCBxv/WQfzGk
FIazj6BL+3xZr4C8qX24vymyfP3vM5+2RDR99fOa54nFxUAnoMrRw4BCt6tTphvc
FJgJEswxAm3hcuQlcpTtQeW3TuLIBKURV+rZxv+7BPjZUNBwv6Hr+CqFluYnhT9E
MFVMpw87zL+Rf3lhZHjKGGgiqRCLo0BEHDXrv1kjZ+HXGBSrqVQR+4165XdcMe3v
mCvV4+mn0TJqHXYfJvnqJTTUJFHLvTXLmiCDwtcpLGIGzf2RxVmQG3SZeOHbjS9t
+WtpCYtYITNMLqP/W7SGAB8LWYNgrhpIr8Fj2FC91dfXarM8MQJKOrn1BsuIroL/
DBybVCWoBG6c0sBBg90jXrxsxp/fEZlTpKoS80E7dBv3pv6speFTlXRbwuxh+HvU
dKFltEQ9kVbpb6LoYmf0wuKn17LRbkU0KcNYWk6ArFkX7XuhJPPA+n0H5n6XA5gs
4AyE4Zlf6cbfwl/sTzOrzHOU8eUeLMvQ/sdKobc15ca+AxDVvjp7u7R/ujYyl4QY
/hila/KnsSIraf8O2Jm47KLdiIXKPp5k5giSkQzNbDYrdmQTLsXfCjUUqIK4biN0
1zyLbmm3ZzY0TvSI0Zg/VFRaJxKgXcilK+LxmZ0+kM+G9daFfbtnahWwTfqmK9wJ
8v3oKHt+G3K6XI1ebj4vije194loHPOgTq8sDN93iQSnvCmM7CaAlMLFVoTQeL/Q
Y9L6L9EvzC8LnPjMrK3NpBckhM4S2JmeSyrQPxrh5aUtMQnOPy/wtS2JJPyHW6pW
GxrbGWQllnd3sHCD4FXb2yZKalpaJHYMgwPumH69YYocisScbccAgScqNLvvswaS
OcGvOsPTxZouDt5En6TzhMJQJxwpNuJFfiaNUregePzFLKX5+FdRjLLthbqhNyV/
dVyHI+GfmSsJYWrNdx/GQ4lvqna4BCZTZR7kp0KBw0rfxpeeVzipCH+/hT8s5Pn1
5oqRym9QS7L9fG25Boqj670N9mxpErFIksi+UC3QGCQdkzWKaOmLKkPEbGnr2xuG
agjNSWRdw58ta871QsxQaVW4e+p9bNqrH47OtJlTQzvWtc8YJsbZMYHX56pXURby
EkqTFV6RXB4wRKSpoYLewEYzzQpupWw4Fx35rUATfnfzYoQPsvor5ndfrRiXeYp/
K8Fe47+W8pdRkoAQMFLXVdloHsYCvHmLJiLERaUtB/iZKDl/bfkfQ9XAerogS6ao
DxiB/+o64eqkIdcg0UADXuc0MOpeQc9ziU4zSIZpTPWSzoZ3nSSf3y9FzA4y+jWM
6v6dZM9WO3ut/82lhOAd2hegMZnmTf08Zxf7dsMnydNE2PIJg7qjffyPdHp4qoy0
IzPSvPVBDDZy/v73B44SJzboiUoi5p6yjsDCrPF/SO7y2pt0GvHLLnm1H/MHJtcg
7KrM7rYuCyIygrhS3aez7jai+wYE251JHakE0Uu6hyhPOy0Md0Gr2fEgptE61nS2
GBXbyiWd1MGz8dOw5i3oJTVd0neWcKqhr/oYzeeSV2Acj/N7lahDnG79y3utIgDf
W87613FqeSzJ/73PMfqZeRtPV8gO6jZ4s1jIFwEh2dyOOi3H4HDxUUjdOXBo6JLp
V9Q6bq1QKMa/pzqMs74hOYEdqzaUmN/H4pN6uwhJQP/2iJ2mnZCQXjfsLtWNExic
Fb4fa7YsNUEKvo95QbEZD0gzza8o3Vl3WUs/gPQw2rO8c9Hta6FvY77bbBlMonrh
rmsOY+qzpjeEP+R6RiUJp1I2px29VwcR8dt8xczAgw/vwtrs/rGqVr6ogUcDdqgH
XD7GzIOHn2yoxCLkIgDg0SNG1JBl+i8Z3sDERcIODtvdEnLL2wDSXTwEp3gI13fP
OH3KorcBz5jx66ypcbNdPM0gMbHolhmo2tsL8VDr8ubdQbSOJlfdbMsnF+Hvccqa
IvPo8Qn7aiPZ569Qb+zMQb89FVy++XDW4hE1hyBSGWsleQEXMuTDePgH64bcr3hB
KwoBG7GgZpjyo2VXjVOTRa6rsyWZGLgmIkNEeEFipbhCw1pDnVKwdGtgr2MHGDpe
Ri2jyk89UbXepAAsDjzhah1qkx1LTlB45y7TmhyvKeFgRSYpH0XfZUCKWQDZ64D3
6DOA+UM/qJXbdTj6RuXj8PB8aWsdpvPrIl+GJMfm57u557syUaJGQT4XYgpOJJSu
aHyjHkwrmT2Z5MDNTng6lmCDXK5oEIwtplmIBGi1+QagT4dypn3J1KbR0Pv7QhKK
laExOMjfHXn1qLftkBB9XI2fQYHvmoaawVpAFfoeJpIODuLnsSxOMCkx5y/rZztT
iJ8UA8q09Zv4GHxWarQl2cFk2nvpUWUWuZrDsXFePTbhb1OuZi6gLqSeKoHfWaUL
QmOU9zYD0C3g7HpiLXHSlQAYoodc1t8CmczNie10ixOjOy9O1V6Y7dihi4anKYX+
GVj5YWXrYW65q2MZFM+xPcqMCoEm9W0Wr57+GDU5+LtJ5aJG2AMWipNtQr32C0OB
KAy9Lfi8x8QtdCdqyK3Y5mEj4QQdZvmv75yY4m88OgPXxIa29FbqYrJ3Zc22Z2lk
SY10MOe6EV1l3vsKnECfhqWGzBmmFuRU6H9LGJAhaqK9Pi0W95e93E/VPiE89nka
w64q6GUs0kbi6xACMt6IdV6f3+qAHDIzxD/HSO/zvlbiXqbPIb/3b91vr6sFBFNo
xTUYB4k7QhzsLiAaqjP9nUWV7xjSUIyglKnsqr1og095LJ9B3TBcaQdDrKZBs004
8vQBWz1GziF8jN4YdImh8eHyt4yHft+o2jf8kzVE5hzfqs1rfOm7TBNVgEbpBolw
jQzniuo++bYu2ESGA4fXo2bXklrrXhwy9OUosSv2I3o2iZvsxi0e5J9ykHb+FBc0
PgvjgcqheoQG+QrUf/gMlq1pr9580pqAufNHD9OCZEW7By7p4HgCYF6boOmUge54
M/tllZAcAAX35jIBiAIFlR4h7NtC/XO6IW8YHTeYt75sFiduMWfW5jPO7YR7cAdP
BXJZ7VIgMK+E0FaJ7KkQMaFARyxv6wYrOX1qXfEpiujrrDOptQ7mJ0Vy52Wc/iTq
U065NWpL4ySFqFk67ImiJnbATa3C/86fz3H4U2TQ89lRKozrAIH1svRkZHCedHDU
FBJcQOu02myXGtDG+1FCYmDBp/BZ5j2ZHaIl21KoJ6eqfAHLJPYJODFx6K8E89pU
IrW3DTB0qw8Lz4E0HIq9vsk2qibtr2Do16qOJipyCjLFbnhCNYcC1vhyPHVAUUqn
Hh7UKkqJekP3zJVL0i4UIXrf2+b8BxcsSoAftDXIx+A1pWhWvpQBkdbU+nfJGqJB
HMlOyrQ52Busn31Zr9MiCkLXwXddLOaCwnCT88uSoBmL9euiaxI/Ct2D+b6PYrhK
nEPFx6EVwcRojuaC46jSYyUpdnmsR1olHTJ1DAmiSty0AeakRRLOTy2Ad1ICuJQA
reb/g7qebGbNs1Spv17J92iKfVC0cNRHWf15lotB5DxdrEMV6T6PLv70A5kVeB2f
QJtVSCg5xv/eXsQgQVJ11nliFp9nU1Odc38PQSf+qo8ZnK5q6gHgepVgztkRjXbs
ERzmFp/0LnyJEseYLEuYUDFVlrFkQYO1U9s/sdKwN/UvpOQhGajBv98hEEB1OGbj
Jf7MqUWhhL1Dy4gTsBJOVbzhrrrqDo0yyD8t22YS+ICFEJpCZKIUb8qNnM/bVlAC
jebeAx1vHPf/LvX9TcIOqMBPJKA4EMPd9jRoUj4OXW8YjtnZxUxZRPmcd3N/Nj6G
ylkE6RUYtYSfLy7hhmWLh8aPe623jhl5r93wYjdrefln3Us1pvqhDU2cQr5yssf+
cOFVgbhrt32qFRRODedyVkkc+aP7BqVor37yPnIOeD/lNGRTuWnuXY3EQLRQTUBu
JWjEVvi/fYk9i2KDrEne1QtdA5tFE9l19ED69YhrTq/Ozbxak+Ou8ZF+fub+FMwd
k8fbv4gxZsigApJoYaAQNuLsC0IuyAjsUU+83PB90+ZdCKbzEX8Q8SFn/QaLPzQe
L/8rD7wRm8FQHmXrTltdiH2wjzyTPtFcGfaxglLV64tgKGBb1FOb4E3Z3i6HRDOg
CHkSKRAR/gCcWRBngQWJtyQtSv0oqfqeou63TKlGyQnR92SWjVt8Lf10aA968Gzj
5S26WvElLIPeanYj+3yasaKgnr6iQgwAL9lTyYW0u1GiH0yqHIT56PrzuCOhOxog
YYD6t0pj17zOylQaT2mYMrk83Wnprc4iJ/4viuH3Y+LVjXW04N4JEq9LMrM06sya
ln8VGgN9t5mcf0rWVBPdK856rgO+lKTQblIfbgKuXxMG0QkSNENAGMZ/so9nuDIg
vH/zDoYx71QvcjYd7qPtQIpJI25a2LVRfZg96BnwIStEIHoR5+yq1SUtQU8i8Ibo
a/6MgmG+/X7ttFY9vhggR7wRN52TsPxKfrY9ORCDxbN70jK0xQZDRxZb5cIPJ1sv
osn6BB7BfDFF6N2YXqXymsLHDxQgik9xoSUwUo4jeWNOO4GcHUenwF4v0mKZwTCa
PSkS1yBiTKRSbx19ate8ng1jHFLoS1rNQPUXhA0pT6TvwCBF3ktaWxT/zG0zjB+u
4vxUfeygIq/3y5M09w3pIxvOJcbwYej6RGTJZa7D6pD7AwzrKPP499Q6snb30/O2
KPVyvktp5X1+F/GiRXNXtI6rA26LSsRUYsi1Hk6FVFrMhcQQMe/5xsDHy4VdffQL
lYnA/itU4vs3LcTPMTGaQvhcDoVV5lAhxjcmkoDIkjeIu5VSslKIAEaXaCrr5Wna
ElJ3ktfFxJos7wYSXjceOxCjQCfJEG3wOEQd8mmCDvMQdB2sWFSqcRteiE/SHMLO
AuvmI8BpgdQ9hI5eZT7BcVtDClTu60Fb2WrlP71FiGc2++WBw8o1kmQQPUll+Qbv
RSpxxCQPNMT59PctEHi8UHSQ2QZsWPjxyuRXcGmJnkk970CvepDo0Izy9//SVfas
dUO3/30YjbuCAk+/b2bvygmd36p8uB2Ged77bdOk6Z4zSHCnu8PJOSVuGUx/x86Y
QLGEHyMJiDTjW/bpNaOgOPcyqUGGNLEkZCurlM4n+JsJQO6CVMT7K4fW9khTIylf
phsrCyxdyC/PiM0AvhEo6cXUHlv2YE1tzM8aCAivzKGyIytgbmtA6CYpr0yDbdXG
M54in3SUz0ToTuqLO7bvVL8S67nNHgKMoxPiPZAR8MWktPs7l/KbQLwUD176v677
Xak6dXzhHojful7YdgSvvZ8FeI0WgekP8IwgTwtpWl1lOm6kVse7nVJ0XTw0Gb7I
Xs/zy/OsFGDdaJhIv27VqPmZT1zEZV8HKtdu+N/ua7emn70vIVtmc687ezXFbpQK
IiGpIR7yfovX/Wpcjg60h8jrDQyNFCreJC1IDEOei/lmxQTsLdVf9XaV3WlOBzkL
NA/LCemWVeYiTziR6PjhkX2hGUIEzEuMsufAcbiaDssoSHHcxLzTH0V8a5zsxqYN
ihMQTHINtJ9VN0+LSAU5c92bCQjeMiJl4RHnsYQ64wRwTMtOJsGccHomtD4YV1s3
2CM3hT1IyO3oLGrpwPDMnSucyKxhNJtPbWbvA9HCPK5sTgviElYPf1u8EfHL6woe
QVQ81yovx16RYbDRlvVm+aTnD/o7SuRvJB0igN2o2CItWfVRifbOnxwgOm8SumwP
z5uy5d5XUr1L6OLG+gpmRo6xmacUwCevIT5GUvTAXuNgSERw6LNFFf0SHvJmN3DW
5h1rzcSrxl8pFmbpp539zZJOZvriBPEBiHSUjeQTENNNpSi19PBG31R6eDu4WW7m
9jNJZ4fIaLcFKm0P0r/6DHLyyUV2ihKBRFihannZ/0X4fyYXXakQ1uJvErbFFJEx
Qu1VimU48cyaXftxIFELIhV5fgpgfsBAh4thJif3M5o2SL8rUgcd3DyUkgwdCY6n
bdgTEf/syP53j7VcQI0Y/5SAHz40tiiUWd3r3/sLgozge7BgQ2KxKzR1/4+RGf+N
ztvVuyrTTMGPBgUwPxrZjRaB+d62bvfB1W/ZjLX7FnJQrK8fGTaESefj2Hf0O3kj
6Lbek0Hg3yS2fcTxIKHrTpXB8zLDULergJTCzET9urikGxQwm0dri4UcEhWep02l
wyYD1BCBSXH18sHlKXQ8dr/10fEyvgBdzMJsL47X2bjwqc3UspA4BrMAwvEl5XOI
v8PQuVcAvB7Wk/O4jzFArNelNYg+rOtDufFinzzv41j9HnTy/Ax6S94xRU1p8iUq
qyF1bnFC0YfJKzU8MStu6H6MvgBHT9bOtiNRZeh1h5RzFf3sWoMxPrXa6SvLrugh
jMxkDHwqTksjKLn/1r1yCewpSP//vBpFJqrpI+0E1iaGc2ou/GkqZ7LNmbntsnXn
5Y9lpuRdXHPCGK99UMxWgEbKO46qBCxP/h1hedhG9XwcJuNpRl6pKL0CA6phKtK9
LQu0AgmX3uPaU0NO1j3fROXrcSicJSe1HbGgCd8QSyaP4aIuqrPw0lu9NLP6R6EL
fTFaylc2snP7ENJa1pfWxLOqOqYWVoBcrXWCNBnxoSuwaCJ7QchG9NN+p/C+tRje
dfjs/3c/oEAiyjrxlZEbKGmtVdnNduHNr3GZy2XTplzGZsrevkJgmoQRX+NilWRg
gEz6BF2XGaPX49qX764eZLO1dVWqV5ZJ2L7wTauoBNtO6FtGMGDCwDct07hP3rRe
9ryZKle/pJgUjz6OP6LBAz2oeygTO+Bc/+DoI76BN4HqVHep95vlNkSwVO98f92F
V3DeVp+kGefg3r98nIaeLOk4/SyskLpLkZxsbkvd+PFcRPz76HdsUnRljezpsPgK
yW7hKFh8NkLnXot+pmoJnVYitw0CdU7sKdFlbOLqO0vkL2EXJrzRdK4o4sjlDCh7
+VETtfB86Xhb3e+BRGM6f9b15pK6tevDu/Fhs49gSZ3d+s86GL7/0+XIQEmF7GGP
1g7TqD7gMu7iowmdENrHHjZwPr1Omxql7aqfKW2aZMOTSpE2CFukZQZ8U20Uu/Pb
pzVRijjx9HbICIyIuHpDT5BvJglyaDZbrbtk/oCJ2J9zXYW2Zr9B8MB547tzRGzM
yGNTFfJPsSY0/RodSJ7mVgBRqBE2ay6rtS8llfhNXd0oK0Nl3Zl3u9Mp2AzN8Knk
UNe93TGCvSKjh2Asp8V2zAG3rNPDaxO9c2CMelbvr0+hOXwJ7AHvhjoNFdZBkjNL
qdtJZO2BA7SIgbn1ntbmCABdjAvt0ErkamuHBJOutVTBfasEItZrdDZSATN4Viky
ydYq+yczffArR5U8EQJT2aVz8utNksfKHePytCaxl3jG58FGa1MTx/LFiPZ1Gxba
7V/7g9/KofGTN2QlTn6XjVLi9Rl9l128cM4MdgalbchsqYdIv9yYhOdC7Q5LeYDx
xcwWV9Gcq+2V8EXaRz0QeW4Y52+grSGaO8IPGsPSuuhS6ir+TV6tHfnObHFoZG3Q
qsem/7xUSPdeFu0TLeH+HDPSvoHxoKT2/eQf/9DQjvw4fXuon2kjD2v1c69fexsb
zD6nk92f/kmOge+CSUD+T5ns2fh1WAZSIiqCEB5HkIHiYv+cJ2kWJawaQsYcGZh4
VxS/iBD3WgZOz+WpvosDz0G1nvetKKYC8RxLr7Ik/gihvJ7JcgA4vrVIgSjTexha
XraeI7EFElRE1fHwIjReOiMPmB0mDs5N1H3k6Pi1Fz18fl9TVLx4cNfTveBTLmqW
GAYoybHo7MuwBw8Ur1f3v0WLgeSYVgdViKK+nxRFwYjTwzrLDPOC9QTDNpisLWYA
1XNF52WYRpGwANE8B5llLP7DEpp8T/kKYiYEP7uRRzmFOUXscNGvTKjbhlTAl9L9
clhW94dTFbVOKnISqkS6aVPJH1FaD2/GCMmzAFkwdQ70A8K0Jaw7ZlexZr5D9JJf
e9GX1TPcRdxdk36prD/U8OnHSk3PgVlvqRrGmXpSjEf1ELn1RupOWXLRav/rHaCn
WWKA+83CzZT0evqf6Gmuc1WAPwo/1TURHLW7mwrde9cb4efjJq7nvkVuQt2pa8N0
OwGnXIsh6mfpUaSsOsih3uDXRb7L+cqCvsR4Grc7y5A+h9262r6S7iEppTY4TCcf
HQmPd32ciW6xxwNIfK/Hrh0/KpbG5AN3pc1bzjzuZV7KzGbujZ73NmfW/4xEwckM
zF3YZSps3f8JkHv6iAlWN0QYhDFXFlv7GHywLjyXl3L2E/FfS1iKzfRNH6WJmmVx
Jb8Q+HEdRZz/SsO02LP3REHwhZPL20qsXDga6rTeWocXYdoV0h2xALdiAHzwpTF9
8b5ryU7v8whwE1uqMh3et7y7k1PUr2fx1D3RiChgIP6bXz/3X7LJtsgRqKDHiEcM
zVPb5f+mF+Vuck2fc8Jk11Tva5J6zLJmHRVsE7mbCM02isDu/Ny6xULd26gH18wY
K6eslzZKExTayBStVguWsd7CHZT4E/uCClkeC42y7XxBtIQYp0avmGiRseli6wcb
T6vgki0y4CV4Ss1XQow3D1FLDX7N6hqsYTHIJ/xr4jtbLro7U/g7kUgu1s992mrO
fALtJrZrVaFb6zs7cRymZ52fKMVUt4CEzck8mSFy0ar6vB+tRxqwoCfC2HHxwzOg
XoiKD6V26gAn9Ypfbt/hyhxs5u+vY5dF7xT+NQBBvjV/lUR16TpScmR13+PB1ffd
xiyMh9W7yEivjSKUGZi0ZCC9ucDvTZe8Bt/P+ob8XDEcvML7UWKomzaDhrb/gJxW
zVcpzS1RXzQVluSkA3pGejQ2BadX9QmfBla1rOVZR+ZgDx9jcSsfO0acA04SesnJ
XE92qPeQ0SCDsIhUwVpxx2V8dMtmFkUADe7n3IlNIsEX+XE4329BRhB8lAf/Pdlz
m4y8KiWm9jpshWCWxxBTeRDXphhBAw93ICzm6bz0gUX+3F/XySF/fQEtrU3Lp/a6
wzfByBUU2IDvDabnYTspKv/hBvP+nHgF7NFhEaSKhiMfRsfEHQOSsNqajUcGPBFa
MIhA9A0pohycKDfPCi8/gAkOAVzcF0gUMLkPumUvZ85sSo757Sv9cUPMNJI6+sWN
TSws7zEv8fQnQSDWgwV4ZFFfCRgsecB3qZjAsdFzxosswiQIbnc/Cdp6fIqWK4CZ
6yYwBumg3C5eMIMDkPUHips/vcvGA07ywWrvL5lSwnRcBQ22543FsHb5CRs4Zq7Y
5xEIoLwA5coubZeFm5Il+wYS8ylSiBG7Cfj7JEcBz7V2qcKGhwK/RaS3NU9Ax0LP
UCL+Ce3ptolghEQzqQHOF/GllzuMfE2RBzfX4To/eEg68ECMEKx2pwl+s2cs/xN+
x2P2yYU9hSaQ8ZIF0hDr6awvatZRy9R56JCFL/pywlBzKL53eTRNyVnEh4AgIIA5
QdiLTgvg3qHnMNgK829M7Xw2RWM5WkLNk/VV9FFUXhTs4rjYfwJvjcaMJzdSZtzp
9ZJ9vKyIpVH1vo7SBqRjlrY7wyPltDG3jFbHciUdBSkVVdXY1jFBeMFIxftEBqvA
ZaETqsdj14tGOVQlXeZFOAyIJW57p/jDhmRziCp3SoI00GXoLx2eDNGkL68Lkp0H
HWr0Ggdd20lmlmdHdNjCT+BIfvo9kVIVTlM03UEQD71pgufVMqMuSnxMhCiadmjm
d/VtLQp0H2nxwETVaZur9X0kNTTR+08AimH0IzN7pDaoiW60UNhvGA6KNyc01W5G
FDdImT+zx8dE3RusEz6mHPPeG62kUuU2ZqjOFLOuGGpXGXg0VqcWo1ER4bLS3443
FBBBxKrhMjH+9ssnBXaX7xImt4vk9DQPvf04CYCxeQgysac9bj3bocCG2RfGFhy6
kZ/PLhxnUrAIYkMWURt0IFOAEjL8bMPfn3A+IGbtq6hSuAhZB/DvTiqfifgagb8s
qS18d8qW1ze4Z1cAvpnSQK8utpTU/lvxjH/y8a8oB+yyZpFHkhajspLfjKBn8SBc
KsLVYJzyrPGTBm94CLlqlLv3hQz5w8aV3yI4AsfEtLzMUm/Im4iCy0LDtBYW7Ei3
BX0zco+9VNbvmt/rpNhZCMFVJPNt5mcBuJ32F+0RMqOBHr1kFAOoexK6cjluUPuW
Jw0kOYubAvEi4tjggHNmTuF/wOMNskuqQGoRS83mvxTPtZH7CuxAunT8MDPqZj+m
vObNGVE3aKVxkb0wylGd346QnaRU8GGVHm9u1tUaQbabj2e7F73eqDFC9ut9K/Px
c1H8enVufIRvAEhTNeLz4DqUc/IRMvbay1cGebyum8Sd2XKkzcj9AMOV6ckMHVQH
hv6FB0iCrxhh69ff+pp7nrQa7oviYsGNw/TE1xxr321l5hXfSdw8fFA6XLPh0Cp6
BKxtety6RIkqTp237wlsouZNALznf6c6iNCFEGgoQxpMpxGDI1EY3DtPN0ftuda6
+m+V6T3BRI+Z8vnGWwU+9sAxGGmIWmpKWiGcnyOvqUg2b9jSyK6godaB/rpoB+UN
i9MyvRTjwMigmjSuPXKbKir1VTsHC788sXn6P92Ct672/uxHUncNYCOm42HDrgd6
IVfrDIIxATOfdhvlJ7Gy6lNFKDNSgBlQRRY8Ufc7EOuT4zhAj2mrBbyuXz0UeTd3
g8RQDy4w7ryv4F9f7fJKIiPy70VSACHBuwSGLGmHAzG7BsbMbGWGuNky+U1H2fSt
+0cJE4MfQ8fX3vGowtik2PCXtKJcSIkdukwFS+L2S43CrFZfHvgXNMnbBRqkyhh4
q9+Kldw52vA3+myu13XkqbSTezKTx7uqu3KBX7Mr3afN1kEiKQh3LzUvBamzqV8H
A1vWCsw1JZPtne02jeAUfWcTAXS0SyCkuHVha6VZWlFtJ7F5UT18tWFI/92StTOy
fi2RCrIm9UTOC41LuqI24UVEGjaIbHI/vyM2BV+WOvRykvB5iaPsjcj86DU5K8Gd
agInD4wh8zBArxTTw+WHA+6AfLN/v0gV4euYgJScTyYK90eXxP9PR91Ev5ZOzP+j
/0uTqYHtVH/onLraKhXDeRkEliiWXOSaYMtyfdvKfhYqpx2xckLzU3+5gzrnNqAs
3Qkk2KssIXJsm2anAQVx4uOUqvZjs3d3bxzzWLzZso+G9BvsScYcw7l+dGGxDy7z
qcWZInbPzhjgC3b8aXqaqwkpsJXJ5v6sMs+z7yIbpM4JH/MJSNmCeFK1NX4MBM2Z
9KwLEc5ErRNxccfqndhyCQiXGeL25tHN5xkRuvTWvBMijSykmRhPATG4YbtDaxCb
M3X18/GPkDk2czuClwpcFzkwVVdqWzNQRC/RteMSP2XeemgMEXCA57hqU1gTIpi6
OOBJDxfAGsQiDp0lNfSP2QTGEMDcz5bCrq7XE2bqe3Lcb4D+kt6Xyo2XclV3bH0f
6XaAzk8WXG/Dw21LfXow3fZYoFDqXfQeLI5yBX6VLDg+gnd3bnxQHz0xdY/nBdIs
cKdBj+64ZobQri/8C9Rq5EBJJWSAOEcxksZeve0AN6SwGvjjY0xjdjyN+37sU9d2
VUPXNM1fFXMLMLaeNQwOqzw5858ivIul5HOZslKOz4ZAYOmHr7XtrqWYWvuC8Zky
/AizHwAPuo+uVCqKFGFWXyeVhIbmQhcex/6dVj81IpHdZVv6hB4ZaULJff9zOpuE
BPw3OOiqNF9YXm9UdR1+UY7Z72TZ3F0C7qmmADI/dkqcKeagWIhDWvSogkdAX9IQ
kcGahSTwmLqvkQL5W2Pv0KJV7ZTJmrkx2S/XzLOH6JixUrhLxRC6MX3iAcYe2iw4
qIVDv02kMuq+UzjXojCzhUT22TALdMnU1ciamOBnxUpXz0hejknhAEpY2UAEMBlQ
ClY0zkP/HQ/SRhS3H1Tg0IPLwhI1moQzDU5naDeQy3YFFPvvMDEdlYSJKslq6idH
4iNF5Zy3JWDTc6XZiKuGMj2bL7dMj7cHnfqyCUAXbOcIRg9uNb4RIFFaqxxgr/yX
Cv8m0c4PXjc1UYutkGR6qGZWi65QZr2kM6YSmFYEbFNUg7adyGXrzV5zSuRIaBWh
jOy19IEMYOdNpdvLzJ4mXGCHpltgHuQ6fS/FcBK38ODYZATM/X//4+MW2hhXlXIN
fe5RFnIHjHDY7D+JmozHUpV/2S4NfdesCNDJWuH/Sb54KebgVo8BPoVSTach3dnd
whUIZBMHt/7nzYGcOUzgMD8U5NmKcOodKvwVrH07NyAGDyhCXPqXm9bnQq391Btv
RTmIOLU8DovJHz3R+FVRHoPaddHFcN8UYFE5vxu6/KbuAunqAsrKp6n6S+o5X2c1
9htbS+X9oEdUMFm1ZtP4y9/AhWidEV9SM0gGVhM7Y6kTUjxcjqXa8hOvDngbAsE7
R2TKqYFyZVWyKq9MMkZly85O/NcYurII8/kNqvUCIJyBewAwNQbP+9vRD3KkMcdi
RtTMJtxY58eO2roV9QytGv7lrOgcSFidDcb4hgeLz7OAe9C4F2fmAvEPv8KqhQXP
Tc/2I7U6dg331dLPLRJoec7u/chPEwypfUvhKVdQKSBBnLt/Mw/ypLyIvnAih5BZ
6vpIabR2jLas5L73S0b3hk4Re4Os3tJurrzUN5AGjycaRXsDJ2PmQ9lQtlzjyVYs
FlEr+ydqYJQ0IKrQvXtFfzuGSBcsZUQRHLEh7pY/g1sfs0BWHx9cv//OuZZ8APvD
C7VxXGPxEGAvQFdxGmZaI9f3/HP210oNwfSGR5gps3Chl/tl4s2EriP9PANfMAeS
tCm5Xe7EtZfQzNAqBL9gLTfo+BeDfR/jiDmidf+iq5ZDBE3t8fhfLKZCVCU/ZO5n
LzDnkgXAVG2fK60u39kz1u1PV2P+0QM3OCGzCC+gC1bS+IzyeyqFpGyBz+vicl86
YaCzGMQc0CEori8lVXPKNczsQi+m2cpsVyJ5CF2ADY1xWBbfQxta93Rb6F2+PHsn
9uqlv5eke2hhRTT6x/s3YuxFaDJby69PfH2mn5YeAFlU7n85Rbs1u/oSE/zlYsO6
a9qXEdhbWkYZSG9dve06yPYdpANvgzEgfmxIJYNVuCIQ1PpOqhDsO/yyo+u5VfZa
GFHWs0hJP68XhDDd9tiz0QdBVY3lw353Rt1H/3jh1ZXrP21L+tRggSta+YyPp32G
c7QZNX9nVdud8HnfAAtkgHq+3LW9gtPCYKqXj0vm6Y/IqE076uKPqM742H7e8i6q
68ifmxc5vivVtcIa0o4OKZi9zxwsgvrKZ2w2dVROckc48lpW0BOp08IlorHT0Fts
EFBnFAeJPf42nQmysZIQAz5voJrReWgMMIfoYjNQN8BK70dmx09kdistHPqQNuBp
kTkhXQSRKDiQle2nAA6hT78cM5uDmYMZvs4xuG/R6fK1oIw9dO26HyZame5hkmeC
SEavFyCARVdZbRp77dsVUgHI15gp7BmV07bD9klTtvcDmP0CUk55Z75PBoxyLBbg
zn/skQDfohH0JyjfrUl2c28YeSW2jlzidNqIjpaWNG5romv8N4aTw4WgzE2jvhw5
94XWtRo3FEupC1aD5os6Izn4XGtlAnsNdX5wTX0wp2Vs6x5cq79SPq5bRn6y5zkb
9sm88WMekO1aL/y6Fvku8/ASOqhbXoQE5VJyOmaoj5FTnCTZlxZ5K2195++VbTX8
VZoK02a+ukW5NW9TdrcF7DYpbkhEquRJcgBdBz2EHDbqoYWN0B/D7xAG7BPIZ4kH
+FO6+7/+ZwRwE6IqkMSDJ55INNCVcPcE2drLNvILBPPUshKgruhm7HwVru+ydouo
v4pOpNSGuNiUOFqytsVRdR7vqJMbS4BhfvsACqbrqFFacxXraM1/vtyy8IV7aOXi
RNbtgyCEUD1C6Oyo4ZZhZPVO4PATbqjPAFbTrcUTtUUeAa3ze5HfLXHRsXx3Upj3
BfKzIx++yShwhKYEXg9oac4xNnt/Xk578rt7cyGd7plyHTQSvlIboINT/AErn2pP
xoDGG9FAfNVQH3oBFOIz3kF8bi2x+d0MxnJpiIuzH5D66TgQcyEG8hI/Gnmz6nws
cEMW4ozxbcbGur1ZT+wy7eS7MbT9q3R8IyRDs0fwx4Lid77XaEdmzLCHcyLg+RIW
Lk+kVcllHYKxtC+NA02Z1NKKieX84UFb3H4X9FjtRbvrL0ms8CwZCnqgbymE7/Zg
3JSttd5zfRGrCMPdeJiFoKs99oAugzD1d+4HzYWRnbVlStVljRBnCYTo0FmL73kp
XtM5tfoF7nPGWRVlPjNU9OVL1Npr/tH7w9ELL5m7/ePor/J0WB22tWSAD9tw6XB7
nkJCQ6rPxKfT4GdzOtZxLoGbyTS4XqwSwn4jVWi1kTTv2TJQLmO8k6URb5ijXEFJ
tzWvn972jjc3qY/qkjAMnju8IGmxqeQbeK3TDXxfK2CYeb4CSOndNvd4G6MmrxFk
8+Z0Kx5UMrXl/hxc8QjW6rs1JinTjM4QezqEEn3i7M88KTJgKXhdbmQYT3VQmNrW
HMAJ19VWf3rw/xTWses38emcwNzQ4Xgz3XMdouiQTnO0MtKx5VKrKWYMIRxUJ0vg
+vfGQ8/6xCDBTM5EZIZY+czAJnZPT+yQ7OdMXtn+F83kWG9Gb9WThXhc5+H2MsW1
Wc0Yj1ww3ultccZqGjarErxHelJ+/yd+yI5m6YPoUq6TSBcUEHFO095qrJRvm790
75e3W75BqWgxifKNDfydhQeOskVITSiMT01k5GXaYiYFfCkKKqLubicU/yh7mvAx
l4udUrFlgtQTIB77fBkyFANnUMoYWCqQzEIDoRvSCib5st8lQBdOM3wBpcBpthEV
ZAt8P1YA3kpWDrapnqLeuQbAtOWSxcLCDmJm/yJgRuEugVoI8Ull7XgVHfK1dOoq
EIrEfBbvFG660ujnasyyd4qEHCq1/5/7r23gMMH9JJmTEDI/cplJclhN3dub3liZ
FrqbLbc5bdviBC1yYyP1BEZmRTU2NvFDTa5Af0p99Jmaacm5UpLLZ1JtYCWOKV1L
hI6fk8uD1I+Pmogtdf61Cv6G8OKH1MRUkN45YbPECO8dSM5H6hq7s2V8B3v9jKWr
5qgw+mJfJg/YwvZp2HabGSP9GTX150VESgSm8R/QD841/bCp8Jz30zJB3H/lASSf
DqDz3TkisFle5VTgXcTBmpTpjA34LnC4DDRyZ6vmAizrxOkiMxTDCBIoMjEcfNsg
FYf7i6bGeceQ97F//TJvqxJ/fgQM+lq3S/MdqX/T/bwuDd+u/1ZCRJX230IOCJ1z
ogNwsbsogpfuUMnkZmN0YD0x2FdwFcjK0ursxovg/1zuVcXWQrQrrMiSvpAOOS5B
tBEL281GZXLgCqF/aIBHqHkLSooIMx86yZ+rdXfP4bNR+3+kPc3PQJMcdKoruZhU
cntIJGBYNMiaNf2xlk99/M3F7EKWHnoDFPenWiQeFgBRVwtLd8A52nz3hv8TTARG
PB+/UVrgxKWxJmJX9kRFRTe2v4UavHdB5up0prMwOSymUNkOCbQU7LBqEClTg7DV
3apQt1JHCx4ZVieNJQVqRMf0Lh/gMRUerG8reS8CnaoqJslROiFYjGMO2zsTjlQY
zRDFopEwuHDrGbS2X/xo6gjf5RCnaqVuAYDk3bqOTOiY+BvOgd9ozYHPQSNYCwMp
joA6leXgzFWLAmIZTTO0OwA6WxGZym2kwtMecfvgIvTGOFZ7hf/jOOGuDzEiR6np
DuTzNTDVHG4hLiP2YoNri2jeUgcsjfzxWaY1C5tWpWHMu5TDZ5yTRlLsA9cqKwHp
oDMMPxfTHe3REcc8fxxKX8k2nzVDmPIDJTYqEP563M+r5RBGl8yX7TnU2NrWLPXF
ZGMZL0komVW4O9K7JclCelXt7w1g/Io9pUI300k3qkjxdLR6PRESkZy/XW08A5vw
MzjPzcXq73/pQCYyuYa3OqCoUd2MKt+YzLqIoKszaO4du8SCE4Z78aA2puK/QgsD
Wfv8vQujNLT1mhc1/F0aqV02SwsLXHGIPrCqmq52sKBvN6WYEzg19lCFplO1iZtj
acy6DHeziCRkAhmqnuAvTs6wcCHEkgPoYeeiCDT4QsgU/NRM7/pdo0TBkk5PBuy4
rFmIgHlTlg3mx6KcPQRIcIIU35+Inb3sASbXvRPa40vvKfiiQw4zkiH051JAM59v
XR/6iNb2pZiS5n1UvJVLzihEO6vwT0r5wMcB2ZDPGRyHA6xCkdAl8BVIJ7ipK7vD
lh/b1jQJrl3KlG4KBGGCUlx9+Q4z73jj9G4xLLoyzXnf1RmuoLJr7gGvRqXSJilC
FX+o5VnMkYTq7zZP+wDk78qbR69ko+Go/s4WdIQOkBjDWe8ypBO8XIT/EHhm0h4x
v/bnh3Ciovh4T8zBqLs5HolL/uF5a4T2G1Qbr2rFaJRH5ou0JrzBJmmzdwf6RDOk
tmseuYdWu4ahwdy8n6OknADzc1YS6iZi/c7q9Xlo1DXRGOJjq8clUiro0B8IWaGe
f7tFm2DGRLHU/gBVc4ksNesD1GyFGvAPOg87vWfx31pqEH67vnjO+F2HQmHdFqE5
VteF/NmKblfKb3AgP+PGFzd6KB4r5ahSHubClYbG+gKm1dmhZxwEJ7G16T3zvuy4
AR556WDCK666aVwE/fikihLkdgv9dYA/7CmLC6eBATGPBGyrga+oPtHXfWb6W7ST
btjUPuxhn8KBKFKU87b6hDBEoYsTEtQ2d7ZdN8TVW26xpSIxr1gCwf7oeSfvHh9S
Tep5NgxV3ZcG3EqLpn07tsN6dFTX0mQ2reZ1rxexOhYgYriu3971y4sd1LdQxSmg
tzgIqe5vrVMH3eoGKpjMsjIHlOkziTpEVDlTPmr5GvY1TCxCd3NY/PmfiCVbYikv
TtCACiul0QBfLpiIhCmb25H90S/pt3aMUpcYr/84lNC6xxZbPtZwFOjIg6UrQ4Cv
6hVu806OfUV8qNBcjYB7ib4MmFFD7NERdA4RLXg+8mFA4OHw3cO/Zga8iQ8C9giI
NvsOXlrfgBOTbBlGEOyFFvSsI+GabDF6wCkAO1dvijMzkTzzasL6szLROEEH9zoJ
l49L4NSMgHH2sd+h/og6RRajDRWUj1+3kn4cXo3qvbU6kCseaH6gqJ/XRCEEO89H
AM2rw6kbegw5aHFnhJug45evB1aNz2/Bt39dmaCy1UtjYQyUogojH5IpA7aCAQ65
SpZzXGGYYDfEkEDuhJ18l1iTAMUiKZ3JhBPYu6z7JuFfYsHfX8ur4PS2fGTDq0OD
6GQnqwyfS+BhBprqyeBJM52XdDcL0K33Pi7vXATUZST5r3mylMXfwQc43o8Dq94P
zCZLHov5pSCRlahly/7in6M2MOhbu+3u4/vBhh40JGHkcyZ3fHDr3VNDx31Ol+Zm
6Pc/TnPWDGorkEEqzcFLyWPLCc1qmfL8NgOyz5ZmOMiBRuXvM919UfQg7A0VZVvu
azJylr5v5ZgFyBwxACqEf8hQpzjYytCzV7U6M7tk3HBmSC3R55X+z5SCysMZCeDH
D0DjQoh54KSM952WHEncm09h7Vfu40muMfsBtf2DCuWYOyyZHEoZkn0ampmtCZ3r
RlE/Ii3yg0LQS+oZhY9lq3XQ6fKZVuhH10nXMiEhtfSzCxM/fRhLU09SisPDiAfE
Xhka++DJ1kY7AtBXwMJxG5JodcFiw3BUpkDZVI1JIQZAD5YQU9j7X+YSAfASTj9t
rQKkgR6/cNHxU8KRVndEIyldWzE+M0CG2/GcmV58SBzhs/GFPQaxAXlrVvsuuydG
OYAtLtHdYN0XA7PR1UfWLSNKeDxCGwRZQbMCfdvTwnjvNFwXFKETjlbGuEVjh0Nu
282iaNAt19X+nXnSfJl+MsqPbgvG5rCk4NzHXoYf0vqoDjRz34/JqED62kNvLT2G
mfpd2vobggtUH1qHS3m0ek6Vw/b6N7eqd8HyjGM5IVGqVy4XSSL+X8i6XSgT17lP
Wz4Hzuf+4I6diwOnQhcvm4tqzlruz04fIoNz1PGa/fGOCHxIkVPYgmPLgOQbvuSt
RVFjpnaxxU3s8wjKgPNQP2itU19LQC/A91+AZ/ilAJQSD8/pqNeie1UwbBOCCSgS
gLG4cJl6+RmGosRHFHdauNCMuqZiOTcF3g5oVLSJxpmWY0TUjmAaXExqWlnnnkfD
1fNzSyErLq0GHP4cyeJRzkw+373K9/+8mvlmifi3qIhvdFtyVLGj3NSzzcbqwosp
5dAu0rJs2kpMN1rFGQ57tXf8rUT07lHMrXWKNjcuP+hV25dY0xFEE+6SGoVXqESl
0Jw6FXAEv2472XRUpAsdAXeaY9+Vwf2Aeb6P/0HcpAYachcYfSii74edUPdKP/93
R/71hRgSmznIGOioJVjTMt2ChUz5dSRjStQ3PpMUeJ34YilS+G7cz6KOq5cKqJz+
pyWd8z99QISwXowGLoljU12FABNYbwZPcKIT1q4B9C6y62YyTmCruHmryeiILwGK
PiLYwD00W4HqyAn3HJUU+jApcib13fxsr4iyEkTw2TgJl++KtZDSO9svJvysi1xh
UpDVCVQFYtCKP7tLxImdPL/TiiyVMRJGXGT6j6tmj6awTKg7/jJdunzdPBz/OFlG
PHN+1lg/2O6C9P1DdDZw9dOdMh8TdSXgqXipJqEp0GmqYMd38KJw9g/TagrEOqLq
nxzYVfz1FRXsDl5dO1wtz3OVAIPhzzm4Oa+0dpPdZcf+TZLapmgYVUCBL6dvTp69
iq4pFmx3TXGKr+0nClAZVGTyPfJFWLMF2Wsv4QQN0bafSQfm5pLi+JVPBCMNEYC4
bNUuGfenqCyVqDdqgfYVtWA9rhvD0BDogknZGSSWVb1h4SqYzwx5BhYLzQAnqYyl
B7ui/r6Hm1ujhjoN9fObcS9o0rNRr1Ei79ZMYX46Dzlw364LeIpQjahHZy5fRFea
e1LYOV4/vPDr+nWfXBPljvTF9avYME/3Knvz0vYqtpK1Y/0MaPBWQv4LH91yBzqt
93e/SEHWPXsE37t0lpHS7s8g0N4JrdjhFUXmnDbEmHpm5zceObInCdgZFwhsahHx
bR4yTVpv7Bh5XHdECT5ywHPhBTsQd0dOhGh2z2f54Pe4ecaE0nq0nBszZIMfwFmL
xJUZcvZnfVMO5iSNr9dakDyiZ6ZCC3WOe9mQddUU/X7GkibwPrRxTY+dWa9bO552
2xc6WebZAirbpLMg0YlVz1sD7TiuKKfjbTlB2su1Lo7v9MldLOQULOAhPTPr6HH6
IVoCKf31jSd7RKH7Y+kB0mUBAv37Zdtjy8ctPJjeZAR5P5QWbUUZzJjVN9/p9yFy
n0gbosp7+kBlyn+SdZFlYI3qb1YCvizdjFNwqXTSQM3W4CWtGer9lKp8yS9brEkc
D31I1QA1EBlxmThtjLQOP0ofFp7tuOMC6EBKs8bkvLavaVRUMIuiy35c6yWdERTP
V4t+nkmxEIFujimEzoc/9lonqJTJz6nmwPezTTGyYR1C4hZbjjUK457R6GSosM9a
88IcH6G8uc7EysaL3ylQbmb10BAxWWD2l1AYukx+/yzDXaHX7Lr20e9gTCeOSFNj
P5+a2GJncs7mVahS/Wp3zLZgZSalIgh+zfFX9rfGfCQC2+racu0fR1Q+38F9hV9b
dXaHAkhB1c/8En+fCRWm0yMCX1dYwiIoevFa88JVi7w4L/tKQeaNom9X9e7ruttm
DAfcCwOWEcCDdhZmohnKmGWvmxJ+sQcgtuAsimuxgxbtdnP2jh6QwdhfDlGxt8d3
OejANeFURa+9PnN4G2Cfbad5OIgNeYqzFK8Rf6soF6OzWBEeYrBqtY47Gbm7DmBy
AWSowS6sz9xfEgpYcQTjNZLnImHVCL8OTfE3XkpNquc36ArUQikMtcArEV3ko0e1
LGSZOJcR+rkiUyKxjVSA06U0MEHx6I4YIn7S7ToDzaJRmAio3sqq4Fj+XWja5sAt
s+Shwceh6rq+iW/H4BjOUkS46jwF7RKhHv8Iswc23R41uCawCHf54JZZ/aQQM68o
zFQaV0/IPav3eevlMU62Eybsr1+hHwc2+kiwvi9dvzzOh+2Wj7kkpWR1gQHyy+wV
aXC0eAWB4tu47rR34zx1SbRdmgP1eHm/sGfh8ayvLVnQ0EeFBNASOtrF4BBCkGC4
xkCjZQJvQTmq9uTgqaEIlqZC7JOPFbwwQgJ/F4vw9ZtBeGzAxednLrw+x4bZXlSg
rSGBzP1g+w/qqXdeH7JVCp+MDcWngqjtgqPmQHBCGplLGdBUNmqeDzwhxhUxcvwB
TBw7V5GHXoq5/X1QLkjrbW+96K9s6exstS83Sm0IOJDDtbB0XA/YU1RQku0MblvH
uAxopTBzchkLmf2m92gpYhK7U9I15PonIP++n4ziUnybbnkdnDTVZVtg4svlZzob
Qq8pNkh6hZuR2onzpicfhSvDHK/UfEzjAI9tffKs0gZynK+fgyJ7b4zqCvZhvmiY
9UMS40NafTL65YFV1C9jDDVQlEvpBWn+L8Ddujqlx25J5HVPZYFUURclCf16uKNL
CWVXxaZBWJaM2cj74QFeHF4TBLTygYxHo4KXZxoNeV3KX+hROG11fHgL8KC7i/FF
Np+tX8j2imQN3S1Jh5kodA60EMmyNbE4GtKVFj94xDSbKL8z9+7vwQg8byWqAO/F
btLTFKpeswxnd2QFR9Zl0Y71KnAU+tJg/TLkcOHFUY2d1gNDV3mgXYFmYh8Mdhti
Yo+cDTVnDiDO9rPzpk6IL/Xb7fJVdY++3XaXXq25lqP0nGk/xPPVBZEhR22ckbIT
ggwvNWjzpUQsAjrOqE9EMbKEmZvBjAN1lMDRtQJPY0kKkWOPUy0szDY1HEsWM19V
h3PgHKRB8Ysmtm8osYNPp7u7lJu8WjYn7CAalUii77GvZHkQm4pDA1cvdm+gvodV
DCjgvrfFjvhV5TihBwHOwE+QWzlNJ6bPmW1DcC6CwXnU30kmTG0dQhCm5NcmBhef
HAZJTGjd1hYjuaa+Gq6zSuCJAOLvd4XKb2iqrUPUFsgbkhmQ1WUuBr1k+OFi3HQ1
09/Wm3YyotMOBM9a0+fLC7I9KFtMur3b9Sji21rw1UW+2vMfzXzfd5A+kOSqgBww
wxd415NDnLcl+xfj8PIm3rRiP/jbRevIZxWqxuXm01BAZU3fouBCnDMWQdAAkSyj
SwysUQl/Ip5D9hJHif44qBAFKOuV+aK/AK952RF62AGE/gBi601ECwNrtma6X70/
34q5j/qvl82TjFCtOtBVVOGvjaRoUhizH6g8DmC/p56ocVA2sNY+xxiFSHaqvzF3
TPMWkBnZe+rfGTl0BsZcNS8GmId7BZooWJjh9b3NY493HnUPaw+xsBsvqJTJQkIG
tG79ejRyB/v2d9yGtMNZaBn2Mu9YoWGq2EpPZv6N8Io16wVjF+dUdD7l0wb83mUd
dTeRudd/2TyGIYWDRbGoUQrgVHa/REKQVlMYZHYGrSugTaYovSEAC/f1ZnhkYr1F
vcOUz1ijUg09sv2BR801GG8a7XF5uirhJs0oNQ81pX4TZn1p6x1uXtxEgKzQswgG
AJDA7b1B2dpnwj9LImQiuZqVTs2w6np2CXkzhUzpsvMMO7Of/Cd4FSOgqgUsFJpa
yKn5up2tcxuDfcX0EenPGQeQcH0b5MogS+BvlgRtP4j8kTtTuw07gpm98ArFHRHZ
CA/eiqwxHwrMq9NaeR9naORi6kWBP885I4JghUTMl4XUD64H2MZk0oyzj6UxDhY2
CYRAyK9J6/Hm40dOmGZkVr3VQ1UWEcVUvZ8wMWDzTWwkwx7lcW9Rl6qclgpmU2IV
OqjJIQRjljL17iY3Jf2yvlKddJw2WKIMNoZDEKEdx9bYUmhndjvydEhS2O1OaybR
CwVOJZYe8UtzBDyBBTAfFMHRhKez0xmb/R88rHnqqrQ2VuS8BpLu/v0/hjGDEvxX
bnAc1t/mkBHjGrf3yWJqmg35AecWb6dK5SnNemo327fE148h4gJ1TMYU20ENsEG0
p7Un5BLyejokbeWiunpYEqAWsk9XHdjKWfZ4ApNgCOShB7AqEiM1K1lVvWc41S4Y
BsFtx+UbFMtJyfPT0vDmdp0nMThEh5SUqXMGD53cCgM9Wxp1x4kLV/0DyMIlFZKz
AZJIyRNGs5eDUNBQXWjK9EIcQLioNVtMiQ/kd9KbEG+m6komUjrZnUQukiqm6tAe
QB+xQJW/vBAP0RB5u/sB7bvZZW//+JpGe5qQXr30mWBiDIH3woh7VdCbbmRsErov
m1+kpvmJQmfGuLGaAuO0Y2UNdpMYTt+iY1r4FW5GVXyS/KqFh/1oj2rOVFFQC19S
P09Ovat7Euc40KtlLBFukzVXudm5A1+yWfhop0opYBfcrP9QQaTA3PhrOsRMpIS+
YfQjnMCpieuzIlVbNCcr68IfMsdSSsAQaTUbHmYvfZqmkVXypKXT7gnW2NL6QwML
qWieBBXL9ILXWE8ioElkx99HN0cmBNk5RW7HpnQ0nIiRuDAbVCUImfts32N+gBoE
8z0n6F5D8rVx8IIM7G/DxGpqyB8U/Yjzp3s3YhpbDMJyN3fgYz4flE6ambo9wbrQ
LWIbOx8hj3IkaIuX1ZKbZHcAKYY/et7H1uM9StN8T7QLKR+n3031YNIPIGdAa2fN
4g+etY/Aoh/CXFW85HZX4a5d44DeK10GO0CSVe2o+98OIjo0vF8deS7/5k9Rz0rm
PTvQ+JzO6t+sq1xmu+or9KQwWhQOrakHMnmOscfjYMeenMSHLeIXU+z8MKjxBldk
eXHHilREJrCel0345ecicPu0KSSoTIGDknye44dSH+z/Sr0pgSMGmxUZmCMM6hxi
owlE1KHx99CsM4euOjnm/leRSmERV4SJ/TV16B5KBzEjl0bMkXng7V6i+/93vgr2
d0ZNXKMAoB7+/oFE13xnH2jaQ6oqA4iMcC6F438jGUKDwoO2wVHbJnQHxkQkl5Vo
RDF3a4cBmYkq1yefVqY7Ygf1pWFM0QGZ5rAkgyLZ1pizaSTm55LfHfexiZCHiDkk
34ae+yorqtvrgQBnNydfZC1QdJg3KNKV8POIIjkgH4cckTDwHkrTIKzFfohtGIaY
YiQj7bKG5p939TNRC6ygKrRoaDW6moyHvJGvl+9EkEjoHz00c+eRrb+hURZSCJId
Egdwg9w0Nwbqy7Nt0e6Y0q2s7lpb3hnBOpfwGr3AcM+SaIfogkpcN+PCi0oWEf8E
uuZMqLnAJxPEWoIVLT5jDbqYVk/qJKpV4bhtnrY6AeE1DFjaeZfaDSsFGZXIARfK
dQAWbwGSajOKAi9q6GRvH97Hh0xPTn7shkPHiIYRK9Ce1Lyx7ksEJjlYotdCD117
TipmEq2Gzc8DHN4mgZjAgMqZkcCTabWfRR2Qo37xyXdGLYm731JLh8xHRLvz5e6S
Egz86KSxD2QWj+NyRFD3j/SsjI7I3GiMQGdrGO+xkrZreZxhLMTtwWIO8ioi3UZ7
jaY7vt6Vm91nNUGzza9JhOubO9fkBLJ/222sfmgKFIfecqwZUR+vooF1shhw4Xyb
LP3LlkTGSnLRDZhseD1TQxWW+aulhppeYo3OX240dKeVT5phfkpVsi/jGix39Q3k
JMGdbyQSSh6k1oyWmkWn0GtuJ1+S/mYHigXVOZ05bMi6G2c81mkcKT7Sxwt5FmTK
xBQ2CxD4e3pScDQ0KhYxpwhjkk7a3ZlA9TpYmCI5/lVvBsp2DPA3adR9KuP0z4Nf
PiUAHMpYT+9/yHLDvAO+1JKInuedrOmwGnhi4uk2N0sLzC168SrNVb6DTuvIAKHZ
wGBY0IMEzrxfIS6eYKwNLDMgNo3KBGds1Gagxl3loK2vx/OFO15xKoRC83UqU82i
g8CkAhCfHYVcVjYJmNBeglq7DatjMAZPzPUINkHr3WpDhe7drQ3jxzeq8MCdv3w2
qPocDF9anfZZiJLDMzvs3pMYMxFH0IU2til4w2o/Wja/EMdZPT6CcL/zgYyLH48E
Fghue8vmOvTC+/xa5lm0TQ64p19ZnUi1QrqO/m6CwNLgElk0COhvjXMl8UWUrtMg
ppPBcH1K0HDZeiS1yaRSAnYlfW0AnSzD97yG556tft8uKTWvUVIdO1eyW8UbkZw9
iKhhF8MDIJTisv7HVGDezuX4u2agxZYKuEEr+PY6SMldoGAL8vIxbCQlzje4tF++
Sb1TyRkfuppUBE7gMay2yOES4xpc/ycik23Mxqafnanw5zN9yrTBvIJQEnFM1oaR
UAvMU3o1zwW1QlPg8SHmN/VA6CaW6FuAAIIxQHnFO1VHYq+h+m+fpAF8Bu/VSE9R
B8osiBAvDqIDOGS5TllISQW1JI5XcYhpT5TA/ujebXWGoR6T0UFG6mDTF+liji9o
kMLqAxHm+LcjWSY9TsuOIgR1niGZPPuBch5n05y1HAFGQsnoWirl2Q4Ufh+9zO3m
I3qukKZT5NGOSB/i3bhSea6UuMxskfk4BweDvRwHVi4BP/DsvXnRpf5NFoQMGyB8
HnvTwC+rvij0bP+FpTihHk81aW98otLovNGCiQtHEbHYadqvDb/q3knH/aJive7R
GR/D1ciQrHwZs+w6jgN+QZGQvg1NM/Mm/YVRm8uyyL+uvC6VbtMniynNviDwJBI/
rTiQ76hHM5XI+hahOgkmAdoAyYQAk8H3Y/iqEbUtMlcXVubMJPzztm53XFg+ICcx
6nqZGUe61xXMkaysxs31+mHmjAA0+6FmsJv02qn+2RWlEWohq7t9Hi6b65DL/m2F
SqJxApVLqekM60OzTd/5W1p2zG6PRcK+YMe5+M+lOsI8PG58DyA/LITQUJConrXN
nIt7DN0t2fyFHruWyzsDXO982/6Z0DbvBH4Ux3qfqbY+LXbMDBbhGbyVkuia4GL9
Wa/z5BpHX/tk4rgMNtu5P2J9QX0ONDq3Xoy9T4L7QdQXrzLv/qQkCATkzYM62AAa
7fTTWEx6YX9bstzu9aBLoJ3/RQLqfPYsrhX/y1tiMRJd/PBWYs33nsu/FCQL0GHq
VfhfxQUOAuYz/EE8lmSIyFhwT1D2SS6AsjToO+OkW1N6fxroVKGhZF837BLrqVkf
m160//eD006tK8Ug5M1WNV4BsdXZfqnzcc7N/+R/37T9Uhq/10U2QdEYpILyw2N0
tcRTn8VkjdreUx50lKgNhM3C1Jn9n1zoEgJueP3WgqWFikEpFiJnFPc9j1aiHpcG
MHGgsHAorzpe8nPelt/1o6P+mSeRLFBuImpTDW113dG67wnpeChsO0VwX5m/rNDH
qs7VPKIWVfKT98QkP4KC/wkFIJbpeug/hhVqHUHtJXvWPR5h1wsg1L4ZBfXybhda
kQzNa7ncHthq+pQMvY92BzWpmLkwdq2aOGD7TfbAWJG/E/50ypcCfpdiFGMrAJEv
lAA+rTKj6qvJEZNbNoJP5nS74dF+BkLX9wmbp59RC6RUFCstPQQImFwpqFLZBiha
lmSOeyY/AsNmcZ7227r6CegqT5HJJdw5ThwzL7wLJcJwKBAgwPN9DvKNVqHsgbWN
cD5CUnZiLr7GUz+EF06Kful6imhl7N+Zcz1F62OEgS4qhtEFOAFNZdPpsz8cCWs1
af0lYHeiwBdi5A092AxpM11oLve8EB8T9GNWoGZpc9PSaROGWVhWBJgRbZN3ysCg
vILetNMXia+5aigD/Gc2NKL/XDKlAX8IMh9Yb2f9MBEPkhsrrOGMrmj2yfLN2ZbD
eSeuI+RitFn/DwtKs/MDtINqSe+MiP6ZxSVLZEZhFieGdWUVB7MxgJEaQ1Jdr0lu
r7Yf0VQdQ6Bwksi/up6yLxYFM9AS/xaJtbAn2uG0d4vM8Z4sPmBKz0SovYEkBssr
dwF1O/C49dHVIf1mSM7GYzrJ1KL7dFcRY4hX6qlDzysFACFzZYNpn1URV7V4hbcb
UOCrXyAPgkrcgwPOnNxKfbBHEbmZTQUFzkgaL4utDMECz4luvKIlqOKRD49Pk4k/
XAlkAF84PF5bBvNNKsSqgNNjLObzQGaUDDavE1H5QerKVdopEKG3dVqs6ViOR7iO
bafk4TVa4i0/NVP8j0OnhgqFB4bTsqWFTW0gI9LBO1Ipjdha6gI3jVQ880lMu/m0
xvIJ+jBpJjJI9cox1sFXXkefTrUUGK5yUqmOP7iE1DUwGUSP9FLy4kuVyHBuXQTV
wfS76HpJhBwCpvudk9HdOb7ao67OrT59GjuHlzvtvy7STnbCZJtWxf6/IIq1HiHM
BwO2iE8MGCIq9VzJtQZJiMoJHykIXWdQxzgm2tyfbG6grG91pigrIHDzZ6qDnIaL
gBpYZcl0zooiWdVoxQ0OMbhP8rzJJ9CM2VbPkX+T/Y8DevKK8OkecHnLqDbiGQ1/
NuHJ563GK/e+kYzF+DFMmQeOlnJlDidGjHhkyaaYjUosOJxK7DAqmBaYN2KFkdw8
oVjWSnaNMuVWXyhkBOBgooxxtxaTEGXzOxLPIg2oE/4Aba7j8Cuo3SF2T1TjXdVj
5lKSoKfhWnUDylWfgbmC2QPAomVHuMrlobPl/Vs5pGa/uH3vZQbu1Srx0UVwrv+o
ACJNp4tScf8gCtpJZS5RT/NUCwtyjes9fORLSnNJtpGhnk4tKVaFwQUa4Lf7RR9Y
sYRfbRVSy1yXMtgbsAdJYEv4J1b7oNn96t0CJpxCU7Fc1Bq5LgzALjQNLtMVKq/f
HejuKZKCa6vd7mN7y32Ba85JhmzPfpFEU7JT1Bp0qdL84NKgHD4nz/nuyIxlf71q
fywoJTerAUVd03nS0O22e4f3z/KInnXDR7LiJWVhjI6DTcGBkQNd86vIFpcZFO4n
CdXqP2e3MJEiN3BANpfbz2A/+dMOry2thUX99adPHRmF2UgUVLSpILkt3rXqwfvC
63Jwp8PZZflgvi7CVW2MhPguIqwqjH1//MMPWD4iVWOqWd715JBaFb0b2RuC4TgN
O9WDOFO6tIf4SEWkwqt7omilk+EMqnkpVz49DiDYA/EB8+dzeWydsDRMD7eK9b1L
uSfZZWqzRhDGm4PDkBofNABMtZSdQhPEHWDIzXB3PsEfVbINEXSrm0gQ3TZJD4k2
8RCWTw4+Pjr4kvpSZ05Ixsv+8j0WZEwF/qtWLxuWIcarT/3wQjSZH87PLxaYjmTY
iy7gflRctUjy5FfsCoRYAiLddFs/U+OCg+qJ6Uh1jmG3/6QQKaqOlRUdk2Ek259r
64rZzhNTVdcvwGQBntm84CsvwucHeYymsVDH/EECuP8DOOYuT6rxNSgc42U9Hf+K
S5a1aObBBSs+3NA65F0gmAtkQ3LOsllilvDcoPMNCwJxnIEQOjoeiapNaXuFKvW0
ADFkFV4WrBicqCt1wcN4U5Iyb8Vx1DDqg/WjspKPO9hNr0KAbxYJdk5EsTt/7lwn
+b1xTy4LOy0JwL1Ze1nYt8R1aBU9aUqEf2/2T4sMppFVLpHaQ0UGxPpi6H/5rc2s
PUyslr3vD6YMu03bNky1ArKisUwsGqVD4dnAD7ld66qk8w86TI0Wvb2s7yJ219f/
JpOJeQvFGXoclSrPq5PVPCHigMiTuEINQej/3v0Qcn2zE5rS3JfRm2QOWzC8uOiT
ygTFR866bns4/eVAJk44PzbdL6wcnMxvOdb8wsDkjIRv2DhDMg3nJlWOLuFmqHxU
rA6CeYdSEARoWfQQ7ySt9rFKSiGKMm/MaOF8Oao3J7MzdMoE96KXl9UlEnsnaztd
UtaOisvi9cbGNbehvGcowMRVaBPu9PYRj8V7MEF6/K2aYuQJ8UW/k9DHyfO76+ln
KpEhGxgqC6AVPqMMq+WW3kEbMbDXigcf1V9v1vrCuPO0UU78MfGIjYcrRPwXIwfi
81t1WK/FD4g/8cytmBytXHb6kRQ46H5Lm5bG7tybEl7kqXrdVR/JXCD0pCms1qG7
DTkOfiXlZ7eSsVDduTEkIRWhjkQVYArQfqwANR2DvFBapsMcQJ/4ODudX0xY/c97
AFpFeH0cm4TE2U5zOHt+nWIFpu2kuigi7Ouc4arXFFNvZY2jtvoOrA3HVnJnwv9V
FwmNJZLKxPtlgtjhFMr6I9m66wlnfNfk+iaFg0zSi0aan8zs5mft2qctOWFbMCVy
GCPHjfYTAtwt8n4LJHK1xpLbtsGDUdl9fevAp+M/k9GQG0Gz3K026cA0VeSnMoBG
kVxgGx+ZW7Tz3/7be8T9YJQm79b6v4zZfVXLb/NpHA7Ym/Ovj7G8CX5U/V1w03q5
jTNtnwg0nYBqupBudUZpE86+KEr2r41EjaaytNLAODSpsmAhxKGB260h88SJ/o/1
eXuXEXIiGbG4gQcrg37Y8a3xeEk3TI8glvP9XQ86KNSpL6apc0oIF8skewE2C+zJ
3WC5OEXaL3c2z/gwOKHOEVuR8YXvmEpnFjLhRED7IpMJxR7PFqjGFITHprROUhPw
HtivK5++dJrPFMi9dLTtRyPz+aazhznC/2IWN1v9yDiyFuoVYUqoLHp8/N//TlL4
MWpZAhXzLuexcQnuRrD+8MvJ8r6Yv6/oKm3Vm46uxAa3kQgNpMVC+s9Z05CI6NPI
563KA9lDF6PkCD3M3ZhZGSd+HeAkaqe7f73sLNrNw0495JmBsegegEiJ6kARjAGX
8DHNPSznoOAvFkjz04VhF45NEgrSh6IYAwj0818XG85EJ0aLqwA4fn4DTHEtZFGA
dOSiAw04ef4X1mwaLWCVnaORV0vh2t4DlPFQxT+NPAw89YtzTrOOoRynRb1qS61O
Ak8ERUozFxMwhQE2jgUknC4ko2Vz/n3+vVZ/r9IJJXABQwsbQnE1XDa24d4Mzd+1
EfNZncuQrU+F49LVXE/Ca95mKngdNqLIIIvIGqYkFr+H9oaZttaZjGvv4KK2W9fY
U9foDFNt3mG+t1SVhgqxV5KHuJa8O/KYk62zV6VKbD/Q+Zwi/1SG5XVEGu8vrTTk
3+gGV8P4sRB1WnCHjcJ+Vv55cDcKci1aZwSPQLiTc7wSUHaMmnrg9fZO/i844+L9
JKTEAtyrdO9EIWftk6l10hGSiXislRXg0Xhx+eEMNvYVltGZ0NFex+b6KL8EXJ6j
AtB5irQ1zINlw1vtjqT8gmnaVscrrhWn0xPZ7u7TBlafq7bqBr9KPLlhMTxiM2yn
FOdtfAUi5ApZ0O6MswUfXyZt4rc5DiyDYkpH917HW8ZEofJgnsYHNhlATVAgftKj
gDHKP/NLx5wbFZNtbDjQ8hoqylXc2iCzdKcY3cUofsM2QwSpkvGjkbFQ88GdwaF7
AbJ/og7yfKjRH4321KNqCsY/0+BQXdFdRlQF1TvZR5SkqTy6kAfbqjbSjmuwkHAG
n6Od6Ck1LkLVEJD1BphD4eO4COsm5Z1+ZoGeV4wB1CY+2uXJjCUkFSc9SUNaqplP
0n+nAuoevpwSOJaGy3d+uGdRHgAVMsMyoqPRB6Zs1mNgwPkuoY02lZjFBTfWSUlc
PUO6WTIXMn3KaNYc3qELaIDXjQKUJXtGrXmu034M0MC33slWhdmL1pqDqefK3Sug
85wX7Gb531VMQSFZOis6ynJRZJsfm9Uwvw/k4v/i2cyKZ1N2N4nMppgZj7kMZjoJ
jGJ7vVlGaK2LU/ioPxeyPAaFKEcNNaWTH7pztfY/xFeXHymrRtAY6dloLHi2J9/f
lBrZ/Ih0gKAN9Ao/O02MtBxae6qbUAwyykn3N4r6AKujsQpxt/9bD6G4jU/KFbaD
SETzj5n/xPcSPDIy9xJrHd9ryLOT+mtbuMP+12j5Bq782weSJlzAPRVP762Mjk5g
KWhSTROQgFoL1HjWIJ4HpHnMtqOJD+Jybk7jbwtWnCI/tEmqyDB+LbbSaSMQwziT
9e+0/TJalayCrEmjiKhTa79BiV7b8/HVfPl8fQbgE3jz/LISVnaURZI06bc8YuGV
PWHw9jKsQD20VjK15/wfeGoCh/y+E8B2txZjXD9vbDS8h6QqM5WMF8zonjhVnMDv
xndlKqydZE7TAysy1+LHucFLpVckjBnhzy8djlca/w7Qqe+iUkTaU6y6Bgy1nx4W
WZP1ZzXsLGUh5JfMzvIn9z1VylS01yg3y01zCkeZP2UmhOvbXOMNNUWqZa43B8/L
gMX93pSfjHdsfLRLhW6/i6N3+I8xReuxEF3slGyW+wdWnkeUY0TpiSZK6NxxgkQP
OxVdyZKuZLjo+DGTj48BV9teAnEoz4qgJj0K4L3p0D8frFUGzFaR3QIf9CQyzo82
tigEPEuR+KTfMyBJgS0qXzN+WQH5HBK6+9ngWeTRZCM5Hj6C2s3l+EfNz1NubSrZ
fnIQIF5H6Pu0rxsiEtLrQQ7fXxO3GsIK2WZ8pna8zoXB+TvU1tUNCYAOeUX7eyhP
j+Sdn7TCj7clx7MZ+N2i0V72WYDbhShx9CZ2uclxzmQYhC66o2RI2yd19x77Vqfc
GS422yBqwQO3sT4vKQbXbacbhtPgdz0zVsnul38m5YxaNWti7dJPFYHYRKzaL9pq
ovPsqttbzDlpq4Aor9qsyTkDHi9N4F8lv9z/fHTNkc05AE/n8O6o0Mu3HbZF1ogL
mrWeX4nMFWBol1pl8V8AvnhtsQWrbMXvvAvYMiFt5OVdNP2eNwTXcz6YfdP7u59B
Q8s2G0fB0xr7NR3uwFvVhYYLcm0p6x7h7fsBJ7SVLqbmld3pJBf8LoH9Zz5DDYQB
FvZs7Bg4N2kMnHQbOXL5R0VP/u1XOeHtN5aDbctxJhB6uZLQmB14R0CrGkLV3RNR
zxP/aDeQfwekNkFmtha0oev3dD4qC5POuFYeb8LVJo6XvmhcNMQGUX1a0MpRe+s+
gEbg0f4uHW+wU+gA3YMlU9RuediHIfCY7mElD6c2Gum/oR4hzazgR2RoZezD6mR4
m1b5Neh27y0WPjnUWiMxXl8wKkGVdklUlsdd7BuzQTWAZGt4LMv742LrbrUW8fvT
FXBFmjk8Hrwy2zF6HVn0/YMYC0/ceogHiVMtUFF/tEI3d4Vrd5zc9YJmm1vID4sR
tkjGC831QEWjDGwMRnOTx5iE3Zda6ggr0EHuEH+JoUOKESNl4IIyhhTwATmY/O5a
UJ+Nt0SNM4H7WnyDyjFwCADqIOTp7G42OHkLVQifLd+2w/zcBZFqfqbGZFJpmudu
XqifBPC3ICXQmQniXn5N6ylXqov/CPz8o/0rf21/rfEnFQ6dNW95Wu7cVNkM/BhB
v+MG+3HOy/9PX0vlRrf+nOz9iEaCWu4TLnvWl+v3G/98NHJuUuSdheQXd3t1CE3Z
2R1ps9hLv6I9+jPclFlJXGwDxFBCGsGdCOhETqHnQc0mPCZjiBY+5BjAgCf9qG5V
9lsF3y0pewn+Q0VO3r2YdPAJPDjOTnOvg0EGKfljFdn+5hxx4EMPmGPIUMRIgiz8
SSN0XPQPYHGjIIiffG9cYfx7ieJF0G2T1igrI/VXlr6ORgsdYuGU5qEkbjDmtiL9
Ca1MxaBguYcJNkGJsgo4g8uYAsyG75nuBiOW4Pwj1YMM9Z5kYmoD8sZY3RiROyOf
rgJngPezNgI1yrQWOiapP3y6j4iKzdC8Xrd0N64s4QbBTed+djZlS68ZEGCO4TkN
h60AyRbZxZfnYnf1d6X3hEaRpobpsiY1ucMIcuPpG2tSk2DVbcQd9APgasRpztg9
zZ9HXvdOfmqHv18NAGL/dh+vr2RFZ/zDOCLCXhm/1zrfSNV9cpcrpLh8yux+TaG6
I185j6NsqQm+6bw5o9GqbjtYQsbaJafn9/+oSaDDFUZNnIrhoPUjSJ76VmhOe5cF
dSsEwejYnqZqOzbMYrjTk6Gbev32in2+oixLeTrUslbEjR1MvD5IOAMzr5jmgTrb
yKnIvj0Fc9fw0wN59ibd0bsXkoWGp1ajq07V2dktqQJcPfMVyhg3pQVI0lXK/RJx
3K4GMVTzhJ20p/bqvLV2fSHhCvom0C0t05MomjU0bs8ezq52Xt/a4aSQCDNMgfH3
A+HOlST1fCmTyp5rT5dy6ys1FwFmSO3MUrjNiIN3CN/GSeOwZQSS15xk2dnk3DCL
JFeaG5hnx/JxEr6JJYj2zeO45gsEpGMYMtN5RrzVvStg5jtrYHf6amnx5jmh4zfl
a6sy5qkQFhMR1hxCa9BsksoYqhuIRaHqWpkWdVoElwAefW+pZS/qyEEvmAbrD2cb
fALNJxII8mDxrdm82saM4yAP75c5T9ujVnNMk+N6qY5QHHzUSqhU5VrTz93PJKcz
ww9nP9iYQaC68yZUPrclCBbs7cAUqMmt+57zxIQ/leRT2HRe2txcZqM90I3B2Sxx
KlXc9n2mmn5a/BMr25E6yPZYggmuyI8Ltk6TF9aYmy2eRe7LYSSze/i1Mr7C//5y
HyYvKuwCddvr8sFN06Elw3T+Ex+ZrY7JYsBTMUnOLK6OgRzerL+vvNYSGd3i3LIs
fYW7hnlO5MHUm1KoP4PplCRR9KLy69l10OjsnYx9dhBBSg4FcDswL8la8+IaLbvx
LDz9GvrIFuW/6nGrUTwimGci8QK+ST+JDCSxxqCk2IBJ7rUOF1s8RkvzYB8oO18v
fDv8JWDqX/w4kW8Kc+2/QIoJsV3XhwytEAUV7lnmAqOXozeDKNay/PLWFPY1SM3q
RVck17fhqX+Av2dUEMBxHdPHGhRhP/03DcXPIeoR/d8IFqUy3qXIeZDtrwwMWNR/
lVguJ/6BaSwTB1GQ0PwftZYaagOAKCJyLGPL0EHhgkMu37LdudCaZJHyZNYB1O8G
o4nmG5qvGDhGAGys90jvgqs6XlpFZ9sMOYgR36r5Vn1rX55Xh9Rgd/t2MkSbI/DP
9mFpndvNVyaa9z36x/kn0H5gUoc74m5PH+QWW5UgMc16hRqkrr/hkvKoCtjtCNW9
QD3RHfAGo4vNfnTPioRTd7P7VfBcir6Xjp5qu2/P8bW27uvAU+lEd1Rm7ZIQPWBo
/WVGrPYM4H5PAeYIVwrM/eqHm5o9Qj9Q9KR7b9W2F5BRMpH4yAIAXhC4vLVIs+DV
+nWZyqbyQ0um1eXCGl4T2atvKbxSa9SHVd45Lx/YBfvIe6qYHMYuxtUJ8vd8yMWH
weIdUb/QAxos6duPbYxGdWpRVlCvfnz1pg42OnYdcDE+1zGKTBO6RpVQ0VARti7v
nS9dhm1st+238DVojm8iCUtPOOVeJ52xRO8DIKsfMh+p14VhXG//xKcJb/qdPmBe
uXRrQaDXuEJ9X1MLV9h8wVrlLLFN+l7FUqmFRUszNzn9D6mZXFe+vxmPDegC/8ct
Ba0SjUC+xqVWDi+EWv6SO9Wdgan5zEM28p4bXr3lEUSOE36IXIoXx39jvdAslThi
pN9+ZZekOJXAwNaKPVQyQmYAHfzQRE1sJVQYzb5V1urmsU2Vv0yQPLJPr8OnDTlW
mGYztB93QEM+fK1YdZ1JAA1T9JcenLG/OLIgIe3r8b7stlhWwWfxXfwLQXDru5on
mhjxlTkhk008O3APBpzgpLsXi+UC8ApPsoWe1fX2oaiFkkKA+wWATZFRqm4JG/JE
E/iNVY1m9Yjffg7ItPATc2rfmvfb1vi36ZvoTpRyz4DvTM4bKLGM5USGr2NEfXIm
jrfafo1Yft67pVOKDmQRqKCBBTmN1tLhvTFrTQU68qog7gK/t0vqc4orPx81zztX
xLXSrchIl+VybrGbAFWi7tCYif8Kvhn3dG3fcuFzi9wDIUlvE7fp9LuNsXG5ROXr
c1QAQKnEUtFB0l+JsrGZitijvmGHP0KO4nILDB61TQdmcaosdgjPI5hR7RTklm8m
BZJCqIrWJO8tmqhDGUzPl2520qghL4hhPZ6CKg8tX+AeQ3g/ec4wRhPYDF17uSfH
8Z7GaURf1Xn6cmcOyR4ZoWVQJNytEtfdKm07ZmgdC0xaJpl1bZU6O3MuNCR0sLlT
YsC3coz/oju6Raptx36DV7YK6DnUzjmIhQj9u+9dax/jfbBXaal0M/h9RqCbwdMO
wYl92Dk3g3prggfRo7DWiv8hg+liqDQPeqrckrEPRyklp0gPUA9b2pSByjq7FBpE
dN+MoSzEMSSXbKmsGgU8ckMZ/5QVxqWyJA9mSBsNIVOg5llYGxbxsAv94coYKNzg
dVFIr5IfTS9KzNFNy+KGpmRzPmMjwOeds1Fwv/Ze+KOd5WkOinXfDgjR+ScxxG2T
27+EXJnTqy59KD+NS+DlwDtnsiBPc6ygVwUs9vXWUL46YkF8fXaxiVvBi4tGmRy0
mtM4R+a+B5pSNXtvqwKG8Fh9kWupsuX416n6BQ7o9RiGXjhg9YCciymTwT6pDj5E
NO9ZrPWAYLRX0PqvcqfH/Mjxlyl+ldXgBuICIq+o+zwuV8PpQJGg7TNAT1c+FqZE
jI/NmKyf2UnTBEhPTnMy+4iNg7onNcXpIq4Z5clonxbFD6VjnTnjqohQDlGQHeA/
Y0wJQRcK8JVNarrXgPYbHfX9Z8a8Y2Y0iC2Jalm0ZqdsjOpUKLB5wIvkJqKT04ty
+vv+u8lUTWDyQbQUR3KMfhVWzj+Od2MiGxmOBV6QaD0JWIRXV9AfUMRp1kQCjJK/
O/rteMdXOkDJagFf9+DTem+xOIkD14t6701PLH6vMqr5StE1GPAoVoyYiOHbKkiA
nQpHIkk45aC7Oyub4/AGmQrO44aEcywQHlU7IO4ZlCSUmkD8M45yW0y6BJtvrrCZ
YiRqU2phjcuw3BBMD04bDk27lMng7ab0xaRWWYAKXKZ80iHqglasz0QeOMiFEPZE
ecQkOiQwdCb0txenFk31z0czcas8dOCPykBQVUXwhtQ5c5G4qSqYa/M2a8SduKIj
v2oJohADrnA7m90NEc7K4Db05P/D0neHljFv5omP/CiqLp/k8FH1U84Ni/ZJorOs
nhBCvqsbb5UFg2YV5cia0wlpTIwCrYqLoQkRfKtg/Jbqef95orkkDwfGTWfNBMK1
7PNJNDz7sK8Zx4WQ2hZwtWa12GA+gl1rA6h/qS+6AYUskR7bvmlI36NVAofM2t6I
yfvcxrqG1n0jgey7JFJ+IL+s3rQuZOwbQtG+jTjqTYqwxpxN4yemcAq7Lixu9MOU
50fq7d4A27il3dM1JmVQFe7XS6UZ0Bkk8NwJG/JOh4JzIx2+pTkTsMg2BDHAVPbG
WPThK5vRqb1JkwwIjE994oN2WRyEtyW1NvFCEczWVs+I5Qw3R3s8sDJrua9dkHb5
2ox4tYNAWkii1NVRLQbjUu5YTyPfF6RI3PZ+7Vllv95hO3vJPZ4o+w0j6INbZamY
t2nFeRrUUuYn2j4wImWp41ouyFQwfHqXGL6aGq/1oHkiR8+eK2p223ePwgFtZan4
dWsYNWl42udrpAcivxYNbzvDP0Vi8GwyNqYq0n3f86KqYmIC33ZUHR1SHM0g+7yl
0EE7G6SevuCclWvDn/ul7VaOJYbw54i6p4pCXk0No2wZzHp+c3UjUaE4Gjc2H7yT
vTtu/g7rj7CrkEbBiHCqm3ZNIFk3sKjgQEhxEapqide7sOGpCYty++izhzaP/y/k
COHhfJrgpgrcmvwJAWObir7rYH8BGk84Asa/q6RoqIOsbJhaEjdaPLamTO52KxD2
EHOIIn6E+ZUrs15KajyQ+3kIu90uLs1IaVpFoY/Ct5CuYoMwGJF6DVSeEshmftQd
tAKMJ3GfAoCL99RpXKI8qSlJT/1r4D+jgSJ55rdMX5HEPKjh70el0x1MuZZClBSn
JY4fHY5euD5a+YZSG2ZWh0hftz69A9VVtykz3Pqi0dpAVZb2nsvChGUe4+PVU70b
CDIDn9CRTNqxJOsLFt/rtvFgqhYcMepqOqtvzsiy6xmzuDnw5Aj7ZRNVsgLNCAEW
zTIWJUncpUHBwQjpDhwOe+xWOPKPASEvKHnyAp6j1hDda5CbHvKpotvUFiEoafpb
9cVuFvmhbK8D7IWUpUZgj3ndBsAD4taKINUSBXV/niYvsXihpSpGgvwjxrPc/KnU
c0QrqdDB+VokZss+Thdbxql3KtxMOCMO6OzgNhu0nM5wF5+zGnDa+lL0JwHCN6SW
oG8qKaEgbKAYm2uKTs7aDnELOk/PnXljbsLPsVQgA/FBZLaCJp7jwzVdtBDu5dR+
mXwy+hZ/V6kN81J1m4bbdxKp4HfihsZKS8AVTK5OL0WG6nvwnu4+YBe7QRPeu9jX
SMKmDlMbldoFrcHOEfB7QG3JGGG6rDxaLQbiHOCyt4OKkW2jKLzRU5rCnE9RRito
DGpivlSwgmc0LfaLrRX5HQUVF8IWmAveOb9CVYkbWDwDdgeDb0wd04WjFUO55HZ5
eISJmA5X/XHMWY9qmfncerRINg3xlvt1AJmfR540zLkKOL7Lg6rH0tfiud1Up+52
A9lLPdsllgUl2Q12wBdM3NFSJGhtwQwKx6qQLSAG48yWcUbwGIzkoPYfV4FC1I+1
rIVa2+FothDf20LXoc7HUGow3ipZf9nA/tig/4OSVIiIQdWqiBMsx4g8tRECO6or
4K4x+VIld37OIVgg/Zi8nBR1lE+ei+BkyN6o5plqOXGfQEaBx/hxhJJkj/4HmGaB
0f7vLfwvUvTdM3LQV/JJUcczZUawPXk0tmiqjZMJNeM3K3RZSDcXY+jc7/HKEYNo
v44MYfp1vJrk+3++7eK791eJJvt4ppZv2D2BLoY/rU+nP1vc+nSG2WV5vUCPK/wH
jYI2ukvLii5C6WD2B3vkE84EfPi+/zsIMw9v9IxAb2jJ6E+A4gCmh0VCSc0AFTqW
m5c1saPd/C8vM6sSHEr7bXClVXAJo5dhE5IMeOMuWRJcKxW1AYYWGWklcXDgIWPc
wTY8kKRmbWSto0uUgFD12Ln8fmgKT5hkARMyuHCCmnFVziMgIFlRm9Sw/8HwYlWB
aAiGgvQcxtsv00PIK6gHOzY3E+xz/b4M0Yr2IhQPIj8nHhjbGKv51FKNdtkPFLUn
hwlS6iB25vAj3Fmg4Wg0EpHKpXXpBfA0ELIu5tt7HchudgP8DZYLRbZZA+9Mdcbd
MGm3iidm8veji8tVpAPWKKIP8WZvERXs7Jjbm8nd0/FoP+mRiQE76AEs1CRoZJPn
/AMqmxG+4GoR5JXdlPYXoX9EmtvmEN2upVWi8fgerOiUGRWvM1kJX030h4GuzbN5
g0l3BXCX7d+9Evm8nfVuQwH5jDMsT7znz6mBDKMirXOBL1jhkdxEZLL5FCIlxisu
Pyn+EV/rkwWMNbk1qFBwsXVdQ5Euj79kUAZK+/JyP6VKy575w8An7Bun4cr7Drn+
s5ioxo96E5Sx+8IrXsRDXJCpiObDt/CGzAaBqPnHwhnxCJIbuPzKUVoi12oZCKFl
qdM3xqeLjlzkXsXCBfTUADlw0OEiMRm5yV4DzLR/th4X4Tkx/zqI0VMtI74ezHan
g4GxpMALOcT306GWl0wy3DrOyTLfwQ2+wIgE/2qEiSU9dz6g+9IdLToMVrBJDo1O
rErce3Wd/U8P2OySff+HJZTwb2lDKGhOGaQR9vUK6SOsxIHZaAZaiOX1D90SyHKG
JNUhmXFEsiYi1Rj9PKm4EDCs7HzbMxNIS259IHGCjdqlgIoyrrh6cY3W9r3NfyzG
GBNDNTiarwLM/FYxVHZle/zjVg35VSoIyx1wy1sJA0d4813MizBwWioMnQ85BMuX
I7tQFvtqxzF96+efFB5h2uR6526Qcgxh++3N0hn9DOLJFJ7yjmZBnMNXGEByBhuC
txJEuoGgolRW1Sud9hz4T9Qj2Qxyt8Ri6y+rywi6TO9tdCNBAastUInnFYYyNhy3
0/tTNAR70tfTksnycvsuxm7n6Qf3ZaZMDcxZ2AdXwfHzHkxWSFOsvh6oJwWgRkHz
nSmn69ccK/8v2LCk8OBmE/DIJuE/Ldyi95oDRckQa1sByvwzrSTz/JZBBvH6v4Wg
z/RXyT1MRPZ4f2485GdhCRzogfkKhXJO84+8Ml+H/6hx+JTKAgFi+TrZtNWFBN5Z
eIs89iq5ezh3G3ARbsBATVAe9KQu1/ollYJxDf8ktyhPhyB/HTS00gp4kqFtFFOU
REpAPKSJPaP6VAaRrFo0MgSIQoVBYE732tDv8Mg4iHiCjlUhNexxF2230u3ndaTh
UOgbiGtJR/DNwBhE8p67mQ1RsBwqZeWLvmF6QI5GrnYCjgVmmpvzKCsuRKn5jZ0d
CAyVh1qU1Zni/WsMrGy/JCLcKC4IdTvtJj3HmDH74+/rwHVTszSf4/JJZFF+vnLn
XruT1V2e8Q3qQvZaCSO16zYWkZBmDY6XXgHjmhbRB1aKDVl8ICZR4U2t4egTtR8x
5Dr+W9fx/7Ob/usXsT619yW3Ir/W1y5DHKpNxBYB+E1rVLoPPEb/DRFUF9vStKRX
Da2GNjlBJAnZAzu3R+oZuuKQH23fQIfFmrezHv3r05zhkX8mjJcCW5hyp1SHaXgb
c5YG0Jv/BDJ9JZG//MaJ3x1zgHWxPW4nOF0/GEP3K/lqInr5u7CB9ucFZaJrBSDt
pfFHf4gCUdhB2loDfRsX6JIzGcKQ8GU7tny8iV1bMKm3sPgh9P/OPtb0w6N2erMC
l4kJgbF9DBNcLbyqdz2Qax9IzdRafAy6qOK6yyFq7ucg0N0Bck8p27B6GENXTdJj
dA4Ef29oymzpJVw8hTVirgCHTw7iIAWVNoKb5lLoxEARzBd9MZNaGy6WkH92LpzA
kLWK5niOizV8amQpZOAKpNwVpY9n3kAPKYCV89/DRGxnUJYX2iZ/ccaqvA7Kby9y
tBVP7domah2YiOEBtTEqnLKRN4nkkRnjC+Ubh/VBDo1axOt3UlNNjr90/cRcua4/
+kUH8MTOJLCi15DuuMxxuhSQPdF4ica0PUv2NNlrah4Fu3wJ9LpjBRV4ZtZpbasC
oAEvzEKsi9Zkp/3Swn3hiONtU5qyczhq62HtvXPi6F53nAE1b6xZUs2Mp0WrRo4f
AXd6UjH0Kp1kbuOfAEVqeSd96BlGC5M+D2ZsblUvih6eOnrVNK0675ePlpMUGvSn
d1sNsuBpUAThsIXarqSmp49Nkp1tYIS7cCJZ2roao8khPelCO4EIFo0Z0vsP3sfe
MDr3HxhgAGwuPMIUkJHxNCMTitSTdIiqAWaba5XfojW5A2Ez6mxibD1MwqN/Qj2b
GVjD3NXrvz+1eKqhjPh0kMznU7yXkR+HE25Z83h8jm6ArEC6UxWevpc/GBcwVJrl
jmQUUFOXV7rY20LFoZid7LtKV3WYTcsvzCEq8OCd+hiZWWuJ73TMjkaSxd2uxYsO
Yh6fDPqt8XTzpu4ejIryK3Mr9nKKOC0JIq7130ApINhAxw7kjmKcl5LX86nOypmU
MGEV+2tgZ+i995cMnJrI8FjtWwggwq3enxLKVcNO6T1/d3ovDC0LIQOCtSuoRg3h
zq2wVL3gMbLsXzd+eUEtAAwU34wLJmNjfZ2yGZx7LRytOXupKNYz2QBbx448T6HJ
cay97Jy07ZpqZZLrZ4ORgB3LD5HmOGk8NT9A0k/NqPQntzpiAt6DaD9qjYF6fvek
VHqI1xCu59l33CsCVgk2RIhoNcsn7iWk1wzBwX2AGQonOJH3rmP4ZizvM/5On0vR
XD0YMjy71ISRL2AxzxPfPIJJGbwuWOatA6yRcb1CSUtyY/Tt6iK5+6EsgpdMeJk9
/oyD2t7SSEGNPES/4gGhBYL3WUrrmFtM/H6wMCDe5JO4ZqiBs5+OG2FMghYIcvAH
5NAwCMZy4vJatFmXCB9v3uWgg3DxH53aJZxhHJ+zvot3omtOAJ7J6eOnx5fSISEc
9yAW9EyRSkayMJpXsJnvQAGkUd3nsxq0wF+fDcSNL6c2K6ukkly5l5nnNJM6DiRl
M5v6iZ291pYxXtOflME741yUyZDWC2Pc/ZQEDNDgzwCOCf9iYkiRHq2Q6OBT0qzY
KbC9518YMtwiNoRZDm5HDEAHcOpulmFcqKtX6tbtySWtNub16Dx21DYzzjTDSEy4
k06R/SuBcC28SDE66xTYTACynP1H1cpQH6Ee/7B2wIVfQovIXIEiyoClIGnRH8Il
2ymwnUUOV9Fojlg9ZE4sofvN8AiXXs6W9g0XTWKgoApHTsPhlfiSV9vlRGMzu2Zx
xkAw8rB/zL/LlFc9E8E0Jozxvno+OgPWF5YX5amTKzM793CTENu24Ta+jnj1FCuB
XaHlpdGQfDdvffLu+6vTEaJyKM257fDoxVd3OJR8062Z7oOmfMYud261RrWKjtae
fiC2bovScJHAzntgPmvtkhY3xjy0it4OHLazXvs1QgEjQatIjZjrRM0s6IpeApqF
WMPDHKwbGsLV8SA6sqoXJ+FK2pUiZGTfgX3Cv4k2ZZaazEylXRTF3AJZr3v5dwQl
+Eliz/zAunNv+wu9eV0lHKy0kKh6TIjBrOmPYAresOhLelNmmZhNiKGi7eL5dxSR
mpr8iBIRbN/dc+08Y9BfB2UzKmHsU7g6xzFCzRDomlxos3gWnPUJCmXx+To3DZ98
kleF25RnsgBu2D5f6yCtZjrw3o2aOMc7da5saqWKutTzK+Vo0yDUNbtaxgnHNSZn
vdWX4NvNR4OUo6OtimFIcitkmHzBijj8mps8g/+Su9USkwq9eOgv6se4lDFEPL6e
qWHR7RNIL0a9PaTWnLngqicLVHCUWpR4tr87ybjMfrP2Db4BtyD1qx/k4HoapGHM
3xqRNbu+YEY5NnWyIuuy2YCtb28pIFHRlq62EhOr1WRyE257O4OIgIC0iSQnC554
aCFbtG3E6mRsp42IRhskJvHlEL+WK+fIBC4ZFOWtJb89AVNX668BKLw/8jMshgCy
hoDlK1rrmb57nfWiS7MZFEdi8s6p8khr4mkOUhRrLUSeMTli3qhQ6gZLwnwXShmS
442xenqKlnOhEikfeRrvtewyflDs/AJbaQ1AQAHkGIaUbeCxvSP4CXIe12M3zZEt
hGBG6IQYjPsvag87O+GEyVtmfKrtlFFAFlzx6ENxYGh6eFYR18uPGHNMsuQ7J5Sa
aelNX62L/ys5j3nYy+cJFJ/3s5A9n8PAZazQEpx1u7NZA87v3c1Cd1YmSORgbgOe
mQmRblippE8n00aXItJDV0FXUOTFIeTGWlvtLUEW5ONCBoaxi+iLZDBS0nFMXQl7
tD0kQ7Koo238jMBw1L2TfLXfKOwp+bp3CN93HfAQITpI6twrKHFoeFqHVPtVo6+X
NRCpeciqKb8HzwmSO70LdYFMwhnNREoE8XT819yveWQsxRrS1BKIsqG2oTS//IeZ
r9+beQmEpppujWTHMf51S43ryNDzUUT9brrx4vlTgrrH1zmiAV2i/1KaOcIBnQ3d
M+JTtYOMt7jxeDjjkU1w0hRfaXueWsl9WQbj2CDV/c6b74nhCXqSDyJxkWPUUut0
WJkOL/MQKbToWklcoCKQAf3TUyj1VDmjQlCWqnCwe6hhhxWHGRf7Bdp/YJ0ROCF4
cyt9AtiXlyChvqNb5SuSMEV5ArLwH/XedRskE44qoqcQkRsJ7xGEUYEYS5CVeZZc
mHcO4wvwnGQ3Dsk58vI1cwH+FyQWkV/j/YARy3HU0jglYAXojmDmoswySwo7/aPs
ixYjxotEij4wn90YganzZV7fYOEw1eOLwMYbPqgHBvpHV9VBG6Zldp8T6032wi+L
auVpd7t0EL/PmuI6NbKUDRI770c73imkRvYEsuOIZ7C2EmjIdruunr02yBPlJmWY
FHukAukGQUYOwyz3jNmTLOTAMpteVHLkLVpekAGr6wMYfp6idkhYgUTVM6KJ5a7z
nDqhUqvWfTcTFnbUOlwrdbm97AC98wndGqsR8dIelG7f8ytEYJhqOIoLrxLmdQb3
YnTAfobzvPHFAN2UgpiNVBktv959SO9emMD5asWjK+hrfzjIUWkl1jlRCD4G0X/d
NJEeP1XfAljEA8jt+42UsVa7rl0nX4DzabVQHoxEDFfUaenfOoL/s3JgaEBjraW7
t9Yq7AzKs03+BAXH0ine7b0svsDcilskNjo+EiDCjzcTm+cN1HX5JcJ+ldg640L4
Sk6Sg51ji3+wJ4eu2Oc70o7EA7QrfcnkYtjPz5FQGCptbFqQ14HEHswmXlcswsnH
6Nt7u+NY5ZMPjRGlsgg7RZtZcGaEutWrgJPROvj2qj7Nh4fU71O0MchRtZHJ9y97
3tY1lkwnAce2onNa61+cP5dTGoAIrkDbDVsFwAmv2TMnmK45YiAQAY9egnr0FQj9
LAp0ZIai7m8RZnkFkDkCpv5L3WkWbRYbpIfzA4F62BdBVlS1JWcnAisAxT2lVe0e
MG+DabrvLjxdmVsURqSJY9eZu4qWJElWv2FU/HBodaDeG/BoVAVA/xFtmw7yZDui
M3r3N7+x+BX0YnJzp3l6SubJSWzrtdwJk60dFlqTSHSSksCL13lFebOf8F8nJv0M
6eX0/FCxsSJ04nwEbFAWZETWOMvg0PDbitPpUonFNIjYYAzkJ7sk41zFgqAcmP1K
zsI/lxUbi2VWNhu2fAWgIeEbh50Mn9wuz2qo4lHAoboH8wATDnIm6mksXGaXU9XG
1cKlfG6ieORmNpOpJ3xnW26wD3D3Xy6Q1oxPy8bRV4Xe6ZVNjxKMbezf7Z8NnPdz
ezi3yIRjLZkV7kiAqs+JztJU9BnrEHeCoIFBxE0ljmVB/QZnfnLRcC82rrCWb2lh
MIHMiau7qEZ6lz4t2h7IMo1JsVczd1J9E0LfpdDd0fDiZOU/5zPbsasapdshtqBJ
KjbzYaQ2wyV/AQ1HiU2Y782680zD+vW4IClVQ1Q1/o8sDU0mWDBLZmuysITpYFQm
ROjdqx2lJci3erFBFFOWxd3llJoBlspL647G/NfUjM7eFwO+T51/f6BYKWeKCDVR
ytVedSi2HSV8NvL4PX9t8OniT5pN7uz8Fwb19de+4ubtAAg0K6eK2qo+/19EJ0Ox
AbpSywZTmvBTfApvrmUnJ234yEd7zLADjufI/xRbxZIAivA9ZRXKerU9Qysw78x6
diDqbIIiasPDzG4hFpF1cKzUialqrshZ8PiVzYP9yOdrQTgLlRslG8Ew7Qi+gLMF
5Bwdqhmphf0P3E6+CbAbQLaD1NPtyLyChVdfhe+HA9mI98XMDWivJvXEynszYv+/
d3ol3wjV56OqFbGzQ5E0vJx1XHjZNJ0be1Hnik7uC4eKJck+G3CwOZIX13cz8Bxy
f/gimcyi+mijBGGdmjUcacieaOC1zqSwwaaBlZyjQTylKZFraImW8gYgbx+2gXsV
pNh/JGkm4xqaFbZhjk6WNgGlzTcAmXThcoeLKrtjOV0T4lTtbKUXw2Lvj4x984hR
Np9itq+g/J9/EGQ30t13pzNDbkCTYdcz/IEMR3S/isaeFUii0LiZN/BCq+pdKz52
J2TXfjKYn7U043d6MwR/ZZiHv6CGotyu1RqGYRuoQKF3gOGpKBz01Mlc22R4BKr2
XJ8tEVjudxKBLGhp/VS6Hp8HTAliPXYX13iLbJ/olSGHk8k+zQ6Wp5v2rfjD+Rkg
AOMl0U3os+IPvn2/ly9GPaM5EcDX2R7hU3o1pGxw8QA2GzW0mz0G0R55zLrfLjoP
xGlGDbAcRINIEpHWenIi6zMvWprWTtaFiYgd1GFLNOZ+6zKFZP6+xZnata3VBnIR
f6YZj7JW6qicn0pAWapOyQf4VVUCEimwns9jQuvxAnIeoGklSB1jNtKbu6Hu1mLL
JR0VF+Xa5lj+oOlOKKHWsdrFltdWYadBERmc9BP5CU1RRKHZuNUpVqWlAMfQSfli
cQfvmMH3OFcHLvVvNWtzmDd2kgNnevj42crtkP6VNYthCNgbxGUef4nY+Zv2kXFl
EN0lt/SxZJxEdOVg33wf53VeKsozkjOsEWZSQHX8LYMKvQLTgZJJL0ZANUi3r/Or
e70CaJ+Z0181+a1IY0XCh626pMi5EIn1as42kO2edH1yb73AvnlTLPBgNKPyHQfr
KTRQUbrMyDn/IsuG5/hXD7mc1GwaMSuWXtN9cXir8Q6AjzM9V5jTlowG6Rot039C
jNR8xJpjVKDBkYGzQ/lenJP+Pa0vEDasPEVFI2pEcQqTZMzF92b9L+lt56x9Tm//
3tNWeLs9Be2t2SE4HQAsA7tQVc9gFpUTPD6+fQ71THNv7uhhqDw7F97GzWJ/tVOE
nVNRzxShnfSfBTRobgJOhrelv2SbvqnI8SikqtbZVLAIYfHLOhckuYzsMidd6KUB
b4bbjkHoLI0Nmg3OzGyCgFwlrJG+Zc2FzGCGuKWcALcAi9dGXH1zAY9UrgzBJpKQ
VjOK1BNcScCYF93lIAY3yqupsJ8MlmlAQVx8f4G38vxLr8F5jQiNv5VJncBNSuKI
h0y3s05myLftlZYsX+mnvGmynvBS4BUBpGx6fhNPagQvZYxeLGD25JX1IUxxZ6mW
3B7dJkGz8pMHsLFOsFyAqGOc1cstNF/1m+o8EwI5KRbRz9IptkWg2e109HttAsxE
6pc5jdQCfKcxXkY65QqTHpQBQ6DmreYeaODROO+/Knxc+xKwJ8/VJeb6QLu7z1PY
RbZTv+kbD8m6aLb2tEyPV2nIDmZ1J2q6DhPVKi1ujRYkumuxrGiiQ0akjpCa9vOY
dkMg062CEThw/3Gqp04G01rHKtcNfz9/FMKzqUv/z1s97c6vzpb+X8TuGUTrOWcl
WmmznHu3sPCkz9ipSki8gui9DOGCweCl9v53lFYAbVbJqA1XP5FQdNjtXEbkizZd
fzcRtI1t62Ofoe4ZstVAfUKkonK/rx6hfssQ86SFwLlakcRISP3dHN0SB/jldtxa
pphm2nQqdWmpgcRPEuTZuT3wZrKN/26+dFBuFmOsFwAEPKsqeP+tzCwbfaW2YVYH
ESk1JurJPK8lxNDx1yCoEqRxQC+s7FkH/Se+NZ0T5H4YV2qdTmEDdO3uisC0V3Hi
q+vVdIZjsdWyOZSTy/JVD3cAiQXaZoXVL3/XZqyhu6TY3ghNx47EyQ5Nr3ADcVuF
m+nMgw0bPGmDtspvn3C3f0+TM9YRkw0HRkYZTCEsgQVkcQ4Hy+5fzbUeCErOXoh0
wSR8Qv62rIMzK/tS36HMrx0ERDRJ+ISAZgKd7y5480A9bR7ER+TD2dj3n95JnjNR
4HViBMkSxVY4EvGxFIrkXJUS0JyK4QTen66oOuKm+ZuNYbQt1cNfsroELEhd0TRP
yh0XC8SitYq9AgCSyYq18NC3Y11Fl5LBzlkezzvQbyQKn7j7sLX2jErW8VVL26bQ
LygryVReKvcM5VrWLHUGILOtiGEi6sYW5cAJJ9pIGYgtvRP/e7BXzguolOFbq36H
OZZvTzkb6qIgMpgGosRBR9WtMs41O6CNzkZvNKH9VoI3zFIAkCshwSnFxVRKudx4
4zV86TEWsqRW32l28XHmyfSPb2FCVuLqaVRGWStphBIhTWKI0dnWZxVfXN2aIK9u
g+Tjiq/OG+0JwUDaAxOjesiM5kOgUtbVW/Ej3CptFzPmsv6IpvjlHikKvQhe33j7
fJ2nzDCA4ESSM/etdF+CdH2rE0D6jjiZRsJF+UNDWHbz4tttQPpJcMVWinTbtABx
10740SAoasZ8ru7Q2VemnN4x7GoAJKSzFxPI4zBVnChXHJO/kFMXPNr4G/JK0Kxb
r9cGV7sVUPqMgZBShkHWW+8OVFGqOkTj26HInd+FuykM8VUEoLtMaofErh582hgd
2uH/t13TUyd+aYMJJ9Vr9QPpiH0E1Q5E6PEcvSv/6FwT1kXS4PxykEtOSinW2S/z
PSHYmFHgUCNNwYWNfCoJ4oqrHBnB+bjcPOfFbxq1cgDkU7CuVitzkNr7XDz+UITu
3KKai4kVTZv2VUuVgjmfibDoRT5IE7puGNaK3Y2we+hFfVtBZLnEuR9Ps69k0GNS
u24D6IuCGGLOx8VGKYuL0gRG6NMgh1UGMKfXWcLzxWzKF4jfd5lX/dkVbXjkUmtW
W//Ino3mo9tMKL+YjsZLniqUmFsVKsAZGfUsB4J/xDuDpz4YrMMd/wxA/TQ27KYf
j2oZNJHLFufEvibjAFqVkjLx1ojrZ9XGOaXPuJR7P+OIMl0ABAo3UMKcZlcRlOhL
667q5hvV0gnoZ57Wz2wF0iOVP/WpjJEQq9nAObgOVXpQFT/NR/2vc9bJ2JF8So4y
98BtOoWJ9rEJWYxyTiZBunWr3t92BbTv9Vwv7YQlciG9DdTstWk/EqKXBn4pqJKe
OMWVCFq74cerLIRE2ir2Ot6ofipEf09F9JoZT2DHBKVtkBf/VrB6IVgWQTpTC8tv
g3qZUPtc50R98XLIcXyFh4zy44hR3nQUz3v3klKuvA6xnf2voP58cwCSJgfch4MU
IFkV1L/7wXgY/TsWLpT/aT3RZQ+HC5CBlXK4/YjzRUjxyL5jGo8mfekDvLjJe2w5
EIJUdOe+fEV9SP+eUxnbO78EfUNrEC56NRRwQJgd7cQJB3IaNzVhPj0ZFFpFIYUU
DXWgRHuNh47IaBGOKnGYG0ZOh+AlBnJSR0LmJBNQ3h/X5jC8MMRSYOMzLdRkKni3
6QoRwigHRbz7KeVZCw31V/Y34xzWenGpiLOgWjQ0LqZozDmgP5tPYjKQy4/kkY31
we9Ww0ITsZH1o2ukS9DE8EVuBQjkWhAwsU9ekvEVNCbCMhppDOjig2mvpYryVAIr
i4bUhSzwxn3urxZkehbnLLx4pBy+SOZ1MDM8IPWwRlyyFVb9jxGJqbKc7UqAbFyi
0EgnU0jmKYGqvPO/6E/wtb6f6K9MIreK+0KV1AWMtKCKGbEQYlrqjjRZJwSzuk3p
6DqPdo4tDpT1bmGTIsDeReEBkR+kfodlrjO3afd3ILB3fC67pQcXLXU95Uv3+e0e
16T2AQOdpalaM6glo5hlEpNWs+/4qhdkC+nJkREeeecXywQpwdP+iwkX4DX/Tdet
0hpGOv34GmvXS4uV0I6loaA2zrmuaDcnC+keKp+5Sk7lwxxBSVmLoHEfH3selqw3
IZ9lMxMy6e2T4WOC/EUAkX+JN6d6gsmOXWCqmCVY0cP6p84MjFzC/mAAuCbZbfsU
pkZ3fCZZ1L1FnsqMK6J3YQFYdDyy+VtkevR5iUCVf+VLZePHVmiLXijqHGW8CpAJ
DT6cYvhSRS6/GVgtxXSN9GRH87Or9Cfc95qRcdflRz/VUOu+Lkh2uRit8TsIJOMa
NFKidIqwuYrDOTHlnTEH483mixRUu+otJnV6FctM70H/0rOzrGwxvAYhVhtiIiqm
OgGv5Svx4JMSvnSqhsIBpdNXNOCTOry8C0lE701HcBD7vXCdP/z+i/+BzKVyJ2xL
9awWpLh3HyFNWL9NZMrhoJ2qsRzUkIAM/dRRSbnOEz3xICynPcb8WohGPuwfzl88
CR3Z5B8Uev2KZL+cXM+KwjAGBhcgGAO0YPh2ULMq6JWw2jJ4zvSF5wdXC1BCvASD
VxVMGQXCA5LS9KvIeTqWMqLp+ljL64GphgTSnEVlq8uFhvhLGgAE1LbcgqkJneGC
7HSCw0NU6V4mvLkJZ9SGa47YoYqxGCzhMeogtM+YRHZU7O0uNkuzdo4yKrOyqFm8
jqz+pmKQaVEaum9fGUGidVwqVbStoSOeVeqEGLBlOacQJ7O4HwNH90HeMlRzg53R
M0+BpHggV0OVEbwvGGYh5ZaqpvpA2JtGfm8sri/ACkaNgGivXPQeYndVdfyZClIm
GlK/YmOJGB1UXyyqz/zxyFi0F6YUTlr0lbEBKcGpo+deW7ecZcd12TNkjNRoETk/
vs+zNWMDlMQqz6dgUqX26yZKAMowwlTgQSg2Ao7FfYf8IVRfq86rqq9KLx4IhNSt
xif3PABOYR4ETVc87BIzHnALyZRNvUbEinSFJsKLbNlc6K2Di48DrQ6wYCM1VtJk
/AFsnSlH1Hhc/r9npZRz6F9BbZAvX9W3AqluoNa1XaDPZwVKIORisvEzuh5C2+mK
JUbtk+LFY5czsakQb3SlYWp5tv64TrjGzZpUgtx4q0ZpBxRop7++CoE6AHnzmG2h
9GKM9H+/BYzWB0TdWoCD6xEA3vAIrgoIZmxmvMMrJi5k1gh3/ZkTKj3k0VwT03le
wNVwpU/LiZ94A7N3V9F9vFa7LSAhQhghWd6cd2BIOnOXHs1r05sqK6pRiA9YgzOY
GCZlUdi+KnU3GjA0neaXkmCTbcAyCubyvNi5LQH1y6ZE67g+pJUqFSUb/dhdBcrh
AB0ygMDbGomjBFojsiyqff0PkFfvKzpRxu+faiAgKetaBI9dEMxtTYFIMUGHbdhN
8kxgKIJxnqEGILrK7ftmYAOxclVDBRgewf+HL2IFhJ5RuoJF0h7mWRNjTz8d4p/e
mRDnS68/sN+SNOIjlULVhteert5OqYAvh8hDh52cTEJP6T2I/r+da8mcXtlhaqNB
MV2yVT+EG8Gw09NIwBMXfO2BrTbIctyoBKRwgfeIAzQ3MtNWIlsjNoLToKc+518y
TKr+MIbQDLExp7nN7DQDgfsvqsRhlMXzSiOh9GKtK4neIYjdqOp70OkyzTLTBKLe
MwvZibyh7OqAxzN/Aa/ygfzUos0Y6cWD7SKYrA9P758JdjK5wjppVDdjN43iDzh+
DFkqN4glFpQBfOPmy9fMVItybO3D5Vop6+5i8jCGU6saG0hCiw9A9ZWnzXlOIeni
RnB4JKNNJ0LIcakzp9VVElWNP+DCCPw5rndjpx9pKGpguIDymlfUg3tbhWlxgTpz
EIqe66e1XN4quh4ktHwbAlpxR/pP7xrHvmAT5kJ9Bqkk/TG2jEFa3gAK2zIBNVEQ
L9VdsIV3BFYZLXnAOU1xkovQuNtP6h+yENb/I9MF99TygdO6FNgurVaZmhrU9cJW
v2P8+lhQzqY6g1vokyvOuVlftTBhX+pOfGo+7PxxI2XK8sd8EIaOkI60InsZQC2L
l5Bb95Ael7UY3WoPMCmQcsBXv7EpVOIB3D0bnl8DvJyVPeL7U1wmbdUgNrGbEosn
x22pJdr1CitrrhQCDSFbm6/ZSKIGl5J3Jt7DGBGswMz8mZ+N2y136glUkGMioLuJ
y6Xdfo1IjamiklORYDsh64QkiL8bf/8TlUw6jei2Pl2jYKrN5I3sIq9Se9GV9nKS
K/p8nvHUwBf6u9Cd/uE0RcrmeHFY7bECm0u8sLlsXeAkHsHc0+g94JWjIO6XgN5k
3LEcoxSKOruXEArJYf4RwvNG1kgNGR7kciVJyrsmdqFqIxPtxXvhiCUKyucsVsbX
gvVZXjbBVR63WvOvoKMOAm9NOEE18Kg8FZZaSmWP3Rnb6iBjJClH9F0yLEbVl+it
tmsxpXhGVNd7Qojz5K6qqvymedTXJqaCPLBy9lfAoLNPBY5ipJm/GmT8iGhA/NS0
fsCuGWG9yrt/0fDyR4lB35r/cdv8PycfW1SWmres4HXuBqK9aaztj17k9iqjXfYq
E8CQFxqp03Y0YPKeIPtPlmxdQbk2dPU6O7U+AmLoM+2jd3V7LvQ3jV9dRwB9aT4h
PVJ9Kztr1pq3qmuuglw7tT+ezRCc8D0solGR7shfEw8uYdB2DFP+aCNlkPRW6Fyu
hPgUFXHgjOKLKz2ClwwEuEYlfkKyjWoSYhd+pw+eapSAa4SbojBJiY4DhI/P8Cmx
NwkBIVFKrWIiIuogBZcFMdy3KVR7Ar9d00DuyWPDhUouwtf1tR7Et0B8myCdHCsq
XAtI1JEgnMzwC9Xy4YgnN4ZkgQsPTVDLUutRAjtyY1ZgZozg7k/2ry/UsAHHJQt3
1nLEaxs8HRrPLzAkuCkvlcy0r22JqT1Raewc+yodxzDHnxsRS4D4kqOVtJOGvta1
JOxZ+kM22tLbMrtGJJHFrfdQp4KJM4926dGka+2uO2ABhmwAaLt8D8P4yabhv+m+
fF7MKPKos9ZNq5o4KFrvIIkPYapZE1bLWSSwHb1pyw2zjsH2Ooh88UXh6s32O2G/
CcLtlxpJOe3af2p82EJmX4c2xnWPIP6fY26BfdpIVhhB/Zxo6V2swtmQcYc8r2Qi
HDYcGfNNGO9GsO8WhJzmom5bxC7mpil22x9h6SyL9LUscuIwVzIkp/H2wYy/kUsB
brZrQger+N1dgeVkDSlSCMBBKbrfpuBAXfUVWnfvLB/lBy+7iuR28//v6alavyK5
1nKl25qL6zLpojGcN4lSHg+rW09MI6SHSDbKrmzTJMeAfWgvO5lubrx77XIgt67b
bLYlFaRlwIDp39llvrqC3Bi8dTWXXMcMbLRJ3Zm73pw5o2PJ3C+tu05JCYO8USZy
zBvrcJsjFLsgS8uvIHxCEDlPbhpwMqSnQUYaf9H65PiV+ODjmALUzQw+jH9hvro2
ZeWvsWTvDx7x987dTh5GrXfwikFPsz09BAAHRsOYe2NtKeS2y6aWoLzx49uuAlBI
MsPVdW1/CL3kNB6f5j38PjKKWgD1oAwH5yKp+GzZJjiTZ+uzjymqD+tShbADdF+z
x86Ms/MJl4LYWd1EMvsYWXn4JwRjU5vH1ZRjVhYLUW7IZUcPytA5BP557Xd56qpS
+klImcAg70xyLgLZodPQFO5dvnPlnXj9wpqe1pS6+AVrTyYmqTx3VLlXldTbpmo5
3lUGwM8HYERvFbIhx9tFn6Vi7H06spYfsg8p7mCemm32tFNWNjkFRuYbHzJZBuNk
G6Tp6xILeOOR3yEfTFD4N6ktJTtHR+duCd2yaxPCLzQguhzhy4rnIXyffssoDUpk
j+QHe09A0/LW6BB47HY3ApX+DAAKPsAQkQzWTWUD6mvib7X18ewO5wUz0Ob2nSIh
YsUEkYNwv+rnkzae5Q0fM23MA2GQEv9m1QD1DL39VRDtEvRyMHcunebIw5XG6W/3
UpEcMZDHXeLFtJ4I/rQc0FPYOOwsJc29DmT6IpaDjFZr+TmHWgwO/ynb5JX0bdQZ
pL53B1ez6fAf4cffPHp6w0Zx25wLdwrTqpjLnGn8OZgedpwBjVcFYLs5e25cm9g3
esxJtGvE3gSWsoVPCUh4mEsaZ7V/JTfhbWDrPJ4nyS8SHsRcS/V11zQVt38/PUuz
rLchqPT3EqI96MNflOYizAuwCvu3QiBHFDqoCsWSnqv7Avnjc+iRWlQP+60NoLbE
BZtUhQ9veIkOevZg2+rqcKPmpZXybTDEVUIK1ueb9kh2zycb8obKqEVReUFhPFM3
W0YYS07FsCU0Mc6Q91OzUpGYT4u6C2PzbogvmiTrXMotLlpmIqVfeXohxBBVZWGY
4c223XcFOOsOYp4KdvDPY7tlI95UQr/xFHoiHMf4YTO2fGZJTvLacHQI7EP8GOkh
EMQY6ldsjETD0nROHac7fKxCdxV1RM8EQ1pQp/a4h1cHNZQ+Z3wPBCHGVjGwe0+2
ig+HVVlS4u1ANU67CbMdnRb4PhntoZgLOOKG9uQSawt00e8S6jGUT1nLaMq+9n9a
4x7fblx4WzynWmdW9bHDfcp1tjyvN40hOdGGCa7Zk97ueQJtpGfwHsl+STcbWYUD
Jlw5CccnfbajzPkt5MlKrgomA7+i3Qau1/xPTXCCsmA4T0ldISEsBtqs0pBP76Li
+WI0yNqrchpz12YvhtiX2Hqz0RSwFx6t76WYZM6kMAVx5n8ST4GMgo4YQeb3QcHC
b9xP3edKEv6drGSdvP0FTalwNn6VXRGteqKeBSgrkaOka9yL+ZkKyZDN+Vg0T7cw
l2WpYDjoQwPlVotcrGPwl9JNzGED9E2zmUBQTJkfkC//RDc+5E5gpi1Svv7/420t
k1nfR8j/ZzSLzH2ltY0G5S0S26IaKuAfq7juBlpw8yTyeYdBh4KXuTar4C2xmPcm
g4CugmixqqP9jBTtBWOsaFbISUebgiRruKT2BgLbeonI1aXHkq5EBvJZ+HgcpU8a
UeDw6X97bDk0UehvjTq3xvEQSjwj5KsvvHUxVnPUcm6Ir/8G2NLx8CTISUoDRVg9
VYeyBUAfu0PlXfHWZhuqxJHjFFrDiLK7kCw9Xtn/1Yeggp/cYik8UPad4Q6ux+Vr
TtLokT0D5E2v532fJW5pVugP+IoBtv28x0dkBzMBOcbctSAurb+aes1bA/EujG1F
5bxCv1nH7h+pL8jpibApp6hsui61WXm7vlPQcClb0XlQSATIqrAjVaw36un3tfsN
Gv0iBQRoDod9JDv83Pn+5pwDydoRFbbsC0YNRiMDXsKc0voGmrYtEtO7oxRKHALk
wal8HzD7AjJivqEY/DfoUvTI5CeG30wCxW2p9ibDLb6MkRmYpJfyYfQ2N42tRdRt
4r0tj9Css9MQGhS5foQEfiqURyO0CPkQVggAaDo00yWmBvkZ+URUbHeeumfOMK6N
R2xAHP1XrKr5fXzv1/v5SslvNumwprQ462EuKsRuvJ8olHfwwajlhGrsaSnvJPbg
GOOVjwgt8O90XiGeg8O/sOfEMOa3k7hDzY0r4ejNOcZryGn+Fo85/jGydVd2lQA2
jecx6OE5UADWInxc7GnFpgILPq9mB+tx906ZyNrxrk4Adaud5Nd+kcCHRAQn2Be5
2MDxnpczMzxuTKrlkNiHNrxXFnx693dyMxDpXWbynwpsEMcljPwwL+l6OiJu/lHX
PETsKQ/ntMN7sTAk6nR8m2SREXVsnVM7oImUiJCpoEKwRQWNdlhroRMa28rkr6pM
ZjHa8dmxlpBRqCknWc9aXwaWtMEA6Qo1yFeBcMBCLoTZ26mlpcZGkoN8LL6OESTp
jHhHf7DYh1vXPBSND12kmWH5+0lsPoRQuRloUOAZNkoH13Y2tHUuLzLcO7jFEkdQ
zXhiX06WtkBgSjbtgp+mIFSNwYeu17gpm+Z2o1PAfhBPk3HXR9JPgwJO0FV4qrzB
Nhs4YmW+hZ6YKU5s8GDHbKfLpk2NPv3AkYTnf4rfr98Rot+R4GqvfU5+2KgsFx6j
b03cJoUdamIhZ1aSolsZmTq2PaCAHsh7sb/heGIoRphlpJ/bsy4DuBJDiCa3fuyP
YHPw3fCZjhXI4GHq3Fiv5eussHAYErd4fgTjB28k/XBhNjumD6zviEJcf62LZoqB
gAsQdNTw7gt3saf7IQIWqrZI94ozP8JwDJ9P9DPZHq+Ol0AKEUpBJQwBEBistXoX
HAn4xk/gdzkBTOC/YOG/61ve4Xg9nDQhN2IrWlJE94eWpHCrt6PxEIFg1NnzeocR
sfjhyhMuKiYlAq/6KZfYe6S+wECO2+DUiaKIuQFr7xjmNW/3C06RAtv0XyavQEDi
20yECxv0fM1oKIkjfsSznu3RS8oXjRsSs1WYfGXoE3xg1HZEEmfUAEzNsKNLPQod
uZ61vCEkp4A3KolNQl6JcZpZlORGWbQzh/yWkMFPjrU5CJQtqGU5cHH5ybBik8Qy
lF7CHX9H2bKX9TlPQplvmkV+E0lviazkfE2g8jfs+fIcGilxSdVFPhwQMsuiWM/g
2NVOJhMPTI0KP8Cbe5+9lcLLaaTkbqDrqR5F6gq2TX3gYL/tRuGomY08wOqokgiy
bGa4+vq65O6ECpQWHBbukvjmFaJ99inDAMPH2nlBTtnzmch1R4dpJmlN6z36X2BE
q3VTrXxdyXxKBdyaKlfu/u+e8dnNpClHqy/hHZ9RrQ03xf7r/iJkUqNpYbA2JfMo
nzHQkju88Uz/y9c9BivOHnCNcBHAxSN1ZquijEKjmSqHV6h/iXMut5TGoyzzbHEq
pI/b6hIq3LqMkAycCOgL2YJkCjoXKqyJG3FuqBaI+Z5bgJpZxuX5BdEqSE6O5PLS
zGqYT3/9TMdmYGYrjHctFE9PM3mwWNz1tKUXOKFXFDMR7+mjlvjqHHv2Cn+J/JyN
1kLGZrA9iBpv8KEhc0GwIu7M+UW3sBmeBDxmooCx8oGu2YDa9SE5pNMn/U+EVH8r
Z/VWQvXFRy+24eRoLCgnTU6KuEqsEJjcOiiO7AwQWmJjGCZgOOJamMhicNRz6JW1
Y5Ks6gbJTJR8s3WIEY598L4zMYax5Vow3+g8Qw3PG/ToSn1JaDKwFIJeEaSWVJ9j
4suRm93FhxFRanZmhF1d11rk308FhUYViv7gWQkAiqbHkLt+f4tx+je6UgWDLBuL
VAqNfeeJlHoXi3A60LHIdfUxTrGwrnYolag9TIO56VBMMkHcK/60SZfxE7faTuga
S5T7S0LPACTAN5//5BJDoMVC6pWIzgI3d8k1qqglTZ/HuS9x6Uc9eetOmmrrkX+6
zEf092G29K1/ILpKnJCaFmG7TTsb4JCa8cvTLnzFLRF0tc+l3X+uW5KE1JTWILZX
2wvjpWg8Zj2DeTnSTZxd8UPt6sQy6ecGx8o7jmDC1e6YcU3SXboUbunkYJ7tYNk+
7r4daPgXGJxcmWOrDytEzWYJGIilufurt8len3dXRcjQ4LSS5KDonBpOxsqPvwMj
Cuu+DJEMjoF1a5/0v3VKKZBkfwklHvBpeBueJ3e7idlgA/uo0XrOD9GExEvxKgvX
90um7mBoO/eNoGGh6+/VuATirMHtMDSbiwsS0oqdJ7UUmpFhAaJW3RTes/kELshB
6JtTpzwhJ9acFL+FP1P06XbtELVeA7jvimoVnZDuAqoRy3rFzgVuLXdq7BL591Ti
Sh5UzcYdat7iMCnzzLm/KyT8gOTNrKGo+Dkme9FakPZt261OOEYG+4LbGQRJLYma
oCtWl9WAYEQP0vgWZdQA5XWcx7FMog7xRYDjO7oaBT2SGD7iK7KmvW7D/GUVNZuh
+VaCdyeJmOmUBS0XABspD8ecRj0W/Trt0707bv1wlWaQozbLPfmb1NqEuvNxf2fK
b7yf4/KsgfkaoFfcfQwtKFbIEy2wjbHT6sL0PzVeDMoz3G4PBp5olkM/YvP9eUyv
4NyOi3rZtvIHQ0hMn3kNlbh0xXmouAKmTvRk+9ppo7vzixe5QSOwmL3xtjqoNHsK
wvUetMfSkCXTKdfojFnSfV5AXffIAp9+2gAUfyGighFYZ4/oYcgJZ6zSh1YrLAfe
ISVwntKSH70AYGqOSRXNLXgUgYrI6VQzvY/hldNNIiO5hoW3Bmj5UcuUwxpQrI70
WY94YzhCiSKe51xZDNkcVfIaUBpfQ/fX9rNTtpmHvDGqCPXYwepuIMuexNo2fl9W
W2qsln18bKy6KbmH3rhLCACnC0bNQmjJu9IMqu2acsC/HNJn051Nz2iznt38DMdq
k0+lRXHtFamDZuyZEHV639zyC40xVgK4e2FM8/r94Xf7k7XOLJNdf2R/wSI126VE
+CbpvArs0lVl+mYqPoaHZa+YALbj9aoYDAp/o0N0FhIBnIGwqMI5ct6bFv+QQiI/
zyqRFnRZKkc9nUh7KilwkMHl12wV9Q1kNHjo+pI7rs/t5585nWa7u1xFYt4ROf1k
dqw3PjG+QKYMAT3nVOKYeWF5vVYghtky7X4fluVaqwypeXhwvTQQX6kkZ2Q7v9/K
d/vCrmW8WOrTvBdWuLSRPUZUx1LpjCTEpnuzMaD3g5FFMuuleDNtI3aLHZiA+JWG
kPQ1LAnj8Zk0f48txbV1puMPozMPB+Mv9rjdjzZ9YaNtR0UaztuEBVG5/ewkvuS5
8rGNhY57SQSMVlmvx/uhimAn66pBAYbQ7A5QNLYJXwno2PROMO6o9iFnTmPdjA6E
J4Pt8uIaPD9P6E5YR8U96vTc5P6GDv7Y8DrOd1zjWz/3GVb5OaECS7henRDm2+4h
IRdLPZ6dMGmZ0EPkw2FpdVJoqowDpX9OW90huEt6vQFUWvOk5h5Glsi7kUMDJmlL
rVOF4KmV6uavFsTzfMiM9zVbFEq1MTZlpQ+aYLkfDnC6W7FhdfiZ2ZN6b+YPwcIq
mdvnpkYY72t0WX1I9zNlN5I1dhMO9+KcEE8cN6mFsJq/1gIVTIv7xe7QCqcuWcXR
cNTosk45UWab8HIoG6QdsZl8FFd+F16yrCJ4XBjTyM4zFBPsPYPoSnaD2avu4hoG
zBdkie4Cm1T5+tY6i5FAuzckVSIl37f+KHS76gqjaezZzfIRVejDk/p6mWmvro+b
DfVJlZ9e5/qwO+99v3J8FJhWyU4jzTqkzYe294WJiIugIG19phmmU/kX5J6loPCD
1W/f1ceO/s8hLLJqCNGW2EaESYZMbOkLWOCMCPDdCd4SjGVQGMoc+R2CcFPpXUnQ
RjBSaKlrDkIiQULCXdpJBI2+erY4J83s6DFnGKw8FJszXqxTXUFuYxH7d5NyJril
T0jyMxtNntlaE1reSVf60stPVyRPs1ls47go/q92yKBIuDxBXL9vJsf4B2jHeFpX
KVrv5uStkEd7+E33FqiY5wKaU54GRwTHcUHuNPzm77ZwB3LyB8K5xV9eUlPt7Kou
uCC52g1ZdzqP94QWzB9O+TQ97DQ/GSwcBOlzxi7SGJoOabvNCOIMeIkoxCPMnWmq
HJPd5BbjVz4Z1AZ965xCiDEanr/cOMRJjkE5q2peXiUjD7ZUowRZMK8BaaYBqGJb
+hwHDRz2XvgxuNe9btJhcG6oO+RLgXZ9SiSTsHExGqIMR3dTt/4nIOyeZq6yeeOL
tbD0qGSF3Gbc+yMHx+veRfVhQrJpImEEj46qu2qxj25T1oE9dezRqUOy4gP/PsUA
5QhboQ7g65fmXAqhn+T6qqzoliv9B6BMAN8Tj1zyNMhtEt5pPc6TuHf96b6S/oj1
1l5dhjObIR0J26MJWPMB4qq9LRBl8yn9uH+V3tMzllpTjyhar3U3tt/bV0MlT9ug
oyhVD4pAfkjye7owOnrmtPHiHc2SZ5jbKKqQD/UY+fXa/IB/qDGDelrv27ocQhAC
P/ADWIv0foiePu0CWKLWgP3OJG0wll08W4q9hVVKL42ZkZ9XhmM1/mvNf2HLgTx0
I21p/+HH/LXETS99PUtJmryCulLg7jBz2OTd6izd2ZD6CNZRQR8/eXutmafn7DNl
A4AS41aZV1zRB+czVdmr5wj8qAyCrtE9hS2eph8KitvCGBxlbZvcWpnwG9nJJh3F
0QyBUFjnl5QxqzwMnFd9OiYev8erUFfv8V0DPa1DN3bD96ZUCqNqyMLM3gWzj7TO
AbhdfDZZgi4CWgjUqX6YZXlTvoTwh0gD8LoZY5JBETPryXw2S9WZs7YyIn7pv4yf
zPdBPjobBpH3M/FkTryF3H1HX+jYdb5z/pGktTlsXHUsuEo/gBts4G5htLg1Q6bz
Q+UWer+S4a3Fk6UUpLfWTu3RgPWulvnoHUbKViM8yMIALX5zEuYBXf3R02ha2YPd
kcGu3FcinaZiU+AeDL4euPHW7D/rvHdBJbwZuQTyA3drbC5VKnOHaL9SoT7Pagow
ZYCBS4nTznbnxU1I0BNwxvKGwOcpdAcgeRavTsMUd1oSUKJnJV1PSV+3Fv7uChJT
MK+SC1NcxsvjL6dQDMeO+DUDQWRtC8pgB2J9GCivwIU6+xP0qJOpiudjPNw0eTWk
sZd7HEcOWL4YkozgmMrD1wW+czPcqonRCP6EGUTnRy8ijxYzk8NKZhuionvDHvDF
wlt/ak7MpGCvToARtsY7tuklmZyFzZTV0cJ92d0ZP5cnIgIXoH/meR461AI65i8x
aCPaCyvhCtslZG97/8+FQDZ2v0uW68QHarR6ezOwmW0FUMeD1vB35uDORcIUtrhp
fdOUPDu0BcFmUgqtpoh4kzQUIyArcZOS8to+txwDfFk8W5X1MuX+fp2qggfyqxK3
iEAcm6bk7U4/4WSATAWViXlvt0NYc4NEM6+IRHWyucuPMBWjfXYN3ipg/T9EO9Xu
IXt4HXwicQo4QqJNP9ycN+BgCUHhXERAG2MUc9kSr/WAKW7kxP0IcV1Zl7kbQBoL
tZFBhNJHtoA7cw3VADPi98DJRQxg8Z5S/FicO/0aFz99EmNUgCCW6v5MMsaKuoUa
nGrL3z6xnOPd2KAxujl52tKYI3FswGZjA0ouORB/+JfeP9EM75UP7VfeDJ9mIlZ0
LEv9SmPOsQqyiV/VTEq8hnoyQWM60cyUnv8bGItKMJTtgQXy4/3jNA2sAQjrZ8Bu
4l+cL2zoGIJPBcyG/KuFuIH9MOLw+3ets5TWdnnqcburi0NFD4wU1hAKi9OmA+vT
rv+ZehgSm/Y9hCcdh0fb9lSr9+9xV7nX1qjBegEVa6FC6JPZCQkdX3sqKJNE5ZBN
YxcpNYLtnD3UNCdoAl5L4QUoeI8dYWCHEW5VXhBd6tl5mGvp7nyrIdojr5ZxmdbC
+n6BZ4rQ1FxE3zZWVr8rVYilw4q/UCDj6Y1b6XixHRF0h+z67IKNwlwPBR2JBmt7
IVGJXStUm1PB6XQqi4y78vP9FGaW30OEUzUAUoGk+k/Qj3viVOjOfLw8p54+Itt1
vlQi8zsjZ4LIyxNqqsjQp9J+94DisF1utY4pU02uQbuBqcPejli7T1UZILETIH1A
HKiqPTm3Z4eVT7sGLFE0jd7p4GeXpydFmGWOx+qEBjjrovTb3esQwo0E2U0bCkcx
IwRL9a2JuM1KNJbhqzOPKveAQ5DB06vVWNdQ/iGXJucUkBAHfsuUqcwRcUIAYnSe
jySJIrGd1vFPDBu/7jfNTbmaRg8ahzfwFhyf2MBpPI/GDhaa9nuwKIAOaXuNXZQl
tJE+c/OncdnhvIUb2nM3EtX08PkCkXpgEDPcfiqxcWVGw1r08HZgvOv2yX0n5074
d7d1PHLMmPI9w9J+j9nMuQrI928cziWuxU3MeLK3gUImNHmSGwh36RJm+CAlIypG
6B9hP9O/u0KQEedfwSArzLbSK8+ncIoTbuPBdrN9VDBrDHXpWqvs6d7EU7wPoXJv
QwA1DS7CXicGGOPfTcS2bDAWlyZYbvxAa7BInph8ADL7viG0bIb7QJa1tdSw3oMx
Yg9NllTBfEB17axr/1u4spvGxaMixsUQMuw0aLeh2DKJ118Yw6hM1KC/lBEOv28u
Ogy8vgLr74yupXH89vdLDZZ9fj/WEpS0kpcqumfDAiNY5Xhh3AkTLJ7hBpWAfNsR
SsetfPUp8dt/ETtddRrejKaa47QHa7o1fM2oswXRayQVKnIUXojlMj7k7SOxXwJw
mDraMClWPYM+V/VDp/OwbAUNmwIgsbGl8il8TZb9NV+mcz5KHTyEd+mnBD1nRYGV
jZycAU/WMyA/DG6o/OJiggwLNgCknEBZ+brvIMlyK+4WoONEGKLYm6sZlBQ9pvZy
f2XTKUJNc9Rgu9xa+QL7lRAf5e06rtcnSi1tBJUr6c7GcJkWELbRqYrXJ7Lb1UXX
G3EzpblkhBl1ytqbF2CSG4o2S35sz8pYXZp04ALrAJdeQmrpynMdaCHvp4kynw/n
7aIuwZfNsLODv7vbNy9xWHn/5FA4iZezh9TkJI/DIl+b1flAwRCQXm+FNVEOREw+
wdbCuOOImHpQxXfmF+WXYoD4FST3W1SyWCEwbBFab/RZV856Xo8NbuvULhkqiktD
2gO5A7eSqpNcdx/idv5vH2z6cOAKK0caWzgC/4iYAFfUJTVjg9rerM+Nc+w8ZX37
qOquPoUhPD9Mio4J3NNmtt8Otd1hk4HK/XSHJGa3ov+Rv4AaB+m54Sf7jxAHArGk
bfwTaoye2gzO0Su4UnoTd7/z0BFPD0byWJkmCEkZarc4xz0tjRqwxrUK02b3sn1X
n4VqpNaWr8htCXGJXTAiyKGPGnl4LtwvCPjYYymJvOGzdLLGT7x0xsIuKVm1PGtX
ufqo3F9vK9LAT/UHg6te5WsnHYJ5Y+foGKhY4EFgc00dlGBiXvlJIZUuyA4xIQMD
Ztly9M3hYTHwk8Chxz3Lo2rKFbw7wIFB1/J9ggOBrEPqautLBaWm+dbBjb9zER7M
PZ/5rNbr0zmHkBXiknDXM4M60o5aFiOiXl/T8GwHjjcOsEXCIhGQzFtGgY20x/Lz
mFNxc+DW6nDj2Vu4PUY+/RXGheU1mDTPavQHNdpeQkKX/IEwU7c19IM/0ju4/qYc
Ty3MAMCbMflY3+2DiNJX2vzS7k7Z5Tu5hsO4xWDTFFirFA9bE5gA/C+GSqXgI5uE
YQRGrDKaEIPD+cHhMcu12C+SNzZAbzyynNH/lqeUrJdgvvMBzFvG5oNJqNvEyzwC
Qae1B8/BluyoAMMBa/sxB37QPJ6N1FTOzFmNf1ABuDZYZarmkhdd2EsO9bi4ooMs
LRyd5Mw5EdZaRuWVixGZtIY5Mv6XLZRR3g8mrRy0VssV39MgQKEhKf/rQZIBqvU0
7OyUYdysXPtPnuGaNIJUsuNJs1vfWhNf7t4ieYUdGGitYLi9r/rJwX71pIYMzo0J
us9sB281rRRoDbQ24AlWgI5PQeuvVGF08FKwkB3CUmtwZKLegEp577gBHNl3p7s7
LtkQmf+J53cjZzyMAgPP+9i9HfUqj3FbBuROMOobptY6wt+vEzs3dY2aBj8haBYc
n7Iy2SwnkL4KPEPeLpcmRVvF+776+nIQWbJDbBnykw8d4mkfQT5axSlDXdfSXVZd
XgnDWo6piLBKA1oYz7+69M9fNjGQleZomOsHegAvxFLZmp/WOWRD3c2J06qFr7XF
mUxnoDgrL3xGqiNS1u5IiPUjAGq7VXoLCW0ypn4tLkDGVmpk0W52nN5Z7zih+mR3
iuHSvfhAGncJxdbU3DUgyaitDEO51WLn7VFTX/8XognjPWaS+Jq+mtNvmjpUR+BA
S0fLyAIe6J5CuaDl9b9lqg7P9hMfnyXHvOOa2RAmnmYMUin+z5fmcL50NJQ5bzPE
TRftPc7TzRJ7FGapEegrlLVHOzlWHDvnJ5BrsZU4ARFNR39RD0BeNTVLy2nuJDuX
W3QRC0YwXv02uCLCWwOgytyaSzNrWQ73QaNAVYLbFuxf9B19LmAfJHwxzLVMGUxl
bV129oDPqVywXYO9HtnDiwHG6v3kkYD9SJ+bWS8SfFTq+r5X081T6Jzps8WqDz18
+l3zkFlCgCach4/r2dHbpxI/t+QbBibfV/G0B/JpuiM2liuqA3rYUXxLJwolVL39
FNUTzLxHdBdxNJQEosCFanDwz/nPAVuzx7e215OrwPagdfckOm9e2z3g8bSKnO56
B7oBYYozNZdaLl74Vtt4zcSowf6W3ZXmT9fkgG0SOql0aQJJHLldfK1gqRtek6Vy
Ywh42rAdYsgGSwKbKgKLTsXrTk16hMKj8pxZoGfRc0aH/Lsx2hH4iVIx7WL1CePe
e++KecBLzCd4bL3V+m3rH2qT4QJ76C/Bh7SPn8wNhqeewGngZNzTJhhqa2NggQjK
GP9WjI7QDazgzc9qUyuIxSYJYNktX6CR8UhgsCf/h/XaTZJKgSMbMn0eRbibIn/j
8K9gcrZgCHPHs9FI93q4b3iNu+ur722QPqFqRYLAqMstTJlF+FQKJ966iS11rj5+
s0AlLLELiISnJ2H0c3XkLIUF+2BXDYhxeXkRX3+Ms5gWXpsmOewwTYdY8GCd+j6M
ieZ0NXGs39qwUyzaYi6tXqao9mxOZGSC+1ydcSQr5VWW3OFAD4J8YxrYYrCXnuDf
gATTTtKbtWDkLhUl6R0lKOCn2Smsg+VU3TCcIHRQy0g8TET0zXS8btR0ykzAJ5mD
w+PNEW4BOQSaRSqPYNHZr9ImSJUzotGhU6xIJppxoAlrOsoICG6v2s1+Kq+ZH2wF
3B4VAoxq7P8+PEcUxqKVXkvqc1riPqVZ2ZRi554M8+bhE/HZLIZAJVvqH/OfRNyo
8pbUsF9Herx4LrcR2BrOQuOV39F8CFcUzTykyENt9ckJlbO2vhm/EVker2p9drLg
0BSVwbegQmwYPYJ1ma5l3TEe2UrnMep+zzUSGB6RiMzeOPjn+q57S1o7xGpm3ZLi
R1MxF1sQP7EUrtwCaFo4BA9OuKMsa7qRSWTJYWkzbZ75NwIDuzVN2qT4Uzq7Kuz3
Ag0rIVH1jKafgIFZYK3Auh4JVTpm+XS3Ur7iREb+s/c2GaIax4DZ+5PsaMy84g/w
xegAkeEt8SDzRtyOn0i/AQbIBuqMR76JjVeDY3Ic2coxLIQe7mjayp1EYc9bTN7A
MySPOXRL4MW+qzzEJYl0/Qk4+RHAk92wEQjZLpGbjbrPgJWUVReZt/JRrAqAQWTL
7qlEqhGxbDEdRK26NqRe/7+PzQ0qZVyBmaznbjIGjfeS7tDCxdrxR5eemT9vO8RT
rKH4kWluZjmO11VwiA4yV92ducS9FcOsBnHV9dEXFBjXDn5d1H8POFdkTr3EiS7p
HIktQdGAB30bS0pz6wf8IdhBKQmIdyVuKvd/KCGrcbCUgQVAr/ifceobRVz5lQCN
S0+3ATpMSjoR34/PmF4VZRA4Tq0+mLoLb+S2DQvWHE85we6pqLwxBSTYbVqcjUXM
E/CKI0dgmkP00YPnzhFWmWoh29KWX/U//rEKWlavNCQpBHZNfslRqi09B3oTWCSf
s+FHsaROKGZSJBg9zyRhjU9928iNirQwrtCl5zAJb9EbDs3Im0FErb2pbah7mF7P
bA3hMf3TLXHW+oE6/7O6zH1RNyJypSsu52a/ul3Ev/e4mR9RD5hI6FfWvvQLIeQG
G6ZhCU1HymPBflEBmI8nTMouPX0Irt8tyMxL9yusRkf/GqcZsgupT6wFWObkLqTC
oYdKC2/scDmcc8zB6qr3PYHNSKxjijPI6HBPEq2NmnzpNx84tmH383tDVLREu0DI
waAHToM4zJ3VL5xr+hQFGPHcQ99hN7SAWkvq9VZxLaJmEA/ds7FQBC62dWZnZV2D
B6FnZ03UxijpXUUmMt7C4PcrDxITB21uatOXqNuoXgHQK7cFWUui5FfbGBfZlIun
RBg8UGLGr/08HMunrbmhL76uhPMkt5gWHK3Fbwtz8oDqDBM9tphZKwLf2QXWRzi4
XKhWvHt23hIvYTsxrpEFOKLzaJK4R3ltadvYED+5mD7Nrc9MZCCHLxnXvWRQAUGv
uR9CH44zzFPDOoie1WAj7XODuB4HQsZv5f+t6DDFtrGYcvDZTFeZWXe1v6a7JKRy
P/v2DhPpsVBlc0PldQELfFSz17uUYcNe2QCVGmH0vldg1z4Ra5D1MZpFx9rorlIJ
yycbgm3ae6XM3XE/fTl5MVB27X3kfoxmdDmoDBl5fQ4AC3Ld90R4EPHohy2cG+La
Gu06YNoLTRrqwx4J4WRQSveAcWvoaVYdcAkj5fumpgFVbCONXqq8xhWwK5Zju9r9
e0ddwHOWt24g3f54g6ydWakBeUHn8jiHE7t9/deLZbIudl72lx/1tkTfC1+qROx1
rGy9iRz4xmfAZ51pw7ZcylON58JuQnkxP4Z75GqRCGGnHIz5cS4WGBvjAJfR0VSj
2ieGu+H+DxErNCk1Z6NMzsIsfmiCmJGcGhx2Ybw31G148WrLFPCTLtIs+mw0a5c9
sRE89IbVhuXzMnpLXaPpUAcTB6okrpBPm2uLRpbAMILbZYxjZBaBKmC57hGlC+Tr
ENZ+2LDscOs/DJtQ3V5uaX3sn+lVPtN/4kL8+hDzn+L3a51nTkkMiqxx5UiCtKm2
wRq8xumqjzZdLYRFtCA5jn7IkIuUSMckcnL6eifCSasNUKPgv+KSxLS+xuJ1lRkm
ffGymXOQnZLIUABngfnLjyQHKX+Xvj8L3fsr7RgPXIF8pwhMiJ5lcFobnQto6xKJ
gZ9C1vMe9EuXf+EHeeZvBAlnNb8H24s6neae91I6K3bngMm9RoKrXX46si91RzTl
HwQZR2My7AcitrTpI+qpIV4TiF1DH8cRLyFJtimbIIu/VEUZXo2rJ2+mBkR0Uji4
SnKCQyqbT/+RCK7KXrTPOxhkNMnFv5SuCLP8xL8D2Q9e1V1j0wKJQVKNJZ7VWOfa
lG54q39otoBQpSAMVSyIgGkZNEZgd/yMWcqbWf3RU9VO7YzhEXvF7u71kFAdndJ/
bBLGZflikn5yGCS1sQrMWW+4jmgaX9eq6RxuOKog1DbIj2w+uAvDYowDvFc8acVP
W/n0eAOTnt5fX5u+xn9Hl13Ull7yrszUzVPxO6Ix4sINK1DqkYrhkXBwEInhe3c+
OZ6uyBK9m35iq7lWQ+rqCzVbFYCENxkYQK5fr3Zl6/cjxwO3CxFZdQCtvzczNRPg
d0c8xDUjRqoVxBRydwnvb/Hn/2uwVRCvOAurkZ2cMi9kug8nnKt4RNGKOD0YjbFy
h5XeMTYc+ZC5CsMYN9ucxT/Ilqe2edmzNxQPYeM3U+NnqcK4IwieSWuVyRknnCqb
tmrl4Seoo0rTjFhHb6aE08luxH9gDHUwQS1NpPDTzdml6JXRR6OrbpntBxedtf+m
knqjljqPh0eVzbZjZXZhM+ZNEr8bL+cpFxvsTsqn4/xX6nGCx0NFC1olhHv0Ecl7
j85HWjGGNbl8rS9Ys4M8gnugZSVJHlTb1mrI1B7pEhYECotNZM9BeAUb1mJjx28L
9Pge1q/wPW5Z8e6ZhgJGFgBT77kDM9EDhyfux4TxTRLM8nJQdgmuvk9QpaxP+Ri3
ORMLu7z4cfCftCd/nh0YixcoVtrsqlBtxDqvK5a5Opiq7mVSOZDJ/RLthX9C7duU
AapKjFdfmhdCeNwgCN4zEQdPSgf1f7wCcvyzTbOghWOi5lnu6w46JAEJ5ISHptI2
7YPGE1yD3R2cQKVMaPPXJ5RmTaZT7p8jSC/lS9ZSVOBx/PfO1C8su5r9NHrLG6n8
DLO/Az+LK1SroB87a2KFT7MaFkBRXVhymN4iCwuvBOhyQhvMPji/GUmUG+KyV/C4
XUXRtbWJ2azRNZFmz5VY5dJSiK6t4w8IAUA3mkwP7bR9txgSRvp/nxUEe2++n9v2
1dz76h8QmiWwMWytorHgjc5M40qkPWpxQW/ukskBxgogbyNPsM4NKI8YGF+WO9Rg
8Vt3dag6Ke/Bp5yXyKEMpvVZGGD8B3YP8KOj2iTThQfXqaXEzm9Fg1AkxT8ORNSo
3LW9jtn5Gp2QiBil7h7mEpDx10J6i+/PV8XC+0Qd1edP8HXl8oadF57uwzJisn/Q
hJWVsohV+/Iqw9oiZc/lSAQXp0BmuFD2IAkSUkQI+TIvZq3aCWc5v6ABJ3go/1Gq
lAbZkULPAXJ/QKY2fgnrOlHEQ0x4fp0W7BtZS0dd+Frlx0Hr7AKsNnZaJcsEjelL
2haSa8SoO2Ovy5wFUE8yA5HeZONOs6j2kYGE0JT8D6Yf4EoIGGO3aR+af2d3RE94
DLE2mnUs88DzTEpjfQ5j/kwma96m3cIS7de1CRMlekeB9eLvgl5kK59I3+Sfj5oM
VLBnjtsveVVA9DdnEghk53ZPbTgGTvtAnNPb8tmoi1tpxeDTRvMpsPfTcUown0od
+f30oRCNMzs4fKvGkGSd0IlpAT8CGw8AWA2a85z/ysQ3NB3nVzz1j1Wwupwb+mXc
9bJeWEU++kMjChzPFOHf+057E/jm1bCWs2RWNeXxS+WIx9MOkpnLF9fu85WrK8so
+z7f/qVIjzdJPMrzOk5i5WbQ4mr9rkdJO8ZFAkGhoxnt257dQdukReTjC3cuSjtp
lCW9e84v1g6DabRBZYPRW03w9RozgzlPdU3oKjwApXMb01NNnHfv+U3whPpxBDUE
QPK+iWpy2BMgWz1XkG49ZIxbofXLIZsHMwbvFF/v/sBmh0pcFaSCGXxMC5ai+41a
6md20tKEiHdoJUmgj/Ko2p6pkW+WSqFy+GTOByiQGpZ8Ct/eC1ETsYQZNFOKJ9IE
vnBsB36NChJFcfP45p5s3V0mo/yBfs8+cfJeV6o2Um9FvHAmtxsqbt6wexPdgRHC
IMjsvR7Fhsk6sAewvL4I4xzyoV0iFnjrytCSHrwwg4CPetzgrsYCf//iUp246t5d
JrPK5aJNPKO+/tRnRi7L54bROJAFKeTLATyVF09dEi6SmTD8kB/ejq6/YPkwjN6B
NZ3FA4W2eL2+y47o7WrpQmpHy5AFg6Bcvrz1nziGNHiq7F8jJ7zEpSdf5WlCt3pN
qTgO75WqrI3RYAiSSW4jA7v0AlnVSq99QbIW0LcOI4vMS3dOWD1KC1BzxWVAL5Te
JG0A+zIi6RnB74QH79NUZ3Y82njovC2/a0PHbkBcRwr0olKdaBSrrmtODm67vxTf
eFnyGVon4uxGc6NJERdkfDkg8W21F6/c0qHoqOoGuMbmVzTg0fQhxMSB+o5obPf+
nE1wXRvmfOdji7LUL8AJQV4Brebb93m7Ks9XlR2+roupdsucukxvWu38Dm25ye4+
nq/9HSLdAXRP1FmUyBmA0EiB7uD8vcaEh1OrZhLwXhNj5FkLSUEan7kFOijylm/1
/h1GTL/WX6s/DXey75RcwC7/Izm4z07spqhY6Wfz2Zq62QU8YGLiLh8E69Z4ULA9
owDfO+LSI8rzvWw7YksEabaBxz368m7fld7XTQmUfldnLhHO0EneivcYJwSGBSdm
x1xkS8fFdYfYhzAfa5oJ9RIk6SJpGOFygizeQINaf+nyWJrhwKBR808GzHycVA10
vb4ZuEIMnd/MSZ6r4KkyzXvgCrbpY48UYtO1YnhBcNjSAnhhiMKlw28X3fro/vT0
4MK0nXxlIFSUVLILiG/SFvgTMqXa8xxwKdinNdVPTbTReus4QoiZtchE1ZVVH3oR
CPTemyPBvBjDfHWwr0Fz609Xq4WlBm2lKSHM8uofDsYgb4m2C15d6bhScOptrzDY
+NUwUfpCD7s55FVZPawl5hhI+RNGODEEi2uFH4weWUtf99rc1bx371OicxkKispZ
G/kRJ1QzCG3nCJuyOS2kqHYWcGFZzrrjGjj/7lYQ0Crv8P9u8WTQ9O3amkJDQXrY
P9sESV7mbJw/E93nNWgF97JszQsX7s/XkjDR3HDm15bKdQLYMyf6U6NCi5U5JcKz
t2k4dxxVd9fq8hKUArqnQVpfm9KBmT3Bj1XpFsebUaqVTLjA+19ZMyTuIj3/kDsq
3aNapc5+QaQxXFo8bdvenU2/ry8xeOF2yONbcqRvhL4YRFnSUFEa4znfpM9Vg0ls
kzZgo78TUm6mN1kYOdRQXs/AGM0Z4dW7RJQ86ld5/jqDfvxeWzuWjKlmap0HgMmC
R1yfGB+iDSyhzXqoAdRgU3IVFfOxFSNpmzhqrNMxy2p9BsHoLFyUJt9E1lLOOEEQ
IB8LR4z8/HhAfCrMtlRtDHjZ2oUoibjBIhNOVDmTOim46AYqHi6NwvYVpiSX9rZ9
vaAeePnyzuX3aIG66cQrMK9O/zPP65pLyT8sLIPxV8Jc6gSupt3g8zD7MtIS6Ift
XVFtWTwUeKPIHZVQDAO1kK4v+WpfrmmsO0hAPNR382mLqL43A14r7YqN5Tk49VVy
nybNq9aqXwjmzlWdAw1c/Wl7WNpMSve5gFwsTGlHiRyGKkO8XqLb+QjyJ/2kN/gS
c60XRZRclgfaZjfCqmmz3KLvVh87hh1l9E/aw3ph58AVyn8ED3JBFelx32uO4E/z
p8WKNmodSomJeRLLu7oxYxaGbIl9GfXX3MXHDJgiX6wLjG3d206F0s+OiAjn8fA7
F8fXY5Z1hKOgA+OG5SqSLaRi6/Di3ukyY356U9De6bj7QUAcAPeQKConLqA6a1Tq
fnwwDrFtxo3AGFkPUA9/TMyLkdvcS7zo2MW0GjsuzIsSh39+nySovR1yFfyAcyyi
b6lbpvD7ditn1q3a5dHoq/XLiSZvOxG59YOznZhL2UrAZTfVaLA9FrwyLNtrDpY/
VkQr8S7AntLbuv8NJb66gyp3xQhTM59S5uxyoUVt5qPyCZ1rv08TEA0FufiKBWh2
tFWqJProQeVRnkFh4uGIcHDJG0+olHPo+kOMvER+8YUJ5813j4X3i6ECGqIhKgXS
g/VVuu6eeTSzWOFbKEmRm12Gn6LQMWYMFbiuHDlsIVrlRdyYPg2G9b2ApLWTjNlu
MEaBAa5pb4ePTEQFijfFpAd4m1nYlrR/P+9z2KgLFU5ZObnRuWUa67Mvt5aMDSWS
JE3GSaFnJwmFqZRyHzdfTfLGm3GuVNxwQI7Qg7sh2ovZ5GzSVVV8MkVoPThrLXRO
GOXelDTGC41/c8zbiNU+b28dv/Iy17krrYegrr4ePTzBnS1LQ4iCpBZURfP5EkFV
03UR+TMpHvjzcNK8RkzhbaW3lkyV7ej2mI2fKckLsOZxS8h8bmIx+QO3/oZv0sz+
7radkQa6Nv/cNDtheRxzvcvRbWQeNDNkVKEn4Rbv5iuLAMc6nWdl7SKR2NijhXo2
DvVcV/mPXAAI0qlD95SPX0eArN/XHfL/teeJttHMnuqzhz3gB4+OBLfjpMnIaYg7
YVzrgBd/WRDzcAkuSD7Uo13D8ybKymzZ4IgrofvuJ2gTyNYWXl18LNUfDB5v9rLo
+riakU1Vc2YcZbDE91qwwwC7BFqyajsbJ5p8K1ATS/rkI01qhRY/j06uVBb4Oeoz
FaT0u1TYJ7wFjwkgMcFZjIs+Ts3TF5Gqz0b8iy8PTK0CidsXcdR29AknHPB7c8Q/
7e3MkjHiumUpMFSjZOjzw4ZdEo+jMCJSmVtrf5DPLx6RMwlhwV7Qs+OpAbDIJyfk
YlS38a+XD49aJbwN+LLD3GtORL11T1oulx4nlbyahHnN1pG2UW6knXR9cJjXMpwq
rFAmtgzlBo08HuBxSSFYELpV4MD3VtWRZNArUxIghYiz3bSBoxS1VgAsrayjdhN6
xGfHHjrxR8qAR+QR4IXqQxT0y3QmjRQ7XZDBVZBlx9Znu/3l4Q3fsEpOwH89/R4/
hPIpjc3ziiFISAxORfjnXg4PE33I29CtvVksGOSCK3wMw275fnghvymeM3UTPUIQ
vy3LOaYu9Z40UB0pdGosgaoGt3miHgKfR9IXpH+zt4uHH9ONiCxlrPfaZvSsa8mE
12Zo87cGb8mdYAquPfcJd6Vt1QN7Dx5txwk40E7Ncg0NCQqSqYCMzLkkduU46uw9
gUJ4DEgLnaQUQcR/iwHpapduENLLF1XJgMVrd0Fyl9z7feYicsD56q0IJiLFDJvn
d/VASz2xCBqLfYvtUuBb7cCXcYkcwjs9EvggcAOnNwAaKYRta3qhXU+L3BOmUv0j
4SKFFW+71YGTC6BfppwnIrhO5V9/NFUcudWiU/MLT7hTxAIFfMcyDACtwg749m5J
I7Qwgtm5I+lfSMXVqiZnW/mQ1raOZoTH7QrWa9Mdz1+oPubCd1qGU9V54jlzHY7z
J5h924L/KKs9gYTscUse5nPHAq1nPQ/sJ9iQJi7ELToqroO4rCqYojr6ilWZG4wn
0NHJdoXycPZ+jzJr2KNpwxcv12E4H/qGiXcMGXIRVbzDWTCvs+YAaOa9ZllBoWwi
OyrX1xQ3vgEMOgqN7FPM3xTCfLwjo6YmSCX8yuo+CzC269YZXsD5DfL2l0Ak2NNK
j6L6Am0qym5EY3Ez0WR77sxXxHxPgDDZ7mhI2pXh3Wdzma6NSr9/ObbBx5n4DROe
oCF9GyKAWPNq4lmRbZou1SymRMi+HqUnwlqYRg9gsurxStgMZzKMnVveVUJ9yFtf
OmD1A8mEkFzVdsPqtB7bveF8NAAthdLc2cP1DICNlAs4iATv94L/pYNL0iyRTO3h
g328sjCVeuNHcxWK5vQw2qB/QS9yUAFiyP1mgMvIsUndj39sv/1meDqsu6m4eOPm
iplBfwKRBszrZ4nFfdIeliwc5LkJbxki9rW7bk40ZGv/VtcLlZ+CSKzb4qxM20A9
h3OBfJpZyaHQH5BjFB5RoKIYaEM+2L8hL6FlxFJUxHNi6i3AnmzHratDPkSkNtcP
0zO+YnrIdp8DpOIM1qNw0DlchLCRnmRnGXOV0psJIh1peg174xa5LW2PZNYS9Bul
bN1qUj+zMtvA3vFg0/GPHVF5x6pteGlCnqbCddxrzWxvzirA0xyxSAtgUR/HRNx7
PfeHScVmjBH8rxEmGiJlmRsk4oJSXut/GaDeqXNpX+u8zFG0BZ6crrk8zt507v3r
+3OF6oo1FzE/oMMHfQJmpijFVglXLuaaapfhUoP5QRD2qme1sbMZh7VpEd2gYfBe
at1xeni4BOcyVtvutT3ykxUzTcetjPG/acQzRpDWSPgR3xRKr5k4Rcnj+jhW4KmW
MrK72f5i2ZpgE3hI+TtXRJKrjyJVGifI6JN2hN7oDsoU2wvF/AsPtZACeZysMsA8
JMnTagNF7NcAb4pcJ6VKm/bQlKMG4M35YusUMBspAmg6Cxc4NEG81muGTFPHcxzy
XEh/scWM9qZpktvKTihzxcAbvrcpqF6Ja/dLJQ/qsT+G+VBCig8e2bGD8aHyCcQO
XuPqOcAzekFkA5cyKyXh+R3KrRuwvxAwHut378qll85uAJfUjLVTWM9eSe3671/k
wLs53Av9NJDzRhK6CNyBrNAItv7nwEw0d+DFPimu4fxFsIYAdB+BhANX0uLVlIq0
tod7TMLQ+nTaddnxUnxXOL96HnX661aqNVif3g1s+zUXizL2Do4h7LLXWH1t0awW
tHEEbOVQu10bibdIpCq4fUHXmzD2gYDiGGkem3VsOj3K/yC75NKJ7G457XV1looC
DdwtH7cerfqef9T1jyHDUo06doQm31h/vwh8s3tyUCPr80e8WAvVeOMQH3Uwm7ED
65VgikVAxWhDVN1OWTXbaUhCRONThIH/S1wyTNdDU8SQX0d3V/FpXoSweAJOBlLl
xxS+EszlQHIL2drLgI6xXR32aKH0m1xIoRfXYiUOJmXAsGlNcWlQVJanj7C9N7sB
ktdBeasoS4n2uMrX5bejjXjuJpf9Z0Il78ZWfD2zMbM3dUQWBUWoIiWQ3iF/tdct
uoTVoMkm+4tSnErDcZAFbLHrGYrzaidvAzBrlxkgtfWyH8MNKACLJXT2jLzMzmEn
UU6DW6vlBZF+2+f8pKt5pqLNv7Lt4tEeApM4A5ACyaeV/LD52Qy8/mVYnRm8AZxD
TcppBo+IUPOAHsWaeNIzOxBcJFEhZ4saqgRUfgc4NuKO5xDhL3ab1kZWuxOT5ZOd
t8MpZuguAaQK0OTfb0lecC3xFdzIssXIFY3DV8W1iR91VCA15rugOYi3CC8x2bXI
HPErwuVEW8UqNPG3Zve6DyjQXU0WpZdt43dyKXxazPDWTQwFg1uQQWX8O7UhGQgX
qjuPS+m3PzSUd/4jVwUm+6jNipU9en5qVyNJZBJViJug++nKua9AE+MGn9PFZVXD
AmNfOkDdz6ll8+dwy5IP7p0evYrZNji7sZ7YS7wm+e6QKGksOAGo/I9o0boYawyW
pyPdsIarE0xJy/CA5EAdIdnihOoBGlUf/YqaNQ6RDe159hLvou2qZfUJjjzV4322
Us/jljz7uNdx45oYtYJnKLEmI1QxI0SmImG4gxb9VBeJMPh7ZS9sJeA3aBv9Lj51
3HJ5dAGy2yOL2yPlcepet7G0ZZpnwLbEw3vhm7biU99Tc2VpNAYpiP7pTWTqt8VR
noU5GZaSpuz3dxSsZ46gSMawkSA0D9G8JYZuDLuHFKPKOD30n9T50NUwwVxp5FVi
pXqn9KJVOBACNbYe3P5YEW5MdvQ9K/T+Aa4HbC4WqB4153SvsncxJI/QDtAQuDM4
j72HrMkP6KnTshpphT9iqpi9hne3UU7632w0TM9fNaxf3CBGoxXs1eK28Zop7qNn
ckt9o2nXIMVy62qppo7uQgJVFCvyTlAm9Xrah0CczsHU6HYJQTLs8ny62Rb9ttkI
wYXSee3sbO4W51vxG6YOO2biCxbeTeNICfZxDVh7nXUvHUG6X23zeXOAz0eQaTqJ
R5iYLI5heaIrBIDyfsY1JtJigVm1X3HOuz2x5T6ZuKtmoLbw2lqzyEb7XOWW3K5H
hHHj0uAjvfRk/oE6dC3L/hkPs9P/mdPkuzkYiohQdDkT0AeNwf5csFBNRS7qrKYh
4CspHD269kezGstzAswTXIEIYo4q69JeZDHYbtldr97uLRzsSKKCWf/Tir0SrxAc
G/JbxyJTCNPUJjrJklgtaBBI6QYVBfv2aTL2Pjw7LHgIeH/P//wHiKu/n+Cuw6Zq
9VD6/DdegNZ1aXxkrvdLsHr8xsuQuPyw5TaADtXQDW2qwEmYhBmgH1klAI3pFmLf
WrDil5WgD2wxVTqedoyrFvj6sEUtJPUVI2g0PrKbK1BkAQFB9/knQz0q1hR3lMgw
mxfgZ0A2QnUwvPHjyqnWb2HO5JW4OdHY3if2X3GaVPapCAMqa8jNwXeTlQ2PUByi
IWpxiXruTmPwgVL9GpYaIxDbIRupmVSE67VzXewv3Zh24UUMONaT1Ns/wqzwx7Hl
G508C4q6X1459oMvyggEse3sdTPQkAYqBItWTknMVgY0NIxXpcXLAWdYNXlY7zwx
GRcQDqODWf+QVlQvdEN4cgICTxsossFRf8r5dlvoFaK0m8qXH3Yb3GYDAa57DVWR
TEUXgRQcpyTFyJz0aDwmBVGGMpQZMOYlMC+63rw9EucY67YliHcrnyrHe+a7uGeV
w79eGkEv/vBzqhjYr62Jg1TXAjLmHaGqxSVrOBlncjHkZ4Aa5m/+bjDJgCqMX+Vk
PiwTFqq7rFP6nzjGwofsOc/CsG06un0+PqvMcvnvD3u1+I8+SZsppOZZ0z9PC6sU
8aJku+OcIylIDwiSHXrx/LxYgtpE1vHAuPmwwcUWhzb2Ygjeg9apg515A5FLSQ62
A/dCDgN3zFwLUEcn5fgQQIG8GaPIHJ4udHg85A44fTl2dzNwh6hLYpZs8waVcCo2
Lef99j5mId8r215ZpFOTGelaqjK7pqjMC0jbJWWENFZNPDRi0m97FsZagiWVzuKk
vpCgg3ezuhbJC9a7r9l38hMCWXkZKxq4mDvqyADt7mOuSaJp8Ha1L93ynP7zSBRU
Jj2tF1Y/iTxm1O8N5AdA5NT4xgp7G4pEbMuZEKiAjhTvQ8Hjc8/eY9ZXfvoDY3JO
WYQE9gQOg1SnrS91ZCXxSdQONgxoBCffsz8rzhFe9x+42YVHhqLun2Pf//Cz1Qbs
wG9TD0r5Q2eqqAzC/rK30zHLYg8nnhPgPGIb9QwNwlOr75yPCFmohNp1jaktbHV+
mIIObi4DrybljCA7KhY5bwLAG8bAtQfh7v4CJY+9SXZ6yeQR8KVuoCxma7qYH9kz
IxIe3vgHbUIb3WUxlwfnx10E/CXZD2tSfzwJpz0SFLIpGXCCWgDd9+YaDgAwKeIK
tKHYFqZZlYs5BxfRfEV0OXj/1O6PTXqy44RP9mXQ+cBOTYMfKsjPzyVehCia7c4A
vpiqDomBRJm4IM3FHAG5doa1KszivwHhhvPjWQ6bHUV3ry5oNhR69zeSIHG7sFtK
0pduBU3zxFierVnv47N5dmNxkgpoUPWcg5OEjRIf1rHqqH36OhB3f1XcoqU+z/IJ
Tw/eMRjfb0y9/qos/yn0WwBkUwZ98NGg3A1Sps3zPQGvbR/7ME59Fhb33er9WT/U
QM4cQSDHjSjaIq6CwIK79BwZGwHehX4rFBombC5Rd2xabfwYg0qYE5Sy8WfI+dHS
jhf3n5xa2mBKo68HLzE+5rsuIirH2qVnuXuWnvNNhYoGtIgx8a8hr5OxkgG/gXtK
3NUzqZ0RT0/Iq5bLiS+oeKVIaneHNWYNZxPlYFudixlEDrN2k8/KauUOs4nEYDVE
nuZV6P0Vkawnd5BKXQmToH+7b9MEDIFeqde3ODwaj4pquDITa/lWIS1U+0fk3QbY
E2WtnCrla0I6QiJmdIqr2sFSgxKY6vhexuvELp2khoU4Gl70AzqAufCWY6C0NWgl
LoF3hpFxVGq3JVNRejRFs4w8bGYeVGxW3lFU/dUvPGtmap4cGrgQppnCJDW9ULv/
wxhHThia1ehh/LNB6PledHYd5C18TuLTjrE4iReBBbMEjSdtiH2bqOxQCxuUzPeh
z/PiZAmZgWdsdQymOAUSoZkT8Ep/D7AJMzCHDQ3pSQ4ziOtG5kIVeVfrCmS9XnTj
SSAi6iQTfhQ5BDgsC/sIsThUrc2YIrOVwjrcOGiAvX1Nnza2HJjNt58eQ/3OQZej
4XPIo+HM18JiL+COrmKW4F09JkOBNh9qilGDGDno0ssT+lWG1bYWJDHus5hq6ViA
ozOWrjL9AAReDLkzs2Lxac7/RxZqtMDqT46HFzvkZQSUCdd1MxOUza9qHmJ4uxUP
8HysbBkaDlmZZufrbKCsgGVrsxFO6jcP+bvl9YYmTIoEpdog6G1gsMUgDn0+9r4J
4SYpMeuJTQDHcJzXmmrjrGVFdYaRGnOy59i/xghve1iH8615+l+zkcyEpVRKSXFy
3hCxE8WhLbcHR6i25arS5OpxpAC5wPBSN4kyzjXXPkbFTMTFJrg/Os0GXpdKszjh
9z2RJNCSEvC+fgFZt0525sD9ivHDFTS1HzzamEcqA9ivgr0IuqC20hSn0CcwfciU
1MPoJ2M0KJaLN1uScS2YcqWJ7symv0I2I81lzALmVJrLaRRaR11Xy/0/R1FXLIXf
A28pdSpmdYTYZTcIs5PoeI7fsId5cj3fjyapuf2shdvF9fZuiwAhuIHUDxDkm9XC
gO/9GIjGCf+j1BxUxZS5C+nJO5OueIjuauB7HwfUzDMLLMGeR/Q4dJIFma/rhms7
hcXG78hi8tG9b82F2YuXkm47Q+6uOR02c6ETKfOAd1GS7i8xitsxoZKsUTOT8ygT
eKr+EXDuSxafvQ3ARxKoYgF+SoS5SrUX1I3tMl7u8D/5XnkShzMXOiB8sBbkyMj+
W7b0nG1OFlQUa1w4VtnJTYJRyV6XGfwY2PaJoGzd1FBrF3h5mziG/SyaQsaOd/8q
R/ZBfoouskxvNJo2LvDwm6CklLkWFPU39vGHMRTLSpP8cb791uzTIKF7ZXa/daNX
qFlVvwk1BfKZk0xWWfHPyFMeria8ODRlNvGfYeNx9JJcOrPgva3k7XIR4+xY092C
iZLux3d8zTqkKor4yOl1MOWEs8UAwV44z1ia/5O36lDsyJmstDVBxk2kj/MPI5oK
UOLF1UmULQ0LfnhfL/7TqtH6VJN4FkFPSc/XyP39vXnubA2DxrkwJ8Qh9rYvbT/L
I9BXw+HPl2R39OCK6ZxIJC/aPeRZsgLLKAu8K7sp0IrPeDbLRHP4O5mJdWXrXmMw
37lE3S6IyZHuaW5VlhOPQVCaf8oXCw/Vm2wVUOE/mnQC/CXVmeLW0yivFp9xESBT
pjlqqVgER1MCtTE6LbLojmrk5TqdDGllDi9ZgYBs2VI2wcsGU6eYWZnkN+NYcW2w
ca6Sak0bEAhJgbxsE43EVFtkbAtqF7k+fLjtTG+tIqiIFJOJGH71PUzNH0K3Le4t
Mzd9mGbEXkvc5NRd1rZteOKkTFWCD2QJg/KgCY8QOy3ag/eRrz6NgCCiNx4DttZk
anHbCOV39CM0XW1GjIsTxC7DaLHu98HMC28d4wFOrIG6nL+rYdtpuLKu2yMDrPAF
8ceOoBrzqIPt8sQX5eXzL7CFRKbo1LOVfjyZZWUa+pHAdEulxeWZPpeEdM4ApCkr
v+rch0vf3zqK6lL5VuBOqg+dBaJuxOOViQ46qo7aUgpgShCMuVOY96eM3+OPvr2t
azs8EE1YhzbZY1KjTV0RPnQezR6VxXXLnrJ+q3r0xiIPobC8Y4yko2mL+esDImBX
ejU769wNJ5quWLdEgia5hUlO4yAExwCBHdyzgf1royJJp/akGOL4+Nu44D4b7Tnr
KYa+fU0Nt8VaWGCZhQpuEJ3wreZQ6oH4+J7RC8nBzLX/iRgt60AVg5VO3mGbZ7GT
yrBxlyqvtsbVaUDB2yxSzqT5l6XDU/L21VHi/FsFXM3em6U4UmIvi5T1zUwbL0NV
ayCYe4PYk+1odw60wABDzOeOzZSmzSHcPf5ZyBAtnORXpVYIEObZ9+i7wgtLG2LD
VrGII7TEJWuz4qjYJCVDEh5qeuIoCyTfxkcCBBfWxwNHMavS+EhlatRWnHu+Xbvp
5ReJnQi4DNJVGvE6tV83Gsu8ZS34q/qAQntqUF3vKk1D+K7O05DQBJybsoaiekes
PWwRJhimCeQGXVogb6P0ObohtEmvW5SqiVqnFhvLExKMBtJcWZmZP4dUbVqqTx9F
FdibkmaoIlZdXmAtImlcHbl44MRjQxCzMpdGOn3zy1ZsaWMVDaoRa8vU1clim7TW
TeIGfa0/nLmx/1H6cDSfN2P/jjIYEen7uDRtEL0Qqjg7jDqMW9PbcR1dlabF04hD
vb2ZwvErQwHUm98L27RaJeZIbzKCSd2juPnCrDVUBVAYuF0nvqgkvo1R9u5ZTfSX
YxFPdKkIkjhzVsgmNc82L3ur8DiDNUyGNft/oWWewFRHC9XR7nP4JEGv+ci47nI4
u7jSMAeep46gL56y1TqYVlps1+r1mJrcIrc9DxMBu0dTGsELzqS0zQGhyOPjM30S
MQmDSfGaZG2GznOZ9wzcrKL/wOOipCcyLjV1tMQiF7hIvwJjPN0TW3ByPFpYEFCg
/m0hLR0sp30yxYTai+pOs/RTU95C1f5Nl1P4HTo5UbtJk2qFYfnXU1o52PYVXTL9
WejoIcSDFvosphTIl6WdHlmXP7VQh8WA+bnkoeKBR/NXmnh2a/6xBsjW3gTrzHHP
+BYGXzl1u3SZdaRIPWxdtYZVdKC2bKb/F8r2vD2d5yriUPPF/mPZ+kdZRv+vZMXA
HPLWR5zGDDI+U9L67Fq4H2KeocI0ijIkWniyufyIe5UIZEQbvLTqGR1BzWatHTBu
SAGJ83YHwc9iCOO9Tar10xMSFLDJJLHwVaAxCiBMREz9KENYfNtMeB8ShgThBxQi
EEWLUWbLJo6rbu4SIgWy5FtI/0KXmX8N66NHySMl+oifXRT7LGFYFIRN7dN0D9Fh
uCG7y7ihGwg+XjUUorL0DjcQeM6AxzRiV1T5HDo61rKrihtzJhLGIZS1sBnihRMf
BFKJj+06PaVX+F/hFNq8sVmFetBV6wdYZZuda8kjIWW+fNbCfyE3R/aQQ3jk/fqb
EUJBZ8sGbd6GwUBqot/Ffdd5a6Zwa/kk/PDTbpBnS7+Be7dkbr8YVvZBMMDJyD1s
BwpH9BalKWoIOk1AlORw91Z34igV7F8u4i945y23Gjlm+BsoYBdi9szG1cjDPrGa
EwjJLh/dDFjjSvJwPawF7bc76g1woeOo/5fw4pmwxWDaiD9ir4QAzERjCYginDAB
vkBz5VetrUuJ5Dyiw/fY8YpSAono8+0EwObV2iRV2Us5ocoSfbuz1RWlchFHsQMX
heHieqLuos3UknyQ5ZyRSrisrZxNn+fU3T1HMbuYGdyhyg2SsTxucHZPC9WOGAWu
oYk+7fSckeN99HaJZw6TTvk1gJHERe86fFduBoIE5eqxcw+9JbHmbzLTki+iaRD0
ZW6DWT3RtblWZTB/+9sJ0byjGSR5dNtDljn5QZAWbw7ILcKIY58BuMOMQpRACAl1
6D8SKVZfn5U85OtzXgxu3JhyPVJCEiFp/hknnz8m+NZoCi5rq/Q82hR5hUnY7T3t
1pAgCJlrvp7oZgh0OORiEe0QO5fc4smZUTmj0UeRHzUQ8SVMURnTzTVafHvLR6vM
3OxjsvTLIrzNKmAFieJPsK1FWhLMkn88QhUG6ZYieNo6WkGb3NHqUnY+WAk/yIOf
pPLUl4wCbJ5nTExhRxR57tfjRv3YrKGRlgnbqmaMW6jTrltax/rjOhMrdJqC3wBT
AQizFfaBcr+WBKp9d4bFZJgA8acydAI/wU17MYZi4842t+U6gVlVundBfcTfILuz
rQ8eP7q1slxS1w7bKduhcD5E2gBvIoP7Wy+ulnSfng7j74MnVpRXjZgSXekVxfUL
CiMZp0YhWETf1j+fLTmIbXKFMGObV+PZqTXyAlJ3ELiu0gphHNEzj6X1gcecsMY8
+3BcsRFT3bCOEpaLI/vUREqZMqREzP2AfeCdyUPOUoRKKPivFymTSaOJKJf3BOC2
CIIRce+YMVEubua6dTcOkC8/XgVVXdOITcwp9nBbOdjMpZdDMiH7n9tub7HHLX/A
8np6AVuHSrw0rliZaoDSl+HexZsAsapR7fEz2f6wyNLIl2zrapO75L2unIOSAcCr
5izlqekRNhtsx0UV6gRBHDeEaphwRgpY+Nyu32Z5ROGEbYoD17U5X6/FycOlS5QY
t/n5G1A7rlOAVJhJ8W6OslMeHk8Eh0zucAAoD3rpTp57W4k79m7YpAgHLi1xIZzz
VMAXEGHa5Zi2CyH2ehtV9P+vm9AOT2IgKWaef/nbBhqdiO37x1Ft34oYGoc+gp6j
gwlpeZtD/DeAQgUKwZrvbDyjvqd6jcMdQTyTm4SykUbol9xwE706rzKjlJMwyie3
eYXUpjQGnS44Gqr8yyIuabO+Y88oL2b6y+RRXPdNv/W6jdLwaiCd+4X7vvQ0E827
kiKhSqk+9dABNDh5Nz3Luq7M9jVIbdSDm1poGmK3uYzHDlIkSgdsQOZB4mug6z3R
vKkXrj71K8yJIISLrm0lSmbIIKeGISWs+SHFoJudI5b2m//xnGklwGe3DqNYc/PI
v3rDaJ/BNY+k/QZ+K5T4GC0DHYffMwImW6zEd5JicqiuqBn6Io2036YfIes9172a
gW8k9MgpIoDrVrzdm2BcoMJ1zPwxO5T5aDUHS3ldiOOU9h0BVFbwE0VpzZwOpfGc
c6HO9GwkO3QSjVmyDi+SKBc0BgnKkvmzB9/usQj2PNY4Vo2q+p9meMo9ReeANynm
C6fcSMPdmdJQztOdtLT5xolJ+dWW/YOdsNz64q6+rrkemzSJWfZnGpbiMnpejA3k
gWwCy+mkBW6mVSwWt6a+0OJqN756MUjHeLF4sxrYp1baEvFnbPVMUOlLNh/lwj72
ew60KYizbk9lBF7jtcyb6psPLWDaBuWpm3D2m6t3JcvuQjvTqxT5Fo9BijiV2GLf
kDnlnIEj4J77C9nYYLaYrKrM29AG4l3Zd3x9wgoKDSbtStBEv2Y7zj7QTt/CgFlB
mkXSHY9bOjQK1krFUcmvtHOoTy/+Cw9GNShsOMwjsxRSD9s7Nldkd/XTnFLh8mm0
PNea8uUUhtqe7kqusCueruaZgNc5ayA2AFiUrq4xE0AKkXRHgEkaXhgPkTErQGco
udt5gqxiexMUgZTVVYcCZ8boHOJoyNi2C3QWNuIMZCs+O+V9eNjNx+oo5FPLgpxd
M6KODw0dcoE4X+OR701jeFLhzV+un7BJV9SZhg4Bd252WUAVseKo3ZYJL2G4smlt
f5pkMBdItXFt6IjxLvc+kepDdmVwwd/3RcSIcbDhx6w5U23iNmfw4d3lz075yrRN
I8mF43QjSSf8UoIJlir8ApQBAb4TNKznhVKxL4rys+6v6BvfY6AVdSdQ4Mh2nmzJ
cdP+0KcS/crO5Bssc5MDI7w0s6vaTNPLkBt97JBMHYJ4PtBLyPD+tIRBdM42OvmM
h2yVviy5EOX4q46YBReK5nWvsgoP/Xso53xgTf1JCxov+KZ/wzBmMEIs0aCzHq8e
/k+ASkWNN4Gtw9f1pX5VYgEENR2JxEQ5Q07QrIvKHeOVvC4gyle1Dvr91F6UTJu1
aCqPALq1Sq00qGJx2nz0cU3oWdcI6hmoDVWYEIMYm/1e0Ekd9bns0ussv4EXPRq5
mBhChnRkxerhDs5p/Uy5WtHK1odlireiGswoXXo4hKiluIxP6CAo0j96Kut61htQ
855kJm4QPC5Ju4zsQc2JoQ/ZKhCmXux0jpktvNvZhASFf57XrXHsJXibFRQbqatr
do4mlOTMzCtCopz9vs3Hf7Ua2WJXoLmDfJS7RG0UJ4NTcrfQxx1yTOot8ekb6Vxn
eacJ14qQaSi/8AclvsjNDoIMneUmaKu5xq6xg5rnWLobEuIwwfK4VNPUkW+dgBbx
Um1I45pS1zX99SdZJshu8hIe5Ft6Pk/AX9fAtk7zrtmjCQZjQX3p/FmETg/fRcjr
7ym1ued6v3S7UYgFM3Xozp1gzVBpAh0u03WkF6qoZkxsAkBXXpwJ8p6DyuM7oUuW
Fgr+YhIYuzwRB7pJkCbZ3+LVZMGc59Izsec1nWCfsnUGLhza/vT52+5WdRVSAppc
3s1CSTCIII6k3zz7YAtRYunCx9uFc2+pSd6DTC9ezDmjTsZviQF4xgqZnHKDaijk
por0dMVApGyb2I/UFQb7RvaIZX7524Cbl9k64ZiPmT28GlZ545d82JI7A8Hwe/3D
Kj7fBkc5zR0s95CffKgCXSwW1YD8PZgvSTwdXxMvWyM0+MsqVX6TSDma5f2NPkK8
8wD4Lfdjyb+Hufd8mS97RueTPEk6km+zIsfbqJEhX0I+6aq5Mt4cUPlAZ6TXicic
Q4QxGQ2kc9qAWHQTmzGCX/s5CdGGwED95WjGKE8BpqZNUVBowyjmF2KdzjHX09Ee
Xzwn6t85tl3/4MtRfuUiaMfBbrGwwXu2hl3o+qTQlw27OYId9ixBlsyMT1VE62t5
Im6fgZzu30LIyCeBGI4KLuu277A0ovTOcPIHsWQZRP7wGNCX6Lz4NeXkbq+KfyY1
tYmDEvWTTpa8ME5lmk1GgBG5iKA0a9ZieuEYlMFP+x9Ts52Ql2TOYrYH+3tsfcXA
76AAuW41BGCSVjOAb8RQwIj6X/jqtjkGY9Hb8UH3fKS6KHno+wWkDcZ/78pF3bZs
JYT07NEEkHq+8a8ApvFrGhVo/1UvT8glzLEymFU49I67U8c+IxJMtSLccP4IyrOI
++PZbtVE4E7mfjVH9Cx7OJ4ldeqsDwAv3ti/ADZ0kWGJCOSJKhd/pTA5M0RgBewX
qEVqNVFBE2SRq27TKEsGVXjI8PQ9sNlY4a88/K8+jY7DqDe60YVQuEO0IIDFNsT/
sC9eb8S1xRuirxj/482NVh5sT3nRrdUPXMCWPgBq8sBikJhAZi9zxP0mX0YwfE4C
09R02PgAm509fKOB7YPDDXPUN+EgR860oAt12zb2A0y9ZS0PNpTnmVdZKZSRpqMC
r6Pq1ObyjNRSf/dlEC4jN636jM5pRwbRAtrZQVkZt+ona1ddTOrcgTkA8epUw3CM
ysx0Yryk9UVet2xcy8Fta68A+XOmhPsAo9qtQRpTDVt2kJ1FforZxG+bRptjbojX
0s9nm4mbrSJH+gNKrEFxeWj7oR5hhFHo+FNXBP1PE5qNQRHWrfEcgaJ70Xz2zznE
gcy4bUb5QLcu8/fgeL7Q1XngnUWKOVarObh4U9yLxCnaBO/vXQwdGxIafHZfaCUF
BNoqKKldvJOlSasDnMWAQEKUaFjvbWF4I7+ZjFtKz1IiaY87mlvMyIsRUlaJLDg0
sziMsckLydMovQ37Wf9R6zxuWT8P++tBwjILgiXHLYwewAuf7wpgyBiRE/Mr+Phx
cWn6LFF52DQNacHU+VKUy8PgdPcRMsKswGERwk0NVOQRsbYwFJS/rqBY2azKZ+KN
bkd83XoCZhL2Qvb13oeauq4tHRaGwdLarhligM90HYFSra8muAg/x9L9pYiv9/9y
NaJxeCfQK3JH+nH1XX3gS7l/IY3W8lr4QaoYNZ5O/16cyp2WahTucCHsbIHTs0FZ
FTVUBnUrUXddVNM6CgIipHNbYYWrA+THN2yXuvo2JWEeJs9Mnxux0+H7tYrZx2k6
sSsgMqW4WL4lzae2AwnHdTrxooNuUX9XcWgnkHt0LSVhyPZQrlA4hw92+Rwce3hA
I+ivFes7O+chJQ5z/uQoFSZNjX4gq04BlVHDiaTlcBquOX3tEt7KIZJztsfy1pry
+TfwvUA88Z8PBfY/MGC96ldZJsT1xVC73c3OHPlMJsM9g0klJ8u2vQBeloQh0aaU
UhJdTx8X6hwj+w6ezSF3i5VpmVcWMw5Jegic0Of3RgD6UFwHCKF08C4kxzZo34C/
b8/qc//hwM/uW/sdbQHAlgz+uPf5eQR6uLO8F2ZawJVYyLfIA7sEb6okOvuPbnXG
jsG9cQr8QW2OyTTk69VbhDbdFtQYX/P4gUqhnad/vvzk1BjklyPuus5fCENg0Y2p
5+qfDOgHkMGGWJWu3erkVwgeYJgfKSeCId3jxmBt+v7YYFSc4jIsvRGbLV3486/I
Ou3skNJYJ1i26oRTVDkc9V5i5ej1Mc1dEVwwdYz0rt98/RsCoeACysWV5HmOwFvO
LjDbKGTbaccmYcsQCBtRu0Z/GUSwtq4z2MQR2ZW+IIcCSUNiFrzbrZp1rDCEgNmg
8MxL6YcqoDIKFg5mG+e2JTiBIA+roAvkycd/vs5m3PDfLNZMgLy1FyQ/pbSmpAX+
RWrqc/J3at/eZizwnDFoBfQGInBVadEviYxGgPj1R1pzU3BTjWkd3Cgr9QA6Wk0P
vWmMwMdCUjE1FFLtwDoV/2vbtW774fmURRWo1voSLWQIxYgjc1FDCPY6WZv698fA
YuF4awP6Bbgv+fiYUxI43AGGehPELgHkmVJFOKhBekX/L2OLM1rImGTj/Br6xlOU
/c1h/cI69Zq5W9T6+miYyW2r2TtE1bj31mk50ucx0q3ZHHZgODccpXmUpCSsw42H
bwznzH28QDx95na5NCSqkjFYC6vQr3jZBBodylAlwQmY4vT76aVwWGYHb+9gbS6g
gNuF4abc/Fn23DSOrrGJximtfK+XLWTK7ylDFz1C6hXFuf3MSb2ergShC1GwWSLa
54oe2qhsy1Csz8D8Vgyjdmx0CniXsLJiPz1LCZIxArJusV3YfXw+Oi4Z1ARV2CMK
WmR9VnjCQ4/GnDTmmgDiSeqNUf/Nt5TSCFF2q2hxTwKl3HGqMS/ikuY8PUTOYarZ
EG0u/gq2nv94mT1u0K2xSfWGHgm5uOoney8p7rx2+X+slXZAkDUZEdmNA0oivlMD
m8xGGkFljiBL/tMjqPxOJQ7eVg4WUvke6ZYjg8jdc4H5j9utWW4mCKM5e2bTUi7j
0mcGn35Kf/WmrxGAqNunlovbLuNEfVaBG1kvtclS+c5BHtF1ECJwi2+nFW/MueD6
ti9u86oddBHs6gWmKN2Maa+tKOr7WOIfoT/YMg/X2teZqRrB+yqp4RCCYuGFLOQ1
zyDBrndk5j8PWUWEGiNRoePl0qDaI9fVExIRuKLHsMQlCke7T6I/RdPKNImTHXYz
8iQq/c+GJRdGLxB902XuES22SXM2nQHMKgIZGAvKYI4bP6iKSAvuS8al54YhUbhX
JazrqAqgX3fTEVaMl6m0uZsficjMsE50YJDGyZZWtYYWQUHncTKLd3mkIEq76cqC
c0s4dTjatMLz/vTTgKWQjY95qzPb1CpFIQON6R395j8cMwtLYTPGOAQEriubYWTh
ygpm2eZJq9vvkJlMDZVRPElQJ1mTrRBADlgyGZfCgC1sdUCYSLMKdxCpZ/XXJCqk
DXKoNy0zglfkHWhqToTZFoKxOHqwgyTaEfZLTos2SXIQpDmhbi0ee26dHXxtFTlM
2WwP4iU8LAism8PdnklwCeKq9V422xsiiZ5CwJqpUyUrR0vG9+2pobp4D6hCkSsX
A6CDa3oRCJEZl+H5EvOcXxfo+EicqpPTVlFfqOKgW8jTKLxF/rbv+y00PLuADVjP
baO7RUjbQf/IGMQKAvYX5nQyOiIpVqgAXR44XaXZ+cqEfplJrWmY3uT4bCu0HPYm
MMUyP0LKtjNyUTr2gE+KaP61Y7Nwa3FzY9q1pTBY3BJC/E8QwW3DLWYPuKVeYuT5
1VnZ1Lh70FbsS0mLOQSmIH98iaUYuyRxpnb7zJSROwXM40xXt6VXUO8hS8pnjfYA
dUEpe4Pko26Sa9luVcsgDQqdS7K8ge7mQSfGsWyCn9Zy/TWi1UVYYZiRxF4nm6vk
VhXPurzHAZeXB8t1da9Iy+Q9Xxq/W2bswx1qJ5lmmj7YXPM/onTabYwnxXGC44zp
`protect END_PROTECTED
