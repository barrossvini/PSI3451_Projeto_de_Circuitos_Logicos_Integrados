`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ghy2NEmnUt1bo7GBn72aD0koDbHPI70YPzE57gvgiyiIqLAcNV4o8PNRau0X8r0x
r35xx3TpXAWwR/LMiyQ/ZgtEupT/LLXrAevpbRRX5DXGlbdrEn14/NZzSjRWc7JA
xTKJ5/KqSEN+WQ81nWUwLnVu1ezYYPckFZLlH3peEGFnmXaRZucZFfDdKUnWbw+U
kh181d/mbUbkn5HZBrdXI7uaOi3Gc/cnMzs4AsFElXeSJskoY2GPKkGMqZipe+VH
uggqhTD60+RDU5+7eNDZ+nSbAO4Azz35K4wmadMeB0MofKCvCT8az6peh9kvtdOf
9sjsrzOXE0CsFMQwGKTrDtzjzhNyTGuiNHZRERRwG790R1/k+TVjQiVJPR953znS
dRTAp79oz9ueQQEjFylktqBOIZ7JzAUWsY54Aeg3BHSXGd9TBz1SIxrgdwMBscJX
qDBh1elfZ9X5nwDShwhLlQ==
`protect END_PROTECTED
