`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KzU5KSow5xtNurr0Y2AYpi8sUEKBnyZkSjHnbN2eFoS7aSgVUDvczm8YhrZ1Nw1Y
B9eDb8mTRebADV+jcWYyPOEbO3CVz39TuIedeLWEP2lQZxWBHuB7BhlivHZkBwEx
7sJ6ulgbTblPZBY2/8plhssR+TYR7sX4Sc3I3lmd8ghMAgfE7dtqap8HR9fRJAZX
bD3RD0wmu9Y9+oLWUZhOrZRLVc/lL92Egcg7FrumGeGm10hE1rSTUpYRgpLuNj+n
iRDcUpD1PfX9F7GPfSvjdSeeY8OjihWKymF7t66bkiYAolyY2P8QIeI/JHDZmJ2t
zMYaM1dv3Jeg+QkSoPx+9/CkpgxY56foCJp6XLv7MjW9LQ2Wk4DzhWnUMOt+zvvg
dyF5Emw3pLY1UedeposKUg==
`protect END_PROTECTED
