`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jexA/G31/XEQBx5RmkI5yCd/IWS1RTUZL3dwpRQW+9WAS2Fwi+4CWdIEj2zfJ1BI
H9UEL4yY4qHkLbyq37j78Rs88tf+AVKSY8PHcH9WCP3vGn0DPE/qCvfMCE+flsjn
MJh8JrjF/1qokF2/xTjigXaMLJ4hh+ZiswUOX41VyQX7LN6JOotjlfWRbjcn/QCk
QEJly8fA2GT/v2f3ibKGfQkDoMSYjUXOT/uH8HCmtOJsuMLjtvOeN6gOYzXe+z+A
+3M36EF5wRzj0nhkntq/fU8CthBU7t5axg26zN3CwfSfub+RcIPT3Y0LdUNSAxI3
vkNGAn2wp/qEcWZFJYUlZgB/okRC2DcwnTTcGyDXyrD0daZKtrb9Mqot2ORgSrwV
gqeZdjIcimChxZP+dm9AiDzvo7+DWF4Mg19NhoFbtMUhJ+0Y5FgOz4x9O5zQpjX5
JLiAecb2A2uKVQC4vbCIgCAbpbZb0guzdH8JxtC8hFhjFCwMqbCEf3Pz0U9s4EHc
PqAjEM2d+ALpS6x9ACR+r/Svge7g2pFRVQVJRt5fA97xKFwZgvPUvxCPLbyhG54U
VyewPAdU4IzWVdadk6vy+HPFQrYNLDQitKno2gkyIcf8KYeQCzCiTISg41gXka8A
WoYGaJS+S/L9DZb5MfYdmhNcy4khQtCGeDpy05LCCWTjEh+XjR8ZZ3fy3shZhYHx
LgUxzS/7GS/ej0Zdn0H3gtZz1DejLncnMHM2MwZS8irex3ejkH0xB5B4H+pteGZn
/LdDSqIXC+BfVez21bSn9V/y+G6zDT7RZGSdAZ3a+VyVpWV/JK9W6zNtN02KhZpl
NeS/k0kqRoPHtpOGkkfLwMvSleHe0YISipv56neoGQT+fmuzK0QENE4GqPjPG+lM
IJHdeyuow8LVfBtv9cF3w462KbA1rIpMbCUHnQqCvwnmCv9YIz6M2VOXKOpWYUrp
PQgYjDoh+MMtE8V4bZJ3knURW4pbvR2kLRNttW/zzfuApZ3yelE+cEQGEbTYTbjp
4SqP99w7v/PRzw/FHh8Cy6yGaSSo5ixcXlNflmN9lNEZBJkKsxHvSN7ksVGxGFR5
kcm+4J7BLeMU+qhsez/zeA9GOhOiT2lexzP8Y1KWHY3TIHiAvpAVFFVFR3a/th2J
HzGK3J58SPi3ygozNyz+LYMXMfwrryQDEbANsS8Ti62O5TvFFRUyEZEDNP+rJYKm
XPWOQQcxRIxRD7j9//d5EEyNVpMm5xHSuaTkvzH9tdygSW7U2/gxINgDC7CoJ0TF
R0LSxD7H22hEuRvn8seZFYyRBNYDqEZ6BT5C+6Kf7nRXWLNPnTbXVhh/mHnzlT+9
2QK7sXaGG0KlTQJhBsZ43343ulVD4DCmRvXcbhvlcPgLJZesQGkW5CiRJI4dwFkR
X9hZorNBWzC+2ZEsmBw0qmCntpJAJ2IBYJ8qIxxAaMLdAy8BUXgWCPjYlOW5Lg5T
yeHbcKrb+f/Sq0QqHoOJ2zobH7n6O16MtGtiq+G1AtxnGF2hkJMaXyA75m/N5qRZ
u7pzJlsbea4N6jJper0jgzsX3z29SW4ryOQOyFh0tlouOT6w5AemXACGW+rv0+3r
NQ8t1cefgOVqMrkmm6ruEgmTx97+fRO2+O9yEmTex47Z9z2YPEXkvC3TRpW9l4ja
C7+zLLRYoK7mDlnDVOVJa5OivoAjn3ICF1FOrAgZ2t8EyXCL/+pMmL3tMMl1ApU2
m61Xn9i1+MrL8H+GwGM3HyIdtW9xT0R5XaHS+93DXx9rzWan+ktzOhnt5fSIlyV+
J1Y2X7V17kaosJtBVKGpOjRng1KIyJ71ZdrSPKQeCTWRzuZK09c9G1xyi2U2IfXA
muKLd1HB/JOBIhj+TCqppBQo2cyjBOoln3uoN4knIsYZ35IOcDP01SEaOBd0xe+B
As5fK4bcqqEvkm+HUEZrY+pC+qqYWSXq8680TYEEyLlLuGhdiRQhgQ6zzh6g5bbb
mNy2kFspkQJvIH2t+dJ7jMijCDConbysHLYMuMFY7gJvAYSgIogLd0OH/1vINwze
+JYOBqabcgv99Ryh8inZD2CCXkccIQ53kfbnDPdq77LGITPCSqZPWi796mx7qaNJ
Cknve8IFinueydLbtFw3np7i8RfYTaoPayM+j6gKOfIqYajyUENn7eySxTYPOUhV
C4YzFIw7B0HipkdYe6EWPaapOqN+gig/XxsLmqF9FVhuo/ii2IhUkgzRGGYVl5CQ
XKQfd/TpQ4hHj8Z2yjy67A==
`protect END_PROTECTED
