`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gTnjt5u+zmXwXIkr0mj80QcVkEyouUJBtfY22yznLkRLoEuwqwOX17w0NxTBOX1P
wUhS8zVIVclXmPr1kqYVmEB6jUPO3xWpGPnPnr0+Fgqij49AOxirBdX6KEEztdHa
60Ge54HtNwbXv5DQuX8+9iM1xLxLSqCVjG1M8EP4w1q5sjeHw+ohFh0RHIk1nhwi
XuN76s4pmiqQi5mAb+XYRnGvcyJSt4liAsdgxa2BYj2ZTyBnbuuV3ZsnPfZAMt5R
zLiwfcmNz6eWJEQmlgH1P1SkTmb6T1yvIldoGxQy43W4u88e2l3p8o6m+hqMURrz
RqGB+D0DzNaMEaIhlNLI0VVylyeXxBFxR/jSr/N6k6aO45JUTGGpryj+1GTND1fr
oEY9rc4s7OJUSC6kJm6Gh2HTaR3sgHPH24zTShTlS4I/CNEajT9Qr0NF4uqcUAQ2
VCeGOBdMIR2OPOjh8w97VYbe6UyJrdWJgw5C8O6xTGVbLnHBdllfHCEMWEfkhJ67
DKBwRYkgm+5dmYvQfh3GptXFZByIF8cJOmwFBIxOGZdl3TsLNJYaGhBTTipoRDIf
6Jk51xhBgpH3SSS9MI5GHntoByvx7sk+8BU1l8Tj2FaCb1W462X/TZm6idnZOTEG
f2KZ/pMezwbCSG3ba0CMLe25P7vqncOcX6WcD6ePtd7X9Eln6Y5Ys8kmDI9B78st
KxR+IrOGYY81dMe//e6ALY+aaUBIwR+hmht4GOV1D27GK3jUNSVkwFla+K9d0z/g
HMapNTOfDzzGvpW+fYjh4KQnVWzhxMirkS6rvN/XA6NtoTzNDX/UrsLdkSVC1ExS
p8aGceMzmJ1E1NIdMCbxZnNaMdSjJIv3OCMgqw108s5cTNlctTFAGOodDeLg70Ob
lZmlY0+F5+J4VIBuc3dGfEdcb2Mzb3u0iIQ/ZqB2SM8sdyOMV9Fy+C0x5oChBb5Q
BGcTqB11KEGWsG/urrzu+zTHnoO/wTS8iSaf2VAAOsxzC16Eoyb37O1MBN9QcC7r
`protect END_PROTECTED
