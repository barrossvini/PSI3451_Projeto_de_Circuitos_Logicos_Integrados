`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
88g2YdhgQYLto0Y+DUjV1LP+W8/HG4ErNa2TdlQs/n6MDrzpU6fW4t0EDcWbKxuH
QQXNvHTmENyR7x+KuBiVD953Hb1lPxfJF6K4qdpQCyg2v0HEpBQX+FpR9TLncHXE
Cw7AV7QYYe0DZw1Nv9qwnLj4bar1c+9bI0nPTxJ0DaZbIQgACzIKR8dLBf8woMTl
sLy8b4oxs/wg83izv6qECuscXFMs13gav2sLxqUUMXjwAV3LHwq1Gfe26eBQc0Am
hQFvd0p8t5IRn0E80CH1Ctyawhq+IV09S7/1lH7eg8UfLuP/WY/HQR8QEVxJYM6W
gAnJeOlp/+9h3GIsMgjjWIoIxAaVtK8LvWj+hCE4V98zj0BBeKfzpOkB5OLhe4VJ
kba7tV3URsujTOE2LA4b+fVdAeHkmSDEx/K/MzuW+ihAoIgTjKT6CZcTXS8Rr7da
sNWkStgFJlsLnilhJlHHZ89BKz+9/RRJqmTwhzG19LE0nwr6afdNAPDa3SI9f0lh
F0G4TzSLJVPJUQ8y9xx8htJcRXc+81ESzUo9kbwhYRdQI6ceRt/4r8sEtXQVGz00
9DkLRtiu3Z+X9oMuqdOhsB3a/tia3nc4G60nlNv97s4tPBRJpc7pl0mRabA+0VYe
SvTC4ZLGRvItYM0mE5h67K361ZcOhOF/xUlHMZslWzyhwnCYo7km/NQzuC4ZdTsH
`protect END_PROTECTED
