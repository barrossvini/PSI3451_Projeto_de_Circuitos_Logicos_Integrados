`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gTWuKNkNnnI67JdDt1gmIHKwl4wewfAZAyfd6BrNuwXZ8k+SYqU/dFd5trL3JuLY
R3cvTqug6SGA0uLWmwRRSuKvCWqcFXHOyhB4Q8elmqgk+ucLhBnG+YzfGHil1dbs
DOgouvg59/ZLT17Kn67y3uRvR12XCwFVDdWYrgbgolwOwKUvIl/aSCgkyiILX+Xb
I+9T5/8U4/EY4h5R1KOcgthISt4RtZUGj5maDNHY91aMGdUPdXP3lq3O0thtp34H
2lOpuMtCI2EAD9AjSp2GCYQdLXF99igcnSSF28PuHknmJZRO4hKI/u521I2NNIJZ
C0dzy05ORZCSyaVpQ4lYfAKOtyBfEog62OyRWoB4wgPIvGKPzWoWknsjCIbab0Nv
+1qJA3EW4v0VMMwihuM22WL78O7ssRSYke8JQU4DreI6BLQJ5JnCSwnIoJoIn669
88KL3ZHG+6xdvY07hrwFD+qoFQchVj0+Jq9NxV/p19OmF+/Gs25nNmITY0XGnJdC
I9C70EeKFp18bcKXkc8Iqf/HT4YXlI8bHz5TitBsfPKHW+0/N1xzMn/opyo9nXXh
43KheiaxSc9LoWNdZJcHu58vbKBMvS0aTe/nKHiOpBjIly3QHvzBG/pMA5yY7or9
jbeZhgRS/nXBaoYav6v0FKPs7Odtotqsgipy0vTrFJFSeUdO4sESNJZdwYVcULxC
abdQ3uW2JLe+wvn86+6eCbQI55l6glxPfdTQkqfIuaog0vXU/pUhcIT2Ilf4F2X0
GT0Y4hU2l4u0/evBB6HobE92RWDr61UFVnU8ASFKisvMPipBH/o0FfYQdcZlrBMu
z0Ghpq0oTig9RAtoU2qjF+//qfoNd+PyEo5e/QWWQZgOxMd5+14GNY063TcVvgLc
GBJMBw8QPt7RaKhkbtu5D5cbdDhOOrYQ70Mi2FlJnsdSuK8zrHBXW6VgN/EjELuv
iRu/tKk2B+JXh8QuNl26UktE037BdRMaN38UG3PRsvzGPN4xEUag/JaFPNP/Wxkk
bV04nJSVRi8t9gh6ffSYalfoaTtodv+p+T48isDg1XmVVeuMiP1E+fLaIxfdrSZq
rZlxxcT2ziOqQk0JHdizbc08XgFkK0pM7eaJRlIDSbeUaVe2ak9+q4gN4tLcnPte
WHnWi4esHmnJMcxSKvW0thyvPLGuMNQMDEvqvmyyF1zfdgBJ6jtYmMAI1/GrhP+E
nOGLBHphLHEt27i4QrwqkTLBFPrFFTvuUucfOtwqrfxo17MphdYNRx418dRZg9wK
US+cJgBFKPxKcnieoAz7nbNCKBwV0nhnsEHdu/99v3cqjAlLEks+XMtHq+YjHPrU
CCcF26qmfa0DqHw7GajDc/LF0mHGiEdFV0YNdzD0UN7Q8n/Gc8kFud7FkgztNcZk
yWJVWoFYl0LHMiYpiUZzcVYnW31S5CFgLeNUZOg+yxjkvLZ+NpqzwuVb3voC6sIp
86vov5jOHY71pJMIAK1KtNyJEK9CQ4KeqQfCBK+ZetVgYFWHqYnyQPiBs5b8A12x
iNzG5u3TcchSMlwxm6mgqRpaarLcFrsnlYMZVyYfrCCCwt3vny3hsc0LsbDLXqsx
BGRMfHZbmJPyhee9VUsmxwYr3dOXFGspOLYSXLSnudWPzD/GwTqIp+blzTAlUmS7
ejCycXLf9BJXvPn34OqNFzHcmuEFO+WGVLWG+pT/xM1l32KasVssvXpJTg/5rMLi
mQ5cXdhRIKD3gXEMISt7VQi/HiPvMdptKYEtDLYg72476Ph2X6yEt2UiNPBr2JGy
S4E4dbHj4jFpv4jD8AQydXL8dkFlqG6/Yk+4lLnaoSynQeaX7qmWkxxNV+AUpVua
9Jl3DwBd0To1ReD0YrXKrYIfbzdvjAUY4ZaXvwcFsVqU3CADeVln7H+pNuZ8rl/M
dymQMbNvFjQ3nuv31bbn+QiwpvxBgKB1J7/elZfn8jaXwBicIX0D7BE0rpxp/+H2
YpFqQX3qpBzagCIQlX4BXwGU2lJ5JjGlWAS0TaExrv3FOEyUFrFlibmFv1N7hTfF
hH+X1RYhL276emKDL8IWQZ6anuLIQ1s5EUhcWzluZx+jv6r+PdNDQbKGjGr9ljrW
1aZmmXGMSBy0gSMswrj0QL+MqUvfddTuJ4IsPyTUTwXQsuscSEmtoizXXSVZnbD3
6SpH176h7VVcmjGao6bsZi6GJr4PieUa2HhSQ59J4XpRA9DiSezjw+6NGvuu0IWU
ajskExNyEfINR9qE8vg0jauFXug9fXj8ZGs3baexNv8pAg4de+N2YWQnkKe/+wnE
gFZYVu13bawfm0XlaubvBu8+esvxXGFxHjvrpH9X2BpAYqhdXZuqCg2EBZEHLW/a
8upaY69wLcO/gYp76d5tQZ/Ch0jkf+pPpnCtrdzn4x4javxaCMiKBTt8tsE8E4tZ
zS+etfHCcjI3V3VTltomuksYBnkgvj04HnVzEVoT7THhEzOFlF1Blcfrc5pEgT9E
7BPfEp4tw5lPapbJwHuJw9AHO3u+8syKOuASBT4/63kXKOsinmpdatXg/VbH4Izj
CbmwvTSEE+Al5WCWaO+FRuB10bJub+cOqk3sKG2v8y+/iIMz7rNXxErenATPdMm6
dT3laDnOrefLBflmTCKU0AkoNA+QpAEj8ogzzdy5kNSx25DAgJIY5YZvZJnqVEcz
exDCGkmCij6Qrj3OFm8jocqRFMK0JtMTqBmo1Eqr/bLpo2GP/fMBIlaZ1OLc3etZ
QHeFtWp+RvED48t5FI3yADFh7nXkjOIbsgQwJPs3o5ho6+unwaHfwQoUu+fOY59z
toksu4fPKGZSQ6+QPBA1BwphhcZZvMya0i+QujvgO3bvHwYV3P7cuahmd8vxoNpo
yTWfDu0bP1jCvexfOd7kkTR3E6NTH8N5rd4JCNM50TKJMQXVOrAqWjnZJY27wSY/
XNN9lmAxgQ52wSOQdDJ27lTvGqNlMvPFyGHaDSZnQl1dA9iOrTfl4s/pZBEgsf8W
kKwuPdcrApSFMVnIH/oZr61G9y7jL2jCyF86waA1lPZ2X3XljkVBGf74yMCVWr5z
+4ctV0yrM67GP7uzbAy7RTZ1k39p+kR7lZXzrySuOs4veE9U6CBoWiqR0SxdF4Hd
ridzaSJE5dUrnNjI2Q8bzfJO+ucrQseiBZ6WdokdebUDNjqI44hoGHyPYzlXPSqY
kJyfHeShmfpNrAR7W90IWJNac7sxtM2QLo2mnRmOTKxv+D6RYv3qaGF1Ux4fGQ5F
dOzJ6H3CSp8JRP2DWL+4V82C+K63QT6Mjm+FA0E+weD+y3RrwYg4fBSOGV+hj1tW
dPxpPnm5CqHyBJRbZsJMbYWjDU/zSF6aJ65/kvmgK0R9DP/Oqw92y0g6q5JerGLP
5Pw3gw19rvLFPKDgvNGTEIe1KLiJcSVZsgLNXATXhs3f8Zzstv2Mc80mRvxEvuoO
ohephHJcJRE8Ldf5bhlPHCwhGAu0Ju2A+iOffwfN4LLsPWszCtTwCWnsQs0YFBpN
4d0gohdIC7JxxBVeQjDdH4KQGfcIBT66bMy/WxO9rRw7e2qMqeZRtKVspReXrfSL
k9sDqcXV/6KlRQ4hYaNNCC8PH/bzAsPE1fmsUQRMXeWSUjtHtkgusP3dGObjodCx
RHUA4dkAoCga8T5wlVIkk6gQyhfZIE4LfpCJy7ghuUrd0RYNo3o3ENKfUyHxv10d
R99QOYidWSZKJOwun1C8XB7NcKS86/O/eCqy4R6DVxJO/g4foVZeaHKa8BRQtg1v
DR0g1ZIYZbiXCrImStjCxMiioNFM9E7xO5Ty74alf48Btxj5wS9tJo3hqOZ3+guL
DAKyiQ0RCeKltMoGTD4Mu6FuYMPscMWP2UZG/tPl1ltp5ATFTWKXERS/XRM68ll1
P6Th1GYOhlxgOkbJI3k9BzlkfH/or0xr+W9GMceS7YLNV06gcqnfWgOpRThTDHQV
GL+x9oVGxSVMSjOw6nSr9ENGqWENxmRJy8BV1vIFcxQOaCdqJLn/EKU/iflurIgz
YY+SVT2jH92ouV/UHC6ezosEYTdNV6p2ONk8qfaQ4/UhV0AlvFirpnCNaDocQZgB
4eMhhrQ/CpEROnm/Ss9eAKBsekXhpZpC71AUbpgtNLrnX2I8IUWS3dV1pCCR374h
hJior7OMTlvssB4GPPrXGeEQKNn48J3GK1kwVk3JJy4uOlkzLRjGYbe5o8i4vt1n
Q3CRhYz0istEfEIqDb9PI5pl5fDMRMWrGrSIdHT4BmVQ+QZRru1ojGutUI2MNoo6
OzaTfYHCuqWThG0jIWH9z1htKUTNAuEX4Tc5/Eoqldl/+rUNPjhj2xL1dZRShBTI
f7ss8djJhRWMtGBCYY9/V1cehfcY532sHtajA7+L86elxOx/F7C6Izhat6CYKGrz
ouioLhgOaai023rIme9zXhIXh8DB44X8u5fSkcV0qmb4/Re9LYDi84LzWc5CqQ63
+LJEVmZxIWjjRfBQwsSRCTHhN2JYPAyrXN2FEKgFYiPttiaI4iUCGLssQa4LYU61
wSI94Gqteo3Gy9RwxgVJwq8MRXTRLSCbOBzuQS26V7lBa8bnUVVPv6zLAnC6RzRs
TXVn5GR6lnGELXlqxo8ieqZBLrsd1MtMUlIyETiAyhoCtpvWG5A0QRhTtw8VZa+M
bj52UChus+ioW+upz9XbEP8xuZ9ZjZdYLj+dIgYihD7KUsqulppA34mqOadoBert
Wo+R4T2xg6gKG3u1+XkJblp+FVWQIVDQv7PKafbqE7dDeNxbAcpHthU38BGi4zHc
BTojyjmM6nkIkTh/aVCAO/n18yf4gL0/6K94W7AAI5c/j7lVA+cjFJTk48v9PNJa
5yP8Jt1dqXW7gTos6C1sAdmT/c99L9HScRJIsxZIjjVuENlA3DWPrsx0UPqYrSy+
PlPJnUt77rCNzm0BtVwj0nYVX9zL3diUMPjsCwzMQEOPud/aXm5kOaqEPJGrs8bA
mofiphOk+dqwoPpdV9OCnfV3znafRHS9HMtC9IytWhl0LRmrQUup6ibzO6Zol8gR
kzy0j1660iYM831ZJDxKq3XIUCjMMOdL6FINp42IghvYK3XSkHk82PSE2GBZXLbx
+UySnuZkssAwue1tkU1xlXr2WjWiC1/xRk8RXptqAH4XMxB/kVfRu3emfEf6h5Sa
ezC9gSIE4EfAb0po6/VWmnFkLeOcmD7o8y0TrX0pqqzXxSwQ2k0uggQEoVHzejjH
fyQYjL8lLaCBl6JShF+0R6vVejfGPI/3NgO3DTo0ibvH46gLWvfUKmEjpyu3hsjs
g+zLVMSuUeWF1/O2FcqgJjKssnOYDFDauLBYTzQCRoyoqT2VPHeHqAUelkGX7UN8
UEaa69osd/1NTL7SZIM7BRXBPmjWf/fYuiGcTlecCfl0y96j8EIZ37diYABiCzI6
J7RmRYQcr+/DeON3OMUjCKLDCYHSC42OW7ycgWBn6FVf+Ht+Z0OO4uuxNewiNcFO
E3dblRzGdVE1AHreAAKffv+1IsffDcirLXGOIEJ1lG5rtIoevoeC3Nl7hhUe8ycZ
EOJXRyzozYo7qSuj6TEbk/C61Utrsvw8ItCJPQeNQEPfA1AM+PywznOMhXv/sP25
0npDEXGLYr0HIUfrRO1ZB+WH52IK2XAIpTJGSrTYmiBOKkwvYhS9RSME6Eq/xny6
K8wIlUvyltqAZFSiBmUpI7p9WiBW1DeiBaOB8ffs60dCFOTpVb14ShoRRG3O0qtW
mko2JnWfARAjT4f+T+LzGYsi8NxT30BHQrCZ6FKsiX+L/kq5LAEGxkwFIaw5PVIK
2boA3SHjn4eKCJLbNv/v2P5QWJ2rCnEB9yi1tb9djF2EbGZKxbDmNmKEdnGRmQST
BkzEDjkweT98dU5gBY4vIcaLJ1qdvMH87dgbh4t59RAkC07YWilSZ0fsTTG/1GXK
JUVAuOdJTVrwUAAdP1xWbxtzz3AAGD5znab5k9XSM4xikiSwhrzHtJCEl4XgLLnv
Auc1Fmff2j1sp1enVoneVTresJlm7KvFjVEaikwhIyCEdm4giYi/GSbf+T+naRQc
cE/6mwAlBgeLhzsTiQRDAewwsyY9Ooy6iTp3ZM48W26BVPA2qih2B13/YgUrpTzM
+/ehQQsIB1zyIl4TPqLn7+geLOetjynS3me4EIGfs0xfDmxGA4vmA+lSsgZk+faA
Kwolx7fgQzoXHSPA9JYB4CO6pbKNrB4YpSBL3IRPkhcfvfpLNe8EdZSFM+bwGjrc
hVB/tChCiPvuIodQKvNjP8NfJQ0fKQMxBBof3E37KDpeyxH539mGgT4YdbSBbm2s
F5AkdDHwMn3qNjy7d2j6IKH3ak40/AeCA+fHXCJniadPVso/rTcnef12uywuIzez
dxCPl1CY8dyDMgPK8JPruxO0XvQ/ckhQRDSK6ijUSdW1p1jkKVgvhGZR7EV2egOT
ddIfF4YqjwqSeA6n5Nov6pVjBj1FilLZa/6g8fDt/ulkXmwXEqqCi9G7fHKjGMaV
UgxYKaJfniA9T3SpEvCvc0f0cNykjPyoAO4UQP4/cof7yB2GMhfC84E7C9q4ynv/
Q5p/+R6F75t44FyccbkCjNZX4SaUffr56ScKXNU0UW6VaShWP0dQhfLZlTuQ8FQm
OVUFwoLcEFMYwbJiyLDOyk8rdOX/ttoqV6y2gnW/Uy1wCZ1BZQIjQzbnrQl3ugwQ
Y+xYaaCWJ5win8TB98Tj42l1Oaz1NGHUqSvySav3+gQ+NyD9NSEWzkE4U9v93qVv
K7cUUZJn98yIMXAtAfA5M+CVvMTHYutJham5sggub7JncnuTcQxsSNi0VSs9BAcs
dL5F2R8qxv3qV9juDwF3qX1Dk/R8VFpVlau9Z2c+XyiosNO1ImTQHsqUc/KNzblT
sr1b3qNaqZZEF+kTJ7xVQMeSA+G1pek8C74/GPFzNndTW8pzgiMPPz5wNNV7p7Y/
IkBD2W9mWaiZcqC4dD1FYV6D/mI3rXxCxyd+cUMvOnJSJ6zqgZc5yQHrzk/NwL4V
2Dalkf4Aktuvzh1xG3m8QNnglojedxk1J9mNibIPrbZ2EWbxHKehDpx3E4tZe+cO
kkanfBNEtZe9aI2RVo/4RQ/ggslGYrYugWk8Vlwv1EQx7GVws5MaYbJatR3cke9S
kBYEKQ74lXUaTXSkAVxQrS3ZNlUC8JYhhaL9TvD4UjCFrjW+GkIZ3TvciQ2IkLOk
QX1lJtUgGrWHAS6fSaunCYNlZH2ouqGJWkgKaLPf/OwonRoR24BCIAc4VYN9PynN
XHQkcgmF/lOSN0qeg++wr3QSYN4JQ6Skhh7tINDZbEp4MGZB5oif320fBYZmXGOq
JJodjUp9kuY/K+4vZggUXubgvoR+DbDMiU7Hj0HgH40m5tdEO12M7vnBlzIp3pAY
Wd02jDvM/di9lZ3bYRUAbPnq13AbWzsvWAh8nGQfgrl/axupKs3NcaKlMCLptgDm
dYTOAr4HjQFIPOgQBynJQ2D4iFnaeMucv2GVSmX0HyQvoLq26MdKJlttLVTjw7pM
LlJPqXyg3CsFZXUgd4b/nc5OniHq7urhirWb3M1vSnS5hrQLh7gFc6lrFRJFmC+b
lwGSmWfU9eGvj+JPb4HmMGEODY6MdcxtmU489Tdzt4KmQF7gby2dWB0XcO27mfGW
LCkmz5zuuRWFGeG9LRfp86Fhp79DJtkFn8+W8gLPH0pZv+78qf8tSgiu3RI4DOgt
Ab/6bNZwOcAVUN2BuVYkeG/jbh85qptPxul4lU0BWbvKSUGOp+EPLJkUpAn7ikVj
fCqnBCxzH2Nh41kG1zH+xiTkBhFLm7cBlMwOxWV1K8gA8oXnCLQWIFQE83pSwXqH
Azl93x4OGZv/BWgLxjq9h4M5G8vnXBaWP+FmywTQFAefYhROUEPLFYlhNvZ3Va9B
ZGTA1dWSEW9hz6ixseQlyrQXYPrU4ZdDwaaXG01uqFgZuKqhwceg0X8YidpmySup
i/JNebhrju4oxxyY8qMxZ21M5yocWmqJq21AOQV8+yB6bu//441T0l9+o7xx8SPc
WZliAd5UQfyDkZPimijVGto65UVJBb5FlciXOEKRETkA3UCiDlbnje0aGIP6r9ia
gQw3yHBRbxCzHwVm/6opP3/0WHoF34yiFh7nhT6ZinWXJVDQ1aJOjbZXJalhM30a
6whaJX4mkczvfOCUVC5TJW5bHOj1dLglLK9wLFUcNDcMWlww2nh+j5jpC4Wjvzqq
R1If5jDtKi9j273gr1DPrjATzG9zqauRVJZ0dq8QR9Jk8V/+i4DJw+MHEkjTwJOz
o4z30iEtP3QYtu6Nu7dGGjFcBZp2mlvGV5cFCwKY5T/IUgg8e6AKYah5XpOfB1ag
LICz6E4XuqvuQuxI1i3ihH9P4ZRYBNQXqNsgoDyT2eKV0YEpiy9LsPrJCSjcOdJj
wOYjqT3+WHxjrz4+m+QtoKWO5QpGiKxcMXzw67+9yiA382Lr8eSuwxEr3sOhFyQ7
B3asTTfmQ2c1HT06LGXPnawiUoaCUvw6li8uOOtRdONRdHJa8l/l8KYs23CSKS5Q
twUmqvZ7JeN+Yy4FEzR8YMTC7BwIAvd7Q26u3ufLxXQjRRoZUZj2mR7Q9wdpw8Gk
q7vVJx39rtq8sRBd3+WloDKiBvcXloxrUpLDcZjjE/jFfZMLRkmqK+CIwjpAa77i
OiPGiUVuF9qpI/sx8/QRAOCfyrdes+DlPcsZP1tPLb5+ZehNMCdOmbufuiHSDTKT
nPg6GfeBARH044UzgHmE1wyBzCz2iQSlPZmMmLW/Nh88KR+WDAVPut93qXMNEDS0
djC7kCkncR7xvyzFaf97q/765f1MOa2aBKS4PifykQMT6jTQLfYLIMc9PYzMaQ4m
pyZieurGq016dh5Y5G6OdCpSdISYyd58Ow8C3RpAwTKr70pr2LHs7i0++RmqhFu5
I3Wy1kwB+RrN+0knxgjlvhEqsebXhbaB4LTDAkTMMwjUaUGEbZac3toWUOQ+pmFu
heCKD+T2PMDbN4r9SCHoghs3EpXu2eyKk/binwYdcohs8kDu/VZFm8TCcxPKCbk9
UWXwEacn+2x4sE9bR0lGegOuJkDCqtNaAZtBum00mujOa1AwBL/9WsXnFeWAROsI
LBtLGXSpkJ5JXcrk4Xc6+N7CmicTAg7m4qaMOLyeJ8CZnyOZaJQB++BPNVVcRfLV
JBQWoV90aTV/ENhv+wy3EsiqgmlNHfoX8Suyk8W/wd1QKgmzPokEGfgw0TNOLFEQ
2j1D8ysux3TAHxmSUZXnkkQiEcoqKjw5UDiuo9/GA+EEhDxbTDQj1W52vg5SQmIJ
ZKqf0zMI4qkbzRP+ix6Okp3+/NSN1a1OFwiFJievHd6jNmybmJbZULgHZVG3Mefe
TdxCVry7xhVzK1rVSfRQOEglo4xKnU6Inaeo6FWsL0b+6CRb2+2pGBqyq2RiBPOf
lXhinc22hWV9P4PAdx7b+3sT941rzbFVveG6P8+TJEVYTxQjsvrferIwevoNUB+B
82nKG/8PeKbu9+xnSRoxQify4t4VxHP2ygkVZ+jD6qr9Odb/EBec3rTYBMkfrYcG
4R5r+XYwtSSprGrB+3dliTEhpSCLldPiVwcmcXg0ci2gssYB2GdNcEA4bKxWdzyM
nIH1DrcDsN9kIqTmte/1NZQ/RFnf/d6PXpbRwrXcn1OPKurjsQrXmHPd/leQqa83
rFwBQmqUsNFQJ5/ZbUzBtqmzT2ijAszGXz44sCuNrGDzOIfjroCshz7C7XyKv/7A
EqW/juipnAIpynkjYBQgWe3UT7FSVKKqkI4xPqD5FmZKjJdTUX17d1z0SN2FOwyT
9l01YVj23FxNTfesU5RMA4x8pQkYGae8YqflqThnyyMatTWffPJok/xGxLIzY6le
535ys3f/cBgNPqTLRHtDQ/SAe6K9CEhtfPIPBWdIDRM3ybD1gUYvjlWmEt0cGpFg
bnsEh6oyBSe90en4TIitzJqcf5TZ965IGOMonkNDWQEO4Tgdv81Uovxgzc1i6V4N
6x5wivjGLGg02mDlPkAMAXUgh3HJmMA/MElE7DmyouMX5pc/9AsuUDuyTggVz5Zl
ha2Swpk0h0drZHs8941RQFkqoe79cpwJ7f00F9I5MY4dKYaFIMVOa+7032fL2AEV
2nypPnrhJS44TbLgfNv2jngnVZs7UGWbLi4O40aBN7H102IZQ7C2XFy+rtGrAwKo
ibeFvSBu1bg4OYlsxOhyxNWTFzELAv8GzKR8kG7sfRvch7a0oLHE1xG2jpFCrioP
9OuC6T9HTbotKy87+mLW31IqNp/+y+K5UT5SAtQKUoESqEYQ5cGv8/dAPiOBDi7x
EA6ia3aJ9d1R1PQHPVJOOrKo0BzdJQLU71yRIzH/QAwBV5n20DVCR4k3MxkwV5w1
ewqShqWBavEePItDbZl5hyMdS+v6S7dogZC8rE5JtlWo1R3jCG9/HC5wPp0tyh1f
IyqIXV0nLx6vqvcuiYTR+KieVzyRykM1tk19iZxQvoctsG8sMWy8S465+7n+hM6u
vrobXgDAu20+mALKhbr197acDYZky0uL6q0q4P2GLuLk2DZk9mPr6yCNr2+CaV99
xih7Qve/8eLVLhzcRN5hE3iJdaQc2fs5xhQvpn1tmSmYOlNbvKmXr0hWmE8yVqxc
U+HsTRRFkSsCbp3/4KjMCrHe4zP+psfEmb7E3JfKq2cxrAEJUUbN4KPNXsCEmwlY
dkV47OJvuvvKQ6Ay27qLnfCZT/w++jpLsx4Wu9NzZhfMx6diJN3ymj5N0JvLPAQL
NqS12Mux0U0n4Z4DkvuKRQT6eDroo11McNnQ0GTBBpaMSYlEWJV0aZ4c9a2SF2wm
A8IotTmvM76QUjMw/C+0g8cFZVZtiLr7GL6QiqHq4j297fYd4TnOQbUkwqcgdlHb
y0xLY5IZ3IsJDu41K5WfVj6uOrvvSq0DCjts858GdJDbf8hqr/LjZX8232+hycOR
mavekZSPN7eYPIvVG6ZGTU4nfPYLL4hHO6Z5XG9YSclgt6U2oeXfOuWpaUVqb8R9
F4x+KEhimGKg50Jr8vaJh3ReJTojHB+sCfwJ/yMHybmsKnCHZwSGiaOFb9LZhgC+
rQgRhEfDfpW8B5PJSTv6BQCZoRizSId4Olau4S5sRmUisAOgWmMJdcxFktk9GRBO
XII8xuRqbcLxTHnuu3QkR1cMrurw63ZNL8lOmCHGYKVbbEIUtu8nosj2dzQtHo3y
Dh+tIt2+9z9tel4dr15Dj+vW3wdNM0Qh0zlRoIWLqoK5QEJNU/XOVWQKaGxJ0TTs
dVVuIevzdXwrNVOf1BxvpE5pHoYxM4vSCZxvVCjU+UeOGNQzpU+TP5f+qmvZcMEp
RpqvmlHUwuVFtrMy0iy0suX+YzTriNTL9tQMj5YS0sHAyxpngW931cazJpoeYZsv
BBhihKnvXuK6xd+hM9Ce7piTABwvvFJyyewWbiKkYcoAhRuxxcvWNjYC6/KDO/sa
67EVfSd16C3nlWklq7B6l6tU7W/Gv2nYovFY2WrJU2L24QzJRQsbfORYuqJrRGXU
0Oe0HJpeyf9M3iEKJp39WD0oO7SjC6LANY+0hIYkJ9u6XYcEUGM6UaC13i7sh7Jz
mqm6+9QOOjWh34rWflLfUrTFklU0VFgcW8HX2gvc/a4xDjf+HMgBKoMY9coXcT7w
FDElzfjxo37e78SC4o1oBdDikAp+3VfvSRadk+U9fpuyOE0EzTJCxd8zx3mwpKFo
NiDjtGQ29CKVk1faYIRDjr4zVM/FcP9sU0/eTVu57rAidc6gPLfkobHoiwZk2Pt8
jMgBm5eDmYqJYrqxu0DuD72ok/Q5DI4am3I6zuhsdi744vE6fGDnM2pbElMx4rIE
tn0iVGDGyzAFyn9o/F9vnoi4Qd2S4HdQC2Wj6PewF1oNBTGxvVkt9AW6TkcpbSQr
pwAMnZVdrMwF4dBboI6+tkw8wSdTwpxz4YG8AC9VcuiMvaBzluaxZ8Ip8u8xVbu/
3WEcnk3lFEk9ZbN29h1uhEyr1waXfBGO0shzVWwsbL4l+PtzZXZzdYprqwdocYun
mwsclN+r5WPX2FSaB5meYuTk9hv26RWmdFpRfBr4XNqMPOslzSXpYjyAdpC11v6b
hyJKXxMxYKz0/WvGtFViTUoZeewOdLRC4FnsusLOjDih5z9YmpXSHTvyZbw4RJDu
xI26YtNNBB6I76Gq/T7ChP/GaTlTJr8tAVqeBDMfwKcBijPjHUP/wICGbrLvMhWU
0Ln0484jaYAMxBvDy0d5Fyr03u5NlIzEdhRGi5f59ldVLKPuJdoF1bWMg80FkSh2
Nai0NhIf5UlruI+4KSvz6lBYCN9iLGuwR/V+DIJuUISvDxzvxeS8khQ9vXIjVDyY
fNDL9CLfKerzqBGivZi2HZNttvBP24dSn7MkDT3iOae6+gNxRGnwzjU44w2AYLEj
vhCpRSEjrQOPrhdScSlwDdL4CQUwlm9JLYTcSoC+DOFRo91AN7j7BcjrWIsHGI0M
yMKdFFTgmKYaihbzetryRNygkR6va6nsk0HDEDiV3TY87KS4xd7v0LNraoSokEJm
sFChY/wOGlD5PzIzDHK6tgZZSJm1EOFjekn+3GuVbtZYSejfIQRWolOwix94bzkk
ZgqsgnHaYjswmT3j9h2os2JLekZsQWNie8dZVKG2OpEsVCdkK9IXTLF8JiMwX1fx
z2ZRV6WuSZOsyNUh0VZ41shYAh4Gi/AJuS43G3otLvF/9K8B739fAOadgCRc1YEB
Jc4SMRRzXOXJcdluz2TvB4PHHR6CwxlfGTgub7wzGoqtmYuIX/GikjQ/pQffWrMG
DT5RYvODDsibfIOq3s636vjZPuMRPMCUUIABc/FmtsFtrxrEV0HvxxpZM5i9CGOp
U7DqRqNRjD3ytq5ftrSFv877vngPa1ZK5EQ/ByGJa+VMmDeVLXUL4NNb4zITTipv
lrYkhunwqeP76xrNmrcbyaB79UzCUTVhigROU05h2UWQNKXxBtvt/2WNlngfaFkW
xu8/eNYxK9UbQU1TQvAPhYLMqOwVxv8DOFo3bsHpuv+Dc08mndZRLMG/aHI2LjI1
JIStf5mkd07w2lI5jjfJOdRX/Rw++ZnVJd0CXRVKWbgxITusYwfASAdYtkMjyiUj
nFzs7n4e7bo3iEHvSjYz5yZhyErLoFdE+jVhg0eP9NIUhrqOGIylQ99Pb+RQq9s1
`protect END_PROTECTED
