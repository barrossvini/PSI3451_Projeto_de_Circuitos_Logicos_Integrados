`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9rfqyR8iquvMYv5NimlrNl9LjuPgWdc7VSrdrOVr6ehCy8CeoAyeUMfcsJDVSBwb
C4YyuwlLFs3Hy68qz+o4J6+86RCjNyPzvU1cLSqARpFBBFXTeFwsXJm0c68/xSON
mPA+tycyuG8IGlaW5Lp6HwH5eoji5KThWgu2Tby0eLVSUEdvhq1iXhbSsZgsBoxw
tOfBTl/dunPFA+h8+00Ri6JBP8fNy5aRwf6ZLl0O2BD3kMa7YjEd5r87wMU45aFp
iZFe1wCQrF4ub+vC7bvu6IsXAesNx4OqddNd7g+lgN8QRmMd5+0KimEeoDlYoiYD
lpWjy+Oeu7pdbgmxKtej56BKbnG8yuV0krsUdNZ6CvU3LKwWBT5jlriQl4/HJvBw
DrWZrwJwZdMOfrPRbX2dvyu2i0E4Or5qn7+8kEHEffolnIyu+5b0LFw+UOAe219K
2W0CnGSJKVhHqYcRngt8AyZtLwSQkDxl94hvTv5j/BeClcAub3Vf+xZ0VvWERx/o
tdoogmfhz+u3wCgeFpCbC0Zmc/iNQtxenuff9mD5uoOBRhJIlJf31I7HnPIGKflk
3M58mlEr/GxDeMQ6mxp22Obei3MZwhMttVrDQEWPOUeg/I8+mQCdKI/ZdS0IzNgm
7FEAKa8bDEQ1BM5bmIFUgvl3m2lTwflDwhj3XeU9Wuz3IYqZiwa5/z7skr8sOaUW
H16GlL2M/eCahmiCn8LYNRMxRmtSea1qWEtmvMH4Qn7CfxicCvI6qTr4I/Bt0z86
lABXxxn1rWJn3Ekdz0RfCzExSHr2LK8HZbv0fHSa0EKo3DERq30++ddr+f8orwrv
jwDS20sU7yceK3ObUPc7cb6GZlZfAFqoAKTpH0UplzollVENKVMLHXqKGSkttQFf
hjsB25f556ghiVaW37pX2VRkPu8aAFxtSRJiYYxhOYHV3DSlwMlmIjbGb2Xvn9ru
pso2efI19LufDQZdOP7wYpC8JsjYMeFlurViIP680ktwVXyKLsoM59bdIJsurDif
R32/Mhr8CF03R1I1WyR/MiOp7qI4ol+N6KgVNGfCaPfff2KkL0JUl1vDYpqf5H6L
`protect END_PROTECTED
