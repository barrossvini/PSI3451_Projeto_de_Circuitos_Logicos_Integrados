`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+NZb0R14UgtltLceYPzH+QCkUqV1BZIfYMu2KMIKzXKeMLMuNMPnashu4++N5Mj6
CA/KtTdowgAXnPkgaoaq01MqKNZerNarCgiMb1V2puvAtet4Eotc2aNMVEsXwHST
fj54ldG0qaJydihp8RXHLJ8Rjco0DxX524ss/msaKLwCp/q2YXlk5TfjNRfgwfiV
ZfED4twOFaub0iG3JzycNLroT8zB0v5btBU05EUeGji7RD6gZOLL2RQKJyqen7Mz
ojngRmnAwxLjBf3aqXW6bXUVWyspzKHo+7G+nt5Hd6gJfwIR/jiTaMKfUL1M1Y0M
yjUi8BRM3BW9N5L8BQ1Wp7sJy51lSJCqSobT8HZJehqyfMjL79hgdFRWs7XxlIOq
Y13ueFjCPif8/H+/h3XKp7cKNavZ1MXGTFGJc+LqkMNdTKP27OAsWlLlpnyptqfg
8VkkAYZR040t3Apevx9zS6R0rYn6f9+L3gIVUldG7HUrSm7PuS/bp290otLaHzAB
sV8jNUI7FcVLOnSR0WWDX83Lj5RWJ1aw9hcUB358dRyCTKcrQ+gDOVWfz35h3m2C
msZSoX/XTYUEtrGRUvZ5CeJq4ZjuPHyN/x4GyUqeiDaopoTNKlctZlzs2d5rtUog
/8jkFa2Yv2M9qLkB4ZFmwIpqYFaVNv/jJgrOaoqDrM02Cc6dyXe5pMch3O/Oz/V6
MY6BliPyemu90Canca0iolmr6ngsC8n6WgAidDyYGGnMpCKEstq4SnD0JzZ1yhaV
6GZyZvW6UHz3xgZNJgClOZRBKOE6JPd5mN5piuajlv4z/XE+a5SwHUViU2HxaejN
tMY3jiUtgSy/0ge1WVZ0tlnXgnl+A/Zt6cWX87WxQ1fbpTgJPTsU+0Mu3ntFxHN0
v/LaJJnjKprtFX7imPuEHR/rb4fydv9Wd2Ndv/RObWAXxuGa1Lo9TINK6OqhAk6x
qHqV/JtkZdFhj5qxt80xMn1x6YLmwLS0TZvwuByLPD1GkT29XyBKX+O18Q5/ALR0
pGjbkBfaqw+zTCY8xLAXXDyC3oZFxeyrVa52LxBfYOI/cK4LMN0XAdK5VAAHLGTa
eZ3r+iyk0xPnObEcxJwTE+y8QBS8V2i3CI0Ei8FQX8qNTU01mOFdNrFEt7NbU5pw
Dgjxpu+BKiD8rcYKSHjMLXGc9Uq9RQrZYDmiZmGhOc/CItnfRv3v4EF0Lm+EbGno
yvtClj89TOqyRbwfw7nYdT15Kr4Gnzc7oCX/PZiuFwmY22igympUq54Grpa2SOCZ
UbDk9Q2698gdqxl+lxQqarUtv8yslqe8KBkINC1gkNr/LwKVhyXF5JjHiDknY8U8
zQwHNxHOdzEPakRXV1uN06HwckMBlQIVVA0VAT6L9VsZ/NobsRtR4shn4qa1ui9z
UQLm3VnxJArLa9VCE+jyj07V7PJAxw1QSMVfQjdKTF6Mx+Kq0o/gnpeuDy/HltPe
`protect END_PROTECTED
