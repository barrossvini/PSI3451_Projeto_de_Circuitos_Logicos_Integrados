`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwPwWZT1xnYkoVPsXUYg+4A07LAI1vhXcx6e8iKUV2HYlTYazMddFacCmVLQfVcI
58sUgm3OADwJ90B8fqtobV70AWUvMfY3+ib3nVyNDxO9UmDYgsambfcVaNhOr9JT
qrAwJKp9j7daKs+uidAcO+JjzdjsxziO2SBOnvg57DPs6f08L4sYNKA8jOsReq8M
suVl0aOAoqnzOuwOGZ3z/4Ylaxj9RwaREGeZQ9mN7M8n9D0FZRSpdm2Z/3TbxjOd
FHdiaB0upDre84aFppnoupOvjHVvB0LSeDU+uYccZEQKHlg3rJbpI16BCjgVezLP
vzGXcUrQt+2LfcET9L0sSvBuZG7WlLDQpJGiu3Rd/TNutOBrkJ7GltSQ2QIMuR5U
egfY941oWYWRB5E1T5oL1sdKzejcwjeeIbObzAxX11nUeZY2mnaUcfKjZd0pqUJs
5rSSN8OcSB0UELbvhS+kP5KKbirallBuLb59by7Rj4wqDrB9M53vXjZNynl5FBY4
SCWccR1LbwIXsE24szkW8tNNlHb2N2SlLrBNLlLunXoU+K2ZNm5aYzsSNas7+k5D
yECykvllg4TxRxMet6/r1M4F3YcLDw8sGr+QqD4nbXJb04t0ZY/hg4lDUZQlRTni
bslvOs6E3/Z6d17AqjV+P+B17BcuAKPzq0hhmRq8wctnBsu45AZZIITTrYBl2ynD
aO8BJ6va5Ce/U1Z8QTLQe9e8j+UhKqT3eXnMMKzlE9b3KbdHxCGIWIQH+ZyJIEUl
sDJk0I6ZX2lR5I1BENABd3Biurf6k9Kl0FAvULFmEkj+GlI1t7pENC6s08ID0h+g
v/0uYjTdBdHoviMAvri26pJlFG4Q5LyWcjRGcRv/Ld4G4SsT9enjFJEduv//pJgP
AXHR2MP1uaxFEjRGMBr6hHSsOaaM1uzVpbj/eeHEGiP8igUJeym39YFDbYXqGI0o
/spy2IZ2F46qkDuhixetZmcQXwD2i58utHrmoq9iXtaijQl+eycfNEHx67gEIV8Z
qmOTosZ4lRwJYe6J0hfTqTZLoPIuJQL6criJN0OQPAla3FKPLg+/VRyo829809GS
3e9ysd6xwqqy5l8/lZq0Wt1JcxXwVC3hhfVbCdP1eakApKVCcwwRYz9YhVDOLs30
sYB9LOwB3idi127SbbANX9JT0ROUVPnFiv4yBCUIackJ44snKXWIZ6m7txRmykad
Xlfpt58E1rPk5o0OorWLwenFtd0kDkxmUpHEFHypiPp9vry81DGvK27PXhtXn2E+
CtpsUu2n+yWcEtB9Z1mew3aQzqPKpIWRPdoU9BfDknukGxXZNUolfGJBBfdaqar0
6YWPvHXa8aVc6pCLbhrUJt+1DQfTm4hQEGqrjZs9/9zM+UaXgFOwN6KLUWQgydnC
8sXHP7gPhK+zLljL/Ogjcil3awKXz+ZAk+Li3Np4YfPTqfA3DiGTFEUmIVmELOA2
HCCLuyfQPx7Y8J0i31coXwhopGvx/BMpXKy8wxxiH1rhHIE9YbCUHubRrdG1jc0r
hQUCtNfG7/S1V/poSP25xksVheoeSVl94zZv+U9Nkng=
`protect END_PROTECTED
