`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QCveHaohOzDfO4mHDS4zD7wY7DrEouERIno/zVvG2fnxkSIg08Mzyg4VyQHKbe2D
+GWlJLCQidoFuSP9/rWm/XZmjI9mOKrBtLtjO9UweOAnLsA6PK/LJ89PttpsepK4
g3Zf0pX2gGmmJx44XBCG0ubu0QdNq3vYTgM/OLEQ7vhyFKOSKi9D2cSKocUep+yn
pczUt8MPiRjJ4UdCSdVoTdiGl7rJcMYEk99/J1PCu+Hi6ToG2GNsGHDhkrlhX0tp
wsZiD28wLWY/E3AF804wly6sF943lE6tub7txs/QvnpQnKnl4T5p1wme/v5z5Ego
0OJxhLBknPJliBP2KHyx8bo9S4PyUj9eVwzpi7tJ0+6nXZ0qF12eLRY3SCiDQeLs
uNsjBdoIqS66Ah5Y4L7ztv7vfBi8TDq18l7C8AavjcuaWsahia0G6EVUiZYat0Ko
8DXSap0OqU4l9NVvpj6l0Gy2okyheBHRxdnmyTU7p2I1VUzUO42hYfRTLaHpdCA1
BdB8fqvLuhLyBC6JulLFCIrzoKLBVnO3E9qoq1cUbtCtrwL5f5ZZOkdw6Aq+Kj5Y
PoYCfjIGDN5Naks8+/7ZFAdLP/C0svWGb8O8krHquJdqRj/Upo9adpOYOWs0LLCu
pF8ASWhQFq7UnQRh4dU6qJZefP8GPJX3YEEeBjVrZcReXMR0m6VBcO8G06nsE64G
ZXbT8ZoliRVUfUcPLyclKHGkxESiaE3a4zhLvXGTrAA=
`protect END_PROTECTED
