`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m2FnV96OIdjabyZ1WIc4u0RAQID5LvTJ0insXv2TvoL8GTrJFUXN8TvXIr3gh1UB
OFT2Vau82CTeedygA+5LWdgdP9of2NKyNOsqjv0fZpoL7uHrT5lAuvbCKzBMAEnC
6TcgDnocjINwAX5s46k5UkLGLsIHO4GS6X7iYABMiwWqTgtRpXhlPa1OGCYhGqM4
HgwfLg+y+bwlUF+EroIVXQg13E5k+TqDuhRMGF27IEtUOWI75AmdgNDTClJQsrrc
VjdbzGWkUyCf9orYrym8xLurmtmqnaMFHWOnfXcI/gUXlwCLrEssuj5mQ0GF9oMh
CC8rRIer6YLhNlooDWqXQZMER8jywbXtDyhn6emXtMaiYD4+Yp0VhboWhhOF/kVA
NY4Zf/z2qvJQ3jHsrHkas2wRF4DgfXRaA0xYknl7tBkYTziygofueaOFn7QUXFRU
HnnrmzXBpjnvPA7RciTT9cp3zEfFHs8qcswt497RzF5udtiJqSUS2nPVgJfQXwv8
YcfYvFf1tuHpQdSYsPx5eO6L4XAjFCJHIgKdzNPKjwV+QIKd1bY1gz5wWxnVMUOY
`protect END_PROTECTED
