`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sinE6+5ogK4tviY4jQVCA9y5nKCTdnsYRIpd5qTVMeIRM1UPgTZTOg2MHpQslnhW
mtXJ0ApYNh1CLT6Z0qk+o0UumLLR9qTK8gZepABtzzWN+t8FDrnykVl5rfB3a2eG
EqeCir7yIVkZFQCE8Z9uRNnCeXfj3k+1Be2u0MRH50lcKAzN2/qDKL5J7fqIMYCu
O9tKfdLJACzjSBG5mZ2dQpYV1sXKb9ICWHR3T8zPCSRXgCoYAdPCbM00cN+XqyKx
VQ3WJvXYu33kcsY/mnbxNghUZ1v8mX1Rx951o8ZD21YN6ieK55fpiOyoEyjZMFlE
aWnEZoajyGI6GxOQtl/UP7CbEQ0shzJCdeqjCX3zS4VhenMUkWrSfvSbaKZOT+g0
TeheH3Li7F+9WdaWgZq3Bcu+6qW1kwAzq3mV5I21i5+I/4Mal8MxjEaBS0xp5sM4
fSFYsJQ4PIq5ylz6FfpSG+3y4XMSz3T3vXo74iQSNMGxHzsSATViLbBauoun3PR/
jdxe/RK58PN8PI3bbB6QHzUKeYHO5cocRMidJv/NhshTP+4zXVsXw/pSP24whIxc
LOVHi/te2qPl7hT+CENlT2MHu0HWjUpplMwsQ3NOk/O5/SN1rBOu3sLd7Uw5LUxt
L9j+dHCjwRIcjfp1WLtXHGj8sqE/bw5kV+bnm6TfNyys00bXVMofBSwK6f8afUAk
O+fxAozC96XZbkrymdGuwla1nGGeYZEruz/CT8rypptFm6WFK0+tvcqB6L175bEt
h8r7BSHUl8IMoJFOf7pl5g/BvndGy6s7F7l0MRV9Vbp0THSjaXDBXx8y0BazNqGx
8ZG53kbkusbY2zhu4GTTCRrUoToeKgK1QiLbD8wb+5ifWMVuPjksOrW+j2n7KKhV
lICSMRdpHelD4hpfAXlkjB6lwJ1uad/o45vXlokoe2PeS3WBHua3UF2wB5azwc0s
0cuNtMzpNsFdn/3d3fHOOMlh17wOPz1vqFGz9QgSQWezqrVX4ILvyY+10Ja/3ZRe
TA4DAMSfRmIITLiK3h31alTMHDXr1PHTJUTxjWDXTjy5sis8MAy1OMRqZS1bxtO7
klXBN+hVhRGzbv9+NU8XLzFm2BmrNSapZh2iBF3GESkwtqhkGv0d9R57gP6uy3jr
pO8yzgF+55pV2LlGsuJ6+jkOfuJ/+JHCJmHWH0TyL7RpDeCsioLp1bJdi9I4Cqld
VR3bJa/3rnUfQMZ8Pd0clsaJjkuyf1EwgUR610oweWMYUNHmGdhEdwOMU6TaSLLa
x9HWqivnPaZJEtcJPmp2Mae/wQ1bfVOaRFsY3rGO76os2CMQfig5cNhtK46m4WQp
hLvb6V3ICmAf2kcuUmdHOM5JHkW2dRSQbuH+pneVNOYTYqZav79m2owYnq/2eL1A
cxtM9rR2FqhJLxgvnZLTJkYZqlmHquQqICqvgqDzeQUhcV9vJN0dc/oqAH9vS+hU
eQoOq4su9CeeRuAo82wXzwgMqbBHhOfA2LNZHWGzmtk/otVrFtI83k5ChqA9uu8O
thcqo3bS7BE63uDmgzrbPGKV/9m0CmaGQT1UBF2X3vGIio7IvONsShwMrKvKJvf9
hFW2Zp7Oy1Zp33IiTvJyAFxuZKBP1OAkC4fI2ZDmM8ZF5Hzgwa1e1CICtGizhTLZ
Dm4FEuo+eURIk1FBIF2R5nN+IBKOOddLK7PH64DDMMnc0s0opBl6kOk27tQVcOnM
NoHL/vXc0Ryn/eJMlf0vbL2XKnjjNOiPLez9Z7LxPVn9Yc06fLFDfrxgrNAF3f18
HQd9wI8xXWefqiTnjX+0LXbiMGYRttJaIosv811BJwKvFLWtAtFrX41oeQgsb5Lv
3B4aA04vgw42nZP/oYB4K0KyMlrUCthaqWtvqaPD7H4YG3DgC9g9SGmE1/y0QSLU
uOtKe4yPE9m9QbIfJPjByaqib75glQuAzN4m31nI1YvQcK9HEv0fnMWHewBQhM78
jMk5KWWUdvXRLJMDzwdZS4qjV78tvXfu/dai9EqzeXN+gFM3xO0W6zACeVBA3r2Q
S2Pl3DtNfT7eohiNWURGG9AjYRldRtaPEMR4kAnWKn12PLuFYFbTpZ5P0CWODSFx
I7NJv+dxMa7sd2CWMRxiYousLZpk9/e9pd0JjIwkniSR7d+xnY8reIceuio6/Cb0
dpn5ZJG3Qvu8DK5Lr4GBI3hHV+OkZ9XGvqTjXNmfh3lxyYGAnK5nL9gznkrc+2Hu
Y2dvdoCXeVy2gXU3bNV1BA48c3QNF+zYsM69mpHXUe1o3NVRi4iKPUuvRqOR6gKB
NKyeNSvZfb9GlXODDI1gymp2E2wTEyI4hCNC+xGYQuACa2ECt5qRoGZzHPnMOWiW
NVygY8IpBPmjuQmaotMsCdzxxKgHFpu2A+EDwmRRiYNIdrVhFSz78sjkD/0Nosv0
dNJnOVc0IgiUSxyHsaSqZCJEy8NyQisSJeqqapXflDnt0wFXaQ1D9Rxinz5Q/ZSe
49h4GYv+S8dQUx66hkCZXqaAZWAAECym2NpohYEl4NtPjFzX0/LTLaAbH0s10zvm
qjxkZ59Uk3DzI7hlSdCW1fihYvXpzNDYZnIX41ti7+MK5x5RfYGbdeXWtKDYhmi2
xFtsNWmMiQGjnOCO+i/vo79b/360mkE+BXHNDXVDvozwFY6Olt1N+A+lz+vyYz8f
TMfVN0x1aas7WA+4GDEyF9xKkQpNAtTi197BTO29plo4GPSjMx431+EPHVZDtDHq
PeuaZPkdfTxsPY0fO0KJUmhvK5yk07Yl3LcH00qv+tz5O3poX6NWWvGwXuj13ruY
1jorhi6bcuqyO4vheJhlfjqaT3RV3MVC78EmRNE5Djgi0EldcE9f7QLAAP3tgzBa
AS1Xk4Z9u8GkV7JnSiVxYQJoNbmnnfZE7z6pfwjEZ66Lb2uu+DwBxDy9Eg98QbHd
nDi2QhhvhkPfmReZhZDF+XiZvc1A1Hp8uhi7MP6jjxD1BoofcteFS1Vwn+owO6oY
pfYwOdL72bs43pI952xxl/AdV1jw9g7e7P1Mje7sz0CK/z4TCloW5ijGF4c39o57
ckoOjitHfzEEUzqpmEqBtYGcE9sr6lWIErhlRebJ+svMZs/XI+jZacI3SfQkLE0i
h7WCWkr25DGkx6I7Hde+CLO3xiLZEoWLiKRemWoZ8pTmHVc1EPmy3nJsKnkD82hr
dsAcLxsqaOYiG/KvXJHo5Lwgm7YagrM3NRF4DVUCzEpEkjkZxQhEGFRN9/WrrmRR
zBE/f7KvKVUTn/CO6su9hDO52+a8kUq39TJA45QIytUp8lnlpEHGfLMS29bebFms
FBv1nKqvZJGyredwusoV0Zn92WzOhyrZpMjyK/a3vV9HSwFuTF+hvxfG67Kou1oL
AyN/5TUfTll0uPHEdC/+9QNGFkQ6hXvbNkYqNKprMpsTfbnPbYyF+SdoY2CVTCqS
L7PZEu9eJARxZl8arGpZpw4EWwA6cCVh0YfKNHphnTntGThzB25IUljC01/Bc0gA
HFWOy356dWVIC85t+8JJobmr8kN50yfidRnP8KStP2rC27jJPEWQIosLio4NCORm
/qUO/EH38xe8tqFlLTfqTd6Kgz8N3Bh5ruVumHZ3S2Bz54VrXQxyHQ1zzsw6OQD5
SYwdTaOj1Ca+LJ1lOsG/3r/2ukD8xq5JGgj1lhHLKZwKtDStYM1Eke5iAYTf6IzH
ZXvavAb9p/xTJJprMgkRjW36v3eBr/7O+LgOYpjl2vRxhY+gv2LW/a4EyrGqxsUz
W5xLyrDxdJwkgzHz0VLcx+NBX0biBZBD9L181gPw+h3jq/gETGG8XnWTvy6tAQQg
RRCYWhleDF8Pjl/4/ETrbPhG/hnWs8LgisoGzG6olaHXrocf8BgmWGheUHstLsIa
x9Co7yq0VsZQQj4KlUh11a64oMcW8kwqNBa1ME4hRZK/HgMczYri23bTwibkZ7RD
TsdYZgJPFxUMylxPs0G/I80F87MkGwE1oFjxA6tWjvMLIdG/xHsVfGh0K97B6PZL
HHtqwM3mid9EXd2SWmAqyyKueNWD0vVNHrgO90aet8/j+Na9Ghs+u/gfx2djv/YS
KiFN4/0O+ro9fk+AYcHwwKzGrGGbSe/m5RQNtAUmO0+hbGPIjDt2XK0kkcC92qfZ
4M60/ZXR1MIRrUUXMhSE7wttJg2nvcASq3YOEBT60h89gE11a5y7axqaHEvd04Ta
pj0Yj9YFHXBj7ButmkhHnroPkNYAC5H95UZWZ5cnjLoRkpKGvAgOg9vefRYfIWZL
/6g6tQ0ShgHw92kyBv64DA8Xw3jcVytp4G6X6uxgePMLxyDmHS7v3jabdt/pEpph
iIutYdIHYx2akfV6OLUMuC6C9nFPFyLoR0tKK4vnXi+ZclcNFZEwIhuuj2A8NFpy
wB/bZ/LGF08ocyw6dQ+XunH91xXI2SIXiwTwb8g0irCeOfFbx/tQUTURg7ColbLj
aMoZ1jml0mlIgGtH9bYQMsh3uTisBj+aF4LkyKSocGiV53USvZDKHsHcljI1rvrF
DvFcUs2+m2TGwJUmYbVHbU3e7LOz/29vxA4FKZ9V2CX/9yLU0t1Qmp9gpLpL+gXV
FbzYwjypBgksqryiACICtqnvhUpD4g5vEnJsMBVJue9LcCcAUqO0rNQrrlethfgV
eK1NPXZ3tWdoj6Sy+ebDwgecBdK8/JlChQPAkx51bkjWkrwOgl+GQ/9CFd4dzYqt
wpuTXfxvVAL4tHLGOGGy8X1khyC2mtVmmVDDnCiQEgQPcrG1WE5QQXbUxcP/iGH7
2JAeoXvgw8V6kitqbjGHWOYLQ8auBoFXJEEw35DbxaRw1DU0soDHiTmM1/v8O/Tj
t7LJomWExJ7+h91DM0oJ0AAt3qtB8hIYeknpWDSbE16crutC5CSfBiEkPRJSqXn4
tQvu5gm6zNtxN+BxxOrnXq7xnvJDUx8UafMspqHRwYcqsnj+xVJ80Bk7WthR/GXb
zPEmlh00SntC6VC0mUAcqJfDzcYHbuicJOY82rdIqc0ezgJ5TdjmfH2uekxa5/J2
klO8hpA0OMZsYeM0sq820bJw8vIU+pHYI91jaVC3K4PrwPdCMSn/BNTro8FT2exC
BHI6YP9cNLLZWUCVTuvW1Z3YLUiVAUhP2k9YytuUx7XTyIrWFRRGEVi+GwYSDn7U
gGZrwmyFUsXQudFmNNY+scu/5siQ2YkvLtG9ixJK7pFwelvoq68+dqPhLw8ufJgc
WfOQ3tilvxltTiGhK+DVkxy+yCg8jEeW63t+MjvDSDRUqtEJy+BNi2XRCHqIX2es
+5vnvJ43nvt58v5+cvDu8rb+wuHsI3457bx4TT85ccvW2WfcTS1ZjOS0Af/be/fT
jf2PH/17pgJR+hBQU2lhb+v7ZuV2g/lY4mB9imdUTZiOJni+CUeWFHPzVxoPnS+6
R6CAIlPlq/dtsziwx9VcwsFpVxAZkp04eTaSR+iGfPgK1aFu5tTEj49sbnDpuC/p
zApsjUdU4GBBOxXplvsajN8XGzNSMzEKvZAugdX8fdyWFgiBlfufGrf2hyVK/IiO
TvTyDBG9lLsP2FBIN/UvjJZDi7ivK9Md9ZaQkUhAFrCqjhbePOY3InbfgN2mas+u
qKhPOT0C7LJ+3sQ+152Hy6ApfBQB+ppCoc060jR0jC25AT4yQE/v/2T+xxoIF00a
t4ltPLhDRUNodxjBqsz/LodVfreHJ6jQvt1DkeFxFRC9t3CsuPFY7+28wmYt/fl9
oTpGCM4RgoS7otfoU+eOksRA2ZSWSrqQVUm407qNj6W8r7PFpyyGF5A26wbNQz1s
kqHWH+UH3GD8vesnRG0cpHtuhkWPwUXIcFjFx0p1jLZa+JOdTub35tXKx6k+UaV2
4nM6pa5canedA6XpQapvMbYUsOFbu9hHtDlAPGl+KWZqM2cnqpvVab/tcIEHB7xx
TcW1Zv3hApn4TPw2Be5FkTnAfy8Zez41cIcQM50fzZ7pskXcsSIA+vPAVNaJ2H3q
cs4PjU8P2t6NTNIg3DPUuQtpQhe1sHU5ZI/lglWoJHWLN2HLoO3E1QprjOasL42s
DD8iBY01weQGQthnuqllggL8nvqZZ/yHe8ekpYOYlMpF8/Be9gynNxXSgDrshWWz
96ggVKGz37R5lbia1JSVbU8MQFilhwfNeNGZLFauv1iqnIhgNoIFqs6VzdozB418
C7of0AQRrYdyJLkVxZY1x9lWtm39dHC6IDrfz4zerfZZ3oHClF4WVVuzdSlaH+1y
pBfCJTtCev7sanS13RtJeURpzlU4z/h+RXoJcQy0thw6olrO4on6WSxlrHnFPgtq
rFLl6mxtBJv5bl3MWRq2vexY1xWROKfDgX3Dp5E4hkSR7QM4nwYdtzQaLLEhjkda
ud1bWAFrLFser7FDy3w3OkIGQLiVHwZD8dghoCCaKjSDSURGuip3LZDN3qplJa8z
tNI+b3yD89bVpinEsPH3/1KnrMM6s/fOQ8kLAJ1tZNcZZk4aMfT5CxBdKLO4oSS5
8oIJGyY/ZJTTQif3MgqTFMbMTn5JY2RQ5HKdmCL1yDeLNnvbXI+icRAjnfYaA37V
XKawItG1S/G6GPMI+3oAS18J6qny8DKcYpMLtNTQhuHfrhM7MeTpmq4w7EIFyJg7
xy9X46LB0R+Rmo7jktdLPLXFr7Zr0EM7n0uQdpiiWaW8cEne47bqKPJIhfvjC7zb
F6l2Yu/QkfMsPZEGQ5SvoG9KzjS05PBtZi9i0zHMesfI78wyZdmcfC8OfELzTLPt
5H8TEUB5yQb994n33sPHDXlc/MwelJBvCv2Uu49h4Z6nvkzMlLGtDsNPBGkRaBxT
J/PqmvaiEH4qd9miIZ2QXr1Wg3ybbc9lhpTwa+yDXoniMTYg3FDY/1bwBN9L74Kd
/JvoNYENBfbjSfqOJhWfwq09hHz5IAmZLcFz4OHRn8uSlajgnb1xeXCjUl4nL+Vh
yQr/RoHnoTKm5vEXlTzOqPC2Zc8pv63YfVmYfwp3d7toPEU/WGJqb+yHG3Apt0W/
TWjsFgcwzpGuCsrtAdQFaN9+DKUAu3etDJcz3RmR3XOGxdCwRPipqzuecWHRFTPF
mn0WxeATEut+1eKmG1ywOnoQNV+OZSxdEkG0KZUqZSNsl39rsZo13d9jR6xNypG+
2Di2My3R4ZEfWgTWLrVQbTcP4f0emcFI7iDDcNErS64HguLLz/ZUhCjEnq8ViOWo
GLk4almpEB0/OskghCRXSYjM0OKdc41pNQr73GBkC7ybJm6CPU3sjA7q+gBGO8/1
Ql+jZpyjIQMXZzhK76IQPmVmWqblVgZCnmdmpDqIbWX9BrabTnFYc7CXaOzg+Vv4
EyB0M84SWdPosd1HN+xyvr1xZ7T7/qv+QZaZOB+SZezJ9DD2Ikv0a55pDILeE9NL
9cms9TmVFj6M/bemoH7975eup1sAtytOAWhoFqu2//Lqyr5fKnZWv8S/a+/g6Fjg
H9ch8Ub7wpTKlU8XPcBem2/xVvkUHfSllthizdwTdEDTKulI9P/I1UlW7M8D2bRu
boh8W5pPUkle07QC1yQE3XM4r+48nefr/Q+pr1898+KMshUUfZQXhtgJ4GOZbprs
npvfcBf7W0WozvDWItER3o6dEuUQYF3RN/YweG7Ge0rGYxXXNBALiSVF3fC9iMZc
PSS6K5TL5o7/keFpWP5c3o9K1uMV6LYXc77pgJ+JCAwHD3692GZeP5VH6P4Ya7FF
Mbv7/qxnu6Bekgf5TUyFzkBWw99Oe56fmcY5IiLJ37DY3MEEx/71vN3Eu7TGMTRz
uwHvpkVS0N+syaNLoh4/M1j1tv/eTGlEXKScCUuDaLwnHPU95KtaxAek/SFvOTYI
r6DpSFtdn7V3WpMI2g2d7TS86FtnCOfQlZF95Fu9JGMHr9pZcYma+GTPK+uZD+xS
Kqf9h6DKAfu0d14WImCIBtl8I6AlVjhu5hIR8oaTnfTCq3eausKoPlCfGAPB4JWK
+UnHJUBgx2CNhfHFb7/nQHXVsiXvqrVsWrRdsyH8xxCMAkuYCiHQ7aFMW7fvdyQm
LIXdwnfC1KisRE9R0DqvZM2WAhgAhHnC3U2XTLC1gzKuX4+ssqFtFLt/6IygW/Cu
7r1wa2pmCqYh0dgxZNYyG1304WxJdMNEzH58ma68gLMMIuquHq1eM7ho1BwEakmh
YjCpiyBWli+2paI7YIwMhTz9eZUe0xnAKVbYS3t9GGijKHEUhE2vop1QCE4swbqB
FtyRhZK2/xo4ubGeYc/dot6qprBu0AcAK65SiXEgQ8wwEsftRq1g3P4uTeCU5VlD
Byoa+OgfuVsc2l7dHmkTrnThWtvFmx25VMb4vi5XpSU8q1B/mlgjBSiuA8Up5itf
jDKxbJ8KmDT4RV18qFVYWJoiO94PJKv3Rfhzg0JERJmUMCmbuMEq0z6DDBpzs4KN
/2eLjHZ4Y2K3/WqENliATw25hvcPhh5Dl7Ld+sX/e1zlsvfDyaLEe/FRlAcsvDw3
e2tbr45I8x6gX4T7sKS2dz3MCxyOZ8mI5Ok6UKxfoWRhuvTN0zqx71g154+q8lDw
CKOd3vgCpHL2DHF8nJU/0VnB0pzpRGkfArTL01lhAaAQ7Vc/oQR8UThmKr3UOm7X
7kw9YIA9cHC+rE5e8LZ8wpGKlrg2KKz6ks//IPPv6JaFQoX/k8FNym1uPBBIRLJ4
XD2F5kS7oNlnp3fbHJd/MuZh4+2cZV/izYQnFJTEgwgvICsRWTUegTwEfu7yilKX
eCyLfXdzfY7BRzWXVIuGkPyar9zqRBKiNPq5lLdbygTsxuXmyD0S8BH1wgfhOTbf
GvvQRSnzBK639UZnbu1rD0p98YFRzzHTcyLedD23q961yeEN+A7Pj+onJlq8CTRg
f5p817eJ30MiHqp26+hqlL6ummzEnZaKzgRgNryBR3wjyDQNwlqn3fOdJwCmDPK/
MGj+BwSW2qzpVyO2EB1xXFlzatxDTp/WpYZdNU8l5MyoW2xn+Dj+E7Fhm0HBPQWG
/jckWLmisQ1k8VQcLQeEeZ7cvmpoQO0r3nst+cpXxJWrxn0cUw2T4ZqpCt1mqPyM
mJE8OKOPGXnIHuvck9oaxCcRfl9pp6aGAVaJWrqOMcI8KdtRNtaTR/Ggv8j1jjGh
YSUpj0+O0nmuJFdb+s01CjnXZd+QZlxDTDiT4kCMr28eAZU0WfLPP0bjKD6KgVaW
HzP+TkPJ8/Ag1jQLtt3yxk7OO+hQwsgO7wzhQNfzZ3yA2fk052f/L+uehekKma1z
7+rPGpEb+gCUiFX3tQxqN5v9ycgGfTsnHBghiFYm62t9w97NBv95AJNko++hgd24
Udv8T8KwsFBYCZKfvfVc3cruohgnxG+Tj8WVnYOliRbQKa0ABxxtF0N/M6+BNe8b
qsgVq/36L5bcSpUpoLy8AEwk4vHIAdhBpnFTleedM9AN+FElGaTJO12YlYrhb7oV
ffpvPL0VwMSaRyTN6+IL28q9yV1hRFcPWBDFN/RhaV+MEMwmfN+UxR8L8dpvTxvO
t0VUEjsFhRHz5JmLfZRt8es7Fko+xOjTVQWSdoLyWBsyts4xbw80WSlpYLpcGY4c
hIi5ijR5s45jg1CFMWWjfRL1a0oascZR2KNeBLDFfjfu4EEx7i7ar7EMqMRy72Ld
8uzkOQNLHFZq6ez87LYbVhd5CVdafuf6bQNLKgkY5OA4IJzKxIK1d/woYsiKqTqd
AsnRI8xkCr0yNR2eos8QzMZ6+3dDmiYC5zLhfYZ5ky+q6/Kza7tVHagvUvEoQlvy
9cR8GBHlwtvWBrLEZOlIc0MnfmuMzbFj8UqPtgz6lzDuFNw5VBFmOaql02rLzeQA
mXKFAhkoknihCvQ+EPUCuHA76BM1KqMvKgLPR4oNGcl1hQf/91nbwjBIj6tZyLLp
V5cllCas2frHL76BSS0ywAHTWAC9CswYGMxzwQrC2ogHmzA+HvT2zM6WlEnsaNvd
wUi6t3tN51dCgkP6/Jp61pJh6mwB6PqObspmn8LvnWuzc/apXvXctygWkiofXCKb
nEGUKIks6LqTog0SQN/eu3xYKKzFUd3Kj1k1BXEHc/jBuZQnD5/0HoqvjAJ6OdDm
EmH1aQWxlpdwCB0vniuZV0VO+koQtosBCu435Zv1O/5gksPFpMFcwTq8Ivr6esAX
S++sKzG2s7Vankkg9zUGAVj/ke+nLtVHvT8GrOUqQcB2SwbfOphlViEBl0g3rQW+
rR65TgKVGgIDQmnvi+0xRZWO9Mwd6TBUQgqtgVJ58BsNF9zbsjH6o1JPLs9ZlSBd
IvV1iMS/CQsz9xAzXQouKO0dv5xS8atmejcINjrftk5TSLcsUtURKcGPXCfIQFer
vsTfzZJT4zaD5ECHNbGUoA8xNK2wKVUzKbEiTKnjfJ3HsbperVeBihD9TGVrxcol
bI22v8relRS7VocVBxEk+oJMfiEruS7sg1tjqYB/mFpmDqDdcGbP7pLnDfhdYXND
UixKfO1+wsrBPXDp86ka+6SQa32NNT3R7C+hiO8pueXu1HnWoDtuyKYvEmdgGCXQ
tp+ZuFEI4o1vxGH/LLC9jf+BX3ZdHrEUJDG4jlh20lZSmcxSH2zzowt3r0X0ifqy
BvPWXt45VL+PWsaWwxeBOryTOQ+6zT2XdpyXOTlbCJ6ULd82jEYfoC5DMySox16W
N1qBdWemmsFFIzkvNPqhjAt7ZfbjuVqFhAPApL2HXBO/m0we0Mvgn6jFPI9pJBzf
Cv+vTvSTGiB1HehFYSkrWMHjtkbWHMAmXNBBIRwSsa0Jd/b2hwfbNkwy4up8eQ1b
zVyEE/JHXfRvBGX6vKBNYaq75pgXeMoWdf4YjYVUTN35u/fCaev+yc2YnTIP5PRm
+pK07htHNM64TuedqNpHVrA/ldbOfHntWQ2IY7tdE/q9DlMZFNnrMkOdhnq8QIVe
aygtoZmhH9udqZKc7cJpVLsQdd3JiOgiRylqDQTZkCAQiogt2R+/Un3c6bqxo10v
zUwnMs4oSBFVYRQqboNF0pBdABAEKikONuMAF8wbZ2e/8hE+qRROVxJVwYT7iT1C
vfxSvKyHxGmEkdcx2Wd3v9XXatc86n9FtjqQrg5bvkJ1jOY8NVsCh2AE1pydFpWk
W1lAU+h4mby936Dm9j8/3OamBI2lHhP/f/4cCSoAFfc1tSL8Wuvwj9Sfut7eFUqE
6mFVDjqhrDa6csezp5jt2TxsDhD+VGqIAS0joS/EUrLfUSWBX9PyqWdVti9Op2jK
o/q62RMMiHl3NBIyTtu2s8dNL96Qty+iCLEccly85p5sPTPA3rt/9HwguZggJVgY
YTzQfMU9USn8J3HnuNEMWRIhi0UY/Tq3nFOLQnucs4xnXNf3e/4dpBD+0pcrFmvO
gHvkwVZWcnbRcKyu9G+4g1xU90NMi1q/n0XXHLYLONisehjvoXxdUGXQIZ5xyc07
yVc7TU+pzH1xf67iaus+80wXMOLnzEJoSyfgP+1HSZeAIA9C4nfaTFjhXG/RrzXI
1cYbjCKI3m+zKmrPYDAQwDQnOz5Yi6zlgqOF3157GxL1C7LpGEV+nvrjqoLnA0t7
ceOjIi0Gl5gAVOz8c2eMBJaA9JSVFKxMKLeamW0XX+WuER1kfXZS/PPD8z531KHH
FrBFuhsbymN0an7qzPJmfK8g3yzJ1CAl287fXsZPF5sqTv6CyS9Nccayembu31c3
TJ7/vVSFVh7vbjtl6OtU0TtP84opCOpmC4uB0Uzi8syJBKnfxJSakSlCHbCkpZSB
ptGFwY8n3YRizSdpQ12So8aQv1Tmo3wzLHOFUCTScfLkF97m6ATU97Xkp8SFNYEg
0J8cqN2dEIiSDXQGw4wRQZT6bAQ8Yqb4PVTMj/WuZ7THU9gU8JXmaFD+ixKxhVIn
sCdOxV+jjVmgBlq4iSkOQRMea6oEpXHBvJ+dUu4wRUZqOcdU3QyKIycAuE6/3teD
5hsDmvupcPtqRxZ+9a/WIjh5WXSqSFXOJy591Anzyoc6tqQ7kroBcoRhiN9Y7WjX
WQDSYZTVuGfElvxGgLn8XSfopjM7bjkykx3qHpwwYBmY/MZaHdUtl1v1KmnGNKpC
x70sXcBTp3mdsCWhmsILqfILdJ6wFCH/0vvMqAQOG7NoGkv1v8OwKFU69LG8fG44
tyz4toLyBvJkHiZOH+gDhkQ5ppAPUjZpeGdlOxrl3F/bSy+GR97UlX/4+Yci0N3N
z3UfWFy9+kylnCu52Bq8tJWoG3nQD8AK/wLix9Tw2PBC4mf58IFeUT9/9Bjx663/
WKGLFKJjo4XjaH4i0OMRWx5rF8tRIRoRHmIQma36yq0+YsShhi4S7rk7Dob+gZky
UxI+DWmGOid0qUPaVDCC2paLFC0aD00HSfTF32wBS/lYpF0kwRKPtRxrF9v4U/DS
rEtMPMXS3zaTyNsGJrTWTUF+qASYxE4tHpZbaMCcQNPDjDhCXf2uWBn419OIyhJd
R+15DaIIjPnfYXValQ00kXRqwG8FPWrEa68jcQP1nDoZwSuYP95J/5ONm7Wlk2a1
vRtBRn3yDtgvAKkXyXOvu5CWT8x4BEZq36IN6GRi0j0hTXv06QgqZC9Ur3MUFCDi
hUeaWrjGfrfJhxjjXUmtdg5KW25Oh+HONnYCcRiPuwsHZZmMLYJD/S18a67DMjer
FRI6JJckNaTWBHu8qZHOkDTPuQNvJt6H/fvvvFkHqpVYYkEqooefM5MQNVfewuwe
AiRQiW5TlD18V4LEQ9tRVcva/lnqcNj3GmKoNhfb4Wmuznt5iyQV2D8nACyzV3CC
BjjKAJRIYUlUYtsIFVBoqWqRbwhABUP+J8fs9sg8DJIUERv7tZG3ZecfhkaMpy7t
aRJE0XWh+ha4j/F4eAOLRbs3+WIBuA8oVq9khN2pgp9L5RxefmnQ8hNs8YAKAhVf
kMDrcQ8XI16N1ByMXGCdhj5jququ3m+OUtNgGwT05gUHyYm/DG7DCem25O1HfxMQ
T6rRYVhv4tuxsE44eU0YIFZWA3LYvYokKgqp/hsPXP46NyVAfSwM+bJdIbWgYpHV
5qYHC3D8LCutYITD/SBtDULBQLLeZbdN4Rq9EdIIk94MkZ9TjRV/Xi60oPEWbjQE
rtifS5m18a80bM8e6hYejP+ctlp+PH/u3eNkQp9tNF9NYIO+xgoVlN00/Ch1/Eew
k7+T7yqOxFpEncBmGcf2LwL1GW50zVi1bEFeiwbbnJMq4DuTF9K6YJ22+QAdp5lq
Mw8Gu1gQmnT6dQdSiZcD1EnsEJfMCmY4QVuciDjSTrIf1P6SMLWbKC0XnABPwmKz
4pX71uDecz1Ex7FwKuzMkaZu9VGm5L9IdydQ9QpBgdb49p+9YqDGsjf/dUnyGN5G
PSYHML2rrM7dFCGA0Nrqn1A1ywnHTh02QQIo3aRj19CwdfTmTeD7m1BtvpPiOeV1
oa1YpDhyl8N7bsqACn9WdimTjj1JRKN+LJ+V6NhJVh8NQVvsShfc0VEPyPSsKq5q
yCnzZxOiDi2Mb5tp5jQg4ErlKpJpYSe3wjoMNLUgojEHUYj2xSp2Ou3H6Xuxw6SL
tR2Wd6JrWetJMnpJvev9R9ZldceMBA2JxwQOjXGA2IgD7z4HYXyf8SzqfPvStnLJ
Y+VeLME9xfqBUOOVGXy2CpKuSAiBheBZUE2vumUk82Z5ph+URtfYqyzKcribtulv
ZWcBo3HB01CW57LBRMHK3oJH0JqdNpAlUqmpV914FmElJUkQIbrR0ffe2dH1thm4
UQk0RvwOrsy4GqM40InI0xvGn6RtW1hggZl9DMzaUeRCFnSxraJtKp+7oyoP3Pln
zqmLAwjXUEIcTjPefMiePCa1yRCssYrVsElbxKaPCJsis4m3Bg0nGOk8tQnGDD8n
72qaZAeiOU46PLFnsXWIqDMETZYfWFodMlfTnkUaFc52/oNEaqQjMGfZtjsTTQbr
IiYfaPGi3WAiLH9gWxKysgkjisj0iFpGR80hVrUArDML5nFBCdRJX2mNUACtGAg6
3/n37IeuM/vkZUvqaQCGp8YYfw/gajR6Qij1+frBbEMxcZCZ+oWwYPKcX3KD2Miv
tdk5uPvcLUkDq8HHq0uOJ8H41f7G0qGsxfrMX5oQ8R3CHPP6FGIwvygHrnJN0+kt
TUOP+c6oqiSFs8M1TDKdfd+oHtrnYEXF/2DEsDLCTAHgOHpKtJFiO4q2s8bLJGZH
YvSxlTzSqUFu1rsR2q33cFqhaMDqO2JvhTYXYCLK1oyAINde5CRBz1w2e30x4RML
a418/By1+di2FIKTCcVl63NYtLn+rY+gaRi9V/Q4fcKJ161UncxT8+QiqN5ElNNy
wxnVFTVADU7i51g5kHUNAmzr6PaZ/Sl5No7NWbbbOoUvACaZPL3Xq/KB7pTBnGmz
Y5xVkHS9OcVqpAORWHvw8I08F5ZqrxOgvXX9rb2cKkDMA1iCVagYlYpm8CAsmMrL
taR9TsPWdrq8+D+qqYflTCR7vAN20tGxp5XUXe6SinCSXGSrLGlL08/rIylm9PWo
/frVSXakuI7a98wxiFnXnZCKtOsWMcUHFNDWXuXn9GDQnDIDkrj/QLKva7UOgRKA
UNDMEuaE9sGMD5OreKKzirYV9hQAHZnurKr8D6eQz4eBSVv8oQCYdJ740psd50Tg
B9jzkQczWyYEEzKrs1sf0VhtTLi6uY2GgHzuZMtKx84cCoRCT1P5K4oEPlc3mBVO
GFLujbkeT9kOoEqEGueC2q25xvAwJ7RWt40p0cL5RCRP8ViiMEQnMnWbUMXjdm3n
NT6+HN4jAgcJbFe5kUFazrW5fxJO5A4ecO1gXk8NcV//jWJbrMQHssk0vrENJW6l
R4gfYmN7T3kRtwv6EsuABtbXM5XbeZ+g0vfQbauFERK8Tv5iJRB9++MG6lBoJ7hn
6kMhDwMqmqh6Eb4Cfr8oYNUeky5ZQ8ieRLfBwna8suOYgP787hoFFnNA2ms/LQ4w
zz0sopS7eBv+F76dm5yfKNq2sjDnu1bB8Y9zjYx+/FAOw/CSM0kVX8Gx7Ra+ABJl
cp0CGugZ94mFzy0WHiFyLlfnaQ2mJFXSVYM4EUxMz2ZV1peSai+Z/+A3dR26NBLD
URTfLNUZ+5iJdhVVZsmZnscJM45kghjO0gYamQ2HefEK2xuJzRhyXc+Z7bMRk17b
25xkUvqkAmN4VGfVwXRT2KRU0Y8B3xYeSFjZQ5l2hphTF9/PIN2jGMQskeUT475d
CkjaGlGObyVAxtpO540GvKuEYlwMva7ErqQEnziCtFYzoCm+C56Rv6wxybKcgdVS
KYCaWPiCjobinBbmLoSi2UbYHIt97lNaIWkbvJeBpunFT8oBrE1qzDDh0p54ZvOt
8NETHf41OB2EyLPjHywhFuLm6VpoTe/9W0vKCik1Qy0kPJASaZu1IAMYDq1bo5Q8
ArozWGQ8Ix201mjt7E14OoZtJG6zth8s7TZXYl/JuukxKkaOxdhOTxgTXNXHx8kl
F67cbSYz/1NHQEjsByCANVbB6QC1pFMIm4+Bj/IhAPQKDBHcrm/fg2Ye/AQ526hi
kFq95sKYTc3VaC1rVD0dWBaRuheIXEp5zw3IC995GRrqDemItvDsiTWVORbHAvOn
+jYsIkKYURrbFZ/8ox5oGiv7xinucgmeNcuOf0G1SMlDJ3f1Hem4TX9dQodEDGcd
+ata19SjsdjXA+tBpWZnCTh4qn8etwoe4/IDy/0skaDpxTGUuOKejQTJRKXjXMKk
FJJ35YtbBzFdvEmQpcIYpcdjDALNyrZg26AwnMByi61V2G5bh2PR5ivp0FqhkwtW
DeMwqySVMNY/qQjfUmsR9EY09VUhi8ra0rMtDQVB4pc5GTjm4BcuiQB7jsRePI4F
8QG6tq4PFG+RJzW9goEMf5fbz6mZ7oE43+X+N75D8uVgtuBM+tr6cet2OGd+o26N
A46hX9AExUKgbmUg7XsuI97ShFw+KPuzdp9RlBeVitTHrQLyOTDdaBk/uFT3pkQH
Jj8170YSMn9F3tO5bOyzebLqdbk+T0oz3zzMdOsiUUrsQdM0SW5In1ZHCCF7y432
OLiWIJnEL5/6xU8e6ZQMskhOodOY+sZknyJVJjP4sFLj3jW46+sep5wI7U8aJUiR
MnNRyRun+AegR1SJUTRG6dlDvLSaPJBi2v3XrpLAw6MTDtddXvpVssYswlZ7DsDx
N/v8mG90cugOU0lYOAZMPoqX8PlPGROUU+59iIzttVDuKqpapKW/j6oreQOrFAfa
4lWF2eqHKWSwLx2AV5ygcEREy6eqRmXWms/JAHIOaBPc2viI57HKAMIBmLBiLYDi
z6tU/7aEpd/VRmlAO3XU3CYnN5ibZnhfiNzcXg4QjUd4XF8ZnPTU2g+R2kYp3bsF
NhA44b0KliK8+LDsuMzMJggsoMK44ddtiaZvyigJ7aLJN7ktnZCZLggGCYT4z1/P
zXJuCXVhz1HW+7QmI30Hwfvia4L9xg31cmCtuIUb1d+t8BYvPimdjEH99iuQP2YZ
kC6y7CPtUZYkordpGRxdRgAK+aarC1s3q675Q6nOQJEuGX7LNpIqHGa+scHJ28gD
lYU9YoB7gpdaMQTGdVpxvyr7EEObrtLitre5+WR4OSdt9U1d1HMSyriiqCLZmUai
8ZbMVx+VFwKvGyzrGiW/fskDY80Rsmd8/c/8JPX6W1Zed1cNNluXyFbtVS5GdiwF
gVhFU6SW7aTADPALsyfHGcXVxeUUpDZH2rQmFSyrfLR/oJV7CkEeRbyBhmz4GlAk
Fpk7MStCN01AuJZ+zEd0GVwg3fzmmEZFnsfvv5zADFhNzoK5Gkm4XmLjAYcKOyKK
nwen0nJQzQ/kg/kZoQ/REo2r/KrRfWt4MQxScxOJU/mbDsjwfdbt0YBAP/Hch5CU
ZRiA81r35bg1NoJHcV+4VE5Mmvcox8mT4x+cWE8nbZ0Vc7kYdbPNRaBCBjiliLKt
I4iCv8ic+uUQZ4FlAJv9m7+6nDVtN5mQ/mcIWsHwGVOMz2I2fdUpCF5Czob02H0t
ojohOGlxWlT5wckailMfJxyBZXP9lzeBF6G1zdEd0XQpTwoBzzk00dajQZWpm5XJ
2Lt2y2YdKIXpOab04qhL7ENTTQeD1mXrZmuvAwCiLxO3YulbblJfk++9ViFALd2B
JrCc0RoexTZnBHMmKgmjPPKT8n3SL5G2ZOn8zmHHQuNVIG0rjuiemcWVZXEJSTma
onkx/ojDJbZAIQY2tTowRcbVRCgSG9h40PkS/4XHtaRT5HHlKNQjvNygcCQaNHRz
kx4gb9gIJS1YCbYIjtYFcw+v/laNAy93PmJlXExJ/+KlZYKA+VmJAvjHM8NSHafl
CDDC6YswnO/HZCReKOFDKYdQRozXSAtBRh3GkTh5+iG38PvWO/tc03l8d+LjfTP3
mkhHV45bc4L+jGKeEcAqE+Rt+7m9Y1AhpKIwukUx6esViGpcOHSoF71OGXWPr/50
6ILT/sRN1vq0oHNdOsi6ccppX0Ki6A0016lazzycp5T+3SHFddW6+QAxDH3CctYr
TUflL7cqSBRS3LNEWGjBctlz2tifaqaN1H9I8gtl1fv6aYaBhjo5oiFXPQUHfHWR
p621GfMGOgHzN7fP2/rumqo+dgbTt0iirJg0nC+79gsod1Iu5h23sHZUzIioT87p
mMm/rfdX7X5BKBqihbUJ/6L3UxTm/68zfuGvGM7gKyS7WKcrzZjV7admA5Yswaee
vLCG1IAjZBlxbi7984oP19E/4+0Plaq+lTS0YMyRTC54sPIH1PT7lTeHiAkzAU7L
9nHujzid8Bg8aZghEI2Lww3sAjITvgBgJG6WZM6DzBkFcbE4fZ7kqOSRGW9H2C0L
pL6NHr6AqzAYa/OgszF8mZfLqeppEauASNPEx0roqNHkUxTFSSQQzi9uxxa0P3HU
5yoM3b4r2h9XPfmwuRQkCIRsBF7QkYiqPKWOs75QYL3DVjMAycpY77sY6MQu3J5L
N8/KaBU2QMousgsL8RPFn+vVicTVkoHWLCEXaYhv1m9fwH+Nfk4+pPJZC4+lUrbP
SDy7kN/pj0DHxjnA6ZS1Lo3umBAl/vWqzY+6bCHzTr/w+OvscVz8UV+RWHIWhHFv
ARBcJ9DUy0iwDiTeHktwBnFN1f3YFvORk7tWDIgSZP7I27BqVCC8GtyIBIO740LN
fqI4wZn1lIgdolBUs1DA2ISgXdRHM/rZbx7I+8Zv0DxWLSYMW4tuLi/9LFPuWHwM
HkwrQ5gb1N4Mq3XBj4z7FB1/qKmKR35y4MPVwVoc1yYx1ijJBBNKr0mOFXXZiL7z
k/nuGeOBtkih4WgCR5gUGTowsvgerVswGy7XtGJmI4xBN1uxKvCZhc/SL6pPiYNW
dbZ8ukvxQvtLNGASJhw6QjzA24T+JlshN1YnSqf4vivMb4KW9uSMzyIPGcdGQAs7
kitq9V9jk+azxqjgGuAnzR6gY5R3QUVMTWXhMUnNO9zLDcxM6RJ754SmaqDH8vPp
DQEl+THrGnJK3PlckwCXBn0QgdVpxij89ZpSgBw7xEI52FXJX7QYWMh6PY3+i/fr
T4y6plK6rtyRHOD31X3LRpcjAaqZZRG+6UYpHjY0lPdVjeaLenfcd4EJH0n31uZh
O2KQICwXTEb5j9MCRSpJJoDNPxBsj9QNUfD0omqg4CdabSn4OozK36lz/4ecAfU8
dltIr7h1/MutnadPzkUHwN17uG/8IsamijMJv+FcUBB2TuU7ZxAxuKJQWCf4WAL/
P9BoXoSMRqdNwsu/LvqWhpdFk2oJ61quVDt7jtN6yIuPJcZFJR6jg19Ul9ENMLVb
6tYabgC7jYrxMeDX9P4VcU/mATE3Df/AuS8WBXoZhhJnzi+FxUllNGoIO0ikPu2d
1/FFU2cR8GU3UI2ZN2+0YQxNWPMvq8/g8HK0tVYlmuCfmroEbseLXPMGg8jd6rwU
qe0ugGYpKj0zYsZVzfqDMNj4PHD30AbzCUhyIMiQDljEgz6ymsrtI9Na8M3ynGqH
pi6QUYeoYRgldszjnSyYIxJAeD5wm1iafVHwSrgshdZOQkj6hrnIim4Sdviz/lK9
l/qii2OGRt3Cwu1vZLtI0HgtfQYzVLYN0hObuAiIk2a7Ax235l7UnHes51ThMxYn
FotXvCUWF+loIsvoSzk5aGZgUoH8uiY8N69DeBs6iZxXWuZzwksELSNQDNTpbqZU
uBKa3p3EQGuRRvcO9siLzwPWuRJwY+wmcXgW3jsBhhxGylkq9Uikv0RZ+HdLYY1i
Y6PeetZ4fOPCUgcualna2QjWiKISf3R4MM76SDlkuA+Bf3ojHnCkeu9eLoJLbk60
PMXBq+FekoLW3P3/fp/o2Ng6bOLMKAQNWHaslEcQmo4tfmTHlAqPUGeSijDRdALH
1D1P0gksPbwROTHjKsiLcFDXPKlvqzNAU0KkmK458xpcZPXiEoj3V+dsDtqpsqna
XARKKaODNWyQiWjtX8tLfW0EOJgCklPfLzYoHPKDUuVNGu6isCWhOorEI9XqK8NX
Enif+Aq7wxWgV5Pr9c9NdU7mtMSttJyvyrBYUvdqWwiAp0BxElizkfcWKmWdLlKo
NqzIzpTfNaiXoetgvXVZM9z7/ML32WJ5lp4NcAc1sYWdkkIlEGTbAx5aZYwn3bBk
6uw1XqFLNCey53ufOhJhYRELllg+op3JobhSt//r/Cb9RMJvckBovYQfswlT++kY
MvVYkWcwhMeiphUEuNG94oX7vRprbjM5ons/1J5TkKdKJAKsrwC4juJud6sIOy7O
I2GGwbJOQAgC4ykJtp/ytWvUFK2x9vKtWr9ZoMtg+3YrBGswH+qwXr65BYVo0bB0
NudzVkH7mjZpO9whN9Sxayw/q5wpYhe7WliuUIxgIoQFtkzZ6hiKXZdAXRlOBJVK
WL1dUgszR+SFUf1tifDDbxP0SXyiy32DVuFLlL4xHbEezTH6F/hL+QdATnNiYUys
I1CLQ5FDJSIH7PXnGJnv5wzJObzNJ9Hk5lb3cmcAy6uCtdXfUYuasWcAkAWm09/j
XM/XR2A4VmrUEhs6j4XdpAVh9fqBGQtyjzKKr9RBdmoOLKNCd7sAjmN/mfqlc3wO
g3wshI6GYFxt6o1hf+FFp5pZkSVzNBMj/bq05L8vcn75qK3/SCsa/w4iaolQNZSa
1TxSscA/e3b8tr5hkcB6lqMXYEYd8SgTlPP4atl92wPHYD2w04zS1Q2zsbcB9RFZ
izWw76CN2SQGKSqJPS48ANk3qnOz+Wtb2hoN7cXXgZmIM9kNoyQ0+Pz0Wi28ctLv
Q2f5rkw1VhTq9eqwo+kAyYeiPBGR/n4KQQjSKdUFQ8lphAYDue922G2U3ZNzvzLX
9Xfd4ynNaAZgB5fTq9ulUIoZCq8INAP+cztl2sQO9q/pduJVrnYcSaWSywL67qC3
HeEuAo+fm2TDqeO4B/+fQlafeAkphOXC3G/kON6Yj10O03itNmDs0GuGkYvvN9ik
ARqvHlEbjgdpAiwv2Fcxd0YHRsezoTASVyWFpI3ylfFSFRRz6ppl18Kw7FPnerI/
dX2oaM/LYu9Q7zSo22iWG1aL2ZtH2ZK7D/ww5sFTJIEMEbesRQFnpzih3j61XiHI
ZfrmmVsfoZWKXHlD2Y9ocOFp8jM3kMvY0rQ6OYgj7hZoRiBc7dZf3mUlTX/Oy3M4
llZ5Ro/kn1Aa0dz3XuOaM/dRsoXKKk4kpPCwFgI7FKC9urQpFFyxKiO63Q07M/sm
cINwI4Lbu2e3lNKOoZqLL4aHhO6vt9kIl/X2fN/EhWu1pZVy1bLWWG0U3NpDlIT5
KK3J/NuOf3K0fAd1ZKBHVoJ2QdFuvPX/0FdVm5r3a+Iyx7dORf0y+HhrPJ+U76gC
IT0oasC9ta0h89LeHLuRTmZqL+Z8cm+vrlpTwAw1VpzJbOkY5uUeM9bVfy6OFM81
1RR/voVX0G7ZtHXuB2YcmpoUUqNG6N7Y9ZUyZJZJLy/RQHZUSOuVEjRfCZEzzc1x
mF67Vy9ggZYDIK/3uti6Gnt0G6TgUQLTy10t0Zk47PseCDfP19IUi/1GubWlfjtU
ppO6OQI1kDWknaPbBsdCzjrMf4vbOHUeQzOmMFpEAzTFZ0PgogdRKMZ7/WoE8DbN
xjxYUCc9ocVNLZJjShR3rYjnSiNdMTgdSP1X0kBqAZQzfpJxbSosGflV4y8Fz0/A
bp3IPH5zSYTdoDrfv2mDHt5W9pQqEIeK8aVzH0dfB7XtfYA64QapBWiof4w/D6w4
2invQiaiSKy75iDzjfq1svaqWDOfZhzl5ubBbe/suMIcH2XzTCwTNWmoJR1x3rQE
3x5OB73cShFEKO9Ej8nhEni20OLJLq4TwJomNQQbFEO6XS8U4DUbXeiefHnirnJS
HkvBqqFYFY96DgS0wtS+0LhUmqwLt0ju+nGB+W+dd/IPRTmCMTpYTq4hKGGXRKgo
3x3Yas90NOgyNbb/BM9dBA0gtMSmI8ZUBADm+mSmQYQbF1CuIKnY9aYSE7V8GsQt
d7BHjzwYMoQ5soWVZpdPuzC9IhK9HGERuBaTRlNSMxSginM18RF0U1qD2GZFC8fN
viycmL7Gq5aPqZJQSGeq2m92N9w+m2EDPWpskbI8sE9MZXkv+xgh19LjXZe5WrpR
UtTgEolAyfXcoWEQBoTV8QRFNtTiGpRhnDHagquACP41ed73cQbFV2yWM0ZONu+g
6356RV0E4uFHc9cMFRsV22NjqDFle+YIE+naLzQOfIoohuyIbtjtU8GoMb8z7Xje
KL1hc/ovcYIO+/cp7cPIp6vVefNCae2jfoVw9oJhnMUoSSYUekoJFFlgIHMl2CVI
AAcAGLood8JFrePX2Woeelklw5n1XBB8FyvisSFBNUSnzwFOYszJEJbTO8fJew8h
NLks02Ax8lbXp5wZUOkh9pMFy3JQBjlpN1OB2LrI7Fv+uFFvKPH8DH5mTDB1ovRx
5VX+7ZzvhMbH5LX1s/rqr6fv77lIBFpphxRZg81uqjc4M8+4urxea8ClMn5PS7cU
/dFqJuD3U9Rn9vHGqI8VmQZR1U+HawZsjBRZZ8UV6XGLte9PM90tIPRap6IXpKdH
GDZ1fSjXM8KrojoVgVtH6pVCg3bQhbNegrEU/i6nPR6B4CiV4PHPzfdefdlMbr+t
l2TJEn9eZiY6DcjcfI16RIdvHWSoAq7OJZhuTzdsaImSziAbc/2N+gUGgWemN5se
mynz49Ah39S861muimFP9mKgEDDr1eeKY2vDvUCV4majRch0/7EKESDr/fvsrGAI
Ikv2NfzYOcXOn5Sl5ffwZvdmeoE1C/lwrynio9sT8Q1aI0DxLThd+qbLzkv5gfUc
Ij6uimnU4C/lDOJbwGmuN7uA0bpEVuz4OlOugqOZmGxzycz9j0g8o4d4mwMQyT7e
AiWvx7NaIneaOCT73P/4Z6k9r3VxuSXzvgMnRWuNMUsv9+CtfgScmkN8uT5dwkPQ
WJQwFQKn8eAxngM20S0sF8edLUvgs+PlcBZZpUam+kIDD+nq7b8aRnJ3dbUOYTGa
bcVz+Mt3RwG+n7VEMiqOvfTcgpniz3hNbAQyV4m5ZLSnfI1QHXVLTJ0cr6tBHhUo
cF6rd4a4gltAXVBTbVSl4n9QcoZbNxTo1QPBI3ho056BZLXA810U4AopX8v3ZuuO
yRmEfLGZ+e4YVBS2oyK9PBtPvQ5+aD5XwGdtvfdz5MPb0crI2RgkCM3mPBuY7IPX
mmr4Nll7bt5Le684/jKVeK21TM+h8l/B9agW3gUMojbSJNSM6qyfzBrxol+2bVw1
haeamHOmGu7OWzVJDymttP8uVXr2F6sB2jj6qG9Y+CDLc+SpyTOCKsP9lalF7ruS
aBKtoKiMqF+MHAcNyfSEXu/vKyXw7cHOsTXtxgHKkqgttogXjTCZodEMcPl/xe/s
ZE5q37086MsLl6aNd67WoB0N9VhVPoatt/ZdGJGKLMIQezww/KQS/gIr9uB7EIjC
23vRyISCi6KY/7L0CVpe7R/paugM+aWCuKTpZJzVEp9kfIDNavQiTq2O5lzyBFdX
y3AFIeBgyriw/bcW3rerXfxzhvPpFbxn8vTWSyoeuE/BvMxx9HPDX+AYjNADZa+r
nQkOw9xV2mVcHDmVqxZf7SY9cHm7uh3UYRgEF+RkdPjrTyYD8v7wjWlRFGt4LdRE
UTIM8NIBYoD5k2CrBnK7BEd5FKnFh3enkE8dTiCDSxHnuXOZokwm+xd63teppaeR
hgzdd+6430kSIE5c2jl8jj4ixkj2bKwvWz6EAH0GZmjhzMjCPU8aNmvDgGuwJsg5
nckv6nE2fEkefIICZ7ELgq7kHxEIFAmH7Qwt14ZqCXTkUhHtPMaSG/66UqOkBQEW
h4OnN+dtp+p5wt3dFYdHKfescOef0KZoWA5VbaYuZMmpVcgprGqYv2LPH9JtnHqr
XE3TtYvpaDhI/UkI8yMHnLV08qrIRolxm4ZdlpCf1DOtko+a3RrTpCcyEh2zH5g/
jmg3gM1q6aKpceCzetnyo36s9CYdAM/0tAO4xYThEmgWztbPd3u8JIwszefkLPUT
ThSSgc1DgjGz+IclgJSDF7FgHj19HICAMthej2hB1qnVF/SKwV3NNYKUbtXbIYr9
KyPUh1S5xKQxcVUMh32VqXkllKANK2qWA7oN4533MZVvc9DlcJ+IUM/kNwzxoDp3
dnT2sYwJ4eNUeFL7dR2Ypa6Nm/xUWc6hBMjzXYYNTsXKkAPIwlsQ2mBdWN1gUwPo
ZxZxichUYser8FNDAat8yTHae3Okmqp/w2jZ1vRACt11p2sEa2ILN3qSsOQ62nFC
ZY6XtSpw13MUDtYQLG1q7l/BvxQWlP/JyH02vU2xZFnIwrlVbbLQWkxW/TqKHhww
r+73cFLKg2WRmKSbavHDhWbBBFWRyjBiSRPYHXgw8HAmTMOQsi6/z/CneiXWAjhk
ga6GgmfflepzNtu/DRBIVtn6mj47U8HINr1WQ5g7wGFKtAtKp85GwRrX4L9y0S7Z
lp+5Oa185CZnWBv2G7PLgn6MnwblsBeLTONCR7ThNzWRVqh8GNd2yQTC36JRgD5f
psXhuWommn5nXlJfk2a46Frlk6959OTn03JdKVV4z1aLXjmoEoTB566Fc8cFRWxT
vt3HpuHmx+5+puKGHcT7HepslAr6tV8bGvnbAhO/yfp6DGr/JZga58uBorcnW0CH
zIhqZbXJ3a++MlK2ggEAimE9hOZCvW+0YMBefIZWQB72lQ8DW0jdAYCLw8BhKG/z
SH+/MJv87ZDAoiReGP3PIOAhW3shmQ+NyBOG3c16pq0W9JPa1LpsdyYEwWpmZUuF
M2exaXnOe99Da6wc+YQId8aNpElRlYxVsYYj5chhjTvce8y6WyVbvZKEJwy0k2qA
X13CY/5b2O4JmecMDmyGGbTpnOEkOxsYl5q8tDOX9iIZztjCrqSl1mfwKYDE64E/
JkSBxiiBG3b3RDi49jWI1U4mczxqFzF3bYq02SJYLBVvtDdmZU3ybsQhQ561QiZU
7FHhicXiGqcPypkWoV+D2t2PK5WxsrqpjNeWah9XbybGXE0yFfwFv6JCzGyDHOkN
KJ3cK76+CttSKLyjUcfM+vB8axhNykgO0PGL7ffFzvUG9vGa4SdsQgQQxc5Iyq9w
1y2FDpRlXI5rpPc9rlFYvPAo4JFxdG3lReZhgifW5NiOAxbe7DkqiZKA19K6AaSL
2EX7fxtILd4WssglAJz3BpDQNVICEQL1EuzbcIgzmPNYPkVrTbAKRAsPRxpu65h5
FjaRmzYL5fECZ5pVbZANWF1CvRId6mPp90FunjTwA/1ap16bMZdwWddbtIYuGU69
p5cGhngxWdFuR16r/cEfRbQyoYjz5SHY3Tdw79s7KmGI8OgoNtrvr1cJO5OvMhhJ
ZDO9wsT68fNfoyQmrT6uZqJYtFtwMFPR4FnZ3jb/4wh5D64DyfNFUZpScvuYC5gk
JLi4oBdvluZuk1qXWhZO5oqTnhGGbj2SXUvZptZp2oq8RNSWr2M/B1qTOIHM1+Z1
WOziDC00wSfbmQZ8eUE/E/02ZnHuyZEUvU07dtiZbH1Z9VkFrLfrK5EJ62jDr281
RbPZGke7sD40Xu+7GTZm+sQ9xnwgwl+IIll0EJMygoGnArsbqumL2CQBUAcJkIY9
vwymCxADr1eGk2lZ0zVcCfldQzhxIZt5lcwr3layGawiyiouaIevNpADs1bQx8v9
ptvMmFERmHkSEMkvB5YGwz5GBCfQ7nI0jJK1kd+wlQww2esKmiRp/Wou9MbmVnXE
RfrXigjaB8UtjyG02Op7OLJPRzJzFfkMVgYXEi/5CxCTgNP+qSTtW11DqfLA4S/v
cH+CYE4LkwkBawWLOIGCmZTvVuahxpHPYQsbZepjfHriQuK9OuPG+vdUhhuS8goX
a9LAsl2AAlxO2LkLcj3f/Km+xbkVLGSLLdkbcCAMFWIFvRM0kuyHDhZn/VtKsAL+
6Q1THi/8umpRR8W1VFZLQ9RyaMlGzqtxxpAOkgJ8IOuD6QuPHKKGVbYaSgV36Hk2
tqhrKYlhr4luwKTYxBbrClrZPwrOpcmy/ddWZlhkXSgU6O24yUaVO5jYw1YzgLvw
V0klYTel29vO59vy7lGaonk0/pexTBAi0Qy0KjwDYYeqS4csV6QDYMbMpYJ0DRFA
r6P3QbpyfJRE8ZSbHSGE0PkYzI6ZGknguvSpqZE4CjPUUhul0zULTSf2i2ct31Ng
/4turjc56Yh1uUhtfISsBIhOL/icMEWxu7dKOlGb+fX8OGutOSkvdK23FWSkI2/z
whrY0pjkS0ZgJ+vU16ASg9W9EeuG7DZOEmMXCJbl+yfmj8irStpcsJ0aygJf+7oC
hyqb4UfpqcROYA/kh1kmfDFkDftoAa490BwrPWNyRfmgOSAqKHapzLJ/FIXuUaGW
TaS1wf2EUWdM+G5oozkume8ae484vhEpRyFWgi29ykIyFdxFxg3jS9iXMBMKWrDG
awHhSWC2YEYCnl44+JIgLjwDXsuSZ+rFv4o0Ia3OEJBA8rC72VZFl2bQVWri4X1h
ZVGvjVd9+mm7n6gRLc7ec7kDk9rMKyR8lnIrF3hnuDuqS05yggTPSp1/Rn/wmHUN
INmPxcP3UDY22NFuV1UEZNVHNVUYIUqdbr6H+7WeBF9eRXsXr1Hq1Llhng089joY
RBznOuIV2z12cp+DIPBj6kK+F+gwVT5Vh3c7f1Qmptzdhkq/D9N98oxqplWd01mA
9bWe/8Udz2KeF0+3vJu0QHDYo3Xo30bqO5GYp5Y3aHF7qZAkTAUSeGgj40ab++Mm
obF6jZLDNqqbnxKbcc5DroiTIBfC3MFfQSA5uFFSZAAcL9d08qLgtxfLxjp+D/m9
RfjS6HfDPOVEZ4msbD3CVFAo1zak/5SNObujvDoMW+kYtm8A4UVsqW/J6zgJeZx7
qcDehDj0Z4DUuvSTsbMik/f2F34F0MqG0JI0LacLYonWiMokxa9dJtcbpZAAw1F3
TviS4Ot0bSYPITfkq2Pe6IM6yZh7sy75zlup0Hau0nF4jdKB4XnUk7WizzGhw9fz
xiv5fYysANaoydbaTMtxtM6wGq8I/tC/CWexzXf1dzBbUEoYayi6HIODyZJAokW5
IXhMPo9eEkj/C5E5Dpdb8OwX6l7N9CANNPxS1dDypXoqUODoqtzI9iZWwYbbHFsi
E0RiaV/TMCQpKSlD3O4H/HCKP4bUyox25T/A+yH7NWvcx43apD5L3IM87sPMa0Ah
xZDgVqXbEqvna+ZBR1i6fq4WpxDwsWXiEMilp6goyRZrwPW3KnB5NOIuLEb8baqP
oRHLqbGjRM/6Z6ZbmCq2AETgm9QG7P+ZYveKWAcAArIrzvOjfEua++XcfMLzy0JD
4Mxa2l9VY9AV05KQf7xtSlVdFrSS6J8gMcEs5SEEgmB1UDpxaQ9G5TJ5P7ooBSeq
6UvSfChYFgQE9Fb3xEyYMX5ckR06BaJFdyC+zamTtBtPoUXrCPy5GQu5lM7STBcp
7qlfDlstedpGaVY9LVdJVbva9hlfrOjcA+QL+dq+tiufAInweiEk4Gmv5ywsLro8
3n14WblLBKOTcEb11PkyXg9J5KkK0cS/H9b6zihI3kYG24MWVaNy7XC2x2ZSvTze
7WU9C0yEsOM+2OZXzmHDABbIP2u4J9MBp+m+I0tRBW+VyTvCto2FLuFEuBnWwL7i
ln19/nkEhI8IXcn2VrP9k0FeU8AQMoIK4Ge0Bo42atEZqt5vJ3yJU1yHNWGC3Ew0
qRdnl+3/NEPie1K74rwyGzUuwdExCxqQH7C3Qf0MVsIpV+2q7fjdyBnrJKgvdmIp
U+XQO5VAyO8rgASyA4H3HzZoK40KckBy6KxUDmNIBclh+6VbZt9EZc3KFePos+H7
4uXs299XGcD+x9gbg/ymGyGxlR/fmA4+X/gKZHGhX1mP0byAl9rThlWeJMZsM51z
w/CIrbOOZjKdTDbG+ItbSJSEgX+EOGbOFRXjpRYD0PR6vQmRXkRUjIOXSCKPIePs
yXtFGo4K4pbA8wCNl18m17IBK33O7DCQ9HEssUPABtsEei6Pa9NQevTJqCmVehrj
BlAiNIUtDSDRb16Fic3t6SwwmxpidCghBiOenizaqLxtyn9Hc8JydD6pGTijcQYS
L6qu3JYayWjXb0tXUM9vbr1bLRxDuj4I+gf+45pLksGF5LN7ymzE6FGM46xIo6ch
3AcPnu+sZ7RWZM5ganXZPjRxvw04H63PAhuTqNgTUfAu+l2WWRB7aDNnOLZVKShO
zLm/0iW8EtZbqfg0hS/G1L8HbDWPVTMvF8WI+x05m/zasfGc6q+zFhV4atGDBjVs
2jSgJaH3DbOz/elhiWFNkasLqicdgRpOpuV44IZMNksLkKZXSb1tasQqBAswRHmO
07A842Q9v0A+JVWq8artXn876eOe+R77IW1I2atSKx3g4S8Zhthi6S5ycC/evOOq
x6jJjhAdSVW/QHyIEazuvi8QW5esZuz1b9MsbLN+eyWQsYc0F/WI/kai7h/G3BWK
T/dj7dHzni0kR76NgM99u60hmTlP4vlE145rOeTqwwyhilM01CT9r1JJ6JKuHEZq
6OxO/8blLkTEsKKWyi2U/Aj8bl2IiljjuSUtZsFPyMGOtWc0uTAqlH96HQywNSna
PLsyicbGIF4pixiGDh7eJ41xChiTq8O5vG8yR5VEpzoiS6UTAPP8yR5z7rcIfsXS
f6eCcqDqaiXB6LB+0FUqSBwoIg4mL34qGXZvq0Cc2jmB+glbwW4jsqCc45sgq49g
fcVkP1mqZSf6VsnlD7tCaQm3sUBYyNUhy1cwMeattN0p+1y/fKnexW0lXdpAFmKj
XgUgPQXASLlf6dDgDrwUlE4+30NYAVkB4kaB8Wk4rU2i2aEZ2Paa9+NWh9ByEsX4
Q8mzGyk/MxgUvbgtywxltjtvSli0cBijk+CmOUsnQTt+IXKgzPxrb5dbUAGf/b6M
ftRgwCzmNEarbJSDE3utjs6LbcHrfajYRjBnW95aDhT0ryaUZ6eA69ySzpTWDWge
9Yc71tm2HxnipBmQ9J3KJAhYn8iOC3SG5vFSbzbJtbgX4O2ra/v2knHhh1mhxm/r
9rmc1uOg1Vg4TIPswEWy8YNgzYo0sJgJ2aLVMUzxQ+2upgqMsNHd+3gKGq5CXDcY
NZzm8LKRjwy82IG7+ejoDGAxPGJihMaoZ958J7sNs7LFTi5ik1xPCftGxj3KUsTx
gDnmA+lzizLj/hIcbj6TqIkg2wtxWyVwtQl9YJzIXv+4EWAbFzqA6yeGvutQyDFu
Byz+dgDLEM3CATm2fI1FeoLGJCjDK7JayFODa2NpbLhzrewEPSJfyLWbgqJtFK9a
1wPknFrb7KbjF7MY5UnJ1o/d69enfXlGLRd9cOfJ8uXbGoXWBITE1oXoK0GjTz7a
EWCMabODHqQGE6TXhG0J3KeP5w8SCcGhjm3hCa39S8zKXODnVt8zwrrkP+CZJTDg
IK6/nO2OcDQgwUujA44ebCm3d1Tfv9ExvarHDtdXgtlchKQM9l0DfiSLfT31u9Ib
oalECimPIrGm44pc1d1eC20e7BomauQ+FlHD2vANQDOZCNvglwqcM7M4dEGIav8f
4urqvVXX2+qiXcEpm4uMuz0c1aX26daaD7CYSPNufSyp4juMcFu9ZN9UItKTLhp+
fh6QCEFt6CaJNsPcCXhRVcs69jyHXn/3pUxHIW18ETUJz7elL/vme7BmYO8EuqnQ
EvMFzsC7hT+Q1gmmycUFfMgx6ZK7g/etOKPLC4ceNGXDKkSiivq5xAbC+pK0STlt
LLU74xTpy9fDoDxdq2jsGH7SMjMOqN1L9b8AIufNn23CeASgDR6j9SufHYunOZj1
yE7lB7dgLBTZTy5gpVe7wq6/qYnooWghjffxsd+oNaI8ijdVb7g889z1yIzMiuNo
zv60P9wrcE0ERxFgMBdqUuwLt+4dn3NzatvqK3Wsh/giFAml2i8mGwVOYBUfP/oA
9ZLn05KtrGCO/33OsdDEP0XI/nQCJaPSVovbVDydxrdJ0Io9xjGMTdb/sHY8wpeJ
MjRXsDFlh/KxT94UnZBOeLGpmV8V7SMprZTyCIIgE2cDpQW/lPktOBI/HEs2jdsB
ZCj4DDG74gkjc2X/6tNGjh8HrJJy2KfChlCueQ7G+7vysFg3ZlABrOcV+8BpVj7Y
6QuLtMqcIlkSUSUO17Q2WAn/ii1JLgGZHnr4HxkQC6uC5taz+HclzKRFza5d7snA
NzWVQ0pOfTEddhVBdhiXsmIk0uBPf5BfmO24j/kgBP4Hax3AiiZs5+L96q75IOAb
J3iRm5cdwOF6wVO3FV4TEfsj/Q6gdzJT/XiRfmEBV5IM1hHrZdTtAQwfrQPjHL5i
ITgFw0wj3jlvfHBxz5VwYGV4vi8qhdXKQ6LZNNu05H7wuUOLK/vVXUYyYJgbMCaw
3KtEL0ZuSeMrOqH6wOpdkNsZdWLodTdlMSU0sikrhXd94xgxWvNnBeEQc2woaLDL
YqKxUygi+ra4n2Zi/+/4YdVHy3ET0i83oJYUAwHZAUaGv3PYmWzayXTX1p0f/8H4
R67Q0KNG1B+DO6dLvHeKptKVAMQG5Jq/3030GjBA20byQmwqoDanhEVzI948Hnbz
PrSuk/VJoF9dV1SzqcZVeVTjhNCyiTLEwNRumOF/xXvzS3g/+v6FIn2d9g8+E8qZ
i014ukCPhVVQyKOgYNFq7AWUpB4LbxY36NnSrMRd9ynELcuk0cp/dcaMI+ElIzzV
tqVL0ciFHPNb5/vwLX7etnrUyXb+GoF6oH6AkeYU+x6JDP3TJpKXvC8jJ1c8yx0C
E2U/VR8H9ieKMaYfDaKfwuRSUp6HAVqwOuykG9vTVq2CkX2ROp+W9q8xBttsZ+WG
jCJkpLRyx5ZIUjN3n1+cUkf/ZOsD6ywDXWqftDT7fp01GADN6b1CcSRdzCAOjHFq
Y1GoPpBntMX1Ol+p7uzxl93cuun7NagSbDt8gazSnd0pwXIao07ylPzmAN60aF3g
rbL2X/jBLp3eH/85XU7D1zBrpeEpf2P2QFJ2toP8yHrNz3cQdE4V1p8ul3Q8IX4G
Uf/a2IvOjArDisFVHWgiHSKsSes0m4t33LMuVhVFTIQH0hS+rdP6XbnvO2EbFzgn
nhBZqAJBFl/3wlhWDrZWL9YMCsPG5OzW3V99HAYR4IZv1VlqrhlkbF8puwAihTgh
INe1u/3GAqUWpjd9/anuDfert3OhuXz+UO/kROXO390QMWtWj0m91zTMU826Vv4B
WPlQ96fibWKGgBdkJkKxKjwu3JxLdCNS+9oj4LlV93PnRdILytH11q44JRGwQbLh
Qamd8RUZWTtFAw4Vhw65iBjjxjjvBB7PtcqOUbmC3u5dIHMzWIhSADxYJpMO3Rki
qyeBF5arzhb3xr7vrfhDPK/nVapg+ruOHKSeQ9ZVotfqfdCK09p7FOKd/sYl0jEz
Bdw/CosQwWqyQdwHBHpdMu2/shX2PLgBKrwSjazKXK4f54wYpO3y/V5Xh04g4R7n
K66REm3RmPPmfUceuqaEma66W7AbohhPkLfhmDhdPdR6CA6BoHIya0TYs4f1CDfj
AwDVclzoaTLbZuVmXy4Lci4Kh2cyKapkQtnPySqSN2SARIKB8IjJIy6RdQ0fItNl
mAFz1Pnifl4xBmpG9upB62OddddR9NHnKlF6Cc8gwh1qL6bprNS7yQJ59LO1s40y
aoOhhuzDSD9uccXm8Bnw7KvpHmSm16M/FLed6UTnimAtvvSae2l98uEPQn7HE9fh
odnsDpNu+jl2m/Ww5VAV0PlaHHRvktFEKkOeG+Pc8h0f93qa5Knbn7Kg/VtStLjo
8bbShaZFqPCC4aU7ECf+EkFyTRFRy1xxlTEGYv32oiOrz216Kc+yi8/xeW0mwMl1
8ZppSq29SK5Zo+1lNk6dEBGQdUtYMSc9G/czMazl63Ml14KhvcteHGfdBR09JHMk
fN0V2nsonl50GJLwNKKvvOWwkjSNLoSV5pSVCO692rTW3VF7MEl+6N1a98Tgw1TZ
MtlJnXj76WVXhZTUjwZbX/BBAK84Czr3iJAOHHNTJuAAiGhieUJ3iPvhrDviJ36A
moR6xj1GYKeqJlCClfMD3Xl8O8hzsXIp4dHn0Ek79A0OcZ0d0Vkkxt6+wegd5u8F
P/P420AYVFLwJ6judYZZUyhuvGy8dnwfLOWB1kwel6/dECUc/oZCzd6Hw/Nb9pCx
epyEI6DP35h4R39cNWfg6wB0sGhJaRDBy5pI0Ajt68cSHwPKyWhszzeJhsDZ1IvN
iXwBWd3toGP9lfYzydqoA4GPu+vE/oAs7L8DrVL73cG0BMJ0G5r3qfkGsc0nhozo
/rbTT4UcCutQpxSAE5EvV9tVfaKcnIUB8ZzoWDv8yMhyxCWSDM7x3m6lw8o/lat0
2ZaIttnRBbNPYdRpnqAt6crk4gsd5aA6+VNGhMgSl7KPxGDuBqswyZyEsZupBcoN
JeLfYLf1335IM4n8p6hzEkKqRxozHXQN7lnHAyr9qTSoTOsDI8pxD55Ew7sPyUmc
0G7cZUeVJ93TJ3in3DFJmi5nhq8xgeuUJ27CXGAfzh5z6FK3qXBuzzP41zk0CQLw
sVi1bSmztEqD9YO49oM/M786HUdnGRvF6L/PwSRoZ7V770BZpX2Z/UuOgT60XB0V
rQJL4SYKyepzEJ0U52JIqW9Y87KW4ErwYxiwMDbmLkPgL88586IpkXC7U6yNy7CS
+8lmXFFIxfQ9HM+zY8pLhMYRBn1DJk1pEGY/LHTP+g/h7DzPkrysgbl5LiMrmed0
wv03OujX/0YS5Uw7cS8RWp252CqfRjAzNdcSVpS7RYxcNKqGUp9OPSjHKZ1eTqKK
sN1bgQtKpRwYi16Opdpdc/BnCrxiSFGoJHWD9OPiYWR02b0Atd4jF5Ie/4KMaM0H
r125aGOpwHQQJkTcTsWOw+oh3e1UwniZX5yZpUsdjnMAMDzqn3o84bA17mt9GxRa
j3WD/P0MJyMLE7DUCTBq//BlJ9LASBKCqeBPSUcV0p6E9HOGBboXlxou3a5Y2gx5
v0DZK80pza+5CkVBjgKwZasp3ssjZ2g5Yh6WMfye2K9DjdUWMKQiZ17WM9XzowN5
OTLOr11036nIYgwpIJ5xMFHXUB7UVpjgkqgfRlRRXPUkEr5p38NehvjRrdVD33Xh
+MJhK4EwkLqgZWvVgJtJjiP4g38HEaQ7P1YBqcAXZOUjU/qJrsAYcjZP7XKjYcob
qVWtGpJYpw3Rt3fJkZi6wYKxCTWQKa9g2F8V9HUKc5QkiCUI2JwAsvureeVolWHb
haZ32dSWcgFEQdy8Ic/tiPk5TrtlrBzmnje7FCjWs0ESfQBgWog7pop0rFrYXEwU
g1wczs7v5oIy0oHsWVPWU8DsFpJoNRAMd+dOc1tXec/eN7G/VNYQQNJ0EdJONtve
ikfpTjBqoPHX3ary0EPLkesfk3nAiEjK4bEyWx28YImIx0JgdLRf8YBM5DdbYurc
j+w1Jj1Z2nNU/lTb2pC1S13kZRd6wxVUU3+exenQRT9aT8GjllS/VMy/Y9ezzaSq
eG9ww6dyXqfOdBVcR2+i51GXDSac6qsN/CDeAMfl2ngLdBkTjvZwUIEqiu4OQYy8
RsOPHoJMEWgX6acK3XQ3U48H7zWJc/CoYEDZhViMq+OEcm9/Y3Duk0QcjBA2Uf5D
6H39EjniiaIffk7f83eafj5YzqSIiGXnOLMUn5kKUur798DqqUQye4Sit5SRXZ+0
JBhpz5e/t+QHMyAL6QM1t528R0jDsoVzn5QrUQkQtOB8Dp6tGa+6tqcrcpMtXWkX
ww8k0QxoISitzb6JY6FnvGIQQrNzVkfXXX6XrcGG6DaJ3KCN48T9RAUMsXs2Jf1U
6DUdFAA7YUAgDq7hPJ8Om0ofNkYF+Q92EUqKVulyOq9Ba2MBL9HSAdWTowFxdoWm
xX1U079dpWTIroELYOnQRed9qDR+DOqgT6k2mOaKN+LPwAljcqw5fB1rUK+YC31q
mCdBEOB2C8gd56QWhvrWDYmtd/xypeFis4r7RTll1Qs7QlmdzRQOAahynIWz+fF2
a2EAA3lOAoeQuNaaxLOqyFoXMfbPkUM/1B3Fe/hS/dQxc9lnAtK1FvLTpdouZbvj
aCGIb+GPVCdR25WcpT2E0Chkfai7VkT6deb62q198qjAa3cvp220n1/K31Z9II/O
G1Nuz7bG8rcBDkRRJOq89qi6arZvlsOKC3rU1UjZ0hszrmEDvPG8VgU50QIc5c/L
8MV/PVCt8aY4TEugLBj0rf4aod78Xh8mJvNr33IIIDxy29pvrpcHtUGLvoa3EDAo
p4toUKWq/GOO4IfWmIeIlWEENNH7Pi9Y9KDeM14sxI663ULRAjeKl2mCoPa04Rir
q0GnhFJsC6n2lBoLjx39nxxDs9xQ3Cmp5pYlaSdyTGLq1gxYWvFIWifLq3EKqWtA
0JttaYNFOmWR+2wtxV4vufRAhxfdx6ztHiu3fOW9FqAuEESPGJu04xHE0St1eZ13
QPnT3eqSZZsDTnnof/udsRNq+VMRPzVNtGoHMHZBiFPXtwIjYwNYDWIj4eygPttp
hkBPjxAc6yRL5TNNMLNBSinrVjPfB4W68PYXJy9/ROeeDeD+I7mqlw2l9ZFeFDso
Xy5fFg/1gCa6poCN9zjHUkw8570XaUgx83tvHccTUPKfAFzd0ShFM1WYq9DC1zVt
+4K31d+7PuDNSt3jEuTF/BwiKqGE1yEC24tZYKUqkXWlHcS7HOKLN3TcqzR+P/a0
nhDBmE4iibEm22MissWwcGFTY7CQtkgyllpVBWVsEalicKKM2s+1ew/bYGFHkGKn
Exrj002qeuqAV+0/AvmqLsPgOawUH7A8Z+Fp99dmqe1RZN2vQmt+bLaRJPu0tWDG
ntQ3u6aVQrJZs0/65SsapsNOzrqV53cm2HHOrFUlYvtG006pLVDtsJyVxrsJEWmj
0zn2m2QsKdYaaumDE5Do79ncHQOp2GnniJhKYyEAOaU2V+FfqafKhfCIJhQJDzLf
SUsMxyTsKKnSmB/mDYNT6CRgpOGGO7y+cZEkoWShHmbpZfFeNN0ZGGd/hm6AmFK2
PU7kqTq3GhuF6zFTNL79KDPXw1VRxPTy00K71XsMSVP5zfUzEwwLvbw3MkE3SGB0
UtjAwnpZihNc4gh3zHBa/fYgbLt9J8HfMPUebEnmE/Kvs+WoV/pt0vQQsTBwYqw4
TqXGhD+EvNLYPXLsT5n27y4Z37u8/NdfMsWjQ2U5BnbKMsBEkPbxM5GOmHFu/vIE
wszGS3JfBm3pFTaYUHnrPCQDAql1wEY8sgGnURk9p9iR5tXR2vUdeQadmRA9DvUV
yiYN5CXpM6of1XvoV4X81u+7jvp0LyI8EOeQ+RyjazVMLQEetbVrXuXfsInFF5up
I7UM/iQvgRkO/1T3pUZFIhvqI8He2TdZfvti5txsGCMol7P6vNOz4fNIWFxS1oPM
zNo8rJl2mi6AfaCC2XOMYj2CBcHo+CE7O1JvbGpcyxhlv+CeGAmhrvrY43P2I+rq
JY5orqg566u6Jtk8Pvk6b1oOuFfyXFkkj7b6+8A70TxmiloKeo3suhaLr8JKhj8J
MW+qQMvmFaV7TZgXVqW3ZMFl0MDckVoNLS59MZLPDc5LTydXLl7UQYx2I5gT0Juh
YiwPhq8JkqCIzxwO6YfA/vzaK0aOqTnEv1a6FALqmZ85J99WSx/0eV4G+Bhl8VJv
Q/hf0uW7qlE+Zat6gOwvpm38yENPoSy7h6yw1yVZuloRlyEGqBlLFlTHKFz2GXhO
zxVwP/klOOnUvAyiOL+Nd6Ns3nApKMn/xSCpogANke51zSBjA8mmh8hxLFq2sPSD
7teNyxGjvzjlxZ2Z1UjjN/+xqS7aAPsvV8lRxwZdobzUa6+Ekrmx9mLJdya6os/l
Z5arkTI40VPjbNzO11wxSN+YvlmRBQquSogA4QAAHMB42jqcliz4llUD5c/hjyw5
vC3/IoFvqiUuFEdfTiJ08ZH3nzO9/VG8kdp1f8Ymp1xzn7yEZSneT2RuQD+DTWQM
i/oFWVkB/QRf+c4gWM+bwY3vnL/pBV7SE6RtrRUQqYftaYLiZWiLIGa5LR0ISXn4
kERL4Ci6RXWflYqscJlopdtG5XGn32E2Ez2VIgmZYO87mQe1P0lT/L9wc8fSpH6s
Idw5PBbWAV71k+6ASRMC/r1y3kWG6ZqQdq4qyoFwB3zbmKJxBmtUYAbnkxiQ9dxB
o7JjN5Jq2+lRgXfypm0S57HSi9Lw1v3t6/YyO1MLnH3ukl3umwCY/Cm3vKz5HG9C
iUYUqXSAdjl5Eu7kObuYTxpQAqDrOduZXLfU2IMOUQz5bAodaDHUXAbmkp8JDb9B
rBGt9WtZmey9zWdfEOOJFUyPLl6W94U/J3WsCIrj/GO/HURTauPLvXW21u/QXB1A
3mLP5AHzNGINIXAagj1v8qBrM2u1T0fBEmXm/ZgnVWkZumcEuAHH99Jxh6zgBw4r
oomVb6e20H8SvHm3tUHNMsQUxtoZ6+s72dzANNi1+7vP7GUDVLbVeelw8QC19C9q
2j/rMoaUIPd2zw6oDNU2GJZlQT8Bztm7AR/jSQJ1xrzqokpn0LjoxyFC96vir2Fp
SYkDtYiovGJREe+AV7XyOXOQ0KSHSdZRaDW+ByyuGPBc2IbxJ+PxN+paDGT5i0lo
IdTzWnOL5jm8pgfyUrARP2Xl/i5CwRK4aU/uP7nXXIKxrOh+byo5aJ2SHrQ7iWUJ
JAdN8OIHS0dljyNL5CM3iYJZDiF7xU0olVtzYlV+FreIxSmK5/h6+pTjLZqoNlAm
Vdo2JniGJKngwMfPTwQBMX1qDO2NhyXVqhusRKddBVx3CvPkNmiUqLshVBlJZ94W
cyY0+g7pHNxtPGay9pxVGTu/RrnP/u69eAkIjLi8ORYAuHX2uL7m9ryo4OAlEugN
UADEhC9kjWJS6uh/iZO7ToHADPcNdGN35+o//nDEpFRKjXJxsrjHVvDvP/E8iDjH
t5OhIu43O6V4S1YsJ2t2KMd1t1yd8do54TgYdyWX7sYxzL6Kbl9soKGI2KBhYnzY
67FBsyHAEAvD6H91JYE6UZwJuOBcLKxu904Aien2vItdeadI+G6ftvauisv7bA6U
eYfgW98x9exbRahQ0CCUXa7hBZCkVwwYnqar/wTDyBO1IRNe/QTVlonXJUf/7m8j
jfsvG4cVWCbGr5lJX89jxVCNNj7f0/T7VjAtkaYY7cEpDrpDPvIrky0AxJJkKqWv
9MHfjWHd1sBNbLc+oh7/KICGWFdpJVcsUSamfGe+g5IgC4MwyOJUPo26dzlgUyQB
q7Ta9KphbazMytxiAy9P0j1RV0xRzQi5DR1juug5+r9RvT14xfisFC4yNKDrK4lm
i7Jy5/yff8uF0VWF2VDYiW83ONs9EhIkgw+6BthF4ipdypbw5Hbae4Z9sF9mSG/7
A/1shax94CRGPHocQ+54ip7wLYXeXJVW/6kg9tUn9WreRmQpJkxGWVdUYo3TwEds
Sp7gHKfIIDQjzILpA6pV/J3b53IT0HHA6FXuH3EgHviE7/YsApvGW+TY0lOujVLq
v+VRjAm9nZ1sUgqv0vlr3zViG4PSyq9YZYU8Ci6J9crj0tXIpuUL+oL79/RWtC+s
YmPYOlYTt9iT/Na8jBXpMb551VplW2luCNYoSPFh9OIfwXjlvRDHUGo48DkRwWzi
pV1NDm+/3AYF1hIZDu+hJ5CcNEUHSGK5O1eBKDUOVUDT4r66Y0GLweEIKfeYhQ++
fdn5OcjIEpjOyfAhF3zYsbOZSu4jWV4PtytWIgm01T+Ug8MSl7h+226kOv67bu3x
ZGEvnHvAiOFhhGP6Wbwiigpa6OmG44WOXuaBf+YopOBqMybo8F+83fOVnPN9G5Cu
s1djkONjPfNd5s3RXJNtU6f8scD8nERbHscyJD7SYP1g3DJEoCdXnY78v/reIXrP
Qe7230p3Oc00/35hwS0yVwBIT0jtWwyiYwO6e5ZXzRpC3HlD1UeaafxyGgiF2zTV
ZdHBOmP9W8BzcYubLvojrxJbvEzjgSMBQ7NK/eHqLV4tjtwYUgfR+BGE9jnB0sRg
YXmIf7tnw0HdwckTrIB5LhTfYWFthar4IqQ0qL+hKTTa30LLuV3vqtvnVUzLUy5A
QoJrSRpgZHNumTBfm6iFfq0Tm0ZkrCL7q9Fs+AtrGm3OCvW9VOBW2HHL8lmgE3J4
0K+EHnwJrIh+iBTC7cbUVP1Mh1KuvZq9MEd8mX1/zEfbSI8fusm2BLpISarz/YWx
Gee2B9iQvE9cyyoKi3EUM+n8T69ZZJbq0esVT8ctFfdtukV80mxi36XY26y8I1cv
YV/hiOvw/2D4KSMVj5K7igzn0g/ZPUXdz+RR2QEDrPnIcDzWbp+B7xqZH83W3/3P
8pKApZt3MyaMtWvyA7lzvHtJOuLg+RyR6mMDgdgNSAY5hXxSwrGm6lkVNvzAjbOc
5bS4t3ZW1R1ceNM8//FXom8jAwOPjkda+5tWoyxTA9ZVK/XNznLgIP4LKgvCXpa3
yPyPilMFMb4sDs7aIVm881AsHgVp64rDQl7xVUM47yanLVKbo0/qsG3GUX81irFe
5WgJOlI8yLhQfAgoWRxHejrKW97u1fDnKhI7J666YGvkBJYcewVnqxADE+t5YFm1
4FsoLCZmJlBjuYDry1SFkEhGVT6/wVecXOdlsBBRKg+cPRkmOiG7RmRcPyK806cQ
V5xMbU2a2L5yzgf9lTZPotywXrvb9+2uHH+9QYLNvUyBeFt/ax0srfuvQjV/smHQ
kozYSZA2lmjb/jvWAFvbzW4VU8iGFUG/CBn1yskvGc/dPSf+OYcJxu6zwYmiK2vw
4pZvm6iYbjhkR/XSqTDenDjD+xx4zbdSoWR3PCIFxTEyyE+DjrGErZAn34pXwOPA
nS+7CTWspQNTFxTXbihJjLg/dGAqrN8hV5gzR1gepm6s7pqUj3IyyCAowuKn59sZ
ZHpsR60BsjLw2ov4z0GL2LL1g8omMHt7o/aDWHmm4gnZyKdFIHVq76/aSERvRdr+
yivqWQJ9I76ztbgsxmV097/W17XrxGlfkRkoxHUlsXCtecqMFdkuo3lwwuAG2n2L
HxUmu9jEzb9li5ua0cZap5QlL9028jTOYCKrXxokMbfUSqRD1Sqr2Y7EkZPJuyIj
8itlsfaOPRURCjfnkba9ZduetFDKKSvK9j74U05rRddpdMZbociclgGc5e0UGnr1
ChE25qyiWCLjB8tvf7TIbyZYlItyZvk3sTqQhNe4v+7LKNKNWHbr5TC9NbpN9Zb+
G1annPkoirEZJ35/Qw4aa0HtMrxELh/bdcWaRJCl5Hjgtx4GHTb6fuxsptWk/grj
2hyVUpk3YJRnTZi4XELXyO9S4iOwqXbRFYnwCN3gd7jmY1oM5lvhCd4Op1z1VZIj
eo/5rxYf2qUIrSc6ey6rdGxmfjDMKbefmrInXUzj3F4ybhkEbq26gpncsLKOzGxc
Rm+43vXx+ByV8n0q3pNUFIVaRyr4Cs9gDnmwgT/KtZFtfeATiYMu3k1uD7fRpZGj
YagjLxfnunFkSt7A8h8l9Qtcr2CoC6ZfwH4ReZ6ukHJS+FxLY6vCPqfY/EQQOH9W
8cK2o8y3/j/WoF3ZKD86ciUhUwAwz5lSQyzn6lUz0QIFIqgTI3hMyBvoyyzlnu3f
2K6mETqv8J+WLMuToKKoTYhFvS3SHQqLgAzltHG+0Y8tviDST3ko+bs6GrX+5EhX
Vwx8+VqEeJ/BxTduzNhwj5pWGChmivw2S8S8bYjA3mkZRc9JtiIHAkScb6xQMqQp
HYPFpHh9h1rUMkeC3YKhNYR6vpw/UZINet6nRxbMDRlHpsmHS6Yhr0kLBrkANtbB
0cAcJ+5VpQQ+ucy2csOlvp3fjJ2oBA95Ij8/KGGH1KBLSIhssyiXFNeXrjcefJj/
ZDkZ2bqZ+g+Di/Zv553smUhrY606TukTb/QxCGSuX+vgkQ6JMyQwlhzAdzU6IiE1
/N7XIIPmZhpJoJ0N0HvUf/MSJwVstJ41aeiy8l8TflGCAqaB5DqLLzrHsWZlKPX2
bUQUfsH/8RGOwf4vgYYhIb4Jwzp3u/aNTMU/nzLlcTSjxkKNMIL1BxHSzPp5xwBg
bKynELjfO/LmwwDWDgdSSxrAQTXT0bI7y4CywQu3nFcJSC5B7NUcTwROm+9L39Ov
FJU06Z7E+D6CwCSSUP3U0xo1GY/MaH89mZxgIDgNUKCiWTOtJ3Kl/yd3QG+53hm7
kkRebbFfCnigje8MPrk6ApmMo2CnWAQnmNtlizynlmKBw0oTNeTCgIhYvEJUUSgM
AaHhgFYdRSnwBawAwtVC/DlGZfYfyaTD8brmIpPZNGmY6JVIaqdDMv8GsYbufjW1
mON5eDBE+6XzrVQQG1kbZmxZktOL64ymoJ8rkX9XTZnoEBMeoT6nlnqauDRvb81N
DJ9HEiACEM8AoJH0cDK8hXWrXzu7WlwBqeHjbota2gvo++0dE4I3nTclhSDmTfI2
M31oy3jhDvqULnKqCPD281xmgMY5qZq/zKpLrJ7ek2d5+8BZPJOzjauOXzcLlEF7
ouaXAKWHRgRO/yUsiuLm/cwELBjHE+bIxS24BF3bsoDg/UvqRgwanXbj2x4jPJ/j
JRZcEp+4NelyEDKu+y9Xlx9IMoJxANkhPcCHJ9Cd8nRWw3fYbcB2xmEgHlMbj1C8
lG0WySbRogrR/EbugYSDXO5yaaIaAqi2dafP6ZUn2wowuelXzM1pn1/keR5GQd3V
lOa4NwD2LCB1PkaS6Q1xbORJLFiboE11zcKf9kqHZQ+ILtRHUDaCL1Lv3xykD3Dh
5fc+zNsvlSecY43qoYJZAb8ONcR3iWa3lZ0zf2dFp3mQucpRTb4u11lEE25vPKiF
nt4HKHGIdNYoV7B2IUMWN7t32j6I7j71hnpHpS82gYW59kBtW9zPyw+CXa6abyuf
hJViiq0U8CuTixjx5Vc1Bo7F42Pej8uTkMi1++to9LG12BGIdG5roM+HUHbb/5kj
CAsXX5wbqg5zaIcksNKU2U8GhXZMPF4hcLm9EXbVERVsAnRWujshHcVNPTTKHhad
4+guvhctzC0AkOc60FfmyQM+jEDO4lFraVGlvPyJlH6BRaI1dX2Q6uS3WAh+/kl7
8I2FhWwyJd/nDDNEbyYO8/jnZHOWe0KuLFKA2vU1SAzCRyaYUCWbLCHwQkdmEp6V
qVZWaXNFO0utWhnpNn9wOxMY2l1G9r0XGwseDJVwwK347C/JBecdsf1bptTE6uOA
zTl0NEijycIiyYCXxYiKcwgTWdCu0G2/zOJWomm1lXpk58/0DOK84KP0p6brKHXX
djvCys/A5c4t8ifUPk9FRpBaGnfbjxD3E3wA46WMe2ZgvSklP2hTihhRNfFZcfw/
R9ZtNOJPOJ/fHytkfRfO6IsNK54mMOja09mTKKK1qEOIFRnbZLgMkmKokM4gd4dN
mUXcX+oWzikT8mnKk3HshxK/LtCPxeVVZKOni6Zigl7ULeZvbbb/7X5MX1iwtRt2
a9ZpA7OWrYcPDI17HEopF9CpGq9mL5b8O36Fe5XAzQY17lzgWK6iHDmLFtJItTER
3nzLCeMp4qcNEXYMb1kUbqmy/x4A8M+UJR6egc41teE3Odb3iAkqnMG8Z5c4nI7n
blCuH3pMJHnEirSQYGgdvU2m24cYbBTsWA87TqrZE9iEMvm6L1toLguPIxY/WKfW
/PDZ86eSysryGM41Wajwq7NMZNwjFDZ8O27U6DkE81ymZ/1x+N2DTa8DKpZ9agCn
HGW5EagrJbPhOU4D3W6ar/o4EAK6BwMOm/wA8R1CTiC52jGiFu/uUveSPyDQiDZB
kC4/+Fr0uWnqPGlu98tHZ9KeO88072vhpiEkGC9onhZUHXlwju2bu48igM3wvQ8/
OckIjTCa61RnYV42BUhm3QrU5XtD4OhyBsXXLMeD+MJQVRl9UEr1epOuk9TapYjc
hNvDGxJ6a24IqwrE+6P+h9mqfF+oOIn4MOmYq5rKGYJS6mjdp7T2xnziAtU5Ax1g
mioPD34sGPIkKkhXrTdqjFTJvjPxsB6AjD9zneBPmi9TL2ZNvb+dOMSOTX/MvMHk
vFd7cbfhBqoDf1IEFVtjtzl46c9OuiHxraCVHnBc4+HuHOdqra9tc3bCbC2QVybT
gsU76+zXwyS32j/LUIR0Ke9h4q5x1gmvwLzlZQzZg8wED/Y7ircFsZ2SRdbdEqHG
pNnxevrEhnUKDSJ0lYAP7266vWLi22UXHjFCU6AUZpXUJLTu7fAtFwzCilns9982
8kHEw09ERFxrfAzwQKwFfVS2rG+K4GuYkMMmwdQWcbWw2pzm23LLzPG+8C/AxV8c
rj8MVgomKF0SC5bw53E5mLJKEsyrlxmDpJ0l7ekEDdzwsUBbm/zXX+DDAwBKc4XS
qQ7X5yO1o1wyRmXf25TZGgwPr5LnxrqN8dJJRUS2B4oDIL7hTlKvX0/Hb4yk7dIt
VX1BCEUhGLpUbV75jkVtP0a595LXi3CoGCpPhrURLW+diT96puTQH2sNxHQBQocC
83Eptbr+7Z6zYXKoP/69E3GSQ9JkIlZM+SQz30FFPvniUg1K+dSbXSU5d+kCPiK2
TihHWdwh0m1iF0nbO3z4HZunXRRNQchD4OFX60QkQUKUCa11dtTqrBxefZxKehNN
kNnRzYDoX4QGQMOvB89OnyThkC8V24zxIIkx5oIcNkU1JY7dAFyQSXeuL2fDScuc
KjcZcFKQDq+WBiGY5qjfxSErwp5K/x+yqROuhtzdmHnHnnK3GrNABxnzuYX1lo1L
kF0O1nUkhdYzK1vVEXajwEGhKplmhrApv7wds61lRIQGdsasl/VADxICxQ/mBhvr
GS6rkL68HmgsWu7ZD0DJ1qLT5LM0+Bz4WHpmoVHkuS8op3n5xk32FjlJNOqEcxU8
5bwQN9Sh0Gs59VWS8Mo+FISm29W8ukzVCLMrHlkq+AAuFN07JNhyUH/tuLm/MsjC
7W1qyqiCcL+PlpwHCiVLtZmTGDr51OLlrFTqeiAu+t/6xUj3ct72FOQmNVcO6qca
A9nthoE6EokXOFH0zcuwy09HCKxuwZs2ZrIqb9As57GLBq4Z5LE5RYzXjkTbode0
xcjsRxTWE8JUlhSP5CfAXcYUK61u4Pjbn9drV5I2moB8/pi3tS6lJWxFHMHyWJDv
2RnPBx3WhU/BHundf7BRXSbIE4cEPrPObN3HAmzpZ7dyXnQisYKU8aR6jaVpx5HM
Oiev3k95P+DTH6h24c6hlAA3i4coHcQcSxjfq1vjB8Bo6yXXmvLfhRKg7UDrUvIT
7wlIKegcyYlvFPPmdg9c25rV79JXt2S9wA1JjDzWejf8pWwJXHh2l41cx7cJX+IW
n+WO0gkgUKR1qcve5LjAUdPBDANfjmeUpzA3edDH/4zLmMmlnKRGabBK+nWweO+2
f+Q65n4hh56TQ1G7jCfCZOqPz7FpCmi1VHBZ07ObZ1ua2HlV6pU0vsvivurMFZ99
qtz66JEG9afY8Q4cpi1xFU2hQJ8Y28vKoP22+21S//ScA9WNFDGJuim/jm/yJQqz
w0qSrLFGIc6c+mzELKx51EMR3F5qW55XUsCe15i/D1Ipnq8pHfDV33IKOEr0fcJ9
LoUlGwE21+t/oMc+QSvjz26PTSrfLb3JaBOyAUlkxGnA86GDAhBUx8WubsqtpPOv
5psP023J4pDwFH0RCPE5cg4j1MS7bLddd5O9QaUpHQHvRSWv5eQFBdTAE6vr/YrH
e/n7RJ8tymFC2FsJXyky1NBa2zireEYRyqL5aS0lXHFHm9JWapJkeWkBsAOPoX/p
FDh7cgw7JlKgzA0k0t0f40JoCxKC2qJV8oxgk86YK/0o5s+fQSDx4t9Y0PUfARhI
fxQpWuqCmkKrpD0sp+ndYIFPv21jbNvLQLhd806vacSVFjUnvzysB8cV1AeaaVHX
rVEwMZlZ1LIRV6YRCGcWGWlTyDSbmVxmX6Oq/ozjBXv27OWlipygCN/w40m/n1Ob
8NuUlTHu2RvKyWyyS42kKvGhlOJ9T3KdbLfCRwm2f06cPLGB/DuVTfIyPR+ho84o
n9HrSV0D94bp+UvNlXcK3un7oYDnmEzrcZrl0Q7wZWBCMpdUHY9cISFeIHm0poS4
DT7rs+GuWpn7NF7o9Q/1o+CIFf5VtUn1v78yK3x2vDHe4faXMbX/ITKnvZ3vno4K
uHfaKmE+COd5s4dzEZsK2gcye/k3MjDLoksAG0AcHuWoGv3aTiAvrhWBL4uHdqQH
e5qgttKIYBbvLf7LxTg/sA+IIwq21MLPdFeGG2x8nZ24G3wmGsrnUMgoLg0MGjlR
N3IXon7v9rw6wbyA/QBFXJWef9y22roSELRre8z4CfH8JNOG6sgJxTMrIeDp0vue
Q8biMUUGG0Q+1T3B+lpV/uPKleuKyRw+3N4I66iTB7Z9CrxS8Exd9PF9kVBgkj4I
34W+rfMv3yhPbii21jRJGvTB3zOn1xw04JUYKPff73mV8r2cJdjOdoNOBCiNNBNF
OcBNl4a3VQdTutQjwaezHgE+v9MPrK/MMty5cqVrcq0DdwlH/dsy2KyszT3mGSqD
nammNIP9m9ogFd+jOlwx2AjN0eEuebZ2GLNRXV2oUaLiuhcbXW0G32V2v6vEm/si
vGsr1ngetbm2bbXxjf3v+b1RU75cYzTnmN8p6iCPKr9rf4M8dq53AzfWH9vpsWBw
ksLGNVkgdyGwjV2QObFZ15p6Z4K8xWp/0HH3ZPshEbLsJ1W4Oeq3h+9aUvLEO6cu
DBWs0nD4Yvdb7byj/OfLExL3+vv3kL7iH8NoPoQ7nPP+A/LjCKqH1H+fuAl58rUf
Aswai7Gfz2Vre1JKKak6Up4ZAbPlmToLl9jZDEhZaqUQsYudQTMA4UrMQuAiXwD0
RXqiadki+HlilAZZLW64rJQI2A7ImASfictUsPqZQh7WAtxGDlQB5yYm9GjN8xp4
EJjTBIUG+aA2QbP2XZBPjQ/W9PZPB6fUyuPcGp2OcCEZRX0VAkHgPLlBtFKpi0HS
OK8reuqs5CTPvIreFPaPpMRgxdCZAPJnRs/WggxjYPmkbHRGqzvjE+d33juQ16qB
9IrqT5JxJkQVfCD3gQTcfzGHr0u72MRg5cYTE8fxtLd9uAj7QjRxv85gK2VuYLMd
fNwQN1cB0UZ/7LwJRLWjKjk0MYQgWblagel/oAOinh6ZWppbqa4w6SHR1Q6wcA+z
GEKG9x7oI9ugCvubdDpbL+j7idkCroZFoXqO2NAXUlgSfF2Zmsv7s26O+SzATjXX
qhIsMDV5zt0MV/GN2kkEp7DM+DkVnDpEgVxgD+DZLy7aoBwS1ZgZ715kXInzAPSn
yngao64vlY3dMpCA0qhSeoT1mgNeL6bXQ/CuhQ55IsXoEVJspS1KtePJwmHkPACE
jFIedVeO+S/L1l2g27XVpL0oxIrLaKOEUxxIDoxXpNM/Q+3yVvXLqABJIuix05eM
Bbv2AqYhCMrdZduclTddiVvDYp3UcayHgPyuKRDAXz/p2jcXdLdGjQZ4pGPfGl0L
vaubC4XZBdF3fPIhBgxrMjHYwaKYWk9aFMVvKOu624xyt47ND1FI+aF2ijfxmC/d
3n2OmqcughmJJkozeYAwLpavwzRv0NkEucx7HdGiNtSe5QfGpYjLsnwN99L60U3h
NplddQvkKpqtdrwOguYvI5lndcLDn4Seh7Olt2Thhroe6PjJjPgX9JHVmuN46TFO
42AtIaWnNzUoTXEhxoaTp/+s48dP0k5GPVugZS5krQNmEif4o14bHc77kRUZbQcq
T5ezpckaqzdW91kNMFpNgkwk7TOdfdiC1eKM125AoJctckyv12LNOmH8WS6fQtMG
XD2xRHYHKliWaAQkrFprBDjyqfRZSAyJLpeiG8hjzweZnzrITp2DllOjAZwC26X3
C21P+35IpckByWb7v4ZELAC1lc2x+Jpgt3qSsaFOGeVhGrwvi2rIcm6Ksce5VEI7
VZNjeX6tHm2Y+lCpnEibzOnniHzpWkmjHfLovaZ0V3McjssogQHceMmoDJNJv5dN
RisVrXlFwcZnA6nyMw9Xq7wc/TAfujT36EnG5FkhH7bcmiETFOfF4w1ELalz30Gc
DmHGBfeMxM4qPP9jjLqI17mIC1UoFr5MMZbb2rbRBgWU5QBHYiuROh25G1IdZdMT
/qbhRFDCI8F86n5TqSj8gMYj2gnFtcJS03NKM4kW9H47D2Aj63/+Dl1GSr1lLxhq
gZVRDPYx8oPJFpOiSkLP/2YJqnkC0z5TM2gSrUowaLNhXATZQ2HJNVIX7j1raFyp
YQekdLn0NNezYWmHLWS6WziJQ2VsI/aJnn9L8EFIQYFEJwe06BPvEWto89QKzCtO
a8VJhAUt+7/njVUdGV3I7yMig3DGSbn2gg0mrzH/jJBTc4OratntxD9seRfssGMz
f4Ivge7xxzGqwiHutwMJTGBnCB6Xw4G91P3M7Dg4E79sFc25b4oTDRIY6UuyPXrY
+r/8ZWx4jadUf+p/8ikjGe23TVT5R7Sgpjv8/lzIoT87MLycsKs4qZIq73HhLa6N
FezyUO5KVq1Ur9gyuL50X5KLUXYYm/FD2Jqu8bd0QNW6gQTKQuqrZv/LngfT6UeI
g55U3M+YYNAiWFZQvXVckfQTpWfu21jipBD+rkLjg5l+pZM8TRA4S1nE8WescWnn
NSiaSs1MQ7RPJU9BL8QLX5cQ2N3x9XEZPmvFf1UB8xLOUeUO3uUBXEXkefbhFoi2
c31KCzvO3jO7sY9j6lYgbc6+NU/cyNkEsbKRA1MTVku+QsNaqaSj+I9D4JLPz70q
A1XOL3ocoMnWAdkW6b8K6uLJT7OGzYC7Z/3g7eKNs2H5D71llNFdyCN/n6Z5NLiB
5ttMnsvcOZnT6grajr2oliLJFGJiOAcQkRghpj+K4fljtvmJ7FtwO5wnV/eS4++L
EBE2BECxMn5EcTxYPt5QFQu6J0P6y/iZFvrC3GIdQOUrqzxdanoGwsdDrTp1m5I5
IDZpKpbx459hWoyPGSSI+lqxvoRwR2duUov0OdCzH6OluA+P6yuLxyxz66Tt0dC6
ljPsWDhm8tDcKRUuTG1lQmeFDZcxNuVofCLao1OFcDoSQStWg5McSrRt/9QcSAWT
SzjSD+8jDiP/C8SgvFUhyAnRFknpdDLVJuMeU5zwz3OfdOr8T6O9CsJHTSaO1li7
zK1b3Z1R+3HHrqfhd9hZ/wea7ZLDyn7hIypwTaK8/Jxi9CxsLNcofdEE1a5/bWsV
uwSjCNE7OGajcvCQipYh8JiL9Gstnf5vW75ROGGqaSiI0Ok30U2J+tgmQXYkTduK
hCbu+hyTWlsIoXJWQHtiq5ZxH5cQgNMuQvFAjNUzhEqfnGqrgJo+N2PNqXhTfLjy
IFER5krBWILCtqkcT91PViWZZuOlb1gg9VEtvku44ADQfE5EUMU/+Y+4jRglnQCG
WLhxtNM/tOzsBh0qVU2IiykDzHuNfhSI0ZlzL/wE8g+s6zmCsW/Dgd/+8+IhD+YO
neaK0u0hDtnmXH3dKC9n+aLnNvh2XF5e2GyLPZzYS7nzNzpI5tCZzgR+3tPnNtZ6
M0lrYH8fBAo6AlEtToU6W1N52PGmTOjwJeFhJvVnl8FH2FNSSMwEC+0PDsXBdqH3
kIKmSU4G3K3aiF+EuLLpBJRMP6GGzvmh9q9Y7Coo9HUqDMnnl/cB4YfNcvga+33h
tTPMXLUGO+E45UgUzS9H7G3UUNV8ezQZNW9ov2csR/RyYv1Nm/4v7oRYNxGtu5Tb
alZCOaTZJeSRBLVVcunYo0IubqibJri/iMMNKogNfPelYvKsabsbK2TNu5g+vFFi
dmJaYPqLZjgab6cBnXAvBR2AiHvFo46Yq7gDe3oPXDRrU1KduS5c9BuyCDc2oK2w
WHb082v/1TjAfiQgZ2LFvHzJ1GJ4dAriioxTEU5YVy3biG2/diyUL4c/JoxP970t
49b/aOoUIKQD7enW82gsn4+fYpJ3bDgFu5CB3dAfD4Zz/xmsXcPP5p/19mLAqdTM
4qHxFjt7fCSaFTJFxoskAAE2irdxJOCUF73taV1IViIXYOvtPoKitjSLJ4ZNOLzV
N/K4tVkH/UYponKlt2MHIfjUc+HFY4z+pMf0rwT9ktiaP7NZQMiX8/S9vs2pjVTN
uMvj4PlkBkO2rZ7iDN2yOHD0fD5rQ3yqqEVqnaYHQgao8FBMf+Wwna+gmzb1BSNq
3NLmc0ufSO6wbpBpxkLQakaus99k66k1IDr+95vmK2MR8/As0CQL80q1VY0r3MNh
P9YQUOmRHGMSfuKnp0XGP4PHvBVPDWWFDsdffeiFzPAlJzgiNcy+QorjsvDcbTB3
42PiXeImQjv4xDW8GWfzpNuTkFBoa5VNfp1kxfxFCv22mZqzPTHoduFzEFhwd6/t
p4L7bLXzGA3/jzHfTatp9QNbdY2RQoq36Kqn538JhWpIaqZ1SWiMj4Aizc9w0beC
l/P4oUTMpcs+oSCx6cDFk2ObR4gR744E8+FYGnxOLCgyHqEn3SRfFqIJiVNarQ1O
ClUGTme96K35HmnN9Du6bD5MHEBsD5zXDsn5mrzrKaSvVxLBT2QLikOsZVox/6kd
4dpPwU63gpziCXreWUw7ijLY683KuOMrEboXZZnXMRIXWE0bCqCxrkUub96mJH8X
61ZvCvQF2/a7KVf38mnHaLOBkY83Dvf9Gls8ppY+vN57Y9Xxy8ER1pSNCphwz2ZP
+xCJZHNt7h7/2DvY/c9ZXe0VUxdjRaHYRt0Qqp41ZSJNJcOaa8UWpFb1HgJGDove
FJp+G7/PgtvX7JcCqVsr6BrhcCu9NHovZuWXrlWkmjHTz+LNGsDOu2p0aN7AvQGi
7rXj9LOuOeRjbv29F7LAvui5ghNtU/6HXuelnah5S3ojGNi+jichCl1on6wdh5fY
gRuwyl1ANsLBK/06NzY6HNBhlLEIfZG8aRwsSV3AvtwaCVmZukkyKjzBwCnMTFZZ
1fY2DiHTcalikmntf3SIHQeRU86t74CIjT8QoqybunYoZS4R3eo40n9c951giB+7
sqtcPDo4vmqeOfARSOsKdKYMzFnT6rpZH2SZlinzVI1prVMiFRl5FGbTntJd0Sbu
eK0+mlf18UfwazswCgtwH1QV7O/44t9VRx23TQBAw+XQzgb6/398ECOLsjv8jU/l
Po3dFJwQ79g4NgxCx5n9ATzUb5qprch+ITv4gKU0TbOXU/dqnsc3NiCxGVGeSCAv
giuwMytlHruBFA3vsTqavxDniElb5VN/DqvjkPcfdij0/ZLzt71Eq+C3KEHigF8Y
DcVfx3JKiCXdqgSQ2RPHHtvSSWf0IYJFuwtFLuPMAkl6JOcoPBPp8Jd/o8v5OS4k
L/9U350Bw3W1GqV5orIBumU9jZHO1tmSKJm2PAlUk7az/DqOBEoT4ZnvDaK/aevK
qQDVrVtFKRwL6wc7mGmOLkjKdXiXDLaC05cgcWk1KzXx8u6/UBo9TaYQnQUeCnqS
/2fRq6+vU67l8XfDCE2JUnUZZkDFh8lQ/wtQTWaJXQ4y5lKniCTG30iMcs+4babJ
Ep+ErOhhczgJNIXohmp0thUT/ZijMuRA6jPWPmprRm8h+fLp+qgi7F5tVQOiY/kw
KlhUUSG77PQIqm8Kq0R/iHpOW4Rcvy2vjYLtCFxcLjv2yCanV+Zl0PvN9bp3oQv1
hfLilspDcPc8os3hrKljiAxIvloZOSnkzRjtLYyLobEiqME2HAFPe9TFLLqKE/OI
9xwtR0BdSMCXqJHilxeFe9Eyv0i6EuiUlgmP/3ypribB0L7MpfLcppdk0IiQMJVO
Zs3CNBpCWfgtFTbEgP24YEqH7v7FYJAFTUvE1jTXN0FHC51yzaCWjt2PkjQpgoFT
lNNhXj5oQhh+nXIi6PU7T+xJCYUCIzir1gf0v06egH36tOj5p73fcq5sXUtLfAlJ
ZjA7XGSKmprePFgsgiJtYIG7o9jTMafZ5HIBK5beBIhUz3o+Oo3gJ9iVU7SolzQR
YK8W3KFlU9+VvLYEqqaW1yC72qdqp1TdwJWYuA9OaISamuyMnoMljC0SjOE2evaj
aXuM28WTD6xm/YGMsiSfrV1oJ1Oq6WYGOxCtkUWchlrOKex1uHj5k7P4c7cddvpc
plfwrqpz6A8Wxhc3T6psb9g/mBt+r2jgpes6sbESwrcbd8RgkiHbn1i2539IOuv7
TekVc/35XtH5YxCnnZcUzn5Snlw0kTRKHeDGHwdmV4AW7U7Bb8ewR5eLHaoNG8Kx
giPzJlXuGoeHrYNBaQlcfP+/8y0eDORheD9eBzn924yefgpHNOXJCe1fjJtD2+2P
gKxbuxZPEYXjr9JAp+NmnrSq9GL8rEzb2EPlM7Hz+Ed9gHclYJ8qJa/u/5IEeT9i
fYLwrkZDrajaiCcMMrixou3bIPM1wHxot+AjavaMaAnUViRUukVWWmY97FmOiECE
BHfSS7s4sgh8CRR1qYW0OQVHRTXvvdCJdjDI4FREH+0H6pBMpdMMEjWmsv4+QNsg
kgFEgZdvp1P9ggfcaw3MiA9jUb4bk0CJ2lMYuQOeHr4De/R6pztMPTBTg1NXHTvo
yKkPBiYVJCN+CVzEds89RVdgef5ChYX5Aocf5+Y9w0qkM6ZBZjAS4IV5s0g14O3K
+FIPj9AuJMMb6XY0I9SPkR3DmLiVemEPde06lXHzgxss2ExacLUrQV7a+Cd1VjkT
kPv1ubtBtx6JAKA2kPbFwhc862TRP2kSpylcG7yfS5y6qxVg7a3zhwQCM7Te2IuO
EYIPmLeyVrc72at5Rn9WYu1tyzvz7Mbd0rURXkd85ofHNJQTdibKpRa/U7hze/rb
5nJSH9SB8BpkW78jrRYDDKVogT4hR0zojyXmqpxdXFSuVrAaAgoKEMT0Tp5NK9Id
d/AYouLKk/OF5W1UtobQjclfSEJ6XlsbMDN7QuNwrhh8NGrAKUIN/PXvoolYK0pR
Shzjv89JPhXclYtiv6SQ48t2c4Ub0Hi4SaDPcMjXwobA/hdU+GA8aoe2R7xn9TSH
4HF1vPicybUD5eIc5V9KDijRuIcGT1hwfzIwN3SltV10fChPqaVXp119B+YPgZjM
wkXfrY2mYL7y883OLLIjGjv0jNHqT1Bj/GprK0pldVxW9jsznomhEvXF3G8AB4/c
dcouPKNDAHggAC7XB+kLYudGVEIHu1Yp1dXDTGMZqamsvQrAn3EnGFkpX37AS8dG
TQ26fTSbRRfYKW49FCypHSSQXjsqAIxaSrIYm7TzwrIrUqSCxy7+qQuutSaESUYY
drDg+G2jtGgAecWz6CWfPPy9tnFBSdQmAeBuNz7VPssFXhF3SogwcmXTTCLCUiI/
jKgByhZNRfbIeJxeFcwvLlXH7w7FPoFf5hJJDZ7Jtippi7U9Jv9MJxGlr9X+QuxH
/7q9uhCd5d0EbWHjGDOHojJSgJ+2Y2zN2Pz5Y2dlMMCxgFeQ24ceOdyoUDkaJiI7
6QXk4/X6x0g18uwXBrwlJnqU8e6/dQWOD8g5g8lL+jyRWiN779jOi8KN10bNMXic
rYbgD9gAvBeJLFbq4XdvO2S3HtNowgDDeZnGi+/AEVLooeQa78+9jMtjIMVISyfL
O/KQWubNIvgjdggh4aQPJZliK+wNgOJFC/Yy5alyTsnPn2zKVcychoD8M9e4mRwg
ZlalwpDK7i7KL/iDZGelb9Z0bXMgAggGSnxlE31I8MmnRLAhuFUWmoambnoOR1vm
b93NdYDYBQPVgUbONOCi5Iv4uMzruDJFx7zI1XGcIapFs6hnKPruAyoOh/Pr5HsY
WYKDsUvNrhPbK6m/2MRu0ohb2sc+A5WjUFvHeowohqCZm5kpkVCLh+PQn6RoeHc7
6B/gpVzJ9PgZ0bIQxzcrYOsetRpbL7yth2F0Lc6amB0rJ4KLncJnaLk+0cJHU1Tn
ET0UzJ5499puPEvPOqHkGmflJurEChYQwy9tzkfko6w7WMBZn2R8XFt2wIkNYYF/
pKhjXMTQWigDPz8PNtdrvQtf2nXtcxOg0CA3Wn2FkJWp42h1z59xL7RWRE59BLpB
9CtPWz5orqaHqiczLzRdy9TN5X3WFo0VcZh/34rJVuYuetWWnSzYsZ7Oas7tyYPo
p9CeeZwqUKibJEmT3b6JbvDjN6kDl7WtwIT55O7g987Mty90KIK/FxMEdX+8wRb+
/gQXu3PAJ722pLXgdO7vEeCl405ATEpDQB66DducqAmmXy5hqnwLm7tk4JAbZcIz
m3kqv8lP4BRiKB58Okw5r+cJH50wGZSsP2izc2R8TBm/4bKhScUqc7GRgs/sW6qZ
haSK5URY6QnYiPba+LYfLmg1/uc+djMahVivn1MwlX6EwE834m6J5kTXxJS3W4iy
flwa7/isSH6gPwaT6VNcjFubS8zmdQFjnFjtDkPDwWDEJ/YnAMJzMT2bbVm0cUwc
kSfDL1c9DbOnuAj6XmwnmECSk3t1x27IcN/a2qhI3XAFY4Dr6LbvnHqIIkjaARMV
l/X+0/MdOKa+8ZqcTH0XIweqMOyhURQaemEbsfYlbZR56J2AXkIhmjna+lXUkOOr
MdKzn1ydSCgFQ16LuVcTdp0LzJbUPGavZmfL+AhtDgLkNtCpSWbeRvIVxYC+4snS
F6i17bovoInZzITX0o5rVGYAt/joXF+LBr2bU2xhgnxz4G4Z436EFp+Njac3tpVY
XtY/OQK4V85+/9M6H+2cjlPOMys9pQNq3aY4iZ2L8PmpzqtTrKGEG7LninwPPiP2
a/yTfqETu+hKosYJZnOWUmfI+D4nhdzFo/EwdICrnpIRC8zh61SHlsOA7+YQLIY3
EsXuP+lb4dGlK/broS3Mn19nT0utt4u5jFiQU+/CUFlqCMmHP3/Vku1rN67NSlXR
PcHeqUXdkwb0d1TyAcBJjTX5V8xekbj1HD9XtW6oSCVzJbvgSd85hj3nsNmiAwME
ddQDSYUySso4ku21JTvAeeICtQr4ZaOKgn6jsOBVp+H5bVy/wg2agP/l6stgYgCx
osG2XuwPkRHlVdyt68eL1/hb9tmYE8+4HH8EqrOinXmFMscsIwdiVyl/IZY0a4Wi
nMRWyfLa+kBgQ3BXMgMqNMaTMsHa7vFzVattFdxRNTYFIpA+gaGwe7p8tCJjyuWB
WkJc8tkvcY8DfsVZU71/g3M0SS9Aiedx4uGiXRrsaflkSYBhMk6uUwnLAilbphCD
LnwKbO1DT8mdaE09p514Hhwyr4LDQ7EP1ozVvipKE+KHS4dONJSJznxm6rFS/Aui
gTJxPfMgKuolVPZiYVXx5O5Khq7e2QDa2nkm+i42dymwbqx1+J812bQEP5yVpKj0
XXBhk2QGMv/mU1tFhPObDjUhgARQrgpmkCHgkM93ASNHMrKkq7b5RgHmIjsi8vxG
PpBMsNs7wI0eRb79hKikI7L2JgWbKYRVShAGa538sofGWzC2aeuzWIwLaKNtYfn9
/jiOgcwJVTm895SExXL/4QEEjSh+K8Knm93eVuZ1mzVIeemwPanh05phq57tuS6N
C289l2oF0X21AZCawRnM6he2j6+smzIVYO2rrebrcOuS5Rh3ispMW/EK87Vv069i
wDaps1tywQ7dzvS+LVM/3uGgBbOyAnpu5hFNGno+fGx8lmpX6GNc2djlr5algb//
Kid7zL57ytioKr8wh8SGdmDZj0GJnyNtjJ047R7BpQ3kJJjsVcTqy8m0KkuBWpRv
Vb18lZWmvjxiK7+do6sfuQwbfwS+OP0tJq0Pp8UofMgoxlzv6XFNAoXN8xdjQxUg
CoDTWuhD9xIw3hX2G9NxRIY4D0NHLI6/RAP6hr24MkZGBgJaBL7voL5UsP7Ewwp+
j2p9Euh23B0iszxA80mRf0j+Q9JG2X6L6jeaqtMNEK0lC8QdLLjwzj+maBaLWKG7
25P4CXL8TFgPMui2kNWFXM06E26KehPYco81IeUzB4MwmnXUabH4pF6wvrRlCoA9
WUIFXyQQL85X9cJUmm917AoRJYEMNpn13CMnmJLC2+QipstvEkUgk4hP233WTw+k
uZiyt/TJCLPxOS6axu/3aW+cfd9S21Wk6m75dp7kL7mpJgQ+i3liCKOondipaD0G
zcsamk1TtMh3ZkSd6tFKYlPv8Yz6Gzvcf/NkxjO1TibTIzeKymWq6lSrBxlNfhy/
3tdMSyRgFd/X7sYpDtIB5OOsEP+Hw7lZhFe5j0ABZjI3z6m2vhFhn93fqOQD5Yb9
V095y6iMKTYFYnTxC/zjRuUr80HpupYpAXC5cs+tNBANZUsxAkMZqieGi6bjk2jb
cINDlXYkdeJPlrI4jdNBVWUeRqxUcMK/Hgc8AKR/Srlqk2rHSAYdzjH8Ptj8RdI4
sRF57Um/+J0sXprt+ANYGD8CWTd5jdCKQXWR5+uj3xtVPLWgnzCPNn6UuZjGmv5e
FtNMi+ro0woVgO0SptDi8H/om+1b/XXfiXIBmQKhDP/iBKS89EkXXxolS0+EuWZ1
YeSfhqbO+4TXw7MZmIDGZzUrwBmsQZvWh4OwuOWJdPbwqic9TbBfGO9nLP5lgeik
kemC6GS0Epy7qRTXd3IHapYO9X8T8VA237AdtkRi43o9mRcLCLPx1XHstx3aVlXi
o1mqQFbrFpXEvjsi8u85ZupCTolwArGj1k4ifP2HPxZFJCLmvHAj99vsKyqf95AO
EXEoGDR1n0OmbtBli3wdPYW8+thd10bu3koFP84afuAjNX4gkACK4GGCiYmxvXjx
b/yUEm8FErVH05qQ2mLHpscnAGmWfMJnNMCUp65ABqwdtw+XWxFjp5MtdoGfGtBn
u5KXtjmX+yt1VfD/IVYpJZNbu5URdzuxkXAovXyGHNiZ0Yds6jWpgtO8Yt2JVNoE
QEI8p28KXKbyjcJA3C6sI8JW8XvuCl1dHh+OcZbPS778535B68E12wcmE1FYSwNb
q0hWeN9CZCs1m98SmjH0tSXPs/eEaev3zfumQPvQm6U32mHvCHqYJS+V7ZBra1sj
lf+bCjRSfRPOTH6Kx/Kbep2vjSP4YspwjlVv5mh9/YeVBTINV+L73Lu9DRSipphE
kI9/Mr85CPQK4eHSGncs15G06T/hE77Zcwwr2gBTjETp+oU1filgC23pHVzcitjO
ELMi0PaBOoUHN1BfB96ubkqESOccVow+kIDkEO8osWJP7cqFgPogEGxdWhb2vsma
Jfoq3ENZGgEveSXvcEX3Q0keXwdSl5S6i+r8iRibK9oLm6Vm0qDiLEutIf6FtJge
0J1Bn1B2mYR1KE0AZynHKGfOfndj6+5HzG4UTvm7ldcqj2+HaObbKgOvDAjdMPfy
oxsD91SVA5vWD+DXZ9ZfX4S9oEod8MrZQ48XtsPtHa4qZgqsS7IBGN1E9jh9m9XB
qf7oP1NIWCJSB/OkUmYMgNAp6MwTGhn5MBQ1ZwcB6+kNZ8/qORplYrzhLLw0ghsg
0SaYODkvN6ut85AGNqBhRdBjbCXl+mc/Gm+epGS7vb2bfmP95QZLvldMl3KVzXT+
FcPhcVTV9t8Je1wvUsR7fk3/XGU9THiA5IjcTSAtLkZjq0QWug4+ecSABECqLoAt
LAn91vqhqSMgdqbHQQhRrwa3OG6Hkc5VLKAH+aHaP5q5MkksG7mokGN3Hx/5rLZP
eQvJHZevXaNFNwLL/woA0s6r8YDVosoHSUIFX1WKyipUhhAoxiJy9n+AH040tdWA
iuhh7teAcae1BWxTusOxmDEnezF60f05PUv66m4sOVoEtQZBTiw5jsNxi9j38Tll
+ccjt4jJ8Xx6QG2QDIBf5jA/p4lEEiTRwt1VDYmndrQPlaKsuIIzyL+N5a+3Icsw
N41lE4FbmaCa+I4NjNZu6pQaccpyT2CzEb5xoE41OEcN+WJFBp+DQa7obsCk2tK9
s2bwbOh4JjpZpYl5sn7VP1iF1sZYV5Y1Ldtd2ou9ziNc0XU/5LAKa1EAulm6zITp
SpV//mCDPzq7mJraLxWtpJUlXuPwzMXMVGQEfrIDwcLidAwr2V4Ke7fehHmrZC6W
OwakH5KJQyYWmaF8gQiwpwKrvzJr6zlU1cvix48KyJu2D1lK2dEXqfKEkJ7Oa06v
8OshVK5A2A/XT44a7ST+hC5rNLxDOdFsIsxcwOakmWGqF+ZPzfa6eEEj+VMHOphE
gjFRJGQ5LTuNGSWXdiAfkHJ9XJaW5+AK66BaDPsgtyccHI/dcbOSRQOmlfN28BwA
QPIY5AKhc7XVztKT381jZM8UdcWaG34q11foqC5VVfpHA39d2SU2RSc5THVeS0Kc
DuBz/h3c59aXWdyPoHPxtmUnlaltDxsbhKWU8iBnVAYfgoYCJzyzDUi0blLpv4tD
rnyeFMDTdi3K5E3MMUDAl+dONkZK0MnmVQkDXTkjiEkpJhbbGTzWxIdE7wpBPv8M
DVezqE68UmN0kj1P3aEh+VwzvJ5gs4NheZor5TjbjHAcngOSxk6dSW9D/K3KgUG9
mTbYhhOeGXcNwfZgc0IcphzILldVXcAfQtye4DXdkYXQnmRsfRFDf5pKNQIhk/aK
pVUO46TXq8wHwDxLNTN70xE5Cw0NhqHtyv2bVv+j3MIia1UdqNsePdN+FizMcrwe
53d/+9Gjjq2K+NtTbt8cxgWFx/nfk/775NXNs7by8LsfQ/to3fLcKKNj5ulEf6oE
EGloHXYOjHSJ9f8mQLf5cYI/uIMlgKFy2cghiP/prOmnapRY0oZ4sWXdp43zNfU/
BjCti/K4gXsIENTUtgXkFSCJo6HyoQlWMWGHs0BHkJ+jheRmOql/15bDz5f5ghNA
mGHiiKekbVryDe8iEX2iMwqFCHGsvZXaZAkGGWCqcoStJdJfY1s3qZWTKkCy6luM
GhTb4NF7dI5HvYQMq7CYfDTu8FH6W3ZzZZWZbAocPiFqpQiaxIybKaPm99chRzLW
HCOKuumsbM3E1mHUm35r7NPCqnGmcclNiwkNvIMANepz7x97f/C3hSHg29K8+VNj
JxVYj0p13PdCqx2GiS9uCRIBvQMeV7Ct4JWHx32XNPvyVA9MMVxzc+biAe5Cw6ob
H70ncQyxfJOjD05Ateb8qK8tGOUXFF2NyHKaOV7slrSAKYRyPpmhG98pyNCTNcJ8
Ca9c0DzEn7WIFpBrdJp+RqMce9o65wKSoNaUIWqUvEx9LyKu63ZYYXCqIuccIHR/
1qLp2X6uT9qPhOyvKQL83Sr8MDb7aypqw71EyHmbaiqNQ+4MOpVyD1wMHHFTHayX
RVRIHrTGvwjkFSw+O2R0gf66qw5cgYJ5lizasgHewM3GGh+DvJswa9lcqJtHeEBR
L0U50GrfALxrbJxJlE+jPYO82DigZrMfCFnIJYWRRfPJuIZBsfBRDmZ/IjKSia/K
W3VChLlNz2jKftoBZb3Hc/KA6iZe3sFtL/KPv+W7mppZwv59qwqGkGZkgqraiMnk
DQN0EZL7m8sxG2QQ3Pkj8uDA1uvbv7taPDSuAySBFbbTNhdBfqLLLcR6LQTtpYkF
AGX6qQbJMSaYzboso5rwpQ1Y1HSLQkyb7EP+V+ymqJsUt9WraeMH21Ge4EpHqTIe
Krx0+iX8pdIfznJPxLkVQWtBfUelOOlk6MmpT57Rj3A2zFbuQIkl4gg+O5KVvzoe
FT6DlIfKNrV1Ge2y3pGFxnhcxFT/kGiHpmMHFHrwnhrZz1TCi+AjqNq43Anq8zxy
+U/fh4JlRTVDPLYwngJPZ5CW7Ng46oyeI9106xCIwpTtWu7URV065JWqL6ES1x9P
Z891/9xiV0WEu0l7/kL7Fep3D9Emouz0Ag/RHN+cqoEK2s6qXsnAKQSbWSd1ABPv
OBd51OjS1N3Mn7FyjZoq1OKp1ctz2ryGubLWPaeNwuxc6AKAjGFGC/FpNcP0bSS1
EEIc4dGk8lxCVVfdWCIrWdNuT0OlZxU4sMarmmsmhPdLqp7dY9Ez5GXQsTsbLPzp
1jNoBW95D+6BJv9XB9v7qwAh81dAjun4F5jhMop6PdQiKyx4IlvEvueKAdISZTla
LaBM+Yuuf075d37yoPUguiqQHhT8YErI8bcqSVi5RtBWxzftjfMe4d7up0txjTHb
hTH0zu2Ar11vuljOdYV5b/4J/6vIJpyhi7riDAfPmchBcaGZquprTRyby6ml6JMQ
C+ogVj3LIGgelFXauVlRJXBlmqk481/r7neN2nikF1ogoPjlSnO0Dshf/mOhLSd1
P/k8zydAfyQUpM/seVtPcIHjJpSwzsw7WR9te+k8Ns2yEyF8kwh7Ghnd56bVABqc
vOf5FB9FYCr5R+D6WgxnxdkadI1Jncuca9JSHeWVkqamIC0yP74WjfIhQ9HARANQ
ptYm93Wg8L2mtYfIExI9G8u9ZUHgIj4yDXpHvUWCkE0SmkNqwCLTLYjkc+0R5mTB
HLRHM30yG/Ppu+KF6aF5rgb3Pwth2PZNRNV7hpDgTyhk7P+j2LHo+Ac+iFSgFOW1
+8yoyQ0uP9Hl87pMTk4N4DCb16yoPlVl4+czLRF7kCjT5bmsm8YhqOe5Unkuuqey
HQ/J6X/F7qDarSKwGcQgHDgxHW+5lZMSQaCtinsSjEr3g46vtjLEPSDzfA9nkh4v
Ogde69AH1cmuWoc8jqaghHFBQHOE5x+ZxrSfAeddLITfqo4y6MX7BLmFdfKcisNZ
BXPpOavbyB5J7p/2d6z0tTR05GhBRkC8Pnzw+HbJsuyHUH59dbWiVzpzVbvslerz
AvYB7cxP+erjvx1fR2+9Yso4ibvruxNoGnZh8o2x2Fm8jjQiHuNDGJWKHk7AZGie
1OPeBR2HGzHORiflekzYR3leHgC5qAdiXlfS4Nx3znaXXoXsM2cZNNO4XRtEkO2J
uBmzn1WViPmx9qtvPzLP3BLa4PJHgo/jBhaTz/WFg5D49XniM7/4khjiQL5Kt1x7
s7JUOV8/DlYU+Ne1ufk5JlsIUGn6ll/f0cLiXGC3EBB3v+LbO1xw5/JLIr7hJCyU
W/x00rOj9njeJggSPofR1fdu1X1kLx77tkTCWNF6mvPIRJ/ZhNyERvAXw40AP9iZ
h1j9wbIvUvjAcPmJbYlGV+++tpsVygL4bwXVNPObBRxRgFim/UaSRjEuGJZccGyG
mCX9lK9BNUDI7VKbVcO+3T1vvpDxhRAd+hIBw0IaSrErBdv4gYr4gFp/OG0CmA7s
SXszddb4qcy6iEhIyYue10BVnHSnJwp1bPPne7c3A9k6t9/hF6kIJhYrwCyk7lzQ
Kdk8fj0xl8Ky7ZBP4EBn9J9r4GmrSnptgh7mUt0A4VUAaeoIDFfIfhdr2GKcsgqT
Fg31fBw8jRhZnfVcFmqnaao9PZY2rYrJ9VggmvznbgOcz+auMVo+eaLJ4IwxJS3/
vMepn4M3GbeqgsSmQ+wnYdJWtzI4TUf/K3dADRT2PKLTLWuoxDdMJ5jwkOd3YQoT
rDQljpRpz8IhMULMHt+xvDHAnUs6vAtCuMfy55P5j5E0sxm150H4g+n6I/CEA5uB
zpxUom9NVwcGseZoDhdf55TfI1YVqfe4GSf+bkzDrPPBsjDKiOc6Vr9BQcDPLN2/
yLaThpR5heCQfli8hz4SbETApAS90cbvfztxSBrUTC1a2+DbfivHq+q9wNPgk2Wx
n5lTcn6kedXxMWnsmHF0W8HBU97h7sK4v96TFbeU3rQe3kWYj/ih4ghpJXvunF/6
PpjsVmNsGEVOWLbyHwc7F2Gon9jy9i7MLGPHQQG/zbn3ahYC2Or8IQErppdtRFZm
3fo2SuDOvVsd3H3PR4FFKfpismCe3EFeFi6JQXX3922qiF3tYuUZLByRwnB2a5Rn
ciNjJOuBs5eZF80PLuZp1Wv2SXd5J10QUx7rjr6wqYrWt1s1u2IvkBIdsaSp8jEL
tXAO4Qu0QdyWY3JKeGOPi3hffivk2HOFpRxGMQ4824PsH/j2Lywho0X51iRgaycc
KLh377rfXG85scyIU6tUPvHi0lWdfRqnJ3XPaqRgeyoxM6L2IwsO6K+FDHb76WvY
h4/bc+x4AYWsg9fUOQ0CDc2dUYwPv1xKH4GPBYdAKe4A8y+H3X4Scxw9L17RQ8vJ
m4pa7a8tinf9DKwjPUQned1bAVbMNtmK+kwvn1i9h7LoMgizGAvrOu3adS8W4VcK
R0fVN1PCU7+NzsQW/CeiJTdccWuzZN7LB9ZsGWPmXoJCGo42RbRKOUTCAJkXXUXr
+sh+g3WbQYOht0VwP4+fQn+Bx8LVDskOr2Kw1FxyiCSp1NsnO4aWpIjT73jC2dAf
5HtlABniqarrEl3SrXxKlYZokhIllHS4LlABo1uMV3PWkFIiiTTZ96PbV1DWxhe3
ruoJZaPuilvX3OuH3Z8mE6HSV4qiFjF1BBIj1v6lNINSjOsGAJ7Y9+67XYP47sBn
KYzR0QLUrAXRUlVM3mABnaMOjLjr5/a3vWKQHMjWvYNlQSwYHEfuWTP9+l+p3Lyr
P+MFJeAQk0BE36U3jCR6v3Yeo3/J97/snvvB2TN6CjeunW1sDzFEgCKZW+X0zI2g
9ECKdOcUK/Hd0Q35jpGPtix6r4cDicRcVwKEQLSXkEiLO9tsOLXM6mEjHEJ+pU63
abu/uLWUxQyUp8DkofFzOLMdNnFivPZVTXL6y0oCnL3FQhKZKX7oEJnB8jBDch7q
uZ1Z0LhG1Gv7u3nuqtHMUxb6BaL1ZcOlFJo4hF9dGQz2W81jiJke+IIkEb/X7Lnp
BLhtraBU+RMFeoZ3uN1wVddbFKXEzUSUg7ZTX+MUO2c4Fqq9TAt6BbLowKZ33JbL
AkO+9XA4WjO939Jgji61ZhWp/AYaBB7o2EKwraCX6LyqM5fPLg/n44uWeZ5aZwKs
+YzNs7Y2AOGBrTOrDHpRyIztMVeJj1oDR4UZXzh8Y9gfsumH4P+xFAbH9m7CvaLb
ssfbv/A16lbAq+7nC92DFtRJ5AEfBLAdqFEF43/0+qlH0ffWyYLxENa451TVQ7Gr
TGNd1ts5AA7gBiYcmL/zYs5m3+rfSuG1ezRTjBbCuLcrH1xA+/mIa9iLPzsA9SlW
tO/uZnQeOSX/trrX7OQqqY5wdIuy84jgM5H2fP2Q0M1EmBa6JeSJGpJn9ZHoGJRu
EF+SrnZ9icYXRcLyh85w7VpAS9L38gMfZIa6I9Qu28C7vnhYQ5cR3WD7amUrPxgv
cDFO/Enj08N08GsopVb0RRvdfeqQPdOr0Jq4mm3E7eV8mZV40ekiLIRuKgy30PXk
95k7/Oy4+JEKWeZrSI5JLXtu3KjV7Wp0jG73T0jm+AU0oNHBF3qs2IIjO1R/FmI5
nJli5txG5mjCdi4epPzxF630itAyIvBq3VRryr6e8lCnsRpf2FNwHxoRxvxd1+dk
MG2ewZaR7qklv5LsXS260TawDTmYs/2SyaGNYduBZp4XP3GO6axas8NSmM3/mUXG
hOut20FCQGM3V0HH0vRsNgq2XkEM0r8SFr/f8/TGGNqF5KjCN7pUpdhvn5MoFbST
Ko3EfgQdGM3c01/BYPcbGKxBsJzFo/H+KkxBwvlWB1j9jTZshUdlU0kHWxK6xOV3
jq0hAIUJKO2YHgljJCodAloh7Mm2l7dLBfRcn3rTWPTp93qdEIbZfqbBF3ADQiAa
qPS4/jJJS5iw99rb/xjcDcMaKLlerADjWYrPyvNklldlXjPRG5wpuFMsfiINe6RW
JGSXvz3HXrW84VbIvAQvqjH9gPAzepB5KA/J+ITTLXPUeWGY991eJmJspJF0eaAL
/kh+TnwQxX2yIuCXC+w2rpDrieRnRtwGfcu74AVKY5gKx7Y4sEGrVqxLiVcbxElB
NH5HzbduSbeGwShycYq7cqfXv5gMLZ7ucPasARZYceQ2O3Tc6fBUokdnvz1YBEtf
gj77wWU/7jkHmm4kYQ1288D6sOROSUgpbqERu/lW2tormuy0fwn257w9cnCbBcVk
6JAiotphiArzxHMCYKTL0Vv0yD9+ptzEet2O7bTxzDvFdipGSjg0WFE5by3nETco
gYw24bHxHWAuV5CUX8x4LpJItxmKCImgtFO0YRXXyEodHguWz9Sr6BgouHSVkiz0
4clj5WVSflqVgx4C8T4RxqEkuuHrp4naV7b0a8VZwT054Rtdo87FxFjvkBxXKHZb
ZHhLFJDkFQX0rPFf9E9K3DZS1Wvuur6ZpGhfhwRdpsXYlgGkTcf2hdY2rzNJYNtQ
y1aRyzKgqSi8wGuhLvQE5hZYImTTlUh5P1v5qwFjCa+lSBputCsNqSqYk36nJujz
38nQkWBODxAMIUocuMTOQJMqSjMxapyPGsHIaORVuZ2dxHfC3oNMLQC30QdXJrjb
tG76qiXx3yV2LFOdzW+rVgqO4QltCtjzdXFF1KAqCadh7VcEeyzscTjtMewGiKDQ
5immkPmmGg9ksEwBYvmNHL2zL78De6SbWnO1Uk0/F7R+qkkysYye6530jMrnw+em
w4pk8QUPaON249RCVyTTDJnnpCGZ3rH2lSeHnbZ4gjxs1ZD2T2k//Iy45TKiwih1
6OybxXTRhHQom1p0iLYQ1fl/3Hz2bnuJYX8kV7CwKZ3mUt8X1aAr9VPWcz/tdjde
3+0bHUhPw048pa4SSE1sMiP/AF/LlVbK7PAEsGb4vjXjQ7uCgckWStM1yEWnb5xS
47pSxGQK2hTYl4beCqNwiUsbkVTw5RHRwhDoD+Fon0Bk5js33wegJSz3NmjxgMnA
dzzaCQH1zeHn+vwDoYO/xixq0f2bbtoAOkDEuC3na2UxqynRDJQbIqPLibM1/HUi
w0pYIspAldlmFcy9jvkm4GAjr9jZ9k0j0RoTH46E5J5rl6gF/DdFqfaKMnO1hWwM
BxvC/T0g9iQIVCeqdF9lQrDir5vGN2BStJxrVcB5UUuUq8PkhHvZNCcTFKoxEIs7
kZ8C2UkjYmX3+snIOtfUVCi7jY7/oLoSH+pj22SHgFVuCdoG0zSoOxAcPX9TN2aY
LcdK3y8GLQcdU4llO7VSROtf9okIHjdYhKbp+O9Ym0RvabwUcQGScjSLdKVJeqYl
sMI6tse81lC+964h/gIHUrcSMnaZE12CctCYtO9g3kLrWkomB7Nb+8fCK1DdDBPx
/53W7X3qVJDNuBIuTKmDddvf7eor0S1tSKvRMmzXNUJ0q6kQwjJ3iXmg38P5xz1w
uToRLClPg4kzxeDPADuo6DhsHThCrU5y6+6/vropUi2nOSPxH8zFSGRaTI386WuC
4yjTRcv7y8rn6eeoggfmEbVHcilE3DL4DK24E45KDZjFx3Toiq5cTyBwqQGWHIpO
tolavOKgpMvGH2DTPjLWfz0IUFnUfo3n+BJ2SbouW0ehxYrTl5hwirQt2pliMmlX
xP1vBXAXw2jvzJZLwoRC9WyNMLNeWQkL2WdRDvQpCIoJ0Ec06/Q8VDd5yf2ziYN+
qZbOihYNG3DxkKVQmV18wZYvTsyD1A0ySV0ofbgalAslmyCVrAH2y8Z44wlwSpx4
pItvWc+adVHP0dXekotD//YNrU83xfa04KeUKPdgARIEkkfUN/tZlH3AHhi/sNxM
bV3q8oHdO3nhN96cnmnLrZVCpifR2QeDugkM5BLrTA6qJz8R+ZvOPWhKhDzzUjoe
R+8mY+cF3VAH3xxY3dAhKU1X6QLPsm4GV8gdicz+rFUoaIjaORj28PZLoZvPcNaA
6xPvt+/bq/NzwxfX+BtHvH/eJQLnhAflVvFhaHc/d/7PG50wJQ+UV/8OF8tSaRYK
rgt7oyvUD5psUjBz3sbfM6wlmpU4T/Rop5NllLeygPwPsx1EFnuRgmNakyQrZ/hF
UGyEYUTjsOJ9GBYc0qVy0Wq7Q215DFwf/WGWyEtZDSDRU1MUBqpEjmRhqzRB7Mgt
6y48hfRPqsEXTN/Nfi8Esd6P8xMVHqymm3zUN7YaI8+8/G+v8mswL4T7y2m/vqxL
qhQazzg3OVSmQHk7wgMAyB3rUF16J1sCAmhDSp2B7Git5Ry6B+19qQBCzXFzGYVC
uHi5wwHb7BUvtoZpqn5FSKelgvH56U47lBORT1CS4yHhoeVOTO7DjEPwhYZGI6d3
PbzSBE2iV2NyA9IDdyyeqeqv7ZRnAnD/npEC+tllMzWKRd0EZpqoZsFD005HRp70
PscwRHol+Oc98Y++hglDnw30DcBt2CYIO7UisQPNKQKMvUcXbdkw4IxRc1mGrcj5
+fZdC1YgjJd/p35dO+24LCSRBOsKo5Hd0qj0FK+GiqfI2F6kfZYyxglx/wcLMAnW
9ChLfN4H9KZXDFTiuPZzSh43X7M7P6npfxbYN36j3F3pjeEQf2wjtRHXGzqVOzMR
Jtr7IzmG7bTNiDygpwdWiUA/BiM3a8gDTFrHPRRBHpWQYdcdBcX4XJ6RY1ANtDBg
+eS3vZXJ87cj4rMv3fIqTHfjx1D0FgJWRMsMrJ1sSCeDVvYrqHsaRdlSGiYKMxLp
mpU7nGFFg8BokaiWn/uNgz7VSDZrR3mEZWLlVvNYKD0w1pPWR+Lkq5D6Sk7zQHum
rylYVFADwjg+9rsLObKCm6hcKMhFmMMDJeyaR/DNq8H9KmZfkRz2lW+40r3bLJhC
kqB5mUcGEFnIQ6T2rQ32RPapMPzuSvULGBqvXClV2eEpCLzdgF4XgATDg+DMf4Lj
N36enSCX2tVpXvh2/QZ4sgXZoxbnACtDSzMNYyF9iM9xRq5r1MWXfiva/xb8Eda5
d33G2OXEmduW+mBo81+3CaPbiht6aQ9PbC6y4nCqmnCiClOl9W+xpj5qZSs8IvPV
0n1NvSFoojNNQM3EpsgoYihOE9h7Q9Xj5D6J8gG5T1oVaKkVlmeQNbca6e4jospQ
/LDkrN88UBY8IE+h6Twk7JjbG3MHbxQw01v9BQ7aKeiEzVMvY4Mkh2rgp0uEY8tu
l+JIZFl4qL+5P7ODfLuXrrRvft4sEbgaoybdA1oipSYl4UUdK57GKj1DxPvv9sbr
EDvKMGOSPggJ1r0Poij5xB075uqyaUgXjI4lZgu22fJ0qaUjemc2EmCHlvLjQimP
Kv4+f01DL1k5mByz9CEXNFKJ90QqXGT2jX6dmADQHGRR0674MYx3xGeZ39q3x0IT
o93QpBZTq91ico5XH6dzo2eCHjgl+V7S8kQu3Lr2/7cz71rp7rI/olOTFD0t1sT8
yrpw8zFY4GUA36OU3ADgWJq59VNUwJE9gDRSWh6t1mflgnL9qnMFP5ETcTVbWoEq
9BPMsbd10DOWzPtl3bSkA3M/CrOvLzvOOwQ1h/PXCTD4zyxOcxZHL7KTpoO4eLau
gxMsfBCnt9rpx9CM2Nc1eV0nCeiobJ3vbKURo5pRYu0ffcD9jVuAxg44HP9P7Z7N
8Yav41r1Mswp5GHuyOHG9XQSVhqJGc1+8EzSZaO4LOPFRAapuJkZxE8HwYeyK84W
8C2Rgc877L3oiP2Td+GJMFcwdW/cXhoxTtt7vEtkf3jaHrYjn1iUpNx19UaxTXbo
imwJyFU9ORLQkr7RR3lIkuN/1cnxUL6nIle5nhJFtiD/fKfnW3MtgzEd8LHL8tKd
y+iy++20SRx2tmMpBz3jnwuJXpbEegW+v/uo4KUQwMsO40X9qjzio4SpsrJt2Rmo
sV1+Ck+OXVpj76IOwgZVcpERXqoo5iyZRlt6GNJg8dvthbJ/MB3k1Kzt9Qe9R3bV
YR0Kv06TRLuCzmwcA8WvBo54/t630H4d6a1ewfKMMYmQ6PqqXxePEBMqw23H5GDw
DdNgxjzZdnJquK6ap67EDR+tU6qUn8c4vufAD0QPLrxAoNg8WM+EGlGlrLlWKqd8
SWs/qLMBtASUMxO5BPa86Vme9IGCUNk2ADqNsWTnUMp1hu4M5I/JUMIzX33X84iX
OV57qlxXsH3Byme/b/oibP8aM4NPav4gQtUq93embqX66zJlI4J+Dvfq3IJHkOcl
0L9YQtxX6hwsn8NTWViWw5VliZZ+gEv404/AFhIEe9pBcDUWUkg5KajuefWxeO3h
ohITP67r8xti3czjUvjZpbLUrbYTb32BKThwSSiR1cJ3FfjwQV1ewGsJQfZmsSgU
R50MDkYTb/tZ4ibsrAbQJWb9DwYS9Kq6f512i/v62IXD+RktQICmqOGCZ88msGYn
AvfTbFwDBt26cIzcmS1R7q23Lo3aZIlJ0YXwJpKd7arLEdescN+AO4bCWhf8/piX
GaY3krkF2DFFRM6xSLoN63fGzSsns7fqGkhd2M88oOvFP183QW4kSwjWNtGXn9YU
PhPzHhbxVjggA8/c+zkhdGmuJoKeeRssgn+/7zBhw7xTZKaYYoGuzOSVqkyYXrUJ
F2E1cTdWxi8C0yOyOR2HnNr+8dOj2IO6dvGRlBpd6Ubf7ZmqAKzclGi+Yon2flMO
8EXqD6ucwg7SEamSTcihS6dMmlhMMl46FZtAunamomHCELia9cMrMsuyksbyru+I
I96tgXaJ0lHyL0oVe3hu3cMJnwA1UEuSvwu+lBJPrXZUW4ju2f4kIWB1OzkdKmJe
M4OgysnrCtaUCgiQ5BuCanN/kryx6kx2oHDmAct1Y4rWAZnJVSa25kgqc5C3f7Wc
xjwHL2Ie55Wxso5Kd5Ik8/1UtnoazB0cRRC62yRfKRwbolzpRHilEuuAEeAJUbUm
y/oYEr+mrX8kaCLBN9/hMsdqCctbEIN077xsVEkg+HWxxwWmhM8B784GCuQsB690
A2HBK41r/6qyssYT0FTQkNEvQJ2wkeZ8iNw6lTR65GaBLdNeKPWEio0/ISCgndw9
+Edo9VQQCJF3N6GXuO1ElThjAllGh/neK9VBZO6W4oMxo8EuJosSZ3fle8AzZ0Hb
iZhPTRtkujQVzu4Hu1FnOmvLoj00vXk9BVP4rlArJvuz9bDKsOd8bTGvp9kKMu41
DZRPVoUf45zTCU2lTpfm+py30nj6v6gISEl+SeA3LVhc2Xa4KfBbwvyKlvS7gs9M
OVt+KHAT9SYHXeH+KqscimHWkJEX7FpsNHCjspmESbOxnip0mllz/+3vYIwhlH9p
c1qgZWPxg6fFV0Pk4ftqqinNLY47PXd4uRm/++iB8IheXW+CtHZ7BPdk2b6YVrqe
xPhVNpQ6x9eiypIf4HfHr98nUvVYy55bgIhMtQQATKWTXKbu0k9yNpC/XY8R7iFx
SOgvq4zJUy3jc6HjTC8oUoR+6SoTFgKMrxTFdVGCfyYwHTRMx2G19U6O8W2HArXo
k9zqWvPLmnNcBB4ib564MT0CI0QzMfRSGOC2BszQ7RZSBvZbLr24+9ZFFKO6BtVx
yZth6vZ8Ebt/KULBoYQsTAlxXEZJN9ZnT2J6hVOIgLouIghpt68CYtoCPxLq4yTI
4tM2YiQVtWxUfEmKXI3WVIF6U3ibX+QX6Ea+VuMP0e10DZACZRlR8KYAFWAW06mu
F5s3qX48qTBmTYRCbgJN/IFkblST2dE9mpX/3FBVb+BgnS5sOXs9ypwTwlolvUkh
pm5dRpx4A6RJ66VB5lo93K5ZHZUE6wUMi7OqdrJgpNYp1shtntBFZBw9fIVfNxta
tV3hRWDBwBN8qR5nRO36tsIPfWuhuQKK99/NhntuV4x+CPOXmma6vD7130p7+yMI
L1h5Dd3WMS2QNxKucuukaaQ4eSznUEqhpIC1RXM2vB3mIRPmId/7ECLdSv0YtI17
IeUU+z7PDVQcMSlqWayk8eGA+JRrugRwbJxycfUTVjEKZhXDJSFqyUw2amwTTYbn
3AGSmgKT1glUqsF8pY/CpBbBXaKA/3PUU/VyLFPs6uDcAuF3tsA3E3tflJeVEyd9
bsepj9jQQNU7SI2sIztu1vPEwL8scky6XxPK6kHiJFryMwg5LWdh1cHGpVqNr59+
iPjQLMj7KT5YDL6TF+2ZPkZEHSB6/RjVxAKn0bhGypnpzDR6LF4bkhI5aTgQ6uFG
be0WgUOwsE6iRvXqIAgRGVsgGfVSH00KzBDjvEGAiQfRmR8E4xnC07AVrtzp4XrK
Jzup7ididR09X+PQipCk8S5TaAFzM7IbUuaM+fVWOm0Ofg8tFDa1ySD+yvSo3Ij6
ucnLdOK6lBZSE5cpGR7dHrsWyoDya603ERVKS1VpRtvbH09JBlBmM45sSgWe0/AN
SMxm9yC6weYtun/2z+Z3UrmUfG6J3PzVeGkpUjGx1sD+Bt805lBdFR5503+fjgeS
FSog1u9g6OB6+i70/csIHjXuIflbHHCQbTPNzXg180afbGNzaINS89axSNtmnOdI
rex+4hU0tABncqIOSOs0nkWOUOq3GTtvDFrJbMjjIyACgCHbpwdQmCgnKt3zqw/S
V3iv/jUxslqn0Nt1PZzR3LNAOK9wtxrfw7e0lLVwwHihVX97HK1m3vYQHayU2Dd0
9f3xL0+No4Ya5t934eCx7YLY24CM1cEs3JtTyTeqiKEMihxTy9dC3TbdIw4LII3a
rxDJTzofPUS50A4evdHyRwTf9KzwzgSBHzibFyts53/npSiUMWOqG3qZEG8eadj8
HDaGTaxb99OoZP6lDfpVaMjPqp+m7bXiocizc/7fdaZFtYxW0CEwudPzIqP4HAPg
8KeilItfp7/GIwNzdcml9b0M6cMtYf0K1EQ9a83tnJCFWgWgy/73V3dE/KzS/C8n
+wR0xV8yAspLwk89ebvASjOyYh9w7jjuPQfL+6y1pD2mj2jX2yPWxvs/WwcGlE5F
C9AR03TTuIvmlMnC8GC5lfly+ePlUbOFPxNszdQdNuFFKUCad+Aod5Py7DZP26sq
x7Q+bJI7iz9ca2c+Uaec/MKZq9Ww2FteHUmQ0SzZZhp1BqFQFNtHWO3iz9J5VgrG
Hag3qPzzPvJp2NNGZ745Zxj6F62blk6VO3bADlusf3QNIjVRroyHG+pYAsdQyzxi
7hixjp32MDQ81FnyJThkmD9EQLHqvABDlEcXEYtUE/TYszemsK6rgRzSvE+wZlvc
+OTCMfRqYPT/E8/ggVitP+SnXj1YEhIheVRSmoc3I2SDxBwaqicqqhOrUbCcbgWw
GGRtYwLVWW5CcyfOj8Tj7V/2VTIlQQitzn6Ptha+sZtlcPzBUJosJQ0Gfvs6hf7+
4SYR4TQKtLdDRLOg8nLsCb+IXdqNBSDP9xiTvSgZWYLZQpXp3OncfB5wWLsvpITz
lqzPcn0ENMpMhPuyZGJC1alYmxhzgNdmfkeXdUpQ7d3sBkMtRbf70KjU1mwa8cW2
vlxOykpLNwxm1xpgAbCu8lWXnbL/jBGrmlhIfss6MdBmyPkpw4AF5ZBJa02osMbA
zNtMsokJj83V36IKYzbWpu85MBgvDTQ6c0J74if7np+vRtFvsDHvcp7BQ6r6JD17
KUay0UQmw3SLEBMe/TL7hXhDMgliGfD45cJA7VnjvwtWfQPlEsOsc5QNbynXUAlu
Nm+4mZUmLGLHz9ko+gqwIT1tN0oUUbqlF1K7TJYm/d5B6l58hq7Z+vnUyPgRWxnd
dp9YPk4AJj/5noA/PNYU/PozU7yz6R6Jc7XW/uUXMJCsX0OX+VmheyvkJnQQ4BCd
eNHOddW4nvVKh2xfz/y9z1vZcz4BhQDlbYVWSyjDxIoPm3LL75xtQG71m6ifZG/2
e9HbQ3Dqlq8So2pZiwUY6iut4qRC+6zjPsTaTczgRqJheWyE/4lG/QQMRYiJf0gb
/0EIdTMdU88ClcukN12BpbbUAE099/hc+RVMIY2q0U3gHg03mVDMa9tmHeyhu8am
Nq6Qz4HkETtWGfDiIYQ7o1SKDwuMt+O+9g7B0gC5aEbdatQwArrgfw38PjkSqZiQ
1RID+QTArU1tAggmMzXoo0SpsmBRgRncPFgdKd4wWaEFwXd7kl1V0VfITebSlU5U
lOMPPXEVl8FJgrNZhPDqbOaj9I7jG0RzXEFoH1NuFrl4Gwim04lrTi/YK94xI9eZ
m8qfkZMoIGh3aS2ciArfENwwe3QSbzD+5lYU4dEMx6qXo7cOt3OAfo58I3WMYEH+
jG2wEs2DmzqLW+u+9IatnfLbM1xoGwXKeWzmSyvvQG62DG0CitCZ9wiseHIRZTkW
KsnXt5R71NQ7nhjmWH8sbIu3lwKaYlM3hNNRomSXCIybdEmHFUftqc4smFCjeWZZ
mESE6xNaNo4ywTRoguSzUzkalrGInWF7J2Uge7BzqcRD1Ptn9wRLXoH40kASAfcn
jaZc32Z5IRqlBY36cr5LjqHF9NEaI2NTvGkSkj8MhgokYAIUWGg7O2hGgI7GLOuu
MLw93ND3pWw5ywTV1TomRlLAHb032HlF0ehn4r2oNgIsN0CkZ3Np+TiRy9wu+Hxy
LsUsZS1IR11ea47l1nCAmRUnGCdQJPiV20beIiGbB0LbyZ1hvQJGtDGrWAnXJWgF
A42j06QMZx05yk7NIMh+Vb6E463W/w9ubhixKoxMN6wUM23jUWyg2o1XhUXAvHRr
vIsH33bueGNpURReEoSgHPyWJVAu4kRVpFqT6o6VISU0vwgTiaXMTIqY5QnI3n1x
SxUnWjmi+mHihWEXO2mycPjJjTHxYMbFB1EOdhybAAm/IlET5ULr9q1fSlih+WV0
o79NhbfXENSudmnohHc9KfJouz0h+mnM9d57EpUTUeeoD3n/6lEwoUAwhzAWN+0I
i/xM+7lFE3UkFpg4uYUw7Dy+FBFOSu2mTCK8EdgQKzyHLwzwQmMRV2e+E9kpB3LQ
24cGU2/Kae+Nr/n32xFuKN18YDycBUZv2hkqsuUmHIkEY9bs92a0PP0uGSQhShWJ
+T2afuEAVUnkiMRcz7RAL+UWtcj9ecdfxOG1tQv0MckBMyj6J+p27USzOv9FlHeT
38RwsWswYrGRGn5VV3eKGfaFfYYPzFUr8U0gd2vVWsMM56O6QQDLndE6AH8in+by
dhGXjxTkXWjSVWOmylEJzjqe90OBjxrAIk8ywjZbpjhLiJn7eaUqMX8wJVNBrOHv
0Dn9xEIXKEi9dnNYoBP7s8LsCP3HoPFoF+oD02JXNH2xCI3K3W/ahIcLniHzBuyh
+ci5gfGe8JK1+0BZi9XsNNmG+/ClD2/Y+d73tsvOGo6adSUHOqj8iG4kJW/BwdUR
ciQcHTUXMH1sVLzhHocL52yaMRbIRE612GQaVtotI0hPrmJBK27Tim8zfatSwKaE
6rJUMLaRa+O6Nn3tbpFQp8ubEE+le6AB87wOUuI3wIYPqTQDrph03W70l3R379hQ
o+5tZUNZnXai3V6vPerML0ZBsHbUEO4Wv74cD4rtsJ6mhxxC9QFMTDDD2uiy4G86
1RyRwZC1mWjpRFEZ8WhXq46kOxxPVEFH0whm6iLSFavqQo/7M6Q8jGCkYaHYIEqT
B+8XYoUuNyYuGXB91EYgZjAM51dVkCIDnlLQ753zzURfBuWwrClxuJk4sW/h51go
YNEj+s4qjqahMM2BeWjOxO2kWafZN7sv7PZ7KwKT2+PM+b9ViA5QyrVQ5xa7rZFn
9EdULjvAhSw6te+qvsYLTfgQH8gLKqdIe/qaiExcYdyCqyhFYFIc+z96D2Btfh4A
GuHGU+Hv1f1gK7PT41pyBfJh596RhAQj6KI98k+YNFEhWo/KOayLtg8c0eb3zY11
2H5CQkeNR7+1hmW0M5kw3qx3jECmF0dbppYLXNPyLSU9CQ+Wlw7mcv5rTmLo+2gJ
FaHK4U8QSLWfW286lu/Pln7B7jeB6i6aiEOOlwjINCReEA7oacl0ySdlDekBkYqB
SyiTVr6rU130+AmEWCplpYjT3oDHlhc1qdDIoX5Hide2xzYkNhlyOEHxTcTGncSI
xwe3AHE/60cEY03zRaSMffcrT4MdGc7rcZvMNCO1zbQ4aPbUMwZuD0RKrBJMxi2f
55+WVuykzfFW4pHYEQesjbQSb3Tv3YWdO6CcojKd0Y908k9EGEdc4S+R0YfZcZqp
A6guecSwYGRhVAkF1SStysuZeCrVG7F3iFUwfVtpCMUCOgJ1lE17qB3p7qgUkITr
A62wNi2dKcXFLU+KH7lVpNnPrRmLjRntqFZR89O+CRGEfzER1+B10iN7WVFThp4e
IRWJQQeg3vhlzhjP1dTk9qbnBKiIdFKiy8jjgb2hUrhlkTG4SI/vMkcOSkYt8uu8
a491ZVMV/lHO5S9QC0h+s/rJ9s2WR3alqknSbLLTA5rUNCaZSEIN2mf9HZLj8tXl
JvzvlQLUb8KTZMYuk6qwrn4W2qbLvdy7s7YpZd/CL2oyVIRAN6OtkwTVxa+BeUXX
oY0S81fPeoaZ70/SYtEwDykUSCAr1EmmjpwoxwNQFfrO+ucY9xbAcoGjOsCuYCJ+
UWVGN+JUAQc/KnwNEZjOhmMV0+Q9i1rk6gXi9HG8vxsl28zeTH5uLflQ6IBdKPpP
znAeeEa+kTx1mBpCwLyhB1fw2cO61UDsd2dziLUx4NQ70N0SUmZDXCHFlLJQE13z
uhslCJdSEZ/lRu2/CPlaeC00RZljbjJexbiJK/OVoUu6wq3jaz+JFpIGyFqvZAky
xbUt47hZpy1qPl5BrxOo3HjmSvVYg2HNv7nibBY7EHtlzFXcR+IGPpoAnrAJ7l+O
lCHWPtVIJI6YXa/FLWjIEC81vGyH3bxVbi8zkDIUQKo/NCV4NF/MPCi7keLaDEZW
ISAFAQWioEOZPnBqwW5xZ7VgsfuyCm1wvChZg3jVYwUfSpn3hQB5XPMrfmmXCaWv
GZtH9/xeOT804jV15YIYHWqQv8E10X2NT3NWS83z12KDyFXAPKM7DBhsaCcjP3V+
H2N5N83yJG0QP7UPE/QDE3Fw07R95txpCTX4TWJ+jfM0hZavc7uyaoBRFffKzsfd
rMFVegDNhROqfoxlR8VO8RrAbcm+s4d0C9rggi8/Ue0REtsbjWY4wN7VVr9eD1en
x1NkWUY278n8NZ1nfDK3rWGIBhzbcxhLTY0eeGbQDrIC5iFMhfCm70XjuB1v0uCl
vpZLl2mHjcIdudkC6k62hYgmwH6jVoj12bvq/p8oGlNcgJrTQ3X+7bYBNUCmnzK4
ElXy1opVEQIaN/ezlC3oFYPCoaPb/UDD+rg8els5SlXIJCl1hZj1hzTgy8Il9aJr
Dkr+sF4mbf/lGmqow8PTMgsVZFM6rKpVmvJ0w8vn9sC2DzTxAc4JdzB7WS246aU/
nXdnCJCrp0bXZF9Oov9GCvbDNsGQUatLWrVj59/iYAfUVxo87EiUTFwpmFLx48b5
VosOMvs0RZA87NSZ3CnPS+ApZmHuBKBcna/0D4o2T4Iop8y24UWtxCrPbLJL7Jqi
a2WLEdRmrE7d/w/TQ8kPzW6yHo4YYuaN/o8RmP/ljpdC9R9QvXB6UC5Z7KHphdUf
51IW+76rg55TwsvNh0zF++Daxi7Da8T9ecLUohle+hWAK4bUikAKltbAzpFXu6fQ
Vre0jmgFL58gsidVqoqYir5R2jyymJKdKpok813qcERbhtlZRSJa319iYfg/sriF
TbXisKt6ZdNWQmb5jr8VfkY3Aarf73qUO770YJGz9BtE+Zs2N9dBACcxUs2/d5Qf
V9bUzfk+U9dV8i+MA6rCVQiZ7BLzI6YKzBi+IMUKrcLY1XrnWcA0VLaFMmGP+Jh7
3J2TRnAJjNr/gCwvpgA1XV4b9Tr29NUXBuNkaM/K7YeI4aXUsK8Bk+sboy56PqDo
RmJY7MEh2RQmhSvVYaLHY8YPnJRYJf3DjEmx0rzUEuTKbA+22M9F02Nd7uCId0F3
yHu/EmRDzovndOzA/TgJxZz6vY0R8OCRG1Hg2zwTaWVMkFVC9SjAiXC8t7jc89r6
cLhpd0qFcYBt0SdzqaIr81mEfKk9iGirflE7129QEG4pkZcpHDzl7v40PFfMbfwD
AgLvU1EbwBtKQp/7Jhx72/5vZxqND4sAq3aUPxd6zeWkIJYivzr4CJheld+wvrm0
iDjXt5yNZ+KaXYuGZHDcNbNFvw1x81OnJQN3Fr1P57gdKCEMmycwQdmtEjXLE4+2
/HJezWnnKDthWYJKjq+XYMxGKtj4JyXFitcVdgDNSsUqtDTjNzal+Veg5bzBFwOG
EV/Ou2IBVU610L+B+ukxvodvkNA3NmE5H8Q9vpq+3LuAHwABmLLaoeie9JSrEVyu
H31wHImMDVaVfxiT2W2dl0OmECwXM/TWxab4IhJWeI28iBddTfzNoKSNJTb1jfvv
65+lMAJLwgxi5ljDnUHUIRTKwBCd/3K3b0k8Wg9kZ52P98qym7GAZQCedWIEgYvm
DGCEzslT1yAOFXovrNzAg5ti9aX1sJMIQOKc/6UiMrAame8fv2OwLIl/gOuQ79gm
MkQLlxxKgOBrSsTSon1iWPdJfnSjPxu57z1TFoIRBAFrxuH7jGO0QFVPpMVAFQvN
16sWNsXzjMxtziY2lmnndFx3yFJ2xqYygjPjKszA+XJlhlXGDuPWOcmyPTW8y95u
M+/QqDopnuQ5meB9FspxXecwZaHV8lYs4u09s5U68X1Z2+eFdGWx8o9DMtdNkr4n
fIFs4s5eibUV3Pf98TaIrqYY6ynFPr+gcPFEFKz5OLEo+HC8zOeHPtlVwThrkNcK
hvl0HccARvP3pNtHtj2bI7dvNogfuyjeAhVq7ZMaxWWzGzx7LVbYGQJM19vjaPTK
k32y556QKzrJVe19EMVbwdxecklQ/gFYzO4kFlswz6aXeeJCdxUGj2fBnhztaAx7
fX634cHkdbz6m6W65HgdzwB4oFT0d1mI4MOAJsZA7/PLbg9lWiZ0ISOFs7OcrFsy
5uH+lfklx3xPQB/1o3voMhTa0JG1Z4BfcTDl86wt3Tm2TbHhyMafBt0JvFkxKrTR
hs3o9jhj18ZgnwON+mys16QZvUBpzZOfjOgowqhlqikA8kqSCzQKfyMoU90PyYRi
Tve0Dsb/a9xH6LBSJRPWb3yyyJrP9xyMr/5wLvpNJ0TIA4B7Q9rvwyRLZzJohcPZ
gCpKT8Z4177ZCXks3U7HLz90L9OQrYUQxRh5qrXuzsxwBy31Ip50W0/paXXaOu0f
bfgQBMSVtxluyiqyqoKHRCmnu/Kzwp0oGwIZfH+c0FrYaGjaEbgcRsNiY3ibrjAk
/QwoPEKW9hzUsqJLGH5/SaSVDE8E5wuRlu/bv2rKNkw9VWWwP0/O3EN1bfXO77xC
KkC2VoV56AjLB4x/G37bmFXxjgWsXFiU/hNKwWHx55f0kz8ItORD7Xceci1Lp/dO
pa+AoaR0ss9qC9++nbA1y5xPakEqAt1X3bsbfM0DEewSmifNlhGv9+J0kjPCO7uD
c1bvg9U2Bql5a5bldbQ0j3CrGxAAwZDr1+wCnzIMmT2OKLqMetM9YM4Ark7riWnz
47LXPqCrlgv+F0S5IWOAwvDmiypQC3I609sSQuaiI5JY09zFJaqyLINjl9mGrD+n
70Ted9xfGlTfB7THt75l1/+eMVdZklTxKLRNH9ltaridMiv25efWPuDKrU27GTJ0
z9HIZ6urgkJFHsrF6ef2ze4y4uvozoNg1iAaytm7tlsSSHdSt0lfs/lIw+Cp3hB5
2rh8TmqggiuoKT/3T4KSQWAAQJtU3u3x045aBlUc0efr99xSkfurVHQPHiZ9SHCJ
4BcLCqdDP6ipEEa9WvomQ4vbqaZYJ0/3Jr/LNWK2gWtWKkANFxtNFU9FTFaiuuaJ
HaPdryGUmCnDWHP7ZORhARFbODQ7iVPrN9WcniZ/UGQxLSYJtZGhDEn0u4ovSLSL
eVKUgfofQ94khhISBXloYSH4TkJDQgIBsxMUvNA/8vDp3IDThmHg3lMUrjg2qq+x
OB6ZPel6/rD3zZGibrNTfco0nlnyicMgGvqcWD/Griy8/wpJfdcUNQ6AQXuqMJbg
vtqZz7+jhjp58p+LKk9XRVVBtlOUz7oNT4+L8tf6wTxLJUJdDLqUxVz8M1bjz8AQ
6xgY1tvierrxlbcuV4Oy7Wj4QFgJ0TWVvy+UyiXZMs0zJnWdeeyF1j2E4Iq2/wXu
HujE6RueEV/fW70EXdoRT+PGq1QyDFnrIk3peRVVetbe8UzQ3TjILWMjZ2WrPX6t
hu5XKKhdsCl5WmJTwFpDiTbrGUD1T5DKURbPR3EBTitRlIyp0WYtvdEKJM8jhi9P
m9v57p+JHx67Yg5cHX3N3jMLFiTbV+QiMAmy2HvYsF3h4EwKv080uGD10k7zQksI
Pp9T0arPDtBb7uK5lPjkjkkiAB4zddba9XBhPQeoxzj0kDfXnoblBf4ndkkTxIKx
Ljia9Dv0gAn9d4RObUH7E9JW9UiFiBt/icV0tw9UWTvE/BM0OiIWE/mLQxI8lKdN
3OSKk30aFOla/FIiwV9T9U5lBY5czt7D1oUBXNrMpjdwH/yNre8ldioFXckokpa4
F2JXoFZQ/+2s5U+xixotFkOJqVo0Vm2T9l/PTF8FL1oVWkRRu8FMsXext8BfAbz8
xRHKEj+WJqCgT1X1ES8R5zewNdJlleE9eM7yLpqKr73GOQe0wbginWa1vo6VdCpw
LNSE7qta1dBf2mtS3RnTJVowLYlJyhmBdhs6XJQFSeI76Zd8YsIokz5Fs1f98s0U
AbilKsCMk6pDA0tK7UuMMysu+JUTHpx/hWVCYHEmb9BnyEYdKMHLivy3N9uHTgIf
G4erwRUF4c8CF/4959fsNS0qUmrBdpYR9xLguIAuJ2F68jKRn1TLRkz5PRyBRJOt
rQZ8N0oy3JdTq62ZZiVIJWgMXAT0QmJT6rh/UQFi6/B0XbK13h5rXTZU2ujc5sMJ
yzBjhaJ3Dhrna0J+Jahcdku0PM5acoDuhdUf5yhB4TrfQZ7L03hHuazc3P7sOlWR
sx+QAxsOJh2Os3dUEvF3CXvrQXIkbdy8x4Vx8szOwUcgGXtRmPoD5Uwp2US30g5m
2wObB1f5Hg8cAecXO18Xpli0rKMtcqm8Hr4Imfv6BniUpkGLrYjIvecxHFFNbuW7
0svi21AAAE00LxUZAHlycwgsESHGd/E1GhwZK5hf0+LHfrOG5cCziM4hXDb4JNLY
PeSsVsgMm/PonpOaWwG7uT5eTf9If8Kp5eOPYBlFoLF/tg13d42MS6B3WNI8dXLl
DUVknroYRvvDs9uG0kg2r2URXBXmcOePuDrFMqfz+B9vnxjn8DNeSrqUYomjiEav
w/UwgfL34bDTl5o+7MPGouaxn8QRijEp8mrN+lszbtAYY1+ofi/LpVUy911iC0aa
uRFVqyDUtLSvr/RdJmkh6jh9ChoaU3GjP6PSXoBkITf1eN468qs4EGJPvY6AbiOy
FVNWG5HqenY8IXPOe9ELa6LrfurjGU6BHxqtFYL94Jblc4AuGl6XmF02VW6uVj1R
FwqsgR+QZPdHI7BL7aqLbbm7yGVuhP2dkkdfIpoPBap7HokMtqtPFNyDQJSNEY/Z
EbOqpSpiQ+JHwYUNlnnT2KB9kYM9vc76VJL+MXUfYPihX66xtvI1dNQw5i3bZLWz
KBEGhAZ/MOH3r8254BTMDqHTU4j9ZOi7rW00LOZon6EeXJ12J9lnKAVgX0y2Qbta
5HrVpQ6b7658dYFJzoST/8X2IICc+qP8L686xGbDZlu3t0+H49+PcWL+5kSBIi/P
eOLmOZ6VDjnilhBPYJSI0IisincKqTU0OtiO2HZ1y0hkVZjst6NC6hWOR1Z5hh2y
Gk760+5bnsHjBS9OuPIZm8nJoZwmWEBP/mW/j734Bany+4eeY0cdPtc7X8OtaICu
I5pIOp6gY9e4QHza05q6Wnn0yaPAzwNOiuw9x/t1+2e8syNrRwZjkgehkeFxpY/8
dQ25Ng3/1MskhF7vb/UkUxFYI51oVsjoMuwGVLL38Lrp84Ojlo4UBq8/4gilwEVq
UC/oOYhtL7hz8bE7ceFrXUj//28kVsFlsm1mq/TOJdSnptZzvZepmAxHZ47nSwNw
/J4DNEiLGAnyFeSGIWairPDYKYYN7uIJWGW5uFIVsv8SJfW0gNBPzyQq0bsV5f2e
V6rHITQrZBQ0NyBdAe980rLDtIAtgJujV/xKDnYm+TnHwVbYhvtrq4IeZw6wCBbQ
yRqmYTaFfxhIz3W45vmVDjx4t4+eImopfwpD+61yrSitdDQGf72qWUDhoXzvjshk
m9VQDInCsDdvfeSG7ghpIxxJN0/5dUi0MnRzxPT86Q5pL4PAIttA6DHr8C0+klnj
cwnbiE60f8M7EdbapxGXTQPOkGImQilvyFWYNqzGsawHZwbRZ/fSQ+olIKoVTp1G
eOn5Msij4iXDdID7I6gWuBommy1EZ9UHzUrAR74H67erxtE+7HZK92BYY7Bj6+9F
fbNmDKnNv82s12IvSHtCbYewUmdCdTzRd09dW7u+EcY0kzvEU4RdptZJqiQdX9g3
jaajmHWtvoH8jGwloU2dHxiwHVSjj314ZaUgt5bkou+jFMpyFTq5H3NY92Hv2d3f
sscFG4t72wyjMNhn9awcDZ2LFltKjlo9CRD1VWTowmqTIdV3/LAlvOR2XURG1Aqq
anTmM/1IocA6xnk/DBvpif+FsH3OLdnT7jcCdE9DB7BSxovLDBJd12eUjMKImPip
yMYp3HFs28xA6GLXhy8G0sTG2aS8/tyKHOxTNj7QsWz2Q5bFYtixM786J1z3/rgW
Ht3MSbqZzDK9jOkgS2KRFsAb6tAHc5G0HZc9kNrigA4Cb5v6g/AyTzn2bm0Cpd6j
xScqK+vz1DWBiwHXzmfLjnUTrfAY1OgnZqXCHnWgveaIhr9ui6jzU8XNHzZhq3M4
g7uz6hMt232sMHRrwG0IQZjt5JYBL/3h8iERbjg4vJFQtQJDDw6CC7vPWIJxcfJ+
yGQWOK8idrIskDZLKKDlVdFwsiUfxNUJYU19JWSckuu0E5QC183GiM9sd7s9knfC
14SxyoRxZPu+5baBGc6YDTMtjQz2xGyutcqhVsHg8tbWULrPkl4d4qtVKiYFJA/p
HRUGNLOk4uafv5CjWYq5mLHPBlOstedm95az7oqcTFkYtyJBaifzIXXbgz/BrDQ/
/oPFBHyzfMODZH+c23EHI92zHLwn+8sv0Ep+glK9WPyWvMK25zMiuUUCemBDkSac
hjYNDwkaTNLsZoG+1JSC+6B8BiOxqBEb3dLMNaJX+LTfhsXvh5WU3/zvaBx4Kj8B
FelyY+wTrqXzB1A2J1nVF4v7iLuAGXKkxgnD44fjQGlrEHXJRnqZeoiJrHMgaV7F
KckkziRAcjv5mc9hIhh+lPR1PND+yCXX3gcd6rfWKsO6MtiUlEWD9YCupOat/rb5
is3QCQg8R12CH9EkSLPjYgj+8ha1idk3TdJJaz9lK06fGuETxGxr3uVe3v+0HgKI
XbVvNBW2eE5QwLnJLrqWfQ8LRtPCfJLRjSSMSXC4MOhsnumtYOMM7AwpSuonJVoM
e6btyF271Z37Ew8yH+AwCGnQLP+np17JvAOP6kl5gps2jBiIr3nXqOCj/mg5lSuj
bs1lFiS/kSSr5xdSH3Im/gmmajk0lW3Zguw+gNuWj1kUH9Cp0xtisGl/qK4k0tj3
UIwxtGQeFSvfAZe6c8XDylphovKvj6MO8E2KHCghkbbK7Tljz1B1m8WQ0jW+Ukxn
eGyTjxafgAbHGs1uHPrNAsnqJ0SFopw4ewFJ7FZw0FFu7O+Q4E/t/FrWnb6XPsEh
C9jfqKeM109Orv5XiysUFEZwB46P+Xf6fL7pdM7mDKlZvDVI1iyaipD/CG6Or1Yv
lS62hZ4IH0MinjJFOslYJLZbaqwrt9BAmMMZkZW5eNC4I5rgmWyLmzh/fooFbIzo
H9bjbwyv0zP0jIpVf73L4HLNE2PIFbIBy8Zc3qIBaE8EgGhk8QKeHN92X6RBFdaN
H8eBIhfXQfXbp9C5IdqOT7J+O8Jrmh26YDyII7aoH2LBJNVXzIHuXA0KTPNJrA5u
1BrclH9ST1e5SQZoExQt/7XdKj9jxJTED8UYcvoeAVNaclnB4uYkvjIi9xgeMnFe
3XYDQsii96xMitAnyDY2p78k9zg1jkbEPa3npmSTyYdJw8VgYjJuiYD8CFD/NC+z
Oae5jXIvevzCL8LNXSDubCSRip4HfLGYtm6DmK6HcQY6RipKmfo8WrIvfN38pUPI
1L9ShbiBhtKC3KM/qX9NkWawWeA283laHpk0mE9EBPtrPf+wXPGG629Xy6vue8+C
j4R4UwqBbtsURKLtEcTt6J92mYXwNsRJC3xMDlDJUPmZLBeatXt1bcevnxBY8TZY
OQ+oIk4kGFlyJN+ONIE9WinjM1HJSYTyqxpxnM6zN8mVyRNUQLrtIPlybwgvKmFZ
KtcWOxGOTq5u3ZRmEyzEiOrR+vpSkchE7bIhoJCb3A1D4Wnc+ly3BDruWLisYetO
4/nQSeQvt1Zyf9YmFARlRwkDjt6ecSg1x6IHD0t3A1TvPN6hrWbjZiaDXQHUTlLv
Iq5vwJIl9YNa4deSdjEVzWbC8H7sw2BH4A3ISMLld7ydBTyfAIQHrGiYQz4m8qtF
IUGDPv07XCP/mkxd8hVhi4mLociTpCYUt1n7sKIz6d1TdeRL4Qw3305wjS+VFRsg
zmSLezT4ckrLx3JgsfrWMilqLvdyqQERFjEnPLYhAPYvzfAusxarDHVekUPmkBOf
v4RtJsNXqbnj8nVQLKovGBwyEYS/trYVx3Vl/X9Gi/8wjzQvoPDH+jDPsmWy/rch
Ht5pFn2P+r1R9dEi0q03jA3zDZ6dM03Yj34+Bj0CaNmvqruyZT3UiMfcHGc82d4c
JPoKQ083w0wN27jyI1atXMWatkjLbBt7E78GAP/Dz8LPVO2tsGCGIPLk+kB9urly
6L6mLruN5Vg7qH5ZmSOlPtRjr4fGkpq6x8aWK7lQRTelupwt1TfmAI6agn1Z8Kr9
6vUu/Q5xX6UYlLyxe47zoEHaAlzDqa9tb48xIOoxZiffzCnKa8PQusyEMIYh1oSv
6EsQXcsW/iXlSUmzLvQxD94o5OMO3+VPMbLVMnzw3B16sv8xdNDB1othFJGhL80H
pf9yqibaNqvYX0xnMadnLhh25VO9r9fwVzT2JNlfN2o/NMtiCEAlse+QjcgslNka
33PBIl1h76oK7+1ahVpKy9gdtldUqYbcTEZ3QtSRIqpX1Ma/XFfM3vZ6fJJaKMuS
SYg21oAOXsgbUUHCX4CJUrBobTzHcxiFBzElu285RGD6BermUDn1Ic+EWzznGFLX
wGGj92eKtv4KbtAfKb8/Ml5n3flfIdFcvQL7jICpJMIC6zPVAlMObt5iU3MFOT0k
33K7ejN6VuEbWmiV+/n3VwAFRk0Pubr8YfdMz8LatgYzic4ere6elI7I4ndfsD0b
c7rBFCRljXXS8YQoILguSLAnuGqGV0tfKj4bqsOwT9pG1zbSlZw4xrQAg2OtwJtR
EpX75ij4l72gnnKYVrG/F5kLpo5jQE+zpluPxeuBg5WdKcuWWBdHdQBpa6bV+ncZ
jE7WDcAZo8JOqr31Laq2eCgmuucMLmEWOlbz4fuxwjLvSXwA7r6PIc2laPxPIWgk
6F1M8YC+Y5vkJopepwGuvlXT5ge/ohSS8UHM32yVH9OgkOvW6iMb/yLVkC/zQdiA
t66TssT8j4qmBTMsr2GFWC75e//zE9H4WNzMbbNlmAkCU2e7iI2R+gOGGHIXXDGy
+LzTFutlQ9c69doCI3uIkJnY0V6SK5bwvoFgwOsBInDKfo1jFwgOz9dv7Z8Z3b6f
Sf8Vxq51cqJur3mEnOgk1jrm3SQc4PSgVkHlmSs+OCcT/tiGVrws2pzcyU0l02iP
6gWX/2ihBDBBYA+Wg8okZ6ao30Nu0xT1S6/hAICF81Mr/HXUpQPWxFOQPN0La6s1
gAUDFyq59+UarXXwLpmtT7P4clgUO2OFSB5jCNcLI+djFu7bmAp1oyA31Udug0Y6
AUUGe+kziftHO/2/HnLiBuQEC8F1V4Yq+C8tYErDAG5/TcciClWtQ63kJumN5F8k
Kkh5h3xMNYz4SfCALWFGmf37GSL+h/QCg+9f6rB6eqYrPaq3zvQDdufAUIe/JaSk
0JlbXV2P4jfYCT9tJ6UbZJWFCvo6k2K56KeXJp+NF+oIW+RhLpoH9NQWYYeKuaAy
Itsm/QdmsKdqdnVhoAeWcviTVnxZssdwEtq3nXrXfzzzWJvzKuu5WEJvGUtw+TZC
AW3cTcWYLalARlodYorsaflE/PyDzoCJxTGbOsFOs8I0kFankVFhKndCUaTDqfcY
hxeexkmTiTNhLwNEwlLsefmWd6C227KwEfx703JdOCh2kyz5pU1Wz+2UWG4X6oLA
OvPOImRYWfw08gf51OI85HIiP/5XgrhUAcdZjkhhl87E1nrYoWr8UhjxrwPwhXn3
2XGi6CKu8+6JJjZ5KuLSu67rkCRPLVkSn0LHff3WZtFtIlqY9pt6zqVOd5DjvW/O
KOyoLTKDMM5ZtLJXcteBA+gXQVEroWvIdnCr6QpnJd1DFzS39pQMF8Rx92sG3Jfv
s5uclFYl40eF0z/66p6XN5rbZ11vC4kk32HTyh1B5oyKpxlvYclx6/rh4HWECzU0
AZeya6MuD2iv7K4KrhEySC01xCJ29WyYcZ+pH21auymxy86FtaHn8OvdERhu1TAL
ivfq2cTpckb2fhkiTcXPp3PFtLHKRCKPuaATpjg7yxqHeGQ7K94F5vp2BuTEVVRp
JX212b5ie4yAsTl8qZ+l0RdlIPzP2raoBwrXmIOQFJ+TX58JyEi4FXQD1CweHx7e
44hKkvPfH4qdApT5gd/SpFKcQWXosSAXYd4nLKP/smY2mpQYGhJLh1v0wOjy0lDU
cCxbAA5fOX6LkBMHmZLsvMka0bZ34OJ9zxqJLkBn9gnA28z55h/y8SvFW5nYnBGl
pqKWnjlWoFr+BT+ytAlAL/bSLomGgOCgyOYEWG0xfOUlLDHLcJSUjrstruNpA55F
3rvIcT1gkD4hpsV1BggKIty/miIMqJa06heVC1LSTUI3JgAQ56M00HL+Vmth+AA+
1EKkjUPPqKmsRJOay6iC88r7TAMSKZAZjS/iI+FaCTIZf3cF+wLDo3+N4jeNE6df
DfiMlA4EbCdPRGk9Pl6QE30K6jqB+Dq51/8+q6z3kbVu1puuhaMbV6MnCj0scqC1
zbTePf3bMxYSQAcc7+e/QrLaCUkQlLZTq1qzQ0ydZQ34/NNNv/GP68/GXibHOy/8
j83HHo46r19zPdZvabUQGG2VzlQBrPNSk039RcEO2FNfEppSIsncqcYQr04DK1FU
YsrlWxkiItXawwBmIwAqJyQlv7u0g7mYbd95KKsBgZ/oJZl7iSttbWYoEfqVTdf4
2CdEAv5A1K454bcu0YTPB+6VacLmJwmgxrtwKY1fZsUD7GDh1VxTbeTwusa93XeC
jjovHZnUx9nm5WK4taMdHgXDXWQbk3CN7lmnlFCfod5/hrwRHaOaepq0PgOC5N9x
D4nj5DAQt79GJDzZ1wS1WP9/fkr7FtoNY9dkxhEYXz0Oh0pLoLJzzXd37hJdYmo1
c7qDitiXjiBrAa/oBKG8h6fgVRCiru6KqytIK7XU2U8hXb4WMJ6lVFiSivZmfb/7
++PVWUFnABFOzrSK2wryYf4eGuE37/CgqCVjmiUmO3+9k8r9onQPDZOWIZvNKLnE
nUgX9KXIWr5wO7eTaOjSy1t2JmEgtZcpE8w+HPnORuseIarW5EHYoM5zihvQ2oIM
W27d74iOU6cn4lt1RsKOpA0ZzSDHcO4AOYl5YtuugQ9e2fJlPz3herr0Qg46z6i5
31Po6IAZ+lajVezwhEdGON51FjgGRRrdZHkCSW/j0P59iYD8iVQhybY49MeETdnj
DNrC6BAfFo+a420rYZ6fQ9ziggIEpSY2odz1HEpMLVRtV1JhDIc2GsI2fNf8maVt
DDS9dczpYVhRigYYYydNzrXVGYHBeAGC1gyJfJzqUWSb9eyAbgdh3yrwUzMKzp3p
b1R3oNHEKX1LDu3JYmBsLxgcVsMrxOblsmK8gHTKKmB2JR746JVxLlVEseYMo816
mShJguQplPeiRIj35l2wyhEJGE1Hm7D9fohEnZ6YQGJZNt30hPa7AAMQ47o3Aldd
FP8eFxeSht4eEQU+LAc4i0/DaEnsMct/3gSE9Kiwkw+4tzg8TrRQgTUjnnBCVUQK
1emrtRy4MHCDUnKmnQzunKhVKUvmEIpcP0eipkl/0TpGQFonXOa2pIplfl5n3uco
uAjg0UxEhKT2K00di5Ufq+sJj6/79hxfdznq/7SonpcvSeD9M4dynRvOPNneSsnJ
JudY1y82J2Zxv12wrxQtVYuBnow46E4oBvrFuWvuc03tj5DK6QUlEi+QLA+xSJsK
KfY+NMRJEjgpEKXWYrr6OEQRlIX1vo7cjPtr5cD4NKttczEEEqxocBgjTv7lzj4Q
PbHdIrjXdh5fbQX58Ea51Tx8TJ7HnGErkq9oOBAxvED6732xNZYHcPx9646iq/g3
5/rqUucpO3V6Xr6bpi7iF7tQTknObd+Gj/OF/7V2sjYgWebWuN1k6HwEat0OIFds
vGfjlinUyGqbvxS1wAw9lvZZcYUSj+SRhKxq+rB9C8lh/F0ioS8Fwb6Nph/fSY+c
5Lah60GTVx+49lGR/B/8iVIltGtjK3PAWKVvuhHDuVPf9cDL6I+UwxJ891eR8n35
Z0geqdVTamhD7LJVT5VzJh5D7wWCcSFcqA2zvAgdipA2iwooZtdB6GCCWqgD3vky
2XWAsiT+SGw/W5QjjIG2p8eYAiRrJbqOmzRE1nT9xwaaMGmlfHE+GXpfTtbJbcNu
/BdDRKaWe+efkyMdkF/cE7uxOiADBZPpeIiBpyvPL14SMSDrMvVPTMt+fM4bPayk
jw/DMf1AJaRZRB3DjuFA5MKmD8gq0+hOkaoDREtD8aFawaMPjJvAPO/wx5oJpG5u
whdyv+7ucBABvKWAj9K9UanM3EfOuqxBhiigbKo5OvsN1oCWdpMoESnuxxfCBryA
hAae2qxo3Llk7zs79KhpJmNEdLAigZbw5ivflTCZFZ5SWHl+pwamhwhrJieTK7FW
kbUSWH+Js5C7FGIlEfA+4XmCm7l3B1I+jEUYqq5TTW1GpTR6RyUkpH4J2vpjT27l
rLj+yANvbHkhRpRLxriZADLayfC0I3EUekduSAQ8MR9iK9hRZ/ppw2p+vj+6bhKt
hk5Du7LpPI0lruTnppr/ouw1pcPkmuopy3P96qkKI0h07VbvUZGS3u7UzPnSPoZ2
i8xnwvzCT0BXFmZRON+XihJqpibhlKmNfXjR0QOiY4OISUMtcGcr+Nwz1Wah/B4a
NV3D718ME7HzXHIYx4mw+sHJHXZyBEeMjhIvYDw7Y0BTMfD7gFAYa0o7FPg9z2MB
yzyKeFQEL4d2ASn9ArPQviHpiSKoSYmXHuBNMjqJejRJrSz1HAjzBCosKCsAJ1YZ
3VxrAKJF+0GYabuVfQ7MfPms2dt6qVNEDX6Mzg8lKA7ER0nz9C/LcSIZXgq9LhCy
Ii26eVgBGwTxbTShD3lym5NTssJjoiSqhWonr0SlakqDXpnrNTR4f5kcKnRK0otY
z/HEJZOPx+svPyjfn7nHhYoqRpyyjej17aOkpbJsCUGjW2skOykIhA4Ts1P2m2u+
rSwtyrtY9Us+wTke6zzn67nOUDJz0PdEMnOF0bZQ/5aUc2O758Y1CPLCP+eyBnSh
/2iRjW1EPakXb5qdewec13ydRSI+gdFjuRdayJyP4dEELZ2z9S8nRc5p0J8RHTio
ydZwgQ+mx1Ftr6wGPeNH9kAvCJ4t8cMKg5hXDbjHd3RYXbKErzatox6NC1eOfdNy
OBj6cKJ3+H0Q4jNasZw6zQzQZv34fHp/7PQPNJOy9bnNd2Ca5VvAJ9hl+tQ1rEqi
UHvh/B8vXoT4AAOH/jNfN9Fa9SMzcdxjLoyW4DroClEU/89rICQRHUDum9m8BKmt
raZsBoa6qdtrrypPSC8aTI159230jTFByZiKtfEoBWE0QPfQ5NuhL8x4uaP77qEw
931t+9iQZAq+dGvojq61oHTLQtoe3hJK0uFK6zLYhC6x6EF1l5C1mvTxn4+M9f8Q
RG+FKZ8CHka1pm2AZ/BQbwto4jAxFjss/mHPydc1VxC3HxvqBs/jKCj+Cc3Hq6/m
TVD0OU7NgC318fjEpQs+fS2qk+FgTZZaJi8oihM9Q9ArmyFqA1CTVAAfdSNjej3D
qwwPmllFSBemkwnz5EL4DMdfhdt7LiQQnDP4O+By9YTygbdvKiH9bLdhSDGLS6SC
JgUUG4voLY0KZfcspAL9hvGAUmZg5dysnrdxH+H8H/42SiQDWKtXwP2YwLJYnXDy
S8FxxvmL0UNMpQNSOv6Z8xTbpX390BO/pzF1B4QF9pwuBNI70QEWj88wnl0bZZ2H
XYSaqO0q+c8EONAcN6dIA/WjG42ssiw8b+B61JQCKnKeuYARX5JzAEQDbVoQ3A2E
vFZCLcmCf6lp6LwExu1GRyIj4fX96Da3FqvQGM6GNv48tDDA0uR/3UOsNHTPAAhd
+k7hdoGLbHN/ZwJeG1fyeukfbTZs24nPbb28czb4o1zEUKXqW5dOLdxPq4C29yN1
fMlxX35lKAPCSChdM7T98vkI2fFGTCmMzpfwI2KE6oqMoAejHmBpiTIT/lb7ftVq
nrnCo4ido4pSNxof6Vx8JiPGSoTGrwZHbWW8+PnaFjYJPQ5N2sNpjLVLVGRYqWJs
/7vq49+ASzeeeFIsrg9r/BxymlIGkO/bnBbL6HHjLmJoqkOMtmFsqOMWUkLZfkqG
ittsJ3zY2QGDmkrKP4CAz3MJC5E1De81MsIaJrbPO7CZriYJOmERot+tbtZXUg0K
4/vluHtjUg9RkqtuZA2JdYMGYhS/rXPRTo3+sdA+p1qzE/9XHXPO/G/HaiFvv8OU
JDrm4bc7rvs8mSrsxtcm7Wa09oEHQVYYf0id1ryxyQqVKwQVPlotcF4JryOaTp1r
qDkvjfcE6whR1jBPbQSVywIjmgx9Lls/rjqnJ5l4G6vJ+tcpLJJ2KvB3IoErvkEb
nV7PpsWHTNfBLYUV/qAXaYCfg7AmeBybfMLCxMX22rYcVgCMZjZjL+6sxwShF2WN
1Y3FWOiavorHetoeCa9v+1g87NDXRgT/MsnN/+lNmoZ6RKFXxr0uhsPDpxz3yy7w
8zeByYxVQlfQ87ekz0CnaIe1PGe29VeqxPIIxyzobRbOM65K11l4PRoQ1Rit6fpB
N5zrht++CPIc/tcC6KY4XVDumxC08zdm/29o9Qi4EqsxwYeAw+SoDEm4Ug0cU0Y2
tZVA1i1LPO63wyi1sFOfEDtX4y1ROx6t/26yKhhfenw0YO0w2nv3pdWqfNfdfp+T
c7JHIBaV1MwieFuMFxg7XsV7/5/XJ8I5l4sM4vwR6pMsgFxKX95rNLaE1ZFYb5Pg
Yu4jgNDHdpGJ1PzgLkErfhoXKxGtL70UKjixUo3Ird8SYlp93qHnB7VjkzywbU3g
dQLz1Elz+wwmIzTeQEsBhpcoiadGGtWBsdMgddSFUNfuQnNDTd2Tq5lFSTyrTnsP
wcGtl4G3IQLREthV41VDfbkJQqV4O/SFfUDPhG1kUX4Yjj9KfzlhNcNHz7Fts8tH
25+eZlKgS9dfIFxvzFuy4gDafFVdY8C94PY6z2NvqulUe+mnl9CeXmaMY9O1N3CM
oB83hnWFLlrFGzl+JpqhoiF0fhPbcXhcER+ctRzacPcVJRgR/pEz+1iv8vCGtN+1
/QoIk/wCyq/UsVCh+iA5JZfp/FNQG5KBVCYfsJmiDtlBjr0T3JumEsjvdEwtGZdA
CgkpsoU2wjz9Kzhr1PbDWoaOplls0WbLG5Dq/qmanbF/KjuHmqlm0wEfvrNRv/AV
Ps1kcGLarjwfcMSJ3rEPi43q4ctv24VXCeeplbSP0pqgP+su7soqOkNXq2YvawTs
nhsUR8l288kPcv6CZgorvV+LEDv1sV0+DJsSqHl9W3r3OR2Dul0Q3FuYIas+945F
bzoy9PTlCFlTu/M5irg+OBHEmgsO1VmgxbmyrsNmfR5UzTxZoXGqa76Lry3itX1r
2LYdIyEzzbIQG8zHGorIN4NrLcDle5XP5FvnxAFTiDJSWTRPa4Z5+hOQSQAQbnyZ
nYfuBVOmgF6sDYuEWrDfUTQ5ndCytbsg/Dq2DRlnRVlo6eTWgosEnBEnsFhVhy1e
BjtrrihkRPsLBekZxZ6Cn6pI3FO3dw1Bkf3b/vUQVwE2juAomlfIhHKSm+rAxFEw
UZShBfq4O1Ktn4ie4+JbWe2D49Jf027VelbzRtzZEPEFRAKo3DMO5kzLWVcMlzx1
WvmHh4PhKIeA6FC8V09G7xsALeWcxxuqpys8opoAel4B6/tdxx8UtksMlIiNi7s2
ykddNXDso/SxSjKGlo/nSpkQjpvH+9HZGNxJrb/KYWFO3IfhCXX4LWJ+KU9mS4eM
LqrDIyQwllpXlgydqZfFGrmpVN+EATUzAI/iQg8a/kErg8USWvx2NzHSQMdyggEj
a9pC2hFTq+TMKQkuVUEEtFIxuItbycSZx31EkGV5rYsIdLCVDBh1Hlpact0dSKEM
iWcbxwcHsV3x8mJIgsJ21nSPAHJo8QgTGd8MOlLPZQ1X3m9xmny4MUQoKY5woHK8
d/L1iZf+7C1GnDFvA4hnLMg/BB8IhFpvOGami+xRyu0322azxU9HKZveCEg2dwJc
L9aATrrrJCYAgxoywSu2W1nLiKnkWUEe4TAznmDojfRlJwkLaLpuaT8l8HqjHX6F
HHMfbibC0ViL3dICG5xgmhhvcKEAKOPb7Plr7WQBd3hj3CrYbzGnGHppHZKMaAhD
g2q2yX7YrL62AMlQvT3al7sXjt+uUxa2RY2Ssq1+ApQV0zxhHq2hPaJv9mwQijmW
9ZloArnwaZWrBEqYu6pg/QWSRZtmRHm+0j8dNQhnT8JcNN3EOJBxzIeQcsTvWPU0
7ssPYGvPKWPYcqWZIg1AHusrKLNEY8tXv+v9Fx2ZtBxOLbt3+tkQcQ8jeTlgBERH
Y0Er0GvTP1ErlRv6bzitPvjvj58XDQty7FF3SeiNJW/t41OANXoEoZUKD6wBBbDU
iAlw68q8OVyLP/2tctuqIIYINht3eYVlluXznuwHz7Fi7Fdfqz512MCDJtJdqiVy
OpjL1f7XLBivSaxBvQX3TpYVUrfUif8P7cAzGx+CI10UIk0sPRp+eVdHSDkqSqIg
NKc6WsVMnC24GBLYg5eX9rbq9Lv9QkKHhWWzqV2P9kAJdfPesH3f464Mam6hCAQp
mWxyDdNNsoilFSEbyfaPLu2I1YKEGzrHxBH/dgLm5l98dBaSAqxGdPcsEabkr7J8
Zevo+sihQRb54P0dOg0sne1B5fx6ZsqGkvI5HYs0XXxoT7Abrxx6f/1YoB2VVGmU
KO+yk9V4kfQuCzbJ8PTA+SxupIcngfMZdwuPUeNqsy+s+B46gWncSn1EaORQAz84
NeSk+zSJIyD67VnlPeSlU76oCayo7yKL2srvt/sqUqGqpnp0QpIJx9H3HodWY0mJ
mLFyq9qYBhJSeRZtqWtLTtt7aeHS24YB+G6TdrGx/ufdaJWNr+hA843Qsl6KkYn1
KqEfjZl2oRmyVTYMTy8KlRpnqLsBfbwmnsgacchu2InhrikJ/3aAt2SKLHZgcSTC
JX0+qwmwj9U3Y6z2Fx6JCGtiDm2RlhzGurnW5GyKkYzw2Akvhh+uLFZ0YNr7he1+
WAEWZ1ZJIjx5VSjK4IAMgvBQ7n+9O9z73YFWbsXZDeO4vMM2MnkjGWOCXaERpiDP
VNvz6bP9VTnkIlF3GMXLQPrtBzMAN09E/A3c+drjp9LV0iG4B7eYU6bWcm1vNjp6
OTR5jl678fDldSXgSex5vAZn3UGD3m5XW8COTqJnjlmIflUNjWY0VeTZORqFJv3E
MjoaYKWNhoTKbD3fDiPPBgP5tcMLEgdq8oAt4DwL4AomT5VCl/wBuFFCSFhmxG/l
H++LVNtIyaTphWGMMnVr5eFJlIan4zbd4AS8AidigPJpUP5woRbJkXmi/xWous9R
CTeLvuAGdeIkA8mkO3/c+uSbh9igiZ4rpffixpdg58tIglyZEKYSeM4EipZXfvud
onhaphGMZIEd4einwKgG4rbbWOcss8N7v3OOvH21V9SauUPcwqA0Xp11ZHnIAnfm
jlK5SJuW0zBjGBplfdPt00HOqj3djPxnAiFj8tJouNExPSwKSLMf+hhJDv3kf4IS
dbCHcVVHmkd4B4FGlgbQ82qVY4ktMRA8Abn8TrHYWITOO6gFHF8DY3Fd+kgM4OXy
HfJ2acBTcbkOGPwdMgkCegzaVXfJ/E4m4EvosBL1ESXJskVASn+NWjcKl9gZejqa
95UaAXMks1XA2A4OzZ7DfXeN0AHi/EuCOP6i//kMx8dFC29b1wr/UFrfi61dlUgf
7ksHXtvRZpgBKVg3rb5JqMfPqdKlfByU4WafiyRXuwM+zTUu86hwGnWnJnB4DQsC
gMI2UAUkK2s3NRaDaIb6F6zD4YSsttqAYHKYBV1tqlby770n4Ts1JBEtPiU/qrUQ
d7nIXps3c1IGvPSxhZGvxNt9G+WL/6/pKn/ALkV0HXn4aubjFXiTXNlP2zFF5/FD
91AYV7XLGovasuLqedwNK50n7MxBKvHL7YWKMkUC1Cje/fRVbhCPdf1zSWCj/TS4
ZM4p0XbJWvLsN3GdADF60zoAZ0bX89Bs4cQHjxD3Mkri/zgvVx6k8sxHq1T37IdW
uPOFXs0ZjGL0qV8uYzLV/B4NCof7R3VH3Nzrlue2F7lek45ze+MBp1M2xMgI33HS
WuppTH0XN8j90Zx6zXWLst2wBVUfuKj2OZltNCSMgpEqX6DcL6AcB3j0ffud4Pbu
E7L6xRvxuS1qNaWv3KNgKzWguqU7hZyFNrpdcfYmKLD/xAanAnnDl10Hm+DwXjj1
BaSshnYhILmFxNeDfHq14/4de5r9VPdr/lReq//i4seDwqTCyDdh0edZZKoz3PK4
A2vQhfr/RH8P7gUItbq0KkYnxWS3rqIKeU+0PO7rdo0rn08ZI0p8cvyZ1NJcvgpy
TSGl/L9b090+ASK8gEg0+KdL12r3dvCYHHs4JH+229jrZe/WU+BbTk6XlPv5iboT
TLXo0EGIiWBiFurXzs+8Ca/n14MdRhWGoq14pPrkM90ztyy0qbQ1PcF/Y9onhDsf
2nOfAewIe+oCDpB2xSmbjpsX2J4QADKZaKD1ikuyAPyaP/I3zXtMwOkyVrzYTsbi
gmvGRSpkozW5wKIXMHQTCkqDATTPUshUevp7+bgBXMToYSNTRm8LDNUbBIJTaQDk
MEcqY3+fufj5T1PJH8l9S48KITkvwKYE+Qs5j1zpySZygkV3m3kHqVyir0FvbHNW
qv4OrFt3DaPwLtlwQR3spIS2G4FieM91n6iwspsNsX6Yf4+gaMZZavBrUxEINdN5
80WxTrqJOWMTi3iGiov2lN+919HDLWDnL78oFJ/z6JbUGs+d6Yjv6Q6udkM+FVyW
OASE3feusvA0PIi660GViDNbJTtpnNvO7EcdngD4nHvKutLju216XGYAQszJS0SD
s0QEn732TpKxU6sbaNLb/bQki4+hriY83NqroXZK/ujgMmVtMN17AvR6MJSMLiSz
6hv5+xVfdg6crMm8PUsvkO+gdI4fk2la2dXVQVcVB5ayvl2ZfGFhkouHsBZ232bR
l+5D5M1F7U0IaCr8uQhucf7UW9daBIrAdEPMKeOkGXGDQ7ernVzW9PFNZs/C8660
+gQPayCxkXtt8vfcORn4W90OiE852RwUK8cmQ72slWWodsFl/KeLQDZdxCPRrCx+
sZQX6KI6S4w6ySHHomxNnGYDomMEl4mJRH2aTDW/1fefuCa8XCSJxQgjd1klZOV0
3EANokQy62NPOZbV9Pst0uJY8kQxW8fNLbXqds87p2NegNxrotkuJSpwwZqEPbhT
Fng8shzsYdETZBBFt/pFoPLbInE/wmnLr4kS1r7vNwm0iwRoHhSHK/we9L1zdq+8
wLfaYAm5AI6EjvjLaPTSpUaMM+1e8d+ynHOYOj5q+WNHpDR5G/p/s7dDWC35M1jX
AmhPd5otiknOjNPXooHn93a2x420u3r0vCLIBgXid7urSABwTMjlBUY13WEB70ua
XMn2pJoxcP2ghKWXnZ9OUCyhEWRnmuA5lqzezUjWCRwcrt0QvaWutyRt6vmFrZT9
EbBPIgmWHqDgiirLvyP96P/fZoeAQlTmE0q2khfjvXSkYqZ4rcDI/4IfnTEf/Vqz
xpmF6E02GCPB19IFl63/4tpqIZ0sB0wIJC7O494sxgWy3vImdAgpjtckGgUjfwCw
lFC5JEN4QAmSpVLs98ZMnWHpZK0ub2NQusGP7G4Djwl9y0hthviFsjbAhEFJ79cI
59wZZ+ZbDN+txjMd/ZSVXL6gGcLVP0NdOmaOF262ugHhf+DSGCNlEeyuZgRZOxLL
Ljw+bwKXEJHnJz1lyXD4HAEaotxUYlyAjC37G06Izw0QiXSw/0+Ci/edJOMFS6ur
k3NMjzH2aCzfIojiAS4Fkm0gZG5sXCNY4a3/TJRAsLyqlYCJI+HsGAK9BkRqjbdl
NsaGC6aQL9Zg3rKzi2NQffUlSqLXzOEjP7VFcfyPGsAD/5duiKdCFu0VZC0sDQUm
raHDPmv4l+xum7a+a3VJ/3wWPmUwct+UOXI2pSkfoS99EI+2E7TVRrrYI86n+8W6
U0y+1s6hRoykH8GZQpGHnoA/rxJ+NtFoIGP4V5uiDORjJMPnXB9EQAIFxAptc0JO
XL2CLh17J1miA33eDc5wlXLJ9roIoiOxSVD4onkqhgFCt85IWr0hPYIGaWkyyHb1
fkq6PxSzTvcsW3r6CTtgSX7fhkikZ4GUwB9HGfA0p1JNieFmjLmbJsCGrgJsGkuJ
abAxL7kiIQRkJgEsb1y0lQkwRESFdPUD4L+EshyhqGR7Ce54OUENP4jY13Pvh1Qh
WXrv/qCzGRlYUd/Z1tNBmg8Br5LdHvteqoMi7ebbcdVyDfEINwBy38ll7fBMnOMz
zZf1ok17QErZy2GbLKhUA9zJgkA6ujJMCLbZhuba4B8lxBeoozgwaRWHcpKidw+o
UI1l0Fv5rqc8oDsmwNQpri81zLfHJmcAyaODXQ+xkHLRO0I/YU4NUrxzc7wsTA5C
GSx76u0fYSofCl1S7WY3MDWYM26Ph/ptstvVWdFLPWmtnIwcwDkxy4vRqEsTHSe6
t5CSspy+UDtlY2HKPSbfYDNCM+IZhOQYSIFG+DAFNwOt4gcg63uaYIAtEgciH84N
k+dOAGcCwlOZc+7nmHNqnSyctESU2Pp7+l4GgUui9nnSb+pWuzmY1FVhZEMg0sPi
tm+jpVTTBPSPmSbUhN8nSm+rxDbcvxDcAZJRPAL4KBpGOdxU+z/gUwVVKiUm10qz
qK8kSnjoL2U2IbiCEfNqHy96PnDI4yYWSvnfEDqwtzM40KIdt9ya9+ATabyvt7pp
ZBy8pDM6So2cSa8TL5c6E8xOwexrDqoVYvfyFQM6a5B6JT4ZtWiGK/q4038Q9LK5
K19eMfR4SPsTh2BSFJ4Lp9XSrm4bW3aAAn2Pqw8JyoQHWn4AqTOCw9TrsyW8eLeI
WwV/qbxqSVy2Sdo3eKrhUey38gKItw2KuT9ubfwPm1pYQ3KCRqUeMECtUjHQE6Gz
+OFdtZaBf7kV/ONI3vGPUIi+zzAOYgo8WeMrFiD4o6le1s6vD3iX41NH3SaRQmF9
J29+7W3fmWpPcIOfXDJJ6Q40OkR590SY910HzTIqQn9MCZhLrNmlqeSNh1xRikTy
m9a071h9RNrgAabJyN92XFQn85zTWFcq5hyHjvlPECAao76FVVxk/KHOo48FQus7
VwXD0RLm2PX9yotvPADJUPS1xV2fdkA2jWQSDzTgZgFkFIkxpm2ixgvq0HJcdI74
lyZO38trWX2UfnsrBAy+Yk9RLanpsTU8icCkra5nkjIJ7E1y50E49PJHZ48076M9
qCCYPi+gtDbSekWWncW8HgHSvcFVu+5mkrm4SDEikdI2Ua2Pq6M+7evKaQ9Um8v1
nwFJZ+GlnAYxRpXLDKQ8wGXdnhSpJkRLKxhwWaWqN7jm5NTtM7sneuUk+pDn1vHJ
VjYcIlKoYIc9hLgmfH01Q0084neC0eJGXFEO7EfC9gXj7TZ1XIJMzJkBLpM/Zm7E
g1lvy+SXiSVBBG4r1VUbXvGVo9JH/V7PcLZleB3C0wn9DGEq7+qepsaZUKa7B5Ug
gDDYdZiSXbPCLEHwr5B0A+kjIA569RzyoXwzw3c0Ms+VkQ2CGAHt4Z7owq1FAhA6
`protect END_PROTECTED
