`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2dIEt0ZtfyaTp9B1m02yNibRNUXsEnJCUGhd8IlbUBSHzJTDqvJywGhowbpIXPYd
L8pmDTYJ3C5fGr8ZbUPP/WSu3tbzzJ3cSA9x30HHEPT9mt7DgDa7yG1jVsc4nRf2
t2LbDCI3V5V1Ns3aaEiV6xIzETpaR3A+VXf3TPrM6zoaoMbMAwYnsjni2p1G89Pb
Qbg1N/wz4NUa9i9ugfGOQNGHkY6WMQ5qdPQbounSW/mV6C23wSkkQQHK3YbdpA+L
joAHJG6jL0dXo1Zjn/Ygn6w5uyVLcqYn+GQ5XHa3/llrfrkx2k4cpN6FoRaGjDZ4
HgeqHZfFeENMxDbEEKPXhUOUMiryXedO9cXWjwp9RfzsDjXn2qO7el3ughivYMRb
cazxxtglHiJjwp811j8BbHwROKbhKWz14x4/QQarvmyC/wTExC/PnnMmTE9Aj4It
mMtlkZ4L1lVsWzw0tRvd0O0A+nJ/aZ+mN6jzr+YvmdWdt0xbj3UgzJSAr6GKN/EI
yjJ2eTDtRf3WByHdTYcIOg3YlLRp5snZU4A5cDE5DPnvgufYnbM7hpk5JO7zpThM
el9sgWhWsZ0hALEWtiK+KFVGC2w7iAuY/gUUG68b4ixFs9XmwoylAOb9Cmnk1LQA
TsXcb452VbvkoApYIgIgjXtMqXx4lGYV7w2v1lcUOabU+9QVl8X0EQIjzZsjAwTJ
E+FZhO78N4xYknG6+larwC4aSes3+1FyrM2fBaYenQyw1Nf6qdz/PflkTdNJBVLf
rj8sp4bnD1keqcSMLHPi4jXxzX7WTEHsFtS8tVab77IgdUr8GEaSThUednH22paU
tpng2VWhGIDsKH1pR5vFskzKkV6yjXcIOXKHQK0orv5b59YXdALap/gDtKkG125m
uEFsUBgH4C42Q0rNAZgFhdj7Y4yeIPWS3L/SThpgLzEh1HTGn894Be2l2zktg5M4
ZeAix8cuvLOiRknlq5glo0wObhI5Z8JHLlxAmCZQYGyvT6mIET9VsBF9hvpQ5PTD
RV8CQJca56X1toJ+y0rIyJikCbWx693NDSmxc5up+Ovhi4E2wgoyc7L2bJ73h7zX
5BH6Bw0K8LznThFyh581dJkvXoqVyR8wvVm1HkW6x7iEkWqRYP4OyrAWIEsMBCpZ
`protect END_PROTECTED
