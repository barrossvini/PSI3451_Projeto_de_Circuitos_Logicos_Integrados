`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/nEy/cN2pJvhjmtdvFq63dS3jyAglD9ECnV94K5Xy7ggWeYHHiAVxU8LDDb5TggG
gI0W4B34NQvooM16oufvMLXxlJEuihpWjRD3V2Fju5MiKrDs4kpqVhy9IlEigJi3
8zPyxENhHGK6A0dXVo7C5SFUSO3s7ROcCuetR9pp69SKcppmdtTRiJRvNzpjClVH
nuU42vMRL5Wl0dNztqWSXEg3YeMnPCeXESbbQBpUyowOHHFYiXfTlWhOaLhYNVlH
e5u1+LousZgvaCPD+MQim40y5gVPSKNgWlV9GLyiDHsySiuBfwY9SD5IfgtTTmDQ
I9iMxWKKSwBqhztiPCNfjr1GN00G9xyueUYCmaHRh0eMLw6ueorXbfdFspieFZdk
WTUKcFcmIfMRMJz4lIk3aZYloSJPk+NlzkMOV2l4egsmNyHcnnjSB8Hrvd/Cxcpo
D0X4RGKDrD+R3gH59prGwQkZdmTpwnZUT8CiOxs9wDds4ym+DV0FM63NXC31FLmm
VO4i2DkpKatxzT4DwsA+v6ocYYWmFVimNuNIPHK9NNnhx9oc6op8tUUuemBJ4EEq
uiHIvADCWabGBrVwpOqKT9WWNZGiPab3e43UFkdxZb3buNLoN+HTb97qK2EbwRjS
FFBmreGxwne2lXkOLoeiy5pdU+SPmNpFS4t9l54FmuwpNMp1kIwSmhyDAYCa+qQx
ZrcUKM7DEzd0g5wMQexH2xWVx/xwbquRMXK/Lp2P6BGFhmuBDOWS69tGyDZRbvSw
2YEyry7t7EvvSOx873YoYjQr6JGdAQLDFqYa1/YOj7125sfAyHQ/5b+dRwoMOLk7
fSmtO5981y07wVJjZD3I5fEUvmH8z+mjyUOywi43ms70IxVdtphjzjavkGuD2T8O
w/GVPLGbJKBe5iePWbhf91nVROWQSssDb9n+75ppobkPVVBv4Pz+ufyr9s64gVG6
icr5a1zE0ZsHTkiYU2VtO7GcS4DNvDoVWr8cnX4qolgZSijYrmTJ9+EgCZi7fYHU
RBDCccDgkz3YO3BGXnz6YpKfFO5vF4CwDFDCg8cNsChScjWk0lraB4PuwkUDJIXi
JI4ZfF++HEgI3XK5+XpVT3iR1SO9lQK6FrhITtTSi/0=
`protect END_PROTECTED
