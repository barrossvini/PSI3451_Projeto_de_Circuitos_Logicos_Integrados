`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vpC8+dVfaz4HoXItbv35j4IZgp+GQDLpRug6gEa1M+BGKM9Zdxen1IL0ui9MWYGr
53HebeKsflqNrf6w38j2Pb2wXTauNz8h7mMZkZpOEjgK2Esr8DfypqglN5TQeXo3
g0tGlxQlpo7AH3K9j6bK9ZA1BY+eqRpL5HX1OlRlJLhacamKRXX+6J7Mx0TITcS1
GYOORhPxC2uTxfJ6KyIDxKj+um2HifvZLS9ET/2aEoKfUbM+zcVzh6l564rsyYRH
NwglW+e7HtYABT/JruvrqXdvNYTNhPN1nFJrEg5ye6121aqAjywRvtGIs0x8bI+l
b7SDGI7caoQ30jG8WRPrL/TfJ0ZecD4bYE3J6DOXp/U/ZUZik0MniZRK6Na2I1eq
GxD9Vc0KKGBZTJ96TJIg93/H2y7KG6Xe4f7mEvt7MEwWN6SdIUhhVwFrPOUBHsA6
2prqh4w2BkXh+U4aug26Qdsp4+UATCXwq5PuD7BjjlV783IuMMLOGSiv69NLEq3P
v/DhQw8z3o1HWh2q5s4Z9Xj22anp+g8m+9z4A+kjpyE2p1qTWPZ3Z6upmxGYvYxj
8B22LXqfI5VPMSp7NAJQvtIqhm0qdYDKRinsZLyto3X/niXeTtYHrJY2IVp/dQuG
DORvfuaFv6yrExgObaCJzcmlyozB2DQgiTtFWyRDxNDMgc2NXqJszpRojLMb3MuP
kq5QOgqzDvk7OJoMUFY+wk49MOFmAqfyMFwqFY1zVS1YOItZd6hA+mInSdRWZdW5
FdmgzLBTK7bkJ0TNGelQNtdbrbPdsrSA8D7T8b6ksC1PDIhXtp2875v8NUjHyIKc
I+JwiiFV+hKQg6m+CM2/M4aLGf9SW5G/Fg7DulqIAzqKo5iB/ENR5w1GQWhUOhdc
H2Fp3yucYZknfcV9kcJc4kiMfPmR4hgZBhzr1FNx7UASMgMEWeBmRT2aoRGR5u+J
nA8emfD2PNZPLy4pen92dYzFdDD5gFC/lzLMVrLCKWTfxeWvfQN4Tpte5eMi/Fcb
`protect END_PROTECTED
