`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RardgBZ/KH0k6q5MzbYAtEVBrJUmtzs2xGRdxJx278AoaXnNPikrPBMsGJhZvoA4
Ee84mQcI5YcAlNlhFknE1VVagMAwVgmUqAjWZBXH8otrtMMHE8NpXCuy6ILICJ2S
g3L37R4st1iYjwhRAhHfuujUpHNP0/U5IR3j0/a8QGSoYumeM0X3MzWzZgWunPML
RaV6Phjb6Fvl5wHmWAjjGCMPAzr4yDB40umXbRyY3mkJCmthDYa1+kRtN4rAeUqS
BztbWJEeSo4bMl0P0tkFptBZwvbN/ZW55n3rPOZDYYKLEM4Xkr3LvOaQmj7hubXZ
HkO1HmImDxZSR1jugi0yRhwx83i1Pp8oxT2q66MnarJZwSpncBqRNc8KuwQTbPI8
5hx3XpJN72sg+YartbioNwNPkZb74uU04O419+K2AJhQqgA7I5yoIoUds59u1EWo
VPZXzZv5rqWclWReSAhXr8ygg4xdf9bZ6NZIoclatkxFOdJbg1VXojhc7ezFFxg0
osiMcrbSoR4j72DA8jcRZ90+he1jyNehXe0I2JBS7A2i7Qcx54szzYWEEKs8lZ+w
nyJ3Ra3Churr+0+cVFmawfEhqtKb/zuvkpJCN4pHRlVU5Y+nktK/EfKeVRZED7yD
UK2uI383HOH7LZLq3hBrmYMW5vyNgeIjaj47iVK1Q5iqhydE03UhlDcQ6/WwQiBE
pAIIUcV64RSKxQM8FFZaljz0OQvUwnHly74Mm4o/QFD1ecrwdHcZUII4FjwjKLVF
z/6yfiQRtKaW55Wfc+U8HxZ9cK7lQ+1gtIDnDFEOWlbtg64oVk4dMf/OvTCerbja
DFNsq+nmm8A+/FYX3IpAa087G92PXL1Xgrm2axTg8ryMEYfg51CiqFBqDkgaunHN
+9L2oprq2Zcnsl9tcdcuwp/mUM3VltaP55/bJePgvNfvdZzpnj/V5jjhpZip0rtR
ePMli0T71IOvoIWdi8ZaVqxJE5YBFWlc+s7uNjQeDVCoJ/c0gIewWweF2PsUlBjO
o/EUeO6mH9EbmpGK8erhx5dncbwpmz9rKsSAzayAZK/wFnqANpvCJGn0bPUOPjYL
g2GsrHbcY5qz4bKLfld9uRGcZBMKxp6y5oFULgqDEVDTTehPDlUnF1QEj5odtsqm
8aPT88bN1D0meklDb6ja5BFleNck8CkO8bTDyovmHaOJM4VhFuzV9UXtKNp8Cmd3
qfX34iIWj7jTaIrwyofy8mx6upXvjm0JD6v78OJh0jD0nQrXqXc7wsLmpMFWpcA3
8MLpDs3ghtHPIU39Nryr0CsCsU+ESb1I8igtHene7HJRhbJhGG48iGpE3ForeXgT
1FcRN04xyRzQUIO77TNqJENOetNcmXa+NNuD3OJFXKM=
`protect END_PROTECTED
