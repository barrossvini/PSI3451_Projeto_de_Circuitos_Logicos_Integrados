`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rtSAAwZjKFHFGaW38VokFHWrfwCc715VxfeuOw/YJAGbYzhJ0uRHail8b2NmRyPH
BoAiKS29wqwRqWKms91NtLrmgP8yrblcd93Rabtk4HBCburQSmjPIyGUhXtkqItx
LMs7H+8s22b92hROY3dRtf1mDBSSMpDwUPbkdrgxvgFaDx5XVuIIGuXTt3kk1tTY
DvyDWrgcGt9Angj4x5L+dbIWTOmWcxybP6XZW7VBbkBO12pk/Bd8NHmw6oR6rFfx
yUh8jAFVydNC8OWH2IPcW3S9D/i1tN59K2jHtkql3YjPZWbtu5lpzpTOc1MC7fIp
leWB8swBjWrGq1T4Vq9ffSNs8UNG7tRKjDpwq6uT5Rc5YDnzSFoRfqIxX1mfb5DX
UUZSyVFAhKjAkLOO8mBT00EJEMV/9Wwwv9JvY6tA72xs6GT8xFIpmGRK4b5HPL5K
XVs2j6tk5ofF/pjVPhCkaZymJ4qUaLmuX1cwf1HSL+hwwjd9UjRP+Hc8ugOQCJzp
bjXsGDAZIEvnRcS6QK6D0rA15SAXgnWb8g65A/psp87kL5Sc3j9iLYzw5tZ8WhHE
w1jzK2gibv1tKb0j7demtIe7eViL4DqBcT5uojSVFHkWey7XfEte+ei8wX6kcuTc
E2+732v6bmfnBut+0ZEHmpfPxxizkI/mOXozHErZq/RVkIGH7KjjsxLv3g68k9f3
jkqBRT8b7dpP5hT3XhgugqrKedvIFrVC2CeeF+x4+ncrE1EuRsh50mFrBn0rPCGA
1ZU8F3EPCGLROMIP53rORrlk+PlhvXWUbkp4DP1ILKMluvesgjyV0pwuyyrcmzvy
kZWNvZDadofxNpKgD3OBdRfWZdVPgfuXV26EDi17Mb94ofGLdj62y89RQS1pcD/t
`protect END_PROTECTED
