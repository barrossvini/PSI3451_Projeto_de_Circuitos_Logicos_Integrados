`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XN1x/JgVaiGWhu3MQP+Ai/aFei4SQrQJa7fzy6qTA4vzykp/MjEeRZYELxGYKBDC
UkoFGTnhTHyYmoGFW0XnUg52xAYnLkxMJRyfJcp1JyJDmv74ONQXxsOG2Wn3Szbc
i1Gi/41vmc++o8C8cKlWA/5uBCMCydAxscK8QUb5z2ErN1oFAEhtToObC03dwsdU
9ECz+h4XU5c5N7LRkXZ7nhr79/My8J8ca0QYJ9nRoiofnnH3dzjte7A0LPx8MdWc
pcYQbBlAqj+Gl9yslaztYlSUryPr9pqCl1dPiMKU+10QgL8jw9COBgMVxJM5cDoD
5+uxPLixsh6COecGYYCiD4d6kIdl1pGy7kcp0PH6iEuqZZPBVvlxTBBucZ2C6E5s
Sxjya94rnJ9fTgXvBEULWBfRnsI/mdRYPBuJBRWoUd/T1ifdNcpXNugtkzbP2kHI
i/ut9dpsOgZzqPhjVKgdlQ==
`protect END_PROTECTED
