`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1bJG4POn3Fq68uT0cd33YdOe3n963ioKp0Py+3AlxMNR7nDUVN1kvWrpmWIgXbo3
gS0cvI6TTXYumPcvUWtEgVBpp4XTubB5W92katAyNz4+q3iSpZBDZIi3vK6x+dqw
UNaRTuJhO2hhSiPFgwMGVnKpMcmYMZ7DrIIEpk1mQmeQg2rdWQxrMXmxrn0zJIxb
sxSGHHCwokZMnY+UgiQplSQUT3x7th7Vda50flV5eC3P8Z1q2HmALXDhB2AfCHL3
xGU5q74EHJp8sofza2NzynxLctM28y3hvs1O1WP/59EP9yKGV+qyPNsLTROm/WyJ
5K2zep0MznTFdrGyj9Yf23a6MKXn/IW+qpzsQ+hj9rIsZr4X8GiZPNDX38tkoSfl
qxVcwkOsNTvIr25RNZF948ViqGSZ1e853FhBNi20tPFbu1C8O9lv7hfUxs0b25W/
M84aBYkvpb7SyIrZEDuTM2KY3HAO11IvjBzSajUdmkRlRd3HcfeO5ObrUqlGXB/F
mO+2czvotunxpxtfn8t7Cy3e4wYoivw5GiamhdbnZBoa7FTUivkLTKEqf7niVdmz
lYvw5ijfaSAkxR8NOaQpusyFZQqtHLLh8wAbc6C4cRHVBjAcyxkjaLtkV8X6fhq+
Ysxx5H/50wrQ4QmcJ8lLKdeAPhn3eb/FhQcoguUIry/gK9bzNeGp8Gghsw5Lmn6T
a9M73FPOqCG9PYxC7UeD2mXr1224Pmid5y85Al2wLarMJZWYIyH1w2PAYtFkZTGC
6psRndVspCHcNoiUfP25lGCcCErnRwcMsGQIYdDXZ0k/TljeEhfNQfBMQPJzRfiI
3MORBC3ADu0mDA5acgG1V+MBJxJ8TZo5NF4m++a4+cjfTOxlqXux3s2nbqrU24Xa
RD4/CYgpvdHtexGs/VeiheffPiJADkYtgn9B5bjanVi4k02An+0bKhFbkt10gaYZ
HGmnB2wEHx9+vH+lPhG3T1oD+ODmAg66ZMaAWtwNz/758ZgVgswXu8GD4Pw59ARR
z0tzCXJGa7oQRxBv7M1rUUwZZzKxS1TvGbfS0WhaRcsey7BEEvtnP3unWxHB9G1d
vareW9aZ5RNqT9UsDDcqUX/G/Azhm/EhlHX6/X1mEWU=
`protect END_PROTECTED
