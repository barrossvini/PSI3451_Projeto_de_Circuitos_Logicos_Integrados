`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MTN5SAIvgZOolmL4keic9J6WqGK4fjWuO830O89RYfL+jmwob/bqhO0/yAUbKrHH
T6XjPrkYN7Dz9HnVzEVcf7xLhHeon5bRI9coglMWoPWDC9h39xTgSXl+WdOE374Q
sypj0RyeoxUiyCDs0IvXi5+b0NmT4EpNkR4rAR4yhCHsAY2TyXWIzGmFCl9Ed4SH
/JCyWLelNvYAqwQzwSC911hovOLmsP6aWo8syf/WI9QC445Jy+lUBGq0/C4aN20a
d/VsFx4UpZfnrdADvSc/2joVjDG41G6fcxbuhQkRzHnwTYghz6Jne9aAnfSfM3lv
0QOm1cMDUvkexwk+GTpG0J+o3A/1sD1GJ8Yu33M+QZ4dzZWfjiALcg/pymMDmuEW
1czgbnPF2/8DzfY3RnPncdCyzaLkSpgyqtjU4WFgfoCCEp6rLMSQaTCmxgh6UzFP
bYUV5fQtDBZ23vuTD06wwyuTpCxwnQCPvyk9rMrMPq3qdPNpaiBqNm4FM8EpudcS
GmskIyLI/wnteGKx8pXbB4TclGdmT8sPgUUcykD7pIicF0sOVghR/RCCWCDHVO9R
t5h44XOcoTH/27irSQ7MVKnTPtt9zYt3J5M/CfGV3rQlfIED8BZlHGXvWkJZYoUp
LahXnfo3sVRCW+eIMh1TXe9p2/+2y4PZSPC9Aq+eOedeN8RdYht02Aji56Ta61qX
B9BrFKhglle4MgUHkrIvTIQfTftvYDhkdnB5LJySwYdNmnE83RdqlDXjKRy2KA2t
USY2XW5Ps3E63ZOGyfo0KjNtWtXzTdtKy5cPSVyifqMR7jPtLmgMqdLWelCIhouQ
I6+MS8DI7PaLobS1Q48zgFMvfjOzeDrv+H/YaBlkOqwgHCJ4PksxNpM9j+aisdcI
4R9l7B0PekN+QOa+OL7nA6mKN7T/jcbI9xPZ66hQ15j7uyJSHSluL9bfEIO0NoDP
mBg2eXFwShwt4/9otplAah6SrjlJPXEQSJwjI67A4KSjbwODWxHTehWBPXASzku5
CBEZDY9Qf5ESPd9HbC81l6LbIQQah5ZKeCSl2yFUsf+O1SN3K66x6tEkj9K/P09u
NBhXc6H6sYp6yV2jeZzy+xvsZ7dPpZ8b3atsPtk46eyZXTGIKbpbC8eHsY82VFiX
dX3SwlrZCP0o7O1IMzMhAI2+w9XUep88FKTt+669lZhpLVLeZauyGn4u5c4mI+7x
FZW9ruSQYci7LycOFJlGxw4GK+Yuelc3YH0v7NZQOb6HAXTjPbef9GxndOvJWeQu
vdKcr8bTfk2rfM0qJ7EdjnpFeNqRlpdQnzYQSvugnbEu/8R+dXzC06QoqG8gSQ3v
JrWdcfKwF+g0NIHPWPxFSLEf6AL52EEpvYDxb5UDsTyJ0JZqIqr6YA0luh0QBl1w
Jlv6jMG/Hg2jlYUS+8TGCPMDgUEToWuiwcblV1/XKvLv5gh5Exc77y+m3ujJjAmT
57egfQJRFpYLTVPBV4Fj2JzhemwosoB+iqD1qvd0ZGLRkUsUbX8TeB2APcUrEzNb
+vMKx0FIeTBZNm+4bOAl6M/BXnvyRdmCrCTvwHnkc/jamyDA06lWm/M46ERqXuQk
HfmQqUke+uNbzV0otL1pGgw+yWoOKavVB4jRjaJOYfuXFq1iT2ZDEx2jfiPsClnn
w8Yy+VmJvl9y0ai/e6OiMtqr7bFSVROaH2ghD6aH4BwE2bn0252w+qm86fVRKimh
jvBlOeTmkuoQQuYQTTyGL5Pum1CI/Dz/td5E4QZn6gnBIPAbhyJW8qTZLcikVHZw
MRG6cEOUq1QbFWk31YxGoZDNAMGoKAb3B6pG4xhdBsmd6FA8drfP+So0fQrt8L1d
7+Lbs+E6GnfGawIiFQIaWRLF5jBZ555+1cRaxFqGztzIfd/sKluVgkIkk9qmFiM3
x0tO4MEl6yyNj5f/FDOne/+TGz9yuGvYtzYf8c7K5dIlHbT27UxwX2Q7kLexg80s
Ud60F5AnkLUuA0i+8p3M6e/zZPo2PzSu/eel/yDqGfsSTJ0elPg1e3YBVnGb/2Ox
LvyklaERWfPXSK0GooIhqwGAJY9oQCfjcYWQH2KGr/MwdkCRJ+MPzJlVit8foiRB
r4/eK789p3dA9CjgW6WgO1jIoDHDNwpThqfYbr00O6G4x+BmB7Re5HBzQqVGOIbc
ZksW3Yg/6u3X3/PmlNU0u9LH2/Qg6WopKQGikBTr77BKDk/4BS7CnrRlvJWYnfqo
n6JnCItk2be8Fu92oTYYRaaAqcPQCzpTYKy46IJQbZ6dqRJ5K8+VUJuggulUeEtu
1p9XfnF+J+8oOizLC6delRrz07hfc3hHvbsHltjsyjk+DnrJIWhIwdZ5lMaKk1uZ
fCJpym2fRMf3rOKdGkgudx6xWTaeIveV5CppPBlFiRDvRVfYSaMuGbhzsM9ehETJ
wlHM6yWPpeYO1Im8APkOF8Pvhd/+f4+idsRmC03mgx7qOamLh5N0QbUZKzALy93A
tObfotAoz84JPYkdjr7NjHpiBmbB0utXkbfwu+dj+Q8mXUXXpW2LctC03DA+01Um
Dsxx2MhMdKWhly/xmnRQmbpFQPKbk27HfxovSfKL5vR4OYv9OZ2In6wjwZk0/b/t
vl8LYA1u996wGP14HRQo+bbgz1nAX2CTWIPKOsOXotGpGl3z5kEFLNxKTtH4DEmr
kPpZzG14z14ouweYDb1lgWi8+NgKjNLmmhGJ5LuX4LgFiUNSEUr0ez2rrnrbOyBI
gPPLfAhpHK6Skps9qgRHyyS6HZh6Uraxw3Gh69HrbUHJd5HhroL6n1xL4HJJ4LlO
LLSxDkqSxA1wSf5kEz2YRuFoW/3DvnH+hnbkhrmb2heDrGgxvU0lLo/pE2V0bHDp
e3jmJuLGv/zOMZoa3cfJ/Esbb96wd7ZGFEj0rrTMzR1yt5wcih0Rj7WeyaDnnzVo
d1S1O7eg38IOgr548cmtpU5qipkTpnu/fIve6VaHqwcIyIo8zJi3L5Efyn9+r1eq
d37nDHiCncjBEah03vPFl9XHjx4Q8B/Uhv0y3aOztSmgEhadB0u3rtB9fqYVd6TR
R4zcOXu00u4NJQDBJtVD+dUjfFQcKwA71DCYgZWnVRFPO2xWer4WYiPsKUbL8urT
uDEEbJy/FLmpJOTzwhmIX59KGVfAb4ilhmlOVvJ0zn0b5o4A3mjQFqL/k56w1sXJ
0LPcaTDVL67iN+koemrDZdtjr/G7GQu8J039P/OeQXc0q+a4693ikUTCerbMmjOX
teV/q1DpbxwJ3bl7DkyKjIS7pIg4MSZ+H0skTN2CMbsiD1hynRcNeHwvVzrNT6ha
j9u7SQoMkqnTEn4r3zgIlq5ZIo3JulIVFqtcoF3FDQTMRFhUSPytveECXUR7u1wd
KesnqHx6Y11lPRoN2A3cxTzRqAeVUu7QrMnfDlV8sChGIDWPcLVZjdlXAce58NCs
iWGiGLX3DpGBQj5ObmiYbt5RhugzSGw+RewmPeKNn+a6aKHcKGw8AXGl+Vum9ggC
iGTu+hy3oR+DyBlHyV7e3M+jPNSGLflNInr1EjpHMfGHTbnkVuuKOWowf97sPfj9
d6yenFzoUEN1r2VEa0CgFQ0PDvXXggJ7LSR9iG4nV70HCVZTi/dBRNvqicOXfC/C
re+B+AuqKCh1UysDZAh3mKaQNAIWZeVmI78faqmcTs0857F8sI3QczVmiTQhJUeI
lPE+McVO+STjCvNjEcmkbUnpNEHvh2GWcFtZmf+2ukNUhTmb/kjFWRLOM/3XcM5t
Vjh6Q63FDxVUwtskXWnrXBYEVbOEZBkMeONgIoWHWYBazkKsixo7M8F9jZ4wEP8+
zoIqkJWdjjSVVQXeZUY9x8pvsxjirCwRI7WSN4jso5K2esISjtTGY1qW2TbrKXbb
eDUEX/0KPPt/sv/bOs0ihABW92NY23PVIoc5nD9euHEsFWPcdg4hXX775d/RTRSa
YFqlHZIaEUAbJ2y2etswbvrQKtxwmGpT/wI/FsEkry7b9DHpxEd4vgCRlY278/Vd
WDWLh+FYNnBQmTqP0FxNLYcGVvvYHaZO2mbRJuexyDdd7raYvyWtSepjbSrj/3LP
/QKuhfeaIXqM1wQHslVWk/4nUKlL1CYOFEQbYc4wYdBDHXUz1VqmGpYHZG7vQgB0
fBBJtjiqJZqkLIopg0niTrciFaj7JG2Fl+5BHSCDIuAYOtIioMYKyNR1klabnXaG
+DxNZehtrxEXhv6jPMQK8gyg9T9TA02HruNqCKYSKhz0ycvFGLdXEoFKgV6ZBjlk
wZ3J8yUQSG5zjfRk3uLYJrTiLEdP/jMUEeI0tN9Kow31uWGZfXz9XjAucNSPRzG/
j4mkTjgECGGho2q35sJThJ4t5+IhrJTeDUC20BeIiPt4DsHh6lkrWftAiyYAiHSn
4KWOVJrH67AvLre45xD8wNQOvYVpaIlNbtn+ot0STWH2Rw4pXK/tKx0T0HczB4Xn
3LYvLCcY1U3fTUbnuPBSXnzOMLlXtB3WgjR9AmI0CsAQTa+QlwNPj4peeKv1Lyja
r7zIJACuiTq0rRyg1xrQ86KfVZo3e/JL76pFG87L7s12kPXF8Ktm7/f36BIiRs98
zx1OmxaUsh6asw9h7VATM3Hv8WxGjAn+4h6or1Zw5Gr+dzLo6Wgj49jppOGI/Gy+
fScnauPEGKanWPHknE9JTvnk3o8w5oQaPn3qaPjatl4HYlbafA/4HjbHXFHlaXWZ
o53RWWx0ihscEPWSK5XLF0Tn8TPsOdCFouMyV3SmBHUEmw2kibwERAyxoSwFO7Y1
XiuvJXpKq/wHS17BAFQTBd0nn3rSCMRrZ+5ImP7AReVwafL4/x+Qb+nVBJrqCfZX
exGmfCcT/e15ECK72AWTI+7pg5mVDPqz8sl6Zkz20ZkujJd/PB70xxVbe+hdbcW0
s0yoz6FD+GARkgYT1eLCrRdKRDvgWpKO03ivDvtza5oYibaK5X5xNY78kXZmLV2I
+EPt58SP1M6w8D+VYMwT45PpBoJPYfoLqJ7tEsr9gLD5fZX0FDP+cD0CX//iwaFb
iA7yAMhHGdC7PbXWEIPvF9F2Zvl+obePWX3FtoqMlWdxDHofIC2pXfjbHJreYtaB
eHD7ijqLJE1CITQL0roVGD9k42vANXR4EEP7LwhxHbeHuVpBAOGTBCv93c4bo08X
r2uFj2YS9GRDIUL0wnD5lThNKnNgnkW6nZEAbw22gvum61XHu9E8cp7Mv9BKTTZh
7wg8k8+nhcQBpYDLL1fPuKefsUU5gnUTM+4DUVuG7HwVPO1wfcdNu852zMf8Vxkd
GxbUZDgOm1R0FwZf3kjq/Bo7e3hM3sSECxZ0HRk3Kh8fEmIL4pJ5q3d7byYVT7yf
YOxW3esVmFgX7p6ezxFOsI0GABPvgiqU4LjixDZHT+AM143fLbAR0hPOtgKSDSmi
xNv7Jm+ca+K/+5pFUoH7okCJcwQSB2zwoCn7tMVtlDT7rQE9CUL6vDJLJ9LWGc8Y
qze6rSSvPsIBaJW/IHC07xg3P6qDKnDKE+LW0bXJ5EhmKARBU5jYFUcan543U4gf
qbt338J2TJm0nuGpuhHykq3El+uMwtIy5ZjpavUHSuYHKufvizp9PYOVU+s02wwK
pH9k3tX3EW/VFlw50NnGHEsZNHAX3b2LqCC4Kx/sLDK5oYkk0OR5wRcQ/nIZ84nH
ortDIL7ZnGWY9TFLGIqwCeCxFOsIcZmVrAjRR3rCiNblWhYLCPeqwDKNtI1Sxk9C
ETaQNfiOAS2vL+X6IaC2LNVxeea/ei3bhD9f0JIRXbygMO+D5tzFm9MdTR6xymOG
kRO0HurvcRV0tiVq24/tW6c4ndkGqpdOwsFUSRTlPIgX+1rghZEzZci0JhrkZ84m
eGZAuo1WuZBk5k7VSfu5dSXlLZED1IjbhgcX86BwGFYzUFXUzBbTulkhCPBApy1x
Ls8IWOqla+SZa0e/lBMBDy5p1v6BUE6FXbG8k16GIJ3VCbmmWXtlbWpe42ls9yhe
E76Pqshvqx3Kfu4ETLKDFfLI5EVjJtCThFJp6GOh+YAXlcKWxXIA/2Frn/K7iHwK
IUjFY4iGMjkgMacsD6p9fdpbg6710GuWYsTn+SpIJDmnH+g7beYC8C3QL2iC3RqC
Mvpbeu9xDxY5tLMFX3XVgcjzb7kVsFgbeeaWlwNMTHBMsrCo6yWyxYrDM5eXGQc+
jKT/axYplHDyLK86/p4xGJgxD35r2Mr/N4Y09HLJgmH+gn6OX1/BOALq9KC3GbXn
E6Q/GlLsYPDnvl7D6n/ymoQlsmrDex52Vq+ib7LSuDE0+Xwo+ARZ8yuK6NVMEeLZ
74M1848NL9HZHQDggxFwymuTCq9k9ptr5v93OA7IIp2GlzYs/p/xQpT7ArDcAnMR
NOyT5cHjS9biKzVec0vB7OoO1+33eGSbo0j515zXzdHX39gweFjueiJlD6yDIwz7
77y6hSeq/CbuUc3nvNnyF9KbIvgMRodpwR4XBDrqyaYk/jPjT5vny9U8p2yKrij2
FAY5G15wTwgjEKfu0MISn1Z0W6WpMAjIYxIOcZkIAGPaqroj9cUGAhuHnW7K5Svr
0sSOPyx+06+WTEnqX35qzmvZH9tdDMdO4JazE72wMZLvjS1hp5NgkAMsxSVrWS4K
nVWFImedyYsnzfc72CkGMim2JC1OBPgjX6sHEhzsR11su6LxOqnqH45hl7MH/qbT
F9xyUGf6e6ifRP8YOmZI9Z8QOVXYl68ueLj4xxazOpw=
`protect END_PROTECTED
