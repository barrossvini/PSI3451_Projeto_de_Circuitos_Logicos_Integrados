`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
knxZDiBsbzxYrY97O/x5kW8RiYy6gKicqbemckRnlzMcWVrukZrB9KZrSO0CNYj1
YNYMzyBGYWZTep3m92SwoiKEHju7xiU8nlw8wOr5ddDZxY1kviibgyYN4nM58l36
L88q3gO4cPeJ3zS14QyCs0yNLz53m8sNvlqcgKhAI09vZGdxMMyD21L0xig+Up9O
H5vkyhq0xLwUQM/FluEXwrNkBwrHf+P3WxkACLICxSVfRT6+/Wh6Vr/670/SuBw8
T+n9VcNYmUWM8SZHoDoqxQ==
`protect END_PROTECTED
