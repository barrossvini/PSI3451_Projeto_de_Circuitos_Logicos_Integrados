`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYr6GTjE9lgBDLirUu7JWR/IgHcWM6rWU6ap2dOQaM+zI5/OFcb5pTAGk6ELfCFy
yx+igvNEDrJO96Jw4Gca3HkNDQ+bCvdD+rwbcCymmqGRZtw+i3mOjTgd0xwAnBDF
HI3R89oNn6s5ALzGkol76l0mYftdwtqaHRlPnzMGG9BQA1/vt0wboGYljhT4dvOW
VFeXh5BekfDkeKjBwuJJOmjfm8rOl5N7OAb1Voz5Gnjw610KIE21HEqlmZ+N1dkI
LQQhMycB13wQWD/DFFO00zFnAjzEsDiHSy6QnrhOQp4hu+xy8aSTnaFn8Vk5syhk
3b9XTVigv7Rsw/ahngGNV8m7XrpdYAJGzOqtfn6+xg9WUcqJd9I+8ZLUD8w5NYo6
ZT2D56Lraa3R4KLK2wtvFlxu8AWhsyEduG2i8NvNTiWLyOYttKCwLAQb1Clt2xMH
UG8VMQNhssf0TCksmShbjCn7xd2QDN4I0fAYFfbmWb8nqTo/1CSY2T/w2rqh4DFY
LXVJE9mL+zzNdgI32tQBfoPFiZfYvIflUsWV2Ftn5Ueih3rA4YNZMRTab3HqfIXw
ODsb5y/YVMa7A8i1N+osbBAuKxG1l+7Nn+z9gdT8supbASFlgs/i/mxdwG9Fy7CF
Mcre1MlTQtbZvKFH+8QhaJz8k7xokxdEvhVCfzB0NGT2NfednFXklkJ0wrjtoymr
qpFOoswhJBlHNt6fdkgSg5t/qDxhbXWDQWTkOxcXsBGU7v5dNAa7thFkOj+LL1gC
wfR4pY6iqfn3g2jvDVgmvbPQhKEE9PEJ1m3a2tLjdfdsOWUUnT9SJZnKWFKUmW8o
j4Z8DtkgXGlxNaOS8xQcM41LgLxS+EZKrKrxfhqCwc1alKzDeOInCKFNanrKleZs
/p+WymhrEu5pkuLzKfP8w12of+w9bUAingiUEXA5ezHEMjLNwXEs5HJSGjTvBNr7
/sTw7m5oZMRNBfpBDyLZqg8Hh4HeZsjEXVomsQ95dwkID17CbLxak979ntJ0zHG4
V7uzoR/GlgfbyS7qSvICs5NFSBIS8Oo/I0SI8/cE7nGCo4FDYpN4p2rNxAW8yHGG
1mGXvR3JdOrQ/tBgrk6TmqoaFCGhl8uhWTTR41TH+H7MkVB7ZDubGAlOXhWwaq3A
MQq3P04LlI6PfcW3yTksFQrXJS8DGjTjZPh2bXmMOqq1ulQTzavQGZj4yC6EB2nG
rN4h9H4L7eIOXRJ5Wkggyw7Ph8l5ChOSoUsgMnX4pDPip3l13mvdv3hOLJqXlEu2
NpYN4W0r6mwF3mEOVvH+ryp71g2k+Smci3e5wKo/Gv0F5Ahu5+RVedUBTN6kRHZe
gZJ1fVJoRdcuxCvrRLI3oqHIKmS4Q0mHptbK+Y8o1/hYbOrl6pBBTUjT8oH4U3L2
l4MSIsYdkbCUdRAiXDAOnV/1C6WqpsTay3adX6jlvjU=
`protect END_PROTECTED
