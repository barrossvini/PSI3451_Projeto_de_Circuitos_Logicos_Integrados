`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gJmoSSti6Eq+8fBvF6rwjUILE3Kv0u8QeEsnc7dfw+6xPqZCLD0R7/5W07WtYwBo
YXDQ+zWum5o+Sl3CLZ56g1bfbWxW5Hz4IJhyAQbRq1m6bCH2c1MhKCenTm4+5+xj
WzGfOxqunOSSUOIpPKWXsP+0NmLrqmnqda1zqDV+MMElUFYcj/DQzJ9qWtdF9Dnk
9lulJutJiJGLpsSOjC2OesHJyFnZKmjlnBgvKi3gKuuJJ9SBEruXR0cp7OJQGWwo
WP1HT6RKBFWZMNLujd7EYN98lb4OGOUUYwFfJx5j4vo/7pbzx+r0MxSP4syZgp+F
IrD9pvRjy8JGsUfjD1pVJffSRrYQFDv8sV2YMz1UpfjNDKxn2xnThygYhWhcvTv1
D1FSvNNmQSfpuB6+i3M3K27beTFauawJ9th18UZh10jG9/vSGtZmw8xtnVKz6qsF
Nkrme96sc7PJvIVQNSAg7C94+t9SM8N9vz/ZtexZYZX0gv2mxOW3JTsDdpIf/nCn
8DDjbyirHk5AUmW2UHxX7uDsrbG39nlfYzJTOgnNRfPxkFkmjS8QbaYm6IWWQTaY
GSuRI1D/Kk2w1BmBD4POWXJA8KsnryxU0U3Ta7LB4elwoyASmnJpr5vc8FNhtF5j
8je2tE1vLfqLeEZhwAkPL7iZJkuu8o6R8mMvxdrzmpidWy9NKCNU3tsBEN0ONY0u
`protect END_PROTECTED
