`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hYUKuAPXwvWUaJnUDapzSv5UxlFFsDYvpum25R1SfFCFHY6w1XU9q/f6D3Pel1FM
OaCDvq1lXkPnCccghYKups/ZmOPaFyxf7Duwqf380WgcV8y+w6u/BqEJ9QdgYQY1
j6PiQWOJEtNIF5IeBRwToUivA5BQ+57TF/fRyEf16dMfPGMxN0W6bA0N17qXzSEr
lnUOrEd+RSiARTim7Z9ljvauFXZQuiwOCzwR2F2rtGOIKpUbTPRBOwtZzlbU4kXd
gHLzDr5C0A/lNxDQBPCMWuQ6GO35TRh3VB70QL0i/Vgl1ITjcsyNrW62r8DY39dd
clLiH/y2vcUqdXJ7+7PJReNihy1XoBSn1g4gCuJUpUIQ55Vm5el1p7WRKqcXuCkp
ZCvHgKvIfOHYTadu+MdCfsnXjjcMWZa2cRLxsaNYh21iTL5ZwX/HRwgXJWhf98V5
6VSyNIUWLDk3nPhPIpT7PnCzHf40M/S0AjyVOGNZYm9wi5mDtObuhjvZm9tT17JO
beVFFR+O6FyJTuHmch81kiiMVMmG/gv7J5OYPMv+kUh/19pBLeq7o/161SaWpDCK
XiXb0tpUthF5em6bUzMmSxIRnbO7kKyefXbA6ayETtNWRLkoLGYJKkSahRagcsVE
OQNOjIi3UpZetHwwTARFCe8RftimHvW2tpCeYT9ErHUjuVMoyKBAdH6kUmxGFzQv
GpPoKGLuTle1lUxLOiNRBQWHgQwQlGs8n5I6dH4bNgus9nAdg8jbyAA1NTXZoAui
TTeGxR2faoSXd2lHCgWg6U5BolmcKb9GVq7d4fHvECrZws40XKOA31EG0k9BRrWB
rkhklsIDX1t7YEJzgwvUvbjDiHR6AT6lTrttwaj8x2F1v9Qns/Fx1Ex3eVhHwI/K
Ph96bk3/J0kBuuBgT7p5RaL6XYyvhJ+LnfHZ0ILAqsDZ/FVLWynpj3jvFf6cYTyW
e5VsrzgGJUUnqLXihBGUvSngelECJqrW6rugFlk2JTyvHO9/rMblVyZ7ceYUomtX
zHoJuSW0aMEczfEpZYnTPhU03OQFKhHOoHP++qAD8KeKvu692TuKWjtoJ3sFhdeL
ODdhuts/z7BkfVS3LvLNc3RzIyDzKQFEw+dk3uGxdNdCKk89a1F9RZQWEc6QPbjP
T9Kz3A1Wc1jlNW/8m+u8xFtQ0OqlV56db3RHssw9MFwsfhtKnyyPehwiCT1fqzNE
Ico6YSv4cjC+t4BCmEvjiBeZdYG0NXTeOZeQpa0vmSianIYpQKvApmLky5lVHb8T
toikbzsHLrvtjb9PgBNojLLCYOCHOqkRfldvSCiMUv/dmHiHZDEONW9pIJ8GVG/K
/dH+biAAu49tEtrF77aAyTV9yFLJ0pi2tbIZiKUJMDYxjRmIMCz7TkGwtfz5eSqU
2FZhUHaYcfsNcZePmHfrY7aH5rV/SMJ3TZGmbb/RgkJBbuUBXv1/fVX0vejJriOd
AqI/KSvRl4d++gQM1wl6k6bpBKgxTwkBmvGVEyawKKLdEF1iJsL9zxsuD7QZRxYp
ATH/wsmoZCkulh9+NNwhJVvDLsNROoafG6l4P74Qtt+HYbnKZmihCs9J10zuTBPb
NiZIVBiEKYgfL2mO0avuUqaa+XbGXkgRvlzyAmhg7/SCXlwFzOeULkg4grj1tdZo
Du4xIgxT/iJMGjrzpNribV4yCNFY68Fgek4CsWVJGyCIM0Kc5qJk22yodNhvcGkS
mnDA9tL0vz7fzU6XS/o0kDfmN0ghOzquQs0KnQvWs+JfSMCBThxFd1ofR2n6Mj26
T7Y1xzU0PF0a0cjxJrCZImpKeueUgJljFolIksWYq6WJHSbUr67njSa9kTY7Y/Zu
5SL0A1pE6HfXQfsXrQuqu+ybpzCfofouRu7PObqXfIiynTV5NQBRV2HTBx8TpiaU
VrCIq1bo79ONH5L/KinT7max65dJE4MIO1NXZCw9ilJFH0pmn+UfImXZ90ypI42g
kvC49rWwt6/OGvmNsp/3uHzcVo4H/fsS6DwBhLdvGlGoR4WUeAZnonDqHx718/vA
upBhpsSucZsKpsuyOw1Hpw4T5s4e00HXzSsOzWmllw1YanY7a7s3cfz6JALIWzmZ
nXKFqxGj4wHUOBUdJ4APdWq/USllod7u5YpnHM6DlnZ8rxrmHcdrga0C9NPwjrHk
yR0zGBo4E0QnHheNotm36Rp2fr8M2zG0Ak80F7OYQS5lX5L0O/rGfhMYJsZ9C4Q3
CQsZcEg4ycxLDZ8BuaITgAS3mpbYASskP/8P7nGbRAyIG1Oqrz0MUCQ9znxOnnxC
WJyekUhWXE6LQ9rOjF45iYh1+gfeuKPegrD4zamovnx9Xtv0yh/LBOqVPeiMyULd
naOvcE5uEW76AJ9jUemDre0PvlPB89D9p9S+AKtsbit6ltz+Jrh8zx2hymxTsQDS
6SdJyHX67dciPaRGXHxkd1pTJzAA0TZUAhqM+z4t/wLtr57Kcr/7A/ivJYvFfx+i
UvXoSe11m/QQXsusuatnk6by8tO7klgWfXnpOkoFm/7Yo2MBMy2HYyURUBOipbcw
YVRAXgDG9s+e+lUFhkHAHAs5rXDnHJHWUn/X9ttlQ/GRyMOtBFNMWPEhE72nGqEa
WNlsl9Rj2bmxliHeZSVFsmUJscwK6XV5NSZIpZkMdLmlg4RPyhxKa+VwKtGkpaLZ
675fCcYRZRgtYf4PEiOqZnzJ2DVypGBS8V2AI9nJGDT5ZiYn8BBWJAnDdMWCW+ov
XXZ1H004DveCp/SkfigV0hHaamaqvpv4+ZgB63k4ME3//os52qN+C/YzLN8ZvV/O
U9bY3cELiGWTPzsuEoRILM/3qBIdN8qef4l5HZwbNZOdOorRfjbH9tO+yU4hrkaZ
UXibZxcesIHujB1g0o2AQh2Z7Z9122zCM7prSglwxEJCT83Jhcs0GVh6pPAK5XZm
PySTYMwr7BC41UOEFbdnxLLku7Up2leM8WjUpzNEmDgnjLmiStE+rLmgLJ6LIEGP
gpz5cHdiGfsUrlR5K7de7u7IkbvjE/Mpjc1zYXk/SO7pjhxpFtUwgv7YhY+CKLpx
DHesI/CcDB499YooSP4eTJJOquDgswUt9LSUSwAsM22H8oA6LhrMhHBDn7/Y8baM
MhLRqFfEb3OPh+RfxFgJxRU80AA4/QjMh/Gx9l1Gyd9mojKyGOhkxU8Y9muJfgjw
Dqn6ha+syOEOfKS+pThe6qmrfaUcNr/U2FJB9oM0FCXvAiY4HHZOwUJ2YN5Tu2Wr
SLdKz7BCKIIa1NiN+z5418K0ihTlO3YF+1uEmutHrvtBJJDzabTcotbD14eH/wVN
NDHgndHARJYe808v06H1bV+woKuPSVv09ZOGOqDMgp+HTJ0EuDqb3LGKk54yxGST
QtgAUPnXdzA3aBd6oEsTCK9jlDloVWQIP4mEz9c2M8jX9iO0zOC6SYYsoLDuurvT
GloXYEwRp0XGYTIyoOi5+uFqVudyEVpC8LB1d6gfuTSYHdp+/P2V3dQgNOmLEjAI
GCDl6GTby+u0sDkavedKLbLNRTWBMuIuqmyhBQ1Y7Sr+SqHzuf5iSVPL/9ZPZsLX
78mOa3oPTdDgZ5EI9tak6u7ZsrokTehi0BQjyebwCrHOfWF1zXoETcqBW5R7TK4D
baTElCiir8q9mrVz8W1a5z81/KKcbOY3KHaD6iWFQB0fZphZrUyaILpz8DUm9Zq1
IG6rZQvWLwzNLPXkpe+7CvW57EQxJI+rwiEuKSuV4k8nTzVB8BS+Y/0dQ2+CXvKV
Ap8QYv7iFmwItqMLbm0HWcj5FhISilxVlF03fYe3CnBwEqLw9xqxe42dPb1cnDf0
xMhG7WGotYGv5j2Yo1mmWCfT3j2k3SeCmHWCC4Q5hH3P2KfRBhvGHl0E7PhxtZic
00wrcOrXNIx7MvZ4hKtuayHoYvQSwqlOnqPRDoOpZANMILE3Xc1a8Nhe7QWEyz5/
w7zO6ecqASBCrx0EFhzfItbdwjTa654J32Jb9JijFtW94Jea+Ab1NuzVus7QkQS/
u7xWZHwfGEBcP3w7SFpRYtjj49ByQH+k3S1e72mAZiUWYW+SYfm+ai/0uSQ3VqVh
PXUskYvGki93zLN3gVR+NIwA8J8kzjVL81LWV3dvrEhvSBJAv0W1gV4L09iH/sKo
Q0IU7TWa5QxXn5OYYIgYaFbum3qhvKm+Yo39YCpIV91nl9P292EIh0NHfCep251j
9X6V0GYy6gizyitnaG/WOuYV35fjCC+Z1B3xsONdB4GX805GgoKS3qdKaNDBfQy6
VaQIAY9Ce5rmRjFOpvSiLgNEYJso6mv9deL4X61ufKSLOWB2FzrwDE2EukXg86xy
0RWriCVo03RJe4r63X8ZJWEmVEU+rJ5R2mduvF2oWdKaKVQsL+Lqf+b1cGYcUGyM
BcIlXXedp3foo/CGgi5T+zf2asRP13N0OYT94NqOCYW9LuDr1lpE+jgKrLjI2inR
ZXaBLBWCBsuj6mUPT7BFZMFDwohO5/hAKyYF1EuiiSwfy4qYjam/6KBwaTjf7KV3
HVJsOxxLO27/DXDuH0eCw1SoeI7palSVVMtbsZUOHFFuXUNQmxDY7hvGaaZcA/Fc
DSz56xcaNMrnpy9fhAoAnYrkc5P7KeTGBokwafSugvOXJM3DtQAW6K1ovITVejDf
UcGZHOsWkTLezJjStzLeoScACv47WkUxKgMiOxwW0aVj00N/eWyDky1BJDra+3yP
nOQUrQ149yx5sUHXdpOPjsP3V5gTJXrTf6Waux4VkD+M/u1aNYAsBCnqHzyghrrQ
5aJVfmNBRHsK8UC9ayyXzxcJJEiRNnvV3TFtqCgXhMDS443YXD2o3qg3xZQs70ic
U1+0i8w8LElFsJ3itdCw4ECaY38MoO65wXEduHyqw6ea/FmFLDZ4yUcfly6N93gX
ykVuPc9Ntc4QwX6ZmuHgsCEQkoHG1pPyIWxj/DFN79Ulig1wIANqBJUhEA4UZv9v
GotZCnr4/Zs3G4mRd/TQUYaNCX4jibM75/1nWeiVWippEeGENPsNjTG1YJhDtJCK
eNKSDOAbg2Difxb61RWk5BZ4Vc8lnY91KhkCMs+UoohHoPxOPJFAvpkED/gC5b3q
cZFHmOtOUujgz3yz6weYFlGo0GNkPR90cewSukmsKayKkm2Es1WsJK4+7oZuefaI
3PyXBfhNWLYm2Mz964gAom755GFCct13pNXFbnbdfPMLbe/5/RO9co9eLXk4FVH5
CImjMlu3OMN0IpkXtTPBopApzt37yGOJe+4zQDS208xLMfXQ4AuIJZPcYLI6ETPU
yAFr3gPuzFqRbSEvOYXAlxJmaaz0FJeBFo/PmhnOKKimRg1xCB1eUUAe3w+m6yIc
ATxwJKihB4NkrSY3MSiGof9f3QFIjy3auTYrnt5wdRrhJ8iWC8fXX+Xfr6NP1ATG
TOAEOSIwyo583Be85iJXvZUjXLXl5i5mQJlrQHVq+na3OclHWqKB/vENefhuq0vb
Fr+PAZl6RBsJeiAi0zzMYGcEydebDavAcTBFKKJQtGuHS+/LdgBtOop8zpk7Wdx6
hXUG8CGlOiovBxRTih81eyPu9SVtco/V1MWLv92X3JZ/qdn6WIubCvMTxvkab7MD
Er/TjUoeXbNFBKB1+EmbyUDB6gUEt4HAZam+1dwTx7NNkgpMlc+v+czubtXHdtQ0
exTlod4mjVeHUEjuDMet672qpwltp8U6amf+5fHnbd4nxqz8xbrLfWwc24aYt2oP
WihxQVgzLn9+Dw1065pwW5Hbj2L2JYAPUq/afiPpCHm4yyhmIdkGYBvON7crsqD6
2q2hBK3fTOPmtibt3VOIurA4bkFBh0jctogGtyBAasJFSAFhQpEEE4tutAeK6ZdI
ScH7J3vxznzivzPcYuNoALZNv1Izixv1KDGlsHAu2z5L9UGKQgS1b27mo7NiHqZb
bA6jwvXSv+6yzavS7bDM4qhiwjN9KGdRam/FQV+Qw348E1qlw1JujxIGGJEeFrkk
TAeqB7Vef7zEsLCyQH9anLD8Gd24AEnn9BO0kK7Cow8jPL/q8buTv6ME2T9FbJjv
qgidoJkHdIJZndM6KcPW3FPzOh7qdmeeU05mBRSZdiLMB8SLjVnn1JGdSH8kmeZC
BsCVJ4pjDK2F9jhGI9o+AgMf3cUdUuqUhIawgC+qXyuvHQ09/kEyf94or+KxfRcC
kJ5tiI/bSSJN39BUkcUbWqcuOhnDOne6yA5SAIpv7JlgZ/Bv+DlPRM5wU5tpGuOO
Q0I2ZC+WUPP4rJFLnZo5A5QN5xmn3aGyWTkc7mEIMBoqwZRaAiBvkcFPAXaqYd7y
xM5RfMblpeaeig0orMyB41E3uNetFwaw8huVjbQqYwJB6iuzPoAAfdkDreZ/86Sp
VLHnpzLB6kr8cr8jgJwv0iiyblbI4By2LoHLwcdazIYTMJhpbJFyEjoaZ1Tc7Vxa
Z7YDjCRJ78LK1yF1nzswQ87dulyJyfRr8EP68A4CeZw26MBajnb+cvcDfSNd7eAx
Ct1e3p2Tv0YoZ7xr+9ya+p1GQya0+w3usPnjHBrpsFWBQhTMrN9CFZGRvB99IkIk
dpgI+HFBk+CQ/cOigSgAIk17r7MBdVIog9G6ztlVygbT+Vc2AO/SsXQHJe1xLh5N
2FsUov32A1H/L6CWZsGRNikkcy2IPB8nStO0ZM9ElH2MRWtttQM8F4tyzbsvOC9u
6ejj07r5MOAxpVsG1uKAjMqWndldlDc54dbXZyTO00I//gAe0W+GqOXoAbLW39gc
3o6FYsxqtEDF6Q50o4oA/sSPvWlaf9785kUDTpOGtyetGX5RUy/jF5JiG4V1eoEa
hxHurJf30zcD19K6vNQDaPyPhDFajn9WIMvvRLVnc8uXSxaRDp+oBJ1y+1erKwoY
BLF+HvXIT62ZYmMSGYy6K4e2NG9k/xZAHVURpGyeqL7J+U92pCEUnfRHscIRke4Z
0/v2QRi0iBJyua6hs0nSs2R0md6kKVYBxEEwk5VdrMPeCRH3FCy0q9uTBNcOkDvI
ZdbCDxkkZGOk/kIM2qYKoXEUfb8L/MkjhsUtEoAHjNn3SMJ9P4+cnGjNx/aN4zY4
pKy8/N5f6p/TTY4HcBFnMgts/qq0oMRfZWWcZJfnH0dMEc4izyiTDb66VkfaVCWG
jCU2XPiNClYswxfgY2UPw11M6s/ZRQMDwYXAai+FXyiV3wYTUmJVbzJwuGu3p3Ue
HFK8efyF6Ngu3Q6y4s5ZrTeIOMAcdj9nzzJvx5X9ESsoq1lF7I5fzk+urS215nR7
J61Uxs8wjTS6inVIGmVl4OFNaki73HgkJASWxI1tkX72+INPINNzDqJntDZGlrfK
IBp+cuO9L97zwZwBh59nMtRCrTiGRmasD9EKuFWV4ElDyifcCELF/6GXZF0382bS
ymQ0f3+zSnh6eNNFI2xeCM0wrG2QZhKsXhtx6rrDGkIOTLb7lYWouC89YVhHn6dd
2D408lxfEVVHvtlsz/+YgGBMIFvDxOhq9oNu0Zh3RCeyglkOc0kNkkk09ySREy3k
+bAsD9+TGbZPcGVwpfQAecBhDxvOeqCI9kAjSSpNKhjsgwvpT6Gaw6mBH+p4o5YU
4gd3Ao6dns6GZwYPTpBNCvXamtiK2uw8G8Tn0O6HP6Mh2/d15RN0thw85Lrs5u8v
+NH1lA7twp7N+qpnGnB/jKC2094R2llcYVX96jdPsoj/Op330zTAbzy1NRTYKkLJ
bGQdw7+ey1EOOfDuIuv2xF5PU8XtkfJaNAMs3tw0Q+OI8Qo7au+RQJ6P1k1BFkZw
b+UScb/QERmVxbnz/z1RFKIvNxV2qwFciQQftqyI3Lb4t0pKvSzF9Gcw2kG25GMb
/jPFInwc3DM+n+PabSs9Uej/aFYD6QZhFsodqBlN2oRy3QAIcPOz5TcDvVibjUHO
aXLk6pCIpUZIdxzNGEGT3DYudjcEu1ZI+MTVd9lFGtdvP+sSXstmHQeq7aEZfSE+
4gJ4xuqdwTQC/dvB8Rh/gOJfj6zk7roePiwCSuCK92OVAIRHrNTXObCGe7X007HB
wrqpcprr1Xl2uf7s9Qr2BeQohIjgWPj+Q2N6q5c7jgwkcd/dc7SH44d9ROdEjfOp
bBNdDbLBQ6Jhy0LrLcQyZ8rn1TJ+QL66lD/cZ444JzTZV21xHJmlcWP6CoiT5TGt
Pnh9zWnhHSL8hHA/KWa+AHKzWmIol3DgLhMIhyPx/kggMp/8FDXGJfLW+1rD8UkP
9SpPuJAEwwySbkd6ofM2+vli3flCh4Y1bX+qRYwfyWJcj/sO6oNjfUj7DktSHPn9
RquYgDKkuCYAIaYXSqmd5jEBQSNoGmMxh9ne2nE/v0bB0rrofZbBLmRtuG22BvA2
2HJgdo/zTeocynrv80T8gHPFoQ3F9c5AMbCgmyrKB2f+qqICpilVfJPMleXJDb3W
Ry2+MgYGQ73VpWBm2qwsVyx0wsOll/01jV2G24qHKqmnYpsXNW/v8xwAM66oaIRi
+1p6vJlisCsSWorkvlDPJn5YlawB1jZ9sCre64tvriUJwpOx/+rBvETIy1E5ee2/
4H7jXppmUX5nraddVfh8/CMM5WsDCHOruBeB6tMYhSVXMH3gbvHbxhsGF5NGpUJd
o0DBfXfeP242HxIWnWG970PJStf+ml0uerRIAHLH3SI9Ny9TMgWEQn9aDGHG0PLd
A9WvFhoOF3LFEGl5dTkRX/YChs///2PBvtQycCtYUUBoalLd7aiPN00RzEtZHOcj
SbhDSlcVs5ADbo6jXA8YG0Fmadc43M6Vgy/PlT3yl7d14f65OH8e2m4Qk35iiX/W
7vv+Uq318DTW2zCtEZeankhZYHYkqKplS2hc5ujqdVojj2MJKsdw+S2VApb9oWcF
0yOaVQl5UClqADPEC6W5kEUCaQ5C9ehSc0YbXmaeMat9kDvY5Rxss0prLPPUO2wz
6wEjEUkombqWVC8emmhHxCVG2EoiiDsLSsUOvq2QyOEUBlzUlVNZXL/0KbeEZNrA
xUBzlo6r21IWTaAEUMLQFXb8ZGo8bQ3OdrLLL9VcN9iZ+pAn4Z51tfDsBQaVIM4M
P/kWdYEOTDMkeCEx5HiEyUZ+fkgGMpQJxu6Cc60Dd/n3fyipMeC0PN803Mm2JoKb
+MtwuqDfGFs12dYcejQ+vP4bZiCcBQXf+B7xVrhZBp10DgUuP/oSvWByQLQgK5TX
/zwsk1oEJ4w41wRIyJHPt0Hn446NHU3nXEPpXLc71aESXPLHKm7j8rFW/c4FKcBt
xfAk6a8LsLR/GOFQurPD4x6OMQqI5rOmLXzNb1Ch/cRwyltra4SUq5WWtMgmIbfV
QTcCPuK1i97Mq1XJgo912ysFDhnb5VfxzCLZP7q9Q5c5MZrU4Z8v/0tYsQ5c8I04
mnBrnY2a0MarQfFTY3k+XirkzSs8DLYFDzR1hm34/ez8Ig9eUjR4tsfVMrXLuDky
BVnc72067DCxzf3agtanc6mGeCPs3xFip2DOmiqRSAsLfBUW0HqfUgw6Ny/tDk4B
hPFd48nlyURjwrlR8arJEwMIh61nHMEJOlBDMW/U6PMhbLV+nSuN/ZSOjCui9t3w
2ZEDyNedlwG/kz+A9ZfiD6ZgIE4GbSH8Oh3c/BSHJilDfCZPNgNR6OxPwybG0ZpS
xvsJB469woPF5NAkjwRt8KQo14oJ8xec8F3JvCJmvM976VPBTDPzHv+yGHWYEI/5
s208bVdQexwf91GJ8ASuzEUEDffRloeB/7jjItvotsn59oVH7YvORXg0kt6cYtg4
4jaEjOUiv06cCbtOcmWAXmp7HQAFmBOhkk+0AqKZlu50dSHdIUpHe8ecL4mKkylP
JWfg97m9JDy2W7JZfqDg+PXcT7Ix7ByrH5dRdQz4uxIZD/PB/QepuP8lwDnO8Z+i
zJqqO/K/p0MHRi5Y0s3QcX0j5CtuTIYWtW0SMylwjNik1aAZCUDmJ9w/750RhUHs
eoIcDbJbLLaGzd5Er/vNdCuNbav9wnbce4LHbEejVD2y9vQxqM32+0HEr8nQd3L1
iaPNcqVXfFSNwjSRgLXjp+peaMch3xg6S1baNutlz4ceU57fJnYeLi4hHAwPDmpn
GBJ6Yre3jiT+URl9AuLOA31qzLPEDmAz2rXuSdvyg7uN6lq3RveLSXjuCTwZFXB6
iiI4V1g8dd3EkHqkq1qtCQEN3sHZRUQd5ACuAKOzA1rqSjJ+bczEtm4qNk+OoyFt
TNHiJd07NEvWGv/hlzr1VmnhIgSP1UXQdrHpn5zsdXGMCErHTQY8e6Mgq3EyXLPo
VGBizZwGL9BsJ11O6aZXNtUDgzErkW2brSStPALYsJUD7FnBYgKqkx9KouznLv+P
jf45GhKjgcTpbGWqo0ds6nhLrrvDDB328CE+9Bql18N+4yg5GAGoJGiwNCNxQusM
+HzAXfUNDWGZbhymXOko+e2bG/6APgAcBqnjQVTFVfHZoaQImbeTyVxxPgCGwAqK
lZLxu8vIGFgQTVSmTGMggg921x9iCWVxOgKxHO1t85PYVu8k5GJGx7E82kvfzoAI
3xuNnsU2W5EpLu91iCT2vVM+leJh+By45kcC3G2PYylJS62qAxQgVuzFwzD/mZ7k
WHHbWYN2xHPs5UEMgPOniWy6XWF0/HRG0EeYqNTiCtuP5rrbB7bfd3aXFZlONQsF
RSehD6GjCxG9Iye3ReHh2O/P+mGLojg/vLYcWio2hXvN6skVMy0LYLxKn9naybkx
7r7vCURg4q2EMo3JMKuKiMYVhuiaPFvIdcrDmYYTeEujeo+2+fLyYTJlOkkFedEP
nHjGT293CfLTi6V7EOwDICamP/bNBcUGc485IEF2ul0S5eKUWFZFhMIf4wv7FchS
ulYEGhxOpNGnV7kdJGYT65gVbLtOylsga2Xobr/Sl2t51NJuZx25q4jItJyO1KA2
2WYfT4b4IXigRdYW9JVDeNnoq2uyPhdTdWUx9pqzXJv0XrlXbs2XRTJz2j7yTpTN
hzq8nHDu8C/fONEQQeuRJ4Rr6hh9ZlwO9YuwLMSJ2VRP7V0scorQo3y32KaTOgUE
lu51DQl4e/gq7X0SPkVisSx87uzDjkl7iKDubSEQukjJiea6uoCaHeOXo4yVNQ4+
2xYAgmKfdS7ntl2L9XYIi9kB2877mXdjAMnI2OmJcst2XVqgW9v32pTYetOkAFz1
c17sNuGcBAz/O3VDnf9GEcp0MzhxJxri6Cm8ALBEL0isAPM83lWWa1zaPM2H0YkU
qehpYK9mE4LXK5sjiChlyZQQX/hRuvpN85B5oMxatnrTlCBAFIoL5ztXjRfJuFa3
3WqayfUffofkP1dhXXvv0PaH7CMYYjGyyY62YMu+ms8AuD3HJPiJJTlQO4BJQMbk
D/2qGHJhMU80NG+CQhQimEakLMjyCLu0i3MT6wHDDzf5LypvReUXCWmOXUf0FhaZ
gFWT7YQgt3QKU9Qv70aO/BtP4COaYb3CGsdXebCzlWcACfJUYRi6q9T8PP9s7vvz
R73fOLQc2toxRpcJMc4soL8nFLcQ6RcQQfHiSY+P3VqG7t8qgJzk3GO0lHNn+13p
MmuAXZm9VKCLy26CpBh/ubQE2gW4OdgWa//hqtlZ99hezmK6uY96DTJnqjYaHgRU
cHJ4W4IkSFoqUbY8HGad6WpUBosVUGA1wiHqIpDSrkOuY6SkItrnLjiH7bu7tl6i
ZHKpXJz6w1VphedkDh3Udfd7LGplAkoncNZL0/38vKkuacSxSsXz9dSJ5C1ghYsH
Nb4ECVgWN8LI2HhPBgidH/baTMLdmzgSD8EpPQcDC64Li6tAqstkDuTM5GRKoBqB
Vu663DoMX3lZ/I0+EUUcaAT+f7VjhCCIWxFapxmaN4IK2v8bPhsuvOgXZW9YA0+c
DtPXhhzqqSVsiQhLU8AZtqFjuzV4wvMz8skdJ4foa/w/3h5cJGdiEqZynxDpsKm4
DyI07B7RCWEkdgQH6051urq8C4v5rSHKxR9B5hslfgPHyeNVqSF2Cp59SvcxbkQd
3gqICGPN4CSo9bAvOpMrZc3FVIVW2EBqjWqGr9LD/hgw0VjLy2tYiTEi2fITAZdP
o2qJCENuqjYsNUl2mT4L5flAshrAak6OqdmOucAUlzYwgC6LRkOpp9N3XZrW4Iem
Gs8Hf31bcpgqZ+BEMWrB9xAGrrR8DcNDKKVPuw/0tF0+RC6dd8AiD88ZpTcXBW/l
ZUNoP19eiKh50NTiaiJ2iJ7+MJbWqJqRMNY02GU+hH48qMUU+obZgbhfjSeyXKmg
3LNT+uALGxuY87iBb+IrOdIk+hDgYrtQhVyq+pag3RtgwyyZ5e29jqyjzEhEwOEc
FVVYjVEXPwatloMRcfrKnuiofmcoHF0tbiXKwEjpjQbaKT6a3O+lXKjho3CG/oTp
dNbInOpN9bQAp2lNzCVLAq7WGFICuyujUe3RPj1Uh5Ht0gEYHGU0rWrdAnY+9M7c
jsgusRyXJoNsHtwYY5BZ5+JYJLKiAQw/IzE/nYFZs9Ts9msucQG1qCfwWQtFXbnV
K9BBB9kbnKv35V4+4c+zA74vmEQru4zBEX29uDfJbDOdpwWdkZVuR00kH8O6JWeT
JyswXoJaLP1wS79nb8LDPofpi0BDc265oBd4jsGT529VzY2/ZXNgF4WDtZfAuvzQ
DtCSK6KONehxUv3PtTuwZUTQWe5MIab2PLogLWlLBRiOTLfR4ilHz5qdzTzu5tHf
XU4h88xYwXARb2+58hw0cFRR8I/3JJZEHknN9ON1PO4C0O2BjEkzp2sBa2UBQyrX
pW9+QhaTywY3vylVyZVRskC+WsflC3gQXqrW301hzqUgeKQUMeqljSPqcxmTmY7L
p2h5RRdM2FWJU8+MOB2TfdMkFeudpkUC0/g4q9V++5C71BShOyKkE+nhjQRjTBQt
a5D9XPQQSof4Km54GG7onLkJ6FE3WLMWM/aq/PFZ7w7K0zz+kMYB6z2kzvYixkQp
4uGkQYl/PhQP8oLZD4RtIvGrWGUCGdCQl8J8zJECoL7v6te2qt64eBq6jmnaBRea
ogtSP/UPm25Q9nyVnylv+Kh7dAe0AtTj79SMMZsd/9/2SXw2cFboiMK96hqGMLdE
KxjJ/7tT6OHUNkwcjR6pfk7X4fZJvOwSMbWE+QARvSU8y47qcqLtbX5ocwEHU5OK
VQ3kjPDhSwuheImxAcBUABbSo7KR1JqL0CFeX2XAg1FxBioyB9v4mSGDbxRFZAav
tXeO2B/qeJha0eqBCcmPWBUxOSRjUIZjWs6sbw/KX8DsDXaIfDVLgw4b2qdW1FjH
mAl65sIRFaqADjleBYp0HgD8+neuoTasXjaWZuNL6GsQtRALGUpvJ4G7ezBEOCcm
HNI3YydVjsibkJmeWx4MSBFFb7Gj7hZLKsrQimFVPzZcRNM7a/KUh0avqFi4XRJ4
yoOoYZvpgbw2pPdmDWYXCOnFP7PQHUGZhSjqO5Vrj/kVnJbCC2gqzKA731bcH7It
J7lwktk9BbdD3KCGQbE92DUPckeh9C+egPca7Aigi4mKBzc3qiZVYtvXpiF8l6VR
K52fikoRA1MkgrhPKHfNQa8dCz8tE9el4wf7COfci8PPXjuaghVY+d0gyGrOM+UX
1EJZvs/F62az8wVffCNheg3Sgb+bMJnS7098VOkvsMxIcpLL+wYoEEgAwSwABqHM
CUmHKV1PEvvu6QSb0evQrpQqw4gjtaO8MX//vVgpB0tSxtkWEtXtLoOr2MqED+S4
JoYb0YIs3OTwwIa1TrFJSY6tAQLY6uaesQVKfjuO93IgH8eLj7vy/uJG+tsWiBsi
QT1jG6DRrxa8lRSXPpWT4XCV5BiGFy5C8FY7v3d9Ob3tlsBkG9Dg04vAQz16UYoI
gcgU1aYv2NoEFxHWF8iVDTSUJyeeIGZm7LD1PHLPpBNQZ1mlQIl++/SDmzTCpnVY
/U4dA0GHzymwKiBiE1rjhd0JHX1257X1ShEh1/nmMqLxkcuglipxmHpZ9zeuSiPU
+ZnP5TxKcTlfDqbo7jLj3ocK8eaO8cCZkkMdDfvFSqukCX7bJ/pyXCLKp1d39vRN
T5PCyuvcMtA1UMmBM5Gb3zD6hwDuTf9GVDWLqyM/YYyMidwXowUZDSdgfvIUVU8j
Hfo5Z/Bfu29W39WkmbBO+eC3XwrsICN8UN7KVCZT1n5pzY55tb4qhwcN+1Biwg0l
VacwP3IRns0xKBmZ6UdNYUrkx0KQ8jq2RiYoe7qdqaUaring0PjWC8aazDX4YUwN
zOc57yqaSm2fCPxHZQ2iGn2YcqZc70DxmbL3dyvsiUL2XdvF+PctgwZjUZDgShOq
33T1Y81EhtQmARYKr/+hYrZUJneYICWmL0OlSJCq6K5T+43DK2F1gKL/rCF55Dgr
/GWLLGcfAPVpTFDcmF2ctOdt1rheqhn1iVBKPi4gHViaBCcmwvdbaZOx9XS8drGm
5gFR1ytpi25l2LfMilTIYtYmAJLCwUPO6EqNCdWpqS30aThbS2es4i8QRJvOoK3P
CSeSNv446HXcZgwCVwsZ4HykUZL8PS1uubbepTfu97LOGxsPvdK7GSkuqzMuJMCs
Gsr2dfufa4FMHD42EcEmT2X/9Fp5vchAXB3hD+cs1cuZdJyGTWQQBdssxSkqGZgh
pH1aBHpi2qFE7VxVcVwHOAjds6xYl8LiNRa8QbFTc7BqdM7hBOaHF5Q7FGZx4d2m
laCIm6lpUzWtvw++u5+CScUrBZOVub01TzXrMUVgSE7g3wLD0jvDf9Hv/mm78dhd
TCfCwClXPa8DkDEJ2lYS6SQJX3MI4EYY/1MLD+ywvtD1BBoAzTHwLQDwSmqViD3h
1RroMvHcRiBK0FwkVOoRV08IqNp6ngRSgtAfF+SzLRauszofl6sR8n3Q8mWTJFJN
4E+UEYO+2SyyxTwSH02+7gTAYhUtNFHwp61yoHGpbztYJaja/bqZUQrYMd8uFPZf
9l0UnGw2xiDfN94Yt+HpHxayAzd4/NBgM+AQDDm+P4kE8dvGgIYKX/9gyD4aUlGg
vkyT/9X0zR8mRN3++THfRNGFhtxV4qEF1q18NeWQqE6C2tY8meW85Th3zHgzS7fx
dVDautWUiC8/0mjC3ssL8w0CetLPXwMXanakbDiNIcBc5PSO4dF3IhRdJPwEjyiF
+xYTDx3ul87onra79Fvd3Lg/y6SaVsUVqecJAqB8QJIHTommiPNDpOwJXm12GZjr
FXt2nDdlPaSNHRMYzyYGuuuCyiWi6b6e4wJtgwtz8xDSzlLqB5ZClxSrN9vgFpPb
BciPsdeqvXfBks1y2tXi99mDRR1pkR8voNHvFf3T5gn7tJHUzCLwkaErr2cVi02f
h2Cp4M10wYNaxYxFH1/CObQFlYIeVAgU2AjXRGJ/WjlKElkGt9cmHFFSqE4Cfd+S
RaVogrdwj7ycMto4V/JBk6Sguc6KNO+Oh2Wzh1Yxk66BEw25YKff6d7jR0gePZxQ
iRkpkana9KSx4cygSYdrtf5zodUAdem+dyx/4b7wDbQ=
`protect END_PROTECTED
