`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DWVq7nq9eXuh0b3Di1LOThM3iQHIC3mRr8efo7HtHhKJLs7zzqLBJH+vviHAC+FG
viGGATdCyXFjGuSLV5f9JBGr0hjBpa8mvZbgGXpLIsB8OFs/n7jMz7sOznvVO/z+
QGSMveBWbScR52tFPeonpi4LkAibUdyJ/zh8qWbnJdjc4NbKAcIDL5si7z4rZ5h+
IWiLkC/gI5M/PjqG7aC+mwoK0mHsKb6a6rSZjjFExGxhP5aYEp0qn72tWnAENmNc
wwLSDIaYD91Y/TkdO4YGayoXAVMVi2qpO+OGb4DVy79fLArSCeNt3Do+I4XBqGO2
8VSHdGmnFi0sVIxJVNjPHzr5H0m6OSQzf+usOSxYU++2t/ypSK5C7fiUl3pWoPGK
YqoGvDYDr+aBDtgGXAwiP/v8ut+nn+0FcGuUKjSqxxkKhr2BCAP9hK4CXSHAbhio
KHq5+xmwAKBVBKvhmy06zkmRUnHpJS90MSkOSE/Z7Q8KtVPVPulWQ4OUFKoNcZxI
VadyiNA96Xmo69f79X1lPJdB90u9FM5YgDYWuDhDKQijqpDXvRcOOP0naffF9uRn
3EGIx0xBwaWxe6EQiqyruYIjpDQWcyj5pZTvmxUa3DxDfjDYnmsmkIE///PQ5x4m
8FQkRktLMZmMk/DHiBz5Lm6lXDa76S0J5z6u3CHS+qUx9vK4NdNNkDSp+AZAe0VL
aYR5Mwyyl5e6+9X/nMgYNsSmcivv4oVj1zp4DB3hdSo+c2jXTkyhM1yOEl3ILzxc
LsbNI2UMulRvO+rY5hI/hpDig+PgXTiXmP4fODH/I+WTsWF3wjIGpE8scy1tWZ3y
pgRN/Y8Y+QIVdQnDUXON48Z+wBJF/cesMnxm3Fzx2kDMuWSsA2whIx4wjO5YcgOm
GRGPeE17B8Wd1n29ng9j2sayVSnJW7zcpJMNkFQmDQk19ps/FQlzT8XPoSERqgFa
rJySnrA5UYAA1mHamaXfH/6Get0J+15F9Sob/4ZdJSmx91jqf/7JQDVQKEsfsq2T
wTC4AIVpjE1tZZsK7QUXg9FJccg/IkxLhT5gH4ZKNl8dfOlDSf4RmSpgzX6BPto+
rzl+8sPpCsBeAJjVm5VamU0Pln03vlgOlj00myD3gH+eGwHlf+GAjWggxBJnecq6
whW0EnJqb6R93zsgLKq3++WkEX+1Ehvu4kbPzqj2CxRCnS03LR5i2cDXKlRQbDYx
id7BBjMqg8QRtyAPQApNObw8LwC8OkX9FcS2RCfwowShU6u1ZIncSMVSgXIWVWyk
B0YZzJeG34pQHlaTQi5rRDFLXUoLkWIKgbW8RkN/6wrNvbod1NWJGqrC7DuB0v8t
qPvz3dptmnsJO/YBA9M7rDEUoKZMJ0ZHDSTymF2xPihG5qS+BGJF3p1ExdB+dIYJ
VikFpJBfIMQG3Xr0m4xqe/lt80g4upHS8Dwiml6rqAt6O/AGyME7oLBNhWi+m5L0
4l9vevf+Hn+ZM4M19xPqhNVPPkGOBZeyD4KjqHcw6UoHIG8ruh5foZTdPq3XSm+R
TCuQkNfDLTr2BKpqgr3zjFfznGZfbi2E/Ve4wl+qt8Xls/VnRP2jP1XBS/SLEBzJ
5nR4s7GSfWeoRBiRLzLAJLLfccZwo07THEKOVmMv07wEckkiRtKzgc2H1K1fE4yY
XZcP36mIwOGswXkP+nX2RaylbnwxCQyBrGtdhcBbBpnPtNUYnJ/AN5n0PwJB2ayz
++JKRMdqwFKscK/J09mfIhchF5i/mBcqCA0xaPlcUiSYNhqqrBTIQvVVObTs3r46
V+8da313p1HDnfpN73sLhicW8vCMr3traZOEkivym39ooMPCn+2wKVSv1tIaXyZz
BLvko1Zs9wCPgEHHeF2HH3PBgz5DhjxcU7djLP8QWPDAKjw2Ne8inXTsvhiQCfkf
/UFtRHTk8hmhFWuXa1zdOD852AN8OVQ/+YgNOZpBDaN7dRY4jlrUqmtJoz3ZosJd
uEwL5lfcHXGsHkXdQUMk5Kq3NbTcExJE7NdDGG2/tUpbBULhsRBdqPcvh49nBAk2
qDNaqI1DW5y6mVqTkUgOi2uSpMKfkJsyqjUveht7uwxBHyAhrdeGOgjxDPca9x0n
tAj/ug+WcvuuUoxktXlgzOl3t9rE9r0xxzSfI2jM3evBdjFm6RnKy1MDCTvjlw7u
DyjR4NQsTTshZJgFpjYycSSrvwNSiQNosaFz8TpLpbWqr/lS/PhrpOcW8Uw7QU9r
sWoQGxg5qPGQ14dnh4lHJTjm/X0p1H0JBqI67lpAT8zPZHSWo1/GYDFtfPGjXDCp
1uouwn+VkhbShnj8LKey8J/Pjos9z9DlvqWk26ygqsIDLzKw/vNvhXJYDgKAvKBc
iZQnNC8kcdPVGpgWsW4g6ZLdukw6eKmDQSeNaZb0Dn8MYrhbrXHCrx8hvgl1u6Lw
k/sYSRyEIuTbfgd4oXbsNUJqfh7pK53x1Bl9D3kVW44eCR8Vlmi/1YcJapF8BLZ5
ETLZ67VakrepnqsF616quaDBfabLy+yBGoU3l93Sx57N66oWK86i+GckTLINFvbG
3ImucYAj6O3/rAavAWxwWleRyQFhWgTNNNNz/BJEj3P6NEAR3ZFRa4wGZrrsgEMj
A+/ZFX7/8+dvOLALWCDM2Ztq+uIzy3xIuMY9XnpCGQuUcUBMdyMxFhyl5MXVWRZo
bU5QvcL2lEeMf4kV3+aeooZjuLo5kOtpPza0hedtTvM+MV1Rm/6y2PsiT37+IjkR
B+vmIESwRk+IK9h17L3OgjPgSqOHJde3YkfEANaZ4XyQH1bCQJGs0RWdIaZlRMHn
yWzHvstnyXhN5Diup8otBpje6fJvCcvU/Cz3MvMCZjAMp70AWIuPn4vFA+ggeuh8
rbzb7ptgsnTRLw2B1YgoZ6a4zOMDcea4NtbJc1sp5ce+hDqyGp0EfxZdjOlK1Qbq
B7mkhbQn1hagl4e4/CFDIHHkAktaZCF5KGhXraeym/0YVyiWbkb5C1fmBboAw965
ReigYPN4a+nZVpY5n1eoraVMoK4Pz3OLjVpZ3LC3GMo4xbtQZOJB/S/isR1DAHlL
hlYZwSbXlLOGdTliiF3U2HLUVuj3AVulH7+ijYHTyjj3+YOJ8yfB3RhmqrgDCGW0
o19bMo8Dv48q1enHe06GYLO1PcYuaW8CiTRQFoLdRFNl58xRBeJqKbxzZVzvKtYJ
H+bCwRb4xJ7ut97regp6vDt58QkhvL/NT0m/Ce3oYUkWnFD9P2RBpVoEizZkdODy
8wP0vjezusweDYTjwRPGUfyCzmFfwQqT+tirsjJJljJOCGA0REbRmvX3WRkpwEHW
Gkzx09Hj4O6bLA3kGwIBlJMWbWMqud7mTlF+ig4ATH8ivTtgAO2RSZ1uz57iUchu
uvaBGv71UHH3nFrp+CDtXe6PbFeFgonAVJ5yQlDCP9n37bR45IyF35LU7Jume15Z
kMvyO5ykbHDJtgezJImxRkSIM9/iiXaIRGhtnUvGLJc0oVePWGVUn8Oxd0hlGue6
cxj6QyooT8PSBDZS5kN6m3LP12w1GBuO12a+Sbv9mvWsE9gUV+9MWyElrRLz8AWx
2aLmAn8jhjRzLse6quHlChvAonKg27/LWduGkRLB6z0tCrS9UqGI4RyeqcY5IMSI
ZT07Q9/CiRenmHlM8199MSgezG+usd3Zw6ZXo2j5oyHXIo214TJ1oH3neFSSd7We
OVL29UL9/pFqTQmsGREoV0ykkizX7G1nkHGqKdZr2VGk9lm+TaXGHmXUPNmzp/AK
Z9cvvqAKevXPgH+gyqk3YzrorbhAIkYaLRNHT800rlfi3h8xDneeymTlwcPO7OeQ
DHbEvVDkmH8lWNOosrzXo7sHOBEwNsKzk9MzUS3ZNc7O5FUqcI61DaiZgQUWUYEg
KBmdNDjbg+n/82vE5kxvXbrsxBrKSyHDY2bMo/gxZNzoArqO+IE8In2gnbZ7A89H
lZFofq2uDVd3Sn9jhn/h3hcI8EAVmjp3zakoMUNZGAf9B3c3zUOmDH4Tzjx2+oZe
s8dt4gno+lBKuU9E18ZJhkErPLZzLgtERNrlFiuwl7zS0Piy/NL/w68Hls3Y3Ukx
QaYrBI1wX0MUNmgbGzB2gfHecOMEJP0WQht1MbPkbeeoCdawvHXWsjCUbkrqIf0c
KmWKrxfpsqulPisLj4L1JgsQZfPBYYBpAJp30Cqn+uSGrL84/+muiXaVH+bvkUPk
s9oip/tZ8WfGIAEKd0WK1aV2k9oNhkREzqn7lsn/kGnoq1RgI0Ebp+NHu5KgxPsm
FblzXfcGEvJHLxUt8IfFBhE033NhwD0SEx9keyTGjIClMDw1uLTYeKZEwWXT9PyU
1EO9Mkv6bsKV+fItf1M0KoLfhhTmTIf2ALip4KO+SM94/T86lqmSygzgEBOAgDa9
9ADKTkFxCoxWS1m569OCPEEQQUv67krojjYI/Ma99CI/bsvaNy8iUjYjhHWESE4J
NXSrazhs8jvpMge7I51R4TdhD9Nd7hP384NIc0K+Vctio40mo0OIR2sXqVWMQxF7
bWnI2vZoznIq1yhP8E9fxlwct83bUPTWsMrG2paG79CyQ/N2G/hMDA3qhW3j3n4j
/gs3lz3chRo349y8575OuZ2mEu9HMTvGQ0vOO7Yn+I/9xRWT8g71OVcyjLR1HCLo
4EQzAajhFUrmvHifIyPE0RVvzeBZXdivf0CKy8M3t/ZrhiGBKef3xgODV2DhpOgx
PJsdJ41ezJoyr29t9DJTtBx6ZwzrII/nTmrKkg04sfEGf20Z/4phYZ0/lULTAcbE
KlQNNJZB9atRKCCvqrweXfbH7soKUKshFiqdZxCSu39bXHT2OSLPDVNbGLjX9PQx
F1wOYhs6K9KlrDX4WYwPnpEWczDkJdlJpa8frizaGRKoyuf9rQi29vHK4KmNO75Z
HUfAikH44M3gOf6kcxT0/wxfhvC3aLiQqUs4BJGDPX7syq0gbSSqUwKNrf9WvArV
EGLmcor6fSN7Gjg9RLKyHiGNbuhlGRnMQQcBdcfMfX0FkGpS9mLaYcnoR8C8DJOg
rAWBOQQVUe5nUHJH/JWRVw==
`protect END_PROTECTED
