`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wRRTzHP95V0Qd9L49qoB+3nZFRXDTMpWJSw56HQv+zOq3Pr8EhNU1o5qYCA5ynmu
qEPSDhpeC5t+i2mNikRbHxi11uz3UqXYaH3yVPhLP9s410dqc54G1w1AyLMu3ewI
id3Xn0nqaxohASm664382WT6WOeGZgsQ32mwsWXka0ZK5Jwcxc/pmjmAWHtxh6sz
DE4aInQoEvnw++L5EjZ/skQ6yKTe2wVaLLkA6izdThJ86zipauwMGdA7K8jLPHoy
gnonH3GXhzKuzxnhGOZinYiiR/UrE6HFsxkUqLEJq5ezB+vANj1RoE5/Fih8gQcR
JHleEDkmIp7tb8svt1cPdIMYJogrRpIMpezDFqDT51TiwcGCzYDdxq/SY5iCKsiW
ldvIH00NGFRiMaaEUzjIVtkXmq7PivmFfe1u07GZGSysNPov6t7mMBh6mOj63xiE
O/wJlRje5ppb7FEzYBeqQ+Z0OMFHevU6fnrwjpKW64/aZZR3e2T5GQX7BdiStDAM
rO2mSZE1K4y8EH/QsWGyq14Edvv9CTtM7C9IJaECmERGlXIFr9yWxYcsk0YNhlIb
KrNEjO/Spc9EGLTAHuXI/pTDn5dMvQGKtx49FlgTA2kcny1EXqS6Whq9lg/Cg3Mx
M6VorNtcRQ2+VmJAMmscaELm1jyUdS3EAuBPif9cUa45vLWJRhZOVZlW4ViS4pej
JVcnZr246I5eazuvsHGte9s+60mYo8tMM6WrSiRnJZCDqQlfgtStjxeSjOSBN5KV
CqswkRdS9kb9Bdyaf2f8/dPwNXCk/SPuxWoWi/lLdQUDugd9KisWzHAv7rC64FRj
75ZsloMVopdhLYIornA96DpO5OHWnrwCXvm8ea4tr63SNSG5YfB+jHRFUvxxgmot
KocTdzF2cWit4Qoccnqe+TolLFIZOMGH7Z3S60coZ+XvKwycHce7i7r1zLEmvEoM
lJ6bovSSGFqNz2ufxVaRRzN2nZzGR3x3B+BnR4f7pzspWQSRXWOoo1tgl+gJ4j0g
skUldgpZnJusdfq/J9TrkYMd0fFdixg1xfZnTuje+Awk2ZLh99rkIxVBkrbJPKJN
BkkOrXSVS/4i14f4fF+ia1qXrakwDWqh3H5JmzwXXqOneoBJhl8F3pNF5vTihe13
ScLLMA0mjdx2r/VHw+EUtje4Z3Z5rLp4UO+s+yB9IC8k8j+IrzCnkYjYteECKflY
YN4+OdudMyoUJ3X7jujt6SIHJLWutSU4q14OXi7QwvbgBanCOxy4xl/ed5IvaVqf
Tkz9hMdfqGqtNfve4iaqt52n/em/6mCSbtJw6zBeV9i9sqi9UCynbWEObCWdNc34
/WReyLnXnbrdu6thmbIYmhPuF/TztPd9pNMd0gDK6NLGrut5TBYfoYHiVoYvN4IK
Yr0Ffi5s8YJbN5C7W8P9HapbrGjJA4iWe3jvjM8YbflE4bNdpK7kXOXul7aCtzRb
qAhyVlBAYM3T+bX6WP+kWhY7LzAPoHb95EnmeMkrvRvaAKwhgScDM+bK1blwtyau
ifZjz8ivuQzg6fxDQCZeb6WKFVlzD0jbiC9bZdjDGSGsYYkJVXq45bPhpAbOxRpj
D6pT7hvgG6pN4fgRKZ5oEZZEHZivoqfMbCJn3qalMSYjaY50vy7etEwC5n94WypP
roYglLLsNf5Fj/1L+jfHMO5NQIb0UOn8fhfmh6Z/dYKleBRWFaGrIGCUzd2w/lRR
y+26NyfDO/CbQ0F+2QIZqTw4vnU9+zKzxwL+h42T31Id3IsNQEZI684OzgnS/GWn
sUfL3i3AHdF7StQhq0HeX/qnXIX1ugeqmujQzYyXznUEAFYMl9fQlGtbMdUmqvc6
yBQjUs4D95H+GLZ6auUkGIn9yRVTnN20hVd7phM6Lkfg53FdFPE0ZiclkkZxBWPC
IZfZh7R7sRsJ1FJswLCONzf9i6jAFBBgXXC0vqtSEVpm5/TpLl+otXdnkGBvKnG2
YwodgQCopk1Wi3D+/kdbidDnyhl/82+VebTj1fK7FrwfVIDDNtUJhIt9iIHL+fkM
4CuHSXEl32+tcZGA8+KdSN2uDI2DIeRwE2D65P9ODmtfdJFXg5M6ijtjzFLZVWtY
4BJ7Mm0WBFRJ4LfG4lAbTQZG9eX3gEp+qM+B79KtDDADUwTBip9UpWG17ia+PIcV
VUh4KlNKfzjhiT/B5G5GjbGgNjTAkz6HE2uIdKBKxLTwLvv3xtwATgFaAosyc0cK
bjYJq+AUKeXqrx5nm2d79Ll8BjatPv9HjSIMrrUGfHV2xK3F+I4Hyen1dBJdRyNu
vgqKkmfzZI9+tpay8L0RU4v2hWI42aunPpdvkSFgVRONXhmLjRY2I41MaPH8B1+5
RFo2CXaIeQpCJ/f+mkHK9y2XsrY3xOOOPbGvjN/kSPq/YfS5fHs0WcFzjsr0CReL
51tBnzAX0jFH5jEtzKm70jwOXcxeMKrB6wpp5nU0VtXIL8c/ykH8AhmXpDC0F8Nl
Vj6a/kqd3Loo3QdkDbWx6zoxaEHcW5/8kJqBR/xjSXy1g7erBr+9MJqUVYBmgq1d
wFfDt9iRJMIzJnZMPSgkNMcw8N96OTS0lBkiw4ciaoeBYmtHTarAHKjIpF0Vgd6y
cRbJf0rcr6N7gZE5Ui0y2LXK9d2RRPmdnir6G893G1Hw6lp6QTzOVZNOIpiPnIAr
3BN4Fv3u1W7l6J7SfHMmgiEkoS3ACpq32yHeXLwu1d2rtqLiOx/W19c4FUY6ryKr
lgAVX0SQTUDBpbeW1Ig5yg==
`protect END_PROTECTED
