`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1ef4OetUUiHgrpocMdfEGWgZlgEJ20vgZpiJi1fe9yjWby7DO/jOXC5vOQbTGhr
W9kUWt2p7ZPQEANK5NZgw3zFGx2X+I3ST9KpJrGkzPpDvmWOXpe8OCy9/R+iX4u0
kTp8QOdqpFTAedkftXkK+gE2ZLwU5k/RNWbXkO7Dn4BsKiSrDMAP050xBn5nbmby
eAKt5mc3iTB9Q5Z9w/3dB/INp5l5CCoqKcAZE/CmQ1PWjp5y5sRcYuAztx/4tRhy
WKHmNKLQ/Ryj6f0LdgReGe5N/5WSh98gBAh9l9fxxXTlbgLAA8BJRYvlJDEw2oHk
3asxCfwWub50LtHsnyM15Xhc3mJVjT2TrJvsF5H4D9kCf2eNpxPuGNvcKpIOrdTK
i60NKUCq4ii1WoQKAa2Oak3428UDOuqSogmJwWBsPnHKKgxeueBUxJ05AYxzZ7xy
Oyo+lHs/e3wh/PdKcgyApTg6aJAY7/P/HeEGUr1FvtNLeHSZBp/uAktV6Wc8yaCL
hN8Kq3HLEQL43suKb9/hsuQfrN5NG1fKw3sfSVFz5WPUlfd+eoha3OYfqfMdr/3v
ftdCzPkNSryqAq4I9h+vT3LORy1td2OvDyOeW0St+drlrl+jcc4e2/QYqb0icZxZ
iZ0LNebXNJyCkZPaFdA41otuRNXJoTSn/0hIO9g/nJ2YVQVl+H4JidCzzpuZkanM
PjFIVaMQKu2Hb8xDmYhGnr1RSdMOM5E8ywvkbSy6nP7wHOm38ni1VgQ35nhIjxOZ
9zzawTtsPQGJ/VUbhLIO2Mul7L+iM2MHlRVZ+BukGjjfleqAnVlSlJ2rs18Hx2uG
5yOtFBvXjnoHf5Pul9EhEIc1LKQ1HIAECQapp8EOUKO6yP5OnvCpj8bMp1pojTOy
4rD1P4tnCf32Jdq4pjMhevgCR4wlG4fQluW2yNnU5hVk57HplNMeDxd9pZ9Z/myJ
7ny7UURb5FvrJNtKe92X766c9j2yhbwpd6m289+ha+q4ZGapnZF56FgO1beZ4NWA
WXfVUOYvqvZKs1GnZPxJOxAqj81AiwGlSqQutbex3JtPntvaWyuI+J4K4VOw6s6S
ofD7mvju1NP3zVkfS0GZl0jdS388AVJMQnEYB1su9oaVxEw7vpEqLYGy/hETIhBz
SEZeuWKsIzXpojWAqLLACN3mJ+EoEcgekmGLVMW195/zP3EsgVUVS3KUXonpBRQY
+sUdzfosvaZlNhAkAqLVulAmq5ZiyfTfacgu4siqzDtWf1+EgJnywxc+e16a7EJs
WKysRxI1V0afdjR1venvUXroS+4yuqezYZdd6mXJ2gTz+9kStsc+YifYLBfZDEqf
pVtjhviKD77QBwGwwSigWr026CV00tSeyNCk/Muli6hWZoIOa8XT5z3J/oGNsNBG
2w1t4zpgTRw6UDNvcSjTj9/pDrqh9P73vPwN3WV4ZmDdyfY9vouk6BnhKHNXuX9t
wqFY1rtdAuFBUyPx8pJR1/QWKihlp/pU75xdjkpWmlahsieyC369KUnH2DzzOQqT
IrHBhXO3SB4aeexK+xpxyg==
`protect END_PROTECTED
