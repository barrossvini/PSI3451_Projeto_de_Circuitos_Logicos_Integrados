`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8dlvS0VcoE75ci92EOYBOmS/4Vi+v56v87vT0J0j+uXmWuUwixZjvLcGASboXkg
HWNvgjEqB7dRjJ6c462CtvwommYK/Rs0DxBdOLLT1vMIiC5KoG/a7gNr9c2CLDDO
h75ArcOtNUzPqOcfTX35nsWzJykUvslQYZxZnKrchWm8nNKjwkO30EyXsSNzalR4
m3otttZx9m0kKrmkYItgmQmuIk8xzmPV/ZWXKSZLZnLjRWmuAFE3u8f+2qrcQFXZ
7bhNEKnjFqB9EHXOvtHXzWXtuv6KFOIL5rHJk32cT7sS+lZDYvRKIjkYKm8j3PdL
fvMMbqj/G0E71EhqIhsDkZud2ekTZ9TCQ2/jXtjTqZ244p9cMhUITpHQ4dCYRtpH
Kd8sk9VC6PawJmo3IJfFzqd5B5qzNspyEavt9Z2cEdTKOL0ygwWxDaYrpVXu9ZK3
9P3ucp8veQ2mgzKg9+nRIA8U6KOm3X1J1GBuGX5Py02pLdeyao7v5vgzaeGym2nf
j8WiILvjIOLgjlbH4Cz0Qexs+Klpe/cAnwfwAOTipWKVbrKdylI79zfiewWw5xMM
ZDZt8X0U+7d6g/iyXEqSgId7EEXE9Xax+yFh9BPa9m+MfcayvB9Vg7VTTGzd9pKa
wnyCez2+EmAijo1v3rsqfYDshX6CRkSdsGiS9bczz+Uesc94pV1IIohychJE5cRm
ClXQ99Xy7tPRK/L8sDG+CaS8RnvROZozDXH2W+7Iq3X2d0tmOqfkVSq1Ytt2F1+e
3SRMwxCCiEVlErNzDsyr0VXRp+zWbH90H8dS86B1Tis1xrt+HUIFFrUcFOIsCNnZ
JqVVxSXvYciLI2yZ7MP5JZfi3RepFSzdr8Kf89YBu6bU9Z5BEZQbVfg+oPiq6URr
0GodR2bCKasNeayU0F2747E8px4xPO0uohOrS/9M7ARCqwYyqmNUx+2na/uEKctq
f8roiCwIC9uLD6CAyUcdGxdQLampP/9cCZYtSQPU18BRrisXNnXw9S6jy7207GqT
eHa2+PZPUNQsRsstI5uZSBpszaHoWAVdRxie4gyCmD5ru2Rnc8tlAHKR6n5kiDW5
xjAYKwcOamMk5g8cQW3d7x3znbuEoMyaQEpr+PmJOYt5A1WGxkuiSLFyic53ajQX
6q1O88b/t7Aj6FM8cA3ptKNHT4CCWlYfMM1QbZRYQ1hL1qBa2/DDPLX0ibNykcFq
pjc3VZxnylZ6aSqQv/iXMb2q5A0kiDvoJ/joL5fO+PfMUAXcTsZuD6T4bimYcs0S
MSWpWy+DFf/3bpxBU7VTaDPsI3DXPDxxHnRe/dlDvT+miJmvdEbcua9dQRUg8XrZ
1Vct/zoXvoAlc1bZCX7XMX0waA3nvnPRUqt9BmT7LMVZ23D5upMibKlZpHfRAe/I
c8U2m6affed0C1Iw3Z3b9x7UJfY/bBAcDRrwTmTeFarjWEJL9NuJVpiBKvqgMNjg
JSVcP7/hjhq71w3DTEjzJIBs0ixNygE3iAxxvrBIjt9Hqs77jKOE4UxmH6IcA30i
SOuKzw+ZGHDc5ARb7wbFNJnf1yf2jDbs5UJjNTau2MyP3DO76M5LlBNEqJQXalnh
VcCBlOqwtG6BhAOx+YREixme6g2Wwu/NUZIoVNF+Y7bdu+1/t0SubrENe6jTkVTO
Z0+6doGtFU4+lkolyUZfkuFsNWWNMP4DQvNgkck3Dd1eJUfBopI6vXb0kXKTA8CP
mEBsIrCuzG4QxMRmUOW80mjBFqhhmZdtvYHrgyjGDzMARAxXOnlammoShynVoHbY
RhHzrUrmzjZBRsadq9+N6rjhzj4SnNDLJHl8A07kYQkmZSmrhcnWzxF9yFVyqLVF
NMKOe5dN5D8px92CS6IaP16G/JnLxKzDLAZnBmdyiNPdrdmnW0ZFV5zYPE9AMqKw
fUpgblKmE1N9zA6TsAB/B4Blkg9y8t6J8lzxALmZKZ/kqhgWn/DQ8nvF6U64xMqw
dNI9IF88mFLN18Rm78DxBkcgz+NVynuKshd2a8N0beNBYMl/1DKJAcftCuCwyaBC
PrrOXvHFyccaopNyqbPKm/xDoWHDV7hpZGd/vsnkoLZ+tkTUcMNSVHSjMrWx8PdZ
/7CIF29vtRiS880vYPlbPHpfG4q3X8RFfFWy0XoQY2qq6BKgDzdRPGYGJmgAxM9x
ooF0dmIPYZ0ErDl5pap/K69C1xl3s1KDlsyqAdno/b+7nmp5zK/qDPmpgiTvNelE
t84WfVf3M6MmdPTIxeGsiu0Yv/VobjqBUjEGVtSGHkYEEQrf9OMIWgaKk+TlJWO3
i8RQEVbZ4K8/gzkYgqLda9CDE+/j3jBYSgfgKUTSYa20HmATwLjG/9w293W1eenG
nPNjBdlIF81wgWmAxjiyORLSKx3IwIPI2phQGsp14GdWN6kBx+0qT6kN93c6Ynqx
6GfCwldgtLa8hIRPEPd7cEf64dSNSjgT0Ekm9/Lg1gIVS/opkDSvstZcJgxohNwQ
dhU7IIuEr1qDzL9bTh6a7x5Gge9FX7vaxkkEEKZwxwZkjKG9XJj/wFyqJv4k8kYN
GyI483h5Bz89ZYsaXS8GNjwDgPejTy/17kmYxVCoF7RdUBC0zu07C5VpRl+Vn1OK
z34imjr1DT9aIPaAsc7mIIP/Opu8BkjSdBzj5pPKrCn5wtHV0qKv9rvTj7QGnlPk
LnvupDtPqrYxkHkc3LxM1QJjpxlu6Xx9miBKSxOpo5mF5X2wIj6j2YOZkOhKtgk2
YmFtqwfvk6RK8ZNrgEsPhQx3mIxacgB7Sm1NjlMgIl2haxd2eASG2C0+QFTwjs4P
C6zEWW9azyyBYcCePJWN84ioUr0vxaWXT3gUV0Ao2Z6WLfc2m5M6zKq/tEsMb6aS
ruXNua5Jv6NO8Uycse7eyo1LZI9sWlBm59xGMpmOWUdHrgFCTu805jo91Lc8UJgz
vF+bWk18UGTLMdTIEmbeV4i18gn4A0PE5o+QbZvVNtLD4X84KPlHIaoToVROQrxM
a9QlKXoabcU2UAoJFIYudUZbdv83PFPhe+Wqe6ab3RG2yzt1dFyOxprdrOVzuue+
OsVE65G1qy1aNPlsBoy9Ha03O9g4KHtKJTy+aj8MUSIMtfQNjnvMHWqPwcJrgoGW
hE8dPxq0iHaz6yuSasIxAh2/0scb7L7BB+3nm5djppdxdDJ0UO9OE6BzTBogRQ4R
78+N1eSkORMV3zD3xNy0PIrXQ/M6bPf+1PNWcfRf0DYNq1gfGhAD+ADtt3vdAYvu
j/+DxhHIP0Wms2v1+jA790TdnIcYytgGBtI3AUiOQBT8IgaEiGDR9iS23vHlZwbF
7jOPr1sqlLsZIb9YedEEHAHkaDTtLChME8wPOg24pyFgTTP/PsxGJIZ7E0k0TOtU
e5+LF/oDCBZP4bEyilku6lWUHgVH5fcIHr7Xf19PpSPd4UJ88bj+uCvQ1bvJuQqv
oeKOo7ven+x1u/0Tc8i5AeXVQGvvylZ15UFOC32ijjLVlcSOk2POqv6flF4Ri8kq
LFwFkv9C7EGZcW5XWG7tdP3zatAdXGva1y1t1jUO8d4o1eeDzzGMVwqKkWNaSzVf
O7+muF9YLDM3Gy7waIUIFErQkR3iPtuzoTOD000SJr5nrjiYyNdS9NMMlrlRqdSI
SB7C1wg6TBPwVpYEbQ07uTweZTgoDhhm/oqrdlNAshVBJJvXQtITJUQ3kkjRmV+O
iLVhpKaA4pA0gKCxLDdHmXVGZ/xfPJWejTDUblofuop0s265NhAG+KOX9gqVejMl
zJ8rcmTjKjucf6oie82PKngHIv8iHX7O7YNUXSb7ZxRkY2NWrzQ/5wYPQvgg6Z6d
xdiiFy+JYtO3ZStwFlH5ZwyySOpKg+XRwVP3fBT/EbdU1K7lDDK6LLgCGY/4qXJh
iKy1zmljrcEXNX8gj1oiz/vQqhdxngg8jN2vL2zimc2GALKCxiDKW+SqqzgOyIKr
/I10TCYarEpHE3Si47DBxq36pbA54stdV0tavtRRJeZ8ioXEa3mIJFZx9dMyz5FZ
i48QI1mkgG99qjXwNjVMjmXtET8FE/wgo01k97XgoV4Mr5utJANLqKM/LLWadxdZ
P2h2kaHN7mB08R3Z8qUwgxZ4ZHd0s+ZQI24fQ9vU85RznM9r3ipVWVZxBpkE8O0r
5e5lFQjz19ZTrAqQya8L+ZR+jQZPtrhJzRQpkemPmiAKLR6KPAfpel6euFQUx+1m
In0XnQuzBs040Ter177fmI1yCIZhwKV3TsiBvnlSpLR+HGxidTjCluwLVdzIWl7L
/McNSOMzVkAa+nv/fRKXBMbB5+zOrZcHwBXkkc4hMy/WsWO+z66a4vcqj1Jb+1ys
JnRhcsVHND7XuhkhX2RMjou7I33zEq4dXhna6Lff1zefNaEt/yRNRfq0mS3GNTc6
j9k1I8oggvqb9hQlZNsOr4ZCou8xGxPhwMdNkBOWXZaF7ELzDKZxfNMq6GVUkxBO
o2Gwegpv0otf6iPAMZbN0iR5uZ26lsauYpe5otWs3fldR2xSU0VepvdjFlpchmb9
rliH1Y10AURn3GgJNsHs8nzievQBu+n6De1085IOolSalJHTelxaBUd2ewFmH2et
4oU5dScFTGGqE0MELFdkUzGYAHVZY3dpFN0F4UzsyCF7cXS8brJCyM5XGhsWa56T
U/CO8G8nVgFx3mZGvRNxyrbQuXoJgB/QLIHc6vrTJcudYnqcsNKV8jMhOKATrXHB
oJv2qesFfo0ekzvld3IEqbJ69ijPCJwcQoRebRrHTG0RFpPPB8LUR/fLRwpFCWAo
2fgE943e2+28qJlzpdmfN796lp46FJ6yVQvb6fVE60dYC5ZPazqMAcMMAHUw1VaS
mOBg9zHcKL6e4fcdFLbqdAiGtl8A7OMlsQnbOt2NhDOQv39ZhN1vZbpTJpqpbqY9
vlga20E/9AOE/tXitEtiETbLgY/mJt1CSzk2AUpHe1qO4z47y/9QBQVIJNlemKWm
sboSZb6z0yU5Cxc9H2PQtn/qPAZQL+TW43to1p+mTkAXmSQP+wWeJEJIM62tWTfM
VAb3lcVpf8coky1DPVOR+cibsN1F4CMVmrgwQYOnUp116MQNrrlH/LrxZiw8PyK3
pNUooucSOJ2sryzDp0podXaY169wKfuMj5bh5S+SxXgMXSjmTv7xqKEXE/UFapAC
tDPs9aAOLzz+SCC3TUdVSG1Z1BEQFeWVSFige9eoXsuYIN12KBud/hZ2VpXxdOYk
sC9vU2ZSVjVoEgGuMZej9yjbWFVVeEuY0kL4IIHKuXoeW89rRZP/wZbbz+xshWrH
0+XjpFmp1KvHqjeug3f54io+xYG7Gq9GVwzX0rReU+Fw6WoyU4okps9Pap3R9544
Qk/17YruMW6UolLboS8EX74TDs97WJ5M8KSzSF6Nc78IN7IV0nODPe+Cocq90Gj4
O6aGBAKtvku0Lybeh9G3L8OtQCtbWE4RpwcaYtEuJ0KKm0awaR009kWoZG5g01Mf
dDLvxkDD16YlEmgksNGSy/Mzw+He4dI0EE9JvAtFOeJfyZwBKtT8dTVqYnvnsZm5
fY0a/lC/1b3OeHYwseXZlGbh+rMOlmsgyDKILwUu+qqSlp3b95Sur9T+P1/TIvBm
L40l0UK8jo5fqTyt5wrcrpWSZhLBnn0UjN6Vz2/vHjOqyJoDcWJCOidpAIFBEpTe
zqAmWSbJnDV5VW9JzQqVqrPkg9RLaiMmAul04GLDvpjGmiliv68JTF9bHjIS0KDk
IYc2iQtXZpF77L1aBLJZGcrRDtfzFRt/FBQkyefYzXSpKRolMlGAbMWnRXqD9JGf
OyiYCwTOOPLDkar7NIKGmXNkJ9X43oB/qVPxOtxPUMfkr/06NVZNEj+D4bEKMKSs
O94yXEXrk3P6VBYRdoJNkT5t5mqtoBIUyUk3PVAFRn7MujOBRFIhuNhtjb1lkKXk
sft4YyJlglgdgsmNGkyy31aFhQzGP2LDFtBqv9toC6V7xtjv23aPDDMux8HLNjLz
szqsoMk1mLQ8v8LAwxq7+ZMbeZRcwkGroeMc0AHGGMYVWHmgP0nhoQArPqXGiPCr
Tmld50t6UXGnyK+mXehK5ld+vUWGdgi7EJccKC/p4vRDn+owL1pP7RGFWWot42Um
/F3B+eRgAzUfyQi/kYtszLWNXMcjVfto3m7AXRQffQoPt8fPaPMBNtWoVA+j6Oxk
RyT5uH7t4WL2r7gv0+9bcQcvBmM/SJ1kftXjXw3FZt8cPO8TO7PBDen3XAS5z0UL
vHVns7O5oA9gsIhMJVy4h3bMc7lobFoIOkimtGiZFPoFjEz0fIaTg0aXJMIjW16E
hfEvbZ5gSYjjgKpvZHj8Kbk9xxMakJAtN7wQh520LTuzKq9nokDMhksgyyIUa/xG
rWWjTDcGSOfIugODLQFd7ARe4xipCkSoT9pBnk9vi2TuRH2oBzHEnRNkpwb2+ddB
XeVFan0Qnp0iaMjuY7W55+nq9TbmW61a73cWXoyRpOHzpMuXvgXn2qP96a86A25c
de+xMZdMcSRXMd3gidP/3h+aHcRTqZeaUev2XAt0D8gwPAkr2uOBEIntaZsVr8Bl
oc9wVxM0Ai2rGNcCornQDbcC7Cj9tzQ3jGe1e1JM3qrLs75MpBzO0vQf+a0caJtZ
96rqNZJCFoMpWucxDfHeqAcK+JJZoMQsMFdWVkJdDN7tGQAJsaIdup8AJCLNoCab
KPCNzUCibw4lDcshwX7Lmd8W1qCUacTVQUQyt9LE9g1FrUvIE1vnugPyWpptP3Kw
awB9WWhQJSDdO5JOr8iDPwfYtk9iKXAy5/qKkYKDNV8skO9GhrwWMJkr/17lIocR
8cGm5mRzOb2XHPPah9i7ENcyZRQh5DbahoRdzHblHGZIUQ+byKxyAkXSaSsIzFS2
lQuC+sMs7wZ1nkRCM8n3RRuV8zVOeTJZ2Y7lpATcpoxcrlpo9XxfFJM3H4roZ33P
GE43ZCMWaN/F4yIrsmdws5f/4araN58nmqtk5nKIwR0rqo+DjgEIu2WcRyD7zASa
2lUnuiJfG1jBGQzuTuWRw5Wn8g63ebu2pGy0inWWji2SyV28eK7fFOFM5A52JZ6C
y2o5V+Ak2E5jB1+y9L+7ftPD/kteKJ0daslR7qLJ0F/ytcDXDVpQ8UzLAi15VACD
wHtPbq8hc4DhXA0IjCMNJn3323QU0RQW3JQ56XZyN3vRkuBiVnajnLpc7UE4lhav
hMZB4yoEHUaZ4GMA4voGAXTq4cjqZQ06qTJE5S8O4qW2iiYXR598SE4liQN5DRaI
XkFqj2eTfcZIgNXKU1ks7e4GY/POv81lQUckaGEkH/q4WUg2C7x94ki74m3SWcQO
6nHlVPp9SjPKr9QI2qrj3cfVDtIBDuRH5P6c7ku+ScZVw9XfAqbQEzbQb4LfexTE
VgR63a6YRh25RWQte39fPtW1ftA4yZNW+nQIwNyM3INL5WqQYq0wKDcXTFYUdzVx
bdraAuBPHSq/0ICyDeXc1/o+y25EzM2dPbp7BHpRlIFsmOkQ+OhCv/6vks1hZcLl
NoItwDmT1Lr5CBWdzbiruh44aYitTZdiasieAwIiO0+OhKNSdPn0/RLyGQVsl0Mt
z+B7sjsNtA2TTCMD1f5CUALmCkbbiU0vqbsqBZKl89vv+KWg/X8wp96FsCnRyPn9
KWtp6YZHJ4fayx9AUFo60F6VSh5C/z8xLXFDB//IezYJ2bKOB4I4sc/K2ugvoeJN
6+pOBEqIuAQxolgq2nL85qWjN371XM0ZvKLOYKu9ZF7ZFWoKviUFFnXEUcBQPygD
BEosgM9XL1Kc5VTjUjnoFO8iv3R1Zv7ARkCg2P3cRU7Gkbng+L/LNdmdwcerJuYZ
Se/DyeCXMTUvaFuNhfqUKt+F50kxN9trpxNoe8u53w1q0YsYU3Pnq3yizmOBBMcW
6u74HRU2hEwtAQQMaRKZ+KTcSeeifMaAypqrOwNV5FoNHXYUAIok9KDZhNf9ZW9S
mCXEtN2UP9olJeysf4QjYfQ3IrY95w5VwWuSQwWSohCmU/+3T0ni2tXaKk4jTvGt
kTIkoPeuHAjEWHErT/gx2BBHplszpIXmMiPvQaSQbXXVRhzxO6UNhQWlish1A2CX
kFgrm6t5wFe7F9+dq7j34MNgASsm4fkJhMKHnAtUOOYRG/4Xn5JO8eYR/5q8l7fe
oJSfPVAHAfBZLvs87oDfN4NnVijkUrTb35oITxkmkg8tKR8gxRGKtLaKOz+dalWD
ElyF+nFdNq8JMol+IYHT5veLSYCoHqR60XU67Q9HWFOmPCzcg4glhqycw2OmQ52e
saMXH/IzgOybmmMvDCpgDTl6SllPerel2Y1+/jGW9aCuf7kbxeJkyJ6QrrGSI8Fj
AiiYT8Jbfaj30nJwxaLrBz8bXzkgQXk3C238hOx0vd6KtylKLFf/FJTbFhU0Cfrk
NQYuiyNFlN1KVW1Fq7i2CjLgoMczdwkOtHkcj1tHsUhn2BXAxM4RKKK6wDdDF7iZ
oyJdt1QOOQW7vdblyerVj8ZQgSWEH3XTGcXTqMNtMqoI8epjKwvDEPfma8yDrP8H
9IttnHf3t39xtBWX5RQl7FnNSLqAV+AvuGrzxHwurKtgOKdnhQMS6sAmttvBanng
2oQjlhDyLhNL7Jf6QX7QLHhwrsbDPXkdJV8lu2Rtikd+FetaxZHZSWVsWHuwqOZf
WDKs1F2MJKulaJZBY+dofA/U439qUpDG4BvATR5UlhM99JhGgrUH6VlgRfC5ZsZm
bKAqNHf9y9fcsehaUh1KDX78tPREITHEA2X9ge1yyDaFzqxXUZw9VW8QL22J9IFH
WMbU1HdWIUPuBmFu7I9YVpWsgmuEEeYNQgswwl1z9VTjB+IsRKfR5MAXbuHZHDOD
QK4BwuX/Wf2KfAbyKT8tYj6dMaEaGShboWtI/W/SIplxCrb0dMwZ9m9kI/wbrdKg
h4MRcC5mAX3YEAtoCLRNgoBGrN/ggMDIUWmXJSllWtzPC+nHh0D8CIchM8ZfqbzS
+4zKOJZ28hWQNW7Na2U/4cjtXfnbHPlwEhxZEEY8pICe/GicE7VSY8ItFtCUr5We
s/c1ni3lSxxTcFCcwbGXVMuZKeFaUjf2vE211hN1/Orqj1ez+LAPWdbxO/k5dyPo
+wEffs5ksO9tqx+4/cXsu7lkd92r5cYxNHWVyBLN98CwyILsXg8umRb3lvPMn4QY
e2hROgQZ3/8061gwJR32PlZLbheTnaO3Et0XRs07f59xIVlgHck8VP6ARtr/pRC8
mGZ+WkkWI8W5I/p4Cp133nM/Fq7YDBQCDQlCKS9TWvqG6MV+U25V2UNP1Kcli/cA
dySN1COt2t74ods3IXvGJa2HlXK8uUf5YXgtLqX7oe6xvJrSlOp3dU0E4FUvaMSZ
H1VrEE+b3/RQnE9yzWriSjG7A2fR+Y612x4V11hdGG2qff4bsHzBTzwk4Lupr3bM
4OB4LMd0iJgSj3gcJYhpz4Sqeym1TJ4Z/titYwBOjF6sCP2sAEzlh8rX5g+2XF2x
kejeZXIvNm9f2zCeKRE4v/GBXQPLd2ihL8WrARn9cYbqiXna9G6t/55lz6Pxv3RX
PCP1Glo+EHEGY7QBkk8CJd07YHiqmcIiOvy6CYG2/OUh5VL6xccI4ag7JU/Aiupe
oRsJ25fStgG5a93ywufg8mtaXw7fFwLoO5tilnZaXjXaK26HLT3uzp3sizQvzSlC
C6EE+gSO3hqqabB3DVa3V20uYXkiajs4OZMnhKM4Ee9VW0dLCgs7etOxmuV+bYId
v7fpWFNRj8+6hPeqVCctTwLja2HFxG99lfXOJPmXTk3cl53guWy8IwVvtB7tYwvQ
sZBUxGiI6y2Q+hznj4dPCivQ9+4ncZdbR+Ohi+h3PjWhAgb85L751oV3vl1YNgcp
WdnsA50xl85ZWtnw0ICJIlm3yQUKx0cCAOGq4hkcmgsID5EYd2KlYWtHxJQg/zI3
qtFUyQ/oHaI40jnO59SUlDmpFTHxfpEfKUiAbViPysOQciyqQP2C7qedc3OK0a7s
5IrrvEd+S7ZVZb/cBmNLzqjPo7iJTLhRa+JL2OdNJ9EBwNluVXf34e8l/jy85FwX
AIFW4NYNQf76obI+LmLxhUHcdWx3s6ysCwBsvc8oHO60qlC6XjDHW7pztaZv2rFV
JJ9qmAw0w3Hnk5BkMNBP5t9/e4qBDzIvo+b0OFB2d2X8/4Ry5Y+3P1r1490bHZwI
fKxtiaBv2QA+KEee9qPz1AOEa7yZJV6K+m3yiSpYJzQzicSOJ9ZZ7+DFKT2ibqMG
ZaerhFo5BuVdJjB3+ot/aV84FzXkLTat80El/+Oal7TbSow+qjM+XVanksKD2cU0
QE5PkR4YXaT1aPoo/hTfsumDmmc5lHzdhC2WTvGgCGsFO/pX08O1btAlz7rn1X6F
ConOj7H2umx4J9SK+nXpMuKzquRb6l9WYbZfe0bniDiek3/47ejO/XIyL582J2TI
MzIEc6qLMIgvaOOkCVAa+or2opS2Nf+7I146TbzJUupMl7pHAWBJiUp1sIoC6imW
HdholV4eJoDr/XkPIib4kvvzzcdJv36yzz+Lm+byZs4gNN5aUvpn1c7Ugv20O4q2
DJRjiiI9ptXOj3TER4NXqUudswBUs1EZrdAu/ec4GoMXDDi52E7zBlOUIw7brzzo
lEgErbygD4RbQdZPHYfXaCIuzJiWELdk03yEgK/Nvomu7u0u+MbM5Eqro/oNyuUv
m0qGYjLd20ovkgvkfZzPUcdLo6tr7SQ7d3lz+jEnCteCkJxdoMIOddsCKRrr5Swl
KSnbxyTbtiT9iwt8vxKGYgpJSVC1Jfetquj5NI0eg99fZOnO4HNAGLL8bqPLzobB
ZDa08d1ksp7YACGeFn76l/yVMy5EH23bcMV4ZmBSwHngREO/1D+YtdU9c/ZbAL9b
XO7J866CDBMtL3hN5eix1P4cQ08cSgHGb2IhImlZcrchZFY2Y9XSpo7szALasv3d
lw0VBhcJAF3vpYNluNRscFRXsciQ0b0FiigbJnOSPzI01HmaL7PVLIJO2VHfsnfJ
AwiQXpd6PnxAz7PtLUmoW2EbzwusSEBpZA9DO2GB23UdFJcSssAmbwvrBfCpA71P
MZMA/YBQjMR6L72UrTuB54fwD90zOgXL2PL6s+p08LBNWfxiOzkLb2+jfZSFZw8h
ods9fylhrT6PmcskwGjzh6gdyPNbCEiagfkZO+7jJJJprSOg4rzjHObmUoVH698S
hW+KlkO4B0tvSW7ny/Rqsbpyjd4vaEb5D4ur5mclyQT/UvQ0INg1O2n9Qmlibxru
7+Men7758/te3j2BXloD69edEswPjRxIhATD1PYWNYf0oiHDvloXdmDXEYlHl9Ru
sdbioAItzxxCPp0ndqffYve/wsMplNHtJekBUvj+feES0xVxmTGA3vk5SSLeLp3t
g89i2Ut8vdKy2tJ+dt3R7gAMXtxsdhNTs1BBQQ4U0pCPXDAL9ebRJUMQM4aYth8t
N/xRwL5akL/byDFS+qNjCKbzAcHdV7+OghMrV7nhEO9CDbsSdIPLzaqLT7faZvD6
BFvOm+dcesHK2nKXloAF+DbT0CUw89/RBNa5Ka/supGrdq79V7ud1r4QqLjOGFqM
PrMb0cnkKUK94PSEmKP9yUianOLNzL6gnigt9hwXHTsYYFF0M8m6McDQg/O8x+Pn
gd7rMsgc3TIoqccHELx2l6vAFdAvg+in6Kq3KQumqRqFVGejtwS+P/MdmuTog7z/
+wfabSH9XzoXxmRaB9L4GHjhvYg7g1kMCSG98jPFd28tk4vb8eLaYHXk6CXxzl/Z
U4Z84hVKH0yPYJt3q/xDAFp4dhPZ06daOTyfVJJX2DmbWvs4QRAm4dwjuZOGHhu9
l4v7bm1/2f+8ZpIzJMyaX127pCW5LwaeealLjw/MhJHwrp5L2zuX3diYvEJMazOm
mkG/yAcgnWRXdMmjT9dlVcCQc+86G/NhQ2i2gq5rzSVLjt+RzeAUZpTA2r8+k2O6
q+rjlCuy46voX1ycKZjUghvHP2ETJ3EZSz+wT2LTkCnzCSfgYfMilwi66HDh72lB
uEUXc2I7S+Yav99kqLt0FH2Bl32VfrmdNv1h7tvKFXUuPOFZZnjyOBkNaQp/CCuI
jesWCTH4irXFhBddaFldiUwXXmPYEQqz2Wsi5a6OXVL9dOntUC8k99PDDmBLqfgg
8t4kWnloJZH37pi1ELzAXFg4UxWmU/s1NtUi8Sf9yn+j9bBM34rAbelVqA/fO8JJ
XZ5Kna/v0lLkkROdxSFx44VD9zOFdU66KYkoB2DQ7TGgW6Xut8M3ScuoG3zsHmzN
0VbgDDXnulRmsg9MzgzfOEuVXnEAFEMocQpJmm1l3WjimBx9HkA8WR61J30H22sH
9cua6xSH41vDCWfFn6QPQwkfrWBn2xq/FWsw/zpWUOuj68G8Vt9XJCwqkIzv92W7
8T7esZez85WS5T7intyHyGB6ZmAtGdNXwCtdA5sVO2M=
`protect END_PROTECTED
