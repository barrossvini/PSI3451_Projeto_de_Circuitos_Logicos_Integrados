`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rYcyBrnHrEhlyG4qvrpS0pwTB2rXzwLPa/py49NnwjevZ5XyM702DEUijai4dzo4
6HXJAWDFhLQ3HdpqpNpmLfKi/UvjVtIh2Uti1IFF3r1t7ADYAsWEpkM17TPxxhmH
g3+9uZLXiynOJBiZzrByXlcBUaUJlC3Xhn3B94ce7qGjvobwZLbyGXj3VEhXHkYc
pNxXeXFjReklIOtOeTaDpQbHD+eHqWAbxSIs7jgsSeXl+pc7i/wv8dtGbQYI6bKk
/cEQV0KY0ZzAFKXYVSAGSIhFhXUXtGKHjnkXTw5usXbXmTRP9PU0ASz40s5Z8iev
EwZZ6kAvW2XTjtv52UY+pPps265MzlRgPTDx56+8w96TvivdHo3kQ3Q9fOCmy1xy
h6FrmL17pDOONlyVwywDnr04wAezZ0IVRf616zfVJ+H2TDiffOIyJFD5kZFJj4jE
e2RmIGTYDRY/P6efEKwnAUCK4eevepN4acMVmSZq0MEMwyC5NDP7HIU+U6WwdiUj
UW44F+1wGcjYZRYMOIM9d7TIoY7Cz28JhHs3/5oyhHBcOqlfEl++alqJxxEJSFIE
CHpYEaIvxi/DC1bPvX+srkjkeOzAMf5FeMQZjgsmvMEaEA6RGHYlJ4er9mM1Q0Ep
jhg4XuKnQojFdN5zKwsFA9NNbrGY/lQhzMDDNHSgP/YHbJa0m0r4f0hWyI5u4vpv
hQTGa4K9y2bjQ6M7M2vuyeS6/amynbiuIWVkAlsbqCyLVNmgvP2JqjNXt1DkxgQV
AsoHxnamC2YICUnk1QBxwbGG7v4WfhSxJ9upbkf5hwTjTJNJkwUqJryhr2fR8436
Dqj5JqUQAVbjllvApAFrUFx0qIdVsrofS9ZSvAL8x4d0H/yutROMJ0zmLCLRwKw/
mWXYseHfPOUCKNBeJkBX5pnD4IqJNoCZ6j199CGLc6YOpfZtnjdyfP2TDFoYL7Q5
YZCha+IjcG1HzhE3TktVdvPHkUQl2LJFwa6bY+oJ40FpOl9Bxclrt4T1DwFsiBoU
dGQXngfAepby+hMISB3ezKC1k+nef/x8HXJ5Fsj9kB95rTOUtlz2/bcaUdNaCNv7
D0Frpc515ygAznmt28Gaqtl7E6zGV0a53MHzgzYAZ6fw+aFh5kb9hoN4AbV+7pq1
atZMp/T66bUJU905uklIH9Kh9OcuBJxAfg96FxdkWaBwYnpazBc0F5cKd5y+tE9x
RqAutPAoMCXsC8FmUROhpWkbrWKLoK6O8IAn6ynztk9O296G5efA0F5emRWH3UWI
F1dmwuZ3/ieITTV4q1rKfqLcBDl/SeUu2CsdV1rpbwoLcAz4UPFeHD/ZzUiH1gik
8M8D5UUM6wV7zR+LamKsFmT0ZQ6XpRcJg9jPt4ibqLwopa3QEU3c5S0crn78yyxl
NA4UIAQ5K6tl2qAoPK2KOCVvGsijQKEbvW/bdO6SmDvbLAnw+BIl3FGoWP4Tayjm
sKQwuiAMu0hSE73XTiJTIj9pUBmMkoiOiczQ2hlz7sIa2BSRuAOujrbFNFiSZyAg
KFiO3AST8iWAO5H3A1p0ayAxJD+OaoQjLcLCa9K6RrP9zm17fkDW5KQWPHXsNj+I
9HU9FxEDzse8M3qktRJzNHVAfGBGuTL7HMGFNHSy5M3gWQk7APEo1ZQecVbgZLzN
3t/LtpEf4dpRvTA++hlNO82Q8yFwWpTqulMi6RCvQJXOCXyFlvKCLLtIJlMGHjxM
DouthJjO2LW6UNEWsj/zgZUhWWK8gd8aH5gak+LJdKbeHsBRIOFIYJ0YtavRPJ8y
ZLmWhALK/Jqn6Jg/i1iGtJYfstIV8XxJ+XgmcXg0a7iSYer2DHJY3sMBpdRdQfOj
3DO+d/iqWORwTHSyjdCDi6iO4ajafmLUEizQgtnObKuFXfBBD723ZcSKeRACBM/H
M826C3XSQ/DVjGo32boJIadrqqwF3LqTRdoYfiPozt8p6HlkIiXuFgBQlOpy9y4e
p4OvqsPl7W0Rz7M8Py9D398HwdEq/9FNOuqXTsl9riV4UxyZN6151DQk3uYkn0i+
SxCtad5i1MSIQ491rWCF+4CQpxgjUFhSldX/1mp9OXBlx0x9zFFq2O3J3BYXqu4d
/ktYMPLfVDzTZhKdYbtxYFJH82Z/MvLhYFCuMNn4FziCU1uqGBcsgJFsvb2qnW4K
3wzFctwkNiBjGUnkY3iq65fVYsHZGQGzah2VrYXzaTcevQ3L5aleSj0I6ajv6DrU
/EM6JhVow9BYFp8IAHhh9GzpZJwXuWwuYI9GZnMHpRTp3WzSKok9y6fXIBGKP3SA
uoN9a70CbH2TQHO9EWbVsyGiUW9qhyeLo7wPxOVnqXlQA/+THuz3tTj7x/Bo6Iov
NyKdc5f76qTowNTrasEsfetZT+Sz10z9CWRVdwwffQgCw7p3LDGQ//kpxNaNo3dy
v/2fJ4w0Ar+20yuzhcQNloP7zNqA4tN5dvelZ6hZbAN7TqIpwQPO0mfVDE+ZBuRf
LSyWYfzOyu55UPIY+QEmemoNicpfZun2h/NGPsQvRcd1LwNUreccZ5j6041fJmvo
TA9nI6lVOr+p1zsns2Vsfe1Cq97BarNTDVh8AmP0ouIaGwxKsVNzs2sbFFI6gGg1
s5XCNyliQ+MjF2S66hPcp8gXzw0m27zImWVzEV9cro5QH77SyQxKEb3y0qiWM6JL
Z3YWWeRtukZH6rankI9uqosoNauLH7AnsEtcbkE2DZd8QOcK21/eH7wzrIydzSVX
POAH5Rrh2QdiVzNOKM8kDV5m2boZD++ftUY0IegLxcAObcKOtFYY7XwnSVV2RAGh
FdERn0c6a/gHAJD6eT88uxXkbydi0kuWJnTVR+wx2qgcpY+z2wjUr24EZoQ80tKE
0dN0phipsejzJpzAXKMNTBuOpV6+UpfPzl59olzYlpwAvXcIi4CVpGJzIn0P5klr
NJ/CqqfSKIPlCnRH6JRkL+V9wiG0XVRZgecrRyQSZ3++D48UHeOUfC1RqQMmMcRe
eJpU4XtqjmyQthLpP4OUrIB/9b6i+NUwKs8JTflZikJN3V4VpRPGtSnJimWUmdRU
ge45UcjxGARgIocrUqTyQ9cgvpmbML2AQs23OHUtSj2a+9DgdvSYQyGGTtgvqCUw
yEUkN8fWYSJ8lhhm5ZNXTO106ZxDtNxlsVjyGBrDqnwBXvXhaAUFWx3FA6HsHFjX
xbLGGpuKpp0BTl2f3MItqSn2X4dnWPycX+RfyKguHqElWAUcHKYsIhGiMNnSIH8u
rpsQEZyBN0rPmW5FIPywy775Q2sdNuFHKi4J7A0OftHW1qSx5Xmmy3LTQnw803IU
SlWgwXMd9Kii4R67TKwVleuCbbyRlFHqxlJ+HZCxPQg8DUZb0cCxboRayt98Ag90
WZj9CBg6vrcJHtP/etco/1lpCP49gw5jkvFHKzOAMfxfRLIJOFs3CSwIahWq2c4Q
j+Lwo/bAsX1Elaa4EmEJAthyEFJUwWLwBjhjEXVm4c7KxY8GaRLDUwQTAPvrlZta
6NOveQP8eMFi+uyfxj8exWHmzZhXs1vuh0Gvc2LHS3yErp9RfcpiEyR77F5x3v+L
fj/qRLC0MVSExdlT3k79ymYa4WGXIQ70EmyDYz2FSpT4z/7SDyKdfpOBqLxDmare
ZZRdR01sTklw5G6rpMTLJHerre4C1qlWC+Msqm+zVVOZJ2xhXmvbQTMGaUoHSKMv
fGzulOVVdRiYmIxiT7j3zgXrAWmOT8fYQVjQfuP0n+dPimNWggDlCQm8P59DfjHz
tKMgEdzn4szCdMN49NoF2aGmE6vAgEEWHzryPsUhoeDkKWwNh5EWuvhNOic05hNR
YfyeFG9b1zTiAD8E99jTzf6FnFkrONzWHkDg2zmKs7ZBuYj7E2coUxl8KtIUznAb
u8nQ0OOBGO6KMfuwKzoO8p9jRTvPmX/cMpv1LoUSl2LkdXvFN2UgK6cMSBHXafyr
y9pUU7TMJTLwhejKtHvnKD4NxZ5w19u4bwvgIPuWFg0+tYK5qum6H5D1WBRiRYQA
+B1MW8sc5tP+BcUcfkXqHhmsPRYy0PrElCGZwwVC4o+sgznWZYQ4ffUeao8aO5EN
nIicILwUkBkmag8RuomiIHOScMSFLz0NzQVWKhs3V/ze3HDpvpJ1WgWoklqeRp2J
gGapihvpbnTHXQ9qkTnTvjmGTmymyjKM0ShYC1GqDyjOpGh+WjJbEblBQHV3Tv1n
ZZXW71mGQktYxMAMxR3lxtUUlSdRWp8LIUG4KhvdWpQzvAETF0cMdiB/+J0sU+lR
VD0gDMIynmxSZtuPjcmiaKiuoACjDsBLbs9bNquG60MYpES9iJUOJ4wdbXo0KhjU
XtNr4Fp/bpsesxB5gl8rxcuqXewyl1zaUwnIax+BEuoUWt/vIM2arrW6S106TroZ
Uwp2NDJtxELPfXICvPwC84xIRjrLOwiuWXZVx+W4wWCFj56esIS3BzwH791if3G7
BkKgbqbsuMawvMeUt8okaTr8C6TUZFx7SicBS1IS+TqTYMunlUPZn6+MPbeO11TJ
UNKmp8yRUX+jNd63/3enC4/nEEQzgBt5UdTTcfu/+fkOAJMhqgxuIuyJ+iY/oU6T
pvVG2dugCkXapIXvlg59oNqe8DGqybZEwzIyjovVkRAg/l/lP04zIR/GExZa31TN
CKr8pbFNun6y7Vu1CyHSFbpkMViho8KKERflmYPoCT6Q9v0BEDQQb93MQeQ33Isf
Ge84y868QpbJYEq7GoxnIBSRi8CIeWyDATcbY0+SomoLRDQYanfzJKw29DbjtD6I
KzxVAlhs+Du7zmkJDExmLasRYDu0vG0LkxzMrWnw98URrPCuq5oQpsTE6v/6pbSx
LPUyppTo9cN/YfhajpLNhcdYmKcZb86LYgCk7KEKJKUxVaNlfmE2fwl2Bc6dYw8T
LwTA5WFCNwWzWVdXt4k2S2g+IVY58A8Ws7ERFcTo1n/gkD/oZI9YEWZ/EkI5OmLH
qOGQxfOqN0VAoCC1/Gf2urC8lPvABSc/tCS2EcmxX4mD5Agpv/YXyJ3lKRA90Kw2
1XOQecaTrP/N1X9p05h6aHm8687XdgtnAGjjP/hQTWWl4sk1wOLbAZnS+rBTBQtP
7g8OAZAhL26EltUCnaKSM4axCM/a3wUNaja3lvhvGSaJ6sh58kK9PTI8O3a5fnpc
NZcEi5haILiwqcfHX90WlHA3jAxsmU8BdjyuHb/G3gvlgSxHN0UoZt6+vBu+wJLz
BCJvs1MEzzWf8PlJODqRemy3UiBAeM//1/fLPqfoULaHhmuB+nNRZczDQ6qf+wqN
T0g+Fj20Pi4NaZpsKWk3v3dU9n30w1GFu6x6t2fsszsWWlpA8VnJvKelwbvFBptH
u/qIJvbgDv6Vj35bFpmSRq39YhBN3PV29tYaCze3FXJZ/lU3qDm+0+TSVUg+Od1L
80QxBvGSfqmUTOhIZ8ALEduZqEf1mQ8VkhUcOFbuFic5hUt/ywwzy4pUqfT5GZuq
8fUVn9M0wyMJMVtYVKlCMO/YlES4S9Ol97gm7TzDt4nhVo8XkCNoGDAS49SDgZkd
+1S7ZfhVUxZKH4G0GdDMHCP9+8w71TiF0oKnuGI5AQGgr7yqagGhEtgfE0m/JX6A
8JtAtaK8vjGYljrEjJKsv45fdtIXmarfzgjJzwlcxwkmF3srofUhrBTq/1usqaW4
wBo11bODSU5y8kRWZEVUdZwtVIbkgqB+wjAoqbBIp7xka33DMZivyfytDK5gIQmo
rIJjhioJonS5KvcP2fy23bWkiy+zi7IEw93Ba6XSflxUfShqCYUAUIK4mSqqFjAa
4DRn8aECbufbf8CVeUCIRdGTkq6JzSxfbBFE9p8vJIYv79/eJuDN0AGf2476P4BQ
aDd3erIrBuxuXHZPnT3Dva1lem+qLZJFOlpv3Fol+iAo5tuMJW8FzGV8mN6ofGuz
0FOw2ix028o+Jc19KeWADAtQeOduuu2BZBNPMmj5LRmTC4X4wVC9i7JVPUoYxdS8
RUZZXIOT3Bk+GhiJF+rDXM6o0GbyslAaN5LHIesT3ZWYUqIzrkMGgVq/bYFm+yFK
rvrQHY3eJLc6QiH5tKTBPVMUDDO1cRN/3zpKuUDbqMZ29t/aoeoAdlkOqB4mxY6V
wmVH34fq9GIvOchEyOQIQPeqnqaIcoo0rU2yUvj/I2ColA0fGAx9EBw3IvrfISTB
6/cUm4SFjfN6L1z3at+YCFQg4tu0tWcm7rfkv/bFncg7XQBX1LZjneUJ+wjFLQrR
5SlzcwJzpKOwfdBO/Q4bgH/8HsLJKIHB84f3rRB5wYvNRA6XREyc7pEPFggx4MSg
1tYEokDOqv4g/+VMDz1BgMDK5YNeTTzqzFYgDcm+YOpKyDY1o17d90iSwkAx0dEt
RdJ+xkbqnd/UUxzlD2hWufXOV1/KJQ8JSag1iySmzhfYBAA4uzABysULMSoMooaN
pay9s4yUiVcVbr1OfPCl75GOfI4bt9WdI/8P/+HwY8qcorco6sbxZsglRm+lQKJ7
INn99VqB9AYRBAkQYh0NJoy+6Qasv8XU5OW5GwftHC3AVFaLlK8mfha5zVZppxBZ
L1F+CRA1NnsSzPF/VEuz65iUhyMBTJDbbqDz5qc4B75OlsjMXUE6pghFjizaVtNa
E2lNo76BzPvEJziuai6zes4uk0Xym4QvY47CohS7UBlp16Bf5AZ2EdKTIraDgmx8
oNqFkXVLB9K/4tIW4QwqfbbfLvtNqCv7B1yG9+Olm2yFW0IhDKluwfzrHhLiypJz
GO5hvC+D25Qz+0qlnJ97oA8pOjFY1wyCS1XsmYLVeM5iRj54ZYKuS+X+XPJNhJVa
3gGKrFQnaFRvazJw94QlwWopq1WPRoz96R0Hm3OYeg+0JiVcU3Iza9F+6s0qjuSL
LFkmm0cwppAVmZf57mhgqVLjSZ1y43Chj90p4+oCG18SP6RHgy5b9TXHcqLVXFgw
mmc8QIXVlefreeEmBLKXN8ODITMIvDeX65un6WxVdWSeB/l3bwLR0rjXdXyhRDJl
iDOCMTW9N18WQD6ZbldPE6Qoy0/xhenNhOhoS0IJRV9wzCWWgg2hOXRLpeOqqPXs
mQ570IIDZTLBRSN2CuenVd/TApJPMKgbbZbOVQyVomNlC6y2m1hj/taiahO9vkG+
G9Rfm40+wCfiYf26tJ814l88NqPL8fLfL7rLswh3PRxmYYTYRdkv+X93SWgDkqvN
Q1Q+R+Fx6RTadAZ9EhbsOxbXiBhqBJYgYEFLni7ZhUCGf3VWQKD3nIYuI0IxyhYQ
suddtlwYsHXpaopOVQcRapNIzVXo1eOUreDmvXLP0HhInx3k46utH8ygYIHndcRZ
CNkQLS5T+0A4+Rs9omd6YKjxKYtxBFlJQFDkNY0izz1tPjs0zp3B1EFWh2kREieu
kpdfIy6zm6pEFDdInvkesXZcmBwNc8ZdxeUnjUMP56H0d2r5RSBgpS3JxyhNJICm
NZBTpqOdYCItL8adKS6x2WlAH8cFLOJTFdhxxZ4pk8RzxAFYqG7gVPnkxUBeVFrE
4wp5Yq5eJJReYVg7H3Zl7ydMdwas/jgcODp6qMFd9OeyI0YjXVKFIkQrNOOQYotq
Rll9SuS9jMlVRJvyVC3s0LLL0ztOpsmgF1t2UhvL/eVtINbhy9B6U77cjA0LgBWz
wc28beI/L7RQaLL3SVe0xc0M62C0zZs/MXBZm9HHn6+lfD+al0EQfhJWiT1WGwIO
Skq2RF9Qp2E/FsFR0ouFnYFWYS9/qFzPSHGvhOn81O/sW1zWDRXAI4Iz1DTojlBT
MxezdIH9jhIaNqY6HKgzRWvXS7VaivVCJGVVmDoAJw9MQmzV7l7rH08av5lt6aig
5PKoiI61qT+outSD3B4Ogrc7KqBs0sz3BqbmKldIU2/sIxJTP3OzUlAKQGv2oMGH
8m11CNfsw/2qSzAOB21lRDm0fIwthXNYZt7ZLyBrTxJZYkgvwTlE9o7txX5Kanic
RF5biQ6a4tuH0xvhjLrZtc2Dian2IQrrd5IKa9XMJxJkIJyxAs0QXGXvUZVcDjdF
L58qcqasnafXSpuabCyyGBffvymRSXAN8ddQpxU7/TD+B5b7+WWQ5dzHaBFQAyfS
/tEJ8+A2s/bsf9FtE906hTkhEWQLPH0wnfB473YIXbtqaokbPB8jBcyylEazkIvm
iVhsR+Lbb71liPdKskqW5FdV18rjTbswTRf3tvFukDFwPbGqbVidZqZ/ArV7RV/q
oylIqffP37ovtrUBc06eYgFfg7KHou9JDKlK5A1sp2lDGFn3bc0NARCLT/kuQQ5b
aHDVLBMnyUwwbnLXtZ6gMZbekwpNf+6xH4+OXEBohlVrBGfp3BO8TjnYkkfA9ts7
NyhF29H1DYkNz5AJ/4l/YQunym+/5l+JYBdTjWUbCNHVk6IYIXCda5uYRPHs0B1f
21bSvo4cfCZcm/z2VLlIiZepvuU+Lmg+rAg4CE39qOIMpg8l5weKitiFljNLd7iv
0997VKs+OrVVL0t3/snpGUpNoxMfda+bMJFFo5wSB2UoE4plJRqWlted0puNY0Wn
70pPGruDHYxpJspAMpYgMgmJqgZqZPh7EZcpjgFliULwcs9dw7y7CQgcjt5T0m4e
3zaq+RCEFfoo6rC+YY0bLbNOtfSqjUkWZ+7SEAnqog2vuP/vDHeYI3btVRcsPZq8
UuY3uD+bUDMZ+Uv9DWnInXniFCXjRHyZjTXbjEA/RHGcRjYBkZj9ByUE3h7sY2MZ
yJCw6cRMSerx5jHSJX8bMnvSnzcGNFGzSbM8GzdL6bDoINBtoZArfmzOz2ixtKmv
8lQ/242dLBXYFwMg+nMddOyGa+89OO/7pKNr0s68LH06SxLEy2fzYW07O8I0g1rO
px1mENoGN7ASKsQ3/hM2zFj2Rb1XOEZ3CkyBFV5fqTEi5CGBBsEH1gRz5CoYkIMh
CGlabBhPm5aVj9pujtV6Jo50NrfdSxfUFO/t4SplwbOygR5PuFQ0eQGMl1s3E8k0
dkOFc51Y+9wI8QOCf50SujAIiqSVRxoerqK/9Es8GMIaMkVTxL4cXNaBiTYHYBa7
zetEPyV2/LnU6l5yDkNUjeIffa/bcnfMOh5eZfik9y58HbhLOsB3zVgD0vB/XHZk
3Kg97FD92OAvAEgAeo60zwgQ5J+bjBiwkr55AtF8rnxccbFmPMohiBDS5GmCw/ya
9HMG13ETXvbSq1myfs5GXtObiDTSJcKumT70ZKIoQsfP3aq3QRzeNVWBfjQwW93W
RDeCG/5UtPxduIlJBTpidUgKYuGeEhhMIVt4c9DHy5s/6PYon4eW+0Bld6bABcGJ
5lYrVc+Ghcy0smUwnbQ8wKRqiIrPDhb7HrlSaP+3PBBPN3Uq8ZVQx7Fsy8uii9BA
wX0qvVuEUQ6JVMNa2B6SOR3qNjVsv7sIszEFlhzHNirodQI7ges3/vSpfpleM5C5
1y6QNADwALlfvLVFjmtzEk2DGF4qHl1FJd58fE3KValGv1yTthE6t0jnlC331sBr
07lOQ2ny21B44iXUR8VfSIPTXDIM9n0N1B9GtbrzP2dWNOFHIx+gi3WcLLeRoBQg
u2YtvneuFOnaPAlFuW8v81meNVDLCou9hCJ4Cg+orjwvu185naL3XpEOHVQFgF0U
A4VncEPZEQ2ye3ti9U9NyR+vKzEZExdGev/J/gaPXQwLidRTcNy2m+2TltL8dl6k
AL6ajqpnN4nntjW6JNaRxBl1Djf6YcBAGiDkuwrhoJSaCG5AHk2kZg5qIjDiS/sM
cLBuITOBC2uS/CtV9tgEqMCUt014fgyhu+ANcgYMKbn0OmisKW+RExvJAyeB79O8
M2h+bAjIuV0k7YYSaJ3sAd4EIZigCDasKE2GkomfXlIIbEgXGkmhqyjOB4DjsvLv
XQ/byORGs4lBY56eL7XBjottbiQ3EswHMQk/48Pp5uGRndEFe3pfAw74NIdbIYyj
fu1aHjA/R4/kpQ3IdYt7eSpBxGGvFiEwVz3qo97nX9ANpRmRnUPY0HV9j+dEpKf1
h//wARhmwqSJcdXr/7SfxMi/umOLN7B+dXiK+LiRfpqsrGnPVaF5yamOpYOQ36aa
kXN+Mm2jm7kKsH8CuyhKSEksL60uOVsvXzwHKdwJ+Us0RE9mI6Rb7YEWbDex/H3J
jtvfDONOz0e4iUf54jSTiw30Nov0nupsoRfMErl9yArD5OCqCpb4A7kt8G9DTox8
QWIPRQF+SJQjP5ZWceJRuI3k9MjLmJF++qjk4Ayf29vX31Dl10+/VtOh1/ddtmlK
RQgo6TyHeuzC4gsgpElzXVhrJ2Bzvde1PWlszh39ntclcRgxFAnjOjM1XRhxGJfB
lQucmBrHfvl5FbCyFe9pKr4qF/oyEolrYJVf7VMt/UWZIihPcjCsxNUoRFVR4ggG
5NVRKYidGMMWXCz5QTofY8RglF9o07ljUoMZSB4uxlo3oXYE55Ynxq/XUiMqT1Jl
RDleFX3OG9FVkrTHk3ivcZ7BaTxBRAAVosUZxlmUsmDPCUF2Lu80ojw/1aCtzCLZ
Fu4tp8ff87qLYGMzcCS5hkbIsyPsWU1y3BtcQZpRaQtHk9losMZrrtquvuE6qXXk
DD/cJ3KsHD5AGCyx/zcBO47mdOBJ9pyokzfRvRnTiVznvFzHnf21mfz7NPQMekMb
xxmUl0IGb5eI2Ido3nycRiZWn2kV6hThjd197nkUffsOjV4c8ydLZQ3z3axBfGcJ
K4nr9sPJ45yROoX7MzRMoMsTB7mzVCffgRarThfMYSujdp05bghB5kkTptbQCbpz
LacRYwDipDAtD+fZu0MZLKKMxUurNutFmoOPbQsaU4X2yvP0MMHAsQshwN4cLc9g
Jwd0Psk+V9JiaPayVnoiutrC7DxmznEOxJRfu3XUx5ZCAfwmdT1fZ9Q4TeZIJvJM
a2ElxuyamRh1H/FKOPrswLmoQwyqjFlPgz/etqfsDqymPVQ+tr7bnXxCEYIpwgf1
4diincanvOiiipd8b0gJVELYvEEXuzJWC4PEd+epboSX7iyFxsIM0MNws2NiU3pK
ic8NbemPc7HvKYAHRkpJELXOrs+QVwkDqZkqD52V4si2ws0A+MT+rLCf2dyX3Rp0
8A3t4lxT+lcFB2kpeOVMQ/g64eH4jkjFfQenMP/hpcUaItBCwvTwB9oZHUa0uVvT
D1kcwcgpAQhvZBXf1Dq+N0O9Qp/kawCVcUj3RBJku1di74Zcp9O/ODH+hm/Kncu9
zxMBBOw+fRyy9GILDKN1dZkGSVfsnVf/8BSnoLRtEsEOc/uwO7hh7Vyz8WBNtLWd
OiBek7XXU1Al08Os52vFNxwqSUWZuF2ebu4tG0J1DgqjNJyc+YxODy4OF0bnPpLa
VqjnBu0vYZ3uUYsnopLz/WLrOpGDnjFL5DeOe8URi/16Io5VfGBAzXRBqZlDgm8h
5wGTsv0jHYpTGG3fz0bAGD14XMfQfHuffz2FpV4v+ZbWTVylNpG5fk4iRt6W+ggy
SnnZTwF9WFwo/WhUAE7Ame5/4HDvnD5yq50kLcLisNO1W/O4CFmWyPEl+Y46Q2sa
ZEJ4kNG0599H8Jfc6NF54r2ATjJpYRmrT5CBfDdq0iz0i2l0s/+R18B+RvEB+O8d
sZErZBIO1s8eaYNQF5Ij7flkJ9jqoK+KVr0tRQjyCBd/inxRqS6Gzb0aWsg6S7bc
wlHyBqLSPxiqSiSFHO4rKMHXMNTKSG6X/7/V4hjEZfuV+vQzuwddSPcH4/ns5Pd5
3HkeboQUaEWadn5O8WLyQftnTLsLYhRLqGMunEOCGMZzzBccGSbvz9QOSfiiwDps
HkhTnfPzYCGSq68oiL8nEU4gw+JGDb7AJqblT8CqEBQiB+Z6rAOcSxCVQX5Kf1cY
hoEdx07Cicas30Aq+HCSbZjVVysplASR4+bqbJCzbmlOpBFLxR94hxj5RLo8+Wwo
ggFfi46XYwuaVYUzywrv9P+pMFrrnlM/o502818NcfpP1CIhVCe2UlkL2RgxsTSF
TMd/CaffvIEV6Frw7j9gyGDwwTMdCK78A3kr+rACGwVFB/tTv0LheEhd4vvFHM5E
tpvKlSBuAJqtBmiTbprA35rKYERmdd0z3P54gM7pVozvvVzMTF8nuLUwSaq9wEMb
guO/CBN8lg1SxX+2vW9us300HMl5Q64rNIzWv/bqfeun9Lx6yiLJosMJ9yStoTtb
yRWf/TCRbwzlyPDTAXQ6kA7CUzam6ozFcY5vk8FUaCSadvOVT1+bFQd0R8iuiA7k
e5ru8X4EKQ03uOle5tjULr45G5p3diZ1RLgPDGit2sKfYdWVGc5IQO0B6MmgdGgB
7PYdus2IaE+2TtOZysb7WTJCk9/1PDECH/PhBz3XRoCypWqgD4AEZSEiH7KJRyvQ
0LvxfuPzY+4xX1BZRkt2xEK+xreZoDyvPhVzrCuYbjJG0HyQeh1UUVjmIuBQVPCU
8ofQGCylIiouyF9U/pF4hemvw/7WCaF9X9NotZeDqX0k1ZjWd4ZD/liqKPD4k18j
7Tzf2J2uD57QJm8DDjt2ogc975pfqNRmemN0WiEjzCy/gkHiRspJw3VJUu1nwbpp
xnadmM1mxS3RMdHnadP771tj44hp3/Mp4xQlAzjTMesI/6HnpgKKSgRprZda9Ta3
D+liZFcwvPaBWYFhovJZaXzp9tfvexBrXL+QRmKN4EjTths41wmIVNhqtsEaOyXD
0r4wAUgBm1ueTiqV4I91rnq1Eb+VSSD4p2MPGAVywpgCXTEKo0SA9nN7+LE1HMlc
/1iH5HgICAr/ZPtipML8AweUHqbEfAWHWdAtoVVgwD9fd2wGebN62AI8oF6MDleI
OZQaMsU+bEuZ01JXgsLFOp4U0FQPBjLpXDI8DL1lJRubf5gVznrjCHo5r733eXDG
pwMYUCQ4ENAHLZACVIxFyOx+obgxcXctQaz9y6jTcb/bWkoktWmmlvFmGHNIJUqx
N7KcFdhNI9bgWe/uOkvIv+Iai50qOlpCH2yT7fSforie+OaSv1F0IMIfSE/sNzVm
kXFY4JmAgE5zf5PK8g3z9zU1V+oD0gyWPpEwRSEA1tladHLbfJLnvKc9zYYUb7MI
4sdpyUkapo4jMH9QZC1U/uNJ8Pero7bFKjtH/aJd3ztN6KzhlWvULLNN2ousOjxo
m/7ZXRXOQwPEM7x5ZTX9j2Ixx/TxU94NJDDPx+Nhaj+8NEigs7e+HCQbmiMlydVk
6ECiDQWvx9EgH30jiH5KcI8rbMAuFE8uXdzDJB17CGBc8K2xEqKK2X29ngY4vXYp
c6FxR9XqW8x65krCvkJ5cA5lC76rHYTXpk2mcZ5qftep37W2/pqDG9+2SGCM9kKl
8WaoahCuftBFLuP3f03xisFxv9ug1/6Ux3w5r/aHIrqZhrhju/6SrKSLNyxDguH8
qL5vusN21mAw61nyQWx3KE1eGayVagFnvuDmR3rkbgeO84SO3ey/4YW2n1TNq21m
jAMaLk30D4e081l6TztBCgsB2gKCkunotQXlbtfamWdGMhCSYbliJtUFUgdkIbEN
P/MfYiYD/xSg7LnGy04D6/RuvuTR5MZg3YZwy22H+HZPShbbxEO9/NXx86v7cnC1
Om11uQiUzlqcMcKphRKbVnQEjwR61si3Hbqabu3ND9i1yzzOWaF3H465HbSiscmC
kGD4PLEWh/AwOBblAyFc80I6++WGeZG2Eno56qymBCiDu80+Fu/6eH/ffHd7u7G1
ZLs/dFL7wcolGswVUzuKsV6sMmqYz3gG6BByIsxMWtzUBf9fkGWnuOxaTI7XimiL
BTmnOvdCTiFXRVeP0bS4rHybiqcxE/Yk6cqDJDUU1lB10+yGoXmaGB+w/yLM0rVQ
nCy1gyuhysAMC5266v8Cfi5LCCvqiNOiiIVvn2/0Dxvo9zyZdCq2iREr/lpFbJ2s
ADpoxOH9LH00C05vBqfBEfy82Ypi2wZ486esCrSfHuJ57fJBatMnOIKs1aRhttUq
Zh+ZpMSwqFTc5AwrtRDXFkWZ8vsxN0n7SpeXiHxmvqc0/DumWr4lh+k+NQ6ukGfO
vNVws3b99vbCozNipU55DUaeocakM/MEKFHTkRxxQqzrjWb+1JY5CWt+S34Yk1RT
x294KAhKUhySg0d+1AGXdJ9mapAEGAnmSJ3KSw7Z+r/Ypb8P9JNPZSiw+GyukCcZ
TlVGTHCIfnfPY94YD6aJaJn+VsGhT0HW/weqizgnY6MmHZycnuDNbXxsxjFP74WC
pNyGscuKMDkfC1UHaX/suebxfhzr1NKUyD8Ps0wiX/orgHwWwfZsmJO3MXgCgHfF
lAHQvE9g6uq0WmtlsHe8s4D7yC9SNaC5DCGvQD5sg67CBKfaQ3qU/7rbEfhFlCeT
cP8F5FGc3CruZ29hfGfS7z9ZTPCf2/YyvLmF2Unk9jwnDxXcmYFP4HCaezLL/wrP
k44IhqgCxdf+ZnMbmBjiveX/QdyyPV9aH0Y//noR4qfOBgHyA6VLvUkFnw6Tw2lX
BPh+i/q+8A35w8D0LYRnaBv9c+KcH4yo6dto05xNJl0EtBmUIBafBA2mbRTeDY+k
NU5MdpUzQXF/EXtxZCW8tKVWXMicpe6I3DTSYSmWSy2Q4cNF5Mr7SfH8InKK7NLC
bO4dIw6QLEN2WXvfvLbwh+AAZbwCDbkHJsqWsj3om9hgs7Nwd5ffsfPUQMtoDiNy
JJkyJrc4E3uWpIdfuKDR0HtRnSAhnZ4Z5yUInxirthS1C5XiXy6YfFvhX5KtI6m3
ywWDABSSOR0I0MUWg13FvVYcnjfk/tM3yG9uJIUmCgkdko++HNztrBY+gcl4UxKf
tq6Q11gSxZ8a2kAIu2JjQVW4baPZO8tmGOgPEuwlNQVVeo7GeEUU06lVBI3tvb+E
7cXmF2y3KCKDBHhKQ7LK7R7nPGpE2YxzkrshM6B0oW+GPd2mNn7o++4odbA2BsT3
dG4+7RASDPSHkW4gWe+31Y+jRYrMtcP98l+3wYL8IIWzSWMJxRvFPBTyFoaPMmY/
67fRJvsWn766AXICPHDUArpqI7VFt6nCznWRQvZE8ws0cybQkxIJKR24kwpEgC2v
GQ/IuaGAQLX3yAoJGT1kZPwcYPFbQyf6CAnYA/vYWlbQ6RtG3DnU86cjTxzf3io7
f6R2oTqzWg89vAPafnLjYBds3a5HKUYHrK9ciBUZoEwC7idf9Fq90n/nxFTKui75
5gOd9Klgpj9kJreXCSH0afXu0sk+lNI6SJTGMSC2xGlFd/X3etsZt9FwiU3UgHT5
LPPhykVXMVrLpfTzx3uwAU/4/qNur4CYeCTeKiF1NkV5b36GGAL5yBGC/OrrzHJH
Zq72oEdnwb+YUCTeMWlCBH64Ej7d8jxhVDwoWGjSsY08OpSYemwC8OTfMJWherRS
+20OaDZMaMxfouQUcpmCPf8VqoJB6RojePJcTrPRf2zW0VGL1jyndDbWwVV9h0XW
Em2RCsyy7jcz7/xPdW7CPxZovffjmeMDDDmmb6XXsMg79GULixPk9E5nw7isJmOS
i0B/ezefJJZ6jJw8B4evNhj+HiwKhZc/xTB96GsSv6NiSrD+a/pA6wrDosrVOzUR
LqFLQtGaFrOw0NE56pW8Kyd2B793kJPlABVr8Y1Tak7Bms2wNnWQeXXkidxpJIoC
JJE8uG81yauR+urtjlA1neLOG08fh9BdZliBSd72RlPR5W3DrncTd5X1SReUG873
kZSgZZAgs2m1RGvj800RQp9ItRVsKyq5FzidjxUjfxkcvU2oShgM/2v6Acw0PpZC
pxU2FASOZL/0xBi6ULNd+yGdvpPsjWx3CHm2bmOtRSjc+4ThY9EMT5KcoKiYRp5V
28Q7yA3Ly9PGpx5k6kJ3tCS9yQeOANPLRbRC3jyY+spMp7xwXgoEbwqTstg6dJLb
S+GBpjhxK5IcnDqlF+d2w7iqIEH3BV7d38FsDE7eXDxsiXvwJBoMgB5oXbm69NPq
Z2/jzkeTtqmM5S0osYDUEkGys4YHDCKutP7FxDqgdWvqeSnCzT+XUbQtWcjXtam6
KMYTv7RNPclweQyYMW0I4mor18tGJ4rGSmLzGUyGmy9M2jNBFL3suEMor9V3jquH
NKuskXcQESwRlBS9MAEcjg/iHaNt2O1Q2xSnOBJ/3LtXsE/erMJk+7+NeBA2SUb1
xe6KVbqMyLrF4EkSDJ60ebmBZ4TMbU9evq3OQemgAslBf74UpfsuumvR//x28oS9
wRTmpi3k/4U8EhMfpXLi5CRLWvg002mFYWfwmWPq1T/TjB7I7CrzC39nxVWK6nDH
lf14jn4fGpsc2vVKNgwldBDbHt9oH4kZUAT8cp/hE88mrgVS6nGX1Ig8LLIWKzjH
DSbJbnXA2enr8h+qQsS3avVSbrWP1WqFbkZVhXCZFKMD2J3e8g+hdGvOEhbmEp6u
rXX4o6ZTVotuaUl4+SHYrF3WMAW7jElj7f1lnqi3HmUokfFoC4o+s8oyWkAgrW5z
E47kib9wjaHJsY6R5eU+EcBX4FLtP4Sx63wnkyHmTbLBUBz00bAOiQWvF1uWQ0+R
zQmW0kggiYfSPhWbP6hFc2RitzSeg0vtg2eN1/N29R5DDM8sFUmUNY8Jkkt0hJyY
SSIGkMDHanx32kT97dM/QX7sHbTjVCtbNQHi5jnmQfyiHNlUmB+ttEjE77gJ5TjD
9ma4O4MzAiiiVBoHktbj6hrkFA7j9Lf51zznpe+y9l5jd2BURRqE6ME+jC3JaMr7
fuR63cQ3RybOQXNeEGdRgvQg619j0wmFQK0UZKwvr8FlfdK+sP8xmVU68jM1beIq
MHI8ST/BNCytEuLyzXy/wbbYvYuVgqSqO4v8oh6gU1Sol48V7GcV9Q+lOvHtckLY
P1shA1zW7YFcKyOyDBfnJQaWk/6oyABhfo6r4AAzMpL6wgsxC1n412WspC4Wr9JU
gQbFZzesHH3OlJgHUChcw9sij3Ce3LkURe435ASTJYCFLYl14ybIrBEdLoH+02OY
B5sZbV5l9PnK/PTxVSR4HSExvXYViYHqjz2HBU7c/fZni7LHuV6/0eGI/GHyjlOm
X0UNPt6RHWa14X8qjkVzXP/3x5IO9Tg9kT5aDvFBRs3uzN2dq+lJNRxtS0F/oWMc
0IOTVUceJktXyclddT2RvHUSUyAZtoWGvTTn+Or5qiIJ7kQybr+zBUIn8bILtySi
VAmp7kpyjFEsswRIb5rU2RgDjim8mOZXVBN8KwFTBll46dga39MdARUkQ7EjfoVB
AAbeAfMmOWaV41yItEQuRDvj1bRbi94ElPUjBymQe45uBcXgLoeqWaOrt/uJhX41
3tAlLASbKOVh2CGGHf/Hil3T89yOktg+7DNtXVzMZ5fgCMJWYREcpek8enP/eEWh
r4v0vXPFvnFUShdhqGZ6DsZP0/9n/hWX3NEyZklalJ0Ppkz7GTqJ/vdUGmxw7NE+
5S5pRV0LYXsPT1Rjj/dWFmB/YKUbpCcY0p0qtGvJCpwOk0jxKkgdOh3wby8s9kNe
aBEMowVO1dXN/a3oCy/n4cueCy4GrtSC7e3XrnDBMwje1L2hST/sSJ0LIFmNSFs/
Hvjb10pEDYQZLpV06qfKY6Vcsto2l/KPaOxMzDbtrJM6M8m0W51/gmmNRHtHPnby
/U0xbZZcZch/vGWj06VSbanBuqnLS3jtagpRWitU/IDcBBw8dAsF6fYD4m5guFmo
hAPX8eLPj9T+g1UgDKuXqmEdItbR4AOj4Uy5Y/Asf4/ViPPQJJwqk7LqmEeA2pOZ
h/w/rGwnhjJQ3pCO3yQg9Ui8vxZbfJbwy9paJY+D9vhq3e61kQK8cDRhbSzEKwSU
jqMgKdbUcSFnb8lHl6BD2Ax828zsiwSFYm2SHJcuZ7I+la+NSGf9nsQ3Jv1QDcxS
C/Hi3XY+mNF+BCXYskd3+eQvfKrveRKXM/rrpM0iGzblkVOmcAaFNijf13FbVgwJ
z8gQUS3sjKH2f4XEQ+EFcFWLdO5ikToAeruuoY/iMRwgWqhSdvsDbeJFfOHPxZYk
bXIzQsHTfx0b4FZgB0FLCgIedqNbdDn4ft1kCCLeRjBt/7kSkuD/J38SLcX8X4Zr
HWOwy5hPbkxFHwCmfhlXomud4JKzRWGFAtKJjGt5bDafhgLUrg1v6QanAQxLnfVs
sg1HG2mGFP+i3DRh5JSj4cjFC+NOQrtKmJEuTMFiEdTzpgV+/9+aPzwngKcgD1i9
SklenbXG/mklCB2101BpjlaYCstiCvjJaZ1AVwyDe/vodqjTZEx+m/KHNcSugpQc
56jMinXlsegAnzaHlMWgb85WJb8yYyhZbcrgg7b1B6foUcbFEpfUqrSZb2Wu3z6l
QheUOl94VXaSkC7tlgvkN8ojea+p3aL5nqHabOiO9wiHV4DlDmuPFxxzClW06+lN
HSPfpsVPspaEJ/is0tMRPMiUkL7CVfp7YjvjfalRNI/Ckn+Lua2N7LsMqI5a0nTw
jIMNhYcMotyeNDs/xFEr9OtCFMl/0+vcToK+WmSDqJtWXG9McyJgbYEus6X//jGM
lLzQ2WoZTDkcbDF5+HLzOxNg7DhnrDJ6BgtdTXQgLCm+kMIT6CnhbtzTg0lQGM61
omR2SWn1dzHjdS0g7lYxNWjAvkuwGjbgGyvKMNDoyA5hCVEVhXpOQXjWDHTWCzkp
+N+ALEbQlpfJ1KeCPtlEZ7zz4SJbAYHgDkaxqEIbOhbLkc7LOqPJvPgzlCbXsuQS
uku3h0+6ErPglHUjkBiFY9PfTfuNaL5flQPtaWdsEF/cXY4QIC/UlZPbHuWehBr+
fr2ktkRXppyY/X1/Fa7Vp6uH9Kx1AT13lQMGOyDxBbVmQAHklC+Nh9R7b+OfaizZ
7fmsIimrO9epErmASK7IPk26+hQS1JR0M8gS3KRNXMKFvW7I8vKh5SgPQZ8SLWmr
VvFF/kIkTucZe4pC1RqsBh3j4ZwpBbfDHYpP/XIYB4ctJf8E3m/fNTWzxi2IyfIh
BI4DgawPbAQ4STHC14rPia9ZdAsd4ABL+CGpE686ChQ41OHmJjHTFEweTc5wUUsm
ypQ28UVS/igqpk+IUOv0rtkNIqsy49lChZWloRKpmJ8ZCjDEylUmRNxugYv0IbCv
E1vcZ/+TNxFkfAItRRr7fGQQViM7GPxjXMj5ln3hNfwBVTZwWRCAT06l8yUgHz+z
l1DAja2B8SyuOu9dspW3I/dCkEqYAwMh8U9fsFvQD7YLpzyi2+k0pDuMA/QLN2hw
apueZGwQUcFCkXS9muNAODP6a8odZek1Dxqwt9FWYKqTHHtGRSwWm6bXCqi0lvLs
lLBNLAkFWVpHFesjplG2tfW840HCJH7oiQ9ST6IP+YaC0NaiatibxNstsW4dWPOU
uZ4gBcArnqdCXQqR+8+Jyd95j/2RUbnv2nS9iPGJLRzizSp8djF6JajlNJEV/IE4
nTspnFdRHkHu/LUhdCD1JY8i7hUXAGzI1fU32q26MzdczJjSquQxHzUbNm56T2ze
RKyP2KS9yCdJvY8hyp/Z6IOnxxF27bJcT5Gg1az11BdD0VU9rvpuLioPyapj9mp1
f+Ce+GIIHqdpO1T93o7338NcCDUhoDoC/1C3K1Ndxl1Bc+mlH4juYOPAP3MghaEy
r9Tj6WfVPaD6cDFZrTMlw7lQ8gDzfFqsLUb3tl/tZQy+/gc5uOqqR+iMw0/kQ/cF
4tnxG8bboiu8ksdueE6CioNsyTwveQ+FHX2HeEva8EKJSPpnVz0hEcnRCf1GrIiE
kX6wUz4hP1hKS6Xy/mNXLH/eVBA0EedHlD5ch1L/LHu7l6pWSdTGg5EFXi2FWcHd
sD0q2Lx0q22lq8IXxgMDCvlF0FjGoKN8CeLiLMFQCmy3Gd4dKIkzivN0Mf657vLq
5yVIF96Q+wJj0+xp3omSg3CM94np+N/L1ER52uunnRHr7yv+ztskUIjUla5uTh2P
SAKRqcLZlyYJZdQqE75HCjAvJVtOjqSbzDm0NmTdZ2wDc4E21v/9GJtaqs26hMOy
PqTMI839CGSUdHokzGoLWGAZ7NbRJupj4SOVOJ2zz+WJsjal7qQuUNbkbUhW1F7W
8iTXn2+J/tNXGibGAUoaaHwZbIocPgEqK21Xwhwr6MaLDuEJSuJv7+sSvgbTbfQ4
bCBjwsPjGnV7CVYNou/Qtu4sVV2TKP9VePkAnQZR8x00JsXgdXxBIbSxfXqBOzBW
yHILQoRqc8sAc5KAQyM8wqR6pzWUwdt8wgz6isLl/0GOOlUTDB63EjHz0MjehRrp
5IhwNSYB++niXxdKML6jJzM+hXkh7qQxZmSbA03ClcaV0Hsm5Zr6r55rIodQelCy
Ioswx6bT0I22RtGSQCQFdEWoz0zpSl8HSOiiBk3xasbW1m//kp4c/bLEO6RU0HT3
uSyK2SOtG/jkwNQ5UxUXXWqv/+uTKspeWaKVpuImz0QVgX7C/vsTAn1rbu7gpxKt
xa9MzddPrXqcNJx9bNeoUIst/WVmbFJypSqLNrPHBreQcokEmr9HI3dXademSjDW
YaRZ7x0dje8qRId2OaMFd+X5Wp+qSmdaIsP2XolTzK9kcqrj/GjSpB4cjTghWzUN
F2H3NS/3emWJ+KuUscrlRxh8OD2LrM5aeFh2hh3FkgvkqteaodhQCezYcXV7q1aA
uTdM82CF2mBNAf7oyDM0Z0NFaBH5i9YXMhpruU3Hr0XzjJuLRVZt66LA02R3xGyg
C/JoppsGupJ8QD4u7XrBNOUmggNsNDmAUcjson/8+JevMsYWgotXR0uFjy98dV8c
Zyt/BuuG8hySgLHG/GnN03KZrLiY39P4JtJ6xyIhsTf6zWGuymp+YmDz/izIgtmr
DEzZ5slfYoxGweAlOY1kv7TvdRTNuhStbZ7RXq3M3RzSZJ9pHhIsS7/UWN8+FupR
K/XZUF/vTm9MRGw5fkcKBSvI6HwYUvWd0R60CSPpDRJBDqK2KpKC44usL8Gn5Rr+
+zpFscz522ZxnRSWoS0XqkCYynM8LC1wnXIiB6GfxCcj3SFX6KynAreSimP5JS0H
4UaoDwO2tHVTrvwCfQgc0dOTKNKbhAVxU4FUpgQ8lb3eFrlWr600yr7lx8y8qB+D
hwtZn6eWPljOdoIiPoIOC5Wq6hNvMQgPTRAcWAUBaphZp+b64EpuOfAxwXYW7utK
ntN9MMz1pqrJK4dNSS4uPxTsgZMIWoRWzSAmUHgdt3IMrsgiuhM5Yd02iDBSTDmx
q2ov7v89k9fd+tB1A0J5PlBbEUaRvwaOGbanvgR0Rve6lsKlK5ys9nkJ8Xgd4vp0
/kg2DGCnb3yK6zdSl3UEGw7BZIC/2moWV136/ufEI+YlCWFGO3FPPnumoo79nJim
YmAoL1W4sclE8Ypk2zdPh6Jy/VUBNPVAlbQ2FVq3tfZDbcQPVnztlOgZgb4HgZ3r
37YeOmu6aiZFQZclx+r3F0I/6XZuMDQ+GErFhRsBLnhE86JdehMn64r8FJWrV1bw
e4DzmXaXaXFfEksipPesMX2Ihr62Q/sjktGI2kqX6TffmTOmt+kdc4p5a9H+XIBL
FwrtmpiXIgYDMdlko/zBc3ozJfMU+amInDCXTo7iO1p6aR5Azqe2qZfZz2gGkOIX
xQpyzT/IMpksJlMLojhNLzja2nAhy8PPqVrAhnw3nUSvnM7+0kYGM3uEYwUotu3v
I7eDgwUN55eEeEbWNu2RsHkcgxdsb3RzE9uWPAxrPqtCxDBLYazqASVzOvrjd0Fe
Q1CvRg75ovwg0jI7lBTsTuIYWN8BwgIUpfbJBHmJjGgLAZ8G/H4IUau5viCJgeHw
kAP78AVRAZVi9ULPDYBOU3WWzWahWimn15ZonPglmH31btmPc8zEBcOfhJfJIHLr
waMgpby+J+kMyrWXIGFaK6s+w6c/xGeZmh4LHmhFiS9kThv59DZMb5R5P1u7LoUa
9tmoF9Mf2PAhm6JK0MoeRaryxHTTy9dZdcGiJn5KKA1dKKDNc/eVgg/DoVGT1VS4
8yJQS7fXO1O7kIQDGhNgjUT9qtnPJrIYl9sJCijPWeZ7SFtLaqMiHwfyze+PpbkM
IHZ2UR6+/6I/L5vC5OwuxTKotLAM/UjvCM5LVTpAmPX+wABY6/n2S46jUaxK21cp
BoFQqiRkv569BaUXq7+mDw1mLGpZuPsSSPkYTb8Fb1WcHJQseM6G/0LAK654ztS2
6ZAyKo+PNZRyZ7L9cUTxx5nrlaOJqBLheCZoSRDv/ThtTGBnOlTX6eHhE7siziie
hnvqXIWwO15njEW9kp9W6UL2hj+urcWIoGm/Whm8gKqwdFrR6JFmVOVQkXPUi6FL
TDwr6tezOym93tLsa9yVHPPoC5wCnfzBtGJHy5AR0H/24BNZoEapdD4MnmRmWB+E
boFZRAMVj7U1p0kaSqENYmATuKh/du7O8fEvNm5mpaZlGG5dHER8rm5hvvLCgFOu
pnGLns4N/hzSHpFuTLRUBgCKtZ3ImzkhvzrYr30WqvfLw4ySSLGUjcLUpdgVjnOL
J5FkCxpD2yrk8YRk42ldMuoRRLCudQEOktakg269czSdpTeOr7cOrg0KUuRsePqh
gG/DrKcVCigIqXZZ2gDd1SYiaRQILYyEr/01VLYb04aS9OTEXs8ayFoE0nr7ZeK2
eXU/f5TG2rvUREZauIEurTE3DPZtQF3MMaisdIqmKkqCIOlso8x+N8zqOATNqZis
eGr7VAGSs1SbXIDshis48lhPcL1XLKXb7An2Np07Onj38RSd+0qKoK8jRRmzSzQt
oT3W6WO5Dlpt8ckqVHeTFPBtBFgBWVjKzSJWJTGQFKks0H/MGDhFpr4G+i83VSs4
9Xx2oQSwNVCY8c5KsJCN9t1nH8oQFG2gRBMOstlZdiEIML75TBt8R12shX4c5k+V
N2gyc/wQ1i7kxSg/hWktdWAb6B++AxzOa3vebrxhHTNuS3VGysm1rfwhWsyKVsqc
gXRXWH2ofsP1zAh1CsBDbFrFZ8ba86EX6M98tPlSnXf2DXgdfWS38VCsStMjCvW6
EMmFrBqu3PaeiOTM90h06HbY9LTjdOIODgYuRazJQ54gCcmKcamT9EtJ7pUH4li3
/RbhxPZZ6Rp8+enxQWg8PU0JadGeJdgSu6UMqXxjAgghMnzV1GzIXMpNphFqh/MM
C+4Mfg0Gzgu7ehMjWY+8/cQD597xJikLQADnAOLE7W5MFu1Ra6nnf2mmLWlFuYww
uF22FZkwvE4rfQXJaQePqJITPlqhkpp9ajbzXIMQicG1sH/h+lTkXTWqlP2ahF71
X1WM18YDgMD4jWm3fXs6KqcSClQ7QrOMI3jgH7+FnUeDyBd9AKQUhLZHNj6hBYUc
TdEncCQGm60mmXiIHbLQ/h8BQThmGFyBDjno/auNaS/NP8V20+GroDRbI+m/ef0f
uF/jRbOIXgouJlELpHUG9whX7HBlbcwDeKP2c7dR49Rufgxa5adk0TiVcHi3j3aI
83w+m8rKzIjPlHiIrqZR8FG/N4UxoEAZ8Jgvm7NhTEnvmecTMk3Uwv74gBcHqD8X
G6+AzO7HOoqOpRizd08vK4YUXvsUjdsBowg8LfK5bBMCyGp03opQzwitf0GEF0Pk
lU8IaxUsVOhUZR3yJ/uTIUjBR8sC2ZcFb3jyzPJFbxyKFlitR4P8aadpCURmUFrU
GkE24mLIkpZnQwZD9V5+/P0IqnJ6ILiJ8s06hY39h2wtl7ROuTLarEODiITZvoMP
J1MQif1u4drPtW5NlpaWo1XZjb8apbfkjWv3Z1EZzklLjXltn/RUiWoh6bxhcaYE
XmYpLk+k+GJG/nfxFECjgi4tovY3obbqC0BGOAc8X+n05dX/amjuoCRg1bE7f8z3
ab/UYkN86w1SgqJtR9pDJsHTbFMcZVqd0Y5lDSty0dQUO7WSGkFSdQg1hAtTi9wr
ZVIstNSh+tK16Zm/VfmlYff2/UAZ7hXEeboYsXda8NZHxothYtPGEIM/pPcYHCoR
qqwsN8McnqztRexIY8Dh/Dthi/z5Vzv77WB11daZfy5rMg+CyFvVu54/x69CdbHD
qrMnYAjR6zt5Jr/vjhKvswVfFEnjX8WcxEqv0mlVCqecHT5bIDKWonz8DCdR80xh
BIjR4RWcqsZunghnltis7ZOwVmOF3CIS7bnnZXJcFhxrqXjUWxNaVeWfq995F1BE
APhsjJNUWk0n+4KCGZvlX4o6i4hv3tXTfcjCA61gq8kXNfEwgWkheMTg2BQ4eg12
1QicPUwRwPMQLIqK/3KwYQ0SUmAIRo9pXPQvHZFK5hwC53J1XB6nuEQe/V4cphWo
9mcvGH1Xp67RXQegjp2D2SHDJtGAc2JuvBHn6EylcGsNhZcDy5NMftp+8O6QWk9t
XcoxHShVKLI5clAxsiA92EOayfowD2SFeeJbdpdNpIDlydC0MQJPOZ0X2nCRc/uA
i6ouW/y1+BNAlPZqQ8CCTthjrZYywafKLnlvZzcp4TDL9SP8O7WlJZaX+wX+oym5
is0tmHlekxTprQ1Oxai43tjFaYCQaMAmffTouX7PhH2+TEwGDEIqp+lH6LDfvKX3
YiIxyGsPopzbYCNMHwa9zyAaHoXfRbQEeuvrNgWCvxgjSuWn+8nNvUPr9CyvRykE
VrAQm/+jTOx4Dd3l3R74EGzif71ta6hhNZWKNW+UnfbxfhMnbU1gGIvNK5QpNwTe
KCfCok8aciDtg3YDrO3jJ7qT5iXbnGI0hknqoCxpqMLp5LzZVjryyMqDaiV2Rbs8
bDQhKR5YfWCTS0V/UhQpDI5gJbu+SCw392ejQKJMmGOac8bMfNZu6MG0PDtkXUEV
o2v4TsBzA5kLEtngc7SpQ3NS5INITo7O4PSziAIhFWkCfxxRyafy9fhJx3Vi18qw
xqVsH17p+UdFJdU4zYyx6gxVd7PU3IHr5fJ69vSV9aAAdfbA8aiTewVbsuZoNLpv
u7r0iAjfnSkSiraT+C8Mg/x1Fuo88bGYppJonWtgeIiyYqwjo+CxNEcZGhcw3CEa
bJPgZe4rQwDxmdNrB3CNe/vdQUgOHqDzGosOC62XJWkm99wqTkeyF6ZBQPzUeAqF
j/kNJx1RxTbcSAV7JUZKPLUr/JUqkHpLMTv9eHsfS3I/unuk5J3hSNIyvC7hMs9H
GsaKZasFl5gxYyO/B+7mlFX/T1gGT1hsxgCMkSUGDgC8ij4NLd2JfZHVMASwaUFA
Cn7qmqyjwoOQA/EAEHFZIBx8Pf2AKK95HyZL1Nay/qiuSvUn7mCn8CPWidtNz21l
fJRBdt4mLMiWCOSRnfxbM0E5cE2BtnvOo5H5drz98WfT7EfCkzN5AUa1WA8r6t1O
i2zqjEHM/PCBPihpgyGWJHSoRcC+yBAJdO3C0XFsRLKUWpAB1/CMPkqlsA+cDVyY
A7DLgvJ1xDeF884aB4kOzcAOxc4B4Nnmvh8BirivdX6GFUVqRfh6AoOd7dB18vdi
iJKQg1vgTh0e6K4rT/4auSaf4NWzO8qahyij0H+udgzivWLyKMhLOKIA12h4xZrz
1yFQ+IUoM1ktNrdnVnZSAcBJra17du95ushcMV42DoG8Pit6228Y9fjnZXQL7F1D
0lm/RPCnMUfSeeKUw0mRTpKCVy7lcWJBS+E7t5bS3cSyK6UsiaKRPHiN82BMb347
j3puj0zybA0KkEGgA5gdwfydE+VG/4c6l7MWSUR2yCM/RWeN9I0WvY+N57kIct8h
BqYyicaEuvmsfzVOdZx8cvJBEwfNaITQkHwe9dFqIKDncagv027ult3rFAK7p1S5
QUDbRuZgnacz3G4AntC23F0lcyNePrQbykOqJ6edKE0FB3FUgqMGjJv1dOAo+9GV
AckpWN8zDRRl29vanGRFxPdvELlntcTWyr2jfTlaLxhWVn+iyPYNcacz494Vs/e9
muf6S7Jv6AIK56cBjdNHLujiKQeaekGzOKtNJOXy5cPWHagp++JGD58gbeUonSbF
pgfGQJEeSHO1KVlm+n/qDjarx+Ezpiww0AFbwKk3JaipAJwEIL20iL2AIZ2tNc/4
kjn36wc9HFXWPn+zDIOuTVrYuPkp41sQq5/7ZH2Cq+bi/Jo7yMUc9QE+2ytgABPM
xmcw5P8mD4MzzEUWjIZW0dOLa6Rpr0jl7aHOLzPNP/akw4pDkvzswW+0a0eTNDEq
nCLpx+S0tazBveZOweje2jlp0DBUSMkhuuDu/fn1aOj9H8VjnAibIdKW+AYRh5Kc
EAZYhCeILUWqTJM5vQMWa6UewG7sn45/hKkpLPmRGmqeAmuUFOiETD48oldoJevK
qdyF0psHS08ew+rKX0jN62l4Z9aGqTjewH8RSovqWINt7+00BgXiIksT0sr2vtv5
Owudu81MHVPoDn+pH8UdQ3/VHB63+HiK8FFWcZmqd+rMt5/pct09V3AfaBgNGmMH
1VU9z1hKRFj0mdDE70sID5E04TLSr2J/ZKkqCLkTsZueL1g9ivN4qqZXknwq7izY
IRBqE5iT54bbAx4dcQ5nXR97Ix9dYgwUQx9ymjNhaOnnl7ejmTX7FuXN+zuyrHRa
4xkC9KbWeI1zeh1ltks6kx12AjlBjJYVCbhH0779rwq3SgNqq1cQQx2QrDtGWXZ6
B3Pcm9leamNxGtrmKEV32vH+ep0X8GNEqGljGeK0Dvn3bALiuSVvpnorAY7z0Ywu
6W0MR8WrD14QTYEGU5P4hXTWRJ00JvY0ENuLu0AQhf4k0unSlxRohraRSy1B3VVn
CzuxB2mD7d/SnX4jLohP+BalJJYAVSBI7pzlpSy4COGZezITKC0bAq6mmgWHZSmL
+j4jV6TFXp1tmCMMOekx9BJNk/6AeJTtJZdo528aT/D5pejazHtV+8rqY7ifiTQ+
gVLZlfbn0ZmGWWMdHs1S8ccgD3U4ktq3T2zu/cvI5xsS4nfW/F8LI4Qxz01njmfT
nh8rbRewfizJdRatn3B6kasYAlnDWhsFKsrbN0cf73CT5atW4HiBCht2TZvViYls
u5HxcFTdbe7V/WLkqxAEwgD9LGrh1Ov/hTtHvxkdmH1w9sPYc2yeLSB5ozSYo44v
zJfptpvk059lDcAtczHHzr7ovAKMyXyt9lj6Ktt8C8FrqA9HUbEhRC/X1ewVEMEY
mfN+hvJaLfY9U4ysNopxiCTCmCKqLa+XsG39uF+qrWiA+2/pNcuh4UDT7qpyV0Js
LBYHIIaQGEx9sYP2LDHV34F8mrRq8UTiuhtV7AC7ayktBICyYy24AH0ip6N9g0Jm
26r/gmA9K7pkxbv34+Oa4gMH6jY3pxQcWjuqtN2DtvhlXa2toheqC+e7cLQU8Nc8
ZBWEW6CkrAYDNpLD8joetfPBQhPnLgpRRjKscZkRBkqBdTy/g9zznYUzLMiSpmjY
lED8FRG7wQtWPhajRyvF0LiediAyRnT+G2nOdvY0+IItMspQ5xcXNfPGWzigVQtc
Cn0Oza8lIJjRt5IhnGoZ5+kswKp2k3KUUq+PqX39LZu64tqaoAQfWqVepEnZXNg+
za5o1Yf7nqm5TNqQLc8/1dYjv9fal6G9PGaclNbZGJvmfqnn7DwdlLURMAWpw3Iv
24nkYx67U3rCLs0zRqc10rd7UA8Pk0Ek0uzDzYuw9+F4dMvy7ykYWF/0Fc6l0+xQ
Ww1mEWbAxggoOxDHGoFKMgzwWKRNioGnBwbum38FjOj7yPuGvS5EELmElpDRguZn
nBTsr74OOs1gFm2FPWpsuSoI15glPb+tc4vC6vi8RADezsOEsEAMl2ROnef9AbQc
8rUUCsBGkXQCHTDY22UWV5CkPO/nH273Y2k/ZLkQz+DsKX22tjrlyp1AncDDOfa0
MbOU2N9dojZGBFglVHaAQE2voy0Ru/Mrf6M8WF8ByUZiFQcVV1QZyKYXpKMomErX
ywfAJSHMPNJYkCdJbZgx2+6KDMYK2q7C61Exs3y+/UQbVLrVkKlohBk+9w2/GKgq
tWbJ4MBdNX06ufkMnEei8CLexrV7EDU4LHOPGu7nsdOLswAnCQIm9bYhvPzlNNxd
vzLJ/h8IV1McpNg5YdCE8yPTAXDApamtFErHXpGLxezCkPezPAAeXLfY+WN7WnGN
IRgRbw3Z2rTrCczjK/ml1iZGohk29rbr8eOwHp06laXqmiMzntvNKsIHUYr33xwG
w3sN7XB5LAlcba+68OcCJnwLDkGbqVdGb1R5NfpKXn8HVFqxp1l7kCOeBBoVD80q
/IBWRITu3IgSYNs+RDuo5expj6ldIh288DCyaQvHE00+pfXfeMhMSIm61iwYZByn
hv1ljoN1/HX54G29Rc9VSEkNWjn2eHsH2rKU6pF8pJNGurzB/UaxayLx5MzhOjN7
nTBfZonbFu3Gc3I70VPfY4PHR8CUzIdO6pShK/aCr//7FyDQh/gNQAlzUKa0dWG6
JFytthgxAk84cSplgkfEEmOrQF9lVBfYZg9aIrf8c3ANFCeQs1lUbKbHz7FzdSFf
ER8P5LWgZ16jPwfiyR67AuHZXgcx5migvT+9drYkrC5tvWxLaijENYrzl5wncCWr
wCJLzasFQrit1HvrjFhdhg0VFsNQZPMkEnVNRcxkbK8Yq9+m8tLkCnQPDNBA+cNX
WsdrLV+pKP4gbu06w10be4jAoD5DtGPhkUq6zO90X0JVU+SHvlkjfrAVkp1piT2d
RwhFg5YOyyUiDoI0F4DOGEHj/V3pCp0tmzovvtg5+NLE7z1EIZRQhS/kQJsI0MhH
B5mZR1U2X20ZQ5ip2uVuIhefD/SBIcZt/cPxdBBfKsM8hOJmXNFvUjfqOIAkJpZl
VrpuSW8GExzKcrEkv/bRJBtt3YD3CBElooYz1dIbnIfUJ1657yjzBNbOJAamFbE7
JUzAJTOpmXLAKaTzEQtme9ubfqMQsC1JiDyFxSyhHxLNZ8sKnSpNXaG2uV4rVnz9
5ainzc45bIRr7tvbDk+Q7uIx+mbEhCluhIORCjIcHssjhk6UD50fkdkZGgLnxr/P
e+vWCseU3qoehM4C1PljFF8l5jFr/87h9/E0SGQCZmHeZ1RSvcOgXJiro8cHFmQn
hwgE1da6Lg4WEhpD3woH2ZOgVgQt0giJz2GkS/iAxyPq0ZI9TLNIQ22eruqEEiy0
ZRdkfL6WFXBXpcRM0IWQa3RhzzrKf0s3Q8WjI6IC7+0tSO3pOZEYmTr+M6MYMrRY
/G+AybzKnC0YUEqup4GBGeWynWTdDpcpQmOsJG89xowhY0NH+esyk9NrCT3CbmRF
sFQAhkcPEORsWdj6mT8CQfROAtTnAPLCepy7E8lo/e/gMoxKgso0V1mfwZf/DpRR
Pk1gXlUmZvnnFhUAr6DWta6E3YtiegS3fWA6Unc0ER8ocf3ZukIa3wrzBkac4xl1
6UiKNaPMrKmH+a9bxEXfqkuz5vWefQ1x/M3J2s8bjmjH/UMh1UeP9UvmQpM89UDu
0SpALJDRu0G3KJSv1t+AHaSyBoCa8raW5lzn9tByvTr83tL1+B4LtidhJ5PUeOH9
Sf0N+HIQfzmooWGNxbDkHs9qhOzd50gP1qjeppNSADX+t82qNV/3oE0GOaSdZiNd
rDMvOE1vohaNt6lJb/MEvaeASBIuBl53rMlKA2nRs0Ni8gasVwerWYLKz55Nqo5o
7QSXHYW6KcFDe+juKXyPXmXbnLLBOya4iWJogKQ5rTyoQq8sVfgyTcd1tD+bBII6
ylmnCr79c4XRUUk2cArg4gGqfSXFt8zGJQwlvhI3muee0ajbhyY/hw3NIA77kiH2
hjhhkPGoOsk+7yUWR/M++l9Ws0VGboopn77B/a4Vy2Man+VB/vrQFpTR56GTW4Wy
xEnUEwxWEcZmZ077alNtTwcUpLVONk/UdT7at2R4FfRe9Pfw9IPR5kQLZ6Qx/ppO
jvKjoXrnCXqNuH0p5tff8qMdchJpqM/H+XDVWxoxKkgLfPIlXipigyWWGZp++5RN
B6D+S3E2mGqiHCnfv18Z/VAgeMImcTj9vkxcuqr3YBWf5We8/bijva647RUsBjIw
C9zYmzBimYQ8P2YXBAo+ly4tF+IKqnbcDNilYYBazZW6LrQ8cjvCieiZ6vfg5aeb
K7YOnIrhvzjWGjYdPUP8nhu0zccdJ7Z3Rmax1GkhpqhH3iRvDGd5F9+EWX+w2R9+
RU0rR144X9vJML1Nr3jzRmTXY6u3O+iXBjxYHKEqgT2yTwjPz6m6F+XN9zsKvrvl
zOrZkLOtgxKpzgvgiqjrX+Z5vGV4qjoX3gNI8Dnw4oY1RcHb1RFuYylpVQ+JaBiY
kgFLNgro8gdm+S3kG4HFsOHPoL789sjwJqHzMrqRCMrWQIc/lJMiWyhzmwLsELuJ
8QOm+OES9UspQR8krlPSmmGmZlBKcczc9Q+sY1W3RikQsmLiVMuQp8OTRnZUmjVA
y+w7f5V5nN2Y/6Jy6vJGFHQ2IVwuAb4iZKNSJIuHGkERr4pHHNyExfG/CwJcXG/7
WqtHwf3pltmlBoZfEU1+isb0qRCSHUXzna7ervghqYGNw3H502ht9+CYGDEX4Rt5
7pqUyUTlI2N/xC4aAP1pLi9PfBL4xGnLSOixnZiTtSPzmEUWoe4h0pbn9cVsJokg
EBIqWD8dk+bHbRYxl5dNlKmdCoJJy2zKQdDi9o/GNsuUdEOSoCBhc+OEfESyPK49
/w6WzBxXd8BTgdu/tjj0i3hYhemDbXuZgvzSFKhwqiE8IbR+Ue5hllfYHpYhecbT
BaYv2rO+3ctdJpU6i5oYaXdYVlLZXFKpNhW7ur71xo6qbesR9sYijqZllvFOJ2s7
FWIFurFTXg6LqkVvALMcSN1DkoiSglBrXFvEka91z9DVSjMgheQ2/mvtxci4gtLJ
miWsf9z+M5g5CfayVS/QaI5qA+X/is25LEWodIgAP1VilXKUjI/r1o/MxREJQLcw
Vv3qhEEodG7VCFOzCRAXnF8rZsoBjr6Kz5J/iN8N5cvPZI9T1Lyz+mp8f9r6R7u8
ZxAvAjW74pVI4bbbs0+TufXmVrR51NAi71DCN7V5MYCRCZKg3ABFDCMMpjey911T
W5wo+oO1eNsgKDCjNtEwSuBovSIr/DfgPLXbZOFJS2MrHPgJWuGZGYYJrHd+UrP9
QDKpavzcIdcUgYcNJQSE2KtBtFkJW6FutjhwKCEwytXNxZ0pMqOQsQ6A8UOtGNmw
C23pqNleIHMX8w3JXq+rjU3QowWFAvF4pkO435tyUKZYRy6ZnYHE0RcVPrlVLvdY
ws6p8PMFzGOgvcNag6RjL5xw5DoqlIPIi8cbXTATqLPCZU3mlc/DMjKGhawvV+B+
+Ir09Wliku/XuH6fHZ8vz0OKymBKUwuGXdKKLRah7PoMb+fjdgAJd7ghuI3J+lyU
5JK94vM0erqyOZSNf2GfUBi9ASk0iVREv1c/WSrTFwcSpIuCTSvGdf9RoNuNf8EX
j8NHlmUVd6954BnH3dhEc5pBMIgV1pPXbJdszSLMAbGiA9rRYqBEQiws5oLh0QNM
Nobq+Nb5hnTVzQwAJkp30LcDPuFkzFyHKB99jF25cN62Hoy1pG6qatbagjPUZ+zj
bmHewL37dthNSRNK2uR1tE774VCb/86ryHCF73QOtMJSSVgIl/5PM23t2fUcZgKP
fhcMzrW3N+ffiGX3WabArB8SzSbEICoqQr+TkkzpH7lRHW64YlVzUb7ngsScfGcY
6qlbngSJQBwSLFS3qV/hK/UO2vqzDD8s3ejbhp4Q4UUwLrd5vxTtF2q8U2AGgHJx
6MTwtOsaK6RezDbz/ohUbqOToxYThND6BpZcuqFvzQQpn61Q0Z3U7i/+fIhtAFUe
E1gUa1iLuw9la6EQoigjT7NSQcY6q7T99owSXY+nUGXLPmrzwWaZsWXU2KKMGId9
sUSwPKBMFe+e3NIUfrFrs6ozQvb1u0U8VSPsXT2iZ4xbx5UI1hdre5gOwfdi7Lvl
OALFD7QzHv6iB5+KB1gu9cET08umIMvXpGqX55BCt02RIFqGtrBikX80eOQ8iesB
0dDPJsz7meIaeumdFfINn5F8qaoGxlvc108YFt9oBi2ImSkYrxu62S1EpFsEjaD+
KLJg8tl9OYRUGcAK6RslBhzt+S3Xhvztf2/e++et9bYWDY7xwZmL3PIlG7IcupMr
Lk5/1w/vDt0z6zA0eIbKuMToaA/OMi7ln8xmNz1FqDEYwLSvHnUmiX7y0aSs32lm
3a053/kzFhIk8hlZKzknd23CGjs6Y+e/8NNhwRHhVzl+te2mJYcyeITr0I79A9AL
aNTIemQVu/oGxqKLr8MhYa1n7/ZB6gQpNxKcb0IAFGEPwPxX27kOQwXBaT/DCTWf
tu7Pyy/hqFQJLeos2r2hL8dVXhu+wT0kcJNpWn8rHSdXscUZCXZeeXTracAlQtdy
L4WqXNO6QaYBSjonQYXthP4Gnyoe4mggoaU16Vp70FPjNwyG9T9ez3nK2Bijixfp
8iJGFw+yVq9KV465VgIBs04yKwec+WthHLRpRD5MmYbji7LkJ6kDf29ghjDWKUcr
o+CONpk3kEFy3T8bYcE3I9jX3oh0x2Wrz4g5D7HtibJyQA6zNF+lPFatLkV+g/wM
nOkGCm564hdQ08diOcJSaI9RbSOxGe5TS1IdURWtyt1Enr6raHwxm3Wi4IWzpKVY
NadsHJgBD6PjJVEE/z3iWmHcr/57rH5F1rVLle8PdtqFCZZuFHO6JAK7BQZRvEXG
1pSYGRPgvGqhPmMVFnbJpyTF7tn9rStxVei6DPnkfbCigqLisnyzSKa2+BsxPecr
Vtg6e6aGfEBp11uscQxt+3De8uAuaL0vl4ThgcVbfqm4DOMulbFFQvMooLsQxQAR
INIa0tQ9uAxYC8QbHcKrxsXT74WjDJjRajnLOY9LiA1bCYAZCz8RfGe82bidgTq3
vXnj7Stlm8LzU5916Z8iA5W9VCNm5/8WHcRbgpYgOkrSTqVl15DSjjMQwIewgFrb
J9LDWLE5gOJcYzm2plDvi2xgvinHz520kZRbnNsoxb5VcTooIYbjDW5+vBICq3NA
vDipa3TzgUmDoeZtAAJLrnkNNIBFoJKGRuw7JLFfl+iPvJ8SJK0CB0BLUuxUDT8c
VpdVgiPgKZqLmPXMdBeZ68otuuPrt5ZOdzxffX2ZTVC4BJ0QFxRpWO1AOxiuTxdk
7IMzIJoyoBuQpZaXwMN9ShbE1suaxxXxYWRzEVDHkV0w0/4e8VmX5O8kH/labA82
Qlcy48VSkJH5bBiRnCjQK8RSLEosJDh9Z2Xt/qnD+Oxs6/taCKmltY+hxS3lhxAg
Yxr1+Bu/FSLWZwBCj4h5id4XWKNRIEv3qT9ePHYkwe3laAnrGOAEKuTHiaHXsXHa
wwAa/SwyVeSTZaTPrBfsFgTYSYW9vNNnSi7FOofXjsjEGNRcrwegnrISoCBD/8b5
v1tEvWB2ELaBc5H7CTQV9IhcILLy02H1O2tkX4SRYz6kurLXT1YeJUkVzXfeE24t
C3/bKAur/82WNo8zBs+/Fgn8ZmLgVsP8xDYphOwjD8Gg/VgQxk+kV4dsmcLO9VyI
GpWiay2fSvLDVI0BL0cDFJEpifsB2L4cvDPfdpwauPYOdyC+DWNcluQwwcSGP39u
O3UFrA2MAOZ7oDSgotFEf4wmny8FbecdrjZkpyRwbX9pUv+sSmIeD84AWi884Ooi
nmQpPIbCwA2UCrqtonBRqUWIUZuAC2KjaYibwBbg2jEGxA4NeJmPVBcMDDhmtwq8
BBPP9IgU7cfp6ZRk6IBtrL+Xl/kEHMx6VKwYy37SAXLwV+MIWiGIUeWYhUbxMLa7
0gIlBXsIJtvfCFPILtuMXBnlzb4d1VD4yOzUgo3EPoIX7C41tWWn6x7WwUjfqVC9
MvZJmsRLU0QW+vXIZOnWXIAQR7GsH9RffLZL7fH3mQ+whkzJHNGkoZtsuy2ypzW6
Y4NrGk5K/aA1LJvkIJ2093IoEwXeSHsiblRFT0A0PSy5buLv95oG9OokoIH1QvAt
mC20XMzBV96NnzmCss7HepKetIsbnPVgfy5kR0aAjnw5NJ81bH26RUUNi4c+RgKl
FLgGlsvwrd2dT3aSgmK2wcu3+9iMVTMUFhGAGfhZNBgR5G9FgZ26oLDL3UNApAaF
rWf4uDKSZ44ZVxfDwrBEmBqI9HA1O2RPJlx4ymmv3hyTxZqv3BNw3RK/4xu+0Exg
CcmqKO9I6dmX1CjStgaLajREXwrUi/PYWSVorDztWzEt/b7Axearb2fMuymNlffp
eE7lXQfVJpca/DJULxJ6ejzZk3Jq0fEiuidgUcnz4EwsGW+M78/oMN7edoRJgYKJ
DQ8DYhZYs0xMG1yDBVsn9ugjKVYKXgmF8HuodqslWXBSkQk/sTGLfgdboZDm+ret
+t356kX2Yruti0uPXEZbDFv8LY6nX+hiTpkjPEhUU3zSHdbhsuk4CxCLlkWsS52+
Sdz6JqgPSD2sTNviHXzc0xZ2M50BIvV5ZfJtauBUBaTCX7wHMLB9esb2C/Wr3TlF
7QOM83TJWx8LL/mkXq5GffdbSIBC1PXraY9LAh+SYnIn0SZTqkwmiNOCTSLCOnhm
wPXvHcTp/No30XQNSr7i27AoPxQfCgi6qH5aqQCNvcaBEG33T99FepoR1DUZX4xl
v02GNpZHp/7mml2EQycyxUP7O48b+zYWk6/JyF23+SWj1RT2K5+uHvYWlNIVjSUK
ONuwR/ESFnMQdfDjX8QZbdRSU3pmNgm3yY8X3jmB4nQX1eSuTRh4fHNB1ZwtCcBK
AkoktRyY0a+keIRJwtFfTd3d0JBzKn0uRWNTIt+EoUbMb63TljMkFGPz5kzcIhfT
pPO/Rsoq2171IjRpj9kvzRdPiFbb6IgvH4hth9aLS+zcpuDcqC4SyVYLubYIk0JP
LBycy/NzHenf6bqngTeTAvFPIj1/kbTgI6JhN5fLRXkZLFYpcC1Y8cswiWXyDgvz
jy2/Gg9iU+GTCTREA883vPBB34U6e7JsNlqARvlJe6nlJkIL2jef8Wc4lJ63Bu70
AFd2+cK+MoSFt2bHAvByj9kX+uEPsjQre9P+Nm30VJXBPEA36U+FP9rQ4YpibEM6
aQtxK+dhRFtDJLcYYZJM0qKZpPATa1iox3wRu7unhwzkEnZ3XFGt+WxpThBCe9kX
MMC4X1Iox71Z015cqn7pe3A1x+WjIg0hCkQhwiTvhtDU8cChhp4vTGjhxTydiuR+
cLDk8LwbDKudn/lx/JpRR5n/Bw8dEQbs9JhFS/R9kEF2CRXRYJFGVBoRjfC3Pvds
AtTSlK1+DWKpWU4/4jFPXV3zonyHi2jTD+4yBSQTV64HSfgMVblzlo4U4v7SnKAo
CcnHRda6zfmQ0874SdDjgLH1q21Ulb+gTx5OaoU895DVqSmoaVKKoBHBKSjbln68
fmswfIqcNhnip/fgFr/HyidF+jDsVAc5Km4rRFLCbz8FC2bLgQQFaurcbYeH2LTw
Ebk1YywyWiVfZDckPTO6cLI46Y8vwnL3c+FyfTtq0yfJbk5F91WkHvNFF0wOOSi7
OEaOuJv4XyHwT6GzLbdt5stwAyDN2f+y+wflXyKZx4qyFYbvKtC9FeCDviOGzXca
Y10BskIcW8x2/+YxVwdOGtf0Bw3tNgz9ma6kTvIqhALqtyY8GW6e4nR9rYVAEhyt
4HJiqzGl85P3PF7wn/4GC+yNh57CsXBOcWRnehAL6SQEW4V/KM8WWDCLdkTb3shK
gTZBEPQAixFLBP+iM5egUn2k0V66KeDw8Ro5MiQDL22+nuIDrpojneVuAk9FBGAl
3q6dgX0araVKPumxz1SDh8kQru/knGIWUqO0opcK+3erB+oqWg0CetlOYYpasjxZ
fyDaLeurdRi9glJ0qvy4Fib2jeMi8rRMdVfru/ArI0kTuHl1+tl9qKM8AcLkGgN+
UeYxXEdsHbkNB/bduFHmsmSA55DN7LnDQNpzE5YjyX10PoYEteu4nn/qYL3dhjxc
5qoGjEAzjkkB58VA3wRo3IYXO8tx+5bpCIAPJyeId/aXJDnWk6ZRdfcZVNXpb0Xu
IFMLPdcZPN84jB16IHs6pxFYjZirR6jAzxS423sjPSx3FJf5dKfSJekFNo+EIeLu
4SmiDCF14DKDAeWniLPanw7VT88DQGzcvZ56i4dTbD1b74mfAofDu/zu35B5Y4VP
yXFylOIqEQ84BfmrFdZmWl2TdCw8u8yorIJw716htWD2J03SP8qdC7Gi4wTdV1Cn
WnrZkT2cg3IcW1R+B3mKqDI7OGtffUhyrrd/TRt4qHZmBwzFvAvXTkQ6EKATSWKn
urU+wj0mRqccqt0kLH7bBf9gQdINqDQ4ijrMq2QiY6DuyS4y85CYkzB/MtqBdoDl
8tyj/tYUNwHMWvvB9WGr3dIvqH1qZtg+eP5KikAu1Yju2bLYGi0oWtjYqHGsfVQE
TjqmuHxJo2YbIhTNpdz1RJ1s4Hg4WJr+10oyE4B3WbZBfbAA79lQ9IwTqjdETc5e
EO1A5bIm02fV5w1CWWfLJyKbJSFhpkUhq3J2ryq2rb/EFhodz0vdC610uSqIcs+7
+mprjSVxYt8m3zHB8CJiukqhN9W2r/4h/hZft7hcAmOBexwvbaRZNUrf11tUoOzY
qiozz9v/sdi99qJQAKIiPn50c05q/4yMUvxfBqKKONeWJzIcxgcfSiLzLSg7F3md
vwHZaRl2fPBwBLVi62RCMP6e/8llirc0fn6lKMl82RVEmrl3IGVLSNhJrGJnw7Wa
7slZmlwIRUAZK5gVEhW5wpxIAF2VhXmsqOfRbo/ibon5EGnQtmuip8goyo7TfO7U
bUNbopkRYXntzbPVo/5VVrt8RK+AYhLVdngN00WGfl6BxARfV13emC0Ox0ngFshx
Ox2WFV+faVIHOv+nfsXZ7h1x6tfkatgxGv7vOBu3nEsYspz6AOIZdw5YpwoLZHwk
XF7ADjU0KgeMc5qP932UEAP0bqhAS9QEF7QtSji6ld2cVU+F1SasJEdbkx6PAW+Q
EOZlzaifzvxEO960qToWFh7HYpYHH5hEoLEQWrpr7csfsENmBsf2LPcEO/FyZwcj
DOY4SmJ3WqQL9bEKfYII2mkE5TRIXXEDg/OpPSn6W5Eb9lnFqn+BLEMfaxh6j7Sy
isgQQ+6cCUJzZpK39waYjcPVGooJkDARSzNmSDdY1zW8FTqo6AnaXhz4eEwbubN9
zq9AOXNvVMgzSHtjbg3fHuxLuOtQCJNe1ABRxSd7Gkv3LZwytMb9+MJQ7qZWaF4G
tqwBBtn8GCqwEVKPEPS8B3cp98ZxXHQpeJ6ryAJtaSQ1p6YyRyeBb6lFUgvGQO7Q
hfBjDkPwUfG93pkK33kok1Knic3O2HC4EZkm/rvYn+Yu1ILqr4q7083/GdzbLnqL
v5/Ny6mjnjxamXURy8Yz3JDg37m5XE8Up2jFj7AeJ7Mq19CTf9SsOjXsMplGV79P
jWxPyMQ9GGZjtjiyYcbNmUMMAQaEEV6UarRFdiFwW9TftICfytsLRutxqHhX8b8T
xWPytd+MmkWqZa/U+YW1jLFBC+xbklk51s5p+EyV9VFkwV0+WFrF/ohelg6U+lOX
nOJtQNveJUaiPgnGP3ipGmXH2LHLY8CNJIU76T8/Cn/E9bIBXrFQUWK+fO6nuMW8
Mr80J/RCB/fQyctm5J0fWJ8ypxDCtiqJmOBdq70jEL9l7eewrONeWPP9gmP6G1Zn
ltT4PCRRkt1zLxWQkwmOaHSXUNYJaHwVx9jDzqi4NUq6ZRo3uXOSt8BfR5Xeksph
dPBMoi3LOabDm4SPfqOGZ3e018LH6qeN5vuCi8HW5yFZ+tMqtGIQrWEtdJb6zIJP
ZgfCaNIAmFAKcSyxZ+qFDGaBwSWNTo3dGyD1CtzZBVdwhpo4qlHfUdGEsFgqMvwB
0IoNixP8Qt6eTeUBh0I5HSkcxZ0m3AQcUOfUfyk4D0CNalbAzqlsvxtDpN3PJlkI
1XWTD4QZDloSeFJrYg54sVBZnI5kegxaZwLhATGodiNCDOWJ0yFD3jA+AfMk9pqr
rmxDOZikszbTo5l/2k4XOkEXy0NT6x+gKNMtqYE1L1YBj/eVVJ4eBsXXHxgx7G+P
mJ83VziPsDDM7uFLZsbXAFesn+pwmSfEfYshBYl9c0oKT1YECZeMX99GDVnHiOiq
mJ8ZSjKlxTGhHrmFI7PSX5yOI6VN5EYHyFAkAfByaPDnKwgfOWAUj12QcFZEzcpO
Mb7waCLk1IHHT8036lwbnx7fXSvdCl5hbp5FkUEOlB8zHaStVc93033B6eomaka2
sbgrM2ZTYwt9vyHQek8SYfSLplikvjiwxYNGo7LrryCb/x3qIy17ep5hsrV/tG4+
XE3royFgTrVOrCU9Qm9FQyA80kunQE3lKktujOQULKu9wtCuPIOCdaiIxaJ83T4W
6BqyA+WjGc2p+d8q5FTCDX3wskckEAB43fhb7NH5r37OxHD36Mth3Ozj+c00y+7K
a0HLm86gzZTi0YDpm+ct44496nJafZEb/9gU3dgFrQ3VOvFzka5DotLMfeUBVev+
qIBs0bB8z+OTmxcWVS1koWPgsBSlL1L6HQMUQd09PJaWvjH8edJAInAQeRIRWZK4
H3A33RGxh6amZCE5+8M1zjuLOQA09d6V7UKB1GL6phrJkIa6GWVCPBVoOlHd+of7
T+JQiTdcyz/+N82gW2cxWFQQ7eLId0+15jbRVzW7KOLHeEGkIWUtljZ72Z72+ZBJ
q3XlHkTdf3vFOXhnsl2Y1pyY//hg+eLiMpI5Nm+gkWuDQIqrtfszsW7dWhaqj5tD
9wU/7bfYR9uSUtuAveuaaKIDnz7+uYuSgwV9DkIRWrgEP588/RX9Ng7vx21Egm90
U8j2qR69f2YM0qyBvDjLtkokf9OPaku2YnYzRhS8G5Dm/rhKMB+Ytwq0DVdeLOEZ
t8ZDDgtSlJKAnoafosP4U/eTJX8+Ae0F16PfCjJRnrUa/LV0sEs0uUELcZKgbP/s
B/fAmv8HZTo01eT68KWuOhZNfbdCPVuTElX2G8bFSCk1RjN03myPtmqM5el5j5Rk
A1vYwdzLirXd0JuHfo9mctPPMlsc1vtoEdJYCEYKsZ2cqiJZPOp02vX6Aj7MUZr7
dlxJ53QHdsSA1bKzSeAgFva3COnxRj7w2Eyp+A7Bn5I/B0Y2QYEBIy4EndmcjDhj
V7qbnaVd1BhIuU+3Z6s9+4nTThIaSZ9NhpLWWTRT6/aD707/kRK8FEZHWhDddYov
LTdG2xu7tdOFOlPbz1gnj9/ew8D+WHs8/x/GZmy3ycqdicfr5oW9by9vyKeV1Gtz
OGCSo1NuemTLOktzPW2dZwtcS5f/eEf4bhdwRkTOtHDfIVvy3Mp3ovm1VIPlKYGB
1V7uXlQl16+3ix+EHiIf1CzTq9AXuBTG3yLoxkvpat5vcipK2YCrOXzSgYr2Sty9
upZvcBSdRYBmfAW2Y6ZZigXfpBBH7AtKOvKrt3NTYHFx4opGrvbBwhk4M0lXIETM
j++jEGg+Pc3lro2leBoh0jzD4L548kXUtScxUSpD5n8z1OWEELIvjcUFXlZgtFUV
OV3eI8fih+YqaAdOrYErqPTlsEihfg+EEPYW9Xd9mwnYlcQCPYfeZ5CfoUN8aqlj
fqNQVbqD9aNid3gKucz+/6h0EyRvZ9JHv5SMfQSvG+uHK7UJSJIe7B/iy9DrSF9i
SARlvsa/vWhUENQRqB7IiO/9Sc9y70d+V8vHqIh0jBE4zuObr7KciPZmc2HgPJ5r
w0Tf8qlpGZTM58Xj2d7IvZEFwvUJZP1V1NVCBLdz43hmxHTxIVmK+6Qsv5mgHGEt
Yldf4TGCeXTzveorOZWs5ZHRTlz9PrYxhVT14ESMUhM5OtdpTH/FQaOhBx4dhTLO
D+Vpc0YZTB/8CE0xybOQeKKAcQ2YRQxv2MtCyUjz1pBSPkPJkYqKbQvoZlTC3oem
nB5FRbuxRiityI02/9daM9llCo0qC7Koboq1Zecvlpg3tNGoc56Daj1IwDY0dHOh
kSfsgHS2/7ExDKnMt3ZMoKWnjTzfo36rC72GKXb3QoPSwxGsCy55wxQ7nnWnLZKo
GiqLePrC1zG5HeeC2MhidF6BxDgoUiNRgZNXXYjoZloUlTgTsO/l/cWpDmiy1W0h
/L+bfesyYM9s2AF4CRbAnpBn3jsc1oJbnbErFnmnhW6ymmdV/j4ks8+eDKeSjii3
z/RKqo4h3Rc4+1sxkX2eTb0yIgi0bUwwkFEItI5qGvuwDskr9XCbLRqQIiLSNxE2
1jiVBvXUaUBFPZXewT9uljkMIuqF9VTY4WwCaxfDmyl8g5c27ttCEBf/RPPslhf7
4hkpw42l4id6C4//2jKOIdHi0i5H4VbA/6p/S8BtgQHyT8f2gMuluzm63EP5MYxQ
9c7talxPQgdJuYpLLMHW4SSHUJkoqRs55PyZL6p9CDpvggh+81M/D+CDXCZfsK1R
G0LlJN5Heg35YK3xWaiNsYl4RJ+Mqg1BxU4BVckcyitCIIvCnnh2P66SGP0MrngL
UCpC6DPUV56xQ+jnHDUo/rYcJY4dW9TO/WbaEDS3gnTv7rMp6OHf46R/IiuTg0W6
Jn6AhKgf0dRWmFgHgLuOraahk7E9jzcRbvmQjLR9wQaqQ1RuPJEO9H+mF0t0OilS
DrBABfWsIX0z3xoU0Clkgu2cF8NCohwIBrsVEXznNbTl8JSXEWbmD+x9XEJUJJY9
F2k317AcQQAmqXFHvZUkpInNHML6KHGEZ6vKXjqnL3H6/q6Q23XrPTFoerx+8zL4
jNlAcV8iO8x+Y7ynTdI2b0q434TfVZAUlS0RctoY/QZEko69+/yIkmQm8uUbSBkm
qWZd6cUpFiPw4tnVhZA6FgDo+vcIawP9wRP9JzGl1y6cYBsllONMBISocrBiC+iv
28tIaSln+oWQyOFAl5oX2FaITkyqMaC555zeDOVpY9FjGM6sIBstrqAafPO8R4IM
G/3G58489VSocN5XzBVaMZyrkZXsMjySRc52yPuro7SIiWR1bWt3vANk4BLPiZC6
18j9Tson5Ir5Pm5liz67O+1zNF0RxHOvDHG3pOSCEoSD0gDAXoxXZBAWShhGQQzZ
7vueJPzFcTOZgDpWbWTxBTAwYnP+9ffJCoP50mAvvj71Mdh27OW0oo1cdJswVTUp
zsLUncX3NZfgez2oIdNCSrVufGYe6GTMN+FGZXDe2kxT3rj3T4wvYFT88VEajMaw
gzD+IeIRdGyAzUMPAfTqNZnJZnTVuSS6KA/v/8I9p02ms5RIKQadn8/znl+lgWAR
3sjvvn103gkywjOwaQ0xzMgqDjak5O0xZpqhzY7Wc+MYBdH8STrQh+HiXt3IlzLv
s6NPdmWlJ4iMWACAhVOMNA42EUPEY2Nl/elzWmGXMpNgRQrFuop0UV2kvv4P8kzA
r1LBVTdPsGEibax2f+PSpyxvRgXswWmdSg4kytc4Ca+u3LlIQvfppWyVhoMbBNP3
YhDdDublZoPO+iEo8FKXSDQwTE0MIznXv/hUBMDbdmdfB9TCMynZ6FJYKIc9a74a
92iclA49trKfKl3d7yvL5zSE8MKxfg75iUsxFrn/zw2sGW5/VOzDwRmMFX3KMZyM
GZIVTRNE95xx3c9tVjS590ePohIaMFKw/Ht2yPHVBAIQa/zihanVhzQZxiEmV3+T
lZa/lEIVURcddz3ieizY7/rMlrXXCKWl0SXizaBfCn/ma1G+ln1+2NdDUj04oiDf
nCILX9F2jeuxWMIg4xZb5QxgIRPqCrdIh0pg9i52RsfX9QsccVlIWY6SxqFf2pZz
r15s6udb7UvoB4d8IkTH/rUhMK575nCnD6gfH52LCAVX1SL9A5CcMY/At9BZaKCo
tTqq+4Jf3nHbKQSDnkHiCM6tAyzTDBn3cwuEuZWpXwAdM+kXHgVp1dxnoIEekHXu
Qh6avS0ju2+Z5WxTliuSmAwK2lD0UoP3FW8aUYcrCQvtVByP/eys3TsSoyg1JMe1
xwrAc98TqApQJ8RQxStjB1Zt3u9zrO77/2N3PKS2SOxJ6IUNgRKqZzLUoJ8eFOrT
d7GQu2LpO+BUDBW75LXq6mtLXLMxnBNlb9TzVNjhU/WeX/E0NIBG6GksbO5ClWFF
/aGV/vKiO9EUZwoHvdQ4kLT/gYVcSzBxHozQ9EXKvJWO5O0UdAE2Kzn6qcgaGMxy
qWbKy1LvEosWMK2759JSrCs7MO2/50M6BVtinVeWtrdfEWPhGrCNV5Ium3C4pGC2
tbHB/JtvnCcmtoVBHKcRx72JoyJ7nlbpEhUdSxP4E3Y1oU1nlX8QvcVzy1Y1p6X2
tJeFr07XEqU/UR49ZtDx/05sxdFXLwhxF8BEX4hRqLuWIZ3RLQ1axgbfV1/YU19u
4jYVL0W3iGN6T1n0oAN8EoWpbv/p36W793yCaK/7pOlAcv8aX0Jo1RcULVmJ9vN5
CHqXtOFY6Y6+Nd8NMtC5AEXgFDs2H58VY+nrZ6yPkTMOPHflTtZOL2S13Vuvqzrb
SKlZeHdT/Hc952ldIC8p4Kn80WvLb2c338O2Gww71RSTC+fQ0pbGuhk/4ixoOwop
FDhmY4xJk4T2CV67tqzz6RQd25+yUlexpQHIdxzO7s9voOnlmdsjwfeG5Q8HDTuz
BZkWWOio0/mC5SceS7ezqWWafYCnpdmys/4UPIq5U+F10aoBq+FQ+dbrLDnEOc4S
oir0CZda1fVW56frw/OD32Nv/R2mx4VNUpAIJnQIdmhB4kvMc0XLonmco7qvI6Ms
mUHqImU/GxOUiEVsr6MbkxBRZr9ithysnwINqiHbvY8h55q58B8WwTxP1QYySW9Z
xcUffvjiAHf+PtLXH9+XUojKYlFyKxf9Rt8QJaDEIQHan5zj4NvlwIGHXCWy5IVx
bBkah3P0/jI2Axgz/FgT7aBDR2kx6fkVGepqeKLofpHHRLiBm5lPFYCMum3Z1iPq
4SppbzGK2bxgzVc86FABCqOGIvyStqPc1/o80Dlh55TsiFnvlFQ2mdTjyyXqgxqL
t3LsxlC8gJxtbwzcPTfjgQkx9exdIFxtYiK8LLehfVoiX/sxy6VOG//DWMlLGiJa
Kwn5N/uOxP0vYFmiyXsha74YbGD0lr0e6XvDECI1hQnnCO+ZWA1FGnhC6wgyE4EP
bN8pe6Bc2O0mwfbqdQ0DHD5b8BSVqEzW3woK5Dw1eH2ZNhDxOMtb/3k8iL0xvZoa
aM7nB3GLkKvxn8Vwd4c+D1teYlQdfK4kB5ZyrXrB7/V5Lqj0cb6WeTw8W12K91O2
FFiQXJL+Tv7phrTaYGydIfWBRTtgfjNstlH0gj11tF3diW2KqH07EddulaT3bhU+
D4Thujrt7JDwplevvJ1mSBTJJHpLOtgxOeo8FsRtV5yX1UizTjOaAr4yiWnpXjlD
NKTXvu63Z9NKtRSXnuvPV0Io5chHR/CyIMTQhpg8OVTHd+DuYfQtAm1eISrwJx7h
uJNMUCcx95ZSp/6abwSZMOBqSIXefWDr1/bHhdMyF6zxkeXKZ4JJjha8g1gSnqtX
D99pVSMmR2bRkh87iiQqDKscs8AN7YhyXOYIdKzKI/8VdkV8JzNPCwG1en0vZRl1
m4KnlRUg6aTrdKI2AdoUXmea/qLnp6NXS7MQ+9GcqI/PknlYIWaZcbeQjJ8aa4mr
MajQQdY//VyJNohUWrFC3/NjrZgjfmSHOQqofdMYNKaKOjSf4+5e9tlI86IeDq1P
WVHRxfLbnJjsAY9bbeZPn8/j3dNfktUPmFJbEwDkZFWhKXXNqxtb33CPQ/p94Bsa
1E1GS1/Wh08AJnkZ9S2H3s1VBk6NqK/ATNOC+4krrXJfHnPnjht8Ar30GvO+9Uwo
K64npbENvp0p3ZnmVWKhTPUwSVn59qCpEueZXvnlvPTYoDinzMVQFcaKoiyGe5Wv
HT4KcT57s+M2cqbwokwsWPR+U0vGye6QWsJV8QangXYt/KYlidHG+YZwvWXOrfZc
0LbaHGBxpRtixcQXBTCHZTodk/tcVrMMXioSQQlyQ3DP7ptgPMPctcB2bXbNpUdj
1zO+g/CVqd+Z48B4Tea7dakUkdIQuhiYJDqK1m0PlFjTrvfTjjcLOGDcM04as2Iz
+NWbcm85RNdFQeEvAKTWrjDfZcvH5ps261MPbhSFuScDWIa2x1PHg/B+s245tRNN
wNp0uKJlBftgJePY+x53Fj6qCXyLz4BfXWz+nTfGYbZMxUTIjsd8xpW3Qd9wCpmX
GASdGXYATO8Y/MQv53nfwu4FWk/OkijwSROnCjJSiGPRrMuKQPHZKoI+7mtA6eFW
Gf9eXd7aXF3QtJYviT9pIfkXQzOE9GVsKHYok5FCng2hkemZDzkPmKAts1cG2N2j
oZvoqN6MYmfahyqn8okgMAmtqV7NEcraMhjMfk32UZ0zS5WnZoKkmItFsC+9qOVi
CZx0qbcosl6x4ip29NRhqkkM411eqiSR4+bsfa8AN4AbICRqWLuhIj+tNaG6+qRY
jCbfBdrA9fngzsIrfhGgqI5ncTAJtaTfCv/2sYf9aZrlrRzx/SoSiaSET4y30FMS
Bqnnxb9VmQQ9LFaUQrhAvlJLTfFLUb1cT7ss+0bRVn+W/9JoqlRCHKdcaGinKAHO
yVL6RF63zjDW+6VUk4zXCihK8zP3KicDIMu/6x42qMRTvQNE+1iWlvQtMVqpUgXJ
EHxBkWPQ1JhH6vpNaJBSRQwgbWpzGWsYiRrQ0uGXABU06JfUsOISi6ZUnAqCKX5z
RX3eG93qIIDLRNT14/Sy96qaUs3E/VXVagHANGk7qzc5La4gaWvcSpSUARt7YWUN
0FbNUFIqQS9eXoWXruNgfHICnZxxbetMQdZ794iiSzgUlWC1kwXq8HyABcRSL1JT
q/KQX3uas1Xw0Hd6DnxdctTf3chW9+QrXuraZyG3Z5N03oirXOmKbaJ5Pgj7kw7y
4kLuf/L/vb52eZw/QKnf39ScBKcEx7HQqnAX3dAt9qzyPTOlz8nWV/2zRGg79oyY
TT+lRF+8fhskK24Bsu7iUBUbmOZ+MiROjnH+RnW7/5OFc1bRMP8tsQImAuvFAxPw
adNHyNAEk4xFLyHzj7K3aAScY/bg82qhZT/1RRdKXdio9a+XstLQFyg0SL467Hah
ZcVm/lStrugCEbn14TDdFctxEomLsljnDyLu0oUjDaojNVOg3DFXGlSjvCGJiu6G
TJ9ezWOZ4NR+frRUfNmCCr81YEGdfY0DjvlAEKHzvVkXYWruvcNhSexyFdof3Q8n
b5jqqYwllP7XNtbkNMfSP218HYTOqZ+vSt/nn/V+2aJ90IkPI2pnSYNFf/cSjncW
2zZ1RHrs/caHleJonsZOmc0ZuHxJHVwcAin/YaYnp6jBNA9NWwL/94kVwT/cnmMq
OamAJyGLVsCKfA3vyw+Fr41Ye5+UVvy4wH4xwUBEuFnX85bW9JSdjSkXBsO9xXf/
1S55IR10SoMIwzLoEZlMwcL8h/ZrQUTEtIykW2t9e6BUsmvHYU7kgqNCr8X6D1Hb
1wV/1FIxKqNjo5lDt2N8s8wqt1FZzIAZsiCL2/yDOeOmmHamVzR8G+st7l5bBdCe
3pJKh8wNJ12ngyjoFViCCrQ29Y4vop7EbQP5jarI8ieU7NwpnX1pWhvWcn4nNbAp
8YXSyBzBDi7KgpxwcmoP+EwwVr5mGAAD49w38OqA8tpRJU5K+iufiKzYkEqcfU3L
1OJOJakUpMh2CcYrX0ZRzN+t/ZZu3qx7u/IIM2CKOTkNQeBDRIE6YEWuE90jOfOV
hL7iYOZMyTFkHYq5Yvfeurce/nxuSjn2kEE9hAe2cUpOefHTB6fOqcdW1ZRBeb/f
4ZKtjlNVUIs+e6Y3eB7PFW4ZOjnzePL1Iee/NcnWnx6zwyGlnrQwivJ5XGmpYIZT
I2ovVgdoje/aydqRVuDOrrPRpegsoQYeDIntT9Kq5QamNH6rwdMI2OYwUTQ3YbvC
K8uIQ+boIZLyS8LdwWazHKdeWOCFGckqM21ASaV3UzTVKzs1anEq/TeNx9z9h83l
Myz9hslzsfLqqco2cGpXFVoY06vru64qS75LAdT66zpj0EY+RvyD6AYeULG2Yu3+
6iKyzQ47cM6f4DFJtick6Atzs6fvQV+y3Zl32g4yDhrnxwZxI2TGEeqsqkA5tWNK
2dAqL5Lhopv5oHrq9whbxszBI3sDFcj97DegHjBPs0jMJjxBcK+p+prtVEXoAwiD
0/TAZamsEO5nHiwKnfIe8hOVYDn2ZtJYv2Zd2EELyiUnHVQyghcVX4IVY5gNQht0
S5V8c5cbM/UErKZIf7rnCOd3UHYbeaaIghhSp9oUnjNcxo779kUDmiltSpgcA+d6
1RF0Rv7UbPX9gyO8jku+J6orOV1/VMFbaRKIEehgrxVwBCJZTO9CIppsidTYDiyz
SziK2y9t9tT94stAgwVEB4cOPY7bxWarZNrCSdOn5hs9eFUDU+c8cpCQlUzNaf3q
in4j2afEIasvPLJXKUY+efzbxOlaEt6ZoxWRxwE+0x9q4cayocllZobsFljonQSB
tNc9CqQV9HBk/r6a8aSYCIkgkD3B2EqBWFSR/iPp0eaY8cb05dF0UsJG/jKDgWwQ
oU7qsiAEoFqgBzgxrrog+SYWyV7+SKE+36espNTIor+AEpgS0bbU/UHUkJdOBF1i
g8WOhbsLnuSY1KLVbw3CT8V7C5ws4PFjojYk2NJQ8oq42hNBHBEicf+pnS6OEFki
5TcExaMBUWkPfBpPqFBU0ClkpWz6Uk+jnETIJwN44KwPhvJmj1p2ywc9LOooMGMA
o1DplFDOn/IAMX50rhosdSga9Cv7qlfRNpOrGIYh6d35ISYdkvE5yf8m9p1jzcPS
z9z0wijHSFki6btlxz52XlTqUQtTeb/DXgIq0rWx07m8jJYfDJ49mdKxJFg5z0ip
QgOrxJnyOoPBxoFJ8GMiNfKhv6YxHKfiSMZqzZNOPPtU5T3EDCzDXCu+W8uffMpb
0kW7mLuOfPQoUsOkC9NXF9LsBzYTbri+nIiIpvmpxCrdYJB5P1LGXNbWHvFgDU4M
tmVLv+3DUQCLzFLwOtc9+JycZwm4+spFyLKuibME17ACzFNoNgytcOinOSuHbOJK
avBpSc3B2pqUl9nU8PXVh0Lvcq2CjQVU8rbZKlMmWxhCNpWK5PYoO3PaIAv+Kzua
7vh4Jt0ZZdDtmU9jXKf45+yDfuagTOY7JZgRsHThfAtqtSfa93ZzoIx6VNyOZc7S
Y2vlijXyvJaO+0PTZWow3K6bcqSwgbBHIHt2CJFIMA4eQbdb0NZbkergFcM0dTBO
sSFhBqQgHUlOGpaE4Zz29W3lzt8mhXSfv7pdBXnev9ksqC64emdVxVHiksJJD4bN
xTumlzM3YL8MnEZXuJgp5rb+XO+mD0Zu5slULOFIabPcxEtGvtrRfWF2mK5Yfcpi
XS2YKKwxZ6eAfk7Gv4cE3pC1VyQl5H8s+BK+oo6TW2flLOdum7wYElhH/XDwHLF6
O/4oum25EZbchyxd3np9Geq/eMt5YeriOKPP7nRXJCc83iUP1qgk74p4fRqljxI3
WMdp3eg4nowAR/2whNvr6v3rU9hjQ5EGoWtyHWruMvBk0jU8fMJwmYJYkANgUis6
rb/FhxYSJ/TCY0T6sIYO6Wn6XEyVHN8OueEBt1vauX3MI3xO/JYc9jTOwnVopbod
hSnjrbJUXj8e+Alz21bsaZrkMpTwIgdlVobA78Zba6G1Fu68PVCDJ0u7HEFIvdmV
Y/OYdM9KzQNzcXoX4lnjysbYrDTA8acOJero565KHGxacC+P71OGVPZHOZS90+t3
fG7SaRc1q7G012hqkSR9dbFVe7/46ahQNGWoVldRzDzRgtBKICELEl1eglo19OqG
jUp/VvcQdF+nSlGgd4OqzyMPc00NUMD2BKsBe0IwWoZIFQAaPxFr1Bz5dbk1AKk1
gdcx3uXGFgwqMHVoIhSztESnutZ266WpWzPH/UHxlJGsDUn6HUq+wQ7NxRdxhGnZ
DzW5+JO+X4Y0lC2Z1Rbj7SEm5m0OA6IgR77tiTShBRlrZkLSAtDsdnVziOP2sKV3
x+JE9OotcdNvN9K1D77jGyLYzY5/YxQRPrh8NEfn7i5mV0P/+4vkQTNvheT9UZ8e
oSqqgvXCGGYHWJjtU/9c244q8lBER679Zz9+fcov7FBHdEUvYsia+YrD05K8vLpR
l3jp62IEBEokOZCS6Yd03Cl5uB96t8XmxzBschB3ONKZMF42vgvxZJq+8uy9ukIO
YYuSDRvcb/FY/+fElbWOo1mO9PWfayrlmlOivw9q5rRXsnOtYPQAXl40nBlc1dT5
eWTOzuggsMHnSDk6HWWX+9C7r9OWdxD/Pb97E6ONte+XOArOqON2zgz+0stVrd/V
OKUFpEaYq7jqMEOmRNPEiv6KQSo6lbUGN/T9Ra9wjbpDi8kZmwBOpCxEjI52vRcT
H7aVs1qssRGkyoyUs3CE4q0ukcmq45jq2b2+YhkpDRcPAN+bHdF3PpDSNTjSwtRP
/jWwlSrU2WCEYkFqoK3Yw2tfCjHiNnKg8hXhtnmVmZZuRqiFI6hgBrwMBkjd90//
/EU4e+4gjDJyBgynHP1OKpCy5qShMcnd2BXhgvB+WMsRxZzh4UQmAetHhCNT6yRU
cNe/zkgpdEiV2c4v1iAOYoZ5YxBSPkmfa7YOoHlWRVeWM3PD0GuQ+gnlFwYSC1Mq
9xUvy/wIULeGx0psUDJFCp8WTYnLIulK2Lswt2oLd+eUodVma+he2FO8MTJTW/GA
DlKoyNpMmX94ysF8O8bWi4orZ401z3CcN4aLBOzNF9v8VGYNyQ+0Fban9+8MfkS5
Nf19z3XLcTyZQ0msdFunHGxlj16pB6jhXE9WzEigyXYVDyJFtram4jxP0ngohsfU
Z1hdaUDbIlHzfA4eHUMjg2oNEERWE34kk/TCEDxb5hHMx20gBsf6CL/0R5Q8CPaH
OKNrGZavXNM+OrCJQiHS9VmTp9fBqvIbCEJTninsP8EqFXpQWinbQEYtIDclzr6n
27Lk2DlKCltGtRElT9B2F7rPiT1SA2ScXec6h88w9rlTeo477/od2iEWY66KZBOe
oZR7ucdPCGX1io/C6YxToL1v6H4BywfExqiVfpyv0blKS5snb4MSBuRTXy9ozRhO
g1zj0jVCnVep4Gxodv5b6zkUfSuYn3KcdOCX05IQsufCQPnSmmxrFcNMk9QXA9uS
geN0l32HInWc9XErZkrcbl+HhEkTQPRw7yNuMxWjobgB1YeyC4DNR9KuIo0VHqso
xFn/11FM9jJLifyb1TkT8mqMgZEI05tEEPIA+7w3zgeh/Q60l9RvM2Ki6Qu1lMrH
7wE0haGEV07GMOXaK/0FDuI9a6CXiHb0I/I6YYy0OFyO175rJlcTsJScpDtCtNM/
Di79xPlySyWRXdX3R90xokP9gpQ6MNI+h5qOxjCNqP4MVfqqIjk8KdJAxHwtDJ0s
7O106jgoyxNfxaZPZH4/GzWdxu3DhXpavMsr4B2jZv25umctzflrJPEDVENNs86m
DE4xJpirLDueTXCumsFe64WVu61+Yv9V7sZ56AFnP+szQBCYqXAtN7tnKOOHfUwy
CPl0fNWWiKfbiDFsbsKHcij+X1DJoUGM1vA/xojCi99LbKtEaxywStJAyDpP1+Dg
BJgYCtn+GMYV7xE8NtK44nnWodVhRGKQggX3ns9Eo+Z9M8os3zQk9RF69Fy3yTfM
jJMkIDPXVE6xLELWD+5F1v267WV/EsUQGcBX3Mfw6Lz/Ts6tbCZVnRV5HEdq/KQy
NtERez7Sr6iKJFRFvI2EUOt4nAwHj0kK7ZjO326Q5aXK4i6NB5EVD3eVmO1xTVUN
oXgqxckb5tG2tko9h15jnW7SWcD2R9x4j0qhxWWsU5ZCZHcqHsWA2mhyxevOnLjh
cM/Hl9R8CSiIiaU+ZSrHEPA/4kr5BY8I+uYf2zcohtFr3hsqQ/aKt5RFdJeZj9tW
K0YVyO1/3aWF9++udOZ1csTylqz3S1fFjxsEZ/JdY5kXgBTGA49oBAXgziL4EX7X
FwGUZikRCj0kJO5UwHABBFjgYq0v6bVUQXtZjr9BbTyVdA5iPUHgh0QGQMU1W5d2
nOGWsBO7JAGjbLqN8vGyoghqNbgOFwqseTFBwKJVIuswvDF8JV7L6K6pKYV+u2+7
ox+67WyltlEE1shfb+JxU2hjfSsyF5/OF55kAQYdgDdCRp8gcJms7vkcuTK2LviI
L9bqwo+rlnczjREKXKuX2SlKYR+QwKTtxqpYfQwjkyJUf733MpwP5YS933Tr6HuQ
ae76AYp4Slzy0sD6UIvgNvaL5+cMhEIddgHS1V5BcR8EcvxubL7oxMorLjUWwqQj
oEvqL4spbv2eWdIYCppcArKMIRUZTVl99mA4+VlQJUFSkWq2dw6M4cf6iD7/FCFw
ktupx0uPd4tF/HRkP3n5Bvkz1vTFbZgXrr3N8H+CB9wY5wDlDZOOGjQUF42xSfLh
3+XQzWmmVtjUuCELQKPK+1uSZDsKyyE7ZqJVU2kl450Vg2V2b1RmmvSQc2aT1qAL
s3cNk+mf6b+nq7zvkANJo+AJURySJcDcN7RO8BrGCLFncIEHddlNebizWTkzLEMN
zX8rVur9JJPvmfS1ODw8+n9nxd7nWPDbj9sb/9fW/pdALR38FAg7rMqfn29cJhRI
ubaM48W8jTtSkuEgmITfPGGH/sGVynZ4ojW0mHUGLS4WicLsRnaHcVpBEGtag9WO
qioEgduLZrTu9BfeZy8pBgbH8JWlaxF00utEfhgdIb/JGtZz/MEiXjhzw8dd6pQx
tk1RTFHF0qkQMXGAnvkce2UxJTrpoPz3R/2Db/cctc0NKZPmY9wMCoN2tz7gQz1t
eGf/Tg7NHs2rJJ6lS/mkiMJK8mKDR2M4mF3sOOlQ2+LjxodrPSaTZvLKbkuyIwRS
AP+Mh99DxI8Um5VxPHi0aGMcm9IQ+nIj32Q/w93Y9D+UED1Z1dbwhHFwjULjos+9
R7iFmpwgwmV+2e1jBFSjCJGZG5w8JDESsZF0XI/uw6Q4arMyzFZrbxhLogauP0Ni
6NCK+wVCKx2XkxobiL5xCaWkOXXBmEwEXbSWO6jZXVsnVh9Bdel+378zrcpGXQNQ
eS+ClGkxNs4gOltotGTTz0BQLzBpuwvEN8BHYyzJHccYsC9rPd7ObBT4BCMOqvL/
Bt8SMfIzjnEAiLcrZIHMhIkOwQsdfPNGVeTYjRLO97Rt10oTh88eiVPPI5ug0MJM
BEVJtMwYqyzKC4UTb7KEw+kaN5nuGBzGcKJbF7u3bIRO6lExhNw6d6IgTpxnPAsN
0xBHw47pqBa9YVPOtQnQJklpwL73YW+jNIiY9rfqDCiErL9nBNCFcWA6ewUZRSh2
6wQdA/I2LhPJz61ZQrmu9pyDPjMqaLg/VHHID5Qx5m/872D9SL8vqOs+s8hBCQ/q
8yvbbNMMvDB2HsnwVBCA0hYMMhSYgeur2lEIXgxFWb2Lt6zCgpk0mT49muGtdxSM
Y+Ta5X5ifQFdMLL06YLI7U+qmGUP0PFty8+xUjdeaIJmVyLTBqAiYWSAbk1Hx6Hz
15RLI++RL8WFtXnbWr0e1lX1ecJ9nnTlXHknbdgfIqWFqGetBEMHJgTzvgCVZl+M
x0dubbyyvGXiGkV/OpBj/sWSTQckJZyOpiKzNFW4m2flT6VwK9gaPkNNSs6D2abt
QS6meIauOdqAVz/2wPUPqUHpivF+lFMjQUY6YJJ37zh9UA5UbUOORgItlcD5Bn98
2vnzpJYH3Wnse4bKdXVKnmVqPIRGS03lgkpTobIZporJ201YiZ929xDuq3N0zo9i
aNmp0kqoutwf7UqgkgEdF9cmmmz01TIB0wgGJT2w3NcjarPAeVRFf3AxzWVPTtXk
mSzSD7C8NkQZd16ri0DpEFBE/PBvaC1v/G4VCUUulyma9DyqqbrPenon6Ev6vzou
WYVMjldQ7rCKejVDUqRU8owDovnwH96wP4h3FxpWkIAYuNWfw+fg35sssjP7pfpc
E2EGEUt90mmp46ExL336Yj3RPU6AhN5yGJfGwGxwDYGs13G2Fx7p6gNyJYFkYb5T
HmFUgjQAMqIpnQnT+MzHvoowgxnY9La2FjUbES/CWkAcD3Ls+fW50d073l2VkqNd
2Q+HLPnWMwzWjyL4sH2BaPlSYIfE1sECNkpaerXUoYYcMCoQWRfH54QEPs12EVaI
xbj7GZ/zv5xKggfY0wxDqQPAyfnlirClqy9472k/q+G5Dlt5Hx/bOO5RUfIyck9X
BEg5TXd/m7BaZ4nGsoLJg55KYNXb+96L/hjT7XWtY/2sHf1bzygkRaoJtnqOD4KH
LKxW3GOPYguMUKMQ39kx5o/vZD9ymcYkC4OoZ4prC5HG/ME2wilDVKu3M6On2aQo
MXNQEOKI5Mk9gPRxCgoA8H/2EP8S4f7alqnKd1Dote/e9Jbvit+Jgq9cttm0Sp+t
WoEeaBJQOtRtkBjPwsBDcghbXvMPp/c8v7Poh4v6FF52m9SdxK7ohK5toK8B3hnF
HGckw/1k+t2LrCyJEqJs62WOjPZ1JV6MMLDD1V4lgkWEEkRy9E6TouNrHWRWhRjw
FO6B0OQk01Ak0/NJlv8A8uQqDLWgUkD+no30mWMQGQhsp+q+t5IFWQzEWsIqvhNQ
/aqMnptmeoJKA3t5+wseCSQxI8RSJHXNHjT83jhVMpbkuk8G/yHKgUQK6tMEhVp0
khW29mam/wlRronaLUdm+4ocgJRL2RBdKDVRIY6KGPi34AGBwoJ3jZBmMeIAHdKb
5yWz9FHKlpRTLHeP9z7IWIMxTuFFhQ452G/Kid743taRe5otVh0yUvDUoTlcXKGL
PC8ip95tmdKSH3LW4L6aDlzqTAemX08Vyix8VavRJMnUFEJqHv7sarX/2nrMjatC
HsT8+Taok6kiVOwwGMT7ejiu5l9EaPrCxBhh6Uu9OBkXpRTNn1eYaNd7HidAHBXs
Oqnnc3dqhbDZ8JQa0uOIqzG/ZKanpY+MZKoFV+GNMMosXhG+unfCjvjJKWvLhNpz
GQrIFnG7nhdq9u38lHaX52rnwTVTUiUEa7ZdTQGxSZewiAobbxOvL2pUB6UbcuHu
sSHpyDATCDfEDQvSlT7xJNZ+SUzQ8OXE5t7O/ApU1X0WkWPp0hBOUTlMgoC4pZty
I0y0n+jz8yNX3QcCV9WGmNdAKopNUz76rhxIMPCuteP8ILE6KDXH5wjxjLXoHgrP
Bgle9Y69GUMvt3d9cYbkW2Zp+5bKYl9E3aIfFbpkq7tP+5sG1b0TbgExdkEGn25k
HvalcIEcxHVpoDvU57/Cn4dvRA8ibdoWCjCckVKI8mVX9fIjVLx31D+Rlb4KWCqp
ESzf/r9nWAUvJsNt7RouNIxWT8gFoERwlhDqMpTuIsJzu6KM/Q5kaWc2z+TJoEvQ
Lzn6ObJe2Y3UgK4PmVgHmVsy0Y140bth+0KhFW9F0+rKNR5VQvn2oAyIgYSki1Re
mXR2t633bFbQ+bsalhMFY12XKo9abH1jiAsG8FdKRPAA251+6Seuypqtnvy7MuvB
laCnVmdNQwjgcF60z7y7KwX5feBdsErW2uUjYlehXtNPoj3yIqlwSK88MsSe21V4
FkUVehmgZMK8LxAN7xF9KIcQ0bKRPWUpspDtpMRQ2Tp+voZtQ1kamNb7fzDEsYFn
4f59xfNb2j6enHaZGlFAHUaTWFSI7Ssr5sgaN4rlBRTeGMCUNjFe4oowHt2YBT94
/S7/CNU2DbQJasxDzU2qXq3PJBs7jr2tnsYHzwverVTKUysSc+7ngph4OPqSZEZF
3aQVff51GxDOzNEB9HewU8PFnsEwWB7h16rZdbExRHiuptnwLCsziIsektB+SSrR
VvizV582ELM5GHMNfy4cnSuD6jt9xmDwAmUwQ76J0mby2tt9qb573d/eIYl57AYN
PkIGQkmJKPyfbMiBe4Iuzczq0hrbLsH9byWqQQJLmmWadeoalrmYE3Wo50EtDXml
8gy4L6v9xDm1Nj1e8QldyixeiuDe7eILlWcDZp4xkCm0bDOVV/nrni653XrPrSS3
MIFMWYnDPTbESqKRmRW0ZFeHn6Q+eVuPSod5ZgFos4A/0U2KTw/YW2EgkItLCwGh
TDNGxtQvUgWP0yfLTIydGp9rRK3J3OyKxdvl53QQY1zSX0YnofxiJArAa8+T1Dea
nn80AMa28yjfs44ddIBRWhFYiAagzZz01CaWrGEjQyO/82TDc1UgqpVtqD76hdF0
1C8DwV0kHpCXHMskofE9L9OGimUjUfcgdFqrExNOE6fYs8QvTM2RUpLb1+jlUjxN
Y1O+23A9tzXanS+RbPzTLugSmmbi2+AdFQbaH9IIujEgYiXjMFiezKWRSJEbqZaD
lWAcZ90uQk/AIONDDUR9uiM6QUxEkwlCAIFDv0/86jXA258wF3Sr7Bmo3KEOBdRC
0VQL2VtGNCboCdo5cGa3U3U7aQ5MiqbJ+qwf7LDvwCnF39XTbEdYnb3Zlu78RjlU
9TqrBvFxaqKPo2GyruiT7wd2tIGvvIsFMaf0D11G1kcIJ6veelHqbpO4ERKZDSMp
Zq3qQuBHtOxqaasaVxtR+ZTxDuTZaw+bYCiDSaApyhiiJUjol9daBHTA0CzDGIwh
0pa4rc4c8IUtVn9VCLlBX6pW3Xwsxn08G3BlvYOWkDLguFA7apzVq+HJ3eJclYi4
hqfk5n9/oEtp68OmHM+oCyxu8HrxwSjtIro0e13dVe1zgsForByIBzOPvaQq+8KA
2BsVz7nsYAQVWG1oJyV7BJldOqRoL3laykzvl/SOofHCdJrm3OUs9SJOFFdgIQul
tmWakqYRVGGy9BZyvRgRQqHAiNiXY5SM3/IwJx8E6y4D88I5T70zy0shYPdodu1n
3kOyCfDB+TbZmpxXBHS1qKlcs9i60wDA+YgV+CBnSvfwvc4WVjLPr+CN7M9fCqQO
TyRc7LqXAKyf65oiIOAeg/fohqh4YYgAFUqWQI+Rl3ZlbZ9BRzZgcDex3FPsUc0L
cj52Qy33Kjq/1byCJ7ddo61K6kqFvIKl6MaSHJ4LrT6ErDbA19d0EFhIJxibZU5r
+m71m0BbEn4Q1YyIoRb/SnFweYoeOcNkD1sfRKXmCpTer1O9BWx+4jUINBTrwONT
5r5V4Wm5wJZmc0Ybh75pikk4dSmG9AzRMAlFe7pLaJSE44QC7SDNx1Wx7WBKETQp
ODy4wANCeLolQGwECA2QHaVVNpVR3JdGmsURrtyF4kmWRIJOFylBNCp5snF9cJyD
8CYTaDwoz9Zd6edtIU1cFDURkpChnOLJ32dbYvk9MHSHj8rQTsGac93WLObmZ1f6
M0aa736iCM/zOXONM/8pN4DnprhVrD190opWb5FjQOKtGdDFrejDw9xNGeJHkvsg
3kg8HHrTN+EmH1lRjqbgtj1e4oDBw3+jFqFYNI25w07zobtncW/vbNYgrRU4OmxL
SS5qAe3eKdTN2ZjL1a/9Ypvu5qajNafYsNJrt+PTvmkS1IrDwUBzDb3Z7ANWTT7K
ll+YTq0O2TKnKbCVbGAagS9kUkATflo6/9OCzHHjFPvaX/k4BCrXbs9MttCFLB5T
M4H9odax5mlRJdRS7xGOVDuWyaJp6MTWL/F4qC8tz6FQJNbIrUzcqLOy1Dm8dvNW
XSXX+vt0ZTKA9YSVzTnu/kJDUgP0sxmXikUon30usgoIdyfiGdmmmasRi/07yuii
HhXfZPK9EYAPjLJzZEe9fPcIID3t3QBROv1qZGIEFH9o8KQAolKloRj+Mhq7WD3Q
PIHRTnv3oQk2eOBSBHJbChjxZkvAVUVrGTs0N/IGSgRRq8mYY1r1085iTGp27Rcl
/vIt1aGzZ6Xs8GhCbJupTXM2YeWRb3qffl1MynNXCmR2QLa/LAwhw+cNKQz0oRTQ
S2zIa1UHVjx2s+uRXuFLQlUvV/ioiaLD7OYoi9knp6+b4fvh30KtJ570lVdYCCfv
dbBYAKLGqabX/GTDBCpitNlvQzoE9m4kX4R+B8P7YxS8233iQwdH9J4SZAP5TT97
YsK9Prh6Gc3iEBHN/KTrrxr5hZF923HokUw6PBxixYrDl0TluYdhwDVCNdrfyP9Y
mlyrxBo+bEn/eADxer9c9bEboUQziCF3df8VxUTUzNzcRqq2vp0aLIm9ps4V/tj6
sqUGmYlC/G6J+/HpSPJz7uvH93IqJEhkcKwuBfkKKqoo9tsfwbGc+xvsBqpfCwIq
S8/GROssVSvBt3uenyMTWjtyXPnyHxu8wiDUPmTzYOd/B7jX2VnAqYpltQMe/mCN
GBYJWAOm2mo8qg3Og52XX/Ebjdk6io0fD5d6R1HJfeeT0rakp6tBClhC5bU2R062
DK56Lj7IzvbiPeAZZm9wZOSMyTKlzWhRRPnSqGKx7Woer/i3pQ8OlBOOZQIWZv1b
6rO+XD1mpVWzrIBTl9O1g6L6M5HRptGAyqpod2JowT6BXyk/NGyKqRc9Tjl5pwRx
hjUKXAjVe3dzz36YHZ3D2TuMczA4fMsGIw4ynGJVhwncendpoZ4EX4gBKsUpj9ax
i7HnMateZTQe0cvvyPW1nHJcjCZ3rgnPiDLWEiES948EhxUbF/LutBJAJXSkPdb6
tgmgAskTqwy/bVmfL3U+3DNsw0c74ivxn1bBU/mqgwnRuBZL7rmW8HXy54JEW1fm
kOHcxCxotFaxEp2wgxpfekqTyIJI+03xVx8qs5jHyUXn1f6wHauB1yG8PSYU6WZu
xTO+CXLT5Hxd0EhcpHM2cTuFCBWu3BBmj01hClTUml+IAQ+03IY7PSso3GYZIf4D
jBGUuuv2tmTFQPufCwHy0Wx4LLbkwkSbZF6dWwEe9PMvB3L3IWUK5CoqQDqoX8zh
6lZALsuaPVa9TsmwyKTgBxmGmqVO/eAKBSCd7gYkJASSU3nSU/7hRXvjejkLFySc
hVRKC2ydtBsLNO1IjHzlSpkH8j/i5x9MnTPsE6jr1oFGrwNaQSS/o8eSIgZcemrd
eJctajjIz0ivPR8laTOE1XT13bjWso15Vt1699hhroUlgPyBEV3/0jIZHwMna0Fa
q3j6o7JxVMzJr4WDtCi82245s0qrrgR0jXFH8FSczXpAcmgTa0fkEJQJpQ/wINGA
J/Nm36JTaMNHc9kgMH2HJ1s5Ix61O37FLiJl/g3dSZdAsvXQRQi57UG7E3IYuv2z
9d4oo6POpvv0758FzL8Rfc6qcThM8pYGz0Q4wBeHDPIZEicr+ObnXFvwwnsqY6un
QtReGRgwpmMKP2ipCXd0hKd0jEceyzAFdCRzxjbETYWTiBt8ykwF6T7jIQI9kL+1
T2UAjX+Kns3bTCtGCo3ATcqccbgQCDrPuHXL95pbehvM+6xd3zxCfiqgqDLbbOQ8
tbEb0SIPkPdJwLN84YnNmgGQ5kwgY8ZmHBoP3raClqKrvEqcq03FC2lIsHbmUu7Y
zHPDX14NEtFd+dhjZpGMx2FBDHWUtoE9DxkzbVPOkKV0NX3XtgIaRXxSyFjQwz1Q
arDc1bqlukYsQ/KgTftw/iDgRfLvIFs1HsF+9yB0jYAVAGUzVEIlvGj3wuLhgZ7G
u0s2Fk/TQobRvInSolYQsnZ1zoc+41CIj3DdwSiYK6/wTeZ442p77wzMl4+g0EFZ
9SRbUx1BLnDbHZy7DjFKFbpFpqyM0ShuI/hbF1+yH+Bgv3QEVARMzpE83knwdoW/
+U5i9AETAoRUlUP6cHYZyrwIwEuYg2BwJ4cIwmY0e7eqeZr1Lu7nZ6SiT7no6HjG
/WK7dlbnfIztZZg2cd1OpxxWaTlRUOUmNn/w2J4gVFn0tWnwyz+W0gn4w3QBPKse
MzelLjLjmUhNn+p/g1iOC+2XR1zThPKcWkcOBmClex1d0DrFFavIu+pYRn052Qvc
XwinJTKL0zVvRp06XuyK8Nu/baZ2MjKDW4+YwRH3nM1fcjstAok8YikJG25JXNua
FnxCwXt4q7vTa/89MQhCuGXUPVjETIA/Trcaywo4sJ24N+7G5BqnE0UlNoNL4/ma
y05lgiW6Ghu1hmCXm/KJIa4Zyg0qYGkHsarrn+wb0luggG2UBioC7hFZoyjhQMAM
HaLfiAMvgr2VnYL3jg6b5f/5Aq0UX2H5lKORC2ZXKXNyoxCXsgDLZ9cISUXYvg08
M1FMkuX0MQb1awdsweQPc0WdQZ7aXrqyI3ZOZGnchMYU/RRmmypQaItmOO/MqtWT
cZJOee7kdXw3QxL2Ns0KZOrrW9cx8MQYKOsjctyT2dMAS6RXq7rJmZN6f0lmcsJ8
R/Ag6cnEHWm5FxkBmEQk+AJ68V8VapPhVSZQtXQPVm26J8gvwHD31rUno+pqDZQY
xKwRH8C0/HzQKunAwUjaFY9H/RKXSy+h4gkvzBX8IngprlXeapvzdVwyADJlWATv
1Tr7Gmb82kIc+ZiL+njfmcPVz5V8DJc1JHXN/+hkPfax0OZMPYu3KNbWa+/GrIVu
880i1LbVA0UrWPt5xyFc5/aPmKQ80gmmu9opw3Uo5YIy8atroC16kaBeDRhrt9Gx
t0KQ/X1laf4u6935eCKcvJePWhZFBREjZ7k8qv3g+V6KRlyRY2As7z/pLekWUfVM
ev4couK5F59yY8BbO6pvFxa5q26/TPVVXvEmjfR2RZX27vUNgphLiISm32GJ6s/7
J1HwTGeQ0GvH6dZKOsqh5c6l9t6KU/mDXQk7p15ckP1qF87JcnzuAKWe9CBoULpw
95+Spft3d+xffgD8kBA6Hjz/6HJNNojtaViLJ7ZIBta/oxMf+ss+YnEs2fEyU0lG
s2lrD4aA4/oaYL4phpoCu2r1rX0a3nmn77oj+rmRiDlYFAgoQcSzASe4+JXYBy35
se+IL3Yl1AFcZl6Uvag/UF+Q8yGJ8/9syOOjbRj7vOx07onjZW/C5xUs7vpjfikv
HQ7ROnmk2wxBtJ12iPjE+avZMGYq54gFKFs8pH3pxJ7syDlLykwgjSRJWksakNbe
bFBRikhtZzP+mxgqHeJ7G8NhR41GQCCL3OA5cisNjBs5PyQiTDMD7EitIzhZhOc3
0GpxB2ltRB7oYr8Mpk0ve7AueQO7WB0L27Tju4dHQR2DejLMSpjd0OXAVRaXxHr0
A0jjJcnfgDlwObI2DfEUjPqtkb4KQGWZMcBKQoz3u8l8ZYh1XMQSFUKtl0nBaLI6
HUWjRnfrc0BhTJK5QD1jMc1CO5T9yrXDsATGfuwyK3zujtkYMt75aCMnhegAbZaH
7gYmBdp5dOmDOJe3lvcS9icufp8C+ZmkVBAIY4dXTm6vao7OtS3dwOBZ1BTyNQqD
KuNq2Kf4JNNcJG6U8H4AxtSv1Kb5J4az2khKFh++/XV1yACFmRhjqfQU4C81nc1/
llBNSjwAvlZ2VAS5ez/GKaIwjiz3wCkjA6IOT8SAH6SxpbwubDHYoZ10ipRVCeA+
sM3DzpjUQwRji+T1GFsNoB1VjfIIw+qU5Yu6kBGu/4C0Yg3l0NadfdJJU2P8El/L
3/tESJBv+bu/tXZo5Hb1etGl7H1SEDmEVlNOyQe9B9+PfLi12BR9KvVlEngqCNCY
KUgQuk3vTOBhNbaQ8GqcK65K0PFOV8OEcmTJ8yCiiTLk27HmxUGvXsCVPIyDBglZ
UUgTfx6jc/VF91uNXDGRALt9Z2eAZSyMqsGEfcOYviBnh1rRNINcsdQTcBT9evpn
h/qDq9/yHV6rhwA2nDMSZyXf38M/y1HYWwFq528iTJaiLSsFvtiTz3sJHlzgYSu5
tkZcZPUgl2Km7O8W4fmbC7gnxXHhdROBr0sE21V3XTK1zCYMFrx7XfZYzEgHbAQB
MdKTy+be4eHVtIXd6CCbTyyxBrjqn/Tjx3YFQ2b6ASz49geqSMu8PhqlLP2BItZL
ZdB5xJyZHRD3HU6i1/WeVVT0gnWuDa7QmiPwUmVukSX77NZgjPvLRK2DONrbaNVX
fOeh5mC5RT8NgebEInqySWlqC9ZgffZlexGdeeG0dUzDY91xSMoPkXB/yqeG5pPY
jf25oxNznowUd9WkAp7p0WoLjjyjcqvno+12ztEHeXvHrdivU0bQ/gDkhbEZYmaj
zyWwxpzNE2mdE1ystpoD6FMtBsVmn1dzekOyG7W8bHQgcBq9i0ZM5J/K/+Tw2ulY
ThJyOqWYqLHjYyep/feF166FTnLQFuQN1+ylpU2+hr+EggdwGuuWp0i3EpwFDbJM
HJznbdYoGQjKBDtaORcnam7JcBPid7DmmSQFaN1bpaLbTUQoebz2DO95yWogaszC
aiwSBznBDucwgUEBHTDe0OwQqAs8HLdUpTRI1bETr4yd+uT8LblolJXlW+QExWYC
WsaUhG+sH4FoIzNUzXiR2SuuMzkILIYSriM+BLbOInrns6HIv7qV3mKpiqTv8B0w
UIm0V4a9a0Qd+HMm06eTKhXOdKU+hRsy/SZU/O752tC7UMhcJuhKBjELwqhWDWx1
lvN4X55r+9++3b+bWdDAK5WaPuOjDiece++RezIFgrnDPhOVqXitbNLxtrHhBjFO
f66IU1ho0qPqifOQMxVyug7iLUlRZptPcYj7bGzHHiDNB79GO4V54YbU3BgaPq68
bLQRDZ8lb1l9UmfMe5hRoJ1eUmwU6HPaKwiPxoJblBEcxVqE0jlyVQ/0NfRdSDii
1Js5yXKBc0NZ6e2/23DAg9HawZ+ucO8+GPM69zT6upoAREN/gU2EatI/i/TtGj+c
riZoDVoVPeb2LzlCaMFZin/ufq24/MTpM4w8ypy7bOG9cExkJVdVyqTRcohqXWkw
xDtM99sVmf9pfDTWSANiVXh3xuwjacec+ddjHhH34NA7//z833MW6gDrVyWOUk5P
9990QESQlG6hLDT9r8unYNdMcILR+jsDllZ5RmWIDsDOW2GrY9gysNhSQb7IQL0k
CcYJyaN4j+1mWAHEpmcNfdzmEMz6c1cyxU3FPVX71T6T7+Px5gtK+qT61q99ktUb
qZl/STslTrBXEqzKymsIte7S0+2VIgPXHrc3nSkqmBSJNU9LJyqDtkWma2Nb/wOz
3rmxQs4maEpv/DcO/a7gUQNe6sid20DNrbwIBjvEcZEDh6zvl8xWbeXgrptx9Xud
U2XtAsnthFeui69ahVyqaTuZG6veitzgX/wydF3dVhDiF3BMG+OMH9zLHPP0u0Ce
VgQmjufduyH/qx32HOv85QInwFYhYQ1dwO19TxUFXPmmB4JAVC0rjdA3A61TiKkM
x410qjbFoxHzP8emvsTqwgMURG4W6At3FiIrdJbaNl3/8v7Ve47Rz5S3TjHgOSrZ
3QRMxJjax9/qw5MQ1ON9f8+akWP390aeqWgaUhiYD0aDpBTG3j6yomA/S+L0AQxd
TN5MUhTHECkfgdYZkxBVL72ZB8g40Jlpb+98rN7VCxB1kXu+IDQcqiWXanuiA5c4
0P8thLF4HrRq+gqxKa5UML2KOz2odIhxr7KmuxtsBJpmODoNuOnYcs/nrrvjsnB8
Ax9/wUSZOwemWnBLHNIM6vKiqH8JZY+c4Qcj7A8+5+m6if8YPxmiN9BOSxlUcSB+
e/QTAhuL0rA1ZeWkRoo/wR+kxz1epLpua5FqZO9w3qFcE5FQ46eyDH+jpMTlRumT
AmN+iPyF63FZu46QQos5bnG7vFeFg1oAhgANWOoTeZ3/eZlGQmwerdq30UfI6gdm
c71IoSgVSXmiOAoGsSXKIiaDxXx05bntPiq34a9fDCHbg6QLbPz8lBvUkb5hh7bE
pHlKyjJckgyMcyECrGOWeZLjPCJoMd9rIOJZqfZbFknkohc8/KAfvsNSSI3pDLak
O7ddxPDT3JRfTBcgbf1t0ht+Vd6FqGnO6zLjzVMW50M58Am8kbgGAbcAVWDU6y3g
eYMlI6I2cGarJ4rOphL/NDBfiNr+8+8ffDtJ/Axn4+2HPCxYtQdkfLqlRCOeJNrS
Xiq3GKYmKpqneFkJ2yVKlVKys+hYPAU/VtgpbMc5aO/OSZ4AYnpoIMHXoZ3C/86O
KRxTPoW//JT+ARch19mxaoKhxsN7ZZHPhIRfkcxmSbsP6avKi3w4YBZOHsJB/m/U
XwNRN+IMFZuEbGlL4EjUIpZOVWI+zZjQO7jp92XYL3iS4PLb3ZerEq/c2+yzsLNS
rADjlHywkC/dQoRSDNce2CHEbHO5xUHUFrE3t2Waujep55inrupgPU/qhE30TsKw
9bVmfY7Z08ZABM2q99Aer2hrLOLOHcVvA04Qo4nnKb5P4gY/c9S4yoWMNSy686cX
LWTPreaFTy7pkL8svEmgGiiDp5t5J5SoGITbPIZfXR8aXGDg9RaJvHNZ1eNSISlC
Cg9V1zQfgM6t05KlpuyVVgC8yw5nuRBlwvcORUoHyXgk5akn2RmI/mrrMNBdq1Oe
k2BmGhDRen1X3iuRToAk/Ygqfsrd12a4WSCMSGBPS0r4IknUy2Qm5igqFivIpojU
Xriv6XmRvY3MDlR8cDqFMwNn6vB0rMdeExggsrpkExzjlcdZoBnmTvASXeSOEngq
JQyIb/vYgd6xTe4i7Mkck+5PS2M9BY1D5sjhgjGqe389IJpWjIaU69RD7xec+Xqo
gn79NCQ/UJpwW5O3EpEw+A7saFxGLIJ8giTTmO9UthSs88eHBUpjEa0lauBSGXGj
BlLK7Od5hR6KN9qxAuvzJ4R2xicek/IgzgMbpw+yfWIx5SkzE8/NyUdM/j9zzixG
J7quTFwzqy94l37jRfIDMl1fr2IVSutzWB9qDgRlxoToG2U6wSrRzi8zI4vb7+hJ
ALlNFR2WvQh9w8qYooVWzb2RGZ3H0soAJK4QSSqglP9+ogqUcfEr5QgqXontPwnU
9CZmJFBqdlRD9djgMKbXYxqNqLYAftdxkij5T5vAI6+mRF7CXk6vCt5glpgkT1eK
EMNTjopYTF4rkz0mFw+Hha6wQmqi8cjQYVs67LQCm9/Vq+JzL9tm0nqvzINU3pG4
T69ycboV935ySvv6K74bRpdoXVDbXSCXugEXUoQYkDOJUAzGw5TeepeXKuoXDs7R
h3rjLUeiwUeXU086bXRD58N7mxO6Hx1znfUTIUO7HzK/YMhHADpPrLOCWTgE33JG
8SXYh/xsoVnLxtH4GDARuZFnxAX5ygmLmKpjxTbCTiffDCY6JhiKmPRo5GfOpLTT
f0M5cu26ZqYJFS4COhQ9W7QpEb9QfsYmdBvyR0kRXJiptbY+jGL1Fg0oDBOCdQbE
NK8CbD22bg7HLy+q0KsgsY2/U5fY2E2LGv8BqK+mBNz6oke55ssbyeU5Ow3b5zfj
RvViKcgv5MFf08mTGdyr09Yr2M0z7ChRiRhFGl3vWLQi4nLZ58r0VMld3dYjvVMG
mdj5Bk02dys5IlzjyH6a5rjHgvP/3af80lJQRDSclirlJweiays9jbkClJMM0vVs
ah+iy4BQyC2A3khQGHscKMnmjW9tq7udV04mRfINJCzJfRmk8VnSTxYOlqubj228
MdcNonoC8nUYHCKTv/g689C9FsiBWCFL8EEqkdlzsDDjjq2q6z2/x1fvkH9Bfoxy
pFVPG0RO2uYoHF+YuOtmyqflhloXxcj9eYqHFEHt2nnu75aV6QqgUrn8gDp8crSi
i3XIOdzc5N56JYo7WtuPLlqP9nOT+ROg4k2Zc8mqh7luf1a0ICZh/TXC8Krj2fyh
lrC3OwqSMsvMa3JngqEg9VQRjsNIbYQst7O0VCO0V66HaAjh2HsbQpbnUk7F5Yds
jABeRtYgnlB4fnfT4Fiq7wbie80V1UvU2lORzpAcAluTmOAEyuK82HVugYMajbN4
m+t6Gi67v4TcTzuoddSdQHEnCkHEbucf6octZvuH2RMQxNNIcJkgShxIElqwYJk8
YY4HyXHeZcmzls4SksqXj6CGBBe6poswARz592M6s0mZ1OIRvNKz/wje31FQfs/i
B6000HeO2QLMVriVk3Rdm16szITQyQxFO+76i99UlNoaR7I8gW5t7ECq6fDcbKXx
lQMIuTKVC3tG32nMt0ea32iLmnqkLQQ8SBwCr0B3WhGc9MOGwnoJMc4wMGoTgQoQ
WFeaRJEkSbGINAytGCoFzwYi1lMgGiC/FXyhj3J7eDvPb8Jron544V700XiA6bE9
DZaEjaylkXQJNmZryCkRxUVqY+IfTrkB5gitqPc6Fi9RvqX7NfF9BTTvfQyk+FVA
4SUBHfxV/1jcjs+17hfxRQAft0ZITMfGGAMv17rfsv8XydtK3WILUHKpNnhoK9jO
UbRvVxQoX+it2XX8VbM8JkiMhpqtwyHpre3CyFVW3YzDPT9LAdG/XBZ3/n62KnMk
g5sOcqzaj3vsU/N/V0jWbnlmE+vHF5/hYW9kjHYQVYG3uDgS5jhN0N3M+4s8mExh
JKBWBfDO9qjT5R0o8s50UyNL/ckVBDiuLGJ5zqbW7Kftwgqu+CHQYznLosUfzyuD
lcWDIABe+idwneYfDlCWeTA0IBHSXtaymk7pDK2CcWzbloAa6oHOfETOhyFWQVmi
y86CHyi1To2hNgtCvt9SE094A6duP1fpPnC4ajzVbVcTcp9IJKvw0Mi4lhGNO8Xm
e023tMfcd1rYPp9Wb5lis1ubeFCs4iLiSW4yxGM7K42FAErUgw3F3yWZBlWSDkmc
BTIX2nLTW6/Hwqqo58i4BibTFEI6ugN0We9dc5h7/GkHI4FiC1ySrw/koL4clWgT
PJfkehOdEM8KubgTN8Khsfu2HwcK0M9b6tsdp6/Mxw5UAION6WrsMrymJib0rWR8
k1NXBEyDP7RuoNK8ds/31unorE1+YGiYgEqKSVzBgL7oxvIwWfDBkg9lofR72Z6r
59MUpts2Xii4+tlAb3/VctwyAsa1CsUX6jy67vGWbtE0gwQZMq1ZtNJbmVsih5LR
ZjImvNXHyT/tf2l1BBCWW9/u+e1McQl2fbSPO6CSr0PwJ+w/z3Hb56sfh3VPZKY+
W7kjg0DR/A99DH9uGLjrQQKJW6vQkPSehu3Lbery5gR4fPqUQ/YKznwyMRkKHt0Z
fhgFROHe9Hr8flB4VdG3uEYrQ2VdWr+ic5hFNW2deYkiuTkwAG6FTGu9GdiQjaBP
YzZLCVDO/Mcf2cNiKRvzYuml41djiWVVgPZhoUrq6VNqqdltiKhVwkhiuGCMvktl
Eu6CTD/c2AbbilF3WawlwKrTPjuqzjI9jhOdPFJewjgSSKD2ZgjKYLXAxK3OhG5e
yesV2sgYnbNM2fviQbjjFs4YVGwnoL7+U8lczXKwWHpw6XbmcyL/QS5F/JJAq2yt
MyhckUzFHn8NnBukclDGSwJRfHxiWWferUVq1a6tdZ+d8qWBYV+qJkysOfrM7i4s
I5xu0VbFsUyLKWgHzZoWixe5pxVoV3f1t1Lwnl2/1hvsR4kNqgOKAX+yMckTA5Ip
lmUDHd74N8+DyLf/STMYtCbMIPCN5QG6ZSq0SrRpm9qDt7Aw7CBLvkLeSOH+8BoI
Uhz7U+RSnmLh/zZOJWZZ15f3e+iNdNgAxpi5KC4nefbLBUdEQ5Z08YjnjA5GqAj+
xLoEe0wjQvmYBVgxsHDEjG1nyJeRQeDYNKneuVpe6lBaedPNh9d4se+CbrqcL/g3
QbmJAPGS4ScIP2p9EdzYQ9FlIU9EzXXAdR5TZHR0kdaFwXVdiNkArXjCxpDg7Y5n
Awtmi/E9ujA8BYWEjd1fEIvP20rlRwfGu5DXoRakqfMtM+jQREPoZN9N8U/NOlV7
e+aG+bz9Rv0v4BtSDc29f9UmhNcSlcX/hqWba9WYKRs2b880ysgFe4FuHYAKmHIe
TqX/glX6YMCw4ltvxiHJz3+DbP9PFBgd45cCH1bRP/6KvDOZlVDmEf02udkxgXOz
Koc+aSsoh3DKUbftXUlKhXssp/1x/7wgkfpDOVPTkeCR5lZX7n86M0HRtq+ljbdp
taOyjMoujjMboTQ4jGq/1fTy9igYc4d6552lMqYgUkMwRTjFRCNrOxe/CE/It9Pj
hK9Uj2J2yubB8Olf2RfAmRcyEE/KD1WU3tgi6kLcXTCawiFDHzHbCSqGd7VNbkfK
zQjvf0SHKAYDSgwPXw+hI7ao4Do+Y2Fpall2A1aMxHq7NtjcV5koIJnco2QVkF0h
FAJXRiU06M4heoPV2yfVPRvqX8ne+ThbWKGH2f0C4KZVNnYRdPrRvTA5NrWpmx8z
lI71f0wmWOYilTHINXPuQuWTisQ+M5KAXg6GMBWagVK6O38JKeSnnAA4LFqhLP4T
zlI4OIhUDhDiaSOmgN76oMFS9Roe7qTbTabki+QMT7m41XzOX/vUQlW//zTPd7/z
BTew1fMVcToN0NOP4WnWibaWUgTeIBP68QIJMCk67kLBf2OXnpBIBVANhVXOsrt0
1qZtQkWUEkU91m9bTmWOsY1yL1cU0Nq3DVeAwsW2/U4wQY8zqBZ7oMgBx3R4x0g4
Zs2zh8AByDnRQxMeHk9jl0CK9h7FfS4njnso4+RYCR73AIsVl24ASSsNn0AjvUoj
EZNR5z4omqVS6TwJRB5nEwGfhGfkxeJLsrYPpiJNo8A2u1xVSQjZDlaVtKcHNVRP
q5USjCLRLH2y7/CMemvnetApps6hevDzh0gf9CJiSHoD7G1ftM9P26TipyhiWHFr
G7KL85LL9dxTU+kLHRvKNbCfPeLVT9P5VHD+gzXfVWzWGXtHSOMkB3hh5LGgTYqw
nyk3VDVC5KPqnNhGB3BN8lxyETbqMClqzenIA/g8YuN6U6eDruQ8A4mDFxU4HwDL
kQHrBvWfO1Vv4KjS7Zgww5ql7DRLmD5Y6p0gO8Ur/T79bShzb1wUDQgqc8bXaWjo
7iQyN/3Q92Me1uYV/awv+qGzSID2FGhQaRf/YawymcZPNkW8Vrpb8sUhCNnliQbM
PKOJ6YqWXYmAgUmlsRUVIS9NxUFntIHNmyH9zv9MTdJ5ijEH1mssHuva31D9Xr4Y
BfqbZnsWJpBfXjEHPdrIhFiBmJk1swXnGf9IVtgLsgmD5JJDqiNbZhKkcyI6wFZR
LAm6s8gC910AM4FV2vEPE+DBRVd6Loo8O4FQqnPT7HSmLs+PFyUqGy8FHnmp9iEI
KSqVkChKMloO4bMNPGpVCAntG8sFBdmiSrZJFr2+CM5NldI8oEuJtxVl9L9tl0qK
US/L2JY1CdyTFksvjgfansrdRVWdNcFi16k+R6Fj3entJJ6aZkn0yTRPksdAQQft
Br+QwHF5hPUxiDfNambFEKQo6ZvQT42E/YCj2UX6Iibq1NvNsuzbNFDC7tR29vHX
/ztnacHuwFwVwyBFMd9PCcJnCG/BRt6iMegA7k9nrEUCx5hXNnCxyg6eKKvIdJhO
nvjSlTIcqkJPEnwuHhlnX0jkcG6DB9SMTS37Dcduo07POHdkqb/yR40N1bAh+OO6
ilVgcAO+A4PTFLfwTnyxc6IRY2OHjAw5laRfClhrQlznLjBQjbPBHbsDcAy2Ny41
Rj20+eLB3Y8L8zAAp4XqqW/4JYaoCz/fYQWOVljg2n24xd39N9L+p6FT4N4Np0t5
97s/ZfHmSJCxWEhmKTG820uu9+5T5I23H/fIT2rueeE+QXjn0ODyAcEi4t8NPafT
HxvB4mRqWCSktNgrK2j4Z2BrXqf8x4HPdK909/z2qxBNQCNw7UKNrMMBzt3hN2B/
GvsYHpdKU9JE6fzgix2XemuXE6/x+KR5e+yn4bhM18TpKKBZxnrUZYsi77wR0fEe
JQ+ig1RHWUIoKcE9y7OTWbjFF0yVjH0de2rJrOA59KHjMFXylINmQJ+Xk1zcvPZe
j40IMmgrm0AZtW5ltZSODywM5L7V7UalcKBAUtd7hQDQP/XsgyypbCzbCS9PEELK
D3c0lel2xxvMhYgPWYJ+bTMHeOtOnfObQZ9RwPeDsJK/PpaBXNTAKklsemFLh2nC
k1YQSCYI/nDV7UGX+cJlgEXgn0VPCHOaa/+iTom2T+LuIvQ/Pz6y6eMXXpNZbDlo
fEPgL72EoG+WKNP0DgVZ/cnq2nOoW3r3/3uTREcNcRhApmOS4ZXTNyaRobhKQ/u1
V01IsugyatfhGHax3lcJeNs9XnaeEQWFP4OwakFq+BcJkoFtxA5mtRdpDYDzuCZP
Lnp5X3byX+W2GiF8EWWdbmZEytq+1o7YTHyNsQb4hn42mIyPwi0xNBz4PG3RAqJO
R9Wnmaqx+mPcAtmjupkuVywyqKTOjWMnfJR5/v7gHwSAaSrcBZBWtb+kE677H8RW
aIRZuHQ1AjfMbHIAKaK09e9kFwq/6rMBwBbxRM2Iz4lkt4qIHYtTaAzu4M5d6rTO
NQRPa80v1T3WClqyl8LPbeVT7+W7H7J0kpRd2qenWJ9LBBLK56zEbfTg2+BtfLG2
q5Jjp0ZXathfZHQdVkfvyxNyg5cjuZ5bt5QkUd1bWRt3Ftv/wXhormVLxqRvauSj
+A5vjBsbf/V6G/ZMrfYu8HLGpKddeMOCY+wjJXxURPAMNIq1YmEDxeDxvhVfLPnW
7WsanEOUI+o2oqEp31Nh/PAZN8a3YJUy3GWb7DYKveZxGlv+AY5y+nH2yi0Ewl7O
NyY3ZTQpAld9qWZQCGyBtEsY45Wt7TRDrPEJeVVsQtq6XY6Y0inBin5RPOM616bn
hODEitEVaRjKol9iErtZRaWJLJDxvWX0OfsZTh2jzaieciXH3VLbQuofOvyWJhin
DUmf7Ry9zuhNofmv5au9MGShxHLkt2zDO2zwf0Z4EAAwIGie0pfavo7YuSIPFe+H
J0+ZnodtJEg2si28VT0xM1KOTqGYoUDjypwI2YZcrGimoKF2axiEVhNIFibHdowe
bD7CsOL+YCYeDewBFJGXUbPCK46KUcGCFrOGzRzddIHELRiWiaD17hLnMIx8C/Zf
SmB2bVgVW0NZmJkyYzfgJzDlOXLwNg89Wwazs6I9CgKtqZJ/FaF5cM/WXN5Ct/tz
g/pMBERBl+W603O4sPptbVbu/uq6xoTdzgnrnEt/oLNB5V7Qn0Arew3AOnDWoR4q
5f8ygLWWrF8kXWYS1ZA4qfofIBdsMpKsxhBxXBSIlzKPUBYOZRymf795yuM9KnTT
CzBPsdHzjf9BQmfzdZe5DMGVtMmJvqDs2XLP2tZzwLrQchL5DJ9pBKD/56bOBsrU
APFj87DRdpIer5gyasS/MGPwG0B2H/naTbzEa/4MvZfQXXl7xPUSa/Q/6z0VIuFg
Uqbt4f5/xrnxrCTsr1PBoiFtPXDMvn3a4jDe7ig2yMPrRrF63ju0+Ohpj9CdkK28
HUEDtsEfMJpIQlE1QZsjdEFVgE8i2ItAZ//fadjb3+1GIiJdnIUQnomIrJelpcT5
yAHA0yiQTiWQKZWb/9Kh+AGkXJUVYP8b3c5Wki5OBzhJaLC4DiPXf9qSKy4xa5Sq
QN+I7CtX6RU9myCNU/+FkQsTMidTdiJmo2eowWsQB3Kqif1/DWwOVrZ7eLa8TAgA
eBSo5KGIW3VYjTWrQNiVVguxfIi61TsMbTviGhPl+ByYm5gGJv5cMScpyT3NaDhi
r+NxXQEVAODs76gwh51ip9POZCFR4oJAWpPVx5omwNch0Q7oBBIisjCxmMsBbmND
nNqTNYf6X7UI5/x4tx8WpQgdLm7FOhn0VYgGxwCtLsWLB/fqSuLYGqA0b7jeahTq
9xLDwRhwwKEFs0lBPmFEWiQt0ZuI0kHq9v52JGli/9XNWlBmYuG/odaRypRiYrwo
w1TLuHkY3Sj0rTwmeok1zDVqSuHYvyuOUEE5ifOjzMsJ7aeBa5R6kMrYMaamyX3W
5efbswK38tFKZRTAhC7+xo/oi/Wb4jzhiKwEW80sKeLtNEk+k41eo/42Kegt/WcY
P6IPyzgShSehG55Vl03y0XopVsrSVLr/nxCzaiaaq/PUqIZ2DiFVL4a15tWD2G+3
IVPvXMo9QUsGA0i3RjpVCRH8jUpCuUaluSaD0peeJT/9w5ZsrqkyqOscccpHwKnQ
eLY0uOqW9LWsMrDSN014U62XOMiUHfRsIICqktylOVTeu+QiJccaGnUPTD1HsTiA
4K3GegqBOIOYUTVvUflLAvDESGHTLzbedEcDxD8sgf24fzey/rrrFd01vOcJ9Vea
wWLOj7GfnhKjfquQfBkX0RkRKSzV4dBllm2pgFIX+UdVVm3GaHGGAUNqp3YIXi5+
gZ6pxFedPJxYRcS+tHRyukKIdyUQckwmXCkwAAUPyQTIgr8v6fAZv9o5gRvwkL73
8xpbfDyTGAgKHrg3OOeKvnthOWWSo/AP0pPkK/63sOpJlWAMZY1+MAn+oMVE+Gxy
lIXiKlIIAjm+ijpqiItZ1iOzb585cHNffiQz6HQGrPZeSQ/CW2E7G31aF9xxEpNF
s91fKUh7KUjN9ZkjWeQjmncDzVbF8NO9hfK0GciRZNnqZw5PqJT6+dSXsmPmwQog
tGViEEZKjm35fuqgINhDudFL1KLciJQVLuO4b6zKzve4u0k3JsS8uUD1JqTHPV+9
moRRUgSxqYkKnBlnqUG3Bj+/uOmAV/MVjyGyd2ZgSVLTT2cfW4bbz96jx5KSFmgV
0YIIdW8Tcabj4JbtbaLSFN1aFj1I8R3xwH5s0zvxWOZhtH8hCF+qQ8kyQnc2k/dc
hKXGXUwh3/+Dz3tQ1xGB7d0fsLFKugaeb29sMHAEyBasFFfkyi8t9Ecx9bRX8tZu
S+dpqseMYhFrSWWwHGCw1dVGiOwY928HNkoQPXjoZCWrA7+Ekp7A2DVuyt6lEFUo
d2+OQKYTroRUVi4fpFrGd/grj21CeEROowJOXz3OI9wCOP6sGCzCh3jkRu0iOWJ8
PuJJRKljuI3qEw++Dg/VX9ZxweMq767OwNx8plQUzu9iI+6vkjBBIWl/+nXnGjxl
Gz8cya6sX8sxRW16RHzvgS2BzcToq45mKVk5tkzI/Gl60aGh4tGH1goGMOBm25KW
J2Wje0GTENmnnKk3eudTaPts9+ewc/6/AlDK9z/nmB++6FbYk5w/2DYTnmhWorF5
pjN/dBtL/zRvNquQYM+TbWhSEHKjvoCxxzc06nwrxuOrk7CFNKsrMJGfYG5kACyZ
0Oo7bXU87IzE5fdNGSVKSGiXUj/qxoRlC0QhXjg+G92KHzKZKuCGEesN3Ji19mUO
0AKqE+Gj7K6mirF3FThiXEY/9pUXoJESiCHZgjO3GG8eH9c/VCcwCw2zcK7Os4Cr
SIZ8V7LEAp3jz8IxeUIw7cS6WeGGPNF1fD0tHBa3aqk/4rJUjNcgmRkr60doziHS
weuIajmtz2FzZDKDqn+zdz72wYPji5NdXKFULN6/0cWpNmBZ+p9n2RX1JHDeNTqt
2RPLVqAJLxmNB3H7V0nIL/hGttfQCdMRKHjzNH00daVIotU696QlXE0tczohFH+p
8U+Psjt13OvMEPstetjQ095KIvi3kxnWsdHNVCoJhdT32TF0LoggX3uYwbLbPUlJ
7+66AvCAIS5ejHTPSSJFnBMsL97XuxJuS0Eoxfljt2IJUQocrGVQvf+W6XlglXNc
LF6jh29I0lgePlBe7CiRJ+iAXMZDvFFvudxgasYGaXzXMFF0dZ5sW5GM0RtJfxrW
Ur5+9akX+GvVlupXeAG86GK9te3HGUmtfCRozeYN4VK0ee0FSLOQZiOta82K+9z3
mB1XR0lSWvAgo4l3OdF09koOGDAJqxPRDUQ15jHF9xvqKbGWr6WEgN+yKPNTkYFI
UvGA1qb8rsuuZcz4N/VPqvhfP0hNkrJFFD+owNUUqm2OcXbEUuZo0yZv3C31QwXq
2TfubJuYa4t4Dfa+wGMCSpgRlWJTrsKk4ZE1bkYqFx4R6GVLeGQVy+gPshTX18eG
tguhMu74Oam92RkBDYZfo8eCCItN0KfGLIoYY542dKAi8KJah1bQDlJM9liir7k7
b21fb13v7PIjv9bN6QJnZHTKP8sMHcfyLhvei/hwNBdUF+HWi5Hb8gsd+/3BLp+7
o43N+6wRR1grK76lHWMCUaMZOe9M6vQv9O5NMLlfpbLfLTmDgknMwkLcESUcWxmC
QYNDRrK+Ljqc5EfWtQPb3ayzTpwdACvDVap9u+5zSDhseWpbVDK7GDBbjBv1WZ16
mnN+pu0OGG148aTLK54+oJlYNEqUzkDGSdMOC2GgtIbQIePp6c9jf2zXXuS+UL35
1bZ5c0Jvd8KhkMoGrsPTN5Fh1aUkWVP3bNVLoR00Cb2pjvrPdCq+ZHqmihbWNthQ
wNQtPbJDa5TMn2+73k1MVDCGGKqhB7gxZIDecdgHGtkXp+mSAc46qZuhHPCP63Zd
bCSAXuqBLjncOAAtQJpih6Nkcw0viXgdcJbftIke7MPcDkG30VknYHxJpisD5HDt
EwVM6PH5aQCybbGIFcQHovW2RhZsmsnH/4/kvG1R2YHfQi431G/UMQl70sfrua9F
xSTxflJ8y5clSYQV/wS5gNg5rBiSXinYvSndNVJL7eQ63yZ5oYjaL16FAajeoqlW
pAT3eJlQZ+lkawGdFHUrzeMi4QHWnfSDmRYR8gNnqUAm9atj1wVUXLs7DHmnwhdy
YKCwaonGachDJDvHS6NF96Prw7dOZUv5TCjIb0epwsRdj9ucthbfoVIirH49LMo6
gEPfF3Mp7wSw4Gvq4Amq9frrqvcZ0N7986aYVtezR3jF+3P2hcklU9k/FiLyqyOv
ceXxbQdEQWYkCwSQM1tRPk1NBDJxVqEH8rHLuO5UKaGLsbjhEtLG85zKThJWzENH
WC/LxZ5R4SqOu0Hxj4ML8RbsKNhf0Gl8pV/RsgWsF6I+pe6y7CA3jrJlZ/P/uquc
IYMn4SKIFoMh8cFNiSL0PEk5t7mphNjiWlzoyq9VJZm89Pk7NuV5jY83357AfWIS
8dCbqCeZ2QBVWrEfexE3s1/w0p6O3irTt1lMZpDABC3E4h+P8dBipFMyECIeifzq
Rp0bYpeyAc80E6eHIVc9pN+Bc2eTJsQoGFnW0DOzlJEEs7gTeUqe7RdO0Hy7sDlW
fMsBbZJNWTCAzC+4Hm8cNmMQ9tWn2M7YF1WTDqOnWjVGp0GO7upg4kuc60PheAj/
ftB7G1Mwzb98WqhhheXMNsnF6p0EuYQ2SzBfk9g2s472xJEDVmZb49k/QxcVfF5Q
nXBpbSgc75i0xLbRgm2xwu5ukuUvVRgL//xM9lvhXmJRPSx9QkhBHHkF93xmqoyY
3vGGq7+iiuBZBymvqZRUQHR75jsVoxcUSv8fSIJWMD85wD1T6b78tPfyxrw3V7av
6iI/v9dNQSigNbqiJPRl//XQ9w/PLVDENOCAJXgSZ7QqHKCGK0laZDI5ofd3F+De
Kg89JxGxjROL6od6a+WvFO/64e9xCPFjzwXueFo84n2nNoCZ9xRCU/sZzkyyrvxr
llh25aP8F6vhazehWsuj4IegxwppAzwcE+nhyqzP62Q29yl2KPx+cNOwLj0vukp4
1GCtwBM+z8EQY8Fn2yfB7HCRCuFxum5AcllLWRgwR8wvx1Vova84eAdgy98/YNI3
qCtWiMCNRgAPzMePwiha4xWmxCnihS9QRoczma5rgPpu33jpVOylXH16KQPicUsN
ZABfsfPYImiZUabAw7cwIyLBWxHwVOV2M1oa0pDyFYUJwy8yJ62T5XNL54UYpLtV
F0eh//24VIcvLsfJaoXaseALBQzDnUd2FjkPunE7ZGZHJkWXaZVL/Ji+D24ilfcz
j06YHw5+xZS4iFCYBjSCxOUlQoDE5WiUm+Oh9Odde79v1KiLCetu/tZJx2D1PNoq
N4l3kCQrWXs23LO2SpYjfevX1rzkJhlKbK0Z2G0kThpOttxCJHjqkARB6pFAxzY0
TK53N/dkPEhejddULIjyqSn5c9mEGpmaUjU2P6F+UF77rh6hAU9xFsoaQU0bLrKP
uVTY8RZwcpkI8A2Brlty5+DaONjgCQz3PfVsMS6BhtqnHABipPLqIRBYelexRhK9
ILLw2DQKapgmUQ/MW9mPcZzZzajIKkdbIUtHtkYGbi9MIlw4Nd0xe1W2Z3W8RnTr
T0SGTQyEJ3rIp9kI1NjyFcO5jRjHe7AhgT+D1n717dgN/rHGZ3YXETKyjZTWPacT
O+5xiX8Lu9BEgs4wOmtcaN9RB+zuxJpz8TmX0tZleZnP4UXa8EsZ8j7pPjD6LZ3X
T/BcSaKZYOSDHTXaEAggQ7VroQ4/xMkkTgYcz9E+qDY2YLeMgww0e+D3wLsbA0K8
RiOodGV0+ieU68Nj9uxU1HzTRWAz7I7SHPz+akzbvkKMmW2j5t/hirdMwTM6HsLq
iGzXAAh839NgxaE+/yVUIeagWqE7inmuo3QgJYb3M3BZLIzI+4vMuxNDFo/CEfn4
zNqrdzAKpwJuwP03fn/o6W7a6hrZrPjEqSa3jXWJG+lPjVk10SI7P+kLpyeGC/BY
oiJ02GQF1eWuHgU0CIVlh5GWnPgIDnYVSafkF+Nu0B2jgRd6duSx79fYLlxcWf45
QC0jQY2SjFEQqK4w3czwKpQ6GxIj7ZQr8A9bOGVuLITPvb4vtSAR7LkyW6HDrzK1
gls+epf0994gHM39lYMBXxfihEq/yOKwMy5JkCKP58l0buI1L14Q8I9ff1lI8AW+
Ta6JIe7Dham909gDjUX6TiyoxLm8oI3Mj1Gg1sXQJ5nPuztZNLONO11L8rtl7Weq
87wIElQ7SoqHfDy5lyfcHlvePOP8dKZXY5ovck1itdTIqE+KTLGi2Y7v3fqj3y8o
mpnuS2+B0eVt7t9+P9pSZmCIBUla833vkIcWCMXvPrdtKWsjqmMgLajB4YP788HQ
UPTXNaRGmmin1307AXzpPrMnC3bnj7n6gDmJ0WHSkYIztS8hASiDbf0lQyrpgAGB
g/aW7/oQkKzxt0AniFh3uYU05BIXZnsNPlDwpOFW7oj1pPs+GlGhMLTEgln55VpP
I5zJmGxOamil9pjW7vg2jLRxj8QvhjNGqcZ+PPAvyoibmPogf+YQ4dvBN91FRGI/
t5P078/7agWdrVvPJAE9jNT575fdwQDpFXGtsL5d/zO7gzIaMRLyXa9A6OQkWJXj
xuIYhIoRaxwmPliDgoWLs/8rIXocRxStVZCqiTmrye0AR4dBKTGURXZnrttkdGyf
871ZaMVgWBiWlqeP8+QF1zoOgiYyIDZ+I2vFZ6BEAAwbGiYdAuUqEXQmBZm5HRVN
vJqmpyc5XhJE6eVPtrX58BBfGNieGSX2DZfBepbpEMPZpQeLdUaykmQaQcTDQMaE
NxrTfwhsAMw9ZZL6SzViDdsTlkKvvXPXteJzfK4ADz98m/KR2h7FAMk1KiV1ZSKS
jpcX/48I4bAMEtARkCLBVxvpl50q868vrG1e40RUrl2kXLmAQJpSvzZ8vtbFIHOh
mfeYP0E3ORGChibt27jmA5gAroLg9tZGO7A8gLHGTc3MzLvzcVmBuugrTasuBWNB
wHHHMv5Hn/81H6ot+vnM10vtZ77N2mBgd2ERyizZ3sCUmfyqbnb7GIOnmsEXR3jP
Q9mZNRcwEFLA+Lc0LvpD/+feB8KeH6NKPqtFPztTOMkzBgpfQPVHjyk+//tcn9rX
UbXMzClCDFHO6ryeNu/NBVpiKbVfN+WVpJw0FddFSvlvikbm7LEu2Jmsw3oqS5dq
ndZk3EU7/bFgUfHH5yj5e1jLwapMLxPTg/HMWyL/fH5jE+BToyto/QHQ7lRHnwKz
B2mxxpTG2wyqlyoWbY7pQHwtfoM3Ptc5iNTxIeAeBBVqUEBh6VUwS1fKvoF5Z3sn
Dtx4HyEgs7C2K/WjTxNY2/Lp6MuxDl8MctBVJvPl9sYc/YUIY8IiFm94m8AQjeOJ
nTt+u0/g9jdnP0+E75ck6R2Z0v9GMC8r0riCkscYB5ZfejrPwNKiq6U4iqleSBiR
Yi9LEttkLEj8pcScK0xPmJSCD/AqZDcgl+hS5PAd6odg+8byqWe2F9L5bJotohQT
yc4msYptoJpFTjLglQLVg/EdcLOCX6R4q8/iMTqetRqzPeCJW8SiaHYw9fLdEC8l
ZRWRqAO1jW8XJsNOfRQNLue406EQGVU4ewpabnbY1hyk6sEU231RKXgxFFz82NE7
goWFkfmIOennCeKZPlSGJpiFTwOXDqHvLUxEj3v+g0i0RaW6WzKryFqHln85A9D3
ko0CqKl2/PW+mXN1aLbWOVHszARxSukarmxvUkQN0ghBj+EhB2BslcX3ta/xnprE
Puyutf1sCAQxqFpLzju6gYfjHxXlyhAZT1d8FLFtAumaT4nSclO/fRfPn8arM5Ww
Ai6CyRM2P+vYN4qnwW+T9qv253jgFrbsh78Dq3HewQO5AErgjcPF3TppvniJV+o1
GqvVdnWAfv3QaYzCuLCSqvjiqNfio+ddiwpY56jNBzSyPp6cakt/i1jYcdkLmlPA
G6RLkeZ1XWMsjgdw0SPrimJRVotQjnUmvl+ZDTEh3IWQV07j0f/xRyAFSHqLPqwt
9U+GukXecNvjBZQEDYyesXK1GJKetKCGGdStQEn/e1M2alqgZ2N9ccZALuHGXFai
OXSOD6LFNnIiVbWFKObvGZ3bVijp9b8VX1dR5IfsDphYUg2sTpDb2wRaX9BSli+O
nRtyXZz+6w18ah893cfxX9C+9t2egHB0VoMO4E1NC9pQPyo48S3atFkTTovZF8Gl
xInEDuJ7yXv0ZSpG5Y0QAC7SUPbeeDusYyHS2FWue0MNoC/NTHsE8vV/K2RXBW21
NmYQN4l8xx/3GskDV7wEqIgLe9x7fGjcPZiK6PXNkTrjFxahvvcnpU9srmGj2g0S
fHkxL1BcAnmRVunP/Ts61s2WX3dYDtToDlCyBCuXq2e4yZ967+g4mtIx96hf+zFY
8tRh7xHihZgfLGxDTiyl64KWQxthjNkUl7pOx4056yZlRSQyAVAFmdz0guC4rpVH
I96VR1VecZNAnv/k+g/8uxzdlICp61VEajf36uwDD6DwYLOGmT1/2auLVbv/tbQA
epMUxq8vJ7zDjNEPdABNESB033rfHjmrlic1RcQRGee81oyX/4X4js0jsMSFEqIc
fim4CSAfzoF/eHnUUS47neiL3Iirm2ifM4x4ebWlPRC/aEI9CFhzyGeXuwV8ZJ5K
fCN9u3sPA+3SLeD7/Mdcm3JRIvoGdEYUhtf/8ufPYkE1saCJmNfaoyKucLDBqYtw
XnmqAPhDDspoAbdXEZghKcslSsRoTZDc+PPG5z7cci5aU/rVP7OjIWtoDAHLYzrM
FPvtYCC61v58sgtqKQQ3pTV7rxbl7DB84Y60tOtP+9OBraJE/M13KKvQyCDq9K4u
sZ+nIogRuxXkn6aSl4aXfoG7O2x+h1JE0HxQx4AE5YPLJK3jHc0UiMBOXyWkpN8p
CkfaxlNcapYzamxmP0iZ9Wgd/24n8rjziJ43saOqKyhBIEZljGFzoAWzXMsyY3YR
BsXZEx1IM/4Smk2xAFjj3wYbAQ2SwW794sdlEMX+L1FNHxmU+rTkM7SyLwaZBhBR
uapUc3/RCOK6sMdGI5rFNP0sFeK/MU2py4xBZVH0pgvRGhfWs0WauDB33hb3SVAH
pIX5h/u5t0SJh3ZHmgzSQXaePGwEvOnjM0BtR7Nfq6iYOXhxcG+ByoWPyzQmciMb
rNWu7Xky7g6zHuRtzZiL57qWXqH1mMmbFfRRHW5+YubAzgzB1tk/gH2hwj3fjZvz
PJ8CIZAtaWv8DPEv62nAyIdaQunT3sHOhUBfjRb6A5mupYhvMtZSHBEXLoqfv7yS
Y5vuRadP1RHIk5UlDIFUechc0ZmcmIR+GnXyhbOd/yjZw+OL8XYb52GTJ4Ygd2y2
/P1ILtd3OZeo8yGN4fd3kiZ7p0PnGCUqh4J1mUPEK6PDuWzPIoh6vZZtDSA61ep1
hBDj3MTPzKHOjbwvTdmTzy858tw4HqTrTc4q4WzL+YDKEbXKcztGG7roUNsi4eEy
0O2z9rEc8DUtptoiomBbrmMDPS65/++yWs7mHgVIf+yIvjrer2ds1DxmuIr00GLV
W6aPrUUAd2BqeaLmJ048QLEUVUdRhWWPLWG4MAOU9WgRHB97MhMRcUmvDD1mY2kG
7QUWfnzMqr+/9W5fRT3nUMePGDmaoSr2VP27xiebyB/TVa/5i2hyvxgUdkLurNrF
eZIsQdcQrh5u8yYI9ChcfHMa8Fu4p9ChxIVnAlT+x8CiGSt3WgDddzYJi8o77eNo
63oCeEntws7Pk2sP86BpxubjQG9K4HIbrIkKSqUOYhDyQWy/xbd5ZDDqX+4PSqRJ
O38adtUSrZZUHIx3Eg6tWdJepihg4u1Qc620aQgKXuhU+EOEPQbnKHK1eE7zYuYV
NVML639neXA8E/Dyn5Jj8szcNF72vOyJbyggW4wpBoIUICj7e7dMwdjsjYErP4VY
mNDuQGJYnA936Mm0+RdZ+42+G5csQK7mQMKdGlFmK8vW7BZRo5WmSN/mhZGAC/Si
ZvzMVyg1PQsIi2kpuKTL/TR0YrQd7NOeQQW5mKOymJDwyshBXc+ZkujOfUKsuhs6
fQRqyoQu9ujq5FJwRGPqZQgd5fouR0uhXRuxN/3ubxKiQCVV+JeTd19UJUlLyJmK
3kmuhywZ02W8eFb4mZvlNx37hIYqnPgWVNVODvWMdNOjPMlVjdv21jqTAr9cNuGw
oS+tD85aRsKwp8FHYqF5ypXBsR9g1bfbWBHHeKxEVFKz0O1d4I7Onn8g2x2r5JWB
YDKso5pvP1s+iEv63iAb8uRXaSsokdfOCE6olukWngeLoUTfUsCR7984M/GnuOQ8
R1ntNFML3v3iik5ubiMR75oW99SYvCVNcQqagoigqmqdzYbw4WqCPsBfIJ+gQHUg
T0RPJIwnKSHchOQ28O2LIkrPx5Qd6BK0CTs77M+STXxuvqoOScSy2A2vjNYt5JP5
9Jc3E/rAXPIDzYLZ9tBmDhdZ3JjbbNFLL04Snf1XwYVBNt30jZuFV9r3bQjyFNdF
Yh0pg2vTTP/ykYs3UP5o4U8uO0OnEF6fIOFvrPaUkl3MLrQZr+on/+lkW19fKQS8
LVn/g3K/D2ic2FokTgmZiiPBTAziTaRvfwjHBXLb0xpXkyg6/9NEozurOl20nhXA
/tXeZT0r4dCo+HIWw0082sFf4cAJPFnQISDn+9BY5KldS+uvJwuYpKpkmAUg9biJ
FsZ19U8vjbZG0VbHSbYm0g1/5iS4gbbrMGlumT+lR+7QUWZAYutVoxPw1lxexGRi
3Q+eTBV1/2Tbty6OAuMjmuzyclUf7bZO0Ckfcvzzqny+lYUNWbVy46bJ7STZitfK
EkqC/8gakVQGPPSWy6iCBkUS01NgfaVaGvRAEWUOLzYJxmdXVlKJX0Aqv3/mKRdN
SkQbuLDkqDc7p7NU9V+jdV/M6covayHMYS9bEzy1YFoIkta1k9sWQvzQfxSMZKHh
ZBZk7A/XI77Tzo8Ue8OW7GJxQi7YdBlyfFHu7pM9ACZfhfYLR12xErTMRVq+f767
GMkMQsjJotI6widoxU5MjfiLMKkfVktvnmsvOHXoQ3UL7I3KKQoYpyK8KEMAYwQM
XmwjbCHXiX+oszSogB2iv6stfasN7sZm5TIlEjiAKcC5+sYSdb5rc1P8lXBtGOmn
bnueFHibW74t7Vo26dmrTn/cYfxiNPEzF0mwgUwIt09CAahqtHCPvxjj4vEbSYBy
K7nbB0KJIFdRxue93FuKiLzENKSm3AS4AKVabbfYp1f05fyiqkv/Ca3R8sLsnA/x
demEyym50ti6Xg9zZGygAg3N4iJ1GpvlMQSMdcxP1z/VAeRGl6sMGFENR+LQrFDP
phveYOQYPKiG7z2u7jaiNDlXKrCs08Sx+mrXrJGdTAl3CZpbIDjCRoFtX/4zXfdv
n5Jq5xAJixtD3eFiJkD+tUfB7x6x9c0OJvU6VXcS7G2glFW+BoX5lC1hzQVRNp0W
plV78tFXenlaS6Wzc41fDGaSyfta+6+xq7CBUsN5rzlozLp0yLbwrtMud0RFiaQu
dBYWmdU0+YYPGlSdIfPGJ2UkM2OAWdzvja+Z6a7RsfmC18Jftx49vyzVCj4MdcZ/
JGCUOpf2zKsSpO2/cr1CsXPsMX8eSf8gNz1I0JiXTZIxEJ/8IccRHu9mpSVw3hlm
Q+dq5yywBJC3DH5TBvsh5ebzVnCuo6Ysmb4u8xrfWeCsnjwrdJnkTm0ZVMtvdZ+d
bL4VQP+JTj2wccoQ2XKWF2WMPHd106kpHLfnGYdkxbhPYb+poX63XtB70KiSp1oj
5kgcTknmWAiRjYTRdIJypdpOlengNiMQn+2L4RNZVo3xnbJbKuBcqEMEMIlT76eO
BTX6vGtIluuXdYqwHNBMnOy1KkggyUnpJz960l0piEh2RpkHXmqOwidMoIVjoTvf
kz7DdAy9McDHEOE33CO+wr7F3MMxrOnou71N+SYm9uoUT5G6Gn6swSdGo2s//Lf4
Wc06vJtG0SepPS96YEi3p8qBtpyNqnOBWBStvnG4k4tb2/3FAiX/6wM6BC+KYnIF
Q+ZlhSIH5IC7UOPKFhJ8JuoMWbM+v8FPKqhlyxB0mpad6pwN3mNAs8vbN9Q9DPK3
ZTdflOs3izQwDZN+C7fFdyAdPsxF5O18cWOeL5yepdMYS4CNEu+xyQMim/9WgKdD
lmU/HxMYLOMRBBnLEH4lndo4oA4qWcpB7ZJ+qXOteCTD8oAsDu4rXi1ptzn6yVz8
ByBJNT/WHtnqSVWScvNeJDOAMM8S6luPF8507PEtjbE/tYFTQ6iPQZd1eEcvVhgM
Qshu057Vyd6Xj8sEFBDrxfg0fSwHO0qp1cWNAwRJ+4jFE5McxiTCnIWzipaFQ3x3
v16Y0DV44+5+s0BU7gKMJYXVy2mFVgQUJIusLHlM3P4ULzKrgCfG1pWjUeG2QW32
n8PKyY5MSNx6DW7hgU1gsNUgwXr4QdcO/SbC93sR/MfWzNkRKg/3E63nsQ476/lH
ePkJ5T0ncakkHuNt9E5FFB6xyn7S4K0FJHz86rbZai6mT94NmqKGvULaTu23K1DY
UfyFdmRi7xxEqoMwcv5o7WLA6qBMUq5Hh874vtOXd8hwbaEXbdh3VJI7Nz9hOgCi
wqXnrFBhAPURliSziy/cILg2kYLBGX1TuCHBRM3dSNospb52n/vqujgGlsnP3uXi
CwQeWg3vS4SjmR0hxFw80ytW8WII9JDr6cq0TXAoxocnDwoLi8OlDD+G+ErZ1avC
sUyLILDKosv8KxoxT6BhUMsy3yHijPz/Z3Uz4l3/eECyJglY0FldKak7xfbXhADE
6wxRE3USZOOfB7MuAwbxhu2EiiwM4Uu9fgod5A6eTTn8A8Qy9XRin967z/INWLpt
WbeOP4HI3Nlo/qtEHqUHKEIqrk4mwa6yw1YF1b2AGmbAfqdITNuzT+CCygK6dbAl
/c2leKmmM2GIPiu9ONkfMKuFW0tBQCQEu97NgEjKtBJa718rPAO6CbuFLU+4IaMm
f2PMkCWbVomP6x8F4IKIIWnxGtWllkC39KTYdSNJHWK2NhnMZ+2eLU2Int13BG3U
XRpB8XXLpxHQO6llhVEv/HO9/2fQtJNKkHHe+Mw9EUmKevXP9ZKr/bbILjWPjUJ3
IMNNZFQDyHoD8XWPgIm+GbMev1D9pLkJJxPv1Gbskt0faTG5lZv8RHIBJ7LjoJhn
QRDcPApU4xGOyi9oPjPJyGVBn98pRj+TJgBJtQI/CKaR7eQZXUCa+zPNuIdqL9SA
REq3HpPpaOLcyxDPffDulbOlU8UOeab/h1oRPQlQVFsAPMkYOfsIqNODhyN/QyMz
avJnri9Mqus9CScBBqloBg48fTQFegav7mwco+JDYwV50xhy6v/5pMcgyTcntWQj
+CjMfpopqUZimx3V3qmVZ9H+lbG7vaIoNAfDezfiW2LMKLkRQV3D3IKaZDdAAdHA
FnMmLSL3kO7QrlGyVM0baVHGO/k0XNSbhdDc/iVRLoLLJnAz4ojPaw7cKwiWHS7o
S8U1Xsk7Tqw2MfvhCdqtUzne+ucza8y7iyNnp9k6zhztp+mHiOMxMnPm54jP9luh
i+1hd1ZZtb87IveSJUF4Gm+3+nDM+8xfdKjRY0ua66fwgKCXxKJecSjIYZYDQQhd
o3nIzMWEyurhHnHnDxXzou96EddlbkJ5xEKxozZeRex4Mcezya8qOl70gY0WS/1I
dbEzqR02aRHvti8o8eVQQ/vgWmqjU3MesaSVe2N3ge19UGZH78okNKQbsPsXmrmK
VayK8Uf6CX5Ts0ggqVamo00Fikx7mi7ZXnTSNkMfHuyPQy9dobM8unxvpuY1ijQ7
zHkxgnjMjYrdrFayWabvC6e5GiCC9/ftUYmVWfIALD6KxzcMQLiLmMuUgwnhms0C
b/paVIcRmt8ZYC4LuFIXGyLuni0bmScBS23p5UKZiqvnJmA3rwZNiVxXfN+SGX+U
8EneIYDs1WXwBEUaCQjSMSOlbrea1DMScHYsksEAAMhji4R53xUa2t2YRg4ggPEz
2V94OAFubOtxZIus9ZuoO4XlTHmDPydBbIqexb062AKKwqT0Y3HsLj7fM1pPaBEp
TljdV2+9CPAV+mWsBsUA1ZCeUsF1v27biCRaz/kmwa/IP8nBCdcm9mQ6aB8fpwwK
2LSXkvMdyJaqcmgQTiwz+Dg3+irJdnenMTjzZiWVtEcML2AMSVjD55VMrSEY5WZ6
Rizr4q7HgrHcaNsXs5ZG1huOoAtltJU+tQ4HiuPV9ZLoW/6VLy49FX3vjJ9M7JB4
VZyxgy7VeQy7q3yms10QIJPtOGDu2tkl9fqDtRNuCeeYo+47NC5ZuLVNdnSq8PJr
90y3VATves9n44YZiFCIdeBFkuP1MiD5/51f0mjgIkFKNU0n0nvO6dTvS0z2U8Im
HR1XTcMCYocITWad4qmXDiRcQ54cpkU3323l5MKq/J422CAane7kp/JPQurjiAvq
dC1sAQmTCF5SkLumDvJTshsIeb6GAznjVKPZ8n0PM376r9N8eQ7eOo1BFzR6rkMA
alvFdjUt/zgcyNUevD3xvPUqfuOCoBsgM6JAmwSXVWLOvUE7J54urjLEXeGXG9ge
KrxE5bU+iUnwDLhTz7wb+Zt11y+SC3T9sV16r9bgnIOSfi5UWXX/3I2khXzL4lmH
6MdS6VUzMPCUemzCgRY4h6uj+Nn4mQ50bw5W9dqEtTSjand+4Af4uc0v0lldpXBz
18LmjcvA1vUVtOx1mUV1RNGvQ2n5PYui2vBkrbbIyh5qVfKhhyMqjjgomKPxgVnQ
GumkbhSc0p58UdNaZkbzqxQ8GA5lEmFcwCY1RDGxMi32TMrpzkvLLVN+Hrh3QFL/
jZQMa8q+P4+Qb6fUXkZUcnEsR+PLEcTO7QR9OMmrLIcdFMc/SljKOWOfpXUC0wOx
TVRH/xhHg1igkY3oD4dDa8CF/LyRFq7WukvcQ2wu/XE9J+iZqKBgbaEh9+OTp696
tkGL2jJnN5F9cagYjT+v19HV+mAR1jRT2rod/0QsCIJywAwuaOnwOnoYy9YqjwYA
nyKMDFZme7Tw8lsgLOuXHyXrkCfudF4Ojdb/UPkHKnmcHsn2rKmtSxwOwkuZH9NP
RCud/HXEamSFXy8KK1ITDx+CRSvYcUOhjVlKLXlcCehHL2/p2qJ0QdvuXWYNmhnj
ZeC+rRiMc67tmrdwm5+ACGFG+MKoPiu+4dpbavDAqwXm9Jz5TDukYxU/XNzLFKQv
y40r2gR9mJ6kKJSjB+XGOh5shIMmY5kFnr06RZKhZbhrDdEG5pNH07UNCW09AZqc
tDySLNyCpxhywVbPT42knpsjHCC7lGuapuzAVvEllnIzmlq/N5sQ1DIf7eJca1J2
JwRowS/MasiZ7vQAC9XwYUBw/sjeTM7XnY8TDhz3kf0ZR7eieRbrjulnHpGYalYB
WNm3DWixn1vCxw2cK0+AQ8QG8x/n8g8n0k2AxHR3tg9wyzHqsV1mwoB6oD4upwCM
+obPeGYtVXCzGhI97FPQ4ckoySa0t1kwRa6oE+x1SdsL+vkf/Mw8NKj5eNrEnUtY
CTozML63MpsnarRxJDhWYaPCRW+dlFL0C2zI/esQ8rD5Y5qm2Ke5WA3+F4LpUYr0
b0HiTpRU1CHb87MTD5QLJ57Ukd1WriaZKUomrUIsJHqvaTydHJpe3WHVXWJqGK25
xAAbMf+0Qn+bA6CHovegxsHHsW96JyIkmDu9H9Y/wUdm0l8GwFdtRKT8A4hywtoe
xg9yHknnbhQ+FS8bPUj7V5C39JGsulQbjkOImmZtgr5O7wDqinF4h6UKkm9VOeYk
Yu4TNIXmAyjKIjJO7ByWmnVQ84A0Uq8dy4axgK92a09f89cUoB3eu+TyjS7UnsSw
xL4NFJ0iAW+/nVjPFjTxr9z4dUZnLp0lKoQhcLryEovlSZvqkoj+8M9YgmRJC6GA
XMXlnYfwFGEuH6dF1dYkQvu8JmiP8tWZjMSx7ZlHhlqUbIuthxRdmfaIvfexJe+y
nF7WU2QdcAT3i//hIh+WFRxlTUvi8FR/ZXj+2+nAGlG92vYp+5RxDz3N4n9IgAWT
0FV4JYyzw5XYkytftzfXG1M0yfuOZAWdu+DGarzEZ3q5Ous50TZWKeade975xZYB
FjgfnkPEo+lRuL0sm0jEavdSn1nFrShU4tth2ArKBezatFZyqBB37BZzM2B5qMRh
EnlNJGzFz7qrx++cmO678d6cttnWjJJ2Hof7x6d4Xi8oTRF6BQeRvsb4Vu1vx2PP
Ey0JKSdBQ+HgxZnCIH995IU6hbZr1mXRzklkYLoV6ep1VnctTozMfD5uvASQ4nfV
jw9huwKvBXWfXwCYqGAfvK6j0B4ZnS4WqpGZu554Z8MK5+uLy6jjx7ufXku8ewGr
xBytUv5i3p1snZRdC6maqzvoScvITVrNh95RcuLWk56XjrxRFC0Z6cFfKXiAHtJS
JyYdNFRbgJOQGd4lqP4V1lr2IfqvT00KvkcpbRAX6+WzXrYlDZQ761+UyyB++xRn
dVW8GaVswOU02MTxoZzHSmTFNBLV107wQZ7x738/6tURism0G+8Lz1FdduPweTVr
M/g8t+rLV+vPaZsi9WcHpbArsR4lj5/GmC9KKHVsgh3EZ1dlX9UDJKmJR8JJcqB3
21q9OyGduz9p09L5J1fKKioxBVP7R5uG+sf7/XG8+sLE0P9biQwxm2Q6tY8d/SOy
7XnC+x1p3YWsK+H72xM07C7bDhf3nFRf0664GwSgbiUckEvnBlkTIekF9JxTQ21m
vXc+3mgR3lihzplHMq9gfmjxcKM9udrlKWy6n+IJDrwcaU3RmagG2PFQK9oxZC18
I56YEgrXJLm93c8IhLGhN23t31lOpq8MwCHva5PXuY17KRPrZmPTfJ+SUJTyO9zr
Dsprfzzr5mP7GzMEwlijqzd1NyNJDVQm57gU7rHENKzDeH5zd1nOIJOnoayzeKMc
ac3qdGK/745iGh4nQuySe16DVa1U76YvIEPIWWuEgr1QBlIG6rxCh9Pcy3HMnSS1
mgDlx4Uy0cbEaAZGrXjzJP8YawPovjYRf7eXTmkLbaghG3FGy91X/a0czqAoEr8M
WuR5mJqI6iaADbjzVLbAq0IjomxEDSfH0Z3vNzBCC15sX9+GkgwGWjLWGNmEomyr
tQEZvV861Hfee4wUtJPNzsZswJ7TuyS3DSKRCNRLJeaKPFwItQ1FQGRYFdPJmIHZ
01Q6ro2xfIYcuKSdfG+AVG9KzCjuU3zLCVNoqjS1Nhk/XA+14GXGUTjOkBMQcPwA
LSbZkvlMIiwyVtn/tEZ9E1SIQeJYsyqkU0b6OdCihhSoees1KuH/LGSfDpxOOPPu
a8kFppTo2bIYX9D6Yo8T7Y+x3Vg40hgSxwMdYiSZeELMM036R4kDL1dAWv6L3lW/
n8UqxKBYLwmL3b31RalUQxpHBjQ4mX5e6TCnXbUXegwS7itZa722Dz+WpR6PxAk1
/5bJgJfksMZb++WfZETwKI5j25i6Jqf8FnmZewEVfUh65ssFIQ2qjWVSxQPUvAhA
qwaLUuMtTqZ5B+4mp86hnDz8DYrSbe4CCI7dM5qCVxXXa3W1Nrl8NW13jVjd4cwv
IKPkNuC0qtc3vmp2IXR6NjwY3mYtez4wb1iajQUH/rOaiJ+9b1XlGBy/m+EZ8kry
4UY4vwQkCRgW5tKijiPK0862XFN5ZYg+txn728trT9i8PAa8uoC8KXwCqgVQX1N2
MY2Zh9qcnJWpPy6GD7iyOKBQWymgBo6UmWK7eAwMxW5osqGIpkSlTPpDb0A94qyP
3gVdk0IIMjyGIFnXUfxNf9pjDa3RAr9gLcCLILzsqsRpvzbNKm1Rs5GewO47cg+a
cVnqL3JbMLoWME4n9+pU6LsjOmzKmRfpH0JUOQSzNee85mYPdHgFamN00dm3VF1H
+PqTYC6IhfUiAAzth0+LWLdcdom80JyRmfwKlx5M6Wfq2oMEwIW9SX9kjwWLeJsx
IedwN79nfF5GptZQImnMkFMwbgMgOVkekGQjLuFufvnwp3joBQdYx8d6fppb90K/
shPLeodH9UvuSFByY+NcUDjwkmqS0JwpV2e6/xb4yjfr7T3ExPHKs4S0ui6Y8VyW
1sUHAsanVm2o0RkP2GjIHArEvWckwy5wXoJ3iW9t6wtKnPEXdut6wuNLhClCLcRC
jkhJkRABNCostgXEwSh3pgNR627xTUUGz4Hmi8QTvvQucQni0CpnLTvICGc+0UWL
N2T16XL5gmMHgik45BrSsk+4z8VqQiAY3TVtmweSSdPEhSTvwBMiT8iSNY0jwmW9
JoCMnmkeZG0sZMGcZyP4glFkP7zxuGlh2fyTeKiIzjXDh+EVjPpkJNLpmAo4EuLE
FTZGxNmE0eBfZrda/ZpLxNno8Lju1b3xqOqCKtz1XmJUAZ1SCl7Iw5WW2q3m6xYL
9jopuo2/va+yAEUVsWcwFNkf8P8JUepixm++hP6T+CriP9jLWG0SXObyvT+J43KJ
5NWCbETFoRtFkujHyDFCIFAggYCC7rKrc05T6kV+VWaFOKlhpqLmea2gpfimx6g/
O56ngpdbaGrFrXsuI9Q8IDxTmst3rJa1Mo75pZGS6hiDevbIpbpAAXG+PFSH7+lT
WHiGZ17obnS3kDvGpT6yduiIYPwgMqFxqDqhNfxT61f3RJQj7nPW5xpcYEVcyir5
0N/G/5NNlDFa+qc5fhhPPFPZHEYURlJpONACtEbIs5YGFhJwzlErGc5kSqPiVgZ2
AhhMLufZlDniFpCaea/lODodPEi6iHS0n8b987uDAjU3twxp1FPDvMAKvLQrmoEk
bEzP63t+3uLcveZWxww2CnYCm+14mWmp0fr6qiM8if7pOZHfCjIrZOtTrAwI23Vl
miIl2rFLw4Bt/AX2y8ehNfMaxBT8ZqyDb+UUTfksQDUkB/k2ZuX/xYqa+wCQwTUH
obhkRlmK+8VcM1nhcF6skQfakdCzFzNpErMzkcAYhel+92kNh2Kout0pRbVP8k1U
M2d8pcwv6P1hKwkC+iAL8uywAbQXmG32lLwWzs7bMjzyciXfG1oaC+iylpPml6XN
By+W2t+RWpAJYqvoiSLGVO58CyUmLQ2qH5j11Gf1m7/59Xljd7ViW4Mgd/D+62xV
LjJo7ZL2XTXOshxUgQVna5J7EBs6Wjtgq+AXuacKF0raU7RIziu3iYxl+MDhUFAO
8pDMSjhe18UfRD1CNMjhEag5QUMppljRRzbJjZGdeZNfNh+lpI4y1CNT+N4S7ctZ
5+h+15XqwHniqbJWP5X14ZVAl3iNsudh9axKfdhs7hjVTNST9i8+3Y1wihPHozPk
DSUvnfPkg/rDBa2KGTNlfc8WPZgC0NWt6/pbbkl8eeks6+YPK81AxN0TWI/P2ENs
4GO8o9zQYrLyVQjOVFipO8Vp7lJE+aCUeYJyySsJJCCA7ZYDThiKK7p+DzT4nnsR
OzmIIV13YoHlcMKe+6By3cKMFV1OB0mqKhQfQnUpgKQMCewL8f8DnP3uTCtc6HDZ
qP0lsUZFH7p3jZtUd4j8NYeFXjWH8yZ7L5mVj/mCgh5f6vKy0km+a5Wj0ieroCHQ
5EiaNJbm0tWQidKSd3v4cz9WMmBu67MQAbvSWogzhO//PJzJF1Ncjvo3EMjjICLy
9yGYQrSTBcasDJzepviJhzJgIwMx3NP9i2CflpnkYbsR5DO1+WWwwUSZ5gvyzBoh
ZHwuFO9DV8eB8usW2CG1k5Y/yXEGAcsTjra+It5Y33go7R8t6CCY/QBoI7IbJCWV
zrI6XKHbk7DqsQWR2XHf6dLWYYjk8vyIIWzSzZ3M/IwAwJNIqJ+HzLrDgSH7I/vT
ZAvi+9dkzwwP/La3gwp0bJiFj6FRxAvh88YnEAqEiddsYufQ4NeDJjgg3yFIabDD
i2mAezP13CWjvQ5iCLSjkbwScT0X6wZ5T4I17rhWducdT43Uf6cP1KlrwsakU9Bw
SzeVaaqRyiiBiOsYs4KvnWpjegXw1QpYM/tXg3zSoeo5t5KCWslq5iO+u2skg721
m8osEGwaAjXemNJQm3tjdNWoMOERtXHAlyUBYj9lJUBJdYlTLNbk6moL3SmQWI6K
0L7U58JZkgfyIXp6tsDNoukEnbObLrEuONyQxmifQkeKNniOf/w4ZwtVVsRFnQOX
FhERF/RvsQlKexCCdCXllIOz2tdojJJ77/NDIDFVVYBweR+IPMPVo8qjd/nUhY7n
nKor1A8BoscRFLDpOEpTsZD04RcwH0x+d+epcHh7DcvX8C2pB/+lHnB6EOSLrgCB
3Orv5VsiKwq5y6xYOlzZj0VVcp+MWwfxKyD/+ADySLKvdjInw511/WYpA7Zasq5y
MWfN7SQVCLEXmuiFjn1A77WWIyFanhsGaiFzm+pWBw1CHePHhPpeKtU4P10s7OXy
cDRQn9mXICRB4wg6EBPMQPpU8JM4qROBVDK+2gK37415ihSHqwcFkaDrd4+AWia4
4wakL/zILEIN5xex+YUvCrRcALgtEyw1SvL5m+Rps+kGdoJ4icGg6MnTYfeRwqYI
trHR98IqW3oiiSsI2gaqS5GhKUQTphsIJkRFFPT7nNt2apsLw9QuTj7KUxibS+CQ
1ZgitJCyY7TH7dYFLfC2Fcj5VjYBl+zpiAefy7ULURyhl/cMA9bJ4K8jqMI5XJz4
p/BMNDWuveQBYoidOehKyR5emgZHK9Hc/Y3GdK1VvVptzulyf4SQqmF+lG0x7eKn
KV9pNNlUcWWla5Cy7kjR6BdqKmuJmwLWUTbqO4fv0G7bTGkQTcA+nMsBTWHv0P3j
xD2cfOBmJehUNRW9e4ZzR/vQ0aFwgNUTzcgrCBLv+HXu+3GloQcD7iZwig/hbK0J
tVQ96XWPm/Bd5HfUKk7SdWEXGdDMB8qo9v134+fI2jE22jqPwXcPfZpS7JzFWiWd
bdKvdhMRwkhvVTnerXKwcgdXhBGv1U6tBzAUGngOOBz/SbEJY3FQt8TB+0hxQJy6
nGYWfhWREihkrQ2OowPePZ5oEO0Qtn5S/XmWO3BgUFxKnbmeSJinY8t6nnh5tP4r
fe7rDxe8gFJNFwNg25r25FjaC8S6oneotfBSH7yFTXvSZ2wNczReeTcAslfY5tLy
co1uw3g7HGuQ8BrRuXWy4oXbCeYOi6JRjH4aSXTFRtQ4VcmYRS47YfgDkPAgZJBX
rgas4wcyazHXjeW0Qmj+32gzox78EmEPdUoVOUebEzeRBVDs0rYsBTOdzqUNC0/O
htnMf9PM1+cQtofMU1fbpOQCLlFP7cAwGzYyyvfTHICa+GCw+Lk8ygRUfMqqsrhG
eFkwmkGq16Mm8fbBs7TpDT4Td2ATlRiHmmFBQ1xng3Coy/QcnXYx4qeFngTx3/BM
By1U433GmSpvTpy6km1gEybDG0cwkH5WzV1TAMEZJvbA+pEIBi8h2CcVHIKdGLhC
oFdeNpMLvd9mtKA6u7DWhUAX9PYdYWddkdHWXYTmjtA+1G212vummAGY+FjTik/5
Y8bQx/YWIQEOVzzcmm++BFtGXgp4l2Zz72F4rnLZ9UEaF78T3vvSTOrKvPFWDOjK
Kb6Ktq7hpqyBEOENiHmBld2794K60wGraCJGWJv7qKviWEcMcXQ02H2nHIDfEBRK
oNmxhyBdsSoCFppo5u+DM52xF8JXMrvZgW/iJz+3G5aMFOpuPYKCWp6Iawn2Wv6O
QjLWbaaG+x08TFUlFlHjAeOEdKT/DMsLMcMLiRIg7scS5SN0msfEmh6+rFeGv3I5
Z4BOsKunbIM2Znuvp7PpNmzruXqkPWH5o6OMuZ+7RsvPcAPQAaGM2JR5Mw1i04cJ
ZyZCXMtZa7l4DCK6k6c7yXFu4fWte716jd6QmKRmi51E8scK6HkZnVwRaEWQrq50
xrzfEpSajcDFuLcb7DAcBKH9pvNJgBjd5+iRbjk3DOclWETrqXh9KDHEP11kGR6f
g5FU+4nJt79PLIk+DCx/vwveiSlC5DyCZ0SvTQF2bg08cvSeZ4LxzWJ2SBg5PDqf
Aqr7+axjMs7XWrI8Y39aSQ5fGMzgy7R4ZoTzdBxjIExvwKbpLPX1h/tNf05XXzie
sfXpVM7TqfvLUH9lzeZGH20zvFGjy0hLkfcwnPXizrVFKOzL8CvbJ58yfU7234Le
Zfcct1/wEV5hXNzTcncs3o1wq58jtiBXCx4peAmC/1yuCWlU6F9OtugMxoZty5+X
yVQsliY29mQB9Bd3Po0aEjZdD05phAOWtuFatE2jhRrO3XsxQlMvs/sKoYjjw1lq
2ejSN/11iEBrS1L3Al3jvMiMUHoItSpU5W63axeZw+Z4Gb6GJfJbbsrm1Ozj0gAA
wdIlQwc2uuxr6oSa9GEZI/MwTzcatgbkZmLKIs9DT/1FQCnJB5lYudUqCSoFCqey
XSKGkWXgP8UDMuZ5XrqRqD0WziWLc2XbsfVnZhoT92lGnCNaaaLTZvPdHwHh7CF0
EhlI2JnFBR3pLWxjmEG8zy2FpXp7tGkHIMEJDbpF5l4bQzqkP/4VpCZAHD91Xjan
LWzk7ncGI32VZXlTLMCl0ebxJFvV7XCqxgnGgLwcDdE3vTYW9nE7hlRJUIZ+59yw
HLAfSDwMteKNyDoHpAOySrUW+AOWtTfX+Sr6urvG3jpuZ4h44a+oK276gslEcjmp
XXJpajA/p6xj15qT3YwWXpx45/K0hO9n2+MT+3bqvay06Ksk70mfqV8+IUP5cEgk
W7ikuV4CffksLXCveYtT7jdVsxnCgLgS5ul6si+uGcBQ82AtGNaNFnFO6AYrHrNx
KbnjlFpvzuzxBQvgfQqn+jJbqIf+XVbHfO7naWOYVfDwZ2z2hG+WuokQcXgH3OdP
uvPRI6g9zNgrDpFLNt5z3qhKhLq0sGfNyHSqmNLX2Ld0rr1nSIKfqrpOePBsvG3i
D+VIttGPXsgYrC5GuBYxl50IjI1+J9xGk+fWIw1CzDLkFQZbATgKJXdFSA+4wbiQ
2PowoH4BkXZtq6HV+jron6ca5y0tHrnuJYyyA4mtJ43Nw7fSiPHIihp3ws/YRbux
hUKthwBPoy9GDSmATe9eRRCMWKIcdJQfhE4OL2UGed2DgX1fKyhuyvTQuogCo9QC
Wsqa0WAybDhOE1adtT1ZXTd0rnR3UyYcAVUse4pe+21gG6A2bF5RZ1/cYgtQfndd
ETIuKJ4iPX1g8qLTFJ7V8Dst3nQ8kRDfG/S0biY/jrHibqBOO5PSmcNp1bkC0KHI
UMz/Pg0enNG3nmGfA5vMyOdrrzWCp3jFUH9XirhlnByRPL/6EUuH7vo3Robd1Pc2
ILUci7ZnZU9oTtp6LQjiYOkuK6nxRqcYySwkv419Za3NpWYXoP4luJ2fMM3mSpEG
ksDtMQvX3+tCP9YyoibRaZAAK8fSGK1WQemd4WuX+ALDJ6DePiaPhGZclPttjHYj
QMvX4yvav7CShjMg9uOJ4kF/5huyY2oC5NcQnL9kcp64hpgHKdpSUNiuXxVnCJKB
wPNJITIaPPGDRCQA/XLoydRN0icqrVymcaMsPQy2b+CAX+1lmRS9LXGPU8T7jXAm
EQg9jlnJPKufgI0RTWK2ErECLQNn3CzlrmwStU0deiaA1zNu/SFJfaXxF30F0GLC
KzBjIiPbn2AcAiv6e7QL+LIZsrdeZ+UP9xkaBFYFS/d+HGL3OEKTuo38WoNhi3CJ
TIEEWGJsbFfU2VF0Q07AB1LNkEpeBKWeitjyVSUoKuVewna2M1THeFNqiGgX9odB
sV/zXSgZ8mM0p+3cXPmHrE329vkmmH8/QMYarq0M1BTidOU6oqV7dNn33Q/7pyN2
xSL69pbLZLNJYiEEteAPjCqLl7tUKnvXcvE0fakUXzw9b8MPWVeiAT92vrZyTFTI
YO2WB9d/lZfsxArUtN2q5UYgR+L+xBbuUKTxYEvPIN0n4HSlimq+XSozY1qksThx
B7uO5O9w0b/Z2ecsTi4XEihABfLH9baOkvlXnL4Pitey4qL6b+lANf0Mc9UrtwZ/
ST09OA2SaQNcVnhvGNxAGt3WsYmIsghxl3RzP5PTFytIX3vR78RVOchzXDnSxHuO
ZweLsxOFAQTzxENt0mAym1sT8Gz+Ag3bMOu/5I702rI1dLWAEnLfukHXx4JhgTz3
ERGMpcqeQDCz7F9GHsM/3T4XLPhPPA9YkpP4Sd0vGnD9E2VV7BOvF0+gQiGMCbXu
QliPYKb1doMMkx4ZHjL2QoktIn6J8Qy651LA1/UxS/42ysf+QsZcZdVgI+c4+xpU
uXS5N4mvoqdGdxiXJRVGGeOLsu93qGbj/1H57YSiLndd1v7Q8HN+8jA5CuPQpMPT
xlEbhI4M+htEKgT34S9jQjYloAVnrZNcpyIZywj3/N/jdtQ8DIbRM6thfr5cO4+v
dHBXKil/DXm6aW/G3sFgWkSETpfjXEA2t3gO09zTFnwBbivUtH7917Ecy64Xpfaq
R4ujBAyoKoyrtJMRVyio5IUNVBgGO83xPUXjBzaBcH1CXSFmsOvMTCSxRLdveiHl
3ypN461tLw1tqYfXa5F6PhYaPPm9Eu9MGy2hAbxL2yDEquGaMh3n0+z0IUt9QSuZ
G6K6S5tBPy68SKc0ypDTsuQa4x1EnCbQs2s5RhNSeYWygAwlUAi4B6Uhz/Yl5s2B
qWJcWvR60U1Naquij5x1S70R0DKVytthVU/0jg6Q/kGhx4mrPX391M2XomE6+MCM
UcDd2u0/jSBm7eQ7O1BYaOYEjI706NlsHtUmahFu8Kq3ChN4sh5CoBLN+TtiuxeA
4BhAtVKLFLw535BH57V3qWvORoNA/3VcMVKZKpL/9rEK60W7+3G7SxgIE5UrQbXc
Ujs+SFOyYPrN0PYlcmd7PP5qH0mscm5PVYtydVrmkpIGR0uv97yG1dO/4MQNGQKS
yfgbJvRQcHgFopRSBAXdTK3Qs7hy8F4eT9PMqpGgahrHVnhMq6wHMUG3293z9tbB
INws2734YfghrrFUHl6+ZRmciKYIRFMPKr4mBba+6aPE34wynHIAg+5bmRZq5EJV
wlzq0Xw9GQQlpIYCVv3avujuvQlnLAAsWg0B8zcZumekYrqu/GeFHLD5MPU55+1c
F+bSa0gYdGjhjddFScHaeAkfB19Ua6m6zQsRmQPkWTjro7rhB2Y325kKAh3QluPO
/Ljl/2Acxyq5vR/DPSU3NJqmUEIrbMNrETDM1zP6/sKKwxpgtMGjdMDSSWPnpI5C
jo2IjXHhZ+fie0ykCk0L5+85To3ieBNtw3IaN98rBRs0dHxc7cPi2rA515h/vPZ0
F6vrC9AfNArvSUw6hHLCguBSo3PFHXTqU20Gt8N7fu7LLTZXFOkn7nr5UxqSyDDu
i0jwTFpSBVdkkvybuNYHlIsc2fMC2Mwp7QuAEMV+yAr3y00tgGJCLDOGgawQxrol
WLs2oSBXqDbdsg33ojCouuEJ3nRF+1VBK5WOueDyHesNkkT2JXYwfnHTm4+Y7NqG
YBS2OUoQTBzDcoF1Ki7sRqcVfaUdNCJIM0T9OuWXuAmKiOzvkkLp8jjCLzd/P5kX
KuiFgxTcWlLE5pHQW6b2vfPNHC/c64GK1mHFL5zzVzqIM0Q2Uvxo5WB/1ieX0bgp
7jus5/eq/u6daI0QAh9cX0dQZhA5Wgx7s08udWugPu8pxpSyJLCNgwWnpq/QV/Kz
QiEpG7ghSD7+gITY0SZvfO16CDM71hwufK0jhreN+wKrKvjEI6RN1E4UWwMCmUV6
MOgLGsRmtwvoVwilh99mDn9uWrrYvPD/3lbFADsIPmemtXoG5eyXL1WGgtMEjgBb
902dUxz6pDuBVRKAtod4YjWCuLJ4v7OOiT1sd6dTELcuyaTQlS+NHxWgmTKdS0EM
rVuw+BM5kjy5/4RGV9TZiZnCc2AbH0PVwyz8nmeyX/0TwasHT2/IOFogiSX9zNuJ
K8/VQUmSAdg5qcaBWOqUT70IzuZYpmWcFBYZ+A+ddMKri/Sgm1NmIBVCmjUot3lq
J1Y7tWh+zkVCOhXQZfJkTAthI3bhJ/At9BtGsyXf0e/htYuLZaWF0exkAd3krDQz
haq7YDh2XD1sJYdIy3/ikHocbgx88t6Csui4tkW7uryAAY6v7SdNCMMaE0oYC21H
Y2gOMgRUdKIr1GOEz7C0KEdFsgKFTlKDQ8zp3bGjb5XGkbHUdaD2Tensrx8rlUnn
LpT/dqz7k2Gm0Ukv9XOHKgo/jVVply8tdfgUT57va7pGZbCPnx4bxeEdQb/b2LQ/
omgDoie1bHdR7oGaNXLojnhA94wvOmOuxTqcYuB8nLEzbl7w5TI3GTOyGRBRSSe3
DCeIRHYevpLJmybwA/gVfwd9CmPRBCqe7s+p8ZvJ+oxTaN6KMqDqLPE+Q6H7ICnF
vOahcuunUnNPD3QeGcfGbUsyNCEhQ8kvL4muhYfWp33MJgktQwv9Of/iXb2uVvbU
u1Q4ZX6diTRG/hSuqQ4MKnyadZpBDjdTrAm0d7bnBUFtHClqBVQTaUUdjN6MvCI/
YYKpDSTgIZBXWwipKgYIUd23QFgvHVmOdNXQV3rn+GJhIuX4jul4HqmHp0HHEggw
5ExtuuZ1l18FhLIgcmjWXx1fQ7E5ex/ViBE5S9UwCuAlm0QHhlWUJxHWNtGURLYD
frCyWkyyNOhodeFWqxEbuYm10kNMp2+GQLaI/Dm+HPSlVRfyGXkyw+tn2OpSnu5m
PfwKsSkaEymWDDCQDB9EUZSyTkn8Fco/Xflj9Sj1m49Y+MdacjJ1L8sutSrhsGLE
Rk2BNuv6lZLkQ2CbQbw3uNwbzR0ZDmmhQ5db0LOqf2q1ymkIwEGZut6YZ9KhEb21
YQNuEfUZby8VXv1EqxRInQLmyzn7uNDmtw4xa1HVoZ0GkPujPAdb8OSbDn0U//e/
KpEymj9H+SdX1csVwWpR3cIn16uf0V3RCSLfUXttlj3jajebUcFqKY6MSvyjiZHg
X/VWi68RcffI7wjbJWDkZuMHdl7tcVV04m9Uu9bMljkI5QYRekKYi9Ah7qCxxHT2
U+uqX53G1dK6H6SCIdRvi3IBqso9eVCFnf4pYbzcBYv7YtFQY0rmIY8vXZZCD6l3
Vyzo5cw/rg6p5CcR4xXFnFcarfKfKm/H2VDsmmo2Dx0ib4EsjVF/R6tboIaBRPsf
i9YtNkuM6YqM6PwPtQKPWV8F4DAK2UNc9RbcIRkIxGXti6K1552i4v9Sp4Sbo2iO
Lqk2aipiU3QStjEk3nfr4AbI00pihBxsSC99BUuTPSBD0ugEbFP8OvDsMsZ0ALHx
9R09V0tpFhk0ALnU95YWkYHBCPcHio0ig/yju03V31298vH91H4EoyP0nmP/H7Du
Ui0vhD7SJS3Xjzt5oDP1z8AgVuyy7f5woNiBEVvjXffVw8JcUkcTQWcAuj6dCH/K
dTlcrvUnUGi2UoXxh0yqHToDK/ZEn0KomVkmdYuSkMAjfrRq5npkF5R9Fao8EYdB
uiDxSOmbT9O3Mn4gHkrJbRSR1NCZ3xCOhYuO9lZqQAwGy264q/FFC9DJMxL0yzJd
qCvnUHZS4wM/QPrtkM5fG3sknWthbY5DFkK2+r9z/xBx9hEu/coFQ+7oN6lof4oa
3VW2JpAJv6IEcxBExmIa3wIbEDEOrUVwwPepdrtqFzFhHZ/ezNZvoyekl7VZ05pS
Tk6Zilv1FPTrsInMRRGZSXmrX4T0nBXPO4BLdMlwfxf6NnDwTvmICSUhrN9Nagcz
2To/xj7ZJdnPQinVbf5jypCQgse8juVuL8CkDToL8pxwzMGv//9q6yKtjCVQJlV+
MKfsOfXwgOF5UY37102WFD7FviWRLloSEDYTcCYAMIJewt2HTUg+/tZ/dxvWX7Vw
kmHoOtXpMvfApxN2CCPORKQxrFLrhg09bbKOJZgETj3/XBA0RM6AGYwjWptGo1nQ
oAmCTIQqn5OFkOFh3UhBc39O1GQz8U2/D30z7Qk9AVGihIsv5Xyxoq+MR4Dua/Ur
HE9LcqWTTUtPtFbR0PyOpBoF9w2zDnxeSmuRIH2EnZDOAHH+wZImfauGogZ0Kdn0
PawzdgyaJKww1MfDGVNghdXjR0iv9nxYn5PvBm8GrSUp7mdxC4/jcJC/c56+NNA9
D1ejWXtpS7hlczWzoHu37YmLJ3c9eAisnQ+St2cxUnbTycgzuPvbulDpMYhY1fBj
DIxUT2XvNKxNIApUH9fTG1uHQp6uD1Lf1VXomqYAAe/pkXYjGDKQzDD0n2a5LfdY
hcx+sSYXqdStZm5e7Z8yHagDzxWlI5QyZFk6+eyWW/imPFBSWfvcGzGz5l4F2tab
pZGoW+wS5D+lTUZkvloZWGmGk5Czw9Vl6aMu1kGdgazHboMOWiQ0Rl6NQbqMH8DT
5O2rx0CX1hWaPdFnNjn2vYztXW3AVPrHXiCqEKcT792QyaD8Buf5B2i9cEIWbvlT
NMcSp08QFfTYNb4k1QOUkLVXgA9rZOYnrSrwd7yU7gAdC23eDOiN4G3uCtIIONk8
31QQGJV+QjR82X80T7l2jv9xzMGC6kO+iQ4EuoxnjlZVc9E2aOzxl6i6LbpYiNAQ
yRmpbVkPv5AxeDWdA5x5MPtadGk2G6rAxyp5ttXAxW118uYJg4jYM3lpwwQ0mgO7
FQ7PFwKTBTb66YrsNk6x21giKA5nTqDEDUECCDhC2ptAdYUCNeg/WsbdW0Bq5IFb
K0NkAT0eHewBi0FTJ0YKluoHMy5myE485ik/Df+on0K2fkKb07JPnL0TWFNoqnBF
8PVJvsDqiqn1Ckql7mpDQswTZdCw1v+zk+MbqIOjQPcCrdg4iOJUKGA+2q3bMa1A
Rt5Qn53F/vaBHB1giL4UCePr9+e/c4i1qY66bvB5XYphDrmWLqyzVBIQ/9K7eKSr
r/3mOhQ/xJ+nMMUfAZgyltDhH5R5rKGLpbzoLxhN1vK1akUKBQKdHRk/4JlBF8ws
tQPs8B3LVH1Fh+h3PetgEI1+WXWJ1EXuCpLLZLd9WELEwQVDyM8Jl8hrywzLVc36
v/HLptz4yzteDLrPPiQkemPgY5kpn7edmssQrNa3ravyTB2joYuQa2qYuSXaZzqG
KwZ5tJQo2meNeBqaZU3fVABH/4UIoKasxxoyAqYa8Dddj/mDf0cEwZzXM4eSpmAU
u7oSPdzqTKb+wgzYYW321Pj+937otNtey6QnwMfRSn77Lz8AcVs72eCbEmbHN2Lo
uYRCXCQblZgzyGNAzmxP2i2YCnSoJeM7A5yOdJYtWVLdMDFuE/Hk20Gh+B2qZMs6
0SJGTi88Fz8THAYL1XF1BghMqUFk4aJjGMOstI0KWutS1BdHFujj0/9TTSXIP+Qy
3E0W7XKGfkXuPKOzMaXHHFV8i5OuziUzqsw1UWpeTSChkQhcmtpK3HsKgwQZvnv8
mz/l2p4N2BhAjN9/fAMvFeWqD+BzH10GgnDU48EigE3ck4aV62vCgV5VeCDm3+No
0XWOKuW9XGrBSjjKqgepYDcvjKE9lrkrlluvOt+F7JJBYEMUbqBdbovp/HBqh/jN
ljmCW/VWIlB2Om/KznBDHCkn7X5Q4cxv0zhJmKrk3nwUJfid8ylx+xs/XDsjIA3V
hDGmtnjL/k+xFC3Zkb2if+JfK1QTLhlBaeDERpheZ/BQ2P0aQMehUNhlYK9acQta
ygQn0qbQQhyd1BbhvBfDRfHW8md89TBENOq8z9Sr1ZAokTkVnNCwgpPofmEJLR2x
CX2HdomrWQ/0aUZIp8s7F9QebgQoFSvd2QCczYFF44lK/GgKH5UNGtJbV8khkb1S
sH4yXcGncuaCS2usJrihbqt51HhL+swz+aS9cGoU2Mx2dGD9/mJKxHq48eH9NErH
y0n56ce1oBsf878rnGttnPWoyBeeOwHdnl81WquCja+GmFkfgs2+r67uvWAnyJC9
maGw2AwL8+p95HJt82fx0oTAfoFPKyl+r1qYhqk5RRMM3pBp+HaIeSMrV/wSnvaN
UD5JaWlmbAh+Wn5s4r3Oez6mGAx6AzQ4CCkhBH3JmiIHPgHFQEYCeXxnxISfjsDw
rzLrT1ER6UjtDkYVgtcqrvZKCIBHg0tYt4LkWYIejfj6PvPOD0MzvdxIGSQjSQ9Z
1ptTHIpTZdx9187xrAJK9gs4tQDOwNH+i4Ko9dE7vFgLloB2jb0DzcIq4mP7KESH
HHnVhHo5eD73AYJ9yN4xPHsAwQwoUuJMEuooSNcUfJZYr6lqL7kpWBInhV+l8gi8
gMFpUiZ28sTjYzxZAGKBQL4Y4/Hdz2U1Tgv5AxLyKCX7/N/jTDUtt2znzuCKA9pn
AvAevfJgrukzUKrfO8EzLVPptAXOwqcdg1eA6jBV0FNf56X2mQfTVCsZgOLdZ7WD
Imgo4ITf9dW29kJaBoOxy5CxOvMQbU7S/LHdbTBuzJbg0FD1LL1FPYuTgi+YD7Qb
in4pE5GnlRqQV3WOii40KweqEiiZMCShfkrswaPwauSkmPncSg7lob/+JAuDEqsd
3QcP5jhXODezcMhIvdQn1pDO8SRh874pfuVGjcGk6v4rHYbtpKDh9Q1q4peZbCe+
uM5xDCvqv/gcliEcOulRGz26NTgzm6BkqyxHIBHQbHXypXP827JYpUaXXlAFZ0ax
qYaKX+dbMKdr7BLSspBOL2YXXzKx/KJ9Q14jKyY4YBJI5yCVKARHdJWX/JSQI9+I
zl92mXUW5G98hyznrHgj1FpN7IRldWXHShb9BJ4fBs4MRYTbGb9pTJDLZo0RYIDl
jVR3Xjv4pp8QWUUf8VrwA//16v8EHTcPYeU7EUS5KdmDTtHrueD/RmcAaeB5nF1m
OYVVD4yonrew+XR0S9s5jEGhEq9lFzHTuQLCtGwsDNFA6fwmu9QkAZ5AJbjP5IiE
mcrN2FvvhvapZPSupdxSoAArFQeFzwkdi+9df49IYZrM4rLoWUdudYgqy6K+O2du
Vj+cZfUAaw2CY1at6Qgw4lnHexBAUUCuW8G2mxVaYiIpc63A20/Cjd/aygWoXW5s
G8JUtft349vzeCeOs6peP0Vtl98eVzdN+jrRnkFngfgB59nICIL38tHOjWWFSqhi
TalnXm5JsrOS51ohnY8svWjvUsw7OKwVZCy/C3ONM1DnRFFAILluEw2aNGMGpHtc
DjyGm9JS5sec7KspaZ5dSaT+fmm3wObIqiZyXUo04QuAWHGAwpYi8wdZS5yI9lVJ
7Ztktj0C/TjWzm8RRtn1+rxaGZNMGBPSRYvKH3NQifVpbKSW3U0XaYJdSEvuNNDc
uQMy5M1UcHQjujomVBjCImX6rwRhFntZObe8Ohpf/MUlCK/PRsRhDmMZ92X8buyI
w+iFCbd4v//GTyDPvN8YJvqzJ7TXo0z247DyYpdT2AuOSARgBQW/dHz0d/m5s1kF
jXe0lbkND6AvdzmmT5R22cnXIBQEeNJy8n2MMHCTW+1E1lXCXE+wi32dERL8hcMJ
L0FCri8DbRPmwUeYi04IJI+JqjBvLHHS5+5nM9iu93RE54U0fi+TvgvOWYLjVdyI
bLtE/n7Pj+9Y77JCKOvab3rZarYQNqVaYRiDyBrm2PK1txj07GNmWxCS8KH9WgLf
3CZEMUVyVWuoNeNDRgl2NpQKBLd5HNQeOrbos0tdLzEEeQjNbUSKR8YiIcSHncyk
lIFlDmxau69ANjflzVGtJfwLw9O+cpAQ6O6oO8J4i85pYZk7NClu3AoDM/z/sPPg
36N4rzWYsA7dRBo96akULIq3VSIxdcyTnHTydSa5DBgubVcj2exTlUh/TWANAmgM
gl81MzUTK76mXhf/l3ICLA4kNhNqdFetR/tLH+LAl2BHalslsYFK8zGZ8iCbpwQp
sUKSLOxB+UQhQIKBVs01/ObjvG6NyPvKWInkM4/jsHO9jCMwYtE4+C8K7J6GByZo
F7bYg986INC9M+zOCIA4QuEMvJEAacm1hK5CnlHX+f7MBpugkoxiRQahexf4PaqI
NjJ5Idow6TUtWwfHpiuaBXL3plbJfDbG6Ih/gItLcshxQcCZEqUKJFoiMY0F0+1b
XP64h3nVmrCxxjzo1yUf8/MBg4lUNs5++38/xuP9C2X5a4KLio3li4AssWsTsrT2
GjJO8htkufGiPDaMkyQ2mz590FF0Ntp9u4v020+RTB5fxDsc1BnOvMJYep5znh//
AGs5TUTn+tzQtuKUZxyxKuZTdsDOa7LljrfLjnSJNh49L9OUyDzxBKO/GWhrK61g
tYAPXrkvrvTQ1eKLHlljM2+d4ZPPkCi06D3QLaL+L00ajhs0F4wmvRPg4nBQMf0Q
TcpzFlY+XfhrlnZ8Xu37xfx5bpaVJ4ePvxICCIKTuOAbBDf3sy8myeESBYu+Z2do
DCs66SscOyw2YFUW5YhgaBwzYuXjW9j03M1CL8zyJiJ4+rR1IZ+NCLvR01UbOxBs
4PKH1Rbxnmgq1FXhLNahv4xc+Xn91Pz2aSAXik2cqDiAfRLI1FXyuh7g7Q19NaF2
oeWxoNxnqUYgQBqTiUtxRHn54yVbe9V9jfUPpbB2wt91Fhjkm06RaBnka99+nlUW
wHhs9PUWcYlKgdAn6BeRuiwt6p7We08BeV/KjhNmV5+ocSkNEdUWd6AHevBtLrFO
Jm3iR6a6hXNihuc9S2yOr9xqU84XuJvL0Sk1ZlFV++Q+flTDgJDKxplR84eiCOmP
WxoqgH307R1lmCLzQb2ANi8xho7h7cLFb+IZPJbFCFCgAjRU6vzFTXrevHZeqflt
/SM7qiYVTUrzWAZfF3EPSzL5OBjos54JeCAYG9prtoc0xdrsLEYIprtJ2WtSBQhE
DdxQCj29Erm+XKqtOU4fItKKHa+rZ1o8VT0cbuN4SK9RSkDwMgLmaWKcfUw+o5Ky
qqNDBq5Gu+vVPK9mOr/eI2GvQmgbqazL/hDp7mJlH0KpjkPeWsaRRdueATWeRzKf
6ci74aPCZT5yjcShgVi3L45J7a7y8OuhrigbKrTrvrnczEKtnoZJIdLbGVKScClZ
6Rh0A3+vEcoqRMR+tsuNxRF1ayoE1Wxbs+2cO7ING48k75gkWCWwWJOyP62Zjnbo
Hi7ym6rd7y0h9nDGPjr1eV653YpycSb9jLoMIM+n3CKy4olDBlleMm5hLCnGGIVJ
TuyXJqXdY7029zxQXRmsjABY46YX8jDVIbMcQa0dv1alRmUqZuB5A6AzYcICoIlC
wV9DFDoW+yWhS6XRU+EwaSYHN7WHMsoVhXF72zs5L0LAah7LxS8vDzhqOMvV2Kk5
mUrMO/KyJGhWl7hQNJdsqZQwm1naEZY3UtaRBLB7tMxvuVbYeHe1JgYWOelu5MC6
3hCO6FcpAQaimBQTO8Q6Z7DLyXHHxwtuvRX9JvAItajVJWm7RmYX6xoSNS+xtI1S
yM4xfUrSe90ocOr8AgsxRmgU/okMoTHnDugu9f9FcHQpj59rGbt0xjhOKdSW7254
a8pycCLQepC2hDOhxMUJiEJ/kCuzkIRzro598Spg3kKbQU0qwUuv4P0AroZGu37d
YplujI/FvbBIK7FbGM51SLk/usF+c5ZfBStkKwHcaLcAGH+mByq2ewV78iOh83HT
33CsAxMKFGsI6f/Yy0Lo8xiIwOlhUUSQqvlROFkLFqsn3odIRRB6KMnVL8DJE5oE
eY+2nVKdUe298IF4EmzLFxBO+wmYTMUCJdHilP2LKbsRbne8F+f7LHoXaKcezims
K8nH/d7W7YKEEbQu7iPz+poqcSpNoJvPUiXKXGJPsRgod86uMRiGoCXkfyMa0+5e
aoRM+t4f1oq4vvgEw8mnXld3HNmxDTvemS23iG+hmdRaFs49KDwqP8zerXWwb/m+
WCjuHIk3ga3HMKsE9aI8pQrrQd7xaE/UVNHxEcmGgWJE2rJCO/mEif5zYsOD/aRn
E2YPeJEGhzWQTGo6WBXbeMWkU+LyGyILeUoCFvrwkPXosRPxKRLhxpc7YhFjwYk8
2xY+RodMaSDV3/fb6rZrIIAziPQYVJhyecXnk5DT8d61nEqyTmBaRfA/nL+HowrA
FLZzC27QoY0vO+aRA+x2eJSjRykv5vc6L70FH3Thj4DiU1SlNC/ilLnVP/6vixCK
Ok+L8oRFiaVGF9w+aFIkmiujghEKnOlijejpuX3znfA5C/EvheK6TQoVFEHG+hJJ
DN0DiryPyWjPH69z6DJqaRSuTx4E55tf13614XbTEAnkxmN/M8Km/i7rrQw0tLET
eck9BJL40M1+aYjtX/lLE9DWPnMow1mHnldSeHyi0DDWhDgxVBrYHT3Fh5bfCR9s
v9L/5EbJN8sAjeXnMq/Qz+Q2I+gMqu2rZuPtHrzAB3tSANqttXs6vrwavnD5uDTv
hVdsFnv5FAy98knoNtRRG8pVaS4sqSGGwJ0uCZO/mddFADasV0S87RgVnhwFapNM
tomQBDn3vTN5O13d4DHSEu0fhK5rQOeigBu8qHPQHG0oOGwQ2pQc938k2u3XCrIM
HFQYgbsL8E1Yi+vRRdLrqpt7V3B6M7Hw2Sq/jp6Ji+GesSKRA1c0toVLTLvryIFO
0c4t1FirPWLSqPVYYSRZ+2wL/7/XHXYw0mFlFpzIebqTdu46frd+Jg/G5VIK62Oa
uLNCONZfCQtM+zEPtzqTA9ndIA8H4GaaLC7MdEIBhb17aOstndj37yea9kD9Lfzk
FnDhnV0XQZRRbRcdIJ+YKFGIoK/akpaNbiNeMDCqNrAZCPZk4fPEagHnGdHxcSEE
AG/EpwzquJ/RrLIyI9ziux3w63UbhfJPw6JJbxBJ5nv5sjRdeZyE2Xnenj3abpzI
9YM7WumH/8kfUlfxQ38McvqTg4ulM961NYRhF5WZJdMJfJvg3VEUKe7rCKKNe5XN
R/uqZIpt3Gl+PP6JGOVULZIYg6E3hsbsYZ3Uqtrw4uZHiE14WPqSAycSY4TMoxKM
l8tammHaKDtr2eDPGCfgyRVaW0URiPjb8MI/KLZQwRr3LxlO8yR27uGiKmM/D7gX
jUEkIlO55NN0xTBfPeTviXIF9Xyi2XyEonhHmcdixe8qJIOby0AhXl6HBgi9aLL2
13UUJKnHLO5eGOa1V+VoZL5p2cyB5S9SdTaDqDwl8oALQvccyF6R6Jn6J+rYnTLY
jU7eIJ99tT5cbn7yjTy4pTwtKiFAcHcmxZRcV6+i0OG6MUfoDRGX4XX38x3vke0N
hhkrtIBEvRceVHIEbFTTTDFfpz4NYmLeUNoystA7TRgFaYYJ8j6dcP5GfASPej7a
wQQIPzFTNh64czjtED2UT6bY9JU8On/TlPFIJ6b9u/Pj6fjFGsoRjkK2voUutVWW
+lDwM1+L/bEh24uSlt0bIZXv3FpB6v0h9tnbAb5RREFNb8mmyIUyplvwLPiu5Tk7
EpvgcGR8EsCEqWteoFH5ZADhieaklqU+mvgoeVMxEjh2q/1d8c/e6DVCuuB4raV+
6O8pam9eprnzUtBIb/STbiTMJg+OckvkRbFBmYB/wkv/nAkABpjHYNVctl+7Wgg7
OBmLB6+raz3SLhhqaAHiz+fYhi/0kiUi3iwsVbpYsXMR0EN69m8Cb4x0kGufKjOE
7ca1uWwakHp54bacHuQyGV3zP432ayVs31KdYrNYyCmU0WghW/ZecPIAlkBdfKX8
QoN4GK1MHZ57z9d28Z9HSXQA5+MuajQKC/+RtwaFMEN+kviKTAnwrwwVrpwd+WQm
St6IiECjdmeNXD64NKAFD1QktUlDB6KdvpQx7+EgnwnnkDN+rcFMxMHLAl2WK7m4
vxqh8Y2xa1xw25T4oPpJr4bJnHjOHMK0zvload+neAWv0tQXOyaB5McV9v5IHL9K
IhILMtWFZlibHeiC+JcJ5a/pSNbgY1MrQnrAwGZ55NwteWiyVLdXeT07nMayUa0N
iaUmxoclh12ljNnWoVKqaRVJMBdvoFuWPdbslMX37QKrHzx2/f4SM26ScimzkYq0
H3UEiykpl0ewC66fA38cdR8nytT11YrZBgX8tDfro6xdl6IT5UO3sVh6/3aqmJO6
mbQwmiNwJfg+CeCfmTIUlBCYHot92IReA+0UCKOtGpNG/qVRaIoBMC5gZf9S8zg5
psnVEpuXv7hYy6TzLh79iEYpdXb4sQ04LYt/xPIyI+Ut0Gap3ejnJmcgH3OtZxId
wHArikzGXr9M22v5HUXj3ruONKPnCdE6ZIP/3HQHJQI1cTEfl8ideLfZ3EOQLfeH
AjVcxCHWvDPJp9eorSHTUP4cWWzSGSnkFatFo6/qG+6GJdqUH7Yj7XhsXl5aeitK
445D3bqilPFxy3gti+YiZvzVhYx1YoC9PAB0RBnAXjYz8BvbedMerQQzmiu1SZhu
3acS+WNxW40Pau7iAJNMmzIpD4aaDh3l2HYCjXsvINuMioJJPhxGOnuz+NC6+I7c
L5QxISxN+LWaH8cQce4RoErQp5MRKITukc8VmsuuLmCvJeXaB8VhQdVC/XgCmk8k
OzHVAOtBE14vY6L41lYrVsy9J1o+mJATHWFKiFMudTfdJBdYLvbCkscQnZ8SxXSa
b9texNnrAKmXW/7MjKxJYpwIvD9uFRRe6E+bjog5bFmCAvxptJpZqOz8KvDUsYFd
aEvsmebElLsMRU4GUkBjs1AIIHRWKC1B8HfgRToB2xGo+xznvGYrLUVND/cWy/2J
UE7e/zZtLhqfYcEasptgqhHTvgoW9hF0AUokcarG2rmOq1Cftru0CT3kMreXka2e
sbVqzcNFw7bqJr69KiXLnAxvNTr/uvlwTiMAUvFiMBymBVozyW0f5z0KaI85X9C2
bx1Cv+0Nq1obAiEqAe4cLOgoS6kpuB6KNnaqFyFyBl3OkUOxVrnaplR9ucns8Gvj
O16cz+WhS2WrIGK8Z8ApaLYp0KPZgxdhvExtVxwNjVl8g4WV8EsvpzIKQYNP+fIf
DjKhWY22DyYI97qxWe72rpBSYR0KjRrsB0RiYGGWO32LqxhGBAr1CRNOAwddFpVV
7bugUFP49Jv1CgW0QnH/J6S0sRAkTGuuvHddhBdbxiKJz7wDFK5hiu8DDR2h7KQ4
Q01vHbf71t6R86MYRT+TQ7r0F1OJKjZwz9zPZhsYkAeTkM7LfaZjfvdUtcp+TxdU
M5VX3F6KM7YW5WCREW0eeL9CzCxzxMe9CcalckPgHF6+W/rvfcKCP3j+ghC9txMO
Evr9RAy3MmQWRY3xSHdAg8dUUewTmVCZ/K1NNzrBCBQrkLM/4pNv7GEiO2jwJIwG
oRXxr/ln9HByZGXAqxzsRmGw5AcPUWp6mZfU4zFDej5Nza+TYrl1ygxlo455Z+ai
mkj4zUwYyUVTkbnogVkM2HbNEJHssYBuiC0laCmd06okjpIacK08oJqo79TgVnXp
3gzuC8iMcMQSO7JjlYzgxOXPeZAUl6VkwQ/7FFwKgJC8ZQbWr22z5Z3MPU0rkEmI
05GkabaJJef/pAKNzkjboxEQspEpYydcf9TqVdj0gVGR7VDUgKC4kOFRCHVJP2jS
si+JqDtj5u2KnjdB1PT7FtwDQ3hGBMZVoeVeTC9AYMdLplmuWslOGaH0OWCZ4Nul
X1WAzagOp6NlCLSrCF9WbHQ2bz5F5GvWYdjozxiwxaHIbMSuImVaY6FvrQdoBYO5
rdOcdttkzyfZfji/Q+AbZtbHLgNNinrwRSiszahW8tTSnbhwugRnRYgvzUrjAzau
qTKKs2mxyxB0nLCehJmB17BiVXfHokC97vsOUJEsbEbq97lwlQImV4zhdTMej1p+
Eql5zYUHsyHJ3DZyB8c9M/jkYfVNZpCQmSFLnJ1U39iJ0ME210BrbExvwgeY+Zad
dvVTezslh3lfjgA6rCoujilAocEqkkoOa3R9GDNfOmo8irGK6Mi0UqRfx+20rr3I
MjgKe1nr3ACd4TccmWWsLyt5b597jpVHOWV36vx/n9wm1YmwnaAtDOwZGmcZdDek
6f0+rPnajkMQz+KGGX1mQUsdLSHofIA22OZnqydyc190h+p4+3+lBcUQduPZ7676
HfvZDO1cJKGPoTTu1+k82cGpdMl7NAell/wPK8I+NgkZ4n5QmE0bjs8SaFiJ5ESw
oIgVdWn0Hp3PSvJ5q6W3snXh4xl3SQjo/JwBuXC7C6j9JZHMcR0X2V1uyrM8naSG
R/E1nitPNDXa2j2pD/xLZY7SzDT9Ud18ZYN6yTlQZz334e65jP2KmwbDO+/Gbo5g
ygDgnjH/rymWM6okQI4ceZz7b2LzKrpKRu8+WJswLIpd65YJ+CzHtk9qKzQjWM2I
IocHvTiXERiyhxhc0+p9aoTJkjQqd+5W6G8gTatyrNyTi+HpaY8p6QK/K+LWWbZ/
vjsM/bWAIUVR6GGapH8PmG5m/aiegS/i4MrvAV8RUVPYUlIbx4fn8dYkgk1feiaH
g0qynjSOheAM+PIWsPV6TotVa7PE+RsB8sEybSXkUELz0BHCIpVs9wUmkvYTGdWL
ZPOEab/1uoV3rJvI48pEoxQUkEZDZ0A8//jpD9t+WVOz+wmmHILkzKXHePrjAVpE
06dFA0k7GhyiNfxz562dUklZMjkA9PODbLrmGN6/d+qoi4E2sCWyyjW3NrKZiDvy
1gBPgX+9e6r8ru240mwNEGdC34eIx2oiwO9KIjZYVZr3V1uG6YExSI//k9AZo58F
sVkUH0dtquylqFxOJdtu+NEMXHHlvSmCGjzTMqOPSeDn3xclbL/SSHBxWw0JAl/1
D1YGv06RtPbWE4v3eFpbpfISPnVtljFBy3nDy7dMLuZMp7B6Oe7LIjK4TldxiitK
uPZAch5cF0L0ukMBy2373RY3uhdzPAciFapZfAo1K9nKKKyfQJtAdAoovTm7WYpP
jnjMMTabtV/g8K41B49y/K8OFJCZ9DAf1ts4NTpdx8yzOvBWnI7TzcOG11iuFuEH
BER606yylkkBL+0gsRfXlvkLIK9fEoXM0v3Ugjajba3B7IRqg8Rtckao6IyYdqDM
ooz/jC02dtNPDxQAzls5Fx3U+s+HWPoSwhkRWHByw+8Rr1857WJ4l0zrddy6AnUu
8aF9m2HRrL4h1Z+oYjgTaMotV5w1wk37QB9Rh/BNE/SQDz+DKYN0LqCmIKhcmwMs
W56E/ykZ5pFpK6DFSqc9CkMqi+JvDF3fPOenxnKI1oevBUz3KmQhq9PIqbjkPV3O
kxKmFOC1VVMl3P5ISWYoo0QRTuh8Z+u6j4+Z8Q4UYH7P0QWJ73MoxEjlxIzUJ4j8
myJk7va23JXyCgnqUsFUNN1aCOioA8c2qEwpcYixcVPNPwR//1yQ9PGk/Hgup/Mn
el7VXgZ6jryMaHSCN6T4ZRtkw1nZlvbHQ6izTuhl9UvTU66f6eSgyEyIMI7dgOE6
Tc9YQC76Os1hdDkkNX2Wv0rWJN1jvM9cpamhM+6n6VYJ6pcGbP80fcwmLkgLZRbx
7rP+ayQJySdUJC9lTBUf4fq7/0CdUTzbzIA/31yesJIW9OhSi0GFPFWluSbgMtfq
HImmXLPtsAN9pXLCKLl2BJ4aVZLh8KTdCVG6nqyrm0ATLs3y+JfPn/I2kbq6dV15
3EOd4ANALargZCV0MgjcVS/O8B6AsCOGGI3kls+9+BAt4M3C5A8WXTIeXBQloXaz
wYX4TJNp9FPo9FtMVYHM7F/tw7sa5y+WjhMwhjp2qZ+vORIqfxxoy6kNp2Ikb9I/
M0cebBoz5/UyWAaMcjdHZDo756sWnATeAmn8MwxJGtxcY1tSd3syn+bhi1vh72Ze
KBbHdsuppsS/affu5nhqRDnHUqnmNv6tR5ahCyrdBN3ycC/OQMogA5f2Ymy5oeeX
ZXcd0819KtTV1a8IKgam3hoSHHl42pLm8/w25sGiKc6UTSVuzED2QhzwJWoNSFbW
kddxJ1xpRQfzyEKTQPmFQYs4RD0KVg7cBA3J1C9lhpxdLPyBTMNYNbImipcx63gO
ndoU7eotPfbUpq7+efBbux8hX9JKZO9Yb1e8JNWecCuN4gk/l2jYB4QThlJoIO6b
ZRzf6LlhoOyvE3EYqrJ/4tqe6ay+sHc9Z0b63KT14o/cpxn+j5YhCof1hk+En3UQ
qtUGwu5Sk5Jy6wm4vqjP0CLPPbVvjwqoLR/OsuBPVta+qxyn678Fr+lPfOZr/N2S
UuBrHTFZjOYhzP3bY0ctouGFXqR3EgVzcFK/rkluup7ZpfHis01c500HFSkXkbIS
Gkz6fTP/lJFGHWt30UvwjS4m6slR7uza3c27yjZ7mnx+W1MGu4vQs9pmwKhGXLVA
XPkPhOmVsTmtUviuk5hEUeFFNlETutcoQLPyx/m977SMoLeWn+xoCk/zgwoeEn4k
qwdRP8oqQGQfWCZAKRe7tqDg68ek4xfziz0k+ATRorI6izJ3dGBD0oAc54whXjxn
sbQLGb8ol2X3Z0HWieXqKllVnkFaWfLsxv0mHkKalNXo01I0h65B3UAia44Nurgi
aIPAz1q69pJIJrilt2lXSQj54Jp/bZspkL3a3+mHX6vlYExJElaQk2lDrBjETJ2L
gU4L41ZtWvtN/kW2ztHxDGm3c1y+Q5d0hiQ87IVpFnQmWN3j1P+vqFWIYbz3z1pQ
A9f9YNaWrhNzk3KYMX6F0gyUJMTCIUoq33Gdx2HgwYiNJ4uM4/gqSB3WQzGQ07yM
lS7tBlGaY1FUfcUZmFdNIsfyEh+fnqLcPBRtny/WjAqAeszGt4MAdg8Nz4uYvhDZ
OTCepVXR7k8h16nT5vq4tBecCGFqXW8FtTxT+Amt3mtLOFm+hsiU9Vv91OVm1Ch7
dhOJk34rFb22Zs9eUZEf4eDruAgIxD8BKewLc/w7AFx2L+GrRjXwEjvnAe0J7oWY
LNWZw8ErG4cP1Al1KYwZa/cuJFNkhGRuYb87VzCe0aFfySHYGTrts2VCzQQGx8/g
oe1kD/mf6zgytMezA9Swl8xP30aSVkXhy11fJS4bkbZoH/FBoJOv8XICJ24uQ065
YFr4Y62Z4m2B3uxXhL+qKlRR0wz9k9ryaUUva4jB2xJ04TFUFVhrdhGvu4HibZhO
UIQJCaWRjO8cTJBPRvFsy3k72TPhXn0Ze95/iEgD+Ixcw0BdZN33/e/RaSZiaecH
y+esVqlLFUPzyt2KVWgdkz4TeJQVvYM26noEPPHXEr0=
`protect END_PROTECTED
