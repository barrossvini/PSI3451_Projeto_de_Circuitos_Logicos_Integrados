`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ukHMkoykkxEv35MnSQyc7+LLUCXHkgt9BGHSyQURHJDohKARLJRBG9S7gPx5GroF
bh7B1mb1ExUOmsjHtPczd7PtJch+5l7DjQ6GJyZR3MZxOCG8Rw3BjAKisI1s7tL6
X9/nbaERf4yCe3k8ca22OAO2OATx98x5sUWNjamilurZf1kt24mDQvCkVn4zHi7u
um1iF3XhhMmJjcke+Sw0+SWcjtwJX8Jg0mJIP1wGdwIBnkhnI4laBbjXIasmMB1s
V9l2rV5VVUHuoTj+pAKOU9VNDXvnwYNPNaepRlV4HeISEdFIVMAoO4yJ2XlTfhJU
sSA3USnxFnzVRmT43C23ri5FIWFGT70iMO7v2Xwfm5dPxmNr1S2NQmj3DzHf8ajd
K7+Us9q0Zfb7L1bxhFEAwkBT800qU9dmCi+dAmGQ2sCbrruQbyHMlaEPmH728fzc
gsi+IWghBYrSebU/yTBBn7sKXrvoNSfam12gnVu9bxQhzFSvKDkIzdwsyqGv+ooh
3I0Khf6CuUHEKkD2YhpjqTxX7L9PpnCsizLbQQmlLF3sD0rJav3s+eQ3Sl9SuIO0
G/H2t8mu0UaKu7o8TRKVfIYudYl+Vc52mxFKtk+Sed64Fvb2WD5MBMYKX4eVvi59
V1e0C6eKINhGuSXPLZ9JSF8VwKoQ8N6fDUz8e5xPWcNRFVlSKPIQRV03FhXwPeXW
p+adCM6BtMbN12H6dsP5XwX+gOPeqoOFzE5yFpFSsPW/BjFb+Cw7+GoeLH3oNVk+
2dXn6IbpHhNuxQZHEpdOw5UUOmgBVYLDxULDF9fZk178TAeu8Vs9qzng4rFcSy9C
v1AC8CXJXEKi8f7VjylLKQ==
`protect END_PROTECTED
