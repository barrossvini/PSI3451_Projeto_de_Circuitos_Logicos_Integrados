`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uLwQkF7Df3A/PT+6UgS4tU2BdFIF+qS25yhJLQdrYNx0WpNi/OfT+Gh8J9Coc34H
0mML8dvwBHv1etKcXf0ui/eSyDge2aduzHOCwjSoi3U3xsoxObIo+vwE/lsZqX5M
2Tavj2jID0N4jgsNJOrIHJg9oUReHPaBt5UeQxz+Grgy0IKJIpNrpqbE6FJkDRs7
o3YNg7ePTBdn1NAyJXYPze0Jr+UPUwZSGU4bRaiAbX5yaSoFRKJtI+xpU1HwR00Y
zcCxxlT07deLu71apz6MEp7q76pes1UZ4vQOuQ1ydly/dzkNUNvmya/x3eSwlDdT
EJU7SKJX4NdZtpQYfXJb4100WeR6e8b2M0VV1b/MOIjicXj8/fNcEndSM3wqCOKJ
NQVkJ7cizVMUzWPGnNfJXGTgfG2ARQTjRb3/OLSMKEVT22DsMrI4tCdmedsTevw6
61NGm0lma34ZLkyqHf6sMha8p9DK2TsBgdvoKXtedMnzQEP8ezkI9yOO3RpnrIPC
eoGqZV2yRQdpI8C3JrtLqlStHk5YIeCMMroVRg4bB/8cnbOm8PzS5pHag+KK3gJw
TdEUR1kAgAK+YYZnOa6FmAaytLBGR1OCCHgjHEwhTSZ283QcyY5SV9q6oVAQkGNI
OxA4jGFpGj292igO6FOMW0VVg+bvgs3gjdN/zOarVhh7aYhShQVu2pe2kVqQVO3L
AvNqghtkoIMii91BUO3ONJ0+lg+yY8k5VrF1PfZzcPQPo6kwewEzP1DiXuMbRppe
jaq+0q39Qa3L7DrVxsCmzlVb0m9MJU9DvRSjTVkRvT2KjzRDLrIt9Xv+u2ClhB10
uMR5FoXAAoz8DJsadVfG+lRzo93gEqc/DUtl+XbuPLNJKGMPWhpYQ3RWTamTnJkW
AqiiCq6f4lwjXVy/uTTuFk7dNRmh8hqf6xTp1fHephuJf+werehzRoo9FyWr15qc
FCrDbSR6GmV3woQvVWQY6Yp6k/ou2IcUB1QTctEpeBBrZnJg9GQqjBCePGeisepe
eXXGCd1KW1AsqCE4j8Jtnv7qFpzlW8lD4baOXOQaP2aNsXPHlJwdB0lph2H+bJ6e
jZTxO9D0xZFpHhS9xdO1XKOkF1akdyv4ya7DUgbR8gU=
`protect END_PROTECTED
