`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/bAsSfuWUJXXEP2qzM1RiNFkGaU1q380yu9xORZM+i7jjxFSOPP/knZ51KybzA4T
LvGqUwZ1JwDrEy8/qATs1rb7K3hSBRtZo4kB2R9W1AaDplX03rZLgd8aWwN/LwuU
rb6k1XKkNw1lCIXPIeQo3GpTt2O4gJ8UjuTjs0dUC/6fTxcTj+Jeh+K62FyBtyof
Gl02yh1Z43q9+qQUh4EDMUPK+n7yLpaSFq3W/JqdIXC3HBsqRTPgU+Uct4zbfNf2
xWm+sMR+4pjOsQi+zmdXE1kTXVr8A3QoJRfVI6cci1G1f14MSfPiJMHLZfyRjvSy
d21b7M3Qeos6Su7lCEaUE2HFDpnn4zPAonAuuJdB/D1aau49NIxC61n8sLZBW9Ol
5IQjw2R4h59uzVyUxviFoTnR0K1ze3VRZp+CnangO4jibN84IgKIXGlxEKUXzhNW
Wyc7d35YDLP9V55vDrPuhKUY0perGQWZ/9xWkyLw16AzPumF0xjtbALJhK7hZ8KL
566XBYmqugXoeH2q0OWGPvSmkUFUFPXT7H/ulz+sMy16dTiAUnNn31R6D/g8QVZ+
Xagp1keLKm6GrXJzCyw0tbnlefN8YMvhEOLbCChZKYXr18hgMN1RQEuLwNdyq6ac
XiY1VETtytnBPJUu2YnRLqDnWFTT8lDKDCfIzxPNKGh1VYVYhi2wbezmez9qqXdX
iHBANVwArTwD3B23ehtl66QkRO/0GDXd4YOklRjGGa+Tqh6KvObxBvNkXxPGyG8Y
zZGYebxxIDT14oFocUjGo+m3Rei27pwe4otMo7VOGoOM5SyxsIltvtCLBwmq7zNy
4VhxKTunr87y3vuKMnaYQUOVpwZR0m9N70Y8SROtvxOcgXKILQpjFS5r4/W+bcqz
8ft9G9fytAR1zAvfopyTNdgrXeaLtW+bJboMCJ2kXNrYk7F4KX6KZUajGvWN0La4
dhGxIXxIIqFlNbFu9WEGxt+DfGynNGH8s6UKECLg+B7ZKOpX98lVucm8M47zDXXl
pVwCSFZ6cFCehs9JyL7J3opRJM8HFIRSvi1Mq2Ww+X1B32p2LF/rxqccblxz1vI7
UuB1NiVNhOHFqk1LgnqTyyxYe3p3ylYBDmpPfC8yovnupgQkw7854xyCAMxdxTYd
L4p3Bs3U7K1E4ywkynvdiIaJU/RL6EgG+FNclifxXU8viEnidtjcUhDx1Zji7seG
x6tQL4j0H2NWcwP5mVxEoLysc1O9BpN/9Asf7Cc8+QaRRESJDb4Yf9wFMhwzCw9u
P+j0gwDyF24S4Qavrmkz1BizUfTtAKNUGpk/qe6rxfTyBn6BGFNtjTP1FVptQ2RM
ptupfqXImxkWgYoMqygvSkAhlfWlEY1CLObelEVZUB8lgydmdssfj1gtvguTta/j
xsUcLiRamzer1K+UOu8bLzwGUCdtZGuEr/ce6r+Pi30yG7RAiYUdRnorSd0QgpQw
`protect END_PROTECTED
