`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJ/2HwTAy243njuqx5WLyUDvPL0szY3yu2gLjRcVDa0KTwE4iI9p3lejNDvz9WsJ
UYwepURko7ZEJn/WQQjutwofScUT63wXBA09NciDfripALRnlL4UNuHdSa+70MY2
LJSEb/7zOMlI1e4yAVIxh1eKAYk73vaXb8nmZpWolvoaJM78bkNRIW5928aT+fTk
Hu5MwnYdfT4Ne6eDGrvhlvCc/7qNa63dQn9RC+dfM08I5ZpICzU4LOKZ3OjJ4OKT
t2Ao/tTHHg6jCyrpb6NeBPbQVpsejqRkiZjS1Be3v1m3Rq/OaDAfac3w+pfqskU1
M2/GCh2BCbx41isUaj6UmTvRItHpCk/F1O2sLnhGgDFZ6bgmtgSCPKGwtmwRod5O
Vlp1umRynyll23Kg/6aqxLpVOg1YclE1k5pwNnKkEDH0t4iXiRJ3E8HF/E5G+5b+
KX7EVtowmlWbyngQnzZp3snGAeRbN0nVVBKqFXjSNqg832/Xz/UyQYvFlnXO0g88
RwiVKmVWdkrT69BdP2P5+66ffynawvgjPLGiQmeHmDUvyedHm3hdIVNZrx3Vy5Pa
GGcCli79SufR5nlEF/0YUp4iltzRxEQK2IzjapWK+OSBg7t4LHvpqGtw2wSQzMEZ
8DIWCmMUkwxE6oSADD7Z4LPCkvSd7Y3Z9czAtOfK7O8e3CerCay3hnQAi4vcSeg9
08HFYBZfllKyLtb935zeq0nGfzw+RqfIHq/5mTWybolMUqNIz3OsayfGMe2YiOke
2gbPaRuCY0UaAYqR+07N6Gx6P+YA8Y7EddQm3jYZ4G0Hyi2OoVyQiHwZdpM6uJ+r
i+Q5x+WdRAiFbmju2VaGP2iAR8LIjVBx501nMoJK6nGNvnFdgKPh5fiffNZv+FJl
4wrXGlbNu8uADc6B+OrV6w==
`protect END_PROTECTED
