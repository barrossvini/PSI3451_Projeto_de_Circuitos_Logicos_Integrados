`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+Z7AcFxzkTGYJza8KraFc+7Ry6Gg91OZZESYlCFRw2VCf2/hzWyFsuho9UnDpMm
0wdIleOT/8MaZ4HYRO8ut2lOnweDSGtW9loaEjGVyohvgrzZ4st4CVvckQiQG5wj
BwHeIZEfRMr+RX3JSrmCykx8rlZHeb8aPVMjEd+MBdiPIt479yvx07g8REIAJbpY
j2DhlKkBwIc3MMspZp1SUxUO6VVKBcFK5PnUQInT/cJD9j6/RJjC7mkGPqYYxS6w
pLZvTrS3YMWf/sQ/c9Ag1U31Pld3tThAsAC92osKONATD+fPPkbfLI1vRp2ty5Fz
o2oLxGpd4wCl9Kl5SvbausrwXfaLFz/+L7ZQU8bx6eh9czN39tcB2QrpTLfhv1Pi
+jgK5QvUv0UQ7DdP82TyokGEVzND+fWDLfeA1fwDXQq/ZGpzhdShWph9l7min9/H
RRNI2WNh2LtjqKu/BVKv3+DdBR36foIl/VJKzsqHJ2oJgMIOlDUMND9OGjPaZd0A
LWvFd8bqOAelKZXYr28mpt/4kYaZCv0E9ZnvXVdmr7WVTeVZXTKLjLKH+I9ANml/
8F7oC/DekLW7jxBT4PeGXXoJFAj631g+hOW4HnXbN9pKlXkUfIonSf/TFbq62Z05
fQofNpY9CJVNPNSDPXzM0zHtOk7ijWn1pOCyZ9R3fOP/JWqUDscj0nIKq6RtOBCS
6Kc8bW4U28CwDVhsW9prp5GNva6pu+vxv0wMc2ozr7O6caluk/90qaXQH+8bC09Q
ya8Ewat2IIgCRozo7LsMeG69E9kwWDImQO0SreY5h1yj2GJ4SjYw4SjLLtpuKQQc
ZF7A+LnqsNBJwvA/rHxcgEUXsxl8FC2IcwrqhxG5wbhifi0oXZPehI5L9Dvf0XC8
//hrwz9IT95ufxzImrpS8G6Ony04dKNipaIL4ujqhlQoAVbihJVvVNCPOKl+aoiQ
kifhWky9yQD6vw8GL0RyMRmt5mLpK75ozGj1uMF/t0MxQqVrDkpPsqNZ25HIgXxy
PklISIOxnKKCpcx1UFcFtd/L0SjxfvSiZKeDT+3vzMqoWa/beB6OCkUVJzVXQOi0
HLiB7pzCyVon03QrFofdi8IlNxnbAmpn3/MzMD01cM/BMlEqlp0g/fHUlRm1g/s1
lzcEm8pFm+ptsHNDRzTS15u6i/2bBbQAdFROT44LAyVZrTXGYFi/dwYg1E1LTZs+
UM3gnwKMNxwmfvD3qtU2QPV02oDZEU1WjNemuCgjs9kfmYo74MgSs3Senbw/XP21
AhN0hfNNp5/QlOcvXDZjvg7JY2cGnxq+fHXh9V4Du+ET5SKWU5ISAv6RcQgQA547
+CjHgf6I80Vow55mncOkAyPfLJ0cCdilfqpfaCJ5kSx3knK1avNs4ITgT5YYhZF0
S9BdbUYQvI7IaRqmW44eZ870b9raG/x5VKWiQXAMLWjcn8ecgb8uj3Z1PCtNNGBV
TF9yWq299I6/AhcrGiDBlXhfxnGw7Ya8ywotLIEWEnP4MuxMJRa65Ab5OAmIGuND
X7Ng2bGBIEqyZHnOc9QDu8Hd1oajadKan+VfH9JKilGkJtg0QtHHqcXn88/UGEtb
TIMTy83MZUSOnCS85luGb1PeJdTeMzOhqLI5tfs0nGxTdZKcgY4xdF4ncC2xAutl
vAWkLPvvOrIQkA8hYsESjqF6vCjflTRiu2wTC0GgNf5EfpNh9au1DIBgYjFVCqhi
yHR0s0v5Efv4AgTVuDi/f1o7C3OCgd4x9y6S0AaR2ZtFKcLr/cMxa0Oi6EQFNEba
+USfk5k+1QVUaHkfQESi05xuUaAGC2bQ1LwQza+z6aEjZ/+v1Ziw7D8gT0SQ4Fkw
MEz8s7HBllJtw7tcZnjdKhCym4AUsSTeMbPNVxeadOVF/XzQ0rhKlXeSnp/0EyRQ
T0mFP7SFoSQwwwRqVZogOcl3zTHZa/0LVPGU2er1SRrB/xwKOuNhRedj6nL0N7Nq
PVUdqvTfHBrVNF9IQj83fnTLz7q/02fjB5WLMlB8RLjqU6Xyks0CLZshP7s8HRCC
m+zRZ648RJR9OfOTMAvQajNqzPgOwkJe/ykGNf33v+EQnSHReriB/2/RagnMbtu9
VpvJ4LbEOnCUTu6ZYfj4UZiZj1dpc4a7fGwskDuPlt8ZHDUJtim+XlzrUseTNNTr
rCcBiEtdVnVye0QwIKVRTyh+jPntJfNQUzSPFEN39o6AN7VwdlxwhtaAmMeBVK98
A76/dnWL4N241IQt4OxCArqf8pEcDecX/UV/TvjM5yvZqeNXByjRvb9wRnhgLZ1+
LXTg1PCHcTjguxV+V4bjEro6pfyWoT3NuWpP7GdkY8TL0DYaFy1Q6VH/lPypnQfX
G1xZcTc1mAGb+C/HnJY9fhGNYai/7XLDLAzqiY9oLKO9qLo15CFpT1xYFMn9UAPJ
`protect END_PROTECTED
