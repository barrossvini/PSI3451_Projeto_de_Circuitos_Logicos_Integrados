`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAoKO/BuwU6ykIHiodTx3+zvM8be33iCJW00q9tUxys/SrXdWZktugZY5sCKfJy8
9gMUUdGmR+WSs00txDWZvrXtRUOBT6GOQGDGHb6nS/iGjoE0/Wh73tgiF+DoAQwY
JrJb4i49CBbkS8IMXHvqpAlpUpFSf2XSbkOHCttRDClWuExNYe0L7XB3BSEpTNKH
/WimWSqqA/RvICfGbi/IQbkbjydmZ1pOkJQnXwclby4DA/HxMNFtRHRsbvJmd/Bu
rFJEmf/TkiD8NsI1hj2k4Iun+/r6SRPZNvArKHVm+FgQt+hN3bxAMSpDlyFrQeEJ
aiCt/F6hrtDu65lhTC4ViHFXSNDq/eFOXOMoRIH5WTE/W+9DUJ9uCjhNFP6fqSNq
Hv7LM4iros26SngjWw4HbxIiyB2HMsGqt/9Ssro3dCmUhLYmMNMjmphaeTV8sSmU
1pHzdRdjbgA4gqAaMyKs317GF0Qsrv7oxA8Tb1S1EDCxD54g5O91meztn443H+Uv
cAg6VAvfFKmWXz7PZCLLkdWyz9AG7c1xUgpAYDoilFwdJ3kcLB7dR2XMsTW5v25G
78IPrAsse3zi5g7UsjR4tKCjkDlq62HSu/whBPtB8lUBbnEQLf0d98gTyX9vQztV
Hu/kSQizptNf6dQbB1n6RvVpav6bY6Tl6RYhTU3w3ag1wD+OPTIbtnUoXuV5sdKE
SjztGQN56sNj6Ig9Q8IPg6hB4O88mOIAA1L9rJYKmaazJ6X2g2upWGA8yGTmXXD7
xyS80x81FhVvAY6eY4r8BSINAElrP3fwK4IpO5e7MVLYqELAWlZoErMtY2rpr6Ba
fMYNiUiL/0RQS56kUZ6FsTWzv0ELlPvaZosMWIOHDQ91ckHpIh1Oa7+B6t0cOFWh
+2mgqe30SEQeFFTXv+RhXhm7clpeawOSF1ISa6TpW2N0pt1Cgw+NiIuEacOQijgP
WXq3kQc8bWe0CuI7pjEwKrzY3SPl97q8IFRmSGPOe9sVRKaW51DuV/1LFL/6ylaT
BEppkz4PfnzWa05xXJ4NVSIPNnQfDgohXBwfP1Y43n8sZfP01bzRDHJOC+sKGw//
A+ess6nja/NHbwJhFFN9N+7QrdCGrejPS7sQyXpOZaqia/9OGqVhTmpedcOZ/OUd
J5gEjJTybMmcpOkv2+fMt/gYBTYnAl6Eha/kfjKUQBY82LqL5bW568+l3PVZHO17
5XTa5ixUIZThv3WUyf4vnEzUMXHSzT25aV0WKiyVLJGiAZtIXhQC26i0iGN1xOQR
BBFBM337257HLKBLtFwfshW7OLkP2G34uc6jWgDGDR3Yx2ZIRrbYmy1i7B9b8GMM
gXBaZbiwkV/HScSMczRCTtbHyhO2eRLWWe2ZcKzZxjIxNZ0E8XiZuRCokMc6oN+J
peqJYRzGYCH/4OXcCjSzgxrDhR5axSkxgAtm7kUMYtWsdExX762uYPS4f+uPccx1
n7GLmDezE8OCOjSKId8BIU+38bdkgzJaynLLyygds3bBlhyvLgNoY/GpbquPbbpi
Y0neghM+mI+vZLGaLO7A/5C9+dJrl8HzkPpLYzijdTkgO8TxMkrCNYI8U2p0ScQP
WK9kF/m2VJTYMsfxLCnp4oL25n10TOonyqAFYJGGCZUD4KjyMN5HMpacogYK8W4d
zjhnWm5qNYxTYVCdC2Jmt9eOLkdjP2pUyg2oXvlFIOFK4tvizFqy7AMEysazYmQv
wmA5Sd1fugo9wuKld/7Aiq/R1VpVVGbmcYVp7EajI9GBvTiL0fYmw1Wd1KXwCdwA
QErFY7NmXGJbWfL7uwYsPT2ndIOvLKnqVfu/SAK7QeR0DjnPNvKU6XNDqFmTjF9h
CmruMkeUUqTfGGywVZ4nKLJEibIAlgJ+SxpRpwvIVXOIne5Qv7mAUxGjrP9OrvdE
vRxBKgfkMJ5x1Iw3k21UT5Xsl63g8ctalZNPJj+mBufNdFiYnZQtUkOPUAg4eNLc
l0mEGnDT4rRYSrleT4txGm5bkUkxwhvN0Eg14IlpKK+JZSyDGyW5ROnRcxfDLwyy
S5Uy8NEaK/juVkiqypkzaf0smRWYn1kscUddHT69ObUyGnESbV89IKipr9tNjOwT
97BI1h+7CgoRHZp+MVwAw1OEIDNsW+5FRTqTPOYyHFsrLnHTVt9GKhc3VFasu1Lr
zO4knvqnNw0XfD4r9N5VHa6NMtrZGJUoWjYKDc63h2fXTbZVTp4+nqKMzjIdZqv9
4y1831prIDVcByg2k1iaq8nQQBJbQCoBFP2BQQKIRRpFylNWr5Q+HKqAh0wA+P7b
CNy7lmV/Y5v+q//5Rf2VuPl3m2GuII17fKKElJHLBQW3noJJjE0RiEeC6AuyyaLW
lG7MCPoQUnF+c+9v8XTEaYGais5EV8ZPsEJq2P2h7hFnFFrNYcNgInyQdyTJjIpX
CHv4eezi0aJBjJnC9stlRkHeSHEf6y2wAOhyGl5yiY3SQp+NheXWwLHXOtcnNYAe
P/cFoepxxTfYXaGUHlKdHq97P3OcR8BEulBtn2NeS3MC8So6WPa3ayTi2GeHr2GS
D/lY0ulHF0PQH8MWsGWQE+vnfNwaEczUZSdOStkr+cO2Go5/HpCa6PWHM1KGSRDE
tKJXxRIA8ZkqXUznwhNK26PXNJQsolNyArFzV0KQYwPRa/SvcuFJHhT/EWutAZTS
gT94+hcVLowtjyiROQvqd5F19aEi0RiV2SGPYbpUynKcRPfUc0qjVreumPVKJDAg
NZa5Frs7BdEB2rZQTJL6pw0BPgaRqcBFk4QGSrXDNK+TppUqdV2lFgX5FrEUqpWG
NQG2uFMh5iOsVOdbME9D6qEemzUoTQVWy4wAlndSAW/4R4ncMntA3KcnRJCfUVOk
FWs1XRfkjYdVOUjsMH8tMmS8VcEIles8VZ3pj1GJ9BYqBl1y2vK/yJ6r/fKhA3nf
5A9EopCWcJKDWgjI1s0WWbkc5Iz9cD/9ZVtzwhbgJDMl0lvEgdhBJlbv7vkgbYyK
Y48Q2A4LPMT5b5zykxGkNMZxZ1PTHEORSkbGLfzJnkUGaT6oIsTXFZs9muFJGkl+
bavX5G6K5W3UWTOZbJCqDtKeWWc2UkuWkhWHttaeDzYSESjs0gGQpjp/GShvOD/0
4yKFI0sfomGC9E4WxUbOK0LVf0G2mm9FopFk7hY1pSWh2FYRxua5PY2e0cytaPDk
p++NeZL73hTAgRXuKt/3smXb2Cn+9tnxuqTPIGEUKMa4q5O189TNto6pGz9OR/Rr
4jfLYzxxt40si7xK96jkWS2dkO5ck4nCtvPg0yPgtTi0GHHGr79uyysPFhA0zBIB
8gWttueR5wtd4I0U4saE+A==
`protect END_PROTECTED
