`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ud/tdk03J6iiOLRLeUhyFTTQmrhURSVixJjTLJbHtfOz3rB+Lvs1l279EUJD2z8Q
OKf0mgqFIfjgpyvRejKdUHzrkGViZPJ6KcDz7Xzi2UuiMvj+bnwvWRkHI80RvzIf
eyf28xL1LbrX3ZbCabifYon+rfzFygPnSwtmuP04hwHQGz36lnvffVqH+nvm3M/h
hh8I9HzWP8uAU12CQVYL+4RBflvWcqIOVjqc3PKfTl2BJLSapqh2XUixORM7QSxS
F4QtaZ6oY4+qxI+xpfjbCBtz8APuR8KV37VD1v+PNKECFHlhl98bD1XbWJx/NTyS
lKJbMZptXp5jEjvVKvH1ajMQRDHJlCe/d7SVKiiMQugtsrHBTuqctaiaLYMV900P
SojqzNBuqIhqjmk3esE/wQGbNReDGaYGuwMkVDvPnJn5SNYuTugqYwmy2xyvVe0c
G1xWAWh2nyKmf0aHzOnnT3Nh1dqcd95h9fb7KoIGlYJllPdZjAebkosiZucXmqEN
aQqa0tTs8prJBWjikMYY64JEkb1dysn936CEEZMzp6THHgT86sgz+6WTJ3oBTS3c
/0qCRaYMieXQJV/2WQDGyrXNnBbwXuEhDCabVs26l3SErzyYf25qqgHcwt5r+8OH
/UC8mnQiS9VBxFontysFrZw7idzprAC9mNwH4O4oBmUZdTyoeqmy8KEV+PAwy+2r
4Jy57Ki4HsJ2x68BoMEVRF90Y1r5xrh9NmRrctJ5O+9cgel2HJmEBoxX13nfEQmd
E68hmSUr+hD4DbCfMawJ5jRGXJDF2oVJFEjJBXNc08woJG29l79zm4MxP9e9gD9I
tAJYA3O91L1JwAh8Pmw3s2JCflWWRU1vI7EjgqiaOU2t/x34aekNwGk57YXcLEGu
uBVImKRfzI6pUXpxGO6Gq9wnOFVb8ygJuYrkxhAiAn8iLoCE533CxYVfiU2hqhI7
hrSh8t6SQWzdHm97o66qE87lyHfrvP3U54zF4/2iyselbDgwkjMZIo03GRr01xDb
TSAlCFvt/y6gov9BZQpEtVx7EgBeyuwb8yp3BAnuYRQeUj8Qh9mJMjFJehpFMgW6
Qiy5qgyHFf2/chrD/cid02IdXA4xlu+U3Xblh2feQUR4dEGNEzZtHpEHKdSYay1J
C+V+i0izGvV8QFX6TigY3VWV1sQJOD5NtEOq2aDWYOsEmrk698+a0NK41x9qBX5d
2LZ8l0EWAw9w8HVTjQx6ZKy0nsUzA7jTvCDd/bWFmWAbrhbYh6Ajl7XRLs6jje1v
sgGPBcIuJFmXsAw8eowwv0d2kXyN3dz4pE74K3ZJmFOdeAkzPmFKgJ11XyPThH1l
qqSwffTNL6WoeQBkfx6W4kipnlQIS93nYBclgyn9EHoAQD3tFFyD4We6ZfAO71Qq
PZ4FIuR+dlzFP7bqK5+i4DUe68BXbpiN3PlcuaRWs95aj1piwpeCuaa5pfdsHKjc
yPRARiGn+RJy5blzKOMUY01InO3pCsEtGnIVJcmnNZfLEafzPRehY/qjOpaxoCtV
oVujwF6bYOwFckCn0Tm1GKCIP38eoOpPO9SNAHQMVrQMkGO4BgfHGgP5sePcp+pF
xJxoRUmDtm/lmvSIpwdUnis3Y2h29HVc5bKDttqxMr0X794sOxTPTjPAMJTeJNCy
Gdie3HEMMxNSGchheBKB0tpaiPdg5q7PaK2NI6UFWLUr86u69+wlI6ZWoubauEnM
oZHQXreLxg/NXknhBU9egegXy7Y06kQonumBaSFEuyOucWWQfDucrrjz8SUTemKq
P0S75DrTwAKIxa2eGQXlYurje6e1PO1pkMiaMDNEu/ECJa5lRUvKuzIhMOJSlqi9
6Js8OnM54AKDvOk8A30GG63W6mfUtpEQvwS4uf07CrV/tqw4g92nRLzzn+63oyXI
r7J9G753gC/GrM6MltJ0w71J9kppT9f9nMsN4V9PGUSpYEBKiEuOzZP4ho6vNeiR
FqccMW8X5aYFngLZE03NSFIzg1L4hwPKR3d2pYjmiQHLgkxECWEiV2Vq/CU+mXir
WoNIEWmz9/qyb9IR3elmdE6zM13kU0a9L3MdR3E4vq9wZDboglXymx4SHbvQ++wQ
BhlHYozZBmaoMvURJMA+hnK28mB7l9lP9OVkcGvHTRzyT3qmcFHYI2ffuXHDDxkA
GjxyA7RI4gvIOCazdHLSTjnNgepvxQUcv8FyeE33O70l0PtmFNci9waPSZvTbVWB
sVyBy23NNYWN2VRzP1+gSv62lC9eK8DHo4dUXJUMK6ceG0lWfxWqXcdTXX10w0El
bx/xtJlVS4Ik3RhH+pXW5GiFSTqIcv6xQpwxWS68Qeaubyg/n8dkWYQcvbFJm0Gm
rmBShrpOrLpvrJ8xC5HTnsaaGUSwPoC/JSILuKDKqpOesP4tUHzu2sHFtBBGnlDw
dm8qywCbyqGzpOVxl7SA6qUL8kbI5rF+IlpPbCUbGMqSRH4Xj651Y2fmqx9vnyrc
UV1e4BI4tpJc2T0tRUy/9p4KGRZA/2p44KeUhYRq/dsXprPV3ZxR+osTqw/ZT3HK
LY98U+7iYy8vTa7k6x0DQqvc4ur4Xf8T8KFLNEK8rMcsQz9Dkojg93sgCy66O7Aj
IQWeoKLObjHR6cQ3kfjN2KXNZNLShO6UnyFe1x29MSQXEcVKxE+k50xLo1kRi8vv
MXxwogrvowP2WU3pLPM578Nj736vlSyWKK8o49Pd/KjqduogfLs7xrM3vOTp0ub5
MQWWphE8Wj9oNmFGK072+pW3ZRiUW15nvyT5kr/kb/snZXXqhkjc5uJy6lzp4OHI
yMP5xj8Yg93WCXTQZvCQj5e5BJpdzk286x3fopPxuFqrivz9mQ0ivZOauHVB1nPV
V1O0CtrRy42BpTNOKGASJxqr69eeb2cQMWWbDTjADo4=
`protect END_PROTECTED
