`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VbV1dyqheoqDcGbKkPgYQsmmdJgGhl7Ttnahs5FY36LwuozpXDGDsxKsp9iaAoXz
2pnN/mdBVpVyfnmDB5c7XKJMS2gaKLbrgNRz5trWnwXShTZ9F4ncVu2qJPyXdmXr
M6c51tY15eqytH90NZrY3ge4V9zH3Orp35fGhDwBJ/r4Dw04B3loYUCWR8uiyg39
8equb+Cv+I3REAEo1my3HfibW24ymY0exg3PnA2jQjaf5d7CqmU1LmBgsWK5jVJj
GrgA0QN5CIxFqKvJZlmdn9VDr2w+PNpUrq94lzZbn07tejNxIdbxISLivVj4vwbQ
g6tiXN22tgMrHgU2RNGWkMfm1lVAiHEw8c/Wu6Y0RFCxlyuIzxAdRVQK2qKSqb9G
jObWfL45EEZJ3/aLCHUJiUiJUjTDrkfVfJlJoUfjqoJ8XOvkoDeVWvl23r1kx+Hn
+iAmwvukhH7SfkITu1k3+WLxmOyiB4Pz0N4aCDaH+ZUfm8WeGA8vW2DzHOmYKSzs
0IWCCpaVAW9LPlIJqepRQBTbFbYdy987QYd02niTbh/5qVzED3vyM30b6Rt4Ivs3
zaQLjywpI7DtTdZ1FviS5sBH7PI1Dm+ttMGKt2Rr6O5J9FSTuRprZ5wKwZN9/dBW
ZGZcbEUpVt/dCKUd46ZqXX+DLC8OmTSuYn9qSeMTUHbalt+BoPsPO+xPpAzFbIpc
fZWd73AFtlYRN0T/MVcgA19JFBJJksA3FRMD+zo/yn565XRTGRUc5GDK5Gp5k6aS
MVICJbIQqgmbQ3ao+HbOYA43ZJr2xgooo7pdu2pFpdzO5+5rEaInYUP2sIzI+Oj3
Z6qo/1qQZVCOY5ztFPbMOhnkFmWylyYO2AmhtOMUPpNpPtmlvC+0KM29J0JJz/Rp
JIIxAVbpP8DcxUHuHsg6tb15fZ+YCrArk4ug/nGnAtr41Rqfimtd6d4CHuQeZinP
VfJqphyxzFX4dNxNfR1/6TXFSEeBXCNNdA8DijodC0sF7KEbgtPNu1J2hjjb/sP6
dRAHedNkCu4T0Mo6k2OLkb/o5UdND2Et/M45UikxYr0ybh7BcrT1oa7A0H1HmRSd
PbU/gOxsyPoQ6Dpov5Y+mBlgaTyBKnNQb7vSIOiHl1jegKiYle4hAZ5lXxCb9HHW
MsVuJ0wXhy6gmmlBIFmQgf/icO0hurFmuhrwmEJGv8+EMYZaGbJZsyYwfefkQ74O
+SGJnAV7fHbEjbPlzg6FRqFLpHfZzaQDPkSp57ziTiljrjo2yVyEY4fvX1cZQBYB
Oe/PV2Sr+YTh06S7HD3Pfq2HXYJOvb/ys9uVMxuKUSoDgo8kNKPFC4I/s5r/uxO+
rxgPfULt0/hr9766JGaSnpmULneu6mXI80+ut2dIpP5w/3O9ywqb7xu59//4q+GZ
GMlzDcvtreyBrLQWvxrZs8IEqdLMIJLUks0T/403Vzltl5KGOquhVds2QKEhbLHY
c7V5Ht5rPvFJ0HfrcpvUEya9QCRaEZ82q1w3+A4SiTV15NhSU8wustoK4K+KSf4a
C3Ba3NjLBRZE8anExQgYXg==
`protect END_PROTECTED
