`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tn1QjjlJZw/7Rplz9i4Vasxzb/hxwXZ9+jD7Oi8MDrBxJS26Kb9MJGjA2A3qniOe
7JUdEFnRoawGriSCjKj0MHa9ViWCvEw2pb9RlS+94wtraTMiEKBUZ1ZQGsYAV0sl
StLqo1PJLeqwvsZ7dHlm8PphMjbS3cterXgbK7xA83NDeczgRRyqxh1nH2wPPouE
Aw3D4rIuuMMW8X+LnN8tLC6Ql6TE9WSXlOphAJqjPwLS9SaOJ8JGkle9+IU87qfj
Rd9luD2TP+VJgqj6qkZCEw==
`protect END_PROTECTED
