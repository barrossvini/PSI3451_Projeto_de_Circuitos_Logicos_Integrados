`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e02iGxAZjseyAHplq9yn9U9wNfVL72FVEh9uMWFpPNXC5APZ5y0xZ5Tg++x7mx41
Z84PB1sLRBM9WsQEFw1SbqjAd8sP4OgdNNS8pcHAyJSxAYa4hy6ykMkKXE3yKql8
gA2WLYa2uL7Z2FVtXysQDIRK6/XENLxsvqnGvySYSEqDRXN+SYDiDt+7V3smNlEb
WMuWD8EE90cGlqVSTro2Bd5fJ02HhHsC89hBM47O/z4+udWH8vAMKrmGmz/sQmwP
TMHV0pzCAs3JOTJmdKwfjvzn/OlJgED1npFzF4CqEDQRUTf5XppAqhiMPfyLZpg+
ssYAEVcILE8zfjipMRoTUc3q+71LM4J1/MoLng4v7hf5oKqBwtf/a9oqpGCH0oIn
C9Pe3fWbU3odozl2CRII6sfzaQGDAnNI/HEPSM7ECvXQwPqgj7LdtyC8DZWoqsZB
nUtyr+Jutyubq8/F8tNNQDcGje/9fHsJfzdU2mXBesAOwPePt8l0Ced5Sd9J4IvW
CnItl1xOrHZIImlICA8PFuJdjcatwyw5Mgbrr/+xXyAVyhXmx+37zPeB0XmyfVhc
B9ZOxp+uVJZvzdSpH+9M3wBUN2/8Zn6qXN0oNIiIQyFt7A/az/GxiPVC3FU8JWJk
I/NLJ6OQRdgbYzcF9+tvsHEsdtpvphEDpw7FEwMdm/PLthyWZC1ncTozAxRrGKx1
pNDgHU1KgTeO+B+TqDzDQtWp3vkvoMxvOExRi2qwVOGTd+C2CVn84/4WR/kxwj3r
4k3j0Rx5AS+L83/Tui/jqrfPsqTZziHWFm7HmUdLkAosHOZP6j8kMWiSAEVDTz4P
2YdYKoWjgQESS2iqqyAjTYENXbInE57Lm2LAQ76sZ1/Kj8KfI6L/0c8maqyUZTQa
pGgkPg6DDLC3LDPQb0QGFRS8aI7pmCtqeHAXUW7MBI9pfOTnTIuzgSdrVWnkc5mP
hLpNkZt19aZJIkas9g8FvRbfbcwBETJN+evqj8JMpHrB/jahUqqVhRZ45ad1vgJF
vnCd1LQkrMVLlDr+m0jsBAmbBaEv7QhHMPmYSIkQnFSeS1rCV9TSDudHzYORNbmA
Ll/p9ZwNOs7B2U3vw3s6GFYRVBT36wKFcGZohYoC85g3GiWvByH6LFw86PLa3Y7F
AsYxj+BtzPCjcIk8Qayq0cvnUSJB8ngygSABzGQlfDsVDqdFZraqzMmGKKH/6non
KGJhBQY3diR7EYzbDnnbdQ==
`protect END_PROTECTED
