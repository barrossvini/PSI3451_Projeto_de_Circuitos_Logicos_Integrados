`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ykqDa8uVDngk6vJxl3fZFmhbe4ACjZ2soE34nM08Fg4uBXavSBaJ52UyuVkmX7fc
7wJrn7WVlbMIG+4bWJn2psqMcz5TtVB39j9IRK0Cy5fNNj+EKFjg5ZFRTBBYibgr
VwjX4qJKUOsuTeV2aq5RXblPc3wx0mtomyTgZq5NBgywz9Rinr6KWTs3GPhhDA4K
HVAmpe/XJ/0SD2J/JScXJi4NssN1k0HYd0KxGXrd8PhzRrmXupNtGf+UYrLnDjBR
WtFtcAJFWhyqFlhZDmUu6E7K04f1OwJ5sao8RZAnovelP9YnvJipDAgI6NXj9byo
39yVNyZz30/nzKXJkPPjcYIZSYvSrgzKUh96bz/+363e49I40ezvzXU+Dc5vePJt
D9quya8AgB0nHyxgd+2Fr9Zhftv1Qn9G9910Y9/y/WFUMnnOJcIXFqLGbI52/5hs
2VTe/PREx7z63LaVR4Myqz5qPxXojRkc2f214W2pGgwSONm0Jb4xD+sSBHEzAxTc
WhHNE/5dF8hqDl6MwM8sSifLeydftQeMcUhXMee/c2KoUnTR+fGc0q16IhNUMqjL
4Dy2odzpV95HL8FLbmrzSjihM3ECI+p7xMea79gprzUfEVhnxGtf5yMsbzzv62FM
HrniZGV/T8P+4tidCSo7210LsGnKWz+KlwkeyVogIplMog2FDFp2ykBsf2yn9z+z
BDbzqd/ohh6/bBYGfKKQbon49npXcty2q/87gYmMmQBmyRLYVNhgJuB1Wd4Z2EMJ
Kink+6BhzJOTs/wisTCFqC622bBZLOrRBHxhxSLkTRL5K682vDgaP9muAll71OmM
0RIn5lhZRsUrF14ayW7Y5w==
`protect END_PROTECTED
