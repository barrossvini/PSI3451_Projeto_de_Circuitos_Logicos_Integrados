`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qPWbooHe8KGotmS1a5LWCXCjrSjZBSf+QLMbc+Ax+WqkfugmTH2GoBaypPwdImJd
NoRNss142T7F9RLx1B3Dr3NVy+0OE/G9YFf8XuZZmo2Ka9TMBPuR5Idm8DS92aDq
48hxWau8i3bIHaPMl8OKWP/6XJ2NsVtKkTuERD/kwSBdvWecOvcszgUkCk1bavUW
wEYBoRmZKNXt0PYIhpVqHyyCrjYA/zVqX4t/m0Oe+Z26k4CzVSH7Yf2Z9YE7W5bG
WzlU6mPkDjQW12K4/kVvkOt6QxPIjm8ssAEE202wkC3AYES7JA58/UsDCS0nx8qz
SY64ppHIO561LgkToLjjrUCKEwyb/JUF+spuRyU9XURlbFYzLFu34UQ5+DU1nTu3
YlLoi+z+CijPXvCh9zQaVDPXi+CJo/WQft+6gNAZTdXDEV2LO2fllDxgl60WmmkC
JusbOnQuOOCgMIj0WhHK9YCH5U1wQBORzcyDzUMLgIHgdP6yIdM1xvIjUWXeyvC7
+vjteFa92sb/f6wGPfC8wdWiO66rcPi7cj5kN50d3SK1nWCS3ceCamXuqd87WiiO
niT7rPWv93CmnwDGA+JyYMikpNyPZUNDG713TaHocn25DCGFwoKpjnBo2ifb2khC
oMraU+xFwcRtBFy0Xg+0AqBTQ9Tx7k1n3uMLtPZsKdLdJVycKbaWPt2RJbRKRMdp
D8sC6C74tyr6bb8GdovHvl57Jqc2eU0AX1sNIA/GoTfQJ/0l7LZ4+gVE6t94EKr5
lusnHPLZH2oAl14Gn2X7pGXLWOwNXtG0AqQ5GXOiuIlLvDns4SjrHrLOotwxRRi4
j2MgSHGyRmM4qtm6UUXHCehji0qZM6zK7MIKfnt0QuY9oO3a3S3BoR+0utvasznT
lyiAa6QX2Xbr7cgXyY+LNkMrQ/W0/899Gn0cv7U73IUFhAuuGsSxgUVv19mXTzHn
24qXVZh1zY2HNuwdgnwyRUyOO/PIbJNze4c/DsMLOZgPDo1TF7Y3hDv3mMO6juZQ
h4p0HX9efIanLZXgaHtRDrVdOY0uM5xbni2fA1RnCy1D+mYvKFMz2zgJxH6CFGpR
buAZloEyOClZs0IhlNZNoKrmL0EhhKZVzPJDIecxRmZ0KjkhGJdzcBScM1nx8Z4B
7RlMNzNFLY7xZZJnBXMZvg==
`protect END_PROTECTED
