`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ya1G/FdxmZcdHHPdqOnEM7RKbnyUnA61tKM6c30dThUW1k6JLTZivUKw5C9Ow9f9
likilAS5qNfKAH31cTIIRLEqMCvftTjj8wYXfck2peOi5YQQLliypDQlgVyqoirC
imWsah2RXj1wBqsQae1x9AN7Qx26N5y6iBxBIXaN1/qXsGihxLzaWOjz0ZJWVLi1
yLEWNo2Zsac26gpWbYiYiXQqD/1p8hwMqjxwQKNEPSKiKZ470OJjEwdKnEYV6+Y0
6/m/PdJb30m5aAu3iSGvIrGkvVjahpbDDU7s3YUIRrS9gOHx1jWU8hATsu81ouLG
L8w9LdfTJYIJ1rBvn5F6zQa6WqGHy/Iq7/FaCsl0IdLEKUOhGBBetdxwlJonoZhP
XtF/x4cn3Tk41fwE8YF+XKc/AGCaiXJGFAVgQTnjcErCKnsMhEAlV21TS5GAtpPT
JIm89heD0IqHEVJ4+OzhB8pB+ymFEY5EvjH1CuuUQs0CdqUawxfIFaiFJH0G4QrF
Wj5HvlMNPsDkumzXno1PIiIJzgOkjGCIx5NYB2w84HsLHk3LbUgbG0i787uvgOX4
zuonz5JhPgIXGAhM8sQd+kwlV/ElmkqViuwjuSJU/NGLZ8UqGTWJP/7H/GEU1AvD
VrS9OIoT6Fl8jhEo0Y/mZ8YtJQCLyImXdgMVuRgU8jJEGpuKJCP0XAVrUYjqrwLl
8JeWrtKyIfSMlJzBgg8Zz8A7ex9DQOL3GcFoOkodY7YOKO9OvncdYUqwb7uYk0r0
C+NMfQd28OGkhVexzQ59Dl3GLrzXDEhwBGFiiJgkXgROwRMf/A81GnqdaChx39mS
PcMgl6evs6mUhDTQ1vtOjpn2apd3qv/FF2eW9hqkcH5tKrMUWxyF6pWNGatINhDA
s56a5dyJpnOXPOWXpASnyAvBpY7AduVhskqn6bvErBcmCa53EQVZi9acfjZxHfMF
scfuk8zvsMuhH98RptdPB8zcVSTzGn21NPxp5zHLBqkelGxB3dYt1FoeblHW49re
10f+nfiB83z4OYkZ1qp+R8Mso5/bD186Rn++CrENI1abfoGpGVpxU9LqFvAN22F0
1htv4EDBoWiLhvKABmBUpA==
`protect END_PROTECTED
