`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYsVbcrTfgUxurfbadi/XVI/hsAtfjtc9/2S6Bso58Fub6fYkLPVr2YSFrSZTONs
VLSzpztuAHHm+As7Ac2I6c9ratlaD4OlM7sXg+dai/yATG/KOoh5DNwG+y+dmWaB
KvGUPJqp9rI3LdFoQ7uNkN5X4GcoPzFdIbX3V381nZfUCZyGJvclBfStfLMy5WwN
g6pyujU0JTsPmU+A+ytuYcdYTyZxnbniF/7J4DGTW4Ed/qPxxbMC1ixnB5dX3hxU
WQ6uwo4bEOplOZpwN22kUwA5XEoZ+0xm9BfNXhBWiS49GK+eux1ysuZMPT0U3IyC
sY+0mbRhBWRyGX4OZuSXFkd3OlSdR6+fP1D3gdHz9eLqaW8Pz1LJjdzn46TN8ZIH
nJLZl7nVab/Xaxu+ehgU6uleyKsHVuF04zfcexYuSRY1oRQUMY/x+fPQCrXYn3aC
r9oOkTeLP5U1W2iEqmFn1svOi5PexlOZk4Ghbg/0OuJu2ZSBjXZvC74o4sOaMPid
jWWwXCHAoyDw/uDs5BJcOeD8N2MZj2jx+9znhqGgmB2cIY3lHlseLs0N9prv1kVj
+vZbBwSmZ1N8D8ovQqifAYUoU4Eal8UUN7BuPuXHJ9E4JQ4Nh+CXNXFtY+fXfIV2
za/kDr0E3Z3iYPKK3x0v1KcV/uK9GJWf1Dr1mBjqpcO2C98AENFYH78Fj6YSFRdW
IHeKE3a9zrdwoDaCmDmpWQqggo8dA2QfZyV3GwA0pnCe14bkGObIcJueOS9XzKdn
C1uEyDpGW4LjRXUDa2tIbI/pva3cG1w0x2ymWcb/BmD8wx9YG0P3x/uDXy9g7iWZ
/8P0xqL7D5KUTgrzL43QhhIaa0G9Gf+JOw64Wjf6LfVFi6+YtCHfpfyJaJ/Q5en4
/Y6x1ht7wHywgbUHoF+RTq2qZlP5WSwnA0tKmCB00hWcQ2ZPuiR8CySWKf8kxWnJ
yHjVSPvA/D+TzTpn3C5MzTHRUdVi2UFumFFveMb/kc4eEUblg6EvoM9abucW0s68
q4Xd8bjEj8VkwS6mOyR3euy41eZPFKQYWPxZxAOyXc4mb6BN7yfi1jLDJkm7klOi
8PEecfQ03PUCYipi6pHlvakRkRXtvHNQBwrJZx9+aAeoHM2SZeHCo7lqEOSFsQhW
jU1eL51w6J/8uHLPBZBpz9Ja5O9sKXeUL5JqZXVxMY4AGemjkaPLDnUdg/SvyWlC
hmIj49gx52nNAlrAyCf9oVNWFTqivVZDzABuJGIB/TXh/nTuV9/xApgWE8fXZNsk
BnaQ9McWauADh0j2RWlqFhdGIzP5BowCUJ8LHWj0lMTVTDI3gPm3V9MxZYQkNhoA
00qR728DuDMfWfjdRfoqlM058OpW0ZWijfLU4EvpfMbe1Ni7g9eRqMgZPLr1LJJ3
krkdnVKfXX3v0tbPJD9U5tfCvDkaghR9voiymd9WIKQz+WKMc7tgGzFhDayszeI+
hijHNYf91ijId5hRyGvBmqJyWwt0H0hqod+4EQlWYUWojlqChwOpaGV8j1F4qjnG
pvhlMt7l/izjcqSjOCvYnVGgePB9PPJYAWf6pcbEMjHx9mCDrcpiaWmFl0C/48qa
b60Ef7oFYtv5V9pBmwfnGmtPoOMIMH4h1do3s/94mSnSyZychoj1/Z9cPuFkWivz
+0VuRuTcDUdew8eNY6TCwgR5vIzJDLi56uzP790oPgEsR7NM00XsM960GSRNm/6e
D8RIaOygDwBtrm6iqX820WPlHm57SnBYh3k2nnFjWnaLDga08BnasmNE/ozLBcPZ
5kvwcY9dXZTM+SLjYvHgTosVMANYretjTYgjEIZub2+T1q2stcSaVWTuWx1lp8UB
XRSnUoHPAkTP0Sgwgc4HJMACg54G9q1YFFEe1JxcUVJnBNh3fYl0R8SSYm7jexwk
nv1BzlE9vGsWqPQET05W93UCG5AbS5inQBzO34+LfC8Fj/fXVzxUApP0NHZsGRlD
X4Q43c+Kbxfl7+zufwwvrhcqtV3aLPhP3d2QyP6Qqzo5SUIR/J979i7CaRMIvXnv
4AlFgJc7/o/I5F9i3hXos787yaD7BNVIeBnhK6Sm0T2P4J2ocJ9JruFy6PQalUrp
s9iLXdY6ho8J6phAamxgKtE4ri0evnawNF8Vl6/+EEaBMiRyHTaVhoI3MjpnuWJQ
GaJEYFvsULhwuDEtXiZSuXK4pGb4yBG4J7spwCpsTVIjePDYZTACMOULeo3lGgjo
xCxN0tNvIzVxZGHvFxbeNl4ddx4BE24f+zmZ7Zq8EaFWFc1QcTegYyrCbjr/seJ6
YEqNuUu2Ra6lsGS2BpLD1tOdS1GTlmn+bcMX7tAvm81MlpT4Xnj76WhpOuX6LinM
tW2R/KAu5kDOmsLRRiFzXQ==
`protect END_PROTECTED
