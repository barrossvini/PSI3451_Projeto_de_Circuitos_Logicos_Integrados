`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VoQvlAmy8vUCNHv1NAFd6EeW1Tf4EowV5h23SuhQYmwdhhcEmvhOn1mGx81WyEYz
odEh3IB5w6dtf2AvEP+P7SPYBqd4avDc2PwEva+IBYPft4vPpm0wltB+C98u0rtn
wwuRlMW68PVLmbTnK9xt8wpiBMx6PzPFcxOggKT2+e8jcKUIdVx+Am54nL34xGLQ
FgoIp66bos0uGMYofrBlNxrVMuAxJVAFj6nL4CltBSdJO0jdI7I1+JVb2Y3LKCC4
oywoUZtxQoV+/aQ8Qy2OXHWxSpQYj0e+mef6yqnlWvqedippqwzMIkYXPGvpelra
K6igA9Ql4HXGGCQdMtnXDTvPQBLRTSxYf7yZ7+o3j5CevX1fRhkCeaC01E1LWtsC
jGakssJeoW+8WXz9lZN1D5+uqHtA9JyYJwfUGjsdn+6EwsVjEz3Izs6bhmosoTm2
bChRVeQUPJE6QeqXJCg8wtn+KwOTQGx6veznGfP+sFZp12E08bayRNERxTDYlYfO
aaOvveBGn2yp3FleMj2AhKjQ0Qp+Yg+XZMC6FLV379nlQ/tWmYdzqWJ95VH6S6Uw
IrshDTtceJG84Y/YIOMkqF+SlKBtoInNMdVvVvrn6oevrCfrQ4acIdLHYhOc3BeT
5sI1uZ7W3otx4SEGpCl5sNy8ZKqvXNMYH8mb7IPg0pMRflHy+/sxSZfEN4/cT32n
5+kLzuXjVbJkdayCDUf9pALN4lA7QV/ly9xqaMsClBY7XUWc2xxgDW4hwyFn9xQY
MFGoB1Uwh8WnC+eqUl0d1a9wogajxPhMgHW4YjY5pTAv2Z2ZE1QbFTxXoyqnJOWZ
Uj1tf4mreikXCDcqXvndYBl2wBpOxv+Sw0Web1K3h7ivmbZfqGN7krC721rToIiy
4enppF4FPI0XxQPzFd0mMMkTirkI7F+VHpNCfnIgdO/vZtCNJgiiinDQdQ3QLFBB
EkT9xZlESscck9P0bc7cy8++D7rtNFCE1zR4bdTO5OizwjX5N/ngIYKNJ76a62a7
6A6n4XUDPC8XhYd8zcz0GzsUpr8aEaIxX8lyvhOb+P+jrEMRkLpuMCy6GeU9BA5v
gONTMTRTTybyO6NS9l/2IVS0ga7Z3lbdF9lefP1wK3OquLy7bUbzIeQei/Q3qbbI
u48z0NOzgWrpzyBNv1jdx58O6W9bM0wktxczM6iu6++tJ3MWH9jBqBtNyRJlvJr8
ZyhfIGgNSu3Aln29GyrIO65jhJe8ovjcuSU8WCilrijI7X8CDXekCcuFjjI9iLVq
SgoiZUNFRxKyaP8vpqH+B6HVOOqL/BUmQQlMrWWYBTPwRsk7/jqVla6lpdGZuwm0
+8E8e5d/gmzlEKIGbhKs7OUEPpnUAF+EBO7IGl3xIB9uPd5BpEelOglGxc/baeyj
Ye6caMcZYkkIprcSSB95uT27o83s1HJGZfi5G3uTkD0jh08cNhjKvzFfYGX9W3Tc
2PD/Z3IYwCqun6LtZWdtGVeLN4Bf8XaD9kBU4WXIUc/3pG33sO3AomXAd05v8fDJ
kYh4PL2kM3+g9Xr750vLFkWnXFcKmNqaCm2zBmmpuiWnGygoqX0PtVryVgO76/7e
jcYGbv2VJSAiRioc/Lj4/rxrFRNITUZwgWRz55M/TKn+IXf/mP1YOtTUbvJZz4fi
RjZzCL11hITdwPpohRjGJJH9fqq6YVwcLCSd2p6bTp42Y1iIPYI42VXOvIQVoIfK
9cs+vQcC9Bn+KcO12OuU143gsYMqPi8N3B/FqlNt9L7TWwhY7xQGhBVgO//Tkv5a
pkNjjw7rKmtrxKCfIGPThjzITq8aTouurmNB5U0d+ev9fbSiRa7WrZ6TpF3mg1cd
cNP0JeUptJ5BJGbrxs9u/1umQdTVdWiYxdTTcGReMtfbWdVzfYsLAU01w32oa6AQ
3wsqXPTiSP0aX2zSPMzPJ/jyh0xePjZKhRJePaqDB3ye4xMi2l4QXY71TT+RVspA
kRW4uRaSlPStlqP5sY1z/7aESNVfM9r774brvTQCKvOOZ6ob3sFFUdWwKh0XRcvB
6qeM7cvMAKLTlpeygqvZe3hft/tDqOfL7Qil4JtqEdXXmAkE4g8MkL1mvqxl72cf
12IIFWR5wA5IevPoAuCwiiOb6Fih/3uEzxBz3QqBoo5wv+DzdS+NSGVmh80rNHoT
GAXoejo9m7ifP9hCMsLUxvOUchp61ZBhgoUZ4M8kfFCDcNLia19Vl+fk9T0xq82u
6kMlK99p1YO3e9VTRUUEB8C1hN6hwIXL7m3FRPIvh0RqsfBo+vgwkSYzOuiCGR1I
jiH95yD9i8fa1XRf0kVFfALmqXjLZCezxMHaS+7AsRdU1qkKTdckKuYk3xMv8aoI
O1snL8H6A9r7ACDElRkPsVDnqUGuAVLgIzguPAD2zfH3zdqx5xjT7ZXe8G9gcAUm
LTSbjrboflMlF64b+/9+kg+Hf62OgskEFc1yr1FMyQzct02DkFbjMuTbGoxJTQgW
XMZaSpxR8+gydGHfF+ESx8QDbdXbIQXK70FL999AqfVwxrtQX6XJ+kQP8r9owp1q
wztG04hijznlm0ToLAvH8AzUtCyDN1eydd4i46BOskYyK4PzQLIUPN4ldpxJdT3D
DLfk4YCykFgaWlfD0ejDMnbe9/Cub0jounod8pL1IPSGSWZpdLLDhsb1B3uMV7IP
3/z7LftyQgRm83Q6cdOh1ULvlps9XHEt41N0K310khMzs3Z+Uu6DqHchIezRiia0
6FlHu2owVcZ24R+ozh4NU6SIv5o/LXitzseUKUbBx2i8Y8u/ttj9bHoWFaNRMbaU
9LlGWtyjnEaLgdUsLmQSugHclh8ywKy8Qh7OLCRTPNUpkZT3Al4CqnXcGR4BXOXb
qBioOTuhEM+0b/PXOF2lL/zwmUOghS/qEKcjUdPXaHbZLlA3M7JRaeAXunQBLrV8
JtGIBo/2bVnCS2QbuBkJTKfvA0t9vkgHSA/ltSSS082MSFwISY78PCYxm3WnZPhY
LxsGEvsjhGTcJUbN4duZGLCW2MM+PsYq9Gn3cX+a4oLX/47Tc+QKYnyoRZXD02LO
htYqbkhtLKMw8LPzOXseorTFlpTk8pDBtAp/8/F7mzyPGXRGkLuUhd9XsyNqB+d8
Gx4Hzct8+OYvCMk1rDDU+Iqio0RjMdUAdeOClETIDXrlphUD1nC3Gan4P4qhywqk
J6HMfjHVftWIGkY9ItKWj3RPxUqe0iBZML7R9AP7LF91DJt8RvJsvXno6s3SGntS
3kSjecllpLxFCEFjT/qyUhAl/wHatXRi6awd0leGtCnn5PiEjcJwJWreVyXHfuXb
HRMkwUq751fNxq4+p/Jvop3O/5Xd5oFwoM043nu8HodIdc7XKAp2rmZ1/nz+bTOc
Zrtap54H6P39gDvQ8wyvSabEr303Uv4r/KbLrMs2HMRCUsI5raz/G7IxQZ393h6H
I+SULl2GxO4MmHMCIB2bIUZw6pgpRcx+MINGEGsh6KrmSlGdiN0qtEG/nHQCrB4y
SqdYCf2TyvIZsAFbJg7BBuk/diMBYDgQIkHF21H2hTxk6GofWqn1bpygd1EfjZD4
PfBZOcGftxTgQOSJCADVO4SxVAQoTVRqn5mf3W0HsRgkk2Fit5uSiMZtmzhCwxHH
sCBOM7Tps3Iw1+BABEsuJpndvjW/niMUB6m9DHjhpkPLHGqSWy/RFf68SCpKDTfZ
Cs0DYNjFiWVA41NCEUSQoGAaAL2A7s7tJ7B7PMP4vuT6fxaSXFo4sER27uyv2yTP
EPkkBU+ep3VAottoy3ctzMBunJzJotQYupTZejDaZdszMRJqPavE3wJuo9Kx8QWX
F8alNM5k4rtoj/te6zWB82RlbIkk9fOR58gTvGi3dI1jWlhbzHQpxK2tZbeE5oAU
9wSJNWvwrxP+mUZYdQVMtMsTCeRxbUVt3U+BobtEXXgdXWouubziHiKXx5jIfWjT
q/KDA1RGPavV7ibHRgsZk3oTElv9Rx9psvyTuz1WCPEkeidkt6oN7+7S7PMaaijj
KX3za0XJUDFpDo/xxd6WRcstWqSzZqEFngSJuFtqED2V79huQVaxfgjSGz9+TM7c
9iVZ2hL5Um4dOIU0EQ21pGryEQG/jbywfqE7VAeFpn1GjtfZj5jtpzIe9wCitAp+
g190HUXvyKi0qM/Vt2H3btcH9IqAFK0nO8s31DEKLVXWdPdzNQCXQdA2lAjRzvcb
qZYGW0i0LZHvyA85/O3WIfYyYWZ6gxYdro/JOCTBbGNdUsrb8nHZv/QU17iT2Cu4
OJCK4naRjwFf/r/O3pve1DlorN/i4pC+9xs0ifB7qEDLhyjq+ZjqBYgzE4mMgz5f
TFZG6Ijq2eSZRKnfPoq0YNRa9ApZUdi8vp2xkenRGvXrsRd8PuJ31yY9PIxmtWZC
WSUV12IDpJlIkjih6t//xzPHeNvdn8N0pc965u+7OxqXcVwM7xrLjLCAFA0l1DQj
98pJ8jTkA4c5bJVCwzmHf0BFpEqLoP4T+e98B96kYu+WiKqBH+QHiP8aaT9gRjxZ
aQNad3khZ9ARUPyI8gc8nInF97otoa5jbkWLsV/lRBRafzP+87Q2xGkqFBdOw7c2
wkCxQKuozzXAhYcGNO1ttEdLbKAZHM7UNJ/pdJ+5S1kt5p/9++E6hdYLTUxTtVBt
0Rw1nRoeoqas0z6kZt3VQ71zPRTsAca+X3JemT1OPmGRdx7rSsh6dMu6Xu1tF0B+
6G7x/x6DtFbUDpQCYeCPmnK6Xjb9snXYLcp99dF1JRupL0R6G3W8394nhaJW7Mds
at6ZBtyK8EZfLQ4Up9d1nr8YX0PuM//gHgAxT5r8At4k2bfPcLN/AJf96GXZ5D3O
fKi67jjmPtLxeXUk/vFEx5eL70PuMRmuDd317TFPydf+jgWElOT2LoDVPu5gbHje
TuqL6vUSIyEEmB0OVxf6o91Z+T05Lf4Dhgl32UH0NfyaYg+jr4DfgLI5e5dpbNEr
Q7sqKxN9a9Uw/UsJFCZDUhmo+X1F6gnFf13xDyUYcll6Sh9xLxJen7UKZP8tWwRS
pyk+eInVDg7YA+vcQnlW1i1CsR3WPYPZmJxbU6Cgo1i47z8sljRxr/48Z/PxGpp2
/FmfuD1kfXHFQ4MHZCEA9AnRe4f16/N3GGnDpzKUfj1Lwy9GY3ZcFcT8R4W+fOE6
mWLH7nVg//2eULV6hITZ7UFTPVZtrmibH5yougFkm8AW/if79zKVhhG7rNy078NT
GY6We12N/2+rOX8gmAHG0gLJ1SxGxlTKnPKmlCUF7MVNFRqIFZJqD+fIhqg7+PWm
Q5YfkxhF4CjOXrIyrdBNwRuggJJkHcS4s4gA9Gxy2KOkaKQE4QbrZTrYAvrOcZQz
Vlssjwu+g4vyysrGtUmlF8d2562aKL5NV1Ynq5EHTtnhSpILgEkDNgx7/xWkqtAI
syHU90krik2ql8eriaVnDr7w80APDfzG14QXI1bZ90+be0zxCirKC9J2QTxudDFD
xIUkrZrg81czQUBwZTepYRePAPUZjG+FYF+7txKmlarb81XbhxnWIkLyo7z6iGzy
6CWiQg+4XMEBqbdOz8DRk34u31D9gZficZOWJySEkn+UN1Z/eJX8pIEibVNOpJPj
KW5Je+j5eBCNG/Wjw1KqMekIEZ6FsXxunhKG5j4Rjm8WsxeHy4mWdt67CujU3LWm
YWOdiQVsuE47fCQkLqUHPOTUSZCBuFyEzlHh5Ra8HrGr/72AXQSZeId/l9Kei6OU
Yvgt+hdKAU+hfUZ8WjlgQQxpH0O3RLTpeUDPzVtNP3K+5U+Kq2gJh60YMyBOWzZe
GvmbL4/AqAVp78Rd74WokA69tlz2ToseHEeiyUTJL5WK9B67ZOMfkbmVwQjEp+7t
O1nLbXVzFNEdzbzo9JJ/gi4imh5PFqlVPiPpVvQkN8wJTZdB4k7Zadoi10mFYrQk
gR9RHm8+3kAhJbHxN2lrK2vW0wd9AHSx8OITN/71RlcBT5lSTDIHRbKeZtP1hccj
NZRufL9gt9/ZpFcKB3x0VfWd0r50Jstq5nnV5glSNo3zJcmqGbSPoy0i6mL6Zy0Y
9lXeiUC5+7Ngzh5hDDuLdxjoJTYoM/GJjCkow56z8WaA/xwZcRpQsL+P0pgYJFof
SZFQ2GhTHw9D/K4HAk2MX2KZ5Dwi1OFn1tvLTUcySzmJn5sm3ODf7I9O/bT9LoG3
2g/B0QrRkV7wvWz0gzpySk5L4bDcXiiZwWX2lMXgQflCMiglNdrBOvWLEfNpcFz2
uQPb62PmiQNdcgcfGAn/+sokOkDv4nvKDYWJgObzKDc89Uwptgt9jso0z5JYFLU/
sbMSsbudBNb+TPZlAonDIgHCCl7RfT7AxcEQsou8ncXerMa7R4gZb0mNEIM5QbVG
rnYMiJJ/B7tHe1AfRIDciLuu4JjSreQvGOJ9ic24Pw2CXVZ6LU+AvJAWb02X8NlA
4TQDkrHM4qNxveCWWX/gi1TVAXE4oeAh3rLDJJwTtHjtgRKwJg1UgY1uQ8kMk9r7
PS4V8+IEmdUmpbDHkqF57Haskln/mKORQZJXQ/lktF/XWC7Y1bedM5v/LoHqTIKO
z9nGcmnGPNS+3BJGCCmwnjT3O8DAP+ER12cEr9NJnI99knf0uoT4/yldUbdfJ1qy
W/NAMxJtTm6wK3YmXlHkkDu5CdtV/LCklaeHObhE3Ic6n2K3RueIeqCKgUYXH1E4
CvNAXtorWVa4WhG6zkSMblrWeC73TTbKu1x38fwnhdzyGk2wGmduUxr75i92DeME
G9zqsz4aVuic3AQiZLneMl2kPMB7/LtVqSlJxBpOeUJM+4KWh7DWgsRPc/nY6Tjv
eMB1i2+UntdgUTDApshhiz9enwZk1l7othyAxI1N+iQugs2CL5Vq105QGyjbJw5X
qj72e+57v6VHf6JMuUrQgBoRRc/RRt5NqtV+nD7j2DULot6qvKQd7oG1QwPY/4EP
xQYCaQytiRLcyH8M5zcTXMAR/E66tD+GgkT+3LBc9YOb+KxULK5zjyH4qQFXU9NU
nouCQAS0oKD0pfK0j/7qqutwqczDluAv60OQyfk1y+mRLJOrbphUnXhlQ+AKHPi/
VuRxVoWq1CHUt6t2Fai3hyDT4RX1vEBKkblm66VrRBaHZ/fmX+uBuJZdxHg7g8zM
2e7j7Mra8BKhFXbCVQFHVwWoYHOtWpU00ph/0jVR/2nm6y1LFzh7ZEfN7OuImBKe
EKJGxQVOavi2ULYQAGSeCQdoLYql12XC9GjKDgqDO50rBnIFiXiDwudyhHWJy9HX
+NFkR28b9/GWTHkOGrA04CN53sqs3bRGYvP0bIpnNSFoeziEA/VAA+jFKoKYzsh0
QZkMfoHrTdIiG9kNM+rL66BzS7Nf0eO7EV2wEXb8aML4p8Lj7Iy5WWTcSPPaJYkr
rZ0Mwj5tku/oHyd6I60yaRkfAw0atUxfPWbqGXIt9c2/8ypbCBE31BDwZQ/Rud6x
Gxc8OXt35Pysv44biiLSjjt8tAVscO7kwnOCbrhahLO1hCh+IfjgySjXbWA/oIdN
V/OFUCJF2SUgsT9zYgwa0/l58hraKxmmgPwiHx+hpYFHWwJAUX3nveQXgu9uKVhF
AhKLE/OmzVFgVyL8jl8/cYGkCwt9dxKu0Ek8RukMx+8OGt6UEHGCNCrfmgYLo1uC
DQcjssCry/+1IAjryWSWA9n3X0FtYZYoc5ENvuUmbF83WJCtnvWT9gxvXudDmKUO
bZUgQicYxSJnbyJXft4QX3cC0YLenpSDskdxwtwJj6+t/vEIRgbuxgXwry/czqCr
lYB0C/bA8HHJFjif+XR8HwAIQqz0z1IpzeLaN0VKoy2w8n3hm/NZt8twyX7ihok3
WnUQ2pbeE9MxedHXS2djaGpXnfTOEc9iG33Bu+72+dN0frzz7dyGnN2L0TmA8HAi
JfPNNulU+8YkpZ9zVdq+Q6OGkOCUUKMkFA/tqNJsuoghDw9TDSxMrFr/CEYi2QAf
Q/q4sACwEPy7vhVC1vuJ1SkLFtHvSKFSKbesMzQYV/FHINhB9SKXNSUrjBUkP1H8
tBUeeoUbibb05obFPbTZj+TeRLx/dx+eiO2DW73QBKJKnwVGe48k4yLhQNRQt8Sm
y2NEfKusK2ANXggUMyL0qEo2U/vWO/NPhG9nXFYb8kMRFYZi2SfXT8/YTQdR5E1I
NlcjMQ0JwAaheNBDJ7nia0UsTS89V/fwK52Uev08zOcdbqsXjLw1TkSS3q5p1tEQ
DZOpYJJ6FfXgcnG7n/yQhdzNJobcBl0BQS9T2KHT9tiXh9r7g1trFzLvhGvwYPIc
NAod8DooZWaKOG6lU2b8jAdmw+Qhubicfxpo8Xc+tLZeH26e4qc31Il9scW1eUjz
o+5zq0Rwk0bOPRCwxsvP2U7izLO0QOwwlI1G2iKPP1FQfx88hSPt/WRj0zQVnilm
0LHoC+gu+3eKQW0CRE1d9DAEc6bKuydXiFNjIWwS9pypnbwE1EIKSyOkBgWSFHSP
KaR8dEPXyZS4dPwkrvQ5u0DqDtMK1O69xxmWBovm80zt21wExY2oiUuUwB9yslXV
aqKKAAsozcJW6PYrVGhb1CSux6Avrl4i7qjuoy2c1eSKC+GgPEMQas7A37E0OauJ
bMktylX+TyEhPiTOAGPmuCfAGzQqXzRzhboFHx/6ONkWhoBztRoCIU4Ri8tV/6OC
MCkm53FO1Abfu9lSAuULBU08kTSymaXteB9iVVyCfRbe8/xI+9/Nfko1P1+A7X5s
4y0kw3ENqr/Q5WBH1YMfSV5GmpxvGIDXJv8ub0UcwwB1hhJ4KTyCAZNHcFqGVQqR
RDWdb/PKyj86tvadJVLk2VWmcZqAES5uAdZZcgf5X6IDLO6kfyonJgZpeUEneJfa
OhtJ3vz6T7bNZ+wRHPGBtRbQmQ+issuCMP/zhombYAHkYvXujTDKaEZwxBQWWbce
AlH1gACTLjEB4I06zIGxSvHjuyZTZSwaICpDGB7mJCIpVEsmkbW9uBdkf8hoRh9F
ktQeXB5z0I5qzpb0RZwtlQAKYp5OpegxDKYnqnFs2TDORGrjlpQr8vFAXIsx0Poh
JwaHRQLVCmIGWXPr/JSu0yiHLHsXfXPcAQJTW9bmpiKUusqDzLkLCenodUuY+VSh
Ft4aIixMzktekIb4VudQUyywFT1zYrozRyKM9+fV9EH+1lg0syg6kehKFP5Y/6o+
+VDD8wdIDrKNQ3OysmfGy3o1aksduMCF57m4UHfnc1GQLD9R32xlkSdws+vUsBEe
RP6pL8UCIXwDSWNpc1ez691PS+WK68z3b37wui6Xq32+mQLjYvPaMUPDtrEE1PYx
l+Sb1q76QdDIeJhltzPjfgTMgEVXXwAst2f96lC7Po17hRs7jV1kOLAYTXS30gQF
1nfWlMjb4ykpdzRC9F8WtIoMrG7LRFdYHFdd22Ijar/uyPPZmfZ9cTtU8r4MaaQD
PxMCcF3B+d+EdTIdywIoZ26D1WK1I3mKDY9RFpv0xtme8I3yrgpL6/QlTjCGNgNl
x5i9Y6LxpAEht8Gd5TlWerMr/GGYkouvPILL9O1LCy1g0OIGcHTLU4Ph8gqPRD0Y
n3qrk7OpTzvWocRJcIOVLnvy57orlJr9K+i96u0xyr8gmLz09I/BIP/NsIuSAbQf
n2N18WXb3OPWtagAlMxh1wJpAezOAhVqDUXgM6Zgr63qDXGa4zZsENc75fm3kYIg
ed15GGsM00sbd+tJnoSC/CeAFLqskafk0K//KKoa22/kHpol4nopTYe91aCu7U30
4fTq8wl3RDjbRcFMOxyL8NrJHAVX3D0XGov4h0GtWKXvROW7UIac4Cdc7PMBKMLR
sY8s6FPJyCJEC9T8xwlOQlULw+xmG58qrv9If/VK8Fdf3B33Aun5aaj6261R1/MI
2/3qq9Cwr1ObjPbJ766s9RgMY0FGhrMrgInvhPgW2s6dJNILYBtVu1Tj8G0uDdtQ
8oXFXwLgFpj0jPQbwLyrRmqnzDNSS+kzv/1prAFFOX7ZgaWVyVnvC/ezsapSrdy3
tfrv4JsovZ+tOUTPaQ1W6ZLhgxgYONfUVEeEaObEo6OqGKSkqr8OZVO72hrzoT7W
pAuEu15raYuoPdWi0bWIzvl1JJi82/cjAu0B2M0RBim1bYzsQU1rSDLSjsV1CQC9
kCnAH6dg9DBe9leL+1EaBFiyjB/L09mU2dyqxWYSrJ/bXViB6U+RDYrynVNctZWB
RgG9Gf9mmkCdVnkVyqCutc+bLpK+p6vVdY/MWtmsIt9DYsj6HBVTk+ZIn151oyKy
fYkUjEhFZ4Vsyy64f34D6L8K+NKzzN36JQ5yfxdhh5WeOhdPnTBKcnc7bXHQHhqf
wp5iG4xgjB87iwSloS6gaqphabkLJvF0XdQhsv1KJ60XK5rh0cl1zH9neQaWjAeX
laLoc9gy8KIOdqkX6oh8eEjtsCViuAdeRNxgEa1LmlFqCEDWr2Ty4yAoxBAzVW/N
Po+fBvCqAGtLnA10xXXIul2HVr1fen+qRMRdYMXUvIiKG+9XgkHCw7Yb//k90Pc2
ZJz+/4n2VLLagOXAlPJaVi0FNakMcSDwVtENedzZ1E4AYG5qIziausnMTXvtg21A
0XjW34vBxXrSFNxoVtXlquByQOEK8E4QQsS2p7x6I1N52J0AqlKaT7b1SZKpCfZt
Xem6qRAR0OSlbut+jFQ5o6yygshXJc/+uoOf1EjgDSRldES+fpKA0vUatN91r4oK
5hlJY9Hj1dleOV7rTnWhfR/lpWo2GwNMN7kgqBlb8jfiqnWYVJ3AEPogjrVXJgJ1
Q3GSepW+S9ySuansGuc8HihA1VnFIxN/nOtricJEA3OtTIHimZM+Icl8f4EQRKFh
MGHXkRdXoqlpB79C9hsEQUdXFiEC/6dOMeFJcHNdUC99us99fRJyGjb3ld1OjZca
8grBo6NqzAsn6g/RILN4UDvIK96DyWrKcwHdFyB+r2ou2qTQ4q91kdL4JiftI7AF
FuxudQylCQ0xabyMf3l6ErLrfih8lRlRmimlq/nt1zykV5EW6DaVZwd3UTIgCQUw
iMvFRN1Pk2AVWMYdwXw6waAzXrMhpt+tagW2QkEicG1fh1VNDcPkoK0RcIiPlFk4
LXuIdYHmtsdWvdqdw4PS04eteh7g1Lzrxd2Ye4g3euCK6azLfahdOPjtlC90x4MS
BjnCSbK+uM+yCcVpw6lz4pteEAeqI7yRCxCf7C7imTuA8aTMbLdo6J8Na17BY9Z5
aUVH2Jcd4lmKVMV9hb9vRycHeBCyImGDR9JTX1ap8byJzlnS9GXryodtTMyDdOoE
xvcI7MufQKV9VDyP+ubhNNw3USph6HAkU5p9R9N6h6dYcwk0fsYNtY9khLm8GCes
/+mKeuE/UTG/4CbsI8kzClBPLEmjPDKtarWyC4I8f3qXlPw3FVjiEEHRhfRJJcKu
8TqXbRzp8rmH2yVIizxFW7Tl0eE/qW/pIjCde04TrjjX9S7Ha4wkWy2d2uO32PUg
ND0/e4airwh0bsOXj4KLDiTgZGQzID9OJ7arT/UMC2f3syInSJi8GP3+UqQG5t7Q
vZNW+xyHRKZ0aUMUqPqq8s26XV6Sl/MEjb7RKQEEWOSRte6KZuv2n+wfdy87IFNd
IOmtvGdJCIN+Rlx9pmMjE4K/dC17FdXgWazp5bGpeYia48fHeJMRF1mdtmIqroo3
DJEp3AFLL4trM49X27o8y0vBbEJlcDpX4UDS2P7DdZIw2E9fg0BSFOui4ywCpS33
ffh9f+1VKsNmglXDkcl8kEk+VjK9RiNtKRypxKn06s4Uk0NejATmvLlZoVhIxT16
Fpmo24/CHRfUWHgjOz+mLkHvQe6BrP9vna4bvYgl97nrj472BVs4rDEhQul1l1gW
wb18teeyjcTXG6V/qs1l1EnmL0YMAV5zYepRhuyeCFzTKkO2Ma4DRbUabxpOnhz3
qcOMGM8wwpz8xCSqA3O9VwJANN+ytW+k9pjtsfIxJC4UK8WJgGJjJGMMdxyUvioX
hCyko9yQOMmqj48Yr9G7gJh0Q6EJ8SWisUPWgsAoEyBeNYNDaVcPpgTm1/YfjSsx
0x0GrSyXdr6T7gPO7YvUTnXpf44Mjplk3I5de19DZ7ernyU7qhoZAorypNI385rY
R0F3gOBL0QUbr/Eik4VufU7wFIn0j0ZAyKST13Ixhpz5ePAbaySVOJFj2LJrorEM
nvnfZzaeixRjDDVoFtdQ8DgXwwZ2i0dhJLCwN6yi9imZ2zKYnpe0Qf0zuVbJy2b0
H4VgjSgeYtJ+9WpLkxJdb8W4iNdmvCPSYns3bGpt5rmXafsP7B3AErlAMaokMOze
2JcScG83ZeER2GZni6MSBsg0/H4ncSjYJSfemyHazH9J76GmtFmU9B1JMDeeiF4O
rXQkB3enrjf+NRhgJVJMUMKLWB3FMeh97sBl3eqSZWXBvlbx661eUghefkzvkqZk
6XeuwcXHy840xUNLTlsWhhu84cN/rgKGcI6HmlOSa+nBHdshyheQrFww/TfuGhgz
e5kulk9E7Q8zj1jIEO1FrFmfnsJ9hxqDoJCpMZLN3Cnu3DTcjvpUfaq3fqjYsiqY
wecSBDdW/VYCui4YLJ/cV3WcAVx2kTqsnkfgLZTY6TXA/9O0ENbbAJd3Uxr58F1Y
Izm0Djal9smGePH2Ye0fSs+em/mulFpnaovH0qxn5c555LiP3Mv8ustY+QgKMckG
RzCvUD3oFPDUUnjnPG+JLpRSQWLdQ4jRG6/2gAK+R46aJ5jw//aBZj883dvJzIsk
LdhpP0eobMGsth0LueKCTW/ZVvjy6DrJqaSFOYIvRDBd4jyg3XbTYYxQERpAfScC
xb3ubAE83MbkehBC95CrfrsApbePIpSZqP+YbXtOuvYNsPXbbfwhULvD7xn8dsaH
I2frRXqBYsFSDEwQzD767qVl+wcQqJNhu3FHqxLMmiNxF8rJsD4gVXvNb/JbrAHu
EKaUF9HApv2Moh4CFetBswBeyNxMxf3fPeb3qf/Ek2tWIaEYs0+J2BjAPaOQrRl7
V0BkgOs6HdIKKWcjzrhDqomFVuAecAxpCbZOizS/MvtHJO/JBtzmrNv4Jzzo5Y4V
fgr/bHVZ14JvTX+7aonRFO+UnlJxIf/XfLeMPOf+0EL1qLym3CRLtLxAf6OSUMq+
9PtsKKvPqK9ebUHffRaiChjuxW0r4biQ5ZcJOai+sLvP6XcYZddmS2A4yifFylXf
K80wEq4JGe9FAmWq7ijVWSXNUpQ55CbGo0pCTKN6I8e85rn0E0aje2VEvzuC1G/P
0WSxr+1BPpvMANZD2siKPfUOf/nMJKpqgxVoVDagWE2kT6W2IoUGKYCUgz3/5LPi
mwG92eWhKlSPZRNZl0B0GdylXdZLrnhUFvFdMYUcIBGchAOsWeZnhWy0RMCQ3GR4
WlUE11ufxEmTzzQYT0EnbmWkGK1tYHvX0VY2GUTUytTSL2022fS3YyubhnZG2gt+
VSxdfpAMoZ4EJz22v/StCElR/zgo782R8CGBEDUR/mSaejnmkPU8AyzGxswc7tuR
F0VDo+7ysWi6sfA4znaUIE7t8ibmU+oY/P83CFqf21COQ+L7oqTk1yUivJCa0d2E
/ue/nPpEdSTE9l+8hPo8fs1Bkw7ZEx5b9LdRbCSQkHH1msY+xNGSX3WFzZSQ+82K
Y70Pt3kG1O5f2V7Doww9iClqdsnRKzM1DoH4VM8GMA9fwTwwEF7VQG4f5+9Bj+Sp
bps29rxBV97SD/OWBsgMiBPiw4RkMSJRbomsmEXcLMgtPOkqYW1OtDRL67WWFlFi
2pmxxKhkXhrOUUboRuMEtKtvvePHivFxg9AoujZEkmV2DLBzsudGE87J8bq9MKCr
wG8Njy64qMifG00eReyzuePAMBEmiNQtG3qacCgN2RTFDYGRjEzIbltsJUbqRNX5
WK7OdqcWlriKQ+8rSPhUFi/9AtLAPtZ0mlEpS2wwEh3hiWx2C4zXqCnxH1pQtoYy
xABE4j3PEehJnQFbWCcvAF2+8A/zUwDn4QugAR8m7iNrxKVWGV5BisoaUZWa5v2m
c1e5JYrda+huEZc+ar7Gz4mQaEiViNPxF4is9EpnIXXVjx8g4SewVBZZHP2y3AR/
UIKv+2BJv2yZ5E6EkLkOL7ibXUbhdr6knJCZak6XJFraIc7CJ4lb4r/V1F8IIMsR
72s99vaLbqacqiFdgQDHGk2U+RgRpAol1lYPGGzRw2iNih5FviSkrQpTkno/5ui8
kJIRidko8T1y04ddiMYtxqOz6RKz+qSvo5EQXVhy+1zZyPL98vK/eTX/cxuyNbuf
b9QjFkumOcSNGDAV1/TbXmiqInBFuTAJqQJxYczs9hONp1z/TYBHYKPRmXF7CYrJ
oelpFlB0kvb5kthueKrDq9oOlehxwg/MvYb7OOxZuUNejrn/+n85/Yfbt7/q9XiS
zN9Zcu012a4J4j6iDFOKbqITJYHZ3ZcFAworVhF/FMLeeCRV/Lsxs0dg5XNW2UYG
iy/kLTfueJqJIgaY+lUbh6vNleWYxNXHIYvUGfTozn1Zve7aQDFAO4UDa6Z+JVkC
43ryntV+t3FWn6S+hZM149YeStVI1LIHBenxp8PADd9Zyb8AwS3tTqGKvzMfX4TZ
bosrI76t3+pFrUIVUe/T359bJD3OA3Tt7kwYsVEl1g+Ty7HU+7rzBgLP1zuljnDI
i+lenzFnwHTm/5DFjOBHGomI6ZaQXhp9WTfN4TETc1TqIr801EMuR+86vaLuCgVE
04/Rho6rgE03l8+uVIbw92K3Bo7CyBmESOodwbbuB33EkNHUpeutKtjx+wgk6OEL
qCTNvG8kTdthGGv0nxLdV3cH0ab+zEPR9Wth1l6eTUAR48oCpXLJ0W+qFBt6OX3A
EKp0unNlGK8982XKfwsntJXDh5Vh7HxMTOwO47YxuS9ke3Iwx6PyaczlwUYBWBIo
Vcllg9HPVduDeuoRIe15jlZd9NpL3Ka2OTzsjgBI0zbmu5SdiyXkiTvUevLSHatc
3mHNxuxavybNnIAidkMr0YRoXEqmeakdpXiiG1EuvXh493xZitQbErtqMFXwb7VC
0ZhZNDZx6rzKkFp5QigYY9LyUaF3nL62jz1SG4kXEhUgsda4j/XCxfMgKqIFc7/c
b5NzQv8vSc6dFAj/xNC1g8vjedpZAqiPvm324BB90o6YOsIbsxROY+rKAqHTzswX
w5uCWUmvYXbJC97fu7AIfuiDJXz7PTGNjj/3Fqsr7ifIuT1U9GVdja+CV338YQ05
ntnkEhC9SlkBkq59cFm8JSAa++7Ob4cvz6OST68JGGIHXSsbfxPyYLb0LrN2KQtL
Na9n3kBJmZs3D1rfZUSt8oREok7MxYMgwfWUssesNrNp/YL0M2ktDkwc/Zpo+3Ri
jzZ3hUhKrzJIlCbtHA/dAy5Y7Tx04Hd8sS1cc1l+rY4CxrnKi+eWj1ob7OQgr+/L
fqcAniTQHRkj5Dw0NMZ70xNWiyGA3YT2euzH1gZRZeIFPAQVuHKsDP+DnNm9RR6W
lDF3HWuWDkbr1BQwqc4S+dsJSCoAJ1iTEMtzUwmGV9K60Fz6g09f5f9edB5RMZOq
WaWvdr+nxj7hnE7WaAhxbAzXuqWqYQlqPSknLXwb2/WRMb26hQnPUwESaQW4Qckh
pIfvrEtXAjgmGkH52ME0S+PbVZ7wq658RUA2VHMARMbw2FJ+ZOD1lHtVp9Fce75S
PdZthBA9CU+/hOuMdpEuz39pH8cJtIz6TKHdlStG0cMhe5nPeKF4bKTjUuY2jhZy
RS2PgOsBlNA+N5gtOj8f9RBotijfvK6Wp4Jktx+HWsbdooPZH/HKsM1UYK1FYyb3
N6oSqtRQI2fMyGVDIl3bHMtreRtZydEyf8wCh+mv+CKBE3MdDWUoc7DpcpEC2WzD
MKDKPdACixppAne0FgpvOUUbYSyxjm7W7LWn4fGgd8IKbKKg2bOMoxMwViBKqBuk
KfthX5s0QejuKTORQBTJzYrL4kmOgq9EfdWh556K6RqviV0ibY4l04ldqyLuzMcE
0y94cI8UniNwvj5mgoAvAv/t4NK0rLYr7ifeevu4caH1qV3bfJ6HTFyDzn4e5ggu
S9wgL3Ki3i9xwPzF0KuJ1eknpsVrmtLwisGtB8f509Br1aDaNvkDTZ6JI0PJlgf7
KSEzhHWNJ59Nm46mtAOt2vMHDan78PcwdyD7c2GUihP2ga5onXK2Obl3Rt5qi70i
CAIzs0jjnq+LXnvddrUQM+feuVXYnIb3frCOf2tga8KkUoKWbdbdR5lX4PAmlrQ7
Gn5FFNMeO3MRLY3b77V9tyOPLaXyCjlo3TBHRkOR4AhIC5g+nMVj8tl1nbhD3awN
IlRyH1l/xPZt6KohpsGWCJB5NGV2sAQvsW+JLm3SHDE+cQ29K2VEoCXnk0y9S25G
NS8PHnSFrPx0o+9ZW/W+W85C7eT+elTx0nvHXfs+jPQimnwpkeu1WpeF2fQ7nYhI
5K707BIpvGeAtiLkMWqf+jwvTMXWHliZ6Ozl3B96qKGHObt93s0xbuJ23klOzS5L
xujI1Vrbo2q/fAv9Tk4VsS4tUcmh2b2pWPmtrmiRdVJIfyYb6C42+xrNtxgXjsUQ
t89mrNcg5GRQk5pqb4g/375+HC02tugRfmmshd5LigUjvzw6QtUwZzP9Zr5PPiN5
ZMXBV+mu0mPGdUT7fXsA7ArVQ0K5ECszOUtbi9X22Bn/Md65HMHwX8fWfaT8oHaw
piTlN/1Sc9b8qBY08ifesbWr4lYy9DY9h++6o+82ftwW1GmCxy0zaXt1JwwrXvZj
D5Qmj23l4YqdffswVuCr5HXjx1brzCMC46JX7rrETgGkLSGXqjaDRFGrWjngIJkN
r37eHUIKneo1RL/qCFQ1Cl/PKrWMn7wOe1yAzePwnGkmjIANXC2WVAum6/6RmZCf
Qx8CRIPfFrqRR41/3jKRPcPFSaLw6dprnbnJ8q2w0/p6GPjZgyJgT1LeGgtq/IpP
lX88esgtDznDn9ydJmEACZIVaePl8+94jVC4la00e9McUdpN7B9nU+lAWM1aBssx
6JRZo4Hy3hvgXktAYJsB9fwST2fMCGOa7u1uwKhgt5lnrUC3UYmBIWzmUmsGGpXR
2/6bnqV0h4/U2jfpgilnmUO9R52YJlTug0tBoZLYDm/C/r7DoedwyqmOS4KQgN5V
nuhX4As6xM7A9F2CG23CfZVehQDnD4/tPDDoL4seY9U/RuMoXgk+PGS05eqZRrpR
f4niKIxvsPszTneLIXNOdlRLPFGIW5UahaRfT/4N55ml53KxZUj5VL4r37Xu069J
z1rqlOPXZX3SfqjLWKbEiP/gBtIvJR80IWOk6hcrLnFGFxJATTMrwohEVPtCQsLL
mCpkDTKjLcBvzSN9onGwe2bxaLk6oGEZcaPRrTJbN6g+5lV+Ee8buylpVbwN/vbJ
CDHKxPiiratVtT3w1RLtlsgSUWVp3QtBZUto/HqsE5Ze/hIOmyB6lJwj2YPSgGLn
qXvlzbVOKLFEyMfWPJ34IuPT4QjBdogWDooJixj97woMPsufGCTgbF5+Rkbz6fb0
9IOk/17+mxrTX8a+d/s2QoRppgE0RVl5rfLUBe3w5l+D9uYzMrNMDkcVT3/kWgmg
WtTNBPW7+uYPBXa4jSnl1Bct4RDYv5BtlCJhqWMWE0pw8cW7KDoDEteD3C2cwVLq
MRoD9/CTxxO1Vhlc5TQYKzwJbPiCOMyB26OpbCzeZECDeKSEeR1/f1g4nr3BV685
UyyEPVln1ymjtwzhKVqIuIsjQ4y4Jcf71sFLuvy6KAXI6lqRLPIt+3hBRqsTb1/U
jvDFBlXFr+4pp/YkRrNotlKZ4G5TZsKQ3A/zjp0Gz5FKXX4d/3evrNWpWTLxyzf3
DEeiMMKqivmK0EsAVppVLUvRbglwzV6aOg630RkXYC5GZvCgzHQagd4wFWs6auKI
Nx+N/BjY8lgPKrAP4ap9u4zjJjbsivgd2xU8ScmlB0OPILEmwB19vQefLgMRv/JG
kRF8EsI2eEn+3WBnD5VtjWtRpTz+UpITnvGnfShVJuT8XPh7RlpP81BwwoWf9ZA5
7Jv5uwBHrnUHEf+EJB1y1PfMpCF1y503pqyg+3YV8Dq84MkuxfP9DTl7CN4rESIw
ll6vFHY7TeMnRvd09iQ02kt4F6KSza+27StNqR0d3WAiCaHmli0G61jzB05CSdHH
0zEa2dSuh6HF16sey+eSf0MLGxTGWxPzP8sYyG2V9NP3BdvVBhnxMN3wNEfJhIAh
V1iFjh9VzHanTPloR+iKXDtb9nYOuX2kcB1DpSQYuUcmv+GZlnZ5SFnn9LujY+Qo
iWkeqhfUe5+s5qcTTi53GF8gwd8BNpBG2FKMfBX7/BfJhbj2nzwzn3VuPcBka3N1
lZhcU9sKo6GNg9nSK4vbRWCmACmsT4J4aEDD5eQ0gmKHK9ox0ddF6w+ONnmnnsKd
ZXQO5DG8PICtfzBPO0H66CP8jxFcEF/1zEGmd5IYCmPjs80tWf2klLfWQjE5Ffyz
HdMo7oLJii3bxExiQQu4L5QGf2wT3BaalrE8QPp9m8mocgs8+nMGbv8R1gyNh7jI
PgAFWcNiHqVvn9JNUSVbEr2QeDcguM+tMSN7aJeiyYTyhIaL5SZ9PuGl0w1eBdKZ
c3ot0wsUgzOajVydyAyNFh69hdLGDiQRwYw3ZSUpWp6bg2e2yilXuyn6UZr+cazQ
f/AUN88wdoGWxYo0yjAYiYUK/2vpbDdV7qWClFYeZxg63jyZfCcgt3f4Mtkk2CPc
NnAgTgqflSynmA3HCPi2bQKqWfWE6SKWcLHJxfxDlxU5eHskWH9Ec2B2l3UgA4SJ
Tc7NJxGjySTbD7rB+JY+MDBoBqUs8QkhWhCAcL5kw7EimB/1Pg9Q5fPt1m4EPlw/
4EB8ZEh63I8rFY+d6djxsBt/OdWEbCAnaVHgjusSQak5tonvea70CkySR0cgp7HO
JJpM7U2RHS0QgZn1Vmv1/w8LByC+lVlO67C1FHyT/XSJEKGMLgZGRxNPTsftgWNS
v2TvLTw+81J5ZP1v19t6JUGmRJr3+KvAKcgVPWej7BTFmmPUtYqTnLCLXI8U3T2X
B5juLejuwHFA/1v6p3k79hIJpYMbEWH8tJ1wNcgZHS/Tlgxte5+Zkg4o1c9NMFLI
dAjUZA/VjONqsbFfVtPjr2w7ysV8H2SrfJVaembMDBiYL0wdKG2pvFZwC+UKV+eb
+L4DMLLyZGnHPt3YpN+Qiut32rj3S3DjvrjgKHbDvAhM94JzRlPL9MTpCH0enz1P
LFq2blr5tiQ+fG/+xDdXvM9v3aHDdm2YM1zxE5d/i/OSXtU5yZjZdk155SrykoU8
YznVBxJsfx3ej+MzoFCoy2kE0h3SR219Bm/RzYHPkQkHS4jLQTH54+YaY4Y5dITW
tRWxao9nkJy0VkOZjIOyTEwdG2Kjq+L4gktwdkAksETrmtZHPmTfLYlmWvAKChfn
1XQRbzlkFHkoE69rXfL7/xHT73f1X0vHXtsCPhLCK7Hbx5CXLhYNpBbvNIw/oO1h
7IdjqBC9MLj2WQ8AoSCV24BdjN5loYHBtj8O6FUQn85Ga2XCJOpS87R9Cx0kzVaK
FYn4T1A+7Gp03HaipAEFpZfAko/a7wqzK//Cc/pbQ20mr+hDwGo7BfBJ2Hitw6+r
FnzURgum9Z1Dd9HpOGkg2PK4xW6JjjKTBAzqH0HJCOticuGjVjP5EzcYP975NWLR
fhS8S9FTREvshHs9UJRrM8z/BQLuI02/TQOMeuZO1wdRIssuTHRyDkJg6INObpXG
W/p0VyBc70rD15jt5VhGgM+f+VLxtqN5TC/o5OCWSLd4fmkghmXvx1pfunmJFfBj
ZaSQ4AwdX2UJu8PdluLgbhaovI7j73/2vexCdACpDYTCG6fdQBuNbwbB0GH5NvCo
iTSgBbW4uJIHE3puvWL9EwtgY4AySz5VkAsFcBtV3C3TQ78Ehf7iVlugyD8d/hHd
cZcRpUg6UUD6BQMzxNAxlLJaBGB/fIX2TC34jc9qKa1jvhUsGdl3smYQVp9cdUl1
yP/+0SNJ58nnn8VMzNbSp/9TjNZ5Fwa89opqRmzRJEAPcq2K2/HFppJtV+d0YoyA
9DFNZGhgtzs7CVP7hDCaHLKMdRRY+hOsDqzTtLNzzYdz9JGQo4xqrdh2Drk/GK42
3RPlRnJhigVYzse3Cstx+TGpBnPgZOrbUXrvE20x5Tp0hDNrg+D9Rwsl3+r26Yb1
EXmAARG86j1PbRMJ7PLfRVqC4tJWyLASXV9W8c5tK1qS+CbnHPqceQecdD9h/JRO
zexSU6O+ZnSN5POGmperGiRdF0fejwWIjQ60kYnDdLnLL9yd6RgyjmRjio1OQp+0
5ALk2keWnVxkfIXSQ4NlbWX7FXXtstdZj2ifU0m5AFgvLiQ3PI1+0ipRaGLbH77o
XMyVsqMfLUVHf5/G8xSw4zTOhHU1Jp5dLDvdJ9Av5XDtCqTeiNjdyGeR7aVIqeI/
cxljHpg/zO59UM+QuJTXbIq2dR6veb8dGPxmlXVxeNa7cd1FMpX70JkMsHNHfFK1
KYbeCQ7vSRQgBK3dDHze5ckT15AqKbjg7galb5y8mmFScS8GyezcCxTYK4OYkhsQ
zCL5Gxs7fRCjPQ7GmYSenWzc3rhzzMirmkzyIFKxaQgJnR6HjCiwnD8Lgc+KFGCz
hMeTH4hwAmc9bupoRuSls89J/IVCzQNlZFD0b2VkYMhoxUoX8gG9giDAp6L0Tg1u
v/A9JQsUypCm81ARgN8535WdJAKFc0y0rD/tM4lk9z01/H8a5SBoPOYt/ZFIhtgz
HtuRbcZ0AZ0cE41gs+AkmitdPe6ahBSkBgoAdkXD0mMN6cUQnZGZ+r8AAIvBRgxJ
lPvcJ7wtAGu6r16nGtgZTbdEo5ierN+kCkt0PTiEVCAkxvx8YXTue1UxokdYRW8c
5WPemr77BLEh7I7/E1AQjgAdZAhsizi/0tyQ8inp6UmcGNCbxQHke5Aa6l0D7w62
Q78OMMxgouH7b2JFOgsxFhAQWucyLazLgxCG6iLM28bK7O6IU2ZW2SxkRnhFcbrP
+AI2RIGAbnKl+r44n1KN3RqaFfeTV8oYMqrmmM3X+8DXz3rgA6Ulynj/ImCwER/3
ch2FCM67HtP1XOn6iXEyp/ahFcpEFv8UCK3UJ7YTaUlytEvpgNv/hCf/6kQY3Es2
732a6vG/TU9mjqAg1c7zJPtjcmtDAa7lyaFzkoNhQyaR5d9EaTPaZ5n5Oio6Rj26
4mgzsGAMP6gg9EJnWUOIFvGtLf/aMXsqkFivtbX5fCDXaFtKTApZB8YaMu29jey5
Jp/Hpnix51Vva0q6hwTPgjR+AHe7dAIk7Mjwtz9XlhLHyw6uaM7gYiaEHLuMIPt4
U6Z3LVlhJYKJXhFOV0FDj7x0NJgrabPAJy3brc+1nNe4xE9Mkc9bqzUbE6lM6rFD
j8utG1OSmEjkbaiONRh9AUVJhJc3Car/puQWyb4gbEV6w5mnvSQ9iLi7E/ppYz13
nLeCYlgdYQavx6P5ChLbM9cbkUci/hntvNypfAkCCMTRNblgU7HdWCdhr9jR9sNu
GxwFxeOvnSfKfPAziWcu4jVaEEtAEKzbi23C07Fn+j1HU9yT/KY1wbL13Y4Ukpf6
bEFhYulAhAJz7I/1AlCMube5CJrxf/9/vzvvHyUfGcedXmL53awiWuxzNrfCks0V
s5yf8VEmmPgYi+1Ic6MHqoG/IJ3tNbS6hUlPsLyOWlHbeoy7lNw16+/W2kr5jK/W
VgA05L+xqO5+z0VolEPbqlP8v9jtQmcQKnX3GS4QXb9x227lDjd6oWrNS4XaOsj0
REVPn11JrXSw83cP+sO0B2/w0ors8m4i44z5SriaosJkT+DSaLTyTt6KrqBJFpBf
RFaGUnbadvqZ6ikIkLEuZt87ys9sQkGsxxLlqrug/ni9Z7EmGJG3QBPfmTMl9bYw
WvDSQTKUxCzc2SnCX3u5fTWfU/DQTERIzYlq3A8uct/uIFEtEiXN5T0NRjMbL2Uc
YBPegWdpuKeAgPf1fQZQWX6DsJeVvhxIQYY73VzdDwJzm52NFd6965dsCTFC6MQh
oWboi8RR9pToq0T3qaTyJbLsOWdsaiUNBLzqvKw1bfvRcwAlhPSfSskgwAXpcpxO
vQz+WRqC1uml3hZx1OJsHdEhr4+906ZRX0AAykv3gkmGzC+l01udt/lxrKDRSckH
XFWiSLofWJyJ71TLVX0OC/nJTHBdLy2+3W2dDGYO5bBr3UrdiOGPUr/MpCtRf4DG
7z7XhyzhNDgHwgce6QxxzNjMtTsUEv2YAagWpfXvtwww/ImVKAU0aWyTWsH43Uoo
W7vLGPYJbDtvPUu1eaAGb9Rtj+ghWg09+GT+ZlQKmleN1Dms9tTrYXaACfpKr4JR
cwmlE3v3rBhZXOJ81dUaLl0LqAQoVqKiJXKil9zf13vtKhxNAvF3B/lGMx5cpwBv
wZhPft8aylbLlpW7Xrx9pBAfigFkKY0nhyhso3IVez6VoimXh9P/HcUt+LJhT9aL
cXrUuwaypvVQy5ZzjIaTQi49mMJQa4aq/dHdQMSVfuniUeNDNu2iPK21xVyv3IfW
oQJ1M79Bz446spZazH6nFUgRJHGdV46D0gXtQPtXhYf9S6EosDx6OBn/a6cZtyLg
KLBrxAlZ8XWYFoA0Y1Q4nKfN0rTS0UgcxkBJC2I8N9fSA4G35MIFYyv21Yv00mHC
WUsW5Vu19NmmFpvdCrE+Vfdpg7xivxtsovrfU6KuBP1Ogf4yEJMZifqBrUZzAhYf
8wWYP6dOTXkSjaFAijvHCYXpijGllGA1j+nPcmSMJE+cq4w/+K32oItMsdrlppZU
Y468aWpED3t+cUS9P1EJdzDW3rjr4m3McUw2ClYgnfGjwjNyLBWTYpGO4+AHDa4P
+U65w4JIAm9i/xZ7UTV23OxzGNahkLy2AYKuQopVtYphTQFcft1i/Vp1gGhZQX11
r8wNa/sBEabvcwuxjoDkFxrHoGBT6CQCh2RLqdYB3hQveKnJE2Qn7R5aiDVWma3M
lot6vUBTF3bMmHxeALWctR0m0BS3XLxVDuptPCNd1d3XuXJbRsfG9xC3MHuLl8ZG
qhbCPlyAKdtyTnh74qNStGUcDns8VpBRhJZtkc4awlvWSDI+x+I/kj5Os7T/RLc/
iIqzOP2stnKfJ8diDVcMovyqNQ5AhR+iaR5g3ZWE/bItw3kzrp3tvCuHeXpzQAxH
gDB6hCFVB1T3Hb/Q+HOwDTZWCZvtPhp61edkH0nhmGSaxI3TnEGLbvaV+gQ0ohDe
wx0zzpqAcvnYD7QAgmOtk0BGi4tT26JMXW18JZ/0kevPdhAQxZxLOS35dcBmu//G
VERBXexMXhyPXHQzKHMSYNHymmy+I32JP3mPjUa7fe8pRo4OW9wq6bWAcI+cIBpf
Yl5030fTg18CAfxKDmnusomQEv1EANscnadIGLwuzf6XxWBv8D1IHnQO5i86PL6V
m8xEYzimUFBgGi3RgdRPv9WiMmAZ19XvV8vTZRq71LJ0DjdnMGmFHuML+xoPth74
L98HGK6p3RDFJDLS+dylSULJ4+cpi4+a6h85waBrNcNRqqYbY/XwqKtXDOxZo0pc
bbJtCxcMGK0BnD2eZgX6whWKARGC12dMFKwV0Dbbn377CDxOyFFNwBxtgconkXEw
aXLoVy4khhpNFhUb2Cag6yXv0S12s9AURNB32p4fwFSjql0xnPl6rXV54xjnKoQH
pTwqM0Ahx2iipPB3ld39OhD9PaRQKzTtWL+cN3gCQ6GIz7R7fcWVUZFzueDTWWDL
cr4ev4FuoFijwPNBJLQG5NCMvZh9WjI42rSOyWuALs9Rt5wMfjmkPd7knnwW/UH9
sffxbm4WU8vka/hS+emWrDJCxhd1uxgYS/qAhEjDAUNH/ZIMg8v9yGla2POHastN
ydV6DLITxO9yUE1uQ1VoYN0A/vVDX71lGvIj1mwN0nTWmllONLe3oM2KN+d7wIOU
bKdarWjAK+2+YdLDSj67fWlREZSRQXZNQ27WJVf2OIefhk9myZmN1g4FM96qUUD5
4uX34Nulk4ftozXDUc113k7MJFR7qHNC1MO8O42+X9Wkv10Bdiblt7P0JGdiaIcH
BywSHamE2KoQBpjlmBhnKvasYtv8OHMEB/A1ABCaSSuxgkWLjRftk100VC3tpIJ8
0RA329MHd5CB0JSYmvwIcawfsZ814WYrbfdR2tasXg+na25wlzL93vT08Q4ONZci
TMiIlLVGXntzBFSd0ifvpPK5dvZ5fT+g8wm6sWFky0lGCPObjqxKOxp+7GOvNmgW
DKYhTvJNMY7zSeQUy928oGcez0EUAKmQLNB9wcTC1cJ4K4+uCCck9w/VBTktcvzc
+Sw4te5UQecdWE6Ffpc9I647HxqUZrqyJiPaMiOAXh0lH+h2CwkylozukAulDD4G
brKhdFKbv1xw9d3qKu0Qu7k3SviKiaI9BxiqINdb+r4SngT5yWtfs31COz4SBPmU
HMw1x/jvIaFPnbP3fJqDBAhiKOStoIwScY5wUVAmE0QRvFu+Gxh2W35oTUjpD58G
9/xZNLd6Ooi1Ay1luYANU59rPRGUoxcSC1/bOoiOqXxHhiYmNkBhQteVC+O86WoJ
GmEglveZrzX4miySIdaA16qcPsHeKqFqejsrUjIlhjHIsI6voFl6UhD3OglPrEnz
V25PeEifuXY6gNuF48q9GXaXt3D+Tx54Zb2iqmULFkYLfs6s0RySLxgXNpGPEuEx
IqnHNY7K/Gucz6Ix0GkHxDOcqgeB5qP8kBtm1bra+xso9VVXxfEO8TpWZB7+M9CT
17SGd4nrDwFP3d7sTq2hyhawaOk6zz9cmolMEp7qDlHbUU+G7OnOYpJ+wJKTktjx
JsIBMUmKg7sn9jACkmoEP9OdexEk6f6M28xvgnqc3ZmOdrs+tcolyTc58w/rkXDi
ttUX65PDXni4TSQNulf5+ihknD1UKHEpj6jx2Bkjx2peSo6T+NMzkvcRn4LARKpi
f64NDUnY/QQcXtgKbLzBor+j4Is//hp/yah0O9hQisxibZsyC5l6OKEC8m/kUkdz
sjwW/gwM89dQrm8jX0LwR95GCKVffB4kqpyKZ+XheqyaZZxIF8JPGvs82mh4g8UT
Cr4Zf+m+q2w1vJagHW9y+qpx04QcAZHqKfe2azUjuoed4InZkuY71XyglA1MdEyw
ZfutmWZ6bwDsyXtpnVfnHGKWu+YMoyAzHzGSRui2hlgvnqB+eVM+LmBooFFz/VHF
PCBnBz0Lu44j57umzd4OoYpOLCKAFg/+1Go9OjzAPpa/QxIRVSBjaWLczlGLtYAz
TRCRb8bx3yUozPwAxs7+lIgcc2DTmifpx0SIefAqq6BBLNALgefARp0IjnA9Nzoh
ri+2fq+WSrDUUkBQ3pkdyAXn4TuW9ZVcRTNVEx4IGNs56yd6ETkJfPk2lyge8Ruu
zQQ0UgNqV1IdPe6FXR6KR8zGV3daZsvzxSj3lySeB/zM0t0UvqhGdriH+vtfSVoR
QlvJp5DnlcNVUGlZA4sVCsw/Z1SgJOWEz3u+BiKisKUYbnXDZ7beNSvkG2ScbFCC
NdpXKsmcPaEy6CtquZfmp4HuGdkEHWs4hP2W7cYP6Nw7Kp+Fj7X5arNY6DOhey/N
KbJSKQ8sQR9rufVrmaOh7k2JF4ACMAf/5XOlS8Mw1JVGCGbIYVo5dgyiFqVX1oR2
Nru/1lpVQ57yp1fJihlPc1abllUyeWyUvRL5hfupqkvF8YcnQM0+HjDbN1J3UH62
WoY43I0CpMeHNzcLnidW0BfFzAoYze77Q7Aaki8fXpn6OTVMPffdQBDylwUelNiF
j1IU8r9YougUoJaIKj05C1yjt3ycmuKPPcq5YnpgRNI8mt33CV4KD6yld5Pno24j
ni5IhfT3Od6GfgRs9cE+ka+0BMDVT3m6r033DqL0uRm6pWoHpG41FkGlHxW2eglx
Ng9kB7lZuQGXUbzeDhBFs891uwI+5Skcj9BVnCKaXNMwzDKYelHTOvfOTr+WSQQZ
QZhCaoi//lgpJylbhIh/aGZz8pMyF2iz5/CEqXvHDChaPQefU12QXptzuyu72xqQ
oSkDKXt4zgzUNFk+HV5P5+2wsXPsm1zwBWsHGUrfNcIdtOedcEuO7yQ3zaPAB1AQ
w+SBN2wQKWdxX/onsV3lTmkLqkGh0djOgsS1sQvCUMA6F5oHGP1Qvqh8i1fBUIx1
ZuUNnTX60h1cegiU64khZ6yh+OjFaAHrG3n+Ob1zlo2HuTKWBTWZEvx2Zzd4iySv
DBS9ZOLKuuv+5x7fiwK0yyYjyw1Tekl/YSGz/5+OZ5F+8WmzyZ2v4bjBD+Zgq3WB
1AqJYuLwxv/InLvqyjmvHM8xOZqvahQNZC0/64E7hpBh0YGjNyGfCZURZz5f6wB9
7+5d7k4dMd3Xx51yfo4qCy/F5+I0KSfpH8JJIth5EX23TtZWiFVSTlWRtpH93cRB
CFclXXP2CjGTYcKwwwSMeZFwbTqSV/48FM3VT4tsgc3eXMQ8M4VtFcUMzDPoB9MA
Gv7FZRVa0BrxKhrYmO6bQ/0I2hulDV+XMZM0Jwgz2qVm5K5/dV22zxc+M4rBTnul
A/aAHzdNnC3vGc0WMjNCQ8XXgBrPGRqOB/ENWgId+X6a9FUUXS1AyIVTbdDJqQjb
tC7BYOv8LxNnJrtDD9Z4MkkaC77bdFSIXQQtRM7NwISlAmj48p1hM1Qf2OBAxBEx
tXXVzVP5su3HaxTgPXuqdiDeo7SoZVSJUJMmWA7ybg16/p6hJY8qnJuO7LOsdTCS
5/6/7Ql+IkJv9Y7MxrvI95VR09rjeKVDyP28B+o1DbLcGQvtsU9YoB1F3N0mztC2
afCVlm29RKMZYyrRp93z7MVoHiRqyDx9m9DMkcka6e8xCXib5TP66F7Y+US885sZ
Ne7abE8NWX+IkIci36o8jHoBF7ULvKOBKogi62Jiu6o/8YXhjOBJeTc7iByLEJai
QEUyEyX0uAJnw+qr5e02Vzy60gU+Qw2ui3sWqZYIMdTQYjRSV6RS03zNOslzY90s
KC+EVYSefm0CYY+le1NGae89cm7uwbQ446Cr9o3JNHzjPl8We4uLQy6lliN2AEie
wSvVqVsdbISsvFKfGkdEMNSdkGxn/Sk8QytKYnyCRU1l77gb0QlMvvPRAp1ii5FB
aVxwuOX1mkBrtyxgBk7lb5KukJu2+k11TgTuAvY1XAUWZKrdQsxpWiK+8Q0TFilb
LQDbgqWbfCb1PQkhz3R9F+koHcv8U9NqUe1xaVuAq4d2rXJNMg+YALXpiGfEuTFV
a/tBDfFSZNNKgUtufPNDU2BDVYrHYXaV/dFqd3Yxh6+dF8fZa/v8c5mVAG7kksbZ
k8cE3MA+RvdVwXjMUm0IEs0UNgK/TOzYj7ykkL2Retjyj/16Wf4+Bpn6bfncorEi
mCS9TlZTI+xlI9P7/6R+rTIGp5WApoW2l3wSAjUGzOSpDeeWUqZDIWFl8DqdUhj4
rPbcfaDDKQ2fdOwz3+6mxKH5s8ZMC1jBZd3VDc/OH2wFDSLXOm0iXpnQl8EIyIk1
RDNEkNPAWoy4N9DO37K5/kdhPQIVRAo/ptpi3vzffE/AzaZ6ZIp1Fp+C+UDuPYlu
GiYI+CFASv64UMIMaWxD1bWK8krwLCqtE4vLi5Fr/rIZD64ELvzJummOiTQXNuDz
/MLHAdbi/6FX051ezakuYfQ3WewQ8P9qB4AV/XGikPpb4arfWykh8jBTyMxzJPky
h6EkwfKVn1gDbBhsKBA+K9MTctDePtDUGwTLkLbEL9lzkLf4ptq/P1V0M/NNige4
w6NLEWQWNMR1rOVNJERBFVERiLznCVLK09s8nFuDW5QojFzeFUlNfR7r+i+xUkHT
owNP2i8gXM0Sf2/aTK9jhKX8X23yVqEYPqO08taA4Z1KS2r1CdFjbmaBJR8lWcmX
YvI8lPllTL4mRMzSD9VaRxuhd2Ai6shbVad4XMZg79w14fEbHSluzjYADhhYKdvH
8kdP5SlPHq0hEu4I1bzikR0v1qoAx9o4XAKhYEHOkQ4AE3zt1nt1tWhVv9B4idpn
4KQr7ai6N3yUDXxBp+HuTOcewEdSPsNkDVzQioRCD6V2u1vW6edR6FpIbbsrQMKy
FRLkX3k8kFVyPNGS7CLb2ezIrf7ILBTn8mfzuTyhGO8jO8IzySycnlG6qAukUs63
cQ8AYdUe0ogwnTE9gIFrgCExtwjjXOpeXGeZ+YfKKdBVbRrE8KCs6XMCqGjl3pMd
yhsyO8uPqXtsFZAO90IcM9KSMgfvOETjeXlfEXZZs6ZHD9aH6ylPpN/UaO7nExx8
pYMQoep278p0R5YJPq16MIpNhJIW9w+dSvkZtLNPMImjKzgffoEQh/QDK++nNlnt
Xyu2Yi73Al0NOfZgh9sqDJo/hIx+Xif/8MMdEGDBW4Zzydkl+lphvVj8cHRGkmuJ
ec9rzCFFkWfOkpP5h7aJt8doEzSl/prh/3RRkhqI9MMGpSDDu6k5HTrE4zBlWDHb
ERGHAQYp9MgWC2q/p1lMBxFmn6vw+yANz9mZiqfZOJQCufPLBS75stP1cfqz48XR
VX8hPdtR9AqyPidWa0INvMB+CQ6Czsm4R+NzVhNtmPhi59vh6ShLIOsqCJKUtTmJ
zzDQZTvYo6oQ9n82bhYTW7pqeef95G+5PM/p43ZqEqLCALuVgZ/FQvUQGb8pnl3j
cc84ksXadvCcjkkhmYNiZSW2hiXlDYHYcR59z46onlnVhynT1eKfuy1ZtjyERyYg
h3jDyg5WE4qIYnenHp/lXdBWBV1Yx7rkOMShIMDrRHNYU4JHWKFxVRBwiDGnn4vO
I+8lGDwSMUHU9Yfatt77lR9cejrCACMX8G+Q8iUzb0G6aSuvwh+ngvDedpKaPrG5
KCnBAz3O+j9FV8ZYZ4W1PniLRbpZ7OvgKC7w9K4maawWS4i6h1/cKM7kVSAvHwrd
cqVkyFYoUm2KqqXhwXX6IepnLtfwNjxMH69tLnmRpYN56ZGGedFvTWX7vB9fgL55
JgMT8KepzKP8itV2+arkzfVXdAM+x4kZ4zh0uT5NghTHQjBSDx2jqST9gfq2zpKX
4ijJ6UFeUcPn6nY2MCiKRHZXlvO1BVCy43I08Cu4v5t1kXrhmc3lGzDYcd8cr3tA
PLhZ8HgEHQimTgvtOhd0f9flHvFhXJyreRCxRLyyES9yVHeTRyPClW9dpRRTBHEU
3yn6yaHYZ09A7kFtqppx19SsN8d4+Oz2aKrs/gq9PDs+AANakndE/OtSYa+hcBJw
orvIq4u9jbdOzUOyfffQ1FggX0erPhr/ocPHJb9JHuWOcfe/MyI136DlqebFQ4pi
bqkiRgJ3Z4SWO81Y+LD7zZQdGWpjkO74Ooi0o0QWXx0cD5LyIAO6Y1gaX9mYRMAT
rC+RAuayHQpZXiA9er8gnvmy9ZzbYTiu9uWuO99jzYD+dH3GiYjPmnYzMyzd+ASW
ENQUiOJXmI08sCcGNC8WgUES4ARDjnjnU6s963KwgT/tmDzj/+AuZ1SrNkMJB52/
JNbeRbIQHnFK4Gmd4X/Rsxy3c/UNYzf7XCx2neSr5C+yzun/2XS9fx8pbavv5B96
RVW8mjI377akWntF+nhFr+xjKA3K7M80iFpBC09QabBCFLtcjjDoVUPoZyiuAdI2
BHdtmPJp/cd4t30noeOecPiWSTTr98jJmTRMzrMnK0Q7nI8hGMajgox+K+fCtTu2
5iTzMoF6hiSr3p117mMAhVgIPIt8VfZQxUvvGlj1MXcuRzMS9Puaqp8lLcDW41p4
m09CUDhEbC5v66s9rjVH+hoJNuuQeO49bjmk1KAncvOdS+oy7vBJqS/4EIMdjkWJ
W0uMtJ8kz3EdPsuuuQusMOHz+UbFErx0r1pdwB3Ocq4KzRKEC4VXRBLcPKeIBjhG
S0PI5bH4dmyr6P8JBhz0HNpmBWySC+YxsuCyFkbyOJ4+5CAHYzlvSPVPlJdQAk/U
UhxG/3iiF4/h+3NRSTwRxACBOwkb+u0GRWAxQuTS+HaxIvJV7iRdPGalytsMSa5c
Rol1Bmbz67nTzbolIw9j7dDIK1w5sT7PVjJKihDb8kYOAnN1B1YmDmJyIy0qNQqj
HfCbsUbeWqzAwNWTya1hM0QE2NIijFSXzHDoGD5w0p4bir/y0dRKPsHZ+9SZer6/
gkVJUt0DPjlZB5eL1haRvxoJ9doCkCJVPw/3KQKH8RzYOaaOErnGoHI/tDloQ3St
lCrSRdm5/exbGn0rOsxUB0a/1AN+BqlCPQ3gq1OSWm7j/QPAc0K05frqFsQLHhcq
YARXxu7AgQS5Ac8WEjlrDsNwhgXUUxkaWGwoJGqOkQCRzeV03rjmUFLeVv1mXvYY
AJntK3y9JOTtoJXgy+FZ7Jp6dVwOCalnIWToVewfYWEl971CH3uXIzsi3H48IiZZ
VJwfStJq76hS8VSkwCoaU99qSzsZGNIS6L5yL+2+8AWW7UsWP242+bt+7fMDQX1T
XFILoIVG1LHdYct6sUqrxqMFcgr2lSuSdsagQ8a8Sac2HT2ayYQB2SzXivR+asBE
hKsV2ckJhJ0O3lL/zJ7/oyTRgcak60mgQjQwfWE4gAumZV37QZc0FpZRUJKq6FmK
X6ghNsvDWpzRAx4tUI0oBJTeWKB0hRqgBSu+pc4tG43iHnT0Q20ILDwU9mw+M50v
VS/tHWjRAXD9Jfnp1tJaREs6tQDxHEi0QZaqo2r400ALxwWi3Uo8h9zXudcPTzc/
LjOWgTp2nEiNXURzm45Fczt7CWVjgedM/vucFa5r7KhmhgPdcDpw7k3gC8RAK76Z
3aMf6kDvr/hILIBGpYi59a9jYayuHEsc+b8RWOBivATvwrXl9/YtnsefTXgoWhgi
XkbO7QVVIKSq95Jy7tLLi+Nan7RAI+L+M+Kem6YkNdyd8/TgVTEFIwvfYIQCOjVi
BProqk92nm73sg9AxqhVogSW9e5IR8QRJf/LldEBFvU9DswTr64y8YHSNUtPIhBT
/QktTJks3+zvrNKGWglr6K0Gkk3QR+6drKTUBVoZkc827e0739jAUZM5ZJ7sAGkO
kDh6P+mmigjD3On22FeYby3h/i8rhyG2ehHNVHGdbV6PqfomIFxYkfSe8sWjA6eu
1yVx199ibpBV5mZVWQvIpGEkc5ycEyAQyahBF/XHc9ng1xy7BE7JXq252kQnPOPa
zeYojMNez1aGcDzsOnlr0Toud/d0TW994zvdLgQeWrCVzvS1KzuMscUQEl9rK5c3
GelifjW2X6ERys+xCons2NWU5/hw4HH10gzk0FoFko0Uazligq08XeqB7xr1OlyG
NwPLAkfAEnRf4mhkQUlDBpPj7Wa1SFBMdcfTAbBF+vFC9jnI5+MRBjK3XayCUi7w
vSnl7j6CEhUPa9znQ4jVdf817TVN4THi3PNWZ+a1K54eaAbIgOJE2tPMTixx6RAU
xyqK1AClW2sV/DUJlexzqi3UGYBP505DC/CJ473CoGYbL/FWLqJmE/ghzKCZEwgx
BeaGLTYrguPpk0sTNjwuz5Y4tAPtwz71ORxVZv+c6qLpap4ChQSo3C8iS6G2cffB
Ev0a3CXiRhaSmtwWG4sodOf29fVwSQIYg06PJ9SJ60VUrBsDVIl3/SxeiZgODpqL
yZAX5XhkWLzVGetOv39Y7C9YBEKZbzN0S5FLc76096ThZGPnuQ3s7HrFaFHGGqLP
aFBl3gAmKg7h+LDglee8fV+mdsPnxFUpzQeWih1FEAxNMoIJmbO42Yoh11wgF/ZD
bhr4kWl9/I1PaArNzL6qaVtCxE21U+VxnaY7twKgUZfRl2OA/9aUlrRj5F9UoHw1
6GtOzIxByiqLM8ApURVMu3oxACE3Iu+EqFItPvYlNJFMfMSvCKctTPxQINotE4qp
GCA22AN61A+2CobCrdi50bYUfPlC+EostBAaN5c402q84fasp1YmCmvrOGwMepA/
qK/nuwbICEqJAHquDUeCU4nZXnJjPsbuq6UtjI2N/Gps2199YJ75iHNpJde5llVJ
TC5pYNJQg/ErVgWs5vprn2N1YZG7x1YPR8gcPUhG7M/zUDk1o/J777pOqfVqGPmA
7t5WihBG4z22z9D/a8NhtJpjnZAgG6lPK8t1sVdLWnqntzL7Y0EjGYCQPGnJDdQp
+EhCrjFJ7EvBy6Ee/VL1GujwPjI2+emZKKL2FDmOYYgAzsJx5H7Sdc1iWG4MJN5N
9VTrso3ZjdW1bIGfKHAxmXh5FURgdIGTiuswrjjYJTJux2n3J+XbF19iYpQpkVQz
ZSJSrZ4DBwdlk6+oHUPOWLlYBaOcOEoxBm+6pySK/actzPB39cqC2+PtYdT7ahao
qabqhCiReiWDsktFcTjUdZwjF+oymw/PMWb6rsYGNbK/P4dMGzQ7MqnEdHdUOJqt
YQO6L5wDO/8xzUzCkSYDjCJR6BhQQeBxXslUiVjT7L9rKRDkupqdVkCkT3K1ysBU
KJfcMJhmaaxKcijEBdUVDp8RLmeMME3LA9l0GpbWQVN1zYQ0Lo2bIhuST6pUN4lF
w8rCAwMC3Z6tR+GTQMax0G1/F+sSSOUMQW54mIUTzYVWMJ6zHigfyM1dkhDtTUh+
YQKgG+c1GCkkUM0Y80CUFuY9kVIuKa3zGi3Ign87rt9/S5+IIZ77bNJ2e1rzbVfw
pMEZzQG+9mHiXy/XbUZUTGBfrlGtSaOOvQGdqApkc6N7UGfUrKGJ/sCsmCty8BHt
ae2klEsZfnikzKaGax6Vou5H0y5NWC145jlAy9bfzNYaK3kLmZdoDIT8S8RY/tg7
nI2R9zgKAadaqd97rc5429gICunQ/vwSRpKmpIfOSikrILI4qiT1eCi8kP8TQarg
RuAYz31sYswD923z9/pNprE2XhCw2w0jrxYDuN7mkAY5rqaH1kFPFDPYRZ2E/5Qg
NmDPgx6LyCAFduyLvh1wT389eQc/6Ruo+lmm1iDjeJK96bjs8PnezKL17CMUOnel
9aXO1mWjn63SgiZcN4sOlTleGjTogxos6tErRo9ot96rlpQkeSgAAEc/o2YTx9Fc
FQ3YfJo7r0NnLE5tk1/bj140fNyafyXP5qL1+obXlPFtn9HBv/2KRrJy8mSTZhHX
fq/dWF2ot716KWMoZSg3buAS8kdYO/aEM9eQjsIruIkIjfanQ0Ui7Ff+Y/+dS86w
zVMmAHR4GnFt8Y4FoGKThJS1GS2F3MmCmmylSNzQVEPZ3Bhn23NGnFpb0Vs/Dzlx
1EyMjfW7KpbPB2qC9N2jnJzrXvc221V4SA2J9GO/YOyn1lvtgSGbMMzqDkXQcZPJ
jK0HVZ1Ns+j4znTLX9gZoDTuzBEpxo2WGsZe5lVPK1//PqfsQVmLlEC+FiY/qepZ
mExTdsoUwvg81NnpnhcsKnYPlYdqsScABnT4E2aq8kEpCvmVw/coi02q3pPuCBwZ
0Wfdih0pdQR8V2p4keNWZy2qsrsPiXXoY7PeGEyPf3bnHoKTggb8Zpj5Q9BEneL4
hXQalm+Pda86pS/1Vnp1rqK2qItKy+f2qbTIFgo5tOZVlq2yvIgdyM8AERcy+Gcs
fGey0INqxDjeS7T+SCL8RAC/1HT943YD5dFrjOoHD2XYVbQea17vAtDqtqGkJf6d
zK+60nI1mQXiApioPvSce24XNcz1Atd9x6Ko9tsAXTG6XnuOAPNQqAbNSxsTeuH4
pklvrDX6ar03PUy3R3rT1eQK+WqP+XoRJM/gKl5q150pr6dJ9pOYAH48mE14wwns
MjWgJf/FvbyQ7yoLlDWl8lmcWlGTixNfjmnkyHUgvQtLMsCDOAx7O2fB+1LbxQAR
Dzg8Sl61NASb6wy+ikhasrlpB00Kc3aVWEe/jXdrBYwmATz8T6+Q+AF9Wb4ayNOI
/pv/cAQrfc14c+dgFkpfVIZyk7litOram2zBp+A6Lmw8t/Fky0oyQZhgl7ob0T+j
wplbEBgsDBu8YQ1pAqGkUvwD4ZLr8sVUYemo2OIcARFcfQd8AiyYNcMecBr88lQf
P66A8+iRibiRnJprZasKeebiKXW7wS4Y8Tz3G0jUImxgxfp3T0tMle/sDJKArFnN
P9RotMnHFTFU9mpVywKkHNHpBA7DPenLaZPELP0PM1q6JPA7ydsRXgzJuZCGSjyD
N1bvtFCZTG7xQ/iiphvBT6ezRv8G7Mrgo3xehjKkF66pbBIibyx6Uj/wp2jmWT5N
Dlbsx5VpfEngpxhbeGdxuo6VKlQQBQ41XcHMeMW/DLB8pwarrLzDlrtKZkFougQ6
SbRKJJOS2Vf+vd9CnVlzbjgkwINJP6vviERodv0ddUtVZXCOYYRMgYXCEygPDTkU
Qb9KAnwgqEK9XgAHWtm6+ivmNSNUfsLCoZbnTxn9x9jxwODgG4KMrWZh8W5ivivC
JPsINPpQb1omOT6sqYD3y+RrdM2L9hYI6hdr2KWx8CzjXOJhex5fAiyRLxlF+kms
cEbY7Jzv6zB0UUiyi1rYflwh6G3XKnQRyU2Vcg89wclXbufuY4cnrztmoxnIb6W1
D5BjvcfC38c/DjvkGUZVn9Ax3xdhBYleV4PgW/OZjP5xF/94ZQsvvU9faOizY38b
U81Y91sLy6bBuugfYWtaMAKA2PN80IX3JFdnKzazDPhpOxzo1ADnAb+SGKrSG+uL
CGsRRMiPTNFlmT9ciT51mhidfcv/+Yzm//6b9w70aEafMCAB8D3ZU/BU23LfAwz3
f1VChwEjEKeBi/Lt1X6Qaye+ZeZQcj0o4TSZskoZXhhu4Gio1+CCuavJrd7zgEbk
ZafumuEeozNi/0NJFBcLRFCEM4JoDnTFpy/lAwbXrV4utEjnI+BxRis239MtzrkA
UPJloIzTQFLmLrxZ0/+BzBPcGFKp3Wg8bQFnbzfndT2tK9IIHx/XRWUYKj9HW80v
eHQoyZXDA7U51WwxufTkTIfx5fTOBCr9cfaEkOSa3kxvgnhunNXbZT2Jfeta9d3i
16bCBOM6y8oWsvQwnXhnwcZulnqQ58wZBu6Hevjb86KGV2YAXGytO3QymWRwSSdD
05Dp6GVoprtNVB+QWS11yZUDWAz8nOlxL7yFDgEBiWp5kcbkr+GIkjbMphoXGv/X
0G5UDK71LuD0MZMGdn+mC2ylBNGaUdGOLYtHMKKBTxzN6rCvwBimNw4Wlx5PfRaQ
wYGBEghDSL4dqiySTXAZY4rxB3s6Hayg3ejed3KHFNpM9oq02MDkIoTQW2h2sxq+
lm1hRRwuqDbaxxS8JtYIj4cwKBGdpql5MBFt2WfRmOCnAqHcH9edc2IEjMc66Tj7
ORU4zkIKtQdRmnZdRAzdK1m8lnOPrxNvSCEywkHDxigOD4IHfuXuPPcZNnW9PPFH
iLbJQOqmyh6J9L9xfSBsKfH2iVvla6eNOEr37PMeD196vIM7KNthADw8s88i6klD
HTiu3Fha9GWggLkrjAHcEwDdG/lrN3hgKIgmTIM81feaB0QqBmXS0OshMVWNU8Aq
lqqIxSleoozevGko9w4X3KrUgGE4PHL4/lLJE21QIGnKtF2b+2pxHfIIDDHuXx+z
o43ADuwixx9YQPxsllkRgLTjZDIRnQjz37WCjCl8wemdHM6GDLzhHHrlql8K1XlZ
hhe5t3iXzuwlg2+itBGACgbKAMHFomZS6Ze1PjLlyIva7ur18kWnRZopV+fGr1g8
A7HzDrQWepApOQ8ONnaxoIC/ptz933iNgWjrUwXN5R6IUN7nutUXFF/YPP30XJVt
v2lVHCLNzKBiwmv2bnI/RpLXRahz3QgyY6ndVkgtLN5kLfHuK4prcFkHPuPJ7SfD
F5RiOpr0p3tik/zRZePDIHwKWWvEzbHMSlGalU1YDT+PZaX9d1CNMB2F/dC6AD77
iyz57DMqbSWMWzPqBmC5AighHoo6tqZNxpqfK58z2U4AIn7ZfwmYTF5EjC4y6ZLN
zAvQN1qwEoW8/t4YHev8abaH7FnFeVRKhDNjWRoxLrz3XbPFiSOdCEpq5imnW2NL
Pb8+HggHbSC7sl/MvQh8dgttmw71henxSHjlZ0/4MsfJstHrjaxDndLkYO5yLQxW
DFy9sSZPGStJRtOmXw39sQX2wym9k0e+JpY00EMBDVtrJZ304Iup+stkaWStdk3Y
bsHbPC9UDuh2sRc9CJfQF9mRzMJjmJ5+dJg4MCmrYTn/2erzlhC+uYYRUk7Q2yOh
KqU+1jlZl/XDrFndw5Tg2qnJB3iKebHHmlgPcLnk1aOCVdjMa+rlzuSCLyhjpVQn
5QkWI1TWJJDuxpO4PZieI1knBnSB8RJb3Ug/XEelp9bYPge8RgmFNn0wi07laplh
LnYoixTvNIOhRDrSlUuk7N5Di4D2cqxE52m1n3FYU7EsDVSK7ptp1rgnMxF+DZe/
jyGHD6K0M0FONvsgaf18qwB4KqOcneAX/spy0PHKFsoGXG6XRGerOTEQf4uJXcHV
02ujSD2K0zhfYO4bjvgLkvHg0lsYDoktTraGOC6eLgRa24ATCietKjqIzv1vu/HF
3XkFi9q3Yych8ZQJ09med85C+LcaOXxvcYiJTVtvAR5VsZBMj7AGkTCNJ8jTuzi2
v+p/vwO91ms5CUF6S5MK3mzwTDeRaTJ4p6G1y4C46izCfFB9TU8HlorRmwubVAJm
3Qd5S2BRG3PgsTbJ9alHf54R3/8bv2DpXJsb6SDNtT1pHfBLTuzKFRS+IOgwVnxO
enhMn9Mq8tj01uxuDrmO6AsyK1bXm/qxJShaKGlwY/GsvnkuB0LfT420AWX/aPP0
pnFx5mKK6FoE4bfzWcBfJreNtaXtYn26fiWoncbu+mJRPcpSslFxvgphgHRxkeCf
9BrU7mIGQOWdaWhBa71UyL1HY6PY6uugEVM8sj53kIssT4KY8QAO/6sR7GxunBu2
tkh+b6ekp9r/AkWwgkimhNG5rl16CfaOxvO+HMlzTf5BPV1HNnKpK9puWEp5NYEf
osXswSaBvK1gSMOje2QwPvfnMh3Kzd7/8HASkC+knjwiAjDA6eK9dpABOIR+L8tL
QaoQYFTtx8ZWX/EX/lh46xsqOs73UzhPs7+1QV0OZ+LNohEW5oJqCs/HdQ7H8VMy
qh4g8hic0OjuEthybg4x5ps28J45A94+IHbk/EvzUmiSQA+WhEOIt9hG7XIYJmju
DEt8uRmAAzdTWFhA9UfR+5/heZ8TzWDALrQpYB8fITAkT0UEcOxyJiveMe1rfnQz
hmcFOGp8AuXviHIvdnQymQVAhxEAIiiphPw9KGmndf1dtg2X+8d4eOF/aDwKwVZv
5Q0U2ifuuS/WqE044vvv902elOoRuRScp2DiOct9dFRb6qQulXdwIJWNLYQlt/Fm
kguh8Fjx094mktg6C7QJ5rOSlgS9O8ixhMGKzkxvPL+Y9nPbA0Wu4hHM7kaxxqvw
GDmsYcrWHXM2BJwekE2FUtA+iCKqIgOBMbhWPAbVtz5GI4v1x0wYBU2RgS4G5+TJ
Gc5frsCJe99GdQvpuPpP+zs28CwXCOt+dBD9zhQcw7edXkcJ/E+mWICeFiYL4g32
YOZcRWCGJXDsqttmUKA83w9AdEws4dEqce1hRPrYM6PMNIEIqNIkww0X+qa407an
9NeI6KiyqIwyqBtXO4I0mAMfq9nRDVc0Ece5OKrrHj2EYS5MuMS2d479bYmNBbwF
kGleYMlGvDrRznAfxf4xSXmx1h3V16nRUfYhcKuhkCjzDG/M3rV6mAL93A3hQFM7
NNaedhrJcMbPHNcAiVUgcGsczDTMK2l4fvV4utea28Hl8AotFrDhMwc5gFOCOkkh
rSj/n1us5jaI+IjcucQISEa4dkRgscLv93XuF4z2W46eK0HBS/Sdy8+pbNw4sY3w
bXN4vIMZ9XuSg1sEyO/okYxu3NTAGgoVjfDt7vR6L9ZmNuWFpP3fzmZ+53skEtS1
o/CJb5VIBCyQQnZN8ZJw2llUIIWSXiMzSFhFmUBYlykQLw7wQGGyoQSmG3dQJEJY
Fh8oH4WhAcmfkhcamf8wn+U2oiFaY00ZVtVhrL8I3lGRSh8Sqb8oxORHdor0sdCv
6n/42fgxZo060ph8bjjPWwoteZiCuuXd8JnPUDTLSoLrbu0iC2AkEp9yNrVO/6yV
uf38HAC66qO+5sf3+pZtn13q1S4H0qz/p0LjPNV7iLgvgB3wvGQxBZqhnnObh/Sl
CHxo3jluyvraTNjlBLDbTi9BeLCgOQgxn1rsI8yWxMcEEP3TwXrX861Ee2SKjF+R
eAKISMhxTEhktrtm485uADgWaGoyBjV3T5udp1qILPyaGK3ZN0OIcmqUekgQln5I
Eu/pujLL1wUf6hb2sOQUKwfPlnjhDiU9IF16L8SQwrOW3/gLyPekYY8Dq/UtOm+5
iBhjeob+atIxusx7GmLsgpBnoqQnn8jYP1kTotXYP1ptXRVMU1TerKlfSI61EBsu
xytrJ2BfyirJ7aykmuUx3dvOi1tJPAPjiGhSOh+pwBupK/49fHGYhM7G0FLW6W4s
fKwo6kjzJRmYyb9va1M4jwU54WjI6b6cmOItrIHIRb4Hts13lTX87GhyvuiIqG5s
MjIR+1ozcdKT23vGFQjCbEe8BWheXoSbNoUT9KZbS1Ax05acNQ6SGzK8slmsPuDQ
y1x5O4eKBKHpDcLHl5ZtVWO5e8Mpz90FejAuaQCmcC8z30Bcuxr5WCVrSRjR/dY4
+cFekZ/1976yszw++zO4Iu3a7UGt8GDthkd3SCxFtJYEj3LbKWKQsAeOrQtVG7cZ
dTWWidlUe+VuCGYdn0enywDQQRAr9xIfakG3urnS2KSiO4IZLsIgJAtsUoC4MM28
mV5GFuGXhucxdMUWw9ISDPqy4B/LSL7egXjLZ9N+bu70gLS4vohTlIr8cq0wDu97
goJwZPtPTUJLKg2gS7cjwuY3PfJB4FwpT1DaPr/iSsL5/B4xUMkdGK5ydF4403+D
N2xVEWyh5LBKmPd0J8gQHiEBR0VhvBHAPsG9ADtWjtIWHRnix8gJKCsjJKEHJVCe
tGEqOlQyiDqAaiIwIda7c52mx7wZYOGZcN/nw3nwysNhiD1Vgt79ioKitRYsF6ZX
tHMZx77fMRVfKYTHa2u5lNTrgyfvXDO5QOGbUnAOSROdyZ+Q4HGwSTPSB5AkfeHk
zLy3qDtt0ZHRrbCdkUVmTtDwLUi6pu14RxLORSOXjKNWRhjOoFI6xQyZGVU6gG3B
Ywj9nIQUZvvmfS9xiVWFTGLP4ZtE89AlETrGP8ze+qmOYY6p2yP8DEm1+PabQWsN
d913aoix5f6xGiEww3eY4Gn2sL1e00DXHjguiZXDccbqpagKioXptTJGJpaELEFc
/Fybb27XeRkMUUBvByfNhQn05U1BJOo3DbzEI1iVcxwLPaibjrYcowWaxq40O4BU
Bw8YVXUOwEb1gdUPh0Z1eKOzb7xWKRn8UbdSRcD+I8MwRMPvGRPgNg8QTqQQdlJz
YBNrgZ9RkrMUtV9gJ8vF5hIanQWQySSqUvIrQVGZWN6xPa0YDBaRNf8lbdNM+VvB
0kiA4yTaiNk4nn1mtDYjQtQUWp3Eo2Unzsv8za1kTVCQr46hpmDOx8qGleWpaM7q
q2QHyK4oIXMZdfanWHZxDLXK3lvfBCTBF1JHxKEgtdJUNrNNJgK/uKM5wDDKWjnV
h1zqd5xQkGb3qQUFL86L0K6QEyEF2juGM7s1sEucweUe8sjJPEmkWKywTm05tRML
mcqn7k/0Fp8QkeIp5v8Ql2uE4E7gpd3/v0PPyEP5LB1MiTRhhdw/IyYdfFjIdhoR
fc7Be9l11vQkLOLhZ0tgpuv5d7AMiCKUO4b7LnqpiS5FU6Uv5W+hZ6Sv2/RNSsdr
+jAO92HsVMDLcld7gj/UwB7IvrpEQdogZeDtZrqPouyhnIqYVBppS/gTLX1j9ZK1
UMrj/Po7jEOYGQzFWC7gkSeJ0vQJcTSwLdrI1TpQN+VNevwFcLUrMWeVHV+k6ann
GI0k8OI7h9u0YQYhIAxfTL0gCsQ8+jpYG1RQuO8lZ8lp5v4uMZJZHXCLzCvVEAwu
r7td5Dvc4YNE0sPKZimPTSeWvP9WCIaLNXmQr5gSMZ7ccfA08k/ZK8rmlRxGKnPB
iDdostZAKqDgbA/c0TUa8g+A1ht7jX9JUDHggRpnOZRmoQiin6zQrlExf1yGVq1W
taVT5RuQg6H0Mk6BdTZ9Gcx84uACV86ngKyWLLMgVDwZDSkMxcIJEnPtHt4PQyrD
yxIBnSkKanBK90NYugCJkcjkVQvvfxXibssP+ax/ja+9HWInWkMa9S4gX5DBqpr6
CovBYIW+PHvEHhtbuwklmozRzyHBvqVgpLhsVXUkJFcZtRhQFAXPIlaBqs4BCrDP
by0su8qs41NCzHwHyiSMCepb/BqUoM7tmepkHjL7NTHpyY/0uTmWtj4NyLDk4SA7
YUIDKtOL5Ox7HYZ+ooGAP6SFg5gDrUmipvKRMBfcWRGwTwHFaj1GU8Sd1LI+AVtS
0ia+Lb9fk3UgyBV+/CoHES0elXkV/hMpwdxFJkvCF2ui4j9gHcBdZrTHh30ZHNcN
fOVBbtmt6aRXB+7hH9CjMIULtvoRNgfc+Xr7/zxal7mZ/dJwUbf+H1RxUaHcvXFR
6QhMg71Z08dksbd46TnK3Rix/HkgyATHP19mzuCNI7BEMhXwVd9NVyH18w7LflRu
crGkw2bzZGYjGf9Jms0VgmVPuQhe81RpET06NQYXFERoIYGe/NVqHhA21HCfbVEs
cAzDkzd+FynoNfZ2S3qveKFpnyjSLT2cXvxnAIiZDGdgKrkfs/q3AKbcZKZa67Db
izoKeO9869VjzvLLsRd9ufdkb4RXtkwfIxCHUn1bNiHdAT5pQqIW8hWt20PB7FQc
A+Mr/e09qywXKIWhUGxhJDibbdZOxOPcJ0oK2JfENhsUVuc4dyziIC22UB3KBkjp
AZUjnb8l40kZb1Rtz4PlB4/cMeufSo6ywfnvLAItF/nNNvzFw1ZRhHKCQK0gae6m
WT3YF/LtB/v/Ck6RMTJ1itEUE3V2iP2PWhH/L3hUzr4IuLUS1bql61i/6PR0n2xq
xH38RAzT0K7xKmd7yYiTnztB/3g9PvX1dgqe5kH5XVmwMoRHTV2tBr5k/sJWTh4y
80J82lp+bdc+vzhFNJFetQQV3f7ZbKVtMKJg0XGJ0L1JCPwMOsQfiSK1jltWAclL
Le856rb1vlEPziUBsvbXykzfdB460v/kh/rsyGBCCuoj3GAv0zGNQQHBBJEwDiI3
CxuEuk1hcKbdlJy3nVT7msdrt/R2X9NsbPySPc+uuR42QQWjbSr7lQh358Z6BJ1W
lzO2Ab+17arPN1M9gRHyHrCnjCTrohs/zDe6fms4Jt7/asffTZwXRLxR5VmzvA7z
/7utc0dbosqefcOiPwiu6o1b5HVBr+rcUXfISU72yMW3XMsNPyKbfmOblVPz2Cry
NtLqwrVQrATgjawWRqRKVQQ/1XqOXJFT4YyowOUqeHdqjr7wZX5Y/yieOXftwt9b
pQ6Y5yGK+PNxDZ+TYEDG6bEyHETCG7iSqNv+D/ZD2LsUviIFSnZe1BnvoT8s00LM
gCloz7x2UnuGRhuxl1N7IOUu/znplpSLZND7RSpAnp7tFng23JIc6lk5mms8ujLR
GfBj/PG+1iz19YoGgUfPv5tDX3WqtchzyYcQKWVXn3I0sQ1CxglZL6aDBTSKYeGJ
AXf6bkq1UIinE7hhU4bSDa6B/HPOQN/fMZhU4lWYyDY03Y9dv4+zac9JWZ7M7aa0
heN2C9I/vXi3F4G0TAtWJmWR78heeEsFdLfoau99JDs1mG3RIyIcUEBPJnmo20IT
BAl/wINuWNwIOZOa0m2oPf3zBHCwDY3ElWlAVKvYGovw0uq2cv1NEuGYpoHYz4kS
S1bU0G3Zd7mpWeYyh6t0WLr8F6x/pP+IVJlrCvRlBQY2xTnrTkrH6YFYBAIPsx9/
dsvngxR5fDhdFesHDfqWk3Lr2YOsdl1uW4m/ZSk9WGKwyfeir3wOEQkPmlFKZeJW
hTr8xsa0RnYKHe6lbpRUf30B2txiVnFkxfVyPS1G6fRoJ0DhrGyReSzVFkCb1Cwu
d2y2FHDSDY9csZc89SmhVq+SETBUVg8we9m7h31LBO6gYMJWQfT8oztq2WEY53Nc
14OYMd2h6AniB4sV0HHR+vhxwrr16TQLO3jF/Hzm3fYPMc/8MoSD6wU+9Vjk5/6i
NqFjje/IrNeuzPvFUQyXIhnUtu1wao3IdiK+eSewQbXImRgipxwDdnr8u7nvCJ0e
HfqBo+8KivU2AuVuQfIpj2AO3h/ewY4+ch94jV+tYGqhFV0PiHNIb0QRZPu26IHq
I2R98jFFruYhJkl8vnM4AQ8B9vouZG8ieyxn3h8JMiRLp/FiCvQhm2RdwG6Pkt7A
UHyMWeYFXxtsDlDjW+ylGvbsXtdPApczKVYViRUQfMB4V6xjrh344RFjRluzLY5K
6Lef3olpHmkFimo47gTgb+1VPtKUIolJm6Pb9AMO1g0hrDxquTs4I6V+2uPRcXUS
4aGfWPpawfwlQ/YcZrj9NLln23ERXXgySbckaVEBRXHPhyy8Z30YDRAOi9h6ViJM
Snc7g7n4bUX4G+ctwhQrHigLztaBXWb1JgwhO8N0ZYx5IJDzhtBOdeEC7mIOOD2C
NwSIZi+tFyZ8f/D4xIpIhNsDS5euE5U5rbDX/rlcFcgapPE3ZD2rlF3zkHy0KlAy
I+ndWRsyE1qKjLtWxCp6rMqnQi4S0aKEZwm4FsxrDsE1Yv4aMOiutsTxzGD/ip1V
MLhL7MlW/jV/Uwth2yxJ1e5dYalmLOKbSbQVEbrjZ4g+bTkzmCguUO1fGwkciwno
d/+RF79eXUSlRGX4QFXQXqpt0LMegMAXmO7Q7WrGuEqYdDgblA+eZAPVx1clVGQv
devqcZAB6qwSroZJzp/DtMe0Po1OCOHHvxBeHXHjSikH7btiTB6Z1BJRLHDOWIrr
FtfzJbf6WeOdgsZwIE1CL70jwKebqQfs9gfscD31glA9idbcP+g/iEkqbzm/6uu5
wKbGVkL2IqqitcG5ZmBywSeiFpNPwC4prxPRJzLaIM7CzoYXySLphnf8pLIUnr0+
T6SIFgc3NU+JSas27MtU/M/s89JeJjSErxEB7nagW5Ii6n2bjky0+QoeDnL7RTov
UJ54AMpJf/vHzv2ogOH/R3yvOaNRjkGL5JH163TN8MybFu+eB7lcC1jbhDlzXSDb
gsFZnAPG7KDlP8SrYHqntN9iQxahMeuQ5shjAln0Tn5BWVkJ4ftRbCxecSsZnhfl
7gM0avndjA09Mnk5RB1NJyTw6AhSDjRa/kNcYLHunJ4ssqT6k9Vgij6kiRy/iiVX
/VP9tc0x4WQhXMbuxVVTibkQVbKIXrLW1MDtcnei+pP9Z89SHwsNDy24gamU9tXu
E4zn4ecWwqU2FqutACXGd85qlAnwEa9EzuzCTNpFtlI6acMjPbwPcXVByNvixyEH
3145RuznfC/T3jnJNLb3wodzzuDpsE9kzDypNxLEuPtcHMpb+rY8jAdeSOiPA7gU
HsMMgYgIN5dF8FuacQXXjOWQ8iy6zr2ibiUaCd7N1Y8T1Gzdy7dsLTfvEhV7LDdA
hPpGysuaFp/H3w3j09Ee0O/9JIQdV7T7+9uOEVJonwkUMS+qHVcKxozeD6Eoue0Q
NVH9ZFJ085CKG0vj0PuQmZYLz32r39XHqClEayiZy/+t3d+NovtYKBkNgW62DPCc
JPPECUfK7CYbw2EoBklDiCUCyLZ+PBJw/fa9nq99Avx49rnmTnEEE3GjqKZHrWaQ
pFXG4wJgG5e9kAFqk19OQX1XpXGBf5yPCgL2/tRq1QvEtYcAtGKSrmgr0GG3dOV2
6fgu0D6H6/8TEGHeI8yn1y0O5mntXs8RV6G8E5ZhfW5Kq2NgC2AocIBKL9APXQz8
yYb+DuDN3ac0kkm6LHffVUBc0wtjDO4jOOVrw10YynYV1AE9NeZzAak9JSPRglau
kzvsPgH2uqHKfJNMHbXXX69Y3o9FQD6UxVN9Psc4xmwB2bqOhC6T+jiWPL5iekrp
CQb/BdRq73mg3yiHgXljBeVyx3mhJetpRNyAZ2sd0uzpp/vmwrrzMeib58vb5TT7
CobiY+Ehhng+gbV9zUpg1nhX9MywegVfBHJ+d6Cz8+gYbfqfENoKE5bxUfLqbZpH
MFh9TmC9XZ3wZsMFbS5dlHL+GZpcXa48i9AqBwXX1khS21dOeMP/G5/3nEEXez4Z
mRAfXIjqbiAYKM1X9NVwgEHnRVHeq58ULmKNI9GnDAG/Kpicc2v41pe80vUHHXa0
0diA5ynmO/1joedTbgyrzzUYqaJClt8jXOeZQkl+TuXXnzpZeujaIOunDj6SI5Jm
m2KTLOACmTpPuDUpQg9vdwUVbiDLvVe5B3OmEWRRTU9z9qMOY2w6FYaFnQRysyjI
SRW9K6ms1sSRif0/1Z09E6kDKXowC7nTxBKE/WFG1Yhrr7ND/qEYXWVoaODUjyEa
aabzq5cvQGYv//uUocBbHiTam/9NJaKQNVjjB+9bsZoqvBiysnmeBOEIs7ijSEX5
yrhnSjtGkE4FYlwjP/VAqyVKtby7KRubIC7X2yoLPX6rtV7M7WGNtOCiIxiyLslg
wvbAn9AQXTAHEvUj6+HuEWXWFsKstx9axLzfW0pyAN96qCM7VMu5FXwupFYRAcJU
s+/WQqURq5NN1h/JL9Sl9aErdCudFu9Ab66AjdESWVXVk9n5zJtOju2zzCeFsOfi
fSEfkzZA5YY9EdnES5Ecq0mRpVTf8QwqbcpVPlfi8AYdyH6qeHsF8f2zxFFf+Vbs
wnKIu/tUhY7e0vZxIfjKdSErYkpkOejmPWeW0OLHcS5Ne083ig2htwee15x/d/Nm
mrMKEFeDyaDUk1QyiE3ktV2FYdwbaAlMmNQqRlPdxFIyOXOXb2h+sQhXOarEg9dp
/WgzhUZh7kAbesWc0rcZI5ufJWo0yx8HOblr/Pznf9zFfRhCUVwLJsEZgbLJ3wdq
h9OGo2Xbed93juodJWeEG32Rh0xjQQvPZtDEMDIDJK7NUm+wGbrsaMLg6zY4P9tp
ou6gcoRRPaIb6zQbfTCmP6X91Pv2CscnR7ndaLwOgtSVKyt55LWorGxHsIXny4/L
FUDZrhROXe0k+3jOMDCZZ/7SVKl14Hk/L+EcamRZRgrP+Af6QsEbinmqLa5f0hzV
uG2oZrXbb2pE5ucRbiMgbizVSi+dxYmuqX/XBCuq/CCzvamYQtol2JjXxAf7gYfC
Z2mtzr3Qzhv1g89IhSrgeiHPYhHqnLuYzqhtNtkVij88K2rwMencsyKjjGA90Ul6
jyJkfyEvSky29T6Fhj2MxflnMgaS0YVBRx5sLfMh2bEkBv9vWpCdK1Pp37qLHFHR
rEXlWbfnTRvaRmt4WmJFzfGntEIqjnPT0gkyqi5LCAth7nwkVcKGD4BCrx1JHvV3
lJRLuJcj+m4UhN07QqB7vScKI0NJirOxkQdqk71ajbFbg3p+kLajuYZJCZ89MEBl
lbPtx8ETV92t3h436BM6DUf7N8oGaagvWmsvl6uoFLI6Hgdd8ltskN75JCa5nXeh
DZ0SwN4ueOKqi/ShDsllqqiDdyPaIx6ArDBe1uwBKd1RWuKGCiffeKbUJ2fN5/eI
odjpzA+rAF/IiNrsLzh94m8jFhd5kix+5Q4dzKaHAT7xUAunYIP4ACIvEJi0W882
1jbV1mWKP5AVq8seZmaaEXKm2t/KQFEbKpklGMSKITNssXAbgXgxh85yFcrEbjh3
rlXVtOAhfpInXCmXjCKqcJAmx1JYVKF3Rq7TkdzSrdmVUGfR62SwzMe4MMHMFlfs
5diSiOwBJiI7iVol/7tWJSebZoi5mPCk9ZlBanAAbbgdTWjzfY5eZhzJDDcQO1/9
UiTbqLgbkUSyWgpwRAyqwRN3n+zuZYSn6CwLahuuSJh9Qru0Zdm7hU3OLjDCdgGv
ZhKGUS9P4HFz0xNG23AwBgWIh4zSDSK/PGsxNTparrseHUTN5xjfOJc4ZLvJUWHV
ggOVD4g0WnDFAqEo774w3bOWz5OC86N9heFN/H/zyJtq/B0pLKWTpEIt6tqg95R2
Mi7Y8M2kdzkax9daPJaSuZprBak8RmbAvMa7pi1fBPzm/p8RdbH/xG5rAft+0X2J
OvdGPsl14dW46DbRBAmz9fBaPpEYqSoyEbPI+QjbqbYUdj7/Pqal6NUlgLiE7Iwa
ma1XF6RHr4qvC195Agzk5FHzIaNaB8+6HRFplysNduyqXRPe/Z3fXnHamzjvGD6m
5NYM0Y9hHpCf8K/KevwvNo9p7IfQ8Qb21+jSq70FVkS74I8OsMor5JsE7aKwUm+G
i6L9Kq56t5r2RPKmHWgmtPejA/4E+FRbXi5ifR+I1SRR9VD2gd8Vi4xZDh/RCvjq
A9HR98Zva07AYXxeyV3v5ky8L/Q29qa6a4bJMmVmpbyrTtWlsvAvkj5qQRq9T9i9
HFiGK0MOtMxkAOcBH1dqZyhOcZJsg76ntsOxFvwZ8MV/fVl8wNIXUi9bxhGSo7Fu
0sxbkmrv0WZLwIH9wDwH0hQl4OUqDP/RfNRNH+xQ0Z970srySOtUUo+e4fhqJjXM
n3UWmhnybWmosBIxxBKmvGDAF94b7N1Ofw8KBJzdjpkKeKS9gIuV85xDDc+z8c0L
1d5mTWa/CFMCdMy7ASSmjuew8MhjSCfk6JTUtql+Lxh0DxrGGqJOymspSQ/+0kjf
AIsS2VVreMQRzPZ8Ej/0QlZuR6vRgFjwBOfijc+Cab/V5b7u6Lus7NhmVV4s3dwJ
ComQZmNq6rcPLayg76/lK9PKC1vpZgO1MWTlbJCZw2hpllt44a+FuAEY8hhCxtgW
b6MT2/myeOQ08gW2X0PRKp863MsQy86jHSJwLLDneob0cy6q+DprxB9djpt2nfuc
Olhdekpkm/oVMpCdtHJ4KsGt8y+j57VhyPz5w37qMvuw5WDPXLVKAzxWyU66SV4+
2eXQ61o1I/PqdNoRO0f6RdBfOeEOmfk3eLIWYmBndIeLixpQPgCIy6c25/6ipUWS
fWYaQP4jf029x0/LaQs1DDhGkXrEOrlNzLBThbQYAFcz1fo8tEsBuWPUPcwCauXO
NxY3HPrHQbM2YN3V1cnisNN6uPFWAOMdMOeNqK6rFb5HE4zGmAqR4opvDI5nmuiT
g0wNIhjUQJzJTgh37l9vTDmzp/ZFpW1QVz3BBbw1/Jk7TXyicXfF9732GwB4R+68
bRbPvKXO+Fd5TCN30/+chHReuSOrCX6gbASLb2zUZl7RI8vGj9meBQUV7Eq8v1/D
gsvs0o597JEeGwKzktHR2mBiy0Ipr7Ld4PLpmyn2ZScOXkFWrNmcBVgKIfPObGMx
tfZF3s5GBE66/dtcdIY/qw4cyUunB0EsJxixSzsZPBoKbiFFxcJXiLVVTf+IJFHY
tFQAZb6yL/2hnGJbWGD2lxn06BO0WeHQsTr9ZSrJ0Ot5UFtX8XjyI+2lkMmqUi4x
fYuYrWkxn9rxflHWHWZWrZqPh1B2Ta2lKmpmm7Uz4r6X8aCkq0lvdfZBlN0yL8q/
A8VI2gheaaZaGrp7hyi7dt9cKG/rtk6w1VDwgoWObyLD6jGZ/0dwQAd0wQR2Q2SM
4y7XtunrzicAWk2ne02Ti317esqyLlvOdk+vpuZFOhwn9vXtEQSnSicljYhIFz1C
3piAC8PPi9jWofPx1n8ofrJh2V/glNf/TJenQpM3FcL2PbD6bEwNezbVDFTnXZS2
TBtlHVbV0k40xXcYl62hxch0rIWGcIFTh2hcDv9NekjggN6F7s+kGi94bajoOA7a
5J9KAFEheR9YLnWAW9KConVo6zOkFxAei7to7TEUA1PdYMRJ8bK5Xt0C44AuH5Rc
2Ysq579kmZXFaQCV/SJ8AJBT5YHN6/uclJoIHJ3e1wlU7TaaKKks4G+3XZ4yj8sc
Gz8q9DypXmkGD6cIdQxHbTnW0H+/+cvrAOZKzJC/tHQYgq8A8m2QGwib65tpDDm6
XcHl7AgJYzqqzKIWQFILiCQI4Muje/B8MCLtoqu7mASrxTN2B6H8qB8N8KMpWkhh
8ULqsUzQb26Ne5IFndNu1KszBwelw3CKAuv1RFlJWGa1v27fEjOlu88GiW9U5S3i
ydRnKQvAb/w57oHzuiFoqggqF2EmJzDk7udpUyUsd3/rXxZpd7K5cbhu2XU/e0+N
iff9YiYAUn96IaV00dss6j5iL5hDB1kr/1YXEiUsJE7DLTFF+ANaJxFUlAGMurbJ
U/3IYfVcQ0nATHhuCLGqfnJe8B5pBcA453JHu8DDz5yReECm4MNzJ6NOFSmKyGRl
jp/5LZe25riLcRfqqAxwqzhyyocIYCr4xcufIkqvoYc3LA/GP4slZuw6RR+WHden
djNxUB4QQafKVg8T5KSnlBDxE3X3J69Wtx83cU0H3/tBiaGMRE4wOdzPq0/JGZCG
3esSdU6j1i4yeTBzsRktKlOL0GjF0AY2HYpB7FUN0lQRjDd6kuyt4VSGmeSX0x6L
Ga1bfE5LBUXcB0gAqpRDRBRH5enyECyp0Tlr9FJqRENXvnpj/JTh0P8CNOdXoajA
OeUR+/gRK1dau5mOte5txnkwZvbXBsOXzmGJGS2Eoe9nX3OKHblAGYQ+ulgcr3QF
Mq02RLenRDgU1XMumQrMjDOXi0zDCjdvB3h4psJdNTltEb47qxOWkuqLioh311ED
+/gz4hyWGTae8COijFMbw4o2lIogWC5Js2jqtOCVHNRs/55T5ZYttPoqBi3hUvre
/n5cQ6M8QRxbMHMrNNg70wY2UE3/DDPlbZiLSiJd8etOrWAWQQpzM1KfX7t5ZBmG
SLfdifM58TQcnxeFUVuHvsWrr+6kbONX10d/lPIJlljDEHJUUdSW3MxBJoTsUs9j
xvPJS00X53dUjadsc63gZzXGE4JhEveHJGCK7RT0jpubtqphdLkYvR+szy87+hLS
NRB4KQq20OCVR4fCqHSjvNQCf6qPpH2j1Bh/xQz433x2Xt7Bi9tX5JPwyHH64Zr2
hTM3BiaEVCdmfzPmCneUXEYavj5SgEFaqQSMY+SvXx3HXbYsA98xCt6pqW5dkYGR
w8U9psTr1TA9D28f36ZGdBcuzpHH39oxIVw+GTlu5N1TM6/meiYLG89NdyomC5H0
18P7C/S3tajS2zZX0s33kvXBV6lYf9y4cm8qjWl4sMnvtwf1QPNOecsKCPXwO0QA
+PpnMDu6H7L9buiNNCfqnpiXLJAPXZak5hCaC3+3OmBEGlRk3aeD2+MqoVQLNjsC
bWGPhGBtSP62OvR+BLx+OEEqOCnB2VvcXcVC3wTdImZHkeHFQb0ZZZD4jaWcDC/b
yM+cc9WCPOD+z+LJyRCvsnznR2VDqsw7nWwSGiY2GFdj2s6BliAivArjCyHNYlHm
uDXItal5xFM2q8I2ZcyKfnF87qZn1FwrxG7qx/41pzCVkdY7TjzmUv4n81OgZOE+
D7FAyaPddqzfOCV85qhuAW+MJb/ZGqcp610tqm/QiXEP0+Q8Csi248cI1E3smgL+
ZrEsSiQnjSEf7q4aQPHSACiuhNXcqfRdYW+GNdFw9ZwrJyVWg7M2LUv5zP2ALuiu
zjMufwniNyzvxqZ08fF4envqHyzvhSWa/3blVcc4KwZJtuT3wy5KllJmUiDyuKlu
8Bl5juujWyQa2s7UVaQQCL+skPEbJG0qcw/mbZzNp0ScYiYg6GK8OWcJWeBltSmj
jyzH8fFtHVeou8EFKM7+Cn80k67JilofSPV0JggTIujq1sDfXvsKmwKz20roaRNY
em8f99oTNUSuCdCiKG2nSsCgkC4B5vtwFKrIVIGzjYFwW3rp6JbqahgZmedl/0sa
uVHvJdCxW1l/0x+MXK1Wjcd2RnrOGABYnJLFybKZR6SwYzmqlgC0fTPLr+GaIGMO
QQnpRAKJ2nRBeqJJ7GEzAu6e431dxsw0NHWu2FuJPRP9Tp7m+TMcoK5xmYg1vKS2
W+cp8ml45BeHnHnVQIrEwsxsjXBEvx0yeOUPlcyIQw929AHWe4+uOMmwFk9P+WUL
qnSoLG8UskHNydLlRHSJydXYgDzQXs9TiFWw5wiz9GjueWZ+NWVCXRXchBaJW8Qh
69VzkBBSK891ExSvP+XPoz9Bxc0eVbQ3WYCowZQvUsr8s5A1LE9xPlVdfZVqUdu+
SzjQZC8tX4egW2p1FLTdAuEhbZBa7+773MomrghgK+DEOQf7UUcidTYBOU68shog
shZnXfyRXdIcdh2sZbSQBJggf3+v1lwDgmBqGOkfrIueW33o0JmiLx/hLImrZUIb
mylbCQ2Z/7Zqn/uirSzWEeSQCFeS6P67g4lXQ4FbJJqChUsfMky4+NTIsEQYDKAa
ohynxPFsP9wTyIBN3G0laNhqVyx08yS1Fscdhda3A/4dTO2bG8yniprqH2CM2Hmi
bPlsjGbVJk44Fp0J0nb855F8tQxtutLGnQG7OXwa6Ls1gh8o3UCdYIRH+cQs7npz
k2bY1CEk7xAtHZFoLePZM+BF1Sv2n1GalQd3lygdnjhUF/H5zS+QOcHI8+3KKI6l
f+dlJ4iVZ/6JAu49eqD5GpiPGoUXSvrl8VyS9aYS1FiMK9QJqTG+Dh6S9/sY/lhE
QjxoP9A6GNM6+JTThbNJ3ePXrQRBfZA//Ts2YtEoiV/iTgrOh4iACrLDgY0v7JXj
eNSjv79td/rY7BGRZdAhSVM8fgi6SFdI8jsb2YSIVusDus4RzMVOY3aUa/TXfp9v
h8dJTkfp+6HYDp/T0ZVNEiRYw7+ItbSVv701xUpPCQYCqQEwax3XsBpoN5C6V2cq
OeHhemKJ838B+L5jPFexH7gyyuQ3xGAvH0/+i7+7Heg5JiOVZvQ2hqqwo2HzqRnl
yBoMR2kWLQXfVUCQ4pG92ppwYOophoGtrBw33fkaWNDL392R9evwFzPr8ThcCDGZ
nGLsT8nQgkw7d+hYE9Z+O8d+xDjYgx7jhIydgp8PTKU5Yk2Pkr4yV6Vyp64bksLp
2ljJyJSe9d6x83SsavRG6FusIS4iEGAYAUQ5n07gzcI5VquyIW5VCMPaDsLmfGXK
x0/j09GXBzM/PdDXRnNiezFXyoh0f70gXUnFWaAAkaoJvLK02gmDsapJCnheIP/w
3DqC6nhTFVkORBxzktoPCZLX/59B2CWeXXSiIeNVuSfppISRy0SUpgpideH1cLwG
PDy9vNliLIfgR0GnKDYSWK7R6zqud0wS7vKmXcHBNbmsZEe40KyVlIjkZDhEAn4y
NN6d9eZ9bwvkSIhS8IfTUzCa+4uK1Pv4DvYNWXoQDb6fRWAgs4owXgB2yTtP9QKd
CUpbDHKgkihZS01YssCkVm9j9IFUDguvmoyemeyulUUId2S1mq+X7MVWSFVfxD9o
I0G/hBSYlprZ7JUWlB6BO8mfgG+XSAFrdj8t/aPEyl4j0/iay018nxbYDTX1QBQ8
CgobgqfbkvU1CLcf9OXwNFWb9dkhpBlKqv/lY7gPohuTq62W7NUyt+MNgMkANiW/
Zc2SI6F5NkjEp6We5eJH9FKeNLgR/KaPVKM9DtfWbDazXaO5oFFriab0CPyRTFhD
kdpYsxLBEv/RkPSMaqJ6AMtvoBIKUFONGk/+96vhs9vffAOtDotVeiNAYG7+d6a1
APjWe1Gu4dIBBIHSPl4L/bfzRaxlLjjMYWUoAe6mSp+rXyywmPu3Jy1m0RW6H9+N
h3dP+C8/zTcrh/tN2p1JQeCj5IdP4/xnNevcrdOlH88d/1W1RZZMxds5hHcdnutu
ouyduuMezie8jhKQdc1Y9PRan2tFrWOhbR633/l/U3SF6u7E2sM3Z/Fk8tM+uGxw
drbCRwiil+HBqX2Xn9F0QFaoDc0nBFNfeBzeB9gzsCYjRGThrtDXbQHhpEFoU8bD
JSrmKFOH6SC/yKfMp4AsM+70yIDhDb3dL3YtuZXvbz5v9pGvZFgwXzeE/QX45dpk
JIBOjnd9gucNw3EAvBs2Esb8iADlFKLcKB5YTxx3Vh89p3E3vAGxbHHkpa5PIzxS
9A3Mxlsedj90nmS309nk5wLSdWLjgpZhMW8okJRBATw9a5TuOHz/JTMQ2/YX6aUe
KiEJP1FMleual2sEzykmYR1ZOlV/mx8oLxGZ1RVcJHgMcYwNp7VtaJhNjVJe9CoD
0AOLlV5IV5G0uv8My84Jc5yNF8ehUYFiAwgB2moAW/hS1F45ReKuoks4040yhOjO
VscIqTj352W7/qCoB89HDzyt3L/Y7bepXM4W2PoNP37YuPUbJ4j+Kmkd7X8jGgTe
Qn4STcFupTXOQ2tewQBwLOhjho5czTDD2LPmYSDgRNbRmQydDJgNUjHYCWY9DcfI
7dNzbZwo2+6pTy1aRBVxGeQPMrR/6SCzNYCfnnaokKgh5VhjM23cFhXsA26kSUh4
oFH67ADHedkCfxsESHq7k2dj4hya7c78XnG+73JbMtoTTBWW3sxeR2zUli032o6V
Kvfz5tfWzVcJ1AEvuK0WlX6y3+dYn2a3b1qX+RbGGEt9rAxwRng8jXiYkcR4r+zn
HWPDddKUpKCdtIHHbPjoratZ8JJUG8H6Rzu90Bk6qtvIQpVay40q9bmU1jQwgQtj
7lXrW1s7cXNOuZctXCruGD9eru6Ma/Y3bfpUG8Dv7Pyqzv4oANP4lDB0QEldTjce
0KMuKpjnCnDgzq2dqr6wznfg/hORGPxMZLDJqDW3Bkwigt41rMuqlrUbOqcmqbFZ
pcWbveXTH9EDmtsoUXjVLRJbHIkZKG1PWiSCY2L3dytrG0U+BkU1z5RuPKtGXFvd
JrQojl73LOkCfh1eT2qRUJ+1ysErNdFpbeJ4NoAOGCLKyszXFgqGjP790RKyQGh3
mV+sHim4A63DkgRv0bBNvOjzcXIn10UdMwNLqizc9LnOvsCwC+St31qnEZ9RRNOd
pUzeKQpe+Zj9HR7REZj3ya+HbAyVFYwaT8I+KhBzLA5ZU+z0CSyDxNMscDUULV8c
/8J/KvrVkWf0O85ocuQY5R9H70jZu4VcTGJHEmFHmnZxBIY3Jg0xya089i9Gwpl+
vHaSi2XrVagHtJ0cL00dm0CBi15BbWs574nl2lRp2hcOLabBdCih1+W3qYRLki0f
9b5WWXTu+urNZZWPac7kp2w/LLibUc2c68iDJFGLwX2zxo1PYeEDO0s6N/z6hu9X
jqFl8uFcO3p54ZQeYu891WTniT6CQ17E5t994OdAV2aCphPw3QastQcva95Zbdoj
asQHLhaA14br0bCpDeAvezMlkHz6H1yGG88EVRpaSAURKDTs3LlveTFpnLf8J91Y
9OwJ0HlvY54UzfJDnOqeH/dHt9mL8KV7P4UfwWOUojuOlu1/Wp/CJzoRXO2cVssF
shW3lzm3iDv7anjRSNjGMj7eF4LH4tCbMY+ZHYK5Bg0csXNeQKTRJx0dBNlSzKwf
UlFOpSyT0LUFpjOjupW7XGhdJrBPBMzgYsRpymmdeJea7ijYJkBhYqbW5XeR7iMJ
trtUK0V2MNk3QK36fUfKfCZIKYIS1+/BNQx0aJb2CE7GPaYa1eeZwdwTjLZS66dj
VInIoRuLgYTWBgmsNtnD+JxgJEdboRqTQ8cR3YT9FTnJdth4LaG0O+YhkE5Gv33W
FmZfOB6j5ZHrrbdpuVNjAVCDDHmk6DO41X8BjzuMz+H0AICkaJIComEjsjea1URk
7Yz+nZ0imihU+cM1s7yhLVLSE99fUHixUQyx/1mK+fW85ZXok8wl22Y4bugQCWmV
36Wi2uN0deO64lruTb82d+TKxvnRS3sWiFumxDblpJKN3Y/m9Yx5lDA8nmn0CbDg
le9JCldrSffgYyRqp7WN/+TWYJggmsYd4ZdxzT70P+vhn4bMS1njsyytOToIeNtu
2hn1IeHeAy91/Ce9FZ2KBEQ2hwmocA5XoXWdPCLQ2a4LB8CsTLLljCEjGXHuJ6bB
aPU+x6QpddtTS5ugXjuQ+kzwkkZYjt0ZSEFERX2MqVEBMSgFSaPgbJ1IEWgOh0J5
ADWZqEyVRitVAr7ZXINQr5sfA6yNd96+oRv2F36e30xZANitSBYhYjhimaTxlC0Z
b2O9XKsh+lflStIv4QFqjT3R+AFvun1lPGcNzSL8OJKBE/ZRl4ZpFxak+ooUpt2J
bryaYU9Kf9WrJpuY8O8spGc0RoO0pafdZ71ZXNww3gtTmUzpI+vc5nbz/4J7haUW
e0fJ9yR/JOlNqgfoKA1OckzkShxXLUzEenKGrzCfby2leK+9bnfHHX+KxconxiWW
NdouhjK8Xdvy8168vCDf52/6dftCxCIqSNPLltAhuv+lYa2P6ZpwJQ3nXwWtenRe
6tf5/pecDjK0MJ3U/wBENjc3RWBHrWlbCPjLG3jBy2GyK1qOKvXMeB7V3yO+nA0k
VILjGedPuXmPqgkMXpUwjmzSdEUMQ2n17XB0gj6d2dOoSZ9DA1AMG2R3TIkbxdjD
EywMlkP+X2qVe0LZModr7XLhdjaxVzH1/tSZaawM6kBTRoLTsiZYGLiAYNmGk6cS
OkVz2wpIEanulVzjNAaNHYB08501/EwWU3cSxDjrw+VPXRfjFkB5C2UdpWLt3BbJ
cY/NaQDWrb9f0J9ekiapKepOKR+4bi5FLfAaSkBpV0CDc1z56N/ZdszvEDBv667S
j+XhUP0ZDh8C4BO3gmvNX4cTSFcacwOcSrXFPnlARONvbL0w2Cg7Dc8sWVvmxvIe
btkE5UHlS9FFdVatpdowvzv1ZUAYQPeDpAxK3MFyNn4uE79gYPluoBOGP9ksIw2i
X8yle15ItoPfA28dQJvdl38iTZHNnKtpyQ5I590oSEDFmSx5MLEAct4EjJe8wguL
OeEFaBJwZJgq/uHbruHN9rIebS8QQ0Ihn1KwQuKm/pMRdORxQZw1IqOdk1Bv7riJ
FcmV7CcQZ24RCpt93LzE69tH5ss+AaBNJ0iUIhPK+zNX3Aw3/Ab8cen9vGx5f3n2
9YMnomxvaJM2VVPdDZZ0vbwuTmIa2PLwaOvtW8z21M8+Ix/zA6YxAvmYKDilEEu2
mBL2DKU7cs9S0yVkg1Itiu/JbOKTf0yvZ7SrosNONtJqZ8MEzK4qaqE5MwsC/r45
MTVFmMmDDan69C8m4UK2Lgonp47WHm46j1Pk7NFOxJPxZp67hw221cnlu/+YLxAo
HdGFQnmZxMQGorrZjdIkBcytxk3PrnmHvwwmX6UAxotIyheegVcbgV1d4+lG/uMY
qqaOhqjIBz8KOMhdsA+gioMf/dA2jrLdnLEpjir9zGEyJRpKBToBIgaTGOxuDvUN
xA2x5B/fzQNUe/73nLQKFU9aEhctYV5OCgmi0TPdiXB3fqxGfu4+H4oe/Pi54O1+
YohAvTjeXho7iN2ewVPk9k1jl+W0AyrUYX3RPRHKFp4J9W45GJxMKWTsh80kg+9X
/P+dhTtQvHa3ByPPnLlBzMSXVHSR7IeUeI7fSU8di7T1dOcWLSL8iwmwcZ8yauIV
8pWb27nlD49n6DdVEtofuV40XnU7G/eGXtLwcCJFpFipxcGgmXA4EysZ46FNYP8J
K3V+oxvxQXs6PApalGF85WMPGvG1bmh7zd1UmiSssJe5DV9KtTrrwYOKrFrjUOg1
CTtpvMMXJ8Okc3t40+o0v2la//VmjWaA/NUQsOUUzUb0pO/Hz51o5wZMOhqx6Iwz
l7x11z1xX6ploPD1rKXuVWhkl5dEyNpkULN7tFRoXWqzUh4bAfl1k1bGz4YJchOm
mW093hzPMLegpGXWK4fuMRqVOyT09kdo5q9rRcj+vyVs84SzEvknYqYcYtKqrF3z
yIEnWwnZHyfFUMpcS+PmPeYVP/XkWKuUZnUOrADQSbWoJrmMQJxqwjQi+xbM4wUj
iKN4N9AkUoLLj1Cz6emh+pCWz99Tgie1m8Z3HMkyMfnAUsOpdTizdGHDZ/V2B0nC
rALSmwSrXJJD/eves050p/5k431fRrzvLtNeoN0alehkdtE98z6xGkEivj5/zFS1
Us2/ebxrWLv6jFjPrrYWJt3zzsQd2NwmeCDUCxlqCSvZQjhaEwT0r9zWs5aosYOj
WiRvkFfIkXmVaymBfTKSNObwnw1xX5bHDKUr+fzPzyl+jfVSb6oia2YmaQK6aOly
1PdkgseB7tz9aeN2+6ShWf8P3TPCvmeBZFLgwt7DNa7uzu1fvDGOvbm9WmUsoTvv
Jfwjw7u6d9Z2n1qUgfEIkGzAiI1Uiy9hhoJ7Be4PnSSsEV9Rp0Diiflkks2kF271
Erw3zk6joefec4nv5aUtLvSYbf52EpETq+99khbONipqw2A+L+OVPRygdk2GvhXF
i8sfXgomjDShe4u8UyJAGB3e5lMkg3X7hG58vIDYR2usZRZl4d9qoEhX9ccRTnIX
gBGTtjfcOeqWoX8eFgEtntWCTVQv0Tn9q4qoP12U52Da0g1udPUFcZhbmlh6P6/K
VpwFeFTfA1xbLU/oPQsUtEsEaYWz81d15Jz9yihML1xl8OjOC/GVC5dIMVwqCO0Y
rlZdZsEkig8bZjloTWhpoYptMB9PBYZuxSueBCEfjOS6PIlK4IxCZg2giVbwZ9eq
y3fjbISj0yqvxvztIAY/TjBozOaCs+UkI6BCaoo2LShBSLX5adTPzqc4xu/vXuCu
/wnZQKDWnherltnvX/G7NZdWcorQ1HfR6jjYvpsxBZHJA5KzlUK6n32IoNB7wZRE
fSinXPcuDwqdAtHa2rd+lyV2OsI/aDP/DG+wpbhWA+1d907vXTJcBxQIlx5Vlp9E
jIuVW2HOhfMdJm20QPCAdgMS0HaJ5unDAiCciFd9h2+npkmW2EZYHBPVT75NBkT6
2umPtDlKYCyt1a12kJ0biG9/uTFlbNFWqLMp6eVzs8j71nRXu0vYwnrbGykWHbbq
Plz19tDAKGYxmcBL36JoakCokHn9ShkJ6EyKtlh3chK6hFDz8749n42CuaG38jA0
Qpf2OMLwvGnLpEjroCgBIOf9GC53aYwunoLsiXsE0WuOw0SKv7xMnNEUocIlQeLc
Pou3mQAZoSqcL65fRonyLyT5u/4VuQvq9VNMY5NLy1rdQGOB+9jLsGEG+nsnP/6s
wmy8Qmm5jCFnYIq7DDQD7fgm/KxFCidAuSTprk2/GsO8BrQPL9QLn+wt12tiHWDT
cWNr3Qpbrk+guAG6pB8swEH6dhScd0UypY5vrHf6m1mbRBHu57xjkPa0lChapMnW
/VdFDthuYG0wgxa1MadY2lcmLf4HLDhJnMt2u/hx9QejbyYPNO+vq9MOmxI4QJmv
A/0m5bS+kW5nXb8CA33uIP0gQfEZsqEsv+RxPk4UShH1WXa8sZGWyJptr38pHag2
vacwSIFnZBZx3Ga0T5hEwv3l33g9fbYzCEPFfPWzrs9TmCMGMmKcki9sge8LU6IV
Lkovx+bNIohXIV+dxKPP/8CH4wXfFXufEniuGbGwoI+yYPC578QRmoiv0tyR2N+a
Zld6sqnlrLnKi0HUxEHkPTGXMJVR0b63s3P8Q2tSkOydLuzOOlL2mhrNm3DQxkU1
T/QGiwWRvvHqFJm0e7RVB3iAfqG2zvoooAzolYNJoPhuGTEtg11oCJI260IeprMj
eT40Mi0kkD1jvikPnfaEKtPjCuhOlX3OAQKz77xUvUsfWExGNzDdX8pnoQH9x8Qp
a40XyiefOwqso4bgQPrwehYb63KT3UPu3rTQm0BgphnfOl1xpVvMecQfpp3a+2Fy
BAty8HfhM9VfudZr7RxfYPyb0lS99ijlj3a+q2YCaYCxBfr+TJevK0sV1RxibKuk
VFfr0ttjb608Bal2s93XtC7+mgx31Z+AXcXOwIhycX7LV+9D2+Kkls/0QHlgy31T
5iZ2i4UMxQX/NQjkdKKRBCJf7mqKgEUKHB+S78nuc1yxaomz2Eg3TqV8Ll+7qegv
teJQOvrViEof66A6OY6EX9Jb2GJ/P6mKpNMud2KMr4rBb1+2i7ei6BzcyucLAUlN
JYHLftz7zmBzLNKA1WaQBbOhP1c9RrIYLyp25FUnnCtX5XGJG2wkW8q5yeR8Wqbj
PnVbN1pPERG55wv19SePH7YY6nEOGBFew4JOkyP0xeHKj53WZhq60rlliz/EfHxt
bqo/L3VZZnm6UpzqpxCC1b3L1HIECH7J2hPbsGWcEbXMwZV3UclQ+rcBcOvpnSrr
xHJMb8azbcclEyfvaUk00tYr8Y1tHbZerFT7zc6BX69uV0Oc7AHPxrkTaxoAS2DK
yq5mDFvZupp5b/wfrY/gJVywakJS03RVlY2rd2hNFBHmCNYRw0m7SdV2uMjlymld
MCg5i5XCVCdv8zdeCgnghwrW41OyIidLZa2U282ZpvwNY1dxV4wUb5zNMjnTZCOJ
OsWMGaLbhf6Ox+MIY4OALuD7QX55zhEpMGcfptAYmyoYz84o4UW2dyGVoKLtrHQB
jMW9WSD1SN5L/17SJxjw2u9ISdOJDxVAMFCTc472mLNtfFNzfZsgzK93t+lC6Uwq
jLpTKhNxx00QZKlIqluxDF3/EyLllPs8mgcC38m7Fh/zIV3tyfKcl360ked2VBZk
UElBYRuVaAmSYOKGIETlWgI/rVouc9OrXq5kTk1i5zzoHoGhXxe1mPafL6e7EGZZ
+1lyuBKAL0BHfVy8wCvwu9oBmOUkTV4tW7FOxc0pZf0EWiSN7PJFy0IuXRUBwexo
3puLDlog8CD8OUg7r+2XH4lKvp6ZHGJvFdeRA7XWp47QQk07A7CK4yaigrqhsAmP
U4odP6dItowrJy+etUeQjtDaQQyDSSOaH564dnhqjx96RuCXIvDsl5+oD8zazKts
r/6YgFWI3W6MFFwOGG0OyH4/8TM52wRVA6remuaGmqJNeFr8lkWkS8w6cPhlRb8L
9KpARNWVON+jIDWryhBbZks6GVS9CNGrndb27uv0DnVFZU4eW1lFMqvt7go+8pbs
mDy2MoxWaLuhO1QIDmYAKNvBiXOEXtUmjGI+c9v5tY7VGNxCfbWQ1o+Faen4Jz/g
DiH7m1H+S6Vrg8ynXy+UFDa55tfxyFJIcQu/vt16Y5dR7sjqJl8UskDwI0oVUVCD
FRvVY2PlGBjAXIA5esxAFlJgWqFhUum2IDUalYPsM4E9evXbDH3OxGZZDDJk/7nA
+R9H9EvhMHk6dIQM56L/lo+tIspJ5yXcLvy5pqMU7qzbYT6L2CRwCltiU64wAROM
RotLwcU0RalCR9dUA7NhHc+mRjhbmiPIkA0mCBYhLVlVbpJPxf9p49rjxGId3vuG
XnhkKVNe8K3myrXEo7eJIETqzM0/rR86UT1MJ1te5YQxThBRR6XzbP2gIryrJqWN
VP9SWfd8FhwEi4FwwCsS8ZO2RUtYe1gHhp+Fuk6WW2wCh6wfK4ViAAjwWjDHSwg8
QRwo51rlnIoojA+3/FzuIINuK7DH6IbTHL4xLZOPrJ0OvwumW8xxc4ND17Gqw6j1
ETWxV/tS03jmNOBJfV742U0CXNw26wreS4WkNSy1YUhG10wh4QvHoj3beE0HFSc5
nodYfGzYRvuLoOL5+ikPLqPTyCS0PMqvUfye2v09GxJaygCXIa64f2eRAsjyoQti
FIymQ8yLGXBEn957S7XgTh+wK7jpiYw2GkwfmPbXWZFkG5TlyCyKONg1pU9YzuEL
7/on21jFV1IRd3maDvyTeuYaCcBOFU0TAFstrBHZn6pHZVyLd3z/fo4K8q+YVjTb
HU6GIpkJhCNnhoqKyJHmeoidBnmS8nxGE90yDVLcOhUQmpc+JUGQk26h223HzE4W
hHuuVA4UlXceUtnO8KrU+G81mmdMR8gU9t186iTK1vlMquanLA99rgxUb4ozD1/i
ZYhNaUrHrVItcl28CmqostvwzViQLvD/rWE2hwOdZJQiLmE4fl4XPtx0su8kW0FJ
gw2o85ZkeI4o4mKzDpJ6r46vNfHRbc4IlNilNFq+3bNfYqmJxMg1bCFSuVwyj3zb
E3ZK/+gNCQqOUpkoa1IGEhstkccXhpWlkInNO9HA+YMaQUYaWbpunQEIG6x5Z0L5
YBTLdiF3v3CRCgHAlgRcQ6/6gbVrlzpPUcCdIk3anCqVkIq0LuHG8XJyrPM/2boz
ARI/+Cu+lDDgq5u12dSmq36jMbf1+H9hvGSRaR4HKO//l60Ik1lc9zVOLVaRYlJD
NEht1pAquIjirnoiRnU+sGTxn/tu2cp9UjCbef/RbEkVTBy9PDIs9YTp6LaM6kj/
hvBzQ8QwyKKXJ+Mnngo33XZXzSky12ByJFJu75Z2gl5kjDuen+4SmgkRxK9EZB69
6RF25J+9A6+JQw1QV5FEnDJCgYUmGPo+eb5Oj1nsAcUNDoKkf+3OMRnb0kZfN6ra
lx0z7kCNLeWtcqHVHewDRs4v45ikenNSsuYxgurrzE/BAz92XHlhCc+9tlNfqEEH
D24ZUPW30Rz13fekY2xZ5FZP2VlOxyppmGMhhsPvmVhQyd1HHa7/GRLpqUOZJLnv
SDQGl0ckP1d0hTRqLDl2gXtFjzRaMzR6CGCDqoUJ1qLPh6TVh2ZI7m166RZ+L123
pu4C/eVxWUV1nxEzKiyk+r1yT39kTQKtKbYIeW7zQ4FrSRw8MVy9oW2+po/5wqKW
BsQpXpyWmbOGNE6ilQvFszB9VDTOpw9nskWu5EtB2PolKwHfItGXrw03qaE4nPU3
WC8t3tpwblmbkZlaRRhl4ji3uhPj9kNyzb5w8GCg4fNtF3wxPEbyTrm4ASlVbe1A
kLt/IwYE5PqMCeOUW0giMx7x/bjjEcerGVIzr2IZXYaR1C7MTIi1SaRG+rx3fu9b
HzEM6jDfSX0odpN78kyfqqCUuRAISDJ97B2xDDHk0xY2ogViyUwkBtKG9EJwZVHn
JOT9q0kDFkUaL3E+DFqQ6GKe5EVfU9dDKTP5zVh93q3FADQbfRO3Hsr7KZnv8Sb/
8btpqLRi1sCSRcGl9rVJKg+E0aiEfjCGxOfetUznYxDCE8Sxdn8V6L3bQPb6N1yT
ObX1xxCA/oniacWdGY2mlifJDIhkk8mbsy4t4DhWfwDtmsEjSPKFnosnPfEC5DoU
JcYr7isnMM2vqHw9iaUWPh68C8LXrnBhHN4qVsx71f+LGPj0PfttMkDpnmMe3ol3
XmOSFiUKCVq5Xu98qIKdQn3yV1z7CGvuSo7dfllX94sxYAJ44XEEFtBt4hTsFcV8
EvBjxZ8aj0hWSBwxRR1RyqFL1ItYQMevPE3Unvhhaf984RctlG0M/BQKt+ReObfm
lITzoU1An1lzyfc5O0OTGEXHumshtDnjBAEdzKEDOxGh1Q0z3MjTRgc5BB4ssKM6
Vkg+8fv65fHbiO8tEL3oRqJRYlmmoj8nNuK/wDlK//ZSQl54zDjiHH4lpg2DVCUT
uWe8yPjMbp/h51lfptjHDsTaD+B3gxhP4+DggRfLA0IYK1gR08YrXgbfWqhR09bX
eu7IGA4ynaI12mMtWZXwDdcd0lCFNlrJNV6TASFvK49tOiP8ACqIWxu3fbEyz/Jq
5b+bLP7noqqx2ab38Xb6Xp+9itqJTdiJYbpjXS4A2ccTk17x86zUPapvapti1knU
NZD3hxw1rlCyFEgSDJVgaAmEroquEtRKPY7CToj1m+419e4KPvFaFEutKkx0aD9n
KlFPZD70tcWh5T6nrfb+tgkU45D8w1kImI7GfNKr6aMoYTaEguIbtMlbnH2N42d8
ATCqwc86NxbOamkcOmm+FidfGOlHYlUyXxvRDbE1x8CX+JEOUXofLMzIhqzLw6Ph
epFJig49/gOiP1LEoc0s7mWNPgAbLotCgdV/J7ZSXyTg+pSyWVpPmQBTOhdkFJTF
9SWes251HdjymLbSVtc5FTH6/3hurUZQmiMXn+PK419Jvi5iyvDzmCwRozrCdm9+
rI/Z3nOjpdUEkO/yLTxGwPefb+HP5l4yJv15rLxcEis6mFgM0vC82JAweiBqVIOG
2OFyfACW6aOzkCsehfhwD0v68xDQtdyb++k5kAX6Bxpq8akL2OPdYzBxaY7iyxjK
l2ReooTKuzaM5JndcrU2rGZg/sFhhb6inc8YYm2imRW2UcAS9a30dZQIV77ivdPc
+kuSNNRiY+gTOy6H0+VqCthoZ3skY6z1yxMZsQ2BzIxvisWe90GIldO56po39NHi
O6c+MRG0FWiuez1Wy4wXbWx/0jBjy1D2PLmY6kkP1Cmm5XD1J4Kx0OneMUe9vvva
fkjKA5OCVjgv9ihtT4hAzxdQ61B4fYSUJLZQqc+3/J1mWq9zAPxwieJ4ao8fWffo
6S/WO2cYm2ThWgM5E2lCXm7u8R9TFKnnNHh8hY4ReYrZ/Kf0UF3Zi+5ex9a94y3I
JJhEZCLmF2ZoJqkEbOa+BuUchAReOIc7IIedv84KHNkpYZ/q2oROANut/8cMEcfF
vHIxb0Gqrks9gtwNjSqQT4rADimlpHZLJiITmZBneTa2eEn14j/o1RTSwr7IXKb8
w//0oU02mP23lPTZlFIPc2EuNJ11XravBnqGNk9jGg21CKG+AFO9cs70BTu/KASX
a2CwA8FBM9a7vV2OU3TYjaEO3/qTqIqJx9K15xSBkMEWXmvcm3WqDFNa9OkawgZ5
WFUPd7jOMmVvCUkR6a54PrwrEiQPryWBnpMFt3dUAT094s0vHaMrHcLLRW9u4XuD
TsGlFnMK47Ewa7qPkbJEqbGb0tfROe410wYIDx0ODQngAzKFMBYGY/xXlmgl5AGt
nQOgujJfKPJM9NOcZiajmN3X+eJs+XBgB8wYf2USBcKafW5DVKOB3tIgGMWEGMZK
RpA72mdTyI7J/E5HrzB+lJ+s680wnCJGin8gs3fYBHDFXncLDX+7aV/WS42L6mkI
HBLEgr+ttXDwKuQOcWxQdPUej2bqXUq0F9vE5yN668cpnJX6cElafmcZfxC0xKAQ
LaxLvaXBfIXvFUgIsHB34165tL+DN3ssHYMcckMH2+WVbaV5dZUIxWU4YUggHX0/
agB3Y7wrB7O+G/Dmi+BVEHb9cErp0r61UA25mBGGgcAJRpWzKnilMkM21a5gTnyK
2/gI7xecHulDCw+InbwoPY6rU4Iu3X8ojEPijcU3IpMeAM08fdmkBBmgX3ONMwwS
4ChgcX1pGVvJvKtAU47WKpB1fMV8Rd8jU3kJMGAYR8VS2FUISkQE/VBRIDATlSD9
eGrT1F54/AjQEEjbEKgF/RbeMOgH7ZRnQCQyye9J6JdcIN+kbq5A0YA/wFvoKVOo
nCHmKNVQlM0rJ0YoqL2+mqTQJ4OQ5VRxFntzh9J78vH8IN9NQ/SGv9kzgkzveZs5
ENr8y2ZexyJ7we2nFL0y0wtlToO2BH/0LJtCwClgv2LkAiFOFm5JAYubro8XGqx5
/vjqqR6mNmfV3bOxVKGrNM1rkjakF02kuPR4+FhfdN//t2Df8I9GBnglj56Pubaj
m1OBu4SiSovSn2+SVb2QWSLHWdCBYvNbM5Xdx8QDa1wmcyo3IV0FTiDbdNhxSkhR
FLj4ZiB9SiDbSrp+atWumMPm4ZLzqh/tlRJWSAtLsFjeS3WXP9Hx1I78wT6XKdyh
YKHNkw9B4gG20nREwUk7kKgj586QD+jhB4hnwvF8nzhFdgiLaCNRvJIYHXTKx60t
U0BvT3AeIq2E3NWIMjHAdXY87eg8qjQt9TTPhySwus3bSZH5gmPBT2JiAcTJr2hF
Nu0Of0+PKBl1UM2/KXbTUxK9bXP9n5jB/drBiNjDjgeHFW3F/EK5yy/zgdkDeWba
GGKEBco8qT4A9NZ7ZzlLWXpNE7hcPkB6BQbkoT/I8sjTABS3OJEgIEHj+GC7vwv/
CKNY9ZgJtp7jjsXOTIT80MX32sk+J05MRd1cIyDOY4jR9PGVGJC3wHL8I4cMp3ic
/Y5UiPP7TUcX+e+Kf6YamAjxsZUCIJJPCNYp6+f2XnVQsPO+bDVCsLuoHaF8VxPZ
DFyK/tExTu60cH4CD9sac2WlgiZh/YKppqHFZcatIGHbBpMedVtdgzM2eqtibgnt
oNYZeo7ObdAt+e8IAmUB41De0RtxTKD1ec+K0bDMdXe7qzUOt3kLBc2fTwvQq2h2
uK3tOHIQhi1G4X7++NTRR6Htjxpq/RybG09A44o2mU04RT76GUUxuLksXJ7RhcBX
+PN47CCuo25My9h7uHUxQT/EDdmUfJeY2x4BTDYYfl0aOdowU5NKBzYOA/aCmTEz
RIhRssNUFRzCJ+piVrZaYtqYtKzOMJXwIzQWQXtZxnSkfHIH5XH4/pSDFiP7UjRG
mvrOElqmrndqM/nG6e2v1z/Bnox1dWpoJB9EM0z9mGgBUxMH7QAYDODsqKonIWo4
qyaM7UkJVDOnnSmC/zpBYjKkqy33x4f3mFsV9vlZEXpU0KHmeTWpoiwI6L1bbyZM
xhaXuirBu+h2CaQ2cLlsWhbqyZbP1vJs4VQMSUzr9D9JMk8YkGIl53aMsqO6c6Td
q8e8TxAbTOT6GWBPBoRqPxvdu6BlTzKlyvad/d+a2ECfm90dGg+8c3qTwztuG+E4
rQPzR5bMx2fPm/KJITdur5unHiEbsInOPl9BjpSj4oFNQe6x6Cu43eweX38BWe8P
vg/2OlYh1eTMTo91BvLjQUkDkG4s97o4Q3ymHjLCEmfvv81Zn/JdLgwQ6PlFpSVc
l364r2C9eGK7qB+aauwWDNQ//YR1JHNXz/UHil0crnItc+k8ZdTrPYwxdFpKw8x5
RihuFxx7CvF+WLKERXLC85RScf4BoLBDh+IEWJxKi2PVYIzKniFBOtRHfHqwUwt5
MLUNOXmqopsGgyBGdQp/T5mkzhdur3e92lAbO9K4TJP97yPOXxCKNuHKdaWzvfyE
V7HcCIi5PxKizhpV33tiOH4+lEe8k7EMUkUas4JXrt7BAJcIRynN9/lGINsRoJJA
U+KPiv9w0hVxy7GGvRtRcNstLxG7uKLkrgD4jreLtNMQ9SeM7enUWYyTaUBKJb0T
M0+hzaeOk7ylJs7PJtHcrqgCxkYltGLeKZ9zWoM2XsCCi4MTlF30u4W1fvlx0R/9
ymU4XFQxkMTjAxMWZ1aB5lHRtXoABGSkDWD8BHKUXLZg95Kc0tEJIHBsFoSG6dp+
gMEhZ34gu/Zqhrd8h1dyKwXUD6rogNx2I9N6MX8rhZHy1bT11v6LsgGJnWdww44j
KfDA2Fjdijs2lfTx0bkcLFKanxaYK7520cjMJGGh2n25XP44EWbgPEsTYdJbOt6W
Q4cwVNgr14/3lR3f2ZiK7EHVNt0SeuzacDdRl7wJHq6S+ZLwL29iob3SZV8Q+Md9
VGG57xa5+pfPRgZxOHGp7CwI5AG+2b32eiqTpzlOhrL3by0FPsjvsmpTTVH0wVrC
Q3kfGH97iw4QRwf0b86KY3Gj/lcZx4z7e2j+npLkZ2/zU108yEUGdaseiCu7iOe8
ZveDgiUVRh2kz7m1OhHQLkGYmkpapb1lPDaGARbZ1mTW06a+q6bBGhB1loqdvLoP
bXpBWde5KClNvVZr+CDolRoYp9u1Tx7cVn/TK5C2RaxdkJ5mIEe+VzqSyf9ln+2Q
B2hjv4DVoSZrvGVcP26Dc70CV2Zf5i086IPw0jISmjnQEI1K79AX0aB2QlWeA6w9
Bo596JXlO1IEODupNAhvlVLG1I3+ff7FtVKj4I/8tsuebxVROGfHGmUq+cm/vP66
3MxopIQZYsV2wwclFNL+be0LZkO2nrU5iyTq0jJXZZdTnf9/LQJfTRu1dyys96L9
VxBZOzq+zqB4XGGtio+Nukmt8CvhbyQHVDnw55Au831zZ6kJdQmnofMt23z48b/Z
cJ2VXDE9QKV7X6Y6Q3SlM4foRgblq4pireOp1fH5Xbhx6ykR8T/K9a+Z/YqsGN8Z
SuBaJRylC2Cdo3xCkttZ1VesC93G19EcWcuO2hAYDkWZSwGcdI3u4ccm5Ut4WsMN
Yw5Q6KU2UDFuBNNPySfGF1rsluYyv64fM28FR5il7rYYylkW2BAqwi1pH3rDdZnR
rwl+P7H2fQTSavnHOifsqXA+pXbASrIrG83oyVc300WmPzrie4No/Gp1vxmWZlRZ
ZPJrd42uKg9i1mSHsBN4utB9Jg+aNOTlEtxHszFH8kllvQgmuwEERPdy+AAjbQAn
PL//VreqgrkJw1Grq0CZrjFR13MtzcyvHHkM2MnJPgtGcE6axNtqZEp0GLL11WSV
I+vl5leMR52gk6FeaA3J8qzWeveeswMUjcWvKKixO3l6XuZ9HTcmOozmlNRiNMAh
bsooZS26DdwkOAUbBEdPz2VVDSTaaQIlcogfi03fIlBdVxQTSJHRGMnQH73kvovV
pDHkRVpoKlXRH9EvQBOhqpAP55Hk7tn8c/ZWP6vDiPD7NNC4T5Pwi2QlhQpPPx4C
WrTpzYN4h2H9i3NtZzTJVLqHsMBG9axBa4TXDPfE30UDo8cv162Va85W0OdpNb/n
66hRf7y+rPyE9d6SMU9rF/hPpLMjXfwlzqgnh0I23naCaVIyV2wfooufxUAhN6Wm
FAEY8HJjEA2GdoJiI93OK3CkuBph4cnBkE3grhlS8iB4sU/1X8aKrsXvEfLZSQmL
rTw/+2HWX741+/UAY/BUCajuXWCjxCJNhYh0gpCjm76wXJ9KW8VvsS7N237L6xiX
qBaSFYupcAj1QuVTu7YXtxnUYWJdLLdbqyQgi5l5vpOTiPR2A5t4gMkhyzWC/xPj
vSuH/MNpG9ay7UlgxV9v7rta39W4Ho62ANmapE14Cj2Ct30f62KhUmraip0aiyxO
AVZ/sRb5MpQAcjk1moSks1klV4HrHTTyQfhvzlczPM2NrtqyOmGPLUaR+nCO/54R
S0XK2XtxUFvcTDhQio+nCIOftlSJXmAg8IBRI/dJeG50yC3UAF3aeUIOpgVcyBFv
2GG7M0G+9o+TyYeFA7jHGV2+wXOaTxbYnMi+chHCjRo7+I2vXDIwGA7njZa7pRSm
CD9DOFUzmoKLe44FuMNYS/+h80raqCcKwSI3hTcnL3UPZlX4nJ7U4/ghXnCrGT0y
jdiqvey1kJPwccYZFw4Fylv5/hLICSuQV7wDG+Bq87FKzT+uNxLFBonO/dWn4NdL
THIzeIOTgSUHWOC6vPixhjhMwxeH2il/AhOU+zqbW0mgsfma7R21vQVYmFYY/gxJ
iNkuEzCQ+0cRAvNmdO6TWDfuqCqbl7+lR12FANpMg5cUn4IlBaJ70eQa3QRAf549
l4wRLmOyJBPUFG4xC00jXhxzr1rp7OyKCfqAThln7VAMP4z8GU38jW8PLWoSgG0U
WFTtXyy1vncu/GG41zw6eNIT23MIk0Jg6tIYvega7x/163duWShmBS59YjFPHz49
RrXlZoJvzd601CjkBzNyrC+gjK5xnkAfah6vTVQV37m2hvoxjNdZn7CpuPZ+TlLt
QtLbdzTlnN7S0ym+niIG4ziUSko2ywDylB25kinE16V1NJaaddV69KC2I/JtOXz/
w8H6uYk2J8jCr1lbnlQrplLJlcZIJeOkxHhXA86SMaLvtmLwwRPgr1dRt9Z2mntK
sA2FxfQlg9AfHE1F7t0Yasyj+X1GJV94/nxxQIhM/QfPRB49HjGXIRO1bMXI2TLf
EO66flUlbPbPUBoGLeLptvrYVFFkTJBPmsVz2cS4lqoy+6e/3rC4R87fjEK9+eCl
qEKxmvwKdKZ6Jg/JgzpgKSdWckVgy8p7i9nPMQxrQHKtWClbmtnN2Un3eIIquEvZ
5E4xhZYZOZ9FoM299hk5SMcVsEIN+dR7babEd32sjv+OYC86andxvc7EaSV997E3
KAHsik7nzlJBNIJKbm0l3GgbrA4SWBOhYu4lsqHYTtMfaBqNImdZL61su/kCYi0C
dx2kpkcHoIWpdQqfYQ9FefQtIn2KDwLLEsEbGQ8PObwx7Yi/ukLHNSgWBB0kT1T5
3kVCX7h2JTWNLNnaJJJsJyA5ePFkk0kKOBzr6ppAvG0DRDsiYmI5KV8qkGy39COQ
/iV4m4yrbdID/xhiKMsnoDu+0kr9/gLGZb6mmimABB1Sv1hlHfqIRT7G4MZzqAY6
IDdcdw1KZGH/FOFTWhMJ5AtusA476DE4jJc3bmySX5Av3UFLaj4qh2Rd10iMdt9d
QwpB04cAe+eJlCYft/vQDnufDEwLUVdkES6uc9tTPnLHc214nfHAJTljMdgt84qd
zMk4c78xalL5KymbfTcNwhUdy7yV00+r0h7VVA4hiizsrj1hlvonZcSTdxxr8ZDM
QkOL5+t/CQIeJ6JkjLKv72tu7PMzMiuHO6+aGGopHrn30i0Y4dfbxbHelJ72p5Yq
EFkYEUcCWzxiq5WIkOQ1LTaHe+agB1wKvtvqOQ5ZgAlu0I5ryOtCgqdS/NQpDXOi
4Uszk4cu0oipU5AX8Ld4oen5ti0G1av60QRIQa4tiheFkbImnyKp7RViq4/+2fUS
8LpzqFPOCfNz27F8MdX9ZgxlhNRWuWGUqD7wnN6fWofV+UyuBwnvMn2bGOYe2rBu
1iVGi4V+MxM6H5jizxQcuzl/ZsOzS+CrrjbkKOHX00G06eQ5uQKjuWN+1FmM2PCJ
dHvGzWZxxTPX9cU48A0ReMve9xrfB9b10fMGQEp7xfycegS4gERwudhlgTWNHaA4
yscwi4criE/NWm43DvS5hOWwpo5Zbz7o4H6fSURh5+VXv8b2uxQ3EdVmiILkCLtW
fE7Ha3q3J1hZ/ncDHx4GwPVp5s4JijPxUIK+V4aECtMvrSO2h6+tVR1wiu0Jb0vj
AqKDy4Ayern7nPA9aJdONIJDxiuhqxSasgmzgtcOZs9BDUGJT/uqQnWpJ9pNCUG2
Hnssr29Hcsw3oVo3uxuXvKVychCKxf54FQl4zXiIohcrhdoY15uVMCuh4AL92l9e
ifpH2H903/949ZGHeyYJbcMeBtciYg9DMkg0TKpli6C8FXpWSXwV8XByi65+W2GF
R9lUCvrhki1mFB28Egqjlp+DdgswbX96PEgMh0dMFRH16hw1HbZLNxRDW4MeMwL8
J6nAu5XF30JFBJd2gxvkeDVpfQVHD6ex9/bKV/D+S1p+/XQgERtNOhYPvfyyNVTe
XsiO9laJ4e65TpAMgWqnR77g57vOTwoZFLjRY/JZnKkYyvQQPt3UmfQZY1Y/tQVS
Ziix8IyJuxtfviZvtsqblr01897B/7BCDReNxuJ2PD5sApVevan0JXu+EZmf1ZyD
pu63J5zVOof1kwpd0BkIr/PHxdPm2wDkNxM9ryH+yOCaawigh6bHuRZDra0e0yMv
V6Mcsa0whuMj5W+yfgN8UjzYg0PctK1iS/GjiBCZViCdIxnCH1YeASDSaQXdTa8O
xVmoSCArLiKYwmVVm2HjppIa9kSvaSQKR3ULrpdsJNDSLCy1YzOti5uQm9+rovPq
7wDsBxtczw6jI5Agxf/WQnvbYkY92HZcfxF+PxJ2X8+utpMIkPmIhHENCu6V9HbT
AXvYg14gUzBuysAgmZiNbmTuj/ELYt9W7rXNNEOq+Hri9lJ3B9pqrO5lQsYecxb3
JxcHDZquzxWn8iqN3t4HRmW8qgucKYYX4s8wEUJ72C9de2a3CJymN4pfWoO6bcoP
QD/2Xel27A17e95eQqDehXclQloLmn0/LEHPPU/EO3ghjV2Utw5OH3BdsGmWROke
6KBwz23JecxzObhsMHchBbZwMeYks9MMxI040lgVxCxJCpe/ouy8Iy437dx8aHir
3oqqH+jzNXqMePrkcNGJeNoZg3ZpI1FifPc3xlSlYD9WcJ4EIX5LSgZ6T85f+CLC
fxpVu+3yurjpJIJ6LSQzQd2/dxgi0J0g79EH4jWiZedIVqFKQcqm0w4QgyEQt3ZV
6I3zoDNhnM8PfMIgm5LMU/zZxcw8d82+pgrYcsqp33irwaGhgyR3kvMXFfDnk7Z6
orEyrUzgYRJaAM9PQ7RKJFGbW2YvSv7ojgsEpaoQcJOldMUCHErSUTPz+9FpkkK/
rRjODH2dZvpecLTwMEsxRQFHISMtANFc/1FmUI3kUbh5fkBV8F+SNtP689ORl58z
6gM+oVfOnlT5j7PNXp2UZx+mbEPdWzpNc3EXRlMLZ1uyX4ajjvY+LeMELXjCPnxJ
KIQ8KsBdh8wyBJhxil3eKJ/q6QO/VegJEaYrozT58TDiqIfdVIJ5k2Rt2tOutyV1
XH2VUSZkLUvrDs0X8ln1tHd/kBayt8+a8Xg2TEiC6XQg7JyETUozh2zfZumd4Jep
iYdX4pSDTCutcPsKnzUL5iQRPaKVWGD0geNLPtAyV0qTCB2tua9rZOQqHLahuWbo
zwnlzJwDbczF/LwRTS2lgOEJhv+LfxmDq5jDcZnqg0dpWx6TaVr7NKYF5KFtl0xd
juh2Z/R/fpxFBgArE80/HF8lOTtaG1yzX6ORnhkpj3d6Ai9VWzKOgGCW+QplLb2a
XyI+drmOB3af/faCWOYJp1tgjg+TF3qpLyMPHfagP4UsUx/ZN6nSML+93ojmibAZ
zChiRET73tWopJSArK3iiHj2ILh5t6K2J2WhynTaqzyR7d+FXUkbm7rqlbHQPwZ3
3cOWBEAzo/rH59simAg8NyyfD8bhfLXuotKNvVqniYBl1YmQhHMTP6XFKcJlcaUM
PIQiLvJJqE94puXPVTblcIoP8KVrmbX0qM6oPeKQf1flYOTeglbhT9Xcw/w1gLHU
m38DvoPfPPnoFSUfvH8/GlUs8XSJpf4kZBNV9GkZ2jIIrDWrOCBHnxvzpkzXV3u5
u9fVVB173OPgg9goGkgPJUJjZLSY5/agHa07pjAH1HxbFejDf+//DeGbEWHv+YUL
DB3TpNSw5KcDt2JZHsXHs/KILwn7HoWbG1k2asNJTBuDdhPZ+QpX0QJv8aCWkpmk
QnoAl/qXnlIMSvccpfuNfJTTNoN6GbERomix6ZntB/Mwxs2XHTiuqLDZatnebxHW
wkdBwqE8k6OWhCFvN9AWfYI2z5DvKTR3SmXlUzDsZjsJjvjpCecmQ31Hp0TP+Bvu
VM/mzOfx6C/5PpSzDb3Lut9Wwgj0kRexcUhGE6JSuN9cPe4xCWLDAzYXPNOe1bxm
cHvD07F8TeLi/C/vhu9thLGmzSLDnWaIWlyfoqEKbzDXoVDRTnw4gWUKxu1Milnb
S52CuDvtHwXoVxl7bvCpPwF6yFiUNLiUbzyJwhYQkppUkINcrsYoT0mJGZ7U2Khq
GL743XToCWvWwGCDdPJDWR7kDeGie+DTgC0k7n1uhnrFpBnzxI4V0tZJoBbFAZO9
mlF0BdB+ujwpsyIsZqtTq9cc84ZvI8cYZ5IER0sKa2u6ST56r8fWFGszAZVUdFcv
fC1XrPeH4Oj7mQTUPLeb42Lyy9i/WXZShHtT9sdgNEteu4Ta0Zne5wulkfy6Dqve
aY/YR8IuFWm9zd+0YSfkgu3AKuTZEChPAa462W+ZfjeyjUN0zwYJc711rlFag4ih
sEddJ88p4p8fGmMdHwYAFO8KM6S6sMtaJ2t2vdsa483mONCZO1Fmomp+p8fmKxEF
WJWlAunjewpnfFBCnKKI27DbgkRN+/5BkeP7c5INVyMw0ZSftto13N25BaXJ+87m
ZSv0A8hSc2Zdm4jhpALnCZgdhs+Ch4soBej9wJACJB3fnzHSaUfJyP6Moa4p620B
eCWAPvvR8UheKghbLhT4dhKoU1csqjN5ge1oppbRJIfnh44ZNlmWQRVPSHyUhnm8
fsLWKKbYwGNDEHz235u6XIpTq9zp6AzvzX0ELPJ+nMywIp9v9IgkgKPA8+exL8FK
yQBi7lcEAf6ZF2Q1en2jPsq0uywWUkE9AaZvU1cKC7XB/0girK5m4WnoSwkHFclQ
5K9nh6vrr9YPfoCRtzO9bcUwjApwfJ6gCsi3gMfK7PbgS29GVEe46cXGdTj5ds6n
OOhL13aGqqMJXKSPdnpmXm2g12FiHBmdvYh5+5RiGzjoY72gy/Eh95rxIjxlYpHo
UY1y94xwg0w+oalJI2AtBF4CK2LTTuvKWyi5nOW98Sr1Lh5UHA2D7/kIZL11IlSJ
A1IXH1YZ5O4sD+VZj/jqXconXcUuL60v6KP+qBq1ZGk0jFJvBZMaP/H3RyaHt8dn
5/xGQHThGGmZSHkmU5k7iS2IR4emysUM6ifjCg60lVRmBJbXwzVvhyoa//rlEYE3
iJDEaP7Xo6EYqu9qTV65kWjudgtINSKBYzIfrxsWMP06smnyktbt9ARIbZNu4T0N
xnzq+iQ1GNrqCYvYxqrbHBCSu8k8Up+pSu3h0R0Bl4N0GyDppRyKUqw7bJXz63rU
/y6Q0swpt3uo3LlAvova33DoKC0rF8D7kVuMuOPhw2shQMP91S6+mdnrzNBut3QC
wdW46OgteiLlU9O5pYx0TyWArBVmzZNINpLDZCddo1jL1h3cW3o6tviBX7fnMSGk
/ZC9wnoljB9mrRF+/rE318ATeSR7NUX40fZdRrg81MBYj1kGC8juwB9QPAiH1Hjd
C77Wi9/L/Jg66lQBQP/qLPsvifu2tKpQoOH1myHHKIB70gSH6JYtmoT7ILmuRNxO
rw23ts69FJtKgP5zb/wCXEpR/AplaSTjh2J+8YqYUJk9TFckzHaAAknWf8b0u7R4
KXXlRr+0ojlm3CxxIT/PqzRt3OjU5DroTLIUPawK+6T6fFRx4sfHD5FPUM/C9r8Y
vJdkqUr8frA4Ss4001jPzktponyMSgciKkVqim/IhgGDpQCm5/cOarKhUILa6PBP
A7U7vX+P2C/ohDLtHyhsXuC4uqcRMRc8RTdrAmRfsXPnGkXMcui9A/uCSOxtn82O
hPpEq/ntrV4mtQ4NMWKrsjgw4uRLIyav1XOz2oxcu5mfasPkBRx8PLLOXO3ngRNF
ra2Q9m1/VMsWtQPnjabOYGLMeeqZGR+HomuqGhlmBqRTqnPQb+umap5JcUg9ynJQ
7xJsqq9hI3HtjRyuBHaOxGbSBFdpMW0VnRQbZx8/BKRfD4vfCZpA4tGVNrIRim96
jEenwDq5TBvQfYQVucfGxoivNXuoDSLnnObsq7v5k6SIlKNc20ycddNmmYWqGTF0
Cd/d0DJQplwla1PNLfUNAC4PKb4X0TlE7YCBs69GZHvamm9PFYfLYHjUX7jnbhac
IwpCvVF5McMgggAoQwAUq4abgik4fXDc/9qS/rNpF9WF2dxIcmVxzH33oyN9ze5y
+AwFIxViLVA+faZYZu1dXLmcpaMnc95MGruSy4TdaHvtngWkvw8e45akIrZPRIDB
sN6pCEi+XLs+dUJP5a0yTCzvsBWPSiVYkDaEKDICqMYZjrMfmW33vH+xmQTTr66y
t2Z3GGd+7DIXmMdMHMfGuidsPNiEYLPtaCupWB5rtovbxJX8KAgA6ZI7Jcs8WrR3
Mc0Vp7kIaQ3NQdmItY4FT93jKsfEvFwuO6TeE8Yg+IYgGRr6m0kFjxJpgihFzJ3q
TvUpS27DXobnw4Os9oV8KCBRX/vi0Yq5sx0k7inUN5yHMSoHgGnHkPl84bZwW2TB
k9VgCsI5l4xrdpR9FiffX1rBU5Z+aJTl+mE3scwVhMd4ujCFnmYl8Go+d1vAvrIH
kIxFbBkJTezGZy4asOiHwnDzNP+TNbKAgXy6uhPUTAdoZFlLk8vIFvirg72TAdLc
yWw9/AwVBiE8d1hvbX8PUda450Z2Rn7T2jya4GzRMRrE4c1mmDWNCWoCV/+l0Ked
FHOIWCTv30JHLkh8jCvs8llxrzhi8UwVfl5DvUsfRGTa4lRXlxqR1b7O8u+dxQ2v
WH0sJKXPpuN6UZOTYI6Dfwcg9US4QdJNTTYL0RJZvDso8A7j0pRtopdDHh2IcehU
yKD94ofXOMbyxQ8nWuGTEGY5uHpGBZfkRocpTl7YAar8pyfufrr2J90sgYzY8Hxn
bKTpzC87OlhxyLzJFN8LiffPFbjhuBa0sfWrKmPhS5wCkyyvTKdduCFePVTtwoX7
RqiSISqIeEwd4k/mXi8NjemXZCTbR5C7Z3O1hlkAqvRtKce0zHFAwoZNcE/OWh9b
FCW3GKVTqmjx6+Gm/mAQBhpr7jnlrbYtlVP059+Mo7QJ04bnWDCkEbX9NaH7/wyZ
ERpx0ff78csGeNxAmYhdC8xzGD5D7Qu+Z1d5DNbhZ5W9chd3UaaD+kDMfvhlM+Rx
FeMlMrvozO6O2KueoYx+Y3tOiHpzRXmDIjDZlKh5ukjfhOV8WXjBoO3PfdLodDKC
krTxXseMRce+VTWGlmTA7FV8xn4um3c1Wv566bc41Ubz+lokGgMD7gFeucRWfXi1
VESh2mlcOenCbIEOWX+yQlhkPWOyQXKt0vPS9L4pgeP3XKwDNFecIAGNI79oU/Rt
rcCPeXXiXEBovTSkcIUU7B61MV948rUViPBKROABopeFNHUrGLgWZJqVHCa8O9n5
ZdsT0Apxg/SAsvJQnuQz5E7M3EE61yWWCK+jemXh/7L997nMSVadjNkHDCHohl8s
HSKBdzeibeY/6bhrcnhXYn490vjR6bePBoJRZl7jY4Jl7DxzkPyzJ3gmt4UliskR
+wlvosl1jJTYFuCwJXwplc4GJSGBEA/Q3UPde43ee6+YORd0FSMj8rSa1Lod5KmP
CjD7iQtwtSP2piWFu8+9afGPF1Drq451QdmNpQBadggZLMYWrMQ9ftl/mxJ2/Zbg
rUpaVDYuSCiFXHX7nk33mC9sJzczrJJ0uilWpl59CMPIZ86fMTQ6jQNhfniRtYvf
WddUI84EBxh9LzGwHIcUO2XxoUgMzQbdaP78HG3hTeh9EQzZGiplNANzzh5KwO5f
BB1rITs+ktFIGk4vcZO7ouA4UQCHrqNwjbnqQLmUcXcHnKp4J+4pBarkIqfCcxAy
FR4snnHFjndpFi4FoygG4jHDsQfbQUutQKgf8UePDubUydPdPd+PJgjZJrmYxzJo
fXfsOQZnbOLLOPiF9d3HJUrZndRejgwRIpuhESx7FWOn4C+ijgHN8Z8P3HGj1qF2
4/cU0CFHNcb6pvG+pEfd36zXMfckhNhMX85G0wZkAC5ve5FFfEZ5+pXONQOUq5n6
DEcQdTbx677IfeiFA9RhdB18EyRsM2r/qHNX/IG5BcWlFgMNms9gH/YGLd0BkwHN
QpG7HIBeAZZKry5ZlcFckL6tsJXDXeVW21qrnQCT1Pn4G+BqFLf/ZV3MpnK5kUFB
DKPsV3pXkybzaCs3HKalSVd6SDgl3KmYcjPhZdIX3zFeZNoZ7zWgzADS1+soa3lb
PHDCXpYDbVsT0FFxhG/D5LE3tfdELWOhRan0HQKeVdxqijD1z1sLrzHZ7uYJ95zB
OcF8uFzq3WH+5v4g0jBcWfy0E6OKh7mr2WAs7CNCV7k0q5Rx49GmYFrPz03/42Bn
Yg8XqQZ7R5+vZCYjWdSGjuPTwMNzj6Ol1O0k2czpCzAc5ZQz+OE4ooRP8EpEUUCs
Z3Eik+qvTOgJW1R3ZBWjB6MyM9o9hJAoyU4gkHvYmzJyeNGL9M2+peNBNcsdd04v
dc/KlIjcVrZgUVf5KoHqs0dOizQDU51203bz/i10aUUKRiejLrEzPCD2O3zh5amt
/83HX7GJVfnFjsuoN2YtxhwkgxmU8VBb71+BpE1LbbmTfou5QuYSuIZqa7sxM0is
W0+l3SmRXBSMUrqKdXfXpaUaUhLMKvD3tar/a087oLTfiqrkT7nkisl/UpEoKNiD
LXQCeOlZcfu5ky3Bqwu2hGhLVi17fI0F1KFbt64RfeyCdZ++/nsvkotJVFe0XjMR
JFY8Nean0QpZidBv+zt15ckEdla0kyB6Tsb7bHCTwatn05Y1gr7eirTrCCtmu9Bi
vYllNwNKiEcxJ5drHPztPK7bfqF0unKlZaE2gaygi6ujeCC6dPtevavsl72i44ss
nggciywjX3/MUMJX+1MzPgWRA9PDWely2VotkLl/903yjyn6i881v/vt3Ds6JZda
IZlRhqEoaOBFPGX8JxGnwpLUyVJV4jADViqFOXt68DP1mplNLs+X1TpthkaWAqyx
v4chCrxp3e4NT6NFjFfndkJPqXdmeveCQGPFAxGGgnk3Iy1bFtx2Wn7xXa/mYzIw
XzPUD2Q+dmT+7Mg8i95Xs4TRUZA9MBIf04vB8Pb4Ngqr5YygTXkLl2Gzb98kyYtV
n7LUQh0onGgwrY4gFxtZJTjQbHeVpnKNdbZrcpaZwJM/QnrDerFnM3DAWuYsfrrl
CWAdX4WEJbjxGSQ5MyVi6zr1HspnEqYw608bM4pihLVLStvwY+aR0Oi+tuXQ6ueT
aglGytf7mu5OUXZiHS9qt6hXxAX0rxoxLq2ygY9kyik/OFd+qKNWD0Dv9/0vLnnK
M5RyKHmKxXQ7KuxInSGp5xHSc6qUaaJu+rClqH7/6fc=
`protect END_PROTECTED
