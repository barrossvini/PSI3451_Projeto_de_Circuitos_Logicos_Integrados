`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5a6wRp+tm4S4DjUVHAYEucVknaJmh9FqeiOQ0XPWyWrEwl29wgs4PG+PmfHs2g4O
Gc1Jbn5w+lQSjRkvXI5BO8hVCyG3jLTUI2Rsyb6b27T9ocdOqYdIqTMMsJGwIfWX
vj+A9YLM2CCj3rh3B95MPuAf94lSrk87xt79A07AY7RPcUA4ZSK32ldt3fRUb5aP
4BmkAJGt7K8P9H0GHpmxY0RFoaGVSWIspgK/KhceXdor8o1NfNActvLeVOPokXYQ
X43DCMtaBnWSbHIEi2GOe1ozU9TitqCq71lZvlXjU85cvkdOnZIZviayAjohjsml
S9jW3VvrDM5c5IzcsINY5MAwAkAQnPz3uYsFlppU9wiXL/+g8dy+JehKDMfMh09U
PjovQdnmECdCVBBc09hLYlj6HUPSkfOhNSuqYerUM/ggIslsfBKOXAOjIuIvpKOr
sAQwCpqZ2GuJCn6RQduAC41zmm/oPMs7WrWtFTiHqIjAPjrwsBe1rVAsrjyHk1E+
xxkITTwsoYfy2NybNO/4Mo5bEOKyDVbyaNo7czFQZMnIWGZBbbyI+65f0XoVPa2L
sen8/4FT0+pgwXVapSMMmKatrHGBv19QwzwZS1OylAPIm2pkUNwGodpIr9xoBo1/
C2Nav291afNFycNLvcAJEo6f9j1t6NK/iw04/94rWwU5kgaQcN44Qbuv0oCOh1ck
yrcvi9M37WC3opF7bXItLQgFVn5Kx1jUWWncC8Lt6Ykq+SA0UEB0W8P2ZFSKRzm/
g7khZoBbNZhggn8kOiHpVzjC+7Q/Z7S4FzQeQxBcdYnAgMRHlQXa/kZBMSebD4Gh
On5MUWHC2s+E/xYn99PG4bWvGdgG/xDxvcurt/mbVfqa8Kj3JKir6Lp2httD2eIy
XPBpZJr0qwyjsJ6ivV/EqWeauupIx3n8d4cpN5sZ3bK8CSWLf2JRFds6lyjW7uKS
JHsGcCWP3C0ysSqSK+ok04PkFe7aAFT9lIz8FCp9+iYAbBFFEqm3E3xpvNwuU/nW
i77v0c8E6HUu/M2H0WyjNJ3H3oMNykvemrd+y8QlW61b67iT/GQmnYes+NBINuS8
cCxJNC9Fdny9kXiXkW4yfGkIpP4LEz0An+gL1tKuxmyFdUJrRHqFITXo09sDpzEy
w3qp6wLKobeiPox8IBv4gPdF7NzMyLZvON8Bbdi6dIhUTaWJOYznu6YFgQWf/+q4
dFnL97Iz6Kjrk4Q7kC9VQxlgcUi85ZCe+kKIyFi8lolcJ9jFCNTEKEtIz0+hIfIm
QJ7jgemrqLZIUGBo3qTLk6Ght+Bu92Mfnq2xIEmzcDkE6Y5JRubFffPZzdDVKrZl
O/8WelGiSaJahNlyUoGE3WjwZmDas/7X/8SnKM91c9MSW1GDWIaTpFyUnLRU5OX/
W3Ff0yhd0gBSyhwehWp78zxdIVJECOxLCBcFW+28LSwyl7nj7MoGkELD2HyybdhW
uEkh/4+nKecGRHNQc7QOtzLyXn7z0m5DwDViJJBJDq5StppdRInpjqzra95DKspH
VxvVIGhZPF/MyiyBIO2G/3vsng3ydAkafJEedt+O2AOKqAOB+SFXi3vXecFaIRhD
JM2XQlelyqO3LacaIJmD2LUnPEoSXiAkDN/nF/QSj2YmPwtw8RfgPIOrwkSokRzH
ulcGOdkOjt8xj+DNGM/TpI0f2l+jmjrVWzaxfsJHUNUVtZV80yF1aQww4iINLOV+
4yIBGtHi1IsPEJhw6R1XE7iDQ1z8Kx8n98vkNOjE+6umNkNDwzCZptkwYFtzuF8g
dHzBQqTtjQNt5tit+2wAxTRm/DLeMZ3CuAQocXByzWL9W6xdnXffcKX0sjSDMCk1
PN72XaVCMYLHBpR3S4Epi7ZEjJIF5eAeS38bG0lpiUa96JVhQ0BKdCUuxAU0eY8Y
RaGFHmZoiDcCqs7zhvSB1zfN2RspEvRvMf0/A9f7jME9fpK+byO3aZN1gA7e5NVM
FPPsCQT/P/gVUq9oXXCYkdccOU99xyXr5NHMxRt3WACrNSAXdH2ya0xX6OXgy6Uv
VVA6e/g1z7wXrHtve44/o3taNxB5EO4UPBIpsc86RKRAWfVQn6bCFOtJW44S/Zy7
K5xXb36yFMbTAFywGzy6vc81kEHBe56sXL5P0ZBrfNOqfg1IJdQp/hRt1OysKoHG
voNfP5JD8oH3jrLlRztChHCj86Ok2fK2CbEUYD7taOo=
`protect END_PROTECTED
