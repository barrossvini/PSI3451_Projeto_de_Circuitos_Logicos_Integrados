`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61SH1Eg4oOtQxECh74WI1gjT2o9CizjBwcLv0hs78HMivaKbAgHpLDJEpk2fvTLe
Ox3mEAeGuLLDmfUFGk76Sw/Xj/MgPqY7qcH5zBvQ5PtEpmAkOM5Al27Oa5tqHDOt
/3J5d4EEf3XLt7P64rkqQ8sgjyjmDVaaczZW+VAl0KRgeEOj3CONapWsd9rVD2OO
9pczrVLKSbvZNL+YW1Jvi7ZlszInKZz8MWUC3kfKylt7B31CHdVlQS4WErk1C2Cg
/SnfsUhIWIM2cxMp3bxi2rEhQCUGnmmR/XCR4xR/RXBs1C0snDuBIa8qYV/eeE2v
nUu7MdMvSf/now3tPq3bxobGtym7jx1nYYH6TeenU2hX1hkeYmoIw0xh8Mil9ewK
ovaPKKt4+UacZFjurUAHqPOr2BuUFjRMG/BjYaKp7Gd9vbCNpVU2dTbJXDG++avh
acQ9x57dkkAb6N46EcVRbzWv8kun6T4oVlpPyKcdp/Y1jWXqu/4EZJGBR98g31r+
+adfe45FN486EJGQKW+PClZUNhF/oeVAWG+/4KoBWMdQ+v6s3Bbdtjt9U7JLMuQe
sScdFVNQezczr5zV97JUEkUDU8TvQjOVxJHRIqOcJbSSerlHW+fr2nnpLdAiT+r4
nltSCs+Heyq+Je9JWf2Sx/LqbLN7/E74yeMSWUzeDMiroJGsNNB9dVcQClXVRbWR
sdMhwRUkQsRVkA03LyiZIVg6E/2BD7Kil5qH2YQokWbWBKyXaKHwPEyBPFBuYa/m
NNP0iMpHchV5h4BZT5yW4VriSFsORGcpM2jKKw1RTx00qiae/CfmgK4L5+Enkv9F
4XO8/UcSPEuvTkPaZ9WkC+S6JXpT6SUSljqEUbaWLx+VuoHATDrUqifomKoxT8k2
riE9EWxqFUVOGOpdnodcFU2WMabt2KiSHILOpeEeC+l81t/IJrdq65xPPLM7vCWy
ub7K3OgP8zSYBKrGc24kvojkaN4W+xnS0aXX9vE4Gec2aFJ3HZ9dy7bJDSL4Ni0b
WGXGiMosm0AXizGFCiis+J+z1rU+YzR7QQxRF0lUQhcd3AVuDcGfgSDI/E8FJRBF
2hB44iRT8zxdMIN5lLFFdDHIlnKfHMk6OMEeUniNm3BwpWOEWva7wFTlRvGHl1QX
jyYPTRa1uIMTEkYtd8DbETvnYZKimYw+/6xyN/glCGqVkJUCtrdh0bWFSQvlOnnm
VPA87zBiwoUi/JP0lw1FyrnWVi6P6/2WnjzWGsJK2wefT/to67se9MjKAB7GxpZk
LeQ9C7lRmLSqoaVyagwgkhMimPQuHj1pSBRQYn5Xn1YD7cC8eUjn35IPJGxzNhqF
s14J6gjBtuMdR7uebIIQa7NcZzvhRyBsxCrKvnrl+z3fbGWPaehK5rd77Xn7kzJV
Gwlr5LpbeEbQgAVmVYZgiBMSaDvf0XG9Njc0ksN8BwYwpBZUMImMAvDn/JTlaRcN
dWOij300jVqs3fL/XO92sbs59ekay5osDVyjFt9aP8Bd4qCHSXM7fItZ82tNdfhH
fAfnOTfRcJEPSmUhII8tIY9wpV4NGonmD0PAAiExKVfquyIB5SiXYQsB7qvHWtlg
CVNHNs7xvSn/7PNl7R7pOCK0XLu/geKQyGSi+u1eeL4g9vUojh2iYj2hyhD1e7fx
cxAOOnzdAqDeutf3EF++xqdmrAiVec5Qv/ybg5qcUM1BHOLwGwpSLhGbJcrc2v09
9at6HH6OzG3JbsN90n1xHMdfz1D4dtT4Pm3aLtmxy2XyVgmK0O/h9s7sRoZNkihH
uqvpsDk4+q7I1Cq/VcfiIwVKmDgvugDMgCAuP2NcO5Lz+gZsnr4zQgivpPqdTdo/
wTHCb6yJKNDO2+7FY3zZqJqVWSGKbdzT+a3OizhP2h88Y2CvJedLDZFRNS6RK1ws
t/TymcFkCpbgCsqxTuex5ruSukqzMb6cnUmGQ5zzFzs7Dx1xNpRbtZXGtF2kcsv/
pklGX7TH7z6tDhoE4FnZFZxCqK5FMH0SRswep+hJkzUtwgs/2SeIi5WHAyoMfyrZ
T3qgixt7+DeWiVPOpKRlG1pmENV/dLmAsnuZUWqQlY1FT0FjmUGU8uJR7agUl+JC
r40l/J51cTYrm5Z3mwRSndiFBgWxqcTy6zeugNs8MOUQhMO6gjNLVIf7OFcpTTvO
tA4eGHljBSa0Fw2OAMu+lrzmh5prz9q/ZZApPKlxD4i3hZh/i8AbE559n4e5YWR8
0O5L8rHVTiN7y5cXYBN+b1d8BoRYT4Dkk6sNRAdsBgn7GBZkMt2QAcJiSJk2g4fw
nmScqeSu53tDPA+dTThuK2psqFGvKB1bARTsssCsGu21N4X/0iimxjb5pxPVljp2
1vCRSCaNqmZBCsR1+EjZtoofKHyCSi0vBLkyuOdT3/IFwJw7gKCC0KaKb83gNQTM
aCzyIq13izDbA/VuaogifErPgdwbz06Lf/R7GZsjRKaagPbfUOwzF63CRIocpKh2
gZju2vSnZbtNGDwAJ3Y9jhxW/U7FcVEwCSASwo+4oGUga0XDMI0wphEbPKuoXrsI
mYT6TW+yusbL2UaDP72/fUGlv9XG2Thk1zAhD7RhZ7j4cN0hqY9SWXLu4/6J5n2W
inJ/kRF1YVfPqQpGDqz57CTqA0gQpAqYgTpcrrOXdrwAOmBGz0NifPz4EghUGFVX
5qsEv3eU/cuN1h0F/hu+xzOZlWCyulOmpTYVbYHvfYP8e1yuOvE7/gLRu9qS+uY+
ywZQKoB6K55kzIDFM/gD85AM/2rIenEjmVDW/PMKGgQEMp3Sd+NfbL5tVHkEAu99
Aw7FQhWho5PyP2us/0P3ZWjDHBPUru/ac4XjWkzbsFBq/4XiTYsAc8W01ZTunTQs
dFKf6j8dtHTvQ4ElC10ZnNUcXg+GdKYdcNjLMnn+FG2YOhFSCMQTz/kxpQEJMtVp
zztBBjUZRwz2VwW//NVtLWYvFVbsmWjqESMEadNN18tsNqJ9TJ16acyTwE6SY7wR
TKmXZw+RzbmVQFCpOlwWv/PfnTc1W+epEtdAW5d5VFbi4fVyFcTmbYJBxgP+w4Kp
WnJ7KJ6FKZfr7+gn30utC2LlQmbxO0Fd1h3Yop6w5EZKOaqyRL3DBU4VxuldP4G1
+bwC9pr7/D2OEEzXowaZa78wej3jMn8pvP7dWFggqBdP0OOPep1SZp3jq5moXtXp
mju7I4on0jtOHGy/nluqGUypmZYjQLBLVTMSo90qb41hLjNwatFlIlZK1aB/1FX1
EzOHHZZlHh+dpPOwowYuRVp20/lF5tEkjGNNc2ua8SfkGUUKmfHTuunQmgNt8Kux
RPvy8KBMQB270uEuZYZZy0lerm4X7UqPvMwGgMH2ShphzpPjSFOpWtPVTxd5W8p8
x15BMIZaN+5+IUtqOEsE91BWxXoL+6DV7+c+PLPD0jBWSzBRZSekt8IiUgxYJhoy
dBEAZQwGFXfGOx/bATnC/wq1MUIdX5UW6Sxp/scBAeKDbMX1TPtuZmMzvCUwl8Qz
RUuKeiKTkgif2uKu0Q+JzA9IjqqKkJpHKmH2jOA+Irxnu6WiIDNUSqmJc5f/QV9X
KaBDOvfhsvuibcivBMnpeE3jMS0hpNqu6cynnTnnvTecqKgh5c4WSaSETyPXUIm7
MBHlBidQElQmZBAbsCoocyLQQcU+ZwWH0XXAJCtLr/FIx/FFdtc0gsnzOKCO+Z0R
FREH5K6C/1doJYqZdrquV/oaK/KsFr0BVWZMmP+XrJ60ciCpjqPb0IJ0LeRPNBQp
GPZSvtHvJjcZGtErgLwgleKGZAVZrmCUWPtjUJEwlzBOUSC3AUVkKCgRqy2r3/P8
rri6cfvO4D5bUE5JhU4G7Ngn11Y/zlwf9SoVZbFTy/MfGKcYR2D2NequOrCZ1lGq
pAq6dMkNva2Wc2Kcr0A/vm84F6c4vOvG1QO3pw5G1LFcLZcEY0iaU5u4oiZJ8wuP
1pBoPRcbomdYGQe3dXAFOQYIehEch3AtC5xZYQzD37hD05pooI4ljbdtwoFlU3S/
8E24ZpSQwc/46DT0SHvbKf0sAZAagGH/YCwK7g3IannviRNgiyOynJjE8s8inAUY
OAU1t+iovZLZr3SkBl0ZIo8F1Er5b1ksCwhT9Wg9v+v83QIzU2yGU9iIjVAnuO+X
mcIaJ/M0eSRxG7S2CmFFNO7lBWDPeuJQBVyKR+GFdafkbPDvrAANIjNjbRcwqQW1
YHgdbhE9bDmrLTY68wq7XeQ6sPmDeFYzw9QzjLXl385mwBmGUNVWcNRML8hCE3dN
/AfOkGFMdcmcFCbypN8yLINoxYbUepv4UTU634VBfWyjWzPjgxdAi99zxDeXrrPq
nKYShFRFJeFLPSc78FxgC+n2ePzxBGQz02wg6jOADOtMptyHot6ym8TlMueSiC+N
BvlX0Pe1suLLB/E9ADHOi5ZQWYj/btff34nkftTNf7WkdMO/QB5oQGHtuuFcZtnL
koEfTlzlUfGoQCRlOecoGKoeZ2GJ47WQ3iJhli7+9LnTTba1S+8M3NQSS6JTOzVW
MnP/yOCrRvjdBJJSNGoP8TJxGM50MWvOJbItfllmaDGowqX7j0kfZueFsRIw/xTW
lymzoMN42v+k6+rV9f5LHA4zF93TDwx1Mu+y8r/2/jdxg6I+X5LxMMYOdMho3j22
PCDWSPUwe1PSYsHwjqNJFky34di8/xWSS/BKx5LzTdSjIZrA1jmBBJBn9bT3wnPa
Tf4y2+4hYsIdeu3a6AEEnsRUSXRbDx0O7nN9kXuspF35DyJ0x1mLe7Ao+DM4rEcf
Y2bsUcLl/0wMJzA6eSa2rl7g7tMhkQso7Wy6izwXeMEDmQ6cFT3wOCMl21UTlt3y
KRFlo4ZVD6+iE5Q/H/zjpldNsqrslTxlH0RV3qsJ4IWR93QyojqKcZycls3Doxde
bQB0MDjMEZLtNHRgrPkXCvQBp8a42xmCjmC///2BXtQetYijou6bFHyuzeZzL+ZP
Kqvx72+poLeKDv093iA0tgfAOu/Ddvf2JTA2uvyJaiA+aAL5whvTWScblRlcFN4W
KDnDESL9PtU5G974zyZw9oMfxH4OtCHjoYHuqgGREUOpf76bgjHZcsQpZ0uOw/AF
53o3QIGbizBDdCePRF7fNWQWOxGiTqo+c79ROnJHmNurZ4E9ynGIJhctEEMjV14M
rADeqdgfMJfy0gCuq62WKLRlV33KPoJLzL4g8HDJXuBCIh9p73EA4d7b9GMwIvf+
YU0jJMPBF6qL6KqdB7cG5RKND62co1kmFnW+vgFtnnVGIHARkDxoe4gWujSyX/M7
6jI8tr4dtmDywsBdOVUVI9Qfbi1a+XQSx018AXWaOlIY3rOHFAFx4smvQZ0x3Scc
DIPiBCzpof1ef2gCWu8UjNWjQRfXoXIjEYfX8rLpflCV+NuqT9v0xFpDVR0rbq/w
5Od/U6zNA6ya6bSQ1D0kbYLBlerjkUjqpMd0e2v74zrL2qofkg5EqrswuHVFX5zk
1/Z8ws1+U00yYeyj8xAbsYuFi7UHXeNh7BYi4TpSEfIAGVSCTGTP6YzpdsFYjup7
vLX3sLrmXot12guzzS6BvhIZT0BGoIK8d6xbzl9tOMFuHg14xNr2V5t2QJX4uOvS
wJGBll1IVVbgA99YBtP+W9mcATEmaobq/F2bsebWpg3mhRgLjBNx2euq/VtBxF4n
R02iNzkj1WMe2N194I0rURRM9MgtOQ0sc/FB0IpJ4ToiT0iqxp2guiJjeIc2bVo0
DWH3iHKulzBmt2NpM4wwARU1TrNEh2xy7on6MQsy0wjHk8XWkshiYh7rohRaQ7ck
n2kAUQDRfvRS5nr0xPDL0qA83bdEpFNhQ09nRlUVt+EMyTWrQhrcnGM7urkCoP+l
Y7rhQTZiHwaQAvyGwBdSQf3wXoVO5TLxchG0fY7ick6DX6ps4ALCGoGY/KJc1Iuc
28lll0AxhBWBcyhsPTPO6lc6zS/GkZVlk0lMo+zAdSOyZNF95rtt2nFysqAg2jrL
ciG6vZJK8zRENq/bRAZ/rNjqzATYur8Zc+747QIITAkxrBw3CYpTLgdZMIObDDI6
GLxnbf1VqomlHWJQTYKsOwr8FpeBIl3hfZj8oU7wAfuF61o/POB1OF9thJV+kFlk
G0vBtE/jXaNOcMK1PFpWt9hu456QscAp0Iv6hv5nZMjVz+K60Z+/Vobx1SYdKA39
O42J+zBffBcELT9avnaiInlfdNrXwpW9y//D1mUjODRbnykoitxBODQMpo/YQfjC
eTw/V0rl7N9NzoxprmRWaN5Y+RFpwrQL/lCEZU3aeBvci1aL1OJRbaAt77APtBfx
KHpniUFU7qdAQs63KzXthySPlXmKItc06OBrCmMxMe1tPsiL6vptZhTsQBvf3wER
C/WW4SUw4o9Fjms1AvxKEgdH0Fl8+ZOqNlQeJ5wtxJ1ytVmy3uH2tSZbgAE8fJ38
8HVbR8lMoRLsRaC7/uthFbC7rxaj93slIYNpVmvHBRlBPikL8vxq5ixDEVELR5Dq
Qz54lWOLefGBw/u+vHvACE9QtPLvQ6M2zYDylGpOvpcHqw0SAh9wkI+7q4jfd+b6
2d8AzdLxzlxiTV3mYF/AEgekfvuoTX9yfH/pTGrb1dGnszFXeGGgs3pcFbEkGP0Y
6m3TiHg+rdzyseiKFi9vk/j/vFTZ/iT5cRSie3Do/UMmVNqfO0aeCr+CmFoKWb1M
VHYVArHakl5Dg+/PpZXZW0uk7RJF+GGWlRvrU+50elnEwyF6jOeTawrIONaLHXiF
TBKBGddiJO3ETy7sl/lHVrnPXo8hJMPWEVJS/WkFQ4fKcuOjNnhxA9chBaLjV0ym
Rarfj5eUJOBwOMNthgf4MSHYDjTJpvf2/Q1M0BR3G4lahsrGnKwMH/4k9USZTOz6
loPZuDlouWLvMPMr9W2p5OmCf5zlOk/Uv5MLEPxqWi6tof8AErUKf4X9aoCSvcdq
khOmTfUGlQygs1+es3MpeThciyN0TNTaEMY9RZN4lrcMiSkyny12FbRslbUjkghu
ylAgSJSiPhuKEmL/iSK3PL1MBgTtJZh+lAJEdELNRPhSk/BQJOAs2tPQpfEVtc7W
1qmKHaeuj2vFvCu1cQw72LGKvy9TveAm5MEU/ESblFy8YZ73Kmpfa88xiPio0fZo
MVZ8Pdpcnz4FbrNp++tGeroxw5S34Ll7u04qjVU//H0tyxkyiv2MRQvy2zsweaDM
Um9ftlIb4F0752H/7owwSGB/qIHfmtV3lmr3IdomF/lsDneCdWXxH6DuWvmU4qPl
5NGE9GKYQcuGrmKtbpkAlQd3yU/iqAvwmqwi2Wh6SMYErpgNu6uALKpE6uACzqrV
p7zo8S5nHDhP6NJie3pAj1XtO7zCtpm+V6NWiSxa3CvCo4UUqZYUXDiFd29gH3xm
EQgEnC7qpxjE56nEzcUf5r448/KEzFkMmgkqJALlTUU2xa8PnSLicM9dm0uzldob
f6dwzBOp1ygHnGct+0NesVnLB/PBdKOWABS+f1Kmq0qmgSu/mVGM7wGssW4RZB9H
1anEcuN4k2Lck6rK0l5/trgMgg2ifOQdA1ztIHSCWggbUeXePvrWq9JMpXClSwrn
YztLt+84r+vJhoenNGde4sGBs2/IUIqlxzg3vpXd1w/1VVYPHsjPRHFOLMV1xjw5
jxk33rYs7J5rqnVtjKAzvO7sYQPk+AotT7Dh1z+vlmnxSBLi1+5MkwcXgTkw7ScC
MG+p2F1ZWv+/0nZwvkIVMU3d1LrEHiXjLxxUn+DBVhUZ2vIsjgXIM7cj3NGrUs0o
rZZEOfRVy7UGj0EQlHuLEWblqIYEk5l8OHJ7b6uw/QfzW5Tio9YjTV47C/8vYT1E
bv1lbUkpUnVKILpH+3Ig7xOEu8a8YBam+Pl1HKe8JGGYZzbzXv7843PaZYJ6vZCl
lgY4dRoSfFIxvepPbALzl+AQKLFYCpNX7H4gnIcid4auuvcKTqeQfBWakta2z4rb
ncl9VpuaY14fJ5HtqJb31ZAnItQThYGxMw2SY3nBB0niDzmxJefPrK5+ThX4Mwgf
kbOYMjucUk9lpQP+B4+AiWdC17VvUDnGEtclRB6+ZmRJ24yYrRn1hU+v+9PXFdJY
/weB2HUVryLuu7Apr5ZFTKrdJRHKZmkK/v50/ESCkw5ukAVnDQJHpzcBa3SfMNHt
hOgAbESHVMphaidagL/lCoY8L1flcQMy/V4KsAfcgljIHOyE7ftltiqAYVS4Kgl1
JeexuYKTEB41b7laxfhSEuHa7Y67AtuEOMR+iKi1OhwW8o0KilB1AZC6Aq8c5Tad
N5BAH/bJTIpRDmACV2fqcCsKJ8cDQS3wevgCoZljurxiuxKY+QDSRWM6PUZ7k0OC
30qO8t+nS5DhkXm6cJIDUfYz1fEFQxi8ZYUQ4hKEfb6i7A6ejCuULVUC1PYF8rDG
1WPyHMPyvFco7XUafK9OLnkjUxKp0tLf7hX0NwyevumMUhCeXuTNR7OjqRINWQ+W
XoyPeBu8tM1mwS6C9dsEb3EodR5zQZQung2cLDDxP6Z56qDIi04znFZpM4G9K9yS
kgkWkD7wb2EMEU/e/4fSqXkjTCAumdiDla4oPZ2OReoTRZVb4UW5NE01f1Srr5WX
xvYn/6QleIG6rba9iwKSH2JmSdD5WvgyZZocGKGvaqUVpg43ibNbgpqWQlXRhP83
BPF1Cuc8ZKbGoOKoiuTEAyG3C0WxGwq9DZKKKv2PYR2bt+yNEeFgfY3Tiu+lDXa5
b1ULocAZa/qx+X0MNbvEzicHaUfKr81mTmGHeLmnsGbgmq8fmqNs1U8biptO5e2O
ohlraiYRna7No1ioMtzFpXcxcPaTPiZ7zHwgOdjXa+P/1gdvuOMws3kPQNCxtTbh
PIZIQ3BvikL/tdW2hPy7+pXVzmLzm4Dt/VKhrzHGRyG+cVSlTKqDprgTa1Qs2YEA
PFAXhVQ1ApnXw4gYEZOgqV+E88dCMJ5w2rf+8rl6KSmn/qz7Xsw9WwdS9Su9r1fi
wJRaPWuE9PMQXil+6MS/8ZudKANHtpEfgkvfU+AfsR/GkVHxGn8ICel/4tRsrJxL
xru4rwbiFFCqZxdtgsH0evu7rVLWLlaujJzTUCL5pQg++WAABGNsQPCeg4QBcVKC
V52MmM08vEZE7+HsGd1cYhEyWoELxOS7ztqUxpvnLLGhG4e+ybqjWjnM5jFf076d
GwE1n9yAqmyckXf/Oi1raDlRMRDSrMWNkpv1Mcbk+uDhnZjkW4mkKuomdp/UaGm+
NZie2pILRotueFh6MRq864QYREQ4U8CaqllfBOXJtHgxeLpQ9UJguMLICXM8fqjK
FyMAuui9PtkxLTFEKiWl/Bn+Q7Ik7lrjqclKarMnQWaTBt98ox4j7+LZWA7ahKZG
/6PGEIfJRwRPwHKhPKCMqvVEolKKKGRzW/9WmfkzpP/oGe9ij6X/Zyar7ZgLxSu1
W2uk/NMEjLepVAzg9S5UvYMr3n59Rb0YTRJQtso5/JFvF3xk99HkLQyXlpoEUkmV
JctOpeOWb8EV6dRpFhTP87Jhd59ROS+XqTPAU4Jo9TYnvUxgQlCNWj2A0CAi6xk2
uYwEKG/4tWyn6TvyUq6oZa6OI6SMSj5fvpmkZ43TwmkUSIqpnilRpRvMxJQ6A81d
PxQGoc4bWi5ZcbtCies4yNVu+FJ9FRtQg2nB/Iv3W+GWpoLg8XcdOuW15XJFYLdG
En/hfNf6mesfM0NnFInjBZzFglG90PaLEOC7wRTmNScaXv5X2yYum/hiMp+eo8xW
l/i7nOyEeC1x8Q3De/N+h/LvRKz5llTj2mpmqs10XWIDWKXryfc0yK4ml7Ggd48F
sBEqxl8MjdxNzk4racm3KmKF+OcKUKaC4TUrpgovSqNnVVuH68GGhCrgAPGhdJBB
mCCQTfXc3DcAJQ+K/UE8PcwRO5Grq5REUPiri8YOON6MhwZBj4zomf6ndoLy4Gbz
ynptwEosIwrcXlZcguNH3rNJU6N5dA7drQATEmOCSyJmHgtTKeIVjnbPkwxO8FFd
i4aDjlRjo2ISsSNzfkeZKiye4VvtkrPeYQu4iYcJi76THR+nmogGf+F4fILbrJjt
wg8ADd4d1Hd6yOIdD/14pZj0bdA2aIU13qObKr9rnvGR19/VoKSmnZM/uDct00d0
kVemjsUJnecDWM5LqkW6E0vlTT1expUJSqnuzQxex3+vzH7x/lu7sNmdXL9GA8gq
uAH7RGme6Q85JHKDxncOQQN/vPQKk89/wlKVKodpmlgeyOdHlGmKz69EWK5epelw
1DEjAvVYq2HE2IfC0kpDqh493IiJ6x7Z6DC7Yf4FMtTunx17GKQlCFu1HzoLLYf9
Jqw2WG+Upgbc6Wy0XUwMGp/oN0P2CFCfuzR6hFBWn/jAO8af/wqQH+cQLvGawYMY
xn6TokMtpdG4/euiFaGCvrLShqNpnUx+5v3kgSL2eb+oygvsCQeLFpDqqZ415svy
Z49GEqEHO/01TGu6gG6phk0EUqmzYtah1YwXJc/Ni64hMBk9K9h91V01jIpjbT0Y
BHM/T0tl1Hai6ypcfIJ3X1wKYnuK1cHjmpig9VOcI0BkVo++aYNCeBvm/m2m+Hg8
XZk+jii2bXqblNQyG2qg8KZTgPpRQ9C+Dd6wWtm0vXX7uo8jEZYe0a/lWJLLD6og
E5FM9JkGJY7U4BJXTrUojPG+avhGZe7gtLCSP4BtlfkTbAlYB08dBja/A76th9mp
mPlKcV529uwBwjR9cDa8nzBX3PAOFB+GzGj3fmPr87IflVnnXFkl95dJZtQxjzBj
qI7O2gM/FEO2uio/8vwoQRfsZ3ylJwL9OJfDBT+8zaHvC1nWRIN9AHY0sk0jVQ5y
jS6NgDqhHaSVWcO09urFv/QTiCoJA7yOSzC3kzKqnn61R3l7nYr6xTqGIA/F+BBN
lqAHhH9qC1eK5y0Gai9enRbbivTV4LnoILqCLqcDMvfQTfgxuzOvaeYsm/Vc/5K+
jaGOUw1CmMRaSL0XtZHhr1GnVMfUCf93x91Df+DrtMnaSwWRQBdhuEGxlGkZdQCw
YXF4lxvXBwmDBHf4MxaEy31pokOWY14WSwlMMVZWJ8qTgGnhOgc/+RwYe6+Ij5ZR
dhsqnG/5/o6io7NZ37NGW+SrQaAK8CDwV2iVFKIYAOOKx6fxWV00hjfXEYvvDsNT
dtfV5PxbKAWkOP4S/yfAbAXVO12E+M1oXVIdAq7L6dIvK2kGDKbV+DUixXMo50AF
UaZutr0QNMk9+mlf40vzxqyUi/4vb12eiZT1YwN4MrNIs+FWrq6UJ/q5KHzsp+2D
bvjjHrGuPxI+SfSsKO+D1XsZ/5vZouFl8vSpRexKLIjh/jo6m5C8GZPiaHWGgLko
enZlk44MOgyglYSVlDwY29iZG7vcVbw83PHxfhzESlScNYP+3Nm1kksZVOcoFJqg
56yky4oGfMvwW45kJFTXmFmM4+fd7kckU0auE34XibUkTwKptsfaQLWzfnmugskH
cKh+jhpPQiP3H8I8gItleh/I45zilui/DF6kxaleoeYvKPvf1NixF0+OA5Ck0yo2
wVcMeU7uZeKJEgW1eEjow3MHpi3Xpol9xialYLuMutSaqsYZXBaU/7hIn5pV9bEX
v4KZhcMNlTZ8wQ6WWWDwjnsefO+v+Lkj1x2Roj3YO0B8W0vEvnvGyy2EP1cEHi9M
faJr79fi23Tc6fvQm7zuvw2ex2UUHnoVnI+skDFT8WYBu7NGfbFiOstktdha3+9P
2kidDYdxhzYMdYD2Iuk/sNkWIKC4fXc5K4iw8j6WJraX3Ji+uJK4Fr0/cwT7KqPK
RVsrlCZV/OCBEkM/7aLozZD6XRnbxkalHa03ohmpXN2oZ+56fG474iLECjN3fhS2
4sgJuerKSMRqbFj4fMRVDsOh0tgtUpdd04OO8848++Afo3Sx8Bzc9KpOwvIg+BQR
+Kzcvwog0D3Ykm7AF/cMoVbd1tTTpTkfNtIDGxP07wiZajHShuAGufYvt+p+hzAu
+mzeVjTroDqXJ5EBU7Djn0M2Xask7UZufHERGZ+4uh3kww2dTL/9BHPK/63mw3WM
I2zyWqE61J3T0PJzi4KcP9rCClx38AHOZ3hn7DPwhoaAwvsLF0VhGXnc5A6HpRql
x1x3Ef6HkgLjXqk3V+i0QZ/gRTnxxMvecMrY9oJ9fjAfcs+hfD2fDi9ccaoLeN6a
ILwRqUp0oU47k8aML2I/kaX2MJGcMedG2+R4YmjNI70rK9dceDHtgwvkFxLEabOm
EPgFQzkrm7cmxz0wdWSffnCccXQnpTSVRX1g+fMNpq51x3QblfH19u9dhnSCfwgs
QLXjvCAfvNBb4SADwbC8dRk/+S/681polqN5fF8ewxx1eReq9e6BIGkBbCUTlyq4
PPLS0fWvJpVXE49q7t8tHmGS2skVobIOliO2CDei3RCFPt1fXurlkSrNHErdrhqH
y//4RcU3S576ZbBD2Y+a/Igu5Fzaw+cJDMEfAXRfAVo5DGCq1v7Itj/YuLSgoP6Y
vvhgQMaTYUZ+pHcQ/WwBxoHTUOPv3lplZT+euzJYRibLGUA8nypMpu2eq3x6rCIf
hCnFqxQp40/Wp4Q7Su0w5WsWS60tlOIpxd50GqfLGzkt4opTxesTMHXJrJcfC7dQ
9bsQX7K5RQBXYoVP4YADwxygsiBpYMw9oleoE87sf3zTwjbgrb24CsvMEViMbcmH
g2QReSzwhfPDd0pq8Cv0tqSJ+N0HQxiw1qaUj7UNKC8lA7EzNbo6ELOgrHiYahay
xbNtgRfmlTT9FlhUVi5B4OhtJeU2gPiwVfRgDiQJ0MVjJv041VjgwNu5JcfDvkqF
+aUMm8+azToK2Uz85zVpbrHM/eJfaydaET+1fpEw9SjCvPk+4PZ7BTPeEZxJ2H3t
5cmfCCh/LOdpoPyoBLsTZcF39GhOrPNhkS36gM7N29r8QYuD5h0fX+flOasFXelQ
mjkOYtjekI4cgor8AyaLVoZSUObkmvBUk7iXm4OK1MdIEAoFq6UdLIIKGcwU6NUW
OZGMmfQL7MQMd++/oa4LninDFRPeUV6sh1DsoV5LwHkCSGNcil+d6bYYj2gHmwT/
20l1AIE4A2q+a9fR90sxpzvlmYorboil6m7UrJoRflqSDhS5Jab7djtambPHmACb
3kaDFUASQCjlAFfpv1yYP3UvAt1TS7wIMIDqmzI1OpzZ7FYLUWIqiTaVGmnOttuR
rEFj3cKTMtCB79zQv6MSqLKJy/cDLVApOaWXVVZdI1lxCIP4xTHiLRu9nB7qdpro
ZRIy5soS4iyPvc9I+JImEvcuR44y/D1Hk8yuJZKjdT57cjTu8eIZ654iTckxUOtR
GndOKuxbYqC8ekP1kdJ191v7bj5G13Ess/Sv5cFQKuFtbQW9aZ2LoswY29SBgtId
KfndtEV5A24xlCDVsTkuSKP81U0OHdsbDEuTXIhCqPGcdD25kSOurSaAJX6nOGv3
hwUdQibpgIWGMETjAti2PlOAwtPrQjus/H13Nx68xLg3aT4lifhi6hwSW77xNv8q
TaweOKU5BVpgaZO4OYeIEX1SrF8gZkib7bGfwMjpSYrdyw0h55Nah1vmG5cauZz0
p7bMJdlOf21c2YnN4wYm8ksWvQSgx4CDcbSrYDWeLq+OQzaIXqmxfVWWXjHJ2x4H
RfUXN3hw2zHtiqYOLSL2egdn9IJoE6OzQ2494UBjU+bAKi9O+G5x4sz3ZrblETdh
9nsbZumZzdbipKsGHpxKps0DJk2mXaykWLIuVoP+Np70261/cvmETZoUaJiS2k7Z
4nkf8ehRmz0OY9v+A37v9Imz4Rr2QnPv9lIrHNMg6xsDF2NUWM3FEBlCoRP1hA2u
XLwdi67YEoiWcty54uybGbotucHUC6j1ngMmBwPw5n3n8WKRTsQWc6SedR6dpjUW
yDRgojxdaYhr+5uRDIIRmJEydU9QcPie5Tilkb39iyMnPRUq0858uCJuPnuXI5CZ
0GKVQUMVHyDl7kziTn9qWXyTDH4XKa9M3YzUl4HzvpEQVC7UprcqO5Ua3Cct3POu
KtPU9C8vXdDTVTO7bPcayScjn0zBFmLCjSik7salA1NuMecKt/frG9rKMGOAURP2
z71iwqU/7AKwJEeEltd2iclFIBaBwONEWpeeWNFDe32FI4Bcs5Jhpe6Zo7rEOm8k
d9Q/3OWrg2vwTkfPnpLSU82komxyEz94rbkVQ0AArG17uhjQ124JlMv7dl3gTEyj
ghkJ4c/YDy9LI9psgYR0nwf+YpflaL5iYQMB6KyhP8YhVBjrNu0E6qQ0NVHYv3r6
JjQ8onk+j3bf09Uhepx+1rtbGyx/LoRCbfheLckPZQSQitxnHIBgVTDb/CZQLcdc
y1Pqby7rjasU9y1hVWCV6RdO0nyUbx+mf0FAjhn361ZVxOt3LedHRFTEi9QA87er
2GmJ2OVkBBP1L9fiyHJ4OXcHWaxl0ZMc5GWTL5HH/vcp+QScssMDyZNgvtISzGgR
hOxM1gdsq1lY+v4UMr5qET92/377aE7r20O440kOBFkCuJR6aVS9CzSUqqRzVi48
BeX9eP5Tx4l2P6TDqcOD9Q9GchVfRbXzluZ8q6bLHW9v1M3EM8Ti1bu2TZ7EmJOk
yI7CRyHX28qSXltC1zE/1IBK+fLChurFnwIQsgjDH+MYvFsh7lFJ5RBfphx1+q3S
RDnbaotoZo0wU1Z9DuYwWpDFdzgAlgtz7VmhnxRGxhJJ0rt3FFqpZwe5rcjC2h7m
IdWCMbEgLEIlrtIh4/+Emlws50lCe8xSP6XhQtGbMNy3ZGriX9I8OjHdFG2wImaA
NhziHfGZEsX46XBp3bwzT4lPspmDJZ7IQMhSH9FqTvl7nfop133LN779NY4tNgUN
wlf26zOARQKQP1rpd5eGIKGZxbwCvR3XAm7qChSN9FSdG+3qLD/tLfAdT3LdyrOj
fCeZuRlz7fNc1la8KSPxOWsQbZZJb7wr39JUnDd67NIUAj9iQeE8CL6qhslKpZUm
Eq3t791SlUenQKMB2gOSAyynuFgjN9R3fiqDZ1QlSsvhcGeLW332nANVEHBWyiZ7
R7eVx8gPwPY+JMkMVgntD63JnxMd77i3ujwTMiE0h4kc3l6p2LdVc37hKlTaW/8j
yRuS+0XKuR+a3gap700OAqJPfH0cp7IrFdaw5PYyn69Vt1Nrv9Ru9DUQWj9rfEIS
men6LCT1Rsy5LNwNW36i9lRZbNLNZkhYosUUwyguktifBWp2DSJLkJs+V8p/K1ig
5UrztbrqE1WZ82YXVm9mh1wyKRyQmleaeNGDIde0MoVCh+ClIaEQBAXsUxZEtKZj
mk2sKSNjuGU81txYribw/RXJIjLgLNjWSosLtKH0QwvKRAieb63Au2qY8Dktv1i4
R34H98jxNNBuFSaEPFZF+F/KC+UQQ8Gq/PudZmGLa/u3siP/QMrKdpCPFK+6EBaS
qMDEUQwv3eAL5CeslFOst3u09Ee7CZ90OOgnmut1iN2POQ28vz/AURlmAesVEZw2
ObqH4F6Y8l0JOH7qGWvtVIC5H0OsGxk2iR5rddMTXO+6i/sW6jUfI6U7wLh5+317
YCkWM2fbhDHi+ydFSJm36xkmLSQwDXF3naTSCkHdSBnnlVrrWV+YuSTh43gwGzPV
86ey/4L5OJbXqUhsr7hqvjeCBABUC02MOHC1YzdXWoLwmc28wHGHE1sFrvohqwyj
eyUVUmz08kjV5AJTFcrUdNWNsJs0YJcTejWAkcEUzOomvsdNJejyn47QUGZLE51W
5FdJHM2Rr3V/LUJuq/zV0iogsxmq2GCreTDW6lHEdM2yJYxCsLD88vDCajPe0ezj
N46if/tENhZXdER3gOe9xdLYUqUOmwk/FddPEEQchhhytwWhlQ7803ocxSQfLPzp
fjtZvdK/R/yQPXgloASZyp9RJxrYMc4L/RdrVaSBaJYadpza3bE2Y+Yp4IWgegLl
0XGzfWhAZw+Ntxu0+wOckWU8QPj9l/c39XyCoSODdPHfrczpSyZ3WTIJEGszLfRO
0e25CAiVYGx03Q7ZIOPo6gWAMzxuZKsteIFtABU9sMRsf7YYZngSN6n6OaGF6Gzx
vJzbai4gFHxHrBGUjv8ngd6vpArTAw1dpXP+OxxZLGZDISbJcaiGDo3a2MT4F02v
zT0soR1h532nE2OzkCJ5no3n3GA3NgZGnMUMjJ/IbXHTWdvq0Ksv1rkQQhaUcDvD
1+VP2tE9VQ4I+Y56PkMpr19mgN5nzEi3hnugDsHRDP55x/rbZE8r8bExcTVW9wHH
rm7DyU8vvqoUJw9fzw6zeCpspminXRThgvOAiF9JOE5I+nbCerF9x27hiokJsGJs
mScohDz4WUO/QaibtUEpNnTjGp9m1V4pyOvAHSDaR9sCTZczJCpgbb7w4+C0QE8y
Hgbozj11ahk2GuOCtgjTuA5AuNU9I/U9G1FkUnBtW4dMFZP5oSsCAkLOkMeEmNPo
0KwsoLxz+G48FE1KrCAhM7dqzF2jpSqTRjTUex7U2JdsBRz8WDCJ5u0vvIIrvxoP
5R0Tf08BXWovrfmuk/gi1NW+NwRLoJuqy9TEbcimFA7oNoRUzoEt11Z9f1gQJGRy
ZBzFmPaw0x2qjS0oymvCOJtopdAOLOrcVBaUKj6RtsBD5M7Gi1Ar+3i5xkQr517m
bl8XvS796rcHXomXl+KYu+wbScOZ4ABTiP/8da8H3jJoGp8oOcolVK/2gJlaIF6R
rELQGOdCxjRX6zzlRe8Za+ysQfWcuYhhXY1goFnCWyDmCvYvvKnbf51+mPCJ/Bgh
bxjO7p5WTCWopM8Lq1OuTMJVbMbpiUkH5DRn+SM5X2U986nuEIpx67hIaozJfrgm
zZ+iUVGH+y3pe2nJc01+MgO8940f8OGk6x2JRiDKxoHKjIJptx7ZrWa8glO5pM8t
WvGR43EPKQqTAt7YTmIIBi1YodlYLy8l6FmsQlQWY8JzFRAcU6SKJQnvR9aqBUIS
gk/obNJuWqoKnZjJ9TLkieTUDR5Lmy998J8JEdd5uRGzR+41oReMVAMw2TPOJ7na
EG87QdU4PmRelnvxDxwBaQI43jDNjxF/VyropVk6LS2YO+XBFespp/64QUmDmrGX
K2Nq6AyoO9QddDehEg3qnwf6a7KlYGUT4yYVid5zh/FfgnH5eNeynSwpcmyfAriN
De3ufs1oU6bRWSCSki+bSRX5G/hZsrN7QWYW7hWVNmzhKdFB7JwlmgDVgOKt42if
UZcl0DD+ESLuYQjacZzluQvo6g0lsZgMESLmzhz4fQTU/tnzQBEaVX+IBnDiqlyJ
CcdYhqr1pd85m/30FlHNvwG7iFMMU0Z9qh8KpZWJLIQLyKWKkfRH8sXuk4AEfLV6
UFPMiXtLTNkZcNZ+83v5x6wqmeP512CCyFJGdVbyL9Xyyfgoyz+1/d2VXp1iPASu
fHIFbhyXqz7D7hkrzShynlD/yLVEzvwovRDczmiDIfml8qpwEzngHu+s0HWDhXeS
hJGS6+4cHXgLyaYYxVVsSJEfOaiNgu/Rrl4wac82hcifz31r3jHbMQJ6l0j5Wt0/
REKnrm1QU/xlJGJuNxFMBCnsl3DeADsZp7+aJpBaEDqG9C9q0C/uYnrMq+NabDlY
a3IYVC/d31TllLc5MDPumP1KiDF/bv4kpWnC3ErtOdX8GwgVqJT9sfJYieT1UdZC
6ME1Vl4vUaJBt11APgE00Oj4Bvx3aYvISsFWJX0T5cTIrceA4rCvztsihAnABSmJ
zAi5gQMGpuLJ6nVYU5PFPo5USdHEQMnNlpQBQkcc4XiNY8IHezLy7IWDAfE/eW5j
nnqB6pUroBaUOUybJ6zhdIe0uAgAYYQT23t50COO1PU84+xMpCrM+ai62aknsMuC
AjIrHn89yqcCshD0dM9ZIIUC4nd4aL9nryp6corRN/Q4WtSZV8Zzia5QsJ8ECopV
7nTQ3ADzMIq8/VJKU+OdCeONutHyJbXl7fiB1WL930WECif+N2O75htWG4i7M4B1
OclRIvXDTdU3YyYp3XSYAvYwDBNA2KPZ7kS0kVejsb0FWcpsR7fzFUY5azOUYIf+
/2QlF0qh79cKHQkFGSNSHVxyX10u5Mn9dd7JVYUV0Mu0gt9OxxBYGD+O7NsHdJwg
QjXong38Le4TyaUNFBuSAL+fDz1SWH6PQhYn6fArTjdX8/HjeEZbZSUxDg4DQRIF
SHsv+1uGjB2sVzKnkhKZHfuaD1nC1p+pVFfxeF/MWQKipw+0uQxDJ8VvuWY/NPWb
bbaojJyFQ7hTJh/wovZHyqRS2deFpg82xfgsSFQ1kfHx5DXGpsM0ypW2e1A2Fjhu
hVU1kM9ejXLOdw6ia397DIjL0kAMXj1M+TBAspACpSV4gF62V4n+atc/xPayx8YN
qE63ns0HWG9MXwf6nKxHa9v/kezG3rTQfNjT6sGKdUaZafYzfXjQ5PM1UofGE7zG
Lz6kJkfbROU149PkngnmnUuFDyVFT3S2uMQgSR1LhHu0qnRBd5IPz2HXgzLq3Mf0
M6KOG3xABCdqxq7ongYWAz2VbUp4Rc3rl+6Viq0D2658cDkmfFkD7f+MqNZz3EEt
Mmhospfp2T1llragEFtU9Dkx8Sa6yixBOoS+uZPDvZyC3gcwE5GkL9nnAQrBaUvg
zdhEQYQugi/BbjNU7MNMzV+GXgXMrvBQ17cq+ER90P2+0EdPfeDA1vCpZ3qImFJb
7bqLxYdRGGm8JlkzYG6sMcU64cu4CMbY4LD5hEcOxsTWck7iLff2OpczrRrVtfI+
NY+yY4vUtVzZEBswe/izLbxOntzH4mDs2hzJsCZrONNZhebY1Pyi2cAdyWCBxDBy
OVQCVrCLGDvOWpCU2b/EOF8yytt0aPO9Oy27W1zQFo3wCEeC6h2bFJ0CLHVJP1dp
m55xse6EcIs0YCftRM6bLC3XrTa59Dw4o6XuHikTXg+RELpRrZ41d48dBiPRsLAN
0bWTN6hVvHAOVBqbXE7RCF4vFglT6JBRxM+hHApWcm622Vpfq6I2Gkz8pbIJcFu8
7ws7/VsH5v0wckkO0uKlzKzNxia8F5pK5xZeE672q/v+dPcJEeg0ZDfxFav81Keo
QUbVviougieznZIlpjM59lQWU5usKaJez9JCCAV8iekfd1kLs0bpTirUnfGrzaHh
4rSJ5etVCrH4EAn8OVxJlpupzKZX9GB8SgqlSUBEsmWmpxqwL0hTii7LSRIpMX2w
B/sX/iGWrX9HhlN3Xd2+ZyA3SvWl8VvdSS/j4k1XfzwH5jvL3ToCpBysuYKDAynA
16t6ySRHhuDoPMiF4cTQ5orbP9ukjWsTvrssCue8hBGi8BsqqPb+D/TqefLhvQ4h
s6zyj3wWjitkWNgnvF4pzoChuJolVsVBuGjJG+iU5w54mNLRCd1kex8N/vAFI0eS
UFCwNlKDztqpPL/BG8M946PlDxzFaOrlPkbBAHSjumUnuuu/LasmwY55p8ThZ/au
9Nz2PL9JPXCo2WXzwViQiDh3zHty8So11J67pi/VpjxbBPf1rFp6YEIKzGm/EAqG
vX4PL5nn5Qaa+xvHO/FXj0J/YlZzTdGChGtbAJgCBjt4ePMGKMeitkFs7CSciV8W
mDMVtMG80dAuGdAsDEzLqqJxJosXxRPcPDOY2CLaCWw3rim5HzBba7UORdXOJl86
0cXXG3VxbQNU4SJUxzfo8MstJGWKRtB3wLhSKf/Hmtu8j0kHIU+a2FvwviGqzVyg
lUNnhCfk7kaRISqCGuE9nLlGO+sHOBcRqFC/DakAtZ6BCTMwu7qv2kvPeKMdJATC
6qdK9KrT2HdpfaMuVjv73zPLwlNnBWBa+twHSbEYYd3izQ/ISf2OwDDSNzlWLH26
MxJW6TaHyO8e+H5tnWhnWMfCwf9tduOFTUVUweSmqqeh8D8B05S4Ek597xlsI7A6
Hn2FcRVTtYy0ajGRO4JoS8YIkz7Il1VET5C6XcZC0HnroCfvk9hd/n5ojwf3LEIR
gq3ko7Iju4Stiaj26Eh2iJRTCK4MKMOZvAQbH9AzBL6V9C6uyRH91mKiQUyJ5iJK
+CNTSv6d52mAODoh8Et40giEIzEm7n/o3bJdhV9lwUYHbp8FUzizZlVrfMXcj6BE
RickeuswHXITAfC2yQbZcerv4lo7tl5HIs+LwlNK9e9xbVrB3mFZ6PcQ0V/LZFDI
GJvyOE30kI0lAKW0FFFE5PxWxsWyewTeSL9idruaby+HCL+ZUieh6Gt61RiMPIAm
Z/cVWR0xL7JTEJkXTk6UYOzcTpzKWK5NizA0eVEX5WaHVYivics5ft1n7GIlj2U0
MlGwe/CSrMKHbqOxZ60C/FzWRXHboMCZzrcQ8SaZBlcIqrFI7q8bYHXhOdemMk5j
RChHkuuxFoj6x0wi4h54cE4HdwBUUXMcl/xemqhFKqWK9mdnkXCPUT+TbYlY67ep
okV2hQtQkFMcZDXqf05IF4i+Xf2Zu3FqxJZ+RbD858KMit/lGaXzhFcZvhHrhHH8
9k8i2JsY4GQwLXGiDAmmnqOb+7FXnU1Qrn31BBLIgclvnpvxMmlgjoL+6xftIRUR
RPcheIX3h08FXtqbbR470pVaE2OKhUEc3YYUKxzLDZQG9ZEBQtK+PrMV1qI50K4z
hDcTBNjOU8zFQECVTFy9PHr8H+Ey2oDSQU9evwsFMFwzxkymOH9xULuZwPzdfWrR
LkOKAm1FxWSYsAKiFsyrxBUY/h1KA0NDxLrXpX18czZHj2us4TU10uCtrdstcJoM
iykOeKRS1kT4lyQQwAHYCl1Q1eV8fZgBdHXCKmyTo0dISg1lGvntdkDCGLIvAPQs
BJ0wHWTjKDaTxpRBjbrjG+s3OBDF3aFaz6kt90CR22YHSEZujmNikXBeFp/xMA4i
nuZaunQebBu19u/WENWr5Cs2lipLc2bthdSkLCCTd6albiCwz1Sj59fzKH+eRSC8
uq8JKGcVeF7MpSj1uoSG6a+M8rBh8USsSeYg3MkHeiMFfg/YuWCZyxaaSm1K1D5b
OBNu1lRlN+8Lhv+oySWZ4ZHd5WVHMJs/6AM0eB9poqIQuPMKzA902Yd+X7IFUAhg
rte4r9yjWF4hzcV/QGilzdSUcBKLDRppNzMKofMIup3+KNAzyPCxaMJxlHnhgI90
UKz8gyHKu3PQhQhYseIfl6n0P17r1C9E0+jXhAbvqQf+MovvTjeT9S+NRadp83Em
P33WmEf4aoMaHr2HW7dLtGOx3V9UPvyAczOui5NtaNZhhN7IN1Cwn3zjzPPMQNvJ
PqEK+9PBGeCP+ns/TWRm+hHK/8oHFunEXG2xn5C4bhHB2koQyWW4gNqBbEdAMKA+
QTozUX/XQ3/uB1Ci81CR/IHt6YIYwpYiW5hWYc66GvuwkaRSywrRtFFvSEnZWaoJ
7iO4Wa4G3Fz2ntVTuargh2hcmq5JLXH9ELL3dDEemS96qkqmmYeuWwEw3Nl87eZF
dpMPByYwSlP2B8aQoiy4R+QIiodP6i3Ktai+JbdK2Xco9e4vV2BaCqa/D39ZxaZ8
WjhTxs0IOStjAtQR8PXaFlESxcRY+3as4vVf1C70nbPyyO/Ga+h7dqXTkk+Wparo
ExxuhBhzfOXbTvxlIgBQnIqmKI0dUgw2Zn7gd310IwGemHSapRNUPb0DWtAP/tLW
QD+yYUPb3UOTgJBsxNI5mjLgMDphLsofx73krxq52rJ34nh25aYPspoDNCCKaG4D
UHI0rRi3swQwFZoAJg045hyrHUkhPlp1rbug3hRIw+hkJKhBQEfVt67Mp0glT9/C
JsM6gBIs38MhHuAr+i0Espc3gq7hq7HmWA4+Nl3IcYzbDHj2OyIpNMtC8ztd0hyK
tyKwP95vAhMcY8jWqeNdc6y+cZxePnUT4QYMKmWh3CdsGaVhdTKAookMp0Wedk7K
IXCr22YyzVq4w0ydVQ8BIPxfjtnNrfvwvN275v5UMA2iDyx3tnUPfXmA+5NDdJCF
u43ap85g2UTp95yJ9jPO/2lN0xDe2Erhp47/NSWlH4ZRuOU9xJJhK1mITGUCWq81
8sEJ9ub+R1KoErqDwSvGI7nHew9FJiEXxHK4QteV2PL7uzuCYvtSabdKGrovPS2w
GxugkQcLY4oy0e5QL8/ebzcYDvzSzt26qYf0oytMV4tk7q/KWtT6GTJYJm1d5C2u
rptg+YM8jL9YM3gCxxCaeh8LNyJFcSGabus5jrG9PXSPNAGQ7veIK1E/1zoIIe08
xI15BljZI8djyuLxnRfxgHm18MHqN71fzEH+yVSPjku+syALI/o7e3VphxBlhZ4J
ipVxr22q34Z2GL/M6dHsw/bzPs68p8jh6Qw3YnSQ+UXLNgYnZkhmvPQAhn0VNjGF
/IvGbBi9FJZTJJG2evK8Q3Xs0jnCAuPnwYzLols77JGCcK/2B9L74Wb2kIfJnjtY
lolzjk8rszU9bcuB7YxTA6yoCsZroFd0QG0VANmpAo8ffihVnIZK3YSE3S/kvQNM
lieW4OeMnsk2DtojgyuTuFTOLWWi7BMG37MmRAlNTnfBUX/4Y6DxMLxpgTr4+UQ1
HdHjRkJp0S/toSYbJxOVqP1rliChiyL70noQ4o5gzP/yKqyW0ttUfZtPYsX6X3Q/
CgKvWhRKCmnPGm+sgt3qbDz6EnS0iolhjvWdV2DhnH5benhSjFVhDwBIf1TnWXSy
QVHbdQNfzFhgqsh1HfJb0W76/J2PVGlvkI6rAHi0+SlSh5wdAICgKSrMlrE+XdiR
R2cDcPBkBbCqF2M/jz1wD1wLmAcvkCY7WR5OOuXWlz8nYSoB1YKSVIpl0vnhQzmd
VCDsdb7xP0k6H+lKLHMfWOpZ52o4tEW2QE1bco1i3+ItPG5FavA9R+akweJTaeRX
GsbSec4oa3tNrR3MI17Ruobknk8j7hRJ4U6D/c3ZHh+W/Ym0ADGe4rgbfpFaKMy5
0fygDUqItsb+4wNl59N1JA1w/ny+M0j7ty1ZbyWsrv6ViuAMJu5Wyw7XMVrkn/JO
yr4VBbDdnCua1KqwtxDBeFMPUn2uUx+Isppya9feKMli9vuRZnNtRfY2DyhOyniE
d+kqVpMFObJa/oby0BTHNdOohH17s46xE/zs7CxHkyzEOcMX+8cIo75C1tbgGjk/
0mUlDQs2XeIUl7bFKAy77XZT83ACyS40WVasbBcblCMwjvjMvobSnUjflrT3E8QT
HNMv3s6IP5xbHH8vu1iisR6BLFkzf3ueHyNmEykz2siaUC7ky8gX4p1eR/ZInmFV
KV5h1mAEjj6YL+4nipjPdpXriP0ceLJkDkvXPw1YybfQWFWtqcBVSfWSZV9/IxNb
9ESyY6ZfoWjEn701CQNDZZuIilcuh5v9KKz2sKOutZca7rONcycjk3Z3EPxVXBeU
BiIZt11j//5C1cdOd9SvNHvTZIUj+AfVes9OMuP8tSAVBeLSH4kOQPEzV8OFH2FF
N0PG1ujdA6uIQRP1Px4r14cmSWcEYsq+JtX+WIs1tYBo9vHBibz2M4e6aAASKlyi
oAsi2us/U3Y9ay0j7NLLsuRxHAETcBhublsjCLCOwc5kFFUhSShUbCZjSwhgpX9g
wk+J3RWFHoNzPXL/lgYXjBJ9iYChp3q9pf+ZvO/QM6VPJtuLykO9T1bns6BKk7Vx
riCBG7cBzH7TFtJn3bgNHG6C18xijK7nmQ79myspgs+1CHFlR0Psdww/zeDBVyWg
Y+9K3rXc2JoqrP/t+3MeopvJ7ZTZPdGKXIMKn3xYCYBy9Wyjh6T9ZWVIXM8hLlZ0
zDmpQFARgaUDrtRogYmvvWUfIdRWOBju/QW80vK9LTW5uS2lb8q//Sw5OodV+E+z
dMcHbMWooRmwySldlXaFJPlp4fBBPno2PlBIgoUlUGo8fF4MVhaT9jq7gGhEovkE
xGIjp4gBWEDUtgoUWbzncexR1snlBB8hB7ph6A5Wc1vVNA3T04sBRW7fh+XmOra3
EdCVqHQ5Wqcudi1OKEBKSzzW6uX90sjC2xC6K6dz3rc8Pmjm3/0NEG8VvQj5Emco
4qG5h2j6c7S9ufvKcS6ggfr5qODDYNc3BFM0KyrgebHwkMdb6iz4d4MH8pBoDSHD
FfskoYPg51sFN2AZ+K4HXwV2i8DILwKP9xGthup4IwuZ5s6NQFQwWMFSe/uLQLwI
/Xp6/WPjYnFHveGkdtIs1duhrfk50HeemiyzXcIO3W26t3+OS/sQUzQYWFHMIuFs
51GIlfUEjB6DSqZePFabgbng14yDJ4mEoBHceOXr9PQLgq2ahkyfjzOrELSvGLFK
tKfzTtm8Pqkk7BOowd/kSNEbq8KRuH4DdX/yMCTC4U2anW78X6NghSigyJIDCTt8
q07z3EHy6HAfykZY4Yoiuz5dAJAbzJxr7dzkDlf3RxFqDf6gJNJysZiPpW3OCgef
Kaf5DFHPVkMSmZOU+W6r6mIA30iK7/It6lfLW8xFrjxWGkZOqF1iBPHa9WcsjS3S
+Aid0vwkZs0UVkxpm6cMSFLg0f5OMxk8voM7tcqlj+E9lTFEARMUAkI+fcmOAWhL
eyWhlXBeOCePD2n8NGdfcbqQ5c96kEKeBzJ1gp/kot5w5cMdOZFPB7/ozYSaNUj4
pqdSnB6M/FANOFMfEBMU5DbM0e67Ped3CbFcxGQR7ZjH3EeHrJqG9oUQtb+Z5XH1
hFcAZN234Ja971BNezX18EcP+ITr451WkX++TaNO8ZGPpU3DpH4X+qzMMJd6R7U5
VxhqstMKqyKE1+9EBky74ZBukkf0yek0Fv1lwjPfiyR8pDAegB48NAA8J8heUNz2
QzR/8ShHqOIuIfbE5ezijU1Li//Dnx1qIgz9FbJ11gGK4GvEOrujXDa9ZIpDfWTX
SyxjhrGDXRIr+3zPaJAjsGxklCKQWEcRuOwMD71sNyLUheh/q3vwxIiAZUXv5H+l
jFT+a7bqC2dwZ4CF6olmeSjb1IyPEQ7VvcNuZQQAQQFyXZ6oX5jW3s1HOkMitFtm
W/ONz588XNVpabCeZMXP+/loKQ41uHley7gnsOG13l1uGZTT3jMJ33LKXmJa59bb
Bj74PPW5xR0k4T1gr+MR+jzAoKhpFITk6UOpDEIj2rOUGsqUcQ6xn0XCjZhS1YQr
dckBrtVasiX7xShxP96ek7vpIXCUK4BQj03XSWJGLcv/H5X1YyvP/S0Upv13ZyJn
0HrsVUsasuHUiucYVFcm6uXASg7zn5beVCorUTI7ZdGde3gx42OUXepexZB1prcu
ieo5ntmhtAwCju7C/jrAE8sB2MBZPXJTsqBfuCXROJhEwyTfBH4ffJvP8rLC5BGs
8frAOOkhANPyxaUVkpeRzVV5aCHX1rWVUwHdD+bmVKItSAwXCwPJ9RRkxKjQUIz6
n2d/UjZATdhJzwc/oKLn9OLZcdE5HoPrCV4vxIajOQfc1TBgPqzbQXcq1R65Ua8/
gxMm0ah+QtKm5wa+dFnrTGVBsXWozgStZR5mNL/1LyUREI+4iwHYeqqJlH/moqJg
jxl/w+LrWu9l8TWs+npzCVPBYYpCD0uq4NhixTH7m5y4JQZmMorpXBhr4+fBVCVz
rncCKLNSFbWaiDMClcepm8XfOi791PS3nc9a/YnDElWDsH9JGKXD4IClmteGB33m
dCfU38HaK3Up/aO3JwlzjHKcShTpYB9eQS4ADy8TR7n71Mao1uJeuS7COj2gojtN
zET3nMeD7lhuTuBYa6/vtshtm5KPohXoSxecHDEdqQ8Ha03aQuXrCU9btyPfHrFT
3VMmLoKeToODp5I6/BjifK8p++g6Wjk1gwH9XLyNKo9gRMOcfhLacY5YVG7gsaP1
EUhWLxPtSRyN6WWR8Wq7H5VPjVKDV5G/hW4OH1tI8M2RkY8OsdliQRKyl7hoL+I2
Oy1PjNOMpsMg2ETwqyMKXWfzXM8pKdRc6aqboyKWxIBYra5zf8l4KRMlM8vLJiH4
zrn7pb598Gnb1pPOKAcU6v0KojBDDIORUnQf4Y80NAs/4UXAe07Mk8ZU47r8aBni
ATWhgZW1IA6d0ALQsWmHXa2loVRrwKZ/m4w6H3nFk36uUie2AqitAAG0dlngB2pJ
4zuSQ0URo64jP16/nLoh4huwuXB6JuB8l81StYNUgAKgqU2r7XJKKf/WeDBwocuF
4htyszBdKwM+IDEpgizow2Qd3b/nkWkcLkOBL6bjGem5dIvrZNOG1hpCS0Pe/r12
7INOQnPeepsxYZV30kuRHenUNMj4j9OSHdSwE5jg0T8JQSismfRQ79l9gnMBjQ+p
MlBcMbf1I5lvZ+6e4G/txHE3eOhjsS1eqbF/V3SB9HDtp7tcDiwOtty19MfZwGvh
oTCge72NQgyoOHlfE1Bhqu+eHEvHqCkcN4RwLUTFyMXRdZX3dQ//XEKDYbGUaXbn
D+ggw2MQVzXO+qQsT94/bNpG+rtI/CcBBaJ2owJVeQfm3567mTpwHCb4hfXjcNVK
62dPW0AxeGyTx9z1iM4EkdzFVYQcClE0PVxjoMsmHd73cQQXX6yYHFFUphl0Ou/v
vclxz5NwiXdJv+gmxIziS3erVowN4qz8sqyQhxM6MKRKrsjm1D3MPaJ1vi0LQg5c
bU1JthZciWzmupUFZWhrJw==
`protect END_PROTECTED
