`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h3tqw1HR1LpdMpRbh4WESvhk1OixK945k/Rp1pFAwxkzrOlZdxUs+vSZBLnx12BQ
RoL4r1YFRKTO6PAbGZQdQhu/OCh6JrWOTxujMR++D5vd2P/4DqPB+r9KgoWfbmZJ
hux83WL/d2bAyp9MJiszyYXJsQLZmca1DPcyTHAhl3mTJkxODPc4P0iDBjSn2UVO
7PGTw/Ed+QYx/wGybS6QH5srPjffcxt3ENMXSz2cJQ3oPz1kOja19nUrpG4NGReU
QQfUJQD62xDRFoMj4lXDk07N9h+93NZwwrg/lcOrQqeXBzy9sSQLMGng6QZ7vAyM
tNayy5+uD0FBVPR4aIz/ANrnl6n1dY5mpoj0Y3yRYeLC1iLT4GiPQe5kQolMXwlT
iGhNAxofy3qBOqTwR5JYNiCvophzXo82McroHPu4biKylbePRJN4YAtnHfAsBO/r
GqK8/Epf4zFQCdI2qtg6bXR2EgscvYoG+ZRL84hvcZOSPPva8lE4pZmsASa9vDKO
BXtsy1chLANAjDeIxoJ8dL6tlECVl/n7DOI6TcvUl4wjs3a5Qy5moxvYPGTrK2mM
Nc5p3CZzPLPFrFCrBS3xaC2QebT26p7T5aFGw4HMuzWGnTkkhlaw3Uhxsrn5FTcu
inOB4GZM/vyTZ2Pg/MEAqYyEhnw1KM7AFNYsa2NRBBAu2ccfLAyJOnTQidNGJ5Tw
+ilAO6ks1k2QWdwMAkxcn83tpXcy5/xrxDtB+6M84fyv6pJ/JPwF7QbZ3VVi0AiY
8J7+nlof9XrTT0y7dR35gDukLN8G3NxjRzBZeGtUpNzuyxh/0txeLxhh5VIxZgKC
Rmj7lir02+bV7MqbIoQI22c03lymYVVGRVk2JBxjMexZUUvBc0eWc0SrTTV0Bt+z
aJ7pbiQyn+25bUBHId/XsTKTAGmXIc8UEN/8h2tgAtjGUHBNWxag4/Tuir1sNx9P
Su8ZTLumj34BxNiywDPlPqCpX0weIkwa6uvMB9+WXNyRIGb82wHjb9cpuGgoTpW6
Pglx0uFYNAGNhA1LLppQf/jfhGvg6PoYimc1xPguyAK2g1BCn35I0+vwClbZEUn2
P2aBkF4Tjt6NDvnSoLyp0AwtNDlSQ6eHaeCRlRheoidr6gI1orQ89pLcK/zXHzXo
Y8/FMu+v99CqDWdwRUBjSdMaI/RLPkPxdy8QbpE7XFZazbEenNPjlDMhWivUaLcG
3ubIvT+uBZ1qO+rXdosq8BEKWVDt6+bwg2WvZ4G8TGSouJD9Ew+JSo+5XhZU2B9R
/44t6flqthOKG6VAgtLFXCUEC4kwPrl4lbp9/d+e6F75NiOBCHAgSSUU+p9bJev8
RA+WP2AR/bSeLKEOvd6F4RoNIk0DROfcjJwwOQ0p9jh7RdwpMovkLs1moputszzo
0r+zdT0dozdvFfcAFc2F4eMjG8hCUJ4PKFtUoRuA2CMiiN2dG4GY/QTEOZRVmN9F
xHUnprxrFj78lXAc9eSevuXtgpLO5DYax06fw2hhCtzisln7kRSU5Ib6yPN90Wr+
q66uCcab+tVIkaH97V84Oj0agFosqL8YpKge9hvXhKwK3w0RJxutWDVoLjBQSM3H
14eJUHVtXhx/7tHS6WP4ZE2RY5GH116AKYYuqdRWBhEyo50TOhosnLuu4S1ooMUG
+h/oSMBYJ9M8R+0JbAzuf6Y48RsgxH1DcYYGlMKp+HbeO+iPsmJSovblolKP8Ndd
AOJuM9QazlztV/woR3gdY3/u9Fc/UMZdfcBAicL4QAStyLUuXk1O2wPBhjqVmzrJ
QhdVFbIyz01eQ+TPnOyJfjnTLdrJB9IFH6AMItyqTo1Opce80jonmX7hOUbV+B5e
PBoSYjt0yIDpV1DKJOlK1Wzka2FALv81bdiKgdzwmbJmeFstbwDV1Gifl1zVn7Tv
mBk3uc60bUfG8WgBdQQsf9OsqjGSxs5S2u5qZhKoWiUWGbbr3N7l6O2Q7AaJtMti
/+SfRC6KeOn59w+NqrvQwJgSHxrbF/9J4ueB08wICGN7RDCe4hpluK0HsG5pk9ps
cDfo+vs4CeELUzLuofhP3EVf7YbA6wjnMD/0Cd6eWZ+tXSOSprgdXOJn2nGNy3Wk
ul/MW0Ewsm3SyJzXNZUlGV3QaRbkTtwfi7IHjqKheMTw+yCsgHQdGpr6neoZeK6w
cGLy+0UmYZjomL69p6NRfOlNEjgIsJGQSpDLGbJeKkuGTyqTjZXW3kmqEM8dFmuG
vzDI3PdZILCfYpPoaZNyzFaeb+oPvN8C7Z1JWjs9b04uTn0GJst5sXnspBwp+aXT
Jd44/QnxdAKHpDiCe+uc/20ByIZx/3h7lrHSvnTDIFWPeyCGwngqeHO1dRYC0xkj
jf2bO8ekyUlOEAvLBAmH9snZgvwULyYL18I2ng1zTK9Wu4qyNmkp//pswK/oDAog
RxPCND2zYDQ8RWanvDsuSiZ74KWFzTbgZrsLhcqBbJnCF7RwUi6G41/1GAGldbHq
uw8Sz23x+CYYlistAHDhU5rXUmG+VFY0JMe6d7LyyqNdcQOs41ou0KAAZU5x6qfc
pgVqyB63K/ZtTULPvsVsXZHE1pnOudfvOVae28sK2PHMPKK3VlGUu9OXTUxYe8hQ
fnr3EgdW1PVL7ehG6HdQHYRcRP7XnyVZDhYv+5HYmqHCyKj5Wxy4Qisxu0nLMwIq
4CsBkq2mJHLGgMgEh4bHqyfpUjDjhtcxRvGWCuYD7cnfGOVLwBljILEvEZMHV8v2
6VFe8PN5Q7PWeNtGP/KMhv9PKBPfJ5kVi/0m6A5VGOl7p5cILtl1P03egtZc8rsV
6Q6/uyxEQ33+2HJi2Ur9PidBBTpb0EXIGiopwK9IRw49vWtSPb60l6UTvzlNRFcf
ebTNzPGsfjqrQaDzv62/72Mj8wp1eCJ0USh0FDPssraHO4rBUH71jUEhoMkRTjVg
QF0FcA3yVRmXJezbGXTZYKI4Z/bWMgwbxwxu+1hyTdcAXkFJDCcQMZel5edx4M0A
1QbJF5CyEFvOjdMQTVl0jwwHbjhsuXBctqZEq8cvc1ywgfZG9WJYrH5Xw1YtLsZl
IfBFVEVgbjqsZ93sTcvCxL7mjRZe9VgROe4iKPh4QjaA3HRwRUiWj/jKY+uYX7Oy
oPZ5snZlIgWyc+YZfcHgfw6pGbrG09h+4nKKvxghpsl98cHErabgaKrDE4OWxU/t
U8OuwQYe2Melh3F2uBGuaWvNqN8P6IGo54SgbBrYYYGG+kcZw8CG08FNKZXpVZ2t
n6wVPr75jiAioiSCRuSguYJqYt7YYTx5oikZA7MnD9JAFT02/Fc7A3NC3MMnbB0i
VpqzIvfhPnoU3JwhkU8w5M/vFYUI5+1aTFrdHIzENi9TcPPUqBoYW/ouMfg/cew6
aG7DATPbafUV5yCi/pP0rM0h6nrMQ1dVBT+4u9cv6K6AFBqSBvdmNnQ/QZZmefv7
78zpLcwXhozAVDNT9mv9s1/hz+Sk9YyLYPTYoFcXVYcLwAX6yPIupjvK5Sc2B25d
J4i58zJjaz4atg+6BZ0fn8beOb6m+jhhsSUYouosRX1ueExplfuh8HW8nblCqPXp
FJwUNMP59lSqiIvpy8JFUWKfUwkrWTM+ZBKbJdY/Ii7E8jQhB9p5UN4/BeXChROG
/WbjQhzv92bzXLzhhkvUIPyaeHu6llBKNF9Bw9v4sx7sl6fTjwj9C6pz1hXK5agU
dOgn5F62BgQLhmFdwGtvrD1QUkfFPcPNAl9T/GXtbZEwY2w2okwFAatoxMaZPD0Z
m6zFpfXnUxGfhb1DQjotMwxdYygZeaztIkR/4J/8paIo/fjzAwGZHdg/HAUZ3G82
IbPbeGoDEZtAM8FZzzxLKLcGgC6/Vkpg2GdfWwy559WkvCpk5dkX9/HKmxosjCFR
8fLG8YEWeVSTJsDS6W+4/gKLMKT2AWBOPpS+n8k9zv4goRAnZfD7jBkwRPwJs527
xknTb0p9c6UxMEFc3AfT8wrK/ngsDhGH2/5DMApt0rnqwxbU7GiXOF/WBFNRzjOc
VcG5iS5nKhPoQPuQKZLqFw6SqoAsv1uDLyWyW1TidPR3HV2nRqSzw3M8K3lZ/2eU
aYzoEk3WxeZRIkkp+M++49K/X+ev71ML4oxJ0QJHit415gaocWzd3jjNOFEpEWXD
ONWCzgtNhyQNvm+w8k4ndPkvOflGBR4QGPGv4rUNAV5WJj7Fnhx1CcMzpvXPuUxo
DJ4ikY4z1B1vj95nrOtRk9HuVjXMteygB48VbM0hlf+p/SIS4+ukFa84uCFxTzy5
fs5QYBK5e0e2Sk5BdLcV/xTE3lIl0bL6/RGf6KHxTjkil2Golu/tK7TxRZhwOSPx
j2AGaa8TOGav0dBw45fmlkeA4e9kwi9CXM6z6V0YUozZkz90fvCVyApC3lkOYUOd
gik/2sKT5sjpgisrr926e1vGDLUi3EAPTCb58SRctu23qRkUKF8G1KbmQJHSSNS3
2dAqyTO1puaTks3TRXzv/WJkCjYiZn9nqX6gNOM0+lG0kKNLfiUddPaHDtI3RTMA
DRUOs6hZl3aRhvZbDRiUo4Cgmu9Ys9AaHGdSG1MCfLfJA6+hjB1K3AinWKviChey
B66P4ZKv5DQTcEKnXCmNtlUqP9SuZcKwbZ5ZXcOwW1DdzGqWtBdhIZSgtS12sO/h
6hj1BubR5qduV9N84FX1mIEpWaN43ZvU/btuplNVePWkeIdHDVOlbdCviZ5EkMGM
15wNY6J+Yq8mYA1SdJDMriMUtQzn1yBWs9IPVjxvekKvFQusc1yYlZaon0CjigAF
Bif5kKXrzi1cz6kr9v8YKg1VprU4MHG7iRu7Qn7xCki6Jlh7hybjdTaWFeFYqK7I
vFw17EjOh4BlZByPmTr9FECvpR5HDPP2R2JoVBe4W/ZhHxESwsrK+HlNUYk+Jdqh
TNBxihuXq/PvaKlYYYiYb8eBFNbJIciESPx9gHJFvQNX1ri5XW9tysBhcYS1KOwC
46u4N/dYvXgx7DDKX+MXfV385kpkoBnHfDGiyPePa1nt4XoKzPIrNOIPaaemlIC8
wVcHfqlClq8bloq2OF2+PNa/qkS4vckVrDaDJDLgyPCiUkfQcY9heSx0xBXTFyn6
tqxKpiIgiiM2mQppsduDygdCeuki8FMbxj4PwQGtPjCHAzEqFJ3FiwQWYEmpZC3J
l4PWuJX1lBalDH/wNJ3GLgohoGHT23O7yi3UaW1VnEggquxm85Bd52FfjIQcwjzT
eiojbbGrfTbnt2QFPu0kOydH6tKqyZGvonBbbKZJVWHEbns4Cb/FPOeIQ3DE50Jx
RBlWwa3VguYfA7USHns2RsE5Mfvrfl6Qp7RaAow3VK8NWfXNYyEPACDoWs2nK9HH
ZCD+5RC3ihY3mgQwHSYhcqEHHfr0VXBu7hqT3/l0FowDhqdjPbwXeN7zxdjqigyl
ALaNssd4Y+LxWfp9lHgFYG8vLCqZMU8HUNCoz3pYNOffprO90nna9660r+puJsxI
t0nmcrYUScpsrsXV0zVoWtE8HlGr7Awg36zP8HDWO3J1z3GtgBE1y9v2VgGOBCcb
3MuBOssFd3DEHRNBVCIHCsAjilUXRcP6BVfI9VRnMhUiV6Lr3BZOt0h0M766USq2
LBiupn4QDpiyvVUF4seajJokTUBhGhK0/50rI0wCFbGvS0bdrszMpituzJxsUKXZ
aW2Ot7ETQmorNMwbJjISH4TjAm+te7o7AAR+vPHa0HkXoBpRml3mLt77VQsfZ9uZ
1McNmoEHrbfEbYWInpzqvoHo3vQQQNymY4sc/FZU4plP5uMlO+5qxTa+t7YJCDpJ
+IskYLRDcmNrO6pIZgu36kUx7v51ydJkPTG4ms1/h7M0jKhXzaPHN/pPK34v7HT3
LVXGl67FDDnXzpibGD5hB3UWPMw9NhfpMDdLxMWzlifp1vaHNOCDItOX4r6WbdIP
QMlV8190IZNlgaYd2qZsIPgKvuij9JvZzcIXW2OwQEQEk8Lj7FbOfu+1Xe0M/UyQ
eBFuu3vTuKM4N35ce0bfkd/rbC7xeKaLZZb5sxt/BWZse/RzRGmVD8tQ/D9IsqJr
5cHNPVJ32VX7RP5GOtGN7004ICKYP7UxZZ9HY1gJajk5nloUEW8/gMomeDCUVElB
MONdO0k9P8lRAZhrTvAmtn1zyemKEhA7whnhaaTrh+aCj6dAY7Jut9etlY6kY1WB
579za68UZ1sSg0o/RL2KmwIXubqK756jSSFnlECA72syAnFfaM9ulgOpaZuW1yIY
+oDxgsT1nRWZNa42HB2yMe2dQTCgvKx+PYs7MHNUnJbu2xmDb/28yokkGzLz1+Z0
WnXhldr/pl81hXaDzeC4UnFAjQZTPNEX+MczTfc9IJxKAa5xHu0d4BStgUVwjjXI
M9BoxOjb8Gf5R328I465Bm1eKSitUU4PAgb4mBPibXpcSmpAXXv3UFAwf3D1HwwL
/opCupbC07J6/Pmc+L/Wg1NwOhAZtKlLl3MVaTVxCudPmZ6+mDlJoU5lrC5WTvV+
79iP+yAGLejUNW0Kl7tK0v9C8d+w0jvL1r6EvDFPvBHNYRPlO+UqLB3jd8PglGb/
2iAG2Q+765dvtw2EQHJhOXS7XA9XgAVObPgpWyIOQZQR1h8E30B0KeoRZDpThAyB
6c1sMjPuqSc5mpqOxojljD01NR8Q7Q/Vn914bRk1RqOVWuh2q3m3Hkq2isHnNR5Y
XHnPW/j9e08Rwbw7oRcc02Ip6cYrDzPCHY/UVV1pkLvtbZXxT/43qz2LRxDt6NF2
6JpwGw+V+6MznrH9nGo5umlGOWEys/CcsrxG0Mpxt+0wsUy+1XoiqymH1IUIfY3K
e+zfBPUpbFu59I00yaHNn9iQHOJqyQcURvd11yYoN+tPu4bgLCyp+eBCazg1vGug
YZcVFzo7rrjf7bYoMo/xpEdPc+hG4/BdSKGu7KB48S5sbstXRli3eI5n+cwbIItk
Y0kj4b9ICZ4beihF36VSotEHdVxdSgDcPNA9ZNvBBjeU33AhDrX/1WVXuQeCBEOU
2VgaaN9LehjNa7JZRAkLbX40fDFl/oxe0v2vOb3Cv5lHyLYok5bCa+1lQV580e4V
R7ZrmoF2ey5i/Y+vjl/s7qjlWtyv0+tRfe78oZ3023wadUUm5DUZ8OYAwL68OiEK
sLz8/6DbeR5uNE5rFxXa9BbyXFgQSYAQbn/53Nj533rmED+FuDN1MYw1NKP/dQnI
egC2oTOlcoFnSzlNZDN3z2K0ibMIIK9bca4Q6njmSlw1iU86wdEN0swgL1yT0lxv
3wPZf7EFKozWDAzM9dTETNAk83OMCQCL4OqG+y5lOCK+avYvrve7hUG3gHFDTy6E
zZWnNFYY4pUdtv/DuBvxoZkmfHKm33ds/MkGGBvaOftPZxyDvADvzWioRYPS0fBh
UNXYCAGIfi3Hm3MbDKq5GVjqEWz0/r7L97VVqRRROAi7pqe65i7420sjIy4NaYQ+
3L4A3ZCYi57lqDkR3dLPMqendw6P8hSFiJ4PSFbuxnmXI2XX5ltdO0XUXE3c0zzS
RnZoPfp52rAtFnAFsqiYCSS66V6kR6WxW4cWhS7daa4hohL7LRRdn3vcGoMSGctl
Bn6oG7jSKOhcIS1lKABr35yfpZqWrnzAgLpuQRVrCFxY3fhiRmfO+qwyqjRw7HWq
ZEW94+fYXENZi+VTApyb/cptvNLn6ANzYxAjlScVmXvhlwXkoOMqbRiUnDQgfmbF
Pg/mInHe4+M6nv+liRX/MGRw7Cd/kzmx47iGSXVnzWUgSETg1w/ZeZRVUaet2LVY
MkKERNbIQ+uo6ecCnRPj68SfwIcesqbbmn0ndl14kSykQNLlHugQ0UpJV9/WtM1d
yuzFQUqPmb+X10SjPBzcJSdYfhwttUmEY6sgvi2SHE4GhT1kuvfnW/c9PhOWFSwC
7PdGZgzx9M/kFnow7eVabz9AX0Ih+0cTxm9fmoJHYPeh+tfYSY7S7d8cQneY1VbM
oE5YcrA7Xsnl1fTzBPAh8NPCllUuY1NkMMwQVNmOOeJfJPu8x/KkITBNCnBbqeC3
3cljNNos+aG+1O/+lfhByLPvLsF9gAfxEUbGXSr0iphPH93/O3IQ50nPQROVHqma
WSvP45Id0TbS/zUa9zKtyf6H10KzB5lNZkDoXFE7yovwUs6RAu7s/pFIsi2bJdSx
CzDuDKMMdcM7WLiJMI8EZQlH6EGTOTQDY7uDhuTACnIU/Vd6U4ZOtmrqe/CUbB2L
FLCAx+fT+6wAX/CrxDr6bPsRl9TuXyYzQOc5QVqYZdGQvZhX4rXGQv4o98AeOg7a
tAXW1irImR6ARzQKoAoJVtRAhftPfcRTEgyrggSitNlK5v9Qo5fGr1SiRJSwH3h0
yW5oORVR6EnJH+4YlX55rEJ2H5ffVH/xAS+kOLe+cos72Bp7dDttE0ctVgRl24bF
H2ZHex088HkWhYgWG/cPkovQZvVkGETe5gSGqbcRjW9KjQzcPezDL2U6KB4cSzUm
qLCWx/KRKQuPyzvwws0iUvhBNaltxFzFSubcUG4wLI1t+vA55zusK+uOO5L7nUho
c2M3BF5KFRoQPABIaUiAy24D84MI/V33gQIYqw/z/G9floDhLyB1uENsjiTjIweM
m7s/eX2Uz2CuzvxOi7EFL/kd4EjuAND2CyEbx9ciB+5MG9NqcpP3G+kzn5TLez8I
q+PlCfPoNzJIRVqr65Oh75L37ZFGZ60G4lmFOWO9D3IFYKuEITQM7eLk6RQHfquH
Adi7T5iZ0ehqU4Wl2egHVy7KwinvNQoMMPbYSmr/ESiq3I6KvFKkNE4mMu1rQ/O6
krOyibdTDTi3ouUMkT/bx1fx35PM6QzZ5cJIAmc+EDc7sh92rpP0GRkU1i9e+yQ2
tvebwcGuSFHC1XwIiuOFMbiVgzaD/d+z5ujcmNAV2TqX5NLcIdUqDYOHPAWlx1qz
K7Jx2D2SnrsSuVlgvkU3kSS0lu0lpK+xjy4VQInF56NH3ieKJvo3IA5SAU3VE8Y/
rlDoV6tmuxj/qMziALsZIV3prcgu+LmNjMVYTKlYrz3JtmqmcbTcDzysO3mN7AMm
BAkqXhRqrspRoQp1S3B9eoRXmR4LvzF9P0UeCDyMnem4k7KRRVkFcDprBR/mJl1Z
yljEuf4N68OhhcdrYepVazRq51emoo0atbobbHcc33ygjQRDMfIXH/GJc+4h2Ci6
tCrr4El6m0Nkx+WTAe40B/QYYQJBxwu+aippj38neAoDWdnng9icU+IxvSr6xAeJ
PiGPJnzIKTUsgNPNss7FnpFxJXr3kVmcDTT7ayGO2+9UWC235Gb1lU8rCSluEzDO
RYQgP121OMTQt4txX/ns8sRc81CCiEBDxJg1q4z5c74zx4Bv12S8+rQSHX/N2zTN
HWQxyqbpQ25ZwbTTgUsOaLllkyp62Ue+K50TUb6hyP+KnO0qFH//wbs7EbuKianj
tyWBZDKFZ/5aNewNsaeoCzsZ3CgeLxXuFIvhx2yWe9SKneXuVYaKRX6GwlZFv238
Bdzg5xEDfXC3rUD0mpx5umDeW2FZFHw7iraaQXQhFkGHqttpYtMTDY7zaVPPojE2
lUbY6b4v4ahnegj1p0e7d38AvCe2mzPI0mctQOkcX+pK5y5N11npQFpr65FcqodF
BQc/x1wdzVRVnN5Dte6flA/yH+Qb3HZIo2P2B8SC2b/r+LVgsJ4s0uK1YMhALgbh
9TbhZe788JFo3KbQPaYM2IY157EyOldEsxTam7wU8g6zVAUyTN3rhNJey77utxmT
Jg2duBn1f5gdxrxdnXndQMgKKKfgARf/zBBtpRTuom418KILh2YoxJSvzsqE8fig
PueXanxgpxTgR0JstzD9rNbTjVXoiZK26bxbIi9bbUJeWT73oIJWZ7y1okk0coHz
JWS2eFEaYMTNSJOcSj0KZerAaf1CpHf68csLQITpToxFqvAiV5FVSxvbGRPz/nhZ
kMIpJneCd4HTII88jPlT2QtkXqOQHKsh9iaPTwNv8xTiNMFTEFNel7E5/a+9x/RL
et2HWUUV+GRjZF/+Pq0mQvBQ8pjG++ZOpqwYx02A4byVvJRgTdUOeGDom0G6dPPk
fMHemI89tjC5+RqfgriVlW3AF0CYcPLypEmd9AwhqEUA51zfTCA2UVWZm6faitr6
2P2m0opdwS4VRBBWowsDphlkxyWxDGKLLM8Ywm/fyf24OC1xo0wfAenwmmsIMjoj
0Um/SWcRb8KR+ylyeOYeXc5LURYJzdDL1De152czIKmEXYN9fLkNHFBn6gnNlBrO
4TAsBrJuShf8r5yIuXbGIp5mN2/Tgnz+yhGv+jfJBpbNTE6G2IL2L6ivL/T3EydG
fcNozqTPkXtbtXCbrZRmFQnbsB7pDBHHkd5uaEJaVc0MNrJ9k8aam3WaiIwtTGaV
GyUBCKhvk5g3WPGXFni4ZW4agwrFjrxXp4zmOzvbPo7aYt2sMq7mcNYxc0TWc2mj
SLpjukrJOF5pZ0Pmg6Eq8bq7WadTyZ9wpRACGswD35XXPXivFDziIkSZcPQ7S4vE
9PKZEOkw3YOJWONalsw/S4a0j8+jm51f3TjQcMPdrWWl0/szQwuvmpCw5SAA795R
CGkJpVk470Nmbo6vEVt6urO5s4fG5f+muQE6q3mWw7nbhdjzcunjhQRm05HKrDiJ
QfvvoFFczuZePAiG+iJCe6CmkIxi/MA2/FJ6wT4yySmI9lNQpeydBeWpZxRDt1cP
aGo5sLP3iv765WduLKVTOBGsK7wO3uXA2xbe99uWLDWfjjeh2AcxpcrgAb6B0sXA
lY0puli+xRjgjDS1gQ5vwgkOwOwFvGzw/+g0HJVJd7cc1nrP8E1bkxqYyQHu5I7x
PVfi2668i04k2j4mqwTMAVq2V3EdlANxsEqvMPrI2Q5wfCxccyQ0dRVnAfsR3qTn
2MUJDSfPvf/MRdBknasXv+P5M4QDAWdFwqqaiLucBmPpMuP8Q3su2TID3RI/14dd
NZv3IQ2lrB2dLPcWRtcr4HCd+2K2O/lJKqAH0mGPJbJy30s8KQySRXVFXWvWaa+t
Pft3Rox3fZGCn7Yym4qTvSxt7XETSFFqpFJqvyX+3tbaQGb3gaB8JwnlgVK756sb
o0i/a0PL6j4IQNx2ksUezvHe+576pG6M5ShwwXD/JuZrXiDtMRBF26x05Yrk0yAV
ab3igAxJtldCYhqv7Iddfo0fuzr0QQjppvrTedfg6iX+FnNSwSW5uHJtOQXYJVbz
tlSR7dLKnro+pNgPRRLecYs+s+qvDnpckGxy4ewYs5qocBKk2ORqZngoG1Ncz7gj
nXbPQJagLWFtvKFA4eCLGzdigmykwW1pURmq7UzqOhi8un+WRm/7Fhn60ulTniKu
HgvYyJbdTWGqYZ22dJXfCmm1nnLledr+Qp0VP6I3fgdiCQnv6iSmk0VmBnSXRojI
oacgS5FyD4PQNk33f0x0wQkxKS/a8D6cgBkJ/YiC/VcA9qrBneSWwudkM0oiEs3B
H9E1gG4k7zl32rgAY2RG3R148p1g0/IgmNksn9WWvpzpJo7FXBSTG/e2xbJPicp6
l6u9m3P76MKH0XwPVyMMh7xV0xNEnx4jwfozquX3shpyzMtusd8vwaXbIIlIdzWW
JCO5+jFC+ty5yUfxyScfF9ozrfihtsyCQcO9ptWSe13+NTRcZJp/PnmyTYEcfnSd
LKsgLRimt3ahwff5MGIEN9CW7fgDAzL0a8GaMKzyviN3Jwsau+xOZ/MbLf5fV11m
amlxNuhyjcY4X/2oFO2AcNlGo88h/a9nQXn/JBezDN6XAIgUeHDQcD3T3LdJx3R8
aJNUH2EHKG6RDZ9bsf0ML/fz+0Au1+NssFHv/nXyqlHrWMm+3IkTWqk4YHXhQFQ1
zRU/jzrjewiHp/ZVRP4QpgwcQFJ5sQF/ESzpww7+jv8dWew4MJk/Ulct9onfgrc6
LmbUq1tgt8ctBVZj7VFDa5hTYtb9ehF1gJG5pKx9mIGY1ua1I/+iH+PDddk2dCcu
YCevkSQzupwcsAdkUeSEncxuwZaiuTQkywWPP18WscvlURcbW9uQ6Mr1H+yaI0ec
bI6rj4dxmgynSgFZNya3d2mos48gwpk76BGxK9AaUWQKm0D9ESm9rfFz3ocbeUZ5
D1OttWLYCgTqYjlwCxqWe2u0/zYKhLzEnmg6uVyo/yY3SW+D1DzyncTK3BCiPCD/
CD++and7oVppZc7p9K5I7IyagmOOs5M5BTF4gNY8tH2jgrnJm1su52Pn3wEVUcvf
lLzk5eJmsV/3ILwA6pKcoANyopXybUS8I+kIXoHlSvTkKVArZ4gfplLPCOhL9MsR
/Xwh/O9t4Ojf6iLr7VbGDfoK9GYJSbY26NUe7GwNBQ5eep8PKr6FsCAAGvt6GZjn
2H5rkp+Y2879Q2wezejW9M6l4MPEyvaOI8yauiXYbt04bulvCeAN93P05UEP9mW4
bN3GYu9j1YZpKJnT0Fh7VgMRKQQPT2R/GlXBDgZ1I96vaRdprFq/MVMdLxRzeL9f
K/BvugXsVeqBb0caermWj+phXKGO1Mh/sEgWPjsqHAdFQER8U0+a1J/Qe9g+aofp
nNr6Y9Ez5WjXah0q11mU0j7Fh0px6yNRMybIK77hkMOH51sCWl2W0GJ5Qohpx8TF
DtNiX9OdIJC/WLvQ8w2UG7nRDpQ2kWaXtYdtK6zPbJnKyUJxSX4xtJiAeej0Te+Z
z8D9xeUhMppPKNGWd67aDFOfHMVRoB3gWpwZ3pB9G1/J5vU5bkzAXV29xLE//EZ/
04L+eLVEpMvS2Gq3JwdVJV0QawJ1Di5HhfDY1FFvSXGxQ0xXdoNfXO0SR7fBnUcZ
ps6vF6vfVAAFXnLoabz2xAqa+73p1xkxgIJ7zdXBH68gQg8F40GAbxwjnsx8F5a0
oRmgDFXF1HqJHvYbSlHjIPorJ6bDIMcDRhpIVkLnjr9FIFByxJBg9mdkca3SJCmm
CyGel0yGTRETaO/KdnPtkV8pgt0/gBIllglIQ5hnWdK9oq3w27vg0RwqYPrA3LEr
l5Px+rtA2/utXb0OFVMc8u3hcRpROioe8T6MVlAWuOKYkmdipNGKD/cyhMwdf9l5
mrsYq7yhlqGRyHrR5CG+rTdGTs3BdNQEo7k+G4L1klYUuTWpaIzQZ0laUUZU9Zqe
fbFKpJIk5EkziiyJWz3BukgXO78n0qGtLn4qsYO7aYEufkvSAhmFBzX9vhECNeRU
mEJmri3EVAZWiMoOM0wvcQfY2Bo67tZbabkdaRJLEpteUNhGL+p0C00K+SSMrvnu
Uu8/XrIbHl+7ZxFuuuOjSZ7C0vVyXdMfGrLBKZT0rHX+Ykadrz0jzBpJrdVaCPLo
1/eYTsla4HDZExJ4XzhKI0ySRM/8fR3UeXrLuk0ca1WhbYRwD1XqzRRut5jx2dYU
XUhnP0TGKyHOkuyeoJrT10ZYUeiQ/Jh/YBxn7nPmoHS4I/t0UjeacrSqM1MIMynz
HIpExcYAC70oKGPIjqd32+2Zoe8tPTr1oSc0PYT0sSD+m+sE5UqNCSGGidF7InCo
n9tbD71k+fV1NwqSiUazAPWdHbfj3Wvx7otNL0vFX3CSlNjDdeI2yZS19kYe3onq
veG1xty6BhrsT37cGLC/umgBIyS8lXEIYZBkDVmth0YomTqlHz/53/pZCduQtQcT
Yp17V2XHdSfYNZR17hNK2c0UA15wYpjTSutktLKfPn7ah7/KDitZrhen1MT90qdW
drS4e7Ehygvn1tuqTf8JcI6u1rQXRqQIWj4WhROvSJajF/mJXVD1wQct41jqEThl
rqYNK0eSe6KHq9THdmdR+xoOwegRyiAHhSe52Q5KoN7UvV6vxMCUqecm4Uulxztd
a5iGuNGy20uOUJlIkSczsno8XDJ94Gs4TdNYbklbvHNWrWJl9ZGbODq5y+/OvGho
IRxBmhv/Y+T7UpMuBjEIf2r/07J3rVeeBd9QFUXPM3POYtMuEnkyZHXRCwXXXf/l
gwvrMErMijmv5SsTuEtVPRUigtADNYcmIJJbrnrHwF7RitmYRFGJA9WpDt/BzaZT
0GOhjSt9kcdaEob1zTBP4AIz/0a6QimrnzGHtUa+feedN9DCscBkndAbEgzytPob
12Kr/BkP1xSPifpLKB6LpmVlPpu6i8/WuF8VDvbCv81f+Se0SkH6ux2JjTMUc9T2
apMzi6fGC8NoOAUePoWiNrHiutnsLo6RvlLNf6/Jqq1VqC/eXSDS4yuydYduKE1z
ejMQtxA28smVV0rGK4mY+DabFX03sYOB8Q7yeP1w31NzsQzTCc5gXjFU2q6Oth2B
eiNbJkn7vin41IDl2Kn5z28D2juvYnIBs/Zf6yw40c4FEHnsVMefLAqYMaabsarD
pf7p2O4+pwYXQyOQxolXagYYIzlYFNG8kuTFv13huSVoEcqA6C0xhcVI9ybeXL9x
y+n9kQITv/9pLiM0v5Yh8vwjk78ZWBNLJX/ENETOoM3y29PEHaQDJmhviGMgJIEq
CFJ2g5wrP3UvMbWr6TMAznt270T2eQrSm/KISGnA6+BrW/0bjgADA+okUnrMRSMP
Es2US3WkossmkCidgtt69qBqGN0+eNmbSsKVjKkrS+8QR38Rrbn9lxzbyPiQlRDG
hzs+BC+vnJTlt9CywbTjCPFOLf0loAmyKfVvHWhTGIEPmD2K7ksMeAwhtuLnZ4jk
BMIo4LBNjoX0gNA6grIXqdSNr3o26sprjWvPwOo9FPa/ALcq2WJy6/zM7u+U5EvV
aViH2kKP9BJusoeCAPx/vDMb5QISXFqZ8JmbKfXAtHwhzA3H79NLIuD6Vuz8y4pk
K8+5MirGJVlxzKbDu/5AV1wvksooX/vF5E5tmgl7yHNqdUVUcFjZBXo4VtktmESe
DrEm+Bl3ZrREBOvLvoM2hZljPeF1oJq4lJ2/g/+YVqCtQYRxuVBAWKpjcPE7bd8/
/6rjE7THA1v6X7S+uGdnjEa2XJQZEd+3R1Rfa2SCGFWIBGgh+n2DDhB8bUTIP5wY
RUdweaf+0VYfSfcxOSA3ampyxl299NUJl3OwhexFJ5R/Fqyx3rIZbN98jXtFQRU0
kIHMcuIq9yFzUaHNTS4g/q6BiVuEZOrdU9ykNh5DA5hLAGolQyF7/GeXTWIyQWBt
F+AiQxLN9jCnYJFun1WGLqR/c4RoAPCDB65E1jZP7Yzk9s8vPY4wARLkgOYj/J4V
pFclEdimJMTtcJkhWHXD9NR3IIbxs532Jvrc+decpPGAXFgk2ZjVl3NKL1vERbDQ
H3/RpPTPXnK3IYcZOwf/CWToeZ5WP9P9grPnJWNaHoAdBep2QivB/GqkWSHrYhyF
c/nB434yVzdAG0/MIt+uAoPNs3DsuV7Udinc7B+bB7C4tnKwg3sfikNMtCc4Eqm5
vK5D6C2TRrKvKRYYmLSI1beN+ApzSI167Fwrkha1dqE6IiuFhhUStjhnM8WZ8f+0
ljbvc/1H2NJitkzGRcSERdpc6UEORx7xyfFYxT/G9HLhU5KA0rxVPyiULEIPA55k
4nlp2c43VQAFVjjSB4KMpvL8cmPMe+qZ0E+waGIjaWCHChswDNCM2iE6huVPG3K/
1DSVu+ooZJRBemH9eppUM6teNovj4IGAhkFa/a/w/TQp6d9PcRWQTpYh5lP2arE7
RHC/loKKzNu+WgEJTSGY0oFU7A+VucssvXOFoHXljNjEoEojNsUC8h7tHaR3Fkim
2s1SUQq2yU+WuAXIPZ7Lfuu5aFwZOfzkwWshtpktLfNO9NILtfBZh6H7nxVrGxJx
vgtmojFr79DKlPhD1igfzpfMIotBaeTgdkm7kysw70plmjRJ1hNGOzIQGdZoJ+Df
6vr7KFP9UImtHHnt3H4GqLyBgJM0fDEM+OBhvTyjA+uvU1U+lQCA4KAF2ncLGgff
tnbu8HJivBbzlG/h7wFPPIV2FLQIBfYZnhzhqioURSnN9LIsBsk5+eRgg44yj9vn
yAMYyh6+rQNJlCL8QnvuI9o80gR50I4VHxWI7faAN/18TZvzlGjMB9yRWFfeF4p+
NAHsgSaAf1pYPS+EEKI7fSEWaK2B31R5i094Hj8Ou8OsyKUV1yWoxxSp4pRdBABd
TLHeXPYzasszGM8tQAab8CYnVmMl7zlJPggGIufN1xAkes8qXhTcNbg25nelavhA
94enHCUqow2ZJ5eeryMprqagIDjqA89Z359/EYOzOaHsHEajYPNyARdAn8Zp45Fu
kYcvcQRkXZhPwUXGkocQ1j/TWhCVmv1uPth/VfZMnTm8iYPSoOlCEHzp1KvFzpoo
kk4SqNFhBlstPGJHk1KDDapaXc72K8IbgHAgbTiwhlqfP5EkNGDSZo4+9RBvHhVW
AAP7FqzP6M9sEgEDiu1GsaMC0w75e/BjUSg/K70AZOe/BqB9njhh6E1jAkE1hnIJ
d69lB6aCa6She+0oQX6EIB5YyJMIfoPo/5ARqNxzt8kbINEDNDm8eg+QoV04Mg2Z
9wZiaxVorlueYAOs7Ab26ITE3LQHUQ2SiapMMAqNgea3ACQ5uUvrmtMrz54SuVQu
9fnV0i5WWVBTEe1U7T5m+QtqFcrblRWUhDOiAa5vq3gobGofqPYhM+dg00lHTy0w
VMMWq2igxukB9nHp4vghfgjjnFmZHGSJdEYedkSOipD0+B+YMiFIzLazuylnxRCH
MTKrQ7H3kkaZH5pB0LqiRMwjSgPUhH2TsLLgTF+oMFU6UOAtdMMVsoRN8rAaB19M
C+ExUlnpPac1Mt5pxsynEyH1g3mgO/kpCw5TSqwdBqs19gSBV1zNmdNXhkxdFq4S
LS7PDg6nY9kqF779gMyzW0YXxVrb5VheDsR9pAuId6GgZdimcLujva4BFPld/Unu
2AL6WCUo6N+lGDHx7XXAn52Jeeu6h82ouMUGS1mQj6SrIHGsvQqEQfBo9zRSGTYH
yUa8DhFkTGJsB2KwajJQ/jtZmGj3EnEf4t76q+9hBahB6mA1z8Iz0LIYsEjL2ij7
ODh9NvXAN10asJiQiWLE1Wvm8xSqsJQDhtQo1X3qNKZvZRfvPhoXfjTGkdYAroI+
l4M9rOF8FsidtItpK5Jhp36jH4zFGv+jLjL+nYk6L4rdhl/cB5375QEgQtAyVWf7
+oSYpZ9Sy518BPaNGrCaDZ2Ls2Cs2uT/EOfVgmyBOJBtunsz7P2yRY15T6enyIpF
x9vqDySuxXK13eOafHzFhJ+xtELJ+mpUL5lcV7LIYm7epsSPsa3k3hpVB0qeE75y
I3egbitz5v1Y426bfP6Je1j9khqc8ybh2Niu4jBG0r6k6GkfXws1Yz5OM68IT0P0
jLk/fzdjgxvHTRxcd9tTnM4db6Kh1mcg7sN3wXRIWfXp2eWSWulgeSRgCUntGCjm
b0TTriTyTE75Ph5RAf2jHYttv+oiIO7wfk1mwD+bEQ4g9ldXwJ0fHZ6pZl4pglcr
c7UShU0CwZXKkVjgEXe9Cn+0UPFaDksjuuwP/zBV6zgvbNEs2yTB+yiG9Gsl0yiZ
Vb+zXgMadF1RLvojDMqHXnK63ITO2k48EktmQj2BiPCZ7/j0loAGdYLNtvHGzDd6
4ZZeuSPa9IWpR78UtA9l5YRNHTdJpx6hNxhQn3lzpWnZ875i8m1xZtv+Qka/bSd0
sAZ0tNL7l6TNt9Av1uJe5lGLR69bUKM5hbgCBlRxxoXfTsYv5wb1xXWGQRKSPg7l
DIWSjYOVUKSBZmShhhgpZY+ryRZ/KINzKaHtMOxuy1BpGfI6bH4Y4W9isbzrISqH
140epeV7/rhmN9Mea6CRvBgSO8dXqOXguO7zEMnf9UCOwzHZTEz7c7ggRgUFyndY
X/+Qihxaj+onL/+An7Q1wxs80LtnHkS+JGOyHjYQkGpfCcrInCtnRsIFIDZflucN
VDBvp9YRhHYa3OS/PagVJae+1dbwx4EHBpj86TpeCnRcwHI9l0iif3XlQKwBAV8Q
AVdOXA+9XTNARba9YooiHyrqp7fcTRDVetMMjElCcDwSidM8tqWFEgADPZ5oJZvI
HHx0RstEXUA5ie/AGjsYNz6GmC5Ytb40ilsZ5X0Ivz/pAyFzHH4ZnGHVOq0q4Juj
bfReOTjL3pQtptxD9RyiZN/YcHZyHzxZF0KGZAyXU0FtSxYIivmGEz7FEwtVviop
zTKGX0nOy9umVJE8fAAgw9EFmQwcAI4wl3VHG5SKtcLbouHNiXzJAgJYyZJRyfwX
QpgyMSbtNZdUgKp6/D6i+v/aoIclA2E8mJzQwpZEhmACF5C8/zZyeU+4XiDOBGp6
gjuGAbCOu0J2wpiDQw1ZMgLH0qqPd8+QPLEoaP7pr+e5cXjnCFr5pigFTCOE5CLD
ULuVac3+UKiCX+bYFG+m1ovlv5DSREFVfOFFTCsr27mDrnbXoLPqyiSbDqypqvV7
7rvgLhWZcVLnAaXv33B0JJXXoYh1UxSbkX3a3A6BVJBfBJzow4FFYmC9jlaWwVFM
uTtReWQyl2SHKIqTgpXRPT7VYl7J80P4nzlcq9k3dhv9xUGLzGOpXJ3S2GD2uXqk
02m1mX5mMmtcghKgwkp9LUunr4RDF+NwxXVO920P9GLwdpwBeTJgYC1vxqj0HcE4
x1ghhi/zQ25LZBwLr4kHcAGofdLWZio2Rf2NzrJ2/y+4jaMg57TGstiXsmXXph1X
Zqhgo2OjncFttxEEKDxdifWvkzexTAoeI3JkXxdMzka7zZbLQTpYPDwQ4yV0NxZ5
5IO1PpqnC7RvS3Zl097AjcCLwrBGlbMIcPKrTzoOX0YsivikeK2+F6PzAg5W1XEk
N86yYLHy+GQo+T+IkxhHod08orRwGyiUHYrGSYkYbfKCWeE+eII/vmdSrrz3s3OV
WEl3iXsQBBpyHhQi1jToVtgGCI24JcBxsEEpnlzH8VYc3gekS54lReLbt4xAvqEZ
p9lEzj+ucMInnOXqH8KL58g7+P74/IR7ZPA/WJmcv3rcrPudlbBQX1ltk85VXwBa
WaqGJa9/Am/VHKA5ZN8sNbfoiblsG+aUpCToKt2XYqeOT3aHzGwMbs712kW6QZxI
YaexyEBrSqGMM9i5PWgtV8Yih3/M9RWeoWLpg2U37OfnoZZhH0d6H5x6NAjallEg
wiQEUP11bewRI63+IvcTDrHaQoa6pMx0zD3gKVDI9AbkKHPw8zWQ0CJcXhY0G+GL
rBtJeVceUM7RRFmhklMOkxCpEj/AshFmpo+cVothat0z1AZGoQoThjbjFhTFuaHl
h54HGkKDGgoTx4NFUzVSMvsKigjzYlz75+3qKM2My6PEPhAgNixoQDeMRt3Ts9n+
kaoVBtx8G00w6BumIGukt85iq4YVX3kvjvHuqRPUKWrIWcBaDJ+NdHARzuUnaMoW
F+3z8AkKNWYqrz4t9eqcDCxOzrzt9q4XP9sBxTWJWMdYr9gf9nyx4It/tge00VhC
34ug+hCjqRyVLdAd3braurSqOZjhcFNxeFP/swNA89RidVAHvYN9FFL/56Z9Ng4M
dC9UZhbcXluOKcN4AJW+L1nNE4/0vXH76xbxQUGcW4C8mYLTLaEbUbvUEuIVxbZH
5Pixc6jaa+Ij7tIHaOrfJIDDJonU4UIlRUx41+1Gg55x4wRT2FHwMONTHfuVt91G
JKS4hWSu25nQEUCkA8oCaAx8TkpsliBHANtE8Wgq48l4e0aeKV1fHVThFB+c17vZ
pcjubzMlld+svqJEcfB6K7Jz33BovYZpMQzqXegd/NfD/MFkI+/J68H6RHXczJO9
1QOElGvb1eoes4ikAVpPyayM19xi+nJ3LYJO14UxbYfHv6BYwEYRIbzgYGGXqrKU
irsztJdCNko6RFTEbtfn5Z9ko35TQvxSFT8rU3ewZ/Q5pwkHFnf/YPef+F3bWKOW
OJcJGY5IIb2d6K2qpdrY8zQxZGb4Xw8+DPfpvZDwnUEs9HKUIt91xY10VyiKHmRY
SNEQGQjy4swfc1+xgInH75j2SGCLKwbyivRUmsxTWba6zOKKv3X990C/NkakQFLr
+nPMAlCxW9IKxSO3wI7lMMjFV39/40PIcq2rev2Y+yP+NmsVeRQARC0QG6IloCZz
9jekrysBxdya6Q+lzf8Dnq0lVzPo6CaYtV4e5dvB5EY/uTPp3806hpHsfGbzq3/H
mSDmbha6NmSO5IwlfIdDRUXFBxx2N+cJ8cbOytxxveyKi7r72smaAGX4AMCfKDC1
Wt2aSfYvhfB6xVb/t+gGUkfRlqBvtw4cENZYmM6cX5tjjBHH8XrvUqH81Quy8ZOb
/ayraTNLNUPi0kSi/DrJ7uLpyQVYu7dEy9Vi+JjpIrwfly73OcGfkyPK1UTNLJC7
ono2RKX/YyjLv4YdXTxZP+2HQi+QvkwN16G1ExkL/vGurBZc128wsTxxcAjAa5oV
XCE4y+VFTJ8xdU2GJPgJXwQgmrijMRzn2iZBJb8lE3Zsqj/rSXNVxuurcJxhnCqK
Nn0mt8Fm5kpfriwCIr0XgFCnaOkVmvqE2AZ5kiQv+xOEG63YaRT6Vjan6hNjWMD4
HHAdJv4uEPU98Yavx7FH3nt2g2QSjXwWueR35EwqzqCMZSc61NogT3Aqolz/jo9V
tiaEVzR6MmoEcl+ydRgSu53q+qIYbOUV5Y/fCQSrXSYW6RdAdn2gZYerIUwInFLR
0hrpmnJnqxfFwU/407SFVeYH/HslytSjxdEfoYs8F2WNcgfobDKMYKZ47pRtn34b
AcUJtHGsZUYPaYTWsPwF/FxOZ2jrsc5AJXrj5I0NI0MWgcMHiHCf77wfPfMGvsX1
ysMxNswaDBitYKmT1aYCawwt4cNegIO7KfGDCrFhEjgNDn/LTLh3Cuc+PbKte5Zh
l+hO5KdeDe7KrFRtah4YOn36QB8t6GxKw076cSAYeqzUxuYdjUL0LSP+SGGB41Oc
CEI0zFBx0q5gDBTdpB9GDZSyfMcaNFxQWuDn41LzM3osYccQtfs39wC/wAx+ifwB
+BwSNug1cO/D7QfCJkeetqWAqbG3bInaSjC3FzNxdVJyUqTWJhU1Gj2bOleADX6H
8NLjtH6+Xy5VHzBCdWT6iCfTpJwKmsA275PP7TqDngxgzbWQ2/GZ1edu9oc0nKdx
KY5OkZ+dK94IQxCfGVSJB0e6OKz+2dc46JV9zQbIp/zXGJxYKWqVPLql7f2JJIP1
vI7Z6Lje6cXvgMIKeCOqe8Kz4RxMp5MBNllJCuRFn8qG+gPXI6+Dy8AyWEhc0G9P
tIZM4fAl5tzatqQcAedV9jZsZXoKUKh8BawdJFcWMQ0ORe7tC9dz3Q7va1sdrmK8
EzL0nBrPn0nwiawC9njQCYO3Cj5ljLj+x3GfqDAOgNxdingYDXS3AxgI4OWiniYQ
Hum9FBg9XkfmPTzuR8ZEJw64TVLhegutajgABoYK5ZbdDDiEYBpeBXsgeEs1V5qe
MgirICu+kLf/8TZUY0taSnjvFz9CV/Ikm6n+Pon2vbB7koCgOoj7cDY6CGjsauGn
FoCc3R0V30OKiYiP0Lsyuu22KCmq4gcwnsMdu/+axH8DyRZxbDqXKus2zq7Rsgx0
UTKI8b53QlOKDrQwA5zVAeQBloEcJ6kHbMdXn1ud7qtcPto3aQhZYFJdu2ZivNNN
+b4cTqigbjnYrShBuC3q/X687dPRcQA3gs6rtdsn1261tX2p1ixfKzaUkooN/8kt
ndBgzM16CJ92oWnIDCEqCTWZEchoN7gW260l244YNPqVScqRKECcTwgMP5ReAh6O
YF6fvGCKZEn9hX5D5JoAqovvy8RW1dpOqDu4FGUje4Ehb9hFyDTDje0aMtZ7Dybf
mwAE3iK4Eqhm5y7xsMPBNthCa81BV6jgGP22m2rHmY8DhFvZtiTnTevvRsYyJsQY
e8P8Y2M5IHv/hAgWCRy6gzdgdTFJzn9k+LSv0xk9R5Cb57Tjf3/gV64o8qRMKLxM
lOEJ8r6BK5RrZvdRFx2T+PQRjHA5MvEZhgrRS5jBF2tZ+U1UGWb27SKyHNAL+ILI
vJUd6IqkPRkzXBbzBAam8l9XBmLGV5iCEUfT8Orz11vwHc9DAI70EtlxpXcvTcfW
MVQsmwSuxp+TppgcCEyyRHG/8+iVgXuXzcxKvq9J1+hJJ8T1nWu1fSsPYxMo1ItR
L385Giw4qqAH9up/5MDORvcpmu4OHNbpy7FcDDV95WPifJn5JY5QF5VNajooFA33
shzD+NF8kOAsSIq/UNayOt3eFqaPbTi8J0gsz+qI/nS0f4yQ+GRdj7ufO+73duUN
+7PKqWW23To9fXNgtYD4wg==
`protect END_PROTECTED
