`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nfTz34m9qHmLg96x3+YYI9icEDOC9Y7mzixw/WFuzDJ/CRkX+cXX/XGzgqdqBS/M
eXUo47KvhDlyuEudQRmNENHJnIa3Q1HVStdGTx9p5ymHCBS3gRF1LD/Tx25Xild6
5exjYG6R4WTCHBdAg3+Eo5KgMjfC8dRBENedgQPxHBvBlyOVo7M2FXAaHLuKJlBa
0sRT8N7dv5R1xeb+ObPBkwOdjuOGY9XA7MrFuF2/g1Zp4qcNZH1EgFEJDu6dVWiS
KeV8iAmG0sMSEzPrgRDBgpoU5VaelZMVuDmZysou0j3YEwf9YT4Lpa4MFvX89wUr
TAAcN53ggSoZMGjAo7XxVe5i8uHsgfE3QpSSULwlphNMxLh0fbdb++hj9o1dwNwV
Eg49X51R68WYlQoXMCV2SawEVFAOYcim7e/9qFljGVXcJzCjaqxE24BPwh0v3uPt
riWtp4Z4ggSfRX3Fr9/ZYVgc9Yp9GaLC55rPQHfuRd/uLBuaHeUvuRNC5+pR3Q8F
OgK4paMtjgigakOuyKLGcrpcWXXvPlSWhTtq6aH9/AYG1EWh94CiSqit/P5FogPk
8KhEwlmSp1USjgmTa8kVEJ0KAIbBUBS1cjDWtJd52IyAEogRKHK9Mpy2+zijEQYi
6SU0UmW4prDN/cjkPScEGqSM4y1ZqjZH1HzqBmkXUilWF9otpndiGrQ6Gw30ioPB
fyEmY2qwljUFm8R5DPsI/KnWkLksS3MIeF2rCEVgWFYDwO8nxQd7mWCk8gOX8b8A
lwmghk+Dq3UTV26OhZ88k2oXsJz6yj1I42RpFldLgYyDpIHbudjpCPJSvT7PKfGo
eRFqOLFfDkEiPXovtrjY5swAfyUrql7oSyRPainG0FTG1CKH5ahYgJT7jCuCug22
LwJNsrnTGouJBJ45QPV1Fhb8S/GQnAxGH5K6IZyNB7m96RpzuR7pcJJVaIEOMFPb
dtL2M0f03geQ4y1vOaLsRjk0q4aEkHOMNulMmVA020vwkOkeVMzcSSS3v3e2dCpK
JIzbN3uoy+wM7D/XRj3NORG2NxqiAwfQE2ZptseWWlc9A6dR6YmALn9QamZLQlWg
Yqv1rQP3qbhDjQHo7jF01rRBfKC48bJZ4AoITLEFee4=
`protect END_PROTECTED
