`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oodv/1tCgO8+SgyoXiU++Se6lxnNdghpsdqwsnkSkItpJ13gEUjDd/z9uwVdtPh7
GFW/R+zwcaCU1dqovw/UTe0168KT3hMNJukaQUEtGECe7Mey+PbbBzvcNNsKd3Jb
+mO1riJcN1ih5AHO2aSPcIeCnNki+aJCHfa/GqhF8Z8Y6HZFVyHuCjzaK9L6C9Ju
oWv1kzhPEwhAfP7Y5NPtRlV037+zCEiFYHfWIB+Es0Yg6vWnhv/w0V8hWZ8BmpRC
ymkRAplUt3WvSXCPvdRkXoWd58YtYgStc8Krqe5AqxLKU4NLujo4DMZYC/E/H09u
K5hN3iXh1Jzd/rrlpc+SoYxY9+GjyX6ngLmaUcE4TltLW23LvgmrYQFaSlP7jdaQ
3AoLlvBpHw9LLSOAESxCizqr18Or4+E0xKyFj42GT68GGjHPlItnnifUhjJ2A/CX
/sJ0Jqxs50L0mBwE1sThw96f55GceLD3Hb9pxVKHU+4cyT3mHVmx8fujG5Pxguhp
lt5RBbk2l1Rv2BPlO884nDrFub2gS3cbvLs8Ke7VPLb7ILVYgFg69AMoeiHbWfdC
7/l45bS8XxIGNfxEHberojVtQxDUvt5fHjgM9YYHANs=
`protect END_PROTECTED
