`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iVsKTRJy0FrAK4QDd/A1UF1tcvDnUdALAFVljRIAhSwyJ2Ehn4b0NeLgfmWuxYmf
dAT0cCJ5iBFBH9Doi5rbcYvTAuhMky1dCFbgMOoP9yiW+P6G1dNaKawEIFVBPrPP
sa9tqLTRTZwWvVI0ZUKRvOge62VG58plf5cpOjaEg6ktEy8spguFApecxiAriqI5
1IvyMBrD5wA5x2exK7GvnSM1WAbdftvZvGSRFKQgfI/JVNlorJw1xmgDbIIDN98m
7zKJkBWEOK4HAB6zPJLSXflSwAqMtn71DAOHWXeHbYXz4XJbW6Mlg8l3UDBpjbRX
sa0XjekB+L7mNZzioqDPzegzlzOtCQ7rWX2qsem2LG3Oz0a7s8cdjQ6hVUwPt3O5
W1ZvIavx846lNw8yvTBFC+kMFCGWcWk6cpIE2WCoThSPrHHc6T4crPYWKupSDhwu
W44YwSEIaLAt494Wyf4zjtuR8cVchVDAY6fD1k19hSQ1kR/egKgWTg3Nm4o8jlkI
eimbNNg6on0yfnqVIg4+d8R3cjbQwKI2aWM8TJlhnoTZ12k7q0+9jbeAaS0+R+aP
UodRNfK59XRJi2pibJlwuL4ZGjzYk+d+tsLkhz0+hzG+pkqtQf5qUPGMRQm1fdgO
y+Y+RZLEnsUM3lP/ENPcMEk+fePvgvhBUpf0XDLwR0YSmHBQCq43TGtBq7yYhphV
wuf3f22oR+9FDNcsjVB8VzDp5QE+YMhOiXU7OfPSjSmVZQR9EG6/r9pwQ2RBjlHx
1yWa5BDAqikCeDVzTVHZ6ntmNjPxdXjj5X3dpK4rruPLsxUG4dHXhn7QyOTJ8pq9
5uXyTuT/un88zBE/M45GIMSgi31wjIL0fEISKXLZOXc/ZjMTkadSGCbTbQJjPvGY
FR7OvhVbhiuBc2Bcc8iB9WG4htmY3aV7Oh6dbGIrYzpu0jC7/XjwtfuBp+eR92pd
sMAB/PlgJG0GGFLrVjlic6NV8EY5NEfXMjntkz2d7ssxYdcQXql//G7T2aird5No
QxudkquI/f6j2JacWuPU6z2iSlH9SAMpeubExcwtm3bTqyXEpMAtreIrzKrwz0vg
y+a7vTHI8p1YWwaBPEHf69nlFc44TwTgLzGFoFPJ3zDyswBrXdDL5ol4MjC2H4bu
z3MmIvfyCWDUxrcJp/Jjq52vepgwK0JdhZnfNmhVYtUTAB7Ioj0qQatZjwmmX54o
E7hAriRJXnIafy4HOao+KsfkeR+DADGaUHatKVN2UBOo9QH8snI2tLj9Tee0km9X
AFwwmOdopGNKYk8sk6AtemolVzBhDBlsPDLQA36Elgb/thBwSrWin6WpqGaLRZno
OnISfsresw+tKs3X4dEJlZFUIUuOxKwXzf5Adypx9st0bluy2A+eR7HdYBpkChmH
Q+DAlfo2fvHGITiOiuLCmaY3vBhU4m5adFyPHQqdJ/Ot8PfuLIZwekWVHjur9c7R
MPK6eENBI55YS5l/QreokpqmuMvLps8+vMiAnNrbnxEYSE6IYi4hCUFz+9vYh2TI
Co8A6vykJLN3BiMuWRZ6efEg3l8D/yIUoPREijWp03YHzWO3QpnDY7ySVU/P3HUR
/uAh9TLF7uowcU8y7TrhZGOglZOI03cnJYl7gwTdERCsyHA2z2Fo0+JNpWWpbmGV
GL5yfGrqLUz0MD6LtJX9oOM175gv/AXfUPM4fXONXuV/E9NiUL3lDiVpw/u08qIX
NBhTQs7moMW/r3weK/hyAuIyRPjoiUceGxNkzQc+DkR9V3kkdGZuRH9WKD62ci0K
gVnK0hgKggmzpxHhKbg3uTv5SHS/u3Gf1qvLdzZLPbg4URa2yyxwlSdw1IDTz+Wc
lsmmgUBxtEjts0cP+eJbT7g7z7mjS8k0NkcVpXYY6YmL+k7QjJXHfNu8P2GVD3TZ
dRe2X1kbrI+J9lC6SGdCwuI4FQvhHPCvaf+XKBwP3hOt22+8DCZSFlbcPPuGy3lx
TZ8/tP2D9wxskv4gv5NeqxTwzo20C8xqwRT6OkiPmgGHEmo+dikm+kgdJUjJG/F2
ufqO7UTi23uopu503r58Nvtrnuf6JeEXe4MyX5mZWbYkZjGjfe3xLEL4sheQQDVW
jydY2QXs/2donA9nkpULDKakOCfOH3TGnO9Z+lP9WC1xnnhv8B/swxE8LLX9f7Ns
RWOkGO8hUzbj+EniX1XukPt1GrIST7ICKqwTECWDOA1TmYI2gGWcKUPr9M/VF29e
KDepLTRVoFSWGovPN/D9qva2ndtao2WBtxOU8FgnOpNarWSSFSJVoGCAsBwf+BE+
JiXvN/suGvb8BawYDm6j6X51i2xfw4dZIXaeR2g9vOnDWj4txkS6kgFr7pVjiTbu
7aISMX/coNGE/X29zlO69BbzlyNyWL8Pa3JeuWjZ/3NTvWnDomWM3C4nD9I+/3hO
KZ2AX2Iwqp0Z3D3HI8VCGTKbT+0IRr0cYOSd62OyGrn2YeCbZX6WIExT7j/B4cJ/
e1YUgYZXyvG9moZIn+PTRX9zjyL0u5f958UOsmYz3kSynPQgscmlZ/n8HRfHxn8l
uW73fMjo3hhCdkjgHcPHKi4zV+83mWHSBUZ5hO3oFU6D/t+g3J9kRYjPcDS+YIJW
Vmuo/AMfMdAkQfyolVnogxLNgmzT431vIikeKqfXgwqQd5PlWMPBo8YYBQL0fUhh
bx70SrAlfcKusKnMiaHc2dnBd88xTzcOGBK3TKgQ77dY4uiuIc7eQ66zU/ya9NcL
8sWlCIpXNU+xrEr0ckZXXNf//2u6HmV1QYc5i9PG7XmQdg7AH5nuFXuKckstTAIK
4L7cAgBLGHC0DC+5j7kCeQRcFZ3cE5730GrMDgDXBPq5ZkCL6yEvhG+Lu2IOScwh
sFGURDsQOlSIjp2ssaSLQRmoLtb06SCbs4AfLVv+jZQSN6Fntrk9i+sa5CDoPW5c
nHBHK5T9FTP/pBcs64pmnsJEv6JqXQcB9r9Bq2z1X5AMr8l3tRxk2XRD2+tCLZmi
ZRlRT+r0IDE8Gz5sYZgdyluj6pj2IH7LiaBAGA0DA+lch3ghOW905J7KDR6ARpOI
BVYfLxQFC7u4eQjbiMNfHOKDw/oS2agNQL08HtQhKEUxnrW/wk2UmqwhCabX4HA3
seMiZ1c7T1T+8QMU45rcwbDNL8ZH6LdUKaKeW8nHM7zGsckJfGhsFFHvrJO/22Bd
t87Qe5UDjd6JQvjmb14XIjp5Q3HfHvqyvJ3N2o83OozjqwJFfmF0yu01OVVRHQqs
QafMAggWZ+qctwFouYD730WeOTflIXAECCHfT5mzns4Vql79BHMrdaBW7WHG64r6
kEzFIdfNHIb6flgLXPxiyB+q+AiuM9aa3l78POV++sJLQd1UbpyapcCxdB92bFK7
d7VkXldEQ4Lvi4HupWJRdVVXRqz8H7DRECOcaaUXTI4qc0g36y/RVVR+vNwNKNWP
GR/b7f1+uw61NFuI7nMn2TNx7VOcs6WFc2WHFBqlNyizEEM7kK0b5QuSqjyQGeCc
Cw7EADxt3/p3VVZA5yWRnjlDYYT3NjFA72nBgt3Lpz81g6Jl/FqzKFFWF6C7h3HF
akZ4Zo9R2pmXqvrG4adZ5/0y6jK79VCYLzt3orsH6bQvOTpcBfvnBFWhs5SAM5dA
Ua6suygQR6CWaY5q9OV3YSWgF5cSayOnCH9jKU7fq1bv//a8h0wUd8L9qYnF9Bm9
xbOslLHP2zXMHY10NR6E2rlNjv/J04EmFm940G15JWb4RKu8l9EWekRSvHFcRZbf
DfqWyX5m6I4FhpO9UhmNGC4vZauMIWp/B6FSxd7VQBAh7Fg9qVbERmMiWY8ajESV
cauGRYyZywLWgk6EeESouxo9OTBx3b66p8+w/hfnmpdEYoKQxyC0IPmplAZj18XT
f1ad4ZRkDCxxFS77xKkMFCsJKgnKbnKnTg0MReGxbRXjf09Yt5RMPaxiGdaBtH2a
65UhNBVMG2TcvSu4yOpeyB1geq47biXkSVC/4z3I0BhYuAzQtH2imRezUXBjnmhl
79r740DUKpV1/6gkQCLLOLpzeYIXB8qL9P2hsiLKL0YmOLC1RCRKegzofRhbmCnM
79KaHOtreDkcXg5opVhG1uXOxk23XdNBRBMtoGyGmZwfHWHRxt9tmzWpbuD3v2Fm
bvjGYkPmBhsvFWepiWk6MioFAwgeO9q2ilfBj6c75ItKzk3QU/C/oOTqcljHPtcC
Um9yEYXMPogjDvBH97L7mD0PLGZlNOJIG56PHscQd6FUsQFAhX4lUzQvuj5Shn2f
/7rKCJX54KKK8A4hx3hh+tSkEDvv0QR3tpA+feMbmhQOKqqL50sM4WiPCyBfO1aB
MvUcL6wcP6DBYl6M0WkTucY+ruNhzt/7IPxUT83h4woAaYvLSFLNxfr/nVtA6Zzy
FAU4S+7uX3ffXVVbOJstUsJOZOBRmTNYoJDTnmNa2OWHie26hWP7pGJiyyHLOcn2
yU+vNFHrVuGm84SRfbNMeXEcNIlul91oxq9I4Q+YgksBlLtYMWEAzWeH15xR7COl
2YhaZJUuH57ZJ4Zo5bXzL3MNWaYUuB6HY1+0ZafonGh/R+6NvtYWQ4ZEYz/mGlyA
DxuUKO8yyxU5JxhJf0J7Q+FC77d6yjeBQndIoFXb1fl6wpnBAGjRkVxs6NZWeukY
XD4DNm5xCnGvhNMkL/8xxI0z53uKzT1K3fI/XS5B4d2VI1tf1UjzFiXOWRlt8cc/
zM2MEcQKpBXLJ6lwA3VB0kX/dpdupFOpFY3/2bkEheb4jmZpivgbqqftNKhwYAy9
y7K9tt5Z7AibF32L/t+od7Njx+m8iMRpQFhacMv+WHQ07zwAEoQb+JPNTULQAnXg
KrBY7V9+D8ZPAgQ3W90DSk9vE+c2/J9TrlnwmS9+thJPTRvHqYcEq3ToUPdt7+kV
qNVtvcCYz1rTuVmwq+4ST4BhFbXJS+C9qCnsvvmVlkawODmDF+krwEAEV19t0yu1
ebc2JdpRZBRnF3P+2hCXXqg9Xry/RzvnAdQg3b4C0qT8YgLwuX8HprKT+AFzGgik
q3hLRFmbXxnIdlsHuzUyFFe2hmQ3xVbfugkm56/UJ6gQ3DU0RjdymhlPrbC2/dPK
N0ZoyxJMmzrB//tpkDEw5yxYTSZbas9WJo9SOx9AYQm+RC+mlHfOVAY3lXLQuX8z
orv3bpddosOke3Df1xI50CYDBiSfNkI4Cq6+cdC9Slo0691+l5e1eKa67VW5mpIK
t59miA492dOO0C9ruhNX5t/7zfWzdGfdzsltFhJMQPJhGwU9gvLPXAFJFBLZuXXh
oVByjIDejsuCAUNXPdECToUwg/M4qACk5Z5sfoXFgAcvQX2zgVYtaXaYIrtcfOQO
F8w3WWunIOk0qy4J901l12ViBvlphe/fwpvCAbMt3XRd0HT5y1x96Cgyo1PFziVh
A6YGGs7LtIiLoBwIE0StUNY1O1f1vVC/tULrQqcDlQLNgEOViCbl2rts1l2dL3xG
OPNKWxTfn0b+tHyiL+A5n9alPHM0+taHBW9JzMM9qm4hxzOKDaPowJwjgXmRiZ+R
xClp7j7/NcBN3Cf2NeZ+KRSnFUIjJD2B6tjoh+xdbzwbZtbECtcYtkGmN+hHkCIg
5j/DyuIjGn8nhmyyYKHQVOuKPIspsnR0gejGbA9DPasKpGn/hP7hos8m0lDT0Zu2
qdz0pmlRVhy09FLVkLkTCz+Q8oMdZ2wj1c41nBvsdba4gqqoE5vI2FNauQKwtxuu
G+ObDSKfSyuXh5H2X0vJmDmwbBtKYhwFmAlViXkL70MtkG/eLJPWa2oSkul686jg
gTUUUMthX5Pvr4BhbvmHYA9qCQiJXj+cbp+zqHcaUdVc4flelkPOw1RR2vSsdrJH
hmna+DhL7C4kHtkE3xgauWX8v13XUpEaOFGzaomQ2hizAWcuMk4P7talf/9Z+5Sw
qMNUq3BGoJwH6QIJK+5Q5G3QveB301TdQq51fGp9/oVwhLx5GcJoHNxv3w6tuPkO
vk3mPAQxuNE9fHDmClA+uuhhkqjAk1t53J6lwh2zYUI6wueOVrF9gWZtcSnPmFYd
sgPofsRFLpQ0CpC2m3A4lDSpt5qjs4eQnB9dqGOaWCZ/K1WfkzrNLrw/OXnDoFHw
0e6lZYOpSQQWK25HPxC0gMC8Dpl0UKzBDHzRKdW7ITbxTGCzdYb7nDpeBcZbzB7f
g5QyAu4vujrBssVof7V8pzgSuvMcxVHingFLg6MSmd11MArpY4XCBE90H7BpAM0v
dcCgzYX9Ahg89Iut9naaPYqygHV+lcoxG9CA+8E5X1HgFljdxOILguUn0tTURtlv
irRSepjszfdsS9RYYdTjouCUYaalU58v+e8zkt3oZKeuHEFK4kval8cJJ4uhDEiG
Rf5Co0MRJ+R1pLQIpl6MTLoH6yB6l+BPsvLQYV9NbJp7IyjL/m5YKcC/LD831QAK
NCZAxFeMpaqTRNOzhzWL2hr8POucqILQJo90tV4xSK3RPZn5mrBVaENxEGXUf+7r
uKEuffiZuRfDyXfPmAy02m9FWVTU+qbRGlBbBvau7d/keWKChHMV/LBkx3oiDl5D
x1VKjrR7wi24+aylXYNu2Q5a0eyGyQNYyX0833duEqrA8j+jcVtXqgzyeOxxt1Ja
3JFEC6E/g0LqI6G0erWXPhR+hfguOdHRzft5jpsGp7GfReQ8wtSMhKTfROK3Wxpu
LFWJMdL0inxvtnCAZgX4+i53C/IWUGeoHhYRRxNqkDdvYW23YeHtiVFih2JOgOy/
SPjmwwsmntjdhcyPP7e9xQI/dvWWXQRO2pbV5J6q11sh0Tk/+TfdSgV0WAPcxqzU
H9eJTdSmvLC/AmRiP/ZHBAidYdf8hSc7BH6y8qQFirwnR3rGa/jAEpkZcd6XC4I/
Auqdz7yxR776+YjQZ/c978q9O2nxZwXyPxZrNkJmPBaNEwl9PhqzacsxgWG6EQww
ftsZqQJH0Xz+zJZIoFTwcuUJCyJEy1qBYIbIqOzYgrKtHKt6tpwoGSzsBL2QvPpH
AcjxEbelgymVJVXUcxW+kwhHeR2y1KIoYBbM2t5oCnMo4A44u5VwuzoHAUMx3rRM
pQGgD7VFI20RMZmtwgDHM06PcrIwKTypkQUaKyHEot361EFLw5YGlpSquTfoYDox
jUvAYhuDOKbi4Q9jLRBqvZMJXrrvMeOPR8pTd+wcBaR/yzQuHh4KUXguwsXQPPXJ
0M3ofNoFB3Z43Rwmd685ldxbgMHh7VGH+FpGGbcQCp67m6iPK06cpvC/fviApTjQ
U0im3uxC4K6qGsdRMx1ypSezJ4kYQ8IyQxApsaqHxKrRj8ETWx07rUzKgNf4rLhT
1TBQHsky0gPZ4UTqyxuwTeqcKcxwVVxVSrd4cv+bpy26swyhEzs4k6qtt6RsNEb3
lj7gtReAcJf+n/aHQKp831bnjrhT8XRg2SCOmv/cCJy6Yz6fHp9iLE2xqI0R3nle
Hvlqzn65Q//xGARFBwqNK188A4v+SjTtCUMW61j2XjmWYcqGAQW5OIvSzuo/w3s8
tXfUBzIvDci0nVQiNhBb8+QZPsgMMVYXO37U+Pv46nkPghkudkueE6w/zDB+9IbG
8dWq4MpyA7BFCTucGyfn0r8Ksz7wQT75scb8Pz2+8SUZ8NTTxA+h+u31dufQoE29
t/ma3zsnH4vczYcM6UGAbtjVRhPvkiojB6GaF1h8TCvZJjcLHYencIpUv8ZyG1YP
9V5494B/SB+TcmhLG/OOFzfvlrgkhwWCwabvMK5SnRwzPrLT5G9B/KVU/ONmVihn
GDKqSUXoZlxlSnHNgvtq/Z6I12IfxcK4K4N7qZmIXbYsxdFiXhn5SVcWUN68RlDl
3nFWR3ibqYh/H4TDFfAm22TrtlorxTPmr4ZIYszrcY622I81Se5nq9unHOiX6NXJ
qpYKCV30AtKkDJW+mN5p8KssQK1d2LQejWncgxP0CvRZG71cLQGUh5fOZSwErglv
0FtyGCayi7SjK334p0njNtg64Km1r/D8r484uVIIOHTW5G8SrIhe00k/pKVmyLaD
RL8qLdPsvm9e6tH1pITfCsiFpVr5iigybkOFDxZa0BPPDE/C7LPkuDg07OjjQWTg
jK0ASixI8xh6y8o/Al6yptwCA8VOByZkb4SKR+wgAO1LCmH8gLa2HU3d4O9hCNSh
kOAFc2BMa1guhwWs2s9VVqP2+KPYd1ZEemWYbOV/5Y2LftB+QUXgUY77OHbHhUNn
0JsH1vYk8BsOYcWcyK3dQ6daPtxbYBse2vox7Wucf8Q7lTQcFp59IhGlg4vKbm79
gLB6DPCEKVrpC6CuTe5ld/YZXLyi5Lc/CeTaZAAxoeRk6/e3NwQUGGIcNk6AYgCM
r2vAIG4KAwkj5j7Gzvv9VAIb5Fj3+qZqdsoTv6hORQBgKP4JaOskAw7pkyRYE2Nn
Tx1XLQv9ZRGEbg9l90U3tsVtGjPGuSYFtkb4j6esDbdkqyN+EDb9BqaJVzjoXAQ2
yOY95Ft9XH/Koq/vB2gMtelSx/mR79fKhnVxJFO/a4B8ZVUGC2/NabRTaWk8yXRn
w3OxiRz3N/x6oIwkSHiLTbWwlNR5SZ90ZKsJi2+WhbfZCH5SdK2MVOl/fW7qtw/a
iS8kufqRCNpMp4TW/MbvYsw0fAM+Lp1xU0RKB2s9N6vLMbc06tbOsXw46pzyTP9Z
PuwtHvOx3W54D4rwX8NxNGjyODHYS+71lmXDT55TRmOqVoaelvaDt3FQ24xIpUzU
ci57uYToVPacyBs+mNr+fWWtJwEdnKlRulJyELSV6jQjc54JT/OlpUVIXpo3mw58
95ewgLZ/2W3dS7+dK/imQyMWKQp/NJao37CZOeO5fWJmInMEWYCJdwMezJ3u3W06
vDK1dlljkZW276lLNq9oF++OTl8iKonPW8nvSSAG4uPN2VD/UUG9AT3d6r5xYgCY
vRMoSg905NR5d1D8TvkV6byPljFNR7st3C6u/pN6TBsVyvl10oZV/mqJyPLlJ3C0
pQD2FfRbfQdbinFvP5MJOGyGorzIRv9e+Bii8AoD/3ka5fOvb1mHV/Ff8ALMxJEZ
20oaW6R47SlEq3PKACNVIZzDCeNGOwevEu1ZODDRuRGWHC8o6Yfcp9/h66f/KWAv
vdiXywpIrIjxGKDTmTFfn3ABViAjdx7ckqAQ9LuBQ6ffxJqgUmgpcf15aVsHeeAJ
Ia7DUMqZgA+4rtEloGOeSm9NyS/DPzg+9TXxAG3mldwBUyjDT280lKGH31+fiAPh
4smrov8++SkCSWrkaG9gqWjy1K1QCTtVednlA0mcIhTKFy1xMHivbrNqOJVsHHtd
gbKHNYsvovUvTQ1RDoEjRE4hwFKMF1q202ydFAfhT0VdF/1eP61UtMU9aQbYFmmt
fTtCBjRbas461lxoyjnw/y6P26iAYpkI+s5tWnoQ5uZ3BvLPXolQMouge8DoRue8
enqUZSzb1x6h1S6bh3RXhAQsAySeHMFNPDiGQwusARs+orGjTYmwXuEbYKVX3feK
Czqm9w/8pl7Yhur9t2UefXRwLmA72IBMgPk+JMr8m+wK6j3x6OqivRKcZ31Kq5rO
cpL4ncK9WzlEgZyIevbxzVtx+tl+Bw6D6+vYED1cjP8gI0JhHZPOl5R0EjTjfj+y
xA0CKSazUqG1QDaumAYdl4tTPwShBBaaj+nqUZCJFM3ZC4qQEgL1xsxO1WPk1797
yOgfCAPc4B/dmGsD9ZZZG2I1PGK+wKWopOSJFl0V3ygTOjokXoYcpBhHxQL5j5GW
20faMhVQhef7SZS7LmHfhwH/XyxZ6K5HGf1Ri/qBVWdfWAPiG8JA6iS8qKuR6StY
BjtqI+m+mUm9pxBeLvrH/y6AMh+Lxyh1+B878mUQbwCOMy8MKK1KIJvePTKbW57H
wR7ct1O5i/gwomZFJT1ZcoqAlLNr52BVNmhG2VJk6c1KB5DAEVEN4IgrpZEcttY+
SsBWMOEmEAjS5EPNUEHvHSMvyPQygH/ui9Tnf8MgaOKPgqiFYWuQbZNePRWjRmJy
osQhFMryYI1qXG+wB2bqApGrG90KAyLOdR1r3AqaW/4dp4zf8KIrbfNEeKxtLyPd
JFHuXpdDtfdayxxAgPd886DJAQ8hpOzeUNLzpmhVGN12A6AbZs/pREyykox4wqmt
IB0zTDJwvJ1F87M9GHKE0VjUMYn6gckCDBl1V5H5KVQ2ZKvHfB2i3bysQmQ6vs3G
aociBs9nvFhnpE1B6U41XnfzFgceRJsNAjjq6XH3/V1qf8/3pj/4ohxNuAFRcSWz
nl5T2ckNhBrqcYgJv3gbBo2SS0O7dQlSuQW64lc7kRqZWQDqbvg66lA8expIv+dh
YZ8gD7nu/1GVd0yXDlVBxvPauYPKdaTTjE3R9AyK/bErUznNPpchueyIyWwtVAsO
ilYqYi99a3u7nf57RDcTmPNcoZqa9txcxWVML43jpwuGPVmYhrV7gEPaGyuwq94O
4vFIgKcrgF9d7O17EvT9FUAm8osjc/i7s/mgv+jaD3CTCH95VH9bg/bub96lwk90
Q4SeCJe9awePWpYkLYSoDPae2LxkOZOGswg2CdgbdAXtJ9J0NosVPFyFCRX2x+TQ
fsDF6balvN5+FMhWqezMWaU2aECzQNJz5kUg9ectwmviUikrML6qjh/QkIOLuaTD
qAvphVTHMIR55NS+01qf3qMvdxUEhcO6c4SNq86xOQuRXpKL0QDLtXZ9/rAg2ArC
pFokQ0JCRZqKeRoH1lbLReXNMg9eUA0r5y8aGZYkfEdC0G40bsj1Hlc8XmE4NrqJ
sq9GQuOUo8bBNZ05N4lA5ZUQArAdzAYuG9iEleajFerZaoyMgMC9ZyNeow6cORLC
BjLkxPwyz24Rzj0xGoOHr8qhlV0PVvYL/EbPWq9vVd17dH1UFNmv6VQYPgwVXqc0
c0ALPoc2ZdHE53tqr80PyJI/DOuP8WY1+ORGg/vcME68T642pkQwtI/7QEW0kWOo
yb9ihcU0GnAeLHy7IV+hClRP5nrY0oObGtnUI7ZO0qKBM3KeW8VKRtYGWZ9Lr/hr
Z+uW+RjcZeXCRNWqhwTp9HO9UPMVa85Wb2x5bw0NG651ZlWgmhRakDC+rPdRFh7j
wObwgW2rB9G/OlJlJ4I6NtqWwEh7yG7EFDoyzqzFvwBrjdQDIME5qZH7TB6m0Y1S
rtp2Od2BpmGrBn9T9fbBK0wbdDxx/Md906pyQhZ0bmLRNswzoOUQ9WcC3Bq+VvTv
Dw1PQCzRXSjkQ8S9U/48W7Ot9NmKLDx+XPORPQ9aIjpmZ0l5Zz+gLsDrHV/J3ANC
S5FTBS2Hj7ufFMRihpG3uEF0EIzBmD5aIcdg0NBJpUEmWywkrX+wlLb6pp2tYXUI
NvSE6KwlEAHGlgRW4l+nqzL5FGcQmI1vW6iAWa+DqRhN/ygpvimg6eHMEIPuJNd2
Wf/fiYhpI0aupUHG98ad6nsXxQCVmasaIXgC5rfTfN4fOB0bFKJm7Af0TbcEYpSw
QLDk3OjzB6F2E8WE9Cl6jRA3CmrDKvcRouqIVp31H4Jo91f8suGHGC6Te2lkdbhB
+1S5NvEToy3rkFWFJ/+L/72UOal69954sQ6lRfxl8WjSGKa+xMQTBmrXBO3/lNQa
FwPL/C/dSvzYAn83zmblCf5VowSNoLHjapGXgABWsYREYZjzhoDSVHib0BHY5OM6
zJTzYd0xJOHOKywN+PN891hA/XlJwHMvkFEegLlhZY36SQJbzJEqx5UqYLvVTm2M
fdxxpMUim3IkB8180Ijd82q0GJasDj67JY499BB3eWyJ06c8LDjOXlFoZ4E2CbCk
hpKEGIIZeXtL3Rrq0rbQ1hr0NfRP1DWdyq4414sS64WyvCnq5ZB9+HuupTBWdlnt
IbtJGd+jashsYVjo0zlJRJzpXEcjFLAEhUeh17evsnt1LKDpJfgqWeTwrx+v6V3+
NZJJ28G3efiJ0OkyDEZMZ/p2xWmqYZ09bTxWZ8bOh+Sjd1JxaFLa7oaSI+dvZYPX
2lhpHU60cYlw53u4FPZCsFIrvXMoLgjlB/L87jzdU3e8uhAI2/T0paacNQm5Kqib
aWCX8Y1LrqIoo95GzBk8ULfR3wZCw2bcBA940pwP+LYQH/TRiRXw4MH8xe9jS4Xd
9fSN4xREBtyR0o9zoKsVxQ8VNiMy/P/JiD07hIoBNK2HCaRTQUBABfx4BvvpAhS/
RN/6W2zWGNLYNh6/rZLmGcM3nPZNR62+VPsra0nq9cwcM6zJyQUhOgPln9ebTn+I
YIXtDzcjISEboSZfAiszo75MnPqsgLHyum5q0JmHZRBPkXUqBsbCYGFwfzCTYt7K
Hhj+2rIH+07pd5p/592znxgAtCxyy0JgqV8fob0UOlMMT06Ej1/hk9+CehloWQtO
7FmVycjw+PG86548PCSk9MyZlMS7oz6EzIWW3Bxm2VOh/XrcXX8/Fwb1ONHmyCs4
qazg51Sx3obZaP/PoWFwnKfa2vgDK0mPwsx1R1QEgR3iXgESH/L1+tLIUL787R0B
/hVW2nxv1Isx0uHXq0vLkEoBHTn9CZf1OgxyIjqOUgTKH6iSpWfm+/urdwPPEVCT
USoNFdXzO85KwnmWX3XpaWl9Da0UfwCSLK2GmxGqz0OF0xlpZ3sfyvo+FqJuuyMX
8M8r5b+rnf66v8GN4XNCQf/c7qr8C+rqrKx27KwqMwwpaJgKH5nCAvLHL5eF1Gka
hk8Gv6KvwcJMALdO0w0puFPgx1xIKvRJOBmgtOii1FfqbF+s8ul52UUSgAe4ivIB
q6aTkgQ7Dgfri95S+w1O1/VnurjLFHfxy4q+5rMiLL5hu9haZllFhBbuEDgA36JL
XSa/10GFIndxN9x2l0e55pYngjElO1Gxq0U9Qed7TffhrtPma/h0Vaa3NRY4n8FS
tp9qC7YXCXQKKKqXSHhLXrgPfEJwy5ionpWnXzH8xVJ68OAP8u+1qVUdEtQjNwlv
6vztZybapeNq0boZN3o9yWYBs7OQHNP9FEdUIkoIKEOJ2u6n4pEDorEZgK9Deu+S
2p40h51dvyxW8Dm4k2VfNolwdjzrQJI2zzH//Xdg+Ve74ZyeZNiDdyFFujdOT9kH
RxC1YHmO0eA1IiXbz9lwtPiio1ELRSg8qIcmu3OfpGsAli4RFBZy12slbUaUDXEq
9Xh7LZ8CO6hPQuqVxxHMxfNJ9FzLpXf6/P2oTPIe82jHlBgk2gJMUQj8ooxJg8mO
WaW5sJhIxfR0imbMJhX1kL/wvnrQ+Ce+Iq+BmWqzPAShP3jtkqFYr0FweEfJ4bGN
s6O0AS+lvAM4a722K45h4l8DW+u7a3PXWWEHDVykGF/6lkC4sGePvptotxLpORkI
okwQ8XXnbn2EINZCLawBQx3H6KUZy8VWBbvyVMj3XOisojYg5vC3S67dIQg1BoUr
naVPUWyUODYk/CUnmZcb2EJxNkGHXB/EOb94yM8cVzIg9Cmjgt3roloh4jMvqhRX
VxcEO/9tjpTjYAHXMz9w/G9aVu1svGUlZRqPP/7rBIIOEi/5xgWCkQv2QV7wy5Bu
WZerV7D2U8fHgtqyF0C9inYpCLjk/bDMc7BddSd9NwzU01vY1XE50Bl2iRxf2Gi9
+CI5wXc1eHRF4cDFTIS9iSxFqRTllmIfzoEnJ28dapFRHVtc9PZsxw2taqWbQN9X
zrgweJr0qdCiOsF5Cgxoyqq+3nba1/crnCn05O6idDTaEYQmJCBPKwtH/ywF5u89
w1dW0X1ROldig1PaSQK089urbmIG7BfyPBz9HXbVn7xOfcat1ZZhldr5CO+Kib+q
LPzOyR3Qm/F4jnVCwx1XXf3G/ox2lkzmAoqrkhrxAZykbQQeL2t7nAizs/AGlEEn
s8AdsavTnq+xqJbOkK405nMyhig18+JdksOTFay59FV3on+kfhCh1gkv4XeeuoBu
ofGfyFuQ8Q0TjcO7nXgl4jovHLR6jIuLM+tmn4reqC1wm20hMxoxCfg1wsqP5mKA
ujcVxDcKU2hU8fxtmt6mBGL17EoPMd1ZjlYtL5h4N5AWuyvWqIvupxP38cLWq9jf
kJgpL9UXng501hK/OWthWx0P+BkiHeiDkzwrWcbg9q09ufGR6AJx8AbLElwoC4H+
7MiwdSY/GxtZqehlUQhxFasIDif2B+u+BewyCwa8Vpn3tV5w99gesQbs8F+s00sM
j8O2FxyCNLdnkPnAbHqMD0xfJesMZeKUtgbCZSB1d0veZKFOSlj6OdFtoQiQgxy8
FODKNDtsWH1bPMgON2RChX81zAS3DCpof+iVniWUoIN7nVbX1w6yTr8v0b4ybqwi
iq5arRqNly+xxQ5nxhVX47dSoptTabpNBdRTn/RabYbP2jI9hZYR/XWbjQjESdz9
4MvvHZuC8pzRXKlcJqdrh2PNDzi1ctQI9KbTgsYvPgT4LUITSNyKD5YVsAX3SNCq
Znc4IBa59PwlaSMiOQCadYUQ06RZk6HPWQ46naHbzEsoNehCr3ZVVOv9sXS9RYsK
9xxmeGTCeQXckiFbZFrjGpgWYwq/IBpWFBL8dUMOay8JpmCk5B3tHwkQPr+ouc+y
4aVuMDU3JjN225/ONz1oAtZyd0N9/aTXN5Ug+BJn4TXaBqEszYVAG9dDHKRsGz/u
ikGmgt32fKajnp1d2XlpJd2KVp2slVn9tDbtuakzYJTqgE6wZbkgL5X/sJNDmbEF
KsQVMH/Q6Poqssd7u0G/TCu6MIBE12lgN9EpECpyOOkcYZnONMJrD5bT9Djv04PQ
Jm52tz2iVViYjOjQNAeuh5vWYWH5/UdaFoozV37noauobFoALxRSNZ4F8yk/Bru1
FLaKt0oYP/jJFburwZ2iCzHUIbFKwvLUJMHyrXEjeGi1R5G0ndSgNu0XNh73DyUm
24D0rFaOeE04+t59BLDFdi7hpfqGag5igN9fjeV+qb35HLMW8g53OYBfCIFBtVWi
O/SUDdoCQ5v6kt8L4a92HABoiGyHsi+a9KoA+Jxcl3Pbhddg1+JwapE+wRcykdCh
JVIbWL8QXwnSqBHRGQn5Uv0WpKyGBpSNckd9x2hxANariB4h5K0g4At3SldbE4H9
/QJW5o9OuuXG5l+BA7mJUKvC0fmIejyJi7Q4o3jYfb3MEpWCzCgMKdT3MhF517zz
RCW0Ws8nraTf7VYrCGV1H5/k/mO3BaD7MAsCgNaZ/8wxZn79lvSV2uN13eABtHYU
qYIl8DD4uJfA5jntvWJHvC5OqhCjMyi3gHyF2DTQIx4BrBdSX+GSVbZoiDOmxO8+
9vk4J4IUzRzTPU5Mo2G4VZtGGWJ+2qUUaSMZM3AzW/FdprsEFHTeIAJynojP5MIq
Ga0A0jBi/n3RejEbWKRMB+bm1dJjOy5+/NdVsIeF7wkXvJL9zbctOoKiO/gBPMkm
2AXqeyfthsXWYYTryxNtCDEysAIhCEy+R14H+2ui4X1XiPnrq9Jaw7cOtsLLYoqu
ZMgNYhyAwm1ZFbJeAfaSNc8ZSdi+tCvPkUeOg/pH90R7A6semCG2ahHl6iKZcpW3
4KR7FRs/8r1ciCphaSRZycD+pO76P8ii6DJFM6oZeBLlB3Yrx0JSDMwPxyW2wXH1
bdwqH3BnxTGX+mXRC7SacYJU8X1DSnuJ70XkqKiSE0Q4JKU2Pwgebq1mkkdV5MW6
IZPPo1Thbr0wUJfO4BK1xvv/NYOvP/IDtS6ofHSlNt+V1Wo/eHJ9dnopR+j+J09o
n5COhjb5PxXx/2WxoXOZuhOmVZ7Y8gXG0g3APd2uv8PF+mR5v5SlvidVaFERoDfa
brz1AxLG5Nbecf0NBAX6lcTUlcJzq17cjV2cCzVJEN1/Z/iUN38KcGO9V8Lx4mI/
/9lUMdp5JDLhYbLdEe0jSd7aG4wGvnnnkKhTFyw//8dFwXGWzsu9/2f3sQ+YVzrN
aH2o6RIuyP0UokKSwXAxlFYjnRloyvIj/GB6LyGKeC1Z2F8VqXtPTJibJf4zAvnx
FmM+37wTQ3ycTv0rcK+lHWof08A7FTOcXo3SSVUUnKbOY7KPDI604KRRxjXacL8g
3WDlhAZi19TP7YVStREo/wNJ3kQxXMVZhFH9wNrdlJol2YtAnsEFSQiuSJqzjrJH
TUuaWpo4m71cNA9OiTB8ciYVTbHK7FCxgvNZbHWoD1T7LGbNVSSlgHVF7SJWlzM4
G4LT9eUg7Mj1QfKD0d/JE+l4Tu6Zpr6Y0oNahmjBuSr2soktC03RtoLdq1qKJVgo
Y6JBnA0+to0CRW5w1Z/ThUV+xrpx4UZNlnWEFVwCZ3uI5NupcM0qFmuIPOErmqQA
kluHWnrZuCFz8lUfzWYU3jHqDnzFTtq9z9MOZj3MWJ5xUXzFJgVzIsRkAyBnD+Yu
+WJQwue1cAM/I5DzQXaUP6LcEuMO4ZSxayx80NuiCpew/SabxuXl4b7S4CmbhDP2
03/TOVIPKr/bcAJanL/6G/Id0pDzN44kPWk6aVjmFkCPZhBMeH7B0rOMBf5TN68i
ctxnk5NdbnUKThguSQVPSDTZyNXxrb82a528D8lLjEsC/xyhqxMvLme2Bx2qb0Uo
OLXkmpRqiyF3pUXY9pY5YaORGFmSqa6XNr1X89Jyi0A8OZbmJNUyou5kzu5BnrtZ
3kM8g78onSdRdlznBS0xe6VTjtLoQ9YxBvAtQQGHVm0v8lhdKYBxU7HqCrdey88c
C2zjieHZLsFNKyQJ1Ukbp6um2hbPefSaVc4die6JsKUtGwutTZ8PAACk4UXSaPC0
O0ITBFgTe5SyPYJOZ1CIIBx0vkUW/Sj8gKZi7qvanFS7mTxZ2I8HYSwZpkD234ON
vatfDex/XmQjQ0aI7nFJRiO5TpV0Fo4bj4ERVJYPfTXhbXCAx07fv1IZmMzNmyfE
CTGaqB3j8YbCqx5Di6DFCJenlssErXgJ5QFl5PJVqBrh25Xbb1wuLHpke10ysXYz
CZJ8lso7VX/FBd/xqp5dOU7aYb+9qJsIrEJ/ZE5MHHzdB+k7FyzlKH9xmmFylbB8
7EXPf3NVO9cNnE752dhnkVIIpMSt+HDKTA752LLD9jYIfrer1vud/Tx5xWVvl/PL
7CrU8vD5mHPWkDHlitQ2ePR6PCEN7pAGIZ1gTEaYMv7KQLBtlPqGDPG5JTTSYdwf
QPdr56lk3mrYb2UJjGqTzsqAHojmEDj8pRATNUQSM/AdxygWjTvnxbQtJLgoIW+g
uO/fnwyOffva68eiirdGbVBzfbP/xhegYu0xSmMieGtBH0qgnzQtQbGJXGMagMUo
xTXqY1n5LDELNU1Hx3QfC2Eo982ZBf3tOz+/YBu30y+xjT5suAGzoH9o7jreouQc
Psjn+VFWQefMPRnLg+qvJ6JBYSO86eLQbNcX+Z9dYXwQix/Xvqhc5530xXu+D5O9
WeA0WRPpo7zmAJW44X+gRAdNqfLB4pHVwDcC/EaBvPbJcD1myR38IRU8x5C5z5by
BKktyJ2R53XIKyhmICBH4IUPxydb41m6Oo3MkW8GfQh2+rlqscpJHHueORSDueQ5
9gqdLnU2mNAOWjpU48PAPdSCB62A3Z80dj2iJ0Ab5OCqXhGJ3RFPvsN8156AXl5t
2u3bkaK18MPGDvd1eZh06Z/Y65BmxGsj+IXexFJQvMjb8tlS3E8G3umCjdPddomP
Oa6RtLTwfxEiSsX4H7sdB+zmZV7NQkSLDHZ09sbxVBaybkl8CEsbHl0SqIzwuIFw
3ybMh1hp6Ct5lJ7cIEFT7b1jDMutB+d3zaF0RGPCv5EEZhExot1NusaNz/4mVrkL
srEietiroqOA+JNKGdsyBbKWP1WYmQXelGr7LiDaCwBNXXpQ6PdtyRf/XdLaA2y7
g1YoNMY9qZdK1YYGWZgtGeU2VgIwaHmbaEFBFC00lLZpULGHkaQVIqEjOus74zoc
YK5+INbXUK6wCOsb1r8XGreGovlfE1Zo62lgkmKVN7H3VNhZuCHsVSz24zSbM+6h
0WFw26twrt6NF4GNBSaJ8Ll9NSXQiArTOFC+L449OcAE7ahkZ3uQr+NIS1hGhm65
Wo2Ae9l9T/i/bMwjJeaZJyOeRW3IlEbSkcLTmewDjHKzj5oQ2YrqOB+gIxNj4ofZ
hAeWXVgtkriXMs3VhiJza+lmHd3lxDwB26fXM4nJu8sFF0l7hxWHgVSWMe7/S/Tt
Mz6zbC70B8qxR/oT8f+eVFzqrl+mNVit4arlhcHgcAqO8ffk8bzKDepuBYSVtb4K
mDbhNokSFF+UbsabAtyZCJyb3ByZf5FONeAuTltCuFICQsYQDeZptYI1Dy2P2kDy
D0pCdB7ZI/AxXxpvMcH/UgcZac7nwK1xlHenVm9FxFaAURp9OA3FB2ry/WZUmiW2
3PakaBVa7NU42chUODpAD0MScueXMRNqmUm3i2G95F2BVZ0F+xEuqTVrsVK03Ufx
xe3GFPa6Wy2W/m9qhB08Dwz7hJBRrXstOhf8aFbj3zOj5RJNac26l5QmPZ7sMEl2
lGMgeGHTloPn12ccjwQbOz9vA/+wFDcrcf38LfZRM6a06DkZwkWB86Xu5CepM0gA
wUC7cL5YdWSjhtThaz1kOb2t4AyW8CwNQ5+wFk/b2Y2VXblwHjdsNH/og2AlsJV3
IHNHjCA5zKz8z+/bPganZ9a2Hft2/cSHKJbdB/RRt1Z+RtIJ3hIZlYXWZTcueVqq
p66MPkWiSH31VmqAFPgpaLwzO9ojvQs5ycJy5WSxpF5TuMMlJKoR7z/lMlEbeSeF
Bb/HH2Q9fWG/68+IArw4hs/uikeTZnRpWYqpSwz6AchaW/UKdqy8oXp7ZxxiizWc
2PiHNlOEfgyeU9t+4KGLdnOeRhKf9AgCTURv/zO017DmO7xOjeQbsaYGktkkQqt0
YmLtZv7BL/HwljpZL6PTYFubUHjJbb7pNuwrAL/Yt626KeETrHp5XbePu0HotmRP
pEz86XWoljZdTQItji/bKTDPR1qOK3Q1gySlSgrHMtr8e/DbJWbjOCXDBBUghyIb
II/xUT0ksYxzcccm5Fy4kV9iVRiPPxo9EP8inPqKz0o4+JcfUWna7fcE5rsh0jsX
YpaGCf7RKXApwSMP7hxCfbEPNdp3Hh7WNFMMHHKBY88Opn2YPRsZSpHh2gdDx4gT
mVvNUP53iQGAXpxlvUEkUbYj7A8cuk/GR9p9xbaJNx8XLPBgmjO7dLB391BJFv5O
0akPwRV32zf+jF8tegvzvxz1ZIUhCPDgbsy0zKH57aYIXlZyUCm4ZUKUOMkiyt9v
M1dqga50Um/njt3onzCnLLNSDnRDZkRRA6hkM8gq3DN6GA/DgxK+m+sXLHm8RKpC
3bJkwYFSqy1yiLTN7TmEfurwXIaHVtLq2rLrYXhFhpJTM5zfJk5v27Ss2QH6C3IH
MUgMO/0WdDo24J/kPoMGf1tlIz8jlSkxouhEMjni4iWKkXL/aj/xs7wZ87oxy+To
6bZ5AEtcQPuNkYedgdsiY5/8i/nYilqOvf1r3sfOTazM3pNDbggsLwu/RjqDtG7P
9h2nXALGT7t5BWxJRo5ybgCuE8hWs4tiFT6fsKurYYo3nqKeWXwdoE1VaUUWnue4
MUaSbiDLzzeEa4ONG7lIwrLjDEwjcD46Wli5MWh0VOp32/8M1hUuR3Ii9x0dzyLu
w4q24aErOnKfl/4XKBpux0/YaW90i50is27H+VBV59jaV9UDtmPptyQaJYKVQU8s
mOPJRgM09IEi+l5w0jV6PuFJyV9ys1AuG+tCi3/9ajHW9p5BK3aGPXWe0EyuAyX1
bP8jJjO2OxEYOSDJDkRBQj9IXYM9V4LrsihqDG7X/Ionj+zsGTcX9qmdzyrYDXqc
GznDHiCujrsiLWmnuH3RTDvDndQHblc4m5wv8FfCuae7QB6V3SAaGwKVSpecX6+S
s4F5CDgFFje2EpS9PCB4hqzVIPl1UmRsgBRB9ykTEJP6Iwq7HXCqcK7gtTRWjkhC
hCeIvtnmFxAl7DODos5jYdMiurS9/llIVzARr9OUkOOT9tdS2UAmkpf4jhwj1EWw
X7Dxzl3En/SS6TYLcJbSGZpcHfd86DhhnxE4Z+76jtNR5bV7dWWTXMCmAoJ5fL1K
2OqYAbq8gvHgo3/DPkbzlQRPmvL47oyipT6A4D/flUXjQ3Da53mn5jc+SxlLH2Jq
m5SsBJ2aj9EeVtMId64b6+lmIW6mOOAXi4ocURqCeg4SSsak/CH7BJmQ0HwUHAmT
B9tWl6vAI9yTUVD1ObjrPBaBjaw7MkRaa6geOoZkCxNlRTig1JUKHshtY/aNWJwQ
CVhr8F6DRDLaKdWb0sVcl4B+GTOyMrMpHDMBWT3MrcJABi+Ui+OY+HhKDDJvg9IV
kBCoXNN8ZNZ+/k3H+6eSYAo+j/QX0z5imR6IqJW89sYIgHc7LSeeG7L2QBtPaFCW
fYvVDto+quJcZmuuvO2b+ewcZsPVVtcpeqDo9ENqY5Y4e+UEFl5Jold2g7nW0Vvv
OsOKjXhT7uUsRdnueN3pTWSP77uchPTbHahDJpuk7l/RpZP/7tLIDqIQn8xhm6NK
zic7hVmoiHFvh8Q8fXJdgzqctFmh15u1eqD2sQW7+U3w45yxBHaI/fgNsWz/JqzU
c67omlY3J9dTFCzNykxCCGfGNJ5AaHW7IbyeXnhB/B6pHKsOi2qKmd3c1VOzAEfl
YnCzN+gZ66N1EgzM95dJr8GBg+zVvN5sifsymRCQJgsPBttAIqFr6ZL/6ocu0LJl
3vY8Hi/gSk0L54s0b86FePSgJMSgp9bPa8G6ckEtGPYcLaKWqb1T3umq2gZahbqX
L0LFFMejVZ8+A5o+Vyqh1/OtLhk1k9kAEckXb997lmX/WVkNq1lw/LATIsECoS2V
+o29jBYN3ccSCW16957s8jV/INAQbyQDaJ5VEjZGYNQ4S7heRCYplogFNWYwyQwP
b7iZFxP4BSUL6Os3msZYP0BQv0WVnaWIR5gV2EZqxR1fRJVio27dknnld6ciSeDf
IjsqSGd+w8PAg6l6M+vYzM4C3h9bJKIpIa1kI+bbqQLil4BNG6qh+eQmjVM60Fo0
RKtX5yP2ueaBYv4W8f67QskhbYWuApPiWrUJ38+Xb6sqq60yW3mtcJYWdg81NT9w
3ZUMra8AOrjCHcQcQkKy0nS2b+idxw29TYU5SQEfNSwJEC2ziQQ2FNgN40Y9xj5I
OiTyT2negx0/MBNbW0PYyZbzZU3zHzLKRUcTfqm+FMmuev/pIEJyADezTk1g5YEI
MIOSMxdhCbT7Dl+dPJvojJrfTHlUaQz/m1ICcd9xqgzF39nGTSqFO3sh77YDa52F
/NrR2e5b+U5wfNkYBPBUUSeyIbBYs4aRpuzgPXfp3cnx61HtyqH1K9iLbeFuU/SB
EoPEyka8caujSpsLDsLnQLxCogsHcYSM4YTOOIOPHcjXZe7jnlpqMP2onbOpdD1v
fuJpAp9MFvmnaM0EvaXI0OX0qGtu20JyQckRmsoLzUsa5gdcB2X4TIiXBCR+RswO
FVdEPtl0zsOUKg6XIpA71TI/g2PS4fGQ55FRugr+LecJrJZOXjNOmDa9iBkJEBzQ
nKyEzccaQCECpFmv2K7haPfkXSc3UdrjE2Fh5JQOEo+/KPVab1Xeb6RNySFbv5RC
AaE6yYXi1zHYV8pNePfpANHI69kCV77jEwhMVx5W1pFz0SibJqV+zyKuIEjCFA6V
X03WeMn/NgvCEZuw76n7QNT8BAbf6ukDj3iLDIs3U0F+E76l6ZtAJ+0R8wKw+lex
n+MxTyvTFeQNWt7q0yav2gEoUnIT3K0bz5if13jRAPpqOCo0L7+4TZgYcVsc2RFm
u9to1vapfLYXHKkjH9hFmZUdFuEHbB33lPWMh/3hQxbBl5ZVPB9HplSgoy4jKLm3
qNSrKz8Ek443+kZaf6rKFT2P+XTVz6O52A7Oys0JF4mx4jCOZQmGe1sF9ZWpU7g7
dGeqCCM3hU588Ieob5wrL5Fsea6FJ4XVevCqIxtRQtkdaHpIzuFdzu4QaxMqf1Mx
dX91pEWCKsutw4V3IyBDYNAFWUXf3pO+B6VmvwPBnpEVWZqHKKq9GFy+6H82bu0y
aBeFLLc2PPVTRqNtwWhX34fTiP6aoIX4LbLktJXKUp5t3UTmhpWAmjvJf3nUlHoo
Qy4eQ9DRBEIbzw15tCNxPfr2QEWWwyAa8ubxIL1EF8lJGOmWK1IteObSkZhsPRzs
4BgiF+Z7Rkf/YEi3NogUgK48Vbco9Q02MIuMvav02lXeWhuZ09TikxAzos1zowRv
TTnlvbf4jjP7JMmsE/X6QOAtsJVyi4fYgdrSDmdVdBf7YCj+ZYvuf1IV+xyL5E9G
5EJGV13BfVSrhVx0dfkSZ/tAEvvBoAglniZcSo/QlbT2JzUg27ujlFh0Yx0nblNl
RFfl4LNSxjT0THrucoD7AGS/XE7ghEw+XH1w/D1zEUjwAhrQxjmgW8brXfZBz8We
qwOhPvFjn/TZFgjpPbvlxqMhV3SUJdmla7lJm5AnhUjFFTtXSJVofsViqlTSnBng
3U/izT+VQYBMJMzCtzdPMAregWa2U3VVfr7p70Wg0rxv2kVk08UZ/2vE5qcS1LoD
MIiSpShn4lW9NpDn4K6dgrmtqQzFwTKjP4fL0nJaEVmi/0+PcFDTYU+KP50XaF1j
0T5wXoVXYvHOxvBpYSzSCBNnjDZ1AAtyEtKYc/h2rIVGtrUWYVesmrPGY4gHFY8d
h3x5TW11tQ1GUn5DklUI/SBRGxXHoHjI+q5UJ5D8ck5rJ6YsSdXLx+T0kgtJpi7w
Cojrq/Vvl+AsSEyk8qkslbXyizzXVhWpPNpWTOq5O4N18Eir1Vhf3PneL8CwnPK9
9qi8YIVGFc16KG4U9Z5ALvWvieDkmUJpY0ubjqRyaqJ5l159XABTV0raYb0As4F9
F5BTgQCGdaBZ7vB2uOyTj/W/ue0IGftNpbUPHe2kvZjHuL1MjlvmHMgxz8O55S26
lWdRfflDpUrIQiHu8x1cx08DsWnyxuT2aBEAHYIT1Vi5Gb4RqaCtduUDv63JHHCp
Dm0IObC2QgsaxuCPlhiLH5Nl3+aAeuoXnVgXqbuck26DK0g4rMBQWdDJQt5ec3Tr
DdLy+oWrddtR/6z4R6sM/3t3IDR2NXQeX5zFDOCQMCaHP8uZJpbPvifxpUaaYlBI
5BHRQKKya+y8XcwpGamnKqvo0p/CKr/ZXTOfSy6ELFfDoKVgm4UpqnODUm4/EDsD
DuL/fGhs265wu73d4nWFV9Q+QllbkFKW4hA04o7j1I3t5wi9QhOHHf95EZYeYjjA
O6aEocOW3peZDLjuD5S9rEgRx/rm549ry0PoRtY6qNL8kFi8fadL1oidbEtM97KC
1poQioZ03OGF6mjPcQyboycTavBYffBB7W8QE8wnIUP8U16EN4TXW/rxLqjWSq+o
uDyrp8SVFri5akdUxLR5xW702avxljM0AtUAOPj1KEOTNQs6Kc78eYGm9ueGZDfx
hXmyPgEj4KCLgR8FsY6gpSUSjIjrPxepKVnAEe43DtXcDtOq95bCmekfmywJx5VB
Fvhvf3url4fUC66r2F8BD7joml45myb6fjpAN1dBaLDpoSglDeKWHx7hWRzG/jM3
xkNKILRJzSl3lF2NymtvOLKiUVoMARBV/1BkBIHWsKKkJZJMbmYo1kcgir3Pq5HW
Ut3yGK4316dSlCm0zvPyJPrt68vPx5CnG6IJfKry5afqhultp1lpXc3Tzw9ZqtA8
Cts18ZlfVBmGWVNVSHfukoQHHoHjFhhhifu0/UOnK7ZgVTaO7eJRwvMQdErk13zV
xacIBMfDK4O7pQN6cmCTy/TKUaH/Eb8kFmp0n/ilO52HRoS+9hW4D3DRMIpon+9P
mGH9AbL3JU0JydtfQhvwg2ZKDMD6f+KTEKiPLwadA3ayMN8dX8Gmk3o/tkc+Yo5z
YHQTu9oCSw6xcQaDyQFh44qmRbR1oxKWB1Ggo91Wy0A/svg89Mo4ydk1nO/GmfZo
yvsBESSjFgtNAMajR21JxklVheQdPKzIUQ6xKqL0XsH4MhCfAlUGYmlKLOkORIqk
r+CIJwxfAqdtTVarr8Fev3sUezdzKF6tOUYdbgX7SI38L5QPjsrQWlwGh6SPSOhs
XD6n3ws5MZNSLC1W5PQkeUrkyJXyNtC+GSFyrKzp/ZQxnUZMmBRzRatzH+VEga/r
y1GlXAxxdb3DbUUE3gUGyPEciEA/3TL2Qonb3EZOGMudYOaBq8m1xhHTFtotUcO3
9c+DhQMf7jvI/sn+Y84PaD78/2mH1Odht5ePuG71dhXYwkgR6/yjRRJIjYno87u2
NTVtWZF7V7kddTpQZJf8Xo0lRhjSYXeLw6Ww8rAxSeW9dBTgFRMdUM6SupJkxX8W
PZLwhRj9b/x7WcmSHPC9ztKBYEApP+/zEiTf6OVlFLsPP/O8naP0HD9W8r6UxItX
+Oc1mf0SJpBACGhOBa3FoEdHY/hErw9zMUEiOAw+i0IFr+CvapH4TRQy5WG6cD69
QYeD7b7XdhlgugibQfi1VReA3fOlUKqLU8YKz5MR/IpMJDr0lecBaX0TWkdJ/GXJ
Tdm3fIJqFnB0XTI0f8xd51a6ODTGGk/gZ6U4dO7ZIeih6gR3x23MoFtj0anICzFX
6dU7Wf6q+3M1XmlcVJUGEQdKKGic8VSU+q0ZV91LSr1/deT+rZJAljzgM0ZCUzdH
QIRUskumccbCLr/lWhMC0acJfWJ7l9rR7kU1+La/bI+G+/OeULOCop2vLFcb2J+5
OS3NHR2cEX0sJ1L8kqFK4bGpuy31kLfKz2qN9CZQxcRDJghRjlNcEpT+szpTCgvZ
QkDdnCrKLSM6gE4lU0cG7cLnoWx78F00PQXY898ksUu7V8MEoi3v9WDCev1XFKug
UK1Ele0rYsSIKdTticD7W9D2qBqZ5xiyJoE+vO7VomoNU47iNsGqM5l/1mpCclWI
6iIn7ru2M8FmdowWx9dQjvk7hKoDAun6OWKp5g8L71CVw8BQYdlSJ4RRn/i6pAPK
1WGqv5G01gZij2I3nTA27o2YqUqB2cbPhVkieIQ1WM3opTlwW9KpN3luhWFajO9j
yNuf82bLj5RUV3ySCKTUM9GPVR9jJX3R+VHJ3aCWbz5tL8vgWul0GRkHKS1aFt5p
FxjCfx4izI/fOSemPGxx4J4quoFDTU8XxhBr5tkQQKFZ2nXMLjiwaEJH8R422D7J
g99QDuWV3gmHRkQK/F+/ZTsSZIF23ZndNEK3wYZbdr+pLCM+18K9JtPjCSuyuS/R
/JfClOSK4PfouapHNh5avKpDpIJQHon3o7jbfcKA6xP03n26OAT48trt2wlDo/GC
jlo7fY02SbjmT38Q+vO0KnTHwRlXY/xjC1wWWcLTQgKvcNVGkEv3C/dD8ovWPq/4
aEzcqHtvyUp/A43ZhWPvNMYGYPHmU1k1q2huxVzZtAIO1Rt3cfm3Q7ALeji/BQnW
yVXxogGmToJcoYNzwdq3/Yy8uqn12rScMpaM+qZL+O2QuKsaKd5nPl3HAiQ1WiZN
eIBStYz9YyZ8lNDQmCxfEiribce9RfUW71/U5Slo3HDJKAgwv+XTUPzMiyo8mV73
n7R1Uu5c7lXxQSBm5uAm5Gb0f6fz1rIUC6EbESaY2tO847oGOrsoYDR+vOW1UpLU
1U6APWZy+XFXlmlp/bWu08ul9e5WWHBN0MSKw+AGsH1rfgmrJa+32bEKHbv2K8er
t+4a7OkYUCUH5CgH8xN3iChpa+trXhyssvqtMz5bfEN32YIlh4NWoCoMWSUidK4q
ylScdWekRcxtYR7qLZBgZExSu82Q5vAcQKot/bOhYaxsf/WYo8YpuV12HZe/vWhl
73eOB8njcF9lENsZV9uDcI2KQZg9ISuvhFHLXA3KykPnWM6DflS7+gSUY3wiJLwM
lTTgO/AXllkLNSJgCKW4rPFJ6VAIVIMRCocaNFdVuJvv178gPDnmsWFvJP9yd03X
FazN+4e8P2jObt452cSw/Cb6sJefJQbhstTllSvqdRmBZcgQPeaXEpkXIYtI9R5n
emRMgxwKRM8NPUf//IXMVcS7v6j6vX8ATiy95UmdN2auOfK2/4Dr8iBBWNqPxAW8
3BR8PeDB9MMvFN0L3wfeJZkzXA3SihHXVyDgfSqemqCb3MANcEOBLkPrvKxhsw/p
OPDGbG8vRKF/OSdB2n7Qhqt3cT9w05e3BzfSoaI6DQDRqoW7C2pQN3Usr3Ar3arS
6eFBOIfPnItyeJ6IY+ioVazJT0b6dy+ppkLEYeokOwhzyacQVWjUUgtASwgAb4Q9
xPxGinj9YFB4FGj7BQAeGB4DcO0XYndv+8gS/fylDCmcNkPSmyIhFGBFcbjQCR6h
n13f5ZD05zvUcTBzHWTHFWDMstArY/h/Qge1X2FDrzyXH9awAUz83cNAtt4CJg6T
Wlr5sie2d1ybRCeVBzC7vnwCrFvVs5iQ2079xjU86C+ktHZSn0Gl7jLe7JqY2GSz
pNrkR4oS0sBELOm11xJGQPLvSa8c02l7Xd0js5HDMAnHl8Hxc7uRV1w5tF8WNB2t
5s3Zvsn8qFDf6/WLJbcZDNjW1TrcsQAOOlbdf/mt+KqmkRIMZWJL9hnMp7Cfi0Jt
fJLjKUwB1ZRqFssxM/XMYeutA0Rydr3PUq43FxlKvqkFkmg8xghzNx1a5tHg3SPA
UTd5galSw3a7ZhPkky3+M6h/7tvrtslDfhYS97xMmG37g0PIVFRwYGKWHw8ag9WK
9SnQRYAbwME7574nyKkDp4O8T4LqUvOcJINOxkk0Gh2s/Xrk7fUuXeBDZgp7G370
nq16A23Ci01yZZ78PkdgVWGGmwtNlWX7sH8VWH2YhjJucHXg2M2Q5ZqxDiZFYHTU
xu3B5c8dEljCpEdpDOloXn67oyd8HN23Nzi5GM+FbU1T59xD/jNKfXkmaP2K6kbE
qA879kPvoPFbDgoLY3Hi2Zzum1R8EHLpXL+F+tYvROPGUgAMPB/rkRVF/YaVwLjj
+S/JGpcBfqfe/gl+NKbq0+ZntZOt1W9HKkFkeh7EWOVK1G5NWvR9Uvc1Gr/BlLyb
kmljyR6T2UfrIA6CjNpm+opnx1OjQxb318+7GqgWabito7BkC3wFTj4m3NkMiV3z
j4Wg5VkfQAhtKc/GgzWHTPWzfPKlC9//t7QNNd7CYfo9nsoxVyF3wSlhtktnz7Es
og4X6gii5zMps5lqey29GlsiuGG8tCO9BSXVujlyChff+BzbtknFk0PXiucoT93W
wmD7dboNLQbmbus88NwXN281lfLX0P2GLYTO3FF8woraO5MF9Xzkh6A9qBqPquPt
LXeSfKjua0L1yEv/qv45VNN8Q7YdgH95Jb45osbiX+uVyiGkGHmFpMXeoEiSfWp+
/ECDrEr/HsIhPnZS3VxjaF7T3dgKtFm0KBOFWSZo/6K/s4aXqgw5JW2G1jYg8fGy
6Q6lKRAunTpOkriLo2+y51TghVLD1wmMB/PwPG+tl6jNcNeoKB8tRCdyGrcrRxlM
JL6jPMqsTnYKMQiLWZwr2/5vq5KdiflMnPrTaQuVSbclaao9GGIe5oyp7A0egdcX
aJhCBeCWtz2YGP54bo93mWG0Naqz2I6YM16IIcDoml6hSa5fZgukS60BXfwBx55e
YEmmZvCEmtmzjjTs9xwWN5JpesLgQUnzdaEQu2Rf6YF0AW0oC2rwunYqeYs5kWWB
dJnHtylH3N0pN30ilMN80gR9AHWjyU6buxGO4U8OOHApXHowN/+HUcqIFIiZ1jz2
5qAmyZ03GIbRwcP7bg9uXmQLu7R5GHvUhDqweUT4Zz6hSgIG+0yprXIbVeDgnxD5
MyALuPkU3O8rovmGEWAxXC+yrbsKl4qarjZZMjQyBzcI3RNtBgsn+Rma9NPbWCFf
5IWAbj8DZGS0KQNesrQo+cEEpbWu7ToH07MJMOZX75vhPi7xzzTS8x/ZdeTwKFrj
v34vQ4/KbpAczJf6n252dxtxkEqohYtGtax333JHDFZxW1WxHO/b+ehwl5QtFqLd
WjumyrJeZbHysJlKsMfU5oz6wAhYz/iZz5ayl8TjQAlRv3qgKnOlkLgKKrvoUSrT
dhWiTUb0wY04fOI6rlwV3Rbxv1q7A6KZHTqUI0L45SvKPKTUagZ63haeRM/m4SE9
klH4/fGU+SH0XF5FyU2MQlUgperuxNIfd4LJmgZHwdPkT0F9FK6CZ+KMXLdXlVej
QBkYD+WpQXn8EpAEPp1IyZFpjfeQno9kfU7wYKaKwGw7AnXDyQCkn+XKqET+vDtR
OC3Wevep8m4ZMgZYjZSSpn6ar1GzjLcpokWudu2EgqO7vcq6gUV2wkR/ulUvmOuq
hK/V8kDR5CmD39X3y3YyKmPCO2QJfQcSbz0XtJi0CrW2hknz3OqlcylHneeDI12V
RtGT4ebmuqU/egEcN1gJk426I2ADbiU7//J/hMaTykhSDwjpd650vVA49s0lttbs
Qx1wSnRrr/OMEoLaMPCCB/sEiYlZpp+X7fav4HAPFBLNjfMwg5lAufbcEu5m4Cc3
u6R1JToCE08wsW+i6MDmM1R1hPaEqgWaV8FAK+z1XKrx7EgIoPHSHk5riFMf8GgG
mA3wjoB786BXqOW43BnmlOIUVybHKhLptlbS2BNgxmsgNIFNRYYMpB3H/+e/pAFB
7shZ1j/blzr0tnOtxR5myZPC9vZOlpYP5rmAxlT98PDUW5pcfjqoWQrXkv7g+LKP
29XJgEGFajxJqkz3XarFdP1I/mLvKlqE/AHKJ+ZK0zN8Rb1f1ktNz8ztBJNcuWBv
SwrxRcyp2foiE8S8MXFqKtVOuSotESLkII/RYkKz0cQ6f/0Fy2p4zksQ4bDSkT3e
T2YKWfQyoJg5SNv4/P+gO9JgN6hVudtuHYfQ6sv4wfOMuXg9+gWq8vTfEUrS5tqm
GexrXMvwyzQjj9kyFeYOTDKLMtmMQtKUA8uzJSovI/KpKkzsecC8iIWzdGCtull0
UCfio6LY3ax+JYglxabmN1fXydLiGZ2Je2isR/eIMFhTpo9k9o3+6aQid7Nc2qq6
p+pn5bl351S68AIToPvVSe2oqzHck3Zwv6i+dWp499y3ky5yLG/nN61ErW3iU/CH
EoQ8ljayZPEeCYNr2fI9d6uhA04bBaTjhOHf6HCHqQOPaATb8lAEjmK7SjO5QODt
/MvN1P7P1FiTdX346Ci8qZaRbl8gWBobdcQHs5Ggs6GK4WrNDnvH8pgB+3ACXtrg
W6Z9l0DALs5yqzIP3HBpdsIeOh284uQP+Yry1DNj/QzTo0qBxZsHYXxqghqBcVVv
xFVprtlC+D4Xse6Jip41/tQvRL+84O2IteOCcw1bIxreAOzitKZXaSN1LJ4Ns533
NYb1jIRe9uGBLcmEWbvrVWLWH79lqYb0YQeSHv6AjQPB/j9O9PjgRyZfzBGXnYWN
mnD3m8OkC9cW2cKaj0sysnpUvRE2KCacMYmIqfUvwcGPGuJ+eY3TyKkOQstOiyjs
/sZZUfjhgi/PwtiOr+yJdqpbs1QnS1bwTWJBU2sCXg2KRVnTkjasuQ0Ul1R1MaZr
dndMu7Ad75pbqjlDn05JoorFhpSXvqld5zDeHLHCc691YoLt5Susi2lBYUfPOc/+
66KXAlV22/oagG3uS+Th9WvjwcSI7VdxSj2JPfe4a/tDbyXuqU1zkbHIXIPIE4YR
SEAFFFqjGnH99YTllTMnk7HK0SA9NqqANGdHphLkg0bEmKY1c96WfiQHpw9ylgiW
mZDKd1E95EbLD52OhcN/c/r2Rq4EWQ1uy24MejkO7S0nNCLbSu79Lnw0RLUXwxPv
5+oXXlIAV3CLL4avQMCPmfW3Y9C4lg1CvDqZWAbh40jdNsvlJVZZona8t6OJTP6C
xdJtgwHtqzyOkWuZV4ZLwNdZnAkdInV+o+/TCLlyXt7ayc3rOpZx2wf2hR7dZOn5
n70E2k6PwUYYinQSAcOGEKI9J1W/CPCC+cRkIWZDC/dznAA0JRlIox8wRxO59wip
pN3FkNOSw6XLKHGovuBQBVlXWoZnU5Syo00JCUyOysx9j1/v74ngTMMEgpX48zx2
2X4d9h6WJ4LAeebxGxoF/3KIC5Uc6VC74ooKv5QDGVpITBYJKZonjsX9xs4zvLuy
DS0hkVw1EzVSecp/DibhJSThVRzPM2YfMYIN7KrEcvWZuGY4aZ9EMkKOwRwr+ptb
fxNP1ohqc9D5yj61wTZseqTpFJoDPnTpCuwfwZwCqyt9dvmy4mjb+sb7dWJ8CCXT
4Hr7VV26IA4iVglM5rclIkir19S3a0/pA0pDKR+ObRAVv7RKLr/0MzKC7UOD0qkL
/gDixUkJm/Y0IW0KmrfnOGjBhCjRsKO9F0tHALDsJGez33z4AddCZvMTxWFu+DMh
lwiU6KAQu7ETet0vShcTwoLFwZfxo4GzI0v4fPGV8fag8VqegtVn0w9ULT7o2FiK
3zmn5DFgrYZEri4b/wbyAT1GFeigAVkGVfO8gW16vyb/TLnJCBCZlZVOBZSaCI3q
9wE3pULQdao3sPLtMu2nvU6CBIQHG9EnNXxVH0gBnQOTEiMVB1KQ3800OMaN00RR
nE2inOEf0IqqunRXFXWNXH9elX7kTGji4iTjcW/7mqXeLp9lxcnVqqz9fW9s4JU7
kkC5cfuQ6trfe3OArQ7XwhFQj9ZToIoVgs1fpXOdKTXplmSkn8E3cMCJy8cOXe4Z
Fr19eJAgjHT0ulD6TzbGsv2QLbsU/BRjH5y65OfQaYXGe8UWcMasVZ7aCe4VJa+e
sGMzupWUHRlzzbTknZko92k26bjPoDQRHRWhZrgU5skaDGNxKzVYUhDBXiW7RxBT
njX1IEUH2HaJKFkVnq19KRI9NkRqCXy+EFJhaMtzdaBlmIFQ1C6wT1oY40ftgYkW
fmxh/KBpwagMq7cl0uJpVznr8kvkfnfO/g1O+i782SA6MekpfnmpyMdfiSXa3g6f
RbHD2hFFiIUKPTvL1yjiaeAm37tdpSB7+Xojl5pLBUgjVSh8rzAGV4EHrqw75XTI
fpsocIZWnf/c8LhC6AMgAJC+scrDNau7mwfsK+SmyTag6w0wL4zwvqp2it8ec0Ak
x9hr4VaWfyviMqVzbApPWdoRBoNXAuQulFMSHk1R+pyJj00RRG7xHV1ICm/czNhd
6P9dEOUQZ6L/yER428NohwjivqkIz8d0/DqQz03oS58RkrfJ7vKSpnH5pEuRWp56
Dd3HMd9p0j0MTtlkvu9iMq0QM1yeWPbDeypeYVov7s3bzW3aBko8QcOpk/WHybIE
sd9AUH7YA3Rj+d8J3aeuyQe93ROrKR9vpBU4lQdJ8fBR8o4Ow7fLPs+JkVCDGoRJ
F/ufk79Tk9nfd+cLc+8gXhcx4AnfcAvJTwUbcPmrPXFu3S7mSM+WyBZNSOvsiUy+
gNHuUfAg/QxXqHiyeix9rav4c9G7/FXNZ7Qn3mRWUyztPUJFR6ImS6HW5qaovsdW
2UcQ0jmVPRHSdxIOHMkpp/KKR1qmhngyvAEzev04zY2R3vldUMPJAoIZEtlRsjcU
rr1Hfj33WVK3p0uPih4kXyBwA1S1dJF5NVpdOvGmTCmioNUZRm18DDcShA2icq3A
SvBSC4Uv/sjST4RqJlA/NCM99Zm25gxwvDjwAH5Vi5evnsKZ7N67uEFLEQ7Ayugt
kjbVK4MWrr0k74vomMlDmKR6yCFTBliB8h9OBqbN4WSnplO941hlNU7bfzt/9XQY
3Ns5uGrYe8Ttf2nV0+duzs11FcCW3T0OZtIA4EgOIYPNPo4tciPsjEPlLLCU6ET0
4Jorgv/vcDFN0sHqOK3Gn2tFwJpEZXdoovEDCbtpC67NfLvEL6UjgjQ2cXDPNFkD
dJukknFyxNDGWbn+9qg59qq/i+a0Zjy+PqB41al8/65UzeIpQXNztFmzXVgrCLt2
7ayLz6wGGnH3Rwnp+FNjZSv3TIYTENjXi+JasLM6pGMtxwbiYRW21kTItvEybodP
9My8MrlHUCapJJD1PGjKDwOarxBB1N+5wwDa3aDSjSfLtdfwgZs7+ZaFYUoTdt0U
dm3vhNtxOZVdiwAac/CjbmaEeeg7lh2RlnG6CCip7hfwWS623DlHfBYvLuZMxqZB
1e6S9TrLqIPLkLw1qvTr/yfzJGX3cq0dYssCTwjFLDeHoZI5CIZJwtVprMnUivuN
/thxwvP8e9P9DHNWg3BINg/Q6+NGWzP60dtm7kBXwVVZvJTi018S8w784wpAsmhP
Fk/0PaF4pE8XMrY5nCb3E1RIlocssTLnouVx3hMX9CFaH0N7g+vCQDOkCyE5xGpe
ZGU3WrO4TMJmspbdfOGHoR2YqTp424q4R119w58sq6MR/E3BjGul7HMwFrEiXB3k
V2OldqVvazWgGF3bE1kebjs1dp3A9eO/UPXNM8pnGzv60WKhL7DBtmoxiqdcfaky
V9een09KmlA4INLQNr2Uf/OB2GLtUMKvPliXrHL9TSzTu58wvkekCUKE6R4rxv2O
076yRnDmdcOHAtp4aAZ6yWlfpxp1c0uhqpVlW9nyAbfwHStkuRg4MAzGHZvyl1ge
QXpytRPoxBvj6tWMttwzQAEY0Mxf/wgHCp6wG5yMcCFRTb9+HeU914zA9albWaOw
vX0j64aAqsrjHowpsk9DhTXXg6oBvtqkWopSsLKNp+ATEJ/g8+zsU2ZlqXO96Agb
/feshA9Hv8Ab3mud/knqnjxBe3gNcE19eZW0MfGEpYbYuxQJIG4s7eFuVMkzVLhX
dvuAozdRuwqfJiRO+YvsfnJqYj1tbVHhUMcvRp+lY27d4AyXNA6Cp6TLIR4KYZTA
yU+5PxdJj/D31vLuSbqtJRs0N1EPSzV/xqMmvBPxRu+Fh0vJnP8OEpuoIQz907Ra
9Ap3q2rO0HsOPGEVg+zMumV6LpcRgzvyP71khk957vCg2BYNLt89SvJf6fjjCP10
3F24hX5zDIn8VLbkHcC/9Y4T66q2g79ndibFHdGwTfYIbIdmNWsmiQZcYBquHhBs
ac6Cg/5fX4Dw9UvF0Vcy4DMfRCbdTeGV7dAaMhvqCekgGFKh4hdA3XHRyMFm3sC0
h2gAPjgZV1g96LO2ASyNL3A82c651Ok7nrt9hZjOUl6y31FAgeALipfh/bD4TGem
ye98xWyeCXdOhMaPXxAc+hYfe43SVv6UgvqyMVQFbrDkzgytPf39IZnhJuOx1foW
jm+TYJ0V9qTep34hVFnOH0yj3hkyCbVqMFiBsqsx4JaTSqN9l8DGGMHIUuxPiw9h
kCicnSaGlSiLMf88HIqjC5jcxteIC8m178OQxNgVOb5S4wM+sR8eC0PaD+6kwQ/I
QomU62h/AsmMb1AZoUUje9v/2apjp7i3+onqEijKjCsJFwmHx+Su/wqH1hLkE0Gc
guZJaqNMQPRiI/dnfqpTP4mf7lKR5cVXcwuE+FU0iUGL3MKuKYLi9iwGF374XyrV
tDiV4ZcHzzVLA4qnWAGH3md9JPEaQL1s/cF4rcn56dX7U2uoMQTryroKY63HZmPP
E8gbjdce72abXB8TlqkUYRolL1m9L1s76x46IgHSKHc5FupZHWkPnWZf9m+8802l
/CcXD0YKQ2slmg7fHReg6ubRLwPIT1M13O7WHVnbCY/uzHeMFCl1R6MOPQThwd1N
gq/b7MhH0UET/GFKQYe9jiI5Hovw978vIF/KL9y/FZddTCIL52fXair7ae1woJl1
wQ9PF05T3Rc+uNIHHny6+LOHkqnIMFwDFAqWCN3gekQyxDlxCTDWMamILr9D2lag
omN2a40XCiRHa+ZlKYS+leUQ51yke1A1NrmaMQnqG9SRMFhJ7QDqc4bbWDDDe+GF
aFH+BbUYk1jQEwHuZgXoVT7H+AMF9fzPQu4aOIKC03YnirD7q7mlnwnYBJzAwa9N
0E3STtVWhD5wy3TQa0YHCbM9+VEEy9q/nN8XV1V/syRfwd9RoQm1GkZIsfGYU8qk
ctc8Sb3gA/oe1k35cDzF16JGSAx9JacKnbuaHZGrdgsVWFr4kuZwobhaJEWwTg3n
xlaUemAHir4Nka+ZTXhqtUCjNCMzV/1Txqt+2JsrIifCegtpt1YcMcCU1gM7UXx/
A5k+BlA+IqogxrofyxCYxSQoTPWqraDFgWgLkINxVx74BC/YSZrtbq+jF5FbLggs
DamuviDUuOVgixAuIcESYOIntruakR+NUC2dWXyt1aKAU8lgzn2rIh+GXStV4Pc1
GwFmpOxCQT6QjtQyGgB4TJDifzq4tL9rtZJhVFgVU6tAN8dXgs6RdgiGmfao/FZy
7pakrSDzkuoBbdB4B0P2H3xCCuMQvd16E05Ocg4mjd2qkIpOPIWZMlH2ioYvzN9V
GxMdFSq/vBdin65CogIGuiS8nDjL5At9ju3FVOIZQIA8W01Dwdl5/zYRZ5ydwB4v
Kg/u6y2VtkzHrr8XqNCbEn26XxfE02/He4iaKBw3mnKt+lkh5+lCZob5aaPL1Dsq
5pd+u7SUNIMDdWaXcj0izHeY7qmdsvwE8bwrZtW1rut0tEMq91+sV+bVFHkVSduk
uKhvtqvmJ8u8vmQk8r65Kr5oqL2LLMhx60kGygBfIXKs3dhP/ts3jszAV+2zu7uY
3mDt/Hd5V5773eVObvBqDqElAfoecT093Pw8F5CcFjtzrAcVnFtW6e419oXCtM3u
EgP0tqO7YFpTBdwib7+/r9je/M1A5QESGaPH5zhCpmb6f5x7QPCsMII7RCNkoTQA
F+YMDU+SU0UYoB4PvFfJWQBWXx7XZvxBwu6cmoPovbBJ1+UlTAxix9aStPdKZaYZ
X8vNmtghyOCGIuNx1Qwg/Mq3UZdyjjvVD9BvpskkZIBrEZbdqzOADfVxuhHCDSKO
+Q2GuwES1GXY+XRfddQ9mQrXxcgh6KRtJf3O1428YgZ3fsApdl4jiKdDz/sdlNfc
Wq4vPdsP5MavruOKJPvUI3rWBwvnvH+Jfc48dshlIAON4NaKTHQjcYYwBbiNwARl
1WEW2mVODyhD6lL/OgnF2aUftnD0ACmiXkEBNtunu3YD0uaJzVfugMbXXP4mO4Ld
vJ2UFvnHxTt6TKje61pfhJQmS+XNGVaOyWpbx/xTrMYNgv5WRdBwaBumpU3qAZaT
PCJybXhq604Gvk3rq+fi8uwz9YeEcUaX9CJ4lLnbNvlmNHsBWskOt+NQTe/tnHOI
Zxk1raaI+Lg9vhZPS2HbmY6zzO9Pc6gRhIxJ0WqiIbE7fKMdOqa4u4PKMMMbUTUV
S/eLtwH++DWdimB7ymeT9mwxU1mZcGgkrvXppSyuXP58jWAK518Qdz8ffeOOFrIr
Rfrrt6P06O/s7cCm60J4jsqxXvOrW9VAlPY8nxv8xXbOTE/3Rbc0TOxdFT6P36tt
/fhxqCnaPi1OQyzF7iETP1ZZ+AZP/SdbxlpRvyV5HK1NsOzXDTogX3D0lyKvYy0R
FiDJQIOR/wlGBZsaQ71ButZMPU+rM2v3KiZoRWpRCuBr/qf6yDnH9TkkhDSexhIs
Sw35hvwMpiz/WT8ZIvZMtXYbaunhPd/8bpq5chFnmABxEeFXdkRyW0ABrY6Tw6E/
WwAotQZbVx43mwhLmVlFIMeiiEqY2XDSxgWmdwuYoEYIynTOZn54t2rm5oco5w1h
ES5kJUHwsCKxvkQibNazJwZykPdYKph5AXog8Ed310lj2e2vXwcKRniR4B40Edmy
Rl5eQxMV800l6qnKe9pyYooMiUdSNrr9orL7ePxmhnIYQNzwaP94vuVczcxXLXY8
DuqkY9exj8zJIANPN8mGdlAGMwkYz1rxX3aoOlbhp3UlUtYLWpmh7to9K9RJIM77
321Ew3wWrMr1mvUYfuNhg/54jiR6+ncTpysaflyqq8lM5F8VD98lMavaFLnUQ20A
hsC6MrSEHY4sal+qgKcMyZqpeYziA19zE8RkS4BbEt0TC07AHLtWpcemcIT0PRqb
S3n5jG750GyXDH8wTCM8rYW4x/H1PAUfyW5k/rEjncrSCtf0ZmaUXDJu/w9o9jNf
20zw/fzS5zIMBp+MCzVJwrp6ld48+Rn2F4RVF59wAAUPbNIByLTUSvZjJDNcTdV2
jqQFy3K5oZ4Qkbr/ka6+hNtkcpmeno85yAmYIH3lc3CTzKCoWtX10bXCf4XuVgH7
qZAkb+lWnfq29akTdEN/z7ROo0qYQefEYTczn1scQaK0zkunJF2xCN8Db3bAQREs
eNt4Vl/km0l6TUVYe/dFnXKEOh/Sb2AIwAGKqRjQS8d2NE+W2Bs0N79uGlennf2c
KC7Qt7UuBJhtqOjvodbRsuqZE69eQgb0ib0RYv1WyWMqdFVxc/ovL5vsTsak+j12
Sp4rd67/S5B7d0ncduFRW4i3Gqqxn3GYN1Tdg1tuhkUH9ih3XRcLB/FA6kXFKRMl
3kylsstp3IKZNKWWJ2SgA/+kAIIoteSJIrBsHxbLmwLR+de0k/ER09/Zgw3NKLXS
awPT6DEzRB4Wq1ZcodjoDaaOWnWFj6wzvv8HLteQ249UOgkFX1Nc6o57xjLM9nxq
7Dg5Myu4GtNW2n7x8BTaDawO37YiUyRvkPj8Nwxy8cCA3m52kNiHqZrAJ+S+pLzh
805xsrRMu2vzWJL8bonNd/pp60iba3V9D8hB1xdtXJ/y6h8dmKJOd37g4HCAo9bU
S9HpKCCwjHvMjOgSpwTCjN6n7mvS/1jFAuVqBIBCGG8GXjE3QaEZnJszQRPAjTmR
evuF33oi8b9oYgTJBCHW7dzNBzJmer2Xz56oaChQxd0ZJXgjzdtoKYxF7hqQLhlU
Ze73EUqlnpGgWNu+nD61d9NytkPOmH0uGa0a1IaExPh932qKM8es2dbnY3XvklGN
IHi5WoSX8hwXLhCi//tGivfPv9bdLqUDRG7qpnctXjeDFKxtT5Sz3OBRNE+xRLH6
IrhBoieo13dxipZxEYl4aoRqrECWQg2tijH5Dnwv4mT5LMsrjBZUMm57fHsv/XV2
LIhrNTYB647CA62jP0pPPe9W7ldUPnTvJSaov7xCVPC8felZJUOjEd5XIf2erKi3
wVwNy3b/0W+t0gKihFo2/VjHo5n5N0lVnAjcYC2LcrnrMeZjF/TeE0rCaCH564RU
7/AzE31QWb2EFl5IEmVKzYkYKDPaCRWinsIlVV13jAqdWZ6wf7qrV/mdWtFkz2xc
tdtATP0kku81G4qqr/Rr268R4hrj9G+i4pfMjMW51ugRt6GGAH3iGoqpsVOe0Z5J
Ek6r7mR6bVFr7LYk/6XdlSPiucp0+rGxHVx//YGLUYrmOocFXe5eoVA25TczYDqD
jaM4m40qVy4znl4+ffcMuUphRkxkpfb71/rDIk5urRqhjb/6GpFZXQC6rsbh3S39
6+FJmTRIUmv/4qMRrRRZxnOqJREyw1IfXFRYeO0/GNuGUGZ8T5QfImyLpm3f23CX
uVBv/bcdIricom0FxRy8DJoRmlqQspwMxdrZ9b1HDSMcZ7JvjAoAA4wwFinEJmVM
58SdkcUprZTyBvL6Ie9BBkrGG9Cc8XrZpmdYZ7hK/6a0xHuITM2hdKXYHDMEjmmY
UAw3FVr4ZOEP+ts2hT13SYRhZ7g+eOJ6aE9ciFwbGmnGcxaJhhw2nkDgQKcxPk8B
ToYKQX6pBKb+e5xeph8d38G4BdsoH4q/13dJtW3t6efaCd1uyjsBwsZHFervXILF
ZPCyECdviXOxXTKPJqoybWBDt8Cj2P+aXwm36ec6jQAqLOUFe9yXGrM8wdZPWD50
W33s/KTaz8QjYPkHt8yZO8Vk4EUfwqJHVK7vHLIKVsJi32xa6f65KCD/NB5WAreO
mZUmDNOqFcMQKNaydKR5kM7DEk0MnTOM5XFIKm+znoCY3ClGGr4LsL8ZdjApLI2k
5EF6+jK8GRq69Gf+sW7xhnYU3UMqqsEYoq8VXuyk3AQO+4/qUTcQiqAZFqst72h9
rtZezuYUOcVFV/e938fvEkOPaGBrr/g8qMSWVpwHCNBdyBBAHhlr5ijHo3eEnWaX
YtQYJyH7yggXqGKWnmrhnU0EtIT+qnobgbGdIHvCZ/LJmmruO8cq9nHTiNkS74n6
Zp1SdQRrtxi/1T7RYc265OxXDDopyd5mQpwYGHDO7JcKR5SEGlqNlrZvWOxddYJk
z9UMt+bejGzTJxTPseVoMVHvQ9xOxXOzvPphMvLVGJoVDISv6QcyRoYRnz1/Y6QM
fmK8uwzIguS3moWP04LX+gZQ6szvfDzAcA3UfAAhJ9ZaBTkhN4qolwMZZ4W+k2cJ
E+yfRAjkx2buzT95mVz5D4ndTa5FtLNkce036CB8BHnXPKRBcwBfPsjzXLY509eQ
p2nQTu7HO3ZTTxg7N6USCpZHWAf74b0xUkeOBFFC1IQ2NwzyTFjz0w4JjYuCRYE9
gYV1S94M42DX92RGkOzU4sW7Ob0ZKgJTJUrvh6JXrYKdhvCjiOhh8G/NaJRF84OE
ynOVMH3aRubEJAWwQsQma6Ryw1ac/MSv8yuZLp8kttRNEWCHNx2exMs/Zcrtqlo7
XIpS+NOZuvrYH6Uc4qu6IHouiuCY2dMRFkZqrGIyDKVU5OY3uc69GE9ZJyiGUe14
r3HASpU00wtM1i8xyO52mcEB7dyFAC4rbCPX49FgFpT6WUBLeOdtvznWAU9w/g7d
OcBqAeGxBibVls90jpMOfBb7L/mwFDfye6vD0FH7T0iAAe5XQitX6MPY1JXXX4lD
NCjWCf5mlBRvKVvVr802TWOme/4llfWr3Z04B/FcY+zUGZdLZsP0bB9F1ug6aKyT
l/PvoLyf2FW46Q0jrwpBXzd6pwequvwXtOK7LGxiQuAuj7J0gVTBdVlzqQ9ZEM7/
BJg/K6SCHshOM7Qmt4/vWgeH9j2haV+EGPv7+4+xhffOMd0Pfy2rrRJ6hmyjidGe
jusAXZ72LVD5jFxZKKKo9GLa/nEi7fjzgjWRQWypRQJPAvi2dGg8DY87Pb+X42kv
WazQ60RRIT7ZYrgmLyVsoQXdT/IZPuOl0sEzDyv1YQQ2/EXsW5qiPPUqg/hV+FUj
nEBcqQ8iJZDrwSQPj/fS61qvN/oW7+qfInS7DZMMOOxgiHiSzY6JnZSu8RMjDuOf
pfa8Fjvg8gwFJ7D6WiGPbdGqkqNRv1knN21NzG4XS1JokV7qxtonPL0Bz8/KQyAC
CpfcBDtx+Ow2WSmkTeQo2/7QqenplCutHe8UuF/hAX/x7r0zkE3yVk4XmMWJN6/y
vRdbHnH+FVJjFATWxMVpg99JJoZ3qpFu5tN+rvbhFbaHV9uS4dAdkcjG7ajJwTrM
L8w6Mr+NcSgapueBUQ3jpX6FUKjk85kkCrm4XmwF3Qp1FTD5gU08q5nRGNNSGTzH
6rHLjNmkJFAYUiIEd6bCsMeE3Di3PqcyK5mHzAS0jgXFRxe19SCfaNZ98IPQRGtx
4Re1ket/hAKVsmJdZfUqTwWuANYNk/D1w17DVqz4+smieocbmllqEhebqc8OvuSe
f0GTvB+vvlKWHQLJmRI9knGQIl89ya7olGRLc5t3n6vvQqtx2J8DsfNXMjQgfU7E
7pIA1Yrc+bmfho+84Dldhl0qt5XuAOXd2hzzsrqKoob0QfxPwlzlMbg5JO78+GjG
kLabY/eZKs+RQqPqctgnXophyNOap9AsRm2JyZBWGulw5sZSeFZ/kz33Cas90W3v
yFTae2Zv+ExakStnJ2O6pYgtMQCxF5Mr+Mdfzz5NxEGC9HlQNLLKdPtR1LZBdFnJ
Af1VpOlBiArH4iRQZWHAp2kYGkfUseRdaD+V+IweNbdWTHA6Yw8dyOICT2u2o+NL
4p3CcmAZ/Ad9mGdnS0wpvLi8msIukx1MmIoadkzTlBWl6LDA40jRF09xEgbk6NcU
YJ//1Z+lPzpIcNq+sXGPRNagjxuNfnh9syzuMk3i92yh/OLCXOYRctc6leFFqS5m
HPE7GLI8muaM2hz2MyfS3QbRwYjys6AsMYCz0SKuAchp//yYmhKeH3zakQQl09z2
QceP/s5uvKcwBTT285VqoQcHYpT6Bm1x7E5YASY/ccUvmRSw4DJMZORxb9VnViMc
YDlmzyvjL0FuFgRZbQWlw0Em6iwGBVRcMplcH9NOpv0+H1uGAETyoVka5p3HlzT6
ZREaQqKBQvEuInNd/xEo/tlvms1V+AO5OUe0TTSgB6ZGc7S9djYiT2MdM1Yv5Xsm
C8/maw3SSkrq6yRk3tcFfCKtWs30sWysXS71PcA+BwwNj0TYcU12QbFurrZtxdou
P1L+XNRea9GAdxMR94eoOfMq16SjhFZ3aisi/rot/3jizDLmeYFsdbf2T17yl8p2
Uhf6uCpIwZmNuADglb5kU6YHaEuDF47WxmXtLDzFDFGz6APTUorEpsPerwfjoB2+
Bq8LSFbtmteWpPSSxJ/IQyhhqs5LrqaqbPJ23fHUVmeHpegHs3hDBLV4qi6HaViW
mBPpDqmd4/meq1sjlGlRKfpBasLXkIfNH4LF1GFE/QSvK1fCNHBQiedoBYmHCiUD
RQ4Kc932EZZGXefVZeItNOGXNPQgmW/ACH7oV3/Pb5Xw2VUUTHR8e9OvOQUVJBCZ
AjLuk9aAq0ovF+9vcXs1GR4Lz8Rne6rpun4Q9VUb9MIQcthCFyA4vpsbnLbZdmFD
5EP2n4sZOX4D0ZVM9lX3posFbXIBpaWtHOBdsliRTNgoY8whdbjyrXUJA626a/aq
dVDRXlpGdsB2cQyT2q9/NO0WXqyiSFyz6kib2/SjxcnZ+TCVbgaOnL/xlN42PWUu
03TM0OVeks5R1AGDUueWLqyUFsdFLfWWvGtrgbbqxt4hq9gtu3+84saJc2ptkbZv
a/z/gOycd8lF7K42MKa8Zk/ZMPvvmcxNKqAYr82wyYTfgx3rG0o4Ki0Oo3WnOwU0
hclsf1gb8OYawqT6ogApVzaEZJPGgoI+Od3iBWbqFF0jbkZxQm18XXbOu0zs6NHB
C3m7vZ9VCbq1Q8dahj3f1rJJVW0L60Bj5HJMLceE6XXC6q41v89ggdJ+s59mQe+E
dvES6xuPtawoksD8F1AEO/KtIKxpUhaEC7iWu9dPJ+DBo3y26hhyf90YPQ7RC668
f+m0KNfRRCbeF3S0Uldwi0wEz1L8VatIObkLeAzVWBwEMKRmPPI8F8IiFCFh21BS
r4t6MJoHILagO3Q9GTc2f26hK1jDolKMxw5WmVopQaUDmHFNBxH8X74wX/yOOdjt
tQgvxhZfIIZ+Tk1vu0YIHnXFn8VQElPg53ZqHAaYLPmvOaeB+Nnl/R8TmuwsIwnr
/x2frLtEBbgPIb05EYpClfbRy8V8ZkXXqw13diERilL0NItATr/snWWSoIyHCK/h
dy9UwFkJG/EsStgW7iqwXEwdRemHosBfKzYML+iJwnqtWy47S52eMjkKs9edS1OE
Z0mzY2v/hOx0dFjKlb96qfVIDHOe9/cQ82FkvchMQmD5liizQqjk8PWzTGl51tTJ
2T3+uDtNXXjF5blgcjSnst8pXDx05twM/Zxh8Q6Ptgdmj28vkBdG1CY/8CWOisiS
SBdLqhQCEYp7CvpbrPgMlr0USMis9KUAr7qrq3k74UEiC+nuh4/RDtRHUL6uIl6/
2u5tNUpwz1j0oMk5OKPPyE/1/Qrh9MCilRz4mpX7zP2leuw+M6caV+Tl9uzC5OTS
4X8bSOiOpwlX1rqSJ5Lqy6ie0ExJoX6IHbNQhbK08S3Yeixxyyht7BG+oG/2TDL5
sZjo1ItqYUcyk8i8dRznL/aD8BFKFCAU5QesCbLrJE2jrc30lZZUqL82Yqpxp3jJ
1plkbJorr12izJpOIhP7dSBbbEzDwHnlTlchsufs1VUd3zkJ7pB0+Dufrmf7NLRm
6Ciu484isAHGhC6xJ1auWpqjQKoCCvZ3ZohEkzyMM1wi3W1KFsFf8k3dCy17olbW
ERM+6fuAEB6xhZEeJ8G5xR2oFVifwb/r108H/yNu7YfdCdrKnsUKwuvmxSMl4GeW
mpEsGG1738c91paKd1bY4wxL55TcQrcGPxYdB24ASKII/PjIBc5KQiLGrkQhRXz6
AfzSw0nlMe4RUOlX5nQpg6g9PJpsCaXw4Px39GDuJFWSeWB2gJKO7JgLOZU3y7CN
E7SLDU0jxQDKbGCc3wlqB8yB+FgHuv/Qyp+/j6ww8KbEul+btW5WvtIdgeFmKiPD
xBD2bYaf91EYFH7Bzz1H3Z6yBaMza8BDCGgTe4HpMrQKN/dZciR8CXw68g1ke6D/
Dipspscb30IJYtCvrkCXEKbobZdegAwv7w08NthMHYX1CtPexlxJfO1RRkLgwsOr
4VZkapU4LIsIjYVEXb7Bizuu9+7AQIEKWkpt5OoivZdpPS2LJnvBPIntlSCpv+rS
1oBjMfUzYxGwbnVSxlyn91MW4sLmzbjGsZoYSANC7EbzYwel/o6gSEcHsP75pdyX
J4VrOO9fGGWGKoS/iZawrTa3C3hz8iYUxwScIJFCaBWza9YKJRtFAJxDLJ3I+HLp
eh1UWxYVBQkFI5VMT9O+petlIQG0Wv4L7kNNcmMmXRVL4i3jiL/JsnpoI8Cdwrkh
E1AaQpIqKMwg9Ka+6xmLYGHAtEtldS2JpM5nUmFXGXCwr8ih8OzWrJ6BH0QH5Qji
CwsAdxeqWbRB4F5bil1giik95xQwEczPhaoa1dlE1/Jfvv/cNfXE/u/LUmVxdohz
JXIahKvmOzbhEO5wWIzQAcJnADcKpGQk3Zn2xuoBgyTdg2Eg9RcJ4owfQq+dS18n
LCiNjuyE51tYtzLVyBLwB+w02M6o/IEUhyFHkW7G86A4oHjZN5Z8Ttwp0Dss7WDD
W2wnxIbWg7BFaEGwRR03OGidIvJieniuNrjJB2K+tuDhgLVJmd1Fj/r0WLHGu0NU
b4wfJbPElMVNPQfUV25lQ/sVTFunx7zgQ26B1+YMfmamUgJXY8kEtNxQRKTeapNp
DcZNodrOu5dletddSVkQ/B+pjKEsMHYtvEr6NaN4tzzV4GqeylvcsPRfaN6tpkvR
f/Rf7ppf8SMdQ4Drt7OFN5XGGh4CNdHZD64vDLc178T8GBlTOlx2gck8+yrUbbzU
23NM74/41ohNYEbYYq+VKgSI/Rh3MsZetTe3u+sWRo/aAzIpftAGXOQznO1uWhkm
SEo2wtqpHEcW0QISoGatj3pHAmymqBJreuD4flIhYMmruBF39hb1DpNo6onfFIch
HAUrGWUObsftdRDpELmLKhOrcpgpqDyd9Q9evADScdJUl+ECQAYo3DIDI9dqM3iW
sKq6dWCW3QXRiyU/7mwkMKuE8WAZ7Wcov+gcc4jI+Fbh5B4TNTqHgEnWQeQa/CJ6
0kFqGqRA1A5NEalKoTEMmnWGCDJ+8Wh2ulIXEJxWMpxqNSd74APmtt5Wvm5UwDtG
MCFM0Gjc+iUm+RRG3Ibu1/2CMNOMhDPLhBSJl57v96c0o/GoETBHas7+NLl87awY
ISiJp3gye0v7dxa2yAHWhFN8OF5uIIsVm/LYi8ebCNhDF0TQAVewd9vOZdJf4Hjn
LRiVUUQzHD5UcPE2VM28LZBtJj85QMSRzG3J2acX4FiEKr+r2fXT5239siySK5ht
U3I0S/B/5j9UpkEnvP5MPBX912OXdDyKz3YRogp0n47ScJZMUeeZFdqB/lApz61i
p2i8TQyUqsV5K6bmzPTDwNddCQOwZctYb/P2/mrDHaYMNZpxW8Ga5fYm6wpKIUSB
THa/c/t8nqORA3zwWpXR78QQm7kEZ3n80GQU1xQelYQPJPwWomtApjv77u3hOk7N
WpXktvjlZy+yQwF1XhNA9ksKDPuQEC3joi2khyPiW6bMTJln2MQWXWQ/o4VcAYmc
JnxoYD/WRuYL5zYmFjI5nzAPmmsg1LVhtrzx48Ffok7rNf8pKO4h2SmfTyOT4jb9
IoVwwYLlKbGrbz3jW0g2IguFijZEfOlA4g5cSdzahB89SMVPl93HqMuJpuQS3ot8
jfAVpdAabR7XBcrnIezGDc5OADE3Seqq0dWlQ0dxDBZqF2O1rgdFqGwBbjJLDRdv
GYA6IQMtr9KF82lUyzCHAfd+9xIALKHUYKitkYAMrFYAnmTpL1bhaJytzCzLY8ak
J+BoznkDPb5VwiJY9id+qzimPe2jz1KS3+ziTY4aDs6QU1pw5BLRPmTbDScysXXW
1XA3kjWlzkw+dw0D3nOa9g4oDBzl7PjIp1YGwtsFPpyRq8namfYYAOb/oz/yPwCM
vwmB9Ae0j8OApRS1dDWJiu5gBZ5/qKGQfNngpeW334Azya5rlz5P2ttADXZUfjKo
WdwdB2nuISb05uvTbR3HpGZVmVZUfXNcLQ7Ab++75zWag9kP366qfPJloWy1Mfj9
yHdw/mohAcCq8Nn6AfSsnLCGlNNZsHHqeJrTDgPk1c68ZCX9HFLxcUNGObn0VB23
1cieJB35SMlG7inpzk6WQLUwMcwh5QH/X0sxJg/Qie0x6ppOkZxTn5BU5eUb4Pnc
E6rwLM7xofZaHZALblb6xIyQ4W5WyG815A7URDNcDaNGL5ihvDcs9cIF8dsPxWEW
GKZwUY7MWzVdcSRdMxW+aoSdRamTb7gWq4GdAWVCdiqIue2KFlMy5WgRv5heCJXM
nJGnbfQcUjR4UTr9TRMcV+wBGsZHZwWqXLaacyR2jEoYVrhjLyILHyb6tK3Npdrv
7E3PY2wcEdQGa8Vuh3d42RvAkJ7HNJuptpiEYTa4r22s74renpk2eCqGBDBLfP32
Kg8SSfYF3Po6N/rChyX/BxaIfhtMUnBqUAoG/P7cRojV1st6F+TzU8SMmfSFY3vk
k9H+O30JnbAoB1CvJ8oXME+mymRfY5U0jkvfl6Z7s+d5QDky8zHkWwbhpT8RLIgt
zp60/MF9EePedLrMmmgU32ckhxTe217d0Qk8FBz0BFw90mQlrRievWYBIckicRdR
RIqN9gTmlqNfezYfNM9mvyRR75rlCrNs3rs+rou3/h08Y/7ABf49MEb5+WLlK5Ex
VRmKo5RBTcJZ24pwubPrUw7VzJTheY5qnBnFLRTKoK8iDScYXLgeNAseycipSTjY
gEoS8ahj/pEw+QMWhrzapVqtKr4JmFt+Od5dHE4/r8inOLvHYVZnfWA99whjFlR3
XMlGe0RrDQNesrhR61ZlSZFpMbk6Lu02aGYOh5tCU8LHNeDh3HX7Ssq4w+w7L9NY
4cK6k9tVIdk19Ebh6ooFz+eZkaYCngmaPFypfXDUCtSLPC+X3mhMzUqem8vEGd3V
UmtVyCP46ExSrGSheXKuTnMN/NeBjnxJidqjiCnbeQ97LnW0Lcy5YvzeU3zMUnF1
uGLcqJz9jZc7uF2Ps097XgzHb+id6qAUWLOOVRwc9JN+KXatTnqDllOBDX3+6BNm
6XqIPGV0nGWtFx/4s3ttWm6tEOHy3FgXaqX/V2izjzsuIE2x969yE9Axpc6HfNZd
9bhtEGaUWLCPINVSJidwo1WfE7tc5E9mtJBHgzjZAamFLgRQco5AWMAk7nTRfIGZ
uXqcYzeQ2WYZu5f08XtDyRXPW7xjinB+6JO+NJqJ4zgZ89vjC1eYseyI3gAdvm3A
1NMb4q7BR2XXwnVTuaij5lTTtttP5yrxm6XF+j0vQKecjPiHVucoFtRGRbmpIlzu
s3Ap1uimg5+zy9xFkvSRFNqienRbEVltAbqIJQBFg5riG6llUSjcbTkDReJ5w2mn
s3f3H0q5NiY/iPboxV+M1e98ZMM0sZAu0iX47jRgqjQOuTujpA/dPtH9rseA5Y/k
/2FZOy08qFGNUf0BxFEBeulh9NkqlhGr0k2o/kFD4Zo4acRQ51F6LrU7aHE4Bm37
nH87lUVMu1Pa87HQ4HURC+rPZzR72oibsM3N5hg1wvb/PdQ84r0xvhhtT+XoZOaJ
ytffM0KKrGLyUGKTPTZpqcIEmpn4ApGhm77EuM6bfJUW/bMYGJOUS5oMuFhTyn8g
0cr33u4oWR1EMe81ukSrQKCJDCCbo++P+syIts7QzUmxZwolkzQiZysPxnA5aBkb
P7nS9RHg5VctgmO3cPeCRjZ1LkCCkcYGOkMoO7uy4KxGaS84jqYRJVOGyQzThxq1
8jPLwfiO+4xq0zp5IzQMvFjNAICQ3YsezQ+aM0pYMYardVupVKdqpQPYq8Vhgr0e
vauOxO6hNUuVF67JwmVHi1B/tXUR4aCovLCEl9YhUytw01GGnqZZS0CDTLum1+Mx
c5JAMbYrvFu3YyA2oT3Yhk/3kyJPTAzO3JKAiG8zqIqU+1QCpiR8lKu7Nxq077ad
KX33n8uywjxBIFLMfaSCvu1Wp9v9FSnMIDDwp08fw14W5rycWfmk7ThjRZfXUnze
4EkK72uIKnizniWbwPN2nbB9Q91H/XYZaBgk/PKQPV44/qouttn/T7//1+wgd4zI
oB6YSbMGUYCRox+6ZcR1Hj43xvJFUU/u+HToKwmtwWUJywFEZxmXwpJbwkMn0/PQ
ILkZKjpvYlCRViWOXa/tKtIxv5sFNbJaKfAsddD2nqmw7Bb+5+KYsIncRdWUwyRO
p0dRbultz1Unw32dTTPaaqKF+1b9aSVMqxIFNljhnMyy9r+AGWovJFzPo5kpXq8Z
NEg5gI0jn+hXmx1F+rbZ+IGph3pUBe3ZFCGj2/PLwBbaJvoyIwUw+rA3mWu3owfi
GT/yfgkydykbil6z7PYBZekI+xuK+RPuahSjcUTVKTYqZhPPD62PsV7Zu06aAkNv
rNi6pYvwzV5lNqujs/B79LOckKFlOoojatYpEhXdtb0N2oKrGD3EQ7ghKjtfZ/FM
ygAQvS40I0WaZhMiGqQv2KAg9bEA7QCrhxrGl9Vi52ViGi+Cp5oDtw8c49o672Is
TunLOfg6Yz+dw14ECLlygP1u2PfW8skHDI8GgaaBuWr90SYS7fTp2U6kZ/cMtFQ2
2kKHrlBS+sP/VHTNnqJ959RE66RYkSqxxZIrJY3H2LB9IX7LKjCxlsIIs5EtZU3K
9tsFSHzp1c2mk/h1ymmTgSqL3G5w3cqtnGuKkSEXtJz4pHyh3WEIM1Q1vCD9XU5v
M9MbhrDIgQiZ+4hXCSv1NhS3FbnOCz3msG7DbHYHBRFoBy6TWhX1+LRSABXSbOvn
q9QUuckedJ3gwmQD/iertkXBehMrVIR85XZ93SVK9sYa9saErc6d/4b5RBMj5snN
sPmJ+GNK/sQ1WWOJO7+pw+gaQVlf05aD8JBzq0UEw8t3Y0A5GbaYpHHbrgYEmh97
U6kvaLkUXBaQcDiOTm5CniTgRjSJtVHu2YVjWp01Tu32WB6iXN5dPSc+TYGHN8rF
XV/+S9KpJB8Hkqu3lK+LeJNDKP/O6y9JjB95SJDE2ubLu3ik7esAf06a4ANi694H
jiSBJvGALlonBxNrNTk1gYaVlmoxqu0pv5ompvfi+RYzwJoNRBlSLWT33xfwYi7l
1gf+4w0MFoFkxNlPQdepOhMpHo7k6kSa6iboQ9dU/6ZSpzPreKw3ln+zb4btQXG6
RplQOQDfLS5uLLqdBnfJ2lQK47DKCcdwpjv8zpU5MkHuNsVXdyO7qzsNDIe761yD
yHgVcatWvllk57vr99wfCpf1t/osq9GGF/48urZW/dGZyn85gBQs0x0lTeP5i9Ua
KG96qRA4MiJ/KbY80CObwKjTm+5CcvRFTOtLkEPA9tnV64PXnJBTrUBX1tIUqNAQ
hT56ttfruc+EHqvLMsJVIaSZ0l86XSMXJTICZ40rZ6xAeKrF4igTD1D8tSNOG+pu
Kcr9DfbD/eSUv2XxlA/Pny2DFlt7EA4oOJz6xK9EvU278FZR8xjUd0LUsI8YsGWy
PNoxy5q3h8squLjbjn9UKOahv2HykTsaqiL1qvqCZMK6ZZSt4vHuW8YpWBjLFra5
NIe6mVKms2e7+BW9At0XxPZXoTfX/OJQ0x2EoK9E6Gc8pgHe8sPCjZqfF+G6ggd6
l0tRAmd8EBcqmnkkbGsq8cRGehUtePMveUq7LhpYxcdDfR4ZEGiDVIumGFHf0Op6
pTix9UnsKlY4ciDrSJk+13qdcUUSwiBd81RYzg/BWdhM0pqw+S2DZSNN4F7q8oU0
MoU5cSBGghwFI88Mkwi0btICGwHXxTzY2SbQZkjLYcPG/yacyEWcVGTtUvszECGF
wSnC6vEV1zHsF5nrj2d7py72qbz2agZzA/IUstG3Qn6fBTMhOo8RMd/juqPs+ib1
FFXLTuW2bPu5+SAyFGxs7D4BeR6uwpCn/hEwAIsfGQTCi8ZM//l3icf9a8/9fTM8
5xAyhnObk8P4cm5YXxjGRnXwTLgWzlYJlLqL6mIG5r3EEzaQFsWsh+yMwilxI4s8
A9TSJCobwX7cAlyp6vr9i0NfgB72HAQ65+StXKVFNabnXkIuKfjVDHT43gx+RzB1
xHcVojwWIrm8ShQe18NcC1eypCfudHfw3sgQjclLGp08yo9p5+C8i+0WSpqQcdRv
TmrBdgcb0HN6j8vHcIcB96agoXufjUqspPG5FAx9HmhNucD39b73TX9S0/A9sfOz
cc25DKeKG/LgrplkHs5H+2wy9JbtwcymYQjfbQDm2uS3kaJKGbDhcsGjm1UtVS4H
JjOsVMJw4uKcchj2QgM41GUCpXk0xOrCvD7STR3VfK79wPfw9EBS2nJENXcFBahO
ccjE8bzCPteSl9FsXdgBQXblskS3XsjP6Pgznt2fXbIicnHg3gpSPQhygkEIINnP
n/voFsdTq5L0Cjjcyph0M2RdIzqNoHG3PV16wwSsqTkWrNP7aZ/AhTY2eQjtzVn5
D7v7ednozYA3YlPZGmSSsCBWvLZgh9ZcZmTdZOU/VQUaN2AHYVB/mnHyHWzY+Qa9
epKyW9DxvMmM4kbE8nxe652iTOI1vYTM+bFNA550rxKcSKVZAJOVMmdw85GZCyqj
INzLOaTL2jiG1j79s2vfCEziSGk+WmWblV1pbcg8t9dLrE9WZsB1HFsXgYnAwOoA
eIxn2v/IuMekbuXugu9mehacBwKyp++n/2m5C3gk0AfLlrzeSxwt86W38Vf2JKZ7
NC2CLYvAjes+64qAEWSQR9QQH2wz39JbIkRZ89QmyhWGO71RrrNVKtyBwbEdjo1u
UnSf5mauAnCUh+hpgmZuPubnzAK+x0yRrNxCHotHApzm484g2DD6mpJC1O1jupTS
fxycRTBhuLYa9UjF5OL5bSWRg8/+wX8/QXrD/E/HXAOb5bf3hmW1gp9kEq4d1kcl
u3eC+HzVC3Rf4GSN8Rn7L/G0Zve8IxKDHE5Jht+4wFrhuhj8W4XlJeKztSc2A6eO
Jrvc/xUDJm7B2Lhcrh0ZJsENyvqcc1mMnDi3XgazlaHYfFkg6l+Mu6PgA6+xTYub
/oLM5TrNTH+wYxNTwgpOx1ynA7mSBnmGekiUt8JRgo8JD2bLlBxg5v6vsNwX8xSd
6xCmzQNN+85m4oOTq4nDc0KUt57puLLHvzWK9IMGB8wPHQJu9iwk+LPmTiSmd+Mr
rAkB9mO2Fo7KscdyUMVhzP+C5IRp7Yy9zGKhLR/vp3JHRwk6nM6IeMffSbwLaP2T
oo8Cj+cuACC0nSwnpHseLYK/2G3LdamAnyahacvRoAao9ruRflUoz2kxcLViSZ0T
NTph+yxAVqwl4yxTjNw68N2apscZymY0ClZzHDngkJxMOBKy2nA3Hqte3AecUcAN
Ikm9QVCkDcQqGfaE+RRIQENC6I1OH0k5oupFBfFVFBp4TM63lOeQlVBPXtXQJlDt
fsXmxCvRad7cetwrbFHtRo1zTgsbF3NyUeWabFegBWwWty51oTgt4hIPin59ahP/
wI4U8b2yd4qnv+ANyn4vAVi+M25wPO1UBwcPcBHN31GvwTIDKK3m1/0s1IB+MscX
xJFe1ItoHRFtC8DB9MscRnEakrQHp0qh8EKJKXMB+1QlzIkqdcHvMOK5oCCHCeFc
FqdKwwf1bcWaM4TJk/5RnfkOvVM6sJBBHRqFcxUmkASNewoo26wO8LhFDmka+e+z
Yn7Tsi7kA8nesDoXGOJwvZVwbJQqeVQeKBrXhbxCpDtm0HjMxdRGTrzc7sOV13HW
kRwnMj3qkEWWCsSGWx4dG0UcQxNYugLB+1R254mw2TlwWv089yBe9xtPCcA1K9jW
26k3D8YV/tpV4/cOJOVvD1kXy1MV6xVFc5SktkWqwUAptaZ7PSHYrBrIjRoB3Hnx
b5bOMUE1vxnnz89743/fSGSygEDRinu9Mtmk44UdpLEwtEuTd8316IrD4rQjVBq8
y6t3avGf2hYFktltcfrOXutLZ4978AvRd3nvag7+fcMuJD/GoIZzNpjtcXdH3Dok
fqZTpc3G0y6wpS5jf5bMbVQ0wm+mfqoGzhzdkS8uE6JDf/XeyY5kehF7gtdgXWDK
bmwI+Ly2T8GLWpgswI1n48X+JPJatSixEwkmQ6KyfFy1GsKLHVw0PG1rvDbIbWP/
D8cUGoRxjZ40tG4fge11wv7wOBzf/ssliw3L0dQuUouUERRYBvFVY1hDBaeFKzaU
zKBnpgUjuF50yfWV0C4f4W5ril+KUI4OPmlr+BbMSs4eoCj991rVmk1JuAjn2Qrw
XCG+OVrHQO1AROciivePysPxubBD8SvfAl7rDiWObzVb9ZDpPDR7S+eU/H2M72jH
K2EmLV/+HRrRdNDu27zAAS4pv7chdWq2hqQNeSGRBpBZxW2vApHQH+AMMPUDwPGN
A01zd1ZHECGjP27py0VFUbdLdMNbgpGmyTse8JKQw2Jok8/PWpmdJqiR+SYcpaMa
1QUfcHHOxYgGa9qY8EIbIHGmhmOxDhiD315dbJsgpaTBR4XAEQCW6ebzDVuOtBmc
IDYF7mKd1t9SvgyiKT2fo807URlNmIgWWOMiDVr/8Nn+u7Sjd1TsvPLF9Pl/+53J
J/COB/neDs0y4ksd29qGhCAVGgpor1JiYWy5lqmQ0lWhWt1fWfYbRyxNuYLAZbVt
7CmjcS+rBKQbEGZ6zlr4vB1Oe1Nb1qRaFGxl3gi6RzvjbCRxnsU98gP9Stzoh2Dy
YWBkU6BdnoECcGO5lHTeU6aj5Gj+kR4h0dBbCb+MOu4BmhS9CGMDxQFk2gbvvzjz
RV1kkzMI4m94zsopNlRYtbjDdl/k4eiadBJSjIycK/xeoIxMJFD43KfARFOG2b0r
XhkwLA4FsCJRmvgJL5BnIktmWTkLDWLAVs7mvb0N9WOWo0V8ZJ0g+HAy4Czph7vL
Xi5qZ0z1ZVIDavWY5SpldxNrrn/PjWWdhuShgTqxc6s7XH5zZvpE2j9ACnJmVEhW
8dMbdHFpog8XquUlhhUG+ONWbroeyZvsF8bEUrVgwtBTKQSs2m5G509q/AG1MPxw
uexGd6VRWaWGhzzD9auBIqdhfJWAveHjGB9WoB82BhnqPkNE/EzNOYUMItWkhyvz
YGyRpRgfXAN7k+2Nwjyy0zKrIH4BU4e8J32daUROqPePgC5rCklEsU42rs5Smc6+
te2dgPZYqjl2H6Y+rxiHbSTd5t1STAaNjnpTDrxLppiQ4SuyKFK4DYfTUoFsmGS8
2QQgCH7sctty0k9eDupVXsxUGxO3uuDiUT9g2cqWaWzwQ+sGFznntFqbtE4uaXvb
3Uk7aSk6OzCi5qZLX4b9kly04do3JZn/FKT1CTTFHq/AeBpY2Uhb94G778BQBgmN
XHnDG0hPSYu9vyDYZuAs3q4ud0A7bx3FGlx5Dh9znmnC9hc2p+QkECvcyBO8W4zQ
eyMxe2hf/EMGwXVEmhPswajLoBn/NIAuvKllwjmZX8uxZ9svOHxhWiBv9IiylYSF
rtrkhOVRGy1p8QpWqHOOIbTwPPOAoWl1nEcdsSrNGb0bfL/khDjkHBX1rtpv2p1X
6BeuT0He7ZYO7MxdJ1SmH7JynIQxPZWJ4xP23vm1oLOsLKZNYBc0ab/UJ6TlUrfp
FhYJ/49W2LknBUw1P+1oNQrxIDxcY+ywMX8kHwBaT5VVscz5JnRoHIaauTKAjcUu
6YX4ewxCPPtcHXgiGpDyzwJc+dS0mG0G9j1X3juiGugDm6OVXwTCdj5susyK29mc
uduFcTzuF32qTxkXflIfcUzmR3mObcE2/eKde7V247s/T3NkMluFliDmq5wBNJqS
WavYBCebifCtQ2IHT4AFHsKnt0kO+L77w2Uz/bb63tvV2nBSJOcZ4mO0Oj08gvJ1
6BArDwMPmS1w77TRu0RxHmnWrHXLoZAx3DuVy8UwKCI95/7ENvsx6cwfNu/gYcNp
PcD9kUV5nERNlms0HO4rzczI8Xb6Mn7/uFmmp2MsaQjUYCop1ob43BG1ijHfN9Rr
yPJ2r7lcJl23TtXIUJ5B4wNKTBjz1FAczU3e0gZFpo3eeIoskzaZCNsHZMJYfgYF
2BV88MYZo2JU/BZHHe5K8eNWqPJbJrtTN9i6XWuZgm03jIgRTVPz3pIgu21W7GV0
8rPG0I97qmz3vMofBo++e1v8alql8FOxDxb9u/iTasWNCo+OtwVjdrJ6ELxL/SRw
AGeIe+MxtGA5rxdpuXIi0RVT9XhiyBXMtckOX4+Ztoh9civxS8CyEzTyWRQQCoj4
YMtEXjk6++s+UFewo7Uu+1sNlBg4Ri6XdZ3XZcJbZIhZerJYQV8VKh6b3zTddmPX
kLURmcTV9vmIDSb3A2VqvB1EzOiOlnNN4ZxclLbaz1QyulR2ypOI4xI5u0W9AnNj
6InhZZclCr+40oFcxYx+yOGFVuhexxJQ0vWnsfqUC1NLng4Jd9c/Eu3TpBAJBB5m
LOD6DtyIuT9U6zWuJlxybZdI4xOWKtwCpuGF51TJOahh2rwK3GWg57HnNZPjHoTv
ndh8YxRDzFgwmMK6L5iz03xdho/8FFb2LwTxLGpAiYZhlMaKXDIrVcMMjdj0SoBD
9uGvoLeebfAsqK4t78r1xSH4Tjc6AabJE1qACWng0p0nKSmIwy5TuC86cABK27Je
41uigi6lEmU4uPvmcWc/5dfGmxElU5KmaaWuHvO3O1Uf+RUWvwBy9GiFkRcUddG3
MbHMrSHIxiGs5uy5YtYRKAsUee4k4be6WW7G3i3NdiNKQtpzCqpNWzts+snNecQ8
UBVIbKkwiB3Tnwkw7T1KRcTbqOI2v6Ecagy5j87VABF5LvgIUsFd0zTgjHdMJKEL
4kHGAPdzHt2jZpmKCmcGp7MUnxSPCscXaxbABdSz26tU42bijB72XN57dDt1VU4J
bBS3xHrF5jqZni/DWlFOpxAfee4XhGSgf6yo9pJJZUGycgXQlXA5cvHFVwn5Cq0k
CbiS7AvUPAkr4nfx9ttyKv6eJjoGQdNL30IkkW7HUg1JtiO233Xkp1le6ufrRXCH
opZJ1k+tZx2kCoA80DXLQHk6l++93Vkt6lDRe3TLoioqElaVzaef2110CuJt72lC
TmqDrTTVlbNm+8YCPO+K1toBlCV4CzL6Id6329pbM7aEtpeO+DndXFGq7sI4ca8t
LIoX/Rdf2h9wIB5inGNBiH31OEoFLsGYPcFXtwkd8T4Wex3EKQ15xIuLHgy42Dzp
N8ZElJVVQYCFO7kG8WfU6PuwCxLKv2W3X9l2X4G65lmcKy8fzrab8ZGKoXzcqAkT
/MSELwzyixraLXwsJ3RXIo0uUpNfXh3knfSU14VllbqWdfnT+SiIxUeot0cfIdh4
3eFk1BcqrNFrx/D4akoyFvdSJBnYZ6LsKqg+noHAJPEy7YSfkHrURHOB6rmfkY52
S+jLumDrUGedn8GcIwY3Nmiv6yJIoxp6Os+uuko3aewxCYx5FJA28Uw2r8lHS15Q
vaPmbITBJzRbObpHmPCtFZ8Y0dMrL2dWNMpgf53Yyz41AbDqjBZYEVSYCRAZfyOy
3RUi1g25CEMHq7BO/EuyCwUVtgHxxeXtYV2RBsKTZkyw2lipmKMRWUDLZrWoBiQh
leUCCYxTXitDr5r8KWAVEjHfZVzg7yWVqSav3MFvXhwezKtdD1KWiYIH4X+qCzaA
ERaGj+ab3YExrPvt215GrckKplTltS0P4y/z1sNlLWIJs9dU4hoNj+GCyhTjY6yH
wm5RT9RyL6a/OaSM0RupQdCibsneYmbO11dYXyRggH/HU45P1xqPjBG71HbagJvP
Crhpt4sRVwG5iG/I0mvcBpWDNxJwsPErRgTwkGgqqI0PwDXDxEVanu9SZ4VJuyQq
r3M69pQixSz8fAK025wxpP264lrh+iWqqTUhKx2BGSWAJ4sHWHYW3wzdkLV7UDQC
8b6Su2dYO9OjgsXBiku8wJ2g4LOF6gh/b30/4hRwgVfm31Kp8cJaljVVHe9pS0db
FOqm72SdGk4TaNAA8wCbEmvf5JonHwb69KdpVaSyf+bVFomnqOOT+Mh3jCAOmAdM
`protect END_PROTECTED
