`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kIULhmkIrrzGCWXWfCoa8hRi2+81oh6ngdYholj82YI84kJdNXgQJaOL4I8zgi9A
DXb+Hi4GWl+SqULczjKvKkPSSUb9VoyxqrjkBJqoCmoaM/dc5buLKAeTH/hNQwyG
r2KGErXJU7pw7kNijidwrRuKf3bDPUKGj6w7Kmv1aU2ZEegnULmDPJiQwwSVHuau
qz5IHzBIONyZv8dZRouAP4rlTnE/2jbAh67vso4AF9cGpD5iviqUPaHOxhAOIduB
rdzM41RT8sekVgfloSl94dtfDFLu7FqXiRCKr+/3HAlhjtQUl1U7yx68LbCAfgRS
LpDyoOATMEdR//Ro3L57Y/6sPB4B4KEdYB/P+k9HSNFPomNIfOZ9ekmbh+kVw4H3
8/2gBAfmQj1ibn0ouYzB9A==
`protect END_PROTECTED
