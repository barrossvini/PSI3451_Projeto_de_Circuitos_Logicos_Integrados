`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cI45YV9lK2WeR+LqjsaBMgFn6V0I+G8G498A0gJbHrHE70t1suk131w4xhUQwC7O
Yn2M1WRRdxYiKEP6KLd4EWwoEtcAcgFBJbpBx5YygU+Z4gco7fgywHpsnuUdpO2t
+NMfttTxP7hsoOZo85vJWvV8ql+b7iXzYnWElcr461LMmJmVh11AZn4aWXF0DLw1
0bR19KEnRKWUa5Xri/xElMJHxLdxKxkx3Q93CQCOw6fLSAbXMX9HbGU5TOfCwfUJ
kyXPlQunefro0DvmQVvCcqBa4mJZfv0GtpLsMbHHE1RoxuASS47f1zkfWRjMxHhg
huJta/Q2gNDoEzNFwUoVdaV4C1Mh52wx2y0pgC9gtBM6ercE4Ct7XRv8S8D9XC6c
WW5lLOLc77ryBe/+/uFceYBDy8cHidGSMZhphZyDwautdSrcMlat1i7FcfKv8JJy
+mJK6KWS1Gybg5Cz595PT5OI4Tves+4CrnoTND+Ld66G5nRlrQInES0FztT3dvIr
kvmWf6wXw0ASmWU0j/It5QttGi4Cup82x9VPQWgrtJsTaR5ufdH5nNjYv26BfW2o
jBRojOWxHZJ5WKjygP8W4laO011wIf6wSZpb2MsChnGWviKF9ZQR1HyxA0RcJCMr
l9cvnBcRCL2qNtYcqNy9ydh91YPfzzAht29RCmddFsTdbdSJlDB+zjxm+l8toM7T
GyIDvVRXfT0SDysE/L9UZVhvbNiLSrRgmfM+drFU54rHNm79zObU+7PbtsnhEP3A
E/Cwk3jYce5fOwXjt2/gpNowg/RtF+bILIAyct5DTXU6PN9rVFIYWJ5bp1WBnXX0
/ThBGFfBrclEF3EtZUJlTtXpV+SsHfkXHennTYoKdzuz2zC7X8k/01H09JlP5nCi
NxmtdXHOgO0NVRfCTJep8d2VHXU0z98hjpgpzV/vYeC9CPbcGhAjzLol1JhPSnJe
tTWhFZG5LnEgi1s8tsv1mwU6U5a/N1P/UszvZHO/Uvdi4z6vl2EL+DnYzy3EVXaY
tU7AS+6zlykhSOQz/4AFf+yUew2qlmzMniwlZ+7bpeyEAq+6dtf2BjeSnfQEC+QJ
a4lBRKGUjD2sLin1ARDA54JqxJbl+X7bx6+SVmvmFLYOznnGIA1M0227y+tsJXCd
nljvp4VHmptaw9RY0fKoD5EaGls3ws66vnybKEcdnYPxbI6ugq5pLlo1lSILJ6pA
EXE0st5uRIQ8e8XfwbPOl63HDd2FMTkc0zOehfB0zdX9aSKT987xyJViFHgsLzG3
2X0oHGMXY9bNP8xYJDUP4A4vCZbn1K80fH2hmv8UCigLpO45jHG8SoXtCrawrOVJ
wjzwqHrfoQWGrUnMNX27JiThNgIEWAxPLT5KfwHK4y6/9kxTTzkNMFP94xSAgC7s
hdWhayAnd7Yfi81PyvRqHd4IF1wBQMO8jNSsNjiKSp/yWjeI77+68WncLJk6PbxU
3xeK/zP01CFl6HmmbI3+AmnGskjC3d/QQbXzFyGu+LkohtfJhWDv+tG2JUVF+Qkc
5TdebEpp+aqedCKzj7uXfqzqGcEG6uU6uciC0K2ha8+eln2OlQPH5BVKmjVcqfmH
ZwP8v1S6VdM+wit0VtI4QXpWysiJkkE7sAwqR4SmekmlQkiiPaAJH1MKkQcjF6FC
rt+tYLvVdVXFyP/Y+vls0HXPkPpfeZaaJIXGJFyGqvrE2L35sBhXSOH/xyta/Ekm
YSPSky4KtOHAA3BxOj5OLa4A1Mv1jwlpB6czffod416TjMBVvppAIX8DkyL372R8
NQioraVyoTrzyan1LK7kl8hH+T2x2tVpWfvltEUDRniojppFM2xTX63H3y4T1lQ8
hWVq0Pe1wuX9sfCLGqj2BimrjxY2EBM3MOwshn+L6qNHRj21uOX2vcTjAKBeIDqx
YgQmiLeB23tHD1WurE093G+uOsl73JyxTVbDiCf6BQvTtTmRoTRJSq+/jth3YISN
lQtG0KdFSPhjWubAaxO6abhdvFelLvDl3gOqbbvepilyhRqMxjCwivVGWQZvNvF7
pp0oeeUfcsWJsMBZa1LYXFnCPPDWVAP+gxbqQ+C3qdOU7wpqkMQSxsq1cMobLCr0
jajRLq3mhpd9441K9WbG9g3hDDJH0YI1ze2TDHBgNRdXdvmjyDBoUPaWQYiBNis5
NhasbxMpO7gmoax8SEceCefG9oeDBdMT1fRU0QJrVmFcWh5N7NAE/41LO/sRXBsS
oRZgk0rOdsL4o5PXIzyYQuL1/jOm46KiCi2PJJH9BhIZsvmCYdrfEFJ3tTdNaLNj
EqgHAAIUa9yHs/NaJUMOZLSER6xftymywoxFJCr6BcaeRD4Mu+tvAbk2/iA2FLff
mpMp6gP1LGRkR33U6T53zsauT+fZ+FT/7y+cbHFg6Tp+u6EnRONhFh/rAiVARfzy
40zXlsPCxtv51CT6wyorrsvnAq6XHMcf2OY+v9WnwwTM7CnfXoPRXe9VfsRyRhcg
G6CmFb3jy6sWbfYNWZaSu12ejwYfpNYai5fZI4GE/kEMacNE8LD3h219o1GGTnmA
VwoWXJX6AnsJjm2XqbIz1PFXEYBno+E5glGAhcmQCoslxIrtbrPVDk3ub+2mVR0I
VXLdgKoYC/IecCCmZPijKlpyRb72vTgnDf7/TPrfpRvxeM8h/SGArhYC8LSX+hqM
03DFKHlUq/uReo74SxjwJ3ieirc+E6isnirMbvHVJ9e2UrPQvu5tw7Zjsir8icsY
d+C2JpiiMuNkUWnRdeTj3CANDpf98gJ79wQxbOXe/60SksMUwL2PeRuuFzdhJlZu
h0vSRq26NDC9yF3ZAfNnAVZtYEdD8V+2dk7VQocZ65+N1N6e62s+TzKAU2hjXTdx
jyjmmhT43eGhgRfdHDafWMa6OfHruW/qVHZla9I05WJ/BtJeZG/mUz7BqUPPjxkG
iQcSOJqn5f2DtSinpYO2TQydpX5r4actGEM94b8kuQIpo9aQZKggzKQbBU8OHQWB
C/XrNLG/Cq8dUvdgnNlCyNOn1mkT6cqTczqiPt/G0N5dNmRMzu+uHbqQbLMN1/U7
2hlmkJ18vfB+8TWPy+6JwDL2Rhz+Wscx67FExcj/gqKW0UaWhWejBWv+m/FdZrt/
dWJrvD7RBtqZp5ruhoc6d9c7Px5WaGhPPSi8VVFToBTpqG8hYKZAu+7m/WSV2IXo
Lkjn72u1kHs1RHUJC/uYpjGsF+koNgpn44LQhywTEd3rhEGp8KiWS5Y409cJjZxg
jNGME1JgtIUWmN/wfsA+sgTfDdoX9l4JCUH1+obxYfHtm5S2RBdl7GarVHF/oa3G
uENevr0Nb32C17Kn2Ezhubzlav9PMkYyCE7hp6bmSedYlBRVYYKLjZ7ADO2u/3Kl
fBwxNXunquc43k9ybC8EW8uVmUh6UPWWJiPQVK2FzJfH8s8AlSICKiSqn/fxX9BG
Bg1mxMyTvtd0uZoQsJe6V3coB2wmIIKcHooDXgzjtYOCccMZEUdtTdmrHMTOp7gv
VFA1s+3dIfHULEP84x7HSSEhNcqofchAk1OB3cMHvde+ihMdDDhhDJ3/4Oz29180
QFPEDhrcaNfAunVV1de3jz+c76t69HCEsG8TXOboAsIll3dBDg88E6X8bOwZKSrJ
1beKrYG63R0+iTNjuEUhGzPtR3rqgWN8XlD8ZyllydeDQPVDaXQHuFbFxkgjrfWc
j3WPLbCqJTmONK7nc5OoLxETZtPfr7vPN8WnmuNP0eKHIsshtCW029y5vWc5hTKl
OEx+t1OR49caiWAudzzqFhqFdCpy4uz//VHlPuTtthJZZCoW4EcWUftSf6uOIzOk
yYSBUb13zNXGd2Rc2D2RzEymirBJ+UZt7jBo6XJioaMXo82dKZANK4OarqKeTz5c
LkztEoLq+2M7q1M7eTsxiv6FaPduUGDW5dgzjiPptCNDe+UU47XF+SAF6QzsEdP3
LK20/IiF+YXxGP2nDsEhMK2+Xb2aBJeZGpIraZmNerxfm5dITPybW3ar3RTweLy3
OAcN8NJ9hBv7sTG9+RPXj2xTDpugKvlansbels5W91UmABJjY7CwD0tCCsSCvuL6
h0nfSStxislhStP188UrM5ZAoZNMTmQVtDCcgjo0juXG51jeLA3lD5eDK2bZXo3T
9j404VojnNJZ3yQCxgnTFuAnAORczKm08a5OwUL7tmUwPpd0USYmKJBgOd9PqIc/
8MHmJ6O2ZK1IFUXMdy7lN2zxJ1XjZuSD/wn4szjWGSMl7yEft6JrB852+1aG1p70
TjtG2rg37f8fyfKF686Wav0vBq+P3XJLhlqoudQFDwt8Dr4iaykmvvCpCC0e/sGB
u0zi8nSLVkZsONxgPphDIUk0eyjIvrA69xH3jurvtKWs5M1qpPRB+usV5lXebhvl
26nIigZCbz7ftzGLs5y62O3h/sZECHllPXr2Cbe7f//d4m/iTalAFYiJS/qKojxU
sBFFKAXE2dnROw70AGe43ibLdeekC+ETH1kdzVFNr9xCSddgGxlp/lSCXi9gHgCO
a6dd3SVxyyGw1g7rO4u5s3ec14lbrfQEHdyV+MBULcmzudEArUGEC0vRfbSAS+Yu
GaBI07hItn+t/6xnxE/z0c9rE+qewy4QJpmcx6lJFull1MUoq0gvGgFIH1v8RV9P
6zwMKfCYb9qGFEoFgnKo5eaV7IoiWVgtwU/e7/a82SVmTBFPQuUU8yZxpZa/Scpp
H3TcgIzTOh9HU+GtTvHdZT1QFg4ntohmCnKMYc6/L6QETdUZxowHCFxwlG9DZR4I
Gmbkf0cuhAN31vT4It4KuZ4S355l5uBk/r7UG4RT73AuoVXq7y6g1HaxXpaULyWr
qO+DHNRvGLIHpOmcOCZ/hcQ0axdYkKB4RZzOGSX3HC0I2ESRVY7xoi5nRVYRlHaM
upMcsnlNU1D82d2vAdN0cyNJ1mlZHlLu1wP9Y4uvmroCny9ly496nSDPaCqNbF8r
vvt2GaBMpqsYpX5NVURssP+osbGKGuYfO8gYV1t56Ada62T5xL2m4kjSTq8hZgT4
OGaqZUZ8PuNHq/Her9Y0AJFsEtRC/bnxUWi/AODlJSUzD8nbvGmfKBe7cmuEXd4r
zQdCf3H8SM9sXonZARXE47yGltZOj9ZmC9bPRsMtosX4IBOOP+x4QaxctcZLFYtH
iYgy6dWcE4ZJo4+w5N8Icnjk0BLADi2LjuaEbnjbnNpXpDsHT6DG5ixYEHIqZ7/m
+Zh7DpXIJMsMtgm9mufXY+bbN+RRLJwN8bPKYVOMBd1YPf3gQcGztciEHSpzhawp
HuFG0kPcBIqVboKbbKGaUSZC9cCftprxR6ueX8KmNkxx248s1llSMIMpeHi9FX16
uJZab5NHOyu6zNrVVA80W96BlP6GmrDN2GcnAfMedf6keP8BLXXR2fyorXkpsF6j
mtdM2qAjpGrvKSwHn1Zmiqzvpo6zHyPisoUj9aJl/xkFYFEqKo/YOsuxFMG1YXeu
HzKQLwZKetIT5A9QwJhNar9Nkf4hp35anzKuZbKVVB4ErzcAQxKSyy8f/ujmDPL8
Ag28HxEb9DhQuCJO5wwiORjPIk9UTIvqTYm2GDQvXvAHfZa+cmC7+T0TTNG41HHN
gv9FYmjdmBEObUNsz9Czl1uStcQbjhk8k4wbNmTwMRx6ovFaFSp/wJjDtD9aY3rg
fNu96FUnwHA+gld63o1Q3tdFF9AzHF/EgvUFlXmI/xnitABw+KsNQ/8UasD179Zq
ZHpQgpZ8AKyA72PycalayxruZk3Pum3Iq8u2yVXZKV4MhwwswvLTF5XMGIaDVPy8
ui9mWfWfXSh6/JCChpVOcye2bIlYA8PTMk2CJorCKke+QhUmHMDW9ymdWCus5Umy
sNJ4ktJXiefqzLJ6Sahr0cd95RreYWK0ILy0ijBuemzdEPlJby6ZBg+NN2eBINK0
eg64PjTAi2cnLLx3ELdnZCZbTbS+jkczZ4L7TbJLy5yR0QfKz2JkNi2FPMhQzRGj
vemmz6TLsainmNTwPvLnJEWP+reSiZp+SWhsBInIuLRRmC8WiFIziFQIgggAkw93
Kc3kuTnZ1JT3YiKuznAczLQmORDtvq+8n3H+j3Tz1Ged6FAgqBQnNfFDOVwfWXQZ
unijWKeszzPnHfKe3TaNTSKUBsLyuQo84AQPsZzNm8Yq+0itDl92kWgudXrpqDjN
z6hJdmClge6wrNOElHc64dkZ0DarwAzCDF5Yfl8rpR7+sQnXF4JmgJrT6G/PLbBn
+WofMWm52EaaMbrb6tdLsSNvElIKVHTgMNlSIBaVk2hulSpRtjnYfs+plfARgxLF
6q/sckaSZ6XgZ3CopiAaiI/gp1IlsjVcHuxYBJds/eYAkju+MMlzfKjuGbX5Hun4
stwB/oAaZvlqygojBqvXwunb6Nj5VBV1zsxzHgOiXld1ZkW7C6tEkRXz33rrGkhy
oWJpbOPj0WN6Mq4z2JdQVy/3H0T/lPm9B1Q7BnhnxHFsoqjuaZLDiormmrCWDjj4
BeGPQeB9SPjDpr/om1jpuc/Mhw+KrIMSLGKNM7pzqj3lzvg5nNx5EgmTlXzlOUlJ
aCzMAqcNFmSGT9GcJkynOlA7DElAzIECbWP+HDiGCv26Ml/miMYHBmfd6P3avxHj
0U5Kk/7n6gfUrIbtilByTGV78OfFWpl65HkNbl0IciqRGg++o67V/hpj7p+Yv/OV
EPqDSu2PYVBjFUTKySXlZpvMhKH/UAN7xFBL6i2vFtwc+i/aivnppB3J4oWjLzHP
VGOuPa6JD6ma7zHD9mDDZf4C/UQZpE33QK8qv454TBendw1YLEDr+DXtVcdu549w
9atWe7HLkWAmqlEf30Cbczw/fQLh1z9A7oh4cd923Na0yxbDbhj+RXXvY++64lLW
358guF8lp1t0lY77152XgRM1ssx+k8V/99vZ2rNMEoPVkmtaY6NOKg/J9IpjueDi
BhqyLDx5/OWWnN94Ts7MdCXYl609XaBCz32pu2snN2JR1ffE4sNjs4kXRIqyH/Gk
0H4C9Q1mp/nS5IAMRL6iuNhNxu2Wgc0wV43nbfIQOZaIx+1hzwvSzQbR77cwFnPf
WMmOzUyVfdLh/dAEZrU0wBJtuZ3jECq0U92JbBDhrgqum3mGIEYBK//DsKwlRGDw
8OQjN+N5ufsKu0g76Z36lbJ89+MLl/XxHRUW1M9yEG9AsJDgqaENQ5ocNVhDelUO
zl0VaHcdWno8j8PT35Mj9h45Kc2iyymczPfj7hdvTOspSMEJ/p7G1UQik3Y8aFc4
PC7iw3qC0gnPsF3fhZBP95WP3KwS3Z+oXbH4Gf5rZr0A1M2F4jGTZSL9x18nsCUJ
pVMaGqYhx/pEqMp+0oYNlpyDjuinbgFCNCc2iIT6aV+k75cjVvMleD5jkCTeK4I7
zZjL5V/qYnqbSpIy+Rf1X72lGvRIBPzRxVavRKzKHkb6u+fjxL926phNOLtBrEeH
FkMPwqpCIWtyg+O6h81uZWWYN7AhAeBZ0CIE5ogSBX2TFvLFnkEgyqyoiQJ8Bhx4
PIsmBJbIybIF7CKno+xinKGjNhGCcl0Uqw2yrd0WyH4Rl1CDwWPogp3mFnhor2tn
wKgjjuNGddmtcq3v/c8M+A7khvlOLb78KmI0s4BN7pr4S9T661ihzS22uOfjOLk5
8427RL826LK576K3gPn8E9+Pqs2B7LzxMDZS8FhQKIfOuLXSIOagBQsJ+gI6UffN
esIRuswzAa8PX58F0YFxLIpdFEAl6W4tVTEEK5BQ48/rzS4OSdNHr+EExOMCX9EB
tLHOn1wvqWZPmwhAEDirlL1P1esCJzSGwzekxVjBTbjrfNiPnPxDx2lAIEk5evwF
qc03kSPppl033sRwiwnfeXoTGd5UDKuRKfJH6lI5EujlV2MvhovcxTrinf+wCBSd
rIMGfpMHc40Ew5LbuNeF+bfMg/4MmsAZAg6nusS+od/IkZ+xq0AuBEU6Bq2204Se
/ggxVNxOf307jMLgY7F+Q58++9RJ1Jo9j8WDZOquIwaWs/gUywUfJSEe+IRlx8yn
klw6jp6ZEiO4PHQYfzdB700vA9vaiTWm8hybKtxmnHNd0+8X1LTVzk70DEIKU+Ug
4JcRQtroCesNRL6V7lsaQ4uxU4nqVtdvgIrmkZ9EWBYQRJ+uj/K3Q52PAqUzefDT
wNRtRbK4C1jRRSg/bojhhezud0YX8QC1Tt5kHlYC20p360ManC9nwhUm+uC+fzkt
7E6i8GFalEcb+WsIp61UJhnlWk6WJsvTW3n9jzJ/j6axI2eMU9QqVEMcDEsXNeAj
qMqWdcaeMAYJCD9/KpTk19uUGlMckJYIFAT1drHtoKH3k5XgpGb+VbsEsGq2gmkL
OGVpWxb1DGpbMm7uQ3V7Thc0ADpFLgtSIMvkuaKHReGmaH2qAHqcbNq1MKmdsPVq
+pX59+i/dJl1GGriW4jf5Ho/wgfy80i0uUhANGsZ+XWxdO+cohmdEm4GU4JJLqwC
JY9W2SE5ZSRivspi9Bbc+L49cQ/AWhsbckunwut2nseAeXXAVEpp34sHN8AjXivE
vqEi1WmZjE5xdU5JiKZFr19R5IROKvvELgplEZYWCXIp6Xui/kKHMZzNe+hXRZBz
PjJVeGHgZyiAEm9ef3WAq8EIahDPjEVsTCo3psh7QIQlGwVzOlOOX3jnxQrqmWSS
OxFevU+T5BYwZ7FW/sIhdrOM5cPwvIqWH0SWIwGudAYSssJcYGgqO09McUniHi5+
IJQwD0gR7QlAQMf6uLkVPCxi/BV8p+SU6K7JvOmF3OF0o9rlsSSedLxR/Tblm/rV
+SYjlXfW0fKQft+zPMovZC9vgVgwBwLjGTq5r244RyXMHgNmbefN7n+EDt2UajD/
uWKwXfCibksgEklNp7qq4JE95DYFX45NlJyJYF/K65sPMhvvcrI3w+/BGcUOuJNM
AFwB4LYukJ6Td1EO04HrXIxAFZnAEGPvZpdhAO8ZZt3MsMft1psbF3Htcs8Ss0Ea
1Hkj5xwJEnnvgntjR/W4XEsFrGUM6qtmFvsA5FS96zwFJRYAsy/chLLDLAmRNwIH
mSUvfhBncESxxEkuJW+Xy4RdNeJVX9OfgS8dzDacqnVmJku6C9BQXmMRAwYHlmxv
UDU7IU+y5De7l1aR742I0tfZs0kokzfduGvoqkJatVW3HGkiabM/sDYR0kNvM9cx
e+/c5mkdnNQ4hmlhrvJdQM3Axo/8V8vQZo4yUPh2rovmc+06ljS7qladrFT8Ieib
pfYS1TAcck1it+HabxuwBRGMFBRvGmnGrPrOmXQu63R5S3bnL40W0M5elfCm6ZXp
2EV+z7YXpLHPAefsacyYSCAeyUnjuOVI73zOIxG2JxFCrnFLmPfadCqRwZ68Awyl
Quj+tOnVH85m9QTriiBQ5JQEZ5WDBRA4leu9QLH2BQkZHpLKGDJuEElOcHqCt1PJ
T8JNHvsQRMrTnZPmF0NJSy94RTSlVXh53CzFQ/nKxe2HpDWIHJJFCG8GRsfAD7W6
QqM1dqz1mqCPU75mpMANwfLBIgIj+TS9plM2nAnRQJv7kUeq5wgGilk2Z0K+lzLT
UIqnbGd9rvHLzwIyfuvx/1tp+kMAECVttYtzAPIOKr2xfnYzcm5DnyhTjmfxJQrU
JKrez01iO2iQ5YZNs1bZPV/NINmyFUZYSqpEVnXGMRKS0MWkXnExFFZEeMATD6l5
HHPfC7ke7+cT6zZ+LzCCdsZcjEWfglMYUG3jFhSAboG/ct9dwhTlEs6UJPisrMXV
XljLunXeGsjuijrGKeQ8MabVdYYL1TpUaHV5JaajdvyRI3Tyza9znttVkH/IYp6m
/mf5n2yz50M1K335zYcUO7VGQPCnORupjorUuS/mYOEIoSPijGZRYbbC0k/MVLy9
iyjzJtalNBsA48YaOZR3Kbh4mXsHlOOMaQmQKqvR6LwFYTTOxFOIL9adya/uLvgU
SDcPYQJS4yGIyxCnKiVEUhQxYj4c4N+U63kxoJIKiOkPHxrc0hkg+gNHDYjJkK1F
njCyT8seiTKbhz1ISRpUcrTnJV/N+iDAwHTaKrY9j7w/ss556bMnjPriQq+SE15X
sHv5kvkCfgaBUuAAlFIIZi0m3Ul7SracteJAyGPQNJzjfDeBx5cZ/GkQhFMsuOTT
2EncnazkWlanvfbJycdWhxk/ue5ktZsZOsfC+tQgZpTXhUYQIivRMju0wzZu8Ms7
2r3fJKqAHLWFgleeLHlKU2nNnhunBcgn8baLfwOSWGk7fZcHv0ZJfVc66CIKvGnr
AP5v549KD/UdRwf6pf9vtWcAc3+W7XoexNxmafUSYhcnlZLw0jeOulExarzfqe8V
wBZtv/gnt74QRSW7pj6CSiOxpVUb0h8rNKVK4S4frNc09JhSloSmmo45YGjD61Sh
LS8PEgFHUo+zb68/hmWZsyO/G1VT+JL2WXXElCqvhAvacc/SU53lPse3rwFInrLe
/htpZ/LHC/vhUpUW+2ic9nhUcX0cQTSJJAHyX/3xiCiQZF/HhqYPHH4oQ0eLgHHY
uGCmNJSVQruufLp1BN0MlDKHgVZXwPc0kdzIa1DIunvbHOf21tnnaekjtjprOItw
+YjtIvAEBWSpdkVbyUuSoyTKs4IZvpyZh7eLzRaqxEXt7VRRBgQlGZt+y7sKhsVY
UTWkkulesu9ViiFrgLNZdbfm0darmttHX2/L4kBrmQxngZVFYSGnhiu4sFAuTKYF
coJRZkcPvXhaXQUQC2L/rRiVt9dbtM0DL8905S/s7ReOUUuOeGqUfwxYOwxwzQRo
qN36N/bjFX9hGlGUkwGxq4sWbT6qwZozi6lrYJSkoGhjF+R9zldEt9eU3jVHbyaX
l3Dh7T3TZNwCpF7+AkpTD5cpF+f9psSQrO5KMkUr00FtOtBOMuBgYsPIzKEgz6iT
UCB8+7dOt8zxyYFzCqPSoLp8CeDAaqFftAf3rftUuVaotMrR4O7zTSqLBVl9ZwEb
6F+qQL/Fn0+udcNHEyY50DG7/vLFNcDYSZJSWqR1MYTaQCHVhceaT3OCZz4cBaqV
9Q9aX51l5vZTbPMWlUW8f9vfUctB1wlE5Uhnf6wDmFIdJUFngAfJ4BJI5ngIpa2x
adGQY78pU5w0lFfBp9vZT2QeuYSv8vs5tg6DmICzZpA0aSufBbmLRoWKpAQPgXpp
bfrPkmngRr7hOkVdDfiFjAj/9eV2/bZeoPAAvTuJA2Pj+BM+0ojbbx9rSaRxKgWM
wO+W+65/jknchmK4YYDpS3TB23U2Gdng8LVM99V3mZ9aOaTPJbUet4GPbEDuYh7E
RJm8Yz65t8TeakZX9yruDO5+Dv0IdnzaHUakD+FdOChvPbtaCbzptl3Aqs3htA/g
B7CgPHHzRylQAXClvR+v6rtqmVlUuri7lQ/noYc1ub7j/xq4ANvTIp8cQNMjM9Qx
xnsShP/6pW1hlddRXXmQ53PNZS6F+qx72EUfv8hfjqK8Qg3XPXpyWSM5xNtsrDoC
YLtpXkhUu8gof6IBsYoBS+tKxqcf7d6Gm/uh2nvVe8ncAw/mRXCjK+a1K8aVW/Wg
ut/R6M9i5t14fjHntu0GOSCn62jxtqydIAAHGe2K5xiC9BZ3Fse/qTaCPQdSKbmg
qivKOQcNgFsynXUhNB9AqOvzseyCTobD+wURwVwLhloWuzjr5lKEwPxbQqNxqpUP
Iq70CebmdbalCfxXJrM+RlOeX9IaRNYCaTdxmntR53GvT/wJmF7A5QEZxYQgPZUE
Ud+UVgS3FYaMAtzhGayaLxCtgZkTcs9KNsI1yBWIfsnYLRVaF99ZKG+2DyPB56nM
uK4E1Y2WQKl/vgaAc/crU5nuTw6tOuShzaONa6C8S0YnJLIhnqx6E0fq5L2dokS8
XHon2dohE5nOlLGOhralkLBgLWF7OY7hRZXZPVtQIJ695pY5N1Vjb6snizjsGakA
j+p34o4GLXXGep4tF6EzbwTY0kk/Ouq5x0ygHAJMp5ReIuELcKtC185cyXxqZphd
FlKdzqmP6HhvxXXZdJ7F9URmsVfKNqp5hsEqjsBVfuYcruD+KELJNiSWDwCrsEaw
NTAC3Bd7XBxqySTt8mqN+gJow/JdZdCQg9L7yaGJ/L34ktKIFUHqjc7NV9AXll5D
T17omnTfr1ZQ+Mt6xMCZ6dYjPZ+ZWjJM+um5e85rVDw7ovLItw45OInBW96ZY2OU
B4CqyU/12SC76Rtp6ojCdQuDvcfq1Zw8JHKEjkubllBWlSY1YG3jVGFlGE/Ldy98
jbQ3A62nPFOSV589aLhkhKxfZ1umTUrqZIpVm4r/3zDkWcfc0B4Z/IhGYlD+P75B
aeEVuiYg/OEAYD4f1fiDAFFJCe11UGnXmLqN1eDSBcj8WG0dCDVwKmMeF9IaNIhT
eJONa5MrpTGsrex2JQ17WmV4jnGa5s/5g0g4ouqhrKsjuQsfPI04vLN+rDptqbko
SDM3khlRjyVF/82psEqQuW8ig3TAJP9mNWlSJfY/ENElCww5G79UhWhxZr1LVim9
2KMNBnyTvkM+RXNBetd+V8+HDb3dpxAojY65zvbeVzs/r1gSjaV7NwfuSh1Oeneg
aFxNue1GHPAazCjl2KRT59MzJKQuXxzhmeKYoKf0e4GftmpsXCIkqX2wfNxgFH9S
fQFMMczPMdmhKZaVz98fyVtg8xaJLXrRiCOy6F+KzZZmCPYxM/m9vtK+B31Y/wSC
BgAc2uvS6uU7g2ixaU4Q7k18S0aBi5h7FvknrAeB22lh0bNDXpakT88Bf/DY8KDL
SI0vcfYCyossIwlO1Cq0x53px15nSKi7mdMArQukCiOuZmtL5jQV/5TvzvXR27RO
o8bdWlj1wn77SYULQMsEPr1foMU9Xr5HzkjMcio6HBQEibYYlfqAFx1HqDdMFfIb
BkkPHHzs3fxQ+ZS7Hbw04mWnXKsK2p1/Q1OoEhH+1+8XBYULNiUIyJ5XoSRxIYfr
nGF1JYNk+62AU8pQNgBOOhbgS2KJ+kBbbZk7GVll8BRj3pvOF+M0CTOdZ1FV2/5P
UMu48Brq5zAZ2KqOv3HTxxs+n9Ov4mTLmRYXp5ML7u+PSg/9/1uzl7Jic5w7SGg9
+uKuziGDBt8mDEU/gVU0M8xLNBvHMqwCAEBnz85tb8rAI+bjNDUtg/IvdWP59+Ta
2+5PbK70eJ7ixpX15gD2vif4UbmA6qVT5FYsxEAwo4AKILIHcfAMI8/VI6VyUn8b
jlb2+jhT8xy4TG9wahJ9G8epnFW4g2NrHeUiUtqArQHU5uU1fM1JCx+bzhZeu0FT
I8FmaiJeBN8gTx9oVgdZwqUGBdxBjn3Nb+N93qVfiYH7WEnWYYeNM231C0Z/Z4Wa
jlcT1frTKU4QjaN1BeZcCDuTQhfBMIku40xtvTQb06REtD0QfAJZgh+LhcZM3FvR
a8BsvfqQ6Jj3W5dR+vvNvZ6sDoqjQ/wXRROCel/d/x/LEp2I6Zxz7ThbZWEF+0QO
+pTCret3TZNJ4NOLFPiAc8dxLSyP5qJw/YTDm2gcs8ryZWeVhw+SeHxE6yWhq12r
s5PCJmZ+9IU3xonHQFvXnm/+o6h2bbjRtZLOpHE3ztOOHFKI8+SKHIrFUx+n9pFN
6afU2w0P7YlwvdloDz6fYtMWpXB4n2PYF4P3f5q6yMNjzHpORAiyFG/FZ5gtytZL
09OLMsmKmv8nEa/HPCpmh56FMeRXWrFqsSBluX2FpG0g6QLZDHQdzhhrkPWy33Tw
jz5vg/C8wxGT3nxZH1/6+GgD8R0lCBmyx9kVKlS6e1l0zAuzUVrC8J8MJMwjEMnG
Mbt3O2iF35xeUyrmUqJzZahdPtCpOIqL3mqmnHWVO3V5Nuo5tFsCWuyRdZTloOd6
GnR3XR6KN/dINmlFIN680r+ryjvvE7JMnscwMKC0HDy5UcUqz5Du6443Pdqwod2m
UZQVh2eqNyp0dXkO7NWcLjlqwOoCaX2U3XCdqJN6TrUT9hZBXBE9AAHCerDSfmhH
eUWQGtP4EKJ3N4DIRqDJgb1U5BZik3nJ+pC+pFRXONIiCGXJwkVYwutoghV5t2ob
MMZrHlSLBy+X4VNZWIzROblQB3i9DtdpbwJ3269IuOoQlmndGUFpk9bNETKHOZmv
q6WrMuB5cYHAaBzP94+2HWYvlle5ABwc3LY2x3waeTDpNoMSR9WrtmEoqE4cHHoK
yOh7tdZLN6MqS/wD3HhXTo2MSZdoOrwywIFQdXzIP2MTkozV6jXuqUsIoBf6mz3N
8WgpZ/BRV9JOSvvKFqFNZX8i5csGj21FfpaxH+jWC6HtAsAwvGCB1KwV12/TqhMV
ELvv8TRwPDRkiagWgtO9eqDA3GnSWffjacMG1LijK+eEqjdMCel2qyjyEfVqfmSe
4CRov/Ju4zGqqbe53KLoNaLT/eRL8YUIKKNJiLn9wkpP0TRe4IcuacH/aceIg2iM
UTCIxi4gue6mHhz5XHvn1W6m7jbR3udl7ZQhkkxoqxYObrr7LQJw4SLL3Id/UKpl
tqVrQ/Rzh0nlh5sF6O+fdakfBAgS8bxdd14CEL4dK5/SXrdkFVJ7J4kcrX+MQclw
ewbJ+miLKO4Yq7gEiu4A/0yICDsdd4sYr1IgRko0NDxQUjW587mPF50uo6l29SDz
zx4WfCwEBv2BmAXRATEhrbMg4+z+1oGN4DaPYpLPsumHoYvJH5WdRup2Pa1SXy3w
7O1fbmaA7Bn5bTRe+AWRruT8UPALfyM3H1ESNYCvtGflHNe0SCpCdfLd104hAmoL
Ay72FBkbGoiFWRiHoKHE3A==
`protect END_PROTECTED
