`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iz77VsRxh1UQE8B4v6RROTzqBn93qkFEJmhgK/JFRvnlpnHUu7ttDU5LMLy7LH0y
vT36WPu3pwPUPtB533gccw3BDKCCTnOpsMoW9AO+5orHMSAaJMAChBu4v0j/E0dh
DPWfQrHKaBlbr9Q+EVF8lgdUW+NahuNRzWbEpRsHnyexRMW1GLfQyyVY4FXgVl3v
hTJj8QZz6j+G4DiyQ97vg87j6bWtYQphmPI7TdlDk/H/DAl6xVYfIwtxwpoXgBAG
NiEPRm2Lcnom6aKGQxS4qFxBfYV5QxPX2uKhuMTdGlgytnzpLOi6zheFkV5M+MiD
hpKxxYvhJnsblqKGJowCpFZ4bejpA12VXrNHKlt4AwE95GsJM3KXA6anZiVSkjVf
UzQxM32I7TfIcW7weJsmDDtWKjYHlJbDRCwVCsG4JMcdrR9op5K0NN0neSOCfx74
qhjB/02OwlqC6cAGvAYrZ/EhhvmzLzza3tte4Jf5znrRm54Cya10xYkhAxZ6KXYL
jxu+aA9fmE5dvz7OZnsCxbL9msAKJYXLQzO9JlUTJB8=
`protect END_PROTECTED
