`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Hb5XrE7is/bKlHnxOTkvn3J1z4ryFsNNCc6Ni5Ftv0ndEyugvxLLNpOQ5RWKdAH
ESJkD4ILRhqGUKRNBzTNsvTKCggHCc9OPuvTu7vcD7DoEbxvyNJixF9psg9Pdto5
BQO87l3O+CIt/IXD+nHwXE2cgrLslOqyhvTAgRWlrW6igDaDCWAElNgQucG4DzyF
vKupx2LxtKm44GSHFLssBXVrwZ/Kq4+KysNoU4jHLDjY0YbriUVa1teBCH93LFOP
5yM2Pijeb8AFZC/4+jUDmubceQtIA+WzlwSOa9iJXu+EpYrHed6vzx071i2PZ92I
4S1oqN9dHU8eCwq9fGU/91f8RbDqUB2PB26p5v5x0op1zsJmp3QA0pLo+MjfOVEa
HpFluMSi+m1Os01b8gt1cUIkQIPH/T2Zl9KuIuJCnsd34ggMBOfW6lq4XUfzmP8R
oTNrw3RCOmeCYlsVtAmb3uJ/n1QpYmtl9P/iSsBtBzxUx+P37+DD47RA8hXMjttw
3AZooEo4BYUyXPMDqxwIBbZ5+HZn64QUitIF/kduPFytCe8N/Po6tlq9kRK2rAbp
q+rgJrjIOgVl5m+j+5sonT05CvKa7TnIDcZbMDU9tO6Jpu+nbkkliwNPAvUORI5c
gCm7kb40VP/ew2DZLGO5AfRFq52EOZl55tOQ9qA8nCrtBQZEXwbOpeLagsuEHzd0
UL5ExWs4GZVN2qGnCsrIYledtNZJwGmoc0LkPDrmFzoD7UiOB43Zk5wf3Q71Xpg6
yn1ujpLPE2mdjcm67dpM7mk1bomOOYVGcTGdqGnyY2un2OTm9jbYTF0+s82cFWZt
eoG/bA/14L6ojU3xSasi2sdFIpHEwWyzpia0scijKq4LztZOmF4GDdggxESH5adI
S7GjwSqVsYjnBokaV9y96D5UNYarE9iuo28d99HSiNoj+ggss4+p7dAbBIkWMjBi
wgXLLIrceRCwsC4DrFlIZqzAzmV9Cygd7Fv+ej5oOs7td2jjPdEkbetatacftfM+
YXkIcZCVarF7GIaycZXVbpX778ZS7M9+TV6n3Q5RMqm/0en881gnPDVCUb50D94N
sPLO33KINBTNJ840fv3hBBNE2DV8OkBBObETFg2+uHc3lahKtgvJ+z72p9bXjMPS
2q5BUnnSQKmjD95T6ovSq9Z8RwHzRAUQZ7+IAZmuz0rDawgkj8RMq4qvf+O1zUcB
km5eoIL+zlQ1w4Zchpixalf2IdcHJK/BgG0ObYRfRl3Ww0vyCjE6gQuGcSdSZ0PK
jOFRjr9GHlCEhJeyOYNVpj8BTfeX8RqjoBxQKa4lxipiv6fF4InLFjvoX5eE7Oxf
l0CAuXv3vJb4jaVy9S1CG+jtySandtSuhwiqSlMa4tdiS0ppaKzVoqvnV1n8AGj+
+DA88jhR0I8EOuKiBIMOS50b9XHSst3YLUuqp/w43YF4ngOWdPV0220JkgLM/gZm
wpZk6IK51EXeIMXE6i4PO7sEDWvfgYbhFGbq/6cHF8EI4QGJIjlCleYq6KANFZ1x
ZmvzACpBaX9ohPLHzFCjafD5yJrMwEe6Pjsul7D6KY7LDR263ZAFTkq2Ps39nU+C
ThEH8eH30qF434ax1GMu/zoy4DM6OReRx7RrZYw+kmwW+tLFPmiIZhkDy9lkAd4I
70ptFkjXxgX9Kp54m9M+XjRvFM0zqM1+K2kEwwqVVtoKQ8Twfapa9UiBW5yQoGmR
sPf1VdgEoneWWw104VzgZs7/Oon/skcBJ33nAIB6BPAgDcxhx3tXyA8HVrANP8i2
oC8Ofn5NbQFUcvjDRE3AcUTEg4NjX9Tv/doE4acBHUdnb9w3ulsyagYOcQKkGvf+
/7lol9vY9ZLrOwRw+zh9Bi5uXT2nr0xe1ywWxE+Cd91tWyXSv7931tnSmqCOlp1p
5X8MOpQ5HtUmN81ZBFzUdQkD95suGbVZOdxyqONxd2MIlZQAysTm8U/IgIWXyzCA
wXzL7Icj9s6t3Is/WLJ3yRJ71QspigBC9cWLKuK1/vevU8tRwsJiSzO2f4MBuyN9
Ft5Sa6QO1CW/9WlORt1jLYxwe3yjVMkz5bCif9dgD7aKOC2wbikvgA0XDSoCX5RT
go1qEyj8ZsJvjJZmZ2KacVNb4J6p68J8rAm+HvXt9XUequFxmdjSN69i8YwXc8U4
5pnHU1CwiAcllMv3oMf0mPilAxBLRJFQqsr2M0eKjJ4iGnmSMVQYdtnECf6Ti81D
ySOUG+PxbfNjNZ22AWDLX7iM1NaRW6c5vdDEyXqXMf3YrIk4SUynOwKeAuIo3Kqq
XyMxKmT294FvWUcknm0oEr6JNa2Zb2troEfMG4Iw7h3rhGQgcPnAPNK/FM/c7gqv
IN2L38IHFWODARKEP/sCYo2k3zXCdQL+Sym5NLlU+YAS7zFIwTQvNOS1esW4t9Pn
CyLXWD6O2x7IkbE89mvoewQmjgOwydfGYkR984KBav5pHn5vekKLMlIUSZUjLUZ5
QW8oJF81oxd0QthaKJC5alfxR03qiFdY+YVBTvCcjMw=
`protect END_PROTECTED
