`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVuqwdEg3QfmWRfOkTa83PW/O+assveEjAMGOwaEsvHzsOTMTX+BstqUZ+asV92g
CWVYoAheEGWO/ij0I1MvqDKK/Rg9pZU7I1W5Fk8PD1fI79YNVS63IRfK8p5zFJ/C
2WQ+ZlZvUbsZeZVwPS3evmiaOFqm4Xv4V6nMbmjnPoMByJ8CrFLzlcZU48yw6ENv
TYtUvAz2+Kx0V3NJYZ7OB5uF5LpzGt9S+ASh860W72yBce3kOcx3t9DRnchOvKwd
QxoNLdoywH3uJBKSF7/Kkit8FEcraKPYslXwviUoHsviUkiFsSrOnjOp8tyQ0+YC
cpfW0OSIFtIkjdsrG98k4clPpJ0edEuE7n1BZ8qCtd6qZ+GYCjjZZLlnHDdLBUNb
xTANezjtkkqt+/Qhpw4z0ixxxhoCc/pFgc/1eqrypGbflSbjGauK9Nk9aYjCu2UL
M9pwGhY/cveF/SR+S7vXV4P3qFBq37ZiSkzAk2yp2emaFl0pb1JF4A6laCajdGI0
PX5DCeHvfhOwzoPInWqK27M2oPCAYBk6X4e+tiIqbgYnKqcSnhgJC2driQpSieWD
xHuisrN78Ml1KltghRmpTVdhUHFJC/ZJie0VvOKDyRG6L9MS4LRAFNM/tBlj5UHF
MIDMrecceN6tC2H8P3rZ57YMOS0SFPmEnEna+9jnf4hDckXr+rPWO3g+ROMHiZwr
n+NIFiE2ridC2PBgLAF2e/au8KRmXVWbke8TXwbRY7P/duoPGKfn5N5EpytjcV5H
BmJiMl2/Y8KtYG/4rG+cA0skJdaDqBGTqeZ/0mLtR9XNvqiDQV0s8C1ey5Ze0Oay
I4m6vKoDj7dtSrOpcO8LttDQZmqtbYZESly6uQGl5/ko5XVXSAuDzEZ8lhSODul2
taR7tQonHwVmYiuBOnncDvgYMII0+xgX8QQPL/7o/h9GBCgoGTYVKEE6FIhEpTRI
8MAgx4scjAkPG47u5PNJsbFFlG6Sh6c9orVHlklTNFE2vfJy8A4TbN84p6SddoqQ
0MOtwtaBTokW7J6Mjx4CS0J5kxODjG5UNJU6OVYODMWWcpJ5VejuUG2O2bmCmP19
AVtbaTjSs0qqqfWH24q583iSj+odgT6rrFr/7VkRn4mCozec+NtDXmatw2pi56Gt
PkTMoiAGk7bs1f88Zlz7mpL3pWM9LpgT+VnkXJIl2VVtKgzzGA45rpbonALSrWx2
MBvZH+K/pfwT53aNDmWGYIcrTay203oMzL/W0VjPFRTnteph5NuDIPUaLVETQSjD
PCedEmbSER0i0ueVIuEzHWtVICXTWLRKj6h/6q9gBZxO9nlJqw6NciURxy3a8O1X
E72tEz/lPTYDyEzCaN3UZJ+NwUWpVwSfsjMfs5CpnBWDcf1aoS4JYmKMKA5eAKck
6LBStJaTBj9Dd4cLvCnWrBPUEhPxUakf1ld2n+xcSjdEynDl3GJZdQgkA8Qt2SLF
mhGrnj444lPvsAXDLDlC8bPokz44yhpE2PWBeIQx1UK8B8XcvwPaklN/pZm5NBOI
DDTHYs/m+TbgpjWfLR48cUl8QRzxI4kxmxBoPV+4xJSCOMpitLjwIDKLYh6P95kH
cYww4cVvoHcEEJ+MCxGCZqFO4tQT+gpcTjSS4VXx6WmQbmtRIzkt/a7LpUvff+11
QUmOKH9BIhm/NEsO6RvcVC1UWCeQC7EliNYjmX5gxCDAaKzmK/oNEQIZ6QYEMKfg
KIBJQh9KNdUQwlc5vQXTj3VzYpivak2Odg6sBXM3lIJ0FbIwhaX5sWFaJtWKg239
1c1iPKR6FL84oQXd+U/+/qfJ1z4d4Qy0dDEZA8r/u81Rljq7MSuZSnmvUZV3nY27
bYP+HcUx5F5dfy7uQ9x1peX/Et0JRyGsyWgHoJzilBQh3zk3toKyGtJ2Ps78edEX
R14JDdZkYQebJacYUZ/puYxHhFulekGO6BqsInvaEWMVC401a15uDEBpybnl7jWh
0g/4B+r3on+e41XEQnQPYYv97UjG9wDO3c/kJw14xZxZMHqV2WRPFVvyBTyKfpYg
s20Tjg4p+UVKIv+CnioyirfxF7i6KoJegCSHH9ab4KYPoM+RXnqjvYhT9NQe8bkF
9SCQS6KJvGmqzukiL0S3PAPStZaDnyRdjtJbzVhVPeUOCbCN/yjEfpUgC6L3/jap
/lpFMST3+5UL5qCKWeq0bUXcfPC8Bst5D81/4nspmBTChEj9CMDVPgAW/igE4eox
vJlAPNBJWA3n3Sw+JkcCSVdRHh4aOMYwHugnZ0Fh/7mpG2rwbcOxMCKZB+C5yruz
2udTJYFwQ7teoxWVuNhNeFaFw9Wn4KpoQsaaQNsNBsE6kcXEh8+jhxDfIBI/P0Pu
duo+1aI5bJO9Y8koOXz5Kb8/lxtXLt16cTXS9ylAVJvXHQdMk5e/sSYSJ/3jc4+j
i6vQwadsV8olYro7HDHsnj+4GR+ci0GQ75A6YQWuj2h/DrDT9DCISHm8KborpdGI
zFj/jZVsQkB/VcihJaRO4HmSj4l2SyhKt9cjM3Fyq9qS2SBJEvO7w5U0aDB/qX54
VVWtFiqC2dkx73pPpRJr8runU3FiyGelNH1mlrwQhF72FqYZnUOOievrd1rvYU+Q
zQYKOH1ECtbky3cR6fO3ebi2kg6Jte8DdwTnTZd56ditVFqETwww2P3bb300Pfco
ZbOdkX85Mf8orV1L2W9UQz6ecNIoxEI7qS3zUkLp+effAXLX2WCmz9UkhhxPXBcX
RiB1J35UzhSrtLVaHYlGHvMaw0q2uRota+eH5FifpMRGU+eb7ODCLg6KQ6/FKqio
g9KFL9pChKDz/Bx58gL+rrJGl9+6m041XtUg0yN7a8n61Xx0hRJYXmhYGLhXJ1Lg
TqpIQ/KtXFAr5SydoYo0r5TxfiRMtcBsC90CMiPttd7bjGEyXQag/WfRPDj8tqUH
RORGSigvScbZLfJBoltjcsSxvn7d+rRMmqWA2HMCJkXF2VAhLdXA7IfYHPbSnchI
Wc9cRw/PZpxO6/eA14FyxnziVk/EfeI6PrvrCkqhux9SWAsc4hH4KFe4tVTpPw4s
cVRCY14GED9BgE4+60tb8OcZdyQxQZbSANNUK06sSMGkVIXQN5bY1s+vMT/SyUXk
jdsarlfT/tHRqcgwnpLqVVLhks1UidF4bssTrBWIyoKUZcfq5GkKnuO7eZQEpqwn
yG6LLwMTg71WFN73xQG9GdDgclCyjydYs5CyDHAJStJ28MokvXDPMAS6K5nHeQA8
NeHmazxn6pdSwY6onorZ2fws/j6BXV7vYSAvQKMMAEj3hnwsUmyZBYYbcegvwfaJ
a09mgbn0Y0vdq2E4x55mpg271BeVb5Wn20tbZ0+7X2l23Z2JZmLGOyHf0AG15dfV
HII7bj3W0i2SZMf0zWdOFbMYEQpqcpvfISarGUV42C1x7X0VaKHbDL2bZrePVT9j
RF0DsqHFbmsSxaZtCr896goTgkmzurnAD8eQjwh2mMgZy1uF2LAtvhSEJV2hniZI
OUiwAHMfp4xbtD7N3Jd6vPE2tmky+mCMFloklI+7zTwk7rmwsacKgPTcdAVDTSPx
6ZvoZ0p+xpJkok/16DUGc2J4Xf7jvapbRI2YnVe/hleVC+5J2Nw08h8WqXpFNr6h
Cv2QMWealTY7CchWnPqp2w==
`protect END_PROTECTED
