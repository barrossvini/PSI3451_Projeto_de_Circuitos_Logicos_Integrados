`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0LBG/YZSplNMT2lEvS3eVDn4aNg1JTx+dllku8JHb8r1ikW1OjUNIPKYRF+77tRk
V466Jd/x2gUnkmhD2qnLZWURyCdyuEYIOIwDQYkJAkzjQAlhKJ09Cl0QEdpS3Zb+
1IBcDBxDoESldWZ0elBcGJG+Twh8Vk3Hyc2fYbnMrymX9a6oPtlYZxzHD+BaKQVr
RDOZOkoxw1p52+aaMJs1eQY/5uA5nSVUbcuOWu2+NDxu2O2fkOeAacStqM9JzBRH
srr9d1rvGpn4P3KrfVm5hLSPeWp1tquxM/T6JFrgEHoLusqkMtBD3mROVIQjoOYU
PV/ugrfayNQhconb2cZUhu8kEDj2SFCudru3pPQ5kjpt2mpGoI9CTWbzMEwlWjP1
HVWDs9zYAKbL3amkCZx8zfqSO6XiP7fz6OOWmQZu/FaT45s1DCAC1CGaUA56VZzU
YfGGspqwPMeESR0BHfazZpBtfClP1RTiHJXGB9YjrziS//On15jp2x25jAX0up/1
zoZsjSv7RHqcY5mrqpk4jaeo0kpWmtsS839ZWJIHK0+VPkGz3u0ZW5508w9abKNQ
FXp5sZ96Ac1DXF00x4tC1h3V2sYdejLGa306p7jySBQlhW+DT5WA5xIqZ2lgIUhU
WNiESucuXVm80l+RTBRsdC5T+bmsJlva2iCVTwh5zExfrLEOwicv+HE1PO/f+uQe
cW2MpoOMwij4AV0MtQQCyGnOLMrqQVnQgwks4p05/4RwQA+5JjMuEXm3HYL/ABYv
59PMTlMWBh/ElCE1BAavP306lurmzb3z1CFeWvp/LU2urBo9HCVjtO/+RXiJ7qZH
Wyd3jERB1RYfIDJZDD5PpUc98KXxh9db5MDqs24f0pHneKlMwdCzfXhVKZwUP/2q
njJBxo9IbCcMreI/VRXcIZOU1RjliNKJR/keXpUgA7mu6ml69oXAKEhCj0prBzIb
I9tM8qFaseVFkt6nQ+lLZIZs6h5wzKbdvmUWxN/QUbrtlamqsXli9LAkw/jMs+iN
3vGNucpaUeUt6obchQkzr+jSssspnIbW/GA3Qrp0m/i2hv/MU8fdrTu9dHXP90TQ
3krwfdaCtnia0bd23MCUvAfjc/cyGPgd3NwYvilmFYd+qYpAU6AnTzRmO4FYrg9t
4ClwnQIgnXG5PWcHjoFXCQ2xMdZZ6ORgAHRo66zfLq0benu2Zf8w/hdYWEsqo6UR
+D5qXizcqTtkD+9+LyHcXr94FPQlY9MK8fYhShNZXtDwXHTticN3ei2NBef55ldE
tMx7+E3oLYWe665aTUOG4C0NOnZsIz+ECNIwhKF6YPucb6veOMuRZP0rdoDCmO0+
Dl7zKu7pFeu8lJ5SnfkFY+ZZ/UGi72KGhVInBe5WDY0KHB39rVwGJHj9BMEw09Uj
uQUU6aw+XA/ydKRdbwsGujdxT4MgJSP0j3D5t+ztr1qHErmrIZvfSmefOOVBKhIi
M/jXyhNyMskHpiXrqiCnL9La/bczzG2ITUzKX04Zk64UxNyuMnF5i5swVrAOOs9s
5c6Ydwy8DRKnvphqKmpPi5fhTUTG/BLxCCIZ0awdCH03+pCaw+bd3r79gFlemeIB
JzvcxgSUpS9Rnq3tQqG55DWUZSi/q8y/FqrhUsD4weIAVvGZYE+PFohxRZ06xFib
5hhK24jz7pld0dzElD8/rkfNMUWYG2UXl4RDVI/1bPun+xdgyMhmhcbOk9ya7BKl
f/7y8gJoxH9UwYb7ib+jfU1gHArelhf2Udj4cVRw3dl6BH5Lux8iDr6TaVy3iOCk
`protect END_PROTECTED
