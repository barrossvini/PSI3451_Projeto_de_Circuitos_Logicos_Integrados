`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LndFmktXrVo6rjEjshLbesEFPhAn6gFuYQhuUXifQd+A5ORXg9FYw0AtuCpcCrYV
jbeDHUF25JIp5dz64ntstKixScSrihuzFyXpGRw5Zo4+lyDia/Em6D4Y+8axQq3h
0H7VRgXh8ORpGMMAvx1DmFMUZat1o9LH3vjRuyrn81LoD0locTDrxlIwBzAhv3Zx
aKecYnqPv5HYHaH3NXQ7z+D8hA6+yQ7ycKlljZWfKFXAAecVCpMAgHI+CDK5mLAl
bHujvNVSJL7UbVcSR0dRPLNl3K6xPyo/ayFs38ag3+TlwXnoX4jVc4nd77jT9XPO
R0A4rQnzBD7OtNwOTOSgMRYh3ItkBzY5BJHoFVtbHXbCOVbk6UV7ANDbXMH4go4x
YG4LYK595YdiuKGljwiGgt1iSAScdnn37YZPnYXHiY7PFhdSKDFNpvsIwojiLQ8A
auArA+yAiKi4uS0XBCLC923hQpyV/XPwzKnCAYFpiyHiFG4Tq/GSDMKkcyGPB0xi
eR2Iyk0DBIRG0wW34CafEsmlNphpDLgqmbn452ewr0VoKsMbEVMT1cce1jYppIoa
tCFQ3H5Ndgfbk+xRmsNW/wnyh7wquCOljo7y2mEb4tZqn5kerR46trJ8l7O1W8mC
UdqpYT78uy24KtfCqFuXbeeIPMhdzTN3YUW4RNbspQnlVTByeMuNjBmrIdW6v8yW
W9UtLgsdmHEPD2uAQPZZ/Q/G6YfUvm/mzsEocPX3HHENSVC3OFGgCjPhhBNfFy8C
EOGiQ4fnOm1psa+EdwBk3GDrnk/G4lvdWiUqN4+DQ2q7wqacuf/rwJtTy+fvnm7C
XTQ2nL5wtc1h6cU4mngdHpycE7Ysz7bLyEGLZfFKmnxhbiAxzf8qeKactLeRnuns
jbtir9T7ztERJIzwGbFWESAR2zgL4Q1GvizZHEfdkFomp2/QkBmzQ9Ls7nZ+henf
Yi1D4jwhsGINwuphL5drEdaURR7yuSHvGOsTs3I0iA/I/w8o2p2JcPmzcEDvWa36
H2iskciZ6ZvmTtNJLE4BzNHDWpsOadGzpZdzj5gE84LzON/BM+BtbVxWhH226dNS
rJ9hbB8W+Jer+kBH+Wgi7F6XW7D82+mfRwol14MC5W1Okh0TD5tECsWTh5WiDycl
BTUw2Buc0UBNeD+g8D5b8plDU4WcCZjDeK9Bb8EeMXGyIOPxCM137c71aHL3Yn59
Ndxm1LynU7D6O/09PMVHcI2W+Xi9QnCPIDh7zm+be1GSxmAmZnTI0hnjPYZGy8vb
/FP39CyX2+G9VGru+FJJIrZGD01gkY9OclDm0OUqmXIibnkex9GU4XzQeWLxuoKW
zs7jt+KLgB1TZVomd8HqgH+pOKIQdReAWoiWg7Z7VfJewe0e/eY/Rp3/n7d3Cf24
cKByIXQV5L/256ZENAQboSFw2hq6dF65RrL6bJSSvGjgAFHhELiDS08VAtm4jIbm
d88WOQQpqPyM3ovfWb2wDByjuK+RZOIQExHWZHWQqNIrMFf6ocI2fhZAdIPUWBkX
IchkaaWhIR8vbXDRis4wWNo99h77Dn3MWAihpcaCxpajHgJ4P7AYBbYg6LeROTJb
RuGkWsuu+K6K/pZwbKLI1HqypaTES7JcEgzzMEh2usEvoHjXtHbHZXoeJbHkUK4v
lCFHFFZv7+c0zFSfzjLC2iva82WgbHnQBOPCEJqbZJ+fKUkFDmEH+xIbO5G6SU0H
s5kuMwCnOAYfFBt65me7/00gNOHdqZlO71sUd/fzJNjA4DRDA1jwsLhpsOtqyxxV
zbSPPDrC98jjN1aFg9IBnJIeZKdb2Z/AIzgrnsylu6xGZN4E/hdS1egeLu7VOrgy
b4vX/uNoJJiVccxFfTGMtKFjt7E6sVslVyWv5/474GIIjKFEjxtgIp7RhiX5peYo
3O7Ygn80/qXYfLwS//PhAJANKmnOu+lOc3wQGufCFRQpcLM/9am9m34+kz06RNyd
sFbC8BRPYZaGK3apRC8U2+APbLP7dnWGhZ8LGqUrUMsHvnG7hoeMFJCfQJ9sL/dg
qdHLT9PDV1isbKNxWVaxiJApovHuED+2KtaWHHP7+EHoHYNIb8EL8p/Dzr5CNkb/
xpwkH1mk2++fhnT3BoOe6aH/+4s+8+PDB8/rk2UCutcpsxvXsOVi/wu3mAueOHa/
HjGDCzbei3X8HOQ2SehMXi2jiw82sGxM6QaniqD+oBUlYcY2/4F/LwOXy8Yi+oW2
wV2P3T5Z8WoF5+qqpXes4LP9AJh6dKJ01qvTfumBmK/3o1RarBHTJoEy9NcLOoHY
p3tylZi+voxlqf/Z1Ma8/RY6+Y+G8g3xjxzDtJCykv7CnWwtBYNdYGVkfZNrvjyB
d1iHTVvnN9BWi4cdU0Q292boQ6M9UlG9txg+871Ha/TDiuFCN+KK5J2BViVjcAo5
zPJ8NhPOg+ryt14en0qba1D82E+G1UiYdm773+qVLP7UNF1xmcd57MBcBmT0UKST
gdhH/aoPC57t6y2Px2Kcv3KT/PkIqKYnso5Sse3Fx+30/oIMMvJBZM+m+sljQNUm
7EV7jfogTCfO7GnVzrv4kbic2iIChYJtvVbIUz+pbRChc2b2GPialNe/d6FMlj6N
ei5S5CkuaCX6OguyjmgkZR2OAfkrW8U7K+miSd99QZIHPM6zVijleI2+WzJ+W7Ta
jbTrswRjrd5Ae96ZNKwHkt/lACQ5uQdzwYBRtJTD1YwfZfsGcLIJH5HDH7K5vGsA
J4ZHBaUVvEPaMiBhpgj2ygXnNrdcgjVCMY2GKrrVerE9GWECYrwaJrDo+tbImh8C
X+Tx3qphNILUfA0UYGQ+0anMVp0Qo8+LJkJATFzXhPReEo0RS0ZwI6OcHDZ21k9B
eogDHOWpfxcxjTIaZPTx1DEYzjkh3HH3wgdgTNRRFb6+jaPmNvxLRT76xrBK6Njg
HrNoGQpxc5ylfcZYyvHS2HWCpmf8tR0dS06FpcaZ0ET+2dbvnO5mVJz4476NZP2R
jkID+rioNyKbrRxqKFBzaoxXSApwdvWdhoHo6x7SpouxvngCYzjxN7WmQtmzvlRx
gTIcRb9CcF1hbFmGlDsWYpaKQ/xvG3mqfnOL0L4ZjasJdvvI9c8ihegkhrPb1L6x
5S2/9aeSV6IJOqdnB1w6ZJBG6LaivlwL8QQ7c1mUfd/RUq2eNY2q8+FKl005t5IZ
4C0wBPrLaf5oL7zU8/NkaO00aqrbs8sJnso0o3Dbuc/VP3BMwXxVf/9o+x735Z9q
N2Pu5/INsfDPRMCuZLMXObDuw2UVZvjMap/lpKx2owS5VCviJo1FtBsF1TZs8OeV
k0ic4B8X2xERxXcqxSF1M8bDujiNVvAHIJTgWdsmMpDFrvXJn45lCKpYuMdV3tpk
ee/UxKECzCPQRqop5oW0i6nh+r7lQeaFOl8meiYN8aqiuZBjieuEn+E6ALA215Fk
Uv6vuIplv8IONtj/3KkXQQEVnzLZCvyzSixqxE6ZXtF1PiCnh+zD21Upy6ykKPH0
JH2GRumz+CFYDOvOIgRLpds7BPEpDAPu3lFJljzuYsG4jhOrP/zEUWYm2EH7W4Jp
0HBnWTJ36Ml03dchLCTAi6kpbf4h7tKF3Vi4GKGOYhguCB1liovi2nR5fqQ2vBDf
HZqiwsOnxMXFi/GRbwNwjuDyWw+c0Or7/hx1ou7164RLC21ynsKMU7jCzbt4zM2i
cLuC8G8TjfTB54A5sFhrRYIKhukG7ajTcRiPqeibSFud078aLX1rhamn7qnnjMP6
MAT65PZ1qiy4XQmwEbuWBucXVzhU9vqjzMsjxXWScwKZHQv6tnnB3aRJ2mwFGssA
V1rXeNNU5Au6OlshKtOvozkJfhiOOWIJYOsoMtgioGduaorx5Dr3hgbEiukgbYyz
sBwfGtcJaR+G9JVevJS6IrtR6ucGg5b9ario7aw3622jMapv4mxIQZSCUxhqb2IZ
sRD1IB/OasAChpvwgP1hnCy7rZe+pId5SBX35068EhYMC2paMusFQuyFdGgAUqMX
xqigSk1nfngREgv/6gH37nycaHQJUT2Lcc5FgMRoYUrvf04eueVX0G3konD7IT3y
BhSSvIMVAQHofEYACL3k57osSJejIypHkWJjnydrIqZqfgXHE0SCU2jXFwfbReWD
a93RkJoHfN+pP7X7/l85h9LtbgpDki3xIgMSdGxckkb4Jsn8hg3SzOWI05cjFzk0
JvNPCUsW2EDfAK6nvwONc6C94ZPiQJVFZSLbfXXPmZfV55v1lvdm9ZL4UGB8E6IC
PvTOB9GYpdievrIg07ihR9N2d7uF5Qn2UrZM3NM63ZgpsJtuKPRB7+yhx2luxPck
GwuCgnSVlMQaaTQE74WfA74hoy2idCsL6dtXe7/vCDS0umiW6g6kiRs0lGzVn7tr
Dq/IhxeCm5jN6VNItt64XYHlSIoHoQCp4alFE24IQ9vssTajFUcBa9HwhDhUWd4i
ki9SCQrpIkn2Gma4VEx8VkThe+sAT7mv7ySKOYz1PULwuJx375WsjvMMpNT74DCX
ax6KIsqGZSDlsa5dJLD2WF5NYU4gd5TS45QdyItZC3mVMQ/0XAkzLWGnMeY9S9UP
`protect END_PROTECTED
