`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmRg5fwlH2ZrGy2zMrH/uRFQaMOgvesrO7YdV0vga66m60R4ikLgD/dpmrwVme3y
z8ek80mGAfbZTq+Q0NTQMn2MFosD6VYIczrBjs+P/syghBFTAWxsaZYQ4JrLIIKv
S7SJb2jYWAXAAdVoAGUEjv0VaMI67aLdOeHJLg4idQDY9Ua9vkTRGUVNpiMXtLZU
5VF9xaH9pgFk3CEsnMRSlI3W9wdJzxaPUr9446t7kx49w4vJTDmwGxXp4hEVJ/+8
XEmuTvg+4Chsbq59aciF1IZP+0Fzy7k/hC99B/MlZQDZ4aGkVdsCTcmNTabeCNqr
DsJkVnsCTCJZnfEg/2nxZMMu99Oo3ivtA348tyuaTY93sDfW8CiJqs87gA6twzcM
gX8kkRRVwNIucl2f7m5OeA==
`protect END_PROTECTED
