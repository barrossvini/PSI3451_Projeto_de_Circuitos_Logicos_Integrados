`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wJHRqfg25QYZ20d6F8uia/jlbeni2KvqyG2nNdcpwqZAQ23lK8GM/ayn+V7WmL53
gnhFDR12fXSwa/amknPiN8fqmKDkycsKjKL5VJY8e8g2W9HoKFESNzRMXfk+Ig7M
15NmIJqRkMaj8dpdhxwfEd+2T9m5kTPEFD098FWEGo5dW4dAbTrE4+bvUkJ5ZKpc
xloQf/W9YRYexFZF/XqMoczl4QnKQywugWx9qcJzscjdZy7mCxA8uJGDo9v6Mab/
E4hsAGXRDTicBU700pNfxxcQsi9ACg3y3wQRUf2dYMPtYWPtMdSUGEfWk0+AOq4I
RMkVFEXuuVrmM16fE7ut4JpBALsUxwtAtnPuRdyf4wXmFFfbw7C5RJ0hjl3tEeGc
2MaXokJzK7YGOA8gTOOvrHMkjAKg6OssgACGdJ86iMVEkN7C8nhuvYEVd7gp8L9H
c9npYl/os7wInEMxRpE4yMH8YE1gsiW1DWQPvy+7pKkGw1vkir+FrgtP3jh3SWCp
8baPs1L76K0xkbSx5S1AOzWhFIkWTi5pr+yQNhaQg5kH0vPdWbiPiiThYQ5WGYew
1QldaQom/x5jHF3YCXncVINPQ2pNLifuKWzST4GgUS/pc+sDYHGrsBi4FZdIS7oX
8EUPgpybg3nYoVLzMx8TgclMfpw52A3ky61/bg7yKqysE6QmOD7EvolbfTqZDDGM
9c5FgtkGUNxliqPJTAJjw2dZQgjO8Y8l1p0VA/QATGdPT+MNIb1uPVve30m8Ieat
WiajcDA1YkTttWNFGHM2Rp57Y2KtHTiM56/usJVap8QO8yvOsZYAmndW9FMcCUPB
`protect END_PROTECTED
