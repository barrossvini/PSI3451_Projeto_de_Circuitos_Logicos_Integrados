`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LPweWs1s+MEn7l0MOkQNSEN0H2RPo3pQrvDskNqXIEwGDu9aPYftRvlAPpz99vLt
q8usMZenaVczaWPSF7FcfWxB+C31ostRiRoQfMLARdsoDlJk/BnnvJl1NalNFDhx
u47R+LVoi3rAAp+CoKgBjItcBMcaxdIc42QDnWLVgFz2iOJuRLS5TdgV5H2iuZPl
fLLTM1evntstU9AR8KUrIhmazJtvgd68jSn5GPtNF6rl6+OKKGHJnrwsFPiFm904
0Qcw5QOTkl98XCkc5bcfDoI73n23N7HG/dOrka7OjvHuuWZ3P9wqf4IRBJ8Vy2uw
IZJ5tcUSjW5sox4sGujkdMxLqmZWpCHj19nTudtft7pcrGLJS9KjYWoofiCQs2DK
GQKbVCkVnBw4NLZG2p+gGsQSZ2xhjhf0pjtTMn+3zArLArDjIqY9zhRFXE1acwnn
5Ypm4pwfX9B/4oNEWCI+fqt9k/xvJd/yIIQE7+A/HeGVHw/5CxZpdeFcUEKUAlWI
+/zTjry+fbsV0qMXK3sn0lU6m+mZKLKGfY823b53H/5YvecqLV974/rTJ3O0Cj3r
vIaaU6jjlrQ26VJC45aPAe18SmiVYtvOd2dqA/4F3RMkUMBCnNiSVpfq0SfCLfsb
rDVXyRovXd6ikixjlKngAyYOG3hBeGEFyMM3SmlNKxm9kRar1gfLLFvmuvnjmDXk
iPje9K9JJTRfxOMeTbX5FWQGmw2fA1JDcB6TQ8sAN1znCXg4GareNhFKtHLh1mPf
Pl8Ezivvvt3Qa4XkM0KafH8deresS3P+6FZ0DHP3/BiTu2Upb5BKW60OgNeBjOCO
aW1aNEGB4h5WlWGaVTcyiQZ6Y5yyQTgJp0y9ia3Yn4qkO2gcT3uqPgZnu9eYGVsn
F7AQoFfBKv5AKm6esI+NkBqYJIft2LAzaCC70c0oIhrMR80dsef1j4J+elUfszjU
mBdDuTHR1ZaC9BWpfwqcI6jb3BIGGdcxq5yyQgHBSCpSRGqh9fR5e1X0aO32mU5S
M89rbuOH1sGUaNpwZDmmBrpI1OORPZwb7Q4y6E3Roroaxz/15SqbJ6PPbnrlCTmf
o04AW5AQWVr2trFo/lD62IvE+96bbxsLDTxEU211oQxEZeId/wKpgYbn0YzcPv18
co9Ys9vS+T2LGdhHKqfL+FQ/ERJ+L3ebI5PP36fST/rpDFoW2n2dIa0UHvkEKWIY
XoCHQCsSPtVO2LNz0iae8Dv0X5TWV6XgcYtbA9nAN2vMnhuVqx0e46fwvb2op+wf
4BMpcxjUGy+1CQJokEE7CclB7qXywAkPgrLTgAUCK7nvKW8gwAPJJunjX/BYmGRU
6tuCf/LcTlbTkzvCLnBoFgANzDDzV/OHqnyXv+NaXYTYPJ60cvqbzcLhRMx+9lz7
00BEyO52lqshOp/1thOnCPBjJqlBysl4AA+g2jc11rB9NCcesGVp3im+NdTwZRwy
sjj+DcehkUH0cNd4Se/YqUHk82A/8GUB0AhGpQN2lHDf7Ro4BideHVVUApQcNNsX
j3wamY3yOCCHJW9OJVlnFjd60tcG1bdAtVI+hAfZGSnGow3e/l26+EYAKX5WAboN
XC7OjZo8evo7ruP/Kyea0qSIJOiMfihDysCFl1XB0yYR5oERThVJAEWMNYaTR6c2
7QBY3DS8agydmAAaah5xTXPMSV/mNwaPamWlb1U0pul9O/y6mXXCShZdmzjwPoqp
70Ru2SOmkytZ4sw49tEiAKuGldiJ0tkeVFTrae18QoM2RpcU3qtr2heuWjU6dJDc
FdE9TAuk/axsd4zZ8mwKhAhF93VWkbs4DakX8+Hj/PMO38Ngv00A60o4npyvkTjS
jJiqqPnSnvrmvRaR0RaLwihLJ3wLUyN4Fi9Uf7iguIClMpUjf+EdeIdc/b4Qdwgf
P38MBpwNZxxTRf0/T8GoAmlxPzbAragCHdpC3IoSxm51y6AHVquPJYc3MT1hwsuN
j0TPU7rdNkgwM47vN4noyMdskTjCuEARNBDui2wIOl/XFtfeK4OYD16pJ7ZTMT2N
lI+zRZ/MPJb0Ft7jn2tacLbqHZOSJAJtF3e5TiBbq0+25pa4FqZ9LwVebLMpqBNU
8S7AIEkZlmtqXv964SYdBXE5rP527yA/gEeLFK/TyiInttqi56RzjNTTgwp15ljG
M/hYBeP1zyyqMp2yRaSw8zewK6cAKgVATU8cAwNtnckuvDakEv5mfkMbhEjzNtx4
fR2twEdck8DMlZIeg3SyqJoOgfT39E9aLjFd7pFnoOesw9V4DvlpP/xFlgMRtoVJ
t5z6j9IT9/DLBuxE94X9GYN1ACIQ+olfeDCOzKSe2eNJRNwSM2ypwCwe/Onm2frA
KGQeihpiQo0ldMR2KeoWiflB4w7tlvhDLn2G0qu7kvIPI9ibDWtmyFk3G8oWuSYy
/DJzQaODjxKqjYpdHGU75CoG6F7kgm6WRCCA+JJP7KNOp/N10F+Gsg4qZCmlbGE3
2narw0+4qhlMIFU3Zntq2tpZ0G0CNdnqH56zn37uBiXq5QG+CLHwtyPZCXmvHGqk
X+b2bhHr/eQLVWDAZXCJ33ZeLSuJKqUFTbXsJ47OqcqibMrclXbMkA95MrjhdFKo
OwS4ga9Ar+b5o47aofK4gVYzJVs4XcnyUqsK1Y8ne/HKse1s9f81nPCScznaBdKx
+7R6GmSmf6Zsr9HscZDl++a3rUqBTfYJdzqBqUHhtBbCQC4JwopPi9S9x5mCZkZe
hD8iYPvhzcSUVUk4klPU3hDN1QbA6VCdPu264PVeUa4hbR7dQ+ebeEAt2zoDx6wK
mCSnsHOSNPMxnRBWhwvnLowZvo3lwMflCYShJLWUaWAPmNoFa/q66SYmIz+hxlvz
Z3awVzBQuGWfXsp3m3Q8UvQSLTZPek8P7mm+5GDwuLxWG2WFuijMIflfEWS5IDwU
fi9kqr1ug9dASe8Za9K2QK3h1Tm7jWrjhb0eikSF4Pn5HPuJj4o51JxVpb+e6Mx9
A/yzW0fmrfdgDSVEwN5rE4Hlf8WLGZgTnuLbcCc0EdwFrHwArOOvql+aAUMBPMQq
TEfA4dFZuMy4b4WF0Xk9jt18ZeCVFirGMIaQAv7MwCKeAkvjt61LGqnmG3l8s0KY
+MJFCSg4kP4ci7RTEeOk1a3TrO2CMcisiBD897lhAQBc00s6XsTF2BO5CSZapFq5
FK0DnPWT+MXKpZMKD8NLHomqjb6yEQzcSIGv1uypUyw0dHbCKYLMMo45lyw8xcdi
wab0YJ0sTxYvECBk3fhASHytANNDsjH2H8lIWQYEfRTHgEHDMlXYsQ8mJZucPnEr
gbYe07LajBJuGAge6kp02zxUEyd5BpF7HNfnBHp0F5LJMTXEOn94ERRQDPde3wgC
f5kSCk3tM3tDcKxDRTERHtJzFVbotheqTRbB7h2tm3XxbxkpN7SRBBXYd9Yk7niZ
ECMfHwO1M5x2a0b7rZjede4wBIoZI45NUkTuvY8J73Rb7O+fEe8dAXBrJ1B8wg/G
qBai/cuKl0B4ZO9Zz4LXmV6XGnXHAUJ1vbwdYiV8X7mvK2RXBYVKh3MtaiMZDfcr
qaqrzeIKaZ1boXO3n6ZKEg9NqIDuCCFkhQlf3HPDQZizdYU6NrSGjNCK3t9SHN2U
C/CNLN1mkPmILvWGXie0gHLyDVyAbFB/C9cO93ezljSCQzUF7OUedDsZwDiSqvNV
1w4SIJPtkRmm56WD2ZdBlgFWxnlLEWNRP75Vhti5aU3VElQSazT8Pj3bOGjlaqMY
rIN2uma1ogbQnGbFu3hWr+WoTheeNok+UEtd1TYwR++fP5QqN7iCQDSGD4UXz14X
4S3d0r7/zN5n60sl174nqDnG6IoF4oCZEGzUYzn9WUqFmaOZ3ViteoZ6nFjwmOU8
2fwE3zRUDWbDLcgqaJx1NKQMNztOKaQ7qzIEc0NT1qNmDKO7ZElSe/vkfkkU6Dzq
MNYJOle+wKl2aGUgQng0wpaIGdFp6+pzTOxYXievoxnCu5pGhYMoa2WTh3pan1XQ
1XUojGciMPpZBXod49vHsxr/Nq/9ptQfcyjhqSjMZ0Aei5qeEpMFBiH28ks6qsxl
UkLeSUqv08XgDBJcRWoRw1RDz02jw8LyfG0dMd56SDcY6CJl0Z445FZjhAFqoKtM
iyrmnRx6rzCajBgUlki1xOGlCnJqwZ3mUeH/oRbW5prn+Mn26S3uStBptJ+BlJa3
QP5njUT09od8Z3/MP/AVrFRk88OX2SzLbHNuQ/zx0GLC/+JfThsF35AroXwgKlII
v6tcTJt2TrYrD5w+bxSWhgFDLfzE4HdY26eoMAIW9UCCVEwLKBk5ySRqR0SJU0Gg
MseLhqYyQm1XGmqrFL9l+P+VvhzWEAv84cyf0kDxW1aemjX9f08F7N8IEI55BMvh
kUIkd0krfUsYt9/SAJNqz4Sxs+lpEuHdUIphR2H5VwdrDTQkzTUolJkuJc6G+hwg
2G59PsC4cMj2G2D1NM3Y03ffFklR0+CY7HINenBpOe4BCZfVH4OPeaKSg6x8JQay
BxA6aPu7MEBAAeijRoFaNqiW622wtQC1o6DXmW5JmOyJjMsuFCerL6EA+i3O1KRi
2HOKUp6lETSDXmyTDqQiO1E+rZpzfg8IzBRjYlgohjw/Jhk7hiBG9NO5EeOiYfii
M075uhskqmKMETaxIWS7TG2SH+KdG7xnb8KgqSV6EOQ2gaERd54L9UL/5HrhWcrj
R5ImLh6oavc+8ZS5UczBBxlF4sHeAefclWZiFbqvS8dw/MVNonr/cek93Bsx2otI
XxVvxayDHe0L1u0bslntN5/Tlx17Qh3F6O5XNadlhD4z+42YZ1iV+ZyjktWDo/7B
jCIod/Oyant8nYjohRO07CKhR4qdaUjrcF93hmm0tihQSMrb230kwqpyklVx+D42
P+G3JEwmzeN5dQrpZYt1C81A0DMUiSEYoRjYhtSEKhp+ObQbaQu7jyeww+xH3BEg
lTakhRAUBadOL20wgzTv+lfmoF0MRKISoo6kbJ4vRA29qcc1Z0ZTsO9MTsw+TTfN
g2bqUVjhiIPWQ5FZbME1NtnYP2dta8ePAqingSMipnN+/OZY3EltfnPctkyrUErm
YC/kCnHqo+v0s/qe/NNBTk655PSA97LqBeuo5yLGspzqARZ/R/PycmDkqamvAo1r
gCnbrgtxxJ5dh0yWB3EfszLKKbfoKJPHyjC2dFBaFAcuEX+dtN6MzWmpedAMjNAc
Yqb7YbP/GOqNngTLq+MoTw==
`protect END_PROTECTED
