`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JV9xHJxfZtloCqPbspH4GFUPl53cCfYvALn+Col0c7EEIG4tfz8oSTUgq8Eeevz+
0xRQ/37qoH5J6l4Rl9u7pytlgS+r0OGtAcWUTyHYGDtwLtQ+3UPpB1trPJBJO6AF
l6Xoj/hMKg7Q5JsF1n89z4iWuN0wvq5RXnj2YAA+ac/XCDv4htQAkMI4gObniMjP
6ZlE8og79XabDRmCU5P1rla1doB9ugs0i5vly32Ouh4ZJNTDIBqkaq3BIWtT4ElN
4VdupYZOJbZyo/CxA5BevA==
`protect END_PROTECTED
