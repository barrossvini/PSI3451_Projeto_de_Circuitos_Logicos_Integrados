`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lX6gc2xLICmFyd88s3nVnJ3IeBQ55ZxSMLQHHlmFkVPjzTv2HAM3PDFjQa0Hh9PX
krJokRn8RXhFgBi8LzKue1IVt0P53FIOc/s48sgYNQFcdLCejqKkNuFVbtfc1uAd
KL6IjBMfaXiwVaOd/MIUzP+6jCtBukkH5l6+Jimc1d3BAQoYroPI8/gN9UibcPHm
W7srt/7nppzg5KLHL5bg4g==
`protect END_PROTECTED
