`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/X4WyG3ZO0MrawL9IhHrRHJqYULozdovqPD+1BUgFJzTvvwE0R/Qfux7q8M8jY//
KHp8tIsj1+IC2QOvM7/CZJPMISWPMvllsVBEOJR10KrP02XlklNuCexak82p1an8
gOnbZn27x6k20rDLRGgVwPe5eqOpMncUPgNVrpH+bdRgYALmcm1NC0Aftpp7R7Dg
27v+ooQAUH24unzPAdsq878Rcd9raWezKLrBGgyApB1lwp4EkNm+vZmXxZIP18Vm
h45hBEhBVZDebJB4dDQiW15uMegBzjSbzuIPZkkhkKv6Ya0jlEa6EN74HGr+4clB
LKtICuCrUUGHGW2lTtmXcJf5Y6F8Fi0OJeKzPMInQJSmwmys8elNOTrqqhLUUTtG
ft3o8SNc68fOKGBIrykgd3dcMDL7NDHUtgL46vvr2wV4RrLdMCvKkaJn+2kfk2Hv
qCurxHfbGOL+5f/qoo996uBgoimGDek21g582GY9ZjnUvjAJ8dN/H/mOHnAPHpKu
n9blsulWBS3cqTcN9D3n8ZXCMWoLbkTmjpxjBISRaqLwqAyYkG7z2tQ1MIkqhdBw
+7uln6SoZ8MTtTTdTW6RLurHNgf10IPbr6Y33wnXokAT3WVEe5T4kJWZht2kwleF
80wgC8yaEK6p43cWrPbS2xihKESQfDzbP3bZsBlrAjXsflhnn+Wq/B2f6FRz2Hqf
ydbKtNq0tyQwOCbhE45xYBVbypkjI2dcpAnXvm0OQZF1zRwLumgB966jLa64ebBR
EQUFbuMEVu+M1HxvkQB9EpAoWTVkN1fKI18dQgyt+pe/2CoTy6afSbQpIKvWWXPa
+wkvPuMjQzyv21+lqbFh4fFlXRAly2+yuzyfXnio3Z3XdY7sG/4mpUvi0zN3Nz3t
mZ1b4nR/bxmml8d4nZ+0UV3KSJ106gIp68/GNrTVMLUUPvv7SgLtxKSAz1+gJW7H
vJlQTFMYLC97h6GdSH0iNcvjuGIOiqNPmZ6amiGeTyFwinQZtHllf5Qm4InEYYzw
oJEWleWEZAPlIbUiBx2TQnjqOiXuRkqZO/uvlUwS8fpe8e+3jVUTU3ilyfr2/Q9V
yrrwzPiKqxTzYyViX4g+K6B1hy+v8Xs0VOKyL1Tb1NtKhTiad7ESnnH/WglykkiH
mBSP6Di9CYAbW4nt/1y7XjfhJTO0wvppSSvpZqmaKN0ZpFrTmOfRAdmDIBqBAf2j
jSmP3lQ0kkADmXrfRUW47WHQdId0qP7KZjDihNa72DMuxds7NYJWu76gBro7g3vv
8u4Mv3byn2s//0NSMKIDaIlSLsvyWufwDCg0ns6CQVbQRjaY7/qe45sv7RrxATdx
tr+1yW7TAtVldyq8e4ZZbdJJVnhRhp//RYMcskjVmDDlqz09k8vTxa0ybnOHPNdu
NnkzmxUoY3lA1BZER6+9gAewrJ8WgNEha2mYOUr7DlxgKlvimasnrPjUNWKwrk4h
dWkqrMYqhUOlVaZV4S8F36kk+d129DOm0DHdUQ66e8WGW6ukj/dgFP+aEtn4cuGZ
SiqkODOoCm9cRR75V55O7mYiTjcBpcZkf9s+WU+YJyCPi6u/lAu6wsUI8jVnqKPC
p867O2YF9OADGkDgXag2146kX7kXx51OxHmhHJe0uU5lkHNYIOwbZKvz2uk53tmv
XNvZdXnZcWQjm+szA52umpcx1Ssgzjet6mbh4mBDjIoDBXCLUQDrvyM28BiUrqqm
R3RkpTlAuQrqYGk2ep43YZAn8J0nicmPvDh6ygu2AFVOayY57Yoa2Pl4/i3r8Keb
gb5/UKFsdMaDEy3lB5gI1ilZewkcn/H/JkuI1hf9Zj3VChpGVJsK2ODvHlHZCbG0
mAgKkVRyPLqmLg4yPsi3ynhdAuu8K37hg8aAEvzHlTFonn0hnTmZtgvR6SXrLRMg
TL5rRKagSXbc1mu5aaRjTHjPf9zxxc2NbgZU2cn03IK49m088RpkbYRiP+yg3kS1
CqZtpJKbuFA+ZclYC+on0C7/RuzEky8td5mt+bhQi7rVTgPqE0dJcPkgo9T6xr7t
JyOwE/gIJpN+iEzM0qPG7iMY7AJ6rh4vnueSky2nHOvPemhRfFxVrwt+i/3uzScu
L5ztITmPRVwVNDXCUB+3Evex0WOGoKJ7mnVNRZZfSOTs4guUyZ4MhwjOukkKo25/
ekUFUg4k07mAy81E0VLkSLBubYqO8xYkIzMNyK3KJSk27wHMQh34f4LpYgqVlaxz
fwt0TakQp646A/pT4psje2zmNzO+MFeMUN3/aB2BxNTYD8eugWIHn3xUwAL02HJj
Q35xYHh6ubs3aN469Oszi2T6XOenArMIAGazucgLZqFm8+kaLBhHFrb9A2r4hqa1
XaqsRtorribgctuueuvt6l2fI7BYg/qlEz6s89lqpbABIFnfwlUksn3f4ywSNLjf
vGRatMGlovgF4AZql4lIveRYWRu5//yvQUrh2p4dJz7oIRcLBzmPvNSAWpRPDxk/
gwVpbNfbwXN6QnijPmAuxA==
`protect END_PROTECTED
