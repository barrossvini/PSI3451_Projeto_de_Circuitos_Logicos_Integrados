`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+u3pqqwsGr+erj6UgC/HtQp1cucAkT5jHfx6wO6T+Xc/g4YT7v222dbv/I6ZL8FV
VOunljitaupwBDniwszvde123iMPjX9liP0JuSp2NJch9C0qRwycN4+tB27f3YnK
H0kfInN3dHIR2r4TioAh9AkCe8zaMrR6Uzj+sXtuDGsHM3mx9yMYPGhr9c9NXQeM
+ezR2frPMeu2Qo9rU2nB9GQKv/f7qvWVY5uTD/Q0A/icP/n6c9hCMZlMS5Tt5gvh
uPQMtZukcH8HpbXTexatDK5FAxpa84D2YG7e3H5ZffPCUuDxqoNY3gMd5zrFtomT
WkDA1Pw5xEF+EzWlYAMqbODKX18cD+yqx5FSSIf+UFWLYGQOCBOPrgQ3k7/jNfzy
iK0Zoq/cOOMcfYxra+JTz54/u6N5P21NFqjJjVLiZ1JHvWw8KrWg4qcMeyUi6tmf
uovKquA+TZgji3DnKAnUBmmYBt2ITkVJX78SBo956WAMJQsrxRwK88GVgwfn/Nld
Zy8Lq6SbRdzy03QlXwlDPS3+gFK+LH90fFwQVcpWgyx9fh+QgU8BG5UiaakM+vOq
ukC8EsQICtoQV7xsAizWIW9HpvyO/oXG74TFx4CBennLnXBh4xrhhSAaw6n1/Wdm
17QXvvHzsEwSBohylvPnzg7T2rr1qz5i+NK+cnunixpCR8SL14LiM0l6xAj0+ztz
rQxKzf2YA2IHQExalHn2N8e1qU5Zc0FBtX2FjayGP+d1XzgjIgE5CDPGtr80zRKH
KKgFtSXNa5LJ/vshsR+7u0DtCDAX71yTnz801pd6OpoTUyX6zDgT8gTpRCPrHHuJ
rkLQnRpAEXDVBrn7r88FYxHbVFtJTeLnxGxyzOm/pPvxPWDHsDE8xy89TKt1+v/V
xXtgbCipZHqVr+74JJBo9TkwxAaM2JzFERButJcy/yGcGysDvsK6HZlnoaqs67Fb
1qGEQJ0Ui4WFmsVwTv9azuT03w2rheV+qPKcznrcyIAaD0v6rjs2Z2JnnFQfEEOm
kvD6eoBtKITGtOoMGqNiKzTrrnTcXyK7EiHKrLb+Lr/n7dyJid78LTGbhIzqdR+2
J48IYNFM7jRIWocqkq69qn/cKOt3Z+izC66odbTbhl0VhassdD7H7NP9BqgT5nf8
ex8GdPk6ZAqyw9z3ZooGcmgaApFAkmyXxHqZfG8il3RZTvm56lQ/c+4YnnScU1Si
VOYdJ8EzN65BKDphIDMZNxTwqXGFthB1jDgS3aRaeSxLDI0+0Cdc5q6Mk43R5bw6
YmyKYHTxnCcLC4F7nr9gaB1qvu5ynCpfglHbpXowjrFMl/1VY0KV8lrrMkFAS9Kx
J/pgctbpGDDMEQAaZv6hys5R/lK3XW+5N5eTd3uoFjI=
`protect END_PROTECTED
