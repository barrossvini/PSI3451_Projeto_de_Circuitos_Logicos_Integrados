`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zWzRyWgEmrXWh2+yAatESk4ltiuOUwa9/au/KRsyblHw1Raz52RyVEZnIgMpEw3Z
oZ7BGNlbNgfa1PopHOPp4j+UlchPFs3NgYiYmSNxb9j5H2Yzp0eGjtilOD7YDGHR
FvCIzH6Y9Wbs9sokK0C2kT8pyJpGss8jOIqPrjcSjDr7BEjE0r/V+Dr1jkNFVrYb
l9VUpnlK0VlRq8+FIJ/i4yJW+bE1N903V4HLisF5ICeyavtAkaAbY1DeJPfEYxNG
wkPheMM6gUorMMc0u2erUNVWp/aE5cWjmqpWHgDXn9bZ1D2h14MMgBBcazLGdlOP
C6uJcv+bdsgzWh2PSaxmlirxILLO6YVfk1GaIhDXo4PLkCT8PQK2jISDzy8yjwRW
PTfVxysKiac5nH/uCgXn7W4+zDltlivqmTh7ZEp7/fS+FrNAlj8Jgja6qcs50RM2
RMt8b0uwNdH3VeWNnMDwvLIdjgBd2h5xVLy0zSzEO9SYTWrC/j7U5bnY2srrQ3n6
TGet/ZdJftFmd9cDuSU8voy1jY1hWoYq+/1DWak4aRpr3JTJlwMwFQYSnDAi1Xxw
rGyRGjiUpGyVZnj4lnEQds+NWDhwGEFIWFw6w/MuujVsWKNWYvab0coKNVL9E/Ev
z4C5ZtHYpqhxFiJwJkVEwEB+PhJCFiQloiHMhqItv1hV7wace7gN5UaJTibWhG7a
C8/rlvhjtDmf0ElhzNRYvS8BpvRXr9c+ZLv/nLj76uAtjc3RS+5y2alHn6MssQqX
QmgzAitdAq0UFKeoun7fBVZMj2ue9MugGgfUF5/FXnoHoc3TIVcSDISddys6taR2
Wa07GHabYMTaAoAC30KWbj4WscMwhyHskZpwAWFY7D/X6chv+9dRUC35EDLu/xu6
Z1K1wc8ciyyGwvxWu0artMyN+Ys87ST6sXBaCIfy1hrN9/3WHtDZUN2taEg52u+b
9xt/3BDGSluzXP8k2E7RgfNGNt3MpY0j0VBhWYr94gbmU+Bs70FvXjKAJNPxtPlQ
cchVH8Q38JduzNrRP5l2PD5e+f6En90DNhk/0FdWHE/iYLuXAnxh5w0cXEMAjkVj
bTh1GUfyO0c/zvQAZKohaxdfPAF2ichW/3exK88f9PE+QzBLiUpfFgps/sOWcbxQ
4zMG+YySI9kZt3xTfT8Y43x7/rzkjUHAWiBI0Cl7ps6K2UN9N4v2TCG9HlCPGNvt
GQkiwwK8tIDaIUNCpShONA==
`protect END_PROTECTED
