`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JE4EAbZK04QMO5R0lf9rdkxWzPIAHYboPilqquvPnprWq3H6L/KzA/2JhnbQt68a
d5gflFm96NTskG0gzT4d4VahiorwzxziDb2UKR9rJnh1fKvBg1osbDF/Go7Vf6+e
UspEd07jdClMHz4fqASk+O7ywm4ZNgOKYOXho0CYL0fbQ7ulwj3Hatzqg9psdMLf
W2YgmeR1QwtqoGQsKGIuogn1LZUlIxzftxfsnfmSxsZxrtCV0D8RZ2QZcDrTVwr0
O7zRCb8ffyrnMXARkLaVe8HPJ6gSrqLuCzHGkobAaxSg18djGo+O01OGEf397YmU
aNW9JwEe+zkKmn5+VGpd6DHRUvuj8CxfKQH/SmRzM+05el894swUOZq3ifnKe7dO
qk0H1uTtSwmedRQKhhBmPRffdzWEgu4AA+dL45GfQI4I+MCGD+97zsqcR9ouPb6r
VVQLw7HTMAIyjfz5P/6CwXuHUrbpsjR0wi9EK5nsg4L/nbscmW3nTEpKXC8+WcCS
jDvS5CKZ60LgJCIzFvWntcUvI1BtgfdiblxJ4KOcWh/okZdo2BJp7fDbN3PV1q4g
d39dPktCd+bMnLSVUu41ONeiuC9iN7920anNmA5QBB3Sh1iAgBDMyQV6DMEZyXqF
if/zmoJfl4+m3nT2Q+SF2qj0Sr8dPSaJPAoDZ3XJBjw1n2THrF4UutRMi3G9IYFd
4oGhtqhhElzBH9x3Ew6XQB66hvg8Popdp2vKyX5ZEqT548iqMcTW0jyEg6klQQw4
Pvg4f0IEbWc7bySwavyY1obkf3m6Ro5xgI6EogiQnLalOf2wGmnX2LeK2/RY49l8
w6OWmlYAjydCxBaS1copOfVZ4776RG0XA2quXtQLTS60C5a//LZghfx5BKpLpxaF
dr9SQmKgE2tZV+FQXto4R1GrlHu3/l4KhLfMoitOmr8Wr9RwCcWbktgckVx5mXr2
uG5m1EgyMbkOovyfvs2/NqrjbCx2qOwigCUX0TNjeneQm0KJlJAZh10r7rxmNjlf
LOdyolbCV40EosULkNbzQA==
`protect END_PROTECTED
