`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5poRiV2BkI4UAj4eja26U/Ex9hM+DxUC3xGTdFqUNvJ4+Fux3htbjplKTw/4hmfZ
8OeWuw853k72KKDZJMQv0Bi1mW2sephB10cM1yihqJreSVsAujwWgqLtyYBaeF+5
yyj42guBl7ISord2HXO/tSsvqMWXCzhzS5r4kA0jKP6+Xtm/Vf0rs1wv4dqjwjNJ
beI1n5rXgXypgJwHtaqMsJnlr05IJdv/mwwnRGztnazoBfE09RsF34COkcWx58bO
rcKTry2X21EVW0CIxyONOqXfCZ7qkpDUKhCDLuucFcs2JeVAOzAggZfQQ7JRCk61
Nz5X2PT/3EXfMXXDIdqZY+9G7PUrxAFSZhsOkA7Nd+Kjt2exgwjkRtkNTwbjkGpb
CpGVKIyx1Pyx63C3NDeGro31Pw5tkPuG2N5JFi8NDsfTlhpVS9cQJSYUqtV/uMHE
FetMfXWXDC4xR2HswxcyFyBOz4WWZtm3YvoL8h3BvicODuZ8Cmkoj3f4/SQ2UG2v
xpUhp4vyHfxoG59iHuzGuvhm1li67QRQJ5h9dfB1JPDHUd4CIRdz+zBkEKNZPSVs
rVzjWArdTXwkdbZzJT0ELbNu5/A6i+JL0Wk7U+uv0eVea0ZpKmXSkNPnNMfbFAj4
byMDIlUUW6tGqsjDy1KzMTfg0cb0bP+b/9lY7gFnoPd/edb9299nsExjNiu1/YUY
G0x0ULN7E9QraEqSHRQX8Mv+9aMEy5rAD3Ydgv2oPe7XU7uwV/QBgqJPNAkEy4Oo
0mFbv/et5NR/PASQ/Qv5d+77bw57JpiiJ5hJr/0v/ey/J5E9BXu7bSl31nP+nQTz
OmUvNE/UnijlkLluegojStKVttS2TTIoeRimX8Rwpf1JqM3ZtkoZXyE0JMlbKOyx
Hxwy9+7OsKivcEn6B6zF6cOrKPbqNaVH3Lze8ze77i5Y1yZ7aepjwu2H8AG6D5OQ
5yWe5k5s3PmQo/B5JsSwYh3Oeeg+yqRc1ZmN/UZpedVvRWZK1H4SGYxlS6UDsR6i
JPRsO5d2+vjx8VZpXx6q7tZWwR/FWBfJVVuY/DUMUxThNdL0fhV1uUNgSgQTqxAd
IxEJtmKoSHizesMtwFN5zOGFd62DdqOh7nfO2p2Bmee+PtL5iGFuzMx+WPYYeX8M
EZZaLpbeTpujv98ByUjyMIy5LF8bios95Cxglq/om3NKeWie0ZGdlXCaj7VVhWOR
cc14a8PN332+sxrCntM04jhEHIdRiWiE3t8KjvwNKOUYs3DnXGiVkjNqIf3J6sXq
3bAQLJVBXbw2Ayv7mijpE4NeVJW2PJ9WRlCHUXqa0lXdmKN1fhUxHsi+39XzPLo6
kxppNq+V0Z4EIDJqMa/RIQ/GAANYA/+ZIAyb3wJsJcX1aoRPUs30I/a90h3L77U6
WNkrFc9suCfDKNfxbQuZd1XyS1L49yIzuPbXo6JBvfZs5dVGgz5fTbV6lCPLcvZ3
otIElc8HOqnOaiPpt5H8CdFLSfp+Cq6KJ2/x17Zjo+Rmt+ki4K+rJpk1LV7FRlS1
`protect END_PROTECTED
