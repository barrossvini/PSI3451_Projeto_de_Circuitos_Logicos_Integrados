`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
80x85PkrFkUtkQATT0daVGv3QNE6nX0adtR4pPbtI0W7t6xcArtJ+kCZpOn2ELjD
/mmYl1EjmCUsinHtqecbukcAVSWoEnd/+mPaLV7RGSqY0E3ulL6gu1Y1RH164JM+
DPy5J3DNNuO5gnPbLqn9d8ibFUe2ik8NrvdbkkpZO1GQr6nSnqw0gk1BpgllITIP
aGT+f2ZeXWocVaPKaut24uP/c3eVoo8ZTcVgf5SOoGYkvcTMnpGf3vkCRh0qezMi
hEWq4jRfIDckHiahKVB/6l13zU/JP7665Fqn2ppGK03zO3hs3bjSC2VzZ0JW0OxG
OTKh3PMR0TuXjfydGqGWOxO3Se5CNVPj/Y2qkKV1YvlOzG6Ncfh6VTy54bEx0rfq
dmTuJB9mPW/SJXcZoTkwPXRWjFjQhg+ckkogkiZ5SBaUTuKM1Ex6b/hqCQ4ZvyRI
vIYP7bBvHz9QGEx9/nPzdY1mXs2p71jxIiNALMfsCSWxHq+4KNcYNNpE5t60G1Er
UJztXY840XjCSp5LN/KHx/Hz04iExbbhyXvWGVSOay0SddT5k6TSJL22be3/ytxy
kVN3B/OilajkdiIwonTBXXMgYOaMWaJgB29L8U4BDFCFKlyKc89QiQLNAYX9UbVD
HmUP+OZ9yH2qZb/qivcfqlpw2W/FJn90abPq2lRQkFnF2+gZaeuuVuFHNnvnlnn5
siEqysb1MyxtuDZfh1ZRnA8QqqoUoGRNX/kI8NJW2dL9YaJ6ZNqGiwgGpXWcwbAo
RZ/bRrOuKTDsoiOO1GqRI+HzdS0I/GDqk16MbgolcJUU1pBksRznfXmGsD+ne5Km
lwRCQHh/NgqkYfqK/+2k5b6LgLOMApyAIMaRySKMpDEFghekgh7AgNnkOpyrehzK
YBP4UuzBGETDwP5FCY83PExNnJrI3g9RyJ0727me5YY37BpNYDOfLyyvDGwjolzZ
8nZhkbWGwUpdYitRQvB7fkjzn+EW2ueJcHCI+TuusNHeHajzVwWdo8SjrFxldeY+
TnzdayVwtnBDb/AgndtW0gWXnpEk+hyfmUNdrS0WO2sV21VJyK0dCaP2jHrmcmn2
affM9247svDFf71PgtPnlvSECDz+9MiGzlTvU6wE/KJVEppjFdJgIAjI6LZy8e5o
Ka29acheGJlGeiubUX4nUcPLDMorI+n16Amy2C1HZvPTqGgtMHqPGBG6C34O9M8p
WLUFLQxioMJS7PyMNJKBMWzOZB9bkhk1882jq0Ysc1GtBZLj4s5RaC6xGQyJ3i8x
uiR7wh4043pdm0vlvDVTYcAIQCf99hkZBAyBH8KNpIjalZbB5GdJvRJY/y0v8Nkl
lric3lL37LKq0KkbWuTxkik5uuiQx+u9nRjLp02LINCBKCJe84/jC8aM9SHzmPR8
E4erjMONhA1ZCuejNJHMGeU10tZ5Ju2m6U+BLQSNw/l/zfpRiLctFxHAKzFUn3Qo
J3VnL73WVbR62AwYo+x7Ir96q6w037W4UN53lZ1WJM/W65RaNcZ2gjYMqQSLOw7t
8iPlgdz3XSu8KrsiO0sT8Jt1K8s8UgATcvxn0+s4yDkUsYQ2iaoy81WnqiHg+h8E
o3YbAAHMMaeZBHo8XbRKEm7TtQ5O5ug2PJrIKGYUdIKJR6xBJnf50GItJTQRpKBq
Y59feSuEEXWgpU5dJQPqSr7BYXQpegFADyrfkmop21vgEmrOI1To3C1OqpuJVeLf
iGvio1ZOkNE3EDt7SuQcFaeCv2hMaiLr64aGa6r0yC20oxOGqxZXidJZ9i2tqwZf
XtUtv9+RGR3MkEpq/dMi8wconSTzQyFY9e/MSNGs+YPvAxABh9Byop7Pqgj5YsIp
RRVA+NqSlVqAZTOkYbWDE0m7IwliegAPXcKcFXExgCYK4TLN/BZ1ThukLZqh092K
CN9+FIHIs5gmPG9p5QP9ErVMQrI8B8k4hKq0RdEu1bboP4lxAL4ZGwznNhdzyvqm
u/ZdZccCDA7/X741JUZzk7hzaBUa6bZ4A+kmeg2083l7CtGBbBtEhEgYuE2FAUnj
ltW4iubGgOCg54M+Z0bqhx9ygxxe/V9fft7M88wuzn/2epQNvEhmAKOAvkmqv6AW
MFSAJfapnDdIGwez0RxXn2UVDCnLAMUSHycdFIcUhj160QuViNdTY8MdOgOBdQ+J
OZScSnxY7qulEcumRmcMP9lwQOzcOn4VxBfYayBmdAFPLPiqe6fHlBcEpV0PUfSw
w4QdCNidP9Rq/tLGlPYS6ntw8orVJ9OXZ8XNS1Ug1oSg1Fd5NW8TfInTAe2BXV7v
BefXd1fS4ZqjCxg+7xzFh7lKWKIfQVsZAN/XbBJ+vOYRf3tCdmuHgyS6iy/PyTnV
zXY64j1xo1VqfeFM0GTffquF63yk0XAL3K2d7bkbeO1IateBtHyPCfPMkdtx5DtI
g/VOFw8VsqYjU6YhS+y/VWxS/BompT31gm94h886uczHVpDY3C6CUIHyyt0SaKlA
IA6OcbruPWz7WFLZnVc22FRvn0bT8nvdFVOpEU15sucbA2Slv8IZeJ5d0ivVNOwU
4OiV5PZZByNkJcntlMxLjhld7tr1ijdKJNoZ07CzfVtjd1w6NuvNog3UwccCNI45
0UbDrARYdzDeD+y8spS6rIIIXk1mtRNibTaTyg6YtBMCa2MrDf/dyDF7PQvZtD0Z
GX8x2eX+HGQE+hJ2ad8FmTPlwW00wVSQb/PKM6sjw1fwS6SPc1ImJZbon2zh3y7r
Ozhl8mn1iRga38zfq9SZbL9rNDDM2N0zpIN2Mk/tXCSyiEy1SMQCKMD41sZjrPZN
Ri47XQI/lWjoJBFfkII/9pN8rqDrrdj7UqMQClYSK3JpxpZTuqK3XYXMWyuVItat
kSxEgDNWTSqWniI742eInhI+zmo9KfjM4nhiA7NrgeJU12AvkZ+qKgtpZ3Va6xbH
dsYML3VTKCifhlnK9Z4B8obq5n4zjYWgZVcAqliG4u4rXJS6wqhWjicfDS5gk7oP
zd+9Dq+oKehbOkxAdgWVPp/5mpMooXW5I5XwAaIAAJYtzACf2TIF4bO8SQ6q7kop
mZaDda46oKptIv44ricuuE4qVQ8PZFbPTQEg0MIDvRy3JpktjJypSxnJV0Mjn1R4
5485GweGVU6Dz504EDEkxGb1+EXblb60zPs3rSKnDhRVp3Is8Lgw/Bag1jDcpZ6n
oQ/X1itFLFw/fWwYfkRpK/nyGS75tlyhZOY521474UQq1DNDqX+uVJMHuL7u0vh4
zZYJK30kqwkhNvhyTHUvBZ8eoUkQPJp8y07Xs5KIn4uOlp9EOKNeMXFGtYqvnKrl
+xnR/I+VBMtvmwIzUIuSN7vbIJP6xpJ205BgMa3IKklwG4Pf3iO1JLBlxApKcQLE
0RVzEPMxfk302GFAJXzfVZcVO/7qrNOWV94swjtPJyjClO9UDt5ZVNZAzBMrahQ0
NF+Qf0sBFdM5wygDftz/nGoO+K99TgMyRRVawVOSNr0CS0V2rR2S06xZn3qWO8ZA
JfOkhOD85j3/9w6O8Z3VDOPEyhoXZx1mBcYCqniuUH//ID2crWFg6ly7jM6QL+KT
G2D2fq6S6456b+ToHrprCYMaGH/kgbTgTyW7TMCWky19upRp07DbcAeDhtXh3hbl
GzZYvOdzOrPVyW/Khqaghe8cGt9zZiI3oiTAvW6jyZ13arPxagUeq08sPfKUmAU0
6grMIPckFo28CunJLvf0mSRf8NtJ+PmRFZJCh4mNX3tx+lxKGefos8Yiqfm8+0up
2P0prsF/dIp+voXw9OpRzZfo4Ihw85UqJE+IrnLopVI6IB2Kt4YoIgdAcyiyWIE2
h2YPSBlJeiDk/UZTIY4C0ESnMSkMZD9ivKGjfW9disXg672QlIBGStNUCvfFmEMw
NtOPZ5Z8IwH1iXtdSOYri6MTWAlBqPuzU4/VoJvQr28ZzQxqqaImtyNuybQBzeEk
BznYORxrUOpstbx1v5RZP8Xao/hdwocMaLzrr3N5VzLQNNEOkX0GmX4J1hFoaMgF
VfXy2TZaul2A69hZ+/YmsR9ppG1eC0kabNVjgdBGILJ1dklr6LTjGaH4r4Voa0M0
h+Siy8sh4LJuVB+0cqI2AEVGkNoo+7sRDtqQCDXT1g3BXrfG2YFwlo8Em07/jM4V
VJS6G7kD1MnZnYDxxomT/NMkk/ZhRFk3cHt0Yk9TLYDNTzLxN4bKKYCRz1Xabg+v
cBFpTgF+oyGLogHhBSeoSE4z9fH25i8x19gP0k0TZcDwfAWzUol+S1MCqjC/hBc5
HxLmJl3NalvIckDfxVJzrFMDJHmpO4X4iJwi33uhED5+7WMpy+9cqnoPK1wNZkP5
8WuRfhPLrSUbouCAjghjJnes+hPZr9QVrLcvkuDyab11Unoxw2RV7GaAxWiHfzTB
u2gnfWZnf6SOMIbwSaKgqnnNgfpuy1vZkU3AtYjgytdIPpRkoQVHAfcNOD4ztVXR
Qh2JuAu6rsh6uahUMk+vrdY9B8IG0gBpgf3F6YbLTjCaygJBuu0k84uyvpsEmXdN
KttdEe7g++BQw3nCEluWtkWSkiNBWYcws8dbXmj8AXqJQ3c6jTxsO6HwbYW/FjWC
LSA0vkbyfwQ0LVc3JL2R+KsTh7vrupoBBmN3JpPwrDY6iCO/OspuGxoK9crSn3DZ
jjyT/U8torHgfqI8Ux9eHw+NBKNyjaw1z9nlDHCEW+cLuNPiVIYE1nl6SUR/prqV
3tFEtEylIiG6NHqZ72RXFde7eeMn4+Wob2rqFMxLXXthnz7ReLrDckmypoML2KSc
OAbYGUbyloqrff5QZoB0RnThfvTUnLk7j+f9HNyxgfYourYQvk1ueEAP0scNJTKt
Kps5mrV+3Uixx5pu4u57z5/5pzmaLgQqe2MxZgOM/WqU6BLo625MpF9iXC+iYcFy
tW6kQMwfabmEkGjD9Y3c3MXZTdPuVxd038FEGhu1xq94UlecrdP12pjg6Q2t+R42
fGmPKQcq2Bpav2BpYY6G1fmXvuXNjbjEpeaeAsblBHNoNSCCVZ+fuaZoazsLhoUQ
BRBAfEVqAhI9mtUkm5EW3IFT7jET5t0lPjzdEi89zQxhAQVPs6CtoObb56UubtcF
H6be8CtLI26mK+s5efRd0sG0bYmTGjWMQZldvscEkfUoLQBgwobfwv/i991USfNR
xqDqZrjo3I+cchhs1t2CwgFsWfEBwJ7cmt5rqyYTVfqqZkKXZ+h3+iZ3v0XtUEgl
t2d2dDX+a5WCK9Yy6iruS6LNnt6QiWPUnp3rJY3uGsXPvdBfmXvosA8CyPXhqVEH
NfSZVMPcpbOyZG2lKpY0A8cAjXW6a40WBWMX51ezoq57e0WASsUvvPlHHmPqD2IK
sFnvhwzE+lZLK+JQ6nMiMqvFKJy/hbLnduC8CjyZVG3YAVJoe56+BxksCUB0vnkV
z0mbHglOGCHACU32IaITrXZTuzMs2vINpogSl2Qn/winlYwJnIfVNa9IYMLtB5AN
ShxGsDOdpvmEACMJyNTUexYtFRgmbxq/DPEdmMNfYLv5bYGB6M/qsF763K4h0WyJ
9x+aEi5gvPj5o9qVPgkBm0nagMyvlhWwXp+HUXKkButS7e3W4V2+q47sEtpSrc1U
miBxLtW1Pn6mzaVPpVin7r6s2rABE9M5phJLY/VDDG/Y3XBrueN+0xtVtt4LwTSz
osDDMh635Ozj6WAssOdwW7sQ7I+xBvOO9GcKAr/N0USQk9K3Q0Aqrgp6svnQl6vm
8XlqNAJgB7O6JU4gfcziWmV93XgrCMTsi9BPoHdB5jtcD4YpwjFEwFchZsqAGjmv
HvnT8ulCNviRutcrqzg2jIWbeyWpbDSjfV2sTy3YcLnes+fFoQSzgtFUoxHIc4YW
MBrS0yU0X11F77CrGOEfTXXzscYOjuzYURuoOFr+9Z0ig44gdfwR7KMAsfRdHf3H
lECfblA8WiWdEP8+rJ+4DWBncxMykoruGTgcoJIOPzQu8lC3aFv1HTYryDb1IbRY
ac+VuQZl7Bwc4oMBixccTCPRghOTmpqTvzdyTlT/fHHb+JKoD5WL11mMAK1tfL+H
0+HgNhg4AxBwfFld7t0XPFlY7e8HxMJ1WIN/1/JPW3HGTqd2AC4Yb7tWY5fK3caa
YD+qP3HNv9YnnCx+QSJ6+QtvK29Sw1pH4i234uHDGDwNJjqz125rbnT6CaVwutvJ
aIU7gaaDCOtS0JeADThl224Q4LzGDGiVpj3FY8zuUv8kIzopdfq8C+GGd/mXG3YC
Y6xmalN+V9VhNvRISghl499dsDUhKRHvM4WV4LGndLZVkuFr2II8nUO9mFBYx9gQ
+Kk4ayGeFqQd9OFTXlH+Gzp1XPQ5gtdXKvrJSc8QmYbKRCogF9DRFSPBiaQ6qZoq
QQ2VbVqzGiIX4pXxNPELFjtXhvLRWffAq7/BBku6a2gx64AHY/Cd1UxwqOzlYwYi
QPWV1RvPaXmyc11rAAXLNsWon9/+76HsppkEJxrtRE0VOmD3x1LID5Zk/SoyytSD
D41KgP2Lp66p28kg8cb85VNmYOHVWtFYBRYAi+jhFc9jPMWVf4QWLvMljAhmZW+Q
HjP1TLIUoUNdl8ttEsTMi2pv/u9NOTfePbw5qAIaeiymCej0kUcnRQ+UyF8KHGKY
jJy/EDH6chR7Pif9oaAzhBD5oopawtqImjKMbfFYCGanwxR4x9VwH1YXARnoE+Qt
FG56hMKOaBnOW4sE5RGN1bhdsw8pymaitnV2+BgQynDqiFks8NnJR7/C+kIVG+Ec
HZ8f91eF98M4FhUgmgSl71vhG8/PUpqWS4fqTSMngdpiQCPQJh6NrxzvnvAMCF8z
5Nqql/moBSdwW0vTlL/UDbYSqCZ29hsHN5HT94BiNisR4uKOEYZIQ7pTN4jNJ0Iy
gWohVD88g0AXhOH6dkw8T2Q9wZMpKBN1n/gjSYr3gFr5lO1kK10mh/XmFTH61RgJ
B4EhpAl29Mlm4nZxExjmxk6VOyFIdntLC+73S3JmFST72ACLfxuPvqkrpq8CjC9D
j4o7vXCGHUY1g08RTxBRSVwXtBvhnr9NHcbq/7BIcu73iYkoQCdYJUP2yh/TH91L
jVK97hMTDTz/xO4Ie/w0wco+f8KBkxPrFi4BouVa+vuaT5qp4LLLJ0CauupFfN/g
MCb9jREyXCRUCLgREmDIVRr/YxgTIf8F+3jupJC4v8C6JOI4hW4Q83vALnClXtff
PaSSSZezvFqrsuLn1xlBDI/IJyRQMvw6/LCK7KxCXKEmYlQ3SpNH1kt7kvED/bs2
BgTq/W/mhIf30EwnEvsnS3wVGIEbRmcCmVmseTQW1D4KofNwSlb/HDdlkRVpXpgT
FdkBgfPH8yRPj1rnmtJexobRQDFnb3X34ZJhf2zSmm2ADbnyXxMeKAxJLP1EJu74
NYGdI4sD6vn7j9ic/OoMFFts+vNLz2IX/EXsTkWdc7jfW8CWLa/+zaBnC3PJ9Ma5
cz9uPNgTeZTtDT+vr8aeFmRDh30UfrcfsahoAOfAEekPRvVhaM+j0+n7X7nd40j+
cLzOBh87BktRWoQEGgsBTz3jmU7Vlp6z0JlqNgDdCwq6LJfsdBP6fTIBe4puYsjp
WD9ewy4jFSJf2a4Zl7ZLHWsatEJWgqkeD7aiP4POi5eEe+Di7HirOizQGAzVTrZr
Rjos6Kc35X2nzuNpdIgCfNfrywekpKJmbKyZ21waT3zuk9VRngcHc/wzLFQG5eUH
4QXegHNQE0tm9n21ziLl7+ULWoCwDNLB9E0l1EZmi+lJAWFCGeti35pPcSbM30Kf
EpNkgA5n/pWM/cBiL8yWJ/uCyrpHo4pKXowP9OLhElAhPD8Se/j/ezL4Eb6Q1I1s
yiUU9MvJtioP4K3dzWiRStp70SWSI+AS8V0rhJHKN0ZfG0NB8Cvmn3o5DY7E3bPF
2qxfkedaAXwfuYlm3+DDqFBIAzFYXQR3NKWOpyPlN4FmGDZddkNXlsftXMC8Kedb
6ACl1cyC9ALko1xenMgftYCqWFRCbq691eg+j0m0JpcG6VW+o+VIj9EHnNS/Skhc
GbHbqk9Q7/u/Z5ePbUDyjHiu5KoL7TAemyJrKjGrCQveBaH302K94OQnsSLvLVXc
hK7zAWt/hDT8xjTUDlqNHsXpNlxLYmp8YkEeLvcGLUmZpJUqs1/XkR1efSRv2XCx
43Dm32+0zlmMHILEJ5huIJ0AUfMUEB8nRAj9c3MRRS+KxI3L3THxzEK1TD/+38lG
J0XBvahAy8Z0ddpnvxKjxMs3YsupHtIRyOoA1QCTgfhyhqGQrm68TcWCupeaTlNP
peo9Dz4NRPDo07IR49wF79JGzPDjkGqQr/cEAqAHdFkTmGtWbo1GLQwhL6WoAUrv
W8xQolvTn8HW0aX1ZSnVsbHo17TH72Sm7K0c7vFfA4v2jjt3gH+TJs0YmojiOT5k
8oyezsm7V5d5MyhOLFmqIw+2cUFLHoFm4bIYHX7+DdfbarVj8FFd/SEKYT1jT3rS
+BKF80Qb3DYHuAS+tk1lP7Be/0Hx+XjzPFzURf2svLjY7f0Ln6KtHGoAhTesmjp4
foN5L4Dre8wgxfuB7mAlrBGNIV4KFGzaOW51sXH/o6TKpRgw3ZmG9EJ3vEbzLX4E
/9yhpwwyw0sYQUD3eJAm+REOEkvZ8CRNjS6ULgV/0Y0RAnmRWHh3r3ehe1tar4Eo
7uyHl8iEf3MkMzoDOccrFFb8HHk5mHxt+DivkSMRtqDQ1a9wCNO1ETfgza9WUYxF
5HIkn+nfEALcDKyA6qsaUTNcqV1hXN84LwVqECl4WpprzVv5OO/V8Mvn5772fgWK
MVC53iXV5wP7mEJuX7sAkKBk+MTkJb5D3YXzwYySl92E3wvvOVolXbPOKA+6J+AJ
5tp4Pc1oio+iBB0/6POLQs3Y/SUGCkXSmURR0XDMS6J9WLjhutSwTbXAViEMXE85
gifKHZhe7QnxYtrvRLz1xK2HbfGhSX8mWiwOn6riOZiEFjcDRBPBybIpVYekx7bC
d5sSu4FZk9RYA/yYdMnXHw4nxdKjo/p2fY1FK9empzVLsMwKc39/8yW/OyN2JfhC
J13KHIZ2sRYssDFGnIN5tZAEpEfngtNtgA1fz7KB9zTy2fTeA6Fb5WzmdjA20alp
uUNsIuRPYlLf4jP0pmSO3wez49gcJCLQaPJv0lDqJrXeAcfY1SzGdStfM1+2R/dV
nBjUwH1Fwms6XzGaMBBUXWBITGLSzLnd0d59kRyhyw2TIvGTq4ZZH8WqOfJ4P7op
fRMbA4g3RV1XZmaqeEHvYEOaeHK+p3xUffupu/mR0scMwoQJpoIkMFfKGLFddVZS
Q+AH1dziJN+oJUe3ZhccI5Lg7URFv8fCMC/x6jYcvMqDlcUD//A2ZPtuPkDNecjH
wppRNkcNeG75fzbwPgGKCuQ4PjJFAqLHcFmwf9WEqS2lnEBAdwlRXHEHqaChudUT
CE8cCVmkbgYN5mGcCMFiqqbO7JS7tTyKaFUEOxEDLfrVknebpLmPxlNPxJqFXFYY
qbjknfubD7ivJLs6vlH1FsLFmzROffnfIYVxaEdjvpa27fITOIH7kRIS7hUw0WVQ
ImMrArUVjFVQUcgJ/AAuibB2LtB35fk8nLJMexMClx/KGqVTheyv/JL8xFlZlBmM
tiIWcf1qnPiBRrN4KJzrOZ4Oc/vjhmFo9HR12/z8mYV+wLtqZXZ6HhRf2sFck66N
cMP4JC6Dn4Su2YU8us12Rr1tRtnGwv0GskdE07SUqnQfRnsXhyLwMhac9jmxrBqY
0PawFZk3+RHSosiRE9kK4PWt7DlDbMLCh3XWd4iV99sE+nDyuYXXHNRl6O4GHyGk
/bLNLFk23YhrFKEfU8+TpeMRXjKNkaioBULQtAOshq4Z13i5CFhxqiGaLqid6gU5
NOn0ukf+haZw3n6Y7UEXly5V5fHha+JGe1neFJqbGJ1IdIU+sTASwfn30lOIjyLr
fGKasnPF//6frSuG/LyF4tK1NacF7ON2FMDNcoMICedmk/0D5a14ZfOeH3MWPDOK
Tx/BYQSajXV/RV92frK8ba1XYuC16tUwLNaKvl6mWMVrs89AKyIq/3bTL48Oupev
mmz7ezTvaCJmGsn7mh2+e5MR76pDit9PNuhUi86xmWYStx37mpW0/kA1TQVpFLSm
Ok/sypWEM9+XM+BC3KghCd7oCQ4sQzgI2li8Mqy5WVS0+ayMxClmlEu4SGH68qdt
OY3NhgHF0nqMKEqthBTc3dy89dRYNDleXEmPtn8yGHbGi1Yu0d2L6sClaofTcnly
ech9mL6zy1hMeRBfkVyJec7MDxQU2FeKYYml8NYi8GY8wePO67p23n2LrjZbDLSZ
4w5nkDPMZNMPLvL7t1s4v1iNhmkNAPDrD+CjXP+ygHnAc+RuqLspPUGuZO7Zt6Dt
Xz2izWXqMV6u8nwcyS8NpjZBjJlwI1ZjBIgy1kd2ohwZHEv5RzUvy2sAcgQqjk7x
oRBe8X8FghFsYUofSaVodrthFIJ+LjhZG/Bx72RzhmZrwcSUa7WqIGJkCXv5v5ZM
mPFGqTXlq86ZgU0YrxPY+qfYaLD+4sphx8qIYy9L6bzC8JVk8OTmlGIyFoXcT1Rs
I5Xzt21yI/y/pAF58HmhDT/NJA/cW+q9YMlh9iXU5AMlWAI7FITqu1Nvhyzd7U+2
BU6XIBLHzJrPdQGIHdm8nN/NU30g/mOp80Dy4HKytKsRuBF2sXDPEBFQjWhOj1iW
SHEzsF6GwZpXTQ4WaTgL8nFvE9WWnrnXhPuR8TnHEHP3llfUSw/F7QUfA27lrNfX
L2NgBxJx2hmssxAf3SPFVZ2fEkeYD6HnKtpG8+wmEhMIIDB6LSmtBYQGj65w+IVr
gp2ps15fqqmV9QVn0FxHAUiT2uM1CbkKeIqGEkN0XdOdq7sxw6s952VTmq2aXerK
G4Aj5HjfuRXCzG+WpiYxlTjdD5orGNpNqCYSaa0gizIUfhPkDvBhkd+Oy38KStxc
sP3I4lPN8Agdhop4cw1fpHTkWVAWgKhIQFoaeQfGvriv2fwhj+vJY42a1Emf6hJX
o1WG05gDhotq+sR5hJc84IjcVp7M6u1fCOIEsEyWW/X760UL/TnvKmeMkqy3bosK
lCjUgxSIdlrSH+gwWbXgg6aMQgHZjCv22TXmv2UTtH2epKM35Bj0kF7tOSTN9ieQ
zKDtP6QqCvTQREIxQrJJFrCh8hw5ubzB0cGOUDFac1tVfst3HEvr+NxXZkTuuwyu
qGv9y04yleSaYxPDU1ooDJwH/H8DEXoYmMJFUnq0MF7JzK//3eSWbnpmUO1SpWK/
1SHnMclRj7P1cOxR5H7KryFeznh25xj/N5bIeb41+JOJ9/lT1HeMJ25ZG3YUYK+u
/uImbCbO5WMf+jel5HC5nqyrG0dJoBS8djmvMt1JJD8rcWYqy0xPxK6lxaqzQb3p
dZtCfiT/19KDNfu/ijVqqSMxlleveOYaeeILdh5E3LDFJMgL9n4KgL6F+W5rFetq
hfn0zQneUfe1AuMCRnxtuU2H36NorklkFk43F8yOQkomXK5ixv0mSi6YTkPsoNRW
PFdmU87WBnubNGKy2krJ7lbHHKQ6PyCs/gkuIK6HxIa4wL0XBQKBcjbVVP0RvGh+
U4zBC9XqKMKwyYldAjN2MFyhKqfFRNfpetPCT0DgRUfeO4ZHDbJzXPV4G8+OKy8O
wlwKVqQt+KOZgvk4rgJAPHRcIw2+EHZsF/ssT/BydT+WO55NL7xLGxQt9JLAFpor
6AXN2VSx2qRlKVZKSHgY5zfpE9fgTmDF9kIOVyGg9GkrNAqFjZP0D2N7oKXnNezS
il/bgDfeGxyEaNaLY7cPlmMeshiSYrnrAENfZA/wK9Cq4G8HEB+H+/SHhHfIVNKt
7PdKU4ZNMsPTmBZXgTZfRizMm/rbIGAXJfIh7LDaYjEgKjH2amV7b4/QCAEbJUPF
nn/CY5wxSBNdMEkYgbgKZuOGO+QR2FDn1TWxfPJ6YnF1lReoewmjlIrjq323cts6
CyXydGUDkqxMjJZQAF6o5ohTK996PxJc6m6HUgikCrrGvZ+sRwH/AiJYK7EyjJmD
NaG606+9lV9x9HhBCTOh/sTRv+rA2gGzhaRw/20bmy9tBnH++EBfSIDkfp2HFJPw
+9CXYtwrycXnt5OZblFO77Vb3I6FP3an9/2rUI9GofhiQPdSEP0jIt7bLJAnE/a+
9ja0v0YZSdraCmU3rlD1QDKIXk80zr2/v+0x2lLyS79cr3gJUmJHHBUHq+TJdrAA
76J0TATpJ1JjcUoawi/0vx02Im3ArIeZ+61M//47QabKVZpSS9tGGX4pOFRC+syy
ZvVjQQSpF9fb12zVuTzRXV3vqdn8NVseoxsLj4GMzlShIcbDRNAZgSUwYryoFKBJ
Q6TLTgXvgXBGDuCv9CaKodpONKaSQZ0P1J0U7zAovjT8bDq0uqwmTlEJpkmJtFgE
aiHRTHga5D1K5LUfo5R4iUHANVMYeXbZZNq6Ar6Di4zyQXzErbqVW3UiKl4BaRnp
41K/8ebXV9bITY8Jy9j0LgSNDFjmtoRXNNGMIErJm7dqrtTmjp02BHM3ts38zM/E
KsCL07OFf8NfIznAAB6EZH8aCEjAnvfby5Ic/sMVJAXjy3UX1a38z/jB3GX2oApu
33u67vyTgj5KFRo4POV0kGN2ilswzbkteG0eEoZcO3yoOSPR8sG1wp1ZYys/R1OG
cbsT6esjZL3QiTabSy5+D7Va/WMz2O4l0ISKgrioerNYUqiN1sVU+63woS9zvVFG
MByUWMq/q4VTHjCRMsn4mzIHLQ1jynTOwBqEA6/R7vck/UTj1KCCc4PvZgMEI1np
o40CWguv0TcgKk6uprGpVMAsB0/6iT1+SfYnz7QewRnnR4GdBSOCBfOMATTErnaA
491Jt2Xhs/j1Nd2aNfvOYGT2OzqHKSOAb7m+UPFxEuuXUF2OunohHyI2xNMvdCi8
gs4tSSuGi38sc5v7J0jww8qkI4Brs8cUMXNHv/VTTMxIBLUs+qfGr5lgcnfjd/+K
YIQVCbMUkVKnWAwR2Nb/7/thEDpM982ARUlzIWiKF1ufLkuv/RfVHyDGaTwvf1zz
j10ZBBDdtUZPcbC6/DzzZMvrPHTXK0YFAySmFQVF3cLATeRJuCpGMMmP70z8+Hbs
pe8RCLCmV4xR1cepZp3+HSehLVpljNi5X4fBtFlVPzKlZIiOu9KYGqSilbWKPFiP
z4tMCf9ENz4hwG+seQWdjkdsfA1cBLyNIm3t+o9PWeOkp1yJsCBQ/k6QDLm9yHgr
WDcRQCrRHBEHCLxeZiAgP6OukSdvM08jfw7zvXTBKdj6vf5h4/5VrvCIzWz0Z7+R
K6XNxdKUOIt3FNp/cweyNvaXJcEtpG5wRV687mqL7vkj6ds7e4vqWei4twtEJUkC
/V2E2qF0UB86uFU7X9MWOe7JTVJU4V8bF3zusmwQFGA5K91+ZCcRr/3CJHGA3G2w
rrM0iBGlJpZyGB7EjV2E2KRMVK/jd6Sb6h+rL/C6Is6sJKHjrVekB8I6fq61d0uL
SVRIkPPY8jWE/Yie1sUpm6T7pc5JBWPh5fWKMKa3qcV7dbsBgErvDgLx7epS3dNc
ofoEB41sD7n/lK0ZM0gDa4EM4eEAsmP4R4xKfLV/nXCTC8f5Iyi6TvmGOY37Ijnf
jrlu0GKm08x8AKK6UEnJDS9rRSfcuuPw9avkxze7ei5P9JPKjkKNtet/TGEV/XFB
cXyA8fechvyFd2QyYhYIC4ElvciqEsCDhNWNV1N5x6M/gGHay3XygrK/I3etUTh9
2fMUhaqDdIx5OHrNBD5Ke8Rg/sPO/qyukWA8gd02b3n9v+3ZAAMdCXPoShHxAped
R8/NRAdtV1wn1UBGlnQ9OzBZsjhVBLKGollRRoY0FjTa81MF+ISlxUDUw2/peI5E
oQqhMB+bncHEybwX+SfWVazaVr2/HtlfaOp7zHX6pD+beTj+qr3VU9Tcrlfb4+S0
ekwwlslqSIdlN3LxvVqiZngSOKeUsz/z9EvX90gbKiKaVARnyueHGE/ky94hK9Zt
3owzbBSl4yzGdV1EWzujPwaVif34+SRMBEm22FvjXqxWHtcgnEFwQhJoKikElMkq
e0kNRaTUe9ci+2hBxFJmqJaIP57F76Lcvvl6FKK/qjoOlLXF3eApK0XkCdvuD4mx
1ZhQCr3/v9jL1vGA70Z+aX0OCp7L1Gqmv49/Cr575nyQqRw04TU1uAKDRgl0lNAs
x+F/pe3F21UIXh0hwLmaQqXH1OrIUEab1qDXwqaz4aKSY8GYPo8HsQtGgssNr5ol
Owv50MzZaT9X9oBNp4ASfSTkSyoEzZSSqsldI3txPGq5A8DeX/XdNrUWggnFuWes
E0iuEjuhynkSEFU0LaL2Sky8N2kuT5jT28sqdAzUcXVmjcZ/In1C7X+Gph0dCiR2
9zauKHVEHmfmLeixKTR4k5VP3F40y1/S88ZmvVl9vDdx6RqAFBJpnHfpvV18iVYP
0ElrOwPsQwGAa9kDIz9JABW0ym2y4aEoYi5AC2AeUb3gz+v4WEI4Q7fPHKVvk2Hd
hfcYCWVTxuAaK+1oMt8OKmNC+OSOakBTDMlZ/Qj/vZ/cD9z8VScA5CUy+3bHU6Xn
Yd+ze4z2OCpRxIovH5awm8vcVJ9v7F5vLH8V1mhtqJ+tqfH9t2gxjFcYboEuDyYm
JKx82kirsCE442hYj1QUqShj3kZK5Efzd3pg0xhgf5HnrwTIn2fo2DmpUR4Y+j8C
7uaPFY2jJU1KC+nGurL5MO/RBWwHd9Zry/Am269mLctWuGT8kbp7sF2f0VqP6UG+
CHPRhkm8/lTVVqzf/iyL3YDMI+cQTkB+1gYydcqRR+03G7z3ZHywVy8O6Js4fFPH
zZ9mOBjgcVDQs51/5M8B7X6MqcaE+aIFAKc/j/fKkmp4/WQ4srIOvXDzHdKhl2lY
Vx8yL7k2B20l7RIaEbrbKZNNkkcx3svwUT4/+YP+fEkBHuREgcrN/W2OQGdpAU/e
Lke24IKxl4K88SYU3fY8dEPo/krJ0PzWXRK08hGoN3FX89F5Ep1AgJ5KNW/88Fg5
PX2F4lM8iLHaGFpLxZkG8sNs9kD8xrZEjDNSgbbb7PMzSk9Gw/bT9qISHPpTB8TE
MWyfpw7lsHTuua61qDcy9UPFQmwQHIj9IScxusCBUkn8a6STmn1CyTa5OslP0cjo
hZCHpJF/Cgck1smW4x0pAskAREUmKhBpSQNCLzV+rbD6hiHt0Vrl2Wo5aNUIoG9p
+CYKrqa3BXE4j+zTvSSLdORr4eBI1GLHo0B4lNwxJHixOrPUyfFHB3QLY2N3t+YL
DZqOec9FaEmhhVr1JmM3hv4Vy+wrcF6p55+JEtmdbb7mmhLNS72+SBb7ggjCV/SF
IO/5E4TPXsZ3FyrlahO9hiGfWYeYIxsxKzxNNB73mWLUqbLhyyM1Ok+5Jz6fIIGg
SuPEZ+Puhy3mhnGpc9cqXwens0Z95cWZizWqPEa2hPQNcLq4roRlfkPkIP/KV4Z8
Y5ylWDZ8SwRTI7C6c7gvy6tQXEEkgTXz0MOegBtpnSKV/Na+8B9nuRSL3CUQ2fI3
LLcqWfaYzwOiC4hJzi4dSCPJq84zlLY17FWfwpp+wC/b+D5dIufxKKpNDj/3Ym60
IiQCJSX2oVAyYnMV9I919tMdMgjLE3o2K/Xs9HIDnWosIwEBcpQh0YflOlnX56Xg
/bnb/bfGGxJaWkZkL199GjgTDAaBQuV/uy9jq5BEpisrlojZCwvtH1T+674t4JFP
CE3/X4VDp3UZ9SYN1LPvynansCnmP+0kyKeZu481r6CaSPF71UmRKQkwwzxabRV9
B4U6Esx9HPU7LmY6npXIXz/aQu/dPL/nrqaY35tjyNY+VcbqGBJxtouGS+df6E6U
zt2RpPX8vdQo0MXwbrx34ZG7+kQG6BElL7IusYnHa/CdW0UM/L2G+77VE1p5i2ai
wflqOkuLtcoiC+VKVN+/kKZoD2Zya4Pn+4cQVdjIBJDsT7BC6FK3RK6RUs3hXy8m
JAV0IlDVVItJli+2djp38SGwNNIiijffUsp4D2kDOX0PfWJ1caiFGokeZybvcnjt
OMct69roHq6pKyaZ5oyD5dE8nU3NMmz7CLn3hAhUT+NlEKE/mUbjTFaKNmp9bK3A
pEM6XEaGexbhuL14n4Wjtv38FFXwkQ3tkdhmdGwCWfZAkaF6xy26Du7NOLMYIu9v
ipfKVPa2+9Nre8yjt4reN475VZ70ld2+yHTFq72UZz8zAt2LEf+CST13Q/YOjOaM
HakrcEWvOYN/uDg+4tN3AU7O4bubxmwX4C2hN6COqiN1cq+AfBvIROx9YyLy0O1G
pfEEHrsrJVooo78rLFsVuK2Rj3bMyHpxBpZr8oN3p42HZ8B4Imyt8o0xlsjLzbGx
jNdVfdhrQxh9L0eYlObglN/TR7YvLaX1G9v2zXBpaWfg+lLSAiO8D0Uay3CRJG3+
5Yz2g/qBzm1O3ZYg/rnvxkVnxGYIXztoxuE8/3Yul7zcQNLpicNj0icqgTgxcK5x
VDE1HnyZo3+WGZ8BmqbIe4/v99RiytYrWiNUQXBb9UC5T0iNH2k8okyXxoWSUCqW
VEk1gPBbt77AXP++8dfAH4We3jSvC2SqiQ6zSVnhv578WAcitdpi81pybUsYnk1x
D4QNdPCXZp8ZjoKKGj90uhkhdVUZtUFC4bpZJeBDrmRTjOmH6NXqXwYb77fPUFqg
QPW3Izpva7o9cSZqXTczV15AKXQOqVXPlV6hX56dqwlZmIs58NV5uJg5PhDEKsLy
E6Xw/ReV0YNgKi7cSdKA7MP/adgKZ1YcixOKkRHHTcXh3xTcsCrUipn/KGsP51uU
j5BQgU6EXWxX/x7R+k26bW4t6GLbYykz1thWrJNRUgDwqkDl3iPmijMgoLjeP4O2
kBd/R/a+wIkZXp2/eaO59cKHSkoYzJraDAx+1ZOUnnBTlcS3Kn9Y7hWC04h/sO8U
dAoyqown3xeh+dfAxZlzks7mXfiFJJEukV9PhWbo/WgMdxD4mPub/fAxtiBaURGA
1u5ipEmn3DoMQQ7JmA1OQZqfLvahxkGJKok3P2ocBRqKVJjcX4YDy1aNLB1lgHgE
pZtKIjT4DNaLMVQ8xEpb741bOLb+tapy9KSmrr5QQyt+1YK9ZqFMjS2ZGGmNwn+4
PbPGCyo07hDFPPKW+s+KRdlczuHdSCK2Y+WsmfersYXkmA3OH8Gkdi5JaV/8Sc6g
kakxgGmaLtGJQZ8BwNq8deyeOpJuw7SzjCvF+s8suQ9XVs7nYajuNyl4R0RHAUPV
1/lM3WoNq4BGGOJLAbkmbbmkNkfcEqFWQTYhABtuJ9i9FQTSjQwMJnAOisCigpUg
RXZphkupSZTiHcAJxlpMWge995CsIty16P98Z+T6QPA72keOgH2hxO+A3X4EmDeZ
amYBErMKUKPuVjs3ohwlMZlsMNS1gAUJuonHZ+RrlWhtI+mLfijqqt/Q+pq3yEer
rh4xKrSY6WQKeijkFraCHhNiMwFNoqEQFzpMpagz+d+SaQa+sjE83Mp8moF9SdjX
QmuUM+GMrZ109cFhlRDxQFNQvNnU3XMB2eyg0i1lIXM/sz4+fl8T9VhptWQlERv2
ggRrxGF3dqqjLh8FWZEe8aaDsDbXFpc91tYHUlz/AmsZTKmjIpwXAu4Lkco4COlL
X6be309UvGl0ht2xEG6bwqWm7H2/X432sbeRbGODWxWQ3/TO5NoCGg1rPYo0vNdm
U1qfY8xJC60wtmfYdJWAT7i+x6UY6KTUuNJqEMa1WHyX34W1GZn4uctKAIifJkkz
yffcPCz+sBprpfAYrafh3ytVjWQMBGG4J9Qrh75RszI/UeH3O6DbXnq6/WgWflye
d9QrIbp8EUR1QOLxXowkAuMtxED/93qdHj2r6RlEPLspXMIM6HC0e5DJRbK+53nH
AadQxPRFLmNkChvjNNU63p/aMKqZ3ltDY80g2pp1bgl/78gPgC7gYE5Ly3+opKva
qDhw5d+HQDGvF8GEuTBFpDbtzIYMb5w41pFqcUrS3SgNDjTN6rUdmXbVHOQBjAqa
rgf2y8B63Udv34rJ2CqIocV0nkj/MuiSga3SseeCt6H/Uy9idQpc6uzWWlb4LGGx
UU88/a3yeAeQyxIE+WOXqTwisSqrp4H8MwB1jvdEErEGQYYop95+D2Yg1T3MCul1
vZHaPK98APBhZ5xl30GZFPXHdu2cF5u0pm1O9SvSkxi/4Mv5c98TYTmByR66wpVX
N9M42AgayyFkFwwoI91mFcqzjD6QV/iFmwJCRe4AluFMI4mYUvmkSYTT/Bk6CHXJ
prGY40e7L/zkeFI5O6UhTIaTdrfkD9zojllLAQEBCtleRIp0Fh6Wr9KOrVSQSm7k
gheRoFrOCQ6Kgf0UgyxzEfn/+5DAC5E+b7NE5xEHQcda/vWKfTfXrjf0feLc+/S3
ZlkbSmxGin76I5fQ2D1eTnHy09lANHoRvERsyUXBkKcNH82zZwHZg5yjFh3/Yyb6
lGYMWunkCIfqhKJRfdGr1Lb3WHK/xDx2iKcFxoL4lzbwTTVc/RzuWiFzDSAlL6N0
1+JAWwuBJnxm7G/jaAXxWy682sjsyrG+FX17tfvgLl3XY5V4TAWCbVV0ofoWAnbb
TSKZAFjDsMZbzBdMeik4SLXtvgyLSH11qDhyTuswzymeUUnAr+f4mVr/fAmhpwbR
KQPGyDOxseLWWBBqVCDzfE95slW71TUAPIO1P39GaxiSUWD+PGIVf47DiLqXKvXv
/4BDTAqwFtYN+oomuSuGkg56NpcvnL7moBrWobKLWD1IGirwBgWJSZTP94qTF5X7
E0sCIID5YU7E3/wCQ3VxwieK/hcCGHTy4+WrsTrr4Y8CjdG5YMF9SXdifRXopTJW
TMW+2ew3akb7lGh0BwQeNDW38MDjUqPyAD2201lF9w7BGG+H5KX44N5rO/+ttVrE
Z0Uhc/E1QX5rx3jZZN6zMe7c5DhIQX3ynWa33JE2Sd6heRGO7VteEBim53TSJ+8p
kXbr5x1C98A2y5137wzQWHLochkM303AWx92uNvjdPNtL8BYt/v/x0nUaVZUBAo6
+Yrb8BPAh7Pzw1IJPDpJy9wm0rcRCDi0U1tSn6rN0dK099cbUWgAFLFEGhojJzfZ
KQhlJ/GGha0ZEytmBou74RYx/lzZI+cW5Yu1Qr6EjXVyNJfIwaHtFXh0XQ7oJwLQ
p169LJAFM7Yz6WCD+Lmfqk0Py+qloA3Ssrxkf3oxjJC6plYTa8tqCFTRVqM10xMc
B4TM1J1bNSP1sd1SmE2yxgLB+6mPBSsSBJs4vVdo+/o8oFNtEb1dIKGiY1DoqpJb
lmBL+jr9vOfXCKxCdk36vsSkrR8Z0cxewF3INvAtNf8SRYKHQyNfIg/Svh8+2Gf/
cUChNZfbvDwpujKBaVdsxhO496MfUD4RWxRteHQg03q5NFSzOX73VYYe72FDK1ey
MNoLOFJdS6ISz3Qv3CVAOtB2bk2kNj+v7WGxm4vYyB0UmVs60tdnmKlaBUzWICsX
PLxvuZhczyCtCfdKRXVyrUlPXpKbIewKTDPtoaglAg28xJcjSCMpfv/wLKhmshql
DoRRd3bWBpxw2z8TzYKH5I0sC534IKwdpx3LBk8o4SBf0AP7ZHHw2pcxSSHy13Xm
2qialva9/LoOtum3BgI5V3aZOEFFHt0ud8Be/z8PR7w+n7r4wbww+XpUgEYR2qvv
lUiMNlfASpGW4aiQM1wvxXwi2lOvmPEeLAO5ncbGoihToFs9dsT4Q7e++ypYL9QD
5CfvO3n/FsBGrrfxXtEqGIqsXm19jYH55kkOFhmxtKZLVlCKyqGWVCdNJRRtc9jU
TP3wRzr8RiIbHf49BJpbEXoKNyOmPQeODK4worXRo4DU3jbzJMlZv1oKSM4Mw8ar
zqLwVuyExq455/C+q+5itSK8ryECti/Sef3pjYODK/fNtyWMjOJyMxReErj/sHKb
bDaL6lpn5lcI4grP5tSyxMK8nTS1TtHCypYVHx5QxbSZ0AY0IKg/kaj/DfGtcrdP
ojLivbVRNragIfSaWEoWS9AJUiG/ox47m/trvFleC44X+X8FYeWBwAmGShYxmNyf
h0UqImtxyQwIXZTIP6IhkLCBY8rMEYL4dzuzU7jygbs/PT9YQK6QHgVbZ3IH+3Zx
R9ZOFmDp7s7eIfOi64Es2QrLLefrqjUNBMDHnk0ivls8MvDEZAE9pyNitkt4apga
K/oy2XgyWwP5N2OSO32qOMF6kcHKFEODplnz5XjeY/mKYJs/XLdU6UhOrwqYJwzH
1wu9i7hmwujI5f7qaI2Zcu7REH/xGUgd0oQ67ksT2jm/GyuAJybXMyPHEC0B4AG9
OuhNyTsRudORUBI7P4fkeNCwltoDfJTLgS1PJXynT+QLWnkebqHUQdR9Ra+hrJng
KuZ5YRKwXclV5KGajy4zek/9ywKC6eV3yZgd7SdxhXmMrp7fdHMqKWQvm68Tfu34
d4rjLV+eqoUymHL8qhS+qAL00UVSQcIGyC5HG2EWDAfptdevaLSzrF026IzHMeru
LJXEEPtB7dPhz6Gtz/Nv5I8u9HHB/SWtkEEWr5j1VX+iBBt5VAI3LP22ObVg48Sb
jczJ0a6Ga7m1ZrCV3GWAIZBshAPNF/uswaxeoobQ7XQzG41ds1YZiYbf+7z2g7qR
jbwjN8yy+m9PoIbBEGU06xLCidS7RBL0I65CDEAzS02rP45xNbqqQ/766B/5fA1S
gUqyojyds6ptGQEQ+O0utD0kokAw6dufrmL3J0EITyHfVmapPQQQEwvldPw9HeN3
qY2gGsDLJy+iu4P9AN6Z3pzc5DizNeFSbU7M74iCMOI3WVXeCeVC5CR4Z0J6NNRI
A/cNEwS8QFdyVswrwHV+P00BQJZ9rGULRg3P4a8A2meNmSPcutm96ezBBeFPAAnk
H3+oNL8p9WlhjwcSBj7ruTh5Q2CSxPGbf2IVluGUm1zJR53BmjDFGII6h2Z3oszL
fO6R5laEv09sEAyBUj9Q7gP4WBc/NLS1nfRI9PISlPKJ5VKQXOHV2I80fWYDWICH
IfGoMje0xZcLa/Vu8MP9qLPEkS96+NjytGp36dVXqMjIMgkOki9Z9gwVqN6L8DiI
uoVqaXEuG/0d477RKU/bRM2R4epGph/tk4N7jrxEdRM36Wt5HcsYL7xt8yGJD0WL
jb1p5gPfl6EIlRfhSEcpZicpKWxfNXV9Noo/ux4sN6PPYosuEjuxToNZa7brbR3Q
+xG+l1ymUK8+WMa4Be1I6PWLMWujkugvmPiLvh7VcJ2LkKZF0GJlLs4gHn/z1B6i
Zt8eXjW4KpHFhRcmbRm0h8hiCmIOtpaa3BodUBbIXK6BarFVloUM89X8MFqWBsiy
HW+ZoEenzoqojYnIw/LerejPTvW0U0XTgKm88roYar0rHaESMot2r8Nm1lGpiMuM
YeYo+AUCrDBWc7ew6qJoO2MBYZPt0fWAzZlsjZEq1fLRjf3QMfsOgTHfIS3/X9a/
yiS5T+/I/e/nNcdau9Yty97Wrn2ZB5iLdVuUiZfP95njLl/aDkaxdtXiSTDd5aX/
61FX66q353XBYON4byGYuXj8NxQjuwNq8KEfj41V0XvWEBqvY87jpmhPSo+jhOoN
cNx6H8b/J6qDRcmDe6Qi5NLtfVhuAt/KVYHYFxs/d1o2+zyMIfZa7uCxY60N9XRD
fAp78hUut5UvxnxgrBA7Ubb11iOAzXsDUwK2L0anBvQF5tkaOTLUl/+q/Y+TiFQl
n8KrOwH5dflDuZSOK6U9K87oP+OKooGKuodS8t3y8fHO22H0sVlbKaHgcMRvjbIs
coHd8l/TATApRJkF+GUxEowA4/hg1WbM7de7w6rB6K6GeOw+fjX+ASToeenOVyUH
3E3w56f/MRAg97Vlw9hCS2sEl1J//82+0xmaZbWQCAbJb4N2gb8sfBveKdJ5OJYr
l5pbW6+EpTev/qz4ZMN5/OhAjLb3etgV3meqCtgF0aCKdaMGIaYdiN2HIpkTZ3aY
fSH0MvwdXvV7i06lf9azzKFgGLBlxilWJIb0Cx0y46w5VX5Qp/3XZuPNxbKbU6UT
n3zXbMrSWu+bBs1q48FLrQWcEbSoVkY1l3nYmTzWjDO3CnzT/aloN6hfNvkZqSMm
majOfpRL9n3cKusYUt5/tRqAF5MREued0Z1tLhOprUP+knS5VPQe1Yi3QbeTGxDT
Vsc/T37TY8uYuminM1V2LNuz9yKQ6/zkT3oCmdwZpy9VSW+2koJVdNJ7Va9XgIzZ
smkYX+Ei6TSmnSuD0PMEs53Ddt1mJyxyT+uOelE4ps81PxVkPpsSXKiwgGMo3EQL
w0s609WM2McKO13pY6IkLqdjHMSXMKDJArqH3Y6OY4dT3Q/Fz7gxAEnk0n1UU6F9
2CT5b0k8U21AceB628rgZJkwZY7fuT/+ssnqU3ZtkWBFvORPZvMChUsikJTebs0f
Svpr4XYVMQhzFTBy/oWbAk3GXPuISUZnDLgG/Rzgu1HrEICNn3ppTuxxHNeb9g9n
QAh1jXWylWL6tDj7A6sMnflbHlM/0DcNJFyxw5KfSexVS5ibOzSmD9JN852MlQHL
ydj/dtKbB9CLRJqbLWzH1w0We9TOJe8iJ4Izj3Mp5d94wK2Jg7UhpA4kPBmcpcpZ
7dp+Da1JEdTnYz+jM5IMTArhuw3LLuG4NPkvLceUMvOAYVQh0oTd9qZ8qnhy/WV6
orSs9/cXl+H+J2iELOcgrZSkMxB4UCQ1zWYLcDeLhDeFZL0/woYpwBAykEkWO37J
QZi5N47aHuCjffBc4dQYc64MA40ANMC74ZdJP60/JG/hpRP1bZljNHXQn6t6u7F8
ciAoGwZUnnjDDBN19LHQFidDOhRXZ/zWb1JtAeRisqRCa8iX0qeq8xizideGLHnO
QfGp/XyLCc2EpW2iGkYbiDed7vyFSC5mgwx6OsNpxP1lGmg6F6FCTkNK+OPJF4KS
06LWEGdhW+8RBvG8AYmqY6TGIspeE67TMS1yb2CG/A3OdynwVeeWwyK2tSfUOd/x
MJ2i9i2HxFkkNbkyfMePVuETuFkqWVmQFeQkQniknEISPkNu3NdEk9rge6D9i6pL
3X9AtIE/skKncJxJX/zeZMLgq58tlzZ7BRfEIb5VJ02bOP4vo9fbHrxesIPxxBmR
06HiqxPF2gb29VHraGqjWnbEWzJHS+3GODJeoXBgVlp9YBvwLXhd4MhtQ/DsiYvs
EhFTwRuz6HsohgRt4vZHOz/rVxHXBPhmPor4pQ9WJLbJqETvbtY1a/op8QmB9L+1
VddjYhEfLQvIoP1tgRHcirx/0pjaJQK3KqlASuMjanD+/LCljgGchc6agHnInvRf
Mu1D2HtIkBdenVxhJy2az5zm1YWekFASHs3Biq2hU4MFbrJlzsLoWWo2feDjeRjq
sdVGopuI1tPmGWk22/jr+vbYUcXWcSr1hpzSs5KBUHKpGaPqw5FyeYh51ix7DNqL
YBSR03bmMZ8KekBiwXN8J48cvFLjtnG0wIpYOD67OEOlJMhhY/AJYTm7+Jvw+RsH
LsO21s/5HLmnvskMKa5bBldTAlpHUXml/4+JT1/vhWgdfbey1yaKL+ePzE/SkV1h
7bqLd+EanjzXSD0wt4MVvZKF27BeKg89rzptZAa3seVoLVUln2oacQImGjZ61UkZ
0cLj331gj9pp2LhSWedZFMRdKNgH7SrF8sqJgfFO608C0o6uac8MO3hp09jMMhZn
pd3WBv5ydiybL2VrQVqKGCpHlsY9oDXZvn9DZfuLT0b5fTyZInZLdlaPMq8kZoPp
cgz1w5is8hyHRVPE0swwnv+gznQVGRf9f+yFZyP2y2yEG2bZtP+2WBGD8EjnELNd
HnioFMk13zuVJYteDXQQMnC/n8y70Tgh7kAjFatkDSs8uRt3kFOPJ0qRz5qzui41
l851Ks8BFXv6VRrXrxCqLFsYu4h31+3UI9kAyGz5w2QIk2VODCCnlC1CnYVD96y+
qcBuO2YNCjs6LKIobrWAxLq99h4Z5tzjHA320BiWqXDKL+IRwns/boxQWLhj1iyv
jE2p5eKJl9zz+FhTVz97mkW/VBu6jUP/kX1SVSXK0AgJhJHwhV46K2ux+OXH4/GB
1Unq6IE+nhx7h7Ghk6ypf0Y3ZLi7lvCtEXPPF6Dnjjg3BFb4yL+Obn2fzKZ4ReUf
saRAyjJTokWGu/XmkmZN8QJdllTEMxXJLEPnQ9IAIMZzvgauiy2rd4g5Wn/2YH9A
cNANopRxgY1Lk1l3Z7Ed+qatazjxlMpwFrES9CTZ+2tJ4eikPRBi1hvF24+MQL/j
g83GWfjDD9YO+cimGiDG6YBa48Cad7CKrcUQf+EI7OAMjmFkYB3cVU4RxuxpNhvB
YDKW6YqjTNKjwvcNx7n+BvQM0ISkhe0Q99cY9sxylz5DC93Y1xBGYEn6iVdC2oVF
Ssb0YHsFOoLAl+4aDPloQ3GesNpxxjfk+LUfqc4+6zQ=
`protect END_PROTECTED
