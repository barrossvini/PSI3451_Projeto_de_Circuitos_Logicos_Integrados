`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C6uhBrGHLw0VQ6W+XJ1wAv6mficIDILh0kQdrrA/GNEp6dlJnpYAZNKONU4M/c46
kzq1yWfVplBOS3bEWDjbkMoWyCRb0Z7coIlLvUMsXRj6UZlD/4uiaSw+HtZgoMvb
PyBXtStRyOYh5hnl3KOdtQzFlonWCsRMkGVh405fZTD2v2qE26xrKY8tRcP069id
vpNnOHkYV1niq/ANNjwo++Hq5BrltRrZucOY8O0FptkUtvXplVO4CqIclvkcJ5ed
DQhGbHVHb5Qgo4+VcMGNKlSOCwUFPjojiBYadQsxgK00aVcBMafg9w53jYYh89Q3
bUQGaoeoSS5BLGQ1s9CR7zrSul8kHRDSN+4j00Zj0204DztFcInFmKxdmsYF25a5
lMz/Q6oyqIbmhZ6ttLdqfbC+2k1dBorJP9qkARPMeLdZryXeAw6nXUKAw5KGfI0o
DCgi7i5kh1AQ5X4fUJOug9PURnoO8/ZwfGaFQg+9K2JfVTcauKdKaUR2rUNCAZuw
9YCoqXf3bFBR5IUuessDbiUbYWdu/SJhSRFGqItwjKa2e5XjIO/046l48AajXCdj
QzAvaUnOtO+hbj4sapjga/+7qrUGWIWhZjSSBsG01z2/UaORkXKxv1l7J9F2aUGH
gP/wuVYL7n/APYuLh3GHjEDbaks6KwMbYKqz3kQb+ArAE9cZYQVOq1wOWnPOLpVR
QPf5JQ0Rl7f0O44Xo4S2uquWpmYUeyikAO4hkdXuX8mbfO373R4a9zTSxtIWpvUo
vTg1fzbV+MauIUhpyE7wAjSjMl8Zg4kP8dbgJvANNVUlMo+TY+aT0+qAFb1xWgMn
JZViid4NtFuHVbeI+Mi6/QU91cfD5STXKkzpqAepIbv0S7gtjKvQ3DBaubyPEpF6
q3ieQcsr7H5nPg3hS4DLwGrxjW6Qov5GqTIFAPKEAWaA+5Z1uQX9XDmsSHQtUNVa
iZFXxOFk+4hXD/IJL4NGSwUqVGCJISco8J58lJSToNbgXjRTwqrcwDJqGzAXZ6tQ
BHp3PF4Fi9oCLuoC990hMfZ2ESfxXGPRKsMgDqoi3j/hUbwx8T2rN+Ky+MGEs3S3
ZHq8QIlNkCovdVlGzQfCwaCUhTorja+2/ufNYsp3tX6KX0rwAyRK4+Lc9zwiN5sM
B67oEG7TJCYcnM0vxaF7cqn0XaJR4y+fe1DuB7vpYW5wBf+p5yTwbrWv+D+Rm6To
LNWtNKub6Jz+SctFOv6fgAMnRXZzPPqAgpCwmK9L83YeyHTLCyEAlgWh/bBmC++a
9tatwoTXVFaG+qXDcNcp3TpRTVaYJTjl8ATmd23lU8TNWj6R2Qp2NDIe7tVAZ5Yh
wGHNxs1TL8/ero8MsqS16dMwJ4zSEDlNWdlamuLzsdu4T48EtO8wsJIbyfmd5Mdz
`protect END_PROTECTED
