`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VjZeidChNmJ4HjboylSgLUxsNfQKGeo81HezMk858s1hZLA9UnslkLtfpkj/aCIf
cPVeP4godqrVEftkuiuqmsxOGjZo+h1i1dk0IXeh491XUcJ3RHe1FBgL3xBhV7xQ
P4wZuv8qs5WYpDLPUWXFD5w/tAct7Fo83dGmk+EG4d+WLWqN8XH8k8m127tDuRUM
vhypw6vmbaei2RSIRno7RE+m2FO3fOGsIg5kjfC3KbhQLaffvqiqMqNIa5X4vJHg
HuBVjBX63YJyvXI9tIdc7robgxaJ9NsLi9gYdeBGqBN7ZRbMbWbGKXZwLunjjuF5
q7X2bw7NfrEqJEsFa+Cj3In4mr/HsKsQ/hNIK/D6IUf25kYpoq4qfGKXNYcKHR/u
kM20PGLdPHMVye6MgfMPlrHx5H8Jo2VR7UYQHOuRF3lTqyF+ZenBWagIzS5DVh62
KSJLuKqXSHF3uXMjjmIZ4ceUyx+bdGTGDltPh/BLlR9Lh99xevdTSxhdfUWMfXkj
Kx2Dlq6XU3t5chKBGK1J9wCCk/qCPNQsXUikPoh3VEv0OU+RvIT6vSF7if5WSk1c
RdCnpmo7LH2RkUgkcQ4zS/zoyC7y/RkvpPvpUhT60r7p9lgIVEW0yZAyfKwaNVIW
2txXvyEWPVjNHBYTVt7g5njgAqAEN2jLHK7MxdkQ8hmakQuGM6AsDRKnLHti5yqL
C3npsLXkFB/ruiYKGFrA3NLrrAB6kINNGTCarEE8n/un6IWbNLXVGp7cDtqCMS3+
yxe7d7s0/Wyv4vsP/jGV3TVA2CPRilPkfnVp3rkS41ZYgPePDRiCQVFAqCIwnHUr
caZfkmzz4GJPIfCbZEaW1CxzuC6KwM12nk/cILunz92cHX74vVZEhUi2e0p0WSEg
`protect END_PROTECTED
