`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HbYcZMtRuwvgW/mm4xzpSKDrKMacomYYuGOR4qsm1STWsDL92C9W5cRc8l8kEtsP
aplIpvAn6baIiHQejSX+akBT6l4IzWe26eY7CGynHWjLYWnvcNSicpyRMAziDS0b
DwM8sEHBC+D59sXnWOkLC3wo8gMJ5qYhzqG/Lk2b9OI7bOpJbvMdy2tqWRnvAk46
lrIOSADjJHkgowpVQQH+EcyIotrCfX49HjhuYz7OGAFZz+IlLfGSJgx99TGHzFZz
+TaBwET2NLBOn+s+2nccnnILPo2EVupLAlLo787jRUvVsDOOBAE7zaLqA29roVrL
XObETPiFyL3Cx6mNNEzvyKGxAyMnB7IaAB4iN1ojIZg3sH4UDdxKXrMLsjEn/afX
AON7jH79Uy+6cCBVOZ3zEP4u6MR/NuZaLIr7h6stXSZUUN7WwvedQVG8cd5n7YIV
I6ZuGBReA/NHPTvt277HdcuQq1+0Fhbq4zUdSJRiHk+ADblbqZXWiOYuqkTF2vdI
VSLFKfiB1JKs58n/wsQkPprNUpOEfUwLULDeIPnKSdXWHLkHCdmkVmOh2WG5h1Bb
HFM77Q8jdSmKvJamNtFyppxr4Jv4RDW2O0XEMFfzKh7dWoiyDsYE/yH0itjIwrqL
jLG0njyPFY9IEP86u1V2etB4JgiVPMueT6Il4HL33XjHXMsyJ1eRgfXJiiC97R/G
2iMmV3l8P1gJo4ZzsTe+gmbbpfCm7xFzaqry9/kgv4k3FzUzRlIxrqVF5DsWZY5c
cADsnIfTrgeE0fBup35LYGx/mrIFCMHNkil7FJoXvV+z6AEW/RRTWCZyPma/3of5
KluAXtfBimKaRbEjNIXknQaT2npgjjCbgCd3Gk12c7mIJRF6sOHlRYH6bWpQhe/5
aVc4JffRHQYD+hNfLdvDaDt4fQYSxu5sz3RyM+kmx/5tfWpX/SJ1qF9RGNT1IaHr
`protect END_PROTECTED
