`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzVlqWeHB7Tib8vtRivdrViIhCp12Wdj+2xKN2TOrgMzm9dMzlMPP213fzZiiFY7
V+PhNa/3wREPuRvFisYUPnwqufZk0ZUc3QlmYM/N1T/svWdaZGXua//J7PALdn4f
IPHA4QKOkC8EKz9+uUx9owPNaZ6svmrEwbDGV7h4zvptkuqE9qSm+CL8f1WdF6TX
qfRVbDu629ifbeMN2hAVvOazSHdYCOIQ9jH+pgjsif1KDTl8AhfGY99XhSnhMQNd
cNDZy3CE1PBfIML2QzYVpzqrMTdsKwg8L5RTteZFdNTIGoUSuma9S46CKXTsnBez
xe7IoZd9nKoUIeBRodqcDmRVzlyKqUYtm8Ju6ZIwj1ylHBz7xzCh9wTjLOVmbYe7
4zSu53H+0dn8Ih3tgAeegz4rEE5XUqS/wGyAduJRB1kzRy6v1FP05hx0IVZEnPnc
pgNEehHhXvX+Xt3LmEXQDwYw3w+tSXGsLp55zgmCW8O7vC9P3QcQOSaZdZ9q7lu+
`protect END_PROTECTED
