`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Fxl1Og7xU7lDW8J8ZE9ynPn4F/fOnjbXi2ZewW9IBM5uDTs7uM3KAZmK9GJw6TU
7i2YCRXV9FLo7g9/WJ5/mpaU1QVMoJFUZ+1E+29JEdmvnkFWpv409MWMvWd+DfJP
kQHKAAJwYqVtfgtTNEBcQAPsR7WbjVRhz6W/fTix3Umleo3wRgbg8K0oSix5J8wr
vmAX76nEd/TzYr6OFgrV64+SRdAnx1Rlc4TFaMoCBnDjFPG9KFDofXyaesWvpQmL
BJzNNnFpvbjjnIto+2JDkSw2r6cQitDNfc8Ed0O13b1T7I/FokmmxgE6pNkUkEyT
H9PipwCIacK4Td1gCsLRrCGH8Jl2RVpui+u3HbILo/LtdSX81FYHbRfsJ2UwkN+D
num/Ro6fS7xiA7UiL2WIcpt0zkWrwx43U2GOR5CDnSCFH9pEjFQ0EH4rBgr7O5MN
s8CnQKcyB33qFFYaqziu5cGZTFui7/J2G5ddCZ585MCLuRX+0ErXuGtWdUIOt3j6
7imvu3TpyZf+F7zOmdqLOPf6/A2HZFYRJM0gvG+naUAD8d4eeuXWOatsZ2+7nbaC
NBmJ8t4Quf28m2Apu7zsbNLTbWcXbIT0RR0DdyAJpl1CrkIP2zsj3sfKf2DN8zC3
lVxVd2bi3QvHcuJVYD3i7rSrFVByAsp0HhR9JgDBWp/TR+51WkWKBlxL2Sy+i0j0
VtYsv8yiE9JgNedrnsBYjv6c3MaPOzdVcg2bSRCQL7rnOyAA3o1pKNNqmcysOd/9
KWDMwsU4rUaYVO3sQ+SS3eXqhqPiqsUyTjpOTh3PvksXF9qve9GtLQBDLuU8/ee5
Ot13BaEhom1yEzYyZJD3pJ/ed5VbK7mE7K0dFgTie7rn6ceYWtUAhFXaMd0Od7ml
pxm0t2cBe5OWmpdNhP+7L81hv4YAmdXRFdTDAB6UxLxiKt+hqUOkOHBRHDpGuquO
WE9taWH7ZHOwtpcMiXyqMs+xzlaSpYZOn25TYoYBP2jWyQsC0KfGDFbhV3SXeK/K
ufNulbnvdrzQbg8A4E7RQ1qzZZusuwx84ysTxEpE05EPHzA14HGs5eJIfcXYNHK1
BYkvqfQjpsHF1yOP46zpG9Ur7wMq/J1qyx0p15YL9el/vtwS6bCKHDI43Lrc3PxH
k0BXPPmc379VONAJnvYdGVWJ2GQank8DLBX367VgzbTWfnanIUxi1Phr5klm6s0y
wAt9oiYkuIFpZ5jBRYn3PWn1UT0gmlq8FZ2OZf1bCI8vFnB3YXgmus04aFhWxVtC
xiDOFFTS2P9/fV7u+kOdyvX5NgMbD9LRYOQ660aG5Oicvh7INpqxdjSYXVm7TI3d
u2jkaGZa7tcN5xUpgs3MlLO2yQ7wVBP3DvVccg7lYgvX51bXEjyXRiilfgrmTUKF
9gz47MLnp6JpxEiWJdxYLo35Agew8NHz0qpTwRUZZ/qDYcjrfC9OPWQLfBgkVvT/
X8lQcDPNoYKrBXyXntx3RXgUkhYYn2XEOj2jNvnOPxXeJhL4WvIT72676VTFoF1C
DQgvJeEevXnStgPyS9RanJoZvSYl7PZvBV3XNyON7MzzSVOBHTO+p0x4e2dGp6WG
aQ3ykaPRu7msA7s7ncWA2DRn5DTQ2coX1SRZSXZK/+nCWR3ldRtwlhJfGFgkPJUz
Gu1nGIaQbIS2rh6K2sF1pnenCmTgskYAejPzlyTG29dquJym7H1N2ZR3ta3L12xu
VFEWlSvOL81dIcNPwvsdaEYRp9Xn1SeN46Tm46X5B9EwTtBmzt3egiG+lU4iCaM3
0SH7RQM8TB9C+g5wmi9kHANJrWBKESBfNgEAvaUCKzYzI8L/dnTHoJsoBCZZnbGm
HF2e7UtUo0/4hf79V1XG6zRE+00yP1pWd65IDj8jkKAgFDx+T1j65bgsZX2jnGzB
3c7qLneh4GZV5WOJsiqGCGN42v39MOYXCKRQ1d0YYAXNdpq94vgHRbdnNdsHkgFQ
s/wJ2EBLbW4xFMalQpRpRcAKWdQYZtaWFn+wBxKxcxD8JN30fs+kx/gwx3iC1psH
pdHuIJZrOIvF/nawDlY+MWxRGO28LWpvFN5dOzFF5H11POOCHIV+yQgghLNvo45S
Oc8V1WrUztC7ggIslPlPvOFIkoxsknGOeS9Kn+WP3c+vKdrjZiDofcGoZRKjirAj
g8Xmy45m/DBgXgc3A6TCmliScefR85el4QaGfkSrH0k5re0I7XS8hnjQOdnpCpCC
mnglXPNOoC2UDh6DKlezudkGHkF8wGavEIrhsr9P5LkZ0CL3EyFAqQsUDeQDoK0z
s66DaR/M7/10dT6Z6GS7OrWEUejycDvSFINh3cO96rKCvgbSF/pH06TKlsMy4qrm
egNADh2tehZuGXCfYCAuGVV4tzmekBVcHRV3vfrmV/3STeaG80kUEqTZvvPqTYA9
nlC8Fz9cVq5AArZvG0YBc1109XgKW6Bg13gf0kiG7diDSStAcCu/t+YGXBFhEw2b
dGwu+WGgFfVpQAOHBn7CGDPZ34kNxfGnlCjEEF8ZlHwF9GMWrhoYUlkz/oeLrvJ8
wbwghI3um2qsw1Izj2y/6ru/tb40PV25MmPvsuqQg2JcwORxKxxJ1GbuJZXlBdhV
3IiOQ3OIQYScUdJGy9UyEkYaOoDUH7g7OhM0uYwctxul7aOBjUhZMeKPAfgBVLrD
QOTDjLB1eUlhWn9u5dFqdH0K+uO9Oe0kBH9KbQWwEvuRrA7M/QeBF+w/LT9kAjNX
XlLtFG5k2aJlKYvgOvDKzIF+vzFfGYMdaqPeBqLzGTxqZy1aQL/AlfPJARLfwvQr
p101vJYa2j/xO6D7w0SHrygqZxR2h+1w3xMDMyJx/1K5MJsZHzNNMalW9aC66ufC
fUc/gX6SkKaSC53Sm9pFG2nfL46pdd3qOCCEzvm/a/vTzvrnsDIR6cIsHDfYgk3t
YjEyFwDYeTob/VB3nNebvM2FUg9w/5yFwnIcMvKO6auam4BBt9PYS257dDe+DyBE
4Zc8i9qcJPLWGxaED5F9akEimPRqwscQ0q0hWJBRO2Q/LJNLyNOHHs7McZsqGSKh
0yQlpFXNNwDVWcBfcyx7bcXjJZLlw0g8sHyweStJogsVjsHB6HSOBuRQe9KyrYXY
KDyMpkWszY07i0a2SWzcMzqRbDwdMFMc61BD3ETbGpsrXlGmzh4SjxP3ZZ5ZWe5L
2EcLzY/dbAxEQYICcGGKCQlpZH3eB5bnNyqXqiKAmQfktjutLugRWVJiNlIbIk+C
tFPeSSMY8GdAwSZF7S67ZxlxirbVvhaZSdrlpSuYhH+VTfehBBcV3d5Z+m5sTvcA
Lea3IybNLZqoQU7b+mTgX5MBgIA9yUQfEsz9tWpcg3DK1FmH/X9uybq81mcNx9Cb
Ew5pNFCALmGKJbon+GPFkBjYMhfZPF0x1lNYTDBBjhxKaT7SiZEAua8v4z9LJMcB
Ubs8X3G+gLqBliptVOsrS28jyiZrJbbmQftYDUVT+6QQ9v8DFBxAdFH2Qti3Tw9l
6XXoyjqHAC1qh/plwd2Ahf+m7M+1RD5LkrPiDOE8slAZWiI3d0fToSkD6bPoS1Ap
WfhiolgD6/SJaFAI3tHC4W8qIU9MydY3wrMv09DlBooC0CG23w5grXEFwTBYTyRm
EzKnASvk4zHJ0S1n3cU8HsZBMAW2HKkEqWLTUu6jcFV0jk2jqo7+o8ljwf/l19gs
SlCuAktaIzT7VYw6g31nljJnuNuxU2wEHnkUv68nzs+2107TtNb2WziR+n28GYX1
PwagevoYX2lWCoWHa3cUuERo7AMJuucX6D4rSFZYSPLL3xeL9or+PITXLgZ53WD9
SDIytTxKN3Kmn1AeD+hDhRrQBVcXbABg9s8VB/piTLESGlRvzmzDbFjdhJkECQaE
JHMVziTfGVJ9UyRDL5bvdpU9SoQUYRLZGie1hphtmhwsVDsKjzZCLBhQm3uSBr5H
u+MnMuoYQTHjsvOhXmQFtizNeg0peifmLpYEho7Xe31eqEqq5elElg9iW4uEkHbU
wKTEcmSB000hdeMHzPBBVIKQm4ngyE5M5NN8xK/X3rzEpyG5P4iBhcLmUcVvuiJH
7iKJz8MaIieoj+nixRr85cQnJoBDS8EFBvsbGu98kUVYXU8dQjeSkz+/rLIJHOGi
Z0+DhqZg7hsAhoZ9K3EKdp33vCIzoHDgzOd9VGL/tyZ72kxZVOStyH5Vz2Y9a5Da
8IZM7aIhq5AYRwf8HPq3PP/za4c+E8soNPa6WXftEwNQ2eg7AXAL3BW5TGhHfpIx
8UnS8bXxXT9CdK03yMZdG0zVcLNHZVIxaJhAcEPSV2KLqgLAsfptlur1h7BjbJQo
u+08mBgEQlO+RKAqv4XjAy6Q2tpAURg6eUNjaJgP+tl8RLBwJgZOcQjnhjXXBKvF
h2YkID8VHYLzp6teARtYY93LG3PxdyGEUqoKQGgLbXltBdcOEVQXQjx/V4DVcJ5d
jSP2KSKZpXnNQeQ2zyv0z2sHwbQBy3IOAZu9Zv2gi3Gars4n+7uXy5vnvXkdTeEV
Wh01hiQKHXbsmgC/s/A91IluJ3O62VfrfrbyddeWJYcJiAiSCw4VVtihDYs8+AQz
nxITbKdtM503m/cRKrHOSWm254LRFlFIbYgh3GTxH6r7cJRB3B2SILZC/NMlaUmC
/0+KWWQ8jYMVK92/fOROLWhf97I6NbiN2ATnWrg4vMkANkU2tHuIb2MU3ZcFE0Ha
DkoSM4FnQlZdkh+MPBbC3ZitQbgOU6LHpMFRf58iNkHOH5KbfOfWDUC30EQf9HSh
IWl1DMsrziAC/vluAVPMVrJnKCs3IFNCj6l0DThxFj+2rEjOZmRx/1qSKt1SVUAh
QpO2dzdQvFy2Y76dvs7uqLxIZ3Dv1uQ0DZ2VTgmHUBLQJ5r7PzXGzjQhReJEHu8x
ln++0QrC/SCeYv/BdI5261/DqXGvuelMAt1CVFl7frEluHZ6H+5enzAWlvhoYQZL
rrlvs2W9zUsuGQAzrm/kJ7WQTvXg5PRSky7zeZt3k1Pp+rdjO2wT/hnqMFEdIg01
5hGVs7W/mTsQOQ5oBXLc6J4AkRkXRq8JfpFe6rO9BzMVUtsJuObzRt9ESqqNx6VZ
aYcL0Bdn3e6/xS5ISHJlxD0ur+3Z2ScP7Y5jQ4UGaJ1WSuKFbd+Gom2pU0UHRQFc
jj9orOt8WNGRuiQxtDP0uJadzUOChsl9R7mpw92cwDFGROWZvLXuMjRnteVbqzks
kg9W/6z6KXTwjP8qwSfVhCyb31CCpt8L5tgdPNuoTG5BcuIh0VIkFopzFPh1Y795
WPsAIiWdvnbh/r9TKuCUug8UDzwEBCZKGchDpEau40enw6SvoYYl80m6/dnW1yaK
hRHo67yRbS0tcQ6fxTDxUpW2QtFyw+r+hDUlxbBG9+awqsfT3pbOvYOxSoOXodHp
3yja/e/AMagrmDTI/j0mgxXK+2HmMP6ceeaWRynp34SOlUReBPJQ4S68oiSYbq+4
bEB7+WX9KiteFfWVBTOrCxlXnF1yiFYytA40HBPFg7UPrlD8XeNCNmAbe6Y5F/tC
mUjotg+PdHsXO8tcqldT3MQyK9JLoqb7TrBQW0g6fiSLMucjedVJQPzZHzvSAQgz
L+aqFymiL++PkP4PjApwohE3vJ1ljQXBAJaygaQMHQNXKVMTx17YFVFTFZ1fbX1S
V/5r0yxNvfjj2qXjRKJ7V24hIx8+5f1PnrRh29TRWQ+1PsCXvDSUketTZs3y0Sbp
pYLjesdM1Zm6azTTOhlYNFc1kCftdCEPU0EEyIkzhu1ivrPiLczkGjo3JCrqGWUI
4r2XBE8xZeZp9qHF0PrL06WoxheCCKONxePOIhCiaTb84qTKfIkp/d7Py+SWCemF
/vtzqAaH6NYDBXlru8AH3SlDg6PQaAh8OI5zUN+NfoXPZW0SUiHuov4p4UrfTcUt
+3oGvXICo/TKKmeGo6GVlO1XS2axI4+fBBQ8wnlxWYM7PiA3s2RDI3FzrOd7Hrlf
ko2P8cS8GLB7atAn+AGFH4M2JmLa//UhUqzU+cEjS9+NOhLDjxiBl1n5mIY3PPG4
wNXuM9c0U5cE91y2cElHmBm98ztPY/p8LOFl/HQ7gPqCTkHceewfj5KV4TsWxSZA
bypzqiCoOKs3jCDEJLUBCUlgAIO50AX040WtblVhnQTlrK7I2n+82t9Cyne87KWv
Gm8V9L4t39UTHYajt433D82K4CWW03kS4OcKmDggIfqL88h3posRoeLfhw0iKFxG
bLOxytMP7BUXwBeFdKynmVuKDMdEK4xwPZo8v147CXWkGD1ICKfAnv6oEyU2Njq5
b2AKLJnO3pR5cvuhtJ/oazviGqW8yQl2Ytc0plWwvCtvOUSIdRlsvaEKbmfKMvw4
l6OajetTlC6AVEGJPldZPv9bk8oqhAZogXJ7FWDuoaFzkaAvQ0JMdzz994G2I5tK
ziykR1IdB5wY3jEy98cSK0IJV7M9ZJ+PROsO27jsqiNSyt2ij384REPejz8gmrCg
jA+9thr9LQ1e+jQypA/j6O1gGvaQcta+VvHJIgxdo8WOpYnq96/aSgfFls90C9ly
ySoMU7zJcetfbLv52P8saB8Ir8nenPc7dtuQ3hs1teI3AmrnKiclYunSv3QRfIpI
LpHsE1kThMELxebkp8W77P9KYzwbY3/853NJqZjrUDZvEeKjKb0NYMbhfPKlSfUX
OmwxrhuBnFqDNfi7Bq2gRiIz40ExRk48gwLPUTTPPGR+Bc5kciU1tO+IabKUb00Q
njf2IRyvr6EFmCsLJlY3uKVHy/Td3k9L2fBAOioBwT6RZ9ctianDzAJNom4eGbnX
kDtxw1wh3IwNMz2Kc0xcBdqsIt7MA0W5H2ePNtxvSydazUE6M73/OGfK7lshqadM
/i3ZHL/JM0tkZDhfieX2NBej5WJujKkHLLKi8ZyZJZ+ucg6jYmFv36CJzcM1pKxf
Z99ptElx6CK0Xz2Y2GIgY/ySvt1wutyKOrV3tpf69/jjBncKUT5kDLYmTnDHPszY
TaIH3a4yvZqnkbWKRqOYZvSzbiM842IpsFXKoQjDjUNlonhZ33mS9uS0x0if2NQE
RozlANnnX9efq4U13iukYf5wm0CGocIHtNjFlC+VyQohg5fEAzpDw9S15zh8SUnx
DSNGpAorU3oRjsjTwiPh4/jxnuzjdAvXB6AaB7Y78oKcigAIxotPDAzJKaGaYWJd
MFFIzSl6Vd5zzuWTi0EwJ1Rg6sh/WvStltxo3Ac4a6xiURDfGxHBlxPAuHrgL7yG
KqcP91cjn4gRhFRmFS8/V/K9YvzvKFLcPLvQ4Kqsn8TaUVOCbIoNrjg8DMNc+S5D
i6hvWvAnohmTelXjvWnhSJCyi66R8mWXgOZD+DZ9//GPuW/R2rmGI7Z9IZddt5Eq
Jy5miTTNsdPcnx8cNXTlOh1oxMhWjcApev7/3mPMJNRBAkIGv2xIEi3iN9vYmb7m
+KCM7u3AXzf/usXs8HN4t+gF9WdVTjYqcmfKkJ+TFR3B2nnz/lQYs3da5F5riMmK
aGb7fIF451/bHfBoBJkZLhzVe6sHoh4teAL+Pgte90EwtVa1Xn+CLmmggP4VclrO
54TBq+3eH2FacmFdH7/t4HjOxEkfeC21wiN3kJ0zmZxOMMrFtPgY6mFHQLjJff28
x+vrDkY3yspMAnbu/5036YtiAyHp+CY1mw3XDHSxAsx6nBuuMFnd6ElUY2RDsuLl
tKR4lrrEAcij1Wm1sT7gv6oXcZSYu/JaXXRcjA1LnQCG8o8O0La7vFt246X5Jwdu
8lPJs07UYFgjfKGJtN4/Tno1mj2FdCg4zuemKuSZRdmKtabyUorbJVVElJtUo+UM
3ynZdx629cWiJciSF2U6bWb8IUce0O4LclSSFSLjtQ39AFPw34A7+nvwFj4bLIM9
OKhW7PgcEF68U9u6vgAM9uRmORxZiD2dvFsYib3Dz2VVeDkXx1tiyVMoKsDxMCRg
yEFi7aOiC4Asy6FZfhE6TqiovvQGn4doDIIzsOG06jIjuHCWW/YSz7MXBUdwcPVO
Pp8Vc1Q0qfpImPIgmunh6J1/Wxt6FMXiYf+gbJ36FTm5oFmBlb6UY+hr8y7/cXiZ
lHqpvjGB/KtRi5atDbnNO6elO6T/r0gQf1MmYj0p/IhnX7hrZ/GbHypO72eakRcM
H+t2tF4rDqRuJduphuuIvjUSiWigSj2pwk0RI2TCeuzGJZwMJohLaMYKJugf+2OW
geQ9OSzb6fFO8hZ7WrhRwYjKDc3Nh86i0SJhoT61vWAYqF9RL/+k4xdR/Db9ZbO4
YiSmdisDsNrVuZed7UrZuqEF66llwxXgaksvNEgpbIUpmOC58MFkzTK3bNEyVe2B
54bApnPAwdAFP5EKTlv/44JCMsUdndYEB4a38wY9wVOHhhyOQbSJ9y8KnSBXtwV0
jwGhGL6/EQBZT2TR6B4FdfJ8F/ty6hbK7bCpqOMCkbhBhBmQh+CxDpX/l7q6qbGW
kDw1GnpO9X40wjeF65WOu0MWY6yXyogBgwgz3s6v+Nm/x9t1J2yYCJEoMRn6Kqwu
u5N3TwzxhaxSdPaWUuoCFCg8xU/uBgtJeODLP/hRcbyAIBSQONMPTmAvZRlO7Byy
3VfwS+DOM/+juosDhRBfTSbuesE92ZBfRZAc3cGgwGnDmxjtUwCwlNUUTGnNOxdR
GzZHk7fXuH/8fx6SEDO2Hnpams3m8IEao2e5mO2IFWWxlAUy3Z2JDTrPerbz2L1v
ybiKGK00K+dukwJSlpfLynAa7o1FSfOgV+fKCQPu+uyqzslfUa+HDF/FTDGn/iLM
J+fZxrVotaGxunT5+TFSAcOvr3TYFpfBdVNh2LxK8p2vN+hPEUzyB291V2gYg9jh
WnFKLyTr9H6kHfJ77VR590tOoTui/cEqfFVl+Fck4Y3zmP9ivnN39XADpSwUjmmV
2RlidEfCu2rcK0BbdXSwgdw/XRA/88wwQCv2YKJPrg9E0CxD4lYc4WtrucKW67f6
0tTTqIFTKW7q85UrHipkJP2dJdiLzCQuscu3pfq6bl+aHVqsmXEkZsveBHd53OBy
EOWtywky+xAfO0hSURT+xwE6bBa8JThyh1pyXDc5ZhiYlkkjky9BrlerANaewmpP
eTurM9kMW08as4pZpEZ8oKHxXdUfVUo7q5CRwQpGJxizCZbQFbcmYIg8kX6tBPnD
U+0ZE9UXJbbKolUzOoFsq3TS56qqo7kkPr/MYn+t/+MJlStjLp40RraWPcKJ2khi
S8RPsAkaZ1iphNvWdMzOI/KobUb1+i7HtKgHK9H8s+gLNwt4npHxzfiXWVwlWeNd
DD9KC/Da2Fd8t0HH5ivNfu2B/KXsx2VRE4+p22OxVZmU1n/WCFV4VLxt5D2yee3L
5cZkjMBxBeLMPDWdcMEXQ6V9MslgIIs/ckspkI+oS1XoLs5NkiP88knFZoABwQ8A
KaKsGxVO+AgOAQjZJ79E7o8VuYm6yt8/FdB3tIj3ldAFT1U7a2TJO2SrFKmXa3zi
bcEdBRXxE7ovLLf3LcxDBcTD9z4Q7B8sqoaXh5tVOyr5IDpRqvGB3GuOJFGTw2mJ
oVLaNJWitvXMABRkXYKbPOlaWPPW94rjo41jeAlN9Ym1q3+JGTZNrsYukgQF8pIB
K3nuSYZnmg7bUViPWQ08G+X/vdCylvhuBx1leHAiK4Nc3RmTa70QgxyQHyFIpGgZ
++aGYQb5vJENNavSb29HBRGiYtWpz34dOujdPuP8u7tIDm4CuiApS+EWzmryOA/s
4VGstY6kZNmIBo1STST3W2QlaIdWHKR+U7j+c2M1WUFN8I35zBvrvcSBxGuzNw2z
XR9tkM9Io2MUTIvE5z6AAVL1YKYOIn4EjHE/tEvWnRelA2FxVQgWnBwSF79DKj1d
/4n0B38NkQTvPEAc+Rb6w7w4JEVt9/iPK26coZKXCh/y1enWPs0fjaGDgME094Em
hpkMOXayrtmOqISXQ7jzcMJN18DwpyNr3ZkgiZjDfLfk/DyIgKRRVzzM3Nzktjwv
QECpoNspk6MUA2mlrjI8DRN157T7m1QKSZhzxylkFuD1s+AzFFgEe1HOz5u3DGcG
SgV2c2tRROt1+VrTG0CcCkMjWwuPTBioFaRvdyHvfayLkgjiusPJp18Tgv09+lf1
S9nDdk1UEXrmE3G27MpcOeNZNq56SGcbAI1Mef4/BXpPnJcMvNS+6F6UTN2ud9Va
qNtaTvG5DO2ZcBYxEeBL0hBsGY6PDPzRpOpRGgtp8GwNGy4kuXTEovU2KVpqOTVQ
MbOqkww3RllMfKWBytmG0mv66pVFCGHgiepfiHT2C9R3VSulKrA2gm2Y6SDxvbFF
Jz5/7siSxQrr16/zwC9/hdfxjJBHM1nUby8b1hiSroPurziJ4HopG1aNesrLJ/u3
Oe4iG6zXmB5SSw+WAGFxG1v+5EVEHgAAvWCM0RRgteYczqyf8J5fQ/1wizRHbWan
P5K+6KL72qnGQnGqo6+5tag3GHjA9HOQoTDcVGEqtXfzZVKEAhlR4RJjgj1f87pP
LFJsBrmVGWNbdmQYKkGqVHyfoubdbmveHgjP3GAFdVVK+cBvLaYSvuJ7cjmJa1LU
v6uy4XOO6botL+d5XryGwhxvvl9GDHQHa7nEGNYS5GQv4L30Ztbh/XIwK+HQQVVP
qIziosaNTrz5X1PkDSHdUGDIbV6kKEeNs2eCpm5vwnd59pnS0jJR0as73AzbknA1
nmqqQ5P/04ne2Os+aeIjFFKQp077yFqUEYqAxFGprTIgU9x39hCitq6usZ+e3kkg
dW5tp2G0lLDSo1lXLql/FdO4Hv05QdkPDdPSVs5IDNxi6MtTMQucCiv8lG0S8tfW
4Lz+19Sp6lV/0tMdjGCMSWJZWO6dqldqTE4LcCKQ26SuL3jJnhVD7zMVbwb5ovSp
2XO0HyrkGFmDijNiWJfBTYAUIvy8rBjsBn8wpUKmXg2hMvXT02/60c1WHvnXMfUG
0dHrc8g6lP0OJ9xLlNlD/UilU+89sMupST7iQymgWfCraU/mK0N+rjfFlg2WwAdz
5udoAJkpRIuwjLDpv+GKx3RaaFwkDbL2VFqGesTR3JcQZ4J//q57ecVBU35ZKizN
ScVgdk6oceQ9OpwPOqKZQZXOIADDm3STSs7EsQCUuWNrSNDRaoH1ZMuxixtmuLxO
f9gIbNAP8V0ABy2nIghwU+ots9h/PYrLcUw3cuTgXioCcVRWpHYZzy7DeLJjaE0C
16Ovl5fBckzgqJWSag4rcf8DCALaZ0SifwbJztqqo37+ConnZJxdz5x5A5QpmTmz
d88Onzc7JmuBOa2JFR+roEtjoVkY/EciA0rOuIan++uotQ8Qs5CGWDsxtlUnj1LW
ths109CDAanigzRS1L5qsIcI78vYlIzm4aaKh8EXq1+jV8ZWL9m8GDiHKUOmuLQo
E0eNp7OybF0Kog9QPHyeLChDzLT0ilnLq583X1PH03uRbLEs1klvXfQcYFhVlNsr
wKERuWqqVgIB2s5yy1oDK6uy0qBbTF7/RBu2lfOwvD5gSr2HgtO1gJl6+Te+ig7/
bB3yX0l4IMdjWh/U8aqp0ciVQ478/6GxAlsk46wk9FvEBzNFE7sZ9n3DwCRh4zap
t+JrZnUD9nA7QsN/hgpETQtsrikJJpB/vy+mOEW6mY4umErQYa9yLLELA4+XIecr
O4kMZkqu3xuxYAJNArzdxJ3cd94+EOz3KRYWtOS+aq7C0dXMJQXBiurRLULJucD2
q0thENwrOMv2IDpLAKs0xKaQOV4PG5hV050oXwpb5GC1CELzQhCou3Krjd3rZngW
mabgh6b8EEKPyI/qAa+wNzyDyUMoEiPEwsgH8GphfppD1XME0JbJ0lBkQMQPaf7K
kECxnEwkzO4NKmdtP7EwDDq/41uBnGtjBAHY1UNmLos6BZwCs/6uk49EyxQDRbaB
ePDvfgHthSIjWd2xHA9NZC1J5xJQGGjWuuTaDpsHn5CPWNrDPSYaQ56Yrth981dS
SuvT03wbM1RHngXPQXEPlk7C0MtFC3Hhs7MofwMuuhgBWoD8d/5geH1Xb2TINE7D
eY70Z9zqd5oAl8J/ri5gWuUqYayG41dC+WJsEY7D46td0ZUPqBQ9teORwRLD9lyw
64asUDrg2qS+wtE/Mm3oy6/TDiib3dXcnTeDP/WAAeU4AoplbVAHpPGNO18sZulm
N6g2Da/mpWwAvTSwnJkD8Gwtdg7Ohd5A7B+ot7fUKwoHC7O8z4J4VUtuUghUPdob
JiNleG6awCh3R2yHv/oOkaBBYW+wR9TXpjLfZ29QsCAeZeTnxHW65P0/RC6j9SPQ
DoQDIwaLea+SNxXC1DXvLFvg8RpsaNreSM8mjaLROuNXNNbL7BJyFMCISXY1FtWB
Cf0AaBth5QdKpJz+1xjSAjxqYO9oIEXUQDufjNgNnQAU4BHZprFgSChLF5HwIqem
lXP35gWxSGUV9vg8mqvPtcatjIzJ0eXqWBr47IZWFDShWaf4Y3oakKGmrGLy5EB1
cukYVqNC+YH76vjW0N1OXBUEx8bkTtQwcdQU76PmudIT58jsG4LwZlUIdjGb9b8k
CkTqAmYooxrclzb8/T9hT4jjZtyCp84QuJMiGx5AgqL3rt273CzRnSkCiLWaWpHJ
bRtZM84lrMUGjxTorxUUqlKQbq+GVp7pG1LxgAUrh0vtpquO3zh9sGO5RV0f40j8
nk8aKLYO7UcLh86nU+SoRQHSEXJKwARhLgNxvXqmQ28996gY+4ZREKwdHeeaPo1Q
J+jID7V18YGSmjkNWaGY1i+ogGEg8LYo646A8QGCcOL5XtlhzvovcsU82wf/IJ8k
+H92zoJNmEpyHDt5+jYf0TnNxkIMDTy83+6k3gG5hfPV2olL58jL68KDAyJlQBAE
HEKNAOXzMvB+OguYRJVSfG4QoboJLGl+fsPPAFyng6rYn7DS8c9avIHHfwd5Tslr
bZOPVUiGjUKM/IKVTXe2tKYt/fjvemY5ZBtrIPlymHJIoSqpUXRX53RVmaXxuA11
vNPWsuco/FS5qGE8ckAnR2l2Wg1tuy4SfLRMIQuDdB+iKQqW/EL/Gvp+5fx+Gi+J
ZjmRvl33lgPMZ3Jx/oWSzX1Ypic9HPixZh8ab+Zsdbk8txivzGguIBfyV0uxVy4y
W5c8xFBvnmAGWCCWLdrnGmgoFRuJZBiO+fB8bDUvgTXo5SFta3DPNMvKoKBZnEuS
9AC/8p1LDLQafXhIOl3OU9li7o3N76RGozJAEbebIyXWR/4+4OZlW3kXiUSi5/mM
IueiNCVx0jcWNFHFwVJAc7/uUu6PrWSW07QTNMKlxFQHAaJzkNSCeXtJVtEc//TD
fWj2nJ707uuadKkW5h24cxlkWP0UZC/ZWPkB17LmLwp4Hm23sGHuxKM3coxi11/c
UL960hy2ia1/YANTHrZTTMJOSlSK5oPV9FwnIztPxp3yf12QJhP+TuBx3mUxi5zf
A1VbYwSVQn5cLup3rvALbDwYxDVSqn/5HpfeAYoazTEAYN2AjEWqJ8L4nMwC3jFo
Iv4RZ7bhC+JcDIODoAnxE3Lc5FIHwPcZkowf6r/zTVTqdpO7XU9rHDf+e65Ty+sb
if3Il/oJfnfyZYSefBfMhPghijhxp1sPSEAYf7As9msZxoUitD6MgiC5glMKejVj
bvj08Akvh4CQfYKuYu44+d/GOPwycQF75maK0h/f9s2CHleNdcDF5RYyV9A4/Bwz
b0CS+6zFO7GTqPWILCuSThG7uqxW3mk5qXOidQaEvZSJOF926igeE16EmVzreONR
CfAY792V6+xsbQnubVKA9dPcKpNF47eZmx/rvw7Bq4VvLvK49zqTOEG15Gg8ReQf
w/3zx1u0MxPh3n0oeHxInAGfYorgNYw7LYI1S5mj7v+DGBtQzxEwaF5Y7EbzjuBR
bPcJ5SXw+8CO68XLhUymdsacVdsOJ5FG3yEghR6pYG9OfLHQbf4BUwC9XMY7pVbK
ecZxRQ84vWp9nwclRfETQ5qz9ILxJnwayjuqQcPS+/JE5OjkABrk23Kv4M67U3Mi
QOyvBHKExSXUdTZflHmIXObnek5VByWRzE8S/h7I+oHn92AYou3XiZI5duW8qoLb
BtfYJEKCvIKbU1Rfa15P12bh3sBUEDf0zUfhVTHC2Ui6EYGzHyrgZJWpv9QKB8Ao
xX6aKQr5nJFXaCEs9zFBSSTnUM0o7XVMA0M0o58elM12lN/VZi/garrdGIwgwzkv
YkdrmvIkiWAXoUgCZVWH3LRwzZbNPxyDEPQdPaTuYCfypiBE7YYZJWm/bWEHrKFQ
xbc+2YSqasTBH9A4ilprW0NThejVfO7ks7Lp6dryXHA3x+npwYJ2BiLf87LzEi61
asycQbpBA1ljr9PA3GwFtSyPWOriiHwnbh0/yamumH1wDy2JaGd/wHY6sRsha923
JFcdVZhwEl6zcSXJRar26YLb3HPwszNaGaMTWK67I6qpQXUhCzTH/GJcxqXAJ8QC
QG0+WHSYzWVFosSFUQ9lVR0grtmowbDAyyE1GPYsN/m6+Me46pxlbOrbZ867g1JN
KNCoJsS9lXLkRT1Hl4tVUvGpQmkftLZ7HsZmdu65vKTTRgixFKasbYv1ApCQ/6kL
17FXjYaReKEUjGGE7nYqbr8Lapk3QyYw4rTnI39GmJH5i7nstS+RygPhkWd/hGul
yyniMdi00WjzbT76fpbkf7DPmBHmSUk/wKrits0MTrcWolbwcU3musEWdQmo8Rsd
TsczSIPDasPGj1I898GQOuwj6euov33AfEwUybAMH6a+TO7SNhDAx14z07PC4ED4
8rIoAb5+PADj2KnN9ULLmCLAXkuSJ6yczoybddEXYHqJktI+YRQU+cymVEyaDrlP
oLbT8eJgR2wjKIDdL1bBAVNfwZCUB2YXUpcWZHnITgdThySzruRo+BX1VT8UqtjA
rFjCgzaC5ypuLMyaR8Qbm2E3Vcsx4lPysWQUegCnEq0rgGSQXujgDtYVYK+8+C7Y
6EJhFqxj7RllPMHjxOI/1xnfQt2moQ7uQ1aErEDMcStFaMLY0cJXfEXOloAL8pod
zd9Z2OENP5S8f1mfPySFTOKNYY6D7bW0DAkbSL4Lakw/xnEiOFw6xUPWllpykTt9
dsJn1Vyha7xLCpopuEwO3vqzfL9+qA2oawrC8mecIJ9odYikvFH73KVBhyqc2CB5
KMnkNIM0YEqz50a615S85BltVEkCIOwLxDJQ+3HqUbv5kVmwievtfmXEsUToSMir
W8fe/zfxXA3GmEn3LmUx7FXZLTJsxxtkFt4sCZOJIvMS5awok2RrOmnoaHw+p/+9
h+mKeNVNav/HLm2M+QsrsTH0AvOnOKhPl9N1CcGwMAA7KRUSuUFOwfn42c0qTkTQ
ZKx4h/94eB00sG/N1f+blFVo/ULm0ExE9P7HCQ7wa2Y6/LNXP0mddKCCLKzxJpHT
tZyX8xeXsK3h+OqwTk3Le7lRK/yNLNc03LHP8TzD/iYGaKwPc+1tKBht/jdmpSAB
/FDciGyMvXnH2kus/hcPQTSbfs9HZyKxJXlYT+M3PW1zC3S014Mumz58oZ++0haS
2yc1RxdmIPjDVk2Mdw5+Z/kWgXa+FW/pCfiVPNLayUI5xGe3uYE1LmWQBuQEoGa5
OUZwhTO0J7jFQa2e3O9iVGdwl7TzcWJhDGPsB56FNh+nYvctWvJKG2C39zGfotJC
jMpQO/2TeE4btO2ba4+tmV9neBz7UPZLpSonZGb7kXfJU/FIwu4afbWCoBeefWTu
21FU8071Oupxmx2s7huSoMTF2P3EfixVagFBBUdQBf7mEeQjQufadOjHGXCD255x
3LdrtFPaJyJsUqCAAXr7R9iWuk1OgyhRfqo06e5bhYcLFknw1OtUKdxM0N2P0Jp2
dUum6uJAtyCUB2Gk4zutIoNbYt+mtLtIJVo7gsgs/wTeZNapo5gOYJ+vXxJZrNvC
EJiBML2PKjaIX9ACoQSiGODf25bfyYqdRi7lLKo+CRu1DlcDR4gaUVOqqJUMT0Fo
yY6br16xai35jn4apLkzFk6hCqmCBHFoB5T8Tg7Ngi+KPlGknrt758xpNLm4tt+d
trOvg7dNInNvTLqZKFjse7+V7EMDBV6x3q3baXmumAnQaw3AbhAOarXIXdFXy4Aj
CIHVwmleC2tUH51k8RzCiSAOSLKTxCD2WzYZ/0mYJHGTA5X2gp5j6O2gh/Vh/Isw
+0m+C5snuI+B9avduS3poLhOCSJjkoW+uLS3wLC5Ta3nUi7Sweql6Rn0pc28693m
Ev8Gev88TEByKimNJbd4gvQ/QZh1KAxqdBVUoyzHJ1CpgQ82MONhomlVIMlsdjDO
NtmUfIkLQNZ3vsYvYTG0IMLg1tzDz63gskJbYjqzzQ6ZqdmQ8LgXlawZYIALavLJ
XGj7/a631ye4L8Nv3e8mF044cDX+dkBSJ5cbAw5lzvXq6DcOcQoc2kd8Fd5XRGE/
YQvppZSUUXWXn9r58fmbN2KP3vxxh/lPObu4wbBtGZny5OD6kbORosCzdxXcM2l+
XNut6S5eTERibsnaMfR3NavHYHb5ikycYwTQ9wR/boR3/T2MEg3pd91UUwyXxo5a
FW12hVd1lwtAb+RmDRNcwmDpx3KSWSJIAx8/UM7TLbeSm8h6BFpIERS9rLH1rWGO
DpRBQHd3mTBK48OZ0uxGIxiKNMMBK+z+7K+vghLS2BVI/cB/yn2S64r3fFEI7Me5
qTccpPnN59JIzJOOlskNPf39/lkXOst59rH/HaT/0grUk0BqmotwokKgsSyILwFP
wXOFcgyWn2FVHWvDEMXaEMtIRNYft3cVduKohZF4ytJc7TWghlwxrMykGmdqquFd
+7rBhz/9uTvyMGBURRxIcU35yMYfZ6BMiL+k1NZzE8Pw8Cbh00f7XOP7k1zKWJZy
DIRbMyr9JIbn0LH8IgB/LXDehjAwr4DMJrVcCzJwvwjfoycgKn+WB8arQeqpUaJM
U095FdNDPT2O2c7PIkM0LjhGwcbTl3SCh9+htQ0Y+KJnm8RKeeoELGhAVXcLfQER
4sGUvj8dnFSAv0AU2lbpuqZeeCFFPHrNcj3D/2YcuS/dyeoVauPMGCfyz6DeF2P4
eCveQRKgBd7OtpQN147IC8RcJpZRusBGNJwFIckE1RZeNlWvT8LfhO1O+CjAQiSk
PONLxcJ/fgcjgeP/v2gGcf0IC7h1Yp9LdJ+4lC4gyBA0gwRf3F52AkbaTFlq55nQ
TEitbdAUzvyEOvBnxln9ZCQw5eInZbnTTV18NFp5wmvSLXeEZTldHvCMGAJ6J0Ki
q9NaNFSzalin+NK+m9KhceuVtnnixk1UEVdyRCEQvKwE3gm19Te1niDEG4lBTfPS
j+7cLNJhpGyeonXmwL1K1Mg9UkToJR1CjnwjtaQhp2XqjxBwxbDnlLXKERCcP+/7
SgjNkIZ1MVJFvWni2hx/6Onq2iCR58WAtppg4bMa1oizOVthE7uWoxBFSoU2WL8T
kaxPeNUTaYyOcwZYEqicAkk7UNmsgM/rEjMXIMOSHiA0TfEMB65Stw5Tzy5Kbfhl
i4foLWveOk2qB2Nf5mlwkcM8RZO4DrKwThFJeN/jLntlIDJWWgWxmMIKA1EIyQyR
40jw8HJeP9z+dMt0GbOwuNw4eQE5HC/0XyTkY9J1OOH5fAs3ZPFtGSd30Kt78sfc
SNx/Q0RQgXTJr84Wo1MpP0+Bd9Hyim1XCHCEqoDMYSFVP+KXxpOgIigFZ+suw6A/
kOwK6dbDrIplg33SeR1qO1YYKuxg+Rv0/KyiXtgXEgDpKazk+ovlucCYRF0ICiQi
BjJHVLLYsu21fds7p6yb0C9GPIQgzSgRel7B8q/jsZCwXSyE11QJdW2DL0k7SGN2
XCNLki26ulyPeopBTSE/DLPEyimRrTNEiMts+TqrwQifw53GxE9KAwJBvHQ47MQl
YCzYbTZ79NSl5Ql/SNMyyyg82a5kH9fjX7qEEkZ1KxmPUkJuUG2Su0jdXgIate2i
wC/VfqubDCEyBsDviPaJkoPpKYecR7WpTLn3Ze/AZkBP2EfAyzFbdBKuDFphqc8s
AdhmBQiKmSbo0bSSzW0/QS50N+P3TdE0i7qtqH9SQ33GhVWTigLwiUo727pr4HN4
+Q7IBFSzALMWkcGvmwGzWxEJnhJeKoIrqiyVPIUyMTrdboCjaOYeUNarl9R9l85n
/r7ZdypBSaRaZMkaBniCUfLmRqOzyjjA99MT6pMGnF27qs8WQL44rtCbt1wPh49l
QxPHDi9V/RqoH7FwTDHef/ymeUzv4RPvv/nth7blbGp7LNFsSGvqZcz3hyR7mw5/
HyTEclQK5MEWeSLoeixnagSGOxPrQYD+xndNngS+5ifrqDE7w/Y5xE6dt3RAio22
VE6gllM8HRZ313p2pxIpC2YFAJLq4rMuWms1/kgtljSLGgbEjkrJ09TuJJSoLeE+
PEFZHV0PomWgT9z07z933DNjE6YYHJLQdauHiH1sCzcLH3KA3kWIsDdKWTSC5s6A
O3kQAuATuHJOCx1MtjTV/PIr5zDVx1en55g3f10heJM9aQOOlOexvL433haQRjU8
BBdrB0+nBsOusHGppBkH8oIlLECSueuE2n6Z2nZSR2Cn1t5QKWX9Qw6TDrQAuPPe
WXHg9eKYhR7C14nWw+520szL7kL+CvFI7HnH7n1uoKwuOfMgozt+LtbWWz1Anduh
iE/DN/qDTchpx6Vf/ytDG9qkY8l6GL4jrRXzWX6VWOfatSi3zpmiynZFsXUhBAQR
MMyiOt7EpPETWSHsWdFNTTLbKMbGsUf5LQyTgc7pWccqGtCcp8Wb8JnW/ndYCmuT
5YS5SAa+mS4iVjxchm+pWjWSOiVFGW2udpSsUnXoDAlzRLU4SRky4rq5bARglEGM
KA25yKgFhnxJ0PpK2kQ9a9fAddtCKfs+1YRQBb+2PHTyeKQgBCE45V5ghZ8cxh4Y
c9R4A36ZMiZOT6HVG9WmlUaBrKc5i1VYTMb2l6BI1vUna1YPowA0WiIDRfO7t7Zv
VZdlBnp1E7zhBN3DMQxHzyFW+uQXIYmgosWfVEIDpbJ9WbXUzucuQQYk8PNWm1Y3
/pgBeyY/7i61ybl3b/IB7Nd/RCkPXKTnaGoz4HrKKkD9rMZB6sdXs/hXw5G4s3SE
35MtzYC6LsHBSLlFU9i0ibYpBSVkomW9Up6KKpZzcjLStk96TL4z6zOg+9ZPNJoG
ycPoMfe+335/9md85MS+MU3SdIfcSn2q52PI0/6qHqSVATrjhtnaMEHPDu9ML2t/
JRHLIHlFlP8AOBxBrkMTDF+DeLy9YKUJ30vqgBV4LWIqNNRdXL+tdPoSZVNXowAB
xN1R6W6wl7TwZCXthZ830AMB4IqozHInlWbAdcmMRJlczzFfhri2jjXi6WEyxuUU
6A4vygW7Bsu1x4rhAtvJfq6pq2XXikZspazcxBXp1fi+5oiWBwQYgEaEIhBnE7Y9
W2TgHDrHnPLLhKGbU9YMTbAGHFl2iUFHo6cwSFGuZdQ3aYNAyA6HJNVFnBqLkRM7
gde/Lob204d2BJxpJyUuXAU6AXzVgyUZMp0ZHE85KerU3gFUWTmNrCrju3ckK1EN
yMI3M+w8rQ4BCG6uQTrtemm15v89GoWWGLWrUX8JkwfYX+oxCetSxpWshEU9uyCE
jZ3MnRwrEMVF/zPTkoW3IOky1i8UKiAUiJb0X54+wfmWHKGJDXkXKfNAXKtPsPdU
KyDQY0FhUdICoxcgVdzQz2wZ1GLl8EPkBuxuuWojcYEKruWqbQnstgf+7IDWhC0K
y/W1busplU/elUC4Ims8ZkJSjC/LYfwFUD8gsEpBeCEnni7VG2k9NQ2HyyipocO7
uEHzQBliApSyeaSp7aSVpOKOm37Z9D39xfSojkReOPn+XKnnAZo+Hdse2aE4ZCYc
8LOXjZrG7OnKaXmcbtKcizkosTvpBrEDdfn+hzZMjyu1x+djHwqxeQgyxxcYTBBw
4OGn69qfFSyK0Zxa1W4izOSpIzplQYhbxPDoDByFl7F0TwQ8hKXSYCVWbjMCz0Mk
MRX54ZEvLW/1OttndpsxgfWkSt+Y5jBXRzqMGDZqlPVAAnGh8qN+bJWu0lNVhTil
XrTycsmDHSl5e7Qq166KZvsGaI2M+z5X00Z/Jvv081pbk3NKboHMiNtNW3ZYaG2K
bQlmhF0wSy2w/Z8siPFzqfStMICTJ7dmnanhO8fJVsTYHAy/Dir91VZbfOfX6Hgm
Z8WpxMDgo5pcHlrlW1d097iXbfZH+KyjE2RVlitdYfBqOMYUSdEsIZ5uUYjjskb3
kV+OjOcCvGeK3nDMGgYby5tgI2xbjiC78lNj8v+BjjmdhHyUKnlUjyr37j7M4FX1
jdSE/6iCtBfHjFJVEpdLENi363HIyAGxiZOdYOeJK8WT528eg9Ad/z8M8YAvyPsP
b2+ERLyheB/8k/ZLm2X7duaFU6bH7WENotI9jVOXwPK/k+qkDAQeHDTdZb2KOYVW
e4ataIDL/Xu3Y4U9e71XyL+qugfXGS13TBuHt8ZtIuwkMfpAogk9uUANNDgSIk8j
VPNgyM7RbIZseaSL/O0WG1ZMI2h41Ae94/DAuLTsjvYIp5oj/I6TRzvrEDAMzoKh
9TRMD3/Cw5jbiIxTGg95s76mEMz4AnsNS5nZBoMK5/GDmN+9HHJRiIp3g9K9JDY2
or5d7vYrDiGqfcz7OmgVjCqRvZOOpg866OMeE2N7lf4/vMo6p6eDvjOeV8n5spVk
6yTOyjkbMBHIGZkCy9T7ME+SwkkvaMS4pkQXBnxVZycCTKrt9JYyY42s88qGjYf5
G7H5T/4GHzDS/HQv2KE34kGvfTaj5G/Ucjhw4FdaIkRNfcCkuVkFZ8KBBorfNo2A
aV3T6fUjSZqRIv9W2siyGxkmhiIHJZHxmvgfudrhmsVsIiac+e8zy6NPgjnGA/P1
Ur9FGRii6lqEoDeErDpmJYL4jknR8Ak6vqDaNUTNaXmEots9NBGQpOqLl+so5nZf
Upa4GJMbYvxsrwwy6Oa6tXa22Cu+lPgYgfeQIoOLsiQzwtiOb/cP21bsi1+pPWGF
WuOjjfbLAQ+S27lcsasvPdd2CFPFjodB74AUCmVccvPTmgxm8T0LsGwzCl7kHmgb
4aE0MHUm8d4mULpB2YKdbn4XphSwgysPAvGbRqSBWZQ9JR+/gEh3llV8H5I9faaj
b4sEsxQCqGV4av2ZiAOk0TnM+T+0MXcxUVPWkse38xv9FakC43XKPr2kIVie86+v
nRGzyUi2k0TtBi0sUFqxRo5+MAnE2MJzU5Z2DoIKaDRDgDPxcdr4HkHhyY550cDK
irYeur4rUC+CKmVXWwzPRm++KrPIM8XXeEmvQOI7Mi8BLgtTKKwktIK1PgCQqjPP
K4eMX8jViTSac6nml3FeObjJImK9w0u3C8ORRd+Qbp7bTYyrTDVeO68mbZDozMJy
cSjwGKIGu41vkGFBlepwOMCLR14nNRmZIrb8/JyTpM1nzJvAEyvExmx09PaXT8vb
M4AzLykgBoTV7yMr1w7Ly59HbaCC3i6092yi4P18vLncWwJIu6zpvznjXW+0HMpU
SWb0HoKv6nqTQ4X0shd5AA459JbqeygdpJQkx0N/IwLbBfuOquToh2ff4zOjsuSI
ppXNNCCulxLzlEusJvySNeVKWk5wmfFBU5LrUUR4EpR86n3EikMJ2+iA5H/P50El
6V1elvopXftz0I0tu+Hz0XfboZH+7PRX7IGIhH3X0GzvKyvHWHigTi9BsJMhr/l7
M1QUxBGotMgUcF3LDhxbY7BAeylIA1LLi1GmAl1rdQ33ZjgGs1a9Ta/v4yC4x6OR
sV1th/LHQC/pYj8E7HNvsAF5LhHUSH8vq8XrezF3EpBOtXuqDlx9djb5LpdfIXNS
4j4nwl/ROftpYbYYHcRgmhjU6CcC6MfJLOHDdKtd9z0fKliOsek3GUmcnVwHBjEA
jWn3FZ2ZRxqQRaF38sMDdA8YKA1/G09v/T0qc0vFDK+7MILG8VKE46uQ0yXjhOL5
Xw1oWWq4OYY9p37CZjdOVDBsuOJLGNZ2zMsLu4RFA09TbdqSXNMMZpnYw4IHOAX7
oIMeebEuFyOKYVJtiRGY6cG+d3zW+yZ375if1tiHujrd9t0DglfJBH8M3ylnq5wz
ONmQ9gMch1n8/d2isHUaLVhkMTtaGfFpo9ywxqRJY+miN1zen/4/12D4ttK+VCgS
wYsFSr3MghzyVt4nRNJ5QKjoWgDKaB/Mf37OCtBrryTy2PIQ50FfGkZtTlz2rnog
SdR23+Sbc1a+CvC5fld+2Khap1LaBCaFrKch6+j5jh09g+imnH/K/fuJHTRlqK9P
lrljtY7mZTLUxr4b2CoxmGszUAtFcnbfTcYC2IWkIVsC3Eptpe3t95Q4l31g9DHP
hqfDNj6yQuoxqKbUKJfbL1vLzeCvmiaBkByijYL8UicbXA5a37rmKpK17Zrdavpm
kZVc1DSOHRJJ2ATYiV+6kks233hXDUwY9/ZxO+hddElRGjwjyyCd7enysjGl/gfT
RnasqhpS6sb2Fj9hZeovHrQ8XYWLQ1+stjLawPzhusg9vlRmnhaZTiSbZz8YwVME
Nw4gl0Vlwu4IvHYWpyjuYnV4z1I/lCI0hgUmCLKKHgZ0i0J19o2XVILESuZPItWM
8l5obiiuxOETOLtY9DiErw9uhpcyQ3zhGCoHfa5C9ZODTW57CcfHzEnh540l4FNe
KuKU85vT2X15UASANB8L+3KscOv9+IK9ozZBnRBRX4GlMES1N3f2XSSashnGi5Ex
X+0SrnQrEDjtdePiREfNjGaAOtzWlQTs5DToiGr0Z+jbQHU0BABMUh4io/4N7KfQ
LZ0BSxwSdHX2ppR2qjleNcWd6NF1FOzGQGyUHDI24DUVDeEYQHiX0TfuoHuoADt5
dqdiT7N/nslDrshIGxHZBFUXmQ9byvrCRFeY4QGv5+H8/2Kk8JE1SBWFksZfh16i
PUjXhn6V0KygglQec1rADy5XQgs8cV3cyiNQB78CadKlj8hv8+sUpwKpFoczk5GU
/MNgZoZprTdOcH7+8S/wGxfaKwfX8OE7q77KX8WqeQNWZu55zTmSRHjybrSDncXX
pyQhTNlWbu6zjqQf50JWZI7GEvKRsNzVExY3DP7zfCJv1H9Na54i5W/u3e7vTfQ2
zNqYvOHhIKJjNk0Bk3lpHi2cxWhKzurYoKMAUJsb9xbnllTcMmk1WU1Zww9W5m5x
Izw5+xW6osu0aVLoku/AI4ONiQS9FVq53Y5uKgoZIGLMH08VTSSU9RJMQZkrCSH6
yaR9jvAnxxdeShRBnQzRt1vlieI43nZDJvUz8lzivOgQdiwsM0aP4htarQ44p7Qh
Ib1i3tTr28W0SzMLF2cTq4WL+37bYqadbjRCDIhFBKTStD/TrVzusedktnjFtAzk
JX/8ZAy4DXE66JijOyf2FfaQk0Ytn4C6UiAGu/Wm5DuR2twQoSuREug75LRj8bum
AZHzi/DQN4XzHYDFcx621hpkqBkxmWC8VWvYsSvUa0+QaQIFlmteiJ35S7HXCgan
OGsbl92nb14xobKo3gN2NtFsqC1OkxCB1fsY677nYQ83g7ldMKdfOaFoGlPw4Di6
jyD3gxP73p8FsO1KZMDjuzPjZGpTUOcN45VqVIoEJYXWaE+VjzcCozpjRmoMiqQ+
OlfNJJYFexQrVaclXtu//ZQTi3oGqUVVgSwbuILRd1saidXaxCXV9zYSxeR1fFbV
DNWLWvevBgecgD51v1Ev5q72b1JXIPcKYObOEbfmEv44v05BI3uIkuT3B+LCiokD
7i7x/GaiXM3MD2Vf1McADrrMTWoUlrCTntwgTPDlyB/GXGMNLSPMEJqaVyRNlmVV
BVRHppCpDmENimiLbijiKms2E+l5FFwkzDLYRAazLJI2f9s4XfzXG1gzuEtzEBI7
Ja/W8kBxnmDlAhiLOOX3AI9eFfUlMRP2cz1KG6b68QXON9u/5E3h9a6t2mZUgj5x
3YcYhhDNO3JyjQ1/PY3gkgAQ/wdBNZ3P/audeFaxB06aDAbkJULFzFgEiHLLofbd
m54XKKdxqd5rHFgKdkMc3YmwLtfNPFVIiHEXi678SJbJa4F7bTxRwG65I7IcgPQ8
Mpa8I5Z5et6zFxYfbJ3HSahKqdLQ8T2D/juPoSz8WbK2sircaJlyBk3u/XI74x4d
lOcg8C6VIN1mz0+YLKW43uttrcuwzo2hG8xMrIC38z0ED+Zh5BThVSsyWiGgInBy
fGL5Y0RToNy1XgSrtKAFCGAdqMBtaMeDoeFzDQL4RPL4Wq/lw3OnJ2WUWOrEn8xS
HobdyfDaP9NgWshJRhLLKmRJ5JXTvK2b2YwQfYJpXaEGuNHbMr/Uyqqo9mEE1rHF
yp1L51UJTZSPE99584UXTH4ZiEKrdMySlNxHaThnmxEb8LBLW0NthORFIxXAIN6B
1LYIGSafCSQ3mWT3R4ZzqNNI6iD0rFp10rAW8W8L5Y4mfTurRCeqHx5ULXV/Zox1
wHF66LrnPxTOSgQb/qYDaoM8RMKuuRswNlqcZt6ESuPHipKT/RIHrv9ntUO4zip/
0gnOQ8pvrPJi2xvUWBObOV3zNtD67gCR6VER5qkCt0O8FpOFlhEAwAv+eaa0XjaZ
2dBYYGyYf1vpP4PkLkQVYK9osMEZW+qTrtu+SUBfyBJnsYdosg+2vB1g/30OIY5Q
BBV/F8I4yKXoAOqDBMr6z37XYpQ/UgH6u6WsFjdzU10DKlspd1k7Mi2GAAx/omcH
4KBYtWG1yCU2FkMTzbuPSZz5qeG+izV0R5ZwIdLEvlIvLfModxz9lrdcZn7dHMjD
H1nw7GcxiSBVrWAwuKY1lGH3GXRSEUeHVYcDDbxwLjhmsDHiXdKtOXkX+Hg7mwGc
iBp+8LMq81rREWv073gRDrZoFflD7Vr2EEhQQdd821r9u67t9MmoZrVnhvGjX6qH
TboVJglHXAjuCNhpt9Ju4zmVPwzjN3+qEcQGJWXomm5NaXPWUyAXwiiv1adL4fX4
NDoF2EsRu4fwXiL95jZNsG4/vB9P3ZwTvrWgyZFMIrlBhAB3SuY5yiBK5oMtW3+m
ndyQMXy3GJnzM1b1IeN813XXAimfUltmMlcE/XtclDdLg5OGke8Aoad5KpW9OtYS
qYSlni18d9nxRao7uM8gnFOSDzjBveYGaE/O2PTYRURunqe46NAsOTsNZH5RHtxf
qX3wwKNxR/DT9JKVLVzu1BubJShK22f677PkKhxzqr5a3hkMjQjSc1gNplixFkad
a1bBuw5fPi3UNcZ00SqkfwrI2tLMaMDO7LfdKTz0QDxPWfAx1tlbkNyvxZ0WOfix
0VMQlOvqmyEa/VHhEBnQd/hYL6x+DbQaHxIFhUlNisBSymJj0t2XdXSni1h2iMTE
1wFjdF/wZbDbpgKX1zjBi5Rh4L336+zB2yPjNtTEZZNkc9uhVoeQIoay5qZbQmb5
3XxeoNEelEvlzXx4awRBcVbiN5xNMtn9cGqZ1q/LVPs3c7zYE0nTel98k3kupfYb
qfop8RnacTc7h6WhrQU5vv4NhFXdcjzcjDT2TSiGD5y6y1zzG9bBaaRXWAQx9WNy
KbXcwf2enABHU+oHDcBy3kbanzlojFJGfKWjUn5mT500ueut5Gaowt3tePJkmf+9
ajSpExF68sCLBoSlCtYnF/KrBiZMioTzdA+ev+4dyVW7dUjld6QsbwvFrsDcq3rE
W5bf71O4B1K6RQci9sbNpOOQYZix+OvSBaikqk5FndcE36BVp0W9i4Mo5WweR8xo
qvY2SdFnGm14wIw/A+zX9cwVmHJmig5vL9bx6Kn3VEkakPoEfkKTcnoZBZJsztTd
p4f8UXgsgSg8EpifXUmsxJwPQw5mR2JnezNEerqylTQ0ONvsTrDggGJ8dYMwTrbh
lAbLzXe7NU48aH8tNoTMLqlsAEcP7pZS5GDQeo1yGJ3Tkbm1a2Q7ls2XH2sAFIPC
XxCfMliy5Jrk2z0EpyL7gpgVWzRDzLQimoHFrjTqOhqoOMq2zmdbVd8jqZU7uHsH
tEI6w6+eHKUS1jdZM7Ei5ttGoOQPO5fml6frQsm3mthK385nwIuihwc9+wejLZHF
QAQ2WsHaH0GdtXU2iYOQAkQsQ1iQDXMNruSDfV1LJM6djKm8XAORDjTBpzbRXvQi
XwgH8OD1wSv+b3wsmQIcIpAvMopzt0MBHOlpQfb5DFozu8koaZJsxIsyRg+UhckQ
QN5GQebHn5Gju5uwTm57kfTASs/fb9nvzBtYvZJQM6bueRMEC+AqBnIH/ctGa7qD
B3JXVOxKo2KyYTsJ3pEsl8ymy7ux5eHTJ+EQ5hZBKoSIi+cdiYgvvjWdLnfStmaX
SGXaQD27S81m02PRetYjBXRDE2ZqnpdunngzO0rEjIepUhN+0Nu1oBC3pFsnhf5s
yafvnaNMTshtIGm2JUVe8ORk9Edg2tS1aKWSweHjwsZi4Ix3q+xnDqd65SfZupRv
kFI0INXE8ZSA+XMmRfC2pmDbuptcx/7KoiGFf5EuAAyAp20ecY8U0NExZYjWKr5l
yTQqk/pztxhOzIEHtCT3h9Px1yCcIz57OY771Q0T5Ld5rsdSy+RMGD8qelEJRBtF
yXggxKhw5fxyxTV9E/WeAw118HfdLGg7fElb6H9L2RIG1Zxa7ypytA1aB0WFCkRY
OAvy2aR6dUxC6+tlnxU0W+W5gQLzPZwXYQAn75ifPe4gmU+UuxQNCQdLJPn2fpnc
C8KpRzsdtOLdAn4iRDQ4HtosDRxWsgt+oVekO12tK8oK4ChsFIYZ+IpFd1pcSia3
0jofdMgQZRBRywV5lLqvtPNJBEwt+F8y/PlIsKfrJrSx0/B8dlUMtymxEQU3Xu0R
I9ainSF/FA/3lQQdhhefmQ77btKuwO7aGB0R1Y0T5saDnPHyfOh0G9+QM1yMaSyr
Z7PYDSwrwB72p78xRHPiXcgldj8twKWAmrvVoCN0NL/ZQvuxiJzF8ZYp4bIgQCSx
ErmROCbHmXKG+VDKvS47hsfvciFGXMObObeOkKw/D7GFnjWfyJ0aKrX5GyR/Iarm
xwTrFAWSuAz8I/Oft9zbhptrPO8vDV+w+8N0HEuLWsl1xtMNLu2aVQwXaboEMGFJ
5nbBWjk8Og35RMX09VQzjYjTMvR2YqXacuclpI7mryvSw5y3tm4VGESCYuid97wo
Sszd4dNt+DRK6NbX9RtYApCOnYmQFirb327nMWk1xNq/knGvHPHk0Qd5YllTL/TH
m6+DfTrFALbHOIk7nVk5AWQDRRRjbdpBoDp72iLqTbjV8PuyxN++/5gyBMqdJ2Dx
CPfkoZoEkI7JMR4Oh+wnEd6uWYIkpLC9Zoxwqnku5l9DmH2MOxjY31ZPEo9GTE4e
AcbzKV2CoBZJTIhCzi5ZVM6eyho3u5XlDWy7742R2BD6+JOUN4cKcbShPH3qJLOi
jjYeNv84mY40V2d+71pLiztiaAMmIRPKQukmqPmaQ7bPpN6OMEODl0osMYIht3YM
Pyyhea8J7YQJw62ZRVdgLjlbe2tBybjwz6wSRIJOuSq9Oa2AeUbUpj8M7y9oU8mD
NUr6VCToaGqfwfOxx5SQXng/f11gnp9o434HCIHy8GxXf3ysC6gRQ34+r1t28NOH
lHR3a29A+6cPoKT6msPxPzeLMT42+EtPXbvokbo3ImOE6v9y+qk5PJ4p4A84deYF
8UksuOcjgmaz4H+J78DayXIk03UbQJ3R2ZwlqBWPxHKjPJ43nBlVdUekzEbD732W
xhpkaeerzfW4hFW/uGi3PZ1nkasC19BgYFmuxROM3uTxXAn3VTu4mMd15wvrwYs8
obAE+op/f1AtnsTdjPvX7dA1PLLL27BNzZDqLseyo89SL4WWXjRa4qhflwHPPD/9
yo7XKlx1GQMsjXob9bMV1EPvps3XVkRwUoahK31bv+iPXBeWLvNfUcfE15ZPMDpe
psc5FeIEoq6O44g4/3h53eqQYLG310KFk71N66cSgkMIeEzG5vUeXoq936KkCloy
OJDby58tAUeBovAPhXNQRfIuYtOyZTezCy/iPmd+ZcDiCk49MoIMrGxLWaoT9ggc
7rhq+zwDOtRP/ThUhLQ2jkUvBAYxNzkSqM45AYi+ZY78UIcxpeqeuVi+URYD6QsM
NTtUgC/AV358MUiqIeoElOiU4HpSRkgzeMcVo9aDrYSY77UlBEBMeYTncvlEbpR4
cvmBj5OyNB3dI/GvEb0iRn/M1nho/KKSenZ515h+RLGefu/GJd/a/+qWW0+qL27h
EsDJ/+EeMfW18Fn9lQJaldLydViGhzwo6rExZk+4wy1Iv5iygGGQxrKHcfGuUPWb
iK6V0wwYSYpn1JN1MAaY0Zfm+oTaPQG6lc6Sp9YQzie9k0JD26B3/Ji8bfinONnh
6h+8YVnCnLGgJ3Q0aK3VAp8T24U+sdUIuSF1jmtQFJWGkU8Oki7z/Q5nHilHoIwo
SdZuhP442oqjMcgqmuypuctAwPjOEl/zrfhEObb42QY2ORp9BHpe2Xfvocs/Plk6
LDX9aYdTOubeSy1KQA40+SsazwaGllqPEvTxTDGxGP97oypqZLecF9aWm3dIK5Ss
G2e7COy40hZYLDNx5yAJLaKi5f7a9gtFTowQwtaFRq7RUKWbhWsQfChSiuOITaux
sQ4SnZQD2ZEggB+gqx0If2VyUXQb7QialROCua//1p8Jw/fnAuhsVOClz8IUbxti
kcLP+2XPWFJvhXtlhXM3Eg9fq2EawN+aUpqVj7/QQwa60PitUHjGMDmDaCXy+Jm7
LXUq/wpWzpsLs29Hpm16TtiX+OIy698woXs/x3YPunutyfQgrLVtdzqxcKIQgUdG
lrt+87BVnBEJtsZvVsh51jAKtgCzlMX5nNlanSYNxMTsii19B7BJhaJtiPZbV7bk
bzeQhq1W2g5ijA8Jl4Go/8g4IPD4yJV+pqYgOxzOBZjCKgEPT2bBDfXMthYIJcHo
wU9rKkM07bL9p4jqWSYyB8ufESOyQJz+yx3K100UkcPr/IN4M3+F/soTGYScK2KR
qXJreMNM1tsK78lKM7pJ8US7Rym/8/SXyuI32ncPM8abtKwL9jagzN/IOlqQLLMb
zqM1MCGyrgotZHb6jFobOaSuRkZ1qyWDvvq7EXDQ0Ca1ErndDlhApfwEH6mvd0UF
/Bp1S4SAClSKq3yDFRKVhzY6kQv/xqza3IRiDXY/yIN0x9o4Lhi9zpg04oMwYo0P
qTMyQEKYDX/hepAV2l+aKxWprLGioBWDBHRAC2KqbP5knnbOfiIShBfxPBS6v0wm
GSmB/h4YQvt9wwFlS7OucQ8ucd0po4ZGrP5gmzNcOYNIIVpytwo3oEvVSNXeZ7RA
dIySk/zBD2S5hQLcWQjI7SYopAtA7dlbDfZRYB3f3BXmUz2oEkf5GlsSUFxsERwN
jZhvG8uGDeTI72uLP2C0H3K7kYxfhGqlcLsq0rEI+Yyxwg3XGKVMwxvsUOA8+CNy
M2Fk691/j3+HlEQWfrAjaJajju/AwHXvkyvgFR8PZ//+soL3dS9NKTaCYla7ZI7e
5QVm20NqQSHsmAVecyoCBX2MizeXg+8BEMS9SYeDHcvc5x7CxM4C9oUjMPU4bFdr
285tVXAQ2zHsCRmLshWm6MvYCG2v+I81dDwebv4+7to3/yReYgzyg/hn0Jb6qQ+i
dma9YglOy8AtL4pWJN89qWzyHGj5NDnSnhWVBSHWmNJMCDjTIGjw5g/vqt7GlPRK
xSgSrOuXS6fXjet0jJ1dMH7I5rgNsgHurq8T6mIXjISt8YsPFWzfZj1s/C/g4hw2
h4mlQoyhfKreXoBMHdH6d0E1KggwI6Qag0X6NUtnDHErfvdnui7sJP9PYD/Jstzn
3PonT/bbVGbb2ikG3r/bovFcBWI2YiuupIaw/T24X6E5nEgP4FsMdNhxc6O8/Mi0
y7DL3cNtV0up/uT873oS3Og5KsICDfCdBrfs95Igtw76F46gAxVWUhgoDEQfw+t1
BkeFwEQIWwYKq/ZPGVD/6T7rhosSvNvAhxkb/sYRhX+GL3T1Sox8o5euJdhRVooS
xrfV1gLal19lrDDXeFNo9Ts308NFGzg3KOAoblOGCWBZTAja1NGAsgBDu3Ga+SkO
qbOs4JdE7C/EXVAyEGLi7Riatr5incehT2J6FWWkvi0c17OzWlEV+VWJVpqOmIFi
qXnKXItfgDIKylvXJaidNOP8dsJ6H4MR7eDy/E1lKwnI73oieaLoM425xcX5DwTY
ovY+Rwgc1hPz/X5tmy0utdGErxAFsW9QQb1qU9vF1g1tMleaoHQqbxnXJj39HqTf
Dp/QJMAGyFaxkMkmuiFy6QXwkOm3WtwP4Z2E6Iwqw45FpPlJ403VBAA2AjFAwMVT
dbQmTHVZiXTrgKfkfnxhjQl514F4D1JHYIIaEcJrmlH0FTl0bA6gLn2YMCoEAdCX
/B4hD/RZK+sQKFLxNykHCNpNF/fDNwmYHouDuZtxpNvntYzFf8BD8MWkdfS5jkr2
cQPx+a/oJ9/ymqruY0zF02gHDfzvFyTdKDET4azRo5ypAU3zYtPMAqAG8CFrzsSY
eLfy3t6dodb/8S85ixzkX97EVWq14KwjOtfOCs2j78wnyUzK37XPZB06KLmNWpVq
StjB5tDQmoBnRLQA3z14cYS95Nt0sisONhG9ZGNBqqPT2OlhWaZnz7vGklN0KalZ
Ro6EkS9eZv39rspQC2ZDLDcoi6FvTEgnK5FQLAHzi2Z7BeHxa6WdpOfpq6VHL1/8
17esl3nU6rQi2lsj+9bmBEukrrnxHJ5v3kMVq0eH/BFX8ZMpvBF9pDtzX/tEJMRG
SkwcVLJ3rloj6dL+jMACJELP7R+o4Z09UNUbtdtkqkAPAqCRRv3HW0LSSqwjL8Xt
bP4uep844ncGSq/b0m5jb8QK0ktIq/K38xB1v4ySl0u1jAwx+nhrzfzJoxgMfRPp
YdMGV8IXN+2eBBGk+BH62WkSZfbqC3nELPEM8UZexvUk46SjwtU/2pIGosg+Yjr1
UacLJKmeIYaiPveCueK7sVoyQCPftlopevIe7QKVCag254E8+fiu6QFwlgzK4haa
4FQoHOb8TOez5IxHffm2NISpWPVHDK4J0E/eY8Inc+82VWNEwCw9Nhog5M4HRHN5
IaVuLgelJ6ufGeEU+Ikw1dNHsDf4Risdbt34pIvNQCZfcEmceqz3hRlgubk4aT9L
WjuBnbe1nSJPG3rtdo4QX3/u/F6TWp/tGXMlzb8WI9mzTqFYK86QwzjcXKAfEQ9T
drXM4emuh2fEACV350nd4di26Y4MMyxY42/ungg4gqXk4t1KfiuFely7BzbrqN2N
E1EOI/p+tZv+Ld9z1ZmCHzKxlY+PMP61kngw6Qp86ZDu655p0Oaf39cDr0+gldez
wG0lb/AvJRyTv0vrPc1w24KaUnB2nbvn3Lj5LkioA3mesHsO7K8iSSCfpguyni37
uUQK1J4EHL72J3yPs5quLLvaZp54+xpj7Gty/qtzFuIug8D77I74EHj/uAfyg7hF
SN58OIJHcoRi9TaU6vm1K4wAXqsP7ulmfDaZ3p1AqwmaJ4pjGPQfQy95yJUf052C
xfCAKCPqd6+p8K+xWCRBJlqawpMXxqRgNX6qFT4LGp34KYJ4IGpn1TwtlGqk/BOV
OLL9Ifq4BhsXEYxq2u0OG8Rs3ftP4MgFhRKBU0RQ4lw1Rr7HyhWqkt2qf0gpMg1R
mXK9De4Ht0okSZMIQN5yofHw+vCJA4FPBQGIKA9HG6BmosJcNo/T+cmDcStzSWee
//6Xt3uLI/70wUsS1tA1CJAK++3mHYGpc+bURJ6poXzVU10V15IEPjpuiJpDqDCV
njPU1sguXfWPgw6e57ccNvpfVL2pFPxSSTEiPAZ8jGjGE3RwqKEuAE9DXH+B6VW/
Fj6PyW/DAkboR8NOFEhKdh4M0A/2QxKOyv+o2OqyTG8mUZ7MQrnpa4RkMvMtnYpb
nAzaj6o6vI2GSswYy/putR2PaAaf9Xbq1MUYHLbC3OR+0twSKsyNRnDG0hv3ILnY
KvVgkdbiiZ3AqN4lxbhKdxqlqWsl5F9ad4fueTcHIp8LQzfHx3XiGBQTQV37S1y4
0i+4V8am2/qdnsdHQMO8IXYVQMZi7/Ucxp+dcL26OGqocvzkoUdgBMIYwxy1KWAf
ZvBfKhGytIRwX1N5vocriSr1bLqDsETaFqVICh/Ei+8URYuOlWz0iBO+AqxNO8bu
IQ1S6jT7oufJ8PcLMk7eaFgRsGJBakeby7lktwQJ4Gllhq9TQy+srhAapeLX8x8J
80zEVVa4ur3Fg4OkUGF+b3fy9hH3vT1FmIR6COPweJkwNhLE4ahftm28Cw9lJ1G1
AfitOMXZ+EyvgKP2Ju0A/PGA9cT0QcGuVTJDlhEKnqe8g+cVmuYEPtEykMFSqSwq
8OPKEBv9s78QJObIFUAY1U6StgR+T8xIkf8jwGvkbw2uJhWn1Pg4Hb7rGPJHJEud
qYeRWqXfe7QXpe9rLljc3stPvHIfEFH6biJzA2YrfkuWE0GLTNWZ1FS1GfJAO/Ym
Gf6s2R0X+nE7m+sBOpZ2/d3EXmlOBziIdOrvMmxyofaiYTtoJxmQ0vSb91QEo6lF
LSiz0lnPL9QKiIRfoT36FL9Mr0pWlGS2ECw2K8qfWaC6tEjJ0JUP0pPneOIjxXbr
faAe885NA1tJ+nNLs2f4gbsmq2hVbsmxPh4I78d3UzzHsqkgj6Djym4rk0JYYIoz
KQhzf/poto5bjWNhlY8/FIqldc3orVLP8GpOywppBA4FWFTsnHbC3YIUN0F4wI8p
ERRa/KyyRmhlvq53m1QOHojl00LwLypYwZLB7IB6GuwbOoDQ8kpdaVq1mkGKpBB+
wuVUVe3lmaohPll4ouqa/S0g89Oo1qYvRfUKFeanAC++qynUnHo+NiW8OEOgbtKi
JmJKifqB83pQaiqAW98tpSC03+aiuOBtVUq6a/IOsQxej3bvUsUj47pJlO6zH7AO
1vwBJVpvxREUiTr7TjlS1jKGe84Qwdku7SEbP7eFtvQuV66JlMQty8Ju5L2RVvF1
7fqQy0A3NBwPy5c9X868LJ6+/4Rw1EYQ63Msj1Pqnt4J2LetSd4SOIfJPHJDJSr0
a1vfD6j4PxWx7fAFeb+ty4WpMF5pxx33tT0lAMVXxP2HwzV5SONu2tnGCXgkxN+Q
KXaeK2/5UU9fRzVAiId0cWvPDL5mUYN9GQOJjow/x5jFQtfUQDYnfCiLAexc/3o6
NA/viNX1jpx9aVkjSRz5Pz4WuyhWt9bP/3HtQokcpbFjhbNsKML4uMCFPB7KUBC6
5h1gac5Ah9JZGogqr57kW0YjsiksR7gFjoaRFSn1Z8J/DMIb9WWIpQN4PWWPKt/x
RqbYcXq7mbxMw6xWAL9bvim6s4XBrb35NUL5c8zBBgYlxBeHcepyoubzqsiUxr9d
CzPGRr257I8GnCagN3wLiAQOCNoCwQeQ2uWwqk0FxY2rrKbxVYe6yAOm0oVbMeud
5lSNPDK+m6R0VcRuYGIPK6dIYdcvV7Mj3wKiQcpwk4uZoVGNXtMFlV0/rjxigKqh
SmZgVDokZRJ3j+8FTMdFHECNIPdQXFDTM2lweg/pfREV4ZT15lVGsfMm4w0YFuNX
IVa/SFWugnspLk5+a5oz/D+exqxMk9N5gwypYH42DGrKZ0n4DkF1oF8VN4MZFesL
8oPQWX3Iikr50mc+T8ZX4G/IluBg6IxiZLLNeCVgcf085HfFrCROEjQwztJhg2tU
zNWRdXCCORVi7Hnrp5RLET7XDWkofav1GRce/5NbMJVAhCP+WaggC2+vzk2JNJ+1
4Eg4xmDBZsj1n4RbOxvehMaGfmTAH9BAKtpNMhbaoSUREgOv2+DlW9YBIGpEg/fJ
ngn9Y7UvWBTehzsSokDWzp0oK050tkMn/FeSAiStO4iiaa38K5KnFrGD3MKXgOQd
XJQ0mfAO7reMY1zX4n70ByLT1CkcrbmFFXXF1uUmBo7Z6deY4Vl+txzYBr6o7B8W
TS5LF5DcCggMvVvGfyS7LWKSj0+mxGrafMDSe47OQPJSdnxMRIR883r4QBrzxZFg
Fpiv78nct0pZ3xgvsgpfWrjvEIri5CsyH1Iy+Zq7BeTKGpOZmAF0CN2kIoQQYMsT
uwWqwWglvSlsTaR+8tC3snX1idQA4C+Vlkg9MhYERcWLqlGOMjuJtIGCv+8pe/bE
Gi/oWYWmkHvYHUQiJPBN689uWGjqcm7n7QJPh6guuH7IguY4CdgulQh86rd14q7/
U5bI6KtOBUMpXUYXF1tktHrNS0geehJuYQ5/doQY4aNHLnv+Knbc4pwfsoPfjdYL
yC2ADacEdCxSIaf5GtKCvuDWQkOTUxHwsMZvcNlFy+Mkh2GrYhFgobPzjtjryL7q
6YF/ltTJ6vwTrE2z3mk/uqEiULyrfxb7fvQfiXKiQFBOVVZipRgMfEVJxCWhjkP0
EL2UCilf/jjQQfjWmCi2TXNI8R2QBt9z82h/xFQXc0mo6lSfEQeNHqyaBKRaBwM9
B4/4BoTlUXvTrdo87vjT4gAfNAHaQhsIkjkriTaSDT4czDxktEdSkoE6xWTQh8JW
6Kt2v8qxAu9QgjfNeAdt2SNaaFGuW6OfqGlKq3raA0heCCUsJldd9UyKkpJU08is
E21Uh4Rotc2R7wRRb8g1GBM+0Ny+WTc1Y3ZmowQRGHY1nINT1knF9GhLDFTfA/Wp
nEZOcUjg2tuABVGH2XfUIqOOgZT7lFuMXjv9GeeFqUXAiz+ew2C63TR5SUVPpPlk
uZyHKAlHrqCHcsvDkxYNM8ManRoPknztONpORu/bcHwhw5iI8BZbVt2rdkagqhPc
GMYRfFMedk33jyCW3gqVDsdMwBdgnyDb3i6SGRcjr4rKJWEQtcsULz+gUp1CWjwE
cRTmeDNpXjQFa5j69FZ97mwRgtrChO4yCmEsgUMHGnjlnMxxzDsBy+zXEAcbloTE
FP744I+rYutcooNVKGAVpTT2nQgi603QOyWXlxIDmBOlzjPYR2iDdZIyZ9Vg8HWR
AfOh4uDCkbwFtaRbEtmSssIuHa9DYwG9kZysdCPud/RAlmpr4zf8BPCGzUGPxiaV
OGg0ifMtdc16J7EGSfzpKJTDa6g0o33rNQBF0PiDqBdDAR2m0JUKJtWyCBFUF22q
CzRjWog+DZVwRJ5h9g83U4pGhb5Nts/yprIGgMbfDmjuzY5vGYky+ijj7prB+QrH
T1DusTpf4rKqZNw7E9ZvN57EXoB+J9+O4ya/+OPtz1sjqlCklHPD5ZWJd4QcjLRw
W9XBB2cyUBthHiqjiq276LbtUG8jzIQP2GFg5YWqEYKa4Of8c6ePdLJ31oRz7HnI
MAqUc9eJU4JqSdNQlm/eG28hX7lIIoATXzj4+HjuT2w7a+UZLJBmiani9Rq6Kom+
eMB0gieQWaa3B4Rc5/wUZL5T7lym3fAhNp2GjcYKAq8W6TicRd7ggfDp/nu+EAsS
tj84yQ93xXt6JaSWh25/ddYlnIrXx0k91uT8CRZhie15QvJwzL5uHpSTjQiAinne
VbRpb63OLPiKU3oXyglKdmpLzVkdJuLa9CzGcYufiXihraNnIoqmj1CYv/KOmBg3
9OnN7uwD+M/5S0aXGkefnNsA/gnoT1mOAUNQTcZ+d+rIp/WbvX17PvDE6X4+NkFr
RUvPocGnFdmbQo5kvR7al2d4goYgM8YqHaNGHMx6SOYduG+005qeFRxdwynKocnM
qInVEAWoHjyGdxX19grZO/vjRP2suTIo9owkaSFNu7i6tLZawX/U7CiJirpHnw4T
T8tK/G+W4pwBmYUAnffHvHSv0o4Zt4IjP8hsFm2oRhh5uY+hmbagkhqYq6FNS1vY
nJAELfNrCFqyG3qjAbDHfgx0yZohWXIjY6Ej+RhEv47QKRNjERz4D2iIcw31j/QX
jZ31ox3Ix98VkQttXlckSiETZYlyAzDmslzKMM+l0wyPomjKD9aEc6y/MY01Z3QX
XQFQxv98LFMOEayVUIVoi/DfzA8avfoeMuk0kqcWfJj7Pa5ocZj33LVnn7Aez5ev
sjORaEkqp/DpvMYIU7U3BIGYwmsA/Y+lgur8V/IyVmDFZ2vJn+PdVuFumc6uPVOq
W9MjE5SDYdVXlO1M+kHSU0829gDSYiATtmJye5tBkKt30NdTaKbEEahKem5QcH2j
K8GdGXHIU8XO27ILAtUCEd6ouQjKkEXN6tZhGrg4Stay4Uvu04X0aCsKGcyVJR2t
osWn2WUqiENeAblqflD2p6YfAcmNsqLOwASUWqG01/kKwM2d7lI+114wY0ONPg2F
VBK1WeuPkwaXgvtIh5ykBvIu7aJHQXI4E1wbcwd4teTdpiTMZaDgWHVjSQuziPeX
b6n4IRi76j79ROXcjJYPH24SzJH5QI1cl//Ws8cjNCHwXZ3/WAtWW3Bers+35vH+
wMSkJgG3trFnctALH2Yabd6j9ZV3kDh7UN/xFlBjsp+j0zRcHgtAVB8siRLE57KX
pnOu8D1RKMvpcWvHmY5L5+H5xnRiiBC+RryRcuNGdBgZWK2AEY8kGjmBxvrDEQRL
89fX/Tcbb3L90qFgYTAlfdz9yX8+xJW8zFZ1mtfqJvTor5BCXJ58RIJbUJexBFo/
PTp6NRMpelu5+KasfgYZBGHAQD8QolxV4Z9uneAlHgVfcdDeINGnWTAi48m2Inh5
Dnr1IrKBwou/qnRQQqCxPFDeTahs1hquTSBehOtI3bn8iuJGBFovldtSTxc1B39m
G+eo6rb4Xt7gPAwm4snAH+4HAOsDyiPj4XFbYp8EbHs9V79bC6Ni0uBvgVhqjRg/
pYyrKLGEzFM7pbtfi2i4t5jDl0LaH0q9BCABE8m/m9NhCggE+fDlyp2e3RFIH6sr
n44UTGX8SXBjZCJS6OBWcq3gHkoBHB1LFjVtypv38a5Kr0YYcLHB2ENxgEaKcLOx
BpL5HN38HQ1Xwf5Qgk/+jp5t9Q/IClqN+RH6KsKfQnMbq5rfqf4hRPmShroRqxFn
B9PMbdiWo36/4vXqTXMwp0gZF0gqKgG0vVwyS4oDCMDHYdGUi7d/Ztj/OBkJFH3K
9nj1QJIhxKyEVGjJnsFyKt3q37dIsD6xUuhMZrnbf5zZusTb0k00JpmRCwSzJC7g
mWGrAuFo0BVJ0843/sTwEJXRsyzFx/5EQl6zs/pl91fkq+rdkpjsm6RmmAji3ciL
wGRDgfcQ/2PZTe7cYnU6YKNmxnriX/7Pc+WvMl/exoKqGtyh3PDZa5HryEYJMcmw
iHFv79WehFMUBQcOExUY/V/B7CbfyhnLsYAaLOKF7/PZJu7kg9mdqU7vJkPo9UID
DuRilvSfWbMlEhXTY2zpUds8/sXQZM6XrdMI04ai+Qst8QfebNfszjnJ58GxqrbZ
nh25xfDuCiV/qn/msYHrVvvNhn2PEHyyuw2n9GnIowyfb7c1GE0naPq1P6McsnbA
Flgsaw564UYurC4JfovjQdZwt9m1OuvLEu2wvqEfOT8Hh8XE+OdY0u0HTxs0zCnS
eihZSCgIad+aWQ449nZNJDTY2s8haC7Kap0EON3VSO0fMN0Kw4dUkDoKX9roWwkj
uBWaGDXqi1cZa2/zRxyPoCEPi57LKOh4ZiDSV4jCBRdpifQhYodt64sWqlHzYIVI
vS+bN7pGV2YBJVSKTuShy0oBei7Q3+ClRfXLeH3oNj7Zmr5SeNaKuu/HZolA+U4J
KeJLxJDpqsB/yGuF7jPsknF8kEDYueElgLkm0JCpi+9zyswycuy7ERGWR4KATF68
k0Nd2Y5VvQeWk1IkARh811GDEmU9NnmPGDOChG/jd1zYG0SX7v7zWYJ9JzGh+SX5
stTCFFp4Q89gFgItpsAe9DXIupLg40RUS4C5VBYPnz4Bbu7DIF6Y4yQXcuhbmatE
dZcf2LPzPyYCk5qdvKUnX3TYyfAnzprfdt9UV8jrGw21azFN1+p3TkCj8tjNlEzh
ov1biC2oaPsEjISAbmBxD1wlpgWK1DmNlL/vWA4C6YiKgYMISV7454slXrc98V9u
P3nG9gUJx7fqig3k4mp2nuyt5a2/Sg8ijQVNZqtZDqgOPfYTXk0sDa3uPZsPOq5G
EDwx3yaNEhEXmavaAUdYWggHuhN7iQ+Q9DOgba2XHfugPKWz4OGZFrlmNqyLJIxt
YJMLaehl7xbH8+YGKxE6gnjbqeBnZaDvvgImSFVfN8RZMEh5Fqmbl4QrVWZIzv9I
Rz1Zqnx8LB1NiBLol1HFqjWGjV+X+K+Cntei/yL6zvjGZkEriTWELjYv8T6pfIpa
5RRumARbtcTNdCXYoO9h4AuQrcwWAHLdsouNBs/DcggFDs5ntQcGwuMsgvaXZ0AH
mFjsYLYTekPLReCvAOricceqILi7xSm06WdElk/TuGXLGFAfFc7v25W6HZ7mEL14
HhG3qjk52sgmQwW0zImxdBdgs7bVEEQ1bupATursmVaV+N5fSpoVD5vOz8qkcGoT
ZnXucsSPFHKc4bwKAaMnv3NWUAOnC2Dby4QAXewJijzRdH9o/n5mQDS7ZoYZhBIE
ZWY8MKIMCBrqJUKM7EPjayIT1WC7PxdLL5N03uDUgi2nUzxF5wQQG+ZUmjeAGkBd
OqUW6h7qLc+ISWazDUuDHSJa7AJaLpKGaiwa8VmbT3sbhikLHEBxM0nnGrg3LSTq
3ph7VG6UIqjvzr6RWlBy/VPJkWP7/Z1eUsFQ2QhcBi8AGuYYagHscDNLo5q2jg5A
IkgBCdQVV12ehJAmFQ79UQUcNwlpv0R7xpPTeJ8FBC9Ztd1I9vvjYictBcCRqW2p
LT3zCPP3pjGLPqL1QHs7a7jtmCdtKkjerSnsLMcc7hZb88j/clK++9TGfKksB9BB
XgLxJQyWqOVYxzqYRCXxd1UCrycc6xFrHOjvlAuaKZYLJrY27h0TqQTkgvZ39iV4
mPC3c8nJM4+bvjHwd7tIyG0cEPv19aXjADX6HjTc/qt5vngEOuLNDOjN4Tf5QpTT
Bxk6Zk40lJeN58t6KdpsWE4cPs5gEYdwzhh9yU/6hYYuErPSfajFtZcotf3qXJms
ROldOrXEuYbfUAgIL074PaK7yNxrcCEKPKHwcd9bFTvI84u0jfOwhwJbmYtR/3Fg
t0H1Ch1P7RIB9G4amBzJpP/6b/nkFhyRmceLhVlNn2awBB3mOdgAqmrLJ8s5KDJT
269NOq5xmfcs4gDwJ1UN76vTPKVY+O7X7N+NzlKBss/0WdYSUiKqbkE9RNRPsJAy
Q4isMIy5aM/WZjoJX6Jzk5BOLrJ3tgCWk2jWBpZDzu4X9XnAGLyWumFCnkoYFtHS
iN8XgBWtdoZit+lG/CpBoJY0Mdalv/miogC6fY+y5aWPvSrCXqtSAiVbzwEzzdcl
`protect END_PROTECTED
