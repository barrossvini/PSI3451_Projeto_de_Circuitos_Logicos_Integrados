`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9eSHDa+1R5MUKphsTe5iG9JJ77WNJ8smmhFm2QrwGX6lPd3v2xK+fqGVWVT93gG
3X62XT+3WY7DtqQ1rF9c0/ungl86otEQB+Xc8ZW9aQsWxMvBLSrPzFs4SwPrLXlc
yVZRJ+68cpgley3fwTD4BHNkTZbJo/96Cw4Z8dYIVZUiBDgg9crL4UDvYph5UxE9
rYGTYCX38O2YoS285mOvRsl+oPNRhFdi8rAD2OBw4mOk0IWt/xCe5vOZj3Xs1q6O
4R6gimjiF49J3ps2XQDbikmH5mHEBV5YoSBXYyYhV9f2LPoas6QyOU7SRLAcBE0t
v81GPezKK50rGy7Za9rRq/ZLr+QtWKLF7urR3lfCkDdOuGeLIGpuJc2Y5Zs88TwR
bh58YO6Tah8GazC5eOyDBvEAjXXWDx/DgG7VDy/gzzF5F9MAH8HTdlAO6kIU3N0I
M+3C5dS5Pz7nb7/jIDyX2lihY1vyKCoBEF3SaR8lw0VNc6CXwcOIAggbgpkTPZnG
4LjNIbn2MP0Cb1j/gETwK1L+Zye46o8/u1GVutZn5N49/7GRxE469puhjnMfvd3V
J+qpH8SrPczcFk8bikdPvRpOu0pvTYSSrbA/s8mKK1JmaeRUNQLw8IGKqGU7GPxY
X52nzAnAtAiusXQSUnANRXKdHTzS+QbSl4uFGd8yj3HTyEP/lhXTFHKgZsFM5+Gq
EsToIEj+vjPIf/YZoZuptwivrt/S0unE04aDZdpKvdKyHrooFqCMT7OdmkBNvjuu
HXPL8wm2e4+Vzh/ndkPw0qRLMmkSDE8tPZyAFq3d9ZQv2C82kE/x47rXne4qbJFf
yweSHlh2COKqq3JwYD7vYg==
`protect END_PROTECTED
