`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hIs0eZA0cUwe6No1/EKW1/LDb3k7yjc6MMhtan09cj62hOSNWSFL7SkB5/t2arjH
uG1czDINY7Qz1Ep02XT3iiaSKuwG75brFrngG0siAv4M3dhhqXNF00EgM9jOXf5A
OSrr5PU6As/jFbrU+NfR22UwklkkNzCJEm9gFiRsMK6/UboBxElPhme9I71vKtWW
hTdlN4Pthi+BaMspAJZBJedfwl2KSMZVKyjK2rdj7B6UnBwP6iTfGoJd12uy77uW
miZBRx/bUdbitciUriunoOG5IMzRIYzc10otg6iAqB/gCFZcL6ljhMExmy/m6JW1
Q18QdjyBRJAm4xn8gL3MmmwlIG0gDrriGlpd2emgCI/tKPMDgvFlVQxvrFPDtBAe
gblzq2az2X7pQtyRcrHi2Tk0NhKCN2Qtxq56oi/5JR/Z2EzYl0ATzetl1H2UqUwW
EnfH/r0cwsCF4rhfKfSghBh2icvvFV8xGM4+YXIzGEl/vFj+7kl1xwPnS4ykqJKE
PBxIwNMOSGtNuwzKX6Zr5ecM7v8ApWhPg/HRIXaW9LybsgsCZtZlwq+ZiQWQ2Hq2
OmuFO7J7fgi1XoMDCpe/cFVMP9+rG5hElCMHgW3GlwzwcjqGJ9+5k1iUBbVrRlIT
UnzYwF0mj/3kbl/ZW6qQG5l2Ed+cl0OfPD6Sl1GPQJyRQsBvHZmIbcuyxPFKiwlt
tveFv0GtO7daHA5ap+VBSzl/eLL0RpVE5EzXZ0+p/EObuawnl53cbjbFDh41kK8k
CZ2RS0aMa61RcKppS6SRKiRLjm1vbY013R7upV/WOgdWhlHdBcESsbxl+XqHQZOV
KhrLEt9Z+iyrMN8NoEapTg==
`protect END_PROTECTED
