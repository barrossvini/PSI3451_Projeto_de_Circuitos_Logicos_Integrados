`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1a9mVg2+0Cw6c7+7Y16a729dfMFdyIfare2pPNYRPmxEcp8pQcUABcEbSrSjh82
KHKaSSwSuF/0D/NgtO6ztY7fxSY0SSBOEUDEE6weTBgxs62Tr3O4bT5yOqf3ZGpu
xhjBBy0niw+725oW6legECsNqlMMFPl90Jy725ctztqbe3g6tdq8SBOUGPFS2qcQ
4gP20qo2b+GX+vlo4F+VsFhe31Dh17CjlvnMASdlYOO+Yf2gfoj8BnFFjGvYvxFw
FSjg0QNZ3sImSVnejtax8Rd2+KJObaa9H29VYHpg1ckGzzhtEja4vRLuo8Vie4Rd
qSq8RdzydrkAD1oiIR5J9f/5m7+shqe1F1iuHx/RZ9CFiT/2dchuYxS+SYuc4UP1
SyNgB4sJCnoDfK0QfE7H+Efh5eyic3Aij1fi7K4/vNqRv7Ge52nZze/H2QtVNbER
n9AgTv8y6TIKe6Yb4vd3PfGidAHoQGcSttRRvuXCmaAghKNy/f1au4bxVQTCokW/
13gtp2KtiXRdpBMjz/d33EIU250AjSvlFBqqOqcRuZz5g9n9k0i/faphIstd4u61
v+RnnzzDMilAUEvhkH4+Jg8SqvNuXrC+eB9gzN1gGT6zlayLtOxlhd5wtaH3CbPY
yHXDYtdA01rth+/GuCt517qi8OInao4J5/bmO/onKDv/keUlbHMRy3UF0sYZCJSs
q5NeZB0SZD3NMzv8a63rtav7xK//DCiaW9G2cAjdbvApZMiZNnhlVVxGtvTAFEJf
/BGlctkkP6D9yK+bEw8RbDMfnPNvBhSiCvi21qleWmOfYqVkyU73xSzYdL3D94ZE
rYWF5iqHlnwLz+Em2sgtJ2sFdhrLx9G1Hig1111R+Z+Uwd2kdBHRzZvTf6Fpxa8I
nBo1TzTmLqMJq5gkDkeQYFOKSAFBCPPMzF5cXClS5bQtUSDhpl7o2/urKorE9Oo2
fKxbwQYF2wpuG6e/duXjUYUzkdBT/NG4tFd5pYgwajXi2iAN4X7TtO2aYxcboK5d
PX1Ygh0qGlGqc43vyqanZOc1WG1+Ze9ZXm4WInA+fLBCAB62cnLNTrdMwJnBCoqq
18XW7G6Sm4WpPfWx/OUfuNM1CIA/a9Edqx8p2O9RKgyNQKyx4Mwk0iPc1M+x1DLi
hdn+blwJ+IRxt25l13+tMRkjo3/yKTA12UX9BRXWy5yYz+8dOR+0VijX5s/fUPSp
5IJeiSIaNA0G89fop46mw2yUPbkTvNG9qNs0zmUAM+tRx3mZbtnZanYphSxP8Tiy
MuI1gej/Kyit5J8JIFS4FfuJebIIwp8WMCTnD+ep2uyJdpvkJ0eKsqULOEt5fOhN
8IeiOiCbM0VFFs2DVNiWXePiE6mTslCXv/yWJgZ35dNG0FP76sLXoM4a8oWPSSqQ
2B89YDlHOma9bvGPEjbaY3RBGGLw076U5u6hbcxKTPzJRIxiCbw+DXpuLaCUHcGZ
uq2LQA3rbyb3Sqazmgk9Xic+nOUfi+byxUpN5mBYECZvZt+V0CBZ3f/2jVS1QcVG
wb9l+pywkFCP7CV+kSjeZUs+rtVpcckRYq4AVLUHauRoWaIG7xf22a66qEIeZOgO
DiAP+Hi01AFj+brdV3wnSAXjMFpwDJWTwqtc5gnx0rLwW9opEkfjFmjtku3aEHic
AUhsFgMF/0ac+lcGHbN6CCSgO8dYWQmw/k7wJSnAzd8PvXQVIGdpDaeOHekeczc6
xYyFbxvE9MLX7ulknPvQWCw1vSNUDcAq8NT5lftb3VUYCnSTWSoxtKchnkpL+MDw
OUPJBfklE9Yhx31Ytz0ObRwgxTW0JkXsLvXSzNa8Cp6LFZahihke7z/Ad6tCkwOq
ANjjVb6Njm24FB7wGPwelJoDjQAM+hk0lWlpEs7y4E1r/wyLyvnfqvkZ+BHApVZT
Utoo2bNF5JZbWF+O+bSXEpPpL1u2Uk2rXgtbeI6FLJsvmDZCq+FnGvaxnPPEdXk9
V4+wVSVY/AhQrlS+Ds7ji2p0+TW4HnEGQZRLpsL9EO2pTzR9yALga0BwnHHBITHe
BtzlWc8IkI2AiYsitekhcywdcgECEgH6FSjz7GHnK0rJAVv2z1B1Xwf3wg6WjYCs
bqg9H/VgAFrd5I+mprS3nWepVCl3VT6nljGYATiHzQT6XYKFM9t0kD5gnipLUnHe
CLYcIHvCSPntcA8YjQ/H26bDRqaCoDMRmUeVwHPfjYrmkGXLHb/XRXr6GFCcKKqn
I/M6pHFBqK8p/tNatrPJuU6We0trWzJ5upQwe6RuMnhc2MybK7HiVYHJbHakMSd1
Sk8P9ZdSqpP1Q/D8ppnrd0gP5L2iBvOeBjY/NcU+AMQys6RTDR34FRexQo3sjkeQ
j7JlHVZTYdoZzWxEla8gmpL1RC15x8I5C4DlJ9HaCMskxquiDOO7dWUgeQWnaX4+
K+QAnevQ1U3o4SHPEvZEYvX5vokTcwSpp7ex9eL3iB6oI9DIjp/vkTtA9LVFx9Z1
ZFBoOt2ghBdlKk+s+ZpHlkbqQcZzYAR6vqCXT2d3eQF4Us3kRUuJYl1cmNUPv+vK
X96EQyhTRi8UIA1QY0GzDkWYDwEiTJIh9F2NLJRcnKU5puSL8xiaNBEBBZniKrim
6t+sDMqghBrQIWEB95aOrb32giYyqA03bf6883NVn/esAmsA7GbIo7PS2e9Jh+PW
4R5WMBZ2Wx4PIi72pMueK70hJ3anKDQzmASDsc2v27a1ws8rn7tRiue4xf4QPb6K
cHcw8LrQJrt0g5SIdPTBV3TPLamUuRjxMfBm7Gqx2Wvmazdh6okZBZ7JsUiys3rl
D0+ZqSlqpVm5YIV1SN+dfSB6GruDmDqofh5BFuE6ZiuebGzRnaL9CfO6Q9bNT8PP
W4qsP0+1K8xulU8xMyYgMyyBMHHu0Li6o6xJokbIcOI6FCUIgdwhlXkKVswuMpDQ
H/2nUftaWDijKwPXMdXS3LgsyYFrO/1HHlAp2p4bYN4dCgIVecpXbFYMDGCYPSOb
5rGqIUkHLteNokR08kut6oPTx4NW3I/Z02o9XJY3TfP2M3eUaiWBRXGfLg1hOxP7
QM/Xq5LNYWg4RZl7qZhMWpGULlVFxgWOlbPJt2OcEaqMy2oIW6lDlBpyVXIKSebL
zfgBk7ejTxbeOatnaPCzZNx7XpA4AYXIYRiLaa1L1zC6Ky9LoUUYwGzQOTUf6C19
Dbv37r3kQ64XQJMFltI6BLFK3IeRBI8tVDY2ezQyuh2xueNO3FjRV9AhJqgL+zNi
e3ps6SNNFIPWqv29MMPwUQ23pHX0kgmlr1JdjRInE80R1QhCGc3xCjMKNZIq4rPP
ocHZhxGXIEeRTHr3QA5dEZju1pKAbSYBUPwrt+qVaaszCdGb/35cBYNNtSWR6GBn
H6okRgc/ohtlCdWwxd9TbKmVBbHURAXMpNmDLrB6LhuIQmYJTOt8kv+12dKbr629
aiJvOWeGeGvgDks42ErSg7rhdta4DsiHBtQEd1dlipG+9HJiWZ9HJVcpc2wIJNWk
WP712Sz6u++bHFNPm5UtibuQEnojA494cWWpPx0H4oJ2eokXgyTRaQwUtEY1n7Xn
Za2mMZP/vDHZUUwU1+i4Dj8dZY3QQmfMsIX0O9v5d+OIHvYH5scv/HqCN3Xk43Th
+IFBeLvtVKqHx/vMPSrEDRkrHaG+qBsg9NymNJiThHpWTQ5TMrXkASkfj7BZ1WW3
APF2jxB1CcXA64THSndwHs5EZ8JB0bmrn+IH0Eu/kPv5Uy3hk12RMvrOv0h3rKx0
u27R0jDxADkO3/KzBB8jI24yETPIwFD2cNsOrC1mLttjTGLVmOXYF4mg4T2FGe2s
mFo4PMV3xNU6fpgbaLX9rJa3nXGuRK6n7fPbQx2c5guUYS2P4xl/G1gUic3tEMu+
1r2O86zEWX04NWZLPIysYKExUAQEWLlPXd0MBe0Mdw0kPqyHQ5RFwnVvxkJfU99I
I3N7yWKdI7uAsfj83dJJPvDPl+C+/Dvh/q0j1aIaFFIrFkPuiThucSp9JiJ6JGTz
xZxvYH1sE2FpLxmKzGJs5xtnOXrdT6T3mU1qZzJ7+WEk9vUoSxe6UCJeE7DMfHBX
QjnwHcm1T5isH9r7q8V2f9Z6LIGVKes2ucLhPsyBWPKDNS/OQpTyxbfffMf0bIpW
xg/yPGH+44MRdePyxBCy7JxdJmRw0KciM7vKLhMWT0NDU0BUr8F2734zLVX9fYJV
rqF+ImwCO6gSgGxa7WA1XEteHkFMtryhl1gtCjLYvdp1fOCWMqH/Gvx0fi5Lj/dA
2Kk/dz7egKM+65+eNB9pKhEYUTVhQjUnB7Wuy9VdqlQhqvBNdWdD5vCaJper624p
frxv8xRwXCsXMw3KgJ2vjuezSQdJ5LzWibTa8tOvmqpYk4zK7vlqvi8pYOkqorti
SUnHhQsvvfTlDu/c+fxTAfrBt0E25uQWj3Fis9Jp6JnMIu2EB4cwuc+5MbBFrSaz
YjyB67bMs9Fd03BjkTIAhXFG2AdM8+1ZnVBpUdZQ6gp/Lj4xlpHFDbj0yJsceKes
cBDi8z+bYpwKaBGc2WGsYhnxYXA8OrQwYoj472yv9dRZWE7jM3vJC586tS+cXbCV
OIXVeqRDp0h721PRhr9LXoDmrKb6pWvgoHbaG7UaVFYP7gyAZ4/SOiOv8ztoI7hS
cjxk4xzj9odR2OmjCxTJ3zyxF0diGmtJJI4XjwQZ54RedlG4GzH0z49hscSxCA6B
FAd/vng2y8k8kVHVXM9Mhfefa6RcbvxYMsBHNwmsJJjDg+Tln/CAjDo0Q/AKXJhe
WDOQCYaA8c4vp+Yf7kGFBRuOLpG/knY9Yywkj3Cx0oYEEH9I2EwhoA7xr8069dzk
mDHcqru/S+XIwADDw5YjmesvQv79ktDAi13jZhslJE0byBKFcYeddMLVXqGfSiBs
c9HNH/4iu6HblPiaZFReIImWuNhk66uSVwQQRYYGyvDIICz+vmagI7NLzHtZxvGx
qj1jkKzNT4w+IKwu6NRp2Sodh647dqkdkOnOq3BOCjCKNqM/5j348hTlAa4a1Hek
7dDZycLj5tzy5CyEAS//r+H2euqJx8SvizEplRTDjqDzCd4zatElUyIeIZCQ2PtH
yugwHSEvXWsh42PWXKwFnbsRa0NMOtGyy5KYt07XdSk2TD0zXUsBfdPK/xZcfmp3
EbXCDct6jOmmTb+7bhSGuSEjgwOWwTJFaFcRFoyt086v2tLie95XzE6nWlcYq+lz
MStNrdlT7yHQrU1esd3Qs6zCAUDaV1p0qmhkL7uqBShnf+5zYJbnGIPW82pLQ+oL
bdLu5Egd5c2Y9McgECViOKJ9nJ9WQhePEMeREiAjCrulX6Uc1Ju6jxCv0B9C9uGS
25NSXfd8nk5ZsiqnBr8KeJTjKa2URVlR4m/bhS17ohjMFCInXGKfQ8MfazoLo70n
yJ/T9mguOOZl1yNS0z3wnMMAL4GmFnWtLt8XDdG6YqC5ndTtYjEplm0U05Buvayf
JHL4GiDjnISATDOYI4iOQ4QNRyYLFtgSmqC1d7eEjmsQ2gjjgJLa3iwJZAUaJBmc
QqVbJdbQJoqrcXwVK1cT2vFbf5YuTZqoQI5GBhHx574l852Zx9Vmi/FQ766uOGZl
fFGek4G9xErSrjcStfWyQ7KiIVoSsFYYRyvbo8Gff0j2AV8obv59oNL+rmwhJ3Qf
Cb6W29bSw8iZZpl1SOH880DCszmL9inVRWkHqh5KFVSRGccytIB+JVSIduGhj8VF
kppg3/gnLwK5oElaTpmCLdS8YxCka1kV/nmpAdD+a/bO4qAjCPIonTWL7MQh6z+Y
XLa6lqClFVEeaH/rQi2ICWTk5oMUrL6K4Ho3eJ2rJwpZERjKCrWaYxN7ObM7obXy
/9UXRjNhs7tK0sG1+5mejBuypmQ2fQK0LUGCIqO5EBIq8zzkP59QRTJ5Kv+5pill
SKXgaB90WDd+TV0fksWa5+VpCple1Xr+GplmOPg+f0vaGvXqUTFjtmqWSGTNYtU+
ak5FqgamTAGZWwyvoPzLtW13mPlIoSJ7nbufxiTdl8ykSd5/e1eprRKu9rMVvAQy
nwL1BM7zUI1qzAOLx535bmGr42IJOcPrT7X/miyUgqEAurXOXzxVNJsQjlFqn/L8
oUIdND1XV+scrJakfUGvAjh2mDmQRT3Zs0dR/i2Pcq8vfGsyu8FPIWtnGmhL7m/k
l4kPg8r91O4XfgHZoaOhYNFl/3TlbYz3Dd6c1seQoD42m2Uwe5JOZmFY3fYw0tT9
0QEarpaZIAQK9VUxuLMfIob4yQz7cxg+6OqTVXxjceJzJYwQqLwE50g+s48UgBP8
kxqcPfe4WfTTgjB+xYne0EvpUC6/w9QtCyduHWe5L1uvCeCSgulWrGVhRMPKhSd5
KPApHwm/Yt8YCG/buNzjT/KNg9LOTFnO7YH4p/xqJhZ+7LTZ5vCvTqJb4B4YlpSM
FHuktFru5ZNJPPRM53Wm1c/ZPyBv4sfNM4KP5BGiMT8PUTgKZkth2YYjzgtEjreT
XnzgPLQsOkRjKC2kZZlhrKwzBlqQNBnA5/zmSbA0tEakJgRgzE9YgYpvAWgMc2D1
MsxXWm6MzO/thdk4yV8cK1K1uhmhSPAY5cWo/+i+EV1AwpddIDFrW4PJoPECUAsD
D2R0qXOq6jLlnwVAtc8f4NTybLZ1fqpEYuOdcNn3WKq31Tn8CDG594iw2IiKFipA
ciEbdRvdkXf/u7g5VYVADz6Bmsu6cVpfxvdUsmRdKHuNZpLAzFVVBS9UUu8jnoh5
/EYOrpp8Etpvo6STXe6YrZ5o3wdtNa1pXFc58lSztq5Czbda0lZVF1PVt+zCKLOg
`protect END_PROTECTED
