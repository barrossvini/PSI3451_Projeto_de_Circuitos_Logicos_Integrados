`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AKBYsGYls+kgYhwzExZnHR+Ywrsl3Pd140UPirRfjF28dSO33346EEsox1sH51LR
85FO26nm0mzT8i97GrpgZcHka+jlEzUIY+JfiQrxgY7yZVPe/TDhef41mC+b3zc0
3dnx4XMTyN2AK7nWUUTLldJM2mj9MOPrnRd8zW9AMA+l63Rrk+cR3BhSbEAXAB9F
`protect END_PROTECTED
