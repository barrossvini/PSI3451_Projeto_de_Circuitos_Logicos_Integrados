`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fcI8mwSjILYemRhRXTzO37FV3bcmjHd9pY9VhUEDrctRSNpXfxDaE89NSAVNBw0u
uZA1cTUHgvRwxNzMyuBDKjF4pBoaenw+UaoawbeontcA5gRWlwWBYiQfOOpLZPJx
ECa3d5VWNdgNhpW6ocx4486mA6JG7GZ560dYb9KZqEmMo+cMV/Hq4UpnidV59jSY
nBu+wSWTWKsnrg4NM5az5SjDrOTrks8JjDIXTSvEbTXG3EJS8U7YsBHLHnRlS8gz
59ff20ySCMsqK7VcZNSIXftGVwYVEqg+Qire7eJzeWg777sODcH+hYxrNxf4Yulp
1QeVCa3XbCCAuYefR5gp3XCs+xhLyDW0ZD2Itija1UyNmQ1RICE/MkHO6XMdvNs8
wQgoeIfEcu+R4nucSOa+/7lUciDVBB7EgG97ij3lgXHyYMbHjCxwUzpyybbQLI5x
ePmOtAXvAYA9h3mg3of+gbHo0BJLImPQ7iMcbfgIch3TbISy7lV5jHKarQ2p96Fv
bd0qivyS02O8uL6LcCN5lP9qykoPhmS/zjSw5AelFwaTm6ho+3+b7w/PmQM6BnZb
OTdu+Hk+v7jXBRGgpi500yFzd6quyOZ018eAD3NLKZoCXhMwZzRcVrqMct1q+GNM
YWvZyzZDX6oH0co7pxK+UKGAE69iVC+y5lLCaACrIB5ieym4o31fI/Y9Bm7JAErs
TKX4lZs0VHnjRmzSJaj8mxMAWdc4tMmYQcUHRGSRz7buDfRTLnTbSRgg9yUB0d9N
tJ/ZLmZBa9aWDeL1kOfGqwyEXa/+IEd/+CstwMGvhD+mjskel7/CUADrNXE+d06L
vmL06QsmdZlqYzKj2y+Y1qtxFpjGVHXr68Gd16/UCfeiGv7DelyDKghAnqBQL5iL
qQyQFwG5pFR9ssRz9q74vj3R+czrwJmEw6wiDtD3rNoGRqht+teARaEdy5uieTmh
vb3cXDJVMO5Q4Dq4mMYWf5ys20AF2BXXz4bJ2f/EvYKv/s7JE/FUZ7jUr380tJ3L
ZBJ4vNmnAQss8XVSBKKOlnWJynz1T8TH2Z+XJhZkcebOwEK/+ooJgFGPou83KwbP
fKNXCumRPaebNy3+o8zT7YU6uS0zQ4vrJOg6YC4giwrSXuKuQQqBMlJonfv1+uCE
tUE+LFD/e6KY80n/qdamLycZGyr81l1rhkbzVl2H41wE4U1hGZVUkTxPrRnfuQqD
PNMULhKbgZhzw256UPiTfpH3LhRK2oJcdTxEiYGd62D4SGXFZyL8LH/smak48hki
ZnMtR+fmN2NgFe+MUZh32LzNy4I5KHhdJG+Pv7sMxFXjPKizsAMOJaonChI1xyJP
DlRoKMpqaW4Vm94ClNHHfHk7VlxeX2p4kn9M7jQUxATMwVQ5Q/cVwgbUepshOPty
39UI0C5iK6rEeRHd254VqnFk/dq4ShQuNQzS+MBQK9MbrPsylDnOqF6JPNZhA+Lt
iPaqzVXgrSruE62YJB9HKMHIC5DSJnr1J2JXAJX0GEy6s0ZBrX5VtIjXNEHRaqL1
ouqbPy8wsuYtEpu15jedE2vZZ9BZ/DBG2msV/+beWF52Fotu6lDtYvFDP0VfB7RO
zALhWcGiWBMLwJUi3zMpl9B7c2mIz52kfVjiXofcfVqBDme7bwDRzwD41CIqrLKu
2iTWhugWPIqCzUovI2kdOvekZMimpOuPpoNUvilIPFw5XqPYFoHC+HVUOosuT7tI
ATI/I6Fixx7VZc/HnpQgoHai8wcGnVs0a85qTDE/XlcsiwDLxepH/lzhgvRloPCW
8UdmwHANueXT2ZXZ6nYE6QxUzrqblepRaDCpdjuY1w097nupz3S4OnkUDqlDdLen
G01lCHF/0eiw8uBg04oKPoauIpJEOD9t1WCJJvHtdk6Mzfm8BRHUvI6HxToQM5A3
+goVrJF8RE2rpiBcL+N1P55Bk5k4olgQK4XlQW5xp0mmqQMPu0YxdzvWrN/yGxnY
zblpD7moAWn9UfMksxKlUxm1OYfMe1Aw1Llt6595qn/cmkI5soRmcAtR7LhyF/N0
08mrLZ9MBiwvldtACba/vU+CE/J5KrK0lZ/0ymLSuP/Y6zL3zr9b/307s/fs6bnJ
vUa8l/AOWRgqjl5pRTV9JaQfjuTBFR7ZnThNMQNdjwasB3RDoySa0VYe8bGiobjx
Z339rUuqND8LvsW4pwHPKnB0rysjR1JJpnz/vNL7utmuGSZF+fjltOyv3RLHxBvb
GKvBzjeIzaZkWmOxewiwxKPZ5aczkupXcgqDdZRrATvoFlhiVQikLs6OA3LiNMb0
AJCHqE1EqLmB2yErEVkGr9xMEBdhGOvr6Z5lx8Gj+a49zRgMLo1/uzAMw008sVwu
SiFm1QL3+BVQYE/kQSN83mqnfNJxZK8Aw0yqrRpaj4dtr8miQbI0svKi4YeSg7nz
G+3ilEpygYj+V8lGANOYz2XaCAbXfGqJVwMYk2brBwFb5CVw9JQWGNNebfLc5gCz
vIr1RYpTffCr44ITjypdZY6y7iuh/UGwiP/xWwG47MJZGzuwpHr7g/uCADPazpif
JzmJjxLFSniVL1IRhBr3DXOlCfEmxUErTk6+ynMl76u32Qex0t/yEYiZMUU7/yNp
RtECD1xYcouL4782OyMgaCMcXzq1W0ntxmN6KLBVcAwm83kACQ2P+OAAUFwAKEB6
tK/M0BKU24dhjGb/YEAZEys47uU82CRZ+OEhheT2szi6z5TNUjLT8GcbBCxC4AuQ
lNXwnkhB/Kv2twc+abqHvz5MusyO52iBuz3c0LEcQwhoZM6O6tLlQ4W26FGSGrso
b/CANDBv1QdFCzRO7+HiodXi/UFLn1BAJI4Ki11alVPZtAu2iPnf2Q6GiRRxvpo3
QJZiwRRIObx49uinVfbqfntZMMONevmh4YTDko/LOUa6sNGI7t1YXrl+Mwcd7Re3
Z/osc7ZNRT1rZoqiS8X1muIV37GDZiEQGV2OBuj6KUdCAsx0bOywcrc6FEFqD2H/
KooRjeBsbxb6Szy1GNoHwNfnlx3uPR+rA3ENNRB4uC62ffu2TT0D48h68YSBE7m5
LIoCLGzNiwL9zuUZGVo2h1qP+C+w02aS95+okg4VwiuVilaNAK+bFk80sBhES75t
EUAvSE4nxZiP12x6oCZrqiDG8d2nswGXap4XwtJfnMXRMLAYCpow9erTqtAX6YIE
9Y1PRGspAZ4BtVpHTMJiAbsvcGkXlmUhuTMW60lvoZ0h4VFvEv3t6nytZeL6aWL3
2D7ogiWEDVccfx+66nsHRE3rQGzkK40klAzWJLrCtxDxNtH/qoV6px+pCLCt7qKh
tZ1Dirsm+YDiARtEESizhL5MR9vWVX8jeyumD2ZSBIQA5eEVvRAZ1ZKnOQIcOFnN
Ft3XOleuemQRgis0Wd7C2vUQu9FxfpZk+oM8ETVHVAYMfa3OyQuni/tjXaajhoYb
DG1E2xRJocZJfwfGwDDooqKcnURLY56Jgg6jlUqkCrE=
`protect END_PROTECTED
