`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XohGH24bRY7zNhK4ScUG0DZwUmCDJPWCLKM3S6X6w0Z9r40YQ9SWQIAJ4yUHahS
UZm2QdH7O3j+3hXIrutBRTI0J+k0NFceUmwXXdL/uM+J5HYoqV/ERuXv0kqZ/TP8
qcQ/sHZ3IAyyWq7hQTzv0gsPf1mSITuTHQOb4xxa8x6dd21Q2kmsw4zwKzq1H4lT
xPwKrmTadA2b2CuHnIe7OuVY1FX/x5g3fiSijKlgnzZNXaMf1PBPNFBHdGlVWdmo
dJuJYrRFe94OVplGnPIpNi1GcOgBvVYtaoOVmBqh9nnES4bPjhdkaXqx93Ak/vHe
uGiYA/fv0Zs7rr1vJrLs8hEAreuIDGdeBHM3Kr0UyU7f3glIbZat6KW+YC55wfmg
U50X4DIefdHs+vI7tvoVvDj1Li4f6cN95pFkH3hieoKFtRBxwCldfj4hJVLUr0Xt
bd7gP2Wb9qbWYhakmFIrRRxR++4cmr4ZWHvVIbTBs02rU8QcK/gcd1HVSkgg1fKa
HpmE86KeSf5NYZWTDaIWKw==
`protect END_PROTECTED
