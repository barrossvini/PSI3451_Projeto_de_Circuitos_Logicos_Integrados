`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S7wJOcesltZICiisp4fBd8JarwkAOaJHdMO/xfsKXB4zcLBTBOcJQ+9c+nnkfDcV
gWQovsAGjxkt3irTgEMDV/3U9bN7sbBIWE2XxduWS6wb3uNx6Z11eHl8C88p5yFf
XNykQT1ntt4sxpkdtanVwjXFGexVhBEb8AenGqkWkXY3hI/xntdkvrDCNnzmg5uj
0e+R6RZNXQCi+i7/GRe55F5tAueMD9sLmUiChoJGO+2zWGWwViL4wE3P09GX5R69
tEXpKKbMML/q+yJFiTAB1ZkFdleHeWZfydblybnIP9MSQdmnqPzdVGjaZyv4co14
vHD2nDSKjURbrsyWeTKOxWhHlQWyjudh/VbK+Mkww9Hcaw582FTEFxvgkqZpM2+I
bMIg3qt+upoMU26Q9kzlhdEkkBeVPbchgI92dFKI927Yy6SHs7s+Y5x+czz2LIny
MKxkfYnIwCasEoE83Qt0k99AkqUd3M2crWgtWPMC48Hu2/a6yokRtjCCbUvt2vAY
qaBJ/Ypqme2Ohho7tugp0qrpGE1OxfVOZCvN5TZnTZbV2mSn8yRNdSpAWa8cUpNl
0hYvkfC5Vcb00/4e9eW1x06BV/BKieACiIBBajNzX20wYpaSOf5Wlitsy/7zKI1S
+43uDBJc9YEzAaX/NOwq3zPqJwniW4CF9OxuXnxMYwHDVJ+/yCgNCjyz8Wj3KDGf
beXJoCfBEzpqIxV5hRAkeeJ0R+tLQXRZI3gyQe7YvdZJIlOmhuw2UGnMdnlkFgwu
N+8rwUTdHp+NOUfxsybgb/+XxJLfwF1/IGiTFvfM+YKPSnicHpJmwOlaOCzuNH/U
IYbjQeSxYle1H7RYGmHHkYr4zpGMwQWHCjOznBqmYKCKRDVp6JPtSICJCPlurSmW
LP2FMa5Ha7QEgyvhrZ6ELQxIR8fn+b2xdcJNwLKdiUlVFiGP/4bYuwm7/v5LC2dm
49uxDtOidH0upqzWK2/SPNShNvsK2PWVniERv0inC3pamo0TTM4zLOagSyP+FQfj
y8ye0NQEi97RHuHuH9AeyPwp+oSnYspH6+g3CfrcdrLrDkchAm0bQeXKs6NpRxhc
hgKlHx4F2nuiYVXvqXnAKpfTC+FE++UXWWJI7aWO7n/HK/acRQcqtpeWSBngGznU
RPYm7vGUt3x8iCwaYBqKPolf+tpRnZEGkudxBN97j/SXTZOuB9TZcF4azNOFtlbH
tV+z/FBS+nmE+Hc4DTRR8Zqs7o+7+qpcJAXIPCLUlf2cP12FvC3UFeec4bHbBe1G
12V2UL9Spdf6g//ivvafC9A3poMe4ahtLf7SuZhBSR5R93nG0ORinDzruHzyHKvD
RiXlTVqzOgZxKj+GLg+xTvRSRoUyWqeDPL+hzBLYHCBVQFqAgn4w4u+A/RRL+yIU
cBQkLxWfRiR4WVzLH+LathlqGJH1seU9Ki1Ql3wh8jGN7AZRlAg6IjGcmS/7Y4df
THU7zUs/p689qimOgJDtY37rd7ULE40D/bEhXzK6/wTyFwU2S8ZBxULQsSWj9jY3
ALoKtN9YUCP/0zQzKlQ5iANaFScl9B3sdvQc81B9LfrXQIXWaapAh9QhcZZs3Dta
PbTPAZ2ihYnzTQlnaAhBeMZYEepOQQd8P9i6x1Lgy3tFBbDmfmbC5+4AcKSM/stU
rQro5e8oiPDC9zuhv4VFd3I0IzOSA3E1wexlPIz0VXhGO7+pp4jGntQqImzUku2L
ByTFfdddQqCWfn+LPLrCZsZK/3jqdRksZwnAQtaGzo9vXolJXfF4eV3UlzMqIJr/
ZMjMrOR3HqJXndH3PprsnpCSbsYbSf/ohsiJGReRy3GsVAo6TpUhLSHVR5Sjj9W8
mttmLpbj6GytPsiGSsJMGh8Un6FfyFugY5MDNZAA+7m/2evMXk7dHTWN5Jmu97y4
0mViIC+Em79a548ag8ggdRBhLJsBAOba5ctR4XxRD088GhlumbpabTTKeIm0ggaj
pZgz458ebMrA68lZyPLNUJtTIz2kBipF6Nxifujf+9az7qtIc1Q5OlcGd0f9NBIp
LpZw6a6lMCgVzaFKOb2Z3vSh5AROmRh1tghvBVD8efBQxrHVZN+6MDDBOer71wLQ
o3uLCAdH1qmnbJ3KBTfedydw0XfwbOAjoNKDB8GJ3HgiQT4OWBwYg0Ipy1Il23jc
QMijrAOsqB6u4knye3iTwailh99InxbRqwDdHJ8ZrCwFVqBXKx0MFs+T5sizS67l
Dk3GjcyB++Es/6nJVLyjlgVtfVSPpcIHkYMzIOgU8A4/G3xxEeeAMi+YdkQqt3zS
9GRE4A0TOngVQwFrlH9L/oaUfa3IxCH8YcNm8aWTYxMSXff58bCak9wBJ7sRPCnw
`protect END_PROTECTED
