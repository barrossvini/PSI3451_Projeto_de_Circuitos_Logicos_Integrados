`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/aTJ0sbXcqaNk3FrtRIDYt38G2wB3lQ2CYBK01ejvTbfzr8CeZI52rrQf0Hlhzmm
ycSOLb6DVvZ4w4Pd2Hn6LKA21imrwgNOQ1ot2cV/cxp942OEYBBRTxTDFmE8OSBo
qgU7UMKE8C/UZYXq+qwl+TcStq4WoaIAnar/Shl14kQQdznudTUhACWbaYY+uNEB
2BryhM4FSiQAemDtaMoCbY/XpBj0FcrKo0E2yl1IFLgaav1/zJdL565+ufdm0mWX
GGn2sQ2nHwHyYmHpCi1UEk8IPxnr0fji5lSFi3xzUu5xGwaA8lIckyGDZbIcHdcb
t5ABLCKNSipyn4GZFPyEPrFQ/qMv8jRYJAGs26vHoSS/x1c4OTiJSmPlkvZHjj9X
DchvHdlDlhfhzljfoRbxm4BTdJbtxUB8mKkzkjT+45sJd6XmlyRcSwJjDcgRzb1C
kY0QFiHyr0DGEZhJsTXY0vYkPf9jmRt/HYIgiEhFQhB4ygC2tomVmvUiKEza3f4N
B2/hYSsxWWpSudAXW0jhttK9dds6V6FS4QHhuwELWoy50HBe3rhNLONK9IvXyJiq
ZR/QwL1+efyZ5oL76pRIml8/KF0v8KJHpefkcZH5OXyePkrl1xsMgx102LdJkmhq
b17NRsU3HWJ0Yt58Pg3CujRIAEPp+18uaDJKTqIVBF5KxpAerN3nQIHk/6tQ3xwy
WB0uUlA8Etko7uijEifz7kSueviVPKWhWWZP7+CfkB4rlQp3fARuH6ao3l7w8KFp
C+URMM4WbEbjXHQH82WGdnzWxxupt+UyV9DM7eLvGQO6TQt/icSPYcrWx2GdvzZd
i9tlfzRpcUhn61nIxKLoGvb7GctXduJlYVOPQcMuNwQrzdncVR+ib03kaJfxYVjk
7Tbcd5KCYK4uZzXFhJSZO1Dx41Am37ZubxjjEDbnA7BexmzaSoKsdZfVwFxmiJHc
7xg7sPY8/uAwA1aWDFNgE0wEbbqASyuQrbC0O3w1QQ8GcvFZrCd2RtjPrZx/NJYf
kgsxAMtRtYXYdSDhCMIh2kiiaNT7iaLVZl/cPFwzhsATtkPUBa8hsNXEifrgTQxC
5IobfGHVRhZmwvtD4F7L3Uugcu4iryQQFqJt3lGNY5wV0JAS+8/XfVEnN9NpcOc5
ODx16Ju/mmhSM9mbxNA5pcgw6V40azb0IgAVQ3AUaVD1KPU12puTD+cIAk/PVkaJ
jKB1a0hYMeUPjX3XutM1NEgTlR3Ynjm4QSNMqSMpfo6MGDPDTou37LfiAimfgKzC
zO4M2Vc0va7QSx8009m8vnHd3syrA9mNXfh8NBVPq5G9liwTYY9A0+tR+O4oCywL
WnYpPujL2czoUmfsi3M+b6TtQMbfJXY4bIb8DGSbMVoCF4/C1Vii5t4ifL4gDWxB
yOygLir+KAOnZooOKkUP3fayPOy0RBNCxXac1EBQxB9P+e+Az+vnL2rjV/mQFAdR
eQuPpfhLwlcFeUk7FaqL1JwB2ApMYUaIEpDyEeaKww3p76qHsTI9lGXMgu5J197k
pFGBBuEcWY95wJ8bPHyrNb8vqE8kyJthCJRo3SSvmbHxl1L43xGVYUCm7g4DpY4Q
Oz6CTTuhv/ezySeCzlrbG9W5mkzJ3dyW7wJMmUz158Att3izupo92rEZQKshbv0K
IGGTBDoohXWq+fU209qzeLIVOeusihoOjKNM4xk9Z+aCqSiXauwtREsMp+4H6OjQ
PaOO47oaE60JxScXz4vdN6MO+BmQl7Vm0aBLESjYwliu+o6RT2HP5zlvv0s0hBft
cs3XafueRm3J7P6Z0VT89sZxSTd1XYkt0GQ7cyDrDhtuPe6AD6Aksj5XYI07l9Cl
TWiH3X5Vhz7y582gx8SqQtejFh3J4dZ6sBAJVsZj7ZUmxXVuVbRKH7SslhtPzJ3Q
oGAaPWZYa3psRPPIjP3wuUjIwNscUvCypS7YumHHZiE/Rc/Kxv1IO1LERljA8+xx
RSIr9cymg8shwe2P6N9ji4um/4MlvTbj2wD0RVhPCaGAFV36dDIe5U496GzqqJrh
gprqyriCWWXPNxarJZVrvZCc9EhbgEfXZJOMsMl8YLk3LMXtxunYTm8pwwAc0oGy
6B58ccFdS+3d8Oe8o3MykP7Zf666Vsd5qGI/mLaK3KRYPwf7vqGeQhwFCzQcny7C
7vkP5SB0wA2VzfBBLsI0pdO82y34vT/GuiLEaoygyf/0bW5SbIjeEttXZMrkJWPE
9/x15JrXYi/o3wNjjoN/y8TLqlp/uSFS40eeBjov2d8Cua8N2eOAff8h/uTO+aqX
hiSDfCEP3o8S55+BQLREpkfyx7XvzMxS7Bw6MJsPDnOPij15ITKmr4D6E2zZCljP
Tk/JZHdtYSdw+LJ6fYwKPsc9Ke8PK+4lBZ/wMdbufpOdHFRXjjZFaBwz8Y1/X/c2
1Pi7G/aVSxPtU+2kB++fUqupmIfSmDKBOani8cdQ+X6+shJbfsgEFSS59VCyVNCi
bc9jnz9BFAB5UPcdzwRuA2BGca9R/QqCwWCfPaHZaHmNtNhYrh15RTZloYJ6A+F9
QeCsMIhsN3ppaOFvebFNhNpoh45T+LgtCUA4mQcukhbFTnN18Ys5BLPM85z82XwU
W7IqKGgT0dsXxOvUC1smkumqOZpR1m4WGi1FABj25/Z8/5lI/APX9wU4rU9TmrJm
rxDgv30jD8/xHbzTPRbniXuj9eiq8y1oxC7whe9AX8hQryeE9dkzc0ulmaXFRIql
4o6w1DQhpKUB/2FXFdodoQq8/Ctnw3SnMsWgNby4vFYyl9phNDK6d0UIm5Qg/mdo
bBUUHEFmc1yG/tTcOfrDhy9Ym+60MnCBpyO2DRdlJc6JEUnxlApcG5CT0UWcwmvT
wQhgI8+rgWh4wt1a+1sVscNTZbDWjYxuUB7SywP4CgheyUdmolu5QI2cbbS8JYEU
LoCacjRefaBcqSse0aSwXBzy8/+ftnzKxgg9J7OqG0uLxg5/cBkjlchLgLNOQr/C
LJOQ5k2Z2V2lynkKfaTjTYq/TfDb6gITxSJBvarwWI884yDaeKo8S1Bwkd603FEu
29slQQeWci8z5RMFWwn1G32uyAJHtnD48p0e4udYsWzcjjj3n+nbuYoZ52RkS2S6
0prr5CQ1xl9Vo3cq1RFwRR1L0xQwBQBjFJsepqy/tB/ziivKnkr3aTz5grPaLRgY
uctkqbUQTCgXv3cV5EasRyl8leO5PfGPul73csrpVmWfwkhoPB6v3wsomPhneXGo
H2pVL6a/Wk9DJTl0zFOWYdpmQkSqMTIVoGuhSv7KlCQmqMps9rYBwFeFFS+EU/wR
WvDMMCyYWwmLBNSRB/QxYoa3XRX2AA8vbDAMQqaUrGiOfepb7K6hOrMyaFVfp30J
3NbROM2wneCLwyQ8l+QA9SVGcRSp1MTIUsauQRrl4reD1U5KqZVU/scAGlj+Mdfp
1FeTFoZ8v/IqXaOhFOvqmRcukS7/3KNoD6OmYQFtShmU6IyWmvKCrMXGmeF352fh
XZzf3EhdH5v/vpiAu7NEPBcrEHetOgqOJWZMIIdZt1o+qpclrvMJraFdKmFsX5z/
mLOdKJCGl1FMOSegQyObfBJqNIsHIlWkX5vA7izLwlCSwkT6dVn6LLmYT5tDGw7h
eP1b96Lejv03AHbOmPoIciRd9iJfy6p/15mCm7mpN4zd0QvTTXbuTn5CcAhjhapF
tLBn62K+GafkQpJVA/+0+GR+NfA5zS5yy1us50nMHGuToj50HdWEAqg5B8ohms3i
e/RejnCCqtvw1dlHCE6Yc13oa5HgV2Sm0d+UxE5x1u43Iof+PlT8eyBDNs0gSZLl
toT8g+jiYeTvVJ7yGhdk3FnZqYRfkfmCOF4KWnPKEZzOVmZcJJ8OcfjNvujgEEDO
ZigDdUX76MfJJgfqNU223sRlJsmh8tUZOgfy41PrwGl1hvm8OXiGNrq3E03NJlIJ
IXanZAZJKR8FO3kogW+R5d5c/9Q7Ndy7+5qrhw5BHJJx5UNkuJ8WfXJIS//qPZot
4J2l6okLC5cHqh2MHBT9IYvK5HO+sr4WGzHwBx2XrP7PSJPVYb75/u036DaVUnAM
3HDHSodv8sRrBgqivljWwesDOQ6POtLy9crMgLzYSZIYKB/SkZLd0Xa6Nv/VVT9/
xHLwdDr/71mPrznns7gmDQD3M4oWoIiOfGGHuRfBtsxm7/NuZtbIx9BiuNt2K07B
+0QGFpjrIBMMy6csW7eogVcukoQizhmqIZZglNNkEla4CR6aRVyMvd2PkiIUtKcj
reHFOWoLDQVBE2e/M4as8bU79bMZ1ulRpid137tFnq3btKBraJbeUsdktNUTMcwr
KbYZpQD5DbIKJ4YaxLxqyU1PuIx1zcFJe/6FzwNo84cF+jLA/R2r8BxezjK1Lhwv
G7KizgIi3LyXvvi7P3EA7Ld36uSLjBI8lX53BUef62YvOHxSTjR5N/2objnqfGrk
0ZGTxZB1Q3bA5TNnOG4YzwixbFgGCA16Beh/L1/R8ub6cS3RSebaKMbSYpPylhyK
lLw33TuEBEqqpBwn7uDPh4k8n8aQYXgvMlHdZJxQ/jYEqGw4KlswlM19EGRTZNig
FzZp6xRzXHKefTEe7bVZC0MfZdJyQaSu0L4V+ZPzJauZXqdhlYzNng7zg0ZPYtzR
iLE4EKyr0wO45+TVZbjpoRbbVl66vxUYKG2dTsPT4NcPP4dQrldJLqGzEhjS/Xdb
rvfVMT2Ug6EvokcGSS3DidV9U2S8mcg0SIyexUs5hRA84SVx5e7lgL6uqFOHHyN/
jw9SfTiflS7oC916pVydG5FtoJQ0yvUbLcOO5GeLUFEmvzjspuBv2kYef8HflIfY
BozLxllvPZJW+joMK5oyMGwuzdBCLNjcyC/ZUhox54hpUJ0MlC4bSX3kjNJI/vi6
w3mRr+ckYJ3/gugO69QnF9N3e1W4gc380+E3XjoJLlMdq2VvhDfXKtF8scWKKF5d
h8088qPA4Pf/f9DL9q18SV6KgzPempi+WGKtcEwADBULL4Zvvsv6k/O6PaxfBQwe
TJfh7cSlQeIYX03qo1776xNI6S0gVbgJBkeLJ66P2cxCXQafLukUdXkk7y0MPOuD
DkmcITb8ZUw3TrZuCHPFQHeKtz6QM70tDVBdYtNcpHV2I+iJUua8tNeq2ehPuNEy
1ZIjuQecy9bmEdL5lVYNSm0QunpNLTmllytG/s8XE4J8Ti25DfSs0Z1sdoqyIA+F
tPZIxSvAyh8CFQR/8u86Y+aCg6E1CkPiIqEAkJ4Kef/uAWkJ5zVXboIFzRB6rTGx
BHJTJ1TzArtHs4A/g5kN62lgqdu0nX2wIpbLDgHuREH0qqkq/hkJSICrE14eJeH0
SD1zAYugH2sZchRaOVe50KU8eQMp5PUFy3BFpFWRlCwqVeQx0QXUh10mzzbgEEGx
jddEZwhWAy2ajX6iSK8MEouqDidcQw+umg0wwXEcSlk4p45Hpk+EQJq4VCmR/weo
wV1qZPrcGmee3mk1Iz00VX+Ib0pruGVlEBBKCm3OBBKsHZzFZUwgWLktCRtJn+np
8yBlVQKRpM3HsUaBROmPW6DELyASEoEDOF4rr16px29LoaTo69W8PWo73pMmbP5l
NcFBAMJmGiOpfNldGeacB94wuitI/pJVrkbEFpRCTJcny9LZl8fM+dXinm45DeQ4
c4W+NrW7QAfM+KJMGiRms37d1/CAfAJqeYVrc43iaWFZjbE8BckPllidDNGoyJSo
DvvbEagmxZnHnwzZbWL9fT1yvC/i5gauMMq0Yg4XgeTto7QsiJPRwcS5Moi0rybN
p4EfEIH/XqyVY+NmpZA3kn2FlF/7JPFFQ7YocM1ThRudMBNNTv5DO8CFLigsl/qp
7NNWChXZE0G0hvW/cLklphWLauKPkhLJ6OfQUcf7Nb4HAqCmAd2CvOj7bc3CTooC
pnPu45Ba2AMVu9UmnHkTjZ/4xQFPAmaX2PuwTW/lHrU93c/MO+shBn9Y6JCuT80C
XxxowEgYRVHZ/9I3nzTIhXiT9WvmOR65iVEoNL3PUJLfdm7PMwX9CDGO0TexlOc9
2n3SJcrkZ5EGhnNGz70o23JPCOHfl/1WbGOm3PpQeCLCeoKmb1QdokKHc+b36kwL
vaooAHb0dozZbtiQy2+x7YCb1P8a+T5Pwmz/Hrg+n5RO+5sxHFn0W/jBWUhsQRkr
QkIv4dYzAOqEZerNzmX15laZMZWwBfR55y7JCjLSxa6CmQFMG+ScBY7yUwEZaxFC
zuUi0licdJCpCi54EE5VWn4Rdb61mZBtd+wf0FstHZFltrxckrJpedAymYR8GzRI
5xtK3xXH3HQArYYU9cxa39BVCwZAiY1msr8ujL9eSq2Qcjn2/IU6DaE22cAtNvCL
kvMxYoVSpaGLVqFW+rCCbjsshEu45j5TWAENtx/JoRwyEn7X+XkNXNiVediIf3aQ
HYUvP8M29JgoMuKUhkleS6bX2mss1/FPwoE94UxzqeJiJqwku2X7cGBrMsntAUwe
Mdz8D4DXv5TEgSe9Qf2J9KyeuxmDx+78XamfVZA+usr64BPX0NQCCFrCLYM4tMh1
8nOqbliLbsvKrwQal3TK/gdHnWGZuSZNIMqoumdRHQdp6yF3rMk5+jcfmrwQvCAj
dVAiEmlmqfsvfjjUEo4KuvwrBjQ8kmdUC2t+k9LFNEeqHeMxFwf03Hsz1gzRvmj3
QgieM6jxeujs0BQtHdkZX9nWRupn3JEFcQLH5lLN/TpZw+pDuBm23nFCP7r/Ji6d
flGXhS5DG8EKxYGtX54LG1VwmPTs0bcIvyJ0k81tlxB+oPT+dYZzrK1J9qsEnpV8
TWmFfpqqLduCJHeYcN3wQ+CzkWUvv71qUCHkvI1FphlrlH1HLI2H97H63L9Abn/2
NVmh3G3o1CkoOZHmyxmIK+lwlo0hZ0g284tQ7r07xaiZYgaFB+um74cjFqeG6Owt
cH22X9yaXbQx6ZSXije1wXhRtq8VmnjPyTBpqL+UBct7ykhOhDb7aGJ38iscWi54
xHjapRUABnubv91TpuYghbMRIKJvPXXhPTHwPaUHJHfWFFhR9Z+F9NLZKRo+W1kV
KKZDllneU6ZqAhfzjYxt0X7dQT898TZrjJZ1arNOaOv43GkhQ/+LDonboTOMD5Fp
1SvdDdXaDIrR/VcU2ZMDTfHK2lp+jUBE5Her9n1Qo+CHzIBxhrOHPudvcfB+tH4K
6ucWtSsT1PPYuY0Ag4xmXLHNEHbgySU1XoiVcfASX133evswjn3cmQA3eHgV2NR8
/GR23HVrD8sKXXGStcsPzT3TV4jMaHZCXwNTwrC24fl07EpHgcaT2p3wu9j8/RTt
ILpUQtZ5xWuyNSg8YEUkded1v1MT+Rw6XvQunU+/yVuZdx2j1oiVoOzsJe2n5+ub
OJYgN/3hZsieTQ4Pck0x9ZludATdySI4uE8XRNcA5PIIZP09gYm1huY0Iq/DwqQ7
xPLzK1Wyx7F7yvugj9nozFPFytm4KQJguiroXNg4xjAhhMGgLUcbQKT1OP4jZGFF
U9XGYJoml9wLaICGFLDlSPpoz4Jj0pDr0pyYcb/lDIrPkJJ3LPDsKQHxbfUvq8sz
CKq42r05zC9/zC3LfEj0ua+eTyQDx55/OllUmoHiL3KjHnUmKRZzPAoLeoQIgWn9
D7JHL1ucOC9wcJWuN2b67FiwLP4PAVMFOWhCmaq5g/4WM5Q9qv6WNFmz2W6nMUkR
gSCtIDQ4Wb/ok2fu5AyXsbotkeykRAHM+imK7UL8csUPBpU9pDibEA7DUPGRfUox
lh62hKUGEhP+yGIoCwkagATzY2F9E62buFgS99jHw9iQtveNNUfD1CbRfUIKi+2O
ymfpDgn5gcuTiHVvnOXSxN2vLb5qrfxUbisNuqqJjavFex6S2Q3mziIewiTdV15e
rzQn8si5Dfzg7N/ccK+FOxNG1snxZdk4qjj/AbQpZJTpuy1PPBaEsuiNKleyp+bT
fH26eTKjmqU42ebmCsqMqdReSXBhRdLsGv/Mxpe2Jup3gEDtChBxG8RE1N8FhaL2
ERoc1ostaljYI+F6x1hcc13VdDojtu+oENCSIoPRKmCpLqqhWM+gTDxYwzw64aVR
g1om9UPD19rs0EqlmV2abfqJ1vrpxCTVI0bH2xefmZj/VCUFT1FM0hk29/V7Ia8n
oHqg23xTWM+2ldED53qI5NaCDuxhVXKSySoNHdalvWuaOUVANmyFjfyXYqEo45Uw
QFWl79jCQK/+iHUW715rGRV/iQNR5cMScnV4OiO76K54KJERYhoUI6ZvFPAxVd95
ujsttqR3e6Ek9umgxvYK2jtg1Ws5pS1AIUDycgHnftvBYldsnfF3SZADELvZYF7I
K5c0sKb7tWtE7zgIZd9KB+NkINLMLzQdueu84PwLvOUBOwJDamBpWFRo4sQw4N5c
VqY1wWyxoiKfNfHmct/VuRrDDTl4DACUDqRFc/Uu//kI/0MLgYj0k5XpC9/n7tNp
U6Umxo2rXumuRnfRGT52Ut9aVPZeHibY+vJxhWmW7WLXcpK/8rl2t1tIkQMrsLVA
VDAItFocGP7nrR+8fhWxTobI+87GKWehUkT9kFbchSRXJKgdXMxFRUzcgxtRdNCJ
m3YDHHWqElpKuPmDcv+Xae3zi1w8DS6+yOJSYFQ9OxWVlZgcFH+cZUMBOt424U0B
cMsFbu3vRIJ/qAH/WIhw8GgXGkrS7+dIjPdeJeHGX6v6z1edSuaboBxp+fbWmOvA
WZOwLkQC98uk5dSB70WiVzKxiKzVH4WdjH4UbzPcl9w7Xtel++dWtMN5xEmS3cxS
OevIidRHA8jXkMhQTgmo6zx09/1DMdgf4xspJcJMC5dMw+c6g062jezxAbQcBLR2
ceRYJbN0drUCdX7q8r5TAJwN/f+vmllq+t3rMOYsMtig8BJ2IhLu0ZZCJhyysXh5
EbUEczq3SfPj2dI0haGOv/paEqB6YpglAYFLBRKXLQ4sIq5IPnBOCl941dL23cO2
2YV2W/i26yxktBSVSIDoSGwBbZ/9/KLA5HbB0oaBwvmNYOuEj3aYuD7Ekhuf3AbE
blDQXg2euhJLyEMO0IYLEG2OAzeueO0l64mMDWcqKBtuq5U9KnaPN8VGqBnWyElO
UDLGsjeK+yP45yhnxWpeB87fL/bIFXS242gcBhGe7YTmtwz0FMEPsezbvxuJYJL1
ivtYD93NpDLusdE7mCtmCKI6Yc1iA3DFY0JecQ6sEuqNcbT2jfp/paaBfv3nBQS2
3qneuXgFueMbxXAtzIh8eFm3AUHDatcq16Dkl4nM5S5jDpGVjNATfNgf3WpBhdCK
52HCUxnJodTXytm7b3uuFwFREA1QVeZzqNnFPvALYxW4JAG+xCghZ/78/97Y7MbX
fPsEa/G4iEdqlP0i9Ll/dc436Fw6UW+Anj1WUdu6g/zVeTOscyBxtW3grAT8pmd0
kMiA8jFyADR8sl5NXQgZMK7RQSq9iZzBPqYM/OPCFLlPBDSVFF87j9latD7Zzfoh
+zpLnOFyqrz+vzHDae8TNipPsBkQ3AGQdU3IuoZ3J+KEqx5jjQCmlsq6pTBOOV67
2tW704C76QBGxhWMFCEdfzSvY3TeLvr2+dRqeZj2tRVL4KmyYSH1e7dvYcfMk6V6
SiUDbDT8K0NCaxheKXjQ/p0HzWUP6tkd29+xoUf70Zf1rq/yM22d89H6gadw7jOP
wgojdAzyEIpVW665AEU0aEwJgV7p5ivxgb/idtrDKrs8sSq4XVpqf5IYRVXpmVLQ
vy4pAQ3FA7K/WJ3zD5JCwRR8UQcmQqoFDKGeOIjtyOKsUdu7QyqZXve2FUY9t2hm
mUkGH2GAXDrU6AzwBnZIrseH+c/F1Tmv0QAzAQj1uC4k4ne2Gdl7htxpvAd3ivNf
r1WKdiXMNbF0DfEPgVPNBbzOBR+kfYZh69I9/b7IsBDNOUQcFWXlrGSgwhFK8VXR
5utxJDb7ifCXcx3RY9Uv7pVXEY6KcfMbwJd3nB9qY81DylnsEl9tvTjePnSA7n96
URDzYsfCTeBSWepk8hlWP3meGSSnIeprcBLcKbU+26aQqw+YeU51jOUG+njnKB3z
D8Hst3tMGXS8CkGm9GwLSQB52QFrnb3LNwvYV3lu9pUDZ+dHV567hJH84zA3p/nI
yVP//9LB2kRs6sdk/okX2y/aQBlHK0I96MxOzLZWNbMmUn7p5UNo50NsX0+I8MWd
3a/vgJz8Xl47tSaVNcsWIdt+nDMrans4HuOk3sPjWDWAOuJzIFSHabeaB5CIyYxV
9NhMW/wUvUBSextXh2vNj2dtL/d1hVDanBWDWhttM6RT8Fwl7ObqaDVHGBtNNE7s
XoLuwaAsd46loIwnTl/LfbQaka8wqkHYWECGMEFp8mUwNXOMAss5uTaK5ErOBwR9
I4Ri+zrEz4aaqf0ZkRrBljpa7puBv4iZj9ma8H7zzZPkZdSlflvWk0a9hzj4lIyX
9XLvbCYGxp6SjL5mL8X/T9x77gO4RL3BHMtw6ePVFs+QdSXbKaNQQ2x/dUwQDA9V
rEuAdnDL6+Hrwb7hH5m1H8zAOFMVPjga7mc29uh0oiAKePRUoH59ngVZBt+U1H9H
9tlHr8t2/xDolvNBqMpd/plzFJJ2Jnt6Nk7RiZmGqRGiqF4oNAyhlaiFHfDAEOTh
P54B5FPwWRN42PJan6FTiWAEd6M9Dhl0eosKFJ/LlTf3ufwsQ7ky8uXKVVXBfr9/
9jWAZa0viKU/ilV5kcZeLHP4e1iJ7KwXITgSe75wFuTw/OW/dqcD2qaMNWluHABg
p2oaoinhKwE+oqj0oSZW97RBPDzb2lwAsN0yhdlfefsVGnAUA9Q7piqw7qHyR7Vn
`protect END_PROTECTED
