`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LtEqjFelG8pqtOOLmc9GWxhLGujmCeut0CUdDql+L+noYsCXYo+YT2aapDhL5oXt
dHecT/HhZ02+XPcyEICmWWpqtzsHezB+yf0R07SBVYKe36RiLoniipOkiDf8xo8j
JiiNeHYzJVCLcGSOHNXrd02uoDQxJyUbK31KS0w4T6/IyGNSTREzqU4cQEdzQ+5H
HD5YrQ/cLz54luSN5fkzfuPtFGZkxUn5aHhFDxlppST1x4K5LiXyXHke3kR6noOh
MCQmIZYPSNZlJLZ0KAMdWyYSz/LGUwn5PH6wBRPdk0KaJiiysnVTKN2Mdjzn5lw7
vlut3RJ6fabT22HJOG1aNpN/feKpl9U3BJv1lKdZWsR1rDcYi+BIgjima6aElPEH
1uXY1v0LNIdPnVG0vu9GoG2tZoXHBE9YbQ+GtU0eLBNb3RTaSfOjgplS8sSVG2Me
gZ3peSqJUtuncmCHjhVR7BFpyLId24Ylc1DLXJgXr7xpc7zFlu3X5KXbx6AAHk83
GMR1jbBapncvQBH3y2hVj+t7QuEdlQibdqfoAFVHtjhrTP/o+97buz9hU77e1533
H6uqXb372150WknJEpvfn4EwTr1BAPemwYDLcHP4CdI8NqK1sUgwq3RyTVf/MZGR
PPhL+rX24OXsRQ/De18iXQIgbRcX1vwul5CeXKfm5uNuZA5N33spGQsLnb90rBdn
w/AfNFH6OVrmYi4i5+OMJnETiAyQ5gG0VVsSPXB4tYtAKecvI++6EcE1SWstCYFw
0o+u4NYDi+QX4zS+qRZ+7wBtDVomdyJffi+IhowmiC0XR+kePVG+NhtdpjPD10nT
4560Jyg0+u9YBZmCTtEGgg==
`protect END_PROTECTED
