`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EqeFu6Q6oMevYT5BjScl+OQev3EPK/VDElIQuO10cvOlgubdJ85Ye8yqL+1514n6
T9GdgISzaiol6T9XZUk4v++jy3bdzvFVSlHM/S2imObPfPOFDAAu/j4yf8WcDgma
6BHuHlZ9RP76S7lfUp3w4NV8gpJJafpJhiAEx29Y6xPyyNhIq3Erqk5NmugTRpjc
LleXoakWSjsP1s6ve3hyyntuDyX2vdlGF/phY4hc8VYa7lGLXW2roJZsx5/XUblH
PpMgmKMdsaA5uLyZus9VJPBvBgqHQe8MET9cxoFM6u0L04ZL5ORXCy0Bc4EvQmad
W2JG96AuVJ2u1KDw+hH5hpSIw5/ovZS5AO//J+4zL1V1Sxen6xgD5Yt5mrpj42eq
8Yal5T9EYfNIlkXUHguRFvFod87hwL6VdRKdwK6qK6DJSWaeY1mBfXdOT+6Wc2WX
GazeSv3Lpk3YAGeRIzBAOtdu7WErZUizTdHJ759yj6clnHba0BpT2TMVkFtox8Im
rTxEs97CZvX1ZfCDtUj8ll/1DIPauTnQetUBKFd6l5zhNw96FcJrMBAM0d/AXyk2
cruCO8RliHi7Jhz7+ogaujwGZ6RfQ5X64nKi59TPsU/fpRur4Uzm4MZ0y6VKBzIZ
ujZs5aeKAf4HK8Rh87IAOjIOyYXLzYc7Io6+U9QCQO0v9uFdWnvGhyPrLv7PPl4T
7xOjcIwl0T0BNxqaP3cHvCfgrCMbtO+Mpd7QgFm3W2KbLT0PjsULL8T+grn1Ie1D
r+zKJd+U9cCFbAyN8AE7e12eGmhv7F9bo41RnOmzCJM46DH0SG+G4z/DVKmhqQSJ
g8nMSqszzFGLjFcnPrvKzi4Wm7siDnVGCfDzVLLdZjByX6xWLvja69NFXcb4SF3q
Ai4NAlOsZCCNabhzOl8HhAy8joIEm0NVk1j50oVTgYHu5uRDyC0sN34LMKe6SyK1
JewalAayqa91ROjBkoVJf/2QvRiVLD1055F1EIIQWf7dF/0ZiJEMAyhpjvixNNoj
iR+dLh+JTjhHfIPivkhdyO96wGT6Vm9ywwVOc7j8zsLs3EXWkASp+EytNNieyAU4
E3C2ksKvhmEIlM88fmNH2pFQRxDBetcmfPyXjeYNAjESLkgql5joU4x1lyhqLugr
a8zGU/wFugpKaQxgKRH6lfPFMzRN41fQVA4DXdEnxG0p1x+tpBBVKfpD89UasINl
oN7ngOmtUKvO6WTu5EutZQ==
`protect END_PROTECTED
