`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BI0Qx8GuDXIS6zMxgg8Qq69gLVI97P7vjPStzD1lIUBy6MaLqlpLrTUVK8EsTHno
MyixmqJCiRV3G0BnPyGHf5+KeRGoiLWXbSzDM9dJyo3CL1LqUU9pqkrex3bJvujL
VMsw9kuSx5nDX76ufTnUKgJGoIF/jKaAiqnVSOWrCJxb+KCJAfC0Gt2p397Ohday
ZbSgr4wU2rrcLbe2527qj/1tuMZbFnJNhiSUlczPzr6eteDujwdW8C/ghTX03eP6
Vq8uN18QF20dtDeyF4AXy2qvVhoqFfKXQ+Cjv33XNPp2fo4fIIyqVFQWOmg8GgaT
FYPWDhspGo8TfgQ8XvLptW6/0/0Vbre9w2Wwg7Wh4rLNJzGo/pUrGJFeFNOJ1l56
o/XCgs0lbMNnpH3GacHakmXAXQQipZf7XPmfKmmt2gGz9SqcXAvtnsVXxw3poQq6
uQxyXFykoNMC9d8idiRrnatfacFphX02kYZbqSAJn+n1sxiJHJw5OqGFeLL7f/9J
P+BL9gNnty0OBXIKcjea5Q1kEzFReZi6d+zdpYlZtfZYgJ8tgeSP4e81GRKjxmB8
vjLGjB5ffS8cByGZVR46Yx4438MU1De1WFDV+ipPaU0Q1Wjo6nYlulrro2sQ6Itm
alSUdxKvEjmhJRzb4ZKKmPPI9LamDD4a28LcOm2r2+5c2n1UBdqEKkrFTyqmAY/k
Gq6mO0rihW98WZxyOjWB5ifUUBQ8j0s7347GlSyl2l3AoMI8kzthFJ63ZSPPHRFk
+9jOHU6wPjVHGOv8wIUdk1jELaOkGpe1+4CzzQLOZP1+2ADvYpQ6VkzIw5F71G0k
EwkSVQTDXYjoh9MLOllsSgG9AmHwjePIyHIi82S9htTWkJML7eVox6kuKoV0Vf7+
Tc8rOoLRiEyN1xY+61D2M4Ee6Oq9Bz0B6pVvT1kNlQZySDxK47mWb2SY8LAaiAYN
HWribAr+tc/uk31lbbeBh8rlF7FrOWOoiLkDgzYF1DLNOIO1QOpp/QMCU9cnzpL5
TyNqx2xg34R45Lsj4ph6aiBBbZja9x9OPECPj9n4DUjVjgbv8y2CqKLApCP/BJIx
F6oIfsSgH8tl9bmIeg32UA==
`protect END_PROTECTED
