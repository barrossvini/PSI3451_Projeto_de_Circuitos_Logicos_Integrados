`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Noq/2WSfDJfJxuJuyx5/JQFh7SEJfvhaXcYmb6mCoS8qcv00V+7CpODYRzY1pvyj
1s/B8Zh8PH2sNAeRM7+pYV0LfmwBZeavXiapeYuNsg+2l3zmxokRfsp4jW5N4PTc
+rNffeAGryMc9u8fcZCDSCqDwRe9O+4lE77Ydb1GDYop+QQMQejjyEI1Ik1ZmR0l
f8Cn+GLvhHJsdOUGJsPDDldoaiWrLFxVijAgvNpmjhiLGsvTEydTZMAg8PHJ3MdL
6H0nmJx/bSsH0FWvhcx6IDC/YEy7/fVQJU0pkb5y8jdusHuuP3Ov5+JA1uf3Oa7Q
E+trlaf3yZJMmGGlAGsaP3l6fjObfkav0lxOYPU9cwK1kGCsI/JaoVUB7DGcxl+U
l4SjtPtDF0no79PP56fCPOuioOao7Oa5Vl6DYjUcmoZNZer3bQ+UL+QInVQyVIwO
8dQoaYiRCLxubpH/iHjQNY+r8j7zR+tRV0dCFT5kotIcqzGM4AEVo4ChF+TfH0ya
r5KtxX3E78Xl26wVeGa02eSxL511kA7aV0Xf9xXiKOn1HzO5HsShyl3bs9YoHvYx
vRwgBsDrQWmmky9DLRY4leKFUi6QfuvecBaqphYL9ct5qZNWzRQn+pAjE7CQqlks
kxcnZlKAzs/xGYP6gTKmzmAPl71BJ4s5I386FAqGEdrNWHz5hUANOYcmtj45NS3N
6SZgvmW69dBtrYKala4e5Os9lJYlcdxm95/C+HOb9GkUG0msrbDacGXMbDxeDNBN
yVhGD9NWYArD4aftj+ya45hQKrThIMFvhBo3vkb4fQiJp3xnFSYK/r4u22jAOEin
qA78P3YqKpf4GWF5s1gO2dqeMoEdiz7doS/rFptWM/UPni9MWZ88yp+uIQH6ZTX6
+PJqJTId3jjYio+5jcFgRv3+XPes/qudjWFgJVhgOtKY3dWyNH9qLjldUyPT7ivC
v/iXz+I2IbG5r7kFY7C8zPv96r5kesD01QUGS+/mPTTmx2dk7rgwQwwDmTvpq+sX
sEhcuGF4o3/sfzKbS0b3Dh4YSMkcjMZpzEteQeI9kb/cvniJtiqRI4EB4lh+4iOb
lt/iZJa01vQUieKa+S3PMWw85Q0mPXq6S1PIjChwLjaYxDEdyLrhWSFB2qG2tb55
K2EaIB91F1cEICx0uEHxEI5h/H8lDffmWrE9cStKk5SdwTYa4ZCylHPiocyaaoKW
opA5Fek+LIrIRCK22SDe//G12BKrf/7PYVkgm+4hZnWpfrgd4RZ1165tTiUab8s8
sk6ELeQCz88AUKFeEdlDeOW6ieKhxvN/1wYTFUN4aCw9lS+Y3HjEYxFwMTJnbVX5
EPY/IslSW1XTm8+5UOnqUsq6WwomXs6eQFzjEhiWD505B+JDXGQCMb5TPnVYEOF4
dm9wTKwFreceUuJqoeAom7Yl9rfZDptheP0qmFJhj3tRnu79C5gSrTbiKShHN7lI
lYGwN/NAuFLbqXYGm6fIc0MEsBATmNeL3Q76rTJ+qEFIGXQqccDPxQUp8DoSZCwN
vmSrGctO/7PtnPAwoDBI2oFO+G2LSXYRE3azjgmnqnA0O1Wr0YBxLC42iQNunOTL
4PQzlpcigp+3YmCqbHme+isLf/VPvcq1KRfL6NRNTWCQ2ZBbkA0O7Z/UuP4rxhw5
xNIG8MMfc+K/RAuPraNQ5Ccbz3a62mMUpORKTIfEXZYIvfbvD5cvYYwLVRLsLswi
44SwcRSgPOkXcuh9Pb8RvGb41jb2L5Epw/fSntlWq97m1UHaVw7OLvpUrGrQbVsd
LcOEWv62x0/adw+Ne4WmzjriT/HrQlQ4jevS9gZE+45lih7JsET4zLX9WhvsWjKk
9rgbeP1PYZpxIgg4RY06X+1YN7VPevMXYBCFSmWTZzKaUH7zLN2V+N+yfFIQXY0/
4JW8mYBhQg6PL5aSka73kiikTT3Y9a0/nTzOlg8m2n8v4LSMbeyj6IHoBvDnFt8m
cbGawygjOO8HDIEuYYPR0Hm2+Q1wx2mUVBevpKxeW57fomYhwpi3xlzuBDCLjklN
6WV8gvADTkfDjMD84JzkXAX8C+CAJd+dDneTG8GOb9Yd+MfDMkQx2bx4bpXKs4pV
7AAzR6qkZi255CHr1qU6E3ThEX5ziunxu9ZAKiD35364YQJRZCVzHV7N4XM0QLt0
N1OhzPhoK7FxlBC6sTaoI8n5zuswNY8UQKTFL0UPHVb7SozyuVcqqrAxuFsHFPp2
YhwED/RpfVMealLBYS0azOTliLk+rHTjllKJhGZyDHkG6mu9GZNq7TR80qGgsdEY
ntDY2SleU0IzEx4949JcmpjtO5sa5P55rb6v6FDvPy4apV7NSY8SyGdMT5JDSpti
ZXidCcvZYZ2awWFK6ka7fYO6mV64RhNCbjVWRtnqA0dyoJUDeINNuZtQq/D0rc4f
Y6M/bxqRADXZaPTTkM3fjwD3ni/YZf3cuoUlVp5RHpN1+Ke/0BKMMWE2QdV1tpEZ
NL2GULp4hMIUKgCWOrb81vNmrjXElAX2bUrBZdQkNYnd6DxDepTZMINfL4KgAgmY
rdgbe/PSghJR+MYWQel1TEJ6/TMds8/2It3JoIqBlCz7JURMZCEMtLop4ynWiX42
YWuUjjX5jzamaVntffbFQpO5z14ZMObVpLzPsevQgBrUSisl/7AlTuPqgrB/MJvQ
TOqClx27RnOMDOtkFuJMv88tv5nM+XSqUDVI/8LlZZJ1PhTHPprexgzY2pUAbNlu
+wIvK/EHyoSbPgnEWt4T2E49DEk1IdGzDEvTKMH1ntyW8O+hZ4JuLn/W7E76TmoL
IkVcOi/ufco7vWmGc/GH/Vi1HxPeTFGQxD65+oj3LYi71Ht75s4wyBjDR8Hjh0Nw
iiwACUYl+qD41LvPI7dZ8Lagf3zimrsgIJZIKaS7g7VHakig/c7GHN2xPKha0G9Z
PVrfDR3k8pz5uliC0yfcQVq67YR7kNzFxcTP/Pb/Jm4TilIB8zde3jIvMDQVycmP
deb97QzWeEZ5gko4rwdB15SVuu1vr3adn16K45f0gDq00ZUdhxNhgt/1qDOYfBAa
HuKHw6JBvgGkLmhgXpPhb3h/cA2rsQ+Vsl+J810p3aBBJ+S/X2HXQWjd8Za4gI+g
3PWp6eIJPdeKQgkR1d7RdYvPtG/63a+Be81l5igf9Wd2ohPjQYV1wCMdBqh8KRnG
4EV49CUrqu6Vp/OjOigqJuFurFkUvC0lr3Aj2hSPJtfI1u/4uw9VzSGtOCGJUBX8
GbQyYBDVfi1nOHczi8zVjumPxmzcJrUYjBAIyS8Wz3lnN+XkUFSHXNVCyL0Cj43X
ixqSEsjUynphOumzzwtZEpl5h0RPGIT0MPdYdhN38HWC4GffL0LlwqrWJOdw3Ac2
u0KYlE+JwA8cngyLeKsF9QpSACErCThLeSN9C6wGAl3XryKQcELbN8Q4U2AR6u7o
9yFwLCkAI8GjahUzn4Mh4pSrlIyCYERjqtUUHC4yiiHmJaszVbBXFniciu63qRkI
zmEqT2cT5MyGFZCVX04JRyml9+GR0/MQ4wlBJ1sGZLpVtpRJ6lc69DothI0ZLEtD
r2qbfB/oRT7E1ND3u4y+LYtchBkQQqJQ/eYf77xFUXTWruaPrhIBam3dgt5bXEsV
1PhHXrCORZ+rW/2gBxgrLCQjGholIAIUG7TSfYyIS/Jtlhk4UOuh9LE0fv8eUz7O
0BZHjGzr7oyL6FIluhfkj6J8OC7nJmWi+/+YX7BNO2PR6zyZmgPHAN0K7GdFSAaO
+VVkH/q/8c7wq+FLbjI5juH7NTv3KMon3tO8s3XfxM7xUmwD4AV9TO8hkuQ0Y6OE
PvmEfUQCTcE2ydn9Tjyks1Zu3G7QwdyrVVQ8u/mWQYVq09LKVzISYscwRqy8apZH
YMbDBfz0JWVXAJYQLfk7F1MCtBJ2aWHQv5jUtT51gQrc/YR54YQ2jbDS2Xf4X01a
ouFmlPL8iIgTwUlDDgTaAE6MGBEnzJHr+iTEodDbYUc3Sm8PJY0TXJSyBmLXa7Wf
IkRSBz88es80jbrUirkNNZcumlcmdj4xERfAw01bghSKxCASdncPpX+IesFEY/Hu
emLMVRdc3CzWmFXUitJ4nvQIXbEdHxO9kzl2tg0ykZA51emCocn1h2cfwNtdwhFD
ziJHuNYHHl3Zsu5RPGYEfHzb225ynsNkTV5Mo9bMeb6bwwSd0jQtwdqoz07Q+U5b
zfXOJNJklEbWzDDYpfSfQ2h7lUP4zENHtsZm0J7b9rOhIONF2YqtlJVMbLVRDGjt
oYykMRk6qnJP1b+2XJCMv18DntdWITP+qG39aQ3FG1zDBRufb+m6BG1uTabZNm8F
3ByBUPe5kuo94Nwx919PS2kTmxJscC8vte14lAlPVQhB/qlBDjROGdQGnRXs2Xoo
2KyFq1ml4GZVPPFcSnBZOISLWwKk+koGLd4xzTX7ppLaZY/6LIj40756evRbCbZ/
Qlaw2FkdrwheARkbgarLCfPF1nST/uE4oUg3Z5qWy1Y5cutdSJ3fxqAqoGS9+Xbb
/bhXTQj3vkdb6KPR2uzW77v0o8OWiecnCRInVwtam7bz5n7FOctiABxHD3sKSTLz
RQTOlOW/aP+1fRTlDMgQCTRnklXsQepUU3544F7TQggfPf7Io57JhOs/LAkSC5OY
ItXLt5OLvl0CKkVM4k4fFPda8ciHLOJ4g9qghwGOxxtxTtEiZH9VJc5wTFel0MUZ
n1j6o+WE7+zMiJ/feiCqmSz0Y/tRCctL0ac1G0lFvoX+sj3wHzWMHxvw8u6or3W5
mGQbP7Z5+SsoOygKra6Dyx41DdKXtduKVgAdj0Lik1UViQj/pbC2IqG5p70v3spE
AeLCPWnncoWhL2BM4m339Nhhpojw+ziJKJHKcfwmHY0DwgmiCE5Zv5FjAkqTbjfS
0fiVITqbvT5juRjhfvUXSfr1bjEf/9Jxt1o7PT/YojQCZGCISEJ37ps7s8opqvT2
kN0gXZG4eeHb7Dm7comIdrbTHJR9JjIxo87fUM8SmgvrM+0xy8iw2fP4K/bRCVQz
PyIcz04EAnj3LGtqaZTmWZo5hvV688yy3+fS5jmJe7/R2zaGs8Yjjma6ATFivs1F
rbHc9FnkwFrvIi8QN/L4ulEIue3AiwIH6o/0La3Lcj3LjbaNLp1B2zc0QWhzCC2e
98Mv7CuOfQrubnXMFTGaxbq4dZIbKFBZ/y5QGppiqXQFv+vwYFX/oEd1ibnZaKvM
atlybW4PVoaeuXktYvmlmsMNjXTzlMciQ5xotHXogNFZDXpsZiQpVHqUr+92a+tk
EDrqBNUujY+uxi3ilR+SGJTWWmKkEyp6jSQBiPjAu4J6uUjjgZd/0apEeHk66Y+d
H8LsG1M7AeaXu0MZ5ZSJDn94IKezk/qSJ073EDZnwxi3rYARjeIgXTvk3SWOsqMz
JfbnzK0YMuHDHof8y3ds3c0kYv3A44v7ruFkoldAzwqEVDX0xhaXOpS5QFpg0IAZ
reZoh7uVsBuFW62pNmkqqPLXHI+7LFJ335eABZJm7cSXypnhK7uigdC1uFOGDxdz
uZpCvGSj7sXljxyP1pxUHv9Z+XyoyPY4KUH0WUsU3x5GmgeICMlUEzbiiNU9fJhk
Zx3lcIKgasDXbActTvSkaJI8ff6y0KulR+dDq+p2Zc3jc61h3+5Siv1tFna+Cm9S
jT831G5FLyOZq4hCkGGYzFWm3xU8ur9lYzCjB0reUpx4r6yQZPgecTDL4CQsh2XT
i7Tc8+y+A+3gSD3q8QGPgMt/7XF7mZ2iNlZoN5nFGRKFQ582ePhDmyRYpEb2PJ4Z
kN9vAFOFdGGID9LyboKW275H/eAj7tSZvpDAH/3NY5ixAkI08GxE6NflxPBey01o
lTBA7XL6Wzf6VejfOS4czMRPR4MuuyApY+ckorhzv3cGHoY/n/gZDuMBydxrMBXd
s/tK3dzUPPf2J5uUgjO1RtkarbOG3e56T3VGCGPcNRs/pF8/J6S0o3evcxgsi2CK
AIAsBeVTT1VBGPpFv22rqq/cbiDkweApkFDhRE83Iw/T2zR2sN8O+rKlEaCN02b/
v7kjTG7xjb82ta2PfFHumssnx4ea0w/oLx2o4VXoI7MXvZInPCJjbXgVckKau3NZ
SOzwFnH/vv5XOp/sF+N1Kw==
`protect END_PROTECTED
