`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jsD5T/BAA2CssI8M3deQtWUxXF5sJxF3h3HRlkn6lnBh56dSAUFfAGgwBAOwgn8I
5vvu2K9VVeCFFvDbLlObn51ru/IQtp9afArvwQc17BxIOgvZj7FtLdrFt0ve4jhj
QaFstMuxBhSkFIpDfgE48+MdvGWVLW8HBmTdg1+RPP0dTy2k6Qyu7gmIxLnpEXh9
chyAK/iC89j1qyLLmQmzN5ZPxWckCpm2G/OdacLXlr7Ze3jHQRH4+mA4kKeL8TcZ
PGbE5MsIjjhGyy1HZFpjYHB3ys4fX7K9dtO52xG82aS7BdBJP4lh2eJaXBFDx29J
S2oZAFMYApc5+S3lak3ITzm6do3h6EdUpguomulcNL818sYFYeFRJofJNRYKUvDk
Z42sOG57drKQv05+o6tAKxidFpDeGG2P3NXNjMixA8Zrcr2tcgS/iYkl/mYZ+Vn+
dKIedbPat2Edt0lqBSixQ5ABfvqOrjkYOnHkJObA3CkBJL+mOFGSdpOnRZ5Pm1GI
Bu2n46eHlMrrLQGklKGWt+vdd+eHGk5C04g35FaKrzaBqS5bbU4bdmn3spWB1DDe
gkHKKivPGWIrhLpVQbSmVIZPuJmo7bTj0lxpjj2snNVmNdtt8H4KivrM2V5gSoUu
4QycSHsaLrfVABe1KhVV+MibCxoy4obQAarkRxJNmSYEB93dX4Z520ryN9gcTiXf
CA128AfRy58iWr/w8/yPIe4ZVYiUBN3ISHjblsSB193aTAWxai18aHZpCMGJdImV
9Yt58iKsQZAge4Lr9DjSAxdhc+wZ1RHP9gSDWp+hFiVVJKy0oFu+Q0LxzvwNoank
V3VQw2GHg4TK9CgzAqqR2XiSGm61aDHPh9nHXVT+kCjLY2oPT1TgZBtCmM4D1oxL
p2ybAhztrcGk7JkLnfI7JhliUqdV42z6TG/rE8I8m2N3Onz5yjOzemNoK7T5Gl8c
mPuJgkerlz7vzZCzr5syqZBjUZxCjydHu3M75TI3FJVyAleYtisxaN4cB/oDzlSJ
8PN+6O23U+oxdZxo3EO6PhbkQOhtBZsXMDH8yCMk3GZ396PAuZzgfIxQrKZTAge5
UY1Hf1mmVgKT7XVMpoW/hvVprP4DUhUj4G3AvLNEXwToKlH9cU9bCglb++EfGvvz
xMaALN4T0wbqg58ytOKI8oIT578On3Pg+eaD2Lrifn6ZijV1VLo7AmRDM1qF2FAr
hCwDUNojQCpy+T7v9YbFg9ywKlK+oyeoYEYRxtbGJhg=
`protect END_PROTECTED
