`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sG3gNMu8W+pA/IN/ZurvyaQxmk0A7OoE21MaDaXw0rssZ6GF0acIUZVZXVL1+phe
FVwQpNKvOC/1ayQRF96FXfl4wfbbI4O6o32/0IWw3JJdU66cH2E/7IycemGphCIN
ItERkvDslLPA+yjbXxD5IKILd8k4p+aXDUD8ykZqIXY5lOJp8JQODKMJISvGHlBv
cSR31tF54VgkjFajvMhLDHrPwcg9KXG/I25qFtkCGRbluKmg4Qx1MC1WY/dKsbxU
wwMrEGey7/3XHXb55JpBTycQSLew+MzO/d/2xasonSJaiNGXBFOONVaueOThNgEL
cF3LG9f1BNbXKV5eXpkKz+cgYbnO3AhLq6tf/BWqLViwUKwz1GHF0d6AWscuaXSM
goqaHymmeJGYVrCjIR95Ak+oR8R4u+Xhcu1S+U33e/tilDaJdkV52WtzUthDx9HP
Juxnh18tyGI8rGMQXfpl1VU69slqLhmpCp4PrMrMvM4MSKAtTm/9KywbyU/zwV6p
1B8jj1mn8/fb1IltZFSZrMlIPnY8BcEVVSrZiAim9EdADyjjm6VS5p2BjDvyld96
AnpdpjEgz+7n4YZvO3b3d6MPvxptKdpdvAcr0GAmTOyph7pUg5Ru4qjIrxUKAQOl
KFyXIhRYYbQibolNx1AkM4PWs3SH4M40xlO/2F+YyzcWOeHU1ccqhnAF/G5+1TVs
O9Jcb1de+iHBn9CqmignLnVMrMKRAnwwA+LMe0nAST7ZwNZ2+JKI4CLtkQRT2xeD
OqD7NHCfLKMEgHlmApslF7snEb74Hp7F55eb+2jXfsLOZf4C8+K04sOhDjrTY3Uk
7YPSAkxdmTsQeoU4GxmvHE++/J0KwBdS7ETneOs9J/xySMDZSx3Mx77d8SbCOW5p
cM2lrpTYxXUQhCjMQmUVFH2kfI2Rsgou+dYKOSJOkv6YxXVABQnWUPeMfOZ4KDpY
t2lnlQhIUWqK3Lpgz978uwLS5DJF+jAIDphZdcN85ndzSy9e8eils+Dofpk+siac
7hWTYvBNyfDKy3tng6IvH/uSoPQuo9OLXizOBxACe98ZZzuRsavIDnUTcx7PmP7P
q3386AhtWQ+fRTo9AlcKS1Zypa9LflPFo8vMYaZlJHJzOzTelS4DwIiNkLZ4qyvn
cyEAOy6Jke6qH9QOvLO3X7aWJ8PCE1JnNBL+BD2weuDJ6NfoYdCYgSjucx/F8x9J
pv1MV80x3djeiAv2WJrqsptlyMHkrOI4OiiBQqnnjgDpiaoS3wFSDMakKU78fsB+
nEyeuRErlnyqvShJpI66gPqBIFv3QGus0DDhEQmL2Ef0aYKarCDqRYc3A3yLrP8m
2j8AgII2wQBh9MIa7Gyy8kFgdz6xzL587J61GigmCe8Xgt1v5gqcKdaxH+vilZCB
9UkdE00iTfbEI8Luq4SQUrrUYFcjQzi7JmZFyze+XGrsY+0iWTi2WNVvnsvUhI4S
G3UAHUl9LB65/DRMzRvNa1SBlLj4SqPVC2qy8pqgpF/IOOrLRizkPoabD3QpgFdW
PehRafhLe1jxOfIjGdK7kMD/L6WPdCvAiBiTy4b5XRSHX0qW05MNkoP3E8muFGF7
IMpeZYsKweuSEGHh1HlXb9k52DzEda5FBWB4qxeZcJDrw+bi1k6yTV1JfD4LeBYh
zq8i+gpwD1EKJRWoak/jDZX4mwtPNMAW47INFkpkaWllu10fQK+T7BbwqmxNi/Rl
HC7KqDbZAVBQOVEf9FRXBsQgq3TRFzudpnua0M+H5RTILU3HpDJlIdP7Nu8RhwUf
Qn3VNXCIjAWa5lCG3Abyyy6vQhDKkuAH5PXVRUOqW4UcNJ/Ox6ib8vVA9a9nasku
3SmnWrg2rJsJ2AzBQaUVyWlV+5eFg5eQUik61Tf6w8sSf7w9XNV3mlg/KJGgbUN7
3m8OO659ZkLG9rJxfM8Md3Mvkr+6eD8qlucE9n00QoEz8rG8IPxfrUI1QXBTCt0Q
1q9EMIHzzKti9xQMT0wgZg5Qe4naFfpUsP79WR4VkSN+ACHxo8ObjfWAoUhLOiO2
pFSyPyjqwYTHsWdsqgvuTWkk+5ar6LgLwIXR+cWG/IMOqm8oaRGO34ScGbjmrfU4
rC+o9gEJr8HtgExraSpW8ZaCp9/kZ+X6qpbdvGXj5TeajDsyCJfmfbgdpS93juFC
SB9kJYbl8JlhHrXfhyV9iWWFprdSDdX+S86xvvrZNayloe4dbV9T8x3P6vAGHFPH
OZv+n9d8nLDvhF6NFpeL1EjKWM+aQ7d9qFU1EVLyaAU7/DzyZPI09OMNlio41VUk
/KEilA8/11eCyKsRlNFGsAfD8YWba+NkDbwXEHxI++VUbZCJmhtXVnwURZ+DvBUb
284ByBxVBUzvTp9gfCBsAe606jKli2t+A4bN+xTjlwsUepcSbARp0Ysi4kXCnraP
/1ksLdsXC5RcVlAUGq60n5RXmMmiGj6iKuCGxBFiFFf+oZGHRXkc2qYlGT+XSwuW
+zqzANE0l2di5eYORish1EKPYXVlWgmdWA3Csv2DZ4M=
`protect END_PROTECTED
