`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tFgEj7AINyUP/d6K15lF5NIMt1MAJdCluY5AOWwhP5kxpQJI0t7irvxcs8zcOQ/R
7GsypFQhChlQQlza3Lq5985YGL4Cbz8Ac7/LTkeF8Rt6ManIUkbGji1sa1AgF7TN
HZiwC6VrhWFrzi/KOqEFC2UBuyDZ80rGEpNHCsP0Ogu8YAAbR54q+kQlNVJ5O7fr
2K2+5G2ecbFSij/8UUtY8EjO30PEJ3yjsDUprRxOQ/9fH3Ea2eUCq9Y510FzL8LZ
sxFu2AqtxfVWYSTLx7xWJ3rcWHUo0hUu9vZA2lYxGBFpGaxNn8IsCwO8EJOoGBJ+
REMDk5bFFUWQFGrV3m4PI1ToLhtiE37RH3q47yfcwy97iYJmcjenc1YTXdOfS8eB
cSxDbo4C54/r4iAjWoeAiewHfbCVjWTwQHR26K+C/KO+BJgJiXyHeaxpQRfBShUc
aHIurdTJvvX4QUWX/sOnA7/VipItEkQCNE/B/McImND/YA0doskMHF+F8+AmBmqV
oSz2kOH+mRu5UaQTrRsSVws0iR88fUJ6QApEAlUzUvCBjgR4FVr/Ejl/Z1jJPCjM
vYGIMnkL4yvhWFpyqEQQF5yLPZOgWj6n1TfcOnZ7y3Gqs5ikvKYbPL+Xx+Neiz6g
kB8Z9TpUPASv0m1lTbwYrUzoWZvxC8CBsfjaRwi1jBWuAsOO640hqs+OzTxWizcq
pjtTNOrDrz3IYNA2duZdQ3Ouifi0cbPQbsUFTM5YRqrXk4tiX6eK0qHUardUyFVS
M5w57pwg+P94FhUBPmxusuAtUlZvmBlr9pEcjLshU56uWH6cmRn5paQ0akhVRolu
BjlKWrcrqUPzQq9IkM8Uyc7an57OvlbGCf3OKkzRIxKFlFlcop1d/qJJYCGoXZf1
qAHjL5eoDRTY6YBkwiqFMOe+NIaTEgj6FRX/7yy13+xqKH3h4kmI0EWm22oaOtp7
s0fWe5b3KHBAbfXScN0u9ohtPXD8cPpafHbUvI69IYgrjsWa0YSQcFyfpxG0kxAe
U/WfjN0/bLTbNP+/TfrxoqsQPXB5pJ85z2dG9TU4onVNEx6HuS8QokbPE6vCDgbD
lwbDheJHCSVvDIN2cEopgSpIgYt1IU3MHwe+85yUikHeEuJrZZl71gyNrtebZJTT
QmpAPJntOWz8iqH8nZPqTcM4JC16N0AOOlqUycAYK4ZfTJJgMjWH74eKbNLuJcUR
cwQKrcUdcnFyqSkZDz89thCktiI0oNqmmJlAoC9N+IYiYhlDNV5g7B27FnYotnAB
VWatQQ4QWc9tzifINnncQ3u/CZ5yuwR5IKSpa/AXZ67jSaexI4FXlQC9UeeJ8Txv
Giq2mM6AOXib7JTew0DY/kDZWar1ETX6MjpINFiTbaHLb3Jjbe74tBetDYtu7ORS
pRLiZjrmd/lpGhfJxE48s4kblLFh+Z4NJU/a8QHlS77oALoDHjUFuhfs8gY5QF3N
kjgHxKD0Rgs9cODTio0xpiP9jE50jAZmt/gFH3ck6rT8ShtuMgnEnQ3If41eCUVM
svMrtyuklG0UTHqpLIcVCW4s+FTgf208j3Y36h92+9WgrZYx78lIGF+Prsaol8NG
pehtrDDtgbOaCYEO60PPlcpf/PaYs/8LZIxIHSUmho0nwddmhqNlP3BTox8lhYZ5
Zrpmyjcxw6tJAHHhRE/sstlCtQ2qfQNOT7FZps/gS7blWmiK8Y39b16iskJ2zBtd
MKwVSNkJT8qmAvrqLNMAMEmpSGHx37JTrR8oD+GKJ158PEgHIRarbY2Zup/ZobDP
N+4J6rBq3yk49GRevD55kLW8vvpoAXVqJh6bLZ1AhMPdPlc/rT460ZqPTT24noc+
0+jpOWJPPtH9XCnrWydIveWjEHlYy53JyTB1SYsnGkCDKbnltS34Jm7LCaq0J4K6
ZjyhObsJDXYgEjIRaLfWSvCM/y5N1qS5mXbLd5+A5/F8akKH9MXm9YkvSx58Fgcj
Q3l5ofW/wORcSZFz2PCP0zT2inOeA8xT4sNpdvgARRafYd/UmusmYIaArLKtQjIE
Gi4vfqxF+GJUrNKHBM8GWH8kQzfPJ/RJ1aPdErZvxL1unHZ4A7S9kjVrJZWBElyP
oTs2SYC5LpYk+Pgjfw0Q57qhxEvbFiVILMvFSDfO5q3kbIvLrmsdOtRaEqUaC+Pw
DJ0AYkQJHwXni3OSVWNNF5atTZAqZONA3JX+N2DiaCkRHebyYL4d/ewiYZKVubq7
GvxuusIffimxmjN6Wk8ulIpMTo/jFtO/TlOuopjPA4i39eKu3aSyZpPBX0irkFrU
ozpT+rNEE4QUtHD0AI/RCcfFaJEWKr9WWZrcmkZ1kQpWKnyJdilhH6yNFtKcCe6A
hbsts011l6Ztc1S2QyaS/du9mObL8JeE2yBlDEcV1qlATlP4KMR68Rgd755/1wnN
VbV1FHiMTtd2X4QuA5/Q0fAIF5zjuXtFG8NKR84J7hWrvJXGqAv9amV9dvEBSThY
N2gdvgfK+0EhQc5yxWYtkWClNPCmG0QTk9DADTlWsX5txDyKtkk0lsV5/DjNSUUk
tOpkzo7ebQWo/VS60DscFAjIzG4AuNZ1j2WW4rLvygYNKDHLEIwTNsdK+PiSnBxD
v/OuiQBBfo7Zaa6GJ60DYiD+kqtOR9p6/VekQ4tH5OZhnL2vuiw06/FdyuA6tZe2
m+Hd4Ar3GFKeCOTauDlt+BvyYsM35cE3F0SZgyqduaiaBf6uO016hGL2yH6QR+cC
BpGnDbiX/15OIWs1rHkJeAwRVW0T7pb5+9lG96v7JNFQRFCHtxmxLAY4yrUIF4TK
wLeun9RaGMy6+Hu+cBdTgrh+1bbYsabZFTB5RZ3b/Xi2dcuSoMn2IAJJ1WB4LRyR
DW7LKzraODrGGSbUJTL0Y6mWf8nIsEZWsv1NnXFuFxiUImXTZMKptqpf2ZuJry9+
grO4aMIessRHZkIO0Vhe+578yo6gxlnz/rgBVpZ3O9XW39TADH5lPJXJAKkkn6ZV
D4+L5tLwudp3NLxFHWAGEPpx05QrJuopIe5idmJEoWRbVwoYE9x+9X07pzhonDs2
hKVqvTIjrT0NtghipQE57LSgOvQfVrh3tcSfKnZQCA6y7u9BdDzPiYAFI8bftXtC
45p5cC4ei2oJGJirG1kuzOrBOFhmdvjXBShm3bj3MLtsGtw9eBqcU0X6tZ75NyXG
5d6413Tw+u79BhArP3ETM/d73XN/2ftOa/UKOs9gYMj/ft1eXs8maHy//NqE7B9U
Z5G0Xt8X79C0km0IN5B2R1qVymLWgW9Bdib3TNYnOM3+ofJvAIDY2iaJbtglsK2v
xCYJ82fdLfWq6Pdlrjca2XIDd26MIWPbw2ha8tqka6zLaJWE8kqWSNztTAvaGLQf
4HEH6gvX7k4RFjFePo9JIsI/Y1lmaaRMoFNqm8dMS+kiGbHtSD64xtZXB+cF2ACy
T305+tpNszqI1qg7laAmsrzvprY4Q+39fncaJuOANGddeTdeqz6XfKpMXVSftfCG
mINJQilPY2A3BdAr06ctbjkFfPea65KVklDsgc3QxWp4M4HJqeGlhfU/RHSLT6wi
9d5+R8d80Xo1mOpmORnb/oezsBazHU142FAiBysFMOtQRN4A2J2gPbUC0UbLKpzM
+u3/XPFqFNvcxt+iThCsCcbsI0PJIjw6TZCULguFR3xx2huwruxbsJSm8iS972ai
booWGdoTOtT1vNkD4aj16u+aJqVpIN8Q3D6bQmfOKe0cadDTNk27v7WT6ZycGvYS
ojKkyXSGd3VUQp8Q4CALiZL71aNCE4eGDWkbx2R55e0Q8bgUfAgpvtGel33uF5xl
t6eSznls1S5BOkMmXtf2gzHuAwvHa7IbWO3KYMATJkl/pwBLos7kl5auoSAy1q/k
dtycfaL5Uf6tXRk9h70ab9JvcwP5fiHvi+R7FI3vnzgk2ofgyCi/pcWV305p/lz9
vBTdApW7Mu0FHGfCS+8KlWWrFM7IlCAk6lv9G4bcgfU=
`protect END_PROTECTED
