`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UkIRfgPob3ULpjLvbqwB2cYbOqB5Mg32SCAOKU5mJ90zgjZRhZn+nVpB+YiwWwJt
kyS8gGB3/317VZHlZK5lNibmDXN8KoXIIXCjG86I1kOnn5juEuyZBbwyE/Suk5BM
0BRKwsvmaAFqsSKU8vpaMRKZvlgnVCTiGFIckUahTORF70XdcWtWkYIpCVIdL0ov
tp0wcPV1agxMASRffDPI/MZAwBwstCi3sm4T4u38CIMqKHukySoyGqXYEw15kXVA
Hamn2WlNvAFtRY8pJzLO4PxTiNuhQsIBIR2EmifEqxZvTi9YCok00EEN97gndY9y
YkXQdnQJaR+eaRqZF02MTX9OjSM7d6sWS+3OkJzpr/i87DOpTbmMJg63Mc2LLsr2
IgUOI8mjFJNP5rulGatBpI5YbchBhe2C8cO+tNGZbBMFmNSkk1DMIIqOduKdOGsJ
Fo7+3YPhhmse3/cND/v99l6gOerUDcJXXZNVW8VHiJJmqawhjrBnUvw5mZobLBz8
dC+wm+CvaE69LmUgCtMYMZPF+VuyYm0Qk9I6SUYjsIBPZs8iYZes9qtSW0BQt9W8
LVs2y5PSz5iSEweILKeTpb3sGpT622p2HoMZCWOxtGit2KWZBbunJNMRrYdsCd3Y
3x+utSiizMO3C4bMhUhjARvKq2EzgOGHmmVklOs5qiKJX5+qqd14ZxodKtQRvNcO
MAr1adHijbAP0IyOIhcqNY8ozUBdLbSwOAjPfZ0M4+6mcA+wKS1wuBazd+/722pD
MIbJgPap5J5pbebLyFHFJ1fNjIINgR7f8Njkq2p6vuyTh5LMRJugDC+fuNtb09qU
joU0dRCp4mi2sRRETw5GTFirIGKUHkMh0fZSPuqd5gCNA8A3CB0JlVG6obk0wVgK
UNc88uO2yd52342B3SI93WYg/suFwUkA8hedMoCLrW1mXbEIllNPRf7MzqbY22gx
vbNSnCwJGacKbXmwqQFSQfoSh25oZnup212SqDNDkpxDenmzTLv5vzgVSvJwv6MX
petqSoflIEOiZRtkq6Es2yFQwEsQur3A3i2sZU+vbVGnYFpl7UWisWIllN+ydJTG
Ysdu7AVoexWhDJ2Ypv9o9Y4wsBuagUW/twdxhciw+0aQi8LaM9lOl5FfU8fd+PuQ
jEFi9lwZ/b8eayH52KPx+7FUJqDpwNIN+Wgcod2l5haF46lPvwAcdB2srEjbyTDO
uDETHnYQanzqlx6mkgxMWV9sOiZXrVFbqQCc2Y6jXSUatB7Uzgu1+PHAPu2U/phy
6SBdc9u5ejiczOd01jKz9j5u1ljsrlGlce2kAwCUgFqYX/5MSaRYyoEo0/p9rGx4
6+x6cLPU8MtzzLL/FNWPZSD0n198Xxa1EG82Vtk4AHYE7ek90mG049m9YXS3fpfO
eDfAG3jMhZjsDb2rX5wiVW/dC05vMiQMWgk/lCDakkGRQNzuq7UKSMDrl/ovIXZd
sQT/wp76FJIyfAlaj+PE03T9o7sJTcOoR3swvs0Z/wFn47z2RF5iXF/Rk+wLYS9R
ONtPxkI/Td4pm3CYdnBhaknca3fENri/pM0sYWIHjMmP1x2MWqX4rFtUlDiXPaZA
6ukbEkRTdzpxE3MVMjistjL2Xu0msiggFCuHGn4TbvaEwNZ6V3gAfW3dZ4iW+yno
a+1CybrGeBg6BoYfvHkVVCpEQw7/ka0x4sSX7sUZel2tCrs7X8PNMqDbZsoPFfie
rhmxsLskTrBfQV1xpAt8A+UpwYp5r4tXACl82u9esmyAm3MShUYI2TR5wKU+qQNL
Eu0LbbCoB/tj5UmETR77Ei8yPDVQSPi4IUVz2+V5NxjN0Zjrh+x0a8xhxgUmYINt
Z+1xNDYK56Akvl6SVDaJ1qrPc5BSKD0QZP0yM2r1NWbE1E5smUvu0dz8pjbIMoHr
PH5+saVqY6EgQCyvi6gw5nkCZDgxEiDeV0zNgzzCg9kjAPkSLJ3FFEHA/PfUCwAc
YqdAWlsfoH0wtqYhnXLGWFqzb8MbE7Uaxlj55dQgofU8IQs5ykMX9XMXAhDv4Uz4
bLdGFBL65SRJ6FpbZyVAoOltRR/9Ziag6d5wywWMl4A/GLkkIXJQ0XBJGMmqou8x
kAWMGbf0Wm3UaEJuHDcfLku6hofRGVPgLANCL3SfNaBLlhC3VpXqgDVSbZV9Jw87
ePymxHIO/bqAqn/1iK5QgTqwqxAZwVLxiWfq+jbYVRIymcT6LQbuQ7piKtezfg4W
QVZAH1Oxp4l0K7b/U4Kc76jtl9Uw+5VdYEhnVTJFSEhz+El9pYm55NB58BkkTqxY
CjS6MILjT+Y311l62zWth0GosG23RJ7KY6K3OaHhPGMH1xccIGnEd5FSuxKKeCYt
6OA2tJmsOKbVhBceLjjMN4T69wLvDy+eIbJ2UWr9eLiV6SWv2k4UxSE61tZqXgAo
Ef61MKc028YBct2O3/V8NNLNNaXvAxkL+wqPqJmPtxRsLs73r4gJTO0v9g/3M88b
bauOsrdR8nNmZ9WuTxxE8X3USe9IbEbzstJSjwOgWAXv5wKGguuzNWuucID6pfHy
PmtxpvB4UiK2O4TmUVyVSrdTCDkwtso7udKyT9N1opWOiCw9cyBClTSfEsFFJOy6
gwTehcfUUGLtfg5Icd5d8f8I5NR9nBwT8zJnMAABzNmrwZ+K38qHYYu+QM9kmJRs
QGz7kYs5Euej/+9wNdvr+YJB2cVewtjSn+DvCfZuhyM2MIM7p4QLp6D07rDS6jzT
X5bKRi8LYIuFxAgmzLH063YofkEUxtk8oD6SOHa/rpWw4XV3Wy3fBrVTtMK3tSSU
WuOnuZ/laDWUXLHPhjejDepvUqASgPoRz7QPBxllJ1ZyxkBLEm7E1DsNa491ryWY
B6fNwyqmnipelrL8Usqk8HLM2G3tD/Eyx/R4BEiOv77pGALqPGovcgND8WlLFm/R
3TZ6aRn8f5p9lxUW6uLhB9xv9qHJL9zJJF5UtjufBOdB6E9n0f3AJuUMF4pM8Guk
SQwYc8EqxTkov9Q8eHTiAu2mZ9biLkPZ5k0snYA8bT44gLt8rJihkJ2q+8LBdW8h
w/N+2taBR2byp6n9J8qSNtbSfjM9hvUmYLu9FFni/9Mx04uocfg29qcYh0MtJ/1j
vASNh7r2HLIFuPiuflqR0K2whXtpctqz0sZjCE91P9LOkRYO0ITtYAymEVD3I+p+
pR6dc2B6pjEPTJg5rcpaSymvi8m+lHPYoWI7WmuANfPufumqlHyxPWJ1x6QjOB+E
8JdvKexx7z0wQAn2nXd8+g==
`protect END_PROTECTED
