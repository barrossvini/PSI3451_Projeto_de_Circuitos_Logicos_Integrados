`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2sQzfxC9uttgK85qhlaoj47wN+QrSv1zKAiOK/SYbSLMOC1lbdjS19V4TQsK7gaj
rItKwGpvQdyi75fjbfzYLC3FsBKE1hdRsdp+XojuppqbY4OEdun8AJfXeFGmVVW/
VnpaEYn0izXOTHQBvGEH+TkiZAdXIM1aSM6evkOi8tFE2UE3lO7zaFv+K+zJW5Cc
2shmLFT2m8H0tuOmzEYll53GRA01+X5UgBmqWA+oHHIklfgy0G1ephZfgJNrvPZ3
f1hEqB988JRBLYrN2ZcioLF3l50N50H5cPWekBifps2vhG2vOpcolJiN7WzIqkwx
ZZQP8mKa1/ie3ttI6w3mWg==
`protect END_PROTECTED
