`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rvdvTMtSB89xSOgj1BY2IiRwlt0EBqFooBoMDa9h60+BRE4MP/lM4Ut/0XnQmW5y
t+FCXRrvOeKO099Nr1OdAvQUCU4+BaA7rw4/mbp8o2kGQBMAsARv5Ji/8yOzUz8E
p+KhEx26iy+7ITxWAUAQ2p4LHDDcacZPZcjA9iglpE5XRAjtul6ouLXxKQPVyeRX
1Z6QtRujVXTeRypf5WBF23eHxBa72nFdiW4HUWGfGtChHhh29BwnfuHpd2+lKjvt
CidH8JJ/9dFjvd4pb2oC5D7BT7pRJzVhSMXvbcB/DyAda+8gq4Mi/ZCRMygjBXhP
LAcvtrCspT3x+cTDc2wiO06jJIq6SMjSy4yZIgjvqcJ7N6ACfuq4F2J3uh8Gu7GT
ocbKLR7vTzAyMo5b4hgeCzr0Nmo1B2aM2Zjr1Lwk+mxQpRbEyE4GvBIM35oM3GiT
ZyKDbRvyQ6XUZ/Haq7+m/d/wTblYhUV8OqC7t5MjO1TEMyOqXmyPDwKunwS4FXcw
0ubZ89AX/4D1IebG5v1KdBBZwnUGB2P6UgNVsJ9PPxhpNhsHU+ZkAbBTlunUVsXG
Jsvt9/YVphRzfgXvQfdZHgUEW5spt498VnAvG1qxH/bbhcDeWumlaAXNLvNxp7c6
kTCyAqP9318gNbzwcPrmFoT1dxR+RfZRmVOaje+XNM740eiOFd5qIbAnAGU7e5qT
Af+cPbTcraFvcZmxT99zSpUD253Cp4znZfCJ30IVcREGkTvkopn80VIj6oOoBxfQ
N4apgulbGibc70pVwXl7wfBYto33FETKOcyE1TtYg8YGhXWNZ+/3zCA2az9g+ord
AivtU8uq50Kdkhvun9OyFZmjRaTzM5huQNrrTSDEcxvMu3mdfZ4af1w6v/zWzG2s
Tl0BCPJyc5RaG7VRa4fLMTVQZf19Bc9wmbDsSC/vguR5nokKFN20pw0KC4yzwGox
vlTIWnApx3S5exlVLs4DUqxrHQBQeYc6HiB/uVAPXYoASaL7vbaJzmHIL09VMmVG
wCqOzQBftYkWSlNg/ZmiCDzEh6woPP00W2J9oHENoy+Iby0nM99dzA4VAf0ygQ7D
uf/3cEtEQOH2HRPj/DRhVfllCzi36LwCVsYWXb4X/uyB8c1QgqVcg9Lo7//5mBCP
nJGZ2Afbab1dEnM6oxZ1kQ==
`protect END_PROTECTED
