`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6nrg68SX8gZ43i3Eo5Ibe4OVHRVTxe0zVTN7WtfqnQdYE87yzCOgYKeQuylrs8CI
9II5UoVJbtfuShdbFDBI+ZSrXoy0qqf/INnHkpc819I/8v3mtijmNNY+egAgexmD
fHq6REnMftw9NsxyKEn7x+3Ru3htsKIpMiqT+NCZLUMYprCore74xcdHZ7oNVv45
SUyIdsj8iQ20LzP5CmUSlnK3FN+PV2SbohzF5F8UbMaC4EYV6Ex8zXzsDcemndcA
ZbouZmna+xhB/yI0KfXZ1/EiHHadRmAPgep9rtfjM4F9XqCXkufjMY/MrZx1YI6S
KluNZth148LJ7RuCQ/Kikk28BF5MYxXSxe752ag3VNj3c/80E7jC89KJlDxWpN5K
/m4jl2VVZhbFfGxixY7tjbeSa7sMqLoU7cFv4BOdeWaaKnYUIlBZyV4zozUdLPKb
aUdSyXoGencrs9HdyHufv5YVQSdzTxG72520a3CfJoMVExRlfwNu95d21NxL0GRY
hZHPmQGhrV1dKY7ODsQBKYxIRx7k3o6oWd2yqlaVY3+Phu52iktK6j4icbpUhSZZ
2CLHAdWolcv2rGKGTQ95KH0CLJuUg50uenUgbIrYJeXknnx4/uFjOxJccDViGe78
WvJbOs3K2Kkw6vyWTtMsInXJvC7tbeQlUhisUcOuY0zc9xY4IZsobGeXxVhoDlHn
IMMBiNraruKQ+R/PoZDPEE7PZ6LmK/hs/pRamJM25LB1Q4aVvumJPbsxB6BP5N6q
1k/+MworAT/ioLlbuINWMC2DZUvm63rWsZce1VCBWfy9gJNbKARTpkqMuHx5dSC3
VnjLnd2TDUpEkWOpBo0F2G07AfBXarcuo6iyyS9pEM6GxttYMYadUwLaBzyEwsiT
gQa+ledmmIaBStoaJHUVydIYaZdThAOwWyjy846els+5SS1Bsi5RiC0EGlnItE+6
y7SEpV2rkzwWe9AnzFd6mgIpQt4tHwo6EHDjlaPmFIBuhnBxnbnMJN+xg8HAivrF
l/X7bfhSaJpcNRmxH0xq1g0p8iqvmAmeLEoso8hfDMDoRGZJnCI9h+KZqSK4fPuc
v7kYywjhsGVspZcqUE92Nu/TZdS7BPfY0npI2IKj+YY8opk3+6yo0ydkltVWSaHV
f98tQDEdEvbe8hcTDVnS3N0plId9ecKzRUtjAYI4POoQQA0bXXUlwCEIC99QGfrl
Ufjp+/zaUHgZk1Cw5NvrXuN7YYwjZCcEtzpmKK1aaMX8N3ndpMIJ1K5O+3n1jCLp
`protect END_PROTECTED
