`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LclgrLPVP6gzfabaGVXIJFEFqFi2Jbib9ep52EV2E9iiH0g4UgigOlqoXi9Gjh+q
yEt9FEnY9E7iFWhV/naQdaVDdi/Q36Sc9//pdYvcOU21rCRCVKfescycLnOmP6Jn
ruH76hxzQCMV4IwolMjtM3h05ImZxXROQJqoqhgpEkW/0M5Kl67ZZm5RmliKCF3l
7Mr+LNJnV1sybyVJOwQx12HMX8UT4PLHfQu3ja4czg6KeHd9G027FE6qYJGVrJV8
uWhm3EuuX5rh7UIro0rO4NP6X1kcOyN9rOAqpvI8+Rp2C0DrcjSC4xVAnipz39VX
0fcb7UNcRGnppacG0iOO8bITOm/ZzjkrhW1NWNSGokEvYMf6FcFw6UypHq71jKJt
yUXdT/4fX4sC+xchYk/v2HGX1O/2eMHGSSVB4OcDAhPl5MMt7oQ3UblypslbGaje
L9OUdrNTivkAe4RAqKSCpLzAJ8MYDEEBf1PFhmNtuBXob8grv1LFSo+CcUtx78pC
qdVj8TxXID2EF7YjgNHujErJYiwaAjoTg1rAl4SgUO+rUH9tUaLNeufiKuxKoGbO
b+1BHmb3LSDQoUoy17q6HT3VU9lkY0TGXfQnj3yR1u2sqA3xejiFQKkJtAQoUVqJ
5TYt2EPCTHDLzpsqY0n1xV0YrwuExuI62SL3xXHlLbYzFf62bgxsc79lfcy+s8sG
aBWSGdvSyp/bKpMI+93SZeXqbsICeYJo63CPWXNAM647opQhAvHZvgi7Kvq6ISii
vIQSXBsML5dbr4P3JEnbtr+CaMdnMYCq1jV21Hu2ZpX99pR1M7KSQjgzGV0Grxwp
3MbHEvaRlG54n31bJZy1Jok1z1wY+eD+9SNP5xJl0dMWygOCwGngQKl0P49y0tfR
5RNclHobrfZsWtIbKkgBE7LJkhptjGHw5cK6/9FbxiUzD5Oja/1noHoMp4PxgGQu
OFKl5cR6EqrA+TvjgRO96opJ6AjuvpesSXLaqMPWERrKn5zgVXR34MpYWK0wUeVY
FzGGi4PSKThAtHEHOaYrX56wcuqZW19vjMegc1cuTHV0X3iEQPNNw2sNVoZxx7YK
nKUZyWEVZ8ReJOH0BW//BmhwWLAx9/IdI5ZEt9KXe7sPgheCEEoGNy978SAH8xfh
vsOPEAdtRER/6ovmYmcPmynqOcFTmdGkB+GDqlxoRF1pxAhAx14qPIbz+gL0scM/
DxgXhcN6oqx0tl27uKfZdSw3Vd7KgMNG2PYdNWuBfpef2MSRHqIOQA2p+CZLDwtv
+TcQSEGLz7cTXcg+4MA+iRkS5+QdnCPfUcZBDMOGvmWtYqsWcJrQOtYG0Ms4ON4H
FteMLbDooKQEOLkiNn8YaufZzRznnKVM0+TeNAi8S73+NteAe/nEqhzk5/VkNb99
qVA2NirQ3uQGoqtI4epJSNP03jirMpvc/UXyVvFq6dpjr0V1NuM0P3GO4vmyCIj5
k+ZtRRoViuCeyd7S8zTHTMAXpEXr4ZVhZwTM4WY9IcK01nExDURCCjd/kZ98p488
jVnD6YLI1xThBLM4h5jelRISbh23eC9udqxygunsnyJD4nXAG+E6XF0HMxU2ss/z
fL1bgEoXtV/SI4T0tnOMHpa0ul+mo/+70LzTptjsF3yh+BjLk1+Nm/1Mm7qkyjas
0qmAJoCSohbaCqZherhNoqvR6mUrGfHUhYAC9Lve1x+nyQHzNnCMmS0qpKrrL4tY
2Nx0f/apELIt1sjgM5B6kl4uZhvvzJ4Wt9/VCc5q8Y9aPcc38SqqpWAI4JEpOnlg
Ti0TcN38y07b2ho1htGKvRwrg4L1OJn6shwFVS786D4FhWxTe5Jgvn5dT7ViYAe4
riG1wBGkHY19fXZ90Yj7L28xpAtjbHuezUdmi10s5gnd/JypXHgE3ePpJjzxE8Wk
72XJPmu2d2u9R/WeBz5fTWCWyaFqArK8YVODhDjtQa0xmkkGCwyTQI+TFyVb4NmK
WzT2DJdXJfYOLZnBXkmDwY2FNmeGv0PAESc+nNq+cCdLlfOJg1oaPIBhv0InuCuM
EEDz70vNx4h+eHJhaNy9YdFKYiEFubP/HyE92H+CED2bbo0IcUQZ+0MAUygiDpO8
qsyuxGI4LNqnIebcdot/+P3sX8KNiAIGl4CkJ9hh+LBu6/uDk+zCspvfgxbmDCQY
yUxBjBXEibz2XdCADIYokLcodPmNmJ8oRBi3Oj2JeNWKsXWDaQWRI2jYY++seMZb
VC0HCQM1TAedKd0jHdLGaUFnzElX+YY6ZWpuhBgj01w/p5n5iLg9A+AgR8sthbKD
Orfdl/9V0xl53d+1fu2wHWv7vNky3U77TD7a7VnnGIG2cAKJX4kMwLVVrCfWIvxA
6WTkLvVSRxyPMLD8ITEb2QEhFUP/8hKJZdZtqpcQCoWbYaYKOIMwPVdXveZX9ZoO
+TOJzFf4QGuLsaqxmB2rs7aJjk51WXnmjZm62cizkDuQmoAK9Ju90H/kPAsfUahM
ZKpnLzg0me1hvFG30JbNJN6hejmh+hvxzk4y4Qq1G2joO6uSr4R5k5bCiK+2+rNC
TmS9INSWaWHXcQt7b+0sdI7lJvyYvb4mpoGF70w/bnfguRM0it+KUzwIUME/SGz9
nliLUt+QUFjp/TedSYrQ8GiZNea4JcIYE1Fuv/4Fce/k2kdJUyuaUtnhp8tB2O97
14pAatXm+9PDBBU0F8Klfwarmgl2UQ0ByJKMJuqDcLSFnnWhPN+6AsfnRuAyK8ac
FZ3geFumXHKp/q2cXuaZkASY0+GvFLSgNyIwaPDukMNyWtfNqIh/nnKBNjt3hD5H
5eKK8JiDOZnbdC5+qqAywNst3rDxlzvuNOGS1b/rrOh5SyD+mOLPTnasNrWUe+F9
jY7MuwjZ844uwrpCiwJAE1GSgOPW+v/4SDcV9clrjXq4S4rXddvI4pyUsx7yetdu
O2vhwpfJFCJVESXFsXAjEKgl5w5mUV9SavH5GPpoXV4ybX4iFR+LgFS05oBGWBNg
4X1hndGStRb3swwCJEsS5hR4hqaLSdx7jFzq29OJYbAAu02QCfGDASKfpU1Noz36
OLTvq9M8s1ze/3XT3LkKbUgeaw7L+e6kXb+H2iiBZFSU91vgmMu2qOOS6Jwr3ZW1
lOF2P+7SDS89/OLuKpgL5Hwn46gpC0dwdraxF0q0IQvgVwbqMwn5V3xaGbFVW+Rt
OMWuV0F1sd/z2k1MExLpYR2c2h682sDdmRgYF4zYR2Ux7AY+F9wv/0J5+cV06ZPI
v85iD4Yc4uc5lmCc5a6VZsI4Enp0cZ33AO1r6rWujU0hrw01UGlJPnHgCI3E5WE5
saentgg86X+Mxh16CEBxECOGp92vRp37kmoMuYcXcmsqDlmv3KBae/CRgKicv9+T
OZmREv0j3vEDEXflxz8XBaBuDNDAYWE9z1dbojbxF9bPAlF4bAAt1V9tu9UwJIH3
9oh3ExRVNGMF4wJpAmTWFhzbCKYjfHIoR5F2ABQ/3YT3NoSNXQSbkEV8LwRu02Fi
z40k4k8j0OozLnToUGf3LeUKB6cwpV7BCB7AiBkxwTjnhJNEr6AeUOZCsNqgEDtD
Id5S8QbrlPezuW5meZ+pwZuQ8tjhQ3U1htA6ueZ2eynnTQOAl4h/R5T0FV0Ymh0l
aAPmyTYZ4vg31g/+UNbyIBwSf0oRHuNosR4mBr/Z1le0o4TJV6I41JiWKVUqHPCT
2p2issJlqywqH7c7EtIO3bjqu6N5mC0mDaNohzpXwLKXvR3FmnWJge7jFlZAskhk
xyie27RhAVVwquQ4eC9+SdNQOnStIzZoIaUvw7bzpoGyQW3XUo/kDmFj4gCDO2+E
0SX9lui35wiALFth+gF/psz8L9kRVrI2DQR87tigbD/mUNxjcuPr2AKbu9ijQrrD
iIUFyCQ3u+H5fUrlHIKUUIwxiMHVDF1q8ZPUpP1PlxfttFdEHfT+i/iJqDMtfc57
yq6Ai+mKSx0IuiQA1hgC5fMUjnxIISHQki4CTIOUTBBA0O2vyhfCmXGmqxhSIQJc
3NlhXjEo7Hpj1eruIIbvKWdB5pdVn51eftaRLSku2IciTdop9h/jmZZg3CMMP2cH
eTf8OUQ74R32rbVqzJif4ciQRnQT9dJUQLmvUNuhmJtoIueiHDVpwnBvy/iKM6Zq
1lwsysRTvrHLybGQcTOlE8ohez31ZW5Hap3hkJM/g85MoCiKqPDV6o5gg9vzCPAs
chrGEzAI9hiroXQMyHGy/G4MTPI+DFtS8OqHOGjIc+6ESNC7gsdkF6SpXGUbrQAp
pzMGtzlYiFXlnYM9ODN1Droep13F1r1Hb5g+B8u33VRlSg8aurobX1GEZ9khwWoq
bUY2i4fTaijyo767Q/GyRCzlO0XHSIiLoOOgC/s+LXdeWyTUV4Ag8431Ex51PFTj
CRCpWzGtnPe1Ji4EJZ7XnNXUr2najHO3HXyLGe1AmNzxcY6CwB/aPj39IvA+yt2I
7xaFcn2nWKpJQj3YcWNc+SMaYYMgzp9YGWFth5Htf7VNOj1kObDxh5k1xN7JEiAf
PS9tdFGfXDo5PO6DnmIFS3YhPmMtZ8AzH92E1CV/NX6DMB1PqKUtaWE+Y0uiFpld
qys+6ri+4EMQsVNpks6a8fIVeVopZCk2Pbvc3P6ijuuEf4TwIOu94GlE5sR9v67D
COpHQCgrgyTP1B9uLS45tjNsNewF5begkgeLt5+ar302WHmwzLpXLpalmBA16Eiv
6WJ9uxpQarEpJekfyE1o/aTVKAxsl1jHr0geapOOLOhUYg/8VWdqMGn8p9rMceoW
FtmQum0nOwmUHJnub8z11yvC+CaZLP+YLevP/qWCcpydnbx95bB1n3/HHDUsLeCJ
eFyBXrSuymDQ7HZojS7TatuL9Dgx9c2rmafcTje1Z2/T1KaxkKByHS2+wcmAfgNy
lhqCg7Tf32TUkbClzfvZwcA84raFaR2nB2ccqVxlEJUaF6PkCIpeUkNuIwG267Kj
0pAGE9emzaBiahSaV7jMJAERU6coh7TGbLPwWRBNtf/YF/jERnYnfJLHMRE+ZaWC
IEaP4zi+SAXfmkU5xWlM/RMg9ge7DmwLUuMYeclYhyATkWN+jXk3F1+rzFCo3HOT
KJUO0wR0Iwn6gqca+JpTYznS3asXKauhNsKy8vCJyXf1VY3GR4mRgcn8zva2cOD5
OAx1D4ARGDEplB5kSMCeaQ0KGJSEmWuMFunvp+GedAF+nvXqblsjq68ChmSLEgsv
4EXsl7ENxmTJBosEHml4kjbhk66dDUApf8vSwlUCqdYM4z/pnANRbZ+6gBwRf9bo
KxJFbEsyDzweTJqSmCkzbs2FCXGaMNI74IliuPCmJD4gr0OHLe6xAZ7wHUH6CZYL
I57xMYHYJMS6GwHQnMKAEbWTg15S2EMzW7ucBvPDJwvx9BnR+4oVSA62ix3alBAY
kb7E82dUBypPJS9C4sFLDnjZquVm60uuK1blc9JQWjHJdRNL8Vi6MfMsuCQ8xpWs
kpBe/3zlG/pOMbSyuL+ld5+QobDi3JMAlgzBK6EY+dIsYvsbYClB2XrYnWjEpea3
eCivOSg+X0jMJwlhEoovEPFMcK30UJXTtbnxBCHsbo5BpRLzVuJwP4K4K+Jb5/sQ
NWYWnltSeIZCwGzpVtS04Jmc+11JebTqVly+aMeeGMPApbO6Cx5A6RcG7RPr1DZH
bna4RmPTkG91zhJpePZaEQc4dPuf18o+BQSEfP9bREY39bgG0hbzm8b7Nk+0Nbd1
mcH1XkbQLnMxudwGaqqsw2lVIJxkEYPgvQ37OG10EqTPMrV1DtGQ040oiqYTmmnF
FfZ4K3MkoyvnbxWKyz9GCHW88izagmO+7qXjD0oBIhU2/KQlAS3L5te1r159vNXD
DJpBs3e75cXEd8Oh0I+j6Mffh3k1kCtVwctHTwFzwI8SBS4nkbMIbMX4tE3EBLyk
9kLaBnPB2akqiewfxH5Yphf7Vjn8a/0IrRhgwfkwu6OQHVS6ENUEELLE82ySjvxg
bAuv668NZsJb12rA4QdfLpLuan0vpFIXY9cx56I3tvW6Ctwjg7pvDMC3KoRocw35
lTD60fxNS4OIE9nEJ9KI5GCmS7ujPDzhlg4TG9CMONOJ0uilzJZrohMrLtNrDbD6
AeurrkzahAmIlDTugZPlvzyPKTv2DtOQLOwzgJ39N8KF8CDhKYEC6jZBEUJLuMPj
ygV3s02VQoCuSUlX4jRpfIMFdSf95p42CXz3N5ZRRV8ebBTA3AF0Ix5nkiPgLYQl
GSqcKYIbOnkH++1+bGR+WuRT+fe2S8GmAcw8pOqFCA4gSUFGnjZ7pAB10N0mGu+L
oel5ozC85oZ8olJ92T3kR6Fc6btMybJOlnQu/hCiPq6Wldt2hAoZzMw/YCpfdYjQ
V03U0zJeR/to+eMHMEs9V6DRbXtXz75DWlMl28sWfa3JXrHebtHXhdw6fC85ct8q
umtRFszh6YaIfiJuG4/64aT6pDMdAa3nWJXQDdUxApBIdIJkAjbk2QOPVXdTRw9Z
qQ+iaFzhvD1Np+00DVOxLyWlUERrTZAoGKiHo6zq4HFFbfQX9Aot3n5W9dngWFzm
CkwFWZj2xgqRezP2mZqADG+BTuI3HlCpegbPAV2TbZhTVcStQ5ow2iVwBZTSwlZb
NetMx2N75NXmSCZRO6ghm9r1uLB8Fa1iUWQPOAVDJiXsiY58A9j1EHxy9RHnXQiL
XrI1U9c2oeoQyatQ10dKug0dSfUV1dtn689WEYv42O9b7UD38OP+dEXIPDDdZ+i6
oS8tfU1WAztRuTmZwlJ9s27gKcYlCASHA5K9pjQYW0dVqUScSbj+XxMI+st201At
PcLN1Ff6MwXJ6Lz1nrjL1ffuy8mD51/Tdw+WuaMy0STv85YG5lg9rf0UXd9r8OhE
gIpUveUVbtzD0AQZJRflRS1dFWm167AWw9an3Fc2Dv9V8DWmhdP70CAzdiVcDx8E
KuGpERPXUX7i5EWs+RkSctS8B4jGqcg0PK0HNToybCPD1TUvnXKvNO+i95prrzpa
4pM4Pr7aHJNqUG/1Ih8T9N85zVYsEvkBkZcGck+kx6ErL83k1k6LV7HltBRkDQBI
5nMmu8nZfKYfLn0xRzY3r8U4fn+zL6ROhvebKRHb317ty6tLUwiyhTd+NK/Ydw6a
7h6A2fH6k5avYF16fNjp+h11UZx4dyrikVEp3pvqKxdgO4Z6+XmsmDO7ho9OLdcJ
g0jtihrNUWzGQciP3FHWE+OnxVt4Gr/xKK9of3uW0wajFFezYvrDzLgrt+MQVCns
xrZ+Am9spncHnkZLAIR5d4FbgigZgQ7ikvMF4RbZ+nPjYJ9hpaF22LTUJsE4J5MI
yci/S9I8w7ZgnwB+0Tdt14Vvt0ZF3TRdj3a71R/pfGhutr+iCm3aGJvHtN8uS2pl
niu1VZ4jePoxRhhk5tzgDYimkUU8MDFvRj2b5JoEj6IyLbaL4swf3eWvyNWXoC68
bosapfIh4/EwBYZRQUmT6uGa4DFKmAnd25XU//eGDfRtsv1Hiwd3TLfCgmzYyG9n
+V+xzknMJygsA5NgGxR8OrUI9b2CwxkZqkwdsQaeYt2W+mGOF3H12oqmfRysTkuk
xUxtVdhi65KxTuCK0p3jpdCt5y9wjDgwlTJoUQFFmq6mkLNxbAE1IGNU7Cojb8c2
Cx5dLPWSCpfWEmLfe3HjLXbh7mOkpTU/8vI59rD4E0UFXzXFIKm5RsltNTl/Eats
+8YUxELvMMyRx0C+1m4GfW+OK1SHCSdcJx59MF7z1ygVBZfh0E9wKVdZTWN2cisz
nLCGJ0/6yT7yfj8jI5qCFZSH1myafvnK020tG2VaqKBjy5GiNd8Rc7UiJogtu3wk
aeznhYzTvTiayE9cj6QTs9iZwU0s7VTW6/OxG4ZvU+zUKagpukKYNpej2pFBTba0
GIA4957V4QZCG6sIexDgpss0v9Iq+tB5VkkQ1jv2wS9PVdzlNO3vdHaSm9jdlbzb
G6zVjQkwt90dXflS+mI/AIEg36lNxTPhXwXyKl3sGkx/9zz/NDC0/RON2CBKK7FK
8pP47kX/0JNBV6D5NNhe9ZenZUzGOv/zW9qn9zqKC7cq9hYGYoyWsTTDXu3sfzrk
6FB+u1tYKiSPqVpEs5dVmfsRaTYy/ua4u1tup0+u5BwjgqMAydzu8wBffugddkXJ
RAVBPUQwBm+s6YQHOYkoDbzugY6DibZ3R2KNYS3TeGVXo2S4Ll47rwfpTdb5D4dm
Pzn/mS48801+m18G8iD0p1wFKj1aCs7lanlKQ5ISonJH5ZrSfEWIhl+/1kPgTsLE
toBV52t8+2S5XgFDYOsnFHD/5EpSwi0xlSXM1wzHtxIzNKVPxmj+IIJxSiDYYPce
y/ueDGdlyqvtPUB6cuwEAzY2QpPer8j1cv8qGpGtaXjl8ywIlsoxyijYibUaVZV4
86r/5TcROtTBrAcR+XEWsDYDt8cBsOz9VW5Io67MEYqSzzCFwUUw3027HD9a0hhr
HGXq8nFflP3wLdb7PqYGVmcCJfCj1ZNMOBIsRAMP2aYLpp/w9G2I0IB350J0EWut
aRAwrxboH6XI2YBrc6qBKHf+vE4RQ83oUDDGJ7SJ9Ygefzuf1S8lrJ9f+fRkcugA
Yt35MG8FJl4najH5nrkNMDXMmAE4WETBMGyRvisSWO2V1cN4EVdtkrpKTe1xoMP8
ytVpzothz/zLk3TxETxhLQeG1YlxXYYjIFrtkiwEJCVsbhXgD1Dznb1vfe4GVXTy
lfJkNicP3gDI7Fxv9IwZFC/cFb8Qk/jD8gpLTaAFkOPqhmN957kieouqNUSi67gQ
iZS1HntS2reoiE9m/929KRNOZVVgS4BP+9A1YWM4OF2brBqUCrtNmdFK3g5ucSu6
CORRUwzas6yhGQUhbzpUz4sLIFX8rcgRWMQ5FMIfAxkDnDWuFpGSEWZD9qa+JFqh
AXE8i6s4NjXChB/1G+el2jBtqTigaRZdyZUCpgxmBbyoG7RkteuLivs6W4VZpbgj
Cj+ApJeZTkDfZhclmX3QST3yNIp5D9Qr3TWJdCAeM+KGgsExuuyJcDzQ+Wokpj2b
XB6ZdXnWHWJX1odBdGHu+Hjbi0qmRzxcIX7ddHbsUyr2KDMp5KDyQua+bURqmz4e
G6dB4Tq6MTKnOPG2ZL5GhEeH1darqHJ+oTmNlCxPt/ZxXUBP9JcO47uoPEVvaG4h
2RuAc85M9XHRxuyXujoef9H95afzAd6m+F8X9FEmf9R9QBx/OQTDruwIG/Vz7N07
4rsK+3GCQSr+cmJXVSIAng7g9OzLhSpshAHXjENL+OCC/zPP1KAwzAvT/L3GVcxN
i+XkddpxCNfukGxssibuu0clHxqTmAKA9+44DAyQ+D33ZXmp3I7JlXIqxXT2Bse/
wGEMnvuuv+9x5ppd4Y2bFIjlGpuNU+kvmhERH0EtRZtQtUX9kVfRDAH4fdkZty94
wTyvD99uzg/qz+JPQ1aaShxtve3W7BXRMay9qaq5KRMAcM0Gpti+OXj2bpnFEA89
dqt+KUmZcpbHgj+cN1kgJpZ7OLERr0BcOK2R0kZftS9NeNBbUKnNCLWt4E8bJMca
qhVAe7fEwKnYwwd5El83xnpTLwgl3YmbOVLnk9uhPfkw1vY3VPdoWrTUXL6BYQAQ
NHutR94Ii7WNbsUTVPcxNjjf+GVuODuUtuloj74O+lduM5zL6WwK6h4cO68gOG8Q
F5ZEODieHXFJpTYPkgw2mpApo7ACR9MTMIPXt/hus7g45wT8rKdILlekUSeyiATe
owNLujtU5ETI3W9Mi1TmWgXA6uRnww+CVdmlNgYah0pdcZmYMT3hg58dNpy7ElJH
rrbHaSQ8rCfdnzPGcqv1z4yKLpNjlXCttYPHUz496uzhx9p0GHSkKC0PQ/p24QK4
e/FAZwiXj0NO7pzEl3vclqIhyELqyZJcapTz5YoxDbX1KoZRt3dn27IdnxdyIqGw
SV6C0eVGIJEs+W36PUQL2lWpt/umhw/cvVtI1g7zT9VYy0HAuHpnoAs32Pl+tzOc
hmkU7vjvV/2kq0fqUvUQe/F3tRQ8AkILu510DIHw8RTR2f4ofFp7hLRI8XWzSH71
qdTe5+7mPlBrIGZ+njl35m8YxFXdtGcwQniGTT7NUDsYs6b63a8/CdOhyKmEQJ2g
0Y508JunPLVatMyhMePiFGD76PqhFD9JvY8FqWpYpbw49e46F35KLuQTNViQ7UYQ
EVduYhaL51Rb+d7yU0b/lC4ETWIqzGyteY1VMsOcDKthpyXBWCH1zc9Wd+6UaUBm
QD/FAdZTRZ04wj1k1j9nXoatYcU4UYxPbPGWc8+0D7qWg8IAW7AuY87SF6Sr/n+G
lFPcMR6GOUTaH3VsmXudeiZK5hzinWgAthrm+R4a0PPYAi47IpeQdgueLKYXbb7V
CvdEUIAE+VfVBaFNFzITd8MBlJ7rDw/MW83xQ6UfofG4hZUz5d71tj1pyCSDONVh
G/C1T8xU7k60aNGnVbCk+u9kaBxjjPmVh5ohyXbEqPFArChBoigS8Rg8XWtvqbx3
RYGFLmXkO8w4dRkHsvEjdLI2se0SqQKw9xJfu460UxBrACREUigVFZ4gtS7ipHTH
fX7k72hx+nL11Ls0nZYZGvbkJXaw1fMPPCdRPGacDSFXTQfFclKlzJtDFxh1Wwv3
+WGSIPqjHS8CeSM8tKBxAzQ/q+RpK/WOEu/wc/fqF0+rKQDKNd0rsiqtBaDqab7p
oepofcYh2si9/27IqLEZ2ayLqFkR613/ghfuqKrwsOMKtNIcB6f7GmK4U7unirM8
WpEOYS5GUvSNtecwMQpk8GJ2N5ZfCZdDpDFjnxC16JJChdEWpuIVK+vQ+c9D341V
SspYkDepJxJee9dBv0hXjuRRKrDUr73s3OeI+eIQWNE=
`protect END_PROTECTED
