`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HxTUQFSZHlF5wcHoi8fjiV42VKutFFQI65tgvtGw/VF8q/yFh/6FL5ztjmWsmKzJ
ihVcRWkmAE7oD/bCVtAKdm13tSlgeVZHY+O8jH0P49Po4UQAIAyKsxQyr4CC9JsO
ZyGg4jytMo01rLeExfDWd7Zm48u+saU553q/Xfb8lrrPZHPdt0maM2riHNxFr3Kl
ZQUq1gPJpH2RjeoM42E+6lM3dfG25VyaQ74pqSW3gdTRUHw+n0jDYq2S/4TI+OMZ
bqKkH3NGywSa5pW2Yu82n1Qg5CKMs2ge5ggXoUwy5qTDyCSW+Z17Bhp9zQ6ACx8K
cQjy5XreE9N2PYnn/WWzGXip3cr5Rozhs1qoxptRxexdAnm9pR9PB/tFxY3eGxIy
XLQPNCxOU3Ul6qKg2xxd6rW8HVLqMB4bAJVqCwx2hbRC54Z0Unk9fmPMG104qlWx
GukhKA92IQqsasnl9x22lA7m/9MHc9KGM9Ze3AYEL9q6wSFwOCAQOfiK0DqZUn9w
XWz+AhI0TGbbYycKmktcSxDb44wAvNPaz3L7cA2ayDXFF71WKqqFcCXhO16eFaJY
R345AlfNwrEKQkhzwtfcMfCn4CYo/4b98W0v0s4UvHOXavFBpQtOrEkhrEP39bf1
2cUmhq8+9MTPoUHgWmNwuAepCTsZ+0HuJ1Upn74VW0mnP6S7/p2x2aPTfthiji2x
6KgDIX3+EstvWl8Q+mXE3qPx7e6Slsq4a8H1bCstWt8Obur1vfa6YBXc0Aoffq19
053sFRamwyChJxRS0t5iZYhvilti5iZCmVoPbcMEgTde1ZEfLUZnyYqjYSXcHtg6
vyB76sCFCNslTLltLVRwk6sM1nQxKYLLnSc24lRgqUtnP0zB0tLzAVIZ7w/WIGEx
9qRTEmdlN6GN/Zp/QWjoMfdWyf8UpgkhV1bppAwRzrBkXkIf9BI+IePs/AR6Kb6d
rB4q7tEqhdHYEVrjgd5dh/TtI8TwVNR+sh2t28VbVmGvb49cpK6SIDNxF15HfP4/
C01ICBg+p36hIjmRA0VWzfEC/aPoziWFPwWct9bozPk/1VpR7HOJO4bkpvE4o9C1
KgMOtchxae5cnDSbt8KGEcYqMvBMyzsi23g5CZA/UOaLcAW4AwhJSFCoA173G5+l
uS1R+klWUzjWZXl1SyI1x8OwNC1Hu+m8sF2XIukHYl1u2ndZ2KN1H7QC+rFJw0NK
2fkR6t9qNUnakn7jGDA/ChhdGbeSdVyk1uzrLgk/aoBNcJ1gSWWqDLhiR/yqGzuy
o5rON8aN8KzntbAevL/FZQ44jt+K+7WBD+hZ9fLnmUambhUhq/PORfyUXbaognXf
3P+tpO9JNHjF+PYpFlmBM2ADGaGeObLJp9I9a+Bm/kZFkcL9xOgm5T9MMMq4nPEG
a1OLoORdGuk+2UL5p5NYj+Kiq0+7oe2JbIWyqrsnbyA+I0E8q0d1UslxxUxBom01
45tIEHoR38m0E7k7ILYQjk+SeA8FvZgmHO4yOBcxdd96pRYP0kGyh0HpIiqJLeVd
L12r5r969BZMm/6dEXaXq+BMRCBj0POrAh6L92qdG99NEhyja+OXDlCDuYmExr+v
hGl6ir/0arzMu5PFbqWqiAQCxapCg9IljHKBxFk0erMC93GEiwa+15V8lXA/Rjx6
MxnEL9tCxIu6ZEpED87qu2if7CRnUh+IReQXJzVEQUaAVC+AAp6Klz2TpY8RbTc0
j1J5Jfn1fV3dvJmHyEOrrvA9PIiktJ3u6AEDDrpRdq91fIAnJviPQxDio8XUvYf9
p1E98s/UWbYSGw7lSbNuruflwtyHR7ThuRzZALQCygCQfIh5IRp1dmDkhA4HG4fo
ZhH/PbtRwFyamt45U1NbGrCmk3CMl9UTu4miyH46My8R4YkN5mkN37A9/XRwsb6c
7I3rLmR9eZnbmAsHsi/HIoGv5YofSDRyBm3dvx/8I//9yRFj1m1ntUiFYCHMhu/R
NkV3EhC37ROP5Q1Ans8r3pX37eguv7F4aSBCVASN6Z28pD+fJxlQvzBadopKvrCg
tgkkDFLCKwHUct3Tjam35Iem0tBc33vSr3mYNYK46ia6GRS6GroYvm0pxf54+LS/
0JYQhtIoP1GAKQ1tW2mv0jqapuTL2MhZ7wHGXcfYN/gmkC0A4HIgZ272jsosBL6+
iNkux5kVud92nRsymFaZI5cFhBw1wMvuBWrsDFYlzuZTjIfVgX8bb4Dj2FYLuQTh
4+iUn2e6vycXhDdtm8w6b+iZ1LKocuHzpOaRzJv+SqQfCWv/zKFnUFH68V+7KPoF
jJds8BHE34iDTwEILA1bQDHYUay0p2SSmAsb1wJZAk6EPX8FAjsZ588cQhr3fz0l
x4yDpJ0BGeRZ0qZCEBV9abL87ObLkvdR2UpFWEfPQlpqn46EfixcEBIeQkfvts39
LkzO+JDtCjoCUo3YEYlam2YGpWMkid61LspQH/wW7+mZOCKsFEqMPh447nFmhDmE
lETfSuzWUNe2b5ney3L8r/eDgR8/1aSr0sPd5V9hwboUlLZp+1Rb0uqczlFGpdaV
yo8fwiP4vJ73AVk+OhCtARH0w/u0WhE+PH/SIWfyo7xOFY/AZp9SNY/Bbj3hu62a
vIG9lMY5P5Q8usYNQqap9ev5L0m5De79jEMmBKMwNf7F1Pug5ZJ/kYFjrLja2usk
tPWjqcqOamnhYZosWuQ9uiVzb5VfWHY46Q8Hfn+P4OmKk656dHSYlAhWG0AP2vbE
ha7CC103ofOEQLXsIv62V46upomWX6bKHC7raVIQ0y/UGyzg67t9bC0X3uoLcRaR
+KsDHXDNpcMMT6HsqiFM44LRne2W2M3ljw/89rs+WxCRx/lZcMbn5j88wOYT0gF1
KuGtaPQ2th+KmnjgXPH7fPCuIs/360RtfInakzEXRJnD9V8aNtmbuwgTVWNG3Pn6
bfxJ51qvpwh3c9yqGm8311npWfDuwcJso/6jiND+Gq7w0kqT8gzu0O32wY4qd8DP
Cf4qoAZ1k+qqjYOQZf+etP/FJqdPqdq0V72JZ46eEz22qJmd2nyIkrv4veqISk9H
YNZPR9H86z5/f/+2SIs+PeESIBteZleaxBgrBeBnXksRhATISVCDEQlYQCwmvE9F
GVwULwKfeK/qk5Dkqc+MayrkTWTdXt89qT0fLSSMY0YTnq0tw9NG9jR/L4kuRwxd
yEYIDjJAlfRl6083wcQMiMOzgp/yG2PE+0M2BSB8iUrwpVpaq4haadAw051+LNZv
gF1reKICusmyu5VQM6O0Z3EdiUowIpdHwD2TVfFsEQ1Ps/3/WrYDs0GMw2TZ5DyK
lzwFMd4EPTe2KxpD+EmniHe5oofR0W/R3yJ7WyAUsD+Sd3og3nwJQema3c9HWMop
SRPQE+KINer+C2k1LqGv6ZWO++I4HI2+275hUa9pMzFapucbSWyAmvd5hIeVYWIZ
4uxrwgFESljF8dnAzBOfe2IxTidtYHfGRX5Cf5QDLT8ttUU+TNaH8E2U4qcdRK2u
uhQVpZ7o/4lJzWy68a9hV8awaGOUIVkB8HWWVmNXInoaoVSENP5FnEScBthfph8e
ApyHUkH3HO7RNGG9vLru2O4bcSqvVT5Im1UxMxBrG1WQRJtW2ZNhpDEndt4dNWgM
jGV/bHZiKycdO+yehhXHeeyttJ7Q8ZIb7HEa3KVzfA4vJDcZRPqV1699CNCdZqgX
AMXZVF5IuMP6QH/mViRqyaDZfU8mO/DGMmR+s1X+XLez662RzkLKy8H7PPqnmccX
4Ymhd9QMe06JbL8+B0uOO5eyXtpg3rLJGx5BqEfCwx+wjGz0rHA7h7FZ4nupeSas
MErAogE9ze9gyw/ggznvOzk3CedQaCyogyxGayM8ZcnElxsayhPbu/54fVvTODkb
XhxOYwAaOyMYK+/IB5Eqp5HkkgZo7MHtddUDdJe8Dc+VyLkecPQgm3/okMGzGtCS
DkT8tHFT3JNvOlKoWIiNZeA2Typ0BJzGNp/Zf8RFckgq5WsJRB7herAscb3FuvVO
zSzDdAF/SG/7U/vsdL3XYgBT0UsvtDESCjKSEfivqi1D4sX9kK5NujoOCpQpc6VT
v5FE4u7SXQ/6PXH/ZRXPZb00k+v8Zf+kQD+5x1GLTCOGp5A3A+P0zYWUqtdB1y19
7I8eb83F+u81ZhG7X5H4vKyJZ1X6BJqENkzRZkHzAHviUB7snJlqolDK5/96WDeb
Dptn/94O+1qK9PfE6tWRNh/fgRNiWLc78TRWUhnzgd4MKExbeSsGsbndWp5+oy4u
2w2+tQZ19ILgBsdnkQEMlptTtrmqGz65FnBjUcJ5bBuqmh3xY1Y1lhJPtSLej52I
5ah1CixhPu4XFKWYHcnfn9yxSMgAzI8ghczoO/PEI8EI7a60cTI0r7vkaSrwYSh0
xUnMaaIOYOxC//wIGisS0GhqEHBJZ9AgcYvpEI8hqPnRzDpf/PUUt2/Jf23FUAdK
TSEilemuAylSYHXJl0n3UcO2XXhNB8/2SbcGfpCs+xqTfOR/SusSS403kn6JHLkn
gEIN+5KKwZ1nUOxo/SkMpqWtQlYdKRwvCmxxiuTar2YigHNNdUPP3gCA+jVaDr16
MwXh4/fg8cwrFFcmbMIhqZd8zsXYNCGGWuw+RbNW35NFomAoJCnH0DNG3vs0b79O
fGCN4P6mL+qETWl/DwwLlO3WjCOq5o4MxjAuWRMtKDY5Ljg/8dp7mfxadDunRH/L
gbE8ZXR4EL3I20M2TR+KmMWTwmdJFhKfTDjkduE35TM2MbQJHWLd3IRWg7g5m23E
wbEs51WhE3HPDdox29nLKmXTA5N0RASbr8F1BUZVQeKXe7kStk5yJ+z9T25C19zy
iwEPjjP4FGF4HuPSn6EWkNols0PAMj4gDS/u95MVs8twLMeRxz898N6/n4x7BWik
NSPkr7E876iliL5ku12B3gNxN3BulCm1cLTbFILgr3YerG6d4S2VKlnZazH9abma
8+9Bs2x3VFC0r448hu4kZuLfnnDl4P70Dupi58r7mLkBYjLxHBf0FFcLJmV7NueM
af0q3FwmCVK0iCsaezqp4M/z4gGtFhPCrjioG/TygUsSIbL+TjbCpvWIMV+kDSVo
RRn5jEQB1TTRQgFqCsuIsLpO6i8mF2tFgnCni2fhMEt/LsotQzakYsJgO6s3EnsA
i4R2Ib1LDIOukW8/3i/JRnPznSIm0xv4OuiYF3ni4vIXCzW6t+AIdgoBhRAW3hNs
Ai5VF92VhSLVZJg7D3eiIZRrI0Hln74fH1ZrXrYIP0Qd4dskk4UiUoFParYc0nKz
S5pPWoujsaio0vJdjlDeuB2m5S+/OnUgLtlJmTnmUZHB8NqWAIT71W/lX4OiVgbd
LVYo8vS5J5sHQFJtHNeruFRBLxCoe8iX1KAPgL5FAiv0n4+GF8OhqlVgC2JgkKYv
Y0iXOVtcHa54wwxynk+J1KxlNTjp/PaxPo70yHj6i0edG8rdSdtzkmhoXr46zIT9
RfrVpMpaVYs+qtYRos+IRhyNwLPVSmOaX+kKaUuxDCm57mru6qCS18OYRDu08Yjf
piy/HrcHhdRWKpe1lrhVV7xmMpQVrFv1e4QzxJVAvrYZcEt751VffXSEmdzvLcto
/Y5GIgBpMLIq+93/mI7FWe4fuf9i3HNYaJm2oP8Wfe1M/XUJjHuMTeSvUwu7nzwI
pS6H1i+QRgbgUm3PRQaooTIXh+3OQ1GNL2j4NZuK0onepwdqYF2u5BPosC475PwH
4wl+DoPzF4rjpWL2K6qJb8hp2njkMKax3Kd2fNeHsc7/EptY3CfjnmRFI/dKDprH
HqtrhrIzxh3YPxCljNAWG2J9JVf2bmBAAQofec1v24pQ3v1ljbgZOOtFhjeA9ahf
VAc62e1AjSileDJf0SxNQv/aRSY13LsENHQCo6Qiw5ag6nvNqZP4bDp7YajXwJPx
HzAQuDP3Elk5Th9FsLhihQ+D7CKq6j+iXTWw6kD2d5rimS8KaCYPxkTzbomSmX4S
cJVzyLtu1DkAQ7A3Iq51NMeWVbKnaEey1qPqMhR5l+0YTOqgeEBiRXMvdaS4gG9i
Sg5KyxIsAOGyCSpjJ3wbWGPOXlCUgw5EpFNduzQGTWYEmnURLL4uCcqHA4tyFgcK
ESDc0qnwaTkL1S1PnFRIqCbIbtKUqMQlHrGttA+X+rzrNUycjNTrLNjUSQTvhzX9
5a+pfyUsq3SmZMJicZA5rRFk8Gb5awwCiehcDSpyIvJEb29NKRIeFpsj6Tjg7Y70
EcCw66biiYGe/PGKSuGn37VRmVrwkkWpgFVSzz1AnPj2gxe+p0T9GDCZ6qQay1bF
yT1A/ULsb/NeyoPDE3ftxj0HddnOhNWU/xH6TceFbx7ZwThbGjyFwQuXGw6/eJo4
v5aBuLdlsRygdEIm3dz0mZc0T5S+xWso/2bz0EFU9V5D6hYUySMDLF3B7fAuW3f1
ckQcL1pPwd54rg2GU7u2370pJrFSBgozc128LlwkowFKeEcQMNHBLNSy+jHx6xW3
DcvGzMFzITbqPO5rg7Xny+RjqVftyNld9tqSmqb+zwzIP7XvMWDj1xhFpZAk7fvY
k99P4FpJP4Hlyuf65NgA4+Fr8jFlab1Iwl3LzqfjvuBY0ejGKKoV+XEMTZh+x1uZ
XD/OCR2TkZPs6eIBhmAXINU4vnZDn79+OVcqGWeZXZ8arJWX8TblU4dRtgNXxHvu
5Cf4PIqKD5F0pyOVpEJZxuVRmLwfpdsthZM7bvjnCln2JXdQu6e5kEvnTTgqPogB
Olfw/VmXLB/neOLwCWhycnuTLtFpbzl6CqPAttt2Q21yC42IJ2fGy5NQDUXlk23G
7HHXh8luF0R3wb1T/F+H7eSpV0S1wKFuwEx1m5fWLyeQ20Zn/i1b/HI7lvR9eiha
NQ2mvRr3wGxSCDSNpoxBAB+63qcwCI5HyZKMOkyR0mqiLkLlKNBTaiTQna38avtj
L+tN3S4zbX9DA6T3RW+ERqk86o0hGbR5m7Ufo3a9xcuEc3uioB2Ac3zmwh8FO9la
my/MxYMzuAKDvAbdOhnSeaiVe5bZJth5NmwXpKVHP2hEYUrzbAbHlfFpznESH+W+
yO62t6qsw/boqaBxUkchnngN+vDnD1T8AimvUG8BBZ9+aYPkWp8MydiGMbV3LCHd
nyAlXpLTpOHCUiZSm4z1UNRrpHo7EhBUvhX4Zkfrs331v/bYFvLOL9MO36qIjmrc
P/SwxqXZBb18iNFuMNrae7UZlN3IVRMhYKVLZHcgssFPaZM7FB+YP/dJUFHO7ecv
g2n0pgT60XYmk54Cs8smxvFZbI3NecE5Df344qwlqsZG1DUKWoHxvraO3m0G9Ux0
RLt+UskP6iLJZzcUqWry5Va4UV7CPYMqta9xAs8WQl3uMkWmFBK/s1raKAOxezcI
HRNIq5570E3OD0e2Vz8ZLO3b79HQ2P2apkwOfcm1BWm51VGW+RpUyLItX6tBcGbd
64TNnwVUypRFQEhrN0YsoF0YGyYvHXRijkl6JrJ7iGiDjJQ5EMCMghuywn2Y1TlU
NsnHFN8DNA6KbssCY3AaWPVilHkv3lL+oYQTglE54LV8BLnorO5bFWZAVDmfA45R
Ys6daBy4R+VKK5TJAcxstWBnuif+o9g+YngoIXpc92x1gZeO9uCHf3xW/EyN/DuA
cMPvGykls5yC8qn7T9O7iCmlVgV3Sm+A7cWkOmIuemoXkoXqTHADtbVEDes1wZwr
6bzxW/sCBy1Q3rjzKeAmvfhaECDx2FJ3QWlX/haIF5BhhPuEk2dbWuf+9tqOpZuu
6+V8V18qPWJpp408yQ/GGPCPlwk5Zz74+Ir6sxcGD7n4uztZNwb2e0RG62DcSEyY
PmhhQsPYpT6YLNAKnLgl3pq3qMeJdvVriUr8BikPlc4gZ8uzaSHavXG3AmbUJnXj
ssOVEgPBdqtwkCb9LDlMtSJ1CwZ/J9wDDo0EQ3Waa+wJSvdki9kH8CnGmhvqy/Cy
/WKIy8dqtmEd0ET4XpRPISzXEL5064PAsWl5mFS8m/IRQPOqKe4ziiSIwiDk9nAk
vWdYsByB7HsQQ3siOKvHpd4J//D1FFJrNhrutio/rwJWOjRH5vj0idLfL9fT6ivp
l2cyJUWyqcRyfGMHAwZAv346vIT8Tl90Aqkf4SqmTMR2n8NJl+hPf/AuThgO71W7
8hn/dWwraS7v3AqVqQ1vHWBV/sqMmcEoEAuY3EkbjMnibvh96Zd4bZTO3P8x06OH
6+I2tPapP3DRC9A/aS5TS1gCQABOgqqxzzU6Char/3ZSpOa2L/SI06aLW3YkyGsy
FuZmSLhEqJjuSuAaEw6DK09cJWKB6F1WxeREUqytrW0jTXXPr4YEKiuFs2vbuCo2
YtjdfztJFMLzkZIgad+UQlJb4zI73/11gAGXneqvSjlZcr/KnNPwPxdkEftKzOGG
5mBxsqi6+7cegR+N7XS3pSAnSw2PiI+ve1eRLgqMwj0FS6mP0W/Grk/poDRRpufy
8OM33GURKYvFRjGkkRhnj+eAooPKX7hJ5IzasYZBQdM1UfMoVt0Qc2G3kgMDjGeq
hNZrbevSsfwKrVGiIQrm5TteGZRXty29+e4kGlS8Fb+w/vOIPsP8hWQla/2TyeNe
1NCQsa24guNkxTIP2wmCjsYeU3r4u/LyPYJeOZCKBTje00Nm2Bq8y7IJTBpECRrn
rukgzVKRfgixzN01xJtcJqXoplxvKxJTj89NSIuSYYb9u8/r18nDEDxKTQSSVshS
K3TqChOUBAh6Ae94ZC2dQF7k7T5qYmgkX2swzYisFJMtWLSAMCSP8ZWfQpO4HPEQ
gAN2SV42Y48qtUWC7VzHyFvH5/WR0DOE8kjgM6nbohq6QdYsE12kCabYNIFkgHS4
hOS8Chu0e2qkDjkEgSNQmtM4TZy9A01Wi50AElsjZI0xZGqXTOeaCDje9VUAmM7C
ulNngHR0Q9AueWl+Fmhul/FP+90VVeAGH9kJESjWbBgxmopZsWETfIEsEnlKr/YF
cCbC0aVdvjHLfX68YQYI41RRlhNVC3qV3sNnK2FPn0XYqVc46TGYUMlmMR93dMvP
jh0sOXP/ffRCvWu+zjJBg1XUP33OpLUoEUkRw6rl8akzmsZPU9Phi0qm9UPlOo8l
32jfm0/Ukbh2OXTtagR2DRF3+r4vAhY/cuQDYmlVOdlknh+F7IFaSaHLlEidjizj
eXE8Yu3+MiYUm/3hLqNk2Gxil6vM5WPVNRBxi7sX8Aaq78cQ0kXUishJiyZsPGf2
GaSA7msuVTes5wx/1+a0zorKOrDQyD+BIYgs9Q5X2kiqa/fhKCtvZgzz1y9D2swj
ysZ0YkdzEVgZk+KHBYg02JLTfkki06JuzdrUZQqcoIWI0DGackiaN6AvE/L0szsJ
gmb6ZOHlBamfKlHf2dp5g0g8zwMYmuMoG7+W1mpAIFy6mhkpxdQePoRy5/Ew8Sep
TZYmgJ/uBSsz/bfnMA9n8sOPhmKGeh42NM4M8qJgY2IyjjEj0xsDTDR3xK+tdUjh
6ajIa4xbOVF+Nut+QfbZE0ihH5VH8OKdr0QuAh5t1O1oFCQio4s9dN9lmXI9nB/3
wW83cTkXN2Ol7Go0zv43SCOZM1Ze4A9qraOpt68nhv2hTiFwXmCt8t0os2sfz/Wt
sJqHWLPUp+dYLAk78794c5DKqxzvPnh7m0ZSxJ6n2Z7Gg/Wz3liMMCvskmjWa70T
hkIC+lTy7ujF0v3GvRNjkH7MYpDulCWQLpY0ElEsQp7R1p3Z60prqvR6Ardh/8WO
kjQ42HLJ3CM4kXxIdBH35sPFdlixwdH7UfUrUDrCT2Q+6mtg91ESL0krYD68QqJq
ZYPnYps9AKPi7ct++8J+7rSVLXoxC5Ovrxbg5oo9G0kVBoRdgdpsb0yvcBcZpWoM
GQF9j+PiOUZACs6yeB6NN+Dp+b8BHPBUQxvhR12KpxkyeRcyXx7051MwWQfC4nYo
oFFOYwmuekw23bmuxkZFbdDxqzr+dJ+VOhvbOBryEJyCOMMctHUSDd3UHNIgPgNy
hxB6LnJvHAjKOPruVAIDdkv14VDq1+py35/UUCxYMHUyRf4YncSCzIhF+ZAp9W8X
T9j64N9NOYjjDWcjp+CKAgDG/0CRRu0yncfmW8RcAfkv1fXNOIV/SqK/kFjo2XAV
BGITNJYYgEVwvwLDaKPAfZJlnrN7iAZtpSsP3wRmxE8dO8P3Pe2sJyT1Ys3nblXy
gP0r8VoY5lPJk1HuzmaqYka5pxYBYh0d+eysakrzWkwvfjBS7+dKoZmrSScyc6VF
0E7qKuXxWvsDHJSYsCJg7lBT6mtlj26uBXu/FuMyBGsA4o+kIctKkO1Mm7IcvwTM
QvtfiSpzarJz2CZ+GbKn2Q0FztnJIErVaLL1JbKQr4R0k1bmpuJyFeSLbmPEWnXi
NT8sF+PL21kc11G1Klt5jg/BWAJ9uc200JtgABG3GfML3rstNq6x81T4TayoCGAG
MAVoR808PVFRAFYH014X8RCS0dNWeqtaf2KnE+lkfadmsm3jbU7PATMzb8Nz3n9r
TTR2J1HjNk9Tdd9m7gpdUrmBWgL+GIHUjIqBh43W9QoHP0/B2rfgqFFgk5iN1qpZ
SlG6tFhpW+CdOEuYlVOe5qMgWavp9fzP8h1SE/gs5Y0xFnW8N4qTLya1nPDK77k9
mrLqqnOEW4K74TCOIghEfN3h1G91C97SmrG5Uf9vfz+bylDfhSLRJof9xAR8coDZ
/K4UC+OdF0t9ZmAL+Uj3i8iAJLpBe7MpuRarKkzcOJWSc7I3e5dVfGxPUSdiwyxm
DZOxClWVn8GAl2oFDZCu5hfrN1ggq1fQbRzC7uhIMF8=
`protect END_PROTECTED
