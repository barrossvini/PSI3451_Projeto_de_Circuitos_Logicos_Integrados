`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRK6tnXHgLDM+9S11mt7J6TsDYO+TRQdCs8S7MxL3r5zyGg/Zymg34CvDiTTbTPz
E5gmds44tqWUOpR+BSlDnbHtC99Qotrp2z1/ZMRr+A+6VcndLX1blAsI+kJOaQFt
ovJliExHPCF+/cm8ipDBU5J/k3OxF1jlcabqGm1IeN+Uy79AZFCkRV8FXRYRMEiD
miRtfaQX229K2c2XSvInLXfs/Olsn00ASX2hFJocYQdQLZ4ym3HoTAPGcRfJgELU
dHpEhWvcIOuYXbJotAyGohRRDdg0fC9Z3uEWitF7qgTqBki0uW+ELHgCs/Hg1wTm
TyUVTmnQprUc4YhYKCV64jzWBH8WCSqV0lqwa4o8PZ12aMdFRX4NjC6c7LgeJA5g
+cW+nfZL6yzl/I905hqf1ORPIC3fayuxAyHC9Jy62kMjCDVrQvor3TmaxALC0a0C
PXrF5OR21Wo5KBgBmX7uRpP/K+jMeYN6jJ7n9mcoYL0ksyjO6hzLBXo6LSjKtYRQ
buYV4efa0md3aUP9R6ccXiGZlnS9/KEFInvgf1Sn/Q1l7+ysSC32MsbdtFaRVjY8
Bk7Tx/xQncsADnKQqBtxAc4hC7NVbKppETuP3lsDIgoXW7qGqXqFio106bd3WRH8
KuSLwlMCxzXMNAX/XolvWON4wopXIrSIpTjtZ18FHtEv7yh2kSorx2iCnsehLBa/
5Rp8+Lx6JWO3uCx19CpHCB53ZRPzj5gb11ayHRS7WbCoHiX1su5bX4H8cFQrVdUr
WggSHGEauruU+C2b7yhnIPbjstBSe7eLUDIAfKqRrixPYg++UxYCmTP2RoVBhfzA
`protect END_PROTECTED
