`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z4tPnXGPLjB9YVAUKir/FAsfW7oGuR3k/wvTCHSUXSwTkcvE4elZdWw+yrIvEnjq
StvkPXCkpDOqgcCuqpW6mqWAsiookN5kLSrumxYoaE7q0lmWyOfzSIg0DAZZU2J/
jENZjItV4tJyOGQKJ9XDT4dzX3sLL7KJtfy3Bq3RieJLro7JlvSvhKHe6n5jTpvx
iqF5Kbl9X2WvZv5uzALvYVa6WSeDg8gl073O17ROKocLQgwAyTCJHJhXauY2QtNI
3rTCYpLpYAdIJat9FP8+PxbsCe+HLI8kw4z+oqaftOQeM3YqyNPg8ndfaGymNPuK
jLhvQugrNTvsLckrS78VEZPvD2JK2GQjKW1gDwkyfl6f3l46+jBucKzASl0QGEW5
mkmBhP8S6zVA1g/UfoA1ge3ryTl7ybhKJ08BQEWkb34vL2AHZC8QBkMIH0NREIAM
kxao2zXdTRhCeBjUEn0FfoIAne0JzILLHnGJo6Ug+MuCl01zlTla4aDjLJhHLugB
G8o3DL9h8O6/IOZi9e33LtWtFBrZhPDShqrtFIdRwkka5321+DWQpeo2JZD658f7
2YKefI7EZfvqEAU+Uah0yXsNL0xaYcNFc0ZLf0tAz30Vq9HkLWfI66ue4o7QQmGd
q28hOb6xtnXSmg5bIpDJct879iXVsm9Y5XEwOGWOuZ9AaNA03RagXn2ueJoAnHo+
9UMWOWH7tySte/Vp6agQN5hUdu3psMRAZHtq80gQ8YS/Q2g5bkikuevUu4U96jAb
iUcpO7XF6O6AuEATNSXgBtY4Mhh6VAGeOIdvikwj5pHwlO5+x1dFnShZ8skFifzD
yc1HrKdoVy/1mkTfGgZcVVmyITvdVkkSD1wE0bonFqw3RonJhzm+TnC7GGPeXnYM
RMOTvFeQubGqjfO7HEUd4RbfmaKEiEf1JaM0cnS+DjwR7fqu7ivLZgQsjHukca2D
LUijNDcqkV/kfZXhSFEY4k/CYa4Czti1y1oyGC8Pqb/9B1Lp/f4I718wwREeuGtH
hyscRwV+1fsjxOq9i7g+Yu8QHNWJWLZZz04nZv4FScbOO4lJ8810vBSyGvpyI4ky
ol06MtzSDbPVOSkuXjDd7G9ZpcV+tMTIfS1r/eZ+24qi6tiiAC2hB3RSEGeqrVm2
lhSJXEEHJtChiyKPctkZw6brtYkDc3IwMtMBzY+coE2/lwnCzkcgY0ErLAvfT6Al
i5UHgHmMdxBCKXv8xvUJBxz4ZlRea685HAf+2w97DxFlhRbs4X4X+taRGZ7RoKXm
Q+Nzmywlg24lldeboJLLFZvbmupgx36IeGMyypatgCBxmLlHwHbuYwI5imhRQl+B
oDNHp/Sp8B8Vj1VtmTcfZleuZtfqfHD+0Or8EoWQefaRyNu0CN+RSSv10nP/gJZ3
QUT/eCJmJ+uy2PXloH2dG0hkPY0zveP39sBVt65GM6qNpXexnqz12eP/Wih/JgV3
LuEWXNxXERk4OCu9WKu8KDzrRqo9PINPp5hEDGp9i6Il22cNYeF8gb5MV5YRGc6u
PLPa7tdpSTtm3rbfk+Ao96sZVFL6zJCW4Dl0J+YCQnAPnyrSEXOcCC3tEp0RxJbb
ygMZBEa0v9wRc2990B+U9V3gXOULUmDxiPoVP+Zcx3hnwD5JA2Ii8wJQO/qB8j1h
R5/pAM/OzjTZnzDJ01XaWJiMjM8WqSsCWvKNYcOdgT5KitDBm+wXv3OV/j0KfTg3
gXTfeahL0MhelQNGuU6aI8Jv0xIfC6vgUqLKaXxwGmztyIIzMn13U5zYq+I5ftcF
W9Z2s6OehMfQ7zJwRkVsmmhzPtfOCqobldtGq6N6dEMn72lfbPmzRh1RDMGxqbmn
YVjId6esgEwdgEtYClxBmpdEleiN/vPQamPqaalHcOfEGamicKoyngy7ph7+TFhq
g9IsPRYWQaaV8XwSmY9vvt18d6I+ffnecf73+zWW3afH6ivuonuWRDLa0f1C1HMq
2pmxp1jx2uw04me72nsADBcdeyh8ZEzF+BTPpn59spMvtEOqfC9EadnJ0VnMfxGP
EHpNofPhYwD8fGiexI0NQ3c8soM04LXNHTGS/5v6Zc9+OqNKKW6oRoqGqs6xrsvk
dIJ3sB3pLEhoVusRUM002lanzRpvv/2WdFZJYx3HL+nEby2ZSA49d69fTzJY8XoB
AhZkmykJlweaUbhsr9VmMQRzzD39oeBXhUtcTWxyH8SZN0H9OYbZwfDxE2s2xNzb
wC2BsLz/TPZ3Q6SCDmT3+ox4UiLdRNVKeZzYqQCZUAkhGYCAb1P8tR6qqeCMLQrm
KnaSFG1PgyoeDZ7tLonkwZEoaG38sBu8T9gyvxXh6JwGcoVEmeJaNpX25r8cpWka
ndaNsXlt9fTihrTWFRNq9j0gHkmRhH9pB4ksuSH2C79YNCbh7QteIj1QrJxbcSPw
amgIKnFvgiOqD9JT2vdDGwAGSa9x17/fj7FohQsUTWI1r2J+Ia95nhCz0K+gXq5L
n+oTknPYbMH3v/mla+3n4S7zSTCitVjONN+obBWOQc1A4+fVKZV//2029Shxq2Po
`protect END_PROTECTED
