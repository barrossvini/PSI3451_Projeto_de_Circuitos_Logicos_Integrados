`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eK5454BcvY/g7igjWoOgf1H7t1d1Pf7hJxsRzU3GoFyL8Bd3J34WSxlEFfX+WrL0
bM3JnSFMaYqDOL34LTtBzTE4sPc1vz7z26KUVji7G5hbpkpkJw28ujcfoy0BiHNP
hRRJcJTnPrO4yo6PMOpqFLJKNsnD8zS5KePOgOVfpLK6Tw4Zd2Lvol0UTOgLlqvJ
G3qHUi5ng8CaD8Wd+KQ1qHq7UonF4sR/kxJvhaTElEnjvLKDLZ7gCP+ifDIi8Pu/
1bao3ALpuZWz6PjQss0Uo40Lyfoywv9DvSRJIYc5z3lzOJacyWNoL93brdZoLzYN
nCkDDk/elXv2In/WFhweXUmjrYxCLRlnJ+t+yBR0PON4uRwMXL46v5fwtMOjlvlr
V7uxG18Ld7BHDt0+nENBW0U1Ax9yw8tHgzZR3ZSuJKN79HlgxkJRqdhlN4qXH26w
Gbd7d5jfK2Vn8yUo+/84k99XhQ3MtjaJHrmgFkGzsdu+EJNtj5Njf7poFmRMoSmN
jhnrzb7XMkBA6rcaP/L/FOW6nr7wff9sZu7BWiKeAGChj2ZOWU2tGz5de6HGw/kk
Vr0JbsgjkGRM1rd5CYY8S+JtAABgHrVdwHUPlmq34hJtJdKFGVzflQ2f6iwuDN1i
PorDq4WGm6lnXVvKFKg+U9szT3yuVwfSKw/XALzOdLsA6qthlVGO1yek8d0uUquU
ZH5IgGVRh8UOxdFkluojg5eKlqKErcJ2eKj259AYILLo8Pr/YCQuJtK1vEdLKlRy
k6+y94q/6WcsYbciPEHSejuD4HhJ/DBN+lUsuEKIfxzzRGpEGryFQN//4I6JFTYd
uA/qZhUKfyNTT7sO+Rlj1Sn8oI0wx7qNztgK2/hLWl602NaQlIPP/d/XDbaJFwHr
AhmHEumbmLFwptTShqldSFc/fGxPUKJTiNIkbBBpXapnrtDuPng9N5HrABZItWuP
qB/04TyyKrL4MjkyGqhc84J/XsysvXNtuSvnlvwVoeyGlrjGMwVxr6YHInHZVfPL
SyEoxPumqnb3MHPBhYGNXJNg+y5Lnb4e5MUFzX8yaSRmXVb5BGEubMj8LFAJBjU9
GZsr7GLXAv9xOo/G6jnUaDOW04bDvmRbAR1kW4N+UGspNdgH3kg0dTq9JpOFMZs6
6/sRrxgRU+uU19E+awVpgJknMuuHz9Wyf8bR2IajmUH/QtAkstXEhyinL3FPtYgJ
nLBVAn3K2OL2BY8shwSatNWl4W7bEIXPJM7NmufcOtpDh9lkeZaxs/1q24dDu5+i
MXjnfnBimYk72UtXrf7E75etWlEcT9vAFPA1lZ+imQUALB3czdxpke3I7rFtwoCw
Y4Uom5L9cEIhDhITkOrid6jrgx4z4C4Jxdtvy5gB/kreC6Dml5MEFm7Wn8MXj27z
EqJRHVK2rNXEDm/NdK65/BAZqgFJRVpKglQkEC3FsQvJxI0y5frumjoy+48xWCCq
MFVhYxRrg4xevDnG9FtNV0HNLuXVJ27QC4XXYOtiMR2MLSO97Lp1NknaxVkWIM/M
EgVyacKU96RJ+9pdYQz+BOrEjem82dWCbpmMuElxgxzWsv+oZbnh8InhjZ+3GwQJ
qRP3m08YFM1/vw+uex2JHqSRURRCMkn1T09SHQHUER45kk/uHEINzocRL7j8fSA4
8lqhJtLOA8MqvBbJdf9gCTqK72q/A2QC1mB/puXAjoiyxjG9iMXsPzd3JUaDIWdj
7o2CeblBd+Mj3mswka6Fk5rAbZzaFnP3/da/VFjud6+vJ2DTPeYreVOLE1lE7qUt
RdeuDVuD5q2570ar5qEobjN9c7lxQYxbipdYC7/2+FW+36q419VLuJOog3jNxm7B
Vw9d7U9hY60r6efmPmMh3gNgTCGT2IcyVZl0um+/sDDyfzoyLorfzNhAGP9pR/Yg
D07p6PJiWm7757P7kBnCgQuGKoVtvxEgNl2uO0shPBoRr+XyJvEIaGU+QVWgQA7d
wnWvMr6kZ/mmeNLPprd5x5z5rfouyxVQFpaOFWWrtpe3ppdcNVe170Ij3Fb8JAfy
c0vNsEMymkVIyKkdZBdLkKG1uyVaXRd8/KicaVx6fx08rG5pTlyw1n1McMu3NBiD
om81FjhZ1DC0hXS3hB2SUOOhw14mfTbLZq+Jd7WINNPhGErcw6awuABq+jYsje3p
cwAUzAg6UvFLLBI2y/I4fqrarpwkHuzzBZCEeQvItwoPux7631yLtE4NyyAAdC0f
IrZ02HMHTY8OwpYTQJQMJNn2m1MxKNKOzrtWvdqTgEax+bXNUFGgfdTIpiL+KeNk
Ku7xxKuC7li9zsU8KcpN8FFAwnI57VAYQtqOHqcsgippLDQrwfVQ3/WYD8sGnpUU
hQK6gEReqfDwCkr/ujh5UpqClBzQBc+uZm46VsosmAo0kYje6LQfCkRTj0fi7bfc
N7blkwjqBAGVKTvAHuZ8j+19jpeR1LFp5IzuxRjcYkGHwK3Uc507pX6hGvwfFGP7
kxdwi3YYbaqz9Ry00mtgFuFQhfCEG4ociBBsOQy3QqhfQnNW0GnsRDHMMdXwA6HS
hH6sef72H97uLbGHg6BcWSxUXRPw8gsyiT5AbcXvoyAOiXJJebNVjuAatICzsChs
jUD50oGbceJHgTLW4fX87n29nCBmEPdxtP3/3uFl6e99svqu0JdH9QVLtosZSV/3
vGOBxed3e+pKLTA5wBjZtJwMhpHWtmEWnlrJGW9LlTZpKzzuQh9+MjrqUhLLnFRq
VMy3eXqMdBrMe/j29aoURXNOr5GBJnWDEyKQZv0qeOOO23MPQsNw+xvOozW48VNu
bPNWxNZ7faKW6X+VmxKeF28qyVzEhgp+enxM3uQKkD/UaRcTRFiOkJfbNWy2lNi5
PARFxzIVhCNAmnQQzeZSjSIifsNQue/hWmzdbMX/fYCH8g+fYvYwb8f04DjKrjKJ
U9bj3HtQ+/HUZRlyvcnJq+l8msHLWcfOC0a45ELRdoaFYp/PSAiu8I0I6po3Yqth
JxqpdO3Blmi02YnxEI53CqLookPvb+s+tIb9V+edcrgwhqp6aryjs9txWymNZDfa
3jlHoadrRQhBDv6rPP5CDLw+qFRB5qgITH3RGHX52OpNQcDkV8ueKyjDfs5jegms
PnTScOTr+V5xAdnTKKrG3M5QEtx3+oovXIuLK2XSR/3YqSsdCbG8BdDXs/Iy2k9Q
84hmuk4WbJAYL4T7UtcnRa7U+rUWZCpA+E1V2yTiqoJ5uEljY1EQNl0k9ZuKEDEt
2AoVvdVdpOXITNXNsOoYdNTqHs4k/JbH1krvNBUTSPrv37LNSqrYBj5jwkd6JZMD
ahulHk7R4zZLkAGXJ5whc8cEc0Gh+g+kSS7XDmiuDn+I6ZGsricXvnp0zg4pGgBb
ivaqCWYgw4o32PjHhVdQgoxKmB+2KIF4WpxNOsbdUy7H7VdnjOGK5depKUWPeWkX
YVOqMBlNKt20RjSePKDqHN2aO55inL+dg6rWKBTBulYOHgov2piBaUCS4LgX8aEn
VdiARAgHPItOSpPVS6/xpM6NH8WS65cPdxMjJp8Txb5EEgUIsSvjFFztCu/j+Ric
88UGxf0NlMscvDHtttyZ9HaZBxIgiKyzfDbWEak2t5id28lvJJlZKyLU7SqNHZ2K
wprfO8eH3I8uKe8uRQLy2KGBjT+aOtgcrwFZPz9RXwhD6xPXdTYE3fVKPYTassjK
70AsmLgCRY5fD86nvbYHF6ad4eMrRFPPM0hKS2xFRropOrqYZOpA64IBNpA2TK/n
8AIPDjp1jdVw0yxsB3QUGusuvOSnfNcYOn7+fFo4M/QhOL3x2eYFAC5ZEcHdj/7t
VzzNafVjCWtSzy26SEE+jdkilQu51PMIJuBo7KtU3Lw6RqHMGaSneznxcEiu4RJQ
Cmyft2YLxCP3AU7E6bySrnH7+deZOFGKHlh+p1qcp9XAloHooMOxxJv0A3WZw0uy
sCqEh0xp0kqPjZfUknrY/i6WCH7BhyK/z3EF9jAs/6/ytvP/8ZVTmZOOiPjYP24M
ZRCtB4RsQKCYdaM5vk3HX+dOlGio98p7H5HSZgEE5vPp8dW4grELH0Wb4ovjnAd9
ZTXHEJDlq/c943hjQJGq6elHsehE3pS0pglnTS1tHKjAhfgIvjKaNYXBPlyHa22H
ShyCAixs3kNidtrFYCY4Lg7U2009ui3grDK1i1ba45jThmTAfoeurkOpQR84sGwV
DGnTQDYDhbNl2NUab2aVUdkJs8OaYhB4icj0IpJonvtwI3CLWWiMaVaxIQzRshUs
taQIHs5r1vvJbfJIOHC7mgGaHGv9pBLBJ+SSV2VEnp4kR8CaMFSjEXYw0bAS72rH
cQqkqsux1dW1f+npVGI9g+3DGegMk0i1nOFNz5VsG7PDng71/plo9DWtYJayN0TA
JJJwiDHWUzxx83HGkFind9bNtiMP6VGiPDo7gj+wy5GzGS/wheQArx+s15O3yBoe
mmtig8+MMmLLvKjEuhjifyfdblfJi0kCwVhbac8ftov2cM9WhJlJJsU1vk2fHMhj
xfSzgxyHeU2jOawGkYvRAH4qYsjmtP+Xmu0AS0sepuNh14BUz3w0KG0ct+JC/ca4
q4xERcJHX2pxUHDITQhkhPbuy3Pb6HI/Td0kGCZhpz2LUidFP9Zig/d3JREqxOPi
dqwYPL5OfKY2rU2jcgrFPZXyR6WH0iyxrus4FWCqSG/WT8qMc94ZMue6KVpH+VIX
WZCGyRfVKQJNDT5vPwPOnONZSHll/Ux+Mc2Yl8YmJv95KflXYnbW0X6Q60q9BJhR
/juBEHQPrzKrXIIDV21PJneQv+JecqjWBsl3gSGcjnOPFkH4okGyfbpqOV8BWl7D
2IrnM0tbUCNV4SZwx584GFJkYTNAbgpiFo0D26CgIZm8F30hCS2RFdG0ktx46QdH
cGYzwnEtIE6kOqbym8VdpUoqFEZYoYVgztU6bWbJ72xusu5fjTFHPYBJGkkA8eva
ZLraNqs0CdVpGFaae2n7NdWeMqh5Hgf4ftJ34z2oQWEa9YA+XuENFQ++TBg9Nlgd
2Rpw6qHHX7uX7W1k49qNOURWepoq99ZQFhpfdf6I2NEVoxID3FoHWIwiTihM77eD
gbZhdDUl93l6NuWyAgFU+wA9NvaWAGawdYOr3et/Auwnjjbiu5yhIK77LFy6H+eC
G84HPdTNt8qve0k2Bymr7KR8cCfEXTml1hDoZeeTcYiDtE3y0lj9YJsmHYF1Tqtl
Dxddk7Lbbc6mSyXUWQXN+ftmaV324qrDA1MwumDLRm83BecTlvIjVBrV2TqySMoI
EJelU2QfhhXSY5uuYcPTEGE1nWNU59A+MGAjCeaavZgVp/fRtiRqfbv87kgqo48x
JImdhHtdv9qBhd4pFc0wmVGmFfYal3Uow2s2821e/FbmNdz5NF5+n2H9hR3PFlNF
sElNJqVyD2aj5UCEjKcz1AxVNzOQwe0FojLtTrEhq2VmlCfTA4uoDHqRrm8Sl4Va
TFU3mHHlC+NkTU/RekCbh+UY0FiUvOlzxzMsNd1DAoaJX0BZAOKQyKy8Las1yFPP
aVHg5U97KZ56SAixNMJUU7VFwYOfqYD3aVWwQcJEXgVtcZ6nsQd1VQ45xV3FqXcX
4DGU5srtL0q4OqQYcnXaTOwHgAJ7ujv2gezhvl7feyoqnxlK7peB9z9qgFuk1ipJ
ba0xoICmwFdY3UoI0B71WgHtDhAM5tX/7UsWVO1AIrx1X36fWrfb8QtYHajXfhxM
HgZrJ92paAT7T+g0eyUmrN7ONaNqEyJXtB1X/dWft93RFw0KhEl0IPComaGzPTNa
RFLGrtALOQ2FWcDYQBFELV8L5VUGxZ4KRdGnqQd/Caxg79Jfjg6ERzf4X/y7saRH
o2P5FVA16u0sdHejTSjYPuGH+FGvhOAMr+9uzYZS7syJl87DYdx3Cf2bMRtnsd/O
39DiSAuk7aDm6uIOZYcuESFkjz9BPoUWya1oanfsfzouL+Je+zAb85CA02CPIKdV
A1XVXCY7NSWhZh/ezQVXIIoBVHg4eL3m2M3aoNMAMJaG+6byNFhzYBPGefARTx0m
6TnZc8E/TcS4Jyz5w2QdCBEEnDV+kMm9gvwXe6W68BK0sL3WFDO80gla8VsMG5J0
E1Vn5mL2f5u7dnmaxb+oaf/Yj3NznAlv+5b0RdfhEjLiHL4vn6tdU9rQzDsU1wbg
ymEG86IdQ73rjI4I5iSYWIHV7HeoppYhGhVGvth8OynaeIKuoyGa2CacuvinwEwn
ESFWPDeNow0nXpEBxKNu3QXA8FWYK5DuIa1SZgqJU42MtpORtfl2v0HjsEVwQDwM
F8i9dE+UzwoZPw4Q+apgEl9UlJTCDOh3vpRx5O9MBwGEW0OOMyFklGwlYt3nN0WY
qNLeYukOWyLTC8A9uCELCmzXpkRDvtjNcSUlPmZC2XQf1L1WYBP7TfnTd2hI5fYC
/CmbSR8ukS00rQMzmkWAwKBBhalFUYLYUT71h9u/ZXuG7oWE1x8xu1IkxvZMB3D7
XuMQpumdrol2x1Tpf/2PFlUecklHuyD9IYfAOWQMmynUnrXq31lv8vAOeY9qd37b
lsA89jGxSFf/tdnR0Cw2mwjb1O6hLxT0BsG3Xe0fWme8Ye04Yjfclt7q09h41Lut
LsS+evSgehnOZpf9rZWWNHOzDPp6Q14wNmglJOX4Hb+zeYCz/RaTEMQHSz3G30Hl
unQcsbBpC9ihXEMfxlr0WbYPoUchk0+PUgJ7fNnoO5HbGnp69KFbayg2AcD0EsPT
B0hx3wVN5V1czVKinS7iKRT651JXmDntg+ZeyvxRVSv1Bc7EJ2ebpNn2qBDADWlP
Jx11ySwzIfbn012sETurSvb2PAGE8IC1WIjGEsbLBoI5f5+GfXR35IrMmcE4ETcZ
pVcWyR8Neyv57DG2CxPgFdSGPwUJZgjpBmtFJKFQ4Y8RkmkoPcubFCY8BINdfIO3
vWM5p7CbNxPnGfdO9ZBMC4tII4FM1LIBzvyQtkuttVSoPKfRkoHzVHJff9eAMxJx
UWcTdBbJW4yQ4cFqLPIg82k7yJEZ+VPFXM3EEvaSbQu8QKsi6jCiN5RHDvAzdtUX
A7RDwuPURuaSQkVF1zUYy4+fDXXaCxTCq0zKAkH3+nHLiw6ph8cp2Okc+mT19s5+
uBvsJWT6P2PC8UexfyzINvPU3erhUw6z01m6lfnA4caJYbYhyWyXMS984H3Oe/nW
WryQAuiEpLKQoh+w/3ED9ySG6JWQ5VA9Uno8GoCCMb0yq0CXklGhzp4IJEWcdicu
0JTQL0urkn5PqxRuJ3aqrUbMvQfJDTBIwucuuK9UgFtqIN90PD4fPcziISmWgi+U
H/8F/cZCbaDYb1ifGqvJwId4mfn4DejU0kuYQXxD3V83HR1vz4XpbbM3VRarkK80
4fNRG7eSE01O0lc8emcPiielm84MehbRBLCFCj+uV3d6gGDQ8kLZz7+uFmOOmY1N
BEUlIjRPQ8015KYSWpA+83SjzGa+6429tjiSx3nmqd+M4hKbuAJag2fRMtpsJeje
U92c2UumJpvHwzrzSfmHUtBvoTTShrNNtOMvFI1jxSTQ2rdV+NLQXez6bRGbc9fg
QvzXGRkC3ieTwoxtAXXhP953rJO+sp6PPGnjBdbQg1+CtgRtDuxvo/Aqr2T2Qi0R
K0M5rHftgBJZSZ6IEqqdzD/Esd7vUWNmh62ZEkzp7ZhMYwIcYSJwN/NVzam+mXGM
S4tvsZefFBWuIV155PwbRpw8pbSDGamqy/9Mh63W9CCsFz9GUdbBLZGRTPGqYj+h
8KlBU2TbehTURt83YkDuwCTrkLOXzxOg+0v1k7hLWmarWZplPcpCoZEsK+dN0u4s
Y10GtzDOIrTmF95mnhwY0qkQyIjpYLzbVNJ6iiAuKn7eAjlbKvH7ztYWKY0qdXM7
pUsm4cemYTSad/FHHX5aYjorWXY4E8jsQf+5kjebys1tpf9NBV4kRQg7loydIGwk
IqGcZNFjsk84F5yGiIXoQAggGBEMqxG8SF7oNwNuXFeVqoA0T8J11dp5ALmpJKI5
azhlgm1prz9A+3wikUcve+CdIiRTutVUnfOR+gKnQP3dpNpc3tufQkPcCuSuJgen
+996gNQpU6u2Emw9mBTkAuecjM1uZaC4s2n3UAqW81u6yQJ2RazaCpIy58nXUIno
TvPP2BmCxOfEmgmcWGuPxZU7S1cBQelxYtxWY8sdve1itLPfaEPPdzn7jNi58QMs
uVPemQJzCMjLIJnXOhf7qX24e8xlhs+dT09mV7isu207s8fT9aESCoS+993CBKKb
FWcwUsGMY+kGYXGTmZk7E4yxWGq63qir7D4UssMBtMV8zkZis0EyyUvNmeDXs7Ux
c9c21ZS5EKy8k0CuRppB7n6A45uvXimM6oo3OT/8OcDcGMrF/O5GAoOQ3CWeU9c6
5GHex8w9qsf+O9CQ4ZUyv0/kxZLDEHsT3aCwAhyI9sGNAMfmigA1PzDutX1MIwhD
BLJq6bjwVZnN/pCKhjkq9RiPH4n0nU9oJXiRkS1sLKzl08V8NjoJMRVhjo+YFe44
akZmwKSp+94YYsMve5SUZ5oM0c+v1FNkBOWalEaJ3zqK7upNjjl+UO0wkTo/dZre
THMJ1cuSdWr4+DJNn2UxRS6m6aqcIijErYfbjF3J5xLcMCxUbKUfY+DcyIFjf6Xb
GqKaIcvbaLmpzBZJ47sGdV8bxDyfx1PgGMsBAKMVQW9urIDwimULgyoxvX8XPhfl
C/zZl9x1daB7dYdBjhP0cNH34ubQzArUAjhW/R1rn6nFJcmauXjEg3au7G7gLlDO
8H/eZ1q2zgrMaZkRD+qssBH4nZb9HaRZUEMsxR60Ccd8+dDTJ4vmcAidDgFEwtcb
iQSq/ak/GR9in7MUDw0nnEeLjeIM0JWhpwdbNvMlbrcbe2bEAQhmqgQfc4iic9YN
WctbNIQAx3rPc0HMH/WU1wzDFYEroLRukngDs1gZ/zuLOdKm/D+byMQ8psphTX69
LM3O3obD1sMY6RYh15LWtEXAlWv0dk09qD5/K0W2bAA2PCh/tvUvT9gNueTGLDlr
5FOYWEvuVIcGbutZdWYac2EOpl7ru464GtwWnEbQy9pvuyiK1zf0rQa5/aAqdM1Q
XJLo4ozTC5WexXx21gXa094li+P9chEk2a0SNcoDva2i2R4PcEA82tWWj1qCw7dd
IZeFo9D+EToSqUsFD9l0Q+VGYvhLFDKq6rU7hulDlr4vuSu1xYAqlESpeWC1ZEEf
jj0SHPPZijXlsKWC8s86dGLHYBr+BOASbMynFV9Qjfq1mA4luIXIYX/oNnc6j9bV
uq+utU3G6nYIQmiVMNNCpYzTqPnEDLZJB1FKUP2nRIsN8aax4jCe2lJEYJTbmXtN
dbvVsDczBau+gvgS77KbNbhOeREA8TdR6Od+88mtbXmED/+FJ6qFx18Lc2KxeIro
18s87oqu48Za0xpFvxvVH6vATa2Yz/VmjXglnIV6++OLwgnh0COv9aEbd7tn9SZ4
CDXnOZxks5uZsPO1iGTSJJlj+MxRcNe/MF3NipHBL/N7JY4Of0N9JbHwLv3U0AzR
LzNM3sAVPHRgtzjxH0Q3lEsdfB5tIXtJfGCOdbyfH+6J/aOZU3AACI+7OMQN5Cmw
dglbEZHJzR5iyTX++DXseFz7Jl+ByZztGYbrvU5+jbxSGRyFeqqtQbAqRvemxLn0
/DUSgxtSAuOJEmpRdXKfbmxq54r61bKE8etjUFXbWKDoS6V0CpbLCthczPJTZYX3
d+YZMUKIfrqQjYJ8fbv12xTXdKYk2FphA0X5eJEKRmwVM6PykUche6jZqimi+R0R
Tc0i6EEyniBKdt2sGgKOWvE0e5tJb1v9UkzPww6rwlazmAFEhHnf1YMvBk9q5ucW
o6NRcUD2/Q0OB9njjzT0k/3xY+3D9HZt73xd/pYCwMtJw/qFiPpsFTZSk09a7Ibc
HcX5C8Osc3s6ug1a0EFeVztIO3n+c/tBAYQDehpMkOS/mpCp5qeFUCY9uz9dCqOE
PEpVrNFK4TuCoL81K+BCuScYG9xlONKsdYk2wgPJQpBFlV+d9gfMBhSGmWIhTuUS
tRJGUjv/yllaYs0iE1X0K7DePumGL8mZNYQVkzBP3FDx1WiSozb1qKKvlKEHYk3j
gZUhhGNhjqsbbB3oypKcvNuzie0KSw3ci7bhh7rd8YwhJahFFL5rNXAw5kAUtlZc
0caTj4AUmSYlsnCI4nBPegx/ECZY+W6hCnaOsvan3I1iNUelEfGjR+EOjeltygk8
f0D3WmV4OeI8vAlNrEgbmehl+70ewwMOPYuLLkHtanDajDSTfuzufFSFLfVkyt2T
C/45geo+hZ1zR/Iol4fx7Dxm7gsYtFMxOAN5Qr85MtRBQwfxJUFn3qrhORzPfflx
LfG3uDkB4kWlsweXMd0yAbkpxLmeCvV2+T3R81RwZgZFa7qDHnvLqbYnSyHyV1jc
GISLFYCSh0JRkUo9ygB5BqOcY9Cqzk4r6DCnC1mPB1UpXl8ateJrClVcVXMEoXpM
546CxUfnlw6MEdxejyR0Z7GGhSYNe84kVQ1i4mh1nfy+2myowbIvDRWxECjCmewY
HmBukvgQ91XQxxBa8dAJLsITyM2vKWyo5JRn4dAAW2SIwDKE43jreF9hgierpz6N
YkpeZMIoNG5S8WYUsgIkIKGYQtIP8iz6IcTggt6bqPQhP/VowFSZJ3mbuSQxVH0E
0niRWzEwsma2Cc4V8ig48iB6vTVM76yXU5dKtJFTvM2+nRjdNjGsMxr2hod3KetW
cv8kSvaA/D1PrVDkQD3p5MRBYs6aMnksP28GrvIg+o1/xw/gXFxi/fz3ditCIViX
fnyJmasuLh7Hjxd9xmuP3cJfHhN0sOBB58Oz4ZZO8Z8VABORJ7GVlMPJ/5p1KTLR
su8RBOvD2qnPBMdRjFIGTihAC77gK3VoT8txZpI9XR/V5AbjjTeKriV1cRSUnmxg
0rRVs94S+KVzpOYz7cbW5JGr3YmTg7hSj8QlmOLm8eUhWf91Z/lsz+Ov4+jPW+hY
rR7NoAUbQTgEHRYZwTKAoTNEftR0pdaboz+3JgzHcvU5Ydl+dt3HawVIwJD10MS8
MyJJ4gbcr6vdX86ZanKaeySaYsAHrD77CmertaMpMg4to+x9PO14+G1CW3Uw/+Cg
sfQoEHiUgHSLPA2/rtnwHkztRKBKo/vPgsCxftVE91JuCMcDiok8Ssuox22wiDmJ
rZHV3ZNCH2TUTcmj7fxclhz5CFn4wqUN32lElpivU0J+XADCLUaVXwH201ek9UZU
f1aiNppFI2m5bcAg/vhntVq/OfWSy3PcLb52LK4HY6Pw/EvmkeztPuou8eG0TVQB
wD3PxLvNKI3uW+CImlPqgOd34AbYzPk/ydcdgCIMx2Df/F1DrNgZ4pamVcGnC57w
XUhw3CPU30DdrM5TgWjJLCetefmMq60dAjKlu8RQY9AOaTTGgEWq3VcuQZrwkEQz
3WvWJMKXmIRFXSOpPZI/4AfHK38GsgidZncyBNTDffXI5QrlqymlVXLrrE2IJS0l
/wC6PvW30uLkPfhcbX+50+ESDE8b7+6PTj7eSPqyoTJHoFR52qmpZcZdYfPcOd3q
Veuiorfz/6QwR/GO2gdkufb1ZqqXsTQ6DyDgLyf5/A9WZHl/NSviXtgWHgBAD0TS
QxBcs6hftXg8bC27vDKB6RNJELnh3yB8lJbIo5lbvUnQeRmylj//mafhx4fR7kyj
ueWEyyT8AFI8DPuxf1Yq5zubV8yKcANqOWrj9dfnmPyy0Hom9vgOPInKrhSqNIkw
xL7ylDBIf8E+4x7FHCIJwpCAzdiKrck3IRyuZQw+mBemL3PFvMcUfGVS4A9Nvxao
QD/5g5AlDzbSCTCGHxnqH/f0NDNVal5bGg6UCBnFyH++B48uV358J5X2Rgc4k0ME
5kRRW4DXwwwdNDA5JVX67PxDouK222Pncuncjm+qeh1GYqiIELZY+mvOBoXTG78w
GIw8/VHrKPZbHW01t9jDT2wYQiDXNHRs/LQYKf0o2PoCO89/8dcxGNWdw0sN0xRV
v5BaBXIvtV9DGv6NP+b/rvyN972JGJQPbsW2eWdhCrjh9lYr86hTiJOa35k60Tfj
AlHBptwybSZ27jC4PuAYR4F6N61FoeNL7afz4AIureNU2r8eLyTESGinsjxewGqT
9+lAevLYJL3ScdT2d8+wEq4kX9Jsu6HckX/zgld8kBECAi6ejzX2V5aIpX/Zs6oC
EAg+o1VeogeCzn1RK5S0PqKQLgvKZ+x1PHLCW7b6sOZeigfgb7qWWwpbyLsNOYMf
ysgN0sRuz6lKx8YCXU7r5GM/j2MYeteCnHFz2ROySZtzLiXqOZXbFZBDGdw1Sqpb
o8mukIo3rTFY7/IL9jH/cBw1o4/v+GaurVyU1+Tv9bEXkOGmqq9WVze6GbHMOEcA
zRyDwz6SktqFYTJvZqyv832v7ppwbOpG73wym1BLCUuvYkcmny6WTFgSed7WmjaC
b35BJih1a+AjwxiTpfqxYoYVHQV9uFsApFErNIhWGBviM5t1OxvqXVxrD8KYDHQJ
jZFByl21PqlzBxnptIzjviSBffzlBP7Q0xqLSzuzq0xzJooRoQrOS+8qDOHQEzAr
RfRIt05yxvIRlL3+GQnxKUdJmOYo8jUBT62z6CRc5V1cl96LMUYAvqkHnwA6UKN0
YBPEHgKM8ITSkRZI/YzZelHdo8q1Zu0h3u7mDkVeaaNXMbO/+IGa+EiFoRe75gVj
lQca7SOr643ysC1bVLJ7gWZs4CtKRjawbEJWfbty4u194BFBfokufMI++uY29VL9
VsD4kakQ8XaqdinzmXkGErLmpacQp7NmzugSPW81yn+Ki8FKFFOBsMgVt3fotomB
dS1xhu1lC78aYZJfzKyX8WbhU5/MbKgZRc1Z12hiYh6V9JkdzTszZVvW+Blmx1k0
nhuyuwdL4d18e5Ov0PgM7NLRA8Y3SuWj9442DdrTcU6etQEATVcfB7PPwWQ47HxU
r9t6GxuzQFqiElEO4rRDAaDSFF6xInj2RAeeKhze6tGEbYUtUexIYuwl4SDh6KI4
dyWMyUoFfZ13RSC8lAdSJ+pKRO6NpV3/gQeVPlx2wC5IbJkZBuwk0tSYXaSZJAWs
hY1obFaCiD2D4+Ms9bJCGOEkh9H2mlhmJ8sMufnzFKrd2JP/fsLgjnAsWGpQKlSD
F6o0ZFHjSVMc7UczxMFqN4UFY1RiLJ0fCdsefACbk64PwSjKDb1gZXUzGK4EEg/I
cZmbQt1NOhbZYdn1kSmea9oERL94O+WPOODjX0dMJqD+Ahvb1+W8q/7QA4KkQcE8
rJCtFWAlfcXJ4s08rUsMq6DOXGHsPQpJCsxuejgHaGSE+3Ol++LOEFj9st/ptOqN
jVJKBvriqo8oX6tucXNJfsIkoxtmo9+elSUNuYW7mwD2J+RwTkQEJB3HQW8vLO5f
N0iw72BVPI8Y4pBlNuTEgnTB4PCUUqxdWvGfDfr0Xc9tf5YFNpi+Fn5Kuau7b5gc
vPVji4u++1qUKKSUKoO9Notm4LK6BDXbMKlSVpOJdTjcaMSlgPchdtbzREhR4xo4
zbHQsxE0QrqzktzJun4NFbYxqrs+XLUG1yQwdUQ/B/NMUkBtiCnjuROF1DPETt0u
Roc9sit20z9tQjpZK9ZLFv/oGN3D742ETDXwkMAlMrpgOSpn0vabFTb6q6BNmwNU
wNZ2Ycx0talkDYnlrJPAqkNp/DQbo+B00S/jK1mImwR5Y0ToOiJ94H0bJZzAKsRu
PEB5KOg8N4Sh+MOmfav0Wy4OzUlyq4Rx2+IBGmB5A4LEpt62YzCMBpxmXyDM5IWR
ZP9knbyu7CSjbeqEYQc6DyO8RoOD4jzD04HEu00OvK2byJOogH8QZnc4shaFTkKM
f2lWQadyMnXcWfyA+0qvprLe7wRpZWhTrgBkl4RVjkZxGKV7NTqcTiTxHoMd15FL
kabtj0fkW6NmktSXOz5kYTLIglLnWGP+SSZeoKxMMiGeh7XKE+v4+cGIr9mIsOhD
slGiIdmahMk+nKZK2185B+xaFlm0TfDloxNcnDmzplOxJ1vtM7z77Mh8Eb+8zdUE
Bx7FT4E6+QQ6Sx7K0tFe8SfOZCMoyvpuBGBRPCJjhha26efKqAaBw34FEyic1ZFX
xtyPjoekXjufY1gMeRSHvjM+mX/qcfa49KnARan7GTHwS3KGm4t+c1qzlBbQvguD
WkjK7pQhW53UhQX3TKkRvTPL/ydQ/klspw8i6Hx2bXsTVQUxb0ywvFFOrQZgyF+Y
4Bi10DtOUnI5vw0esrqzrqI5tMSdmkbiZnO74xbSSOpLXDle/isfrumUw9TYc6Kp
auEpqNo07/40R08Kj9ou2H+4umw0FxtxdLNG1CTGEr/RSK7Mi4+DcJIWB07KF/Ki
Od4iaX65k3duqBCdA3xFC3Id6gLn7fNTGSe7+pDzH79CDPDN/+Rc/hw+5sDVSusT
uqgaPBDh1MN2QgRPJ1/3FjTKyxeqQsJqyaNbr4bv+H7zswZ+BOHNKkP5XYJ/hH7X
b50yQCj8cNRarTKxeqXAdg4H/c/SRV0YVP94JW+wK82EnlLcedRrdJNM11nIJbAO
Y989Hht3Aq/XVZo6K3M1/U8Y4GEcgV8WZ0X2PXe4f1jdULa1GDeLmw04OWWosyFZ
xHo/MWL66/u5STarZYVpJIFK32XDnjItuF1PZUXBspHvn8blBq9qp7gpm7rzfCHs
82Z69fB1CMMSBnxaZyIBnXiU0yIgXsPN6koDXBcLUR9qaEWgwnibVwTOZurZwae/
6c0Car8UNaqFjKX65ZjTlhccbKDOg4Fw3W3GrrohnCb2TuMu1YRSvj0bHFg+KHPC
GoWe2e08rdMXX7Jdw6VGxIJDN4eSmAkb3L//EgHVmxebiSift7PyMTeT6AmzJjBz
M9MvE/kxd5T9a0ylrm4EKp9Xd5fczi6cC00Ix6T3r+cQMmAEhTE02TjVhn7Wyw5v
YAzpFF87nHXPJ2bRL+jv77TTf1zaeppjPD3ngSxkuo3TXWV09soprNo8Ljwq2NSl
SADK8OPQoSX51DCPgdCj2WycZ7Dzdkk8B+CQ6ZV43Qb3HU/mJHatifkLljrby122
IlKsMKtMLae+W4eMc+kisXFkvEgBElvVHYSA33LYig1Mo5AwAhIH/KZJbc0eB2YO
dVvmct8yMbKKDqInFn+CCPdZgcreu25akrKYwKilh/taDl0R9v6AsLngC0CM8Ahd
/n5zYN6rm5Ih3UDyieazU36sjmhcnykfXyaqfm733EJ71PGzmfoDB1EVp36lgXzk
+4+x6AYXjFjGAD5AfQRpWgWQORNAkwHiMEB6rwy9aeq18h3CqfVMJ9Y0B0WZQCRb
QwrjY7hvBpsL2H1KUaMnrEXf0MsuAfVyjIynsS7OL2LOLxzilS67r7h69LuR6AIZ
/XhMTG8/0iAyHgWSmLNc4mlevrhh5kuThhyg+kPxg+bmZarZKERbDi+4dop66VhD
u05U7npkPdOJvL3JSsY03IWeMzB+Fbuu4E33Div7cjkmY+IGhdK4RvI5b569ecKd
AVJs+cuQkbnvsOYSXMJ6ZzNyis0wp0fU3d66hamqxAYEiOjclV7YajLemYuFOihc
TaPXSkkkQo784SS1/xrpoGDtmah7BGBKeLTW/+WhpUiTqYdxy7U7xetjC6B7cO9p
plyZj8nHx6R8aSe2P1Td0eXoYRk++nuPEyfL7dvC05hXsBWmYu0ZbGZy3Ip8U+0L
Z2kGofDcvquonaWULq+vlD+FjqqfUMak2VgBZmWUN3OnKgE8kY7qUBwXCLLFDtHs
oIC6speEQ6ERzO+hLh17XGoWlzWs9dAkcfYCclIjt0n+PzumNoJqvo0DAiMq+VPJ
Y5YeAL7WaDZSI66W9BRZReAo+aD4o8bizjv487hRdamk9mVx3yIYxksFYzMQWASB
IqgyljxF5CkWZhTBw+vt2d0ajFybNHSdUVLtEAms31lJpR+TY8HQKNHEWDbsfPFQ
xXdDPYyNJFlbm9sje9lISsTBthf5oRhRbG33Mop7+e+70VTMKsrmbs6L0f0ikMb8
RbsBCC6rnA+WETev4XXH8jAbi5nwZI2tkmrpak63DT8++oBQsj6YaFWoP1lMbIjz
v1sufm12MOhENTDpaW/1cOAOm00qS2yO4rxpV5jIE4KHB5csKR/ymAvSvboDPZz4
o1Wwg6dLhaeooQ5wGut0Rg75g9D/nBaV/AA2XTauIV5SfNasNPSRJHkKZyzfimp/
tpagf+lFC508IZ7R2QJ0BKCDvIqRi7CJslggbA+/fvBe8m8gQiWEGXRWUrLIr4ep
ctG6IEg9kBh1I8yqFoiGqk83XIcvrvLymuljJUonw1TU9xgHyP3Pc974gK8qbd0R
kC3JoOv5hRJwPLTbE4TS/CKQg3H/Zc3Ybtryj5lRXAzJbMF0ybR37UDL7Ixzqnzx
mH+XQiRdoy0CMmGiD1IUclusxW2VuXyMWTP+vboWapJe/rt5dvhc2SpiLlz4hjDI
85Jm6ZZ6wMhq/y8Avy7yUrakVacNSc5hPwan9FsbAekWSnv234iuePiT6EdrhRDI
fkxmijSZr0PzN76rbPZ3N34OBy3TTfmO2FlPJYNn+tyuW274eWf6YCXff5egBFZ9
Mb9hESHXdF6vbaRxITp2HNzMiJHCrM3+08CHUDlTKi83yYLu/YyBUgzam0aFqDTh
LeaCL7zfz+zwDnlG2PKpKxq2F//53F/YvNml8IrfyX90MdwSur3V10GVAaM+qSxj
ur86tXWucqZzHbizlYT6chMMUCc27KQxUNlg1UTVn/6sdhfL4xZvWDk0wDAxPQct
49uKi3fLkt/YN8VNsrQfaRwvpiP4jrIRL2xrLt1kbSlqrCi6flFjyal+k7/9Ur/5
ZCNVrjcV7OmdVByH+HQWozlDrRhjo2pTvTJnb08OgiMpsS4B5yITg0WNvOWsYb6I
n0tHBKPGFxFBgnLzARyHW7kaplAoAxA3D8X8DVDQnHTTlFPmhrEJsmiYtCWnvZpG
W1qqfXh/PPdiFdZqGyC1wAMPG3ljRnrslCUPxsbSl4K5EtO7MVni9QKVtgjeIQJK
Ai7DzQztwT5+JKeLIVo1BWhTCVgmwvbkuOz92VHzTqTNM23CjcYGZTPb7KLhUA99
BfQJce/036CPwPZATWY80dZguz+IWXSs7onxlpCtTEKVtE9NUCxi73y/OktkwIEW
SKbzrUCC5UsaXFG58clFiEGdgd0RN0nhzLXJ2Vhm6mxZYrVEjDxkbKZCQuDEW2Bx
/qusO7fhl6+k7QZn1xZlkVTyp530/bnhgMbQ6jDu9/xykM8NzKFfsC8+a6b/suX8
hg5DLNxK4OblVfyFrD4xja4fAwBTR/7LIKJxvJ2K2Z2hM/1C8cVME4NyfjUBZugO
mmmHJHM2evZuURTqHJVJKCtRNWtRZFJavOA2au5qkioEgPVp5jsH8iiiHCkcWsMa
ZtoCJub5pGQiQ2yE5XxpleFvDJvdo6tEc6lITfgxMSkR1CqHhvl03MF0QismoCS6
SgKD5UbWrTgjZvVxVff5RpAlrq/J1+H/dZszmcoubwF9to3cFET+VkyRxm4zkAsz
QuJi3FKi69OEl5Kg5rmKZAPLyWjJTNmbK4GAW8JJr10UBTL9mOUoLrcfEfKXCDwM
HkXGp3ZyEjnemh+cnRi21MVFQP1M9nOoaNaf2KhS1FJcvyk2a25W5ELf8QHkKHDV
UBD6Xtd3o0md89lV6VcDbrG1FOkz5+9k2HNNp1FYz79tYu7DxxN53Jbi4PsPRYy3
oPS5ew+fnjtI9jQrz1Bu4s+h5gtok8vDa+V46gQMEJNQ6fjqPO9eXDRrxhMu6lQ5
QCC5cD8Rx17SnB0WuNCLoCTXJzxK6N7r4cjn5o7jiDsTo5Lln+KNETQoK4ASb+qz
AzGbtQTZ24UmiyQlBASqaEwbFpcNeipGkvrsTLi9aLpahOvnMOnbS6/PhBdoaPt5
jMR8EGVw+4Vi0hQoi59E/zlG1qhlkd3bZrG4h09dsTC9qf08l+xb5HdAHqmovpnk
sgGybvMxLGKybMAWtbHqVlBOS3/tt/i0c/a5+nyZjP4StQ9nymKBNj19wJHNMgQg
Ag2Erw8kuaIXPstMUny0Ifz0IOMumB7/YRUKB6/3ZW7bEV2C30r9LPE2ijoHNRPU
jw4QtCpKKkoVYWp8LCOw82rDz8h/lPi+x82SkuzEpAxR21+p5x1Tj9mO1/8Q7U3C
Ku1hV3/UM/7SUtzQM2KvNPMs6ewPcD+JqVHSgO2eY/gZAXRlVmT0WyAk0VKh48AY
2Eit21QfC5XkodyaBPjehU26h9BF6BBD3eYzbFT3TOOLIXX+GRUll1MvtPOQ0vT7
0n5rufqdP83mVxKgAKdVnMjHKKNz8ZNnW/lNZzuoI0Jh04NJJIf8nYNyZrokoYyu
cIInNoqL3wzs3g7qfwgpkiX8BbosCmBwIrJ2SzMLw761A26AuvZybQU49zRMMuMJ
FNn0XVduVu2RGsyNtLOgMXCBgjvZ5yzGGUBPSp7PB15QnJDuJ0bEt0izjolbaZ2i
KNUYxgai5O/J8bxItkwOhf4jpHgsVKu9YuTK2uf4OdS9UCwwUvUlUXuT5i6FUMwS
/mBGfErB1ybUc09KDi6QDWYQPNkw2OJXwcjR4BFl0TfcFbGUM3tkfs59/va4Dhw7
iUpgv7k6Y/5zWUWLQ+2I4b08YIhHunR1EIbHQ+SGJV+j2YMwCbi+aanCuNfDeZCl
+qvtgGr+6J9ewRXeFTPe68uWeHfeNenBb2Q4fbxV+soIyD8R9BORlzzM72e92irq
r3w2lPjrkh7uQJPaUCVOd0rPKm60TrS119ptseLoUdI5fiCvTUq2DauBpzNd++8/
PrwK9re/kdl97PpxOd3waR4V/k/Io/eCn3Eo2fxLW/nTMLYe2sdTokLpRbaSVHje
+B0GT5wNJyAH0ZLG/G6BWrGVgU7tXeS4wOq2Hjb/X+QGwcrZ4Ncj+py8u2wLGaKx
0d6p4c4EmifiY8Ql4knBjs6hmM4tC1zxONAlAbsvhqUYrHd3m7eHiyaEdGhS7JtQ
C7A0okVknbBdKczCSOgDc8U5q8PwSc8tn/XDgTwMC9EkIy11qmBP8Y6TaEAS+Owd
dDJNcr5XBXR1L0IlPcAnOAs7/GmXWPd7EaWUtocJjVOs8VKVhGt+pVpH0/5OvN6c
AZlZ+OxrHhGyWEn6JIV4T8Y8aTU95Ej789J31TK5C9OT0JpTMCzliA+gFzW/OtSg
hqyRlU0zySXMUQbSpPI0ogCxN0CygXV3igVkexrFB2ZxzrRPwlS2ju0u5ttP1agb
rSCV+VKG6g2hXnjFfC6EUvIG8z4bFivugtSvxE/jZdAABzgBX4RIWdZCQSYAs7OF
qhLGNDV+IWlG2dX2NgTiyC2XRQxqq2ZQiiyC93MoiHM0P4ByNFenT/FTfYHFy/Fe
kMD7KmfWl8nSRx8Ofm8zCGLEA7mjIHavU0P88297gGMMoVxZqMiMUge+/x5WAYfQ
bLQhQSp0RZzDzKiFRPd6rJuMo+Q6uqwzkzKLubGsXHI9zZ99Dij3BmJXowG3iSay
JYONQN9pz4jBd+IJ9V9kZnkGKQgHK2JFUsh98iK2z5JyCqskfrggZAdrpqwi+BRx
MnwOG64FE7WxDH0oyBVETPDAKIoe4LINjqjshPU0uSkJiBsfcHk7Ql+x4M5SNgMV
sfLZd4t1YECmX4AdD8Qk92Ly0SCTj3Irn6rDh/Ro1r1QT2BKvmlebzggR79DUu+C
HkDt1YGz3CGICWs5GFz7oVvZD47BJKQzgJ9+KMqsvCvyOnaW+I1gCVGC6/mq1/Bu
ptqAXondRhKTjdCCQFS6o8t3WK39vo8u+sq/gyDCZl0RXHo24BQ6LA3EavzuM/7Z
Xm/YxCerKxommhhm+5ANPkeYCcp9SlSaNYCk6UelSNvDBbhhu//oiiOxSAKfENPl
/JVliKTILmPQ8E8fUlsAfVxxyWytilV+DxSp3AYW4aS32g/WxLNOHjNvlAqvrdrH
FLg0k/iiOb7y6iS7FYLrwJwD8J+8CJm+HHm9c+2607TCbJOA5alujKxdRyZEXrrP
3ofOsMLBGUN4YU9oDk5+OpgO4/WCIf8SokArCQn664Ys6TYtdB5N8bJNxLtONRxI
8H6dE4k6cOqCFPJjuN3/NnwtnnYvItq//7ybe80yaCtfuT98ZYrK9y5eO/nITpnd
kgYSwZX/ohyf/YOn5pfcQcwKbwkhwEiZBtlwZTYArkIJ9kxWajPDcAt2T0AiEo1j
u0pBw4HVHz1KF90CgFe8xR4x/eehJsBUxye1kDN5cbyDIjrDm+bnc3HOXInVvRPj
aDxULjLieZR9LbTfcp0RiQqVleJBu6KXxpgCA0G0WzdTSUpVyRUsLwILb5mcMevj
3LxGdW1whyPXouY84G8M4wEypN/qOLFFImlMVg9lxl8qpjMzU9wyLb28IcXwwOAH
2trmf1pKAKjyeeTdjH0DPOE1O7ujDgCgpCN1X99o2OVxFJrUbpTbD6qHSADQSc+Y
Xmy+4VJOo0BXmJ0FuxI33c/YxNlyp3Dcw3wITu2Ca07ZloHlnLR/oqvq8Dfh/Rsq
MLQg4CCG4Q9d+Gko8ACbYR0br6X6+QJlAB4ncPeGPxSVHn954bMuo+nopaZL24Vv
6L27Ih25e0ggTuu0fX2jnuNK7sEMl45raA6GA/ACXhrboxgNJDuHzBX1A/kiCmwS
Q3ccban77pthQs51TU1h0K60MWvnWURqT/NWW7N/Ld2W5c20+Ir4sasSUVk2pXYF
Hx3r7j6PZxUjstHmVs3a5UdYMDkbagGCO+1V0IASQmcebZK9+0zwMRxPt7F82Fmg
xxmH+HE6A4CEme/3KWqoD8mKd6il8zPd8/NbW8zQfFroCnSYeDmn0vkkGijthlQG
IJQg7J/QlYtvMN+cspr7RB9x0DPSWz08FPWCw2SpJFN021pmwheLh4UivSgAh/hP
unt06C+6BmlHyNutWtsSxS3AocLpet+C6ssJLghQd4kY2nTcGFNJCm1ZJjh/jztA
NGOAckTDAnQ0IS2kN/wL9JwWX0OG5t0JJewyeEefC8kUAazg6YQF1XLYY8dbVxmA
sfyVt3D77CU/jX9IwgafUhNcgnK+UAj56vhXn4clO1Wx5aC8VxgT92TUQUUWKN33
BU7peNzriPloVRenWcG/k7Cz+8MOWC4nlMsEvbUv2t20XJ/OOMAqtkUuh+5ZIZ52
FGcHDTlQEv5qdfX0a35nTjMNBnFEH174ysjYsgYTSFY7MsoaUwxOzQCkd6PjqNW0
dh/541I3EN2b6ilN3rFJNZ8tQthjaZrTur61TXbAhLH3BvxtYOFjyJlMoRwnG3To
bvY3EYseG18ODlfPcPshQgFd+5DCm+WwHZO//HRu7d6CCLHOEmGiFvru6cLxtuJp
dq1yChHaBEzbJpjNLzlUAAPMPfZPAxdk0xBuRtDPNQBWJRtEleZjGtHdekl+NVp6
QJKgHTA6yCB8Fp0EhU839A3v+TUomgqlzle88jhsUk6VjyV/AqLPR6qxy5AOq0cF
k9Bt8m0kNQLj5KyAf7qEd6eq8ex2zkzJKzSk44FAUtacg/uP/oBc8Vac543j2uDc
Mo2u+4bGGLRPS41jw1qd17OUHlPG8zFRhcnzk1SZtoha52B5/z3pnnCkcbXN4jGg
DkAYHXfFrHQazDU2xU39jz5g12BXi1E5s8LZ9pnbOnusJsOLQCbC/J1HFJ8/grto
HnFLcTG3PLKc5zE9geiqq1Bp5FYiExHRL2JYut1Lcv5eTuUPagvljHsMS+82DF9p
QbbA+N1H16CtjcF7dczEKU4XvHmL9kvVppM7BhmIM3aEgmn5CcWkBapQf+NrcHzn
KujvHEBMj1FOSw6hxpWzsl0k/JjlTpE1qQy9GR32fpPcpuOYCv+qd8KEsRSMmM2p
diM4R+GbVGCvL2ePCIvxEqCJxpMbsWbuwSrreXUFZN19jr0s/EBORtASsRxlt4KT
zdjyg76b3sjxEtjHeWAJcYmInRe2xh4njaaWYf77ZEl2rtAbnC21joISueTFEc2V
1TXbN5KLoZlfBFLaU5E8o9togxWafElnYJlyVWMmB3/pCGrml61rzb4mU/41Lyjt
OcQtAUcAqFdI1ywJAKncnmnh/6heI5B+/BXuGjJmK4SQvZ2cxDc5XPJgGwjFTikv
bYhz4dwWG8g4sG7/BZupK/1nFbEmghyBRnB+1V9UOSW9Z1GqyQVebUB1h6cB7vt8
8kPYWo3s2ZBs0dIdp8kfszozNnqCsW4UWl+vBIChpQnnWQ588XClgZEyjz/Cfs68
+QECYmibUSMW+gXwPBjLn0KkKF8iYGn7XUj/w0Kw0YB2D2jENVqGW6m0+TYfMQvr
6nd1jwWLRtHWUhjUguiDSuqFyGT8AZ63HlWzQhx9XTcpDYvDvCru/u7Bsgi/u2ZO
1NI2YDXmGjmvhzwx6k1BC5Pdxgtsupm1ydxEQMwwvhee0Pz/7z5WSRvcjbwuQm12
U0ru4XKwIJBUUUaxFE8D0jYzY+1rq7pM2ikdcsr39PzXmjG32EwxtO9f+BHBymfI
xSj2p481RZsHJcBbazmhJ5kjtnLFta38e9bbgJx4uNvzH9G2j6niP1YCOv45305T
PmkCuzXcGnUH8xl1SgPncpACwsmITaOX50QOM74ErJBvPf0Oob3JYr7lKDPjishH
iwGCP4rb6wdvLO7XlbJ4ECpUPaxmb0/Yscq1qMzXAltfodFsNYWVo6q+jxk05D0D
BuaW7S4IDfEWfTeZ7DI7bI7dK6XSvW9ndujJSmZZ8wwnbnHMcYkMHGCc4cDYCI/O
RcauqmVGJ32T5/lTY+4zkgLDMRHA97uFFH2zVlbSzG6siz/+8zce+90fNhuXiTw4
G7UiQbUJBYKkfr36ValquQafmv59PvF/kG0uuR+w4jTFcNVSFR03iUB7vylIZMc6
SjBHfuw+k3yjH1bpzBWiTgzzvAeJ2e2upXOqpO0u2lL9S0k9FH+wRb7S5ydWcvwv
M+Z5JF/Qw3qXsSLnsPxy4Vhycrgi+r70OV6819Y1PZScM1JS+CV4zRMqXj6Uo1rI
5FgyV+RpLwWlxchUn+Wl7O9NOhEPry89k0JZQDjJXjx0BPtYChWtGllNsAMze2Gg
VpENCEKFyft+uFaLjI3huWnmhbbcvV4s08SKfzoXaoPhBE6k2dKq/LU5qqtypY9J
4O/s/l50BtQoSp4fMrdSYiixokeL1wOKs982WbG48O2Ea11jZlqBLqYqF3XfgWdM
qkAu8qfZeOL8EU6bHkQxJAJRVmNfGvcGKMw/clX0o9/rr1vD4zO6jy9ljiynZ8BF
QJQKwb7WVdDklPpYmVPWH54VcTypj2EtLVnFRyshkyI3CAMtBGa82wbLC6tzx2hC
EPAll78KSIXEB5wWOOc27RYK5fTihKuJp7PycUtkfuaGs5JbsOsDeYvWl+haUsJU
rVyI52gAVSQrK4DHMk8vfxrTBT7yIIG60Pu9FlTpZlytUDLGNYxZoMapG6ovi5+L
tsZ+6moOb2v7iHj8QTGvXylZKrKis0GhkJbscopKH73IVohx7aiY0O74tX88Un0Y
a/ayoihMaCbmXqSt32zpWhE7hdU+evT+Zsg6mmVB1uwC9/I71ZfmLNeiArXNtbcJ
r7+V804otZA329ItsgS4qpKaQs/0z7WE+3Bjil8hBP3Ejw6lSEJ/cv+YUFsux+fm
brxuxBYeg+BUqjRkg2/vo9OtFWdAs11dMgAcwta++27Gx8Hoz06hoPQMeLLlvhNc
YWxMxqT1kV0RRgosla1wVI1HoIqNMatDERqJoDmewhad2tOKPiRkY5u9E5Si3b20
pF4HsPAfy9r6apVsAQ93jH0QbtdFyj0JUnJszG2t+2lRjVoN4FR4RsTkeA19F8yM
Ai0aiXSJlk3RPm0ZaqpHXR1VIkE83MQOlxVPWCfWI5M20ViKET/SI7N8XDE8B6wI
PZtX6abR/vNjrlzVBxARdDrLeG4LbLVjUm9ILTP5pmF92Ktefhgb+5UaQgyaBQSs
pC1fsLEIAGKZIf+6K/Ass7IVN0uiB3QGHk2U0r8zUchXMCXL0v4vUVblZRHqq4Ye
N/qsIbIiLVeiE5gLfsy/0iPfpFv5OkjhFK5YTd3Vg5sWAnbJlAS6CeK6hbOUvCGl
vMVjD1iFoLFCFXzyNhqBf0kwA5qmQGmMnqR/yuzZe/A2Ys5RLVrOXldJ78W/g1FM
MOd8qQgawcjpR+koIkEq6Pu9oFB3aTPw851gGkXI+hceogmnkPOAwldCZS18qG2a
WWpA9VEdSxXfiv+ltwSrcebqlVDNKFdZiKOxmUNJjPe7kKDxfLiormQigt5MNSxo
3UgwYq8k1JMpy03QW57A9Gp/sAvMvk0WW3Gtbuo9opOj+gVQXXwc1haX8URY1wEP
khVYvePcf+J/tpMXOcsVCdyQpHjtAW3m8kHL649WJXtSJKme3YYvKLe9BPEmBNi1
JvoAw09mhksgJnhnusrc2nRd6HQ2/jjJM4P6s9oLhVoRYt6hD7tezRnSUnMOIBKN
d+YsifpFzY7WHTff7Rd8C0ddONSCImTlmsE+ieqqWIQAcrRr8rU57wB1qO0ZST8l
nDzuL5rO88P0To8ZmdqhDOo7As/0ItdS0eFkAalXOX9BGDHebA5fi8IqqdjwT0HR
EdH0LlkhXZT8Dq8xsX/OTWBEzbxJ+8IiflDtzjV5Y2SatwoYsFw9p+jStT5J5lku
fUbP5RNci/mDdXNQ8OJwVAZ9ASTPsM1JNQKHnuaTXM90XNBUo8PZNUx37jGb975v
TiKLIdgsjFiqFEYQacZHv8fcXpscYT3egLma6UIU5maQ2+nL+zVtXrPVNP9zc9CY
wn5lOtG2RIWBfjE4cnbKT41hiwfSOuYGS8gX7yPqdvZTQPHv4MI2JB8zPcR/YLkn
IKkMYkNdlc/IbBX2SF1aOAUQcVPRXh7qObexkP+zNc1KROSRoR6345hE+kNvfCxx
nm2jWZAO+pxphuUHLMEsCHOn0PY50Hr8eKmKWQaJsVCwJEdmt0Y85qJgaUgBbLI/
vGmk7bQuVxVbEzFMePUgNJHTzZwIgp9NsoAiKEDYy68NYYZgP7X8ycwb9EDiAlqn
L6c2Z0ngSb5W++uYEyzeLF8JIQkFcGyLEKB/94YW+JKs1ORlqpmAqwa4zVYkvKtq
X4D46F5/w+SqhhRlhQtLKVUj2QCss+1dhOet0Ixg934Hh06WDvADeANK8qnG1P/2
TJwGI2Y3S+2XSN2qHAh1VPpPsIFMJem3z1mrMoY9prDG40NDvbKQny+HbZv6KSer
8N2TB5yiETsHOb1I6xInrneWuu8zr1uqZ4OkdWTciQSaNCzV0JIrdweNFPApA9+b
eKgGRZK9EPSB7uvmB3sqKCqAXBgcb6cmDRItGEa696bOwDQdu3/Ox39FO0QGjhQf
7q2GatN9P9weSoFIOWFnM5HMqHIcWx0ygZyH7cwlQScVD+2pvj7PmC2pKVqPinJc
gn5Oo9bYN4BKtSp/RE8eDb0e+ihEBpXZpe5VD/HNzuf6GPDLK8KYmelXUSvvfM/3
25jkYLgvVg35nVy9GFtU3FZb6YcHbCcBsV4ATMjkD2AhDdbYO1lkhhE7tGPYpZS5
xHCwhtFynmt7/ANH1bpx+Te6JwZnwQLrXtLDnmY3PAz3C3b0K6uXBmJCvpc4waHN
TciAglFjFegfZWTnVyikVN9SrBr/2ceS5X0Mpn9TOr5CcaPombTmWKsZ90qvIYGo
z2lMib6isgOM2G/VzJlOEbPLsWgA0OLunUY2x1iUsjbC0Qlro1ZbqMPRBEX02o+q
Kozo/IX+INy0YyzpWOyhns6K68SsX6J6smGaeJVnOV0jndoRtTz8JD+3pZrMMOM/
sEpTAOwHmcjlTv2x73F2N+KCWXyyTyi49Bt+im2ewTPIAL+IwavuD5NRTDLCjqWb
/1dxfwoqxtJSDej115ODkD7wurhhwhWKXyFiL9Gg6+OpIXBgMURkhL6XoD5GOlz1
LCmSP4UBjvYROvH/yUye0jABNPWmhs+TK3f28JnS7sH5f4Z/6Q0umEHWX4yoeSFR
hPTukyFs7R2zTI2VfFyqYTmu1otKu1wBuphVfb1INPY+kPoctC4QOqKo3RhGZjHd
KVeQcpxhb4unn4p0s6eFi44ibPGzaMhagFT1q5cDEURR5+RdmoUHZ/4FLfNFdiZ4
BBeDH7qugViv9uNt9zyWUShpP2JMS/11enKgHvT/3j6biofw/bRxWr6WG0SRzWtY
GsBrzXADgxFzLKzmFHUy1JoHMlKq39k7avvzTxElGvX8t3aZmMGPemHCbTsPVIuD
ghLcN7qPzFQRD3FvfgMOnUn4rn/FIawjAJjfFAL13wAnqM1c3m3ELGC64PU21TCm
FhUCWMXAIXlGRFtSYMCQHf+7vLrnlEhPxwTb/R/m7vgSmz4FnbaLEAUCQWHqXMbu
YSErP/UqTC0zGbEiB646TOkCrZHyLK2yKuS/s+rR9+BBKKkWsas7x8AbLVCue2i0
YrUPyzSvOuFyrRjWMNZBl3R76PGC++WmbTTZ1XJdE/Pgvm40zjZl3UulEx6mUSQf
91kDmfmsvLnfmk0BcrhHZ5XgJMr1CgJMIDnM6hvJiT7YNyGGNvlXbhZM5RiCgYe6
+4rrSu4TxXBu/U95qTVyimlqN+3h5/5jTpWP2NHxHDY+kl0f9DEW60S7N93zJ89M
qWZ7ijK0Hp8B6GexIOxSGLWxmfgGGcxRTFs2/pkxkdpIL6jWavyq9HNby24G7sG1
kyrkr7ROqLKTIVgxIrY7u0KiddrY2wIbi4RZ8l8fVskniSXvf3dkg6MdH+OgA/eF
jNJeFrg0djV9mvOc1Eiyu2KgJL9UgLUUbBdq8i+GOL2XP+P5oz1vTFSPp0PGGayc
k0fVHWf6Sf5AAG9xw4srXzLd/wYyyJnhiuE6NdFrpPMmLcoLwIBf7U1n3aLkP2Au
rSGcOHWLT/HHTexdFiomENcMsvECoq2GH2svE9x/IotZVngJ5cGhXEadiHv9WnBV
buRctCPygwUqAL2X8XdTBnRgRXp6MbEiLZRbNEG63/8WfR6GCA7qpcG996zS/auY
WeKMPlrghgNPgE7sVUChEb5mPEY5/TgTBJEfa+dT/DrTD4XA466/dWSHIZ2jUj1V
OiNSFd5LTHli2G/Db1dXVk6YHx06SI9wg3FYGIO91AdsH05I6p9jY1wUg0NrK1Cv
vZwsOXxl7vrpoELCR0/zneXF1PuhXMoU9z2VXyvJEPm0w9E1n3OHuUGaGy4gaFmT
v+/8GbEsesIG+4/ex6WaUdpLH6qQVhiOlE1WzaGTcFaUcNJnaiuOGVr0JYb7ApOj
N1fTqYzTNxyWjXCPktctQ4fuBeF62xL1Ep9Eck7hEvRpuYI9tXTTcGBykb78pov7
qzVVbrMm7tv6uewYjngqL13zZx0S0ABcDnZZE1m4k4rTGXl7p9dixLysYO918OC/
1H38+6eqmjLZF09gtdCdTb9cXX6PnJ/a11yzFYcgrIK8fM00SkNVcTht4lCy1mAO
8sj7i3ixC+wKUplsZeIMx/T5EilPld+UEVPJ+sqziH9R5Fk/xneHune8WPldl3bX
uGDk0fuWU/mWuhH03/yTeMK+EMUEF5gLNmGLe8OZhSVCR/KVZTYSLG5Kr3sPFEsm
UrgqpS7rd7kwgTJ1xKO1JrHyzzzcZ3VYch/gvb7Rm6kGE4NMwZqqjcp1U3CL0dmS
p00WWPKXThSRwGE+9iVFE0efZ3wyGpTxnd+VQiYNykzYYNYoDcvVeWEQSSKSYTX0
RdauX+K8pT1FpKEHcAUjyyuqv38Si18fJTOR+qMrjxNGM9DnScl8roZ6S4DqXQ2x
5oR/l02dpKym0DSk4Ci4QrCoHebwk29M3+4oUSmder7zz1o9Duwg+yTgDHB4hoBs
Amn+Bz6Xfa5qspWQy0/vIv10x+BjCz6HKYjTLXqIQxUeF6Y5tPIUElSuOmUFv1SN
aA9QCyFkUCTLNvXqzPOEP4kIWw3Rxi59FGBA+xBqfIUIMmrT/Pk4cAW+R0LTo9YX
tt5Yr20LBOR1DhZoDzn1q18c2T4Qv6C3y5dzdy1LcHXpEdrwkIZZHAhYw0H5JkUo
v+a1M9FiwEb6lLR+map6ir8cW0Vl+ayGpaMfRMTlPpD1h4g6CI9dSq+8/ZgFPKhS
0IbfPi2jnWnqzMxJHTtQS92c27JoXtUrybElgS9wwwJzu6RR3s58DsxmB59ID5jv
ssGoOlmE7GaoThzKAezmWCkYEaC/wnCQKl1AR64eVEXf9SD/YuF4r7ZczbuwAX9M
KqX4nI5OH9pPETsZuMBkLXesZgjqyx1u247V0BTW5nSXfDYuKfcqXYDIpV/474Ob
QDaJcmI0eYZ1NcHeBJ8fCa43pMYz2WDNv3i9/1TS1oHNi9gbQnx/B/sJ6uCZCrxo
GD9NnpA3qQLqsNjjLzsayDD/XeFW6Xa5qvJnF0KRkjHrittQMzTX51Z1Ob/oZPfk
6l6iYyBSjz25A+08p96HKI1BWqJnzdWyCNGUYjGCyzIK/iP3wuIMXrGbdhUe3V+c
jvvu6I0hCGBxX83rzay007bnyXL1bXiyBIw0b4WNfORpofxh1eSPoLdTcTc/QLiC
gpPDKy+jsbPfQdFaaV5ov2CHZuZYrqI0vfxo6lv0ixKCktOfZbXpne6gwmSSQ/az
wHGWRSujKj9KnMylmCV4cIm8gDEmdMWsJr5CI9yvRyu/AvE579S7knHDvlXkGG8T
MAAj8o+TVFVdc0jMxv6gtTNKJl1EYUeG8yBe1UDO4naVx7/vY9YxJZ1z54RpMWdS
ctSyWhs3BVCXUKLcmOonuggaHOy3gjdCLWDUtfAwyw3PBhYJrji5pi5UYGiOquVy
m0HDZwFj0t5f9ngHw9R91N8rVJ4/7ufObEOKjTfmc6uRsiiRwS+N8f8JN1BrHkgn
jUQLMCPAzWJFoVHZYGhXQUF/yRy23zd6YFIZLio68PqX/bD7NdzpBTmPZKiobnhR
LAP2UpZ1JV2rhIr7FXG+8amPKCbk97Hhrie6FdtbKbhoCR7/VVvkT314XxS0OIiv
WAzeGr0VUwbAlG2RXqBM1v5g6t23Rm+c7EihZDzGvDhB4Hk8hbmXLxp9SvIX+Gk2
ZJGz+0v9O4lIWknyrYwVmu3hqXI+lIRTN9LEXQJ3jgKkqsKpRoPtxpnvKaGUjTW2
xtp+QDB2sEL/7UKmF8POkDOqGAYFpYOU74ZUfr7Ba5vKyK0wn16RmCSNLKYWBsn2
eghTZeXSP//u4WRQHKGTHwoY+N+Rr98CLPDAFvQOfooXIuSo/stQ6PlxEEbFeOws
TrCytNg6TXiukgl3vx9qR3ogVNsUkp1yWAEb60CSMZ7n7tU0lm0oX2sFv2ddDadv
JMav9rp1o18jU6faVwSAUovIhXF9wlK1mQiIQElgLfM/DwYvSkIErYdxdDtsVhVr
86/TeFiMQj+wD6RieF6RTRHJ5Pwt/gCV8j5vtdtClWM6v3+Cq5irpYuOwkYg/nD6
XpXaDYGpq/HnmTE5KQq+RMOdVo8ziSdHRf8NcB3eALYHmPdAzUZo0DcZW9YfGVbx
V2yB803wHgBrBmZ/cKR0i3eC/EZTeWE6ad0C5u8JLjKywglu06NIwnZjNb0RXtSt
K5Pxa9nAl46DUI4u+fEGV8PgxOAMIxD6+Ml1djtgynAK4FBonBrjacRyIbz3PMPE
ku5WoLvqfHv+SF5qOcwuk6LFuhBMollw8sZ+habcuaFSETZGg/Nad0TLnP3wT04Y
F0ylVTo/NiocbsI87tvGG9FlCUawRENj44CJyWrDXzF50B4RFhXUnvoQ80UA8ru3
6E6rQk6TOdse2Ut9g6itaxrAHw4cTXgfqiCjOWCW+1MvQbsQYm2r/C366G9/nQBr
JUCdPP3JMu8O4cHWDXN734f7bxnZVbGDklSlwuwSFV/z1Julu6XYSMcPMzVjt1wq
I2xkBeT6uSfZlX/8iYR1BVfIGUlGNvxADxoW1oGZ4c8mOr1cIIGILCQsTk6fqhT8
bX3Hf0erAohG2Iq4Kuyc1mlG7bVlowOAwitQffqYhqo6ITjx5Kp89ysFaoxabA36
uyf/mO/l2RZFJUcNMNHekWcmpTU+216o3PBJVQJsIX8quTAuuBoUBkEMJpM4xPpU
ajEXvMpXaej0aj/JNVC+81qj4o2wzw2vVM67uvuG0x1ljJD3yk3f8cd0IAzds+lX
j/VEhfuy8CoVRbIw1DISOAn90jK7Quafv1eVMLyS948JnzkNufuVW6px0kviIotZ
+Evo0+KSC+E0ousizwC3zJ55l7O7CNx0URCqCKKXDlyoyM67MDmZVq7Wravl2e5G
Tu0qYqWCM4/fGbw0eOL35X+dG3KuDgvQM7YxGdjBNiDBQYEoNDesMrDSKt/2pi2/
ldh3OhUrDb7556EixBuUNB8RJeG5G0NqyDKGtL46z0UciAWsrxZd8KCS+xFhiL3Z
QxepfET9uRzx3MzIZq/Y2Lwcu/ca8Ns7f3Is7UDfL9Gxy4gbPIg4w21Hz+yHa0DX
asBEqvhhwe6YLx+CI2mnFY/aJ2WjgTNfvb3VU9rtCN9oqK+tIlkJiO7gNqGDslrJ
Tg5doKjTdsi3GxLZ/cdh9vt3tNyTHwsHcEK4wqmR+aqCgRd2/WiIk3xrc4j1bLa/
EqDVIonCAzl0egU1i9B7er6X8SSkFoyfUi6VKVN0AcfKJHw/0plkeOhEEWUFO6kD
O5sBQ+mqNxdySDGtrGMxI2XIHm5ANI7qQTA9YRpiWk14vk093HPQ7QmkZynst7aJ
OAAZk9G67KHHXcbRcvXG5zVTk+KRMbnVtWgZrbQJPAIqTqrgwn9k94PvpF4iZdwu
0Gk9rt4jc5VNg2e4tbqhp3FeNW6AOUdg1lenTu9xusFtQ5TveWanLwylY7+ApXLD
U60nOHvcTl/v8z6jFAvQuA1R0iEtBBFhJrKGiAva0m2K4frE+PZTgOfUTSseCcYV
rAMIyt/g8NnaqalT2YO+sBg8cs6CxdMphzPQgQhpwYNdn3SbXeh5WkGJoMN0VGQ4
7HSDfS0ib1BVzcwDWH1aokiAuFeIAyOCkg1UVBnrS5XjdnA87x2TyDG1fP5NYfpM
GxJ+crugddQAjS50Z9fA8jZOg9qmM5NqJf8t+GVCDs8qW7AQEsJ3vtf59u8WuyzK
QadjL2snFQ6ltG5bwvDrH4wD6AcXp9MxxdeYaSP/UrXaZiSWdYig2qM4mYsf2nQL
NyKH7u/tpKBmRS3HOKIa5NWvhGvh7sOr9QZiYVMxhyPO3KfhKgSj8TP027lHcNi2
tmhCtC+XBuwYrituqYX2SMwNgCGG1G02Swnf4JYse0JirW8zv1COV9MqvGoIc45o
kQVQfBGnm10jum9YHsdVb8fFhiHXP30ZmFai3YeAT56SXUESXiSgtqbMvJ7oEoJY
FabV7860IlRaqSbMmp2cDYCmD+99Lm3IkWJA5dw+9l5FEhuifTIoPyc/ofUrOXVt
4T1P9pbNAFAe29cqSKwCBm3rYdxz1A7sp3IMSyVSZKAsK7X9lUrdN6W3U7+W86cw
1/T5ASdvQaZ1Tk+8VPt2ZJa0Y9UFmxoIdonfw6QsdUgbHO4qn6+bs4OQgyKDmISd
P6PNd1s08Z2sf5mzgRqZBaS8fYJZxR8WmVH/nUOh/H+O+RpuCET3HjPv8iV7ajBP
OWRLXt7YvklU9czyun1mA8SdPiiSuP4M6vj2FxneL07BKa7tzCjFAnEvKHsKUXXo
eGhd2ROZzLFTgm9LSWbD0q4VylV5rnuPw72ZntyvFurPpkv33QSvLgFN3ZH8cuRD
BJ5XH3Z2S/dI6WDDolRUPyY04lc/xaEHVWdE4xiNfbtRqrxoT9VcVigfOKpYdROi
jemViWjgpTJ8r6leu2uQW86ILGy/gD4T2MksQtQQCsWOhzR8XDAjL7BLgw+Rb/dy
mqxLgJLprVHWfxzjnzfNPw6or0AFyd/3bB0z6IvlngAlCX/JvE2UXiVx8hAELnqM
wfQ6f+xeOo0jC9ySjdsuGwSJJVllfOUjaxIxaHIkLj/+J7nDWwUZY7xbSFI0wlCK
BBABHYj9Ujg1yEM2H93PCrNrwPhVqT2INHilrFM3HqVq74eOQmPSMikW/+Ow3TY6
sHutes7msZfXl2Hqda2TOkOdkshjV60TNk1TdVn2ZQEetn5g07xA7IKdFMu0iXfg
pIpFGjoDaRF6zE88vmVbkg0+KeCRRkO9I7A5g07JDpZGBBxwvcToBt8FPzCYQj1U
qq/HcyP8uwIsGD7pITvNfymA+gzq1U326sttcVayrRzuNCVXr5qK2iru5ff+OsMM
Sh+tuGRbgeCHgON+VwZ+ZvkLg+sdW24U8yw2ReLEv0K9R77+0CnkynOZ2B1C/qRK
jQCIVSeH/nRvz+p/SqCSfaIzixe+PJ6+UY5dav99el09LuVgy7u5/kj+19no8WQX
SpGUU6kterJgXHx9nt+/7u0V6ZoV2zS2Zy0tDbwbaOWDmFBPLlYFC6PjE561EwkQ
2zlfAhs9KkNGUIaSZQ2TncPhGovfb0t2qslXXt7uyrLLYncba3DJ3t47H1YbqMx4
tJ0EoK6d4ZzZyd+uXaXdjxK6/Cd6Ym59t4qyDu/EkQofqxxk+0Y+Hl5fdR/8V84l
bS8jp2Bxf4AxkwfI3RpcNoonejkl3voT7d7OmWAgDFc1A/N48L3WDTsE20JkW1HL
ZxfXefI8d6SCcAMAYa84sAz4nxIx+iDiqwQEUgbaE/j72ByIS+KHMDdkl2wyII7d
PDsKPXRWYaKnMiJ4+gMTgelE7LE8l2zJUfcZLy1fntaqW5S6dVl567LKdH7Vq1NO
o2KChy4WfzeX+UpwFU754Y3474S1NNakTRLXZUbMOMtVbogJMYe61vEa74Yoanvr
moJVSe1ctbESqUgZMBCtAkTrnf6nvJuO6a70PsWN5sup0DivyMfrDCLFYwKPQ34G
E0SIoymz9potVofO0YxPv/5o2RUwcfZZQcf1/riH2UHK2HAN7zbOddRR+8RdSKbq
0rGl97v+oUPg1jBjIvv4yPGyv0n+gRuiRqPftpNJN0Yh2g3j9EOItZ+3iHEYLtqg
Kyikl/tAlo0i4t4dHW46MyMRHrcQ4iJr6iA+qTQpXv8iYJqR4H3GUYguLozGn3oE
1EcpbgG7lUNDJol6+0FVggsqgxk2cHCOdL4lCvXWyjo48UsvqApYZO0pXWIOfoA+
G857cSQn1j7vOk+Fwj7d183UNWX6tw841EwiEkvhQhNsuObv+CAKDiBwf2Mgoti0
cwdrtHLWAP5Q6EK64RtqXJ/vdg4Is1s5YUU96rbfzMUiwnC9dfSwhdccSopFKfpN
7+Uz0N4KtrYelDdrtkRLbilaIifIxLQEn6MpCh2WhgTYPYa6nH1tFW3Dq4T9jQKc
n5A3qLfHc398oIGy9TqN/zdEENaKh5+aGGRjSlBonpFpucYFit/PubiGoDqDcgmk
+0396BjqjiyG5eagYzEyrtDP7c/JNej7kY855llzRiuzbap2+Z47aGJIq5mricil
5jY0MZtWSmK2hA5cH4DZ/8QyOTxThtYWm+nLf45aL5Y4EmcaVYotgOSDtkVatsOv
oqSHPJIiw7un7CFSozw0VE7xVN1A3cfmdOKkDftFwBpa6SWfBBxsfyVz+8FoNPWr
IvxJI1ylA8OlOV5UqTQXLSpFmNQ5W++oIw1CyrRjR7DMxvIKMok/KlQ60TvtO1NN
PaNQjvg1XhIleKuN9mwKP60lUmXYFbjlPc6jZvX0u5ABFlU2uNl++3jQNaOsnKvO
nzGvsvPnHgNdOS/L25K1efrAkxYTPz2ZUgL25KLVY8Yjc1WSjIejKFvl/7T+tso4
aFsrlUBd1qioG/B+4llWt6z4rxhuJHaqYvgON3lWAItTF6g+VL1mFw597rKuA/PR
NdG8S5Tg/J3fSRTppJ7yr58qYx1yTmsm0+jXnCREA9g82F5itzfU1ttJ0ZTi7DYk
oNUmlBjtqFZW+OIckCbnrZGSHa7+wv/FyrLoUXBy9raqD9yYDiTAnCFvN6JXGZp0
K24S3vfCVphxVm632HRRxsk09rqNzrpYIV4SSG1Eahl62C1jw24q/5A1iYdLetI9
Kg2Gcx1/8kRIJVrl6kaGhK7FAIl5juZu99cGOb3fLvCTiC4tD0a1HdA+3nKyBCPh
n4KwAHW8qEq4L6stQ2alcjhOpoAWhywNQhsl/blTR2rfy+FtumXvj2bzPm1gUuke
HXmHEyvj93vNpLiP7Yv7d3PziAv00x1yWJLeD9uAIskh/UPE1yUSTM9JpkJ1DihS
Zf6XHiKXtoKyvdc4ZeUBZz3sWifC7hRPAooUsNTCtYo5O+aGPRsfmHwrOlQDCXir
3b//aIk5QDNCXAu7nkVTEZpB0ePaAW8WCZPtrXb63K3dBcxMUsZk4JTVa4Xxfmq0
XAfLL5f9tOZxa1bkwhtH60shfs97biMY6YC+0X1FMZmGaPaNlWT8f7PnUEJiD2g9
wDQIRfTFO1/0ApDGLStNiRyyV5WRQE2e8AaleDQsit1Ao62RRcscTotvnsUSbluG
w1PhV4BgUp49BSxiNxZfQTuFI6tPrlTyKJCYSLv8+7roC6ZWjBcth1D0nGgo5lBc
4TJs6w096V6kRs+If5HD3G+z71dwwD2JnGPpt84JB4g/06D5HBO1ZG0Jpb5hKDh2
NmiQLiWA0DszDrnJuDcoCMYBDXMpBZIVopQtz8WymUu6hNdeaY4xxIxGMQbwowYl
/BmQ1Ovy8uon7yDyP9F2XZD/T7ocYzpybIZxZahSC22YBzRc4/EZgCkYXg+ZR4De
D7sXo8tt8XWYn4x5A440LtJfbFluYFqsgxFyuZJdjfvwRh+ktcbnWt+fOHEwdH0d
irFU83nXxB9Ab6bPYI3QeKqX529Otcd+/di8ScFcvcCrXTvWeYGszF/LGXx7r9Qu
S2WoC7WuKG74LNcKYY4p14pA41mqO+7LF8KuEBqDPDsfqlaTIaOdnnEKKf8OdjRz
GCYRPUYE0oTHBhQEaMTa0yMDQIZ5Y3dzSNG0eJVH9crXV1o/1mOZ6LpG5YsyEI5s
go74swfnRzIGWO9gd3Xe7ryIHp5Qs/WkkZQ0Xpwhmc3j9yDKKAE9BsGT6uZut6C+
oYs4BXCNrAFamYhcrC9mnXbpmsroK4McO3BTJaQqN6SXjaGGWZdr44PNnISK6T8p
6rXYsLLaoU9t2CzZDm6ECqN0MnckRW2NiG+V/E3SBjrDyuUzDHhgjeubyCSyz+6O
CXweaFTALVhoy08OWKF0T/vuQpvIXPGcFYasFT5udbngL/m7Q1go1AO298SsK8Vm
Bf6nq3+osPD62Edrn2oyzzS/joMUPYQYtJhU1BMhWuCt3zhXunmCoUYfxFXruThT
vW65ZUCtwRW8xnAO/L1kV/P6lgfCBusWyjRj6SoMi//GMUWstb3EI9hetQVgwlkW
bJ49paZs5nmE2Jg61cdz91WKX8H64hXtrkX13z3Qx2zBLNYKptUnIJu7/BTXiouR
7tW4Yw2zOrGvzR4vl061Xp9LI5JssTtUUTJFdaXkPttqVhWFg3Mb/PpkvYwgTwR6
SjXo6NNNjbvHUXKH3mBg5neuVLgI+52LysUxlXor+RRMLuNiidKQVIH8MAnQSU/k
s/1nU/5QNY7eSS2su6XuEFHIxiEbk2rI5dOj2SJ7epVKc+KoWl/Xch6BWiiQ7jDc
GFKsi2hJLs9Gv+9Vo3AukV+sggyN3cD9sUNlL52xVOtSd+TLBoe1k+FlK7PZDOkP
ST4Tch6hmnVtiGWMP0yMz1oXkElmBzw6AV4SuDHLr8vIFaIYBUsFcWjh1RMS3Hom
/aPNKgev6aFHvC+rYk3FiSATz1bJ/+7xxXVv6C38zv4vocgiOi50ghiMvmqh2zy1
pu11RiNFrw5Z//iUFnK1889nxcnFqts3A5y85kSGnrtK41fe/viSxY7jV3pt11S3
y/bVX6Bt1eaV8uyZ7nSZU2BUaYOa49TLWffyg2E4eIuhiS+P1uQVIDIv5+GIR0ep
+zVx3SdqJZgrV96RTVqD/xRAvrOKthUhL+GuhY46FIgu3vYybFHDxQZDiyHXR/x3
XuvtXmET/VzQhXSHRshCzQ3t/Rx20mzC/B1Lg3TIr1yH1U0y7DUOA13Q48NCUoWS
e6HHz/gw80WGIN98seV5E3AHkBJ7j9AtgGRQyArLhBmmE4slZYEiLufg2zmzJ1Fb
8RmYmB8/a6TFX/p9VUenXRPDdJo6Q64T/VCMPlxwnafpSxigPug6dYlUOf7MF+ay
hzNukt5B+3ilLFYYcFiDULy7QrGmBz1phLNXcpPy4z/DPnw0+jRob2kgTlYBT9Cp
9caBMran24sU6Eia1ymwrvAjpN7YRxvsosgmf5g6SKZBj6U4EeA68d3RKSkMEc6U
AFBzR5/PgaYqNzuGXX/DEuGe/qhP/nh/0lK35rt6YB9bdFscjFwN/qyIh0i2JTqQ
8A9p2Y8zvhpsowPSGJu9eGlDzBbd3ybH+iocma1xYKIUlQkWUUUk1vF1Qcw1Dj5U
1+2Xa0qRlgijWaseFOXkipbhWNAMyAFuulB55BhxjSHvvTviY1lPIiUQZIpqpOL9
h61NKDuKMiU4194nCRsqDU0xxYUGUlWo3tbYo7X3jZGkS2KsNdTWU1g55R9F99N7
s8IJLCInM/crI0hinUXpFZeyARBnY+0R1ayBgsIyOX4U8hcXCO433QYvXiUmK4OW
z9IkGDQhzwf5Uq2RwQDxZi0RVWA971NExZ+f4rQAhltA0Wubx8Y3V8Kyut2/CiEL
zLLOzOai7ohpBhXkRRq0gITm0Al604mDoIMCfkQt7Jgn0ak/SnftiguNzhivd+Af
NsoQQgtz1FtviorTC5GSxvjjVI4jZLv++aACjN2Rw4J/ehASfaL2UZQ3yGzBdgPt
a9TqBsUY7wSts/cfFgs54Y8nqEgxX4O7bdhLIIC8r4ELx9ROupw5oHYup036dFb9
3qfbg2y9xEGil18qKjMJGWTkJSbJE19H13bU0ZUMrTVoz/BHH6KCCCVJzk1Zniq6
tOJq5jcy1ldG92dV6AgR6Wb2byDgd6OGhetUgY4LBi+8oRdCWE7NoBaQ0npwP3ZT
IzfiwtZSQyT+KwJrxxPIoiFRUIsYxUG6L++6NHiW47klGiuZf49016vHaaQgQeYW
hUbi93cnmWg23iqqVtWc4YWnNzvfgOsgWIp9MTpk8274whFlosqUR+W9/5eJ6+UU
0aNe/19W6RLKLdC0nMOTJwUeMnM/p+q4faWoxsFMQEZHL5BrXQBZBUmv9+jTmBjV
6BjnREBGM8GxyehcXMFanlW6AffsYECwXdb5K8oXmDePvMggHNAJwOs61qheREfT
GVJJWwRlScUHWDATemEEefVTNL2g3klFWjDki6XP0Z3PoUe5TNy/Qya9VByy9Lc6
xjGiD/yTpcB2Adz+0j86hLy/k0sX1HoiTCIxloaz0uzusCWyvixmbOMtJwpMprJT
BM/GPzj8NCS2sdFOZntmL+oduROXyIlGjvToEa6y2Hd9siSlav+XPbut9At9vUUO
2/JROlQz137ldt+kynzNSPPhnGu5dqNUFt74ThCzMXpD4D255FrjTMDaFq1AmGin
xma2phn7/rUeP304eX1QW3UBl9btKB62NywfQRHCVYiCyYxkby6uP+FHtb4goR31
EBDQUuXqtG7/wPMb0XWluXekDkKh+9TroKlljMdjJxiP1Hhq2XR/+OjBNTqfI2rd
ATWiyj3gl5tp+QWz2qMd2+kfstXDPgelWbIhARTFI9ZryD7fdO0D1IMgG2iav7Uf
UTyRBjIlq/PouIGauWJyHqIsADaSPTHmR8CHdEPvZmropn9qKmV8wmwxr2zYR5TS
Cotgp7PZ64arOIwHp8o/La1pFJHrfnKK1AzPwAbm5rfjZoscZ1QRDmYAl8nKeHJf
GfMaIzezU+3UsprhCZqI0B7Si+JVq3T0lJdso/7SSQVAzfji8E7bj6iBFZZLcdQu
DfLuXHF9EmvPYxaMQpWjvfOzPL6FnBgM+QujMEFrPDY+KrtLKrQ++1+zOBnrxX4A
n7SFJe3xoqNH4fSvo0ufLLpIrcqHjuONlWFaEjyyaEh4UBOvRqJ2mp+mpZnaM3g8
Q+ayggo2qrlHQ6RZV14jExZD/uacH6nph3LUvD/IOII7841l6TnuVUZMQDB2bBRW
LPWLdL1mldHw26AblmqQ1vipJ3LYAUiwradxeRNVaNeWT7Src7MP2RCf1QCZ56It
4Cq11hIGIipPrWuWgkSmRxazsRCDKK0UD8I7AaxXpV4+Q105mJgQQNGJry8Ccf1l
9Bqo1WPK9dxQPYj04zTtFCChtsrFrCtaOAIC3SsMNUgD98J0/Msl19Fpybl2Ec62
SOedqoezHSrWxQNNnjWAFmQxBNnFsQ2+GJa+9KjYxxAeMqyORw+rDYpj7VAmLjH+
YP7q+pN21FXOcz1K+qDdyTWTBiPPUM3TUITzvUy//QhGPKygviKRfEwjs4sTjRlU
xHxhrZ3BbpElveYQG6AHcEeyy6Is37jOjm2+fVUMtsAD/AbbXnPwXvHpNnL/GcWG
QKPzz5NcbzO1R+Q0JOWFektRv5dWV7SeoDfGcbKrJMN0KKWjPl10rMdBb8R64dvw
78GKWVvUXzARIF9o1JT8BaL44meF50cXqkvhq6LvKwZZgLxdwnJmDzNjuBRVr2gQ
kjGHHQ0Ln3D5r/bBL8MzVGT3aTc5RCnvRvRj5A7zvSSVD+zlq5jtF7sLgc1N7dYl
7ZHqvYnsQu+q7P7WvXvxEKiwKIMunmR5HtKaZqcNL4lxPLOQlLc1x48rXBt3xT68
Sxl4D7JVYd93h2xhBJo8id0DpFMrByFoSBhpxoBbn9kxhliWjqqEkhTI+8pGlnQR
x1+NFsnN9KilMYPkMzRus+vZM8WykGD7V1kmpf+Z46SRLuRBdWi6yM1jOmxQjLrk
mb0pb2+rXPV7zHtZXxyEoigP8ftq/FdyrJdRLyWr6nK7l2ktqtgpJMskYLsdTL1h
WSMU58+rUFFgjRt92yulh2dLAMU4ERI3o68ZXaLru5OMaogzBXwmBOkUiY8zkaVX
jKU24XD+czqzH8YjyQ+BxZffUUyiLgivBOgJ8tT6EpxxRXe/WVW2t6Hn5cq8npJz
0WPGHt3MLi8Hs6J9iPUKQXuZqh1IZKGFb6PG/nQeWS3vN6wSJ6/tWTCGajiFCdww
eKfTD1lnWSPc7QVKb0iQD/cUbrPud1i3fNsSz62XL4q0O04BAyPgTIXWrmXIWAzf
wcxzFHPMkITD+J0Jx/ACbAsZOJWlLilTum9CHO9jSuD8K7XIa4xP7cAV83xSULq+
ytHajFGGLAeFNZ7RovWCYB7xAn6NNtobC56UDHrbQnvaHulJymCa22SJJukEdqb/
5U3qmhDpcPz94+GFg05OL6KNw7ZuuHbeSJ+IwRJFNn5WhDnsD2QF+lM5Hq87uOcp
qIYTMA01mVOYJDpUw0fMNv/sKyCoydAPqOeiht7GSSxF/N8EPe0HN00Osg1tHz03
xIaruT/ynB9ukr3S+jKhTd4wNSkPfTYAGVTFPa6kVU7JxSWZDw/mnRSDQUFlZsVA
BEk9zTjnL6fma5nXWe1dYkUPmoXao2z1KOITgsxUGDYFHdss5K9Fukl/oW+He4A0
hDxwLmgqs6h49AZnLo7sE7hL3+LErb/yrytz+GWZ6pC+miNOrzfn1B8E1FuYr8kM
JalxTtEiS7DKpjks+H2sjb10hKIeg4rFDz5grDG/16UBfaesaM1UfS18EluATYXr
pYkr90NZiKTA24ZLebvi/2HRkPCdt2+uIQ3jyBzJZ+4W0iPorelGsxC7r78ZKTyR
DVmb4/RMjNEVgF69Ji1/Zo9cazH6nz4uWa8qb4aZTA22Gw2mPMBuex3AQfuBQtZg
8aPiaaj866f6t+2HFfXaPLwHZuFop2kSAdD/QdAnE8lBN2P6Uf7gNNCJBaG7pSEg
obpbnYFb/N/Jff8vshSJUQvRVdsjXLWj8IbOaqmxZwEiA9U3EEI200P1XmXzTBCs
CEdENYtS+1Ux9jSGbyxz9PDf+fhH5pCAJ31gvsaftJSJaOkir12kyIQUDkSssa4d
9IWOA/SSYtXWq8Etj2MJxPDDdOyWf9sYWal1RgP42e1VPv5kBoNQGVPzmrXDbfxD
XWJSIQzPdd+3aG1JIF0/ceY21jUzrC7bkFQY5JRQ+4hKaalk+xLDTsNJ4anUZ3SJ
jO71i7r9NBGBBh3bQdL63oSH8TMq1gElm2o4RLsPAFQWXzM+V8ucpToFZeaAZ6TF
myizIrb2U71EyxDzEDGcIrdAiC+FAcvv5GS2wlJr2+A9ZaTMkT96h2oF9ZBycAAG
ePV20T5/UzguUYZzOtlpImTWyWQRTl0r/Ps1ogNMdpeV69oekP/ncGA0a71ji9Dr
ZwbWFOJqCs2Ite+Nx9htG0Av+CBB5zK18zuxpc+ZLa3ThYuZ6HbD6HmkgUe9IhBc
B/KJwlff4Pl/+3EE7KGpsiHUIkH+m8MVjttDtX76/+ynFQ7Hez4ENDwPieSprSV/
nI15+LmIr29NjhVM2y2xdJea6Q+uSsemL4Gas+BPv2fO0m/VkzZ+VgJ8lLCCb63n
giS7BVIhsyXO1KNiVFIcVdQt38WVBAi5YGObTBHwW5hqpye4YBrf1jqUN0ddnc04
AM/mEzj9+c9Rr+jIeGLJaIEx+hGgtRwH7Q2IBT4Z0JPDi3n+hKRBkPSwpjWBO/+L
9+7Pz+4gOJ6bnHCuTJWZLU9UB8oqnyDWc2FPJb33eMmYjj/SK2Jq1vENzhnlSDb1
yO4lAioqqdpt+7a3ky5WprDvz+DN0j8BvrFuvsGgxuQPFz8xMd1yooSTmbiQLkod
xf35q4sAvhqXMUD/odx9+4mCDvVFCe3BBxXNILtE7nq3D115FDva4HVBiBVwMZsq
hQxIMeW0/9WHpCEqYpZlfbpnldxeepSCHMBTm3yoo9a6EFKjnRmkyvFF0HA3uMOE
Ov3VsOlw/B/AJOe1+4C6QszQN874Bw591LB5XZYkoBJFm8q9wiUgKqAHOi3OjuXt
iWUjRobLp1rZk0ID+vx/pLFxq3VU/MTKPVFRhOvC9iXbG//sKTUp3fCtrxb4qaXc
TmO9CS1cy7naOUjoz9fEFjqRmdGEHZjExnYo22JZpZHC9HFLXi5Ect5OsKsqCgPw
MlDnwu/9/v+Bvv9aGohiaj9uqveLkkEAx8COg3HVIqycAPgQk14Cj84pIa7/DrDv
O0SLaFQI63/cGhhM6rVdOz7+S+EX8zO4n5aqFt2zAGHc7FWNFWQyK0N0qIaVLlMi
CQMWfuPmsAQxAO5rBnfGcHGKtWx67RdxhGrQiyJ67Ir9LnRjCI76piyPxHl+8cEv
vel/pL0xCjnqjSCOGP+yQ2vMXT3ifLJK1hlDO/dpab1hOpUvFRjOpVxtZny+N4gv
ivYX0naiqLEfGH0GZp/nt0gpHz2+Y7hWBI17k+60O/JBcWLTx+A9K1rhjvqKmd/4
MOhosF75QC4zAe3BKlquCOEDZ08XTbVoypmVdEhfdn4ykSrfOZSH7dRuOhtQH1us
7R/Sl+fQB/8ffgQvQx+X7bo+8d7pHUztgDok8CchONmGnSMp4Xg9yjliERMWpK4l
2g+Mqy6NJ3EH8B7XuJnu25TPgtkbb4D5fJx2Vu8mWklrBpsSq8DQnhBj9bc0/H2Z
TPkbxNN49/zqatyx4F03ZF7xbO9CeSkFr0uI5TLvug1bFDxRqs+QW0SmN/dKl33q
TqWRS5ZNtr9/uV3sK4c12RttKQx+QHN8ZDkAdk1mwYe4a/RYUGJZvwuSjS5a1Ypq
22B6XdkAnd5Gp8ORNatfE1+9ta4TnBxedNCd12Pr4WGaVmDtkgMR47gsATIYcOHV
hyyvpN66HaUFxhCzm6/FGq5D3OX/cSzKkxWS3H/bmCFCsU4htk1nogESslg+ZFsj
onoNSzhpIiqUCiRKB+nG2LHTx9NOIWG419rtfFKGVFCAOiWZmYhid1TmdMAD9JFB
4VSWEpgnwLUqY8UA3bE5ucNj0FoN0SzSAhRPKb3ZKo8oLjQ2Y/a5zYbQC2ZCrTZy
zAfDbIgNwgDo0K2EvuXoF9lHttwzOVbHILOlD6hDI9AREl13mdozZWS0TGvw2yar
qMDYSNgkH2zU3ujmbd/Gg1DpbuzjDhneEi+53dhMKvo+oxl5bwOYu18kZstUf9lS
KS8mzy1CPy7bBY1DA+xfdx4dM8McMezjmfH65hqnKB2QGmPPq2BUxteHdWnX250G
vp346o0P0pCqiggWBnrdh5eXoDZNE+QbyY1rCwBAT0LsnNKef7kCSMY1zfxvXNQH
+SxagLn1k3h6WJqaXwhqh+8c51wHsFvPdVuRkN+ZLrQovUzjfVAf6mNg5XXHepMY
55kjClTO64JNdlUCycGQc4gcZijHyDMHikdkaxWkmmvH3YH6CIX5JsQG90BsA/Ze
LgewePd4EjFQj0mkHlycXZZie6Fg9OxGe6GLmJlMUF1I08bNoRE8lxQp8K7Vsa9d
U/A99FaAcCYyMkqqTlvtfXrkEzbwJ+8t4eB6TxUX22hlRozDPKVVfCGKDZmu6uH5
jmRMoHjQ8gX00HCobd1thFYRChmB4e0IW7YQHjD3n/ZM7Ldmbx3e8m/2L6QeGKXl
jB3sbeEzv8lGMzDVNL7DPGcq2P0sY6SCFdoR+m6jMsi5bYGhzls+Gc0Q/AjUD05J
BUda6zOu9JrA2g9KkS748/6Gn/2B3bPXElT5AahgZOz8yPIS6c37I4Wq8sOIuww7
8QP9HYacr+PR+oMjr4ElpegmdJNi/+Mu8LYOcMo8b0AKE6EUP142Zf9tGET/0sUb
kKXKnPo+r6NLnH6VfMvqs6VLKWCMhRyoHybsK1Nhy+lZZyFosJW3OdEEnZ+VRpDX
CorX9PwswQYGoij7jeZn6Pyq/SmwehfCNl9VbWs+UVF72/Uvn1Q/vWKiK5nBF8Xc
dLJM8QSOnl7LgSGd+rLecgUFyO10igPX7Ogcq4kDh8sVgOH8d0qmuOEdu3JM+xgA
5KxnU5G3H/VkA7HXAd9yaRjb+edfzWoPUIbzt/rHtUH0mYpE/cAfgQN1XdJjCsCC
9u/cTvtTBXY+DpmdHyGSpzOQbjCmTSURgUpwKacEJfqbQPtr75+F6VchL5BbdIvG
sAIwzNsyBBXuoFJgnBoae5P7CvK+LEMheaE1aBp7qkqnWRtJYhpQSFEwzYJBiUJh
jerPjz75sPvguHq47IQC5QVn/swg2LGk0jyqFByIrsiTTXDhrJrNHs0/Ij7mpZH3
WXzr3HkjpYbIYQVutzpzgOo5/As4iyEAv9oKzSbs0eV0/YOs8xUh054LN2Zz/d2R
lUb1sqDaffz+TKyZgGOFA1IxoTc5YUMwnBwm9Hf91PUr2nhkZLw9fmZB75U0Jxhl
oDUmnAWS4lC4Vt2+jCavP6fE2FwzeHC508CrjaNZfyg/IVpor8tQOvvFoVXRgc4h
O2JZ8XCXOYsfDkXvURzTHxYbjnqnTTx6enlHphJhP+gOdOAre1sWzzN+5Ks0aOFB
QxPtxwm6glHs9fw0iYSONIBM60IvaUK/8sq0sbekBtv1v4I+lbXt/0EmDjTjQsHL
3xYEy66JhVC2F0HWKL6MmoPVowrwQKOmE8J7dBFbS6IbVhfFbr8gESPItIO0wJzs
HfDUDSilLs06yD8B8LTUqA7NC2O6eEkDlOu1roDzXW+COoncU6tSvTNDuGS1sJmB
nYoddow0PjTp9i49FaBCzEFEvkyJ+eCifGSNjT5jAlH4IKKpz89ADhefmEh3CuP8
BFeowS/GLQ9G60XB9jPiAURvDoRpFrQerM7EZhHMwpal+Exx3aNH6iMv6GSybzKJ
PPxGjZAClcBYtEiVXvfYBxdXTgvJrTQ3+ZSUxJSP9VRtTJv1/wtg7SqT3ZvXnj9/
34WlaYQnX0hJUvBIqskL27ndSt6CE2kfUpxuKO9Bt+KDQajtlDdQH4hFZPK6qWDV
mynGuoJmhzpfKmOWEctLWKNBVntd4hQ6FpAHe/LnUpM+I2kU3U2VEhEkXqeTb7p1
YpxR9X/CTi1uNHpn8FgkhfzbwvmvxHTM6EBmlNY2nLZR4jmtm6CjpCeDvtKltj6B
8Cf9xOISMkUAICl9/r1/uMu9DoshKqk0RxCTpwqRAIsDSvxwCTkyuSOZiamrvh4N
MCV6JMtZsWaG+xNo7rG1r3M5+q16Ff72zaYSF2f3yjfTJIu3KWtsAhs+iiSv8pKR
Y3tnncyoUsPuMsW+SY+3N8OcPNIuzEJISINfVgx42adsxbpI7QK/5HgW98lkeh7A
JO9dHvFcbSR0bZ1yhjWHxdB1n9gMCGty3XqYbMmk9SbVA78ASneIQ6ZHhbUbp566
74QrFH/GkLnbN9wvTP9CdsLFtlyVzGwPsdgYaWZo1x7VERf0agOVDwk7EOGDooV9
KZKemNXSTaOdo6QpVjAxgsmWBT2k2pOf0/vj/sBMdi5BwaJ02gbqhwN0aPBYJYSA
ePwK0uNYVJ0i8Pfk/PWhRmJOX39ihi5WUU1gorE4uMbzg4YYIp7oCvhLeQlrbouH
4GP7AaQFZiwUQOF5Xrx9xrgdhW/A1Vw+q23QeQpU3XSPQDSqzLRoHpRGctw0TTqu
hDTNkXsVgD/QmmSWAT/EwLiOy+Yot4w+BnRj/Lcsz7wFpujccTqcoGEg3lmtOL8s
RpI5qjpcKWROkF1OAP95M4KW6Fyg6ukwpnbP/qkV7rnvCF7RBlSqeDF6HxwJpLtv
Y+tuX3vm6lexLGF4QrfjnlVHn5oXiZsYi5uFCvgo7Oty9GndDvexDnix1syvogy5
aDe8+XUBRudF8/8FdZE3T34Iy3B6OcojJsOdlxdOSGMvkAZDyvK4mhwQFOamOBTk
oYPcuWyBGBISsBlRu/5qMH1SiKifuU6PRQNoyKHyJC9dSi2laC3EUKMYzEjeMoF1
Quz2RfnvcFYrnqyKwP16WLV9LYqtB8F4QfmjHUpHT2oAq/G2KLCec5QQhmkxqh5U
MqzNqwbLeXyXimqwGiqI7OivfTfSP6g1tL6sK0L+t1UziSC4oczZYDnZebjsbmdS
Nc3jyazeIXi6bVMw+itIOW8T6A+61823S8XV1fua/2tkqT7iOPMFETpvdgwA7dFQ
JFq73YEPm516XVwKUv2qqKZTGGlTTPuD9uObrJZUpT7lT6xAFxYM6n4B+eoh7/vf
aJ1k6Ie+A5NxZ67BilMYyA00w8YnCHTKMSe5nMV4Dj9u60lVrbXzcIQBmfBbWE+S
jraQmyukwqkq0ZC92MLwpS2sUGeQ8l9nS7rAdyuN1gyq0p/sVd2tNZoZHp1FZoXv
SB7UFF/cM1RAK2TR9DJ/hNMvFgGKK4DFSji2x0/tBGlDShFVcbM4PWqvbqixtuzl
TMRvww+2xqW79BDGr4mwdGO7p3gmGlDe01o+LyA2rZk1nM3SRuoJ/psOXPncquTL
b7wU232pxg79y2y7ekEVMbKmnWBCDLTrFFofwvA+YiItFHfZrF4o47YBzt4OPdUI
N1I5WF9296BGbf+r8Kbxf8NrLHsHQ0Xqxv7f31EidMV5olBakLSIjZFptIqjGoby
Lw59MAChH+RzWvPtt9YRkV8vuvkWypYc0OqCzhD7T128ekEtKuY6/cHs14lyYY4l
FdIrez5/xgwjU5qmQcKdabFEc7mXLqAkSNNOjwF9CSI3JpgqxcdXqZiDKP8v7hrC
OVn+pVj0WI7E+WhuujVJOjiqgeIq5LdLejFlSwevmNdL5VVDkOsRJcqg2UwPbehg
DJ+I5th9eukHSpSo+qmM+sZGPBCubNG0Wcd0XygRAhFDSNp8p5QIi3hMIed6omck
cFuGYXwaP22oYP9ssSnVWf4w8ITBtm+QagKMcUCv0Ha3/1nX9mh1bJA+c/IQjcUc
/VIlvfN0q24T5x4Vtzp7nI67+bJ81uM72OMYTZ4SthXNUYMDrRa9V4mcqtpea5ks
kyA9doOPmIlL9iy93eCfx9Gq1lnlZzxHoHaTrvhCIRpk82nDIijyb/7pbDLqTEso
SrxfW1K7Ujja4oNF4ubzGZXbRipA68X6x5Hw1Ww+1gby9n4Tullf9fFwrh5zptvT
gGcwdTl5KxcsfMTsmIYJYRwRw8QEOspErn1Vn4gAGDkOV7/6o1q3GYTk4hoIcP4Q
ZZHNFRD45V/Dr9VEB6I01nneNNgj8oA4EXK6QDPZB31YpJ9WKjIJj7mpE2Moz9ts
qp/OJc8u3wlhLENc/AOeg/G/khPcyhpskbI7fuI9KRX1r2/kkZeAstW5KNWarcsp
hyHfLo8ksthYgT3XGzjX3JdQ4JBaVVyESq1rjt9ASeEPhpp6e6L9iz2pNdK6Tc0+
66dFO8H6b6mLoGcRp33qVmu5lqzxp/QJQLbq0Zclk3b/npwkZjgoQEkn3SJqlZ9B
ZqHuTjheFhVSazw70nl+28foVCTnQNZ/ixEel4W0QTkfDzGz/8lLA+4TlXBY7+Hu
0jqx07UNBzwYLKRw2eqtMN8n1qGRd3PotrYCmpS+vm46Y/WyU+7jYKPxClzE5JUm
I6FzaVblh7lG0nShGYE7HH7E4CxIQPwOojwfu+XXhXBzQbNb3YKGtPsJ98G486Ou
EntGyPQUH/WflG19fO5TXL8IHdnjbwpnfKfogkWanWV6RJ1YH1ggeZxNnOtgjsvp
TlRDm7A3heQszoJGhtJyJVlbikOmoMjNVCNud9bYPCyB6JxkrGq6o9ESB3RKfYEk
ScudtpNUd7n83J5hoPRij6+C4lrrApHkmQB2/qgIq/XLIgYRHW5iBVCgNYT+w8UL
wFNVnunVMelnAZ5fDp2gOhyCrzUku8xu2lTL9rWY42RWcZ+meOIhOtSSchIJDqfc
ShD68dJ0SfcqxEi71msaMR1x4xCB4fcdPtvbp/0dvZVL2eJXQs2u9XwFz0pBIMTX
+bRDH8qSTeqeHepvvwdnh9hWYHuzJqJ53Xq2pUKLtHmaqrks0fNocXTG2DNJwBeW
Ajwc2+NgMF1wwkHXobvk4X/Xf/rBPYRJjM/RKxGYB3nbEqbLT+mLmsbruEbjwm+U
Zf22bQWZRFUZYWCefXS5tXHn57yHcYvBsb8yT77TbWmU1CSiyo6xf5Pi1p23aijH
6S5AEaJPmHb6CwQOTHSHnbfM4cxO4hBmAaxsjCVmsp+JlBZMmvhCX78sIEuXw039
dBBFFFlZfeGOLZDMYkMrDyt+PQkxvzk0V/ivl4AT2mjipXefN3r8MIxd+bSZo2od
aR2sPeYltw3e+ZowFD4aj209q1t+J0m1Rbzz9XIQzI4DVw9xpbqgbZHHobxV/pcd
PIsgA1hYI/YMp+I9j0MJsxxsJhAUd7nwizrl++Mh+vTr71Y9294LjHwSjL1NCyAe
YZhPnYjV3wG4z8tWtODWIkIpfUCLrK++AoUfB82i76yIfTCU5K/+7GVxnyFgg+HY
nEmOEUDFnUsGjwDv0WKmn96ThbjQP23zjJDoe2KHXIQvtHYbxE9dsnunPKVtfHm0
Gvw8prVMAZf6Txfz9cOagApZ2cG41NNuwKnxNKmzcXK/mRizuKCqv6ARsDY4AAw3
7oW5DlOQjjrdRgryyOi9yOJwgKM30JcuPaxOs13vKSw0rxQwRvr1ZDqyPJjz/CHh
aMAfHqtZCLDVqC4rLOS/nVf0uzYpfjzXPnZ2msLgLjxItDlEdz2oIGIFEFJRG8ow
Y3GMZm0JkCTn2Koagg8HRNXpQ6MFAPpg+XWX8djfkg4HRu7mhzCI/neZMqkxx/6Z
JZSSDRIxbuZPpgorNDWYXIxsTubmXYEJDR2C44Kn6+bsUeKWOkDQQOjMdrzu1FvL
FMY8iDhtKb8dEvu1CXdm2/dIhX+a5jsw7q48jVMCvpXY92Ca+yqLAxPrNR8U5qlV
tdhnyXkh01tVO3Fn48eyj6KCyXp8929HsRl/FEVHNyUNem4ws1cFAHLoC4r7Ci7/
02pAo39WUw3dnaPbVRBkFQ8Zy/+0br6zLExOTWbzwv3X9pvngy3OxAfiegUzMY/U
1iyQJg2arTfVkonkfftmu7fEHYZ4Rx1vbaD5bDI3fBotPTRAepoKLq8YuyHvLErE
Y9SvfK+rvHDw3EDs8G65NFJAuOYuvbcG5Zod1VFRWjmxvw38dN3QYwj03ByWF55M
YvCTHrvETvVQ7W5jtH0ytJjiu3B7jzjcRri8VYfKTxNbbOYt0X2DlRH4mOU1n8c+
Km+mQbmbYYd2cOpV/IGQi7WaUfxkpvXryf7tpVcUvjF0U1gauwLsEpzalZnJ1XeH
XD8v3DyprUftSHqZPWG7kzUR5P8AnhKhHneWKncPrJDX/ErMggvhPpS2W9eEvF00
8OPxCNdO5E4eu2tefhwVbGAQd0kb/X9gGdATu4un34DlMhtYqbBm+8FQSzxTCbMY
gqolPtj2BTrBkgk23dz2lJvt76oMC26JomaA6yz0M4PM6e1BIyrMw92eVS8wkgcH
iThlLa9wGh8Ray5F1TX3MvL1Ef+hmSlSawASoaNF6a2clgsqhPaC4wZsFnWRFzLo
6E+VZEv/loZ2ptMRPeo1GC1/oOVyPO6hSw8vO6ER3O5tkLHninT5H2fQERvQxnxj
j31XmhMxeiFFrLzgMM97IciJNbho6N/znJWTkExOjfMBHI6ZWziPoMZiDq5dD6P4
Rh1Mc1y4w9a81nYIjuUo44tKUoSYVY5PnQzGn4mgUCxv8Jcf2oXfBPTgfw/p3BOX
B1m1cb6XedDkpZv8PKyVrIrh+UBUAm1riUbyBRtpPoSYym7kzmrUwqnjpWPuTP20
IC9054ZPidlrvJ8ZzDZGYNCwyPKeWGaESfLZKa7wIoTYHAIbC5ej+6de2fwcP5IF
PHcOJHLDtwgr2t/a1TE+RSkT73X8Xc5guLy9SmJXQfYEU2cBjSZnjD6laiLnBKRt
DAvc+3NiMnNr+/4AELSv4YSlxa3k9MwApbgdv/jWjCL64EULMxUZgqhqrOaI6WUj
wnYyW0/HXyB/2Ecr7z5W0GEyYkxA3KQ9q0/KrNZjJbMJoPT9lkbUSeGiiwBGHPN3
kWhBblzQdBbfoah9/sKw4wMj8p5EHb0YuPNwZoYqLXYOq1Gi59Upyw5L9yPac3rs
bHE+z6GnZ8OzFPR8HHptmju4Cl5XNvDPUJxOgqLIP8R/ftXZ94/mHhEZn8Xu3QwE
3ZeOkwKqM1xnYUhd4WJJH6l8WGq2GCcPQGaJdyOqi6Y0sBfvU9tjT8vRwuvGMn+9
j1l4U6ks7C3YfsrFryun3GXWj8YYw5x4nSW2mKzAxTA7HcgwqUu0oFpyVfNROynz
DCOiqO3Vq9TuzifNWI6vVQaJuUsiYiBB5Xq+bITjQJqy1tRK8j4xPg1SSL7WYM/v
2hjph+dROCXHsvbGG3hkTMqtEJPAJaT8s4kHxJznsAdACIOaj5ox3Z6gYc/kfFU0
T3skKEeh9LCxe9L1JZtuhm1boIOlDCnU7xiFLQgJG3/QqLBx3bECU6AL4iYsj2WJ
WcCRmuT+/QGCLpsENldSLK+kf+zQSuUTYdwu84Y78OCYPog1XMyKgGJbJ2jMxm0h
HdbFJRdgB+b5b69FHl/FbhHbsZ5B3IqHIBvx8QQl73tPYJnuAB5yzbMmMAFV1KpI
h3t0xWkpL8BlG2pf2f8tKjUgQ0U4rcxgtPT+x+N52kTvZWef7cVBu3v7n/KXHWuw
reEmUp3OZek7nrWhCyvn+2Asqi7FMLcX0r1efslO46L/ab0ylBaIu2G5eI4QSXuw
EA5v2heggr5+TsknVwBLrbx3W7wLhXT2YzeVqE4xPpszkfjV7F7sUmuZNKonRPSb
TzVbKkaJxMQzOkliD8TMWPIfqB+KUwaxexJkkeUa/n1bY2SRvl1ozhlYgkn+o6Hm
sb3FqFbcA2//pWki87V4YFJPIXcyYer/Ci57nACcQgvd1dlsMVszNMSxtQRPb7M8
WXhFOuGvOkBkuAfD3TtzJsqGBZtCjU6CH8tder2/XjpWcztv5iwQxurgWZmvHOmx
QBPRcMA0/Jr7/vAkA0p4ERCJtiMQO7f/prAVoSdyW+l5sDgz+X1xG3xnmw3z38qP
tNHNAyHTRUlgdYWrrvgxKHsSyVIQaacGCUw5cZpPSIcl571veW2ec6kYfMFkiTvA
EIMzpwykgF49tSKUvoSEierg53LO9leiweewD3WbFMQfLTcAWKtqyvvvY13Za0zx
FXQVJ5Y/9a0xXoMgD4Al94eWuN47njVC7ifB7V2uKukTVIZeEtBZlnqX9+LlsbVM
JQqdMo3WLO0fIXIFfNrwbG/ogThBkpWrTHMdBB76oQvo46QhDX7B+ZyFwQOwe1iI
xQ0VGhi7hqSRcoVKTM+KrX+BDEPCdw65+pds4I5s2ibXhLbyAL5axKLs7ELYnUi1
gzMpZRRlgtLxXoBz0fU6t3HCEw//5V5IXz257c8uJ2DJ9TETI9hp09bhpsmq/UuY
bf38n29OPVnR3/QAKv24hmkZREEBiHY2ab6RnYGcnWlJPzuv9LXbfs8+UZ7+GOqV
TJkhP94K3qbpgHi6V5bFQCpJPvm1YgjrbkX/gYfx9iZH7kWOfmUknEbVrtlIABGA
w3VpeV9ALO63dxPE+hQ3XmYIU/BUdl+3uKoRweVCA8dLnX3JZQLTfRetb49WpAEl
FZylRRYHsxc7Vu79GI+Ok/bmvhXFruG8Z8W1g2A6G63GjUm5T2w8CztahyPkKsl2
5oCQiaA3XBb9TdNBFNsWwSO7l9ILoCvTJw+aHog1to0PrbPuY20kk4V+E9EGLe8+
gU1n868kIK39xz0Uth7VV/F+VO/H3yKEz9z37rs65/vcA8DB6RCfnaNAv+9TDKbq
dzxW3U7qsW3MMX07m9Ya4ZyjGRH24DfRIfblmgstKhAPqJhp0Uocg7fNl8efwxTq
d0UYmb8QZMT0koWD2sicVd8zzR2FiUp/a020xviX2G3g2QgFZSZuapdlIvgB4dNI
jXkxnZogX7mT/G5ud/BsKCDsefJSI+F/lSNCe1M1abjufxnAXKZlm2OfKIPAwhlF
AsU2LupuosujIjV3YW0piSd1l0qAFmExN2ug82e5j3/B7zL0E1yIxyYTfQzWqToB
tqqv8YhCuzHenlUxq4p21bEkx5YHdxAkieKKq0dvZPIqQW9Q2oN/WUlX6nDogXoX
sAMVfnBnderqBNdfg29+wJYBkojbph5VwR2GuLt9RmQy+/bwT3o8Dl8R8Cr+vIPF
zCZROo3Vvc+2P9/lXCDhII02lkrUMcPMwSpWjhMePYKpqXNGLM5HkPzSH1rPjs3O
PiBYtD8iUW99FAezAJnsmMrgxEcR70z6by8UsOL3w3RUNgA2z4XeKcV5aF15dGsW
5G4cY468dDgqo7CGrG/3Zhjlq0ygKUT0wJQrLm17QBkPbZ0BYo9s0brjECiBQxZK
TjxZJhG7C/xgtoMN0wwIX3VVM++UXY3KuV8us1oei24yORgFGMWmQIo9Dp6Gi9Mj
HvMGvGN+0uMhXFq7XGMIbWHiLnP1/koANVg6d9q5sierPGayFzwzuuVDNF9YxDhx
O1HSoqc4zssnejQ2dQbi+XTh6KsEtG41eiVTBjqhtrxlkcc0PVeFXAofBDjuf/zt
D+ucZODrrVsCvBJRZ7FqPp5vFLZRomMnVQHPMh7hj9cXV17sdWN8lQMvl7xQTCgQ
1sCV16d1q+G9BeVcQcZXfvBuh1bJNaRTyDy4uGh0tdqK2iNXhCDQq/WBiVvflCV8
jkfZS01wlmaniHr/lokm5RpjWUSt30kpgpjf7AQgIls/uKqI+s+Wi5wSlaIB8yOb
v0BRUq+Dxi941/nrY82KLrkddp0xQ6p3WcIKt2oAFL8HmG6T+MxT02bmaN63kRgt
WFWIKCA2SYnr5GrqiB6tuoeTWzwJYHSwI5V4+TEKnoNkS3XmhRMcHKSPuuuNW84i
BgjR3ItYc7rL6WhfRWEzgL/NZcXUfrDYtuM0IdEitZB4ePcMhQjrmILvE+hel/XK
xKLnIX1JNmnbHeAmA4TdW919FA2+fzjoJkyOI/sGJAKwfphAzAqlgqRsVPozwdKd
M+idxaXneolDo+hMM7+ZY73T7DyaPcSn6lDgvW+k9Mi1f842XqhBj8iMK3qQqBsO
zuZDh2tXwctCgF8/7bdekQU+3q+lm1vPps1Vynakcak9vPs0TINjPtl3ac83vQDq
HMDQbTF4PMEuJU1+HbXLF3Jj6XlPZfuSH7E1AS3uX3VJRvEF6evsOJT9Ch6+nURe
S+6WZD9uq283KBENaHNPqPkwzVakzu9x7otSO/6EBt+A5xbm2SwFjXAzH3SPNdqR
aD/cza08oDkBj20bL9jIiHBF9AfdB1GJt2G9UMlokaRxp00LUCajcjxD/Kq6hIYs
kPmbuwo+BxHcfI/OILd6wOatq9VMCiS32Z/+KB9GYRqa+YvZoTf9cp1asEUGxmQm
Wd88LUJ+ANgBp1bf+/iljegkGMLH76sNtD5GwWMa4ux+j0Mmy6JTw6Be0d2PhOjk
QWVOebKwfUdKZtrHamQCS2ilRUZ6YMBXPE5058I0rq80rOZH4Ylv/Ep6+FQlc+uk
MC+pPE646SSjZ+y4bEoDnGpOgn02TIS1sK5BDI6YPPeE50G4f+DMS/gpF66ZD3tA
Rdi5cx5ugO4a+WFF54joI5Eaw1Z2rpbhiMo/gmOkjGobtPOnxUPs5Ng1SaZjJlRs
VyVm1NWhvOgl67DjASmTTZcrLFhUD3eLGNNzOyNmdFUBVNsOss1OIhDgG9TAdWqE
ibmoFVNfKvJFfmFNFhW4XIkO5RDxQa4To4vW0R58W/h68P/AJjHF5J7dvAVoUpUV
VkxPLpj4f/oEuZSZ1PZAJrTCNvl04ht8nnMfgPM7KFYAQ9wbacRzReRk2MHk8fTm
kTWB8uHJ31xxNw4DOtWtmSdsJF411sPgXUH/0Lkyxa6+z+sJmv8jGd6F0tAg5Sjk
2RYEBFJ0Y9UIc38tUnYLbpIqIDSQJvMjDr/ONKtPjBkBQpgBpKLgcZrbKZbOnBDR
CW6iv7RvMuUAjFELf2XsW59LfuSlRdfRWuJj78VyFBOii8KlPgghdIdk5Gw+MEeS
ncMtgbGA5oEl1o67WGRcWhdG+tow9mHz7v+r9r7e74CAmNx3lrXRT2u0K6EJgGQV
kXOX4OO57EU5PQ1dMcWuHnqSmByPBThoAEGoHKVvc3TTnkPl2n5ym21c67IpwKeI
S8rNlGE8ChxZbrV7N5Fg662QsgG+m6dBC3v+dcMf/3VIIk0J8q9P1fN3la17QJky
Bwtu4Lxh7iZfzsYjQ+lISp53j74GcV7ogcJmb+lLyNG3mks8aylwki9i25B7EX94
RI5cCLdUfkO6SYDo15PEK6bHY2G4+ojN7sz8xpfRijGSBI9zc+6+Mygt9jzE5wDK
+4/QLIQ9j6OUjJqeziMs3xn5NeIeJAmBcWHzolUWwOW6pFDDs3J2R2roQruBfAal
aVT6wOcLjJKCv5tukp6fSKTyH5oe1cGk45rEiIdRu3GLWu5h7g+8DwemrG9qfLtN
bCQ77Y9Pyu58d8m2M4OmIzhZM1ikAJIVKC77ZeSZVwPbXwtvM/1/i6beT1RzwyaO
aKamof1yD6zxNQbiVp9zmXcz3bVprTq07Z2qfOU+zWPwUUsx5AOoCfnA8x9b0inp
mBA+47Fc6UyPplYLpmLfSrUgcaMI6ILyYOS4MzY1+4Qw/3ND9r4I3S/AKnjQ1JHC
cZR6t6YVMfU3TruMi46WITTasVjjSvokxFhpEx+0fGbAi1buBUHmQAO51lamWYsW
VJqNCVwxK5Bj67V3i9YiaY872JV7Avm5+vezcho762CtRGyKX8qByQS5I/K//mIv
UVRTHgUAA5joTcYo1B50TTrw6nOrtX2o7/IEzglKfjS7o6t5iH3wSw0r0GEFN/IM
D20j3bomN23CI+aBdj3J/ZO3rJggtUHbaDJBHu0r/xefIoyrgIeJmT5u+kBB7SQf
PpI3R6e4XSHAP9tMSvfX66y7x/B0fNx84N7PZgk5yKjm6m/FJClCE7lBnfi4fxb4
OS+Y1UPVox1dBRUuQiwsYRnZ5dED1X599pyaxa+ls+zTWkV3VQcuUCePOgGmgWB+
ZCO7MRQTqHfk18XOrPciLE9Sa3aOd+iXkgZyk9V7jmO/f/BMut2+6kawontHaZmk
DGPPprPHJO0eP+M+BXk3Z/TXRt9MS7YJHZSZzn3vFh0KPHGl+DnSRfZRa8zSNy39
CkPhsIM47Fag2h5sz6DpxQ09njJbZ4cNYSCHp4GNDk/wc+s1F/11YtHMT9AaJMLH
QS1R0HJZ8+PTeJKN0VQrxqck9JJ9GwfQPfVv6qlfBJ75wm0kf/MsU6eWy1uBld5w
AgQzTmKu4MkJICCZcIUmINLfftek1BNxyTeRE7gOPzrj5NtfOgrE4QV2T+tSZjQI
phx4RaA9w9crHgtbdLSK3KKuAbsUfi96nwI6obxNXx/wBGk7lcikA/Ftd43KN0wu
CPwrskr2OCwo5xaEEK/FEpHvR5dpz6AdRoKZPIXhsxMYmgwsn4khg+yIjaXswCSQ
EbzAJdvDZhw+2HO9dyhOs/1rUzNsInsaBODbH5VnvEn6ftxJWkHsqO8QXHeGfUmY
FDPHO1GGkuyIAlr2wErwrBCh/VATPuP991twTqd59lu/i/R1vjcOySaCFPPFguib
0nC6yOdaHLeMULkf+PL7Gr7obZhkA53Dg0us2HVRgP1Gss7m23VXPO6AQ8aMfbSl
vqN39m6aTq0TguYkRgAqm4LGI9fhU+W5DJGXF2Ycf1V59SapUixSNjGdvn92y5QN
bDtFKmotOtYrmnbHR6Eo3KPIBPxUMkYTPv5xo4pRiihTArebb5D7Weetd1nSFuys
eqvhluUn1zFcFM9KFLQ9tC+SSrWwMya+5uxWUIzs4C6vmZCh3Nec2X5MjtKet0pU
T97byrHKI6AXjDP3nHm2M+c117ADgpLCURs89cjh/7KKYR+dJRHgk+Q4ZzglUZUX
lJesgx3fCeDIDWRJsOLkOa9H8sfE4syKMB5Rf8DTz2tU3UUaNKBGDG9FYEkRmbm8
/HvoDjvCVu9OI+Eq9k/TQFW1ADG266pxoSea3VobflFoGMEulOCpW8ZVNxiZvo53
z3kBnB0Ol5wYI9pr8EFlkGg47W/JNedvEbz7ZnZ6xsmodDWLpbIeOzxTpYvUH5lt
L6WEZmFenviTyyKfuQp/rW2CT/fHInCpeiIMvu51pUfnlH7zN9AoF5/Qxv9rBzrM
UiDqWhV02ETWjikCkwxSaAbk3t8+pe5fSI9qI7M5Z/kvUZpE3eBDPP2A3XuXIoxN
qTCS7jDDJRlBkUoKgkEGlimAtiOdUJsjuIpMyqvb0T2gZM/CZcbTSTkv1u6M+Rd7
iz44fcodfK1BYSKtBTgcpA2INA/BfkrWGngihK2Y6nrPEBAzw2CRtDydU7eaFnbs
LCz2UCJkL11cmLgpBfYPVDJzk1obZtCX6FUexafnSeROJC4eUTGF2ikq4RRVJPyG
rxxbCJkAiEdELEC0GaEVGcA5oFIZi94komtMU6OCxbbxUpWi7SiooRjJWCFP2qqo
o50aByNSsc5vjxROoQ8zuZoMnMi79C0xKyPsL/pwNyGSrAJWnomCoH/DOm0rg3ky
czn+yqgymMZNQYf8QQH/A0NmwfGXoJ4sy3VJ6kw61WAxvLmmlkt72rgSfgYZB/ny
Nir0ssD1MyE3ZsklawsTfqo/XWxDuuJr2mhXWleIZ/n4JInNHFcnqqWT5TqypGWq
UigMhOtzwetvK2TKiao1UzFqvU7vomBOTk+Gk+EdGvXPU8pjsI2Crh4xcZIpXTT6
txfwQ9IP7o9Xp/BOwBSp8KJKOR1Lq8+1Q3W+eSAdN4z+jSEfUHORIj1fAdSLw8KQ
qndAjReIrIsTJm9ydY7Zdjdy5t9UtOJjiGrJOgxEZJXoiLgIbFHOPvJ2zyWN2M+p
3DVJzv9SMN1O+mPPhl68z/R35dpjpC1lOTniX3YTq371JGT9e9ODd5KOjIko2fo/
XIAE238pW2qKpjZ6OGpR0hRKtegjtY2TOXEU0gzXc2Ik7Z8CCJR4yEV3ijSEsV83
lw6KDdQX07QbGDMS///L7Xcess5PcNMMJXxDF7W6ulfFME6NOnEkNjLtgSNI0igr
VgredRBjENwqnrRU96vsOzKCpC2ny6MFsTgqHK89A2bXlo7pyvx/UGnDnjdCqzaQ
1rrNBppbzp6aqp/WWJmzcMiWxbDX9mBbqiovkKd1heKPE4oeZ2+O0HXwDB3XHyxI
tDc+JcuOvAqQznHMLARjDpDMSfQBO3xc67cVcVmPVIx5SUnjYrOyERVvNyFWdxZA
sweaExUzYZxa0iZWS5v4SFAII4Ye26/I17WJl7fuNiu4gsaH3p3THKNZbQCE5Hc1
dflz5gQSFimOy+DBEotrXSH/2SvrepMBzsXY1eCzDR3+Py9XHI6CcN4oUpSCZP4Z
oKerhY5bLi2GTK51cQEAES/Ufk4rx97Gx5B5HiT33AG9SqXtDACNL5tDQrq589mb
UtNJzd9Ewl14PyHlz1vmSIPaXzSGM5H1LZm1NHdRDodquNrHDsw6HjdrHwfK0u+M
NazyyAkyYsfO/toOqq0Rs6J4yWWXpMdGKzPYUDkEqwHK2G7YAt5hzCNW1OAKr+0S
+u7IvnGlpKc+6Ngs4DKEyuuEt3kH59PLcZpvI4q8lt1m7BImUuxORjUnDlS5CrT7
KTVoPQeN0JQjLvNUooSW220m+9QpxyILhpIrjw1Oa/NP8Lg5l3cX0tyYtlKiH3ZS
KKOIkdaF4riIciq3j99N88LwBshy+Ib+87EPSGyxkXp55ByqODQM8OdnxQZmHSdq
dqT0MzY5p7D3hMCinyli5rjxArz4znGczDeia5EK1ZLucsZtMfPrUMOlorYUouKQ
yPLwrJsiazzyPJhKf9uy/cQ2bphmqKuzgHrhDl+ren+Qv6y00vul2FazCcNt4Ckn
hYKFWxBKedUZUGyvzXZqxouKKUmL7fMFj1N2D/Az/24JkZrBD5c+gH/Hf8BEeLLY
F08kfPXC9Ubt5SmrrKLOu8yseeioO7DLIPZrOwYFWN4Rd0JAIkVBdnsCPeLEtIAi
so73+UToTTDxaCAO9UoOJujqQkp0Vwwv2Af7fhxswxoO9a//ala7dj6yG9fCi33n
79cpEOkTwyR0gL79FPLpjkDESYLR6JEw2yCIftOWrE34HdPKKrW5J+XieOPntQlh
6ha8OXuMrGDPg2o36mioBrxQbzOzSYHSeLmTTMGjZjoG4httl7L7jJqeZdhJKMce
taoLvoh8NVPX5m1ZaAzEXVx68+/Tvtx54dfdmgqeM710PudKF4gSWSq//7n1rD7l
G82ZGFfT1plngZYo+r2XIcxVnTBCNb9w9KsUD5EcxUwWi21q5PO4uRzTKRZnLzZQ
O0k+HX5P5CHoLkQM3b13YaLXs8cl1vfTVgE2tEOsj9VWAQnXpBuxSZSqljd3EIdS
ZPO+3zMMAte6uDmIQ1Id1yx3c3+2+BLIQQ3OYodgo4F78XoD7/enEqpNWRAjVNju
w6zTfUvIzF+4zrmp+D/OoNehDQbbdkQUe6eC6zbOAd+vVckGVOls7vA/HIdyct+1
74N7MkdtAcRsm0Z/ZxUUGJlD8AaX5PJ3UZ227CPNvzbkuvmy9IpjPfvQjgK+kLpI
TbGRAPz/r7c8D+WjH7TpJ5C2XUoxb2+AeaevRXzb+ZnkboX8LMFgoyyYJ87nUma3
e5KvzAw4rpfK+byvO7/fIXwpVqIa8cq2+bm+hl0TWOIi1LugV8Ucvi2F8MgaaQJ6
3xip6ZyM0P8VS+rMT00cWihREHLIl0Q2dwLvHn6qEuf4ywlWAbUNkCpsTTATOyVX
phR5GGiA8Zz/msxAZnTvwKeShf/cftxh522QLlKQgd7bCRt3bD+3XmUst1CiWZsg
yq+v0FrLGAqArqzGCqV8jeghl5giXDsArRsNvLB8FQY/jBlCVcEO7pZzW1Tvw8dd
ZQJ3pBLKPDMFG/508NuKtDEOLbw1pdFg7fNilCOCyHqKZF/THl7CYfTtPjHNdMZ6
q8Q7z+hiRszLqxQf+2LY1u/BaQbDVaPHv31sY6Jld7T5cLlt0i/wMQ4SI/lOQPZp
shxKAOQFzwM1wKlED1DZ339w9vqOdqM6R3svSeGixQB+PP0mAN+Z7pzCdMJPPxAR
FerBIH0rJ33mmP9uo07rWl9h1dzZ8y911EwGtczFCdNzyNgzOC+cl+i2icHNP1Tw
CsRM3jLm6v4+DcFvtrir6kymnwOnbyDDWFrobmVAVwQ96J46CQbSaOTQfw1gyY2U
g0EIbwjQnT3YmpinhhBUGKQwczai0wio1WG01PtyQv9xtB9Toh8CcUMKkKWxoTMO
L9D/QBhYzjz5COCvEFtp7aVtQgavNUTCokDDb7/w8eQSqY6sT7sF4EenXNSsmdlR
PcU9R+NIu1aLo6/JvfbouH3OxoI9M1i91KUuTRN70xTikCD+0Z2XPrtiX3DfrRzP
pL/gsudktZw+YKBhwLKrSHWQbYfr8W3wzkgayua13oCiU9FX9l1doyIyF51euMWj
ZFMNujcFRqNPxkLWclEjRpWlRQVZeZHZ8xxBhPhdm+H/eAEX3jET8Hs32F/BRs8G
13BS8nZfK5A5bzQLLqIqYY/smylZZq1MkeSAmntaEAzNFUUuYS6AOB+0EjkSMdUb
igAbcCti93aexuw9wvaVInCGdI9eA2rkThhEN56uAHjLihDuRqs1NKq11tbPIvon
j1DNA2P3YZa+CDY7pj2k4o93q1f1pTcAHkJTMXa7kHPZ0U33z+Rh7RSDZY7rKjWd
LEZInm1dLTDoblE40k0OROJCrgRnJE3j9k7/387oQJUCcO+3dwrXV8QmE+hKahEu
UWRP3LxU8mub2hal1kba1efWt3VaGC5EZH64xRwU0nPyvWF8mgMmkjhUX/g2U79C
oSEVf95tlAfys2X9tm4BjO6rYckpbRE7OElmLL39dHVEqAJrEjeefJzRBJwGg6C9
T1vNHAMzMFKSAbTppz7i34Oe3Kgr3GEK58LlMLqxEjwwY9tL2w9UY2GSu1C1Lm6B
NVX43gDtGLjb8HW+rhC0bC2b0Gsdyzdh+3Tv69cWsD8f83z33akicmHXKLkQKPnc
ts35rLhoECk7sKmRBZ03JbVYP/jLhNj2FDvh+kuQwJ6FINqnOdrLeZGcEvgVpCYY
LvRlfAFlR4LDK7k7LaJeehiiY392b9N6a3uLeo6pRKSbnQANbV/pUTer7VqPe8Xi
8wGvFMocoeaKUI7Wl2UIkTrikDCalk+BliReyk7AQQnAGVQdtHrDUEadKa4KFEtY
bTqB3MCP2C2D2STMHW0E4akPgmRmv1/6YtfILNyKfk8gLZ2v4OmvaB9yL5VfawC9
VNZl/Dy0TairOBQoUdCIA/knsjHZlDL1KhAyve3RXbAoccdwuSk2B+EfuIoWcFRG
t3um5suJgBbRvcujIbAxPwcINh/eNdhoL0akuoPXVnCjLc3gt1tm2sYGG3rjOKS/
sJyyX3DpmXEExrNiLZ15Dt1BC6qDJot5LwLLnRl1iUEkB8eUifHs1UR6fkDqTsQm
8RS/YlZiTatHsVcC/XPjTKWRDqYipgyebMyaGySohoILm2L4oCMS417RmmK/0DNN
ne6RjSAFQPC8xSCRf9w98AzMwpEyELnsznltrrQDIF2hLWpB88lqFrdrpj/yJvgN
AXeAJkzl9+y653GMb7TJNGX7sEHlMciNcE2BS4/i7aeLvhisRT1ADvrLGDDyQM7Z
wbUzKQqrrDSOQSW6HQFQw2IChGLhCQjj2I8k/DJ/beYoITKx4hOS14aUJL6N2SwJ
1sRgrxcvdSRwPuSN8oMkOUCr3XTUSJCKmPZ6k3AfVUsBFCDOLzi/LvlJJrN7FreN
PhtZJ8MZgwN8hKPSWSE8No8NZ+MDWENZuFsr/j+PboaLdIddaIhKJu7CaDhfjk1Z
RP0YJa8fsxBRh100RMwnZuP+QeuB+MHSRxCDV8d4NiwAKFBcyllyR0vwDyR4NdbO
ARxNEfxyLEWoBImiTk2dqbvxm9q8WfMlqr/EZiwkAxieoh5hb+GOrAQbdRxSZ3xJ
CKjMPUuwZNBhqmCUSE7zFekSD+3A39l1VhnFMbRwZUBGcOm0x4f+jrhRCmrPt+LX
KnKna9QQZD3KHKvnn1lMhAA6zdRnhttxrHlBKO3RsLJi9kdnCAxK1dlgd22KKyCI
KQgk1vkqFX1YrYb8pfHuoYXeUJ2KqpssgynpDMjfTc4sSlW6N+TVv5qsPJWWCKhy
O0SNGwRXuIRYIqaZ6zSe/NDhK5WOEExkxE16CRYunjETA5BEVca2vvgG2FaETIuB
cFaLrtALTyBT1WoBYMN0vrfhOikg804rOMXsZSKqZiMo1h/2SDntFtyV8j+3iIRm
tYrRj5ecpAQENhcUs+g89KAqy8pHGInQQxTic6uP/xKKnSJ/zZwHlNcT9knleFiM
cyGgaCeZC68j6wmiAbjPn98UiKYc6fApSrVdn1rC88yo3Tf+WW8Th7HJ+JcrfoNG
VAgONEAK0JQP5SHUbwU3ND4jULb3N1FfRiqRRvGAIT/ktr5RTS0wWLiyz480Dk8M
OjtPlGXV0KQMu6QcpODiicLlJ1EswxIrprC/GusnTr+hPqqzqcQGor0iUMIuxB6b
e7GI19nALsNPtRgiMFwqksmgUwFRswwuZ/gcfrsGLTzsfLcvwRHREk98nJYl8kQz
v88yvcwDt/M+Wb6VxzNIimR4qCdsn6Bluh7NgcOsKjC+zG0JMApba3KS46GvbXLS
hhd+8u69c6D8nKBUorEQkRZXGqf/j0yQtWoXxcbTECLiT4i7l8mxruuw6jWiqHQ+
vbeTrm9qbhEbi481ZtDtlQeSqVLxsXi2svZQM0Wbl97x7KIPsk8ZRCPxdf8YipjV
Y0mW2a/ZXBCc7ehxuv1VyI+DKwE1ZHAv11XSEKcfD7wJxApbQxiASwUIZrdOvBKx
w85pL12RekuJGra79dFYtJPV+HvMf8XM4CIA5fZ3cEgqOD2M8yF7llJv2Fcr0uLM
EZbu8HIrdQZzgMyloSK/hB0gk7U62wR95XHx3NA8KjMAsoPb0guag6GLwA4XUhqw
ZwV7xbYbzggMCX1EMXdq/mb8MRSwufCSncNFOZrtmjlFxmMj/s4nZz3FYt+hUPAf
aVat9kStEzOJ2JK+6aAgEl4EL29E1XFPN5L9T1U8OrDtsh7GHNrqiAXRlLS3Gvrs
mlp0NtOD8II7HxfEo8YlylYsozz1BOV85LuwrMdyUANV9nbAy+7AGPbACYoaLwEN
tZIT4aI8h7dbyc70+ADuVa5OnPP4nBZ3+zIlZVjIfpxWDsqc8hv93sgXxvM2lfU1
CMdJ0ryKCslObp/1H4HpGl81Z9Pn4HPflepsMYO/Ya8hFRV14p26alPiozMA23X6
vpS+MzVhzxGxcdO4MplJrqmNwIk/OgqsLDy0zzIX0diBZkC8J1Aa2Kf7jBlGQ3i1
IkIrh8r+0C/xgIB5Z+A9eUXvBoB3fkzL5sa19FStCMGd4locTZAJSfTlJH+1/RIu
qtJ8KqVMUpvA0SRBzcVLtXUY5d5TTVoL4gPMDwWqVVw+veSZSjNsNt4fhlcDMIgD
aKipWwM80O/cbvQHdahz7tr3g9PjMfaDP+1fJMv/OPT+nlZFVHJobLW9WpJXNY5n
ahAbYJmw3b0MF/WtKXpr7DS7F5d5qRzkKgFP8wWcVGPa4x1YcZgW8QVt7KZm4r8t
Feu6FygwBXfyo30EKGMtEJhLjsxB8fFEjLOefD48VTiul36EepBKdjaEggJnizy0
8MjI5Vcs4nXN+cP325kfepbb5ZXGc79R6cDJJ90TnPQhECwamFC1Xd94kgT7EpIH
b3t/P5+arFAFMXNx/AbYtkPPn6YyPzc5EDqFqD8w5/U1Bw0lC2sBmCRpGDTEHJdX
ntdUFpnzG/BMCRKkJEEoHRchBncf2o2huFAcr95CgG0SqM76Jb6Zbg5Mm0g06RXr
Lo0SpHfaGFijg1GeNW31h/8aysc8e+zqSz3TlEKRZsYFbKkVDxtQqn9WHk96zZnj
gszX0/MbXpn3M2kpjv/Hzu3HuSPyVpma9gu7CANoTeHm7yBGtawWLSQaGYJheWx4
wpcdjebCgjJRhXRNpUVKNJ52pC7EUnazul3nFnuPuy6hoAc3QOUizI37a5dnqguv
UfaX7oCvt2wSNQBdInj4Ba/5FCsAMZ3tJ4yyNSd6EVGkuFEaHSaC6l75EFvLtLPu
yeetKVtctQ5sMIghswsJfW9BSV0HM7LJBHK3EwmG2kvySJlCCSDj+S5Eoj7L6qMI
WRjcbnd8VTTGcXZMjCN/fIg0f15DGFT+oLKVjp3GEW2T1JDJuVKSkIwdDw9MqaPv
scpzahaM07TG2zO4Hx5VDI0Q/t5xAss2sZ06hGxlPi89jtaZBvLJwoVyUJrE6/cm
0tx++fJN28ZyK1Ms9sN7/TtQAEv8mkwcV44F7j66c6pdyDWddAKDkBNOUUcD5uUk
BAFNd08Irrr0tt7AG6x0gDl8G5UbGDuQlydEXwa4dfYdKoC57eY298JWBCrcqisB
+dKhBNVAj8s9m3lAmlRWtzEFr7gTIAjV6CVPeU2Kz61EwjHDWDXMAkVzB3772VAe
JKjSRxaw0/UHT6KSVuCEdfKDTaFMs+/EdApKnJBeLTQ4r5D+YhAbWwxHFuAr8d2x
ZsF9Y9MOR4IZ5nvAfbteXtvIl0aHZ7sTQ93AmZUDDQG37NpcPp8ogrYJ+ENiTZff
4CTLZa+VlolhU7JRRhLmRe7GxbxxYU69gbrrtKhiCQW96IjwNsedq5YOnEC9avr/
LFpcuQQCbl4/t9e8bZSIc/QHmpmnSRV4KbNABDlAL/I72SSGa56O6//ByH6EggKg
ABnQtH5C+chpiUl5NCIR0+A6b5VUKr8Lgdk+R/AVO/UeyzhtinGEs6pNH/xeNs0w
uDe8OtOH2/nUPl24cyW/tG1ZogpfHXeILv0/hBG9gpIEZ7ISjUrbJg/4srl+el5H
fQFAzB9ffxguykaKQw6RW6x3dFbM//inV9IcxnSFsRgXLbrYGHVKZH3m9kKvq3v8
eCByiZZaVnOZg+WC2+TxVJomgVP280rqJj0ppjqMFxkfl0yaEX1f3lzutVgMXmMj
QYashMlQvIzUvK9CjMraZcHFcHb4/sFKe8+ewKedCV53FzfEwXCnJpq2r0agY2q2
E/7SymJpxZ+hs9dHv7Csk72zTGxIEg+sd8sWMA0tt8gvPEWCDpU1a9pCcw7Pjf9N
4YuLYkuZrWYU9brnIeOcoKqm7jiRrMjBojEaV3Q8onYQBZlGkzWj8fhVGTrCZ0ur
eSH8OcxNAMH+upbv6PkuIwYUJL2ymBX7JBI65OQa6C/gJe3H9w0aC8dCU87tRoub
WyerdVUq/glEsuTE6GdA1JOmZPP74ddfMVopkuuQhf5yN8prfU709c4jr305fPQh
k95l4+HhE/cxh8Xa6b5sED0wcsSHV7fF/fz8ZXfKxb00AgFVFI1rDPbH8ZDWzJv6
m54x8EuWeDYcEit40NqZ2lmQnbz5CNIBvET7WrNxO++a1rO2BTRx3unCH2IyHIK9
x6RxOxlsQZxsMtlpoV1Sp26SC04kgOWxfYEM1LqjglQ03nyaY5pYksgh+V2Q+lGk
EiUbIBFM2yDqPJa6sEkiuwLlcWFgf2wcMLUwJ7Y6qMztNFuToSY9xK5fwHXsF89m
LaGTzxJk6MJbmXMMekVVbvEgbd/2wSlT7Ur59V9J2Lq8tecRor7M0SJ7uil9y3Vs
ev6XFC1wtJoclA+rjrSkQYYdwJPFxT84o/L83a0L5yTDKBa3SpUSQRxY45LulZ9f
mUow5et3fTdR7muSa/ugELeYl+lgsRKxRC3JJOcrMu3X6i9LLQ/YbN1OflFsW5hO
FDIO8m33bSvHaJbrICoryo0JXMfVVO4q/mglPWgt8m4eyXUceGebducJVyF2WCRn
2uE7Y0ellO8rbQv94iF4L/zey6bODn4umV59uakyZd88rfp5CJU8GAUcSqZW+l4g
9/uJ+S+WAYkXzg4GIg2wvKVmgqcdpqLG3VnHXM4z9HXfaT3AgUyMKPGAyhrK7Gqi
3NcF6BxrYGzD02Q2W45rjMQ+R8jg8fMRWrK7+yuNTjDgwRpdjPrYl92n/d9FuavS
SUVkM1Xczx6wDXS0tQq4tpAGtkE6d4T+WOPKH5YiVrQNUrnbIi7DDotc8DTkQpki
2BHv0EHQueMAdHX/nvYnViU3O0h7z1pAO33DcOqkJyOdc46DhwYSXwcmwIXi4JEb
waQCRRG0H+bXkXWXjAhogbyCFT79qiYG0x2QFJY2PfLK/CXpungPOYtKqrs1rkJ8
o+6dzemQDbPmrItVwjm2XDnowSiUjVVSKRsH6bP6vq92NQIF30sx4tvwQG+htvij
NqK3um5BQHLxaeeCpkDReW/iw6hVIaKVk4j6bJQ14yBAwxS9pxAYq7KmXnCKVdXy
lKR+lY32WfU15+rSGJFrl4Qrxde6QnE6liNXpL1Eqr7IFDbNxGfdaoPNbjgDk//G
odsjY/NdXotD5eZcThcrifC38h3DbniKzzjFlhQXLlClvPOoXz3g8vRC+jCudu1i
vgiblL2i9LL8GX/2TSFGx/pcP58UHw6EPnBWTCWMiTgVnEPLp8TCW7vWYhYEVpoY
ev1yag7aM6DT6WBszjECJw6oCBmwmx2aEO8a+vLpiKKfuyvX46CY5CDT0kYs+oes
hX77Hf/qLhdN8heaKXczU6oxmLIXJr/E9f9Js/O5ocHhGFn+r36iK4iGm8ka9k+C
i/uC2dL9OHnVdrNpndkl10B+livEM/ZbWV7dgVHXkprO/NK5AXoyoGKJTK0wGqub
4vLikfVpF4R9yuVonBGBO+DlntQ8vJD24iVK0hcIf8Zi9U21Pv6WHj7fN6S03Ajq
sPFDA8NUmVFC8xUHMWBc97w/YWLac5pF20bDvf3fCyFLv4Ir454o6fIULNQ/PgQM
qm/hAcT+O17+aTTZzwu50oVjz6niyMZQcndeBdCMEXxnb5lpRZPNmS5g7XDgSVmM
gXUoFs0drNzggZrO2nfHIOH2xLAUfjslJbtcmYWTnn4Czaq2AO7xWt6uGHPFmjxc
H7JeNcvqwrUggzjGCkk/k/ZrHjN8mgIvUHPudPo7QQYjp+TeLeyVv7XWBZjxjkd2
RARxgmNB9yZvrWz59Ixct9/cw1CB/NNZdpYymuxnFhqajUUni/+LTkJ9kQ1lkBYJ
CSPKxb+8YqxNfn+YNaaLBIvhj0RJumduDxInJ8QYzDrYHGpn8w7D8s4V9s2T86CX
LWFswVstpTKak6lE0XGxrxuzec2C5orpyAu/DkxUJrisorZa3nKmU4e+7bvD8qN6
YLWNgEAZxsOmZqONMOTJuYN++nbRbROPy8Q7MYpzFogvWAnKei3Z79MqVNy0B7ZB
WTJ26tk+J4VDh63B3piWruI1977HI7MedR/cjkYQJuB7odWrXUWbX/Ghcs2yQI5p
Fjpzu57YnmSshZ5+qjRsmOVJIBqZnsNkjuzb6Yv83ZAHdRqqaZTdbopGAHxocXhJ
+VVRcgnD40z9um/tjOHqQgptnUkyzXi3yJEdW4Y3mvx1eh9vgr+sO32KdJwZt7UK
JxeLcFX756Ka6cT50H2bd+LqwCm50nDbmA/Ut2Nnpkvdvix6L4MMRSO0ZwB6106n
UMdlsiBVAoKWDV/NnUSkhAHjSUiH0xDVeFJ2mRK7YTP/jekBTtximQkZFVg5MlGk
hTpAKm5qMgJPjnJGuGyIWGK3XqXmh7qsBaX2luaonVuTMlAs+VUurVp3lDzzmNeb
NQbbpAYCcBPM+eTgSXKlZPaDKLTC83pBmFTa2TlZz9O8JFa5l9vaz4k9UuW7Hqez
nt5M0aNQrCFZQxt9P2A7e8GJCYA1zPzPhBGKC7b3SV2wTU1CwISpBKyieuQukBN6
9SUv+cQWVM80gBELZxy2yg+Ufjq14XWHvCxmvwFLEbEOfLmBENTMf73VY63cm65F
aapBtThJ7uJN8IokB3afqbbfEK1Ay/vFkAUH4bAiAQPa6yYda1lBehqbecE8dat7
pAYhbCyBayVUf4garnBx7SMu0e4InHWqEtC6ASeKMWHXwtrbghojjGDcrpb29z2l
5gbcj6Zl4oDOLl5pgTKhCfvw5edO0opJFF/rLzdSKVADoI8tsJydb+mHAYgpNohm
SSkhHWLwa6YW8wEGv0hJM65TDnHo8Kv2NY2+J4z4YBZezt7SskjuD/Ti7j7D/nuH
UXz/HVsuMUTGDrMnnMvOtFlarq2ughM9lGAVp3emCbqKkk0pJdLDICeptNHvl1ZE
1Qlm01sARcXE7QCGGeEMrFWLgFcToKaElZoo0AEwNV82z6HOkhlqGcfopUQ2aSDr
LUWgqqNkPP3uT+sMNu5lN7vZ6qDRwWCmgpv3ZAFtuDLBCB915XKnbQDOGihju1U4
I/zxtd7O9nzCmj+Bw5UlSmy9nhCQ63R/Z3OTAyyZwHTFRjhGsX2V8jvJQ7fPI9p7
14kq3oHN67MGXDt8JYfvzUpFGgbTd6EJZm7ZaU85ZgxuB37soklh+khfpXQRG4LX
0Po/128+R08EtBO3hgQuYb/Ag3ewoUwp5qLCi3nLz7BZQIP4ROgqvcsOOTaxcYc7
s6gAUjhBF5wmwpnsYup6gN+gdddBdpmIOQ1pITdJJunDkUCqvqy+2eCR8rcbk8CB
0JLNjQwoPZuHd1osw+oBy36YTCJsz/QXPt4GTIH7NWJ5Jr/Vo5CT06IbIS2PnXv8
lkNiLGBmpJL0SjiVTVxeA7M1JnRnT4BEeFMhzk3XP2YtblymFneWsxWOW48bXrPS
dWEZAx6nQ1y28vA1dopa7PW3cmrlOVnWBSdrVP3jWYLTj8AtHIStdHbfPiYsLjHi
2YU/6UMtOAbtkqfNXLieIustdQRkU5AHO4RLup5/IR4Xzh35yp/GfMqND4WR1KwQ
Uxq7GPfVfYu2+MSudENHXTjWwcpQgzDXnpXuOWd5LllcTv9gGkn09F0uXMkmNUVX
Qvo1vKpecv2dAxcYe+YqXRQPrWmNJyiq5xGzvxyBYwMbnTTIVBkV+LLUs/wW3/1o
Teyp4HeTrCT1UKR98mD4yZxW6WuhGQS3/rrW10givDkM8N5hkRXWr51bl0pi6+Q2
koqNIySmbmuuyTM5mpUzaNX+t5IprYPJvWpVQd1cNhBcajmogHRMsCe9ZzIurxXn
J4RAE8vkRhpgj+jfnm6KUg6R/na0m3IBY8DOMJ5psaE79GM+o9OMGBEswSwml9Pf
oAbtyN3NA8uHuE87T5b4GyNqcJMmDjfYlSRirMD0SaSAub9lE/PhFn4Cp3mgVo9e
cw2TTKz7o0hkCeSiyYvOYDqNl5T6xLxZNAu7GyOlkqsiC6eZc0D6lLFnZ92CkL9K
okVQbAdpvYPV4+C+rtQCbGDXJjggLEOLAJPtT60GBBrET9UMWcC7cjgExzkS+qyc
Mpj4tVEh5vxTJMWrH1NPPZcjpK5mkcLgF5Q3QxBwNkSPQKHjf3t3kL1TTZ9eVLxR
RZWca3Xk+/cINRBumb1u0O90j5X2bTNVDSz+PQp1ZByu0PnzyIySfNn4IKpXA+Ku
Z6rKh0Fn+lHWaP14yTECCsHRNFusceCyWl7Km2sZl3L5H12/1UU8WSRR7RzKLIUL
iTpw6TBUR0gOKI7cyDBABPS8IKnNzxhvkC9IBSGfgXMwcvi0MWwtfYcKhr+u42eD
066jY9layu4s9W41NsmxW/0hgB/PJEnQhvvVVoqtwsyI+TECTUy0y3+8vOHqQyNg
HEUINa15WExkj1D3lBCzhQbuZUKsQ9gA/EHjFgYjZHlGchlbBl1R9pmDCA1+ghuk
yZeDxlIFQL9xJPsSADDgw7sAR3WXeBB6d6lryuqvlR4CgXTgS3NW/qk0DE2sFuze
ohriutFFlkjLJv2GWIpqswRVrSZtNJMXEKWDhLcDlqQaUXr2QsDxkLysoEoaDseL
OkSIba/cnpYKAG2I02EH1wwCgh94zws5zRsFmJLYEv7lkt/5qDOwt7Is0mgVlf0w
OAEeyumTJdtTKAp3ywW4RZY3URBKeuzNp1H+AVJsPUSfJCk6i7pwkIqMrx/9HT3/
85d02XDMLGUsas/TrQVMBHcEljVdz5AOxopb0QYGcRYkW3osfmjv3RXeolF4b4RC
IYXvncKuaK/AwxFqxN2L9vCkRnAC0r38Dw5S9zf2Z063LOhCTlWomR3aMUJ2Zj/L
4RF76BRwt1LmQdOztIQkExCpbUQPs9aez/mcWqheHsjJp+hWs0SZu2gc0qnolUca
Fi2jU3XpfSfgmv6PEk528L3i52tRGA5R/ipblL87kmWBW+pZe79dCDHPiyJRwo0H
pft0pV9y/Sp5r3TNV/scvKcTeQclLvsAxl4H+eBT8uyURjpUh2gc13VTOrdECakc
VopfktBWCWbHiOuFxfBFq17Iv8vWtH+jR70sh+Lm5W8i131SOjKg3nWjLCmspPZq
pktfSn2bg7G+lk8B9Eo5yt76kxfCQ+cwail7T5bEHgARhUpfYdHNc6L2ecAw0+tT
lkMZrcVqielvGTG1etIaYCb8uxIeXtCgy97DiI2gvjjEFzwx+XUpDxuNPIz6g5gB
KQ794S0/7RB1TYERKvqox3nr86tZ34qUp4pO+36k28s4YeSMidhcpBokaOkx1Ed3
2xV88okvL2znilaCYsZyfFX+gg77pEG0hui18lmD89xOTRyPOhhjepMf8A+MDB7a
dMDLSg4souAM6fzCX5+El4rV1Pfk29ybX/tiBTqFXRycy/s+bP7vM+eJlSlyiw6p
TqTU1dyAAzH++5uC6q89T+4eZN37QsEv9t5+g4JdDDF/O+o8TJR9Yrf19zePbn5F
ZYi3vwXTqVyXvWjcq/dKHhTJenczmGgkhxdrP7J7823mRhilYOe+/8l2TIDfm+HQ
woVT5kL80kcz+6NcpK8SXHyP15Rbyodb3qlu8h2AovxqQryhWiSFl5Q3We6ummn3
MnXIUFiZufcCrsBuHm67LWEsq5A4O8H148VLA3AIUnKba3WNS+qQxUmZfHYDVawH
41go1bQAMItDkOqzZ2D3C4qfQ3+fl3We3LFmBg8JBV5APl3R6Zh+KswuYXyZpgvw
Hoj5OIwTGVczzjQhr9LKkrYzXJoDKmOZDbmUdvDoUoiUWIN/O1ndQOuJ0Ep4t/Le
xHw9VmF+9bUI7rDuuinOSZ+8Jlg/FEEYsSPRvAWqyCIl9KtCK5XEZLF0L/ZlQaNG
o0Lhvy6US1S5K46VI8S29Zx19s7G4jc2xvLXwfYTzViZtgFNQfIiRXXnHZwKNsA6
BAN85Zq9uwMxxtu8FtQ2DJ74gEWInHXlQg/KFVBo80WjeIg4U4xhGAhxO5ROhJ9M
GecwSLibV07QfGWgi0IgK0LoUO8QocXHx8oMrRJfbZnSUrvj/odPvEYs1WBuD9T6
L7ZRVgpfYskmsz0tBfYgoyhuh02lOUjmwUCgS6DqYHemDmAD8nBbOjXLqKHkY2aF
gLBOpFziQrmTtoHmPFceV7gIgipCn8GsBhxVe+qUyEpnuDfKGaoPuReg6ujaKnrg
P9p3EuA9F+R99t2SbllkYMJjmN+lKClFPADcHZMToMVYwm6nOyQD17ovZLn/XAB1
VgOq9nDKCWVg0vwyTJSh1Codfjn+R7SPNrbkJ3PdS0AmZR9QVhckBIwwM28Oc6f2
HjSSPSXu0uM9yyocpfw0MQCQuzOnwWvqLDhH5tAZuAE4ioFMIp7IyIHahhlPFLss
tZZt/F4xahcqjrAXIcJTymutCb7j6kjE3WRliG1sZyDYZ2ybZxno6K3yWlNGmLeB
7FIIUhha2jbXQQqAsj8c81PLAgdGwTAYWgmVYjTMBL13WibBeO/BYQ/lSfroGpYK
8KSCaxc/frH0uNOfwtLrjVJA1JOqp5namyEFj0xonvMjOLrwuBdq1inW0WC2Oy8/
lvV1ECjoXDePvAFbLK6Y6TodC1QRD+sR8+4XBNGT0d7PJo6i/d7ny+fKKlJUs+iR
SGHCe/8LTsIB0yFwsUwEzEUMQsM21M68LAMwPFCJlAla/XoYoG3guij+LvmyhQbw
EZMip9OqpX3+CDbEtMCbXld+9cuSXQIyU32/PebeJnQPCLtprdgse4aoa6Ed4Lca
CVtIpfRRVai3dILu0jiBRrOFFLzaR6lp7Yjv8ssHZc3GyRqVmZl0qc1GaKn2PQeC
PUOF6KgHc5yRj0qvkhlyNrH4OaXVwK1YC6h1+F3IhSB30zPS81Lp+Tsw5x8etI+N
7t0rkA6qTkVrqZ3hNvpEQjjScDazrLaG1KHVvFFxXX+E9qvZAz2DoUUz8B7a/tyC
gFJKesG4G0QnixFV4ito1zY2SU2Qkrz8UOPsml15jgNHl/7BqH1nQjqL11mUK3IY
jju6yCK67c7WVg1IYnpjuGI5rlSIwS7ePGafcIhQph+KFy/KCK846rIWf65t6pkx
T3lerv1UW+dP6z8Fxgd3V6pF2PS+2pu8z+CePnxXm3dZx2XHaZ3FOoJpm2kISp7b
txdtDasxbzwXxeiK7y4nion/6Nof2MGuM6FvnLbVmW18jOYagD10H2gDAdUgcybR
StPEeBCYm/UP+8T5+vMMOoz0rgpyz0rJxC4x/xOYehIgZs9t47CYwy5DldPQlxsE
4imp7lChyvm0EDEwx9BUVpuHFhTlqfV98ovz16bxP6CoXYuuRxE/QEqfxUtZidqv
Omom/xUYtOWw1RtXBMe76vm/pLaYa2SoQvojsqVR0Kx313cl3IdKXvDAFNwNhQo6
uV70MhwlTLHIhdwel/gb8wtsYKwSu3sj019YYzm5pWnP8yTf/O0sYhef8T8pOkm4
8O86iJMGrJzNI9f6iox18+6IhbXRbCWAfCrY+SLJoG05zzgvmfFG7dlorV3R3hkZ
88yU7nSB1tHnwBZF587z9w42hnrrCffAj4jvQnGPV37/DMb/QE3pILuE1wKUAffC
l3uccnk801V4CY120deiB4O/JS9XmCkfXrVusEIa/fYAazt2YjXeUErcF+9419gR
N3L3GiqlV0CUtoDolHhfMVPdabBPRu7HbgunAofu6mknxvpS2BMOwxis5KeR/01b
7GoaGj4TjUgoPKHY+LcNRAziosw9orkjBbyDdKQ39JIcdihWgM1dfLWoDgrBlINf
s6jG4VTi0RT/YkppLzIZR8nJobWZqR/wyHz947qPitgcWCVTckEXpZDpdEPDugA1
Erh16MbenOzW8sY1nT9UDQR7lGM0uuFhrVRfsKdTBsOFPCPVJLOxMS9EVTXASRZk
8WUtt1ulenpIoX0TwFasQ9USCexb5IRXs/XBcr6ZGuhAxV27JLyBJStDQbRTas/a
amHnTTCr+GW3pPe/qIolobXHbOzuNY5ovSoGP2hjot4D5RBLRoYxR44T1bHrqeka
DxgHIGU/D56naCSwKrAHPhX+F8hDtHgqJAuuBGZRbWgvX+TLxE3cPui857m0MHtm
n/VvjMMtleRyeYl5CEHYPxQmv7r3drbwtzhDasGsn6nvYsxTbTsFg39RGM2yHqXW
B7gRXb7wPfUVP8dWY2mHB+D+70q10GyDKt9qk/xp+Yi5zzF6/T+JE0DXWby9mguq
E3Xsa5+RXlcGTHaa6TL4wWolhQ+zzIH8Zfps3ZonFBIxCuO/j5sILGp3TAkzeR1V
2grSHsi2w4b5koaSeN1OLQ//xq4n1ab/isHQaLAgdJTMpUxBKLOd/aLZYzLtvF+O
aNDH9oedJLQKKnCEL/8Is1a5sQ3zo/stywbBtOiKSqxJoeUMKzk/RsQkL84llm5m
HjeppPLcig8Q3qy1/ZPgHNobyuhR4Pq6KypAnS0HWflhMpe0DBhFjfPBiDWtGMjm
V2mjwtE0FoDBiCOZKeqE2yzXKYRkP0HCUHdUMryW71Nlg56tmzeIYmkapc6tfJBs
pJbLqW672dcvoIxzKCZlkMYwR3DYyv80kSgtmx7vCOOgVUvqShjt/JHdWN0vHpR3
Mh8bhrR8flk2oYgT0fRXD7P6d5OuF8hzxm8/6monEaYjmkD8T4qVE/EvtyaG2U0v
Je7CPhvAp4XE8uFWLk8bZP6HiACotc4BfNmRzE8ej1ouAdEjShTvbpfCtxCJujgo
N69+jv8HNfdqQbiDIjVBMnD39xiBtDIpxskYRierkBodhQI8OiMlf0A3MMC+RSLB
FNRhD9zL85ItdN8/jq4tQ4ZOKZ0i28pSjET/Kbkkj/4bdaBw9uXgV24bH3xZ5FyQ
gDBK4KRTiuG/cz9IwCxWk/3zUZn6o67cWHv6YKerKcAZJRwzWbQO7EpzE+TrByRa
5Teph1u318YO5p8jgFOlrmoodfq29B39/Gfgf188+kMba7FI/qZh+hoXHubWbZLE
HMNaR+RSrCNl9k88pbF0l96UGBsmDKTuiYrHkJRb/QiskuAcdLsPzYGvlZ9qFWFg
lllE9HLSTzAx9YwK4XE6LhM0mAFxKFlwvQ2ixVP7kSCAGi2Ckm7zw+j/ZLbPfJCH
yJX8XZDyGvhH8FOkJ+t8RBT9jEO/+CdfoNT5AWUkmMWdEPj3biJ1owIrLME7pWBl
NWLjnY3QAFYjHYre1E9nWevJlNzurK6AfsOwd2AOIx4DpCdPUI5qN2Qek4FeuAmS
fVr+aBipqbzWbXMVYA4Yome6zXgrgAcMkpx1Ppe3XcmTTX3tgfhQ9WmOU7ap+MzL
rXlMytEXO2mpuZYFW3un4L5N8U1driEvtHc89I3It7Vw1PJd5gwGAcrdcAQsxJJ9
5DnX9nTrz1yRQ6uP5ne7OkVL9vd9aQYh65J0VIVN1M0OuFJympGmYMUsIqtwfBgi
Es9KcCYon/+FvvoRa5eI172sMiCtYidwoi6L7E6aGl+FVkfxrogHYHe3++lUYP5F
uB3d9tkuwg+inaT1xXU1dhTWnkXe6e4LVIsXP0Nc3nl22y56/ZuC+SXqKAu/K8JK
h31WXd/LXVazqboMAx8GUK27k9CdONoR5MTadqyCs3Bt1Y1FRT8Bn3xuPH487DAA
KgmRR+Eaw9YHYEW43oGGLaE4wEb4mhHed+pDDG2SjpZbE8BjLnv3mZZf9ArlCBk+
Zn6Gp/rbsCWhHEQ3B5chZS7s8M6cRgpO4pAIu3SlETDvE6/yPurNhMPMj/8zLC8F
77ZifeBLHTwawk157HNSN9CgOT9JFzxXJ3m1qeHnENDm7UT1DIQ9Zvu76LtAUNFK
7+16WF3JKv+HA4Uy0TPQzLsqRVH+duo+2gRQ44bvP2Kni/jQRD3+Uh/OKJtQPq8J
0AS2CCl6167IgXg+dxw5rPg9w1Q/8j3SUSNN8Nf0EGOQSTm/Ap7KWC974BEVqhiH
DLgWZcQ31ZUwPrWU1LT9b8zrG8QN2r5jZwivf8h2Kfevi2ijUI6l6gE66r8BGbhy
EGvZmJEjZ3i48bT9SXzB9LDNBvIumgmafMtYUWW6gZsgwn7EJc8iq3LRJFu+qEJq
WZrj6pr1w2yThyX/YSNF6c6M5InwSoa2WztIdBpOfCjzFdt3zSAT2UEDjnoKCdEv
SoRkDlzk4y/J7FhQp4dSuaFmGcaQVLzlq059fKTvCELASVU1zqeThQFqkBO7FXdq
zVGtO9FOmDpIWEMJWLT6XbFEj8l1PInoaJjIDdkckpN5Wjxm1zGnhlk1A7rxr0aK
DmU27bna0MOnx7GnWISIvJcCd0Tn4KIj2+gqivcQW4IxnRJVqu6ITjoGQ62IvtZs
ot7rgQ0n5KV+Oav7VccKtcXcqQGExgy+q060uuWV+KSogJU0i7dFfGogtxKb+nlf
edeOpQmZCxbrTQJoDpTQasrm1BR7PbHj+8cYXsYfOwJHXj/cAnaAR+tDb7N0byXq
Ziyj/pz1aYsRxsGYpslO8CW5Kr/hfegTswwhArQVJoMpjhiq+OnxPAApvdrDBpTE
3NddO6WAaCN0gmwwWNmKpNGkXvh5LGHD8W62oees4g8z+/23hvR2v2cah88PJDAP
moZejht8TtMjjj2tG5AbUX/PFHPWIrX7vqhp8kTflGYeYs90c+w03pJeW4D9XbWt
51nOAQ7zudg1okodpTwKb64kGfN0Zt7ReQtZNVsVajnPTPbEiD0slMxGAQbD+J4s
DdFifV0ULnD+FuLeErI53JBxRwR4ONMurPnjfivuKgeXw5btgx7HXJ8wf1ZY0hf0
V+kZKvgW0RZmIG2HFajfXysPV6g7XL2RGYz9rf84yNRSJZOSZL3+PmnY+1O6n87h
CqNtEs1t50WLUhtOpvdU40kQN2AGPa8u8MynmPDR3Z9mEQq9RQwd/hSI6+IdUn0U
oMkvsNpXbjfa8HUuFn+mRYQ7I7AYeV312er13ZI3oJHaiwgqgrkuG86TVkZeZxZ4
E9QrzNexC3j6LSy5gxIVlwcCE0kLi/GDTpG1mF9TjyU/XSgmmlhiUHA82quf2g5K
Bt/zwjH+PclcLFQTXqYGgY0xZpuN/6htpy3lcvPoVeV2/MlwHDq2hhTPsKEiljVj
P7mctTMqBEkn/X0+KU5w7vbv46087qBp7NNjD29GfA1RcrWi+7D01ahZsVfHzyof
iEtyDb/9Elj/xniOnrZNUq7abTY3szezgVqScEyNXQRSwhfHV0aSaYhFi8w/Rbbu
eu7luf9/xhpW/alhoerddveAzfPbbSsRM70YvGgEKYaHPs/wquwz1PMB98I1gs+2
f9UkkbWFqpzubE6lpSS3iB2J9A2y5pAklUWGSpcLqtOInqn9q78nZo0ZaXPRt4dD
XlZzSiTBsFhmh16ejGT59taW6g6Zlz04+SXIVMjFQ0UjuYR81yRL0YvdWq0r5kTC
Vl1PCsfRVutmWCdPsVTr1VOU739Nzx6Asr49vYknmWw8+/U4F95cy4fAtdFhn7uw
5CBDWhp1CKxqv4LiUVThQE/tWhjvZwdhAm6IIiXNp+DijV119vzyyZJHkomI75PW
bVNHvUluPb/G6kgwgJPvx5fhbVoxJbyKqrGS37Bbr8B4BzPUwbhE50PEKcWDFp8P
DYN82RPyMrQqsN2zv9WC5HqIoeS7/9PWR1pFOwM0vmELN/O5BRxJLzcy8jcAiPn9
jqoyjAM8EBRZqkYZUooTBvbLHx0qi4mmY4I4IufGkBFH/wcaXYlbHZvYeq38rM6A
J5Zmblwkm3PK+yvvnioZHIWJljxp+yda5MrbLE5t7Me3753eDV+hJ9z5ViWyGoTQ
ja2Vxf2BDH6rV6CoWIhiIFao5YmHRXM+JkHUAPBfHzBWG//vDskoDWcOf+w0bzGk
pJ1nIglwQaxtS17hJjdoyjX0cFW96de4jGu2yjLq0MCXNzQ7e1qvuhGREj1unDjG
Q3cY8j089goXC9OU9zPkwzV513TchdtqRRVYwAvaeqKoAos5c1K/DGoS8zZLDzPP
Q2KSQIIua6O5PYaY96/h+wnHjwQrAKL3Qb/NlUP9Z22kG8zECt8P9yY11OLqESRb
DLuYZyWYF3UofD636QdlPc2uDmy/AIJX5me54Ex4P46e7W0+lRNRo6kc36O+0Vxz
P8MERaAkW/woDJn6Fo+yVpOP37rdyXNdww4qY6H0tVAsWfJwg1pQe/kctorULCbt
JXXKt4Jr6Q+4QQxx1H/gpP2FxOzV9i/pKj4RUOrvl4Y/Pk/y/IloxX97AqpYJHvc
afUFUss8zgjuqzaVG9zkNGQqRzL6jmod57dUuegidjq6gHswYsWpiqjuOmjfmnMV
Ww9V9F7NRTQ0iIzBEtaY6t4eKf1RDW0928K8+HwRYs2P6htIFzTGK/wZ602Eg9rd
1TK+PaNY4UvBvI3nGYS7zx34+MNBKp0oYoetxb0Kq5jA5BhVVxBMZpw9rIgt8QDB
4d8ycHSZ2byP5BTWyCXFBSki/uPBFgjjJcGUJ8kzsWxwSUmReLpBOePyM98g9V8K
9Q0FVZEBu1l/RQMPinGUaOw2Op4/Ex4FScNM86BdS9Hnv7S2sn7oFHdwty1vKLyP
KnIkSINlpY7S63WlfpgOmxCs7vop2+ElUDlt6TmM2a24rEkFk1lTXpA6JUSjvmsc
6JFAoUojdlXcKLc64VZEdBvcJrzExf2JGLamercT/SL8uGWZ6n5Yz898JqVwd+7B
ft+qH0eUGm/2DaWtl9mBqI+3+pQwY/hNVLcV8gNn0X+i68WBhJCj3zHJMrdeiguD
7NSCYM1LrZFuNdJXMG+B1Hzu/EWh28heQwwh4cxzA8gq2PFVlmt7Fwufagvd3juh
djvael18NGLWMmp1fQawAcKnDsnjEimGHUgZUMsn8o9sFeZ1Trgv2u5lVNINF0X+
zD9mNjqP2u4Z3phHhYxBXhkxOIfscgJgWzCrTselhB3tsWOOzzsWYsyShhrrCBLB
YEjzXI51QzPwWvi6uw7HossZKVhe9B9MclVTRzGhckhI4Q22PDzJ4Eul6ynNisRa
KPOhw95/nkcbN8yN/j0NlJz6+q+8v9oqps61xsuslZ7k/Ve0yJDUTMd2qmL3fVvO
d0xOa9o41Q5Vcd0Nxvvsm1fK85sDaSvAtl7N21hK7YM8z6Bq3Wrp9Vv8q7yFYxXM
Qvwu5j/TCjl9Ij8NPp33MgS9OuCkCPGmbYxud7Qhl5JwXOhcixk1CHx1KBNy2HF2
/j76KOr8MEouM4EKu7bp/rmQ8peEC5cbG08r59Mb8Uyaj0MbJT3Yw3UKaHmvtAzL
a7vR1IO81PZADjO7jvpl3BrT27dJG0OsJ64lSYe62NxqP4Hdikv5otTGyLy/D6FC
f6BjKGzVNv4s+qkNjEhiDpKcWmD2JvKirqMjeogSdr05ZNHpPiQ9kMEbgcecdCbU
+0WX1Nu5JytX1FAireckleaAPde9aUVet0uDCG1UokNwXi1bfIw/L6FM1CHd9iAY
dvdwzrzqny4vIrq/X0SeMWgRD4Jdort0+mxOJMBGXvulbAaNj4uEsrddb9T78yk6
cIXyOtxzPrTppiwYdm9Li5HrA3MJyiMWQYbxdzbVlhZdQ74Gmzq5uh/skhI5DPJI
lmlSGUiY22TRgyg8hvuF1WEWjf1jYKwp3BrE0Z2invPBUSUh7VGnZalQVU6Ek3XY
6rVSkIFGDfNFIDDuPoF65pwRr3QHD0gSuRpTPloYWnExEABJqLLzHPnFCEfxh04M
vxORzhWJN0TJVUAcqtWv1y8xGjeicOxvwOZQoLDF6/6Hw7I4a0B1Mt0494120K2D
cOpdjFWVczvgmw0DQDBpMlJwUzcTa5F3uMy8/diVWRXMhItQTFurEMqD1PTpPn7K
IYy4PfkQFoX1cVx+PoBVNlgYayYpV+wXGQyY3nDxFv9zW4Xp/aofqSLmZSOt2LKo
3fobrwyUS6VvfUWRPTxCj6ZWo0xIKg9M/9l0gpyhNmIue2EMDJU+AMwMXBhGxhGu
irOE//lqlhn3h3hi693TsDynvUuo96XPLxdJqMFPHFBdYlJtdpAld+WHrKiWFNKD
5ykaMyZ28EO1zWk2r5pe5UZwQRmIThSgL3wxnIfqxK1bnqq7+Qa60uU6CkZYLSqR
ieRZKzUae9fjs84nfgL5gQVYXZd7kBlbqPX7YUCeTOj45dGsVcnUvBEiYStV45tW
U7qfWjzFo/JsUVkqa8XdQZRUYw8wscJPSRJvgtkiHSWdupHRo5qXqMRGp2e9buWH
TwF8rlNwDUg5lbWEHoJgXanhfkAxByAZfiBsI2HbovbM05es8nZmRuKACgPfGx6g
COnu/hCF8vnlFNm4W/MflXgCx4tVzh3Glx2qljENOOYiMNB/vpwveV/nD53sFZJ0
w4cz3A7tq9ZvBiUTV+3CRgnH4m/unt2HxJznBGwJQmDDYxJxoepVCzXKMdVz/Tig
gTr3udNaMJ/K9CZj6EBGuCUo1NrJssJap8SkEdhr2v1uGzmP4gHFRaoF7UyBVJm1
1dcabd3kdK8NmojObCGBfcyOaMNaohHE820DN9gXfXzkztGDEqlMpUxw4zNM3v2z
sCilcMBX0kbzxJqY3ybKJQFMuuO/elLWGOypBpoOWLWXojTrZ367DHFw2hSIw8R+
OSNXKB1Z5qNdKexbwjhR3LNPbCjsvZQmaZMj0TzrvOO8EbpAo1xkPPNI2ARd3lF6
jjbigpS/KnM+AehAExZ+DLdaqH4qtCGZrbkeLn5Bw+hmmDJRycpjNFbEq0BEhG25
a+0eIBgYonU0m3yzVjWmL3vkFrupXfLRpdEV265LwmKw8ccX02brfcTWGMMomQzC
CS39uLA6AxQ/oCXPiI31p8lsLJT7DMmS4qKjPxkvO3S4kXAYescISD9hDGT1x3eE
VG1yP2HQi9opVku5m3P10JYKf/95AendhKOPuk4/T8az+76+sXxS3FmLiyzF7xfL
KaJV2aOQ6NNGM9BPp03njGH0HVr2OKgxLQvMhGsrzN0AU9PpmqAm7eSTdvsI7qmQ
NT+hkQKAdRX38tJN4ecaVIGhe7yk+i7I2MHYPdM5EV6Q+D6TI9zY3wXMEj4qVILA
8QFD92mo5rltJJjZKlIlmlSCZTGA+DHhp0QthgMmuEaLa/wt64O4Rz520Tilgl6/
xtSlrbO0LTaHXJCqW0NBvi67a0AWti1xYwpq1qZj4K7/YqWp1mbLX3aXPY8oJPAL
m8NcyF/zTsIXH3WteMks//vks9/XgVtPfdwPUEEvtT9YynWg9DLNJxr4FQuUAXqN
MJZ4LpYGtMOZ/8+tcD4NFBlbqJtLKl3Hkn5vJy6o0zFd0qMnWvclseXLEXOQtaEZ
Tg0g/Tn7lksMN7WW9f3G39zLHv0Sz8cZclDCV+Erz+OJBf8YJPQoT8FZWbfaoiyz
2f6zSgrrGzON1DGk4Fka7tJOiAg8i4H1a2sXb0DjjSvUqeaCoMzX0K8plY1WyDol
mx6O+DxQrggcm/J/SIXDw3NbbbogSh4DHtWwjrilQMH8VbNbR06EU9hmq9CibbqP
OSmGDlRbg8ti6bd05ZXv1nABCU3xVoDd+izFCYFaDzxpddt3JZ/vMYcp+EVmJbYF
vxQA2Z5Yu9FpLUVoid5RdFX3rlTpTqoyubPdyFVLmkVcqLqmojGPvQOoBoE6HPeN
Kx3t2S8Nwsr8obeDLP+FDrt+B1HzK+lMqaF5qEi9roUzgE4yeBUZB2uMOq3ewrJb
rGqNGOj2Tr8o7mcXJFb+QCgjgILgNvzRDb3qJpDJ+hbFHxhrDruNLrcOfMBp/4ES
dP0OlNYz2WE03thsdbYB4Ewzii5wHKUx9IYiHXSU1ameXAF+3TIXMiJSEuOQHswD
6YN4Cpkmx4YSu0u0u6IylwBfnfHVROLU9e613Pub6B3S3KQMIrels69UKTAPYemC
cwkcc2FF2Rh/fPkCMTXsHA/wAZBzOTgY4JnThnUOifSVDiB/HFh+OoSfjSxG38an
Ui+Gyr0cNdUvxPxOnfCLBgUX/+x97TR3jceaX+LPOaPCxyo2k0k914fCzTdNWKCQ
bMGK00FKhC5N0Yd4ZIh+eEDs/B/KhN96ySuS76pq1MOBNSiMValXOrLS/ZlTj/gm
fI4YHEOwS1l1BVmR66c6JaNORL0/sz03UJ9oB09y/uWjQ7VSWQ+KPiCz8zq/SZr+
QzhQ5YcVZwUTBduv4mmrHuQh/hC3kofh+wnY0u41Xll2v8DC7r4rGvrstT3aUYqP
m7mBtUZgMF9K+jgZ/2qn1kyeBYrAg5fYQXt8BCudiGXxyuPYc2OtkJ9zmCxHhaSS
n66nnqPpxi60YT+guvZxztetEQImXr/NAKlXTTFZxUmbLec098oZz7H8Vya7DKi1
PZ/3sF6zLDxYqCTKKSiQVczebkmJvGvX3uEHVw0md/oc4bIhnXbG80TbAPhy0rIJ
spBKU2+LjYp3y0aRu2ZlPKMF/fLpnCEFaQFeyYhWCz+lChudCycYmnYX/9FUkLqF
FAlwyl+pV9f324CbjY8A6Dezsr6FIQyK9eGLoJynTxH2srBUFCLy14zcWlIalnF0
h4/dKYeoix3EFY+G/zBselxPvLOyf/wjgfkICuCxN45lAjHU76ZUJZJIpIsBEywR
5fXvW7juCY2qMHA1J3A0kK477Su7uv+gsaH7BRGH/3loAbidM/oJAOAoTbijUTZ2
5q+HYpbjOu0MfFkP7l5LudUTH4SoBNJ9tDZIQz1RGvdmTJIICYVfv6CWXpRH6rek
sPexM3mxTu0rsCi06Vo5wLrYQSL60+syED1VWDhEv2x9U0nSOfTL7w4/Tm3j8h9N
NaLii6VuZgkFS9/4nxCG5yl70qhe10J5IhLiZJW5fbPgBSnEroxfUO8VOLKRoEWc
egn1nJ+sXb/sr+J2UseImcYH9563ymf1R9VuzyIwUDK4RfktnitMz52Brk+UkBlB
+o2UTABYTUvG7q38ENskELILGnsv9K07kQrqHJs1RfN4xwYf43cVvERmYX91m01T
LwcdzfWAM+Eh0+4eKNpqjL6fSS3WJFM15t16bylacrfEF55njg9rJlRuysTqiv7o
HzRlDCSyHbEeinbBH9dpqVmb0lU/GrUJ/hWBLfxYHrbeVePxCKYfHNQfpVXy9NsN
5PXTXnaEkjIZ29qkGQl52sq9rrEJ/Wlc3DDd934fVMsvqBWhvF5jdVSDCWlC0yZ4
3r2s9gGrqenyBzFwzyWgQgAfM7uasku6BK+blAJJQ/sujylXWctZyz7YmO8okJ1j
3fWfg2vMyQK2xUdw+pCxAwtbwWJ5jUwtWUnWq33k7ImKCB0r3iMnovrrCPnK7Bj2
APEANwd1xBxFNk5uVDOUl6I2PKEOc8opJFu3xjQ1Ocw6dFi4qxNqRr+yIGQ/MRDC
DkF3ncspC6soh/4NGf+9uo89tPk77OPg2rrdGNbq5eUQhBNTHZkLV0XajeiLWDfd
AOLOCDBdOhrB9FdFS5bmezKzCxIuc77KthUWahifgtMQIVHCCa3gTNKvoaesgPrW
tIsQh7AUBgk5GidDqkuAXspUliZ8Qkz7Fs2+I2i3lhYCO5IpTkuILQ0YlrshBRKz
+JtDsoZ2Sz4BdJkL7wZh0bmOZQmm7/WxeDGWAo6fICZUYKm0Fga8l4l24/SHFyq4
iy6w5fYOUvvTyguX1gwxBegMjBnieHoSjypgxL/dopeKuBSgCcFK3d2z1rRfnLeh
iFyECPEDyuTPRsOKDBZYvvmmu3uHyJvOkov4hTSJmsf66utqcEXWisvV4FvAApXz
0wy+otkKmKQAON3y2jFz6v5lOsIOEDmhKHoXNZV+OLWKj0RxKoNwy7ez/3oEL5Rl
TMF10vEVBZ/fKI6HEKIy7tgVM5l5jyzBqFJFhRaz65lLXhvuvlhbG7nk3Laf2bm/
TDrUxECD5aUrjxwZ6lSaWQBXJX/s84nebIkjExXMosZkkUxyA2Z3NPB2z3ypvYlD
RSUxR2qNRy4TV+wA3MrLdSGBAO+AWa3Xa8wU9Icolciq77YNGLUcjT3wkqYsDt2h
YIJCrW5pxTaSO/7BRj5lKh1yKbn55tnK44NSkcbVHbNQif948tGTRfdDO8+0oIVs
myu67ORBRQiSzg8VQv7TWCqd06nDxkMD4WwmPw0qy94IaKsv1IbLy6DPnRhTcqNR
mZk3l3MRlxns0HmlAOaL7FDmnQ1MfhdRBbHLcpm2P6tvktuFhdjwGHRiw+e0m1HT
6pcicWtmnCfI51iRoGrdS0KswTsvAtptQVYGOu3cbxKDskSoawsysoY9FHcWeUoU
X5Tkd3VBgHEOY2J+ywBK3c4azr7PKfnTA5IInwWqNLfFTRCSLKqTXOcNNEL7yqAS
Bss0p/iEYKDJNKlyyFWHkqEZ1mrnVg9lNFoF0Stv5Un0wf8VSjKFy8cxEL03/eic
T2cQoPAEl+OugxWDMRpOaImJiD4SS/1OrbUozKW/ZYfCqqXCkaJHG7mMUwqLjpi3
c0JHfIp15kdAuklSCTkWPWBI2iDSR5sMgzLMKOe8bbmfYwLfUuWTXEQXt/PSwnhP
1m7ppRY0FBxHMadY7TpH+xXvMz70pOnldFs8Ejwml/n43jT0z9gCchW1vvuNBRpo
aaMmVxLjs1xpoZxJ6ycJpB7/gybHMwHINGClov9vvj4VCBvgjQ0djmyeY4hs5bkA
FrS9q1Cg/mLOAdHMe/6Q+elnkjMuf1nLQMYhSde667wK127lCdhXCUbvYJ+KeT+e
kwnRaqjSjqwQEyaUz5CFS0LIwBxfRwSVyGiW//6UVy0IRZDTYnYdGwmkDESRzG4r
3hOcQAjTkk3gxXyepU7v8fhlmdnrdVvQS1JRVLc4gQdNqVPnnrxhPEf4C3+vk3eZ
mg548xjY3klUns2m8Y0aIgGZ8TWOSwrMTsDDlJr4I6xjxEYkG9w42gGvrdepwoPD
Nu6Ys7GbM5qjpZjXSQipoRxUHngO/FZPA1Y4Vq4jjVC91gY9bOHgJ1QoupFz+OCI
v0BY9934qxsJ6QzKJSOrOiacF1WuDMs4mHyECZZOyFyutLLk5x/HZ1+vHncSZIRZ
Cw8maVfncPwNxfY5MzVfBv8IrXnfNvfszKmULDWrt+M11LP3ftNp/5iezgRkAHmm
8SxRPVbzdHMdet0tkY/K/DUoyDwOuwWSjkaka8pZ82iSA/oYMJu1kGfqe+1Cs2Vy
7OjFk7jOtpVF+T7TzZpv4WFufey/BPlXpG2+lWaRBeQtYK/IDCvl0RD36/o0E4Rf
8NAk6dyYJQRKG6VMBClok2fVQ/fNdMOA5SeKng8YCQt8UvGE+pDE9bqLde6lFiTw
XsIOZ+hDiFnMJV+JIYpR/KSZLteTTB8wOa6QOX2bIKtZJvWAzrj6WkhjTkOaMzTM
Myd/Ppav4piay1O9ml0V3WCIf8GNrcGwRW8EqM2GDv7qzoIflsX024NOc7YX7DRN
0u+V47t9VewV/eNUz+O/S6duJ+I+fY5UktiVqvJIAIjhhrpKAtOKHUV2eRCG7sH7
cfA46KSYYasNjIHbZHXVRSeFlzrPXZ2SJWlGq9fNyYL7c+YG3kWBeAsaKnojQIrG
E/GzlMLamhgpaI01ltSFvMK7oVFZkfq5nJw4lAFDi54gQ0YUlx8bse8e3B/0U5KD
r3J4fZ1GlNMpN8bTJYo5zMx4eQbKrX3JNsEJKRQ0Fx1gUFX18YEPfozL4LqfUhxe
hieU3YBlAnkH6glQnhRgAqmxlhoD5HbMF8SO/0W8Q1+QFrwd53zBEMEyQuMd7tKK
urcC03jSsUcGrXu9CVCZ8uPKRt2aNTz98/GlUa02Ws5GJvPKSTgreIxJJFKFGAct
e+UxlLC/zcoqZ/775S49JLvQk/Xu3gUeKVfnK88A3ohhpygcls4+AF4WDB5DbrXi
VWt4GZdTk0suDEZYWcgMIHnLkAN4J7Ffyocrhv+dIHxxCpGw4o31kLsKmvMNH+Dg
Jx8X7OjU0J79+fA7auL2Hwn5s3kKz/H0IDL5x8AgkKDR5cWaKo0P8nVi0VIuloez
kbHJ8BnAUA/xWyYR91uzainaU1TtdFPos3EFVuvzUp/Xc51oB61Ma40W1aJTfSCg
PBL7mplykE8Okkjd5YzKRUYmFB/hsrOzu/ZqSDJdNiIrEShvBh5B88yySiQQruVG
0gh7g4bNbUvB+iR51+qMpAwOnk/kYZV3kh+dEYSgc7LINgSrcocjjUCuEG2iRzGh
uENb2AaZzw2szy9+YuL2/k9UWuPc7vgKkckrcwhlIIJJbV53ml/5iLPVcW6nfwEI
GeaCtbifZN1TVGL/+BfA0+2SL4RKo+vY/NWinlftPW/JQIIp3pZNyk8fzql5Qiuj
egu+hdVf25Q2zyTghevn80If9gGmKvN0QW+qwOsM30FPoQ6Jcj+MKEHOkDzJg85e
HDPrMfo7joGiyUJLYZ47Eboy/OmWquCVMxbTuohfS/d8FNiEyMhiVDcTl8lAuVAx
sERQrmJVQYMCbiGhfatgG6bkX+hfv9U7qSgzE3xepUhLAC9lyfyhFIBbvA1g52Zp
EIaUSomMqI0GRPhyeqLPbslJ3xnxN11USMkKotWY3XkcVmQjMcC5rO7OpMP7yV9C
6uANVEGyxKU9gUCzTQQGfA5C8hIfaVuueo09Bbz4wASGT50SLNcYTZ1VdH2n5fFW
V1gMasfw4Pxfgy0ONoy6dc1YzLuhnX1Xh+F2BwRpIFDX6lTNFPCGhrsVip7a9Dik
Yuf3thx3c9Se+mLVKI5Q859VhJW1QHLYDvVEoOc2DRIVae0vw1RXV6pHWnL5Y7NF
Az66fL2AKVQOWq7Ua+JyMZeLK97nlt6serJUHvIlnr6/EzJkOs4vGzAvPs5mphAl
xybc9TMxeZBzTlyazM5QHLwVYU3D3l42cZkcSs0p6rzj4TaBPcebZzV3Cn+dlzvv
JR0VIKBUOzRh+srKOfUsxM1zbie/h82/MNhVmjne3BVBENPpYJ6+6gsW86iRyBKR
el9Nly6kAW2gQUU0kicO1us/dd6kNLhO2+3xQDDNK0HqAZRGCT2dRzI9JdeOvch9
vfpdzoBp/sMQASrxC3GQhnBMAr7tdAr+n1HEV6AjkvCp1t67BpFZPq2fBha3NJKK
zGZmu+z/PXxh/IbLvg4zBGRFr5o2XkzPfknyE6BYxXm/W1ETmasfuya0fRxN9eo5
AWpQe1R0jWiu0/jZZ+swMeZfBk7jN0silSM5v+9gHEeuKt93Yi8PBO/cgPE+GG27
kvTCNTuITozIyeLrahLaMSsaaGvdf7YN5Ild4fnei3Un46PWZ0ZTYwvKOBFBZcPD
XS3PMGc3y3Vqbc6LU7nlNE61LdQBsj6fTLb1lCvChiwRH2yx8verUsFtkElgUFra
mbajsIF1zO9Qown5quR7DT01i6pTG9XGkMHwH/7M3uooRYH918zenikgzKO3zymC
MqOwCWVSMg5rl2EGmZ3grdTf9loQB7VjNB2H0fywqU7be1lzYbqZEHE+6ZgUrjs9
9KyAG6lSlukyhH85vJJuhBtXW5gVaKZ8YUEGLY6uf1+ObgEEDE05In62s8VBmlej
kBP7PP6fb3F/oX/sO6j/K1PPuWupgdYHfJ8+TB3388uIvC3eBEik8NKf4pfcR7B6
0Bzp5p4jMreXcHrgmq3TD8VGmXmTKq5OxhwUsbUVo+v9gwckdGffxXcHvpwHbWZ1
+DiIJ2AbNA1fD3+B4M1C+ZJBBpZgoWjWL6PA0LGpVhUr2aydxxXvlhucYXd8onB0
pIGvITcTT+ldcDVB3VTDfOGkzleN7j6/n50B67U+fOEYSsBaCGIDS9KUFPbSW/rq
44NwWKTdvmntnXXqJpap3igosRBxlUGdMGrYrY2xADqgh9HtHWNDzZHSbM9TDr6W
+A6W+Gi+qTakj3AAWSXjpKmVnQf7VNabnKK9OOM4oz0BusfufEoxT7BlVzgW47Kk
fRdbY/Ri0VJGzq12pB5NpR/h9w7kdGQMdTVFkLsXy8Y3V7zPrSQGiMWmoJFxfne2
Ygpm5YUDUDGhbaVpJj35obzDoF9rzgrws6vyT/3AwmaSSFPrG+Hqv67ck6pqkuqJ
TU2mnPRw5TJuu8U2bDGkPD9qOxSOSusUrFV7yusNTdfzKfzqG5l0zSudh90xXp/s
IqvOgASdYB6oYpmvUNqpfDn+Eu6c++uM3R8YYAieIU7ch/vSiY0P4/7Fu6JMc/RW
oopkBzpN3DFJPvFHsKKg9FYGmxxeAIi7e2n6hf+Xri+cNN+9yclLZDT46U/kQfw7
6sDNcDIcCSBwGf4JOQnOZ25d1tZuTsfleHHaxPT94gA+0rPH3lHTxAzu3yPhcXjn
NwE5waxBsPkObza+xnEqf7KosINtGoC1vpU4JdBLB0KLBpoyT05bD5x+SmWi7CCK
DsNGTg/wcGzFjD3JrYFv4ApyjvFOWE4wPS966ubRSu5tJrZFIvLY1jhbm7Lnpl7U
UnALv0y35x1fgfiOk+x7QUUrlyCaXz9jsDsNdc6ChTYjsQRm9w7Aup5egqq+ZrOC
mtpDwN8EPolxz/6tFpE5ToBVGEmYjRtMIfNXFfJFnpk8M+NWjRDfCiX/x1DDNbyz
nlNHw6PYzyPgy0fcO17y7xSDr3Oco1iGYjg3K9i7jXzMeCJZ+HdlnAFE3EtDLocL
DmcedvZ8FmDTYj/kaOHE3DtLXFUAvBaqOO2y2AdYekBK1w0ZBlxHLekZZ1973TjW
gzYwXVB9c2iYk3pXvkqrtHBGg2S+p3p2QgaToPQ7czxFtmPOXC1Em63ZcRXTLM6N
FonSW+NSzFtSUZFzqBcjHmxc763d5qhSvoDnFWDTNVsoiWHCIANYpkviVVIM26Pq
YVLeTM0kieBWOiH9Z6VsyE45Uw86uPaE7NN+ZZADCAx3HQ/scFbuiGS1u8tK3UbH
XK8acGUEInw1/Y/G7aXJCAg8XIO/1D13kSa/APQoPdSVM0AjWSiQRjMagFKtXEUA
oJnw6BYyBHqzQ7XWA6SDidOu08cGO3AwxjdAFJfb3rTCVSZmjdqVE1JC0mcVc9lO
YZTwLxBxcokgVCatiLRwuUbR3Z7qTR2ZiUVsapbuYuJu9EL9Gj+brJbZ7l2lZ0q1
e1kHfFDlXUhMM8GM9bQtVSm2nyn7Ef8F8P7R1GyiQ3xFCtLk8CgPzNVKW0BBsfJm
4XFOfV3eiBzszMjELACUzRDo5HhnkHHYIFlSaC0sK2BjuiRXAZx7Ax6SSR80cVdQ
iL5pUq6M3bfzBGAX8NYEXUZVU7KMd0LEs4pfqyrW0aGCglCtTEMdMpH+xJey7oGc
4WG7qi8aiSMRjmV37A0rwuGjgHxKmW1pHLUsukqq/oH5c4+6AgOGkLKJ59yuxbvK
rdv1c0bFf1yRjqB3pY3XfSXd82ZMdVsgRosuhJbYC+m3gxEviJRsyBYWmpfw3rvI
zTghC8o4RHlxi5ndIAuY0f32gRhaSOfvTtXVWRSANk51WbvLqdv68oPXo5Z1jkvc
VVmUHWT3SfuKvDncpHxt5MYuZr7RJmyLZJlbhipXHaTR+STDTVTPFnS7fcVAqjQP
zTAD3/Z5ht7FxSy+3CRSQp9yRZ+PajURb2Nhf58pR5b7P3Ic82VZxoKnndw+kxlE
thP0b5ir0i4Rmrag/uz38jopWlEzD6O1/W5objrdAaeWVj5eSYY7oEpZFzMUZ9y/
ybouSHGgBwB2DBFNTocDv/Zv+0KDZ7LQxTJ7TwnP4gLgHUWZSwxWWkczXNpjD1dO
Yc6v3aEXyJmCU03YuFr/J2C9zwivUs18blITzsG5CZyNEZOvfN4aS7WGnMMYiETz
9UGoA3KIBJgARGXLxiq7MLzep2K2MraltRGqyNbBhysn95ghOUzm2RNACuA4J8Dh
zk7lxCFyden4Ecqz6XL5rxlXcy2Tjwa33pnmt7iX8zr2Z1/6/mtS63FiiQPC8JzL
WYtMrXp6QJ+yawINF5XPDIK3a+K3pD2aKXjmXsBmL61IOc/nr6D2MoyeBwn0mxSg
Uks8U0bI6G91SaeLvfe7DE60A58w6R8R6XiM/aWuvx532DtQbTVaRG+BIsSMKsK/
OZ+32I3k2CgMKCGy3gg98CXW+nmG7//0IuDG9rtKrYCI+7cpJ8j7qIMwFky4O/YW
u443zNTMMBG0qDF2wsxOBbaanJaIyYSXPkYPzRWOd2surDHkNMRJLDnw9+0FpHtn
NCNCcJYvxMcyJEVvmlG7Mqfs5FsqVay42hKlRAwNpw6adWbdn3yTzO38xVsSPSJL
1muaBIKh0L5zc06RWVjPmPOOkZLM0Rjnx1Rjiw6gaAAr8miGBQszXoMGiaBW/Iy5
9vjmcYMjsD5kfi/OInFE9gjlIgu8wWb1JbyMwe992YzxrB/CUFNnEy6OA7Pm6tF8
9TTUwnvh0X/U4+EJYZprHdEviVpeINSdqMs7MSol/2lqKjrmfQE3toa2xqhQgb8T
O9CP0c+wSo3HMWzfNdxZzyOHvDqHKtu6geKGnam7g3SEiTUi9NgmwEnzGBcKhG1g
PleAaK1Bbx0uMr+1sX7y8qjdPlbDzw2F1eMc+3w8P68WKUQcERiffyIi6mo5GXEN
bFOKDMDhkwGMHF8DUA+zre/QYc+LFuTOVMyzj5n3cnSQsBadxC1f7s1kYdQsjO9C
Uq6c7Pt5iaHB0spt23sWB+M6JmSzKaPSn5dXqBE/TN0mhV1tlEciFKhOqEk+oezi
o/ICYS+TWVO81NbVZ3pMApr+cEWICWw/ST0oLu7bWhirbbePr+iKtKe60pTwTNsU
bf8mCktlC8VXfzRFA+y0AdHxdc5ZI5EuJxCR6vIdYM1N0cPPE4ItEoH6Sb8/Vabz
szAmfqxDj07oWvCrj1Mr0BaRfLj8DrTcWY5i0slhZ1jSfeE/hsono3sPVbjr4K3q
te3kZC3A5MNc4+BvNI4KcEU/xUK4RRzhh5TQ5bDEyNskPgdQVMNKYITciCY9/s7W
KJ56390B2KWPcu3W9D2hFbeOqRZuPnsRIkpxdEq1bHj6a2F+cQVSIO8JAhkzxmVU
scMmphq7LvQ9vBfQJBdW/+NLfCzJoCNnrUGfSnl5u6WDn9vC6WHOshmZvFlKPcel
vFKH0GNd5rKX/nhmQ4pk/ODR1fvM5DWkQ2bSns6s4TcgaynN/JTnnTg0FbR1XmJV
29DlCNmXJv75+flZ6Ov35OCfTBg8tyLNDASou9TsLIkc4WcOR8ekWDn3LQv+LaQM
OCjxyIAVtz4WLdVyovFfdyNPcb7pPplyWdpV8k8//t9IiJl9dYMXKYQIiXZvOc+P
TbfoDq74pCDm/OKrH9maYbVnYy6vCsp2d4p1NGAOjCRUagxRGBZqhQl7Q9EYUBa8
syV1U2ujVvXXUq8NuTGwGbxqhD3oV0Q8Ilwhc1sIJjOEoFfxb62Sv9kkTkAA8fUZ
joEMeFf14/LjSCMySdGFN81yW8Qy4ZllNPWr+6Pq175vOsMW7/cNmLeaV78oXa9V
U9LjJPlvKUM1zMuMr8HqRSEppLhHpPe6IYgqcKVjDrR76V5fKrJdUnMjxy1vjnrd
eETFCrG4eU7mHpeQ9HVP3T3+oUa3F6NVolriCYge+Re2BMWNB5PrQ4Malefqy3Tj
lCZ1b+hqQnB2SLI0YVzSkFj5sERWelJog+QeGh9wWVgUbIZh09BCmQmZ/4xD16gd
s40zfpNQA50Ppn78L7BvUDy1KOdRqrPRGbdzII/LVAXjMm7/37RS5nS5xfL5oiKz
XXJTN1mwfrHNBC3FXRKBlDxUaKw6LU8kJn/qKIJyC8qzTj0TizWiezG6Hp7i/N6c
lauJOgYTPasRlschhorf5lWl+UhAyKxj0MHHrfZh00uaZRl69YM/llO6ZARsLBw3
vOhqnUPA7Wb7KOuSD1AYQqvKiKKkebBAZfw4TGmNGUKYIQVv8jf1xkeMZ6w6nZ+X
pg7bBlriAOk7Mfp+QUYjM1WLYsLoXy4VBO+jc2mA5aGvS3/TlV/dGAPE/l6DmxJR
oKbyGPc3KZ4kty96JqPj2LaNy0rrT8sDEDwWmtL1WJmMjQx0cfkJ1cwDAAOAFSNl
OWaXlfS0QVi3FMs9TdgxCTkXlbaw3MgxKUH3OYdsudJ99sW7uHTX2WYOQXIYqvgq
eyZfsyPoVzO163A0IU8hCdwXFgxq6Uokn5jzVCU0EnVZsRb+Vzo4QUWDzn+bZmr+
79wFzXtjDmr7KrIKotVLO07k7dyiZVgLEMIOj3wTDByb+HEmIPPY1Nnm920AzNpn
LGCUmeTyrdmObhS4JXrdXjl3XM/Gd2x/12qlphJzRcWNFpHIykRBlExKGO/4iRcn
QkSsLy0EkYD5gcXeOHrrM+9iC2QKgQpfbUT6kAUvHX984//7yDrFcSN9Wds6t6sO
cu4Qig3DH3ezUDNWOfFrW+n5decgvOGGqHpI3Pb8a0a/aWSnuIQrvcbYopZuoRmI
vkcOQ7MAXJyaYMLXUTboUUdJWWjUQAtrlkSnT+HpwmtW4QfPGTp+SS+Qk3xqy/cC
mrmz6CMdS2+yWtpN+/NZpcHEO8WKuHlJuVCE6s6l+Lg+fIZb4lAVP8EdTqtToeNR
ppG/mSP9ejmmqCFKADjOmNI+sDn9QWNnY0bcGBN2a2igijQVBysoV45gdokMoeFR
AlaibF8BRsKQ7ZG5LJncFZM8OZQW6PqGZdSldjyioxLJRsuGdp1+D4hbQVqnOrXT
hmuCYayD2GJXCK1Z53oL/GGPJ7oj8Rd0Czsy7+gZmz0RU73fY/JRf0O/83xBSmhu
rZynRTALSMGwsD947R9SSnPsS8FMRbCrwVqMrrTxPZNsXT1MpjNWA7kdZtfyENa3
hXCleVBn48BfS/CbAcPJ+AtcmRAfouDCqKi+aQXv0UchoKpNbw2QhfzlOW15Z/Oe
0es8Gi6xdTztivtu2v1728syz+8DTQkO0FAmfCu7ldBJ0RUVg+WJuYAb4PSn5xJZ
S+s2kuVUXck5OfoDI2xdy+L6fWOcMhWAHNEwmrgdqciZvu5kCbqVJrybz96FFFrZ
pwN/w53+RjJrFo1TlXctVrz0GdVr1Hkg+ZYDPvhxduFhKqxW/tHggwF7t6N6JaQB
x/VQJ0MLAjrqGhDxMrSLdKr8qF9DwqV2FuiaqxnenZZ2qwoiLL8UkwOgtgqlgk2o
Dbgfe6pUYyBb1CayzA2Gu2G10PzR4JiQQJTLbD9hngj6O6LLr0dc9Z7sy1IW+Tv9
b/qJCWlgF656VZwwf18jkrWTd4fwzAwHAcTR4tFa12IBktjWxvlg98He/5RNfA1v
fMZVdYzOqFiv4UAXKB30oBJJZe2naYBLWlUnXssAn/8rGz8wOlkVVw4oC6Lh4YLz
+O/L5erPKVL1e7KnTcQBO8pD8JmfVW0nR4GR4Avo6OIJ953JiyJuANU+qxUh6mJZ
2UU3Iw7gDRJ+Y3JBQCmUscxspsNBvkoY6z+a/xKN+IBQ5D+EsiNdmNeMstlP0xG1
/sGT+Kipt9Hapa5Qb5f6d+RqHJ8PkrBv0D2v/gLrU8MXvzY1yqM7/Tr3B5urla0g
0ONX5yh7Yh9GGFyMy3MvL3U1q4Xc12mRpJJhbAkgp+J2rdzCmM83rKaqRq05oLn1
wb3iJuR8/AAsCMNOE4WjRuja5921Oqxf4slUitQidhwiadQ3Bo7Q6SLZQTA0HAKE
ZnkRhHG+0gFRftDMhv3IuICAKcqZdMHZUGoyjrfWpQcS1vigj274AAiOb2QVI7hq
HnATtCZy4J4Dp13ECC61eNYWrkhbaVQL4E7394iaLu0nT3dGXYGf7romHFGStPAh
aeithQG0PjEM2ntzMifCOMcdfEWo2rnObGoXmGqMkT6hfUB+x8ufLmxv6AAIR+qk
FElrN9uwKkZvycpsl/3C5NVO5AX0xNYmnRbRfGMhxHNy+CYif2mUHRO7DJKDcEC+
ECojzI+9WIEyZrK3L/ySlmexe/63ERIyjoFgekHSk8+LfQK29zdWd4zAAVywhvCx
9KNzM25BkNg0WGWE51kOX9Me+4/PnZCEuMMsUxa5XqTtCHloqOr/oLHG/54JVd4I
Amtui0tv7itscERgKCeK4BZTRbagbYqqHQmJ3Py+tg2dZbyqjKzMOJZaeelLg+Y4
jdbQIzX516Je+QEOnu1ePJiIU052/1yMcfCeRVKNo5Ixf79AShvGsAl1PUTq6ifu
DTymRH0jN2eedRtmUIqh2CbmmauZnCWU3IgxAIq9IB6V8Y0XIZCFJa/tPOjoWacc
LchlZEboQuubBbiFjv5ZZ6tcoRFL/hh7ffjTxegfYTlPms1AKqhClWwbW/Aqzyh2
QXGaUKEqwCyrGOwOADDlXpEIAYI5UjrJv0odLVFmgfy9h5b6Q1EYkGbnUHVl92Cg
R46cz1D3k5RXokE/7sFnfNyTrV5l8LsqbliDWYSB1vzQni6Fii5ekNEk+TvCxAm0
OeLcy3bZZkDR1cYt9W5Vd2N5zHUVERpgExLaUPlUfmIOqa8lMspsYCN8fSJNPc6G
mmhrbOSAELJ45o6JDm4A+pVz7yhoX8y7kJQPIhzeEbCAtf1hhpjFDDZXacR4GShI
bVCN++UVb5B3MT9t3mTAc9zHjJMekYc+ma/mrMKR2hW+eDeNOzKcJS3f+QIpk0Xi
3GPDhb4bgYlwv5yRjj//l47RPRDee6EQv3wA+9fvjQWBzh+/Z1GXIYc2lV8YaSHE
k+mb2D9sPGVLnVufjWrPVziNQ1Ao2pp8hk31hvDQZLDHxOmI+FOi/fBu68YGauOu
oiLdsKQt/cEkW9iBAMNQvykGEFojAjeulQWZ3/h5ILbMZWCQv4yJuU1xsyEEeDcP
5JNr+hPvj1HCrM6yuO3j+wiUi+f8Ih/LXrl8VHfvo7jA9OAnq8B0AVDVl5DKYKEQ
bM/X5fSnslDxPF/pA6Ynz9T7y5iM97lG29XVoIRaxR/8HclRFou1+jNRAP0T33sj
6KI0LY+xzS7xbiW3srrezIhSrWVyJTZD76wCukT/QBpycGp3erm2GA8DHZEWXmQw
v+dVzy1OCwvQVMduZCYS6VDIrGSk3b392cR91my0TpC8w3b9JH9wpcJfbNWpXluu
wrBOukw+dpiI6Re1wZJ3WVJVgjyNDJoaiCW59R7l7KDjrSY5I7okMj8QLZqkiqyZ
Jr8Q8G4SlU+tCWg//oH+N4GQ1eyVVnu4HBvkYRdoaLFLDOiAtbFreVISrbHlkE/t
jhHEPTOncfh0wOuIQm38yhMnS3Jta9bYcWXcUyLkWTuc8cAmc+nqpvfG34YIMLlr
tmaCp5fqc0BRhClnbmoXuZf2blJ9jsxOFExAHzvs0K0yz9k9i7yXsCZA3Z2nT9G/
5PMyzYlok2EKxPQ5bnHTJUkBObZNLXhebrP7TYoUWKRxIlu+ppXRxcYEv5FKUJD3
BICQ4O6Qqlp0JEcqvK9JCAjWZstIbh5WSaKFLnIp4U+pniUMAhBVF34y686qgBa0
0EqbZeXrw3vpMJ2JyNgQZ9FZoq4QOWiZqRjtImeGhXANsh+Hu5BLCecX7b/P0HX0
s04Lu/GFSNKZZ0WVLLjgMzbq8FjTGYsP0Ym2hhIfSuRT2W+K30YwWn//X9m43ber
POrPUTEMWsOo8Q/XCJV5ePYnl68+29z8qzvdfd9LvWjUmAOD3UEzyU9jKVWBMasD
IiQm1y5GBJTySf4NZKSiTfcMXEyWo/ae69f/7bsBTjNd23gX9vtXptDU8MDVoFWa
xqn5toUaJ0IAfBZMCtAmlkY1qxh5FErML+DLDf1CYDgsHmvOCJiaiK+tB6eOJJC7
0ifvINecmsgSgh7FV12ZOaH9+C5zb+WAt9Hitz4MT1F6Txoqr2vswKG3BKPiXS8M
9EbAiYvQNwlBKs1p/VzZG1pqeiFPx3GFRvzwX3H95jrTnK6WzSlGjzA6BKQtB3ur
ut+Kud2ASCG42pFGVrAR/B+jEwjLzTk5c8ha1fy85mWW8NPOWRrvZZCAFp7ZnuPu
kJ5W63/+WvQHW+jcLKlN4nwouZ5DK4B9bCEICot+Bv7xTIqnd+FqPK0Vid+VLztY
sA30OH+dgE6aqb0Ju+5lgpdpxCRWox0z+9zOGBNvqIiCRIh7Hnvrnh4UyhHLf8dU
4gX1QAGTtvzB5vo626TLxyzDlOp6z1JA5qthjhgLMtmeTSqOEkijp/rLv/dgLfFp
`protect END_PROTECTED
