`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c9YCtqQFJ9It26UulIuPmVIV1fI/EVfvzx356a+ujOhHj8gZB6/fycGHnfH+51Cr
OW56DEkijOis/bMMyjR0u46kTqrt8ZhQya3gL9OUcW2eNr+TDLj86RI78SWiUSKb
rMn8y+7JkN1N3izo9cTJM5xVc0umTCCczuOc7EEl8YFvZ0EyL3cipGXOxseUW5MP
kyOkuUT38uZdI4AAomIjLodEFDe9cYerpIpmapTgGDmut3LU6M3x0L5oF9aOIdKv
ImqmTaHqMTU7FGpqYmjaeOTEfqgyK/seYF6uhAlIytWGS9EmYPeNX/bogrzJiAhB
DKmoD01dT0GTAExwpZThRedIdiUab4WHuK+Z7Uvij+S0W8MTNjlcOjXzjZ1iLXnQ
v18lCSKqRQvEjMlOF2MJhiH775/Bij1Xg6KsVHsmpxKI0upWN/pSbJHE8+Apfdkb
yN+cq0RCWKfR9Q9I/axcgUjU6PKDzCAJeRr2lcaUW7M8QlGwsE4kmOyvmfbJHvzV
BoTRR6vTG88IJUjU6stotIDZw5crOHdWILirkn7hih2gRo2gwHBKQmSYgkeG6ZBg
WLDcRaoTVBSsgWZ3q1W35eC1O44N+w6ALics7YV42sZTewmuBHoRQQO5OzAOyzC5
27NXo//5+FRcI75CBv22ACM5w4oRv95kl4qj7JR/Ow3cZXHPctbL1PAchCZY3smY
TmEyWhYbk7ezv6BXUKR0iH8C0GOdpARegP6PYrbPA9beCY1aGmoJuiy90cY4B+yZ
aNzxIancT9Coo4xuiHTqZdulEfmlFN1QpZElO07cSR2Ddi9G2o6Irn27jyD9eqz1
8IQ7/FU5FqNsqwt2Ymac1rBWGkif8dRdHEyZLVwPOqj7Is0t3YheaKVFpZVKkIHY
2vjMk0f5LbRtOs9wR2XLHmt6j5dRcs5+03QWX1PuUuCHyQLXT3Uz0brRzazTwFXx
jy6aaK93rAF+O5y74AhZLIyJA+xp9Bj/lHJ/p9janJAXOXcXO/nzVHQ8Tiq/WMgH
m+vgUAMDKenieX687AND7NIaIIBTnuJTMAG4rg3MqliDQaDVX+f0dHPHsHyd9mcK
mF720bHg3ufr8H0WHW9OznJPjuvtr6eq7gXfx0EOaPUJVR5iyvh5tfh6GYLf8w/+
WaMErQrvZm/n+q8rg5lQ04uReSgc4Tki4KJ5X1JsRP+wZqIpQLAUZtE4Nw916Sqc
+o43mxa5TqMoXH6f2vOtxD8UEqnc8t4ksYPs8lsvfaURBid/zJXjpj//MEbxnIco
TzqpjyW0KOfXCZeGEkazYV1TIL3Cd7tJm6em9acIm3hNRCM5ye2HtSXvka++IPar
Zlna5af2Ln6nyZdxtEMin1TtqgTKoVZxbjdT+BZWJ1pAW1ibOdZjPM5V6bGsRT70
TFAMxFB3U6Re3Fumf0M6NabkfOIZigUqMyBjPMPtIcRZK1QYHnFHSEiMI/tS/6sk
qUE4v7PVS5o9ZQ6WkjRnXFnrN4xKW0r8GrC9FUMdjFP56Z7QvE7tZjoB8Eblbo1H
dO4cuq85v7eAoJDj3XUTn9ScH1YE/PzXpj7D/rkeTTtGZGBSQIBcAeifKRtAJwcz
7kFfXDfK6y5vtUzGlltbhp7KdU4n50IFrY3Gew2qJ1OM6Krt9g+LtiRAgdBv70Jp
Ma2ShXzNgIvG9DAoMUkA/Kz65PCNdYbrhSfANnFQYoN3K3/N+98x4+ZgnEkje52M
7QicsBySXY0n7/6O2uKjFA39qLT61W+6X0scMk7U96LLgzOZ+K/z7Ct68j91rCNJ
aoRdd5kNAgu4mzkVlqSIW9rX+ug+xPo9YUl5mfs+yC3ZB/sysIFF4nN89fnNRY5F
p0ZUnSaaMMSNV54veBdcVxsgZx513c12hfTuFlb/DHXNo0IiNh9hFA+x5Q1XKR4V
KcKSKrAdqlqEDKDxxoUufHLrgA9a0YxCmzlgmqJx+SF5iDpF+AvNdaLMn4nujvWK
2raYq1il9ziWPjp0TETGwePAH+8nbiCzKX7oA9rjRzTq18eSkG0vejC8OgQBkfwF
wB6wUEq2WCr98KsKAaTneOi3ahEWg2SPu7xu/NM2hP2FJiMNJTEw3QIH1grquc2J
DZ2V4bCPkApRDBjcSnTU6woCvtfg02FpaVwmS/01ovDjRNIZXKodZDlIEwdscypS
qfrbXRMwv8VMAjdCkXAVA3+HsnyBtwBwYAVOLpfGiTz+kQNJXiOeY5wd8MuWfDPI
8QUSVOgBLFrAipJPxmCkVHViNfP9ivMtwG6ryXuu8pU8z83kawWi7tSyYiVzjveD
LaR2My0N1o+G5C7WPpwEiMHFDL2neLRsZWsQhRFksoFMk4qxk3jqWv9K6vRz75Ud
13JZAFMbRpunkiOIVoih1S9N5bIZg4OHGo1NB7jxPv8v5o0skinTqLpIXGELJGAC
suYTY36Yv4PNFY3wLVPfuWYhkRiiiPNxDaDlUUcSLlHOvoAjvAcKdGS6LvrB5ysD
5UnlBzTbS0600Yf994dy7m+rAbr5CpBp6qdV/4WD19tokx8OmfzOgRgcA0B7dFjw
wgzjcKsD9VFsDzConuX09KFwD3vtAYPzO9u0naGjaG8zKhHCqZjWFk1C7h3kYC5x
HGM9G7MjxMNxS2C8gXRNzpoB6MZeRCjaID2ZCtMIutVzIudwUbs8LYe4Y2Ucvi4S
rGnqi8b7bqFIw6oaP82/UFeOHKuGdYYnHqMu4XqY9NVxxq8I3IwdVA9lbFWw/p07
lx1QFJ079zJT3LsVb2QzFrqx0kB0A4lCBpntrZj/HaxwKPXjbHIwZWAO7T/kGs/3
4p9M3xqbTHlDES1nPSAP1I8/Q2ouwdesqlgPXptkRaJR7YZUvH4bf3B6OF2rAdC1
TL1qh+ovUk/Bi/3eJy0ZrjeVt1UNsRlBGgjc2KT9+edIwRCobjnfgsJ/A+F1U5wY
DohBusJBIoeV6zoQXbKVU+RnJn4YI1R7wr/BvNhX3NAUKuFFepsuEev0Pj1wmQMp
cSOPOrOdgLeenGgLH07ZdnNqz2cn2B+msJSroLK5Bd/J+etwN58L4C0aRmEROqGy
sQPQf5l+bUBqMaoyKbWVUXoLVPEHxTV06yFiHuvFSfELs7OM/6WRbRM6lGWP//GF
H7YKvB8kB2rcy8+FAFvcsS+LkNucvF595rVOqIG5TfELbWoijy6TG/smhScQNY5v
GWI+6+KAoQ6lOcTy6UM2wAhrIO4NVOOmA2WUkAVgST4JXBumnNYDa5E7bp2vWtcj
UsxsVm1diACtAAH3fweaCyMklc4xWJhG8rJANcMA6Vvfxlz/phMv/BR4QPzys5PL
n7otCrN1d2oskUGRcjhSr8XodvrKGzQjs2Nn2xrN1HUsK2xJ5zXqzWasEqIiLbHG
bh1vQivTGp/Rt2jgFf6l15EDMfnAJMjW6ATUVlQdbUT8yAZH3dYcBqvnlOH1ZNo1
7m/ut1emQGdpLiRSzc9RDIdUTlt+EX7k5LbhFpU+dZGAv+WoA7iaBhvVDrSP/TZL
vJJ1PP9bkj1q/zuk8NtMbqCcSqFyq8bQoQ14NbkY0jOg8IplV7pAB9of9u7KdTOT
1y5aShfDsh9L6YVF8UOyY1WeTWknvWK1EYTgh0GjSu41twkScAZF6EUA2ZoeFK+L
WYZdjOfHKrrJYnGVj0bUEwWDP9qGmgybD1HbTzmRdaQftadqFAbdcTX08ozRw0IH
gZFu3jtmZp9mgeYBjPJxzSWZuqRowSCBVxNZ4fGbR206xsK/QGHCVo0MAzyR54ol
TI3FsEJw91P5kowOMS5SJl/cjJIPUZVA4mEe/IMm6rW91D7gO1xOyO32XKIZULD1
x+iW6xK4Y/vTO7r7HH286XiHkKg5nD1L/Q00kNxKdCDK5knL0LafuUIvu+8U4qGD
RzbKKHWGsYl+lpdtZ9UzyasqTdxch7lu1fWBE5dMOBfvgjfPdgHpbQwkycheDssj
ZEtDaLnGBzx6eRGCgyWNYsbuW93R51E2EEysschv9lTFyna1V3GigfPC2E4qcXzC
vKN6OmaPWI/QMnVXZ0ZKCpu71Avj7ZSAq01YvV49Yihk/FqZ9r6W11kV4CNRGVak
P37DaFlZcHbPHZlfe9ILsXBPDhWv+hV+bonHZHVkBV+Hfdp5IegVyQwx77tzc2LH
MBOCxG4YJ7Ee9vD+H15Du2tv8h1rMgyu9pQh5Prg1kNEUeYporO8EJynhreqzuHP
giLtsjfFj70HMSI2zK/ISHGYOGklQNyvkyBuIdIvUH2GtyR1lKImj/7dx//cT2Ci
h/ZxR5qJJ1JKRX24ZCSe6qX3vX4cppeF83F03fSv3ixx5enECnGxW+hUvDuELdnX
igEB8eaN6OMFE1Reg1Lb6gJSteagkhS6RW6cO6S7YDcmwU8pisTFXb255W6uxdAD
8LsMJW0scLBLKhOZW0eELx7GmnFMC9XDNvrB5y1UIi6lhgI1F082HcfcKeLPcx5l
qo5BfnBPrZ/xzrbrCNdbjt7OowUkJfQYaR/Aj0d2ykKjqfI1UASeTXIwrkNKImOx
j82VlIFThRY2SE4HpfMEymxONjcLUj/CNdhQ/Dl3O1DtIqwLnEC385ttTZnu9uFI
5xRYd5m7dDKmqMR5TNBQrBYswbz9bx8Ely3ATdibi7VqYVrn6A7duApGhj/qjbHP
x2PxEgJlf2k4SUjyD3vNA142CHMCjP6ttO4W1LfGGUXksEaSzPk2usNIu8r2GGoK
6PqCa2g7BCjzqztHFt8BTUIpU6sNqIAkt9mLPLCV3xNMAVx9Cf7x3vzTIpqjeaYV
RoUJLsYTfuFETiZHw1lnWzbCFaLXpjH4gAH9S/7eycsPwPWRXkEnmoTTvL5DXv9a
jziwm8OHHtxv77zTCBy9h93gxPExYUjuyEFStlRf9Kl7xEP9fKiCoxYUa9YK2nG3
R2OT0aBzU3ZdzXVuUFc+zPLs0hNbekDpl//ZRzhK5xQjpx1Ku7MC4fo8JqiRW6Qj
jXZyJOEZ04ncEx1ZOTlBX7j2fifoJxfrL3YQmUOvVU0u6R/b87f5T2CiBEwos1pk
kSCszj7bdfTLTdviN7p6h/wuIHGstIDfu7zlN5q+aZeOYIjgN3AYDm6ggaBdXeqQ
88PNT5NstudUqaCP0KXVY3aLzRL4eysBpJDjI8Q1q6+lgjjCgiMirT1jSdhlkkMy
cZJslaBz0AYGFNM1a4uTRd9KnnEH7aPbkwoY4wEey++9gL7KbUsXTxR61qlUo0+1
FxGkHpj8byxi21M2xnsgSm8yJhGMW+ykfQuQLXx0R7ZosgFfyYy+CwoqCD1Z/V6n
wv9odeWSY89zhXixd7TW03NIzoJ+A0LS3zPWVsQGbOYCXa2tEbch0KZI4OxaLjs1
WZS9fy48HhO19IuwZhNFYNKlqE5xhtbjLaWfZVdZOfV1MMEvhI73F+VnYp1+QVZu
WXa13kRsZUZeyyA3pHFfXJ5kkGhhPj7QBZJCy0a+GmiXmKqExMtmPNGxfoV6F07W
fimSMXYZ8nGfZnFBaDahFS5vVs/9lpMS+ebv8B2J76NGK1DeVxHaEti9260w1lK7
EqInkJpLfyhOtMBchrW/Z+P34zJqi0MQ4QYaSRu5hGxvEnJEnEXqB5SfyxP4nqwO
f03gkPHcLjnsmPH64jUYig==
`protect END_PROTECTED
