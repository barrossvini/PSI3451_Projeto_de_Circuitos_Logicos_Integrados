`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTb+lkR82rNPfXdh8zu5X9ZULBCxhDP69et38kiHd4EZJEkxM8iPTbPdqZ9TYS61
iMLj9rPt3PRm5lE3qwGBe8pgeVxKCGTZKDcj4+Giu5ydjmVl2/wAOviCZ1zn0Ntd
ksf8ysnr3cqCQlUw5sVuEcoRgCDoyL5eKqRIdbOTqoFWJYHKamiqloYdwTnZ2XFx
FzQi1vrQtBYnvr38ES6HnRmmm3Uc+J3i6c4NAxM52lRdIvGWf54tUoE3fJlxrrbC
4ozIp9dKqcdl/Ht+WEdwtusL8SwHElHSov0kZwoNzJyAsW799C7Xg/x4coct+zK7
tL2aPV5I1vbsgvXJ87vagmmL37jUewuv8wYPPd0JVQznUJPwkSf1Cwd1DjKHjLb7
pHDtdBkgPmViYcR0eZr1HseGbkqPHuwBNhBLdybDm4WGQv77gDJx2s8F/JwNIrth
8KeDtSJnDZ5R13287rle6xlb8aTKW+Ng3z4UqiIfR9hCNEPuAv4RTsUoAeWlcu9f
wf+5/A+UdmsxFQ7CtK4gbmoSHVcU4/8Bh5zbOqM1JIkq4uzHADlj1NSXM4KS1DQx
sYfOptxLSwBDUjauyvyWh0qxkeIqVHZZGtjn7cxDgFCYjn1xuZwffyYbxtGfZQ8H
alzQwd1GvlYP+/hfpkGFPwypuUWTm0E8/41nTckDfbAouZX5a77ghD3dFPLEhz90
Wh6kQdWIslo02WEZQTEJ/mkIvs6clyFRMH1N8LetfHFlRLz24vHCl2vqJBRE7x8K
5PsEPVLfiRMZnl8ivAnSWeT6V7dYpwle4eAj0fBZJTBrkgyLDEfhNN36rUfaZYpk
z5khDng9/BwxOS4VKNznjQAkrRX3kLMSVzjJL+xbSGXJTNkL3MP2UIOpdcyfOYGp
UyGxsaDEO/SjsmD0CprxAif/iOWC1LWHpjn2SIeCdECE9MAE5Pi239NPm2RnBaA6
SoC4E35n/v7nIOOOP/k6pCWuNeT9jWvxEFBv2ENOh5YrCsfxBb3a/B8zlcmv89k2
+P3bQPbjAubs0uyhBGWCz12paLvQfopIRCsMj66mbxlcLM/8s4Ehx0Qg3o543sLK
vFuy5HAufIpBjYJIlKSj3r1ilmcgmCBau3CvvZH797BhJMCC38izwa+CQ9nVlZup
2yg2QatgoPWO+gy6pYHjzQsg7pX/NZVaUve9aD4dM1yAkHGV7MY5HfIqpdFDrfg2
kRw1z+ou9+USzTmD+7Eud55BDCqNTzaPa70vocnPOnPs85EIfuwuywfvKner3jl2
QInQKR+AzpTnkTcr/eJICJ1HynhnQpcRTGAqsjeAuG7VkrcjsVXntMTt8Ln141nJ
fIddNhYcZnJYD5SxUYztObpf2zb64Ojq7RuMROSgHk9JFvyCUdI3lhMy1isp8XWX
+1zSxcPraTzfHJads8ZN4v4teXi4YRb2eWxMTXyil9Kl8hqVxZKxoHHy1oUsNDNi
7ZhVrjHQlDbvcCDk1sAOrnfB0sWet0UQefmPsv+zTdv4INaVf0HTn2EBSN98ZeWT
MdsERjIh+HMyKeqQQczOaz9I+FXbX71C425LJykbLWb/zSCZ4/fIo2UeZImkrnYN
CsmoH2dulsrDuU4Q62imuvuoShDb5howFldmbmSZsjfaNXWm221tAEoOT7XOz8nU
icOrP/Yi8eBCxCLG1KG7+Hk3IeWVoww3CbrqYbNog1uLo1/hsoDFY9KqTjTN4tTH
YTXP5LXPN+kOf7wBoW3qx2sZ6k+w41JYabdsg1r9/qg=
`protect END_PROTECTED
