`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDMk93NIlBhse1Pih0LdIc3ofyAHUBhYgGdUagMpbyomxo/8ZF3gBME4L6edVnC/
9y3+FUaiQEc5eaaT9pFnK19ktnVM0bBonSHELG7Z1HchUjKbbJjl53ZSM95C+SLh
SV6OTUBW2Bh3z1Ef36z5z7FYqJj/bJke1ns6s1BNL/lI6rqfxOHYON9ygZ7Y1B+r
VLvcVGlour41q9zLZPpEKFfF4GeX/W28Rl2UzMMQ8l6YRMOrKttImzTu4PeQkJzm
f9Ago4EGntncshl5MkKhOAAtiDw/ROFfNbhx/Qsp2k545yaE93HZ55RIyC5xomTU
+d8enRcoG4XGgH539Ha30tbCM2Di9F3+Vjv1jqekgI6kUXy6JC8siF2/7SyrSmUM
pR4gadnMtSk+jRZGbzt2MiJx8O5gbRKzfdhrjlGVVl5PlBTqurP8jJnYWaa+QyHB
AhKtnAgrPtws8vCjL1XvVL/mC95lsehsSiOJ0yWY7F66CU5klhj+1GaWcBkOs/kn
CRdh8Ac/6C+N737iv+/FIVqC/vk0155nBT9kw9bporL+/4CVZFwZZqRRC3TcaFkp
/03gIIqJP6LkDctsipyD0cp645UMGo7EllEa0g5+A7XgwT36j6D2PnmtiO1TlOs/
gVVT4h/Gn7YEeeO/fq/qCbl5oph1WoZJ1067vL2AYJmDvNsTlct/h89EVuvwdevx
l/bSF/KczP1R+QrzWvEZSL0yggaFiyDTmfZpH5sr+Z0gAsZFqhXt/Jv2+Fq2NQ+9
wOka+mqM4oAHG8OsXnFh9lpWFR9/QNDU/I4bmocyVdR9vlGYhjmfPIC9e9E4lf/8
gqyLSU9BaVv7xS4CI27huA==
`protect END_PROTECTED
