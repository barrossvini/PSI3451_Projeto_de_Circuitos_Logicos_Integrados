`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDNj/SVKL1/6p1htUU1/pa2xOJGuzo9BPcIpZMPzkyMAY8qrxopAxIeqaLEEnvhe
bTdCsHjMP/Nr95Pxk56zwrUkl4C+E/PwYgYFiyX85+OFRDxYD8uaExMp3PlZognl
qmNq1XmKTyl+oM3g3+nVl/DHOkxV0eIkEccrrnWA646bbXsoboa34mNk8u0zTDoU
9QHWYAqDQLv10b/X5YllxA0uarftneGrmT1RpYYWgv17ulOEijgbcfMzTrfNBmBo
GtwJ+CC1fLv/kVeNy5EYht5MKOubrBU36bBTi4WliqNTmkD2b3umxUQ9KVr2tocx
hnm5S5QiIosZjpvlUUrQhdUbMkq3ldo43S7emfnCsdDtDAQpkIs9cK2C5ZkKuwoa
Ef64XrDQLi0xD6skJ5exXw==
`protect END_PROTECTED
