`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yoENkN5VwmrZt0tXRJjVtlnNeEGn/Lba4W91DilzbYSJwU8o/1J9nISRkR/dzetM
2bknougeUsGalNhSnTPZWVbe5PZztwOYBw3Io6Iw0PTSWSp4uENJwtxb3zCuYuAc
SGLz0q3LDJSi+tDsEb7l/n6fevtyXunl62i9IEYkXhVdAB3RGiyjPvbwXjmBr8iB
`protect END_PROTECTED
