`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8OUpaN3Box6btt8EfSlo9YCj1QttTA4JNRhdxPYVGOJUmLoIT6JKxkjqt/TtVzv1
Yh7sYjr5212QhC5k3v11Yxli2cPCwXZg/3H8MHBIYdZ/NxmevxpdtwcwFFpiRjWs
/WGg741DIJKvk6J3PSYkhNI1QNpP3saZSiH1+ZKL41mP75pFc78XaszZWZtVBveu
InK6p+h3S45f/4X2hDyfRy+hnUnszYL0nJVqexKs2YfzYkdDErMX+VGbQOTTePwS
sYbUpww5dEVsRZBkYXRZrImFYh+d9L+wEaO/VAVKrRsp2v+PrN8Kmz5hP/5Oh3l0
7TSzZsyFGK7WZmCZJoBBrq4pjIdMFLGvUZnxH67FkVUJQCSZP7cbN7STXbELZ8FI
ss5/9ncI/Fpc2SRQ+Rtqgq8+ciSbVS/d/wFpDYcXbsWCifQEkVPjW8bbed8L/IMt
7D6TOnbOCQrhsQK4HVHvMtwpFCMgizNIYVtvg75OWljTJ3OjfNtHT+3twmPDruGt
LirtB6Pvln6pHKU2HOwz2Cgc03jYB8N9plgb3fcqaT8JN8lmKO6ZLOd8U9GH2Ys5
/lFvs6hvj1DNL/A3p3W3ysiXUQNADkg803UeAAtZxU6cRZCGTma8F5Fn4sdmQYD9
koJATFYbve+arMmiLfTfv9FfKZIov+/+s9E0KH723opOmt3+ssGcF0y33x2CuoCH
ROd+JXTC55Jdyh29dD1117K0fuqO7ZLGo2z4cSEq95LIape1gZaijMgUvEHAf/+r
9UUwUL+Yc3Ln5qJacTDWoiotzl8ArLBfAcLCdA1HTntth0tM2gEsDzkNYap1gWaW
eGORGBYQmZp67pdPG7nX34P0VoLP887EKksaGXDcSLN+qLttCcc5Vx4+mTOdV6ip
C0fm5ACD5HNka1GTrZ5iCgnmpPQkgI5Z8G7ZLuXb9Ls7KZP8ilmozdd+k+TCDtq+
KCQyBMw4ctdBJV/epyQA7lZ1OWzFalPDUJO2yrQJFpCi4NYiC7REDgpfBAlK3Mfp
M6QhaRr0+JbZbdZmfgQgrA==
`protect END_PROTECTED
