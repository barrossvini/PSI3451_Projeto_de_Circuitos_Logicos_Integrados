`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPp1LjUZYph3+xD0jjiyFucotf2tj9RTBpTsWOyERTqUSN0+38Etz+/wKheTP8FO
azcXEAJ8CYAgwYxVBvjaC3eeXwKs39doXSoVr2ReSjGF/xCmlpFoUQv4wW2XOkdd
3kzlyUA0VtDG1Vrs9VEZ3vv2sYVEh/OTrMBJttY2ugB4kMtllAzjYj0Gd8yoy4bn
8kx4XRXwlaT97mHLm8jJB8GBTQKBQY1SDhz4DS4SAnK2I3J+U7wa/QRyWPIkwW02
nVIWo1D2duu3zdkhp/FneXxBVn+wtbixDamHVFjXIfFYPrJNr5twB1kggjGKnIut
uPyW5UsYusuCSr93Gn23bhhrh3UxxGoyox6/Zc/edaAisl6Cc5RPasn2xuD8brv2
W/gSP4WOT1m+JPoopxvfb9Cx/E8FQAF9VJuUAEAnsmTIuievSCGgjKeDm5+pKtAv
LpbMfgcL4sgguNPsiPwfSNdeXU46MOcUtiX/WAFdkExyQCx/XfwXM7YnvQQrnxkx
anmFiFiRndy55hkx61ZMiMCeUr2J9OtD/wMt4FQ8EGVs6Hos01Cw4d5+YG1FDjwi
Jcc3MEmjRwvG5TzMbjUCQ1DivPXe8XdELCtEcsVb2z4Tfy08aOIAcVzr9AnU1bNS
HK5bZgtfCjVmWF25gsEpKxJwsl06jNlM4VvGI/d2W3ERLyjPDG+p/h9SY8EbvM1d
RzaTj7EJnlL9pNNabHGNEe2pio0ERwWGTgOJR2KQWhQFmsMGTgMwWZ6xmIOtNmK0
z5KkjYvMwaApVxBDoEsDtREQyfN7HP/AbKuC6s6clZsGerqrypMxTiaLSmrrB4dd
b6Mq9S2htx7Kds8E1BmMx7ft0tbjn9gNnwmL/aVLKnREPz6Sxmi6zQl1Aeh+OpjN
bRW7y4ZbYW/9benEAlr/na5RikW1Gv/b2L49dZWRNYsx0IP3bjL/sWGEI1nfsD4c
XGf1iy52a4A5ORT9+V7LxNPu0h9An1zdohUyFzHe+GESSMgE7i7ORzR99835rE1G
qi9/0lgFs+YdN3U8op6i4HdPRV1ZxzTytg9v6+L9H/y3ExBFvVOqPMMbwDfMF3s1
OzV/dOkT67hrj7uK7IBSFCTXFX69Ayde13X0tjQlUWKZ8mIW3k6fMissZ1EPTkqN
QI8ewTQJcQ75f+C7RqyhOjDyqfqm9umJ81ppL41FE0FcM+owa3W5gWyRqI/DvMIQ
mcLzMRn0nEDRK5XpoPywjhsXuA/pf6NOxLLYnQmGbWhKul8tmLSASlnppHSFFqA5
QXhGfc0qh9ofj0JL/vJIK+YfsGQezAreUgMKQjlf9TSfAitSCx7TId/4biOrshYM
7qTHWFrwlGBaElteZQhBFxmHMUbxY4BE3/SxWS8FCiOjmpjoi4IeFegfv6EPRgmt
TbsqI32yqMpki6USWlzYdT0QpHwE8tre7DNf+ql5suSRgasrBxcTlQEmYrsOdQwI
NZ4j3XfIbqfZk+1w0QHnYRyno4IsUr69NlnT/FyBKkYnWDGYNN7gDcgX0B/srd11
pIUztyaKxc7uqY1jNF0nhdMWezZvLip4vBIBuyH7SZDMrb+NgqHhha9GQDoy9/hi
B03KA0QMDVrZiBC8erNGMrlBKd/LuGcnzuQWY0xvekWTotn/OBrywrYdmxFoK2Ng
DykiN8LhpsVwiYMY2IzYCF3mw8JLh3sBBlucgbzoCExZqMKmEWOX0MsBkw4+UK/S
3/XicSgU5TnxfxdbrMZViZEQwg1KNWdXP5vyKbnEkwvv9Fwytf1OGEkzXLE+GHWA
6yGZJCDcJ4xgMRgcpuQE8DA9+yc1/D1DnUvL3CHRSE40GV6SJsiHcHRXeTZqNyeU
tohSWNsamyAMpVh68wSk0IOpx/Xg7/Ehh+Rk+T1KjDebAE9w4KlaUBobFV1I6O+e
Q6AwdwY/RzJu2HFKgHem96di9dt6yA065mUDfQMapd8BJ3Zc9GWUeDsdqC8ZpIi+
eax6YNnWKXf1xerXEQfrP7DqFFpAJTGL91/3OsBsXnDjZIsQMQBHY06OK6gwPdzI
MaHjiNWCi6nlYkamNqrVNRY0pEDFxwQ3IKQgAzJ8ObDBZgSW8ifl/eHo8VbB64YP
1zg+rASN6/HiZqvjGg+CakKcmTnFPvufsVvxG+ZOxF1SNnynNgVQkrLxvMsCDliF
jRyn+dpWuvd//8x5zGkApIrNuN6/2c3ItmQvRqix5oDhHVr9COz7FMTvlLFKb5UR
AlJSuxH1NFNwaNBffzmDKF6S2Kab7I2WoWrmcIyyzqjOgIpzE9oIJBK78thfE9wb
QIkR8XUNJavu3Dlius1rsVPp9l1ndS/ltSYtj8ucrShRdPsB0+KWjy2hl9rO0jwj
AcniTJedAJwsw4N3HFFTjlvReBKxLsXLJHeIeCKp+E5VpKQCDIO0cNlAXSsibfRs
LKnEz+4m/sQKq2yWeB1DUbClrXDEsRweHpNrYGmNr8RAsCWboLqw53xzshV2CvJV
caSFuKtgqeC594+EDjeZpW9yhH+Atxxsjm6cXvruMSMspaCkzeqyy0ABPHP/e69A
UAzOmv8qFAZGtTeGY+vG8vNMPPSlUW8BkscbS6GaPQ2FcBsuVzKYlYMqVHEwt1y5
uVXta9pVLTlgcvGsUhz+w/Wc9eKNnohMZztWTW+jhiJZdyn9qUgmSkOAFWM6O4Hl
SDX34xW8jeZikL3VLJgfaoA8Ir7fEb8UcusLmzD6uLFKv5LQpeYAfuBXyXv4cQam
gjDBpNLXMKDU62E1CdqTSJDeZg41kiL3CEaqUH1XS2TRceoixp7uYuy3o4RqbRJY
ul+HnTYtcCrURL97w9/7nF0PSL8/2s8BY/PrPJSCOr9TZs6PcQC2vIL0FkVSO7MX
y7upQv5x2MxtR7fY3y5q0eE3m4UM8sIPK2uNGRCslwcWlBmN4nYjFam473eSnNyq
neFWoDRJYKmG3AfuZXxKpA0wpB8Ck6PqmwLK0KpsCQiKqjh/hF2fHt/T6Gt2HGRH
BgSeCsqxqhUyD4m+fY9K3babrR0QoZCE6d7A1+gqOwYPhUV3hqYdEpgtTwuQEYJU
vCFJgAwA9nrQ9S2zZSeStVVd3qxOmf6wJ0stTyJJo98R4nOlbJE479Ukg9gRTpSG
LZx3MZbp/wrqH2s6LWvP1xDNav/mvLaK/9tLJ3kQKqVFLx9chL1HNuhJ/l13xAx7
RzAxMkWsBvyNEjk3RBultUVHSedL0p3AYXxD8T75y3MeU9f90dGgV8rAIDW7nLxx
Qy+Cum9Mf2Yk3QT1FS1fnGK/AaEdLAaEB1JmZ0Fn0s/jf27ejY2+vv6x05wjmjDt
njjvb9woSzIn02K2GN+L72EiwapCKgUCNPK31cGqJyUlorl6uS+c3geYLfmD+yBV
4mqefy8N2VjFqPdOecWzKP7ETzeJxjXZdogBb10sWfwJdB207BtU0Zz6qgJit/Hy
6HRGQ+9W0hGN3zN6CmHfRHw4e9oUwQsFH76sZMdMflSrrBLpuU0+njUVzHIeh8ta
DqndhXT9vAAa6IwZbZFEnAN+E3eH/P8ieQVrfPn6OY9arIUKmUF4R8xOwkimHWWN
n/LfTNFfwM+0BemeZcj4o+WmhB1tk4JVFWEu5LBsWLV4h6p1KThhM74Cr8pOlrZ0
omdOkrTR97yc9rLSO0hILGwHUyHIWEU7/hpIo620anwJwQlsY/UnoBG7wLQDAs44
dVr039gidnJ/H23H8ns7/kCNB33lo0FQS7B7aKyd0kDdeHB82uaQVP3g4Yto7FEB
fcrTwj6pfseQpmsRg8CYsbtQ5INGxSM1xO/e5G/cFA6hlT8HPOik9rRFR6xQS1uE
oSDN3F56jqhtWybXm8uZ8fm9oTQkIpTl08nlmuwfaqZuEhQdM6qn9ujl25wo2SBw
XUzxgC+CcP8I+R+E8cHYUIInwMjKgV8OhSk6CDgChkHJBZ9No9gD4HVrJUZF/Pos
VvYmVoeY9Igm5pNlwJcrmcDW+ViOSuFOTkAmZA4aAUgEXFsFlhvSV4QluK5SpE9+
ntKO8UrRbs6NlaDqS4GFLsf/WVXSWTzwuVD0y9EwE4gh+Unpv8Q3atzJrMiFpGw5
z+xly8VHzpuc/lA288aAZBBkidVmYGNf2wk0mIFz4qpOjU482jloZe7XD5y6HMnT
Ebu1hdDaAZC6JEfyaO+khY+lhmc0MTnAW3xsSlCM5i2uDYematPo4u0mjtIkxRGW
8d6MI9k9Pjdy9OEXA3z8Pfqwzj/6+Diev42OmxwdTLNQ/1b7siM4s9XiE8Ds1CY3
Oy8/xBf3NhXQXgB1mh7VuSSvI+AAWrC4iTL0ngnAS9Zp8q5oXYyyxIL9LYF2HfgL
zGbgwnYo55pyQRMYDn3508qAfsqi3zmMLKITEhVgup+FvQmuq33Ip1i2/SRXQZ7H
hBSJ36zkzzr1LFsUyPiIOv8dbRQ7yNzCcuS3GPSxJsJplj5RbwCzTWhEq7cFg1cG
0fad5j4/VxPjPz5y86EWWOxenaOltOmuCAXwnDoFaEekqcF+7IvGJgd+Htq7Wzzr
Dopa6h036O7Dd5PMQkSFZFvlOMgxssaEp2AWBwt6WZCEY0TlS+ZVj1AP41jiJrmM
Xiv9dvQvhSh6Fg1R7HIGx827ThCMHkdJ8aJdMvpJjsN7JoeyHscLlEMpOxwSDX5P
DG7SezNF9CSGSimgn835mlJsRhxH5PyQKFe1YfjARkNXep4t2jmRoVeQqARep/fQ
c/zDmA7s8GB8enZpnxqXOykcp62WjTHFeqnDgyw5KMZzSRn6n1LJMyhhqdf4VNga
5OlQRTExjXkhKrMlLQTmPb70SG9alEU6JYXivBqIa5yzwqqUmPP56r+HrzOR3aA5
AZiowiFXcaQlMNyIzqxzdODKjmBAU61rumTvZh26FeHdh0p8f5QqQWWa0uGvGBdH
5quQuDkoIFv8KDrZqv2HvLtbw/Tyh4Rah7QnWFVcbNGFOfaGMDMzX517ZB9kq7p9
ftPAoTg7ECoIwyzChSD8pft+D1E5+hH8rW10G27LAW7RbyUsf9a81LpVE44f+Wev
kwX7KesFVc77miEr7Py4/fP2XLNmSCm9OnXL3QR4xT/fFgTNnW/Uy7q2KGeqzK6D
/15qFGGswbnUG06Tj3erUdXPOO1bd2pzxI9n+Bq8wB2N+Pp0PpF6imw3D6b1Kv2P
Gy3OBJJMyEreF6RN10pUXVkcTxc+M+1jEJpMs3eFAwJJ1H9dJSTOr4jlh+w9kv+v
vviRQrV5WJ7MaFXyoR6CssR0UihWFq150wb00gNHAR8VUCA1Aji216JP41bA3FEL
FkNjKdCc8P0+SO02aOH+09EACzMWXagUjRwFL2YXodP43NbXUOhu23N0htE3Aq5o
psoNV8VYiE/6tWu/ZWCoBlGsBuWoGWXifq3gDovTgjnKaA5XEZrN4iGFFxnF9V5W
KoXDgiVAzjpmwWkNQcmss46CPJe0zPb8os2pERRmr4z3OLtOdn2RqAsJmpitfyww
E8LjHz1x/5vJQ3li2H+gNX1WVacWXnzrlTf0YlaIhf0d8ys2BZgO0hAGq2LVLCCu
9MHTVf6oDDJcgkh0NwEUn2kWpxc1dawuVli8gNzzYsFryRASz/XefSN568RPD/dP
A6L0zBZ707VBBk+D/DHRilLrkth99PnutlnH/cNJP0Rq69KITC7xpOeBXnkao6ou
hjM2ztGvh1rMX2tg4kgJh5N9G3mw3tzskc4+QjhFpyvxmSGt27NXO0Es7m6ZoLn+
aq99dsBAhN6Azxm6TU+4YKKUfKIFTqRPVWfyOAKkoHraarpR291LNysOp1tN94TT
cciRaAjdMiedefRmVgP9aaJMykEM7Gg5uYuXzgOJgw5sSXJXAYSfgQYKFsC5QdLa
X34UjKrGJTF3mBr5lQJholV9GhXCfeNb/xWEERZusSoixgM4x+dctvDdngLluGT7
WoywQwhIXWo7+pHpyJLcyCcBUcJe0sjnv+SyhPg6/BAKBJZEERibULNyCxlBo8is
JRLmLVl/QRPvvztOxjSDKwwkTv+wFuTAoYmnviC4k6LLY8OCv7X2OJvTlNtKNP2I
Osc+6nAbs5IUbniixdXMinmSh1MYUGTfaaQiBlVFxOMO6R6fmGVY5EHxp8yEvQD+
W/wu81tHnpdbu5M5rycbxGoNi4asbljiQvpNDN5KdlG8pfLvcTL75kOW27pv3NMr
gnlae32wnMhaHKbG9GVUmfEwswxxjPW3S0ZT/5OyQTTg9FFKf7G0A1jXbdNRY0mR
LQN2ltF4GLzUBlblVXGUIaz1O6s00z/xKoRUCWS7xfXRvhxcCyTSPaFv440Qx0Wb
OiUiyHP0cqe24+jBky8RS3lIy1YvW6vhUTF+Fcu16uKZPEk7T6e77NEWIAmwYxjB
ofSC9unNt2cOHLDRcKKC++2vLRMxrx+l5H62E+7uV5agjeXR/GVF75ksn0RXGWY9
ot6gaJuG9QZzYYbTbo/J3Ekwju5j2mCO5VqwAD2DfvLmtuXotEo1NOtO/plFOoMS
IiIAJv5qgjvUemI3HCSuUsYBbvaddvbcWbGTefUo5+QWIvXBBuxIels76nTfsdnf
p3K1H2QcHXOOnoRvPK6Nf/fpx4485iNIcf+Bt4WCwyculMNcVwTTY10NTjy1ZaHu
/X+tmni6oWLFr+pV2IqwEr+9YsoVJWCXhzCmDv9w1dHVv9fVY2W2+CpFxLKj+Pgr
p+yO+bQOdB2fyhzLO+cvhkTn3xKg2nPa4qvQrQ6UgTulcJqtf7w0br5f5Kf4IOH6
VJ446hX68IABxcyZ9Ie3vm0Ker2V7hOhtBvJcfiE/I8U6Qhb2LNveol963cKVqKD
0wwVrk4eo1Fj+uji3peeSloO85pqKt8M7KbRwDqq+Qf9IvgfPBxuGcH50627SBDS
P0xhN7EgK48Si62V3ICYxeRyjQ7KSKArSjK+ubVxibIEuMJ7fqrO/iE4LMrFzL13
immKrLWKew831gmtZQfIOaaNM1YbijSrRFs6hxW4NVuy1MRn+IhtFm6R9wyguRgI
9XyWUqbZSAoulEX4xFQxQIkzN9E+DJhR6QDcdv0aIlan2ZbAhYv653Fkn5mJzmdp
ypZqcQBWI6wkEAVZi4IsjYyZYJFlWhBZm/kPY9KBagnCEQ7KYcn5URAmn9WpvOtP
n50mKl+gQ8WmIvCAPOKD/zBMhc8ZgA+X1rn98+OMq+17UaLkFtDyBgw70b+NvDFj
KmpTUU3StYJc1JExgQc/byXGRcuHoLoW1dY+a942jcvWUebEKsr+MF3Vm4Tc5yA+
19GiVhcIBhXUF0xp+rUBWR3SD6XQds2yoT09DKYe1jmeFRXZIVax5E5eyehm8GVU
EduVTlsal9ban1ZwhAkTERlkSif0O0bRHj7vq6eywMcK8I3rOK+mO6N7cGktOvoQ
y2Uqc8d4VDp/M+Hlix+vOekTJF9o9j4kYKMSwLiG340REMpWQ86jEteta+1MjeM4
xfWYiUqD6gBXaOmZ0MnHXHETQdLuWW5DwoezQzjHDomzJHaTFJht2qR7TtiEBTdp
W+P6h7PGK4W/K2Gu96L0g4/T9Iyj7Uv1Q9UrhtnmRMRssOcTH/b5BT2SQach8V0I
1aaSzO4p7XyrkS/BS9apee/20kkv3xlx5I6qMRJuC+bKp4mFhEEjgB6l2rXf4uRM
td4RwTvHeKp9RedPjglV3KGR/EWXxLQgyzg4a+nfZLrT+AvK+JLACMY3WWIyYg4/
3SynOsE8wB73Vc9EqDCk2K7tohj3vvCCYW7hn0qTOzZ6DlOJeS/MaSD9qg+JEVMu
YtJR/n9LXsVVMU24mzwavSq7y8uh8dRBvJBDWoIPeIDPq+HNXfWVyxBvxqCi7buE
R++uxEvfW1M40y7NNioB5tx5Rd+Q9zZjdfSTs9EG7jTxa6v7m7zR39p16wRkqsUX
fCZTCwDr+wCOvvFgGmeaWvUBhYFCnx5MEAetLoAhKdEqTuxtTp7REoX/GCuONQxL
0d2jkzqiTRLUshpBoXARLk9cEEgA9eYFXonFx2Yj7hFzCGHvEGY2nTPrc0MNI/PR
59CfLkJL2lormSxagUN5EMte0CaxwB+5hjmLQRhOKbYU9M54lf+ArrGaQdapLMKe
PKwu+vIx1baM4FtBZTw60WGvAk5VD+JvThXLlW2tfbtJCuSN5lU7P4IEotlKl0cs
rIA2fOigwPNg+7GTPrm9flHoDDVDACle3W5bXV06U4SPv7V6FHKKAVbcsqFNoLax
QgRZMZAOTYEhgsVVnKXwv7LxvzCS6HsdQkx9mvK0cAuKbn8wVDXnfIPidaNAjED5
LpcbNSRSwraAZH8MEEnHkMfar3UxjXCYSuEAL1XIJTCEjistdZ2MvjSinX2zn+Km
+eGZ71N5W54xTA0QjAw3Q8CWhvDF9g9orbF9IrgCSa6sJoBAAG6sI8M/aJK1MS9I
ycXLlAqcJhuX2Wm/avBzeqPHLw/otlWDjuCjL9tOm22Xy/pQyj53dO0mtwXyskuW
Aq6hegRIYMIIY5j+bxbMhJfQ+sPrBcK7OBWVXeZ8fioxH6jEFtfB1TC1+DiDmQog
wqMKPhinu/+22QRgPczFGYkssg7Im77oZRzcKZH3v5EY1cf23UZY8ffFc0c1tmfH
Ue6ZstImtgKxih31yXsiGgbANgX1mn/aVN8s0jeGhfJVzdgp0oPjAIYN1bmDoj5S
Qba6lriWJfWj71d7plrLFa7q3JM3WV6PDl6Ezl8jz3WQuMVTNmPiOveTZupud1dU
5aD9S2x9qpJ+MEUxMN0kumbQGVW8PQ2P6rYmsW7ou8qCSbwdAbW9PsRf5VTb8eJ3
qgpx5lKbvNfaYIhQsGec1PH9ObQ9JiPxvbkodOSA91ITdtkCa1owoBEWaMvs49sV
lU/oa6d2Pnk/vBkZwPDQ8rXeG+jxxCx/eNFibphs0EvI/WQWt7xjyHmdPeVR0xY7
9/XSK+svMb2e5jLuqss/y1poXvGdqHkoxdHnAR9AFtFcr3Jws7vP3STKtZAZyG2f
Uras3kfKZBjYGJWEy6G/EwKL6sX45kgCBHtkk+LpDwk8Q/2Z+mh7CqOv3PEUtYeS
i0u5v6WBTO8WikXbTgigfrrP7XxwUIJDgw3g7zeta/4IqcdFqExiEPg2H7hIJ6W5
yW0NJc67ZLOy+LNDkV/JrWITiKVOWvVWJwszRxC6V0D4xKzwRWQxfTJdD8SLtA4j
Iua1MzuX643QEL61YOZpqZ9eJJcY+0HvrKszEigtfl/LRGDvlTL9K4xBbU2XzDyX
zhNQGGpPiNPGI0BZqx2fBXzW82wvBzYw1YvoFFYLQx14k3BfZPriTFEeGvU56tAV
zFRiNHb+no0xrkYdXvCrv5jMHB2PDnv2XbAunBGeAfAGOKMfsiPwzw879teNGV9e
h/p25xBxWvUbFrxNyGh3JnwU3w5pH/R2Jd+PSE6mwVDRBHz/H5faYtEYakAk3QMh
YT274DWwRzlj0ps0VXKpE6Yr8RqsMH1CbsubZAHPlbNsQuwA1qpdQEq/0SbVKvjh
o7l+/l9OgTsdotd067YkmXkcyHNInhnOWcaO2yt/J66RO4LYzStj/Nx3q/otFffb
qPDmV6zOiPjb9MnnB2Fx/3sLvXO0bvuxEq2Ib17Ma8b3YDLFoE25XcNTBbsV5qrO
74jdQkDaEjh7za28CIcvgfDpMYf/IbqFk5sax7Q/SuZgfkJkO3H1b7M9F/68XUrt
sfJro2Q13z1IXcVbVqx7ovA63HEIK3j92ThMAhADcWTgalp5YP4O4zrxOxHX3h6n
Xf+S6sBpXpXiwv32WMxSEnWlW7ReA9RgmdOkfxfgxCtty58uJLvL4CWuoSMyBSj1
iDq8l4wlECAWdp6J6DFKZZRw/6xKjNVMKHeOMNndrFmeMlKuNp2sIwk6uHWDQbnR
Hqaun2XeOoJlAuj4ItV3GNzGQIgW5rW7MJ2Bz4ALfjZiqjHnGAmOqyYNNHdROZxe
EbPM6kY9/NTWa+VvOBVGdoZZs3znensprF2pTMKgjP2pNSczFNjyQ3iGcQI+g//e
fAFkDrqYLIa6++SrSbF8Ym1svJyb/DuLtf0Do1X3lzR8Ks4HEXXWTK1wMl0iSj9G
9OVJkLXnxveKLPbAY4fZV2nq6xJMlGYPxQ/JQmGs0jROx9mYM1g5fV9/K9xmDQ9K
gKcUO4+mAUuaSGtAEjYCsArBp9CBD3Yn/yDhpmwEKWs6zKWz86fp453lEi71jmD3
QCX/RkKLRAbU5Ir5ty9opmyMfagWVuuJqogeho/ioaIAqAUOb8z/h5U3KDm8LDqU
PV9mcWfoXoxOlLoReoutinTgNhI39k8v+Q6em+N+0mESDHnwCd0/1Wddnavid6QJ
HwoCSPIYlxDa2qyQL0JXoUtPkJgfUunRrovj/ddGeBgequMbaFf96BlJxOEugZLq
d8+GTEZzIUpud0fLYjjY5unViyhaKzsUWLfZL47mOQbcvntVr9qOCJXBGZi7m+zM
Wz6UKjBW25PbAG4iJ2EXSDJ/lESyApolCyV01e0Jb+qBoPFke4qor9NQ+DuVXlUh
43pHEY6DjKUVlnAn6vJdzrQT/GxOvbz69jn/WRwqHOR0Jpjzn86rVJco90TQheyP
VEqKPQpt6CRF6FP57x6qqYqS+y5BPXIPYmT4awm3LZkC9qXr6AFT6ADj3QzzwWaf
zJ72x6tscNsqcHUnQc+u3MMIZuHvAS0xQ0bNuhJdgoPbGU+1kMK3rN1pRhimyigc
yIeIWXVfKLgHLYwmpXFvZr8wGYKu40g2+sUySRvdGWiV0M6YtauKg7Lz9ihLFZ5H
4JZ8gZwWgTQH80cn+3BBzpgMRcvtrnox5EwIKEKydEnv7bkyu+4NMdPCrgA4q0TS
IQxsBtfpIc+9MTDSydQ9tBk4MFK1lkuU37C0JAVGtAXiYWfxO0wtHJUy94QEie17
rAvCzibZD2UMog2PctRiZTKAB8eMrGdPMiATbHo/Yve0+aEWLsmsHWeufxvBXNC+
j4VyXC2wfv7tDtcGUkG/wBGqMGrcdJigEwDrfPQfpvAj+7ScUSZuLEExDBDKSwuW
9ibsnmRrldg2OXEDQ/lPHoD+dHxCUylb2HdocFwpRX4DVUG50Jb5+LrFhWktsB9W
5Ge82kjrJfnxMfUbx/c/3toKyAmTu4HKuvjMoX6R4zKIZ9HqbX87yQ7/1COHN6SH
uBr+hZqcgUgXYiyItbayfGgHsKU0RlgAf7wfgpLcR5KSva1IspAABN53AS5gw6S5
ZWy7mo2wXrFLq7QnlMmeFz7jDDy98/c4lXoXewhLXaMJ/VVfl48b5qfw2H7JC/uC
Onv+HoUVNFVCaeSICwEI3uWgvc1csV+9viyYqcxzQuvl4xQtWqvGCKvwlMUW7qS6
bkd8dQYp/Sy5U3kWf/7E/3qvdDhbq8yRTeBv5aDaLyWuU4RidYT6pSFTRANjWvma
Ij4JK5Y6hXkqvNqkxe94vY7EyCl2FEsRl3uCBl9IPXo4c8AIGDHN86HWQwOJyhFI
bD+HgLih3TbGLDI1C+6WtDJ30zPFnZfQtizfQQ7cmzF4ggkf0itcWRaj7EC5J3+G
TYpMJrbBe8pBBSR5bJsxghSgFA15mdzatjDB6RfyPkwc8RoWUi0mG8WTn/DAwRJo
gX4vh5zPx7u5vPI9pHW2ih6KlvU68sMW+O5ojKt7AwsEW+rZvTy6NvNjER5DnsRw
rZvZyqZ5qrFMACgdHKJixb1eZbsOQusfok6Tv/CZeD6aFVUJtdWqOTxuz5ff8J8r
31OhKx+KYvGwLdEYEXJ5HAMj4JDvzpPuerlAW5R14ufTERFppB5YSqA0heWsTSZm
AgfePE6/6qCPcU3N42dGJ6mCA2p3W9wURoTWubCaX0q6uAkkDBICtyiinmwQsVtY
DGnpDStSfb8bq9wynxC5jwn4Hh2Anez75DchOHQ32arGcC1p6fAXKaqzNuorQ6jK
yBvSo10kwv1wCyIUbQsgLIc/dplVOnbgn6b4Mu0BVw7nS2ZhkTxM5u9HkCb7gk/8
XEyGkCm41Ik9IzUSsYODWeQDn4lPJ8FeahNEjL066R2TFAmtHHgvweLxNqkyuRGZ
iZtIu8A6TUJucjE1scl5EI9Iaoz7OZ35l5qnvvMjcaCTF6ckqFAw8GlCeF5Nog4P
FjVtFNkOw21ehXWKvGA3SRw1fIldvFVtmU1NoyAcaLQ7KlSsjYCHcoYaCfE+cvM7
/ew8yANlysplY6PL0YZ3zIsZknrxWFqtFK7VXF8kewFR1L1cfntu2y4PvBDqvk/W
bdtDQ+n1k4UjnfhSI+Y/JxC28bvJwCYoJXv7WlTZTdv3ONhV1+H/iZBZerTNYyut
rpv1oAftUzTvJD2JuVYMaO/nS0GV71mUVqpmXZtak97DTzA39b+TTpBvHM0F9tbm
Un1Kl8SH3bGOHQyInhtAKKuWBX6IcS2IHJsC1fCwsW5/N1xtJxowh1/k0gXxOyGs
nnieEwwviDmgJfYrl/Y8NXuF+OfQr0ILLFJwGelLvEGExl25FxiE8JPH/V299qeT
YhevdIGE6kwj8RyF4/fx9ma66ObYgTwqaWwgPIaGI7AzC5UFcHfuZnHpsxuDLfYJ
RE7GswN9+adRAilo4vIqa6O47mLE64CQX2oWeVrsRYIyagZZ4aa/DLVzEqrU/fd9
6Y6mDahfZmtuHbYh3/LPWLZ/is98RRWzgNVK1QTLkBIkyZyt9AdMX70WLO4tdgpX
HIbIGQunY6/IKJvFqx0k158/kNlLZEQ2SyZbHu16AlZM/Tcjh7ObktSoNtCijPxe
HL/QL0x8r+BEFG6YIxScHu2mjysQRyrMQJW8zUvorNr9G6Er5SJ8M5q1iYLX7aRT
OyALwxxw9N0IPSVlsdY+apwg4f++y3OOWp2YhtL76Jp04d4DPNMsT9VWCBUMgGGP
gRiGtbtmGCXhuYBBvebB7LHTMotZvHpqLeHP4mBYCrbfi246ao3DyPWyLZ5PCw8M
JNGorg5QR9t6hOxNyoeXmZJqJyLUoSE48Lja0EBjKN29wR2kl1ouHyfScB33MSWH
4aqqR0VesruXD7yiXS0xsDmKom96ocSSlYppJgswtMBeH608ojtUlMLaZw8f7C33
ltNwVoLt3JEIUAQIQW5RoQh3lTh11x2jNlIjzcmqbu2Emby0MkP4EZ7OpS7it+3/
v6oLy9oGfkD9AIcNrrY/ki+LIM/322aX4ySGXIEdfd/XbJUsghMGijoPBezdNNmw
ctxRqr1Ez8j0rl3Wld39psKqHw3IFuUwb1f9pofLjS9WaQVdPtgLXNlpC1afO/yk
fHJLIHT30yjKJkIdRwOjf5IJrApU7hS4sJBaVQ9avN5n2DTicJZf9jAB04A3DMlW
dmSyUosev7fsxlI2ZfBPdtw5SESGjSX+sr9fibeFzW1TGPTN1YJ2CNozAyM7rtyF
ttPfYus9yhWkxsUl3fvthIO/IYACcKkTT4DmqBZySJpe7no0oqhgogOCVXII2ciO
ktfUvV2Qr4Gf9yeEZlfTtqHLtZkTccG5+qV1g9+2VwmrH9HOcc46zrTwBXE0FUZG
c7lw1rNYM7OhdmGMBvNbXW02zhz1j6/vY1QyKdXX3irioR4XutE4G2n92V2zxGnN
MyqCAP1uU9qyJFN21wKq0VZfXOaogYE+BkgW8zlrcCHyi/nLm4hpP1ZUK9/S97xN
9UWtI8Kmj99WynFzypNCJguxicJ5Kj6wM3080s4tq1L9vY8wLqsvEj2ZC5sfIUop
827OqN34sLmPNctEIBbGuQRrfqruCr6DstvtrsHUxZ/LNs6J2BHeod9XAnS1BLJQ
d/62W0wcI+qehDFne2svs25kbqtBuQ19KSevf2yrP/aymoy49yRuDU0nI7KvNulQ
3ibRt8MBaWbljEZ1ARYPB1nis85YGAl9R7+2+xou72mfxfzyyJZLHTHISqtPb+G/
4yYm5N4CIdc7iMg952lgTWRfGVqYONbTwuqM51mm9cHSZyt5F3x6FeCb5jiEffRq
OupjDHTNLcs7llgzKEZPPYWQfkaSUfmSX/xUKONctkrkdtgGr/poGydLy2XR5A/R
cn6BcS0kAd13GYg7+dnAcZ9UqnIQHnJxiunZjE/X+QF7lSaRO6+nO1qvef7rs8aW
xRBAAXHhQDclq4F+5ck+lmA3WmqE9XF0VcbAv16t4AYORQZBXmyIZbY81f1tQZz8
3LT+zLyq0b/CjiOOMWFEfQPTlazqqff42emdANM3anT3+DoZXITZ4ddc9WqXpPcG
bAdmEKMWTuugZwHJWXPqysqCEFI9OjHfhlYfqI+B10vsmC9GCAmeIJQe86GF5B1J
qbgub5ouNkTyHuUW6jy5QgaLmHO3sbZUcUTfRmtfhV0qVnCM9bQVFg6mq/81QyRW
OA3jLAOfvaS1VJ+4w9cgDIIDKuTnVaBJLB+ma554kY3Z/B7BFuHROSfmplq5MFkk
whs9FIEDE9NvDMEbK8LASOnoDCbW7PgSLWNNhVVKODsLNJoFyvRwsuaG4iOz5oWP
aRVtIc6PWLfBth28cEDIU6TNdll3RHO8AXIUu6vbX5aeCag+vgjsbAGm+4PxWzB8
+jSEdF+0LpaaQFC8V2iRnsyy8H3y86vQNEElGucwaDLqCvN3oaFiUomaOgaft8Zw
1LYdxV1jEml07hW17tEnPJEtufhcwSq6L63NwexaAu06PrfdQ/m3HyqDZN2oLK7y
eR/GXbVqEZBJ3nvphLPEBjQLaxkGX0AjCeSi2FZbM6KJc8YLr5Y56RWzr8WPyOoC
ZMw8TRlRhnIdssoMD2IqcF31CqJukksUXLIXBdyBUHBMdPnHwKUzrGsI9AxT3rwG
2gF/aci51Zy5/mTrSSUWRxGgajQU0OYb+eqkMli6YK7dAweSpJ15inXsP39tUt37
O8I99tQQ+kH+swgSErSosBQfsoIlBqq9u/joHCNF2erq8Vi1VPVLH/7PnRQpCCV8
IZxhznxPRK6IzihnmkBr1zlEuNORAMK6AC9NUW0Y8i3prA30aVePFEyeyZvOaxJm
cxj7Gh1Oc6R7Oc8TAap96GGf0Ubk+E3LRhRuJH1Ty4S/5sTPzS1Dk1uyZMJZimll
HMhZgmubDaEyURrC3/nCInLRMg7JQjPvXH2jNs9r9EjVRbulgdGL3ZoNlRxguOp8
z0v6Kf5JG4aO8YPCnB4P8YoRwWPOtGOdj4wZYX7TNhUS23BxSH5dX/egU5iym8qV
/NqtDkxlob0ExfOdHOE0n/RdmkVS182y5BZdF+F5ooH0OghKADwfC0U6+85YIEBH
Zh+LlrCzDWEC05B+zGEJqDkzC8WzIKX/zKeFd7OnNrxKVHVElHHPMgYtvDEXUUHQ
u57XqSj/rXNuDZFgREP+Hgn5PvkWDK9FBJjxmzzmiobWyyh1riY/FxbhpQ/AHFlF
yu3rnYdEcpjNk7Ouqwe9m89Tl275BBFLMk9bIyjW4eB6Gfm114CziFNjFeb2gV7n
apWXddVX4qu1xWxmdR03ngx6MtsbiCW2YtQyP8ZTXmAZgOcZiUuKogkT0mNMGC17
Hf7f3obGAK8+UpRY0gT+owToR2KjSZ+YbiS9sgY4lqe4PgWJcXTT12QPazspmQEG
PRfVATYk48HpojX7SM3IM7YTZnW6sqx2o5XTRmrGddfWYjkqMNdfJTFg0Ovwe3Sm
EETp87UXqZ+m0uJV1DroK+GDEkB3wT1AIuMm1RN1cRnYYD8yUksmfGCKCBdG+KVF
Mn4mOn1CE1nLqSV796kdaEkdx/n7y8jEYgB0JBoR2knvY0xFikpXFLJzMSJgA33Y
Y2KRNrO1u71Eu/NecKAeJJhcb0ZsFFQV1vTzMCRsrpzPzYijCMe4kAFz3fZFZLDd
RsT5fnfqeByetq0GVS95cqJg87yxGzbLE1HQRK0ErsjRBuRx1spyY8SMebuQSU2H
DsYzzCjFsNsuxMgUq5ZfmJbOesu76jyEc56fjEg1kUpELPB90ZTtm61Oy2OA7YTI
ISqwFXHswsB1VU2OE0DA1IZ5SIJ5m9XbkqX+FTc1rMrktBu+EYAvAlw1vEKetGy4
4Y0x7RKfiuqJ5ZNGIDcNLUelQ3Ud8PG083zTB4OFRLQA/X558CRLflRxve51CSJ8
N8dnesgyM3TsphZPT0kI6qMB1evsymUGmgV0kHIMNFJv6FMqDLnZeoRHRJ/xmWL6
5JESqTJT05/LVRY3GrB46Tvq3K/6ivc1XFlyMcq73pKNGKXW7Z+1b5Tt5qH/qztZ
uxfdEzqv4UL9CMEiwTZ5zAhs5+Hn7J2Mroe4VMS1pcUjox/yZwKoZSbmTwPCTWfY
7IO0MrJq7XCkq7qeN8/4NWFqY0+GN5ueDqlum57c3HzHvNuh5gvr00SqnbX4sJcM
CkICQz1ow8uGlmVYlq6eL0JwrbSieKfR2a0jjhP80ypcE/K3SbsdcNaIy1ifUYRI
/yOtg88mNIoEWXuJmejcN6QOLDIk40iM/9Zl2cowKqOKzm1cHLN7KgCMf6PuaLat
CPXVCyX7tSpwSQ7cQdQwKvpcab+q4zY5j7cdXyYHtpFrCideILNLXj521Q68cyjv
pkFLvK2IHvTzno0k48BVm0201AZiscdjmjxWamlc4HvVn9XXo7kCCbAKmTJaB82E
/Ja3CaE5rIDKwsMQcnFK5vx7pCMrCbR1w2VrtLhSSLQWCB7hgqv5680TFto8/iBy
8osZdR4LKZALhEzYzAggw9IeO1pj4VsZy6JVI6jz3htzG1yEd39NMoWNH2CkCART
HzPk7dcDbsL1yWcnndkyg7Wn69IqG/caWlhbolFdUMhV3eOgNOPTI0QEzN63uVZY
nbj0SqxleQtWNNjtUpinm8gOorKAMCdlRE+rcaY2XddHYnwJgjhQaHO5zDdoe6Xh
MaipNQJjuxoAJksYViSXUNTvsbR+0eovv1qRJ3RXtREVGeTn+5buhmh2gwmwgQeL
BbGoWZH5RcGdQIOTxv24ITHPGR0ZgDY/5V1VtKwyITrj5/Gpoy4NZFBcFnpwOvji
Hg4KC4qCoQBNgK2XcZB+9wto2MNV47NeM5idp4eht6INGU2N/+AI7F72zVkSfV1n
W8m9RkcyLVat/tUTLLHsxtSRBWFCyH5zwgnScHofjRlrmAV5lO8mJHsa12eEji5h
D1iIxcbeopzPFt2hnbYj9HSfkfP2w0SIQ6idqmvJ0IxPWvoHKDwxhiMD/kFe08ei
8+Lmpc9od25rueM4TnWigwSV0ptiUgt7APYfKmZbjVgRclYGyiFjAmaNd0PTyQgm
gP0KMmiQbbU/ya71mg8OJqBBvJXiEptnAxTYjiTKq0R9Z9VV+FnYz48iTWXUVQ3s
30Znt0jQ1455LG5+cT/a2O16JyJfqaJQSJc6Rn0LYulIBRmlp64atWLkasDKjWMf
TOrv7lfnpIHjxRWqG6HtGF8N0Q/3H+CRmM9g03GMQxzlyjrR2fFMTzmn5OaW2iWw
9EGDw6dtqst4qiZUxU2JptulSXsI0BE+N9I4KqF9etsVR931sptwu52bVHn8W4EY
mSQoF8zWrj8i4O5RXCANJrMh0TM/2zNSRXPBsQOIujNCBgOQTqduhs+GkPvX2BMx
0D6YadZ70hS4kfq73GugJwyTYyinqH085yo/txSYz7wZA4FZ8VZrjsvCHP2mz1Gn
WGGdSl2HHi78R7B6G2z9C04rGnx71SN9bTKIWB/IUuPYBqivmJjaQ56UoFpNni5M
2lSCnmFb3fJ1VrmM1FixR1COLXjp+QYivUrWWS+c/XqKKdssiH8oBZvktCNeqUAY
iANnnje0S+UxMND05Oy92XSoTshwNi/fyJdTcb03H1HdzmTrA4R3My9esRWghmlE
h0V0kwrvKb696QFbXWmlCc3gUwv/iztszfBqfxMieLt38/kGAW/jr5232iC8P8E8
0kKAUanfNmp08I6L1klBl+P5jD0mRTKF/FPHIwYk6uLL7968de7g0IBzHTCjhJp+
jLGN59Tv43qnstHAVfmu2SgMKRLByVYq7cZE89oXOlw9S5P17E0sXSUV4GaOhZFr
GtJblXnxgRLC4VzzPqpi3JaEtFah1hCpnwsIFL7iYnI0hInTFR3elYLZjo1RyxTS
cKUbjB8NuJBiisd1ioo2X+CADbkB3EFYwjKlZCqkWtYenhLPSjQS1KnvMXjkKquK
fB75f7vzRiuw0BPTDrleQPIgrQZ2s51FgUfWQnh+ovXuaombmCljU8KLtXporcQE
WKwmUuWs/EfzP4Gf+nlGM15MzVWE0kA54FzshdUifKCMyJzWvwVXzZRqPlivXJ+R
MRHod1j6tx9nPazn+i3SqgDxcNGSTG7SneA542dZavZpHMYDx8bxXnLfDDo9Hiyd
Q89TmjhKEX4xZ4EuIOl7cMly+XkA6+vqCdWllbfoY7JzUBlHof+K/zBUDaxkrAt2
o+Hi3417nIhFaXeTW0LmO6/4/ItnOTYHsDwwM+eWuXdQLYdBJjfqn+Gb1Ycwe2PY
YGS2tSakTxpHxZdOvEHZVHg0kZpUCT6tuMp6LMxmSgp1rVf/84F9fzlrM606f1AF
eJA1SFqcgqdUChX8onCbMXOmOy29byv4EbNrfq5RMXHXbEcTNA3cWuq5nb5PntUI
k/YNTrqJZjqunrhey9osTXayC5TBxiIcsgB3TathssQVmis/XHBEfK5G1Bv1yEVb
wJclV6wP0UZZEjCAgcBZSz3S0M4+SpD7rLEbJZA40GwdRMn/ICIRCWtrOet+NItN
ev4kdVdxfyACFn3M4BZPIWBCkTqTcfS7gJ+0M8QBNW8Y/yCNpRBZLWfa2xbggpd5
eHG0x+2NmrcSictIyCzBNLsvEHn/M/5CQG3Q02UbBUy2eR6reCpC/0MsZqM37VU4
Keu8t2gBPnZfeRwuCGSE4/JYmUhom8vOCEzqD9siPjhZVxv1rwih1NkZvLzYaeV/
cJxjJA5o5ztabWiAYCMle+m8RhxJy7GelMbD0b+UCCFix6dI06UDXHhEb4Y6o+LV
j/LQXTz7LkZK7yj0muYI94+dgl7Y1vc5ytLbXIkLEGl+3WV5gTmAJQx5OdQEeWod
E+3itTOTlGMvkNzzO+2qxsFNyBC42kLbH9Z+F0Wvmoc/t0mSxJ6GOX14+l/dSgpa
LrukwS/Gp4PAVFiZZ1JkuBJECUEJU6bMXwHxXi5Q4ttVsn8XfMSAqsyRW/ej44Se
9j56chTdZa13HCIObdTznsV8BrvnmKJCsumJEt4Hz1rTZ/Vy9llisLVaxMBIx5zW
XBmbTFFrwk6lckR7qQYCL2PiuOSNB0VqQ90DHSfS79x1IJXyo/i2dwbc9E7fdUU6
b0LNKVwlDtbERCOXm8r+DuvPIT+Yx17xyhYP1wqwbMWjZXdKNKcfBMMPWQkNkI2a
6gUnHu4NMaB/foWU39768Jq78xHNkinIMpMcbplheVxQISftIUASizW53i9p53f9
qHZGmbTrPcMe0Ky4DLfV09tn6Yu45RL5nRcE13t+4W6i6y/4/XnTpWLAZPMDnom2
nB0wftAUWqs9HmqNSJZt/49jqs2Sbqr83Zwa41yDkLsNet8OGTVTuPWQ2c3mCDPI
o6Tis46T6hEkUjAX5LcnvgITxqhnS/UAwlp5Z+pe6m1Yxrm3KSx+k6MVq6WgNOES
riCo2EDJzk5/fj4fA9t5k5n+fTWqsp78ZZ8eDnv+Y43ptSiPSmrnjQiRCzv7xwTR
uLxRsciZLjB+AUT6ogf6LTa0bvXJ/BgdPSe7hYdIkYzVns+lyslkNHIPkV2Sas79
tQEDh6VVNjHe0Pkl+e6jl08GoRhUZJQQVWUKlVpPI9Zvhkon/sMI4v6YOFq2Z89f
FCVaqXcqFgFwODVB3qTKTpr+FZY9PPWmL2ooeCdTNVG6SASCxBIH/GCirOkZBIHz
cRifpbPEvIfAG9YOsY+A/Ilnvlck+CwNf3+x2231BF6xfXJ0MSxZ5n0V/4W7yBrW
MIoKK/hJazDkYKcHDinA1AU6D33Pd6ORGkm74etg3R6+nbN4DkPqFdqKeJ1VJBbM
YrBMkXlKdWIA035t7HrkAe9mPj/F6w7yz8PRFThKK1/JVwL4ei7Ks5I+H1BYhKqP
KKE5jwp4CJa3hS+i9GvTiYWrP7VliihJO9DBaAXm7SczcSBfqK6ubUKpagDaPfzk
zSXXcH318EfUI2Wseld4UwrX039u7y2d9b9Y4yuJxrZBkSrJtIqMAxMVEtW+97Kn
wQjJENm6faLw1AhY61Vo5RbJJ5ppjeV2Ab3u7xhv5ytjkF6/UenWqV8y8eOl7cbJ
oaeneiewBu+CFs5iggBUhcbnVJ3UDaLbmGO8OuHYiSaUA+BWnliuP63HxUCjXcyL
7D8RJg3ZpIM8VTDrEu8AT2C0y6s1eyNK1kgr/gmFXLzg7FfmiASpTO9Zn7bFIFIF
L3L0y2dId370nR3iANLm4S69IFqvLK5kJIEb5dBQAbcaFtpVHlfZpsBQ79CITttG
jKRzFfh8We0NiwS939MfvSDXF8a3GPIuoXB0SJZsEbpqcy/7GfGUTxDxukJr5O+m
PjsP50isQfo02XHs3a1QUIvc9x4ul+rIIdrIYF96X/W4CnlNxAAlxLjfTIIOn/4F
uveK0+l+tKjjIuK57JCO4MDha8vFaMh7RFV3nCbRfPTTf1HcZOlQifoZW1IAd6+L
soUH8ZCuExFL7OmgxQm/qaFzPcQzUYlvr+zNXYzoOvTtHssbna1LNH99KmYDftNq
OkXYGhZznqdSAKXt8GLOMROycWSParny10tr5SFtP1W3Ma23xgzuFydm8G+QsrRE
k/gJD1CudJaaQQE3XJldUH5paFsnHw/K1gIJ6WC6r34RhRhKlhRPXJWFjs0X6uVr
VzMjmBAuB9xmwE7aw69rSAxll3RigZrWcs4pSOJeGlSRmQYHsat1v3uQoTEI4RKS
ZqbtkcJWL2zk3O2qNJkN/Rn5zBSHPKsrIGQ868jCWKxZHXD1dHxbJMFqwDJnd475
1AgucrWxSzhdZ/InPypDLlHcKfL63HdjFyBWF9gkdI3K6zeber35XOlNrcnCSG3R
TO9Il0jAdpG+7lz8vtdyEG68KXWoXW1nDS7qwbngXCUv7IMBW0p0xYOzTY1Qzad7
gzsxs2u3Uz3O/ScmpO/IWrTOhgDwCU4Kt0bbs6qtDcYE+R5/vai0/8IAOUri1+tx
CzYYTzSe3Vnx0TntJYuCkuMdOzGWHEi8yHzi7MrvBLFHodZjSOyrMRhnfGrPofoe
GRvmYMInDGAfBlMcaOx4baWezkE17n6/sZ6aqyGBh0BTD0/vN6DCAXEvM6j3mUy6
Xn0avEc1IwHJPgakkb/M4LsCg1eYnagvnRs5E9IRWhsWEIUYNdBk3M4/494eXSiV
2AyAspkPHDOvqo6TCHDrSdJ8VRnmdL71dY4IHDvl+JDuDojrKxYyMo6SgeacBk4B
uKs/AXK0CozzgbrMeBpNQoP63cle8qj8lJTOeRM3d8jcNg3r5dAOWD6MO5AdVp+6
DSiN5nQ5mBnQRWN3xylaJAkAXYNadJJnWsK/m/wymHL4efghHtbtzyv17QpGu2RX
kUuI9V62S5OkeZhHiRJe7fBB9d+tKr2Zt8OBvJA8plNzxQGeWHYREi1vopm7TnW1
3cuCogzUFp8bDyQCvnr9sW7DVkQfFpGGw+IVJu2IjJDImy1Jxu3xZhJDqkvsmgfj
rbmqFNrSb79K8/8B4vDtFnw0yHUfjp2IivwfxzB2DFrNIxzjxN7VDM99XUh4VWjZ
bjDr6Mg51Mpn2bPk5hSnrsnwOa4eK8CU2DSKXb6xd7JsT4UWXwuFQMAHe8gJUXQZ
HDuSAye+sAHu1r27hn+aqXQ4j9UETag+WDhJfbZ7qmhrYBtMiYIMc/9KCM7c4Kbt
pJEJtj/JYoVMw2fzfQuKV26aNqB4E65zHYr8YxLVACbJA2k9WKSfhdyJSSFxjmhI
iuqTVhcFbMqW2XYZ8aRTJpVieywIPZajkNTXoLW5GBVLxB/vOV0LUx032RzzZTI0
HlxUucAUahk6mjuCJKn6Q+89ZW9RJYinPG8AE3ucH9EZ662l12xQjEEVrcaeCzPx
IXSg/QHfQ2Ua03+Uj+7n1YUPGH+JidLniR+Q8GhKzypO+xtdIzvksGfkPrFHtpOD
V32DeJaYv/cd14xiI97DT6cjxKksJfFx8zg4IZarqP1pxgeNpTDUDEBBXHMVMjcO
0mtE5hCD5YEczzG15ll+v1vYCEZ97+5Q+djP2OAF9LEY92nSFbLkwoJDbbt+iTyL
ydVJ4v/wmDETWRKr8Zt+5Q==
`protect END_PROTECTED
