`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ggIXSyEavbBar1XrPnNvUcW5//Lmv5yLNXPRCTmQEn0Le2AhStChQ4LUkJFUcst0
E9r392mMybSrGvKPtYN+bbqSlUbLxlPNYfnGFuRrDe1eua9pLq7oLn06ocFtuszC
hb775572hFaKnnC1zcBiJ1d4GEG31d7OtdubvVMFuJIXCmZi6BPluErexnTSD81r
O3RJZ4831k/fqnN21BW6PcM8Npq1kfeIiIAh3CvHheWP0h39UKxPszw+8FGUsMCd
DuapxnsDQbg6NaIlGSv987PUpRbLG4/widIG17x6pt+Xwivm8AsqPJZ7Fotq6TWs
HLiG19Q3DZ5+GeitcCQ+G8zOwY4y7e9wrPj5m5A3aP1FodNE2M6YPLBnz1PvhPqP
MxP8W4QAW0NB8ZWOPgb2uqD+Y0r24uJhQiXAiEm34XfCdkWybddvzGw69mosBXuN
ed1/odsul9s+P351bQFWkK7DXrLHuFHoTsTma6KnjjAsrXG1G8pr0NGjr9/DWo7K
unRq5pkZEWMKGSzByw74Hy1oN3Vr9/WK7neAOCFMZLxdVmH9OtjaEW9C3b16IqfP
wzeO7z2KG9+xIHZFOeC5tBDaLHlx/L+7sNj0gx+UmUSs1MOyUFTbrwPiP4BNCz69
vvzT9+tGSlvqsJ79Qp0IaC8NwY38DAGJBnCVrZ9jchPc391/UJEoRo266wUQKtfB
DBeEx/D+TcUzoaHpXiJgK6K4FMYhnVjc5wJb6S20+82hYrbJFA+x3unnN+Ix2KDd
+33aYdIfutoSfrIHx51Vh8Ahk/xw9ri66CHWKBQdCWXcCgeREw2bWbNfJvaILIIV
vqybbxIxGuUlxBz2BBcdcUFKOG2aVocm4rW5Op6EasjHGqw3CkJ/Wm4YjcFV83gV
WArglZ6kF1ZVKmGYMVHnI4K56KG7s3ig4axRraQqe5HEQcAnblKHV8ZYfJI0OR68
HNpF8ZVQ43PS1//3ebBJeCWrjXFigsLj2hoyNB2Q8y25yo/YMftSUSabdyNFGRyT
jnxa/TbMYcpFWltiq+oOwKw3l4Eo4gh/Wuxyvj4J/H0Feevkcwswdp4cvZ1vpxlU
1OD102d35MQKhGUQlw6a8PyzEl1tjBy1180yfvoUgCJPzuEvMaKy/K7IDdLTV0rV
kud1tnZTX17qfUfBJhD0R0T/QcMcsiJdgCUMp/deyliv69shHAy78GxC0OiGZRgc
1spY6oslYp8f1ePPXP7eWvy89gD4UjlM1u06z9xgz42O6Ccs8R63Nn+dlh50oSts
VMMEWBUCo9vuuwh4ap7UmI4GZh5jd6gG+9E6E3uuSUywyTBSXCj5VFaTVBEnftOU
xaUNT6lyDK5t/7YG61LOHSlxvopwGqAXXMDlALuh793HwmxSvzreCcGCsUY6sd/I
NSMdxDSXbvAO6RBleaprmw8EaJWoxHBVVIrHnyUkLoryrgiUJlYLIpfu7tk8x0+O
88ObA97lhEPzWWqYFoH9nHimWnkgAvTmHxOlZFHlDcxtZDqvj2ah/8EQNJX1NVpO
+t6ai9A4h07m1sifN3sM5mSv3I5e8SYCB4SOfW7EhCLav/C/pAhLSGwm0uEkkFwQ
9XBAEAqL/FfbHwrHuHGvs023u/ZmmErcG2v4N4RGbGwj9YC0MbrzghiODInSE8cH
CBVM8Tdoey2kOrUAhfbpMfG06an5Ojkg5elWQyCGuX82go21PXbMSQJ7xRDudMW9
iPhh0ZmkfCjqPfL3vYSkDQlmkc34oxh9iU9xL4ItnUJZAniL02B7br3GpH1DCCrE
fCsAwfSSCHeWQpnXEq2y19CRlT+U8h/ymWo9WPDVxAxD677DmSnlwO3H02casrbL
q0Iw04vn3BMxiem+p25P/gR8lS2nNdpZAScwMiSXh+YUqCUK8wAQyRLvjHTXzyLS
upbrRQS4Sd74N887h0nXKG3suBVU3rr/NRZTIrIGq20gj49rVvd5rXZsdIHoQ2jn
OrrpU+HfU88tjPTA5vANZ5u5ih6oaY1+idUwEziKGOaMhjM/MblNQSgmpJ8rZV8u
reDsmVeq41QhBX3czTNfEsOcxSmsliP2AbGaNZLS+0Kkft/tq6r9XxUvyZGv84fM
swQCqQ8o9uGJPSDafFC1lXpK0wglPVy34EMe6tRaVRa5TOnSH2tKjH1BKr04HJgx
T+WL8GjbUiDiHXpT8UbkpjdBq6TC1SGS+sa3bCPM2zgICX2yqIefiDsBxXBgmmgS
VQTUuAPSmvFZBavBJKkEmDkiWohvz3pIaBYhEiawi9RKyqlT3UK/Xw9H7qvhIJbl
BqBerWMKf0LTqWeRxKYt3r/kpk4sofrjuq16FayT2/FgpM9LVux0NHmQYkjEdZ4m
5r/9Qj/o/oFmZwaoKPzADw7bzC1hcrFZsN8t9qb3FOP9Nzobllf89vXulB/SRKww
Y5vDrH/XrJ54GdwDDvlg9BuvybDTuYtQ0L3fpDGb4Z/YeWviRBYtzVmJ3v/CZ5Nh
s2IxYUg8mCrmFO+TDHl1QdIEPHUucYxwRmZDpDmdEtCONnNXX9s4Yb+k24xgb1qi
SP5Y7tr/MUzPBZ9asGj2oQPkUXBGwA5oT/PLilX1R6/xu8E7eQbTdDbKIVsR4HhK
FIfvKV7Jfp4fiiWArrynK6byyh2QtWXStcpcpiGxg72W7tfIidNkQVav3BwMccH8
LAAGVTiV3c4Y4ewmZ2snCwtdjYf1p43xzFdZF7A7ZV44044dea+VkHizR5XGVkZH
4mbURr6LKOZiBesNxlMI6YAA/ZbSx4HfZF/1XV+RmNe1fN749t+xt/chMMMYsoVB
3det0EeF5E3MNvS7PQJz83TJjqh052aLt20DCTyRUUi4IflvvrrO6s5H8UoJmmCV
mknjl1tiwVOrmHiIB6JX95Ds60dpU3HY1TngR+qwDVZrth/iwVI9wXvTOSZPZgIT
TpaKDaUkQI/wBZViin/jVWW7da2SENMr0RWE235s553KdvOuYUU8p+CghePQDlNv
06gEn6/OfvzRi52trQwplItHAcqC6GGGubBt/V3uJKEScTOFwjMbCUVw/a9Mo2yw
eNf8eZJq7wa6gjtzmXYDwLTntAZSp0XHQiN7CGQHQIte/eY130GXZ948ZJL966Ic
ZpmBvM/RbOLgAxxAMMfw7EsIQVlzGWb397VVMxMYBNVpyuEoAatYh3L4yEobp4+I
Ddt0t9gmJlP5Z3UkdM6QVRz4JTZEHpQMfGCD4MnGhZRXJMWrTBKdPq/Je2+/OAOS
MZgLytITGpq9svTxpeZxTKBOq+qRGn+3fSsVOnae2/gsvJpl6aDLpsH/yG/IQN7I
DzItnoQcFikigW9MATRl2m3oi/Xw/bXEZ9snS+qEJOuDjUOpHzleNwF6rzWuHIIm
2hXSeSNtJOjrdbeVCDhi3Gp0ik5CW4fc9P7ArM4yaZxrb1l+S1gdoTvRiZoKcrD6
IUSq3EXKkCKOOKHd55Z3PyCXjupUNedPporkZrGuv4ojXV6N5hdHxu238Sw5wffr
GD77hmHZOlvkGotO5r9RymBKpcqyvRs5OJ4DnDr8qq3Zd+6HKqUQ0O/+UqxFdC1U
pDNctRS4FDiG2Zot+Lw1yfQnAYTpoZxoiMEc4Dd8Yb/N+ToRuf0Kz49r+W0O3Xpw
5RWLjMWwCZPvI1nBu5e7bq4gH2ocgISiS0bbA3MegzzJfsYzPJq6arFiwlcPA6BP
0GQcCyvevxa0cFwZtbQFaAKkPPoa+GMfOdydfsYQEQ5JacApDof9W/KsRYOEzLdY
217ikBIknzTtWpWwNXuJuPojm7X1a3Min0cte5Nw/xOZVmJ9u1rJHzVTzF9Ma6AF
k7myiR8z6/GRlmyfgFwp0jCyBisa6ztEuaQZxJxm4ZncoU/e4PRJspPOCygQ2OUO
xxM5gEREO2ZZFPYhkPH/2MSK5+B7pzaF75tONOf+VmzkQdT1nq07ejgKstG98gSf
40Krn+f74CqvZM54nBOXfV/xNCmPbglsi5B35aNchnjczGq6GsZsR2+azvvrfho3
VpdGDSCqWyvx81RAfJBNKyuji9r8OjLL4JZjR2wcr0q7r9AVJiXmoOpojHd2MDui
d6gQadwvR61HGtSVwWeFDJ4centr0IaDwOpVAy73OAu/BlV5o9T6a3U4+AcG7vRJ
vwks4LVZKmZEwqA2iXd92brNCaBMXq5nbKtt92Y2Q+CpAoJ/zwCEXH1wRJfmU3rT
R55v18iBeEwHYzwZvjYgKX6CptoxwyzENMgQltbLJytetwbqlMb25Y03sMFbzFjh
1TXpNtXKqyRFtTrNEUoe0tUcOdWbooB8aRFRGwxNxZBTJSYAjtcCXfMK5vPsPu11
RoLQ3SF9KiCmbDQZGbo95E+uuOY6eKi19vmc42QlWCPzb+CWJCo3v6vR0Jgmb2Zg
Cf259b1R42NmTPlGV+TVXKEJvgOgPD7LpJuzP/dBWh8ArL1mLz0SqNyi0QgESnrm
w2K6ChNNCnuu/4Y74aDwdeOz6P/hFcGL+5RU0FGyQyKAJpO0LJGKThgQl6vxS2zv
4wD4KuHhx2B4HSLZb76rupN+CErD19wQ4VGpvA04N655mod9AaPBrrCsMeZY3C6n
8FbUtizkF22dGjhWgBWBoAonxtc/VW4mT6DVZAQPbGZumgocEOgZZ1w0/LNl1zEI
jR/DlwKxu/KCpbk57Jg5P1fqG1AkBPy0MipicZe21nkRkn/HqMxu/xupEba/an8a
/QCDbouC4QEzqq9Z/LhxqsOS0SGZoa+c6igbCfI1mxGrlWeMEzAKxCDGDM/+4rUG
7gvstJE86A1aS/Mw6fJg+ELlOJt2HAjyYaxABVj+hxw+LScu1vokyhordHBXCmFs
SCM3b1fYpemC6zjP+V+q2gNY2uUJt0T560N0ZMy2jvenAcQB/MYBVXEzIwXMNiS0
5cJpEqCNiFN752MR21Fn20ftsewFvBh6WdkGDZvPf9g7WiKatUVc1o9bZAFzKsgv
d6FIxjtqTHAfT8I1Fb/eyvpd7wGI6UoK8YOWbITYDzGqNZUbvLTVfkHzVwKeJiQL
gpmR97iH093OqPgogmsihTt0sxfYINPxn22cUlVRbARnVXOf2Xh8F9ih430mV+IQ
iuH2ixoilj8iqGsZQEpyYBbQ2bnFnh2xmyYMsGEf4WWJ24nlxxIMN7K0Ga+foVfd
meRDyyTXpZNF+VK8MeAI+N8lGQuf2h4IWcEbYTta/G0E4XSgq0ZKUqsiW+ETQK6C
3mdKf3PjlTflXGK5JW8Z5HguA6I+c4Rv3iDR9cWeUtug29D1Op8uw7d+6PZ2fe/8
u3Ejo8Kl7sO9iT1mZYd2EcftO08BB3dZTsjbFTUjXygljBIPFTNEgRyfwkYxQgqE
V9Fj4ZEgR+xEKt1JcxL3gRFYHE7zKqZ1R2A0A2mdYDbCazhLrDKupyH10d+KPW8C
z2mPtgm5C0IFuJFbvWPD5kiG/ucLL2tqKGzpOifUzilFu8WOumDkf5iIPTOR6Heq
pIGGBG7ZG+FA/CTqPuun5Y+8JffjPy80T5/6BrtDHeHxXB7e2Z++XQI2J43nDm7m
MkiRpLx6M3wSD+XO2lCPI6eRfZrYf4plj+GGv19R6Aiqc5aYPEboz51hkihvGBDA
Mh9lJYmd472Mc3zlkevwvaPVNy38SIFUltyMlc09uN/KNQ0EiL5VxK+mq40JN06A
1n6UqQ0ciRUP6/IFZZEkb3eyK1FngSPAqIbrQqLurqhKgNTTvGT8fJbxcwQV4DEu
f16U/DnCeFD1mCudxczNQZ2JVdX+Nrxyjdv2L55pEYdGcWnm1IRbFqF+yeAFrDhZ
4mDVuo/XaAsFruoEqzu4oCexcnK9qi5CF9VLg+2cIE4YoNo8/nPBGTL2ILEsR0fs
ECn74BP60oPYkAPq+x/0mOt4yRpP/C9AsZh0KlwVWBHSPnBC9iC55Qjm59JcDFwo
mY6WDOqvhTTxT/xeY02kLi9JXBdr0kb2k7MzokncoK4uESZ1RVdyD1CmAU3kfrRO
0GrDFsa9KacggixSVA8a8/hFRra8ay+iO9RwSiwdJs/WZkB1CsegJMmAW4Jw99vP
gUq5wbWlgOthEv7yibsOkVftRaFMcqVsTBtL5YGVlkwTHh9/KlMZeTqQSz7esK5B
hhfjr2CcUUfXkdLsPfx58WPHFnS4GXlqdIq7bQEAbuVUT8SUfdI1kxLx+5RSMrM4
odXSLKGd68+f/7rFXrG0Z5vm0y88SomRIS1JbHV1iMenC4zkojx53gWMN+Sel2zz
ZDRuBFgP7aiZZHeHyfRoWcxaOcgg88w4CpIoGl0p8E6Eu6AQHs1qUQ7yIgsQmf2C
8fpYUcyiEeTxC2ffUo4UcD0hmSnNbsdYwu3iXbT+Y6ZgxaIWGzdCjQErOPNVqhXa
MNFfrc8dRnZYyu/IHWUqppNJbHWyCAq/rwW4GK17IIZSoQMvMlg+/k6glQD8/oCS
JrpqR1d+FV7VBb84oryAjB5/PSN17z8IwPo23OWWYOKM1PifiGJULYL1o+jOGPkQ
pINJQFPyP1fZhX/GUz9dE6WhkTmdJt122+pvlA9Hw8t7qIP7xu0FuHwrQDjSopD2
2fzwVqWAKSaqMtGxCuPnpKZ/Pv+I4ivTTPfTox1huKeugnQy5vcK8OG0X6CH9ilm
PJJKB3hR+mMBIjKohS17Z0J6351R92/+cXayT5yYZ130d1XlvIHq+n0X91wWmgwG
t2f3QfjX5KZ+6PXTKlJCstzTspQ6+ekhzMM64rS+6pqNksTojM6EIdmWkLbGLyu9
PLriha61Wtshlwful/Seg8DzbCxxtEq/fh0f4epQq/yYtsAwvsnLUKSYhGBcyblK
KyVqPjtRwimG3xI4VjHBF+dd8Vice6cnCRdFSzMu1cSRH8Qhj9vCJc+6ueFgX7SR
p4YQKWtU7r8nKC2wRC1G8ijg0UJ6GBOmqWnS4SLwgoV7xhIl7ufyi7ucV75+4ugB
iL3R5SExhlAqzM7RuhuZWayCPTtT0xfhGqDp8NVka6H73v4k9TZ3g6EjJfVFQpTk
BDNAjMg8WKbD5+8HHS9psi8124s38d6zOmzjKEWXU4tNBo6Dm2gEYOU6TCoIQFdj
0TUsiZ9xz0wk6bi6rGAlVscD/1GuOmuOtrkdF5F34bWYoAT6Mqq2ZDLbCuSkHY79
/T9rCutokMjhaI4QfxgyPdBl6Joh42JV635MYsOQzRqex0ORmsAt/0uYLvPAke7p
dUZIgpH5NKEb53cjgtZRKyzsQOaFwhXKgu/JRes43qqPXNf6cxFOTQ9Bu5YIvuET
69gdzNyVf3GTeZ2/wVkjGR16YLzg45PQNs77xEK9dRURt4WyPIpom3sCEbe443qH
oKYgiLAgM9Y3iDEycCc+1McKuAszym0D9kC1foEuDYwS2W8j4gqS8voK3uoLX+qC
x6uQCBPmdSWYWIsfNX8WpFVNuMnHCMibkEhx0brMbNJ3tRvIVfbPDW1IDFdJdWMi
wxGF3A9vvIZVvZGK0wdb5TktVismsRu9x8ss8gJNJZuu7fbN/QwxGFJhIATKpui8
MQfOKultVHZBEaFaetQOauqFyuaF9CDw5NsHo6J/0bavxm3TIUKLrRn33HeNNhHy
UL9y99TGLA1EddEm3A3r2a/hMrX1y5fc9mCX97nYo+s9fYlRl8Jf4122URzmGPwL
LkQV7jOx4+ihjUgCobgNt2kmRKDliEn6Z4mmO01yGQeGoByrZU3wMlBs6lgPJSL6
2glI2kGqKSONkROt8+bgqlOtPJTl9vhZF1laI3+HJSpJGDqIYJUyoFaEEPzUG5lI
eMHvDSTKLNundguaMECxKAKUFpMMGaUnOnCiFRBZ2t8js0qLMEYz/gcPTLEUi+ND
1VBPoCO+ej4aEi9sYaILBkVeTSej4Nc5qO4hLI3xD7QUFaRCnWILnR//QtfdsyBe
YkVpnpSJ1RsKQCPqnt9BnuRqBoi+yqaipvYMoDWsmCtscTkDbOs1eCQMytN6ad4x
hyj0bWqyJQsNp8WPkbc9Tt4Co/GCRnhgMPOSzBcxUaeNGwaS1vFtPlXCVjZd4VcF
gxgDssbOw8hBkCFL2HqMvYltDH+9CBAFlhgmzXf+G7X6y5T8xtijYGLpRzsy0B+T
MqG6hbAIPcWwQR4Th/LN8dOn162EYyAzc/7D63o3Suc7sm0dtsLVgXTJKSRVvIl8
NHhL11rhk6f26UaNZx5dHXAyYmyEK22Icac/witGAQApxYrgf4eYN024Itp2HgTT
wW05KEp5xU0RAwjBXjHSqEEFj3bhCQhVARNPo3NH8LXqKmDaJHosvnnT1Fs+Y80u
Ggr9OorjCnS+flekovsA+8ge9ek9gCHxoPWpm2zKF27coFV6qytoxvHwAV3XUdZv
Vv/+m6cI7/nazsbydh7eeHgV/tZIyo42WzG6MwU+cn191gBEGvbNBLGGjn1DTPco
rLMC5sfnvNTpX0bLoTl9JiMCWiF5QZ/akMvNE/RY7vxnLVDXcyYuyma8k7F1Gvab
pTiBCCFqmM196G155WGXzUfGsVJCS/gUnK4dJP+x7bexG/sOrSQAFSOo59RuPFw8
McMHcX8Btm4pUCFEYp2flyeCujGelLPUWN82sPKz+LgxzYeFMSjMXZBSuC/3fi5r
55Gg7azDk3EGqPXJFjlN0KtKUj+N0e88tRta4lsWuELyvhm+CE9hH9pOHWiNsCJX
PTY91ZPw9BEm8KuZ/YEPCwGka6Xocg3aMvHA0QB+ImJ6HcsnK99GpxLymhh2RsPw
wnhEE2aKyT5XiX8T8J1agGD7FfnZ+yW9gyqtxsi+MXv1J5ZxTMtoO1wz6o8BTpc1
mbfLFMI7nIa5wBOahB62ezkOWw5Ks+BNXj64WmU1/yIr3y9/GoDY9cFRBNfvWZ09
FYzfexrh19mt4Y5Tat2/r45mfKomxKg7CVGMmNMUr15cJ0gW3muEUSuRffaraqjD
p8i35klFOuWIlHu6qMfJGdVhTOYxA0JFhAaAZfHBsQ+iP4tzmxrO5t7v58UQevT6
UfM9qjILAwmEiIM/vpFFTnmYj+wFLH+HFEYbKhQSkN0egvUUI57rp3fm3GXTx4/6
ASSlgpOtYHUW5YyqiIy/cDb2MzozrHBfs2NeRdnfPfrB/PdU7a48LzOxjzt39wvT
rdVU+B/4RiJsmf7FgHbRhrrqbI7UdaO0KIK2qMrEDVmozbGjn04F8EwcJ0eATg/h
dnqgC5/w1oMsgq5U0/LU9xfnTRjCEcu3uBB5VmpQvwSAmD4vvjWV403MXim+21HR
mae+mC+sbOSR3tlxCVHLevaDsjVDfzGk0gYTGBiUdFmwIwFF7LWQ9aySv9lZ8Os4
y6kZ5SEPaskLDk1GnIHbkHwTpbYO/2nUdwU+RpmDgIzJ769qUmXSewL05fHd4olD
JP4rJ+wL3GnAo5ZgVV3sE7DIiTHpupJi+8YRdjTeSEtf+D58Vkukn6pLMq2B6V6O
OSLIL5eVkUTAd9Xh2NLCrDBQKU3wWhRKekEYXIFRFVYx0vHfeF2PyFul2SLtRBI9
iAVOgITtjtFl5TJGxQjFJgoU/+U6gjQlSdtdHnxN/TOXvp93Rr5ov+5MZpbqs4wn
HL/fmkdGkH2wtoFRazDFc6EgaQMnEZarNZQM66Vgop/hlUDKTe4UkMTRdC0QkRVb
nrr2fbIjzZrXQSB2LuE2bWmRjBdwx2o0l4XauSBfTKG1X4uSqPUp3FjVvUYTLg3D
28baSZT2DK6nKsiEsiHCsXtZyzFn/LzqVxFyxUSzBm505H8CZBPkCa7zMyC/3yvz
Zy6DNYW4tUpcrqrrjsXbTS1kmVPm9XvHwS7NMLe2/O3ZFKoIMlGhLv87CIBLzUQz
A2miOmKp4hqTn5wOEBWk38DeyoNYihzxvdtWk1OqYlMP8vYOWEk+S8ISLESFBGBs
mnALxJndethUIPBjxWgPQkFGaXogIufpGytOzn8lfSYkhAxwlXPcrW3IfowFBPAR
yD3NC4idG3rlFbCQe2nDoPaFhKXptOrS90f4lK4NOZt0/NhmkH2kABsxg6TzggHI
KX0xnSW5Rq21a6NAD0nVf6fZ0Z237ciH0ZNSQWI8nt8FqmYjx2+6ZhGQLzuM0eAE
Ac7S5aZirAXjG0mzed/eTgLXX3NKiCpN0+UCmCvw9OMHykx2FLOrtaIIhm48KekA
A+xxoXEYLG3E3xs+UGbYGp2DZMCE61viq4aXZa6JaCw+9iRkAFN+PSjCqbG15m6w
UZg/wrR1psnNSJPjqxY6FuU9g0bxnyDsXogaQgNxxklVEvYop6A62MehEeKWJCjh
zB8VlOYJ9+vV3HMdYW6D7xe+w5jonBQ1+EDOgjS/M7zHwinT4yAxkOhsAERXN37q
8SAojihmcyJT1lKwXrqXGWFLnEVslvObZ0A3/RFfOZsWT7gH5iXgQiWIxJ0u1rvO
aI7AL4zoNiY/BQBRag07yEReYUAYvsFeR/Fe2ZmwHbxm7AGW7WQQIM5M8ZAb1f5J
YkjH6D19DriWFwqKntzkh3H+bKXIKOCwEWwHfCc+VS6Mo91FeVPpL+ZESlx4/LhT
jOXRNLb58Z04vgzT8s0LptRra5cMpGzP7DM8SaF67fPpwsaMjPkzIuDOYiU7yZuO
qBrjcRhCRVkoVJXdhem1qv3d0hChdCG62dk7/ZgFIheNoEeDCMWchg6ZNHebFv11
nI9Q/izhX2Xie52ckaiSdm77y7Iefd/ldrCLuByZVltYgraPlpTizPOAeaMocdYx
5GARGHKhDQz9BSC1xD/eHw8j0P8lRZ9QqeoAuhed7sVtENCQyAZ9x8j2rZgGzEmP
AIMHH/tqKFc22FyiO3I8sDmIVIMel/d4GRpKgcaREMCtxCogSSxtOhbZ/Vn3OslL
aIli8Kpi/f6dTTNkYxsNJTZGddglr3Bi8iLhADXRbco0AznAqNdLO7/5NZWWQI+p
jJIDwZbeV9asrT0Ei4mSZhKTUdqD+PFXllm+2GeSPDmpJzMDPIuCoUn/XUGK+muH
my/LZr4e36Az4Q/+c3WJQ8qmhloxP0YWrMJFsrGBM0wG7gTxWDXl0EhpQsQp8jUN
IdTwHn9p04Oub69D3FvkuvOQgwnx2EvTFPRRgiJdmsyFd/q9fKOOHg578zDoS2uW
d0n1aEqYjl6znk9I9m4TynN+/luDpYn8SgrFO6jVoDdHZE34KFLPjEiysa2znBOJ
9i7o6fBdAFdsSMSwiPpClqmpwZfOCU/nRAHLfi04raFRn7HZbUFnu+VFOwoA4NKl
jKfN6O1d9zD3r3cjClsMoHdorTrNnwVxXSuKxCbziLIlUgimLj/tsuFXbwzuHT+c
jLcmO8Qk/N/c+N7EX6l2h7mJsLQ3stmtK1DAAAE8fuil2V4OZviUfy9lRvTGcSdK
d6oL4xlabM/l6FUwA32usZeSifhH/8vVBq+Gzvao/+vq49lujJ+EWmUUbLxOydnJ
OspI5kdxdZD5M32Ky7Xbq/zqjj+AoYuQfEEFonhC9wAtu5TvAieNGwCmFM1Ueb5I
4mdMDJXb3in0n67SXDipB72ASjn5gwQiIJUJM/yfmhqp9NYtOp/zE3NGgi95svGf
RN7repipswltjQJcXzyGgpQ9hB4fWPVKaQNKAhJxAV2KNYuVa/WPpIqL8yvPpTp7
19tbKacLLlJo4OzmSBEo+Uilh8XsSi937R8rXeKuUSMIVF6v+siOpJrOxNETWI++
7bEFKYQnaLFRT0aBvByuAm7PuwxjA1UGLpD7pYAkvmDTr7+eD86gztEjfkQRxx0f
wcmzD3fx41qg9Gp/KNw3raI0CCuZmDIsQ2B1OvGhclg8FYwlN/yraTgiJn2Xock1
b9Dqh8BK7Q7t8Yx3bAgSRSLGryzFGl9kN00TMYLsgIzKbxW9XF+h/hNgJZ6ICRe+
DYEYJty1fARKj+TVTTJk6mbKten1q3Af8JYW9NPirXMlCV/KlaOFlwrfM+YJRuDJ
wu5P8lObNbpmkphwVJEcS1fLf8kAL2TepbeyRnX99iSRy6G0FUGuitmjHD5yRXFf
eOdXnkICqgtP/Gggbvmfq+ZkjU2CQQJ12VDMpMUe8muF8SWjxmrvB3IslK9J9bUf
CdUfCXuxTs4lJZCzmatRcvcKKFi1J6vvvA4lV87q/DheocBvxdbyKXO1BpzSN8zx
CotluyXgzmIsI+pKhJq+jCE+/GIqJq+LISceAjQcYik24g0xElxVMUkS++UesKbE
y4qyMisxPLm4ellOfUGPR8FbjXR/gsBBQ8A+IsbmGI5tkey35XTVC0NrCLyb7Wwk
uoJYLc1tIcnifj+KsB7BS/2dIZDb+pJaryw9gauh8AnUfXXosDMHEsiB/6UnNB1n
9V8BNkdE6dNV41sC5ry6ZsXnQT+au3b3R1gEym/wDfEvnyxyj7i/aJFrvXuFl1sF
jIRkq7CCd9ZJPt/UDXwQMxgxupoF6C+RQeT8Hf+D7hGHZVTJpq2TX8/2z+4xVflD
cIsWMEo7eFN5M7w2tcVBylPlvbSE1nDDi9lzZ+45OxeLtqTLo7uIjClN/o5a1IYt
T9UH14PlKPOzCbHdHctpeSQvfhCRAX9fLU8HfaqOrIWaondNpzRmD2YF1XOni9RL
rszq7CbhyZ3RC5r13cZPz4UeaG7+0im5JH8SRKp7Es7QyvcMZPO/OvBt7vqOhcIb
U+xd543q/RAOyD711NH9mU+8OY2nYCnqJcmUd7TFSWLQkUEROpAhDbGsVk7M2zRG
/P/m80QRDpqthILP4l6whiHPxXzLlpEeygzjuV9JjlQUu1rEO6zdjNRvyPrdQUhJ
G7RMn4n+wrIH3pWJlfpmMBl9xnvj1z7xMM1J8/eR/MSf72l4/YxaMPB0hcLFDFZJ
UOOsPZya2jPhhtRnKB2FrerFXXswPSPzdWK7TBzkN5Sdy5VL1wIdu9GKTRvrAmBg
nhUkbt0e+wy/aAq+PmYJwuNn3YeVlEfnCrUH67QIBuw+W0ZqSFnh2/Fa2fVD2BE3
rGiPLsH/dMlO0F2LMco9a/WLpZH05jjdhoZX9HbIK6O1Gq0d/HlgC/X4z/zsmQq4
PXaak25t/ebEriAZzxufPgAJSpkjv8pwZEkQ1WIshvJa2i7uVCf8RNq3jFZmZ2SI
gmN0bAJPY9Qq4v76c/b5c0Pu6JOrfy5597K1q0LbErx+D9/PqzlfKXrXDWHPFD4d
ugEmAWYXebV3N/OBDVQU6Dezr0+MMdyOZa4jsVOqOgLW1YJBmwTKWfu53xcn4M/K
VQVT2ve/+4HgtkzPzmsDqr1ArHuT3xSKlBPKr49P7DmnG3GBbtQHSFw0xbexKPcR
jucW/CaUHK/2lAFiTBZjd9aHyI4Zf2XZPacRyabmS84nZ7wRGw52eurFkZGd2EJi
gbUX7DhvYfom17TJlu9UeR13I1vElOHQrKWH8fTM4ZZkE5MlY0JsYgH/1w+R1soA
yPQdy3BTZtAL6QQRMrLt9rjDC4Tt0+ZG1N8kpOXBlHT4C5zctp++wKiSXyJPfP27
ybqqhFv2u5ms6w2hOE+G8dCjtdRV5QL496pQ04bOnb/fbzrTczk60bw5fEgJwSce
tvjH4MN3Zoby7RbA8FUJ47VYnQeqiT5/CqWFaOd0XKoVGIfDPuCf1uWBRSBxJGVM
+pAozmCXorkhtTrmCUvnqSrZB0R2n4tOSEFArgX0Nv/7nbJV7/wgiFnvM6lV3yWw
VyBmK8aFu2IypBGaDAIB81a8kwwCUch7NpFT6szSz2YcODwB3l56czQkhwh7wKyy
x/H1hB8jFW0T+H/GnEfefzysoeOOuvutubuFnMvbHvp0oZZvDojGz/YppCwwZWrn
WoaCn6FRg+bg36KuflT/NbrOBPGJ7wFydXRRm7XbRTqpiIAYuq8/gpIzZW9JsSIi
QABB62WT5Sd+3PrxcWPQxdkGEFRcKWHZZQ+8VPVvJf0LCDvVeLmzYGE+ciEUsPyS
HBdN/cfAWA8rpZLN09CvMZYDIiquyX4WieIWa4RloF4VQt+JopAqRrwdQUGuJK/8
ntLbHLKDd0vg6N+qogcVoVuGLq9dBMBjkAPRwT6QG0hCeX4CUBbafb3umaMCv+Kx
G0u2rTgAYsFHxKsykhwKA2faCeUZC5kKz0hiDz6dcA8iKkVaGmCa41YPrBRYPHZ9
NGv+1U/TMU58XfmwtglRsLaIGxwar9aJOrV4PhLxtI/RKy3ZQDo0rR8hDvqmKsQt
Bsun5VJJPJCR4dJkpmP7daux4E1cwSQoGjx6hP7vOkcoB6c+yDJytBboJZSN6uj1
emkOHJC0Ij5qN0rzJMavSwYktBAIMlBjnrVrXAWe6gGPRcJxdaWocNzRKZd0/6nn
2ZsngGW1b28nEj+pHfhg6rEnYFZrbtV2YWJbBcfcTr9iIi7iaLeFiUQ/NnM+ny7y
mNeUkkJ+v6xdyhW7NdCc7U/oFsfUQfvTOjCKkg1e+8cR2GBCS39OFAbvhVHYQDlG
C8dOeGFUjH0xahIQBcicrVCZEKjDaC5jkpIhdXl5TL0aVfWV2TTxY/K03cOUcPo4
vN+AU9Ch+oL1CNg2LdJ3ueIqEskWIngm5an9kG9tZVkz/B0jZi0WgkdTtIYA4r3P
Lusz2F9ymKQK9FddhorGnqueqMNdfon3ABXBDUMAjmpWacRDDq/Yt/9tWD/sbYqK
dha5H0CjMz4l3mo7Gt4/KyggtiL2wW+VW0Eu7CHT7engk0BBX8Qxbfa8GwZtKrTT
ZDZnqGRHIKMOB+TtqpzJk22xX/SJVGNwxNAm7LrlcloBwkKzAD9K5WE7S9+O5h4n
2grxIUqDtdMH9xAX0HZAb5HOmwru83OQmECLHJcFLslNgDHQoXxX4zWjl0y4muhv
a/Gbx9fpjktp41LWgbcTciyTE6Lo8CUUw6xEBSGhpmRDQFP/Es+5RLiClXChs8YL
81aNhGhYtkrLVhQOzux42tUNweyGxjhXGtSbAkZXwjDlJHHY1Esq0dH3qmYP9IEg
WciZQEwV1zP5KCiDHe+wCZFQAUCq7rrP4Nuq6jmY8R675Nr3rIaehi8Ttg0RjJbh
qHl/rSdkZbMfHuFj68AnnBMp9IEXyccsqQ1UQiYgNlQ2zBkB8/aV+KAbE50LLAOU
4vrm1eoUqkS+0tNplYpL3AR/ZfqfBEKlSSGIrZ/VA1fOACFv26o0fBaGN1f1Sc3M
9Wabzqw9RZANvVluoNbif1Yne8I77tJpMFlA4tGrwH9tTNCq6HNtNSKK96Ihf4Kv
+aXSlb3sa6WjwZXcfjFHyvLTOgutDWpPTaJQ3CaQz7mymPAOuIuROU0qaT0mukD/
RDprzW+3n1tFmV5VdhpcC3FdHvrf70NjDw8zFoSeGQKJrqKM4Ma3Y/1wdOUzNP2m
XlJMXTTgYRrpX+gSn3w8Jl5xbkIpV9YWsYwMqGHSQpsIfDFMsdO0JjlqVxIESz+Z
mQHsxut9bQ2L98z7sRqJ4Z5a8rtOOHqkMa2IRiCQ+tAw3HO+TIMeAJDD68Ixc2cG
M8yNiHWyFrRHH8LKLCAApAnkQlBSMgRBKpYN+oAJyQkBQ9IcimoxtnTY6QFAOKtM
xRzoFYQ1qgdyCYCuAacDuTfHLAUyOMoGZDluoQmtuaB2s5RCtjJnPZfly6cwhM9r
Vhlw72d/9mLU6qDlPDR1X4SZ/lMp7YHIaMo8srHcTPzGnHC6pb4dRubKF1AcAb3f
MpxWasNBON6kmTtf1RvfdrSvESnFG0AFROGSOGOJMNV7X49BBcuJ6Y6dCRxTi5ET
ep+9BC5mSmzSmUJjKLkKO307phF+I4/TGIsYcZxZJ9btX9Oi51mHezpUli/W1fA4
1j/e2C8BSHfQM70+1+7Meb0zeUIuJL+x72YB/3SRd6krNLhMCJIxei4ccCvTG6Vg
a0J5e2TsUgMYXctslb80tIiEj7rqyFOE92qmF2YeoeKtTphK5EHNpup/OsBmUvWh
1oSSfoCPRB+q2DFOhYy+U8axq994TLwhuO7itSHX/rttJnkMAfiGFzHRH+OZfq/K
Gdh/41Pf9Ke328jPkWYL5zZXBi3qEov90y8XXy7D6DuVjJ5qBqPCNVnRl38fDsLt
MKFZXZvXpPWEjBXgZa1tsb5OLYp3iblyVfJrPeb+Iq2brBi5dzoQcDCCqJai6nsH
DRMybxu8pWfZPQpXtzk9A5F0yybtbPluOopKH9vimdlX7g7SFV/DtE0eGrjIbFyy
7/BexexAWXv3iFvtHSpL1U9Q7TiTv/4E+hwVYfCQ5Nbq3GsfBna7quwXjSZdSl+w
teuI8JZkBYZvL3UIy/QgJXLc/iq5SyNCwaiBhDMVuj9ku+hoqXD8JSx0k9a9NvUF
QJN0OXc0NkH6PNDCUsA5mM+w8zsEPvPdspv3KwjJyfxmird/+EkabxlwVZ9sSJEB
CntImL0zoYl41a3+401zMcTTBtbqd3lzn4/sOKl449iFx3sxSVHv1RKaB9rdjpdd
DZPHABIf52/6btwF74BRyrrXddFG4zdYArvXNTdhwIV07KAGctj+So/MvJ/hdTAi
oV0JXzWeot7jFtwgOmZvzR+PHasGI1xNIc2m9c7fYwOy4A7xy70py1weaIFkdGKd
pw+rc0oBLjjuiDDAjR4yMiCgvx/k2lBkKCI29Q28dWeP3kli6YWaxf8dfGDBN6z5
G+FS0aqQVWzXnyc621nJt0nktGjdCns+2+08rGB8Ja7DQ0yM5bE0yLv8gsg0fZYn
dCZQAoSeGCEL0+lz8b1mpuLAgbM0wypAJqfmSpqgLiMuqnXzymiKYrPKa6G/eZdM
X3QzUlbvD+C0gKjUyfoKumaBsbdp2f+39apw0Z5Fp3lq7Q03DF3xJMQashavVQsl
oX7N7cfUc42gP1fU6q+typko0zsWKMGpg058qVxng0Tz9E00BbwAQJO8x8VwTbKp
vIPe0AjL/7DSdzFQrCJhGvpZJ250TEvewnqy5u8WnPTPZb3I5SYk6xcOQ5x5JCH5
P+xv/is4fLun76B0RX6L9rMD3PGA8OF6yrD1gb/TCWRq8/2k99d1ti4roUNbzXUM
M0IiY7d2AwXriST1UvgzLtul68f7oI/8TAFVSc9g3wpYyw0Hq8stXS67PT4n9rnt
bWtR4UsvX7mivmx6jjRx+6REA3R+wsKXiNKA3DoKcNJXTZ6TtChd580blZZlKlAU
yQOLfkfmHbQijx5QY7lUY2Ek9nwyaEZqPHgIJ+5xWbksW61sCzkU8tO1lNDBTK7U
Hz+GizBEtOxlV8+o5wqk4n6bDnm5coc51TSm/C8FO9QVoISILuC5yqBICbWkMV3E
WcvfSwLRXQtwiL8dTPZ1OM1QZnQqUcbr/lyGrkiZOTZpD1xdTdYFQPe6K5SyGtGY
gbsgJyaagR44mJ84T9FgZRgi7O62HqNr1jXYV8gs7z44PEuM50poP566f8LufDUd
kpu3qX2hmsB7nYRvGQFJfOuv0qQqOB96nkucFGR35RZAT5tqIznFUiFoUwCbkNZC
yNnODkSve9fzOtil2j6/CLJ2NMA3RFdZcQQIKi2yuxdKbi/mQTz3ig6UOj7mE8k8
gDl44K0zg7TQnIUuFsEUfgZQxqQJxHR7gWzgw+ogPv7NgcymHx8D5ghN+vfE/oSw
T3Ob92aOq8F6+tYcOdecJhvoNGJDZgXTrzDz1kQsXeiYqUJg/F3KZIUtMa9CyJE0
QN9q9D17uGCgNDJWHyqY0glyOQQKE7QoVLL7IKMtElfCyMBBid4aQznCi3E9lAWv
aQIyUpfPVqmh3KMa+dgMS19xJZbDg0mnpXUSZCMBg512jIBAfvJhZB2960e5w8Rh
IhDY4e1xJzk1Q9gdmwdSv+4l+WCCblh06AjaRZCCRmTOYqk+EwYbpZkpmr8YL7A0
Q2JD/I+8fSmsJUJAfdsCkZAov/27G4pp+enAHz1IMAhMuAa0EIXFI2QNN2F1BPIW
Mk7VUjXKveBu5ugkFEqo7pa6VAOh+NfIhiX+bHedF7L4ZO0mo4BOIZwY/GwbZmQ2
X8KdYExzyGNW3j7Zb9ao86CoXCIz0h8/cfhO0Zj9bkv43cG0is8idqutbyGmX7Zl
sbIbLzCl8Wuy1dQ5807fs5/RMwAFKnerDCQ8exNZW02+UR0uhrd9CJzZG1CH2ymM
lBViQn3d0W1yQ+VeCSVc8YMR7qt767Ujfj0G1i+X/TZgA2Buc0HNYMc5TWSzYwJx
jMR8kuvw5gR8eehdb0CFJ46ljycOiAdfC8SxdciFnJz4+yvkg6NpW0xtPqz7EKjt
RRk/6OSIwfpsOFUysP2+PV2V6veHqtgTD8kCTyzdW/AwvmP8GpeBh6+gwW1wNH6k
vqCmuaYGDDXv3cviFa1ussj5VLC6tpMrDkh5nTtC0TCBxOeLq73ph54uVAS98v/m
NAbd95iV9OPxQMDNtlWGOv8bEGCZ1jPxmDSxeTL4AmOqOJ55Q3TlM1SI1QvZh4HN
iK2b6Oe5L9/bfUPISVvmFxzJTMQnoQXYwy7K4T47gaeDazd2dbivPAjsinIUenGR
x5BeyKtqJgptL8hlEkNIu5p1b66AKqjYEiAgBuGWCNC3eXeCWaWsMV3+o6Kt7A+v
B1wrx+FgVMRy8Rqdbx1+bNRhZgYVZVx29toc3FRrWn9r70MQIb2+J7o/V1ZJz5sP
HMYdxnrGwXh5oz0CNwRQSXRmReP7xGucj2l3v78A24CC0i2vNHfUzr6L5y+n5Ora
rKWhESqohaefbqMhIx6zpqD4Cah4rH5aeFU7off8Gtk7sTyZTlCjdDgjRxf2qfRx
eTqfAv1DtGz+YyHrBuS0KcnWHCxVDPuP3ifCU23doNf8PHWbi38/iJtIRjHXV0U3
OtDKxT7G2QDCXkZ6W5mDFkMNxnQyJxTF/YTeYvDVjIHboQQe6YezRZpgwzXyoMT4
jFyDLqBMBV6POGnvrjSAD4SPOz05OrgO7qXxwMAMm/1QIge/EJMASaaVhsj071tM
FIGPQ+3MXKGmT+bfv1/SNkRwNYSHMGCIW758fciXkSx0pNdb3jCfJLMHRX/IQf1p
Pc8rJZUTkCLxBvlUdM/Azn/yqTVVWNLx1+LZ0ulYKxaw3xd5vixDLeV1fc4IP/O/
yjs9zfgUz86GKCDVCC3Lxop37MrFpJW8Wza5ADxBb5LRIj4q23sU8ytaC/1ujmm/
kn9GdF0NlX8FKGoM2fFF6A66GDjjPRmGjHrpXxIsvDe75QUIqBDFqmiaB2BfX8Tz
IchzWlrMSVhkX9OzGp5Vnr7D1eL9tyBESFFdyuz+ARJYm+65LhhBg5tqUxskd7sb
Fk9ZhouosMWmyh6bIVT++cGd963GpCvbc9hgOg7I1iPFn++XvpPYGi0MK0SyLAbH
6GBTygAMLiULdYIyw/uKgR3cLSxn1k16+08FI5vT8mgLSys9BKtN7arHIVxydzPH
s+Yg3ANCyxwIIVCH6TRc5nw5JhAZk5V3vUEQy1PuhVc6XIVJGOh4yBQVj0Caa4+T
rA5Ukq5PUC38HXTg+0gsnu42kEyEn+67AvWLjZReHD8xo6pQ19MU7L3FKq+mxMgs
bpfpDLq6i45CnW+FHFFaFsOt4XvVUEx3Mtl45KQkQt3yVpjD8vgNoxFF4xi6pKqT
Hb6/I9/Vjhy1WXvv3LyyADAEKpbWYtTKYztQrxGEywebqpZEotSnf1OdTVukNbbQ
7me+XvXzImHpc+xAPZ9I+ELsQT5dEoycrZWsoztLK51j0ExCirewQxO5BjEZgQUY
TNw31Mil2n6J/vn20R+YsAeXxX363j5TEKV3wDFZo8SMa+d5upAZOeYsspaH1i9j
36r1VpRvD0QZViTWHsWkxpCtFTBhfjn8q7b5v0yzYPWkSJL5K2fl4190rauCW0T3
UuKO6ZyFV8xW7SPudfLIf08IsN6qOYStJADrQcItwoilRtIOd/5EoYukvYTeb056
8xCBHI28A02h3K7cjyjrLTqJJ8vcMkP7tpy5lHiJz818wOBKZu19Ylk3mOtpl51Y
klpQRdxMswa0Cdq8lpwbwT7ZeAoGLgEbI0jybMVg7z9PDmeyVIjpgh5NJhJTTWOS
l0xZDRyLFrI6bGe1n1gvokR4YIlx4AcZwWpAFoQfBTPNhuXDTciKn1G7mSUsR7yv
Pe6AzpKloM2k/65JvxBMkKcZNQFy0nA1LKh66HY436zLuaXWWvjIxI6ICwM70zLj
LvRnb3QCN+YULuq1egyRUGN9Hp0n0OuiBMtlyKLz5+38orFaEy49rYq9JLeP9tq1
i2R65moTjHIwwqyd2HiIYC7yOdrNyXNWfR/alYVQ5mu/s9iSWGxK2v3+dkSy7SRU
G1F2GhlRWAn/2SeSusQ0A+dXgz4ABjfOLp6ACXfImWcMcjGcxJI4w5NFZ4tAnrkZ
MAqYuCL3PdB1bySfphZYjPfmaY6G7Zn0Zi27CZlkgHerB9viQzB+oHgaOdArEfbU
5/hjzzyMmqgjW/8/1QdFjsPS3wjqlEREiRKbAGQ6vF19YJkXAoMLGT/mNKX17qnN
480R7o6pkcgC6NyqXP01S6eHSMTj2JxC2sfPhV+mUmcePaRmYtSRMheWc6MdBDYh
6elVKE9oJ9ez4HO1BqgurXaKwURdNimOnSzTFZM4JZOdZmBR8yIjTVqxTc9Ipe1z
aNh1eiActFXRD/b2MD7B9mIj6IQtzBl+XvccMC85WP4mcY899YWiODmkhc+2k75M
JorZ5UaOe22G6AdmdLsJBgiQIotwHbP4enbEKM/81AAnnANhUXpW84Oh8WHO9xIM
CYQP/CCloFvx17jI9Lc8Ug88f+tow5HV9f9wMK2Wo9PxBgBuVxiwXYXk4vGnKyVg
AdGKOLhRFghIkMfR/PNJDCxnfR1z70olTb/FkFODTJWIh1Yc9FpredO3d8n66hX6
mOwIaa5WWM/zCeXh50g3L4NxiFzZJl5sCxk65APJvPxDndKukxb+gqtsDCfCivbu
N1jG5q2wrOPadGfxeEEFs+e/vyw3IVvqDqnCXQAP39G88LX/f0kZ6c6zgxCO8rRG
X/haTbjC+O5UuijBaRGIjSdJyBH52ZxQaCOc740fmWw0Rh49fRVCyC8S6ESq7d6e
plob4Oe2QnnWb3t6wNs26EWAeK0x2Kq324SDmwexH4zBGeUfSn2a2WlgJmjzCdY1
R99WdLBK/qkqdt9fkyYQXrFqfObLoTT0AZTE/2Y4hEo0FfgB7xT+Icb8a9BflGdj
SZuuaK3NviVO+LbCzYTlF/nKi1SVLKftFDMmCsm7cFAEHEZ6GLkrvqb9qhoCffYR
6ZA2vtWX6wJSG5Zr7+kfjlFD3xjO+oAjbugZDweifX5jx80sZGaatQIyK5a/gsoU
uSshGmUhgG51hSUymt0SvX9vlJHBCKDolcIpXh/g6TZjT+a7WQbtFjDVWajPIJci
5ranMjL4ongqEly+T3wdmhtynj+wUuTYv1B2xy5zMsgoY9SefcSMbw5wFk1KTUpJ
RnixpuYNAI2igBVTdirXmsf0SnWpo8YEWiJ1DzQOudICBPXXchjdRQgiQrHAuU2n
H3iW6WtEevqZGB7NrQW7QDlLClZHiZVoaDABJQ1De0D8fnnnvx9xEXhCGrJ2SACt
HrA87hgD71axAmegNvXtXK950CFhpAt1yimAAmfV5685N9Okb1cjvarNUaREwndb
KZtWMwy8paXWT4e69HjgasMABVPw8ajnoIN1i/0Eu65C9ElXxvyAwY5zeolPmvEw
2h8cSQWRABwgNqmIAfFBI/ZKrUvm5VTCFJi+4PzWLo/rmjLISOByEt3zWuGSpme+
dLt5CemYiQa26fKTw4kN5jM706Ec6tAIbm0aNdtgt9ySMolbLootNviqIbvkkHDf
ph37IugtfFIkL2ymcS8NEKzzjhF7hG8x62MC8hloXltonEJhgJAA2BA6Uqm+dUQS
SRSYd5lyoC1ZxDJO6OrM5BysMADqWCD4cuJOxK50mlqvykGMxNw917bxgebeJAGu
j49jr5QztsA9hb3dyZhIIlkQi3EB7lMFbRNx2EiIbxaPRJ6Ct1NmWojbwtBUMJrP
35BF9AUi5/lRhHJuUWLb2Hlxl6fjIwl0pgnwLybNEft7IJdabP7smgd3C2dBB/34
i3qImu4xq1n78JfshP/4bnCiFC9UEgtlmLeRVDuD3R8Y71dPRQH9e8psEzcZh+f2
8ts8hrYiAJQAboBXfMhzHUz1bWS7WXFsyLuI+7Yz9ekW5zRK1gsCCgd/49Oo/kfZ
i9RKOk86jZjo0O9vvq07eClJjC5XA3TssmBtiZl+17tEqPKN5ePvA6jumkr83zDg
6cbSZYXtm5u44At3t6fA2G88+TMLX/u2WWBcyoW90YFnWny0KONuWDh1qhY/g2Kj
k9nYXBu6zmgpwgs7S1/gSJGOa6R5rpJkwkReZVI3txoIAKAouHgZAstDfRmvH3qL
4hJjoKCvxD9KDE+M/E1kWCqLUMGHFu/2zHMkrkrVRKiErJNubqagicWZw/ikWieS
+pL9x/LGX6NmyCCsUujLMfxUK2BN5197S81gBg+E95o2P0hC/2stHDjQ/eNNSfr8
H7rLnCBDlcwNghIKASo0GdvgsuZP8SDOhUr6DSoB7A8W7JmRNgme/UFSW7oikgBn
13+zDZkDI/C9mP1GLiK07otsnk5FuOC5CdreVdGI4KH09DsMBqGiCPPiB7uodof+
NzDOGucVuE+wVzaJTetGX7hAdqeSdNOMwELABIKc9CUmRG4g+mlQGQELQ3B9A2Nn
oupTL3Y2ljQe0QiHB3/QASkgkjUqZOfUnKxqzHpUCtalnKIbPRXuXiwOXXVwZ8dK
Y01L9C/fqW6Q8QtwzW8gM7/ZarO8x2GuMoJxHLzp80nKghUnzke4XJ6oB1xupM1f
e8k+EX6mIZ6A/KY98Y250zW4iOSBgit5A337mQumOQthfgsB4fXP7o5R1z4MpqrU
Jxa0YUTp4en0rPvVVSOQfsNq2gug7/1Ltup0zCw8vrxYxLxh+xEqHZ42bSCyZk2T
KHBKaKK/t4mcZ/MwKa4FqRb0PrIuV2VLx7O77QhJ8HrmWN0KFrE0JYpNdEuFqFG+
qtW15P7BwQZgs9q6hc8CUXGs5sXN6u9wB4jIDByJ9LBOA1V8u6oj4sJMEo1MpugC
iCawD1UiEt2PIsBU9tTtPkSkJx44zSfC3fa2jUxM3AHbkgUVbpHFakwsFuAKXXyZ
LpxmU8gRX6W6DO7pDvIagWcdIRVevvNK7UqO2zFALAym+kL0R+XuDh5kSTD2hEW6
x9T0fUXhjAF5LSjZv76KKJ9Qo+sBo2laFlR/npLa8HUFoCjHnGl3t2UlD+yBpkeI
/1bVrqeAXL8bhmqqzgJoNGWwoyNGEd/DhrtXZEIIomyCQxeXLVN1m/s8CUaCRSWC
Fd1FMQGrImxo6V20Nq1FsaVFs2/T+ERSsihtcsbWovjkFURFzAYzLJ+EhKuOSfDn
MA1pzmDffKZjjSci1c5QbTHeoMzZ+5AFnSSRG8JJwzmpt+N1rzwsQWdhQfXJSmCC
G+ZlbUvBHLJI/5R1W4y834F7DFsxmglE5aI2+HMINiXj9DdsJW8RVgbAgISy2YeH
95vn8nzRCLpYe0SbQN5WRu3r/+zrlj9jZfAPh2if3AhG6bfGwlKirnMtzX4gw0V1
EvZwh/XOH3tmODPuJuL3qu+9T+PQtVW9KlSx+55sXSTMvHzhUPPMuuALmeJw1FsA
SLfFhjTf259rgzYxu+zcG+BRv4hvYMZd6MtUBbYSiDUziQ4HKnYJxq+bzpldFD2S
jiK1HQuXapZ8cqTUsYB5EnOA2o8tHLUeu96OeBFpSlZXwVugjzUJRBzMnYg/sdFx
YAh1Cg+CgLsFlsRga0Kb5EoNVid4u3AOcqcth3HO6XVYcPRzV4PL2TCKnQEWClxy
861a+GaSp8G5hdaLRj8bVZ97eR9J4hLQHCX4TsyTTGuaYCBMNgV7y1D1lzYUOVVl
zW1yy//H596eUEKM9FgEO9GWzsY65xzOLG6pyMFvaEFN8vF3KbwollPXKaGi3Edc
hb1XSYl0H99nHBHB18/y+ze0SFaGh2WV6zcL2cBsgJUfD0/XoDytIDtSlTLV2nLa
5OnKB12mVTKh9uezOk8pfDHPQLxiRKycqGmzB8C2zAwpC0fxX13oPcXlIWfa2GZg
Af5rqKBTbCZeRtuIv9rwCW38gHS4CwuU9Cr31JkY0DuLWTLD+jOQL32PJNRiqHm/
AoN+gyYdyFfJ6FrMLFil6Gp20U2YF/xwos6S/ZY0dhxdWHdQBMy6Tfn1j/VMB1LV
BriZAkpV+OwWroeMYtiwH5/RmyuxVgYJu+hpi8KbOPSqUtrhUKwzLjf21ope8z9b
lKSIAgdmdNANCgE6uVtpUel+bXh/O8kv/+tGhyeHFa6tS/GWaVD4btwH8VjxMmYj
azYfjOVPOJ9HtuTHDaEdLOiOrF6qwhYCHo0+Nlxqd6TocCucXvgqKvRr7n1Ra1Vn
5k80ckEH/9ajk1sPasQHowumgj8f80bQ8sSL0XFG/j/iEejqUy2eUirKf5zpU2MH
arShXeUa8JQ1DJ5zX1Xqkxz97eXCrccNhk/CWTR6klqXgQ8VR/ngMVk5Ig7j0OeS
rm6RA2jMykXRVCaalKx75O6tYb/my4FtZlbi5GknVesce0cm/CuAanh2Eb29mll5
1YPQS1HqTn0i+1GOcxwD1mRfbS6bHOang2YMweY0/UxMABnOCHOFelaGMURdcm0/
WIuyYrFbpEo4+qgOYAoGDo9DJIkrUTro/kbWfqQXrG+AcLj0o+pbhJXFCbEfbWUg
bYgC7i/rppnx9BGGKC+AowbNt6uy7sl8EqEjO90ZMS2V5jX1SN38S0VwnZYeCM1y
FZ+EGCdBEDGSeQrIDiMif1xtRGUbyDQZFAItj3x1kFSpxg/I2Q6BB1qaO8rQHBRm
fOdF4+7ajvE89DpvhQSk2QsHIcM5MHNEMqopvx0jvih/+N1u2tSr8owpE8WUQgqW
5c90zTJPwLXkQ5Uy9khpdb6dLONbDHNBtSkOAXNBXKEXSoqS5uA1/JxRxJ5Amdr8
9DOITEu2ZhpRPQtUHh5WrQy8yx7kbOKT80de619eQc/xBZp+OxXIhwSzx5FxWLxs
1XoIw4iUQJacxrQCTOeSqgq2HEHxFTtxJwwyCl/kJQog2HOfn++3SZlRoV4bi4pM
u7ku7Ox0GkTI560Jwl3qPeBlu8dM4DYV3aUVasUoaV+fOZpK05iZvGZUPuaCK45H
pSKfcqrJfC+HXr9SNpxIBNshnaqQjJ0g9UB8VGSA2i3elK5u7g67zcX4D8ubZCmS
PviMp/JcNXtxRlzhnlPJkD5snIwzljL0/Ii3C9eCtfwykm/NM3oS5mX3vQC3HT5t
7MCwL9vg1a96OzciNc8tncVYhrHaq+82AKEmNNnAj/OMt5LR68wIfHQyJlEm/S/d
LZUSZiDR67RTesNoQ+gPyFiwccEcN8yHkzSOSkaXJRYSpKjEo7Ouq8pLiWhG41i2
ujkksGHoOB+gy3D4u+g/dNL+szpet2+ViFa4vozcoYI+On8JZtddHoVHJXo9Ihlc
GsOovUzr8zEUTyguIzlPay0VoO3b8Hbjb4AFif84nDV11bAj3JUXEzPaeVK+Ndmb
+WuhmButSfoHq9HwWy/EzPfEnCUAZH9kAE7yO/DZO8hKvbXcXDcvX1g2VLvfMzV6
qOrn/uKMGcYNeL84p47ajNCvuM3BrPn/ud1SO4M8Ohl8rI3GsPQRP+SrKb+tofi3
DSWL6M9QgYKpzchpVQ5dur3CVacbIX4K1OeXXXik+jayz6/5/qYGfvFUK7AJVOql
VEv8uzcSyxo2kADSTiCLEJWY89nAkscTCmttIpS6dKnnMcfem9MGulJy+gEp1p72
u7m+/uBraBOwL+/fNB6ZbCt/U4LlIy1ZmFV2Wj+lbyEC95NaAxpbvOT4lJFBTtyD
x782RgY1gDhFnSo0YTn0OQzkvtr8mtK8BtWGmcOQZJZQqakJi5BM3W+1/rJs2Qou
fvJVifIiazq1TBkbNiAf6kOhToiOtMY8VJOZVsEKSkIpFxU5aLzVRyhcByQv8EEs
D8r3gEFC4q/w5OaTNifEBhR2hP5wuO94ppblUyLq4vXg6ORnvBKCmdV1qkmeg2N3
HrsHH4EJPHBzXepTQ6tJelpnS1JVBXwQOETodUuH1Q5aZrpi4OAJAGUxO6PEDb1X
4OcM+CdDXOs/TbOGDiqAWhHg6jy7RYxbqx88KZEbpozr28d0RUPiRwUxUyym5KAm
xL8pX6Qr9aA1HHGZ6gimQHdMEnXnWf4CRDEKXXkDC/lHN8yDVW4V2sgUYGogaOJG
jE3VsZTFc7XSj7hZvU+EI2mqgB5HDR89pcPsXZLdfV4OM98E4w9QFz0HI8qwC01u
oeABYa0DWbFluborjNZqZTrklB1m+8lFLVfdRCvP4Vxfw5Mr/kjFTNTGt8iRpc8R
3yM2GnrgPaut8MQYlRFqymIRclpQm1GGUrGbWGNuufppUYe7HIrB8f+FVutGjaWy
EVbxm38Sq95m0kreC7iMcQ0vsztKgDQdoWzsTHZrkXyF7TFP2yWxliRl1m0QhhjI
2jt1alG+Ho0FsElhTWkcJQOYIJpgKADabU1lp8xiAlPDSNsYZdFbY6lYxQsNr153
Yy4tcesjeUHfbuEtyq2Q96Jo9TW0oW/+fzHRDGE3EfoWqzpVKXljvxoaU8I4l3NS
QV0XB6RQ/obt/33rRYeD3ZqacfJ/0bSrOgwF74gPvSoKz5YvtlX9mdn26qkwJ8AX
OdeuHZXCVM3k/S3XhmOIv4lY3doL5/0cQu30uOW4Lw4Tz+VPSTnl1qitT1OYg2Lv
TDMzNmUFM+GlLizrGtOMePNWCRErSjnbHbCbe+gblFEwCjzqXA7VyI7+5yTiNCzN
volsLwD+P9vnSqDKTb6lditqK5p9XGZ9RSVTPpbT1JSTnPhQ1759Ydnrx7ZfavG8
iX3e2yvE0QRUhaBJwbi0Y3PoQF61BppDcUUSvLmr3oz1J2mNrM+Xg0zZeuxxkBHT
1YWqqD9tvpUVWo4Ynj1oxL98GUaGoQjULML4wzwNxgVRd900FlxpXIh/uRWW60JO
MwYCTbxrurDOssFSTpIxephH1BDors2h+iwg75iTkPkYTp5k0qAh8mqTnuj8b4ii
WGc+Nz9ukcHyK2H95gERSfwyo1WS7z3Ny8CO8OYpXVWW3R8UWuV2IZtDGeDqoawP
deH1IqCu0wPSJ+3LFb9lXNzMTtFKb0Co9ZxEbTC06siFH4y1mZdVX/RD59TknyUg
mTH7Ga2SgRAbw9cSijirDblorl6hwKQx43IPku5kQFkmKxA9+g+D2ufnu/zEyxO+
F+jyZh9gGohXNgBMZOlttYYVBPycdGPG+qUJzt3m57bAQ8dfG6PQLtnetqP4Yaf7
ex1OVQ/QqYuude5Vj9ISfEhA47N47D9nHP1fWr+bvECG+sRCASPDUsy4dAoJiD/O
bTtFQk7do6a/hEvzjMw3cjtcnOK59FwsySIOZklaxI4KTdFwhi1SPOUN00eG+ijM
fVLfAi7NtFV4/JH125THYmukgJxVyqy8nDV17n3Z6CHv/9IUMqQc3xFHmR/lMgmR
gxlLaWnSeD8ki6hVRAXEKohi/wKqX/hdjKuS1AAL1lEkjuD+Cc6nl61MsHobcHuI
lWQfnF0bXcWN+d6HJjp5alBlyZ/u38jUFhV9PFP1N4557E8g/MlJl0gRS8Xo1pSH
BwH6c0QT5a8z784liWTR931Ogq1a35/AEqiUWBuG13dlDVoQXGl+ewwoFbYiBrvV
9oAWdm7V95ntvULDncsnlA8rPLGP+2NIM1ca9U20YLasnNL2NR7lLVsnOy8FKxDN
qDa7mnEXadF9LQ1jZIy4ImMFfZhgAac3sE702yx2/4XJjWKLaBoN7F2+TCf99tvz
bAbvUJiSHQ+AoqmCdtAG/QeehpKlI0mEa9XJpzlgrBrrxC9nOn5D8k8lvswSsgI3
AmkcPKVdQpwq6eNAY9kWy3Umd9dKev/ddWWUCGbJFqG3FwCLwsVmqE8PIjk01sK3
++lma1bMQskPbpaVe0g+5BZVcWOuTuXcsxXP29jcndpC7izR89WD2UXzQS6KGI60
IZYnYhy/fsfMXEFvhFU0PXY60ZY8yAV/dvG/GGf2fij8ki2aAD5JJQFB84VozkmR
ZwhnoWv6ziYZwxlIhkO2ZcDpdNIOWW+8kKcQgW3RQ4MWPD23Mvm5WFyG/O3CRSqG
1Qkr3Q1QeimDZvMevieh8WyBW7Do+1NpByWGFfKlRAeiO1kbbv0Y4dpZVKMqfBE4
FmPW+x3TK4TWOqXUxviAzqWDwz8SC6OLtyppKhRnIGbUs3uE5oru/qCAlvpUbX4E
RNU2V3Puiaky2IXtGsc5DABvLql8n9ni+Gu5tdKb/3i5DJ+Nv5TBad8f5Jrl2w4l
2CnP+7Lpupc3EcDYd4gadelH/DgaILtotfvkR4p2MWTFmttUDvMPBEb3B8YEVdbM
YCBHinUa99sc/UMv55QMiD3fjEY2OqwRn/2bPMmK3/+kxyJwB2aZh6vCBS/BJfVX
pK3ZPQ9Y7qiIiA7nIKSQLVYYuJ9uciWI9BDV8Tt8BYKjiUR4eeVgltZvluyj5cm7
QZTqkd3X2ZQ1NhvZB3Ia76farQJVMxqIDFOQvr4Ef+L/KvqFC/ygEpeJTHa8IdpS
KQ/un2b6cDWTRKN1o6mm4fGIZ7lQNYoFsRsW4ufTHyUJBvMB+XrY77s4CdSQCWSz
/ikg5B5ShibOCJVL5z7K2j/Ojj66P35CmwAkciFVqOxwmB0nXlUUQPMEqgIb3eo9
NiWxmRRfQ/H7x6+Woa2bFhHQfwyaaGIMsVaLt+62+kjyh/Mx3nlDh0XHXMnoG4sr
MUf9B8XamIMrUhRc5QYPiOgnSskMw5qepQRFAa36ABXScpWO6AbN7E3u4fkJvSbP
8r2kAJHz9Ac+9ogHAL+K7OqIZn4w4gtT8I8EuB9A+4U7Ht0wEn1BkrI5jUsdpShN
8JWDOf0mYh3qA5EAeMnhMpRCxN+PIHowpviZR63b2ogMUOcROG8rYYNCKwkAAqn0
w+bOzoYuNJIdEa87A7MUTTQTtcO8JbNyVdLemb3oGBaWaOb6zmCLheUWCxBnKccS
WqPzmuKzIkvOvLin9GmmSBXKisLT07qACTLB+rVvsh+u/IDuFcbq6kDpZMcDKkHp
JDrF1eOy2XDdHeMCGWHSQpRYr/X3dDMejOSh6N30GvE4RZ2AUxz9wOR8N5dq8ggo
KsENWC9ddND+h9GXUXQGEl81nwhz9fumpO8F3vNGDee3608VDA8Tq/kjd7+g/tJt
oah3Ct+c/nIseQFAy78EWuwx79m6mYtBS/t4gYlyBQKSrpxAV2wMgr+k1QVHGh82
BpRee6QxO36GnJVOvxwXW/MC8GcpOALp5Kjy/kVGN7n/d1gnAKa/FlX2yZY4SWqV
4D1NRlsE6BQwScRcDNyVyeLqbb6e5WJvs960YhhaNIO2qXJb32ZEpx1iWgEFy9P1
ZtAJFhCyHQE0BR5r8+kHdUP61c3K1a8mWXGbp0+fXVw/Xxjd2fbF2pgdRFFSzEpa
77YSTHoaUms4mgHhUWZvOvIWyz3m1/1Fz9e7kKulNPAL+bgqG5Po2VopbHHWMCuq
xCqqZf11R1fq70OuIwkZHe46Tbf7jXSy9edLl9ygZWn6OqG4W7uSrXJFIHyAk/I5
uiwSVf246Q4Ca0Ryuj+7Daq5GBRmEjSp526OZdcNb9XF9A9cU2PPycTmSZ5SV+vC
NuodWFfosmnZbvTf5cImN6n//+xWxgYIBgXo5sMyPM6oCYsPQ7P8cKIN+jkCUv61
njvDDeKMab6ZfZmVf4QOEKDzqodtZf6MamaUkDMqqCcWavKch5eULlqdMGXwMMc4
/ffjkh0FrAVJm/sSZ37+SP9Kg7i6msIoPJ8t6RJFFaWJoPmBbwP1D02VAtMF0X6y
3hRoOyosQqVMbFPJdt4zpiG6+e1I6VBQGvmzUS2bdSmAozo0DRXX2p9Qh1DDPHNR
/UsdtaDcxTJEmsgrDYXsparSulHra33//X6gzlwQaCQz9ePArCn/LG6jvH3wDGZH
crkYKb7izLyMdD/zTtONUlaA/CLUNmkeTYiETcR83n21NHqs8BTrVwd+AUsOFTWN
rbo3EHXHxUexyUnuA68tgxkVx2atlPUTebnqH9brgKZNFT+Cpng3feRyxGGUMODZ
D2lWGMpjOShoddV9B7tUzFRx2JctisNxanQwKJe2BW/x7C6XLseZtH+l31OPJ1JP
2SSSjyLoRjx08QR97Rd+ftQyUeH0vrEOwanzJRVx+Na+qRxqu+Z8AIeHJXg36vy3
Hhpv3ciii4JA6iZLYhR2MVUDDl+Rzvf0XO9cFtyOVYV+nJpA+Cz2Z8PkfL8aVOAU
aqehD4piesUKX6nttzfBJVeAy45EWSfAOb6JxHvZX5yeVqIwlsw6LrUgHURW0R6r
22Fs7T0uUHaJGyqkVk2YmjGonc72weS5qjna8hPU/N/oX38C9e6IIqi2nOUPHztj
XImyufDWeZmmU+Nb706kiSvhPDE3WA1NowkfWNFr8Gtwo8u6FEprPj7G2rtK4YrS
/5Q04vcioC6e44Pc5cARPYN1/L18RDqgjpgKfWnjSIPTHXXToIEByUc14YDd6JYd
7RDA+EUdcTTJxJBpx82VtwVm9lxmuwN/tOw6UM+jtSGDwDGhc0krwZkByUggFkPb
hrzNYEaALuVnnXcG+KU4vP38If4xWvuX/gZmtgBwGuy0Ovz0L01HSAjYXghbSGUI
qcihJWYr2LmyA5BCB9xgykYwawVyKlHvEI/Q/4Uc5MVuhniwsO8qOpEr8lzPHgmI
uxEXhC9R2m8tWtHUxZ1DkNaANRF2hx/CWWd3Lo+VTYPRMp2eSOzWqmiPn3sN+DCe
HfjRA9CRJ/kjreawVGhQ2B1J7UJc9gC7s3ZDnVWgY1FlFsjgzEhXnwAGJpjzs46o
Xbehuu1bkOiEeVLLjj2JHFxupmKP+TVl6X8EaxBX5Jx9pk/6uJTOSSmTWLtobzNG
MJ2eb2DQEaJopIhiiiENbrRfiZXQ7yOH9dG0QesC657k4WmvweHBdJKP31+Whfhu
XaVtseIJHRG3JAHbbMC9Q8JUQROrbeBMGZCKXjfthvi9A7jUtx1lwQwpzlWwKIHm
WkhIFGSK8C8pMB2XNgRP87KlNXG4pfae+GIDODtBuYNHBS+IowyCE51pwJj5FdDF
pmmE4aJRjZ/PDjyRlkdKLxDT8KBYdmq4yHYaMVNshHhsuXxhn0EIsHjD68UXlvWx
OMibZWqcfkgU2j8zFVCPUv8V46qs84sqjzK9fYBgPvgFLHvLJJiOyaQPlRqQfE4P
NrsDSxE9QyQIzeH1ZPL6y+B7LRxXZioQh7rGnNLkVNR3PQH0Uc30CgFCatTMA77M
ZTX9WL7v8TTjIPKGbYboxqU1wqlRPGmPxVDtTe6b/RbslWqWa/QU14yadWuxtOqf
QA5mpZpq0e3osdeAVmwCoLLthhgdTtagVnBz9fCi6L1TMpQmR1oVXPQr59A0Aw9W
G6EKFLRumUjJ2um0JGm5goacxX3LNvxLJepiRKmbNp76lBs0eDXfmqVsdYZIPPwn
mXz3JdHJ0y50sRmLljC7HJ66F0FHEEmsGBigyuE3EUvM5QQtPCGNxgjRqIKOhA4m
nsYhbTugrgR6NvaF2Uu57kFEXIPx/P3/RkrHMYvtoErLmfkOZ+4Qma7QxNJrzfwX
+va8iEjoKbYicyC4Ze+iHTLsDfh9FUBRIyhYnn9ZLiVvPR6BgJ/8sSg+J18ID6K2
8clDLYp5MFwrazaCgbJCuYsbvKjk5e4W8SVNcbcE8uAb5D8t1mNMdGK9DhZuDkIn
O/YZSOsKImfyigfnSZbgBV6nOpmUdgg3treVgaUVV2rSobWSBSfDtUpUHhrkmgGP
hc/946evDJlFpDPWbUo5R3caCy2RgnZLVs8fKDfbFV7fWBdfM1PpLq/ukJqUJFH4
3WwEl9OG8QXiJHo93VS9RVlZyU+FCRRP0oQK8LegrJSsS3A1jRVzISCS5CHhnhA/
9UoCoz6PPWhSb3tafiYv4g8dYPuII7Gkebv1gTiyHrWLZfmjaTrxA4ogs/Pefijf
wMOuk2c0NDB54IORfMcFlgyUKcP4TsM0ddAgm5UupMpXG4+pMe8KvnKQ6DmNeyiH
jSkGYa7tK0Zf6UHvEL2/h+duJ4aqM1hPQe4/Pd8tJCvV61OpVcDx8WZJIpl/jC+x
LZtBYp7yDOprf1MMUdxjP6fTAIPiB+wW45ZIS3q72QGpjaTX52pIikTaMneUszrq
YIoP4HKWGAtMqQC7cQmDe5DdYqJyTJnGv5GLREOpO+sJgH+QK3ACpTYkI/MLmmiZ
aCWe7CXYi9CLSMTSNZKGIKnfb1trMyisEi7xx2u4upw/Jzo0JG9yk8BRMS4P4n/Q
aggcEQvkkJZN/AOgA+ZIUkGtIAIFdYlbymJ7iyHWH0GwY54YSaQnOpUzbjPagkb8
Behd1ED/tfQAgo6RoBqvGByC9BmQrVzqhO0AkNfkdXy1nGdCGFOKHb4ynz8NiC2D
1NiOfr/oyTCWP+FqM9Yoe1K2RK5AGRMFC4uVjWTbUCyvFS8F5tfguhiEJPFkFGwT
+gvXqlgl5B6rFNQc2arCZEg5CptPEPqQv3kxM10VUyc/DnljhBgtcB3SbhachJQ9
XwCjF2glVND87u0Cb2A/Bf53mSAw0DUwQKNH1m554Ii9PZPZ9+eZZit5WBc4F9sX
+9XBGTQll+TQy1MSiZ4uLYtDnSa8D07+glDgnFvtOcNjATjC07V6saraSYzlUPyB
XPQTAhZ0lMLR1dOLO+tlJVdDbmsQiUXb+tjvCatWINT1OJQDXOi6F5DBlSjJpN35
O+j/UX+rfq5olDh60atQQKd2v9IrvfU1msbpltwZUM2GDJh4E4JYn7oncLofcggq
kJPiHbBJYJIuzA4pUFZRJf/c3Xka3Hbr5e8oJOuqVlJTg8GZ+HdF9sgpqpVelWEY
FNdXlrB6ivI723PEMqFBIyA7Np2B/8fxp5X5fOBulESsZ59S8PJ+QQUIuQ9N1wF8
uWw6G6WplMZqOI+7hlRmHdkAtCibq3fRMsYjT/dy5oiweS+dB3CmsUiyahdNHk/l
K7rQUSdPs1bzioO1Pe8sJcAfhoantGNTzUbrBRrIgO+B3akXreVJTliQuHL2A5pi
brDvU8v7YhJLGqPpoCRrHEHujKVqIEOtqo5qNdLrJxm6+dru4LVjE7P+XkRaUYgI
odruuEkFnVnohlogXO6hXeOSH4PL/hzpuarz80hrfHMAtCiSoBJ5C5ywiajg9MUo
aH97LN/GfAPuZX1J7ojFJ0On3rTnP/dTZmPFsGnPm1UUzxLWyit0m2lmEbDNxOSR
gyYB/ysY6Xt1RmDN6nPrMSCKFyyTj853W0e524wlv3CLVnm0GIDzYT57vSmXjv3n
9skdkVNL5TzL+K2o35q2RieBJzQnYpH2/j+BV+5WDUdz2Bpe5EikT41r0ECfVztc
HKDggNfgSAoycSZ8MLUZeCXtFUTMyACjKf1o+tD/ymkr4LthlIc9sSawbi4QbfmM
N3ok3Bbga5rfuwUX7gpFS8HAkfkKW8Pue3TN6RLQiUqFZVv4IsTFJa7G6g0C9/9F
l6czbkBV1SkKa+layExpg1rcSK45KlKwOsv41Zw+j2lbyk8571IN+XFRYwJN/yGp
9RV5i7kgoNSdLZPk2fsE6+w3JBuDh14vEQ2mMT1ZZwZxxEmKZvUUxoMjwMqqeTDy
/1iofUMeabwLolVrAX18uQVC/dbpNZRNf26Qg8CA5hFD3IRTCgX4akvwtEgfs82y
k8SeqqHwF6atX2sBcfnz3X02okNyaULE4LiKkaA3MXbL/765aRzM5J8/PZEK79/a
IapVR6ar5zKFKDnUJnrj82Pu+XhT6ivem+SYz8oTsxUiWybXp9X0B2RTJBPr3dxT
8YbqPT8nbRRY+aixjcxKNB9DcXcfH9LpWwVwmKyNvZahMGsjmKfhSfJ3Zg+2DcAC
hjnBw9qlF3T98VSGf1Tzaf07BTVE5yykWbRRQ0vSUP0KcYLtGVCFLi1zfHzlZW5C
CSIhYwQO7YSu7RBBlJJtrBqyAHTFakM8D9ExxoR3FOAbV9I97TJCWB6QIVnKLzo4
PaEbRzGSYqVHW/duQAoNsGT7OVXP4y/QLKTytaM9QmTQsIglSB4m/anmU9G8FLKR
XQ2AgVFEkIO0BsMZIVSBwW6mIVViELiA/RWAOHpbntDil4+KQASNgwwJQZ96ajYG
o4AO33PbZLfpaCVsifxlblrMaWYWf/TKHRsquoho0U3ExntZBU3Z6t57iD5LfLbU
QxUVloNJPvfS8cKffe9Gy0jiJ7wo/Uwu1qM2fB7sV9XKvTjRbUSl0bU2ADAxYiVq
V5ylo1X1i8VamPxcl9YOXxhkyFNl/17213s4KPrHagw8Mu8x8+dW/IjyAOkFRDUl
P15trOgU+cAZfQWXEPwkIbA19wHWHWz8h+8lkytl9AmIaK6JWiXLkDn150xZ2ZVL
dcpzG+xDE1PRLqbbqrDeipnaOeuTOJ6Itw+aD4Su+I7oXRDHflfzGTCi1WnALiyP
sk718YTvh3nV+RmvYMeW2LBuJKv1eWY6KlQFnu+sc6Nu7g++UcUYdIpMgcDrj5Nu
Mp5ddYgAIAQTHcmjqoaffCOtlocLtzXQ3eXcfzIiOBn4tRjedQEFsm65Z76xdSLw
Pqv8axHcoNUhRx3wZsL0HwJ4Ztb04QL+L097BivXb/3z/gTbwok3e0PBLUbmf51C
rlH2z03nUpvjWze+JwG5TqPX7KoOB4ryyVBb+00gO3aIgBvEy9c2FZGu970rTKMg
l2dDUvXvkIpShZiMWSNFlDrOnUfU8bUEM1HZ4HXxhWoF56ngooCtdnW92bVWoVQq
/PmJ9yLs/6mTer6LkXGD3tKjwGtlNBGDM4DonMMjZc+RwwHNzdnOFil0U7LMVNI3
djIU7FcjNeJqh2v1vuPESoRc6fy4pj9v9e7v86Uh60ZOL3p/Gy8abrBH4IhFcnF6
orwtOjrvXOrLDmcc7ECqLbOigCUOyVy7LMIaBGPuhWRqkh589QFot+KRBjMF1f7l
0LLNuvEPw9KqWvTYS6JWWLi/JJx85XaOjKCaZZ02Mw0Sk2fC2CqdcAvjltZ9l3cx
4lRFLDFaiGW9RDWVr9gDuqYdJjurUVuL+l4G19SXDsmw9LjKVvb8U7JuY+UUQj1H
6NomaGKOhRJwtkUjpTimp1EaOrQpVF8fJPHTkcufQDnr4zc5Jh/y5j+2XXU5HorC
EuSiKy9w5lN/AFHhvvao1SGUrjAROz9Mq+Rj7pKiSswT8mHHSKUsuHx9qUEfK59X
mcblBdDKMtiYC5lDu5asMmAPky6C+NnMMJK8AhoB3LdY2F69M7oyVsrduFC9MZwl
ZFVQ0S03qGMcXyG5Jk9fhesNPrfFS298lV/E+bV9o0ojlWTSooXLUCi9ezs25caQ
NYlaaTBv9F3Lh7PTTYhiWedgvCPZSxAViKAdvNdKCxDBkxFfBdu4/5FhtD93aBFf
EdBHspxLXfMNdQ2v/qSmIyZTTGzyXDZraWnL51RxBVgTpVEFZZgZt4r2Wr6/aE3J
5BMbDo/+gE01F/Sx3kDYyBHoPIwJ6kZwQnvTLSx/oMQQb0syg62QyKPd3BHVlvQE
Un2Oggi7B3K5Gq4BcH1aIOLwnYV106Y8RibVK75tbvuMUhyiaEb+KXBHSb5N+8V6
BhoqCcbgyzG0vtPt9roKOqBYQ+9rHG08vx5c33Qfzr4DpOgUNeztWDkoGHd7Uobo
Bl7Xlbi936BIFkuWrJybGs4YHZdlWygK5Ehc/XU/fnONgK6GWc0G4CFBndOLIWeX
Nk9ZY8WNow4g6r/5qrI+bA7pPrYPxKHisne7SIZloMEop3ZAtFjC5sCHdChFxqNG
W4TcVdxmtgNUbm1ZN3bf8O+8eTJCrA995vkVowZKwWi0gsJqZd2AOkGI8VFQ9IWq
CWSkj7P4vMvX4Fr3oQlh5sDnIf6aUNCQmYpGHZwixIotccshiNCPhFtHOg+v14sM
7DDZ/kuFKr56aROSIRMfWvF0al8gBcPl6BsprpvqqpCIYerbIW/E/boXQVXzX7AZ
cUHjFK0NpSak4nxe+AZ2n0ZC0VtTFh16tGrmYkbNKmryD/RZ65Cnkmp4KRKihImb
L0toCRP12JjqWasIMWf+8ji63Xbr3ezJW1sHqMb94Jj9yo1pOF7g/FedoAdpoAmJ
iF883qgBziQRLVI5KBtj/1Ad6n3Ulc/gV6ioIaKJGNpy/K/6hH0T8alBXP34D5Ma
aTMiJBC1VD5rGVxSr9JuSPXROI6cpAxylPQyTBXDzu8cQLYqnbW3RMdR4GZ0vYC/
XD8SGAuJIqwUBiUe13pwirGPuRkSB0ZI0AQZdBUSfuy9hAcnEPTKDvGtR3KuVo1r
bse5oIuCU7DcTF8MHNgwLvuCXKwMyna/TlAHJEnKTdLzfEr7Nqdz9b4Bw8EoISsC
7SwBE4t484eNtjzE+IlNZmJlA2W0c9+J0yvH26nEPXb+32noNyGaUEr6wfgw0R0s
mVwxMLBVkXzYMGTL6FyTy6qddR3wbaaTo/gvwrBW0YN/4+gefjXirwfkBDQhe2GS
H2Jg+lEUftje1ydwGNjmb93dCTwnv+F6jkRpKXqWvrL2fSp6CU3sLKn8mvZ5tCU7
c9TbFq4adwZt1UIgyLbUPOkjAA1OD3lmlJNxX40Dtv0cUEDw8FPG3dE38n7Lp8xY
1C+jnkVMVoh0FIqlUAVyPCiZOLs2hF2xXjm4dw/732s9JBqUADAr7gqVhFfUb1FN
ggPykyyjx7PxDqLm8UA0DZr5mKv6y54D8drToTB1EE8Oky77UFu8kOISvxVAXCAO
E+EoqpA95F67F8VpWN76Y/ztFjNSCnXmIib4zKZV8Z4sl1sebIS3HRPJYd40P09U
SOPTPeRMbaOWfJzNq9vBnrqdkDCdubT0bVVkk2uvig/MqZUBgPNNqllFxC88POYW
8dq5xbc4CQN9Kh5s/m47F2ZJPqBre4STxCf5X+bZC7itJn9nijGtYrJj6IJoF3CF
w2kRBAPLVpU4FFVo38+U8nOmn6XbKluz0N/zSIC2iyCE9+0qL4+/Dy2OPQcoWZVE
GzaoQAMs+9yc4/USiljWHeFW04EQ+dKs/dOvSAVixYaHACnLJ4RjuJeGrQsxffdx
AmSRPj/4HB+0cBUCrhUkhzaqo5gXWwCYwkQbTDrjquR28ZxBz3AeBjtQ65zxZS+e
vHLx+iewWqADFRU1R7DpTr9vCy1p/cg29pVnKnGs4sspBGtFeM0PIzaGNEuj6wSB
kX0nEQo8ArEJ1wfW4d+o7HhpPzQjliJdboCMqKv/OdN65AQoZI5arPOw7coKtolG
iYbkv6Js557j1JxJPCgNJxKTD1kbri5xNI4RGnV8kicTfyiJaWag+YNAPCytW+xC
lyvSKYpY/LMVEFTwYwXgqquOto2zXinVa0/CeiGUXhssPwwY/Y4ByIYOkFWIKWL7
4SqzkGtLuaShZw9jSZCAeqLeNXWt7wE1iS8veOhevh9gZzjD949IwRQfevV40lAj
YzuKJwC2xkSfxIxTlyNaAMPCGUDi5XYwY/bAr/qKDdsbX0biNCwS4xzZClSCUPnD
zubMSYGgAZalqtMrLvglu0W95zAJ+W9xjsp/ytWGLIuHFGvlbnGHcv/PErOd7mi9
nKSEu6PUk+ePmb5sptdKJf4Taow0Xo9muJRo5CYQBIML8zhUYhtceXAI/pj4aV1r
jZSi5Hd2etKY/JVWdyIq6+iPuVa19HDBRYsLZiKQVEoppdlRz87aUThcUbmMdd+8
fIztTnkkS5sAtT+v15EzN00hRp3mgisreSJTt2UY/yWeEq1A+L6hWpmq0zogi9Kb
DLNSS3TC9VIqygsRZ/nQFBU5R/OE5WYU8cy9BoX3g75M4/RNKscee/ei6c+37a4R
k0Dh8mUPwWv7zlHrYUosjtCJavW4pUcwjxV0TqPgsIFZUyjYCOfKoWSFMeKk/w6Q
ZWQUU0RjdoI4Pa2jZ/VCw3BhxJF1YiORPWEdyR1My/jWzqXdbgwKqwrmvM90+BHM
MIM6VUkrNoSbmIh/cciwIHxMASXV4rjRQ7c4m6RTdXKnLdsL5vV6gn/S2P1CtaaF
0AOsZjIlThUESbLtOnSBlAKQQ+zWEVTtnCPmLgnDDcpADt90A3NTJyUKGES+5bKm
o/HKYIT4pYnX0Z5YmHjQyZFWFyMwEe97GeFh5x5D7I2eTNYB2tuicEFViptj67yb
MXeLE7gWdEmm/ziJWmP3GZmFwMofTLZElpAUv91zZ3H+j28HpN9pLjZi7N4JJ9tv
NpFP7/+KNaSJPVJSQzdgbnUICd1eju5lYyn2ShGHBDTzmepgno+A6BEGR/UHZWKe
oik6kOTq2Ztgo1yOXPKLKnRCVLIuXqAtQ3XKB+cuCAzFIcXM2HbbsL3QZU9/LCkU
ZtKmLykTpSLGPCQUkz1gVIe3T0oZ8TZAsB2Os8K0w0BIeOmEbWYremPZZttEdCw1
6GgQClB6xmwqu42sIS/zsl4x9A6NFMrvL+y7xgp1PYNOjGuqQG3rlsze9/LjmQN9
nC+uzwuzpHGCYICt+scmCbk/X9lXdjd1TW4Kl9UuqeGqqM+61lUcSG7CdNxPtrsK
SfL/oon1OlW+wslI76YVtkYfKWRU2geZAZirA5emMDMLr49L2ISfigHjTZAXSP2l
CJsebqg3ZaUY6xMqnsnhr+jL/STHFBuBq+QE0Cpt1KgpAwHvTOU8HDf45fFKwO5O
F8PIN1wTSNJG0h+sCYlh7C6J8ykC4gYFlNPD6clh3ptiJgCXfjWbpaUpo3u7aEK6
3bfVg2NgE5jVMYFGOofQhukYMA2pQsaTx9uAYYtnG1q3FlQysBveZbyULZ2ix/RB
0KzSiaJteP9Ng1VVEUBsci5vdO8ISDe9sW2MsDpCz6U/ywYAfBGkK285dqSlSyb4
Essl2CPqVJAZu1NbmtpKtb6Wbk/A+4nHVxkkesC4eas55QHGVtOZBewwowHbhP0r
GDPUU9f+6KBazqa1tz9JcyKSKuxLnC+MsFq3jDnpZnG/4/mkL9o6Z/oc6L72IXk2
+ktyUZBAAIlVHHGn/xgV72XxqlC9vmehkZuJ5IW/8oVOItLAmOZUGphgZuiu7rwI
4OP3utZ/SKuxkEq42BEAQZQwINml7T/p2i+vyOfd5mEyr+wgtw5OBqk3/VCi86Ka
hnNlx4AYJxVigRjFy1L8riZWYHq4vy2RX62ki4ouRrWRB/V7VhAkpJ+gcuRlIvBw
s5sq/XGcS1SRMgxbB3KA9E+Xuvp+IuxnEPQqulkHjLDJo5eNEddB4IzwkdA09+jg
JBOIq/p6a69/7XjIWQV1dJfORjfggdTmMyoZRdeNzOiioivMx9H+2bDnYNw7E/ag
PXp+fWPhw+ai7oGQ8VAuq3F0vXzb9BZ3keLMDRK1Blm+UqUZMhRLZtwTInpJsCjd
ni4HEC1p/4f/vpdzFuNYxFwRJp1bkiSj0D+dmBMooG7C8sWIujxq+2rZERLjgZ8X
EpAiRfzASWYk+LykmCvEgVZEkn9XqRiuGjy1TsgKU0vmtBxgAhYYsi1zzZILlmug
tv/WmgZmbnQzxcOqdNpORW1ma3zv6r+P2oqquhUPs82E1tmT7kzsKy9bQSLXpysQ
I+NJd4i1DFgXVwKa1ar7CjCuCzt1SmxfATCGDld516bJK/5dXIRLaDYJInCkLt71
XSMqF6NmXPSg52y7FRMFHq6LtCUhSCSJrGOIBvQzVXWYqPMm/XgiRLAwRhzAXmA2
6z+mTtJJmQcezRcixaerbubt4IMrazxIoYyrIo5ujNIMPU+S9A7z6y9blNNOi8WN
I/uLY8Th5XcfxrStk+1NYRBH/WqwdbJIi83eDLMblXQZWQxfLJ/89N+S27/94ZXU
98PwHxyi8LaUJVRiVvt2wkwts2bVVgQrCE/UAnMJBmCyeonVOnc+O4ParHAwQRTY
SdIaiP1jQDJEQhDDYXvl0gnib7JFwwH+12lfMx9EMn2yR1J2eGPZ3pdDTHdKD6gV
QR5O6LS3+s4LO88yGIwnEudJ/PeboX59825GwVH01wOjZ9efH4HesxstjV0OUsNw
iZK2po8OwhR/3GKiMILVXilCHhl8eMzy0tQHN8V9hTdrCyCVQ2OYg5mS9BVXCdwD
p2If9xja+tJPes0MsXVc/BZG1O2X/5voOyitGccwZsN7tfe8U4FvMzA1vf/hfWyi
Ggke1J0DoPKYdOmza94NyeYzEjWErGd3G3oL/6vn2mab0DF4Yk70J5BGq1lbesi/
WzM8bVBd8NiVn97HXo00JY8eTH50QxnsEqD7doGsm7pIbXZCfRbeQ9bE9OQVxLm1
wJtixrEBICL+vmpBy9r5um1Q5Nl0dfE2DsY3OU00ey7OItL+ju8OFDY867n3ZFKC
tFbkeKfpt4/i+E6pIrhziVBk/o+6UZzpSwXOWOn24xoybWd2hxqQHC+WZvW0eda6
G5Kh+T+caiftU5Qpvz2VO2Ykq63ea0ZdLVnshcWU+9iQ02w71Br34zf+ugYEdDja
YphxpQcCKwsPH5UT19JAqb/H0vjc/+BREvZ9uehx6uNHJtmW5leF4NqC0y8Aa0T7
/J8EqhBsaz18p235avrOjKe9U+gV5Ue7CcovsabGRbApQVpf7tst5ARyBYBEs92b
t44lbqXDfW2BLOSUB2suZzSBEnpnpAcZ7G4i4DHaSrCPI8ll8jVEDmtfzOkHWaxu
kDlse7CbWGUSA+SGPQSy5+I5GwtjWRnUS5JvbXwkJnMV8Yd+Dd9Xl14dcx4Qx0Rv
UiOuC1pfFBGy3BxrY1RSfbiox6YUqMOIFBDt03pu98r19vHw7Rc9+QH6gFpjAtX5
RLKCcOWb6Ts89ZcaFjOfHaEVRq6NrC10Xv54yYmzhIrU0w9ED7Vb8al4/BqwXbNZ
J1fmr/ONSmBLwradgqKekfgc9va36oa7ehrzkf79CLn/ikSOaqqXh/fyAvBJnUtA
GjI2CHZmDO/Spi++L1BPDk5KcD1K0jdKkRkuhVkqnABZDv7BgILczSvqYUii3/Ky
ADeI0kAPIS1K+UI1bnNp8L6zj2wVxP7+7sA/yzllTXlR6lgHZGPliBgde8qXyyIq
SlwM9Byn43wwcTeFRsrDLohsKQAemPFbt1mqyRzEXyo/GW21cIu78dsZDDjDqpR1
fpTdK4cPpN3KJnfR80Zm4RfrflH/LQbbXQWaHfZJGDjkrU8qbYTa87Ui3VmLW3K2
LsQhozCwmNsOaS1xbKiyha5nQnMI6DGjARrjoAtLqZ1Qi6XCUfDV0JtSucITMOzK
gERJKtfL6PAry8GPtz+oYNN4MLIT0qIBOgn1V32l4wxemuMnoOVHg9/QsflFBcgc
JQ626xQSIYku+Wvmgw8E+1QAxUd4VjdKyAFoPMHvKCt04Aqmr9wJyOq9BGTEMlYs
HNdyzww3vpfePM0kfYXvuxmP9Susb51g8RHxkofhzlN4uVT40izF6iukeZie1Gcl
WltKr6EtdIatDx61S0WMESbRXY332nLol71y5PSHtr1e5RcYkfhS/WQk9iTdtAkr
MqVB7nRZjTOOMWGcXUsEmGrHrKTn7XCczJQbLc1XU5mQro/IS9rwX2TnK0fa6oWb
AvxZerkxikxRCjxWpZPqqAqMYaqRzWzEFc6Bro7ifRaNv3dCleEO1zID68/cEmWS
c/oQlTSlHrw6NGxaSVHFLLHt4zwfYie1oxKgzuM1SqcHZYsaVBK+31jZTMM2EZs2
YtGUChQKymGkN1OPJ+k7cGExICEqvW6o6J2Qq7MwcMbBvEwELqPrE0umgQx3km5N
rkp8JTWSWi4dTKK6QH7Z9wjEtzN0UHnMygIJY8hHHaeVO9PIwr7lnfkuHsh8fkE+
UcvULVSBqjwLQhPJel1YTsRig41onJrAkCBIaZHxTM8UX7vCIjVF/89h8vJ9x/XJ
mNtAqIQCuoswWzxa3hYNLxwZh5RRAlYXN7ME9CxBb9lDrtX08EZGZ99vJ/p+IQaM
ZKFRH/tV8Uc4HFzHJWDaS/FtZTjedvXrPBsRpMYDtvkl/b8esSG/tNBw1qJQB8BY
RA/fZtDsxC7E+WUWA8QPm+ZnO4gcE5aIBXWAjuToqcBrU7Jh1tKfsAFB1p4x1nn9
ePAb4/QDP3/jCAV8iUZkK7Vw0I+Du4+yYVsPBwOPbb5f/8+Ia7MbWqJK/lGiHC1f
SWImxUleh4zsWGOcFPaYLb+DTQScAfP+gcj/j17hDZVibvo7qDo9PMRM7YEXOzxa
+T7WJWtMYDWBw6G090o85yEJIZWTn9tP8N6zmLuPQ3yDKOSsAfZU11VV3WsZLBXX
G+/BG68+qHkV7RRLMlQ/bZBBvPeS2hELUgJD4z21SAlN9H3UsHEVR333gAX42utF
JeMmnoR1FVYrj44uQYBI1U+YlnGaHwAI5/rmHuVhlN0VfMDMmPmZOyTGb34U2AEn
HLMavcikF17tAN0MISZj6Es3pdWmMZhuFGhCQQn1+Jc20zB6RqKGxjXfDfBRR9lt
+axTMylCuPvaM6PpJrg/8Fm8rkOZfp5dwk+mBjt6iVyJjaqfe/7aIsmqoeonkbtH
9X16Em0z8vbWNzJznysjbEQf706RtFb1Di1aPQDNa62f1Q97xpCgGTlk9M7Kh6st
Hs3Aw9pj+e6Q/WbM6duJUtamfO7AWWsNa/54PKjIXMmqUDhfz7/m3nJsIethzymj
UpfVhu8uwt5lbgKYCmYMBk39agr0/ePCsqo/z7Ds5OM+e6WejQe3QJCmdPJasKCA
spPSCyLj+3PYO3t8D8b40qs3ij1hQ16d3jiSXGewpZXnBcSMARXwqccst3gnG7Yk
ij3vVk50GCEYTvdcixgH91Gxbgc6xyJAitwpCw20P+B7OcjhR/4UQsIuWZdCTJK0
p00DzGhG+mP0Fz+cUiOdbfxAVhUZt9NwsLbgn5bAmA4JYeofR3hZru3JNE9Luqi2
kQb38J5eNwIM1kVfuCdC11LPQmgHEsBrh38GFKWXy+B7fy+9qxa3KMj/Q1Y6vqwD
QVOZiuoZzuOcs9FwvRO8PICUg6sdetZH17FpJ7AgrE6K6J53MDDfjRbDMBJM/sFm
4m6tMbdwJgo7c3K6Uzf5xwq9gdGJYlM7s16BuO6rACZAnvm2pwqhcjZurqHz62sR
E/agnRy6zNiHNuFFR2C9ml9KwJR1fRzoi/HmgNY11mnDy3ObVJQ4TS1BjkEcdl8C
suQTnaJQJBbxwiHGc+6J8HfurtGrho7S3P8MMGjEj7LCLciyQ4fm0Ee6AStGmPhm
mGvOTM5lSO9X2b1GjP4kRAioglLqPD3G5ayJWLzAsKRN/fYtX4p+iTenhEGcRtBf
rbxurUqIUKBiamo26QEl/gTEbFrx4e5Z3WEJTm4unsiV8fDw5J5LKo2jozwAFiuJ
CY9WQDTFFDfcSd88ML1geDyDT4aXpx9rm53RefP1moECd3Ohh01ls3XujOgCNPIu
KhvteemtPF+gVBMKl2Ux5NL+VcTAcOs1py/XfU+mETssktsVhBdJgH7Dj0FAuhmy
Oyyu5uVOPKpTYsIigR6zeehRdl1u3hLnpE/QOKOwM41kpubMhlpsQ8qAwUTyBUz9
5bjHCHHrNk+BKKI08Vdgxjxyv/8zpA6jMWoFMIuhz2qvv9ouSQzhsUPr+CTtN1VE
ERgt1VvzQDz4qMro34+c5ZPW4lG80weDijdSzbW6zM605yFukt569r2Y5BeHERRv
g6bbgcyaMgO8T16x1lGcouBdXsCK9XWhBHju0DUEJTVxAeHND26KWafoJZzHQ5yl
tF3h6gUfy5scU+hUY0nGmO3ErMZIGYiuzsKuKLk5Zrl7WCCgjYFqZrqzM/xjEdV5
aF7Ob7DIqYSNxfQaJQj7a9zwuWY3dM1QF0VV6vqvehecCPIqgrrGvcSDllsMooEF
IvS1wTVOubpGSTeMOAKY9xsJvYqw2jx0xsFsCiTVKZxsJwjTTQI5qgoks5ycRqIZ
CbyqxFT0t8jLRMw2qnd9GqoGXLzBVIBp5MR6cxe56H7bbG5OlYoZ/6U4xg61YC77
UpulUrRrEmGnU6k6QATXvrKwbwM3xB9mFT41hB/iAvR2OpWSeU1cMlC7G+73NGi0
NYMnsS53udZUxmbXjtKLFGfOuvqSqX/z1y/QYv8IFQHtRkydRvLNBSjyugJ7cC4z
ZBkyXWvfyHJgs5CEba4A+6bEb3oL3QhHCz2cYA+8QzMO/fcE3dxPLqBfXyNNMpuK
pF+7L5CARd5nej/k3rAHLeTtCtJ+ydppc+YbMEZL+GRhAVbiRsLJKl/rP/QZCdRM
DT3pNgcMexA/Ve6ZaMHhyne83fpJZsEJUx3z4hETjIJ9NWrFXgeW/xjNmgNuOXW1
79RWz8jES+WqKNW6CRcORSXuMFHMSPOScq8VTOHgr2tay+RqvMjRcfZxkN8IMiBm
cguRMvqlkWq/uutpmFsagx9+Lx96ZW4evXR9Is7LWNnnycFILdqqRVJrWwfNUeyp
uwN+jUSd0el00RQNKXXTGXcge3nVy4q20dDzTAhQsa6sphUyepMpp8epsYpNq8O0
nYnGEUbiCB18kP/s8MrjPq92gIigqwokiDwtvX69u6KahXRHc4x8xcxXhC8xMTBr
v+RLXJtkYhQx6jSRtVABDnZ3wrou9mNTgCmhCxfGomTEpVY2pzMvLZ3Z+7wDuW5E
s+ggAwJjr0i/C5yiYzTRIqDgpY/SS03XbR/fIdNVhmQJTlshan2cSs2Z9dCSq5MI
R1zUkzI3R6cZD9WtmdPGNg863W16teUGpk4LZKq+pi+GV8pX8I+OszbhiyDh6u1/
+xvaaQ0+0Hhrh7yw2zQO+8fqlijTdGOO1H2RvvSUyMtEYcR4N9DBrb1Z+fk3LPB+
/ApMhTGb+XWjKgxSn0amI1z6b8tb9p/6Uwc5/RGMDF7DlNIOM4yUM8WviUmzgTpy
1jxqMi5vFtP79muTPQ4Lg/a07z8hjEVFVqLxZhhF4pxPypl1ciSZbJafhLu/Hyrb
v01055zkjI1oZxLfKLv2gSMBHPTboPylHzXsqv7wLsADajm4lr+GUENAH11LPUo0
QM9wB4KgQvRt7luS1EWWY92DYIi7fohP/J2duc89+thCEgsCR5SttfAs9F2qUZUN
b15slS+1DdgEMH1J9QGN/qKsx0X+yigYCHRJW/qaS1sAcZ9i9IktIUXLYIacHkub
l4inNbg6LHY7ekMNaecZ4bR2V0+HR4tMClQ6WZxcfdsD/hXmLZ6/+x+PhmHGvy4a
Kg8yAfb659fVE1WkE5KtorjXcnA6KglZ0/h0iLQmm7Daqy1jYVlAtAqrIP41XPND
2otngo+7Gxj45bjQ7YmNLB/YJvmNteX+sS6QfXmsrhCqB3hyRhhL/CxkOd0NWgk1
TUxtDYKUnN1Z87cwkgOsQ1AF5JGNxM+Vm3iBjGnIXLW1qwnWnDWfBEnrn9EX2iJ8
g7zkDY+j/opyuIsInD79Ch/MK+p3UBxtXipvjqd8sDdzbi21E8t1JPd8W4Oapgqc
nRCLeOVLc7DENegnw1EJ0yBmkQUl/JUeaJU6zD90cAepCVkHMr/yqoaIG5u02vmc
Ybn+tf48iMkNCEvs2RZ+/qCBuxgUlCSBvaTItNOTifb9tqnSfsDOCSOhbXv3LsWl
rCHs6uEtktJ4RlWhpmosMzGQ8vjpcr8S7QyEjHnA/ZwoVSTLArY0N8s6JBJv7bno
cSc1sesWyfNqdQfrkbX3guUM242il/9Rp+5sSj1Q3tJl3j2fLmVU2+/jTP7CVhQc
KvlVMUYuchC9A3WlKqOSFA2QXHfFnQtOJIVKTYY2zSWdb6lCyDMYAc9n/iVUFbGp
zsNtQAfiCC9P2ySDZTZvivzkl6DMKyTofL8W3lemg6jxFSvauZr1BW4wQv00aDCn
Nx3oD4yXHW9ARlM3HX8VLAZjaXJ2s+GuAs1YQNq20T9MtyumgsTYkoBuX+CIMxnZ
garNC59dj2TjsS2pGpSvLc6dlMWE2D7BbP2sjRinQ13WF+C0wDx2ok14fkxnoA5M
uiexn3+2h6MPXUj3FlH2i0kIFRO3AcTYMuh72YYWFIOpYWE/4CPOxlbUaaEmGr6u
XKRoCpj4xXBIRfNYIEnAx2kvhuaZZEerm8rHh5OhzXweqhXEX8jfHSqwQViBge92
3RKA05xpde06WI5dZyQqHjUzHFnRUvGUbn1CgWr+XkGA2vFf5RNYRcB9edhPkoGl
XSWM/UOihmW8qSdJg5UDA9QslyRSSZQ5LMVOOTvgSCq9bFWUxb+EoBePs9G9+wKh
V7Yl5GC9OVKa0LQOTVVW+xM7a6/As7RWxxNK+ZyeWj7u+d4Req7bbzLWvTMcwCJt
oAfrbL2XpObvLx1X+il48sBH7QDqhCYfr3ejBogymRFH094ZK+p9c7Jyl7eJPYoe
NGKnW1AmE5TgITd98H9Kg/1/k0A1wWw7/+HFAM3gxCxkMdshszJknBmYi2LGqyOX
g0uGqAfhgazorXFeRQSP7TSVOj575+VMjNmZladnKRNKNGfZlrH+fgeGwPdfs5Ui
VokPaIozYGuu3MkYAMswNkOhI+R22G/IzmQsLFIt5pCzR3jLWrUd4Ho+o0JiExGC
mcp5R12xd7W3G/E7Sscz1n2DBkXYdbTcqYMaWIkBijIY9yXP3QANe4pJXHt2XvDh
8gW9rJdCHbjFprJTYWMqKYOvMI4NWIMIoWxHfP+ik3t262hfhRBYnIVfRMTRdPYR
qVIqN5o4ZPQ1SnXuQqMOatHe5p2l/3IAfCug3ffaV4vvtPcqRc5EZ/j4nQUy1rJD
y6EVp26ECpSn6erAunv/uMH8bMTPgrB4U02R0Q4aeHHEoB1orkZxsJWrljGZbAx5
Uc/EiOiU/hBl/9+qEgM/72ObGnvTgCvSU2RujozPjHv09SdKJh8QnhmxVA6ECcb0
pBYX0fniYcDHxJQ6oWQtIB+gcJNvC3qREKN24Kauvb4Sekz/3wPOcUjanIhD+OCv
jl2qoSu26AuFqOhGmwP/J8T5P5U8xw4/VtghCs0FwiF8EGkIN7OjggXqgFQhajV6
hBlzA4mGH5VDT+RBTRC/t+plvNVrqonMQIqcib4aLru4dryGNms4CUUvJho0xI/i
0wrT9BQATYs4kyvog30VQtYMgazfSrCUem6/4Cs5OOj5Rda1wf9URC1n8i95Fw+Y
DWl3UFh7Stm0p+kClJCbw99bXyGI9Js3H7LDxFVmXvf7OXhNds7djzkdzELIyK/t
H8G6VmuUPizov+p9uHYRII0H0Any6Syyrkgmb0vBYVvr88iWKbERMh/1PdNgIC0V
0FlIHNvY7B3oup3DQWiQWWY58Vr1pMDfwZgD5AmeDI7F9EICWJA4dsCXENrKaR84
9bQ5+mLvSGIgAgMbIupKw/a2jtbSxlQmxrpLW+5417E8ySIPe7fLW18kb3jHHZdq
ElQhWSj+ISuA6VkKtTej2dKnYCNKGHIJ5NDme1SdOvYR+ySd9ELWclYnAj6nWK1V
NwcGe2r0dYs8ZZcYyh70HXjL6KOI3uNdZWYiVX9WKWOQgaHWS/DYdRindDqTftFA
aJEDk0u4wmlKt5ZgPGyATgh8rqNEl/l9mmTpClBwX1HIQxjWPSzY0Fpid78G/KLr
9OO3KvCbwWoapNyxbsvZlNyClRYUvjknFJhCN62ffY5GfAP7bO/KcarvC8/KGo43
K1DAi8LJF0bw2WE5rCLc+fL7y4CuuOz9oviCqFwWfCmOK6ybaG3/Hvw359sYahCB
t2VU4/74uSapze7B5HD7Uwnb8cf8+rW8lm8Mo82g4B8mjcQvLD8xxAEge3HP+Bjm
jY09iFf2x/J7gzJbnyaDV8mYrMjr0kHEKVjPVlgK7sV+J2hJoJ4NM2ocSygoem3u
YIqkljkmUn/AHjdT15i4p2XZjIvsQDLDAUlj7ScYeFyKs1FFDv/wCmjlIK6GvNnD
QjsHoC+Ce0GDoGeKHcFBqSJMyt35tIfTR7k3qI7CL6GdUghaO1K+/Od23D2xYx/N
Mt5v3x0l4pEauekU2QdeA+poKQ6QQqqnI/RlPB2e3Cw5JYLEd44BL6YtHqrINY74
kz42lnCbC/UP+nchTx/0of1NSww2lMJYbc8Y3xafVW67A301GXxN4v3NQWvYHTTT
s/nQnd96BfB3mWTWEgff/0LG2xVWlP5juAVbyNPumjZ8Mr/+0tA9OlMEQ9OQIMA2
f7wyAnVCsPMnqCt+zv7gKgV0HZ1L7Qu0ZLpzBCkrJ4ppTO3ZgiKhp1mGpR8shwWs
lWrSrcGD7QA7VG4zFSRkh1OMGP6ofnTVZL2v+gXxK21VWsNH/OzzvOOyK/HyKOOx
vnvIujoRJFTR1rPrPX/GAGu4bKBX+STmC9ZNIGJW9Ivzu+5YkMdEnkDrnJUXCqIs
RLSfSM/kB5GKmP7cCg2lnbKIDrG0zswTMS31EY6sJ0qSj4s1xwy2r0sDWfZ+sY2i
teCLOYwTKzUbkI9eFSn1DPZmIIk2Kw0FYOIhUuZugc+wn1qwRVx7+GgXbZH0fH/l
MTDtOWd3RYAyNWk13slrdoSwRi7Ws/eim+k3P8e5R2EmRcrH3HsTdNHvQdGbzcui
ak768Qj5/nvioZrSdUJ1t9D/azmliK1qdXIOpPmGf0Qpcd/sfyNPknh+dmnSy5Cf
XplI1VMjZvG1VvjxXWS5KEuZ9fhZ2/oIzu5R9F9nROvAd97f6BcSB3YIkgWLD55u
LZFn9M7gcFrAzJjTJ05RvoKEZI8gv4OXx+1DQIu7U5WCklveIFGIkdRcd2WB5Mes
HJCjUpY+jKUi+B2NP5Cf0KA0Rt/U9wENZzqFVW7V1nJf47Zg4ltaYtLx4dN2o6ZA
DI3QWyt2rRuCo43LrDZp4cEbB2nwBlUO9YtjlbXD3CTMbq5w/I+JZG3b1Oiv3VAY
sOqxAufKOEFIupIAv212JH42zEWoPZG+O6fBF7/rBVpBuwReZgSM3AFycH77TldY
BWyeh+Psg2dDTO8lOcddsfxF62m6/bC5Wl9i2dg3n4YDR82xa/BB+UegcQyEHbCY
lC5iQJRKySvqvF4WCbm/pu7vKeAedcvciKdUEbiLX9O/hBcYUxYZpRu3UN1jPfCR
1d5eK+PTs/fJUlnj8cZuwIc3j5YWGRjPW1NvDCkdDbChANiA7YTWeaARYv6mRX3X
XqhpM6Ce2KC8aS2I6/9dS6oUI5p1UaZA0LX7oZuRfbJr1IG4H08GbuCo+dSW40i5
bW+CqBZMIx24nsXr5AkA6CHd0fAnUCN5KR3kxl70oVHPDZGR5in0K7KyuTa86V+Y
r61VJu6MQhVaSH2nXsKXKZC2m6eCHo/4ZAUjFyM5OX3inzkpo0AeAH/e0SH1KYTs
19m0d7//FFR6PMYDf/CL7Hx5imFHby7dzHKpLjrGIHnOGBRyadRTxikaI7RPnFSe
Pt9KUSBSxNR4DFTSkPQmwp78C+X+RLDNWb+h1uEDch+MJgb2pE+B2/TXdDxOyQ3i
lFG+hN56drSCZMwLdW8+jarn862QhF6nJtEVzKFIV+vgHgMtveIWq4Qp9EDZIRHl
Qnq5KB0WWP6ZqWXOnUGB2WsU8McS4y6rSFfzbzyWTwMfIHG2gsx4/sVNdesmXnXT
FcRhzoHYUfBheWUCTbyy78ZfV4V+BC3HQKhjX/mW5OgFmmWV3DLLmVsodhMz/ax+
ljxfIOC8pOU6CmlmTrhl5EggJlXcuv2REhCdqHreDceN26eD3iC4BUqC7+wP6i7h
p07J+WBJF5vbfwN76v58CLiRtm7PHZhjwpdRpNf6BLYmGVxoyK7sjsaIo0wVWyb5
y903OA9klzLIKMiLA3NMqGhCYP7m9lqrdLXl5zt3Pe6lKNRDe/dVLr7NuDV2T+Bl
2cB1Rasl/zj11p7n5IegC5ObRkUkC6ida3epRhEyt8mko8XzhyZD4Wt/S6Z69Mee
mf7gxoeoYDr6UihU1SdDRrIqeJH9SJCgoJdmgOIOw7jHdBVVkt267bfUodEWyXti
ZpUG32koOsE+MSA1LZKxiqVG085UukIYd+16w2fHKdF+72zWN++T0N1BoPAktjgr
0AJ6c0LU3o+5eN6ksMuwkvujA/PdEkMKvP/BKtodFpY1EOa9VtCUELVwFTkquLjN
OZW9qzOXpQE/Ka3iXBDsPrYTXH89FgWNRH4RVOm57OMH1iu4NflOl2td7lNiP9IH
eRJEJ0hC5wXz5B+jf6avXp0uBVgFqx6xOwcxp+xdPiHlb6mraeGxszu5i71c99m0
icoLMkGqtdXm223BQNjt9InFF7uqUCkZKku8XpASGyDxVLusubI5+0w+n3xSvIhT
pB7AdylSCqh8iFfncOp2T2Cu5/AsvGVNJKf7wbBEjF7vajtPJqV6Uyw4BlY8Up7/
QywThb+h4H9xYhIQ9ItlrZ/sYwv9Y8nCrcwaxSBppFgwFKOFEs4fcnXJDYFaQ+4R
i1be1zIV3ga4k1amOCOR14Ps6NsxdWQsbP3Tksu1JJpdvJ/arsO7QnNRZ6jP5R4z
vccEsVG5KzOckA9WCShqGszniY1OnE1x87tPFGGYdboD4XSrObcsWp6FCksIYJT9
hgqZKy2NEP9IlBMGOeaeZen3ibUPHH7wyXLmoLbAFQd6PjC6+POYSml/FazFdyYW
fJbIwPL/HZj/EnMM8Vpc//ElLL+JfkjdDRzGS/a6EjtppJ7VD4RbivyqQOF6NrUO
mYxBAbM5yOgqTLg9PmCxaGcRFTxwshiB9DSBKsrWn9bR1az2zjXwV7aJDISao8OF
qUsnJ5Yu4b7i45vPojiw+qvXsECf9D+mIHno4hdMPC1xOIQG898Nynvlkb0Eeiu4
ZsatwY1nXApSR/l64Z5qH4KFhDyp68NOSIQFIgeRnn4L1i27w1WbqPt2CWn/9zOx
7QYj0cSbzvYzHwotS/Jw1jSieb4WWyzMFB5RwW6uTRhwXUEmGs6/AG/VWXnmGZrE
C6RZ0V6AmWANJnduxKoR9QI09mtgXpAdY4Qa+aY+N85rWzc/+gmfPv1eQ7VXTsaa
AtLX1opmse5lqxxyen3bgW4tmi/lZA9viSmQ4Eqy4TS8uHGAbXWf5V9bJ1F8pKrf
b7Ofv2+TnuLtppQ7Z/k59vCN3h4BYoJIdyTKBztIcB+Aei6jrDrHzxs4JsFV051M
D1oKKbAok58iz5dpxqG76imZJiuQN8tH/YNdAfoHNwF8ONqT3OuK4lnKUWLpmJfu
gL1SYndHH6AtN6u/Y0bpBw0Oyeu+O5SP1WCgp2MKGiDu9nPN2VNhpQTVH2jOc1mI
jSBTvDroo2QsmCEWBIncUzFCm+9C8KoNOxTlzSjcM+KdW5aKYqhg9pD5+h76r7MT
C2PP5EPkX14fe6kCnPKUPRGuG/5NAKVfXz1HZQmXRicUVggGiAKuOB5AHpKoBdHr
sCM5h89QPW6XqDfwGqlm22MoAn6AlIUqWZPUTVs9LRXM8chDOjDQun7zuEOHhRxe
pQBhT6TkeX1tWuw2PMRBeRSq1nY8Tn3S+S8kkxTjTF/j0l1D4DJM8L9idsC0ZTT0
m7POPwQSi5LzusviBzDhayd7RDEZ4Izpa/0rLB//IK2HbPPfsdxi/r03SsTo2twv
UFTbzUDFsEtHife+0HEDbOlISkmyRkl7cI9FcPKnRQsIOpUppxczLz2dfZ1R1NGt
NyFX6Dsf/Bve7vmskN97m/F18xmPR1sLGmcLKF6wD/zAWIekpW2T4s/uprdUfNWl
7gE6hVgj3D24JQHQk9sXg8oEbdljxuPgFAjzpyUwKb/3B7K8pK4l7n9a70nSI88d
F+ZtNyIIqMMpZHIA8Ucm2GSQEvT1Skz3Y4GuKQVpdICn6HAu+3o1+bxFp4Mye0pj
bTwn0l91cV6emRL6/4u0bGlupFOeKfqZcW3p6zNArbr0VJM/QWYJDaIHlo+B1+Fh
OxcZfuhUUIbIYNkh8ciXYgqHx+RYDtF2ZXSo4ndm8TGU+kw9llvSl3ZbC+J65+vc
u1BkDZDcIfAbaBA5fSgiXAbehc7pqad1dzmMcv2dehrr/OsxvRvOxJlLTNL2oB9T
epjISmpKfRK6tWAYhXPhvP8YJsk8ueZ4Q+uLSz61EIaQS2AXq3bjnKAhlHFF4EWw
FsUpVEg4PM7eNSVjdgwRIWwALiLJ/KpXsUQf78Rb1et2vQlkUm7n6c6zzm7yPMfV
XYe/Q5rWZ+cZvA2mfCzHYZtGQRNJkhWSP6z+qtOUuToGnN1twqmBy7Zc6DIq2wye
ESOo5KWkOq40WSdb2jd59UHmKZ0U1yE3FBI7Vm7uQp4kS1AjG/d6AMyduaKRSkc6
IMHqNIPvxGINcnThDBNbeXUqfMbWtsDJ8gfpZYd1kElKVqmoPD7V3ffzHrhuU/7D
gO3lAzGVUba7ThcY2Wm5mdBOHb7oRcacyyBRi8Uu7a1+9gNIK7ikys2ISuNbFewe
d1T1BlFYR25SSLuzWkyEPeJiQNZKWRffEaaMdNS+ks6VQy8qhIm73NF31xnUgPXi
FQwpR9r0UoUusXGqSFMpmOQEH4DNXlgjF+OPbukxy9VqsGhcTb8KTRGuRA3HI4Wl
Yl8bQ1yxwWHPQqxnmHw5Ly8OQdV/AayoJoxDgawOjEUuwgiL1sd/2i+iQ8NRkvGX
LsL2fg0dDVdVkghdBYpX8GZFmVO6ceh3aFMr+uLTpVY8hjayIZ8vwu8+EMaZyuK8
+QIo67wdoUvO1vdCdKYGbcEhbVe800YTZmIYYR71BFIZ4EsLlsR96tfoIaMzssdz
HVXEv4LSioBBXOrxL2uz84mXvUD0HtwGtWPnRwPawTbiWTpuFZ5agco3xYdz/kdO
UXmPTEZMiUxk5juwK7aPU1x8mNk5SozP9ZjYrBA3mLcBxtb2VrNx22bL4GGGLM2g
6JUTipiMFuDM3Am0rmz1OVqTPrpYMxHCK6NZoIcC3q+f/c/xoASW2NoVCCJHYONm
6MpZ27N0dQcMs5AbwdVzVpEdZGI/q774Z7F64F58NICj9q3T206SErLKfvlQgSxE
gf77MRYhKjEalWHTxi8kwQygJJT/flDPPORcML2N2/HNfgBvwHKmPppmzpOXD89w
qX69lVu5Fb9yyFLRqTQl3WnAbReTk3pIxSd6AS1Tg1+bydfB92bkhXZ33/MbMtlq
EoyDGE4Vtuk2/CeTQZSwOZN+u4UK4U4QiDhjh9ZkbFmj3uCVMJ3Qw+y9L4VKfVVD
mqfKiqTsRiyHvGnywiTNj12pUuvphutDFlUQBAQv8MmyRlw+B8SQwiMSig8KwUKi
nCpO/eDjXY7sJvbBoj3UVXy2nB88hqynS9tXaZtKw13ZYghc89v/dfJXfC2UyRoL
BGIeMFI45RlLNl75JjbipkCqQalL0b7v7nPxINEolISwSiAT7BEn105ALtO1icxS
FZjCr3wS3ZAeMRriAA5Mhf+teXdVcyV5bvgPs/FEXjyQJ6VbQ/oqBAvF0sawjd29
s36IGlxJFwBp4fn8pHCHN4sGIzGTp07BAr3CbGBcSoMYzo41v840G4+wNYL+MGk7
MWSiRsg6ld7qDqWsbs2JEkqlR1PKazuCkP9fMSE2IHh5Q010MGY8yLF50PnzJaBV
SQE3gAhfI1GWyVGVDtUpRMSf33jjQGBlOQ64wZR+avf5Z41vUgfBpdbxJ1Ok0Edy
yi3scUc/2i4hwn/Sl1oshTibos1kWlgyx9MCXaJkkUQkcpqS7mlpI1up5dgjpCBT
58hklhRSbOYY4cuFEzy/t/SpYFHDvP8FjNAkFl6S8/bsu+dkWqb3MGW23Q43dTSq
PUoIduAYHgPc8Lp6Nsaf6CYGEJ3sJ6F4wcdYMDJQVWkXLW9W/T4DqzCwP6sVs0q7
QCZ+vPpvdNTss1KtbeTTZuiHA7MKuL+iMOzgUfcvQNzyKFx7KnLWLkAvejYkkBWh
2FoHWydJbumtxs+vgiB66dDuriCaVg9cNYaop0KWTaGhFFL/w84g3T6exPywlD5m
g1uydaGX9LxPl7qTeogR6QUpU8ux6EN0w9I5pKpbWCI0Rcmc5APgOLTUzRstipGt
RmNPdzGXViygs0ZCs7WRwN6i664U6RgV23gGr2SZzii5W4RXo25zN7kcVxhg1Uho
aHdW3aFAYrIgw5Dg6c5Ndfc94cqC9Tcrns9eBB5B+Tm4Ig6omjLSnsZQ/s5MqSok
MrSv4e7+tw1aEPRiykUly3OFBdjHeRl0Spadirrrr04oLqFAQMzv5f0UGeCMlbVQ
t//KEQdoROhVZWkQIMTrGCG759q8MqNaOWb23RCUI57mD/HEVscg5ikpFiZzmlmz
Cm0wxgEQWy/PUJFWXW89curFgcVJUMLFSkk0lfHR+shVVx3hO1W1Rl+x6UK+yroZ
URp4sEL/GwastTDBmBB36jB9GVHk+Pv2RlZDPFCmfmxV6p5fb03xNdhV9C9G/goY
qSX02dlemMMFgN5yM0AknGYT0SkjhsfhVNyseRR2lcrbSX6P4ulfuDxQGVXkytSp
evPqvKueTUX+d4eHrHLHODikKyYo6v+xIfA122W0Y/ivvnYIpSaFggiewAYW2Erv
ZFHNmme7ncWev9s9NDcboIzfPKTbwgi8ZZXvwheyK4u0UkMBSg6KDRORHY3qENut
Rxt7MHM5XjN+wosCPYNZAlyLejkxWIcpV9xrloUlD95mDSBO+oG0IIbQprdw2WPX
Fa/QyD8A6UsM65WDJUuiOYx+Ss1RdKfMQwFR9bJh972iXmieBaRsIrLf9fhBRAOk
kJZZabYNJsp5cZjvDY9NaZrjZkbWZgqr1uUqLJMjOTpINOsmKdNn9bWGQtpkb6T4
diEzBKIW9YPC2jbO9bYlvtB8y9bDIYhTSn1wbiBRxWa/bQLjeaV9kQ8D894VgSC8
Cnvx1BQ//EOLXrDapA0B287RKIKJM27VeDceP0wPMolS2BDDb+FVFm3tWdqqcT3C
PiHhFo8euTT0PFQTzuf7tKHf+r+WfySkbSMMNaOYxIy7mHaA//EnbalxXCSiINEt
56TztK5XqsVFEUtAvDx04Lj7C23RbyoNbpjP9PhUGZ92g9W43FEjXGutTA85lLtK
K8Mh+sDt96g8fsYU81Ka9LpzEvqeNP7C6SlK28ozQeZq3Jx9cuxL/FrDLtQ5pJdu
xdx+ecPz4Q5mCfT3vy0U1rJio5YLwYAhafDhW5yNT7BWULs356FJLDCcwww5WNGq
fI19BLDXlBqboDqFkow741559z/I0NL3/rD5kQVXA+JS7H8qNubPi9kblLINx9BH
4Kk1eRgr/4o4za2F0ogv29zCCYGEF5OnBZXrD5tOxmPX46fuWy8Z1N/UXpy8+TXb
3Fjb2mLII2XBBzWSG5hGPFcG+k4+ScwlImYfLiJWiktaDvcnQ7ubQ6amtA0gNC5o
mV29PcOVK5K5ZcMv7pJ5DAUNtybthsBhBHajGz/EYOBMH+Kyzi5m+FhQJUr+flrX
ahAlRiGlfYnayZjX1VrlIXwGDDXT77c+6eTbr+1G2C1xKR+4m/bVQKEVYMHtoW8Z
vgUwDyU5vW3rGl6mW+7jOEfO0c/BDjXhwG/6Ra0hesBdxeqBW3lQHSXSN6jtCGHS
Wx85jGFJgTShMNwX0cxfiJAfXB31+jV24B+kAO1ubHcQbKo6ioiWwQ7Uz6xsnZIe
ws1Te7bd4R7P4XH6LP9jlul8sOOKJwGTyb1aa0BCahhrp7GXEczw/3lDZPgmX4Fq
gl5C7Qin+3B+/9HDL8h08uui861MyYV5UTai6jlnfkJ+AoaBdn3GSLzoats8wNQq
IEre/ipICJ9j8UTJh+GqSwL+7R3t352x8L5IyAKTZQuLuf5WHUqTXMW9zmHW3zuj
ZAw7rFcBKe4jUad2MpeJkm4eE8LX55QOH8pWmQP4RQlbleNUQZPOXEVEaICT+N52
i+zxkvUOHOaawUQhPzzVGnewDGVC/XE9p2A1G62epJ7BwfC+9W1SgRSD6cMLWFwd
iFNMQlFlcCQWMZLP5DnDqMkH57FuUzhOU1abjf5u0JZxzbB3chE3v5INnc4ljSGY
DtsOIT7P8rrVS894sEmsaVHJzHuiff/jHee7aaMitKHmTcRPfIg5NuPuUaiE2VCn
XsbazGklPI9sxxjgs9UT4C3M/5VWn4fKkz4gWXnLXWQP19GYXyxck6BVtFWMpLyA
/n1JCc7ODJcaqSTpgMMBIxkKg+dUhk3Ledt4oI7CIYYyLka4DZ4H0JaqvP6WDFzs
IOW/cZ62kep35YrqBp2oqvAg4InoeRqaj/i4CCk1Gc1iDFRXl3tkLfy/S0dL5/Vp
idKI42Fs3Bfz4zzyxJjHSETUwrmSe9t7R0gNj/cTACQ7g/J5waB2Yvu80Ky/wM/R
vWIWFZdRozB0LJJ4KAA+qZMczfVyLJte7Pr22kmYNjP/PoGs4c5cbCpysUHdHoua
+Um4F6KG4T00ATQ6onWGCw1dBWJHnwhzt+D9sdLRHjh+erqce8GZ8eK2C2MvTWCk
gMr33+T8UhWMNoylTG2zUKdY1zQXgloR+crYBeFvKIIIqMRNSOpEmp33Ep7ZATZh
rGEmLpJUwcG6RtoTUOBMI6IVi14634wYcxDKr5dD87SYRMHCERKSR25dFo0GlZ7R
ot4CZEs/hkEj+ht2FWqNuUl/oN3tkWtEepzWS7A3z1uEvH35o6K/kpY7eM2bg4d7
wEt6UGXmHp2HM23cfRHoaCmja2yWz4yT2FJ2RGiwwequkay/xrBu0X0qH6Ba+Jcb
iyf83hXUBD2c5/xlV4eVrLTHPUP02UMwCwhUEgryf4B/PtyvLJO3oUUb0rwXPIYx
JTPJhIKiFWxsaJsHRtfnMJB2zXnCtArdXuKqro9rw4rjWR8eaOLLbAzVRoA3qk1O
fatcWlutI/ESGuTyjVH1yXyUwr6UbYC2LNrF2scRpRe37aeWHyDX3OTP/i8Z3djM
tIl6OK+SDJiHsS2CK1VOwzksRq/QyxqFSBPLa+OoBnASwZYHzGoFvf5+mvFGNE/+
cFWMpWhyrkGbEnjmh67kUyt9iyU46x8Dpt1mqcmig67+uwl8dGB3Ok5TdPzKO6Bj
CMRz6cINUY/DXEYHBFW173pW11DUUxn3b2rz7L6ZLYhingEmHBGQYaCs5jUI09rB
3du15kz675K9esVQgyuGHXKUoCmG8xmYzXg4FH3E6gw4b+qJhZPEG7sKSJS5CeTy
ISv/LcnHjSmfOI30Pj3EiBJg9DCn6dDenEFqbQVKiWO4u0pMP4ubiObbD+xhPM40
29rxPfYdF+b4ztSJDJAzhGFS4oVRRdQoNcyYt+QiHF70uPSTQOkbObXtNNuXneq7
HiJxCvsqaIrjH13jnNKo/PMGLjlpM3e5MyGdvClmgxMAkI1fENFSXbyPZCevlgmR
AOQ79p/rYyOrdzkKu2eJ9fr52kY/lM/PkwOm28RgFGfmtZgVOcgjiBvIttHnfXKn
lhDKJjpL/hm1lwRzY7vrzuOV6B7Ow2cMhpGdNK2zHUo+C//Mc3yTbpphopFU1qTs
7/hzXt6ySrLNSxYRkBZLoMnp8AtaVKm1PM9WowBKyYGai/m24p52r78T0AfFDgp5
Ki/p1Uj3pAzybiS/HFah4dMiF4bYgFwnNJ0olHFFeUoxoRE7SIrs5VIya8Y7b2Du
/CpQqVkXL2aCHWVZPAREeVs9pQneADCB4U3AcQbtZRqhS8lKYSYUFj6Urk+LUUnV
j1+MhU0htcoLoVXXmsOwIUYZ/FgxMSu3Q07UZn6tfMV3eQhq0Edsee05fT9h1HWf
f1W1knRvCsXGraQ7YwRP0GD2Q1Njs/J1dDHoWtdngYHjSaFJxnSNqrkmu0peGIMT
sgzRpAXFq6yxYY2F6Gz/YgGllgzZkxjnOsfmLOLx8dT6iS+XZtKmYtm/BAY8O8FM
VOCcxFOiu9T+dXwCut6aMiKsB4725HjfFCou5MUKIIBJcVBegylYYBj7F5OCMi7W
XxLhFV9dol2RGF7UYsFaCtjcuMzZQW5y28bNTpX0HsoKLf+2knqkW9Otco2IKSZO
isZBa6S7wzK/z5sjPTi2E3mPOEOFVmflbFguMDVZQEzDsGGG+YVLlkkBvdzBIPvE
aJYJDVmUsfyA+7U5EvxkkZQcwmSNcc76AA4rVPFdF5U0kuTOVRiN5s+QGCLHioq4
fGPSHLj1jCI6EO5kuIZZ5xy5lEDjZwspV5dyJbyveUaOhAyvSTILVwj7yuclN1ch
PGEMoYKFGiJGxflNR4edTKKNr2p48OOOQsTnkSfWp+6XzCx3/cVvUyiUzhqdFBR9
A4g8Dqsx5TusnMI6IPGOAeFEIicPfo8eFbvva6W+aQdMIAptFKlxkHmX2Rt+ykLq
jj3EPzBLixSCuk3NcPpDK1/1U3BA/sj+j1a/D0w5dxiGRm5hCrlRs5UZ0A4838YS
OP4zLDyRrvESpLfyHl6WrhejIUlSTLi92KJ7wRiGLPcBxHI4c4BDEkKL97aiAjuM
iy3IcckQp2/8DQTi2Ynn8dn0WsQlt/nAwDrVt+VOmVZmNI7J78I1A/7X4IDH9mHi
DLUv3BIVshnlpw1LQeIVpQoxKgDKBIATza4UE7rYPuBUg7xH54KL7eDma+WfHm9h
y4Ye5K9EaLzeMaXx0tqZCSc1pmfjbunKmDbBN8TriasnI9D/FI10Urjj/lI01UeW
iS/yU55p59UX9Yv11NOkyMmBLabVl0hkPcaw3mZuwqsioah/EX/R3YvWOksHg0R7
PCaAeo81cY18fsd7GrvmON/6W1bS+llCzomYjELwMBO/gHLgEcGrly5ziI76+z5e
r+WXbK2LDaN18O0bw5CM9mXo6ALDpn5Uhgf+FaVvb+1q4sXSEtBaaHnhtuQYpKYd
Y9Bicr6HygDWK7VzHg2R7BMSxUXEwUU5vU3RT1qP/vkc3XVVvrp/95QaJEVP3txi
sDCeu+yte3n30Zp2DyU1qyaBi6v6aRwHz8BjJJfIuKZKnqTDP4HaZobhbg8oHdem
kBPh59Df8pxDWqu8ye4zzpXH2W9cAKrmftu3Elo4iA8g+P5jTpT+jOneuvLmFGS5
QZtdE/DZHq4yEULPVxaj5+rfU8FPCb7x/AI8efeW7SamDrDDVCAK3eRudWkDHQ4b
XhCM3KbEQrZQwWyFGVJC+Edmrm65wFNiZOjVdAhSaawhoN7qWouCtFaeTR6EGXmO
ywhEULU/9Bg3iiFOML/blAkjp2IKu0jQUs6hkTt/vnT7aC2W7RNj0jLeO1M4Xc0C
+KSCrk0j08IGCkUX1O2tFdtfNHN4cVy6PT8wzuEzW5KNKfMvGN4yVA6CZAy9ylkj
UYgQ35trGkL3XIj0RFPUTExxtjPFa0eF5XBBzsbYifBMEAIdU+R6ZQRXgu3ettTA
fWl2RS0CWKZ3gIxi3NI8K0j+LdXcXpqnxbngVWt1AQqqeWlBcK4p6FZTWEX9Q6Hp
QsxTQ7I30B3n7sc45W+JjoZnOhc6egWihciW+GEFU+fG0s1V4FMhi+cWOP5WRYi0
gFwtU5AvVJs9FhpCBWMLMLCaSDq9fNncvkoveK7ZKF8E85rm9qOfJ3Fap7Bs+rHf
t6m4KBlzo5GtaMrO3i8e8WUDujOQdRdUL1xNzBDkmauGlZvugTTqKS+sQdeA/ZCR
sSlbbB5SKinkGG/Q/CRQxLAuoKBFQNYp9C2tntAnJHJFjkfFRTEd2AoW/JuPj3op
dB2f4p5b3dk5Mg5WGzQ0GzZXN3NBMMbBQrfSwaFHY5U7tLetfXvNJCVH8LAXeqRN
e3RAszS4Y5QTVVyI48pMP/un1Ei87G4j6CDaz03auvwDf5u625X6ER6a+fzFBC+a
0llUbrkRhexHMdjYWSfNVGNYVVJxJ8+bjKroLwexW5M0RHOZ2vqejspIhEVxCPcE
/2DAdIumM+cI6Dmgdk3xW+1Sohe1gHWjhve7P4Y9g2m4oel6vZoSPe2SCz1E8Ery
4AM3vyOlWW3s7LyXeLJluQQxfETg1BWFm51GTj+EbOTnBV6bakel/qNx0fn/PCa9
ihDoWLZAe2kEfbAbXlXL4EZ/IW419XtV232fF3S84NkVJ3/4QBFbIG34TJNRHC6d
QF2DFkg6G5ao0aUFHsOZy2qeXpvTJx1LqIwu2slj7nKI07kDbA+FGYEf5loHPJ43
Uak7AAeZjKbrSo5FoWCgSxsfH7KYsYh/gCvcAOw/wBe2shHQCp1wnhQl9GqM/0sC
75jz6PvtL+Hj8T27qGKRmKs/21O4D02rpPnCVLvhFbSSA5g9pS57g5AKjGJLIDtr
DAU9JpHp394eLXY0n4VDMeRhc0kATBXsweeoLyGqo0fdeRIQk9axm3ouCNRsRFM3
EtUO+E0xBDJIgMSgmkHTvwyqJWJRQXED1c4dEd2tEuywDsg3lsQ877PbtQ7oOmvY
uHAtZ8g5qTEsTkrOcxe9CypMIDpTv0tL76diGPDxRizKMRkPEIMdzThQIBrIlYXl
dFHT9tjhOechVTrFQKDUYRowseOYb7V+sLg1gFSMwuxXUajDgkbZvkIXduQ9gK3F
sI2UWtC4/Zy/SGF/ovjNzWxL6Jkerevc8hupaHB5ISeoEm5ZFOGmFgWY/Wz5Rl/6
rCPY9TtirjTMKkj7BxxDabYUqnheHnF+L5k949AcAlKd4Of62AfMdBAwzXGFTl0y
uogTV+0V9SyE7aFtqZmootrg0999RPsJFuCwOhyoseANp7sDIMUoZBARUENe6zB5
a0HfkBZDI39HPsACaui4NJ+Rk9u50UdYlFe1dxn4+fV3nzvSYfSiXV/XdZdy2yUA
nC3WtR/P/b++8eSJvugU0WJQpcdXz+RD/PbBDb3uL1C9++dvK3I6JdCkqmINBd1V
q+gs9ejVE7cLAZIWDWSLbVeDdYsQEIqacMb5WOW5Vmb0pGILzXKidfszVHl5YEhf
9HrZSer+412lTkJFoRok8HZurj02MulYcv5lUlWhyhX/FBI3RInq7AKPqHvPx33A
1Pmmh5uLzc2zw8jrThBIcAXaNP6qInzvpzCgJ0CnGVP2bd3A4C3I5xanKRuoYCrO
v0RHrTT6tf3gEf4zWb0jmHtjI4uSnP6MsJZoexb3hodcY91fMM7h0s7xeszyXV2I
tTiJb7Tn7hh/FrxWEGCXTQS+SL9P8gbuxd4h/SihA818qq0dAI+Cl0bTsdTginYO
AlOi5HR6FLSPIeijY8E5MNKh4yPx0Hl0O747o/0KL/84L+w+hOSmU7kIizASekB+
gkMT/paz5T3OPFLeg21D4IbMxneJzENuAFyXlMyHLSCj8+9+NfVJuCeJ4Y0TRCRX
heKZmtlD26eTcLjDHXErIb943lFn5xQVVXR0mM0klGMHmSlBQgS6KkStEvof17H8
svJIyHVIjtEVdAmbEzdc/Nx2cBUuJti77FzkDJCqCD02d8IQSnNvUHqQU4ulJr6q
ICYkw5KnecrkoFqcRFYIOaX6o52K0gs4krWk/QdfTVVNMoAamzIvsm8UZMC+LFIt
t99ctLQONkhA0jNflKmK///mrJ1njYSZTM/Hu3mLlor2lK2P3E444VmSPPfxe08c
R9lB/BNxEiPK4OPwpMRy9rhMrOxEwGO2UsqVm8JYyO8y/T/s+ZQnAwZIWAZ/2aj4
JB8XO3GmXNGkhiehJbURhBWuCZl6FONyfPii/S1Ci5xkwVZug24qjyKXnTeL028/
paN2sWMqGzqTiXl8iihqvgtHjzrkLeceWqzbYxg1z4WK4LWf+uzaQhLTIP+G9KsE
dSX1n8FQApfL/hcV7n8EjeyLfOHcOLpsD5wskAWxXOiKyCXesGNurtQELohxOp5V
Z1G23DlmMPOsT62s+STLbZU+qs6Dn6fgy5JvBUk+DeQf0905TydT10WurnkEBL2B
L1gRFjOYsMoCIcPugXruTznsaeHswSj0B3JXJmboESRS13GAhd1na9WWQ9atJL5H
Uawpk8c2Ftxbo6UDeRmKXlc3TROfXt/UbQn43H+1Y9ggsRV4HHDN2dMBFDsOldPp
Ik6kEORLKz9hkTwA3ARH34DmVpWS278RhSdsFvbX+zHLyjzxPnekJQCQzNQewMk4
2KwWVxyZY8wGI88lG5HgBWU5a1o02ZqlyCch+mUkRlVDtyfSq6+KAHhG1GeB4Hya
LDwO5kSn/LQQpFSRLvaTpHFG2d3OnypnX/KjwSyQqI5/COS7pxrXcY2Fl8VKz7mX
+lfMydE8nsQjs+KL4//oKuepn4EaNfQPd/5P1/PH0avlizS3tfzV6GltbsAT+dP2
zGKCCihsNROfMBQ1cLHtkaZuy+eDXcvBvidy9kISV0XxftJKcZApeBc2yTw5bOat
EzlHCL7qeaOTpC/q6f7r1zhv/lSLKppZwAZenR9qJ56ESlcaM3HWCykQyO7AZkss
wpvvcqe9DrhIoy8FtxR7F6hvHNapANqDyYoCIxsDpMWFcGrmBoehChEEwjjT7vjO
AlxS1c8WE6auLtYpOwRT9TIaAoM8ujiALqrpNejNzNRQfsp6n6hxJukZRnHmlsFF
leXluBt8HqgWrLLzzcilulcMmHUfO6PT6sLQOl7nBTLUDV8sSSO15p+cRcbsfV7s
4dsoX6ACNTZOfFrclyptUJxHbRxjy8ZNBIT34Rm4Revmt6WeYxQQQsDBOg57IoGT
tWYakzN+NuTbDbCGbMrcu//yoPr3vH0vaU5mh6wpAHQeq+Dwb5siPJ1TGHSx4QWZ
DkN905N1OvM+mnwlzcrig8VW6FlF5cXyZbJQ5z7J4X53svZO/FBhcYhknxZxUOcA
3oo9cUe9656/449W8rwZWa9MwGPCbmMk2iyI17C6m+7xN9ZaDunqlrDR7y/sdzaf
w98geaxNeWbJkJ2WqvwBRH8Xdou3OyZDm/W8dAexVmI9y6gRxMgbZKb2O96Xztci
IQWvbGYUJSNpFcdNHrLDG8x+mnkDylhjsQ3FjT/rBGFpnqjsxEQlrXa7TYFxbERl
Ne/mL501kl5tAqxFCgLC0N6M8fdqHyNOKwtCVpsXxOL779qquwdrLSM2gVFLRYQL
nKte4wG8Cjz9aoHpVmcnI2tlPT0BP1B0EZNHhX5sVmdAn/s13ei2DOHE2E57Oc1V
RhBJRfVSXIFC8zJ5i4HjkqHTNOyLDtmEJrEm+QBiUyqd+oALM0/X78OM7Dke9rem
M4qcaD8eqiUxakZXHQ0ResiG3Ie4cJZ+oqGhAKYN6StB4gMquEuIhghFKEivosrX
zhU7TcRnb5swOAc6vefcBj5qUOTQKmjkc4CMyh7ny+t4Mhi0gwKA9KYHNZZpoG5i
iq/py2WYcw2HgKCNRCbGxFVwqh9p6qs5d+UgUMaRGYCJYBXoVjvo/cKu7uiqDHtR
mSQBQixsNmnDDQFLqf0JNKvfR08OCSQ4KluV+aBAkp5dHoVGLrAxST/nnmtOByXP
DnNvy/zDaLInfsxsuT0tx6vN2yG53KrwN1DUHYG6290YjMjSsWAPCjvdaJcAqjqD
//jHE+fZ8qfoXSXeALxtXDNmAJSlJ+K5OGW/w2M/cJTvFvNU9BMNZVmLA5DXWTDk
ElX88sqYtR+gHggbbjz4MP4TQM6OYaIjT8nG/E1TRQiydAriUBkCijt7GE8q91tQ
RNJ/geG9cMPzHp17NSY4fQSAMKdyjAmD9ESQ1Gs9EoNu8UR2rNUHV/MzfKungL3X
yea4D8RDWynKct+LdFq+Cehp/08RqbDn9fb5io76JBBA56PAozfdtkXpu8xwRYyJ
RFXLXtLf4GDSftRUGlKTSaaj5GKLRhRju3mTHhvKSZIUHYttlYceeMF4UeqpYmn5
0+9aeroLKZFtWg8nTfGGFUMWlMZnNZVh5ygYuLC0bItnGASqLlhIW3DH5bNMckhZ
rSlKR3imCnS5On3y9Ag6z+/eMZJdjEZ0P1kj8fP2xtNwJhDA4pLOgOi+aMknrzR6
m/Ch1srDwDBzvOeNIIz/dlfbbzn5AiX6k6fFt29Af89tw+mZrxnXO2AB0TPWorW5
SZNR0JVqvurEQJ3YryX1XkwYaQ4tAVYP27SYE03uofVCrvUxcKxwL8pilQGcKdwO
1lpaKlSYbbKkJKLRtQN0GY4y97Ks9Enp/IFe3ahDJmQqOWte3pPX2cdKDAn4MQJB
6ioQIZpaFBaMsuyOGAxWl+meIaTmrfXuxLmHlt/rjc3AEUfZROmmMZmAoVRBeUUy
hHdqKooW0dH5fFk+gmzY3UDO/o09vRCtZX000cI/KUcWVd3vojTgyxtRCcOh22F4
j92ClNlCfdYGdTu5KQYGpJpHtTFNnPVSOHEcbPfddhZ/ddUs6UhynNk02X1Fm5xk
ZUY53WntpuQmz5RvBiOOKwMP6sbxoWJzAuAG4DAcPwuANYz7LhkMEBm9j7GHEf/r
1iBH1KUraNGXtl5gP490yJRs7nmyT0+r3gpNILe1V9IWEXUFOXY711RLp4QLGp1m
g720rbirBlzpnyWyizgvnm2usenHuCGLuHNrgPsShX4rjd561YgpC5N4LcIAsu0w
SMlATOSi+Bw8E53GB7uV989oSv9XkhVEdOIdXxcd+m3jew4q9sBUpFtwk6QNj3fM
h5kfhaLgu827+xfbjuUxF+KnYiijwDJY3bFCXKJatsDkUQeQpah93cIuKMxZMqAi
v794mHJLoO7tttwy4RmqQ2AGublvtVbp+ehI9PYyzUY/xjijV1+ObOcT+RhZ8XVv
GEVlHJJmM1zN4GhIIZMu344XlL479Xw9rt/JJxt0T3k5IIuEr1mFTvZpbGvyYb90
GV05F1KkWCxseVsq/HL1bk+nCUezpIVUlnLDYKWUOfFTAeGT4CV+yPGtDzOTp7Eu
eMrm9YB1V115LgRMS6/Sj5DH0+2Xql5uHQOdg1sSvOVNuhLDL0gUAmlWXy6/iTMt
kAo51aIXhhlzu+NhCCYV6RU2e1z+jFrUZ0zwZGd1ar5FdEN6dLgJ8uqEctgoZQQC
phwPVVTkjPLPfzotcKWjksEmKHCyit3q8ZNV4jTzW1ze7La3jNLt3J+zYbQw4NVO
TWPbNFx2tWnLp5oINjhAjHGz3dnVG2Suo3Gpx9dBpl5HgG9NIKyJJUAqNDoq3Q+2
CEGqsm5bZx0huaUM1cYzctYZrHWkohNhCVoqGH/fB6amU0V6T8AdiwGtieZJtWZK
1QfCBWq7KN79lnk2b8rwyp11QD+aHtRTKraIqqbcuOVAgD3qW0taoYCPKs0DOZfU
+Dy6hc0ZmWuOCvpyHOKrVrQZKXnDHtiDlygUO1Nd5Q+O+jiY9d6MgCTSiZkfk/+w
QejNn/vRXSx/9qv24Bmdkeiec6zwpE6WC0a5OvAldL+X7sidljY3Y4CSsrNCjYaJ
HNxMLg8xGze8bJIGnfrE7lVq/ak8q6nr5s4l0CDLdkxn655Vos3DTo8vEDCUccw+
+Zz7gdH44AQc7d3lILFzKO+ieR26QqgK1nC9uZLoJGeeZogvtVp7DtjNua62YBBq
gN+f6zJxUBRL9aAJJtUXqFOgaWsKvE8Gl6s0H+FZgKDmsqfqSSBNGSVZRlE8eK9x
Bx3MbPXm66rz5pGdtINzK75RPI8Ron39fQWGib4Xa6bYU+eAqmVEJl73gMQOBbp2
xLivslyG8HrRhBAC8N4/ptMwq10BaaV6H9s2Oc5cJCorjb31cKbjm/LRBCcMILBn
RqLZZ1BM7lpVHUF5U919hMJ3r/9YWSVQ1LL58V3NDI2ow9U2dRITQ3XOU9Ydk7Pb
A+FhpBKmzG3UkWdeNIpKoUp6fz8cKqtPbemGcdhe9neHf8QFpasyKmdogK7uHkQW
SkJq5bw6U/hb80eiU92hsOsLQlDkjFDGrurL6UKPjN5uFLgb1K7dQqwXSgDkVZV8
aEblIOy7djPIitVYAYwI3GzSUAnw+IlX8fr2JJYg4EeFzXYk2ip8AwfEQuKxhQtA
HphPX0fR7tnDADeNT/UCqFE984ab2uKYcD27XSWUenLQae7cN3kXM/HQq2EsSBbe
+sLzEf4ohfqrA/DHv9t5SnbPDvrPfBRMlnPTPmgQYF6bgQv3koVgRiJmd9h2yR0b
cyh1SPuVG9a3iuLcowJMMyBhkm8g44t8ylJTzzF2yvgGiR8giyv/12ew3Pwk6qLa
SCe0/SD7jlq6EdnX3yLBcrpFqSdaQ8xanTNQV+PhXLFVx1UPyNn1J7NKVojrFfqz
oCuNDZ9WC07MGQuSnA8E7kZl0a1L5c+EIjHf82s/MrDkZSVCAA8TqoXEhMNM25Vg
aathJ5mvFGxl0HeNtV96T46qRtu+cs7kYVr3njpC8Sxy8bJQE7kOGwwOXXTP4q1m
GOh2MT2xNEwExBTXFPAiw18UM+o4if6RS51dY8Jn4veiP7rViAQRd1QbZE5Jovd4
M1rG4T9GLS/kQmNq+o0tylfXb2wRBwPtET4peq8QEOhqaGhU99A4ZNc/d22jURp+
BYML5Y9XZFU3JZhR006K8p2sFbukq6OhjW5oK+i/rA8qocracerwxayOBNbouqi9
Au2JdIG1XU160Rm7HY0B4DPq9xw4dQ1LtnvOj011kdMlVh9gBb78sGlRpyG2aveM
VLxrp9DKgWTfzqWUPlXjB1z8sDt0oUbPsMDJXQWe/YwFZgl1OY8qr0Fr5Tz0yfGE
jGBtw799YzaE8gGG0OOVwkhq62wTbM3EtFsyBxp+fAc/xwmfBQ2kiFNQBO5xyWRm
AlGw8Hs6WKqrMVM5WIdp9Y4yZ+nmKw+AV5ipicXdMP6rx83IOlqwzRaYEdzQiVT/
5CPN8dLKcOZJRxykDrbclfEVHpS2j+Xf/fABZ+7KQEzdyG86OfWQ8i2ZqKIXwM4I
RFSmlt24JD1TBllxWsCshu4hjkLtm0nO7JfNH382N/uNRVOhORxGzctwXDk8zWqx
bdxYiWKHxb6DkalmrR12De5mALcPN6WH8DOOvxVkpciYlS/DpAOqkkHQRAosnnWb
rGQDcMRPabQmMrmC0qEmye/CH5hzPRp9xseq06ubwx+E/02HEGS3AiXCXZj0PFK7
1PMQ7Y//547CdM7mPC3g/FIwmY1stb+UFmPufVUeYOwkGSUdrSTk0+ueYF5bIJLW
J6FIEbV8AQiUTI9SOSdQfUN9TW3nXNtlVgCqGVis+R17y2GckRZWkroO6mpSopCw
Tv7CgAXrUFPWYyh71K+8FpQ82EatsLsvSZzqTrUhrOnS3vDR6xgE8AR9UWygBbV8
BcRHxAIFnR+NTX8L7sQr1Z0HEifh5KaXsAmETQZ7jDsb8sHwhH3amjowQfzRZdoH
TS4J1bL8SYdtKv5em7p5uH4oSs51nSSjCB9SeFEB4nTNsl57qLVedA5VhWxHNwHO
rfYoqconcmB/zLayHOgTSejxSeYEN4fJ4vMx4G/Bb7K7LFFfnvtj5MpWsOKjHSSz
rlMXT43eCa2gK3IpePDmEmZxaWOTID3zw45g6kcRN9uJSDbcf+dplHuE7DAAziYU
uP3g/MfUVHkShLkRD03h+NwxwBCsFWvUZ+6LAbsFV5/dVSIEBw+/r3l7EkKR1uHx
Ik74ZiQ7F+4SG4yX//tlTzMxjcfw8zobOw3bpvqRzkvEa464h/7S9TQhNMYo4jLE
QaTCXXyGeDT+w79OKqbQ+mT9somQFBObUqG3b2P5buo3AAtIR1C/As37KtVOjt4O
BgkLbH9vZ02sK5KhgGpbnv6ZUbUyiM7hwBQtIWD66QFt6nQ0M7RfW8qKsChNCu2S
I/nNfJjnLDsSy33y7fShkYIbKAz176jHtFA8fkkYX+rXl+zwXDlXK3Wt//mxla4b
vH1xK/1bdfZegHz4DrrJqvPDTB2oaYAds/vjY5YGnWjyTytu0UuQTXDNAX5wdB/P
3zI+5IY5IDQG1wJegwIBT8cyVDsAnIHR0SVD2Qpg0taL8mIoej2h//+r1SV/cgGR
kFjP1Mc3fNbVqzqGeNNPxJzmDaPb7PSXhiI1eD5KOKC7HmDkGSsB21tkazGF/6G3
bwmTSl3AuSNm2KWOWRRMRr1q//Z72LMvz4gs6L0ngZzo+X4aPHYeuqUyOwvquFiQ
nM6PZaZZg1CA39RyhPhFB3o7S4I1Ey3oLY2b8ACYPXawtHQ6CIXCCYEiOhHdU2Hx
d+uEE68+GTCUWN4Vz6m30EC9qSnPpNolS7ft+7REdMPU8o+qgk5UjBo0vitHujFK
vN60qYQTUKs1b+B0k0qK9UhBga+t3W7GNq0lwc2YimmEk+FW4lE+7nXfaXSCvatg
42ttxyN1i4LgVolkcCDsT70oc7CWTMKgw5yMUbRdCzBkqtBUA+OoTFC+aeZcSOvh
/jr1111C1JrEk5z6dqf0P6rnyR/10PUppqcRANpohG2M141/5XU+unGHJwNb6mCy
ROZvMfm7oeo5YVU1sxwjx8GyVZhMr/Zrv7Zs3yOQjQGuj3vPXkfoYlqxOe/V48pA
H26slbwCbs9ABNeuknLDfeVjc//PIK0RNc/BJu65d3WpTBTlY7tzGRF1B+BhAkRh
soIYinf8YAbQ3gdiEGtSn0tsm8Z/m7iu/dKUcj4dUYpDJg18chm5LyTH7zwhBZnc
J9w36oktpuETZJYNekQURQttOUTwTiMk/hC8QRDVXocikKrZPRCvgTme3Dtc9RDK
OevF6kyXzAUbS3y5eIn4irTD5BA9PNtmNTCN3YDFZacPSynm4D2NtiMwxN8Jg/mC
LCr5NIsJv8tpbo4eZd9p7UjmxdafQSi3xE1WrpRHAzxMNc//Vsivq8Nz6IXx+mnB
l1mVYgZ6hB9VfanSgr53dy/H7rohC/RvM3L3UX/MQ0n8X8aH0NvKJJXgDu7W23e9
rDjQ0Mx17JvLYmBJpcSIhJFyk6ptrMl6QbdP6hh4ReM2xMK2/9/Biq5ut6yvPVV9
FISTHxrzeBwVcTsVg+AooH7e2R5L3iZsXYXAoatsi9AMMRiUUfEsNilcW3qiZ4IX
vSuSCc068vlC4xD9XvX0B/lzbyd0hcvZxoRVbgWPRdXIxaRX0v717L/5wlRr/Jvf
EOMmwwGwnToss+Fo+Z3MBiJdmdEGpr7mismYy4Y2Jhqd4n8m31LGog/rL8wuF6gq
8Nk3k+OCVQnx676Hyh9y0xqOqY73cTkllFbpYSn+PZ9/FIC0Us3zlUtnwHPJlML5
lLTixRr2D70dlIFEorT0IO0qOHU3jX8wJBYN8pcowO0CY2eAXCwDQKoB3XPsE3TS
WmjqK8os8MPAiafcgbAaBidqMe5eDRY6CMQnthNbYtj0DfkwM+mkf04cXEGYndtO
2JB6n/6HRUBYC+Cy8Jcw1FotSXKdV/uzEUHnnjKhqxscFQiJyr3K2UkfCJZh9muY
Fk31TZs09u80o2tzAT2Dr4gxZEUwLP0G7JDH9v6KZDUndm/Ii5UjZJtWvp2aKA3P
vnbkCtiHKhUaP1fTMcp44lhe5ueyTzSmGMFzIUe1v7e36AAyfjnkxxYdqRpyjzyx
LcpG+JGy3dEEgjewjMJ48KHSXyGntlOPnCtHben3HtTv0bSqeeRJVwmnTs7NWlgm
eaQ06FzW9lDCb1ZgAa3rlZWrcoFRFUI3O5BXVydKKfb6DH667XMT3MuR5NmZqgMq
2xzAKuWpo2QG8xxYd25crZPU1eG0Y+z/OqYxmkbS0K+iMBfGAutmAw8+UW1rp7Fc
Cm729M/QSiDugNdzDnnH1b3aGt/gA/ABjTHpGNBVHAuIs3Y/4ZFY/BXlVwu4q0//
B5Vd1mndABLxmPZNRd9j0Y0fNkoTUKzfQzAGUhLKNi/ypxBrnB5wp3Pcu/KeWsGM
t942ARuk00kx5WBTtATQZ3oN2TABNUcY9nQviO7/AXNYzxPTL6lLMM3+KM2KNM4h
dvscwzilGDUBmkWjUtBN5nccPpvmYl2Z93vHhsuatRAzykKuC6NjZOpkO+G02zVI
loqI2eBxPgrA0gH8w45wgcJNs74fkjYiqdahmCFMecA2gH7DXcbG4Y+TJUiqZW0M
zTioRImwksApcDjPIs5sI/YVa+LFgE24HWszW7YCPhYe5qx4H3h4+igs8jmiEqUV
BQJ6tePC2K1uHcda5bsqNq5HvIRCylWDh/Zyiz20DmAUZeHqjU+v3Jq/L2jzrH0I
PBVuSCEziwgloDTl4BWgAJJeJDs0qD1VYOs5BTLOucD/Ic5jJW8TECW2CX3n6Yvb
5sKFdXiCNX9ozPxkhCpeT+NjmO0SCx7fK9UwKWCg1mW8OdbViy96uFHta+2LNKbF
rSwQTd206b+oRN3RzaWuvAsag3O/vjRMX+qWUcNaqx/MSbOwVUpXpuRb8nuGh8aK
BwmgmmSWCKlPywMuY1Iuk09ykglTmIQgtuK6SiPjA4abrlTWd04ldoN0YhEueLoP
WvUsy+p/dkHlOWT5maDw9EwbcRCgZnhL2/cirrFMzvkV6A7BRw9PWom/mVMSkxyn
Q8SCwqkpXB8iWPYsPM8HzYnMnPKdiEvABEFo7Jp06jQ6E5Li0PykAtRj8dawTLzM
Zn+hjZZA/W1YVYPvWUhhS2mvw9W0pApVgMyxDhFxj0X/dTW1r7Zd8Eh0gpFR4ojT
hCUTkEYyMlFlmpvD5kIw3C9nVXnOliiYuHTOdW2avrcNCWkUmOmlWM5yCNOpvhC0
rYuDcXa/FZofrIygqjIeCGVElS3guiaWpz/mnhpUPh9gd8Urn2YivUkgx03/A+cA
c/4aC5DotXYll3fP59edQ0uZc0/ItGiWG913Q1kO9U6V4LDC/R4C/kEwGRTmLMwV
6kvevaO6TShtr0P47dCojc0WcgXU5EwQEdaw7jI9HEKdwEoCX6P0gOGvjpfiJ77m
OSeq0C33B6UdaBlx+95+KlKfcMDbGp8XbzH48ynCVfbproR0go0XeTgV1kVgb2CT
jbJmt0NZ+ayLUMdnHsCOl/ilpbAKC2mIkVa5UQACmmbeViijelKKCTP700L0ZrXw
wPyWFYqufKfXG5jUaBm6ptr5aq3UZfU6OI7xruU9ty5B4vPJLWp1v3VUUx7ZGvxY
rOAau8EigEf81LKm0d77KIyve621wQmGWEAC0Hr/ClUNmWK2C1KJyh1sxqw8lQeP
oUwTK9Oh6RTpQhwNw7DxW5L5wquusaTMGjcB0ClmMVdNqAjtI4d8z7ZNN9vlGoWf
HVhFARNqD2VWHCh8hASKg1liOaYZrygRzzvogVeq4JpzQoaD20QyNHuEN4FI8sUD
44loobKV2E+AaoUP7OXcQcpJi9pQzDM3T6epCPqGYgSgihklhBEOJl+RVd+QFzIB
+8urVHJO/+DsRsLKy+1ocC0RidYUPWDeFmc4Tx4PF7uccPhZhp3nNdy9p40Ezzcn
yNruy+Guv+iG4plVuFC/wtPh7nw/JKqpjzVQbyKyX2AspQc9UajfX4p3LiSu4yRp
iaAqEa3TjcHBZ5fRZvlagBA9+ksci+Ngt0eN9BJrwykNz3KUZOWCsoJrlC2etH6t
wYmQor2T0vXcYArSkIaXF1n9mU+ZNHxVmHSdPJE6MBtc2gNHRXh7/KLHZJ9q91DE
LFLrMrioLjxRCKNcltbxPQxO2G6F/3ONSvg6RNI4bG3zGARQPZ9qTu5tHFjPcqPD
MQrSj2d2zPARIcsKtUqewmRTzQLb7uJ4zZ8sWh6ceCwLBdQ5Tii+McGRHRXCvPSI
K05Kz+NmEH62SbBUALbYIhOXtU1qIcQCwnCS7PHFP2I0yOglAkYppUwjl4e7VW+M
/E95pTHKtshG27Xw8gjypdeS0RKWy9e11JupcXIlcj6mTXc4VHF0YWuRye2aVlzz
sAaNNeAk08jpj0wuu7cto6QJgudxYcVCUgh+dD52L5vFP4txV+fTyuZV1yP8sFJ0
TcEcPo1YDDCY48Gi/AkIXuuZZaEmIq37ig8nL5jtkgo6GucFm4UM1nRgUodOn9nU
QUsCJldT5bDyoeGY9k3uXex0jDpl9zO6Ix6gHk0tRjRTmxAscQjCn6n2Rnst/In/
OfVSMYbRMfiKgDUTf/Eiweg12wxBKDjI8oRqn+NUMxPn7M0YHEXPbZQB4vvEH31U
09Kwl9SRFW3KuXwt93RMwiUmV9UeSr5/ihCN8hjotHPyaL2e9Bq/K07JtVZh2BXd
8XVYjsu57rIF+UTpO//195tvhD2tsuS02/T6rCpnAJ7FVWCrt/+5TN4ZXApMbIrU
oeFtr/jkL8mCjGhzVaiggrRmv7aVSIyF7oYAx1zFoNNJf4CwZsq9R+3G3eF7FGf8
PBrUuSR7QObYcjGhgQqCNiCEkuYZsomBlNH5ZSpyea/m9BJpnn4cSORmU0J7x13Y
8PACqZ/bdHclQT69/41LdWHCjhVZnDv6NcVPvU2q8vxKAdEIAUyXLpG6NzjU2VG5
nuOELLzXcIoLaNbDFnkEos4OBb+LsC/6Fsh4cACdbdQNZtmwgnD4viFp8mnrUT/K
QKAf0Dph5wadm4a/t081CK9YK9KotwAuvGCDVNwAwNKWLgew4+kwCsxQltEayAYo
gU8FR3LT+h+388OxzRVTxULJNHaG3kIoY5j1w5RWZZ031hNi6GUiXXBVyZFNFfUc
qVan/uWKICGKFU4lGhjN4xhEuJ02Cuh1SZh9MaBBP+cC87kPJZvF1z8me0EiHMce
mzUJbowl83WiNaa4+/odEtivM94EKGm41LCC3TISYfvTljNb0ttRWtXpMznsWeSF
QpEF9HDPSNFlDuFQEawBqyJKuIBHRyQdmmGFAIsz/lz8WB+ESYaRQOli1N8A4kTc
8NFHKRUBGa2OdSMoMRIvHAvJBhbMevGcx+JOHzABBPy+ntM5lnXh51Mb2TUIr+gG
jideCvFJqge4zT6xwUmcz1eOFdwHCU0/D9OlCB0E41oPKOn41J6X9vxCPXrh/+GE
QgQyGW4nnRO4YFxSSlLxAZPZdOuYWQktBuXNc5mCLQG12rRp0sdGhz2+k34Cm+HL
iAnFdZb/3nQ85I469kMtJZFl7k0yPysXYBMdAAv9IniQRVkBMJ6f8OKpbjRGIkP5
H/3GpZ8+EpBIQSPAeIjz58d2XYAjYSHVwbfc2OdGo082udN9NBocXECBSM/UiXO9
8IKWbPOYbPoOeAl80aCejvck2fFdOi/ZWVs0KxQmNLvA8SD5KhB4pk9uhIXiaYeJ
dIbjBBeRwei2tc4zY3FgfmgAJfTZmB5Kjp2h3N7yoEMZwv2r/UShDIjMtTvyyKu3
cn6ovU/b/J29r1h7zfh0aEUW1sirdaT29PfbaZRZ8g850YBA4pZezuewHGoEEIQ/
PpPgU3jjYVslUk86sOgNKhjZiRFXFFx8HIr+7VuvYd6AC2v1HstkH+TKbOtvRqED
szObtuWrIWHDwlbO+e/gBf05UoKk9ICTqn4jyR+K/NKNiDCKxF966jSHvpEsthDx
6aXyH2b6EQuCCWguehFuFiJzCIl+Xv9GU3ysMEzVNJkgryDprxGfEbqGfYO634T2
Luc5S/NVMZJY3xFDHAuutVb/hwot3+3T6kn8wNdXWlK6pmMTdsOlbJ0FzFTi8U+I
mLAyCR9ftfaIJPtFDgkli31sez+NCahSxLmnhLvGBUnG19bKsARg9lRDq8Qd0imU
ZrAL6TNm0JIa61aDQ+/l5gv6XTXCd0bzxDwE5SOxo+LoULfI0ogYkwoc4lSDoCjK
n9vD+87RNv4lEFBQ4EiMBCCwbR6Gt87m04+REqevuoTLMhVi3Ya8I2s8WcbxHhGa
a1b1J1fzzr7gPVGWLGufivqqK70fRqBB9KUh/MywpoCzl/WDL2tV4GENnm/FOoC9
AyGm5vyo508JAwcL0gZYh/pVIdesjf/7SR8jnM39h/2Bs3j/tI2DKey/5a2BNBGq
rh6b1MLSBARD6PEmtZ2YCyBCoHhusHApklZLPG8oyc36lyrrJfs/dOwVOkxnVVHK
Ar5kRNh71uXkza5ZitTNx+5M49E9qidRyY0YsqlcBrO4wIrebnH7/p8AzcwAJ0iR
pJA1D/BhlCABMucFBIDVzmHh0nMvJSXa4wdUH1JgDtSk/MfZIDxavTaLZWiFfUVF
eLtXxxF6SmhwT7DrJKiNVi/zrNoGrrysUTjZLLVIaSEW4Cizp8vRwLqrmp2g5tP5
88ZenzdPU7tx7UmmSQldJduIaWJPhjyUJ28wV1qyxfRiMIdPYEPIFCmnnVV3uX7v
FWakIvEdo+3Lktrf0jUyKKFl7+7g1NTc3hY+TF/ubvV07341ZuvCv7bgKgRFVsSD
Pn6oHjwymIGl6nRh9x4HySTIAGCrHb1KrOYqGubnW0TEHPfzBJuk38AjKIeYpBwZ
NM9hQmyCgYnxc6Ox+d1TbSBVklYyG1rhsuOY+Q6dNQce9U/VSCaUHOQR+7yszsyV
ZQRg6C+t3pA4fBmUg4Jl2ZkN7a9E7QhD/BabeyvHCSdq9x1MZZUpBFOTar3KWv3j
X5qZFO6Oaq1XoJ34vIwV10Xw4IizlyaS6MXndh08vQd6KomyTWZ6MTRF/teDQOQE
4CJ6+0RIlTrdquFRKSrw+gARTG0QYe21B+Z4rH7k5AB6ryAXAG8XzFEQyIE/gUTj
/NYKzPTb7atl0Rqr3imYfgEPEOEqwdNEKnmXL/kzMSn0ePVjGSw0tSvA+QGv2cWw
b0wxcnu4ymSGKfEwQ1UH7plLxOH+g94NSjt+6A0y8lGwk4BHnLuDPwKBY831ZqwM
nRjSgWaAQ6C+6C733kNKHuQfWyjV2l2LpjgA4kdv8Pu5hpKvdiPafF0uKqweq7Pd
FC4dSLwdQxO47marTJZ+aZZ9yRY/wogaGfC8JdCdMhzlwKIwZPpkh7aXoNq2Ktkb
6QRztH0RJKgmnEC4aVPqGuSj5ZuF5y0pRk7gAvkwjuBOjgPHPkRSmnxw/CKqwnzI
QcaP5bnnWg5jrP0UJ2t9s9UUxTHEzT7KMlXOwdCWSd3oBs5PoqIYAiVncTgP0exE
OfKzbj2QtORHGBBiHSx8N6N06necD4OXQpeXql2dC01s9LZe3I8r5Ff9Ly8E0MMz
I1Iygy24uot4el2Rd9LGrEz6SQoL70bwg9Ttf33VIzHZ70QLrxfveJLbU521G4vy
qGvCNJQ4gJjJmt7FlS39jTc3Z0FIii7rKrELW2AQD76QPMB7+DuHKuWdUC+quM8/
03eP4QcHGj5oHMbDCLUA9QqEDhemSJ6fpsKT8fFn8jCoNUfiIrKnbEfvwT/9fGuY
zlXMRfrVBiC4nBRcRm+6Bm0EQTW9UtFoxLjDe9PEHJPeKSQkBw4xxXhhw4bhRS+x
cmHvC9g1VeRFGybNhy7mXV5MjojmhBld9jW86iA3nmE01Y/Qwiee16/MENnOn9d3
6CQL0WkLP01uXRdeI4awwHj8EMflFGQmb4hBVcD637XdRwHyk+7cusl+/ozomair
hWbLTqkxHPM1CrDodX47gHA0DrztckJ5IWqD1QPczHVNdRALqcAHvz8RT11bw2ec
bjFD+OOdFmCZ4BWz8VVla+8Z8cl3GOvHpqZbUEb/OpwG1KNDaWLh2R36gBr7YA90
2NuYftM/Ob/8AVJvDAXsoPEk44JOMTFc0hA0G3/btLm/pAp/DuNQMsL1z37/Iho/
03o6DJoe9undU8k9OYnpGKfV5KXVVogSsyNipudSeucw+h0+rbydQhNfTPy8dcvm
9Sz2Ff7REs52vMZdGzFTEkzJ2Dkk6L/+yPzYIh+2wpGT3QDHlcSr5THmcHYXGJQc
XYjf75W93BLrzo57QCCg3nrjtGuUY630VL9iwmWpbTR6ok4OPXKJMWPOx08ENkpO
jl8/NMJqof1XCOeZYW/jDeW0q66v5TyVlXzOgh1bal689kJ2RXkiU09Fptz4M/r8
cNkMyuJDcGLhp1Fhwwbx/HhwGk0zVZoqT9CUy+Ohqy/Pad8+Bx9KimTUUjg4+Bxk
jG0cAHP7U3HcGCcx92nJeZDsVCXmFa0QrTlRPqWuPMjIUJYUk0D7so/3IVSKaeQA
+kiA+dDviSOcCmBV4FsYytTsUe/4dYvM5KZOb7WW8ORDrHjDMhgEmDekw0d3hU2L
NoB7417hHCx2+hDEa7toL6Vm3Dg/jEZlZJI1Sz3qQ12R/SG2sEXr2jAG4Nbe9knc
VQiZHLxQaRRAZWxadWCjV2uAZU2YvX7kDUGSQuzZNzwm8DcF87J/b+qBMTcP0J1H
/47WKOzq5RfA0qsgXgQIwonPmqsI1XFQuBenXcQk+O0n/P2eKoyMLrLZCoiQDlR0
ZJDjujGuWKFCbyfO96wHcpAA6eOVzqIEq7jDUyMfnFx7tRfiK+v45XRuAQZzY8zO
adRAhzt+jqKyjjgUf4A6GzTKzmDb8Sg5XlSpYuc2cT9nBapwncm0MOqUz6/BUrfy
mOZYq3btToLQYhzEEHclzYjMsia3xbFh9iT4v5flf9sJWqSKvcE4zvq5MRs+5DtC
KqZjpY/JoVZe+sMkcTF69AG5URVm5VS7a6HDJid68i98Cv2DHj+engWVVmdvROyh
i0JhbPQrunH4Thsuf0bOZVdsxW+gtG9UACBMwrlVy6+ChPfW2YFChcjbrwQgQUYg
xFkOYTJoH5ar5WwG6B1fW3Nxv7W8SL94JMxzn0IKvA/SThGEXO9nx/kKmJolbITX
852FJX1NpH0mY605t79rSA/y+OX709c7qN3tOpqxLkVpFI8oDCiPy2RMalIwDjeE
Uz9QWaz0F2UXPMKhBOIHOKOrB0HzJ5b8LpD8HJYZ03hAyzmpJAF2l2wk070mArx1
3ZvfQs87nv52GoBZEvPKOIuKWzYWTXP2hV9rZMmlgaaRbAqKbMkMNRpXNDYkEYMs
JvBNLB7v3NBR0WaFAshZTYIHnU1H1eBjjjUTd44jkajuAyCBOpU6WNiXQ8LeGMMr
Jxg+MAnTPVeWr/A3ap0SwgLHB66Q8c8LPIk1WiG9VAmaP4XqU+iLnzlMfDJN4EN8
hMSCoHR4oQRbTh09dCBdeV098xNdvXnrwq1kIK5ObSo96q+FhK4jk8eABDMUg1ZX
OhLfct2rLgOCT5oKl6KcxQJrKrAAOS/Imya2MSI671YxdSd4bTm+MbORpCNcQeIS
51rscJGdBJyo5HSnU8KiXsYGSjwLbhKHLR1jjwokfSFzfYNRZ+tT1DgDdKdfujMv
2cGW64iMAcUfZVNDKc3WxWCY99G8gAoNn5grmrdUBrgSVZyDnxtV+HmwGjSiYTiG
b/4j4UXuj2cd8pujhtoUY5a3GjlxYeFy9v8NjBhwUVkn4x2iffjIYJs3GAqO4Vok
/3s4R8N+8677R3T+Ko0k8mzGKg1jgj8yzB7M/PTcpaHx6zz9tszv7wdRBkBZpxF3
bCGS+wTPLXjW2Eg13lgRxkCvFolFAskJVU852AJvLBRfryzAbaUbOwvAyErXztjp
wLb26odKmry99IMd8GZIIl320ENLNgQI/9k2NqZVsX5AugGhaJ6lrepVYuL/gasb
giuEzKzB9rZl0Th9OLO7uFRBHIkfAbjc9zT15q1pPcE3Rz6KzgrM4cGybUg4fn63
Xo+qvRQxX/CTXmjcHQtOtjX9IUzly7GjGorQivmsyTZtsHyg1Lj48wMjruximVci
CgT6qF3dBuVOjlpq3C3p7yS9KgloXK0FjzN/I+arwaS6RIU4WZ86IIAtI9yFQBxi
b3XZDLO0bWb9vso/nfnAgK6JJWfKtFkMaZfHLXqPlHm+cfJK2/R+5G8lp1qtn/qo
iuRGkzShSTGag16juCw8SmoIe+IFNo0+KEhOxUunUp4+qVQ0J5r9kKtKVHBn8u2X
ptoEqohb99SlIykUnLCHvh8yc7Fbjc7mQwgVoXsHUXRp/FvzIjyEftbHx0FKeTFQ
5tmCwHL6tImgQsyMj0Oc4AZwkKevLqxTr/PJ8x3QOBUCoB3RetjVUQvR+9eue3Fo
p718nZICOsKF1wDJirPVESZfMokoCfpTUC351wF4RcAvqlBOOKqYc/GgOh/8he30
+RLgpVX+owOYvwWRKgIKpa6lQJpVAT2mjQWjEht5NIIT5dIBw2xnRHE3I8T346Yj
stXl4CVu6NmdrrSJDe+Fib5qG+GYG6sHDe6j8wjiTm5Egf/tUO0sz+hSrTYrVuoV
uvJQ3PG2jfKarnd9footQui34PpXfyxjeGzKo/yydpKurD0AD4feg0gmaIm1SVIG
fM7uAHiLX5grGmYoNbptDJCLp7PR00c8Wghwx5dNWC3TbIR6Lt8uNGGjCzCOEpwE
7AnmEWXfLsdgyLQiUG8K1f9jQsGaoiIiyOZWYUGgONcXaIKvWWR0xku7612O+WI6
5WT8TbqzRwE3xR/TKJ2VSYWsxGGH0zyPoqsX3xW/c/0XvNKGAfpqa0N61JMis0Si
pJQdJxeP9X/92itzUvh7EYjnYVEHepXlUjL4Rgso2eQxdwqebQmpxP9Y3+AduC9h
k77SYr4x6WhGQQzuiXCXD3pB8qimeTsx5NORvBxn5dabpPFBp3daBHQR2kp1yunn
DmfzHFKvZ0oooVyZAzTlKdCguj03DN9nTh+WLEn7QROE1cz24h+3nCVeJfi2+2zg
axMthSM+1XcTXliX+XDo5m8BbDt3ea8OBgBDncPBKPS8xApYNWGtvMzffuvybpNF
KvCag/mDH83cJJKVjtSaMj+fwZKe1R8R90xgjYUTCjIqwuTOs7W3D2ofqEh/psg2
MWXiJ5QZW4G9sipJEgkTdy2RVAwi8x8+f9PVyZbxDw1D6limlP+jCQU8U8iYIhl2
WcO9t2mQhsXMmJNOeZH8xcBHognfsc+l8zYSB2bJtCkh5MQ7/4ozsTNN03kfYbzg
OBQrCnLLV+lx4qj28a8wudhr7/2/SvFSk4xvKaugEJdltTjOrZjBZ3pra4YlY8WT
4DWah5i8ULKthKPqyuKTD1daA0YzagEwsBDnF+YG4u5L6AAQRMkn8KR423GQwItR
UqH0OQg8SIKBlDa8jKw58LguqAqc0ZSzii4D9bOarwkChCiJy//gfjU2AJoFKse/
O2eaays7puLVzndWUc41Qf5aM5wL+vjiRMC6IYMJqitIIwDbB2Lvb/E5/GWN7x+g
bQj7QUDDsKYjigLjGESHp9nfU3Pz6uDs8XWVPFXoivnygpEgUh5YjNcY7aQ6+7L5
pdUY6bKszKwDd4vlkNju4jEOu5icwgMcsAVqwURuzmgTs3UGJyq4rLPKPPdwMfaF
+umgP32Tx47CmkS7Zix65OxpIv8raxx2/51dcrNpJN/tlfDlrBpZAvYtSVAHW0rv
1oYdZtdLYdT6tO0OgiM2jvkVU2ZqfptoyxSvQIPpELd6RJ9hfUwgvs1LU79lWWzM
HX4ldm7bbecCDBVTNFGtwYyKAVr7ds6jZTwyAgsJ6VGkMv3V+IlEWJ9lCREzZEhI
z4/9vL1Yaqb81OnPUR/mhVj1odX/ZO0jGJ5EqkN/H1ZwEciSiiR5W/OaEZPO/Qay
f1naEzaBVqvyQrTopUd31Nw+zRyGbc4xY6RLAnKgdSBRUnq6XwOgk8YfaoRxdA5b
irO9/wZjeZOF//c7OIbYsqy5Sk8SFt/3KkaJorpf0sjD+4gmG1ofQnkv2FkqXTs0
fjAxTkVK1ppDTy6VZiLaT3pibqy9Hvi0iZAoGraMhNWLkjOD0aUaF3cqKMMKO/BV
ivBMjJchtj6c92O3SBt6k6NRCF6qTha97JefJiWn7YOT2uZODS5wVJGm5Dtms/Vi
4c9zwAKcG/5rMo/WElv3R6T3en9VqNbwQ+d89bE5/9wfaEgLpeGPMnkmBqESY9+6
Evp+7J3/cGH+EQ+Pd2vxZYgRU5iFlP+tS9JsgPrh3vilyDjKSgSKkJFn44q3VG03
E6RwQT1xs8MBin9JLgTdJTTFi3h+rHXVQIWZDl3A0NYqoXbSM2wU4JpwIaTl7J3y
o+Aghw9U0adgv1KoZw8amHEdUQpaPJHebOGp5AZXAFZt5B2zDjiXlsy47arQMVMx
OiN7ML8nBbhR0VAF0e/IeDeRoI19m2nyFwBibUIdm2bi2ddXtkQiwVw/lyNB7EYg
FTHDo5Z4MoNl2SPdNoF2C9ERO4vs5XoVusrO6Eba/86PZ3ho4PRDpzXTYZ7GdWh6
XVh2TNFAht2/RJ7tdX0Tvx1jNnLHFPiDzd6e3OjmBaLmmYsPr1cp6/XdibF+IWga
7zhpNfQWCMlxfLTXZnEtxdel0Teqw3z0Np8PvvukXiVA6R8XdMgiMnpG0vhVdS0x
Bb/ffurGN8GqmRMAS+zJFRMjKWtce785kAzv9IC2rHhVGPJB+ow7zbkZAWTEwe9M
Qz5995PcfNAAPRtepDNOIlxBqoRnmpQw59ZraCFopBPMF7nefkXp8HTGSg3N/Y0a
vY3w0nGPAUZqPV3jnA9xlzOz3OVntX+4aJxFOFTW1VRhPOSpK7FjvKzdVf8hqH2e
oeG1D1eVaEFo9X5COhh2jDA8AkFUIjkfpRQ+GgCyY5kHkurtjnutnl+AoBNZBBZh
e37NAok7Q3famYLwUdWCe1pSAhCp7K78IztlYJ4OUDgrwksd/4CP1G9W3V5y2Jd5
iQtQ1AwqKuO6Ghbp0koVlL+OsSajOFiGPPBscVr3t7UvsFh+Ix5RUdOWzJLVHBtw
opHRIOxZHVDh7nJ5h/VKfN6i671exIButL5Zcqoar3d2u4w9FsCqDQLvHR05AqIr
28bHCZlhuMfWqrV+M3Ig/O1DrdflJ8aK+XsXNmP8MsrCFvWPks6A6TBHxVDsL5Xd
vKarzn17NOGMtB2o5jLN8BamWiIldKri9YGEZgJjSuvAEdqeYjayx8SXZ6UfaOGj
y2clqC2jfydjKXTfA9pGHE0LSoXWPfm0h0H1Ld5iefnAwNQpz4mt4wnWsgzYCJ55
OXfA2se7DukP9HvBoiEU/BHc7F8DyHIapuKSBXnhqmtAxV4RN9mXdxoihedqX726
Mag0wAXprNZsPusG/DV1Q61h0F184dhVUB7dmQb1EUIzE4B2fPSDmtEg8A8jjD+G
LyoSYiU11gPP31Tb0KUhlrYs5PrUAYFH6KYmPFNCIy5FXr+zqlefzkLlubY6uqbl
rKC08ETC2/jsDvDGMzdNOpuizB3kuONQRSXkSE/iNdL4ucNuztUBmjchKYFp9zlo
XZMuP/pYPo8TsFRssqNXyPnOxpcDjjpeWdG4tPpeZhyoWSJj6SkH9+GElEFjd3Y8
a0Q6EaUG+EwnoA/jPclrH0qtm0OQm1vi9sd0ockgNTyJgg4kt8sfO1OnY5Lysg4v
m9+gLhjiSNkKlYn5vud3VpiPtRMmIBkDjlM/gIPNXitP0myVxd4UY1OUxnsaFk9B
NX97C7qukrWE3mH3OZYMOQXd6gYLKZ4r9qdcXkYcW8IltdW3fukD/CSkdxA07sjL
IqpoaFcTLx3QbS3IwDtfw+2Aa1BpTvGLJFSDAvRSb2Ga/6dWsmKK5i178z1oiYKe
ZQXMDSF7ku+lkJk7hQ1I1oV+a5lyFze81TJi/daeribLUQi+0sG2rJFhdX3bA7Rf
C5o0q0k58CYz/0nqLwXVJEaqRJsXQaRgxSQLEH3+YfddfhxXCDDxmLGRONkmgD/q
vTwVysKhLOwXU5kb4jL92E8fKweh8bziYiOlx+omWMRyKuskO80e9/wvkVUF99/s
h3FBNgxI5Ndnf4kegEOe6iXIMFibU8xYeU5jXuEQlUOuBHuNMzTnxBixRM5eFR4w
xQwnTfs6OG8nsMSTPOzjztKzMjd43XNHzPBHDAxfNy+4IF2+AOOC7NG/82Ieax0s
AlqMnsxsf7sRzzxC/XL/i7wa6DstPhxhEvPzdlnp1FY9NkehevVbjE4N1HSu2mux
rOvH5lgXZQPEryQTbQAeQMuGmo++7BYSx04kHoE+BJhaEo64u1UVOTV5ph8zjiBf
D89qGp3R9BYdLlp8K6cu9F7Uv/felhW98FB3ECbvB+fLNT+d/1B5eJYT9gz+B77C
9dMWo4xcV10/U8ENRbvX2tO02j0+wsi1RbOXlITvpmvgY7qKdjEazHgw0Hvp+Oox
RcyioSP5CXRnydsMCNUuWb2ageyR99FPCsuKsyub73W6DB7k0kRK4eqzbZe8BPhY
wfa7N0gcq7M1mrjBEOc1HwK0xkt222cMz1dGrao9uGdC3eupAe48qhWCCPHrAAtl
FGMtp6hbi5NC0nRrrG3fl/ed8ixmFOr+YwAylwsVE8vC9UwkMs3l732+IjE65cPU
b4rhqoIpy3xwVKmLeIG9MmP1TZpSpAy+jWgdp6RYJHnbVakHsiYSUe64yqOCCjj0
61J4mMZZPKUojRDBlOZiMMLdIxmVrUKs92E0qT+wPEB/MxV09oXIyLBwjWbHvqNY
3Oz5JTmBdtZ6lDAI+B1YlrhtURHSDVc0Syhhcgg5PJ4StXnk6wzNizXwY3quZFDf
cEjiD0f/gR6k3ub1W8wtYUeYTTsCkkSfRWdfH8tUDcBSLB954KqJ4hfujYG8MwF0
eI47mfIgd64cmcYbvTLSCWAWpOH3Cyro8ggfNk7YZExsojDsMV5BReYsJWIjEtSV
IdMyNSaEt/W2GKm9GRP4omYRi1D5eO0z3hsHkxiCQFokMB0p4OwZgJctNpake/Q3
G55tIEires7zTA9XYovhgGgwAp70EnXt1CewEG6VfZmFxs1u1yur0qZ+AvYk+pHW
q2emh3ywr65R1c8lVuL8UudihHKAWXZ00hwk+7TLj4c+suVzg0JXYnmJ/pHFHZXG
JpaOWHIeeLmfx3swceudx/YSBES0bv1LoDhEUbOEsRswvYCpHdrWHHaXYhhRQrBO
G9vrfjQnl8NJH3PWVaZpKiXyKzcshBnNjsNb9Qll8woZYdFvguyij39U8djXHltc
5/M48USr+JmRabOn4jYu7YWXq84hGDO+KxldLCDpTlZ/VsZQKHnmDQV22cyAl7Dw
4Z5Mrxm8LAUNsZ+VPjbEPdhBB3M7XrQY9hxWoVvA37nbvFOw5X0ceQIgkwRWT7Z1
579iIc9yJuRXw8q3Ro/Q1zngRrUlGbGQqfdwZ77CiTeY+x1QH/9hkukXD4Dk1ojv
RW6XQ+iDlURrUhtb3rUI/YN1blp5LF2UCrcvvpJtim157jy0AFEajtpOSUCF4ObQ
scRbi1hjPJPsnOvsRd/XweWegIb5zZ17vn7RUfo4cSOq6mLeXNeaYA1dpEmRlONh
jr5IEF5aszxKpdQq4dswcqJb354QVzn1aIjrS0z0hHAdVeE9IRNQJUlYkCqJ23pC
YRmR3R3z+lZ2xDZjmnmkGYe8fEN0bHU8ZZhfHrXZd9BkXyKTriCK337B1jp2G+Yi
kIyWErPCi4SmuI6u/iCulqTTl4C7l663PX++HVOE7LFXjNa/xmb1Giyc8tJwQpWC
WCmfXF/Y2z0iH90PQD6+TAUD9oexsE0Jp6nME/veS0ZAuGlQ73sP3Cb2xaabBIg5
1KvawYHky+HB0KYhHGcKSbsW1BQQqzIL3cwMnP5c6sAYfWRnSRBEKBke7BTwvx/9
IpvOWfnlkKBDuWVrZacZw7TzIdRW1NgF+lr7k5x9vzPYqo30jK/wWrAcgZQbOGeP
BoeTm/Ps+IsMCeShzP3a8lklrW4JKGZChErBPokiqyXnTaCdggKvTyoYm6tgnSMK
0S1PFT85cYHN3STTcM7q2QwNVhJ9Y6DVTqhCxqTvwJ+m5A6YKIOAnEaLt4IK9j7/
mhLwfs5VpFmg6DUTTNIjn7UpAi8yF3hGz4yxQ3cSa4NagVlkcWZE8vOCjoPNGeb/
zqdqzrbVub7JKrnOgJQrnnSFSMaS+lccifOIUjnQQqz9AzO/5daAh8qbIFDPeeey
pAUY1v1fh5CoMb2bl6v56bJGet1yxQNutOSLj7BWL92ZywG5rbfMMTCYgjC1+wnD
9uig38xErifEoqkpQRAp7TOvTaa/t8unB3mTvGA+cs++dYMx2fu5W+3AnZxFrZ9e
OgudFk0yatcswd9wRWUi8Bma750hEHQLG8fdZfLUXGCtXGT4QVh/NqYz/AH9M7Sa
+OSwamINLcmx7oMDpkv50CfpQtr8k+03EIVJWf1jZDM9ALfeuuh6m9S1RQd5EF6+
yVwxmX+gZZ+Y77JfbxjP4QSxYY4uVAZ99RdV4gLGMvCE+YZhfJFI3qkw8402lvIt
8Ry/A+kCvpED8EbZeFLZI+Pkdv2cXmwahLnzMiWPEC9vbNu3mRhd6mS5YW6izd5R
OuWV4hdeDc0Kd7gLkFrYOjZQzhZzrdDG3UY0S6pp9LGQRQGr0xXDbrC3CzIthTkt
bltbwAWoH+vqMQXSA/FABFdzASF6+0GMK1U1uERIUZTz9TL2Vd3DliXQAfutxcA9
1Hn8wLvnZUUGbXOcZnIXhOPJ3Kr5tCWEwjf0o/iLlnmtAloPLJamIU+fE9K+yqfe
nNM6CacNrlOtifuwHrFPUWSeT44gFBB1ucrKO04lHgvVed8goVmzB3L9XnMWPgvx
qjdgPC5WL9TkkOnPpmsi/KI4gjYuel7/pegzClB0eCMlQYjRR8CTJ5+4/i5AI0F+
lQbf76/xNy2D+0iuQrc8kZ7v32d4Z5I510kZ2ZUbj4ZshyxTvx74yZZ6cfOIm+Ia
U5QmFiQUj8Z7uct9V9ljP4B1HKinW+5BWDzmPKPkg/Ydr2o2cXl7mC398VOmZsH+
SruYaKjG4hhMufC04DJ7qlZK3Cpmt1sIFbdRHpUIbE8qHiOGOm6hyCQjLEyBZSCX
2TIVxoUQDA+HZKj54T8+CfZEKRxYih+pqvz6ssGZcDEY2pL77LP58bHaslvNjnNa
DRC6s5eZuSG5wRUDB5/hILcFu8a+zHHp89Fh0gbBV4+nFxgQKD9bkXU2UI8KAb9I
m/fyPYbluttkVzq7UYEQRGTeT9t2qTXCljyeBORaVz3i5063QVFlLvpLRW/6RRLQ
l2HUGbqUznUWFUZGPyJe0Cd8hduqVfRWfLRRAv+zfNluNeBKht96ZAIX4wzg0Th4
cR9xiXopRv5nCTs0kLADpvn4JkoZYe2wnMLVKkZyTbXFO9VTJVaXT2L9lRHuJjuV
qTF4rTZsEFunlYU+A7+WnRtEeZDOwf4U/91Wx8Tl8+jek3WwwIM8Q1RD6WZIagHS
IbEteBNIRKvVTb0K/mx7zYv+uBPg6zX6DGpWnJYGyWqWSxDRHxY9WNR/8UOXZ6pA
R3TxQTBTc5qo5zx5IFWQeibGkiKl0lHzo+7WXEClzcbe9jj7ncZGkXEbY9DuKtYp
/Eskfx1zHuAb5ttZepiMp2Oh6daIBV7WAXvpH98A8SVzbah4fR7vUaDAZ8WLmafl
4BcriVkRuFXzpjRWgE2ibQwju/qI5rOJzgs1ZPu83OjUHZNdacsFBp/KXOwcGww9
tv8XUAy2x8syzkJM+LZDj0cl2YGXmbf0w3WoMVNo04ZEy0G9Q7/8krSdoa4/x73M
BksjecXB3ubpQQxYsg2YR+yDYOYsKU738SW8184NhJxUkmMpwoXw9/AIda6+XNSF
QxhyiMi2cfQPn89aWmje5mwyfO6mPbXW0rCHJLHXZsUX6hzeyujqV4f+azTRr2o9
Q+8k4+m/2d8KIzd/1MY4gRRaOs4xS/2YOuT0ahn69oI/i7sZteOaK5qVoumgVFdW
FI/TdQybwFjCuqvS7RAwq3Gdb+5ZtrgVI/pVss2oUBX3FGf/iAC82k1THkFJ/IWo
6bJIa0cCmtXNoIHBVtk7GKfEgvmIuV0ZqGHo1WnCSlJrdiovjAriTrgYmPtJaKOX
qk1nMMFph4eO0rBpwc9oUWfhIRq/DsW4I/6+IUgUoPMN1/GBqa+Hj7OEUvZrtHcF
RqqAxQs/2k8EVPvCrlKWxpY7S23Q9UjjvJRbWZ2ufCH2EB7zeQv0yf+2VmxdWO/H
3f15Lt9Gyst2dh2mgBvQ5X7YJZCW9MVpbhHyfz9O/u5HjYqWwiXQjgiUWFybOATi
nsUyCLb4GnGErbaRVH/UQl8Wyu126eNZYf9UaQBwbo6s6dmFianSOZpKUvGSbtDw
JgN02RQW8sXzHWWHjdJXDpXc2yz7HIpC3t+Axo5SkDfpzo2XRMjiDNahJkPPqeHi
hFJU5LvgN3dNCG0zyfFQk+nCaT64inWLZa1IQJDiLwQ8bB28x8DXrg6+nXgL38jC
+zZ8RneqGw4O73DeFnXYEhJlOl4vQTsVgBjk55VHln9beekojCsQYS/Xw1u+Q9rW
C3l6NeB73MhF5MOEXeACUdmb5VsftdHUVIhwXfZIvu8mvvNgkmo1MpVRQtE0nFdB
4C2Dn7sZR2zYpQ9nQffZyaVU7hrNhd0w7QBv6hrp6bSL++Hl0ms0VVmrEIg4DxUQ
QoY+KoAR91egGNNqbd9Hed5P7hn07vMrV+C6YWVydXP2g5wX2KLaYaluC54w2TJX
MD/US/Tsh6Y/bBGin4dIPYdLHW5ZMI6WAuk7NafiREVmho1LTat9stYlISoqzvG4
tKDBIQPXfl2GfhfequEVPeoZtTY50BB6zNI+WQpmmR4phc4rWvk/8EUr+1UrzwK/
Kv+CLyKVLHpBDwXBI+5tQVwEeRezDSsdSX5vEGresrySfWR72HnWMJlpwbDwc4KO
B1t00Zxk2+vCOor4SjhStq3vBhMNBH152zFcawKsuh6Llp5NUbjjASomTHrLSwff
ivPyKlMmOcjFnplWKybA4eLeMuhn0X2cHN0pusITki4iLjNTKpqviWgAAD4ev00E
64kzKS1iwkTFkQ50VauGZqu2xfRXUMd1/vDFLe24i4QVp3lFD1TiRctAM2cDIUxv
qQj+baRSSTkcUx4vypYfOwSS3+snNQ0toSKrYcfw435QE9JZ3U6fY8kBhf7HB2li
GeRA7xyVL5AENzxEZ4IEbeu3JS52Nx1VRG/EerqunxBsO1GUX7GhQ6JpkP9aBOAb
HphCOO2/AaREETRESy+gRtrGlefZqHCo2NwL3ICqp86AJwxwhgjD9hcoPSVvCZVq
C29SMT1RMoUiP5eoFU72/GPlVI/elvz5Ux/9F0R5K0keYztNeN0EzPlD7BREp8st
Q7f9NQ2oaho4nIoGXdj8dXlEBqwfGXbEANWYmTpOFrNmEAbzOKQUAmKgCeYK2eiE
Sj2T9FBDZ76YbUo9T+WjDVlLgnF8nGTXHq4c1be8ntmyQ0TPruffXeAwGd7N5FvW
9Z0fy/kOAg42eD4tGbxDxfKHFPj9ocl6fQbCy/Tdg1mzd78oysvUggdYFIO+zBz2
hnELUHoA3Bs/wVegF+yaTxK/1lHnJsph+CUhiD6vnEQrWP8GHsX4PBuG8spP8MQF
Osrm/ckLqQt7xk0QGLlFWOhJK70fhOjFq8BHxvdo4vrwJsWgw3+iQrQ3trHvD/tp
4oPwK7/nA4OVhEolecC9MEVxhP/MY/Wspt9WaCOyuAmA0jteb1xehjPbeEvSkVla
bI2LikFPvVnH8+BHXyW93l7q/rX2aTIG535+6aVqQNI92tMQ1ekqNK1dQotORHiF
CG2ugE6xHGIvL0vD4oZR4VeLL0kKbPrGLJUdLUl6Q5BSPpVrkir/rCgSkNB/eeC9
FdF+KVP0eGG28szCcgomSRO9/Q48TMzygoq6hT9jIydLVKnHZCplUmySy9hLYHEj
DFAHmBcczugDaOFiKTbgjc/OkbK9wy1SHqblttU/BrWkoE7Wm8/+f6Ed/w63vVob
c4QaB5zIZrpeAfeZb77yMPzTZcRAUEgnQqSXQkOtMHPGqQwDaQw2yc+RSHF4ZF9Z
otTDlSilivlVOmJKu+cImjDTvG8x2MLiU+ijyQFY/f3k+WrMMxseI16Nwpo20yT5
CrpwDCWBU6nEXZvUE3bqSLw9uQWb0asTpti+R6WfzckpRc6le4QiUT6nAWnDTmD6
NQyAyXLjZxmKGbr79j9/BtrfxImyFRmwC6JM571kCLALLXkvcUjb07GSBaS5qmdC
MRAT/8QVrjtvA2DrAdcc8/QLOT0/B59QuRw7S3BAg5vLptJnaKzyIghuqCrwQqeP
dEBpO5j/qqogHfnhawh834XVApiZvF8429sIcBjuPNXAAzxJeLQG3s8QFhNfuEke
21HCAylOWUFC4bEuSuVIQ+oQ1kfPkurWV6GRp9qh45lMDuuuYpGbl7T0m5CQl6oQ
Hgr98USfJSplTQbhVzzbU9qHnTBqdkXPzgf7eMfMYC6UCnI5Mqk2bJmXSno6joWI
e2wyYIZMNAFZ/8xEFQe+hY0L/b/rjeA0s/uKRZMfKKlSqMqs7rGT0GAPCcdry9m3
MYe8r8j+FOjWZmlYJud4zBqs5z87bd5xm9Y2MqZFzd4JjGI5XwkhPZqHWCoJz0R5
sefkJJx2zlKOwyLPq0OamSLeP1S4ra7LnHLi52a1DCBTIhyrRc2pbkzmUS7xsBN8
EAN2t9t88KixZsw+T/e8qH7tjaHNKXoQvWsBzBId6jHl2pfdQPx1FAt2MiO+O2g0
R7dRuhuC3bENbTsOxrQLhYKH6hZnpRDxAxvQwLxJRGOgT1R2RluFfhnYC9NUXQiN
JaRp6g6xRFqs/Iy1yxKtATnKKMzGfdbXUeKpi/OwnEftOz+/w3/64PUZfnOD7eOd
9OmoVi2RjseP5qPblRJX2mOfjCFRgaS8kbBs4YR+rqKxAjQYSDpO3aOch/yevSrB
OO+ZTUWlcqfuQUxXuYQgQQteuEM29dOts9Gd7ydgI3n48XV2RWv8VzwWSppoKhKJ
tfyoNR60vCKTp/Y9zpS55jABbMhoa0mgBhkKJ/ktXRRZEXVZptLINxGpDMD6fOYk
eXUWnKmLXz0EDr2TBadpaFPJ8ZLbj+j2UkgI6AIT6nTbTgS2V8M7EIXyXgbNtX9f
oHZLhmRE7JNH92JJ9ATZbflE+gATZ8U+nMAGSnK75ud/fIvLOt1DTZbg+adjbH53
9q4eLD81qt5xHMJvc3Z7Nh2Cl165QAMsmYlUnRS+ofzXjbnRX/DreZRLRsbZd78u
kldsHeqcYGZUiayQX9AB9/IE3NPpeXCOG4GA5Wa3SIK9WXzBrPVjjnyVJ6raR7Nr
H4DXiY9de7fy5IHGY0XSzzQGLZMWT99p4GD3KwWUkgIshTqRKV9Y+hWKBomks4Vm
kcxalR2iiErKHChHfSMF74d2ETfhv6jKvFsSNXshU2olrkSx943V1DFgy9ufM7gw
isWahtb5rSgaIb+2tLjEU15k9+b5HdLaWvIWS3spG29i9NkYzyEj6rJVbZAA2Iiq
eBn1gqADFX31ed0D/bQzbEhxC+ik38GQjjshenYvhU2RTsaXXwe28PCVspgO4uDD
W6jaxNhqaVcHdfC0LIkSjPSmU124M1tnyQSnmHhAeEUFYfflmsXPL0j6sqnd+tJA
ka13+rKhQ2pUK/DiXRXIvi0cyghztvld/PUQh520OwTEegWT5NptPkSvwQkElBnO
iotfCvanOp2ZaHaARHYXZ+3WkUn4tfVN3g6nGO7UxXPwyHgrrWmPduw9cjV7SGJ+
8QM7mFI7nyqoYMTe1zjkEHkdkpJQTDQCqhIVyBlOnKZuX2k8qD/di9Pw2lfjKZgk
ehuvo5kprJ5yftooA0l4ThwHm5Yianqn8FbYtWmeDOdH9IWMoG9vgOLETrr8lNfA
0ZGaookQJpT9fApaymwLTeFVN58JyijdbAVaMwHO5MUBwcn2dWtsajdCubjkQrM5
0XcU/bWE8DUt/MzGNOxfSl3m3Ojv0q+AKYNWhFg5TwOL0guQIa06qmhFII5Lbhp5
FbZpUDAPVDoEb7zRM3s0s3Y+Hl+/s7klxnG+vBHfAcVZExKgv5JG6QS2vvWbRjz5
/VrlMBbNChntlnfOLSj/Oa1A2akyXpg6s3DQ5D4P8qklMEyVkxwTjFjtcP8mHJoI
YCoMIHqdkDXo7xhJjWm24LMZgSo3dra1/hWoFVG4eBd4rgvFW2vc19bVh/QHLar3
lhdH6VBruvM56nY0hnZM/UaZHJuXtzEOmF8MHIEN4yG8Dz9802+pBv8P1MEI0Nr/
3sVbq7exgBnxFQaqL8A5hbo9MEp1h4UQOvZAiapFjlnI+Me4zBjCHHK3h0wZ8w4I
Wcx9hGIK/Mjgk4WXxPDq94YNlfawt0FefN3OreCIN3u97ucCzEq2VpVhuyJP7YVD
ah/OSBHPluWzXjHSgQz4H4x2QY3P087s1OabpC8Z1Lba1OJLVfADQc5CEEeqoCmW
FJpIDoBAoZWHus7yMj2NLgzDUUk3TJlSofbBxpERkyjudPpAqeESEy6bEXyIxUmI
IBI6l2/MRH9ptyEK5XRbTpPHwuiNXrtEzbwtf6YnDL7twdcUs36SaUml3HJ6fF3u
ZHMiCX6y2RS3fAfPBgar2MgyBAgC17s43z9dk4qJ0oQ5Bl+yK5iv42GaNCnRGEI3
J3dH7QX/g2kYR3Ys1nmlSug0uZZ9UiNdxdFCKmUDq/48UAqpL4TdqDSrR0wGF+O/
8gPBIwASAPgPo7mRXbb37vSnESzxU//+/7qLrF0NS/zicp/yFFrSqNoB7jKgixb8
j34UyrVfjUG8BkXXvVX3E79w/0cqhk1mpRuxmp7M9uNjRh/15CcStxHF9OZlAznh
l+5bOhe2rERuK09WvlPlekJ3XE0nYER15lxGEJNQBe9T6rmjyJOWz/PmYOYq/6W+
4Ve5yVG69/pMc5XRWZjMkApu2q08BdyEUO6sAlhXFDAL+Va0IH4aFnl2CMHkMPzk
exfT7KgrXZMU54TzOThS8CtEZn49wYq2m5dbrYy5SHN8S6Pfrf3OJ8iSpQJgZKCQ
dyOxQlcQMyE9R7IYPwSUSpZC5ifgkuLKSDRdkOorIKxZ5nRSYjOAfsUBu8q4MrmQ
SkdPxwJhRNM8eCVz3tQtdbEYD9rHdjtrsIhhhW08Y4Uv4uYWeFUA2dkB3IkOSB+X
tIqAyJxr4EBJUw7VXUmqjiAZbIRY7P0sX4bIVh84AI0yaf7P5B2YDNdiWIGK5uHn
c9Xn0JqsgTVjo0j0Wz0vZMtaNL6n4EKrP30JMMhY0DAhQMzhYpyPwUaveqzvwBLP
0DRstWWy8CnxXTTfMUw1oCvKOIc3sZtRVlI1GW9bZA71wGYmmUMXypRn9RZKxV2i
IXMgdkw+R3cyS51Reo87pC0/VOflk8mTp8ab0JpGLG6t8cy9L/dy3KdlB3J90aHZ
LUX4mUwEXN3Y0dLL+FiU/GtmgawnYl9r3jP/F43BNmCEOO8LWSgldsCYY1Axjg9W
oTo4cQWVi6pkVeMcAgWX9XfPSTGBTkqXfGZ6MTKbyKZDJ2jUx8PLcdwKUpqp9shf
oHXts9AdPtdvoNmwjbo+o4FNcgYJkVPXeFGJLFD2Kj/cMV7pOevjLQ3U66DMhidy
5N5TTxReX5ZFp9G2wJV75MGblJc3qQ3koDVits6lxlW7KhM0ympozlqtEOniCA8P
EyxcQrHaLXouS1VLz/gXzztCLLE1cEiW0/Ls146KLmw2P8WJ2+rd9oeX6SBPYlcM
8Oxn0muLjkDG+rO9JbKippogUJbzE/VymaHTUFBoBRoQSg39YoaNw1/oLKs9Qg6L
lhP3dq39p2AHYat/ZnCiOYsXdM48TFRB+GZNfxBXvjCNujSRDRf2ryuH/XcWS+9U
eemh3IadPWEOQAE9wipA1TU1kmtQeogPTJ/Qxp6qieMsl0aC4NGZzzmNu/n2jyg7
reUOVMqh9UeyYO0NyYbRc0NorPN7/FzbGMODRY0i+qfY0CJMMh0dQqImdP4GxnG0
j9+vFecD61p3arzusiqY1rpg6OtqlbUnYedVrfyE4LcXB4zPsiZO35lqtIVoEAYc
xFa0DRq2r8hWINdLKc2bqyFEmdn8v+X6Fwdzlc2Whp4zifNZsl+gYtVvES7Suytj
8rCSfwowHVwYLoWLSNqwGQ5tpE70tFJo9+iDvh+sz9kSWx1g3Nc79oAKmwnLiEWp
0BOz5O3qUDSkJawRggYwi5qMsidA6EWknGE7nddKh0pijb6fixIagRURvywRe5/I
fnfyz5c2yB7shSfGIqNUNdK7OtLwMdoHB3tfnTm1U5yzSEgQhjLQYp2MbmTIFMxC
yjD679GwnJyZQhrS5+Ew3j6hqwxSwnVSPkG4UXmjbk5TA1BcMpjt2d9cnw+aoQWb
oJFhET466Gh5ZdZVORsw3I9O5OIPHfZBr4E+1xeoJ1IMX/zRwEyBdlY0Mf+GiTGz
UcrtI5sq9WUq6gzanJi1ph1e3AIyexKkG0ZfxUYgJKydyVaq+aKmjcMCZxwzsDca
jxHilC7nTO0qXj/Eo0uFkIrIDpJB0g8ZbcfoSlCCS6eiYu0k6qgu5u4swZ6odiGu
Q04XX/fDqeE63PQI2W12EvETW0kE9ajaitn7U/ioNeE00Yq5rAslJ0mBpKbPPeEp
NW6u6kJXp3eRvmr55hNgzDzbiLJCCD7mPQ8iBH/ByzNHooVV8hPSQn/RURT85rlu
9/R+490KMY2CtTcCm7Sqys59agd+ER5iLCJuLSqLoaGF+COgx3tqL+CmcOdtkj01
Whgtx3BJpPAPPpT2TZnaKANDGMzGm5l31Lq+lp2hA1vptHo4dcK/0LE1ZGf3ToAn
9awe8QBarUjPHx68bxIo+4n4dBDaGiaBRW7UpGCql0Oy7uIF2rHfE0kyQrWa4lwI
QM1VOkJmdXBd0U3K9pW7K6MYLoMnuZQpL7jS0tyhu3m901XPEZDq2Nn3bSlF8bA9
5o03ua233CgBa3Jwg+uB4cDM59rLqnhHzARoWqgn/MvSIlqmcVSYRrEGzrmrfprL
m2U0/6tQgMtds899I1+k2eGZwuK16JVuppKGLVZrF9/p7NtCaV52WJ4P4FB5WL9P
lgeEVPlt1gzvvN7tbefrFUqOAO3hC/3IkMIaaAVAkCxLnwv0cvyrw2zBK9I7OVdj
M0rM/DqojNMEu9lf7/HAGYKl5gPVJNsHOgxnXmqmPwNwl7Cn3Coj2zjietXcs1Rq
GkOEcigW8y+CRp8q/F7vDz7Y3ayQSBOh9Xt95vnI2Rcm8nUCEdarOq83r5kOTL2U
MI9zHTjnSX80E+V30IiuCxPLePuZ/DLCdd2ZMNcx+0iQF+I3eaiQbyjLzpdWD6p9
oiwvOzXq5KLj8WLu30cZ2UDDk4zDrZujOkof3fOYedretXqPFwv+LRVFFA5BUi/m
y79C3qKFOmis0MNc1VyLr8zScEco1FUI1X0UBNjg9wwoJqoR7Og8MBh5gc4rZ/UD
IttenSlU98rZDd/1dZn0MnyDdRFuDE53ngThg084lCC2+UChUla9cevIDTDgLsTo
ZpkpTK2aqO9ePe03bsEcBvnLn67QrBSOD2PiQr/FLITxKCj4/TqJm+0XTHhx4X9g
Q52oehyTfFp1l08FwXxo6pRNI87GPLUSdeoxiufHEl/QbO/CvFCMdWGdnXRh52qM
y11VDwiYgGVJnBCxwMiwbr25ejX5OdhWwFCRDmzvMIuxUjuFcOwnuFwSCaKmZDhy
rT40HMd03DzGfqBINkp2H0lzyQFjQaE7tMU80zqKkjQVeoOJM0ufssjk0PJ5UVRG
JZ+13lMgPnQfrO9srpKK/EEstDBBHX3iIuFE7fRosbwuLaS0sGhF9dGWB3uGX/3S
p55xx4iGeUecxZKaLJa1KcP+H3fjVs63MPt8GncTN4PQY7lXrPh/6+C+L1Qxzb+w
XHW5gka1TtRzm7H0ENclTed3XTcBU6xrWNUNJ7jN7o4KlkGWAXXxYFJiyUBYKISg
F1GQAnEp1WNkiC6g/n51XSisjLM+JopUh3D8KQ19+men/YZWqlIjIdwBLyG6+j+9
i+e2xy3/JuIsqCW85jrMMKyyOG2ho8C5ogaOZkYmTj7nJTciPoD8MWWbFpLLXFN4
`protect END_PROTECTED
