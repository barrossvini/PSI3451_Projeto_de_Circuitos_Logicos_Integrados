`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfxGkhaW0wtY3ZSdv69AwzQCUwGeX3XNUxhoUGDbR5mz8F9YQjEfStwZmx8IB8Go
q5Qgiu3Wt8AQ4e6eVEIepKfLxcbO3TwE4HFKziBZLCrFN/fhlXbeSI0zjkWOlHFj
RfV22AegHgJ5eE8n0A7qX6CQFizOeog97MWArIrndtYPTQSta9S5KfMxMZfknfF9
VnOb5ZZjBKzAMu4KIZD08DJHVYtmiWnm52rnOd4K/tkPE+8FYS+tqsZ7vH3tCmVH
2vIvi+Lx+77OjeEV6Sw6DVYqPbQHUwdHUdhikEoGNgHfItl9KSYWQBGdinIVV7Zm
pv3VTKgjKGYjNEOEevG7VYRXxEGzILsw50v057wDNVU97PECfG8AvqC3kOuETGQA
2lpaz+c5y7qHxzbJ1mnaHxR5LszsyFXlhqpIy3UAWiwA8Eo0G3h4DsL5AC/5Lbf5
yKuEI8PtE7o4fm/At+6JohBJFfmW8bg8Ftl+y0gXIqpE0/a6AmBH+c3s2+3HfOEQ
nd6WhtrQBIzPm84OKNTrArcU65JOL1AiX1Kz4ftj2q+fB3svmgJU1yOeKdyL+eJK
GRF4WnO5DJEwMHT9n91sKn7vPUAnBNxcVAZyNCMk8EeX1G0/1b3G7LQ+S3+jQVgR
/ieMx2EqRfl5KjsrJRGnmA==
`protect END_PROTECTED
