`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jBAaCEgx2UUq4iZ7yrilSAjgrHa7wabkGsuJp/wFSm2IhbvLAFjW25Pk5kgDChPB
zG0NOtBiGY80kLlcWSo5ncQGGzF+xWNaTv42JZLXN0q+fS6+c/KyX8EqqONS7e1d
8oJJf5K6orJ1VFj5hy68/sXjdTPWyUV7n6uCkLWFumz3s05eBTzYYlyB5Ka08aV+
F5oQN/A6KjqcERgl7eoQdKI0Rzxwvq5WHxTU/KsxH/wImLEcKpA/INm87QlmD7xw
7+uZwV8FWXqwSWPgbYUojEVTqJFTPcEjQz93eSn1Rl+gzVahs/ZNJAiPku+m996P
nVb7p9KZOmWitWRLb5aKf/8YbSWB/rVfKHriC2yXPAAcTIoWgT1uCnEHBtLPMz9i
ZDIR9eRfSzMczbM2DsBN4YvI54JRb1jLsruKpar0ixU5ptC6i+xkXAvM0KTiFXcb
VVg4mQIAVRd00JJhWW/tPF284JZCzSBXe7ON1+O9WjCbN6pT1OYjn6ppnaSk0kiN
dEw9MB5KtieNXGdaAoJaBySmCqxz11djrz3kIt3nmBRvNvKSfogzrlfNhjit+Oso
ozV7IeX6BOztMrrI9Qs8ooq4CPYHW8ATLwVgCFsjVj33BJP9BpVn4+0mgHir4GkC
wzK9G0q3Vta9IQo2y5JEvusiOdtibSQdiShpH4U4PK02AAdhCZnmslEyExeKsxeC
BGl0klDDeXC5ftXR2ySeKO9vUk0nlnLRWrnDh1QmCxmiL8dm9bJhBSzVJiPSWtOr
YRvmKVs2sAdViQKtVXHCl1XrBRrV3BkYtxlGjsZnBPUhqd0TGuQ6JIzDB3j+dWMN
1FlRQZWU2NRdKjODg64bBmhdAKtimhKwRd9wMXFXv6DyqK5SfbnEsRQ70FmPPYve
wcbY4kHHdiV/IlF5A5BgJ90bpyxZ028GU82AgctiYYF2rQYsIegH3Z9yvtr2PoZ2
2dBIkZrMJIdiv/wdMOz4Txsth5y9IjUat2U4nxT25omTG8WuUJSDK7sgDqyXfkcv
yUSfTALcmoQIH8eiDhmr5rT8vgui20Sov6awkazRp1e44RKU+tnnazoERWXNDHge
C6hyENrhZEBj/hUwWBGz7BKyWxZ1PJtXSZnMoSLagN3b2gPQJwk5deWYo/2StmDr
18wUoPfw0JHvYPIAwyzLTjgqCuIuKx8aO3Dmxvw7etcHqoI23KTorPLUKU+a6EEC
XToVOfgOQV8UnIYDk6cqMLX73Oi1OO8a4XZVqGNTNDkYHmP/BbndtYAG0Zd5pERM
PRaWhhIRHcuEzZiB5Fv0/V6h0aNBQqi1Xl68wKJ1LauXkDEu38SZHXGAgaS47xdJ
6TMMdQfnGLIGoqOIXPQ3cRWK3kE9lQt73VmRs2zdEo1bkppbGlerHq7zYY1/2RUu
lcylpHrjj7Jlkm8bdUIrSD8TyaHcN4iMonS8aIDhMQyQwBbgY39n39rmjGaVWunq
n4r+Ur98uYWcEY8208c6BGgpCystmH29P8RrAM8yW2LpTJswbj0w16epvX6wT0sP
kziW+r+/uFasDaueQk2pR2XutKgaN/ILH93LVzThwDpJnQN3hsgiXNI9U4uV2xL1
uzHZv6ovBI1NKv9tBhPdd1vOTm1l3jobhdtHrOJqaH+IuVmFVZ9w7EtoH6NTAIif
IUS2J20QMFBFu/b3+vmBAs+jjEHPPWS50ZlEe1tGFL65lEQpkqkgBZGfCH6Uyp0p
4NmuxRtQrBCMygsqT5Vl7hkyS77WAr96hBElUBwXw6FOVU9vmRQbzvgLkImrKVVC
gDr21oDMnEOKJ8jLrpgWvEvIemecZ6gyxQ33FV//IkGBevrbY0abW+nCy4xdAA1p
VTcN6ZXa1Ml8IfuYg2gim4Ixyk+CLap+oUw6w6MzglhkbwEUrsF6NlNBVrhZJgCg
eXhQVZk0fzp9bkauTtv7Q/cjGohRncem6OwLw3nsWgWVA+m0mShTv2EwmwhZsj2F
bcWtZWWKf/7PbIEhRADV+sOyCd3tPUJUzsEumadDW3fARvWN+zpHA/LDWBa3JHZZ
JdgXWZwOTIvWFGNk8IWzP+B5EdEKEKCtKcAgEiacg6UmkuKX/+toTgrVyfoSIsHk
o0cj5ofSjivtMHSfvNB/l1iyD8B5HSSnIPOykUo7+oX3/qFwXz4SerP9yXZX8Hxg
dS7Bprb5Ete+lc6dJq2+bVEGEGnsSjsSFr0rAE7X7CuPxgClwZJvquYK3+EnhCWf
ubPyPd51ME9Xv/Vyg0vd7k13F5Oq1Z5Z6E5QWJtdJPHNu3se5r9Eu17FoIjjTfYK
eSN1nf1f8L6Zfid806kvR6g2FORyzTyNE+TavJfNAxf0C2HMSd13jn5+K4a57SY1
5wIm+Q7TvwswbFAu49/VZUIaG/gsODvoLrqddOQmW6NkY3b9Aw9AKjvDqWcIzAkg
6gUTMcFMZUvr6f6GzPMfaCF8vHgz10KDUNaGOaZnv6h4UoJ+gpMFZnNmpYGJ7DY4
rOR+PQ3Dua6l8Y+wDx8mQLyqkrAfIaWiZCFx8XTgiEwYnIw+b/8PMsG0n3fsAJlb
PA0olIXKhb9cqjHxTao4FvBglG9UX8bDB1bq8fiusg/emSiXgn4NyG70hhIpO8fG
y3AjCgvGH+PNVpZ8UJoxHFBxbHhcC9zcgaPrjAhst9+PAd1v2o1U9F7kNN/t2c3x
DXLhlfdFCSvv7fe39lykzXMH5Vg939HUpFM8MhujtUY0IDnzHJCbxnIP3R+LpIyw
NPOw+F/hhvKUFsEjpHPD6vNjgn4xQVNYrN9E7E4Sgyf+73pVVI/ZVXjDnMZJ+R00
91uBFeSSZz/1jZp3sSUju1cHI8Shf5XeE6pXgWZP9Kx7HI9TnqjSdrk3vYLxryf8
D1f+QVo+Yw/pmGrpG3mriqXvIYBccYPjuBGwzPVM6PPsI9cSyvhV2MYMoVPUSfar
E4xJlG9PwmKQm/qiaHx1fJJAijFPUXcv4Gjs+f77Ti0dqVsU1nk/wARqAgUC0zdx
m3bA6xbp1287itCFnZu2B/I0vIHgK4+XaDwyVGGd62noImD1Xo/86Gnb9gfLN+5p
U2VluHHuWc4WYkmSeBPq8PMI4ninhUvnonYv4QuVdo258OTzln1TOzvwYjkN94Yu
CIgli7zhOtgONqrk/BjgWmICB1tu0wXUOpK0dJg5lErOlNubW3ZCU8VMvlSRz95A
PgHP3S/GpIJgrZ/5orSuI2S2FG514FYHuGf8H4M46si30fmyR7Mco/DjjWrsyY26
XEy+PEiv1xBVoU15rapQKQ==
`protect END_PROTECTED
