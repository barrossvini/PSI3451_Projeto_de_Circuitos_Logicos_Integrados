`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmQRx1JKCLXCw2HbKfx3VPqn7MpW/q/1PGbuZQv0qT2GM9FChnzxBa0l8WvsdNLN
nq9lIruKPZggcX0RfkyAz/u5+cMhEjvS/wZpSZfHj52f+HV22gtWNEHYf0pUDS4J
ZpAdcwE/4IxolJRQaDg+69DcMK/2//Jsr23V30mdFTfTmNyM4rCcfQ2/uN2XfMBX
yMccNH6xqNeIXeEFgiU+rIY9dDWpvhBiRZrvfrIrmh0nZcZc+aBgZ0WKera5xY4f
IZbUhVZ0q6EstWkBsEclGqnGNa1S7rwcG5KLMEpaZ9p+w8xyT5f/+XUYAkMkRXaY
l6vxBbyMW/K/3ZsklKlFSiVA+04fO9cfts2DI0MRgb/9YC3qkAqCzpm63eI3BKyL
9nBrbDg0hcpwej23f/ZbZ2ruhYWeAwNrA8oyYgcZgloik/MJBT4MLXsMTUNHv3qu
zL/b3sEBL0FULG4SZKgG965U0m5POc6QAd4DABQuV6oNJ9lYmWBiGxXI2sb82ZUK
IPplt/Ij2kHkZZxoHbuq0LPMrOTyW6AGB42YNr/+XOXaQIpC9fOUDjgyWyGH++r2
6VDzBNwvX0OSn+baISFg4wNRSCcOwV1nRNtn2xHo4jVPulFoSRvs0A4wYHAbc2K7
NMI8VElvuYdKPUPY2vVKQ3IP4q3jtju8FJdFwMnQBk74AuXVj2uDXmYeUvq32V1v
NmWrN9bk0amkGa+wZ4M/zkWaCQi82wX6M57EMlshcw0mwi5zYCbJe+SwZPCkHDIh
Ch+jQiljO+jqnlLlQpNlG6yNLQTw87hfPdRWI6wU5gAjY+9fMRy3yaoE2au81Mu3
hFne8n5tc8L5eCvJvZtxkRP6AXEfyBwALZDp6s4XIAtRGVV81RQc15ZUvMU96A5V
OpuGOQj5lhw9jifbT3GzIti0qUd2k/2ZmXENYAmkbR23OotCNODe8hlCLlbPyxHT
Te6HxgP2sVyySDSSKMp9+s5e2RTTVBWR1Aem5mNCiJy1l7BX10lT86imZQekxynY
+cCbXny43lo6dR/nR4axeo6ywVLq8iS0qR98q0by1oFabPeFod4gVlVvWAtiu8K6
ai6CvLBTcahqoytdWwaSDkQHUHpr8+Z1N1N0Y7RaqzmTH9ROjtfGgGC+SmGGKJAp
bATFw6vpsKRwXwjI8V7kiJKMzrx7tuENGDee8FUamOmiYFeo77JXZZ3zgB5BA/1p
/vprNKWdOwULltuI9EXEzTGxrG0cWJYzN1hFfQbomTwFb4/aYPm18SCPZVT0uVon
Xn60lkBUOiSFDnQRCKHfZ3gx+/53mIb1Q0+7noo09PwgI/CzbKi0DyrY1CS0hQLT
WVSE4/m7B+8x0A8zsTmrrhMHcHe7qjLy7IsjwSW9Kdpn0ezyQaU3X2E0Oyq6sWNv
u0ZxeBNV/a9MBlVc9dqYjxLwz5Tsn9mvo4oG3IA/X49rCo+SoPDcqXjTRr3zSDiR
DgMs1cJrbzhYdLaeNW+BJBlfUZnetqxmU5f2qaToS0uq6I02Gn6Zi5mc4KuQRuOi
Dz24d4PclTAZPoySvGlr9dxsBVfRjQUwqxBQXSlZvOaVH+jllxA8PiP46E9OQZCv
/7PqcujsLGilyQMjjqkcVr4MDyrDUPg/adgEKEe5ms0=
`protect END_PROTECTED
