`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hPDPZdIqHLmA6+efiU3b7/bXdFPlnXg4pymVn81jqatHofhSXrc2zj2udG67BtaU
0ZZKziIq7J9LukkI/KunMzHSKOmU8VCRdxpcoBJy2rVsBfsxZY2jioWQD+yZ7D1j
LsSXH9ihbFgTQJIPwbwTD2ziYVINp1BLUMIhxYyUqzgmBkZU6BzCw2+f0A6y7ytw
pzrXRHqK6vp0xCwxE8exFX+f2h2mqEuUIjjLL1xT9ri8G+gCx1UEroivUKtsFYfk
ZUGWyJyOgMx4k1zi56A/F/AhCNaPS1h9k0zE2+Eu3PByJKeP1hfBtPgv8pxHMdYI
vcJu6wF19Jjqjkw2Qj6j9hFsp8m43cCo8AehU9mteMDVMmssGhBmRhwbjhPWk7Cf
BLVr3ACYQNivS/3UsuUd/QB7pkJGpSjEP7+88s75nZblzsaZa+TGFVD5MG7ufMcf
zi+8pz+MYhTW/n1x9tBHzW6PKBA/sRXKHbW8AqIh4hRfaf77qgolD+RFkQSjq5xk
A4F2U5qawGHuYKjelHJ4cnvRuDUdXmKpFNN358QynoNHHWURmA2w24dMhx0XARt3
zA4Pn3g53uB62JKE5bBRWH+FbBh2wr086djKnuIM1hpfSF3lFsG0TdpFXSyzW8d4
fYyjzYmd7oORLL5A8dEujuqX4iLCZpugECkrUCq+R7Qjgwtmxoe6i7oEwf2vSkRn
TAk/ARZgWj+9mW0rGWXQ1MBsJEjvQFOUfV76PtKo9V/3RdpvquYJrZHfy0t0UJt2
M4MnqwbPqujsHEE3rkuz7LLZxEPi7HEx7DiAV64svhp+1hGH1xBy0utzGPGxUzlZ
O3TOvIkWScNldqRgSz817HyQpVmrK8KeBVpl3g6TaeIumc0YociXXvUCQpRovQjP
XqYcCsafxGXweLnvzV+U7m0E+Z2lx42sovgdR4Oi8rdsqZ+LjQhzZINCudn1TQIv
+q8hV3MZrVSCwskcPcOHtSNidnVyyJsmsV9rwodTp/wiruYU4Fe5C5U+sU9rTI2D
WoDxJ/Sb2jUUeaVBEU47JHejlN1vlrNtu/RlaI3friGdVmMBWh4ek/5guMnQd5WO
0WfyKyNtKucOVad9WbaJswuYt4vHEkk0PuK9U0YDderZEcQry66qnGyAFcl38D5g
0vCSq+CMfKjx18ifXihd8aVaRCcrHV7YLXeTKODdjkVKnNfF4LltGFkCfZthWv7N
caM1o/GC5od1sJNO1crma2MqxlSdpbihpcGJjuUAnWfyUEwNZNAtjDaD9Tn2u956
RAAdsy7lrVh3j5naHPyE8hDdIpBIbnNKraVnOTcpEfJ7QiLqw81ALN1HxfFCEtBJ
hUpVU2xzOLA6cn5S7Q8GoZKmia7pbxr8fL7wUPsnuZi6uXTcaXyfxBj8tYwZUlS6
oioA1qVNoyhYRpcU7bThXPom+8T/wjPbYAcI8j2aY7t6qB3rFfugK4G9XfiQfPrf
jyT8rxhDWStdO+fsPmKPCD5LXlpZetB7gUAYGbJ9bHPMOhNVaJOz7LjeMbvrTvAg
MO4feP5Df5i+JuHoxhv22lNgHWDWkaQBazwFTYhB+WfRQYV4JvAWFznoTnrAjL4J
`protect END_PROTECTED
