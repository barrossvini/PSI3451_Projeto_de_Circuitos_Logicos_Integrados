`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wvquu6JYK1g/B0FZhAGt/iipIc6TGwxELksib1rLVCNfNeYkre7HOqH/hCduUc8u
5N9k6hX9kpC+yS8HtEoCeg69QFSG+8vwabHq+TVnCf7EIDW6LG66eJI2WLcMDAij
8s2dhAUq17rVl5+8CkNpjUmfAUJSI4KMQTPheZ1fGNxD642X04JC8Lb0JrQe++uA
5Tq8+a97vM9xPo6/LpvgQCnBaBm69dUj+6PW++Z+IQx9/rdQjw1prA50p2fhnZlJ
/crebhCi1k+FxSMVen4KWSvpl2aMci72yEZf1toN3jX3R5chcHd60YAqtwPJlJdv
jgggpPtPfLI0j07CS5JTmqc+/hhgR6PfZ2TuVxPTJargUX52dSiAkesRrnoZQ9qW
VUz7c0tSQOG28aCWeECBLgXZH37kTMwVYt03X+ECoi5ySN4MFPV6cCqweNGQKprd
Tt3wyzWZ2yM1/PkWsigRHzIi6XHD7Ch02jKHCxAdmEe5hmac8tIr0cDrjCeU30TP
ov6PBmpC8RSDvQUaWVH7vqF/MR4vsYnP3DxY/gsQ0u6jJWXcHr97qAOrHmKSlepW
sIebMW4AMvNxq82zGMGYJqT/Wih0oS44nq1WwX8cGMQlmhe+jz4WlKnhD+a3oLD+
vpCHPfdO9jI4wTEmuSqc5V5rYqLx/vrP+2g6S3h/WSnrQyGCwGNTTsLRmVzSoRle
3vyuRF6uyOzhnYbYvOEyVvD2x5BjOimc+i+aBOnhzZr5kYoI1nKUDW1d0G22Tp7B
ty6xPZNtewdpTXU1YcQZkVACRyRo1RuylaZb7SE2tPCg5RCFGs5GxoJ/Ku6VQXCK
s8eGj6m/hd8QqYLos4IPH8q2StjScXb8oUX3y0Yr8U8db0AeH9Hhgv8rX6usSMSe
FvOg+vJeHCKYmYf7lhNNgdTg6U4CGqx+drZzvFTDx3kju2LELTvERpw4W8qk7oI+
tP7kw2kGEwiW5J0yASh2DBgdqJVbCdbgv4aSO7dMknbpLDovK1YR0OZk4OFvU55v
VnQgQ498H5jdUkecvx9I35mTtO1KEDKK9e2IupdcHnN3oRpi/YwgOLyj0oBEFQbd
ok750aiv9hyq1GjVEfxVekqcyxp386yMvDsJ7E/RePQTEoCnP9d/NP9U6qtzRJz+
UUERYRANIiPTVQwyPc0xNf1RUmiBkcIp54KqAMFDSrl3MfWi4PHhEqw3aCRkHZ1D
05e1eJa5yyQRzZchr9MHw+OhYfBv6Plf54AnIheSCVZTAM9Hgj5CQPkRHqGsCcL7
Pgh43/LW23b3xHonMADudZSdVlFGhHoBtU5trn+sK6xmsKZaLVNho9Tlpl3J8FAg
lGe92eV3dP4poomWgqV548a/T4k3nxqhrDhs+1oAhfNeWnFVgXPjhLpqjqZWcCix
wUsIvTvppgNwLDZpQAmZJYakMqb6DPSxzmb0K8xRbG5mBhHmv2yASPxExjvq8Vc1
eLz3+QvA+k/Y2kJ4sstkm+JyS5rTLlqcHj4gD1WoKcw5FnWXBAGKeO1KgNOCQ0GP
IDNvth7v0inYQVzyh0zW9NHolgsyXdiQ5GLOWqaxUSTHJrGq1F3S8KI4Qp1bPT8h
xyBPa+9ri9EUQNuixvScCkciskJWwPOKIA92jc0UavUouShnRhXaWWi1qN26rO0u
+dCGjfuDX5Nbq4eu5TAA5hiKhqIaVuV1qc487DlnwEfZVPlMcw5DLw9ncn5+MsVi
Lb2hyJSIn1d0qQ015Mb6Hz1onovOTZXB69EUTTcpmJIkLL6Rge94b+ifjulj2Pbm
hL03izfNFsYFcBMEtibLszj4dFf2R6kCo9yfAwuiCPX1/QNI1dc5QciZPtJN9Bc1
mJWTW1e43fEUdumRyRpyMzva9HRUscCWOhq/T6C2M80PcVIbZRrb1rhKV0RQL0TQ
pWg9O4FE00aFxcukq3ucRJNPOam07mTmwmQ5fA/9Mf5nWpd/nnY2A1BNWLPa9wdc
dEpwHmiCJqVUkR5p8zh6iuSdVhtKi8hYxjlmOK5C4Nflm+iEiqP08ccmF45PNgOJ
Pz5hXMr1r83JxL0bKD7EjJZ0ZgQogFUyXYddC3M+DhmHrXlRwYZgm/xTPPtl+TNh
IYINLb/wKL5Xt/HUqQIGJ/NXWWflDz7hNdzi/S5+oK4FZc3FsImqveCTId3Q1CzZ
GE0KULzAVjww3AEstTyK+Fw6S7jy6VxsFrirjjI1YVUBjuJR0+73DY98Tq7fjxAV
48fFZK6nqnkmpEAS+w+47DdsWeRDFZthbmnVGizSycdwo68GtffvclmNccmW8goL
sVyjRrw84MGdspYAPc2xEw+In+5SZNgDVCq9pe63cqiaNUr5f82irLVraIqY+y0y
aH8lMF8m6hyBZCTTpKbv1gpQa/pxxZYLogJIHL7LIr6qY7XemeGPFWGJ07kDQ2pL
sATpw7Hyhqk5b7YDZvyPxLXqdQDdaPsff3Vdr7QtQAqLURArNWIS1sRvhACs3tTI
xyEp9cmuxJq2kKxskXngsjqnrHzyobk+ro4i81mJieTCKiKG/wpuH4fQDhM4kN8T
5xTHQCsw6T1FrNIEq019c42ykicVWIJYvm7tM4uuUCTskTGjrnNPOT+73xV9PJjG
RTz27sFlh6lZ++vzJ+K9POMg99KM5OBk3tl/ZecwkjCJFr3rRheFuV32g/4V10tz
NO4/JkNifV0I+z270WaPvlP55XtLR0d2xUXcuegnuYkT2ga+6w7sGoyOS22KHRIp
jK05g57YpjIQ4QfzoPAxOzzq5nKCzicVtn1wVvG1bPyFHE50iGy9GTNN5bJMee4g
LVDLHu7LWtm7+uenGNhBiGWIHhsBQ4ZNcg6Q3K4T8X72LgPFFmwfog/a83SoGCG5
ZHUjR8gIqALjZI/rmIbgfTCkDpfONZuxphXN432GxdsVeVJM0oS7qOdNYDfCh5tk
uYYfo9+GE4iXKs5SrPonLXnXStujUisvl+reP0ifAiJ4Jfm9HmqMVoYj6SmLHLNX
uEJJ38BzPNdvbnIO/psQ12MZhmCRIxFwnEMyOOZK0cV6ES6oUmCehDSKV1xWynRT
WOZaB2Ymvzy7rYvHQj9alurPMMFZJsNV16u/8yHjV280jwVG5DcsmSyqDba3WLAK
JFcd/2nfXGoxCajSgeYPgGA013/HCbvJ/d5AhqKlO4D3D9YYjyiHDUv0TmxGObdG
8OoRKY3OgfQ+Zv4jzf+2lY8Nx8dhNBi5o16sDLiGTwj+DokLIAT9kkU7gi8eP3GC
ujAKLhzJSmD9MSkZw3lzYyaKJ0xEwrgynKKB+Bk5cU0nS95jsabSeu2+Jxcj75O5
ljasB24OKe/Shy4+Ey6M3qoHJ6lfMVbhiBCGS+MSTdkQkDjku1LA4uxob8YrQKEk
CQyuaI+ZQeutR6+27olScy+egsNRGYQQIjP4wHp8aUAQqWNvrq0CIAcRo91FMAoy
BChjUf1Jwt/I5o7x7fatTvIX4yjdIliGssXwb2tR9WfxSjzD94gRLVsgP6m3LG3v
inO3GEfrVLC5yMzz04pNfNEAU523F6DxjXBu0VO/cD/aybNFCDbzd+Pro9SP1IjY
OpU2BQkYzA42JBIhPs7YypbQJnY5LLB5SCL+wPsxcGI=
`protect END_PROTECTED
