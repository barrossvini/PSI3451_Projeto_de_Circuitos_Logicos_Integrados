`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wj95LIS6V0KdYbCe4OeEuhg+kujaOASH9LP0zl9z62KXhHQ8Vhi7zL/gUXLuQrU4
hAdkqiRhnZjgxTgx00Mve6WzeM8B+sgvZrDxDtEAm0ebXrcXZqbngh93yPx8sucw
7YmlUvXQUHnH0f+x9yhsmNzra7mNLib5MVXnFZBlwdHirsJyIeGkZFx6GstluwIM
8PMc0CUn9t3L6TQhmDcRUYrB4QtsrWMciCIpTmTKWj4TKA32YXT2EqNSoepebz+1
iL56KWMkqA1jBp54ftDyS0DXma9pSdM0ySgL/XRmCMEtuTI/Tyfut1XqhvrVEaCa
yOd+qTsNb+H5hf+TTegxEV9lkC5cU0py1wtBetF7PnBqjNYSoMpBbEWLcNNpbeVL
ahiEHlwc7FJxWoXv2a3y6DGCWUDg0PW70aX7TCJ0k1GBS/AaRXruxi/SnmI0FdK6
dvuh7A2+9pigsMwYh8fOIbp1HRarxXn+xp5byNfl0Qm9KEpIDA3N0v1zR6DNGCI5
d2Hjmy8MtZJdUlYrnYB106+1s0XyV7vqU2+stsJgqqJBQrvkyEDqC96uhkHi9kXY
AbCmZ0/KfBgz5L/RtjI6JdjAqe4+kEclFWmosneDBKC7SS1+Ab5O6tOGujsie6LY
HmDDfq3gGPbSG4M9+cXgHSBIgmw4F/hvGYOd+OwQEAmqocjMiP/tZ6w3L3k5AKOO
4uK7xmbnYPDFHdHIZ7d4/VXUW7NiWeud0F7BCjwhlHZ3ap0mpN1tk2go1ZT8rMIG
PVgl8My3J72RKIOT8/VquZXbLdpT3hYD6Z9XcF2GnbDt2ASPFdM+RfEC0is/WV8R
L+u7YX4f4+40q1zmLad2pPal6bVYBlwMQjdmSXAjH1yoBIRK+nD9lI91t5rbQwCn
V+FhlV6IdjSY/28+i6dJUOyHdHGtHNpNkgelIu3jW/ohxlpxq3NvB071x2aTouis
SSfacQpKponFWA5nJZlLN0WLJ6xY1br6RaDwBNhGrHvRQJytC6qi4658FwzR9xXN
Pbz+iGF/5Bux9JYqRrFkWftSTGiPgTfkbB++phsuwn3/Oe/iJCHb+D43U8sBiIwv
vAn4J9s5A/QJ9N4AoyCW8CegOE8d64+0JZeJUIvoMOQ=
`protect END_PROTECTED
