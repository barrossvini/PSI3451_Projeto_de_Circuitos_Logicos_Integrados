`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3BuWOYHIx6PuERYi1ZqE/ljz5AoFXf/g6m5ZNwwpGh6FwaOHrrSm+eR3HvQgAioI
pEDov7jQdeIPymlA76zSTrHl5z9N+cvRW4wZMKZDTGQyScmDKKNNindCC7ssvBxj
Sy6xTUa9BPa6gEnutqS7C3e5oTOfQQ+E96uZwFJJgmDjOOVT4Kooy9p9Ib3O2V7U
ZZtsshyAvUPyaGWV0y8xFeMHKsZP/nhrewoh2GanXrRGVEJR+6LB4qx0lxHHRsj6
frZ9ouB8+l98K5RjkVTNgseyCYbt2JY+gf9xVDJ33GEnB+3qAXVRwnmk+nNzfmum
2I4/81SC3qlf0saWA9J+QE0C3b9x0UY//Yri204rf9bT/lBqkNYv/cwOMVUQDw7s
KXfL4qXQj/bz7/iypJZBgUaj8zkvXWnfTLtwzCuHz2HX7yIEUaxIgCf8z/3IwFgn
5He/8KaMvhgwd0k3xYS6TThiqtz6YdDD/MuEfidsHst8SyyvdPj7c1+Ao1yLLTfL
6XHjZdMofnRlDyod36M+S1H5FnKQOC5ZcRo5/Hw27VDLoibJy/KbZQ7FTP8aqzHe
klEpE3D65DRqJS6zkIcY95WRFNv1CxkVKCqMpZHeJvN3RfqTJRxItrN546QUjsPh
5RALUbH2flHebrDGKSrBy9b4sd1T3Qm/3oEHXLF+IUDYwnR7D0ccVTnqgnUCCjph
OotZxqMY/i8pKrW0+P+f5wvcpocfPUyugkNiFg8+7AwDDhallR9zxlTwkSxXpj9o
jPcuFAX9NFO7+GticOvkpW5Kx3JZy6HeaVhZ8jPcZ0bdgvgSmGrECRqbS9FfOf3h
kvP1QhLLk6xd2gqGP8tVZXx3KOwpf5TCRtm+8CApYzsuqcc2mtZZaVIEdNrycS5Y
EtpvgQkAHqwRQwJBjOnBvyeMmk9VYzT+g2piLFyINThzWe3c6ZJQ3fQRU7T2PgCv
r+7/teznshym2pEzSVMH68X9Tl0psW6B69QCk+PEOqSXwLrAxyziV9tJXMJHTKAi
5eEuFOnJlJKUAGlLBUAzgBtvRkgMCbwXR/PgWvFyukGmNOgPRFK+VI9pQVUCFuXk
QuWUNuutU8JtLfqQ+Cp3SDqkYhIgPBNtLh2WDvQtp5d/BBljIXeIp4I6IATlhgLA
7gRbrOEV3egUjik0WHceEAlCNz5a0PRQGReugfgQO0Va6/2mk5gf/ga5rJZvYLvD
+sSsNS+vhxtpuCTBzsWjPx7D9RpAGApE0c/sI1xR/8/bXCHTDYI+GvgsEgyYSVu8
uvIwGV2bao4yay2C1OwOFK+PoCv1kEiWB/EmVs8OfE5FuCPYbS4vLArR3cCrHX2q
Umvvti8eLMdI22Vdtz0aH/8gmx24LHXU2AUufdHFTMl1OU1eBu9JBimumhyog6fd
R5DDIawQdCaFvs9iPLCEnKBfRshbx9GwODoq0Py9F5oC7KAUgLs4z2R8ZcPtXZQn
XAOnuoPHU9HzAvEN8PVjmTv0dN7q8KvupKThqJZMMZcS5CPfMZ1gIOFBzNMf2nD+
NpQB5Voq1Q+pm8m2dygCx1rvjxjKD6mJ9Ld+guVRYm9O3hzVxk/M27vLtYGDT10s
Zd1vkMqJGjjglZh63QXoDGwb9n+T+SgM2X8z3//iscXbyWU+BVLtx0iiS2rr0NtX
7j4r3pSldbcWzjXoF2YG3YivrZSddGJMwQ3aR8tC8+dc2MVP6Y15R992eoKnid4c
tho3Q+BvkaiRQX8oSAJkDzHbpHJlwkre7AlZkc+OSChuV6Uul9G81qozd8bPY1nS
XwYzX2TYyAcHzdXy7Yzu8YPEKPsKlYMF1ZwaGJenm5SbyerAc9WbaY9ccib5A1Wv
MCGeDVyrDrRMfbSGfsyOoi+Q9X2AiluIQoZ8jbtKrekyChg5JP96s+rWDu+X5vko
N6A395JdADPL7smLR8GuJHqS5UWe8k/3xnr7IU7YGrrPU62Gu4KUn6tfRFACw4is
QGIpAm22XPngu2deMf0jm6kmdE7XHAnCR3ffE7KdQ6XKbh69aKasTkOY+VDjpBX7
BKRgyWffnNTzx6ZHQKY2jk2OfBE8BBZadSIpTzChxl7DGe04bwtNTZ1GP1aIXmGu
0JBGLPCgZHfBOeVEkgT51FZbldlsmghyWRFgdafH+yYs//8XJd1zqcdW84du5HNp
PBYBFxWxTADM73xIRAN//wLXuclTttlMFIlg7lORzOtM9O87KDa4xsr1HlMP5GEN
4FTTVmiE0/9WtzPMBVjSZmc4L7kxEhafQGvZw9t17QSfnE2Ev3bDODeXxnXpsaWh
FfEeRwbngtz5sTj5Q3jxZWiWr5EwIdRSDMMn4JvlOH7MvebyFNzQyZBS8LdBaUY5
E/PMrUtJBy2yZWLsokxYto6vL+6DO+uCCXIiZqDot4vO0Io+pD+7okseCW6zTEER
UdHcIIfEeY+LJ4cJTpKl5fONnuB3afAGZF8z7wtGLSv/dnDLIP4/x0IV9rPN1BzW
6br3XwAIXeBqTOgJqk0TTLUot5KmoGR9M+/mq1F7jTD93domIrhGgKiRIqaK8w1Y
zYM/2udWc+X2Ofle7iFvj6qpeINewHEndWRGokjUKV9AsyQM3zqxHmKMaYFNjhAf
HLN2NgQ8cYUOQMUAg9hngCVSdG0JPWPv1CR0umJc+NxYIy3xNiH75d7WxWZnKG/H
eC7lvDz+kEf6O9k12i/JU+C3g9hPy4KLk3zpOY/TOv6H4+4uGRNNqF/afuUX3qh2
D4I1dQiW+hn19kTUZup+GPFRkJSJANuwOPVc5eK9E9qly1TWiGQCenEjO7C58plm
edouAhZF/7mZIref3IjKXzR/aROQ9eT7uydedbsWy8WyJCB5N4X1NBDDAsvnFbfX
JGeApq0RRWF054dpHu5buqYrNEYUahifQEa0OJWHOYhRwesL6wrnaF509Wpvw2AQ
3kiYlJE7822vG/xDklEkB/TUP9VnesoviMAgy80yuwyvC92SQsnWlKjWFvFuiCnW
U9G78yAL1TdpVV+zgv5KTFMmU0I3z9CjzqQxDjazTtqlEtp9dB4rSDThzBNZkYHo
qvld4Z7abIzNy8BBNKRoSuTlRBKo3M7hrlB6vpctD6JOMUFoiAzPRMK9Fux23YWc
7xgU84l4ndEJn5qgO/DcRGlz5Zuki9aUPGNTfnEiUOnTuMj52OSzHcCk/xfLKdiB
mAa+pUYiMdNKbkSSjqo14rNftbb61WWCBmK+FFlaMMzv2UtyT35+j5fB/aZ5R0jo
Ywf17qwBRcxNbH7iNRQ4F5iSRciqD49+txTL92b/nyOv8sh6PaQE4W8fCTqc3cUo
hmwA7ornblTEJ2ZxTj3qnQ6lFo/JCLniS+YKboaTHnXAE5CKOzdt0M5wlH34f1Xg
sRV3OOC/UeQYjdIHoah4jkoFB1lw/lq5VxjYveRSkJnBjUNokue01uwKR2yqdOBS
yaqjvJa7ePk1/9hGyqIAqY3wIA+eUDqc1mNzo785ZywLhUPdQoRek3uQM23by4W3
mTv/A+iIZxGO/ufG+GgRnKA7Y7y9Jp5p5knoVOz9mz4hUXKUtjWEZsSSlUu37Vjb
ibx1CIiRzo7RJajR3jXwlf+haRTJgx0FGXsN0LdFh8SSPZAnnH0Ue2MnjS2axNmE
i6gBKWnSSoLm0SeXmkG3AjvkfNssY7bk6mA0IuS9xt9jRSzxVLepRy+ZRadHB2Q4
fLlJaqKUMiqBvF8pOqVV0nJvBF4m8LZSrYoBJLOtWBxJCoPRHYmwxMt8LKYuMo9S
GKh3NMHdcUJ6yqCSaGXbA9dmw5JOBbRdax0A1Z9iL+Z8v8L5GIchT4tIdi0niosL
dy1Xj8g0kt9OmZUntjJ5/kioQxZIkvW8pWgjUrM2avbyM0KdrvEdCtHeALNJ4eNl
bCEQkfALQg0x4tFBMDb4fhlQrvNuQSoJWZ6iBnsGgIV9mHF0Sozu9rSg3Rts/MQo
lnlX5djpT6lgND+MTQ7jeD+63S8bktTAacuCPukvwKxmeyGOd0QsriZMm190/UFF
P0Wg3TGR3egVL3RPMr9EP0GBDy6iaGBZiPPZEHo7eXYR7+17UzGm2RhDINK164Jj
OtpcgHb3jqfWv5TnaZw4lXCICMDwq94P6RDf+0jqGneFvL0NlnRPPeyTim2uCTIA
zZYebux9vgDe5ts6j+21GbbQ1OJPnPAjNPsVqWLHiTJrq/ZJ7UtiFcT+ATaB46Mz
OfREVH970o13AOz/R/ESxaeqjfV11nXbncwxh2L+Yj3ANPk/utC5M/PbuQ8xYWlg
3n0d1W58MAMSLnOU6v29u/UDk0EeV4udSEQYVn2EBJ8uXzuggz1Bx8Qn3d2x6pIi
O7ai2C0h4Vjb3AZ5+lQIRVssW6N1F+kxNgBOkkgDqG+hQLlTgpssZ6LzfSv9F28w
zvEc2xK0LnfDfedOWpr0ZScggGJE1goXmVuB3dWgXbDugnPyZVkkq2H0fZZPUP8k
Bu+xIW2bXw8sILzPhxCCZnxltseR9QA/E8/RPb2JOetV9aSoLFTFv/gfJ9k7USJ/
iV12xBcgJ8KTPpoOBcGaJ8+RmHhLnrvjrOzebkSYSGzwtPf3wogDfYt93NpdhqxX
EbEXUkKyVn4v3J/Ge2NXJS9m41PRds4MvU/LMlLp/Q/ivQ+UtcHVgpqDt7L4z1SW
uKzrrfdGgawSzNSck6CZYaZfKReCE5U4tK1LfoPBeARJST7Txf7Li5dKb5k3iUf5
ypTrpCiB6umZYM6mt8GMRA7UX0yI/o/1o78HF59jpyjOGo6nWX5uwEG6y299AOLt
+MZiifUmEr+LPAXnFkHlcGNt+xISb+38QoKcZT+RKwXzcgRGa9vQD2u28196Zegl
8wiDy8YBB7AvEXLm5p5soFz1yy9Nl3zCKMIPgoN0vCczp4YDA+/RJBUC8AK2G1SJ
ze7ErQWe1Ds7xm/C4tI5bRbPq1eM/K/FXbpJi0GJrc3W8imuHaWV2QejwRN00ntE
HhOJRjrrbgwxygIUuQsdz3NzS1qQRiCLKGNlbCECL2Nvn42SI2f58zKFEXOsjsRb
cuMKHA0Iz4kUh1pEFRzQFjVZRMO5/Ipr6J9ogmUmbSBqXEaNedIb5TPKss4+LeCK
Ezjv7DFOW1E5uAtxogaiXrDP943M+g48OBSLerzmg+1rBGGRf8h33W4e3hDSmODg
nzYIvtorTShaLrOgryUieky9IVCTErjApxaneZGx2QdgQJQFkdLnz33g+LhM8mGe
cxFCRsZaxZG3GZKntgybCzJP9/JdYEAl1WoyL+1kumxhIByS9wq+B17h5d11C+Ml
92PGHoPZbNz9CYlKLyNEWChno4ofZ8njIkD3m1EhIl3qObUiTtIuTVz/yOuZs/nc
ZYiDpbbxipWiERTODgux8fKirwjS56uqOE+Wtha76QOT/LBfJLMHZ1wWaYl7nXZi
vPErUuj2ic8RJx2t1EL3OA8iwCiLnTtWzcUFxatqQI5APkoBJD+PCtB2ylx8tDHG
JLg7eyIYgSJDOugUp9FS81V3defK91yYZlSLFHl3aE0LIivYLt9vywr/k+ZKedCA
82kR4RUO0iBtgouP9snzikXN2gM61FQlkmbh4V4JalxdIla/uyDJvQtfxcALlaXa
1kVLjXvNoRh/OJzlCXSaa6X1xPMQH5nVQxPj5qDVNPCpGL1r6myKMzmOEBS7tu5V
XSw4Agc/CMUDI7cjRzBCfDX+gHb3KGG4Otw60VKwY4RkWDFH6Utw5ubnGtygj5VW
POyZQykcBTA8RoTqmeArBiylkSSlDwl5CEp33R2vg5/EwhEKTnZBuR8csdUow0Q0
MevevFBr/YNzBzOtxa8jLRIHhQnLuXZmjoZyJypBYysp8jTZxusb39MM5jtGFRti
wuCfpWB3rT6xD8LYlNKLmG1eZD0JqquEzDLmMvp/bU6E30c1ODwZqFGcKDdASCX2
xSgKF9SOtFIn0Edvz2XJ2a52W7Q1qkr8gF0lK7nWYHZR94snTI5fzXApUDi5/9J0
5srLieo88EISxbpzFkSL2EihDmBXH6RlPywoMODrj5hEEAa66OMvV0mHAFFSFHki
afm4YlsNIDyRuMXI9mUCasC2xui+d3yI/Xou9k650WWYilq/+9zZD/ignK0rzXlX
Th3ocuDhDOHJUgIyfizYbGX5Y0CkELvpWJUuS9q5VHbk+2YNYMqszXtwVAxVF/Z4
RXO/SCTiZFYv1gWwFLgyd4xMLDHxT1M7OFF2mKh7qZbQZTThRgqb1LMH1flDYgU5
RNJ1EJKR7KohJCWz5ibzBJ08utBI3F7ckCDZdTtR0unW6gq0abGP1WS6IhilY+eo
KvDeCEZMBGk1DDTNnvyK2Gu1P3vJ9fbCFwZawEiGq2ljfzPpQ6yEf4WAtGvgJwiG
Ifg68fpiAej2NExnkPbYmG5udsVNvndbQ/cSBK2q+oOgUhPGx2kR3rUAx2cx42Ex
Z+etkYfq9EFHNO8xg87kDkEMvZK3cQsvGD4T83BEtE0Q3ZNnonGRukPpDVa7AdSq
JKG7Ze8VoE7BxrJW4M9GLZ2qEHZMN+S/NWxNf1j5BsNEo0FOweYRT1VD3lDEvJXd
WIeO9Sq1o9xTefA6RqMwhABf0rID2xmMUnvEiWvA41Xna+sqmJBCou9dnrurQiIz
4KmgzjtFkkQvgZ9FAJ58AWwlJsonEzPhfLOmmZC5reu1Fx1Is/N8nTK4qFoMQP+I
Rly4YEFVOdSAu1P+r1rrksVN5AbfUvrknCNwb2j+ijg=
`protect END_PROTECTED
