`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
spTTWirNXq6TtLzDCKL/M14dDXrEt7NDkdX9U+Ym1el22BYZ7V6z+CMXmvg8qurk
qPH0rCKb0Gbpt8FNE6dMrMGyNgPt42Q30+/3WWSXCHfEnL0hR5vivUaxIg0zEU/s
f8LFNPe2e6KQe5NQRi6197EYcOk1dLJeETPgoQU91Z0YG/PjSrvnsO5l0K6aMN0y
nP0P+qAhyOOuMWGNPfvIQn5TUxiFE14gxTRpvYVaYLzDHha84/m23oZMZ7odyj8v
Bqo7IZxopJNotZzGceoL2YR33abB8wXiz5tmQ4fxibROAOJBudgG3c4EF+YtjDMs
aslrdYejAYwxgjJHTRFMdmAzDavPy4KVa9uVJi2+5puM1Qxbzo9oR3X6XbaMIExE
Oeywb/2F/tKsM8wa0rcL53XUxC0GB0KCNTCNExGPygR7+ui4Q+jfy35uLcW2DG78
7bjblUekZlpfaJMwpyafIRlrktd/1CJUt4SjC7h1Axq+TtgxbRi9oo3VGPEq1SuY
8lrixNp+k4vvlASCcwz4FFnWD/7CGdTHyUMWDA8+rU6lnrsAnGFv0+U0ralo8tsF
dN2H1na+nI4VGlPjO9DhsA==
`protect END_PROTECTED
