`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
noXmcDIv9l6eQRwUXHr7uq7ucP/D+lmILQZvDusU5tz29aS3ZewmprWIoTzglNvz
eCB14R5BEnZvax/WkpBqnD7NyVn0iICYDA82DrzorcuUf3uyt9yUy1kleo+/6sGV
5BBwRdyhipvFmgOctLQ538sG9Pit6Dhjc369NfDsjuml7Am51stuXx7iPEelfwAd
GTdFmMjhEOedBYRPYBGwstyaH7NFErJwqFMm7yoWg98qMnos9PP1k+SLPCwvfSYd
wr2E3VV1Cx5jNRamSzLpus10Rhw5HCaz/MaT0PXwXP0LW1LYrD7DmYpvAvm1a/oO
D51FlXoC7HNu7BGQt3zfrtMtMf10q6NhaicXLg9wmqhu8wgR7JMzwwZv2L7/kRCe
a2x2jYJFrd6C5DHcZKizQfKgi4vhFrCdr7J0MfL2SX67nOS/S/eoKABCsJUz0Jff
RkfqYhKFN7MfHRnPbVbwOolbpR5n3OCbhVo57kCXw9ej3n3yvjQH9vz+ZegcxXDf
ui5nGm7h8uDdCA7FM5Hq3fBEKWmtFpffdcyZk+lTYFf8uWzyfGYd2fs/UjsZVFwi
R5vR2t0ZZVcd67jZMif5DxVdfykQMVLdbvJWVDVjzJ3fKRLTa9krvjoWRyrwIm00
m1yK4xAP1cPqzHJOMrmLifmLEzkupZjxmNF5shPdb0XCJEYWsAo6iFeQKpSFRWcd
er4i4KsLhlst443BjJaoQ0BE+968PWMWTb+3HrhmDip8puIIAKagUztIct5eIWgh
KlBsz54h9lj3pfjRSKNxLS3dcpCDvW9P4myWo/XgkyGK2PJGHOIWZ3AdLX30iL0x
hhpoVcPb34SNI7AYsf3LW7sWkUC/P2RJxC9Fo1385MyZv9sTRO2GtqKRigVp9OPL
bfhqyy+UwY10TPhe49Vb/obbodNVOrvqojtQPVM3yY2R79e3WQwaCxJDKXTwL4Yg
nLkwSRlJSoGS9uPaCKRgs7LagB7A3ty2sqwrReduMub9esxUhxr+MXQPOUDnt1zA
pGmO4HdcMtkOAdiY4BBlsyqvpx40zlSG/YFTe1Rj4+nHigNCRPYc0X8pOQwFWNZL
3jAHdj3PpGKNVYgzYK6lmhdHJ7KyTyvYmHNb5huy1iFB1Nhe5+k/BESO6sGu3rhm
+x8YaW9Wm+n2JQXhD8CFPwfNHRT03CPzIihidhk1pXQS/hFJxBHmMCawGL/NGNKn
egoSyR7mNkWwlkk7fzaPx7nPPcwmJpDIYbNu+h15c2ZLO+BI3Ye+5goL2ktIkxUY
YF2uWztiXYBHsj3svdQxNW0Aj9v9B3OLrNLZi0erNaNpy2Waadlfuy7GKa3i8MeJ
US76R9E8x05Wa5/zLLjTekwljOWCCxWIcT4/AT3t4411LZyE065h5WRFb4ZDmaXs
3QFjjvziWxLQDFrAE5TmHhOcJzOHkU7C137y9Alt0JX+iyQQ03Q6PlpvqhLkb8mE
iiOlQctj/+MEkSYKcfrpiktVHQ+FxwJoIqIlc5oKTWDX/QguT4ArQY1M/kD/ERNf
GNPZQNczb72Nz398nw7DSvMJ6OJZgQejXNL6SthpC6vxZUynxk+paXx7FDYrRCnS
CCHhHvaPIVeoZDOhUKXqAB9zzgJU1sU7GDlZLzEH5JT4q14LdzvT+5SjWrp5JfGn
pO8maPFQmVjwfZp6FxLzCl9tcSLMatXJJ/vnTM/E8mB8cLI2nhVCx3y0wBAnhcUj
6cHyFxS/wLaGCQXs6HbvGm/yuXLP6cFgMTyO7sNFs6HTZ1JnBFMtWQ5noWfg2+UP
qZ4X/myvMfanFAyjux5AQ6nFosdDRjd0Wu2jlvmm2uU/1wlPmYjGvkiAvkpDsEqT
bhxPFvGgxku8YzV0z2CIuNZ86hBdLFJKW57WS9Ne+5nl6y+OjKmlCqcI3WGwHHYf
7tixGSj9fT9uAznHryfx1cKxkg9KJZQ+cOfCObCIgYbsRrZNYfuFPwS+WrYd/XLB
ZWlzQh1qn3xakwoV/AWD3aJe1kd+dPQg1QraThdCEDRCDeZyX3JFM3z9JD/ViAdf
Czr/wv8foBijmnW2C9piOdd0Fka7AL0cCH05kKxc3MZ2GkuYdkwheVfj4158ecPe
YX7izOzppqrt0PvUug7uA4CTG6MZTZlGEipxg9s8D/uP+ykqEiN1ZYIl40qRStEj
t086WBsRieHFDodoEim/x0wrvLUXsLWhDHR9nCa9dnD2jchvJyAkZa2Bcxap1Hma
jnEyTURNP2dtuOIO4ZrLKB8gFNPaKCz45dyqVXJNAdEAi+yDEsxU3Tohp4fcnPyM
J4kZ5rp0BhVTKLok3jnhNetE/YYVUzZ5IIrAuQFC3rCLkaVyqioMTo5VDAF2/KTd
DzyhFhvHrwxXuPQVVo+I58+ZRAjURI8lfTd9/mVXgTWChknOaLsn72p/vj+9gmCs
qTGSoeRqKuTCCXxwSHI3xAzSgq772Hg4hHad+LxIcWaLMty4MuOf1kJubHtE22b5
zXXzv16ygHbVNPBb78ckX9z26rnTFnEBr4teUNrzggxPwr3SuFdXakt50qRMoi6Z
6NaHHp7pCI5xhllrMnsnhpHB7huM2jvdh6iBcv7c8BoUtdUatQgZoY/fE1wNgLWg
ZGBPKGsZnOR/Cl9cr9sWAnBiJjB7RPAn8IsA2OzjFMvc2U/+PKKHui/iltL9Sp8i
5WdWh7tG/GMOr5QIvIBMvzaMmMGDoJ1gt5eEghfsbdMeqKNKZXCCjMwlh8HkEljs
nEnRYYcd9dDFYD+aJDHpkYhPpBJhCYNRTFcTZIiIXhS4PblfEhk1EjT2nCFQVAxK
vCgfj4QJkFuRSjTnwHhpqsPDdQLBbX1zcSg+NvB1Mc+jnjSk4Svt1KIhaurVp/LL
RydmL3forjd5UPx0VIvwPUcTXf1MKUDlP9a41OvVVTds1NH3zi4YQryBtJRw5yYR
r0mCt24ih2ZmpHVTEH/yN1TLiGL5s9Mux09QqAwgQOrBVe0RV6/QK390VNTpn3j6
YZb+Hpxp3H85rledBRr1hj26l38WnkXkWI3svMRPHVBseun6Cnzt/ACz4CbDhUmD
dLj9O3dH2qb4HmJimO9Px/2Iadkrt9jbconVDFa7MOGAO6C5qcQoESxRY2LtK9pP
uk1m7GUr+Z9pTQqaiNxKSkwCogZgxqvfm+drPOiINyS4J1IYGrmaBfPB3lkv/54p
j9qm0YmhF9DQ4JD2JfXDLB9IPwB50KVE/XH+OG2LmzOLII2Lybxugh5HilfMou+3
g/ToxFmj8JgHyt4wHE24s4GDmGSA+yyWyRSIMXq8W5Zy/pKjtxrb83laOBOTxex5
LvRnQHiyNpOiEcBbfwwpTHl+VdwCThpoeh1H4wEe0CpyREoUEMmWHgb+3LeLytRc
nlp5PAgrPiGwbz/jh0056NWwaVHwjGE3pRhuFgqFM8gCxiCp3IqZYzYYlrOnUOvI
Yl//4f5hA4saxNdbYwyybZWy4RAFstHLR8gcyO+4uJw3hY6i7EbyQMgmDP6dsThQ
c+roUE9Cp+/CRjnEM6bM9bcThhEy05k4OBEe2NDSg+jkPh2ZuSL+5Hsh/JnA1mfC
t5PM4O8fg3+LZvLCAXJj2AZUg1zu9DEa0kEnIqJ9uxmSbfsrGVh9HImXKclqyXMV
2kAAIeS2GIPIUjhyA871kjlPBTvb4q5SaKqyN+e3o6ezjY62NZifx4k8z9B3NOZ+
PAJqGXT7Nxr9wVxroPrpfjSWxfMaw6j6pFfjRhc83tctE7UkS9KuBx8k09IPzKSv
2Jy+xPDVqTT5CmV4rYRQoF4u7qEmpReoCAF5HXrrZp4WL9yizqIj65FxVUqtQO+h
EyqfUcSe3i5sqVNBcNg7Ypg1SB0xHIV+4dqp5E73rTRQjF2UJqIu5teO8lXk8ntw
aE6qQfauT17Fu222RFmVi9x2Tzl+AH0fvaPlzaQHEkUxhiH9RzX6CwA++lHPs9hE
fCQzLluNUrHh8Fh4weff904qmM5sYhRyfJb8SveqXajhhvktWy6Zh/+Ub4U+p3o1
KHvkSVQXraANhC6jRLD8/pxdlZZSBMOiPU38PEbWLpyaabvAAmMICkfQZcI6n+nR
HL9kPrVjR+m5YJ0Vzqug4CvRBxYZvZtIHVBnA4kKFmatWLxUWN1x9LrZx1z/E+Et
w3vs4IQ2aKehaxsDjRN8Y1WV6euie1eOKcAA3r1nHZwwlNeThVhAHXFuRxMEp6J8
wEHXVMYEOhNK4JhU8QCM5oGnBfN+dZDfQo8DS+jOh/d5NWQ/VPloStumlFeEtzDP
bbMVzeIGl3O8PrWkKdOqwM7et5qUTQCE7u0cbyCQI9Nwxq9c1mNwgT4v91MXJYdF
ZmUDsRtwa3Oc5apwpKoPmGHYZn5LlpvzNszV29aXREiz6GN6J7/nAUq/nJ3HBCWS
bgVkWNqOhStX45l58xK4b/efqcKHgAtjZSl9IYqwfBmKB2KDE2yfHEVgwdOkPgrx
6zIH6nWkZ/KQ+5NaEyqBnUArYT1W8co2Im2Lu1WlnfgG1i8g8FlHtr2kRR/z2eMz
cs/ORUKUhHgvUtwW22QboJOh5gKfCxO74kwNOgyzQKoMtYPV0EuGy1NJ1xqBDTUI
WgmugNyfvS/8N6K3KZ466HUmVH0I2kI29wocwCEE7Mpfx88rrrOymGROORFQp5Az
sA/ZQGLFqrooMwWJCnOvZfgUTFMTuVD8FFD1Oo7nTJtZ1AISBEYhCNOmrfanEl9k
SKmhbBbEilsqTsBGVSyGlj6VRTgdm71S3wb/227vUHEoBR9wJBppRSZUZ0WwXxFD
wOBHlTCiQZQVBCMD7oG2FYa7NokGyDD0gdVExcoaR7UcztfL03j8AV8O+0v96PLl
z+34NMT0dv/OjcJSO1H03OaTI8ha0Qkp4GwH7R5/47zmNiw4OzrP6xyXUl4JAx2o
nzfdoeGn3vQNb0ilUrASyfwdGtbTDe2h8zVABJ3biAvbf+if+0ahTT+axHJeuV4Q
dSJVuDLpyFSsjc2jb20b0N4noaaYF9Sq6rRu0+uNpKYxjtyow8ZIAoWr9Y7+USxR
X9NYAfE7MbubGw+MxZ+EFREPXyTVkDymBdByUiJiLEsKYNdR5f8LcYDTRbMGgRta
mq2z+9NT4w8d+D9+qGTmhsY9bj2SAFKoQ6fe0oAw5FA6FUFGAPgKAEoPcjnPH3u/
Im/dO9ybrKu/suLZfiYg3VWy0Y52oHlp3KklYxOEkTkafXpkpkTmv1oaQcI6C/Ng
Qo7AvJ4V1VQhCCkuVd0eiKER11C70TWN0Ip9w933C/D4LZBPtDsrZW7uSQeVe0gz
hpB45Xk7no4r8TMdSrppzbLHwVPeNxERYEiSzMfszEUoW0VptxbjTTs8QhN4hedc
Cqr88fzBFVt+aJCvZ2E38NAcsrzXJ1kW8Im/r2ia6vpsKq84OykcmAKp3vWDKJyz
5u2en16SrDTRsJwPxtadlVcD/ITUcpnB4Blf04yPXAQasDNG40keMaLnWUDs/E5s
sr/2M24ESzmF/TJf49V/a3BYWn9DRsBlsV2MpyMbVbBpjFi6XKPjDHKr3z2n3A8m
lZJMPjHpFTIyu11JLG4ZlrEchIvyOCi89gVpMD/dUQHASfFs0f6BsRjRci9Z8aTS
gSTpVpqUwGFHNTGdXgn/dZvslvfaeJ5HcVcV5khS7+giP4dRYcLagROX2A5cGuvH
cGKg4EONk0PAf+jHXEHIge692jC7VaekAaCHTXrHrSSeKs1wIg1wHSeKOvy0GjQt
U3fN+4ekUma1mAFJh57BbXC0SvoSijf856zlflquSsB11+qOCYLbeBvMac14KYQH
KfnUzQqI3oS1xgIkJ7TjL1AjyX/9Ij7dVOBLDx7TXmyKVaSZufDGhFbQUCguxEgA
PdwoFFg3mGt9n44DIULW1H9wav8Pk21hsWqJAv1Vz4UOjddyS6xsLawXiRfbpvQZ
LZCS1F3UzyjXX7ABGeE2mOo9fd7erIqPWpwkxX7WiNNM/Q+5P9vmQS/ZSQCF5RLP
1XfPE9ULtEiYX6JEf3HYRvJXNngYNjeHXIsKPfD1r3Gz+kq5Ed0aPa5r/84l5fAW
5AR/3kxgrOwvpTrUu8FWJWc36gGO4/rJL42bO67/JXxyKQoyrdYWRStTj4+FkYG8
5WN3EfukaqubRhw4lTrSn4yk4rnaPJ/5CRZ37MzzG+fsOhcTiL8O7JCw5own+WXN
dxPtLADsnYczYImtPEptTG32WVAy6bDPSjP8WUpswTqzoJF/4M3hNI+ynyC1/HEB
5v6mTO/59lbatuW97qLgyBD9VgLm2Ww4V/XFlVEQ3ioOBQ8ALJpB0DM2RZqRFLTJ
t0CiqDAM3VAL9dKLMr7PPpmccfVV+ZXIkg84JEkrLHUSpw6IU9FtBzROMppdPS4P
BjCsOc6KPcgdP3xs3KH4NByQnI1ZD0sAMMIpOff4tTlBn/GqhskOnYDTZIBNfQu1
PT4NfIG7pQL1RvdWqxAKNAQkmuzgY6g5+e5tPly3gqmlX+zxZpWwgxx5XLLIOzvd
IfeesR1WzeBOU0ID8GQeYSfILb+7QWzh0mc1ZyzUzPL4lcaTjGlLrf09bhEr5xZg
X778ceLkoQcjrEVUODogRq5zwHQHvd+5DV5vI1vwDScTWUYjFUODZogzhTEtotzN
M/7F6wKfxm225emqJrkhQsiQsTlhvvBMcdQGlGZtLmNnm5SOTbJR4Z5jYGL4hhyG
+816lDYkahOFdv0gDItqMxU8vpl9bB/5bwAJQ26FSOnQvVyYT251NWVrO80xonPq
iqBdMJ4uVVBkrZVq69g7NX3SyAjgKc7h/h7snvWHznO2WQKRXkd5lloygku+fBQ0
f9ovp3jZNnPq8gJid1TeUuRoHUOP1+b83ei3uB/5wt+igWDCwgmSslIoJlFSG4+Q
QiQmeUAzQY//huAIhYMtsLyTx5Ot+FMHfHmYkdYKayNhc1jEWfaeACVZfBMRdKo3
ejcRIoqu6hu+ei2hTAtOvZSkyfojBhirMEASqaCo3AIRkHpn0SPWACTgljBl+29o
HtzOKDkvblfQ3wqsXfU4MSoYF3FYCXmMcgFYOH27gbgUkJriy2VK17ddyQDkCdI+
sBDR3MTnBn8/UfL5e79+u2CatwSL1gfQuhXFuvwvV4/u51+h6nufrjUCFfU3T6bN
4GPvxAht58HFrc+zBcecsgfzy5CxAZsFud7/u56sVNJCiWzeNUHz4qY9XfoVPS0G
HAMA7oGT3+G4AAgbpVYDqEvlup1SJlwxi3wrd+hOMYUVTYpCbMNM8lCz8ujt7wnG
8/elZ2YiRhjeWD2uNUqFMSsrGUrW2oohKLNiYdyqyemeoeKs19cqw+TrSJVecTXX
WXpsOrjNc1RqDhK3zo45N78Bmn/wQ6LJ9YA6QKfFGk59oKpYQP3v232r9+IO7f5j
OSYu7xfMPKahszyThvrCVkz6WFjk7hVdavG2OGgtD1GDIrfs3T2qWz5lud3A2M+C
I2S3VZbo5E2yyM56qHrL1UMYL/6qHgrKRmX0SeaOrGGsBFndcYs+1P+eYHYjyDBL
6/t+Zs9PohboIxHCov36xjGIBfBEccoRB3p4IIf7aKQEWxN4FfE2aeeVriCzpZXr
UjHebfDbl97LRUgZlXBZ/telOE7lsKnWz3B8a69xL1i07nzBAAYi09L632yVKDK4
cnFbKAgRVKrdWJoHneeM9BQR2e8HiRCuUcXr1laPQv/sfstCly+F0SFvlZ9R1qlg
IaZtDE1V8/IoSDIA5ZuWS4EHVkuB4394WoemjiioC7RAQ+oN5qELX2HFCg10Lr76
v+MxKAmmcDMicE7PSJF/B7o//FHf5ZfdOcVRdygnK5I0IR2ih/MQ1NGM7283BpmT
XHvWU1hC+im44fJHYIN8LLbJ3fkL3jTFL3LjTVnhLMm+7T5uDM7jbrgRyXfvIKEW
RpSlvNQY1qvoRkITHWPVbQEYH/F8y3xu08iyvRWfK8mHhNwfmWK2hLe0jQNaBRMQ
BUsd1wIiD2pe2eRGSVvteF2bUgJwRi8Cln8e4PcISWkY8NzDdx7QVD0Gq7Bdk72X
PO1TC4rnCBQSoaaGHvfQAnkZ/hWjz4zPTR/5KIEvkR+Ra2OTsJ4sJ9wWdicl7Xp8
b7GIueyrcmzEBCf4lvme1M5x8pFlftDzTIibVmedOiNrSE/lEA/KRXpa1s4DTfOf
bO0z4uao56T55dd68RabOhB11SGg8QCO5sq5GKicwBRciWglq4dhKnsuW8lMb+Kc
ea3psXFJHKAYoPiILBNGWkdzawG6v3Axv98FayoVy9mFG1U/k7QIWI/nU0vaaWDy
cBjJfDuUojX5guW4SZSwChjvCucOvLiclq1gsXmcXy2tfwycSxSbutEGNOOv4wX+
4IPEgUPpx7ywrR55BNbLc9opbs+j7DZg0MNBDaLslprEAa5OJijoeu4Uo6VDoq/o
EHypS8lHx5epLi2XsYToiQggWgF2+AsktX+Mrg1Ka8VHP4/VgJc8mKOTqvveY7Tv
HBaDMsOzqhD0RQEjJPxpbS8+98sxRJfR8GCSVLIq8pio8WNEJ3PG7fWu2/PxjIS1
OKvxmKUVBZIxePz2XpKHhe5a5+ouBbHIQV5df3qDdT6cHR1ZqGUpUfnGGxq8W0p2
mNBYeahrqdq4dS5pSpL92Jo8OgEfoe4Glsk0ySAcyjqbZYp/g3eDIAv0YIctQV6a
puaxMasfczyY8FfTQHBxZ76vgITKQAvuPZxlmqQL8DLlS/pByxOyd8T0FdT/Fagd
VwZnLTUxK0DZ9lp1929q/FcSPpo7F2mj2vtoW7CV5Pk6FWXhp6cJbxjXJCInKJg8
GU6PQGKWREONbzO7IfkCPFNUUer7yyH6eluYCjtP8dMxDup+tRTHC/i34tomNdG/
AhzL/XP6zwyzUcqFGMgbOd6yj3zRV35uKm2BOptTQr9dLHa94XoKzM2Iy5r9JNGN
t53tQ8PmNwR4zqrXMzoN7mcwq914zPyjn2C+LMMv6Hno4MkjG/dJT1yyyx7RqTfU
2ohnm3cj7faBfCahbbAXAsAcWEJZMyJwUQTA/R3TUMOFzf3etn3GjACyezxhcUGQ
e42wGCBsCwStZuos0Z+SHD+YqdmTMH1+o8EBUVcETZlPKseqp+QrBqJsFWTEF4xs
gUZsFNRXL6iaYJdIfp8zqx7WSkgpTCyTyeqNYtuaBLV/uXMLnjS/JL8i+oY0HZux
LrK5zkMNAu+p9eo/NATgVw3GHTMW3v7Lktaq5SsIxcAYVbrwGlQ2dJA6kxLaz3h6
j9YBHl2UrvU+ZTA0QSoWIyRnra18G/YNwkZ6bh41FYPKtHEy2zx/yaRRRBckdl+z
NaTMx3uaouNzfziN72WGdDEQZnLFlyzB7xT4uxuq0lxYs3mhPXCHu0cT7HRk4rzj
yISysmpJ7Qwq3L11D9GIydKveFOZSeDJg/K12hA/5APYrDxUdQN9arhiPX2yO6mu
5RNPbXc3IDVPI/VNrSlMKE2y9ucDkt54W7xaanqhwSqgLXsYK2cQ1JYvi8C2uOk7
bvvsNLku7TDo4CcljbmSKawGy6Sl84kzsdnC7now6dKGffSyhT2X0aR6+ceDUQmR
mlJm8VavOQJcOhGDoIpwKOfpqN2mt9hgJoZiDgNyUyS56DbjboNeF5rIb513WVp9
DY1gnfQ/ouTZ8h4YPe9Mns6Vl8XjKQ0Z8mpvDLQJKZcUDDOrQgrNHcJ4msorKsF9
PuspRWQMe79qbNjFXkD9HZZJUQ1Il2GApu8pHQ8cAAQn0UWcNZqgvyJgh69WjL75
viLzQWMmaKNyTnSvL+/UMfxWYXx5qaGzDROJAvk3rounwQz7hX565DqD2GsW9iSq
pf3QAT2Otp0ysRKs8xh2Zmrg/e5HOV1tiUMr/ItjEikmouFIrRKeyzYJEEVAzon9
NxisDmJW4FAryDV/ZPfAe1slLkG3epCfJwDqlmg7tbh2vlZPggFitVlEj84787HS
RWuTnHEpkmq8eGri39m+i7vXvShmuQ2MN2uy3XuZ5TcNGFN8iXKEpW04bkBr9/zZ
1je/5MaNjCHuL4U6jF13qYIQdnjKM9iuXPHynFb2swuCjXVuSxRdWROkx/sE/wrI
tdimXXsasRcv5SlBDXWsnKPvPf8900gamK4ZuU6uzU7DPG/5vMl8A+4ikSGhuzw7
uk8WnFPoyA2wh/wBWAQes/Q8wFu9HQM9P4WGsNKmPB+Hi6h6SNMdf4bhy0nX/oi5
rabQU3AJxjDdTJqXz4oUSx1LAq4m2OWJb5E0dtFi6rsXj6TFdAMVaH1ZiqOVOW3B
DzDPuumOtwQ29tdveTOwp+GaVFVJp996vsQK/3qsL3O3rWh+2+oTyTNrZTAb3fEs
f0bVnascQ2q0crHCUf1KBtT9YPxdUOTXR2b88CFz+lkZOq6MFogCgWRU+AcfvwlV
2wjnRdatVBOhJ7VskHAlK5ezdukOPUM1z8fTBj/PaWjRbRbVsYmNTeXhTZQXc0L8
vp/Xct0m43JXSF0sPEDyuGOhjOFAmgX7maTCAbb6xxUp0iqH65yOMukyJ3UG6e41
HSa2dyUmGGo0iOqNtPYHA1fPXCKUyE1AJ7g7h92DzGP6zu+DT8w1KZyEkyVDsj7Z
RbKwlcxf26y1upQvwR9qaYfhpXAgFgV0A/gtVv18IDHwkxr2DIkh4OoJPrxaH0By
yKeY265QAxztH9/Lj8z1wqGWaAyOCy427jukNITUKFnhcdZ0Cs911Gz9s0VXMTgA
sqRGzEdUfKVPW6YJs7bwwsxpMMAN0GzDX5ruCcgQBeugzv4hwOv1KCtCM1zgcACN
Y3bxDkZLvTO2a5W9EFR7w0nQdYLQldcJ7mvKOIHuF/v49lxVNCeeL6P4t2frMOiM
831lg7xdAYkBQN6kfsf92M/OeFjRoE3qX5NCc/AfkImUuBQ0+X+EUAExikk2hg5W
F8KeEPbsgiKoQ1pUAsinFiZxcd/c5/0uAVEgg9ynagF9AeEmnFD3lIIsXMEBAGiU
wUzfHOttwlx2+pibSFh2pIJiYYNZLwW534MvbWHN379Eu9DZOaNf5ghr3tDh51L5
ptBQy6F8tj1+mULrRQh8ksJ9zEOQ/omTfJJrCFAydoPQfoe9IWqiKJlO7AJ8sjv2
Olyxsr+oGi6s5Qw3jpG05fxIryUaadZHgPZKCyGAHeo46Cog1P0p/Aly/HOaj46G
pNJ35lRpST2YH0Wh98cPvAwNKLCjxabvd3cFxcN8EldK0amIO1AFij4an4yk2KPD
eVwtP2M0f86szgO7OvIz/tdZGm/rWM22rgT9L9eix3NSlnGGdQ/huJ/TLLApn7me
ZWkkwa9utfo/1aa+zGgJ1e6jfVCdR31WJaTJZP65dLFvQu/laxyguSW8+zsGvnR/
JnVoB6BMvUWwfiibyrDTGimhftQYQIv6W8ovAyTWdR5/8cIeTZyCJmEJiwsxpii9
95iAGUhHVhaInp94HO77wTh1DzVmA26oLeiZHIBs2KPlh8poKg0pqtw88q85dHEm
Gev7bIpKuqwnPhSr5PB3JBSc/alhxWgrtvCRtPwdpVNWFy9O2I+SbLxe1QQydNvb
/6lulnDCECi/tX4uEHF3Bk77tRU1b3tirF/Ix+oumU/0OZN/AuNogd8nm+0Qymdw
+g8n7efiNrQ54M4HsjpilDCtXX1pu0l+7aCHNd3l27hCK53fQsofpCtYKsZGEe5o
HhpELFl63LLeSyYLG0VybPDcZjPlU9T5ToEIYEuB0fcGzTYy/QZGAlFDb936o7BY
cjcPepTdGhR46NkQu1xJkdrJfd1LCJgPg6CVW57ixrVqZXzWBzXHkRcjWhJbp2JJ
nPR7nKln7NQT//nU6caSv/ooI98OW5xlWN6whty2sI/mn2EhBXced6h1DbZxzTWb
2AIElrgFJyyvJYatSh7O7zyrfX65TwRIdDPRvdNdGOXRKkepWg26wBOlHllwv9CI
kaPVi2dfAjt8TZYEsSKuZSjKHxNVKi/Zd6WWnOh3GjHTCGKbQqQduHqzs8OoLv7B
fUGwoXcLIao4d03e7h4VAlpSfSFSh3gwltX0ZOgC0xpY0+YHdfPLqdoEstl2QA2O
w+6kEgWJmB3Dcy7VbYL3p/gaCp0aHFRgAz2PhkxEuRt68ZPVT9q4oql50u4RAAPK
Jg3gMggq6AR52SIHHxLmctKZ3zBeel5W8bObtCJRxiSYuDvSR+lrjlJVacrE9K8/
6SBJklhqpQb0fA6j3QvfTIOYsusOmLg0IPMHAWsi7Nj2DEQsXkiJxB8Qd82HnG0I
pb63wxV44zVAIw5kAOELa4o940xlGNT1T+f/JQJ54EokMH8aKhWhvhfNJdhgrDAK
KSzACMZ2y6lHxB4mFbRyIsAnMxS/X4GN6C8kQmutP5ykj8tsyHdvsfeStMYMHjY1
3zYTKkvBFs4/hSIUJvWnOP7C/WV7Orsua3wb/+XjezMTMwZjzS7ZUDkbcKwTrhy7
1b9tpbfWQy4uQfFcrJdzeqxTdjT+3QyYdvyMgntaaA3cxMs943nl+VaKniHLViIf
JQ92zfyS7b8Up6fRisIGLf0eQChguXLzU+uGk0Qqv8Hm478d7cT6872J9Bqn4Zi0
6OMPNSo8sKmAYUCWN+HpN/YJbaZ5C0zBwcso+zh8DLS58iOm+czcWevoIP2/kr18
g4Dh6aOjoLHyFh49Wj5h8YFNm+yjC3FSQDX58z8aqxq4Njbuc0mnQtLkjHSZCOuL
JXI+f5QRr2TNgMEM9TV0TpLMFx8T9wLPzVH5O15q5OFsOuqt+fL5NvdZrUgGrysn
yhNKDiW2aeeDUXzowIHrQT0JZc1lq7aiAh7N6jyPChB70uDT5fwhYEuvbvnrFNIf
MB+R9PU3/K9tySWlRV+LKxpEshj4bK+c7h+6oqgTrX1gKwtzvgjIMlWsKWX5urRH
kKlmrGX0WNyHPyIPiZYzUOWns4ZZA+TkUZvCs/rmb7BoW+RSuRg+XtZ/tclduYxP
Cmql0B142//gqKjvQwvFwf2RDQFSv6kzcnjpp2xpYnqjgWXof+m7dEeFGWf/ablA
P0VbatL0KAotK7yEfpceXPwR5uci2JMYc2sGwjb5ISz1wOpzRi2j8VSgpX89ElWa
+/mvu7X0A4lHYOMvbdaOXbQ3wc1+JfCbajPltKnXtLODb7lqqQPJu8j/XmRXBO4D
3DWSwQPhtqU6LgIJ1bDjMCgEydPf+x/2S41im+6ggwy2f8hDEWxPZeHylsnnn9Ty
UVRonet9eRv54LU5sfkgI2bGzHUST0PtSDpad5yqXs/Vko2XMqGhsBL8eyYdAmqP
jfpekfM0vKq/4QmoG1uKxqTOSnWvslQGOvSiYHtb8E//l04UE551uJGYvec0EV64
x3UhMjapRxApo4a19PhL3O95WuARIVzJYnH/KasB9LGFl4+zZKczfluI3blm+nvt
g35WfrPNZeaAeHxOdtMEVJ9QGooym3KC2QfqRKPFfom/dMpIQj9rv3IIIY5g53VN
vSPQUkd5NYFV/sJGu0I76uvXLBgC6iRQRUyZk2ZxHUArixasYfird6LpUYUaf3Fw
O9PeBiOXh5fKW2AFrJ31tJvw1i70Mc8ekZ6M6s233bwqktutaqmbF1XLXDqSPXJd
ryxSXSlla6BMoDy7cuFnnhieP8fylkorZvEhCRMfQTmtrDvxao7oEXgj7QWBO7ti
hpIlkCK3vkDpEVNJtYpxxXkU1yhuU8aPGHxR9bWd9Dq8AyWQOND978kLZAmU1YgE
q9CiBEGAYebc2fDtj2QBjc7ccsdV0qqFBlV0t2Ps+EOgaRiibi9dJ2jSdEflNtpT
0F5Zc4Jxk0lE0+O9VFbkKlEAdnRQyiVtl9ELBpUbADQ9JLwp8z0wmATgcZDjVpjX
UZyBHNZSVLBdS1FkMVQU70/02N/shpYEJftptYZFWWTiK3Xn/7Z1CDI/hBm6YgLf
efIa7T8tGC3iCTmB0kPB9mAod+VC/+b7PZs7+kLd8fVKKML4IQAu9aMq+Bi9PAit
6/x0mcdeQ9wJXUM95pMHcLrg5m6CtgW5NWA/JMugS0xfjuJf4nCkOzF1c5Q80G0a
i8jyZZz+YxVZOnR9Ogi4ovUgOrrcWoNzz5Wjg5p/ClyUjuXGmcfphf9OokeyNH2n
V5sY4jlo03Hs5UoRCqzKPw2uGEm+niytUWnnWItH1Dp+gfjqa3D+N3XXj69xnyaw
Xfv8C9DwfNDWCG0vaB1huhgFu0y0aXTZoq9pesQjnaiAA7oQm0+HwgCuNKLyUuHJ
vde6rhe6Q6Z9nAMasxDdSRUyv8LlsrFljSDYjjCZl9vkM84vzr3f0pEwxDKZZ4MH
H551udtiIbu5RmBUAUmQacTyCckoj/w7KieuEBEe0T6cYI+Tac2jPJx7fUVbWhyL
ak3O8tCUicSOYjk7epm/gd69OvR5rYuoSPzvDPaMYBJq8qWPxW+XVAoElJAgvO63
XVjREgIOsVr+N4YN9ZsBYv6+ithPza5T/kkTHLv6xrR2WavmSyz9CptC0lsDpDH3
DBqBwh5ZRNDqNDJi2BVkauoyPIhqblrpbqlA2J2e7ppxSXpJ3GUQjzMJNCqLUDKV
hjeuia+RtI5l2Ofd271GJ40UaiiMP4QFOvv86oiq5AHg6LKGB/5F2ZMF1Alvsyum
/kfEM2JuF1MxbVojOvRZiBo/nBLN752yt8H2NYkrfGX0ExaNrkX4iIQ6oPrFQTkk
U3ZsCkson5+RvCXcOX9DwVxMzhCtiDLXBCqtfcXMqgfJkTVR2M3OUDZNldnAy9w4
izEV9UfLBCcBeMv38wtNLyIL+JOSvp+Slop/8f/68E8d4BsuercIv54zoQSCAdgD
oNKZX7yt7yepihPi9me05dFToe0/AZtsEnikYbn3x2HRw1bLIe4eJXA9TIGiil7R
VgPKYgVOJaqLn58iygAUg3uJ4lXsI5yRMbMvjdeXXgkfR9qleBUAYli7ju0Ltsy0
XE0pYV40nKDU/Us7QXku1iPGRRWZRDah6GsST+bO2L3sY2zQHaNK6Nygpg1m1SPf
Q7jcNtVB5mVI8y240TqPWuNCgwWSB4aeUc9kCD1WXOEbW7tMtETJY2FaIXXbsC2k
CbNJ+iazrzCbLGjFbJ/34LWbfFD3+UDGi7/plJ8eVMOtxu2V9VzCisnWyi72fowd
CA3FEfrlKKUgDAJVLjBCYNvk8HKCDkT7ilEC4I5BdbzyPEvsPNj11FJnNRRcxVaA
VKbaVaxCm+lJcDL4ZSfAKIMxrAR+auo3bdmRAZqH0fOSCuBXkUR1JYWx7phkEjiZ
1go7HwAsa71gi3qCC12QPZ3A2AmbEtJ6qWdS0NBw6DxINOg3x0koSnDdb+kuUxfo
glcI7tCSgOlEGLhN+HoRWaL/X+i/G07Grxq6VPB+40JXBRwLxNdbhE+P8DvC+QEm
i6SOSmR52hIr6qvy+ACyakOHWWpZe7S4tFlWfI5YBQqqjW39HnHRHRVwjuM2pVny
Hv3O8MOc+LddDPy48PRMksk1TFxpoT7D5F/rnRo/hOr91sFuoIpN4105KkSP2AX+
1ky17ubRxyl29XLdSnztesH6eV+00i1mHri3ptUi/0gUG2YINndq9cvbqMR7ICQA
wZNrK17JBp+zA1xgsmD9AN2gDM3fxpbUceG/W7CwsS6dBh1CmbuCjnT9vV/5VC7a
h6kNg5nMxRLH+iaaupC1Hr2KYXBtVunJ6tOFO+gtDPSIrGlhKSNKmHlcoK7WYlAf
AuO3ap1WmvV18ejzoHZT1C8rctBODmw1k7Ux4/xCHLUXNNk2brHV1ujPP1UJ/IMR
llMpOJxs3PbhGB8lW4TkVgERVrhrMQFo+8lcXyl11OjMqRw1g615KK7o22NX5TNI
cYLgWfjS88rwMG/8NF6ZlOigXqUMYE4aeZLpVaQhFSk82mEXAavCdk51+gXne1qr
BEtTQSt0h1gAfRDc/DTBx0/neG0J4MvTKxn8um3BeXpAB9PYxOcEdGkCxAIPBuiA
xO9okpNBkLSkH7VQBhAuxMffbts6hhTgFc6vjWD/b38nW65BXqDdyJhK2JWfU0WJ
dEfzsTusgIHxpDsRPuSw7B+w1XQOVzCF4EZJsnTRaQMlnH81RVJfc/1ZC6sTlRIl
itq+600Icw4RKmfM7KCG2lLC6L+FuFfwp2j6AAvFyJzbmWXvM5S6PCr46JkaNoAp
slgzFysgZY9i2FFE+mZYR2Vkgwd+NEYerGgL+jlHXRKyL7Kvwb6Vyu9W4LLvy5So
UxC+/dnqUjhpt/0N6ZyRCismMeAmSXKQOfhDkkUu8J5TbfgVgl6Eyqmu+aeq7Mql
Hu7UGo4UBNmo1CIxxrtf0WEdGxNMIjudP0AyHUM2PvJM9+UaAiOX8oAJiMgvk3FD
7uHTp1wsFRhoZ2vkBaEyZoebnqRp2WIuJkp5dSLGfDhdVa/gPodltqtZfHK7ChSi
R+lkAYS8HMCvFlQN6bsOFio04yietqhY5akMzg7qJZz6yIRH6BbpfX8jfkof7rEA
QfderSBG9YA3j8kqI/bYZScpbyEyoyyok0APE18l//2bX15HG8fI0kWFgHbzVELN
zJPtlfqf8/1VF0I0SOWVLk+V+gIt/Lp/fxSZF5mn6NTl6qqMyr35ChrjwkGBAyE0
F0WLLl5cMISWHT65azeEk4ofmjD0ud50bHsH1dZ1h7rMwpGizmlMJk+zhPCRpk8Q
D10NAq+K9j3kqvpw9KjEQgwQQ9Bzu5aV1odyRfce3HpakrkoHZGQOEc5ENwO1cCi
3F1pYbULlQ7ViL7gFlA6Z587JRH8pkC4afE/8lhj2v4exu14aVsj0lSJFo5Gkxts
WvK6jug5SxsZodVhfKqWB4FP36t37RUMLlWlnmz9rIG7cjB/1WurC5IpRBunX/Wm
iLFoAv/yd/KrvzXddP7TYPZJ6zr1HwqgoNARH366w9YSHCgBEmgSYPclTnlPJQyN
Mp6wSWfpiqmiWghdJgPTiwV6eR7JKHEAEjXkPgTPO/epZ3ELl0+r+SMHIW3muOtb
KP3zAbyZVTuLJyl0p+fa7w3h2otgh5NR917a/7JzLZrX53XnCiF+Xx/FYYXtBz8c
wFyEoNG1eNarfzeE779sjLFHvMZ/9HGd9XiW+65ujIH0m3ak4CC2cwiN6n8Idl0n
ty12gVNoSylQLNCsqNATWdSu6yM1tEZQc+I4o1bKXgcyCbfamBOvQ1+AkIhLz2fQ
cZOZXEz74XFBc8jE2dx9zmgOasSjQkGiabaKBNgStobkK/FIf6SfJHqShEQrX+wn
VsFBas5/SnylMoEUyzYPXNFXfOhxsCuiKp6EKXBywZFKityJ3YlLSCe6ys+aHNOl
93gd/fBwhR0h+BpTQ+zTaUZ+OcqBAuEp5BxgetesJuhIhClWwxHdL7FvqIDFPTss
wPmM8M5KfIvTIh8PYrD8LkiuqI6VS1xzac7XJK5Kb+r8lMSpU8J/bE6qoCqYn58Q
ZwkUSV40W5acpYvstHQLokxkKrMYJr2h0HTKTPQqOX+qP+Ya+lhjNSuEuJuqCWu6
VwaxHrpD5t1qTr5fNjogsqLqbdigQxYRpEoiXWC/vqW8nyF357lQ434Dr2jeNRtq
hsY5GCGcJqEv0VR6pSCbNlQyK21Anr6mDXswqB8ITfg6WQrX1ASWfy3U10ynQA7K
KcHn/sYyfULcXmiE964pMV9A5WZOIhCrn+mnI0992ROLkFl0l/3TUZSsD0HKAy2a
fp+E8j6lAARV/dzrIufGa2yRodEJXrOVgXTsTVGC7M/QToFNC87z3ca1vkZ1NA+6
JTUR08VGBy5sdWyFhePIxgB/EB96RiLeT+FqsjfcUJsgHrWts3vrSCUO5/FXzUAQ
tpqtNU+bdfF6Vf3FZpgAECTSS9z6FbiXt+C/g+hYwvVaA2Ovqf361cHQGPqzOKRh
MZMvJ9psV0yJfk15UrBPpESq8TpTGkXAtDXtk2JmHO/SZj3j6ka8WLsvKQELnl6K
38lO0ovAsCjXXIFAETZ7TDJJ0gn+LpfM+26uDpAGoDFeENUEtQ4iE74IBLry8EFo
EOntY3rGbxPLc9E0WDpHVU1Hgc9hGn7whrX2ipCwyQF21E5wfXpC1gi8D1qcC+Uj
gHZsPPAhHmoCb45AvO0g1ECINbJWYmYd8yZr7vxPMNDt/Kszp02yA5/NQ7ROrLL+
gG/EWvOiiNT6ezgIGjzxZaOJuCd20Kj5Vh0myl/WNTJ3rEmPXfu6t1VeGH3J6+o2
U3LIyQoX5+WuOoUtXmGNGGtbVltQyPZy0N1PBzZwYavVvbOpF5jpIPMLCmGGMlaZ
iYPaxdNE5QmMQUm094G9OpiafvPeRyx/Q+dqnogiUkBSBeKQ3+ZGr/c2bE0Z1J8E
WXUBlB8KBwhk8/eySJq8UsXX4FTOiZOjSfvj0G9CO7IoHhNB54k5M0GhQph4lLAK
ypWEw0nQXgQcKISIB+ZjsmnaLfvDBil/i17vwmqfj7B/RWDJDzQmXuLmvrACn2nh
9WELJ1uhfVSdN20xBiS7xpWvJ4axrA+GK3vQerisg7TycqCdja+W8ul2so6E0d/k
0kUe1fk2r7x37ia7DUD0PJjlG4+coYw+HOBHYD5+WNUUlSmTdo0Ljaobewn3qcN8
t6DGWQnPei5PoiQTCOekcaLApGDRvwoAflD7veRp437rAAN/W1WVHg91U7umbsUS
0H+3NWGIP7TdL/usCky2UwXGSSHS9aloRqIprZDYrlQ+oqaOxCYbYOOj9gpR6tWS
LQfJPs2OQmx6Eown1zrRQTdenHtq/ENALyWH31+uYYeMmStEygaEF18V5WspWXoT
CyFlLslbH/cqGcDI6hrY6+vEBhsJXBDIN4cmaR81bNmeBjtadPLm6swAm0Ryuq56
ynQNhk9hNyviRnTgE7Pa7KZqP+DHSCjnHRjdaEpNul/DD6oT2BKak+62r83y5qFH
KNcn+CEZTAYr1l0HtO9IFaYIkY56Ym5yAkYwDHDJP7ir0LGN0YyT6wsPY7e4sonM
XU3b8a5iAqWGUUASDbVGOiZ3ShGlg+HOvcFfl7ZXyujbkgKPi6xOvkOzq+oGKiy2
YEXWpOx3EqifO4J1q5gGYs4NBgKbT0+whvIXfdWPJ5/XoeVkOxlVtA1LubSMCCKu
PRLU+ioHL7rM8j2qUdOMVcPyh4tBmZC1cEJ2vzuH22vHeJWMXch9+IrjjutpeTTa
QBQp5FZW/OD6Tv+/GHQ+6sRDmiHzQpWfB37ZbT9KJMRxq9gCKqeHj3lOmm2dZ9S7
glKgYuHuaOBJSDu9UXTqkEN2NsezFoQF9dF/9MiJabn32XFXjnMcUJe83BNA4KEJ
4PKhHDWcpCjAuNece1gKDkanbJl96B9zK5CZwCFcG1Y5TFemgngv21ZRPp2/gWQE
Lk/L5fxb+syzP2Bj5YB8+ZwZNcrwBnBRd7A9VAD93pezMzJ7doaCqA4i7KqMe8eO
o6qJRSNK/hijbGWgl8rO7dbJAeJp49A8h9XXPRTcWIOsF9uklRT6MXnb7i+W2IUt
mBEPk/bl8SjR3oo91GyK2DmyUIjviToW2IgLtS+WDL6NFZ0T/ayQn7e78QT/eqXl
uBhbG7GSD4ADZwRFlPXslYd+/T6xr3fp9SUHFIjv/isnb1J5XrVkutkiMUsAzIMu
T0AU3kNWTt4ghGszeVh/gd/vmCcxhR40LDzIc4GxgEX2Bh44T9uqCI/m5LS/a/G8
eJqyNf6bVPdus3zxjN7QyeoO9P0ZqGjI5G+VZQOlGT9eMBCW9Yl5dULP7p4qLgfC
N1bBT6YIl8kg/eDcPqP8M9amG0+tdXyMwROx0Q3c/pe4muubbmetqH3VN33gEOig
7XBBrCNcUKD6C1VmG5BuTpmEHmKCYWFDh7C+BZpn2eQDxeaia+LoVTVIsHXvMwn/
tIM27WPMSsUHNxJ9Juz+IoKSb4DvGjk5xQL1hvQquxzhLyHlQNgs66MRByujJqI9
TML78H89gI2FEPPC5w2aKuJ+lvR5ff/OYyaUlyFUfF9lFKOBIb8sMlcljwSwqR6L
au8md+8G0YtGkQqzBYqr+GhtH5DyzrG9SuzjOsyGU4UuFoXNoFAgQ4nBX+2B5iRi
TTuSkdAtyf3gFUP/m1SrWbjcpf1J28ttF8YmDKc78es0PSh/RHVaLmCSKjLREPjS
9aijtmNPBOGRTLZhd99rIPtNPjLFqN1UtAcOcUnNsMfyzkTFS+M1jzYEUKoe4bY3
9Xu2i3WB4YVDNFdutbiESnu0Gydc1r1vU6d0MrY4uRSK/gOcJ/MivuvSKVtAFZVU
omRoGk3FTGO9I3ebf7RhYM7B158vfaaSQn9nO+qI2Uf9Jn//DzKyxr5YXMfeS2CD
Btd0KU0Z3TUpqYREcKrXQ36DKDBIz4q4pt1hpuVQy8utwt8lFPvvDMEP+D+/HEQ3
4DH8e89HBE7YNdFw9urblaxBz7INnElq8x8QlpmcWmB7FsC9z9HB836EXMHmaWZK
v7aKYaHTVyZlESlqY1n2qlPVVI3yLINc2ITrwDn1Cqm/FSjqX8P356zCvuLvzRvz
sTMkYzqpX4NU2nX7T+cYyd8xy43WfaKJ7Y7fvREtuN/TumNDuFhOCHZh0EfVXXUc
5K6dSZIChWdw+Vg8WOtTGoMqy87nDoOES+wchS9AbqBCPGVvMoeBCvTbdTx+6VoH
WZcH0qra7A5UnqUR9ZyUk3vt/jMoRkPGDq7n/6RBjtARnzrBxrmowsWRqUTUFy5x
ToBHfYskmNQmAXlcTtII9qUl77XWILw4fCvi8lY9UenwiZRnb/DISFlKwvGElnId
BbYBIyoYXRxlYTAGOrCK0XrT2sGUrfJYKNvVbsGjgajBXIVcNhIR/YAWnnbDiNsB
k9fkH2sCP0X3DGGiOxsIim/EZMLZaMA6ZtIMgg/As2Dr3/vcO45+ltW4jE2tKF0d
9yZLiZkEyCNyQt9UvvaNUnpbmeJ04GaWwb262yQCUnHTkpdZbU7nlfyLw6CnFDmz
YeQIlwpZmNIHcFbQEnd7H7sQjdqEs6vY+dBW+zZqDSax70jgLzIMj2nJxl4vop+Z
IZek4kuaYCaSBUuDhLJyJIcuSJ2C1aSmMqCiaqR8i1fvArgryOJR7vxxv9I52SOV
ycZgQz69c2GKM1Zv4Q7+o7XmyoZ0rPcwp6d13avhMOsdjWeD0f7CGDbsBOjxRaYr
yFTdIHsLWOytdXqOGiq3gylib9ph14e8iLoAu8Yl2oR/ycw+yDPJ4MrkMXUdBKI3
7XX9y25gNZMsPFvuVwH6jyd0OlNODbEHL7CKQAtji+/RpmHM7K7/z4JUO/fZpUEl
LBLbChWBQizHoZhMTSxFeyOJGHEdFLBcSy88lqnNQKjJd27yy7mkUYzYjmjxS6Kh
w7dhb/6WfLbVF1vfCf+y/2C3wOaVCSSFhkseeLxhbRt2SvFDlrLJYeYH5SGGW7HR
Zd81PQojP1YPGsDV/dI5m2sQ9MFBOSbw0wyijkle7yYN6YvMVNfu4RNK/PCku2uP
XNafIXHoREe90jlEtIYBirqFc9fe+mzhrX7gJC/M0Wm16yWF6eY/sYQek/NM49Pv
mfjySYo/Sq0f4F9MB/kB66rOJVGIK7qICOXYsypgsFloxwPC2jwxsjYeVN3j12Yp
xB3QKeLK5dCzrb5CyDvJ44trajE8KEdbIaP89xywc8Q6SeqqJBT2cBrrWn3jX0kW
SHy4xIwrOxHVkajhhf6VQpTJ+dzWen4enAxqcd/IkdxbStB8C1HQjAd/SIPChZ4Z
IzUZigFvHIfGB8XXg5o73d1uh1LGfBJA9WAMX3pFsvZ8wpGt/0qkMaZCHa0skqGR
Y43BRF5XfJKmZLHFMGy7LR8ll+Dk8Q/rl6c4tfFoA+A5YAqtU8iQzk1QTOrrz1qO
yhb73pxC/4kqKnfg67PxX1gkHTzNhqveDw8ZB6SUBsmgSeoS6mXO0gFVFChlj2ql
PWQlpXSnIbpT479mcV9EoLWcPgBQJxFuBOmtGUEwFO+UbtiGEheZgkirujpXBwFd
ahCL+P7B0FknwceNjIUB0QU5oJTlBY6wLbar/weMBUdUedPL5dbXOIuf9BdvIbi4
vzCrqTXVA+eIscbFMXv2BPxV6KNYpAj/DooTzDL+Iy/Y1QJWq2nIJ9fwPUHFF2AT
dtmurbu5zIVUYOzaVQHUBbb2e05t3cJiPVolsW5r/WvQXqmmFT1okTl5lAs2gTMf
2VuFvjldM4uEuLTAH8xc2msOQq2o83hOs48nI6ZgmxZQtxTCGr4dJHV2b79DM843
fLqxs0rZfVox9MXI6nWGGGv3B3jXPq+gdr7hOyxyp81b3i0B5IXRjd1+T9FyRLeh
rpC+/75QmEGUmuaC2WoTtzd1WDeraX525deOuSlzSfUqyXD8ghxHALylRgYTevaQ
luuO3SM6Arp15ZYVAUviImmuV6YReNIYGf/M4lLYABpL+gJci1heAn5ECvLW0UYc
hmlzOQ5hBQtZLetqXgZyFN+qGH7A+nMYjM/hPVI6jAC3ihevU0cbQIr2DIN9YkcL
mMudTSbI/jWcpU8ggUPT7FceNsvJH4r6yVOHCx48CpLR0WvMl3Z+5q85sBHYqRJO
Wi6EFFYdqkNlePg7V1roh+1DpejpUhEjEVKRQRsuJVnO1p5/9YBCkUYmBdMZedyj
FCxjofnHaZn7oYEtGxRoSb00hV2RzVijGU4DVShYM6S+S6cZ8YpxCeZlOE2cUNAT
y8JJL+7+lG1ls/5Nv/fPwE+LWthyKScT/hgbOmuvhtnYmRE3xgks+cKM8f80cF0j
EK3VZ39WTgLhzTCDYa3GZvk797X7VIOPd4T+B//UwL2zu3Cz0vZJUrZLTSBHdMPi
pTJNX4ltIbdc8frJlj94KRQAZOfrEcV+VIp9mYTzSgSp4QFz00SZ5BLPfeLVvZvm
BPXMfyewoTBtzt5u25WABovq37BnuRTSCtn9YdDsRCx0qMh1PUJIHEoZ45pRRQa6
Uehim98ljoHIVl1qZe4HyKbv/TT3/TjZmap4GyCJuHxMsQ9FG+aqpD0JoUqbZB1H
U8ld2VUXCRfOVDE0UrVuoTWU7DQD032WxTGS/W1zRv7ItWblWoanmk+MrRlFe5i+
aMxYoM9AqxMDbIGeVyt/vtdyJKTI3/uM6duiTmfUfgklhEoU1e4mAhKwMNttddgT
SXXk0TJ/9ZUCRdA3h7lqlPS56n6pNTei72uHbOQlJqsTaO6EglrZWU7nLHOo+BDY
XSrxKpuRmz/Be6vJyEDc8WSlIAte90qaOK9a/CPDOrMr2T8Xy05SNBv7Vi4nRrK5
4J/5J+RBINzVU4F48CwH4Y9+1t8+ii9YyH7D1hXrV+uCLVuo2KiOmHi8tV3J5Rvg
p3GlD3CuryekjwpqaPKuueY3KX4ByAuWoCGCmVdXSxOiovf30w1Zf4rlithWoq5B
4ZUUTmht3R1ZL4PsuqHjWHDAqXzUizBfIHJmBx3qsEAkidC393ABMriu2UoBlHD1
9HJJwYq8z9ijOXHp6lijuNBCYoGOQRBTjb7layRxxvmr4orKqu6y/Uq2Jq3fiI3h
NANjQd2Acg8ak2UJy21QS4VoC3+83F83S5PZt6o/Y0ARcqh918p46ZlCsYrg9iBy
VVBQoZGkKWJsCYsp4jfEoVcgOxSzGF1ekwQkMt52tC/7aPwyVhBrlMCJ6HLKMLDW
lXtI0bTm9NuKTWtPaeO4JJTSXNadNuDX/yUnItzyIrzk5xpOz2mM1EqHeGQ9N9o/
F16kmRtoibsvj3yH3c6WlZ8MNPUqu9WzAxJB5TESgoNESRUCtgwqBpEVdZnVYRbu
JF5i1o88w90zbwgxoXNOHyhYVcHQiiDuHfdv78fG23j/QGDPFTazNeLCNHPO9Im4
uKP6mSOGz1G/gkpaqLvQ0K4gp/nXLLd/BYHSFSYpl0CqeFsZ2u0AQltU1moEjZVS
piT+xDbDrA1vj4KVs0U3uQoRFroJeR8X8n5UVHNpkqqeiodskaiFtb7SazXR62Hq
mzIhCSkMFLYb4qWUJjemncSp78j+7CY29ewrWXaZg+nOTnMBoEBtSiLykyKNjWoH
Lvs0B+NwYMomMCOrS82cHSmdzbDOPNIB7NPDhT/TzSei0BVJ1WQVYjcMWq37Kkk9
zbvTNsNiKicCBBG7GggUJuNqBjKHde7lM+ABRgvmrZWgVz+88qEKfcxrf5RxNmNP
LVeyxAu3uMCq0MO9EQ7kJg5pyEye0fFVXIsVv5UoFoiM7j6jNrAU6fJvICnqRLcz
hFE6oUBG+8OQ0dVZT4x5hoggGpFKzPUqmzVdekz5w3vunulnLHwibWo9zfolZZIc
kxszFyZQnXLOgRa28OE3US/jLpHp7fJFLpuB3N+uohgvbdj0sNb0q06pzIvv20ew
ufDq8ww2DW8dbuvX/TUFRn/NEaUp/9GoDOcNxOtvCZPnQfbShBheycZcxQV7kucK
meYJFbyVqgCoSsIBx3AGeyWd2hiOxjoUdQxy832FGdFQ9p1CGFkxb3rn2irHqQ1l
nIytX0EBLRp9A4mdcxnr4CgZs2gzeZLNXa0mvlJyygZ0qP2AL9SQmJTCYk2ohAqe
s1NFuXbSqvpj/sgfLbwC/dLjtEY+ck/Dzxxv455VVcOKCkSkYuXuonJEqzsDxkPX
pnj9eVJdue8bJiQRAmZqU4jSVWfTJhEHrzR1pyfw79jLR4FgQmoFWG0Z/d6f2UFA
5M7wPIApRRzNF6VTUArNXPuYL1qrPCkkFOthyiaVeSt94cGdjPXTQ89qIlOvKu2x
JYmnBF2jgWQ4TrfRxCKE+ieqHuLtf9uNq+9pg3FsSTyMl17HRmy8zUhqdY/OpqQR
mDG+dxnLvxNkV6vaL55wkjtgqyj/Kwpv6fdePN9Qg6Cs9G2M/dHJYUvq8+7OZgYF
C3hBx/5F3ivdsBSt9QqYf4mluaXS5vtS/sH8Se3oxVjPfwvKuv+ZxgsoXKhUDV4X
mx3tMYcwtQ9O2Z0wtzH/0i/lwzL/juX2WGrI4fzjc3rfgbifKXNWoVPtwPBHQE8N
c/17TyENqHRtqmK0hPBrOzthvbCkiQHXSBcGjVupnk+pXsUwlHNc7YCPUAzCvh7K
0+b8doNNIm4p6m6osu/ULWoImMzPadXrw5iCNU2yGPaL4shIENoszvcvJXf3XUgp
Gey9xyeiO0/QYXfa8H2ZW5RcM02U0Xkmo/yOEvnjGqTOKtVhvhhjRKc6sL/moyNj
rCyJ52+GzZhAVa1EJcluQq09duBURyHt49fefzN7JImhGX3g108VNKJSm3W4BQxW
SrRUOjit2SA49V+ZKFzIwHLaQvr+oMsqkTuSb7t6ozRlHnf0Z3KJFfNd+XnYKGL+
N+jufYaODbXlBiV5PhriZPKcrKT1Cn6QeI9X8sprzztlgS9qeL69JGcfviflN7ej
b4LEDTc2S7HAOtN6hLcR354SOeMZWCQ31mhMsxgfLB3/0uvzZAIO1BKzOLTEPL8o
bWV+VJHkNUBR7x68EuRzib6e43ke3bMA5oK+wdkTH5DlaFzmdRi//NPaybzMYhqD
vhRNhYEMqNe50i5qF/AXtN0fu56EYdZenuoMCCavOxhtCaGhxsJRSvFPi0saMHZM
aVMVx/oJfj1UgPTQVlwfjsyrdPMVI5r8aoClmL5am6uP2sWK1YDnprwM6ds/nv8N
a8NY5PkX8j2u3cL8TOV+OykIfkXbM+bz6psE/PB1cJ3Ef+mx6McLDq32qYQSffdg
Rv9jZMQaKywmPrtXFBnCnXGF5qRvd4dTrxUvmuO9QqE1KfOP7Dz7HaGhUrrPcdAk
/qnevWkJVb0+IOKDldtkPmoJlGGeS68D69AM5CJSJIHvIY+b+nOa1xcr7lwLm9q6
hBNJPEqSBOnWaSH67FrW7/Hmpc2WeP7KMKcYaxJYGGFHyCGAyKZKSNYfTc9+ezxa
+4mkVjza3sbZ4knDiC/e81j4P8EcuKCl8TU+YCMS5IgUK4D80BagO/DlnIBcJ99o
81jAc8DF78UdXUVtsiG6gg3Mj07CneXudwz9t4f53VZgBpVZSEoKKF4Pa7ogDjej
Xsfgm8W5SdWa9qdgRulYHKEAWDKea20GACg72aHS/cmpgC/2NLg8AzFyu6p453ib
FuEUbi4Io8FghyFrIdzFPlkpO+gS/aS4QXghn6PcoIt3JC6xcESRZoOmoy5Asens
iLy3nVRH8CBkRAGmVnTy+MWJICHxge0bJzEv+a3ufHwOH0v/GmRWR0zEYydMUwBJ
BDAV14ghy7tkLn9Xte2uT/aSKYGHa4PnHoj3tzTlNI27PLvxkFtVJisdrKQoFVI7
hhIbeQhnNBkj2zd7oRBX5MjNvNyRGlkAnF4YCxSQZCTLEotuiwGCtiHDcYSjhQRN
X+xle20zmsUeETp9LJIK3AfaHc0WB+J2FNFjiRjesAaKZPg4eLWo5WWboMxPJkqG
NIRow7OiDVPL8+FYbh2HFmce4L9VaYdslEf8TApLF4tYhQYWmzNLd/zFOnHkIGM4
wmMxJLeuXCrLS+Ir3wPNXYatKOPoji2G4I/C6h/a8EK8JX8FcNAhEeHnp4dFRT+h
9nV0bQVhBkXmGO0Z7dcT1G+NragkGx9dTE7puy3lEkNVWAj9bA3MxcmhVTM5aEF8
mOaC/1IEKXqvEjjEYJPwOfVRL7VlVNTKA8pTcfg7L5pOx4+hbI7eHCYgAaGi3xkv
vIhMgoeWPLV5IBV9iD0+p5KDL+P76xDj+XsJsiKaUr+yuW2ZWbWSVfdBNNrKgW8x
3OeCZ1TONGfHqkF92QjcWHvTgyOevaSlPEtFVi1YHlMR2WFrErxK0hEX6PabDjds
Q65TmxG26j7c2Mg3Fxg/z2O9a/iZKwWplYcTRmNYPnFNuG9CxYamYzRky8xiugqm
Ono21RHW9yFdzE1huh8o7b9GpSALxGQVsOnVF4WGA0dHRn4TOhs8w8ozzq6PTL9Q
sZE3pYMjFQZGEspAsvXqGkq6H7OktCR0EC8YsuBiOEzvNARNPGzZtztm3xac+Awl
b98gGjMNVXGWOqy0lhoDeFftAdF/irEk8jVimsYxjuAJHnoeUuLJsGS7EDdDczdA
lzgopZYoUxZmVdbbZnn8M8gUPopMzD6gzAjWQYF16TPUsgV1zmAi1zmAqWLKhKSw
p85UYa27bvcwhqNYeiwe5k+8CSXtxI/ewIuynb1lg8avHk88oyceU3seyRKy5RRQ
xmezJFrki5I4mgoZUO3ZW1/i7Hl8c2yZRUyZGOSdlcvA2YiXFC/7CG1HiTyBfmaF
xyietr+XmOFAwJQu9AD+jcCCp9wcn/TGimue9cBNbSVzcB0t2O8EcFAO9Gjkcmn/
pklqacmnir71Dr4ykHT/3vl3xcYnw5OuS8FFo2MmvC8TUokD+EggTlHliDDrRtYm
tbYJ1ozKi61o1OxOQ1pO5oWTFqCd8Qz9hp2oEVdhzFeZxUrxemaytNDiapUWO0Ti
PM/NnX36+MmxbP2CBACdeDunDofZ213Qs8wEk8OAJy2fsHM8yCy9NjfJyEMRKwLP
odwADdhmjgBqKRzRG7mhjCgwmyvfvZ9Gh7YYVMHjqCITD92YOkpXXSbPWGIJnYfR
OAiLxZjsH9Qm1wd4v91gTkOxcryfp4mBPIT8GwNPu4WuEJRPqSFarxfK7gby0Big
MBbX8XDETT846kARt5vbhqYS0o9UGNttgB8j9FkQJMz602eBaf90NTnYDZqDAply
wBe46d25R2eJ/Xk25u4qTAdeY3w/GdB4/QaNT956z4IGB+kNnoDy3j7wRRyCp5dk
R3URLIBZRWoIVUfHjlvdLhh0EiUdqoabBZM7lXxH3ier46UhXm8amcqZX3C+T2zu
wfNKrWa0o8w4SiwpqxOlR5XsiIGxc8DZJ41pm3iwsfl+lzzbfwhWzCf64/JJnE+g
h+I/p3jP9XdnBq/YCi2lPFtElJeIdQa+pXPHj1iIFbwHkCTdgv0KHHUvqD0PArcI
kv2O28lhDCxA9ZqNLhvwijh1fBPe2SPLgXNdH+O2O3ioyqTg7WT2joIYLFuQaFmP
gKP7lPVnsnzfOv9Y5KSzMAxGFDW7Gw4YXeMBcMSOg89aRN50GhInxk2HG1KJzbx5
ZdIxojMDab7KF9cZPQ0EAIdTDyg9fcSKkdhhQ8+J99R1HqlRx2hlokLz+KwbkqA0
pIXN5jfyCj6qwkv7W7Z1sckHgPTF+1u63/b8/GlcbCK8DIoJ+1CtdH2I95IHDXvM
oSA9l6PLKrQ51x31Xi6jLpTViKZSOiLn7vGrg9iQmW9muXE15qsCA2w4pMwLJ65E
W9uHD7XlXrm0KiDpZjpjOXjkj+5c65gGsP5+jNHPh4gerpUKVLUauNaEG2fa0ECG
5CeybfnGq4ZPWNalyGWav5IYL/utQo29AG3sA9FyogY9HMTKTs5RLYkH27If8g6C
e6BwRDPXnTpvu7ojCf7/VfPCdFGoyKF761Yqn3qlGiWM0uWhXtUW5hR2BAKwhedK
R0HAic0L1hCnLa44Zj29zktrzwl1s+OgIgymLen9vec7dO2t4Z69IXMWVQO7ty/M
VhLuini+bxb0tP3dj/f9Flfu/F0aeljXRyK5yFmNT0RF1ulHcQyy4UBd3UZ39F+q
n7lzJQyyIpOgdyO48UvkLfeujIeQyxZNdI67F0B4bMJYQeicZwo2Iz04UgbBhlWg
cM+l2sK5V+bqxB4MthMRbkspPAxyX0BXS1viul86nR16zPScm1JUih7Ydj74G1Gl
+amn6S0UqXWwzT+bsKBcdTmBPBBN2oD+sdK2efIeWRIeYO6G78e+1IgQJoLf+Quc
3NmVl6gwcT59o5VncQ0MK4P8mTOByrfizAmGVwoKh3hYhNSM8MdGcP9ePejn6vt+
rMzsY+3FPXIwbv8P8vpNCnf/QBu3ay4vZyHsd7RiH5MTxfdEXKQV1/7JtXXNCk0r
OiHsn+qUYzcLtnlKxIFbfwvA7pOBpGKEyf/Em11NjKYJVpJVkdjIGSCkV/iXwjHN
OiYqs+8fY4eDjHKusITv+y1pX334hEXosTFRaB4aWe9/E8xKBAMh9OCXaoWQEnwQ
DskX5cRKYb66BvH8e9+E3YnQynqSbTc8AvXmZMPh56xcouiMarQZGmGkpfJA2csu
vdhE87AlqukA8pB9FfVpFq+qi0UKtOMmpIlzKdJh6oMR6ZQaKMc4jAABo69skzZj
srdVghtMgUHpnFhTekSYDvaoCbNFw54ij53VoE+F7UFSCPKepqapn6IWGiH0jYMa
qIamFA4FZoI2WMFJYJdu4yBmxwtW+Ay8StS3qRxb2EMgj1oPboerjBlf0a91ywW0
bRHOGZdCU1toS/uoLVpA5C7R2EJ3f0jrDVpFhA2fbBtf8LpQmZxK9Y8oom8OgvYv
P7Rq1G0my9MzUF24AeYTZB00gmUhgeCK2gtrHe36RchnFDBPak5hpgiWqddnz8uV
6d8Sdgmy/9+9Y4cayK3Ry1ObMPcmA4lRGovAZPM5LVfOr965vqAhdia/V84UFzTz
VwMd6OHq8O7O2Lcrc6DUWLVWUZztnmZlznWNZf6RFK3Up4Nwlz7/Xjg82fLMAk8p
8PvD43M6L71D37084wSKEITYfGewVdfpk0f3Jlmii8U3GT1XG3pKEArZCA1AvS/G
tmckSD1HF7emX7hEZI4VG5qg7CBMnLPWm80C8yWnaYxSf+JxyHDjm7VOVLkgVHc9
+yb1gFe8EYhQhXjCa9yp8BcZOeHDNrWktQtSuqsi9CbEbVz75oNdQOCXJ6u7VHWW
/Mj/z+5INyTq3RElbvB3sK+r2EbQZ5xjmNimNqiU6cjXpydtsmCa9fR40Y5FYq39
deWMUmDHx+HykwBQ2pr+s9lVkjzpoj8+59WRz5UMRLfuiB/p1Su0Mgd2e0OObNlq
bncTgStcdI1U0atC6DdaYqZvVqADqOZ04L7hIHJtH7fSFOOROdG7cRVeVbqtdHXF
732nv8ZcnImn729b9K+RogLm7/c7PZfb3ArlaZmSKcw0y4D38izWh0sUjFNDFESq
UWU5QIOjAb8EnzRgKs5nvOD8d+ko02IEk60JBq4DSGBlKFgGxlFyZKQ/yykZThvl
6T2JUuIT8c7gx1Rcrz7YCfYIDSAgBXCeHqUIV+Sviz3cLWQjeyI9YQ1IQU3HX2J3
GigNh1b+DUcCbXNqRYsHitJAbcq7F3AdPjHhFRMf9N5xIxGvKNYAcfSmkdSwvv1c
JSYrd28uz/Q0G96fywm18VsspJOMSIl0X4OSZI1zGXVfvwsylwaturRUnakgjmfR
tP6a+upLYPvnTWhasejoSqI8ZGq2SxbgbphM4WlkBdf+lJUbD8qulJLt3A6gV/Mu
o1oi6nSWhkkzhrO3FCHADHd+JDw1z/4VLCRqafHZVf28VH9kzHrkzMZd9lneEUcv
oPBTV+qvpXgULWL/ElMdaOtNRJprvNvG+m5o0v/8t+dudE9gAqXNFzj9+0sVRoz0
d6h318kHZ3+fizKwlX5faLMRhGiJKOVqUrPxbqV+p9ALbcNIdk0EZzQ+8IQeei3A
bfhUe9JrRWFCCLJgD6oPq81OLmRo8Q9Dcd8DYhFWY/jaD89G/G67d5Um6aoKmFvU
DegbxPg3rd617oN1axz9prV0vRLKIEinshsJNUf4qvHCRew0QivV06eduGmIwLpn
Njy00eZofnUMNK3+y9XfYK+1Gq7MeAsdUOh12iEbLXraGx06nYKpZew7yhkh4bZu
Ml+HXxkxC50SOQUCAwI65Rsat0kBqezxi9ZX+4hx2sdZTFKYtoTrfB9ahFDecPEc
RIuIF2PpX/vzOYodWl29wKDERGWcjfwjln1g3DeM2b3eky7Hv0IHG5yLg5gj4Yrh
VFC6NJdWx9sDz3xF1otl67SvFjBgdc7e5+fviFR47oGf5rrDLLSPCDtPqcs8OwH/
PS0BrGsFXmySt8HjOLTgmX+Dt7xtyf6FlhbI2Q59vN79SgD+IxLPu8aYQNiRwnPw
fT48p0Wu+fyDnMHCpDGh8LhgxClKuyvML0UXc2FvNY+Buu2P9Db353I5yiYnVYpG
EIFL7xh6FZ9jBKrF/B6Y4Xw0hf23Io9bpr2p8CHvxxz3U4tCrtu8OgnqRblHrvZq
pyvgI4QwsRZwk7Im/XqGFI0boFdyb4YDd5qcMaK0L1iTXK47FUfgt2oIObuiklZK
+UwWyGIkeLgBEUjpPYzfUp6EQ4lcQe0Dk9kJyFiOACBP3CAHpJ+eLRNkdcn2lRcS
HhQdLf3Ajb6aVJiJJ2tkQ6Bz9vw1sG6Oy+DbKfeg+SIbfQC35C++OL9Ox8ynzqtB
1ppKPvGGIQcgYelxYhUvNMff+odxEHjtQYxnZH4ZBCwwFqKwcQFWKGChtlADw9W8
7QQnN0y3wDJYFDqeqPvlWCZnozblPK6QzqD60nvoUmCoP8JpZVjq6P96ZngVzVLX
NeTUq2GHHelZtmD4nU0KSgFTWfrI6roiITpYAbleHxIdbvn97k6gXHEmgB/DEO+w
XleXpzuVW83nhFxITJKoxwm0GK+/lMfZMs9ysxco/HEH0bDLPNLjyAV6cl2pYljR
Rl49V78esVfQ6mFay8L0icNhNRB4jgq1iwpQ4Q7LzljkhGiSfbBxm9dcULCtWItJ
wski/kztaIN3Gj5Wp09QQPJtBRJ0CIi50GI7AXb54EYg7kBS+sHDPrtjE2ZdLwQc
mfE4grjNk0nI/0UFEdyet+ZPT6AlQk+KHZPSnng883js4bAMdzXrPg05RjFuikCW
TmNtDM5HhkpnGlPZIvQ3ETeXDqWn22Trtha9r37xNL/nA6GqcBVlJ5wiNTFtxOeq
tkpSv6roejU46stqahF+d8TbZKNttQFftJSQcpaWYsd5GPUD9o9jixevzapdtPrN
qq8RQgVYNtpiLljbtYN+0ZcADKcRCwuaqS4shaojqtgwNc6MYvfHelm9Qx8mtmdz
R7UnJiUcNQyYMTatUqPPK9CtMf/DsfusQZJEQCSViWDi7MujlRW8QS2QHNWSjByu
lJiLms0fr7B7ecziKms/O6mTiRXvM4e2Zo6dNsdrGz5woPEc+Zon4gHng93ILt+a
DpZ0rOdJwOeyg4rGI3gWia2aXL5HbISFwpawwQGSup9pWMLBioEmYXkYycLgf5Gb
h00Z2mlF017BUsferLNT1OQrL4ucFI1++LqpHTp07POpJvUA2hPG6suDLvXFjdT3
yjMPL0BoeNSWxrhFGbPyjd1qbEZA0mjdnjh2HtmtCnBsjf7RoeIXxYeJcjYo+Hp+
epCyNVw/7YHpwkIizUxaXzt+8dc/sg63ctUg73hT0eTsaouH8CYk4XoS5i0Dk/uW
0ESQNpARmj3quBPoC/xo55/5HlBpdPRnjRsRkwyX4k5UCtFntV5XFXd3URVgwp8b
n0dPeb8Y6ZerB0L58pSo+wkawQT1bTrqakl91YBTCQbHahze55c9Ek/GqERI3cBF
ixLTkcczGh3M6Gc6A2EIxR5LbjhKh8crwLW+2GDMR2WohVna2kgNYBX/i6DX2+Tt
A5mFuWjTiExnfoyT8xptyzNHzBxOmKFpBkRVC9YUEtQxptWbPooWQkw2BnWWUdXT
8NQyI9g5Dzt19B8bgTKifOogunbdIh8spErtDpaG4MnOWwSKvDtNh4eSzQ0fa2uT
wCw+bJkqcRq5aQoN8BBKuARF0Ur2ogqq0Vha4Xu+z/qvhPRNuS2VZ0S28jyRiGyR
m1seyBpS3QlunEr1HWPYh7SHoYDMM52POQc1F1+UmLCNKU2ohPzpBU1tN9zOB/M7
p/S7YCEmEgrZf60Ti4EYGdfOkwb2hLI/1f+sZAZ5VM6y0rbLEVhHQNsK8UYt11XE
5IqzS5sjycqZ5Xk1mjeHiyhVjtsNdGnni8N2cHkaj3ilpJgovC6kkbDL66RctYvE
jw7eoLmYpQl/a9kJ09+GgLvMjwr2bZDaTH4SBqn8IPwaaY0aLXvuW2ZIonSoPwxG
aTSwK4a0CEIupP4buKBNxL8JZZdvttfSlEiHLzPR4K4hwlYqvP9AuVetbPks3QIX
CeeyRCOcJOUc92Z/NcqBNdsuiQcjunxZPCar0HowfMz+DoFKn1axKlZt0F/il4Co
mzQacUyr5vXHD153/Waw4rKwgRHxKWhj7JZH7d8pa26B7SI7FFn0aXokHWNPF82P
DISGF+nJfLp1IODv4gJgi680jE0KaLxpPB9MBU1i54LlkSEcDRyRdUTabjVo40bX
aFE+FGLWtYWKpQrR9Obk4tgpdeJItBjl40iKi/vF3WAcaO5B2OFRLfYLQU08jgTC
KGLY5rxLCSsXjicSHmajfmsrbckM/6FrXq9h7NKgmALuQLBEgqkTgr/Cil+aiqxr
2CnXckvSyTE2la7LqtqVE+vfUAefVneWWQOpIo05vIHAT2oVJr2hlf3L7mrhgK4g
rBENaxfNCQd6OObnKali7IDSN2dpKhU9/0Sc4V9U+bx8yj2r7ZthKntIL6tZ1iqH
SvUEiDc7xOOjiDlen08RQmk4gvMa5xLmESUjDFky19U8uV4T7jEehl45uhh/jWyI
NydKJJdT7/zCF4zbinmJ9YgFPIERpf1cKgLOK7Oi+tmUhoCdLYbTyhCeMFMPG4+Q
4qMiPCwVXe08/65TuTCTVgWwhedsZLTAe0qML+YdLKUfWVTJSldp+Hc0H2mhBq3H
dE8uT+X/C6gUfP17VbFHUFATPZagkFojLsIUzp0Bh3mnUZ+B7+SEK9fFpynTeioi
d/DjlJv0pcI8gLzhIZnCRkVPCIwq4W34NPMUgtcQ4Cu56Czm/gqaHEsa08BDDxae
Maz9JjGie2N7yse59Aw6xZURd1JVRjhxazaL9x3RlRu6meARzOgx69s2WXVim/os
eBvHwaXbLAMGCmiYIbDhjw4zPDbF7WYiJ0RDmkGmRiRshSMDva1wtgdfPd2+kj+2
zUoEWm3/a3arulD4UPPYNzswfXEXY3yfNvSXe53SdWoadlLCWHia+BAYp40DlZjX
PhzHelpjQQqBB7hz9z2o7CnPIla5/FBPMWc/daRU2meU/7JoZI/6e2EqmaCtzhSN
Op90C8ANqFsgET1rEfkd1ziSdCB1JLId1JaP/EEYheSukpmUPj9D1vUkDxQpEpjz
rzynbxzb2PXFDjf/JdR76tOns00LCXaSVjXrgGjuzt5qoLcsQ0UxwD+Ww+2b0F8C
vsSdbzAaG8byJ2GFVWkNwopyB5PjqnF2AxXJ9bsqLTzrYyAPBWMgebPb/IBxL/PP
3fw8mlZP55FU2Ne7jI/YGs8BnNGk/uzBNCrQUs4PdOcLFdbLW+my78UwEDANW+4q
v0KA9lqtGMvyx1UPdcrTRFEW3J4DSOuuQBZk+2ocLIYUTbYix3hBbxlkJrGS1hsn
RNn7C5pez4QCPBaAZ9kncs4FOpDd0gWlNeRuRFnZz77EdBW1sT7hU/zdOlKPEfYD
ArCfVc3ZJswbmGkYzq06/GX1RvUpDV6eff8n8Nc+Ik0M4WVkIzYTbz/wB26x3HEq
8oF4E4uFP3tlZYtgpOz1CjUhYUeanuA+m8yzEK8imXR1SLfr0jMLaDWh6r2xyAHw
9J+wsXEF/o0uBVLL9q/Jft4KQE/41WVWqpp71oytsWcLdOGI+U+cKIFeXNG/wB5q
5VIE/M2Go7Y0YDqbV6Wg/d3g1Wit9NjckSyqNoxqT32jxIdJrO5j0so3zYtHArk9
Qec0d8E2iypnbwzs+i31HqS2sXgVtN6Fgl7Uy/Ft5fckk/03UgKxCWYYOR41Aby4
/tddzRn8b9Gd4kOXeCIxBdy6hPbXebSHAE2GC5NE/MH03zNNoC8gHk2phaCi2kKE
9Gh1zkfOPQ7vnS84BU3/n7aH42eUJeRC6Crf/tHUM1Yuv1qjPQnvHKbWmMpk8aS8
dj1gWKqKpvdgqtqlgKrOCWWKO80TESKgOWfBcLnVw+J9om4XrUSy43jpsYLxFvc6
I61xQ2bn0Q0ZNAbrl2cK9hCUXgVz69Gzbp3+Vj2NG4fW6/qKCm9PNgItOK1IvRcv
DhYle5gKDz9pssFTiQ5QR8QuXm0YhKWmuM8kC5TEOF2ILkDt+QkpHWP6T+cdOGXr
JgH2trEBmU5SkOwM4J1V91KqGLHTMZfTAralLPkboXUCTMf5uEonoZWQi9ygQ9r9
f18CN6ZNRSK9BVBl2K8RwXj+5YxhhSWEDeYSsvp5qZrMrYsgaSb7hEJCfCb1vhk9
inhLMmRtqCzHseli9g6CNhjYbFKwC7OiKXIBnTHb0KMOJj8YtVBUm9Tmv9watPRw
2vaJb1Ax4cA4KTUyz0yWvc+XJcNNCZXId1XOwIX971p4W8A7NTt1efXQVaOlKU+f
Ef5kSAtx4jblE+fD7bqSpYExC40Nl2cLlMtX8tD9Ywam4ipsKveL7swa2gBN/mDO
MH86FMeY/EaJ4lw/hwj++aSJUWLNPz1yGE2fVMx7JLgy5+4h6VPlRmWy6JcPSkG1
MlkvkWpazbzVAgW4xJ/mJaZmwDg5lV4VOGIbNxc8JBeCNtK/IyvNd3VyMqChBj0e
Hz+CkyWklJV9HhIFSlXvunIyFSm19TIgbvR5vpf9fOU9RYw0wOnTP7tqhdKTt1xq
9e0AuKnW5L+oj13wyIPmIAOmgnPYQYBOvin25gnoIJ28X9qPLa9gYjmLK1l6Ue7S
7xzY8h9ogljKN9NUcYeYit4YPwzAWBi4M3YZbUrPMc5AJaqxmjLK3gHKuKY+og6V
WqM3fItQ+l+d1M4S0rCfzPJkRNDZd3We/Nt0a1cKAgihLSybsoAkNz1Z3XwjLpyz
bg+08vE+38XatErjCAyK7Hsi5ZLq6zSOyxyUVtOBoAhXtYG7h20IKZ/N1wUGAyoK
TKi08rOfeXC0Slu/LWmA/C31us0csEELxYKrh/EbF9nXYyGanUpa1tMPu/Uquqpo
s0VLDELWdzw6o47sAgDyfdOJJzn5fO1dV0/R6BZW3mQW9lG7Sc45LzSClMzlxAnc
zQvB+9c8G60Uq4CDWzAPn53YP8JUm6qtPAYS2NEW1tL+2XpuAAdi4Otipn6uP5HF
qOMHFnGtRTvrwXm19o+WvpT4uFQsXyfVjw7P+WP0Ce7PBIBNMQDhqyUO+lLE6llO
4GW3NPqhLyeD2rCGq7RWMzwba2z5Ie/i/SYbsfBaz6AfXDQ4dOreGItdGxLcjEXB
+t8PEFlInXmPdblhvmFkcimiW2oZM9mtc5VqQ1AGG1jtAd2jyLtAcBv2MUW3nnQd
N8O4lpHZCs9WCA+ORDdByqwH22lbwW9c87ykzDwE0boOF3gKcTuxet5KcNEu/32p
74cvOJaeWrv1f4fPPsdlJP8QlEZeD2P0OpzqfnQ0DCaOpPUZW/aOczkjoEhzaV/j
gsNxqFWdNhxuTlqdl0n/d7jUA3TR/+lf0IjFHwQFY1jwTttmDr3J5m+OeEC//ggz
uKbE7zyr83VWBKSOZXyDBiAprxrWAEDeo8emmcAUOQEfqxnwKKeED2v+jccKo+5m
gxRlb6yPvWpJgusXKZCsujrckgFgc8eSYblPirZhpxORlcr3wnXAHkxTdCSijNOz
syeVVqcGKIUkXmko/1A/cAT03Okmvjb7kS5at9O4dPDZnjZ34surpewNGiZOeXrj
ybkxquEql0S/lzPfOzhLol/BVwV2NKkLiFL1DlL6mYlGHKZK/Tay+/A9t1stQcWV
0ZazW0S5KogJETWOj2NQzj4OnWaqG55FcZUh1qBqTluXEPiuuQXFwcNmBOHZcYCE
6BS+y4Y9uRE3l0UfHXko5P3N8EzVGTD7lCbNU4/27vMNboXmbJmAoJ/fzLQnr6zB
GhIc+e+tbIYFxhjFstjUEfKVhsfEHviIpsRX7X4PmSGvsO3pTa8WQNSh+rlZYo3z
z0MXD68y5De+hfP+t5u5IcVY2z0yPWQpUPoe+VIJdZHRwaPukdADIAqTOPZQPZU1
axYnZYdSZfWT6fke5XHE1o5WAs3roZO6OQGu2aVAswcTD+sNHsw5nuRjkUiN+Ii3
Vgwv/vCQPBGz/B8bUK3MdNaCE1vxf4g6mjo/cOeA2KD3Y1hepvcqurN/E52zTmNT
gERIuvv9Y/fm5+5iDKk+Urx3dnbQltGFFRKxxxWnGNaGQJXN+x8y9bVJwWMSghNr
+PakzAzD4L84m4Tl8gzykc8TUzHjsyfTWAzfbyx1OoPJgPnc29RRCpmyc9DgH4W2
AFUTvbuW4MOXqNXc24Gbt2suqV8xZ3smQEhYGdlFpMN4GT5VIcVe7TKXFzFG0oAE
0/epYI4v76gCKEtv8WX2ZXGMCtnPWpfOcHk/2mHzLgcvq1NSiU4S3kVl72iGk8PH
FR+zkFnmKpyDafSvpeS4tilbayypcTUP+QrQauEm/wpU6nzcVOWtDiD5DnR1JxSf
BvpVSs8Y3KF07lon5BvZzEMpdldRTm84SPiyGcKjr+e3qd42FrGpXdbIkYOwvCac
vKoqVsxc9O+qWPrLHxc70wbN6f42bLSPISrWyaX8isDv22lE1UM4f4zJLtAzUDbL
5e5dPw1JGRLKlHSLaudKIt4tJhD9IHkbAIIuix2gR2im9tAsH7mAhZMsR3+hZMxG
1RxSfKXdwLXBAaaCPRXVwyZIOukwy4fVQfezHbC2Yt8TFekK77lMnxWNrAYdNsQq
pEGEfgheW6nOq9LAmyUdJsbHhzkbHElWEPjmcNKU1vM+0EDtDRXuBfOwKGtVz/Li
o84TeLZz8KYc6VVY2C+dHm30X6aieg229nNWZ80A9psUnHcWGwKK8ZEzl+lDjM1T
q7CEi+31Dv+07W6ux0oKHIhq/HxJZYUpk+f0AOCTbRJptDs2SKa971I46bKGRSUJ
sDHlDj8A8vAvFcdRk+/BSOw5v1b+EHiSp638a79C+ymuhyYU77pnx/023hXbyuda
ta80eqHk21fbCYqxbM57drmPag50WzlNWZi8J7AJYgfLqjezYAZ89fuMDUZIuZbi
udjViUhIpDofLpMLeYdRU7BDg9+5CsU4iU9/k5VpK2Q6ejwoza4Es55tbKP+qHJ7
9pmQXJHGsEyHx6WtdWh2odeo6s/QLuOEr7sKgqf5CENEaUcLotKo5vkkNdiJCmyO
Ifsey99IA54EpHujTS/1/mnA71m/XE2vrnCmfcGBfqzZDCD+LHOsVIcQsQUHCoyR
6wbrn604d1bfII+NZeU4RJDCxem8eGE7znsUWY+SOnyAV65/A7ItrZtOM3VAakzu
cultU7ts2FxII0is6CUv1QZywkeELQrGHQAOKsoLoKOBUJpkkuuOEKblW+qGlGPE
1HlMSlVWK9+ywSbugw+iX7TFdExIPj8UrJlGPyLM83B4C1lG/5Hf+QNFtdPXlbHj
tMzgzC3V1QzjmlMUe17H9r+9No1+AH3F1ISKMeZwjOHyrS7hMa8d2q9m2jzRzEZw
aFc+HUa4AESK/yBTm9xtHNQkzgBczNS8oGq511NfuKp+ufBeiUMLNEroYbJBhC1s
Xu2Dvl0AG7R8aBwKvEBGnatIim27jfJrSlyfuLAXRFSUIYxFID3nrmfJWLJpm0tV
GzZBsXAEaw/2TPsfRWD/3aRRly6DVOdEJPJL4sYlE9I144abMaVwfjnC0QGJA/HQ
ZG16F+WjHwC6NVn1mk4VVWE0PDqVdVBVCfZbPvSOxWFt+Rt9cgDb3TJFBv468KHn
izZXMmzxWwjoGVaKcPusem6uSwM9i39M/QkidEuhXDp6dH7FY69g4bFnQBk94/H9
soa2rhngHtmj6FNCdFeINg4wvL4/bgNK3vMqvb/Gu3cs9Q8F/bwfM8uQC54U3+YZ
PyfnVaVzuRy4LVncGsHxCycr1EvZWhcwHDgT5h4Ooyzex/6FqAJlFsKGC5HIL3YL
r88qJOiBORPeUNEZpqs7gRZ2wOxQuaINP9pGlGSPA3hVf0CMTi37c59XCE7pa+x6
5O0YxgndhfuUMvWE0VUHRMSw7VNefk/JeVn0IG4iWH3FiLV2nFn5h3DWdbB7Q2cq
2Qxt74ZSG3qQ7ojTbC4dMzGjsDbahVuOw2v87xOEgE1cjw24cFqlYDdnqtGA2QEy
mDQxoVEgpSNnvIy3o+7REso3BAi4VQBCf4RXzFK64+RcZrnWLhKvT8nMk+M0QG5A
lCEcoCC5v/qmPpJyDvbhKBDsq8sDW+W+6/+OizMwbiWHXzIhRIntOZY+P/7sLXkg
eitBFDf6r6XO1kXUIaGIJRa76+DfNIW2byyr5ife2JErShCPGZwu0Cwc7W5YZG9p
rAph2MQqGbPdxITyx6Wd8Owtt65IrzfveGaX8Ft4aKqdPVaolfs4siTmAv31Ivqx
qRnM//91mukq6VzNHl5J9mxUIYzYHQT/VsCoxP8Adl21+6pl7CumknZUZ7wDOXBZ
EGQl97OjSPvK0SR6aS5OS2L6bHo1IgDE8pexf2ixOlK1soUR69PzdXg18R7sU08f
c5vuoS0q/hWb8wqJUNprDBKyXHednOqftqhn5dNDueqRpxXCAZUOYFczUaoBhIva
XmZzePQs8HpvdlMJxznwkSZrfDvdhBYhkYy00du1C5ExwA0VMSEfw1IK+Ap2jZDv
iNzq5LSM1n+zfx5I9ojWfFKMioYaEjQeQxWUECYxfv5PjDSquLQjSaBpNeyvtiHb
ywwWI/6MjLYc/k7ibgdEHYe10keNam6tNjiRyg05VXVyTgGrGf6mQG7VDj+Bcbeg
Pkv13q7SfcP6fCpvP07xaPWXKXRBJWXlPvzA3z857fNr/lkX94oalB8rJNiXwpry
w/vJdvQ5mQ7QVaKHhozxn1LrGioQ/XiYbBROIIiXXCpsomoJHwuDqVIpmNq5yQQQ
LHdXAKN4QbgY2YWSehmqWxKbRlFIHAlnxpy+hEvQIpmu3QzNx1wvHMHjuR+B3W9n
xgMqtMqXC77wYJiPrD3S1qv8KarCv/bHUVZl7Z6D2cHRvSGF3WTvzzZOWr98BU+k
lSKbdxVFotAgy4OW9EEXQYLnb8dYcfayOSdC68OeUDv9xHzmKHGbYybeB8M7nMdi
pvnN9lSZ8S/fi2P+s0o18md4B7QSZIHmoL8BdvKEJaZzACaqhFZsfcot/0kSUpGI
C1wIdhHSSIfe5TdPpYqaavw7c+gWQgjZy8VWkDyYV1xGVJK58nkwFkMKYqZSoXgn
3ubMX8g4UVNI/pqW4Kcr1ivF3FOyBy2rVEsL3qNnStr9UgeZPKQhq+lDza7JUuLw
jUIMQxnblLBcb45AIbsZBPLIPkSkfGT0n3cBhBcBqOrCcGYXydKstGx9M7F3AhuM
Y4t1vpNZYxiTpOIDTokzrnH4VkbAfXxWwfL9lMbFhDO1CFp9YXrJzYIfdoy4R7c5
IMoNRW4x9MsIL8aMmxq81w8/LPZg4L5/VUbHhpo3NLWSpP035CiTd+UCVXDeqabT
80xrUs0e8cqyVOqMURnvOFwtsaxtVWEFrWgPFXfKfa61uZi/hHxPP0UEmCVjqOMU
tLzif7Kj21iv+9fKy9w5TeHZ3mCfZaPbQ+Gk21hsK53kTe214wPgpnHjX99OecYA
SwZsHzWLD+zr15lY9E62JX3MkHInts1L32loCN9QaJDr0Auf+tnGWB2v43t3M7hm
YVvYP7dIcZ3MAF9J9xe2Zc+luJ3eklpXd9i/1u2w83B10T1xhruX82aXPcySansv
fiEKi8M5ekUrtK108O+e+zsYiil85lmo+l8WFJdrobcZqdzb5w82N9SQkioKSBmh
p1hW6jZF/hjoRJ50u0vp1snZnAtf3miANSiu4qeVTynsRes848tYfUASS75/CNnM
Za83n1ls2J4UTmnx1ETTgffbKKyck0msYj9TuJ46JT652OknHsDzJHm3dzTwaMdu
2l7Tue7ikjTlYhVfZPrxzWVhKVNZfybQRSlCFSNOg4GJOS0YwexgP+llBCelA5xV
GCyF+mEtL+7PIK91nhtqEo4eFHzK/vVblbCbZaUOhW5HlhwFTC0fSECLj+pjlgeM
Gg41OJkX4JIxI5fh8eG8S3Y+QMppRak6tr+IBszUl7bF2NIBSKXKY4cR39nSPVvd
d14/ex147Z2nqeI2A3enOS3GgCpwLc4Py0QdAcJ6LAyVbv2ej7lGWkJKPOjFWuY8
OOMmNEa/RHFgsIzNZT8zqyC/Ong6EjBnlEcy0o0LO/JLzmn5vOOm110VCXYLpisZ
AFOSzWqVHUCEOQWcBQw9NxPft2IVwPCvDpjeU3JTka2U9NJ8+x0bgxGqQ8eFga1N
wNWzGa13UNpH1H/DyDSSmBjRtJ26so0CQfZsmHtvpY91SkaLGCL6Q7i+ut6k/xCt
6K+3Xd0YiT/AVALRh1d7LoiORYatpfGQVCQ17AzsUfx9KtEHO1f3Dalw0PjnN6TJ
66Dlir1gjEnwVEUZLKz1LFVixAqCpT2GS691Ilgv3HSgKBcbLnS5BRfQ/8e3GWGt
p02EuRdlyUsZACsY6r53FEflKKdsYnzZmY2wb0mDmtfHEkvdOtpCMlJe6yS+3NRV
t69HwqrKkIV1u+or4/nAdx9xEzhuFERmd5jQXM6spo8ggIEPwdmChF+KqjOcVRKf
cvANcRptVFwj8tW5MHlsL+IDd6B6xr8uYlc1Pyuayl3r1K2rgu7TXwc5bL0Fdhxp
8Cy/nuEt7ToSzkjz26CQB+HQCbjx7UQVkBTWORdm9rPYBAprfp2UJ0c9Gex/iWp6
MXkDRHNm3nka/N8CCz8KRH4zmvoYmLEKPzvOjMqOXbv6JvkPjXAG5iBbj5wnNKP2
ld0KkjoQsNct2Y4R3kFlKW+ZPXNrv6IhyX2f9SpnxQkzIwPE6MmKHxRw6fPZbkAh
rnHBekItUg7Ak8DM8k70L/FyWiuZa9Mq5V9+GnQw8H+i6HxgGRk0usBToe5rQk1n
bFcCrKjDFtfqSFpuAbrB7+XXkf2mUzW1TnqOhyoeAJ9agm7tlyosFOXvplm5ChAg
RbpcuGjTgDD7uehHZupJpHE+JsvLT8CBrNkDtv8AH1zEBQjh4QwpqzjOx/Eu1hLg
sfQiEcG55uJHPF5S58XYPq6xB1qf8VMfUOPEgoI2QAghklQ4AW/txOKHjON2GJwK
EAQpEp/VGff22pBuvPxnbomFqXmishCyDvPRbyi4E5C8x2f+AbrshG4h/w0Tfuoj
rjv723egk07eDH2WK44OFANTRROCEUpi2eYWxFo2t/LKsfLtUj4apNEt7LCqMdbw
c98xiZYmPtBkU+WeZEV7osoyfxmic/sC/pREDpZWr7jRU6d++MDf5ujNb2A0rkYo
tHkJP7gbWby6Xx45zm0SOpZbHQObq94j7z3OzwDKIPaTh5SunOMGSXwRvaQesnR/
CzjSsmpY48KmuGr+9aLLi6dP0BlI2BtInR9z1cN5At8OnySP61gVsvyUjDOJNzW1
NHQnE57wMTXY8yL1l5fwjLFSSRgSP5Rq6EbLNPICuMjytt9lgQbs/yGRiE6rZ/Ni
YqwScQYIfHkPjfUHf8gpluPz4Ea1tp3zDhBdEjduwAymFEKXt4r99UndQIPVv0BT
BVg0504RFJ0FIrKR2/tQaRNH/n9RCUjNQV6TboKbNTiG5EJ6OS/2xf+iDiVcM3+Y
85dV82NccIzXU2iiv3eeFPvc71piW8C0Rpm1fwVjx4CGBjyS0Jz6K4Mx89jXb1Vz
lexMLT1zFlKpNd5YiViRGR/sjpITzmHiu/9UXlCgn4+ouVqQymW9nPITxEncWm1u
+pXQ5FuphoeVpmpQRqn7FJeHIObashYSGAH3u+HPRyspbZnr1CIbgC1/9cLCJ2x2
B6mB8PfP4BUTHXU8dVQ+wUBzPrpb3NQadaviwsUpoMWTQ6jkXyU7xvgMpAZAQBBZ
nzJQVFNi9njYqJQ6w1Aq6zcCXke9lfNeYeMUiGFXPdaLjg5gqQvDetukxahjKi1e
6KOsgsXsiKhwrl+FFtD1616IbEx6cZofVHeEOe8psA5Qmw7wNwqwnihZrBMPnrpZ
/leG+KPPT4nlaGWPJre4/DjmtY3bjKW0sLLLSyGSjIBmtmVssDGAjsqo0dRbLlmq
cctmgtRQfMhGkOyGkLPtUSldIAxmodmT2FPoz9Nf3jsYFtmcG9nqamYaMe2p1SOD
DSKftr8qgITu3gWK0eVYxdOcjcTCEwP6q0Ns1kHpEqOOYyuV0CLPRMm/nbq3xFN7
z8rV2ZLk/8Rk9lVzI9cizVNnpUhpa0QZaecs1uluODz/U/KznX/gFoE6WIgSFPMA
r8AL/s7AS/Bq/Yw/UmdcKQyMMsnMUG/Uj1sMjKrR9l8yb6L0f3BIwrvIIAXfFbXr
GDXnP8mz1NJV9uOabfHNeCymBYzbysgklzz0LGKu5BBxUJ0nRNKNc3PyE/i4v4lV
Tv6GoHEYg5igxBE8g9Sa8yuWpsyfGJ/LW3hshdd1fQ3lbXu5wnakHP3HyEYFpSCp
YnAGcSmOZc1iHn292EXuCG8PVxR+3MvVtQBaEJStKfj+FEJ3o5whYbYCDmlL8MtI
qu7bwU7hicZfafR/wtFycySkOQMfz+iu5ZPqpiheAe2FaK7VkcFxhccGXZaUH+PZ
xJ0SBvLb/b9vdfGA2Ipgrkzc4oRt6KoQ33+l+aU1BHYXBUsvSVM9Ldp9YdAEaArV
hNIlT/U7sc56sdzRKmBAl2Er4euYk47moAOnXo4U+edXVyvZn7hwjipFpr/IL3PZ
VJd05nUX0tR6A8VYFoXSBbcR6K3WrPUdX//hqoucEywNBYPW+40yejV4b1BKZK9n
TvPQf3y/9ZxU6Fd4Z7zXDwHfUbKXtc9uGHG1mGbO96m7/D2wJHL2Rmn87c9X1k40
ylsT7TruEHfKzLlbZY/56mv9tWJuTAp5A4mVSDUgb1LSGyLlMW79DkvGekLFB+bz
/NpsqWBHc0Ej776HDbJvZr1GEdfzy0qJ/jYzq1Qex5GBmSXpIxfTfeenisye+wrP
BZMCtUKZvUs1TzDyUXS3aR3JOc2zjDKgBwjgiiXHXI+f6NlhX0DzZDjHDdzTPp9M
3q6I7kt/fGtqNYGDpcnPdz6ZXRZCnWXIFrzQgPM6TkIbN2X7MPXr00xF2j9JAiHU
P8HfV4eRREdRdRNZR29nMU/2P6RuoxWEAwk0b3uNPmLJuwMNveQSQpc/Zug0LQ8c
NoyS45o4s2zJqXUOEechKdZX2n52AIHpNTRIbIuq96ILm3JeYbG9Tl1XbKHST2EA
Yg/rZf2OaudYek71xzHwDVlAqQVtqBg14Ot1zxdjcE8AoO00VHjiMAEJbbJk7aoH
VGw1FeJKt+xq0+8qBAAYzD687E0tXE55efRzP4NTMbQ0UUrWuG6TONFPe9FcbuHZ
h+q+jecXgGSIPzyACM5NPLDrEnFwCcoW1kFVkyYNz0YE7rQFPEZr7qOAJFlKcqRw
LWVjcxcE5X82bwLdfgtQCChVWwTjPXp8dIOVGHWbGjM/tyC1LN0nw6eifSZl/rmY
xu6mTE8Jzary4kbY9BiLpat288Al3CPUokYXcNsCIl9EdVRWqJWZtyBsQSqaswDu
mLA269n6UoR8Q7n+O7KNCxhktJELBsF+tgWcrLyAySf/PZsuYjkLzY4QJykTII3w
p9R4QggNSC3MpudY0EFTABt2m4xU5pqYwAlWaOy4neO5wkr5PNlX7AEr411ebfz6
HdHswnzcTPp9CjRHh7Kq4FDdijaivYmtgQWwIpqH7igUx2SQ7ajG9U+CPRUCr5r3
wZu+6nUpM6edNCFUQyNeDgUXAer4HekKQU1Vu8VHoB/50kkjPfbIvRJ620QcGH7Z
ClfSERa8gvXQvS1htn81ms5r2bhk86GdsMQOuJBACKj+tndWnwtAcaWyYZAWQ/vg
rB5cwD6ajeVkvqdKREWby7rpZXbhSksd6Ad/MMZ1eX3E3fGuCaNFy2bnqjQkt6qN
JjEOtvZ57P2MSgKXcRYmDW01eBeO9FDcf/sWZjGmNK6xUOQuwOL2O2WGO5PsG3+x
YpVja1u4q5FK4saiifIIp6fFux5a7RYnDvIEXMB/sioaob7k6jp8Fpq+CAXjoRFH
YbLpJhPuNMOUsMVkOt/gnM+QrVMFHHXpWUzGpp3Pu9KgEyBS9R6L/ZRB32NOToVA
fTtDHF3nxVIFpgN3ascMdOigf3AHPOwIJe5FTvJkIQ/cOl3VKXKIUOY0jt3EAw/p
qcdDZ4Vnn35D6RT2eqdy6L67M+QSHZfeQr2ddP0RWp4SlZjuWtYmrGCDMUnmgYqk
QA2cMO7luUy4dpy34a7yh0jhBMoMsKcsAJVzvOoMAB0wpjRrbWT2tNfI7c+2ZMyq
d2kGbKEChzlAjU2C18NeS19Ha0+FUEDW8HGKXwBh3rAm4dUM5YHUO0UjoE0UtITe
5G5DsU9I+Q/ZIOJWCfKZdrJmn8uyrAdNSRjU/sjiz5tK9/XXifOvZFLAMZ9dKZYm
q1suoIF14J92SlpOI4naEkEO9O6IzkFfHrE4NVLtRLNr1iC/Sky5u5b3hC4PJCVC
hOcljJmuf1h2I3y7o+rqJC5EnkkE5MPH1BGfjbSQRH9a0zIwb3AmazcRpPDgJi8z
XLkAOkCiWaxmgL5u53qVTGuMM70yb5xsixh0XRePGNlaBfGvCSszi9ilq/X3tcic
yKx5cu+/J4FMTdilvsyzigOU69j5hVCwicvuhovGpEnFg5agRv0BHqSAwRT8X8jq
bSlr8YJVxZ+UTQ8YTVqvWlT4QT8hyl3OUHXzZlUQn5RUjIwTaZJKAPiHwChXlP3q
Q054wCFC98UHhylW4ZL9CujPbxnN7MUTBOwJKCVb5Qv+lIY1UhNzRRg0oUJ/jF34
7WXgDYWyiADDfOtz86zc+G+Ot0CepHk4lJZLe2aDaWDdBLR1ltxjyaYbc0nGstYG
8PH9omfihskfkruuoC9iuAgvKk62slP46Tpl6FODCQPVIIz0kH2yJNi3+/vqNMUV
bOh+c5xhX3Suy0oDp8n+RXaoXOBJv05suEPjzJ6rKAKaZx3r5lfLHD1Y8G1dtWdE
8zTNMYc6y3CNqkcItK8YoW7zXMoQ4NsJqXrxmhey0wRL981Pn0mhKLJNCx+tmHS4
qowOix1M8qpICufDUnfthDVHkgsHcZ1mrRi8h7DksZOW+E7OSaM5LT0a1dwxqHIa
Hd1HXPpvgjWQsTM9F6gh9L8P7Q1EKcUzgqvdC2G8iiUwowqQsWYZ4u7PLxGWC7gZ
l5tIu5UTIl5hsCTuezavmN0mXi5dLcVutUpyE1z1z8t1uETYZLRoepiLNebHnbXM
EhP7EgeQjjudpHxbpVkderwyYWYX2hOvBcd9wVfG5jsCYyQ+/Pl07rzEUjdMLzE1
a3q0lhSoIgV2mNwC7yTE4nPVZbGh0wS7stf0X18eCFSYcINxgCRXo1yebn0mEjL2
xgarmomvDFujdfx6fInPkuYX2+PseyCAWcTtPU+i64A=
`protect END_PROTECTED
