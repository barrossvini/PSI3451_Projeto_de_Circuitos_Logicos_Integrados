`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BPwfXq3p1byci/mm36wDn2hnlV+otvPIoTP225TykF2Ohz2UQ9if9iupR6EfWe5r
zf1drMq2XP6CGD5zHUrSXAHPBIDv6xWJGLJB3674guVgFKSAw6KZHo0LV6rOWcel
XUdWbey8VPcp/8tQlceVvOCQ++luInSGARf3ou9BkPIzp2cdcMwsvBumeaIlFu/W
i5nl6BsEN8Im+8KkMgm1huZqfxpGKvJYNoAW6gD0G0RDg6AXBOmo5STQHMiM8xzP
/769Avt//i4Mt26j4XBUU1Un8Go9Hh+OVopzaKRgVOYJ07zzWaVpZEJ4Tp5oWBXV
iVNYe2koQ8XokiJB/A48pVcSDtcI1SJreXiEgIw2vMknmyQ2AjYRujO3EDbiXRZ6
ImIFzo1S803Wkob7/z5qdesljuamgZQTk9Rtu2gVV2Gh4Yp9a8GW5fV0kq4QsY/i
VFQVLuNfgxM1lZ7tbwT/KwmipZIAlKlm3Zth67C24SSpiB6E2nTnX0vG3hOiBGKC
XeF0trTN5x9RVW++UPGUY2L1l+b9JSdBx1uwRkSIWhmVZ7wuHlk8oOrDSEwHkwBm
sYfCOV6T5w876F6ELgL0tVHU7Ua7j//QAqb5X6bI54Nxxptnmd7n6u/2XL3hxVW3
NUH5QqM2SKq+QQA5ALAuH2Z4N8qTJ8ufTZVxzvzSb3pzOZy18LqwkiQI/WJiwBRh
YnhjY153Twz1V5gBm7+AxkbnSYcwChj0lcYmSUJnhgr2gqsvic8p+1eoYuDKwLn8
nVepMDUih+0+7jzL9ReyB5kMqf1QD+vhUQY1m6yrEYdDkxNQC/Itng/zsB2POued
Z0eynvy92FonQ3sQul0oWwz4X0WliqrbcvR5lbgMUEh8dG19l+y/seF/ZRViRl8p
iixLEeSK1k83Y/N1zmZsyJ6rL3hMRkJ+jYYveUpdKfV6wn+duCdY9buKoqEi2phS
sHGEGOesZLaKyRG8Z1calTznPfaDGZkcClCnMUBS5N+RTlgPlTUvoKyjy0sy7M/w
79U9zYtcwqew0zAeolICo/V9qZvP2+0onStfVPv09J5quwdFKHbmPVizZyXZNZ0C
aHRI2lGrT+qSMbYCTpNGzXviyC8pWNbvziKM1TjXZae/4Je+Oc0XrkeAqo8CB/m3
9n67fYlZHDYdxXRVAEw7Nu9/0wRiQGkLDlSE8+qzIZ5zZI5mr9tsRofIkjTa76AJ
vWwQrqzcCgGo+Dobpeo+5uJPpEx1PR3T+WivONZEgH5EGxNyEfKqtWRiZQL60+oi
6Ws+fPRndZvc5ccwONs8D3HoBpeMHcy7aHSoX9Aao/qNz2H0WADrg/NittYvufg+
GH1E634Gbd90e0sb8qMK6UGLmQLtUgqvcFBzCNvnU6YeA8mX4prVhrXQmjhYAf9X
mHwdB6K1sir+XV41F2LJnsteFaaFN03YFolxDkiZuDh57tAhvzUASrUfABjhJBNh
y6bYryRsH0E5NqpealijHUL0sRh5UXqYH5rrBbDhoPD1n0q3v1vcoLChM+FNGEhk
74UHjNUCPOxiniwAnClN/c8Po4c/ebsmsqgUqGC5KAow0iTVBUwv+daaZHHs0Fw+
NVhWsCYm6XAdohtdgEA2WgL2Qpopzf87yI4iMpIQABnXw0PX2A/V921sDRaeyC4Q
Lk/r5nEncMDtWHsDHYsSy3TKW+qaTQ2RcqgyoIR50HS/X6TEr1JvMnfOdE/zyXie
FZx1m0a4V608PV5XbhEvVSlLwtrlHe37f/afMu+Fe2X2MnJbGXkZJQIhPpAXgze2
`protect END_PROTECTED
