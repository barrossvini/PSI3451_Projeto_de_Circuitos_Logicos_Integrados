`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chBDlYmTfkAuC7+WXCv6pV4tEO8ecyaKHKnJMckuQ5gt6hPJEO4byqNpzYejbNtH
DTKGhPEHOUWIjDqX8HYUN7s1S9M+32hh5dGCUqB54GOaR6TVBQWXZGiuxsVi8QEz
W6WoBTRK40E/PvRaRcy85F3+lm9cukuZPoHYRMJNDhmnH9O1FQobi/ZU4RC7msz+
K9G5U0lMXkDJ4jyTQjs5PL6AsLpA33WYvsqx/gAYNKqiMnXz8OEew9YAMl4Y1xZ6
7PMsNL0ckDOt1Knh2SOJ5kRJzh0H3Tlpi1So7GvjNKL9Q1gGjA+HRtkj0haPe4lk
gmmafYW9tbYR2D++y2JXcX1gJGBCfR26sn/gGLWRuCCUAOygapGsyKs316S7MJ2P
+0rDVzuRtW9plde7OSyLBE9r2bDOoJj+uyet8KVlY2XcdwttZeYyec2Sm4iY7EEe
eE7bJI1j5jg96LhmF3KhhsHoJ1PTRZQ87Th4a3jwO7nYeMS/zwTXAFDBwmn6WYCq
Scr6Gpju7CCO+vf7Se+BbV3c/myIT/3xEXcK4BrxM1EbMLfrdqlLedT5enm6PsBi
TptPu6QK8bQdp1/omwmueIhyhHHj6feXe3l9SIPue22XWBFg/cDlBVrTTSWrHPpz
ddskBAtKDuCLFDouL9dM22/hBdj2R7KFNOo8AGFLCynIMVlDFnGRORsanqFA/tzO
JyvFFdMdeP2BuzTL0+O/0F2zL2HgmFv7RYGY0soFQVVyuJECbqMyxCVvN779pssl
M5i73d/Bo6Nn/h6kzmpwvqtdHjZ5W2U2gzcbhE/bcFxCTEq2HiQMHkW0NJo+7tnE
uAS15vrfGWPNxCZcfxpYqv6LLsj5tB4C8FJk3aZOSprCezo5Ah+31+qHb3deEQd4
P2MW+QlaTuB1yC0s1qxuLwPG3VsyxyeuGz9P+oJgEXh/44N882nPZ/g2F6tmooru
Ixon4wo/wvAa8/wJYIItm0bMCg5EfAvesc0wTXtFdXbvqDT6eUEBBmfN1bu/bfU5
u8GucAwweOIgMH4+k8ZF4hdYYOR84N2zDI4dMbgqCXfgrwF2VzxHhevImmcciEuT
Ni1VcUOHQXgvrmApyTa4UHA6zsA7oM1nbrm4PuIZ2ccu4I206ayB83KxQBFUPAfr
7Axqk46QNSDqWA8UkN9NORShUh27YP7VynhIKiAlhdyI/DuMKwoZaU/1Pnc8OiIN
esfXrpxhqULpWw9WVtvcuD7UKpwUIiyesZ/1vjITYzeV55thNgE7khfPVGC/UF6V
Hyg1m6DS9xYa2GgNrvGLLIW9xOgYeIRRzPom9hGNhLWY+zj/67u2RBCkG3eYykyX
3i5LNEv3zGz8HkbLQy8jWvs0iiHcJRhsftEr08k4iX5qtFl/6mEevnGxpJ5D9LOz
F4Skl0sYr3hVl3Lv3X017yI5Y01bG3tq9n46vCTuPnyq6S4hn4L7UwcnxAsRAJAi
f+S3givk50FX8BWQ/QVHzMybYm36Ax50KVnhzb9VVs6jXiK93N+2Vi7YormIbeMi
uOQE4KHJj9YCbhbyxxByDUdlDtgvMYFVhb3S1pJijz5OQPMgSdMPkDZSa7h9yZR2
IZc6xV2SBvQNeguXTwXqJTKKmb8RFEDZqO3Gc0EJIHXCFH5ryp/kXmRpMSnHMXZZ
a5cwvBSJGJIqQvTGu9XpTcOZVJs5qG2G2uE7mzZ4kv8VuI1VC+FovWiBufQ826OB
yT6ftU3DcMLrYXUTvE3K+Kx4h0zklgFpodPW4psxdDswgDNudVXLvZNeUfHefL5o
LC7RgO6HOp8BXglYQc/Ryn5ZGpY0lnLOrlBOr4ibsLpnAm9A/iLZsLaYyYIR8obc
xVU6nOF9ylvmAHkThDFVyQ7IuP9MhfV3rx4OEK0M4gVRlNdXKwKQic/IM7YBdby1
4uf+kei2lFdge3FZC/zGamQOsx71IkLxCIgElt46INpLA44o1y/gK1/013arpAiP
W+z3JE7V5SyyCcJaTfzjhPPqrerkv3szncVAk2slOoW0/1+H/o84EJBMVR97D1Kk
bHcQNpFMBpfzt909OCz/f0cABqZ9YUJGf3Y6f91C4Zjzb+kYT3sLIe8y1GDux1QQ
Tfk7OyympxodW2Svq7B3z3/+hCu8QKvj1sytaDwuRKGQyE7Q0twha5Gy3a5KjRUo
9DSqYzELEq7Viy+PFGAgcfY7MkDx39ZR84lEvze3w04bIO9BKV1WVBNdOp9H2xF0
4HJWOBKd912eydHPZfGzIXyEvQTOtOjvPXKhSZ9sQh6dDfr5ENGsqAr3YYYVzelR
dabXuO7VhBZFKyaUbkbNXjIcI/I8b+hsjonOTZYxWgI03KyD2Fp9iwwVglRa7/tE
4NnU1XkyMEyASeUXMi6tyblLOwyeot2U3xU9PxTWN+r55UgxcUtJtR/Bd4fwg1NC
kuNgrcxZ3C+XIEs2tzxx7l2rONK0PTe4VGQvxe4w9qw/ahkXlQmbNKEmO88YDzPO
R9NNYQCTv4zY+4RbfTvMQlRsh7BXOFXeWAqsavR3vi+l52Mi/VJw/ksOaHcedKjP
QHHKIJQLsIJlo4Ss4W1AJnoISHLIdkGlWYamg63k+zRfhIBDu8upvH3NUiM+dCMo
i9zGmg/feViKwJBrF6UDc0g2giSjXofkLWRwZ/yf2DYZs2WJbiBwmpLhrBZYH55T
TXb9l9NRLIf5cdZwsdIZXC84p7kfqbQ/xQLC7nMeVA71Mv+IkRuq7/xmH/ZBp6T8
1d18wmh1EMN+DjU47TnbWhqg92wH0oMVHgjuQEXU3FzjXIGlgXQv/KR44iMdNjjo
bnez/CLWUfbtQy1oVKPuWbpUNEIhYImyuGquQImnV4RVqlsN+l2E5bHO+j78rYtt
C17XFrqtIrVNIql6G4sQ+np8cEG7iyYnzLuJUKHki1bBUOCN/VGGbR5C1BkW9C5s
HwbLoRZA93RAOx7bKiutLcCECMCMOUhtgR+cBnuPzxEvcgLDFOBmSH+hNA4Cg/12
zyXL5YmE8sZkL15ZkXWtu8kq4VSD+sry7NvTCTuiB/tNXmw65xUfalJrNFHoTd0r
/xdZIolaLm2CCx01MSm87q71cV4c3NtXsMI5rvl9FZ48H4zs3oIh9Y+nVS6jdHzI
5xtHM57Ya3lGkP7WRZ/Flp1wIj2U0VSMlve/OVIVMiFya2F4W5J/CASC+xn/jpTW
jz/fmv75RR9Wk+xpQZ65FPqWoN4snmLy4L0+IshB+wwreZAHiFmZPA+TEt7G4xFY
4jSKTi/chum9p5/VFlP2vc7FXaau7LkBAactZoG13QIt8+9Jupdz7omA6yx1qhbf
gudiQQdtIfl1VdMif4dyCLasCJmbVIBzKkwwgarFtexJm4vLTtMOUFl5GL4offE2
ISQ25xWVa4gyeQVR7Wa6pQO4uWUY/zMNpyUWvEpP/SU+4iHBhMVTa0808rqrS1Jf
lp1zHvp4Mm2XpFdCj8jiV1Iyvl2f+x2W5u24Ff0UVHKU/LV/6n4Dajd+ezhFAmN5
evDciXQcBZXLJbNcNq3VRrlYc1kbO8qG56hOS8cgWiYLt1OWTu6pHdIY/vHu0pjc
RuereQWrffetlU8gx7rOMHprQv3xM0EFSiKfVRFOWJHfzDU13hU1BDsAxmzLq30O
FpyqJQTq163OjWuZONBS8Thmqp842rx1U3R58bGyJysbQbIZ3aRFuwHTrtuS/ueI
jFcquYdMFBflnZPUufYx2dDstchAWY/HDezoVxfEGh9ztDTZItLRJTV8A9aMBUS/
fUDzCI5RbZA3W4gqGuhxMEfwrYWhthTADTBpBLtyQpJSUNcF9xI13qNgJ+xMxzxt
VSeWZMxLipIWwM5quVOQyZ3IXktjVjlLlio/vlDE9FjtFNjRDttKdT+pyNs81naz
MHVRnISVZT2qyLbtooAGiHarG9qnVTsFGFAfIQJrk1yl5Z8z4XNq4J4cl5J6/88i
2g5efdr8xkZhNzKAGz2TCZsMFL1zSur+4bo2J60LYqiuPFd+thet7EDCPRI8nVzO
9RSOIyyMLZo7Ufo86eyAbGTM4XyleMtP2kF+TjN1KKFEhkzupzswFXrGccE7P6NX
XuGwpRS2VcHYd3icvZhdGy0xjKi0kHAqkswW45H61CLlD1hxtIZHQSCEeT7fHXUa
s4/ZLc9aiDjZx0nMe2tkb0qbiHnrkK01Irg8Ga7bBrBVYQS6kKMV9xW23+hUntBg
G9tfNW+O4ZNvoov9uLLpOHH68u6h9G1/K6CRAPzYJmGdIzLneoUkDORep7UQFhGE
LZ/rM+CY1sIQpUT6Y6+VQnPSpGQNuj0IpJQ6gN9XEBc1qcBODJbezvzcb7OX7Kr0
c/TBpsgl3vU6dcDCmoQOLawPyUPy7gYeDHKGzJCbrBQqFT30RI4bPApIQH5k7nyL
OeZnFolRjGJKKeJUg5O5BPp6TWot2Zc5gW97+RhKPtv22j65/nMrKhzEPBvL8yEn
wku13DbPfk42gkSSKVCGe8Uq9DHMKDJOo9J6vg0H4LxEDJkh7InNwyw5UBD7HH/a
BgY34IoWLN+hZKdYN7casl/QvTVmAixFXGawlkDQ9bmvxDp4Gz9sNxQG/hEapHgE
f7eDLHyYo2Y0m5O2Pgdi7OJ/xt9JItPUstLGv5NJ5rpvmEWdWAKT5Va8co10yjjm
23j4nrPa75YnX88t5dc++5kWTadjYFzc1DuBiXNDeg2jOWIq1P+jgotqAOhgmfWS
zprmgXlIoD95QV8zQmEMaVPOzQSUwRqA1mbSSzwfpvekylYkrhWaD0B8F3uL4H68
vHnthMh3zBHbfxE7OrfFmWtABT1cwoI5P4VsfBCqENuTHG70IAfNOmWG181dYQkh
C76BC1SbFyX63RzpkUEic7bSm8DrUBbkGteeCWqOXt/+IPpFI8Zl1oMfrkV5zx1S
HM/w6C8UaEa9HAgiUWhSsx9mA7oEZygqX1X3+wBy1Vlm5HrTX3ar6Ql5XGopEJik
RPfnru5mE+pJoxm1YDKnzyYQzt9nPbf9bbhaMMfP3Jpw741ZQdWa1a/lrJ1cRmPy
24rrrGuTqFRonquMI3E3KDYVU8QxnpbAmRbBkCgS+Vq/ewPipt+YB3IUutI0XWFX
YECj9aihFk9nGydGaGRmtixF5bgrDd99wp5FGsAHqUW0Z9D/qrDXVvP4A/zn+2FX
xPB0crQFXFppiKhipuwDI+oxrppMK7UASRGxFDBnVcziH+MWqy8+bB4vINeSleIf
pEjfF2NOloeIox8lz5XBGbWA8OkYIySbU1vnoW0W0rzjwY4L8ME5azi7QYsSWVle
jko3wpx3AFi67cQ037nESj5t28Ttd8fRy1c23IileWifnjy308oFEZwukE1JICIk
dfDISEUAqWG7aEcVmPImeun4JWKhF4JjG+sMjmX4mayucBd84M66an4wqx9jWvas
IotbESCbaa2izmTXG04DwdN9+VvepCkMf8zkac1rZpdglA6f6ELR9kpteCcsP572
Sj0P7JHixP1mHI8d9RcTf9xcIrKr9NaboQ85m3jDENky9cnfch20YvQfdaZxQVUB
6pN32Q6n75PEFttf0kV+87v4XZju9lQ7QdZZS8Mk3Oqb6HskRxEi8HCqO1YSsAXp
+5sKq/iIyiRg9/+vVkY2/MjT+/081PFFToyVRSSS+X+c7X+pUb8BPp6Runql2utn
RUmKqvILSl0BMx44n38BYq+oOBcnHXMdQ6T9Ct6XDn1jWmBybbUtLjh4BAGZDvFd
jwS99O+iEXC02ZGqPaj2LTx4CpkvZ8Ajq5JAxKLNOfSdK1a/0RC2VrDLHloIeGPy
HL6GEQlN+f1C/XBMFU1rxZsR3m+PSyAJQfPv+xiM+nFulACpp1XNphfL0iFtTK1v
fZZfZLsNeeIARC1sZIFpfxkqQpSalBYERFk4LLoy0MeUG9Psd7HIOCUDRxJOfXI7
+RhtbUi8dHh6cRVxkzWxmq+GOx8R/BwpEzb1T6j0ilLJTvC3nEgp1phTiuTYIny7
tvFSuB35TcQI0bXJZl+H2U+r8MQBQzfsDRA9KxcjSw3c9Vyze2MxBIzHUb7puLLM
9YzxmEZ0pKWrvywvLFbpdGatlPBzoikjEODdSFnbvEE1Yp1s3MPcNZrvOCXRKxM3
LI78/mn4lAi3YS/ryr7QjQ==
`protect END_PROTECTED
