`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P8IR2UKNRJmhsrIHTvuKMCi97sutXra48mFl9tUeTBZs6TBjeMJtouhmmWYjNO9S
/SEfEM92yV4Bb/cti/ddS0/UAeuVJ/QE+xB4hZ4V2VKeA9RSy8N3lIZ9GC5yzuy1
mBe4NFMF7ZmegmY2hWyKzg++AZZs+anzM5IemQ8ycoBemRTI6hBzkBdJnUgki/X1
wNb1S9WWNTS0tTkVkMvDKtGNd4fBwF9ZNA9q8wZzxhX/L0JV9X9qV5slvqSwscCN
FFH79ry82++ADLoYJFrnpwFT0313UtBG2n7tCaCKF6r9BGMltKb207/sBvebgff9
8meOH/+WXJv5JzyfELUgGPcHCQ5A5DohjgNOHCYntJ2iFilxFzxfBTqflw0aLxNe
euONc73lLMmJMCi6WP/i9QF/nS3BtFC11H1HMr41yEt+8bv1UQeO45Zt18lL6czK
5XazS0tFSfkLgcZy2J9UFILlypdbmOQD152PpQKeJSvH5drpx5XC3dI+RCjV17Ky
5j3lEZgoQXfIsLj7jkvrODakwrBb8oFTunyW+WP9GvNfiau18tHEmcuVIsLF9/w+
BatSlyN9Pxi8AKfrpAllKgarSScV7P750bZJWeuHDDiOHPDoqoiZUJYTMWchuSB2
Vyh3zHrHrm3an80mXqPeeQd1uO/yAmH+DNE16abFl6VMfAmQnt5Iovfq6dxaPzjZ
9spfTDrz9S3JzCEX32nGMYvreit3FYrDoL8WcuTW7ts=
`protect END_PROTECTED
