`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ch/arZ8Di5b8y8kSEmv6DkpSpjmOpeS/1+aKUBB0WHjtpazr6hylzgYb5lxpj1LA
6NUWLyQPERUNFyuKrjvBkXq2Z6pxfl5cgP25jG9Ru1NtjzCCTMODOwJ9kI8HiVYT
atO6qJQkjjgtqk+QRQ84IBCueqHppsKtE7tK1doJti1jhJu4MkU4rPdugsjjr/+x
Ox49P0t3BADUDGXUwO066bHLA+isevN8rc5OSUTFfHzcDbZwxgyHDMpKZpce0Gym
k+sFQ5+WYwsg9bNW+DzGyQ13GQghkx2ej48m0SDxxKVm3/8Ja8wGtrraDMUxu/m3
sVGBYe9Mz2QYebnn0xwfvId6T6xDljx8/szeQs4Pi8Ug8m+RtoHIjfeDwZtURfiX
uSq1fhV22UH47UV4QPmVqixoZV5nBT/PfgZOsNW/KszpK6HTAY+J/C59RnVRToSu
jlUe0q7ZIEODFCUHeJZ35Hd9EJenxhUGqFT2K+kD4ylgAdaOtPdZyTmrRcBXHhZP
6BArx0K0BOZSg7ZjGNLA8Wj1wuvTM07bx8gR2RLjAzMDsaLONHFruxnR/FsMp+O5
jOB/2ZEz2DxdziiMd9sqQuhCxwdRoXd49etvv2Q+ympFA4f5wsKrff7PXF7P0oB6
51Vs33mmqaj0mhwtjFYhK8SZQ5PpFB6hFeMiw+B86AFX/Af5cFcA1UuLLIbNNvny
OwDiTHtMO96/bcX4IRP5t5EXaqKGrj1Jy9S6cogwkE9l2vMSTJIpmSODjHoo8Czj
7JwHGpcQCe9w3QloVdDFr4vgrCqXE81e2Ag0Xzr7zFPRV99mQu5ucvJ6f1DEgpvQ
oNSXSv+s+1I/3MWd9/Izw/TlNmNw3TkaWv66vS386A9dQOgY14DKhigAxYxrLpEF
n0lajjXOrh5vGrBKBg8rWNF5e7gFUh9e/q2EkyNcloRRzz75b2ZoOpLg33Bn8ckm
waCLWJx1/PTo8i4J4fJUtJ9Ql2Y/WdeuTgx2+MDkA7snbZ4AGfAJWj0UEvsOxxRN
Qo1C6woNb/hxYGYaZoWfCAedlhO/VVO0gV62mLFmpWvcTHeg9gDmYpnxuU9aZtGq
gCMqnId3SQLm9ugaHN4pT2qfohC7DiQ0YGzd/EHyW9NlD1JLxUfKAz4wQ97lg/7a
VmNTHLpOKVtiB5J3aFIf5wAW7lY24cAwyn/rcZtEUc7izPty0xRlSbSv0H27Cuf+
uFzs35/eXRl62hjoRPuy8Ke77lWpaIuCjzX1RKNyiCr9ITEgH9dq4BJy3p4hEY+l
/Ivbfp5UW2EbNIdc/jXNGjdxoQ55km82cVJcRDlxSkr8FEzg6VH+tGc2v3a1xlKz
mxWvcJuDPmZslqRUjQpVyKS5dGuN8jylClO2XHqyRExUeBm93IhmLxbURsB39wAm
vqaG4xoGxz1VP/LekzbBO5U6ym6b/PX/EkeQE6suHb424Rz0+ZOIoQAKQDWdACD7
XJFzftPqBk4g/qxuZnJkJiK/vg33gIR73ypdf8is3caFynxm6b4VDCDhDucH/M9J
SSoY5TOuJgpBO/46Mcs9ynLbtJpCC6bw8Eh4KR7G42514ZOTnAc+TyGYUTKnIkqf
zfhSvBteMwdHWqvbIyGM8MTffC+qUOWd3fyjk7X9oAliBj7kJCO0RxDTml2KgI6O
xdWzCbmcHduLmg2OHY3Vyaj9sPWDGBMrWuZoKspEaudgweOwHxt36wfkBCDvsNw4
2pyY6xt9vZ5HupZF7jAndYrRicYXKDdNu6tqRFfCnf5qP73XzeT6UmkkXqGGoN+D
Ty4L6OrNi6K5VjyMWyau/m3GYXOCIVdLFK187MPcoklDkhEO7z3XVQpWuWwauD4a
JxS3Yltt7wCSJ/rw4mLyznCTjGr/GoZ8t/oLyM+R7tCz+sXeYSM6aAZMtwnDjKAj
falyImlpkS7OgIVXsVhNASFVPgN9F5K1kQQbWmgNu3p38Sm1q/+sDp/nVv3WhT07
cWLbNkrKlzB2ZKan1YUjLPXBNeyALLXfWQPl0O0OpANYEkvDwatj1eDriaddL9e3
0QdmOkvWuLa6Vg5I69J0syDVvPk3FYQxZYvDWoZsJrnMcIWTirUKir+vBumnQsE2
MoYxPpYOHOijTksdsGeCZjhvkiH0yW5160GZW1B4Y1BkYDtDjUHcNFD0HyQR5v+m
yL+ycpMc5+EwqMbcv4nA6yqXG7hlKLiTYzYuf42LSnA6y0q5p/3VQog2E9ZgpKQR
AS9DgMC/BdMnIwI18+OafWDN4MFxUwrA+ViGdz1UkMPAIxuczUjPvcnufyfz5C22
iaVBNaAa3K1gsPlscrMeRQm6ASjvzoVBclK1qTP64r1Eea+SM+/9GFL09ML7JK3f
RINrAW5XewvMEALGya3PTbA3fgG/hWnGSFENYmqn8HC3oRsP4bCD3QEHqwEVXbdc
/DzY6PzTaopbhhxnk7LTsUta2dqd8JRfeBiRDJhoU3jP2xnIIgZ/ocpGdbHl6VO0
us1s3ixmZCGRCMLNvIFPY+ktOkShy5MuUVWcISbSp/JeiCviDb1rO+FueQ5efqSU
VBepmV5b8SZyewGxx64Ku75HkK/BZKGhBTdHrUP3IgK4AEhuoQFV8Q/g9iCSJXtI
fSymVgrIAV8BJSltaL8uj2h4Yc4xeAaM4GMApTWirDjySZ0tPaquY9YZhH6d399X
OtHyKM1ozKjSXhKvEo35IAzRLWZvhAxq1/sAQxttwwLQ/kEOtR5DCJvtounR9iMK
G1dborafGUR1UBQHzJImANPZWMW4Ok1bPPwF/Zj6fHCpa02GWqA0Uy/xbM+i6zmF
3Rf8DwTzMn5KDoyGl7H7vcAV/h3kh1Djc3aaYYrdVOILrMZ87p2+rTArOFrS/3xF
dSCHPYCaqvCPSxco96JMHQNAEtGZ2/oo2f4aM+RIVM+RLIuwbhs1n+x+556QCPiG
Rl7Li/iTxMupP+LRLcQvoZp2y23WQCOVGXucPO26N0J0siG3rY3SmpMx9Qjh/eBX
bfVuETmm2K6hsQf/iz+FaiM9loR2qDpXlR9hVs7MTo847d0SC/HS9KRM7e4aXL0d
1j0cjt/jEVsJDweoS5dK+kl8gluV5nZ5frCi2dcyLE7NFVLpRQ8d7C9rx3NEvDXE
4bjXcnpacRjNJ+RC+JlV7SgV0NU4+vyahu2mAFup6TBdyZCrlRmrh1hxBsl27XCK
/u+Pf4IpUhTpnJ9zD8BES9jfO4KZw50rakmovDxYqQvbe9ILMzNwmMjuzUszfTHF
XWVcFaooku82cW8GecoMdTxXQagteRnyYVKsiVFxZV9Rg0IE5t8Cq/pN+h59pxhq
G7KummI936WiBs4u2ScxNCAwUqk2iahiL/8wWErV+pwqwHyDhhOL7CnWmIwwe0OK
80DsRO354YfcfDphg28go4qjAoT3PLarb1KGk4kLuR9CT22VI4Uz/D+ZUzpFmb2f
1jtwE+rBptdCAQc8SSCqDJijZMAtkvpeEUEHsr9ZBESTjz56ZvXkAO5huHeRpxsS
hspHUqzLdUZgHc92SupX7G+i6IGe69XI6NbplESNJNuydzEE3+eAz1cbicPkdIaH
gkqyzKo4kvDjUrvn285Xij2r2DYHdt5tT9x0s9MqHIyuOdNJCYuFsvu+uYivTonG
aiLO5x6GUKabIDjvyP3TlBjx4shoKpizCenZgV4dNrVvw9HtAUYbR6MZFGBjY7bu
fGoxU3YioUAMTUE/E5trHE3ncziQI/zxo+GL0rXQFyAc61LZSDkNFTJQHeS2Doby
+XXyPDZZhrsIswudBjt0GIsLTM+zBGD8cdG1CiyUnO8azsL/irzgK7x1RaFXYovj
uZHBqCXw/HM/XZtpXLO5Fc/3WDOLquWW21ElayTZYpxBC4Am2wBY239a/6YDeRjT
RpgPmkPm7yk8Blg3BTRyJxbU3o3yReuAEIxp1cl0tBgKwcBHZV+HgL5enm8QP3e/
i6L+lZQqzYhZsQKPVYJ9YaWQvUfmxhoB+HWUJhCUjrlcfv2+UEC1pdFrTcQwqHda
l0RyfzekS6sROiCuloy0stWnmcUtTRLh66SuTWLezUSnl/Uri8KwCBlwEHFtpvoj
ILaJmwBKoZzUlncPjCN/NSlFbEmxRU4uMCCS/HNOEIhGcEmUkt3T9HiFk5cnMq1B
c8jat+5lOX1AZcuAeeLp22XUmsg+87Tapn/gRJPIniwvzpBp8/8qDpgCuPrRvNx5
3p7UggOedACmtenaNxPB2QRDJGXaYRqZVc+msFEZFtzQbX3ocA1HgHIDM/aRoX4y
4BPhuaZ1MIuefyNsroX9nf4eUd3wO9JwD8X2t8LBFfZmuiqMx6wOOnHfumNvWuWw
j/xgJQSgIY35kPj5itvaaacBUeCvmUFcSQbKeYR6c0ZluUmZmhZKU0m2iO9Wp4jt
PBjllOlLuxsq8S8Hyj9iXkNZDzVad37ZYPu+pBQYMC6qDfVWJ7xnkXjRBHe7cjwM
QkxscglFoQEZmRg9l+J6c3nVE9ySkqfJXx5GtQOxj3Eo1l9F+HgD7xlYZireywN3
FEcupsBrtirJXx2N6oqpuwloUcO+CYDaMR1e88GWFgkB81rDd2XSS24LrYEiYp8p
EaOAmVRbjQtSJ6wBgMtdUrpuxRmENX1mJ488A9PaxcDM846OqJ/n47GuQB8+TGVO
sPnsdvDPNQVAXGhNA1hVXFJvNCxXmMoKEY6mT6iHMUfGB0s7QzKq8am3Xr6H0loD
pglT/y3c1g6s/rgQycjPXn+cz2Xd3iYeNS6HjDgfN0mqGSg0j85Nb4h1Z1SQM9Hq
DY1kQfMvP455K4piULFMWRtrruE45IPet+5i37KooPiQYCx67Zcr4hd/zsD2SV+Q
mk9Jp5PdKxjyuMc6+2Cyyp6xycCcw2SPqhhjDO+uKzy2i0jlzCSHqGSPNpHDcbnR
9kGphGAYN9EstUvaU99nhWipoqFNHTJ2ZiaH7rGcHgz206cUKRBCaLOdcKZkX5qa
esT+yO87zU/oRiKdY6j3QRgfJOXOe1JMiBDIxlPpeajQhOCGQeohFw+UslB+xqwj
5dydHukfcVyoEBC4n8u2vRDPTNnqnQH+VAOtnS09syze+UPFNWnPH5RG0AoBNdA0
DxlQNFpd5M/aWVv0xJfbEuJpHIgsKTuIGKy+5iLoA9p/RiO8emh8L6zLHdV9IoG4
aIX6dYBOrrj2VKlTi7mcYQ0TUEb21iAgNwrZPhPirir29UsmYHVwmLg9OM3hbpz/
7CQMG/i4WNKoxTgLD/yp1sd4XpaEhUNTrKkY74XAjnAszP37uiAATLEb/BzeZ1QN
kCoRjA0R0ApGS9znxUDiXaahgsg/MiwvZKqk7bFV//6xKHUeLDHAXIu1wk29/CPr
EpIwFxxwlJKMn10T2Zv2Fao1waDFDMXY6CbEmVV9F+AZr4GXMVfRJoOuzWVdkyyH
H6TpBY3qsICZ7cGDjwlsBRf+sC/zcydnIeXsDay9xHRHbAtuCW8Whb1Pl+6M01CY
XbvxoD9AQ2GcmBUDYT00L8pcoZGD6EgopJO6AGLo87BCQnSSM0ZNOwkVgUTayx7J
xDJvpMWh9Mh+RzNkaP1BnUBKRMRHaHGzJ0prM+X2sR2oyLBCQHo/YkR/qPnhg9/l
4zDhTiZGkOHOs/qyZPnCaMMeiGP2itTCYo2TeloptQojkp5z6cYSJCkH9mTlt5lb
68PMGAPyHnZDyOYJW5mKcNGuDqREF7R0t7X6slJxfARIjHcd1BhEK/C/hNVs5K2N
xUBYfhTtWNPtsn5XhmRBQVJvsHkOChjOnH5PlUKYo6QGcjomgbziLoQ4bQ3RJDy8
f7SOeArOltw2K92onEEViMYEY3me7s955OJfwBNBRljSlvTHUc4t1iEorYUdDoPR
NzG2RlFz1IEzFwerFGVJWvUl4atwnB7ED21Gavow9aztbNZVzgSP23Fle9u4ptmK
CEjOobwbevn/oNUofdPmaiL5HvkM1lMr3iRRayp3EgH32AWWHC32+qYRQQ8FMjLt
xCautZQ65ZVrvi3RRTsCZflJzw/FkvjKqkoHs8uFpqteYNOuK3whv+IFJup1Ie2T
MzD8r7jnNSGGg0CUHd4X1rGsjBCznSzkv0a+wy086oM6vcWCipGH+AeVVUw3/O+G
+1Fh/lQ/HBqL7+B5fJzQms6h/sruYBRFlg9SXCBTRD2Zsx22ZRyCyBPUREZB6rZO
uQxgksgEtTaCed/cedl5+Oqd/GB1aCJdVCofGNsZL1vF9lkzfaI5MD9vKrT7TBuO
6rBizu/NSnx+xV8on8GSSO0tDSaMos1k4pLCzmY5TP4ECCc/QtGXpL2Wpe5OXcXg
F+HekOcisUokJvsKYD8zQpO33tDCZFnJ3aJr2CjuA9Vy1RNOmQyPBdeU8oGBo5sh
h0VSyjIRXIzkIma57pojybOunqS9a3ny/azcddExpeCtwguCrNzLilNyaXHnueYg
s1sIb/w/KVli+Nr/qFPJe/bukb0XiW0TeSsXChQq/VWIVyeHE25m37o+k6qDUUX2
FvuXLT1Z3pAJolC69ATf39jMxNfpscf70mKStt+Dp8TGlllvLu1KPa0bXDHclRRK
y4MdmHLd1jJnGbHl63E2vcHETFH3ZW0ieW0bTSVmmg/rfvKtjH4jGKDF3L0F0DAN
sVnhGUcia0vwq+ctPtJozrC6dfdt425BTY64P7brvsXwfGcILtYE7T7IcsHyRras
fozEPuNHb0IB953n+d3T2EbnqxFiudXF+piBEZT/vXEbLYzYYmv3HHb8r+bvoeh6
tg4HHvkJwtilSh43FlCv8cqmuchaiFxbqjrQgpJiJHBuoX6iSEBq7iogFkqzGJHN
RjcauYTvqv3GcSPeHUfocTQvUsm2qHG2uQILFcIex143b+lMZndgOXtNQb9+9nXa
SRwQforNibyhmFmlTLtetqYZ0edUVJS8JXQjGrOiL+AZuRlwT9pW41qkeleQK14L
jUMf6XLFhmo+K1g+rU4gGJOjNhGwI6xHTCcLHWQKzXashxLuSNU/nHZu6gAF81Tx
871t0kUORQvCSNX/u+P0OA32r8/xbn329xd4YPmGlCjqALqv8nmTB6tcACvNWryB
Ilcd+tvL75YGcE3se0w8xoYzp7a0HG9PMHN9G/nQXsW3MU5uz8YrGrb1IlBjJFs4
9Iv0vn0dE5JYT83K+5xEqEqKIGeUS6cSwLLnujHnCBAKFtEwsyHPzeCz0gbE3Con
QSQtTip4USvl5yuOYKLn9waV7At4Oq1uq1QXTPLOkLf+3vu0+XXbDfs+5KE0URp7
bhA5ZQrO18sjlZdHjpTPxQ==
`protect END_PROTECTED
