`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mqL6MvA/srEPywFsQJUJsXSjJmucUga6U/jZj9HAnoT9pRiD08SG67HwL5t71UzM
5mWbh+7BRjaHNzsQduRTNd3D/43CNdf1+e+i19BzeSJvW9huOg/rzqbZYwC21q1M
CmTMQsx+0gWgz984I5Zxnk2L1adJRvckT//yb9nlNeUiNsDlIMaY2nMuh/i6Vfb/
VGt2YCkWN034dOcpEQI/g55KmzalfKeSXyUHBWgXWWPFtutTN7UQHSfOBNLGpCX3
DhmGm1MrZDHCnbl8L+l8Hw==
`protect END_PROTECTED
