`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0MhuQSQxKKmzLTEb7ye3cDSP3OZc55Iie9rwPiUnrwket3boHmREfxyQOND7oQd
QYFu6qhhkpoYa6tw+oHsA6228Ufqec+VMgSn5xxOPPa94xu7Qk3js1HPylEQ3Yhz
Oe8hViDD5z0IqHg9EzaxA4KunRt6bfPuCNUbij9uI0TOYXRrtZseErOoPWaxz+63
bxO6gDGH356XXMthg4rkeVFphfyJqAvpuemabT1ZVSCILyVxIPKkoQOtSD+8cjmv
rst8PL6raemJy+VGfVgu+zbdnNTjW6ZmVNEJIxvjpPATGRapmoVtxteQaBR1s716
+5S2Rs05VPVhE+cw/wo+zHH80n1WjELJ13lJ8qrXYSINAweOo8SaDBYbl5runb1n
caTlpF3Oq3LBwNw3k2Bn30KE6HA2VgwRQVH7RV0Ee/8RfX1TMTtpfJU7+gg919D3
ho+RzQFbjB5yoCWWXshgWOGQydW8bQ78uqzjnx18ziqyeTOz/xvD5FieqFvB5SwU
00K2IFljBVb6G3JmnpBq6Gisr9JBbNzCV3NDsSsK/9v/wi8jXzItfQODmbWUiMqn
EVdr7LPZYoOk852Dp44AsZ/CsSjAH3a1KwI9n1L6F+XQRsH2sOi4cmao5E9b+9Jt
/oyOgNCMgsMDlJocoppXltC/nwcJi7AXcV6tHtRCqU3coY17EghXyxwj5nqZDfLB
OMFveI/fg+kh5Zvlcho9sJGUfB5A+BCzmz400N0n+YdcAy3xLa323aUZCKpmwjMK
nv+6rui+7jATQYtAXNuufHe0VuOu+kdQdVyY6TSCMCvOGt4RWdf6kVacZVhwASLz
VH/1cQn1tB1wwnFigoDaSuV0h3Zfd/d50/b8ofjtI41XMceyr/K0Z/LTWf6j0VsL
TiZk4WYc2Yjy5x7ALtXiUPzpimutDyYzBd2BHqgMk6M2m9P6gN9qWWvskCUwV5Ba
3hILKYw/tveAS9MnIK9uDYhbsIvvxSY2TFAiNvJPWOLpEgbr86lzkwWLf0aSo/VW
cVJeKBAIlV5acuaIsfCu4/F3bA1eB4o63vURckqqdlGQM3TVyB/PYTli+LKko/rz
syDUio/6pTahV83Icf/ZUCBmpCoivzXsAg57ktzofLboP1POyvi6787PefKRVO+k
seeJGX+0Kdjh8njKeeu9RZVNWyMoLzXi27qgu7uYNXJi4Ilxam06rIlEmyrsUHbI
Umbw5iABYq1SxtqutYHOtIzCutbpAv2tcrUYoB2tJi8unwZSLGf/ZwikeRFscFUH
m05G216SDKo1YgoiptUReRNi1wd+xUhZEObZY2FMM/rsUkZ7JlFFEkaVFRMkQYb2
nGaGPRTCHmqrJ+ea2vSFWe1e4Vh9daxqbEwNJ3ux1qqdOy6X64uyDGYUPFDIOkBu
S27PQMmYhu1R4xDlPnC7+yvlwuZQcPBJenU41hmoF7wpS0O4NbasVk1eTVSqu4De
XguOdlP8YzgGOc/hfnS/XbvPNzYC2Dq51c4V+AMk2mxJaaZCCQjoz8Q0hkDueac4
ApUf9vG99geTRQkTUWk5yGxwPlTcZ9Tb9tfByVIEMykMf8qkPrlu+VVRJCYkWYdK
z+Ekq64XzzoRMs7TQeGyWNq2TNtIadkYiNWR0Px09dJUh9gVpapNFq6vJ5o39FCa
JRhDhGYnM4elhmWH+phENGv3CaQkX44yzKg+4JoXfEewJeucKnZfPrw/HKYJdcKd
`protect END_PROTECTED
