`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AzoqxMbwhZiuIfoWmGiIUWB2ka8l65BhZ7dKQPl6NC8s1EjWPuF30DWy9VDpevsR
88WPPFLVy5AOqVjrvvNurJmHZXDZV/uWoWoUo35zHSZ06zlc8AITpHbNQdkSnMEh
UXTGNsSVarLAOhKL/eTbaCSnrFZfbWIxkc5o3nXzkdryAWBEo95Fvj1NrY794zXc
qTkDQk1Q1zUsyx1WJsqty1iGRCfGbhVxsOYhlYTDlF/SAWHhiOyCPptQNyL3iRiA
TgL1CEXlnbM8cCc42Jyn+S+GFQGqvfOs3IJsM4KUteUqgvxPCnsw4u5MjNxNYL8w
l1jx23jsUzl9LTEcMZRiAes17Ogseg/JvwSMSM3jzMMUFga2nuKCA8+jLoO0T7l5
XbWM+yYhRxZgWeC1PhbW0XVjzMBb9TlAoGqZjCBi7dKZeTg23uWGt6HIhIz1v1Cu
CiIHzmut9wfBEQMNgwEavOFChINA8czdycIl3BDsL4+Ny5MN4YTMPXHQQOUds9iR
Bv+qigvtFCK0PMVE5923+eAp470V3UcbQR7eYBY2N+PBWvMGr9FgDQQZ34c4VLAF
ZBDyGsKW0WVejmn7O+KiuKIt+l6bIhPolzeC1DX/ChPIehuvAczkc4izCnBvp3wA
iYVTviQ3z7Si8jZzVmkkGSHl5Ws+JeooPkXgxXO5Ezvv864LrSkT0hQBtBAjuaxm
oXRNk9/y0gGApoOvt3bMrkLABT7UGwJ5G21j7Ra5BunMps0czy/ukUg0m12S7L5p
pBufa3RPb2Ssewyonar81XBvCMHFyxOLFeAOMa8NFDI/LUF903LfXYHH2FrZlH/U
AAGEDQHElUfoqiEjrovdJIltVZ0sbHnlefeABUTukWr/jeF39bV48YFUMtzuQgGf
224v6sy9wV7rZK5CzzKDcdlkDV8UUEvJj2+3SIRK1RbGsnh3OesBuL5dQyQvXoRu
mSfkBpXJ/eA3VXQmqnWJsk7OFHmJtLa5/ya9p7SXqElzjnMoBBptdnL2kluOzaOL
hcMpvB9fexfrAuEi+U1/o8z7KytbN7I9++XsdaKf+8BOmC5PkIbCGpiv6E8KQfrA
8vJBpWKKr0Jtax6TIrAuk+hYa8YjTflOAEyCoFWDqvp+fdXODZRdxoNV1WCDxYQe
9IysEZjmfpbr08jFIOYvvVo0rIR8rQaS0c0T8SmpjnqGf4wt0yBpfbF/vuaJ61G/
pD+ds9qCDOwEX5XM6bP9LEOPbLdBiDk0xs2geavHgalJU8jbk0RpE8TDFAFVt5qP
7jH02DTXK2SlfUzvmdLOoNhq4S6S63Pq39URq7J5p3L2smCbWDwFtSQBCbujAPOr
72ob05CbsW5U1EqsA13OYFN4IAvHZunpwi8w2U5pUq4PaU2RakN7k4ufO7HtiHhq
KF1snPYuZ0N72QfuMoqcFpm75OueecVnpevGgkGL3fywALxZQCFMk4bMBm4tkgQ0
0JCH67UglVWD3ZgS9Cy9zSe5oKPzyjzT63KbwtHuHm+EUKTwwJOTtMwJ3C8NpzvL
sUt5s1delFmVYZcO7yMVay1YgJBKLqTcghIi5k2jc0bqNECpVCr3BwKMURo4v5HU
d8wOUKNlW00gHpb9Mcmtvy72aYZhKr8lMqXPFc4lFNEjFouV5Y0UwEyylLLHNO6C
xQKQ/9fC+WgKyrkBdQa3WHAVmd8xP8Af+BNGqFmwlEYFZwD/8oBqUWvUe647IY1x
kmQCwVQvvoeV+cqiQPLm75mIfnEkrIOYNjGC1PYranC1OKOMUrD94Hn3/rFuLDK9
ttng92fpB+ngL/GZaX2rxaIkqyRiRj1UpYfQMRDdR7OVjmdoz2RZ3KPcR90aOZUR
Ppv8EI1HQj0P9ntj8t6kX1JMsznGJFYvx5izX4eMT9ANLb2g9/e0+VnXRhS3XGTt
rl5zxXt7ojd5aMBUF4CBWGHYmsd/tVmKzwNM3hEG8K7ngYgHqama7ON0U7lAAUE/
V+TOVBX9sFQ0An4TD97gdn3TfEYv2Sw4vIgUEbfzxilMbF6z7MsOi6oW1KATDOtb
/fex+US4HCfspl+foeViD4J83W8ZtLMSpj7nZk3a/dDBoJhLz/NPFd/C7P26clVs
q8Ar0wwaTv5ebSEFPCJTMPZmRt3C5/hO4KkY+yFmE8SFBvG+8OhsKPjHjIUPKNPe
e4W7XEyNfy8Ow6yo82sUQZZWj/JJEjnVRFc4OYz2EU480eVhLZ7i0K+GIsjLLZEQ
JkzDGlNWJQCUONFI/waNl1TVSAssoSMTqouvmRGy/dTtnia/Oz/yZs0gGuUI15gi
0xV5Ar9e8m6Mp9DhjYNSlf79t30YryBdwV3uHpjfD/ZEZbmPGYHJtemJAzAvc/Vr
MtWa0/zdcIgOTQnICbq4xM+08sWT/ulW/VXkstiDr4rAUHYpfe4d4eMNNZf0l6VP
vM5h3go1st3qZa10MBPLfg==
`protect END_PROTECTED
