`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rX1aTlNmY/1hH5Strmw/QIkDgxQHvS6BVO794gSxxErc/fbWXasHgzEZ0X6wgC0m
XSqMNd60YS2Q8VdSd1/Ih5yVw1cHJO+o30A3dJ6Wr4rvE9zxCtMFuCT20bMakHjN
hrERDZcX2Zhlso/dHnhbdzOKcpNw9qPFCwI9PFqsTp8=
`protect END_PROTECTED
