`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9eoytuRdxV/Ukr9HG8fWl6eOUaD27JbSwOR1o3NT0uvLErMyIq9AWpsYZd5x/31G
oAgHjtjIfl9s/cfnOMKS4T+N2Ga4RvpvFWRRr9g23oFyZ0puiYF7RZymW1Fpi61b
eRIa6dOOuiJjJKs4uMefW8rRgvxjMw1fVzzF8FoYdYPaewNelb5mvxGpLOURnim5
/E+BIlZOOhfjhugWkF8BKZKxCC13/JxnVeSvfC9mWuCy57A8Ta139Pv2jGmFBeKK
EqKKoOzzzVEW67wZa4am1gPEQQAUs0Ke6Z3yvpkS3zgP5vuJJNRgHISHBlNCCyOd
rnO0Msi3xpHm4OAyxyaz860PYP85qfKUZakJaVbzRYI5P/ufUJ3DiDF6R4C5p7rQ
mZ/MRAQeVaYgle7cmPzdyY7/TvlgdJLuCbmNjmnQmFbOfYti6oo55khQCo8SPV21
ht3kpD1QIwqBc/N+ZsacNvcbhDnbNO+XT84STsD3wfcQtOQkxAgGz1gi1UH/pPvN
9zeEH40ADBkQTM8QuymLj6jdLdZU47vfCYzhg9ec+PzFbqFNoSNeRzoHtUOBvQWC
WrcdtUWhRowH25Po014kcUA6olWhlRYoPCVbkhYIaxGbKIPKLyzgXvAP5EgRjcrI
Jraohw7TmTdbML0h71+K83a76WUdAJC+F9+WwUnS+yWSUxbSykyil6EhKYo2va2s
`protect END_PROTECTED
