`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5cQ52hfF4t+hvwRjTXqxqHbqWBdvVtJviSkx9Un/IxE7eywUEVFk7Cot0SJ3nadk
zWnL6FcnCYQeTlLrxJFkteU5sMa7V4sCuzCxQbdp6GdzSQr3/FRl27jutwp8gQ7A
+oCN4iQ9nLlyksh3deouS8RpanqD+LGAz9hVKvldRypFOqEHJfFZlXEsMdNLCDqY
R08/e0/0nBbAb7wqJinqfrJkjZUKqlMGMRs5HY0IapQKlCfD4Y3xaxO+Gp47vlV6
a852D/QsiF/uyWSxCyUknGrkbsfz9pCYNAdN7sLp2h/vzHzST0/K+7j2e1KjGjO+
jMQ+ofmO2M0un1dyudxA3sBZR/NH/Pix2YBRuIDKxpxTnEFL7mrU8WlFt/sw4lzS
CI9wPVM9AN7HUwB5fyfD496F+SEkpLS4a/b3nBZrk3U2q/y289hXmWEjT8+kQmZE
Gn2hPwVg/PHPrtDeITS6o/HySK1JnnY06JMKdP09Qh0REWn14Fdvl4EKUSHyGYyV
plRo0lxBxSNWvYKwwZyAjMp9c+okOQwKwSt6sHjXmqmIl7mwvUpcTayXaKvyuPPp
/OjpOG7RjIiBlGRNSJI8wXBPjeoxoDapfq2VFhAWBkTdms9Z+5mxFUe4qWyqAYvQ
SRZEPnqu1yT/GvfQYhZHxHrMEQVwvoNCWUwtAFzrLauUEe+9uxIcCwDRXzWlCyrv
TeyrlJHFeIe2HTigZnzqDp/0fSMlCvbphAbm2Ad3r4CERsIT0QUi2m9Y9jmJngVZ
kPlja2m7jD2/OFo6CmwAz0vrdYgmYlc9Pd6h6xPgQkm8yteWPEIlpXZ7c5kEo3Ec
OMsILguJ1sogq2htorbMxsXjmVA//EkdpDifLs/HmokGeTL5L5iOALCJiSqf+rwM
KoLgzUTHXInx+qVs5qd0srUCaHRGhZlNOBELXpWAC9Oxb+6E3PgeY/XLNIeKlQA1
09A7yD8pQkS7h99kzLWhv6L4AVe60nWoNeGazb+2wZeiavT1QbP86wKaIt8HhQuT
L6msggu2Ru05Efcc/MZDkMfymWFCL3pUZ9CNoxquB7uCiHQSTqjo6rvclX8a/7fz
L/QKHyGNEfb2CtorgQvfSTBCOrppLvcJgPU1IjA0B42dc6sQdCdDocrkT7a/pRrQ
hhW19/FnEiRA4tMoIUfQtHXNDFnfaz+rC1aiHL/9G2u/LFH6ff7lE3KH+dyp5eFl
nKyF4pIFiZGYFEGfbZNxlPa/EqCvmNY8umdFWiaIwlZj20Bws3X34bMufypStq4o
2jEAT3gCC/ncMnFjkiwV5VbhvH3YPbsbaJ24Adey38ktGQYGaEBh8ApmnZlTWOf6
OCATs7jvE8tr/sQHdtFDO67oNYX2ZKkk9m5HnQa6RAy4TulqSqB/m+06LxYWMkiI
mQWxiUDF3r/zkwW5eDg7swlEs1at4ITzeORh9rSg6T0yhwWT9lI5GBieC3ZDHRHJ
6XQGBE/xC456ogvZOy3uyiVINmJteeRfTrSY9diiMjNkxoHMQkP8DzmlG8/96/jD
vcbn97UZOL0W+AahWw0bBpwXnAkIiMr7AXtTFV78RobjqdOCAYuCpYgc1whLE+Bx
8ZaLo8EGI/rIDLUGWwsASnNr0mm+BCkBG4k16UTjGVBlm79zM6FvjDZAuNHMwGxm
54eCwd7IQj2CfVtR2PHgqBjL8ynQlO7VG+kZwPa7ZNgO2HaORvCknfj9IcNyrMhD
YQJqkjFDfGhXV7cH/sROKsLbchZs/66E1u1QecCQJBz0yPEnCu5Nc8zHhlA8x6xs
1q3qDf5JFjN5md4pf3uunlbO+26F36q5IrurLL6xh3IcQ0wTcIugbPq4tryoJHFT
MufFdBFN7LwhHb+8pJutjaofExgpjib66qAqwVje5DoudfbiMcIwHNfBq6HKf9Rf
GKGRIZFW1P6ZxWyLuoU9ZQ==
`protect END_PROTECTED
