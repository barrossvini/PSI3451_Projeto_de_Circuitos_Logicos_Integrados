`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PK6ge5h4AOat8Wj/teP4s9LjS2xF1ikCsf65XwWmF6TFVW7a+pSzZXIjJGC2X0eP
wnSuWnvUWUlwGCwbSHkFitfToPk0i07+rxQIKVMRrDEJqd83Lsn5n7kxPnKsS3Vt
dosDT80DTL/z9Dkf5pW1OB0ZvIUqg3rAFdG/sb6voecdoIcIhBJhSmnIhmV/GFOJ
7NewvHDFCuhXcjEgkDDKj976w0tth1veXERyVJYe2E9hqD5NXlA00w61qDrvSB/f
JR/nc00OZKrYdASEnnlLVWFMFQpROqt8ErzluRFh4K5tYkvm43Rrq5kF7YMjpIER
AE8S6GzPq5MC/3YiHhYd7rGxuQ4cbb4BgeGgY/J3DZ2zOJ6eeyGyAOlYeRV7S/Rz
WDQQHoGwEEfxQPNl6bgndmvDdJT1reriST5xIjEl+2rQrBlTDdWeBwY9dMtV9sWK
KjVqQHBLvHSsSGOTDD7DfqpPDGWVKtuxretJi1YgJHW72kyva9oPKwOdo2XEM+py
WYcGdXiVdDDMYmNaqkVIe5+vnSCh1kaTB+lcIQB4RGVrrtglBYYjeRt7cwRbZihb
0usPym+ra6wpI1//OdIt8Wj+XHphGAKHaDycWWHAolF+0Q0QmaJAmPu99XG1ALtM
84Ciezg/oJ+PHGeSzOTUDzE/jMC/abKPHfFJkDOCkFecMU+/3kx0k3r8qhA4dQut
jgUzTTnIplSh6ir1jegeAIdVd/auzgWQ9ItN0ltCKOqoeS8heyKAdU66YbPZ1nzA
byT44XuyIQ7J5I51hAKI9zTq2iDWAjd+RH4H38TPlyFpwpS/+J657xQxaexQvJBd
Oax8u51XC0l8CORG5clOqUNzAVE2xHu0Fnc1rfqfJXrwjWIsUDxfBD/11hCnW0sd
UhQSKWmA3kiU0zLFJYxvwN7mxVnr2WEzg7jNnti/1zd4oORMaAjSen96B/uqRK1O
+OK3f2O3gMJkkatsUjHMNdc4VhoJojiiL+sQrcpRjy2Tt79vOkr0U2IEgg67Lf4B
UB8vw7rlc9kbpQyQF0QkaLjFIvQP5rnTKw4szGpNicQRtRfJa53HgV7HBa+xumae
A/DW/cZR+pzJUBY7DhAA74kV5EjaovCaSNIV/me3HLQ=
`protect END_PROTECTED
