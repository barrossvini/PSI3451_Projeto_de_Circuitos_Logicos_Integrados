`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
woOlJ5irsr8FcUEmyA7VrVTixINFkRL9qMRthjBQ04IOKHVHEBERGM7rHKPdl58f
vV/HSYvfrjrng7W0s9TWdlDW+hLAMyGa9RyvmXcKPd5MzyKs1AVbyleqCgMd0FUP
qENtE796cILnvNHz2FhvrSJQunFD0r40AzpjEUVokK9/HEs4mQspLPx5QJnUHhYf
ymgHZqVgJO8MyjA1IPLDR+xnu/OyOQQMm078PPKgC0tVjHP+wOe6aFfneyvefX2U
rsQEtXqVworK8WLbDSyx3STRhK1MFLC2z6YviDyEtrhMf70qSKm6iJzY448z03W1
xBtEzXVq9Vcwhj3/I1Slj+gckpmsC2CXadu/V9eJe6PmZLMX4OOxnM11if6SL55F
mHIXNG/E7hclk/UCV95egOtXcUW2viLdGcG6U9wKUodj5iHi5eBcK7KWvSwnnGOc
Q6eGUwRzHqu7p6M6rsGjrXkFuAOn3PCTdoKlfwhrHVHs4h07v57oMTf+LCV3bbax
obcHKwqLqHS6ZOLn8/RkUy2qR/zSs9G5dxUc9P8LIJ6apxaA/PnbCkcIZjkAE5SA
IuBmHysTFCl0mPWVMC+FYv6GVr2v2lGmTmLoGDMyTUJDIX/D4Wa03DGvZ/220oOK
wO5yccicc+7PFjf+MYx75h1Gq5EobmgDT3051dKr41yRTfRI+2DD7r0+2RzT/bbN
LzBshPEW6yM6BxxQebYWIpqLDsZgIxYJHC0ToZTnUUMP+qmmp4zSsvAVPavAz2zU
DFHKQ49BeWs+rimb0a/geSNi/VpVs0nzegEcxJYyuD8tCYesg0wk9lQRmvlJhJbq
EyeWsEkM5sCynkNuplVz2En0pcr2HTH7Loq/6mLzWmzoMSUlRQy6qQqlQa3Txv82
dHQ2bt1o5KMU3iRFeq0wypTYabz30HVGQZWmp7r1qKB67KYEkvgohOz1QZczKK/z
MWLwOTcjfsShqZpVMdTXjeAIF7LcrBF5rj1oVDcqCxPfCHTvSFigUN4N/c2+wCxM
0Hfu5emcczfNx3gZI7F97r1AVke81tX1QXhHa8hfW3zm11rQjKeqa7BMbtfqpU8X
`protect END_PROTECTED
