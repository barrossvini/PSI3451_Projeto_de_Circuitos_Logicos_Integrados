`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bmrBCffS8uN5WapTTv+mduHdEg9DXuZaVMzxi9vwAtvnFNUdjShMqMAFwZUlVbTa
MZNUVsdnARPsT6Er1H2c5SObkMEoNpx8uqj43eBZfHZlXnkysiMGbVmpXe25RPVg
2tGyK6X9S9YbdY6ouD4ilFJPVZqb17tsG73vd95wky7FPvyOjxMqz8HmfZFePXH4
FS/caYbatrIETxz6+lQ/kEv9LFYXS2QOFxmkKYUkfX5HkDDCdLRGw3pktp5dgdhY
CQJZc8UxB168iJ+e0WTDebNSShTcHfXhVdbOGtElWq9suMT/uubioh4m8C3xIJJL
Efx3Hs9F4cnTOHpdtRE1j3HjMk7KrhvIBm8ECTFVjkWFrCPIoD6s3g5ZXzStxrJ0
MdSuYZO3KGNfEb2uPJwk9Pk/VL8qtbcSc3ZMRr10xTUjoCQw9RHlIzZxj3AObt6h
OnX43mPkZi9Qk9+iCzXTetFKgP/rSzvLHq8Dhyzm9RfGLJxtwUwh1yCdVwSeffPO
B+XDVYlGh8TZJFVTsJFe7CWuXUEd/jb1qvx1nqH7i+MB4ZD1nh8ARGp1SWN4ztH+
+aT7GytVm14hGOSB0NVrEmPGXHyDxAAPzlobdIy/zpUJh9l0cnou1Ip/eDPG2hlP
aN8FCumH1jDBXRnZvB8sG8fb/+zVUE7zbIdLbq9PeKfMqnF/3esuIdVhZ4wt2aED
rQo9X9T2dZhDmxXs6oTdAIVhpqOPpn3TUaB8vflqozMkZ3JxHCPeuNYCKRYSAEJe
RSELyZojleMWG/+/VBid0O7Yve/9hF4KesygSOpEyAt2rLgeQutsF0CN3SSRzUZ6
IU1BRXTwPG90jIyecrxhnAwQy7XnhjP8wmsnPX5fyrKIa4DwrpOjIgLx38+PsgiF
e5S5hc6YKWncLsoOfbJKCak3NtVHtS3+JHBKYHxv+xuN5pG0mcuUOVVZHMEP9yLX
4vf5wBuNx66qvQcbjVXBwqshhpp2gk/N7cW6S+4ZrwtGWFs+tS5By5wG2KjMEJz1
CHQ9qdcRjc0md2WlUmoFSsbndqk0i7LdvaoSUM4KMDUB5YxBrR6iwDvOUkgvzNYj
VdnrLxGAu/cjDDvflYLJlX+tTaQqRn+G1BUfcoUQE7VRq33hHv8Qtqm9j7aqz++w
c2dWTyHWOkHGYIf7pAqXeFxxUvCoaIqd8OoOWbfaLHDyNS+3glUnZ28bInVYYDji
VumcXMiDiZjGvOi9j1aZNSOqC8ath7j3vGnEEocKKLD+swKKaNzBUTjTF1klalO/
BnXb3pLDzXPLzoQWWPuOfqZcpqp3e5A/hD2EahJPzgPrz7YW6Uw0SD47Y/OBXlm7
1gtwsSiyY3YZB3FgNSb6i+mVlrFT1Rcqi5q5JxE3283KZLfNfUwLKj7YQunB3u0y
P+2WSOj+A5HE3lyy195m+E5RGd5GsCD6ZsmP/h33aIRJDQgGkfD9sXsF9wm75fBa
N+IU5RvtbvsrigMdHaeVFh56CpPQ28nxcS+XcZgaG0qe/R6vjfNPUe9+pS0b50o0
+sAhsBYo7SsbFtFrPX2mzlTBhdAZaQf3qNj0UCTjck02pMuGS4x+U4S542GyOuaP
6L9jWFL7RuldKIHSoyYQBrgnx/VpGuVMl76atgDeo8ht3VJNYEk0Y7mlgKdgiQ+4
TXnY+7QdcIzKy0r2Sl/fYgz4j1o2BvnIRnpkk2Bs1sAeOziwtXxrJSZ2SCljtfva
ZHERXBJ8YAQWfeguuC0Q/wCt2YRzydvoJcGWjmtS4Op6GPYUNmBHhT0QsKEK8kBj
e3GcGgYB0ZGZYzDxx56VqkCmxvMgXhw7GopE1I73ghUDzpely8yA/4S3K/3hiZje
MDbDJyVAmKXu0wbnS+n8ttA+iBfdEw0Pc60yNnyGG9T3d5js/4ssCArIhKdEfJa+
Fy3YpIbisaNYU/00HzA/6vIkSM3kxkOzHwyrNsxJiUo=
`protect END_PROTECTED
