`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yK1O0Es204jtNZik3CqBUrrpfcDkzQPmqBpw5ycohMteAGyHrRRsC4rMBomPrBne
G/vHxlsWEJSKyFZCmj80PV6YhhQ8BYnGHAFs7YsEC7IypEG8ar0UFWRGZCRVuCVY
etit5oWy7bf0Do6FUeWq+7A7tACsqvuN/98ljkDQaJcMmWg9PTWPWIrkFBk9gTGg
NqzFKfoch+npqlZ1YsLfvbZ4shOONNFv7XqYjLUN1/jEA7/zmhHZGn7/xNFeTwnl
PDXEOy+b5EZyVeV+/TiLhGdAwZPl5EelxP0zOg5DwRXHnbS+9rcCAwKvzNkGORe2
vlBzHnnOqi5rUNm1orlaCn0voPPWbI53+xL6QdfB0gMIJ6x8+6Q9drsLzospFRnA
eHfECSGBE2aBchkGaOtUghV/5TbM17wscFI6QSj4O0+oqbe9XelFmFUZTmBxBoi7
6rNwhdGkn3zGX0bEZ9xzmuWdWuRYoD7ZVFfgup/ps1YOfHSYgEbKijNr8KRZFSvm
M6GxSTU1399C73bR7FINKzIZPd41xsHHlWe3jp0a2FPwdqwZMq55mDAgClIAYAXB
KcQQjUwVldKQ7ht1WYG2Ln+Lk5uwP7N0NVAc8ENfQGxbcVb1Us33xbc+hbguVqNX
/AfxfUymlHpjgYlxbI+UsgyS5J+yqZs4/P+zo/1wEOgxO9A+yAKpAsklQjgqcBRZ
K+NrdU2AomwfyWEDqI37wcSDtPnl8DO5EBzbDk3INxq9nZ8IBizQg+vg3GpAokNZ
+IXyZpAAblqU4sSQ8kqaQwthdHTpEtjC5fuyQqoGmIQV/aE8tgQ28aHRr29ku9OM
d2PVCPUyYG+unefyGnZosnPNayvMsWyPac+ah8zpnhjMiUQTEkpLzKVT5eXAnhg/
bK+xC3kP7AwheYR5YMGVtj8WyF65539D6LyseMbMQIIiEMQqSp9SSA52WDgl+Jd0
6TWJD7vam4i0yFkyj/Ud9UCsX0PAEAH6eRZZZ9ZibXS52yY8s65wCBUq+SLRNoMF
QocCu30r89IQGCQ8kQKn6a0E/amQqEsa1BV8GL3kSmZQ1Ej0t+N3Ca6cZBMKoXTg
L8Tyt9+9KrvLxKN1SUUjxnS8Kagu7YokiQRppFelotk=
`protect END_PROTECTED
