`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jF3YXw7zjrsXhVZ1p7IiwTdTMTiEVnO0vdGuUAJuMZhNtmiL8ulyivqurhLCfRZ7
00DxJu2fYodpHzOqxXaPnpR9AV2/mS10UzVnwyNaJxun15CrJJlW3DUdiDvJOp94
fMLcPZlcJb7oUl0OHoJIq0hHDeQzvvZBG+MIZOUeMw1FX4JB05srx7NpHB3n1cZS
UIBcQ/RKkwUUACdrulE3tA4KSfYR54XRzVE3LO62yjDadh4okFXKvz/1cWq5atoh
moENeXcnvppTX6gkAQ1PnHKIvoMTKgDN3/7eGqvxS+W6mnfeR1CvwX+gmsNqBpLu
gN6Vg9iXnpC2wV47z+BButqsu6Tfjz78+1wxE589X9RZMceiIS0oK5B16DfgpD21
hxyVahFNHGwwRgDswE5V23ZKVsc5hNCfmJrwo9TtJaAC+2eTedKIzi2nZDKkh8MX
pGf/dEn5o8dpq6GCtOmWYw1Cvpx0qNl3MAj1NOkhrwUNNzDIXwzNtZglgdo5ZfNb
RhV2gx3i8A7QMH1svgJI0qqkG5XBO8aC0mIi3hN4VmEhF2cLycIiiQHO8C8lev5f
g6+fKOjBwTlE23RWpUdqIM5Z1WerVufhb5zmUrVJwwg6m/EcH+t0UlvzJG6FbDzz
DAe+Y3gAF1rx7BdomoMqR4vfJTh+MRDmnaNYxGVpiuhECoBghjMgRLxdkJB3gZPS
Cfm5ajgOYzKN7Agc2eePcW7yQowbQ/l5AAL3trLqtjDi3izmISlGVUS3A0PBxf/C
feNU8dluYgKWQ57wA+KoSjpVm3AmHn6ysG6is7LbjapVW3U0CCkbm95OqUieaMUM
gNY6RB15ytD88JYPUU9Ve5s1AM8BMKHbyWh2SeGsPYlcVfsp43rXvsGpOi7zi8i5
ZoFobV39WBnB8uJ3TiP3v39dyPSCs6bX4J8ndRMg3rB8o93Dz8d0pWgvgtoY4dcv
9UGpmqah+ISFCe9K3Evc1NNQ05OgYwEhCPQgApU22WCSxj8CVV+0jxmLgPBxH79g
quHgAtCOk5G+lxBRtT/qj5CnRx4RHymatJipSgClgjV+ezE7HDu8d1v3dUleUNcX
SQvYUS0D5fTrR2QNdqwCvsyRGmP0BIboZQdSfRhPWDgeGHiqhZpzL+R2nb1hBFNU
ywPbUVmktUj/jYFuFGowtv+UBwdfSSNG9LlMaXXD5fBFSnuxAm999UXA1L540D1n
Nohhikvq+di82KUVFclaIc2jKIxgvyhlgan4POsafOxZQl7KaoK6NSFmCZoK+Not
CKsbothorAuFa/2mbrjOHoV8xwvPIgtBxobc19/3xlE5FLHUHKCqyYryAzt8+Wrb
ERzyIF/bw0wyfj+279PPnE/ZoGX3EZVz4NrNBYc3OLODslTnCBUIT6x8LWZEic+6
+feDxKPHD97vApJJ0m+S/AcWCc+t4OsZjDf2aaUzPdWjsbLX0q+McZj/sjQCR3qU
f8I6cJsVkWwdMbZWaddpZWFfqh52sfFj5yocvYlsGED+dcJbNCDQdurTqBTosOH+
mAjEdUcy6HY+FUeibnTNPOAdcLRSC5rv5aABBop9T9m/+qelErfCJbTkNQCzJz2s
+JyIonPgeWrGMs4A6Q5YrXiL7zwRzjU8bJmTqaqgDPAn6fm3VXtRi4WNchVu+0Zd
VaqNfDh47QsChNbRXMT45sU37YHe8KFmJViqxZxoNGfGH6FcUwV784OfyiOkQAjX
gQrD34tjrgx3Vdk3Zh3VX+Zmy0QIDISRNOtRfetAT6MnHf2Pn5dS9eDiJ+WZLDZ9
BBJncD7fhxwES9anM5Am6JgXhDyffiBemSkeJkjlrCciCGwXzM6Uf3z581IvCfyl
4qxYUKQwJ5aZyw+tp8473MAgYSR64X4Qa3aBCNErVEDgzIXFG4A0OEGWYZ+g6o/h
Yl7DO42Z3AWVekS2Sk7/huOX7akHnMYZa55FHmWkTyk67Z3IObZ1iFiBxLyUzj6z
r7coXSPW1uIqQZE7Zxcqr9t5txrst1acOsvmn+ir24v0StZ3hdtMwGAlzk8NFFyh
ePDKv1Korscsrlp6FvgG9Bp4DNnhZ/hODKoOMI0vkrW4CMJpXc30Pw6qmAvQAsLX
7uRoNzLcJoQojaduzTeZCJuvFK2vcWRMvCVwTcDg15CGkVmo45G3W8rSC5B3pljt
bv6wcDnPg4WmoOM300ub2TP+to3jamr16xXPOoQn4x5N0xQIIjxS2zT9wszrKSne
/DcL3l7pebFt/TgkYsCKP/+OsSJorWUuPPZhMEixP0UmyvOpVDHvjGgcZqqcB0zx
s6ajo1KvUxXTaPwOiwak9H9UnxNQKuxy+nm3k9AqBTVpckT5OIcFmCD4Yt+czkgm
rt+WPaLSk3+qGtlT2Vc/6nFDfJ4kzaf7l70JXXoHU4XjxL/XUZ8JV8x0uO/MMzbs
hQHoXms64nnhz4ZWAYP4QuVdXPxyXi9+LV0rLqcOWBkYPnQfEuVgrTOJWmAlstKh
icv5Rv8zHQejsJijlCTqRl8vW71wVKnKO1yh29hAvJwIt5zDZ+O/4oE0xIKh2bLU
SfY8PYe0ZHdJivzc7rxr/HOxuSAvl4Ds3pjG8PVvC+7AtUAp/uP4vRKvxOdqxkg1
+4BZunbuckW5Mpwvpqldg+rhhWxXA0TSQGvyc1yc+DvhI4uRMBpaMA5CfK4RIhFq
w0iB3P3FPbDVSVjCUYcsL4Maw0Z0m/jKV5E6Drd6ecgK93zgWrcDTnog2JdOFDK6
/LkwkAdebGt3s1j5D3DUMBhLk3Meqv1G1BsuIDW7PW+MpU7X2RsPzDxjNgO2ROdV
aMVsXcQDE9AWUT6OpXHs6MLMg2urF4c6nYnObvZyQFP8R+CLFsovXdDhiKNE3mQp
hr6xaIEhZTcZ+DOHnm67X8Z6bNp7S3lCgnxZaJ3Y23FPZnr+b/FGPCHug1b82Fft
KVZ4wfTZCstIfTVIw+Om1Rl9wZRiVNzJ1t+7hkFnzhEq2jObkzAqMt7xDNLrf69t
YRG+iIiTtnF1uaS92es6cK7GhaM3vOuhGCPNr78mlnvQ3xx0hFPzFrPjcjtAfyx5
bJnYh76n4HSQFaqovrtmALutUVmZEerZzml3damWZjlUV/GBu12bSBDXyiwqumQz
SoK6jvENX4MA/R5D8Kv4yEEHZY6GgPafdLO80SkPIry8sl2ccoZ16Yj6p0kxem6+
hcUOLCvfr6d89AmOS43Z7c/IrW8U27T2+mHRPQ/ZlLkaC8lMl9dKedHeGVTVbRjC
LbuBOe/wwVkVXNvv2KSIBfEcs+BI5QY2a9BPaBUPc3jPLbq5Mne93BHEYhKghdvV
siYXiGKX+xgfH0cd5P75qCVMhIQVzzM3dZe/suHPomzhU+jitYRQWpePNyQBn+sn
6IigNF0ukt2UamssFw26Q2ZnmlJIOMeCm0Uk0BtuN5o3PWLyhwq9HoAf+f186e+9
qUe8FJAbNcM7I/tjTNS07Z2UWZjMU/D7olbXiaL0qRxM6q9eHVZfus6Ggssm1kk+
nfY/Z0g/aXmRtwYu1TzznUJlqVCWJ67lQd+qC4tr+45O89O9BINsUdERRbk207Pz
b0tXZolCDL33FKVmptmJc0OVbclE9u+NQm8QDAOHEJu9qXWWOf4Zd8MThdTl/iYx
IqkZYPzUHXCJq1Px/2n9jh4WF3KFna27s14bOU4oxDfWSHVi0B2SnJ1+OQTLNb8X
7cJKhMjDGmdvwr4lo5vn1iPGMe0m4LtWH/rReokNoePnLq0RYLVSAiA3MHtmXiad
fE4z7DI11XTF35nYSEeLFp/2XY1u4KfTv6gGNDL141uax/WiWbc9eulKQWThAhcD
g/OT56KlzqJizPa6yxTuzAK3OADhL9OZTzP4SeZcnr8qDY7FM4iYLRD5wi9FEuQO
Vl/Mhnin+6fKXfhGx8MR4fuB/GNqT6wvLawglEDlQXamTqIEDKcEcS0thRRBBde0
YL92n1sGTLK9F3PKjeZd+V44/xVNpKg5wdbZFuARcLtHcC7JpTulbh9wEDP8KSbj
sejTchKfGxqKVHsJNPH28xVVe7VwWSaEYhHz+aDv80MISLUNc1q/Mb+QIywUz/XA
RgqtCnbSzV2T8CfQTKG5GYl383pVHwE9ZS0GjHK5sk8bT3f5JfQbEmAJIsUE3VwJ
ODDjI8cpYnBcJ624n77b0bxrvgSBTy24lxYXIp6+jh16uXLsMdXDRJLaUtE9df96
M9KV3sEO0AO7NHQNRWS4AnjGVdHlT7udt4lyAVGTrj+V4cwrJTIcaM/dYObffsTm
lzkMGVYsYTeCO9KkhC30XvC5aIkkdc8onvJyM+bEIKxX8HArWY2t8hVBMdVNJsjM
GbNgMmcd7qtEjfn6z+ipK4GRNmbGuUYmYE63xab7xklf4vf2/OVdlzkZ0ZK9Mxbm
2TMQ795y9gcjp+PpAqvZf/VqgK6MO7Mj68OmC300h+wvgnEkLoRbsw+11mVh4AIz
rhCgGZ6sO1ujrlgoEmHxPjvocVLuwFJUVsxraBdw5bVNx6SRuB0gQRZNKLyZeq2/
nP3XFZkhQSKZQ6lSxiWDh5afsmN2Y2msEK++KqFJTWrGOa3RdvQkC1od9iLf2+yc
8VKM9lVa5fkPFmUC2l2hyA==
`protect END_PROTECTED
