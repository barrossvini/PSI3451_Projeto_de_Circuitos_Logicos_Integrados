`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Q/wOu1nh/hRpW8bLMp6ypSyTJB2KMt5lqD7mWEUI41KcWvTalfoY312YyUoO0kC
Xoxd1ctR4JmaWaGcLc4PC0ERQBbIP1udfSN2Y1oRfRPOfWmqxTOH2enQADYJnqGc
M3eGOjdjAAx9eKOwprCwiPk/w+286ZmfBSpvJMxnSzXTeJZWeDZnmfZ0ZuWT5oFk
RH4CXfOZH5nEbCXFO87bwvJvtlUcM060R3n3L3l+F8n00KIruBnkvzwlpiymJjlm
gAgBuBsxs7SA7/J77CEIESgajDu2xaAfdHVWTPTmmpgO7ScdZIGkzp07Ox96K2X4
zuzlm4zAP8jeF8gWDMah4AdbQrWoitu/pXnzIsnx/BMinfICYVqiSi5tQr+8Jl7q
e0Pk4Vg35Eg81stxhbUWgwjq78ubroDJ/EEgHob5yShtLeao4upZZmcJnxT46eUf
QTimbUK6Mo79An/t/8GW5A==
`protect END_PROTECTED
