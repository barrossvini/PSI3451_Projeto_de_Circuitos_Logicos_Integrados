`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q86Hc5qIx4RPn8xBURcdH4ZyTq8Oqf+yfX1iLPvcqKvUXPrJxrVbYdtbMXQZY9Nq
/G+UMN5lQHn9M9uvtjQVzU69vDLAQeATFPEX2tmlmFBB18nblxKM5QXp8KoNAEgB
mzD/NfoKb1ZG07C2XNCmBKNvGxox2l9+O5oH+h5NzvtxpzJzypn9Nef7lxO38BlR
KgIU05YQkxPA0UTnmpO4Q657FHnU+O61MnqhENhUouclU9NOpdxuXrH0yDgtp2ge
psqz+N1hF8A+Du2S+PILEji4xw/EBMacMVhOJ2/MQNkWnXusgtsjPtN5jpHjmVDm
ts77XMhBAaugXQwZ0fKZKRfwxHrL01n/0+IvXEKenldQhGIXZM+vUbP5Fry74cuI
d0nQA0SagMjGt/nIQQLc037pht6rf0FDAcUiyvAXyuDK0cgmRodMSBCcSHOIKlTo
SCvMeAvHIhLTEV6ubGNHr88ww+urAvA/B/iCveUL16A4lxVSNXgU4sVyiyB5F89r
bNCQxZlBNiqKl7VTRXzc4G8ipGd0FtQReTeNQDykTY/s8tO7Ftzfb4B/qT1aWdsH
b0ovSPulCZ+YJDJA4/gRaC4EZV4QwmATUJz8XrlCcbSBu8uyQBKa6tFRAcLBX6J5
4KTbGtfgZhi7l9JvlHiEsOcHLT5RS0Y7jbgIG8LDco7NKfWFbDRVPsXX+/kB5SA0
Bkkb+0jawCv61nO+PK45ZLi5icm5pEkmZn+UFXsOMyKlLud8uYjjftTWFDvyaIsv
Ox9gqiCex4vrP7SO2G5bAqaWFqy/EVo/TIqMoSp8m00FO1o/oRIRUKHn5uAEcg0V
pm00cRy0hqj9yHyzWYZo7OeNhy7XxRVUpogUPaP29Y+26EOhzrbRFCayi+ts9VJD
1ebqAsB3frRbHhM5vAT14V1B+WWgcBXQmAF+AZ40P3MU6VuSmIAgJWuTHPD/Adtj
3W6/cdmpYHIVIg9IQ6VyXq3kofkgfa0HqrGFiT5AVvjibFc+aWl7jsKbYLzNiDmo
vpNbML21GhsXGneAEAxJDeSPrODOU4TRoGGSIjpXFaLLvTE9eHqx19htTIv3sjmq
pJpjt2a1fRskvMJxyKo6aoMvMxPKlTtesc7sZAGJSJcLByzgI7z+V2g44xnw9aCa
d91Unmy6czFau5MKUpDS1v5QA5N9IurxQOcy5nATO0E6pCBnoYJiNScdL8NDrJ0y
ug7XdOgm74tn67xvKfrzq7Ttj/ujfXrW63nQF2u+T1FPmAK3kWhv/ZK/MGR/ePXd
Bt0+kwURteQaG0TN+qUijK6yTZsp0SVJxpEtMXSZHzv/H1T1LqNTWjo7gx/3Cl0k
avKtqcZgn5kQU16aSVkYOKZEWUGpeYAd5eh09xX5YfAMDK+VTrHBLDwp46ikSvrN
P2tmfsJe9luy7GLiYHobpN1p4n6zY1cd04azttJHi49A6whsBCUQIZBuRjHfjJpo
Rmmf3lSI2/saLZ7X4u0FvYB0lSM71rU1PWzPFnqdvM/Ot+W128xAGT/s7JLmrO2+
h4L9xH111fGMl94sXuXoSte54iAXVGjqdVXL5s2mlLJND2cVZ4vqy12LeSHMOSm1
C4npRsgLqCoG/HNd8o/67jjq9g8URZdvbspUXX9qTnp9RGHsH1e+uk2dkJmFMCNL
F3QPq9RVThnGu2bSoxS7CerpSv3W30EjTS/y3STM0gLRF4gM9rv2r6XBg/+eVVvU
s9DIZEt2Vf53Mkju/XL6u6yJTtvCx5x1H2ujcPrMzVs7WhW1I2f4c/n30VZs1WM/
BhJNIkVyW+HADpMYWn94KNThZ9X+a44/qSYzmfNYaa6MyGPb69kl696tHa8muGT6
4rjBudocCFryi3lH1+FFL+thR4dUcg35zDLZplp6lrchhvbgR7m6J1iI6XCmQFbz
2ehJui2iXawHudkablevbKJnNEe62p7TZkCXMGdVs1RpDJhl+MQNu2bsRu0j540N
Pvo+RxBP1zt9EfDTvgHDo0BTH8Mk022JOmH6NASERPOQQcdQBIRhz//QaWLwjpzC
EmgZxuuhVDuOEg4ptS7XNVKhZIQqJK/bZl88tn21L9ZWlSRsrI5DHsDHNsrVnFqV
wLKnKUtOGiVoEYzjj+xfk/UKgYTEPTQsQqqDtnpoNcvVZyWXkxkkOt+OzFGQ36Fe
eo09I9wg03f89ZrBNsZQHJuU/hhz4BH+bYsQ+hAtwoUXnNMZilbTE+S8KbdErnwk
B5V+t/RroOfLLcpHwaIuEwhsKnsbGQXfxAn6lx72+ETiGNkRZUe1yowaiR4zB74K
UsOBjDqSN71BqRGsgfttXaHUW2D+CyRq44ex7Y30cTqxhX9lNSrNwznSX2q00nka
ebNOCZKaNa7xwRnlcEKDTJN5vG748IQwwEXyOV4OGAmuU2vZ0hlbyjy0ASHlp1Na
pWgeFfno8aWGrfxkXQLVXrAmPPZloizH0HMSsX3ImPDtqcSqMPk8C9tRhrJ0AO7Q
XSzXWRjtfP6nTLEn4ANtitrPOitXjzucVMykSjKn9/V8bUKTFrsr0+Ge23MbKhTf
F6PZ1zS1hZilVQx76JtAT3sPgtYdEeK0AVmplmXZ57voUz+UZuIJ3IgxwHc4iXeU
qCSNL80rY+aeF4xFUwZo88y2KOXsJU1NNACsgWhCcK4g4PK5TaGSaT89TIZI+6Rx
1QpCWyAWFNW9mF43UQ4gjQCCt8sz+lLEOqg3aEZDEfwj7EkP7RmobUGjtnJE0lUD
tokUKblPqjKv6S3ObJUrXe0p/GzqpCm6CpdJZJG7JtHvgVbPf5MiS+jy1BtQOXJn
EsbbUp0LX3IwUAmjZgeZ2DEo0EqbPbaa8bAT2Zy6I/FJqaQJ70yAgPjvd3lrPsDH
xuBC63asmuboTm0sMcFANmfoCALzeCB5aGkbhtxZaBQjtLqT6h6b8BY8M31Q+Dza
4217qgT6bSuqQDqmPmrkJxzZT7Wx/qreNlKjDg8CnWMHse+G4HhtITw2NXVTsBJ0
QbpFnd54F0pLZy2eU/ZxkCGJ03nmTtfWTR0jkpbg6/XC5TcpK4ucXXKg56aKZ+/E
ZtfwOLmbOip74cjG5TI1IlAXK48DHbAh/H6M9Yr1e/2D+0DD8Nwi2Fy2EGEydkHV
smyQRD8HX7jY+Qqp1pfQJgAtq6tyfTsw+b8sUZiT9IEaWI1S+8biAcn5tvuVWXiQ
cUpeDPK0iWEgXKZIwNTNHEK3rAyd7t/bkzZEzocCnI/Mnw5M3JcniREmrast42eT
0dNj5+GeF12xc8plD7clAdoZSnXHxNcYHt+LJM2SUA6iuIYDYIlhJPF9EBHh4ZqA
cJ8IBbwQ9GSR4mUfWB83p7qbeiOupGsVDm6qcAUIIaexTXq59nDOj8Nzap1q+MZn
lEn/IUmU1nYhjfh9DdQZwoGNcEJib4cKo+qPAFm82PTWT3jeceov/nne4GQdR/FQ
pyRvo1awZUeNgoCoAOD32zz3TTng2sEMRbxdGIIuENFyoZc43z7MmLaBo4cpr+Li
XnpKrW55HLxGl3ROXRlfsOZqJEa4WZtnsAioPjSwirHc3gI6ZvBIwVdBsGio7GCk
8M8Im57SnaYRLJ/L3q444nC0b16qTFYhHaWWNOIjy1WtpBEEYZotMC5oRY/2PG6j
5/gLiPQ6jxKUHObgVLmrswHilmHZRQS9frztjTkx3zeqaT1bq3CbZUbWPjhDs+oj
MmYVEXaESsP1U1W3OUI8+mRxA3YptXhvS8YP1ylZT3/OtB86rCJI46Oo4ocZxOe5
5flR7xjbHvxU+dCTEQQVykLX9A41gSlKXQXR0F4rfmIOPjRmaDHzkc0CZdmcZQ0Y
vyFF/uqF4epAF+K1ZLv6/AMv+1EI/DGSbkvEKnSv/eNwZk5v2NBiXM7s0dic9hK5
zToLDr3n0A1vBy5n7CXpCQedv93yce4VP58RveIsa3UoNrk98Ww3ra/JsLzlN0Ok
oqNBq2Sng3ZGCwSTfUOp0cZMI4Ra+4Cj973vg+1qOab7z1sTLKIt6jdkG5uFX/3c
D1ah/xQTpmMHHKai9RKmDQY+GK9mSR23ceV8yABGVI7WLNb13fJtrhLjTtvNHJUT
syTkXdh5qpSowyUDfNvi+P671rrP7OKF8SZJAcMBZILYVhkcO2TRyn+AIEvIMr6n
Bs5Ifphu3d/ie8s31KQtTyTUEiCWMInYyezAmqasF1CLJV/ACKTsbO37OtNmwCWU
NafyHNNypglIl3apLffJJQX9FYOLSHzGTVEqN/67P28iDLhcuOmQ2+sSGJDlx9bA
rrWgbY2LSO+Wa4/glSpO9SeizUirXhQ3jJybpejFZwJQKimfhGamT7y1xWAtcbcG
A2cu85IktDeWoTOW2V8251xKlNDXhFSzRv3BvKIvnqiv/pHX9d2l2o/Cmz47okaq
fqSjB7fopm+10LRGqnsCWl9zzASdUzpdeeHfyEqpI80UYTG1gwGqyNfdPjTIKb+V
ZX1ORsSbI+bVPdQMnfVwq48WAxNZQko9rav/X/2NMChgscGXJc8UrCFD1So4N2My
1D/v1c+NyZpmY/c4Rvf0PthQYGv75oObBM3tsgo9zH1+mSgjlBJBdjxK8SRkWDgL
9KgJar8IJZcmDB6XVNS/60V4wU5ZtqNmIs5SD2eHUrf68OY5up6zb8TxWGWj1wHW
QJKu6OIg7PGBTVE4pZtuoVlX/PuABkPOXmWzNo06nwIBhJ2UtBbK2b2gBYMK9eE2
8EEkDOW62XJzRgEsBF2csBd8dtMQdivV5ukIiaXA5Nj00yTUVGZ6n+Ab3fzbLnCd
njrcOdHYa6JsNYUqVHKJwdECNXMknAA3ijSIZaR/D3zdkGK4pMcVJLcXR5oaIh5R
qG4X7YLzTj+soyjq+csHTTAJJGMBSjt9vXxKd8pCvM6ubvQT/E1qKi6ypbcs3L0T
0NAhWdqYfqnyyn3o0mPBsOYYwYWIlG/6g6eaQW1IO/4QjOSMAODwsiXVQn/qMNP3
rMJvIA99piTVG9MrFt3JseVWnwwx5cieCuZ22gnBg7WBAifmz0diEW168bla3g9T
+SZtrvxwTX6vTl2SlG4/EVfIxfh4YOP7WGJnINcVS4CaGvTiPu/y9/wX59N8F7AO
z+loK81aJVCDV1l9tSMdaxDotSd/2taG0324Hkf9UTF+OjObPj6oQBAH4lBkioyI
NKY2Nj9y2+L7n0IiaYfMVz5ZJupnDXx5F/jFA/rjNurIgZTQ9zSQ25v/9NppWuZw
mOammcfhCIB8nWmhGKVOJI5Oy82l6bMRBqG6agtEjRxlaIiSRT87eRtPNq/DNuCV
4415+8Ete1lmG3ECMnZnHN+LaVDjW8iD+WWJhdRlCeh1a6XtmpHNddbksZPxty7G
aUazambwa/HVku9sYA84UQtCORjmwE8xoREDkhx9lLYkDxg1ulc7ip+4ZRD2KbEJ
Ti8PVercA3tYf7MG506Mwxh4VRx+XEa8Q7Io9Ukl/+6ZIMNigcnIrpFU/E1CqwAX
8SObbRZsQ9boqKGzAyfcSqUmXueFiWZunc/l5AaAHR5GSbfsbke499bTSAW8lYGd
HK0CUX0mEZkC4BRPR1RvFRBqaMfGLKIrRzxG/zQam4bHMXvvysAoPyFoRYsK71vC
vuStkB+2/BKQeBZoh2j+72JyU7NatRQO/kycpXF/kUdAh9n4A72i11M8zeQwo41h
A1NHFa58xv9M4ZWX9/jgj6Ot8ZbxU/Swl2+Bz513UnVCb+9TVfUkG6dAxoPTaWn8
Auquaw5map8UwM4TvtgZ7uF4eK1udnOc2db425FdFJUNGalrAJu+vWCN9zbW0Tf3
0jC2BHKs0FZ5bNIiHTx5sp/HJND7Qwqr8lfyhVTbdqoOMCvordDhuaa5HTa50ArI
ylFaOzV7S5s3+v5gSj9g1EPBdodw8ZmgHsRhvJlYWKKWCFe8Is89KFilXot3Oe1Y
BIhcz0XxFfy1wunpEFfkYmjq1P+E67ZHEyyU1Xe4usq84PtwT1WZM7wKbY7z/vHB
xq6ARtWEReuf/FaG8aAqpfymNiiM1Z2Bpak1dTUWzku6lrnAimJ+TSD+5SFLxh2N
PoZ7WKgL1kcI7WUqBY+xvG3aF2wm8XCQ0Qk4ItYPu2Sl7uw6msWwF4htgItxzBNa
OO32+Yh8EHHScQOqdZgkVCC98yxzswK91GdO9mKR5vHndedA3KzOjvbUrK+JXVei
Pt1QyOsUGZKogXpZ1GTwmZaJE6tA9AovrJzJVqMUzWYN3k1pXThxRaZlwQuEyKAQ
fvHiGJXYUyuR0H5ptJK8rKuQOzrmdPVXDGk8Y6kJ2/OwWFBxU9iWJGjj2mh49bi6
dxo8VphQCbMIkXABiSDSL1QjEBPlPEIaon8vuG2oa7HSU2Bxi1z2+w0pxI77LlbZ
YtD2G1T7AJd+bb+8uYyH05J4h2hY4sxZFVQbQerwg2aj2sROcimbgQMVw5J4TjDO
g+wVpGB9MkzxEi3OVq+o9XNZGqM1qOJ6BOeqDgmxD7p8waVv5o+PPrNo6rCJNIza
leqxKjH2ivBOIgBjkkIPHTxFvPwwVm3E3k94tOnjaj3V4zvuju4gKYPrT2885DWT
BIBNoPeUF9pSarYtaS5dHF+tBBi2Wm0/iy9iWnt1vj+C+O2bDJ5PxkzOS0IuDN5x
1mf2Vf5dNHZKKg4Xw4CKazN/+0T+YspteGAe6nLDDZtQJxsXsux1KD3O6GH7RpKk
pzRp7cY8R8ugyXkym9/ulG+UwPmPuHjOHX9VZYHnV7eZHtk53bKcHlinMps0t6HX
JQCfe8C/0mSYiHj9/ez0ymnRDddvpOX/1AZPxxEy+OXUjRBrsu4NE5TViROVHAzi
HFJkk6GsiNRc33FkZUPbo8SyQ/SJfcuPX5akPok2rzoRDlkySlk2E4Colh47o35U
u2Ad1lkI5J6KOQirPze1XE33mKuDJolCkzKU/CkPRANuIzbhsttt2ysoqsUNgvBj
CLtrgDW71HTrpnEYNSiyvlgx/TBiPgw8riujZDu7o6D+EBQN4v3NaYIrDlFZyEKV
K682vxaDwLu9xYqWXhqGYKlTBb3GTVawpuFHVEsI4vcBMnkGMlZKO9x0nc/Ggf6U
TbQXrGv7A5q30A2bRYfDc6whMtikvXBiIhm8A3gpwqRYXBmf9jHavuCNcnzRY6fB
PnkCsK2gwsH7RG7hGm7z20HBAeYIglRArReLkPAN0jWHMtnhgI9UQOBtA48coRl1
BvI4t29wPz5jwq1+cQwg+Mag61g618GtsO/G5MeY3g42dPhswT/z2TJv1uxL1vrb
jjLuQ+iejk6WVnoxaqjQagrLfuZK4JdE7zOE3g7/uHsYJTG2ueK8+WRuxi6l7nVl
NYESR5axMtqTHcJTPCRGIMBFQSxt7dG+Q0heNoi6zW53KvTVucbVM6Pq6X4YulPS
CRsWcfVZeYeCpZPDN3fdPwUqtLp4J1XosgvrCIEA38xeaLSWLb6H6Bun5IfHBguU
gc1LvcQpyst2SWC04ermEBpEzsKIUv3qsno3FJK35PWr11njcH7JH+fdkQkCwYRX
VXXiTCiPckci79frm1HsUsegw1kLAFnnvVJjp1qklm/76WbZQaKiM6dCGuVHDcY2
QAzPy9WCSQknovbD1nzbta5PJ+JmII29wUCS+q8R1KESkOyaciaoLefnvD4PDTDh
WpYBwNfR2jEE8oxd9Xn2qBHvwzGL+11H8oDBWNTTqWoYumKeAx/Rj31tW/+McALx
HVhZAsYJuN219x6Kvy8NL5r5hM9D0VtCPMq/LAH7iYLglfbwhCAjFV+ZztmBDmzo
5gKo3NvS4EJqQnEVfj5/09Zx53xrTHMQ0zQ9ckr2XzTlYz/V6bZxEFcoAHN6cIvM
c2B+IzSiMFqk2ENbrRqiksTMXhTnmK2Zn+MOPYyxcA0+1WxjoczcovfU4u6rMk00
zZEVuvcsrBjYdlFHxYx08bMHQZ9MFaHsRbEMp/qz8RWg87iSKj3SSo79kPJG5Y3v
Ju90v5BJVUDS39e4WpCWPm8FF4/MesiweivgJn30TWUu5enPex4sdAh4cmjlg7iD
yLmGLrVV81zlEJbCTCTHWTu+sy84C8nv6VymY6d8v9xdkk8I23DjhatQMPBo9c6X
1SnMpIdKTlJHcNBnHu4InIMYH9vZE0w9LFyOnb0qZduw3/ZtrOK8dZg/MTGPe8pb
6tH4i/nQWyljwwXLNlZV21U4eSuZoLARklvyLav64eeV4cK/+mfjR5EeA1IF6O5z
2OJv7R1XOY+gTpAZW/rVhNlwETy+6tFUSgkWvNZrFKKitJcWRbnNaoMZs0c+BgU3
6KpXWGpeEJZk9t3hiCheP34tYcP6yoRA7WPhUnEvBBw+nZR8GJW71fV49mylpKJg
kNY9AIuDxG1vLtqM+wClQPNriPtdnSf3cheVSCC6abWFCFF2ORp6ZLEoSFC3j3ms
BIA1P5eVpKc70TGplxIpBZSwXIofdMzqf71DbtVIUp2x5h6lgzYPp15yCiye3Upm
HFX/oQbbGFbwhV6pA85snpu/Sy9tY5T7GhjbJ5sSdHUGx4rxJdegeCjq9DlBQVOg
yQMOCcepUXS9f4rNgrjJ3PqMlnvknaPzIq75hvmnMqNlZ2a19TXpzvyLeGcUBK0H
Y9KGLgbiNT1STt/ZEeSYWO4PiPojA22341O4HtZbhwOL1wF7SMXqcnpVhXrMabsy
VNbxSOWm/XCKc0ouGg7Q92ZHGkvTg/smQxyEgENTbCjUlFtik2OBtgcxJ2UfLFMU
hwKOn/rUngThzInFA/0nZ0rd+YnvynS/kk9OrnzcXj1hPNqWo6vzg244iimHZYg5
RPmXXJKsfqT4ygc+iJ4/jmH7UF6Rc5iGGV5JKCqNg2QU0CtmjDw4c15AfnewR2Lg
JiUZQY+q7a0ITItdY2gk/sGny9v0K6lIIhp1Sx/oZkHqF6Lq9UY8CWnTLrKfLffm
WHEii1+a48qBmQgYX05SOIS3+pq9oRiqeyGeLl/cbwS36ExSTE4Fqccq2NbGqhZM
HLwYVBcUMhl0w3mhNRoaDEpiVMqr5VinRxR286Qk/dvhD9KDiLZ9TtavW6knahXA
lhRnOmrdyGd7cTic41rgLF09L45Yi5DqvuuCq9eziIHm06QuaXPUX8W0cuiyMdez
0vqu42tQUWokGd8o8JV/K30zRQynb45pqy5UwD6THcpBIjzQ5Uuw/7Z00JaoWmnb
rxtMbiJr3dEILk/eEUv58r7wfv1lihIhoupc4xa+Tv0kgImcnRlMOOuZ/5xC6uE/
YJe72tElcSjD8w4cDEtAbgjJZhKLQ52RE84UAWVdDktwaJvzGTtr/238w3/sRLaS
b5Nagisj0UcInDoT0LK13SZKiPlbTxsiCv4OzDXxr7OU4Wwc/HUhvqZILse153xG
PDwRm7tG96L/MKVPnWSPL4LJsBjYILmr4fgUQ4P/ltuGki9PSsxhqqe50jfQXsen
jHD+7K1UL+LhniOYgRz3CifOmjemzhCVdLSBcIuXFNGY5EjUSmzp2/ImkxfCZBVP
OO3CVTrA8cnc6Hs6vo5f6Sj7+mTrqvpXYLkz68zEqgDU0uRGngpbjPrAYBXGLG5P
k8r3lVtMk+sMbAYN5724aIe/MCuBXGvOi4/LUB6xbTwo44anJTpES9PN967EDNgs
CnMzuNZ+PdTvUQejlNc3X52v3K7rpuWzO+lBh5K6euNF9zXYSZVdXN5c2Y9feKxY
5iOxtzToFnan8yGxWaDijAE3kAiof3yXUKsgqQ0zcXvbgwhs5A1nRYuvip+Vxb4G
ws9a3tSnoTj9kVJP2+pdytwW6qHnnYH5ucHAy3awmWuypyT7rxN6VSHzX582GgfC
oZ05pQ4qmFN77k1WeUFMAwPSWqBsyDElTBdEQDPvGAekDLOic+4Nymdl4HlcG8mZ
+tJ6xcFwf0d/AwB1QN6pVWnScXrpFGfuDOSeoY3Zn1xudueEJl2DlAl04EEHwBjq
1bPOPmbVZdirxhM6JKQMMs0lCMHEl6gkYl7RvNzx90CefAepwrcQAEg9TP8rp+Iu
46+DgiN0NVTwa8DlijXJIw+dvQ4hO+msoHqmBbClq7gAJ7KndjMVyIzSUtbPZUom
0nGGaX1hAMd4emOyg/0ZhvmJt1Ai5TCJXy4pkZmVjEKH5F7zGqPqZzWi4W74Q8Vz
3tePtPM9gmBhQGfBnp/G60qIYEVeidHdvJYJgok1Jmuu7xUko2G8Sdp8w7J9ISpn
X66ByeB9Zs4S6TdLkhRCm38lhPet6+oIJUf2Adb5rHLiB/w5wsuoP4elamYhzaXV
xoYq+oQfvPgoKLauyn9sbpBtznzrzh17chVoRx/YIBg3gP8Y6THAqovWsm+ZA0E0
TaH7rfMgcKR0mN4YC0FcUfPu9dsgUzcoZQdvaLhyBb/hV1SDDvxExqoHkVyMACcQ
znqHSBzCmcdIiHgn7+Gm0enogVwm9j0WUpaLS/UBIc+dp18CfGjmI1suVHNIXMga
kzBf+ux9G7tcNTrGc5sxdJMaZ1zwIarqskbBVVOMGwhRhp1nZ3SsOOlRIVCTYLEi
DSWV+8LESpIgAr/7X1xIcwANGV/eseJyJLAQ+MungNtEQJBRXDayvth2UUc3HsPT
B4+iIaAWgm6clX8WHBbHGn2fyK3qavKzCI3UKtlWfMR+pUmbINRE9pu4PUZ18iBG
hct5qzVfsh6INHs+RASnk+CtB6ybOaA2amFkmfe0KjNY8T2lePUmC/FERM4Ni8z9
I7Xuu2mTQQGe4awmejgIoIrNOSQgOWMg11Ycausia96gkrn1gKlIptSdnAcnKVqm
mIEJ0kX2CRV1cdlo3fEx07zECqjkpfUuaBqut1P6LprGT9GeRIQk4UY4j7T/waK5
RerWqeISLFHYuYmrKsM8+UtzRARattPCbBshA4WJ8lpV25IsZeY/v3/m8+khABUs
mYxxYeug/apCt5gf53EksGFY1Fa9rE7I3I8RWqY+mBwjBfYIPTlRMdvz4schtSSt
tpLQgjfov2uhz2/YdKBBv63MpRDK5WdmK1uVwd1FsWldOGkT0QbdbaeJZmo6pc3H
NiZVRDD/Rq8qx+B5MItM35mNh9/CZOB3/HzmsrccoG01T19iLUbPbgmhG8acvUs+
+ifpwbz4ffZTikeI6pQbsApoJy2PoZQMvj3A/NunlGbhy3kVaJuoWvrDmQMB06CK
MPtE2c1QhXcgNri5U+K+hM59sAsVK8QzbDL80GUHqpKr+rjf5YNW2oBHvPkMHHkO
QCdmYefv84le9KJFTKqMuHoaO0J+BMU6qhI20ciHjfx9TvyQkUaj1BvYozIs11Ud
gDZOGyfsxLCy2V0j7hiEFOci1jX2N6Cf8bQtOnQs0pSxAy+rr2MePEeuBDskmYyc
x3f5MqDfeUPW9rd6md3UHvIv73vUZRPQPyBYLL3lmbDqCfpOGe79kJTEroC6hFJ7
NHZULnlT6s6+KWSF28AaNbssf1lhu+baefff3UAFrE9RpksvdDu/isYMUelWw03l
k+yn8isJpjoXOnwCaQZiIxi7euzrajoKhQLneP2vQgs+1H+yfe4XC8hWb7yXh7Te
XsKAWrens9AFmZOdfGil5ER81tza5E8yv1kj9N1pcSzsBS6xXfOSwj9/2KXz2CYN
qFthlH1ejWqtJNkElUTsqyGkF8rQrmpdTywg/UBVJlEhSE/x1BZL7aNTcdD8SPek
ND5F0nxKTz6rsuIbR3TLShA4KAVshRYNl4on72o8Ji++Nr61kS13kgrT6cQ4HD9y
chvh1SM9a3G+KxKxZf1/TJuKNX00ZOU7lEVWOlSXrkoJ5cGNKWaWnqi+J8rWtI3s
4ociQv/F2XWrtn7zskIogJrJ5LaVZsSiXRxly2To7j8xB9X5o1PpHwxTw7qa6s/C
fjUG8OqAJYfwtwjfZ/rCGCYD1ogLeH7DbHj/lDA9n1et/vP2tOE+/d995aEKKpZg
gY7MiC5JkQAIrKmO0/6SqXFqP32mgbfkInUU98fIZ/DDWghAYyMN9dC9CB2WZexp
NUEsRVuTj698hU5SVzO5nxiYXNfgCNR4rBtXlMdCMdx4MXnsKxgWl6Xfhi70wNad
ADkFJaK9bedQKA/EL5OL2yKQLjfWmnKXFAbmh27bSrNSn4zgsVjyA3QXMkXyfVQp
cOXGxWOQKd/xN0h3gaR/Lta/Te5kyCvSw6dnLCx4zqN5XxCEKS7rxb+963L9WKk3
oCi3nFyiFYOOfFKy4tEmnVpCslsCSQzUCcCWczba0FcKhKQ2MRfdaVTasZK6Hfsx
3RYM6kIjUe94Q4cDR749+p2c2xvoPQOabZuL2liI1FGZ0VFNE3fjRDHCdjHV1c5T
nNCSFnKQA2P5Tyg9TASKrGBndLRugOI6R6WpyBCnFOU6mRigUs8jOWCnkF4bs1sj
0Xp6LhEtxYlwLOlsukEcW8jeaV4WVz1bOSvHO+QDZRTcQLjELBVTyQ/CsBsMWhR6
jaV/a4SKHoy5lPR6IdaTskRFlJnRH08c0/v7F6qXFS7d+6NuPv5BE/sSiFLBsXUf
bT+/9XzKWG3o+ZhPiDpn7ooRvRUD5G+7TCXst15dhpq1Hv6iFm0IMRc1/WZmNjTX
/ZXjYsNjarnFOgwYo7reP1EVQbERwU3jGr3eKmqCOpLmYmdw7x1qSMkxE1AOfoJy
6OcmUtJkzT0Z1WKzn0qYvB/eNvjS2rlTG9AqZ7UTy2bw2GODdm/OqS/Pi8T/qYUm
Huf/hrZbfgoSXVbmw9+tGjhoij9IDREXBnTmY4KYf6nz/6ccMHw2cbsOI6edkXBr
r1cz3FMylBZHWFqe679CnltKUsNu3+OWxj+HCUqLlE24PFvqRngKpHSyrOu+40sn
XikslHnSlm2N3NKrvfk+nIgaTX9vRw0M5stUGeOGk0ln3a9HiEW3ACJduqe08R/G
h+iCGTuOCjRUiGDUMvd9zJM4Q7ms9MYE2W/MZ0n0tUnb/fyWofHJiWjDIVToCmAQ
+Re//Yq84hNtS8E8YCb1h/tyZzYEpIr4uvW+zER64jh0nK/+KU7dRjFRS2Bdxb8d
lfeOcspDogJjZrAdf3vymkVFPFYwWQlRxqjm66uAdpfQebDci8y7VCL0yOSmsuh8
sjKUfJza4426wpCbm9qQj+GIHATaLD3bfAGEvEA/wN9o0AKSBgw+Q834ZebInhvK
y9FQ1Nfx81+YZhybqVUjFyBCLjgejGcmMdOg1vf41eo=
`protect END_PROTECTED
