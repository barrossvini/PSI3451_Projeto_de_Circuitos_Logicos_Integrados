`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRTKJuMpdLJzqtANcIw3P8rabC3xxin1uKNX46bhzV0ISnVwqVtWFpgkyq3DcBrA
20Rkdb2qD16Mu0ADYBE3MfFq0Z6FNdT7nPSHFdRpsKlYFh59orRwYPznbGzrDEF9
Db9ceJOmgOLRlvYcA9h5Fgb3R4bZxJvaoAisG1DKhuKmcxIQJn1Xf/rfxDW7Q0am
lLbBYargOA3SQE11C+7WjILWoP0rahqFjaODwL1gcOiWtzUeRUWUlb4tmr7aGW2O
WbTG3sGoxWmVXHw04V94CBD+0aR0B9Xi1fV4YtySIeB6RcgeeNST4kQP1RsHt88E
ljlMo6giHQZFXgcbesQCiDqNI9pabg1I00BZPhEZbc8rCa2S8D10edhl0+c7ShpN
uo3PxUMTUnvsabiq/pwhOO1C3E69ci53Uwppw1fhGeUkPIDZSE1BbjzEyl9CRpLJ
YElGFkRnenfsXf+e6szRlpfZa64KzX4uWmno5BmUkn6rablXAG+iAzJbDDFZ86CU
oKURyW1mmxSGfWuf032499KaoLmSj1kUwanoTje3/Fg7YVjouLwg5GsHY/zNNcWB
1nZOg0zegtJRZeT7Lhkc2fWV8JDUZXLBN8iN5vMH3E/4a4+Bmen5Ico9T3rVcw2t
LrI9TpTf0djpj+nMG3Y78boYc/n3O/7OmjiuNVutdEyVnqHlQdRBIuIVwkW3QQB1
shWzjWFOpgNLXh67pBpPc3CVhUwhijA4QD13+45c+Y72+/PgI1WnUnYK5MmRwRjI
k0zzyuvt3jbiw6E2YodoylCJTDD1MyBy22JAgN1CUAiqNe1DTgrZ/BXG6vGFGd8u
YMe6YAL7g3XKgI1GORytXSrClKWq0C+GlfkmonpSkD3NBbSNy326jn/Uqr/ERG4i
hU0PMJBvREW6ZReYTfzIx5MOaSi2v4l3ydN6GMmuc/XT08UmhQdXfqHOPqQZ9gdh
U5rklmjspIkzeDcoSUnS24yF596UpskjGjZ2paU9bHQIttLNpYAXhMsO6WfDwQT6
Jz+h2sPV4RO57kUNo9GoeyWtlLVWpbtzmUhXNJXb0TvTyojwEOmKc2WvY5K22ij7
fNHnNkEzd5NUfSOx4d1Z7RLcNBmnGWuRjU6EjbCWitfyBm5Z34giZ8Hj7y98M2pa
5mOq2bgGu31pDu9jPlXhVJkyisvZRF2C5vRjiUXShlWsJNlRNXYr6h/eafx4gwuk
bUs1cG9hU6tajMrLO/RXS0YI5fLBqnjVkM4m+TxG1ywbrHL2/XmluaVJAK4rE34A
wp23gV/DmHKAhUDhzsHzFp8g7FjS565C3oAHLRRqBQ+8gg3kxARsQ9IPrUhw+kSL
RcVA5ku4iRRtY54p/Ys5TbHX3lurGkhcjByqQqVH7xkfcdXjVKIjC9KlM9Wughdr
WejpZU7hmfCvQx8dVXwkWPlveSwRMLi5lW/C13A1N2drAvO40w3fL0L82cmUAF0H
xxnflRfIG0bq3SWl5Gi8H2M2LY4SUqiE1FzKz0IYqfdro+S9ViwExWteo2PGzW15
WyzRG68b0CFXwTI8b5aKmjZ62pbRqfRXvBhlXPck3haqInENG6L/J0wR112m89rn
1BQ/EFwlI6xu47WwafXtL2OakP2Vp7Yks7t8YrLTJ1+XDMi6GntHbSZWVbIlRx9o
77cLlzMHaitABktuIYFs1muOlqftKpqxZcabm1mjWYhvw/LL6Hnm9CRo9N6/j+5n
WtzDTHM2b1CT4Xe68u4O3m7K0eiJPCJ4/tFx0zX51f1AR0XaoOdo7BZIE9TH2h00
glPA7M0ToVqPoNm+ruwruo6il1ZRcYLNfuT/0YrwykNaYLKdvCE/1lnKQXMjvQ1/
qKCwKL73tmobBwi1p7PtqeucFOn1Sli0xam3gHAzJXkqtg3mjn8eC47WNkfoYiY2
YnUj9/t57on0agycHn18NQsnTtup5T8j5iJo7YY3XzepzGtYG75Wxgm194VY0s04
lUNO2yvwVneXbmem317qCwXJ1JFyJ+Xxr2Bpf24A6C8tqsBHgzCv3Lk1d6q9ra2x
WssjgZ+GjvWmjgmLiZe0N+kCEs8I2jShofBq+hPD8VYwZFllM6mCQrUXGGwQzb2F
COSGA3UgBz7B76pvsm4mAqYk4NUqNGiVKu1XYySfXn0Y24alM94WVwNr4ygbviDz
Vuyb7M1TQ1DdFMKNulwbPKqmY+NAKPqbA25uB1phdWWSrEp+8Hmr4H6/3WzgS9gL
QTfV+1b3WjrHoSItD/nd48JWmjdV7n+5gV7QcPTw9+J6xXP+0VCWVH95s62q4u9y
+YSQOrdeOXdfF4tsoXOnqdBz4BHwsveHICwvF5uHe8n3HO8PwOuS7gdvw2grxs8r
+RYqS+xp9nrH7TOllHnizUyDuFfJLw65myEcaKvusNWnaPCb9iSNjar9bqOteoth
dinOHIVdt8K1fs88PrG9evP+PHy9cKPCHOyjjpeAPDUvkcL/UHVPGBWXJxBlldH6
w7RGtP65X9ugx3TckoKumGqA7hmzweR4BbuT3OvLJJyZPYiJ2dIrUhiPgCa7yc8a
ivyX98TQjYVCLLxsfUJJssxZbxi2GPqeJbX3ZqepHAFppyA/TB6HQNeE5/lkcaZf
9sP0VBEZ0Cc1+r0FauMHUwY4VyTllde0FlbWKgCxjvd9jv1O1HF8Nuv6jZ1Zz1pC
/vEZXLkQJE0rasEWUTQvDKll/53bp44vU2F+S1dmP+ntX3iJVd7epCLYg4UhCL6w
/qs8G9miaO03kzFXaWIlz+ne4fLv72/rOadaPsXcYTodAhSzZUU3+0ADQIEZnMQH
8+sCxoTMwSChdMiw0HDT3kOZD1njB57SSNZZAgdoqwAp0+R4RKGvUUbU2/jC/6eW
BTzNVhPahpC5Y8Hd2JCT23QM/ZwCdN0M5OAj7umygxOwhFQo1sGp4r6EMEYsZhwh
iz3S7OTrdwQMRb490b6oDLAW69fAB6rTct+nN2feI1cjI60JnXXY/U4tDr/sAhE+
m/WEgP4l75GODr1AW1Tk2iyPDh+WfAYXv1p2MZvriPfrOlsgng4PeLrlU64rteQl
bk/IqMv5DUqppytG9VgfL+mwelHjlHzbaBGMi0SNGtcWoZGCQlLf+Ftf711Qz6Bt
M6r7EzZiZTsB8OZ7udv3ipgq+GP/fuCJZny67x5p7Fg4EVfPbZLvN4/lGb9KILQ0
8Zc+ifQ9bNmN89AAuKJe2IbHW/hHTvQW4jJr0Wl82PqlaRT3pr+uuogaGowp5dNu
vNwhEszJei1Ir/nbL3ugkISd0kNWnGMkJKx2jny26idO6DEBqKLIZ/NFb0/pPCat
LErBww4D5rv2TtZ9o2QzJ6UhpYqZlzC+5wf2491sHK6hyRAzMccxqQSM2O5X8doK
9hi++6GOnz6NiRrRTmP+LsHIxQUcxVnppoUH97cWcEDsWAgduAjGwpQNN47DdjgR
cnRpqhXa1hMi7xHreV9sWsVhOzrr/SuUna1giVNqAMCNF3AT+pUi0BpDnbLKRw64
9KuJGYqLynTDIdHrLgSpj5wMBBbUaKmJF1Ta/lNzimb48sjmDSB/U28D3rDbHWmG
Gs8nrRtEU+s5uScoJ27I7O+p3B9ua9RVGJwUOMa/Dll1Ry7lnKkhprLs46whyopX
w7atSigDUjpjZU6eX8CvtFnpbXl+UUiRxiJD1tTVObkuCdZ86NSG42g1H9A+kunQ
JbL90N7YWnu5QOUx+BTTnHNUyVvijrBH3Ygo65FnzS41K5qp2+MpGWaOXTv+drvy
2X6rwJkNmwbUOuG/Ws8IJDxMVNUlrstiP7Ddkc0pcwCemkh6Gzbq9w95sIKnERKo
sZNy6GLY5rESJboCH58YfTfNuzgCPpLyfJ8aBeh4EZU4SRU01/un0pXY2tupCdaR
BWLyETkqlVR8X4eFjekyg/VfHHP70CaCchlldORd522y0Ggo9K7HwLNtltkCCgxy
DlJp8/kRo4iEGLiLdPkVxE3b585C39ZxwuBIggmb78pSTlKekGyJV/AyKJ/CBY2Y
TbtlvFLq1L4vxRRmQPzZYAHJvz/orQ2hUXpr++aq+kx6/n9V0pHjqeTLNGSQ6Zav
1jEhtb+3Oc0X/MJh+uiQLS2K31ge//YV/Acy2KuB4ZQegxWFJdI27fCpe9xs83io
oEWlfRC/WlGc4OHNX2AgvVe9sy3URgn3nJOmV0igZ2oGKyaUDsGlLZDKPcYaHCtM
7Vpog9v/uhJYiMBhAWK5cQI/FgcVNiX+1NkAMGhAX10oXq21y9/XbtUQdaa9Le8x
0SQadXgUtdvme9ghX45jYwndlVD/hCWL8nMIc6Eyu7JQijD3g5w8dRSoz063tTy/
iAy+NOiC/jIclUfVoWI/7rMBWEQoQmjSoGu0cqYwDCH7ALjGjwTfnAT9FgE+0JUl
SvXrkYhz1v14946ZCG/64EAswK+K95ERh0Zz0vI+NWXIvEphL/qUhX1pGk8AMLRQ
7t8kOcDucIrOlIShYGndgzqj9FY8uWblV/R9oHQZpmPw/nfJdqLGEnOzTHzMfAsC
qOmD6ptVJ7+MzZpe9+D+0A==
`protect END_PROTECTED
