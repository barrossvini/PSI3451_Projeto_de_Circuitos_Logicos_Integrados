`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SSfmgaOxFXiy1fkr77jM7SznC2sBSsVQLBugKYOiRPjHt+CBebFFmGcnizvPDTac
vgN5sj5NKqShdgW9Q6HULEez2uWwWfGqm9AXIrYN2dcVuBYyvp/KOlElTU87MoSK
keIY3Bx7gEvDF19llEIeUygm32Q6v89pCY70dv6S+FFS8rEQ5dTL9H04bp7xmd/M
sa7WPqy+kfym9KY9KSwJnIwmnpxE2A43Cemp45Cwr1uZ2Whugai5JRvLOH2eNtfW
KMRGrbaWRsqL0cWjkpnOZM0z1JSvHUYHTsAHz1z9I3pQLaEi+8+Le5mm1CtiU4FS
C2ErWJJvZmz2CzJj7tlpVuY8Z4ZkDo2Jth0dtxN3x/iXXJJiEwZXYbsQhi+xptzv
gekZLyQJ3agLkNszFCmUjX9Ed0HfAjz+SfJxz8XN6hxYitFGtZkTimvHUwMW8esK
A/iaGEryAEVb3GISUj8LFj7sLbRRo/jf631I/noYdCvl6ZRQ7urooRATJPVX1HhC
o5g6xj75RS4iKqySQaVRbmJc3myR67lHsGKCVMU775NwPOVMlCBiNsv6NB74sCXe
NSC6nPMIfy3F7AouSj/1EVIAwQ2mqy9Sez3hOCJVjXY5qRYiQQHJm8x/stvRUUDn
W/Vpkuo4cTU2uIesvzltEZ1KiXDcWEmn8OwAgvrgEHEpgcwkYJaBrYKN9NLUgR/u
cf+CB/kDOIpBpgyl/ZYPCR6O0YIGe1bAuMveo9Yse5UmvQ+hsKQ+/TpsLzXtk0s5
ASKetQDlphMRGH+dXm6lcvNAhBbClz97cSw41AYrAo6gDeUZcZu/eaFrLgBwAfbi
yfeI0eGaBKEC/SFuflF9u+sINypwXBa9WOJZRl7mbM3Ka8dqcbpQHol9W2aAT8DQ
LJNXN9K4WZQR3OM1PCgkXsV22kcGzeuelZKEfXU+4gGv8Ifdgyn6LCu2DyyTQpGu
L24w4W/sXEEAHGrpzB2bYGXS6Mg3DXusbnssGSvDGAa9upUIOMlygmu33f84lYy6
julos/4zJ6XGiY2NX20panq6nDDMzkdWgGgAYMKwlbE2iD3MEu4o1q5LicHHIsaa
JEE3VCvneuM69HcegbGG2eN8BEWFFcIL1xym4BJdzaiHBLjL3pWOIVXNiRQsSAcq
ZrpfTXmtAMx3F0fb3LiR4KKnyyAqHEBilKQu2APTaafXb+Jzior84pD1EiC6/iGE
PvXFTXX65YVUb0qtdBwGL157Eqr/mk+W3u81OFzXfVoGq+XkVJfO7SkGjMDwhhYA
5cKhWvzbmRsvdopb9OkVC96fI+vgtP4RSvrG9myxR1StE6zxNHryj3EvwGBDsoBm
BNGwHwg41ZlqiFey+bJAWURZjI2pOE+Fcch9WWBzahYqMFCiA1miYdM+sSRsbF0s
7W4rMvYHRMZELcI8AFUGm0sxQ1NPLXXrD+FANNic7v/yz2iyfeMoCqjtXXQENfNf
UgBCihFO+jGE8NwXAXisFPbOlZFqQfqKkxzMVXaU2sGTQ3AVBZh5KOzSdZAR6+ZO
YEfMgnoroUnPoSE8PYwJBssPBqh+ev4nChX4ZpdHZFSQYZ9u1zj41x3W8R/hQpGU
2jMUnZaPjVd25u7WChVGDNwTfAQWS2Q1KaqQnq5jmfADQW7ksY5BX/sVWS2ZOIXG
AaNcwZOGrF9wlQ+tkhD94iSu44CRHO/ulydfz3RNNxNSfGcFWwTsvcJk6WYx+xBN
aYk+HpSFH9XdO0ganoYKS3mguTTmU8tWUFzBwkXhpR705hTb+NSsU8pnZtLMqDBr
+4tqEPdWw159TcYhEyD9hGcEekH6QJiei+RHjCpa6igAoX9VVKEFNbptzJQ/RMM8
CE3hufb8jICVSmWCwkXfkQm57kr+fDKUzEF22rFmNlhAKTVjpMFVrSlTlci/T9kq
NdfGhOb58lMkYjf3e9XvHiokT/mICZ/zM82jgvAJ5ONbZzcfLedz8tqqPvg/ww/y
5jlEsW+tXr8sYoH2M0kd+s2BC/VncxlF9emSZud6qxNJIl4iAY8fvkaovklidhCX
DLP/qTzLBJ3CGRJG9F66VjERhc/ZZG7H6Fza78ZyIjXZFM/tBP4+i+yfP/g/8l+X
anjhRlk4d8pfaojGU6Th1TIQG4RSFyGXph8L/FiyQ1uW5dKmgJxiLXNC1aZ0qR44
54xUdgm3oWpC2kVkHwUc8zuvLO0rffTj2bPYtgssnURetFSts4ofVS2SFb4/g4IN
FWFF3ByY3ExO/5lsgGQW4V5AcvM9RWV/qtkdWCZ7ZQ6WnTNs9ja4HXhUOZ21tO5L
EDs971dVab91eBbx+P6zOE3UjpQnxBp+lMZTFoLZhYPcr6Vg9p0vmyKbJanPl8oz
VcvtIUonGTIR+hz/CvdUsA3fFK8uPPw67RH87ARDb+b0pDZu2x142AsYn3ODjnT0
uZBkveIlepQDkLShtLIPjsY2aju9fiukkGHSPCYwLX+AuLCr/g9vOIJ+/gqau99K
9Dzz5/74ZV0dgWWeaBKtKg==
`protect END_PROTECTED
