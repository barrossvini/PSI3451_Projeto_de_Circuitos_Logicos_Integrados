`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R3D4iWEkkKqZy35JfSbSZ4Xn25/raEgo1o3BDck+jQDPk7Y0jJU0e/O3DxKVTLhE
/1heZP6VWE6EH5UpGRqfncgutzqHYajn7xjsVDMe+L+LyiDXwtDGjxSRDu28z/9U
mj46HlZBF4mm7VI7E1MpM+3iYrVTuCwW4ESonQjYVc9RMpBCPtsXWm/fn5UyGLpl
p1w0Yh7FpzVKJCGHl2kUvVlPgjc1Crk9DF72VfWWFpZV770i8J7cPEkvaRapVhOo
v/0K37IUcoKx0QA4o1NR1Z0e2D4IYGv0RnEuqCHxvBmAo9z3Rf5cMhazOeCh9gjz
bk/VtJd8rQg+IFbPa4QAN28F+NywOR3CIchRe86pn+YQnHNAv5mf8KYsvESZyDSi
pkDpfEwlsYEyOg2cgOYAy79mXMSZbzIfXcUUIEuxXjbwTvdRd2/apeZSkykRoxvY
mhvIghaGjFeU1Lsx58WROXIkFJeZN5JqBqyG/CZWyg4k3IA8Qy8l656NSOR0+L59
v42RVP1/GFpdvybhQFEtmSyVucnMdM0SC3naCHSLQYDveRI13EBEyLmnf6qH2De6
OoS7CRfTkHszqACDL/it8Pbme9jY8cPQxbvQq3Da6jh6hWVqICkrFtqwvzQ/F2Ha
9XPvO6eDDnLwFAF6YeVYdCIxn190QjbE0i1ikdfYYso2N1q9lfEqQlGDiv6cP4cO
PesdNpLUpS9Xr0kxsGGeCTo9V8cm1ab3q9ldqbDBgEFty24Cwyedii+mLvMASwUN
XFWJDcN9AwfrwD+J1KbkxM2dnprwJTsUSWeKFKfJhq0Q4+Itdzr+vm+r0D9FSw1C
lokfV0YwLWFnKQoYb3xiqRS/jXgD1qd0O8ambB+c1Wtjym8pLW0f5RNz5lw5CFyo
RyFq70tKFDeK99fZZh3/9wIhYP5bYZfrxUe9hEX1XoraggcPnB10+T9ArNXvnhvK
TgX41her8nltlK1Rij+xosac4mgStcbrCLgbmSt3VGSrDZ7Yhq7Ed/T7lhRRa4hV
cs33xnnuTmlWczaRBybuBW26kG25aiK6brEC37dtLJGxQQ3R5UCLxqxkd/uko2Or
vFqJVnHGsd77yyg9af7EVYad0nyc9+tbxTzQ/MrNfRz0Wq1BNUUeTH4V9cy0YppR
61oEb1xby5LyUM5vOPAP7quc5UfnRp+6BixQzgwRTMJqiAjHYSuDEP2FsU5mux0s
V8NOhCp0PgRkPSRseK7DAqu44VQ6MJwC1PjApuQFy2ZFXq0/Yk9poJcEes6nTFoL
YrAqfJ8UFYkIqNh25kL90/sjduBwPuc/GYAlVUKTb4vTonGm9/w6+J2R85rQ+Myl
V3nISUchf/LRtwiW/tRVv2C6QzSc7LVLIIAF2iYHBWyXeGpjJhI5la1TnSeVdqoB
KRkFev2kCop5A5LXw4xjdXU26izkx+z8q2YAg3Qes6VdTDXdsRUbrxU5WGTKDxi8
eVqN806ueWILplVLCejckgoD2l8M+8YnkZIssonE7DmiU/SUZv6vaaAYBgxbm7kk
xSDtG9s6ZjABuyD0SkcGdPBxpOA9pJlyhKHfO1LrpD5GEsS86EgwwGhQ3Ym+8MvT
H5IhB5zZSUxRT+cl6WG2wQ3T3wbB8yE+wTRNl/fBaahENEpy68R5i6rCj3/2Ghqx
pCaybh4uVURB5BlJ+H2UasMCfBKNnIO2KfVikbvcLzv07fXxR1Jw9tt1YwCPEDCq
VAyO5hAayAnDktz+JEpoksnbV3289jfeTTay+YPmh+girS8e4eEanh1N9SI5ccpN
Y7c/1g4CHm9tnDTzz3q/I1M0TUuguDCJxZ+lBmQKdOzWb0p2R5x9ff7t8fYOXH8/
Qn3dCEi5eMnR4DEx9YBnJrtXPjlO0QEI36F8UgRfJ3AurJKl1XvM7IS8jFJ4yNRg
i9WoNeL+n8DKhdtiABsbGrICd8XR/qijk7Wg9NHXI+kHSo6/++MkugGHdEBdUGBu
HBMCD7sHhEUeqPxXInDra6MSaSI3ew9sWbiV4RKOPxQ+2TtfX1/f2R0l8PNLEETO
wNwcF5Bk/OjoDlE5hrU1CJ/59f1qIMa2VgfL02BbvNojq3nI1P0T2Qe35zQ9Lzkv
VXxJ1VMGQRq91amj1FK8bkXVaQOwkXbSlsJ08VDersxtSfr1v6htYJkE7trvpAGc
2kPwjqmsAD0JJHZG1Q5wA7pwkdbRvSKR3XygyobnSKmAbMYUPjnwnm5Nq+iFY+yJ
8zTdNySPIE1F3DHoHCMNXXWe8zT7PPh60HoB+EQoaZxlLcW9SRS8V088BXrdEw7U
h3uIAk72iKkHuWaBxg5XzouVkcOOnD9TxpDTsDtcyqV8jiKmFiZFvL6VGCBPRCT7
trfRZ2prqVRPKeK45oGie/PG7vcgUqbEEd+Uq2MjowHa968lxEq7JiVhoAjbj6Xx
EUCpxannAKLF4PvK/CgaLqK1jsBd7ZlqLLHMGL62ADX6mJCWCG27lNc9nkM24Ob9
SXekJ8LVAVgU3FCLqraDMlP3AiDAJnJJfeMN/YPf0qDEqiTT5wauTXTz5jGWt9vg
pJi3ILqH4omdMR/tsCoN+EzMEcDRLLmJNUVTaCPo0m4vBcz/r7+QREYLEUYhBtw1
Vo7PyYsf2ZrAJpsjYjSSpd7SyswRmVYYiuz98S7mzildgsX/YnIeosRu+Sr4qnB8
83QuFR/MvPXu3rk3mwrtNkJI9Sg6U+z20kF7ku3Cl5vHd9atKWS9llrwO3V3VF2J
nZdA+loJWarM8ARYd/3S9ZN6SoRPo1S5hw4DpxNsPMwhvlF7oAzbz7jfNArTfAEj
cRxg/H4A6qHJLYvW3u0s9ITKl5lwbQTaMNLA7v0hxpAihhUFs2x58/lOGrhXIYH9
YeecDsCm9YfnpToU/JKynKw3s8uAYF/yfnW5Ckjn7usUiL0uCZv4hy0WHwwhbrG2
9DzSYUQ/2S8jwHNGoVv2UPPDWJdVi28CHGfOO6h3x9xCXU9yvubxHfdgg0QaRvBb
1UAM1hvCmBh8gyVhTVsJdQ4sAmVJdTvFMdkr9Tn0z68PsPzOetdLlcS22AltD3K4
+DSJdM32clV/ciMVixC1F7McJ+9pCrIzOBdlZq72CRBy16IX1Yni+EtfdBJkaZ91
chsmcITNCM2u2IbAP+AKirjaCze3IJoevoflXmX/dE2eYJtw5Bn+2QIPUKZZN5A/
eoHyoIb0B/sHO8Opi2gU2MjEv17JYZ5LuVSdq/14AQcAMA9BjkIJJz1HLAIiik5V
AkGrKRORDYcvfTMCXfPIo52MZk2jEwZWti89ssVtMucwxNH1STg9pXPGa/ym0vLb
MOt7kfoqEuG0OFCIfMCPMln93yjteXdlFAKvFvi/3kwysA/oPNoSBV5TVVgPsZnr
b5gEnWJCxlGopDT+8AM2+KMmRGmVAOkePi9Dra5BfR0eLyTyONjQ6oZG7X9uMxzi
29O1jhk0CKgoM8Zk2svmJ/cDlxJayWLahZZ/O6h5r80q6yfArrNMlLSKYNjaJlus
H2q71EcB5S30VFyBF6QaUmchsCDxIiFjHGTSvZRWgfs/bVkrK2aJ7+yZyuvbUY4T
yiwXG4KxWlDMI3TaQnTcy6/NxwDE+JgWTjNUuEwSF4vVtRT4LbDulpgyyliqhiwa
9coraOV13iLQuJYKzJ6NZICu5J6OymnpAQSEkUJ0wYLIjB/l8uld9msOpXD57ftk
vRzwlLdvKt/QVaiV5kPpDSCyYyEnf9eqLWJ8og48+RkqiID07a6dbD/TgYB/3oCU
vbf3RouXSVEvFsCZZvOKmT9VBIUGyxDm/K0hd5ijAcRJW2zLPUTmZFGl7MLnzmfq
QTIBQ1rO8LRpxldfgr6Lu2XQZ3gDdB8k5wT2y32ceX7BRpFcAebVNT7/FR4vyCnW
geMMvAobavUlqrcwX6MHZcvOmRCWBuIS2/PdYbQB8DOn+YtVHYxs+dzi7AFWdyXO
u54exEoY+69sp4aREeYR4pbWUXcDjuQr1z72Y2HqLkIQbULhg+uOaiyNkDouI3qS
DY+fDYs6duPGXt7aQxrbaYbDGdYWzVBt7xXVcYNKEqzdMkTT1u+h1fR/n7nm0wfo
Y8j+lBCx3OcDNLVfIQ3Nvcxsu5hbMAXp6cBd3r1X/YUB20pjF+IV9slb8Vst3yxD
ByONCee8hC4ei9V+mxyYLBMN4OxKb3f+NXYf+Z4ISxNSF5vtEFwPMM2Lw+bhWaOE
tOyUb59PL7F3Rv7GJpy7a0C2GgI2bVFOphaNSy4oYCrbieRvYQERcCuQk4lp+y+b
5uOlPFg3UNNrSZqVbMK1kS0Pv1YUQ4IZeaYR7lXx+DlMTNTubfOM9bvm1eg+Bafb
ItBEjH25Jl083vI+RSD2ZRGvwCm3YRIZbrMNGjdzXMQLdhHIKmq8WUP8XsHoFKSL
MKmjOe1e/ggLwoUoTXLxknTgPvAGmrI2uyjZGyyMzTlESuZrJlZNZR9YYodsz8sk
orvKzyF6981H6HMNOwl8s23Ls4F+xugkpZHAigDTsIYIAGo7Lg0i/jOlk9EI7vUz
9sFe0pEO3ug6s5//Z+MD7ssb3dlg6DLkF5dPnJaCkfGsOwoLlYpXayExnzb++3Fl
IieAd3PhS/mAQsayaYPrmDDmNMi+XhcOzLA55+THx9ZEJeMEX6v/4PWWYvP8bn76
cF/zNLYav6rXJfoE9iRckLKbUgaqFaOUh8fJwu3tYOKDx04JmUbkbW31UFgQsyFK
RCy3eXPgHqDkH6afkL6ShZF/zLk0HJfa4fjNQLTYBBJy3rtzuX7GaMk/Pqcglo0U
GplGRiYxa8yUBYnchmfxfFTzp0Sy/gE+kz9oGVrV6m4v2JxH/GNm17+aL1TWDTKx
IAfrCqLv6EQKO6Z7JE0uHlFbIKt4wkzxDDricPLNJRQqUxVtoMvdjNESHXubZE8L
kBm5XepmL2GWqjIFRRJOpu8FZvPT7bUQHohU0wqH27GBsqKo+GVugFxHJ5KEQ7Bx
a2itf5EHuvYW76gM0G82c4qpMWnMn4m/Ax5Hd5xddlzIxOph+U4a0QUdCFDIy4JY
aUGml0R+d8kQrT3+XvX76F47VtCFLgDl6nTkHNY02rckWvXVnjRjskL8ulggtU8c
9jA913w9/Ry+n1e6eX8IgjO9PdjeF5wnk0DCJ5Wd5ykGNl8FDKZIiYfg2T2++u1+
aRWN3oVWT/8CXc2peG6cEf2Hc55JgD0I5cFIaYwXUU8X+KU+5k2+uBmrdCGSpG61
uL8ScpHcfIynpVIHk/sUw6w5vfcj9QKdpHLqjr+IlODwCmhDy+YQBjq10cw+Paxf
yo9tDFK4mJP27mqDhXKaSQ0vgSyG0imKLbO+QYrldapf2avM43QGNXgnlEx4+vpe
CqP3AujIr/OWRbhDKoU5RLqVBmKLBLH2rVW0pNN/Uw834jT6kI1YzxZAsoBUUD4E
A6DIzJZEbbVoQCLgHev0ms991RXrYaIaSrLs72IJpKs5x1nynpnss0D7QYR/n3K5
JMHxQja8vJaTRfo5Ng66MD2574QFZXPbIZ1KBEZyUUL/2WRpFmWtMgtQgeexwqsR
5KQiHPbxFbMYh4TuFDx4xyftBZl3TH0d1AHcEFpQyu1eozphBGX4/Iaou97lkh4i
vAZwND7tsn+4laUZe4RFa7JqqNuhZ1EgcbZGfWO2M6RrLMDupn4xLj8vQy+XposI
6V+ONlVElajPdIB7NXfZID3ER0/tNBCzLVhlzRtYXsJ7+TGzWLARLQHUTuabefjR
ePm2O5owNVux5+gYynyMm6fveU74sP8A25tYdtIAb8wIHBCnFqciF4KrwG03SmMd
bGTlXzcE8Aowz7PUAGpO3a/ATqpy4kz9iea7HpXF4gaQlsqG+riXy2a1uOjt4aVA
W8peVQUDsHP2G7PuIaaVccOOB2wnJNGZvmHkNBPY8GnG+o4jfFrmRNcx4YpCeaxw
3VHl8FIfKJg6uUnw+ZYKOlRKcTeGD1yf4OB6Zif8fj/ghzPT9B1KZMsCKYtYED2E
1ok8mSTdhtGKD8UGSbpNkF8ubWl51RHFOeLLOwmMXNwar4rWZwa7XFdicUH1dRvP
f+2dgHD+JZut/P3Oh+Z52WGwgGvHMa6PW+yprZYI4sWKsmmyVLXqpy2NYXKsd765
NdS6i9P5BIxst5UIwCLahM7ffVUZbKHewywENvwwTnuMx0QcVq6DP/OwQ/YvDT3z
PYMWYGxX/JiHhG2srrgZItXhIZkzBO9GEAzVYHDq3qYxQ/JDlD6ZChQ5lK0raPPC
zlNuEhGb+e52eLDt6pYCG8cFKHGjgyaLYTuF3aIfrV1S0Z3ggflgQc+jfrWowLOq
GYLGXgtSzxTjWToZmnUb/ULESI8RhVTQEy3Z2Hr+PBRk9l1o28mguyi/bhuE9PQS
emPTyYMcKjlIktU9HX25eDjm1zbOwbUWrU4yqikZmSW7VJF8xUluNMg5Rw89bkoe
nHaAuVL0KcVgtukxPWwdvE30NjTrvKK5MTvjVhrnOt5ECzfZ4uuGGE62udyRFA5U
cEy+I6Eb2yYjQDnqn9JsJZ4emewMvxuP4qq6Cj5KspsJlBZARKr2+NBwrcNMA44c
8wLRKxF8tzF5128P/E3LhstFtMONHbYLfm63La0AlqQ548Vz2ACNAAQyau6STgTf
MGxrsDLUBGKGUFFu2jVg7EJ3UCRfh1+/0e6hQX8a30gVZKX2UMpwipWNLh8nMW2V
wSzz8FNivMHbuIs1hn6ITQSnVqhnlEvmn3+uXkf4uYzF5y9458p/Ygb5axMNIExe
uGxB0lGHBg+SHIT7Gj2PH2BPK7tVY1VaJnFHVFxvP7DfoBocUkE98zDTwxKZRZDp
POyncgThlgZYKNMSqvkhAiGNcqZ3Zf2eboNjs3zaKEcj+1DrfFg6057MqaR0mM9a
23sQ1YAeIoJ+3tX7Yw8bVWSJS0O7dEFF6fVDxXH21eQalEaBYipseY2vylrQRAsu
6B+Mr9C+J8Na2yZsMMFxu/sM75lo+86lhC5B6RPrSy67g2kyD1JravRRfz/nqoID
VV9Rp0PrNH1XmVWEnzh/M51hbRDRc2Tdik/oG/sIilE17blNcxcgVe0/0UeoVLBc
0Faj7trzjU+qrmj8+5Qdp9mRtX18e6lbzR52dmAQiaWFSSEg1q+Q65E3QYDGBTjs
AvZxXkta6bmY23q6JATaBFWvdaIa2hg5e/H7NhsE3/WiaMnrBKc/Gz92Q3JwB25y
1TprvnTGmS7l73rE4z4oUK1s78mlnXyQcwyHpIH9G4ow67WpVo7tEDtW08YoGIUh
NWLOYXdor9fn1voPR0MoSRbhhl3yXjOSIK3UFfYECdvS+Pfst+cyzhxh1j9s9tG0
K9x0iiKceZfJPbt05aa0wLXhV7bgaUnty3q+M5MJPeGMJEbMQ9L078GdUl7iD6TE
3mwjAQcB9Py79KffDf43DdAme+bewFMQ/K4b9p+Gl86bR1sNkhcq01rw7QLOXsNF
K2uYQeHt0p99a4m7XHJRbtpdgn6Q3F1AE3tQwgtj5LYdJbctoAzNPNF93SbqDwr6
fPeR2hahi6G+cIgrqanRm1B1XiZnSwS0CLk5EhTpqkeCnKLmBVBve5/wHl2nqqDG
DJHGq8oLrLWtj7Srcz5Bv3Kesu6MbY+9tr7bUsTimNyHhaaa4LbpostYmiNergob
5FRYwBUaoHeNNc86LtJUlxnlrCQGcf0jLx/HtRa/hj6PO2CAt3CRoY7ejR08Jaiz
q58mqXd1q9y2W3yjHfnHrTj9LZygZI2RDZofVYKI6P1Jamzkp4SNREqmAoxjsWAJ
qrF9QI7Aq/uHd3ny6ZbnKdEI3L8JuG9nDNZyRNCHlR7SzE4xSME5m7Q5AVwxdrqV
RR2V/PcjCSn3Uv1x/4sGGTrUQLQWP8rDdil/CccwWZWs6jXFFhjQMBYEjl0yRQvh
lQeJWTjv5oKk7jVXwCWUfWqkIhy/CGYzp/yW7jiCXCBv5iZ0dj4QPe1nn3E0cplX
MP9fQDlXSQoQw4nlzvpyhlaA5IpJT7m9kLwHfRW94Q9WRpO8IXo2pyRb52HCGpjG
+AM3Q/mWZJbR5AecdxX/A28X6C/AgaGHQlpaW0w7MCtoIPShkzPK5Ap01t6t5jZb
r8eq6ikg5C8sptySDnMqgqHjtkGByJ1ek9Rh27+lbAZ8brwejUB4hqAneou5ZomO
jSHlaMizrgjqtif+jCfRAR1JqlSJg7Ts0umgEBDYtNQe8DXwcXnATs4o2Mq60FGq
XEWCaG6XhgxnUd1BFJ/DG8e+FX2welNE21OKaffpAW8BaD1hoNQtKM4lvgLCnbz0
603nPXffQEzsifFW2lz+Aw8bKcnqNDpd2Mp8VNnWmdwL17mzgzZ4yRdHRzi4JLJt
hYRcUiKZDTK0T8SJcjf/ITbV7GeSFWYu5xCSDWX4jmonjncDFNrJG8wP7ZfjoZs7
CTTxRIbxKmq5U/kzq9PXwHt5sRIz0bL7C9ZxqyWOnK7XgiXn+SwAzOy2/AP+YGBG
sRpfWriK8EIPVolOMqCtJ6Zm6mZze1J8q9kvUG38l6hUHdeV85FsX0N0p6GSAZKR
8Qg6tEai98KeDOWIxcqvoQkPUDZhfZk+xBe48FcSRzLPAEApyDUeuQ0tvrnI312t
mT61EzBBQGE8uXY3tY0GHyyER4NaY/v2E+cZkB6AOgrOywOyT8lsa9zSgQDkPh+o
uUmNgCK/9KjiyyejcmJaraptnrbeou2gzgvyb/3hFbahE1FAY2dghuQUtdZBj26h
BU0xzxa6fDLx+FX7ulbJ00pUf9aqq31CAcvrkl6QWuqn+B7tlEAoaTOedogSo9P0
zf40lbXw/uyJLjh/YLVrBz/wtCfNCzGY8zLzAHVHTNHxG6Eu9vFX6sZu5+S+XFgv
0TJaOVOsDRzpeKnv/aCVmQRVscU7O9nEtr7CFJFEfLOMDWLUMbePdgiVmLZzp1k4
KOVy7Apa69QIQCiD6yE317TtIyYCnKMVtu5DRCIwkqMlXhcUFJUtXmxjZH8X1vnP
X4ZpX4hM9GF1MOwbMRP9Tlnz4Q9k6nRQ2siOQaanPv3yqUThyB/H2R3lIjTmSlQd
DNfOWemyUyukXVTTY1rDGMeMBgLV4n4AUvMaTtm8rUCA8eBUV4UAE/3GQuEw1Hz6
n/w6ShNpkWn3DEEWhySSU3/MHLZ7JgowiFSj2BSnYiHLMgfFrdlcAgmiioD0cryu
D0zF3N3EJD179r+swcrJNOU0CEpHs1fwyrxEdFwZn4f5DBr1rqZCPgWKRpX/Wtiz
+Tmc93kNRMHmUsLDIYfvkx8a9RyKcI+sjzIqqQPjhv6LD0XD9H9SPsii03HKq1nu
yecELDEJfcFDp4EKuwd1dmh8Md88VQDwHyl7C30DXAQJZaKZoKPxnA4RZzxc3HwI
HcWRQ8Hf289bl2nGLTqog6X/7IREltyq75aT95F49F94yt//PuTfiP7tF7RhEukA
81mMJCnACVtUdegKui8gRrIzUNu0YI9MNjvvEn2sA6IH/wk9qptU/cwwjF40KAn1
RV8F4OMBVbehn0zChRJzlc9L5KJ2tts05t8ptqtfsQKXt+6KOd4HV/y5T9HRs9Am
Bkva1VlAtIuVZdg1g/dR0jEvcpsLVbAmxPARioalkqHp9O3vM9Go4VcI9easYMdl
NstMZOOUb6theXAGXyMt77n+K2F8LF+c1X/rynyAPqppbyGp+8/JIaS4cGBl7xfZ
bjl+10MH+hpNQjtbaNkySnh0QPmSh4gTv5N1btl/2XT+uf5BX5AUts+fyw8m8EWq
zIYFs6ZZMz5XambJkDBOrUFrmEhvhRyoo+SB45bvFQZ4JBSoI56XbwW6daru8ieU
HaRs3TsS0I3RwdPtseQemMsZNfsCb1m08oqIkOYlBvVd1J5zIz9cCMyjU11Mxx15
g2rnjfgjRK26LTa6BqFjTPvCuQK0LIWsYtBXttNQzfFrHI8XCGWA/PkjLTTVLxNI
4rqpqf/GKAVcL1oLrc3JfSrRGo7QTzRyQJrRoKfQGQAidhK40je8H/tvKfO1Ok1q
n3Cq5306cxA93PW8fg+Ws1b9RPt1V89SFGXXChx6EWlxMX/sNORUS4ak6VLpdbwi
qBf6dhVNsPuLHfMPi+G5jViCyFd76awVrPK3a7NVTR0B5a/EapNGqu57UMsT5PwE
javMzHfaJCep48wIWQrnPPXlqYa2rOpBIr+rhvGAi2/Fevya01tXqM9pRuwOzdLv
62jxq/ovitGOVAuO2MUZsrnE8Td/M44zf+01x4+MXJ8Jhqupw3hWP8Z/vYAm+G+q
vUlAunyJfK0ExWBUsQ1gttuXbrKh0hQJJ12631GsscDRckGImGzKpPpGP3hRzdMe
zhyIZXhu26ycMDb5djEYdrWmbQrnj5582uHa6dJ11s7aUeigIyuFSyeR43yzxruX
cF2oDv4ZAUUq2or1STena6a33YTITNkFdJeNgay7KXSu7ddXC9vBDdT9NFtOpREy
EFGCPIgEIQBvUpfjIFPm9S0Bylvf8Tw+n3c74ZUTna9OlHbcmHWM8XI07Z4iTerb
K7lK6U1A1cH8Hcbw2I3BFNMBddD/Nm6ulDIC91IIwZch0eiW0NoX/BZu8CPrHW+P
UD0pm/KLoiT2AlNdGWSQTIoaNI8eVU1iXOSaKo1zRflPR/xAXz+X7/5zEmREz6l/
gNYf/5Ez4BZpaj7jcq2mBZeBOAF7M4JRUvL9fihjKbAfo5Y9AiNp3JTNJsEyYLRT
k35hVJYI+tRnVKQbBaS0CPrugXpAV9pNCVh8HgNKqoiH8Z9n3fha4Ly3vi0yE+32
6RgLl7DU/ErXgUcWuxEGdTNQ+gSAX3kazpJ4XKZzFcoDGLZGtoWpJP2LhZcSF1Hg
jdyMrVxpGBT21u/9vt3azVDinmd1NMKFCL9B+Ld7HQXBesgyoClFn3AApgwo3++A
ttVAMEb98EJghVYNeriYxG1zIfZKku8Xk6c95IPrAz/+EL5AOKWRIllk3w6R0f4B
CxWHxRR1xMU6Fbp0rrdnToOlf8Y6JAn5GIiF6QxP3BsfwTKDbLhec8R843ozm0xk
szL0CNaxEkzxD+SU2+XXvadR872xKQpWCNV6ivHRzoPQGGOrRwjziQ4aaqNRV11k
hIS5yNaKiajupHV3eIZ2zSRxJ34sy3my0BAcv6foy6wxLZr3RU8OErlwfqwp+uuH
YDseCR80+xN6vvDLtrx6gaM9Wf/X+C7MelBpGCxnBUc53VMQZ+yYLll9feTyHUiM
8SGfF101gmSPYe+nbdTcZxK/VHIwcHIDLPajpOWKoRna7ZvLA67gnIUi0pxwAk3u
FCmQnrWrjgVSKmUY0IFh/mvO04mXpEw2pfh1JK0QrFHeaszX71db5kNUJN0SLlOE
eHTX++L3PnM4CUYaXfSL3BQj1SDF4QQKnHvP6cmVc2gkTmKNrL/Vzpr1gniTtr8R
YroDF4TGuhl+EesAdvAkLAeEJtWrsDPmVf+VLRTXmab96sGiSU5tAyzDSx5uQmMj
nwaEyApZRXuaxzuDOacJQ5ePmmwYgJH+5pkiKkD+NZ3TxmqBfoHPc5ealpp89oVE
ull97UBWfSE362TdNuuFv0+A5TQSDREFmzlTFJqaXsZ498MRD+U9AP/ZJs9nxJ8e
u113Myo+wVp6yTipSkDujbJGqdnWUH57QQ13jMdivtqwI6xHc3/Pxinr8esWhDi6
bkETSUhjB1eMwIeTXxm9vZjKVl7WK8kA99rR2bFUJmQ3DXuf6koPK5R6kk3Xy5iE
htxQJaIgZM1Q5LUxKJ0b9qQq2I5trpndSxvDAPUJa9AZljH90iGAw3vO/I1KgHlP
uPyODydUAIVbUqNhxgSu0pilAHOJyjkS4p5+tbiG4/TuJeBB2C4hx9AKpjyTvQzM
p8ZOlU+nM3sgOWxqY65vY7EuK5dNqXfPBoWdwIyKg+ClmIeh0lNmfXN1B9AGmELJ
+Zf/PgFDjLe5wgbJltypY1YFpw1RNtpajf22YTbUxwfPSyupQF0HRnpvTz27ocKC
8VMxIDcAEkJgE5yGRMw3Rudzyutg1SROxt+itkMaavdePRk3440quJU+vbInvhYv
UJX8Fzg92RyF4HaEwqurpp+4YLvrue/+8WAcpAaYYvEpnc+La8uVjtrE8OdB2Hb0
KL1SB2wc0EKJU2sAFJm9dXPZsvOqJb9cGS7kGIROwCe9eux2we5OCKuaJwqOf5ba
8tZMV15ERVDN1Cyi9n2khiUYbUXzTkVgF/q+IytQ7Fkl+pxsvQtqwk/IIAHdPMTl
0kijuuw80vCXJdwnE/QFYYVz4Nw0OKZl42ts7wUVivgVGeQJKzT+eEkGEFjJHZvd
/8BzHww9tUOeJ6SWM9NJNrEgGGSPdTTzJhXWtVQuEoJcKLg1wWapU1awbPHz6qwI
XedH3bU3zrACQRIgXzCkiOmTGXf0qgTHMX3uSKsRjiCNDcp7q6DsK2qDzPEKZiWL
0Zw2T4Q2apuRdjutu0BdmrJmaVPQvk7ILlgxDDJ5uMpZUOAbAFIanvVVaSgzVhvc
oh9gV2qab9ptlwMGrClPPMYB0y5Pw3orRTJxcY51KiyikWzT9r0wWwyoCsdAaltc
svJC2zbUWs1EmrJvUVe3pL8MB6waQBdVcXPQOvFd52o31Hn3OaPxqmqtdyba9R9r
HF4LBoAgeW8oyuzBmnMk++zyvukKDUR54iNLAKka6VeHbxPbl2pNF/LjQLrAoJ9e
BYRX9SBFK8Oobi8W9wP6y6maknzrlM80/7tnXnrd1fbUSaAMtJbRmOSoojCGsJi1
M2Znd5EjbM5xlKrG9NESdRnCQOlqkki433/LKuw+2Nia9kQ4i4nuUP+87OVw+44s
dkGRGPd/y9QIglRhmtvDBuJPaUcjzSZaCFMYSc2Ps+/C0KlltG9Z0SpT0bAFjw0k
lFGCKHlCQaIyBioltCPElwn8+QVnFvogvo1uHdp7DnEoBWm/jdOsuZGsw0FeoS1X
zO4z1ZHbVGdZJ5a7ISUGxj4ZZqg+W5/9omv88dIssL36rz+UAMKdvhSqkjzBG5U1
30eJJMez6RZ6PXU1TzsO6ELTKqH2tRgsfMlFmGIVWuk9APFKpX08mMe7p0b7xtjH
bjmjEn5Csl7E2lvC2mGHKZUjHEUn5JvQ6NqSwE6HtcucAsRrjm/TLKTjZEv7Wodd
plIpB5QQiW3EFUjThkA1kzz4INX6j+6G4nnwgHe8Dh/dW/lnnccnHl4p9s1fGq1N
XwQxJxiBtUW+dKLeBfWKeQlXTmzW6QRkTbri52TErw8a90T3uA2JQLxhh0M6WW8m
U3Pbe5hySRW/A88UIaWAiQhuvg/GmKzxm9dsrzuKlYSaHtSHlPCm5qpFUU7Y45qN
4eBKmWcjGyKb0ZaRaa6nPSIyO+02smjQfNb7WNE5QTHRfMD5eF4XkXnE6vOKpfry
F8VbXZhAdi/Wti8ZlcU1FZeYPVnu+x0B+FneuDpwPiJPL0JpNJNZLaWn0KHk3zQ0
5Ku5EX5byIjrGDsJeqpmHNKCyFg5YPzFZzGHdHm+aVBq0sM8ICZHDzTcOq8Wmt3+
HZAbD/3W8SzRIi6L2/AdI0l452bXXz31A6Wb3YgmxX5v2U9miANYIdACLTpsspht
e1JcCoS+iCAqKHD7tBA8i5N8GlfJrAsXnRZwzHP42CD8MJHiF2dkw4hJwYUHvuSU
MjXe8nYCwGqCskKWrNrz9IytQ5i38iQrTXzTeX39lYy3tv0mEQfhE4BvQ2hj1P3c
LejTWBjCpPqd+heSo1WzrkV2THKkBogbZtO5C8vFFbUPpXx1+b3PYq6BswGL2WxZ
oSsdSBitW9dI6TID3EPjcsguzS859iBBbCN4OCnmH996nqJHvzeniqGrwVZ4pJev
4xzPl+k7VVAe4uZutpZuKLQcjUcyVoN5/R3pIPBzPctsY8N5MDEXI+ziJxDCb5Cs
UTkB0ydtJzDnlbdZxPeNXvFvbKFu/ay4y2S9jXhPe7C+MrBH807UhJzusK80MYCF
DEWlPqHofdhalxMJFEvmWrQaOe9RxpXwz0PN7VOeweycgYDA3eI/ODR9TMUyV2f8
qsT3dep0w85TYRtMVnDNHL9s5NHsM75uiwPO5I6KJHvXltXwZu58UMyMLoNkfjqq
YnSC98UmQhDnBE7Ya+H97ROiZGhFkyUBNMY7CzUW8UZSv2Q2SL7qRxKyQRV/Hmbj
7wMTjzKBtKTLDWMeYIB7hSXrsF4fAlvVld37KwctErkhp1ljdDWYYs7l4BeGTS78
A75nzcJ0MScIX0MCFzHjtOSQj0p5kCaeoiVaPzwxV23cwDykjO4Dg1UZgrsBEkuB
1wanyU+9RMkrXe1P2mFgk/DbXjJxUdgJN5G8EQOAZUrj5DVJ0hhnEq2xwfRdzw70
4jvIFZnKsX95DDlr22xid4cP6MAXeP41T1SwIDF21RSgY5rWt4nZfVNnQn22DSUv
gLmFTgSFR1CyAE6IjkN99JWVVFd+MM5x2rhUDFBY0KgQ10YWbf2q51QO+jYuq6Xl
o7THF2qc4mdTsh3PznossCLUhob8x47tFxu9TrRzQ1fM4487TEUvMHajqcNpizAI
VzTSHMu8oJ5sx8s4YmRvbwlFcrDjVcNXnvthggsVRD91HzJ46H5HiuOoSpXEnMJ+
vzRcGIsnAntZEPDCuW9NeDcg3bE2K3vxxDZnLCER3vWKZKgL84x//dRh7lCUUWRF
D1PjPYyRJFJDx/kg5V6oFYfQO1cuFFF6Xi12WJHXGANpTnVeYBX5TYHLszNArooV
GHKX5cfwdvjQa6H2mtFksnw7p6ZZSVA3oCnsYhD/GntQR7VT8TBkiAZcc+JYTSe2
sJoVKeaxPIRS3xEDXYOKxZBGoEGAlPWck/tIVaZyaunBDmIxue9OxPQ8yCACxE8K
ExgVIBbtNsTYxLnALNUvWHtvPFtX7leO+Ka2P5rArrf81mJVz7NcXwefW5uXJjGf
De+K4ui7QUOAivcdccaHF920FfuLsVp17AejqK7bkxB25F+BWz926oG3W+dBjdc1
GAb/NC7Bj5ac9VpAzahdYcBXWsjPWCsngdzuPhcUehfV3qM/ogRmPixJ8PHOpT9k
fURjw32FjaJMq1s8525GlKtea6/QjuY5GYwQssG+t0Shtmxt0kEW0KoZ6zdC/6OE
IBsGBJ9NhQzJmEtCigOT30ElNisabmdJi+GZeVW9cYpF60/zSpKVaU/96cC+oQ0X
maXoOR3PgcUmJY/J5eujPuIVo4yaAUTUubUZ5wayZXqzcVKiUzpkZJN++nA31ihM
u9tqK9TH6BZwkcr9k/fjpA1pGHrPS9V912zGhWd6HDsck0njvELXuiYzrV1d5mg/
9cHFieSB7nunq/NTIJnbKHx3VEtkCZBgOVZ4V1TO46q0J7Sy4PDHBU82EKw4CDic
9CbHsmU9DrGLHmFqXhV6IWZfoUgC7nMat2QaZIfNu/qftM09RftotVxv+xG9Y16T
ATWBpMvd0NabDG21ifgiD0LKpGWWZEiTH6FCKqZFER0sM+xjjNvevMQ/XH8JZSjK
1Va4ZZ/nSrYr7PR53gF1we0fFda7sOZWJ0purIAqUpYJLbJk+NF/eNC36HSmmqwv
jLVR0XDgO8TN5eI33JH//G7jMplcp58Zc87oL27DvopeoWyYdBJNqHVzgjWkmHi+
hRNvFYiXmF4mBFvjUkwM1lMLEpxsvAFIcQbL1LKZZTajWBTlTYYGhxPY50Sqv/Je
kWthGp2URhqWfcN5kfrnWJduuSP0bMu77zqzMHmuTb6AYFIsvxpN6G0wBmwd8Yi0
86Be1KL/A7P2IyxfhfjUuVZgPBA3ZqKvQpFfYyExwqmubfpCts0TAslHLqu53rvj
64AeqedaNSOCAZBrL6atxN/U2gDP2ERmWODWfMOOueGAirestRQIXH53JReaNokP
0Z9Nld32pWdLAWfVywLWhT2/ufERKlnDHsUkqHvJ5VGZ0b2I9ihvx17B2vGzsE9R
6abFjrtNWJr8vsH1e08IEx7TnIzxDVbnu5osgG5+4FH6m96Mgl9709VjD+ZZLOsn
5iT9efPtm3scx8l/yPoDUqYQXCtrYkPktWNNXygxx3X4DThH/3teVcfgKddALUgX
5lx/wdF03sThF7Y4kihHEvaqZjR+Q3IWa1pBloWk1eeeqQ61Sy/cRneVLZQMPH9T
5ygDjZ1+wJySkTvKI2F4zFRpPxIfJRWfIXN/Xp+2icFLMchV7bxIF6R/t4qPtz0i
z/JD7ziamaMUnXx5NPUjrVwt4kbio62Eyi9sT+/Q5s/7GFo36JUMc/El+1A0/AOR
m8jK6uMK6gVI7Y11UIwI+msBeaFM2Qjkn6VrY905U2n/BCsfSEqD1hWTvFv0ikM1
dT4K7uZt2pBeeGIP8QXIcQ2OnBWE5xz1rcNECEtlCNVDs+8kmOOTCr1fIo7W+1HN
niNXtCiGEVPtMENBWcuHbeHXe3NC1KRJQpvPasX+9TRfJt9JtljhVOnv/MhvQ/Cx
PtAdtQTUwXaT2x5l1BdNdKsLEduPGje8Fr4F1Uwg7r2xqcv6z/9pd3otoZ1zUAYr
HDoJFfmsVLx0/izaL5deFf0GKiSDf4Tfn+HmoJPnWC8euSVjefGvNHdCFHDF7pAn
MdHeAotUNWMcCvNaskFf+oTBFD9m9Jfm9OXbDbP8PIwOC+b5AnmKaFprW+stADOa
aHIHXLwPHeaZqfli51J4B/3UzwTzUC+KeBRDp6eYNrdMuQs673f1Q7TSlOqK5fk+
7HSld1mCysaeYVlB14tGKBrEsov6yoyo2z7qkoj0DQ6apiPk4cyirhSQ4SyqDkYe
Bk+TSaRMohXDcT23Z0doyOkeRw/Fmh+85nVwnAg9Qsh41zGt3rq83KQ0m7X3QhGu
EyMy7ykOOGq+pOLwdG2ZNUJfY16sKnIBZrddKeTgaFq3UXFGCukmYuVNACAYs6IY
+jDXGz2NkxARk8u02uGe4gq+8jK7vn8xY+Vi7mMlDJYbDF/aQ/fAC/AAaKvg8UUy
WLUUx2YjffCUwZU6aSOyXr0AimvRdKusHgsGtUvD1CcSbAu7tJiPHFk9C04QmL8w
TvhMtX7VzeBXf3jYCP2Aun24rNlwU/dQNSa+y+2LTCuE4fsUrf5j0dXEYsAspWbl
rLFQrNzfH7yV841FH4hOb1b02F+OUZikDEiouV2+de0XfYWncGHdqdo2SEqrx7zA
Dhbaz1kxN3E8RgEsxIjiqh9ory2ozf2jhdaWjcW48pjoYbs6DcQrlJJSPk0idhnz
9THAwRXhMhGmdbBNubvpYfdvD9g31cR5AfHBM4RY8xestHR/ZZJlS7BisoNXQqHJ
PMu3kPEb9BF4MKHprGyeIj1kWl67JjiEnSBi3p7mQTzKd5hTxRo7vviFh7Qa0HCT
upjJD7GwmVef6VheTUv4riGgH6wA4b0sezwZ95prevY3uOAooKTK2JcNwVsVI6MC
WsXrCeZ/p84oZfwPmH+mGhFq8FzZhFXiY4fSVkajI53Zb2R4CC/H20xySRAYD2JI
2Ny4sSAWervBwEiOtE1OaZ5+pscPZelfu03zE54cgsp2UvoSvVv9UT0Uy2PuIOPB
WqWP25n8sJFTiDYBoNiAR3TtYtzBEL8dLuzLEf4S18m+t5nwTJsWm0hlybLz0vsM
UGRmDEZ0qXcGkGrM7XpDQP4Q3b6Dmmf09be2jugOcz/ppj/S6Q6+qeMHHk5enR2k
Fd+yfWFpTHjuM4y2fiWxqcgjA4IPSbpahWak78RxEX7LRpAiO2riKzRWDp98mMWT
S/fT2R3B7C6rSfwDuXRgqTgouyZECDcPerbILSvx9nLarO4UqZjr+Kw8QI8MGlq8
nHXlKC2M33HgD/5hxRUNiYu5j2KtFrXYeu0emdDfREvfJ3zGrGxapR2Qm50IdZeL
60Xwpip4Ka3c+q8Xto51nXsby1nlXMf/YS6PH1YK5BQhKEphFfy7uxlwQ49anF2D
3rvVZZHpR9r+JebEksmrfgC7VX8kCaPD14b6X7VDEq0st/SPrtEjqeANrYPV4TVZ
jmPleuf2coXXI5RfgvBO8qB0nqkILz4cxZM5CFUI0TKaQrQUl/EpYgxWwTh0MKpf
hsenFMFkdmxytEf7HElM1u4mClJVPV1z6SlNWIMtryCyc56KNDIgwmuudZ7n6k7y
iqYPUpecZcGDCoMNlGewLkz3EslXFayeVHj55m9SYvFcypgqEyOASPwBzOR8iGz3
u8A/r9U5mJTeGyM1zAONj7voJMzS33wuU9I/jh+yozN4+IgWtTiSfx1yyfHsT5GX
oMQkn1aINBq9X+ml2CKJld2NCXwyery5ZpzUOL3dsSpkgQ4VF0sHlGYT1PFiuTBg
76I9d6dfN36ut9ZK6sP13hSyf3pAg30TatkngJKtED5BCZkSxe5VobyGI4L5GOzi
O/b8uFRsFSdSL//8Rsr0pVz87KYvRHWGtGWAHGm2G6wz9XhkH7LSPFToGVSd6QuW
0siWzMklWiy1BTZWxEVbuc561QjGiqeDt20iI5AE4cG51057j+TDjhkVv+720egx
TPcMilqJPPdkHMxz1WRFAu54jZXnPa6O2Xf4WpUG63+W5z73e4TRah7AyEvDz9jg
T+6f7dIqExut84O/TLKRnaBz+Q2EHeIYPkU01BexLG9XJpn+XWHacrhn+6Lfss/e
kjbI1JfHen+pT3NgnFSLrylYc50PLwVHjRB63VF0V260EqJCkDPiLA9vwrwh5Qg1
OQ2MuX1mBcoNBiHIoR0uOB0fR2srPDU2dit6/zTW1pa4wSIdOfsYxzsNDZsYlrA7
ktCIViz3T6wmx1w7f8X5y1PWY8/dnaJ49X8zJXvriEuNPxiU+ofp3QuEBBomONYx
Lsr24ZyyfZVykYvpX1U2aiGR68UCzEzXbvQ7YyE5LyX79lUzHrNCyhtJn/egiwvq
touiCUDRSXpOFshsBpiY86hctefAGPAbsjd/wtOEZeTCvVS/L2mTe3sWPCJgN7kU
jD1i/Lb71OaSHKsYMiDOFk70YHP31S1BTxTpFwTFlMV9H9NzyfdYYbqGRhMpd6rb
6diapP7HZM+7YLbmpYNWWi+Jj4WRnrtC5dQtURmiSndaqo3owVM1pF1aJM1D1rew
AvMGS9A32wMAGWeWqViQC9p44jLN/76xz01CWhwepN0Axtzzf8uKUhr2rtSJT1ti
sblHD13Dqqp3FP2cJh/kHW7WH37V9y5nY1IsS8F5ENtNGbIO48+GBdv5Ejcxc293
KQWig50T0ZEXnEeBPMOCVdIkDE3Uhbrj6RX7itYNa2/7445t3i2QBPoVLlOouvQa
Mfa90rd9XgfWC/xOfPojLSVVaGkp5TKuwTs5mrRLNBGGNGUAEyqyp+9/r5Fg9xkT
Yakc02HvkTRsNDqI704oCqfWrHqdTxVblB939Q8J7kcn6GgjN0nSqfn3CmsjLdI3
td7STW/9jJOKwc4Etoyfh3Jk/WQvPs4TDz/KJ+ymPj+ZNam3cmcxn3j/I789qgRk
NAxTZLEQOYbV5oyTnFuSJbpjOBaWKi9CicpRCq6JbSk6Ono9CX6nqT8Iui4Qr7sB
O6QLK7MJ9sIesPODXp0H/5/J8Y7PiaQNe+nzceW/8WEAUFNWlFtwTeNXf65lQhll
aAMu/Zgw9pl/WlBYcQ1KpYhFDFgxVeU+MK10Mr62UTvnc5H0uupD/Ms4W8/Yt0L5
FT87evaOr1UPdKQNp5meU+y7TjtxrBwg6szunb2N7M5VGDjHQYWd8nOQgh9Zlyqj
ecK9UM6SEOOxE17MXJaQb3GPbCYFKWGrwTJHi0gQ/LWoaSH2z1untzoucdDCNJfc
IG0eF6hnGpG2C3t2KejlIhkxjL/2mgJkXnFc7OrE+SdXWXdWtN4wakNEURX/jg9D
YE6ZWTSvHgLf7e3W6qmG740RPpE+JKgbLwXSxmg0/DoNVQeB+RowvDIHlEgELDjV
RyYQF1cLT9uKZrP55CKd0d+16n4FUxPU6yLEEo6emE8Q6JBKsl0vHaS03x7EJtU5
XxOayoLrbsYZ8w0A15QlG8kZ/BmKZhZLsWcLMPK6sgstI8A15sMy+spb6dJT6bsV
OB4f/daloT+ywosstWQqEXkIODeHqVN0YYUiRk17A1yaKTV9JyZD7f0B0E5xuh0m
wkKcdQAZsDs2munOjGqkAanHFWmRIPk0/uOo29eYSQ6OqUeMVQOHEgm5YCHx9+pA
u76ozyY4+FON9kRbeCGGrrgIU8FF7y/RkZu1+uQLyMWCQWvf9U9me1uVD4a7iCWC
VkA8paxxoRehi2VhB5rLDVLwAMuTBocWpQilJH3k/swuAipR+4TCItV27W772Z0O
9w97FfbwUzS/D0u7lIobp2bLgqpUaGBGu9df+s1Nk6oWSb65CSYNnARSW1M0K55D
VJSghJVyvKiNiWS4oXzwVp/xiCql+bXDsev9sw5xIfL6DyKdXmSjtsVYmaUHLrNl
Ej++B9cdsICzfA/gT/I3n8LzApwDB3beWa1d81jf72MCnCoJS7Q7zJcPTjYFh1U5
RrEwIil1irTxw9AbRXIyEK678FqkOk9clI9hCceDwitmN8NXRBbimVy3gJYc9bsG
o7sBj5pllGLLSNCPGV6Q8fJc2kJfloBlfu8cV8k3UYBR8YsgY1m5NSLZMJEPOHZL
JtMbI/sXQcIi0WMj86rPi5KWKsto6FxRjh32X4xWmS983q4rO4UYhl+hXCMSj7V+
HNk5fPjKTNFa/xwRjluuVRuc8L3IwQROVV//Mw53+2e+zavNS+vLqnEuxklYTHJp
nUljANrHaEfqJx9aFWw1h2gW+5IOCrP0XVWmn79WPi644tw+CE2syotPEkgmqtUO
D7caFrBGddr+lpkYW0sVFLWLiakA6SnxKilE8X93HhXeW9HUQOmi82dnjZ2FAIId
uLKfZEbWm335K2XLokYEJlbQ2bv6d/T+Tdx/pni6HPZo+Jokoox/KdIueK6zdiGx
iVSyfomc16Caxy5JmZGx9i4l28zN4rUtU0NhmQCeRltEZgI+Us6YDRbQgMO69vYA
hS/yePocgAVSNmgrphuAhgZcDnSApoIxF228VFkRIhRMEFEFzdG0uOWexSwqxJoS
CCv51Oi4Cs2Teo2lyI5Nz7QVauxOHGbBBUryk0BfSvvuZA9lnM8wxSqgGHwr5xPz
ssRh+n0W8l0H3TEx9TKtdAFX6Rk9KYjqD2RuNXLJGRe20usYKkVvG9JbHAKrrFaF
dnFq9lEdgwZsJk/2VF9nC4ckt+/8lvHFLgtVnOEELrClE7E5g3046J4I5XiRlDvj
ZCMNvA7N6mFuyGaHzi8fM8vZuQv9qONVtYH59cmlQzpSdgH+pJLcCSJ6xMh7NuVa
DiayahDUyBUsXxjtOlU2XbNJlGb+HmtdOZYJI2QavS+Qyy/rEA2dt0unofRy8/0y
r3iO5n7yLf0fKMHJTb1rRGVBN8jwghC9SDza8nPcrHvtQNt/TjnhVPSGX1JVEmmr
V4sqKtJ115GWDGjEYX2d61iPdsHBya9f52JhPlVlmSRykMCwBIQHmt/Fyz0R313h
booYbsgY2TjkBzxOLHKvVIKwdIRxZCf2GvxoE3A+g5Fnx1JY8jcSDhTubpSYv9nn
a55ECZhqh4h1iW2+el6JLAqJdhsdFGHMOUeYLnbiGsMcfD/CJ0ypOn9QQh10I37b
TiG/lb0eJP/KYfqqt95GXm2t9cxSiFlN/odnxr5adgXeqtZElVsrKo3MfS0UX7Bh
yeSsrI8yHqxc6lnOI7r9Jukg7XzXQ1yk0uqiGn4+1GC8puPtAJZWzbikzphy2d0G
OPy8v4YSAFcw4ArpBUYyjuK+ziB+YpYgoFpAoYL1fESigs3zD+oU712frTG8J+xE
UR+CjuxHjM1bn/esXBw0IB0gO0YWu8xLz0UhBK9pLpKpGlWFR3+8N7a8Mt987A5u
njWb6Tlob+CMRSQjmq+rY6aS5qxRbXIvazC1MGH82ksCfFO9fBslh+HPtONHZgXW
jI98SeD6Sj8BRr5OpvwOSyvXofLbyHObKCqJfA6FY0c4L7NABPzk0GjHoiS2xMnn
j4L2IKLU/YaSZ4anOP2ailhHoyKW/lP58W4yke7NUr2XPdf1WXhobgZ7qDXxrjWG
cMA9VBHbEzLobJfTiHhZg40AusafVEYu+4vZgIW3Gmf1zdKI43+x8zu0siJSRbn+
YpA9FNak922FONNuC/PcOyPGhnaRs8KLE4JTr6R2lNtuq7G86oBAA7/azCxI74Bq
tK+UhNe2U8N17FpFDzMwWcH8NmxYdcvp7DTPtYoxNvas6mEsXSJCMK+W5xBUxzfq
15LUq0kOqdY53PtkKl3qSrAOlbk4s6oDKznrAMzRpIqRufPV72l+26CR4wj9ZgrP
JLrGkd9TGNTMs43A7MLcrPZFK1WeaFaLdlDBZ1v3yF8z7l46YvhZMXwNrXAC1KiV
9s4+5pwEbLGPZPjHaOJutWEHxz9JrfChtR8tFBkz99+HrwDPcoyUGXSvDqQ70re/
IJ5GtEqdsVKBe6UZI2T4GMF1cM8QVbpQqZ5Rizye0mWT3FMR0M2yGsHHz6ZSMmAz
/Q+tGCYFWXIPRlEvV+Ye/Yscfe9nD8IGEP1CbMBwiUczlyCppTfosOWoz/SW8/NB
ZzWb8EqQhvBzeVWi/x4flBdHdfLvap2OTc57QhxNtLFCxQmm0g9S2J+8Ko/eVgwk
OQKITcqUgQBfMcPhbvUvMjwSjlnFZ+qKuR6wxjW/+dV6Ehzw52mOA/iB7ZUACL+4
zBsdCDSIplMfbGLGv2bIZdy9R7GXvY5j4HEt2aiEcPQoI7jZyMTB+dDim/LFaBlW
I/HMoXi/vhx7e3UUpLU41uAbSNGPXi1DnwDFmdtQHWZEo+yaXHAc9X0xn44T2GRX
kUI8qk8nGTGqDPIlbw7PIovxQKsNMI8jUx5lX2SqTpkUUJqBp+RVGRR0F5tsIvpL
aV0BeWSj9Wh1Hj/oeAON4tHU19EBz7EI5oQuxCHDgCMF4ebHFTyDs16JTcxQ51zM
7E7tiL5/2K+AaaGUKm+Q7lf4tZy2WWKRk4Ab1NJJ8BVijwTRPX2fmlS/vmA9Cz/H
L8nJQK0dhiw6PYwct2C3s1rJl2UQmyJvje1u+oaYbldYxx9s7M91Y8k+H7OSc+oZ
k/woxjqlHFMgloJzUxR2viEPZueq6UJurr5A8upJYPn6L19eR6od7p++zvobaT2+
HWwTWsu8tkeJ6L4hE3gi4ChgjZ30txl4OxJCGJCmb/iQUSm1xSeiFCc8T52HMVAs
ZV+fIx/E6C9nkVQtoVEeLwP7N1HWCeM61SBSR8CuroksiP+61N6PdlPxzSNPMrzC
5KevYa4AHEvv3uoNIlexYnl9SMtrAM53tASQtELKgFxzRDtUQdFRpXaDjCRHfRoR
06AUSXrlkMswXNGJ51epOkrRwZJXzmbBvfI/Q7HcTqFVywGtGCafNDI2Gk6PuOKl
IjFmN7CGq0IgW7dUaQePpUHp9uxAs8DtiHrStVMK4+UAwKzVRfEoDBbWg93YXAsC
zK0k6uSfX/kCRS+l12+ESoUc89ZuTbVDm5S3MjCl5XS9g890SihY0b5QlQYWYXJR
IkFp7bK4MUwp3eTluWOE88h3l1acBuk2uXphv20pp6Qh/mZJngcrpYhMDwXsu+kU
mjk0wLxPAiF794PdGiN/gVaVWQRdpGwyQ1T13iE0GdPgmPl46NsUtXfgCA7pUXC6
fHLkqIf+iVY2zKzZ8mgffCOXLyCOTFQQhlB9sCB9ddVyZP0+jRlaZmj9zzO61k2i
2YxcE8UoiIU2jyq6lCh6bbKMuVqjdirVnBpjj3kAQvkHnLa4xBTn4Z5UPxtL2ohq
4vXCu8ikUbHQzu3zN7JmQEsSz9b82yTxZ34m1dSIRkHAR540hLJxHgm0xdmk7jpe
kfbNCYNza57ijQrwc/hm5yfaLU7+gi//mRW/NE5LFEjtCQff4MDRghF4eE9MCXMJ
qxzfopmYLMXsxuqFPtWGLoPQCL0Z7DVxVzvDGTBSdu60kJMZ3pbMwTWKsuObqUC+
4g33uf5i5PmOFzYzYqcpX+0dZFPB4VXL6FQbWuoAWeSGcQhKbIiOi3pefXKE5wLG
7XkHnXsKL8L8XlwgrsV+oWFL1xyZvKvhpr6wQy5F1R1GqAG+pMH9LetfDoGNd5gx
LHNsghzkv+NdaID2ZIG5cKLBFlfPIRPuYty+0Dbw0yPy3VjdFGV3h1H5EWDxkB2F
nEP1p16nsWfKUwWi3RLbHXpJEK0ZMJYn5dJnoeT49EW6xmcIqnspBpn4dtlflgvi
ddOy1YrGk7nZCOwzdL3jf1pnIblNMSjssMOHUddgHIo0aCOzUE0S2b9eIPQj2/UB
Gpvl7a1OUzqiGU/D9bQhfg2AIKr8hC9RNOhPfjPnzBgm/QhptUKfpcvW0PUEX2Zi
eTCBkj2Dr7tdrxnMjOfSPTEqsuVChmMHPTOktVaYz477gUalGrqEHpql4a5S/WIK
0Rihm6yRmSiA3HlLf+TDQbk0B7iXThCw5mDgO/ih3wa8QTmwWpn02WR8PA1xY8b/
1F7+WGIIzdCK3vaHUu4Y7FVT7A6oTp0UFGZa+XQbd7bWuKBzJGZcIUcrmug67BCe
n0ACllgD/0NwIXUK7tqKLR/aQBvWVHqEhRJM65GzLTO1u589e3Qp/s9g9jOiyCo/
x9RU+Pr0cJ4vH5eRixdJuiNt8fVBMnVBAFyj9bLpWoHb9imDs/QSVttMxbxNWPnA
KbG/6NZ09iZHs8etAZik/uYhqUhO4oqI+PETyt/Dzlm2om4Ya4LsPZciqwL/a0l+
M0ds+TuTOMaVba043ej4iGIKDE+KH5wlFjK77ZnP6/swMWch7UcEHrkaQR7g+tzO
vHJgYRvUGlLymVFSpN+GX5xjA6YC6L6euKfdmM5V2K3pnfmHOOoQ3UrEZIhGov5f
DOeQWYs5VyHGMKw5+bnIHvJYMZF4mtqgtmdBnPViZUvPQi+G4DEMUG4CQYxuUs+x
FmslB4DK1u33hv1oPadmSPHhppCgrRAiqg4qVOgU7DQGpAH0Bgi/op7B6d2kxV+Z
gwhuv4+y/v9Tf/C4SyN66WedMy0qjihGwOiPkoKgVDvfX53ZObybWIaUXiWFPJK7
R8odWPGPbhFOXu6GR+LrR0os504+lsSHjPKMfqb4HnR5MyxW/jrJ2Xzz5sWDwNif
88KQaiOkzmy/FhsOsQOj1dIQbVV6+M2C4yqWubhOsRLbXzH94z6zsuLf8k+pBG+2
qoff9RMUYi161GfRW3YnqzJkGOPA2rIFvfzVJYMp3Ej5gxUPJ+KU3rJ9TkKnL06R
nNyQvtMuDabmXNMkMVdJQv/CJqUbofFLDq/h8qa9S4s1HcknIVkWbGK3Zko61LVd
1juLWPTbHTEoktpJZPINY4ua8iWV+tPAMFDSsXh3q7pci/I6XJDbXBOcl7tdXinb
rcvMnmUC7gYBVCsK/rgBKTTEkaOQ43qYGZ+9oAeoxB/gcWpKiPYwfnM+PzgqLmkk
Lbqp/LPTeTBpc+XzZMh/k/ETBujpsGp45SwSio5lBY9BKoANmGmuUR4m5lG1A3Fo
GcAoxlurZUCHhbxkJCB1M0iDh4YxUVkqxby2lQR373Txd2qj9JYUkTTtONlyiczo
aOHxYsBsgSesrC3qYEnJbxvBU+5XL9mY5uZE0BAXF9ee7QK/LHfUItSmEwLqL0WB
mthTc5Cw3NZN6h9kS/W+Shv+/pJFjXeAZjtCO2T2VC3ROY1HLlVHaDhS0tEtUqBx
XcTC+VnizE5DGX03zvgKKeCxtLDVVNCDQcTcrPbPNskdGou7elZxElFPtvZQB2TO
qZIzK8G0cb1LTNwiXy/OR9MyfYD8gwS6O9tASglhho5YJw5RXrr/9X0UVwmoaPrB
ypQRoPuVDb/7/3ee1MVF4TM5RywH24UsGGZolH9LQXC34qyMPv6vm72tFnE862lQ
fBgi7bgE2wrFawEVe3bQyB2rq9nEz1yPKT7xWjfgDOUYLVVFzpIdLpKsVvZsGzML
ZGLt8YHpDv6032XmjiZauFZKt7ALmThitpxa/+BAGq6x78PEGfAvovR9Cz9zJUrR
J79tL47uTQh5zCjW0gWfHjm/xOxVtVPSLRz57grwvUWV0vxR4DhT6G7ETYQxOXoJ
a4vON+cO4rQ0gOdEvx/mCUSN+pY2sCFeQXqcMgTvJW6otu8XEJH5E9zJ8ZEiQrZn
A9hfYv0loy1ft3zzUm6DaJpbgLclI6v994ST0uwOx7C/+kiPqui9VJfqgBn4EQez
6rdITyCe5AdOfj/90RYCmje2+2Jzgte5KKsKTG1k913/4hgmA7mD4SmSW6O7hUWC
kmO2pfRpJToiXJCfFInSxvZYoF0r3UqhVw21xdcy2g+3iZxSh7Trj8DGAjaSCjef
q9i5SaFUJhKTeHcH1Ursss31UCTDiTgxYqULQd32CeZn3byuHrmHCxOWsrJeo54P
Q3zgtoQYZcyw1pQV1C2y9nQhZuD4AKTP2gQoKx8jGpwG1AFlu6I8AyUy8Z1ZxCli
kdMeYbBrf5Y3MUubNQb+a1bwv+GCWIp1yESylrVDEJBLVmS8hqfGHFT9bHunEXX4
JDv6OE5exzhPVp5doKIJkXLVbMO/WsmgIlMnAQgYaUbX7n1Zwgq/Yjia/coiov+1
T/wOFmu4MCR9Ih87sHSnW0WpQDDr6enDWuIL1o8j9rL23MbrI6EFCxwCEvcFPDVr
GEWiAosgSQ0PZe1PmmoOZC7ULkOvKSMZg+BeAxHZdopxR3VAMg6UiLio25KmHkdd
BARnMynbyPeOwAjaYcY2HWqifrg/tt2kcdlCbXFuSGjwm2JKdz83H0HQggYMVxmC
B+Q1b97RiXzbEZhY1VQuJPdA1dmWMXostYOVWyh0iHpofZJaeslShYrZi9e4EBFp
eVMsLagylYaSNMHVNrGqgrgK4CrO5r6nfR4O/81ArMrfRYxhCOV/wSQqh9kr9v2H
xqQ09B6LGM7JGch5QXhOJmCAMfEz40RbIwmTISTxevz7j8fEaanHMPSx4D8pFQVR
FxpNKSOscXRW2PVic5qy7frC7XOH96Ak1T1i8Jc4/2muISvGx2pFM+ypTGJAdMht
s4nLx0RBbQuajgqscjq0soziA4gHOIf2mQwQ+aYnBsdoIYd4KgcmnW2JxDLBtByT
lZIEfBO3t3iV19+pXkp0nRdQZAVhm+EiX/6NO/2G874VevGsUdVxUgAxwqtKC8os
IjuTEKBnAOiM9eKHn2gIIAW7GJQp7NswMsAWyIeCT2VEzTtdg05TuVgU9vhCJMKv
O901gExYHHxGOw+3u6osWaN/QYWD4ATcc2a1cUi3tZiLqdb/L5KBGizCSQLijreW
0ih8pALB/TG9JKPL/2mbfAjSRZPUHOnRuUMljD0/OoN2vGN6fMPXVD7EIxVlOm8p
ywyAiPKXHtaqJo5dm9pC3Iy5kiFWwIXi//KJHqsYHI80LlpmrXQjQRM+paSyGyCG
e6smCF7ZC7Nj/V+Fnv93/IWZ2JczaYppflA5OFLcEbnNOsozDJVEtDaHL2a6KwtR
vewGcquvMX/rP6SELKqNWPZgQ8J4BWTCcZJ8tpKlG4s8ywTi2x6FjjWROE4mQ2Ow
qIbD5NvAx+wttPzlsYwm9vcKmp51rsU6bcw615GMEppxUUxBd+UAJQDMEU1etnzs
W5BfOc5l6+hzhIRSUjdzRKbeRa+y/hynzaEFJRSs/fN/2mvjSm9LN6nb+8l77K1b
wzTDHVDCAlh6RW6oVV0njiuFBom1u+7cVk/XzxXoNBm8qzp1Yld+8kqQq3VuSQZF
UKcYY3pSIrJkcza6IpFgcXOw04eLF6aLS/fTOVY4D+r7BNl2jY5b4mSc7i/0umQL
eZE/UyGbcO5R/IJviJUlL/0nLZGibVS+W+TlCwAFchmvlD9e72QmMGh48brQaM7x
6OoKrUNibHlpCOVb+1JRQG7EQw2A/5VE0rt53R5vC9STI8WbY9u8RcwyiH6CdKtN
RCXBSCBUvbwHe4BxA/j3s89w3QgxlQLvcHtjcyu4ifGz9dGEdZwZok8itoRxSTYU
DANgX0bKvGFccjwtw/6vme7uflLHvspYf6Dd1d+W2ofdboAzEhrvJjfJvVvKL05x
aIL2ujC8USISe+PQFCMVtrQZ3jPTKXVYzhUoGj8siDsUtzZPDAHCHnbVRVnn6VAv
8nZTUS7ngHFaJes5BBaW1VPke/o5pFEeXDyzp1HYtdTeoOpzUhGconBeMilQ8+Wf
QoAgd3PiyH8I0tbpva87bvXBJljHwK0GYHaKmaDlwTvmcwXvtBvtJ9m1ne6FPxV7
1ZWJ5FS5sLboQoCl4cN/5cGxLnB74Vfbx5v+jVnNEjHhjiDvxH1CU5G9Ous5F2kh
0aILv68qMN6h6v09dXO7lksWgrpHQbkavrJCxn35fPDDNgBoobWz9gRwR9tYJUiG
GjAhrQTWU2KKQxYtZnvH9O/uYhe2wdI/pbp0k/m0M6ivq1mvwytDWoY/6gxisCew
6yIJI7jRXaeDJK567hkotoSzz4A3hPVfgBaSkZpz/X/0ose2Vjp/c99L9F2zKQ0b
WOs9CwNKS7hXQo2yE6vmANXnuPpM6QswIKenCQn8eOj1LaEZIX9/4AYVDpTpr92E
WRBR745XrWqyDTCWgKUpsYwFuYIT0BtD0BnST+Y3BR1nQYLw972luxPVmTAhjMtr
/n7zNZV71FXvpQK5KLJEtSyvGe0+ZjuLEJ8B773YefJ/nCEFFujsMEUVK+Q1hsCW
F2YNvF7HlumSP3GK/wey4Weuf9pwiBmDa0hv9SbW9ycWskFnDWxDidldRo8LxWjR
7k7eoNdw0hE1/VE5x/yA/Y+KoTEIdckJ9PMIGYluD1BcM392rvjiQ70AYhpEkyxV
Y5ji1SWOGmSOG7sTF6AXJIbAgeDQXF4R9Ku1JfX3MyuMbzi3x2cpS+TtaV256baQ
0yIAzEHiZML6KlmFnSy4ra8v9ESbhxPGuMJWXSMlAo0FNVeSJ+o4hhOOCHztRJ4f
xvg0U6ZG9IO0ViFxnMFlohFbvu1CHPVmzBjZmNk8WsIZghsy/PTp5wnTySVBLcgy
ZERKl7cPhE4q9I7DzHRtM+bIY3C0FnL0rrZU7oXy7cKj+qSuGHYpdNP2xOxKB0Jp
FtbmbJkVnle6XFuOqYGPGmrpqzlxT4iuY7FxNs1MfUsC+7xIudeeqLjeSqfJOCBV
r9S8wqxT1v4jLzZUvwX78qrsg8P48k+jTfewAMrFpo3bUkABaWPfnhdLD33Aej9G
FasKXKxZ8cKb3e5fkPXBi27NrP5rZWhzJlQhEVphPB5KMsh/74hmc+jtQ5NWPRJG
4kQfJYQUWKOEu/+26yusjfAjkMh/9BPgRHzZT2ujjqyOU2S3dO/B+IELLaSqeNTP
61jmnnqX7TKRG+Ju3u5rs+QKGE7kCxUg2lwcuksfMFQY3jn9NSNth54lBMSP964P
92p5NXNhB8oqPToFG5HHJ5SQ4SilRuY921aURkqMHPcQlaU2JrZkVYSuFJFp4pWO
wJLHaa44M3Z02S8WlfVmgGmpil9c74qHqmrr//9gCr3EMGfsGmAigKZiqISHHLOV
PLfGocabU38JM6sD4kWTTSj/zDaIEVZpS5reqDNxROvMZCG0rhRVl3r31/uGgcsI
npl3aP1hjDJzp/n0a8AISg+VaqfKYTgtnVyNB8ZP2AgZTlBYFsZhPDQhYHd1ST9A
qy31YqknapXTr+wtUxIYy0jnf+TntiuqSIfpdIip8LiFWGpvlp2zpW0j2trXvppH
SqCcMz3AUOu2AC2z/Rm57D1FXRNKtSNOfTwJaY6XUp4FCy6Mdrfvk54ObYi+HnsR
Y31fv0PBROwx61YQrOFPmG9Fd038FiEAx22LxP8774SYLXHZchXRXt6oeuJ19tFO
+ZSMcYq2SeXa8lRHEUB3sSrm7JjFTPNaVWAVwhk9o3b6M8UbnyghhujjzlGB14mz
GPMZ14x1Iz6BH7bfJJToL3d0qhTBpfWiT2GxOApwC/V/8jrIU/d4XWAxL0udV/Ux
69Psd11byCM36uN2Xwnm9lutfVejby3kXsPXOSjZpmwDiy6Kx9Gxob2Ut3Zwl79y
Y42ovOqNe6dpyYDCuvEZftz0zAs0ZCB7z83ddEPZpp5qejc6dE7KPMwfempKGvqg
kYoo0rwi511g7ioUwpXY6jZxnqxUVTduedi28iR9anmOwrzRetwSUvSTZ9T6u2Zt
DSeXju3OwFt8s1SquQWcD88PjRhxQRImjNPR55w79J6ILf8A3RJphZVoWt+ogle6
M0t/B4+3nRWz2Cj7/eJatXq+jBWPo+w1J1T3f/M5Sl6SetXLD2pIoo/F28UwhE3D
Q0osaIODfQbSOg4tizGcoQh3jorEe215WOmWMd4Q5HmbSRAnAfSgkiy9thB/TKVy
Z8sT95sQjh7usKinf29cdDLO/hXu6c8B4OtulO6YsTTa4eNOmz/GZXTVSiiEa6Yc
XmIyvQNrLYqds2xViKtyyysPiDcZNNbzwytgBCsr58wg/eGQaaS5ut07Vre1Q9Kg
XYS+FfMuubrTdThXp1zoevCz6JIYtgBEx5WRsNIVsEgCQfjij0qqzAFCEjCL/hLJ
GUzrgYGb5kKL2tNsOh535KumOyguRiLieLNmG7vP30xPHec8dxV2oApE1jHE4uSc
eZ7ha1N+pET14VJsdiXSJWFcnGlXV38/kyMrNeg7DHlzdTDmQ9xcsAbBMXGDL1yA
DlIhs1J5TCfKzGOjWX2K7ez/LhjB6rijEOBhMWNes+Mb4DnHRww17I3g0uHqmu2w
oU7O7BUSNgFMsC6m2f2XTj5FhDRGwv+8ctdi0g0Ms3hUPytxB2JySv5lk5qLz8kg
ahmz12UtDx//E25OgJzcl1CxHHfmnM21/gfwoACfFqSymJ31FKZr3tPcASCbG1/5
zaxvG4pczM47lgPZiPfAuSbP0AkAWwYEltLy8WDYNXsK1T7TZj87n0KAddFzK11F
bHI45lauh0HA+wIswOprs+j4c5i46eLFSBbLhhyNiTPidWXgvin/0/3Mat336PqP
rYJWeIZJX/58f7tnW8PSWKSYzStO/ZUjstDv2a6szsdeO6Ncnmwh8pn0Q6YYGyOE
6Ihu4gY5KOLdRkHnop1a3h1ACh2gEFhz8jC+0G6KENH5PTJdYZhni+BXHvnKdwjN
rjaOtIX8qq0i0a17rYP5I+/vxphRxCHoTe4mRHe+HoIF9M3vZL2gaCdWnP5pcxxQ
1L8tWuxicj6saQ2AtNL+n+NeleSUec5qZq1hLm1Yvgr/xTL44dZRbngsJYS67X7i
/ZxNFdUmxOMVUnG6bLgbca31aD6FwPDldM4OYV/KraQ+zPtysB8x1mlaFA8JVPsT
6ndQuzFRRRr/kBIJLFb+Zr0jT+yQlNwWXQku8bxcIHikvS2LCxWqzT5APraicI6l
IsVQdEpFBvsS+hfxyqdljEUeVv7/JabctAFOdFXW1X936cKs/CHisoIgBCsB91sV
jtiTKEkqoTL22d7UyiE7iEcLDtvILCQfyHsg1BIcoKvTQlvrEoryoqs+FCK6CqRK
XmjhCZuaHtO1U04LIhCOXJ8nptlAznTuNhxB17FnZzNM5pUd0xH/3qKRg6eEozoO
gEtDGpA/hYbRPa4AGR377QF4/klpd3Opx946dKErEWBM0z0HG8TxmBHfr3h76Nnv
2pIlZDiIiScwfCJefuIjHvFqQJ0efTST6nDt9CecqWb5fdVw7M1NSqEZqG2M4ULg
id1lmsCtg3n0Vb6FT4iEdrRPvZnyIYJLTuHVtKwCmj8vzsdBO9trQqTEcvGb8NL0
QjEvIP/NLXMBL9tpBpcY4T8zDF5YShcSNUPwYtn2Xh0Bh2KpLWd0LN9LTjGThnzv
9EMXkbuxy+f8+//pV0TkpnstEJuoHf7jD72aehHQv19dBlHFUvaUR7no2y4fum5k
LNmZst6HO9JaxnUcdtLH938T0m4iZSX4vHcM3kEaQnhirpAY51AZJJIInl0NFQKm
cPNsixV/tDfIUH84KPLMx15dkgZZkMmb0oMIB8S/PaA7yX1N0FTC7rmNUPXAJ3rM
g7LarzaL2Qju4oFZznj38LV7KKT1XU3QPRFpNrinr+WovAw7SCg839ZIJ0N+U3li
dVCIoU26hRiVXNgCmxqTwG9DvLYscI6/aRScU3oxoAwbBKJfqnbKQK3iCbS5SdrX
kE4wOzRrwvAjC7/RB5YUM1INq2oNtrLdhikbgPB+w/g90g95JEESk84hoKSPfC7G
U3W0CqhgOfh9uU6vuLPtZsH8NJqD478AFqdxXMtSCryxq03F7dR+2gUpTGla3clV
2JcQO9SZb4XdhcFMfJSPVcpXjyzPHwoOA8ALdRKd/mHMryElljb2hl2uv3SAPCQq
korPp0FyFYc5vauOptPnu5jt+xgqPzECb9KWpfyh5WK7CiYhAGK02HoYilTyXgV8
t1IzYg27IGCx98eqQKILzcuNV8ZLnGpGZAn18N+uDUiLGoQUZWEmezrR3dlHDWMs
K8fgNdt1Ip9b8+PQ4ymkwvagMw/e3gvqvGr5BVnO+fJJunBW6rI9200V4Abg37lW
XFscpIcq3bgFXVLEz8YggB1lBg/4vvV2QIdUfTY6dfNp0au4UNGMIBHcH5wKxlfx
VagEwp2ZgX40aOTkuc3k6cRBLrIa17yewCrrZ3T8d9Wnfz7QpfUPAMky0N1Fkvt0
H3LIF3rP24D02wDaO6Zuw4JZ7+dYROXykfNyQja1aYgAH+k94hHda0kuUON+lNXl
POr/WXi2+MgVwctfMMLmyHzlzs38AO5LlI1KhC7NguKtCSsJhtcQuKa4KCfPLzQ2
qi4U6X4QCeeOd2IW5ll+6iZQJhuD+YieDdV+OcUJWc7NTf29xjZimm7tL1yZb5RD
2eFFuJE+B/dOFgWyiRcNVkY6+52NpgqjJH7mZTpnbVPSCa7PEkWJOzHlOoBXqnJs
jROiMGh0dD/9uxpnxMleQMAqsQJkHXEVFrRFuqox1ALOLuITItpf2TGtJDNTGyFf
VdGlAz7kC4/GC9oYVXoMcP+SKaRxzcQpIkl6AZBaSD1T6Dz6a5zzXhZddbFKUK87
YLVFPnCVPGDEe8e16EPzJVsR96Q7Zz+mXPqKrQxubZ/yW25tAtfxw7skjUyG+Yfm
l4w+v4fp1aNxqCZgswpbP7iCDy8y6agMgkU5xi6hm4YeHKU39KjuqB/+6B/otdmo
62E58aL5nLsM2tkZ0DQkIgtLrOD/EoNRGgGArBiPcaqjoCtn8RO/XIskbNlD2G2j
WhvL1bYPv1Jf0YOqqucuEUeafYgiYQUFQmY859X10ocRi5/AWJ5BEuR6pDdFseVI
+buN1SSPsm5N5Je1zkDqbKp2iQFbiic4aUPKQOmAPqMv7OMUZFTip0CKfeNQ8/1o
9MeuEnL8Wmlhhr5puiQgV7qtCIXcT4ey9/PtMsj99Wgq+183285gBOuPOkB7VqVg
SJxaa97y9XNVDp6gDxQmTM1JyKcWG5eeDJgAzxWkpxt31A7Kr2Jln+vkS1ZzlWtw
au3eQcAcsgNlVqyAxTtmNAJJRmt8zEwIdkGVslfQ5rJX3+VhYMksTDNIrFE03tno
qttYOnswxOuwMzJToqYZ0BDlfFZQ7YubrObxT1HAe4eP9MAI1Ldqkn/cYjmp90Ts
YmXTj7lj0tdKPAJmmruCztNpI/VCrs54ETNmlk3D94S7MBXypSHherAaBgl8XRhV
IOr7375LGt44Go3eFN5DOJ/KDk6x6TMXeVd0CRx4Z5Ylv1VnjxfPzH4G87tVibrW
q2XvNNi7USFqxdmnoMqEEMvhAhjmqouxt4jvcA09/26e5QdJ6HEi6TfdB0xeO526
5vPGOhcegMWu2evgy7QwU7n8h0lTyeOVEps2rd4xNyzlufgCb4gJMLrDNGh8yqHX
VDhzaaN2sCTBe21KiXG0zPBYoqXEeGdk/1b6GlhqkkZh/+p0aLk6Q+mKWj4VdMC6
SEO9ie06QHhaZDNUYAXzzOJT18mGsncslVuKZwoKNb4AVsCw88yeEt78NhJJwLWR
K5QrT39+n5yx7Qe1BpW8QPxIf7yYfTYiNWvo/8Dai4ZOuQsGnp64/NxgXezRgKVJ
UzTefhvSXBz8CB5juZPhTJxslasnTJG0KdoY5mFW+hKfWcAVLED8OsuoKJjsJTfu
76M1zeoPX7T+jRG0+MFKMR6Xt7dgSxfNkCpERYNMWmEyGA6O474LeQShQK/4NnCj
HpMbSYHI2hT9eWCzz02WD4Mb5pOEzLAbM+Bs5wV21XA1USlqNkAbGS+6t/Xu12d8
eZ5alYSLXZNmolEJ333hQZ3nwwbg+MwDKtBfDzg01P//owTe8K38zKSk3SOaq91T
+McM6WCt27G/8EMZQf9s/0MKa64p1AMi7wLkjdmmui0/M1F+OqY5dEtEwZVJ7VDW
E1HLv91YUiz+MZrLqA01X7mOwAsJvKoatrQaCJB+vU/tege79omF6+JbFgqWdKso
zn2iuoAqBvzN+Trm+srPn02M4yh0aMoGYLNkw623k0/buZHffDDrKP6MXnj1CnMD
ewIjgGb3ZQa/VWJtCLOWSIibJImLrj43/CKQxdfIbqDW26k0Ta2qzxsuTA0rVDQi
HguYfbp9OQw+844CjIJrMKEsfcIaxTUBVgJYeANC1B9gJOEfPR9EyJOhEKPD6hX9
rE4kA5JLKEbS33vQabpuFWaEIcOb91K+vLHe+EKShXDRjzZepoc2DK5pSRawrKyx
GT3NH3nQ8DaxvGPFbo24zCXWmsaYCsw8P4DepSjRKOvhjpHVei7Sy7RRKMo2zdJ9
CyNBVToqNKn+ClWlMhmGA3DOnzjH8P1fWh7aOdZdfDum4pO4mtH1okp4Glok5aVZ
kVxczPimKal0+SABFaOXnSvfzMvXYA4XOPEkS4GvN3Fnwdh9X0QuihZNIOfz+iD+
uTiu3nMq0WGrbyQpjwCeo9QUQ4deqWr9EEXMDnu2gXg3RwXKE9t6EOxtPyUyQTUl
3TO+60CmJbKUvjJokoZaeh5k/m7r2TR17/2MqieBVVfUsL2rpfWC5FxpfRQEparl
PRwloMmV9A1kubqhRsU0WVlRQKB7E5n47XScfVMXWjxbLoiWP8e/7SiyV9Ym/LGB
nLIi/2tkWqNsLyG/1GDeHWfXl4m434/NaPXUQwXdhNj2q22qak753zdl6Td5u668
TaoBVMYgPMgj52/H+E8xLMnE6EyeSv3aGgWgjoDQonVn2WPuX2HKGthSKDnZpguA
Q/c5zga0iOFFkW/lWXEDzKkkwkrHhldpIv+Cfa2jepaDTlCNBN7VoGccZabbVjSD
TlRazczbA0cG9Y3Zn8kcziXK5/vIg1m/sn7kUDWMKtI7Trqa8Pnst4LZ0yLah8Xr
nO+uYECTmD9MwuPM9U3fe9d18KGagQbxCKAFWv7SaA+fBrwaZ1mFJIQPuX/VuU+9
0kHDDsLGyCb16vrbvZn/q41/JJuop0h23col0ZpRvuYvDPzpPjOiKxxL6I6OSAml
BPf+lmq6Tj4VaTkwSex/g28i8R1XqEZrMQLpmzmEalYus0S4R/WLoTRufVGpcIjd
2wEpCZDEtFDVCmq9wXEvUNVtbHBPBa0IS7Dy0DH8p0GDqdX8DsE1yT84T4TSoPFg
YkOJF7pPZ2lxTa4dmB8+APV4UzLTWsUbdWzMwskL/rwIVKt8PfArLZgCqbKJtrap
P0793La7MqzaIUUXJHzbEGKWmrCLQj493IQ2rlMyrZ7ulOw78oMPy8IwSiI0B6Sg
SfBz/rEu7NBB9RcYW1yM7+Nz5nmGhGhiOMQ42ty44f2pmu4rw5JpBiMyFi2+kxKK
Cp5mvIl4OCbLEQrYD+AqPVWMFJDB1RZhj3v74I5Z17eMIFVnBjCPcWWW9NuHBWjp
QOaj6M8sxGauZbZChOLKTLRtvmPQba18Vjoclmlo/P2vSW8onmFPKyGxhZlHXe1A
CSOjO6ykakNMQXC/Ono63+5sQPSfS/K456f3sqlxDfwgD/aJNiEAJueIGtyUY2wk
rKZhn2CaPBSaA8joq1b8nM8v3mvXDCKTy65ZCFhiHpOVJ+YRGEoNDcEUIWUcF/mn
3t5XSGA5+XI7q1AdEwwt+7Dx8v6kAEpaFpgwLg5vdiJ+oBlDFmyVd3AIwFcqDiyc
1Vft9VjLDtrYbeYE5w1Y7zH7yL7vshDn60J3VFoC+ZNn8FW+trHQdQtF4UpQ0c2m
5HHWpMUbKNuecrade3iQUgNVlcz7sTaDuIzwdkCyc+o+S2Hd+/wdyBArEDQpmmq/
2/lNzQUXZ3bU7sIwQ7+p5aPyIpTpL7Hq7YCNKJvgu2VJDmIyzyu/6pSdeVcDWvMZ
g5QLLCX8IkpLo9AAcuHY5/Sb6qWdhPFWM3hzYa7yEHQoCEz4f+ykOvUfOHV/EbEr
00O7xhZq+TEOGfeM5D6IKtVJRaSEUPyBsCbIqbjNOAM6ZTCqOfjoxfpsvGRw+cWs
kY53lNKltlxuPjbHe/f2qMNbxtQc3nIa/TCKn+bJJXQzM3CSqvHTfaXQ3UyvNqfE
auJOL+wcFe303HLeeeb7B1thWSXEEsIJeXa9yEr9cACfFQNyl+C/G2yQPTNGjvlL
2lDKzG34EOHL8lNhKb5tTL/bTHOZ3rkU8N2aItTlbwWFZ5qtJKuxdKC3CcakJDsr
f1pbO0ljbfXQSG578BiMFMuopHfOzcd40YnQpjttgTWfxlRDJt7jHnJUpWcEgkwn
IOMimuzMSXlXD08fvoD+TRTdZuElMc7vTvuwepwEVndveJsR73DOxmWahGkC0QzR
GgGJO1PtbcpSPyfRwJKtKlOtvLzjtUUBZd6bBJdV/3kLveUGeYJeCY0VvXvfNAy8
DT615h1KX1zuTRW5sNLTMRhhN6HkQVDuaPfs7NrX32QLdHNmmybXvQiyggKXgIk1
1SMETpI21aWE5KrLxMqEh6jtesSs80ga7U79KwqzLH3ZC/3vDesxDKk+UnN/LisK
6jYMtrNr37cYo5mu3/YY3DGvglKHsyumvgXi749Pzk1p+edOuE6l2G3DQJCm6ueD
OqJ13krf1/KKXC+IdXZc4B7RDtfc4N7l2+hd6G3E9iRDb/rYKGQ0Z4viATG9ViO2
Rb5OzgU3iNen2S0NOy0H0jgK22oZJq2L0wsf6VXomZlCtqq3UlMf/edTB1o2tCf2
w/chU9eKMuy8KmMRCBPjMiYQClSmjuemX9eaPrcx5fvRRSAiE+jPozyYFUJWfRl1
Bnc3kPTLd72ejq2tQh/Mm5d0Tfkn52hrqkbH5P+JKC3Ujqv9nhuFSJYliRinrCBK
6muuAfA4oMbHcsChlERJgRnphutLg1eVNIr3LQma0rZSzrecUnkNTYXNBCEZaLiV
aLuPE+/ePRLDh9lYq27exFxzR90jOc85xKLjDvydg0P9UyaNdyDh0b9qaSCPoLFB
aus4SH8jjR+UL1moJzSb2lcyB/KVRHeP/6IrtEIJxo9tbPjKP6NKXLmX87sUqfhi
7TMd1DkxSzhdhbOuh2I7X6CQL4w5oSAECQFPF5CPDkRkCrR/ZAS1T6/PapI5CZ/V
X1Uwv5mPGqPs7ElHUP4u5PhakY7SzBCBis60v77PPMaF8UAATT9Ffp+J+wvHUfrC
JK5vcTcRJ3GzzUlRmPSjGih9DwXC8FTUK1meNRXkoa5zFJTRtcugxiPOXDhgprWh
LlOVf7G8ruT6E+VDuSWwx/GW3xMP9JwYWMhtxFdPzATO0QjJoP26mbhtyIvgC+zW
g33uzVVfu2zz+gx4UDMkLOOfMAwZeWDc1ihFX3Z51NHsreyD1GuL3eit07Gsrf3P
xhHJQKhuncYfy8dpjqrbOAea7g6HIn4i+nsCxVRfaEVsxzlKmX1emcYqDloPWbMI
YrTDU0uGl3MwUxzG+eJbxIqRCqiCFcLutKPQvNb++oKC4zjKi+xI4VcUvF5VmRIq
I+vAp1wY1FUnlfb4ebP8+kQVVRzpmWPYf0gMJMfceeVc7bXuBsm0AHCP9DbOq9yC
lYBoNNFs8w+nYxZBZO9w85C93EiBht80iWSoyrrrFvs+R6tTYMZ+hoeRoNtfIxBH
hX/cdaGmdEvvdhKbVMW3aZDoQQe7uwONZuk7vd70fyde9ECRvG93HQXjWC8/8UWM
3J/ImjY4sRB+VSP7hfcdRXh46hmuxUEaO8skQtlGU0d2Els8BjRMzPY1XG2Llwpo
8gUW21wqwJ/9eQQUDSHPdn9mzt1OM+e7lqfWAGL0/WehG0+c2zPRUzreqZO/X3PI
prM51f7z6q68rGyxsn5wio87Pz8QJ5HXpZhRjjXGdB5bTtTfivywzwYEjOBXoX46
8BK9SX97zglkOxw25ULdRGf9zstEU/4jsVMvdHp/pl7q9oidNZ8YgbhfRQsBNgKo
7/ufmYsNjIBlqFYL/0A4zzoUxKaL+zR1wiQpXhwC/wu0e8/P+DRma/odGS6wydMb
eK4GBKPlv4ZLFbB0171zvy1tP81vEmUY3MrwAUEAUD2yYZ6tptr52osWKrnmQO3h
qYEFarX1PgwGEaSXHKJ1XarSO+l2NM7XAujmmrSSAOOhwwec2ZiukL6z53zMkgUN
fVKzRqa2W0Qf5jcm2A15mqF9FLIHXe1ls+/a2aZ7mcfgY1YL50+oTXhy6J6k5FKb
hiLZy7luLwhXX0lREfP1NMLwfrbf4XqbTjR4IyX4y66ZwAhJyM1HLyR3ZTs+aNA9
CwO0Gim2aVcnxhdnCfaVmQP+MI/sfzOIYq6MR8zWximwwVhWR95X8Vo0ERLtt3FS
Bxpce11dctw8GaKjlugrZYHhiOXCxJhuTKGY4cJWoDNoyrpik2SJPw5WpL+fUAt5
oi5SGrdCowter9yhlOR/W6J3MqAUu9aKRoqWz7oonf0vFPw7BksKs9WT0bBsfpRQ
4nLhHtPbW5Z/7RzwlTUrqe+UpEy8b0zFCwv0uZgiSOGDGGC7aq+MTzEhx9Vt51SJ
bZRV3nx3tTofJGhKt5mfJzSetgcPwCxS/GBxZDKQD3M7TcbPGryu+H5n9vbSPSFr
1d0yJye4bNCO0kQeJ1mzyHensmd/jlwqEiTJ+Ajj9smH/Hh7r0z8sWHTgKhFojX0
+2+GiSwnD1vlfp5gYnZ65VwIJbe53sXw6rg1vdwbb4BYJ4gTvXj/Lad2vUdy4h2T
ge8l54ZW2K7wdMqEBbzr11p5OHZUh0ollDB2EEyvVU7BAj+bLuLNwBZWpXNFzpHU
45c+gmr9UnHicJCqe96aVkBqmyuCKpchl9HaZCBbGKeUhDxrkE602OQO3pZNtbir
qzUEtHrxSKgKymXBKerV4hJEYi3htAzslxIBwZoIbk6D2XaWHxUGClRWW5ZyFRo+
CBF+7CAvZUZcLXfBSorv8zQiLLgDNAj6g0IO/tdQS//VeWmkWna0pZUZKzByPaPE
5PczvYy96l+dLdwV6597KrP002jjtHUozM/99BO/1f/U/bedlIanmbfgOm5/k9vH
fAtcUY6UGAG/byPzSpzdubAtMNI/0PxBOIIlBVyvujDwxER/mfr4Y9COl8ncfYmm
PWYjIacKp+BgcJZ+f7k+cmkmKJwmkwkmID8xGqFQsJix0SWZ8lgQolWBSpYsI5Y+
NoWZf2pBE4ORuROmZHNN6UTYdB3B1K7PHeks1APiUhf7KUuCq1A4zXv1ZOX3hYeI
uJ+7QOy9+OnYwah5LjLRweV4rG8LRBFn8uzP/9qLsGIarUZ0dokK0k/Nwr5Rk4Oh
qjUFGLBjFe9Y/Ax5OYVDzUgvmkj+6Lv275933qSZK4QMCDc+wq+FOIx0vPdWt8iJ
e3J/MfbqXFmb+cCXY8M28qQClQeiRYzpz9SMoXC+2QP6hryigpgkOSmf3H1IeurR
9VxmF+wFrRucwn4fm1pQCkGvbr3po5Viy2pUHvJlCn9VgQvPMf2TGihTJqQpmHEb
T3bEEP0/nGwDLvrlseo1cafCDJjvS1IQKOB3RoDm0TggFAAv8HdxYs4gogBqXQk+
UNWaqEh6bN0JKHyjlXPEnKx9z//kJOkjq/oy3NXXTzCbH69lQYemBbbVj3oac3Mf
C3fkeWY+HRpvGdmREtlzCDY15a/kPfjkVO0BT+dmPbQ+G5uQw7XwUBlwnT6o/DMQ
V644+QGNyaHdM94aQq95NMmIijPjnc9eDB5AWvqjjAK127tZn+z9O0oy3cI2nmS+
0CvqvS86o8RuhOEnMQe3Jixn3YwY0ZDqH5VCP9zQxHdhDWaz71WRLK+aUw/jSp9n
FPFyIs5qHU07a+FSx4kTNyXAE5VJykHW8M84kqfCxQQbfCwLxUKxt72ZYjGRJW/w
QCGiilMlxrO7XIzBHS2zYEi48z27u2XvykiqyjFLGvUpCSx06sJJyuIQi2lZRJOl
B71u3rHk4vajQVpVZfdUc+dPTYN5tgTNCV2bkwl/WwEg3QwKQAvJQdF8wWGV31T+
7opQK2CKK3AL3ZRQpv8YcLdIlZ9dg6lTH5SOaCHTbv/HMLqwldFhSsS+JMqcW18e
gJSJa8JVBSfBFKqqtnngjd41lXUS3CNWVt6lOIhJTIAxhmSHmU5cTfjJ9SJTF02y
AFFxy7nB8cCrwx7PlOpzYYeNaF9+gIooduB4OayABXx4gjyF0x2sMR5b2fCtJ0pm
N8z308SLyXObwYWtA/1lP3zbg96T8gBZuEYk+Ww6vh7GUmmn2w1xBCpz8XZ9ZKx0
sKP6VsnaqGnOAesBQAb6Xo5Umo+bo3ZHEmxHzbqIoNKPDthQEtvBnP5sWTsVcL10
ej56IUWFX35r0gIo/myOGZ1VCzbk9p32RCb3SsS+pLLG0BzO1GXmS5W3rSGLrg2e
nx/9huOeY7/Qy43GLb8gFdDdfx1njBuEzeUk4vpzWGVW0t8FuyTSw4qfRwAVqZ8B
gv+gWHDMnVgMGywN/tkMhiKzrwNDEpYY4ZPM/bqkWin62rC0vRx/Ej0UcoiRHwVT
tR4hAaJ0/UwttiKQm3/8DYA7RZgSE29NH548Wu6u9dA+L/wcrviR16XkEV2jOK/v
DzbqqF5NxO2rJ1hLVaIbgw/rjRtpBAW7ymmzfRo8B1bDrDfptTgnjD7mHaYNDX0q
30AqfMMIIWtP7QHdb3O/AZJchxebv81ZBVDsFpDmsIlCLc4cfR+YyREKEKmPTiHn
Z3HKZOqw5vCL3DZGiYUua4isom02XLucFo3pbXTaGNfmiJaKOzUZT2p6cTjP1YbT
zlaa7WTJSrbSKnQGDp3eVwu5UDLYc8mgF9LGnUT+9Q0iMDGOkA1PCqVXzTm9HTNk
buWx2Qt5qmYyPskZTnE7zgRjC98vFAVjW99NHDUGNWpVAdQPnUlhC10Cx0UPDJHA
PgdEqGBK2yoIrx7bR3mgQLhpS0GS+gGvsbIfwhqWuZy1M2oibbMOFrKsRsCTYE6o
IAdXD30cLyGP1cwFzBCx0j1FTp88CQFcPzS30Xo0vpzdUJtmb9NvKPInrIpsixNg
MVXLbYryGb+K+9IkI8WgITwA/7FWon0Fj8mQKX/+d2fcbPRWRZQrnQN7kXN4nSCA
CL1vhapUtBNYl3QYN5C8HMx68P8j1gB5L0/trbtXuWlpnruNm1cIQltGzKeC2bUm
GO80KrHLsbUG58Uhmc8dv3mRihM0txf7iIa0oFSV6gM/RlAXRtuEWTT1DseQDf5W
YO4TnsDZzwbRo5zw/vc0bHyBv8oQ4o0r6sUaNO9lLQUsttrpAXbSPGvQSTRllB9e
k6de4w9d9V5PyL+A4QE52kUUotPtUGZNdG1Vl3ygqFoB7nbpzx7II2xxxQ0Ixvta
aUsG5laChdlM9KGEzDOhHAIWH8PVh3HhfiOrhkcNJq1PRdk78mitugxUP9z5VYFS
FSmbkxiwackNq3TgxkMOKcgpnjq4Qen7ZliMr9in/wU26zrMyntn+ogYzU3oTAVW
YF3ww0qj0wXNwQxscIOGxdVfv9ENxO+5qHLCZ2lZHI/Px8/0eSZPGOQso2Ex9uvG
Tq1E0KFQbnkVPdiseI1L6PeczvRxoJ+ceIRjOwsFXXQh0jW/ocOXpfKJNbjVumgH
NmNvfE2/UBEwAkKNzf+dMljDD1oFhJN9maFSUYquM3ycxURcZYjxVaN7gQUNcFh6
k+uQwRnAeL7aAjoHxXogDWRXVrEuYDpebdCzRS/CqDeijPakN9CYTDpWTvWEe8Zk
7GM4neSnWrT2ikgfGMQbt2cG4cD4MPsbxOV0lPOqzy3tAgxVPDcFSC1RrnIx3qLB
rWwjbvDURxH1b2N7UJ2m7qV9LVJCoYautG0wuuLo3TMmG88xLas0YhPrBmd6EY3u
ns0nIIuswz6vQ50mPWKzYv7UcZ4qreI+/Bl8xJK82omVF9pf2neBqNZvGDKt7Rzt
lzO0rv/0XDhK6dRrV/p9ftVt3BN1Rr1XOqoPJlAJ87XRbh0TNRfc+ufJWqL6Tati
bI+4BBBdDbFRAcp23Y5PCupHJMHEfEalqUtbOPUBmaBLA7QC4uoqL4Vberw4xZ5b
vBKHfWDH87PTUbuvqp/JoAXf2qV4mCG0eKJnwKwiOWWSmMt3A5mJcUsCmgOPPCu2
KExaxxK3jE8dmmBvCH18w2z4ONfwyzbKFbqPdSwRrYXpM8U1ofwLMh0/ut9XOO+8
U8fG7v8eRxWGS4nLbE4DM1tjUBPt8OwasCfE8qXevMP2Yw4Um7M69vVYaTbIINua
HvHOo54zKIMqqVTOBl9Kyb0TUzw+mpnfj7ASMWTloc7iy6+OYkUzEcDRYbpUkl1c
+oM9Pj4sT0d93/UA5jYmHTlW4yAAz9e35Yio052T583aNUXTGnDqw1Ba3kVMseZr
0qW4SeuI1RCX7I/YMSuMTx34fkLtOcoqQTCjw0V46Z5mHy/KY3Cn04UR+SebQexl
c1shVMoBp29GA9H9K4ESvnXHThiYTnwE2Y/dgnqSR2idbPKQSCKTllZzzIoq/YJR
lQUSxZSIiJqNnlNygyTosJs6E8UywOQ72vJ6UQPYHm719WQK/X/XEBJtN7YIWX0K
VhdhmdPm/VK6oUAqovz1qWPhnoHGdjxrtHBS6RgQeiYpsWIyNhoc8gq75gAY+aRL
+ScpI+/YRIw1LFx2hgguYyeMMhifLrxS8thC0w1qEcjDS/jIvvO3a+p8wnPBQLlP
LoSQuHUo/bHJYJsa3XQOtsNLGS8Szv1TceLy3hM7vlI8YA9DyJ+uEIgW9LQf/aa3
UrrSXQehzLDtwtIUMb3wGfmAFzaPTdYdXt3v7qE+Dkkny9Ib42294r9lpv7gDRV4
VvdbvYSaGiOu60OGLMIJ2+7bcnqnCCd1+5BWJq0TxGYI/datoMIAvM7M0JNT8Dr9
8APXThvIB5JxjWS2X4X3YmIGppxDTzM74QIOmf+KOP8L1D9jIsbm85QKM64YKtM0
HgAUy8+QcK9RdmEXFhHfXds50gb60WGhtdPe2fxRd0R0jfstcupsfNuCfD9gBSIe
FfSzG692JXVfLPphGEvj/caTgW6NrwaGJyodFlkIGzQtgFj195L0fjFFbsCgpym2
vzSCaqpPV85eSDE4k+wsJtJMNaJ8+0Cw//fRXP7yl6Ftt/AwxlLl/dI+mniTfrmJ
uPidZoLW0UM2I/73qETDuWsS9nQhidrfyo1zDthPzgNGYm8R9DXlwJgS8Q95PZsH
u3j0JGF0jcHHvUsoNKtsBQ+W+dMEE0iTivJM1yNipIAcHWXaZYevymyU9bvQ+x+b
/aWGO0vR8TqKF07ZIySBg7YV3C+G1l7UM/AWmhXeFQp5H9r/yBz5X1QFK1xNrZSS
2G/QPMYUVhHIMePEt+IKPBrbWp/tzCYOW3BfA505VkssgGVaFgOlZO8zwskSRMc7
Mq4DnkxQRrFnrFzE2Oc6REHm/Im/2FZ+H/tQeCTtp3Zd66ZEeabDHX7gC+6lXkgc
HNSHBMioKwygRJL4RKUShhaWUSOzSPx29SlysLJyqt7YLc8y0lvMM23CHQ71O419
r6HZYf5t2BHDqOV4ZLJIviypcDc9z58nvhaUVxuRs3J49yO2QR04ULqQEEgmFFfw
mxURETf35Y16V8yVRFSdEFH802KFTkFEnH2BPoLGkUmJ4UnVDJhbtHam6aukkHGB
s3UXQxMJRqWPHC9lxkghkwH88DTnU3iPhr1Ik9ucB643/hm28Vcco6CpDHgb+h6c
UIw1CZLIfHfqPH6+hsAh0QZbvc9tYar6TsdvQrnAqu2cQsRD0wjN3L4Ylzedng17
Ulm7Q7W+ujp/m7nGVsFzIJZf8BbhXbc8wirK1vOk6FKzqUBm8cyVeNDtnCevBIc2
mOIFHY1pKMX0a23q3Yfu6S5kV2AyhIeBvCk2PbDtfcUVbPiwNzjLwCb1mK46z9M6
q8HybNeOljKvRbOJDVcpVZBwWiK9WhdczYYSnJCt6yVS5mj6GoW2qB6z0Fv89A4J
3YZ29YK9NGbKEgNsk9pEE8c2DlkUQZBiPbaLGvPzGExMuqQjwI/D3EyB0FSnwEPe
rz+Swke5KBTWKYouyTbsRloZyXlzz7GZ2l8BmlnghBf0DVQLeW1+jRnieKu5TUNg
Tx57ZQ0nhw6+MJTTIR4QNml6unKjlXF63EvP9IxmPj2sjVxY0lRHa0NOBYMVVNjY
3JGOCD2Be1EATh9PzJL3FIKPwMxuPEMCVKd/QyxNqUzvRG7wTW8JdER6iP4XrXBJ
vQMspNH9+qvZuCuXGmcjofW+RrK36OKvX0GQhBf05DQr4VCws+hkurWzSuH461wF
eygk6Smp7mw9w+dkLsiELQPmqnv1J6f+HpI5c3ujSw9UV50cWhoDMcvIPy89iTqj
B5L3hdXEb3OWJm1VfHmIkeQNz04cdKYAc4FpptluUIWA2ZlbN9w+wRMshVr9fFwB
BLkDSpNtLX9WtslWdFAAyApm2AbDTz+RVdCSc5/EN3NyRqWw6RaUVML9/FkL3QQN
xaVA+kYqD2T+8DkVYBI6Sn2jAUsaQRCpjvxYOS6gV9d9c1LRmdX0mVahWZRwGitZ
GMgVsTTrBq5Ca9QU8b18AkyEr4m30td1XoATTY3U268FFptq+TuInaIToUjSkhkD
Vfmwvn555sy0J0VVcNmr22urodMNEQ7tTo0l7qAhf3bgiVqmgwlk54kxLnEVwSyb
+9l8gGU8w8YQPodL82xXZmuZ/EnpIMU1lXvM/L3/KAoP5gIuwBkS5nhsmijc7sZX
XQzAFgd6U4TBXQd1MRzvSSebHl6Ys7Pb36S9HNNhhWBTGsh0yWmvusTEIg69GXpI
EZ/rJ57yYPtFpsh27WKA5yb9akLn3J3w3jd5bDug5Hlkxb0rZPuJWgt6MoVMKR9D
lAOvhtBWa5u75/E8CmYuCJcwbNHrVfLKwriA8jprwDyzP8hAAyOc8nynDi/9zJ4k
MKfIKgN5UJqOY22v7teVllf74wtThgxlq5R9rpo61r2rF7S63dTuaFwGru6fUDqJ
N4U2Muaw6fFzM0jigOE/2XhJib+s7t3x1T4rIhAVLP3Xu9S1QLsfWON721HLLvHB
A4SqdXovvBCBLDMmRfipuaUhrpHk7qei5e3Q7bUgqg7eLEAcYFik5IfdpbgrVVIk
0gPuRARgDCJLBsmeR9xe5NrkgbufCxxc++VhkNyyBep3k5TdrvGKtwFlydg9Cazn
IYwCfL6AKpLkFjs/V4UyKAxI+PdDWfEQXfoG9d1YWX9qrZCSHQwGuZVO1O1zlSr7
1V5PwQ/Pm5fNxh2Sbqf7j1V42BjQqHpRJ9mW7stEGNaN664dzDSsdFtXtrOEMlNw
zae2X5iggTGH1iDMK+BlpFGIoQFa7dAYWcNJYGYJL18UMkGo9XUuEoxHARMRpct/
9V+zN3OjJ0ulg0ML7qJgFFGDXXuDlSeJvt5b2mAiZZriNrqe9T2YnM2fWCmHlqcG
ZQWkCfISSiljTGw2YBK6U2TPiUHZmLIBEFdj0YQCRdhvkijf3txNItd91PidGlL0
zqnYHpDkts/xWsxzWo+gf1vP9fwttzYqpMXx0ZgksckeWEp3MkMZi6jeNA0BBIE2
70Gqh9N4NH3LReqU/XSN66Zwkf9WdP1P6fOkYS39vxZfOL404x7VN7l8oAHL8PdS
NUE9WmSzEqr8zW8idAG/qpkp0j6Y/gsw8nV8HcjdxxTIlu1t77i+MiPp/BxuCVkk
VsvWMrpStQ/yRWpajkdx6l8Auixt3667hNQh2TFeN/cVIvxHA3JHHRnLgkGn91gS
UVNT5e+wBpgSxbN9gcpSdbDSJUgXC7bnEPFhTwYo0nbrrTCE6+t+LAebnnflvBt/
szXD/2wT0Gnai/t04Mly0RNyaqNXDjyo2sbkX5fdt2svqKYSOdCPrSezWXs/k+KC
1hJ80UgURuXcK7VvWfmeRieBGQCjcZOVEzZ8NinhBRz/eRdaJ3Vy4cLIllFT4noH
MFROx3or0uFR8cwe664RmgqaEQLEgYsc3ciBhqkyZeO7cMfCLVZTG/bSYUrWmH9i
gi03PAkpeGL77ZKzusZB4TeYKI51qdf/+qum2sOwYm4D4guKtrdBZZqWOG7ZYXbv
68F0zypdCbvX5ReUsj7gzAMQkFY1S7H3ydlrQ7w1Q9l89PE0uZJqGlpyK0EO7Np+
Hi1o5JsSE7rqmae/zdVqgBnd9xrgCIQwZ7FIsAwpDUqf3M+ID06L82/vcNr5Y2EC
6Tde3+pJcjf7XN4Q2h+GNs1KlD8h/pK5zAZBeL9Om7fLWM9YNogy6VFcvPyTa9Im
yWIdlz3engbbFF1nhMMINbEpctd9xIID5iw94FtpY51qSKFin4X0DkvZwybJSp51
i4MYYd0q6WC0acogq4+dzAEZxl4fnSiFY1Wb8gmWrwjXNpiA8OAlyEjDIvD2Clio
W+QnxuCCEGkl7okoLTGRHCfIFWqjeCeOANpN4WG0n1hvFLP7kj050qBDpur+In5C
yOCzqpsfC32uTL5J9wI01QCdxfsd3yDhRspQqoYS3ouXYIH5iDwDX1cyW2Mg+ohd
XJLoAVL3yRl3boPT5kIlhJuH8PlUXtZjilSbhiGGcZ8UiThVqAGa2d8mCqeSh6Rq
wpIZdDG1dywBYn8sPRen/T394yiUzaDUVg61mdvyayElbKmu4dgGJ3z+5ETBfj6I
HlhlIP3R9Nd6r8D/AGR9IahBRe93mo92PyYabFxPI0o0Z87f/RDZqPNkuaP+S9/o
0Trbf5FPPvuAasfXhO8G4gfWSPXuXFwopL1kpJI8Tcv/2kO9jgzrrkSAPAs5MWsL
dF/WBvruwycU5z/VDp3hM1qAwUIbWydfGWU68hyOhJGzB1nkBt+JHgimfHYNO9ht
Vb3KHHFmrJPFGKhpqvbyn5BiF91j1duMIa8Cfv6+5w3PAZouytiOcIIasMmedfjF
UYyoY81VoNdg+ET2TfMcLzKPnCjLSxT9FBKtoDKCrMofHBKwlQpYHbVIxh3RI16l
jsDpEQpMFgV2pLvxQqVK38zZmnn3vrze9LuJu8j7S30CIToFf1ao0EJpKe4a9iUO
PjcH1PJMxa5IUi7m2ckjk3jEtz07DIi5Epf+jLXrfusL+GpStFmEsc0Edtd+GJew
iT6hqnSu4VkvpfFfbmWjp8q7EANyvCAVt7KUE9Af48VPCCmXgF569RI6qpW87dlR
/9dMQoODWNkPB60E6BNXl1JV+lS0HT5NFiAmdde4woL90e7kjK6D2bMduJFqeyDj
i5GHI/qO/cBvXPyhu5fZac7inKdZVul5sEdL3wLfBrlmobzy9TBkui7jJc8GjfIU
2cYaOpvRMe5T9qPIJE/B6dEvZMhgtAO4a4ZBF2DsEGhYsYBOkVLReVxCN7kPM7lh
AIYrgkzIal1EkrGvlsQOEaUJNwOsUX53HWcQOLvoJWPR7K754SDrxsOxgqzOKVfL
lsSpzzzw1KVhJZjWSrB0+i2j9lAUipiFEqjC+0ZI1eXHBXAS8SeX0Nxfjd3ycPTO
JVQPT0En2YPT4qkQFeAJscGlfau92g3MmRtPeFHpZhHNVxlaUssdFsyzI74CIeW+
Wu0McZ9PGBgOKGte2Q/ivhu18QocK2N8Dt5JYIFcUB3rupO2J8Gnzxy/bt/+SS9k
gT7cfSXV4azhHrZlLsUiqiTFm5lE1sdg5vHWX/ny/Hk3eT0HHYYQFEJIyk2uoRSL
ysiUuM3IvgEWNvYwesQldZQqXnM/Hx4vZq8E/Af/nAm2iGnz4Q0hLFJ6IpUVwmy9
aM4Q9wZly4gPa3ObyRuzgpXxuIGUEEaz8s6Oqvcb9OQoYpox/u/3GnUq9FbuDNJd
iLTZx+tCS/5pgCjz0q6fYmHX43O7LvMYcTCCUkvxWeezapzOcMmKuTur5CB/7HD7
8zSf9zhDWkOCnFHbw0pItZdqqsNM9oZp0NCx7g3UjIZ3CQSuXR9TN0GDpEreU1Wt
6yhYU+ozzag9eMWvYugJOedCuimlrlSW0Ri6LCFuTUboWSdfsj7ERIEIpUzSZfm1
1PcMYLSQBNkwMnpf7mTPiyCGYXzDHtZAHcdrU+l85yAwMJk7tgxrLTYsLP62d95Y
s7a4Com8E6d/OTvqRJhIGD5KITxw1zhTcP/bl1JfOzCwo5GzyjQTZvptBPuj/YE0
Az8vnbushbVJk1tFR4LSISL+HD0QBIsKKFAGJ0smmbRlhVdtW+4y58HSNOVg4x2V
jqHGs3OUNOzHlXF0dLgPRuKHpdUCBX2sLXZpW4tRUB8fZNqH/aRHaKPnhhkuy6+N
eps39aNhTrhk/Ht+lpcGW2ODEwcvALXWvJLQlpFdAtwYWp9VjNfl/iUHwO/HUItg
ISzuYjtRSFU4EaAHbyVk3luLDIa5YIbvbkY1iaZdSHx94CeCQs1dcJGWEk7nYTYO
GrXgT+f8y0kMNp/3BJBU8OmhLY4zGvTGIqGEeEJTUE96clYoocKUs5YFF4g6Uudo
Er9qcQAu17OT/wspsi2Dy8Gx5SODZI1KqBN+jwaa1s7J7+enNgq4b8lG7ygMOKCQ
szbhLDLinDPvZNQys9MVehFo/83AFywVL/zdZSq72v4RkBAMB2b4/invBQRV68DB
4P2e+KvvFV/2gxqWBIuiVL8zUfNzWC+5JjXk/GkcMW/AE/iAEQoDvrhxj5InK6HQ
ZSpevMgrzNzJU0snhObMRE0bUgbSBiLDO9aRR63wEB+09kDLuxsDZGaZ70eYAfl/
fN8ksBGy5w2ljBVBRKLU7rNcJYFKLUADpsgv7llr2BwQeyedRnHrn2pVpRerDSxr
xmnmBKGr2lZ7I3G34DJZ4+jsutnWoX9kmNtnXuV2NafIVh/qCBXYEacWZVnQx9+u
bALEGdqBVlKXbqn1VAiI/MzM1qQjthFZgxzx+s6C5IGSsZzFSTzkK85LgnXHM0t9
i8GpP4Pk00F1EOjS+efPJkXfn9uTbAWuJe5K3dvohLssx+OJF32um6dtk+CFGmTl
XB+xce6VWhYx54zpupLCp4Wrw7ucXVUVqhmavO3l31WMiQ4dNXIIK33hoEi8UepV
I1TNIX7h/hcjQvCVHSKZc/9jNIfmn5DDbEZIZl4WCPNr/Y09CyBOVPvfZR0+2C8t
63aXb8F52LZS28uwIjaJ1pCV1md+t549LanPdpncz1NzeAmLDgUO4M4dZOeixijM
d1FRxjb6BXtj0i1OWeSri+25nmNSLFRr0zTal3tZEgtHku2OPda4WnACnqDSIWDQ
QaDObVtfoFqIRF4BEYygewWhMCJ9ckyB1OaRv+qsEYjsMOZr4Ar0mkkcmXLRiu7c
ricfVmsiO+nuFUfIvvZmuI4h70MXO5fCkJ+uW/WEqAvE7oYF5ZWb4rpoRg+MaTK1
LdAXH5Y3hHLxFsjbaYt9c5AZzq7obblLO+CxNnhzWE9yRTJ0a77vI0hcWd70oTRC
6u/8ef48bY9RrOPDHrGuVZ4YlbNrOR/GduXn26gjxfOf/uTUJyEZPEFLjxfAwAwe
CS0Lahc3WdGhc57DOv830zVx2ZOoZd6o/Gdlyyp8q0H0+GPGOKpc8gSwbOSTQMEi
/OJ3y18vIsI4QqYl98ylLYb0MYTpVEhY0IC5/v4xyvKGAo8XmxSorSJjp0NgN915
lldGgsmepl9UpIzEBkaA3fNY+p3A+X30WLkn7/aP698t0L+NHqvQsPbOMA8/Xyry
vhHmhEjRPKY+MDztV8dvNuNDA14pqH8QSU2VRXcRP2FdtT4RhAsONcWbsaDs+ncS
VHdPZdu/VF1Cd8u4uaWAtmUc+kthnry/xwNNiJ4uIOICulPw/4BUEeVPDx79Dk85
hZXDitjPorOC6V7Ke6qN9BUHueOHbhc61n3yXxgDsoLNx5VMQmEssQdFamhWISjU
iFJ5lqzOESkLXF7IXN1/0JI167VTvRLAvdZoBSZhgRoEMDGj2Kb2lYDKFhmYIhQk
yjdaYyi5Ly40sv3EH8F6W3CPNmNyILzf+RXVUnpFrIt2sXWOKFszaYk2q6B1LFam
aOtxcFDjEJxxSvgS0N1MB8Fb7B+0yDgrs1BqAVbg+5Yehlw00hqGdWG8eIvxmqFr
1Jvx9jzKF09P653cHncUarpkgJCXrYhDrCCvMIIMpIo7t61OiHIF0dgSt4qRqPEM
0y3lFqVzMoLeLaubbYPSpAa96DWTFpuA+9iYGQKw6ZSmlThyNd8yH5DK9dmEk4Kt
w+Lx8IC+kN+VqnIZv4K9BUlUwfQYGsfrI0Rud/kTiyc3rlZ2U+o4dKAhgAk3AoIz
NBqqt333w3zOLStjEDLxAbofPWdPX7erO0uAA/x3k6uyMRBHOigULg7KNe+WWtBJ
eIxwe15emEkKLOOBL7beajlV8ld5w1c2T5GABvmzNvVm3WfDLB70hxnmqkTuTXxd
3Tji1/47G6/47yynHnYv1TLPtzy+2PkiuEBsbuzCUVMom15zKtSiyzy54DnNerjt
PPpWwxYXK0r1TIlVhTFeC+yCbIXI0SQ3v5EXknOTaThqC8/LgaOdQ2mfVQqgS/Bk
zjM1JiPwiPtfWzJmfJVDpRXodFnQCWj+pO/BtPJL9YKI2aWKoEp1n4QweSiHFORT
tWtS671ashuaFBW3btpc0ZEfMy3UFoupK41hS26DseXX/PD6v3xdRuIA/qP13WPO
6L4gWdtFwjIjYlKDG0tAEGqg8x44CdiazVpCAYpNa9TGQ04HOIAMiZpseTaFNDvn
UoCTuqcAA+e0n0LVy3LHByEvRS2pCd+4Jm13z8UQ5od6uMIH87zod2vIRQMggUeR
wSXsBPiN8hgOuZJ4wUklxyJkGO4R4CtEj2Cl4xved3izBXt4VRziEyWtY76RRBGe
+LmjTUdzknBzQwwhz97C9+ivKh8BQ9ZmYsvkdG0vyNA7kJ+FerZ1h5oA/QCdkwfF
6iXTnj5nfxNz/UQE0QTLJndQ47jI4i9e7nBZzErihWrUdTfSv4Kfo2FIJDkKi7ya
7hUF7C0/N5i1hJ06jgUlUHWSn1RER9a7NHOms7sctz3Z/tc2aQHsTBPuu1X6V4Aw
l2U780GhJJ21xLJeVJ5ODw+UUhQ6nJtA44FZ5MOzaaHMCVimQ0LYvUVaSyrlTQFt
Bh6Ai4h/gy1iTDBaInIDW027t3LipfE5YDzQrAT0Qp+G5VorbkaPDsKbDtSOse4J
xi1mnA7ZnHGvUDRtqlJPQjLlRobHdIGgIxwXHBdeg2juFVxb3mcEwfklVR3w62Vl
0sGv22dsCg16O6wNzXjDiLDBwozUs1Ar346CJg4Ih1glCJ2TCKEfH9pyjxLdAqA1
FAC4VJI2OSMLI2aWIJbE8JifuZkoS+r9TvDXWBqX511A3hAev8iBt3W/SrqHgIzq
mTanLlE72hRsL6WQieyhsJW4Y4mk8UO4pVhc5PmNGhUvoHcUf3MV5G87l9EYXBkA
9z1K7M7jj8zwXie9yEPhSbo+8oLsdAwnqfE9EaQU9FNJiYbMWAUgJ/Vg8SgStQ3V
Xe5KDEPIzeZ2SCXhzAzKOwmGzuI4aZS5nyuiLeS0GHwNLWayyCkydeqDuBkDHJIt
Iaya5bPinuftgM0XVWn5uGea5t26x+UJBe0qDpvcZICyTETfv7nr8pdB+wOh9ITF
VByyJUJ/IsSVXG8KikdfizWkVw/H6YqFonjHNhOdEnTWion8M96+1ajdHWrehRCo
xeO5rYbiOdvFPTYeXkaPIWwTJ7rNtHTWxfjN7b+M3mizPnsrLaNKCW3or57M/R/1
vzgFnmnm2FDkqRcze3r6MRH3a7fi41bofhw954lZiu+nL4OTt35uh+zaZShTkEjT
Wdvm+FqdXZlQyZWZgQLfYUgpF1kl3iosWieGwAPubgrRbYvaIpWMqCpYF7+gTOJ/
1WCrbXi7eLEZ2VQQgsbu5ij/z4t/mnP/wSUwrKBgV2T1HxA3sO+LPKIOCGPCqVaY
80nTde2OREWdEZND1CxXHllJ85VWVYQ48lMKug0maqQe5E/xjNirIFVaqSJWoaMI
I3udSZNyE18/N9BLhPOtg+ykmfhUjC1bcrnhjlC1pdGN+9t4TIU3SQFqgADAbOsC
EX+bkUgAfJ0j0+5JHnmed3FKWRQwtRonbVBTBDVFJvlbMbsr9gIlB1K/X59ZJFqS
/4bRmYKxItgDcA2KlPNx4R7qdz6nNqjRb5QJ2iYR7d0lremkO0TGmUS4RFQT5Ls2
Qm8s+uGh6LVk2VRRtsT5nf1gv0Fk4tUYYIMuNhgdtoYydlzlE6sNoeQrKqGlt8iv
NUmoQavHhm+d6+AGO7NbMAfnkIkme3mBEEdIM6k7VgLL8YuKBh4wvtRKvUKZIDLr
lKuBs+Jzo88ZNeviOdEsYt7o6LkSjrtR6Jc9uBU7hZqNqtGLsq2xFdimkoKcBrfA
IkpQqZp4ngjxhR1WOsTtUgsO3hDJbOrmtIZS30jq/YCRYLYLWL5vQbMbdYUhEtoc
PwOpK8EAuCWJ0rNE95p+GjvHdJfTDaZ9dEMcn7uR8qoS/15Ui0KHjk1P2M7ag7th
iSuRCBV80eAG1nZrLFteSMLbv8VWSFGHV/LBlJdEpoQJWIpqJ5WwOodCU6tdKyR7
tQr5oEzgL8by6RzFdJsrBhzBcGTKce3Fr4c9JxLa0AlcMUz35QafDKg49P8u4fBg
ZfQV+05ThAfijoFZuIGTn/PXHinbo/OUZCROs8xGz7gl3Wk68/qq9wRfpsq23Ue+
xtRLAERMfVnS3vDwpdxmkRS4bhWCQtXSAJn0/EKhXMtHjrXeZRZFDfjYl7XnttlT
Z4XJEEIBIT9QskKn56DmbG7tWC/hkcGTAfhh4lENkx5ygFUK1/JWdhmJke7NM8OC
gHMpgAFSkAqIQVh0DUqA1Y0Ny1yUKGU7f1KbxEHclFbrqWk5dQn5koC482JJNTOk
Yz14iKczxF6LFFJp4VQAoe59qZPyxFfSIv+NPO2/7QJ3bqve7K+TlH5uhiDLiUxT
7ZUYilx93tVTlF63WiRc6+AqGre0iTI1En7QGKIEjt09WKS/1BAJ5d7smR7/HKvo
MRskKz7BZ0CNxPWvaZGKOblwl7UOlRFyGrTf0YdsLk2x6sqwLGD5RHmajNiDgaRp
8ehpeP1g3xZAODjId4x/WC1GkhVb6NpiSmsXoxoAHhgFcss5uNJjDhpAjgFHrEhk
vo4NvT6GZkS2LHhHNkfauhXfBIjkeniK9unn5F/KxVqmLger3jQHCuZjl7zZZHHO
c5+fBZ2Y30nhQXIRJIsWVx2SmvAM1W2LPuH2x1FCDINUyxroCLyoIdfn6hOc3RgT
3h6e2IxFGyXMLRHC9sSRo9nYxOAR746xARElmA5C4KAtEu4+MGMt0POaFnNWJpJ8
Wkp5qox2VaPW2Msg9CwoLW7gmYkvlHGYaNWGnNMt5YAv1QZv+PJMN1X/s69t2ITL
kogO0+3Lxk474k6XELa0s2ZJh2/b22tHjLhZifuLxVQNue0YoSA12n/yss7wJUWj
9ufbkIHV1vRDVv5Iw8R402NcmcG3dU9dXUUuTgjFVJ6d3MYRKk+CKQ6bOZbBilCX
FYc8HpdTutA/ufrtjEZmz4Tb7gWx3FYzKvpQEOBuC7ZIDOaRBijoCMz0Jt8GC76v
VQDnl+s/Es5FHDbgVNLhniRrwM4JNUllBsDZHl7N22IasiXIODXYAHUzhFct+75B
9LiQraIGO4hdgoveKdWm6yzeSK/FQFI94MOjOfvQZkddIOypkeDDedEwszDprjAv
miCSyxmd8JNPQPjC/wEvKK4ZE+jQa/PhT1jKJ3VDs0uwD5WwFC1yM9Tiwa57VbPo
//u5VEPH3DUWyOXYExsJEzmBLbwgF9sPjQVOkC0HeCrBXdyJikzMM8Zrfwg56lYD
IqsuAPXd+EYItlo2WMOxdouEZrVjulINLIrISoozDzpaGezQ/xXXuhRliQ5zzKNl
pC92KVN2CBWBA+wOFNQgUhPeiw+JAe5p9NCNTwsgipzrgt3W5Yzkl3aQ1kKGKc+Q
B79Th7t0GHgCW89BUkcEYGNp/EIGSZWhOCyKeEs3rWF/nD/MqjEvTQaCJ42SzgAT
p0zIThZYMGHhDUjag2WLtUa9pQX45LLzY3/1Oy3/1xyZyaAVAABC2uASGUyjk4q1
s0QY0ae8ubWRPilUVgrL8Ks9qxofIWAuxCgAGVk0sQh5/eEA4HsvaH3I8e4LnT5i
uoWNEk+/Vtp3UUN3G78sguZwQqdlCchdHrP5CUDXmUL+8lt1o9sZrN+0u8aevHxz
1jKjraOi7zPxZHHjCX7MijRGm8cb6v1BGzyfv+q9Dxzn9TqUyRsTJGjqaooGZRO1
6RxJqARn+BIP1p5pEP7MNaXNh4fcAcLNONXUMvJDrAcNl4m8XfvdqcNBOZqhVRcs
8nJYE4OCmIhPAbSyysKvf/iG5Af/zwxokKtSkaijGGPDDRsdDHC1PPTcegBAP929
6sUsQpWWVcvWLojJp6JCsnN2ABgrPOIGQmGCgFurWHGxCUtuJBMxEbpBagqcLnL8
P6S7jNIksstKOz6O7vRNjAdnq06kC025QeZ6SAaQcN0m0R9yVaxHIWHMlnKCyPeN
3zTgCDGialkTz8C4mJgS9V2cTJv6vd86kDqiC4XUk59009U1XQFmQydr8YA2V01w
cNffwGGUnWZRXAFvBu11/nriiWTo0nQzwOIHQbh7eiMf70VHjdERs1eosAa4/e0z
vQAosZ8uAJMS7vV+qZKkqWzGtmzWGwGD+8rtUa6UiQb6Np/snPEi7x/kINpZEW5r
HZSm2DeRt4dLAb7zNks3NGf+93SszEJ25HbiOhYtZOFWNSZOCX8/kzIbhtRxDhxr
N8Z2TqDbF+JjaWsKm7zK/0iOhC3YFtqgcHVMT3+V5n2mVdn521pzt7g/hhuTRqle
6G7m3kur4UlVs4M+oesH5TKWG6LDLaGInssBaQDq91lXPvhx0WdktU8OiFGQq6/x
UWkdjhQSHmkBDPmzw+4VedNAU6ODpbzeHIyjZPPSTF/1DSSfsH84WX1C9LhK9UO0
GhQD0jYdGK1kRt8fIGMgUq+R8CFfDOC1dOa5laeJd8uZmYRBffHjekKg0dbWqSlm
xq2xJnKZWPz/qBiidMqC6VOs09zbXGtVt7jQp9dizRU3lkZyTPrmJAupttpKDOUl
c1a4WAOC45NV7e7Nr7okr7KZt8exiDmVfypioWqDdmY0UhkrY1uy1l67O0B/ekqF
1LFlTU6R4DX7d7buH3uQkFalvWL4sIlaYJnt4wfyBdp/A7tPg61BjzUt4+i01wcP
B8qN1mJ6G159Kzt/9pZ/su6ZnOFAq7t1uGBhnkw0x7tWUeniuoEmMD/GTGmT2ba/
r1GEqEPLi1kpkbtw/ABqIAeBwUgZ6NNeGDwf0RoRTY8G3BYEJaRTRxSmNBGy46cP
cYzDYyDoEdFEaycB/Wpc9nLx4m4wNd3SFuZVwJjaxNapFbqUCdoi7mrLEVkeF0mL
+VQ5KuUE1JtbvBIU9tS22KbUVqc2TYJpA+4/MGQMQ3MexQLLW+8veK732k9d6L99
NrbhN2QjbCWyBVmDiUGIRjoeFhDaJIBLXD5yQc9b6Z9RmspamQImZeVIq7ZIYqnv
kr7yvtVX4xK4T63avbQdWFhGGlZGz2xfonKailW49KRW1mq5ccfIzTwsj9jF7zAk
f2wcrYDl7OZSUAFVsqf/qM0eBVeMAeQ/YEC1m7o8sBnhzL19ZHHAxc2/z0Zm249H
yHSOMn+Fstsvaq6kWhEZi2/B3pyNKjl+9p37Tn9eTa3N49H9pvvgXUvI8hdp31B1
JTM7dylzMzjk+JdH3xm5vM87GZ9c2C9bUkEqWqDxNCpg1l7b3vKcp5nicFzEvyEa
ge4yIH9kjb/6WcBZvsmWCrq/SyoWBSIqVcUwLkF7AWq3EbplRSmRKo8TvfzvX/Jq
sh3cVuncJVAoyllCVjtkCMG3F5GZfQ0RMDIoBLu0Uj/buGzjv9NhMgHiQT7+dRMt
266fgcgc8yr5CxfKwaZ/vyz9Cx6SfpQDo+5RPLuY23ylYx6kIG9HxRrjHZ72yBxL
eEaeEZFBZ2oTmF2qi557MR0qZBoYqhimjrXF5GS6A1Q91QKe38MkGYaQa3CW9hCy
qUjKWhmQ/OjThF2Gk9agYC63zNnf90y/oFtm1RHh54zH9t7rxgUQnvjo4e3v8a+V
OJM0JXqRr+vlr4jFmvQE2I+xizztofWDnckK+w5gllmqNo2cbN/4K3w2n0gJWts3
ZrmE6kv3UKsJh2d0cyPR167J/q44pAkDkexJboxviAfhWcK7sN7Em8mBb3VVSF3O
RP63ngBvXvegPX/ElzHzx7VItUBuG/Zx5LZjiSuzHf3Dstu3EOHtYg6M0IDNWqkO
YUqdhCPIHgAY102pbp0hJ4/CPq3r514thIjrFcznI0K7na2J2b7yE+7xxOQMZ9fq
ce4DtizXm1VCfL6MUxjRBawjHkKv6rIwekeIpJOZHGLsxTqbHKJM73tywEnWLX42
843QMkNBRMRbqN4QKAXwJ/VmStOnCzxkfGhqq263rjh6u2CoW+vMg+cSY3yjis2D
lIO2yvQU+hkPJjPUoW8kQ/sYyd/LmjYg1iB6zNLHv1GvsMuLKGh3JqRj1q29iYRS
XV9Um0T4gE1lDhj6TMb1FWLminN0TBEqL9cBE0ILBZu+jYVEYZj5ox5AE7fygDG/
h9QHe4q//nakAL8j5cJ30QyTrBRmzMLneeCZ2gCFpnEfy5tb//W/+9C9AeB1oVl4
h0/TyBZNOtK6pkcPI9fpex2M/NoFWiPdF1R2DWd2pchGQMXdUHqqWKLZlFSWUec/
7AiU5i9x/OygZcgxwW+RWKh2vlq0yjNdr4CTBm1uaR9i+if6w+Wn7sD1WtiZ5M6f
Ds27FKtHKLP4jeFEm1WAMn8GXh92Zv8ZEZp5aCykrr7zGU4Kd3RD+zwPmE29Fo22
6/7gsgi4sFAqBD3phdYlBzXI1wxYKIxU45QYWrOwKv0hwGXY188cVJqLLeamprAi
6fpjkXTU7SCVFHHuTk4micyjsWiro3KZd3uXcN9fVSM/OdMjy4axBfSk8O6eisaG
sGoQVqtK1y8lL3a2Bp472lTG8LnqMBVLrhKF9eFGY6GhHX0MQLGJ4PJVORhcOOzU
FkpUG/RPuzOHKNutyOHsfMhW3WXUuUnhz57z/8uygs+KBsvtTeWsJcn6sqeM/sfy
cewCKtIhhuX/aIO1tgo8ZnRD9SJxf7BiMpJ296i8Uhzt9y0o/d54fj5R+bvm/XDa
+GZpfcy7FEWPFBIemphgomfi7xfS0Saz/4mDe+JrdotcInmPcaiVoAYpInLzawcD
5tc4nHSVpNEmnUX6MVHBy8hs3Vlb6UyzAUn6c7yPkAuAxd4nASlfonkwo6BBI9+9
I3mhoYIrNFN+EyG0ZeWPJyFk5vPNRkdCstpnBMtVORRxixM7IsgGUfQ9EbFWlT6V
BWgFnmuS1a0gGHhS7Z+rIdVjZ+rBPcKdn/fypuv+tgZ4W5KwZq5iOtLbbivD1VSn
jiuW5gsSCSQTwPf+hEh7/jHz8n2u2FQ/I0yw96U8fdt3bdBo21avIJUsvIbC944b
5PXqCFP7hON0Nnh0sBkmUyN4bY8zUVsMJ43dMW4PFb98mCB7dPUe3K+vwWwfg9+g
hsJUNWTm4PlskjWy9qS07CBkFK2Fg1a/dNJ0/vCrh50+vyeIKxEUoInZEcwbxNNe
r1Advbut29aNAR25lhhxWLXd+LKAHUrb4jrO4DxzClyJHFUzlfYGVHraj2cHAhNf
M7AXX59MzwC6dr7QvT//i/kbLJbsRxiIbRzvClQMV86EytpjCJvenVwXWcD3RQl6
HjoBnQaTUatgcXP0ad0ORF5I/o88q2P8557NwMat/GmkBgIg7rdQ6W/SuVPdisiB
O7Si50zn4bcUNeDAjI4qlSfooeQ5HZYkVpnKqBj6l/W7rYcrEwZns1SqAf7UWdyZ
UVKqoPn6tGCP+RQGMcOydHw+tVyX3dpfVLWK1LV4cFB0WDyKsfe5XvOzTgR1eGPl
rkqKXiNtpoL9KDxTXnxNY+ZrWDByIwvr/ZBO23iHGiX3ax5ySwQAvoukeFmBmJ73
rgmiOSMYDlWuuYtL/jV2Lp2Z3vSN9j5bOXQRlq+9xB4GuSTbyHpuRG7IFGcEmWYa
7/VFjD5p26AOUbGzQR8lncDk63EPiEyPi35tC5twguOxGcaSy3NYvS/ijz1scaif
eMjZnbdPDjq8iw0qOY57uqfqSUTwHVzMT7Ecy4ndUKt7FwrgxKZcQ10gHS7XKVuG
sgLJ0WYXCZjdPtIP+O7dFTzD2EOODdWgjlRF4rxT/rWM+oDcHV4YM1dugmKnZELf
AE5GV3y/Sytqyk/JDYjcs93ciipJv9CgJBkRdXdAuNhO0exLHrjyqg/p608CC+XI
RKpv3FLeTgs16WLkKItNdASRc38ZWFRHfR/MMnde6ZzZkhSb2ZL0ikfTL0oJCeJ6
+rDZz/VcT5tVMlbb+LVx9rvyR+Lb81lptem0C8om76iAmlMxt5dv9MedWofLE/qF
WeyhA4jqqEnmCSAuL4C7HAYONiqy4PINfJG0wTJIHkoeDAHjEmQtFok1NgsOTbP/
01pPQIuN0g1nCSOIZTHN77h2SazixHN0+8RQYh2TCsUJcz7eEF5IFyqTUj09Vsnc
Gy0cJnmeOhdA0s+I1u+8LpkewdtUI/kfEfB3puADA6/ZnB0E+E7Q232wKtpTvmOV
Bi0Xan1ZDxhkHjtVnLCHEG6tfbD/ZPqCrkzATm4SNF9Kc4rOGP9D/QxFPIcDP9/J
WPtHkP9bcWE26/eSzs09LcCdpebfauHoBhdVvy4eWjidCqB1JDdvjsf4ZsUB4d3m
SKdFcAMNc8GcICIDUCgRIxkIWfzoDxxdMB6lpp29XFOhQUehFYUeExKpAmdz1XW4
Wmb8W1vwILeFdGgKBtKsnUVDf/OCNLCBeZeIXhDl2MvRPhjhyOj/IDlHQYOfjrya
39a7rLNL48nvW2dfR/ra/Z8OqI1zXZ5brUQV42RhlH9kMZZIcIEZcopd3JvWGzp/
TFMLIzrE29ZFffAkynfYSmfDVuiDh0KbmQpeX5CWQR4m/vwIe6/n16xNQOi2Ad7z
2DRmmybnN3PGyFwgOCLgomzxImm5zvyMLeVLnx0BbZKebravrsV0ji001pDlv1LM
6M2y+whNSYe3Kk+NW97tbkcXA3H64EkLaF7F4aSB1B4pRKYtcvvGMQwWQjUZimSB
gjf8AR9+9HlXDBhVbriB1GBNUuf9mupEzvRhsrveHV+bhV0QQP+SJJtJoDmGDKWm
mwr6zjNvUzli4HjvZwKlJnUfOGFlcYPs++LvfTzFTkmp99UL2+JotHN4NJuKyjOK
rALpKJPSjXrMdpdG/3fOhK0Jo6FDdsRFUp/b6ERylAPvZxZBOQplDU63YUL8Ffsp
UXJGJ+Qin1x01LryaKro0QuJZsxYbows77WzthANelMU1SfSMeuH/++2wcjih7L5
t+vp3sKRQcjDzhhe/y1pyAut2h/sVbliS1+41SkSvDhOUWO080M3MYzAvKmtgIxB
KvX6ar3U9/zuFKaq8/PmFeIgUiKzzR+VEE8PSOmN07DzrgPC9DsV9hWYG9sPhtQM
B/RFRWwY0uDjbAhmAbZ1xpOkmvU1WwmbKThlSBNinkPza69s96IzDJnAWRIp7vqA
E7/a0jSc4+b7g/gtVO3741pzxEXuAIOcTrl01hICibKokgaJY31r3J0pcc1FV6s2
YYim8iEq3nBIXxabQ0mCoclLl1eoxHg4PSu40e4JHyI74F5wcLow3bWB7NvKAw+k
lkvGIRV2pq/i49B39TfF8lxx2NUxHeRtmohIEXhLceK6RezWuM5PnXyQY+SSYLjE
UzFD5PBTwuTNYScJUKs9dqBMQX4eJMfAgZ/FeNsZb1VLXdmLL68zVmanNR3pvqs5
G5xFO2K8soi1CqhyXJqNqaKi5sTVOpnJhUAF9djvzKYAxQptivowfgpYvxZqnxdG
MC+9ng7qaLekbsUt0/wWVeQWA6Pq2C0jaEHptgoCV/FNLMEXaCkrj39XUVJ7qaCv
ZOfRdHPqFCXjYSn8meI18WqF7fPTVZBNbjvcEIFjgJBZtb+LD8EqVAq6JM0485r/
hW0+3F5H7VGySgAiz3qj/UrmwT+BusaIN3tFQEUjrf6cX9XDP2srTnXk7vGyvpgn
pReBPjhMTQGc2J0i0umycNC1MC54vdDqB6Nh9GApaXFe7uF1ewVnsr6Lk87D41e5
0ibLQPdKSUJXQZENQPKAf4Z8Lv6RgcdYk/KnT5kK6yz2Ccg1V4s2dqSA+LTw4FrZ
J3zPIaXWNbvc2vSlfWpjEQHEWHiLNy+QjGZu29mQmKlJSwHMnlNyGDk4uUwpUx+V
JxAx1XjEcNy0gLOYH7lKhtu7kv/3Co2IL2cpQx8yKlOfb/MJWlYq4gUDyf5ByUdl
oRaCYh5i+YSC1KHaakgIIbRiTtPFUN4JcGHMgXMMKshwPffTYT5RlM+Y+eHmeCMl
aEhbiHx8a3TLjSuSDQMR35sJ66d7/z0y9gJop1IfUHgFvkd8AhPeJPCmvQNmlnb2
+LiNECCKrehVjKRCmk+yNakXgkUQ3jqfnIhgAa7hKMiZc6JzyDIequear+B7Di+x
bnEUWLydNPOy3cPyycSloNg4S8gd0+GM0bV/2Od9DA72bCiSXS8eY/jNJhl/w3aT
GQ4IbFh5e3kgkTvgEWN+beDZYcJtfmGBXKKYEfPck8dlzsSmwKcvJqpMIYH88Qx5
7XOEposgQDp7xFZjA8zRNlRWakXR8PZqu3TM8dwLxj+/IOFN+UV9yWqwru/n84VC
uhCKa/fDxl8I3i22qSWiwS9FWYy/5zsC35oOzd+yuT9Q9SuoSRmkxcEzRUNU6WDp
xutbCYKmClBVRA8vDO0ZEq8YpYNB3n3JPqYQms3vbTzdiu49AsAKwHxJcl5grLJD
PHcx3XgLE4c3PVTsMGhd6R9IrdzaFBeo0XD6i84MIljm6SYE7j4iVOG3vnKlMPe2
DSESVfRN02VfrU8yEM1iB8mWD/hU+W/X3od913L4UzYy5EENKOh+cL9ayd1Gh63B
lXSfz/yqWQ9Bv31rV9w85OphTTMdGvfatXYbHboeVgVnPbXEuRA8L5dgiAYXCZ1p
Cvis1CzFPqpz6BtqO5XMNx2hg8KVG2VyWzGiIPjTdjs3Da5nVElD5I24gnXgsoSN
I81CNFqhzOVWP30cmJWCKYWlYTGqMJwyYkFtUXYylwPnkIQagTPC1XTfOxrfnYcV
zeegliM733o2js7xtHclfK8FU1nUQ4FtzNspPXecLr6j9O9u0qWnoe86LpDlMlyS
+V0HvsI751WZ8ELqTI+o9UdGpDDLjGety1B828AKgK3/QCLR66X9ShNN7DErpjjA
XLtXUPrtwgIdSlD+PthKFPF4NIxraPXvabxgTYXWoU87la8nppVyfP7W7RZS108K
M9wzy4Rgl8sbsuVAZK6mEGxtI3gvUWGtcg2r39k+iEVBlJVzM89qe4hQ+Bl3hkFc
bY517//h26vAjQmi7m3MSZN1g8C54bwvHaAwP+CnyrHEqWbhuojEJyXlub+ksONv
D6YaIRzZ6ujHQ2EEgmofxCNQ4Vs7qwqc6qEF9/0S9/u2pckoZO+XtVJ265KiK6kI
ZtmiDMUoX2QUHtzsQr2vrMDg7Hv7hBPQOfLd/HPafkUTDAuhLR0UatatIwq39e2p
OMIu3PcRE4cBE5ZJAzy944WgLuwc6sE+8tXdUrWtJwZcJ6v3klL9dA1vU1CNM1/g
YvaWZwivifXlF9cJeTB1f7aSR/z4vEWJWJgLYgQuJ7Xbjznd4SuWfd+DyuJh5h1R
S6DWf74e3YJGya9xtwnAy2SZ38a4VmmunZFhJ8Vd62TBhXC+uVjT3o8Aa0+oUVOK
ajZg5Ef+cdD41tFDFYbevlp07QyZTI8fIqozIaF7lGFY35IGoz5cjloVOaW/7Z8g
Etj+Po+Ydy4D7v7ByKa0yt2wD+ih5vTLd6yYD/Kg7mKq8ZdZ1IszKweIY0qM9xIO
unTAuMdVS94bGx+LwYWA0C1vbj6NPTglphbHNsE8E2TkHmF5440qsehnzZoVWRH8
80aeb0S8negdQeQyhhOVi/05KoZ9J56YVeE4OCVoQCiB8Jer4d2NlsEGO5PnzZhg
nLryXwWPCLnP5xGEg+FRTYAc0cBQUYwKWXbpLDLM2pL185Q3bzmln52l05ebJYbD
9S1N3iXKkxC3fgiQei6CuwNx0sY9LHYjnj2bNYReVT67nA2nPiVhZkA16i2Qs4c+
HNeOxa2TouC6h6CV8agMtsyuagQQBi3I7FshIMgDzIQr6F10/XGxBMw3+pcGptcM
GWHDVA5MMsd26mq9hWvoWDFTKa5828Tng+LnK8Fiz9tcZ4GtNf9BfXw7jC8mHd3R
pC/jnN2xM9SZ9CJ1EvbFcf5jBsaAEZuXou8ov949IKvxrj8cnMB9y/8Q1DKggpa8
60RtNcVUkXGHo7SKnA7LjwGR5fsw2JMgaPbiD7yKs0Z3EpqsSgVnL22kBBX0HKTg
UFjQpwy3bAkmzsN7NRLXmjUtWFMh58D4X7TsyWX1mSm6rLcss7HFpLpDqJdAho+s
n4LOXcEBgGl+Dio5KBhiAhc+1HuXbi2RmqVtQsz8p2XXKsbzShLK3Jr3fug/6uum
oDkutJxnl8r8WlxHFsodbeWQ82QldYCWSyFcXxFZfFbut0EYF9ijshOmkaFEMbb+
S+oPuy9XicLa9GiQlL/4zDn1sRE3783D+GWeDSrUotbMc0Fzskx5NoqSOERewFQV
QBYHLMjtuwgjvmw5vWUdsR8zTd7ZUGBQdriK6cOU7SByZH9isKATLNSeNkWG1b61
2Btpl+5hCNIfbdWRV7MjvM7rplzbAONMdcwjphJiLOvMSG4zhECLtqtuBET1rMFu
uX78lQUSVMyGKsfTQGykBaS/6+tUmBZlTAd1gdWOYgzyIyGcJzdtGTHeUhTvNYI0
V026O9MZnMClw7ZNYcWTWXrsYEmVvPopCvfblai/fGdbyYhlPeOBhIGiUCboDxZT
c1kHlVgMRsfBH2I0nH+rP5fBmLMIcKJ+1f+bPrzDvonaIgb2CjYxIksCgENEgHg3
ypBJiOUmoGy5FeQyadBfahwszXB1PElcFROPpqkD7jeJRZ+AkE5a2CnTvmB9XgFy
XVMMSk+Za3ItHGHytmHgEg5CH43AcNy5xzfqXbSRkuLZqU56ZQggddMRlLui1aQO
dFxK/ZHyUiTOQngfzEkoEmd2TIokKkUKNk+yIf/tttJPs7ESaeVlXyMvkqyZqb9Z
6CFoyHB9yD/OfyvZ9I5rC9KGV71Cn3ySJ98hJ+pfDh7w1rv+4UQIRn4gXFI3rSIF
p6o1Q1qhKmmfc5qad0QKYMgn2cTWIXPggZLTUB/sVsJ0Vrm9q/jPx1YsA8/YBAHd
xo15BLKefgKaxR6fWvqtLvmSlJWW+mMI45Lu0OraaKF6YCnhPeJkum48alOaGltB
yqCakZaWz1uthEb9QF/sPzYVRMb1ictGk8GugHEazG5DetX2fm3uzwfT8Qa1coU3
6GkhAr1AjQDiKaxbg2fhOtJGRGHo/wu7XVmKrEBMEMA+rrKfke8vkbUaldJy4brE
ggs9DRg8IXKsfFTqZb8CtRjhQ3jOcrMhTf3eK+sDmMcfvjS1HgNqprpU1O0+ukhj
aWZ/hJGbx/33PS33Py3cg7ZsGNey3iXNXrP9kBd+q5VE7Own1lYeiWaOWcHB3+Or
FD67P73mIpXCyCL6QaTrls/b+DcOGluhgc8iNiVRyAfJ7OZAm/1yjHODCxrmnpsx
sclOV5fuM50P1rK0rOYzCLONjRZJxRpMiCeJGhFOdm0PvbBkcM2qqir8D/klVQ3X
jXG/clepSSBAjRzbbJahMUMt3yScuX7zgu+MSKidKVJA6Z7YuE2S2yBNOMfh5Q4c
k1Au2594+zF9hFWh8r3MNiOTmodHCEZeTQQV/VZ0DuUSxKtgUDF1gtnJAAFV2tEq
udqLyjxOyJ7E7z7IR0DI5UKT/4SwtLcyed7pubRHdGE0V0WPQT3QP3nj6izwcmbK
zplPfOCKPrDlle66IUBpm0/eGHfY607jsJ4NbXpZOQqpwjn83K8NkrKeGGZya4EP
EQgfO+49yidKh6CUtBwhNaV+0PGeMocW40NMZ7aSfaVdW00/w2UprAXp+5HzxIpN
3K5qSGBXQ3ml2bvq8nTAgqBI0jRNh86ROKbjym6zAr1YLqnjzv9dAAcPFS/QQEES
17318H3/9nDBfzrpZex6Kf5Ny7TjxDn0iLrfBz0EkwdCywXTC7t9RArvS/4kQDG6
JokL4Yda9R5JjBGtVqJlUQ6r7r7CP5tW+Jg+mDJpVI2GaY0AfQ5aXawto6RAudyu
1MLtMZ17w2i2ZjBQiJUCu7R1TOkZHFN2XTQHXCqp6qp3TVyB8WYN3310CqO7MVTa
/zviDE5mYTUDyN3opsXkrQxyecWcXxKK6mxeaUPM7Fg6D6Y8ACcnXdN7gWxCkjDh
uG5BaWaNbJQLfGYSYWMIpR1W0W6xLNRM3cOg1lJG+HZNAC8OCbUmgGtvn4hpOzKO
WIoz3i17WNbMZb3sC1N1J8Evh6fovkAogmqKl+Q5gN28+wMc0JOavWAPLpQZdv+j
bFC8rrX8OYtx3FFWgZTnpabJi8Pf3jf6++otgQbX7qxyKG+GH+5zDwgCobOCa4+T
S4b9QsFQbFGs2P4L0bLtXtWj8w+aZfjaDgfDxHsZe0yMRNjAUXplRw9nWeqKq8cY
pXAzs7ainZ1+YhHslGAmEnEki0vDoUxCRI4nFMc2EBy0/JBZKHL+Ls9y5gjAljGG
fMcDa/w3bRGww+Mjvx2ZZ3ntAencAxI9FAPuuUPcvgawVDdXPf6ukks1FzsQqp6k
U+rm+gOaNgbB0X5A6sup6OfD6rwgr1uTuAQqH7zdbbizLevBX9JXqSLpbYANjf4z
ry8kDYQyIaPzEASFiEh2Mal6gUsC0s3QwkatPfIuyE8JQVJFFJSZFcf1y7coK9Lc
Wt1gKKoVS1hg/qwxYLvE6tTwn6yeJFEqhg3LcX4pcIzHCYFt+zt+YTUZNqC8CAb5
Quuvyv0fnEcAVzddrydpyWYf/qaBtd0CbhyLyjciB2mUzS/kOxqWXD06165uWKd5
PGUVr+Xed8gzB9NUDNSUUpnd9i692C+NPZ7xosA89eemav2QDvnJHbvfHedHDdnI
p6XE9yRyD9RcCZUXh/IrAYLmHnEtPre81vnBpiPb1f/95ETeH+c+QfGAeQbHEZCc
nBs0PHdnQjHWO6e7xDPtap1+ie6B8PQNJH/osPlDyNZzg1BlT/i8qtFqQvnKm8Fa
a5z8DqXUnrVEWEnmBgr9E76VrX3ZoMKidQryGSqy6J/m5U6ZwQVUB/bDRwgstI+h
/xKQGVPQP7y9DCjv8h0VShfoTw8+pgp9S82I1YpSbsK3vB3JVyTe+3Zy8gEkfksZ
ptK35p2werdVPgR4aHX81k3GAqT/50aCOldvAOr5OP67GAhP6y4OmZyUSBWmJWww
hpwdLG07JVfplcCX9PsK9lWl7V8s/di8RpSe/XgJkuyea+HxfuHFdR4eX1BK2/Fx
07eGB0+YYPAmcjS9/9KUefQf+7If2cXwO3pCfYWMzjNmwMxgyvNL54h1DtY3gQha
1XUyIxAT+oTswIBXaKRbp/1ePP1rhEVILyPFmiEjK9/mGAV9DO7/EeK3ZUBIAlZb
y6VaN5HbGPeyWQXrc7pWjj9zKbBuLd8pRooW2D6NzlvvKsH9AyzGSW73gE+OEgSz
wuhrt3fWMiIhO0t6XtQiOkyJU2Xz+EQfeAg+NNztIRlT0m6Ai73w+g6VN3f+xLU4
lOE16mpNBv+Dl/rMVg87VxdoBekCGtaCdkrPxTcNfv/ezvsakmEfg7Db4nmMR9sn
lqL/MV2C+Tmy3lQuwTeQ4UBl9RfIQuzRWMniZJSJfS+H3gAwZdUfylpMIViYuMnQ
B05L1e6AIm3q1ZQkCtfat4wB+2Jlm6CeBnvjQwmpiz8J1b3z23I/iCXe64vWhuFT
uDuWzOfdVYJ8DIFXdnOVbdPXmy0RoYnBP2DJBYFZzki8YKQruWrgnlSADxt6JYz7
ilCjzrjDhJDBwx0J1HJT/4+ovXhPlKMn83mNcyYtE3NmU6iLt2Tue/vIyClFHiJY
6id7r4e0l1zdpu35/P8uHmaj6ffT8/f4NL4oUttyhOVjk9NrWwimlh338k2euq9u
OezpexLxG+gM8F4mlQkrXom0bPli7s41OhuIHXnSfdZcbAeoNIXfSURf3sES7I+q
JiHLk9rCuvcZEMFO6ccxfyyfj5NY2UPdCByXQ4+zJ/0MYWGfcr4D3ejkRxIdoZXu
j9Rrl9bAPXWVi4ak5qdJ+CFzmY4KfkcGRYdezO0dgbaHG6UvZQkZ1HczOaU/TvBq
GN4z50S5nR0Zv5d7AgDg7azDzM1qnW8hfrQu5J21FOdLTOgjjFgygiktcvVCxbXo
IbkfQxj15jaIj6l38bD5jV23xXEPx5O+6XSI3fYKxqsRTUVTctPQu4rIoOFlJmRn
5Dr8yX8eOq4ve6+bSdkayD8Xy3MI3deL4fyIu+Mwm81KfQTAWQ2R5bICEh9sKpeh
PuL+r04sk8jyVjlI7nO0epPbRTF5wnoutnLksOuD8pEwG5Dv0yqmKlxndpELbnix
zPcOLbh0juz/poEjzWBvNXxzaJ7KBubu9XIxVF2eKvAYPCK5mnkzHATltsS2YYpj
1yQjMsWNOvDNzc3Qkj1mqMC7jpcZ8+ffp8OALGuACslgfhDl/ftZ7IbZ4eo1L4rh
ja59mMV0nefs7q9F8JjKWVKEIDP88sPtdQ0dIITWE+fzEvxTtOspbNBhi5Twzccy
xYKSWjpicylsAMUf4Uwlw/0lGHAtKD27cgSKPA30zEhtiDPHo5nQfnwx6mIOuydG
l0yqb5jnOzB+SWsIpNADACLdDjjM0lByWiO266op/Qk+QmfTsk8Q76FuzYuD/rZ5
R/flFrDv8Pp8ibWHzBCWuUi6AbPc9u9XjqwBt2LDF34U7e0U3pjSjkqwZqBAqSdK
lIspDEzZ2AJWP8RevTciJzm6P2dyXJHa7ZdcQpR4gO/0JYfMsI6XasNjFCn5cvXQ
WUE95k/+9cmNt4cNJ6sCw+m7soXu5E9VHV9TZeBt/Ew2URH9rVTH4rUZ85/O3/ua
1RADnbtzxVgDEX5jTXI8mY6VWodtIk+ULqgrB9sOvasBbu+HFaF6Oz6JdeiSFtWe
GktXo3RblR4tSJvadzzOEVq+lJeOZ2Xq88YPkzPepACrLDQnjBLnBlloDeBFVES7
qFNg85LMhV+/rOESIEzMHXvSojNhih8Bdws24M8c3Etw3AlCePngQQDnOgoQIOO4
y7vkyW3HyPPl/0onwIBWcwSKcMC0PeinZyloyv88NO724Q6jfyz5Cs2fvy17uIph
1FLdmqNMDqWHduN3mIBEXCCItB8KJonVY0yuzDoLQaHqoh4zFH/B3rPmv8fJNO0w
iNK2HoViv10xyq2/EYO7zoDcu50ZWw8fYpQbLjvEMN0N3LI4p0AwC9TkYPhdZPaL
jFHyA6nlQ0L/HrRke+R/9CQ0AkmaJLlTQz8aBuicwNtiUmuNPA51hIFQAgYyezHO
MDEZuo5Y3XZywdT8dVrkwsI0yK6Ksd03EsPRYVigZ56fhqKbBGomE1A94DfXOK02
4wzIYmhmi6OJ2PtvQ09KC2SslZLF5iX79lo/etr58laKArC4bpF/g2dQjA1Hnznz
BIEsXQMgdgtEBHRMq/aNBuzJFVsj3idZZm/vJsbdChsLrEiJyLIrx39ixUFi6XFJ
0d4m1Nfu16buwn52sr3y52YDT6197b3LneWR/vkQeAKrwtCyJ+Vu/ffHaxtZB77R
qXlr7vnY/R9YltSNPfTsYefeedVm7cxQ/hynjTk4YxVWuwuk7nmNVjtMjRp5sWQ/
ed9fvga6BmmKVCKdOFctwmjj403ljtdcukXhSpfDVV3dDoNKMLT7pmdZS6l0VtQo
AcpypSZTXiOkIjNSBM5apR/+eu/aDTFZ0p1fYVd1KOLeGO82iCJv5CpQsSyruk4S
L6y9RjMxLm3kxRlg5K89sFz9ZpRYvemDd1W9jElhsxSOwaddMB227TO58l7+S+00
l5q3CLno8Sb1JBN4G9SpE0vz3ZjjHS1QZzml0FRE2ytIIcnMWsAz+lJxWqgFV1Ma
iooVaMLTDbu4lFLdj3AoXO3ZSX01d5eFAIy8KT1tzx/bOd+KvLkq/xfuxEEb3a+p
+U0k6+yxHpAQjEAlvEuMeJg2K/n2QS53jZbJ8T944f7avXOvnwKgRhFSbs7sLKXT
hqZi2jElpz2cz7pDm/2RVLQHnbyDUl0yYqr7URUAzQ/u8YEQvKCz+nzTZd2i/0/+
0CTi+lELRmV9fdAHtXyMLtNO2gCoUOokwZV7PSrXXIxboBlYuINNargMzoePmkfa
j8fpSxIUdRsXKjQ4bsTMRlc5wP32iTTw7vDfHawk/IcyXC6Xo72Enpl13xdIAgh4
QpeEJVHrA2zjBTmwWKiHSHZ4bR3fQ6MsR+sujx+VO2uqiaHb35PLUeqtgEyrD6Vn
Eq7//Nm6ZEIY3Zkp8A53FRkEXTSj1fXncqJm2KSKM8bp6+FYVgILOOw4WdoU0opL
bOAbSsQjeWew1WHxGFU3fnKl+/TQ203rRYikJkdvWZbtUeYr6kXJRyrG74yNytAS
7QQmHSaGciTP4TECWtCK+JbClQX3ZD+6XpuJa08OOGiNiBDQxk5f3k65LkpoMkkt
9+8fgfraVVbvlVry3xIu7yZ0xmZaCCHXwCDiy6zDfz6UnFAoY4ar17Kn4LQxBcKi
7LkAYhbQid7jJqnxcbKxCJ7d2nigTGzHpJss1piwtnk7bPB9uPixakzydlQ5nDUe
dKNffk01nvONbZ0Ynatk/7Y0CEvN7PYy8KiWGN8ZPlLkHm+QFdz+ELkGggC+Gspt
yDTfnkv5Q+wNEr0xFZ4qvkou4eVJLJQKZ7B9b1pWy3n61cg73DksnAZDF0F3uWcs
yHbwfrgU4CnLRccXFP1T36wWJAVTBHs/UQrWg3e5+7I7uNoNqNqUmgyxot48dxZ9
nCZgrjN4yI7YEBj+sCZKbGbCuw0rn6pLM54KRIlRtbKQkXMAzlkV9525KS2+puAe
AhLv7Kd+4SpnOGjcFmdW/fdl4mTuVgA7dFCtowKUDWcWSPGv48vAtrp7T67zERWn
Vj6UvkQG/uOm54pE/3uyMMk/V/e/hO+TSzt9bZF9jNHGxQ9V/J04Jiujoclox9KQ
2DsOo/l+bxyMQ/MJbeEa8mlTYu4GzQ8SSR2ocslLg/bzoN/yV8g4yFcUODPo25Zd
sO5knrNedyJ1RKkf8w3vPzsKRs47xGFoNos2i9STGSrv+Fp5PS/lHiVThnELRf9N
GAEzGaca/pvj8x3WGQuAEqoNTXP8OAeZTFcAUXQzsOtApasuJ49C8f6JSYYisTLI
FpPPnWDXMzS2+2EWTDuyO3hTJRGTXjjw2/V1QWlflpvDesO2E+KSftRN4Qqa6OzT
gbWTevmWEHiJdp1ynl5+HTitf2MVCPoqy/RcVUQfA2FZd+nfUC/RWDtgNLcHf9r5
ESE32l2QNu8s885TdmPQC7WMBtAb1Lf6Gbk3C0nzdgDKqlrE6gk1VW+E4jM9M2dm
97sfw+0XSBPBwkhoWDtF/1cKsIxqealHFJAGKe9yl8hzK29AvcZrTCdO3JJpJRex
4ThP39y8RfiEh01DEfdS9+tTRVa95e4WQS39e3twAS9t9z944cqpVbv2lqfl4Rhk
Znp9weJfL2J08U3q9NeZIaTC6mjiLawT/m1JWB1Hvowo7nBRfJoxQgb1d/CAKjGf
D3w7mFz/CGwe4nhkhUAiXTZCAG7YMt1fGoTzh7crMSDf2z17ekOcfONlEWdU04tB
BR1AZlvS4TayqX8AWFpXQrmegTFxMQAeN0D081ZNYQbxb94KJ5QlLKYkEAFMfK/V
9kcBV1mdJJwLZZldm8MX8g3yvtr+iJsurj/76Lt0XTFH66POTOS1duCSuRRJtI+B
STQsRKDRCbchKcHBIrIJ0gIGOI81nDYSDtARiIFrQNsUszE7cm8b2Ofakr5M/ID5
BvTcaFFBKh1PBUn2usEZXMfPEb84kkAIJELDrCAbxsuTt6aPJ/bAheTzJw8X61Nb
krYtuCtqTfOvvwhYhf5Xg1JxZ0+iAQHYG+WUPsLcg2Hpglu7/xXV61MATL6LVHbh
M3lL9FO+xHGfbvD3UpM4RCHVWQDnDsAODYLjHmvxQJ3sT95b1U5idsrhxbsDj9hg
XCSMkBirb6miI80vLVKhkN42ak6G5eSjfMXI/7I74p1t5UGVHx9Tc0gn+M4ZGaBG
BmxBt5loStxE7zKIUJavsqiRQOCKGqUIqmYe8JccRdUQruDNLwe6f/nJsEbdnXNK
NLz/MoseZJ/zhjdo4sodLY2UC6CO2yIl4OLqjIQE17CGJ066Pqiw4Aga3G1Rfmsk
4FrUJGVis/lpclDHkE2SXGk3ppekEPQI7u9308PcxoZCByaBL2vxl9qUbT2unk08
rdlWeGChnryUA01YLWxdKha3ufTr5p8D7I/oKTXTC5slumqC0qqFiTMBS2SwHkJT
UBEGl5eZBMZl6ifNEHap1823NpdB+gUZXi/4QlZqJ9o7GbncWv4H/P5xvlOh/CFH
5ZnQ8/jxaMvJYj7T6qmjRTlij9T8gm90C6XwHxaHVGbKKfueXo43WiL/pzdfjxAd
Rhb35xfyipvz23E597+zZsroVqbJU09e9udo5y+Mmf80cLnjXVUaxau5vEnyxwdL
s5fqTcdTwZVE5pWCihoWDIseisevX3mR8ZVKGZ4d/XmJ361VPSXCJmlXip/goVGD
7gbJPLJgK1yQErK3kAqz0TlD7Hy2mB1x9MxeqypDufjCFy7faV8rzRtHAnNRFl9+
YOR7GNiRavri+ey7TazMw14CMuObhXDH3VdJstDmia4GJ4mMM3BiyK1BUAnx0sMh
EU4apbz01cXYc0m64JmS7SMvhO/xgGv0Ifp3rE4rRGPPvTdd6aV72upNjWiddKC+
6NCSjMyvloeWP7Gx3cHCv+sMHczISzscnIqCR9G7O5ZhfA3cREm02pPdZjx0dXv7
elxnMOU0r5JHZVDDV+RVGGA5/AQbquTVU/U3tRD0xcLcum8shWRki4kW+86pFT2G
B0QEb9oqDJBjPxT/jCa5bdJhBVJyI5XJzlNxnGQlGyHIOHFw+YEW29jJqWU4QFq8
R4CKUdwbW9iZuCdkytRNBwtM6wvifTtqU+UQDAD2e2IR3n6W9pdMtcFMhwYJQxpW
7KQs11jJfnTf7TQI5niFS5w8wVMEv0XIkSu1P/Z7TbqFL5wS+MRK2NBMboeBMUWP
2xjZih5/BtbgYNdEnuRx1PtkK3HRH6X9Pxk6ki8sRYRPFU9jcqD9S+cpdhIGTpRk
H65BWIXtXn+DRPnrD1j/ommpVSaeBSFCvsiyzhSV6vb1dhvdFKHN2sXdJI0yg81t
8sePvCNgUFVKDV+wbhhiI9efwaBKc/sSoldaK16fHFj0hJMWIvaYakNpHzXW9j9K
OjYoLuoiVCmZ6v38ARrmAvskp88Oa8TlSKVCmCNi6Ew5+5duIQKP8rZe4DdR3duq
YMkFYy+Jn+hv8X5hhedrIfMV2kplT7DcvY3+WOz7T+zFOrw4f/UmlJ0HkVeWIYZk
eV5YMvxzCjKyTkgOks+xb+Uc9kqb00JsrjKuy0SC8i3I6S99KGcur50a8tRBRFwr
TmS//CVQ5RtAAjo3FI3Dl4iSIG2kBHPHbT2SxZTnZcHoaIbgofe+Rob1ziLgRAl0
GwRr5SfwLd9Ts+wk6W6I3OwqRhBsMjNFsI3ZNTPvipm5rZVs/MD/JK81CZrXmNa0
IOlxjkX5ozvVwHgd9L8gJ5ldgAYqS11ulDx4sPiBJubcsdupz19Ka9eOfzBKDLli
2whxCIicfTL4Ucw24Zl4gs0IYgNiQGklo6eDOVdZO7yKTxJsKiYwNaXToCbsR6+t
y9KJxBSX4WrF69oX6OevACMpHmj3bVYt5MtoGrt2JRKd+i15jIKlThLaZ1d0Skxy
RmGh+8FJJ7BzgIV7FEAOHJ8i53v7Zd8dWTjejpoP7hpBMAm4r+sip2eRwMTc2AJa
uV+gUTXyxQmOf76NTKJN6KXxyQLc7EDugPYw/lHUijD6ytHhcWCAV4paMAfWUUoU
d7LRuU27mQT3G4Hy7Hacbac+Y8mmDcyFUZ9wIz2mG7xKXEUhmAA66NkiRSP/eSme
WiOUbPpfcVSltmsHJz7c4SAK9ulbShHQPDtqb4dsDKxqdkzgZpKx9Tcq9xqZS4CZ
eK1MKapIweq5iM8SFHqSZXMEDVlxKj+Cgo+5bW2ZhO98cjtONukCpIZhU7flb8Sp
LYEUIROdLVxGQjlzd+DfGCSEMp4WgpT4QfUch7pXIKrKSNPynNGjvPRMmZECOhot
ZtpoK+QblBZhBGuAda12by7/6WSrZ43goZKZUKXEh0djriumBpLHrGWFwT9q02SN
x0gj8RVgEWQimr2LZUO5/DcARfyJ3aajhX+uuEBioCaa5PLZuvzi2QzuwZhr3rS+
DZDxjcGQDUOru16ES6Fd6EiMv7ntrNLuKD/9+BZL8Das1rYq+6DnybtASopmTL7t
CF9hf9iF1avvHt2+HWLqLBNkp0x8OEF1sXN7JAnVfr4X/nG13+Tja8+OjlxhR9rE
na8agDTp1sCelxxmg6IZJbWsz9rGi7udq1/u0YlJwEaMn85Wod1fhiPlol6KbxAk
FtOFMqQaf1T1SsLiEdTPDd8tFlzaso4FRAIqDCKsfeBepS3h5pOityArWuKZJCBR
lEOU0Z8u/irj/BQQPe1qTs5Ai376teevSs43O28kO4PG4KVkDvo0ovpPvCYeZ77r
QwOYcXlw7T/STz5LNQ09jwE3q90W7vMzejYw+pu8DCzftF3b0RN7sMxiBsi19z+E
DWZk1HXSXPfHOYpzlF3Jlfm6pEcN36pDmRFim3Sgjha2zqJz3dTUbWDGAbuz1VEa
1Nc01oRQohJnMRF2N9I4Mbvpd7bdwf3zfWmioLEmoJMZcwfI/BSbB+wptXcYhEyL
PW+KGvLowgA/lZIxSKLKRj82fr3uJFSbNnvdY0CzgB12HHwkPSSEJW6itnq4rk2D
AkE4se2vioMBxFgdih0lrO9WzorOl76/UHJ29KSnHniZayvh7HlF6H1w2fxaDWeu
kgHKLR0PAymTk4bUuThdTGVMtPA6ClrFqr1xuaaonSr1b63X64lMUUbd5Vb0e/bL
lsZoe8ba295SYngt6DuadK7bCEMoHV8W0YObTOCxw4e6VRDsA5Is/g6aBJBnqB3n
bzcR8MZ2t8mUG2Xv44ddXKfFGDcxM2CgTidpLU27M42B3WVXIiJLddWKnuzQTNtY
qSswf9gu2IHpltq8Sc+q2yhfepCLDRyDdh4CkPtKEZ/GY+4rm+aPyuh86B1JHabJ
WCi1twoGFChXB9NyVXsKeYEMAcahpUhiETdHm45a3zdCpdBbuLTwsoK0zFJSxfqS
xEb7HrdQBuEAOWExuZ51B/fohvCIwphp4cCEPypxmnYyjhAw/bSPhWhYztqE62gs
NZNW0mXFNl2kH4KLa0752F0WwKY7FQC0rXfdBZXVbYtsAEqt6IGU1PLZFEfBqkZO
H5iSeSjBbJ2AGD/vVAijzwiXd2wmCm3ao6Q94OI/n6c8WLS8MxL6IDwFMjqo/Xci
aIxeT5OMSyWBgDHuid4aVXABE0GzsJNme9ykobdy/mFjUvWFM9yvCLZHoUgwWLet
njgt1vmdR1gLaQDdpO2lCy8xGLCcbqEOFirVcA2YnDS6iuFjV4L8dMk79y9bVRjZ
YyjA39IaygG9jORJaJxxitc4+g6+40ple3RHr5hRmiWos6Y/DMd8fZ16J7FLyQoh
1IWItdTJc4A/LU5lqObArUkBGx7iAC9jNhTrUvDKw3+cEpIInb0FJQZRR4dVbK7Z
4Zy/jCqSe0WK3S+Al2HG3S85LESa+yZlOMbybYQ777tsb+bjdf4A2ZjwEtG7vMBi
TuVw1f6DaLuFQUrwD+ocYhBidqhUE+IgRr/YOGh3ohgQ+zF8kxuUZY16GnfH8jRQ
ep2D4ZRJ86owUBGy2tCEJgcKQUrbcxBohlVZtsAkDXrukL7Ajgr1n2DT1wBOT3G3
KcoH1x2Ndpq9+yeBYoVG36mR/mGSyV3UZcGz7XBqM4Ya2gAKi83PRwULhJoUF5Gj
ePftWJpqJ+WJmhd5IxgogmRpnqeCB8/sUjtE0KA2fjIDn1WUJ5uuq1tpu3cqMgyi
HWXT0CBqMDMXdn1wvRLcUf5XDr+tlLtWliK4NM1hhNbr9YWkw+1bnWbbtoiH7D5j
pG5+C8u+FcYv68+Dc+o3iF2jCEUuBnAkMo6oPFZJP7/YggbLJkB9XP3l4LEpQt9s
5wfPt1WTny27tu8DnpNUw9/FuVJ7BNPUO7J1+S+xGhJZbEuEd96aGmboiQfIXc7e
JgHJ65TViOPa2Rma0GsZan1T0iTYQDO5GwjTFCDqc7uoD1WGIbZu3loR/aJc613q
E4Ng8l+PhrIO2RahCM1OSR6jp6QagcdsqXpjKvDS9vXqOQJ6g1CwXuw4+XHI+p4m
lcTEYJNifpMeoHaPxpaHv2t+MJnkbRmTAHC29dmeSw7DFAsEsnXGS7MM11Gw6kQ9
kcCDj/nBDlkWtfTr6EUfeSIF1Jl1O8q52ahZQb4/7kubLRPsLwJJ+HPNVKgFNWvp
xwF8wIyClKpN2Gw8T238bC/wtp4HhiVgETXR2tExXgJ2tOm5IYDPSyqqMzcC3Cyl
8cgbo7M4SmvWWtiv2oq28mSKR1QdGA176dc+BZ9P8hTnvyjZ1WJPdrFOeXXM81GH
+eJ6xmnL0mJVXh+4Gba/7mD6owOCU6os8vXwB/Ryv+ZpD7wS3rIgbxnfSmfV7T7m
H22c6LgN6FQclcs66ZnRBAxK6oG7mUp9hTxaHaVIE0/OR90iFK7Zh7c7VEn6EPWk
QAfsKPyi8ot2X2j2c3U7WQXKjieLo0/5x/ad1unlKcgs6b6nQbbHvDz+b6yokzFh
UjJKuCiSkQ1sZguJgW59ZtZPP+PC/ySViZZFq0YmSbHtk20efLxYN279P9igGVwt
KwKJkFxqEJp+Rtha2dcW0oWrIOAHLIIGOai+v83Q12GlYVYhG6awMbmbukkEm4IS
kP/gYb8YSwXlmhrEDvaRztMun2JoM0VxHGhvrgniEl/Ydhe/wLtllZ86HK33/U1/
52ToHALBt2qRB5HZZV70BkAyjL9PhJ7FiB07R72r51isB73fgB9bUgNJJN/dhTQQ
mdOOIGhqRkk9KVdOmC0Uh2NxEMlwLt3dD33arG3HKpUJHzzKsTLUPMmdISLfvf0k
FR/3+cDy1do3bb9Sf/BY+o805cNIwezdtV9CVBK84qrF8hkZnaTXgu07cgFE1hfB
plO3zrxWzJdNoLO1h7Vhb9bHARBpHNFdjbKcPNQ8WFWHQOs4E4NPz/J1NnQFGQ1n
BdLRRSjeEpg6s0Jtt7KnArG8BSDuopAC+0RXABP2AcXe7+YAAlYwyuMJ4xFbYV42
2U+S53hiW768338/s/DGFUCzrb7Vq+dtXQFRzr3MSLhacOwGCbRXJzNqKGlxMIa1
jDPyW0Fpx2MMbSZLZ26d1EIUusChim8c4lXNKDCnHKlKPtaX3ZxHw//OYJX7PVTK
t7idAaK2JyNW79mJ55N1KNOuI366Rh/US54m280mH+lxImgQKgdY+YZGFeYphtaS
s/XkGuhC447TXCMsFRNQ+bNiMAQfOslGAtIZftrTZWWxM23gx/WCauEMjCfKSzcc
yBThsk9Yz2ZUGnFZ/ICB4Yez/3Y1bJMFBBve9ZtIQx9GqRH2Y39ewcYxhevdNNFm
qo224qV+e3xR+FiiHHzfP2TlHGA+QnFT5x29QVHAmy/GWlGqlj4H5P1yf5hXBOSv
t4k8Kx7qK1THLc2hTavVuBu1Hop081Wv9k1mezEthyAxBxfo3izh6JCxXTeL1aBr
FatoprPWnYh72J2INMJePwPLT1U47zQ9hLUbGuaWKlO7vMtSRpISULmcYnF6OeOw
ZqNzbH+j8sAs1w2m+/ITi6SzaOmlrD+K2acs4fPB8bHVMNcmKnZtOEM8POuKxCEv
XKhfQvM++wIrP73p8Sox446qow2uK/w5hDdc1ZsMnmUUj+5egoWgt/sGAHclyseM
qleX3E0s5xuELzdhlhjsltGpSgF7jwXp39UzQAcFP/4wbbqxbDXJtj+R748ZDB/Q
kxeDqwMLC6yvl4T1v9BuXXt83mksNr7HGEtoCbMYX8dHsvmicA11JJH2XdQ5+ZWc
63a4VxRuxxJHCJC8fss98Kf6ppO05RNNU0h0WpXrszZWtR88aKgtrOtJiE/ylkv6
AG83/qpk32m3A/f1c9C2pcHNEkXEoAbesX1J/HCQfUg2lIfC5NT/ajCkA74PlR08
9lD68Iam/bOl93QyNiH4zEH2Nbe3uzXJWtE63Y7k/kYN1LyWuQpVEw80ZNTkMJh7
9ls064hUOaurMJ+HHQ6Bx74sk1hiCH1srKAcfbtvYAd53fij0MouxhFUGgPgDJgo
JmStRHxA2Weuul0yHH1jSPyUprFkmiX8uX9WaRQYSbvJYBdVfu4r4DThg2PkxCuw
4MEo6+3TtefBDiP57EkCi9gIDT8Mhfygy2ylwqzbWDCEjJFNmMNzgy3DKjfwu2Ef
s4OXlVa6Qzwn0YBqcHykiLDlsC7ekQdtABQ65Ecn5EpquYHTD8SOy3Gq5b4JQGAO
DxTxVYcvdUIwXfsXH4y3JZZZQTgtl9IalPpmEnPwK8dyPZzBUJE9PPZrfcB6g8oC
gYS+ekJIo5wsM/BZ2BRV3Z3OBDmYg8Fm4k5cDbux2vtdUAy5u/xwW51Pg2TBd36K
VmTjyAObs1qNQnYOcVYtqv4QmrM+VJPZQaXBhbmB3utUszquJL7lZy0RkOrwKny9
9GAU27MmNlCe4ePHXUV9rltY1jP/OsIelD5S1lVo+DBOWu7kUmKCwsdUkQYVNTuX
/XHHA2P2txciCs9mef7B2GJ2S4vr9bVUVQ3+U5LyN8yXg4t4CzcE1WHIl0ebSIlw
Agq5gMJVmMTt+Zmk+10lZyunZIYeljvlPo1fhoN70S5/x/jmopZfPREhpH0MjtAX
EFazz/YsW7BvKf2DU99tOnFjo+6qKrBGnmJeDPxAUoRFEhCGyStzuJ8BzRvm+H7x
9X1AA6Ih1DuK1X/ieq4GpGJHSv2FVRaoxbVRPviIk26DU74dT9agvThpvXtzZBJ9
1jsOJhaRDj4RKWCdP06FyYsUE801BstGx6LIZynsp9HAMRWWaBZSS0HduCiSkPqY
v7KdtJV46YuN+MRaZszTkA1W9PxgTdhQ1QAsyWzCRcFq4Pems9h3Ebo/IfvQ6Gvc
a6RXuS2+ooCYmTKdzkVJ8fCBsD9ReVvM0vNk5zyuHFtuHto5Rbyo9rW7ux0mKxrN
Zn4wfMYLUq5MsUsiOBd33o7anc5/V/2bt4z/0fxGJ9UF7Z30OCZJ56RxJsDTIq5e
f4+VVTVJDlkh41TX1WWjaSyxoUVzYfUaW9+oI1WPM7FUVE3Y6ggcyiTaZvo5UsTD
yIzGKqdlxf6Hp/L1Mxi1Jqw76cbGjqL/inF8yJAiN3hd8jmOIpx5jpetUZqJ1ovA
U/KN9QZpJEJhZZj5vjrj4uZ1Q4I5znI9Tcqd8FuuIFvkTajAW2dscj/z4c/9EADx
cIbfefiLmr9zW9asp512dgwrqGPd6MfGy+BEyqx2jR32kwvy3uROvcNTqFtMd/U4
4+/NnVGSvqF/u+aWwXAI2vli7PJtpMx83pCkv677URsF/sZ5TfnY0C5HGvDxqbiP
yf6/oZ5jtJ0aXd1LnZXLCIL5ZnhWEnPoguvhpwVFF7cG+hIb1tdfciFXlkrpblY9
pae5V2/IWbBkYnoaP86wN5p6M7P32j5szna5EGaH+HGclkIh7WGnomdSoHLCfj2J
4tOh1kTJXV0Qb+OQKyN0RphQYLH8Bus4FkBHeeaUnsyagnTPuOlElguxfW2gVLjc
98plh8FWu1z6bnAnF3EZxiJfL0RnXaDFwdXUa8icBgdOeKHcMgLANSZJyt3x8glC
CpogktEp3HNmypxS4XMW3M6obbT8TIWrUWG6Rs5wrSdeZ3GsqZgX0l17ccB9TI7j
4WrRKTXDAZbgm/GHrTbMdVoEK3rLuTI9V7/kqwUrc1PbHKxGWoDq32SOM5vq76T5
wNq51ZX2M8VjmJyiuakSNUByw/4kRjdf8+OCE0Vsv9YrRUchH1ivJBzNYJr03AIH
UDxS5pmjhkQtUpd9DRZX3Vn81ImS0+eoSMXjWBIM5aueyUus5C1S+R6vSj4FZPWA
rNz20YB7GO3tlxIlRmw3quSqKppceeEEtwffmfNsq9hE68x/Kg7OGhD44mwEo8qy
35iZknirnb3T5tkWoyerENMemJUqq1tAQmoqpGpGtRBFySo2WuH9q7p7W695lW9h
osI0y81HYQVbbdbVWYQcdoIef1pQSuEGfJw5KnrWHWoYxw3qE0+KN6mr5hQA7xy2
TgztswG6nGF4FMng0ClVz/7MfW1TeG5HV/NXljXk9E6CTNB77EMfULwtz7zDYvZh
at6ztLb0f81WdZ9h7veSlb7u6j1st3XlPA8+OvjRdjSl84B8+SWHG92/yKl47qBE
FTUz/VUieEa7TYfCukBfDTZY5B374Tj+PWXYPODu0tvSEDSs6+CxjmX4dIA/nLxE
qOgv98E8ZeyCMoZvajmmfCFbtEUS53/O/bgpKU8wV0NnhdwYJ5ftv1q9u74OYFNF
mdwrQBAtQ3xdNJU30juSFhLzWyrEXbNGsKIEaoX5nAFtd6wobYuSUpaD8vW8TX/j
XyfPRFUkbq3sk8EbpumKkwdfOodZotNcmcDMQcAURCt8XPieRxgbzEMtzbh+Wc4w
XLKvLcyuIvBOZlE3bvhC0frKUxhLfiW5YA15Ep09YE/KDofqRLinhZ4hpmL0AtAP
Lp2Se81JlxK/2/Dj9ynVA3S/gGzotdLVpvnhNxXu7/nqODG8tqfjAH6q1dDokqv3
Vrx+0bx0v3nPjA/5rF9J4JBOORS13j6tEg57UH20BEWrujTcJ9ZPd3lV/N0mo36Z
fBuzFKxoriIOAxLdMslpBkRx6ugX7L66sp6OX6xOpyPQwzGS0ADdr+USO0A13T4R
0eX2WUOLsyFqnOSwj/IYurGw369XnHe24Cm1kR2876alLMrNeLyjhvHJk8FWXIyW
8taIzBDhsCK3V7FDlwku2g78RNayoKJ4sPXp57Th2gZo195GhEXymzGuVCGEMgKu
RbBfvnMG3HkufE+41B08vYtXjaQom5ozlm7dpuxaoi5uUwogMYNpEHmo3azyw2fz
8gYhvY/jLRohaIX6jx0SnCPTi6+uyD46+nYCW3WJfD76Gh8npKr6j5KYAvcvBsla
vrYVFwH4uDf9tYQmYXJasNmWww1+YKiPp9o0abBqVJ9hL1lUaFXuW+NQqRGAyxRn
AUdlGUtUHeatZvLdyiBk/URK5ZGYD2wNCArwQTIHK6poI64+fGSCjqb9S8gb4E44
hYSggghGg6FvJcP/5KB66oPG5hF2uGBQgXajnXf0/diadocqava89go4FfrMML2a
jwFDxJGMYfKNvBT8Bf2K6vdaBMx9KzzhjZNgibZ11izHIF3YrihzmowowIAegyul
+FjeAqBbUildHbXWDZpWhbL8AK0R6YM/6MoNxiFzRLA5xbfU6LN0S1dzQTThFtdX
qs89T2JO+2jfPgpDqM4V017nqMQFdXdT3uc/NOOlUa3xcwGmJojGIjzoDxf2h0HV
bnae4mdzPRTByoYOrTA0Ou8xNMFBfWhuJ954XjisvKpYCg+xzXshoe1/0s4vIstE
85M6akVXV0uHWqnrWzr4tye0f9cSihGXf1Z+z/UIkzXo4UL7IqQrkZ8rxPzQV/0O
6HsoxC570IQ9gBD1nvvf2fKxU3PrbNgv79CMiAwqupyqhMA21Cpj8TP9jna5pAE6
tanhyeEDKoy5CoXHf6behsOffmXHHr4/ByYUvZAjWCUpzJXsIQ/40l73rp1LtEqW
wQjOlBcWYczAITlwXK2+jlhp3ruk2STNr60J5Vq/ADUuXFTiGntUeYxtPj3SxSp3
TDuN21sx+5LI7mHW+P5HYs5FCTgi3jn+BehkQDI9FrNe8yVofo9cmxZQJh+I/2d3
WTWBRJQwB6gMY4x5efynwVNLtB/P3VbGwu/1mu4V8kaEsCB93/ruLTlyrSrTyGGb
kk6miXtFVq2MkJCoWInF+0mERw1pi1vUWQw5N/NNa8J6rvxtYLiEDVr29xl1Awfm
obZP0ChxeX+Tnk1s4bQzq2t9kE7NKwlugcbs5LuXd9gauvLAJFEqx5NL4w9bV5zU
xhVZh8zTU/EPI9pAmp/pyXIivBeTPZQkHKd6tFu8iucifRgSkRUP1tRuFVJIfxaB
OZ9oKA5qS+DJnrc1jRZy6IpPtbnzlCSbYYRrEW+J/kNNItjVoZU8gE0T58kbCyRl
w3to4D9SPUE8GIYXAPJ2HjkUwTtwLEWCZwyErbByNacVSJ2oBBfrSu7b9z1HpyFY
ZZowyYh3giTot+jcXb9BB628HkacEGJhQbVJtH2Zpwg7puYNYI0llS7rxkLDnz79
3FYTtLLbv1j9O2ujMUy/4xWNN8TL0rpCATjJD5R/CMRa2Vl8LHZ6y5TnS28bzlzH
ZJjNMXEVxhk1N95/SSK659qfalGiV0Lsaq4Qx4aShhr24g5Z1SONTTfj5HJgHMXH
U0d++F7yM2BHvkH0SlL9ZuKpqcC4R453qVZZGKq3KA3AGgfLT0LSy2B4zZzmOHZT
hxg3B5WdRHrR7kJJ1H7ComiyA6sZ8pZe9iVBwr3ir3XrM7n2HCdmTIaGZNAzVHyT
gHbw6O1wOdpI/3sLYs0GzZr0iFVrpnOe5G2xrrItkaGrosPNZUA+AKhHG9FAbn2o
jVaqMIdCysxjYj1ZJJ/FHh+Ev1/SpyT0uO4LEKKOwkzfNxzcMp7aaLnTgaapvhRM
zGuaX4/OuzB3p+gQN3lrK3EfmGrY8TGiQjK46FyN9rPR2YTFId7YccQbK8t0CX9N
efHI30cagoCi+zzmlLYV0qWWMK6kPNhz0kT9AK17vcn24DbztjtGb1JaI58kukLN
LX5FpRfglmHtoGxwq7T/AsuTYHYPBGOo4NlbVJ3AvBhSfBo0ESIcKDETirTZ37bE
2wvacplYpfE0EmRAmoZYJaFC43c717/V4+1qbaMf1ZQAZLzNeOnwa9ElJrexTo4R
0YZ6sSL436rUziTii0DkgQSFwfm6WettjEld/qxhBcW9UP+M5gCvmOCne6rKEGH9
cOVjelRaxE4/g8tQEy/mE/m+e4b5LTt8DO5vWdy6IFg2KXHzvbAHHRhlU+X2daIH
Tj0L0gNxmpTNLaMUaQoZqGfB1E3MSac/3E8oAjtdh4HIsq3B5yVy5HGygFighos1
eMua1YfsypDKMAzEEAOuiM+0xLMzZHhimsPXsLPOYbP0zUbyJtgLkxcSJyp+MF6f
aL4uoNbl59y/acIsM69nMjBuILytM+P0ZYNuF6v4cl09GTDyJOTRtgzJr/DtWfme
1BLTnRk/oVohqr88NP5WkEQ6C5x+7eX0zOa4jZKuRZPsaMkTEj1cSq0qZGNtyeXa
lZgYr5VruLUTiJCoHMrEuNzNIPSVPVAXVwiDHZL1M5FSpd21GH8B6xnJXYvXFc+e
zs6KimqMDY7wSt70fBi2QmVzL7z/XdbqrpTxNU9ATHgYY0IY6Bm09EP6LTtwIwNg
7hTr+GaMAE3z0EOAsLgxpwCPmbjoqcpKkpjM2oQaRhtExbo8M5J5HJC9hzAMdzlf
QoD3ZHWs3ASnhUs2Ql9f5JnWRPTSsgQX4Ol5YEz36H/SzVhkysYooBz4gt9HPjjB
J1cXolBTqOcoJvOmx0recoE0947Gvj01tzk7ukgf36dADiUVeZBJmNvFGr6u7lN0
u4kb8NyMA6AS4mNKjeK1z26da+/XT/oWP7ewUcpUZJ/dwHEmXE16POwkviLxbyU1
1LcrhfBCAPKnhpacdoOwgzoCKFuT8Vo9g3pbfxDDtoAUWmshDYwocFrCXnDdwNsP
G7DNGSXwr2aaw9ymtSR/uAL1axuYvVMgTWdyvdvw9y9Qp5k1p1WrTtxyT0TaAiIX
iLu2eRBTdp6NmMR9oKZ4GZ5Wwr6yAo5SGQ+AYaHkeVGXtwFLnKjCc3y+UkpbUKCh
BVGN4S+a7UeBT9DT7tkK678HfkcI7EAc5VWbEJmmZzMqkUUbdk2gA649hFMnw1Gx
sVojRaKOlvQH/i/ZWDfrZ6H7+r3IajFblgh9CZg7sZX0Syv4/rTIONc1k9Lk8QTB
o9f6YHe78TovrwgcmDoVb6/JehoLPIbc5pTGxi4qZv4qUvpDJPZwt8J6sDthwYLJ
Va6v/y43IZaL6Xpl8gt5ftTgW7sNsS/qbyP3uDWHza1AyqVw8U/QtsCEy2ZeHgw/
hOmmsZKuO2wewpLmC6FAAgQPzNQRN3CMJbOidRCotvT2Qt/RGdIdV9kclbBmfO+u
rljz/kDA4lOoI/7OWAgzZGva0TAA1SnVb1TfwQjVqQxxGDfctPqA7Ltc6YcYOP/v
33M9jRxvIQnWTjy1Jwd95a0L/STQeI0va4SQ1yrGMgpGzwOj+4Ich4+A/3tJ+hjx
mup8zOxQGdMFLkaaigNCaTnbvhuZcUSgRBhqqA1E5WZWBIpAgrC+c7v84xO/BssU
wsOFrhu53qkP7tnJin0NOSH7iH1N7C2odtI7/4Ti54qOZqYr1fEHOm4lt4JRgAyM
Qms8dy7E30HJOjJ6/z1pRG6XmnCBg3sbhkj7o6CbE0AZpJNSR9NOAEu6586fPhjK
AkDHf5e9qVpzJjYzM/q5lxwAaqIZd/C8pgPB2hxp/Kzf/23pwGLRFTuyBI/lx6GP
+fA0+nRn4ZJglMFM2dwAhFMfEUfOgKBfE9q3fH6vo9zXBAhBJBgZbvg4PyGFSBZj
HMJEHcExfmzcfWgGGd5EVKu8KNUjsSNExGJ49QwuRIQQWOcAgk/gGex0Skhv1GMM
JGUsbZKHZzmDJf0gxOMRMaOauMLnZZG+F9HftqTEFYN5LdBsJJHokAU2+elJ0cWC
xLkQqbNZcRGetu8MamScHGks6Gxmnkl8PRbqF+IE+FCEECV1kz3fzXM61rWDIgOM
HQPqdNVBxgditMOu33o7JYuGvEzQc/zg4qBNMUDkIJMvcNDY/CMtTOtIvm5tY63v
d2OEAGxRy28Dynup3/HXwbeXWpo+9Galzmp5SM98c2LFtpRuYdUVLvHcYQaBkD0p
f3m42oD1yTLg/jtcS8OYstd4YVNRnOJDi2NXvps7ElFgnIeI18+AONH5DY5vDkRw
N5xoPAS3i19JFK5kHDWdkNFQ2y0fl+am4Yrrl9R5WOwiQjryIhoSvy0wVcdtQ6Hz
rKtLDcY6iYDU37UZumARbvr2d4pxtReyO0JDLO2RJRShSqI0mBBGqwNoEtNTjZ5/
HPpVoolXtkBo4e7lkjD6mTkX1CvEKBTr/q8ck56QJ8xEPUzs5wOdFyItujlhte7v
ft+VPSKhq92EpFO4YergQ9bXAeXm820aGABhm2cOhpL0ov0GPcMnWpO+YHhnNn8t
w4kg6hMeuJsUskBcIDFwr8a2EbIXUp/nFC8Lyf9WkI+37r1atp3TASXWkrlAfVgI
QLNrbsZoBnkvMZ9iKw3GO3ELOeqJGI5HF/Hg0aNJrY/wLuII7lozKU892ng/bMpD
UruhtjWCGI0FB9bU6ghZFYfBeAOpPpBvO7aroy1wFgaBzftjzBb/Xt3P2iSOicxS
E8s3/dnb/aXVLbwtDP8zd9mddagcWG+wz7IqGAv65BnYx+jPTn71R6SQyo+T6uNn
mMZOaSA/um5n54CLHPtKzp9L/QTxOmU6eKFDcimHAGBzpAO9ihOsPzDxyJh6mZ1l
IHFQO+7MJqCO6WQq6BGEq5bzBEIRtHlKi4/96iKkzNUHmahR7ql7E8nA7rbhyITF
A5Aza6yqd4SqIqzAe+JaR3CNNhy+7V0PPLWOtt19zYtKLYLss+DKTMaP21Lm4SOK
thLHQZ4o506xMeINVDssBa+SA/WrE8K3L1WhlzNOEX5BoU/Umvp91nF5u6ZCRBcv
C8EEg3AKOp1MnX10yrdC//rdwrCTCPuaah7O1EG558gyrI6iWS5dyk06dxA9YUxr
nvfEWSy4Gjye9yaocFQexHTjcSQzq3qoxiaf4YQe6IBlgJyHNhB4B7N362xX4I+a
pwVwMknJylJmoAZVYnRK3x7x8iLMAupWCM0LaihkfTx4gpo6EE33kixzfywfCq9q
0qfz1W3UVq8J3sfBTpAoMMl5dNNWe1+kW7i6rIcFBjRkRivpyNlKZvX0e400VJu3
tnMSvAnGbpmODnx0QgTqWe0IUk1lCksA8GS2OqMHfmxPKvIwEneYqeqYDMKtRWO4
u4OQgFRomcKinaqLQstm87SshCT6s6UM+fmBDoXi4v+cPVo3MMGZuEac9aN7Rs+X
+mmQ9RPc/34MBmtD+wW/76VRf3mDkv1dXzWqBy00OmiO66xoJf18UVhob511+zJ1
ZQ9l9KGV3o/PHM3OECDkbYnY43BIasYER7Vw6FgOONUeILRSSf5ZXF3a4vBpXr0J
millR16M/t9IQJ/V2a8qZNqq2KxYhPhOBliCdaN9vKMR2SmuokJMVYjayxjgyZA5
499zkW5wL56k0/m2If9veqndmxh8Wl4terzDBTofi8vg1OvlcCErX8N5vonRkj/s
RNJxfyJ84nvDJ+u51BTTtabaB04SYf6Qgtrqa2L1jJHYGQiRX1mYtoU1gT992VwT
h1hUXB1QRItNzKRRTmugHEWaQb6pZDuOyJ2FgUm1cOjxuJSDYYpJqX9pN9bXAScc
Gow7MGI+26FdNHKMvYa3AFw/J7BnLx0enfLDkWGHaWHeD9qUcT4cTRAAFM1CNFVS
U4lI57JhRr7+GlDJkrx9seRTEuiyLJ3wqKmgeLWWk2fJlK+evL8hZCVhzauGXkxo
gRVpTKaAwRsqLK3t6V939M37SHQPqQPIu7EOft30rgQgHYaVNeZqVXMpl3L6/3mE
ktGQc58QrGELm2qy9cVv5XK1OF8OqRGVVOX+oh4L5WG29xjqzIKAzWD4a4dWsKH5
Hl1alOmId4ZH/HkCsgY7P0qhF0ZSCI9NpmekGAU3MuREGtctOSBJ2kk6bt4uh4v2
Wfw71gG7RBeoN1SJ9hBZadW5zMXFCAFa6utMO/TSFlHLFT3lM+5tWbicTs7Olq/9
1wApY4hdxmSfRxwUM5rnYQVlIXVVFQSDNQxyRc0Ex8bDvVdB/2bxgZzq4MSTftj9
S/lpREXat54juRviR1X3bL8rF/Feev/Z2HtnnJ/RP8SDIs8bZuHB2A9DijA9qijM
3ZykpftNpndh4CIWb/1+9z4Yxtp/AXuM0vR4u/ElPYg7ipAG98NVFswX247paXFO
y2PehdX1NN4lmptId3Q0t6VPocZ9XecNgrOBOiUnp8icSW8kaL3UTHPqUuKJYZFC
OmlW35QcUUDu/3O73JQg6eolKSvBnUT3W1Uk5strBkC+NQ9U4G4DG6ZRAyvkY/hD
ghVJMwDMDsHrGF3xUjo2cNKh4rRZXgJxdl+Ti8Du1gLjHVIschmuNYKK/FbP/3BI
XXdXcSvMfUw+q9dbQdDUyQUSRwW155nmYRETtwxb56a0gmKL55tKTgovCDYjyYV4
oYs50hYDYLXV8vVdC3sJQ8CIERWWPl6REcNUH+qDCqafEzeKLSylIL6J+L8EFmP2
9mRcVkblPA68c0IMaOA24anDSFLqcTZdjWSNLmXNDOhHLlypV6v7r16BZ0BAx9qZ
gRB/dXRiF6vgaN2U9U8KZ7bCNjUmXKVanHOG8RBzg/D/u+P9gvRnFwAjDwz7mWOY
kwDkoG82HRolAtx8bI0yPYK5xbpaAgedwXImXuoZ654l5cWSyxCaArLhFumnoZUv
UCrkLlxq9kX2GGAAywi6RMcOpAJ08/egXiByPSPJIz6dpda/xuFNjgVDLI0Zib58
ImtqP6TP+bUB53ozV3I0q4DDBeCqZYn7FoRzjvqHNRrSVSbJU4ZhLcGfGjK/5Ihl
b6/tCxInc9TvtdOdq+R5tnZM0S0MLnddoxyf4omHrXQipcWgut9PB9ayUaZmwIHm
m3SzkPW2mF4LhqAfG38wWQf6uh1HAkx+nWtRFPs9LeF5s3gpAUjHGCIHRgIq1pbf
mNfsDKmberol/H8VDFQwKZCuQdpsPe+CZ230WOvuKKc5xC/POUydgbtJZPdblZoF
+qG/fdR9jBJtpue4GC0R667rRMwzGcpFCCQd1uN6csjewh2pimcBuDFeOeOFIjfd
RcykQwg/jY8Mr+yRQC6q3XqRGVPtrNAgafN4yqYtfoWvbtHtzx5efehdsCixNxv5
5mccnfU6Ik8gx+cFqRvO9jg7wzZdmOMfu7J6OEQN3ziQhngcc8irchR1SYTl7EQM
mAXUzqCmqN1LSrSpVI0izJkwUjdANtoqbzpOWpsQ1cGjzh5JPT3raFgwmKNysDs2
Tm2p28CLNrscSlSao/ekmRcRnxWGGXuVbI7xpVzOqcXTSJmUoXM7HZc2jO7wjD1/
ILushSxTEYkMjf8ixvgOzwXJRb4jIOa2eagszvDwAdlXJrelQYIhS60AzdGVXHZk
0P6Z++wrfyXJzKRPVSQ7y8m0y3NeV3kcZg2evmM5G7dHYz/nYQ0cGVDtxvZ9CUHE
+XW65XnirfRyHon3Vug8oMzj/Q+R6Yy5U01M8Vjcx4YeOsJc85K8N/f6jzh00qEg
/8AHcWS1FU2Wu2ceWpbYfTj453vhp/EZO262tK6sVuftr6LM0Q2rVD4CRErXa0jB
FVErlseMpUUNFsRzTjPXHWiJdXHNYAqtbldzcRx4X0M100m6QtNxvZSN+cvDaSs7
QtGaraPMi0f8ADVJGvXq9E0CbpSIwCCRqtReyWpWWw4Mb1sI0lVGnb2s2BJi98In
D0WfVlPIEDAayyziyDpPAOH2/e96laAucbKLzXCNCk547qBv454nUk9IqUTYMm00
oDIbJsbQgn9vSQvc4R3Im7JaZw3xcvwNq6pu9kfqHISkYMWOwaKgvCIcgKFcEtUr
KTzD4gkooCsdZ0MIJ1JOh7N3Kwen2YLBCPERJT5Ce7ciJ0MRy3X57xskDrL3RmJM
0s54Xf7jYVnOSqZJudSumrm8MWGwbEXME0XN4zBBZ/2ZosGPwwzeU0L6OCxWkCZg
5opzBkbFgLIE7vKrx7iKYZYNhONQnska6eccYke7zdYo6JQJUrH1ebZ9KPKrIl2D
ZLfiwf5hEdqlrzYmkFPe/dT8rxODA89t6WBc5iOIsbRm/ZN1tMEA1i5IwvZuFAkP
VSZ+kVRNIsfvWxRpXg4CYoSg8sP7FvCy2b9omsmAh6SvFwugiADSe2SQt8TVvgLj
pWYNtpIef4A3D7ZASa76qGReb2YkVsWNxGAztGT3i2vIzv3rEBZDC1s6VRPLDl/r
tbCSR35F4v0SQAdFo4UesRylQKXHvI7MO/Flzf/J+1G3rnBy13njN3lcB3nypuqT
TbZLwlJJZqTCeXNX1VeoKIFTyKB9deA4q1RLI+ZTDOJq9S43p/PSHdfST4fMcpA6
kTGflcbqJJvDlhafAe1Jhhx9YKK7KRCMlHqaiwbl4x2VIAAPgOOu0O/eBMUaTIf0
t9wuBduiOJkthTtuN1LoyRYfCYHLpS0hY7v08zOvWky2YmOHSFVi9O7VPjayZO6l
88U/DrVm40fqavE/nGzY3eZTUC+ecKmSHzwq5WSljYffwEcUJ4c8RbInbDjDW2kK
ILbsXhou1BUUwII5ERZt/QwP60Q2adFIl9CnZCj/baVXpGRaV3mvswGQ8ByCbNFF
FAsK/dBqHXX+zM2RAzAMifiqe8tFN97K/++POksHBqoGfnN4xLUBZMSoORul44/0
0IDOOfT79TquCdINeOS4IgTitmXi2MDttihC9OUvPpBthaWWjC5sR949SDFSJzgh
EOfrCqr4WTOsfOLxWmuSWZRVhTOq7DJkc7WBAYWX0gwYgRr8AjZZfh/GCcRTrMR9
8hMiWF/nTKkdo7NFu7dXM6Bdn+KofCf3MVj9s6gnQgaalThCDH7FYDIvsaIjQbbA
IccRwRF8Cp7Ellqk26nUxP3zCbxanua5cpB5lZ8mdGqgQmGyvEb1MXpSKBCOOgy7
CKMnHiqaTfAh68KvYk5L+VpsWhTwZuQ1xLKzK+fxMkeoBXhGx3ls/3ei0UZ8vl9U
39en9B6WoPjCxQCPP4EQ/ZyAXhG1oSdB99Uh4pwxyO3t7bhGY19YzeqSe3gM0T2v
LUOzQWXB191vQSRRz3+swNnn52yelOfJSGp0iXagyM0+H5MLrvdckB+Kqe4GPSlU
vz5lTZyjvPUPj+6f2Zl7ijLin82fLt5pqE6ULItLd32Xsn4TtTGj9dD/oxQGbuy6
8tYemAsMnPeLH9NeS6q9ALDmxT/PsZjKnQPWwxH54oIY3rIa0hDsGgcMWeAFsekP
gCDNs6Jsrddyz8vuNUKv1Xaci5PW2i4zEogrT0AHHjyrzsOKFWn27L4OZXOki5F2
eRg8czdxJc0YGd4eo6j1Y2+hPkahuEPTUeiuxnLi0NMhTahNOokWTb5IzuM9hXDi
fWCSb1+mte28KtxiPPYi/zTnQFlAVFyBDcu+LYUMQ6+SIM1Ekqf8a+7qhPk2bIyT
qvdAgPXSzNUDKfNJvBjMkmQeEfR8e+Yu3uT+OSwwThm+wuGF1eK964DIPXTbC6T4
XC3e7qHiP8AAECovPV99R7gwvlwHhV4V+ljPlnf78V4EfI/ZwmFmsKTAPWMIcIwr
DFggLkZi8mBiuUQkReWl8QXWPtsAz+Z53BbCFnMfNnY9atb6BNowtxow+a2DNGRK
rKRIy98mWDS+6OP3cKuRDXTb/oG3ItO1X9drz4i5YIXPz0QAGIjRUhnQ/Hwsn7mD
OUVXdh3zL6520ezUpO4y7tinQNym+kROkl6vKfMl/Z1+MInLMR964hibTgU0xUHi
q9EImVfsV5bPJDJpd0I4RG5vIfg/jVPm+EllpdWnIPkb+0CVJh44fff39qBiHDOJ
yADk3ANBEsq2dglBxxEfzk0/vCuOh/lDGsslWqO3TXp8D8LfGPd92YxFcwcU03S1
it6tIIynfErx1506vdqQRKDHLKRUzgG6rAruYH5k7CSo+320LVBL75v1yMB1IwHP
1pjGQabPRivqvn/ccJPcXgZNy+89cy72aQsky0X+rT7anPyGXbIhmkIymbINa0nW
8WzKLHqwbwETWeK2WgDdQA+VKNIjG2wLFDIcqzf+gYnoDo4zIXIsRp/pkVyEey9e
RtMjLyU8Qc7nAZft4KZOBpcyItt8T5JdS95El1blz0yVGJ6MjtUEqxnFumU+VZN1
fwButJhLrsQNDaH92KUzsUR/6o8jdRpxzb5Ati2y8Jy/GqyjEgAN9oT+iLYARqul
octvOfhN0TarIkEfDYVpwvtSr20662S0MFyScO6bKx6XnJxTMOYmeNe/8YNNT5za
+Rp+XvdHSxoAOJNPJDTanahXdUyiu62/nvoEZTwFA2yMMdtbR6fSVHoeen/H60b7
xNsX6WlRPnil/a4g0Xz+cnsgzuvu7A0KpnHRqF37xkQlsC5Bk/u8dLKSzN74GN65
V79AjZPeymTfIg4WmIEFnlc8DHwmMOG+o5HeekY2g/GGgGxWR8z8q0DBWuXG79bD
4M870vimJZSqmMIfI5ydPQ/eY6U4RuiWqjdST53i5loAwjfIvsAJRDvoXeGi2JFE
K3LBffmJWWg2h6/iMId47Ea5MZgU+yeaYgzBBUinq6ANs1cERgJgsVxtKXTiVCrd
3xHGf44MCF6cY/jZU2x//zkh2M4nW/X/qa6iGqaUA16dW8EpHFRokgwwxfQOXbd2
XH51l+BRZJov7/82zv2DM5VjFCpbJCR6Qc/iz48WBaxQRgXYZIRoqG+WvHWXvX1x
fhOejXjs2xJLBs+GWBoPO0pT5X7rK5rJ8zgn8rCHf7kevRaiDgGIeGMsuVe0eX0+
Nutg+7CpGY+mHQ+IsXV7oBc+WdqpIVQiwKBqFx16exEZZOP3mZX8n35o6rk7wPhy
r9fQDWAEExQf9gyZgDL87QOr45jWwQHfFBrqhM0O6RaoWjyiKkdztDD84AqOzxjD
VS+3eYmTN8rDDyc0ko0B6Wd3HDTVg2jBnciP05TBq9EcL96ZDR5l5TghmHBcZtHB
HL7pssEKb/Q3p6OJSAcVtKtauJcZV6+CON5YwgaybwcUWY+kaYAQpwbcetA1fD1/
3OM39kDd3PYdLhDMd1qYrE1+AKwYlqg2IwnthTYzBG86Sj8yucSMvW59/luWTN+A
fCWdYrXVC7DayhADPvkP0+drUcjb21eRnFmRQflnaFOmUXu6aqWNkfAnvFXX7kfE
/1W/hINDfKIvt0BkWa7zzHZ+SpIoGWNSziYWGDiTu63PjAPNn7wG7ERPx40SRvdx
7OwVILQFzgTp6HDO3XGGmih7KMdHf8Jm6fLoxpXcNRxUIB5wusM9LK83+EKjVIdr
1GCTSQuTnjNuCzTVDjUzX/i6vL5Iu38jkgAwSTxevuxGpHOC6Yh9V8HcSgaHzxEt
R7e5r0lybq6zV6ZwSJPMW92g1763DKnXEmnBCyOz5vsy6qG0iuO9CKMw1FC5eayx
ZbrIKoG+jKOs5sNpFE2TY2ktjxoO37heYbSWHklvp/F/fIvS7MaPsBUE6mGZr0ku
WaR69pluKeV4JvVQUR4At7Ra8AWqepomq/wE1+3kTpWZOI/hgT7//x8qbkdRUyiA
S68YBZevPsnc1g89nBdR04tud2z2gzOtpo2ZU2Bt0h+bCKJBXtpSCB29rMXDNiEa
sF65eNcgQ/7TITFFj/b2OGWoOk9thZkXD7eKwAcZJzRnt+nOcNHVqD4y7CT2Jej5
XjKLS8vWb1j4cAHgDQWp2NE7GveeQi8OYDSuYrYSx6uKtE39vGyzowV6nGZAZAms
VrCyEXJDxqiMEf6432jLUKGXSuFekDwpOScgMoR/SJCTfWe7UMpUPwHjrpI/qeMw
2/L1QuU0m7U2KE+A8Hgfs3XCRHz0Gx4TpYNFUQmaUACVM6r0d9O4deNFeG++Z69y
GOH8/vFZAxUyisAdbQR60V2HthBNHRe+0OJfZR+9S8m2XRHry5NZLA8bYJGfwmUz
niDuKK21Fufu6KdDfIeV0rDYWzWwRJtylMlR3FMeuiyxEpbLD8dQG0UA5UPvSsaZ
xpc+TyoHZ9idnm7ax4UUdKlx+erVSJQldv4KLi7mKeYaSnZlMMqKUP56DOgn9bx5
AvPcuI7dPxRLmgHup0EBHbd4X0aEpT/WVXY/bUsaUDicXzEl7wB3gsJUbN7HXKd0
3yP//rJP8rezluEBzDCNFLERiW7FpJxLU9z5fBKShiQUWj6esFEAS2mvNDwJ0Gvq
K8PujcBkfTNbe41CzIdiyJiKWlWrr1ft54W/uAVikBrAemkPwVNtczJgHdOsTmjm
okCzyTnOO67sQ/YH+XrSu0G7KkXksvZOTkMCk//BPA7VzaNOriI0mHsnXwk6HoVF
KEGJ3O+9JuWHfh7eXOrs05VXQeeSbRBfQR6/DqXIIgKhdNLJryAmPhw2cZZjcBDQ
a3kXmpf8b6sTYKi2B4WCHsDk5dWGhKljgwCVY1vof3UYM7aNnmKsreTzqKSF7Pap
SoTSy+ZLYiMUvfLxcVyYTSBQpx6qo/clBYWfATVi6mbkYMYKgmcO15yxcHZhvx2C
XENkd4s6HaeKzM+CXfl7JI8IjVYvSBxVcmnGXHXVlrnweaTA5XVsbkbVaiB0eXPy
a46yMBdB015vS27ux98eYd3hXWOoOTbcxVmXQnqzQZ3yk1ywlBe81DrZsAnHeROe
vN/5l+5ya0r1kwRVtpyM8DCute2xxF4j2pA2TyYIW548fE9ZMU3mOApifbhgqTpl
+/Knd2WHd2aUX8woPlam6MjPn9Suc/Pyog+gB4nY3LoQ9IRoPkKtwvdPUF9yTtm2
cCqN0P+5gyqEDAw9GmQ4bZMwYi7cIi4Ci1fURhU4YagecjvVecpBbbSFK0tAzIGR
6nafUPXBPeTUXyUzMg6DmmiYwkJnkTMIJbkHM/voEsQ+5szwhkOcIAM27gYWkt3E
7RinMDGhX+XbXjfpXKFtHH2sjGDKjDhO42jhczq+NvWdVwcRL+MhJqG1QYSsjxZJ
Z23EqFmLKMXdj4GuUQLzxYr8NtWLIdd5bPqEadvqjbyJtBiXYPGpyXx5dUREwoZe
l9fMrbtELRBdhylPv1/1e3Xp4F71hIefxN+LRo5ZLie87L1rk9RTZ7n780zveWq6
G7a08Y7ojYjVrnLf5bAj9kFK1LVXHULKTeAxLspT72UtmAYWhmDk3/q9K3FtSxFE
6loTPU6Aje67JjrjSNeJp3iK3t9cZ8EnRw7pG9pfLKmx8CvMzIag7nGQgbjSTZPq
tG5/tt62iKGgbQW3qWPD0Dy8yZKaVUQAOZ3mKm7OMjUtFfZfAkDmgj9/JtUTgg3O
wfroM4rsg9ALp1s7CVIglVkoVwt2yD3eV9BD8v8937+NDsIgTobfpIgmEcTXv7hc
AQdhwDGKFwYP0tlwQhxCNUIkcFdw5KNiFTBowpBPY0sDGezBLdF89YAuPBQWsmJb
4mwyiQvcsiZW6HmvbMjmo3KHM4mno471nwUvLRux1X/CVj73xT+MmfrLI3ZGj8yC
MbVWqRp4w4yM2FcH/nSohsyc51P3CqSMPH8QYQNooaFDDatI8z48aq5/P1z0+dCv
kPSte6EP0/unlKxAeZM/Qd1g1PUDSsCtTA30s95CfuDwMjromNQithNhZkLVcofK
ycN7ENRKH5LW44Wf/RL1kuvrzyBNL8uvYA2QW2+vyAfq0puGXOJr/FZpWjyNLOAy
g+drwOGNGlEx+RFiVnXThtU84F5Vo+UjAs1MHg3czgIhFaUu/inOAfvf7vC0+qD+
GG4cH3Dc4/2NNLQe84YuIKYphh53A3jXOfa0vsBcg/BAsYYYunZ7QXi4big4qRvS
`protect END_PROTECTED
