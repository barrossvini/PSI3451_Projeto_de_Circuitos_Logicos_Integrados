`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iTs2cHL9hHy8dcT8crDpHdaeyQvez+Ix5wxTBzMVv84BkT6LGKuxuzxpWr+eeBt+
OJH49D1vQ63FUR4smhVNSnblrcabVGr3bs0qdkClF5TxR2RoZEGjqQqNEwMPQJYg
xqdLqhSMxD6fQV5YxR+Ew0faTUHJhM2MVhsaHlRlWKE9aRSWgwgiCI1JF/9u5bv1
6cTUZAEQrC8hbosrMNmIgHTrGwIKoSOuzCBbEp7keWe9IS8AWvhVWVx7RCkSFLmu
Y1ZWPUIKGnhcx/l9bU0FGZM6y4foR18fDrN4C04lB/6DF/wXVH/UZxMd6SX3Oezi
12AqYcVQ3Tz6UOMTsdcdscOXBJlZ4msw4o7g3MObW9hz4PiOuA4Jl5am22b648Tk
Wz+KLnr2IHWztQA8EA1g0kDY+Om+wfndDDl2wMj/FYVX8iTvK6vt5yAGoNyVHXcv
j8S28Ex8na0D/9uzvCW8Hyjbs//mgjhuCSMJ8zb5yfsUOg42CcuNsEJG4dTRB5ia
UvAJPuWcVDVKrCnDYlFpfS6NhBYK8aDRCR4YxiEzd2bf/0MX2iPBOLezyMejy0Ab
SI6J4XvA+je9BrSQJCcf8iYGr7bfIEV2H3K3HFHHhAC7bUzeG+LdzZ3VqeIPlvtW
dQV1Wx2hkZHUfT/SE4jXTnfYT3MHzGEA6S2f+I2PsehvWTLL8/N80zYtDj+zYem3
P3h0ghuuyRtnT3voQAhzfL2EKSDZgEjFDXy6t7lmYVLiImIiJDdXHtDHi8WYTuXP
+na7m8laUQuF1A2v4O+lcuEJnjdNe/klyGPNTUo3cnA3VMDp3qfrJaMWdisTqifz
PToquJCWUPJCT/dre/IgaA==
`protect END_PROTECTED
