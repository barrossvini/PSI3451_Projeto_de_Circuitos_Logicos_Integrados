`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NP/LxX4+8QwYXDJQQmyckiz/pKcLCbhLqH7q2Ud6DtSKQ8AtdUrj+Ps7YlWJAffS
kXUuaZ7a56a0Np0/DsZ4H/p5YfNof38BACIUcAUXvkZlR9iKRNnP8UM7ouop8ERC
E3kRfTCZXorTMO1VqTkrLKtIicw/Zv2aPAhlXCuVlfL+5XcA3pL+rImwAiACQQ+7
PzBVsChVLqYqfQzI+lwrOObGq7If9w1AkzCL2jgwQlXXOa8IEUEf2+JwUGBTiGt4
zOBEQqPwQ36fI3/ADCCs3s6KNsR9WyoxFfGr2Bl+syuVGGO80hINwQ6yasy5x3je
ro4KZxyjxaiNz8THZ9JljotSRRJRifCpubpPJHeAFLNqCxIxT1nlvU1djZPLbeZT
z1ZH7/ElztOJz6kCX9l7Fv0tSM7ccJSJnzEcIvMp5JFvdP24jdS0AkGWKBFH12Hg
vBMEdagW4IdwjqEfvVkJzjn6e9EWaFHhYma6oDZkhp7KPXU5jJ+aGPzntXdh/o4d
8u4u85TVk5fPyVaVjTwJcq9fZSSXC+txLrDkWjIVdu5dJ2F+bu7LF58omqT9lwVn
qQ6ImPcrQiAJw4r08/WzNPvS5CfBYMkAtQgtDqt13riHrbjUzTtvItp08xvqW1/h
sjPsc13ApsFvmtGuWmHnchqhTPnN9zH4C1Lo7bHIwNAhSfd/Eqfw8GCuDoCAPR+g
bUXtB8RQBltSaqfpIIHe6o6ZpoJlxLYpMgh23kaewh6a3e5owJXB1oOLBgkMjxzp
8gCwJfx3B8TFME4cFgtgyVuVhpJHLXUJ9JG6LN6VqdKHIe8kVpWuLzcvVETlRmvj
GUnjbQgEaFh+Osq/0RCOfzRb4/sduBHC2+pDxfi10JOgsxruhJ+eB0LPCfTnq21A
IlqajZUd4y/VRcfMsQphnn3NLQQI697MEMi9N6SfUe590i3C8VEQ9TdhBm8sUsiP
6Rn5jQ6yijukuq2UIFMqfNNJmplPHnMPx5+QSFcRS/3lX8uKyXUv76/Px1wXlAxl
VevQmsWizl+CEpcY7+RD2ewTpBXj+4uZ1RvnKLN6C7gCy6ntYXYeJzy3sh6tjVLm
SE01GqzRohAiGvfL8P0Tfz6wvIVijDBaY6xD5Yh1Po5ECuiMJHiMRLSCmjpKJ7Vs
O0vFD4/V37lOFdrJoQCBBennjsVd/MtYVE1GnN0ue54tnjjt2+eaRU8aIeiKyqjA
nSdqnl/s1SI+8yVi1MJdYPL/qTYxjr0evLfBpPleEJjZY0LVEO7jifxnejMmMibJ
aUlO96Dd+7PPOXyPe5ulZ78Dqwa31cGLf2Qy3VEIulBVP4akL1dkH8sRncAo5FTq
O3ho4DhnxtuL5/3X759oxYfl2epl6JwFdBbMezPnMyXbYTm/cSaP4M8QptTUqYmu
K7GIbZuKGWfjlC4DHgDVqFjIiyrOkfmEvz/NT2sbn5GkuTXUx7w48Wl2iQ0AX7wC
smXA8JJQFBBUFmqlCXJGWY3kvLdWN+iGhzpPHKARQwV+D8u8nJmDvJmw5uSfaUuM
4YJnw/sGGWIrpDUOSKstQwzg99+gNKgfZFqoD5qbY52+jEHo/u5jRayapUZj8RaS
31Uw56AGvBKZI/wljcJXMPCEvqgS/6+DOqw7e/vehcU=
`protect END_PROTECTED
