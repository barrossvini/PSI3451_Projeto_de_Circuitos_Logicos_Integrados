`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2uply+Rc7Y181NLkSK9zu06SxaEaGLXYk2aQdros6ztEDy+F9HkT/WhJG/UX+BDn
mLG5TM8hKd21syBVDZ1X4NhZIeySs4BSMaFAFri3JpYfR0c6Y65tB1Ij01a0DkCG
QoCTdPsUpTAUK2gNROR74QoJrnQOPvxZpovKgJE5Gf2ILlGdWnWB7AKVLo9f9eTc
fb8ENJ/u0kn8bDounFpzrz4A/wGSUR2MRk/KQVvZE/ed+APbpwyI2fHMXFO+KC5w
BhlofkXVR50M1tga+htU70uZcd5QbQvbGDO1zcnGNpYQgY1Iri8CCOo9GSopxSSQ
EhYiUCmicmZVcpOW6BsamQ6LNAKPHH/gxGBO2k3qcvs+V0Ej4aoCEAX17e42cKXj
ryIMDb/IRl+tphoNawDvTXH8PQwGajgvfCYJPCOlraYaryJACiGM8Luzqbz741fh
+rq3wyXq833icAyx5Jk86Yo4pml2siGyBp3xmtCNl/I3kg4JIlz6UrP6V7Ufg9ZA
U6hn1iACstXrPcDBwn/L+wIP9RUFEv0rvkOZCBpNk0pKEfzDYFeK+O4qtdby2GXq
RpneLiBtEXnZrP3OmTeg33MvlidmvL5lOH+M++d1xKu16otGHTN5wh2n36k1uCfZ
C2lvHt3VePiLW58olz8p2LkXcBBgifvlelD3tG9tCwsTUQ/Sy45hzjcf+dhCZ/Nr
OLjKbBebcypFVYPbkWmNZwZmS8ZEUi5hCi8+1vEflm1CyODJ7gdLw9rsQs9IqiJ4
1hmA0rzWa/xYhgruXmKNGaHRvxP1FIiMgBix8APdlpNgxB0TzSufhM2t4Wpf+iAR
Aktr11ttB5b0MuhOOQna+dc/e5DiBTv3R/eNibzOEzRtkzux1T6cQlQJmbCX2wC9
e7MdpL13OWowC6gsOS/ID+2Z++fYGDoTAqlmDcPnzr6UNeqeXD6JWKfOWItW/1Ce
+ofqmfx3o34DFAQJPGxfypFqAjexsqZ8g+AdPxqqEZ35Hh2hPrM7kY/pl+4hE5jR
C/3j4jCxDOAzsXeD0KRartsNiLZYPyh0N4Ffp3CAdgY4tnajuEJwP5SfcO0gAT6O
4sFdS+tXYjAAnyavXR6ZiaAYcCxvLKE2n3Z4wfgbNnyZA3odBkygN1SYa69ZAHNq
eQIbPWwd4ByIbj3bgJdmGp/Wvvu8IGVWEK47IyhV7AJjpwG73nbtlPJhAfl6hE2H
B0Trrj1+uhuEgxFXw6Ot6PL+tJ7OHsu8LnXnYU+HXwqp44UMtotz2YkRVamrWUd1
Z2r59YmCJ012Dm3VC0rwupR0QPdHG+NqKKLwT86pczstqgGRTeiOi9gz16G0fyFh
+QF1WHwgzwqJTVcTX75NCOOVpgSVJ7tvQoMmxtiJdsl/l5Cdbk/jJ+raV29aO4BD
gsX2fU8rBdbNHHpXfqVYNnrotUQsPW2mTwHSasEZJBct+o/0LEuPsIET2tmBdIB/
VpF2qbn6yAZPRfWqb3azuOU89tCZES7RP8+7aZXwtT/A5+qqTphuiSDTcUq230lM
FpAMEUf0xuVoZ7rz4ap5wdUz+pni9+VUS/w+7kWmMFSuvGJzqnomTPJmKL5Vcm3b
v4qM48xo6lkTSz9MohN+K02MAU+RXyNhmnAtj2Wqa/LQtF57MEPkRR7J/RjbM4SH
By5P2vuJPDVxuEskzaOc2eVlE9MjKmFST2mH1h4N2CDhFYzUIE1KphAWp16AFkHE
Tu4XCC0vLr0K5zkx3pDUNFYDaP7ug1Xv4q69f9dHpyRb6k0jsvyXJnSF+i6Q5Otv
mEJZ41xrvRyUFCtR5E/k7xLVoCZLGCCUvC8TN9p+ScfDAwTEW27PtXaGACrVSayQ
tjKuMr4EJimcQ9ElsZnj7JxzO+HROoFA67Ts8/BuRvvJuyH3WbV8l/C9U1CevyR0
3bD8be+t9lAQARB6yUi2ZnNiwgbbp89MNcWnhoBBBFG6Mw8sLXVNiaYcWPDtpxEO
5CP3a8/5ijWH7VjL/9F4cV9O7ixy5cfiYUkXilcr9+N/N27n72NJwjlIjYbECQWW
+wX7FCrKyGkRslPtXfx0YtuoS8RbS9UeEnhpMppHfCV2O/RbhdmMFvvUd1TYBGi1
wdC0PoMuQxbLLr6C5NuFLELyAqOhpLtjAdzPRK9+QhanLFCx/8Z2OUEWLKl8ZF7Z
9O/j9Q9zQybTXllq/3SzuwjjPT0JYNbJ1petafCsYNyZ1+hOqd3oj/T6eb7akfOy
sElH1kvnRqlnjitrw5THhSnGrpoh5kGj0HXd/e0YgjcW11eOAiBFzbZsLg7KY6rH
icJVwybBb7wJTDbxtBRIEtnJ6xRDy8NvQgLY1JKNq9jeJyvZGmllZ3BrypbkvPnV
l+dc9aj7W+N/5LaEjqTEo7uBQ4YcDiQueK3sppplbg17bMgox5u2uWVGkIPLu028
H7svA2EtzAaqZ5c6u89oGFsDwFwLh+sfPwne8+7n5Ags4rU+l1gHM5tdgqwLFJvZ
yWL5lRki0HmqJQFK+gYPPg==
`protect END_PROTECTED
