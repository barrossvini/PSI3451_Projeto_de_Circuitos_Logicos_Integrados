`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8xEwtuURH48SBuKncWvQiOVdehfir+zFt87qkmCV2n/NaYTz9mDbzUDAb6MDQbnU
ZLitYbi9TuwZ+O6+FMF5rvGhsYhJIevsS92f9XKaxKEdzsYj3qRHDeiGx/ieJyTo
2vksLmDjSy30tuoAKFEzrMQNhJ1i43yFFZO7+NIhNHaWTMj2xOejch2AbhnY1xZd
N5gBN+SD9Le6IxCE2rc7e9ypvCeV7u6AZY68y7EuKZbyZ8RSQdy+1hBTOX9nwKob
SzhLWifEz7UyMoJjqQ8HiwoglLhfPrGUbQ3Xhd1AnotQqTHB9QNBLrimxWqL/X0m
TZUMOjIeh2d0o32U7gV9TfcAZk+PlJJdmOL/qjqaSeC36tlda5kCBq0VFNVjEUdw
auqJH/hAY7C3fTVA3p4k8WwjewWaeMBmb+6xKBmah6FdT3rQH3aUNGjCB6m4XaGr
gBMQWUoaUI6vP/daQA5r/O3EaF123dqlXq+Rjab+cM2p09UT8Z5JREgOeMk8RBWW
CCt4sz0tOXu1Quc0KTpsCBFSacbNbcEuH49S7iRFqPjIHlJWzWeI1jZy5evElHMm
3OnopnTa2yf9OaWeB+wtO/Yvz1oc5TTrbE+tAcFLij1LMxLEULuI1yZQUq4gup0d
n+uDLu3y5RQzW3gcJUwveMEufzxNkwBUwDRLwApHmWsFH2VbJ7DqAIiGrJOn7j8y
dqQcULsb9fhKkXlw/jro76LmHcTck5T1L0hI0yGv6NvYD3wZNhIMQLWSwPkRLATv
Q4B1idsHGvMCMNXwH2posue6e2xXThbApCZkLzhecRAePR5eO8ZaK7MTUmPoNzl9
gqpeKzrvhyfKkqNVKV0b9DE+o2JZoQbnP7aEcNnkMqOsxTdLCWe5p9RlrUOLZUsF
ccmzJtLX61rKEm/wMO1V9Aj3FFraqnueko+6ee66hOCFIPQYdh+2IJyBQRg5Rs4M
fBmPtJNmgBU3HNJakrzfADxY+i3bw4dqwNX+zi5iqmAEHp57JW4AATtoVce34Fkt
xNMC5lL9BT+eQ3oHSLT90x0C0O90kWeUyzMjV+zTGFGo/cucBujKlb6exQ/DRx95
GWbCGWoJ5z/G5j+NgTbyba3EfemryQvSthtZ5lW5ltdnex/XTbpz0waEJPpIDtgZ
CAlM0ukBst3ge4P30Uk73mH3rTomNS2ZsFNsmWpDpuDm6nJHDAYS9YmEkWwf4tYp
Ma9LUv+e/2q+8dwep3qRwSB9XFbZ/kmCCZCdUfd3SFUOryNoSO8v8eTI+X/YBc6V
FvADVeQ0VmKGf7eoOwPJ3/zRzqV2OiimWfwqGG0Sl21CZ5heTuOaXiKH7NzqPVoh
d7jmF+BFvotHizmOMeYjtXDfZQfTHQQsQPR/ZnAFOL7vhAZ50dthoVqa2U/SjWXR
VE1/MPSrLb55IT/kZgqliLuGu8yCtW5VK1L+0bdkJU56MwLhG6uedqCOieWYpVmt
36Vyh0/5VZVFTj+SnH5Cxi+/HyNUnzqh493pbPZ3XsxPpLsIbtnm4hdUzLwJc288
8Cj8qUpBAB+IiVAcAgMvaQuFVjw2Wdvuujv+6qI7ay8=
`protect END_PROTECTED
