`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bD242fOTfSSAE2aD4sJNFEnTOAnqM+RnBj053tjly5vPWSwh8lRB4RS9HxpEdkqA
pF/Zd5E3G41uLvy3r0fB/KPQcD7dhhRNxgyfPDhIl+Y5A5xoF0an9aryMoxx1mtt
17+7mif1Mf+NRaKxS+OuGElXzEf1XzlHmNnSq8UwgRPF1PFnMH+A3565HArBKR0p
EJTnkKIox/OUsDCA/Vl6mwSdKKaBic9MgdjZ7t7pcmcChlpaTMaQxvnzJ06QNPF2
XV9bZTnFguzIBdmAPUUEix9XkLcVxz9oOEEapqE4Rn46IPvDavTTXobqybQ5pS0y
PFpUvnaHbSIlewn0YC68ErG7DZpXZUjSEIC9w9SFA4DOdiMDrGcdnAMlSCgPefON
PYarrGxBQ06g/FdFq7rvqApetXuZ9EixZVwJ1BPTEQYp8JtTHUGMLy/6SGeklK4C
fG1PR90pz8Vec+Xafm/12c2XJmw4ecyJi6JCyj31zK2Yffh5+4uAXRyCCaGTnbQT
gnq/1Z4wVL/NZWMt4U8FMe7OHXPd0XAgG5pc52PsgoMW7SKTXvBxNyMv+AZF3WHI
Y6yRVHjAWHb5wNCZMd3asShoE89HtH9qHsp4vpefmgpuLu1vVXU/Fek3Iyj1kfI8
UEw5uqdeljFl22PGoWpUR6yWWz7zjQlLexiOHeUB0J6RISROFzIY5NEVtt4/fn5c
`protect END_PROTECTED
