`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+djPSUYOh9Wo4MkaS6+3z6cGx8uW2CnTafeUiiWQ5QJHEobvtnfDY3WTp80ZeyrX
ePaQoqskmsqWvl1i6CRjcbTGRJ+V1FWjpNycVwr4SQIzpagjKrMeuw9KT++I1Ae2
worX2gchJGjHcxEK3b42nGoGoLX3TBV/SmwKjfmw0dfSVWwGCr8VikTsjhUitVSw
I5EJwJflR2FvkJn0XaL5TttxrdqlYiUoi6Q49TMXw8y+PxZU8vwns2x95g0Kyqqk
PxAxCWh9qtOmoSHVwuNeOHuKez3PQ4YIYgz9d2wPsh+mjtd/SKXpP4pCzDVkBk6H
2ldor0MzTM0eU1QhdmPb/Q7GMXIADuTLApsTgJv3xtlf8/5rqP8k4NtKWbvxTRRa
nqT5saPSeIKHUsMyPEkzn0d70asMOUQrLR8spMcUgxhan4mS+a68JnYG6lUdTsMb
NlK9q8SBsznN8ujugY4Fe6qdKtQoLxdLdgRfXdpBxwCMQzJWo30eKApDXvWGcpu6
gsinHu/02ezb82GsbBner/UtcrufdvYWnAw6l50D9qEobGOyBRJ5C8u6DBji0kfv
sHkI40uv72VPZKbYj9leHBO4cZK50eGijL6ZjNp0kEcNqZ3OdM32Nmn9zjDMkDxx
fXoA63A3GrlgNuL+juHfhLlUJU3drjfM/eMVxZtlCVRPO2y/7wT9awK1kLXnxzEj
tIvReSXb+8oTPvvEb4tFfIQyGwA8k7f4Ev3TaaNxseEdQiImjJkhscGinDI/5Cu+
jAF0diKAB4+wpc2r5yfxib94e+j69SBre/XVH2C0CnI5R2n0CkiSr7V79U+FBQG+
zUHWGAwhCtjoc0fmeowDRg==
`protect END_PROTECTED
