`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NjAH0GUPQ70Ak1Qglb1XFp19quSLQjbgmmp4WyErKK3B8UkkAazYAh98EmwpttNW
78dYi9GoKoBYvFcTxD+d/msRooitufl2vqufax/GqO8ejasKCPsJxdnX/jCRwq4q
XijMniwyIMGFmQObEIRnTs9wXEWi0QA1FjO0SU3afApJ3Zk+cd6MdMywMMobRacY
pp5rlTZkwTNJMmfEMar5oI/IZ0d04H9CbjSaQ1C7mxnDYhYaCdc1Ek/2gjiG/g0p
D5yN+I9cwB22AfZFcgwF0B6zhcWkxHyowKOekgm2rQKk43ejva8Lle7CoENDpm9y
wfn96hU0aRKkhzJcQaFvta7xoQKAxrPjc3bRYDR2EwOHF8v/gZXi8BNHfYnIotkj
PpwrfAs4LzUPX1RdOcCWBFMIy5sC/G9N59/Atr7AFiw7GBFEiYTCR5cMpzNfu86m
iVCk2jUhki9CBndETF6ZWMGub7O29iYeVLtyFKlzUZV4eshRuT93xZZ2I8Ih9ieF
58dtWtIEa+dQk+mwQ5vvbDsouxP2IzCCvNgXHdSnBukA3C23NusOIkGHgrnU5E7a
bYwfgv7oMaMgiSRv+vSZ9Z4uFeYf7pHb/YF3+qMXwEc7b49DT2ObmCZbHdRurXFr
amrZILJqnkFLTrDLDb+Gx5+L2GSQJ4T4pMKNZBmuPgKtwPqxDW3xQAvLxTXdcI0x
Cklz1PwqYCcEuGoNO05mYy14tsz9dvynd5SLskCu//veK+dbcSos1vIkF/eWT7Bl
NkJ7IGDz/clLWNZxPvYClzpj/hD/0qQIHZU0kVKrfgzeOkI4fBE4oVDeyqPIk2oh
ZnBL/CHfNgIgly5AIwj/9K8Vp6aWGvdDFHFzfbQfHBZ/13YCEXZztvGLC8GfPb53
lK+tvy0rAO+jXWKqNN1W85dXQbsvvn8UGKrANkJ2UMOrW75pX3rav12hh8bJGUm3
qxlR9btlvysQWAwUKaC4dZi4+q4jUf2d3Ik9Zm3tEvfKwUdrapdpMLI3Rwu8CtO6
iw2dn4/t5hOq/BJCZLJtXjsuBOtuewcHr8L7jpRYTUYbgJuQ9zEXVb3jaG+brE/6
5bkM/KcR/gBqgvT0+nW00MFWQTiROxnWrUWjHw5JlsXAtoCWi3WurfIqhjRyXP+v
wMiYDDN5An4gADC7yrkI8jq+tRcHmojxVwJCnjmC/VHcEi8btzF7d86MSQz+MQoE
gg7lR4qsePXyYGDjulHbnr/1ARlTNXeUWpn4zD576Erd93VDPEtHPX7p9XcvhGnB
V7bXpNtG/5PhTMeaQEd19jZWs2Hm1ucrEBfOPvtqN47tfL5WNwZ0Phc7+xNO+IND
YA8KXvHgTL7lDYV+zQ/JXSTzHj2a1oRZGdenPGsZQqUtXxEHPMzGI2S0wveg0pXD
dz+PFjF9d+HCUdv2XHeTWQ==
`protect END_PROTECTED
