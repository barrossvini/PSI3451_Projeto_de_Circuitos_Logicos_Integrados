`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qCCTDhA4vTqg04RNB847nue2i1Jr0OkjT5xhPkl8sA29MtTsahBAdId8U83mjO6S
FlLHSyXGHmnFyImosH0FnNpL1wFVrp7UOJkyFEY+NLFZR+fR/GFEbV58et4vfGeM
D809X6oabrXaYzOa0XwwtJUEPwKtHSDPH4zjMWYXrLhBasX/kLuvzmMTbIEU544l
bU+KfxqIyDBMcDjARnLn+44m+Qr4rDo1OdMqwtvxme2H1pCdtowmH9UGgJjUFbLE
k8/khPvhNuxl3xrU9sqX/AR053cCfUc8Di60lSNz5ioTeQG5a6wLomppWUHmpA0x
MbUkUc4gfB/amzXrxr7Z0LI90gljAzLAcWq7XO7sYEnsyQ7ASreqeJoPmXOrebbI
JTTFzehqn2MNfp/XgeXUqLCXs9Zupewu6Vndllykv4unJLFhBR1JzfQnTfZdBxEw
oBXXX/7CoKZd9j/XAksrD++IUUI+Pi3yW+G2//CYtQ0hXinW2OlKo6dY4M0B5bZ/
hai4wDtZDu268eGPdFR8xHscddw1BT8w6QTCEmK99wmSdKhwZcVKj0UZLFcnyo4Z
kUf3B28ZwHqIiHTC0fc5DXUUrdi6f+1pktBc14qV9m7APLWzUDntVl3FxyOG4vw9
8IgXgZqYRyLOTlqp4N1TfnFBFTDv7TAuvh8L+xzhu9+d+PHRi/2idsur8Fudqrjm
ARTOH7md6ElSyEytJTDpVMlFFPWX2MNA5xjN08rXUh6HQ7GcOeWrgVSxTkn+LOuY
LXbR9xSgLbdD9M+yoSaz10xmpFpSa6heTqaUzOeRkdPzwV3G15sTRWcgR/6S+Z9f
ktckeBiyPU1fgX9ZmED4sKoHKUcXk9s5srs7VNdy4/JIVeCTpoJ79sQ3tW5oTkIb
5/NUqiF5y27I84e9Uo+qSBz/pSYOMMisuB3a4yuKzVR4WoKu/phGvPY7EHn6VCFi
OGRwUHweO7AqNgIhRcY2A+qDEiOtp8Oqf7klA7XuUlc0b9LoanIKdtNVfrMNq7xU
eQ5LeIvJOfgYoPZVlQRkLbWccwKmnv6F6EFNxDIV0Z21xnyfFwA+4+IRSiKCoaJo
XVJD2Y18VXKGyuw+Zb/4Y0O4Ue0YLHs4u3udT+8tY8l2opbtZmCvqCys8LvfBM0L
MHO6OUZC1FCkJRhGeEOYukI6LLjf8k3TB0CdWpDwOVUsGzGUqSCizwqC9T0R1sOo
qV64WsH+rCkU5KZWffDiqyhqQrAXy8T0mSY85fRbGzsqdgMzN8ejKR0nYuiL3+0d
KI3zUJc9gxrw8lwyTmRuRBWp8O0SUzKxazEEQxlvIsLxV+K3rzK30Sf00TmscYvq
4Gu9MTLqvnTVWChUnOsGcBr13SztbMfarMKWf20cDJgAG5y0IZmguYJN7TQ+H08d
f5h44qbzrMBoJSroxhgQw+lJGfKxI+Drtajs0epTEe+O4VIW9EsQda6Nz1/H+Bnd
KQdbzjd7OE/rD+IsdhPToQglMVLuS2gaE7HYLli2FLlLaZAOCFvp/7u445t0yVtp
FYYjnj0IxuMd5MgnsDcMTgLibW8hCckg6/3BjNA9FRCDZ6r5PdfzhpWEAQrtZYVf
t8+W1/penAiMhL0G+hsAd0Xrs3ZtehK7fAo/gfY9Pa6DIyaPZ8+RZ00OesWVGmMF
aMJqJBAL5a+6wSRyetBv02hyRo6uogI3cmpJmvgxd/x8xuH3Dn4P6O6U9mL1H6Hf
WHa0Lksdey85qcilm74NpAVdMXPUZuC4yE9tmbhkt0Nb/aO/m0ESiruclFMSghwx
MT/JeIp95vdW75KY/KncR5FerPz/5OUJQHAjxcMpbF0dQTXGxBmujYJobXhQHeqI
91XMaQ9nyTRgZYo9DlKa6d5gymnlwoWBvhU7za2kSOWrJ2RaPtYBu0R5iHP5sHwW
3WQfOe1xQcS4pwDK3IpR9JlKh+QB7tmSKHP/1JbcfucPpsu1GRgDfhOtKQE+M3qP
TI07mGd59NSLd4msBS3U7jiVXi4RehdxtPuB/lnEbrDjHoqacuywIh2nW+jVU2SC
TO0JMTMjszX7RC0HA+93k38iX1muRgNqrPH8nP+RBaCG7U+h1YFWAyfRSj210mCP
byQ/Qu+7h5nm26QN63j1Uh/7M6wAOBAkAqNnKn0SNKA1RcnJcNCgGQGxhwnfo3Jr
5BXoPh84VkOFRwQ5eUTWpyUDoeK6w0eIACucC2X32WU+rviqXyEf1/rfGW/ZQv80
5B8LeQn1qXFRMiPEdWmU2FBFHSAgM4Rx6TMq6eCT1q+8Fex1Z2rjTVF07//iYLuS
50t5JQgeEtbHbmK0MTaMMWBUUjwpef/gJLyMhkYhsJaoujBms5/ciA8BKO6wLpJd
H4fOp+v4UpFskZ0jR6lheAnmwX9CwMW5/XruNI0YiTbTu5y4y5BycAeJ9MoHZSXQ
yT2VnyM72MhuXNiE/PFEYw==
`protect END_PROTECTED
