`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jAeOestp8i5tkrVTD2vyHQZCBe506VDn9Bt0K5+jbC8Re0RasDIs/HoGQsD43ext
t+t6sIiAbdkCR2P1FZJfzlUU3Z+mJFAqatW2KZT5jjjCQsH2B1HSGM/znkAGFSSR
BcNCS+mJ7gxql04OVNrxW5Kr6umTOQekfUry4L5Hasc8hDXFamqRjyG+woxVqIsc
iQdjRbxKvBlsDD7SwKdosZNIfNfWmUjpjfVgmOH4qcRBK1jmBso8Jz+VKFDlBvJT
9TEsIhhJkuTiKUpWcMR3QFRASJxNGoz9wM998hs3CN0jkow3fLgs4LSTPnRVmDwx
bbicH0xn4rci9HZTRjXOLeBdu0+2YVCtUAedrXXNvk+KoLG9uHYToB9Qkd4kzsCG
1f/o5Sr0VEGM76jgfskzgmKPbKf79YQFxxlmHVHN+iCswWfqhxX2dQbMh7di294C
C0pMPxhL6lE1gku3QQEj0n5A5idmBuwXKYSPbe6JtEfV89jPqgYAc4cp+cCGs2Pf
tmF5ttukkKyiRFKX4cPRAuo7VZOZ40eM10AaawxQ+4wNtFai1Qn7o8Wvgv4jd+J9
6IRO4Jd8xHJmR7QTh55gYciRm1xkgxN/igr+mzC1CpGEfzySRLSKMSvZwhn0FYvB
fga7lgrsr3y6KMCMvkY5gYEjiO71eN1jS3gPRRLcBhTKsAUBu2kEdGbO9vAKmNOu
3TE4fRPq7iJzGqK45+7Fg8iqW/28dV3nA4ITExTdC2r9I0ubmt7cAModFO9nUpLL
gHRGmEi3YIDsUKRlM5uCOtuzYgiFEj6tJRT8rbbmPN3bYkDiILSos8/xvxAUG1bj
uk58TnIjpQR5WhNuEJgLwK853BZAwFOaaRBUy9cFEFVa5PBusEqlJUP4s9ArFe5E
ULW9H4rOH4ZUbbRJx7rtZgAg1IIlwDy1wDUPSs1txBsU0Ouj7LO5vjlTmnOicwYD
DOph/uwqqXuvOOfcOZxw3siK1L/2pYaZZzsonlGVlOczWY8Lp202aqtvFt81x1F1
8qYJoOiWZahf7kBR36fJbxVL282uJrt9ZxQ7Md0cRZPUpiCACbpMqgchWZ5MxnEv
Kj+E1EQc6IFHETb2ye9ZPAVmHzlBFfJpXfi+ZxGB3AT3MbA/hd7E4OXBido9bMtj
+cuhasnXkQIiRwjKdaGbans3+N/7OMnJULtgYgbvbhkljcE08aLBnvcpdMgNvaJM
V5cTiBf2BbiWbpXSnqQ98hApVYkz7aBHJ+O1v7JAzgqeEgoVm4BeF1kgKzdYPn27
nSGsHz7hfqM+u6hHjauffLzBSv/WYpA4+pR3zYrmIBH+D7TvK7lX3f/o+q1Vck1O
HG09mz0afSKTX0og1q/8NrCuNMBplQBErhUWnRpKGOyxXkJ1iyZpuEC3UCPqjxQu
aoF7YQUfnZpPeLkDmam8m9qEvPq/veEix8KBMJoVKCG/hME28urTc3E0oKy0pZbV
4ZXmLQCAKX919XXfttz66qkM32eu/Ml4Kylcg5FTBhJrVDMlTx12mqf3rPi9+8RO
7/HT3Y4fNUqNPFJx21LFPqSyh2dROOn66Olq7i8DLAMsFMcx3N41x+xClZOv0/o1
NOkoLt7m0F38B3jvbcGZUbet2j4TizpiI6oWyxFx0Gq2WlfdLoPVQjBKtRIdi2gQ
lvpqWteL/XCKjVrxD0cScW+hvKKTLUyQ6lJPpR1c2tziBfrjdM07UTPQSoXrnEUE
KaQ7ky8ahw5LuYzFHS7erA==
`protect END_PROTECTED
