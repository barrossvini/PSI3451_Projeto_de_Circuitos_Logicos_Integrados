`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jHkpucIVtdgXvXeG4cxWIMwpGJRnrYFJgMC4/jAQrgB0sA7kGwtT5wOT5aMRdva0
uHte5j5tqSx6nYPtOKYhlEMhqh4M1vF06pOkc7kvMXBaurxf43ISeQA9Ns9gAYRF
UDKfhIppS721/+jT+L8MFhzJYDDB9DOawjWw6/Z9HFjg2xUnCZquHmV1opgfgFYU
O24N1rT43kGxOhlwEWsOhc2n7Q99nlkfEZwoX2kVSZUR8P1tjssCWx8/ZhhsSZh9
cG71+bkqiNEDZMwWmrlTKveHtJm3cDo4olO8JRIGEEnya5T8Jw1LGxd4uBuO7R8D
07kCqRDUm0TTg9IXbQy+j7pNESWc8/D0UvbNbnzer0Z5fe+u/+FTOC1oMQjXUVWb
dPhciFD5qqwXl5Gee9ZI4Ok58m+sLu+zg3340AsNLea3Cg7BV+yuSi/WFC3UGc3U
9z6sEbXihmRlj8NT+6xGR2RG/Z+U3CEs37ipWJnEYlTOJ6O9iLk3KXUxD1E9/GIu
VOkQrQsUlvF4U19oRMLud7oxLWaJAJm+4YXdC8ye+s5a2sHcQDEsLXEQ8jsKCX+D
kKENHhUJL0302Ax+VvXc8NQCAmVQbYx0+oMJwMqLSp7Sj2ZEfN44pM1C4Y+znZny
CWyHmVzjnuyqlg7d7FiudbPamRLSg64501f0AL3zxxQu+jBtW1MOeXkw7urIraGO
qsbhw+q+KyTYFT/Tiac8eKsRQfXvK3KionDbmUNYELLx9BBBuqA4I3II7HsAYhwb
zL8txEJX9weT8bX4f4Tc6ncRnQGBIbDI6IBA3f4STAuA7fUCekwRBr3tsuVcPkbn
X/GiiPo+7T0Ub4pjPSwVZWV+MslBWhO5u535arzrKDcEmAQtCnwR52LBdcleHCy/
maIfnNt0Ae6IEyzywb4itEUDu1xsE1JCX3Ei1WxgEi9kterXejaJHIIKHHjW5RfG
4CXJn+cQc0h8ZjbDwQ5O+RvJTM/17fl51Nk0s7sLJcnYWUNVZC/LpHaC4LfjrwRC
/ViS/doFED3sqfxyw8LP08hjAMHF6MEM/OWLNW3eIIWajIsqM2Mhfx9oPLMaHDXz
j+O3DfBAj/Pz7J33HDOmNB/EtNpfY/43O1+7IxMxj9REJshXQDKFtTJZg9vl/Pdu
/pSzrrPwjNm8gAUQ5POYqQ8YKs8c0pbMCEbc6621C3qdf5m00oUhzNzJU/oGBDdJ
wzz8HTKShgQKRggppNwRQvGLt3EXngOYJJGHBnDGj2JtHLJdKdssy9uBfC+lO+cG
wKnbLkh+xQ6baCLPxPHybrQ9R0JEBF1sXMGknpgDK3U6ulVrHk3i5Jo5uYAoeyTP
BuczWZMya7Xt7E4HfVEwUinZkDOzyqWoUEwqOODnTU8HGnjQf5DisPJ5FAFocE2b
L59TPmGDkw0nX20JGE0eY/r41llr9/o/Z8FUeK5nqPK4kzHq3Gjgr8D0vRMQR2+M
lDvub7l7bG4JE/6Bslklf+XNUjHGN7SZ7FQ4X6W/WTluR6ZONfTMtDL4mBEiJOrI
9XmyeMmKtk40nbstoPt9NzqCWQ4vb9KqtD+7hbvPyJMPiw3WYZeB9RUW4+SIjrxG
4UPQ6qD/k5hUbmnqG/UCdEyWT0bs+6Qij5+OjD3IljEnyj/KAn01/X0o6e6p5MXs
HHO3xN+3X+AClGZpSUWZSfVYmW3lFxzIfMvUJpa96jbxcqSScRxo/s2P/0kGtJNQ
lGJxSyU7eBp7gqJwrbaQRk8dPtd6LVI4zz2WJqF7kjKUg1yBSgc/vEUYlwPQvD90
I72a6rYrpXIM8uapzJ/JtxtVin2qBxTL6OWnWr4L7ZgF4IgLNwfWhjg0AYmWjzLa
R/PHpp78Y4vvN2ZiWxQHSc5XmU6GjFe9eoAnsn6G9yithnwuCzXnzyIg8AjYzJDw
bOxxddMJmynngHgMyTTNhHQZEzC4bcr/ceYiOfQgpEZCGJP1zzxGNdiKG0K+Ildu
TF3J6PSIybaPc56dXr/6due9rA7pFSoq3gOsyXEPqFvVHy3G0YWKi0XqdJA0yaLs
rCJvnnHTPZOrzr3yUYySRTG4dcPgnTPz1eb96g3L2hwhCg626b3yn68OhJmBB31N
R+jwn7Qn1KCgimyAojLDJbuijf/NzWPOV6vSSIfwKFxkDYGhw+havbNGPe5NqZKN
BlZV590Gqy7ZMG8Dwx0qnDwwflEErlv/wIXwkc0GljpWd3luesnfXMQuJiLSBOsg
Hhwz5LGZ0N4XrWBwgykR7UOeFGSfYwRcc1iCFMLTVbGovgvr679+pDe6C7ucEAQX
+SF849Mefa1L80ogNGOWSIl7FErnxNJYIQAGh2cD/Ai1FB8FmrkHyM8tVRvonOpQ
cpRQrgQmb3eNuHpq51tIn2nG3xP06ufyWCEETKnvkj3oHngSBVV5Jwoq1tZMxHUm
r9WrOEKCxvh1+UkG5M3MVWKwV0P8magulPBQH4GaaUwPEsLRIp35m/Os53ZuF1+e
74ZJANvFZAerntDVQRNkm+4Vu/mrutlZTD3Jt4Bw/Y67nEd8QGZN7xnUS83s1lj2
dvEdsDbUOJhLqnbrkwec1m102LXDi6krzyrqHmsIMfZcDP7Tww0kcQAqYaA6nlHz
o+dcX6coDJBWIJLze5FO8MjAJW4lsCJqC/M3cAauNg9ExtsC80nEdavqwRywT7YM
UvtLN+Hl3kL+LYZ2OBPmFW4blNBqr96Lg/JsUwoe0zfWTfKaMtr7DTAnEAMI5fX0
5i4skcc/hUYvWYmXmjQuRDSOiQpheoVvy3g+ET0XHt3ZdVE/Cbazec96Z6TXEtvy
FwuFdz79LI6qL5PdPFzRmfzVzSQU14GNN8/duiHA9WCyy9Al/P/V9seFGbQxYYBm
YnH0WAHfqUbSpgbmkBANrWzfrNkeEBRcFevVSFNGSVW+MLgZ2mQZioOhuzt+Cxam
lhkNzeLWgVAa0XCQdPzikyfJ6Puq5tiMAuqTXnY+Xu5Vw3wY5w785vdIBu0T45kj
Iq9RJ+4h8q5yKVv9S0SR5YvYQvo9uVZcm7vUv3E0DcPBwHbNW/oim3aXEWVBFDlL
d6qX2Ik/P/lJjKiTFFn5rhVyPF1/+g9p2ty/SU7zC0T/HoFlJFgqcctYLQ/50QNe
3hZqvZhs7KWTe/CS+35VGgLizSqY4TC8O6bV+YRGVM7pXw9sU6toDzZLWdaVFZPM
Y7/hM2tzSfurkrxDcKwnG7eAC9IPb/e0gGyWea8VKJnqFjz795/DTIGWdUpgDLxV
8XFzNZYBMTInLv0DWbMuATH6ldy+bwTr7XkyHNbiCa500ztM7T0WbV2dLV0qb27M
xqy0CjZFZsChCDiBXP/FEgcYKGJ9OBjKY58SKQQmAleGzQ4q51PBaDdOqtOdZejr
KXIuguSXruiMGziUtED//att4av6aHsTri1MlcFsQXmT+zBF5R6TCnEnznUXITYA
MV4xD1JKRADROYZRPeewJoirbZShWnpqEE9aUw4V4de3ijDPhlrS4qXQ7Re92zyJ
b1EGAn26YQoz2CUsa+KW8w88Ggeli10gaEoACSf3rWWNYfiftVMUFDKAU+adYH7W
6HdyFmZgFpbznDnnsLZxe3X3RuhhxNYXVZ5cBpElL/CE0OZ1H6Di37MToDD+Wk8L
TnzkK4Zzhz1NqrqFoveu5jgR2Bt33G4xnrZgom59YaEmmFw5oFjPBpLpQq4pE11f
uS83XOuVi42pdQ1GoH33do0H8vEgi/VC1nfPVZdAQpvB+ROytHQdkFWdjh5328M+
UzrMt+ydFXn/qb7WHk7wyR7kW556pwmv7K/CAasXkV+12zD9civya8DSpmmvKL3K
7FDSj0vnyv981LzRpF3KzmOo1QJEHd3hy10K7HjE36xF24T+n8adYSOg90Af7cv6
jcGbz0MTQ97F5K9DM8OgPA9j6Ny4o/yatqieV/tjiiO7xAnA34gL9Togn0MAVmIZ
Sa+ITBV0xIOFF/zaiOacade3gRyem7o4Fiw7SucKvHBiIfzoF4jRyMDGyzeKF1pU
N265DYCAcJf+Mgv1dvM7KsKZ8bhQrHttGBArMEzUuOx1Aph09QfzeBFPf9pRZNKZ
q6szvubbx8z1wTI7YDGLKrfTof7mVXygS6XTlxCHHeXR0FTWpAwJEXTJpuAFztLP
9XBnk5RWteFPQF8nZm5XK2+szJOm9QzQHkEaVvVj3n4RmxaCi1QMAURBktYCjpnM
tCr+9TAum5Lpw8ejBpEta68zCTdWQ0jZLfuGfMMPnWWDVBUuvhD6fP4q/zO5+aBy
4x78juZMkkiQSnx/Z7zUlYOvt2D0riWrcnmv1OgVt2Z6hrnyF7DFEhTAhIqnaSN3
nJ51OglOmmVbasywK8f5O5CufAzRm7/TV358cQQjMyWer6H9hpScvVx6ZCN4K3NU
EEzGqcxxhx3ipfL+Xy2LOnuR7ixszPu+jxNRSnORBJNFoD2rmPVsZWAvyGc7Z9EA
JkpywMC6H1BLd8e7WMSVK9R7wR3LWw84jBoclgvYgvbHA76wiy2D/K4CHwvihrRu
PtOxDS7bBALI1eqFaRBgSS2KmGDxwWJeqq9QGkjGUKNae1rh+jNklo03xAg/mrd9
6VZfsHKM1s3F72/No04VZtjFQR9B5bCG8sbAcrQonIZD+OqoCuvs1CI+olT1yYAg
joutTvzt6UwC3k6yUPo5cjTnxv8wti9Wvxcaj+GT/WHOOD+UVJnRFGNWXfqCYl+O
6FdYWxqo7s7eThIPVXrt1LT5HGpmn/1m6tfn6LCq0wkSwFWBmIVtyrjeVKPxtJX8
XyKokPeIcjzqWSO+SIT0U5d3KROCk2akJP7jHb4T2osuUF83M8WR4PfZanRRwvnt
QffQiZ31b/oGc4A8BcsoIt8ze//3FkIweM65stk89pmMzRLBML1BlMyt1bjM3WE1
y/SFPBkajsa6ErZrUNBse9yxNUMKUnUYBBL/3e/2OB4Q9/6dy9rZK20mTjdmlLls
EXE13zDpxf/xLsZwGpaD+Sh72hzMK0y/I3j6pZe2cZw3rAhEa24KbxDaidjfKFCW
CwvS8g4XnmQ0dLiEguVK3ZwELHUp3yDXflb4pVRdFElvrAuVjWGRLLXqYbevzMSg
HvzuwxXQTVZSH03n3VnXmYMuW0JI6xIYY05Mb+gEKW8Es9rQlZy5bC+1HqpZWuys
pmUVDL7BIm31b6tPUmOExj+XpRuOGpLIFtBIoXZfdnrZwK2jfqfWjNwNxkHoRCtq
PuGspRRL/g/lQySB3qXC45qg7KNcPZTmWpxaQv8YOI7Mj0SZXlX6LGyvTRmZK7H2
aSvjxtbUPv5cTIGE89veHg4iY64/cb1pNyO2STiqWf0vjySHjXcVPGMPKmPLyoZS
FQ0iylDLgBm8y4lNISJWxHCOu0wiB+xc7GwUB0V7QTwvnBS5K6mEZfn3BMtFfMPy
NkVr17wrQDS3L3sfVxCjtq5UDGZPzAtGrmYN8d3y0NcjkuDz88hvsZzrk2nB95+l
KF033GsQIKH/DWNwE85y2V5Gar/ztjsUPZr5rVIZkUfNr+odZP1OpLeo9Yc67UZC
jHtcYIS6cjSAH1okicIM6hrT53nKGTJwd0TV5RKNp19fHkrzykKxGwgJb5gzmlZt
UpvQZ8fWNBnN29WGQZHaJEa2iJYae8VEVhXyHquh7I1l+h7VvsImtSoI7AliPb5o
PGDMIX4RBxUjcqme3361Hr++Bg2tXLYSXq41IXHLkDNBpo/FWhfB7iIyEa6OjjKe
ouHN7fkNEvsRahYV3hCZYztbengcWlX6V5SRFS8Fdyf036AUezdhiHW1yqPPwZ75
eAo13j+QZToGb6S9VNIbGA6ETvw17rTlMwIHwTNO9ga5nHsEE9pUP9Ka2PnammmS
c9eUpzGmmOeEaklRvU2oWsWNqbTxl6eEWRije0QRbocfxl4+NWUEwb8/8z/Az/2D
9ZLawAWrdy65IWfz1+hiFD7hOU08wH2kwbDB34rA11NoZSBLs3rB9ZluohoHXtKe
xsqeMrjNnq4fvE4Z1FVoYoz9riL4As9sVzAR3rZaU3rHzDxS1LyeMS0UMQuPdRpn
BQoyrwr1ZTlKyscWJ2Yh64oxGKwlv2hmkW3zqP4Ji5kNbkMtI6NK1Krc4iTXldTc
V2hy9jnNkTC8E2/TQPrQlMo8hxX+PHQH3kbXl0crKd6eYAmrO64I67CQiUDgrfho
rd/YO8juZUqRjkh6lcgu5OrMssmyhYh5OwTDk/XMGDt1iu7rzcBYpDANBPxnePv0
dPkDrXKExH5paQbYZukZ5s4uJ3FJo265a1OI2WhGebZt5f7MInJeuIqWm80ZS0er
0sf4rFBfo6KVNbCjcKtUi5ys/dchPFdmQ2RNUI9MeEZKCRG/Ib8UJ8EZ825jYmSy
p2LAaIzmXOjw8lPZppTvmJTpE2AHwcvU6qgR20e9BVWbmQ8WCWrJhoKQdxGPfxQR
VG/UNTE2HoMCO9zZfNQTHmmLb8xfxRMdx4XPXfxTuIsgUOiYRkpMLEhBdlzuz9jK
bmsR5g1/jPlnvcyToVqBdvPA062Ag0GBkWRczlhik7vzyWBcfnneV32a3av+ZLfs
N7si4enWyk+GGj0WNiKdHulpbbIdMsR+SzGcjg8R8NPH4h5gJwHOyWVbikxXbUZf
Ko/dkclNmJW7fFbg1asbNCNFukJDawDGLjZjEtD4t56n21u0tVhv35lqSIhsQgbJ
bCCLrQraO/FQZIpfERKY1shbVZ6kFyIyfUI6152vQXlo9myzGZdBQoXMgVzwPrHf
bGjMk8Fcr7+lLg1ugby6DiOMHBUKGSx/vN1IvphcO5IxrA+pCTubxYYrjdVBQwj9
xbhVFGky4nOMP/Xa2CNphcXVhFQxFoUwJHA8/JbnzqOKmz6zMoM/6NUge1nNh8An
spz7cPvalNmehMgrJEsZycnU0nnu46hoNzbcez0pstXlBRmWVW/6/A3qvu3OxlV3
GeE+pNTRXfPFrA1ruBtFSebF930R/PVc6wIRkSeci4s7Mv/kkOGcQg4l7zDrjm/X
R8LLg9aj2SEOYnU63jD04eMKhGqMKH7G2rN74D30MFG0uTzlqR6g6vbXVcCqQ3c2
YK/JCgo1NgQflAdho3xp6Xh2Qs+XVt1k/EJPZVJkOi8pdP4WkjFQcHLXPVuw5SDg
zhQ1BJw1oLOc7+sWt20oTwokw2M2JP/ttqUQ2hLqtnZRnIRX1jRGPBwFiDX0WHne
bT/AlHEMShh+24OGGRHeUP1XtEUBZUu0+mbSRSA25sciZqv93TsIEsWCmax7Gkc6
V0ANJa39H81Xd9aQSc9TbYwYIvCcbJZ0FJPLPrrK7JV3uWQlqeGSmqpN4KAn4khy
Jt07t5d6/13WZBgvPw0BnbhyM2+EVPqXm+4bRJbOyRa0s8v5zluyfaIL7dtb2xA1
E0aE8+SKpOI0+hW46tfR11N8a+220/sgvbS2vWs5K1yw0Etydl0mmx7UOLQAGoZS
i4AwzY4Lq+XO+qhnrO9dg53qRbdbnLgbdTCSdNHByza+O4Q3vWMReYUYcuQQT9WD
ySlHbiOKkyMGmms8F+5/WyrXNVryGuE5GkUEwJ9WQilUhxLjU1yvz0ipht5TtPZ8
cQ2qIF5uJ+gcC/kh1VkFGIcWyQDvzQei/z39y1ZGpdfX2Dx3lsRUKXSXbxiFexws
2sqjyWHDYa372HSzAtCvg1kcXPB57LkwpcbVPYmUvXG2RGngXy+Xx+gQTJeA5IiW
U6inYpTTVtge7hTI2LdmpCNYQQgD1xu2XQLvly5NvQdG12F3EmPIPULhAs8T/eOG
anoGUuTXFXxPx1vR6wJrIssZG02oV7EipUBusF5Una2bTVyZHBiQ4Q8oAxVx20R6
7Y/kIjir0M6HHPMUtFCBSMf+p+CtBtOHd2Hah7RFNlRM/l9Br/Asj1iAzn0DEBrW
rk0BJy13qSFe4gMFoeeGWEn+9g+cRx0r3vRRsv96CAwmSQqGrRW2PHB0O0HjENiG
GVtqEClCfPPMGdIiHaG0GGUBmyXBQNrXYM75POoZMPSjoLv/jnkdDHla1KKEiY7X
VGAFXJ3zHxp81bX67yHFxdb53s4djLeYC/gCAoya8qPz/3pt1YL13jDdRTVfNM/L
5MYyKmph5Yeri42FRkBtkE3QUss6JA++V0VjFwpNbdOo7ewc4CmCDYHVzIDOvZWQ
mogirTT6w391SjH09/oKRE0Pgh+B9Yu16VlTS2qFzEnBKLuHUbQjaoxL4JFu7kOQ
YRI9YH8t5rySy1qLeCHFV+VBxJB8iOTZaCDwu53HJA2H0FbOmSmzTwfoB04iJI/I
ZX8IG+GCV+jzzhUT7nV3FR7R2tmaGjXmSCEUvgPG4toBe9yQtckWDgBrISPJp2+V
s6CtTWl4++fdL5PnRr7V3knafMg6fr5UMN6ammLQSSIvsynhQiEA7ZCIYh2zbicM
IhHJh3q2R4RGXZ0V42lIS6LzI2N3wjjimdY7E8+dQWn7vBa71QyvyYwYe7IyHbz7
WgXauv938zyka51oG5dg9U0tEw0rxHcT9+tks1e0+jYVzVYgLkk6vnVsN7zcGrhU
5+uJVUN+AQlPPLcogG3AfsVcNScn4CKswnvRaguELwx3OG5zLXpeCIvVmSDCzLY5
X386JZQkkQD55RjtsstIYKT7zVi86AdTiBApGl8RjTmzsTrzeckhhfZ0x0rTAVHl
QPDC6GidaLq1TyFHnetHYU4sbPbASAePidjmpTs9VAB9qYL0cPOCUcMnbhq+HzHe
7eEkpzLeOyaGP2bzcbJWsZKzMs5ujfELko/X7o4YSF/8VLSyc6zAwKnOYPLBsZld
eTJhZgQ/otrn2CDQhHS6LxTv+70/Zb5EodksAfGn60vKrO3vmZmQJVCpD0/+yJlA
8KbdeF+S5jFOKaCwRGTh1u+60a7g7k2jvZ55YVGsz+qVj3kxkYNFzOSjJXP/BjkB
A8UWzpVRDnXitTHaq9fdnq6JZJ1yRTCNX7FnU7852Mhq/sqxYN3hg27jRT1WSb3c
emqGUEQZitYPH/ZKEzGAfJ9h+ORTzzDPu1lQ4HVHVVvxZF9jw5jMmVJzENVAIn7E
9rB5IfbgWUN1zv7yQKagTcwdGpt/RnuhmROebmAT1Lt14pEbiVWnU7SkE2/UU7vT
I2Sk/HGlmgsm2VQW7n5d7UhZRPAWXYQUFRpA+z5+LGb523/m7csBWTKuB9LGSASd
bYnXUalDe3IXF/Yo6Ki/0dp3CInxJ8Qf+Pjci7UVXdd1nRR5y6YlDKAN+F1eGxks
JJeKBl1bJ0WRlGg3z6VwfHxzKj2mO7CxZeTUEI+WDkHIGfQ4tFUvVHNBLWRQjOxA
Y6koH4WmXJ274AKoAeocBF3d1ujqD22t0ta5ef2g0BjVebs1vlCjjbRubQSYFVHG
/PAmtm+W8iDaww2gD1X/HWPVTmF+Aeh3UyBP2g14OGa03uBfA2eA5JYhdUdYyAbk
LN/ZZdtRqkaZxi7YVPteTTShwuyDU7EIHRgxK4V3zv5Atr2W2qD8STRVi18zrtj5
97/rBozdpXZ2HKB2/WlLIOThEQ8WQiYy34OlxQEXkixlyJ8uCg2ToUN4umTmcsJk
O0z8RRIznS+4DNriH3yB0aO/OilwHKtRg54UESU/5ehlO2AXBkq5QPGKOffbLCnq
jXxPcIqeUDDHyGVKwVu4NRHULSw1zm9VIeF9i4358uBoh/CrP77IP5K7nr14TTjJ
FofeFi4hex4QEPtD1soO7o6TLBVRO+OlxPrX6JE7yGvBAqwwVS892z5sOML6B/6Z
Di+9IUezPDYu8RT5ZnaLZIorjKeKNt3Zee+rEABxm65X9kef2IKvKvmtOauihZSS
BMGisBUoozFPFouufCafw9iazy9LjYtWmTNZWr54Nv7KXOuMNqZQ49OIQv4Aqq8b
y2BUPPTb/bGLYcIttArMdPWBW/2BDfZXLIk3F0LddsldlDfMaj+Jc76nfB0ZpiRA
3UEeQceQqoy8Xgl0JuvQWBkJsxw9xnKQFVXaV2rXP+oP7HTbsGaM6sXpgVxGXeM2
HKY8d01qfsKqnGtuKXjg41GbnEjyydevPi5NHfBI12Snzjcmz5x/gFnCbnfqYpom
8uHw9briqLezFsgpPhx6Yc0x9Ch4yu7AnKiUlNwftrcYddnzR8K6fTuQnbVyWqsa
ys/wrW6tMoGD441j0SceSA980CUdh02nB2MJIyTZ5d1DlY8iDTXA4aQ/D5ny1lnj
Gw//2mgv3+PTgtr0KYq8nAcbu/XEm8VpsofBDVfDdiqum81s5AQcMCi58lvkc9c/
T4sEhZ4BQJkqpsxM8MfDPu9kQGbeebCyiEu2GxymXDUrxpE+eSUBytScAdSvpU4u
Y21JSBiF/+6dMF3dQwZVHrARGptsSTF+LWGa6wyrYUXRj+AZpLK/hR9FVfNjIrGs
0Kb8XUB8LXThCB0/9d8VvzkTK9FGFlfKmGv6mY7iPTkK8hwdKyZpmviu1zV+BzCK
cibDqFjgdw4X3KtVxHMqo3NirWB0jXYsrhwiR9pq1qai0k0L0FgHTYPDrQYTX4pt
GvpPSsHfxs/lmSqww+pPdFd4vQ2QS7+nmducR9PXZRFStQ40Ns0Jug0VS2Ri1arY
0/SWwPm8PX37jzVEjCwlI68BvRFXEPzMFvF+UNhKwjDvvEPv/OB4Ru9mTRadI4p8
ZdQ1YmykEn7R0oWmyyTifqbNiD/nqM4zEKAUFijrca+4DkzoAHHKy+6XT3uvAvuQ
alg8OTdnUIQP11SjTwKWTPZWIhHnaEdKbB1S2dFx5tJukXuQ9UPh9hZ4KdHBAN0H
fzdC2i2OEiKh/qFkN6jX4zo9juB2DDgIlGgiPQheHU/tcWPhGK551beqY1iV9tFf
cGtXJIVyvnaJuBkFRsGOx2o4vXugyrcq9O1nUI1N29x8GCjxGGQwd3UV2HaT2Q+j
D+VsH7m87joJGtkszgMlYJ5NsH5mWgxJYSY2Q6q5n3O4SUzdftbqqx8vA5gZDlil
FoxzwQHs7paix1uysGv42p8vSbT1CFwWq+sMiNUGKdzlA8cOBQ1OwjJY3aM0KAA1
3qKDvf48O+wGu4BkBKL/Ag5NTbjGlznQaswQcOvROKOx6+Faj7BO7gMdCMZmnZ4S
QN15UGl/ykwCHDXAw3pjBhtFo6L3A7dBvRqoli++VurdnsDPD8F7LCJ50XGpiDjb
swYFJs71uDou9GUAOhPKXo1O4LVlsSuCLaPtSosi0ed/Ocst4YdlAn+3XKIMUyn5
u4Y3WPFFf6QsUuJZeU/iwYhN7CXfAXfT2wdQsMSHN/a15k2m37nzCi0v1NNfXdzD
g86jv+TPcPvMP+5v6rQ5Tp29VXTVYtQBqDcAiJHn3GKfR3F3SnqrdorBlFb1OHPK
AxF11YBR2ZfNRKbvrCMSa6E6qMYpZpMBTsk5WSFWUx88eYfyeQh8hMHXZRqseGuc
0ybE6NSVkdBcPPSB8Onvjj+tN3NEQkoQSiUV58c0krxTXkLLaCk28TMbEmGZC+Q3
/3HmDr7c1pJRseJ4QFXXmbol6ExJfiPUsl9kiSrQd/imYyrCDsvn5sdYhNHOWId5
y8JpyKeshYIWhEltxRG5jC4kuJaRGkRHcOt6icrT+Vt+xopPK8sBrR2ESR01WxYY
ebdfTzuYz9s7/sr6qWeLfhBLkmH5YSBQSlOKwQ1sij5ozAecRycAsuNRHdxr88f4
NRFSrVnDdkC7pAqr8XPRFqFYOft47fveZQ3wVy9xVDqY2ceYx8dJd+Tz5J5XqXKn
Qvj71zz2Xxf0Dc6smzY7PIUe+j8OHAyamAxUlUEi1cUjD+eAWJ9KEmwb5xKUVejG
kCTDPfLUaOQO8iR1MXJZiOHRREhtJsNmkleaqEfEdp/eaHW4wKsAcE0sExvwm7E1
vGcg2VmKEqSDRJq3mZoyFW1XFQHmcCle8k1E4dSEf+5wLboJPzEASoOsLq9seE4R
JgaR7CzTjLHvlsC/BCNsCYQ7NWpLKmyv24vMw9BXPWCHJUE+DibWG0tGzcK2JP67
K1qaM8LIq4N0t7G0p5jubzdac7hc6lMWcuLhNMe0RtrFrP7RXtJ6e0GgLuHSKSyy
p6S91owY2KkhvKnY9pGoRyrGLa0Jx2nAux6QR6sOP2KwVNcV0jOdEbohfBjbnbyf
Nz0HARNyPYrA/bn7f13UGrMG5KtsUuaBkh7eILYw3UjZB4Ff4MDQbwNO9rtcP9PU
Sj4rKx4M2b5ItofdxykhlRtn2WwVJXnzKe3cLOd7AxRmpXFexTzptsfmjDQvkCAe
Tb5/7J/XddkrN/VqM3CIyypkCzZ0Mvygfu3/l1vGJw7ebxuaxLpTd+oJhfW1dGAi
29NYlBV6UalZh225hsHTZ+2N7sQIzr0+8GaegTJccJC5Rt2ktdT8onIbZQE7la7y
egIt24RnILPmVFZU2V+0vVoFBbBpGXnJfd34EmrylvPGO8UYcMrSVQ9znGUvRxEj
ISMZru7NCvC2yk6NMyhC0HVVF4KgJaqdK6kAGvL+IRjYD5S6JzGhZE2u899Lr7AX
atjkABgpJ99vP/s6pzxgZxudNUx3xYmUmnD7Wk+BcIC00YeeZE54yRwrtTiWxNk7
2bzAMTiHBi/5XzwuYDD04gNz3q24DbtLR3IOeEUEMDg7Mfrer2Z8qikRZ6CsiD7z
2lq03JJnyEqYYK8LLsOAIPlggM+puXTbtjvJBvtlvcDxSiw3omqfoqiMwD90i/kg
6lkjDbVd6uoYKvlbtbRVOl50wCPCk7Hf6ziMqZhXwa+h1lgCwQ0bmfgEdvnl7ltN
xbkyncXsk+sSLmcI9kllBFhJ0E0j8dgbVwd5zemUByJMlcrPeROuWQi7Cq11apf0
5Lrn4YzVaEaE9K1CXnLa3XAoc5Fx7YIAxA6BihCvSjmLxpjsps2fr/fAnqr2e63t
0VYTkrmPpwGfxlabHYMDXqkg3aS5Fxeu2+m5C20hTTxFeizx44Usb3snGpr1RtVH
zGvlvcifunqFoWy88fE/xKa+dJ1ya2mba5653CEy+3vTshDfHM8kZwaIURDkNbAX
6x73voqW7Pv9tpf0vFdAUocNUJnGCun/puVoDKuHD1miZsXHisKCnqHfeAfcHov4
suwBQOyM4ZD8uuFDUNl9xaMZ9N8bTXACo7rqAF3rpjjqhXykQF8VfyK3cSKcUiCi
asSnfjYxrOkoBFVS/ag7srpTh64DDnhqFYkq4kNjgL/dL7eCevdn5cMXibDfHZ3q
aGdAMHiOsbFpit0Qnax5PSpGPwGFP4JV0oc9tb8GUgLbpkEm4BMOypLmDyxXZ3UN
tXTYdT90QcYHibziOXo7D3N+du35B3hPDkfEU6XfTBhkKoq5XAB/D0GcLyq0Y4yC
Qk9hNMnWp5GVv7W4/tSjdd2ADRZ7j0ebI9YCfF5MIM6+skkOUNKvhf2zCm/uiixZ
llp0d3TVgm3OS00l6G5o+NHnQDRxk0+pAMl7uReq984u3PcvXMmKsPkBjPmuJMpO
bXCAzbPX+kaRwCjZtj2IlK2RgaESCIQRXVdvNV+8dN+x0qAzjKEFAZUE0oqYevzN
HJJY3IoSeItdut3rhMNi66IhIinWUofjm8YfpJ43EpwvcUd2a4I/84ND3DF0ywe1
uuaWVmF4Xx+6Qud7Ax+AzgiZnCyGxIB9WOesYdjdXpAlpvXirLQq4QF8ytscb9b0
dZRam0uPGAQF8L/LFLt18toiRcEOcx5bjv6wnUhw3CldXcCoCN5Vxxq27DTlIHUX
L3t6cgXIvYJdXR9E1XEEqZy0qN6XOWKZ9JUyJtXmt7JfECXTioAV4Na8O7jDmPiG
wnRTsJ3JV9FEZsw/wZQYZrmA5jskkjxfDoImEEO7A/UCDTw3QPshqSnQV+xVymfo
z72ibmLJFdc1diLmynHPvI832ufgXUUwWbtx4XmmALdnEazjmd1cyPE3FLckdZHF
yWNZT3pI0pO59EV+e65SfpJjqwDfEpkkEz5XlSAqzd1+WdxWrrqVAyIWMu4iJye3
JTfqjffWUswspWKTxk/Y4Zc+DgeZ/WFywS3Y+pXoae8J6J3/pdy0wHV6/WZs64Tx
qi3A0qCi1NJ4j7Ghp/3NMegvbpQ2yNrp/iwkhBdYMB4/VSIFZEaqTy024g5CzOs2
drOkMqVwKKQINSAZZS5l+v6vOu6ahtxoGwHiYxtJrxn4cnOwBW3wsbTOI17kz5CD
93jH0/hASgxDTx/Blxuq7EESf+5OGasJb+F7fOxjqu4GJY+3eHhAVtje+7Cl83Ip
cLjrmpah0mq5JUuuP+tTvJiqlN24IPx56vJYLIQvCTlFI3CUpH53Tn1G3FCCvIUN
IZfCInWukJagcAaTvJKIJ4yHLNL9ohaq4pWvwNKQMvGhe/1O7ulqjIj7Ww1XNSOS
p/JNUc+o2L12FminhoBlxT7tqyCBEx1hikZw5DIrYuSgJabiC/O/0JMMhUOa0nXJ
c4Ui9wPB+HJKv6Pko41lFAm4ySrXiTTXdIhO3ZPOOB10cgWLsrkCmUJxz4e5DpAt
2kKsf//XQSCccj6y1TkcajnU863q8qCOz53rzyhc0Pqh4nMPIShqiLZ5onMbqcre
YgWfPPQY/p89xQRGCHdkwCm8Iw6TFRi9vH4URWL7RT5IEGg8hinSxgUOnUtB5ecT
z0lAudQ6nv/Dd95aLB7I8D3T4i9pJ1moZT9RxkJFLJGEBQPkxvWvfqUWfbfWCo8h
taqZmD0wqEdDuVnbD9NCbxgC53HaYOgWmo7onEu6S5vzh1HNLcWtG1ycE7a9uW/Y
e4dwzlspJiO7o6LWNakhSV9cMGDl1Apr17xwgAzsixZwil1h8sNVg7z5sem6BhHd
B1GMZeDfnxM6+k1vDeDEFls0ba9ax0GLxvXc9XJZvdA3VXyZwnQMWsIGyUiN52tb
jpZPnTzVGK5IFpFAOkAkpJx3YzyJWgkqTk4Bhs9SFMjLorqShHthZy7WGwh1vikH
9HoRMmSw7gvq175aE/z6pxoBXfDZpyip8Su/Tu1J4N44b1qiASXqqhoBnTa1SJ7B
mAW1dAUSJFQ/KCGML5cEYeHOCPqgx8XDK/D37orIBp9qkGklAPwXMICr0oh3hx8j
zCBiB2VYAJITvdGxgJ+kjOr5LbjijxaD/dKyRcbcmmo3XVn3lYueXLSUxP2J/FPy
o+vIvDEuMPoPvsD8bgAOmZR01WFvhFv92c8lPYve33Iz9CISOy81uBmicIDivhWV
Tj0gxc/55oHbnuY2b6xOEiXKJ0HAsaJb2DTYzkZpkW9hAOBbhuVMxjoyHgAv9Q5j
EFN/lSAf2F8SXKhHiAMVMOi3lUI/O8UoVjKZOghAxfmSWmXWOkLuQN+GVLQ8hiBU
PmwrRJqv6PqtbQY1m3vcYQa/aBTi0264KbBOpTWoasf8942sl4N/gjxOpHgCUsNw
PjMOmBl9EnRFTPdiSqxDSL8bea5CIwuvsWAS0Z9VTdkqAJYw3ZE76vuvwDR//Zpr
cYfIy6CVUCddoJmF65fOkmGD8RQ4Va8ht58+aFP44/xJRL1Kzc2Hf+lPhTr0/gZc
GuX9A8SGeYC+E/9WbXI9Q035obFUKj+1NpZe9yNNdyF2itRw3vbZgJULB0zlMhrd
9dUDojZTfBIWhAjUiUf2l0DXTGDyV3RvNS8s2B2QQhtQdozBje1h68i44BDDiaLx
crbiLKGOMG6FGd1fvm3gk9EyGud5YerbX+4SQhJnae4ZxU7j/AcyBoxnz6StX0Xd
jNC0stU5dX3o5m9i/6Y4W5ajkRLI97al1tYqLq4RCaf6IOAHL/8Tf1/pLkXqE3n5
SXSNJ9vZMmEM3JjKjbLK/2MJgLDzJFZtos0K3IvHJ9dB2ml8Atn/AoT3q5JRs//s
C6jan6b0opfvOHejQ8Ueb6D7erzT++eojgrX3KFV82cQodjF13dEPhJCm2qYlVZO
wdKSYfA8cdswA/qV5Yj5DglFJj7p7074MQZJ0WSZmBRpwKQtmjSENIL1pGyW4GxY
H+7s8NJGm7JijuIUsAnW6AfF8ArnCjXVhqmzUhvgmgSbXUbfnQufPyKAgPeRMjdm
1Dd7r7Cvz3LSOb48x5Tzi6cNLSUIfOsHxYcL4HY50JSeBY/9lSXEJoy9Bpp9XPXQ
BE48ecvsqy4Rq8Gqlbob1/hOsmJ7NOS6zC937rC0t1ug2sk2l/mmH6FfRzF0p69U
6WFkzv2j28dfErYYr1WvzQ7laC6/x+85QNL/p0L0lPVisJtnEAOJiEuTm2Nacs4l
fr/HdeDe6scgUfEhcPE1toeMh/2MQWv6NV+3t9EfECxkIOR9vqngInIXEuBxfnII
F3xjhQJyoo7Q/G87o18q/HGtV0JIAmnNF44+pFLcNsjCCUbipx362wZgP772AXH6
RWoUmQASs8biWoUqeVP74B9Gc5gn1x9e+sdAhcQzYBSRourLZ69N/wVRBVnW02Bm
KtWzSX9Um852OVCaDaZjZyTcpQktVE9H15FaY7qMt8l7s30F5F3nbF/SnJs1Bi7a
uQKN8FQAmZYi7e9XlCmHdRwxqNWngu9q9KTdct/QR+08qnThkO9VpyWjEHyTsE7A
eTsk9C4k/MQq/hyTABHCY2sGeIrmfWFigPUA0XsjQw1OZ2YxDbURPbJ1lcU3bs+j
9RhvbcohNO+OCeysVAUmyFmMEcY0XKJqbGpQKNqI5RwLx5FRG1OhafSi0P4lpmcK
Gz8qKWZoCooPsk0Tb2M1hUTxPXVfhvYk3pk/5vzG7i+ls7J3DZS4U11dZUdSvSdI
+Xp3tjAN5yLCv8HLZyeg0jc2uiVzGv/KvKJb0VPH12kxFoM+w3hoh+skUhE3uqQw
ZoBVmOEPYJ1mzTzKlgNzAX353t7WD/5lovgNR4n3rs/9q1iySuJx8aKZvVp5ziVN
AvqNarP1awYF/EV/XwzHeCWpepHRP7RK2VFtnCfk9jkb/Y2J1OXa6/GIKDwa7ntI
QSIzMYvSGcdYkKSNcVBDDrwreqAebJlkX+bcm4Zfplra1byDzF33dIweBizFWiR2
9zVYsqfLj5AHy0U2T3v64UNoc4N9cgr6Aosb8LeZ/HxogSlEYSj+Bp1LsNWL6fqO
q+X1G9DCpoYG3OHkTPCYKOJkUIKWzaidhQtIkS39AkTzVvCj2wzqj5mFutfc+qmz
yIMfgF9djvO1qRhqL2tmUvjEIBCoghuDYXoM8oH1t9/kK6O5n8pCsnfkWnAP8J3v
gqR8HMX0JGxWtiGMoEvaPenrwNmTncLg+WoKLOkjV6dMa5DjfMfkDf80bZX0U6no
0lRIUPL29KMYGN0klm/5HQdNsFmQEm9GDE/kMU5cNo+iovh+cRLEa9Kvp08y0HPK
XdpXxrjli8k2f8vy77Z4hCIhEO+78et/pkGFDtSP8m0MLfWZixVMqfKMysmh8SSq
xmZOni1nRL21WLUzW8q+gxAmkg29sqTHZP8jA+RMg34sSyqL2kpEdmhBVQjBCSDa
iRQg3PvNNtkcS2p9uN9Zv45EsnwLcazIhe+2g8PrvilTZ1I+0YpHyw0gw8r9+FFG
7IHQvmJUH9U+pNYrsyQiB93s28qW4HMBq0kOA99w9ZpH2CdGPNvjx+rTPFhfmDVq
9MjTv7S+EJhixLFxtMvdBdyyAt71Exi9FHZEPy88dmUxcdfytXM6bf4n3T6aHPZ5
iHeSKUL/twpnzVY89DZ8rDRYfZXZDAr5x096QoHGiYjVWRgxZOi7KQIsj0pXCT46
Q8jGuifqsrdlMmfnaVjkfTLwUfkXNhUfWMzbts+skS6hu4ymyOEOfU4zVOqShA59
c824sloh0Iib1g5G0mUn7ooEZMHsE/yTg7nPNoetiWEx2Tluab8sSLXa25LmfUB2
woz4k4jp0fhW5I4cOcC0j1TJ1xyrOIy4zIx+tyEopsF5YMsfQUjxARaCEjJBUAzP
QMUZN6FLACRriXifCql1rtN2TBtkPcZrk/kl7nS2GLk9fO6DMZGkDyzA4FHs4SD2
uWpK1ngqqYl+f99IXnVxgmmV1VqJ4KoX6XSiNB3q68G4Vfsbbgj9QM48J8eiwZq/
OIrO5SQri1xhN8YF/lp4RSKhN0f1DlvoSKcbF+sikJ8t2iIFrYp2Pyn/IxhWy5on
SD9nQrlcjHog14GsGcnl4RXv9j2tJ7oWNnJ79M8S1FzBLFahTtQoIozrxA6oaJv2
OC1fCIwsJmHajPMSj/OUB2MhhbjtV92oUNSNzqH53cTtOwQE8e0ehOmjKQmMX7tf
O7176NCY3nTIgSNr3Kyvz0zjvxPxxZ2mJIUVUQTdTUF+kXRas1Fd0ftsJrd9+Pz3
6SamSilzuRuztEeYRv2ggdVoJ2RmwTnQT7BQCSPQ3jTczEda4CB9sOnVP0oiAbRt
dA8MTl9ljqtXTYZaiRA55J0HSDo8j6CP2LjU0hil9MB1EGIz7Uz9THhf2YEQiYbI
Uty3wtFDTCQslNP54Jceq6mXIDMp1TgOI0y1Nkr8aM1+5OwNw6A8iLUXwgkEjHba
xGIIb8hgdzbsUXI1dnA5UGYkLE/ennmG7rIKEhfF9YEgZ7DGMoOiNt1DEyBB822z
wy0lQo4Fuar+f0EMB90ZGDpffJVoSa5Xz//wyvhVbTWotEcgUbKrWKoaojamlbYI
PuVHd0lTJJSXi+b+0Mai7R6U33BgG3uItdxTxFIIb8UlnqNAUYoUbNSmudOYf/Kp
BxqjPaNONgkLxkf6bzWtYc2PrxdaZngxpZJg3QZkidTwl73m7x6Wm30BbSqqOMkW
e++AEfy7iFPGaLNub1zZCHF2pQKxL8K22GiioZT0NObjupQ12nXsY00m8Zbg+u4U
4jJuOjkr7i2aUXEIR05esn/K5wiC/ZNrsgwfVfDzKIkT4davi0xMbQR+c+3tVSIa
ln0sKa4gCbzC4It2a6Y/BEXGYw2awfTTpYWpsdAzmSinnHukDybkL707SnJ4O98a
XR45rtyYbbrQMve0g7BkBIYWzKkD27ZOP8h6dWM4r2x+cchvYtiLfEfyfRfJOrbg
w/12805UWKjxfC5w88F0w7xyNO9HcZCX5iP9UzjstuHqSVWvIY/JtPMe+uhU+pzz
flTJZo9p/b+u02oaZyvDSmZ6HlzHenDFMrczIpZ/E8u1tygtbWmcVV8D76XFLMiT
m8P7vc2+a16HDUQZ5jvgaejftsUwq0IzwydGBz/HdR1XdXEKAwE7qZqTfyXHFoIO
pLTQo0ycj1Zi+DLqwsWlbvq7trJFEiFh7FdnKwpVyTwbZf/UrKVcXlCSLGhlE16S
fgFZcE53eBG0sDeJOwVN0aTcja6KSrilzargW9qtp+MOnL7XHNyWsEzxzN67KjHx
TZR7osy7wxJ7CrBRRajDrh65PQT385CNtqxksHN6m0jNWszs4FSbEC4fIksxWY2I
zQSL/Phk1ZGeYPtgvqbcPRCuWbfC+cgywS5i5/ZZ4orlJtiuL6xqPmyN8pQd8I+4
MAnx4JzDmX+ATiqypAl8CPbIhchA9AMqScMDbKidHXZZqDchaGvvVE4vM85qdQAP
uUAzXZr/MTi1U87AQok67v4ur7xbDNVGEO5HiFrh/XtxGglD7bXuchI+Exq4f1dd
WbGl0Umfp6GUhWyds5UapcKFZQ8plaKYYuWCzNtTNz6197tlQ0IPOQZfkw/jA4JP
8J1gtkMpINJYjiVsCOVGmu+Hfa0E8KCTpZvw2yLMzI5ps7HGgswofoVg+rkpp+Kx
v7oAazHCRWMA24wHPjCjPnuvCp3g/nKtIDUMrGp1BlrA9mDvktazVo3N1D+1bF26
GzBT/KEuxEpX9dLt6z2VQhRoJFTm4bZDssya5wMVr2nNuHJ/IohyDCZNISWSk1HG
DvoAiGJCaRj9ii1dq9zUjOYCJRKzK59c8SGUlnd0IzehpaEci98J2rKj2qKNcunR
42kYxcwTcdi+XT3CU/xbpGmMZ0RhhrQ5ZIKORBukMoUf4P/XSf6aL+NV5JKEMvbb
kxeVlCJFHlB7csT0DDSEXX3kSDtJeZF4Jv4h7X7Lhf0Fj2l7SR1WH+WW9F3SCRCC
Or7hK9ztt4DWgpbnHgdwsUAKv85ax0R6U2FODy4VybKBHhrhXQgqMhduQoUJzkZI
TOQJkrjo6JDKhFvw1F67UWDJh2TPOsyQtGXoN0Gt3stBKBMTVnCs953cVDQGauW9
0sZe84KqcYaI//QuZyGmJVTd7tn0RDC30UbWhZuRoRow1khswFrG0HIYP12cawmr
9hQ3yV0PMugKH3XWmwYKM582ZwxtfHkmzWbe2cAeGlMC+S31568QvLN60Pk2vfUu
pT+PW19+rzrqS8kZjYv6Z2yACGPD8aX3hH9OFaeYp4BIsi1A31Dd+Z4oZnK4Gt7t
IDVYcMFhf/JjkNq917gejHa/WR65bvyqHDLocWrOyOm7Bt+Jeak1BwIZuGWnhIcE
agT3rllDvjFczt85MWF0O9O+R4HvJgPw3BuuejaZRss/idEjPTD/UDxhxVDRtV87
0l4SNZoYiPAymHBMWniH4MIEtVRfnZi0oeE09NG6zb6tIpab3kTF7P7yAXS7EhgD
tMrRUl9fIxdnW9oN+perNnPRPhCRErlC2IMEC0WpJ+osAWdX8H6iZaM9ADdBawa/
5VzV1xrl0OgGhETF3AjoGfKHF+renw5Iu+g2ajEF2Z9W8aurnG1SOz/I1FNrn8+Q
EJiMAu/qHXRPIR/uI6Xo4zlA4jUMfee7T5D5+OX3Nm4M97x++jpDTMF6d51/E4kM
dELAU4waK5TFI8zlEfxz3oCgyM8TVoqY/8Dpkvg6BXp4mN07ZFKl5PWJxiZ4sdKX
Rao+NY1qFCQS3H9vqk0QxK4IyRAOA6va5Q5D3tTxYOxTrVdo5vtBpuZL4pCAWM6b
MbjNAHA9WHzW1qrX3rtyAgGOCDTsXGoNDRPh+cP3p70/WOP6r8xzk9FQLx42NuiX
QT7+NGtKkqLE9i8sUbLYBBsc7RfOglzTEUKZKUFYEY+Z/olPsw12bCqCHAvftXnT
LbvTeM4W4XWYkjdW5z9qdZGzfAtgIUTOnqdn8f8DQeJcn8QGiWTVhM7bsIUFFU1B
zAdYvZtDwrACcENTJO2+qkboehF6e/9InwjtKBz5cT6YKacuckOfcQhSCDsAyFuF
nYL4TidIBmLX2m260lHO53SUdzeyEsnpR0+CrP+kHj1EneedyyXMoL6F/UQ35yED
uKq+oHoCp0t0umxPgcYJ8VjKEXETbA8JYSBKK75lIFU2J3PFvXYa2+1/xbEFoldS
QuWg6a+ieU9WyPP1sP36nUb001m1seeDA7jTlRDhQvhbiayCVkJKLlMeYgerAuOw
9JYV+RHQAMZHYEVhHDxPTm32VYv0HWF8SoRvGkVm9KgIfa0KcJHJJZiHGEbKyBgx
jfseyjGVSYE10SamiMadYuXWAwMAsBddYa2IsOEHZvjdA/t0S2CqW0Xpnf97Ymkj
93zO1Bi3uq+BPnKfD/H3IGR6uszkZ6zTrzdTXTpa7xaDcS5fw4fdCiAdxvpo75Lb
fpnf2/5NbunXC61V8NKeyxxypPXJbeEUrRixpwNG1zVHRTgWj5I3dFp5JePPkG1P
WefIa5Zd49eCdem35EWBcvlRUIBkgr3Viq3Lh/swE//d8snYhgtbms1PccDe44EQ
OszdfxJSU+5Z3Dp4ufHXAgMrQJr96twsr8OjT8A/nm2x+YCLM+CyV01fZl786ZgO
B7C04TDCGlis/boJihnMh42HuWRTJB4pZN34WddtgHnjdDaQ/g98JiANyxF7b9Qt
tpJcbGpiDrkAUVHGQlpTLiytdxlqmXZHOrGVRR5P8kVBeXd/xweEszb8isE1yNpx
jvSnD6WiM+fsQqdl0dyoYw9KSXdNyUZBULaBFcl7xrH0hthqnrvntbe71dIb/BVD
jWW8ne3QDVTeTX5LY/lQ0MMYFmqfdT7FNGoZ5wDW6rX6WdWnnddrm5/vAxedSowB
QUa8oHChRL7iiLpX+p9zm5iJn/Qn+VnGaNjlDpAq1iw65ihommw9fq/IZ3fIg+DC
x+6y4vfmUwfzuMcufyrS40NPuXq72rOqAjZRE/2HK3lirdNKwb4DeA3qSsJV3lJX
qjqlMc6rHoSDP30coP8cEGlO1vYqcAXZUgmJBsbTwBe88yC+3l2QjcpH8870amvV
aXUtzNaC2kpRD2WhxsjDx46kLTqpuPm4TJBdz41T6vYytI+CbgBd5J2hrcLz5iKj
tvGIIAe7+tA6/iP3FIwSpAA48XwltV2J+fgq3kW18gqw7Oig+N9IGJ1UW3OeL8jO
R+YH4sHWAD0RXpZFPCZfpxM/vudOdrf9LYpsHZ/V/3UytCSGSt4Serk6lluCaE9D
w4OPS4+L6j4fzbIzenjJRqLzVVevd1k3XBC0nxUlRwzcTAu+4OaDnmes1O/+p5yu
rZ7HdfVSdo7q/u4khDwaZwXqqa09D0JVs1HiPNX8CJAXa2GKJ0+xc1sdYcDGcBoi
WKJ204WEsJlFJoQMrUqcgxcAWkDtoS0mRePLfdoQ4vy2oUJILj9opy9vdk6IShF2
8tWKg7wujmAjsPxsjOiVyBU6n3GAE4t/e0Yh7X5IKqUvwntekl/JnoH5Srf6g+K6
fm4P2T6taWWpxlKKdCMFWeRmX5sMXZrhA7BqHD5pDBsOtOfPwWgFzflf4UjdO+Hv
0l99Pkb7Tu6096+q29CqO9RoJYQoHIxCLACeHpV2akAdrKqOlEkmp5feio7NNEQq
0DdRa7TOGpq5gzHdQl+TBR6Htmv5quXTwsuvNFtwnFcnlwzq4r7rCXG0Iea+S2mf
GlUSnsT0LVBJIzoSJPApxyTNRAhE1lw/GfG62TooR45U0Sy+lnd6GzWdH/WOrj+b
+5XP7FjX5VbvRTOaC0KUnE79bG7Aq8HrjFKIVAqAJjp6B6mB0l3se1T5ZrklrotX
wUhaSaC50/gvtxqnFIlWElsa569XdYnl6SZMKH0HnlPjqgezMoJRSkgjqlAJC9FM
yEWd+CB8b0Ta5nfkkh6OyO3WsSNx7hcAFG4BdJOUuUdqCA8fK39WX+wgEE2cTrkt
/7Mqq/C4jKXDiIbNfh2Kuc1hQQ5OXICmuEU8dvKFILVM0DoEA+fL72+bN8eUBX6g
7grL9d9MrJa583BiExRpX0l5smtUUWsTpxkUbKud8f9dhjtkg/CDzyl7fwbukOON
n2ezQeUccPOfDDyc7ne+RldiCSLSsrQtOA+CUTbrN6iAqREa1xOn+bX3/mKxQ44R
umtvcawXdwMc0Rymol9UnrSQMyizpqMnMVKZoM6N3we4FyY11kvPGyXHichxXiKp
F1k+yi64iDCfqI5FwJ7dBpMLRHqJCQYndbzMt3usTjQzRav3jtGMOKBGHBUP5jfT
0cVSItti8hDOuWGRT27v5ioTvxkQm5Sjic7RaDvisN1oUJ1t5B2+6ra/8UiHtsA4
KYCZhHP7X6ZvU1D5vRZhaW85wjnCcrWrCvz1y4Ug7ZMkI4eoBImU3hNnEMuGIlZf
3bwmzsNmS+IN37dxo6L5apOFes0Q7Q12LOdT/PpSuwi7XOmli1AV4uuAkRoXKUrm
QoLl7oKPdqY4TnaS4OdkrXhpsTrwQBlV11NlUf2onF9fNOR7irPfASUchrN/a2mk
skYcVlmtGJO2C7eTnkJg+4AWVctUUzhitHpwlQXRhTtMFU1KAetDJmdqJvo6ufcV
IBRNxTaPnYgi/pTE5ZQKqci5NtRTBuVNIJfh443z+U2saCd9JSUG+wgFGV00xsHk
PXjmfJSn8VmDUio3JCK2UAEtE8/ZA2f4BOLeE8Om+Z1L8ILGdOfGUQgbzJtX1vRb
y6tirbxeCQpqzk8yCxafnoGElchMK5tazJzV3sVtchJhJcSQfTppCnyRKws3fLuM
TdJPAaTeSmCH1jqZ8g1D9lZdVluumTo0+0NFy5TUCYtLkeddX1TqqsSjabqa6+0J
ef2omwWwT1c4o2obsH0OxbkDFLx/HyZW+es9yQGM9tZDR6dQRn67SCun86JAhMpZ
/w5N7RPAYD4JxI9jgyLJmgozzvKx3nqD7W+GfOAoCzfOyNM35eRgQy+ZdmNNvVUl
d0PY09PnRaBKLvznEitgCs9rp+iJNE0e/nBML6yOb+//moz4fKMl86rDimlt4GUV
XjN7yPyED7l+S2SRwtN8td76ScHAeB2y+IkT1IKn5kxRG263NmILvgs+AtZauVSC
uvN7IFjfUlMMEZUHLzu91a+UeGgrEe1RP1OFAWVNakAWg1920+pz19GzM2Rg08zu
h/W2cr5LOlugPnTkpAxq1x4FKYXDwb5gSio6nT4J6y8fyDydaNf0iy1F0X0bOCbQ
e1vbATEWQ1vCOO6g0t6xnnbk4iF2gi+UPKJy1s4Ku4FzKka9pBZHFGsYqqvl5vHc
0rEQxA57LUqeYwhsj74I5kpFQZnvABzVDSHhUKCaF1065+zL1gcv+yi1hlvLeppN
jNRoNHr9B7rs3xzSKG8Ui2/2F0le37StW0iWmKfHXgUxA0qvOYGLHtnP6cgk11vU
Cf7WrPDUFSrpjfiJkRbfsN19qgBcaiSNVYvwjmkGCe8AdhoKzit2dO3+Qvd+zvs7
8Xv351k1tZ87pA8vS5MLMK3mA4sWaBrBH64yXpvRB86v7EfqyPhWguglL/u/tIiw
eOWM1EiILvGw8EbEECvsRNYwAnN6LpmkmaeQUBaeKhoCTwVZiDRtkp2oycKkjVxe
UxmcggKhxD+Vv/f4SMPxW/cDoYziBMeA7n1fo+vBZZHA5dZn4c1lzR6kISEjYg4I
7RJkerjwJAaslVjKZG3VheeyIWpa2bSJf5Tzrd+ruq+dHIWcy7q31vorAyVCdKH1
ndTtUezkL00yaSqQGLCMe1nsUMGYCccQU+ZjAgkjRjBfbWZ4lFn+cWeN01aqxlup
tblDGUwRRIiD6cqf8kHYp1Gsalp9reMyJ6QeNLC0ZeaKdOg4iQljG0rxMCehsEbV
Uh5iZyWGMQ+ttxrXENb2jz8BJ/pu2JklDGM04bq4XeEA+vR66AES5Oca0ZxvI/PC
zeqpR4P5j4b0d6CwMyyjk0wtghJchANGh1McuhSvBoJEHQMkPFiM13FcIxsdApMh
Hki6A/buiv1UYLfmhH+P+bfjgbTsY48eNz4qLDHXNDfs5qQuUwpUhR6kT3jxNzKE
AAPMKRuTGfXNZNV/I6na1ans4XkDG6F10ska3yiP0OUvEB8b9Xyp+9xnQiGxbYKG
rZn7q9t1uB36/ddbKtwomXtoat66QQU+Tbv02Nv88r2zEK4506kZMkAVch8ISCCS
j15lAf+cuSlCGqkZzVDYqPXW2kGyqwjjSc9JS+VSz8kT6AqYxYm2PR8ZfZWei+8f
ZoZ75Dhz7r02ri7OcUXcoVIZ++5hpoQFbmLHLDDIJPDQEEpe9L2p1rDliI/VSp9P
35gaL7GcPC8js33zGnYAcgIwqxemEFXmHeMF4BdvFAoUDO36Lc5cgbAFw1JG1Ygs
pNJQklvD90v9yIfxEx3kEEvmJGC31BTEACknavALRDToVTzsQwU2ogSZLqyBgmPL
I73qvs5bReUbuu0UvaYs03elXwhKYOwEb7kZdRl8E2h3NKINmIwGv9zIESZ+RzyO
roIGqubMBDNY2A+r2w5wOK+6uQatmQg/p5OB2YrBRUx+QD04NWKPpcrLM7qknA8h
GDJAocHmA+vn9H5uJP6xNbTrcHUvRpFDVG8v6hjgFB7VwiqSPLv/huDASB3sW6jV
7IzmWBShvUgv+DlavqrqzkMNQqUbkPLEnCyhiD/dl73w7Fy7PnW7ff9nXUYhr/hu
esR9XIIjEfJT8BcCo29S4wHlaQ0SgbGaTGMoolnDfIZF0UWxGZMIMTO6DD/aku4z
Vj0X0ml2u+cDKtDjbQOp1xQ3ioovdSYYuUq58O/1jxFJTkHSofQEqsFgJWNXt+VS
jWZ6FtyTBr2Vyy6tafyTTWER9OrugoLQhRa4WMlV1GomwGBB5I+eoqUYlnK2TCvB
K36HucC+qDqpgIRwP5nlUy8Rs5dEpjnlxAhXyN7LybbweTp189tXCRxfUZbsgTyt
ZctTBUdE5Bdse4hr7sAVPQcnemuhTgF61eanYUgRmKSqcFfaIs0ue6ET8QqUfP+q
KsLdZvBoljnE4AGIv9xc6ny2HKctU61L3Sn6xuUf33bchiUQph7W0Miylovyxilb
OoQAzOSzE19PayZQhY0BWCBTaotHvQia5PoSYG9nMwb8bOYdP9Bsxap6WEtb8JTW
Pp0foIXALnWphakdkQbPKz3GD+xuPiNJlpiQFgqjiEcJBTfHTvLIn06grMIW0Pvs
DpMvFAS6osT+6B9n/mQtBn7jDUWFE+XEHcyok9l3Zm1SKtIWqd45QI6gF9lipYzl
WtUZozh93sxR1vHUW0Y7WNYB8qx7eJ3nw24y2cCGk3/9JoAdnofCfq/xJR87ff7Q
gjOdAcdgJhqyGRLcE9Wjj/PjQa3Aes+EC+XsMEpaGMj72XFFTwwmxhmIfvLWlmZL
RtiCA93v3jrXEmmfxuRyPMB0z1jQuRyCcx5wi/7uTOkNtQTvIiBDxORw03RIETwk
EcxCx9r0aiRy2YRGH5WS605o957V5xj4NfJeZ7aNHDZedQ1sEQPf8EZeGsgqejAw
sRlQHZ+FgUukdyTgEW2sTtIKb/+HQLqzEJmHdjzV0oYPZf4hfPmjUPdnWADanb3p
tLO8kH+RbUun4OQ6Sx7XeOhcuj/zLDOip3dRMyYEwu141PADC5gSoG+FNccjwqfs
iIGMmf5XOI92Ft9y1ljgCoXSAt/XT4viK/bNoIhD93g7NqG8v1/DYMU28cGlf2xA
Bt02HYk3TTanuC/FeI//Bq2mZIVR6PccHyax8q/QdnKiz8PNAdcTjKb2ndBazHCH
yQYlcbvhrLbLHijq4LbCMWBziAowLV2hg4vvkX8aI8acQuuO/UigArUZpweCzPlM
y/kBirw+H6B+hQqylC3Q4A5MyDvBK5Amm8o7lua2R+JyX7KKFG2n7CvWbgDNDl2f
LUe75YhOnzwofjJNb48Xx2B4NtskbqhDt/CUy22o9YOc5lXQKQ17PdfgzLOY15hK
b9tNbl+lpb1eD7hDs/CmjiOtHnsUEcRZH1OhoMauPvJ1XAhb2+kfa3YXXVFJeS90
rU1Ed/z0eAQ1S0pcimtVDaS3htWndV+4DIMBr6Bd2c5KEJze+UnNsGv//zPbyXy0
UvISLIZFu4nSYu19Z1izDuXCjhCsyAtE2nV9INP5ssMgUXH/U9FtwNJDmv2kMsdO
PCucmu4MPV2JALvZmnACqufL5L+R7FCrCDOUet3a0qH5/DsZ3RiOQqqI1uDh/Xdf
y15vANMUfUq1WhcGMtD0XiaAwLQPFpcSbHqk5wW/0I5YMDXIwqcOma43/k197TKY
PLWGdEaVMup4MpaQmoJZVI/zX5ImBJLixGsSRWOpAs9qGSZ+XCIF22J26MSC6St+
b83Ch7Zol2+wRuuweN2BekkuUhlB3BEshuKgm8F2OYzfkcqzw1zWespTBrf/loRg
YAwWiSk31Ysjp1LeLu+M0U2GJzNWTbtZEP7CNwLqHYA8EHVS04ZreVKCjKcdyr4Y
ZpX9YXRr5DiB2sKZngoj5zFzAMnCehAx+HbohvCo1zpK5VF/Xa1u3wMIiUMUZXJV
nMdRGOXVAUHtoWk4VJ4vSjC0h6KTR9LuXIm0dMpakzUN8PYyo7p8dAP2Rfe2mIeo
mLS6fMrAzWU7Sh92zZ3vRxyok/JdzmOUhrp9YMnBdt0ORvA3/YlVJGVWAq6PW3Ou
geg3WM9mAZ/36ZWEGL2PmM8ArnTk9FFzvUqrxV6hhUez487B79xZ2hVzrsgh8KFI
5f4MR+8+tEdu9P9nvSi9FPcJE7IeBE/ohtQrvS2P22I9nzuYZMsX5VU8AGnRSdEr
rOM6DZeSfBO6WPYT5Sh/2ZgG7VOD0Bpq4X4d5D6JH7A48HFTceFIHFeKgnqpvOyE
3+NBcrb/xBQJRZrRpntdrFMLCqNgB1LiHxgzxIco79FrEA+gGQMHpe5fYAFJjWQt
0qTUbzO5+eiXQdQQXU4oTO6BmVBuBctRI4ejsxcMu1LHTzNsPBoCj6rlGk+eLEk6
Gsdmf6eTprE8qfvnNY61q9oe8ev4xIrMcz+AV49RnkRdB+fmMsjkyZUG3MIkM15w
e7T9Y+Qc4GTotBKP/MAoHl7w5HWU86GIqFgPdqmuF+NIQp22k80uTnWgEMRWElsI
KXUIE2MF5Ops7xDwWxjcIOPtfvQImMuLt3n6e1RbIyyA63FfRiz95BGA12qsROhB
ydnoQ3q5NG9I4BftUjl3WNHWMqNQLMrzrPfyg+i3GfCZwgScq2WRAf035L6Cyf6T
Gc+oSh4JNRHEL2oQRPFVJgZCP+t4eVEltfOf3UbiFrJEaR8IETowPF338tDZzrr5
mnVJpdIoqsoxZv2Jlh69kM8tiz4ha+BFGfKcLnBvQviK9zXXMh4HEJhq8TIXgQ0D
bTl2w3DM9584FMSRh27BPLhwU61kOgEd/gOCtfhC7WnOKyOnNJiFBgP6shlDPbqn
pNNCgG7Z6zPcPkYRt44G0TE3nJwHd/B8o80SJHjD7Q0RCnnE3+YXK8s7skbY0d8x
Lu1I0qkXFuMM0AP/Sq6ptP1ltTYHeVwjys4eQPHFAE3NgLOVBA6XTq4nffG08egc
3rmDX7LkmQLWjUIEgz3VYkmTC+8PqSa2beDT/o5B8KRSVrHLCpa9Z6SO/gU4Ht8w
bq40vOn2hPySwCGpBvfNoSqI5+FNScu/xgAMWTgRhP4pSxH+iMqcFJpJsL9hHcPB
8xypxj40aTodF0YOCpMx7VAVYFmOC517/Ca2nxyeWc0+GJIfTbLMCASIGbJ4l4PK
bmwVbc/HUWvGWIqCh44kPsh83RLtSVXZEemGBlvnaOcV/4bXYevAjEvvXeA2Ar0d
9L2b/T4HGTui9M8nTVtweono6TplkdS9N8E9vCnY9NZvitsSXmmPNDMNvp2U5nWz
1z06QveDbX7QJxpH6XqL+bEmLARNQabGx58Lms0p4H882pyDNrT4YRV90f4WVOVz
bhpY0zEY1eEuqJTV3/BeTZS3rPIpZotUGw2DD/IhQ5hJR4sliz/knUc2tus88YKL
Vprqk+8txTY52CoAi8Nokoxg8jQ3WqVPZuZZcqXtvmwmcz2AOtCLqQOVBA9XU6uQ
jQYfDUiMZQYO5rTCQHi1GEZSGYGb1GZqJkDtzWeOv9mwfS1rJJKtP0qca/n/kIKZ
9GtzgNi8l6NbPy2fOePMah8gLZg3cgOwF4Xmlu1SBWTPTsejwR6UBpSK3eSSCNtL
QNa795NyMtAmlf7gcmWqcFhNl7SSfdaI+ERASbASzFfjITKd4gAhPf4lV/40FxJR
Yk+e0X3YvCdvxW2jLoLwYeTjvqOFV3R6CQahOva751bNg3Z5yEcOsHkmUV1ZEMv4
RHdPokcFmGOoEm5ILG3su2jDUmNQyiySxkid0aw1qYa+SLonLyy7xkjQxm9dKaG/
v89ZM4WJqxt4S4U/gCCL/rr/OJ6gIkOpocwlju27R4rhR/vPiCcIoIH+ZlMczWNL
8mxPH25L05Dv/4sVxzwbXougcVHOrbs2KFGOAaShjBnVpkPeGZkApw+vbyqlW371
bAHaANbosszUdcvj1IkeF0Q3XnCeg10wOwSSlElLbHJXTNM+8lprUmx8jrrxDpYq
SeSYBtzOFADDhAeCagAtAmTx1zFH8P0DCEYHT2y0HM8Xn4UY78TYf9/1RdmZAKVp
jfxa2j5Z+tXWBO/ApFLfFGeg7YduBmkS8AnlkjPhV2YmLaDyt8EZwZBrJsNfpwTb
QgzDbm4XuEjZEnJVFRrQN7VSB/0UXvq31uUx2Xp97fnJCkoapfI8yj8zdzzhG0hp
luqjFUrf4tv5+BSNvAWcXbwtx1YMMr4DBHRjZuDGvt9UiJ0nK911RPwCHKzexLR3
944BzggSswoS7u2uwMEZUG21p8upqJuGu1apfQLwbblzy9LAyf1bFJ+W/0usik2+
FTbjG3MTg8ekW3N2vIlMV113MRfTldKA8H5VHImwP6Z9/1G3NypWBSUhukweubGx
0CEquzQD+WO0VPFx9c780LYlWqQYvZjPTI8o81J1DbJJm0CCehaotaKM+Xralb6p
moOPcemzjljSVzbDD0p0T59LwnP7fhwOxHwZjRTjsl2sWBwUJudMYT4wtX7H30XN
lg5tKsUxIKEUmUzSXNrkmIuN1xIRz8rZ1rS87+e3ZtAxBKZwCW7YayXnkhJkOIlE
n1P32yvgFv5rWE87Q1X36JpYQU5spdaDSbUWO0HbUr/22UtsNNejf8FnX4ogVbro
fFBq7Ai6orSNrHqDlvKslP4xwadewyOxHaPB+5eh7QO+9XMTk9NS3EuTl7ORVcnK
E2LrXZMoS7hH866cttzqO1bpmRYki19AHrGXIkd8Fe0/q4n3llOZTrE+yjoHUA7x
bFeCU5KcM5Hz504MEZbA7soFmMCTKEKr+xDU+wliGnHij3tONpD3g9z3BZVJUSp5
6puu4CkIPbLnavTnzYufzZx5IxZsdYaQYl51allG41/cGOtv5tEOkL2A4rZyqFha
V1oa5bV75stX6rgRKtimSmX74y1Qg+C5EiV4052/ZKzMUtT+jE+xnq5EeohKLp10
yEQVvl1vtssjPOgMtXgqqA3ECtwSJPPaQnLkVXI0T7gmDF148hlm7ZnAF5ZDEpRq
pdp5+9N3FNF5F6L7VVo88/LvjsGLbGSi94D1KTHzyjBzYZztA4F8SCgirtwpeEa6
jVOpZ5tHn3JNMuUq1Nr6M13/qTDldw7yuH4HJoYqa+eVZ/8ZuSwzqjkFVFgK/4Jw
kCzn2dROtf5841DKdqOlA8rdXVP+LtJEBPHEOYJvyE119lHyIFG6w7eokkQ5oI5J
PugSK46R29zw/R6gy4Eb5GnbvhIhgkuyMczNzJE7fKwA/Zcyh7XJowGQYKOHNmRP
y+jfpsXPi6jQWRX/q2nJbVhk5H+KHI4xZ9hpDLuSB4C0wTr9T+ezSunQTrzptQtq
Ty/vMsoHWPSuhZExA9Ug8KqLqn339yHsSVu8k1oomujhEng1889QT/J514mV6CLe
tD3r/ln8vIxMuuDi4tIoKgYCNw6dsYhdChmEpvjBCui+4X7xAIUxnDNnt0U+PbeJ
jaP0LpeCnvZTLRe1RW5SPKxJXzim5ctNAfUu/oMuSxsiwhVJduLYSR3crvWysK80
3+Eg2rt6Vw3A2v65daeb3rgoThsmF1u77JG3Z465El31Uv+z993vAQPkP+0eFJQ2
jX5T1N/antzcwV/18/2IlnRiuw8c1LQpiNVxa7Dv/6iQNYslA1lttEvL7V2jV7ws
1GFmgtinY6Cxzkr861aZXmLQd2FUUbxKwNLtbju/XVyDpklmj6eVf58aUWkcpGTu
2dECmf7vAMWmo4+PP/0TSLODz8+f1smXCXgnHOjxtk9J+5Os1t3AKwhJ4VqVT47N
qsd7iMEcLfHGup/RO+fWQMP6Sr6x7cWQgtiR4gOMKTKtKOdLRyIQ8AC1PtYq6BNi
PTLe9CHqjAlanoElT4AzUnmSoruERoW8YAJGeDcbzVZEEeD9+kMjmLu1pAOBJkBD
Z550mEupJEkPqFO4Dmu2DfofZWJheaO2vxpt4HAMpGzcnJHSxcJgzdw2J3SQpJkl
rzHmaAWzdVC2apvOtt/2P0d0E5a0FlFcwGx3Bw7wPkJ2N9d2JfBUMZ+Sapwh2E/r
XoGzcys2QIinsCikraQySW3OzpJHxvjvfyJb8PIUjWksgMs2JvTDgtrVwkNBd4fx
FoSjEn66wF7H+15LAzXaFu3m825eQrSkuyBWmq2aboKHe7Nbl+853GSJkP6ee3jn
gedZL5e8sC2yrnkyWLkLOjkpOby4novhLogaqCCYFOn/Hlz98FXe7q3kK4lwb/Iv
rjlUgrWQnFKIuui8GAijc3zvLPXUA7wRkrFsgxsduUkt7R86s2H4h3hNuD/DU0I1
g+d7XF1Vbk7Ro7JrDP7aD23JiOWh8ed/C0VFrOFdPtVCgCehZHyVUvUCsBXAYSMm
JMFDLvoT2PEA36DoOE1cJo0y4/9cn25m6okBV3DjhqYshVPgHjSaF32SiAeB/9fn
C2JOF3on6V3TTuNE5eYYC2QHJ8Bm0C1QH5iG8nfCFF19ppSWewLX8ZPxsLHXMMD5
UiGQ0IIZ8T7ys2ZUzim4fAwl0bPX57IVYyxQhisWuNKhswyNkeZTXWdSgpKASvQX
x8NFQuym2TwrGWM4H/ByRY+JkFeQ3eKZ6ZyiadlJ6bS4xpL9dDE6lB9HQKj4KcZM
wKcmmMcqaJGMUpFDmaiY/fWwtoDQj3/pLdb5RqPFMHZcWUZ98ze7jBZVI61q/GFy
ciXuecfIN4U3TMOwwQG2eTUhsIl4LtuU4WMH7YsRfUblgZhyGoH6ez+xDzXaibVb
FnWoCpsQi6OeGm9QnQDio1lmQ44NuZShK+hYNgN0k+zf2DETdForiTLd3/t++jmz
uQjVwZqsryLi50m+3LV3oS2fQJIy+0F7f9qdeRs3NEUq1cTWiRBJerpeulShyMH+
XXUsf5a/Cbiylfjuf9t9KhoSaeXAr8VkLnaVNikeJ/0dhuy5iUa5eujo94frF58g
wcyRfMIrT75sLQHwLlv72o7LzLA3Fe6PmwASBeLQmtmE+5/lPxtJl9g6WVT0KrFj
YdnPBCNXbCGacWeQssGb8jwE5OsxJO5YnmIJ529l9eYWqR5N3dLwPnTMDqnGHTef
eSY6aKzV+sGYmN1+sNt8+L+R3eprB1qMOKzbaTQ5lSG3va/L8mZ4yg84bmTgkd+y
k5VybS3PDacEBCpAnvrTiiZdHoynUGucImXrpRgIZgb3dOTnD0fVKcAsM9AloUzL
2VgU8yo+EXf5KmTKv7zO7Nzv5n8AGsNChGYXb2Gju7KrPEjdLjvLGvxWjby9ft39
XOxq1Ym0bN7w2ujymKL5WU9IyZj+G5gJr8xFfdYQANQk84jF4h8R45AFq7/4OsdT
yTqvh/HL+iQuJq9JqF4mMdqRp7GBBOqAj5+L/k7jxOml908I7/JOLd6d1Qu5ePiv
LcbbNnZ/mCrrZi70ZAMYeNs6m+m0+26dDCLbV93/FcAecdBqcGzpK8xTDPC0A8Fi
nvgRdY+ABG8RmFxCg/nnjCEvfr6OsPBnrJ3ERv6CIKW94oA3raIYCNrJwt4oUfeb
D2mGJcHpp7pp1obUpchAT+V2tl4KXVuuFzXQSWzzGRi22NAyeWngDInXqAzTFMJC
+GyLZEjnlKlYqsIhEf468sUgb08kM3SetS9nwZAc/Ra8srHz2+hwgT04F8mobQft
lOsRfMPVyRpW+63x1pl7akdHM71h1pIDrhQb7zWm7laPgFqmQDWk8ruxZ99VK3dX
x33Qa8T/OrUD7NKoXwpYGp3GU2oyC0Spcbj+ENbEzC/d3CPDxHtOTeKiWFTOofQ2
ejdgp39M6rcEpcpHTvH8+f7P/n9nluEDwHLzVUDASvTQKVO+/rygJo+5CtajdEZd
s3WjW/D0Xc3yT7SGVG7RQDCi45yrhz31OKKtim+xqxBEvSYLfN8+CJfJJ41PtHNt
hYR8JE9U5JeBkF0zidbUpTFxMMyjcDI1sNM00jXUKK5yllROn1uy2vI230nlnHgG
7NXUklTn4ZEHeNhrhGeAFwZzFzzzNsY646jkWgg9yCtYi6jW8dMbOcb9xUwXhnLH
9M0NjIWvQ9HS/vi4Vm/oP9DngFUwdt7C+Gg303jXdGYR2U7uKWG/tzZeUvvQek8R
RFLWUxerO+AoC/H/6nczz9BiT+B/k4h42ESN2OPWNo9iJ9x0oB4g1Y2wlq75WhYv
R6mAtZpNFTsxzyu5qb25R+/R30nKWyccV3rOw85K+iuafBX4LNeYtq3oB6b23nRa
uYsZWPvLX2lpKrINQqF6coUYm0NIriLVlUMc5gxuoOtu2derwXCDE8yByBDkVZhJ
0zy+0vcipFuHUEmAgjpiacMPiY5pCozveAqg1tUbalcdHCcFcRj7iodXi+7kvqv0
8691PIVkWc34R026a+/Qzc2vi9CgcmQZMElkNwDUfaYUhSGOYZv4XOSSEzpqf74d
6AoLY3Jop7SVi3as9iE3YVq6/xO0dg9a8ac5fvvt88Dsgwvku2oVIi9UA6J5aZqp
hewoY0Ap3vqDDT4CxuEOAiDpKa5Zlx5RCUxYFWUqUyVNwC2EG046MgOKe2QIre0F
Ok0ICBRm+k2u0TjtAD7higwBe1zi00b493a71j9r/RInPWWZAAtBIwCPYaIhj/FJ
AMtpZpmyua2BAkBUD6WRc2P9FgBdjV371h2dmd4Ekg4Zr3z+GAg3KQmhH7PVduAq
s4Ijhn8m6eerqamVI2Io/nJDbPR1gOG3UJb3ELFjU8epO6ti/dshnTySthBpe9yH
epvBfIlFZbJxTJUjdrb7+fNSzRyDDVanD9xyjMqDIKiy2oQX4ashYuQXiJLsy5kl
f6er8ctLvVtt80ykossQeFGMb/s9zwFYnq+oD4nyZTrk4riaV84I2Ok1FVwTBItp
n51amJSfjls6iR0KLGXmmvqSZQJYU5PHxTf9VnBX5aWIybXlfP+8wZJ42A+xkNoo
aIeFt/1fJRq5iWb9LrVFdOKS1ztqmfo7h36MrwChj5x9Xn3QVyhIP2FVGJNiMC2y
ymhukkF0EtFiXKgJ9kScWZuzobXMHP72q3oz7TmtGzlvAsWyiA8xfEyms6u6oj/F
2TwX9/k3YJeKvFHEs3Sq13/L03B527roEm8Lud9YlCcJi1Kv+o84Bn+2OIollseC
5Q4mO8ZDCa+02XTw8+0xeF3Y69FqFZZuQyfdti8wOc9a6YpxQNeyLvskbQO+t8tT
qyeCV+rcuAffxtBb3W0Hp/Bh1jM1KAulZdoNpBrLWhrSJtOXV/aXPrVt6EpONLMj
oq6EmZqXMB5WHO2Xyarb3PCyKv5Zrj2n+OtHPihrkhy7I1q449FG/G2ypJaxn0zi
8ngZqt+T180XTFyZqZYzBBTVSm1aLQ8J5luIRQARZSppjdoa8n/54yrG2ygQndlh
JcGDNWTbK9LaRFo/JFde+FiF7PsFGNMP8ASgMpgGkVFB1NuChWBjaJD/vTGB3Pmn
aKvzGAIlxr06KzzzzWiLTm5yhoXTE2f+N/h7ySI0kb2CRBVdp4C+rgdCw9ke5366
rVrFe0CvS9jz9ZWhnp+qLdzgCZmSub5rkISyNI8YfDW7dOSBF2XTaNQKMPaUCOqS
Ew5RfBwf4Kqc2e9b9JpsvUH1KTH3RYWJv9Al0fl0ZKtEfA+bYAAUIYhQSwgkCcBJ
jHaokEJEXyLNuNVEEIBY3XGTB7UwDZBFvG9QugKmN9ZKpNOY3fL53hNyU+d1KvMC
kIrrUIohMPDEP3gvxiBdlsyj6KgegMbpc473Ie6AGA3L/lhZqkC8zMsvVGVZ3J9U
BgPNGY2HOIq+hV781KJ47Xk+rDympE7bMzGKqdyZrfHxBEP1VF7qIeMivQaDwl47
2Sn4qTI8kIyaiock2EzE5OdAJPn+XFJ/cwyYNo7mvDvE6eUoB6r+gb6vW5BHbi3t
y6lcb80Lrveq8HImxtJ/HP5LcEaK5khcFJaSmSNYjuwDtPn42LPHWJB4O+Mbm4XG
JLzd+6DBpq/aGyjBVEEpotWKfcPJkPoLe0r0pPt+VREPmrzepX7cE4Eea5bKO4r7
jmd3gauVdWoh8bW9lRaJknjNzjkUUZd2IQ7MfXjS8Xl869rw5xBgeVwmbf9v1PGD
lDTKexXtdGq5hPxM3tKX3YOk91xhGDSQc3h4lC8W7NIATBd4eavHr3JF9AnGaXis
7B+gZ8lh7ZsaLx8df/GtMSTmyPyryqL1pRQ+ej53X76k9iN4VMdHHKGuTG/hk5Wm
ZDVBl6LBNgn32H01JdP7hbS0L7+gE11OzYpVoAQyTgW5A5Ruz70l5XijSm27BbuB
KtukboAzLRQpDWvkmO6kyihJxULpzCkFeiUcbmzyYkfrHV2cQ8rDT2ueGikXpTkK
iC6RFAPSR41IjPcLkZA/T0yYS/eZUhrNUc4P3N7u7+HLQkNJHYVSQS8//wj4zjzk
Pr00EMutKJQlkIQoKN1XsyAUcMrB/vIbBQRczQhvQ7B0Gyo9oUqB47DR5kT+Mexg
A34bwZY7ZKH8Yt8L01Xbv8bMaFPEz86+lfgzdBupHDPwpOa02KCjbnZDjdAGzR0/
C7KKp9XHJGgI4pUDv+Ml0XM8fFPTqF0CeYwdjjoVCTsY3qGosoCp9E9sZe6o/1Tl
Tjr8w15Hti+7Wf/oZaymSgm3fotc90tkIdXs+DYvrReWVXSTcRy1rK230URquS/4
e4GX2HaD1SaXNdROFlrJIvqy1RW84mwAbxO4gNmu+le1S4LiToPynUBvvJdjD9n5
5lo1DytqYh3h5lKbMegOfTYQzBki7dusRUxal/+JDAN6nFb1nBUmqsab+rdhk2mc
jIWqQvxHrZ4yum0Lnl5CWPmcKVrM3mjNpEKoKqVztveAtkUlkGdGL0rfCS8iAwv0
5FBhoxI6VA0ZlEy9sjPdQaP6m3zKGYXlue9TIt5nIRIOqGOrgV44GediVgI7UG3Q
b50aS9H3a17MQUBlDtgLAPiBFWjF3s1NMBFdM/uu7G1pHbfEE716OueT0T2Ked5J
ALF/ozoDNo7yB5zcyq5Cz44iR0XLhu641doXxbYBL4TjZIgmAR8i/KCWUdub9OA4
Vxaz3RuYJXDCEkwXlmPrm3GgLOhKnFLQ38wmtXTzHwegqykFMTF+vPQLYJUaFhBq
zjMVd4o3rmMuZUdUgEBsqEW6WiEDKE5HGtGGuRrTgdByvtOg090aQoA9NTCtTBa2
WFnceHRw7b20p8a+idLWSltOhJwHzTn5ccqVSE7fQhECTBsmuxuJ92RyVab7DaqL
JUfc7D4W6yFAhosfMgB4EkDA0Vg/sZSBLvgK8ktkyeUJNibdULP8Mmxbsl7RgG0r
4jBO8XvAHUzARxY1CvzZBAho9SXigtb2nrCrfqAjLeusxHI3JTUCae8Un/Kkwj2S
EsoVVJ4hViVi508Zc2jdht1thk5UYEm2TX/3xScuLurdJxGehmwjLsFAl+elNxsr
CjZwqSE/BLJTf+A6B0YjtGsT7shYPi9Yt1UERJ6lO7W5VEQKAV4tGUdY4o0fQjAL
F888cTqfHgYGWSM7ROL0Aqtj60QRbXtqNCE8bn9ZUS2Y3CZgNratvVXstn2MVifr
oyBNS6E4HIcwUeD6kUW0ZmHXoAtOY7ux6UwqxDKCgqu709XhBjJ6zgmwcg08eu2a
waAaVW964DMzlOqn4/SFuw/WNnWPCUjIxdMQDw+he51kIJadM+cyS7iddP3k6YdA
yzNOmdNoFI/rKmi81/sGDgOcJbQOfEqliv7sxOegNAQVW5diRPuEjJzc1//fjj7L
K1XAz/MiFidvnRCO25MgSyk13vFMt4ZdMZM8N9T3dZ8VK6zFrtOfzXGDve+SiU5I
H9VmXW2gh/b+lBTU5ZtP2wDdhztEBxiA9kdSMw9SPm0Il7FJdxVRtRMtkiCBgm2k
zDiRwlbnraFc7eerxYN8Fsync9lIBh9XyBY7Tv+2nbWJl923UXUV2OocVyC3yiUy
xbwTOEB828CLEzqA1Vfe0oQIKT/ZhD2j9M0JxV62JldwSFrMzEkjhhPCLSioXc7x
56yhAwUzfYsAu4bKlvsONGrgaC7GSTKwP6OKcOC868xicvmc8RvO4g9+1KQQuSKO
5XojlSAYXqvlmqBdgjDE11g3Q9XqMj4Q1+sR9brjzdRr3wWgmc5nXAxTSvqUUIJ+
SSqGVdZs3uBMpJujZ8H0Ck0mSrXQkdlBhr8c/coW5fZc8mH/hfGG+ILML23g7Bcx
EE70pWNu+/ss7uAUBSJNnlAFF5NSu8GmLaSuAYgbeZkeu4ZfhInic2FdWlXMRABX
dW0jFY8PNZS4+iQPDnEy/oNRwlaLDo0AqS8vIeShVjx2rgEevLVZXuWpcuY0BOI2
J94NF/hJqmI72xzFttDE0+2atyat8KK4lKY9bbkdPhyDD5h5PVG9iSHV4JSwE792
UcRnZRj/t0prMfAVEVQzrUxhXRgr0hir60GAH5gMti2jxGJC0kvsE6o3uVYbHgF+
771D28IoSdkjJ4++HTqj523BMH/f7ETeKrW4Qn9Ej09VDx2Z8ekn4fv3QKvAjr/j
OJXBOiDMD3djMsxYeiZ38HS8VKiBfXao4iRJgk22M2CkGCoQ9ji9nxPTyAG3ph6+
hovjDuciMUnfc0jzW7AU8F+8P7uiD8o8TfI0eQ4qwcMyMhNr5aBUXu5TRIRfGCXM
eL/ricTvOsCk34q4sE6ciolT3wNhcYI1UJEWHWoljm2NirieNMx3pc0ckEEQmkcs
/4albX+xAVQL1zX6bh9evbKtvuEBzso/GXSL8S+QrPF52hv8rak/b28pIQQJTGD/
i/NqIi8D98drCAHeHgJHtMcoQ4ZsYs385euDBJzT6NPYgpQ7Dtf6Xfv4wNL7YUfv
54vueRAicnKvWItG6l8DsqtkvGBhfBwst6r+q/i4GA94CxNd42q7evyYseosw+18
Tv9+u7BOlpUSxxBF5zDcELBQsNyP5fWePMJfVkbwaTqoo5PS/sjEer6BjvhvL0Yn
niaAbDhXEvZRdtn2l2m8zA2/WaojaRu6nT05PMpN9wrF6WsW+RTyUHkIbgEppxiH
WwrLewmVeIMt6ov0ug3zg8BhZES4yjnAbag3OoiDFy4te2O2bPHCn+1xc5XLSzWS
aIa5PTwVlf85YTV5RcedvC+x0ZjvdKKR/PeZ9hn1HGw0PKyLeTDUiu+EqBw6IL8M
EJbCnth3HXluhzb7OdFlymU1iXQvEhJLeihTbUk0XTiisTVtPuJLcOwguRiS1UPZ
f1+vXpg5ymFBg9tXZ3lPh9XnSnGjzN2QNYROvUYliG829WZjbqvv52zHYxwMb7l8
13LvZli+iWnptGjE6LoPs0ZZfP5IKK+jHmvRquUg7FpsC2BUuJ84+RYEpwjHsh7n
C+sQKwCKMaBvMEeeUYZGAs5AU+FlSRDzeTMY158+u3JLKkP4ACfBq4cKeYyYpnU1
sAhd0eFvRM3u2y98ljx282uWEa1iA4ckUBhmuI21oNIMwEse4G39neENrt/FO3bn
2qjPj0ZygG8jDVB7WapSPb5yvFEozOAFW0APgYWvCSGzEHwt7Hh8sT8ttzp6YnfO
CLp4ebWlSbaw5N8kyzYboNizC7dZW2Gw+jN/63pdU2U5p+ZVb0imLGI5sFuPmw9+
bllMPdyVAwFpBZJ6WLr3XTKFz5UlGQ+XUlRug2Z8q9ExWbDia+Zm9GlYdw1FieBI
854sqKlogpbiYyD3hEPRaA9u/VQvEsXat1rLbbqFZF+HODA6ptu3kdMD2S+PHAqp
1c7z3EJ5C5BTXzFCdiIEcf6+mMPVYEW9eFW7/o9r8bM+XQi0KumwFyuZ0EagZI2I
Dtw80iqgYIIlai3QHzJf3RjB+0W5fnOFSdFGtlNECqLJmMmfI7LSr9v8yNPqfnjr
qnz4fCGX0eR34yjpbzlVcPvkcPhmbxwRV9BGmNc6ngXh6gqEXq8kjYVV3utVoTDh
ND+OcUsoT7futfIofaAxgEr3hTAzC085Vnr1e6oFM6n2vfI1+owF1mQmMg0gg2nK
XPTMl7Jh2SwZ3RHF4qrU24tzrDPU66dt54y06ObZRvBILXqLOCnc9SfbTZPxAwpR
rdUMQBWYHhZLiA/H6R3+CVu1HJQwf7waHewMRLQoxtKqiKq4qle4BMoijqAjAA3v
khGmyyUg88J3TaSrDv5npb9IVYnELiuedfdUI7g9oLLGzQMGdAjdvAcVhODAJUKn
GxuXJnbl7BZdHpmmYUfH6+WDRDQ2ngN1eHo8a2bZdCBSs7eUcapvKmRPQj6s2nkB
yfGA0vsUTsCc3Gap94VCZqr3QuaTKqWEjj1MQ3dzfoEjppi36QsQorGUTe7GsjvF
VWRfyns2i+Ps6w0ETcdagKLFMgFlmpQUEsdLPX2Re6TsFNxMPOawQHtLFznv5WAZ
EKkLk7hgWkUbeF9ZBKUmmNerH8B58MHiRpZhYyNdNukxFEOaW0S9KfIr6J5WD1+P
Sw1bzmoy9Vd3OtW0/CMAParqRJwZMJzyq2f1yLVk1Q/Fsn5QIQ6FacXumDvS4GdU
Ffwt08WOkS5qDDO6FcWSWvNyrZgfdbc8xyE12A1eyxwo3mqyDYtsuwFy5Zmmnux0
nMzXCbahdor2dbE9+Y4hjiC56oEyV8bT7/ETM9A52t3XNv96UhIefCBCv2EGb1k2
JL/AYcEjbU9iTcENL9z6zx38tToQg00rPZ6x4RX/nGxMyqDxcW8tP0MCD/3+5utO
gXadTKpvxTGlHMEOQ6wnfaeQmD6mMaHmWJo7XoEzhNmCXt5CCs7g1A9dW8DfdFeg
qrlgyx3IwrIIdVF5dTsG27cOdlUTKXGRrA6a7m/DjrWywRF5F67cTCbkwlk5aCUO
X5E2ZQko+bbczN5gisdXjEeipCL5SYrcLivaGPPnrPu7iupINxPeIUzTWnUnGoji
mRPhLS6isSE5+5ddHyzeSdNIPrLryUnfv7uMArKgWfgF1gc0licaZTj4qNnwsYZc
F8ZNsgsxywE5Y/irW33RQEDJO4++D5LFkDSOSKPAR3YhQ4xbfN46+rdF2oSWvhjs
rf4Xpj9DLy0ZIywhm1ZC6dr5FnF5TYKOXH9ibRxec1Ov+Tb0YGnOXKI+1coy0lqc
JUYpV0ZS+0YpijbyNb+C5HN0b70SjxMd68LbpFQ0tWmuLG+FeqBLntKh8i22V2aD
R9vU7+c7umr5edk5NEFqxuX/QabjJdxTKzSBlmODfOOwdsfgkA1eGAmgskhdnc+e
G0DIBbGoIYy/3m6jOxYjwcgpHQ82jifcP5xsm9EaQvLvS5ifV01WZA3VcuYnPOz+
CPKFMDJXOmjqvCzTwQhlaHHvp6Ni1BrrY+Azz3DObS6FR9HEZcHuBMxFaz5cprlk
LZh05WuxjK6gVltnEMIc+NC9HrjylyysM0SsNeMv9LDHEkSvxmrt802Tx2e04iIR
y+vYJhBFumOzW7/hbgw6W8WFlZP7md8qb5wRWF3J0HIAS1+9qqd913nU2Q38FBjK
bNGr0l/vaHH+VyEbbeX9jUCwPQ9qeCGK4v42rBOelA+CvFAI63ePyXaizbOPheRT
LjXDw97n14XYIKqpKIk8N6azvPPQ3fagVA1kNBYW4R2qAoSWCsA9TRtOEKpRsBZ5
w3s24+S/piKdTWjnNUqaVXLNy9Dm6k90rKFBr8PQDH1WyX3c3NqN5CLqXLR98RKY
oOD4UB5w0bCWl6foz4BcmoMLeAdd+pDf4tRGGHAwwLkCaAJFKjRqYAz5mrFNMs+y
2WTiY98PkF7+1Jxx+eQsbo/G9/Dko8io5iVPC2LoIe7zHERLIEJv2gK1FyozUQoR
m350luL4I0J3BErmrrr5lzLDHigXkCiCgUgzvN5hgO3X5Bb0orCqiPruG5azfD6A
zxgTfxqEtezIMqJPnhaWu6a8D2wukmQIGkB5yoQJDnm3uHiyOW2XpXrugl3/vZTc
J17YLAn+CCXzRgrQH4dEfyIfllu8DUnwQozY+wdp0oQs/7mgiyVcOhceoLvBlI3P
ppg3COd4gCT9qNEB32xXbSFW4H73NfFE4aEtTum4BS/fZrUhpmkbFwqHmc4d+5Dk
cRfRoyuANF40MoRPPg8AMz13+gtH1MxcNFc23G/MxiKUqDH6MhHFqUL425Vg4/TR
KcxyhhANoI/TiTr2SGBzmFVmGWjU8MUsk1EhQA1OKSSng7RXZg0ArJyU+q5/GT3Y
ddIUJNz2HivsM8kRpA3LVcsjhkeAKPvth/VszPULdl+ImYdYNrmmH1MxVpe9Nj4h
bRtfOoDCPzYUeGQ3f2QMZGEBFE3evfssDSuypJOFGHug2Z7CuqI8xEuW4UxYCV1Y
ubbADN4FcTURB5t11allE4Xk3DC5L7U2NiHOyFDT/z0JvohUcGBGmSCugm2shZiD
+EPsddbA7+aCIZAOGPUaPukN4ks3EkdpET+TPwwB6FvHdk3FWgbriCzuAEHomZ5V
RpRKIQV+iHYH54Gmta5tBs3Ny4lVP+bqmQspLAR7lFngalISH9dZCH+MhnYc8OfL
viB6cboZikGesiQhR5CzYbi5pZlAbOBBxpqjeyHGX2shcUvd3gFcJRqw4r8KhKOJ
nUUadWnZ2V1x9wNldizriEAyE1DWIh96Xw8AXttb/W3jphZRCe8t3TxsXGwE9Ulb
pOGqX6lW5zfNTAGJxzXVdW/NCimTg9m3xOaxxo83Mx5LPIrzLhGMgqmawZeORxew
yMVwVU6PH4eaAY7L1/l2x804zEU+ynYfxTeMQvxMgM59B9NCkR0HSnGOW5nD/Xmf
HbBBy7kpZ2ro8H52/dZeYzV1JZcTYzs1rp3FEmHiFolKhp0Rltd5D4VDvc69Tuja
VJtZPccqR9dA+V8++0SX0t0QcMyO+kNPckTgtNwjyZxHgfSyZEuFE84XdXNB7Pyp
94SRL2yNABvDXhWekRL0WWPemvf04SkVAEZOuwNWJ+H0PIKSikWuRogvRl95dUkK
Z06qu28+8q4bSA3NQyqai6oe1LV4Pd11NgnZS4WNSRe1Ijbc3Lm8gIcthDTw46HP
FiH4Z2czcEDUgUxDUTuGbmd3otZcWZ6cXzMy+CMERmhJK4g7/dTxoELUqen4wrBe
HUrwXBjGgB7JVtKbzcrJYJiwWSEFQo9SXNlg2e63rvz6i+9sq1+zHQz8x0cLXY4I
57wT1aY4ydq+VmYa+sKxMfkzJ8YqBQZM7eVDlBbYru1gIkLygl9sh5NvL6kT0IyF
z+CjZ0+4/25+Z+b1YGXMi433nsRdK7ldgZHXO4z72k7wj0VQiIfagvRMWzd4IX40
rbLbZb2pSU12UR2SEq7SEzrtEY0lkJrjn9+LXu80lJEiXT4xiD+N6YWS+Hj2k9Vo
YlkXXOD5TPzFpWYOoD+n1Feri9bmozjNzaU0yaWStNv1o7nwYg7Vt+F+rj4tT+BR
Ywn5ZpoUbz/wVEz6GaPX8GJeQEjgIKEPyXHzr1HrDSy9jpgYmHeqxSkTdUNSwN04
N5HxkYCbKLV+j0tlUzr1PqkPNHFcVlDoQC6BvyuatMV9+zJYiFrBaci2qUCZg+cn
Mo6K5eV8EVA5F7iEormP0B8sOJmeRAJAXY3IxD6QzGCCgzFMEIa9ItYFTKqG9XTJ
YTqCLsvknN1lOfmjD6aN3hXAjp+dkPisjTkYrGVsXygCMmHaWs/V6uqVj0rab9ii
kKqE5kVDV2jtjbTjK37NIBG9hQp0+01erHeNOpKEcug6iUYjXbHJ0pqX6K79MBDE
ZcDepoh4Iq6SRu8Lk9dM/JmI6KD6eMDgiD1/eXomFMfwuf99dtzTxsNabf7me+IZ
wwMmAAttc9TkAIhiJUb2GlbmrHqpLHGcsjZZ65IIuk4rCz0Ne9/nhmI4PAe/wQ52
umimUu6iu0NUhkKVDy4rXikXM/ufETB5dng9+P6hF4RpuiB/ZSlF1+nePpRRm4el
NiNJtYNeqJQxdJzyEs74Pqugu+je4CGWZAOabKqh4BmU3k1qJW02kMUoqsJfXk/B
ZKxlgeXRfsfCuCyy3g/cLpE1tDInfcolP82l3523b7B5YGK98O6s5wSSMNXsveaF
0G+iAfcpMi924+mC/D4swaFlccMu+a3KqWbTjUtMxMgmb6/FLyknufQoiqgu+Y8N
kISNp09ajvKhmvee0S/ZvNfANQlEsFRDr1rRrKmfVWhoUQWFbE9q8mgadQYoC1cM
TrJbJTgDisdDDgTdtqMJR8rcc9pScXAWBlucmcHN2MwPmAnwMJvZigV8Xxurt2OP
9ArerxzIq1adnbj2Y0KzNt7LrSLYKS3e1bh8Rig9UccOkkEFpXpb2RRZBrXiTC9w
+CF6Qz6d75FOLPE/lGJ9jMK5DgNMwR3zInC9LqqwzJUdnQHMbMUcov+2FynleCf5
AIpu7V+cOd3j2YcUcgpYNouMPorgkiUMOqwJCEOLXp+fx4ZHGT9TfYTCfYOCdGtn
Lr6rq6hEAOvmtZuwGp2plmGRIz/NkV64eV2ZKlK6DgC1nu4IfpnS2YV4zYw3Ustp
1CkT+XXDLmM1nFoFnQCE4g==
`protect END_PROTECTED
