`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5MoJ4J3rv4ABhtcfpPGJETXMC1e39y0x0Hq3bTPMrvzu4Q79zSCFAdTfIdmmWGT
1x70KSz3i8dpS2IBetbAcc3gt+0x9wB6dNrEz79jw4dVQRcSt7NClX6dK9ETG/4A
MUE2P2g56iF1PiewqAo7nWTB4559zyJry/dHiLkA+9dgBvdN2CDkxJYfcR9ZxGw4
Jy7Zi9YMxUnH1uZwPZ2brO7/r3V6SfNprnx5RPKBe1sosJhAWBdNkMljz3HMv2Q1
J4Jfh95SFgSYKioRXHnlSpHJhk/MykBT30imuiZHDohV3pPAyuap7nn/P3m+8t8S
W8cCZxs5CiEXcsAwMdS3To0Sl+/sIMoWrkGcZk0aKyksz/Rs6wxGfLYnNJha+G92
RpCJ97P8WSVo8ASFkKVJmpCF1QKFtxp668gtbXirB3QFhu70xtQ/qtA89ro9fouI
WPdwXCGFWW+ZZF+RHtQ22eRv5oYKNeGofbCFAeHi3t2BDCSqlVNziJkAKsKPgl1j
pooVJ14kVnEWTbCK54WaOGayvlvqvHEXYjWdfXFs5fIxaxGL3HVsf3OCuB4eEmwa
dB3dPPJYG9sODBycflz9Ft/LtyzZrYVGaGUXsS8TASo38G+siPXWsQd86XjjTVjJ
BzZKXEkcVdCkO7DOJMJVqHPNCQ+C4HJOOwTUWd8gr/PUVEdODXbnAAxKZXPjYq6C
Te6wx80lBvwcNu5zo8mabUqcCSqF4H44KQwsfFft+XyuXSRO4shDzZNnjlSOqQWB
3vO+FfAtdHGChUXB6Jvj93nvppn6efg2c+U2LMwMpHFj1TdbZS94CrCvh5CQeBNZ
cScN85gBA+lVgDKye0CRxvVas60y0LCNUtk0jSbsclMIWdYs+2sxN3NzlbZjbyMb
odQ+WYQgg5BojVAIbETl4RDPSieK0bI5zi2ehC3Y3VPCGw6Ogb4CM7AX9vmZ9p7u
HlDmCIyLIYNVQNoa1NvrwTcRXj1VkOwle7Kg0OdIpWYna9CMfJGQSs7z3u/UAKeC
BvViOtRaH10Q6XEk7mI7Kztkm0PfXbTygNtzPeGppEJ3QB0GGX/XfjVzTGp1aaLU
wiLfi+2bPHrg7vM91yrTfDneO8VBK6vLR/qsVfXdFRiD1cyPrACh5/zBmOr/jm48
fYyopZpYviycMm5dGsO8abSLv4Igq0v9PN1WJkW75y2udHN4xCSbhR8JEQxHeTrr
uv3UsX5HT6wnj4nAxAcviV8skVys+9QLL+O3zIT6QxQTvjUbbrQ71zsecd2BWVZ0
cI/+w5gd/+yBFkZsPcMjwQv/SWIU2bhA/S8Q034YfFp4hymeq87YVCsomNeO700W
5JcHwqT1nVy/pGG0toHx1A5mlXphfCL6WJGoDiP3S/AaCniDY7+Gy3MlZbJtqIMu
rDinJSesoqpYXLl+NAK0+THVmeG7F+WJMm/kdT8x6bX6dPYBYZAn0EbDgZyCrNPU
KMNOI6/vfXGaenoIGuiffsvCB3Nne++1e1tSLI99oH3PRpNOEMAYFOgYtJhdrh0+
PBYUYH49Vm92rKGiQulCwegWdXe/4jEnlO4ZM9OYLAtlbSpZ2OpXy5xGy29GeKbS
i+2XtHVtLLe3EliMkGp9tJhmLEL3HdAFIn7cagprFOHR+xI9oCBXyUghKh5V+xar
HWbH2fmtEu48KMiFJT7zkp8mZLuh8twbn9pfLWalLZvnyNjSaa1oAewI432CbbAJ
qcjO/ClCLRBethW4GiruWFpLwEyaPik4Rg/ZE9SQjKQgYbXDKrVhk8rr3zEATTrz
ruUzLKzJCor9PA0kdKNHE+COx7/hebr1N8LYC3WJzuCRsFptbBlOZ1jlm2UFFEtT
CCNmjkQU4kNMpQFJp6PCbaZZA9z1xcteUwMfxr7hQV6lpyx8307jVWU3SoAd8gIv
h7wwAlGuXprYB/VN75eunbJ7kVzarW/cFdsKv63Do4AkfAoRd3PHHmqPZtCb8+nI
F+RUxXbCVwi5pBTv31tz+jykzNf5qhjENEXepvDmeh9oDEv1MVZH1aHQHNe0jv7P
l9VFyvlyzKr9fG0GjOZmcFmCc9bKDAv9SrODKPtyG5xpZTrtqXu8jzDX6iQfP45J
ROMhn/QGbPG/xT7aCUg6o6rG2jR5tv59Zsfkp8/o48WDPYKAdlVI9OlIdq/pykJs
itWibrhVzpYDxSgdg3C6qGeW4c93JuzEZ/HUHAKSxJV+moiXT9Sw7MJlMfqtPn+F
C6cWMn8gIKrY3BhsGd+iNQas8LomPUMndYAGVqbhw2N/383hTb8j1jXKIjv3Q9Zb
ki3XonNRj8iZXbK9oGLAuLd+IcBPI3w+KDWwQ/5d8+rY97ia2Oe4wwQ0mWHGAQRv
D+jNg/W7G9fr/I+/yIqO+lDbFyLapvEcY4oVI6QGRq2XF17QSKr3+YZfPe+S7v3Z
Pka36JIS2TiBpoKraX2rC9WDYOrpqe4nLGRJQRT6Ojv4S2UM/886NdA9/bcAw3w7
9tE8qruD6LPy9S5y1Zzn22p+NHC+zk5T73SvTQw7IwqtBxJkZQmWvJk4lpYyjBsJ
+cMm5kQLo07+zHT/gpD9zs4826YhWE1SBZVGhQ5zXYmmqezlPBytw+bg9x/jy6fT
LUuIe7mYVPPArAvU3kEdvjWoB9kzH8Wq2F2Dh4MjJYmc8sE58J7aWGqTzgTVSPui
xD8jS8qYDsYH3/ma3hI1+Nmd21r2gBaJZuVhbo8R4cGeg/dXYGIWeKEqbvetI1Da
3B80alQo17xcCL7QU4BX9+yBUpk2I1ZGTBCTw2NkppQsooThN4p9BEwojcO2D94r
mllt9xKI4jF6KMn2qeoQz1/yvrh6g4S2V9XiaKWLKfrTpWZl76XqN4E4kbpPrfKq
Gl4rr9a+ocg5WdCuHZysMkw/KK9PkavVWjdtCTW8xt2gd/BNcHPRlxU9Pm5wrIQ/
Hsco6G8dtEmehBLqD/ZokJ7yr+N9AWrjzhQwGV/nUzELsiuO4x8h9irxZ7XBZzep
zIJJPCjFe4FhFRgtqOi1jSn5d+qOF1TiYqLdn9j5VlG/dKNtZpB1hb0dbnzxWz4B
5QBtA+aaBcKac3HBXVHHnZUVO1FXf/7zvBWmElnEYIi01uC1/EUOGIZWzOqZELcM
v9cjvW3YVxEAQ9fQ9aPpMfoS24NIOUwUnWrT2Upo9Vf1K4FmzP75DeboLJk2kC2L
lyAyAzOoJrZUScXVaaq5Or20ObMvuJ37+gWfQoOxmo3K36ltr15Xye3/lyGmafem
vMpjhe2QhK5yn65Giujb3URLUBxkgWpEj1/Utv5k3kJeunVX6aMJywreLZQJaXmr
CHSZyiq9/OwzwCoOFmyZ6o28Xh6diu6koA+OA5yaswjrIvGK9xnBi7jv8w8WtESF
N56Xrte6JnyS/ZjBEVCNeRMbuhMrt2UfXL0FMDbSU+RSaRkAGYC2UvZQNcCGDipO
RYZvLflSl3tAYKLqnI8hRUTkiyosh5a24wnr13+EdlTMkilZG2upfg8B0mtN9Kbx
iGI+VKs8UqxRbAZT68t5/Is/2AhwwiyOCcbk6hMTr3rdFDZfgWjWEeHxisZJY8uf
mjZGF0SCK5/A/rZbShcyg4SbluqeGQJx+U63zcFbj79YZ6Br1s0BBaSbxVic2BAh
LILMltXGjpmkDTTRG1I54s4WEyLesXZGm3oG2OKwBIxHOnL3GhADwONOpKOBAv8D
CD0UenWZTwMupS+QNhxgfqM7hLec9m3AjfKsY5PTQEl7bs2K1XMDpMIYiAeCroxg
OAEchR2cuqn55v5MxXcU0xwzXBQLUhi9BMWnw3Uf3JxqJXVdLE7qCAn4ZDE+byJF
aKD12FaeEKwJ4rUieGpaq8MKWVJg1Fa80vLZ1D3j4Ja8KUsNailn5gGm0/hsS0qt
RhZihLcovK/cTA0EfIZGeXjihf+qQkB+N7PYStNMfEkQ0bETMp4V0qXZ7KQshSqX
ydZLdWJqBCdNF2YrEaKsV5IWAFgo3e9S028gdfEnK3blUCGX/JT9pDAEhzwG+cN8
JJPlnU/2TfVMuODwqQdNzxmNSHiVI349nVNcytprXkzrj1Zch5m123s0UHLU3y1W
tpnZjFwM1JI3yWFvwPchPYnyUFvVZBukISMgXBhMONNJj/7CSOpYRYN4pA7mY88x
9aTt7aVgxHLaQN6ojVP8NrY4+D8ZPxfFAE2VrazUfuC6GFutYPGHAPMa6Png+cFE
7vLGUnYDx/rBwnb7zvA/c8fnRwLSNm+WGSHNYCQXk1SdIQl8+ERR32Ks1uswE61h
p97nIaFroF8UiQ+uS2XvOCHHnkSue4Ycaz8UzM8U8CPyh3c20DzVDHKyr5dZkrsr
Qxdc8HRdDIpEPjhIYgSXHfvvA3+lOZ/ctpsESUfseWL8vPkznZeeXHCxwdCx2ACq
3c5objXku0UfkXTHQ8ur7dM9TOxTLdf5hctiMGz62OU3VYIoTltpS/RVJS0HcKkc
w9XLzEHyuPLSBtrhOAGEo23dMHt7pDUCif8WjDW+wzOMvIXvgKNf0QQZdy9mAjI7
MHKclqMhvdg88VwKMmWr+ANhmAxuz7JJxVlrzd4daM+WgbgoOzbiOpa91Eqwfaq2
H4UHbw8v+K/aMh0e7wnkhKS/AIJyYKPehjtPnIzLsE3yK22YKdFhOojzFansSTOK
DjuqbHyTmBcdyeGjDExpYfK6cP7uN+8oUMXfzNbK28dFqigLmoT7Qlq6Vx1bduK/
r5IgUXUUdHmFwqP7XLxoYWhXB3p+2B0YQYURp62zayeQXGmKWJuypbYiTjncP0ad
`protect END_PROTECTED
