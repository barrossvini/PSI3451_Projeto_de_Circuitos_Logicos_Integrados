`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MJgpePNcaEUAQCD8cpF5Qsu14di6UD4CGOxbduA0wqXKkni1SiRNPy/Ks5YAvP+L
dTj0LbBnc+EKfp7Ow1AH+QLZz/8atZ0Biyv6CfyKQoISsLz29B2k0KTKgTA+MUhg
oA35bsblUoucabX9oCW7jn95JsM67DVi0qPZWru0jr3381Thkwa3BqycnPqt8o5L
JftmTiHSRWYRdQ/hAGxVNYWRl41dTbQc7JVn1gJbSVYk7ScQ5umrjleV6rNzKPFF
JWKJC/cTaKYAVwDoznXvAoK+dh+TsC6eNJ982Y9lSk7ecaOdEEwjD4I88wUhmfN4
gwc8BoutZJuVZvUYMfAmt3EPgcidBt4aSKRjWGoCYjHcHm67c3kaEkH9Os3ANWg0
lAltVNXB+rnVPiQrio7/S2aXSknYegegeTbDCaX8ggyo6OXUo/DbyLtwq7cY63XW
mNQNPKVkpKEYvFqMNtZZf6+ZSIXE1EFK782laK2P/7+Gt9JtfJjm+6lr+PdVIlEX
dn7S2r9aXc5o/vhBOekg81fmG2WD4pA3U3UexJLFO2o89gUwhzZ2Ntkg5KI3RGW+
D1sZm6ID5JnPn23IQzYr3KV7+aCX2O8JPSxVmWc6CvkOCKYHx6+vp34Oih+xJo3K
cbWWM6dLWohdFvks2NK9Xn4SxhQJCwi+BXtsQ9BAKbzwMRnYmr7nG/XsOd7snc8k
m0q6u7r93lT1ibLb8y21Iq6KJmfWD1PXADjRYuOCNBMGRm3gY+SkrLmaQicVki6s
rUJlgt6WRcw4MI+ansOmoJECKa7d+Rn09N1U6a5f+VbjVxk16hjsm7vv5HtS2KUT
dXWHqfgVhYSwmEwt3nnxa3JKqgbsD8NiQoDN3gQNwWSJwgCqmUAKl+1NXf0YNjH9
me0mAo2s33+v/AbXI9FswwQQkd04bqRb4Cn0/Pm8Kc/Sf+9c22lkTYI3Irh5IwDY
awr7r3mUXkXZB7gJ2f9DsE0hW0Xfn8Vic6eFLpyUG6Ms+5M4RnqBUi7r3V/T8M4e
cB6dUWE3T56oYZDPIFw0DT24w/PoP7mjRkh+gGNsmuRvxl3LWf5KB0ri5SdJTtcN
SM7p/vZCw0L9en4XpMWDuUNL5/VToQjfS5qIDyFzGF5ujefZGUsPe2KBS+Q5GiVH
EPJsV6dWDupOc3ay6iMFh+Hd2K+RYB8AdHQPVXsuwGj0Jb0OxjS/EBv8yYybvbrW
FnA5JJigpnzZVC62w+F28qX8At2dGyda4CagppVPWRfyKIEUGr39bTwE+lujiEhI
RqE6zI9rD/4INTyElp7d3boSfaqLWHKn9KApqMcYgMx3/2WNcBQzaC/R7U541xlC
PkzAmi0Ds3o0yMH5095YQt5SBoSTdO9CnpJbOOz4XeNGtsz/T52Otl7Jmega0+J4
dKWYworhyoj+OnJvde1Gpii23aoZTxkhkDzGx4dAjoQX55VCRYcuJdRugyQaj04x
SW90Xxh3h8ajb+6SoHf5OvOr9mujIqVuaauNB0gbnzeYbUyHC2lNChTszgH4J8/G
XjV4OtimUmTlf2w5rNFzCtXxZq/U2NRidqt7sKSf80aG05Tos6wxDu9+xOecXkOD
tq67GR248sMYabYq2zlO63xFqsDnKlHXZorpc2BRLS7P638P8Zq9bzRXbnq4HxM1
UsEaux6XJ7VBIB8Noo/0mnBQL/gaZsgrE58SLLpZNHGEvybJX9wjs2hlVqFKUrJw
ER+5b02Sru8kIrN7zuNaRDHIqLLJto0AFxhRO2TyX1qxX+QfuI2JINHhgNx7slVF
NcbXhS6/ACOLomIZmUgCnc1PmQPiWtAdzwohPrj4sr/5jUz2okT3mTbOc6RwPrZO
6jhIdhOGd8/yn4YUfIzAx9Vj2F/6X6zy6sH0XiGOv+Koi/6XtNe9ooZkNr7Y4NRu
qVG1BBo9KlezTIiokLWnAXqDl6CPuoPumtV1yu9cViJraEtp6440PiF0WvynDcFt
GpbA9VnEdQ5ffbteFiOujmhxNZPFlHEpgEMw5kPFj4dAKv4xB6c6lDNCpQFo2hRw
uWHWl2qNMsfQ+0+TrO3qM1Z4CWE3iMm5FHk+YokNwlWuesSJx5cCfWpkPX2WnvtQ
IPPDKq2lcPgGac78xxY3hZlalhi9d+4TsFZIgY3cHW7EcrOk7Lc8TjmPk17BvaiG
vohyGIeNUV4eJt93Uffk68QEDCOU5mLkpwXofAdc5A+sd0HlIU32R1XiQyeHJJm0
DL0ZxBpzPeGC86GkCVIBc+FGZgRFbHSUZJuB1CeAGNOoiuAwrr3neCDo52ItPd+T
x4SOPkFQtlnnyi2aDxbj9rHxSLACR1AroY9AYPPbg1/0fAmPYl3qd1ve7hehGNNP
u23IerObKDVB421rCsB1ca/OGFEkgDBSblXm9fk+5E6uZhbRlh9CaBXh+uYasSYX
AIwpIiXSjfeovvBz/JxxRLldqnbEfILuE8U0NM34LKctewzXZb58m6rrCBAl/+AZ
MwTc7u3xAlHvF214VjuDrk06arcjk7PZ/bQkPiiXvjL/kxEgf1fq9EjZk61LYtDA
Dio5heS4MtZaSWJysrRK9qsmpD1p2r8kL3V1M38l95LGUerC6CzQK7+G+bYxx6Vx
/FJ0TBPbU5t8BXBAxwqtII9Izc9RW4brAfLx20gu2YysOHFQR8mWhwM2Gsr6vinV
uIF+C70zZn0zQKNvshpuno8kO4O8Vd0DP8hX5EzQtj8Rxpq7CWNFz39haSFb3SwC
IbvjXas5fPDzS/zIusezSl0ajI+ez/zI+Bxa0gfIch2gSNtgkKvZxa1fZqVXXPG/
GuGy7lSaxMmUdb7yH2UAMU6xP/8+D/Y+TEpllQ3y5eaHmWLzGfca1zaIavuoS4eq
IkKo8gK3dTa9DYO0YuKZIiigsTe+Pm37RCa0YuzY/3k3ciMqS99om6ExbcVzYSU5
34asLhe1/IpVvz9ADPuYnQsXVv+Fw7HoCB7nW7nsjSWF2u1vd5xnqgpbIF7JiX39
vydisp4UOSqQb9RPHs204U9q53MwvyW8cUMSasrMJFbdu4ompLH7z5PRjOwK2JjM
4/VDKSVNTo7YngGFVof905elcPd8Wthbui1DdFeh/AhjYxAfkMjjYC2zU+3Ws1NJ
Fnc84p/fUIqQXyyUpjRr5xHZcGaO/GfohOuoe9WJZF70fkDColh5WnVEAixdTX6l
MUo9u1LBovyxeW+oeWn5NY4Zq6yTDS9CMxSw05piVZqKLqKj2bPThfLjZnnWFlFO
HTwRiOWhClrbRQTgGo3jyN3Mh1z6UooDbserlSnmelGgIKEXgP4wkmw6oDdX+hF6
RIb2M+P8tb/z7mPIHnZclD+KOD7U+s1dU0UrFaIeklUXia9LG5u5JmTkqDcRGc9s
ozEuPzAHHMngvYx9raoalSadXx6/ySNXJhBNhEo2DBiE10AcM280TFjOVNpF4UgW
8RVqFmMgqRNKBqXAXSH/ekZuX7RqeUNpk8TEBmpF6w5upscnZmyjKIPzFWiqAug1
XTnqknnVFZU2soi3SUvwxFMvGjnc4pZimX59g/I1APhPZhXIBkoNT2SBLeIVrQ4o
UD3V/1MrhzRsXmb+QuIVcQ4Y2mOLnwAlm7B9GXinPVAJpw8wTa3QR1rw1cyFTy7x
lGGuHriukYOmv/NwDhPQPQFNzlpq5t1SrOBniNdAfunAYjWiQko097m7+l5rKXcp
WoR38paJFkJWLJVdvpGCL2TcHKDi8SIiPqYfHxGCQDjHgNnzlxLaXYWpu9vXWF+t
2YNvatGJPt4DOCsV7otSVAhRU6LGQlMGkWEvohyZiVf6OjhzdfPTGBC78OLlquWt
9zODBeqvnk++NWmWLI7iNGKSg3kqOOpdJjRGy/WNN1WtjGrwoVIoU5co5YRqHCr+
DtOlSI+LhC/b2o3mPDE3MN4h/3g/5jtrjYHWQ6eCZU1F9kTOrvhcshB9d56XGDio
DjWqN0ZdjI3tq/w9HUexy3zu3H0tpR2LE73Rbfm0P7Brs/YFQzh8Urs3stVUyO60
+GNp1OMMxOJORlBA87UQgOzj7nDuqEb1tQ5WdDGMNmEoS+/cV4Al2/O4cSBXI+5S
Hrb9dBjCpc0qyxurav7ZAtbo7N3OM+yP4ZJqcCjJYhw2Eihfai8Y4X5FgK5Zt14j
QW4EXXr/tRUcM7EUss0YaRbFjpEdes2d3iyPQR7vUR2L6wbsR4vU97k/VTRPOiWB
M80WeKqLeU/nju5bTFE6FwPAh+ZdhVAskFxLDRSwGBlQhFWu9e3NrORTyfr7Mtp7
SOGgSEmXxKShH4ZWqpfiA1PRHiOdbLrED389Ab/PhyU3fHVMbFz86tEf3QAo6aOR
Rt+7PH19Gm1U03a5QILEoudcE+E+ORo++IwJtZG8O2x5eaQZvJmWv7JpC6cOCo7v
tWW9Vk/1PKfJkWuMXHjN0sjeyY6L6Wd/Sht2+DjiRfHxqOSh4rRZRGs7S1ypFdKM
YhOHLV9UKAfd00CDkj7rW0UdcaQBX4F3mNV9sIS3iHJNjlBYphLBQjAsvxTMx4++
wOaCKCHmBRMPsKNISys8TejWgodw78Mofu5iHSMfM3qqeD/bXAhY1Tzsv8VydtBD
Lx4agoxzufcXf0aZdW9WGpfGaAcZRpoubk5a35VsJs/z1Esd/qdfua8f+doP6ab0
DrIYt5Bl8y8ejFx5lJAD68/iFfYq3GevO4oavDqt0ljaFRJjGj3aAWOg+KnnwO7V
nmFKFefdKmhN190bTt1NsZ+tfW2uT98ymGBVSBRYQN857HtUvQZni/p1mvujCIfJ
ZXi5AeCcMtgpXiU7oFeQIo1hVLsiAJRvhPNLwat8QpemileEvKFEj7beL+OWSzMr
9iLYb04pmthbNaDeaGcQAeUFOqPkuCgqOqeI0PRmzZIIW5MC6TKkM/uTr4csDQtJ
ptQ8HpZ2Fp8iblqXLvNoEZ5OIHF+r4My9VlVbepMTL6AYyNGGbAh6EbEpjwc1S+e
8lwOB2AZF8xxKdJTxRKRsDKv+7paB1cKKLQoXoYExPZk72AOjsnDOoalOhT9PA6U
lSmQ9p2vpcYA/w75iONUZakgWa01Cz8k/L+Ffz498BRrH8wP5g2R2QwPGZSbd/Ub
KikTQiYy6Q+BBpxTt3YMVcbNVN0wftsXC4uGEDtC8GKyjRCGdA1e00PQmhmNc4TX
D74oUyDfeSVvXRHfFEM5wpQVshSfLcYeqOO5+CF3Y9QTCSFjFuYHILuqX9v58m2P
HGdHbBBiuCTLigGXhPquOJhgQQjkA1NQGIHn+0Z3de2ZXMnndUmn2e6VtJeQ9uzr
hL8tnwP1Zreg6l21gcDFLXQXXP3ltQ3ys8o3H2+6K7N78kDFiEsjalaGT/CGFplt
yXpyeelp0iGUYcz2U5XiEnqEQn0bTIZKmVCCYuhSQSRZAZvtd+qbkrenzJ263As1
BCOVQxC315oTOjNbgaEj8vAoWAn4OMATkcn9R/qHX18sLx7/D5Jz2AcW5ZZwrX+j
V4lMgNrxYrOZ9myb3Elr3ok/UaL1WInFMVyFiFNmxLtvAJBdplPlJsne02T4Kj+S
5NLddt0knv3xcLi9SKDCo9OfhKluITqLeR0LtGGa7SXIjIkbOWdZ8cPJBHv5zSyS
M2W250BMS5JdHY4ueq+zN0m4Njk9/6M28Bw9OR2uNBf7i+rBHYli8BUyW6Ywky/x
sC152Ts80Igkz3J9Y4THvQC2cQp3rqW02dpy6zVQz0li4/OR8PGQDgZyJvrgChlA
j+bpO9QkwVMyHa/j6Ocny1G8zhRvptYaVBd7jd2T1dqzMIANTtT7SW7UabDUYTBC
O8F7dWGC7AENWw+ka5udm9uNvdcb45hZActziVqJFTYeFjgUwM9NffaxeEoMizdn
yr404VEGAzlFfNMNlbuJDsma+LyLRGB1WsDYOLAquwbirGWNDJgty7pwkWjvqqDA
kQmgD925bN/U8KMNLgF+1m5ZY7KSOB0jcqZXhCwdl0zRTrcBYqOcyJetwEMLaSpA
zMelm2yoqD+24SLRcr26sJ5D1Gop7/USQFGprzoEEtWslB6OGmnnKu1t3Ws3Zupo
M9W0ebqJG8tKZcjk52iuarS6FYIMF1KItxGcfvdmw0nydFSype/6AEyYUI8QHn6O
8OwilKVw14Z3rKcHkie2mUFA+8EuLrUp2EDNxsaiIX2bpGsZ6t6y/SoclHAVjBbp
KN50OgFx288vo8km1EErZC3stQ8ks5NzJfxQXBWm629Dl6tOYj9ueL7ASF3mG5xb
rrVyDPx0AlDEJctWyLAFcdLULvHi5Dqx6jOWyYJbbWTHC1AhFhvEyULhipLqd+s2
TyQrUHazfJZZzvw0vK5rdyW2i5N9WH9r8C7EZ8edHmXZVZtkcWQYu/eZcb3A3xqb
WxfuJWPC0bwaC0gyv+sXAxfIUoaGpcYtvvSUTcIFg4+88aS/UhHVAfhm0DquJv6W
sq6ZvI65kXYx9txzuJpJAB6Kbj0Tc4xEtoepb9EyDuqsAzRHUp7sI6A3IknrgfcH
2sbOIXlsJn016lFGHIu2/8foCHaQihIyi9SLCrERH0BR7czfFituDRi9fR9hh9mj
/kehG7io4MSm3UJfFG2FrYxdyi6xNm/na2HR8H00EisUyZl56HH+8zieTN6RfnWw
/0Il0pDVhdzQjZxZQ7BL/34QM/3j4DBk2cnWNBiaplXUJ/pp4q5HNH0cs94V0LUk
3CMkXUo27NO14VAFWy+AwcsruMeD6cvfSoGy1m/oY86SSq4+LkIx61n6P9IsHYyh
LDGME7Y0f0Whxb/VfROF5Z8dmQfh1kSpn47t75NF6nJ+LF4tW6euk2xStbk3xBSm
xyS8rsLbTzSf9wksP6sLlwMJfNc3oXuvelOOxwViOrCfYzmSMHaLm9vGPfSoa62b
9mrSaEMukUEGUgwOl/+vQ1yFaVRT3uEjgHGIIfrzzP+BGgZTIcyoQgmVxyGVhSmT
dNuYn8sdY1qUre29FKKqr4iRsyYKSjIH/95LAMc1DoNEJB1B46ORpwi7fMPmbDlr
0IgZHWJUc1lf7B12lOqJN2w1ESwNU5Aq6K555xqgmLSZTkXguFdYIYe4kyPYG4I7
WSjtcmI0dZ6gVzzz0a4eFEeXGLz4m856SIaMbIS+Fx8vDyIHCON2T/8hJf1ShkEj
zKnCeIMsC4rWkTy6BIWUIpy6HuL20lKIedrTxmvVBE4ONQQIJoxjasGs5IqVkSpS
08vXzoNp8UFFGwMn6u2uNEqLYH3D/7KulEHv6LBtojZ3vEHZzJ7IjfYY1PpPNvSj
oclV6XcpbSMirEU4xPO2Q8AER9SQVlmivUzIn1MGtAug+k/OFsm7L9cdIPVr+R6E
LJ+d8RePMaFqEwl1J+EipjYJPkanbAMUv/JlCL4Xe5AMy3G+ryd5lLDGZ7VP9v+G
eOoyP/oIHDa4s6np5OT0MCDKvEAVY8z0OgLTPuPGffh1mcKXTKO304rnjcRMvhJO
ELiGiEnrIDpN+WdRJVcWFYppxQqtuKkID3/2FyKb7Gc2ZC+NoFB9Bdf8eB91QLAG
vw/PGytAx26THsaz6Nl0LIwSiBlRyfMBNpNDPUIQwBP8m+Wf7Zqf7OMixvwM5Hjb
SBqC2cg3c9KZg/cKPadEolST3/4oNetSgdA80aTlHWlKjEf3CwbXKH7A2eq7DsSD
oCz+Ke479lFHiaseaUssbuInp5wOKWNxce5IeNZtgRcVLxbKWba+p7ofRxlwFc5O
5KcmUKJM8BPevegS1m1embfnzioK1kjFBYps6JsEZeBN4ompWJmH+6EhabtPs3Ty
FIBOn9zwOmnwqYyLsdIUE5SJ7hMtNqLuT/ZMzTBSvUV4qZoBxFLe22OzqR1HsOOE
JmpzU4rAq6MPzG7XxPxxNJbIJeoEpz+jhCfyLau2CR4xNQrKNJGb6f6UGRfD0vX6
TfBgyAFboLaAOYYl7mLcsabqhMO2BWXjeOyzxPVpBsuF7rdH5eqI7mHW+8Y8Sdag
pfRlnlPBGK0Y/YmiHzQ6j3iMNFJ4pdzCMmLsRPGwL6ozcBakC5UV/zvViGwwN9ME
DdcmKO9sAhV3KgjDd4z3+zPuUE+lkb0pd9KME2El08+8tkr7XnCmPe+DZ1j14AKS
9FCfeXAAd1sGd0XUzzLbXCZqge89JvgeEq1QMfo8Kv+Kv2AADjrB2ovZ0tTT6mdz
Sispa0CHPN2Jrpat0pRq7FhSbDtBncoagnMImUF+VOaAnU2Ov/OaWC1TWvjjGjws
AK0KJ7pY2qF+9ePE3XwhfdJgUwTOyXI5WXY4sjVZNbkWGOh0gAZiT0Qa9kLPuIdR
UgyBwVvLLfj2ubvt4brrT6TdEK8mrnnD78Nj1kGa47lHPHho8IwyTfqR4i0QUI7D
rfAdh0i1X+EFo/KPbjazcxXNd7tVvZmUfYbRud6sKFtWY36gefz4l8+oIry8USOy
9mdK5ikPoLq6DQh+S+Bnsl25FJgVVON5/LgnGdt1NxjhqWQcMOmOAKJNbsa3IrKG
26WEYqv1YJBWCn2RGxXHyr64LAfSS6fWp7sZkHI9HBn+dmq8TU66RyW95zkySpXl
HrKuvHSHG37+hWyCIYwynUSeE4LgZdJ1nQ6t1R3nQFFb62HNwT1zxcMxziEhd5vJ
oICMeohW5MNFrSK3hbMQ2gOPOCbt1HrZ0DHYE5kOdDDgdU2qbS6evJVgEhW8MtzH
xBiLU7iteGCSVCrsTa8u1e1wvOIjqpaC0v97ltoMAYbOcTzC9OvfMJu1rQQKScbZ
CaCKNGs7KFCH7mX8/ztsFKisOvaNQ41RL+lmAhJVLpezPjEROMlbl3eckOVb7Gi0
Zaz/1oK2nVZROromZe7ELEdQCIFgP0yilu0y2AcFuFTkEQaPSrpUozX7hFhqxTbe
mR42gyRH4XI1iwqwMkvylmx6ha7UFaA1NxcQAuohyvfEf9BDlLiOytTCDq12BE7p
ffMewXZzUnAqjQ1x/wiZKNFAVemU8gQ5Ukh0EApOLjeOsF4eCbhrg8QQUvMtzw5o
NHyD/yq5fzRUOxzi1JdG63hl1hsZqnXAS5rK2QICH5TfwxmlnSip/Q+E1SHklV6u
MzldYHsZkckjI/TALHaSsSQJ13Xb2/9rRp61o2E62gc+kHwxsw/mMWr3WHzm1qHD
nHg/O2jeo+qizeSV4w98DLKnomiZzNY7l4C5bdX7kEPzNXlEvO5Pd6oyyWPuQDGb
Wd5W/eBImqhapqbNYnmo+vf7YW3QACaSI3kcnuXJOV/aGY7DAB061SM9Z74sbe6c
zOUGLcabB73OGP+3e7d1UCQqSa8r/5sVQbPumD8Zm+53ni2f5A0P/yJY+vXcwvay
fcCfwbnSa2juWP7GPH+McFDLqQ/J+RDzBLu30JtyOu8relP+acT42ATUGMdcBRYZ
leFr5vuCtavkz4axK3CUv5XCKR9GgQEhPN2LqC45XxE7TYuoV6VzvR5OmoNzph5k
KQ5zsJsAGnB7S5qDOeNygDZ7ezxcLoGTbOCRh9Cck7pS240oiuMfYosUJ+9nAR85
qS3oWYtkI2PSRdaQTTWHboeEMarQ75RnC6XFFSDMymQCyDXkbmMaACfb1OtjV7BB
d0mIkGx65Ll/KpLJYNeoQRwTWv28G45DdlR+UGp4W66IxlI0Yn+d2jserKg3l9PH
UPcxfllWeGlF5nEnaMI6ZNYJsX33JvQe7/ikJb0PTDNn3B4lFVf0g744d68ULxoG
2+dAdeElPryS+j82jYu9SpfxLhp8Wi5yzL2SMktwKodV64ExgkJyYUJuX8C+F6Vy
0C/9kYOPZoEEKV9IJ6YY//nCNLH5bAMzczE47ri74rXur/9vz7hTcWOni5uKEU8l
E9DfuAk3F7h2rPWVhhyC3oN4PAl2u2O/ritxm2WGFo5BmsNZlfB5jpFirelp9xmd
XHq5Njiu74Fc2Vy/2gWsyRRSbjmwiLgLhloWGZChn2b+8A1f+nUXTdodYSxZGNF8
4ggu0hf/AENYWSLgq2SEUV5dENBJDJPzqJKtxpXbUgKT8l+9Bbd39C5prLwe1/uO
q3Xm9cYQx6LA6IQz7/YEUw14UQiT8IXLGkrX7SS6uZTcGD61mesKU5MfGFmwNN1U
BKcMPyUk9t640mFLU3wi7T43rkJF3GAM8V4Uj+47oMIGNBz5rODu2CFm17o5JNGM
kwfWynRDEJIFCm8H8B48jrCT9nG8sfbwgE1jLASNZwneScM6pDuJQtNn085xJQeM
myHQ7EkjAIFDCtBgz2JjiTYIZ6yBEtrEaZAvUORQJWAhRhScildN//EzB3E3Mn8b
J7lwciTiT1k1vLn4Ljc+O3kRMUDNgymnzo2Mf5PJJQ0/TfTNvspJaRVE/VZ1QrA/
3UY4Uj/HMZJnYxQL9KWp5WD0OF9MKDB57FTul+VLoWhdVLnncd86lW6ZNFksdfEA
iXXOEsqY0Z0Fa+dOtYAb+ubJ7MHAOv3KFOolArXMVosU3wK43bKyieFOG6baxU3p
4GihLKHAyNtznHkn4hUAMiZl7qfCPJO2KollWf1IsrCV5iW60meyBPjvrcAHYXWg
AiC/umg9/LMdyaiUaKs6TTvxiM9zAsOAi16Jn02gS9NkhQJcOyfi9Ua8ZfRhkMWx
BI/70oWTaT04xFPs0soSsLt6ClwtuCZIkSC5AUIRGlwOYe0Av4o2RQ8DKNDAil7e
0q3tb4n2akFK1MLRlaS4c31aYpb5xlHp4G/2LiveWKstISEeZmAG1FGN8nZ3ljGC
SGojCqxOaLaflDrwFfCUOF6rb/VLd6ZvuFscXaVbArcR8GQ9f3ddxB5ONImodrJx
/uncUCY8sVrtghOUw39jdjrUxJnArZba95e5wZ07xRKKq6iD+fkihOb7J/P6M8S0
ZQ2wcrzxXVDT2PCONT16tFu+xHg7fDnhP3ukmGeIhfndNbF529786L608xtXMSPT
M4jmRs1Y9aUL/wQJnDegP8FZmKKqjcJ0WwcwNtQ1yi8mUw6OL1HSN/Q9Zxotstv4
/W2jv8ZaR4pcuggJEKNOGysoSGoXkDWwWaCCBNYDLSLOxtabWGcET4gLg93sLWKR
AeH875TjFoH9MwK0XQ1h8siihE9eGJe7cWZ1wxnjYZFzWZg3FD40oPu3tfAzxMq2
4OIcuQ1/aoT70Empw/b5+jECjrqKRhjolA8Vk1Kv4fvgPo3uS4UFiHD2zAS8dk+F
aQ5AlBeBmXKklVZ2AvHquGEnk6tWr1rcaQChzPFpai0vIVJRQRwdQcwVyOEFklUM
8IOvuNKzQhSdmIHjW7V/IobnjjlZYfn3y//gyT24e3kVIAqQMpDYcElSkWE3MaYG
egp4M/G8vkgq0v44wjMEtNRUdRFlbZqI4j+iPrlerrlZNUBhuUDXz/rjFxNpM6Zy
DUvTYX13+U/dbwIPa9+ScqsaObcekCL5v7qpoT2Y/E5B24spxM2PmOOD8NcxeDcp
axl0n4+21BXvHTXQ4DgHZcCAMkrNm/G0Xr56GIsX5J1dFDj6BbdDJ2aN5pdsmUpj
Wf+VeBo7aL+Yc7S3qD39BXjwy+IE10yfhgT390fI/QP34mK0S7lk/h9PMInBcQL4
pJrPrlc44jCVyAHmtGg3LQuv+ZITNxg2RPhlRXfMPWpKn5KypQd8JDrrpkSfhhMb
78fvhGJPUcNgIaB/iqe00bSlm/wA0sKs6ZzVNhOCP1guWmFxnLfU3L1A4JBz6pTf
Srg7aGtXivgAdd+KeAx766k8EcRjzhJK7WhhDK69mXq9bYbhAxIC/mkZ4zLVWW3J
E3DojlFzKsJCaM9WCkJeKdPybL8C+yj7fEZ1iZcuUfE8NnhDtUFGeawYfcoAYi82
lfa3CflaFa9P9UGhMqDYEhyS/2dHUj4R06kSf+E2g1Qu09lO0lMoz0kC9j0Moeix
XxM9eltYnyjX5RGIrAU0ECUI2rwM2P05egxDcwTqEPssAHx6++9DYplQKlA96QhM
nlNaROFjkrxkSXWTOn3vVYJMk8Vrv41W5pWk/vVq7aoJoYbBWPxKL+gLXFBjSlYb
S6MAKO5xlUKRUoYkGuivOs9Iu0vQeiLiw+jb9Ojlc+5kmQJtjRGdQKKxKIhBzwbh
GLDUnm2/MWl2cW67bcyB5HLp5CivbQwMy+BMhQUv+/eJz8hnurctjEC9HmnTrQaS
9YFhfUOWzVaQOJIZB4A3EMYRaWsNqdTaT6LZKT13UVl5aarQDBdCZWsMIksqxAwa
FcbLvC52M9JdgLCCAxi8+AX2MQWmOEX69YDNzMSgapd4+BWGDlCgovu4SQtXM8NF
5CDJDepWXDfLrkGRT56zlyZzIp3LFeQ77gomzamiLJIMFES/Y00hZIaKHiNhge2t
aVwtF9QScj2AohfFzTIRIO+d7W8NeulDYiMQNBO9DFC7OEX65lOa09Ti1v1NSakN
bauhFRR5n6rIYE1hIpoTttmJ+lP2EaXEMisimhMVmLQBoElAs82FGF8aHSd06jhC
fpUcQ7OLT3IIdYQa8yZYZNeoGxgwAbbfzoIOagyNO/w=
`protect END_PROTECTED
