`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Ai+3fRS73Hv6SXbxdgNj+jkz+vpCllSAgpkHNJYTseDl4ylWZdLnjf7PMA6nrRd
Lo8zyAzhqZpR3xbDgQuy6y2qxTm0AfbQ0mZldcXPvo9Aa4HTMePvVvHQI5YpD0B7
ZHAlPWMFCxcUdV85c3k1squVv/mBu46Di13cYs4e95kuGZe/zqCWiF39SnmhOd4v
+J7Z8HGT/EkxYDS6epqHggE4jM2GR7LY9XOhyeEqNq7UHgeAifNLRLMaSqC0+AfJ
rkJXG4azgecPtEeJ+z7S3ekSNnCn/jiTTt41zGo60wIbw/hSOERjnnwDMDiBqy3Z
G66BQ4z0yN8XSJUfgAMLx/qqkBBGzlxOG7BiXooloS3lwYUnyeCmw2y/caqcA3qX
4I1cnmFdPVLAFdAuiUo/DviWleOvktrTTRm5Wfn76qhEyR5kcTK4kfbjW9BL6L8M
4m13GLPgGVQc58Ni39bzLdGXbeoWSUJbGUYgHMPEDetEAa4sDOImNvbOpQCZ7Wxd
pHFP/uo1H4/UyDeoMYqeQ2IoJStOf7rY2kI2Ho5tSxOdOPBrAah8RZvRaYRl6Xta
tlmg5GTqnSo85VHHo1m+1BchUIGFV5TRy3z+VblqaCCs+FyLtYz46i3/0snJA3dG
8nGf1d+GzbZvgNE5EpfJN8etKx3Pgm2NrJUrTwoHDV72hf1kHPbMEnfrW15bB9XF
S1qowfBU7GfiLlVtadyf38sBeqtNQEZGW0cgEfFPHgYBVIldmktaZQdGFlsKbe3M
tJNGDUIeeINQHecobWnV9vKhIJDV9dUIZpRfvYeHVUSpZGl/uM5ijTl7JROTulrC
FEwjD+/3B3VBNEcKXJuAW5ArRjuPGEh/aJF2PXg8CFCveRmQYsV3Biqw4bCRhm2o
EaqhnDCcnEsblY3b6ooJGBMHNWcFv/Rg2C+Kg4ymOEARYSiUu+pP+909tCj0BX7B
tYeA1JblpCRydfQxWaZXrGoDrEZ8iuVuGVLL2Og/yUkRorLSh6lv3x9Jn2gi+zXU
6iOAPfnfo7W0zciWWYCiR85YGa1qygoc6nSKfq3qHPGZp1tH1unQhL09XK94wjwp
CRys7X/gUql5IN5iiMcN3kYNh8r+N5dBgZqvwtOT/lHC9YUl/ConJoSsab8/qkHR
uZdQ3Lfj7voFCIe5xkzVnGTJyPxpBCkAJZDk11qzCXarNVJJT+ZYNqUXZUtAdvsp
B1tpDr+6hLx2p+EOw5HNd/xiPBzCAjnHvveNyKwf87gJvf6XxjiSxxnIV1HWos8+
PT1SWrQ5ufq+MqnZUoR7T1sIsWJerp0JK2sqFpb3JFwD21YkmVtiIk252buFtDzC
2htzTd+fubyD64Zhoe0RAVJz9jfsFjU1ELWg4bDfOZB2SjwkctCS/ufPw7vQVEcf
xESdkq2wBtQ0/TU3/4urzmqPJcWFuf2SPRntnMeoD+pXTQJhmXkQ8sD6ab0HjXY6
OV3WL3ePiZmcSKZw3m4v6FTnrGHPV8STF1hdgMpdJeSKWqQKSAuMmUTqTQhylSL0
0iS0u3QlM2U2bS8uqYdldSBBlKZvQNT+dPPUcYVeTQSuVPEfDVe7kb5uvBaOCz2f
Fe0yO3oUMRV+dFTJsavSwtHrInK5CEzyhuyHZBC0pHUnKVPPeMiRTRTptJxMAbui
U+Z5/2HCvsaZxh6+26gcIpJdkE7Fgss6c21zIGGfh1hUgPJv4NdXKAlY6i2b8IvB
StFOBHZpQRF9E3oXgMV8ALGW22cKJkd2Z/t8MuNlL/MgH/ANzU/6LQKaIbX0OujJ
3X0DkZfBzutRcjcSJ2K1gtYDsgBqH1SB9/6QwwoSxi3DOdMjvBa8Ru4ljPoGwzpZ
cNtHnaLtEh+4HYYEDAiWCw3sVTbhOAh9kS7pBRi/rReb3f8JCg/g5F80bUnUIoQu
VlgFhvKbBr3Mk8d7Lsyym76u+H68+pujlOfNR5X2u+z1p1G+yjbQLj+OqSuqwruD
E1OT/2xNmqECGwmLN9Fqn3B78TmN0kG0UhQ7FGeN9KS1IODPsjak03Vu9NHcllzU
IZqoNdApWvsS52IhYX6cZAHimucg69x/hwqPBMVIvfPoAwtyoXPl6bxHCmbeiM4O
E4QO/6iIZGvP/UESVM/cUF/UWuJBsorjtY6H0CJhck3gqsasH2jU0mEAKQOVP7RE
Tzyc8/KzY+dvl4vPrDf8Kp3CV8bqwarmSXvff7Yi5284Q1ahLgfuhUKM+2dzlNwG
OZoQ1toKZBpSYiRFppV+UDXUZ1rvdCDjBvl9HI2ArLU1mekderc/SgbSFffroRcR
op+SPeW+0bBiVZ0BkyVPf2V4J+rxPH06UBk/MjZUlA04Q1et2srIzaZeREb+T6P/
a3xMUEHHCa9a3+pfoGTE5nFUen89a+ZEceVycrtW6OZ4U+6eKbEQ2vTZx4x+V0D+
82NG5JKKwON0+TrUZFLZrnZu2WlID5sDqOjZnsgoDq5VAnjveAzE3GZTmVJPyOdp
op7viE9au3/dB2G6WiKDmROkyV0CegezYEMmHhty36eGG7NdoDnRAKMZ1U7VrRuN
TZzgdQ9dYQlfh5vyqDLIQMjmT08k5j3rORwBHuI4EBmcvhZ5Gl+lmExohcF8yq2X
nS3cziFBkGeURAvLiNvSg6DcQ8qj1MlbvKEVRi3kksrnI4/58Y2pMZesvt9mcx0k
iy6+ivogZkUuq8YTDdNZ0ehgJWgWBXvvwpzufVErCCzyEXYAObhfrZStEh8EmcSb
rLq6ERyNWZTmT91JQLPaLlsOU/sAizD46TXn5aeF/7GbR3x1MARY8VnCHzX8WAu7
6DWP1necrzC5iYbGTeiALdHU20gdjkwj8LT1UrSOH0T8bU+rxdF63OX5i4poAMF0
iX5/GfuzBBSQjyx8VEXLV3RmCdIcGBGNIpZ7+Xcz4wFhrRht+teWW9zfSCTbCmXt
X/w+7C4KB4mRJkHjnszPqkAknn/fLvX//lEMsrQ94JfR4XURqhyBWS2xkbCVYCTm
98NKbiBbhlbi4WdPFEjyVTEtc2x7sZmlq2pLwOyQzbtk2E5P0XyDi3sm8ut7oZl6
m6OR6y99Ifo4nc3SsMuO9MqFerSQo0g0jcJkYz6MQjJTjUa+YwatC71exepMh0L/
gNj+N0dOYqRHzaiD74ezPvE9Y0pmVV908s+8FsFuudi3NLe1yAEwvq8C6iMwryMp
OnYNYctC+Z/1VlHWn5sselZIeF8EPO9ifkSbpTqYyckdTulLRvQhd4oNFGcG8Jsc
MzLEwN/95U5vITN6UEbe3IkA7EHeTuOikbs86myH44bbp+ZenOIqodwtHMI/2015
JVAdT2Tf8rAfZziMcm4Zs4+3HPE81hNFkkhf3syFy632zzQXEKZH3vVvsliubV4o
vafQAQ8IvIZ2FwEHUhGqYmr3bwto4VFUtEkCZGAYrlhLQYBeJmWXfKTuoi8VtKm3
OQ/Oo0FHM9k/T/ooPg12JT/Y+Kw/n9bLlfsMiAIb3rzsWoKB7JQs3sdzVK0eksAd
C5eV2oybXsLp54wdo0KOYqC8Pin8Ox554ipP+KgZvXl57AkUvShpCYLR2xwmLVID
ktHHfV1vNQ8j+Mw46IYV30X+yPFg8+3lR6myzc+J5L+oouTzyelpvJc1b5fm4sue
glm2+L+FYwS1SF2e2m2In3KGfYk7W6Gy9YklwwDxTZlT3QG/18yLD66CTuzRugA5
irG8VbJYWzkV+HLiOktYTwl/+wBm+WC+imlAgGKPagGXy3Nz7udcZuK5hPLvI5w6
vjeFxyXprWqIl8KoSxxU9cc0lw5ugwsl7f0cmbzKfRoMoMxLffa0I53DHopiy+Br
HjEu0ZZTJ6++dO2qwsZW0DeeNfwT9dy1QhdyHW97iqoh20ggQhg+Ynw8QFF/Xgdi
/lVg7sg/KP++ocIZWvuJa8nyEYaYKPFjEemAkgv27+J//f1RQGml4ZaXJK+GYMc6
13bE/08zozx6wPTZ0ILJf0ZSJ0ziZbafvBJM9wVzZYyCmwDTWHTWGxCUaWmUOiVg
QyGod7RHe45EjutbCNMf2gFzzVhHXzVYr8J6BpblRaJsI+aygCcvv12gWXPU7fr9
xeM6Cgkf4GnHfq/QofZSU9LiMbM5UZvofD82/y8NN5cUuowsaCY4IL1GM+4cEYxj
xdHG4VKlFXpV8jGxqvmwoZ92EmE/GCYlrTq3Ee4ubdTOMkfRuLr/BCj9KSSD0Qm1
jkyap5/8zWERLDukflv5joLzdgWEFONk+PaNPPDd5jNOk4HbRukw5iU+I9hC81Ur
5XQpFYw+Gr0sM+lS9wikwALKkPDwg+SovKa7hRcxGuo9Zv0gj69BrxRunmHyu1aE
KACp80oa2femia9fNJgSp/1DfQiecJXaodfNvzpE3eT/4O32U+kpIM/0h2K/l5Xi
2PkT4VYq7LM2GZCZ/y5sws/W3sO/EGHzFyLt15+intUea4GkyP2zrzKSG/kTMZzg
LoTuxzien3c24HtVONAF9ZnqM5e6IpbELRbNwsipiDrw/myu+Aj0gbQOo53d+iqY
OOI4foU9x6/cTGDQ/prAjXMHO8umSt2ieZxx1yY0L5qUOG4YTcb/ma9WNK7UXXv1
/S9KwbS7SPkdxWF8saS0lWbeQjVzurWy4YemT7EXE8aKdGoqKlzVMk59QiWjFEE7
ebRm5al6WrAs1fUutm0Xizvn179hlN7zuRpy+VREkdxtpHJFAwKGtwxiAYpUTNfC
+7rHYp2mlHLKAIzWcFqZarxiRrvNO9l1B7M9YcVpOdPUluZp6JuszvmgmpcvA772
0AVesR7DI5KMq95zfhIv6Cqq5/NP4Y3fazCdbVnH8wPlqcwCe8krMhv6bntb8ns2
LgAcCDA6qD1BSWRahlY5MCO8FXhoUms+MWcXE7JgJEntxlwQm8Ze9sBaVFJtogdf
5rca11im+yse9hrPSJOz8aqX+8brxymHSZ9BYm+Dxu4ylOYClJPFhZF5WSaHDvE6
AcwAH7u5QMfzQ6sjOFQVz/JlvrltNblBlxM3dJuLoQFlnn8KRXxQ7jtEdc9UwJ+b
o8jc5RIrXo2BXNRH0wa4TTL1BSY48uudCKeK70RhDDIgL5LaXwxIrqWGWdxGpDlj
PdLsYiNAM9yXqZ0DV/DZxgMbG6M9ElIN/nvWuOcef7GWF93cJUYmRmTCjsJAY/+x
UwW6MBGBWX+Qz/Dn2YLylrGBhwW6XOiYkzl7nb2UG+rC0XZRngpmBXtpM0fGECTN
h7cFSOMSR6pkqUl5NEIkNu/JFekzBPyGiHQ5WclzdSnwnRFb2vUcyfpSUiBWAF05
n/IE+6d0f/8QkQfZTQSlwUdfNpyvPlZS1eRgM10Gy+8fXsjJvqu2GX6GGZAZq11t
W9OS0Yd7K569xW0X4QogakRL4xR2osq90ad7AaVhZeuRgtrPbTK3XxohHG1vdyev
T/6ar/YHLeZT5+naaNw951aU+yXEpjo31/1h0/p8EuTrexvJ+wHGJD6MoS5ajPbg
Xo1XUNPSSQgG6ahuy1rCqb1y8SH8mhOp3vwKns0Rlvuttf3upa8+gosdf9rSVlaD
bGo6nkfbTWgDNYd3jxvoaUxgwKazdIsYiBPCT4CH3NRVZFjtc8gjfGVfrO/3aZRN
IMXy2W75Eu/gnMbU74tlE51p9nyKHMpwYYfZAqTcGS5a/mK6I+9iiO4dJGT83DUC
uR0aX3Nsdr1/O9bDFkHxOxjrGUePKC0HiU+Z6NpLYJRU8xR3L8k+4FbNPqfw1kd4
AUr/rKFF5j6Ut/WnjHIGbIFSAxuegbYVqi59EadfJIr33YoO4kcRuT1azZ6IAR7H
N8l9WeKtrpwD6wUim0ucipw57QdmJVUrOSVVz7hLsZ6AqgB/Mr+7qYyETcOBt2A0
p047iGJr+ht5d72VjwD54LohgH1q6+lvhMK1rnfMMsy1KGWYJ1U/9UNm5kLcnpJJ
MXYo8nzEBtbPmKc6rS+4LSAEThGQMbnTTADxo5ASIXr7JDnemomf5xBeBd4BVvr+
NjWMnw9kpjBnNcCgwsSAKpk8/OOCM8A6bbQnBD6A9EFfSqEP1wDPRMT4CKhMn8G7
MbbE04bECEoOq4+Ntrl6Bt3qOJ5xm0smWPFrObccpnmHw8XG2QLwftg1CKMHKuJA
s+by6uGKvEWnhv9rn4gCcEGe/uWxppOOVAzLNlwTYNtC4bNp9Kg4nvgJG2PjyI8g
HweNzbBIhAukE2orx72KgX98FW/3tgnS3zRlRzzEWvEHvFt29hBZRQaOEmL6m5C+
+x4aS3rHZPMKFOlG7CrNxlU7UBPxEzGoJ7DPfLnNDaUtK6GjyPwFyzao0EM8rccj
8q4v1azdKmVz2MPvt0urmxOA+S927KmV5SfyPupwo9MslwW0w9RfRtvAl+v3qFoN
2B3tMgjCN1C/3Th+WF2F0mC1HlSR1mhiDsz+rKm+JwXFqVi+gO2QlnxdMjKlGWkI
VhVkzVvrydrUtNUHxeb4y1atkqw1/c2oPG5H4hCe00WmoUe4UeRLPl5nk39uxVoM
ylPx7EL4BBkj+IRPfAVeqCivBrh/j8RfLWTkHzh6eSJ+gp0+nCeGsepvx8akHFhB
1vkgogo3ky4Jxe/GvMLs6duDjViZDByz/IjIZlLPeDA9+DjiVgGLtpG9wAp1GOwC
S/smYZv+G6Bl8wvbWii2n5fxxPEoWrKGfFU+DXhJR6dFIA+eUGgFLp/c37q7PSSF
hxMfymFJdXYgpOsrJImkiOPceyx2mljaHlFSPt6AymAPnwNERKFySfRg9y6kl6M3
EMDog6b7rVbo3GkiPSCS4PPFzcxRamp91XjozQVVDDuC9PLniKaSKZvptT9AmQf+
SZs+SeaeYXVsLpLnGi+WikVx7Unia/f9jpLP+zn3KxKEYtaYD5HH6GKsjTllOJNy
5fm3HiP5LhhMqQzFPBLxMjb4wbCfQQypum9zNuTZy5RFoEtJe9TLMJiRsahXtyNN
Supj+8ftJ6XQbHPtXFJoRnZDr/Ab1ejpsvpxjYqXd7PHMaXm4emqx9+88jD3jUh4
lSJl+yXJJLwtK1m42UmN71gGpqn0ShoIqvo5YoCplcrzaVGnclVXgJu5/3TYiV+A
TP3xrDUh0VNqo0NIWsKn6qKySXGv22nG2v8mEwhmsBEpwb4rsqnwIIOinrrnHSwB
MSYWN0gIPQAmWRfvsz16SkPMzdR/3hQZzWol8DzQzju+owAirVQTn2EZOO5j2gmN
4XxYXsZS//kzmUOq67AFaBXouKdmig6RlrR9C5jfeEVKD/E9LupbuiJU59Binypi
YAjEzfDoYjBb+wppHolDs1uETakwicVD0Hc0qRvrLdLhRKh2TEqvwenNWvHPTKHP
cAOyO8qSeIYdK49YAolu6Y/CzGX21SIOos8XdgKD9CQskOkK29miYtGwmVQXmRti
gw1KqnA7qbcGEK8ybd42XQZi4QC8NwmJvtaTHuMHPWw3wXvJIncZTC7s4RjInCQU
ExgprE4NYVkzqUK3f6Mj/bj/8izOCOQca3DSjeOHaHZu7n5/Qd5Bz0LLGbh4zE1X
7ZSMIbUpDdLGAaNNXrpwy+YbKk479Ps3ov0BM7nHfcJhaSLQeuS9o7qgwvdmJ3Mt
BYQtoa2J7pvAkdKADLUCqMwmozBvbpVcdOT746detxNmIF3Zj0Ky28IF38UaHhJf
ClDDOWoOUU0czBpYIPe23Wt/5Hy1aJpFbkW+tDmsEsTZQO6nCfbZb9xSbpN5nEXw
rK90mecwSIhHZVBtnXI6uz9av9CodVZNf2VOkcKA/VK6NrvTP1NWdN0obtPhqIYc
NPzuegmHtuOkMlJTUUtyD2djwJOx/kE1ADWqTbT2K/dPFwrrmTNa9h9WYrPEvx5g
UqXkLm+3t+aKpXOnqMmiPdmjZ3uma0wsrw96seD9bi+UuD2mxDy5KqrD7UBBxUzk
M+FweeZxGmZdN6HTPVgkHnw9HrzcfBZkNWWptoPdQec5+sHTwQB2K8ZThLwkQUe2
B5vHFCN73wNy3K6JcqsJJG/zMQHDiQVO5PQJvwhVo9Z6NGfz7Zw+X8ZPK+FonlTi
pWRmJOaVh14xgqW8dRlxMOVN91OLDXajxUAcLK9f4TQFtGCApkQfp9LSiHp0FD31
OxzOUswwv3PVnwdaeIWhfaamMcv0qnadgZApd3t6ipHQWOhTFmmq331mweoulA9C
1Ta184hxuocYFx57JR1LGpm/YUevP/97OvxNN+2uQYLNWUW7ASjqHUvO1b5EcgHr
itG9DK6hkdW73evGiFBdBqYHqUc46bMOC4q5R9T0HEsGpMuCmSd08TZY6B8HvYk/
t1j7X7/cjBfAvQJDkmcYEkIqVas2WWH8br2jzH3j6bt6KqHAueGMC/f2+lxh/rGT
u/HKDd+WvMoUtY1Pr0+Yqei/+Df0i57ZHWVh53VPRLRDH31hBzT23bJ0L06+5Yph
o4UoXtRXzbJUQsMZmJZlvzumlfkVqS0W9aIsKqOiQepyzyMDACAb5wwAxPTbE1J7
mJz8N3JBtn7yjLY8Qtx/v8nPQm0BWAFLL3/BSrwRhV/aSteM941y8J2Gf8d+Yah4
6pHulZx0mKIS5BO53L7ffTDSjRG6VdChsNEohmOAUh6Fr8KDLtl/LZnG3lpH+JWD
KHaQeknzHqbEIwWlj15nGoUFKkGNz0Ok0Bx0aIxScfTuhRHjzDGSgiheGTxY7Hn+
+/VW/NybHzPUFi9cucYfMYs180JcTE/LDpzh6dcdAewqz6cyZCF68QY/H5LqLxtr
ElpYh2NFgOCOYxj0Yk7S51IZ41tUhzMpODBsje36rg87d0hbO4q8VpC4EilRESeK
IrkjBe3KvJKkiwdJ9p7fS//bWjL+QpQpExY8ic8Unk01UZbsUmupzv0ISdqSfUdM
m7BsbsmZVhGohyfd/QLguhrcighEiMLa5E6CEvhFuCb7BaEoj+k9/ouhEM3gVuzb
Q3+tDBU8+XCzCGKqqKAiKJZ9fy4oizb+rVSj3OHEViKgyuGwbvHNhAdQ7mQ7YTyD
WSbTd1Y1Qj/srfWBHPSUnetKywdw690vo5g8/2+Q8su62Q+fo84vAWTOAqk3MjwR
ZZXeq+lx3PLHVYfF5s6M2HgC004Cxs6GGKswnJ0p4hpoWRrC1oz3tecssDHv8Fny
rq/vj2MKfez82oSuQrElNM+W4JSEwsQMSvA9tk38R8H1LpqgTQ19MzyzDov3JDEc
WarNBc9DodbQ7IrbVROuZm8ViDVhjxllgiJlhvUeBEkEewK1unulOfXXyxHZynVI
pEgzsvUTu69Tqhdwij+u4COR+olryipYJLjRh9w1fIiahfVNAwY72hCcVtr4euPD
eOFWzCPB0Q2nY20MFvSEI4RY2d3MOhk4uDkJc3tOXgMfFGecUnRngtIOYUg9hDHT
N6n7me9LImiUkLLfpc+wkFMvHzbQZhDVkbldDZE291vKO8RVPNF+bGds0XhcaEJ2
+jcQ8CPdGTER6O2hIlxq+qoAhsGuQxbGeGXPEX5UEYUq8EMzcaoUlq/y+1K2AEj2
gwVhiEG5/2e/FZbCIV1rTMp11H0iKPQB2TInc441oeRCgcL3FcYOTycsSlHCINou
Vmk4Yu3KHANaP7RuC9EKcUZ783xp25iTV5bfcOo3ZSYg1AjW1CXjLHEsPQVlxHGz
61YcFy/nAEq/EvuTsj6Szk5hnD7jvt6YLBuTFMRnB7ZobW+rB3x4NyAaDIv6UEpo
rxmfnnbtfGMYi175LF8MebKZBZbIK3XJzPQ7zTibDfC1gHQuRtReVorsIqiyscBQ
2qUQcfu8ZxgPaDLPtPEZices840hLnLql8WoG56xp/qxdszKq9EdC2pBynF3uiRZ
YV7T7V4Z6yA0kDVzZZlVG99A5HkHL4Dg3Ag/pFYu//ArYkS3bhKTwKWDvWTD99f6
cJzmbz7Uj+BX/w/i0htCNDn3z+ThdOxYacDvKQ1LP6JGJc2LxtMfVvfSjYiOkj5I
+19cjGnVHj761m4KJvMiNZ2pKp+ftt5mSuJFWARXA1SZW9qvJki2LpQyu9SjiRqe
mhWzGFsKywOsf1HCprf/eUpjzFKP8V7xcxmT60+CKAjLaq5v77sbvqBkECt+8uBe
noDcn3e6PhLbX42qgrrPGbnrRYF5lIVPJo87nAmTclmxJZdMcrfXYkEO3ciz6QAi
BJVBi7lGPhqnaSL9LZw57S5gQW25riK209rmNGbt2RwtCk6gtmgsoQq2Da8akcZY
+jC7b3BqzDmJV9uNX8Nd1iqoecJ3JFY9BPuBzAo61PzG7QQ8W7Xx4uzgjidQBD5L
MEWHsrXVPadmx0910AyvL92CqgXvqjST9toQVqNUxj78eTupIoHGnsVwbBO3HjTN
ap7NtU+biN3N8jIOW6wj/lZvjcDMzXPCixkdnxfWr6bfM0iTGXxwhx5GDmP9mOoF
wxCUVf9F3V4QJcFYQ/G+i0HIkOFcokC2aMR3Cd+UkFnUlXjYbmt1rNhHHTTzHhs4
BZYLLVNhM5FOCsa5nRw5kFWwubFsGN+i/HTB9ydMHc/H2hJQu4c3lE5/NNLglOuo
COuygpqy7gBsruoELNjEHmPqmRBhqEX0HLbIECnHRqpmFb9CWazSUKIakcmip9Nv
UFsqL7e+PiOxzUnclmv5/ec2Nc3ErS2D3W/tFHS3ogGhdFFHd7esavY9ZxiyuZbq
Dg5PAKYqLzvgEdMhPauZ/1FWyPERzA3a0FoBP0TFQ0QR+Pthgz6fZ7z5GenLTY41
K611rV10A4PrgdenuaogyaHnJhfektI2BQ5gBvwvCXs2aLcW/gXFYyb0+HRjC8/K
ImLk67l1ETLUkSL8iCD2JHTqsNoxN741yIVWkkYMhBQ3EH8DHsHQFuDiP/RkcTyg
GjEU1TawSp6bsnImUL4YnBpxbNICJ7B7GyNaIrocQgiCz+qejeETYAwqeFINz6AT
eXqJBkBIA29h8bX33NfUlRoxEQsx2bSapHUYqDYWpQLQipRlfe7faQmES+XtaVEm
naFJiYUqxBZz3ofLYneIgiXWZfZGdL0vvKp2ZlOrHCvqv5DcDEH04AorHKG/BELO
+N2Y/jcRmi5jwBhTCGtTxjSWhdZy+pFJ1QVvPkzVqkyVv9Uz6AKXP/Rdxutna7IX
//kAkYgcxdncYn8BeomKqtqNvSEMMoRExDa3Ne/9wCVKKPposSfEdXwwbczuv4CJ
wRRf1fg95ZsczdJ2Y+0ot7Fy1BZsdQ6RXalIGq1IsvBAFz/H+YopEEYJo/L2BDQr
ixgPNxZlc1HxULp85Sv+1T3bj5s6YQVXlINuzanvfUVULVm02Djt+56g+abE169o
OhfoqbrszSV6AttKQIrOsYNCgpzxU2wiNyLndCRHZ0e71P9bp+eeYW3tIHCKeDun
6Eo5/ZATKCFggTAAhJDVlwmkuB5h2yZOhAadFY5PGCvcutw8WZ8omrVSYpZYzHXX
5BRsHHFs8mEsSjshAL+PxdCo/evvMJkmsWt5qA2cDFVo5tvNPNN9nsS1Y+Cez2TY
XDCDfteEYvViUTsHhOqb5HPUTHzAw8xiXvFGn/kqrzRYqDUZuwm/Z92LxIPo7POD
FLlrRj5tO6ilzsTHTa9wDd/961miqJrJ4XFYzVc8firpDRHelLlXJjgXDwc7z7tE
nHRzdesQQxNu4ecaoWCjB+ScuWJOwTEKS4sI1KiAqM5KXpz3LWmqagXQLoJGOVWi
HfpIf0FyZl23BGXImkNxfKOedwZWFEDMNwOLmsq+GmFXfNXM/7X0P24ED44SW4D4
8H3e/4F7K4yMGZMiqRmfTFCzaFMWWdjmU8Lpo7fezJg1VOFzvRBSBEGmXWO0eqe/
c2vXiFOOwwYI3woWHNH2lI0u3RL6yHCK+u2nIvgmeE16ExjyydZUH1QbH5WzEkT9
v79wkK7w/ZanpmAqEWc1Lc0eRpNmUzD9ssOb5M/FQBuFGOJM7fOwqvFRsTHC7oOa
RRpAVHnO8k1QR14AeujjWfBYTxGBNJ6yKSEZ/8KweV6SAYiP5c+QPRL+YM13U/Sy
kJWT3UH6eht7Wqiqjr73RNNYlYKcY84iYHFnMNNcQ/40mJNIc9b0I1m+cQz5CIGX
VshoZ4JZtXUxVMshxBSsLh7d9l30KIgH4GphK2ukgL/cO7OSkzs645q2S0GLYjkJ
wo9t4y/ka614XE+XKvzyANWyouyN7Ucy8DuTgTl+849ZOZvQ+kdArfsZpaxDXZv7
56sFyEOY0MxVwo+RedB4LYlxLoFs6DLCcaA2glJmS2KGk9awCK8Lauuarv/pXcoQ
iUAqF6UBVQIxggXGATeWbSRNm827D+5JQEdhhFJxZERNQvNRcln+ZlqiZ1jflmlQ
DX0URFVnjFl/bH16iQ3Z/2lEjVdg+I0Rzl16xaXyX9xXKbbWx4yrhs/rn0zlDAB9
HeaOURRkoqYK+E2YXRL7Jb0Giblj9rbKXWwYBZMOV3Jtoh2FjHBZ8fB9lMPAgY+x
PxtQV5YTobZ5odWPBDuKWGGhadxewZwxvg/xnUBrmwGjyyNSQmU7CYnlrlR0taWF
OLv3SRyxH8y7ZpMIbwiVShA4xhBBaUKjYQ03zsYp7x1FZHX6xV0l4xZTD3S8/Uhr
qQPYZ9hFgP1O+bWUt8xc7gR2K9iQ8cGup/2ZzRllHNOZvbFd3+NVOWqXKbtiiYrO
pOtzcOtawwTeEVxODUmqLYBvvMdDPFcPOZx8y8v2bdnEmWzVdhhPJimjmCZcN9zZ
9VgH01OX7q/DwvQDIfgo4q7wL02lo+TIC/Bw1Nh2BUZOG4RCZ06RGIUTuwGG+JIr
Pd6QKyZdNwK9Q8ZbsSdGa/+ieom6iqXj8esEAmQPDDFY7YVY1Lf67/7Rlh1dOnHo
ggcWW49aCFnFz96v7HvzQrRxI5SG2dpeeLNeAuYslx9UEHMESVx4pzidkhQ3j3v4
Weh5ch9yk+mNySqyKJaahgjNW1GqGfyxm73O53LP0BwGU0Bz8boWj4+Huvs7fUwz
B7bw9KvDBqC/W1Ss2Aa6RrtBJdprivBEDUE6AfRJ7dMKjSCmDjzybW3Xp0WBO20H
h6dD3VAkQcnh+W5ESLfdTWN4NJ9DOX4jgC50GG9ifWgYmCDX+HGtWXDbA2VCmZrE
ZQY4172LKpBh02mhebyFjkwTFyTcCyyPdQO4Uy+bGuxzOmuh0DlLkQ0RuGAevHrf
IEmV6S0xQlzgHA8dvGF6v2wIYkmP9mZZuWOtl2vBgtYqnKHpgiod16huAMoFsCa1
mqKoqgSoVTbw01BXedOxPHEMR2K+TTvZzTpA+ndBiCcIDBwZs9mqYgZGW1vf32x4
xaJXsELKuP//AD6rEmP77mWBxoCJ3Ae+RlYvWJTnI3++fOJO3j81+VG3AiEpNRPC
4CTkChe8sJXUcShbJjE1jZiDKnkCgfFENkNVIGhsAHgQ67VjjnZ/7kM2vKzbKBT3
gJhCSBRFSrkMTyvAQ/zVszYnNYhCIqCCcZJD2km8K9oFDPVRxrAt8dQAew4BFXTg
UflgwqXj+lTNLNeIxxBfQW4cFJvEBv5aMw8sVw18f6JzuXt9rUAO9Wzrhjf14aPg
9hSYmEk3FhFLf5WIaOCaSU20hAWAx0yzPAHdcTTeQuX38X3A3Eb2vvLCok3dr+Wx
5SutyahFeh06oTZK5/5Nld/ua0pf9UnjQOnsEwV0WlJvKiEpVAPVgS4U9KxNEArm
pwLtRuUFl3KC82JT+Us1s3XrpfWzU2y6/W4k6TSaEI0dZ+gmR12ctcsWN7VzzbEZ
MxYQxmIC1d0nFlDskp5VK7BXk+MZSqcGB7delE+/KMxyuL93zb4qvPHgRgfh9ZV8
ep8Ca+K2kCmt++10fpUvhJcP8acMVeU64lkybMsP63Svn94/O/Q038fQUCSRsMLC
f6D1bxIMuXptrtBUlqPpZIg9xEwFVpI37d4PbaJ+93KdN0OpX6cCYubTxiXDNPp4
fm0Kw4PF3mHso2bnvo9xxCP6LzSnZgA9bWr7AJCDH9L8Y2c0Ua6O3+V5f/9pBaOf
wpv4U/gD/Zbr/YIIj0XYYaMAVK884yVZhQmZ4fkckq7koQX43L2sBrE5l8Ow7dw5
/EJ60yUJMnc3hL25utDigPFpIBAHExN+DPnZ6v63/lGEgdr4q+1FK8dKOt9krojS
4lRDv3yIdQ41A8UciVSOT9XEnQcUh6Sa5De0qyrlbr3hgb//o+Oxj0d1eDHv/Rk/
KlRsvc6s01M/iyo2QCre5bBC0VY4RJ87l2HAZTLV0+AToGJuFosiI9d1rrJp1shY
Y93xi8nxtd8DfBdeWbI7k2nhRk77xz+RQoCigq+XhuSbXbmVwtb4pM3EKf5cmWp9
buPOB57yXvL3jSRRgd7QaFq38+vNo+kGPhLarCeSJDF8ehi/da5airr7T+0v35R/
ReqWXEk1/8e8Oh96HnxU2asFTFj03PPLZ9mKKHfAJ7bHqIAZFdILW39TnMc88f5T
AioJngTLx30RlAECP2/ARwwHkujeA4VXxsocxXlkNB8yv1SSWaZkfJ/hyrNWVKOa
2gaeAAtsZCr2XZzT5Tudn03uSotJXyPDrjT4bLsxpiPw9PmevKbd+S1PWSi8gKUV
LfcXftaj35scsgB6I0e9RA3y6kGyrvDsxkDJNTzD3hy8ETdpG4q8yWYMvYGM6L3Q
WOPjGjIj87mypf+N57yltAKjAjMdybHBX3NuH2zNDNT1yBlOrElj2BHyeSe81ggQ
/6/603AdkQES6KdJ/Xv2WpHyzM6y44Z+5v7sW9SO0AcazFgNOU/7nyrTGHegmTaq
vA4OntEFpNnmS18pwDFvuD6swkOjdcSWZr2PW2ZY1pHlarP9LeC5E0Gb0I6Y1T2Z
h559AG1oW2z8ZFqIJmYXUECxZWeR7Tt0YVDsKTfEwutOa8+EEbWD1kqlSn22MJVA
zS4BTL+Fr3q2jy76mEzuj7eRSpSSHhY9wRWK/Qh+uMr09JBNQ3dMeNxweRSm/d4S
00L2RoqHyOOYA2/BqrLCOfNgMQ9KxH+ZQmTQA7K0x9YOGz4MjKujaszqrZ3NFqhz
J6mB0kfSKXXPmIgc5UoBmO5C5/IjYwd0PU63NnKrgvMSFGkVWemcq8ol53cxOLUc
/AG0Hwhhn4yuZggez5mgAy0O1PtcVRgaCt4Wv1NsL/1upu+svWRiSIHvm1JtlOs/
yLhbp9gcaxzXWnPNAe5XJhqnVCltyFwfYYV85OGK/SDLJy+xMUERdqE+O4v8syIE
nH74uYRv72bXkCP3mvgBBx9254Yxo6f6N4LwbZM6fZgIs5hpjIeRLE4t3nnSf9Wv
GUoheW4+qcdyDImbrHbtDdkf1IUW1vXkfuTh1eUdUFeQVUxX8jGTYi5+avFQuSbL
RWka1yjR+ZhR5E9TtxQHqC72DxV+kc+7U+/ax2lGTrdCdIYHt/fzdvCXX6cDbHdI
ADh0luW1vzUvV4sZkRnAF4JGSLJoWXGZhVOxRLliofh/AWV2WKsgZmA1fq0g+MSz
hCTJTt/FuDOROjVYKDNviRM+p+XyyUREbSyldWlDkH2KBB0IkrioN7BapJPtcaBS
LGEeUTPaCTF2MrPaSxK8GbuTah1l8xM2RzHAWFewsi3B70xHi8yf7zCtGvBU3zTx
96UX6ocLmF7xWz4GVbxQQWExYW33HU6uSDWbSIh67ZEuzd/xJvnMNnUEslIxiyHh
DLN54Cuj4+Q/dAi+DkHA4eBeYH5WHhTMmowV9XWN5cIm5WxVTy8GpOS/nYj4/NQv
XSOIPwWFyh7l2+OW3DHszvCs3GJ4ZKD6sSiDvGh+QCbWaXvAATspA3D5cm7YLMx/
e5/J4W8UtxoZLdaYas81yOrOIVV60Q/TFiKjLlYueBlYy+I2uTm1qSH+HB7NFaUi
88yC69vNlMK+zXPebWjmmmLEHlg1FEHa7hqvsi6ccH+rFuq7Qwh2Fa9evyh/vuoi
E6iCC77xHqFwkZQgd6k9F26jlpZ8px4gdYNwTzGA1tWXgK1/6yJZ87EXS2tm9dvk
O7qccLsWhIFzyx5j046neTgVmb7uBg/x4A5exHHBfNDNHEipusW+pqrJBMgVy1Da
lOS3Zs23afBjK6iIfm5xMPrfXKfAwvzhOl3xI3oSBACnzKCL4yd/ZJ/0pdEhCdyQ
9r3fGUawP1tRnGhZc12IMe6v+LOmNdOHanqOAy5wxX16Wo0sA1ypAKrjB+NB/Ghs
ddLlvIaYCeVRW+huFg/RKOwqSuLiRzyUOmcDzfaOmz0a5m4HryyxXNh0y8yeSr14
E2VSNFJWSbdKxN7NARP4CBb9krxSl7DukHiUk/rwnRQUTNwUMgFJxI7ZvNf6IYYe
T205T0aSZCqokedwXXC5RhaRro1afLaeiVTn4ecCsUqpDq2XhGtU2Lzh1zBmXtz7
a0r8H49rj1YUfaD9UqCz8iFcfB5UAj72HsC4nJhbhXgrQcSkpsg/dtTGNqtH2s4t
o4eaZXz8ysDff45gt4rP9TJPGLYe+KJf7C0e96f7k3As9U5LHw4TaSrcG5YkR9F9
H/twCXPgpdpL+7iCA0nGDLT+v9gxjvuHSCbiYaFfGfFThqc16W2/SRzXeQOPloTq
FoRr8Cnxc5Nn9niExFuGmqpGZT0VQiS13lpK0Zetji+eTl0NZchI8e0yvLQM2JUl
Rb6NKHfqthJOyB6P20UiO/weneCQuKOdviegwgwU3gal0Upawks1+CSsOBmBuDMP
t+5XTvotRKgVmVGgGkf48Y8a4D3aJ2pxQ6lmPYrcABKCaWHDw5E0+RqShlcnbdkf
OMmwnOQ99SrFKuseqwFColiJRXIJEMFYRzA8cG8Rhaa5D5PMHhIlZkbFkMkq1EdV
GNYtNeZm/e2wuCfXkNIQqxP5c+hTEGE0WRbaCDL3cH2fDIF9GU17UCiBe2SmC4DE
HW9wR2TVtoYlXykLiPbPyCSg8/UI8WSpUW1X86dZm9ft+OuPJtc475jnGzH+5d/h
t9te7MB5LrP0UpuOXtewqMIOcQ50xrctriIz6Mj3hCZEe2nKSrn3nVhl/QzBufGW
5RG2dJM3dLfk3MIL3GVoNdVQtSjJmHd76ILtVOtHO07fV794h+8h+FWp7H2SutoZ
nhLJeUaWr5uQDNnh7B3t3j+dvYQCoD/C0/k374jX3ON6cLTJMR5b14h+fseV714f
fvwnKnVdeGpZNqtFakIE0acr4vZjyLizDv2sD8XCeq9UeJErYcU3mnzjqY+nEucG
V6p2K+QtO3ePtshaNIWxKyKO8sEgk3fx3xtrVMNIFi4UvPSQIzSkFtud3us6SPdZ
5SG9dg84aCvRoICs18/80dQJSIp6Fw8E0569WNbI9CHkUJ1s1tWZ7cIu7tcz+oNs
T53GkdfAoBcm8/pmnZjjAsCxpSEiXMFV97/23/E4U9Q3v4DLA6ctvuaNeutyc56L
vCtKDfts8spXQqDJDXlWNcYEKZyJ+p3F9lBR2pUC77ngzYJFPWt5wtGrWCkiY/+a
ugaFYFG+0bqta1MCIoYg7vUpIa9o3pPBVKL/UkWt7hPePpo422p2rfBZiluzmNDi
mCuxmlJpL4CDbHhzAcFdSVly7t/IbWoIhDEHmOM0KOUAnjqMfYR5tgLvgYSKWb+6
bLB8Hj17Q7MwbNxF5DpdnftZn5f8ZnLWX8ru/YM0Q9mDnpX2zJ8ehkhKXQZ8Ugcs
UDn5H6rFVNlriJqcKQ6ylPz3BrwbX2ozurfqpQpiliR3di0i/OmhPepncRzl2Nff
CR9kPdg9Gr6BYIC9OCLLTPCyR2VKvddKSFP3b7Dyq8mo1bqmTB9iBp4+CdWYXk80
alzK2v1zGCQsIgypT4gdxRFXUf+EPCeO827lwezI5M9guwkr1q4wRaCANHucgR84
Irbbbx6vWZAWmNCREj8MvtTK2EfA8XJPZRrkMbF41x8o6ASM6XCVz0RMkLIpZ0gz
+ZVFY6EmUBdCu2q22nup2RftmX4jISOqUKjI+NwWlLT1euC2tLfp+Rex5JhBMKHG
b5jd1JUwauGWe5EcMkBvCJlcoURP9hjvHpQVkeYk9jGEPB052Tbe39DcrZ303skd
6Dzmm93igH0zGWKu8HOHpiJoNlUYHEf0B6s0+orZJIlalRAu8YWGAyoRUKg7jxBk
LS7O3A5XhxgLy5TYCpBPsPwrCaWzzmZiOqOqKpJm4r3mqi7DvkLhYMeLngQ60EwD
FBRHH5wsZv/WNujIiuBkO+snbFfo6yMr+/oaSx24D+YQs4pmfH7NUzjYsANZ9VaN
zME/joFzgWHL2sHvQgjSZOrLjSyiYGBiSqOotWrSx1mA9jo5n5vJWuZNc+bmDwXc
JanqN4e44/cxrIlJl8JE3pkXO16Pe9qFnFjFgt/bDrDTn9TeEMpmK4LCV+5z242P
u1BxzlayF/eqDvGuoA/r1LsvKOkrN+tTRX3p7BbSiF9v06cm6UM7uf3CYXY/QpbJ
x/AJhyYjq2xzjBHHO70+S85IDZopJXBuoD9XYNNxXT7zQ/zWNZgZl7wRMh8wqrDO
xtpWeuqyHuBwMPz9pQIWpFb/1RCheYaSzD/qSnHN5Axvq57uPkhPf5fqJuuQHl6x
8Wg7rFvP5k/XiRriY38NokYUWCxtJR8A+rmAafOo7C306AvWuNVIus+XVfvvJqHA
dyq1tXR7GCxvMbZjgmS202MkV23DRweK3kzvSmye9PVK6YTOXLMG5YNRaHk6EYbp
IHKw1uja/auC9LjTM5qCTUXXSJiZJT2xZygL95hYEFx7TyJFjl9ImgL4xsiArUl3
6ZfKqtT04bcBKba06b1uO1ejExSC4fbNck1Ct8I1FfnLEcHSpMMpzHDJ+Er+imoS
I8BY3GyhxOKBUK95Kid+yCNcOcE8CzHPXYd6V/8fC/u2xejTh/s8AL35nFQqFObd
PFjwT7oAXTG0l+KJw3jyAwaUkH8pZezCocyqnGOYqchRCQSa/VlgXePWTHhTJnR2
T8a82bjybqceWZ01iqWNF9rZ0BXkIEl5aLFhIDKnjkTBydP7kKrV7M5hagYHLOCQ
pQau8QeyuIxRdn4AT4RDSaIW0DB7IBr48jmEr0VObtD/XjgaEdfK0CGVAf/iKQZf
xuQG0zDyxC5bptp8MnSSDWgFNuVeAO9lAhq4nxKLhN7gO+yLNbnvtMOzc31nlfvD
fmJZpvcahJGovLYy9GmRQildJ3697WJlp5uH8O9AT4/kU3hOxdgEfhVqb4I3jr2a
iKC3z/alt8Fl8RGC2/Id/hDKaXejCuKVOfvWDYLQnFCNZ8Yi+gPJMGf4bnsXVEiY
LYQkiBX77LfZnyj7kksWEC36ZOPSeBNp5RRE9+jzTC6EY063fSMYo4Ads3qwJvgm
U0KlNzwjscNG/W1rLMY6sNzL2W8HACGgWErR66lJRuERQn4wEvl/tyF66C52PETI
f4K0Hg/e8Fgf7I6awesPUAvxHWPD+ChF+pgq0w6JoaBvx+RS0EbqiJ1sAdtdDxg9
+UasHJpZKIsaN45Dj1u7bdL4g6IZRkhkZPD/8ib1niZ2ryKGVSUkArfiVC8t4aOW
444xk7cXWBNfaRSW2GcIgpjkwbKQ12hgxLACddJjv5fqyaUmYRoEP7cJusi+zgor
vFuGLUOCu9o0xbcmFxvHdDvZcJsZraWV71XczyA0Jvr2H9iSKZ1t6jDt3Q2gwzGV
6nqQ+MHoGxFdVoQhWK9kCaEcb5oTOvmKMIISqZukYzOxs8YGx04khaYIMdOdY6Zn
tjH4Lk8zIvTF8kA7oqSWoYRCBk+fBU0fh/n/MmDtr0kuVtC9Q/qgpL4cFg6Wwb0r
fbkdN4BBEw+mF98GIrjKYty9jWJRPb2FZC2+pKlmEJBkMGg3A1e2rB8OSkBg+BP2
bdMeBpF2HEYGRdju5I5APXOhR8MiY/K9kL12s6WhyO6LnHAyxs9Cwx/RgA+v3rka
FQoBD7WrUidzWP8W6JoxYuLcqdp2AcHDO7O4DpttJcrHrNxsgfzlOCNA7gMV6lKm
+u9kgV5SJBD6iEyiEUpxt07F4U//P1lxCJTD9uhraCYh3oaj9nuw464t8+jfdvAa
CoWMVN7Ig5+oP9oDz0C8dS51LUec8NYWQrF+bznUM3o9V4ItuurQlAEA9hTwunob
Wa/fW8CgczVUq0Pv2r1BTG4B+ov4vadO37RO72jXIWq0C/oSZdDvKFIHKHtvmzSn
E2pUKtixMRG9Qz8Uc1FNBYFZX4ipB9swl874MsKBd2JyxDTS0JC9yS25z1ClHG6e
0XV84Fxeg+uZVPDoPDyRZrkzv+Okhn0wQBei87zy1M+iytd3nC8AvHy9ImKVEM12
jROFiRlfxSiCfAUpEitkEIQTXczW6asr1vyZUK0LoyzivmNpeoSJ9XAr0w7bj7BZ
cr1mTapYmxby5zgrKeCZuUXnoK5y9W8qcD/KU78LqA6CPaMmXdRyPeFrW9A/k3Gl
+xPreZz3lLzqog/MOuSc6PxBEfWvmVbyIr3IA8SRFsYOg/Lbe4WnWnI/g4I4dCCp
EtWOC5kDCySDXPH6hBbYYSk4QYK8tbC1WA6uTJWtNS7RMNeNrykqUuWtqzGa/i9O
xfyVK5tC94VmuurPyJWuP9a3zhmrBYB/hEbJa/sYl/tmwe6QWgZCOG79LTjvHxvT
u7L3zBdiJrkyZnePeEmwjjvy6zwykuG2/cBGNVtiTt8pcGPIOynoXE5+qZ8r0lLF
Qm//8gt+ou3Qg5btcSSq3s7LTFzsQxQOSS02pKjd623l0DoMh5XKcPgh7smG+9jz
M4CKk5djbfCrk6SRgmSsr5bjNh13WvLKq5AzCCXDAGMe63Jqu++xtiD2lnHtl9CC
vQC3zb4Xi8O+rvXsxLJTeOKZuDvu541X3tJzR1j+TO4ZehwQRCxxcn5HdoUfvRnN
lHsqu1kT5fBOkAsuRY1WuyNht8Fh1HLD8PABAUoS736HRY1l3eUX+vSGENRoCyR9
+CorjoAxBPp7IX5jg0bsZ+W1a1lGs/WPULDin4Wj1e5lhESPhfZEdLsLsj8PkRty
hXNtRTbuR+BSgA0n6n8PTu+1nAiQq0Oq30KpvOJc4PqnSTzvD/QAtzc/AS6Oc2aC
Qot68J/QEYDccJ6pGdTHIavVDykARrh6HnMBIEEAqzmgk1arOSPRP9PoFZsDbs4F
766XJmmfkF/g2L8Y6Nxxe4IwCoQi5KJZsoh3MrBl/RSqnX8tz3O8eXpn/IR7ZWW6
+mekn9OH+IS+OWr67qAT9n/KOg6pQQUyjw2Fuuvoocg5EGxg5SG06BWagBiMJSZV
XlajHzUGJjyGw3h9GoUNIMktAQTfCXMb7BkqGzeS758a/FOZXd8FB87KSEelRf+t
3X8sCrIRxQaPQmi697kT8uGFn3jXiBiBfhEfm0HuPaSGSr5Y4FRZQMpZcFXapEPj
Lyx2uyRxSnac3DM/N7keX1leqT6s+NkLn+q+XlSGRn5qG55f6Wfesdg7K35fbg20
e+yo+vHCevD5sE/so84Z5ugybfrtWVy4c8dn6WH5pcSNlt8IN9sZeS+hzQz5mpDH
63sIrxOO0yMBurYc30cT30MfAcIt+7rQlw6ezfJ0NOJOf8+86O/kygBtOoOnHVT9
NvIuj1I5b2RMJpvM2acWTGXpoHvm/L7zOsNQl+HzWg4dhAPf3uuVgDEXyj3xhPux
Fb42BP8BJZ863RHhVsglzXWsS1gr7JSNMxtUg6gvSzEnajCKQYPZC61i0JPUpoBE
q27+cH/xvaET1bHmvlSR6brz8R1zECXH4YXPrsAXn+lRj8vxRZBTCWc1CrM/1HDH
K4RmaMjS8rjdEaoiQmJvUBgrffWcgUy3UFXtTB2JTnXz8BY5IOzx/tqR2Ud0Qvrz
zEGtHVNf0yU+RzA9ZcPefimyre0nhIdxDkZxRiTWDXXDvU83ciBhDjCQaONSoptY
eGaQ38i0XCGWImKZ75o8dHTcgnu/vB5d4sOqnsvjDZPoSAUDA3tdJjo3y/C/zVeW
vg0heYdoLDigcnxiznvkUo2Gcl2IcQ3S0LVrvuOJqevh9Po+LEvqZ6T7lwk1APRm
smB2RZ89uMaTQs+JhDdaHqRUlQrSc+sxtCf0ubK6FdtE6gDNME3rQxItlI0XePzP
nNuLLXDVgwRy6E2uIF80QsRS7rnUkmUO60VK3sG+WZA8GgCkydQi2PQP4y5v2D9G
j2NO4qlmaFAuPdnLO3bRQmUlnBw+KswCBgbi4tZcI1xJzb8/3JPicG61NrbHay6g
O53IO8/6TuvGGsBXurmZdw2CRgw6iMkVNH/IEvGPpCW0OQd0BmuXj1zmomaKnq24
NgUAQ0p52HfpbdgNrCOdjUpdvdxDJd8IJga9ceuXcz6t5uaS+R4CVkIeIBj/dgZg
XqV1m6lCbs/GJ2vwo2WrEYtOrMRETFVzdotg59yvrNgpgChECHDOxL3+5WhQbEJK
6m63qWy8KdOzBB3ReKjPMaTCFgQipzzR1pB6LHnisLAmF9DV2sGIfmGe6bCpcJQS
Ekgsz3SQv4hU2U3FcR6Za7RB+4jaZ+QnhqMkPN5Pf2VFxletsSGY8P68FvVfNC8G
IEItX2wo3rVLUfvTEdhc8UrCQw95XeZNCO4TBf2k0rZI5i2g3gC1QrwKpXYIQ658
ojm22384Vnfpm13X3Fe8YEaZm54tKcw699o2KkWXXMCDATuQjQZP6/CKSIPxsj64
8hTsiyMr+VUCqzm7PL4WGNj1TlWJkExlMXW5Wx+LQXkPtnep/3AgkfEv8LXAswb4
F6N7Kp8irQ+64+1gwWb3dVOGPoB7kWqR80OJhLsTl9Byxm/wX4OT7qBLWQGXIPKh
HK13Uo+4hxVQOqdAVE8grCVLvr63SQkciARIVBGn7ubbHpVx+7WoK3tx6g7Ymlb7
43XTBt+S+LZ2MXKk1Cy+1G8D1da+6KPlmctl40jfpS4bnLSnoAb1COFjMwTUxheX
pNgNCEvXrE8vu5MFKe28y7IaXs5uBplXvEOzjHeJC9ZQ99pOlgQVKInkvEoh7bb7
ZhUqI9kVmiWKXtevwb8bsb3TFvTJIXjr/KCniJqzG9feHy60UuzyBXmTwcE3zaNh
kwtYQ+jGeWD+Gt1QCxgDoPHFkPj43rtybeqMdI6rdfbWqMqQXt49m5D7raWedr+7
DcpqafM2/9kM71EPzb6WtmBiItnbvLKO0Hj+OJEnTf0T+TOr7uCdqdFkPuxOkJkg
8WVuVDH+bHrnAb2sttbTcmvGZkSvydjHnB47g7fJxkqt255sIMOgehZZSruo7Cg3
+bY5cP5tOvD/npsO7kaz5QTbepS8MkJ2EMOwC+VZatFTDzc4EPvtPveL/qtN64a4
gabY4qJvn/WVxIYdBJ366f7HMQD75M8WPA5SBS0KAbpWHVsW/doszrw5cuXCGgrZ
ahUHBStpp0mKOnXbLjYsN/4xT9C4CXKqBIjiCKMVL08FtDd6D+Kv5CwMR88gDUuT
9KfDVPWFFILLrSq+cEZiozr+plrptcdagFDGvvn41kgRHejB193f60cGot1xMWtl
cp9BrygQGseMCjOb7aH9MY6UjFKytRm6eMkGnRntVCo+K8iylTe6zlTW8iwKj/qf
iq4gnHh5v2B9MV8I2geaLgGXY3JyMr2/kAWO1EkLmejbS9RJsvNlNjLe74s9cUDb
+bJcsyVnT3cVJNJkApGDMC9v6wM1aV4vK1LXRW+bF3CswhGxm/Uq7gbcSfkgVxZM
Qks7+WbszyToK44DQS/hekxbyjQ6LnGLPviAkgG2w8L5a7EV8BCV2z3jgrfHd8eg
BLnkBzJlGDa0vQ0SEM4IgmyMMwKuGi8aKeU0SdHOLWnFtJzCnf7JKrXI4Wo9yctD
h+PieWQkQEf/FYoFvrXu9lWx3zemwaTR55RtDbZqLlO7zIM0e0FVhbPC4+Bu51Bg
phSmn5rJH4mfUiaM/bHp8PMh2YMsxdcHkftOTS4p9TXTKVmrSA1cxQ79mKOfHEum
Au7SYNwql2qXOG8GPBvcuHF/iEBu/xVHKpBse+PviSDnEnqsQJlIEv4gzOBSB6hl
Gc3ApGiNM8+jdEmMrKVjqwhMmvit0yf5/ZztBw5M9wvFe7I8eW7pyQQn9+kqC6fG
spOwa5Yy7hwqmbAv4IsKR5xlebNNBDrjfFm3h3sJrHpROTEPsAljtzzN15aZhhJA
QCoXOnFfdw+ao4Q61ObwkaUdFLmUrxLM7jhwk6EECZcfYDolcODP0oALdIHxShv5
8oNq/XN7X6N8qtCRWCSC/d1kQLRzRi1bHGP9aRSMquCsPOmsR7LKTErlcmbS8F8X
qsWB/SSGYzUbR9dTDUNn+s8AjtMkU7M+BIErxMAv5VDw/W/7lc4oLSpU3/yUBp76
pXAhyOJtnM3J16T8bhfVbJRwOJv1UcJN73I589gQZBkNfqm+pqDlSwU6g9bY74+B
qmCrfuRFJCPMnFStORKbpnHdPLaRzrY+m7ZkgqB68W6wlGpec9qScmzD/lH4hJcq
Ia3FZXy3bQkqQEEsec+YMUq+0ntYSXKfhyWGv5nj44St+9pjk78pb46DKDtGeoWo
AhnbBmgxKfCS0oD4PExsK2G+BcSOs1MysiIxz50x4eqysKLtW7JBviwjei9/WuVv
KhWSZiEaw7ngq476msZ2Jd6aZztOH/Hzn1ms9SwRik5I1LK9Y4T73OpnClsNgNEs
Jpgnlbz5Oqe1pEzBmFm4RUAiSZBzQV2SYpyWO/Xsaj5MonqqC8m27Vlu/p7TMu/o
ritRMYFwJVtxukQqkvlCXIKQQnHWz0MFsEdAQqQ93cU9lO8HEfRwMnBQcEqDjOul
IMSZ95/GWf/y/mfJPTi+WHDHgY3FbdnW23Jq3rTptpaGwDJ3vJGsNYXfRlsj/0hi
ypoOKvG/mU3SVJJoDsDBQJXE1NscGBt3IoMLPpPxQ7e80AJmL2j8qTZ+Nunl6fno
V38G1aoHsELpFNo+AKkDgg7K0A5Nhn1UyEqHbPO2PXm5cn3ytNymA7sDODJvG1Yv
yJ15hcEICZV5zGoEJbzMWog2TRCPiO6Hafzq4lPVNFtsaETqW7aEiVK/LLpMuPgr
PRCTxb8DIXqXse+exOsnM+9mgUiBULWAYLwNnzkLLWoyPEYPCSZZqG1flcjOzbbB
7zMcvQcOEVRlU/2poJcyFkwsxNykpxK8LPfNgngyNY0dLRIlEzxwdBW8vq/5cNya
Z3VycUsdX7eyEfhd0P6Ew0vaJ2gINuwXZtU9T1+BQ0UQLuUn751M5HN3jfgomzfX
WpM8+6GblGZY99S5o20RuaBF6pKBePO2Cvl5vMCLJb6cx2uG2yn3D4tccKNQejKe
1eKCHXE8yvW+J7ej3sZiJCWlgIaKV1i/FpZhHAdwWvLNTziEcXs4Z6gAuXCNFjAF
jyE0lllFe9ti9hFx/noQ4M9OiSCm5Mh2wjmXFNwzjOPZM2VwpExfUL/AQ/TKKrFk
Hvd8SlaCxHLC6IWTVSBHb79BEbpB+zTvWguKvbZwG7XIxog71RP0+aFBvYcUiDWu
3Z5TQzt5sFv874opSnjedkDGoh6GEKBcY9YqKS0LF2XfsDRiupQzNRUJTSiNHl9v
14ENw6aB+m/28Ev5BSMJM/NnNpJBcCYlhvhJaV3IDAQf/uMXzr3oE6q30OHswOPY
F/B9oIpi/DnUYYZzIrle0AipQ433BHTJZRvQ2MRwenIyvq5agVVFDMCSm/AQg3I+
WTHZhUoq1j/6tA6ETRsp3ptFOap6699je8J2/C6Kt79FAeZirr0P1QkOfORWkX4l
UMyEN2QOaCyBM02E7tAM6KCLQzNF8sZHRnZu5wIzUVmo9MOH0JLrgi4MW0b0YW+l
LFCY11W+LTQhTIE6RAikflwvxTHRovddlVaoo25fLlDAzcpPsuyQE/GAskNwuXfT
kllFzRycEmgIUfjo4XcY+0I+drCM6E+YCY4gsbeHx7OyOs4Wf9llnLWjiPHjOn7A
3LE4ufAGE0u/0t3BoDS4r5aSsmb0YC9YZIywdjIXUIPC7QsbeIs+oAME35n+fdGE
OewggruaRAdye5eoAI6IhBeIw9KzUvQwzLBT15J5hz7aURFqznDVzc2B5CIFBwTH
F23Cx4VniyFnzwbVX5phUK0WBeYOwIqisZ42NGWqeSsVbEN28t/r4zywGxVj+mGZ
aEoMwHJLDFPnbh4J/CXMjm99EC3pTnbrT8cV8MrwZq8hrneeNjO7n9lr/PrF5v6f
IEiQMaF2ALq+mB/bJ+gIJZqVb8cFHgUSVXALYmBB59EnfiXgnpte0Bvf8UP4TcMs
f0grkdHnZ3RkbjTIy8um/3CubX3xf0MFc/HnQwqOd3mVbZOcZCEWLtiJfUtTrdvK
SfwQLmXwpg9NKbznWvEVz3D3X5O5O098QeWiyMHN45+DEDveIlVNFBP26NuBqJHB
UhX3M4VscFldTWUEpHJWG/nbf/dcAMnU98oy+3kJYc6mR8YEmJkGPAOv2V/hfnJV
8quM+hobEBscPQ/OEl+JJ7GVhT7Jm1eioG03uXykB2+tXZC3jlX27naC9CavEw1z
k1mg5lICEsu01//kcfM/+uo0b5QuQhoLJ/NBSM+/zmVX1iZWc19WsooNaceZf43i
exxFDJUrk02UjkZ7sXIC9Pouc7MzaZ0rIv0F5qv816UG1opYjpzOfk8ZHIqQnVaq
lqNOGBiCI60axSa2ZG+9zPgVwKeEPf6zg/PI4pDNl6wsTg6xkA62bA7zDDXRmQpc
3RlmRQE599vxdFrsG1k/V+5wN0OkVCZ5o3jchK6HjcQ/n1RzCnXGsWegCDvxw3y6
y8jvPBH5GSqj6pt5pgBboruGmX7o9dxuTTEZShYRKUSYMGGwRIfTzxrlY7BLmDWq
PVcqWz6M9UEFL4dBYHVfMmq3uGXomraWWe8V1R+UAxDGth2VgUCx3s+ZoSxVkl09
geeOJ0PYALFX3FeWUqa9rfotvkxJ6722K3KTvMYekN+5cHVeYveebvmSCE3kr7Cg
mtbK9dCUzcEDGlE86cMKKdJHFnF+GPZjARD0bYYC7tK1yowSPLdf3GdBdytSZbC5
tglzPeEoVVa+X3z8ZkaV2pE/k96xCEZ4eXC3QAw+fVPf+UODov/EbVHk6iZR8Yel
aa4ERo6w/9pPEBysR4BPQpMh+2YSnj1FAV3PZcX06wknQR/Yu+860CG66SGEAxh7
iteRqw8mUyxbd13fRWYLIsyiaPTpEBY6FmTTaRDQFeQDHO/a0AljmdO6jXb5ZpQN
bSMldSyrENp+B20ow36nLeQJqe1NzQaOOu46MCjI78WwFtRgM/czhLAzM89KjmEQ
vRXxg2HdyGAZhBz82W8ESZsFwDCm/9zliObyGP1EjdZGNiF8Ij5a1FitexTRjhuu
Sh47RWpJO1tZbaChyhXFPmzlejf3s0W1NNIDEF0lgI6T+s1XXJc+RMn09uOW7N+N
KXYXN04cI2u5ekZmFsHdtviR1pxYmQVNnZKZjQ2YKbdzidaq8a/V4bRcdXyX4dKd
4Of26z76dpJId3NYsXwYQSPcAQofBgpA7lhwcyLPnKJGicaNZTPKN9rGnT96fNnS
o3qLXEnWZ8LhzLJhItvYNcEkGVEI15BMMESL+gPzmxo9ma4qNk8/oYLcPEuN591A
NSB8wwI0XCN1aAZJcsaQ8dH/YeSBRGdPsw2cYlrv8m2BjRxRbAeJXNT8sR3BOkIQ
s80HXzlTZlwy3m2Oct4qTLG6sNqsE73kAU2RP1RxX3//vlVDv7/Um5DUvrBKNvw6
5Ic7EsOudTiNLdSbBpE2HSKY3FLvHaZZA6YTm08gjT7PU+P476jJNzW7vAcBiyky
28pYGY6hoDfJiyJdXfhw0Ucb4eGFsDZcsi4Pi342ZZKsWgtE6G6odBhfb4F90rtf
RMk2Pr9GJyZXsUkdge8jW2y5wZnOEc3raGT/oKPWVpvK+MDZcW16RfGTuS3zlAxr
DckY74xAh/IfmOE6+OsQ78S65ifpYkXdfHZRpZ05xd9Ex9ZNHEWImUEiFAIYJ9wK
1Sj7G8ot98CohGwjvCUCX7OZfGlKD5Ouzzl06AZoFviy5XZg5f6pTPtVrB5Fm6j9
c2wgYI3fDFINUJQx5T6OfzRjdDryrMgc/0KUlI79mlshtkisWKH2xE6SUsne33oM
ke6GLyiqPa38b2zEXSBO/C9RnVHqZl8yovlpPv7zYAxOaWBRZLGBn3BY+rhTeqdE
ujIGuRxigiLqQYN3zLa/3Ov9KFffhhZsQ+5qyXE8zKqZCrebe0OysxCMJR7jNpZA
aUWX7qdi8oDlph071KAgH0Zj2e//gkvjjXXY1uEeHswjz1BEmQqXNl2WvCgseAVl
36M6GsUv1lPoAZoMFu9jhtsrEYmg8ZXaZi5OinowROCPOP/hKGdmcNg7gEG5gWrz
WDYmqOoT+mdWk/IYnqBtzXbIpyr+/saYEkqTNfjG+elt1GPfHKRdcp9WjxUt0zGn
nGAKrBdmsEbLfzf8VdlmNZU5yURZNkolxPIcHv9aMp6NDXTFMNxOz2LKTYeKwsqu
iLaHpXY0qtbzjCkoY9JVKIwuMXBdOZGGFHhCETlzFUNXZcJN7wH2tH+kdRELMu1h
akqioaxvlsiTkTg21COpUQxrbteGaSXnLIZGF9m+OQe56vcFgpp9WF5EVqpLDf2Y
KefZAXT6ilEBmaiBZbIXtJy8cc+8E05RoFhDZ7aTdvqEl44apMk3qUIeFEMx/lS1
rKAYjmkZsAvyXkMmAso8papwQo3IWwuUxwKfxmkAWJe911mEGX6GD9bwLrFtcaFa
0R9GuKF/cv3ORdOjp+xbS/e2NCX8Q4mS39qAmgHYMw37dimCEAiw0EGhRPkVh41E
XH5EKNojFsTwVlxGOwxoEdAVjl5N/uJnG8HhAHnMRCGqVc56TJNldN3i0vV7mhEl
UkNE2bpjxTMSMlnS2MDcBVuwBhsTrSRqtXeOSjxIf5UW21VFKD/5d+/TTARR/e9t
Toh5X+EpJ4Dvf34lN+M20cxXTOft+AY8DibjYozqIhT3l9w6dfUX8HfkRA40ggJo
zAe9dy4/WtNBOvpDXg5pIJcwIFXpabxVmVfcujNI2yPG7eaRL7jX4xbeeeL3q9KF
llU6rEy4UQzDGQFOU+J3+jm91YgoQFwzLrzC2AEWU6DjKzXc5kSwe6K1wCWWfomI
TZqx6niORuv5HZrBreUd+scO1YRyPVqJAIEuemCUz7Xpb0Z3VrcK/BT5j9FPZjR1
kqi5MYHSLujd6nd4V4i6XmpedgggR0MQYdLzbicma5GEwwQ5RPmLht6YlEqWWVV+
Vrh7xSDuTRFGzTQYpVJLvnB4u97cPTR5845y8xQshldlhuFnmDNIjXABQX6mKFeM
HfdE5u7O2+nQ8vyLVWkG49rWmcPFctWyi2DlPKbHkPRFgb8OTQmg4SXOkmmB8Dk2
OE7pt3XGcutXSxhNPdP9H8R/5jGsvkZih7RW8eiUZHRUjNqmnK0Z13u0Ffy73kgw
CGb5oMV/6zjhmP2jtPGW/JFnLPJWtScGDc1B/kZWWItPBgzyxra6kWT9j8G32pMw
/+6MCIfXtiG1fpgOCgt1EJ6WjDIxaEHbRqkQduK2F0ZDtyuwD/ePyT3yhExO1R2V
wPQE3S3mMJCzUL0ZP99ZmVd2xdtyNGxcoctstPvsWIUZ+11R8q/HgN5A17AZ60n2
4RuubaXM0yOYmHtXaClzbo2VvWSIpb+82BZiNvMiYtP9G3xkErL57mRAEX3KoMqS
AToED2R4zks5miubxWA7YYl8vZJZxd/jr3Wtd0ibPL4+BOcIRsy7R3fw6IXQOAGY
2QSJ7AvZdgmxE5+bZvKuXumEymRLYsjtlCCv0Dlk9r21WAaGw0mo60qUscWfx/ym
k3XhM8fylGxxX3bj4TTiyZgQGqzNj3MPNaN7miOpmoC0+9i4IpvWhtqI22ETSP+r
1qSCUyV6RQVugzF/egTey7Lq5Np3/fWypNF81L8gq0KcCuTfzfhOqvLp8qfxnBcb
ZgqSl6wnxuudN6ez0IK+VFXVcsayG3wM77eT2cWJfqEVJPGk8Ih7VpE0ZEv3et0a
ppsHCFW7maTbtCsEuUoR3WnfrgFwunqaM8eIRR+ywC66Fv1Z31xU0EdDNQlVdD5f
398Gr0LtEId1pedyJIf4n/RTQ5GSa8tDSj0Gjt30amzigslGtl9PMwkGGffL7RfD
hfMAUghxtGj55xptp4UnfauQUpe5x0Cu8oZTD9ZZjH6Su1Z+i3cZm8yU5vVrhlDV
vnGPBR+jJjTaJFU3ZHhHDwPLnuFrrvoDdYLAA4o2tbidbF8xKHDP/zI1460T3VWz
Jf6bNDRxaEEG/g5vNfwAZuv/0fhCJ6z5OYhXP50CBh+XBH+PbYJS76x5gMLX1hNl
HQ/JXSgeXom2j0cdUsDRrQ1n6SlUypVYJyGXArGrpC4hM6Izi1LLm8WeOlukVbxC
Rw5POcvVeuHEUS9BvR+4lV/kDZF++qAInd9dmtJ/urLrLqxZYYe2mLWG0ysgP9zj
JF6tX95EFREh7c7y9mSRBabkQ3mz+HGls+Jaqh+UAocecmfqw8+HmP8EX08bNaX/
P+ErvnriXe8RvuILW/23rF0d7dnKRSA3K2IYJB7Q4RSNeHAI6W2ex28WhiS0eVh3
nhECVAmxpzjrCUR+qOZbRls5V/EucEpk7J+5BtFveMd/V1GL7J616FiNg6YVMr2A
oldDWtSVSk8ekOaJPe8EHQtE/xtpvEiVVx3QYPxxc6Ky9Jffj763qN3yaUMaj7CW
8RmRddn0Z0YPMZb02krlxnDvXdk1QRi+4kYbaOQMauZDovwM35HEmPSwAL0UVw6b
X3Ol70eaXL5Zg82fnpPV3z9A0HVefh+aJ+7QhGrj5ltmx0sfnFrPKKNiAd2XxbYa
MBnyLPjkGHAk1VTONiXrw1c5fp+RsLRRpihLTrJIiR2TR9h1tJ7dzGelmrZ3Smq7
x9+l/pr+M15/xa69F79F7BBHEVgW3ux4nvoc6n1iuoThMIW3YMus6Q3vzIToh8mT
MKJH0aCFBnJ8yJoOFsE7tK25s82as/iHP+gtF6KKzN1oNt+lRqJxrzH2i5KWUlLk
Z1CmIUUVWANU9X/oQdOICNzIhz986aBBT2DGI5qpKHzAIgmlQmBWLQc7Y6sCtCdH
IHQFgm67tWJ269Wvs/z74g7w+iRYgel9afbkpyvPFOT3gARwQj+3MP0+ioSBrgoz
vj94vTMXJavQJUZBvTeAj7gtz9nUchodxfCvplZFgKGDnEnGETleoqRQ89TeBKQi
e3FLR3fW6CwlWTa04uwhWSMbLNuR6Ay0dstbz6ipogxgMcXQ5MoEkHXEOiGbeflg
+WAnpnrD2weu79siZnkRvYf8PHFz503HTqBUuc2Vzy1x4zWQFpExkIpwxkY/2d2x
Akwrlyo/vg5So246z1sybCR5YpaXv1Xqf+kSWzkqQndr2Ts1s8cEtFfw2fTjjEO3
oB8ZJdHhU4I5b7sN3s2Pjwy0Qp5lA5xrpZHLOO3sb0foyDbjecWtl+iHa8yN8+Jk
ynNrD/3teVtP2JdaeGyC3nkfkAiJuUW+MPgU1Y19ddN9LcCGPsPWSQ77MfIo3eyj
aUx0EoZfCp5YHHLyTXXROvnEFnq33Uq0vBvdnYBg8pnGa1YSLj78Glp7QuqprjHz
SiZdnxGQAiu/gNd6/a6ACBMT/d++Ow4UGpHAxxErLYp1BEAxDwr5YWB/JXOcmvgG
njUeEEj5E4I0XqzSZrB0UtpZQ5Kg0o2Ju1VQC4ejvYKxzJh4JHdcSW+/4Y62Eu12
rjrT17XLVdLccY0Cd5kMN/EoTrluLogFjjkvL3LophrjEUfA6TwG/HB4iihM1cha
VmgbMUaBlro+zEi8VL+Bbayw0UnX0YXUZgBTDSBvruqOHfC24XdUWrntX1TZNqoU
puJopx4x+wzNHNH/DXO19BJrXF/6FAP3Ci6jOiH44Phu1DL4zdxFlMrEV96RmlHB
nLZx1yGwAvZhHo4jueYX7wdl9aVSNpoa3WEikDjaHd8OsOuFnYfmQ95HNdcT2Grd
R0Ujy0bv7rSYelhz0UKE3XgSfp+obNci1grZASvPRDCVRKBJNhvLa21fRClvBERl
B2aUaUudhW0mwBPxBHh95zvDaGAm4wRp1OPIRXM84OiyeBu78HCPOALiM44j28Ub
Sf8o6c0B3l1Xzh0l2pkjTVfNxkVIsj2m0ZBrU2Ur/Yld++yiQ0BrVkT/mkSM19xP
CMy2hDMEjvLNKRW1fVFIpF8ph5zpeAG9HbgieYxfpX7My8V1s7kfTPMKGgEXKIqA
d6KpVZD7YS/SFI51afIKg3OR2W5uPrnk63GuXMPer4HOiJBFz99k8F57F5n1Mf/E
fvKbPYusf/A3KSjRUdWj8DZDHiUVyNN4t88E7UOrpC3i3Pkk1TIIc5QDxoCv8GRN
OVqd1Ja4GFbB16p0/Dmcox4L/+X9VHRk486ojILgy6Et/oGtucpg/iUBCztzH1gv
1qnCmz3s6l/HcynM+eYtw2aW99wMlpzbqir7O932LcVQzcdergPJeI8dB64uutSA
5S7uLPaRzUuzkn5tTYy3TE+kOu7RnxgW4c66D9wk1iA5zuYgpvtTPt9ZnjF31L4z
B0QFGP+UQB9Xuoa3wlqoWH2Z8DXI/I2gmJMeGcfzSVXrb+ydmKLafnun/fSksheC
PL9QNIhcy6W4mSiC4F4ClC9eqDnN8OVLdW/OK+Vp1lH2n8EDaVink4j8yHtocPQF
3JW3Tb19vf7hsngZjWXF7TDnEY2kPU/nUR9ji09xOQzH7FTLFhnLx8ybVcTPvuI6
zcbTw9ufQZRjEsw5O7GZPIefA+adU5cpsgmTI4fNaDU2pAo8uP6HBj3P7MKTZU1z
BLpvA1mb5i/GBNxcAGG3EQBkuIngDtJqI/14C/NWjI7Murk6HqSl2mWo3yWuHNbg
DmhgzBcQfm3AtCZjSUZuF4qHLx2ANlPNuDilq+5nX1DCf4PMriDry32XqBeCV8gw
gEee+nWLJo0OtgOpFVJ9W3qFJpTU+AYuDIYmZqUAeicMYO9rb8AQiFoG7gjASQb2
EqOFzswMrPqyOc3ciJKY6V6ZFPo7ju7vOywp44NGtU3EutZo3NGEcjGYyxElQycj
6VKJi+j2gDqPoe/evUfCyU2lth7GSXbTi6iEuVbcdJK8p9Fy2cb8SBbteePdduHt
9kV8I1eLEBaPAqxMXRJw2+YIqWcf21ELK6an+h7mrVUcoi3vKnWQYj2Byr3vwE0x
bxIJpF8LbACc7AeTmkcpBt0i5YkhhjEejl1LVIqk2aGlVrvfoMACfeYTEObJmIs7
8dS3kEO5YGRYHgpnju0KZ8hCRt0OAcceZutt5EX9Yh3obefcG7G2NUKm5PHdZsYh
SUgu5z7KduhZMMZ59XulyLb1CofGhmp+jmvjxkjgihQUxESTZ1/+rDaz2/BR7paI
zr26rObnMFKABNFJ2AtX7BGZrBFj7by9S2nDXAn3Z1KL+GkraHPOBtKPOOh++ufa
eXUHUbeYmuRFWIcFwWKa9b7gmNhlMqCwAeNqJvnvltPYCWdwEdxNDla+2xw9DbdU
BqTBYbOarFuGyC+zjzhhtLuX169+Swsp5bxGW1Xqrs0TVYqbi5RFpcZ06/p4/2JF
Qy4dRglP7/goBgr1xEqjiBTdpWe5lf2GYp8OLN01FrMH9cTa6g1GN5YcQ5F6AAyc
jFxl4qZQBfP+S7AHULSg3Gs8hmXxCURT5ulLGqS1suW+/HEfsiLGWFDaSexzZl+6
Z88aDn3sY/F5UzeABzwEhH1yRSq02OAulRKMW5N48iwHY+TEhu0fYPk92umSGMoi
+jUJd3B7BcODoddEX1Li/A3IzTfxZ/igsH0GMNlZiB9/VEgyz4/VMcNpR3Rwelsp
0TfgZVyQ9HAxIoqQ+/tf/HMLVgZ1kG1ofjo7w623cOdJthc7u+Ko0K8E0YtQ5svu
74Iky+P6cLQ1wcR3ElUJvDmnpR+fg2S3y1itfnoY+VK+tHiR6erxcj41JILAzzDJ
aISSENpmW6UDHKImTJsJ3IljvKH8Pdj1j0FhiYvaQ2dvq3qTRyV6jOCWovVNB2IA
X35OYa0DQEGEnlU1O8d55eeKJqMABh+MMMOV9qVOBORLmn/qZcmv9RCE7gJcluEH
pdN4GYWkhNH0FF5dUFzWMaRQgNFZgxvBQrxQN6VMercaCz86nkhcam7HvdwQydQ9
gZgWDdrN/YPoa0qRrSekup8AJObkx4w5lr59h9IWDGvenMRfBOwvKfZiBsWqUNQ2
vb3w+qNVn+gVBHfhw7xpt92mKX+bGvDQ6nwLp+soJZ5KT93LQtyp14pLXERC2O0c
U7QHrpND7SQsnjE5fQl4g4fSckyEopNTWhisK22k25cDAC8AF9ZxXTsFAJh/NUeP
ZXj1hb9c2eGbVxO6xfWodrUeXGs+dNKj5+nUc8Hm5w9tjyn4Y8OZcKxSjAalWQpH
wx/BGLGqw2i7ACJKzPG71rJIs+xyMLnuGeRgFRuOaLnihn1Lme3g0qY/cyBt5HMU
8pCzOdQsdgb+jE5BGYMg0rrKesBJSkBOQ4DKn9uk0O3ZA3+LXWMZUFlT1JEJGgLP
+OkNx02S2qf96eSN0vsljSWpaR8CjJ+KvToRCvy9vTO/cMp1YoxZVC0DJ+u8zg5m
/5WF2DIEu+/EjeNEOquk6vQbOJiR7maL+so2KRmmSlWjkJR+v2MrhE7+5ZdqHSSv
qTiO69ZoC0QSmMHFLtZRt0JCGHx+Px5umPguq41YiZX5SYivTDkCMBtDpEYJDukL
ck5K+5OALesjyDEAV+dMqfhEfs26CE9nhIIK6L1Nr2msHe0JAstUrj0nfiQH/5qv
xdnQxNcjnZNWgpRtm6x7fVFMCMJifLHlwnSWjJRFjKXVhcoqKtFsWm7wsi0IWo+Y
dPWjEH5qsvk3xIZWJvQiVo+NZ88ukYZClt3Q5lzaYRsZfDQbztaPv1VpMaqwbQHK
mYrc1mOMEI8uuo9th/HiHYEaqDSsd+7KBf3ADPYnW5Ilk7in8zoHrgDEZsM84AcL
GQRu1IwaW0u40ir+UjNZ25PfdJzJJW70aS/OuoKz6dt8AajJwwS37ozDHnSglvvH
K01Nm3f1ks3B3qb9K4fGK1fbVThYgmOmMdo2mobR+TkRcnHXDUuq1nGOLHbrWn8A
cpXEX+CqByNPxT7TseHt6SFxgREGoz/spvlv25092e42bL8TdPdPu4OOvkIvNpFj
fkgT1eIeq2fdLr61P1P3HyWUxO5QUvtLuXi8Ur5hnW+pAT6zKULg9fMd9HhgZHwG
ssLHryKcTkrw2xAyFY82bVGrPMyZnIyg1NmoBdcKI/zGMLOto4oAjfCVk3mVTEvX
z3K8yVthKpuY8ryoVRu0KFWCg6RNjz+1ir/gwQKHrrUmMbqj+mX6aFRWNxze0MlI
QQVC3E2NudQCq41AQlOCcBPfMFoYWFuwbsy/DRRGlbR2CjtDOMOc8smMGmQfqD8Q
jIahvmGuaCqUO8T4jWTOX8eeTZ1dBZYzyNAhsIFgp7ObdqWHa7B75yDjA63QL9wP
BnH/axg1ygxGi0cNEvogYmewkmki8TlX4BXfV9Bbpy2HMuiH7JBPqK98m+7+VWz6
0fT1wu1z8JkFCesO8FH4SVFewb0LQPS46srJk9uotTb8b7JK1I4sR2lXOMDLofUA
r19lWPozMoe4T8TLBttbZR1ikY3x8gz8q158KqQnkiKUTCw/bWw2W5pnd9WzGtw2
tRNFl6kM+DZ7/qcB1JZW4Z1Z+hYik0Sh8/ng6i2w2guFmAGdRLilxZs8rnADsjGt
fYVWRlkSwYVkERr1el3bu9N3kDUEjx5zwaWmEX6rE7OAkykhTVA9+v1TD+cyjjEU
AQtAS86VVe55PpxAlBRqmhPOLDRCQs/FGolcmNFktkRns2FMEcIdj9Efu3HPDKtA
HuAefEsDFfHd8mHxbJ1G82xC2ZvC7fJrsBL1cw6amxmqoaIz/VIYxR3amF4FRMv5
IXEq31OShDAE2bsvQ86O+mUUInGtrsB69ID5hcNzTm0R3Dxk5qbJYgRDxrhMAod2
/ZBPlcBsHmOXRVFC/3zkiYJaIvliXiKfhoT7juLkpbDUQq3T/ZlO2WOAdhl7JBkc
PjJiyhRJ2kA/xblBRve3+OHIZwBX282QDXCCswUnSVjJAXHGRj7Z0+xZNPl0C62w
L5fw0LzjGmRj+G0BNgbY0SbNA+Qw7fnZqMaMrmyqIx68Opb5dP3Hezd/j2o+DG5N
cmpMraOHG6uP95wn8OAXXiv+eUdbnK0+uuFXEpFDs4vLzLyy/SJwn9oZTZOHubva
IlzdkY/KHOzY3XzOSVTtDSNEeWyZ1XJMlrUo/RucXHMvLi91aROGhkxV3rhoPj80
Kt/rBwYvsaesPBGqOpPNH8y5Ocs7xL1I98yuHVeAMpxhpm+urjAWLHu1b8cHSz1t
IDCRV9NVeBxHqMJpdXVyQRR/bgzMBUypzBgYRq/CnGc6z11eg+Oqsm8IjuOybNHJ
YylDGCTcAxD9xJMYCeiH39vFiI9+1s19cNnYiBZSelkYMDmZZOV4znLSaIJruiE/
UQPa9GASBdyIBnQ3sSu7hwEmqJqLUEMU1l0+wZUTKjB0Y5gV1S3ra6RprwQrBpap
FOx+Nd4a/mlwnWVLkxezP6h1NZYccIMbtCP+PXmR3FpW8VEHb86euiC7xFZ0rXxg
f1E3m8ys2WAZlWJAmBpQOB+bzglILGcumJBAdKTzAk9sIyKDxOE+OcEd6oeZfMws
fTe7w1hsmGP7qMdyNpNeK6vHb8JlytRyqjRgmXRyNwQ7OWF6TT98ZzMFIYuaqjmQ
Qi12ZtkX55nlx8YfK4+f9rfWQMaOxLU5jgcDf4SxCh/BBxMZrUWgktFiJJqh/EhH
dn7oXqTqNszt0PjXStNbMIcNNGYMFNL0yN4GZfMwdPvtOacnlVRGPRLzsOrQ9UFH
eLAj9kbE8Wv5aMaMkWoOWx1FzBk8qFJoBKTIbw4pd8LjfOvzD/VyVFn5k3ACJ6hG
2+lrQQlC/KOLZNposHtDZ4h2u5kIpYEQt8S6d8yoMbmb4vtJVNe5QmJqD2tneOUi
AAc/rPWvekX/BPWXJ6S5i9F/SJrykh0GiBre/F4kFsFzKaDFd4PzPQlg2yb5G6YI
4yio9/S7DfXL0K7oGpmaih1DhbPdIYixDSEYZCSfE2EaNB8dKSrIWQBlMo3KmErA
bOZ8uUKsufA1FomIf2H4EywUehonupWADpKoJyoTDRQNrwX64c9GPxMZ9i9Iv24v
Tc/v/p2dlBu1YMPMdgQZp1Wxrvo6xP0OX9bmAl3jJx99aO+R0LAAH9CGzfiL6Zn/
oH+TShVZUglBnwvlH+NABn2WWXrE6rDUCKutiHCFakAN3xLDnJoYrWZz0YAhQpY0
o32Hry8PgEZjRSfa4sy0ULLoNTPXVprM4lcP5Kkleq6erLuNVXBZxTvFX2eO2/xI
iHzxLKqez+le27IndqqR0iDoA8nXP7JJCIAijsOjP+PhfivBICPWeBL87Poz9UJT
IIde5UAOU/sHbLbVTeJR59UoApHUBHdY3L2lt2vTb6wzwGhN5FqvFzZZ3DZeClFc
MA0gchnWIoIcsosRsY+Fjv5MZ+UDBIat1eXsfZJaZWHU9dCNTrb5IQqqNhknyJHs
qAf/RDDo6Iq+ZZunlGZD0bznM9OdB4Z4LWcrBqDfZd1uBALmb8ZXB/4eVhbOYnsD
EvKJDaPeur4znl/frjsqsXYbo59AzwX0oPX1uJSawNG39Mdsd7rczvPNbHFr3lvk
+9IqOBMh3PYvurpRXUB/A7A7261kiRyfFgf8FUoIC2O1/5gFOzP0d/nWxsfRn00i
lfJVh9K0eYSC54HYfqwMMtHtH2oE+yQ2w44Fj3Bl/4FZZMrmkBdjILM48E76uVDM
730jMzvkLm0Upptw//pPMLgTY9BoZIYIPWtFW9YNw5CNYkl/3fS2uMQB3Lkr2Ii/
IElllGg/CpL5mB/NCwSAq3dd7gFaBPUbFbMSATZaINuDV2HM2CwTSEfII8RwOflv
bYB+N2zrc8EYd5M9jOucv0v/0qIf/DKi/qR/6JhwxwNWJ44wCzhaoQli4l/j1w0B
PWkWkZw23a00wvkwLHD9z3JL7bSuFYHBax6ReS3+D4nwZRDEJAyWc8IGLsCfyknq
qfv8ljJu37rL/xkaYQOg+OBz/JNiAuvjkj46Mh8ed5+wcixktWyTvC3m5F+3vm8w
3aRrlUWv5K2DbSQ4q7TjvKE5vushXfIXDGzCxCnR2Gs2t3vOvzTMtDb3OFs36TBC
Dl/Ui/S1UcQc9xbp3SdOceL9NAXj7o3z/KHL5LuUUHEa4xCy5uP1K4oe4IqwG4yI
MKE3S35UPvZSZHc4/uN0omxVsjPaU4/fcYE7oI6T1PvGwuwsDsAVL5JiIinBis42
METtOz4DsULJx9GQK72J1lKJBhsCtzEI9ENUhkcsD5EbEBS/FQDUDJQaqzXQ2LG5
0sIPLpDICUHPn4QTHh844UV/8zrolWF+gi+Y6r/sOjc9ZZxl0wNer58rywDkkDXt
kzIY59ojo5NyID+EMr+M/v4aBuZBfpwy1c0k3PfZWsiPPoai5//D8ZQfYTvNk49C
Ak5UJDxtWGQyVHH6TGJRuqyeMnczMBq2GTDlzWov7Y+ecHQONhfFeH28PHmV0KMk
JiUrWWS/HzzpGms9BPxgMLzWJ6N4z1KZa251bdymf6ZM0nPDMNpr4qoDqRRUf8/J
lavrLMOV55qvmsXPu12eZBWr5REdsOsYbhTQlhntbqKY8/z9MIo464iniVAolIQD
VAse55eKkZWHyK/63X1gKKCF9Y7gdwAwTIsiggjn7ipOYOBgXRHDekFrnGyTQgJs
uISmWmVO8M61GaRkVj76PvW5gdAq+9yAJWOtcjtleJNT4fFOMwe1LSZ7oCREdD4e
RLIzRkz7w5xE6eu1JJlQgp9bqLP4SKgs/1xrTCPpsn8h5t3b1FTVIWc+XWzmPQ5N
spLLQOgL4CQvm4SDT8tVntSHMVqNr/Hxr4XZkQybcBF0pNthxeD2GvKhF+rkodEx
Sm9nxvABTkAOcpwVZS4L5yt+bTToOf70hYWiOHoTmr6KQYpJCpD7Kyw+LkdfY6Jp
okOGXyROdPIDs3vIDwOcCmrrHmqotdONlh+wYj6NGDbnbNijwSGR0lCZhpmG2Ptz
MxbAIDX91YDym1zpE35E8DKwYRA81DBMv3KOWmj9s6gQSoWPqSB8BDzvb1FtDqZN
3xYwOnkANZo4rQHYRZxKKD5BIVhta1JBpIRpevNkjUcRZaAC+xGBxiORXRa+h0hk
e8vDU0zCHdloIalb1fEoEQuPibUatkYVrAT7X+kPgqSgYUgt11hg1mvkA25qxfp3
2Ie8KZok2RldmJIsCK1bdQjLZSgrvqBYRJDFyu1jKnRZfEcfQlsAQP7n+RdBgDLD
4NhSkmHWi80jZoBXxDRRO/ZHAEqyCPMv2z7lKMDP8JrAWQBohWOLiYHhi4LmND0Z
TK3cUvz/PDFggKwbx4nzVdqG5UIRRUwOhUrw25NTJ48yKke/qkBYfkKAgWsg1rDz
HjAKXYGAgtO8XuPuO2QLw6c0SIprl/wINTGhDONstMUybq309ZvF0mYCmEI8gWWa
07R9o/ILoWppfu7TERkyEmdtzLhC4mu+eyHyeTLEQSne+LtrfU7pnzOe1Yvn3rgK
1CXMdj9FDAOHFPqJcxNA7cMKHGeIiEnTEDRV+ThyNgaBKJfw9/YVE2ARw52W/hml
hsLDJ7tOOpULxen5uCL7q+GZVEofsKXWbR5kEnm9tQcRrOaIMzOXA//IXrTmu9Ef
mefiwOsblIlcc0Hrg6zwS6UCrs+QnMDIDw2xCAqB6Coi63vPgm22DC7GvVqYDqnn
JNImT+cCPa5ANH2pCzXem6T6suVNEgi1yR1LqjQwtLRcmgGwTLElCuXZlyIc3cd1
455SxMDd4qT+tMkNqaCCAfOrtab5/dUNMfP3vce0KP+YwzibUojwwQHndPWlcrFZ
kJvpw7KDM5d6anhgFiJlCPtKERiGt6f04pXBkoeEIpYBpq+omSssfFkt/SW/ylo9
9vHqSW7gG7LjXSyVzzDOlwrq/1RbMKABwSBFQg+4dnLzLj6BwhIKzKhCFHxHLTiE
WZyAcXJ4iZtcg6jCkXuWStykmg0ouQw5MQVyye7GX1B+ji6obJMc+rjFnpWlCEKa
YlAAmC74/KLCKdjKcRXislO+lUNCdr1NCCUlUryAjpV1YNSVIxoxLOGehymAYyJn
+Dfhl/vK1/gph2O0NaymG0rKGo61oSz9meEPIjG6mqAKlDDxX+NC3hdZ0S0xjNJW
a4hAv26xrLZxVfJscVNdauhvqUrmMX/PxbhJLpm+PlDc+S7CBN4reJ15NBs+xDG/
hN0BtkdtChyXlAFdJcUBf23SduYh6erkFmakCOjnTdm2kHudQxgrAYb5SYuWlzhC
g8r/uexVqm5qDWCwQdyHkWDmRGJTnC1UPOeKbOsVEXxV6fzGL5KvdgqALVBZDQhF
q/SU+iUP0LwqH3EAx5yHEz78svF/EarOIsMP6jfmCYBQNzsHNIgBD+bRtZJmThxV
tTXD5BxdlyS2LnNBeU/XwNt7qXEits4Mv7+WSvtv9ZVDXTu4shrWoXcuEvlmApYw
yrZMGhdTvXCTPcFyHG9utQCba9JcjnRQB/4wTaLusLEtACo9sVOuDsx/IfOeCxjK
vPPSeSmh7NRlVCUL0Ab7wSaknYmdjrVUYkdfmbssjtF8dbIKUBkBTEF/6rUYXhEs
JxHWeHs94yHYwVUW5RVnzlVc8Hca1i9InFhrYQY/Szd3GuSL3aibffO8dVTtxZrp
vOCk9jB/J2Klyl1OhYzk+GUkfoacTOwyp9RRT0mMPkknugFWbudO2fLC2KBYRsmU
Q2vqck969qN9fLQVt20L1T6XIjpN9p8wYze54/OCHfLSeCY6rzLo7pHo2aNb6eeV
zbbJBCSvMgM98QVNsSr5h6RWNZr6TYv5zLJ5yrXFc+rw6EtZbY+SKPpjveIUhYrC
fxoZaFGJmg24eoZTwR0L8CB6Rw+x7CPYMK6/MVPr+hBkM1Ve45vqqjDEOQMqpj2p
bJDQhky7kRoUMu3uVV73SDhtTF6bLFL6u886/abGl73sb3t6ZhB+PVSuXWndsejD
RZiw+FOwDxbtgbKii6qMKCEkwcjAfpq7KFW6g/msrhPtRYOCVB8FJwsVacPecCez
5n3YxekRebMIBvw2F6QWvztVzeiRIVacaGrQp2GGpXaiNs6+Dpai9ARjNDLpIG2U
Vr1OH5l1IQCD970FQf2HnvVxPPRBrrd89LD5C1J9iZR/YBkzGq8tR4HG9HqadW0d
ifxylg1RuozVfkJc4lswGPSK6hvQ/qMaQF7ljA9fE87rzMoj7d4FaIA3DT+s3UmN
2mAqTG4aZeNVd1VYdPgquT1CGsw+RRXbp6zdw+vSb9mEKZHpSVGtRWV+1IqwhbRr
bHv0pz8Z8aBHGloaixF/FpnJYK6hqFMGiAPxWphbK497j5wPGbC94ypjiLZI8slL
fb9ANCfDYFbNfF2UPA/COtEuEeyKdw1NV87uJJpXQrVKUQYUky7i0xZoZ7DYqz7Y
2NlzIWBpFyd2YXEBAg7m6c5QhHF2etp6+fHlYCMKEG+arQiS4QXXXjfFBs5rQDbr
oaPyv/CJF9NnxjMuia7SRnWawBxg0qQXTRrdhDbNRJ/dLS469LaKgU9nyNjj0sVG
wvB8BJRBe6j+Nsu/GYQMIrbyyXPolHVbgGrd5aRi1nnp7LsH0ZLNwtJAqNXaVOi1
sS/756fe1cCcqF18uTW3M6OYIpUu7mTrOjombTVKmmUNKGeWIwOxmpawuJWa0zBw
pqTmfMpcGRSlZ/MePUC9zYbb2uZyFldUiwYKT+QMT1/EqleYjvPS4FqogyADvQZg
eDXOqjoFqxj4hVGItkHxrh2eYOTWQzHFSGd2CP+eLqqYRi6kNeVzDfgomm5CiWoK
5IRq4gV/L5srazpDyAPYp6gD5ZRjvXSV3rR4Tucz51PO7W6U9y564g/QI9AX3b5c
pUHxxtDxGHUgDu8v1N0e2nE/aWTlPzJKjL2SrwZWawX/Ui6N6XqbW6ZqFD4ZQpAR
HxrysTvTDWeMIlz6urJ/bjaNshzBcx47BuaglC1+e7cIMMOkds3/vgkN9pfsL6bY
lEiRZIjk4NscmXrSidrpdPGntLTDPz9voBN17fyxhOO3ULsbDHr4bPF0JanczkqJ
/FyHXSaGHw+busyWojrLbYASA0BvkXLckgadrw+s1m2ckdReVr4b+YiRX7eYLk/U
l3u6vQFPekFOQain9SnFc36cvRAmVVoLK48WbgKut22nyHrErIT7IKCaGNiOsZEU
+acnra4NZsk01JJ3PL6E13l9crPxol61vMXXYvFl3r1QfupDTD0Eem1zIuaZ5jCH
7NJcVk7/0vGCMrOH72yrCdd8LecJ8N4bJvon2KnJK0L1mSzLMWh2618hwOkUVg60
nGmnSy4qiRxGtx9coNPWFoqCIJgeXRJJL9g3b3Ycy8nhp0Drv+Toe3askGs5NkOb
nEC86lNCao6fPSHyo6z2rbbpMYCRrwfHwhut3FlUOME+hUyzG6MceaU4npatdPOp
DXSkM9gXCtP27dqc25VcCroVlDAipdKAiwspqpB1UPfAhrCAMC7nkSBYnwMUjd0z
fot/9eeMJXjmQOhFkdbA9iMhHU+e1eAocq6xJdxPYdhAUUjpibdGtX5RiZOim/IR
jZNwuy7Fos4fNHk5x75gABUemdl9HtB8RdP0mQKJ4h4c1PnHQ8I5tPg/No0C84qr
k9oETOSsaSZotFwXUPKF+WiYVyI/nE1uaFKCksIWgtrLoEJ/Dwc3hp8vbQ+0/P0b
0EhayQBqeJlMfab7UqmkZfmqdn9yHRKPylHwZLgdXp54Wvtc5J9p4z1WSeKyhnfh
NC6GIn80pUeIwA+SP/MVHINf87HwEhcRxIVxH/pgOReaqhukToDhC+HUtkWXOG5z
/0C0PS1TBEboX+GoeJCNQ+LkVFjAYkff5IFwN6Q1XpxIIaybuOvtTDT6OyNGIeyy
Y1zEGuKuCUqrjbVuzbVdHwMkaZAklIqbAWn0KLvPqie895+aWJ2g1RU2n179F1JE
TINj+XY9dYES4lwGTMdRBtXT1RN5VFzO7ihMMAxn+X4rltyvswgKpjLRNtp41V/z
xVyxyGih7A91jM+VS0O/nnwayVazgzvzN6N1tIazgt/WU5kjL4UoCei7rUmM7Nuz
w+ZUBrFI0oXJ3/0wHRVyXpAU9+S1N7Lm79eD5xmyCql3T0a74Y2Vt1CbEuA9aBnn
lZucuNni4xneDdhr81azlN9WImgccSZzoUUeeZl6uAW0DeeCpIM2jdS2xaWMtEuV
dR+h0eaHZB4ho8Nawp/aFzmq2+i7tihzhSwEsgQ2az+rc5I/5zyOY/gmtRpd/MzR
TYGD14TVT7NQfWUuRWxxbWbuY9us/GygB2SkBhd1cmcR7RKCb7IxfMbNh8mYubhY
JhtSmZ1UvH7K0MwRm3DKOqCj2rsP16Z/gDrAA0HePuWviy5jPvkPznmFg1MgFpS8
xXHhcQI7Utl+TJadb9jShnkZELNbKFEJFUP3k57vbrDwDcdZctWZohw+WcAkDh1L
JhabjBGUht9eMvm4EjiZECQTSp4y2AfxFKpEld0r7PrFuY5iN7mOFNyHWoddb5wO
oeH8T2dR0Hv5v8dJu9nW3gQjtwXpu+8F+fqpyvzB4597J2BNzVZLK2j9FC65OYac
JVN7G01UCLma9AvDfYDXZK7PcU6G1GuKjbgwPYOEiKTlXR4lzkIEoPJXSx6Adql3
Blsfo+h+p4ck8Iix7cMGtkVRm9NjPo2KWGK1DM4ptwaU36z/a/r0o9QZGVd79IQL
aW3tIjBBx8iJ8128MDn3MlZ0AOOyi9bznMiZIXhAdQ78OsgUjpK2mPHPD3RPJq1N
ArQ4npxMOsfcU8dGr8Iqlhh6REscW7gmetxOBYeUKrz6W6pL2tlGx5Cb0lFNzDho
AA1sYdOUd7X0hua0fPt2fPJe4eMVdhRDqwbsGwJAPpbaCCRc98KIqK5pDTiA518S
yTwbJEiKNw4NyVrmpSIWoW77/WTsdL36HG1ADW+W3uJoJ3pTIuAfM7BhCg4IYwfa
OsKW23YH2tcE+DEjThKxaCJO0uVB8R3SD5NhrQ9U/qB8TfyEt3cEP1kW83vhWqEM
HEApZUB0TPjVE3IKHQF7j7STobTmivTgbbcrVVmiL4ZBNkbXHcaX4cS8g9Te61Do
MBSYVzGn4T7TdMiGp/etDS1wwLPKohrqdrioMOVD/W023U0w53rMZuDSxa34UMO8
SuRf6W60b7YspOJobVpLl7+tPut8G8E2rDn0dcVZHJgUXfx2ubLKNln1BAiJ4CfU
sQmwtas/DXaVR87M2WmCTvlGMYWDaWz0FKwSsxS8x0jOj5dQHnOWo781CE3W8HXe
gxkIdFwSOFDx8Cpud3Og/a/sQhG1At6oo1rMpVFmhS7+bl7VTh355lHdZ1ja+vNG
HLTS6zEkYt9XIAJSE5BXspUH9g244HooeOcuAsaJSUXQyklAlQZHh76ObyhaE0rz
tCfUbqHoYa1x3Laz0dgtcFp55X0/cwVf6aGR9ShJS52IjLNasQjrDtjsoaWX0jAg
UCN5o/gdHmm4NL7wWnOXyMcFJrn394wH1d4zcGhVJBtJLiQqv3srmbupRmsMtEkT
vKZiLwNtVOQP/32rtAz3Tb4aPf2LpGKmqA/4+9Vwvksnveqh7aXs1dj72sVEigRL
0xdKtZe4ljO+FpygFKYx+5sBAj3Aad+bs/kqbM4SDacv+YOdzpgru62ub8hhDX5n
8ckxhqUx7p4ftz71ZygmT1R6JFg4UBAyUbwSAKl1cjnuaqlzrikcDWvp/sCbWNBr
px7DCubkQWtcyUE1rRiaeoEKT6AiFdGQ8GNKCCf1WRokio+DOfTFwNZnsZivd6MJ
mkop4uFuKHM89mfjxgb7x9Uk3DcfIzQSB2GmLrZn71ePoUq02qEM/4BnhVBWIZQ4
iq0ifYvGQfq8uyT+7ZlTI0OYTUrtMFOqACdX6bHeJpnquS1Hgp1FB3wwIJ8jskFl
3Lmh6fgUVCgiEqhPzIoO0lAA62I4KczB335KT5eppVVU2EaspiSGoZnLRkA9IBiJ
MXdPzoXvRnA6sP24cvXOqbhso7RdemIJZHjP3RBmhH0aGxLuhbtfOz4CVk4pXCmQ
aA3fYzJDkDP7xxaJz3CuNV2AHxojK01mdLqBGuPMh/WuJzVUCMPK36yDc7IhcjNN
Z5v0LAjWvh4J2tRU0WVTUdMY6Z6eiMtTjxkLRtP+5+RkFw6AGxsOQvXsbLo4Ol4S
eamVyEcCosd7QbF+qEwsC5JT6iYTCKrr3VUTyCvCEvA0HMHDXY4t3CwhHrsn6PlC
nvEahFGuCBKO1nhNgvB3unwWOjp+Qr1usm7wuZ+WQhc3D8BuoeWUDNUWO2B1bCxR
zVjkJJs9BuV2j1wBuHwq1q8sIZKHltCvhvEdsbHZh3hL9jHutQJWUFrJCsCMIs9G
9qZF1CZ7J1dBT44ZoSOI9v6/VIcQl0qt5tAdMsg2/0gXG9WfQOzCfpHq0qu5oaWh
TwyWIWoHsv5eI/l4kTKAh+FeZbaYObpgNLGdT71+58KEcdIrUHJpUxKGm7fJE4Ou
1kDBotp7WMQV6wZlLHh3zbQ0kQPvRMBGkfPQ6dcmySKV/B5dneooAoFW2fTnc3vN
LFf9iQGnAtl86fToQemO7dF2zqSVqQuPnX3CFzIV5o2UbigGnF0DWgxTQCRKPY3U
0yvUKkaiKZyLsB7N8zHCs5x92/Sli2P/RvB/rfQNlwriGWizte3+gYAlHOeqjBQs
iKRK3R8mPaFpgqXAtyfsVwDxPIXEXHIN7PCWR6AUNjrMET8IZqsdBawuzktwUzd3
MWEtq7jHqlK9oWk++3O3lv4TgTrK4LMGaRx+LcApdSBhDYwO+i/jIfwrx53a0c9l
zvWUH/K/963D5Eu9i4742ErPRKLBpjrrzG7wbkMX6Mc4reEqWcUQ3UDbIMRWMWGJ
58i9/bCbmw3kx58i0pNcCLRkaPU12meezCTU+7X7W3SbWRU4+vS5dMlTpX6pNt1l
+/j3AO7M3GhCnMBKiGH5Scg7RclsojcjWuhgsI5H6dcMw7E4XKuYXYb1l3ClYKgn
jAfj7XosdV3DkR9ImQKovvHgtgN7y6L0lX6/JOTu+V63UqjQCkKEHt9zYhJxUO+z
C29ErIw4uF5vmCzy+lYbsakl1PleScwVsCRnAEdxIZeLR0Y1MkDkB53ZNNU9E8jC
Wo4S/KNAkEO9932IHSALWI5RiNPeiZ5EMTNASCU6jQ1TDyXx4dsY4g7B5wvZCS/B
rHcGG82diYnf5Vy1W3suTYBWS85d42rOFTfT2HGWWNgOnWBnCQp8HPRIc6epcdor
U+AsaMy7lV3bH9X+qtb1LGv6GekaYPwC7Bu+WuUE8IsDMccYtB7/7b45k+pPQdeQ
ckoXrAywBlJlFrzj6nL4HOHERS1o/HoXbciaY4oThM3Fv2ngc1hYbfPTucUyvFvT
X4fbO0IxmbmB2DtUvI98Y06sXPahGElmmQBDCFhQlltzi2KvN+R4sv0ReJD18BHc
GUBJL/RxfOPbVrsdoWbsilwxS2EMGzFEhkdBu/Zl4QoPAx27/N1LAh2gUpXsSX7+
P5101zzcISlkgUjqKy7DE+O3aVzCnya4NOVyrP7eE7vTNt8wUoYgMx2McyrNGtZe
kx4IFulC/saQqYbxO/63tKKnxFKCYe0s/fLuPk2DYbvYWiC7tzZpevW8eHZXoDRJ
JGh4zM/uZ1i9BvGnHjT/UwH73aWJ7twQAF4WAJSCFBJiU/Pk6gJ15cyE/hIQzr9k
qGYdfQSMsgWSsbd4rPetr9LKAHXxcgIbf7HU55s/sOEQ298sYRHxl0hXf+vCViGg
LolmIZm+9bPbqBnzv0oAgwhfq+KLTEwg3d0cNEnpku1VrfZZI6jaB//G7HJRHOY1
kYMOwjF+xpL1jp3rCVx2pmUzEHsv3wvzAjchvKYQ+5YB9gBvQqxw3+vMirBPoZ92
T7VKeK66iE0zwXupDtv7tt0Cz6Hu6AZ+9vGAOoNiya4NQ1yRloLw2Himr2MkpqX2
w2Jh9T3wnvsx650QyD1j03O/R1u0sk/LMLPSV1S9Qla7sdASTKan5X6LS4QyEw54
a6ZM5+23MAAJoL0KwSAlzSdABLbQoFwrvJVpl8359b0irDmuYsqeyfc010RKpoJV
01m/CKTutsQqtZFyH9Thr/zVfDVqaYUyGHnwg3w3LZ3ZQn5VAjEeKQBKr8zZZnlZ
VHMCEpgB3owxBko5nhfnOqzWxuXXN5ARHxUNOtx8/tFQAEEn92yyxcEkGCb/bf4E
444AWjKDfg6YVKDlFIDqHkBkgJMjr0ubWNdPfWOSrWUQXQK5lxzPUJq3s/d/B82x
Zl+cmprVHEoqARC0OByO95t5XEg7wCfaglv/ywhGhuqxT1DHAhrhW89/cU69tiEd
AdlNm95eS7Foba6tnpAhB87xQumaBCQt+2jU5OhWPJqQNayozWjIcI8B2c0sT2f/
gjECO7wfoHhUwf7QUlY88J/wlHtoqemWvxnc1rjJepjpwc1IvQwjM6L3irU99LHG
Xjb4rmql3Ms5eiwKTM0/zvAbcin4i3o8p0AjabrpFKLj/3lGamtIpYjwmniCE7Bv
aMdTvCwIwiabxFz//ipqDGeONcYzq6x4iVmapdaglK6b/G3XmkQEpshWsq1fkQRC
3K0v+wkOEekvhQ5+H887yLevj+xjygqNbwycU6AlTLCQBi4J8BYEu8b3pxpikAdz
FosYrqHrjFEC7bs0ZUOU1rsUeyAThJ7Kl7XwOUx4109FFUHKOeYhqFaPsgiVYEaj
7FzZwxencwsaOJdwHY7kGtasBsq3DzLo1tPLkYSQY1cDSzfLkZYtodFHLJA5a7Ur
oucIKeDHQrhhwxRLQOdCSKhQxLughHu3LlED7aHkCmJ33xEDzWTF3hDfgFhKfF3p
ghOjZnmqkBnzi4SQwzBFelVHLFX6gaPgf7X/exyhk8LGTZ3AdmDTvGZwRbwhDHQB
xR/d0Lcc0EeeTmUnzEx2nbsiDV0bT7XtRckg3Xr9bnZZGm5z1csk/bbxC/QQe90m
TRdAXbNQPc412zaKoJFFB3eIc7DaL9RD8ysCUP3WKp+ahxJah+0U2PcCIqXMDUBB
no4aDr8WGYR5dT93AvGXCoNihZwjYEdpDgbbdKeWwaUNrCC7/dDehuzdFGJGiGlT
NiY9tvmmEyi+PAE3127Inm16h78o8aws8ujFdSfVv/dvdFAWCIZQ7aW60GD/gfkK
BYKva6sn00h1iTy1HwFcybNj8V3vXHp0SXdJRccBgGwFAKqe94Wh1GLaEgYef4tj
jRUzuK/wM+Wc4GSEP8ZtUrKzILolH0h+sYoJ4LYBQhjuJ+Z4SumlbaZnkIxYexwW
zLg40EfeR5/ronJBaDMXki1AKid9tKE7igSM10BqSZhahJbCEZuiVvmp1035Fsme
fAqAK7YyVdbPpr+hCGV4QVTwoyVNdUwlZrKpLimFhVoflv8fX51isnrG2yi0oIMB
f4LqfSXNpZUjBB5W75jk24m9Kl8kU8cJQxs0TICo14B9Ld2CNWoTdhPs3r3cj03t
wCQAYwXQsMQ6PIbhvFgAZytDG2u4qyG7Cz2l1d0zsOf9yKpcrf+PmWGBAnPFExXF
YNvs7ahpdrf8NIN3uWuyXdME+UtrqAGMTwOPI1qe2//J8GQ6Uq1i3ofYZ0NQg4QZ
LIPXbWyOvL6gkgDUdOM3RaL0Q1jI7laJiqt/vJMtKROiwkKNhg9f5HC5tmCCFiH4
IHX4kzLb0UuA2NMzy9SVO7jypBdjvlih2+Ghtl8oA9ZQnr0NCkbfBIWhxYIYeZBf
/WeABVJWiWraZE/WMsNt6OdvzQccE4jXkmO2qdWCDrP+SjdZp17EZJWgyiGa01Tp
jYxf8LyPCM7TIZUEvLaRuotWjUFIa6T5PkwWNs9Po/1RA3y0CLy9U2Ol9RbSUhLO
+R1YWjc/P3IsUX4tww6UDMnqOQuBzEf5L1ZsecFaAB2lGE6l06EcK4aqERr5wkOj
1uiD3y1jjZbdGt6wsMSEiLrj9vYTVwTKoqaqMRZP6hDhCW7pjUqbIJLTDd8xArdP
hCfzp3HeY/snk1xkuRkBauMqRolOzWtzESY/4eLNHfAwbr4kdX288Zy8AyaIHl9X
wKcr4mNTUsTFpH5kYzdQJU5KzcbO4cJhovncdeJ9gLFJ7/9UwlFyID5nANziPfKQ
GNzpB1uEtjVOBodFJ3+xPjR7XxotV97zvl2c9irFKVy14gFjqhUzhgcGMltkugHf
sYOVvVMICOCrbCkwRc1Mr+xFIcVYykSVRsCrVqhvxIxUEaMTDx/0wxbrivOLb5H7
bi/w7UgAbgaihhVDNnZWap9fa49Ol6kweERIgRbzVMwnw3bVUvG3RFOjPpT44i3y
zS5A/xzSTy/OQdysvy1DQHi6fg4EA9wfj9HAi/w1cpQnURH/AdwB9qwVKD2klFXm
QOD9oOhPj7CaV0njK3MO/9qLEdkscCJKclxgltb6S/UGLclPKwYQY0jIylmMQ5mh
VsmXeEvk37lVbvBGyVCbR+afsLOKkfdyacQ0V6aSrRT1vTC2qu0nMF2yJDNMJAxn
RBOeBYbp0J1mEdhS+88Xng8Ln/XSIR318mMzG6h4wUCqG3sH17iVIvQSKLBmG3cI
69d4Y8tJ0LMDqAlh9xICD1P1AACDlHvQO9Q41BSciyEhopLfCxrRXptYkYh5iIcP
hNTfuK63ZPKThE5CYomrsRLAQudyG82rkLG+hkkwEJL0NgLUsgzRRnTBNchHDo8J
nCmNmytih4CPTQB39wJ0y2+9L96t58g0wp8jsSzQcX3ERQmaR5P+apigASOeyXCy
S/UudyYTUs6qRf9B2DpGkdLPR0a37UfRXFTJkmDZwhHRioxQs+JWQUIhRB9DeBkq
M2Cxli+OT8Ebd77f4yJMNmmX0Ipiqz+yMJsGkyAycMPkCEa9A82QiSGyrqzKcjHV
BrImJ4a0IzDs8gsyWguAV5xR4nNbhscK7OuIxRr9AOE10I/kR+dM8lOjAGMrHS8Z
daOie8+FOJiKYFWfiFM/fgh09IgVY6IzQvHyVlmixmXX5JK3sCqGB1XdxMV/oP+W
TK/uyesC7T3qwzMgVnaoJvicTMiMcNDs+ohLqJpnGCg4LOcr3Wn6mhi4v/iRXnc1
+PxPgd2NxQEhkbyi7JYnQDBoz1qH6HTOFbwxjdvmVUApb4jkPaVshGlx/9RpeBBU
Q2WhVpDQERJUh+SjxQzzlWuSO810IIo5PkR/725EAlYq1WX16x0cEOSZnMzfvuQQ
0Js63/HQz2QfQX1k236t6oTQphwJFUIaKf/ImQQskfOqLz8YUEIoSZoaiGesoUEp
ZRXnxGv3pp2KdZFrxUIPg1S4eyAEXcS8SZ83q9XHUmEsnQfIPzJiwHYEVXE34J4+
m7+mZF58IMffgMC/B9O2W5R0FnT6L9mKUiUT4SQLDqQ/3wzH2qY8VZ2CBFoTMy76
hamKheqVod8XvaGJfQDN53qsXX8soEPawoqSQ5AbePCDL41n61ZKOSMbUrgdXsKO
kpBsk+Wj+Y3dR8vDNqnHdEiRbIgYDyA/nqqTVt6RJXukvXjjz+wMo6kYLQz9mJnb
nr1jxzBh3YvZKfYR/UnB66WdgnHRYL3EznIPeleLh0PnOsX2TBv0g5IB0myj7p9u
IfwstCJaYZW1rUzO+Rh9VDQrmHib1J+Nza+hWj4kBR26xkOaBhjgOgAUg8vaWRpB
VwIiuRa8+rzWaqJvXNrKYCmsCqIIUoyjIma7JLJV1wPdckUIleQZWktEx/K/EqdO
srf46yWhnR12QtNGH1G5i1J/p1NIsML6mlcSBp3DH6K0J13GOcP9dyHlwbYfP0cj
fwJVHimtPVt37TDaKTeOM9fHCDwZ8CU+P4Obl6ih7Hdj1pqf8UbWrUtzYoHD2UjD
hEOVp+7WW1F5Y+GXBzXCtJyQ656wzcwS5DgoYyg/B2DlnMB7OSO7AE/9HwQbaMHF
liC7Imwhp+TSfjLnZm0T8nEZPWBdrYkl4y4DDRpP0dOjMJqr5i+PMIP8CKYU0PRG
yNmerQGgAt+rx4gcRoPSJzJynkJgr1Uy31v5a8F5HIR9yKxN6AjDqzffsrYBBJkk
ck8HiwbEO3DEeydNi1NffOyukcWct58eB75OrFH078unrV0f1VAcOg5cEhGvk0lH
/UTY+r3tb7u4WKCLQxQ7//TAquczZ8A6tpL2RDh9/0p+TAimHNLV7eVs7WAH5T3P
h5yEaekjxWg7wGeKRBaF7RW4/LdMIkrPsLLkxomyySqawnB1uglI2kPz4cSUNJBE
tKxIkMfuyyqWnaSM75dmkN5LhP+QJXjx+vRlho7JBfg60vL9Db6wDpFKKsLLlJgg
DJncppJOo+iivJQK7B906yPD6T7q9K7yNDD+VqpYy39nfJV14IU/TQIfWwmRM9Af
fYcAFbAO3ye6cIZeMmi8R1Z95CLgjjDF9T2p9/OesaRKFuETKREzvUE5voTwBx56
wrtzPx43yyI32xqTwS/IC0FpnPkTPRU4xWrXG4NdlPE7c9mH/orXg1TfS2e1vV/A
Sitq/IPBjrR6kciNuQAYxuwO2MKwfZf6W6euhxAecPDN6F6RtQGntm+z3NGTFYid
vr1FvzAyqcAFIXW5ixvMUXLz+CVk/gR++qG0n6uut6IT/exXeZ67mY4o0KoIuoO8
8uDsZdBf8AqcccPixIg3kXQzrAr8gUSv3K0ctl5EHJKwclVhnTsuU+yMo+KAfZ86
Qb2GT6sLV2kfJC/AgDgaASMguODK7e7ngZEuMrOiSjti/uvDSK/0NTTSt+uXMTmv
bWnOqA+AZM7l58Q4rY6TnS56Gr8308M2HC1jvkZvPN+b4LW8mxDKPjazvAv/Ff9B
1HEzOr/QtGtcT8jcXNQ75tIGBi4h8t1aPzFS7C8C+yReaM+zw4xSQpMqAbdbWNpb
XusakbHb7FI61cF75v/pwvW0lLJkfYdO8rb8A4WxFXfPTdLZtOSKZ5LUTBvvH2Kv
pNJhvU1UCWEqUW7HKuY3roNuZQyaGU/R4oXsOhg22W68/BnTMO/z13PZVReStIMO
iUw7HvaZ9ghOOYvL2Xl4NqvzgjdLcivTxtyfxBCD4vzg3gEuXM8W6Xs9/EnrWGKK
SglUiLPxf4zphzYjShD05mDq+WbmaHwdJtrswR+U+WB6V9VrirSg229alg3YFsrO
HvfvbDQmJtVF/wyKVeDiSxqo3MQ/duVcaNsEFhipfsQHPjDFQhNgVnuj2dBW0G4A
NAhc4VJxKPJh/zSxuFoxwsZ8otehxndxsS+8et0qrNV/Mf9RpzaVi1bVJbi9WbT6
hV79Let6f1LEsmEZEYuBUJqy3ENhNu827OsR98Qwh48NetR4sl8+nIafXM0w6ffA
6RHcict84tjretrW6HF4mbdZg8EZ0BrFgpJGy+YmdXlPyg6LduGlQ7ZVluRSOm5e
JjdwUg85RbjrtfdQDZ27sast6RMmICcFQcRVZHp7ShZ0luAFHScVx+AipB148zU/
Ldoh37B4W1dJGWmhxqxwR3J7g8gKImxeJh7DKhQAeMX/ud6WXJ06OB9zHgvNfRn2
pHrF3/RGULkNZ1VleDx9amuuXY2ba4tNTVJXCSz39tgfzH2XI6DcCuz2XKpIk99i
4r+86ddCHkByOBeCeJQDXYeV6a43Z1FshwFwxm49sYYSflj15h8Cje9O7CAQDHPO
ZroVnpf7b+nreeyfiEHd9tpRy+1LwvYYIZnnOeuYIW5TzUsputzm0cb0Ry+MNMGL
IQkfl4dNezb+OWoHPGUDqjEyKyA+BbOakHyOKUkGBH4SNyrpNi3bio7DcSSOUffY
iGj4dRO5x3it8GAZgPMD1DeW5OldhVB7veuP9RIGi06L2uqAC0eLdwhSaGi4ff+7
aS3kPPmokE4q1oURNt/dNspe4yIEeYol4nL7w2BGCqj2vaxDMZygssvScKoocqXu
dPoJf7zciHqs4Y/0pjMeB9eiQzT2rtxmmFHXCWlvt/a0W4+ADi25ZwJqz4Z55MkU
ZwihIlMojOdh65AZNt0g/yUKEsOpebOL6/zsqZLLJ0lzL+a7v4SiMPEP7jxxA4NO
T/hwV8Ew70VckvDldlkorAZVodvcgKRAwhrpWyXzSiVwXg2UUVEjg8KEr5v3UVRR
uvpGjMyPE6UIoW26weGHsp8NbHmd9Cg1m1jidJkEd5ft48HaS+xlolYWrYWGTCEf
4pe7KiiQt1pQ6oYvw38fxcWawdrz8eDXwvaXH8khbpO6b3vVJJ/1tyuNVA3OpbL7
Q9fZ5Q8cAMxzThyoWh20eNxpbMM1eDCKJF5d+3vBHNAzGxPT0wSzgP+JugFRYJ2z
NLoel4JVxlF/r3Ho8lG1ZLw720rRg2EAPGzLYC2r69N1ilzSuXsq/OdVWC8SIdtO
L52TJtX0jW0lj7HqXW59jgQ87y4H+D6RGFfjVziHYlrTLWAnuT0Fk5DtRrwFaHXL
dPFN1Doi3JpJWwnRBtSr0N5Y22WnT1R+Vi0b/w/wK9k6sAsE37d7qzErIH4Q+S1b
FxYwzlUqs18QataMEsFk+u579ocQxBYT1F69FxgZt1paCWzAo0mIS53mjB4UhzKh
+wtwnLo61YYBdjmF5VXZkNsWHJuwUK9Gv2xUFs071zoU+kwa0CtDEmcFLr/2iU+n
+VUcguHYt8/lFVkazPJmeBhlHyI54ZuupwHGB1A6w4Ujb3cfjZEr/ngEcNbm8mSz
4uXsO9sK5NZ1lLEXJldI+ip2BsS79BxGy3uSPSxuKTdZD/Be4zifyG9vVjvgYVuX
hf+9QRsOONZO5NyWCMX1EoRjbASTn6PlZ2zOpcSoIzrzFYHh5jr4fptrCSBTCGbJ
7NQF5APw5/qGXIA4zbZFDe5jPESj62GxwuD9QwQ8QjMnAiLSiiVdTXGUxUnSKZWS
TL5kn8A4YLvaFn3QNH65L6Lx6e7f2fO7yQAN9nwm/ycZoD6xbNbAznykCBMVS6Zr
u6/XlLHotGZbSp0ZkvkBeGwpJVPC88Y5IKarckokpjF4ykIm2whbmHof2FLJsJ9e
CRaaEsZ0H/ik+OSNMVlE/tTr5B8ay7OKWXAzfPuG4APs2YOo4UhGEza1sUuYWsC2
4F5VZn5bMt6mdVZB2Syvsr+f2qUJh4cwZxHpwwsv0v2iP6O8Jcz5LlDaovCQY5B8
SBP/g+1uU0KJR2OnH6EmolRzoKzJ6OSuOx35J1qaN9sx6mPyZTxHH+9gX+ZNRvqB
/LvGnx67arFn9hZ8Bm/iYwM2pB3WtkqwAadR1x92gEPVxyyYHp837bMVWa/RW+3e
nFkR+RO/dw4m4JA17Bzs72c2GksNE3WpPCvXEio6xflj/MzN57S6LjPVqrHHMi3O
75QBGa6c5L/1uGnmMpPTJ1bs8OY+F2/Wh1en5mPYla2vrgwx22aJHDtDA4r/Q5Oz
2Rbw+h9yBnpG0NthwCwPU5wjzbp6C9V6SYkR7jEFJZyOXKH4hs8Zvea8fymvggRK
Hd6/5l00a//B8XKpBG6f6mp+DGO1370rmEe1MIRvHwYjcG+/xjg+jwkYNjiBrVDI
qOdrOalvnWY0rcV+oF66MflI6BrVFOYJNlLLTSpN5ILkWYeRTCl1CFbrlMK4Inph
shRirn5oRx7fEsalfKb+q02Vm5cJKGwKbRiql7hB9PvPd8hrTadsrIb9jZ7uqEQV
aMoxp2fRUGpDfDfXNIz2RJYiaJSBjToBTHEa8huROJ6E5mSXzOx4CET5M6/K0srB
mGwQoR+vkTCuM8pN2Xtnbi9KVz9alg90fCf9/hOiltHoXt6betowPsTa3coJPwaK
AQ2U0SgyVq5pmG3aDjZVcZ/D0CV0Jwp1HrTOGSw5M5SGD1Psf2d3RMPCV8A7eUfk
qI/teapP2df0pWgOOWf5CBgiL/5nI/qGG7cmdnyrp6c3tynnW22bob8y0tfK5Rea
OLfhpd3U5CYqP/91CVb24jdUEotybxKgUp972hjdU9Y2kwIgB90pxKpq+bu8NvdM
7b7+Y7Hg7ap7VLcMLJVbO/dz5NsoZLo+ZqgNLv8rNtKQchGe8wCtH5V7TlwmIHEt
VWPtLunh8q4rVWdOwU1fSs3IagL8/VC5zDQEYDPvmdpHdOkNP6adr21fzK7MqvyU
eFFlKNkTSugOyVyEYs+AarvBk0uLBvZwoHbi6U5g6thGZBGxSsvVRwRHWZe55yhR
nkdAIMmzFfEYaZXd5qYCntLIFpK9g7SJdI9lXlH+U45utniS9xvA3Fj1JqqHGfk+
NXpIRmvw7kGC/uMJa2sFv8qMdttmgNUXDIBRFoKZgGbPyHhO2W6k/xVroTPkVqTg
IVWzLVySHWae0GeVZMUUiDUUQ3GqfRnRQzcYs2TT5GgaZur3Yu4XyemWRMaAohiB
/VKZUzfJEHRV9XNMqD77lksNUaXjq4xexIRuhIZ8FT48wHEqOR3PO1+uiBPnV53O
sSGF/YntMOSaGpkk7vFWByLLP69TvTGdtX4b/ygLzSZERe9W8q/goBQQ7sVU1PEL
aXykgABdX1GodBL7HJ+1Ovy5+hu/2Mj+T+hA0ieWj+m0U1NgW1YW7yFqbdN28PMD
bmQ6wCr73Z3dnDA1x+M32KHWLqoFGm3YF+W/MQ0Kn1BVVKcqcrTDe0sdSnKO2S39
p6BQcit68Y9PZoVXBzolWs5ZgS26RxX6w6VrthyxlYkWIR3Hfs5gTv7rkrRDadcy
AgI2U0br0iOJO8vNm1uei5uZVka00+XUS18MRj5Z+rA+J6E1umg5ehXpRzXUscBz
bnfocBJxrufMKi9KsihgPDKJ1pMqCLZC+p6gUm6RZ5Z8bKAoNj/BVFwt+Ut6XsDP
KsSj/GygLkOnF+g3420lJ2cqzce1v1yedi3cetEElp3xz+WpKYIPkjQDlcYWJTft
AxV5gI6vxa4idtTZ9eDP62afNAEkBYIc8otUoCwpSOM8duE7my2dxy08zSYWI+4b
ohS+Ec06oLpPvwVkYjbX1pGh5ZuoWRaqOXXEo4wNA80hUSg+oBNGhpUB6XvUTj0P
hHiWzHhIuy0LtGYCPGBB0accHprtZGVBCIrEn0C6rYZgyTuJWoptaclj0Hc/lkHa
y8OhcTvoB0/cmJyLAVp/bY/ENqL20I5W1UqwbDM27PxuCyyCCmzailTqo8sokiim
MWwzppt1SzyfWvm0z+UJsHWS/8skInu5ftT1UNoCaRepouyAsN66ttRzYNs1zSY1
J8ghpDj8TgEX34cVmKD4+SgOiNQHynPReHIxVYoO1D6kt6gUFgV/QSz9Wv8t5aY3
fjl2MHgqt0zue5busChFROiYxgUU8tv/xS6dT+cAokEWFKhKYKmarz5KoKbmWlld
15lmgLKSgNzuFzJMa+n7GlZhMKbe4sjNvye3fzapoWIvBDLL5IHJMiTNwLkJkDbC
NDJehDf7Qlzjx5DU2Kg7FqlxGKpDOCA+P/h6+2Yh3O7R1hKZIv8jzYcZsn9dz09l
gy1gouuyQGC07KxVzUDYJaxCuwkCNCNLnjp9IYKuatpFMMkoetrD8Pws7qRqKptk
SldYhvTdNa+isMnSUdtuun6X2gv69fPsPhqxpuOF4p8qHvx3pNCbnw29T5Qg/Goh
b80gKEANmP85XmGHbUBp/STc90bq10jtrRQgE2qBaNovsuSZ5qBKzjKoF0Ddf5Pp
bleNjuHWgf+7A2Gg7y/1VV7EEi9djgeYR4q+uNj35ttSGPzMqQ+hAn/V06B8IYLS
Cjk38AajBmvwZq4utzF/ZUEZ556fpFoYrUTGee6qyrLs+J5D1qXQBQjpEi3INBWj
1xP/2lS1aWK1pyO+s4BPMm4vh/QwcSeElmpfpn4y87gx23v+aMXvgIB6xzxVnKMS
sCF5HE+Tbhg1IFKSBDpcMbosMzJnNg/GXMK77bNlfJdqNGjZtjXlPmllOoUDAFIW
fD4dc3OVq+hsN7BbJqFkVfZrL2AqLoxvpaLwkrVguQh+cpOjhbB9sMiLY+0/wBCy
Tb6voptWsu8xSPqMoqQPEA3nLazUsdDDcJiwnzj9/btbh/Exu1R2Jy6QL9B4VjoW
8jxiTi6O70IzEmcvLm5mhjpl4NoooHFZlXCijfz3DS7rUr08syeOpcbDxWmrz60s
12Tv1VQmB/5ATwOZbuRQUKgNpGUeK6qnUTmIoCjT72r6QC6lxMCURpwkqO/7jaa3
XzKfyt9Bybacfw38f1gGZAdCM0t2j3hjw42BA35UvJSKPN+f8UHNItU4vgzNJSvd
8ZRn+/+8UMmv+R0NSkj0gkYC+6U4Ik6VsexwSEcHl6CpmtlwyqOegNwxEBxvlfi2
SENYa7sl6Y/U7F8jZDnnlYlJ7lmKlfdlm6vFZoZoo4UfqJpYRvdKoYKjInRyr/kl
YElEUg2YxVbF1NR0DDZrvq7tqXKcrAv3MG4TOtv2DD0uGb+WH4qBn2LWdO+sdud6
cKT+vTGFFfoVxLcWVCKvcXxG4eir8Su6nWUMkoSC/3LyNRBIkk/zOtTOHT1WonZB
o9tiNAiX7/0/X3IoE8Qocx4aYi3Q4SLB1tXqkW1aZSu0CKMQ5TbqoGDOz+IPcTIN
ORnMC44cEd0ft0gR42FHeLTm9ubcgPkkBOPNkMBAOX/ySnsbYDGRt8GysnUzM+7t
B+KHsfEOv1wRRpV4lDiHkukOnDZ5to6jS7bgOH+rEozQXA778h4S+OxXVzHp/pgg
FeXlhyUY+vJX5At56WlGPgH0iQKDT0yVBaHulQLb0Fsk4X76mQyGDfViwh/kS7u+
Qnor/amYAbrDrdRaQYji8vnn05RzMIR2t3PophaIfAud28GqyBb5QSRc2pQr7cTw
VIInMH+c1mDvklZzFQX20phGNUxYtKVdQWEYg/6Y5VtZIODebtv/tcsyRSuygo7O
Mar5lQFXedWU+cRmk4xOpNmXXLQ6nGmwDcysjcFbsDxk4Ippgd4531StV0d8fuI4
xgJGwm6l01dYWzDup3ZM+yovZp21oLzgYp986+tG0TB9qfhQBILSl4BKWCRJGtsG
dv5lIBSeyZmAqAX1LCQkUviSacA5xWfIS29KWaLxlO2/M+PqoLTrEQSEOr1RZVJa
/5J9LNNrLsh6L/itD1bIGvJmGZoJtWQEx/DgvLSwFgCozy98+ugv9mUtPqqfIZ+2
ebd9XMTNzvaVnsGP0Xe0N2z64It6Vo7vb1a481xMv07gewxhd6SrbhQy5bnRTMqQ
tCh/KDfz9+HjkrvQmYvpWch01OZ4LWA7ZjbnZtfemLjE+wf8WOyjWgsVUfbrt1gq
/MtcL7SDs+Zz73Qq/aPg7sZtXIsM6VRwtrR5PUJe6p0rpN1zZDySpATT1+Ck+9Mz
q0p9mgf07nu+HO1AyVyoLvQRznbAeJ3TCs61LviJRQ/qQGEY+joC9vCD3oX2E1KR
5K1XGtSXoTyszl4x/6iQszK4FxEmjDZY8ql0CLPLkZNKU86lp1jlboP8Z1qQyr/t
s31wtnRZ9MFC4TWAbiIPlHI+QighEwyevLnQYn5/bbSzQ6cd85kilPIsFVQRJsLU
hWOHuGCYODrDEsWuaFOCqU/4Qzau8Q2OxI6hiH06LmEDVP3bR4FXgfy1X9jmNdP9
5ySTxpGc6cSRPmztnLzaUCuyb//Jw2VOCfYCF8zF21tBnQ1u7anjE7WkFoffwbuB
0EdReEsE93GR7hKuoDRvLSEuYPHz423PdsV1nqirY+bkq//QQ2+LIEpU8XTuDuko
QU+oPRee//V8V45AvVFZf4zgMJWJAfIQ5+bYa9LWKkCkUYSfEXTAOmvg7WTa/zfK
a9RQoS0HewybqMcK1VKcKeyePsm+BQPMxgOVJCKRBF+cAyUZqw2fWbkRglhwAw8G
HY9eBtXxliC6Gpf0a3nbwefk67DLO8KWeOBDKUnpU+1RACRpuw8gYzLWEYyvMvgf
/psNRjPBJeycSUx5ZbOiDSS4iiH9DS+KcPb/yPtZ5EWnY+2AAbgCWbJ3pSa1jsfq
YRlDlkDcKHr4UEyFZwAVFhLbQAbwC60d35Tr4JZa7SuCgMVuAUiP2sQnaAwUA8vk
6MNpFHFs1H/baiN6CDrqhCF+BiP5DaTOnVSCzkB2vPotGAxxb2B4VPtPDy5x0Aoe
DZvtI7W2YLPsyvqHxwe1KePTuAcSk6hJl4+KySbho3FfAKJZzrCGCs0WiAlEgwSj
CnXyCSeaPDE4urPzR1YIpcj4XWhQlJmvqUg5kSNIMSpHg703V4+RdJ9BsNNet8oZ
HMFzrDtQwATX8KyRuhNk5UoTwt4z09VK7M/pxGb8MGrerMlUKpTFaZ1myHJlMVsr
13bGWf/LNzsa7dHYAM3Hu9CZfEtn5Ir5eYJRsYbfwEmtrfIYuWdn6TLWLZwf0xvX
+e8EkhrThKbjNZB0CPCpxmORITtlMNwqOz+aejCMqwuIv6ZTFtAc98HLlijbQ/4C
nq1yT/dNSeVPpMetGcDyIVRLHbX66wBVt3hJgVriaG1kHOge0YXWF9uJF75CUsVf
5XASvOej9Q154tAjLhjmB2SJo6Kj+5JWNrjbpUBJi+5IB/VYOt7H5QtfTzcUDRBL
f4PLK1pHnqvn+sPegDOnfYP9EuLoWLaSwPtHmB4tiHw+WV0SzarTYbv4fh9d+tIS
6qO6uom1hIGL5zYF8oK7ZejtF4B+tw5ysjSumnbGCT4YfVqEzdw2/rn6F1CcK/zX
Fx7EQiQ5Cd0mM9KjMhAMVY1b+oAaP2s1lM0Wtrn6XBOvYj77eb8Qx27Urp7cqDmH
M6eJYQV3T5vDJRxl4Dt9vtG6wr+BwoscDhLP7nvhj/LsjTFSSPBrM9xx6m2C36Zz
C4rvbackOEOsIEYFNErqP2+sJ4E5U4GG71nRMzFdUbg0LeXsTT4ocaU5C2YkXGix
BQ0g3Z99+k/oPOCrj3rCgdDBp4JpAJn91p3DGTAIxAOnJngA7PF7MhmIaMV9KnAP
qq/FlL2WZxOmoZmUgIsXlU004yw5wLdBq/zX06SHmbEljf+IyCLQby/9YqehQCZ8
oUlP9FmANqteXT0fkJZLGozJn9v2VkjGCQ2ELgg6b0IUJk9dNMYXtxEscJ3pXynj
FiOuczQALURw9MbPGADax3zNz9mpIxuzoAwNJE6QUe2klSZffJvbqUhNrT0COWsp
/4OGFSugGep4VJ1JIGdQuKUeQseKYqK3ar3hKBAys9Mqkub9Ne3+UWpz1NCOhL5x
nFQlKIMnbkLta5oBM14LSh1c2WRrASF9jAlHCW76zal9Es48Ym19KQT66Tb2I4o5
Lw2P7bKT6MLcoMB7D8YJ+v6M/IuvDhufjpdJ6TpV5GsfB+WdZbzMDd96CWIsv1o3
jh8oMzO0LdNMseBGM4JkmZCjIkezEzbg3Ry+zavY8ZcW2s43mqDcDoHEdqh0NILI
NtKfc1+R9ZnE1vLGwPQlVTUN0mxrnFL6OORikB718NPwjRB5guUjmLAqJdrRzvY7
53nHXTSa53ELxk/uYbFJHBDUiafRZ71f5N/ZWhF0PYbWle6fr3CiNPQnvdeweJdO
fetUwKHfGvj3AYKq96eLwSPAweHhF9pmxjtXNmE86VMrbjNAfyImRls9QBtiA7UI
tXGCuRqH0lRjLNx/+SYdiU/UQn2/0edeBHg9G4PSvZ5/d1IFBkbnvKpIiFViXoTf
0tY4elmDUa0o8jdxFmYQJ+StV6yNHHVKQVT30Vun1JDW4IX/bfAvTO3Irw/uC8bB
7AmU4BwlmQjTlEkDdIsMXYWBHH121TVFlix8nlgIMPEnX/JtfsfEpaHKIdCXrMcl
91I7DnUTI9QxocjG3Q0UMkrG/YCvBO3d1K85nrm5rcCmj/kobDlZgflks+tblJIk
wuOfikjZ3DvvAaG59GdGVPp5Ss+4qS57wkykKTcPv/oSAqkB4QVd3H4kKN8WEYTx
6CrqBP4VnCFG4d6GSRbjrygU4ivDZCnYc5APPBEpzMXAGz9pSkWKd9f1W2YuAne+
UeZReBFhsOwvyF854rinzi3p0IwgiymJL16AhQzI0T6deYuknka10PA2yfkoQB7L
cohKfkj2a0r16LksvVsOHKy+gHVJzgHtgiT5VjEqQYBtCxS+WvjV2TIQe+lfIJDv
TvkOIaqqghg3ScZy5aVeM1EIvmZnCSQ2Te+7bGiyM8UCcE1RCPExZdYI3Cg4mIfU
cyL85VmYJk5BozQX9Vx9Ku6qpbWSk7uwV+syuuxWYj4cBqVblEDhNwWkg1dlzVO0
pfks7Iz9k+CsmAqlqhXo3YdOA1dNPIls1mLaSwoBqC6M8zhy5gfdRtlMY85H9Gtf
rxfWdKJ4yjXRpf0TiFLvJ2ceDY2cq/+K1UXeyYYpvvpQSmkVtPKPaq5BRMJsMzJp
jNYGawVBpyOfBxjYguLJZ+Wd+EzRX4/RXEqTTcx9UFyI80Mbg/k1zIOcdx3Qqbff
199SQDj0OQh6AEaTVCSDi8PFeL3xbkLDuAPFCgV58cs6UIyvNMIV8yZvwisgCmtT
rZiLpLPK9I+x11hJ0Sx2NIqGht9oPY09XMBbDfuDtQ8eWahJMhNeR6ZTTWFDWXkn
SyU2bpAaXzDs8EZDGgBMpOwruRC8VMKIPERmOcBj4Tjlxuko8ba5JeDMm+yPMfWO
8cSJhcLB42jozvdIgZg17iemE6+uGJ4cCXqooKgqGzxvR1ynMJuKHYRvsNOktKha
BNwvXpTlLoe4hBeSMXuxyRaqxmHz47bvbzpbdD7DBtaivYglvk0w0cpFIdZLpWDT
54KTfKo5GfVSrZlpztYcTec0/r9UJNx9JoycC63593otlGSaPFE2p8U/hzasJf8o
KovsevKxzRvKGCwCzk8I21XAcJYh1XPHPEb9JGuVODgTGJPzD3yD/HpFj3fA8yse
AQEfZcxkaRk+pyLR2yj2MyF+b+lwOBxhATbpvpWW6xszPgHj+KbbfjiV5TSBVXdQ
okRPjeLjb7OKE462ZKX/ID5aaL9kVyiEVFqARPhQCArt0/he26fUEM7Gz7FuOGkD
YiK7Euxy0VLWIpp/MDdhW4b9uJe5D+CElVw7k/g2U0B7YQvLV9FZw00pe5ua3HOd
JpAcuRPrBm25nsi5qx5cdNxIojdYeVcfSLEa1ddtyGIqMGLTzFt777DleLIdsBww
1KMh6WBmRXQxhxYQdxNkSWj34knXZjQ7o++4PVxhdixrDN/8Qa0JY9nN58ZbsK3o
nDuCI+sURODind+ctgBwWsbefLsn/qnOUxNm4ZqERP7GJxzTuQzfHgKagZRTEU/n
C0WsuyG4jfcRiuXmG1gLoPvko6fxtl2nkGu1KJrBtCG5wHRM+YngRKjlQcfGFpwV
bDsS9D3jclrwwLfr4KXZAG6wmAN3ZmP6raWO1IVXquIsYGWOQVOu5R168LEvTEsX
g1A3Q+/YWekYJSyg7IsSZLtqSBz/KnL3QTfMg6a7CHdjWj8B+XSW9y/vUbth6m1n
Slaf2jzdq5lYdN4v2HaLzOEMhojO6LT6UFXjptmfSecRhiJ6YEtU6uy0MuQM+p1g
PsfwX3ssq0Bp74+t52t2zsBYK6BeMbDa9HAPjFHEB8TBCsWr3k3PZ1zgssltgJZz
NgH8MIVjWVyff5Jr7FBa49oFPAtQ35xSCVmefvnUQRq6sUcQxsmEgkSYMB0as9aA
mlojyv0V9FyEooye5fZF9DZfmqInZ3kAX3x1NpLC+yEaAVZD9X6rMYxsT/uSIu1m
JyXrL3HJqvi8FBwzkyZ4DkGwnEFtbcG8cLkkUiy4D/ByHrR81Fnrg9oVswZ+jHQ0
Im6KHV7UWHcDAEbe5GRbqjm8VFKefl9ByyWVm2vTuxcKQ4ZNgYBbWelgSReF1UOP
G2tm2+TUc3XUi1pCpZOrgTc/aJXf9ISN01i0odtpHexG15s1tdDQd1F7gUx2LuHq
H5v7IKTdKGhyQFQBs8euPeVqeYDOBIl8ss4h8t5tyyn5ykVbysX0U2SdZEN2pXgL
V25AmA9gg07/UmB1j0a8NJeD0W5xGThwiHgNbx1ivYo7ZQkLSt3Y95b7+VrfPbSX
pm4RfrdTgMCYNUDtcsZL98mbcynLgzyCEMCGEPw7q5mIxsKlYXzcLZ2lDN0/fZ4K
otvsZCFkZOMi4QHsUgsFQEfRnUgvM7QsV7ymAcj6OeMVz+c2p+hEI1/8hcYpZmV+
30iNn5KME/uE24G6s3NxvfXoGYlgaloXL/OZakxV5WesZMmNqnwZadbAIRT21sn5
LVNVRvtz+CyFrTn8Sm4rU8b2XxCBBUBpNJltUsltstB70GWQRII08ne8bQaRWSHw
F/DbNnWZZGI8em3Y59x57G1n6UxXn3e6KQDtKcV+UV0kxRcPo9tWZjbeTSV5sLoB
zV9HmiPpfm2htiUTFCackcaOTSHoCvYf4EvLuP4PyauWZ9aXCkwH30h8KlpOiCXZ
vHP0Ala8fQzTM1MUAhAeggRSRw86ROdkgAMKfqeiBFjPknQyQZszYpaJE54J9BuK
XmHYeUra1NkOLaGxNCN9tfJRpOetbTbEVx5eYg4rOgeoRSJqDiAVcbFpcHxgNQCx
ZoX+XsXwbOm25UjV5O5/dPesnx0OwpKSz/1xsZKaUCw+52esMa9NJp251qV9X/TE
6iqOjR4wzDJcsexVhOBdI+Uck6v5NXDMoTnRGNZuFGuezrhvkDMbQVOT0xk3w9bC
78cOA6uSVwZsrPFgtot9lv8jXZ/Iy5HCjiq3W7RfqoNAcHDoW3zauq6wW2nAK2Cc
n+En7lhJcrOOLgfoIV+mrO6uavPxFnJrse9Z07W7V68dtZh8bDkP1OaVMjNldPCh
KJIznFnfF0RRY0mXUtTWX1X/xUoLSaa2+nfaxHwk6KIOSNdwgbke/2RR8FZ2k5GL
khaA984BjV5UVrvjlLa5zwohsJFWsw4YY6xFF3YP1pfrfRSGVIxyDdoi/TkGkUWx
YGJI2dXu+KaMK+jXwXUUh1LEXj9A1/fs+axjrnrw0D5MvpOgBlUSJTTLsTipthDK
efWXiLOff4O3Z+Je0KpZ7skyEQBWa/xXRgRAaEI8mHcp01rz8gkoFi0FBqzRET8s
M4anl+OQARAsbtMkQB0+lpqcWgHaMpXp5XnGrDZVvCGv7Gm+um6TEunUMljZhf6z
kcQyfze9Vv5bev/QA5dSG3lFlHMf/8MnPG3j3p/fJGX0H6H2oRGCKmcpo2vlLyCo
f9DBtSn50kLNK7/5gNeCu44lsuYLgDvS6TcOKsqmRoGPjvlueWWiIbVdzU/q/LVH
dbaxi6ZH2YjuYXmQKDfgk0MyTRjkCRLAVKuKaNkUn858pUAzAyefVI//yX7zLu4c
7jtQo0Frv4EL7MNGCghBP8FjwOkNLRhnENyzAi+Vpnevjbn+D7Sh9fXQlPWSnvUP
ppT13mRRVsbsXtxhzd1CdJKyRcV/gPESzYO4quRaVrFJuD6S3dEZiOypTvfFpgIu
r7JUNWkh34Vb+j45fVzdEwZC/zDEtDmIwDWZcrT1X08oqExl+XsNjY320I3ktG9I
U5dQm7axF0CJK/TX1v/t9/Bf1vx2D6jpRSR5SSgrbc1veePLah9SH32UNlcFWTR5
1EFegJbIj2wN+nL1lwxKrLQFESeTY+U92w0sQeA9KRwHBRAhGWHQCasBX9lCoECi
S0wZVLab+oOL54wxBN2sWKBgBGJeMtXxnrHFOwlRpe6siM5PDc1b1U/fq3eBaM4F
cpIAX5dq4X+IOyJolWWv6cguTm+vG/21FmgZFdgnQqH8i2dSi2whcz50y51c8Qeb
9s4Zo8zXhdZnax4NxXUp8YAGTT7cJQILwnooDj7gjqA3FCtbTFQI8XqmkZqHKkVg
OVX+ZJ3po3rkzkvU61+XVaBsakiAnp1qpFVv10Nrrn+nAliP6qu7ZMFpsa+b6sJ/
WQLgl45zI3rra60+1Iob4D23eNSMRNR+NMiyL0bX6YDWlnN0P8LtsUQ0V4EffDbN
ciDV2qoCb5nslGDNlE0eZa1B1CoX9CCvkLnibKuWM8wrLpSxQ08ycMrXe9dVmI9a
aUfbW7a5m/0iE4Nbd4oLR2nUxQlZSrUwREJHqKs8rjFsoI5Rra07g4lqoFdfPmUp
PkF+lr+l+o8/TaLUjeq+9c1nOmV7HwEdtj27aEBcB48PrZ3gcUiUT4T34CmbHEQf
hZWTvNkr/PPOeCd7NsDsZ9tstc0bSX5cTh0/IMYRR+4owbhVLGZzjeRJU7uRKw/u
06UmmuB6OMu0CCvRQJSk7oYvdAhwqcTiNx3h0CXS4WsCRS6gflMYMeXB6wJtTuAa
ZYBFxU6X/ayy4fyMq+5zOIeTgxhzigqg3liCNf+KLzxHdQAdZjFfgjI+zHyEiY0v
pIpySf59SUxXdfYXRep3USdKYxiIEAjaB2D2IA2kLmuBC+fF9MUx5iul7yJBIV8s
urLbNYTSxiVk+c72L8UgDOR5lx/TM7BH2SIrIbBDIoTF+KjfCW+QOUUGQfCXlDgF
q4yTUQWHQTuwGrmHPY/OepCKk/QWBuudOtaezhzLuvbkVVSLRiZsOJKDYPf1zc/0
6zphXcicZd4xwrZSCctxhDjZFhr5JeTyJpsc8mYRmnqs8C31vHZLgi3bDPYkYc6c
G3aoxcbAAJhtuHz5TiN8bFHrTeZ6cItF9F1R3yC2SlC3/GSX0nNLp7st1sdYoOoS
Sii5KXzrcNfT04dTA9ANVDhq3qvtfOsPbdKMNsVylil6EJ/Ak+XB4xjSSWPZCj5v
Ko3zmBYnrCHy8/CTgStOu5sUKrq+Z2cRp2RAlddWOxjxC4o/xDXwdx9r5f+jfk3U
ezy7N8Uf3EdSm3GIhpA9djTcjcWhYM7LGaqC2QONhvZGWdiFxco5BKM8qPk4/IGj
1eqlhtpWa8hpPlZm3LkUb1RdNvwRPJkVn5sD+7aPn33HXEcryhQGYdT0I889EbtT
yUqJyvttIaVwnoIzIugzup7K2X4BnjYL7zlcJomY2RHYYmSWw7nmDtIq1sKsTQNc
ix++LIJPbZZ/8R13Fa5pZPq+eRDvKTmiBN1JSj4r0wrXumzmyWtbNH/ADW6oHxqx
Mo5rsQD+MtX0heUSlN8fAqyP0whTrjqtHr5FcdXkP8m/eTrcu6S4F7V6hXs0yV4c
qphth6Rmqfbrrtjw9kx4UXt2EXJkB6o4tPAyzP71J3n+1pNNGG9z+fPfXqL35CNO
khKeDqIh9C6PauK4+pIYlMzx5A6frJlUIutidiilpO8LpfoRjSI31bKKJHLYqnxh
oRN6iBfTrVOja7/ohNlRCCrfOrA3PRRNtPPWwh+yNPIhUC4pIZug4sUa37EbYOPV
9D7QYAXGqHisfEj3S9LseittklXkMkmylTPV7rlKz+0sWvNic5bQenHOERQotai3
UsXDduH3RG5eHhilhNTLAMlPJY3pLFULnNvEJBrvTCPTEQVwKiBOxTTq8GDcw3HL
FS3rCAHY/wyFGH4ah8nCxIuCK/UhvUNlLvGo3SLdoX5pLUXMuASTliGCnxWN17Yx
SiRSABkpzQ2pyJB3O7KaqQUg4I7k3YG+jKgLjs/MT/Hp0mJtfvsHOUSCesNIlniF
VnsvvPtx2Af/xLPr8nZQM5r3qaunzKcnantjZyqdJueFUCvAMz6dYj9Q6tqZOcCx
uJFBMXgunKEiPwsANIHFjHKe5k9+cfwwjykRrBaKxV5355U+Z8fltfd4nupHzFzs
4LeimxG2X8+OgtNyeCnrPL5O3q+H15h7dp/9ZU5eS0zrKQWB5oAXt63nnFmfPplV
Qp30UWtTHsbqoyGLbtt/kYVq4gfr0t41ukWHokf94WuMM+ASPODSGUsJqIljp8Vm
Y4SzJhLsB9dvxfH39oD1wfDasRisFfycwB7iSKucavKu6+deQT5FFCK8Rjwec8fE
vBhv2nFPYWcRfasmtiodPvEZYC70FnrwHX2PyJU6v0xVKcS868AAn6V0l3eVPvPL
ZTinxzhcANYXbOA2bWugYNfC/YbM/8GGSIQ7XKtr4HBuTutd45P1b1hGKozRPI3U
gYevTFuc0BL6VrCNtmxqqd/OGfsXKjXvciv+2dH/bOh499w+UisHsnFcsNCk/SXR
vLHuwDQOXEqBHD+XvyjN0hyujKzcXPJsrnxSR5HT7ExEjgAvA5g59Pixu18rGTKJ
u0PlnVw3C0aLOoaXZDTp4qn1puj3HZEYuifhkFzsSKTRLDlL50db3ac3qJsLF0mV
MCAVMw2M9tTEo04FvvyIU2xebC1w9OGovRHoCbmAev8H0EYYDPiZZ2DBdS9NwH3f
rwFlwBq1rl1fhHIbA8ONrLrS5etSAhr2+LWmLj4HlWV5b21c0INJHtoeAixrjmaU
9zVdhdCH8e85DVlgpxJKcEbAHQGGsHDm2+qo84hgXtCjnLH3JmmNm8nXFBSZNzPD
6GYl+QCfDY9iLiUU7I8DABBO7To23y+NFGhy4ncQ62VpQ12oRwa/a3mUsk5csgbN
KjWBY6eIuNAGYwxTN0RG0Bnvf9fN/oy/UHkPMA1LtRBEx7RkuVu/WjToDC38BxEo
3Lm4ENx3L9EGaSR/NEXUg36xu5Ug98A52Egg0LRskAiwtYfkc23A99+kYw1xMRHJ
twYjiS2oJP8WTITL8JU66KqsWiw2rJPyUZ2anXS2bm2pRf8vTc6iscxBJqke3Ctk
buMJprSr4NfMU2W/tfeWyDsQq55hMkxps4xRuITw5hOcdeOmAlNN7RIC4D3o1lGW
S2/rheQOkBPbkYApxJFQ+XUUq1tmlqgGJCPwx1HTvT9qFUHMXZbPg8ryOUOGA+IE
/b7AmSW6y3LOfJe7ZSnHHgQt5qqcpuqHYYWgvfvggMAaoQY1/0EEzeEv4r59o0Lv
5KEYTGev+dIGzCZOgnpjpn0Oba+YIu7MIr+RlicCVbkjMFElLnloKEgx0gLJEVql
M4Roc/f863vpaVkNRMotgIamXk9gtPNBzbMWQ6T9E1Vg1v4BO+aQGLLHoT8FsFJ8
cHz6UGUDH0Es9VrdyUNrvYgXrL/sZ5tc1I+qbdAsNIcKcc3MU5lYdKnBucZPymml
TyMp6nfFH1ojOXyv4AIhQ3KTYAYz4WnSTRN/dGURMXmlj/+0GZCmYT6/UbHgPd4+
t7nF/png6Duidj/bgiuOIxDV9iRK9pPskL4Jec/jUXEDMdDw8dqHjQ4aNr8i8Jr0
7MY9t3qFdxUyHkc7InA4kqwIgzQctSgA5CjcAQs9LDK03vUGdT/k4LKLVlPDl5VS
tbKCXUlMioF9Q9QsKAMW1t/EmTwLpEJjw5amtLNkaah6jjkWH1Fr2bHeG/hBaCyW
2z/q3b9JE0FSbL833M43bxEwB5fHCTWfLNhvoNV1xud020jh1JvufI1mHuEGCrRL
9auuFDryX2uY4BX/zPR41oZ3XgBStpo0yinRVfUhenlLD0KzhcEYa+Z9w23jKzTV
Vz83RQ2ddGCoo9d7lVpCpK0GtaEl8awd9bXgmhyFnRMKYd1KEsEA5VeMTZUvoXg+
q3L5Oy+cz3tm27/yb/J5c94TwdVCiDeIANhnJgLJWLoeNzMfoO1cWYYQmpGTL7Qr
JEqwP44sZ1skL88YXzOTQtkzs3XUlTk+FEr3f5XP5ySYP3Jw/6AC9CQWhdRtqRdM
onuggW0QJ2AzYyg6a1/5L2bcdr4XnjFFhfo7cVnF8A5KW+TZp0CiiIHOI3l7oRXy
YM3yH3ccEUSBJyoTixdAgBeu4nAm48i/UHVdfL95lXVKbRa7Bv9m80IHb/zGxbqC
5RXNmFeDeV9215cx50ClkKADPZjx5AgOaOYJS+J2GiQK8WLqNH5HhSTL4UoG3i+q
LNJXnJ7FM7yqGi4TffYcKyGMZCq/1qAZ2DaXhnkae2/q25t2xtQ7aCgNgSUIhEn3
C4TMkZVvcaVyJZMZKkOMQ0myCTthEvFoblDqhrPSQquI6LG+7saLNEkX7x3DdwS/
5zrw4VKlToS4WmZ/Zirzr9msrPu+TTPgBRtrY9rbadcKsosoeniXOKUZm0j23u61
OImT9jYOqh9wiOwhwjskzLKOdpT+mXu6UXJRP9YOOpeq5EckshrUR3+Tx7s/pjOU
9hI0Hdmdy3g8BkaE84QbJpGMVPzwiSRdjTlJVrz/9qJj/zNExgTLgXTSdlctXNW1
6l8rr46tMNLJXcAEKOH/9JVWxEYf6nEsdbbuiuoTHlAJ1Y/yE4GDgr9eErTiV3W/
0AdjJSa0NWF/gSECj2ZcBIh+IcHW7k7aPzIA7WIGZ2P7OAOIt6/LZCovAC/p1C2u
URsVVAIrUe8Ggoqijf3hFxnGBfB4ecalLd+IrWtDnOlLriyDJbJK8fJRgsqfEffK
AhSKMtu1Wf0VxGRR5Yskawu4Qj7dR/5v2+CLR6apDr7yHXeS+6R63H9wU1JUdOkT
9ACAAt8oa7UNUrnnN/N14b/VBs1Y9MWh6GFiVWVcWubZHhFMaUPBSXyTXHNLNvcZ
FGepxB16fOhVJ1XyTrLscFkQh5CH4krSFkzBt7Jkrx6NDI7lS3pcGE/aJYHqVCxn
3ZEt8YM1bbGVof0dqQxWYOqnpnKUTgjKGH+DQ7N9i6rNZf1XRbEXP103/NhL3RSR
//xxNPHfnhkcT5SnfFyOaGBb6iog2pVi45VosewKDVyarINgW6PX8QgHQUbTDe91
hWWOJSxLYxNHmwEe5i2kpq+VNysIvXGW5f6eI1rvarumPWLhiYZ9QSHvD2LDQvN4
bQjQhCOjF62+/odfbpfzIZCR1tj2FKJ8gWctgqlywaVsliWxVJZcKeyWubefjc+8
iBLbAIeVoirsIatZU/4iKveWKxr3mR+ZqGfqnTuNfqHVbv5y3C9Yk4qqhQhPjy6v
45yaKpOJA5+uen7RfsaHLqHXv4uPDcox/DZpBQ0ahWVc2tbyqal5efqnYi4mF63L
aUe0pkfjtzXm8snptRDjYK2hmH6q4OC6Dwq7rq1llCyx552FDBCYRiAgkME5cSck
BadhDPWrY0z+lXytt+8tjpQgqlvqBq3l4nJNSa0MOjs7/JGRUj79J25GrWjPxBOr
IlCFtmip41tmViBHS8sK8j3z6EYcpQFpD5X6hKQoFjR/5WfSkU2G7N1PZrENq5Ot
XEjIhCYnBDaUGsrFjnb0umpfw2tIOjaAZr2WephhutOJCRNt0f+Xp0Lg3JiS1vXr
ch9Kq90AZ9X50mFnIE9WpWGjqpLsPQ5IW6ud60GBmlM/OU2HyCYQkgPLHAjYPwjg
+SJ/9NSJ2065uUKomqc4KisRGPYKwq3EU/bju/KqP3J6ee4Qd4yJMEmOZSfiVdXe
Zf2skL2Ibvwhz7Ow3w/FyWSAhgRedG2KWqgVDYz65Nbu/6LgheUPjKywIujbxca/
1fmiDZjsRXQPEmFHF2zHax9LSnvg0lQwThuu6FyRphGJ5N/ny9N5VHWoTf7O2XbH
ek8TZIyHjxnl0Hl3x5xmnrXmOhxZwVi/5Ft5i+uhz0QCvMCqxB7Gz1xxWxHkyBz+
ulRRjzg4p027uYqO2bugxMJHVhVeWrJct1OjzXdhkTsLgXl2Usg983Yt8KKZc66d
QBkEwi8FxQjec7zbQAaE8WWTWns7liTiaz7UA8QiunBkZQp874wcOrVXpeCl7zNS
+uAhDJayZbeuebZd4xFyVRRZ/N3r9fy/YsV0QFuA9OZA5QSLj8zg8FLFDqajp0d9
aUOEoxjzjTOlTRnTYKZSPNg62Wd35JwV9LNq6J7LybJ/N+ZWDaSZMNWiWUQxhW0N
jRv+jt69Jn74Xo3ly2OEajOkh/kY7sXEw42li4i+EJK08wkvk5chHOtnYavdvNZa
Wr6GeWnPKomOAKRXZGMlOaNQlySLLOx97D8Ky4NVnbPcsFo0cHLzqzQS8bFjBpSh
eo6fFG7M6AbYmFvfCocmoBRgryMeE8vyJWg5OQihT4Za4Ib2oihyv2gz7zJ/qifg
zXQcR9Fmx8cPLl0+EaqJSu3QbMu2bUKWu6rP/gazzEgslpmkYnvb0UtykgJbTLJb
HoxcFtssynAXGy8GEYoHfBncHrrXqOikJLl87/Sw2WfpzbqzY0tqmUYfq1ykqFVt
mFHOlFFa2C6m99jLDvj9vfy/bgCvpCxAjr17uzpICs+TEK5Rj14DNvlItBTAc8lf
QBRDfpV5oObzZKTwyQ0V7+pkRrJd6o4XpOsynCgnS0y0Xh/jPL7tSH04hnCDGssG
xvK1ywOF3VP33t9IidsG/M0kdt4fo6FU5ihWM2Wz070pD0itm4gCQnp07LWXe+lt
tfv5/pKhWu2LAcq851fENqHfgw6nQJdIp9PRWg94TabVI/vnv7G/eGBe84rwEKS8
t+aI+tRgJDnwXlOtzHSTYEiR5e0fV/MmmV45JgoVG7v8NgKaLhv7avJqavTbq4u+
x44DgJNU/5TxCirJgFoPhwAekeqStNb6ExcQ1g9L+RBkq4QmSZufJW3mekCWk7B8
dvo4FY8+pJrymE52J8IsN8dALHzbmZB7N4NyccbjXZGJmaWZ0CpL9azHpYTEQpqF
4gOn4tBZaySx1Rq4MRC4TNzqzemIoh1FN4MMBdQr3GwI1z3iKWNSzwlitjaaM3qR
VQzRmiVlyk2dsEtpEmrWhGSM2UakBBoxtL6dFMJbhIPeIcByOLmT7ZVaGzqwQAFf
4fZURznK6azGvawavPbMwyf9NTUtpfB0S5vRSebGWftbbtzuSJyVUnR60JAYLPGh
g7d/vhnE1P6qWnjigGR1TE+coqCpIhHLLXXWkIQqO1V35W4/h+E6h5NyYMQ9jyL9
LCOIFD3UCgVJ+Clgm8/ylml6dgVTfln5h2WhKKoBJ3hRyzXc64fvvMJU50Fv//Gq
kH0Tx6EJGNJ4/7kE6oCggX9jTAuM5FdaLEHZ0fdBhN5xgfiFOZVZNcXuygOqwgM5
6b5ndLA92YE/NYUkpBoHWJK+e2y7ySvh9eThsSen41Gh3XspDle7HCMbUkASFlpl
S/0+Oae2RKk9+ErosLGdF+SFIlErXvfEVYuP5FFFdvoetCVmMODYuXj9UW1nziKj
okr/CJTopaazXBa4Gcjl4aYetyxWlgSXEBIy5Qq7x0flj4lVdB4Pgd0wOxEnDTgV
ilxeg4FO6T50Wf977gRG0etBt/nmiYYwiUIsc9nKM9bnknuEFcA0mMF7ZCzv0oUA
HaMt4ZBCX9JzSrk8qKY1t7NKemsLAboifhY78cNizAYZR6P7ACu0RMPtLeefdXmV
VqD4vBHNAHPpSOPjZLF+lygL1Xyq4+9WF9jpvvySJBLct+DmUZ3X7uajmupC0gVP
/IDkWYUCrMY324ZwQ/aCFVkTyWQgSd8QmJUXsvxGKqBpZXoySBLgB1X6vkUaKQy8
dUbxNidMqaA8daBUUWcqCT5hY5BORqsDZ9UVFo5criYoMFFkLOXiroD0afHreA8T
Yo2SElBtXnS57gqxlvfK7scUoLcmoF6a1GC55FMCvpXpfbTdNIVgiPctAdNopvrR
g/UGzKdzHniE+QQ56r42wya0fTyr94WPdIgDLYNssJUVim5wvdNLl39yMw6GvOpI
awIaV2erd+fSMgg63QEbQTov+tOwuHA9TxcoaKC1kBDszbWXDI6ibgm4PdvDblrG
uuyb3Wz/+qGsIj1U75otA6BUZVHk9nHw5Nu/BxD5HkFxW07gSNjg7BNFTp7oN4jT
i0x7/szZdEFZKaZYHkIt9YCojVgx6Xd/+4+Ms6w3lWyiamNl3fYDYfIfhBdRhdj/
DlgVIj29AO3pNwepVvSUcTYLCE3gQJ36djNdK26CepYLw7/VxqJUfRSj8GRSRYF6
CHNy1+HY8T9NjL/i3o7mk7TVLx+808tAZf9pw6Nla7zMZIHV4gWk1zcty1FGnrsq
2iqZKRXhLOxx6K67yDUQ3e+VH/C/R3a/AE6c63L8EIgD4lx/Y3E1Y+8KP2zOr4nk
HI1JUk/Y+NvSkToR12u8El0Ci7osmk8fvVTGEZvZZfHlaYBlFAHTOd8VNn/s/wch
WYrsnK2OTQjTfcD+GvXH5Gm7VgOOL2yEZzOrII0jdV85lY2HtYlDbTwCOxbgnQ80
ZIHTmfzOZ8m141lEONyAhDv76CqfgfOGddCYdGz4RuCpklNuQql9Ihs5AdKiSCJT
HhhhuLrnv5nlPVIwY6sKZDHpH+Awf6qzBHDDg6PmJdU7xCbRoq2/pFtG50q86nXn
r25Dz5ZBKMJpltkwYZZydp10httHUvdPR0N8nOppKEO/uQ7RtO/tAY9sgAlfD35h
UbkeSguKeHATEvdaQyRb8jE2QSuyLbscokhxmUiuvHeaf2MkPlH5SJcl8pa1uCXT
yDL0cJinwfA2nWqSCR3aUH49QlNL6Scta4pV7r22dQKZwZh68fM+xPexkMbG7Jvq
emHBIJ2mqbeTHFDcz/GW2DdCnOeqzTQpqQ3yN/cO5cyIa4lxbTyZdj0r9nBArccp
cgdAZSEccTp5OBlcRDKCdHi0F2slYJ+kiOT6XGRk5+5oQ9euR2N2KixkG6ZGbUGe
OUwbRSGMzpwf3ujZUXuImFgtxRVzd5Gf/KCk1Xof1WvuqAzAwXvk5v4tObjnKsFI
eyQth5Jvd5+JJxvsHuYDnYC8Afhsg535lXnTOQyTj51MLjghwS0S/6U1xpYp0ji8
dp/QEuYuJ9unu14uDwdl4igzg12dH5II6PSBEJcy1EBZVDxt1fPTeK59zKc9lxyI
Egi/BNFspvgldlyUG2jvT+ws+FejQz2eDGPiD0A5q3n+idZiLMCuNfNR+xChQm7u
d8tvPK/rextriZOMOCHuCl4pKQ6vqfWOMjWruv9H9MfcX9jPoGpyj3+36Ejkgxjz
CVXzGQCeL0JNzppGQeKbejiQSMriVbwgnSio04W8aNCDQlbLku4rQZdNKVFeuudF
541WAdmG39fqsaFZkKfjbBdBw8WtbRxmRNHINXH4Aopx5Af+5aNJyI9GhjLqc/zb
BGfCMlQXMh8TToVY61SiuQH0bd42fk9iUkzibFMoh+6zZUdBeh6PnTdG12sEE/jJ
WBSZ7uNEc+2ZaQ+PjrPMLkzSAI1Sj1skU5cdWmFBr9X14QwY+9P45sj238qRLkZs
Dx2zVlXValxW+hxp1erpoqKe1OmKjyc2CQYTo5AbCYqwXWdvqrvAZJhFrrmSfXYf
PBVhX7ge2ePNWExH/tx1ufXC7ZPKtt6zspU3Yq30lzene1V69Y0FoOqbRKkq5HMt
2nPtiIQHh39rdAEmt5JMMC8JutvXSv4UE9B6xuZzT5A8j9In91Xk/F83lizZvdk5
aDSKkxkrMFwZ08DlIHt8G/YXzQYhgu9z91a5c5UySQ4+4LQrY7msWhk9v29vxFmi
AE8mcA+aNa332WHUjwqj2WQW6Gx8YjBnSHB9fCbUF6WNjRz1SgZ/8DWcbaKlzPxi
rCXQZvlxm+5NXRIJAgwI7vHdUemf69GvH/SoJguv92PaNrACh5tMFKHxX+vAsn/t
ogvGNZwvPBLY5TdgB6zKEIKNeSlqgNOXeL+4oBa6zntCPbHbkQHSgvIu57VfFWFz
WZ1qrzpBM4hrNpiHRGJ7Ot9oy6R3L+3IQ9KMAAlPimgG7wXztFTr9CrVLW3FynBM
L+S9UGZBvYnmH2cSLO4MVthhWY1OP60YGwLRBYiWUO8cJZkk+GBVWEyGnM4JNYCH
OcCQMvsZchR14kK7skR0WqNg/DDBm/wT5XQCi+8gHzm3ulmiFdsKPVhoQJB49Fwm
JrJ20ME9PVey6mDM6mSWVFWmSoygk6daiHm20xsCVVMnbNwlvDsNflcgfzj7VLYF
I3J/2aQEsE3Qm7Kq8Qi4Y1naXrif+Ftb3vnvQ+7fhvl0bJsvyzHHVBr3DiXGrUf5
5dxNgxjA5J9zIqDxg7HTC9ElxkkMLojZdEguoL4YizXXfTc1gQEUn9AWJUzIqSFD
QhXU6h4vGZa+yvtZl1B+n6kaB788+4RWEKmXFkRjveoH+kvZna0Lw50G+F9leRB8
fKORD6IK5zm9HjU5hSkGpQ3pjS14rygOdghMS94C+1V+95j7eZLORi00TLr1WOoV
j/z2UhbY4htGIFmatxZOPr2uRXlQsLl00nuHEg/j7ISDO8uyA8hYFIKboBH/HK/S
Cse0ciXhDm4ck2nQqfPlZ544iVnmQf53mMDSWc8rCUl1Y0zPO+0trgXw66TM23o7
7zg4IL0SrwSysZD3YKAa7lZn7DV1GSGowSADx3KTXN9aym2fjqW5EOcNLgw1IxBX
TUneOcYCgjilPThAmvr4XZLp33UPqO9d1/da6M6NCIceGRYB5UdZPCsKnLseoawt
dwTnC0AOU5fUAE4mLinVzxt9g7KKqaqkorxbzkzUZfmzLhByvF+w7NrJ/ohHRu2B
hh562i8mwfZzaa91TJhwDfzLKMXr1iyJVmAx+m+n3sha+871vymvl1zYOgunsW2B
dnfnqTWRGZPrrKNqOT2bJXSBdH8D4ndUxWkpi6iVkg1B6sm9WTbNTyoN1DNDkdyU
hzMlmMRzgZWqLTOzIWjg8YTQVqHSlaaVXM7LEiN6XVpQ9gzSknSeQjNla54obvH5
YBfvsmO04glPjlJCZDcnysH8SN8r2wZ+WpnGSCyPjRT9mDoGf2aIG9Bv9hVVz2l6
hNhwOpH7IVuEM42NbMCDk18omWfOg/0hcUHauL4NgFW+TG626O3oHOmBGYrBOQnL
xsZe7kf1C+DublejE6BeNxlqFoSSLf934W6fpw/pjY6BA+hXuJaIiT2CEnpQiB38
OMHdBUfeNb23eQ3zObKMrTPqelKXC6UWRMKoDYMF9Ip/vtUdzdoD8Q4g2lWE9ETM
LZgY9SUdsFXWiY2Uvmc1/yBJCi71OkK3DaBDDxxovvuVB7szhB6VgMkUahN4qLvR
+U2MrfX6eyh4t8hTkKYvaycnItKM/oMbZ9KdWylBjf/wyHZ2TgM8Zo8X4YEpsBq+
n0PdI232YIiVx0mjAJPFIASmIGDO0WXL/y12gGlPhXYjjK0uAkqn8pGAmhmyzrqg
LJWIiwQU87YLJR+L+IPUTgMRbX5baYFkLzr7tH9k6ws1bsM1qDP7yqyDBlr4yfbL
UNlSc71lpbdHd0AHXwVUk9+1aY1BJIjaH6++xBRUUI0lvpdBcrrWm3dxMik+8s2K
Edk0gOyAicMK+pcd96nLWn0a1coWo3kGqgwa4mf9AaYZiqcwcyA/Cy/FRvtncH+p
wFBJn14VAJTpRDoHzXLJswJlSFsViBdqU8YiAePyAznm5XDjuuPjOK25zMpaqCRU
Ix2Vh6Nv1Fq/q2KI4J27es2rp65rVmQxLsqsdnYx/ClWCmQWT1wc3J3A1rxueiyW
JixCWyZjKnN7EwJSaXNtgvNg8/F6aqJKF9RZztr/6izEMQ/1keFzsuGX0rKLqNEz
qkTVRQ20+SIzTZfJTwaHD7RnkxMIkY19BneADaWa6A04MwrbH3CpROpj8dPoOqiw
bgEus8cXnIIzcSX/hFDvTbojBfKcptGN/2VFXKEbb+xGDjUJCn3byhVkNGt1YimD
2EMUs9n7UWbjB+j0gTsqrOW1JHhm5BrLNfyQFVND7kN61Qioe58yw2KNjelSKHHB
grjAW5dk5YgMlCjmfEyAWSYQFSK+LXbY17M5DR8cl826Q2MgilUAlC3Wy4oOukz4
gzT7TGu3VtcNp98zwbPKNmqov5/Xq0804OttsfUEgaj69Bur4+9652CWFO2noKvm
Px1uembhGscZvEKvfD65rg3B/8cT/dQ/hLw1TcuHjcMTtI3Swt3b3tVcj7xU4z5+
69pYXDFOXFhVDRXXvv7C8B1IKzS2yvA4mmB+HYAScjTjZONyFQZLTCbTVnZVUcbE
B9OfjwCFuB2joEZSMZtjjzHyezZdOSbOJUcKSFYTQ1YePtw2fTI75W9yDkmj6+gA
fsIjpUZfNMAzFu8Tbnd0EoPCmyYxQ03aaqdVCsM/O0KU2/H3VvnfBSGgmsyvO4Z4
5095elkBnUrvl1vyjkLumAjxbAOt0xcKpyB85lPg2jxCgIQf9aNPYIKgmXv/WB9w
hQXfKRo/SXOfLCxBVL94f2G3rN+0dUIndJtTZGsaKeg5hl7X1jCuLnGh3ZN0YqC1
TpJqj66NEHd82dBswEQhWUk9xVnOLR58DYLOeJwryUfnq9qkHvtDOq1fADwOQFZc
3HxWbrXNVGwZFF8D8XUeK2OFC2UX7p8kWeUVg9VmhGsNDC7JA6WrFmRWLigF/ZR4
kQeUJB/vfvnx9qVH+Z3USYReEYJKlAmtQQOfa5eiE6mpk9OjggBdItlL19CvD4/0
Al3jTsul72SRIBbWrgIsFssGOzQ9rBRTMOhbuk4JKED3B0TkMlYrL909xpATXiTy
kGDEeBoXpm5pas+fVvUNbWrbKyCa+GQ4Y/TJ8WHwDZL2jAsrRhJSeHy8Y1kW20jz
jWZesEsuVZ8og8bQqcvz7Y7pLjx03rbw1hoLjgTFD4F9SXhievdEVDyJiUV/A9x1
73PQJm81Z36kIm6w9pYuqliXv58y1pgCVEo4uwBcKmmXsaHr36y1GxphKyxyjtzV
x71EWlvo9dP7bPhdV2xgdnhcxzZwF+U5ZHX/DhusLlYOAbrXxEWwKc97HTrLXcDt
S+EQtbUahfOsFulH0WCdFRbootX/V+nsfeM7sD8Jn1oW+RBzrUKwAeT6YmaZzU21
tdXsFAucrrTVDAofjH8dG1JvG8UKISqnVflTLM/+rZBq3zSfClrAqBYIsExEFqB3
AD0yW9PWNKiX8spDnVatPeQ3C9LB9Tm3vO64K3cSwL5AaJBXeHlQd3qcTmbkpB17
Z49AGSqYeqareXUMilddBTLGXQT71BTCYh2D8zjtiQ2pO89JsJse/u/10hEuDNsN
BNqUxwHxi8YefdxXvrekiygpHNflbIXTWkXaPNwKxQFrVatimoK9aHdn+cAPDyRA
1tBoLL1JVbuU8IpvFC1PUjPzuB+fgp1lbK6UxLqHZ+o323y87fW/VwruysIBDWqr
XOi3vo6zP4bKgO/lzIot2hWI8+s0OU+0al2j4Y7OZ7DuTHOaaCA1UzWmofpuWvJN
CHbclciJ5vyt/RhUfZRN+q67Bk1XNIBuVZTcVNbq9y6G7qfhjzPMC14ZjSe+Eq2s
IrOVOGvVBgLWWfT4SO8eNWmxWkgngpH9KIuq0JBRUtwFzGq7PNNx24xqufBO/8vb
8DkTISlqsPL07gD9NBMsJtWbqRkh9XT/v1sa9NzWsYSv89f47p1kDiK7nDpII0q6
jxWsesMLcx3Xj1N1VfyKq84VXWZWe4DhVQdzl31oA+T+IML0GdhlG7K8gu7i7d+n
BSCqq/GPOAYViJ7bQ657R+aTjRBKpXiKfyRd8owN18gH7ULTRR2tVoUspN5l3aMd
49cO6xGMJYlY/0Jcc58EtRPvBU2WyoHJkKtSrYEwVv78Mc3OKhUKNXpdf9c5YcjV
Ew2aldTWKQARbMmS9ChXv11LbZ6N0a+sS87N7mZZ4LPmQ273f8Qc8L1WZ+/uQO2+
v8Qkvhq9vcUBPFtbdCkLs07EfJSl6rhgYRcCC/vzoQkxtanFPKUV4wDjbBfccDSf
/iE4rae5pYeGZMAZwCXAafzYYWTKmWLCK5aEdfGpEHEW/o5LBDqJ4aV5EeTOQFZh
pxCGGII60e+D1x+Twne5lOh1qGSBlKcfgDjGPav7GnS9z1h4m6558k+ztn1jB8Je
t90epNA8yhvbWHaaVPUUSDt0Wb2YqfS+EVCiA6A7wtZh1jLdkWIfA6bj6FzsKDOJ
TM8QtZcU+A52pAueMvJx2hf3rcsJkGN16+r8ysv+Edph60XtpBoScFIIZfSiCr8f
PWi219FzusSxpAjL9Qx59NhBBs1nsOape7NP+xFOYnLWCy/aSe6heXPWQzcCyFa3
5pWd2Zy1Og4jNQsC2npP0U5hgQ2bTmQ+2AdqZMff2E6RzKZWgUrMWbnaXZ7F53To
b8txD+xhZkZ2w3S4ytx7WtvAQGRKoweaZ1+wmnf7P18v4NfqJmZcBsy51H6qetYW
UtcBiGWec15G+vnj+fe4n5s2/XDJQgBn/woC3ektrCEGKeermu53qc2Hrf4u+zOB
mglOncqvIFveOSov7vBEJv6f5iv8yl0IjPptCim++z1nPOxocjX/EDjDv1oq6FkD
z6utmcE6ggCyhhnrJZjXZ4EBbKzAdWOdEZNzTJblh/71UWo1gEsTbKO4iEtOANKS
86xs2pynIw2jT9TUziLgvJYn5ysXUKS9bm6tKqbBzlnUxIA55AldaY3eEq6OoWj3
38qskKr1hpwyd3qYh/cFo7AnT+8ifnukMr1S1QAT/YL4wGMIwlZxdw65HtV5LrBu
7JXYCrZn/C+p8Dbn4RWTRxQ5aG6RF9O+v7DBWU8uZY4NZT2EKlcgnVCugu2AHOto
I8pkadvKbXWomftpeaULfExAoq3D5sqxMz2+n/HxnqIxDEWx+HUTbXSpQp7mhZmQ
zDOhCwrYzqBjhzuPdPNIt1Tm9/65UiJYc9rNFb8jMdFLp6JqgGTg2YFmbViKmvyX
rQaZ2E0w8OnE6D6jXnbZS+yX/JcwtkS+NL9BjGRgd3rKYux2YfsJTrk08tWkJok9
QBF7kpztMFQe0FvVScgDBH6zrh9EUiM9Ll7r3dD1xFQRb38tKqh8nE7iHUiPSXjf
wT998Mq+kg/vETn7iqnDoP8+MWhlQuvNMsf/6syGDMQmBCPdz3q7nNuFzpooSjFR
3maaUWBxRvHFDYrLKVL+pv0+x57/ai7oRHeXrHprGO+AkhNJoJXSbGODh/SM/wQT
3KjVp1ObeR52yuikpN3iuvQpV+GXVV4TiFQGYT0y1ND8CScWh93x5i1qZF9LCHFy
1tDid7O2jNCvBckVXSNZokHpONuN5ihNG0gLjOr5spmG3WtXCQaUgee2+ZdkRc9R
IeDxHGIPXV9I0QsSOMGGMJQfcCYXsgBfwDyOSVa9pc+ohuqHkbHIlpPHRMvoW9lD
YA70uNBl0gRj4KVo/Ad+aywTDMIzhpuV0/2o+lkwARPjyPTjHGuPHn1+g9o1ldQY
KSJOci21FZNxnvpyn/HOF+f0NqAJkwHTgPdETvmZpTTIL8cKNMyNSGEG0b6sn6Lc
UVCKjItD29gvdjfk4bSXKc/TrVD9OSzt/oXToJyVcGX+Q92gSztVif0zoeXykvM9
X8MEnwpANJfHGN6I/TBo7eeNTPdK0KCUeHgg93DzahIA4wZxczSZt4H2V+Poa3Q1
PYMj9P162F5r3yipN99IVFZb1jtem8WLFEYPRlj1LkMMPv9cKKy+KAawiyXyNnHN
oOF1yAiA8zvZMfFbcOWonbvW4Iwhflv6hDJ8aWuSv9dLqtQTsTUipWujMqu7rIwJ
GPfkkQuLtPP0MFTJQeevUmZ//FWd0N7fYjIyp5mYkkVW//8Sn79h83I+KtJfmUSt
5i8gj5IwYpCcqMRewulQivy7O7EK8TqWD1974qTKpJgG3SvfveuuN43k8b8AZ+RK
zmCwASphy+0+Dy76pUobpW9Vjq0LeP4TQPdI/WQjO2NbIx9PChc08bbLLyVVQVby
ZiD4ahahakhMBYDyBw2AHgubzEDez8qSxO+UKj8n2nQqG3Jt/9aTrUtux6VE3fZb
6vxAO33iSXHOuD4K/VqKflua0CqbkpNML+MLQ7EtGqdq0TJxnvRsSOr8vU2KDPKa
VfoGo07zjvjnykRh4SuMuvF2H4fbZn3gTU8RmMBS8mx/M/iTbr5edM+pjz4dQPUJ
oYGldr8pxL+8vMVYtcsAWDTwwtHB/6/RbUmi8VNOZf7UZkvS4EWs53qcKwXN043n
kBejakoRhANpjbg4NlLX3q4rQMUcGwuN0hf5uBuSshd8ei3dH5I35GAJQsPAbwgb
+VR7Klrsy1Gdult4WSqHwA49V1NBPngIFV1Uyl8xlZQmEn7v1rMRt1AjX29aYfpm
+cdZKhSqgKoml7D87VMpYFtFxixfwUYpBWnX3g6hcGtmxkZwC1GpoOfsc4MQWpRH
aPAgi+uMKuV4XmYrhtEO4L9yARmhkPFWahzzbueLwVan04qBZEmxQju2KqKHMRWx
xQD98YDy4841mMhmpM05TQHNO8vrNi+aEbloI5NVbzroE19iZmVy0WosMT3coF8m
NWO4o6K7QDOu2Qwbl/NGP4xT3gF1h4kjG4feYiJDAw6buWBOmpKDXLSqsdkjcXR3
zLTgYMk+L1gsusUqEgM252VHVm6wCGZFXNnNfUxEyhthn2i15xmV05FYJ4Ftb/Bi
mm9fWdH1lG5mtDUkUiBPeHbS9bjpaO/tko4BRlz4ewcLo7UO6tb6BPoP+W9eTf7A
ESmP9sKv8HuejtCqRfGsVVHP9HYkXpYOgMZN3MS3nUDr57KAQ9vchsLY5/KUO1a5
n30HRPeLXkkMtH/fIMxts6q6TBhsXaBHZENu1IrkkwVjM2ksGNzUUsYF0vD8HMBj
/hmhclFcbkhbtVfJOBNNhscXKi+8zOnw8jYtEMg7q93MdtOd36KBKuPNhmtOVlwh
OSb4BOUSVHxhNJUJ1c6HmHcd/rZApt71KTiKtsUXEaWqWziqaDku9HluYo5eSJrE
6cljSL7J7KHi5rL05+qAyjxjUKDHh3c63eSW6qcQclrAeUY51mDIfuZOOJJ8/wh1
SWfVO2sdRD2CFEMMYu53pk9ZfhyBzYas022aDtTtPgdX9uKn3gR0H7dDZqw9DXEX
SK2Z1k2qWtwlqx7UPaqNNuEm0Dn1kRHEIKIr3OVsBB5jL7CdW+7IpejawzkrjkHb
ANzYljCV4Xr3TPB7qRIthbHjtYMyqbTvky7oeeCngwNI2yO/yXB1azDvH1TlNs5E
C01lDvs/fH8fWTFbCbSdSrGXTUNn/MFLxywu8Z3tqyFg7skLBN8pqW8KvcJIKtn3
q4/6s2T+KcX5Sb3HxRZVj6IPNz3TXDrG39Jspg+lg/l8tlcYvGZTIrLJpbaRYpI6
YRCxmKFtAcDCKycBGG7seO7/lxY8vonDz9kIa95/bpoSFF+O8IJNnr0Js/Q11QV8
R0oqR2tCViR1FwdXZiZT7Ll+hNe2SflJrYORNsxp966+HHhldEX2N/FMvr3NdUmG
21A5pCcUZs9goFDUhCPzcl8mbmBGx4EBPClA5tTGt/Ufaceh8Ig6n3XBgGm5Y86U
W4MAw9KYxYjK5avJ1ARX8ehZmT6BZuMezK6IjTA9nxWLxKUzrbQnDNQExN8moLDZ
gzs1B3T5np4IZojFmryyFMtXK+1UWIhHCpA3AMuPbBHJWWI41HQ2HgIjvKShEfCQ
DpbCLv+pAvep2am3QgIsvFJ3KDDCcWT08mwBUHqCh2LcG2YjjlMKGestY7mLl6UG
MIx2CoMsnNaqh65VkuGvXiYHIQviiDHYAdIRGI/g0B/f/7kk/KcczDsdRW0ZwENW
ZwrmZ+tM5fWnoZ8hTGWi36lPhMXQ9t/t1CrRz23I+rDCP4XzuATuw9QMPxderY2m
1GQQskiNVy4WHZhWRjQMyU0NzHyaYUJxdYMfD1DrHeAwuCdaYISqKOSC6VwW4gM+
YdkFbSW7wxMmC8HoBvuOb+SUmihtQTomANHb1sKfaObCfSIrR0lXyfsLOV5sIh+o
vs+6VhCyZxNuNsqzvt+rjwhZ2J9FELQCmEvn7hv7wUgsVw4uUBOsPQ8i85baYCJ5
ABfz2+OMdJ72SrcMSEv37JugJbJnQ/ADPmsGp2MIwum18tVyFNBcjeLy9UQy+5Il
AbuInNEQi4rk58DW9Ovnr887sbQu7mniINSGprHHmkezX/n0smj174WusEgVroec
Q1N4gjLKjffVWr977JhJ/SgU1J4gPRV9XqquslfKyW9jCf/FUjC71rY6PAq/IWM1
XmEchlLJj6dpTEgq/ggY4DfzwuSETt3wBnn62F4ldk7OGBB1xMIEVAfyZHabqBF7
lUhdsBnbQ2jl/RnBIbTvfTIbKv6+3MnCrA6V+voA9M6UnF1xF5WFE7jQRKPcuTFl
ImGA+yTjbAJVo+7yVDnbKl+TKokqY4aEFTsYh6yO+UOgJ9+jpCeuGqspUR7UDWxe
jQxAYhrAj2dgYG76DJSQiEzJkKr8EjKC74oi038Og8G9QkcCH+b+5wSFnWAsXWnq
bHwKwCypigSRs/IvWzSiNchQcOxq1o8tgWgnb3+GQgsl/DesGCgSDn4xwYgZ7wcC
LdHktixdXEpiq0KZZctPw5rwReaDmPihV90kTX7DvJMwedzQuYACoqGMqETfKZIR
4CPcDrQz9b320B2WZOfBV3VbcDShhZtefWuSjlmsPTiD83BoKutoeK/mPDpgwcNU
mvBMnRfaFTLL+Mx1u731xS8+QYmTxNMR08zv+4X8zSt82hIBW657B2G8Kf4Hokck
9Gv6VQwg0lFWmjjK3LuYRjZqeqVRFm1/MMYTvFiyTdkexSetUV2Ti1rlg6Dp2Z+/
JY+GicliT5OJTVjxOcgM6qZqr7yIXtbrug0BFVHjJXfF2WkXp86Gau6RK9HbHwW6
WFhmSioyoAAgRlNM0R7/NkhhmRFeOfn69eb70iKNU/e51TpywF81XwRDlt7fUlg1
xAkb8HZnVTUi1ZsBDVgQWjkv5JS1gMoVanK3FFJPAUmrx6HEvJTFxT1D6O0wmHF0
5Po708Xm5UXuersdgDe3+wMSIZq/90rgvNRvTHeEKcuO3l70fw3U3Xr6oBdZJECA
9HCmQNCCfURFHytL+8yF76m29XnoyF8aD+YshLXqNAJ+ZepXUrpylyC1MPQdlfYn
iYnRljKY6u/EF4K36zPzwN1LO5yFJ6zzfXK6FnjVyAe6Qf19HyuOAGGj9feUVZFA
gBnnlVTEOXW9pAcy/cpf/8QbX39yc0o1Z2Ei4ZETyIAkwJhUKAmaPEoz5xkJsVLX
tcuhenwpp+MU+q4odDcac3+gENHAySxCubdjOZWS/FzRDnqvVNdmZ9mZzmPl3S4j
5Ssdw2IirwNL/T4DYwyjMVfRvhTODH8vUtegwuwfgiU8e9TIvnx1mxpR3XUknDPG
TPvgH0EB55Nz55YJyOrejivvz257exWbo+jvckYRtTE8YKM22mDgs/acEUAHQEBa
fKqUcs2N7fOHFs3tr+bw7mJm+GiEFRQhFI+8px4bt32RO8M6k5jKFiBGf30V1UOh
pXgf5kOSuwrD0wxNQjsdHaW8bT9Nq9ZjnD3KDsEvH4SmK2djDQf3wPXZ2r8scOhV
cYgiMiPlA75x+sHx5j4upR/oWHX82s5aJJvKBr3GIUoKFJbEb3eumwRoctdVmK5K
V7QapH3urTalSZC2+v101LJRs5o8O2hXV3HG0/BpZgNpLfAoHbh5hrGM/s+HUAMY
rI2i4ixPJHHmSe66q73fUIhAf14mvJkJ+CvW8p31A0NeVscRoEU3z3P5NB+U6/jE
6vJt+7EhAEdE8RqbvTKtxUsuW7fVrtf40QEuhTk5FOV3xaiMSxEd2XTRAVFsviuj
BjydBFhuRl/uPItJEPlt4Ttfb6M9hcBhsRZHHk20l4e8jXXIprd1FQfWhj10W9nF
EwzKC58DNHAJOD+IvNymVrOqZgOpeJ1Ui8BjXOvnPupAcyogMW5bRLbvkm9xWluZ
w0I3ijPR3OmS5naPHjD1j28zTuGeEn29lT42jac6fDy+UWEj5ZY0M2kkvOnP3A2T
tjjPMYcH6qKE4XQFAp3FcS8jeN5CI7beuK8dUjPPNhJPpGdofyyR0lyUqN5QvBpY
3SBzVE2WFe+Dijl5zDByoNUC2jogLFat17WE/eChtDpftpJAc7GYeQanc0VkduMw
XFfCVIFDThtPPrs/4gM1uZHt1erKg+VmRYmpUHCmJ06hVilAR6If61Y9S7PUL7xI
6pw//lHAWOND1WIe3KvSdgjKHXP6XcvfXPD6ovilqtzkz4/nbykM6a+w+oF1Kl5J
5T7xZvidc/CBMW9zyvs9akEvvimrQsRwe3/c91wXJE9p6UUw5A3muc0VDMrrrc+O
jEH8oc6/eyiOb+B1SWetYhCsRl/zSv0xEqx8SrTUlDb5mVRtKCer3JPjyS0ISsri
x+t94Y9wlzrG2MTGSUpJWa19XeDfmBRKz/NcFFZWXOq1PXKsxslF+BrIf4Wfwo3o
pHeDqiclNgjy/dzgLeh7d+aY51H13bNpcIivXM8Srwq515N8yLyuRvO/fnfVuTRg
8PsqRuM+WALvR/4wa56iVJ6r5USL4fuV5qZk0wUzc2ZZbBP1q3Xu0cAH3CeswYPT
hrwQZ5Bm3fiYQ6y7DLgV7QKm950gjrmUuMGoasL9wj3nK7Lkhhk5MrH0SXrNoYaM
7QQvW8tPPrzFP6s8MVonQAPy1Wr8CQR+BnPfDS22FeSDDivSDRCvvY9SR7+TXE+R
tWZKvO2P+gWZcAM70/wtNQHUqzyAYicCMXWA7kfLgEZ/PJLiPwEVk894YOiaxE0h
XUijK+4VtiliKRWcqnBTrsyUiyEHyRCgeGEDu4aOm4AGLjE7LEoPPsy+wcwTE6r0
BE/1cqRA3/IuqSw8zmpGa6eZiN9k5byy1AaNja6NKxSXUcAFzGtnBX9oilFhyu+N
xBo9mxU+KR6yD172ZmKfg1+vcq4qjEJVMBmStKv/5gR4canHvMepxqYHMMbOP6Lj
VR0JWmdDMyvkpQVIqE+naEH8jXIaZDnkFTzUzOglun525ynlelRnZxNSLgcoYIsm
dVJDiCKnhvjXA3mgEdi9fni/HBNUDGKVHlpOLLwTeesuPteme/jbnmiGiqALQd80
AMaOHd5AaT0v82MC3MLoqF5CkfwIWJRhvm8kdZYZhoJz80EHIAoJjdjoMwf61Jzp
Poi8uEDL6ZeQCn8pcZ5fTv6tuLXqdjknqAdHH08TFYpY5PXcard+Reql4W4pHegi
DWq/ATPiTPJnXoKVrrWS6mOrdqQxO4hRwvA8FXo02FnS0aS2ly6VBlN5CrRkoLPM
Wiu77dH5P5pUHdI9xdkkv04Q3jYfIMGVwECeu36hvt/smEsInf/s/gS+J73QN1XC
MqSpR3HeGAAfUfnYsFKCoTkV7WJlBQrPsHli98Mt97J1gfX1hzV+EKwmbgFuxhNW
lMQMnrzQ6xZ9SjxW4mcNZyD8ZUx3Gl/jYA5NADh/X+t1m+n5D8shq6HSIf+a4udv
Pi2qB5u5deEHzI7P9PmsVLvy0fDZwbwqoX+MJcQssiHT2fPQMEO7dlWox2055mp7
lgPgPYIoqcrFaN2IZVKUA4eQm20Kgbj5BTmkB5sSvjECvgXNPV08MiGcooFgGZlN
MZPOIApKswjD3lW+483SOK8OoBn99LmIqAZO14FhbuHwRIG3qLymJiFeZaX5qt3Z
5Mj6fnSbbG2vhPP17k1T6W2rXRYtZA1j4TGkueWngTv/cOl4MEvF8lsz36IvL/+B
8fJ90FtNKuXFqbsdKuFyyXRRrX/U2IHyyjC48z6rZRMizcoLAXXOgyvHULV1uFtk
zlNMquvPSgZLGP78mdAv0ltY+zOH5QFbxmF+igeZ/RRaHPkkz76ggy2dDEiQJwbv
xJN02ehGP1i6qa2va0bnpCc3yoPHrB0lA6g/NSd/ptpQz/S5T6T6Hj+4LPbD3mX1
MJEOeSeVwPY3i7En0XcWCYHM6uOXq0jR6H5mlHGY4eA1fkYhXzFfJWCznKxac+wf
XZo9vkj3UJ4Nr7ZlCOa062JhctePljCp4BJTWw0BC41hSEyLR01E8FNpf9WCy8nc
8sqFNQdncZQocVNCNp2UY7hD+Oo7FHgNfdgbTbq34ftnhllWnSVE49cw2A798uW1
JPzZheNrWLuXVN7677yByQNhabk/Er2c7axUThJ7G9nPt9xhZjV8P9iXn8bA6rJF
odqtUn2+vTg33RGkJlytrEiwGWSuD6gIA3h5BIdOFSLhjKz0mYocRNc3fZXXwlEB
YsO/Te4pxedp2xmCaSnDMWP5rYtcOl6yJlLnvviUE9EK9OaT+2QqoMpiryKBPbtJ
L2AotB3WxriUK08IqtwRNemw5YLpmaOebMYDzT3YUKgvHzA2JdzgSY+8/O8mg63b
PkJ9Nq3tpjGVaVZgViJwXrHKB5jHmDYovwuuuvjNS7pFtIpTagjo4cQhM5kTPpnq
Gg7oPfiUXWz7vCKrdQqJRCRGJrQ4NJ/3B69kZiV5RvYMuhG+tf17Zoj2zNJ/PCSI
Ijgl3AFxFRajiNTaeYsyos5CDc7W4Ahco/KJtbyyvTctrhArZidrDeDMSUQ6T6Gm
C9qcqRsgX7gVsdsBP8eM/0W63CwjKW6zrKEXhyGjKFa454NNh+58ehXyotc3TGYm
qaijHiSutoYT2SY8sI/3+O7HgH21cTHG6goN06MzB/6sjWqS7Wt1EtIdZLOF71qc
3AbJsjwWceTeLMC7hnDAVzoO9bzEXSIyNxLqw0b4Dw8RiAZXtE/G6TZaVDUM8OC3
GgFZFDVhnVYR+wIkWVKZ/ekUjsgb0LrZ0FH/aX8aLnONUo1xx3KSrxlRBrKdJOvc
LndvfEm5iY9zF0zgEW/Zd1d8ALhVI8ZVN4KK/JSe6d7Q6WuKSd6QxMbtd2pI11jE
Z2Xp6TKWRetyZuq06Dm6giZpKhCmG0LM/tvl+QACotRxKdA1Z6umgeBLyYZI4FK1
uCTk/cbJMkxB9dUmMKyf1AQUwK0a0nfx3XdPv34glH6bOXPuqysY9Urma6e6B7vY
j1wItnPJcXxLIqfW+UwbQuzqUOzacqJVYJc2EwKu4zAXQjpzl4gPCo0303L4an7V
3t2ob+Ke57TQZLpkQoy5XquVfZglxYdAbjm6CWGO9fSqdnrX4zYiz23eyt1JATd3
/OgIqFkHTBdtwviPcugZzoX7m229fVAJzkC2I/spwtKZbMk79HUb0cBrwbP3v8rV
6rckKBf57OjcMWNDx3RxoHXEs60zq+YRk5pNJ9jgDs/EuoNs5A5DLIK/pBEskA3T
iyMdLZbH1GvJt2Y+Y+6FzBxhz2qmhbSEyqO5y9MIVh9O7vibKvgyMT0gmYyUiGUP
LvNMIm9M5Fj3RbmHPNQzkaXExUdnVlZWjBw+JDwWCRYcuVjjNzXqXf+E8udRTEDb
vpgAw74wYxuFyfh8IimHRYMglk4jke2lkRxrpASSVxrbrOmfBVF2aQakngxpUQge
CucmyzMTbyZy5CozI3yXks5V/TKvt18TNr7tQDXpqAjQYNsvZydnCoL4fEFrPxnh
LzTdcRKn2MG6RYxHw2clT4TaWfJshWOXFdwalE7odSJkEXkiZcNfVv8wg2Yf6tA0
ZARaXXmizE33SP2G4DAV2xi56ExPXQHEcM+wru/Sme5CnxGVxAoj/qtEeDO3dm/+
1eNvMnrxaT6lm9IzpZnqXQVy/Ho/spFpFPV1jeywo/loNbyLLxdmU5oG5czrlI1v
v8AfiYgdrB4bdsejPo2Qb5pPBSe2CKxZJRZQ6afAxaqcwEVsL0mWppv/IQl2fyMz
F9G38ihS2OyzccB83qT7pQAjHvvo4hpoCwDVIwGv2pMY75ZDgozWGZtt2fWOxnz4
5cZTLDHzNtWw05DlJZmY5x1s04ejWbpdoVXxl5x9+QLw6Rw3wUmjEAEONI5THSU1
+RZT3SeSIFGZTOoyhkRcJYHH8JikT6jKzXRIBzuYggKcJhLUEPmyguml2Nq5FjQJ
y3yauS8DIkVdz5vZw3dGOubsRgSgoFo7ORtkk13gFb94Mkafp4d1U4lwL1mtpdax
AluVdtlIBJUcU+TFwkBIPmLLwFGhe74Q6s7QSCF87Ybz2+yuH4+4krp1op9Nm6I2
5lmADIAPIzf2sAoyZZFiLgIl0tsQnr/yUybICOE2T1m5XLpCPX3boBjuKdFSQSHP
usVoXH/TQDrTQA59+2sKe1qRX5fHZZt1HZDzQvW2zZRD7BSwZCspwslJSJkNyl+M
WLcuofWbpswkZfIyhAQH7OU6eyOZLMLFsaHBC/mh2o7ncjMZX5a6QO6X63dp4vyk
q8bmw2gLFc4oRVc3IEGLabtTtZ5+S3Jlt+tu91cWTcmaXeJZxJ56EnFylsryBPrO
6o7F9sACpt7t2K3fnVh92TXSC2W6YowmHICfjgsc8LkncB7TvdVn32tlE+tb1t8O
RbVzHpHDPlrpJXjoUxEs8T+3L7kEb1+cmSW12eBses7SNHPhlQ6B3tnxhTm6+VVe
Z1yAzgVmFt45rEY9yqehjrLcI4POA46uiMNmx6owJWgY9o4h+5AmloUxvjhXWY2t
nknEqjLMP0kf+gKqWqcEGh0f1dcHxBq0G3Tvuek1d4TEsGO75AyDP2ZBb6Jf7bmp
kiFSzggJl2Xu8V9ytiR0QMLdbU+B7lQAfa42SM23cezdDxRUC0ldueVV1UUJE81B
7cS+xxGoZAdQOZltRTAI7QqfL5qaqYVtPoLp5wFpODXpl0TtrhdxZsS4rihX4dTW
hvcCYuKhzMTqWIo2UB6tsmpKHqagh149xyzMlbRdsGn4bewVepShEMWXCtZbkgHa
M3KT8aEtmuTpM8lcAtc98wEgwDv5pQYoQdjl1z/zW0P//B4TsvS9t/JetxKD2WNN
usksFBHtojlx7Ltj6PkruAhzI56eu/MhItlHHt17Gt9ryiskgBHuokS2Y2TXB6Oo
QfB0dPI8j3Y81ZiZT6QKBo059Q0PRDWI+LtKAA0cIxSvujpK/LJhfN6ETnpvixJn
ZrTtBW+XJieg0O8jkvVnK8AUKFSeDEWsQLU2yWFwIARCWzpBb+T2ITgUFYrxKnNr
ogQyM9lVM+3mEql30jCICfjURBU/HkXKjbMkQGmMJiRv7i/cFzh1lPkChqpTtgaK
wjDhY3dwiyoAZIZrLUbqhbv4v8v5G1if271L+Tm77/rhi3fnutk+ZYkUYarj+RTK
tpvdCJ2IUPcgLED8sUAq00TuobrRUyeqo1ZeNbauexBTiuMt4k12RJvXehP/Ze5G
I06wSZnNcGLKTZ4nHiGyJs79pBbOGIg0r3v9roNNeNVbVfZPUFttLdt7zdz0eAdT
dGfIj0qi759/InsP4mIUONLBtk9TiRMDSL+x+V0XPezULr8XsdKXA6R2f6/GWqX0
NIrA0UHF9/yb318v5U4ofFX9YHBWqn0Q69DG7MKkkcX6GFW4fjl8wm1B9XcvTf71
McmDaFQq8M/bqHBnau79LXkGAejwwIU/gx6KYSEm2YQNnDVvmf6prm5Xb60fA2W4
YHFah7Jja/yEeVD9AXewT2Yr+xkELW2r6vGrfGtlKvT1S31MC5UQA9f9qbHHkxZP
YWz9j8a1jfO/fhKlMzdF4Xkgl6/IavpX+ZqHB/IF5aPpxICAbQrJZ7qGyfPUd16g
N7nuZ76jPcdS93Ff4QVUBK0BROApFzJakVQB//7kl+4+Ote0GHPX0bNnC5mt83hB
zLfSiCBiRA4SCDi5qgyjTksGDHy6evWJh6bPHQfWHwyq/CaRHkzVgFvBslEdfjEC
DVunmDObsKSzYNBI6MJOldUMGsO0DvvIKGTbbDWYrIazYRVWfgSX+Pq2yLcVi12N
VJeA1porDA/7YNVrqTtuhFpNey5wZR+/3+g810f9vzyafesvDiWYkDiR1uxQtfsL
m/7ShN44Khl5A/gP7B+My/s3DsnU3qOvd73KogYwQoGZIZg2RdYaP0o0XdrdtQUM
CNX0gs8LmhGXFtHXdIgEBpMHiuGg7CYvWd4bJtgsI6RwlxwhhfPwbZJK1FCeKHM+
iK7i7a07l8E8IVvInQP54aB28VbaiOqN77UUWVmKc1plZUN4gx1bSDvNTFnkYt2Z
93MZm4Qk2sIfyWbFG1LZGFCiIo2GKYNwKP3mVQutTHdVav7JGLaHWmwP6Zd6eSD2
sdVW/RHjHSAacJ3lkfM3zU/tzws+1JbgZyXojFmm7XGtlFKW0cMWStdUypdZ+U1I
6fp56M05+U8hRiDG64UUSMk47vJb6XQKsKYWlHR9lxPo2VKOgNVvXyBaLQrH+Rg+
+pCYgY9Aoml0ZNblT/wt/Il6jt2pPmSYQmaBldL7UuoR/v9Zfdgq+Dwc45kNLZeY
+0LKjucZI+PDk+P3S9tcQvMyafkUIvd3YGK4gRPurJYsWL4nPclyJSz3XA7h8zQ2
ET6wev+kmAKjEevV2NI/dQDVz0Ss25lgtej+J5JOo+Q++fvTfBTu86yahN+FpFnI
oTSBj99ypSBeMD8bniYyk+FIi3nRWib51913z55BYdyVIqNpeO7EfYx7ITEddS9g
bLjOHpX8AF9bTnQ0fJ8bGK8gU7aua6ST4wc+Nl0gDaZ5KU+aPz2c/LcQVfLVLOJb
Te2OhL6961YbR245EahIa/6Hiy0OQx57QCMk+XSzs24hX8E6YVBG5CRvZvY1LOT2
S4V5A7yF8zhLJHcmgWuVWkC+9Ka6vM0ahoJJ/hupEtA+Z92QDVjnlyB8HlJoJJkJ
RMsSEcLXOJ8bwKZk55GJ8dHtSxMcS0wlUxD6p04ySf9/XESKAVeh51al4Ccqt3M4
KtYQUa1AShqVufW/xrVQrDwTIxx48IT8gwtF+zR/HiuLjEHpB7ynb9R6oVghhFBA
IqVwlaYsUynsyO2QyOOdrZxMvJMMBMt2yzOyYGEHWeX1jwSTdEqCUDgDtuu7RbEq
aJxx9VUOkkq+3kPMmMePncJNN6FCkVUX7NgZ3kDsyo19EveY4jeVfHS/+0K+PVSJ
X9HD1hgKgc4MZuvybrprB617jb38N0B8OTsc16tmlrFsLqEa3239iB+86gyBsqSJ
bd5P+utUTOHtS60DuU0cQ0F0pse1gEkhG4HW0ZffWZCc2mCg4bsrJ3w/eWxz2EYo
Ww9IIuFZrwK97R47TpabfOn2YVtXne/kaNVhqMW5Riu3XRupZVc7eWN4f+SmmXtz
eN6XOVypa/eFgUCBJ/n5twhCmG2hTaXD/xpdeM/Z4Pms1pMKb4FbmwMl6y04WUBh
hnby0ftEXlxSQb6DgzYhIBsj8G12QkSTKUPugmYgKwCu7Kq/UltIPJzfNXvkwoPO
WJgKuXSajX8UZzX6qTNXFTInI0a0e2wvQbOpmvBwxUvvdtctCw/r6aSAjYrufEtS
6azd3SFQ2iV4FaQFZKUubj6oNEHq61CDDOAhjuLuXxrm0u4bVepAWwsAnp9Rj+wt
ytxg/v7k9gq0WeDA2/w2Z06lj2tRQtRoBCFdN9PtDYabF4Bgy1h956KScPYAgAtH
kEvhR2jdjzoXVjT/W6tbZtyXpJCknBcOb0K/5OWY3Wbn5Jq8FHiKUt6ryWPmocHd
5/gYNCL8hfCf5/TFkXeg/6iLKwswVznir3JdnQch3h96nJii+MeHBAKQC3WGVcTa
AXlPkWfzErSF1nIqrn3KcvDbSeyd/9jeDZUlx3xdmXu2rm+bX/MtJCPX9+P4P1nw
DgQvmZv9H/Pa96cqc+Txh+JIgbox4LG0DVrzxf/NqdS74HVP1n3Mh4UTeXgIn9MK
IS+lHq2wmb4omMvx3gsmOXh2LgEcbwBbqZHbEpSscAh/3iCJAUo6pEn9zkv5KHPz
15HC9O1mbwoexAlzhZFYTmBg0DeEjAc046h4TN3uQS62tkVRAge5IeNljfSEPC8+
t1BIHvrFycLZ5TdKQo0I+YOA0c4woOpysPvu+pYkp8/T0TfCGZYTI3z3eiVETelM
RR3s8P3wb5x12pmG3rzdzIm+wyXum88rAW7vwsIG90RuEZVMqbTRt6Pgtsm6Qu0J
+W2NMUq4A0MJyzwfzoV34RIAQPuy2CQATxB1BqviJ4wXIKYJMgDnfmERuCJbeFXo
8an6DkX/CsI5GRfXDVcJ8zP8GqVF9ZI1Dq3yGtRVyxxA/RTWmMS1HqDB6EIaUyiM
c+BU6155HWI3eShTHXUWlelvrnXo5e2Ggp3If0K4mXzBoELP6xljX3RkEYF+46eZ
lVogHMMl/VUGHp97JS9/wtD3S21Am5z1uzk5KeiDK+B8mJ4uXFasmsWqSR2c/opV
v1FRGuhZZq/tlp/So+fVHR51G+PwvBD8UpyllPGXYlRgSpVIZrTVIttXcpA5hgis
J1E1lAG7r3neW5rVXSymc1H5UFZoG5NyMyiZ6Q4pjy79FQ/nt2XB8sa/fC+p9JzD
OacylXPmiaCbut/aWv9ICdCFkgSxGtEldPfeeqe99w2k4NaFur6GKerieuPU0Gin
AXMCeN4IaRYevr68OC62jVK8wYMp2U4yftI//L9I429RlgzJ4bzqGHNXeL4kzjbo
ienhlGbK81iu9cPTF5qd7Lhof/q/lTGVi0CG0/6J9mVnHfOhM+hO4lC5KkU8xZpv
shnkgFsO60RzG3H3HL3gi2dsNIah5L8cqQoHX38qHnUhVBMZ2RigiTpUxfTOUHBt
swbDmHo6Y7P0fgbk9ikI6OCne9YZG2a8+HAkJ8ginPeZGievEz2jwZSUvK74kW4j
ah6wgSF+1ZvMMf5QLkHMHnuXxtssU7Cj4Zca+wbNaz5dnTFVPp9GcIkwvvUp7OZK
9naIbI7hcZ8rld45NSDQIxCVmyr56jOfZJ8BYARWl2stfjaeZhclUW6C1StySX2E
gb0kngUSop9MxLu8hxSAStqgL39a0USLIAzJ0CgNRhHt4N3C3eNUsgZE8kfq4WKi
Huc9kMqdw1cg/P5SjFrTy4H9gmDBXegUhUfrcxsiB1X+0TLDkwgfUs+s9IOhO2Y2
Gl7/LxaoBE5Oq+53LQFXGmosDhBNd7qxM1x7lEvazSc8IkaJmdAQ73uSPWUPdqmj
QwimlUhe9+v0VT25RCrpWZ/m8ptomJYVSnd4qvXbW4yQwLV2l5Bqsx3/Uj+eKuWY
BqUj1LeLbZcrQ9pLRrs1X+cJ7Oi2c4kZawEcJy0n0v6fMnT4pyN6L4pqBlFz7/Ao
/Sjk/3jeD20RIvNF24+yUc0mzNMo4dX8JBu8OZuLlYH64HpC7KKQTkWnPVSRFi6I
+vSGfpV5AnT6WPsfmnQdRGzs7w8hzK+zqlmYuL1b/7XEPKAfbRBQkzub7aHVlPlf
EG++RBL9kxIbgsyD7OGRDsCg9XuSyy4mc6RIWCZ1JOCP2XfCB6itw3B/GxOmhBV8
mA61SUmylQERw+LZe3ywlSbHJMHsHh6ZQu99z7nTL+8JAOXki/6r3UNMhKne13ej
2cbIgfEOZj69elq0WZcRTAo+UHFFH2BvuLs/WRtxgVcWqhgLSJQdQrxb1ihd6M/E
DfCNDssBLE4HQZhXGv3meIFJZxKKbvAYLfbs3xjXJHKfj/memSXHZnWO26yq+YxO
WB2wVBZD2dkb0WIW1q7ra9Y3s56Cnz+pUHtc2FCVWGpmH/ECTRsj/hByaDLLADkd
OhsLyDVx7M35LeWFCvkCWjuSDxjDEZ72TGlaiKppfHYt1mOs4DIPk8iMLdSj2bmS
9a/05+lV0JV8u+br1w2D3AW6B0PpotfRTynAF+AWv2DP9ANb5uLwEU1/SfCvZVDO
RR+d98oyU91tDn85DL+DPBhXRqGD9bZhOHew+7RL/WmYKw4ch9CbdDmL/pADPx3V
LPw9cIdNftFhmWKu2ToA7rjO/XApl+lXb6PoLM2yL7LmLO4YGmTjg6xIHExwvHOv
MM/JXovOffvIGvVRbiDxGIcnOJrTTB22qoSMtl93uyxpHPRwDSCD3J18sQeIWSNK
KFSGi/sFozTCC8gss0IJNtHLPX1zp5nKGN3Koso60SFRncoTV2DcbbgAGcXFao9O
cSLm7FM86vb+evK8iXANuwinE4qpjtbt4NUecfL788xRBYD/8Qd0SxsCPeXIZxkG
CKTthezuD0+EFMfpTbs/vOXgoEpu5jxhQg2oo0v7RL8gJv+VHGCE26nHAH5T/38n
SNb+hcd/n53aIzdK7QINGkiQfxjmxYQ0BYlkZzmiUoO2yhsFV6FNNo7EMT5qhtou
bqqZHw+lAskxe2yejuYdWq5UoV1vYJc9z5i34jbUIR1Zd07UInk77AEQJtGxNr2a
4D6mPWhLaZXr8kgZsegxfeTXsmzeR/bVzvhej+2/YoAdwr3Jv5OlxK8QceirmBOB
NjI5F/PP46/8ZLOxOGnkmAtWoxatRjcFuaT8DExJ8KvQUgnA74vggoPgRPhq9sWz
PaH8I6j5RHKLwTh27beISMRlAUKD1MW1aqsJaiERMWp5uU4wys3FJi44X25strnn
eIpoZMiFNrHvyl8VeLUDg/1/WHRQH3kSh6lvEhmArNMSIQckrcg4SiUwE3AF2JB+
QaWKjpufdke36XtbjBKby1QC5WgTnaNNYFpOhC4lZbRPAY4BBTKQGKvmid3K1Vle
Pz1sf+jB/a2CDSCRd2OgV4zFKdIMf62/y7faMBB0L5Uitsv7Bycf5ZYfEAgQxd0Y
MHD3ayGFO55xbgJ/URjGQ5Q2vfVG1iZX0THLvQ7yCD6gS6LHrNHNee3+djlxX2yJ
r1DBjB0g/qs+cpAO8zIUrOBzRbb5wW2kaOb/mV1cxHuUiO/jkRNgrBoTDIun3c59
BoSi0wjp0V9frRmvuzTwJP6FRrBKuhdGndfmYnuo3TMsWgFPqptm89+52Nq6AoPs
3rvghjn9NV9go5H6W2Lc7CUW0M98s+zGqD9Akdaq+HZFiLQgkVApnSZL/oEdBP0s
4mHu9itykb42lLV+u/TB+vZQ5uYHbqA3KqJ9QnlXC2/4LGM0IwQgoAtlJMr0PkpE
5WT5u6EjIfAIlIaK/VARvfsLxeHc6cl8U1ivFF1WwJvWsZABv/lEsWvM5muQc8fV
mRBw5OBVlfPojTUo7vTivvxOwDoUovuQoMWfzmEbeU6OX6raHId9cQZnjU984GVL
ROECZ84D7Xq/hwZDHrpawVgh6AJOPbSBT1ib4PgcSpfM2PuE+sZdojgCbV0lGlDz
eZoJ90/lQu3xAB5xxy1q2Q/maxHTMr114ChXsa9kj/MZbXso6GBIBDgaVEfd8rTD
IAHLo7bvcO0HZyTM5YM/dwofdYGLhYE3ljaR5XUnR+J98o7oJ/Myu7LS6DKoaZCy
NeevURbRzxEw8Yw1PCavC9Kiz5DqueTwxlO+bQZ2Yx/s6ssaaTnSjFVj41Nc5mAR
P91+0bKhriIM6i0bTlLMlvwtaI7JE+7BLCTGahLyxaOQ7DtNA7aOWfNzMQ079v4/
wwDUJ42x3qtE8yhV9NywxfBy6PAuyLyx8oIGZpbuDgD4342+DMdF8hj69JyEnsfE
//QzTFWZ2U/Z9tSl9JUQEH6nxcXSBx3U3T2da/tWPeYi6evipzuPmfRSuRCuDbun
0vgWQAGTTL9LUERvXagM4VQQUz5SvwiL4zfJ5GtZbcgBb5782Roan8wOJDdxQdRN
EQB/N57X2sjcMW19FG4c2AFpkFJ1Fk/I3a3mBhZkWFAmaj2enrn0mhe5ZKAW4BEI
PnCkekiENMsM+4SMCggibRbxlxckQNJ5IOa62oADn0q2rWXCnLYypuyzVxi41L8K
JZl8ue/gJ9GVVmNovjSeNc2Jn5l5j8yChHuy5KWLONWaVz1Lu7K3zRtH9wVLVQ6u
A9rtwiQpar/NQGjs90fsJdtRD4JWWicu6juLrWg7BKnPC0ItJONb9O4gp9eKR9y/
U8JnhOG4S/EqR25aazYmp7MDuPq5PQPQPvgKZlm2YquqyYY9kSmrM3EAf0nEZWEH
SfJSnjMMz8/atmFNt9gUtLH0bGBaunsg4SZLvTcAWe5ynnlCA40RQ9xtaBwOAqcA
ORLN3+78I97GJG2Ld6kvfP8f87OwcBJVwPgfpsr2pdquA5aHTg5TiMB/qYjvtGJD
fNg+oDO5dddkpSYcx2l4QI5dIKThVZqJ+JEFrnhJQnUktEaaIb6MpRNwCLxQXPLm
AvOOhe6aJTliL58XGxxr96ksSqhyxqqv0rFzk3ZFv3iuZn16D4fbJ/hQ071jtXMA
jk/Dlzx3dUFct4AtcjWVeyYQaVkdARIwFcte/EDKk8VI6ldkeMycsytArvohqnEA
H5LrMYC0GMVhUtypMrNNTAspYiDTlWyGiIMyKf8ggUNaN0w49uXPxCX4hA+Flwxy
uedYRcwFhyUeQBJCaRvpx6jDZf8tdX08ZT7qVIToAuHd/zCn0wpVLMdyGX6sXXSe
L4lQrBY74RFIRWcv4lTYMMKS8lJU0ly3sgzYr8JbEWL0NzFyrvPargTUqKhoWX1D
TAnuS8VabU0PBPGQtWfuTlItRNclh6gMxKQ80CStpRw+QwpWfJORwX16u8S0A3zE
InD4OqvFPLmesOTJKCDBRQRZ+m5UNMhRkU6+nbS0rrZBMYtcCvmUwgu1PqTLB08o
j1jcJIC6DZuZzZUJC0kFPu6ny4tv4TeCAH/Ozp++lq+++bXsQAKUQv5PnZ08ST1H
eZyUppJ/pRHzcigkSZorFj1AJBTuVwLJQ1mzkgU53mOI7bPGYvPTAlEtff5ALRNJ
iilJRBZRBME/nEvnIGAvoC+xLe08KskGTyMzglyqmEhgvqCDXs9iqUj6BxO99Qhl
3poIt8GH9AEX07Etrdv1kzE/l0S3d8nncjEji/5cfPLQHm8mPbgIOLn+TWWix+/v
iDsW/5MB59JU2kBMKow735GCZiEtAnOBGmTpWPoVNn1xv2cJ+4cZaMsiWRz1x1fK
Uh/2+K5LxwKr5xT+5dIhTjnt3oKAWsYrOZZVk3J2vRFszZT8Ij5j+Txxo0SXagUQ
GeK0mWTUBrcklf6Dwhyz+n1938NKAzsnqA44FZABbGqiDJSxBII3HOUkYEJApHcH
8n64HrA8dUDf/1CbdyT4z2rNnUfJjDi90v/WwksSn/z03xHYTTm5JdZ5u/POk3sP
49iMVDabeHlow73R8KtEbDIkPb5E8xU36m6nAl+2LpNFJmP00roKf1KCJjJeA2sk
GDacO6DwrzfXWEj7pyMIpwaefDqJjb48IUnSNmY4WbFXmGXrdNTF0kJ4PcHZeuVU
CFgj25YfWGr7UT3dMSPRxBmn0UUbqYfaofUuOKWGeqiLQuhII90juXFa3S3ExZRx
LU2cKvmoQw/mRSyD2Gnttzy+Y4qwkbAhXJ6ACk5mc47fR3SsEmVPNLMTeGFV6ekC
v2dvBT3MfdWistYzDilvhOvMKrTa8oF4kxJmk0tmEuD/Hg6Il2u/FWQHaxj+uioI
9nIGV9UcDVDi3ToE/g2Tr1etTLhUzSUmfjC9JUyvazBSag67NzhUSyuHOy/FUL+k
9nIGdsVLf9clWiv9ajzjcYdEf1Mj2Dvz9Beq1CwHJ9SRcn2FjE3uUkFsEbsLgq0D
s+YeO42ARID3ERf/VcalClrHbuNilYQ8hDDxIIQzDcsrypgy7j3cBcYkw5lalRnS
mFbRfFN0U8aeIprGQYxhKBVxMs+N4yDnxseMQLhjfhTactZ494qk+j+gLIMDrCEt
MgQhthH1u3gU5S4gYaAxl1W0qYz2876BUcrY9OiQE9llUUoANgfZCO69iIsab0Bu
473s2nzIFfnlMV7L21YW1PHFH/CISCYNN9DwXMZ/AErkxeIyOD6hqjpzMRE1yD7V
gx/VU5zQjS+vd7onjXB6syk+NWNmfTJLZj3eTB9vB9L1e51hCuUFFEvtFicMDQUW
y2lKH6R1sfb+0ZWELCdRQbfj7CpSgXuX9leBEA19YFNZLqfKtmE6Dn9XbekasBuj
qf8ji17ZJ5a8+yJPVkGVehIPyc6ra4pig1HIaldR29AUQRcj+pmmFqWuF2HpRMx6
r0WGI8obngIu1rYEQQDnUkRJRA2++5vFTZ5qj/vi3+PZVgEtCE6mkRvyUbE/aPe1
LFRZiIKrEo+WYaA1AyEtwvcUiG6ChUmp0/LNaAJWwtEy/bC0GPiLl0bTK8IQxeAo
gTKhMy8jrvlABWMIUcu9QQCYryU6ny9dh5mmygUhnF6ows0GI2QR3Ly5seWcd9he
/imvCDDOzSF2unE4WwvgiWPV8g3u7YVw+Ic8K3T5YyYYbCKqk6XCzugXdEQWL3wq
HJysLvoIbQkWjYEjj6x0LtdPugMfNUTlBKC2g0VUpp6uwZq83hJ0RHwMKmB1AkjT
Zj79x3jCzsRYRE/b5jUgpElFweB9uVsmYtkKfSY/3YCtN7KYYgBw5pp/BjSQHOiO
rhI4vyqug8doZRTGtbHChV8eNm1S5Bh03ComOAhqhA8Dv51ysPlNDmwOrz0mXxkf
mMZCUTor3r+hL5sidSIslzjk/EW8ViwZU0KtMA3IgcVLvKB+67lYMEODK6cUHDRJ
xGydP5CvTC8JZBcLgrbSOFEQJ8rSCBGI5vhTr7KmDu9T0yY+ZzORiUHf0KxUpSeQ
/tSQxJn8gkvLw8W98w1O1qXdTA9cr6ycXhOBGDjQ+p6OGOExv2g44bnfzWMi/htO
a4MK7gCZ5htWdIPA0Vx/or9SHITujTI8GGxGpryIGwQSVDn6iVr1TVzUls6pWEtF
iESIYrgFHGJCpQHF30BycQ1yUQyo8TMP1PKBFXxMJq0tR9hHTWBT1OBlEW3INRFL
aZQ1/pcjE+/7ScS8GlSCn7UQ39HTR8L9ZCo2aIjHcPzwsxpPkdNUZRxlsKoRrq9R
snKtfdYUPnDvcBEKTvh2lQt6ABZX/bG69vkzHGDWsroK+4euN6+7JYyR1XEaX2Cf
LaUk8112044+Bw3z0KgyayKTLxv1EkB07/3FVcKLCzEy27evjZ/81Y3HReHvJINw
w+1eglpakZgt5X+nr7d19962sa5Xxre88BpPAHo7ofQAq0sVoQ7p7MLsFsWr0uUE
8biSqlKp5X3i5SdtPNB5SVpI5SK4G3vWLEVIEbwA9ytEYTsmtR4J0DXqUe7SePnH
t4x9oKYKvUo/L8b/AMKpxgJ9xvgSoFeVQ3Lt3oYLpFEUUWDBZ+BgeR+zQGEOHUco
cF/u70vOkINfCGXkmbc3+qEeDFohl0W9UZWfM2djfhkzXKR3u2OSRfaz9T85UdB3
+L7UsTxP8If1K0bRijNPJC5RqDLIrye/n1qYCrnHpwEpAhDcQ0j1Bqvn5spzWzC6
J0qYb82yqM6waignOREqd1PuMKgdLVxCDA4ZIgzLifP2AY87+Bt79V/pbdZ1gaml
tL3/CLcNeQR5M+FsXcF0TwvBSa/MQUq4qFcBbq44ZvooW2xkwCpf45TLRoFX/5rP
kjsd3FkKGOCEX+X8+JkqqfuuGEX11qfOWpWt3643Dz/Zr0P3hCrou0u2bipvJeR8
cpRorvCI9t1m7SlKH8XjotM4d/l6h5D8nUVCYqEtj5dT9mQwMHO1W3spTbgBs0iD
FUa/PEKbAcSnGd6sSkVEHz0aIwFqy6hdkXpH8fNqMyC6+KE+rLbe7Bdf7FJHuXIc
7nirluTyKM77HiMcCr8lKKP3dbHtB8nJnqZYV6Wpl44sCT+X8K/osgjVHgXnD0Gt
nuqKf0mBjKd5IICIwVhH2ROvKFUsE8Nf55JdtvKO+zD1T4zn1ojLkd/oFP//4AJ5
gdaLnoMyUk7fBBbOZna8QsZatbihDhrYOl0lKMiTTNYPYMXhdkPe1bV58cONnltg
C6rMNq8X0/PcB8ZK1t08RN0yfk8Tlh940Gc5RIuTl4ttQdE6kzh8Hkfk2e7/kRU6
t5LwT04qgVI4CRtmuNpNo4jpOqvOMraOUFGAP2D5cxAsqsHJ3xqU8Ufeb4BhsDHG
DCJOkPD+ZmcraJrLoGF8qObitoW/pNpi23i2uvifRPgfkoSbsHaheAiAw1gT0KRh
LfYJFkoK2ycxg6gC0Dh4egtn+xGwtQC0V6R+DV7VPbylZgNunn8GMOgwfl757YOG
XKM2isOBVk7FXYbn5DTHA0cWHA2QR6Noaxa3O3j0Q/JzXyEQtK9/X0shhJalVYVd
cSqr+aQH/wTUEUnqsvGQ2ayqoyu5eKXHzDGeJymRiJu3S6oMH90bBCXtN1JFBz3U
lDHocAFHBjJCk1LSUEa9PFfbbJ3m9h+RlKUKLU8dfAHF6puqFLR+K27sh5CUxmIW
Z6qY6GUqU37KH+3xl1iUn8kWvRDGDaBJSK2WtyscNdDiRuFgd8CpAiXtkTXFvATW
a04NEVQDGkqf1watTBAyPXmE3bQ4wxIXCHjPxjzGYcTWwaC913RS8OX4xhlWm+4G
jbiJDdy3yjaJVSm+Ha0zod6sSchxhGAiyaTPP/CTJxZmZ/V/9PZowKz0Gva60PU3
MdlrBvSDVE752izURw9NsYHh2nqOrveOt4YJm1LGxmwJVYNJ8KGbAD9z9rmudfUy
Qy+quVtQJ+aLt7iEDUfrRo2bES73mzagWwI0I3ah3dvMcoruRsDRMAVk7ml8NKzY
yjKdaWf5/v5EQn3RdhJM+9JOHnX6zPb/tvTEbY8rYl7buO1aG3/WftuiWhZtRRUa
gSaF/8lklEGndrMyEOKJX/thzvJFxyJb3vezhShImYrXRrJ5IA5KOVCCUEHKOsKj
GCAtjwHVuvqbD7h4ZnO7zCvzEyPt5f3NF0VVEjqpV0QMQ8F40cmy54k7nCYvxyRx
y1LV1dwZCCy3lrRQHK+4HaIrx/0V8SiAId/Z1e7pVr6NjZfkx0gHGfOGDQ/F2T0s
hDVewhfhSwQYnXUGljeEMrcrgvEao2/SfVBIuBLUNEo+Lwx/MAU8frhVzFOLnfhs
B+RV5o2EJBVrrb8ttDBFqXiPMzxX8mZ35XjLZqf47fI0A0NsQqlHa6pVd91fbFjV
D4IdljJeYT/3/6yO1A9pJCbHDhCee6Kywz1bRrSc062SkxgexJuDZXeCmEXfObpk
1yqiMxcJ0FazQqH/swhJQSQ3BUHCjU1h6Z+rIpa/n2EI8LyMSsIiWX3ipKWCc/du
49LWBesZeddqwKN7qR4K6n2keZ4jBjp1pNL3CYS81wzJqmxwuzoBJZj8KpNPFYtU
zQknU2wKU/XEPkbUkiCeG8iI847uNYqJaYVbsuAk5txXNeQdbFL203U2AMJWFZrr
g7uQDcu+v8fat6d2qJEpS84eghsbhGgBUh6yXPnLU8o/F+rMwtY4FGUSJdUuWlGs
jENDbNvPiRNi2uyXCNfap4xVtYwq36+CFLa6Kna8agfy6W9IHnWYGBj+BWlXwWds
FXtq9aOELmqDeSV0c4tGKg1DRiyKxRpWx7kqTPSEBfJsBEprAjf1mVsKaeU7NWvQ
6dMf7BzizJOFrtmQSjknTcyfWilNPcSBGxENOdDlacVTi2ohIEwhAtwgJ3jaJKXn
sbwcAhXt9vE8oxAod6AyyWk828GAZZUhObaew+wzQYFFPvHei8IZxKoQKLKoz88L
wKpBp3d6YnnxSB7NYluiOvdetUvGPu40O0MAy6xOAuJVhGM2uZdmok5G/3pAdCNB
yiBWAveSa79P8Dd2VMZLhQ9ZRpX5dRBQUJDBYalMvMUfB59GLvdmPXENklMHC/Q8
1oYwf7ixi4Vp0hS3IU4Y9YunqP79vOWTFjxC/0SaIM59d/K2KPdjbzKm9mEtEZs+
Wb1PrNkFqv8ryZeNyv7RvnlS8DTAYUulY7JXz+6L/dDT24yh9OVOPKtxl9Knn6pK
NrRA1U1hZAWxcuk4mwT3qGdcS6qoYcKFiANd4fY+L91fkAJrajgZF2BbN/p6+ETn
f0KJCYnMRDVVq1i+xDHR4wBBDWVsg9wOCirmTmWlHAXB+EZoaUVKE4DVO7Uk3wLS
fj1Pvi0u4ioAVolQe4LrzR1dwPBU71O/rc+9RywzZZTqCoY0wjeb/ZSRBzNdQlSE
tLSvPRbxICFz2AJoaVFoY8ziw6LUElJjr9Hqh+kjDGfQph5ICyFKKvdOS684f6NG
dWpgT0Quwnn5xR0yERTv9rdbTxZdlBfMp6U17X1C7GNqZ/sEAIaScz11R+UfnFNk
BqonScwZSAM9IL1mghWy17P5CC4b2COvFwsy5nfCxN3dAJOZN5S+dF4PAaHu1vMW
Nk2DQ9EwkGeBZZsItd1YVcNK6VNPWrqGO0r67wesUXRUyr+kNMU+SN8uPR+KFg3O
ZXyQ9S9o3ttADN7UHCOH3dkSkGSO70Rn4GbTeQwVXvssF3qf945dOWXeDHeMiaBc
o3A8xRI9QFqEZZCrCYV7tQP3w4FPICge+gXAxXPx4CH0ZjXMt22UTqUq5y+2Zqj6
eHxCg+e0tJArQXZgDlcl/z+obRhTlxMfZXz3GlTVVsOYZyMfNbw0eHMky2bPsOjE
cS1gBled0YT33gdXGVmdh3wvTozYdvjwtY7PpkL4A0cy4yV8Wy39YuesEsBYvFG8
dVgSBcu7wNGK9qiTRMnbVpbEg8tlelfrdOONFuQGREkebk9XZNXKC+sJhefwwmBO
TMFv8D3H7taxQzdeDHjuTO6SEzii6/ZYBFwJmYg/oTeDbDaah1au3DyuUOq9gsi1
X5+rhfZPxJuJ9qlwwVHxOraruvfLtGsU3E0253viUZmGSYX/ucUf5dLVRfNN141u
3SKQieLPHWRjGjgZ/0Yeavb+mHnfHL/wvBVX7/VOc9jb4O9aA818+7X0ihVzXRpZ
9WIvI4T+6/C7GVimZoGdONUiRLmdljz7XSKdKDhhibTkl3ao6xnwLGAIpSMz/X0M
p0QW0uqXxC20/iE7CbWvDGVlpoupyLa7hWIiuQPf2Sb+unlFKzz2N4EB7JRHvR0H
yEsJ+6pogSaXSwY6M9Wu4tBJTVY0aVRw0+RxVitMVrri9bZ5GVjViaml3eQ0cQaW
UZVf0ryunH/OO8dNBg0n2VGfBrxfb9Isr5F/7m82ap5SL8s5Vi9AAAIhQUuxKwBc
pij7sOfeo/C8RA/mBpOYY4jbq5vYWrSsCA9dJTaoB1d/gZwMc7jF7s1cdBncAGrs
okS2NgFOXICvtUvpqhAEMp3ChhGuuHqU5k/5f5XXnj/9LHlIUJV1G/YRnQ3fru02
1sgk0XaXpTkTa92koag4tkwozWOsCYKu2z6NujShJUBcxL8MAXDm6Wrwjl4MVDEu
tLGfeMfeMqRlHFIQL51T4GVGNUKGQu2ThLLEM3vetkow0Y6/DrwWSUz5trJHUQXk
Dqcg8zTH23oQNZC2yIs+0pvefQbb2SPwwsEOtMjuFHAigUEkKV+QMiXZvZ/gcfr0
izov9ECDkMup61XjvaIs47nIcwnUqgMFerdQOETqm8DkM1uZi1N2CPySWYZVC42O
d2y3C9TGRHYM1wezWS1vaj/o2luA04R31yLba3DO/QGM6em7+zWrYRWa9ZTS2Qh3
T8XPPfqcm4yaigb1lzPfJJZdNup93pxarvoj/33WdVTcEc44Gh2Mn4YFwX3z4RcC
LUvVo4ttiShmsh5LxNNxD8GsQvXlKCyjQEau3bM3+KUoc+bxlt/Z36waPskhyLs5
hDDNJ/dUbvbZUGH/5UrcjRJLA0vYdwm4plcDd8V7wiNj1jbWoxNaS0rr6ndbYY+o
qhSWqlf6hdIJG5YMZpjPnkbue2t3LT9CA2rLnfyozzZnjTz174h/eSoajL/TkNFI
GStNPGz/7AO0gjXMqXNHFmtWejNmB7nADJaIlSGoUXQ84kSWyUpacca5FVzVSQLw
SXkPFPqrg96MPH44eWKDHaXMs+wEOLkEBmeRVSg/MWEWNnIdmkFUQO9ujKOghivn
0o2Su9Juxr7nO7Nx0eIFm1kX+ZZ69/o/++z7zlG0Q//xq/rc0KE5m3SMx/pmU9GY
U34wsxcWdkJ2/V1L3mQwY52QJh0jO7fFp4JkJvB775va3RKM/QJtcgEaxCZgBSvD
XJUcxlD9/12A7Pk+TBb9PdEssTK1DZ1gD9+/RMLETt/5R4V28A8p1ZyjcxTNAGoq
re09U9lto/0V0nZQuHp95zz6TuOhQ93YbsKplT+wKYqeYV8Kce0KL+M+H/OQ1Sv2
kyqzftVEN+esrDKc4oH1fjiFSLvfWITTLfhwvIoj2/TA6z4h+KnlyfJOEe9yJIsp
nVVYrRLCSBLmi4Jz87MQpo6o8zAckYemvkzYO3r780coRTZE+voYcG1zOKkbFp4a
dtcUZJ/hqcu4xiZOTGDCk40eikCUKd9VYKP/eaj2k9gX4ayWTVf4RqgARk30sXOz
Aw8qUMx0wWc7CvlznBIiOe8/B2Jgyp/Ao8IdpaZDSGN6RluTujNSahmJv0PmC2E4
5xNBEspnbl3Z49NnVgw/YI9KamBm+WTKqK5sGj8vCdiU73cLJaWbY4M7P4ujasHT
yUsOhRzv9B67Bb3fSfGxO247txwtUKbPBryCkgEleJ2p/2zkfDw1EDNXehb+NgVy
9ZkNuEnlTO8iX78LnA4dT2LzPXWqh1tv0a1eLOBgwypp8g4k4MTvGAxXXCtLC4QD
CaWHaO8jpOwR0ORCIHS7EA4cyMOFlWxKJGxYHcs9V3p9dxNtL/zNEZ0lKcdWcaj0
vxwcwAAi0zQqCkikqcvCtllz76MvRCw0oJNX/3GzHacm0O5ZpSjh22N4uFEC2icr
w5RSPfylTruMBcFqte6jMrajwDvChkWNnzUqX7jtBkPqCa4sW6f8y/W91RamUjm3
81kGtEqU+XWpytFnLXWjmOXKJuld55XyxPkRpMN18VQxQJs+9PPz5WbHreusylXK
epMs80SzRZ6z95/xIqmPdwvhExXQOE2EZU3pyo3v4WYmpg73Uj5PbVb535A8n9ne
B4y0hyablOD3NmjekBFpRM4T6oMb8xLXh9SrpkmfZ0Pwm8n1F1vME6LBF00LWJz0
fH71lqmzby341LMvGR3p6wK3FRuS0z9i6b4F9o9RCytGTYvnzbRxdsQN0BIJTJvD
FZ2OofaLXMtdcynF5NtzS5GgvYaIolFAP5vB1feJuT3+PtOOFg2I6MtBay47PdDr
yz/9lgI9y7x36leFOXE+1WmEsxE/8GcnjTprULj9Oue73kQxOllUOceWPpNum0Yz
5PdogEXouv/mjzRI0mFSwyHKFeoCmbMxceRzOK1x8cKAKOuxB9R+k15jNGhk0OX6
vcmoEwm9hDw7SJ5PbxvAginde2vCzW6nmyxo7lZ9kcGlcvrM+l53uN/CSVrEUowt
Xj8MRmCyUa9ZRYU3cEj4Z6HE3MZF1pyPl+t7N+jEPQBa0QctCpnousF15BwflcHY
suAhzHCBHOw37o7Z9uqri5ZTv+VM5wJY2sT0PGWOffuOFQ2ilMIGQECFylT/c2wC
S2KpSjU1mCOdaBr8ulUP9qoONcg5yb34YkJUdTuZgyUyEH0nsWl+FdUlMmhoUht6
7/0Vkdk8rK9+678orjRtDlhobWi+Fpol5dG34sQ6lv3paqtyoVLmUC6bu+AMnq1E
+sIRWS/BhxeMVv4ye0xVDDxnENyhfOmLqiwHmwlLrJyl6fm//gZUyWiH4Y/Tv3vY
trMfsSSAZP7XPz4AhNgt+Rm2Z6rWyBavitZkqGlJmqbowwS6kxPLE2dqvXitA9Hf
BALUkgMSj1JLs8OEXxKGjT7V9QXRy4VXiUmHZUG0p3+x5OeujiJRq1OlwnNVSv2x
KH4Ki2Yhqnq4U8ht3hoEM4eX0/cCW/4HVD9kBou1jqZdKaaRhfKpBgwA4k1OHuaL
fDTL/s5ZwqG8KkykZLgZ9XIF95A6QuF2Vqfi7fIHP+n7rrRvM3lcObk4hp/HMZqV
LHznAw4O3Dv9TokdLGJi4IPZXajNd2ohKO9CJT+v9T4ffxMrhQhpC1NPA3OKxfQP
P6E5hEOG2QbAmRfeRkzyMRoF/NAgXgiPg9P8y6+yFLgkkyIMPyWDdmlZyJYZG6ST
K3jiY+VQDmso6Syd/1ZQmzCaRZr7qCAdn2CtNYtid8Q84ZSFJl/4jpRj/B6CSGsD
ZY7gGizdwcelRfTggPsZVi/dkKoVScCuXLdlZE5TtUJrZ3d5OpqZaxtkzV8gcJqm
CdBieNRMo2hXF/AFR0/OTx5knFySNKs20Anxydc72p6BECDLE1V1/X2oEMhKcyyl
dC4VzImd5e7eingqA50twMY/NnCmU8U3i+qW1SolQefubLvDyFLSsL9Xwr4O5qpV
Qz6cOvByCR507ojfSnQ3tAfsHyWYrnpolII0ogg4gtvJp28Hs2i7QVLOIMSjpkuD
KYicl8TA5qWEaeQXlEvqPYoTgD+WzqJNB+trRyXIYO7xGNvN7qc6c29ZHmpviKWr
balv//gDgM/ZwTV4PFiCAr6NIsZBq1Q91dv9hyBDFPMGTaSELGEe3nWZfFgyv1u/
9LqrwmSWJ1f6OKZ3L1cDoRaJeNEQKVyuIYDPTj84onUS+qMhFsC+Nw95NhQOwIhc
ar0weZLwS3TYKV7MO/yLUtlabBUveF3x0bd+YzDoYZ1V44/AsUjiRGlEwWkcmlCj
/maqctRwDwbJILhu0Yb/s/yFPIoaFjPhvaIkJczCE1RZ8hyMYtFLnOnN6w2D7kdq
7cvlnDjWdz1AV6SiOYfkDfE6mf+Kay1Ws0k3iuw1/VAMiO6eCRPvxpIDdh2rIQyt
cru6c10ErT4+KXrw2ZCjASIjxiaYgfQjreWcPl5ccZXobBLxIEE2FGXHa+rVoDxn
0fZm3O1TubRoLlz8DvttdU7oolbLnH3FuNCrvdmFe2tCX0NdxGOzqQdNNCndLSHb
ZRwC7ejJ0+16jG7KnNtCPltt7FHwNdU0D3TBtyC5km0TC/7ei4gOP+Dtn3H2i3z2
vuLHk3p7/Rxm4EpSU9iSIg5fdRIT5gEsYVNdSKwAgo3dN5dqbHhogDIclWN/QkCf
PsP8X1BpD6uDxnTEBA9VWXGQNd9/rX1e0cGG1FyC5F82w4bJUOgmZtpXccmgsEe7
rccmVyw9oEIIbxGoanggwxDMSVnz5DmpByoDi9UVgkTG9LVQa9rKn4YCc+B+YT1A
eFMjxDNl1f3wzcULSJxfpSegTVcXDR/dEjcKk+COx7uamdHgEsq+d/Eqn2VhYGtO
Orf/6merYnYIggxGaL8bf00fVB3Y6kscBLEDTr3DKbFoqDXN0Dxo1+ZJkj6zHCBQ
ShUa+8qsH2J/rWjmoKgNCl1GdonTp3yB2USOaNAuyaYuR715+eR2cnfb3A4FdJSB
Yw+J4oJRMehyMCPtwdny5wYdX980R8cnGr5J4M6aNeGZe9pdtF9g5cVe+LO4pQp6
QIJJsoHeCem0bHCNneV4FhtcAH3HwmsDNm77a9xh9vCbd0bqHgsVHPPSvpqy5CQx
/t/c3pcrb6EUCpzYPlJvlKSNzxlggk7ruGM5N/1k4iwQ77B4SLsaGcGGN4cKqw0G
p609rZmCIKOKG4uhd+2y4HOFFdnBkZGOmRNIgIJkNVI8xa3BrXX6UBk5Pm5b1VBE
oIJLJHsXpHYoABKMXO20J+enHmsjiJtGa6GQzk1ayBwxj2DEjz7C+761G4M2l/G7
saye3tlDcZNiLWLMnzgixtyIF7D77erfKqFJo4Qo0OH8GFlopDv9uMw89I052s28
xtF5n/lFNNIlOSI5ID989zGiBVR3b2zIdDr/xuNi0vIzWze4FPeBBRGv7oULNEZv
V73D7/H5F8kZ+ZLbfZvG91s00mHXnNs77i2C7o9A3z/cvUehmbWT0DIoz1Wjc9/a
oSVMU1cI+tBQFsyJ6vScmzZdN/IyaEP5UF2WT57zU2silLxXVOfF2Ehdlos52nEu
/7u9e/ODCR5cl7sA6y5ZlAbWIaEtdkZX2gANURsZShTC9EdSu4n+ynVvr3R4/ryM
GBTHPE9PLBD7H7t6ndHNJGfTMc+tf3xoubWoHyapfFBACEGm8D/WZmy5NNDAuKpP
A5ShIJ7u8tnsIoXsjOKhHGjFWwlga+ly35hjvsV7ncPf+fMgP/2gGQAZrjACUkF/
X8a/ZXth0iqwZhiSgC7XHxSW9LNLozGkUn2JmkUV/AEQT8waucIKMs/8kFcEgqWr
T5Hge4Ig5ByoJxz9URHHb+XJngzBZXD7jVhH57LpYjf2cQNaqfLN9Zsd5voaCzkG
ipLIX31UnT9ftwGolxusFtWu+8kCD8QcOh8HMMLUoHjT7jfDyINPKT2IoLVko241
RHveAc2PY5uwOEBlqW6CmloDGnr/HklxY6Ve1g+vGSqfoS6020AJIzEihka0RbQL
GuDggX0ugo9Y+8cwtlatgDRHv3qlHxIxEuYrkW/9ovxZsF9Wi1sJiBSxL5y+m84N
MvFTNFUmVPdZ3pyWJyYwnET5u5z2UsFz1Rd77BRRiwa0dSITeEOAxLLf/q5/dHNg
RfVSu+fyhB4BfgwhIddEPFBklXAqyEDR4mwHJlZuO64JsdVeKdFyEK33IKv+Mhb7
B7x+udm25zIAP69MWyote6jYwHN4bhdEb5MNHXpwVUqxtpv22qfjegoXkw4hXckF
Q7zKCAdTo4oGW17uwNvv6kPK4YzL23t5fXDq1HeP8guqP6je/47d5LlH9egrf0Gd
xKvqZDFmqUCdU1aSwZd0N7MEdfgFFubimjbNe1TJH6sbH1XmoVSTR2mwO6IIclIK
ID6lYoTEkeAke1OvaNzGxX7wzuyID8xSgSlYDPHJd0KIMINja3qcexAHk1086wXY
OhIWsEjDBcYwMc9YLU5cM8DSxxaMvqChQ6R0O2dt3hWQn5RnPVCPKM1rEGBBglVN
grlwgFmsjVpb+Xe0lwAeqxYO9Ac1+mvt9cVsOcPv10wRDSSOq9Kc6OJw+Y6X4Z2i
IvaNinPNblOs7rIOP2Q5YPVc3w9o2IoyziTQTugWhoi6LVScAGhfegGIiP8fXLuj
sWnqb7nWgJ3x7SPA5UxOL13lgMtBKkJjOS6Jc1xll9hyLdi5YV3lcbIl+eEDy38o
+IqALWUFkjgK8e/8Z0p8W4mR7MDIN/5zl7D3I7UyaCLBk8tZXpRBdYeRdWppQ/iA
/b6yuSeOyq2oPSqsmzeaAqKhI5Tth13iTGPXGUv60at6GR1rcgwK+wYYISKKbIBC
gmTuNd3HnbB/BRsXvBwvzkD0DTTNmwAfdrLiq7BPgg2nHHehBTAyuEZfWdWkkq7R
TV5np2CXYzpQcxgZaSR9Ujl2kSKj3AAa/1I+8/aVKpCcDIoM5tGZ9/fjZ+H/ypfU
4e2D7ikmOFiVOH8av//QBbQ+XxqvFYJfINaWPPMPDaoSRxr+Iykj9S8/njuuekyz
UvZsXADrxQgpeWWSwUe1UgttLBqfaQxSYE/WR09QPEWeUg90iPvWdZ7B/RaLJPiX
W/30v1mqJ+4CNUfOByxtRxTN7o16DhtY/bRLH9r8vkXE8Ub4M28UYMkJEXQp4ek5
xP4Xc+YVs/jbOZrChiz2/uO2jc9yDg9k8Y2KdNCMiNSu1XB1b+E2bp4zS3Rsuryu
kSyzi/5QMcdDBcqA5N7hdQIBWHF/Vb0NfsXH3Nb93TvyvF15LNl0KuCZQhxT4GL4
/lecLeVLP2GhFEutKUeR2SSKfb45BcoHCZpaoNoQo/qK54UlHsoW0jIJ8KKp3NyU
I9tX/6Om6LjK34cTKCuBcaKme2elqa2blS3FC7E5WU3+sXg2wYRhUzisTnUvljoV
67JZwg7fU5Qa9/wq7ccc713Luc81mG03uD86F5Aks9cAUe9rZlgKbWYqb+3XJbr0
DDoL6dkEipneHvuunfWhoAFVZBPfztZL4S59j8HjCQYonbC9udaLkpJZfAf7l5+g
UuuXcsDQBDH5PSlMMr0MMZpcTky7TN6lAwQN/AzqXAW7AprB8zNzHyupfOHXMuOt
YbagMZ56tWawtQ+BA5/4i3Rs53nZOvBj2eIjgUqxEVAeW2vUMS5R7a2N+HdBYAya
wZ+LMDJkD2Sen97mDQchHs3tE2i8CIr8BL/yHqqzqXrtOYlxC0SiwEopODpN8t1R
BPpstE5rvRr6axpzyrjX9knydVh3lyGhkqCoFtruPbUh2HuxPFrWvrNw/4bNOPx6
7C9r3VTTe/v16ONX9oZRB2tWKWgmPYWA5x056VKrt5bZEomxQZCwvKDzktRfh5IY
POvClmme2/uKBc+gADwHO0T7812x2vzLH8J7+t7Y/E0MN69eyNIDl/ZHHjZb51ox
RQs2DIYG7uQ59f+RIrx6VFPtYIHYvLzA/qwurnvTqMfBPZCpRyuwpwHDleojvUTO
ybzRoCxuaWgZd123YTCNxOboPhNc/UY8uF033K3ZClQD0BaKatWSKK/8QUWqdO59
XdBkNU2WezWZAPh6iY30PI2aXbNoqABCB+TnLEtScfJWkRvNF3q0y02DOnSFYZry
zrinlI3bOpUhbkN6ALz7mKqalHdrfvBOmW+4XvYyyznL+RnBp8Pr1fhEVz/MxFFX
lytQhMIiBqhSnEqNS8hffOXyk1FkZ0xB+/AXdh0H4sf+osFY35UFpy65ArLgnI7l
ckyAh9CLrVjjRBSTbEkEKRoOhtqwoOWgaVYQ2Ix3RMVpavCZ1JV3TFzQaLKDT1xW
w9AxLak4Xle4R+g7mu5w4DvFSi7RYlM6VCguiopx1//s64RUXujjvZ3Zt+To1CMC
PEjNVpCWg57+E3Z/SiZkJkEYdEVtBq8O4cMneSJUqOcBpQfAbvP4O58C2ScsOpZ0
mYi3crm49PIV/9hJK5vi8lEj/UMcvm3/TYEeHYEf5YaaHlt+fPb5P81FnUBKH68X
0XHufvujG+n+Ug0dxPV/Zs5J73D2sopqSpKT/kGIioZz/O3ZZAQrN7hRWii+oQMk
NMwS++deR/cNGPxsxGCEqKi6NaJwSzwKcJk57ScWierlKJb7aLwoVofcIWCVt3M8
UjlYnKaQIMkllHW0lHVwciXMpqRAx/Nwr1NXAheRBe8JNQ4AXn/SJmMsphEid4Ld
cXkLwbSozmcLnE/X5FOpA/nqMJK1+n+w5z1Z3JH65sSBW4dLCA0F13fDwqtwTa7h
oX0hy0nymM71H9aoKPUHYNS7WWqHxSSFiKoobC79byOVFRaqO+R5H0XCgk1e26n/
YBtLsvCvkCUeYW3FEEWncddeXBN329jsrXsZ6oXgONhat+JEwbEirZ88o7q4gLYP
n0xN7BYthfMxemLlA5Da1P/JHBYUzZM22L6dDeBTfxrmehOyhtnRXWcZEd2Dez8B
cyldNVSWx7XdhCr3Qwk3EkUE6birmi+pRRdv7eloMT02yWBvo+ImCMgPjKfmxMny
LxV7LwKYbT0mFk8PPj6yWTVBE6YFE7CtqJRed0og6uim3Jix7vcDg6dsyZjeEqqj
ZWmf2gF44jU9uSmdhqZ4UkpRFCWCBnMXXl39cTopxaUFDTew43jlV8knidNeGXgI
7OLztxUxmxRCuF1L9g6BvYtGXS9+9Yi4cJGtSGAbzzpmpdMKQoiWO6qdjKJ/OSru
w290TPh1YGfP9aIlH5flnq3K4hwWFFsU6+VqHCDx8EKr6LiPmJhFz6rnsWmHtFW/
buNYxIhCxxoKBTBGuToRUGCZgzZ1xsdIGLdeeIkiDGGTdAbIUYT98P+8uaQGjTbP
8cpUq0Y2AlM/1W8+MQC3+1gb1CvE64axiDpQB7dKfZ+uDg329HQ7Bwsy3K86WWP/
RJCnbCwBnoQwmCisuG2DBWiT/8RFb4D3dwPWf/dLBovCJSgD+DfVOQoZWzE+hz9m
Idw99bX+2/hQtrFK+BOUNodAMjidwSuG+18DhYegA2G2j9cpooxnE9gg5N5lPnGx
yL6Q0IhscM0Ag7ZoUwRUL5ccGFAGqtL4Hlj/7V6lhTUVTbuyWk0IOkiDu3ANKOFX
BVwagZRdWxiYrlpm9ANLLxH7itad/VqiqjnTEJ3lyabomHMdrN7CArXR+AU8rabW
adlk+gRbiItKrQZovHd0puKFTN3HqS8M7i5D7WlBbM/zm3TmBhs4BgPCt7CCdDz+
jpTn5Ts5pu7eLab9JAZZ5qauT8T6bZ74Vw5X0ZGJTwcljPwMlgRxH7H636h7EzcK
HJw/5ej21Oase5GXBSmCm+6wxJ+L31VGaFBtUHQzSwNeZ/ss+Nk8COi6ZwOs5pvN
dbDH/hKuIE1Yqa4EBghbVuE5Jo6UK/LvEde6rQ0NOFnx4/cBbDjcBQw6+zNAtuab
WmpqVETGNCKP9ulvU+RYJwtiwaZ99FIHPazK/BAWlJtNlSsqiGwrEsHzr8XEHPMq
xAVdefUJL67gLdWzDOyDANf71Dh8MECplZoXvnVY5PStUUW1ZLzAHvdtNQ8KNl8v
XCEAcynA5QnDYlzLfLhtpOMt0nf08EGuc1xprpSjvkgPNziG2M+2kB3Gd66q7pRk
oW05duhV803B4UyJytECTnr0ieEvu913xkxzHmbavFfHPgGOextm9MBzeGFqYO8+
SxEFyTlw3cqQjZxGunLyRK+37npo8K2+8zs3DE+hILWlz5wBsI9hVJGDaIokIlRV
Bcstu9jAyNuNvNNd4hvajX/gJnNGZj56OyD3f3UNUf+vfDY29WD9IXxRFUp+rseq
tx0j2H1YWyB//PCnoJONC8aazA6cj+CVsvR6GPF4RsJafWk75PN6WXQwcKB98ktG
2LpwyzOwMIeqYh02cnkSUPJ1yAgA4K/iTs64cEwF7dqzOvRvcngaH8Fl3mQMxEd1
1PIvP/4XV8VdThJXaMt+lPXvGqfqc0dX5dbyCWfsgZCLRDdqblY0dx1GRmCnO8yF
CFUWdtthbUbPprA1hk3QiYHLNydelWy9xUgobkaj2KM/x1ijchG5QTpOe7rEjNR5
smLmOc97w9MSgpZ70/dGANnohyfnvhSlpr2fZvdLmNwwkhxbISEwi960AojyBpG0
2xxREYwHJSriX5Q2z2iScVpLht512rHEIr0WqYQq9x/hhJcBNUHvH1DboIjrY1TB
DbirxwwwNXCxI1vKBfPVioe6OzGofT9/JZysnXUQeJqkVVRceggHxPG/2Sz59T/A
NBUwYwnLsRgtnNOrx3V6mW3gq9Z03Di4jnakO0V/bqahnCQ5kOVoA5P6rAhmAJkn
3wYJkGE3WRTzdQNVJTJqw4TjjF6rdkSWVv0OKceCXRzYFPXlVr/YDw3/cV2EAPaE
brSRRTHFLKUrnLNSo1OD+POOiFbh5qffAXYebYzYz8HHHKjd18T5aC5E4el+ACQC
cef6R6k5lRy5HE5dIzXK8IT3BohXq2M3c3/3jKDNH4K9MMSYjeNU8KdFkCI3nnxZ
SX6FCKMmbbKrLKpDOTBCYYQHOOUcrJsepRvgzxiFNiBKdNNEz/SEf5DsrdqJlBZ6
VJPHwNDQVVYrXclHVo0XGbbXQs956KC3DPwc0UZl6H1reXp8xgmQHmI/gthStjQw
+lauOpto2TSCUnbwr1FaWI2Kn69t1XtbAURouCRALE+TVe5s2vvCv3VZTURl9+8J
JOg/Hjq3TGiEOSmqKZidKrtlGJiKvk/ZPeuWZjcMN8ozfYI50LtOAOqmJLZahOUJ
Uxa7ccT/82TCjHRCAIavYg9pkMV+dmW0BVabbZSUCfIG8mLKOAB/S69W7pXlnO8n
WYRcpYb2+KFRB1a8BWkOTfH6mlvEsvos5xouXdy8V0fVFORxjAlmUtL9ZvKG+fxa
A35m6xi+uNzgPlotdBqBoJj4v1gGSzPwp/VGJlG8GBeF75T2B0aqbTEi5KwPb7Xy
E10wKq5A9x2P56KcLcNnQ/lavLQTPT6zuruvjMxORv92BGhIlXmvm17VNso1Lx1K
xdOYlm8xoIFuFZ1zVrrWXt28j5vJNhwutwmUFIkIbDgLQMDeV6aZzwtW4lNwjW+i
l3sVegGxxDBMc0AtKDRu5j7unOiVrEckr1jTFRt61xF+0fctvcktuyvoZbYwCfJS
GskIur9Vx2p3OtX9wWJM9hJfwBDmcll4WIW0zTtPJ9bN30FRwiNP0PChnV+3JFD6
Eo0zJKm/o2CXa4U2CGY6a5c6IFvbiXIdV40AH51ZkfTvkgs1zJUy4LagbnLE++kw
Hye+yQw+/QMMMjUMlmZIvfu5hoIf6yK0GBUAjWFXReU18Ts1QQAaHGg2LCruP0LQ
pfLgk43tQ0YsdP7yBvNju8uIFWeM9iAmbh08+gH6Vvwhce90frtOWHgDoz3CeMuJ
3LENZqWYsarevm+M6EB+Rhf2+gH8R3QNhy3u0lyXWJ1MyXPEig7fxx/zHQcHDJfL
WSpYqubBevOOEpfswtd91BZdZDZbyGJnLyDez/ykxxmrjo68EVJF3/ppar6rcpiW
DOLdl8Xcv1RUxe7I4Bg+61SmLf/uT8WBiMLRi6hd1NXjK+AkXSIlC+vfVVXnJYg3
4rQ+Mtf/PwlvLEW8wYtmbPXZzL/jFC9A4zFG5GP6TUSVWc5e3b1c1BErHpCdG7E4
iHgitl4xsOo1efkl41Jv5tKMRKKIkAGGssafNc3qiPI06obEEl6etSEZVhBxMv4y
UnDs5ScuknI0Vn3043roH4DnNzEevRNz+nbTk3ysyT8ewauTegd1vxMgLas6Jvjt
GhyDLnmhoTnC0SPGCR7Fx2xqsbSm+dC6b4gxHrfsYSZNkYPJSsJZOQAe9wUP9qHg
SRu/eBa2MyCFaLrKIPY+rVRjyB3iFxUvCAH7ODFcJO1w8yXWwoZMe5pf6MLDqlzf
7NVhY4qM06xSFenZ1CYgyUZXuyvEkTINt1qDeNogmAtuRua8Ncd2nrbHayas8ThS
4c+x+56egHyLps9H9gYIEKai6d6DKu7ow5EYbeucbALh6uJbOuC7i8MYr7tqOrCu
Qb3vjiMs6Zx9A5ebLyGI3Rz9QNFNZEEnokdaT19K6rrYIxMmr18cv5SZ3Rjeu6K9
RoUfEQJUZk3wSD22G5EkaROfs5lv+JGcRDNPhpaMY8/ePtTy+wkxVuMY1dqbuvxO
O8SCE0U38H3bP8sGOJfz8UCxzTAG6XO4u1+egpzJ0MJ5B5G50Oly+5LCHUF+CuD+
Yw9j8tz7jAaIgozeVyVPWkxpbxLPZtaXRMT6On9PDujcBGe0xxeUM7wARvOuxiKv
xXlro8mKClLMCkvHbeN6MH3mjMVqJRAv0LuQ+0tmmIYV9O3GWdZFPQ0qcrewWQjJ
IL6QOaAntiZlzx524ztkhzA+CIBgl/Wr/uwrYaM6ugr5k6qOhZ9dlfpfaYn5U8cS
IrO8RpfjFzSMGfAZOT54ambsM6Y/rE8NWeMb1gz8W8zGWtZWDkjKFiaqs924InIn
nZOtc8DVzrGWEmuDC4m828J70qCEiuaBUP7RNUL6dGSbRZuW7tQbZmX8Jinr38yX
KWCnhbzX7CAucj/NNLYJy5k1mJYWz0QJmQznqyPsn9TSTXc/OfNyGpqTCt4OLm7E
y9JAofjdq1QQpGR76RJg8YDnXe0uI7PFhjtIEAVTI7whEd+Cc0JavvGzMb8SMp7U
3Feyll0xqosKqY36hBuNNO6kM/F3pHGJ2IzqN1RhMKWKSMiTAFmvAdvY1dDpi7Ms
hoA0hNWNZuu1Qv819MDss3H8oeHzHuwpj5h3HGcIIwg2G7D/d3tse8TLgZ9Xd3po
eToactnHUAIx/BSGTpmiy2tvgCx+qAu0nNxe4L0a/2N9k8ZA0pp970shkRlK6A6O
H7LL5BlhNVmxYurMK4/iq7PM2HiosA8p70twDeMoXt/bWu1724nM+hcEW6iZ2Kye
McTZgVnj9MrZsxzOx/37pqatM8SYOf51UnDTFu1agBSJ9R42aCNxT8tCZq8cNX9A
qVY/+Z2OC37F/Pib+5pF95k2XLjt76e5iYeDxauSzZlyHRpBcIqeZvxV/Ph05I4X
tw+zZTEFDIouAaXmir0cX91LWg3hcUnCdxDDWyoIC2Nho8QlbhCeRlAPYOzEot+Z
4Rp5Hif/ZClZ+a6OwnDlRWTnsVmirzwnjS09a1WPJyQmeTZz4SPrCvDe0vEXrTzh
vYRRbyc7kIXdfCZtjqXjsaXY4YTowiEUPzim0Tv3op1nCegvRPSgLtCMFEAAhava
uoUdZLk+VbpZAhnLU3jBv1IT/7pm77/fHdzfuVMiFHv6WdAAY5URLBuPQYHF9DJE
4Gw22aBDLzsKl32ZJwdixfwtGLhh4Zz5UTKx5YqQfItVK59zFCVj07nRbdfpV2cp
Yx7d1ec3OLAnqmjUDhYwh0MdbhzqYhcVdU9hAczU3ze7JeQ2A3eLChvR6AspCp+4
GCHNXbcggpwZmaslCYm8pnZvqgzVC5Qmm6/p/j/3BP9EoGIdU3YamKdDqjYqak3w
+0C9FACOoWrFd3NW/wetR+bszWyYJr96Zuq8HhQ089OeICWvSpnj2TWhIw7rsXfR
wJFHxwSnTkILxwjMr4mHL642l584yxPKbeCh/BCozN43Q6MfLGfHXKlJJnLoe507
XuROMVzEgoTvdTwr+CxplsnpZFG1QfzrTGN71i2RPzeFcQ+xslQjX9c+YJ8LaXuL
1dqTv/4Pw4LQakBxrmGfygy9TkSE3RSTR49e99gUJ6IA5rJkcS7qZKZDD5O0OLr1
YV7LUSkaLlo+soJvuWcfjoMlaToo9u6dkHOA3DmKBJfQ80HlriP0T5w3zjG6TiKm
iBH8MecAZ6ROvdMSctS8yePXQ9Nqyo/uJujx5jSo6XiNyGpMI93NDEMy6SIykJOG
+ICHB+vdltkkpaaeGVLtswWyGWSxxKAQhKI+g7w9jErmbzrzu7AQnqSAuupIgbBw
UrWhPUBno1+cra0T33w16jqZZt5+RYIjh0ZP7a9qpgkQy8APfvVVVfIAsow+mjZm
S+xhLSMWVXsPrBiQiQizBuelOsCt8HrOcFbKx41XcFtdIrTtgUn1NoDlZoi707dZ
40WMhvr4wh3Mlufj6xps8wioHRt1LsLPF5QcQa/0+RUT257kIod7afSW5MLCgpyy
civiqdd22JA2JMtnbkuZM2ssGK5KsVe9GROITjghRkJCysy+rYRjsGovXvyJbqsu
MCxx+BCGb4vC4/h8iwyAobdgBUJQp9XfgxdOW++V4hs2yzBtBjXDaD6c3w6KEsXc
FcHAwkwQ7B0eK64zcWxPP63j9AZQEbpW5fv8h8dIRdq5WvIZ0RvNPRXfil/9ffZK
Ra5XyDZipgpEkUvUqaOjH1GwkUCunF0ffHjoNzgpvOw6n39kSMJHX18QOVoGFL+5
9JIsh46Ic8OA2oijKvR8KEK/fxUc0DP2910p122db9YM4o6rB5O7Pl+F84v/2hkd
Lcs2DBb6TIQ9lDMqny8rTklRqQ7dFl+1S2t1GW895jza+jwNuSbHaFzlKsQgA0S9
wBbUCrYMMkjNjk0T1F0CeYg79BVGOrjqheejzWRbHwUFyAAi9JCKd0p25IvppQW5
oxJ4JfK41Ah7ZtFN/v91s/xmuMRyR37QXpWX5ZyNlKDLU++4JK1ZC4QCS2XPZS5z
kfUBlgkb9QpyUMTun3ngaOU7WoGLwkj4IS1qNJAJCZ28nGq73WxqNTTzVY2YqeeD
HZ8Gi7lak3EswT7RQE3Hjsx3kQ4ZSwVXYmf7C4QsjFMvNnmTyFM8gvVBwhZqEpd0
X9P7Kzeekk9vDIOYQQZunfKIvw2CPwtS5nGW3AZGwiYFDHuUq+KCIKg9AQaIy75i
9cBeddys2gaNW/UoKP5ZBvOXWWgcz4DFeJM5+crxQ4K9WVfNfA6ry676Bcg+JY37
VnrvzBnV1Yjt8KjoD0dg2xTbaxYl25zaPE5rD/o6BDCVInbsuXPi8qmcg9nliWYk
1JDfQE9MP5PygqKHnzFAYGbVtk85SMe1hqp0cHio6VDwBaM4hl318fmdus+RpUip
cO9ckUnE38WHmjZOE/mkeOIQ3IIWbbEm3B/xm+DKKQnFpq/SUHN0AHIvr7FRChoS
ZNjj5N18F83OPLRYugRehvvdkozXyLmHxRphXLOpEMTocliNOzC/OVKcICZ/yc4u
Z7MZqwRbgaKXku0D1w6f8SDbaigkArkVbwIJ/nDSkJX8WEqf8Ix/+ZKO4lqXEEJx
Zh9V9wOCTmMjsCWKF/0jft1vb5clfj12RaD2bs3bsTbwkDyxF0rYNayCizV0xA7i
lxOqf5YSgVUTH+gkVczMY8RUgJGDtw6whkFXbcn7ciD/YCu8ynkXTykeN5hsfl+a
tRvN4RRQlOfUi1SyqOJ/BRaLC+KPVatp7wcN9oocAGVaNzHZkVG+WBTEFimjpjsj
hsk1Z9QMHE7cYKmmHywyCnUk2ztbWaDpf4BQovRpKCa8j/2UW6pdbD6zfXkihB5a
/3DF2GCD9T/09dCvrsCGGBzT9adl680HYQdafm0pQbQpjKHXkNvEKsjv33Mn8wdo
cuxH5vcPeFrCIUH8s93w1P8Yal3BuyK/PuE8Bk6avZMTpGGMp5CYv66ovyokoA3A
5xozC3bm7/T/HeuE/m8mNF21w/ch6G4/yVMxz8h/db1pYKoIGg8mhjtRLwifZuAZ
Dug9qh/om2QnwBFSZJ3IUnTAccN+KrDZHf1/L0Nlzr4s7FBVN6rhZxZhX+WeyYKr
f+lFsriYcfa3OCwO6En+HzZMgvRV+okQO3NOQKB5bzHkz6FYG6RVhc3SElemv24b
cMZS+tKl7aS8EXnnrUpbJAKsXrySawOEiEQNyk9vxzDf/iSvYIm3YuSIXwPCWMO4
WdZllL2aRHurqRp2EaAYWA2+nneneDlzIsvIpeL0GXFOWDsEZp5JQOAzoXdnTrfJ
SP6xLmlf3LjxV5eUle8iGOltEI2JybGCLZh4l/hSQqtvUEgD+uK+lD+3Ul/p1X+K
496PZ8bQ4YQy9UAsvyufvaYztqXQZywDH3sf8NVd8XsXUkWtvXusoScGiEFA0wmV
zEP0jO3TJ/Zp5W69I2dIZZCrQjeZb91om10Rrjk9Ho4DXGJx6blbYTyWZ3ksaef0
IRrSNcF+MGD37neUMPOQWy5gAnqJ9d56965CkhXQrOYn6ZPrG6/7OAuBYoozUHSp
GU7pSnM0tJ7d93olDoeOgCONf6aSI0f/KZaKA53RwAGzRfbdsXeWuoGrbCDYg4OJ
4V5HK7kqWOcYNa4g2lE/cZy+QBMRmPADVApV5ZLQ1PCDSS1UZ8DuCuriw0E7kEHI
nCtvv/kkGVqT800YyGJrr0fb2pQGnQTzaom6ugvYBcndHPU04REhoa/7yefP94fw
stNLJpUgaMppno3s1mU9/Q3bnhN4qiH2OScu7TBjYYYgFRF0nKdVy0afHUtA79Nv
RKzPcm5hm/Apuqpn2kOsKKuFDIxL9mrvi8bPe7k6229n2gJDoOWHWooQlx77svGI
1JxpWUhxvURaC4nAWGqv8wWvCMu9b67TJGM7Tg3wwjFVTJ3DN8AeYJYh8j6lhWCw
fL9nrA3lapx2FNHP8hpkLDYdicp2e8l8iUcBlCjrvXmIP8ZQ3CaJjPM2BuyWe2pt
Nq6pTF5X9MijbINrT/g+AaoldE4OqLMEzgO6Mvs/o9w+BiQzapVPlCJSgOTcWJEQ
ggE+pYjJRP+ir0mXw6rEoUn6fUlBJfXIMpuEi1uZr7BBkb2DgKOA+yzoaoKNkAgm
GlwThsedZrG4ywmmpmnikdDgwPss0dyCA9kwK6XVM0PsrQYK8zP+IpIyOrTiSknu
vxtaWqNRCpHei5wfbjtEK4IgzyiQhSMDniNGvQF/sTdBmnTYQ4pCTxV13qa9pp5x
yfyu6CdVf8Hw1GXp0cLF1wSaSbxxB1hNS3NDzfde+v/ExU7zsIpC7tuv6Mp82cq9
QZj9HGRgElGSNLqV9nrcedgG2C3tHOx0gJU4LActt3hHnUS/nQa1ABuxNAHt/lLb
B1N8jZSW+L+wm4xVrDkRSlR5tB3BE9A27VLZPbCLWUDfEBQO9bc4iXYNV2dKPlKB
Ha8zCLxiyx4EkZ/LOi0atWpUCaWOTMGm5XvrFSz4WlGbcSYXfyht+uy3+W5g6OUs
gBxyDrYCVW5P5dw6dEM3VtzJ2H9V0c10hDIVA+nYfUfRS/seuWLXv190PzteFlOC
klMTJCGvIJnxY2o7fAHy98Qb/vQtFm5y2/l973kAxtjCNAGuoR/8+KHMo+EFLuN+
sv4uFXlT397g6wylMdVwWuOW92+3ebiOfZCa85j7uScftujX6Y5qX+7SFTmmXSkh
hhaMncXjsvIJShCExCw2tBkowK/qIB84PyAtoIQ6zXkuaVMQwCeOLAULMsF6kt1I
EsfnBnKlh/SB5w1v3Q0nf4RoiJP+pJL/rh4F68AM5F4/2UeKAPUkoDT7eMHuhB9s
pgHGilDhWQ4y92MTpwitSLR9AH3OTmSMmsqd4i8mZBlIADZcWAUsKAW6WG5bwt92
j3yJ8DL7EjmOtoDyFYvAv1R5+z4oM6+qxqnPs4VX8U88hzNfPFrsaYXfnTEExXoD
KuZAJG+Cf/xK3pmmgS5fENEB8hrZ7KI1E31iegbMo3vmjTltoCqAu7NJVg2ihl3o
nBwTA3sBHhWzBTKTmISO88ziVoAMIANAq/6nM/v8ULlHD2iXohf+xQAaTAiDJTK3
xLeC5kLdUHkXNF5hmZKeq1/I4XYh/axF2skAIHH4QNpKX/9I8mwEsu7ZA/hLBPGu
o0MyEJrRwJtHXjP0w3u+yF2+++LaAdWMw0nFRTdyrAWmKOQ9t4n1vj5ud9rJfl9+
jKDZFNcEucitqjWByA7YHcfr0DKXFsmifX6OQoYY/8MSu53IQ4wCwIMCuzPKswSM
4CLPwxNdl6+wd7DHFlBAY+bQxtvm/bblqruu4J5nkAc/rJS1w6iWZEmBEuo2Uc/m
05lJClZq0JUuem63DsxmXjSlYpeGpG7ULRtMLG+b9Pa1S+XAZrpTCM5C2EOR6AfU
VT5bOrS3fw6y/OVMqa/Uip0rnf1bkgOTG6GK3XYNDzt+xhnayxsSeUQIfZC1kpRs
3Y296Fd6LGfGknwLCAjljCv0kEDLi3bB4W64mXSFKYH9SMi11b9xdSjoc8BU2RAF
h2liGeSPAl9y+JUfyRjHe02qCX0JjkFmnLDXF9zp1aBOK43WStar9Tm+iqhvvuP2
uvEXuJkzEB4L9yNLe3XpZmm+v6R3lXO761HA9q1UTH0hwV36oxoLhuoti7Iszfyi
Nj4I1GOzDb+944A+duY8DbmbacobTqnCi2/rs/Vvh+nEN6NhgIhdV35JOm8JRez+
zq/23ejSNRiKFvg3xAytgKxRSKbRSovycVSA6M62n3eIDW9Xe0ycDZpjyV1KhX77
9QOkx6MwcRU0VPHu9sEtdFROqhSi/i7RxOGdXOQk8Qu7w1gUVgTfvF0zj4NcKGU7
XzLH0/pZdNsP3L6jXso/7w0EPysK7GYmHqeKu8E3BJcZovwdB3hwYreynDQ+ywaU
wr+LYXSbbhfCQPTZTToFw9jwYAZv6o8CMCQ5btENu1pv9NHBSEI19Rvm6fJ9kpXZ
HUbE+tkQDeFHPFipI2G21WEDzaciM8rGgGbAsOUxuIMQQOgVOI8voOmSl824SRmx
N4OsNQrDIF32naze0LZlwuo3q6lcDHFYtwavrRQUaPXxOcsy9xf2gQuLDMP1nMvO
IeciIP+GJ8fFymBc2igJ6FxP2+VotwrHHbn1bRdu6UKpjXOpHpNVx49chBEBGiX+
+UAUU83osBK+307fgpXDjp1VZIJjgXQEeopfKVCzY53FGDiJ2t15/XoKNB467BKo
RiopraNuAlW4Fc9+o68Wg04VqataU+QWlxrXV/EOM5bKnph/+ncDmLiXttY3P/UF
MgMpIE4HhCBqKQaRcpCyIgdrtqnAAxXT3oTWGZiW73erMPGobbPcGg48L6eKZOY9
i2jC/JKrgTpzxGVqE2477ybe/0ybqdXuO9/Jr4SCE7/Tq9s3iFSQ1adkqitRlCqQ
G6cWXWzvysC0O/9raCChut52M5pTEpB+iqi65RH6WQlC9Lc5oLHyIYqL9XNUysBo
KhPuvNXOQrgNMbLXTcyGR8JC5N7xeaeUSNwxuPmSyzK+gHiWF5E3cTfZQXpeRw74
YDcjqBrjbCowkOGtp3LlpBRd1P3ggdmiQQUvHP9FfEK41/SGm6HmsoWKqZlXYgxk
B25iBtsljL0oO6KZqcCFtc5waqwdsLd7rKwDl/OyuJyE721eFWzf9rzlfjBTn+uG
jgozKFb1rXij0yKxeX7jhIQgx0FKhLZmZsdzqY8frzrrtGjmn+OnkrGzR3q2NeYG
+jOmQ1gottPGxxxlGnUmcR3M8a0G4d4ZQWeg0H5xHTQqKc5gdtZPmJ2Fg/gd2gv7
wrJ0oarXF+ZgZp82+1tGsHfooQTCAAAKpo3nwIDTToQFgEE0f+VDM59sv8KKc7Hl
rSR1UfYllhrVUwfzORPWszuupl1Y8+WM5qWX/mf8V/JCXJ2dhpdFseDPMZa6YH0P
OYCfH206wqDMtAD9ZF12mE0/nmto5WS7g23ZVbz2Co5GgZnmpZ8+p+p36vQxKI9g
ZhEQpeFWErGgiCs44SFxA4xFvPfDKOLNDQpHLIHnx1v2QgJQZtpEuBVIn93hp605
HQT7MUF0psae1olotKWM4lxNEGgogKiu7h53ypidD7WrmAqAaJrYHTQt2axPtHXi
RGgryeiS0mweo2Cx0MfXpGk/TOLR78mGCHWKqkOPHZfzG2bN211xYUrLfMUWfS8Z
Pxb62Bc71X6TGXWc6sKzu+9kaqxLz4PsCNAId8v/NaNjGvQ1UJmMpjjxiAJHFz6N
iVW4ws26VJy96pipaVzqhHWyWBgrLzi3ithJ5chkON/h1U1z59xAzmwqJ1kK2o4e
ftfX6Snr2csu4w5YbLhxKvqVOD5fIT9mt9anWWc88ymIfWmMkrQ0DnrwbyLzHhPF
0HbC7uJBUkJ6Vi42flu4lDGsB3YEdmjenbqQaYm18BnWmnsX9NZfVHMRay0Bo5et
Pm4sUTwP4eocma9EDuu2jCPNo9mxRsuLQMQadOyh2Zi2kb9wYqD6EQNxk5UHFtkD
BJnBgWWGxfE6xoSZ37XKydO3zd4qAutT6IiiLGzjGFD6v+eJuP1b9+ZgviW6vIjF
FcNMhbUgKjGMlffz/b7Wai51pXnZruYeiIo7bblZwPxWtB1+KzHWLHWwOlUH06hA
rUKGiq+7UnFSl3aMozZ8FaThzJLY+WUtZZzvwH5bsbiWoVxY5oQkJ+JgpXPZr71V
uU3FD39l7wjtDvlPC9uximMGh55V6sC29f84e4KW/FeQ+Sy2mh/0fmtbnfRRlXZE
dxUbULZ9TUmFTuPk8HrWSzAqG2sxZM13MAY+w8/sP4h4OyYkYOMDZvUna6v6HB35
w3gSvZAyn/tTQ5NVXz2rHQBqD5EFTY+NlPqWJGyKMbxIVPzgfF6i39/K1SXfZk+U
7M/DU73rBn/khLwehgdTSFebqbPnO4DXhFg5gajWWikU2fp0pqKKgGrdXygzxU77
Wes91qtP1+zo1za4SB6FZR+LoowxjBOUB/PNVPVOpoPyxCndxebfoeCMu4v8UTor
3ZJSuG5rL8s/9/XfG9ssXwg2Jwo5zMREZflKKTRGfV5wpMNpfXEGByok5+Dd/IWr
pDr9PQ+BiuhkyWQUOu4P4wLCv3NEuxUuWmf3LIK/fOkz9JD/yHteYX6AMKm93WO1
ZRdqn+sz2C6s7N6ppzk0M9i4uJnoWiJ2mlaEgR4F7kRBxCdrSzTSk41aRGI1VDz9
pqMIo5msTUtZ3VrvXGFxg5/So6RAF5YEw4CCj7m4caTaZK3dDIL4QljhyPpefhjc
DD57svcwbLUfNHdqWq80IZ89fq7kjfQrN4wTjMPTsf3XTwhnN0tA0URLTpafnNw4
LLe7C5DKy6QTUJMsz9HxfT5YcXyf+sFdf94nhSBi5EuInZYaFG8jaMg0vFx/taFX
tWSAnDCNzxRMrva35MFzj6QyB0Woz+gbUgIu0sbtkQ9hZ3Bu8/G9CgQ8lpElLALE
QKfQHHLZ3v2ZVji8uHI+Ui3bcG3uTfXmuMUT9cI7cMsIpZdbHWk8UVWflzHJrZXX
nRlZkCptcaRvaqdbwPeieqYQpXDtQ4SYuP2jFbM8cB4Ifb4ISFPYG/dEJiVPEY1S
s1Xx/8JCLsC/BhtbAZedloCzrFNGiEDmkvafZKTXZqznOWgjVvVQ+9r8B7TjHaP2
nO62l0XvcP6PSKamcYk4qllefx3+34FhkwtODPnwd3iP4ipVCXUk72AEyqVNONdV
yiDQIJ7b+cH6SXhVrYmEjiwRi2Bp8uje4VtnYWQouRmZD8TS4cdBnyIj28a6YNc+
AwsOFCvERy1u38uKDW1bc53GFnx5uDcz2oHBWt9DgSrr1yFqq3+Il5auadFb5tUq
gc/TBuZayd+Im4tYp6yxTf916pu6GING6dHPXGz6Z60e/RlN5W5DZXZFBOf9xbFu
7UqkUEi/OHQSfUUNwcCQM7A8fsaV1hGCHWoC0sU5MueToQskJpgKfSoGOTCfAQqF
h3E7m4U7V4n/1L7CYWDNZiKkpGT3yr6RUtR0e/ujO+4LsXPwica09FB8xXoW0kmg
+Z8Y9n6ne4zuQ2FBgp7B8TRwqaUI3JKwJz6+oRx/Io3nbudUMfKu/OROi07K0EH8
ifwLuiDrak/RAwwO4yNM3NQfNmQdMrZ8eHHGGXbydH/cmoaePcUsHwkxrWIPl0oU
YG5WKdi2YmIpzA1z6dZENO5arsDjJ5JOaGlk2hLnHRrW0fQbKwrwVijMU74PiDRr
EINMxLtoHaly074qFBeYHtqsSPF0Ig1iaKQyJn8vDcSu5UdYex4Pxb6lwDgDGlQy
+0HG9qNT6UlDHR9kHSm/W5OO5F1Mll9Hw7jCnnB7zxmx/WkC5SEpqcLH4Pk9rgVP
zZsF2zLxudqSTUoLdcDF/ej2M0+E7bQm3010d948kFfszY40GHWTd/85WVPBOZWj
GP5Pi70Zvc1lfuCxoRd45g8ZRwhdbnu6hn9e5eMi0FkCa4jD/aIrL8Cj6VvSLR2t
JrX/ZR2UFmPPTzczbhIvCa57alKTEApQrRPuV+5evVQV5vg57unaeyiHWskvUR92
PHgBdB8yqeEr2gA+Gp8TZ+BLAa2u3Oai8zL//C9omywx81ChYPSO1NnsuarSPrex
KtIj2CI5vKwzpP9mCyecdDsLKmJMxn+rWL23jZKuqT1Z3Sp70CnULdzEjcHf6vlO
uhCUqJ6UKj3RXfeua/zRebx2kkQalbyDGgV2N/kZVuwh8+lT4VL/mVNMeblOLGOY
1Lb340vxHUXPqTXiuraelSdSZ59W4rDjneY9z5bOWe+XQ/5mAmpDQKJO9t6yFdYu
I/luYgNVbxOyq0/7Q6yDG2mr4awbxNd03RDYa7u/cfqkhIEHBZ7FL/PF8G3/bHRx
68ElZhOpgoBQo8HPBvlzN+NIKxbO3FwRz3vfhW8J/mgkEwhk/0A1X7q8JYO6kPVX
HnoRsVUnhQEyiKFvZL5VMqDHAMg9GWYdxGndG1G9L/thXpCF/Rdr2JpBmEQZIYTk
CfmAGXX0VmJzPOnF/uGZWKiDPCw2P1fQYC8gAhMCAT3Hkm6Fq6mQTZPJf3TXwkXM
OIlxTdI/bSSKJWwJL5MRIE6OXkoz3BvC165N1Z815nHz66rZ1ilB2Cc5LWnUjVfD
BrPMq3MDCp7qFhgkl7iHCaiol2DEDKDk7jUKk7UpQqNoWaKWn5di8pQhXpTHgFU4
3hdg+t3jvTnbAtOBcChPmCC3IWcAQ0TSgtnp0JBJgYZtgKpaAM2w2PKMTgXXSOPx
hmdQgfj/j8pZT5G4FT4doT70kVE45fRK+gXM80Q65HtqHJmiXbAyFkBnupsKJiLb
ZXma38kzAsKRR6kcjFldGG8mSLvMC1fO32lHkgUxS2mtQd6XryuqWQhnYmstRVy9
BoNT86fhzEdmMQrI6wRCdu97Fjy7BNLn7obusyHwLrb1HxGkfM3V6trTZdiWqTnG
x79sAWPZPZi7Wp0fRV/HAiQiLutjSok216P0RaoBHYu01Zp9CwwmgGrVLYJNhFAm
4KuANfH6l/Nxk/ZtgHx0IlXBGUhKrrxkAl5QAkSLH9XB7UNd5RyGnTilVcPYjQ8v
dn32BN83yhLri6yqOTCNb4cvW060wWsAOmAU7GDuelTGA+dj5bWMQCG+VDqI5TdF
c1Imw9JC14Q6j+Yggv16+65Ncx67czItO+mD3C+AyGXszcoOcFygiwbcsB3JQb+k
YncAU1r+z3J6eo+o9fs6TFZXAFmVoa0ZtIEp2WtXIX3mTUBQncte2cUuy2HN2THv
U3NGN7nWGycP0mT6RwdlldusjvusT4AWLUavYHP9QU0ZMGr95rn11Hn/ybNC1FiD
okjlaaYjGrsb8yD9hd36IPTRfxA+9SCdG2znzBQcdYdL3D6N+SAJ0FI1eKRwYfKA
CT3m4WmCEEpwX40fxKWWyYEbfWlW0GvvTDxG3MpYnt4C0k/0sFiS8vcW9UgTXb2n
BUj4chFwiHgVqkNI16ONj263i3aX45twKnoa3l+uwJfkRPEX6AkD/reb4Qj3FQDu
/APHqNF44HIhKfjtE1hUyWkx0tdZCBWAPwcIlZcrNhYA+2Vo6Q6vFSGnmv6zEOO4
Y3CTnWaqcEza5XnRmN8pQoGgKEXRfi3dP2uezAPE6NhERI0gBfcUPx76M0lc5bPt
lZfjZI0eVDx+NhEwlBS/dyt32UmCnC4L/VgeBO7AdXavB89STHnH8VHkXxGup03m
L5HbFmBiiB/w+Q0LXsFs+oAi2wwGGDVt/fqa2QH5HqgjjkOOQQ9TuhijIv0g58Ts
kRFDnK+ffxe54i+ooG1Wso30XjZlPvnTYg7WYvaTdVxNBDHtiltHfFgO9dH97zyz
lojWWculbXoTkYfFjfRIl5HiqEMGRFxTQjDmsFS7ufEVQ+oeZWKTZV5tM2VfYvDC
srD8jw6DhyDvg8sgwyUFWP+7QpQQV+9UdsewReS38T2lN7RJrBqcBWc6jdzyvwuW
Cl9MKLuoyV3grzUzq4C8qTkLZzT7Mu+xeMeP+SNwzSUW+JAZF7st4HpCR+MAwwmD
AcHuRtMEeMrmJg7o15csaFUgY22YNAMnMrdhzInHhH17WcHXArMLHRVfGuwbh8Di
0Twh4lrFFHlhnINGb8xlOOrDV/nZlvx4Ng8K6ySvIfrKgrXNzqDeuL18Pt+iddNR
nxp3wmjDT09QwXgKw3I5Rsk+tNWpAWvy/eLxTSxKYcxjWk4P1v1faLwWYl3Nwfpl
ewI1aHG5pd5HALFVgUjcyFxeIW/loB3HG7AAlR2CqgQEOouev7np8PSPQLpsVllY
r4xJKIFhEeqI7r6XZAyzwgCN9GO8lCanGgUQpD3f8E+vM+2+rpGN+XIEuetXkx+U
66pEpo5eZe7mJ050ITGIYgOc3+uquBaWEeBZyjPqP7BKB7AxdSVmiq1/uUYAu5Af
y0DUqv3YYxTMik9eMV5cD9AhR5slGg1jxh08u8Shc6xC1iQqXEEj53ykmlSAoWqi
V3QOvi7a1a3lpbCfKV7L5vlI2QE3Rwqi2pRo7c628jZUJZkNAzJEyhtCuEckXliw
fTim1yc5XdrJ5LOiiHEzVDjMTpYMQnubv7u2MsDkCMKo6VN/yltPDBv/oJpvw7oq
BAPeaEGt1t5aLyrs+5CNSXeO09yW53SkmfzSorAkj28zuvEwvQX6S5KicHz9v5ii
4wsZQJ1ulHP/x6B0XZuJXGffkVOBxN4KATZUAYSj0kais+WF08saHWi9BM/FpUQ8
EQ+jrFRamXFXg1mvDl+c2lRAG+8gLP2kljXdT9ulqOwj+wwJ0XNG63prw9pADga7
sGK/jIH9heVkiltcxldiZQ8P52GOwPyPGNQ2aQJN1F+/oreVlUDKKiEjmNDJVvhJ
elwXuEbTCkajEXlnULvXVZanusZaAi92no+Se4UkfO9ZfHaB7mvH4tkxzvcvoi4P
yRDANOIuEbNQV4wYNrUUF5/0l5LN3HJEw5geQdDHrQfbu7d8nfDdE7ebjpDE+MrW
Qji5SPGZdF5nq3TXM1AaGFkpbzdO9v1Ui5dZorTZudPYv374xD5ewaHKE0ojw5iN
p+mrp4w0AJGKSvc3rBBKBXMOcu9A9VSXIBkDCsuNpBtD8K/AJCvRgLDUkFI9EE02
IJAoXBFgpJ8vMeWHOd+kbQBSLO9XYpKZzt+WSv07lRCVJL8ALxhahyTfCbQ/d07w
QnsUblO4y5+mJZ7EHR+HUQPbbNZmtYp5s8VvOXQpYCDRD7lkeG6R8en8rbBkVGbE
+mZjISTlE8DqATLSKQLa4qk+oZGz4sgsLJ79idJ4nu2lDbRZk3hmqmp7gBOK0uTt
Mrfs0ks/AzxOdu520GdasmUIUAao7aocFkN76oGA2LOEYpieRTzC78qkHSgAvnDY
OJfhZ/jQMEn8Bx88yUaeJNZu5bHUgk8/wES+B3bQpJhR0J1qytZtcLLV1wXMz+0o
WESsKITISN6XPm+LLhU2ufU5tZZgF9aLJXXGaD+JUyZEY9qbPdfybG8dV2ZpaSXO
/iS3XCEv/feh8lwA+wTpkqjDVMid+llvZQDepDuj1TUyz/xZtjzQA+/r+lKVNrys
+nwB6+nDTmKWvLMzpueCbS/6+znXwUfIsVfVRphXJuNJ4ehG3CkQhkYXqfo3oPn4
U9Owc2b5efrC9vtb24MXkXWHufPguBlzvEzQqjafaaK8ugOBrBisSOZU2AQymdYD
oPO42eZzLc3B7+2A41u8+JIh9C6sLPI9cs1cMsy1O7SXsQnbgrQWwM6DaOe0ZBWZ
xMt/RbJBw+5dMb1samjDyKfT0mQ2fyufpNYD4sdRKINiXWnV9hKeGmVj/uFZ+HWo
lx81NKjw8GuhSUFuA97OcY959meDHkSJNruojxpZlUiEZDYg4MJnExxIOY38G2IZ
olwGidopAwTH8QczAx5T3xq1CHoky1YX8VskfJ6ZXJTwf4g5v7izac993Vzh0C+/
Vn2LgvMceC9U9y91+Lf53RMkr1GbAlkwGOWBkt9IVsA3jbqxwqXGvgnc2iWBdnTp
HQYeypyHLf6P/yKFoMJC+MQzkeujmeEq1bX9xWAFaEBoQWDbkNxHIdfZmBwPepS2
qSZdA7ucP90v9MIWXTlD90bGfaivZ20dJDmKMNg3oZuTuUhqge2RVUyhxYde+6Bt
sDeVtuerhJbiceSegIC6D5gNvHRd4+TbBUVK8gF9e91GxQrqOJi+9aikBEx6QbT8
IKL4MWQMcvFkJpLO59UW9gDfz0cnT1htsAzjjZESOKwMkttFcIXL7HTEIH+Wuhvl
EWfwZRt6/FYpOKtLZh0nmWwv41OrzbRc93y9mQQ3800/zkQ6B00Eoenu+iHu0Kut
mcvqoanuo+Gh2inxjVzO0Lfsn7rXMHREUnP1xU8/Ww/xQLvhWcTwEEU5d0Na5wuJ
c7Rj71WFerdzFK+5k3CEx3tX4JEWyXvTzYRHGutE52YKUmEZLT7GJC3hOII0+2kH
IDz2UOyR4RIwWXuXPbwZp0gs05pc1i3dh2ITzGNQ1+hWtBcFbo9fHxt6DJAgURTG
i7RcLbRTHxduXxc0H0VJDV+msEsYcTVdaAOHhwIqHWtz4GLR4yOog4v4IV8CTARv
QHbr3gKYkzPX7nM8xQkZeRQgiMazk/NecuxoXIMkZevtf6zYpH1Wan5rwOVzRKWS
J8xww/ZsLxjGVaGPttTfQS8SRr6nbm17+ZvU7Xy1Lu835rY3i+Ky7zyK+AxeQ5J3
Lba80zqedZIaA1gd995/5dp4KKHCUJPbA2eBlLfpin0Rt3jMnjpJnWTUoRiRHhMu
I1XXwOKGNdUIB2P9g84uk5OFsSRaUfcMLShrGRR32qzy18ow+eLWxWuDK0rVCCHy
f5y8fKyad8ZMQh+RXY54UTTGyMlJKHjVrtN9uMaOFJKN6XMQLAcnuX31daF6zS62
1swZrxDBdi8DbaVNnrW8Pn4GaeaJgtILtWU1n8apkYFg+US6DzYYmaQnkoCkHLwg
3fZbl5wUSqsoIwJM1tcA5Lm8s+7WhHlPb69xjP9kkFzEvLx0pOkw/UmMZkDMtqEc
o32w7d6tjFicVLwBrjatdGnytaKApw+VKqCtcSNbYJqWB/BC5i5Y7leNAwvBsYXq
xyPDF8Sls5tekupUbUTh+D+xpaQGWK6N5pFbeTvmA4FVGuU/UmqtY7vo9RhniP8L
AXYMcmQfS5s6Za8luvvSU5OZYhk7z6/3B2uT44uYRzGMN1M2hWuUW8rnmIyU8Ozy
DHHY382bLip8uHjWNlAxDf+2ET3dztLkU5QqRKElcA2aFcQvRQbfdg9phvSh896a
9vvbSFUFXsasPqbcYbOQQQSK62T4uE01pfISpi79gmeT09rRTcTM8cqAXQj+EhMW
AsKfNoC8WIy+58aULGkz4HS9quFtVckGvcm4QvuTAohJUf2/OU5brFfW511rCqZi
wC+EAH4RI6OU/zF81iNm0P0ZXfZEA4KEMJZ+beYVFE4xRzCpZxrZZ/0Btlz/d1s8
j9DiYn/+7GiclIs7CtjquAvIj+bJm4C6eyi0L+zmw6n9DrRS/MFhMChh97TWUl7/
mJV0ZDJC8SEBlUly7anaY6VKB5O4IdS5RAyIqYk2fOIfRq6ooCmB+c08EjE8SDvM
AIqeYYFdPbkD8xO7PMG7tzY8f58Cf6GwB+3xFupzSUScBQF0qrrxz+1rkPmnYXuW
7/7KhrudYdMvskEFmKClVU7+2GhNW12mBELJGDkNLHCMw3AC3g5cLcF3oZa5l7oj
Ptuag3kajd3n/sAbNyzMWWdlUWKi9RWYzy+UMVW0K4xVk1blX5gHERVQ4Yf41g3K
7o1mukmR5RdZPkjXO8skc1I4Wp3N3zNZ08hLPLYF+hx5pGm+FSekpIy8t4s3l2IV
aXUokpqD/MJhqN4x9TSp5qc7jVD1gMxng9BewvxZ3J8/cYqYrTkeJpXxMzs9bEv2
HjsW5gTmNKlPhnj6uM6oJDyH/E/IMqhO1YTk+w+3GHkzBRxVZkeAb3GpJZp5ICyT
Liu4henYIB7f6pdszagatZIFOCZr7PIFYOLf5TgcRf7Si/8Cb7d2wObzf6aV/v5m
4acjGaME+Wpyvh/XNCFrv5HqAnofErVax3dQ3ZxDi1AAYTznZMGvf4TagQdMg1Om
gWXG3EAnKOAS/LoKkiNrCckxKMehJXLp8TIiYQOkMRUrQjA4a219hD5kDdaFyvLe
KmYRru3DW6ivz0qIwmotSMUiTn36scWJaLPvTFGxwDjUkGnwREwR0VcbqWomE3CF
2isABkpp4cyZ5iwxrl059IatLPz7pIM60d28I4NHwo+qqK1ftXwtlA3qOMHOJ0DV
rsHmHs7IaJ5v8LFL5k5t5dcbe9KSfizK3nOEw3C7RryvmKuxZKVfmQiG1ONhM9k9
5IDprC6eZXeNGaHMFJqMHdmP9HQ2jzaxNbnDTorsyDs/RBXFlX+p4atoYl0ztwGz
KspN7VxchKOtBaKwL8L+I1SZ3vE7CruxGEfF2T7jHIF3pvydSjltBkitsj/z0iU4
s0uN3DWl9ruGFyrlYSqo5wu+6zkUaQROrLJQdWiQE2U0JT80wUUiH5GrMfDlhOaI
339jhSKkLX/cjU9VY1ye4hNogOGaF6/k8yt8mPIZoCJq0ej0D+65JsfXToFFiVl3
YKsRd+UcN7zZx4FjqMLtIDskUaAHXC1nfpmqxCrtcp77nG33J8NPBn/vyVrN57Mh
V25ykKq/IXnqDgHz5TIJrwd5VrScHPs+ZxAREQnsTTWVSLiyWfK5JXVsl2mLB5Cm
+Rw7M4QtPiB5Z1HTMiT5Zmnksv3uhehk6FURXNTfnVIj38RfcM4ad9BArxfxZDQA
tG79RMB8eTvtSrcxsc9eDZ+BjWoKSk14BohL9ssYGt342perX0fV9V8V5byCkxma
Z7Xcy5CH52SBzbsRInIQmmCiBs/kBJEIJGmW+qLacjQBADheFy0hx8t5FIP1ewzb
w3iLkuKH7ZCokGFUphYF1WmEV+pWTJtzDf23V4X/qDeOL6S5eTVsv/Z8cuTd0P2/
li3cCLWowu0ObdSPX4qBWbadQ+l2G0GrQDNhg9PxpJUqJDPMSeperiYu/9jXXedp
zABrO9s8B5IIjYrtAyJwhiU5E32QgxCByq15ptPbJLtLZYY96zqHkJRc2A9+iyqN
B2JL3WLAVKL2PBKXTJE1eW6n2ofzHvXFBBvtk4G17r6aBF6B6dTCcBqiqNcMqs/c
ZTeaHGI618iHIjvsrT4CCGHobetpyDbl6BXnAlA+5RqJaleoB4612FLi4Ld7ezFh
dHO8rlV+k72xHsSPCYDKm1GXdz94+wYAlejOMw6uRjMh5v9lAC5LaTFtZQ/ls4r5
p97koaqg9tmo4WHwHnePqVNJ00A21oNvN+0V3jsUklvUWO1qGYFiDm39KGor0Nnx
y0rWpNVgIEvCLVtVzFPvnbSRqI+1RZ5Q837c3LI21B6ugYoLsF9KAmRv+mSnw+jt
Goh7qar/7qFb+PHCTwX+8loTJ0uUoXiDe1LKqg/CwKj2pWmrNQvrPQBM2djZbgls
E62Lz+otmdujQmoOm9u4s0f81b+xkzLCONCl4GQp+4OF/4/y5cMhkBl+pTA1n6tR
NY0zvh9Vd2EaSm2P0pFdlTszGFcUSGgtiQh6YSBQ1YIyGdG/U75Hj/NgcXfcX6BK
zw0hGqd/l/NxWraCi4b8qMSGK/QA4oK5cSFLfS7Pm2Zud43v4vH2YYotqNRUMD1+
rKvC4b4gMh4qRrdzH+JjUeKv2wNSYQCS14uyjroWSOdLfcZaiWazsXtCj5mlzSla
Thk+G9czV6O43NtJNGskjG1tKJPSUIOdZQEiAZWYdOlP5Fybc2Uc1nODJZyCTsN1
uUk7eophFStJaDTqEkr+wT/858CbjQ95SuW4zKEfid6uSfwfpDZ1/z8PcRHuFpM0
GyropZTmHsZipa/mkb3JyyZ3t9W1I5MVN0iT2XWcN2S+l+5m+GIYf/gq5tqsP7jy
GA597MuiP6ONMjMROWHWgXsHB5v7d54lXppVqbunzUHOlPKXsIBfsA4O7JdhVvGH
oe2+oI8HY09+oO4AY8ZPBwJairdkxNTyeUfEQzdVMMSvRdT/tu6r0OGF7coANvLM
WXUQDWrRyTJD8m79WTvXT9P650lKNDZChXpmvqDIgB+8bKXR2iV3jdgebo15WlmX
F5YJp+rqSGbLMIQToJAPl8TWxpZjxZldxCc5wZNPEk1OeRgZWfkM/Kyprg+f/yyG
lADl3Q39/VOHETtsbpPbuZ6yTrdz0izHuLEiM7pgoFWB0+4kQXJ0UpwaT3TDGdxj
j7L6FhVt7/YD91PC4fka6XFPqgtyruTX/g1J95a7sMVLSglKowM5ow3tsnzMHgWZ
IGcB0BhVs7MDfY+KQz24m1vLnSsJxv6vJSv0QMdqzHkKAubcFCQ6kthzjxo+NYEY
1Di0JW6/hdNr8o1N96XcJGrRCc/HUyUuRuft65ZFvAJq8szsJBQ/yHaIzUyhIu1F
6fcAOIe5OcqWr8JRRUvG+eim7v8oJfT0XtsfvYgRmTNkx19OtixhMROhDQZDaobq
D6WZPUB4Y4cCO2+YsV+7rYBd0FMUwBt/QCSOhWRrT99T9QBGE/O5tDJwsDa/74f5
9jhW252Xmz1cbli0BA4NZ6dc641jIrSg2djruRSSwKZsW4/FAOeC6xMeg9FQ37YH
2ZTSBc0sLCsDoyxmpymTOOOq15QSu+SfXW2m1aTT1aTGU5c4X6cHdIjByB4Qevsw
NGwfP4b6j6cpU7Bou7aOd0/AhwzAS7NJ+nOAp5g7pxMJZvVWbqVtrYkx0RYSosVS
6W5IC+XOL/c7yAh4LKojDbbrdG6/Zw/xHi0UeKPs+hsIIxy/RCAxXEexV+EKOEP/
hWmqLip565hO5C0R06cFvbZDzSya9X4ZXf/zP5WYZs3FTJ8zuyYoojIOCGUoct/Y
n4KgOCyENXKeaDboz3CCXIdJXY+OZWlEJlIlMV9XzH5r2xB+6kHfeyFtrvOLWdZZ
JRYd9mMwqKI4dRt69XpxqoiqXqPuWFFF3MNY0oCDrYWiiRWktWLPGtEyXd/LbWX1
I7IN8AZyMKfkbeE1Vqdr2xb9udk1GwydJ2AcX/MfH1qNhQa3eW+MHWxFeue7X8pn
8qZvEhyBeQjxszyQXIfn+lf+1ILbpE1wkVEz08myjO4z777IDejAa3jvvsXIJCGL
SN++0vP5jDybJJkxTee2eY0URfm2QG45Tnnb/Q4ZkjHLz8vy4rH0MRrqsFrGIiA2
bwVrUQmh3o4bApbM7bQ4ZQe9LLzJZxP8o2iYZVS9J1tcCUZO3ie09PlBDGiU+2wL
FezhKhbzmZ6e5RKgt2GTqicVteWJzprcoDg9u5dxxAo2L+KiloFRKLzsizxwBGSW
cxtqZOyKtfPJaHbccVtWbCrDvZEOpOC1mPcRNJA3bw9EozV4No0KT6vKvN3BPHCN
gCYrjCbfSyrWnCrM28GjVVqOhxBdGdcGVTzbL3nhnMRPHa5OLWrjVh3UYheKQbyH
SVyqKYrfURaFBbZsIYPJ9S0YTYuTEMJMTeAsH6GnRDR/P5oU5lW/OMVP3TLng5lm
/EOH6+rpxjuizx5LQYBWCvFVe294EUcGzfCujIVTuQW3SCgw+nENnVwHRtkIAsGU
PuHkiXD8pgazFkUIocIEPPvLnP65DdpZkQaY96eHOPxBYgFM72VJzO50WgfLKdIj
YIaiyrBDFF2DhPDbP1AZfBngqELhcXm9tkO5Ibg4T7ONSLx3wDgmu6USazxzyKFv
Thxgr905hQ9oW5DWDAGEjud/5GQt5RlI1KJ7c8YO1Z7ehwGM6eM79t99ua6BISVy
2BuZQz6usXmz+2IdffPFe1UClkfdvfTW8VQbHvI7CbfFo1B8/WjLUoOHadwG5EbW
7EOGzVZOJouhej5dH74lZa/ap1FSGNfBLTOuwYLR8una2cwl6pJHTo0Qq/tiMYvQ
3R+0JY+aEe0edNEFmd9dy4ocWK6+TKOR2o0ezugwPQUFxvQabUFlKKijUK5/ZIPw
Rew1TPkFonX0mgc55fjSD585kWp8xnWb43VIP2qoPDjh0XNW2lrRreAdByziZDjR
bDJXv2V3VVoRBU7o/F7LN+2WOw6LZJ/aJw0ebXT+0Pysh+gQsAjYZZC8nAGkz54D
pv5W7jG/sWjigjjobPVbG86pV3aKURlQ1M3NyR7JRMSbcnpNgplLNn6IdAjzoYja
5wYNNFS1K6VlM6vEXlgp2/9xPOeGKmdJq4fVDiSzXjgxjy0qCJhkitGlt9UpcTSj
IeRaEe1KBgU0hgM+zWah0YpCVJNCJY5SjHvro4lcZ2M4hSI1LFCM7H9BGXdxUoav
Ye66hOM9MrPIl677vzCh1iQ+iLEh52lHEifdNkYmw2sMORhCXVJr2NZCygXc2UOj
cJvNPW1Rng4e2sRMUdCp9oORzX+WLogcbqZ51ZCI/fPFk9wzPm8qSpBii/9KojeV
2dRM05VzWlEA9rUjsn5HHnqSb93sBoYfZgI77mZkIjZXauksjoUgBu4e/q9o/L/g
q3BeyCSbQwmdyI6M6jNI6NK5dziKM+RnAXuzfo+I17VGJHG0HAapFG0TiLD3Je8d
LsxROACLDPDJRQo3XSOMo/adnDuROhmGv6A+ixr+5vG/a7aeA6tI85xcWMTvE/1X
ByoPewa62flKcfRyAHAwSlV13IOyoGhsbtDPZCf7L1oplZS4uBOt2qGhdnwsoI4x
7Fmpajl4cO9V9KzkC9svTyLxGdn/LySCT8RUL9Jh4JJdzCIgcBPU4iOKsEIZM2y/
a2IzEmB9Ep2w2Is9SIz2Pa3FgiGkcpIk7uri8cr8H9w4/BQ0JdUaUdzn/10x2dR9
O8mtS3CVR4ja/py0nYk2q5MsLY2VOTWowSz6jOhczS+jbPQAI65QrukbU+6GA+Iw
nPyxY6ICbI5hgKVPeADWms8CURU/vKQFKyknMUIo6tMq2lnlhNCNmgRULthUby1e
PCo3EASNRcMixrxNHI+E1daDacm0w0bcTAqWfM8HPImvDdprEcGGFD1eLcj7kBig
aC1Dnr/6GkESSuyryC1Llqkx1rvMr+lmwdwbM0568761PXllTvEdq83zi5/q/iW6
w+h1vrUSO62E+5ckznB5TL8Uqb5nTPsVqHbo0UG0S0lcfzn2t1f+rWuLUBWl20+u
UPr9J/qtL4sKXnkBE8DjjAQXgQiiSeTs1TakPvts+HLWL8+r7oYirhamgYAcMd1+
cuvF2rVlQyYCCCWP9xj0lLf4doO362fwx3jXfL2/Fhj+ucq9rjbS4ixGrln25g1Z
af19RuwZPmTy/uphqhwCOZxryTxMi76t63YvO3IWOI/rS9VLKHjbcjnl+3oE4du1
f51g/om/ff67fJJEb+7aXBpfvElyTFk9POD25PkkGUj2pzWfm4Wd1YZyiPPiVP3Q
qEt23DpV5/erNVlY7o3GeGG3R0aS1OmLSYlmotAro0vL/wa3LP+PRIWxXCSSKijU
YsVK7hO+dSWn+qmec+gIAtppyo/flQ+Y60oMh+xZxZ8BR23/eyCjp3sBsqM7M4T4
VDN05Syhz6pjcVZOZrasHNQaLEdQmo4uNn4qt7Cbe116TR+3eoskxKa/vuGAEE3k
wjmh2ZK+JiMsKQycCDZ+UdyPWZZntnNz0fjaRe5tieWTEDywvGZ66ZBmKEwIHrhF
ZOZxtTHt5hR0+P3jKGLfPguJlHi51iSmX+tRq5zgbE5QcVL2cPmfRJuw4W/l2Q15
+1gDsdYh2hqJgPbCmqNPw/QT/PxpV5xKbcEDsE2XJCVtpcj7Fwc0SyeTX42Fy+GS
QdSG+SggJ+l6rFhOijGTcCuImfn8upDSLmbDo7MzDvvwTqvDo9Z+p/aoGMFVYj3V
H8OOkS5KnfAoWfGtxxA3Y4MPlPHanGSuBiebvlgxqi4fcb2y/VuetHwSSTLvl3g+
LcvVVcu9Mdis7xZbmf3Omill1LXh2OcZbcRWMgKKiNI2iZvzIHLs6QKAzMBFRZsN
yubO/1HzRbVCaUBxC8gfItQ7NLk4C/J2Cty9rtVHxAFpeePakCwZQDpNS6xxcJS+
66Y5RiUahUyr9EcFFWPtevZgpfsvTQwpk4ndviPQlcCcZyD6kJOm16Z8bWd1DthW
y+22nk/CX5tXYoaZxpR2sqEILx6bu558aE6F9HUQaMGKC4FxFrYReI5BAQTl82+3
t4cPHlNInaXw+QOtXiDH3L/kj7L2W0fqfnRnQlVg/mVZKZLD62jLvJN9ycT1Wp6p
YelxeKGFKBgxx7A77KX3l+p3gGJrcSUde/2YldFNQeskxreMM9XYVCANHwOj5a3A
9Rie+xh1bP3TW8U0L6T253Azt4P1OGnz/El/Me5QQL4tCG6o3SQ8lUnTwt1OcK5d
Ju+Imn1UPl81LcqdoqXPo5/38x+hJoc1JsHJbJrArAATfweyeSFLjBUshZneYgJL
Dk/BgriwXssM4o+K4f/38TAjxwQm9rchJ2UoBGCbnzZO0Hh8jp6AeFB7A40Rr/HC
Q6hnCg1NdISxm19mXw2w6aW61XtyaGqWvlRmfPHpeVPuAlqNshWypOC9gkUKmRlc
UleuTae1K3CuSAXTNa76scRx+QJe8wG1LEw/IMMinfiysk0AgDT9Rgz+kskevEZi
4bcrC9qfgzDyFibcRey0Myp+VLa1sdac6zc+i7bpZdneqKUcKJZ0d5kJb/oQUrj7
N6kMmksS3mSj0fuiZJ+a048OFb0Zcn0Xq4k6tTH3c+OKGjAuwXO2f3LWZ5EVw8Fm
6KnDNZAcWrHq9QzlC+M7QvVgWxb/9XsaBxMX9n1yIQ3tzG2EEj8FzadFmSBuMsq0
j5opvpjBJuvod8kjz17iNOjjBCxkmHbEhgJ6QIDQw5ImoLrIzJrFGKDTDLzvWuDL
dNtZuxNK+RKync8osuYUbK3l+WHvzSdcdc1n1ceypIGHsMkJAaFOAkilu4Sw+e1H
fLvcGRcJj+D+ywsUjC3xVcSnJPb+Fmt5Hnyz82IkF24UjcrWXqQcvdLx7BSs0i49
7c8PfKalhLkyqO4yWwuiveoEP+T8HmoT293TcI4WBjKSlaw6XKx3qorkAUW5N14o
4jzEenhRyAzHkriWeRC3mL4dH/Jtxx7tr+jZ/SoKBoQ6I+wsndMSVHtJvVuvAggq
UIcDNpQDPgnrxwyMPIwL2vvn1Yn5bMugu4haAuEL0qs/yNQIDkCqLnHDTy5ofZhz
CkhmAiiZThjFE4cWPjgxQWe8weDtagESbNB13ixsRWbcSGQMm4RYSumRKjriPpJF
EijpYUgYCj3zm2/+a1uRUkb5BzJkV3FOYXzmsfI3nxVH3xs1M4gqASo+DWxXv/jF
3RYage5saE79vTmh+fDCXuNThEB+oRgsJa56Rkg6cJJ86luEX96UJyIdEyEiGF5h
Bne1zNcNFbZarBGwaCJrF3GIQzHCUW63eQLWE476y5QyK37IvTaMJ/R7wBw47uRQ
0l0Wr4rVt/u+z7huxuqS6UOnpBMN/psdmha6NDGXibh9y/5TP+3ZP087uee1NrGB
UEaIpj8nXHakryMpM5A0TF8UEx455L5rJkkrzcU5qEA3ldPqh1W1nuvH9p35EefL
ZvkoFPIyA+y7CC86F0IVyqaD7qimDBMUCrTQvDFHH1Wqyh3MRaHGbi51Q3skRb7f
VxCcdvEtLN9vbpvUe/WCf5zHLpLKOmUZp4VL+9k8+Pi5fBCsC0qWMwmglLZ41zrm
4430OXcb5NBb8SmPoM4QRXDT1kkeWX66lHdY6IuuGj2Q6GZP71HjRjvF9gXn3qh1
zdKqZBwjd6s9IxEylBO7gdRZ3zEL11YChiNqYqX9HcUziZcezF9EP5hUKVmIeZU7
KgYzubVTMzgBct3mXN6MnBSC0qIvJmmMksxVCrahmC/hFZW9eorlGjdrOm1JVR64
rIgqKECAW0F+Yx6k+qv30043IsIHAhkrfKnfVr/dn6La/U5fRl/+EbtdUKQIhiIZ
R+/LXjU0QZJ0qR9TpupRfEY1UCB/wn9L2htykVL1uEPiMRs8XfeqUkcMEGZBi3Sk
zIIdDqwiVsgQPyyPd2fAA4COz8rez7k34xnre4BcjhweJYKrQpmAskCTvNHct4yI
abXMLePFsXn8l4noyMFvHAy8+CBZg+AdSCQHdzw0QSOfo+WLuMJ20Fai3iX3Ipi+
Es7ULeoTZBDVW04eeZuT3E1yS/Dn0VXA8ejXR0rZm0lFMOCgjtFrJTwyCz3eZQGh
ao/LiQC/D4mLrt1Ap+yhP9fNxfQTqt7YpJg/0pNzzEH+quXAt9TBJbOlXKSZUmwt
InYhcBJrchy+o6Ei+6bO4PDuxtx2CNmCJDr1nWQ5JZUFvIxTCHgSNpd6rXGy/NKo
HT43qiW2CqGgQZ37Z7sKv4NFJRpp0kyu5uSe3Kt/Jz+KhtI03kBtGsmYCfG/Jk/Q
Y+LFbMw+rVq8okReQzUzcCRtsxyz+5HlIbnnh48UKVHySShCMxbEmU/hm8jE6hJT
F1u3CXdtgZvCUEDn7I4jCLsk0zO74jyCuOjPLCLK0xdaAPFOtye1Zi7kQdpAHiQU
imEqBf54i568zg0iDKJCH27Ok8Vry1ql6kWvRXkr/t4l8twK20fbcWQMoNHLITsG
EFYU1IUk3FiD0M8cASyuDdzORMhLBbkea4+0BRB9C0jvUsci1vJMxh7X3wWhs9UT
0KNpnhw7SWBbkThYfPHEauu4kINeeGhWFuGtXjB6WIpBGUvGV+NPurJzZdpHiU8m
DBpYUlrlQTgrQGlxh9yO2uhXWZFxqV3u91Czy4poWCk3NOKtAeyomDV2sUvYR/qG
xzmRP4mVDRinGizQ1JOppcYKoRnHVvnTfy+Ldf7fD7Xgxnzs66updkO9/tLS8DGz
HlP3AK9AKyv2iCw6EXHYr8vQYvnYCWxNg0PAcw7l0PvaB7g1C9bIuwXbz6Oq9cF8
1a+W/j6u9huPzonb4/RSESO7WwA9/gzbBAc3xvRoO46VUCd29zgGQlaGKuTLvccp
zwKkF9CWJbQ9MkfzdAu2PNMgJTpJF8FcbGG8dJml9aUwgHoDhdZ2VEE+NXOWJOrh
d1job3dQnVl7xnjeUEB6zKn9tehPzcDz98N2arbRbvsJLTHgBZ8r2PTk3RYZtrbs
qqvtk04NHcaSVweTSN1mFlkmaN0hYKgGPjxYpk2OERzKqzKFoBXXukjhrHCZNw54
XtholojgieV+h39YN3OuWonwyTlTOUJC+eV2Q162oU3dSSQE/RMPJ81WnfacJIyr
6d5lnviOIls6FPC2mXT3z6pzfed+IOkVRysQeuBwRzwLHr/rZzhrePy0fEBWo8Op
yrMmwYlMevGZ+9otX1o16h2cYjZyjf2jiSGmdeaUNkM9L6leCm7+oz41sZIpVDWy
2PWVgKQhS33pTMXiXB0pYH2cLr7DHWILD08unt2N5GHAu70VJ8sijaW6yBYe70XR
Q/tfXeSQtQ+T5NUcBD0fs0YF0S4iVlsdcw7936yqtJNWv4MwSH1ulUpV+F5p1bIj
hR61ubdTg5QwYlEGY4Bgp2x0RiQquR0r530D3Vx+Nw6bc+bBI78yx917ALJdN3/s
wQoz0xQxySxZiqTRn17PiP8cyzhRWkcwRqHEnUxJSsUNGLrG/MNLIYi/3CIxi8M8
ajEOEkJVnivDPnbpCwHjOwO2+ozYJE9Sr4aedcJTUwrv7CXUauitx8UYdds2mDg8
YuM3ImW7v9xCdksLEniytIGjKgxOUE7M/0IoXkibGWHDQhddWjYgY08PGCO2q271
CCEiX4Qq+dBTqe0HVAsfxFoZLx+mKcCUSK89iD8Ezef74VEbWceU562o+66HYogS
XLreTxEwcZg8eOkAmK/gcurHp0PZ8SbtslOQ9fbS4FoLoQfVpLHDVe838Ll8A2mu
ae4vxggWbgxog64s8bD7vR/1LkzCkr0UbBEwpBJADZfJK4HGPUQeRCTgb/Nfqe0c
1xWnU0VQpQ894G2u03T6rUIRA+TC2y+RoXbco00setLNlhIsM8H1xZqU+kwOu7+6
Eexmvx278zt2zI7UstVRJEf/Q7h3SMHmjCQlPZoxSrDpm9k7AtYw25P1dIuovht0
VcP+8Tzmgx0dXyArDYSF2CxmTsNApnWZZpj8TwEaz76XtjkecXwpgPqel3l66+BI
g/EgzfJWqnmE4VWvbVCnxUHoVsIvhnFK21ikw3gjFR2i54ltHv/0xd4PTw5/uzLy
SEETh/dapEwK4oSnfKRgA8ZJTBNnV1iqWW/ELR8K6JUWfQaBjug/2enNwFqRY7cc
XZdLN/eoV44W/RfH4W+iIjUKtT7QBCPXLZVSzF9Sy8zfp8lr30nSNE7yQsrfzHFH
xwlNZzwN8xZPR2enkqE+9RzLU21PxoRlUPt0l8qzh/+OpbrIcF8wjLUfpdS9ET9o
N8tLQ7Jxai4de1uICSacaLP22IaQrQa1PbSrpQ4rKRy6nzmPWcerZnzYl1GH4RLW
LQ/AL8eV55JfmM59Jc3VHfjEGPBmHiMMf+aAGuYOoA4UKBDkSn67elDsfEKIRxfS
n7UQSVXHHOggyEhKkBiua1GY3kRSnvIRaFg8y/bfr8n6dPVpbr9h0Mkcy3ScHr9r
W4vi0UUaihyFasQx5ItO8GlCAqIMH2/k7HabmX8rjFDWYvHqF8tWTXd4PDQkKHWk
fI0pbVkulhds7DhZQwyKmAte7n/ocgsV0TbwW2JMDAUi0vnyHcxxbbZ53+ZP9zwy
ljbhgZSPau1d9Cc8TlQeeS6k80juiua0vTOfdoIg+Sum4dvhhEzIYhutYaCF6MjR
BD8+/lN35bpPPpdiXolirzLhih9nT2ThmTSQluM/D4kfew5Zz59lV42zBu8yo5rH
bS4P2Ok0cltKgu4JOs0mgi71W3X+2eWxVcm+lBL6egvs4CI/ZOFFvyVgQSO3CRGA
ywI/ATAKmgQq/4o3VmV66Wx14yamshhYL30jcDYjNzNdPPSQXxEq64vfkuHupGqb
wCnHw7752+gstsmAUCVUhcV10w7xPi6HmqVUHZTJnpSrZUzwfcujDoLnSBaKH+bx
FybUqHEs75tdPmhFCMzqWPYFOEGQTI5/F7hVLfUPeFpoocC4tGwe9RTPtTWjSnY2
7nEfFLNO6cr1lVkjw23lKlXtoyTwWrE5wQ2NgDuiC3urwnVKME7puGmkxpBPT4Hx
iCsyqMwtf2Fn/L/A+8JsBGHtnTKF1ZcqD0qBAPHFSetSyHBiOuJRpaD7jV8O+0jn
kNcTTo36FrMDuBOLys8JoDD4YP91N8snNnBRd4lxb28UbuHaZ5Xc5dJRO7WMjH0Q
9BlGHXxACyYRhCm3YriSddGrXwe/te03WBD3eIvPZeBXTNYgUewq/RU1dVsX6H61
54HyT796iVR4j+kwRg/U2r48VkGa1eKHQy7LqXVB6Ja+ODybze4vMVCMWdOTn3Sn
x/0IL95B2ocSkSQugnZphvkaRDYF/YPaw4+rXv2v+vEeUKyCHOJMipfoSJkVsixP
XQV9LKN8YiwPQxx2ooBI645UWKR3TiBOhWRykmBx8ISE2AKm3xkqzYvmYpiqJHl1
h9ruD4toI3S4bLfzSx0rP0dB2HAMWB1LNTHAegGmmWaJjNBcu+tpNwqEryJH48p6
Cj7VpHQ/H0uCR7M74DOd0TwLl2L+3A0Zp0nO7SP5wjqNg8AsXIyFpAhRFGPuAVY0
Os8sY/BET3CA62gPiwXXwiNAd1LCLQgh00lYuic45sbqxafrf0r5I+k8CVEvMqO+
MIZAQ/u/lZoYRXe7K6mOMZACO+RoR4eZ8lxm/mSEnAwYRjI9p+VQEFYmg73af5Fe
0Nw8AOt+s7Y2cBPlju+Qa35VZmm/Sm6xMwxlqXPVR7x2cCdGF2ftAF2VfazB5PQP
v8AUNXF2DlHudP9js2fxfcFkaLKTkxhk2f9wDInNzBJRyGRqa/l0b9LR8qw+OWwL
5ofv2qnwzfiFFw27c4fKEboixCZsH3W05Luq5CBlT5VEsM8OMAyuuVBL/65fwVF3
1ykp0+KCWtN9R5xzRQhXnmaGVN/VRbzIzhXlCMnFowoh8J/xnwLpixhbtiBYNpK9
nUpN1S0/m8xQo2PtAuBznvGggveNvxCIpRu93A/F+claSeZsargg6tzdDc7OrdQ2
6LIR5GU4yeUNV6pnbVKHqdNejOPkwjMswFpEWCxOAyD+bEpCglTET/Qc5/zRNRMs
nVcN2r3RZvc5a6qfvb+8TE0km/MBT/Be/HUmvRo6JoNBAPJeE9pb114qtjROsk+w
b6lSupJaGOvYvN0u3OIWJYbfwQv/jxaVWvyRDm9QqIA/FM26l7meXpUn7XECLqpk
azqO22qtKXIBangxviFfLU39murxtyAjsBcJcZV6+KJL39cDJl1ejqOUQPjuSJhR
feNW10Lf0yAUOHuMEFNu2fd6k1n/ATO43KfEVl/Btf6qyvH/+T8srVI0GjOyugtW
yjaPP3saOSubxSjQI9ZrQKruBt+IkCQ1qN3Fncn35xSpBencREIjAweYNOegHBQA
GPBtsgEARSG/MDl6LOIwPxpBZnIMiOB1RLaBE7V97e/iO251AV2LDEnT86lBAAPN
hnzwzr//eWSe/mNNwk4mnai0fgjMCXFYC2dYrAUhqPMr2M+754h8XkQzZK4A8RRW
4+JcGQ+QW5KpxH+zShABiTM/vina3MVJW92wDrBgUrXHbRhk1QpO1/ju/DVW1SKI
hZfX44wVDV2mhLQOZYFO2kmovXqZh6gllyB/0raza0ndBS+/9cbKK/j6tO+j1HJb
0Bb53pc2/3esOvIqtKNqDqVqbQizoSM3nZtIXEBrvUUIUNrDecxI8IsmYZvMHxyb
tGks75yCwhDJo+mQFy7HDGDKMVW22ZtR/mEOKAi3TNOJ62UrSrmyr0jwxLNqUQeX
r/T2PT+3EwfkZgI0vC3sR2hHDsmifbcKJfyCTXThAPc33GxpuDne0klCeij2ZFeL
culzdJJftSPkpt5kiKYRh+yZrBJAmWlHFb65HdDarRDz6T4+h5IXCvANltu1bZzM
fvp/3wgJrsq5jI8IcRpuJ/5yltpz0gav8dXwpoZzpBKaAZlMc+tEbCQH6ddMjWef
USJMPpU9MRcDwM8CLZaygjUh7YDofckTKdoNZa4XQoKL/cht2LkNpkKFPTyzCJBW
dCfjGrktQ8y4jBezB3uShGtg3mttkzKmRAIWKFrOWnI00yxoPaC+49tghLb+ZVo2
yeT5LrXPoS+v65Q2gYyWYDOrwMc/82vnFzKTxulVb8LFoESUCg+3WYdKwKajMEy9
Zo+TxD9mYtvorMKzMhvgp9vW0kQUSaJA9uArTxR77b8ba/G1xkG3qXx989mvCeSM
G0Vt7Evj3vGELcelZlBBpe2CyLnTkYKxhnp1It+6m20Rs5kcm8CGz/GCQtoU3FSb
UETEpHA+/4GaAEe4wfcoXAGV2DNJePNXb6nhoz8y3pZflIjXwY5GlegCmun2P6hr
7+KLypNkaZsCJflZkCNRd78lmJfXLK3qJyrZPseca6tAfAxQu2iT6iSPEjKQBnKN
P/KqxEZtnlbHhYmlyiQ5rUekB9v5nqNCn0VeemPlmkHJyTyzhrGm6PDPDmudGQ75
BjkYQdMitF0cddoyCwGSR/rIQ+bZpEHIp0v+aSmI/TvpEbAQJWKZKsevVbZx9u28
EwsNh3DCC6FMOoGru7NqTuvSjhnM8M/2ZeXUmMspQMHvNGL7sdy2kP3AishAiByk
OmwyfWwozpesx4yUTCoMt5zqR9GfK7znX2XmxB1RfW+VGh1bTNIunyyQC77owDHj
U/yeQncvcWy41z/toCHNkQ2v9BqJhY514IYc3acOyZ8+LzTuJDlciz01eIoMbl7q
lflRFHIyI4moy8C4v1tBm2BUeDVHjwuW9ge4d5LzOFbK5xUy6XS0pNXMzpc0cTgb
d/Sr165m1BFza2qbPBb76A0cQOj9ZCl/eq9dY79VJoaL6AoJUqWky9XutxbRTnAf
6dRdK5sQH0QH1JI4Gjkr7NcOh/0TeUw9fs9Mx/WXqOOyDDodRByu6oMKoUaWYGb7
5tntl6DA73AQdXzmnxVOmUbhL1hbCRWZJqXTQiYsSaPDHFAujWp4e8qtkf2Mgivj
HH8pwn6Xo+NgRcx54hNIaQRuze55/1EsR96WPaEhG5ZLydu3EcZWoWEK1oxhBI/r
V7JwndZ6LXi8qQVOonKhDDuDtw6NUoTeXAunzWUXCxSTb6OyOkwy/LUiow/H9ZsO
NDju5YzLBo03Ov+O0iIIw3nkKRKSLaz5hwka5QIkP1o9nwpZpeH5cRhKvyLj6z7Z
Tl+FcpjNES8b+hnQSnjT/DI3B7zBQyizVF+PULRh2hiZCnRksfeE/gQAcGf7jPj0
SaaLtERp2m0y9ZO7lbyzgyH8XHWWAvrZMG6YtZdZwL+Wq5ZZgrv+reWqvAwvyT92
TGexzbz2dsqZGpGrRT0E3XQKdGeBnifLgWmmwL2vb6NeuJqUCyOiNNwB02fQVvJG
6uyL5C8ZbVLuxhipE6PI6u7u5Av6ghX6Ih/DWjvVkvs29LTzIz7p2RU937mgUU6f
Y3jT72HSw7SMEgjaO0HJbkVL5rK8XgF47svUB7GVY/ZLp14TYLamBkj5UKWCfX23
jwPfK2lvkrEWCPDqNXZGzZcU4T5RvTVz51NGb2/VOqntOnYvQM37Uh7TvJciObod
+QHzw7q3EeFYJuwKDduIMeaCRJlGZLOmtEASGhI8mPgrzmbwSLsgLpqByYEL67Vv
lhNGFCgYffDEJ+8a1pvrrb5hkrMudTfl181rcw9amWwlihmGaGEdSEh20lyUQZWD
Niu5DxqqsuThmiWH16tlQBLTQmrhfmieWouD7VaXN6oCqbTDEbngfP7C03s/YkWH
Ppaa6/vsAUeJzsefnoj38l/LycRy39iAk89r2XYRLOLZhn11H+F8lucDiTF47Mc0
TpyaqYlxb2lYUVe9Uf41XFx/YX23Ojq9MOqkjGQ7+iF/TkbwB1AqZEv1xh8WdbTj
DaF72bZMsud2Og+c9tb8uTgCgb1k+zs8Vb9GrWQWAVuSOVSN7wheKRS/UF8cbGYi
U0gw66wOXPaBSPWtydlCZFIOuezeoz5v2gRwJ8RV5cuKrDvvi3GhACqUGCq9qbJP
8St6lNnwJDhEV7QUgV/eHpNxdVB2OmK5vacISXEur+ka25JUyTIG5PZKbAHmYDIz
tLvj92SAt7qdvleI3EJL7LW4aj+kePPm46pR1CzkAN44e300oWPZOHv5BTD97xkB
x70D+qyg8GpuWOmROt4/hjB5d/XjD16X33lrRdAX1TL+NwWv0hiHkOJXQvoZChgI
wSEGJit3pABTkqp3UA/QCn+p2NIVZhlLfLkQuNA007DeO1JLfSRLowDB+hL8W2T2
RoNmFYvwR2jFMCmAKz+qIVCrVgf6hrWZBwAI21cThmsYQNh7vmB4oxYQHBnsUl4I
gvDxOZT+729ijVgMB38QrQb+bPMnNbtln03V7m73ybCxE6AbZUPpg7CKOF7hs5xK
CJ/q1Jl9H4gH+2ueXODs0QZLehaJnFln/yT83PCsSEieAHIL364xEy17cHUR5jBk
zxKiU6GPQXaGds6ya1T0pTsv2XY7IFp6iw4DlO52IMT9kRuD3linWLW3JWMNx08+
INzecovBzGtKfyn2BE8U6RqboqcLb/50PK50Ma50ZQSq7LWuS/BMqvvhcXyvwCnT
0R3qjeVUr+qPpovzmwJAhVx4TBp+SIl6pSARzO/Pqbe0oU1Qd/IC5RHFsZXeg/5P
ugnKDaADX+5dazZEZtSCToIN3qfOojHpns4tpEJrEjyJlVurXEIlPkwV2Df1hJVs
pm7xNc/HpyXhvfB2g01iZ8/xkRbPZAf0iOokR8JtZe0JtVdmKg0LKQDWj3CXP2xT
4vzqAEVDV+rKmj/Vuen5C7WvR5OzYqtHxPfswZBQ/AVP+a1miv0uhc6TOMXS5BWe
2+1mxzaV63J5XPuJWsT3zGCDuDx4GK3E2QGIsBVo/GclwVDDj/PZUnRaFAM+F0WE
L2yJk9azJLUZp9+4nvobdtR9QlXtQ5l4e+N1SK4KnIYsL2VEZUghWQIIDUi/c9sn
gDMaOR51xaVKRSXs8NNxuk6IpXz9wGVbi7hrEuTJeya48Xugsnpvz5CHD7idTtqw
KeYRqneYBZVS9+ntrlvBHg5EO+uJ6gfsZ8EB51B6P4HtsDIR/A/6F7Hqv2v1cmLj
FHVih8s/RMeRGpdqsQO4NI3B3iKr6sW5Uo5Z2QOjhZllD1DBCfm4XU1i1sOmSSF+
4UK0W0RI53saGiB5bVkL06eQ/XQ6rtQXWPi8QHVB8aO/wtabTQUUdlIOatRdMVqe
oBIYcJD8dirXbOFK9oWwlCRpGZtW2byn0x7R4cS3nMGubpYujlbR8Q4fqiiIcS5T
yFV9VvFNvhAqaYX8IsvpbVOvBRKpKT2O49PtYKBRwQnLuf8yxkPDnNt0OcT2u+TV
cF3uH+JzRFYSE8GMf1tcQDqoH61CSEjrwgcZuE2fCVDkYujj6x3QUYC6OFWrPuXq
iwC/tT2x+W0JZoRX35OoK0dC9OLbwhV4mLdEHtN5SLNZniyRUkm65TNyPPJL1Ezq
uGCMET9Oar7RknG86VOo2q1VN56sc7DBu+HhpGzqiwF8J+bANNbV8ghLwjUg3xR/
MgkuHLvr7ae4m4mgkb7UTdKzUoAj8rJZuh2c+UWXGhe8PR4Jl0YgrPWHkWXRS3dq
vo6BDyUwD2YDhrqp3ecsZS/lRkCgeZ78v1zffgwf6mNZCL7NJ4ACHzCDnfPfUS/q
V0UdZdU6NfFfExbh4GtvnwDNilYyWQUZkBi0icQNHpkAYla7sDDukolewf4pl0GF
4OudhvRGt5CnXBXsGN4BcBWc2gnCJL9/boeA2+RsoYhASesNvykxFJBWnJwsHBDA
YwIuYu/IRrlR0GNu5AbD4urFrbxu1WYIw6tq5ugO0AaEnxFN4IE5sWfXSQ9C9btk
4XHbitJGD+NTBRCl4l4nZImxTog7RWN++fGRXc1rMkzGRDECJsAvmxnK4dYxuxjc
eOjEUTSqqQpbq/j0EAkx+QEbLB5OIhMovN/FGNzRX4VYHB/Lqv7tgW62wSKxPI9+
7QAHtt+c2yMRsPdlfeLrllEHgrgCgaBwioP7roWufETniWeqr1KDqCwGl76kRPWP
NtHCDBl2Vv5HUYv3Eq1BjKpeTpZsmDlQoteFOe9tg/Mt0Lblpl02xdZEOxvniwm6
iIVNyrq6Gei9zkoYwAy/0XhkZil6a5dBiKH4mZIlYIl/gbQN4feiqbjymsKFuUIG
VrCOkyj/bT6AR7MoWJfojdtqbBP6MkHOgFrdR+UMVbXonQnEBcl8UX+CP736hhsl
m6J629FN/Z9i78j59uCDcMXGBZYzDOeQjCul2AMpx44iAP4hvRCRKtRwjh2J++5a
cEs7ml+iyIcuu7eKBWxPSwRDf7phH7sBmKQKyyBR/FV3D6ucXr5baJ2uPhlpnO2o
EZsTMD1iIc7Qtcn2c9GJaYdJkYWgLHlL6VCWXTzCxQvqaRkXVe4qvWifPS3UErUM
TcYY2iAx4u54OyW8WoJuakKn5PPhpUBHAMDo8I08neIhma0P8QDXiXN8MBGEUnsg
i3IP9JwdmQ69AG4D0IRn6MSi0ugw7509MTp+8eIfe4s0sBHYHnRZNiJfY0COdmIE
WAxXQAfftUFoe56xBnhHe5kfvIWkyvY/PexsSGvmsGzqNvKTUP807WP4WbxtZJra
N/1yKoM9EQrUdFoN4QU9DgGa+BfNPBG8Qtln04U3JvGWRWKCvPaRat7D43WMrXXd
18EERF5+TL4U6CuhX4wAkCJ/F8gnc9Nek6XVtXo51sD5a/FfYWpLY3LcKKD/jNG1
EtwyBXTWk/y85+fe2jvpcUU7+WgpGbjz+UmHg1Baya9M1HArMytRel2xxbr/bdTg
Gdtl7bdjyoL9Ve8XsvDTIUXqekIP1pa9IjGGZbAJyphfwYvOYpyySorbrEUtZGkq
Mn8KTLIE0AfrLtRoDuF65no6itfWUUBntvIluy6lzX9Nn+XigzcUZ11ZCJcPzlTa
G4GnGSTLk+QKtaIor6ImlcfXwkxZvG+5eNZS+MVhjP8q7gKHKvsauP7XDrPh6kSr
AjrPzhpKUiCj4DUP4bXptT0JoPl88Qbu3JdH5g9wM7pycEs1t9Jyg3g1koEEDYSI
RDbQaA+TGCUEAlTt3lm69X4aT3lrBXqkDDUlHe7EpbD8SRK/8ZLcH9Mq59+tubx4
O1e6EUvPy7X1bLlrAKq5YTYKuV16lTEiBSXEgdTbMSWeZwGAaIOC4W1KsF6tGCJt
ZyjW4MgFuDg6rdEbKCqewqnq7cpqi4d1yK3jg/D/fa/p/F9ncqQft1PWcsKEI5Zq
DefvhZqYMXU/OaztKq4xTAowNvQcFtIe7aJXzj9dH8mq9RVRaGNgZhz8lyQ+dIoW
rKQ5QIRVRO60OENASuQ9u7secNXmpC8pBCZh9yx/fHaEYwykisz+jayXgXSXCURq
JU/ewHoHI2awDCsKgpq/O11tmTwWZQVZzqiX39oN1VQ950EiNSj8OK/C6a5uGT2e
dFwcOmF1PNOsjjYwF4+/cMiGJ5tQe4fKzXKZKsBJ27vk6DBv+6BlKyERIFt3blCg
b5E7mJ1TuU8Y4ZM1MkKPX6hv5bUxXmf0in1Z/tIj5s849Rl5QjE7PbkLjtDEchCF
6vWCBOEUZgd7spl0BnGyAUjX6uzlXmt4Peu6H5biW3vjnYNe43UdJttsR7OGwQmm
M63pNgVzCD65gPTkFFhZhLGGiU+1nhArnsgBhpFZcU9NnR6MSaee2+Tjo3Emf0gr
HkX3tE8kOLhAe1Bf7mttYu+KUE4NHofPJxBzL+nEnGXscooUcPrixie5W3l0xh1Q
NRP3vAAZI4KwSn7iJoV6ydN7frWYdkeg2ZZZv+qbPzigkb0uV2PMZ5XUtVw2cxgX
LNDcbq1O+KnaDtDYlD1BL0Vfi3Vo+pLNNMGfGX5EQCqeIH9I5JAVb9qiM6XPamSS
xSkRTx4ne2/SHFhgSel23aduFpPfU3d648EiEOThrTLxkxJ6bP4Ya2qKUDBOgkTY
LVnGtltlMtgWpsClZBP7kkBcE+b8NelfmKJGqnKviJWCZbDfM4fWpL7OTUoT30KV
aXKiXA+mw2UzMQCAAMIJuqhV4PzWQqrLIMCZXXZcljK7S1thPO8dYY4f4JvCXmxg
i6CeSvNOqoBFbWNSBAgK88cP11W7MhI/RvgCLlwnk9JBhHwRxrEE4+AllunU8IgI
RhVyUVWomY7yATPTUkLrzcblO9ZXR2KZt2/DuZBtnyyR4S++sjmVAA3EavwEkImb
2JXgOVgOYutvbmT7+u7DXD89xA9IPy+dxEOKmF7z0m8U6AKSgDSVEa9JEhp1qjMi
FtRuClCewiGSwmxg/0c60TVJqOwdTEO1XxqVJXWX8WUhkqJWl+MyRigrzjtIbFp0
3Pd7jCAEGLpLYW1kpi3GE12hkroda9YzBCKQJetoGwd7feG4ezfgQarMwuLDEReH
e7WBcd1riNnBm9jpQaxgDWsx2ZsoLbCMGrnwP2Ydl/LR/fHBAc68CgB/HU77Vt/a
7Wks8st1j2914Yp3XCqMHJMXWh8+z5yGVGl10bQXYGGx0yE3mv4AeIqVBMw+ggcy
i1tKUTNLZKyx5rE06SNIDIQ5fUYodiEwrhigQNG4Bimo/yzocn9ztvkEZO5Wr9KU
lGpfvz2Zhd7fltAh9x+GW3SdZgR8fQR86zyPb3e0HIVZmZBf4R3QZ4rWJo1+11Wv
tux8ZZmtOtAqrg5WowNEYPOthoKhQux0WdABRlHvk3ZjmGXVMCj5Nc/vtcRgE/rB
zMe8vCHZyZ13FMcgE8cT0bev+/kti1wBVg1ez302wVHHbOjBFg4zZvJJUfvYAn9s
Hxw2RHZV+VmQtXftp8vecUCt4USWFcOoBlVlFgIc1VIiS0mjHEAOI9oyk9TZrQhX
9U+eglpNIeEYPYuBIkmID0/P7YAZcbl8cI0X9YnoTJnfPofQZOqF1f5TRs4zSO5l
pTzf6wjZO5wNTZePhrUuJLS8+0WhNlQT3iHFemjMf2LvamkLDh6UstVv+BJWao0q
K3LhmzjU9dWz4FTVcUzQBVCbwyBtye+aBNn4cuSWqw2i76hos9Sc4QNzuSJoERUx
2ipMbawegLqqcpYfaVGkJ8xpckrHm31GTvEZ9fU/lsTD1+k4D97u3o4XSsGKM72q
hDAiGoutF9tFNICfLrEbGilWAPZkUVgK643pUvTrzz0w9vWCv56fcZGXoozpP8xw
rfvOjymIK8OD9sGI9deCZCa3ufhbdUuSBHuQl0Ca83R1g127xW4MvQgIfRn1ukIe
3RRLdKyJIjCDsPioD33WPy/hZv9uzaipcSAWYLgXf4lTzM6pwegTx7untutDzfXN
//Y5i7edf+TzfjEb1OcHso1xup15TnxSRM76qQSJdFHpIkB649KWB4SF3rAu1gUv
7YWu8DucNIDxxfhI90awVKY2h2lK/ivwAhqSViiA6waM00w7mYp6QzrEq0ldn0e8
gFNyVMqgrdWLp8BWxX/hUTOsr9DzmT2r+WNVCuLtcquLuk8sxX40JuCFkBQCh5Cw
+JUqG7xxyQwAsAe/rW2wwTZZTHyrWR1HrCeL6pCxLlbbYQJdxgapYpqQe+OvwxYg
gsdVr9jC7Kf9dzHsaGbEk8aigR1tvc2Bzxrl09utOmRzGCDAPCaEmUnOKRT6R6RF
GMpYApjD8XjZYA5WIeo8CNdywpYnxpnL4xc5wUPi6Eymw61mdOc1jM/8A131S0gn
Y6VgQWKkKkrRSq2JES3rtj9FOMq7pr311O71MHhZFzoQCVFuM1qk0j5wYGRd8z0V
JL4EH3rj+yZZBgxQ40z0zYWT6p1pPhJULJFqd4aJvUPnpJilYkDYQMzqworHBOY0
mfeXrubxw7E/3xTJP7aMV/qYryiz5c6a1VbxSb7FOuWdidtjCPJmkRLokmAdITyi
geTE/yPd3VHUO1kEJwlv1ueRh1bEtF0Vh3nBuSd2Mg42FjxcpccuRrgHHartS993
wcQsXxfNkohNzmyGVjy8BcEUl+auXWo1C/rxnZDI6Z1qj4wjOQ3Pa9WMHggb8c05
A/Zqw187yjHBW0fQxYFbfA6tIZPrQ4+jMabaYg6b95WnoTiNz2Wfh058PKm+n1PA
v9Pr1O0rukfKf1oyk2qmpI/cbX5r4+mmfUulICdBJyFcRRkJc8K5DTL+vI1xCj8y
JoRIjfKrnxBAqskS1nqVidlgmToW/y27lTfHKweXzR2xeGJ+fhhymbrotaxk/uBB
DXRW7rh/vqI6ceruPnPyUG3QG4hdmEnBXnBge5dBmQozESFXkSxk8a18+WR/X2sE
4AnxJoaisOKoZdsZA2e2P/gm2j1tZOtj2kPN7f4cTUZtD+nBBDCvS/nbafu/3/LA
pOpPZ4QXOF/CgPoMPqTrKL48n+2U9O6CB2dr1NixQOerfsu5gtMtj6REk29v9UUk
XUceHX5E6UR0eg0TFi1pTN1rq3mJv3hsnBhdvNDVYLzjL5e21AZaHSV0HF+AKesV
DTxYD5fbaewvXD7c7TSt3c2oUkO4+DmfIe8r2XlZs/3EDuqrLG2uYcvU4ZitLSJL
x/bf0wcRFdMp8aHUDAck4R1nLSZkON3ZBhvkXD/2SU9mKZ4b0Kw7yaLcBaf3aVOd
zQKgbq1422FvCFPexbTdqy0YDgeTtL//V+4uzd3QyuEyouwhwl+X1K2P630DGRR0
C2o/N00oYgH9ltwVV3pfSt/Y0Wup/ewWLpZhzJs4k1K7suMoSW3w3uXMAR6BoUG+
UqMCuqOLI4St7pWgDnnFNpnLsOlg5OK77vdM4OuoYSRFHxUmqQkXkQaWgcAdXFWT
nhgKwmansfZglyB3Kt3aQQiGpeWLw58iMGg0+1fEvNSebgAX+b9SxecdGXN4JvHO
Z9ufONzHjgdFytypli3YCgNc2ziegRWsuGyhZRDyRmeYoBGf1NfoDAnuubeGOm+t
AVgOT+zOUUajAOb7JKxBdDxKq89F/q7r1qt2pdh3FdAD8yE56v2zUQWYwEupq5Bj
662zC95CB4PmryyY4YtWRWxIOnOVAz+SeJ6PdOrpjgM/f0I1NzhqFYFBYfPNmQe4
7Hj2hM3fRbQbOpV1xvClq+ayJMo+a9N6f147A4TvDM4vTpG6QN/A/O+Omz5FV7ap
+yJzntwz4fDVPLl2GkppfZj9/ZPktg8KgGmXQcsdoxojKSgIqyHgxLFp5xH7hNim
lVDBRVEfCnwHd6U38tT9ldtYd1UO/LZ69S6QHHB4P1575ZlAEfMtrGDQvS7c4r0+
4c+A39AR6NIajc+Bf5LIk33aJmwMZOGjvwwJo51QE6W1BURIxJiosNxqX9hWMyYS
UQTqwqG2DEN9rnOaQ5s5I6LR7XHtcTkIzPC6BoDM15uTlqsswBjOXY2QF46Of75A
8JCtRNWSqkBFvKWATK565N9iUTAaAM2F6R7l+WRTVaTwlpkmCIDEeX2gCINM5L06
Yn1369aGd5xawGi393/kJSCCVqi9qSHmM1QfvpUbBmL36RweEsh55ikKiAGktEqa
pscFX/s/DEOA2kI/+HzuHF6qJjwOAp36kz5CFO2dYxztVueXXUB/FufsthiXzDLN
U1tPnxA3yIo6S3JbsNTNY5Qfh8RWjY6GTB8FYXa+ZK9mX3o7lqoDQxW6XsEpZW6c
ydW8zZeORSwaQ3Ht52byy6V+Mz1D/pz2aOHKczsPJwgznHGjkRHXJDLBRzPAsoB5
pySbIULJbi4iKr6pUvER6TvxGf4nbCxH+2Nkjl0gZZod/cHY46l83LP8MTy3Fnox
1cn3oVCsFrTDWPfqhSGsKioi5trxdFpaF+g3eLFeGyWguWimeowUWKD5y6Y/C7hJ
jG+h2+6Kj0kSCmqakfNURVUu6jSabNLlOWJAOMTG9Xx2qu67STU6GegljA7jc7BS
QVAYSFJOa4NJxMOSfl6YnLN4YeHCaZB0zx18J8OpiBu8XwgVIGUNouZklKicWHWc
pTZNWAuyWCs9ABEUbcZUhxfoxtx2JD6yqeuFrpLeJTuJeYXKA249C9hVRfliI8zq
xU5dYR5EKVKw3vsb5v5T36sekVf+UqtbzFjV38ua+keLHei1Xu3nl1AcbfwHLBPb
mMAX3Kaih1ulIvhXzHYTnXG9aHIGdMyWxdFz7HSf7dsBlhZffj8iCGBWYXzEFhJc
mRHVE5Lhui+y/SLh0KvJzXAegzHzltk94Z7dWAcIFHgveufve3NnAgPsJlagQcNR
sblq61vS6G7/4HsjiWHK/dam+ue6dJtaBZsV0TOf3yhf8v7gg8GDeN5Rj+MxZLop
lQtyXHeFb6zYnGey92SbVuIhKp/B/BEa81T6bb2Xy/dLreXVFUt2jXppfY540coF
tuyIU4cHQx0k9OffGEp/zDcEXkm1gxHUOkw8BqewcEyHV2YA5P8GezKBLbpyIEpM
o3dMKTicOhCg8o2l6KlOatuqZHc61i3UfQSvMhZ/Us1+VDoem9eszUx+aDytguth
QZfNsCM7ihLcVz3idrUZbchzZwY+rNay3TxU6W4Ni2si4nz0yuDw7lT3uAz8Vfdb
rE92LTb6Zfce79t3JImGwmlfDMqYgz/tjzb+EsTJLGUx9MbhoIHrDVC4EqwRNhdC
QeuLDBO5bVF9Q/ILkJrgO/vOHJBu0Rx+r/Ujs19jMfuvXxFYxcTPBwm+kxejYjci
F7KLfsG7ldvgGHugz3SJr8F+IytIkuPsCjudkSNugYxB9udmSZkimWZ1n1m8MrIi
kSAp5jClVSOV4p/IMMCTtGgra5J3hs1ohyUofTFoh+tvcD+vj4Gb67BDXqJIXif0
1IY6H2kIp+LlGOc1f7qIm6TswuKMs49uCGLoFRbguKFp1gwM9E+B/rI+7/nFbOhU
SCXRDYDDzgtKhIIwy+/msNc9Jf5RSXTFqnIudMG+kCUAOqvmICLwgxcT+M0rmhde
jqk0aID8rYlWLogPoE/OvKFOYNbf+P8aZnfcwlZzqQOGTkeUvrLQ2DrhLBH81joU
KeZ4oGL3sDRNXenVgmHUFVcPOpDJk31q5TbDOchP5hxUXRP1dXc26VMji0J2Lfgb
dAVTGlKC2PkFQLWhssMydGe/6XN4brZDKhWSs2f2a1ls2+iijCQoLr5dI6CCjzjt
k+jBm/kGh+44ZwRJIgP+UdZKAJ1etAc1yAXL0xncynuQhRJ4BMwfHno3eZTofLdq
n9PayZC+HaFW9sAf/ZvcX17cxfKOcF2Ltn6iimWAPEXCdBsdB1b9HJU9LZ3uhwUE
0FReF2M1cB0KOA0QwXrRzlrNG+SLkrnhWeXhNmeKjuejMhf5IE9MTFlXJL6vjyES
Wg3vWKyIWkm8PcYKMJbL19+nXNV+lHqzQeOD93XeKIQQ+BYDXPK2+r8z1WbgkpDB
I/8d07kQO9q0ib3BPOKy1FDzHqt8UadiyNkBpFlwcM6CDadYP6p3MyYfunt4Uqze
x610V31u0tNAvCCM59DbOzF8Iq1C/+5mzlTi9eJaLr3SbB5h95fsR49G290s6o11
Q2I9eyFW4vXaIVyk6L8/U98BE/RbpZ9qHkMvCl4NoAfhvXaIF7QX6TuRY+rsSskE
23Ve0DjYGF443mAdGcFzm3gNP7xZrMvbwYnC9cB+n42KZ542PA+FLZM+D6SNdg5h
U3EYtYwg3idLo7N/14t2XRo3/BW84MEcBhbrU/y9rs9zzfyrU7vBkLh0zsYF9zEp
241JVBwgwaSRG05DcIYRBVw01/xL+zdhU4aG0DVjVpObmvFayVW33N75rPRUm5kk
Il8L+bYQNnPdqtcq8bt9IDuVhNIIeekQQ0qtM67dT7nqi0aH4sakt3toV/wcGwgM
OuJ2MPo+cLzt/+zAkw43JGulfQTXMRwghn2I8IxpyJRBbASh3Hb3hSksyIfAzbBE
0ft074mZghenCREpR8Trv9eSKBQH6mnymJAsWTh+7oXm4SkQBKqrsILZ+ub9Z1GJ
QY20UTYxrRE/zmUODts2VUeJ9jIbdJobJgpb6RUhvNkIYTCATp77wDCdzHFRBl5v
N0YVjggnAtkvRZWcKwhyb2onvfuMbV6H7tlAFX50QgWphN4HNQKO5Oa/KQhCmj8T
vXY9i0jlPSNmtDbX7NZV7i4e1teEt0cg3Uy174lfI7TdbZCr6RRTG3C87aQw8w3c
d13D+X+TFxX0N2gWOkrIOjLK5Jhsr5Oxmro2dG7XmmQ7noQAzEeD5JeDJ9mpOQLi
lbV1/03Uu8angU9WICjnznKLg8tjP4ZqP+H4C1ZKHgndV/USLXGYcIsNNMrStGxP
+mIleNCzmRgHjyKA9vGiIw1lxCLvfqmPWG+0htbcpW8sdCUML+zivxTXVOOcbOe8
fEMUYHHiFdY6oLGIKjo8s5w/fBUz/XJXBJGOfBprINmD1/ERMV7BjKZbfq4zSY4L
dSkghgv3/yUJ/XMbJL/pGuqRGE2AitCfXdxLxW89W6ulWovYPFLtzmDSpJMC0+6X
/mdln/uLUAw5rNvw8Pp47P7RRzfQAUuSHOhQu/3hKr3nQIE7877/ZmkYJxZbYtZF
33nspNTvlJY2M4/Ygx4pzfYy3HJ1XQyxbW/VgX9133JKgrqLDMsuMtqVecLzsQNO
dshnif2elIP7Qe5Sr3YQHP7nzN3/Z20IrF4AXwQhd0lmoRu2Vivht+FpP3Qls9+E
/SxuFU5qYlFXkFZGGheMPmgZowEBoHodgufEltaQdtnvukOg9Wv/P4baGjV3K3tL
LIos2NJfHrIfZzEElhQucPzf1iVp+Pf50icpSVmdARHHYhyNMn9GDpFhy6R2gtqw
VmqQwEeGVszlmPRXpy8t0mqx/rrilqQ3bxg0xIVGNvWE/htT38+mewoXbSOBk9jU
KalSiveWNmy7hvLQaiT4ee3xlV8xr9IOAYTQlXIq0FuTwl46lbnHXdo0SEpO1bq1
gLGyJkmsX6xfsomKfD0WKqgSG5oMeRlNih4UYVsKn8awTI+G4m15D1uxamdR1tuj
uFowFyd5un5C9QfcLA7kaOe8gG6H5qKcwCcp4OmTsKezC6pasfo5YgWKjTMilop9
QeOmapxq/JhSukjxeTwviw9E1SGHdDOaxQyoFd4bV+91RhLgjIDtfeC+gt5N/rvt
M8CBAej/LQWYgRxVuOVh0mS4t1mjm38jZ61FYLz8xbgEBOYo7yIEBC+GEimZdAaO
LJ1K+aY9mA1HDuenfkfKY0VZqG+EoYdIOzgEVTCV76Jecp6fGN7noCUCLU5HUjgo
b8A+x22cOTCP4bVKLX7t5Pgikiv8jhp7zZpAFEBs13oKT2/8vmNRk+6AX+TTRRim
QuL6yHnbxbtIkjCUobG+iw3XWYA4a/0G23DEwPlkX+sbqcAs1ySahGCQNQp5feHA
3CqMLpJpp+Dt/PJjLQ05RJCu6CS4g+K3cRiRT1xSfMkMJAaNjnxdCU8DK3fRWdJp
537tCrAPFcyYWfQ7fvU2rORU1OSYWqe3MzfN0XnoCFHDDS0pjjSzK8JswyBie1AV
XfT+3Eaftqne4lvtrPovu6hA1s5DY+rkpiuBivRh4u1y6bfhxyjKZfYucEkCH/jP
I8Fu3/e2Cp4brDQNlOmN1nlVhYjge/3KW65dPtBSbZWPO2a/jgyYOeUVIU7hzIUS
l0idu++RBsoYJnvrb8aNfER/cBgeKZRImBHfLStl0FhWVuyzxJjOJ8zozj0O7wiL
2ZMx+XNh1EXe6JLUwsXFR24uk4DO7sQ6LmWvrq28icCEMZ8BrG3DpBrSidagpmNL
oYcVmRQ9Vcmfb2tPI25E3Etd6G6fTx29OszV7aA1brE6wiIZXKl/Dh6KSPT2pjMe
QHOr6S1H/TFLYxEliJXpO9vZfQFdPXSqDR1xdK370bVjGywPIxVlRPxjHLC8qMJY
dKgljt5lNZdBt+hpboGas8Kn2AJF+bQ4w95XkRfpbWpYYCRaqbZY5B0tW82mbGa8
C8JQzzAjjZxh597ER7zW+CrzIyMGy7/3b6SXoxs6ofeW/Rv4r9SJizuLB+en2ScL
fvU5V30aIVKUJY9VYxaCiIOhTsY1RhGfuzwIyNvXV6/ls9XNOoqeZ8wct55i+dPE
tzQhkXP5Zqjxj5eaRkTlYQEeSe57g5H5LioEgo1p+hJ6kyzfktQmuKexXUIUfNw9
a/7l7ZTI1Unm8T7E1N0XgCLhj0CfyROqaNz7/pxRvz3lGUGRVeNQcjaHaTLxl7gx
VrTygaJFB+HL8bl5QQpXXXmfkeKt6/XOxj1PMucNKVMw56vDDJUyPXW4Lty5Z0o8
aEx4FLfipueCg+622QEGvi8iXx41aq47BblJo/gFdFK6ukFV+3uhjb40YvwF9+Di
Ycd69ddwu4twnfCJDHV3B6BBDu96f07ynjhP3ot8waYY5j46ad7UBk2zpXU27HWt
KiPtM9DTRbflytPPx6sD1EgTM8FZaZne+4muJwZ6pR9KVz3nnAfVesgcSEGMKkUd
mdNPMKCXxe2jS1VUalRFfwU9X2QIRWt3+/200q2rKac7sYt0yvYowngnmnQA+bpj
Z+VE9PgGHwC8OcqzAJaGJyHjrj+R6Z4sUJdQdIGvKQw91eh+tRuQ0V7TGTmSorJS
S2icOFTmQr+BbX5fjH6E1kDmPLj6ZO7mUR0F9rSCl8kLHDbCsgEv9MXGeI/K3b/6
ZdubXqYpiOXxaakQZz+pVlKlxsPMLdthJh5rEU2IhxGTN6Sf46aaC6vliDlq/uQQ
Pe5WR/orMoHZpKFXCvvBiHOqjZBUl3z02ADvQAS+FaQhtgjLUPaxhjIfaE6sI+P9
gT7sjrLYIrFAwsAlpMRqjSaEuy8MNuse4mHAUXvYAG1ZZOVaD0ToS3EoNjeePd7v
Thnwh53Y98wZB/pCu3bbfiEKLe9zxDDRbw64+0/axRrNBZ7vsoSIx09OnWp763hb
0M8O99tPjC+O1p+4VEQeIYvd1tCSu1ght3IBiFH2E167Yj2DBw9ApWKiC3fX1Ga9
Jysesg6UYfJn4379zEw4tkpTnRBgQfT+LsbR+wXGapLXXJ9c5Z8BKfXse1O/yqvp
HZPu2azYwrlebud4J+JVI/2ZBOT+CHwibIkwGw1anh/ZJivsj2jcSgDQQ8zC8MqL
ug1+h+1zYwwynTT1t0oNx3ihCLXQq6iBQTrUr7H1iHnT/uXGaNl6cwYhLL5LsBkL
T0tdYSr1oX84b7w9MzI8YJGxw6EjqSxD05ojER8RQyGOy80aFpmIzBzVAY7T97Ms
ZeWe/HDamDy08i4gSGdM3KgSink4yqURakxSRE8IADwpi8pp2PWnm9YVke1tbIDq
7xdtvQD+xUU6QcPzUB3PLpIDUtU+fGCGQCvZJwjAByThtLG2Sx4N9cWUpqFRsR79
gLPAExMmbHtyMqjhHFJqvJiyHr7wjjFshR1zqa59c+75N77Mbrj8kVKUGA6ASkOI
hXT3Am1J+37+kB0Qn6h7nUMtN9U7IK9VhsJGJYyjLZVN/lPDegec+c67yQ3hpMLo
QBjmLJccVG/ELIr4L+Of8mLl/DEB7ijKQLTMr3RZSOE4s7ZTo1eygudBqm6IZRYD
TgnFY5DubO6hnC6rvi0oA02/dAOLhZoAORUgwxzJxdhkJryFrHF0NM/xuUY1POoe
Lc+SgJYNytjHuKpoprON6mRcHKKkxtG010ipBOhLL7qGeph9I4dvx3BfPPp3Wk+4
vMN8OqTRBsi8gdI0DUuo7gJKAJ9yB32vCQUjXO5ZAYJD5ApUbOStkhN6742AEw2O
7RWZYjBtjbvuArlfYz88mnoHBwTCuBEX+7fXPzsD3LLLzwXA+x9//2iE6AkH5zVt
g5RM6hlSQU0kdH3TX0qrjncixBLnxnVzL2HxNCKEyuIfcky8clh6aDaNdETe6Ibj
u6h0OvfaEfs9vu/4bzDmyMRfTflvGQx5k/irgHOTUmMy2HJ8/D8XKQZKUhsf9e/F
am2giSc8XFrT5+QPSOOSlfNkNBeRHysU6f3G18maoLbrfp353EfpJ9Di0cgUFQ+M
WkjglLg1sWbBA8o0Hmm0IKmOwMh/Jg0a9P20ZNds/Vpv1au6Zp5nbK86N7qxrxcx
DtB7xM2KdRkDO9WoC3moP9s07bu24cBbw16qWOfllewQ817cyEvGU1Jsl5Xtn/Ew
buvU001I9NLwQUblhM1RJMtqKoitIUiT11O3fzTsUBrFacE2m0pHqxIfBh+EPpDm
PcsqAiEeZz2sZxqub+ObvWDsfMSYkvLBLACrs7BTj3YE6Pc5O8mlx83Zdw82Weou
4CH34vEhu72AjGBS5UGwSE8Tj0ZAY6zR3x4MOvws+j64JS4sFDafVNDdUiVr7lsT
tNY53QDbbZ8rXzNaWrEHbhtc2dSjKFvURH0+SOXcjhqzJZ/NKxUucUNNjD63JogV
xlcMFxHKzby/Hhh/FTqCFsZHcIZdbsu4V+83lCpLNkwPrPt4N8MaH4yLujk+rZbf
xGde0TPc3CmJgi17IjYxgD6JeD25dv5QgicZLIl7gwFneQ1Bo1JiiqPJVYeZ5S7N
brDStwVQHDDYw+0RaYyyF2B8jdHDBOMiEAKwgGUMIeVQYVdOvleTsReudUPQlShj
YBPzU1WV23BrXmLkqbevGvaaemSOt/PHzmAIM9A3qVyL5qP/wyPNtpZv3TVOKZ0m
BrB++34vMuibnZ1ZbqTLvkMyaE6CV9zC+FTKEwvn3qbs74E1ihnp5yfIumurFNUn
U83PtEjN0Lq1UkPoIdOwyM1UKeJrsXyLMgrwiM120tco4DyPrmic1TmQleJE9En5
N6DLkwg4ph6WWv7lFEfCxRxppXX52ggftLVtLJcUqlU7kzzxt7+ugyQy2nYRmdd3
XsN/huq61MAqxo+x3k0fn4DSWw0vuTHKcVnD9kM62Wz9K9i8g+0xKdTH/1bLnmAe
MwfJims+5moPUCkUIAi8U8JHctPFzIsPDbR7x3ZYsiW4/OxZcwPUQ7F7QplhKY5V
vFZWHLMwRL2eR8jeLix2KwmypMBr5T1/AGVpbZJ20z0YlqK2Rnuc8wz7blutqNQq
+bzuETeujfEnc0FIov8qAR1HBwd+OfnU3c2roB+ySnTT8NWhYUDuWwdv5B14B+9k
SPqy9SVaJuRnaLIX8COcoAx2xizC7irzm+jR5PYmlCQNl3pcY463aIIimEkACZda
s9ri4hqTSTBc219hLVWZdGyZtaUCm/iTktFfgetUB7HNivXiHiwWslLDmuNSuSN2
f0l+S102q5LY2/eLqXwV1DtnxWUGgY+a09HIvaVtnDcujEGS8rS5nV1FjmHqZwFr
Lcs4rFIeZSTKjlXBT+HC0A5eHUr25mhkygklO8w9WKpdk0NSnj+bbqOyOV+ALGZ+
oF8iG4zjd2PlXL3CqjEyD+Q5ZZW3ert4Tq1OnLJR+i+jl6SrblMPiQVfgIAiS/go
jhYUT2l5kRXjbCu56vbRrCKTGkmJCoTKkZb3hNmPOrutYxT5aqednuR8k8LD+uWG
dQsxGya2SgyRzGpLk9sLCn9T9m9YNhpr4/X2Hb7bCJ9laHnTFA0T49em6VJLK/U0
OieKNh8rrZwZqiLqmDxR+ucQk0ZOYBtbf6/+TBWsPSw8RhpRaLjNASrQYo1SPC8v
bvijZ8NLGMh7lBZ7qQnK5zjx7sAoNz3Iax0XpxcSLNIowxvB3thST5IElyL7V4/R
j3e4L+qoDlgnCvQ7Bd7WaVQS9vZgibUiCtq7s9Gp4Txo42cYTN4mbj30VR/op436
O473Qw4WLcAMlyfACKEd87ohwEMuRABm2yqBP8TvbgvHELXwghx9qgHz56LxIJgC
0iJAZCw9Iy0BeE3kkaQ/DkqeaqAqCcoe7YOO6MycAlXkT+xgHIpR60YS2b64XZFb
SJPhQvANsMIp5QhTgxdM9J2if6tiIa8nZ+kQilV5Zj3Z5wlX1QM/EMgPq7Cs0qrk
WXHLolNFOLjlEdRIQzUZ18c5LXgC44r4MRJjo1QUi40cexVdhp9lIwx0EbyI5t77
oDGem71dWcdSwI1apbhniCZLPwooT1gaz77D/GHK7yEjVHHRZ84VS7oLqW52IPc1
eivQrCRS0ib29wXV8d4b6uFgTqi97iZrugLSyC4EArYAX2jxzHYU2BDjDCxq8RgC
TGabUFIUEzS51BomcV0/f42oc56EgD8514LiEY1ZbQNYUTHgWLHco/JnpfbNQHr6
W65s3EzuBuZAtGW7nRgHwoXSX06Z6GTv37qs/Eow8Lq8I0Ge2mIuLT3tRsUvrAUf
y3MzHs74rYaGR57hTuF2oapSxUQb9E8zkH5X7dsZeX4AQ54BgYfX4BuT/R0eFqr2
jKeY7SM6O/W3m9g3g0m0eQRCFYEovmxFDa4kGR+4QvlD/e1iLRuMoHYOiTD+1m3R
fXu88BV/4TY79RLahLkpGQM0Par+jqE5I0l4pbtI2WlPIfJObEhgZZ+vwkC1uVKD
KUjvwxKCKrGNMWSZqF65xAzqfVjC7dSmkRrRHFysynwMQyk49DxkDPSPWYgPK8rf
ub9R/HYiwvMcNb7/5ZEElq0kMTl2YTS44pZUgC7RLtS+MtXY17rAoQxagG4n7xvw
fS5qV8Rm/c42fqh73Q4KwQyYKq580T8Bua1Kmbrx1RPdkW6UZz5BwnPEVP0rev0B
akI63Y63az/AAmFrqXZZ4I3hvRdiWvEvsHlRcX1hQIOqw0xDu4krGks30mSMz9/t
ulHztUkCh0wl9Ev0Vckp9SePF4BPrq0JEwNlShLZb0ib3VRw/JvBF+5iMRfVaw61
nV7NqQHlXKy31kNWiX1l638WmyNyV2+x7yIen1Pm7rowbyqXY7OAauBHUB4gntKE
5Puwd1TkKtSG3VcYx+vwWxrqCsuxhLp3MuCcneG/iTlYWsGGksxy5DtReSjp3Cbu
jOkbstYR51jpGmmayR+hOLEtXvRyUM4f7TeJ0G8xQEtZVKmW99EWpXFE8vhSYUGP
x1uSSeB63hmP6py9DXTu2BPvhRt3K/2CuoOK9XzdEpO5Lj+DZeKXFWR63bpi519h
t6KtimSzHpZgqZmlhF+68ukL9qTqcWeUHtoYmYMPFi0gsCuMAUxgjeBTo1s3ERNb
qhbrazPSYDj65qcAvIPoIzxRy2Of3qiL4YSG9QSDkdG4F3NBo3Xm8OV3T/4brBuN
VT1mwjCyJVKXnkC4R0ymkPHZqknuL4KvWBSs3/k7n/3kY/ybbxGPvuBh4Cvd1+ie
lLeBYxKiYCcyy28CDlPIK7U0gKtCYZlc06edkVCi6SLQReHfsc/D+6nuutSatK6F
WTSGCYsxBen3vDlsDw6vUaUieKOIk4vGS4sqealRcfuLMv/fU3LiVRHm/j5PYSIR
XeUBv96A8hJ9Z27kWSTVAUVDUcWO4HQlVK+lXhen3ozey/9HQjc3ia/f6q8BpGDC
2EEQdFjiokxXDvvWy4Il/Tuw3V7BnNXEUlJOLzhF15KAgcHdghlQF0CX280sUXBm
b8PQcuH6UHdq3Kkw/u+SpC3VmhLI/x3yAqQKgO5Uxd2wHWeqrGN02aNLAVt0rD6Z
7mdSXKVcnvT341LMfbFXV3e5ZVCvINaEoBOmen+0a9+xsSMrHaBJS7cAuD5pVBhj
ZozuD/P0W6qnPjrm4EQFb7yiYPQcodrbH5xLVeIKJrZNzzyEgCmAayNGH4Xj8Y9e
uoLjjnHORTI6SV0kyKMiZIDf4NpAfceCML3mVEJBCVg5yxOzQM0GC844Vk8N95cr
G/cKZnLiItUqpxU5i2o95HVSoUnv0LhxnOUI0siMq/xJkAKIsXrLnIkjIQqJDyn5
+bQ5m9PfZakWPaIegbiaGCBcCLRfkCOtFiWyCnOkbfudVneZuarKI7R5SGprgDNz
TsHQaP7vRanaIM0ubV1i9iOZjt6p2DS0SPTPgbARw8GATQDehlgLJ3x3rucb4lRp
UEaZldcu3rYgUoT9P//xNujO+sz781yeo8a/PSlkDJAFta6pUGRSaR+Xr7uAsYlT
awqGvHKyLXtJDakcq9Rd9hPAK+upoNNtojvhuB5uxi6GY3NGjSaveRHRJnlxpchL
6Y0/cO65RSEzuiTvvSzTJ+zFAAMYgifAv1YCSE47NsmKd9KhUZ8V9jcqq6Ll4tIC
Vf6NBIsUqFI9nKjydtB8Bubavd13mmeHt+xN0X8kIi+9L2McvugfuOtj9rdWf25x
E7+V3jUh+DzYjzrndCGXG/BPC9v3laQlgg/E7yiK6i9qV/8CLeT4omG125z88aXU
LVTqElmRJ8WSzrP4VnMDWpydssPsV7i0bRNbYdPngaUZXW7reFlyYXdEpFK7EqUS
O2Wi0O3XvN/pek2LNRoMGkR3iy8/etGgjuD/yWtcrxcltM3G5XQ+fRDpJA/kod69
H3sxVqxjcgGUTamVq9JEs6U6wPwR+KH+EE9lz4knYBAjX0t/DF6NLky7sCIot3zA
FrD7leSuWS1wjJFG52k2oGWCUePkcYjyLH/nnNHsK91GzIVlg42q0wwJICfcbuj6
DatW5GavVzEEXLiY/E7YYm1zclJzdXthzn/hGlTN41Ig7Yr9k6SXiMwPgHt+45yI
5YDM0BUCAcND20W8EQL95eFpxVYn8ug2EkcBpTo1RNuXZ8KpIqO4VpMsPDMyvNwg
JZtuGpKeVGJLMmHOgvTx5fHK5rmYv7rVn5FWwNPAocBDIquAWtyg7pIECJuVOxcl
S10nJGeh3y6iLXhGAflJcYu4qhK0NvftO46gsMx27omUjRYbRnCV/CCpbD0Oofnm
8dp1SJ7pXUNVGQH/W0NJCuB4OkVwoooVstYkZJBAIbdhpseSwy8rGmBfTbpDodLR
z8+2ob5zJSN40+jLdYckbBcIkU6ipYIZ4Iy3qDG5f6eIn0pVwevuzzuV5bYjvepa
07rIT1rcLsdEom8hjEJcwOj5KBMSgmq2z9I74aNhKSZLWFDVvCbWgGhvVp4h+TT1
1dutEdtsR6KrO7QFPK00ykRvC5rwfgmzDxBDRHWo8Wli/U5V8ZpwBcq0dL3nUz8o
dPkK9ZgnufYTg1zJDPZJOfTTrp59XaR7GetswkAaVXod8uLiMJSYa2x3Ykfgsc6d
f9zh+aP5zG5K1fE5dqyt29XcIIxlJtvjfB3zzK1tuI1veYHXKrlhjT0fwbkQ7riC
VU3olt/gR+e3RUT7JaD9EAG/JRn0wFRsAA4ogh7nF/TgTQFGdHNawuIcZJ0Witgk
HKZT5RaHMV2gxZIYzlhS9PbXMhirqzYSSwfSVRxgiFsSBsA6izetyI9TGmEf75U4
TgLIH3EkpIRpaK0WGLiMko4Jcp0VZVEQ2BKMT7QApqwxrlY32mm7BvyOeucq6j79
HT2IZmbRQUwJxDvcOplDmpS4VXPM3gprtbKrcfdAlDzMAN/7gddw4MMxB/R7Piic
nV/glbg8m8g0h81owQCSVmottUkZXfHp1NsxhdNH5azZ03975riSvzb+7PoiZccD
1dmNZ2D3OljNgcXUpNt+2v1VDRKUfBcQhymGFPUBqcU9mXC+Q7XEW5/6vsCOOWuR
/sF5KFoDeImyDKkgYDt6aJlQJLEYlhaeK9NiaA17NTw9Mbb7AO2jjAA92WjrIE9f
Iu8yKUBQFpDY+LY3jqNVfEtnRn0OS4KpcwwrZfkRcRto6K8VFSFY++KDSFnwPfpE
nW28SM6Sk8tGOGjMav+WOVPRDyIT5RxhBiaQhs6sFiPPrBuywaV4/RXsvN+recOC
EFtOQ3pM/WEYiuWXgbuxN+NHjlR7ujoQEBoaDj37R3j9HQVmMrjLcTisQIqVOwGb
dn288EXc9KsgmPucoQjV7qfZPwOdgPbKV0JR9mYSEYquit1f1URM/+JUNjpXS0K7
UmRcmwuyGcfXK27PrgEZRhGORfWmua1JraKL+gjG2kD8FziDRrhqkFbzXwaSu86L
XnschudzCrWgxXUOACcY5l3INXTbbGy4dQW+BJLMA+B+Cq9HThISGhZLBUNKQPgO
84v7/LWI/t11Y6ThnWaW9uOkPykQjznOo/sX+9LbiWj1WFRCAF4S8CdQSXbGlECZ
n3wQ/2npr6AdBlpxk79xcU3Tlp60bkJqwvmZIQyyMynBBbvSbi7CVfUQTvPdUJrE
2Q537BaPLmvwFbIEJx5pMOLaFE1gymnVCF/d9L4akpHLlZXR988VbMQk0hJOTqdJ
LF3jQn30vZ8y6nxd6NBn3bVHc56xTfeGqwwAYYUp6WjFCmkLnzvAuY7n4S1vIDGh
G7ryR36idF3bGCAr0V+I7bvxxSS908acVK0esKYJ9KESXMEVPUTcJDASxQ/JEU9P
FmqIHM9ZwvEaXyR13BAlK7hzRQMQ1Ia1uDo2uHB53ypAT265SEAzt3bJjeLqRAio
w5dwDrhc8GUl9fBwCyyY8IaHad5nQBOReVuH9nu9vJUnWvDWmXTEhD0AZY0ad6Sg
uDzG74zUEGv0gOON95bO9dxAm5lI3INCKS9j6eheIF5O90rmxbSqH84MjRDcfFVR
wFHDD/sYLNB2De46oerBb4ih0HwUSLX8iA5CJydBxK6UZtHu46Aap0nte1kgs/rY
SjCmYvQChzPpBWta8tjM4yQs8CNnWChNR5AvAfY7Woz5xt4sb2wVgq7Qu5igAsJI
4qOkVnuES1s4g51d0mvCDAP07+aYmJ2qFShzTO/Hol0j+nYdc2v0XhiYPam3zKVg
HfEe/xDtqIHfjKEi0wnkUSGgyNZv17EXX65CSsC7+YrUf27PhT2COk7aUhQPYbvA
1p792S8JEPwWNhid7K0FokKA3wXhMVxXMU/qhL6ulA4GTxWQ94eNatevAnOmuiaC
S3ZfpDdqcO3sSGLDbR8XV02L4YbzQkCmF3zONxhRFpIg0hlmg6SENZZPy7XowFIl
othOzDWwlnzk9j85GoDqPDJ+qfqR8qk+Mp45TzGee5LPn+S6zViva8LVbaKGG7rs
PtZ3EJHelWnThQLyNi5akRtiKZ169vQyUjMDllg3lb7x8XcZItOdhq7oKqL/daJZ
WKw2pcy7Fcv5DZJOQvSBo+ToroVneSKI3CTPzYkDrALQdhC9MaqUcl6KC6Sw81to
6KSRgD1JHNpCtnQADyVRyKv0LYd8QHeGHR3y658XagvCLsE7h9pK/Fq+nBWxmg01
ssImd4Q/MXo4s0rQW5IA0VDXrfbweGW8bICIgOiVgVlTYAJNU2FOmm8u2uCB1qLv
DsU2VHfzyDM1Qb/v7UG3fClKGdGjn81Zg3llSFGawWQqXbAqnoJpdFqBbcYGP0td
bmT+b68D99MZGt7jhAUyFykdzESsE3wcZIxW2JLHi0yh2EHmTtinrH/bLNWslv/F
F2wUsbEMOAbeu4h0A+f4DyMAHZ0QxyLCCCaUJE3LxUlBltbjVeQWtVKJUzlUdl2L
+C9t1PLpbrYMSd8xHdtawDpLkPs6A/tlsltlLsCaSWjwIR81fwqwkUGr9YN0LU3N
zzO/vHEm9CG8tfoHXSBwxxM39UZKM0LL9875CleHG6LCgnaLXd0iQyAe6BzW/ijl
JVG1K5v338GDng0v6xldpCN+FPutKjiYRjkl6Y0tEwu0Ou7+C9kESAvrtPsByEWY
A/O3IzbaM7+bC9dupbnXLVbEKXuyZJ1UfA3FfVTHhVpr59maxrXWu65XNlcBy8gF
ntaZfKKOpB+pVvZ/2rv6MKDZBSwA0J1ReFX0tm6X81XUiIgiwJqzRx9q33W1dCtA
ONQH5NZy3Z5AuTeY/zXmT/7Ow2nW/HALWs8+uLIRVlymTFwNh+vBFBCvvK7gCeGF
gR7Myi2A5iT4zYJ98zbBwn43n1jj6JxWDrQZV5rbpIiae+/5odNaoowOWTfPKVxR
RLv3VHgp5vYIQWuqnHop1gRhVQ3DjN6ojBD6X9KxeUaSZqxZlM5FFsfVrqce6om3
qahS1ox1108tjYakJ4BJrZ3WHarLS5b56E8WPtPq6YuJYbhlR7mYuY8tLnjXCbXp
48IPWv4Aa9OdJW9EKk2WCz1KMXAHTChQ6xNPNKEkMdGRRe6UIMnQLr//XPos5gCI
h1PeuCIUCcmhci8VCB8mPsyabAMOiCEvreq2ryzGi7SCz72ylDDCLH8J9hW/93Nm
ZHpbE354/RYEbkjyWhuclg7lYPL0jFpBfOy9rFRjAfe88xIH3A0YXJCLVhsgwaS0
m2tecVnzxOeCCKG8urLMYAQj9u0ErfGZ+XZzDAAmsGu4V/mrT4AfsJsB2r43PGz5
unn4sbvp2vpNhPwPAKK6KFReaChx4ILRkf0JTUrc4pLpIz5QefZmQ8ORDvn6Xu4o
LC6I1mXiiICwDLQJGKgbrNKsGdxjXjFGHVsZIHsXAcn1Ew8ABziLZpezf37PyqtC
Sz3SBfXeNJCORxVgIb2TNXex7B8VBgLokAwV1ax3p0cK9YTW8GwldTjuvZcxyaCf
O7pLdGGKX6y0tzO12RWsRua9MLHJh4u6n/zVG4FwHV8g03VbeD7P5S9ajnSVNhb9
xOknxaajhARjX5QFKUheS8ZDA6YUI0/Zo0TnxUlNmMXLj5r0U++eISadVIvkGZGw
kOnqoT2FFnYNGH4QeTMFzSpBS4sBJiHfd5FSbeRjbidvKTtjC72Jgj+/reL3RIQe
sYoqO6W9a8cH4rkRwneiXO2u1XDXN5ae5WXuZoaG3Ko1UcawFIwgeQRc3gG+HKrE
48D4svWeJh2W7bVKhDMOU79clByHX2MJrQR+olAaZkmk1b8F8q8cZaAiJMVNl035
4VyRq2QfIhCiqemmcfnPbwz+jijareslmVWIp48DGJmODTgvSq8uuL10A1LJy9On
1r50pETL39m56ptWxXgbQdUnebbBiJcRknJS9HXxzu76c1mzZkVFEN/HUb5Wsyvu
qkb3v7KUJneQohPnlUTUVH64KhZb+r04KGMqCPO1Z4TMle9rFXdkhXqIL/IIHmil
jfvvHs6QkeCL3x3NI9zrUxKRS4QeHqP7ITz5QF7u554Sacjv4EAWkSseJXlJS2u+
CrojQvb53IF12Hs5yO2j2r5Ay5QZiDy2zM2NyKpfPofCdDHP0xWwoZiYQ59BkQ1d
GI316opqnW9Z1SfQ74sa7Yc346NT7h22B2Rl18BmuqtgW3HDccGD8qJSGKA4kVI5
aJTpjfkNHN+TfQ18Dfy/3CsbL37o4c/fE2sOlWoUQedP4s91qZE47upN9qDl3nEQ
kLgwXq2KWqD5FVv8RnrUQJ0MkrjplBMsWClN/8mv/dMUPmUj+cPZ8cuNU9pr94aL
3/4g88M2sUi0mlUZ/bqI+24VsHJdoG2LSWeZmFFy7jU+hn3tv02jvFGuJNaEYjg4
A0bw1aqmUuFl6Nu6hQ7wx7hM4ETVFQo2GddNhMgmK8KSJ5inZ+QXeomloCBsdCqd
76v+grjd4HJuyw81ytePMyKzEuFg84rmyljd3Pu9zQX01hC3yS3U275wVNSHj8qd
8oiMUB8EyHTMCbzmb2qxdLo+DwwywYFKB0JavdRIIYVNqSG0uqjLLmBjzlyTIMID
C9i1nQEmmAqs44UO0585h6BVw/gRHwc2JMLyqPZxQgPAKVWDuqcBsymhAN9vbTlt
UROjJVaiydz6mzO3Obf/3Y8fMwebPAmWXioeyAYa/SdSiTmehrqJLbkSzMrmMUIs
hXmiVITyMSYR+kGdEzHDmSzvb08ZD4aKXQYvao3sJ1K4UIrWRBDOhYMeNuuYV3wo
FvdN8Xy8FJ+b3LkP+C9c0ELrLyNKbw2RvjOnEKHQaXCKxBFxaCPkStY4BHfjaPIk
iotwgRC18GCoRNsoJkQm+AVrwxFEY7p/33a0wl321w9FhV6cvc75fXAvEJUHx9EB
mEwBl0ULFxe5yJtJw2Nn2hS40urxVAo1R+XSS/Hen6re13o1/67N8RsroaJEVyHB
TX/l7ShP+n2lyOER8VvHtJNfCCwjy+hnHQCIlhkkAc2Mki81wvvqpRwo0kluZ3Xs
pl9kEyceujr/KURDmBKHhVsz5XNh9rj4o0h0TrYfsrgydFMU1oezoxOLoGWTEfRC
86TSmNRWVV9fP6vPgEvNu046ttnh/XPtzXjhoiwbrASn/67Edj/Id1Rgy6qp8BbI
HBPD8Ms49DrfYGvNKoqTDRnGd3k+wf9eXVON4gu0EW2iVW2cQ4V2yPFUe3WBEphG
LdFsjEw0xeG2DOfLgwqa1r8fXpClkb2Z0zVRPnRUNYO9Yr4ae0wIyv72yOw82iS6
hG8AbRbh/a9/psg/Yy9T1xdBRoxoFi3S1CSlMSnLp80SP0BEzO/BWl7H6DPw2GY5
rig3i3x3bySUjTpU2+kSJo+r5kxyXbHGxzksK+LNf6iYw1vCH+UtdTWyumvipSuW
0L1l8+U92IaDTG6xXfu64WIUriZHFrmuVRFwdrXJGso37bzupDluqCNrg6rNxjCv
8eugPDDY7i3dpwv+xSAJ+a7yRDqHj/U0oRXwMb1uMf0JIuO4tGeyAabSe1sOXyYJ
c6xCo90khSmnt3YPn++MG7C9H5LgMtQbXcl3j3Rckyv+SW06w4T2e5y40GhyeJwG
HBhs9JArDpxDTgZx6XlETo84TBihe1l9sPJwyeXz0lXIvltiecDzbMbq9voNEF2/
iGVmXBo8HdAiMVkFOQVhPVWnZctHa/xLSz63+9cpc81BKbnAVLtlzCnxO0pIRCuC
xNOBr2OtucCTexy+9ohsMMTvNyTWWsuyOy1QxCpPMNAfhtYDaWTYZ6hIomeq0Qht
PvewT0/ocnkeTDI6blA9trk7ujFn1dCI5A5vHD4P65np1bbNuDo/PGHvFMcMg/wZ
MgaL1nKwinx+DfxN7iIQcO1sb+ymDyVfth4FMOGarqZF8WsM4k+KQsCD62BIOO20
U66T9ZKRRyvq2K7TScNqYZzZVIJta8SoUoArIUWEuqdmtUTbiG81N+D+r6TGhDqz
jFQJJmOexWZ8gfLVlIolPOhwdERt7vyh4ZaQ/IDn3A/0r/WuHRuS9YzriM/32rE+
GpOdPQEBsnUZTg5GDTdcr42okouQ349aX9UpeoZQXWD2EczKb6QLf+CGa2dPpnT8
i9q6Qtle62XHBCM4LTVo1HcBKf2PoSWOPLnY8gjs0ToMbTEpCQr3qwZfCKzg0peS
8ENjxpeoCIkBqf0dkNG16fib3E+hdG3ebjq7S/pN5L/VGcMmfEk6+GRaobumsVyR
z7fRylKISef8+8dqWUW65KLy7saNMbIkN2BOl00/eJQ+qp85jrEUIlEqt0b3b245
MDJGmR4O2Z4NGjBB2tVEC/OGwnYQZkkNKwEL67HIavQzPee6VD32IQ+IkXsSYWPG
pI15KcsohANfXgDrk2PwHL3jCrFAmUz2flHlFo9ioMvB+108LKBjV6RMqiLVhUqs
2hGSyHMCyyDO7VcZDFf529TUIbbWMreSsd//4fwChnciRQYMM56EcBzoof+PUozb
qAoc4I7bCkN4sTdX1R9MfkyOuZ0n8dK8zTsIK+RGUmaxTDP331pHfRqenIn8si0z
8TmaJUBoo+upqCIlmr5E7YZq1UjqplFDkaE2IOQ6I53NiYXQ0Odz8ii8Hlp0YSCB
KyTJpKUxi7FpELMR/IKN+Likw28WTX+rok2/SMMLBfN6AYwlfhYsze+PvwwYttrc
LX17Uo+O5JSoskacbUAvgQ0ati07aBCNHHxy3CsXUjbadGvLlkBHl2c0nOQOeoBk
Elutad5bb8/es/kgg9AMe0eKKx6j0o7Y3lVh/ByPu3OsP0RyCIRI72pCndNN3MYD
NN3h0ml5lK0WP00Ic+0VopGNXuUImTmxIgQZtr4aYJaeBrE4NnPZetDZDIDsZAe1
c/bt4obc3ODf85abecWstrUXxpZRFjYo/Hy3Lo7cAaHaWa+jd7P+m7JCLuz6DsWy
ZledJ3pgBJhJTFxLiAAjPwqYmJ72fqkx4LS7+/zbya0DRJQba/olSYE4KRHuoM1H
7eUq3PYvcBmLeRg/qUWrITfRy7naNhWmRFoRg5ubi5JkJtdYk1dAqgEKthUdQVzc
+SEbb+F5Te2E8c1O5G29ipQSA44+PIHiYCYCRnBVFt/CXkVC0wjxvGTJUDzIpmUe
wWGAaMieAWQIz4IHDiNfiu+CBaZmX3Z52sz6iDPhn9knaXTupBaob9BhCuPaHnWO
xgGSN66QLh3END+MjDIqMB4CSwfKk67luNcOWaaZe6H3xi1Aopx+APQTCJ0bRc9m
dYYredf50XBfFErZCAZJMhNIayuHkjEicnLa+HxRvEndnnT8muA90heYred3HVAY
hZdUsF96Mm13Vr4gd5PZPoXVWnNYl6ScsA2Ga79mg3ynUGdybP2ZM0JjCxOCKiKn
L9SGjh8BCWj23Z0+R/P4FDW8vi+aTdwUJ1csnqV7mtdO9E//MvUI07vAUzJn5Tdf
d5DAOLsurBe8BacCdjbg9InI0kS1e4PZRjGkb9mnZ3rn9iLtLW6ShYFXGssrSEo9
PVWuxv/DEcNM/l94DHwUFJGefkltzwn2uAyt/fpniq5y03kp0ViWZrc2sezUakkE
3uADnDnU+lfxWdsqwr5RYNbVW3arlVpWvmzpG1V06dB1mfTAO5gasvNPbOqu4ZEw
8dvpL4D99hHVifebehSdIlKDdQTGZqUBZwKJUpyCQ/xEB3JrxHnpl4ISgrMjuEZv
ixz5WUUXJYuAoFqBRwFZSv+IacHVfiMPGNYgPL2abm9xRmJpiwkrIug7ni7ARi8M
WVeHqEPcsYDBlriq+NRN1MM3IOgOAWnt4pAtxxaAZqde3AH8CaOXh2Isru3UjG+f
x6odJxk9D7olqVMtWnDjPBrpEbo9JMSHpq5dsH2+Tj/UBgl6Zr0y9NLXxeSZobrh
XhVaS68qDlpGPZoBO0TMuSMBOLyqba7HdrjpRjAnrGnFXP6jC33xdXW0wtz622/f
NE7/Sxr16ZNPSAKgJoBsL6BXbCrbpZ8TEJRZHwPiXjtXHohCJYmPGfa9SArtzQdg
MXI7TohkE6WqDTRO97H+QOT4r3hBRKqQUEaD6UKhv+d9q+nZ/Qy1fvL2Ou+c8M36
WgxoUnxfRYaPP/OuFei/fsHQjJTuSFNw6GjdY2pxUFrmQmvCE/uOnqWGFJr/Td/0
2SviKmmI9nxQ9q50bsH5y7sL5A2F0auhdflLFytp5odowagyJDdSNvvBQkK8oB7x
5UMuBfC+hfCY+ws3f5E8zhVD6juafaDgI7xIt6VGE3yXOLoxaG9OTNoXVdTpJsfk
f4ezkqHbIs3SsxNOqKE9L3bl4qAGf8roOIyqJrI1DhMgbhhWFwOtq6S2ZHS4ZQmx
iU3OjZIXT9D/x2cv2g1rmoUqTN3gvqW6tdZDlQtZiC/YyxFJPaap9ngJcSqLA7po
VQ4PbnwiyM3zs8k2IpO4oIiuq22btTp25ay8UXbBPlQgxlFbHobpL/N1lcruoCaT
U5L1TdYS80RDRWcS4p58ghv8YGFK0nThe0+Apc4oiPPmikXTrKx/g/XkwFZbL4Ua
la6nG4INbhzjg2eS1uedLPhMVTirVR0bMWdlcozLHs0Y8lLA/wlUJpzhFIwD6A7m
kCl5bmdXTWo8rzBUojsLxGchLYZAP2+1ap8UfRirNY1wQ+fzEFKsQwwmY7WRd4R1
zpjRSjUmx1NPbkMdJkk+oZjefAqihXr4nbmJdtXauvTRYeLA4vokYog2efDv56MZ
mMw15jCGOeGiudnEC8+CIA9lGmKnbzw55NoXqglw2Iua54P+DRMzBIBTP+PVb5Hf
/mfSbWAWGs06JKK0DUQZVAYOm/kBkzvOO9vHPdhy9Y+8pTzNwCj2LIwo3tUambuU
89Xkom7W8mRbfWXyN7Yrnz6EacyfEebRpuJm/yvWl51M77jb2K/zaiJAzBW3y4Mh
iO2lgo0f4SADAeaXrskDMxd6xmqByOSpNgyI3+uMqhAl7mLlTycvpTSkQNivHT79
Pf1GcfOttE1hKJ8kYxwFkS+3JZ5PKYZKD7Nr+Tf2b/3o4nNV/BvpM2JgMBUtD7QR
fZ8N6CsqelHCY6DQoROerOTcuzZC8kFAl3U3IfWbPvBsBZzo8lx5X/5JFk+WhwVx
ffnIN/pT8w3+0onn9sMZp55xt1R/umyjLx3BFJM87oNIBpHaQdPkyXXjAeTovwcl
gnOFdbVOkvGZKMFiz3prnljlvsxf6uqzvsQpw7vJdesFkWM0ywMWOCrj4zm34nzU
iUOhuqREuJElu2GDE/ko/FdNGcFusG6y0LvVSV7yypLvJlctKCHNjNKPe6uGIB3u
2HFGOfPcjJ9PLNXAwun34nQmAm1Dg9WYtP9raqUXaowTcF2ckrcq8SSDD+Zf+kMo
TVgzNObew7eINA+60GalQe2a5KMTelYxhSBMlVrqiyM/T7qRDYZxZW1ZUrI4vkse
KFyjlWwAhGVaPajCxDjK5RMc0rM/QLb4nwQYTor0g9w2soIYvgGAlT+9tj92OH4C
DNBvf5836Zs5nupc6Aml96GjNDZN8yiVeMVdQ9EhI+fLFFWHdfFtgRdEdki1FBH0
7AM3BeyY7aWCOeObY4HmwqGbvor/eecYM1MlBdU2c98dfFV+lfF0zRHGcmDDI7bT
ADNNkfxQOaxtnN29kkL+5kLjmA70MOUCfvvZ5lSPPufQ3LbEpq1BgyasSC8EgpQQ
BFIy27dHSARDuq2wBhBP7qEk1/dL841XXVXh2OssD7yGbWu7/h96IgAm7oJvQhtc
t52ivSc8QKIIDqM/IpjJ/+WdE38Z+n9L+cyZTKXUc+KcsRLZuWRvFYLP1ao0I/9o
/meR5JvPNDwsCN1sZLvfdoCToKxnviI3KwdGKLJ2oxcj5NMdg7vSwLwB9CMAA/1w
kDWYTU/npVIxTHlpsw6vTgYPEyv/M+Bq5y4t73hN28zc10GwUmYXmeybtafQXeCc
Pd0a3jtLXX9nkciJAT1nCtdVaqlJDgPdsp+hBwOW7pFlNo9Sc3EpMMrNlUKqyPIv
Xj0JbGOtY8ZdnaPlIaavhiGuhANGx4d+DZM3x0+5lTif8xGEJtj2CmiqUFPskDw4
mbiLOMjdWrYYl0p7wM++dNeqNAbfng+wDLDROeOeusQCDfNEpJWSX7hWkZdCg+gd
7iZHArnaPqizO21wzrWIR4dwj/mfk8Kx4kPu4ySvslPisgsGx8BlBCStXdUzpkj1
hPcThOcag+3AOIGmal8epg6HFETpiLREFUezeC6WlEAim4UwQDwpUb9QxreLMWb4
6SBZFsVdUAbajEJRto5qcVru0o0fBMQU8+S9py/DM4hGIv3TtXSx5RJC/DR/GZO/
z9KnKHQrpR3w/BsCiyRQqLEhJ2ob/yNqgTTjPICrigdPFRPiNVUfUrsXbmYwRkLX
QZo3BclwpkCKRcsZp+PBE2pvoUJR03O4+EenGPlQt3Jmdb2z9ryk7Gwmi80dxxhD
YatBNytEygAseKWLJgNt6dDGLSzE47epAc4jMi+u+PeJtTpWNWnJjSMuzUPXCE60
c5K7Yr+vh4sKDKdubF0p3KmiqC38XkFr/X1FQXK3SggmJc3MPtfejcfDtwgB7p0u
9MQxWGNKnGBVjrbaOwi424yl6Y2Pp/Mc8vrIIe73Yr/nRZAgrNx8XLtViYG5oGYm
lagEj7yF9fQAZKj1oZR2MLeMWnEYJ8hNv8RYnwd8V2PP2Hjd6Ymm5eiHS7wlSko2
P4lKKGypnY/PVU7ljSihL0VpKaytrpeIkMiXvQXtKrdeCdCnjwLfr+AAwcgcmj8+
tgNHuMlVZKe3xL8xAgGIydGCevz0PXLCgLtcS0f7Fdj+kUr1I6d51oxwU+0aAhRn
G7Q/6T0jrlDjAzjfsR2TbQrH05xYPV61uY2ztEyC68eGy6LwMEkx/mpdBfm9Uq8n
aC0ZWxsqXBN6zVBDR53sXTYySih6WMjKo198k0wRDVXvodgIb80zVsCVzdOy+uem
49U93YEQEsjuh2nBbaQv8QUFG+eFtY0xL0tuO6H3ijCaLgPKCd1aX5bi9mI9iLw8
0D35tLSD6yoK28iWCvH8t9J1I8EcD58VT7Mkf+DERCoDICtPz2NjW882gnulWYpv
4RjCmdLmm11V2oundYKPafQK+dIt0V8tZxS6E8O5YLKQnbhdDZ0Me1AYwFHilF2N
xuK2kg+H2hg/FOItp6hVV2SHarnryMpIDC9foS7c0h0ZaKZKhYjaxugExYOhHJnA
Yr0LcdxD12hTfLLciO5Dg/5y7iDSd979xtLeYTOdWO8uegM9QiMg6u02bAdJyYlS
vNDicK81WbAjlrTQcQt+oxDy+KZFYTg6PKVG1fL7S8v6YvbwLmRNXPPHWbjSXY9r
0dcuEBIZpUotwjQnPLLov39fm9l6JxTWxQwQXSNgnU7focQqhFqwwH6sXte5XAPk
D6xtECaGm98s4fc0hqjHAR5P058jgH+mL05dOWySApwPRGVbhpXlUFbIm8J+n5rl
W6QsVBZjAQdSZdnD8DGljw1F47IbrPzir8l6HRnELZxw42BntX4rHNADj8o+jnmG
V43M1eqV4jdtSwkTOQ0/Hk4hSMOE5ad9Anuhu+s2bIrQAtp35d2+nVK7fkN7VsN4
+4kGPyObg4U8kdUAxxAIMXK8poMLIM5Gj31Bd2DdJ43/tKKJEjAoJvQWf8dGlhQp
7e6Q9VA+4AyZBaK5GJ5IZVYhLf7TejdtjkXfv8cMgwgPOE062/973abzBMwlnPuY
GHi3ioeJ7l0bt7OTmyiHqKsiGK8cpQxSbYZJ7zWd3oDWfmyRZ40KDjJTcTZGiD9S
VJlM6ePCXHBeCDGf5Td4K2b2JE+ctYXNPocoejeBfJHciv2sgxcT4C+oIvccHHuZ
MZ+puF7r5Z1ry6/l+sHr9OHWpoRcuRStFKSi/y7hSOdZVPYsLklL6fnJFSZTYAxY
6pmF29qAf5Z2UdKKeuCSIo5JswA29YXsInIBrN0VxETMNzVZadV3EObOOSbCA1W1
UIX73bD2eUd+F5XYXxmExQZKeVnGHTJ8NhvEnrOw26ISlmsYOw8Ytw7wF2L14cx6
HEXJvMCwwZHIUmHzAVp9XObUHUSVDiJJFiGIDwkhUxcPjxXKy+auhG3wL5F2Ayz4
7zSds6bw6OzVIDz2eEAJa5NGlglfCvkhnMqG2xctF5Bf8D0zAOuJziW4FSj1/FpL
4rQOzZNFC6E3qPhpqHat9qRCE0MvNvNNZ1To/bGI41auVPqLgNNfhI0HEFOyIo3U
iqQJannt9x/mBmMDpcQvlhB6RVsXN55I4OIT3wPvt+g0aXjFhK6G3piYhZgvjYDF
XfIbN59goY0QBlG+gAg7Fmd37tqYMAS9qT7uleoC34mDSUmqOqy92MWPgmdD5b2s
vKjjNA4UddpSVKLUGoVX+DfI/UPTjRb2DmQ5XOQQHeJw+0JM0nRkQpcIE4fUqTVz
qo2jjzU++B4OJ2JylmxUHCHOYKVrW0EVBw6rLyMhx+dmFKVYIWTar78x9boz1SEG
EqW4eiEjnLFr+K2tyER80YiLytoPHa4vaws6wZZRpwOpH4H8Lprpoa3NU57+D4RN
HH8expz+R9jQAZkDnIB1koC6H0PEZQCbA4FHXGYpQCYygM/A2ec7gc3EB0j/pKQN
wGys12Yel4z6CJT8gCxlsLt7oDCgDbGpZAQC0DMZaYLG6JRjxQ8YpQ8fHDfbGSQz
J0GxeWS7ahdtJhHJPjnGEV0QhOMiY89zrP+vfx0pTYHGz4t0MIG/S9XRIi/yuoy9
f5s6cRc4PHkvbLj3Z9x9QXT/IKTaETdGj+g6nmUbVlsvzJn5a2oEVxL8SNfTSiZG
Nxjw8zQRjgtkhPZeZJa+P4b6sMdw1BTMemsACZQh7ir2mGY+pfywaiCNvWcT3DeT
xxUyL7kbb0vrFYkD1sDtJyE1gPwBVFiGf+oofFQY3mPfqpVH1/+ux/ocaM4aaJXH
FCsF2X59XcRnH5N/Mrzcv2sFEAS47T8KIdmIJQ62wYBUT/XCaa5nZAbLA0WLvXzy
/oQvF7zDPVKgQftFTMG086ZIRvAPrMsl1cPmRlu1qt0H3zKcbGfZ8o8Jvw7xdmOb
f9nphPYGlprOjs0arYXI56vNquDLJzfxdvFEme0YJ/HCLfHTzDrQWY4dsJ7AiF7u
lJRcGrGHiiXew+k9DA22Mtc0qrl7H1rjrWwkMKp4YyAoKNl5EzoJ5mAM9sFktpWl
kJgkweUyYOPVmCoX6rWuk/aK5bwymE2CKwEvbl6F241xZCgW/yTdn4LUxVT9N5Be
KGvbIR/3LH22IMuAwabLSBkAWKKFCv9dRWJ+/wKLKo+2fvKJnlQjozjsybyiP72G
oJSHGebk6MRscbHNPa17GFAz4FMeyhmfCoeunUXasr7p0fqhdBCn7cYrYHTr3NDP
CXlcr/PuUjeI/u5Dl5G+mQdliOITfPPMynVHlwUZAQdlGq6V8mSB5PeFksxhafbi
6Lvmu2O7i4vIjBU10+jwrqenF4h+9OwsCJ/pmCPqz0Zxf05OWH0NemITs5mV8ACf
EArPCr6dwe4Dxp8JfPNXR60a0Q9uhBY7O6cyueAmYOkmplU+AIsZscCapL4EEbxm
gHZ5lUKRsmHWj5urh7teBPAdoFU64USfuU7I5wTPEcl9g80ZReIoY098aT/wsuFM
z8kHLYPP+T1rxdw8iJU8cmhcJnKo5DpNwwImY8CnMSv1wNyTH47fvv1vC1tkOXw0
p9Xf8aJT+hzTkQzYL7pSH8VPRvZMbydW1DqDKZv8nCH/YC2pWUvyEqfQWwun69+x
utdnrjqRT64GvcAWl+OkCHG0B9BdrnJElPJHB5+k2fLe2ZJbqDpiqBPtsI41U3Jx
G/yOZQKz6U9cjUoi80rOV79ygGr8Uema17lfniWwPx6ay5jvKpVBQze/oGLZ4Y1a
T5A4hQnGyJwFLk5f2rYADnbxLwGPlF0/UUzExlOusUCuDFU56HceqgrnTQmhl9AR
3QnxjeMCEMP6iB7QCw/QzXou4nlQSkCTlpnqVukrYW+7W8+3WPp9Q+tK6BeGRENv
1CIBjL8ByF6R22Vrm98g8K2pXQa4Zirnft6f2cmfntzrOoJqaCT4Wwzm/nmHKYFL
uKP0Pjljsh3QghPavicSLdyLlQSvjErseaRvz/je653jQPoxVxPlhisV4ILrYl9e
PcMDFGftwUce62dcQb313qV85xwEUgL2rLH3bs4iTEnn8aup2zXdjppUyhgDVetp
8mGc8lgalNYHcb4Z9zxiFn0MLU12VV3eZptNjRQPrjrx+4JAKYFoijT2AsYSKwXZ
mL27gkip5/j5X77MlS9VCZagmHSdPFlQr/n9nPDgd4MvzIICqTqRWS11fkudBbbq
U3LQyLmP4ZBlD2FMVWfKNHnHkKgeH5PRsapw/N2/2ZVqlW9HCPL+PGb8ZU/tlU7L
GsEausNK/J5t0MsrmowOMHZIqUHdBabZG9vZcXViI9IwydI9ruQfb+POnXzcUoYq
K82nrZ+CTf0jaBm8l0JMttY/9wp9plqIFKFAByqUZoFOoy2IEfnynJFF0dRE2kUX
BdNtjNrIFCweyAE5rnMN4JQ7u/gTFOW/8xtmXhV3EP4uRnqRRks3hGykBxAetEeR
AoPWkX2yX9QnfhrMjoBv+L8vLj9nIyj6OCxrX8LIwzLq8Ovh7TwsoS+2kLHCtcJh
rWgthCbHmia8fuGemc5FUu2X1JPSZZoWc2BZ3/EhG7R3WXsUTCOwDvBMvuzztxZA
rzEMBWxPGM5y/nFrWPeuTO7FSakUdDmScQ5AGjKZkuihG+QWbJeX0CaNuCyajpmP
3ybBkyBEH0/DWkY38Wj/lEYqB5RDYdi4ak5X2IIX/cxPjmYSz673wGfRJB7GWEdE
/EbeDnGvmjVyJl+J/fLFfJUTwdhUyE47cpULAZYQ8mhxY1pJ5t+jNGxNtdxTr96d
Zf1Nb/RS5qC1L7giZViEAZs6AsHBNTuwBhgtqi0eq7fJhwUrxeQW7Z5Ajd8zlqHg
o6yWUpbj8HnO6JXjk5RQvUrEjtWIBA0UJkZdS0XwLoCXlMS2z4bdD6oFXDAYrQPR
76GQmGhmHvGWgDUhK4HLKFS4mgVuxsYB+m6WD7A7QFEaawmY6mmpSqXlJsqMnOsL
CR+WLAO4arHaiRfAM5HG81JQjzrm4WmS3RPuIiYXTvV2Y0o0Imrs8BEbCX6TvbyT
zZRdn1SCTeWtnzHWdKJ1DqS3Bu4zbPWx2lvfAxjS0flypbzkKf/5l+WMazt6IgTo
Vv4ndEeW7i/OiutAsjG7Z5djZrsuLuH+3cNHRZOHBnKmY8UPpmsp6QugShdgBJSc
k1u/5oyOQSgxYjn0t0PzQPZMXZpS3Cut5zffa11ESjNmG/gtDH2ccVGuattK/fXo
U9WbiFTSX5s+UM2nXV/4eGcVFgdY9755k7X89f3PNGqrHy+wrU9PVlReILWGOFm+
lPpUa99U5M8TMJQuNGwYHHRBluUwRYFcM5YBIuuQeHBL6pZkaR+BM6Zk6RNMjrHT
eaiOe3FIyaSF57i2DN07tXgtr6lILtaMlzZjgHn6/F08lhea7E4z36aSBgsQH8X5
eKlHkiRvvyiQDvI5/PEitNeOWWP7hOP2kSbgVGvBePvak575KGLo9UofWA/Nin/B
nmENmu8W8JCxCEshvw/GDOQqpVXgiIqSOQExWAi9yS8OCh9oI45foDsp7REuIQvD
chbR6fxlhoQlqo6BskIl3W0nivOs8iSvrGshv6TqagiO05qrcTYso17eNP0YP/HG
io0oNOAJPNeYqq+JlNz5V3wmx6f1bFOW/e47QSmTPRoEf19LhIWLqk5ldPY+lCNn
MpPpWP5zQeHc6vWm6Kwg847jHvY+m8QaHJvhp6FenVEsa+msV8boB0QKZtqOvhtH
3cPKcwG62p3VuufDGMQ5rTtcBIiHVunHyO7NfOZWfmbclQi0GqxqtrHW/vQYbI1L
cDh2UFY1fSq0XWL821LssOaRMHQl4JNuSZMSpkeo3ga8TC05jqhI+g4HpmhMtksx
ZDlL90l2U5EcXO2QQz2Lmd1/YT/tpvY17WAXE1ELsuvP2/XgkcL/v0HkLHfcQHqa
mvw+nNdYM5Knz7e434oG2Q7c85xZEKcYk12/Cn07UHvCq4D6dSrveumueQOE2Lnc
5xGUXOEvgu0vfKIsTwGdwbuJ08r/pOcEpN6muPh0UL8wc9zJ0aarXIWne7q/6Iyj
gJHN+Rtd+90JgaRobFvO7msLQZqUopWqP8OAcPbaIYl9F2Ly/Oik+PQVsbT6W0Xm
y/bSxHrNbjlYfuJkUkpPHM3e64gqp/DB0bEHnPnRmMKrD6mWOMq9pXVD5nL8YEgW
FcZtqef7ncXTulWAb+Nv1DDogfZBoLB12W9SvYExfngzdt9lVE5a6+JxKiYO9vUa
LnhWn8mWhuECV4R87Pyi5Ed4aOrRt8CNipiJT4I36MQ0AqB6jAOFdkAyCzurwiX7
MG5OapXfwtS5tMWXSxEjd/ix6Hj60F36iBPPkMUaPLxZ7IVjef3gPsfGW6BP9dHH
w9H4kR+3ZmvQO1PObHvgAuNW294+ICCKBq/8nGkmfGcANL0gB5/li+2kYDdkc/Xc
fojsVXBDQ72n22TKUSGo3C4Od0uKAfgoewVtdDfV6iIdSf00Cejq9ewIFV+tNcUj
0KzGfe11/2L6sYhBFXVDbs+OPHcXvpGrIVKSio0TINDKj9gNR8crDL6StWJMEmru
SFT+mpyiQQpi2dA43fzYKvtfsQ6cuSloXKq5nyk7SC9rJJUi3ignVi1YDcH/SVEu
/GE6FsdDESEWpgh1Nz7rEicZ0woabu2lvT3PYLj2sjmroPRvAsSO+8BjwraulIAX
LTISbJGzuGfFVasPv/M72IWHyQNEq44MyLNVGxZDHDU4Z29QMjoLcPB4j47xNHO6
R6aonMBpXoYhyRZWeb3LJ/K/SNDe/iGY5ywDExNWY5J9OdU52labssknFrGN2ZGy
nP9xzT8nhCQlg7F2ZPLTRofh+Yg6Xf1PJttpythu6BM14er8exFxusqYEDCoxWzA
fL57CtMAaK14ooW0yxLuDdzcJKT47USyf6xD+jQFCf1842LGAdH0AlFpaMSyZsCW
klfE4e6c7O0cW5djBI8oCqtMam+1hsj1vJWJhhnp5pwLHGoiaM16LGcP0KCecofq
B4Hs7pjzKE0CatHJpWyNuRs9xjPnMJVjWZ0QttSS86VOrhesTQJHuvEYFgnT06fL
YWHpNgLd8Hn+YydECv25RTSlAKYQhc9VYv5OgiVdBj5fpYBryXhnyUmM6q1FHzFT
QWU8af2MnJZrWEGcqQV5jV3GTrKVZo+aexoi6DuS8V3D9lbNevmZ9GLSE3G91IeW
6dXF1g9mYOFWgMNXuy/in4pFRMyKlePqhJS86cI9nBSq054Thlj35mexpubwsbN7
qv4HKOKpV2dWRKL8jcTloCqAfEfpexWoxpynyN3Kb8/dlicrHNwCwbFwkn+SzqXE
15P6abLKXG/okiFMho+VZWJNRIWFG1p+8xDn1tVjHEO8qeqD286RAvI15zN7qYdA
kWuhGyH3koTxOrC5Kif6NrwoI4kcL4WGo9gu7lv6mN1zGe19FwAJC7IfqgygrUHQ
aNDmhHgk3QUtTFpPIsoJygjIKn1XyJTbMmst/r8Y8iVhHKF3VDD1uPhy78lejAzB
rgkI+K+p8OOtGlCP3jTi/M2avNix3KxO6mvCl4PGmt0G8V1XMb+0ckp7vMghRdKz
kFclalnZ70WxBIJzBFUtaBCD8lvBvJ15iTGw6hTFwgHyYsOQH7rxw4oQeyWcA+S0
uZSKAYWob0Cos9YSikKe8fX7MRjY81m+LYOEy9Yn63mnbfkXarYJ6e/fVOsicMHK
JDb8LpSFC0p0GWpmZGQ8d3kP8GkbSoSpEPrxLAEn6/uYgPHuUvlspWDyy0GtbJVa
qb1uWRVLS9ibk2yL4U7sI48iR9ErjnAwMqU/kbvyQ38nkqYgGPs+wCUwHnaP32b3
1PjOsCD7RpmYQxbyukB8UMO7uQZs4CH/B8dsBUacaCuRUKL23gbyAQRL17tpZZhP
n1ULbkQ5c+BMbSN78w9lrbIjml+lPUFGhrVT8vfPXekosrQkon61zx30bEazcvj4
cbthIoKy7kVTs7nbbtkEghopFnTsEBIiQ6QN+KMGYkx/ig79eaNOq+3bYEf05Tqk
S9Lefz7wnM57C0hfcQ2uzCDpVHbSFNmBC0caiV6CtiCQ6ujzRlAq4UnPotZXGMTw
jWQ4cSi4mj5Vu3dnKa5S5A33k9TN/lPcyE3doB5U5PAXls0qGu9eOsLhvPLwmGDP
UtHT9PnrWaDazutgoN31UawwSYf5QpbrxNa7BNJMW7fy6QEnEO9r9OcN5naXOFm9
H3SQ7hhUwFqZZSsmny4OZ6aPBsXueqFmR3rPmnm7W7V0WMVFCgo24nJdVHrpEDak
ejbicp591VaHy0/gMlgvEQdzEOI/WiNr8qR31X5kIFPb2lQD0nykEHiX9HOUgDqJ
OOdo8bjOzwZ+BGW5lLVL4XOVVg85AAlsnF4xh2HfJtEIpuEOC2wWqG+lLxdM500S
OQdLSz2l5nrpepqcHGTQzAFBBxUt9biCq0ig/1zZgU5fF7xmCxuxIqIdEWJfaLRG
KVqeu7Q34litTPzf7mmfT4QsiokspJ9vYlrDgDaUoq5UbMiXiZKVZXK0/YuBQTCj
9JjIbhKCHpl4lXMUjlSTK9mo/LpWH8QwbS/5df5R9Il4mI9qsqxQ8mgXSu92+k46
qMrVxd0wwDrWqyhFeMbPtSCiuF8Pl01FHMh2Q2V+1E0waC+kzyk+PmxHBB88VeiR
DpjsNFhMZ128S2IpvgSwOKz5jyYV6wMmweN0TV530CmrfkZy5kcXVmioBqxFR9o2
aX30b9t/KPUv3IUsJ8fj9CQ7SzU9ai4Vb5pvx2fJx46jrHOhlPG/Kil9in839Ktu
6CH9QgMlX8Tj0U1PLeYdFAYGyBfSr2kT30A+a10NF33/HjLFpdp+C3WdEnrLVkx3
5sgcgS7eoK+iKBcDxN2ejTJiACBi2wSVhHQt5SfiDin3Cl9S46keUQtMKuQ+QdDw
4kQYoYXWe1XB0T3jrErGQRNitP7wIkxS45zMPBefgGDs7QBCBrzeKYeCJTSxvOjX
k7Y76Iei2fRnbMbdUBtxjVrbPeOODFK50Xqw6H5+cMlY9DHu0VaRMopjuIsNYQIQ
4z5BkLr9wH9g/3Qrw5phhcfPeBG76N557SAN4OaMk6g/M7TghvjssarD/WsYsIP4
ei+9yMoPQyaMnWMxTUCZEQknq7G1/FerPXvL/M5SXPJm6JDsOLx7c8eAXlmH2pjJ
ptNUwy7OcReXF6wP66zqGJCyxHAJR4h6RbNq+lGWTo6J7tgCCFGonoHjBs49eSwM
ZEFI+h54l4wl11+ty/cR3L7QQkg0bsZfEPM8N83y9KDMMIgAenQl5++EaWcKpIm9
Iz9Yy6Z+NTv8coKi1rj9zyGq/vqK76537GtQZNf3+2LHRpR8s8P3JJCG33CbQQ63
bP9bfNmIml3v0aHTRUYpqcjiKEV1aJo51qPTufO3cNHpsDXpRSlj9IJOQ0KrEm+B
hDevdtgWZ2ywqkRXGjyxlhR8B7IYagmZjTyyTAQgq2o7Mc3ZT4xRMl3QpX3tBBHl
gm/u1FwscO1Mbi1lJ1i6/vTc0F64u5eKOZp9v+6GBiJVJb/yKHbHCCKksWyNp818
tBCds0nMit1d/IPMgUTpwexnKESC1z4DVj4Ke5/2NrK+FEBxkwU7NEUAaJtHiwmI
+E7TcawS3GNX3HiPAewKgSL72PUVn/lj1zB6Et82hOsu5gmCcuIP+zlxbh7oxVf4
APhetp4Nz5VdLQ1pWfg0tIXLZHfG6xiFwhq4BPujrNyF2unIWze+dLFzN4cvgxFb
6d819Y9l4kKYACccRHbwrrhb8n+Uk4zQuYTxlAb/1iJ1vSFGlCD0kXFxfJ5+ow02
miJ+VMN17IIhqpTDL2lmofqyxt5lJMStOF7zX6/GW7N//yA72SzhE3ZyEhmf8vod
hS0NAnDAi9gu30oOvWJGohzF+4MIuBpydUtSpIGaHLJzRDp4M+NS3u407ZJQ+MGo
/q/Xx1ioV6wmvuUnDFSljw11sdOB9oZxSP9tge5+8/y94lzb6Ie9q8rTM9nLhsxv
0S9mmNNjxjlQ3g3iLsyA2s6TlHZ3yjpzy1lZrjsvJxaGdy4DFiudizWpY3pXZb30
ZJs8WPdCPhrkga3NuNb3yZWBausiFued+sxSeUVIfI1moM1aynV3nMGe4vAks9X+
1Fz0gXdfyr75qLG9lZg4yCBW886/JGtylwZgMHydHsc+kAD4/wZcRJV2Z9DbZHWq
Dkns6/EltjtjBpQ0PVcrTyrVebQrcWxVB3pYr1F6LOI+rGufbsqnoUPl5w1AKPZj
d68TnkBVjkRyZUw2lK/xI5UR8gACBALP+0KseODHBJjTp05U9RZNkDtq+ISsb8t0
V/8lHJ5HW3ShnWpw76AnB4bfnGHsrmBoNn4E4/x5QWX/2x0paubTbrk6ALTLhgq0
nHkAY7CljkLZI6svJmPjI0mIkN2EPZpKS7LdyBS1VEuNcCj7gOsXWSLljR9z++dO
GjmLvlXAgWvKTYPBEKvVE0hkBNoTjVYziuqTsooqEJ70TAN8ccQKPO2Xht7jEl6G
cQl4j49g4GyhlGTud1yH1PUcSS4mfwal2+7Q+/wend8=
`protect END_PROTECTED
