`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e251fCt6NDUBIRPSE2GdXJEzBuQDVOi6X5vynAP/8x5QrYRDQk2hjuX6nZbDUgVF
B9yTjVo8qYnVD83/qrp70UUoYW5P8IvoLtJWxQba7s4Qfp9qfY4uV2nFuchmANHT
dgpJHod01a0H16gamhB6irRT9A0MBcvh134U/8flYoy1HP7GjEjPCCjqU3H6b+u7
zpw8OYwZHNLKy7QE08Q7M8x/ZjECsSNEkiiWaru00VDcRPf/GMcPPzuhhfe2yrRw
NV4mjNis2jOPDaZRIPKZR6ALKGNpTObsUIPNOgShEqEuuBRW9J1TMevFoiwR3BI5
Zd139Di6PmdnaMr7EhFzSYJuRqNScjx0/YDEeQTqE+Y4Gk22cC5hQFvVaH+fc1SW
bFALjpntLKkp2+klNNgGWIw8fc3F5pdgbF7Gl/2nNWDzcjtyPI4G16XUuy7w15ES
HxcoZd8ZiU3lWkSsu73IJVl2e3LWjNKWysHiU0W3jJKuENUKt+EvdwRlk/jUNyeg
K1Hzw8FHT+ef1uHNcioz3MaLu4tsB1t0aV7RW9WYF/KfYAu/3DInTp6SfCPBviJh
OPki6g82vWay4+ArIvwzINXeLS3Hvp19z+Mv2oaMLITBIpUNs4IlxdH2h4tjp+Rj
u7DVP20sQBYGjc9erXiJpuWnXnc/I8qBZR5svZd/0UuE49wIpi9zdUVYZ6eFhUvl
N6PfeKwyyaGNwh8NIq33KawyBt/hhSpVI6x8mZeLmQpnr2wejIjC4sZXSJfqglQb
LBPgL85JkFnNrhyv8jpO6ZQCGlWD7SgqzMgt0mzCAlyo172YJxRvgPg2VeaioM+0
9EkUlDQpm9FetoQmbYcj9gZTlzYJ+uh/RUpVX6b2yO0=
`protect END_PROTECTED
