`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/GgyhHrKQziqEteLpE5ywTxmTLhaF75BkpgfIll1y+z5coU3spm8IzkYQDBq0OvN
HFdM49CbUCVe4vNDsGDuQchczh9AmRo5atcFeVQ9S7ubyBMGzND4yXt0JUdeu17P
iTlTt3O7rT/2G4eVE9qZZuKVZuQipdi7ezYPDP+2XE/5ra+bKZi+03WD5HAa4v7X
FVdwBiB1YHM+WrDwh8d4ZvPPz/pJkbiYIYMhL/CXbp0uDx+YdC69NgTmCOlIN1xa
NomODh+qJMR33Kt3hHKhdIHbpRryNl3BQmMYb7XnVDtO/yfyWVEhMC9YUGleExLH
C+dQUu0Mst5o4Vo3YgpiY1L2Jep79ReJEulrTTCVstgidNFdLVX/tSvH+Vc69qCw
9wTVbcaW4K8V0XBk8kuGocW+wVTAng3Z8vX0L43NyD7vzwOQdeHOiJmxPfaIALqN
1881kGqe+rRbydmfeqzjb7mwknp76zpr3tHbGrZleVXfjGVvsb2KGIKzP2sgk0Bl
8wk6nnUo3EErjbVXZP+SO92GZXTYU6CJqrP1xDoKWj5VXS/xkZ7gr4yj7vUtpDN0
UmMMVK/MZrX/oB14ZXnhERCRwtpGNxjylnodgpxMoudF+Yd026pI3sXMpwIKw6kF
jLsrfDYTHlfZ8/qlchtL4Komeg4PlyCFOyjvR1Jq1KHgV//Efc7dWNfIS+q3pglr
p6qThHww7lVggkly/wOEhi8wTeW8pgfsmX/aketftufISx3M2BGnszYDKtirrv9Z
DBmC3Vbpr/vTxT76rVO/2XjEG35ir0ebWc/9t94iau3FmUJekKYjlkD94DthBzhN
w1JrkzXAzXeaf2GC0EPHVg13r7Jcl545Uobg+ltR6z+ecZ4963zXDXrfwNGumjYU
OeHGaudd3Muii2NI5jYaCm2EYKe6DyZwr4p8FvyEW1rl5LV7tGvF6mKh/pF8L9nr
LjnCotMHfIPReG2ROhZzqNuN9IvJ4s12dTugSLeytH820NpoQvKEf84V+6sSqTuq
2FTYVyqpF7k4mWP23xUO5ZgXfiVGdHgSpqudtSGAqlNYYbxFmris5WKvGGDbDlqJ
xI1MEIKNV8m93F//EFMtFiJElCPvnVqIEOmJKGjQwN4IdE7x061WFquP1O7Sh1tk
6agWr0k7A+c3uGS3vQWlIkD89XeR9hp4R2dOxyaxK4gCU6MrZkdbuq+wec9cDiwG
W2sGEykbCYHO8AvB95XPK7ae9eIgVrPZATz2aAOC8IlFGN30clyjF0S2t1ezJwpA
FOv17vY2sMkYeqPbsstuTpiHxW5chAoXvHka1jGiIQZGQrTA8RfqPEVyA+x4Io1d
qd26WmR9uByE/YUzahWGIHVldESwwRUsws3bIkIIdSSmujleTJqjb4y3QtuqlAgx
u/j6v5W9zeaAEPLsqbE1KnRyK9cgMjqk1oby0MNl+gXuusoOSYfukJFf1/8pd/T7
czbhIi3jzKOM/Dwe1vWNu0IlIrLns8iBLV/pAtbo5p0NfRaIM0JPGmeJGhq9u6kx
CciiQfK/rJeRIdP3yqQEZAu0Mc6h3GWReCNvun33FnX7mgjQDhsr7t9n6TQiJn6g
25GlcWX5GcAuyy5t6vVhUIWxdMgatrCcVNygfrhfJD5SxRSxh8NnLj1NVX8JNCvk
b+ncGerjJQWimg7amZhmWkevk72nj1CxRkFa+11nPXKqXCRjXRRz2FlkhuWk9Inl
sPX/of2nm80kgTgXLduZw2LMLm3LAD5tGogV6NM4xvJzjEIr7eCH6wvak3KPJH4Y
+advmdf/SrM8PiQApo1pys1k7yl1Bo8siWrw4bOZeXoFTPigXDz+UYi/E4ya5Uhj
60xo1CHzi65/DaTKEU4RivD90Dw5qaqllcwe6ixURLXG+z8Tx+lMV4P/IFUGTc5M
Jejcks0YLxZtLjT3zmCNgC0uC2bhghSCzt3lRZUl7iOgHv3Ze302+xoIgcCv1jBf
HiPKwmxxE4RFPmKknpI4knUeEktpAkcFCFMlmvKYNaQ0zQk3V1kRuDI9414/HKNF
KEtbWomlOiD6hkBKowlsunQH+QBARUyjK3d8UdxVNSYp99kQvPbrBTfabob0FYvF
I2mGEDhXnijQ1vjNhiUgssCBE+UwVGC8I6v/XJIOZ8Kt/F3hURY9qJPfDGzT+EVB
KUZ6VtP1Yg0j2hPfkQXgGBzouXsLkpcvS62o1f4l4wly3aBdKSFZms2GI9tbOYCL
ACSYnaycAPB+jjooXWTiE2YqLYlKO1cS9HO3WxxuyFCKNSeLoPz+RG5cg98eb8DG
Qa8Yun6RxIEZ86yEFGaraDfQCtJlRtzGpoKnTx5Z82rr6qhp67cyXCpQJCVnag/U
D8zD1We26BO8cyvgmXxV5moJek6ADx4iJy6Qf/QmO13uh1sI0X7rDVvehU5HQg81
a2kFoTy5f0S6jGciqTHwv5F0qehUKcPyQS8dIf3//DpAklx8Yc5xJ7v5s2ESbG6R
rh7+IfWATMDYvaZoXWrlRhICaqkMVKRyteg5V09pOaKtnPux0Jd0GlqUqUjYctrW
FIDsjMM4o0MpSTZTTixjg9HuJzBuVafSFX6lRyyeF8xpvHWHiK7JP8WQ+Nrgln0s
UjmfcC7oE4rs+Kfdb6WlNXIjDAnLZeU//2TWbo/OvAEZrFt4Ig/e2+x1wDJ0Dxbb
RuCLvZNk7ZroMHOiX6xMDBd6SCvpzpkyuzxw8rmBloGm5c7N0uQdqqjapvw1/SAG
ROv5MyPSU43sGA7lUAr82AUxb1qRD7BfK9++PquM0VTon6SdgCZ7OxuKqS9XnGKU
jQzPjgHDSEdQtwJb3MdDCmimFgj4SFmASTg7CzwWq6wag8wseRGHquEZ5dRYlTPD
hIMSkzCGKc4ywebPQqvsf+pGzP6V0udW2uu7K/qapZbUGGq2YOvLtb7lxwlj9B84
eRyCDZXzwIFtew3ruflEAbbYxTRQu2QrMR6P98odsh7QusQNhOCQ6bMe2o+pI0yB
hhvhHEGOmRQFiflXMcX8sACAtPaebMszOXgCV0SXwzv0/yehLdw73hQEjCayrv/E
KJl2u8KXC6aqM2ENmBXmbwnH7oQ5u5kD0gtGPG6Lpva6rgEzjLwP1MosB5S9hMuR
f6bw26jS2kcma3Iw1fPqm9z6IBprqGvWsdgt8WenxY0jV1SDVXbJi3t/hl16ir/M
yTYjg6aPqWnb1ZOFYfIoA4L0WhDzFeS0lB0pq5DUioXqJwAvd8nvsvK6E3Ni8dWk
EvoL1ZDN0zuDETKO/mYwvMXD/zEKwA8jry7Vv/qnl7xkv+qPUpW0eq9F/kD6+HX4
wYrsA/fPEVGXJs7Cntb9G1brR+ObltskI3PfBeBKH1J/+Jt1ol5nnklZwG6AR66g
u5O/atHIlWfjk9ZsXmBWGiZtDGPMaotqFCVZ5HcRGXynzg99VMmQYH3wZ0NjqqRn
OjVHRsqen7oIyw28gjU65BB8a1OtISuXJOPMLi/ZRn7rDfrzf5ftoWcwTdO/W+hQ
k3OpLv88Z1+5pKk3ecXkBso8p0fuopNn+qx721OBsnmMc6Rrj76Q3n35rkRuuVLj
GWGg1lSbsEghqHLwTsyHyh26VpO5wIziUI4ggeduIgNCUKzf+C8Ohnudlg3pH0cq
daWe0HQZsOLMyPywI4OYNtXJ8QAcgVCdI0TwJmlxuNGiQEruPG3n1WxJE1wRI3yh
FOaavfhNklKaCTltzqdplIJ7CJfE0vJGWX9sEl83FRVrwJAvFm3ORkzmDVSctr4G
paOZ6QHbb8XoK1rxuL1ROG4gcd21eVyTVwE1WwATQd4RlX8zTaLCGnlF/vZIRnAf
KrGHDvCzpaEcbgcmlfpmZcK7fBfHX8AFf0RYsqjd0hFMGJhTLj1B0HRUuNFAoZmR
qV3HnfL2z2VSQ7nop8Og9kfDwDn4p93zKiYfj2JEcVU7gVJ5bqyWyYcyRxFS5VzQ
qFoiorM+OCH5oqDoFRjcgJqxOlS9dpy4UdlJ2pbQ9Z6+44GFCtzm6V4Ug+A3+HpD
tdL1gbtMfsTyrJLM8L43FhBmYUyWuEaIj517JzgM0tu8F2An91FGAXysPTsfoYQ5
CkYDxkmmSnwN8C5L6LIjwWiSQa0sqwWPAwh+qI30TzRqUJk2LCNm27ctEOzOsm2Y
gXhJRYuEd0Q/36k8IllIXkIdAv+6/oorKm8kgZaPFa2Jg24QPZ9qDgmPgsX6XZlo
cWdCk8wWln5Udy6gns3J6nR0xIp/NDnvmcCaPFVylHg/Z0T1hSs494mruU9ivMQA
GhGaZO7M45S5OM/v8kyh+k5+8uX2ghPIOZBUzLR9KRibB3+oPRl4YvHdlTUTFI4m
qZvqMBVOw+3HedRzrcRq92l7cPZ0XqnND71kH1dC4laf8FJnVj3Nr2Ji2EzvXPMx
GMqNbgYokE70ArxwdQkHlm0a8EGpCScHDb4nUERuWAwIszpZO8+NS2ylZcyVKSwv
sY2uSSRMuCAPrxq0Nyn8Vn7h6SQdLNV4EfcIuYgYkCH8ybv0IjXNOzcEHIHUaAdm
/a+kmQgQWFBd8WX1R30wnbPNJWzeeSJNnF3fQLcu17XgK5KIlmWjo6dY2teLWF5L
5wXJ3ckXg6mODitt9nTK/g3FKQMdpd/m6N/lqnxxOcnXJ019JJC9vu3r3DLBYdbM
PpUx7lX1ehjTb1uRiaQuLGgY/V2SCHg5z7j6TYexwV5Rb/YuM2u8EDHIuVUC4+um
nw55TXosb/t9vTfHvMGUgUBgZ5HbfPKbZdxMGZHQoHCrTkxvGM4VhBByswyFhxCH
ditjKrZ42QA1IMzP63GDof50uB0FQyQ5QHbAt1R9gyOTClt5fzQ1ql6WqMR7k2wF
gTdSicbkBQCR8KQSuKvEpFR1L5vUdhC/lR3Gr69TMFAHwKYfTxFi90mjQ0PMWx8G
y0Mu6v9eymQQRLY/69A0GhKm8AHB8q1IRzwhhYF91foRW692JiUkJRfP5r69E3pR
bTNQ2yXsy4GqCSBoCq8Gy1ulXy14KQd8gslqiijxq9LhyiwwQb5/e11+YcNC9cqg
0hMn4lNf+xVlKVsCS1PxfcHf68VdWSjXixPgM0nlfiwCnLH7Mu1x7+lpSbxJHVi2
cuh7ztGQ2FY+OHWMhrZaHu1qYM2YrMv2G5GCARHqItrrOtV/7314M574sVKjx3v4
fgILIKRQ7QyHy4RttknDcCRSenugitPX8OjCW6xn51btmQZmGGdyv99dOGAw6OTx
BYif7FYKY74gD3u/gtzdz1WnDtsJ8Dw+dpXofbt7EbOTnH0r/4VZWQLAZMyWD4Yv
a1sX4xoUmq9xsi9kKa5Bgf1OmNhoekgiG3R4M3rdCYTDigDBrhMeXHI2adHtV3kT
wJQZTsOEFk49OUpQBFrYUYSZ4tjM3/WgK2GvpbI2iCdVpq1NS36+uNx8SOF4QXuo
q1a6Edd+1FbXHGWaIzWBHWCaweTCte3eRWvZCQkxhnwTHgNPfucbNloDi6GVR7io
jh5vZIG8voXt7NlLQCt08coiuQg2k4QuHDjuI8i4CRxcwdPSwVRBbSmQceuvqetR
ColpXugniMnCG+IwMo4jJJfSlWtVr0AFlmWy3nuJa5bIfQ1tb/6H0URo3zC6H5se
QGieAngquDBvkXObe9ENbSqaA7T8os3pHjHEYsxF1NOVy2xYIiqopIIq9MIkP0/b
kzcWQHTZqjb4z32PPVtQWnjRbvKvOoeV2D+rkZL65snn8Q8Y/ASOFSy3lC1ehw0d
+UmhDSqX2LpEuq4oJ6SR75wabyPr+MENhJBn/xPrnWAN4zBu3ni9jNQ/vCcUg+52
KgGZYHwX+cU60uRlaOWPA10eYjXyzSe1U5jTcQptWgQg567/LPy9Njf2KNDzzqNG
uZKCoHIo5GSqF+VnLXYAxlQK5oKPszF85RGNeK/yesQZG+N8MHdOm695GB7GtrUB
3MJUXyrMKAmlnoOU3SnrNORQAdBXGlinmsXlQajd/xMz481F/CgQIQ3lCKxVc7l/
ubOIreLjDJHwZUe5dcPACfuChskaDGGdU0Wqv7e8pyAkVjDmr9aQ+WJzSUx41PU1
U3KtAjo9E01D5EsoyMNIfYRknXQpzMUWWVQPY8iSBNxCIm/gI4TIyJ+uX4x39r8s
kcsaiK6aSLWp2pkGuYg00lXbrM2AtE3e1yMZgEjJMHE3uIxMipuglCLuy2u+LgBU
5nci1W4132fwoVEkJgTUrvSADV2VbipTXHPoaUQlLzSQT3RoPsudInhpl6AKdzwN
hwJlqy4lS+eiFHc0qWmpdx2y8lvjlVB3znw4phJ+TtNu5m4KijQRFOivu9mf5ftK
bhRVOpSQsOLPK6gdXGbYJKut2FUrIyFrsGIwvB0FTnZPYgsJsBFpE9m2ZotgGBjS
6HTnmUqf7LfkUu9hpboYRfc8/wASGs/pb5eiGWQJszXg2RFBHnOhzHHf64CnBd8B
BCeKMVt4dlcbVKp0V5Dpw57YWtZwJaWgttxdhCEYCJr5drpoTRLBJ1lH/+q5vz8g
aJm1V9Fsajg6+5Cwr7i5CzrM+pxd3yzk0pceZ1YHwjB9i4tvhz80noQJZ7J93sXw
w2jB2PA/DfSF18hb4s0DRkonUrEYF9DMjCt8t1Bt9BWwKD1ErFRQT6hPVj11Wfgk
3cSaUhyQD2EbxahxYeGEtWvAb9lmwpeWvWcN6OQzLKccLf07k0qLtul22LTVqIJX
/4F6WRFxrgizZ471hQvlO9+BDJOHUSdLWe4IXJgi1SBfRj2KtXFcP7CAhGhWTnU9
8Yvq1dTUHe+VZj6gfR7ZJcUBQ7B+1GAniEdfiEErYNVhQloyQunnsb2nqCl3Eqs4
WXgY8KCwOmmBW3QZgvenzkgOnxBtOR5sGvoC2YNg4qQaCcXV0Yu2MIq7rjxMV6DN
d4CMvm8/CJ7F9cxrNvsuZc9y3by5v7kiX1bHh5UCRqi4bmPC9tkhAkPjnNKqJgE9
ngU3jqplHWvshz+ehK8CbNxRZuLorgqaBEE7LBCF9ZCEp4sLW09OAbcdqJwEr/dg
6SDLS+lUxCd8SHyFNLhEu9wfbQFFDtkqGkuwImqqtdv0mULYGpoS+jiTuUMFYc4N
hRsFzBBNwyy4rCd5levwBamu+IixTb/bNFHaf6ka+HpNyWI9rz6c3l+xXtrf6tdT
BenPizkCNMjGlA7Irer9IxraQCLCRW5jhr6+k/Rmv+cOy//OgOjopPn6Y/GedADm
msXhoITo4f4FGEMysMuzuas/Kru1fDAswPKEry7NS2vCr6n+Js1WK9dJfoQuIx1g
3BTWFcxDyBok+xmZt7fNOYmUVANUSnotwUXe6tToJWD3xUVRFxmMFyruhsL3+akH
kRS08C5ePzWyIdCJMmTzCHeqX3Ru/dMepMuErqM6Nd4Xa+YuvCogaheFMW8GIds2
zZpuYZCqh8/LFFajb/qP/Q/EwtKy/8pJYa1MSRcty84/T9jdf1qKcIVe0X4HS++O
3vHIgpjV4DGhU08ERE1MxSAG03/D7cFmkpd1WnVVSAAd0mng5fdEBQ624ot+IXeK
Ch+KuOr+Gz0iYNICmmPX7NnEA1/ELHXkE+19/V2SVVOVPsen0uW6jP1LTVP/ll4N
9SmTEhdaHh/58ibDRHY4rzFAk3HD8G+y+4jAAZs5KKmmqjXmzBfiXepzlY6hRqmB
L58BVL2sZy+6v7GXhux0r+brGBVnc6hjXsRXBTTxZRr38hyd44Bk/RR5JeF5krHA
ZxtNQOnIh4eiCC0pUMM0r8FwIoJmUUTRsBsPDT5yDV5RSlWsyykr3CS7PBFSjjL2
F6vZi8Go0Fztokyz9cDEohT0Ekfl8Mi80ujd8qvGkVyPOKAckyjIHGO+2DzQ4UsF
QtQKhcKXezvA5cFVbwppQaXau2Ra31pqhFGUArznxs9YSbShw/GZDV7sA7CyHGaM
tIcjpF21I9ofzEmpf9Qk3fjIDdMgPCCmapmn6ZI+MSEca3sRfXDTMXaq1HBPOEgd
R0c3/Q1Dd0ujue/Qi0qGFYNRRgNO1ZXkMHPZeHsl3IJjTf78sD4GVaUd6ZITPMWz
pHwMZm8dvv47vB8cBxuIZoN1SzUcRBpi5ecrem7qyYBFQljatoCKO+JtToF0KxO3
2nMO6DKoAKu5GNyl16AgKqOxs4C1UR8+pI/n6x9t6qK41xleBnY3EWhGG3ki/mlr
p3rJwB0nNyq0WFw2VRlS9egrkirIFQ7BCfwQJfcHuHsTdSxGVwoxOhJc5LxPt79J
Ad5vU31/WWlB6awBNgXFphdw4D1c/F37lSX6KjsERISbNLSkLWn+jKKArzKP3pfR
2td5JY/N/1ar2kNt6yDTeM54wXb990SxjkqYcKiDi78ZcBNDxN3bVMLZsaMOxbVE
JtyESaFJ/gpkdqgytoyJzo+G/q/t2tEApowRAh5xUlQEHwUhPcz/1g2DlXWTvQ6a
IYvV0YBuXDFqPsaWDfBTdhZHF1GGHnFMuiI5jTov27lx2OGiVWChXPEBig8VZvJx
/IB/D8hECJxi3KCECcIc1kR9LHO+isvxtekfH7Es5y2yqLN9xip8yHkbw4/cO/MZ
BKfmTGuJr7MHek0wrgPdZc7ryC5KiPQEYZxnk2iPQj4GWcl7k0b9DNb3JkG6qPTO
Vp9ex+q+B635NI3EiwfLG/chuZwgiZcme6fOvVrlrJIfqyZUbSZH2+SEhPCUnnKf
e18WObGMjqATk1deW04Zv+YNxRli7Pp2erkJnvUPebZQQnHZ0CHJ0TE8tFaUlzk9
m1qJtF8x1Y4Awwrlv3iXEt4JAxbkI2LNXzNCq2v8dBiK7RaxfmRW2Yo7Xy6ub8Pq
gZ/K/l3RcGpp/Rd4UdjcUaCc0O4dxyXUDapWTPmU5HDhjL8wbGO85rH1cOhHt1RC
iI8F9jDOjicFC38MCBjcsnEhTAIjimFjlXZo+GTHKjrShaMquhCWs38e34Zn3FX+
AR6KwY0lQ6aST9m1tgBKd06ivkz1k8Q3/5FgITZLn6CiWXmEVn0mYu+b1d0yH24S
kvbTefJpHOd/UH1W7aBibBA+OI6t+nhkjrHwu6B6Gd1XJ0dgQ3WsuyVky5xqNiVA
N4d5gNq0bl/8OPOqCWYdKT64xlQt7jukYRjuVsPsz/DJrM5cRZViHjUvUev9hJda
dYNwNN5KU63AkFHOAjw/K9APkeZ+FYnw14GDzD8Uz5fl2HCYpLjkf1YYP6P9vECI
Buc4vUlUhRO+a5Di+bldkflQNAaRXoUNTbBB6u3ef/Q/r2j9vHEZeX1vQ0mfCe6n
Lp/1JKXoGLC0YO1b1Qn+jN+yIIJd9Bzo3pyILDwAt8Ov68ehFlNTee6cC3ZIAb4G
No9RJItmYFo6vECetuEo+Kp/4rMdfbkuKwyJ0PVkHaA88ZHopmjc7eJqpT6QveP6
r67zVfiAy5rji6t9BBuAFGhnyEDMss3UBEw8dXrLtjaeF21f1lfs9/FotLrFb/cL
SaP3mkynh/qIKzjR+js96mNsEMcqfZlUn46isvPNW85WkJQu9wJ/2UHq8zo7GWF7
Pma35gEBBhUfJthX0zkk5dXzEvOXawIUaI342L/fBnZnBeEcztkIoaxk1s/rnuVW
IDf4OuT1JtlZWUuDibV32lkrG0CAO1JLX3BfhnPFguVr7hPyqi08kl63Yud7yga4
nhmUnf4jB2nvqp3x7XuEZJhJU0TOy7g7LM4om3mypB5Tt6DPcIDmJP8UR2JxiQjz
/i0PyctGd69WfJex/FPJP0vQx8XtjI9nE80gL2IJlHVSy35QXedC2U+VrN1RrdTh
Dgw+Iu4lXdhBLiE3EUOxxx4sP/gAY7hymTTJt0nj1jMagxbZr5/1flYCmK0StGrC
3DOwRaBRN5449GhrNI6PtY9a6dTCzRvk8LYzCmFSmh0rELilvteIJ415doLQAqo/
KES5vE5iJD5wK+N1UNr5kX4xi3cwqPsebo/muU1QhFg5XeK4aDi+YhRi3ffrwjus
M9KHfsUjvlfV2WPGRwINhTKUvSZ2PX43OnssttYZAunEguCAhzFHtQ6k44LpIF5G
Xhx2V8JLlzJoqZlWlbChHeYueLDQN+WvbCaVp/E/v/a5k2sCzY0zvvKPkmfq0/rH
KwwFPycdjP77BI2TEZM0UiydWMpW/H9eH0Y9f3hbsxS84KF+zxWX41spWUre8mga
b/szf1Ghcm+g+yA5H1vXzmzrkU2rWMn/6f8cgoGSnLY2VSi/uH85ngKVxuL8tApT
N73D9yDnYjiEgHVUH7zSM4c2gsH7CXZcJvx775Zm84vSDpR5NrqbS6ZgYntSZdUd
t7OO/RB53h82JJfEx4DN+U3Sq4HGaiJiKr5F6hJRZxCJbz6GhxQ5CwZ2BxX6I6Di
rjVvkniSgZhZDyaNsBlpYanDMQUOOYazY+AFydREF0HmXFfl9VJI7xGqP/vrvUql
brvG1QHYw40CjKaz1gJM30m2HSL5Xswt4iPDFuQzgkoIEUEjFR6iFcHJAgoplaRr
6hnFzbV6Seti6alIa5xic0jC2kZQcEr36/BvTMyyXrQB+ufdzr+dmMfNpWlfSZ/c
AmbtaNnth6GVtGtZQ6OIzrOWaO5KRJIOhYukEc6k2FNDY/OcrVzGLdoOsHiuDl2c
fXiK01iOZZJos/0tZILvyMHrbI7TzowNE81JA0abA16aT2vzrDsGNzr2+iNUWTrJ
A6SKXxl5mZaaJBoc27oxU1YWBLdaQYb6+riuOWaCyWPJALF255S39/SStG/gqkmV
Xb1A/PxYdsp5rQziY+Tjf0AsC45ciKiM2F0dQmP4cGYOJgDdE1vMya3RCSLkPNdK
DOtyVFcam1Ki4sFlC1cKRdcnflTYEEACRwW3suyvZDGmIf/29iCExWmnZLg3OxXQ
YsmYhduur9FeoYUeTdRD249VzF1QvZtWAnPcUNrqkNaASaSd5hmmpI1gLl4K5PxY
d69noQ0irSzJauEcTng5jd+/h94qEa9+O6OY9+ceJI50Enz+GLhv4aDqjYfmqgHq
azRIwPch1GWurf+vOJEgs161UUdLpXZz5+iVLjO4rn8HbGI9pAgpKq/jC/FV7aKX
Fb2raQ459Y7oP9rGIvi+JcMAKsBkryC60ScXv06s+KL98jjnrTaF/ggw5lgJjN8o
sPWUqs8ML1BvpV3+Q6wqNkajrfEpespJz4jc8TxnZq87ig58U5bLQvd9RBOnEZeP
rgMkKjCkefEyEUgfMvR8bX/fYRn1qONOU5WyC2qH1WD+hFAl8uM0a8RZqUZiF2/5
wvKIGGLFZxxl0FWQdmvLG8+QHzqHgbwx22ctuvkjRJ60jp3xOK0AuMb8Z6K8gWpw
xpO0PUU7l4/TzVftprV84/EbMlnY2nTdvLBqxli16KSvACVyWLyeykVakja6s+Ye
100t0ZFTf/m2agAdP5hf3B6swytVQhZux/S7hZlINXljl/I10BSG60UOR0QSE4x2
IUi1Fpd0osWmdOeJf4i3es1CPgwGuR6TqAq08cw+o316Jk0Vvgrd/a7ZtVLELssP
QDlc3kY5RhOWWnW+DZlU+XZYpc46D4uV63ocUeCVRh768C/ZezTIn9YZQ0Ht0pT8
UcLHGm/5jMgS30jUsr7HsiPSLEByGbRjqtFZhHWvs6kFWVZBVHCdV0FZRD7ybYAx
HmpCgEH1BtIoiuewdZ6TxuWFqyqGHv9mx5fWM6heU/MyUuE18akmN8DOMJci8pP0
z9T3Ce3Nt4aoQaK/QByAdQN0QrulgcdMkGUNqv14z6SWO8CtR8lWftUZPFTMpfE3
Ho+lm9q2Jav4UaTCSJD3mzT9KJj9IApRYFzN0CooCVsW9XqSBP8DtbpFdpK5Oeqp
NqsLn1TQTqRKEzij3SDxhcuj0+5FqpiYrN482tiy3scrxpqmID7ribNTCKxMBXEP
pl5MoC1zntLzoje/ScFf9ahr+J/HYXyerY9JjF0qOEgklM2H/Lz+aADRNxHoj0yA
MAOBqOcbnjgBPapXYFQNfLUhr8/7Vnx8I173HGLgngOIc3Hx2Zv9+HbdCdaKYIFw
B9+HmBiukvS/0wHf+a79zENt5GjNwPOU25hhTg0mWIrhV4S7Xxcd6uaTrJkqYfa9
EmszDa6B+8U220A05ouMNf+LtvK3nZmGrMpUL1xfzgF8QobmzBwtQSgyKnncbQtp
GeqnIsRAwySnAf61oeiZrcxCnHh1EvsK+iK12xbnQ+ZZw+6vq5kuc/6QMeWmev3j
pV5ZTsslyijrMUWDfzMQbBJAgxzfIvJAXWNzeaj3onY5P0DTU7Kc2JME8oI0yzTl
Nn4ElAoJIyz79FYCbqtsTGVNPaztB57R2CTbxQHMGnlDnaEoM3hB629P5oyQcZHj
ToDiBW9dghcxdQRUc3pXtoZ1duKrnlY4sbouY4+L5iHaFakvuJ97GxyZ/jk4QKTe
HnEUxhsLj4AqeUSxpUoFnqrAS6I0WW4QTtJi57ZBUbYdB38Le8lw44J9fOcxpn80
wAsayAuWgCdq0xI3/pPEuqMLZebCzKDzCXWfLc2Kqod4lDhEq4pAr6LEifLSg0Um
BtBVH7Hw3oWjkHBXWHygiKpk+TWYN45hmQTsDmmEmT+AUBr8+zy89hqUoLLxC9FR
kbnO2lbPKV5ox50UDPb8m1HM4KhdpjUwmFyXLgbbU5EJvjJ3HvS9yfUpJm7Fkt9b
yAIa7jeHcc9dYHcZ4kCVTy1nJwU/gt2eN2L3wSmoq/giVsXeCm2FQwCu56kO88Ns
XNdLFVDGSdtRDSy14NN2fbGKizi/pof/T5cdCc6L0RqVP2vJ6XzTjJljmwqTJDIU
N5xDoNjbmLeP7zhOxWzN5j9niXNmHkmLzFyqMRDRVXuoDUPnkRlYG74tMIU0EB7e
ob09CJe4/2DGxxQLPWHrIBTozpYy5K8PpaN8umoqzoYqw4L/kZRYh/+myaihHI1n
usCr4xCOiJXmhJZVl9wl7/jO5khzl2tVMwt/TuLkTXQ6j0k6Xq4X57cQ1uUBRthd
gdkxkEo9L6z2NYttlNreNVf38+zSBaeLZ3mbUX07iQwxum2kI0EwFpnfjntCuJbn
4o8Izx+qI2sog5oLpcSzjRJfebOypjKViydDZnuoPweYI4ccucI+V/c9sUFlKCRs
SFQZsmWrYJEkEOQvydFZc8Qi0jHiPZoJAx6+REmHvM4+mEtCNvEiGQMFodGHfwcU
0ShGyJBxp8067Ty3swv4YMSsVn4mucCsHaHFHqUoNvdcEYluOj2Jt4+vdGS16HjL
CbnBAevp+p935IKVCP9yOhP+kJ7zpxgEO4qt5yByNu1xQ0Ci+CuTsPHk7BN0l1eB
/S3JRwGyKEicj0zNClH6xQI5l+iqwbtbp6i7C3V6PCaKViLFjrtERlBUdE5argoi
I7IvFl5M1bdn8imeDXPU5aRkFuyKgIT9XvzXZQ5ElxTaYU3FphJlD/57bSNov/Dk
sy9xCJfuPXGmcEE47uFySNPkMLXzBJd7qPsK7y/3WFrQ0TJQRCCG3FcGMKaC5Cff
dqptU/gcxMdeZO5R+ICOSz9/298b+75pvhjX3iYpAn0+WxspyPEdr6WW8CxIz99j
TJTsB1ox83MLTk2myfjtx/RWqQJABW1sVdySwx7J3JYrvMAEK7iFBxP+h1TxriU4
DBMBLGqhN/Uwgj5wvMfjJKURdhl52WBTKCAQXy199psUBR0XmJst7YkBpeceCEXb
0/DQrrBG+PMzlr9k+iNXy41DkvKKzpHzpTmQXbjUgGbiERNrJ9j++VFzr5i9k9+K
1OTF4Y0ghAkMUzX/oCzn0H/GRmSasEUtL3Yh+PwafPQgKB+4SXm2yzQTMaKgtoTj
JkavCO3xLM/i9yYg3GDjrRImOARN/MnTprvZsgLTich3sfiT5tlC8EMCt/CNZeBX
3yR+7Fs/mp42TPH9cTpJDA/airod8O1sOkV8UTxqBJbASCz8qkdEi6hcBoigobc2
by6uvsROLFZFBaD0C7za4c+lvXoCHFZk0IdE4LhM5IFzGSypCB1aFYHW8BW9SOpx
RXv2nIChSFl1xaki8GTvE3r36q+yyV2byXlAvJryyymz6JZV3G/TdAxXQCzzo8/O
v1IEM4h3PLh9IkYoTs2hWnuM2FDWi+qAKX8O++VNK/emz2VZiNVsf10T6X821+Q2
AB+xRQkcg/GJ3b2ze2DqLPswmmSF8KQCRIb5hNy4niBWb+KUNOYG4F7dHIehf56p
sVs0VIqcWOCfsJ5FnXVzAXlEo/zWRhXtWXjh16EbGoTqvcvM04W+kHjOtrcO4TwV
zSqCIcbByWK9U2K9aJuchMkPc4pNPsUxdPre4W+wbs7gscHcrTSmIDzx+gNdG++X
t0kfE52Mge7f+GIiGMda7uyOsHriR9SNZkQ5gBHAdGyL1Akdpl24WxsFMM6xa2Er
pLy3mbjp6bWLoSC3JmAZUYkoRP/XHsvtwy8wu75x1ac6OhtxTuK7yI+W6nFBWZMP
V+EEixGcuQePriOFasltipjynWvb4IUuhdEsMRjILhUx86xA01aH+Xnvx6/8/uBP
jBh3wjLZMAEvDMQI4FYOLtClcsshbYrN83kpgjG2jUIAJrNMNsayvk5IgsvMAgPh
/taYt387q/bLKEkQ8yruovb6lmFfd5BrH3ftdJV4k8g1PFvO8Io3LXxgfO3MmMz8
n//Kow2QDVnm+wOsYtipSrWUWtdFjET1o/yCnfwDgINRTV/QXXO10e/50x/LMOBi
Jk2Acw9Lj7sTKcb9LE3evBnK2ntxaCzAzYSANbk3A1V6cYI3J/Li8dQd2xRT81z/
PcQf5b9CIJdkQy6HIAaV3ezq7PIN5dXvpg5GXoWwS5CCRA7q9jvFvG3O0tzr+9h0
tHUo0x2v1dCGj5YJT47YYmR0zCilf9aWyr1fQDsVcc6YneBXK19sYEMU5scycRKK
UIoDgVfeSFBjPyO8BYJCQLSmqK+iHN4MAkAa66VjHQ5uLCIkG4tOWE6QaHbufXi8
fzFQLOw9f+qgc50VqL07Cfsbe2ME0JdDDVVJG8II7JdDt20rEXGJIsIRNtu4qOVJ
gNQui76Ra/q+izBYgxXobtcagAPb6qL/Fl77S/6fnYzKIzpzhd6oPDEMY59N0FZ/
jvWlqZaMriXwiTU/Nr42DFcudrELq6KMJgWeuIMfObQlRRZr/TgB04XUrCciKJqc
vrsL6m65etTIG3ptxfRUwOMEosKg644B1AxaJw+5WmLIrD8nADa+rdvufe0SAHnf
mQzpooaHwsN7AXYSP2tSUq23wW+Katk/dmW+Qy19lcnBzk/BfKi0BRMbEWxdowxt
ddYSwa7tvP9gIE1FCI5FtbVVEsjRHAxW3bLtlS6ztPCJ6L3dTk4Xsyoc6dINeTjw
wwFG8RQGsmYjYlerikFGWB0jrRy6kEZCirHiiqvUbaTyDF1gPG4kaEL48om/Yr6J
ZzrfCLGYy3YWSvWV5acNa9oInZTmhfFH3vSYNdgyuAvsRUuIpcxOCmKhAO+Y2FTN
KFvBp0/1/G3rBk+un3GWkMInLdIZPWggkcBCSe5PM2YiCPVIrSNMo9hlfr6JjZj9
p6Lbblz0Wc9TBzTT8EQYv9jkg+t1lOUpih85XOlFVRZtPIQGNURe9uyuGZgZOAf8
H9H26q4LgtuG8NEzeWmNpFYwR39DGrxQshVuW6GEBG5crBAY+kkflQ95bhipmumQ
UAXkRuC3iMG7BicTryHHZCgUDUrzxX2cC3heBzPL/pAj6+xql+1a5WDMsP0pqrnS
30KMy8hckMKKf0r0z36O69AyH6Ycsv3c+XhgKoVJXB9WSEU0GGF3otgumJg5hGh4
EQ+bpkjgx1kom6izQ/RLqlOEH6fobpj6dHyEt2e0Ev9YSc8hITzS7cqox7c6vWt2
/ZcYZ0n1oxFx+/Dq2aZSm/SkxMwDHSoGrxxGSq/MBhjoSOpvSBHEm1Fs00tQ/ri2
I+yssgoOhGDMs9q2vYATVNgWWKPnz9ZQKgNM0h97YSSdojIriIAVQ9LUmHAdx9LL
pcqKMoPfpIgfGF6tJf/d5+K5mu9YdTcQyg9383S7Doe9K2t08pUcnoXd1XuRQVcN
ntWe9rCUQ2kj5bSFcotb1o925yWCUmMu6JySQve4vOzP8rPLDwtkkCAioqJIESKj
n1tE94VZrqxqdZtnIJE8cmto53Il2ICh5jMePzL2ExlpdNIieeDy4FJOpuBLxgCE
+BdFtfmsHNlTWKDOd7suCs5mrWF8R2OVddPp21nLQ8jqLwWYONMOBdj5IW0wsefE
FsCCvuZiG3r/ViXHJDPqGX873Hv+1y1Zkt6LZj0V0Dm5CCtwR6hfXWmYMNCx9xsp
HRkSvvK5LoPPH6tOyhXwI3JIoGVipr7qLCvySEGk9molqTOwQGqTNtRVvx8N45Bf
o6lskU//q06W8v/49654OaXPBUcniwgdqE936CNvi3rON6rvwExnOiuuDa5yHK5f
16YWJR2UUIE5VB6/ZgtgUE6dNX2yKMVlo24s15TbRY0fOylTmzn4DD9tG9IKrlwm
POARmzkCK79pa9GATynWnuafuD8BjAf9onPYenUw9Dzemc719kw1B2IuDg8XHEBo
nqkZ5sMHWxFVcNTORBq9j0efOhc2lm3tG+ZEuTyWaEUJU6dO5C+nPKe4RM72vk2q
f9dJ1YCDG8Timpwu8ghqYuWN+YBFdGRzsaweEMoEr0DKXHGLGR9E+8tEY3RKdznW
jQ/9zBYe0uaeuXmfSxxTosDdo3HFlf02vX2ScgT/fMAwRcuvWNMgjU2Puvv9HNI5
eSG57pAgGeraZKs3WOPGKBlGZmMxyhz5XAVRHKDOPxYnGiGZuC/gV43hesWtAjxt
j8oQKBgdBdri+F/dm1y8moMkPY5zE9s0zpSaPCpSM6lJAyi8iLcNphRoTIWKGuup
g2hPpOa/7RVedGjXlm2DuudSMN7yO5sIa3NCG8jFkocMoJQWZoIQNEWrnh9Vas6N
6IhC86/3M2p0k4UYIzpzTWdlNq9ZoAXbQmtI1DHwhkZl3UD0hTbZEToRdJGY4bum
1EWGIWu36NTcLkydOJ5//7Tem9iYSdr48YD0+kN+Eeu7JQdqIqiYw7TjJLBZqBXD
nOD9zyEKCYvxeQYJtzD/HIPiaugbUjAWopv+8k1XZz02tvUrcMTOBkKbjG/YPvqd
DDrTYpuIXWrPoWNBvbXy0UJSgTbxn5cmWehzJ6vJ5ZqP3gtqBgmUCLadKiZvWUSJ
/KTmOFGcimRnhoMA9gc36befKJatRiqtfXuO//k76X87sGAETK0g6VheWp1YqY5C
Hp0fm5/gO2/clX05GXDmoAc3xWDAa6dkc1g80P5KxomH5uaDIrgkCPoSPX/iNtsO
yJifXotEnZaYzQBpuT3JNzDpK3MTmLpafTIEItoen81tCpsAxD0hD2oCVpOxpOny
TUCrPihYz6a5R4ja3rAn5PZovMPJvX+WWQvwQJrbol9ql6Obo0tod/KLCcXxX0XK
5DmRcuUKCoLbveJ8Ffvc6J5keTRsFBWOH1+oCKkL8aZPMMNuU+lRu1YtJb8SRaZm
WHdflnL8+i9KBluvTO+QX2Rx9JyH1fljsFEZW50LD8FKm4tXiZR/sQV4v5l1L30t
UzBPRlGblKyXmGhgjSfGATZ0JWZh6rmpt+kOTKAeSfSTWzA/yq2D5SZez7IyMBXD
adX9rSUGXMcYhCHESlrJAvkoMpmFfVD3IzV5ELriWhFD6Rx/uT9l/yWYhzQui9TP
Sv2idXCsQwf1gTDbDRA1bMCEiNaQEFhy1Twb5MzNLToBviKxSwuT9DiH1gr7QgB4
X69UJvJAR6isUQmuN/ocsz9erMDzWORvWDDQhqFE4G0ulsLlLdn4VuVLYmCH6Tdy
eGT2kOd1ZH1jl/9rop2YNeoeZQd8k74qqP1oTrfCifz8vn6dLCOeNcUZWEFBbVKE
KqrXnObmrHoYUSUD+pY9+82zrcsV9YcuvsTCAy1dnOxJrAGuzI9t3NBYaC3C1kZv
cg7hpbHRut3QTVXxwKi4XvIZt6H1hHS6z88FnlGsfdcdeziiVjQF2a0KdPHzkkHY
6fHESEo+NAf0B7oHvm1hPqfNYL8+Yxmk6cvL9eX4AoKAPj7Wihz+D+LlXxVkasQp
e2tkU+FINyU31QV8h+5TUXNLJSc2V3VyC6HmzP06mLMn4i4V+InwMrxmCKaSlYTI
nmya3sMKFJu2vMlzbp5Ik7rBIJpjvLFsmr0HjXZKiy6p30ZPILrDLrV0T5oa1fGv
y078H+3N5E2stTT1LFUocbUI+mM1sl8tFb31ZNuLldDx1HI5KMPmDrKFjSSV8jc1
USYRSLx+xELOKQ1AMmz762RpCD8qcnspo/UWEHoqYJ9nlgCdUdCs9+b1y6qBNJhs
cRNHkjY52mkEFFLLEvqnAtuJSl2HTmDHRPeJS2hiDjiJ4560dXJIxApjxqOUcaT5
ObkdhSYVMI3I33kw9s/4UW+z2b5bpaDre5cCQihcWtBEweEdKwzPE/PG1iRSsoZq
HwzEriCLJtwhOvHH3e1ub2+SxN1CeNEVfSufmjbEGmbo5SSaFgkzvqBSyyaHlDob
q9tQ9mxTIYtUn6gk3HXJGKzhhAKflUo5A+Rw3/ZUlmJstWgta7at1c7XQV0Vev84
E4SAEK3iwW9AyaE44wkqdRiXPE4myha2jVDGPGgBlcN1c4AFb23dHbky+ynqH5+l
wdRIl0rpaU0B+iRIpy1+qKw25giQy5/SmONxRWs3HNV3tihIo7b28/FYZT8us0CM
PGA8mUlNSVAEq1xjQWVpwbSKxHOgXL456F3t+P15zfAp+P4qUUQ0RRlb6HDkynct
HM6JevInZPsPQ+rfeVRgqge2GVyrmvONqy1rL7QjaK6xbJHmQTvyIRty6nuy2Bx/
4i7koUDvxYn0IfZAbIrg9inDeE+BCn8ZKlljvJ2K7BePMQrACreH5G+WWVQdkZaA
9CPOr+yqvnyDXoILbg0YDfO1ksQmQte/OI0MPjaB6LXhVUSBT8bF+/SpZoURCQmC
lUlGMsqPTK0DYQA4V4PjyMk8YdSNmj+zufEEY336NA5gS5Sv3O2Upp1GmkB4ljdC
AAYRdUHvbEnIlnowWJoT2FD0Jk5O8uY4V3NZcsoiG+Io9YbZx3GspX6GoBsME4OT
780vmKksHeFgmUzSAJAIS0j5f+/Ay/Y0THlGr4gtjlVTfFYSjXjZfgb3XVqYfp+D
DQv3+C1jCThyhC/Sx+UEkefLrM09eWjOtxrSur2aQYpHaV0DI7guUohlSvkisS6j
hnoNfPqZdR0DEGC3OHy0hVLDkvfrJ8AUSMSneeYaN3YaWSqQOP8vHIcNSBRudSIa
JsyMmBGaOkgPJ0eoaLpYl2YUp4rOirMD0FlR2pK4bt/S2lW2E3bZy6cw/9ZMVUtV
dXYkPZGyy5O5I7HzUP8vKKsrdyWQa7jDAK9MH7MqskbtPjDrR9jms1VksznXRjC0
vsWr76Uut5geedmxZST8i3tuiluzhFkagn1KjlhdblqdWjB62qv1c3wRJVAJ1GON
tdNmXqi5yixjqjYVIje/aeX7OhJAB4bT5EeuIj72zGWs9QFoG2eS9D8U2boh1q4t
fZthReafMgLQsU2nPIzj0GzZo8Mi9/dpnpNlq0tAd23qvjdgrDLnWOrxYp3SBatz
tM33v4gybuB75detBrBdaRRxze2qeuDkQzjIXr2fRqTudOD4OnvT47ZGPxI7MEz1
L1bohvDpoKnvi72AWSj3cVJ8ppxGjU4QQb2noJKFPoQ/GEoYKD2/eAJ7j6/xGYek
hVM0BgK2g//Fj9E4OaYinfFdDME2RIRcn+CgTKzxVUYebDxSW3MllEqgfP7JlAwe
qOpIJnG2Euaaj/yvzeDaz2oAPU4eN6xBkdKRqbByZEaAyTsQP9s15rfZa76zx0ro
0/ntKoDPVWEzNn2n6+wn1PKML1Z5jh1ngLdAKjlTxNwpzTtP/+4iVORmzwh9vwEA
9QCZQqlsUxmpo+Xs7VMr6B4lCnIc9GnZjShDtocSP2ABw52+QyEvtrNM64DPNStJ
s987ygQewQcw0KwNErxtSu9qnvXo7J9tFgJIiwMzwF4FX6K/vsTipjIMZN0WQD4u
y8u5iOjXwHpr/eSeAU6qSvXV6moGdzl3cPQewXiQTXR8c+IjmcQhFygk2Zwr1+mv
nImTWIRs32pLJU/VDa7wpYjzc6bGiZfdnNZYn9fcn9DXY0m1l8he6p58hKxhfv5i
e0wM5KQl6tAnCv9kpFymxDBqsXJM4TV39bCUjg6B0YIepIK8gyqaDcMlXqxx03Rq
lCaZnBE7kad0e5UWsGkUJZeDNsN+J5keoHJuvXnbl6cWQ/PyTMdkhFLMZ3sHnP8U
hffkGulaXOSp4Mo2wn3YGa2pV6d55IH3X4jy5/bvxRBUnyg9S9UndVOPb1LkKiNK
zi6o6MEqG+4Txz/ORTVZYeCdfxvhxNEn624yJH1kfZcO17aJYjv8Q4s3G8RY7tLz
ZjO7joxNWIF8awxVznY3X+EEjrM+YLpIhBVqNosjEFdNuK4/U/NcK1s79a/Us9MZ
w7czlZ2ad7hWkKZqX9RD5fdNsBjT/ZslhHO5Oadoi1s08yI8Vz+VmNLCNXkUsk5Z
iDzZ8KrmlcN50BpDUylS3gRy1ivwnO7OiUN2tHM5ePWdLOruc6LDSQp64J2e/w/C
tTiKZrrO2S01hwOJ5/Qi5uLV9Da6RnRKybHty1TfAkg8n75ufPkt7+lU5SWZBQrl
SgyPnu7pQnNN/VCJu5ygFVGhFasmh5Hv3Bj5WzAgfrot9OORdBV1NUHKlb6r6ZzA
uwTR8xmXWGpNon++MLpAkqSVGnULnlvAJD5nHQ5xPyKW1TABxUJ/8vxNT9IFtkU4
2xZh2ZA6tY1AEObx+jjvQVp6Lvn1kmEj30DPIMmEvxiy2MSrwjK0jPv9YAhEnAvx
NejVqxGkcjDnhG/cOBBhu0oWdRXJNYJNHXifbzIWggnA1T+8dgJfwI1FfJViyDls
nSnPB4V7fQ0CYFQlT7VzXpNezkR4WeazQO1SL1mxTDT76zVcQdnBT7ivKQrBsAva
fypeVAT/HZiOzEr6+ohr3q3WFpY5cEEGDPPUFZzTH0Cm5fq0r2Q3R87Y4LCnAlNo
TuK7aVetyYxiJEV5NJeMurKSYBBi1Tk1lY8RzYfM1Cs2GMkCx5eGQqIm6m5YQYac
Pv7v3peg+dq/KfagOlJTeEKDRy0CBBegY8/uN1tYZaD2s7tEKrVGJir60C9FBSm3
cgt+nXXtt0FB3mjz098bYpmdKXp+aDTQckL6+tgPvloR07H73Yhhqc01LtoscE7z
NSZFlifm112sXKBgvcqVH8LZCHAuhMC0ileNnm8SGYEHKxetqn0IWjFZi4mrsv9G
kw361RJoDnECtNGwdTXl2vBcvs6Cq4yUsTeTvbdLsLSdb+b8HqRI2GOe8HmoC0bQ
PLypilQ6O6/awnsi1wqs4JN5pLmkYkRUKThsy3n8SZ812M+E9Mu4Ah2jFyiGyoWA
lN7s3VL4Pcc+EORofC5Cbxa1qxpQoNkX8+GFn4jCPMfydjL0ahIqesc+BjN0ansC
JoqSYs+zQvhVU/D1r5N5UpIifRKG3BtP/X6I0bypRmeRBeAVtiMoJa0NR6uP5e8A
qT0EnQSYUzdA+IeRQnbtZdPf3/3SfpmaDM8bzsTBDfeXyQKgFKmRoiYQ1YZpyX5a
yVQLI1wZuf2rfzWsxaihWO6JsQiyD38pY2lVV/PnmOQMJgPNlNolUV4yz88huQXk
vVOpy+SyCMTuIgOVYrPLULvIzcA0g9iq5PiPiSIvAQ7JqEa2U9Db2QWSFPqkupL6
UwuexTSVXEPF0jZLsyZ9zLpW+XkLQy5QlZKZzOypG4OUQOle7224AAJxgU/BexEe
N2XjEe9YdwmP0kytGxRn3JVFvf+HppMEO0IumRYx6g7iQN9LWtkb045FZlwZlbWO
+0BmyLo+l20gWEpQ0RTw9dncBnhiy2EP//cDKgJzUtrFQYnrq91lC77ww6RD3Sbi
bjnL6mqN1QkwkdYGLvmd3sUhdyXKpOrT2aM4vdjU03beWX0yeRDTAx8MrTmYgpeD
jEhHrDfAC1vtdfzgB6BPdMabnxKmqUI6P/CgQDlbVqF4lCVZojddzZp+zKZK1RCV
/Kl50Fqupj6A/JnyUmetFP5pTp9JbnrdPQAR77yfspBait94AeZ2ZvCty5isblO6
42n1TOVQJDSlI3KI2UL/0yX9fEfZQxPXkaZRk/HnlkaaqzMV3yHenTZR48XSyZkg
LdjSZ+P5f0t1sCS+ywCATETsphw8VNT78JDSW8lZtbmEQFy6xs2e6TyBAKsM65dj
DRcqP29MXwHZyMDI6cP2jPaW3ZUbPcpt2dNUVyf6CgZNBCIaI8mr2j2TWAUdWI39
RQkFN6QC7d0R/bYIU4iqzpw4bRu9u891i2eAjlYNiC8OR2Otjr74aAtUMoX6Yub+
ws5D45LXw56SDXUd9gzUjd1aGXqKyTf4Mj9IA89H07rHmZFkoj8BuRfPqKXHmphz
iSc2ieAXAc2oEaY9dv1OYfEpG0ArPR3e6EYPpA/ssTe9/g4NjIQXZURFQuO36wzn
vy8++iWK2FJ/3HDw1KT8zJ171nec43+Gul5j5Fx+zLLRV8kUxGkEUNzaByFsDDqf
xtlOE8+Tsifnv0QUH5gVObxeNUIWApJn19yvYjIjiPEhUyXGBmrU8k4LbPOyVUMe
yfHtaW2Kzw29B16yTr+jCKCzjcWKQr+a3OweRxuhKO80lftSDTJKKSk8f3yiaxn+
GqvrjtzJI4N+3j4WFAfatbSXiNO78czq36s+NLP/YK7g41736FRehz84TOBuv2W7
5hyjGaCHmQoFAKlvkokkWYixxvQAj+J+hBBYLefovMEF8msvcsl2LtM7BZh1IYrm
OW6sNeMM1ZYEs8AvABdYN383O86c7++DC7D7J1rfdUz2PcjEldOLwYQC9B/j0vzh
JLg6PiL3b58wcHlO3Gd81GTkohlM56iABEA5xI5v4IvBkhgF2pejLkCampDRKB4T
tZDvWyEGkSAP5KVczOPzZAVK67JA6OPkbb3PcpTveM3GQI9LCexWLDd+j34K+3hH
6ioM6sYYMgFuPcfF3RM03vh4EiQ6MDWm9nrw8li6bi+3iRY5hjhK28prL9LjdWhx
W1iyVEqQCPJN4iD7F0znsUJ0y3b7GyqylI2UsFuVqp6D6o88v0Wa1sKrUK5k7O22
XIpPP3E6/KagxYuBEPEltzClfxiWI9Cih9IYkJJ5wX+lB276W3mxouywbTxbZr9A
ayDSgKLTRLxWFR5f/V0e8Co+DFBfylTgxDmAIFnIx2QN3MEqftP0YANrzdAEQ7gr
P037WrQt3ZzCGbozIHzkCChcOha9/CgoODP4Ws7yQ/7rzR1ii+L88FTL7Yd84oak
FOcK8PLBVVLuII8H06JhvA3aqViK/m/SXJoSt3r0npwhebdfcKMIC2rzCvAwCWnu
7m/cFsmU3yackoH2ZS4qoR0wuuYlf/aqGAjgKt8N+1Izrv0uRCrRs3Gb+JB7MOGI
mkoeXBY8OxncLvj6D5oN2oKlfO3n+aIi00AMwB+ANoJB1ZoTCaiwolBSSdtikHsF
J9S2IopoQyPBs+9imqkM6+vfaInCxwEfSWS94ezCPTt13g3ZgzXXuKqe1GxC6M8m
d51tbl4x65TQP33/91ZZbCQNQKHIT115Lj1gT1hYp3rMFi8Q/ky5ZsD1Sl6LKy9c
Ov8mkc12mfEr8bZ77LgfrJkTmeDEEHoZRMua+V6E+iMb+B16wJOo909f+vr5RZWl
3Y3YwwSBJWIt3kCAlNiLm6sv/4/Akw8v2b+9uZNrbS3SXHhBuhJ/bjrIfBVqHCkP
gfyhGgqUAZjT/Sd+/M0hu3RnBRyKkcrlqZc/yttk2LhBo3jg3LPas8VUsZ+KS0Vu
4JnViJEknkhUGfnpmiemciGVhlGcFrZHKUy2SQOvWo7IOK5IQLwW3OvVl94Egy6U
zcFTfZ8WLy0+4JszEbhvcYAiQccDy4cTPW7Wjg9sbMEXhUxyz3D7wvjtmZV/57Bs
GvrUgsqCsBsfYAovN/pKWovuYZqdY38WDStEbbOxHqz6Q/BfK4QuVMbF3W2ePkrt
k51Wb8ktUxV8lEwvl/BPivGPT39RbrYJnYK3dtHgAeoX8QktZLsYLEJAwWTci9kZ
RJLBO91WRcc8aTcX8QqjYrXsvILVCMkl0G5MuHzbqRtYE7k4ilDNxkEHc4FMa7jO
YekBNbryLEy0QUe+MOc8YnjR/Hi4E6EKQcrSll0tQb4Gmb93En/7dIfeKKrMkHP5
DoGDqPmARMl3Mgn0N2eJX45V1bAyBq7s3ZiQZLr7ttE4RAUPxA05C7O6nkt9WESE
nQGBRLVA4VOlYJm21iNfymKwfBRuzx2evwDzrZjpC43JyRTNQqHKg0kQs2QFfPly
qLe5tYZvekEKYqi6bvrlGlNC8XGnflUf+jxtOO1iu0NB7QMDcCqKGPHvxIHt0MeY
KCs41ky/nyPZbaUccKYBMQl9Dk3U9wpHSTx9BnFiw04=
`protect END_PROTECTED
