`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DCCuCOnR+r8L11008ZUAqJdVcjaQr58CJED6M7C/TtVRuZVz65y5Y0/azkNAELwI
9yDUKsDZmWWeo09CUW5hmVZfBsqCIov8ptpkBQPbSMg/K+sW5ygXS5a7N+WBeudT
GC6DvDIy6tk/287yfzARKlOMMNR5wU+YFoBAgEWSOYT17IDp4O88PfZelVKz/+gn
cKF5uEoMMOLI6//iNhAvRFtWSWX0DJgRYH/mnQTotAef7tPHnL9v3DpWwxYX8ayD
GrxMLcg8a98M4gS+Wl9dzPUt43tk+VRJ6FKJlQQrHJA7doy+6Tyege7cCj4LdJt6
G9ebL0Uweh76YZThWxb27tNB2MKCH/lXgzzwwXcyndLndVuKN6P4VRh436UTPn5S
BnKWk8lR58uCdxz5Rs+TMd7xags2af3X5vWd0wH0LGwJvlXf5n8xaE0RylqtM0Ka
rDiJFQq7uYsfhLUKOwY6tUwoIn+fKVYM5YqyZCxD8VCPrHaL7W7lxCj3c73PUj5q
3TqE9HnzbwHKCNPahOV4hNWj+Uplh4qxvgWixM6NnTT1Jz4Ws1dnLnJ4z0NZtLLh
MqaXEa7A3mNODno3sWle+ruelAuimLEHTnSXmK1Yz1HqDpaRSW9Mx/Jiw8vuwl0U
OTi6eJKru7+0Ej3mt1yClAjRiYyrvGLWPHkR8L1Q3rWts7IaC+Uz0Oyvpl1Us87o
Ri9jrjAGbvCd8zq9z14KhcMcgWhjWdvTVWq+D4xIMCpe7d7HGRSHnx/dPAqXX9YE
ZpXn7OqjzM0YxNlto1OIXv3ZaOTdfxj/Ak27bjhddterJBlIfCyydkQC8Fbkv538
D01987B0wRmeRULT6zFbhXde55ndBACNcB/HH3Oo4L1LWDppunVx7S0KXKSsAuCP
fVMfGh/dEhBUwaVkSXN83Qs3R6406X2YWO/cpdeTmGWJavKoAowEuqIWZLCMpWsi
kR3lUFpSMbSrcnb9F4jW8yHEmqJVsJcLUToEVKI4fgBHAsMaygPwZO3ef18AKF92
Vxqh2Cu9j2eZMAQ4gsXEBrR+jWvRKENEdUbcrQ2Fvizvx4PHaGDHbbzW4uERLNOU
Y0NP662w5c4vuqbXtLiW/t9jPEs76Kihyl/UhAOuw1fjz2kcWKOxac/xGOyxwezy
S4x9irBDEqylxtiOw/xtwjmzsRK/urRqM/UucHQ7hDSJ+QIhkfn2EyFhZrdtLRbe
TryiDR/fnlZyKoHPlmqIKKLAPBG8mJhtMK4e7YR1/hC0wlIreH2BebO5YRs+c635
Jvw6UCbap39YjHbqxwcnmcuzn2cY3H99DV/98zB3UbRQuLjZX7oQZaKEmZyqJowI
Qnkk0gbzKx7GF4kdK4YhwBJBTY3QRYCVe5yHpU6oyQykmfeX7V/g46hFACyOEC2W
`protect END_PROTECTED
