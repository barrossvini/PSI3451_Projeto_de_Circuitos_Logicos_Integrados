`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ILWXh8jmjgZxGYGg/wDxdrCW4QcBvFTVcpaRh6HzW6CI5/cbaecf40EsrvgMnJh
beETo8ryX4pmMik+BeV4awII1KSlCvF03YYvnYw8f3XC5utSdfqwVztCmi0K/eUb
QEVSEBuUUmy3Emaabp259GKii7i5RFVGIuu9XS8uKUAVFZs5o4NuOBVFLa10JfB7
RcykCC9HIyY7mHPlRCvxqP+v/PcF9IH889h7sKUSB4D+7I5AhDAp9FjdMNE5zYg9
8rRQmz/+MwKv3ACQyPgW1+zH3mE36+hhXdQVoThmxIWqhxY7M1/4L5H48bBUNn3m
QdJCUM6sGZjtYpWfh6SV533GmmvONex/MJeKuWa9V34cXPgtowYMEFuBjnMWbNJ4
pwu9hCtMfFgiqS2Op2xyXVrH/2Tki99L4xVNEOT4Bkh+Eh3MgpXLGeORrOXHLfK5
Y6W8Rj7xhtJwtEJZBhcQKNyo8dd5gFYK+KlEuY0rN+EJfTJ3VsilbOLA6btZR7eX
KlYzNGQaYnI3yxL+I+0AsuUSkI0/KcO2kLYkxqzczemKpX5uK250Ww6qp6HNGFXn
aQ7lbATCJU04IJJw2r7m7dQcOdhZPelAzmhHEs6iT2w5JbUABfXsW4UlBOi4MlK1
cIv1CRFYBp+uB3XeDtxhmk4YMHeuxvBZZ6yBFwPOm3yIkJRZTOHUdnjeINN0DM6O
Xb/vPsZqCDnaoE3VI9fULq7gwmPBDq35f9/NTS1Om+s=
`protect END_PROTECTED
