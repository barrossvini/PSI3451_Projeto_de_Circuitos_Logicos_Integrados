`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HlHCN2DKoi9XP4znCYu75VOPcBADSGaIOpMJ6TemhmvwHoWcH1Bm49071LeDtmzt
+0Aj7Yj1M8ufo5cb1z8QDyQ2Rp9WcoqIj/6/5K9Q+PWR024QPNJYjfDaud7I5GNH
ScdOPQeedaC7VWAPRo7nPSFORa6l0lGeJDRa50jUKiIj6ewrbExDMm+4IMCFG3Ul
TyCAXnroRYTmTgFbdpAw+8vHkDctVDAHLPa+Y5d5I7BDCF2SmxgFlQnNYbuRl9gO
C2xELxszd9+2ysCooKKrlJUSADu9Smpdq7Zeori19UheL7DCYlNd1nMNjGid5HJ2
Co5gjDWRV1cwth6sPkBkNt+lslQS910evr4zPCNfwrkBdNF73zuxCMuZdgISx+Vy
yFPsIUlv3OMSNTSkI82CFdAM/JwhZPGOICCam/+EzN4PMkwCiTqflsAxJZfHLPLn
dMCUErFyofsYjU7dV9oDshDDexnPZGTH1d5gmh5IinSr5RPgi7mI98Zxj2FIHUro
lhegKmSnvHQk6LecCfs79SzF7seo2EH8dBVdl9swha4uWfy8sQrtLwxqyucEbXI5
PrMXjmnVum64Qb2zMPHQYbosWnAjjj2iqG1JeGg7xEQ0bIET1pd/ZVRNRnEdWS4L
G02NFXfD6OLCWQIsT6nxC5oifKQ3yMryNvme9gynQn2BdFxMYCp0fu6egWjQsTU/
olQUBUPCU2d+JytAVZmRAOVcMtO8AkAvl0eposdIVQqtLWkgdyRqNkXF8C81MGmH
GvqxoYGycRQtKrIcN0QOK/c3MgoLWXAkPDJNFYTXoKPMwKRB3NkhD5UnmLojufuK
Nz9TTzwtJWd8liOd+pc+Sw8V4Ke61AjOsvfLMGoVfDNm3flKNBm3BeBNxSCnJ34z
IDROSbW7BkV6Z5SplsJ9eOAZa9Cu+8VuudbW43imuuiz9WiEIffpMSqQ3BPjpoDD
W03PKqH3yxr/zTfGehaej4G+s2TwGmzNjAm84iAxAou+iKCq60TCYXIaotPHbocL
CEl/cuRWuTrgSg5mHePNICIJNtHfo/0E9tpTVrPUGOfWwyicwgQT/g8SAxdmhaHj
o54gpWftVffUMgVn6rDJEwpo8s3kbqEpz7XBR1bj5YvU8+kiSK6N/n4gCJNlBxyO
ikF8Qz4p+3By4jbSDuCWlndNxY5ZMNEXfnUgQPFgu9oCKEHf4T4SspouW0i7h9Vp
DdrxaLv/FzPRzZbZi5QeZXwdX0PupdRX8zFs6CMT4dYKiY7yZDDeRV30+qN5/i45
0sGUv9NMLSpp43E/Qwj+TBwSBy5fSCSe99tIKwYig+8WeANPUo8lsqB/MGrUvYd+
n+hAdOOnp2IMNFmtbV53xx+XnhOOtp5rsBS+tdI45DtXu0rwpp35odvIgLxxTifB
kbVS5Vd25w5sg8wWWnT+xn6C4LVrDtvCDSXI4Kr0MRii/CyGjsvgRQGjc7Wt48T1
luXD5JEtqJ+eqnUP//AKDyGsOmgFtRhQol6dfJrZU9LjobPQqGs5vNvw1IvRYqRb
cxiTRRp5M0mNNm4sFEBzTGzR+dRsyz3LeK8CUSUO1304BfmXdlA2zU5CbKzxARf8
7uKOLVkno76ivyFeQc2X/jdCtD9dfX/rOLzDxlcu0yagiCPv07XXfLVRHIfRiLG7
hTTn4kZnu+CVJlYrtBRQoJ9971ne8TnKzbLiryuzUfGL0FEje5zJ+AQtj9EGUVkO
p2ifgVUMLxBZxAwzykR4AGodzoceyem8Wt/iHul25GYeUfbs0o6ssPWKpTP0M/f2
F/J+wIiqTY52+otuD2G10dR9N+OEPNc0YXFKZBEGAo5F3ZQXhpNJtvh72lWtrpMG
6VOQiWxXL4ZbxF1NGIaPFgb9qDdVb67Y8RXgErM63zndgfPcy6xVU9f5SLzHN8Rk
cwimaf2BD7kd/GTAT1atyix8pveCm/fhxMj8pH8l6xqYrhIwh6xJbT3ybsFKQb2W
mk2E/6h56F0KKsE9UZWdyCEtOEJaj9ViEda3PrGWBMsuAqOp90w37wu7OyK7NzC0
1BBYVOi96xg+tPuQjpijL7EiBAPznutWviJezlxxENp5JHgSfC7NzK4vQv5qnOW8
DUbiwN6WUsqJ08haZ16MdTqPHy6v6QD6ySia5aFQcOyypKZfMMNrjjSa8E69X3Gh
xQMkkV1WlBGwYSq3Z/DWGF1HLJC53IsdoY3Q02mPhHowDJwziqptgnmQWxJt2LdD
FWL2dxSne7pLk+2iQsZI5luzA77CCvuSHzgSoCYXf/kICKCiYv7huiEzksxjkH9f
0U0qRpTqJLTwGrbrJ+OYB9FydPzkh19KC//uNY18o7cc9EDQVS0bJTYyuMBRn9T4
Z3Gx8fhKeK9RJhcpZGxzdvzEa+OKmnNyHyBEzSjmzGcBrs1I0+NbbQNh+R3xpHTI
mmYMuL+tehwEMyr7Q7UNdS6znuRwl6Rvb6oe/sXMA1/tArv1m5OwyBZG6sAuBadu
QRAZayvu+EigKz7sMfPVw2rM1jpuZLmMSplSO6DAFJ0TFnsxw7gYJH16SmbmR2fI
3dDQY5GuzLqEWVbdaRmhpmgeEnIFxx6Uc+WmG39q3aMdsbh/lG0x3tIdepmcVpYO
yR8OQc0ENT9HXL4rTsfgYdLI/4sYxMmdj8QUC09NML83swAOrI7Lu0OQHDIaC9CM
Om3hMqLEgk5AMCJF8t+PcfELM4pJGPRS9HFlGukHMrhFGiXCjqRhE+bCQOYVwtPm
14roCc2VX8zy+5r/fQIEf1xIzorSpezLe6jxlesTQq/0Rso/UGeQwWbsMxEAGPJQ
VJ0/6O6E5ZNgS0uSaKIU7Bza7Sk2l/Nds9B2kipC8XD1ZWKP8oBSfDbtsnUcznIE
H4xAgD3IXjjoPlh48OGDWyDjlQQNbRy9uUIc/h4EYQvRWwBz7JhVx1SN/bgVO+4n
45kYYnjZyfg5nQ4rw5S3x68FgsUlWLeL+E5Te5jO7AR2DPeYrGuUzHjalR8lvdQA
3sEcGqZ5l1SeZXl5gDu5+eMfTlLDIJgojCBIYZTs2I2IxxdhErc6oq78ZwksfkXQ
cuDLELy83uIsT4ZwNRLFOKjYIFq+eBacOuLzEyu3BklR55kzHqXtcH82749NCW45
T/PBOoqXG+b4YiJ04cl3buMRgglvvcEXgZnYiWfN6nc4jgYXB7kdrOLr2kuDuGxx
8B48OYYLCyFO2Jkt2Yp4qju/5GX4arCGoZ4dQogZtnryJ5mSu/7QnCJ55EuBCYgQ
DVPaaQ5PwVkTGNLcSUDRocYCYjGVDYLBC44AhnTnQaErMLliufOvJM9/mMC15R4W
P17v+aLM6HbGBDz6N4nl+DLDMK6czDH+EWyYMVxeGxxgZEq2CoPdtcVm5/KAOSxO
5QZnBjc6v+GqbegZ/AHaLzr9Oj4iWNvTQwIN7FMypK/EmUEby9cAypO4Lar9LUQS
d8Rkd+pWJ5dlFeIYq64dypVP9QFuQpXDHw/FjkKYPiRYf56cFrqLewt3qQFKh7lW
zU6AuyKESqclI7OLxs+D21sSmuGLCm3FVlHZbpXIhZuEsEihmW7g51AjyzxC7FOv
x+cX9gIjlpufNOFRXdu5HCtFZ2jpn3KoMahEkiDyO5zO1gVUQLEbOWo37beK8aQS
gk86+hs9voaUZ46cYd0E6mdYUjSm3inIOkoy81AoEsIG6TlX5imR8WaUE/3vY4Af
95VGXaJAFOAEnM5OOq92HOUTS1lgS7tISM7jMU/qjAxmpkkXTPynfHJtN+FIB7b2
vysNqRS+fcn8eBPQQfKM9h5uuk/Joo/v5p3Udoc8jyUoNnNC6n/hClG53zZGxiv6
V2mT2f6u82daZhb0y55nGn1rn3tO1yD02n8H3S8G6Lt9quDtA7bGnnIOsiCOaeN0
RCjvaZXSNKOy/DdLGtn9fQdqZX+mwopmAzA4OSAffAz8xTmoHnYhoAus4jKWHIEr
pjOx5MnkkC+GZ8TVi92b93QiXe56MrHsHXI7B2DpOC6ssGa3Gqjv15BctddcPMlj
lpDTi0HPbkvYtLbhwXiwU1hs6hHH0KHLNcuAiVWFggoLtHGffBTqHyaWdky4wb1w
GcFFS2WJwOk72FulEGFf5+vOJF3h3YoZ+mnjRSbXhCCM6C5vd/wylxWwZJSLcxFi
7as2jZrCmT+5kdHMtSFV4R2is1R03UnaYN6TtlXLAxFNqOQNVajMxt4cOszwfZdD
12nV0HPigTCQcUzXiJGkLlApbCWIf21pcjHubwhxb0Cy91tIAfZ297uddUUD95Wp
risuIn7J+88CfYAEwYx1NYSiOsQ7nWM6ZKvLz6bjA4bMTd8+gDrfHvfzJarqO1I8
EqS3xk5qJblb0iBnyoVEPELHYYLP2jK3mn6oFYn0xS0kN5DDcRPBaIzkSpySdWZI
LLut+u1dzVH0I0csZoQpacb68bPZ4vOPAJlOkLBtqu8KBSo70/97IhbYjqhtndKX
iYjkJy1K1KpBI6dWNlpfbI/2cW5sqRJ4y6vaLEIMXKQrgDvPKcRvwH4aj1KMNjWw
EZDKQWEK7ZINHf7Ck4hWpnwb6lwCdkk7fnwEx/TxM8umzbbCMR30U8tfFnpwsjZi
5ryIWb5IAEIGRn+LP/VF4CFeStq2133nWxn+KphMIk5+0l0m6AVRidY2wI9sRfum
cjpiVBNoVIIJFkGU9U3Dbhk0caYHAWY7j04RWnhQT6fm/XlmehL8sQaJUJ79Xxpr
3yaisEMBNWn/oI78RdOg04cIviXbwSFX+tBDt9qmwOHp6YVMvi+kIcjZcBkRZOer
OaX/+kG+G7+HBT5VD8OtOY7+VHi0h4CCMY8/xzNiUmZBURz+q5E/bnF8Qg+RHNLT
dyf3osNByU36jpI0APpTpkw68ye6eYWBlD7L7WI+5DqBV9SSoVLSw5RMJxCpWIyY
tnWGqsjkU+FYCFUwsiY0LtTEBoGbnE7Ijxm41hF96mQ/9biu4mI25qhJ1SNOpMTw
jPjxZ5jN1QkI7kjtl2v4waTDe4d9RjRJGijs5uHZ8Ej3SW9AT7xjl8UaaUurrZU/
s5L9v5XHy4aqPASHPicAHTdvjJAYp3cM13G80ieJfPSzMkpF2MWZE3nN0Dd12o0K
PA61MoFfttu5vIuIlhiXlgphWGIKXjVyluR/VE6GXQchjPZYV8nLcB8d/em28Co7
etupTZTyo0P5cuubh9ZP6iWjusffYsetBPwJm+ECwL9QK8azIPBVTN7C6Ac/Su1C
m0/LWN/R4gS/TyaPQD+8h1nHIfO+YiyNeao9LKxHl0llcP9oAwXU9codijdmsi1q
mmPVuX2UZuV8xQiYgToZQXKFJMqQL3Ed97wIgN1Ao7swdfmM5oPTdAn8gf5B7ky9
hBc/CjWgg3ly96KEVUPkJ49zeH5aJKlB0//A9Y8h1RbBYq96SqBeJINbUPPaPAP7
kOu9gK2eOyo682afwfD8Ja+gR3S5x8PjHTSxQXY3IW70DtGFt1KGxtY9CYcJEzSy
ANoottS17fpDjMLmnwW04rS4Uq1Z1swdnpYEJYRsvTQloKH9VJYiVCKmjI2V93Ov
kOM6KD667lEaMExeNmY81u5ujCo8fmSgpcvXQR5VbsA/p/whiOSY6DOquathiIbH
UG3rlY2vqH/YR7wSS2Taj12yzTjllK2jfIvuayrhJLR+KsQoIXVPaV39QGfUTIHR
xLKSBm+fLjPaXOdPZQEann+obJb8UWgp8vMXum/1TT53Bz8v7dWP84WByZIwcBX4
62ww2MH5Fkk0mfuij8A870B0p8LpMDS2zPNjPWerHkyv4z4FBWCAc5U7avvp69uB
i1ZX1FkvNCnRahQekZqF848k3e7uQlsvcpbQxvQT7fC2HMZg5Ph68VRTqDkCxfj6
zJZyVIJ7slniY4pY+DsDHm+kEp/aVOCfqqDMoRzdyEkL8m0ZH5ywNb3FTyvl6KPy
icSL6amTZJqUEscwo8hLgRDOpzTQ64nyjcg44cyYMv1aI1iC+G9P4W/rNqYhBy/j
BR6c4DADo27RMuQ1RhtHBwBRvkivXcB90I9u6Dc8ZizeQRQBPOefvmJqhQO/jjuS
zmU5bNLzGcqorOYOkwqlxI4b5Yovs/Rt5nP61xl2nMeuaYJB/LJs2iW3gEXRuikQ
aVUR/bdNJ/KbQvH/Up2uCvK0iAsWQ7MDbZCCildI6pyjtoE/t7KaYy4q9PIh58tQ
+g3m0ztsuxhBfL9YU4Xa+QRj4Dl0ObSbtYRYVXdAcNWbQkfm/TAhY3iemhhXkWix
lY3PGlbqaGSjQtAbMsXd80H/Mq87t2kc7buZ4du9A0pvSSFcSDsEMGE36Z1oFEq8
7QhZBvn9qHcuCsMVqV5kCJWH7v7Z+VGh/jsUKehAIFNdp0yWsq+A0YJ49IlvCWiX
WUVfnNpeeUYLAgbLp7yVvrUF7Xsx7hoirzhoSZX723zPcJsKYxT/tbmPF0tM0jc2
pi4e82N5vO2pK8lw/HDIJPPu0a5lhUfLPF2n8208LvxhHmXAybaUov7Ljc9jk47F
wdotHpgsJyOIZV0bwfWQ6tXx+Q2ZTZFez7TbMEYOvho9ovbOXimvxFpt6vPe2kaX
J+utJfIKrgM0q8RPgIk56A27TBEmrWd1jDWdm8BT30iKG1taO8cywNanxEwN8XGo
x0GUza5TVjjvjCG6/4soYSm7DFpYZTfrD/6RCvk2v9R8kmJUIPXjPn9oU3iyuilC
KhPNBDtJVGJVTctSeJEJa7/Q5HvH1RgpHHfD6cwjfblX4uc5yWBt91cPJXjxYRxN
zy9Ij2tp8ren0wmvb3INUSQnSWQwKAsE8Ppf/JW6g/Sy6dvMwF0Y8yAuIE1Iwf/G
hHAyIN/w7I+qX0oAeL2p7r+QInMc18aQhjk+g88JFBQF5II6LOsJQ/rXde9ap2dX
TuwZLsfwhTl3K83q4gIMd87HfjkvUpuZgB2qbxWQBYefSepettdtO3qCwK1ckzVM
eZ4umQ+3dDCD7zrqOb1jzGlg1qeLtPQzP4vT2mT4W6mNpT9ZES2ReU8i5UHjtVvz
WwSl2MGE0b5O36eSVSKnEBYTp9+JzSIqy+9upQlKgXYiVJaRU6xGRFvHoW6NMWfk
uDwwmvRyFlNGhbN/1jxLCRSteHyhQ+86nkfuFDECKwRm4UkCKNzsKuSlDbzvVNWq
vhRDX8vVxf2L7T+j+yvEzujCQ4nZwnsrKowdgKXm3YZyb08L300T8Pc5PnyRfnvi
p4/UHEd4fJKCap8pJDJtG4C2TbGjaFwbko3ys0EXRXQZSiGIbv5weK0t8ndiFIPl
eJ4W3PrIBXhME+PbBvieMX1MwzVHeuiLsvfPXKrsn2+tfgoD6tmnJKKgISC5pMnU
MdMmwLr2NmLzwfw0RRB82wBkAQHULOkZWG1wHsoO1vluEcyn9GnFSlRZRlCD0m4m
b8bcYJtWhipSlXh4rQeSfwprZpklxxbBYEXpgj+lRJy4/Z4txLHQKDTB0T6HM/+3
fXD7eLzQ9qxozwVlLwCFVkZcnB9//OrnGF3ss5qRkkx6mx10lVfJ6dSGDB6cW4SE
FeR2nMCJIL40stxfNF10rWLnAoXBHfSw6guQmAcvdIwEX8yZt2SBQJwZ89Jg1Xya
niZlEG2qoDdc7Wz1oNOgjxIHZ1acG0xBI0W/o+nCpNLRSm4SNLpKSabmtp3ZjO85
KgdraljQ9FvMLLr1lpByG/XZ3gij+quvXyDqofV+IUM7s9/LHVrWfPop7W3qJjf8
Z3iAaPOJ7+CiWGwJulfJ+J0fP8qM7x6exu5FeZl0SiHoU/m14+l9A93Wby0RkShS
5NDhEs7SA6r7tA0BcZgUdIbsueHWHV2pT+qkvg02NEYsTCvRvqrtsi8k4gN1Da7o
+txr6NbCmTi5bA+CTAwXY5X/oR1YqoqBQihFSz9M99Jq+EY2O2eAnpIa8rd106Bx
Hdo0FZZh67C5R4gciwVAWRJKhXOCmmrMq8KkEb+EpSTysyhzVvYaRhkiOImp1gpp
2PEgMWGt00L0yHly12CcOmIayAOdUYdXAFb0O2QDFImdtj06sbzRoOm6GzCdVWli
Af5SrqYfFKzXtny53etSITGVuo3pGvmoJEXNm2csZUb4nggqEq14hdezN44Z/Mlo
x8VdUjo172dbopVJA1OGzPf4wpQm1kkt1a8Ocy6iO4+VY1aeMSkgRHWpDys2pBid
HTDsE0kuQSICO5BMY9fud1FgM6D0LVvt39ZlxO1MYTz3g8o/rpG5oKJtxCxKE86O
hEbgrd196tuGfdCPG7qelj/8fBPQZP99pX62ttinXegPVbblPiVVXUOrOjcFftau
KtnOYTSnb208WAiizyZyt5vtOt/ROEAU1n2sCIi0JIyRzOmVVJesDRBBNF+f8duI
GYZpbJYFvG2traAxYWq8N0RUiRUi7KJpS6XTs/5fsV9/FJtnjwXq4hpzr1wtDPln
sVICYLkYOKpwmZfHrJslskQPPXUQoKNX4Mx6uAAjpcTzJUOJ/5KfU2coUCDvcIzg
SjLYmNl7kMQn2sBNdn1fGLktdqgl2+eUYARwgQPVvIZJhtN2AtaIuJGDNX3KXaEU
7VD6e5pkGrQIqsqYRVEAR8edD4QTOVXuG+RUX+OQZpU9qJqVB3WjjmMOAH/SGASA
Ny68oI+Sh66YwvncT27KXCMEwD8221p1Cr1O5frfvzHJT/N9pPZ33GT2gFu4hlZA
lc7/TvfVOm2W8/USt11rQXHgc28Fig0oC7h2F1ExNSBh+53mVonPZGyMfzUdUg9h
gNZ+MacDh3Gr0DLvoA6cUvxUcomJ2OaOY+8Sbwadd+ERSaHP2boEUqiQnDc/Tszr
hJAKJk525WTm537p6zrVkS3/wdjWjRwhjy/FxGwnMGFpmlNHBYzDx8b8Lm8nU8VO
18ph/POOzm3dR7ofqBe2ke5lJrOTudi82sjMQBW56Ieu1yYXCnk0Tsjf31iUCKzM
0VOyCD63qPZr98MsJ9lEzggYUx/p14dx0Wn23x+0sLelQfT0tFRs3HumWeMzdsZN
vers7R1VG/HABt/XMm2IHaFPQaiHiynECkryLHAQ+EY1kn7SDhZtUQODeeBkjRF4
Jfc2P7dXsgYJ+LMyeHCR+se7IXISmVVcSlnaFaMXbj6ZVPeBK4Upz6MIg/G/DrGx
MuN6x8dSMbB06meAkRf7QztEmSxFl59svKNJk9odLF0hzRt77qGPWuac8m7hnkHn
eO/kw4Avsijf4jhDFNMmnlG9G3lukXwoirqJiHEpStcGaTwaqZxwUPqlp1y2c8uc
56jQgpiLPuFjK8oIglKJ+yLIHMY3w+B7iGDe7gfxHF14eKF8Xy6O96YpEap4SVn1
jZYG7QxNZf/oDFGySqMnDsb7VXDtqE3WErUrEEu69P5Zuprld3van4R3o18wwaTT
BDMqHesyp2gy/2cE9GFW+xt7IdNESVKgQ6KHdh/clm7Eorer7p0A8afqYWdDRSOR
5nkjUwvnQR2H56FPLB2ieBOG79jVN58nq7AGxZdJitmmnki+Qqezx0mbScpzVn92
0trJknIx+f55Eoq1M7yUvLGdOu/sterRxy8ZogiqtQiU1YNJvb5a59Z8LhrcTIyZ
ZwB/CIcaj28yNffQSC9aDwPgBPFamPaftLbFxq26DJTUAJ2hNh52hs3J1f5c86DJ
UkQfOdDfklCxFTUjqzQaLDXN4FtYeCP6Z7rGb3AGH5J+XoS0wUUhnUdNzdQGRlXo
bv63uFFSGkXpeLl8jZ9spKjMFWTj/LyLaD7y1G7uodnHj+7wbjVcV62ytEl2RsxK
PNgqgck1b5oG54m/NJRmP0RWivkMaRBHh7Xq88tU8vkvZlaH6/DOklrLJN3Bd1Rv
3tdtNpS6HI4haCsLZeqg8TH12ikVLzbLpcBb1tX/Xc6acYE2NQamDRwQR1JB+lpg
kFbvX+XJEkSEyucx9NZWSkPYkX1+1PcCtLEHL7K5nubl5PV5IQm+Qf85f4kwZSGl
PP+qGKL2Q0jz8Y/OnATvxDiI5r1OafFB3zSUD2mzMQEIR1euLCNWwbrG1HjQWFnh
TcQCRUBiU94/edRbl68PZQGLuJzdWJ00AoyRzQFoNl9lekoKTlp0bvF9SKVKXSWl
CT4Q+CW/CuTmIkIM4Lobhm5ScWcoAxwx7r+GlvmYl8N7fsj2KqKBuzR+PpuP+aZ8
awHgQsJVnXSdjvgpcC2Nk0vMiUNJl8Yn3iJ/C95C2hpoKW3DjmuxtoxvwSCuSGch
7/zjJEny5A7OhoBpjWORuR8/6b4NIfFLKY18ld/5hsDAWop1sD8yruLaHI/E2vvU
J3U1kUAsud1jeiN0ZdNBY5rFwV14UuxeDTFJkVy/eHP2locuwBRNqET8XmK/uysF
HBKwowWBUfUxkJoIsoJknkaJ8j1vZJSHARGV87lInyqlUEoxvQuUmr5WE3Ff71Hw
cUpBP+JVLcXEEzrr8VlYW9zyvGPp4n+EQK9kGpTRVDuqjAVtO9UOK/NPWwsJot2E
tsBuIb+s9mcEp/PjfT+kkjIkQ019Kj6JG9bR9TM+dTfMoLhm9JXXahC9Bw1TIpFA
fdVdmsvdkcxHIpq3sukBArctomI8wXIFlZZxNuI7jC73e4EeBJyFKy7qnYeHtFXD
QEe8MwKWOHSxiyJpj0dVFVtp55AkDU5pOMVLbnEazt97A1xJ25+Gb76vgReK0u9H
J9cd7fBR9VI8UvtmaLhrhL25oOtMLb8vjL1mDVsbC4S98BoELIx1AS0s/5/YGiiv
pKaN/VnvfKOldtuPkJTiOr8Of1S9NMCq/GvwDfChc8g5rVVYFmfaC8VkH9YtLb+r
CNslKky0HGOi4TjRZtcWqe6L424fzmOTvfA2rqEQB++q08BR512IHRyzLWKN+kCV
xtcf/CN0Hu3IqBUMkvI72Fg0lbc+AZOGIe1JJjYdeB379g2rQjczn0MlY6Mp1aPm
RwgfRGGTMqr5T7rCPUSvRtPcrO3Fqfp8Zr3J/CQ7QxCeJjmrzSY55phK9M18YSQ0
CaAc+k+8sPp6s3of6tcw0xGxTD2mXJtvL0bRkwBRh/VktgrqajvMpwMS71SncBqK
YVDJv6OHeb8r1d2vri94JPVXGPCDMKDS2ddo0C2UDkY7yzQTmzwJehQVi5js8fYG
Ser7gbiLisYpndjq5kpNnPspq5b/Laqd6XU0bG5CbUf6hUm09YO4mcwZSghU1iXi
6ePqla8+TRcCgmlFdjk1lKz36zYgk5jf7hhezpuSKMHtkDIyz/968EXRVtcVcPjw
SUkDwc46EKeiduaW9NckdGCxOXhHLMIAJzx97JAhbgM/wh1+cUGACpGsCPGC6Q+H
+7/O7WCD8e0/h563q94MBFBrNe8Rlvm8pddoJB0GhYAaZ2Tr/UcrRhESWiAZ04Ng
LfLveIU9XYX10YDKtsDLjnii6U59VFs3lYfu+W7vuPAaGSjqKSRpwu03dD92Dha3
0GH8dDRsegeVBt0K8qFoXpiR9QQV/VpMMrTZBWIk7DHol4w2hEJw21RYkFenLvpF
vpHRyYcK9yNLjbZMFu9cF5CB61kknaTwuw9iDC1TXEPnZwLH8Iqy2gKnMffuBDV6
WT7bp+XKUznC0LvzMZzZSEERTklsXfFVoj1sWSaIMEGWRYzCEe130ZQ3LPxhMzIZ
g1BWwhcgrzmthHZDrPiQ+V0t2DmtHtK5Xvd1y6NEPzPROoeQpuE/mNaZFysOn5cB
2fIixug3RdPuhCibKavnfILu6J2OVnBemnDKz9cwAJxE0dohIzT5/2mzJvCil6bH
Djkc7qcVOrZJKU453goj9OiYNou4m0djqRc5+Az3y75TwnKCnwxg4M70aWr1plBv
luENxQOOrkfrdaMeoeqJ5T16oxEfP0Od4TWmRCddjI9ytXnUKGhuIIAFkHi1Fy9C
dyxsQpOml+FZso7uH13EQc9JUTET5TOQGc2/iGfUMQTr90dLjs6YTKE0OnL73k4g
H71vnnOkQTHqHoliOcdyMJarI5CluuN1PfwgPuFPrDGbS73aEvfYI+e+KkkFgpC9
lKQTnRuOaAEouc6ihNws5K4eo68dc2Dr+jtONWqVrvT6TY5nZ6hQQhX2a7KgYZgp
zwZzcY4Plm3Xag4WO9D1Lihnx/24MqGaxnLHXwJMSoqBIroKTG5UyKFSU2FDvfOo
3OLZQi00zaJqDVpG8z0PhRaGrKOzNUsXbR5V046WD/4o27V+mmOghl+clUvwfKBR
5CExmT6PrS8Edea+mWwbXnoRfn4ocieItmJZH+QL3mn3y0fP5Hqtjusf4CftNvdC
45LSuxYTiByzk/HtHZmwbyQpcB4DROJIzDRf+CbFShKhuL6XJJu3uDqt/SCAeLAy
ZQgd9iG81Jk6RWdUQI1b7qmWuGynX/jbknEqHHdpSx9WRurfvCJXcYSqcZylhks0
fjOxyC+9cOE5FPGbRPFL+KeI3OQTO7UnF1OnvQz8FWBAW/42IZOmTHlEPrYqzDNB
f61WFHmyr5PrNkQxhFJlyU2qQhUwO4aA9/Www10pd6kxu2yMK09AiHviJxYFb8IA
1eYwkA5jX4jmZY0JwyAxmGbywbPtYIq3lx8ff4zWAMcFsfuJvBPVn+3is/AtHaxp
naHWf51TsLyNUX2Se9Fng6B9AFuoxmG44jbNJI2tLgnnDrCcumbQD9EsvTzWM27n
yRezN7k40QillvJzezKKUeCEF0GQkbHZnftVsS1fP2lOvrv2lBnZ2Vx48hhfbJ1/
h7nvgmvbGrfucpmwNoabjICuJ6HDDnNf2sZKPUvd78bUAIxi6Gm1SJY6J7/Ob4XR
nR8VFno9jH5SEpYWEZ7FfOZ+aLGB2pohFVpRiU1QATonLjolY527kLIZYknjvFe0
KCSiWcX2EHk1JuKX4k4EKlpp0SMGPNse3r6v6aTZXoAdQy/dcPkZLlL4fNQSBuIv
72byn+oXGjcdPpfKY7sL/u8uo/scTWcMPOBZb1t6QsiBt8C+mMn+glTlTEDgudL7
CAtihAazMHIxuiNas56F5fHyMQCbtAlCQW/z2AUVAivB1tw4M8pTEFBFc9qB6yyu
h0HIn6iFjXeXghlWsp6mZ3YROLJwZygRTnnDKJHIMOtpF8p3Igr9Ow4PeohCrj8m
KsPnaJkci5MD/tOJ3OzJyNJ1aYn2mDZ/Tb/ZnLmYhVaas+burvvaO0q4X4ctJQkv
GRwdEXvwIvEQmaSkUxrsgJpI6S+G7Gvt02VRZrnQIQmSj+g722+ke/IH/algxkrQ
SlDIfKC51OFYcCKy+1KoX8GVpU0Z774CDzvbEC9f5I87RULbNdYhBPVwLquauQlt
Fm5k7yIjGqtygiSCkkPf9zBzXNXv5m2cns3JNboqNsom9yH3eq/ivkSfftsuunYy
tL6n3JTSvwsuMwfQBf4nwLtMOb5YIF1SvT97HM01knD/CNazHf89YMrkzjDAHEv6
1E2OSMZgPG0jX0JDLNnVAMMVkUz+PNPJTJ5zkWWqh848MDMjNCTNF/vFkR0cUq45
G/Uq/NDNlOAXjKJ0pW6Nxe5wIi4mt2utJnbFEpc4sHLkIl+9PeWmxL4zorigcCAu
juq/07HcozLL79U6pXgEVUSmpHwA+LRqANu4/DUZNM26i9Mdjwc4HRU63qbbVRZw
l2XPC+mDWVqtoS8OcjfgcbdNbstxyxr4WYY01HOsLc+jyp9QDry43lSqVdEEE6NA
RDBYA84XlE2/9mckpqoCBPQwoo8oyxhY40JI8Ixng3F9jLlDpdNhL0TSxgTwlS5e
5LuD4qLz4TzNouf9t1A+8I5yFQ+DpshPrW9ygOuSS7z0OgYT2uOmoBQwZHxAOwwy
8NohQcLfNSqJ06BVBNHWrqaRlTHw9IYKPX0igHUJmkqzOFeu6jqwijNMl7sBeTFj
Zhr2Mys4a+t9aYJLuZWha/8nlLoRtTf4ic3rMab7FDRUJXFpkX4uCztw2JmUxE8h
r+DnPv1UQFvv3RyWzokICH3ghQM2S/PXgRv7LbjtJA5t4GSbfb0xz/s8wHxnK3hL
pdSr5lHiaWK49x/hPxN//lUdbQZWz6laKyY4rUxwpeBA+lwOmngAG2/IpQeSvgDE
JcyMunxz+BMTMsWYkfPAhCc460DGf/n8eAA46E7KSWK3HQP4OCDqRcGtO2a5vE1g
JhdwxZLvhu6M+K8Y3pGThl1AvGSH8qSY0+mUEDsy+W8qCwJVsYkfk6D3oTiKECnh
Gw9raVb9pPkW2X6mTtX1LizQADoE6UlU6r8gYnKUZccGutfLGUByoyf5R4Q4mBKy
68BKQNKdy1MctwQcauAyb0IHZU3xYHOpI3NPmpkBnqynhu3BNTkvOfP6Fux91PJM
t0K8e8IkPC7E3FCtoVtWMHauZjejpJd8WDmZCqPyqWJAhYBmbrOwqBNpj+UMtWTJ
PxssQpML2nrjLcPAllJkUZ3BbX4gvEXdvN9SSgiPVVGe/F/VTsrsjMNdMaVVlaLw
rV1UNrm9gEdrW4iH0FJV7ntXISzfXCGHv7/VsEm+ogiwaikusDE65s6QUagaGy7j
CxtocUaq58ulJt387jmGm7Ckh2wvEw/er3BVk4d6F48D1xNinXbcNTIUMTdOb5H4
4KZdPjXVe1ftk76rU08ra+FWA6o+k8dP5nl+sRvsENtdXCoTP2QT6uezcLijT+F/
RG4ABlNutsagiiT2kVPzY2CXHhkkkoJyHrNLJjqE4pT1Uhbczq3kr3YLx47/I6Mz
Jvz1YmoPPXdb3spXIxnT3WxbbCiH7nRbJFpLHbO1QTIxB0GKlSyD6JvObeB9oaJr
5vFBFut/XxS99WXw7w2fdQ==
`protect END_PROTECTED
