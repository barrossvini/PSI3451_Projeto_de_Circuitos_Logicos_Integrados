`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gPFGVMjU4/zHj/l33+1SY25rKUQaobUsALh2PYOrW4SlyxKenzt8o2Hg7wBt4j4Y
jNKGz+9LjJx5Y4WKMbnGZmnojaVfBrGgqBSDx4PQSKGcCvqTMLBCJakmtaAqDfav
Vz6Df/leUVVfgj4CmWmRHLyQPlJEyCphX5UF07p+PCdCSV+tyaAUbKrdjXD1c7UB
LJo3pBq8My9dyvqQyV8AgVxpSlEzjRwSnrJXQuCUJ7eF98VY3LfRDn4cc3f5e6Tn
4r4GJM1XeBM8wItiyXJouMQdKV7ICLnr/DXRLXEJBTbDbynm++c88bJqv1eaZevF
tbAHgK0kzyBvSYC6bnHWiS4kmE8u17tW6tLOA/AGDxrNjnkL1sfKJPOQx4CLWMjY
Un6h9z8DsVjinlyJBo7C8BWHKmr8W/AgxriZe+VZB/O02GcJtAuNudpskiHQd89c
ofuk3U6f3viqLm3LG9iqSgxf6eeEGJ6vBAkeVXRLoJZJYjcWk2CScPX7rDHe0lRc
/QoAHVc8A7gN1FjudXesM27yOV/K7/kpAw+4oXFYHsmNaPp82alhghDQ4jnBlE7n
4gTEV151f8gfHUab1EqRf1BMymrsci+w5LBxtDCD7kq4wh6SfAQqOSlt8PDsqNfA
1x9toXFvKWf1QEfyLi+its2c6gHxFBk7mafphy8wli6tt76ZEZptB/BPxnH9xTLz
ynNXd7vSFN26EudG2Qes7ZuY9B18DcvJSPR4lybzzSp4oi1W0Cd+f6JT1D0Z0a+2
aMIhEITuLqTlGGoB3wjpHCTLU0l9COXIGWlRIuXUwnBSNprVVyD92hbXA5oYef+D
RqZceZGef04sC1K5dJpFspPPf2jSLib/3W0P7ohlAe/YJa5gE8uAVdnMAD/+YJPe
btsbGin3fLEHjGQPZd8CpHt3ttvTThASCHhm0akREPtS8rWeytb+7PvGXYiu98y3
c+0d6qZtl0QidlP6Hkm9jJgXdXAlQF/44T1R1vBHA6cm411ZY//RaAE9okdWVu8a
saMFRWoaka81FLIxlrOXM9yj/ffaJzauITzDo+lS3mNVXbmncw6trAB4zl3w7qY8
nAb32didxkOdYhjabsVIG//ALaDd7ClV44dnrChlr3Z0HjK4e8f+KT+QMAMzyutY
VzZlEvkHMwPz7nnrH6vUsFfNo/bQh7hmAJkhfGzFS0UtFIzDztsP4lnQub+BP4uJ
rsqhQB4QR1Qsl0YKWfN+uMKe3rVPEGO/Gc3BYgvK1YavkbTcnbKxdl0EHhHiXGbi
`protect END_PROTECTED
