`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NGL3eODUvUdRgpRw4J+oGKplQOHYoNsRV+uFzzWrnTvl9hIAjYT08AyaBq5LI/bM
0Pk7JB6PC0BEIUf3WcZD/YZ5OYO0Krlb0UN7zWvW5Bl94o1Wa00JDCNoqdQBqkj7
waNuoCCVFbiqsxrcRnAnFnEJ1NXzNIQcx5axXgZcOXGHQ/Y5yKziILGXUhej8ZzK
TcoIIOusKtnC81X5554MFyFXXNys4MEMFqygW3GVsNqOyoM04r10c4YuQm6oRtVg
K7aoe4R4t4VnXH9XqmNHHIJvYyxCJsz+lIrcXdXs1i+SgVxTukRWf4M2NN42L7lG
1o/ZKekTGeUlIzLuFsRsHcpBchqVHME1txk29+gFszt/CvXlK1j550sxvezUExpz
`protect END_PROTECTED
