`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
74ri24M7tx7ndApdZr3cw3S+SzlnssBF+trYbtNTRwRcO53OuGmE6NJMwOE1TUmk
OLpdAC7TXn8DKGlePB9vmNYWT4zvX4dqSy9EWjBtTPXDe/GoTk1lJagi1Ln+DZGE
bmIgzeN7BgDVPt1IYAxjaJMFBV3h0SjDbSVyHojm7MZU9bQfpo1RVEZNtLGI1/5p
UIzLdUjf8zxlXgUg2Iq5K6ROo64rynEFAq8B6A9Y7nUsnoE9MgCs8YDwlFwSlYY7
9zSa61+oHTef1Iy5zGNny0HyPu91LmwUpm6YZdEc7uQswO7Ixw4NWP2FdBnzWVlA
5SD37ejEYZfJIKFbeDkB86oTPvtZ0KurHVrfhhQQLqR9hpoYQqtESqJVW7r/eXAu
EqwVTf1AbOO9gh75zluVSidKzowSbgZsgw74X2Uv5+NIbbcJ2Yn7FaA6dLwVviuL
xR93ufgXLCYCUNZDa1mjo9o1qv9Qi6FZGfNCLDX5m+vhh4gif5MgJZS/6aMncb4M
j6f+INAqwpVUKQtzeraPFAfwpcSPdvqZqxhyGJNsk1yL7efUYaZBFoAgkK1FqJqX
xFFTXYCwb4USFJ03W9r+8TwU/PFSK1h67dKmFaXB8LoucOgIH8NBgydyvmxt1YSE
ghLnABvlKHWNtHClOpPvZaTrXpkozx1u9qFh3w0U3s0YPUr0pPoSP7qowXXXwsKt
DXO2U/alewXdoRz97GknXzwBJXtobWCYdLG0d9pwDvLisVQWT8qusZ+re0exvAjw
PkXYMRK7FrZHnMQc/BQJD9iyOITnJyeiFBDl4SEPFm1NxKLWifOvLksJl1474r6b
nGxTMBF2PQu38Ns7R3Q8SZyClGjrSVmtMTc/7OBhuXDGYpq3cXHvyi8gXgIQxGjF
SvZVaUQIq6mfu4i/EUPRIo0XL9nmUHnEVfu7O1mPrOXB0ZMo8gy+39UsI8OjZUUe
T6OWc2+me2nad6SRZK/niaTXJiYVTwStetunUOxsuu0XiGFh0B/UDvR6Sn0d2CKx
4Gx2J4ppfSd6Xl8A9JL1GlN5ncX/7hVEafc2qAE1QBsUjoRzGrZDc+oBCHfPn5YC
4jajbw1V05bcDQwDYlK2CSi7vwaWlIxN0NKTX40fDXq+UM+sfhwjcT9+vg8zJn7r
n3wt+EGHSZT3Y9ndB4TCxVFmkS+F83IOF9GOL33Xqg2mbzLtMO8bM/+FFgWdyGxj
daMSev4ZYwYJdYZWAQWK3DOLZxxey/KjNMcwNoJWf2YhFNUOv6/qOr3Z1bSgRZly
X/t949feDDlE3v5gHOIwLi7YPdOIz5AukTVztYkeclovIr7SjU8TMRLfuTNWs6Od
+27bdFkdWc3GbHPTMvPiDYtpXDc/noFRQGxbKFYTM1ZMo0+BUdqXCADnMquq6154
gN77NRUJ4W0UMdXe2kS75VfF2/Ue2vFjo/56fauzurssDX4Pe4EPcttUr8T1uOxj
XAaeKjQIrhcQkd8ITNgNudNXyOOZ4F/OGZKzdb94dip7PixZpohmB292ZZWHT6OR
CmMVWae4Y0WkRiL64yHjHSxprDhgZwigymlnXXikZl1xwkJvxSo9ONXdU9mAmPPI
GMgzIr4CdZW3qLljykSQVulfgXaiXe1R94DJai41D4OHm3LPAjg3iGIcuaUgY1Lb
tUdGeUH2ymIQ5evxpKbuTw5Jgrmg+xZfFnNa7kDctzlFcxCLIlFsJXcd+PMR6UkV
2KrLYc2e6ntElirdIoEhazsGI9Q7lmI3tsfD4gfChmG5n+G4MTN+xPvcyaCDSh1K
b/s6u51QV2wkMPSoT6ViT34FjmeUhIABkQXwZ2ugiifoIgpbAB7PqDYIbjr/K0if
ZamMOGNp1vach9/m77Acl6fKCyH0vSUYoHXpVRciypJHI8cr9EyFvk7oOPap62e8
UGGV94wj/AqWXM54Dl0N2b5FR30D7/ljPLyO+HY9+uw=
`protect END_PROTECTED
