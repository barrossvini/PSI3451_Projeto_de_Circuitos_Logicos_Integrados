`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BjyLMd2gCtzGnp9W8km1uav76yioJN26KuSXqk0RMz/80lT5An/nI+iDByesR3MX
9rI3+z6EBr1tb1toDmUQ1/Q7TAZji4yAQkYD8ZhlP6DHGLt2g+7R5KzMsTwxlDZR
MLN+L/NSa7ZNYDE8KPO+k2kKVmocPKWwpEBVLMUM0wSu89J8Zp7IoTIaoydIi9fo
ArjhGQzt6L2PU6jfOnfUivloX4FcRm48JyJ8uuZMtYyV/4A/9u6avUkxbxDyzxFI
Kce65XDJnG/UydOP8qxhKweStLQAAzcS4gxrFUd/hfbIyE+HLOGc48rvNUK3kdpx
DHESTSeTAlJMYqttxFiwdC1Wid5VOY4sL39WKUSLbWPdBG3PyZ5Fp2P5+/gSB5ms
QcOl3Rw/vyKPntSOkTNZoeYeegOHmmgN4JersKji9tFuGSuR7ImWg0+m/vrm2LAe
ecP7vnOcwjvIH0oFi1zUJXFMGNcuv9XlQk1SyZgbCaTUAPRPoRaGmUxgq/+BITi4
zXSbXJy+/3K8Bywpqx8AGVKHDH+y2deOmsSOfhYhXFKR3LYb2rcbdUVIAnTcbcjx
CNh/Gr27X31yIg3cCEtIZ9eCQaXadLQEqNA3se21ex6eZWk+AqoYAgXZbcLfl9Aa
Sgb2NQ52auMU6pndsVG6Z2EJAY0d9RvswbWUDHGkCnRnDcF0KFFqRALnBphy38Bp
roG7uQYX3JbB1pjeWNU0iwZoekEXWijq0oGxjck+7tPEr0ar/LJnP1X8MZ0uMSiA
L3mebOfy6HxLxLT1O0SqSW7PF2ZR9b5vVSR5wlznh2G19Lv9No3tc++lp3j6WnsU
6ajXHxaJREPIbYkup0xsFqZhPCDtabnggN0kWLHHjXBfx2iENZjgv7GmXqDL5uc9
cj1/F0UQNGkhQX1ijsOR4qwCqQ9GKr0zTgug33mEAVjeLtSz2kOadKZbbVkcd7+X
LGF+GX+Z/fW6UDCSuiJt5upTrxV1j+ihMnQDyVa+nNlWw7fdyz9WAiTc+zLDgYhc
RFd/4oBrjRajwJ0vDuKsESfZOZ5tOwIogeXG5S1gK3a1hJMsSR+eqfloG2Y56+ts
VZ+0lhSMQBNmohj1gAMmhw==
`protect END_PROTECTED
