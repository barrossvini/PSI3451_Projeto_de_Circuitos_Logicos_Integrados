`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CkFJp3sQYEi9IxhGxvqcl4MP8xLeEVFrZPJDh8t6ocqKa9ZiYfC6K4FgcMTp82vb
xav3cHDOaKEfJ2ai7tChTcAY09XBY3KBb4AYxNzLQ6IvUZKA4d/+oZGFtj7S4nzn
WM92CtT/1aaJM1N2qvFtMQaxAlmjlp0I0V8uB4lWa0MSS3jBLz21rF/acNghuO4D
8t/Dn9f4jJqWnKhdfdIqC9V6Z3RzwOkFaaRXdUP0IBK0fHKfkADMhkS9Ty2Lg3/Y
gShmgsMUk/ebpK9yJdZ7h3GhLiJrKtZbqPzYRwP5DwZ1Mk0OEXv5Rww0iw2i3m+F
ZxuHcQQhOkM+H8etwsYUlxP7KUcknRDilGTYPTgPgxUvp0v+vMwZt7mnxlz+CgX6
v67L1W24FTJuQZtVQq2lj/u7m9aC32Any+CIz1D8GXgvYIiCNfk6+cS1N1adECn+
MpktqwVgGplaNgNYkDX+i2xPj2gChGwdNAyyekwEtIKh1TR+4m9o1pVPWWiFmqqq
BSMm3UCd7Srs7nwHnCmfbw/CpZPrpuLAkeTSWmEHPVXQaijuHDfEp1ObdkEVkNrU
JapRV6m5QRRByA6+Wzf8Q8H82e1qQ63fLGcrcyKc49nwFaFDxDF/3Fs3A/ZIisMk
u/fn3HZcEWuHqVnOOgaG0Iqs1ykTtCeRdoPIzhGapM2YNeEFLh/QUpneN3KkO35k
JpW1G8TJls4fZE7BoCRz1JkiQaVWUWel5oGBNG1UYd7xzblH3VJMbkjyfXKeffXb
Mi1bvPxPZhmChjxhQrFpic2ptMdrQSL5Dp2J3CNJtgYBPA2Ac/X+mgwtuUq4akTL
VGAnWyk5RmwrKK8kDZ+fCsym6SyTgrTMUIkjIC/9H49t9CLWw3ckfQ8SUMcZwNUv
tCQHfQOgxBsvzt/FaC+dfCs++KY8voudQV2ebX+JVzAniNJpqtMFw+tSymPqLc/v
Isn8FCFdqap6xEHxBz0SWubaoJ04GbPW0VbFWkEJpfoet+IZuPGXgWXMmiPoGdtJ
GLDWrwnN8Z6UTUwM3oHwn6daYTPH5e84mobe8cUSYxBNXCP9r/esLAsrh9oq//De
HDPYKj+qM3WjVluziyQc83+kZQIHwMVjnaTXv3DeeDPJQjc5PISvWFHaB1yOiLsb
fz4lTvZVrCmU3PdAVB1N3RQ+PXeNlAOTTVX2GviNpjswuBtSyoF7dnT4Po0wNiOe
QbP2tkA04g0KsU9IMWzFN7njP8oxmmm33eRpU5hRCDd6B6ZSfnUtlh+Mp6KoCipG
76o4kKRHtekXhzbg6fgLt6zehzyem1cP7UsMuvJvzPmdog4Mlvikstdn1ccRTNQg
NM9UEv+JlRWwe+twPUgXSqDdg3vCYI+S1GUmY5Ew3RXk/UX2KAJSYT9f6H8kyPIt
JG7CWYCVkvsg9WVOhwSfkIUfFCGYDzLGzpjF65cmxY2WNnAjV+UIT/vUbnQxLXt7
52oOUXb0ceivZlYBPRIqgdJUK6BgjcVAP5YcUhlPK/drCTDnpxPC+JKx5NpEO+nS
1q5NuHPMitGNHPGp6B3iUoZlpKclKDcQB7vC6W7nxzI24zslDzK3jtBn3lh1sOxR
RD9394SmJ7oeA19E4mc3BaPW9ordKW3cdkosNnBdr3FDGPxgsFISDmm/uD/U6O7J
t3dh38/nsT10QLoT/nE7+n3LG1sul6XUBVVdw01vcY5yJH6RwcUiRqeVqyWakJsD
+g3pJSAZ5+Dih0tA2pBTceoGVOlI0nOpZuuFx1Bo8XVrSNgso6QFVnmKY4uRKlPJ
WZAfhbOHEWWHhzgU0EXpcHrDqpgeGRDk8RJF8YJ44Lo9krhtyO7GV+an1eA63A96
Ff6068RvbXfE+p27/JnNUpbJE5yM/X3oemUJMoyDYDHUhYF1oC8Z5TDmf/Zr0dmX
RGX23tWIkCEoBqDiV+pCbq9wSjdOC4W8DB9DQtUrF13WUja4BzzmPVRwf/oLqVUB
FtOcMZyCdwhWs1vTVqxNwQBD/pN2apYiEZk1sI6Msm8o2gf4Y+ErlcHC1DJANyUf
8z1ONg+S4LjgHpuieBM5BGukgTiAZcYCtTxSrdVRxlR5H+hXbLrLdjrpxkJI+fQd
JvE4jj3QQmisyxJ2cxENj84g/Zxs/3WTirMDh7LcfKGRz7DExSkgowGibduHURLq
1frq7qNjfuJ3gWKgGEZYDXUaCPApBz9UIndU5WHCCCqbIlAEC+Q8CWLwppbfTrMy
2uTiDtn/WHdaP2Mzo1gnvQ==
`protect END_PROTECTED
