`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wCEVzRzc2oHBOaKflFJq1yyDqo4+tT/FV3FsZJ5hNWIEpbHsQesfgJjS45Olllk1
6psapw/eWSpXDS+GX2gbVbSK42ircjzIIrQJBwoeLlSCZxo9QL+ItU4JSRW746C5
XAd6L5STZDRmRizKZ5vgpmglfYaG+zjGICLP2fB9WZHpLjkQRDIji7TfT0C3HY3X
gT08QxV2BvUu0i3rNa1sziKrpz5zYbi3WXYWbk7lhmanNmJ5mx6RieWi9yE36dQr
/WPm+rPJQ3XHUueWRO6eVyXh4gZqtlXMnQhlRSSMH3MLJG9MF3ndWq8hO22NhKan
zPnLTlzhq29xDYtNiay9ks22/hn4uBP9eCWalgE4LPjXNVMsImUyM8JEPOJyRauG
UXh2fBuMaDP9t9f+wVG+H1PDejRGngfna841buuX9DjHkV78xH3lpQTbBxKSU6pL
Hgbtl0g1dv9qnGh0F9Jy0RS2BYyHz/5e8vch42URaC0HUEUJw5xjy8QM0Wbmtko3
Y7C4scHeq/sSfhFrfF5G7edRE85h9r7GuNdax826hA1fsrburguKgj5IiKUYNNCd
mS3cpUCh23jZxBeEhb4zT5wsMAzyI4TBGyNi/dYIDWIGgUAXwkLDhV4O4FO4orWu
Z9lEUbRJpyCPAky31TrThivMPz6EEufK3IjJAeVzb0rP141gQ2VhATvYXqE3WOYj
fbwaHuDbfUd9yxx9SqVHuB7U/llgyBQRlwuEI29CRnMxxCU0G0/gYNhjVrPP1qBH
EwEXOqZbimOCOzpYxJG/UJ4pNA/aBr0iLj7YB/pjwpTtTHWi01myBJh/jn1T42+D
roMltJv+u2ClkESfsh+3bPrrJfCIeiizGBkhp5k201Wnt8D75RV/X21KNBoe7t7i
hOBpX1zNyJedRcq9JJ/oCTGHq4wy104lZK3U1lDjoR9/BSI1zNlJRld3+NXuysRm
aRqz9WngIuF7hlCUPC/zSDyYGwX5X0FcWXTCX6YV2bZXy1Jy5Gju9JCQiA3MzOX6
FUgRADW2WE4Ru/rgPg/pIgS7p/wYe7cxTZVArWE4ZFmOFAoeUkp+V25nd/sb4I4C
QnTk6Ki6M+6rQQVTMYPUv2cufEU6j61iHX3jOWGn8ryOfp5AWwfmzNNR6oEBRlf/
yuL4JAG9SAuzm6ITmSlF8WZFyTho6674uF43eAMXiBH40caKXG35tcVFvCccFrLa
0EDu0wgObvxQ/ZHapXCPiDnGeZqe0JrzhAzXjS+vb9RoAp0Fqu8A3P+hGXQUEcWY
iiD36D9Sy0d+qDd/p9dXt35UE82JATfy22OlG646yTTyaKlg1Jc2C8ns+B96s0F1
C6wKlHj9iODilfY1bx3mITg8tt+t1Qw8Ts2Oj6tRk5tQRFc0qZbNIOyPO5YFw2rt
THiaGj1rTe6Eu6bPfb9BL+lj8ZaD1DOrnLz0TDVixFbYYSwrnzGiciQO/LsNKSYI
mJHKnak1lGNObbdyE6NQRbVrDR1Rr1vN7Wm3YLuAlxxDiuQhNbM+dTmkW3GfdeWk
0eehuXaGkpW2a5xG8bJeVZcYJc4i1V/C5s4+XE3ix1nVHF8dSHSl1nV1T3O4JIMP
CBW6pvKbwZvMzDUnyJTgNnSYEomIjMnKtip5zwFYUOO3qb2ECSILF3b7Ar/U1uF2
Jcco/4Mm/6ZbWP6ViMFNC/iuTN+tiLPDhLUjsFA55z10iPQFEkmD3iMlM7PJZ0Gh
do0yAztRVfv/K10RZBVXKfwsCkKqRYjurzcBZaSXK/6eRQEmWW1Rx2svS9aj4a03
D21ecIUjjLssuyQBoRL7OV8P7N+TdJTM9/s7XMtYsP/vyoNM3KY6td+HhythHetz
nrdFuY5BbObeZ21j17PbUN7IvElG91X1y5kUaG77iki+daj+bEXS/9nWruiENSTP
s5xl+521KxNFSuu5qe8P8zbptNYOyFpJFtgB/LuJxiXUrOSFVAgzrC1333HZPctU
LZcLnSUvtdgnMEXLcw6528IDKrfLix/qrsxpOPf9LqZRNe2EdKkQMy2An6gUVQxZ
edASBkYSY29rFj17Cfw+AyMjQFsmOb++Gagi8TGLKA+8xUwxxljqjx3xYaJlbqzU
crUAwVcyU7yhCZOzQM+p2+WGMVvkZOjm5oXtd++tYLYANIhTfNwjOpNyn8ue4baB
qwAeMS1KWSzc/gmrAH5HHo0xSq2D0DX7zzSpEb+OB9czHNuYfh+qFfhT6eDZGqcx
X3HzGQ0OlbylxdnBYi1Da4QeGgPX2Zi2nDQ+SC7CX5ZjPd/RDvJ9HZ7mA+fV1FLw
rT2ts1thm0CCHNZSt6Kjn+yYwBDisqclPopAuYm54HU3f3QFcNMcWfUcG/it4snJ
a4ZdRntGfafaMHn1S82nThIz1TEzajLWh7h+24r9TWumFDtu5Q/VeiNeuOh5gSbL
MvUgPwqa50NbIAdnj9SQYm03SHmC0QxcQD08iqAJSZdtAAldVX0/B47vVOYEk0bC
nnUO5y4ud7MHe0fnrqHHF2b8wQ8SlT2rUBmPGIDXrWg279RMyMsuK0YxwdkcRuhW
q+9OnXWsPQVTtEq9VI/XtnXa4JQnCZBBfOvO7pgpIV3FPGCifHlvXwTDOJQL4O41
9PerRqatUoNZCXWY2N1yTR0kwOa8bo73Ta4sUDSxs0uJcjoUo4dohrydlVrpizDZ
8msb4NdmS5ZcAVhDFh1tu4HI7ly8ZwyXg950ilyHdC2gQfnsMMJeXX61JX7ncRES
Q/oLk2A3kohqO2Np6lZPvR7ZXJa/4eMuyqn7SaTTeRMQT/MXFy+cnRF+Dkmb2xfS
ptbvOI/n/E5BCKzaJ85PynRPTia4wu3Y+wjmqvezjfhRWaoU3cJmb3FwhBf20gYW
z8dnhPBsNqnwAbCuJy9lyPqNc+4oaccFM6MFnMabt6D+XUGpcApVnX9Urj/JNTiD
+1pBvfr8OKndCuGv3xpGszaX5uFsWj9OF2d2FLS6KOi69By65PJToF43cQeOd6fX
QM6zDU/DREBpOqbE1H10rLHOdPXJPjaEsKqGTPhCB/Uix/NiiWbXbb4/n2FqbUEB
veQNPuTvVn6vOq/9cX0F9/uGNnn7yfx3J/wlVEVdQuJJYY3guZGZzXDJf+pW6942
/SKxdLa0CEqwHqj4LHhF04YuiUUoDQ1YJ5PPevyR651+NE/mPgi3cadSd7l5GWMR
ogzUf/vDPpmtgyTiJCk44NkFfYrhc6i1t1qLGX6q0fysp7KrYvRcvYPMq3pGS4qn
bKOP4tEbEfWsms/Q3J3KC0UhOh3vbmVLK1hhw4H/nAZNXPIjH/vR+xzkzWkLo0ZT
VERoirD5KFW2N8yK7pi79eiSlaRlBo7hp6dfJx12Y2LoHPuP9gxCj+RWukFhqsld
JcIP/2b2KvdPoB0v0LENXvJ4ucGPL9Q+aYAl1/sy3Bv6tAVOo6XKuEoV84sxjTLc
CPBrMxyR4EwAYDnX9FTM+U4j5ZIpuecyqewrO5VcAxxN7mF7ptNFxwX8fLKjp++/
mYXmg7Qx1Sae09YWP2/DmXmN7iImQmYaoI2vIuqGpLpKZuko0irqDHMRvudXVWE0
4G/UnZUWA244Wo9/tCxOd3j90lK+8AhgRBJZKn5toYBxfUjUxoBC8uthXEB1P3ZQ
Kqa6rv83HW8TVZOpfscnnaa0Vx3aYFUFStLFuh2zXPETmiNymWXCFrgFa7gK0yNx
cTZILuHbLajpzyv/ozfhEoDl79zunDDniLpsMi+zSNZvyI4WWamkkPEEGDSrXmE2
l/hF4Jqq7K7KVmZqXfKSx3NPwLd2zOCL8/HAWjorcwUzBhXn+jjUVkonusX+yNu/
tUqNyFR53Hkn1LH4n55RqTOjPHuQ8Iw4xjpGH+INU62oRsYty0efrf92KVx5qlbz
TgHpmwwFBnVUJpKSDnXORXyIqw69Z4zC+Ku4i2KKv++RiK+qMVrFfTmnOS4C2/Vx
8dRV1wA8ePrBGsOPGyFqvh75VFkwGLf6ESwA2VS6rcux8e5M/jJNSRYwPGBQ/mga
Bdz/wsTz0y+KMDgMwTliAr1HXmW9CaDz3auI461Q18xvNMembrjoZzfSnh6+TNa3
vUa0xTiQ383pTqVvbB0xetDSNN8BS42qv7bOlQUtbAaXRuBbRWxFm8wXscBQqCwW
2wYkr2OuBe+k2KDimdWfTO2f0zvDciWXck9qdVdzyKJNCNAMcVZKglI7e/ulSe63
eLJn7whaoH+qMHG+rvAzglmejTOm3tD15HcUF65J5o1kUqbb2V//BnTDsGcng3mj
M6jukqTt5dGc0wEa/Q/jYCbzd1faEZGtBN9KYe8Zkov/wJZ2NAoX+K5FVQO2sOp0
/i8a2c6RwOwGuVlSiLhzDEGD/hGIEf9ZIsHYFZ9F674GkOoylu1m/eOIT0xTSTgH
1pJ0a9czPBp4IfWQt0LG6EATW0/Iw9PtvHsbfVjxyPnFGKwGQae0eY9t68CPjk9Z
/VyhRi8+orkFZl/g7ax10s7QoAXG/S/5HST6yB72qqoiQKXAsCEuwhe1ivcOoDDB
s40UOGQ4czMN/M3WLp8PfyFabjZf9lGZQ3omewPjwHwvSl6+oeAhzP7jZgcLLACd
EYt6vh3v0QEfMEmowaH9+Zy6jktNDjok2EnkV09RyCwq8YdedGQO9BoLQ376li88
/NNmeqN66dPx5hsTW/0YKU4YVgHChe1P9gOlAo394pbScj3MAh1vDrlKtvUXAQpH
+ce1ekw+5Iz7gPNYB2rGWk+Xi8ILZy4qRl0O68Mq9cuUodT2flVKI5Fv09Nbeo5h
h5QxintTTLnq3yEEIPPOw2KO4eUYdjDAlif3acIleQpXP1ADN8cMKc1GVT1FgqCU
7gXJd7XBos1DH2gMX5AYHlRqMHWk3mVpfmpDJMfAIiXqHwFa4pTNDW+Q0SNBySeG
KTFEA8+YriRPGHDwqfUcZIgixnWR9Zouy8DF1Jn69ju4bRMlABYO3ct3xk7X9I4i
jvdnGOCXO+64VsCyae4xIieMex5XH3D61lKO7/EuZF7qbmPoPPBMM1jRpZ6JpDtb
p44DHRPtBeBDc6P7FWCPEhqBd8qrkvkkusbLejYNOosrVXwd6CdxjZejUEfNrRxd
TZkivq2UsdMea9w1VNN/VBIHHsAwlsnDQvp4cob36kGnQs84WeDsYuER6qU54v+8
Vb7PadzWV8qMpzCo6USLbUE6vZcw3vgXMVpUY3Anb1MmtjNNhwGHxmYIrEBw8c4E
WNpIQBU5XFdHXWIFpBTmk+yDEsVHuoxuQQN/aRJaU9PMfkW6lYLsSUUQSh6qJP7B
PGAyKu3mYlHZvIaJN+S5KPs0YlkApa41IzmjCZMdxJLNhqjUmCmZ+7jsNJFkzDmd
aH0oK9m73U+7+VHGEmoFQefZ411KRnOHVJ1LGF4CpJcF3+8Q0gWErOFo9OfumFMo
ueW4P1fIGpLXyIFomkNMtns5Z4Y/YkypXUgbE1Pzg5iKp98fNjDsbPZ/5e0shzDg
5wU94j9LDsBSSDtqulVa9jngi5rxJWqDyk6QtRL5QcsRspfreY69dQjRT5F22dvk
wh0Emz8Kpg0SrH/XdDcGycc3wanuNy267PmW1HtDde2FAdPtfDFSpYQB19D8ifkU
FAusapbdvPPVt3u4kDDcla8tQfPJgUt27L6yQzWXD52N6hu7sE/BoweKHPcPBKtF
mf1TglJFceeFAYBt7hUZWe+0t1fHIxRksenWx0U0bYs8PEdwljpbpsEBMq10nyr8
DQIk053wEvZtP/vL+VNy400gGK10Z9pz4z65MepLr3ExZ49eCHZ1QcafjrNppgaA
WrAKTtf7AF+UPy3BrJbSox8lPOocHo6ZycnzC8y6qOcYnZRntAq3LwWFozsU35md
yjqK8rpBVtlWSRIKJxO6nFfI3FHls4gos5oCJnsYmMTqH7nh4nS9cwQr/QOBfJyk
SV8usTcGJPYwj+sWeYKFkFNDofMH86O8TPEjXzMjenU=
`protect END_PROTECTED
