`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/FauH6rUFGYAjc1F8qaIqfVntLhtGoFp8Mz2iYMaaDbklv1JEC34o9ASP+2FIbk
xF6Oh5Iaz/HVzHtVT04W1WkuNMj9Oge5X9UVO0Nleo5vV75ZVItGIcqV2z+K8+Xz
u02gquiOEoozkMpcU/FcCX8a6ueg63gqgzg/qnfwTpXa0EE/+CAurRxBp0jm+hln
MKHNOhblfyNp+J8HfJxzlBkwNALnJCKPMwYWrIRyUYRmQ+ui6P9eyRKeRYAuE8go
jMTHkUctj9RT0F4Xm9u4klc+aSHRvIOIMvcCRh+Fsui9F2MERXVqvgccCn/jkMr5
o/dfFd/Zx8K6pJui7L1xwklPXJfnZHsjZ7+95lAfw+FLaRTpWgs8zn94R3Z896Ab
Rci5IxncgYukuwS3EuH8f7fda3cwbwDTHe2b4zq29J/OHZo7WjQeY2VfeVu2mEby
ZHzvxyvfW0UoRL2wyyBQNjsb7MlNyA8uQKS48ft7RL+tT9tP4qjiwRBFPv4ByldJ
UrBKVO4Avc4aqfkW7yZVzBqpJBCiePy+x5rTtlQqxQtbjlN7e27iAS/8GFj8Qr+G
8dgPuVgWofO0Dy2JlD28G7rOpKm5x7nFKIa1FSA7JEnoC62a/4RpjN0Rh5e9wMQe
0crrN2B/2IOHG7+lky0TFjmPoU2iQ0r0HMvVEEqPjWfL3lJauJEQoQN9BtN4Grvb
7SwOEWYyFte+FNHENWcqSxyda3qMWjmrQuwFLOm4S1L59cCC1eGlX1oqgEGBFxz6
o68gIQPXzPXhAaaNoyE/W633gioYDDH7u6J34+v6PrrbEepFOB9NYHmgpuXmXUnR
33ltXOru5SsGFmQt9EYQGBk3OKmhFTJENghi2quXx9M3NCzVRPVqxO+s2GunUJqW
J37kMx/T1vbdvSN4FJwo6CxQeFHsyvJwoY3vXPwOP/3bJHb5zCyvnvyAhqsy0OBM
NJYrFsh2Vq8cSrij5Ayfhg61qFY59Idzo96rhRmatrPDlHGWlRsE91Y7Vgu8ASzG
SNiqNJJrtBnzgCL+TboX6Q3tiksgjq2wO4xfYnfS1VFfIo90l6OQcjz1WAEVZ1Sq
aJjHKE59FXVplTfTJJ0bpot7KWYXyqTwSYczS9YznsLEqphQ286yT9zdW9/jSxXY
HSRAnjoqGkL0p2EfnXnlGHayrDlFCP++OPtNFr+kblZMLWXWLUJzEbDZXN8ayq7Y
LM16n/6huYhah7oO1TrAAs+8wpFTII+Z/YB3Wm2CRFW9aDTVHY/JSkyWS5wf/aVG
GBHjJRdoZnULn6Q7OhiKFqEKK32LHoX1snn7sTI+CcsbNvY6SE+cMCSEdS445u7i
jyBn2iJ9CIwWlhnaSDPyVzs6OYKysrISAe4iqHrtMZg0JCiDVusyOEYEmF8637Ac
fRQbOv6v/1b6kOQEp4l3jAX32JkVyqZ7UX288O8o5YYXyg02tP4yswiojxWzlJrk
0Xsa9qE5NPH+aCQNOUEXHhdIeBtd9g4U5iZii2Yva0+6fW/d+7tiAQUZkl59W24Z
0W1NMYjwbpqY1YUbhbVzmDr+o6u7h3+2cDaqgt1bjdTSxKCmCaBJxB9hDZB+GWkq
3JxnsSBHDXtF0fdVsBxB/6GyUJVOOdzJ6Ktt55l7YnhGGsu8zddcgdVRUxgNPOsZ
qMhfmZQ7/gTjYyU3rJjP3HIcq0QXgIVdffD/F1+wKa/gQJJr7Gjo+AjL8v9Org6i
pnDaKmCkJNKffsFeycyHEy/0Jw9PZ9BRd6LFu3FbKvvQmqeAI1iTxpwvKp9M5XFG
/OwqSEL0c6bHuj0L2APaWQRSzq/s+lmSZ/PoWMDK/+pTbhFOFoydMLaZQV3oIDik
Hcdevv4yE/WnKj9gewS96YqCY7aDAV8GZwtnfTK2+oq/7Vo7YKa+rz3Cc6JzLWls
C86gjnIMMUA0hCXnq3W8gZ7NeMjsNMSFC/CFwRVOT4U56Irt3bUxjk0025LRqIRy
XfNmpYD8BAP/NsnW4I+D05+eHjfgsAY71y8JZ8CBeIqzJZoyKIsqyVCXKEOH6pi6
i3BnCHtX3j30NxTW+M7zru7QkW5PBJdvCIXaBD5UtDu/fIFkoUOGlUlXC+ttIprh
fUK24JTYweqpYF5hbLsDqBoN1RxQDhJWPO91ypM4dGJquqcx/NVEpP8HIcHrimJb
IbTiYDNt/5gKiOt6A5tTk1f+c35dB89SatLdlT79SQX6hnrn8CjSTNV4A4knx6pc
KnUbuOXGisMJEVr4d3PZ7Q7LG0j9wE3gyv49rlPwbVMgphM95CsISgTHf5y9dwnZ
BhRVKSLQHz6z1hpK5RS0p+Y1S8FgzwwUwG58UFlBmxD9BHfkWZ0AiLX2VHLNlijx
RJTKArWDEIMf+HeO/pKI4SLw564u8AlRMyrrJT92HzZdyueZ3VNppPuBvjaPvKvw
Bnqf4hONS51WVYLy5BFtop4OYeEtwbhia94X/GTLx0yFztQxAs1xxDqogt6OxqbE
yep8hxnWYvMxBdwBk6rCI2gjZ70obSKuHit3E5GgcV53X758SPHt8ivLnf6l+QDi
eCpf1g5o3VNi2lH6ZTatyoD+zn+5LpUjzcpWIRg9cxxEHVsCEKRnwmVFmIg2b0vy
1k6nSqYcV9EciE6KGhuYy6BzTJ4dvvPBQxab4cznQ/3C5JMbMZvMZtUGiQpwuNh/
ZJZwP6D686SB8Q+GcYoOG+yEG6yRPM12I3Qz+b9iIYoIvDG2LeBPZf+tQUOoIbXP
n9NhdfebMR4LiSpip6Pg/Wpf0+5zRmxS09DhsyNSRzveYy97q+bVP3e2v3KviXjH
8t7v07nrWK4v4yunkchfiGAg9xwNkJe3nBzJm8TMgThwm2416jTntgZrLP2WL81e
OhRHMUNd/UhUeAdw5Av4wCHrS8kgM1mPmnBhF/IaVf8G7WpX6DAOV+TP83ZGvvAR
9VrIOtCyeMriQh0b8WX2SvWm08zKJwZQUtKqr37S8OEwZgmsT7DQthVPxOeQkZEu
dD1TgJOIgatFFPFDKPwPZrd0IVgwhZ/0AHSS86yi20EfKF4RrYnBU+3pAUYKKxXG
M6ftXO1BYA5k0fKfi9WeIbMpCvqJ+beMt4sTCHGv9xfAiqq0rOtuzLgdeLD/xvpF
K2ZcLOn/xC1f2PMlmAXoq5RDrnwLJtfE65q3SIBxXL+vpBxEIxlc/GuKOeSJz1AZ
QmlQet4aWdvweCqGpssSEnjB8szylQivfIFHR75rlok5Gnh9LQ1dPBvtey8INv8M
UkTnujbJ2VMgFtZGOydDxtrS4y8j0iL3G+ngWDIM76i+IUCI6SzL8QIt9YV4ukC4
dmgqiFEwZFP/+Ian5CmAzxnfSbrcL/uQgU9O6ipmU4PNZ4LUifDmfMQ7dJD70DOS
QKPZv5anBv9oeSmLmoIBSm2OLG4m1zau/r8iq4vMyC7KPMAf+PRxdmB7/tp84PlA
2Pt1ou/8l62pzt0Zmb6sqh03NUDbEk0On6oxmcAkfxXXbNp99rLYqG0Yht/TPuA1
txA2v6TmHMUJH5GS4jREtEWGXCa/oe/ZAlNeuPEWAbS1wmwvIIl6Y093OrXbdNBv
cu9NPQJqad5kUKXFa/EdIWS3PBo6A24Z36KzBiDLZvSF2VaMtfA6LguH4VBl58dA
RVJa2a6ghMz4WmVF4QTF/ZKdyD4kVT/YmyIBdFDOV/R4dH+UBkVyEY7MWYPKAaJd
DHC8Uge0JkrxoBoN4eIEkHzn3ZV14I6D5LQC7RHCuaRAoI1FHe9ejHIYCM7VYikx
l2LyYrPnp6nvfI05OH8NZgQGIvAsHiw50YBUvDU0WJ4WNIQmUj2qoQYc6li/BB6f
PYqQ2hVtiQigibcoTSKGdVNSq9hba4G92JW0YfPFZ1mzVMk8SuwJQmS8kqgb2GAx
m6qPoW0u2Juvu8UhQ+70X10FrpFgGoMZbyDbN6muoOlwq6m3rU7e0tgmqcE8FPw+
uFoWLrd6MWW5bFj5Tq0yC2qkpgLIQULMH0uk/GMoA/kgrK0/C1PTM7U3yMELFWHf
NUKR9NmQajrvmk+MMQp1p3VDH6ErcnXZuACZ9pjHMi8UR3CTs9++ku1xip0BBzjw
18U5Uo6wzZTyRjklVN6sIuh99zUltWWtTv7SXnowYErg4cEMoiq7eEcmeJwNZOl1
PpmjgA2tyIJfrCag8IShUmFrlsW88z+8FiuQgbURA1rbB3cClhR8B8crxCimVwqK
PP6VcSe6sipU0IkQouRsarRsYI4LIL5f8U4tbgtECkka/pHlez8Mpc1Y19hBrZam
odqltZC4gHfPIeNKr+I8Ib3bvUM77763g3TsAByH6XAsTzgnJOs/3Y3JrJe61eIo
eVc+AUd1Kc6qeqbYSd7/JgnJosIk3KiLDukNPwdjPyAV5Naj+GwgLuhb0aNyHma6
51RBKrN714DFlaO/RnpMBxioMcuWlrxMAtDFL2j8K2JqFN3CF1wDDtnJntK8sekm
gEJA2fvlyQLLpoAtCwjXFedeNE7bwyLQVoKk6t3T16eprECGrXwZWjbT27FJ/Bjw
US0YF0IOif7eUhNL06dLehUfQA4rbRm0YJHzlFDhsMRrWz3mybYwK2pyZuA0edv1
FGhT7XE68XMB62bEzH1QRiqg2JjZcG4IrYLvhLSyD92jiLNoj1IEgqBcJ5Os1g47
YuELXLQGICHmF0q4vKmCxMxEwNL9XGlJbPgUQBbfBDlvIt72MbsCY6vd9Z1KNBtj
C/G0o9vbrnfaqJkeeZGEm3gA5mshAaIGRHOzlFcjiQM3gGB8QYvD2KFJhrIzQeCP
TfvXNsUyg98qupT9vFp8ULQCbAKywGo+6/h0kutpjjsNZF/31kZ+ukcNSsCOuIAL
/3t4DaYgNI6L03XwQbFnZ+nJdhlDARTsoAGnoyaYXU2/cpfCN5aIDsSm0def9f2U
0gRyZakY/0x8JNvOMxsv37470K7bdMVgwZErxmMaPwv0nU4ORuh7kMcINJOuqhq4
bPhBL3D1hhIlnBTA797CmRlkRWrQNk+oxR1IB/3dVQD5hQ3ofSZMSbdZzli4DPNO
QRLeQqs4AyjvJ0ZtJcBtBuTSekxNgENCNVqPUJgPU42FcuM3dMkRQyQHv7yil0BN
1g6DnOuFbpAYj//GbmguKoaIbAW86dBs7wJdjR8tEueyHdsjh6uflK4poHXHyRE/
BR2Essr6RNKn/rueBxOEkjYx5hJM3RWRwJxZph96ucFvYcgFFhk5hMUbcYdp0+Lg
xlwp+e4I54mzACQU84PSpapEDAOM8JJlNm33PvBTpNorR0o0hSaIjKNRZ5beLQsd
nTlESwQq70DTrmfnxQfHB7v+3z7uG7b0+7/6Fi7wS3ckFRrI4B6d2A8kNnZR1VIt
1MZU6VYeFUn6uMY+/YfbjC8k4w7l94U0MupQlOdXPnFeRfCG/qseIsE9LvkXuEZZ
aQKgGrNL5Ma0FvtAIX6CeOJRWRFGXg7m8NgPYVaAIvLSWI4Ugfmn7ULpXKZKximH
L7ChAa4cdFwnC2Fxw9AKwphe5Af37NfV0eg+b6Gfpng6IvO0+7pSQETWl6ZrdXDe
zWDRGDXYOVvA0Fb/WnsJcVBUH1DTYYDc3FcGqDQkrndMmNGKV656SUliIFOn9QUE
StdJqleCz64XjqM8yGRT0c5LCmTxuUDSuC3RjPnFrRUWyEVojsoPShGKOl8dFTmr
eGfVhwv9LE1BcFk/GKZiMzBhQtJn6/Qxai4eIEYTaZrLv3VHxvvGf2SepxoJvXDf
WVqthzjT+WaK7evnuJwP/lc7bQkccEmiK6i2erOn4S3eOGOT2YP20AcgXLrraYkJ
VTOjaUzgwHgT9h4khlMzAYOSJFBqIhefmdnu9SDx1c0b8p2xwlM/xC6j7l2QY0dm
jt560BSN0yTpCzScJT4+D7kA05AQpKOFXUnRLSGzIBgpRkMPWzwrUBDT9tDI6DeJ
tO8vjW2VRBcRvQ4vmeuRWz61zHmpV2NEsSAZevhDWBBrYUh0zRdKaI+9zvraCcpy
e+bSNcBGN2luha4Ov5vws2E4B8BHap/60Rr/sO5FprLC5dAhZv9MxYyQ8n7sKCsK
ZW1lZDqmsiBaFmXtrh6t14cUpgAMmQWEExFb7x3tdxwg32CIYH4WKZe71pOwJms2
YXstyaSfoMGjlUu5qwd82FfDsXSCc4hfU0TtThR4UyyWbrR/KOV9+o1Lvcoh5KXu
daj8kMTh/i4pxV0yeYu7k8JBzxMrs3gUL2umqqslTcYsAkvNkKGN/0LoCxu4no22
mea7rG1eyyXyi7C1ZTha7ueQSGmpcz56s7ALqgn+BiYtN96bS3g5KXl3yugl3Q31
zPqNl9hhk8qc5DjxNbsAkaFMtvGnxhV2aJu0ZJhO5gPTFaQy915JT/ngp0AHSyYu
EYQgIt8fl2QZpgLEbZWI2t+DHwPXSSyPFJU64u5JWt897YCKVELW6jzZLasN9sQW
hnRRMCSzSeWGyu6G+8C5MVD33oTIpNvSebAdoq85zIzk0/w0Ts3bcWXU9VvpldN9
mVB9gihahSfhDFxv+aisUg35w1kVclBCACLtc6W/V7BKu5Qxsljec8T/TmXHkw2t
1KwCyZStX+oEN8HXG6u6UOFQFzjL8W6JxXvKpFsjlc/6xsXWphXaI4WaNk6ytMQC
KyStR9Yz3SXUjP2f5wdGkKEHa3p2HMQYWMezBVmll3BR/9rxxd0CLao3e/YbqLgn
6On/InPePU8likLjW4/DLDb0H0TtjNweJ/3U/cMmr2E2uF373P7tuM50oqAHyqEX
5WLWFpACkWeKq6WU+Ja0DYPkk8HgDovxSXvA2LYNIyQEFwgDvKKdeJpK8JTm4MT8
iGoHRp1WPPaeRLQa0EUM3AtKl+bU9ugs4oLiGua1X2qgMArf4CA7fQvAycaoQehT
QwLS6drYjhzIowyeGQCFhUnjlTrLmpEw9BUuiPw7ZUZDmEPQtYykSViQb+S60Gza
L18m3FCPerlX+S1D/rQ1URqtedA8APRFKKCFy+cR8iq5Pw7bFjudmeIFlV4wdSEx
IvHS3oo2gZRadIhOsYr+6C+eJUa07ywcYm4JWqbMW7M8VcfKEcT9TfU3QLDMtR+M
29ByFjonCmkZrsCQcbhaTeY68/i2YkBV5Ie/fD15i6SbX0o8uCvFi2C5VJph1pZ7
CAIiZGybrHhlZy107xYqOkaXDbsp7N++OblQ6T3iTmZ3ZaFYtFwcOydr1KTBJeQZ
cAJM/JNsibpTkz/8ubdffPkveRY8TyhZAQaiNfUl2nHJST3Gyf7h8HANlq+zM6ZA
rMIPtfqXvrNEe9aE1KuVgqjC1OcfBQFL2ge7P6eNeJGPIBG5jZaWhlZ9szLlhZDQ
rb39QPLdVkloqG648ZpWttbUVAKRM9loFV2VGS9FmvYHbBuH/ms7DKzFHB+xTZrP
afNTkn7WdyaxYG1xmFNdasrYE3gKgvejDDNzT7gCnVLQCxVv56K1T/qm1SqX2rpM
1gGQWjlZ5BYja4jz9BcsQB2zPdKhCA90ylcJrD2NGV5H9e4uaQYzHVnD/UUV/E6Z
tLpf4t4GTEZ27Bnqg5jeh8Bjju2JFYcnq0ceG9dlkRxcuDd/5HCV4tJTD7IKDoWw
t+m98j6f/3WwzmCMYv1I0AABWWLToPIGp/CgGYQUWwXcj9oR2Wq9ECyCSBcr6xKa
uUTLfXzPEZICEfayt94x+p2tQaYGayC35plU3qTzYD84KR+v+F3K4+qi3maY3Q8g
ZokUIVxfmhYIt9YkWhyxVw4klbShpPPqVfJO+yw2LAv4rtVG2DMc1bfr7Vy70nWm
v3CDTfJzxXSYVjvd7jR8IrnWQ8VlN19ClKm2qDRtCnaiO3GtLZx2YmOyMk9q3KxL
iSBeqfMPWyGJd5IRc4WagOaK8Bf6Fg99e1wFnTCY2rqmYBz49uWOHI/4FWkxzYLg
6m0lH1vzrHrWBqKj5D0h1rGgNVlAmRLDBNYLej0CBCxq8r2FYX+Q4dH5MHPYE25Z
SM2lUSbdsoYFoW7S4vrybLQsybnhnr+FCrKNI5cB2XYHNIjLyKzmszvjGxoTrgqL
V0SEqNj1mixcbeGTAq0U74kGj1BYWBgJTQQWi78hMitXg1UHp/oqq1PUW8+1a3r3
HkXpkCBEK8ZcHYBt9O22tO3rzx6fwigksxVBjoUe5ywYRzaVciHnqkXF3xYuCsXw
b46wNgOTekXnZsq+YsrM6tZ4++CaiI09z/OVga2DT29grFMArjuZ10o1YzdWNls3
FtPUWxrvxXEklga1/a5WUlocLB4pDN593aklrdjJ6wS52L5OmEXtwRGb3jU2NUHn
Qo7tI2vLNte7MStkO780ZTxyL89xWioaX85cULBF5qOkT8t7T/C58uTQ5PKNJngj
Bpo70kOgpr0FmoEPdUmI1XCCk8jtr26tO4E8WJGVnN8xODrL+dw01xTi7rajYNAx
UfSDBnVKPahOKJr1VJTyMcp9LSzRpJowHfpFiaiahJirldZc9DJVPwxe9JbGiLeb
rtVV5e+W3DI/9xwU4+oSbj+bIaaueIKGmYVM+THkja4o7CEDGFSSzY1RoU+/6y7u
AtWZk7V4zEZY+FiWob7Y3xniEyJr/SGjjednJvFD4iMbSlNgitxpd/93Zjum6G2R
fJ6Q5wCJ3UsSIxG3gweR7Qd7flY1o3V2bJ1QB5ghvGvi6aEgUbqBXEtgzfAEiS6F
+O6Bz2izkwCmEB+VNHKzkzfb8IJq8CyYoEKF5aixzIThHO96Q2nXgYGjvPUAoN7d
NCN9Jol348Plpvb2oqTwNUHLE5vpv0fUKQDdPwSzjTzvg19iMiz/08uo3OBR+L/B
ZcncKJIvmihyq2o9Zy43ShtUQ9V+YdwTA3EYBS+f4qXPCw0I6R/9lgf91oM7KjKs
ekT6QIyDVPeFePuTAmYJDCSnOIzaJ6h7RxB4vtcivpsVM5r0w/YXAGDNunjwpTNC
uTWd6MH5IkNrCXOLSodD9u+US3H10d9hqs6mJ0d8l0tFrh6o6DgoEX7YAXp4EN8S
XtMhvrIJ4+Ul+PuAj/cX+wpQyxj9TooLCPo6HNvxHip8KG2qyyO7jp01AO9WXROE
KJ23dywq3gguVT1VyHPEXTqJsBYDoEzqLBDM1lUXWf2CrSA8M4acO4mXf9/GLH3m
UUGQgI3uhZiMA58h1i439Rt+yryaY7ade0Y3j82Ibb6DjTevGT/54DygkrI/mDAh
Tz2T/zHnD9N/+vYdFBpE0LEVISUajK0x74jpeKcccAmfZsn9g5NibaksV/g3eh3m
HcaJ1tWTRU5cH32gsYFSBC3PuQUjhBuRL9my3F14OKcTSzECkuR4dNWUIYYEVO99
f2lMK91JTPsN8FxdPmKdl4OrCPLw+D3yIPqVd2ncyPCy75tT+wclsUk9p/QEuV6h
bgj0quPz7Cz1srk2X1MOmllkhE194PjbICNOxZZ5VeqBBjCBLFFvL30hCWW7qCFd
sGHLFRb+KbyJMiqM7qEf0lwZEA7gujM2VeC8f2mOXNkxjB39dcpu5m8N+kP0mR4x
r+dSzxfxSl5zty276UNIDeAPCtD4wNS1JsCUcsOlazV3/g6r8GDZOJfzXrHACD1Y
Il3iQ9XQh7qAEQ0oZQx323VlGEl5fkknRWUrljFLSlkzQjJj4C24pXqT7+A3lVtd
4UQIgEXWah8gcHzHL71k/0G6fZj3sZmO9Ca7mIr5W1ynhf7WUujVE5TPDczQlkUp
mXy2bb4rbTdxNdWAc7wXZyVA8UMcz5MUsKdCEiGCjqgzDLUeVsVNXOfxbMFzFtI5
OinGNdOGcAys11DRzfErFKyMcCF95tlGYKGazRxs84/WeccDc3RQfboGGid1a0Xy
fEZxw4pjOvAcrx355JJmqdqoryLDZrBnq8/5sFiuL1tUw8eIuwq+MdFDqDkel4T7
S/HLzcdABUT5wUeyPBqNgGYAJxiP3VONU/+tfJqhVH2+zIq/OGYRkWvv0BPKHekv
4VHkkt25PLMhHTXIaLME1wWca7MoLEONPIz7X89gcPeTKNTFjneQq78wXUL6v/3m
H9fzL4PeGuPbrEIKJ6vnsNDIYsHhTzdrPOl5WXSLy0jQTg7sisN6qMIEQcSXgmF9
fitFmG4JXOaWH6swemCYDSFZ7M9BgScasVLorGO8GHJ7pRvxosJUN1RxUe4pAj6e
Q2/mHBM7425e77X28TY5kClzuj4lhqMd//XgLxMJZEQ4w5IgoDTG4asxXv0w8emm
UkO3pejF3gJfKAd9cp3PZJa/Js87i/f5TJXAkJrhyfmhCBFvSgmyzx7z7ZfddrjV
ApNnlOTSDhxGb2/q8JRJ3gl30Ly0l1bJqAtTK8/qGHwV5pYokBZOSDfcPNWCll7X
wNsevDmfd/coy8m6dayCWLAN7lyU4ToNhEI9xILxh0Ew/DgyAsnxmU8AeJJoyElz
sGEs2Ib/14x9he8e/31WCkHBw4UGzS0f8dfythcgH2T9pRPT88omjP9y0eZ/53Ya
WnSqcXsi0R8I2LwIZgBSq7JCAIshBzdlOcIV3kNQqDy6AF1763ssvIYoScyu8sNs
VTKvoJL0aE66K5viboKUnS6rBxWRQguseCqLuw+Vh2Z30QVmeXwhAD1TLtfJwUYr
XS05kE15yDoXUsp/ONRJg75UbXIPDqx25ZAa6jag1Z49sF28TCOEf/V1V87G8gAV
CcBvuK+PAVJKxhF0totVNmBxKFAv+OgTBJYPh5+zpy6tUqm06j3U6ZHMG1uDMqqM
nIfL7/aegvJnSczuWoNUmYfs5OVUw5lssGjSxpFpf+wUFsEKULI+jayOFWIuQVOY
JRNfoBXFmDpP3u+/yr0iGgUXN5mUsPC794IzHqwukjc2uZ4TsJ08dAD2J3rSVy34
8/8NVMKstOvZnPq1f0xug1Bg0A6TJvQ7rvr9TqHYoiU0RViwqpT86WCoUKeYyz0V
BRogxm5uCedkmW25eRNWwQhrx4mkeAn89QmX0ewbIlPwp7xkrPjpRm7NmE/YNDPG
HcMvPQcKegsX5kP6hS7VcrzyxhEt6wSC3nwYXVSIl5EjU4LS2z0u6wT76PEIXxP0
FmnSn8hg2IZEP/z1/rS7ntX/PKj3aEJByzFFSRG9PqBgNWzI9TLMvcY0k1HBJahJ
v9U9/xs+H63RSwyDLnyzYL8V45TincPQbfWJ03rxO9n/Z8u4f1Jl+RVUzO2phetP
Pw5TTupSwkaSjJxyetfSLBdvUUAHSTAvZyYAkx78gzhSU+//xPF9zFh4dCvWFak+
7T7/8mwzZXsYzKsUJwCk9xgvTTw3u0q16PIHSsFRWWvies0gdSsNWNQWEIfZqYa1
1fDsP7xTMgQ3/tPfoPNY08plSzexIBYaF2LNqf2MJt4kZm20RE4piJUC4GVoDmBc
xt2oe7rWXa1M2FqXp53hfPwlGSzvs9H+BDy4wS5OPTjBkMAJwxAg3hwjiiqarkfm
NhvmmeGO0wYgUX46WZLLJG2dkJXtgrt4S721EUSE/F0KD6150/FV6EYW4w/gNOCt
7mDZ+kAtGPp1GAiZNIMsDTU0I9VsNt9osjFsVYGcEMA7VGQjpkV23WXGZMTPMrhj
JfC/q9d1fBFpSCHyqwTFi0R3myTsb2haRo6K4e4p7WGSvqgWDPfw9iKYFrd4EzTh
dszkgsM+76Vb59Nl+ANGZ1+SkcrD7WfRzuQ7rU8pai8+gjRQmuE7XZx44X4FyrS2
BPfz1CMz34Iz2jRE3NfVODjotJYjZM9wIS49thd2HGDmmR97CokkiZD+W+XrPlbS
aY92gJGUy9a87IrDeqMqjqsKI/nFzp9LRGaMQDP6uwi962PeXxl90UPKbL+o2tOh
27X758y5Tm5YV0lh7xwwdXZ+3hc2/dxXUqSbZmT4yL0pJR+4iqldfi/OF0ammbOg
tKdnGgok20Oq17aRO5AS28YrGo6uKzFy0q6gdg15X/b+qwWUDa4WWpQhYJSVMdII
Oh4hJkeg1rrazNpp57ZPC6kaQ6Kz2+YGIc1u4H0Wrws4MAyRnDQzwSducbQkwyCA
jPMAVphkFGL6CjGkmxFVNlrtcACOVYjQ0ug7+97TJwEgXb5Qb6FOyB/5c4bO27lh
xBNEd3nNSg7augsMbl/vegUflJ/NUsz1n9N/4GJ4ZTZIXT0ESnZyzi7AcygMHL7W
evCqfV+Di6pu2jByFoZEPDOeFuKpMi36UhJ/mpJh4uptMNJ1a0pOFwgh4WBYnruh
rIyMDhhCYDW7WMgUKF8B8vzv0KLdtPI+mei6G3MsHxfs3bZac3R6zaNiF7rF2dbK
OVY34du/cJYWvLGcWk0ci8R+Zoz7ooHUfNeTbO2uMa4IpmXBO72ctMvyM62VJSyS
iTufB53AcJtkIbOBe7QCfSnxFtg+JAjv+nRjwAisw62RUW1NHJbtQsStsfEugnzd
3L/rTRURvqGmiiwnanpEV5ZvDrHwI6AsbBxI1wT2O0+d50JjVANtehN58+qPxnzR
pRKpNd0oY2aJ1Qq/L/zXBRGvc6h27/aHG10QwXW11Lg9yyGifReIUoJT91vbfJ1B
bmWLhICTi2t5al3fpQtl7DsBA5VWPnEhcoaD8tWe79ohdJx8bOSOjUjBy9N+Gdr7
nE2sqq9MWBbwczcr13+OyYuSMDtBDbcrdMpu3Am4MfF8jyddM4UFnHVubc7+00Au
F4ImUJzgBWLGBHODAkN7zKzDpCBAVd1aso5sigWeyVuXRsdQ539fcVllDIWQdYNR
B/SJr6DdORuMPQNSxZuei/LSetgEalWvyB1yKEU4jSVOEhCYiBuei+A4//S0HlFF
wqEpHzLIA93psYhB4Quqba2bgjoS5epC0mnV+PfVzmGYxz1XZFhAZ1V1SIG8z0jE
HEtDtPFJjUd5FDGjuiwzJBx1KCYE14pvA7bXOZhLJnLu4O0AfqyoO20pUzUaO07u
RF7RdNsb1E6muziJi7zYU1Hi0q5O9MXlrPkMjhh2erflMkAHHQSj1WvcjyNeukzH
m7APGYw0c8wNjApedpdfEsWbRpJHw9MEARfZyGU5qmyWoZ9GwByXe9rUpwSchbW9
jzVLZr4g71Llh2odA697otGctu+DSvHil8wV5UskX7gDcyhFuNlXijJY3GakB3zp
LnyMY2mc1REE3zZNaMaKuVa3EaUbC6VObTyjMAssmj0thrub3AEGyi8pTmEC106s
wVixwaf6QEPt8Aj9loLbq9F7j3RFEQTkUHs1mvxziKrDofK+0SK1jwnK/OVFWnLY
TlQQXZdceJTlFkftYuwAf3eQUa9kIz5QE5QDC9J+yd1RX7j8BvCBIo+HQ7R/kdzU
8gKklJzBw6ziXaW/yGw4dfq9MA09x/mFiRm/EyxYNYcNdP8gpffayyR5ALes3mVb
EwjLB4DLVVBOEYT+gC+xsimhWrSH/2WxV5CyE3oVLb4+DuqmZ6ynrjF5thqGmuC2
g/B2hvji05yQDCHkdKLGpGQs829nK9tcLQpk7cDfRJOSGSpqTqk9zu8d2wV3T7WY
CIJM5QvSHqWcEdaK6hqtKDCOxJ7P2hBUh0Qvy6zdOifFfL/N3wCZkjragYisvyIl
pLMyUkt17xvyzdVAfrkMK0puPfY94RsKeZHjxbjthx4XAqcVEmMm4u6PPtH0GySa
5D0mKHij6nH8JALMZuubLxvmUEb8DX6c+hpSt67ArTCDHjEzqNh/jysdz5UN0No+
/TbQ/n5lNPA7m2MmnC/z3MPCtMJmP0EiMyQBoj/uXevZhzGXv1c0yVS7h3rWSZPs
UFSDRCD7om/LFXnNYHgIh9WQjrxXXsz1vG8TrJiMwsw/nZ8u/AvSfwhwgIzikGzV
Cr/H686Snw5IwseUmgaYiKV48Bkt4HE8PDlBYdXhyq3vNg4ma+nl/FNFJYb06xIF
DgluG6IGxh9wP4+m2LsfiJrayt2YggpViTe/jKFC5xrpe2U62+fG63mIkQ/y96VG
b46PGdVZm0G46i7SPCEKZSHVr1hLU+j1DHfC/g43EpPt8EW138Hq6+PnE+2oXVaO
SI7pfbR2WQgnnQEHQxFM4wSYLpoey2x5mCICXBoe98rrLM5bb97tpifdY+9pKsqi
lUVR+RX6FvBl+sI+qNcu0OUTgIsGq5Dr7jeVquO58gVnCq0SePbBjlZkJh08wNy0
pAw5WurLSPSglxZwkmtbWg9i6Ld/PPELH5TL72GBr4+GiuDMvnhwicuOIRm1cKXP
zSwfk53LGB0s7mFriXM7SyChibwfinJs1p50hR9jdTHkcFdBQYG5G9UTfi4DJx69
772oUWkc9YvLOJJXDBQdkM3Qw9tTazVCDjCkjC4WbPY8PVQSSA+1OmJ2OPRe/ngW
M82mcbGEKKqt8TBNKRSB57hI73hPoJKrsrzIXSfkoBGLFGfcpA/PQwqQnOhdbWE4
F8Qeo3jmyNAhDgAs0xu/sKG2NNv03wuAsdR3lbQCZN5yUm2LRWvw1faNnI1tCfSG
SWk0Ye44yhHx5xJO7ILVJYlCRwxlrab31PoWW+6363R3t1ycqm3T7FwiA9+yZjfj
mRrulbunNNRPJVlmfCH+CCkivM0KKlG1HOGr1w+3dB+mY/TZA2x8fnDOUkT/8zlg
TxkKU00PJN2tVbw6O75i38Nt+siHDQv7uvQi9I7B1UQgBbz4p7q1eUhlGCSYnVu1
ukF6l+zLLq75OcE4MTDoF28Kl4UJWTJPOqqpCZUipUMPtO1H78KkK+iVhyJ92a4E
JtThFKrrSOouzvr524/rO0VW7BFwj958+hhh+WcNaXOp7kidIDs/ati7xz32WBp+
w0vvreKMXxEnKpHtYohE3lJtOUZshPa2CeSuenn78+BNmMqHLfNscvhzQDnKy84X
GOTDB4OCh7kTTxM7UfHWacdYbFMeG58gohMDfk3BXNNgFNxIXNB9+t+XobXKDlIo
NxC51dZ/3zNsAEu0ftK49orCzzz9tisweiK3CZKp7O8uF+RNkBq/yhe1rF1nej4M
JMLmd+joVymbZnZEiNo9y70OAsKHdc8gLWJ3GeK4ebheSS9JB6OTZSf9MtelAsEG
v4PKouZO5SfClb+kKSkKNOKLFG2VVq4cSNYWTHrHoFpzEMmQZ2vDo8TTrjJdAfpD
XvVjoZJOwctlCzYKRRmGWI42zkwmN0tYT6AAAExFdHNzUE3RnUTGnSHQciHjyBvf
yL67J6Es1G8sYCEmZUtoIIlBWnFHrCBuvgKN0kve+cezeeknOqglZdGpN0o23XKz
Kp8/nWKCNAyKPndHrEUwhs3E1hYpKz3bO6H92KyLtuVNUbnCj0LUv4zPSgJWc1Wa
y0LejS8P5iUseDo3eVdJgp3XpYXq2PbCP2K7nL5QLr9BEa37A+1LXfMlGy5qicZn
1g9Ou5y0U1ekQnSl58wxw3rdj3c/7l9zKfrPXeyjxX4eVpaaUSWqO8RTOzyseTag
8hDjKrSPZrKBqb21Q+lGsO7RWUzUggFZBekfCrnVep9IAI+bXL68ygPp03u21jUK
7lOFUnMUEZtHP6n3rrTFskTi0kbG69CkdmaThT0nZDnNuv2ysZaTJ3JbB0WcQ73H
JL2gyAiclIib+59irKDrwTusQ8f41IoZEzU8LJv4VuN/fXvs77GCxihZd6RBX9uQ
HXZKRZYNX4f/r0P9eb7Alelw/lE8MOxWs4kBhcswGrksJD6f4lNSNw8etoqUWlAT
Hy4fvyp/AWkLM1BR8aK1/Nyi1bXKd0cdl5ijFRr8I9W1oLcAHlwRmQmyPIzvOMnr
HVdXwvEz/D+uNyKS+mvxZADNakOCt+Z+8FPcBwR43dj0/ZYG3NiP7g4QqmfXdwVZ
gO46JYtAci7zcQaOKWGrVwouvxAVFdzU88gnQm/xSaNYAOQ5hr2dSqSI65/O+cVj
rZDMSP9FzVQkcHQ4yxhTBQReHInilR/448njM8jEjLKtL/ExieqmziLt3RCnV3ne
/Ol0J7VIs/c9H44L8BbpTl8W3Hos0D5KoknPhT2zy89kaoF5H8jxo914a5veK2CS
1Lf6pxiYWi8CGEzToFVbEGeswVj7wQonGB/foigAcwmMpVV/NunuBqUhqw2MMewe
PTLHHXSf3y6LhLKVqdfirNF7WgsgvShdfl6uqynoj+kxevsE8FYEtbAATCF65D4e
sjgCGRAB+RqmtO+C6UHD1EAkMNv1EfZBCw+CA360TVnsE4FjGLdNUYjiOty+o196
9HsYPCgE1KG+rRbW+M/AeYrh4F5vuXJvD9R6N+P1uXJzKtK0tPBGlIA+a3Q30oWF
g/k1qu4BMU2MbrImWJVj7yJNO3b5VS0DG3aerzGCigw0rfmy1Tyh5SKyUeVW2HHi
NI9x+lBgEaVBEXHT6CsO/5zDZqrV9BjMmImJF5oqf1AcqIZi1C9Tn8XbP6d7ehdA
ArATGCORQcr84RPHgtTYpYWbrCt9BVkr49wTSwW7MoZ3auH/l0olD8InSy0r0Nq1
7GJBOawGH+cULh3MfAH9xJmYjXsjsutmhYRUfVMlviC9E3BBnbze3Inafdt5/GYy
SMG4X+n8I0iqre6MVgFYOB4fDVBQd6D8+JuUPgi4LpVjHd1UPjouzrGoviBK/6RJ
2L2soGgIZTQk3x8hqtQu7AveN0eDmo8WpSjsUFAp6hRcGfIBzeNBmiugPg1a7xmC
+sRaofwxgqCoGopTHrGzefeLqS3I0b2fTBLXPMpzg99WPgkzQ05tEg0cG3a8s29r
bVfBuNLDaiPstGBz5SPh8F5KskLp1lOTrQqyJzW2af9o9pQFOdmquf5wWeBJPKWz
bq4Z6I69h5pldXb7H61yZ2ks1ShIUF3MEnr+O7ZxEie4m8qzMxISe6/B9taCGtXk
MzDDvYlk3sqiHcMSeJ0Ebl0qoGdevoDMRC8hEtzjyRie4+cdOE0flD5I4bmtr1iz
WPyC/YBRhWnKEGQX0LlhtBwJ00iAasH190eckTLQoYJhOGkgZjS12EynGcz6MGWy
Sh8PCgqiAccNtE17aKmOYMt/gZ1wRk/3A1GfPh25n5eIn8q9A//kfRHP7pj1nb8p
soNswa89jTsc3C5rOWrx5rBPso4GBCrJPsSAwO2peYMQ2+abcZ9eqsY3W382aq36
P7bMG7fuRIAPEa06h3VtHHzXCMjivRPHBsRJMCg1iyMskLL2sl/oVm23QkV0JkmT
ThLMSx9ysa30XgXYbntbniCHsJBjUx2Ei50KJf6EfltGVHmYDvQEdf50n0rIplTp
GCLXIh0/E4o96VFB9W4Ztf4k69yEaQeroree0pn40kvrRdIoQ8om8pubN/mNEUKA
SgxPEyoD1yhH3zB7FhVJQJdLplCHaYK4E9S+WyVFzjaMPZWB819WB9hMIFgmlL8g
Vo83Yf3i6crzuRXku3ODxBerCSKwotC6a+0jOXZHzht3RCYrVcD3XeLt8eiuqyUu
k3U40raiG9hl2uD5ofRpRYBSKKTeQoBhEx2QsQzvJwq09WsJVADTbOd3xsYLSyLc
5VOxzlgbQDLjwYSGsuORGpgk2OBMcLeeMYX0a1A8FsX8hJyMGQiFQfQKiMeJjr2D
nypdO5UlCO2gct9Wv4mfmA40ND0/ZP8didc7wrht/LxjK8CJvntH6HJ/gRCPPuOK
qGpCWUQLioXva3Vl238j940un0eZQE3FqTs5R0+lR3VdASK5iszlRnQd8GxJN5CN
h2qN994TPH8HxWsDcJivegwCFIsitTR9oIHE36llPKqqLaXprpZIpU//GvDMNWkh
paxcX47AMjkxUQng6/3EpGSwT0H9EagW+WRCv6aVw8L1v+NodSYCK26j4W2FmFMG
Eeezdv3L5Mna4PtYAd+3XlK6CR7yq1PSnP1gx7eDHdwVvnHko65hRuDyenQaxlRK
UL9OYRIGgpfRPGqAmwEilgFNQYkWZd541zlHmAWbAdd5L/aLI/ybENqeb3/A0waD
h+wsYLFHJdyyeQ4V4pgGitJp8Amb1tmWVkkLjq72PvzG7fr4TW3Gl6j1r4aBxXOD
rXpAhfKUSMoOfLlmzxFN6fR14L7hlH4dbjDHkn+XNvh8see+XsW4ofwsdwuN9Yn1
9ucSLGTBwFFmpH2B9Jjr49HSrE3VGd8Gd/6FOt7asIPFxMdjHNH6A+OcV0836Ka8
Pc7pRcYT8zMusQRIlv3Qxu5HzmB8AghBS1GtXGXdT4k2KO05NcSxzbhFj8S3GUIL
0vuehpwFXpeftFyWqWbrVfvRXQet6nwD8TNtcPI3mqFM/3m3R2No7wsmmWU5b3K3
dvFdH7DRSg+tSFkkz1llFOM0EkMcB1v2qEPB4Dx41W1UZ7HiDaIzgljbF2rO7r/A
EDIvVOrmNjffr03tYNAbPUEmCGSWgdv0U8OWjnW1sTSsHhfisf/3+mlxXABdgprQ
oVcts6z4BDu8NC1ijpq0KZwQ0AUgoMjhU7RH8f2OmfBR9XnwWDn85EvSDGtoe+xh
byHorYhgjXsmg0nIeuDgJ6oBZO2v46E4rJpsNQVcrqioPtto/E8vYQvzt9Kpc6zb
ImNst4CHfPYkqUb7iI9+N01afW4ESMllCHSEVPI6AdOgwDWGVj7EaPiJBYKegGG8
DiJq+GVd26YWQbOx0zNBBJI0U2VnH8iCjaLg0Izd169E7WOsrikZgxc7PDV7bEG2
Xl+M9vtb+d/fiPor1IP84vfwOMAGuDqrJYoIJzjcUuQ6OvSuN4OBsiNxOtY0lmcY
Jkf8qzrKNHw9GcTzUbEFDRieUWu4UePfMojxmWYa5hoP+b/8IGim7cMDgOYCNeax
0BLKuDhvbkNkE1kADFbbRTBCejHMpnjesfgGytz7SXsSGMgpRZmd6xhmFsBgWQcs
0Qgod17qvd4dhOkk+j1GBd33U69Oa40yTngogu/pBi2k22dxv9J5RJ16xoHCwJUn
+du2FyPHztMmMYgmEqDaN8EWbvw2Xj3rdh9ZdXRrJvO6w1OPhvXW24XPlT9tEZyh
puJsYeVa6lNXW8DYYBylUUWEEjPsbpJsxGJcfYDBWjnsxWdVJMQBsUy5Vl3czEWs
AZ8KXIx5Dz3KBKrca/cqcRKjP8efmDSmjltwGH495tOLddvsBZ2jG52ZKN0Ydoei
iEKQ3xVHtvDhW/Pz57lgyhhPPvoe7mg6d0wkpNJVfn/gHHWaOhqJZROs8dbEMYok
Cw66ACqyQ0KUrb4gKodK7gsHHD30bQnnePyYDAw016U1ZzsAtQI8EKiqCBL3reyA
k727/aZ6fIL1Cy1sSzc34vJ3Qe9NVUOHqBDur3+5GenMGcd7Q1ziXxLKcwzXZ5Db
YdpgaHnKUpxBMSFPycU8AIoG1RdxZyVVuAjJAHltiqfl9F0c8QtWQqS2y7vM27nd
sjmA4+vUz3VFFc8Bqdpvr2d5fGy2Kdsm60/U0zAyjra7aya2Rl1HcV9laXqOE66w
kt4OPkw67CAauK7LSQB1NFfNN5rpC1SoeFaWzsfkDZFDRB2Wpnwxq6dkE/j1u4i9
p9CL81guYmEQSpqIWlXRmPK71bdaYvLy96xVyWVpyy8GAG0yjnRmqfDvFoyxKE03
Rn+NeINLynJPPSxKND9iMGMNsc/1bctEJ3ik0NGiC/Mx4CYHve9PAyn/VR0EaiW5
GYP+XzUitt502Bx1BLSTO+mfXXJck1QOEWXlsYpDpcr7p8ahelVBI+SqJFU7KdhA
GrRIERX7G8iyn+7JqEeut0CBOqus50eP5+CE7WUR1X0AZfiSRMOeaSPyP30BY/pv
HvOvGiLkyNMt9rmz/plRY5rsz3nIQ6U2Pj8YnYIlXIposN8jTe60jGHhVgAzVc5T
SpHqMDpzIP2YRUpkc4vaqZ2gat51Ts+EkWIfH9ElxTtSGwhflGLnxk1ORj7vYSPx
0nmWuRK9qAtmqJ+FoObNvsglbkXdubPduKrVoFhtgxw4uDY5wBceOcmA/4nyy9wf
Lh1Gz7DDhLq1AEm+iCqL+yCpZ2vNv2sxsQHWN+Q8wCGXhsy9Fb/r22y1UYXw6i58
n8Qq6sBzsT4MhI7BH3gj5Z2qoGkTtqNca/fgx3CygF2GlDbwgj9XvLM6RHaIsRS3
D2+pBytCTIQJI+Rbm/f2PNFAafmWfFrRAPbHY3HkxZ9tRIPQ864AyjcVG8XmiAn1
75fu92XTQ/Z7d1YGljBv0cERt9iE2cziL9h8KWNW/L1Q8cMcYgZ28KB0GwZRIpDl
pziCL+AzXU3yhe4d1DW4oQfYYeM+PgaM3PKdS6elPK3aSztyXOMedx52QQTYmmGG
GEMXXVDS68FLOjlYt8oTawC2gJQA2FLtrs0Bfaa2QZJkCyYFiHTPpYW5u9OfEoyW
OKt3i4cKXu6HfEoJsc6BvTqfWDwBDE9Ey6cygbbaDi1978r9qvmuyiOWK0mvhCXt
yXt5k44KBuol8TBrEqstjnVhhNxbYjKAaGlaaSOsl/aY2LL65A4FNIrsqockGGpk
qpdVE6W1Qh2bKSw4wtv+15pE4iVaekLJ3B7ZYs4Mj0a8THl+Bh4mlEEvSxX0d/d/
U9TZKI/QXM8s10GYKejHHphcC9FdlSVBwhfvrXaTADFeajrqIKVXiYsttAIQCKGp
5MtLJaXCezI7dzpdIMtmqz3NomH9N59PibSGr4raiqsCSuGZB9FTH4Eh7LHHlbMQ
FiYULzpn9YxZ7/ZFsrN0f8S3vFS9uynBhlvSfN926aCBBQYWFM1E6rXgxmugT2gk
1sZF2MrK/oBNFNiPbGcoblC1XCfJz9QJEkGm+ou3BM73a6f/YwA8sok+3fnu0RDu
K8sPjrKOL4fQOYpXrme9SCMnDdYQdIbNhYkETKkDFFJmBtcCR2R4Q/vacoPI8lD7
YOonvpDqzZ5eA1u8quv0EF6v8XICgNiJ4zIcbjDfUtbbXKAHWB8/iJRcXUP3rNEY
k1wskByJRortj2T503jg/xKAdKNemS17jIzO4fgvJw0Q2VNnOfOQnO1nG3VZiGfJ
jjsvs024mk1sNgyxpbCjGUxKk8Zftn7VdUoTL6hgWUwyyqnN9czGOr0NeDsR/IO7
SylXbSlHQz1jd2Rxp62XemBRJ/NdkhfEZuZbaYNJQ7nzj+NiK+tBP1Ti13K78ICi
t4Fixk+lbIMqysSDjOoXhC/IPBgOP+/5NigUwcYaZhiHpnxeVoSqbBIYgNMUPrII
syDsnE1iSWDYjAX62072jdml0vL2uO5FlfkjDszGI3MHRR8lMe8Eswhj/GYoDGt9
sEUdh2kpNXFcq5m5gxbNH9nAfUXqV/iiKJgc0YxvkS4e3JAD3MRUDqLx0hQD5w7z
ripiTYV0Qq5fAhV/TIvU5sDl2qxAS1L7mQ8D2KMkZXXisJnJ5ZiSGtV4OnsVY99S
okoIoefstiBQgmlaCa67CnEPuOhxUkBfaSogx5JDKLIBKWNdNjVowJhZKpMTrenx
g5S6Z4wNW/IEiYf+4yMGcffFF7p4wermBK6ISPEu+9rGgpEpdVpjiLByGivaFrZZ
UIT3H8MhtHM5y+POj+O98FRLq8GaoFZJ6MR2Bx7smwjVPot1FQafS0xdhW9GRcZ5
RdErkJC+ZH2emhTrtjf1vvN9x9swkq3iS6GQg7mag3HXwtpRghTZoc3CBoNgHFZ3
uD4TfoMt0usNk02jbbHYY/ZoU4tnl+6v8xgtA6P1PrqKMqJYNKt7aBLTKPKNv+0I
1apILdtXNLCDMwPoWh08iLRITJpg+XNY4bVk1baOU2MPM/Z6aAjUoL47EyGCJ7BU
vmY1m+A5cRvsH4MUHtgZCSBynRHw7LHRCiWCiCwTzaZlLiqgPKhGCyig9UrI15wN
xE1GzX3lMsUGDuriKhUisyo+maCIz1tAm7pH8uw+66bTR1thyJoMTgGvNbUvF4QP
If+yHHF8OLCGlUQvSColl8x9RyRmFYZYbpKArYhWO27+C8QwAwEBh1r4qZnkdmft
QcHcKinm7iXfv32iMXYSqUplFuPy3DrtgTCmZAEKqeVFRerCRXlZh2v+zbFIugRD
edtLTyj+vlgtcmbhbURofw/gPKzgZ944U5XA1pn2/CyEzAAPzAum8SnxeP6yZtB9
eqO1nULmklnrPG+CM2O0qwtaXSGG1JLgOhIbuu75C3CQpjHZoehmauUecK0cdi14
tlsPPCabgeMz4eCpCJJGxKBaUfpIaxBCPshbysgfFxFieCXS8Ew0Ll/0xVQzRS/C
zLTrU/4msi3v4trnkM8zqs37kkm5ec19E/Y6WvI+JIYRfyKGz2u1m0INJor616R1
lXIEZlDrgSN9Mts6OKLPSSTSYTWq3CR78lwI85+yDCqBguEfGJAAPd++9RsX9AV4
SWF6fEcxgKvncq3jzkTJEU0cY7mfS7uLNdx+YF68M8qpZLKZcq57+IbwyzGyjlEm
HkzFKI44DT8IowN2IQBwOJ/ZjhLLImE9R5fdDtGlCdx8yOdzfIryeaVwQk1M9vqc
x5sdPbT+m6/Z/YPreVqGvBchzOym4jkl2FRp/5vlv+DKGgcOFPMVB7PjKTbxC6B0
V7fHaxOdI7V5oy8QHVXfY9nhpn6RgDsTRYqTkB60IIjvVjL15aBZDJCqRMOupGui
C+dbIFiQr3kR//tZlxgmnUijgG1c5xa8ViwI6+mBMA+NggZbAUb5o1Ns+fnh4vHm
QRaXPm2dS23s3F6/2t7T4LV/PHub38enSpWN6VrlxYEporjTZQvhPqd/YfFNHxQ4
6/LzZ3iARrcA2BO1GUpcMESNx+888JG4miw2CzyNSLXiFm8D7ElCEpyigCCjRbIw
KNFKj/R/jbo/XIUCk5CjNYnbRJx7RoCQ+eaWQ+Di6wt1zZjlyZjGOj0inIQ/rJZS
lqgnKIQTTYNMdNvcP7+ctf6S5TnopBzS+2pPU8bgbQ5//wBP7GPrNV0SA0V4AzvY
waOHMfai3yds8hvo/qadTSnSL86M3j+HR/TXD1XhhG6C8jU7aTpfJKd4jeY53+vS
nwXlEgnftKd4HLWMdFpmoiCCIEWoXghmuNEVwG2Y564fXwVnwe4kJveBCz4C5xuO
1DYjMyDbdtAial/Fq+LgHdSJlP6T/kMKe67gzDU+7nMFcOFRqkMg8QIFQZOCpECa
Evwr9ti4oQWfYQt29cvQzzXXCt0hVt3NO4GrqI+GgKVNv6ImzoSpiI/ihc8BYOAU
yI0DW3TOHWG0oeZZUZwGBtKWrbY9gMukfS1PYV9igmqxf6Qn5BGTFtCu+hq5iKR1
9f2bVuNPKyWSfMaJ+LNlls5S+X6J9FmHfRKZ5W8BxSb+3TpXQ81kbY8qAt6GQmab
treI+/cb6koyRkCpkL3yOQ4Cw4kGQ7S8MEI+CcZEOoSgZDuXU90PZtLgg6n7nU+y
f4vvDfKIpuSatQIgkSdUMu+SaRDD8snW+jqo/vTWIqZUwq9HFvtG84zoPOQ7r4Zz
C6PRVZr+ZR7Cc/xhl8t1oPjwUkrnQmNBouAXe1CGwKRfHhn297X7goytUwmLE40W
GNFsWH+i0K3I0w5iJNe20gsGE7rJvqqtFQlU3LoqUzKK6RXJhXiPxnGEWVWr9e3q
tw4112f3ux6H4CvP6UnM4Fl5eAWD1OyslwazBFEjBTXfiiiveA+lt9UqN8wt8jj/
aFSF7/fnMe5dbHvEAQwClnO6Rfbbup+cD1NchK9bLgBgG5FvGVxJS9/4ohexakJm
8qCfic7WD2WRsF69YVnB7ZEYQyx2TY90C//AEJadDmEBZFah/lZus09Um7O9Bstp
56kQ5oV7TAbzVNjlbTLwEHl8LgCXZmStQgiJmDzNWvQKNt4ZBooQpEHHNYgCrK/O
PBI91D92k/CHZYZ3TQeMWziFkPWzFqTiEiRkz+THzFufjyb6GtItIkjEMosbShuE
ISxBQoEmHjcDegiTvoX6GqH8eZU18qDJmDelq+Qv9Vi9NLTCjwG5Z7YCZsDLY+pV
vhdyI/wb+LEQW2dzjzaQjGR+FeEpkMYwgJRUiwL1KSqX7Vm6rM+c0K17kDlTawwF
c2kg3UUTm+BZ3z5mNEKo7fVSgQ/mbl09oT+dyYIpbEwVmK3hwq7QG4yznfNsrw2M
3kRQNb7GDEqjPAwm2Oo2aYyjtf8Sh1MmPTgfI1JKVgsXhW3D4D/W5d0xLXde9O+U
f3mpGdJM5A/GzQWyegZehKcj4pln4ujXXeU5utrc1ygBbJXpRQAHnw1y82c1cZB9
GM1Y5p1wXIPEAc1vUzRBsBYaJpcEItLymYopn4gfTfmXbOKtdGgzwNh0XgDPUtEr
brL5SgTi3EodzwmrYsKzVFnmYMEmjK9BT/VitZw7tutc1JIheSXCDwV0yKBQsqfQ
EUX3sqminYJKZGKqGjYkyhyq7wqnCLfd7/wT+7f68sHoHFk0ntEB6xNNrh7ZzH1d
H/8/zoHo3QQQ2HR12GlT2lXNXlNdh9r+4SZDAWScon8kbfgUwUUigxm3uY9Uc0a5
nBHzsc5zewxJFIgJ4GqpCWG4cPkYtsDVvVVIrziEV+aIAprl6Cg0sSLy4q7kMebr
LFws2xIqc4jjpLJ4CtjhN0rG5bMF5xAesohjsqW/T+ofgwtr9OLl6DHNCe3Fz3Mz
nmZyoF6IBuQaWbnVGmf8QLfeEi07mLsMOoMDPpBboMW6MtKTOBzQqgJkbO2tK6M2
LnQka5js+nXDxj5vV3YfffXGsqiveSoONyokflm5EgTZSErZ4UPOGIRUJJk7TUYt
gaJWr28+ZwwdSlakI84FTP4QUO06qJM4c68p2jd9xNDscCrHGxJWeOdRgZhN4wKN
2eZDV/pZYRiUN662lmDxN5H9W1cHm0PuVLZhkZPYnQ4drFnNn9ontOcIbD6GtdIt
7OP0s4qwuC6vo//g+KY074613ctW40AClImA6+DZCVfAdeTb+iy4zsDvwH4pxGU4
j9qC6Nmj3NaEUM4/shHeQwIxhvuBFwj1fjhsQa/+/exN4Omway68hoZ6qMtEXzQa
scvxqUv1jkk9gUocUR/PbFmO/BlmW9FSEpmwnVjZoNycZDuVOBKdP9TzLjLcE5ij
mgrBkZ9lIFZtgeOLckqhWKXUpKxJWcwh7ppSsJZ0q7ta54D1R5f9QXQyCqmtRPi2
ho3ntptim2/DF9CkV1eMpZuVc2KGw+22c5pLJ4jBzgcsjWX/34xZI9nwn6/mQ9Bx
+01WNUG+29OMpbMpfcw1Ee3unryY69dqKqaROgfk8TlpKPEvzZ2U+0LzY3h7+AMy
G5FF2JBMLyr2gJccrVX95fnvFOG81MNcIsOG033vyBrbxGIghDdteoIIrIrE4anP
DCTs3Cn964YQslAyYZGOuA2ENHCXycXX1jeIPRxrxZfi+m2CbLEzElA0r0i2P0ik
SLhbrKWfnsJWWzrBzxL2A0P/cL9/1M0Mv8ncmt4+3CfLxXpMRh+FXJ/z/VJ1MUte
uMwnfXNHeA0kzUxsobVDGkPKPNjI3DG2Q2zFK0qPZjIB2NsBwWjjVTLDwtcCBtTB
SwaefZpBx30yf3EBCwywl2/gDgHBz7KmkG+d4c2SqxEv+xGVRdzie1eM5CNPIp1F
QOChwMV4WeRzU97xFsPkHgpY6QvYlOjgPhUftBa3eYgfUqIEj/gUqb+UY00+1X43
oK2gUWXnTNe89EeQbmD85HiEcpmGClR0jKj/B8wy/IHu3hh41XRuTBNgBTlbGvhh
HTuq6cM3MYbqegKe6BFcfiKRFEWLVPSFh+tlDHl6E1CVuVCkarY3H2jduvFrvqCN
aV6R37zPSjolLYI4trElFmX0qL6uZDUvae6+f7njQZlCWdKd2ogVxZc/OrEcmZ1B
dDtcqPtvXzNL/feBQ6j85DGB0+6nD7/N2LTKxh75MhWv8osq/dQYHBickEQU8X1u
KxUYPvyorO7GZULLyj+MgcyX3oE05gOaY14H0LaCb7lgRo19aHD5+WryoYlqXVcO
ZEKeOBxhPwbA/gYKQQ6D/YAO4bWEnO05DDrIEfqyyTQa9DMXv0HZ46tVtny8Q8ee
BZ9UfgAV6bAZWoN1RvyWd0Jgtbfp1zpf/heUlz8o8FLzgkTxpEtTmhwRjWBLKfLS
ZKaele4+SbkwjcfDqP/RpzujlDEogA8/TzF/NXhPfiUx8DS0U5re6hI4GuNZUzRt
nib+LTAYcRrHeE7IVSUmMBNmEkHeW8PxshtqnNQsS5eDO+trahdV+Y0qBUjqZC8B
aFJqVr7tTHrMO1cVABkJz8JGzX13SKYPJGFJVO8IeMK5RelzlXs+fCZyC4u95QAz
q5Ft91YiH5JK7I6M4ZnhUAMyGPjVkNV74VAUZJSnvnlB4rKGMS0qNBFY68lh5/Xc
EcIhDW6cfMB0Vw6nwMh2sjmpVpRLjJld7DluXyV74imb1+ZNfU7k1tCBeuUBdZiJ
t2afolihB0zByWk/ZtWWsd8HTEONIY8SrhZW4RvK1K2udlWbf1CxcYFK5r/hgkji
jB7LLhInZ5rtuFYCZtJrDnN6G8DBCEVS4njXuhkaZUBtu+olrD73DeVt3CfTsPlV
RkH4w3E31i49kxwWfoUTcDM3404x/neVk66YXmzcL7z7GS1bD8SfTcorn2uNvSIM
X+Sao6W4EoUYWuH+Mx9zbcmATUq+RG/HSvTK6Ei53NS2hU2IXkBf/ShoNJIwQ2E0
mZmSx+q0/h6w/hz0drAkFxmPkMUsQfu3rNddM3a+kCZ/5LhWMAFEnSDSAF1Tr1wi
9xkgGfjp12qieM/KuuU/PQ==
`protect END_PROTECTED
