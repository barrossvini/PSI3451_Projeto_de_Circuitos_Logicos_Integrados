`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aPWBRPUFb8h4T5beiGnhcediF7Rv1aYXbxIA8Xd0CqIxWIvlHZdSKHLzDLSiNUdG
tF2kUihErhfAwGLNe6aKznVIYH9SNYGChnrLEKp2fu6HrGQUtEvQviEza8Jw4mfV
aEh/M6eSe4T9B9aHp6vGBE+zp1/nRUOHZvRlLpXyQjpwL+cbjVp42UYfuBjkq3TL
NKbRKTWstEQ9yWbIsrd99NLpvv8HdQSRJQKex+pYz3MK44lXde3vFhWLxBXV0P7w
fwARG1QonI3+v2J7cHFiITJcVu1DXRP3N04d7PyBKSB8cXXWfhF9tQivmfJtY5/5
4+3WcB+8ZvYDnmflkZrEWFoG/JMg5/7GeUkEWu3vP6L3vnlC+ar4ZvNJa72REYlj
tCglRmuAhoA/KasdoZONwMStvNFAgp/2IiTvdXrmHAY9ojxq5xOuWjg1IqURduac
rRlSBfojKHb/u0B/0FaQmnYLkitpCyEhbbMWycD4TQus0ZzZerpdUtkE0JXgFYX7
ya2P3vNn/aCA55I75qzZa+3OuwxskLOlgzGlNa4+0xoKYN+rpgZ/9Nq4MGlWLmTw
O88uwodzwkI6hNyYxkSPwrB6bUb1tvL7KSPJtufdODwyKuOBIwiNj9WB5VwfY8HU
PuNHrIAtpm3EbawHfq1+FwvuMggCTOug2mmatrnBRbAA8f3Df0WzC5+FfBW1TnZC
HltaKl5opo/pqXY6MnVYHevPMcIz0ebxkw12Jqzg5B4AQVfrEyayWXHs99Pxjxx5
GprgBfv/VM9Srs9r6c+3kl/gDhe1ZOQC5Ppk7sT56qjudUqV7sPt7Uy65YgRqNgG
`protect END_PROTECTED
