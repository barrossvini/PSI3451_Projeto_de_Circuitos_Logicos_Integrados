`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ZL3nz28Fc/LR2GdACD2bOBTJdVoFnIpVgfsK5MWFG5saTtfbyrlaEoSA+e+xnHw
XgddRiEwk2lVpTkJLrBEenXn+AziVwfoIK3qyPXhuNE8dvH5lbCQesQ22fwGqbyU
NC6/IF1Rfdz23kXNJgqlbBHHBxkpJmZ1SETjNapnrNG7nF51K5sGIh9iJ1FPqL8x
zgL15WPYwSGE/jZcNlN1A8LudPQQ18AlTuSaaHsOw0MX4uvRk1ovz4UQUoGm+HFd
NEZ/JgxviLPntvpcKFQdoOH0gnfPlQlNBbcx3da8wzhppsvQZHmwoaHMS4ha0VI6
RzJ782W5DmLqooJoxGVqix4IeC3APOKgEeVW6cTvj0KDgwUoZQmZxIWMHhOQUs37
F7wbi0/7rGaBcDgHXSzoia2LO73sawfTmV9V3as84Bt9nAQ0Pk7iNaf1uwlCK/gk
bLvq3qucZIVRlfIuXmAnJp1+ICj+Y5MQS0iR51rSe/N0/uSbXZtuIa4qr7cTtSR/
z9ukL1sOBVS/y/gYcGPXv2Nubk0S5yit8pzu1HP65HD3x0hxitJdzIU4FoasjVTr
6iKv5m49rZJGce3gNvwzn9kRMGcbc+cVQc6y70j7R35H1Tb5+Mk1hcGqPE5JIyrA
sjLhCNRrQmVHt64MatOfzuEBjipPmgkHlgGVUvqvvvrPEhpK/wTsr4tHbj6qb4y/
Ln4KRLgH4654PfArzcyfsMPvypqbq9nmOJMGhiqR4VEqUDSK8Y5r23m5vo/D8z8Y
XMbk5HAgWy8i1sQVkap4JlnuSmEh1Lgt4wE0KP++SmmGAx+RiQJgN+IJfXrADpDM
15wBV2lvXF9ivs+ERt0isU1H2IJsXyqlVt5kmd2kc8VwD2ES3dwQXHZ4sRYUMhMP
p+KtsP943WD7pzdTJ/FxECBHEnEeQwCsgpGDEQlvlTuDjUHqJdrUJGERO01W8bYA
Q5JB6Se4s1GN/zj1L79I88JAJotB2IUcbxBI/qjrr9GOY5uiXYl+d947aB7c9ipu
YjimoVlv/Lovl5im9vm9E+gpbMsBBmm30J3JiFMDcI53NcrvCWsfBcJ2XYtkFGLX
kwoD77LAUeOOR7Iai+2ugavz/kPz0WVVUnz1jFVEiWTHlikvmUPJATj6B2HfgEGK
hDsc9bRF41IaWJaNyDXhgZCHilZY2hJ49oJN8/Ti8SnJBB+Lv6QyzQYpyWBZRacS
jKHnwFuBzOEFNUMXgplrs5OlwmcCebiv5McouM/lX6/Ec7WVRovk3LSchLJ62o74
sGhyj6WwBORepaVzd92yUIevUwZm27HgJDVF1DAAWKX4n+kK0IKhyA/mhE7f/OZW
H7kIGyp/wXySe3f0vv8/mbjtMPRXn3Pu51jo7AzFMcKKUC55l586BAUNbFHfClqN
jJuCBX4ewhr6mBhEM/LOitAY2NDYu+GqlvjqFcBt4EoIrwT+te4ncrngNkXjThqw
e0sxnR0FY9Ib7A6Dx/J0iJp2LTAusluKDnBVRBR5DADpXBVW/Pte+4u35YMvAe4B
ckzYFayYl/UN1PFbdMW/crlUOi7ltO6BgF/DeW1vP9IWWTwCSgHDDxUAsAbJ8iow
D+j5TfbkOqxU8MdV5WPpsoAlXdwQubLH+rXw3TK6IPMRrXAfmcrrwLQZsK09yigA
Ocqkr/cPL39aZbotQlSrHUBXjqlkAA86k2Uzvk13vyVNPbPcJp8umF5npvfxPyHk
4Nk6wbwTlKIXdkm6asCwZ5i+55FwRzqHUAKRDz+4qc3ncdn0hCpu3EfxRSmBAXYv
JPsstlS3kmlctOtET/k3+Dg4f2OSmnpEk+pslSnQc+Gz7/am40Fg8c5tNS5J6juC
1X+uDikvKYnrQV3lNrI5YRsqT/yF3FdRx3WzhyJL3H3cPF7mIpbp7CUrVVkab0AU
wMskyfjYUWYqvDH/I0WtSWk0NpZHCgSKz5LRelb/aUstFLClAeiODAQ+qDxvERUB
ydX9maUoAj4D9udyI97grxV1n/jBZZPuH+IUPAXu3YYeQApEGJUnZfoUIRIEpAue
MuiE92hdgyqt6o5hJLmtZP++pdRZ16ZL8oW10ME7PHJdgxqnF9cW1u1O9h8Ghfio
HwiOWe1liF9kCBHFO0Xs3wbfajSz6JvCiS+/Ay2pwcwam2K50YcJnN8PCSM2SE55
Zeoqe+OkMhJkgwRJRL/7CIKTNpet5Vcu3NnStA00H6BWDYcsvFwYm28qqhp+m7Do
v+4UOeXwZQMac50LCmyFcNffV648LgiiMiuSlA+HpSADAznkq6cjEhm3+Ue90zIP
10nRFR28Yh0s5audfTP3Djw6jskS3OvENFXEvERxW8W9R3T5QzSfLbxJKLFuaSEs
764GMGb3t+yDkksAl6j89eVZ2Teik+lif101MbPzVdtsppP/M+Cdn6d1qdGHCx/o
PehALUNnsKKAoBWcpRR1BOPnapsYzNLCC51q3Dys3AhwlRJ6W24awZ+l9mmMR7as
IwwzLhYJkpuT6fOBIi5hg8YkgPQ1lHO6W1Gu5A3E3oLfPwvb/ElQo7MbjQmWH+ZQ
b7qHDDOXRHUFcCmlMTF1Hubvfhc7MONtROYi/ljnCtDgIEmLSp+FtSgjn/8ZYeMh
gcI/go2zf3EfsVdpjay263OhN27i+ooekQHgFKRpdpt+/XPnw3flCloYmw8VRv/E
L3wJPattcSqm1N+AQZhU7ZGDDBZvdNy10qEwSCClZq58u/oiujhUpB+C51v1X/16
9gZmtb6yKxoKl+84hsPNqPIaaiYL0D2hRGZEIExFyG7229cNXWUQsjwhL6TLUPBT
1Bu99R3PRLDTWQ0K/w8EwR8sfOf9Rz/iv9uK/XrySAGkuKmLwBKw7Y2mXN87cxl5
Mc9h2cBctNxQlwM0CyGLU4LlGnJdWH3S0WDWAlBhFKGeQ+sj0r3eZ+UrfMhhMZNC
DIeUqIA7PeikIqQYuykHBexiEgDGafvubY8p2POeVp3uQgQHJMWbtsvXitYlf9yq
Xxo0cXJIavk+8JREmJ9uFjuPEhCwmnWhHiZGqA5PmtpHuIvKxpzX9RKAPYkOOhnI
B9BPddYP+KHgTavEOZVUTtQwsfw6r/EdB6825V593K/F/llOnoAdaOsb7rQwcrY8
2t5RLI5UAJ4UuZ5RBbXQTlfh/CYr3pPPy0pxTBSeH+UKn13le4fznhRUI/m9napb
Cz0S0jXQCMyBUYyoHqwcFvOCK/HOvT90wgqBbrY1pwYQ9crqlQqsMlDZbJbbNGSx
WtjypmTALjti0ZgeONYwv2lLWaAcafoG43x4Nt9S6hIr567Cy1LW6j9AE4xWndF+
FASpxlLX/mZOPjegMPRQvxpnnP6anx4RRp5DgPe6dcDGrZ7YHlX0A+C7pJrEPn6w
x/+oUYhlgpNcUm/vLlhnwKQWtihXkQWOJ0rYHNzsJd6x03O0MgPYvdVO1WXOiMvQ
QrLThaXaPvd/2JkmVDcXPuqLCkSSUu7/1t+rqOBfTeEUnK/kcUG0jbQdLZVEN2sw
lwsSC1NjGyMa9rQNvy+AFeA0ycGD1V2zofHjXMJXdKH0qOIDlttAaTPTNokdREY1
k/uQtrgL0aHB3L5nIENq878nLQrHcvONzivMDkC7Xq6drIG2n4mmfvsmD0CbE4M9
tEGkyn+Tb8QJxZg5bK/THHEsPP7DtLtTXdnKrNKYLA+wE2DRNeQU2AihVE6G2NKu
bSsgobAh155MIJxUbVdlMrtPJCUlJeFGUIqFif/bQbT4/rRjbcO5I2gjeLC4VOHP
5gdGhYSTElBBa2Quf381oOjAMfuiwiqV7nIRzkIf5IOsmFKZ9sEvlW0fxJU6zGVt
/DQ+Ad6OhU5oJWSM25WbJ0IzDhQdsvKDCRjuNWZ6l9+g5fuyZeCOpXsSC+wIMyp1
bx9T42YvkjT7QadauTJKNS/nW8GxtoBilcCizjPXXDehCym4FrwQy942qyU+oo8v
OUerxAgykDahaxfWN9UI+hK7e/IgXTs3uuNJs4/g8O9AWeeaVA2IYX8hruyPzqU9
4gxCREetL3ktGuj+Tw45W3WlpnOo73koosOCW+qiVrcroSpheBKqODYMWhAbHEF0
J6YwfQXwzbEAtaqNaIoNWIq/D5x0WijVf9fnJys6cxqeVsJN9h3El6cFBLmbYovm
D9SmJrZaKTVI5Rwflzk74JONFcPH6UMQAIUS1L04eB1I6NI/7Q8XT0P5gNnNhspQ
fITiLJ+2jzO3dLHpMmglTtX2R75/7n33SeXObLz96YOx7xmA2vz1f2ya4CurrVXe
ARG/ewgggClK4wywaEfggLF6gWRAqyDhL3PSBO1dKmz8X9BE4PUvQ9bIUYnvXmuO
Mp9VCGtwzI/79lKgbNsYY77hb7thjwjUvfVjS4HvrXfriDnRnzxiQkawgQgdc9UJ
qoR+JyUTMxy+m0ZEYw/jVh7R0upoGWGAVOwkyx30Gk9R2Z02Ah1+PWyMqfY7Dn9Q
/OmlKsbQKjhJm5GhR3KtBfYv5VXkYjyLpKKwIIZs9zdV4pY4jyp2Lf3DDritr4YZ
BnEUtwQWPNeyhRgPmRGqv24n4s9m66m7IeCEY9wWX4NVikyDKbdYpbxgPxUSQi1N
yya97FDDAo/YzPNNB8tZ9tUoI17/PDTzESA9mQKAqz14hTFg2deFIxcRgAqZEwBM
ssIzR7Vooytk5j3zGH9ZieXH/Qukki/IFh1SiJhlT9ilXPCSDvGeg+sfV2pbmJJY
qwI6Bf/5XQFRRNBeoiqqfHi6g+hS8kWHQ8yfFCebLoulv5wfPdOqZcusUKtEhKQN
roffZMKUR0NrMR5IGxzPLamUFBkX+FRVgy6H40yiyG0owI3cgL+sg+LkXMX4Ys9C
ezA+CRtz5Z6kq1o6PA8iVuaVdV9R5tV7wThE4ezKUzhuHoERmycjdEcH4Em3UY6f
2C8t+fvShO16fERc4kOsSSuYE2E/iywm9H/TVcsab9BiQyiBaQoqQD5GC+0IWTXi
KrPpNWns+1cE1R8EEs3ajcD+A83oExk3rGnbF9NTPNwqFiH7X0XpqzNI+44QyY61
sEaFDTvq5H4vgxogXwfFAQXVwrHxB0Obl7Lp9Mbm6zONhIpCBIrrBcGGvKbv2sWc
CK97oLiT5Pe64vlhAW3CT/zumhRfZIQ1O2BGmRobvqiN+bNctZ844xAFpekjcWm7
31AezgQK+htUxRZ9UCFHy+9DmpmIucIBU8ik1GK/FiXsm+dpFD4ZPsgcik1sslZ2
EtH3DntO17oim8NXWTHXPzM01xHlQKL120Lk7785aW+FsowYTXMyUpuZ5Qe6WFWM
8dmZFOQEVdsVUkt4YEF4gTlOq8ibkjLTQB5WUbNk04B4XotTHR24edGwgoAIGnfQ
gmkSX+/WoBZB7Wu7bewNN5xr3hD4r/eRQkLQ+e/xRkzsAyHPj0PshkIRnoAw8suC
FOn/2idAj8Ap1GAFbeRoEfmjdmsrCTxhj0d3KmF/lL+zWKANukDTe4D7q9eSJPRo
VVGmvV5MOWuIPxgPdJ2lLqPc/fi0AprtJxvL84fkMdHK0FWHegShsAPGp9UoJibv
L9f2h+phBGGonh6K1AOFNmqCwGc8UIcIeJ6akJ1Kj7TzJobIngRY8beTriecAkVb
8/7kcnlARdO8Ez0mRAbajQ==
`protect END_PROTECTED
