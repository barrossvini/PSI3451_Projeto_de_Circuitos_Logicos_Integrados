`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Bd412bGHME4MrLwQ93pZac9wF1uhP8l6BG3OO1tcSVcJqs9v21wtnXXgUA4ak/m
FgMy5dRuakRPEUn2Hq9xxZeeP/eLY5UwSHmIbeSscN9I2VYnzlDxAYxJChtda1F1
AapVJZTYFnUqD8v5fwgpMjNloV6g7HXvCUUrVrULrwxv9gbgOZOeVsVtR34qfzBX
fI/xaR9HuvRlH9sRcxinH1TPGMawR51y/F5BNUbcaxkBUM+sZ8swPmV4ER6AWtju
CryifMgDFdBiE602JtP8H9kGIMpAyxHZ1Q1Du7rXareVVZUmmMkInERQXMaqpJ8W
zBKq7lmG2N8dAycx91fhlMRNmrEnEMiwptjRkuyI6fE0NOllleNavk457UbsqY38
etVOVCsEiRPn60XAMRs/3CUyoMAEaUX+z0/h0ylG/AnYdcL1t+MHweAi9vpj6ktn
lSqLF5Ukn4biIsKbgDJ6pZ/OuIp0zbff65CIm7YVXw5sH1taURKd0LNdus3JRc5B
zagPp1+igShtd9J7oXZwp9IQnDa6CTblehzjAJh6RXT6Fnt1/NxKVMMa8hO/5NW/
RJR/zVKcAkqyQFWbJL1s08NVkuTf0S6Fwd+2ou4aM0iaCZPswjVdrs6vOf2gP4fE
EB7HyCrgploxPsabTeOyI2n/T93+mLPCoF3ZIa4Tw1IermTXqES5zqctjuipPGmf
YtOIQ55FHtlsxu1y20cbRRFU4R3X95fwmnbeQVsLNojBgWJosXhwoaWO7kDJ7g91
tXinRtygL8Tl1TqtIZVnfhDv4HrNUQ0RbQ39dV63oe/GCOqFsSo9xtwZOlN3xycp
RhZ7kUjRy66zrhprT5Bcotg2nrrku/SREGvTPYIRXfxBTVwB5SEyx6bR7teX7uXs
y84simq4IITVtcX6p+ZWEQp0v44DKRgTf4hj9euzalMleWIHgS3lq9OKcsmyOBW/
375ZX3ChVkwi9Mmg2+7NGfJ10pC+uaaYsaypqQke8/ed9fmy2BP02tXk2mBlYAM/
2a46m6ox9u83ljelCcCcBdOkopWfTa88C2OVlF48aPYr65tRNq2sT7irLUXKscqk
VqnoSeQSfHoyrUG7eIp0MW3aZXcAqqWPZiVmEd2D096JpC2kLdf4XRWZEFgP6ztT
KCFnrKYZDNu3Zz9agFh/DkyIJ9OniIpNLrU51qeIMNNey9d3nCC5hJmdaFHgwflY
GbINJDds7fpzzH0txtNQKAe5Xp1bzgiO+OcZynltT5ngKbHakx4hNQh8ZVDkHKGi
aiT514WT+0cvpx8eXbw3k/isDTZyS8kL+OBoDM2Xbp/RUXteUNc7KWragfbvTWnP
BNp5Xwh3F2mp7uIV4c4Lqyn/dGJqUnavEtB9Dq4CEcKfcCPBoxLhnUoHrSB0dh5e
ikJx99Uj9cMEH4kDuiudPdsBRpUo1y+xP2QFEZYu3h5u4FW8jUMjccxrSbb2GX5P
ka1KLBpTpbcUOSKBgLh6pNA+adLIJKS2LyvsUao6ad4JTkqdOd7a21aYiN7pIA3Z
B7qbtAuRK/FMovAQbkfSD3Nk1fOIK5jdg51YeLLtRe8ESj06DTjhL4BYUsJp/2f4
PtAyTwNoWv3Km0UMsaQtP5aaSyTEAjIjQ4CqgOgNpKfJFpu69G1hIMMfDAn2kmAF
NdHd3u5/B9PlmFftJ0+QhaeF343lPkx7qEcqFvCtzQarlxYhQN3MLzT/b79NrOpI
JutOCZ81M/IwM8ENYxfymvuZ13tmchmrjLpDs2VkWiIAjO1RyrZ9RNZVQLUWySwk
`protect END_PROTECTED
