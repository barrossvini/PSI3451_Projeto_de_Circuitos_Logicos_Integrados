`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0gYkNsmUPs28Y+/vfP8/R6TcP/nKFTmsPYUQAbJXxwCud2oKCITWnxI6+wJxRM/g
pRg1VfeojN00NfkkW+Oghg9hfOKfPdx/euhvUzZxVWLCoVDcC99iO7DZlYhp6UMN
nPtS5Qb3RTw1DAmbw9Hh9FS2AQAQh280lw4VhGkB0LRvNuD3p7hlohT66zh3q1fW
Vvik9hKS2id+C4u1MqANbX5/Jl3kJPSPRXnOJ9zCgN/mL5im4wQ8noXweRqhUVRK
yLtERd73bXklqezacFALRx3xxfurmXpeo9gK7UQyAlzsEVnOeh6KfQvzPepMRMpU
EinNPc8sxqIP+/uAEu5e7BqOfHGTUzg5e6CrYanW1Qzre6y0x/P35TiHIh/JTfhZ
bU+AqVKmcjLb3Vel7/wkSc/agQa/XHnNEtPTiUd89BEmUb3b4ZClKyz0fVZ+3BN/
fqyX9yeRgKZmdKp+ZuBz4EV/+jVctgSs1M/dAZR7raIOjIqrSIy05d42adz1yDc0
vrEmiq2ByYnn2+IvKJZy0SjQ0PGoZkHL1miManlOceb01RT3WNjZjx56vdq48ZTU
3hL4V0rLtYMlyxr34eCOnAi525JU3RJkzz03fP629CntR1A68JMyxF2P4IyPjN2A
bhcYbFrfmuq1nb0aGhW8kjV64l8YyhHSC0eWPSLPa0npDKBfpzkEMZv9zFe8dvEN
hxaplmuJKMkU7ttr7keojbZPpEBHZcS5we7Dp2dAEVDl+rADN9kpCkJWDllqpTa0
/b3FiBD/MxJq002vNBd5y+BpIaPwrvB9G+BDC/xEQhwLt4jn3DpMCS6sCacRGtdx
eJLnq+1RrZrYy9MiHtuFL1zJsXc4UTl12oufKbZXLzkg8EpTh4E9ePqBQs/yX4Zd
dKbxwmprO3NHSQOMztWPYIlC97vgZ6oinnjjgD9FOUwKKRHZ22tf1EbOkQ3UZfGm
VCwfxR4BZqrUDVt1ndTDi2IAA0HaW0YjeiZ2lvccQV3E8E3a/pa1jbTGa+dHDMLE
w3QO1bpv7XLwQEutJI1Xht5fux4/IuAI/d9dsO+hp4lrxMybGqKxeMp44Qm4zCCV
0AFAI8iPkNwbGwz3ddwDERlMN0hUL5czhw+ViWRTAOrJl/WlCsw9AUgutYhCOUH2
ZLYmPJKFqOgQGQX4qfn8UpjIvrGLD2BBe5JFLcH1t2aWVHbvsWvhLM/ZC54tVJ26
N2lq3Zk9H5TIYYa7f7bj/nyavFsHcqLT9swIVpm7gRsbWpqIiJ1OhMqQGq5MPorF
KSAHqVVizGuwy88oN1ZaN/rXqP2pz7ta3fXX+nwhR2DvKr/AICfFQziJzi87Sl5q
gUevFeppW+OaKClIxLct7ixXHLA3Eic3oVV4EhfB8Gg32A8kuyudBOwMJ4BaFI+u
gASQPIE3soWoNEbwOwBJW5VHE5YgqXejNIz6Whyf+aU6LoYbPhXcRw5L1Jn+QT9U
YYa6w8Iuq3706O4l9mILoSGf7FFqvnZ3h2N3wwHdhZzngT2G/J+3SNofucEGfgTs
ZJDkMh5hwD3C/O4oUc5H8IVAbEawDjJuBnwmRj2eyZP9epyDoNzNruukBHB9QrMQ
ZNNjjWz46ykMDlWSN8PfpvFJu9XpYn4q0l3MfSjJNzVfzXSOm4MfU9RY3T+kM640
R9Y/LZBgldY11a0VWUGgbxy62cvTiLXS+hpP7IQedS2DDDohzBrcaOd1BA+EoOVN
vGuGws1NLxHN8oLfCIS2oVaS9ve3NS8+DUpeuoTo6TzrApGRlHyQviSwQi5e/8vi
OMmmj9oE+oFqr99tvG1rII0wCIMsmdQ0V7baDJWchXsPJ+p4ruJQ5JMKRLzeB45x
BsKN5PLWl6MiN5vqCFUnN7CmyNOb+xOhZKDeb60YxmOroDD/MdIhliEF4ebqJ+t8
KikooDwxhJ3RWXM+6K0SiaK3iBnIo29SBv7vcYOAD8mvLx04ngWk1VA3zNtqlZE1
HaOFC9fxsGmXli170npagDR9yh6bp/eo/Yu7pS0updHfewYRrvjP40+JPuCqAxqI
bCGu/jwijG/CvAQ/8rNfN60VCK0y9EDBqWVfXLfdHwi+F83CzYWZ43crZJ59gZP4
TJVeQwjQO+iXQeBNF0iKYm9VIcDB+R1OKy8iiKoyUhOiDGoLixbJlaQWUjQQkDjG
qv2J+zxCfhy2hY9zaF91cHeIprFa+v20/OuwbB3hp3l+1AYPGN5nGRUoMZ4Ye1fL
NYXyaeHjrcpEjKI+oTtW1Vkhhs0RRS2kLWcZALiSwcDKiIh16EQvLs0bxla8THBq
H4/FV+dUNXd200dVDCzGd3tz6tHnRA5y5lgzkbBGexLM+yQhBPi89YOoDq9dsqRf
UxbpgQ1ea+vh5/hIuGb1GqaTzQ0JDYyVhjSDFG/VsE6Prp+9brGF2lizNDR6iqeb
DGZRRhOYOqQjakO9x2Y2wzz0IXk3QUJWijAyk8bklXnglzyRg93uBPYleqFj3M7Y
p4VXbzHKTI+pfWAB//1tPF/0hTiSSVnkrsTMfphj859UK1e6bx6JAqgJHr2B5zUX
zsCmCyaqg3zuXtJ4Z0YvKSMfcgrIgc1BbqmyJsRlS/XHCE+Y+qMzvpbgLvLK5f9F
R8eGEccc5oYSdmyFyW44mBCElkBd50SRqPerhLqaY3m08DTO+JKRgYpj6PhTM5ER
FgLcy+yadqGJtOe8zo37mxLgjibCTdgFboO4+28pcFf+BEA840U03Sq1ZVe+n625
BNE68xnWvyupcaP0LEBPVcwO/IxPe56q+UYEwtt6X/ShOCKpeS4/cyLK5lWBPJW5
mkuovMF5W+EKGv71XljndHs6v3u2SPeX8UIbtT5mtVE60xMHDPBOZQiI+3wv6sbX
e+iB2lq0nJYwFeZP90b2ZuROsVbs24QnNP7+uyDHIjQRjW8g/2RptrBayBpyyns2
VxC6peHbWLNTGdmodTzyBpYzGww5IBRnkyFmGgqN3WUwQMTZdqgJEQJ+dSPjRC/2
wRNOqmnLSDHOse/xUOVXn0Oo9Px2s8keOAaDdk8Od0aHJEqHZgfLgRXPU/Ciklqj
qOoZufSEmwDl4fExaXvsK2PLlr25SSOLBME+CU14oH4fHw5W48yiaL/x5XobDPdw
OHt8+RmUA10RTnh1csTluaZnJbb4wvPGcxDiIt8G2AkrnVx0vihcI2H6VNQRIQ/p
7gCu03mcpht1DnpQW+km0YLpfdGlhiAImJUDeFo79kqNFfzZfv/DZ5u+Wfl2LNAS
wf52O1VboWPidpj6zaOM1e1OV8C55eoL1TGTK3BfO+LhBEhjjxhWVmEZKU7TEfYl
XiVsL4X2KixTGZhJJY8R0o8vasFQmvYbK3IMxsLr5rxD+SZ7WB6z2tRjXmTdINSN
+N3YAq4oiF3bUSIFgKz/odHLl3y3SGN2GoUnaGrQLEGISnZq0WNOYb08lw/+MLfj
pet6QGgDMXG5LDNB4DpUmedTM8x2UIvZlTJI0pNAr+VYX2ZwQNSvjckBwRcxi/jd
6cjz1YG/IlLGGvBj1CmLVmz8ryv7ZcF923JhLVUFBQD1NMcrcInT97qo4E6PHNds
bJ+UlU08wk8XA1070Zccn7vVkonxeyZxnXxKK60sU4KPUgmgHXeGCBb/j2wqJxFi
RGzE5G8lsFru6OXz+O6JyTVlKgx6DocfNe+wFILIN7wvpvWavWS12qA8zd+kzZd3
Fl0Mpl3K/lK/UzdkPEFrZdlafoBaKuZ4Y5Pkh38fQwbnDbOWotTvlYOQ9ohv05P4
uTa+DZJrSV035Vm/eFVBrojw840Xhlh828u4KvLzDi4mgatNDUWEchZ+ZtWUzP6R
jsKzsJ48UnYxexLD+xpRYv9hRyqtfZzq5F4GFUa/m8v6C0IWO3nxVxNddvTdPlGT
kuWbUY7MK6689S1AZenIfYjJxWdAwLA68uio5/YhA7emS+XnZsRHZ1OrI/PeXbAT
TnF1L4ZXvtXPjQiuzT17GphPEFjTMZeULKegDReYGM+iz3vR2qcXLkef/HsNUJrO
veZkKc+HrKmu4nnQ6bYkXbce9/cLDuK/aAx3w1xAhLl8KHxUyY/o449Hu6PDPdqN
J7IfqSfo/9CzAXAbxPJ9kGbgymCOgarwq6DlPkHALNJK47+7iU2vLWQzHzQSzau0
le+dtI+sc+iRu1r2S9ztuH/0hKdgnRcr6Eoh2dDqQzQHbM3F4/E72xfaJZteCRTj
StrWOQifvVnrrOTwTKzh7I92mz7nPbqQaiIyfwPaDE2ulNWaW7I9p43x+Dwnuf+w
yi4oFkPzOXiHNmBnVEWqHqieFOzW55jgHIp2iFWTZRTDHg+mYMYlvH6h0hYB8NO3
UJ0GR5ekji9ygWhJ/vOSnpqT7U3l77AdQ9jPVjF5iP7ZpUPwzR2DNxoQnWH4JoFo
2aFezJLaBjycK5i4HaZh3U6CcODPJJYlnb6Oul1qdgIVEvPJG//JHhq+pECbZ+xv
uXz3pVcI/A1FFnGsEfxkEUyPk1SB26n4RgDWJy9Z526ZwCnctz0RYZqsa4GBmxxY
r5mYCBk/AXEdKNEFOpZgYBoG+3nEI8Ds8SPQK1Eycyq1VVRImW+rjtJtnWWlnAjJ
mRfeYIZ8kqHHHl63TAbnhB/qhyoSnS3jU3r/hKWA0Yt61iKW18WVhxXWMplwt7bO
vDgX839YDeDZ1hb2eMqEcJho1QNMuXOEnSbO3v3+J5xshMyCRDgYV1sUSxxG4z2M
5zyd3xddFSwMB1ND/m4Np/QPDJtLa+7/QWQF3zxgBBH77kd+geWgcb3ecYL3aPJk
DAGKI1nBqi2l40mt7gaRZzwv8q0bBAy6y36MLie70GjlzLdq2/hmAUnuS1FIuL1a
lDeXEqRD0fMBoJx3mom3/qZNUA9ntm/RVpaIPVe9U390+Pr4aV3QJVczdDCiLsEE
RSrVYZxcBP5GmN45yhkQqKO8sMxbQyUb/ub2mKMPY98=
`protect END_PROTECTED
