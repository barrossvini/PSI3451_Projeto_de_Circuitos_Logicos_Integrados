`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RwVnkePDS2B4pm5RwA7rx8Gx6JfhIAuAzbqSkrGXBOXF6lj2h9gQlP+oK8o8/yUp
dl07IraMw7ShM/4hTEbhSInR6l61vO4za0geMk2QdMpF/2BN1c2/qhLDPOpMjuaw
k1Q14ek3yuRL/yvcMuMHfJe8ESz+Yc3Whfd2rLN1gENr4dpziMc6bEwtivV3Hvcl
d6PZeGaXUo+lhAO10lFVTz2HKERxPwXlmzgFvGSMK+6NuhXS5CBE4cKvo9uDoEz2
a3x+sSjr6e8eBc1bBLdEOpr4YA4b6ljuXJYTpnSxwez25dPLK/QhNkWjZl3dfFpK
3eZtsPnO0Ge+ZnN3qRXvr2EujlZ6pqpvb6B3KL+9KG2Bcm2p/GpxI0rHlJysqgv+
3nZyy8Zgd5tFpXjkBkmUDU3ccF6kgCFvsgLPY/m3cQavFEGC0oEXHetRV6nluILq
Ci2sv/t8CG0ADFaTC/W0Xnp6d5Q3iEgerF5JRyVfQwHRNhKt1g+okp4JS/uBxlHX
TUi0qWDdyQ/F3DjSrDLqyId3E5ZozoVLNTKBuKemw119EtKiBfnNOS9lhLR4lVcl
RgMZaOW0DMAdDJvo1Ccer4qXx2OpK0QwdtY+J9PCSMg9wMqk1GCRC+geuLpgs5i5
pYuSfFFGjKfCrU6fMhx5KMXgklSWM25nX56UYUe+xRRPgHCTB4pQiebFAt3w26p+
xmfExF7eRAWVhOxJKAiChPCM7IS9Ydn+gDIjzZQB1kk9yphX2W/JLUZoLgWyKxZ1
bzvPEVF/S3OMzLoasdFm+uppYnKB9O3cEeqQWVquiYr9tqgvIHTqX2+MixFShzj7
ZRiqM3BXI4GuETuEfrfF/oiCXNCVogad+Raejcq79KFHjk2g6LWYAex5fqxIZrI+
JBvPbUa7lRAgwJMCE3bPpTMz3CfNxL5JbYfwTivwfoaNhEuO+qKpXavHEaCZxrUd
VgewuVJtm1zUyrKzDBFKKGS7jTsTMAXhHv9WCWtFrI5yHF35wNZWftxlK4wPa6ud
wkC5TvdzZIAvw+culI6/J+e+p2I9A0OFFOKokNMxUXkIKh/yLjwDUet5XwBFgVoE
CGYnffrxC2MikOmHG9fHZ0Fj14atvoCyj2OFe0LWBfZ+oSecyUdAVk3wgaKSI64e
FKOVpAxpzih33Fccjd3Z/XyPBYmE+Sh/5RD2RiJtvyiq2vfpZe7RDXgH89kGiDYK
iJT/CgVZvrW7Adq/h7OWkVEG0LkDI9Gh8hmS3xdoQBvqMBZVpeqZIe4Ph7Gsp1sg
69Cqstx1BRHZ/eCZda2GXBRakyTDgS93A4o6F1Iy0LNOSyMotsgHsRwCLqRq/MyR
gQ+MEBtNGI6aYOdBBo622FSgKPj+sKrNud4k5QmdHTWUOlUXjvSYBdZExAd3NQdg
+5vqrEfxWdvRw4HVK76hfT8k4ZAzchYt5LLhWI4qecIsbDKYJeb1TAScP+5+kI0w
uVXwX17L31N+8ZJQ2b8QMg4fVGwtABFz6GSYwTC4KBwC4WaW1nmvxbx2Xxtcqdwe
iHdIOXg0O3o7w1U0+gjC+ohw6pnF6Dgo3sNlJnXdgkYsfJmZ4rdxO39FJSmWB4u7
4FTRasygG+d2FoxIw8D1QJ2/MPWcxWbMC/H8F6m24wGKCzI308Dffz9IjVGliBXC
ysjShTNl1GtEGrxis16nb/WHV2sXptpyddnqhok3gv3WEV0qudt1sxoBPjvReYx7
j7jyuRd5Q/h1wHWzI/bhprL/LBPOh6UoYR7dEZxWdrfLQN/alMOTDf1qWAWnix1A
Gwbza0mEaHNj0XbuXopBUH9BolS4uL3TIDe3+HkpITM+ADH+RDgyYUkt6Li3VBMc
BHn/OCvY8xJqH9FGdrQ1o1O8Ibxf7LfbD9hLKFLlgsBg0Fz1HSn+tJl7I2EImdFH
Fs5eGMxN4xoETph1p4KKdimoQcqgncptzuFZa94Je9G2HQ6rXbjh1odrFKqt/2Ma
L5HFPZyom9ldzewE6LugSWiflEes5bc20HQxag5cVfuu9x34FYhefD6I90KJzcqQ
JEhSw9l5aPuocL6p2xgFb9fRINUzi2JH86obTBOtdlu4213P5GRtBR9cN2vzec0v
UnFk3aLUtqzJA+i3M68WvsSL03oR+z2niGtUIGLPlgL+KOOYMcZrr98eHiYMTtmB
LUXhyyzFY1QG7vmILGB8cfaz0e7kokSucYnwihReuEDoM3NjufOiCW60Mu8lxP+/
ZxrS7P0uFEy80od9pVApRa+DwAuH77NreVzzlX01M6qlTSw+HohsfPD0jCJ/24sm
LwlVMzLLUNttVshmkvfplurCSKfQBUCdXZDZu/efFKiWn/gBdDYyijOT5wbpZ6+d
dXWPSuQ2MPXUDNGIuxBme43V9v0EH50tU0HYcm7yzpJ75THXTEF8EelGHDIB6Hv/
ZFSmOngM3JzQPP+ytENZOI4wGX5iEYW73kYl+ZmwSxM5fQenOCKcHXorD/aH9NkL
nTRw/HAXyGhRx4V3KTAfpemH2o/L+wdaRYKaV7E6vmL+37cDQGBnrYO+ucDzzPlq
NdT8yhJZ3FTHFEj6Gmd7zLW0NnMEvc07rn+4HNWFZj3s+Aq0/vZRBUokntveA8jZ
m1bMsuDV3v7Y4uWvgXYxK5uzif5iVn+uhVD/742+zlE0FvfpsecHsAXIemCMofHv
MTwAS53sj1iP/XzXgoxsrQ94/HJFeXsHSHHBOYbe4PRHWTMrXuFjpqj1ZmHZQ7WG
xiQKeagYphcdTFZWIcPW5iyP83k3SUf3JRYMuLw4cLvbNzf/5vNweojFQfnhNzlY
nlC9VNPLtDVMp6EI1LnO+K9W978YcAyx0M3Fec+u7jTmZW4k9d7+QD3wkAwVbdLJ
4eKGBfGtco0SD4iVjXntymUdLZHA0j/aLsSEHAngpLSC07XeSWACqu4m3aTRy2Ko
Zp6V4x6I6qesfj/uE5bi5xncezOtk5IyHMLqRf9d62Bk51FZfvzK2CdmcqMoYL9o
zPKI5pmWHXxo+0OP9fvXNkW+ScrG35CfuBVlutOnCY77GudrOP9R+HgDjTqSv1Kr
nBn015D8WtdxTwm5CpNBonaAfxYNTV+lSWdr5DBp6+xrxDWoHWHH+NAnhH3iJ54U
J2L03IY+tBrQmZY0BmHV7HzV+DO93ZtY07SxyagOpSyjnjzvVSZCCjWLl/Sm0vRA
l26QEFfkPifOGpQSJ7IbGXcy+d0I6n7DlY3IfX414T2bsPPhUX3qev/fvjE3vNhR
yCM+lFcqYZG9pJdPRjfmdg==
`protect END_PROTECTED
