`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i1dimol02dlY34Yt5fEiw3hKxWxT6HV8m8rop4NSYRH9OH/6P4R4UzmxW3HIM5Ds
6V35HSRdnM/JLeltNtMZjYYPM4d/uIOt/c4Z7oUjdm3eJIIeBsOwhAsYwPX2uyH/
lV3y+xTbmX0lkzxKB8zsoyhCl3QJQcOz5BAKYYqYRptjmcdIkElIgVGH1ENUCKrK
zSg8I7iKnSYM+uiX47SiAXm4LzZwdZn7tBVDvQtZ9CUtPujxKLnOZ7IZ/OhgQoFR
Q4PwcM9lYQOi1EvKLxGbABHN+4xFVDb4Z+SIlwgOc9N3WKDO52GDIW2I2wX66PZf
EJHocXvyzmvcQ4jpM4QpzRoTrjIcHYVVXvboyaRWAidJRufMAcM8Y+67rsSmxUBs
+0p0DRBK7PdNoBCyljiZ6HSv0ybW4KQM0okcvK9VOYbwJLXeZ0dmq+ARY9UPaayu
QqKxjcT0L8VoSihsznN04S4DC+XwKw8r+BAKTWYi0Hr1AMX//pIynmSC5eEKaPHb
b/vQ2qVUqoAgnARv4y8T2AmIPMvZuZbGafyZcOUj99sZoBSkZeboptsV7xV5HpbT
nxkxIOrhN64BGDmfUOA5HPXpq/TmPtlNG76LJr+0BVBgKB3HiOFp7MKoHrYn3oP/
/C+7xsBA16oXi8udRIWdNWoUDepK4Yve6r82QRMs0vItcMyfh9S2z9bnPbid9U+e
C6fUsH5b8cAoNOJnl28/01NaWuWaGQAPO4nyMCPck6q7tQpe/Hvu6+WJMq2aotMe
bqZgvIi3cNbO8QFlHo5G0oFZ2kcA0wwe85jJiCYVW8ImQADL8hNOpdY/3IJBdDyN
OqNrGvrw5MHa68pU2abinAcA8EX0UP8b01juT3ARi+oeGvga/Uc3NjehDBSTCD8L
MeqCrdBkz3+c6wOsBfaadg2CgcFRygp68CD21DPiC56Ml/3865gZc1luQ4xVjmqF
JMFk/pMF0OboGcn9u77DLi5KYXrCbdgl8q6oRjmSNcjjTuNVAb2l9hQbN5Rfoobk
qIC8zFc+40QR/LqInQEoMkViWMdMYBOZ6Xnpuy/o34A8uukzFxJkkf4IwTerNxKX
4qlvXYQnTuP44dSb2RlLga+MADmrsElhQtkNwECIvdXh/e517csHlFbW8AwaWRp/
E3T4qTvvNhDEk1eJpZGZSfQRkR7hoDnV4XAwHXoPFXgYLrk4GLqs7eOTu2tby1Dt
4vJZ/+J1bS2PoHP8N8OJmDM3A4/ZkcqhIi+BUrUJ4roJCS3ipaSQFHAekFrfIoYx
pxa8Cm/0aO4JqpbULBlJJatEfOsq1m0nxwAWZJUOtlq1Iky6wI2apcSOyLyLVBQf
M2knMnBWVhFOf1QdzUYwvk7+HxecAFrL3HaA3r59ApfGcMYI3lEiB2shVArs7ViT
0E3+NY3OD33WYhZw+az+EMjPbWktLiRoT+wfDcHGm/StW3e5bWV9DF+6sOLG3FT9
bB7Z+Zgp7uUonv6lOpIEPZ+IeK97zGPDkP9VE+vsaIpcHyepUY+Rq9v/kZXSn47y
HXcQQbntcbKQcj7t2w97PKZSxJcu+D+Dio1Ue36G8ei32iE4L4DuCTh+vhHT59Is
WOZoupmaLYrMpzcMr54mgmZM2KAKqe6wELwbmlrrAFxWVZeqMNy+gqh9MgIkXfUZ
Lm9wwd0ldTWUYc3zOUhn3gp33xV0xZaSBCBSN5RSnSlLuOLjf1c6NkYv24OrA7A4
aVxDehw53j4eQ9VgjLlSSRmwGWTkaUYLuzsyeg9bKDcit4yjlTd4PFLhp2RGks4E
mjEzzXUB0Wu8SvH3ThjkH0V0QsBM+DpUKfds5mUv7tZCWKWQsT4s/9n6uFq4eovw
G/F0uYg13PLfAMKW3ZNNPR11VPyqZkD31ELfkgDTwR2acSJP0yqb6E8869AxtDlw
4zXO1htVHwurOQqt82+efvM7esBuyH2RS/5lVRQXMMYwHBQMdQPKJEuBetvJ18r3
5ZpxGKniuFhlgehhGoX49apKzczTRcb87qV72eTd1Geh9qzz9ZBloSt4S5GHwVVU
fdoE36mD4Pz2pQXMbyYD2Xs+EAi8VUTFp9EVIYAC+rfCz88L0pIWT08mCUzscaC7
z/d0YqkSy1bD/ppHW2UZn9uNyBayMBRi91xAQ3s8UR0F8XxovI4eJLeBpt3FsLuY
nbOuc+qSnix876tlxhyv85zjXxnPaA2s79roZHfBh4FSNJD+MuO/WIyRGbRDhvwm
PrFcWobcSinpg9L1XxAxzGxjCTDkekIkSu4TBaiuRGXOKhfGgnYJK7/aKLq6ys5b
NttDIZkUGlKxB27ATBSotf2hu9o8bUZDhewovR5eGfT6IGNGKMZ02UWeOQuUgR+e
zRI8cRngCpdXyBuW4gAyYqw6L3uF4MMymZahHMufG8RENqQ/z6VerBTiuRCOD2bs
kUySERFcZqB7B+tNBq1kw5CvBU2+TBibXjBhRwxbIE24CEz83WNxKaN7rNA0S1uk
ANtLBYrUhil7ArR5GKWEfRqkKfq0clxF6bnrfhToup2rljNrz5dFuLOLH2Qjujla
KmxBRYl0dh9jCH9vi9KadR7cDYzppoqbBtEmuyBn0XMKRQqoMrRj0R0bFLOt41n7
4nplz6eQopS60CUjxOpxjKAADKBA1qHZ6Z59/mQiOCbIpsuOk8ZTXFHU24WEoY2q
GjEcGAKUO3YxXkziZKLVubqisWFs00zSe+myr+lZZUnw3m2piGXZMJuqUwswNrjJ
N8BMgXkHJfuL2JorzLLRpB8O2twASfGwKr6DQSO6s5K61WDgDYhakBQzolR53ny7
BtJ/ZE7SEjp6Je/UxFsr2CdOwxEyPzOMiKE2nkEBY+XLxsL/phBOdhEBk5WpuV+B
nwnz9FqT6r0hwCLgvL8CsLbtDjk4TrG3bpOPYy/NQiv1Vie2BgZDoBFxdnHiy3o3
JfNFoWrqENyGDvLy9BvENsE2Bq0GLEbtVMO0pf4RByneaF1xCGhIY6c288sRNt8W
V8syibSNNdx3OxwgnFeHYnbUq0ky7OrfTysy6wQ/7sW1YN+ZNkR/qF8SA1qhDSne
dNSZ9fc+Ja481xa+l83morJzBhZT/6fLyrSFnvy0DAuTWGRzLM3rP1tpZBC0Z+Sf
Z+M5jcegEmWpr3N3wCRswkQ6ePa01iWPUx1L/0FP1AQm1PJu92xo2ox+g4elDFvx
3rGbTqnpxpBbjtk/7D9ZkzJXTCb3uZgKIv7aDU2naymkM4xu936Jz9MqWyJ0LD3d
ZXWVJy3OL/v5lZKjIAlAewcdPdnfIggvVdaMijxAu/sas+0qPGJKrSjOaOD+9Noz
fbZV8Qd/UbM7hXymOD/U+EtUYoyWxDPK4LvIFScKDbN7QRezCm5E/1FrH4UeTyLS
S1X4Z9mp/Tgt0FFl++QSVnAYRuCTFTbjwjWAJHEEQSgNo05p/AIdyxgHJwYSYFWd
ZT8LWSXegtJaXLQeF5zNHA9n6/0W/UkIB4EHnIaAGdViYAgGvPfMujwZMrESNtW+
nXllSJuVx7jk9NFU+V35LRumEpNz6TEzss3GF3sS2V++jBye4j8VyOoBRGy9FOjd
yycX/XYiQJB64GM0lqPM8p66yylh0YWkoDj8awThoG4PvvOZBgbcKW6JS3wT8dsu
g1Kz8lNb1PciYFl0MVKVfbzu39NXmmG1nD4YZd/x9Qv4Iwm2MD1cNX3tAVoXHqeN
E6QPyNhM2wlkXSzLgZblthh7Jkd2uTBkvajdiBEdonxHhHu8E+4tRT4fcSOgpENf
p3ErLozpsn3ol7zyiyj5QYtJHFdJGNZYcZ6keLaS209bCp/bGbB3OwXsCFcLk6wS
AHXOm+ifJ2Ehn+Ovb9GSo9Fd2dNmZvJrY3+4QiUtrN2xNFAs2dojh3OmmfbPZQGA
ZskC9k3ovEJ01yzwUrptG10qs55qEDH7XrKuv9susem5XMrZu9SfjVVgr5Nmj/+7
1XqpeVaAHydk6cDAZ2LCluQ2ogplP+8BbPR9HfHUTnQITSN3sPl831eXY5BqOVV5
/cEGBIeCBLQs8Hyh5Gz4UchHvA5/fXH89B+1YIYWpta0ciV8g3Lwx8BpG90iyasS
rQB6o3jNoFmEfCtHC3JJgdkqPtdJLABGULE4PCKJcsqZOe5RrEdzet4rB5X+hsp7
xWuTP0VJTfyyonTa1AVL9/OGEZE4EZtG8zwAEure1qbyUKyJeZJld9u31BEJVzYE
GN43G21+/BAi3e2Dj/jGE1vxg1n4ZGtE1uaIhuElrpqMLYUrwO5UJkCDM1XDSytf
e9in5VszvT3xzKQdOy4/e8mjxe1bqTTbVk/Mey7bM5lexwhqTbBpbybHCOmOoEWE
XLzkl/X2ejFRu9r3ym8F8b5KsSMF5WjVu5NgsAetEv5cUO0Q3ZUOdPoG56pG4Nz3
Oy/OZdPqpr2VUmC4ynnjhfxFIJj36Dbq+xij7Z33t3uTA+T65dwgEKaJ6W6y79Oj
rWZsRv5OVWGmkzIwwazFH1PUjKwU5l7qvtcv6+MIrAaog7vSXMysviIKeUtMZ8pj
FRcPYn1npISyjaAksSDGH8ZT2nz/z8CVGVqvK4vKSbf+C1K1E72CbkkX3kQ9PDNe
aoyCFc55B5NZ1LvT+ntm/MrEpmH3BSGnQgtgFUElqFE9DOtD/5WuKe+VqyeQq8i0
YBSobDtV6BWS/ADs/1ZgwemJylbyF/FEdTUGLrnOvP38J343Lml/qC/XXPz+9XXB
aY5FaJIWE8Ax3p8TCnMF1IENHPHVRmJZKbAwSiHThEEDYaSrZC3S88Aa/LNuF2uY
Cihxjus6J1X1a4lkNZCpMrUIRjtFTHRxGAEWV4AViz257dpyIBzWQIQw3OOWQAEa
QNDBLSRLCuAXbF2L4NizwYdMF/amRrIxJalMR7XhhssCd6O7QOknwwWzNrytNjsu
Sw5tYgfD+va2zJnBi64+EQP1rY3YoiZyfPsRXQ3qrNF2tVexB09pczOQbUuo1CMY
5zdn6DZodkb4dGzDurIxRpUSusE5bJoZWnoXc1lufqlxyvz90hIkRRI7wCkLqNu7
4kzSxoZ5JUtozbJYjAKD/rNFLwCFrn3W5SvfrxNWVXpLELdDQVp2qkuU3mf2ZpPr
q5eqhjzNOnDjjkwQzGAxkPgTaVmVDLzxKzJSIZYo2Wk4kTq+PwAYYCav23Ta1V1P
v6mM9Rv2MWpH1k8D+DVZDqXceqrBQMFmjwuWN73nSmM6wSwHUf9Q4MGg0OfEj99u
MELzNSTk1So/lsrlYdDRuYtqNqNLgSZbr5+NEX1pvO7eYav2FSG7YzvtiLQd7eGR
Kzw/YfqCJOEJnQ/WiG9Md4Ox14yrgkz05FhuCPgmVv/WmMyXAP/qxZ0+J987w5GR
xwlmtSo/YtkCtyqInMAEYmQqIhVY8noSJlbl21Ltzs3BgD/Cs7mN2Sp1gwcwzijm
yIOcCq6xKjASBF5pj7S89r3ZyWGZg7tKmLyEkyLbBbjFgOaL8MBgr5riOPWIqMi+
Yg/jfel9j6tRQfpQsePSmvauX7CYO1wx8LKEsgTacAfHZErFsOPvI7RqmhC9oM73
e1pHuw5vi9++DkUNlOup2oPjD6NrShIdmKwmECxatA6MSiqn2PqAAqRgmon7kHky
NcG0U7zYHF6VXl/iLeDa6mxCc2qdKI6FBI6INKqrZvL4VYnrh56hZs35J/0R6p1B
M5x7n+UQfUi4pjcgfOsiXsSgAOR6tymPRDag8jyw4ly5nakYX/1xNPMwpyWNCNyb
zZ9YBnAeaSgjpnTP02oexdPLJlCiFhQZq0GJJpDrdWyNvONISzMcdwWR+l6tRVZ1
/d59CZBtEMQY6FhjWqfqpbCiRQV8BZnXz7n5tvtqpojyzkcRPKKPQcOGah0dy9xL
DyrC95I6VmeF3MqJShXuFAT7YepEsgloodyQFOjNHD05DDHqnxgOKywZPH2DCMKA
XQAQywkA0aczwmKjLzHr/bjSA5jqLBIbA0qV1kOZxLL16pScoiD7j3jk/9kgYEkt
m96ymrpquA1vt3iP3ulk7MnWAJFUuado7Lb9egT89xYKNYxpfQyUhcOc15/pXtgc
BUGd9IMRk2FEw7QkF/G0M6uEzrsBfRpPm6IFIEpFgC04fC1igoNDF/zZSwpcZTsO
j1KXNk5RoBGz8Z584eLy1VQ6zUA/Qx4jKKznBV8KcptdODPQx5MrqoESDEa8td49
VgNYCClwcmiW7ELES6X2TxWOddXCgaRrpqqIWfSjOc4hWHJlc7HT4p2/ljOtV57k
Y0cqucwwdn64WaiMZ2k1lDLVn3bSPscyK+L75RnLS79HpHjrjkuKbPRfCoKGiKRi
QcwEhls9BDtz1Oe725LSlzqcIGeswqBBJNAPpOgwex2KjySzqImgfXURfodqnTs2
38dK60f+XoppDdP7rgMn5zMa4trYOz18UtJwffNOU6pPBAcsqPKzKt8E/sRmDBQo
BZwR49nSPgYx0cx7fnb2P2QRYYfCe4k687J5XCQCuxQFas3zhHaPulxtAGqQdUkK
C8M+N1IEtqGZzUGkkUC0aqGLY07UA9gKQ+DxIGA7D61Ex7Lm0Sw+rXIg3U/Bz7pW
BJuPUXIJcPf4OJzd+3CDPZ4Chtpg/VxFrDOuGI/GddZHcgLW0D0fJxtIFQLBVgwW
3vcb9oPifAFAfohNrviKJExVfiswPPHVsRloYCYAkn74r4p7/mjNjUKhsUkxUnh/
lzKNK3sOJSqZ80txC52TYMPgmyjkxzdV3iSXUE5gNO88QEBrMi1kYmTm0/frXggT
nQydbSdHqfJ/Jlt4E1v8+b5jI/uZp2egpNPapBwvtdb6zYPrG9o+ff0MsfhxNKyB
F/51eX+y5FoONSj7NYzhiAZBJ9uNwGB7Paomjc3UoZK54aJp7qlq8D9ARqq/PXtF
v+Znc+5ZGwhZC05KMLl6M5XGjqYmNPUPUrrpRzkg1jZqesBQEOFpLRe06ZYIm2j4
P4kNbNiJmrGBiItUi4jufDTZ9L6iGPmIEqY+ZHzLbSJrCuYO1hxL0C5I9uzyDHdx
ZUMa4cN8qw34KeLxscJj6SSTbWwbANhdUquu397ExcFxZ8eoiSt0AljaGETlKEGt
pKoI+ZaEFzMs27NHd0FRQK3ToUsW7njYtPdUQYwhtxHMwibcsTAHneG/hkNG7adg
g9tueBCOHD3iCYVRTJc8EUPjCbFOmW2gAUX4q2WAo607NE5240TECZ09SIeNUKOy
RYSL4ejMA51GD60PEVQKrLtbBQzks9lJFGkiglGB+VWp0BHW3pQBAJ8+eX31KX6u
1EK7CtSSfBqUFmah5Wp7KAPbZbxhzxPoOe/nM9m07QJ6EFlYPcPDvZEKZR3Z2anL
E1MI9Q+sNG/uWiG2+NwuaCzSLZqLj0GaVOq3v5NIUiq5SHAnkJLovkY6t+4bgJHk
/y01ORPLkARJYveB6aHuKvc+d9eNeOh0UCp86DkBHQ2cd2J2VdsTZA+HUTZMIvOb
XZo3auQjAO9jp7GWj+zZvhltQRvzp+PYQlG4tDQyxixo9sesDOjkwX9PnyNf8krI
SCE0XvKNGr0ryZUPTJILHM2k5EQVpjYqgVQzKkvXtSkk1FYiPVPxf0rvt44eAdc9
mucvja0GOaMWm63wh7+cB89KSSDqJ0lkcGP0M8I8DdNLRCPB3pHgr3/nO6JbPqMo
tm+jXTcxtZ1wsuruq0XkmGycXJR8EHfZ0MpXqzQR+qSf8NvsoJ2GOLK8DTg0lvtt
cMQWcRUY+L2fQgJKVvkZbB/v+E4A/VqpqaPnN/kZHBRuK21HgY1M26KHOJXmmqi1
HwfvdihSAYDja7qP1GzsjWyTWY1Dzxluwoud5jNwN8wOzQtf5QKjIAPdrufeMkCD
1rrXLeyT1EnbGN5/fuYQHrVmmhi3vIlU/p/SjO64wx7zPzlqfnyzZH6MgoyGXLQb
+vHdqXannCVNLZ657BM+F3+0EZDukKxk3Hd7k2+9zw+wQOsyuWCWimfBPSH3m1xg
sokdGf5raiY/rBWk270inDuWeu/kcIZZaRRR4h3qypZnv2AqT76M8XuOzdZb27KX
wr6kzaWVXUttERg/5JnAM2pfysBLMOWOj4s7zfmYndo1eDVqGXalGykCSkPNdfPt
XYRm3y6Znm7mQlBk7IwQ3GJrd6G35ErXJ8UNQgRrLnURbf4fsgb5Bsc+mQxUj+wf
N12zPuk11K9HMDkLlGF6aXj8U940l0ryfnAq6nO9HAWRLxXo9ZRGi/enocu3am5z
yVeHIOoHyMW3F5PdlhbcxPBiOZ5mf0c5ZP5Lg1aR+gl17nBlLjeVZxH3RzbR4G3p
KrJ8lmScjf9ozGPUDJN2rwfGBlgKROYItV3p8BINZ9blvOWsRFO7qi9FXTZE0fjM
tCP/Zt9abNmLfTkLQw92cYJPLWSuMkalvD3R7veJnMDv8V3HET7S4vOKPO9PSxgn
oj6soJcWs2ppzOnqQXQgPj4oP+lsRHRWJSWy2hO3bsXlTrKgBaoC5ro2npEtRHWP
4hl43xk4LG+ALqGXM6XqPkzon50vyyWF+cYuYVHBydwO7X2mvk4XQQkn/wrPH7db
Ztt2Ivx9g/rEJSsVBRN2FvnC1PZUoePId1nNMDUKSb4lRYiFOzhakL0uWqAOrrSy
KeQcAaWPLD/CcA4KRUGbWizrmV7QQIxm/WN5TtzZZPA/oA71GolPbnjLkIPVET3T
o80oIRhr2r2IAerB4HmkfzoVtmL46oOPLxjkoNbTywfa6R2Ij66NG/i3xMfaZzLO
UwmBKw//P5JIO2t9hWMom7WuxLYMv9RLDImtk4V8NR5X+C3lBzSjRzlYSUJdEjgD
uYrru/edU84+ybQKyv9TvosOso1gCBYzbB25nXSPnu/o7NrIoZAFtvdLxjBE9dH3
E51/uXwDPSgBYcLYeMijy28KlQRklOjC5RP59T0ZGCxWfz3dfJo4UEdlhJOdDJ9S
km6PDBEuTmEzx5dxslrnRwjXAc+4ai8+qXuj/DcYQEc/jGtTh6A8bpcATw6J+zOG
TYvbr/IvSEQd4Ssjg2hWWb5E1t4NmLtiNu1whsFWyhHPIR3qK1LNGFLb4+yrQP/s
zyny3VIrSMmA6SgJLqj+/0MVI9eIpWsxFk9gGsNZD5ojp673zJlwdx6xTSGXH/uy
wRKtGU8tw8GjSgX4OzQnIEzLFd8JHu59f7haLJBZqOY30bRzPRYqdpetQvq6qTIv
x+rWTHgdC932/fdYhB5t0KPdIM6dPgiIKR/4O0Dhd0nrSV4RlviCjBCaoDth4vjE
Lrepm+clkIuq1d88f5UTtaN2A5diJ+JQeXComT6vLqnq9ZSm75Q+pKGVJHHMQAWk
SpnQbSFM48Be1A4V0nOmDhqfK7/CtRgQLyh848qnXpO4CWvX7AZfdQTr6gtyBJS6
ysVAiXyDpTNtR+NSoVgpK5uw9PN2IzzmXO9OOHGk5wBJhZ37R4DKC3vaSy9onNgw
/ljgN/Uhxhqll4IpBeQzM0S01ejQSmkjFVV6ic9nrpFZaNwwIWOE6r4d/OzKzdgU
MK6810oowjSgGdHdqM7od/YxCb43SCzXc71I5Ij0G9QwlzPwyfq50QIGD2tObKd2
kqfhu8fxb3XeK3VzcVRkoIo6T5vYtR+YfnOuojibgk4WfQVVtqO2KdYQ1/Wyq6ef
tpxXGTgYR8H7UG4a1ysL0tjeriCSt6mimUN2mG6myRC2UeZ6OcD9n/kmM0v2WJPi
wQSLDv8cmn3zt4pHayIp9A0Vr7ny7is1QZryyGmg3TP7iuhyd2qA/em97PnCtxtS
Aegu0tjq6rNSIzjUitutYlM8fqZK2PB151wYhlezJXuIHAYsGR/ALXnBUUvImDSw
DYZWfZPzTtujWUD844VhIcclFo+yxjREwO8JtYjgGSDNv8qFoBCZOHrcQ88GIowr
YR0VAHPmXRhCZoP89HQH+IIiePqZ6iesq52SV/7slMQd6ulENG+N98+oh5Z9Y/vm
IUS0l9W/Vj529JRKFWLl0mP8Ayo+FSJ7ywIUWc2G4v++ZFHRh92dPJ7LOX4EGwsc
ebUo3XUbUapYTIEQRwtES944dmvFjBx5dFk3r/ht55DoIEs1D0uqMUbpvk3BXJ43
kUe71hpzaracShGCNT1JSHTc+AMnkUhD8k3tXA43QiFmR9N3RYShWi9H+3ui3hVX
lDli145/a+Kp7FbsCEZ0SO47ZdrSy9/KRqbaVdQRtKNa+smBJT3zc/4JkkZCLzjm
8uv6SBrCxUbxXoGqs3RBnAlUHSZQELOze9W9BR5Q4UTQeFsr7YkQI2t2i0kjUTLT
cGHzLXNeTrzyk7XjY/iif7ErofAppAWTQD7r9hbLI+p10cxDHfXy6TkizQSFnICT
sV+fP1xQ0U65U3fPu+8Y4Wi9ZTGCEkU2stcRwHgSM3qroM9zEHxTXjYrD6sQJLq5
mPXu+rwJxYYwHpFShKczphc4U75mbadThVULmS0Mq8QS+UEf+6FBPyCrYITHq0pu
GvMyyj/rbGDPjpPYyUpP0HECO9gu/ixu61VGw31kzqPjKgZHpH29zkTdZ0eYAsNl
7oeLa98BGKtSGHG/uG3LSU7iZo3/ns+mK/MFyTLLNLpyWc3yxuKElu79ad1wPoDW
4pl5q2/zxztWQqKOihq5I1DvF18305tTSk7tnTgo2/If/bdGx25OiaYz6N4z5dqW
ZMH/aCqQRuDid8srrMdu9BzNP/WZZ2S8i4tMhduOSLJSwz9fZebqFURP4K5chrF4
EEwiBasBxNPjVS3BtZfHzCLzKe8EsneKpoWQL39vG0NIvDdsZEM/aV5uuvdE800h
HRSF0zkltk7OfvqUWCl0grZr05CjniCpfgM1Z5U7JXe2R0BvfQ3IHXo3ZrlJOq+p
j9Oz+PpU4JHRu2JboJ4LhwSdrQzsOXlYtuVC5UrADjza8u+u06Oi5xCYB9O6/81a
Cv4eji77VKprbMo9rWKfpj4yffZ86XP5CgOCyZitvlkXmvK2McutT2UgYpv3ZuTD
/WhEPmipbMEVeLtho36BwQJ1x1hjVYzOa1V0N45KC4POLzxUISJp/M239Kefe3OU
OIo/aAU1veMtWFVFAcTMFok1ClD7miJ6WpwSUrf9b+/N9kte8tJvC/NJo9YZKkH5
8FH5dRepWmEkZqu3u2wv2huGr+bCljb1/AiWdrFa+LU3dcID2fNELFSVuZk0enNW
ZDvYbSbl/OHLfljBx4/wfooLfuPU7kQAEunXLx1ipT4rtpmKf28FWFU0onH9i+gw
8S79qQWLtE4tTN73DOTlUUUUw04tv5rSvRd650zINleFej7B3fFCMY7lTM5Dmcp7
bL+vvoFICX0WVkl4y81qUvbomNi1xKod0e8Am4ecFKtPnmUJPBEmr5H/urG6gHCD
Fr6MB+uqyqGJrKksA6fZU0fEApi8832NQmYfCXtZ19TCVf7fLqy+mHOdmR2Sq1IH
NbP17UfpcgO0sGe9yHOwexwE8vF/Ake7NRzbd7JkX6KVTon6CbjsF9pwF8/I7DJX
83P0XbSKraczjfwRTjNZrRHATiL0Ph/N9/nKhR8pyXstSNrdGF3iUxXz767LW4Lg
MNiFpVpdY7pAcfZNMDuGV2LInSdSIxqZoQQERR9hgLaxzfZMBdNC3Es3phE5e68d
6mDa0bcpDwN3Nk8i3nY5g1J1lcQKrzKt9kR/wUP+zDDm2Q9WT6wB8aYpl/pDFwf2
Y6UDJ7DRv7YKjOekOopLRzsYW6iqyS92HS9gW3G+wk7Ezk26s3F0rqcRK3k8IX0t
DR8F+LV9UJkZ1GJoDBRBi84vcjz2+0mgk/6BwaJvvXUZSxAq6ZZFs2TuizXXtUB2
YQ6aajAueDT6ge7NctwJLDsCE8RwEbJ2x6xjpLUmX0rf/TrqmL61Zu0u0iIH4OPw
GWf4R/T9A6bLgtKzJBl7V1fLvWMd0PbILpNe5DxLgFullFhbd3bktC93FwALX7/N
jsJC/2joTvw1XDm+dZS4Dck+7UQJVc1n/uwbVa8m5HfDFmPK7uESeinNkysdztn8
522Xg8MKQmUKN1MfNaPzV+y3opJECapziypG70OxFE03sPJDXWMdtDhHfv8o88b9
+r8ZVEj/ltStyACwuhGdMbLgBNBYYrjiEz5HxOYSU8kW5eGPMVmIT1Yw5ZgieSAS
QEO5NZopoGTVjYi5dnTNAcUlKuHdnkTIQybGZsNwtBgcpojlLCNLcPnK0pzoDq3r
YBm1rjmEDv2STF47/diGqMNYZKG0oug2uHUnCbC3ydlQZW9Njlt5fJ8PVM6H8oiB
I5X95wHYozRIjLHNaTHzZAryWgFw+3kOp0bdgeHvZADXWnnYxDhslLF6WomKJkIF
tSd1nYAgvgllrDpZEEYNqkX7LS3Z3DTznEHGvMLRgnP2bXbQtKXfQeEDm2kVzmJ2
ZLXBUDQYqCp02Oav50cpYSl516TsRKO4hsFsnBX96JJTGm9OYhyymCSrRAmzW8Du
F0i2BYsJOJb3lpBlRObmIx2Sy51KFpM2OvdIgelYeUUCbUx+Azt0ZbyGNX7usy4a
lDxNFKnvFE5mTrvdc32BjNdHPDMHUuD2py23ZQzO5y+d3MWL/tHW6Bk6DRL3RY0q
DybH4PVpD9mnqPpT/xuYZUGo3+5FHHw5Lgds8oiOpr5mGNkB0euEGKJ6gFX0FNri
ADBP4eBuUyQUywTmr+fIYi0hm7KNgF65VLpw7Wn4bB322ZKn5mKgo0fQbWCFqMtZ
rbvIcE8x6r7zM36sLKlZinAjvSOdnTVqFHLuBuc3xlSVklROmRzbq8kmDc1AFlpJ
myA6NK1pP0smJtLLdvoA5KYb4CARbxrsC4ML4tINMmM2duS3zZhLmE8n6IXeMMQ2
vmaBhnDSHrY/QcLetH3vB7HD7Y/xnVsC73BDMTj3MP/SXCYrqYvWbqNfRvvFWUKa
CgMfZVxzYpKOhj5dvCSBwpP0iNa4RbN47J1Vr3PMwauV+B0PanC/Hs6i/SNuOrZx
Ppt/GoYGjSWOKLicPrO7YZ4PFf4WVebyTm8VkBUyMx6/ToRukT0PdcvZVAZ5exF/
6k70tQghkQjPIRg03Am2CrxEVRDrjbHKBoqOfY2i/uxIWf+09EoeuNtsmPCXELLd
x2WD51pMP23E/gl8Ox89b8+rhwZVho+f2BT39fbSFJQFeZwPOx9h82K4tKfzo38Q
mgUfOMFxgYh5uPpXH1PzJQRqw5Twa/qC78b2qhxh/0TzcBPxsBdaTUgAWq9QTeBl
Sm4aiPj46vUY6uyANHSHgOzUM885LrPYatMPmqmJKBJ4Esun6twh8weBnBymNJH/
udwCj5oSLblkIpQo+bu17TL9lD9iJOEeW3Fpv4HUy9v1KuK4zxrhnaJ2Crke+E0S
IY0MMO6xHjsG0hTMYLlQ3chpwhPQJmAKY1ADFYLN45lgJWX0jhUdLM2KdaYj32Wb
mm1Mba5dc1PXL7NIiLO7zJrHrCWE/AK/LuNfOsBFyNqP/xzY3JO+e62zuhTm1obi
apoF6bYAhYw90BnrBekJ6qFy1GfKDCniDXhvmU9ogfQ1fQpeSiupli391Y1YNiQJ
mcNLC8N86NXjug7XhaOu2BSw6SxXx8X1bxjCuv/qk6a0KprSy3a09S30AbpN8hWO
6pRbgArM23fTK37ZphVUFaGsKBmYSLnnSIjDB4S9127MReyMeWLnG7Hch7+12TL+
nMBgHbW0PUjZJXAF38m70XsIQ9NzgQOq36fEYoV0TIbLeOr0hK540Y4NvI/Q2D16
Jp8k+tl09S5G+IPVaZMExd+oydrSbrJmPbhF/sz3YAk9xgZzE13Nb5YjMHbJVzAJ
/spTI/gpSVfr/ae4OJSDs0b0lnYbTADwkeqhLOmAA88O8lyt5Lwv1invfg3SeEjK
V9kihcynjDQsIqF0kgX6VNcIGb/IVs76OibOHp8Z7wd5HxI5nVxbfKPorQzf2slF
GVFAOS/T/xKmGXRyVsYG+s9FFI8smIUbMZtCypKTDjW2YVRVPZIk3ofOcRuvXPqs
3Q0zvLNSKemL8+oOVSlWx7PNt2X2c3MhOd5qNO8naNWhb9gMmOQnK+A0JkdwS0xK
P7Samyv7/CO9ZBjJ8ouAxQjKBCUC5hBqR8KCk4hv6d8DZoH6OOAlABS5IKg89si9
vKKGQ9GGyulH5cIaKCHgsa3finAFKk/03qxG3PB1ax0wXocO/tPlqa7/3VrLYgq5
3+BAi6FXf++FCABygMLap0RNWQwwMJIpMMducThqxA2mE6eXtFpf2gSTciJKuT5S
tHo/ruujR4D7TZyD/oq6QGK843pXGH2VZdV3cdVy0P8r4Ggnhgw2gTi1K+REUVdd
W6EX9IiCuQOkI1MAtJK4/8bXsKtSJr9t/OI5iwME4jdy0XD+UArorzGrPSCLLpln
G49mK8ZE0Rhnz98NjCCCTaBE8VC14bp4PMtVpXxRFDEGsGd0+Iw2ThOh7nQ3ZtLF
yhhjieUKwVTcHfGh/cJoxPPib1nnAVJPHLUqu35JYXw+uN/NQzetVU13114J2x58
RQPLnOrhP+IFtJRTeOXpRaY5p4kOjT69I6WMInR+AzAhMtwG9OoDwKl3zIPgKNjZ
6VRWKMbcKHJP0MKfK6ZP/JYORWCKZgDb/a8jieYX8RcDfCeZATAIePQ7689MB+gL
nepaetnIul0MzWsPKryZ56CcjaC1lsT+Rq9C0WXwnbKm/plEm4Hn/nhuKd++4t+D
TQhYjLNszjJO+PX+SwxqUSnZF983SJXYXLCLunwcTGoj1b4PKE3zpykKOIObKhEr
oFdm66J9YqVfIhzOfTanolRSYuBo9+KCoOYxc4+IMdCSncpEXnJ/MmryYygrUCs2
+dbh6MYjHoNw9z0UAhE45lkYzJn8fEL2UU9Bh31Bn2b1w7SgyffQwru3U/nrTjon
VKQtidQqY9ZmoDd2P4g5n6kT2zRKROz+LRCweGcC1HDF1tTYAKYoVDNp0UMRjfBa
sd4gtOzcA+qL2PTTRpfI+9BA8Bdm5TR7V0msnDIGnm4iKKcWoPmGXpa75YPcR3Zb
NV372eRBxAG4PxLhIJNkgOrQxwhAn/BWWg2xAfsNamacI81ifPyj6/xbmjXnL9Sd
3OTqRGpNBUWkuBClhvpRJ1UCH3aC1FLYUONgQxfpwd3CjoWWD7L5tlXjrrG0UidF
RPeVjnMyxwWXmxcZIfkF37iXc4E2Y9iqnD4Ge/tChyE8Y7ZSEVBBmYPGgETTm6Oa
6j3dIMxmqrpFx1h8p3N/QSoM5L+ujA06pHAU3zReqC1h2DQ9x39MOUIe3R72S6Zm
GLOpYKNXBWnZ3rjMy5dae/DqfWe1lDF2vfwd0Vxvb2QD0AZ4WyFYo9jEEVZrpeDm
REAUfGaZZZp4UEqX/GH3y3VzJZG+tjncbGTa2LTHsq+1rNtSINf/Dh+iC8DvulLd
POyR3pv+fOw3vq3uCPXWA95v+mgBeLo53RNtPTu2nwnM+4MZnDl4mVjZZaCoFnp2
NT2Tg5auigmm8Aw7Dywzme2iwQhWB6rSEbNN1KBRWGoW4pseu0hYksLHEHV04ufZ
rAflFnpBisTxhn0CF9RylfvcPKHS8gXALDyKr+FTkDWK8MfOszIFoOeaLq5ZmYP8
ZN041acUp6rEi0HYls835IALji1L4Za0I2ydunAkqY9SYlkULEmyMl4419f9izhE
hBFHj7PHKSF3SJDWnAvO+jV9HAh6s9zWabP060Sn45UlGbBIvgIzGW7xKdvgdK4f
Ti+H3DOTNHjmzCyIRy+tPH/5b0nPHoCGLXXm3yVsnOx9brJYyRFNccq0sx2rn1rW
FjwuNgeES7XbP46edU1l47+vhpHgqHNifDCK5AAJthFMFOZMuANwlr/E8NSfl9v2
nyYU5mCi4fmL4hCCKs1BNi6Hs2ce/ywRjx+IrO5iN9Y8W2vjZscZJCwCCvDHqjET
U3gANdC/TcwuAUAPOx+AWwELlQ6S/g+8RWUvbhzUtuRciCKp0w4mwO+B+LsHFrVy
ga8r/m/i0BjqiGxyDcwAXkpcHEZom7wwGUrXnbN2ykf17gO/cQeJr3FTLFfHCU19
wGDTrI1RPY446YfGlyZmHG9gE4cOWu975vYvoyKdldG2AcY78gT89K8085QSd3vV
+5PjWRVPIRiUIZVHfZI1llR8l/Q5ZodxdDlWp9p+OXjS+hY4wqPsTv1pJ6sZEn3V
DBR6x2JGniXr9Vk6IXJofV1T44gIxzI80eNg/mPOhPM2qcyAAV8Oqk4DGv6InpP6
SFasUXdiQNTuQajStSWv0j76HVfT4EPfbqEzZO93owsZbB3jYwhND82NpjNoY+PT
77iU2W8fqvYxCeNTlQA9cMNp6RP2miFdpWg0/k6aJTIngspaHIvU2NLjw5EadVl4
W3Omr84f/rudYw9hZ7GW2kLF1lT+Ce0KWik0oBCasprDDUrokerLlILCOuAvaUiC
M40ZuLXMqLAtafHCBAkmnl7fhHG4XQ60ag1j+eZ+geXz6Acio6CHtu0LTZtMigKu
WYhfLg7d4Fdk5qWT+k6I8blW/FJPiF2+YVcZZntETspHp0TPl5/sEFrSEDTrram3
l4hp0eu3e4wX/+5MU6bcDdAaaSss40TGUxriI6y9ewBCdMmpv18glWieP2ELHf0A
ikLGbHZDIpT+QPO6++vYFk+2TmNTWN90V691QENCTBkoQ70kXYfxYSj0536BZdMx
it0xBLVkqSkO2ApKZgic3aIWGoirU8HBCv4jO1SWH6y7cWwhudstRCF1aFVMS48g
u8nA91Xh654BivlNo8v7EWsMDnn409K5rfnuAPRuWyubm3wqoz6j4JW2TQnc2bqQ
kOTIKWw0glr7R+sV0T0zRfszskROxHM/Ysgm3h71Wpd9Zo9ECS7ECQv5/Tc4HpBr
WIOIqDvzzbXmUXFXeOuADp9LWF2UfQA8qP7VPV/I+GUvZaMupA+AocZh7/So97uv
SRiOJkfrHaVP6h2wry/uTJJcdX/mG0qIBr92cCCeoKTN4RzX4kkrEZEPjOx4G3Fw
0JDF2rIQgoto0JQz4PP0jlXGKQbt98NoecWiAFHY1WZfz9QgkEWlO475LSgulL54
htNFP5Cgc1vxastBV96AFVBv/LcY5f7S7XGX9WgqrXbd9acTJ7wU4d0FL4uyP+Y+
BWtYyQVzu7S1az3ZimAYMqXpCk64fkmc0u8lE099mawLWbNLOW9kyt+cmA1gHjCX
H6hFWzYYjcGyyPvFqkiL0f4QsCwijV3uHa9PtR7R9JDdnCbouPylwxCSt3Zw4YGs
HRFE78ERzoDaYXhMvL0UOHxgZt5v7Vqp+wjYyuvMbUhCBAHxVfGKVYyWctwhVwQv
rC8boPR60LCzL7KJyBy1jMiOAOb31AG3NBrwNTpVgkyjW9KTIudUWCt+BGGFzr9m
yROlE4YDnZ0r/VcKrH9bfACPBNmSmPaTVDYYNvK13jLfZvQjIPjA2uhABvXbuwD5
ojvZreHq+VHYhu7KO30g8OltCgtxF32yLONFgfSrB8mtlj9E/eufuTN9nTnzV0K2
WGpoDAdpN43ioAlJZ7h7p3bPFqtV/4noqQ9rBS+fZPGeuxcCHjVYWe3cJ/TRl70B
gn5wZ8UGQmehkAL9w6ZdTdHzjTsbJpruw5wtgk7MXjXPMeHhKyMpgi5lsdq6bF7b
genPKqs7MpjvVtl1Yt0Hn/ZUezxSA5OvtaoBjTaAbrCfR57yMDWRKDt0P3DTzZI2
xfLUeadRuM1Ut9v1BlNIJaibNwYQ0i7rrah2jXEG0lu4TNPd0MrbacfHNdPuIcCk
9S1mBI4RBUfQ0DpbqS2L8O7Ts+L60UyTU9aAkKLKmpyCZkv2bR67Xidwyfe7WMnv
smA5l1T8OXVGmP50LRqKm/GMw+I1WkZ5sMe3lifEuS3twBKyRJ09PnHwf/DLgtZu
pJucgY9J0V+5KqoDIkrlbjMC9DqYEq0T8+kMK1UirQdnWdI5hEvoyGw5oDPS9ZvK
5Xl8ExPepp5pyy5o6VpOygDFoduwatCYBKScg4E2pd4S0eqJNEgaOGogDKqn6vJV
3fuxvIRpCmWKN09PrDRGyYgeA2CcthK2sOfDXfgZdcOs0xMEP2WdSahL9SqwOe6w
ZnEdWyXj0ZntSBSZnOjxcKkAi1PLtXp1vqCdJL2LL7Z3Vo0D18xmEkLq5qa6lW3h
NpUVmyY/pdXROofWcINjC4wF+LDXinpAM8GFTJxED+JI4t9RIzeF7LjP0ienaH4k
cFV2I3ZRE34XfYpLInDdtj/LdonYFiPa2APXi5SdU/sDOWzy5zocHPX0PlLNlOjk
4cxfSlZ5/TuypCeLZ1heriZpQfKW0Pxk0HdoBtMo2BYZWw2e/1oujsrQEDVjedco
eL+ThyhyiyBZgyMNIuaHLeSDSJ/3oBbRS6d9GtV7Rquk6NxicF5FGIkqOx/kMk44
xpgQMwBeSGWsmVuJC1VGO9gHXvQnin6R2iJW3MJmDGWyp8f8vGxSzNwPl9/ky/Bo
dxpSryCAMap0Mc3K76CJJDKHLkdMW/vd+/+1ckvLE8yGfDaoOfzMwYHOcRNz/Zi3
6nTu8YAJ9hC76OHCvUOqcXUH4PwcqzOoRItSvQTMn3shYJpuh5tYeUMiLsESlsNL
R5UMcTFp0ISmnPe83VMnJjAbeHAQV+pZQKMN9MUIbo2P0kWHansUbcjgJzBvrIBi
9UEE+Y/q+fufB29U56LuvyKs3FPNfRtmbUSRD/vemHu/p0ljowGQVPhFHKhxoMoj
W6ecq8Pe1U0h7p+Z8lRvDGLo98g75Rffn/Yq3ypZYdyhwchrJVyu/qu8HQYEQhC8
Kr7R9rUw+OKD106jBW5OwEx04kxwu2IgR0AJe/Azd6NDcME+PgiwFFjlzcNjDtFn
blsVWnU9qpIGggtDZq3sZye/UkH81ziUIH4SDkIN2eBQcpmxJHIaf+dBAxDYiR64
nC5GO9OpQD4/3H85FnpJqA+GbSNMcvxQVa1LfeksfVkHZRyHqFwtf8NAqWPcBhBU
Zgc2YE22Gf+pFSOJW5Pk7xn66DQWAP7Gt7iOBK7NteYBZOvzG+Np4FKc3vYc2FOk
VbFe5fFiJJTGn/bfDrFsxq5UQ0iEkCBnEOY7erJ+PhYbz9qfDvK7ZkZ6Cqj8o5RF
1CScjzh5ylefTsfsuJxRGNWizcK3fdWoL9uyP+aH8y6bCnkpmPFtQy5gRthb1Zua
w8JtslSz9krODBrtCk9mTOqFMQDVmqksOrYciax/U+cmV0IVyfAAUD2kqQd+vWaT
sQswC8ZX6HPvXMGqRf3W7X/DwFuAXCLqa4/zX1QCX4KHlsMRu4zx6yNStr/j4N2i
FKm/PLvQ8m38pCkpPAe7DcIptk5g33cVuNRG6QqHWCDTXrEjac0f7sOI0C8PN+RR
LWIgJcT903L8ldDmkq8dm6ev4h3s+p9+395BLCrp7z7jUVNi9+WFW3WAQRd6ueY1
YDthmMtHG+22wwEtCkQMdWMosW1ulekLW4O3x8Ih1z6lpl25IXBAE6VVU/9TREjI
F01dYSmTgGdVLEIZsHfc8FVMgV4U0g+ac2QetK97oW9fDr3t7AxbHj+uAzKOGsaU
aQOO8eQhKnVuWySbT7ZtsN63hR+hD/pYzxrPNLSdt7ayCXUoJtI3G9XE0tVQatn1
czud7X+heAN1L/4gTw0ghJWjYY4f+P2Mi5PrOP77Gay7Deq+F4ZTJrqhFMmM883b
W1CrwnYJiCD7Oa/FRPka0eg3aXsGQVdwvbaAmme9KDh2X1uL/2SSUbqd0m16J/E3
zmkRywRjzDl2LKJWVLXaFBDEvR81znBCY5gNemgg4xZTqvdLQVIkkmlRPRMNFfTU
uiLtQ9evLyDD48VmjxEeKnqfmPRcAx1Hs/6CwYENF/5lJgs8Vy6Ziv6YFOd9+/VZ
Y+SqjVjdfZi9PY+q8gTxFPpeVVw+w1Tkye6U4+KtdvwZcPly6MGMQleODJi5pe7t
bzxjy0R1ukiFLnY5UkfE/XTRw5JJIZe31RgzaF8OqlXfA3GkBjjJu4vTH22rJhSi
jPTTJnF3hwFakIEPX+A7QDOj72RPnVdai7ui2DCkuucPEZQ0yRW8za3nFYBCASLF
Zor97kHomiCDWoaI4WwRSPgVN/vIJqup8jf1nw7EiMQCY/wMxh9RJW557DvTjWJ4
DM9Et/OhlHi90c4mWhzWzQb8eaSXwUuIJAk9nUHWebfbpPObDKIniHPgQC2lvUMa
Zay1tb0hdJnMGSR6zqEhG8NhObqsq943BBRynLSPpKdDs+HtGck+2N0QUreJhhy2
BmUVkUtiTQJumTsegH8IUUJz5tHEgGNzbZKaWjRB3BQeiRgHmeIbj7Pyi8HcaJvA
SMG16NRMcPVShx7qRTRz5PKr0duxqULlxCNEQk54THqmIJo95IIYEVikSQkIdYda
qb85WLFJEy3b2bjCkrDZKq/Xd778yjPFq15cWJuyAdRupdp+UyYUiUCfYCgbquK8
tjXQdDIBByKIcL17Wt0dGSa5/iAiyF40iQb8PtfZNDZ1j+VG6Vlgbqdk7PbS5bIZ
6uvOldNro4CgJbxgO96gGZ9PDJRgNg4qnp+tCyO37TR2nkdjt9yCnsH+3sMrQuGT
6Cx4SFcENFJK0+I788gXBYJ3lTVQZeytJTTF6r4gqzBY3KEHVLo/DyXBd9EiSRan
Ik8PVDB2658Mlbjs1uFupPGmbKSXG6IVj//wHTxZGz6xCvB7cZLM14lKjUl6zts6
xTqgZuu06ShZNCh3v6C6XoYj2s0h/68R8p5dlblClPfesW3GESg1zeuOW+uPEBzm
6JOqcaI350YcGms8QnsGmwe9AV3fOyZh3jBnMcEWRXxUA7tnBM8j6pF4fcLJp93j
VDzsBhwqde//gf8otiHw+Tt9oGoZHMBrs09Ohv7JHRB2NuO9Hrk20Qgaye98oxNZ
h3v27I0g5wtonidUtJ73XtMeLO76xVROLgBNinb0MEBGlvads+PCFtzZ0gchLqll
ebQLgP9PnAvc6qeQPNvdxqV9Shbv6Iwj7kB6gvpe6J8c+oush6wj2WTZ0iYh+XUk
amgf+5JGric+zumLaEaR8KTFzlRzfbb6V2znrdbWsYIy0bnYSMhvg21rxvwdkiH+
N+yXiCvwu6IeWUvIRLRYXQHYxSWXrFIZHz/bqvIActfzL1UD2hqZdGD6RlpQILai
RQEdhGu/5px3oLHREcJIbyrPEhtfvmeYM/V7vaiQT4BHIYyaTBHOgAdGpRN1w2q6
KvSxw5AD7W+QcTlyRkyPy4u43NHcYUHNmuSMr03ToErAabLUAA0tFD3D8T+yX/K6
n55UxOKWqkadNPWFdxqO/8E7EzRAiCeuYY25M3qYXm7+j+iWJrTG+YovZYPBQLzq
+AOS2uYr5VaPP/jsZg1iYRjQ5/cMGW7WfxB7TUj1O38gzozJOB2ZPdAKpkCKPvYu
srKLKUhL5iBYB4YuXRqpYRLJ9Bf1hvhBeTKFpFtAVtW4VTRegaus3w6J4mgakteE
Vgt9nTlRLYC6Q8MdyJejjJmHFqq/swXSK4Jrrc857xnJiWxtQXnvFnc096tGjuu+
u1VOXY8Sp0t0O8t0zZIHR/bBm3fZOkwKnbOcwYosyYOyj+iFVMC1nLChYEtOwmMT
CLPYmLXtNNmt4pFvGcKwc2mQ+KWJnyOQDriHuAaZuSxI6tNBmNHjLdi3VtITmSH0
mfyNQ+CGe/lj01Ui5kp5/e959/mO1kziLLpNRDX+HIoQnlM2bGURvhrbdM7imJFi
QFvnsAJ1P+zsargF9e1ZfbFPcMqXRLZUpF4V/ReaQtDny6mkocWz0qqUPHVw9LI6
o+f5jrmkyB/Of/EFXQyg8DciBFFeG36IGLTd8I3FueOTdchH7sMWNCYpkdu97T+Y
ab5W2JFscR+IWcGLLh8Yd/fgap+m9Wx4bn5Bumm5tywcjvE+/oKolUo9dUFCcsoa
lAL91xeMLC8L/iB1tj9aod4TYDZ/rKErDU6Sm8rPIxMpSzkwlrfyport+l++xWVs
CXP44NfblqP1K2gHadDIoSebZ89AQq7oAnk2L8LLNI2r/l6WwJ1gZXIs+uh/g0JY
r47HPFss4u/GCPGUBDF1MneEFbl/9W21BPQEuVe/LQUsVmsfUs94nyFcfF5h1dsE
YrhGTH37HaddOZQAcMLvMxda2W31fwy48ZJbHlDVk56zThdpgqDh8b1w4sYghUKu
6hRMqbP5zw3eicn7OTadI0QKXJ85C+fJ1VDege1SxEVSXa+x0WpwWLuRSKgnxuDT
7nHqn8N6txasgZOlT/KONYBaZnz1muQSulO1va7kbrhMcUplPQT5EXyqZwMnqMdz
1X88X2joiH0s7e7Uvz7peH+KqQ8aR4i8Yv52f10ejvx+LMIXmYX0I4U8mBj5+msM
wrz+hL5Y6eFDzubBbWRWS65adofo0rcC8RM99fKWQIKkaMSdUSKwzb5h8Q5yqj2r
o7vQPL0nFJ7ogqLUyT2xQZAwibwoMs6pXc++me7f+owyJkMxPP9sNp61tb0Pudoh
0NLbsBhv2svOr6fZKje0d7aHX0mFLreYNOGL6t2wO3J8PZmChCBq2YqfAMwX9KwZ
oKGXPhvoAKwKtxnAKPzknJ44+k4guqK8QH/mvGxYByw4PgVcw5UmA4oMAy+7gHri
KanZSXYW0Fpjml+ekEFax/EOYk3f1dVKdoMZvkytNOE5WKRctOh6vy+COhq81WIG
F7E78oV9PN9tI5pKM4utXQMMI2eICcNkS6Av9kbS2glrSKXJHt8cTb3dSesLjE4L
zTmWWcfc262jmH7nVJAwQUqWqUpkRFew5+HOoB5q8yII30jcmMBcw0ue4oUzsAQ/
bYoV0h2VGAJwKl23YblH/cTBDKNhi9CqYRBkMeZ5InwO4b4YXOVDJXgz8DYovAmG
VQMrtRx5jCYd0pjW91olOB5H3d0iWnrdkgeWwDCfa3w5dOzzYEeqo0VEo30qCxIY
BYiqeIs1ya8SKJfp7r4k+XcHa972f6UwZ7fQMH7f3WjDWmZcgyVzJBSJJNjO6ZgT
aFwKiZIN2V2R2KO7eGcjsz8uC9ZSzQn+WKZHl24Fc1CWCqz/kwDCvtQ5PMe2Y83G
w1yDDvO1TeIUGk6zTsjxCjjq1vl7J7lgypE65g9YLdk1VXj85qcpnCVGDBDuITKY
wuS3+8JEGw9JwAohbTnyLP9SMvTfYuzinKik03+hWl1+EHlWfwMWiQiz2vnRuEBQ
198gzLaY7AjXdL9dR4iaeam1XPayFgmwDltPQHOh22nDCGMxKVEtUjPYYpChyIAq
WkGto+1hb2zyAl/FnGAOaGgG3iu+fgoyg6Zkdne6pBMoW8BFf//aEfG/zTqW76TY
Hr262w4BEQgnGD7VSCLdAFAxbn7oXt5iY9Y5ze0qbMLyCEAJZVSN721J7rjmqvza
FpZvyZ+bDCntSDeuh8rfzptbjEBsQfpo8z+0OcpVasEXlHWCvCm4Uy50/EuqPLVn
Gy/yVcyMLXqdkteEhQKKLsPm32m84gqzVggC9kNXXAcZJwSxfnUYhbafZPqBTBRd
CtsgICZkEJRgPCFRrbvWXQtztKiTXxH9STBaWl6Z13PuH2bY5iESQUJLuWCGwjqf
cjh4BZ7hnMLK7v9Ton2CmO0sO2qCU6oBETM2ldDha4FVuCNLXFumqVwb8i8UhsdC
Oy/afCJTDaxgwdZ4r08r4k/OGqWtqTx79qnFJAJf1O8r3ouSG7otA2w9BW3cCyBZ
tce8M8xbTaLn0CG+CmJcR63MJjAhPl8Dwon5wkkCz9k5yRXllieoQ3QQEB63UP2/
JjXnvE+ElObCQhxKbcE+naRIg3CZ7cwASGvvhrQwkJBoNx8KEwJBE0aOUkfYRUe/
Zq3qOAzWiXpanNZyNioRzRbHRsx8h0NdzjAT6zOCejd/HCCTD4Pq3IIouYTTjHD5
K5cOqAWfzAJGo3Kl3/pD2vzT8M1G0mtU8C+9ZcsMwJNjczcMyQ6zlJlTs57SLrFX
4adDDwHVyCtyChyIYg5BtaIOiDII/raDmUmlaBV9YaSmkovi+WGcMsb+RCrWPpwu
3n4uQgvjgkY6iq73Oo1/mMkEkorMIkmAGcJTmSSRPm5EZGTJ3Y+lUe8yYmyextk3
T/vCQpcVq9SnKz6xmwrl3hvYaOs8KmvxrcNhYkOqU0GiYoS9ArnyhqpdRAeADNTG
3i9YvI8Cx/hMoygggieTFJ5Yvjm27JZT7UCZkq8PZttSYT4jZND2HFi6w4eMHgvO
ONxW0ND8dyRkyxSpmN6SLgplh/0mriUhNlqCcvlVyHfEGJjNwFweYNsJcvps/vll
zYsJyJHOf5UltAEV4q7w5hcw6QgUxhHCz7In6uGQj7rBvBJUJYoGbtmT997quw3u
wNoN1uPqz8i3k6ISO8xgiak5oduaDPXwhkCadurTDUFOGwxWfBIDTyf3zoqOSnuT
CGIhw469BrQlxX9NQEi8E5gF32giANUdirXVZoza06tzdYC1ScKuzOXFCPEfzWJN
ycQLfbB8CpLHh1O6AY6VwQBjA+L7FHPr7R5K1BHbNItIeREhKIBubZalbz3OhRMw
VimJGFSxtOZT7zVVVtzGSuRLWZoKPyGyS9imCFKV4hTj5OJc42aUFjWR3QjoAtog
CwDHbzypuU+qCDe43BNQT5vA0d2VWvBagFVAEKDZz+jJxUbsxnrwqqMtK+RNLfQm
TRSDVriMWow+cxcpv71oFzWBWXh9uMFvDLKZaN36iGQi7s+ecBbobSAfNGuTt+CA
18oHZIBXcPyLSART/qzhuFwOyQmDfnMafIe/S/LfZcuC+19NUYDJU6PaCIeGrDjm
n2//JSh7oj1gXOlNV83jywEohvJFGN5q0tuSdXUCzaUOQaOMYLfXCwUmvwmRtump
IBnGHNQ7kq0iJFSA+qydPiLd5TFZ4/gNXKxkbOkdwlO18QstbL2Ukvcta3gz7iHy
Nmjdb3d/uqPnSQsROfkj9y+MRnyYv8XQU+PWC4+WZholi/ZyKlRDd6W8tKMflfCR
KdG+2wlQ5k7ytX8nohJljdsg0y13Q7FCv1OxvyhtDicY0OCkQGHR2zHpLHkMSUx+
Yan0JJ6WFDMgauoLrH+tkKibhjhkuq4WpLEqRcsfzUFSoofmhpytYryKN0TQEONr
YbBOX77VX0vUspg6Tbq1ZWdGHnRHtK91zOJ5KT3Ms8WmVkPZZcHkFBEMf3KVI1nj
/WDmUkJpXwWgIpb3MskdOBR0u5kVCMn5HSI2rE1PeGAR1Jcoek2wTONIm7RmTuAT
3K49qno6HE0agBrpHufxojRGr6j7P5cl5YKTfaTTh4dJxYNRyRBowUVfBlPmXWvI
5ndLJpIBQYRIDQ5QyfW7RYyEqjBYeI8ni6/OuF2+Yarxlki459rRe4c+zI/S/My0
w6r1Gb0W85IH97MiHqc3SHJfgl3UIxtg92m0QDrcwOyhqOl43AWYxWdrQ+t+b0WF
FfDaDtstW5wtZZGFdHQQu3JmNgpH9BZfDx3OQ9WeOnjGP3o4++9dxZsDF3svDTfK
57MKvZROiHZbqi6tuC3aHYyBMhjYjp3Zbkl50+uOikvBjMW4IsUFAbBn+WX3kpNC
aUJVpQfQzSiT4H9+p1j79LWKfyWrw399UVkaSfaCRs3IM40i9aEIUyusVGs08IGV
9Bf16Ex2v03wkn26wns2ZgyCglhghMtJdRCjv8ScoBzhLGJDbp4uTjHJvbJidK1G
pPktnIRDilbDeHuwqVcK3kXKj+Ezfu74lNZc99eKQJ6S4ye/Rdjv35moLmdzmtwF
se/b+Jdb24dATzj2SZ4AQXKcZFiUTExt5mr36fzRSuDrcy73GWOaLO4Em8kgvdIt
b+PnUX4IdpEU7m731yjdzb3kp26wdyxaGcwPuyGOtbm6AxAgo7YuQJZ5Ab2kTTIR
0GFC+3cCpIa+RnbSO2WwQc/MLeoWxtD25H3gi15GM6L2tO5ot1b3TIDAWe9U3Nxk
e6i2Z9Iug5AhJH9irxZbeGKXrc23SIv8PDmMjSL8M2b7nTtA6qxgVBSzBeKKyaij
uxuAzL1ydo2tLkpZItO3X4LAHRqTsr0gMzwVi50y80AHHKDNOLbAuoltYT6jBUbZ
HZ+d6yzPguKwXarq7Hb88JPotnRD196BcwFAHGFwtmrQ1xROoTOK+xX+vMlaOIb5
/RdchIfs0v34KS3Wmbnkmf4qTbFc9nexqNs2fG2jrZNK4Mlb5DOAkgpa7KM+jc7y
BksyeC2DBCJpjvJGZmWqq/ek5YUVCKm9LnzsTA1/NTEcNG12BQjiyE4jkKfmoRw1
h2C5qwoai0b5JAadzjykjOjDDQSvWd21hfv1YjDwUDL91V+OIRyn3+SfrjZGCs6W
gm0YKupoa3v9jUV97XLRXp9dn+TMHJ1JAnkweE/rYiBiqgjrO8dbRCv/MsQEvEz2
lyCTd2hqPGc0iJVe+1E/RnnHIyUT6lZxPOfTKuKO5jDwP/6hZtKWup8hx58sId8d
vqomZgFYAonic2ZAA9vnLgrmG+753YlWUJjZ9YoZVL0q1lFNMQdmAOvZ2A/qTL8v
IjOfpWSLuhD1JgRxrkb9CFFrdWDjDj8EQXK4MlX9VCfjXSICsh891H4XhjcDy5yY
eOSiYsIravgkVQpG5S/ohaf+jKPDbKfQ3lpmRd8nayvG5Dw+zxsmKoDNwbAVwXjf
Gz2sOTZmnz/FUcc+S7cWQ9nX3c31hVgkpviWxBv0JKmwjpY7KaU1L+Ckm+NSY0kt
0VUe0ZBAYNsrENIldazabIASbQ0prpUUenKxl3Wo77UGOjpe2mMVAv7lS0n3/LaS
PR5V2Le0nq2CuehbCgybZIKBzmI8Rl/YBNInGUemdKUc1iO3ym6+MesuGukJSh8Z
P7qZq45A3ckviDH9evqVMJUs1f6Ke9FoTSF+m6sL9hrA93RbUEN2eKKkFzwz64EH
k0OwV7TbySAZuU/B+zL+TKNlS9TppiX3wZlmSW9233o1jv//S17Rg/KO7KZHXg1E
8HyeZmtxclYpMz27oj3DI8GgQMWG43A2ZpTZzM7FRSH5hrF2YKmSsHaQB8h8HlDU
WwEgftZcnPpkhBq+7g7JiZ/BftLWeml28Z8YlZ0Gm2TpUcr2U0U/y1TMgyVShGhV
MzHDi8fuyhC7hbWqk4NxeXxI/bd3lPQmdGIV/wyumD4exX7G+AUIanA+mjjoaJ6I
M3Fx4+LGqH3KjOK6YFPfuPGGMC9J2lfB9uvQTdzBOyrhLSkMAhvTDCtCYPhhUKc4
JBJ+uY/LXX3mbcd4h+wMpgxml/nRS9T7y54F/OQNZBudRGpisGuHvMK7RNfuUoPm
OYmOnQmNuZElGa0FKwsK6vWNOz3MGWtCwG4KhzuBqidfkbG36cSea8/EInQb6Zal
cAln84Ctwj+S60Fc5eY8x1WIlvl+7hNbIbtThcYPWRZuKRZ1BCIwqLGQ9jezTLrB
qtwhAe1kPhdZ/kZoSQcI+Z54iyqUZHD+fhmlcTFlPHB4eK9gNjPyBoT7NFRmM/pP
DUwk5Vmyc1uFxrqi3t0Ng2kQi6EQ/CZglxmCuCMc1VvWtpBqgllfhs+4il8vAcDA
oAtNuvJt6YpUXNoNQt+muoXxykiqh/TEOP+gf87kmUz3Zpq5h8E2rcUIDA50cCG2
tVj5Rnak8+GlhUDzVCTqU+0hjom75GvweItZDdRxgnBMAKc4wSzHytQHJjuySPCj
YC7J8tbgKWBhKJDNZi4AYfZFhjTMLb39iXNse3z5+UF3k5nmM57g0iof7NSb7f9g
y/Kc7WEFve+J82ZK8Jpb1NoxRY4OKmiILE5HVgQ8OBR/lVK/7qvS3Ac14DcPPGfz
SsaiePM4it2Lc3XG4GasI/GF8+izW42rhQXZX/6R7C6rqx3a5dsEAgX1kh43nx7J
qu4gULqNG33oFzD5U0P/Mb6MrXXmBlf00oU0njfSdv8Cz1gub8PNr2g1tTYLGJHw
ykIt5fhmfTP3I+xvRxeUSaxT98N7vUBJK1uODltNAgm1UIHp8p4IJ4Fyl/S/P2Eu
sV7DcjMlh2wIuZS1rF7Uc7MwlHllTx7fcaFc1k9fxcCRdd4ePhe0L/pkTLZbfn+p
B2aaFtxfE3AncgNhEHYWJvixH0M1Q0Thwh1mDQ6FMnnfqu3Uxt/MC7fx5C9oc/Wy
V3UP9JZoYyykvGdcnKpmm0AKz1frncfsl723dZuwAcRV11B3OJ7UaNS9Mdn3k9xd
yuXSHvZpURcN12aqwWUbGrSOYvFDWaZCDuP7ZYFwNFX41ZqtA2tBfl7rIRZVcegc
5eTAzpGTpv/xYxxi0SsLz4c1Xcb1BYV+w4T9BFpVR0hwoX8mRZ0lotuFpNFhlZRb
KUvLN/SNG2LN0oKxnCXjxEOzPmzJXcW0EvqfPM4dqLlQMCi7QdhX1EgbhA4JBX3W
/CCy2oyH3x8I7CGJX8XXg/dExHaPGDlXFpA4G+dk/pEGqXXHGhGfZpGgBuyWBIxm
2QDimy29Tdqd1oCGsDDGTGkyX7ICXCZC+bXKtKCzDRfFXHckMr425X7XPVGboNC+
pbocXRUJk6Ql28g+rJzBAyjxKNfvUW3dgpXtvfjDmJNw2HUiP2tEad29ceTDBP9X
bEhNcfcxKHoxP4+gr2+3dTxxe6Me9zQX/VtvqlcQcLAAYgnKwPLBJP2ewoytSiVi
OipTRVq9+/0XM2+76b7xrICJaPK4E+64iJzes0hYPXELxPGaR5JclUjJpnCbmBFZ
DVeN+AmcbJUQwktqS+6EuBxH//fmMvoR2whoRqmro3zPS1Krfi0qS4Th6r6m0Nl4
z4ik2TayLpBI088Xh4VXWM65FWwPEFfAoCAJ2fiQe7G3iQvHA2yMe4JJqEVFPLtL
zfQidN+BzX4kwPFytr3paeL0DbZUVeEYE8QehaGnN2OC6iAYJy+5Zh+mL5GGBnVK
JkIGVJOaYWlb9SpEqoSYSYDSpjs8hcYz77q+jFHajteqobe5rupJCbNjXWWT0/TC
IPPMO07yWksJ1zUdWfNymmB7ghtHnCW2y+qF+WfmFCSpz8LnxgIkf16/Di/nSZEX
Vu9ShHiSlkzPSfBwt1wYlIxUuGTaSKpeUsqTwZ4JK7Ip0n5F3hNfS1SBcD29Oubq
59EPklwUZ+v9PkFTNpHfYPGj8gVnzmwCL6DXjbCzGJZwd47xeS/Pzwt9N+CjR9Df
aD2dS0ihoaluFR+eJrS3PU9XtdjbkMrL8ni00FH0drpR9dpXdf3QJEOyitVmsr4I
p3iNQTwQnBLZYPffVwQQYRtyQgLFCd5H6NrIzLPc9eLK3F4FatQ0lsq24Y5xNYKY
z60nbAB5Za5Gz48Ig6Y70Fi4+qT8KJk6r8z4y3RRCyVUJrXvRiQcbMU4zoGP26ed
4Ee8VtRpbnA2GqAPW1tcEFxwJ+iMSo6hBeUxwsL8uUvTuCYYntsA79DibCUK6bRc
/Nvk1+ateZpR9agnP/SXW5QTkiNBaFspc70aOdI/PCJX/YDesb88B8NEvoLsBTkm
0MgCv//RkRIZ6YyjVaC7EXFbfsw1mDhZI2bsOAVXOJcGIZ7xPcUwZYSJExX6zevJ
LudzMh28843LvjWYHLnC07IWFc09rdGE7wmmzdoITNpjImAml+/jZopKQPO9oXRF
qIzwpuvWlEOAQqP+H7fXehRFBOaYVT5nnbCb/O3liI84Jsn+TlFQBH0vLNcaRiUC
qjNx6GTq6xGpcwYfMdBH6VG8uai8U+WEE5EEwPxVVAZGXAXA62GRhExsHRp4a7+Q
FXpSBg6CEpXMLc9YLtswZ/IiqZQ8DFLLHTEvVFmnaqrn9GZbKeyYSwmyAesSMfrF
T94ovSNWs7Sifugop/99TF8XJY19SVMcF5m2FK0//6/OVRTKXtDJNAz1qjQZCPpi
lsfx6rStDrH/gNlzsHmzObkcrPgQrclIKC6eUaYKTB8pC+O+6qoYCXvlZKQk655c
aKMUoDBgUmCFN8k5JwC7JxTD6wMo+DlShFuPS04+aCuuh7gTRg/YNFdrf7rS5XJB
evNV2ByeHR5twPjIE5vgJY+/YGAhNZdFiPSS3sPgYh7NxHlazBzdgJo2GrHgbVCu
dBNQCAESzSVMleiW5F16YS2gF4b3T7MJWecAPSq7p9WiGI0nvGq6HLNyflmuApX+
hMstAFV24lNS3jBplTR+M179Iu0SC+/wK6HMbRb5XEFYCiOdHkt0nvSHy7gLTbjb
VI/bq0FUc6dTvWGfP/MIS3/tXkYj+hBL2WD5wmJbvqUQArb/WmqF2uy1S1Bs7+WC
oJh1ENcasEJ+MVBAiTWHZEZ3iLrDJcU2+h796w4LwZcZOJiZf72q13Uk9qBtYrcO
05tTH6bMSIK2v4j45n6sMbwmek4ulyg+fIgWXG7S5t0v3JT3Dzq/jLXeC4EO6ULJ
JVWLop9CO57EF+XLvboJZiVGsDSBmTC2SWtHdiET2gAxD9VK8ieZ9yFDqCyCBSJ/
bOYNpIrWe9C/f6Ei57V5TWsF+qDB+/95Qoq8BlbReVKeWvfl6BHrZJDUFkhOb35R
fGeAgkjCqhYcFfvpqY7Zy/+i5+tJS91GsXkEqq2Dg4ng1PpsTuIJrNl/VoJAebAv
HOgHRVKHlAxnQJOxm5TzoP1wf7BfiY00Ghkq/4i1eppyICrshe+dM15IW7NhWskK
PbrEsC2/zx9gQAAqe4OS4kPhrn92p9bLrzUxXOW6G0Y/Z2yTYUWFa9EK306Z0VSW
II7fqYpxtAf+kVgY3NdNk1pHAr9zzBuaAgAYGICLvLUifIjSjaMrQucU+6rlG91X
fyStCHyrGDiLkxljL7JLCdlwMwXGi+mDgiy3Bh05LqK5VhfQTJXeZtLWw2t6yOZD
AK5Bf/nR5XqDaWvIweHJKop4yVl+ynLmulC6vhrvi9Mgu0JDHJmCRg3iiyBW+NuH
lXhANiR0z7wT2kyeYT2UzFrQyAgnRxn1K12l6ispRX1nCqHhKFO8vlLhu0Jr0l16
CpIgXDgf/EzApmy+rLBwxrjn5Tj0+REuWWaYFqQOWi5DUp+Gld8RZbTjMdj+VgGh
cLG8tubdfSDUqgPfdpRRvqqZyvJMq3UTbQAu0+jCgHK6tL2HkqdQcYWMP4d84wqz
uqFRFKixC0Cv8o2qenRZyhlP/flAp4vz/6c8AouKupj2cpv6pWletzk0z+3ZXCOG
bm8UeB9z5/ciyx9mAdyRhY3fPdVIh8G4E9qbNgVlMqPZQ6tasW3dJo1+dAq7b84Z
i2HaOrF/iRcE076EMM2YVl3nw6fN24fsEDxRUIXt6CQWUyX4PyyYBruNU2AVWEsU
zSJHljHJwUdxOYlEfdZj7mDEZg7BPDTBFVNC5SJGLL1EtYqlLmouifvQTHh7aA72
K+5+TS0HuyrduLh+h0owWPGZavHSeyftcVqF6tr7xfT2C8/wb3h69rXKgHTSYoME
FBmklKWxj86Q6KDW1bZxwW9AJV7HQ0hPZi18eOP3GvSX0/mREuVKIuGTR+RoMtVs
SgydfnnpCOtX//cfOn78N6duKgWDXq3yxGAqOSXaCK+9FPVvaR1gophf4gHbs/sq
mmVJdbibTBKJEpYFKxsSbMpoJ8ltcAg709etiOut37zEF1wo/MQn68S73CpQ4V5l
l/bmRMX9EBU39Yc49SiAD5r5bkdZAFiPeGqT+4P6BlR8jnWV0it5KN1efXWQH7h3
komd9dLwQ3Q4BaxRf6nWe2qN/vw7v080CiHcXFeVr4uDupnCz+PuJcf1uLvczStv
lSCd/yWWV7rjKzX5+IuCH19vozzOtMCk6ofx09wkhQjADn0ax2mVDNroWPx79L2X
GqSTXVDrG8daDEB7t0VtlCwIA+NB1DUhR6hH8I8LGIWZ5MndbtdTQGM3fk3E8Vco
5ISp9LlDbQMiFF4t429hfeoyyW09XyxO4M3Q52PahOjbLz8Y2+u46szwJrHhPRf9
Yw81ohtOqfAAX0YAljGgIOnZilBNICAQWnDS/xcMNesdgH8qUSXvYTdOhildFPlh
ZnUQz1zu85y6I+AE2qwW5DeETaqQQGsLdeB6nvBxH8f48W5Xgl04OoeIviZEW/WB
Zgru+iJaiUctDcWmn4jW1Y4sQg7wOlAS2w0ZQYgqgjJVEbBGrJYKa7P9fH/Cc9TZ
k/M0h7rNuTeaQq5D5gFa2i16Uz8dxh4upm6ELdMouQLhLTAQxgffFnbZ8A6553Sj
pE3sjBHVoZxV6sVHvBEpZKRAeHgFVKJR0xlc2EcEl3EiBUmvD7jXvEzpwZmkdb5W
sFAAAfiKIVO0A4+dcPS0XU6eTJqzqoTdgsirwchfxsStdcJ03C3skuw0QVkI9/4J
VcCm+Vv9DiS2HN9tFZFRbYhYDmwX5RJFapelJY515kLr6a3VsBoK0183Uesxjgll
6RMz1DO5ikskQLqhEBxbmZF2n6w9TyJVh2SZAFzW0kd7E0+bJ+aEjHDMN0ZzHU2Z
5i+cYuh8HlL42SOkKwQa/01H9HzB84jZyByOtfPP4B/2+jaLLN0/3U4Jr8Q53S7w
9jB8Gm+2vtr9d52D/L6o0YBi6cMNw4f9Xx7Ys10FDvMltm2UXxSghPHeSQN6oLOi
5hbxvhaghQwQYCmaSQU7FMu9fkL62gkXSn2x5zR1+isvASezoRLCVnqaZnFZgXA1
BIHCzdbgQSTZZY0MtKnlpnWdyhaxf8btRdzmqv0f/8NGI4sV6GKeuuuvuwj8O0Nv
muZEgXa9aOukogH4hcoG9oV1GmxaAAWpMdoN4P5TXSDE4A/CVma5KvKs9TlCWlXI
vQnYzfCt404o2g1Yy9lq4dEriYnh+W5rlOUENFa8J+oPIgafdtB/FP3vCrkXV0MT
rGscwjwdjPmNCJfDSQ4YP4W9H6vS3Jbw4i5N7GLP2I3DyqBvzlQjf9HztVPwRBFV
FaZLXPJAFiIbiFcfD/D4jGiJ87sGl3fBu/hxj9qDWwne08BnP1OZwgoKTKstFQFP
8U2pZvxfcaFFgeVbSLXXrRIMkHtw+gx5gWwQb2D/6WOuP1PRXb5dKf1IsIHQ4ibs
z5QLv98utWdHJbB+DYZ9C4efm4GGzzQFFwviVBezGbbIW97Gcxqqnspxwd9f1U6M
M1sgNE73D+X/KKv/PFqko9JZXD629NnfpgR4uvfsWRbIYznwZXMVA80VguNjPkSO
jmMU+lNXempAy1elCXK27A0X+s5PtGgANPqcdILRChWxEKfntEiTyN5VVYvuvuXL
Mp5vgEM6adXLmHJUFTWbwaCe1VlhFsBx4ohFJuz0ZMaLs0xdsAvd0YIBfDfodEWb
1O1olWqt5CgicF3G1TQNFjgGQFjazc63zEKbORxUXMzbsjruYkxlxHVr4D7paYc1
ay/1zVMvAJ3N2rF9VUBKdeS6hypwWJgOuMpnmnop1REux8PxvGzwC0RFfryDcwMh
FyJxdas2WF/ZmIekCDyNOMpV73LIJ3r+3VpCIm8PsZNlSx9OuhY4avkuolJlSp3C
7//Fp5OgmW6OmszTOhutLY43y+x6jPYTKBBlxJ7mFr2E4+2Mn9r/FE+qW28uyEnE
Yu/NjTh4vdsPJYqJ5yrvEJEO0P52tOisuY0AMnG/UHoE7i69cTSDjJQewhHHbrxj
DIKVeurtng3L8PwrMzvkib1wjnhFGYMEcCH0p/ZISPZF36Kdt8IbzJhAxbMVf3y5
hhQtNj+b7U1Monwi9DJxUVnHEM25wfhXuWq4zufkp+qaZZaVqB+Tf7IzKcyV5k2k
leTlM0Os+kVsg5G1cBLmrGqNwQ+ghxD6RMOy37efRdMOTsK39zikV3N0BJv9m+yZ
MIxuACP/GpXrJ3sLgU5Pb5dTdXLPXlFudMAkPnMTB9wKVVdXNqYs3MUvPUxZc0f4
jMXmRouyIirQS/z9oi/yRATpTH6Z5wA5J7SBTBwW8TakQouMwRO3F/7RMS7oDESm
dYeyeAc1uqy4d7gOAXGW4RicZt67YIJ/AdbMCbCcKKQT0Xqc37X4cy7ozxshFiWd
Jmt+wQ3O9CbOoWi/eIXKFbAN/z6neElXDrP3IkldlGnHq1GI8wFOPCi+AoKpmBI+
NfeJKMi8Cw9MCiFLjH9gc8cUtTrVJQsVqBbREdK5YqdE6RLzl/72kBfSC+b3qKwL
O9ahvUbl/8eOJ0qmyDTe9a1fS1GRIoqZej7OFaOK+bDk3/ySx2yamQ3uI5NZyXND
6SoIf0XTOXcfCWAU6Fpc7nW8EB68Q6rgk5y9YG+8iFrQBLxO3ik3Ft0t9QsvX1xV
QS7Nq1OKLTwOTwVaX0N9lAcHmRz7TJkoVkONG57cFH5TRd4xWFgJX+0h1V7qyAla
5w3AfbV4sWzTO6rTFQnFUSsD+hNUaUN+Z7Z1vs/xTCUc4GGR7DF1o4ib6H0TxjQ2
gGkVYLOWGcHHz2oEieY8EkpQYh6E5Qh5Iaznh1imkF2U8uCNIKjk/Nv1N/ZafFuK
x9NimIsTom3zzUgG7i28zz6T2JDF5JlDh7+HbQThmRdDe0kxPt8oYTqXrnJPQfHL
oW/eGiDP2ZPC7PhYU7aVSUsRofgII16QaXJxDiFg1yHiCxLeJDP+rs6m/YgOYJEX
ZGz8KZOnPNiK6uGKovsqWKJDaaj6IISI+Kb0YLDVhSIjrDQLJJlRUteWrTA97Kz2
UxKDOR7xmo9pPXzXPvaOwhMbcHJBx2kmqg42KdRvr9V89UgtOUoQNkW87yfNuBNe
Vo5MPOxehveViVkCzvBMJarh1R+Z4MbrGvlJLgGs7kjL3TAeqUdJO8eQXzN4XjF/
UlO/ZFYfextssfFZO6NdROMoG7uNxMVpUR0H+1VBPcvmEiSD3tAxsvI4hTm7cBdZ
jM8nRwdYnycXanZjDA7jRngIumQhpiqQdXCqhK8uwzdHuIMAn3AbeMEx41Eb8375
UOPThPxVLOSiLylmn57xENfgj7awdlI4BuekdumxDmeoTh+7ioBWCmiQeDmVVXLd
MemqtYMhMf0CAq/4KR8VWjODQs9cD5k29VmwI7bLtraTN0MsNX2VwbrVGx6l0s9s
pdgDDlx7dISVra6yP/g9ha8skMoSXs8Yv1s8rFgPEXRTtasE/R0/7jNQBdwTn3Jc
OjKHQrc3TZL9uGlxlCikZITQ8Cf7GWz/0RrZRfPMhQ+W8s3ZU+7pkICdIDZU9wUV
h+KIYQy87DzsbzuvC2npEgXzEi7a3dz4ZDSV7JTXmcnBoseq2jgte65Kw9tB23oR
nR6BaAeo+cAGvzWP6GTfNsbg3LZKTJm39JwLoU4yodr1Y3lZqyW2HvCt8kBA5+Qx
2tmRrOSaOleUCOHGSWGold2GphUymj8RWZm2w8P8r4Y13ZkqmUTnoMRPwgeE09Ru
d8/xSkK8TxYcywyZXWC/uLecwKK8j4syrWpEaBKp+c5PyKV3JjaDhNJSIXp7VfnL
cXsa2KaGyKjgqbrTCZCfUVq6R9J8T24hwRXw0m3fB3PaZPxtUocDNtHwDlxzVYPU
UQ75MKK0T0fpmgb2Hio9UQ+HlfgI+8Z8PAz3UoGLyb8xMqiHnlqZ7dupKAfO+C/A
AcJ4bAqfdrtQRJs80I68TDsGJXi0n9wnmahkeBNBwfu/CTX5C4XXlmFSJ2By0orH
ldHcH5cn5RmEERN3PuN7tq7JynZ+Q2w1XBNTBJFayO+RjhPgY458Ovzvon6UVA/B
2OzZENoc5ci0m2yVCxPT/rcgSDypqrjEoK9fIFsaCngfPMwVDlE2ZmtZ8halfOnx
jIRewCton9ke6pjCQDjr1lhDf82hzPckHYsjWQW7KbZVjNwaHil37L8qvuSOa4TR
5TzMkJUOtYMk2uyrvl8xUH/rYQCWxWNcCj88DN1u25uRTuGuhZwP+0hJYkomiAzu
dJZFReGiprEtGI/cuWG2KZWVP8MBpG9zIPBYlh+K5jkjr0DLFgcBIMbNDGqq1Sc5
FZL4jXyPI+sE/9/T5hEu6Htn44OVQPL1Hf1ysKTtgBDN/PeuQjsF5LG4IKzfNH4R
ZWzKRQeDT3qeRFc3KW6iwoV5HyczyKE0GXHDyKINwHoJraRpkkYfQeG1qgJHtQFC
UyYumeZJzNkcmWAvgXufnWjsvBhVqtfoMCf6Pn/zzqu4/LL6ci/m35AXQySGJ7h0
/nC+n2qg469VaIv1a/g06H4sMu+XAUYlzqVQTExjflga2jKfC5ClnCqlrevwIVKu
1K8M2AkZ78LZxCYqhbif2EOm+6slGjNKvmcV96RRQnW1fWp5clyX2KlyxT6ygD1y
R41hhaxu3Ip6U1zUXdt0h0JLkK3MMDeeRw46ubTbXXlzcHutnGYwUQAROOAyNCET
BQXi+7oKQlgch/mrtxnS15U/ZYF1U1JPqQN7NkpvPW2GeZUKz8u6q4ZXiO8n0qc/
GoIb3z9nQ5kqKbvwOcx1v+2oHZezaId725vtobmceJmcUbOve+RdMkeXa3f6RU6H
3lupSNh92g68ersDIK5Zsltz0ahLx6byMza4HJkgUOWMAnT9hKAYi0GqVH/TyatB
ufH4UtZe/KQH7skMBLlhmLTtYdgy8Vka5jMe+u83GMB70XbSKdCb6iyuKQRlnk8K
10C+244MDm+7bgecsJBPGOiMpheIhl3kRNWVvRgdIo83csYuRurxEE6gva54wYwf
16Go4Svdy1W7yHJypSn7FQKxuMiHF5o9ppisDRPzY/JNtfFmHjuyEirTiJUoAURn
vajE0JdBucx0P5uGVNaP/gv+d+0GkFFJN15XzqieXsTX5ldoamNzrXYWmRUSL761
unu7QEtZeld8gDIWJ2d00vWNqkSu7NdRQwJfYWLqQyiwDhcGQ1OtS1EEZpP4ibTz
Fag4+7fjBsfR3scdBQ2hxnV0yBxMGnpXxpLY0T48JcY6AmScsyrKmtvZiK8gS5mH
RCUYd8P/0aBAXIGB2SfoiNgS22/HQ0Np2oZYgBBO1HOujcA3J3bB7qVKavfY7W4I
k9SUdVJIaCbJobF0eN6qzjg3GL0qeBXhQUKqFUy88d4rrRdVRXRXOzzuQGGwayNx
HYXGb5KFtDsWxB4/Dza2UUA8JnqaF+m5TP3Tbx0r0BF2j7S9guPl6MG369i9VV/z
mAYyI9fyhjlwR1lxGnopMUwBLCddkDke/ueTQTxuXJ3yhpPYQToofOdoxxltEQUz
HJVBDQ90EWqbcrgy6CtHtkRrz1Wr4xcVb3biQK1V7QC6SIw1MCxzXm+fNQLeKF2K
pxEiF6+tC7CBjcUCKugiNjTLpPsSM+pE3xO/i+MRViY7tgyQjMs5lBIVlUzYdL3P
M1YUTUwwpxXYhKNZSyY93oh93e+2zXlW1ppxpu10DDkLb1jP3XWZoUK7+jlKSRjR
SMacEMumMwKguD+x7by3tHocgOP9s8tx7tMIo+FIbnVbc2fw2ctnI9wjlrWle9tH
iA3XE6Azbh/+8KBnlpWuOOkb0T96UkHLY9TFEmmHm5FxsoWeDiPZAi1flBQjRkxe
nDj1nwgspzeJZ+PntUK6K4mIc1D5JCjI9Eyi3CepauW05so6Td3F9dUIxR1OmAsm
aMBNZTEyk0Lp0K2gjFij63J5vOSHDAHrUomFHvfny5XfWQWRN7PGpbNwA91gWtzl
bpx8nzRt89NcVc9d4u93Mc6A61YI2SOvVSwcm9iiLxuqNVpKuo7YfaWxngmTEztP
RWDkSLPQBrZZmwPVP12Yp7smeavlOIGUBDoAsnne4w2roGUU90eehvOeTQLw/x0S
YoLrZJCoeOy2M5pADe8MQN7/XSUzulEkn3dNUQ6Je8Lz9cTcs3EY1Xzv84NZYj2N
CE43TMK6f7YUkVZ9qP2BaEbmh33ofaU7PhniDCnqJ2UvrIMuePqJDwdrhdWWshrN
yGXsyU2ntwFBoFCHBOkxtTMYwxssia8ZhXZIhRXLEW4IxCqI9KAc/hT7kUJwW8Pu
+iFWdRMxkXsK3+Bvb5ZIjF38wTbvX9dH/7mfQfdQgJBcWs5ubp71z9qVZJ2DobEm
Kfim3BrqCtF6DqGC1n9QXaHk7vle0Q8ABZkSG5/DrVQmpGqkOubIgu9bRh655GmI
kXvbOjzI8CSKyFUYTcqswSo+nNv2y2a6oq8wpUaAQHOeEcLYB8GuI7JcnW9cF3F8
qsZ6Z5qWHg+rw8YdZ+iAsSVKPNBmvsc45IhBQGgb4o37rcbJwud9SOT9qAs0h2kK
KES/OX7L96/lHJ+y8Y0EgGpWIHgvPmc8WTxqcERalq65r1wl6x1Pbwi1PYPT7CB7
Lm7UNucMHAVwaK7VmOlkaciqvBo3bHA/W3H3XNIvaa/m0GvYt4XqFkGQ6Bcs0B52
+GlZi9Acd+qhKSqOHsj4tFKCCxuv+OXZgCKYoaeg9fCfnQ4LYIYTqIJDwkQ7o2uG
Rna6Mh8iw3/Zh+trOcO+v7RgwW5+hHeGkvGs3rRCXe/cFIPtvlumJf7YXV/7mxY9
cweL2AH6MIaZUy1bDpG6gLEbFiJ1R7LkwvKWgrpxjgOfRrmW1CKRj1rbaooKLNl0
RzHjjbn+anJ/ewIvhbewuSWwcFf//zEqXUJ9Fq4+KjIGBEwct6odIYYaoD+0G61G
tm+LSHW/xcmlqyjhwzUYv+uZlp5PnHbemjpU9NvvbQ6Oh0DP9pkUUqn9K7FuiKEw
VZawiEyBqH0JPHkTV3LL2RH9pWC8pfbaI0RbwEa26zeYIJbY8f+XiDZ9bZSUU/SQ
kkiYS1Xk7dKCxiw38vhaKKo9f8Znuc1NtF57Pvny9oSKNh6vIXbFdCB13BnpgCzi
WjmmyjFNXFqgT7YN6NY5x02VX6N0OoIsAK0yjlap7SohNqUXCfdsC2yTlNTV++4i
7uHegzrcADMSIZXnsxVgHQxn8vTJ3YDBySNHWntSF/Zr2Cz9NVY68iK4ttg12jL9
M49u4ovPbCaOziK8rNrpqHW3VcpqHltE9pYTxCPS1T8tZ3jYYpm65tmjBto2kV/V
qiKpJUeK/+C1PMSo74US3EQqQPFs1h4vKiTPyrYajR1vtkuLB1pvhhLwLam10ZIf
kJjrIBgOMjeMdb2wJ9K3MqLHtisd4fDuG+OBNOx/IBE1clPwXNilEZwzwW8jFZkZ
xW0e3Fpm2cyseJ+r1hkCh2ZGdHn3M1Odd/ce3B1lf+wngeM/cQwkKKyky9Pf30/x
+fiJI4qu3R59Ju2KiCXryl8+D2NWWN7EuXCqCg5p15odny/fiXm8pxfDLv4QQt9B
pAQruZBs3YbLTobD3EMChR0KQB0cVDSfcVWdVfEbB+LxE9C5ukD8pb0IIaBW/9UP
NI6eGL5kOomkblVsyOYO+YtEz04Q/4v8a4ktfuLNHiNW2uP/zOfJgShCRJshALTn
GneG/pwMa8aRhawS3FdvW+mVWixsfuqL9A699Od/NrOnmjhV5Rdu5+KYQ17xhl5l
Pnwa7wbmLNXLH4Zprp5Bpi1YvEe7T71URQXhQgcXrODn77cCRrDyUIneXwFFhqoP
PyGgJs7Vn3s+NW46Htun1jLt+GZSb2LDtmZNOjtzYKqFPKzL94wNoBb7MnE96AEF
gTcUiUuAlzMoVgnk1SNbxmC24I8MKPHDFiCfB5vBZj1yrnRNcd+IMYX0t881CfDY
ZvXBUpUSiUDZ9E/eEVzPj7Ujixzrqk+MUGZb+jGNFROlo5KNQK+i6jg0VdD7ZS7q
F5TrRPbfgWeUQRn92JppKT9Xc1980O6w9oEk0QNB/xaiedRBlRYNVihRYSfR7zms
vFV3wHP554J/MtLBI/FgopeP0awTADsYFw2d7nx4stozGkfHaRP7U6M41LC9itXz
b1LSY0mq5G3gjo3XiJ3MSBjp4zPZte1/q1pe5T/VmMc1gKZq9G2bHrvOwb7s2M/q
ayQ0IcTJN+GsYmf5Dm+eTzU0F3s0YJxySZLi+CKG30m6IccgHODoyjAgK0mWGfzq
85NhzR1K7lXCD21btZm+McS70kcG1JxThKkiKh+qBwXOfyRQwPL1x0pj2VXmbpL7
f4Rp/e/EUXRN8A25pCSuncDbKJyeVJW0txO4UOvClxAdEc+Aj8JHDObC0y0RLcNe
lS2VKlti/2UJyK87rvVpaL/9rUM1vSwt3bNBaGOGXE8ukUVDmv1Xy4I1rHc19lbt
jmQjab01JODgH2sGGiZDsjBhLB+tMm2oTwFSFruyqr7c6fV5pP0oXVg0KRK5sTnx
AmbOLYDFX7CrDr+FC49qxnGbhyy7PoISdKT+aLcenxhooGFtdD2PUCT7NyOYsfDS
K3f+9nEMdFimYGl1G1HhJD3JMS4QwuwoWGhn5YZyll/qv45Ssw+BQRnVxPVTm/3k
gDJVLbknMlSrznufVY28R8O3oO2QxFKWRLEy8RmJxQSYP5B+3J2uevw3TfMYfmby
hZO1K/mHUAW0InY9TAgnVh7mFQjtG7ZlL/fpwioX8d42c4UEwsh3vZRtUvhidV5t
Udhe1qtNo1gqv/mFQDugspiqsEhKwEVbspkDsZ6B/sy3MtybCmUGnohyJX+1+jSk
Y7H6Rgpevo31KAe5HiBvbabP1o8igMyZYMp5oriED/AV6/gZIV/sVkCM5b8S84Cf
mvZLjaeTcPnPJfL8YUUDhaSdpyXVKotdtLgRsXlTCZ3lsj/jlFB7QbnYyMHJJoeU
zTNGN0lnkFJqgeuya5PfFd5sx9Ek+yAJBSAjd5D6kR2WnYjNmh/FKE0yOxhAF9eo
tHgo9kQZNbqBu0OpHDni150UnrSOACVKomavrHm27/wlw6ws0neKYm/AG1O8bcuy
m3tNDBOGPOUrfrw1QLPBlSpB1h1+ejMasDjrJrPxggRcwxvLCk44pr/Sv+pfw2OB
sHd9rWF1Wo0gac/1NpeB+MbImQpzT7zBQxxxj8+AuThOVX8f1ip97k7oxCIqhWst
mAcLIbgtPA+atneusux20XjN+ycYMyT95FV91nrzj/UA8sbtjWLqf15/KPwsYy/E
yuXHwX7aJ2uT7fGAN37rCVWoAAcihfXPn6RlqpVoE0f/PzOgoijmq0VKnoJdVMPD
HHMmZEi4UBpa/Ore5WYrna8u7esvNx7W40xvkxYRZRQFl/BclfSoxGlfegO0WDez
bagMFIOIOAGFi3W4IKo0GMO8jC+6hKaSfsKtvknllMhuSzBVHf//5qJQ3o6BZ68e
hCEZVcJ4bZQmjN9xgPQRc5wX2oi+P2GNN5hEO66KfdCpTTSCQLV45azRXCFqVdVC
w0keDwAmO5xrx29Bo5mVKALlIZKOGMzskrZBlHfE+rpx8Yty0BzMJxirrM1vIfEC
4NZBW1SCc15JhGwZI1l7iim1aXHWD8DOZ8yVA9v0InAKJ+B7DNoCtnX8kWMJh3at
V/Za5l/8WjbNnqCMQyM3Rj2BBF9Qqec0jnWCu5WpIOm+/gDxpeF87E773DZupGRf
W+tIa9OGMsFbRKBw3XeSswBg+so1XucfBVzYuepgZJHhCqh6svm/ns4EqIWuh7O7
ahMvqORIpojUMQoxMJNacNtwByI5gS2wySbFWzgy2RQgSsxm3/faldLOUSb0bUDt
jx1myyv0iCfJbMC6KoCDQsY2tJscGD7IhOqXi8orf3cdqo82RsH5NNuHQHid0m6k
9cJ4gKHvGG+tPkELqtpTe5YPwCUqq6nZXw0uz0QQGWwVhXL/XsNDf9WjCWVU6fv+
csfwRj4ZMRVSTMSxtnmyfI8918nZAsBVcJnGeouZrsxvygkvVJUU1ovU4ZI/I5wq
4FCsqQgq+DQukvlVhRC5MAuJdgW0qJ0EAno/jJO3wtWuqtujTnQc2aBOol6QsuJq
xIndkn2CMbY4etptYMTcXlii1DqkaHbZh3R3de1C0GyYv5su8JwbcQTP0O1z71b9
oR/NbdzsP2tQfqk4Sfem7wNbCxLLCiaIowBdgZcBje6XJ/3CCf4btQUAokMeHNQV
gWfgACpCAZWfBqs/ktujbsWjx7esBsbrhSD+P3GyKWXOKmw2qdOVC/Ml2TL/+yor
gbWlEBrsByQwWK70mbArmdSRR8HJ4JfqU6bH0GJP/85HkwDdjnkxShxJCAk8083s
JJJbJgt/XIGBaclzP1WAy4hSnvX1RiL0Iu0laVZElKpgGYrlkMcpGlGHhiFm+91n
st5O87jXXPgeJ1khUAUhJ3UlvzSjMb1iXpzA8AMRd5tehYE63iBI5bkrhbvKkwQt
ujm5fcEdGRwL1GTUhaiB+ol6/A0n1zoY670CdHlq/mErmLWhd465Ji+as38CcypS
8L4dSHEuYx/ehepbYIM2UAWD4j7jWguSXE2UvReFI3tG7o/iXR4IK/+4yb5srspb
M+cICyBVgj5HNI3HYa4jpLWnSTBLUImixS64DBHz0VpQ/ZYD4YotGb6eSZXw2aJG
kPCF/IJ5xTy//D1wEzdD6FdTrw91oCUKlN/k9f+tGKOCOezfMakK5gjJpeVt/81j
7wrkoAhlkkeGS2ivAiRtH31hCpyXAD+oXJWmA3/v+7sog5RxeaQciTGYMlWJRyqk
HX1ZtgLzJrU3v7bRSRjrAzWMGNkSN7gvFMiXHSQ5wgEeRwZSJlZtca3Tsgs8BT2h
NJbWQ7OYgaCx9fWnclu3HPvMCSQWR9Cjg2v0DA+n/P0Jtv3UsCiHup8TRdK6xn9n
PWXVqnRSoU4q7ZnnlXzZ/5lexYApX5uiXjmKUoSy0Xbrb8m0rVPMS8io1Z4R6dDU
LiJdFy+rPEQMfP7NRf5bP/3BGoRhDN7C2ImquPLfojc9ZIY75uz/yBsYPN/LgnxB
7LkSRo6uWPs9UzrYHxOUoe7OcKMoSdTAJGzGTmW1gjRFsH1AgIANUie7GmLMRwdi
TJsh7nussxtagOOsxMnit+BpmLa13VsE38izLT091nxEXlq6MRtIphvX3qxSct78
eAnX4zJw5YscoZrp0+QXAOJ+QzyhJAcAxMZMybgS/8HkRNCm2fSOlAPI9aapi5ui
eX2MTNJ4BZ6FIB0dBbd3cJnY5Kx3jz/RvnawWbq8jD5IKse1BM2DjYMOPXRscoYC
fypGH1AwHkgYzK9vO7WuWH9Q43oLGNq92oAxL5u9+Srw4Dk8gDiWO3MSpBdew2yf
bazzbSW315OnhBaafbSkmZ7I/mQXUBtUjBSCrutR54BdNskWrd6l+OmWDBblCZFj
1mOdcSVSkNfs58NtYRZHKi4nkwKPPiT2OgecrOZTGAIiSLW1LWbrRvMQ9wOGZsGc
upaZia3SLKKDqYzXEIeAE9vyaisdP8zLof2JPWippO1hXckAWl5FMPq3t5KTvFbJ
3Cmf/zrOq49C1FveE1f61iCVUcAebf7op5vCspa0scqoDjPR/Sv4TyImrfp+nMfy
VB3EUcZVgi4TyZV3K31JLCoOHe3uGYob3vmGlaj3AcW9BX33UOUvVeHJOaJROBqa
lpR7E23bDrOfumosfrSr1cTvgu4Qob+Nf6Bgz5XKrT4RECjVXgcgTQ5ADL3lVzkT
pdhVs0TOe+LbNrrWixl1bI989DhGQmjN5tovSXDaS4hbTgSknsPSBtoY407VVYn9
V7g9oYDvc3BPCM5srDdAmzeJYVKG0R3rGAHyVDkmszH0qncMRWEAybQq54NPB0sz
xSJsM9OQ7c5QjT4RAiCtE5L2/2VrxZFXG4yW5m+hQuPQmPn8ulmrKZd2yat2rAxy
xNMcbceGqH65FVsaETaqFekPVTNJ12XQ/cHzsu2Ln8jDFnkbbEhkcT0HHukpiecV
/QPmtoDI2bv+O2EIaXMBgjDBADaGyFqlc5cl6pu6VZUgOymH+fbObCicmd/IKUsA
TmB/w3Ci7v5GCgVICd6Sps4+MvslvR5hC+w1Vi11FPlXJ6m82HuQzMFJLuczH+cO
f0q848UjsxCbuhue7SL9qURcfpcELNUWxZbCzSFCopHW0d9PqEapKS6yM0JTb+7g
AJHjq/L66GJqASZCzNZVHCGew+uPGabeqtJe91xOIzYXGUJI3u5yUYJTHaLA8ApA
nPFEKej4b1+4DOSF6jIGFJ7CPG3xGMeDRQsXgdJPcezJ0mpXoUdVYtzQFB48dMF4
F2CBlCsMb4e1QUuvVBtFdl4kTY7YCop2twsgM8ycu13l5HrUno7Xs1VpAI/YWggI
4uL7JvSXRZ37nUtiqQH10Fzm77EQXsQhTCUSYhzQhXoyCwEEATpwQ7JgAAhZ8Lbr
x/untOf5rByUEwd5sV1QXumYmxz9BaQ7gPyCLElJM4wQIRAvqulrmyyEnv9bimR6
2j+hjFsHRGF++DH0hhngWA==
`protect END_PROTECTED
