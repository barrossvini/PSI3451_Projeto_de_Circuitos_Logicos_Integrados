`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9DbOeFSaqRXbDCDpkNYkE9IbwHdiEEIBk8veDfRC7SueRrwoEAJVtOUz62ktx4Hh
IsKuWPnGB7Pax3ZwnW/91AMswubXEhayLMYNK4oTRbRM2c0F2hPaTuLwkS8ZIQd2
jgnGO4+XGKfnrL0VTve4qYeYCBmaxtCbcFApVP+awuw/jVP4LNF3HIYLjh+n86Cu
Eum5XvFeYEghnwKfW8aV8i6DsUINzb5QOYoKegAsI+QMoWmcU8ABntCFojWFWXTG
wauomXBIHMf/livgKwRjK9PauUrZ8JS83iCBKNpmVDixJC/Fq+Mf6idBjtlQgZKM
Pfwh7ukce0YK7UOrBVQ8NgzBaZobLNMAmEk130R3+vRucXXY0prBF6H2Zp+tzYez
J4sW3bJHEpSLsyWg+W3k6muwlpga3mT1DU6K1lTMghAboAnKx6NFbD+E+0SgCrvd
4S4HhBb+Q0AFnkSTXCrRFrvC+yL1vY6Iv9yGC9DO6DA7PdlAGEMlpknpLZ1jc+7k
IdSPyglCKiueexm9Pxtr//N0fpJb1aWoWDxIX2vzsem9MiSsd/ksPcTrwdDumMfB
4EHjUQnq4MqFZ04Un9oj2P0gpWcsbVAHGqmbqCWy9spX2JQaxFxB0rsJD9jlw3fI
8nMYlWeaAi3SOR0kW2RYHHSW4W9W21THRAPm3aRLoCuR2zkgWPMlldqjNDI6I7OQ
JX3W9hI/+eCqdDBT++3WpdJx1i7mogLXnvPkxwYYVSCUdvVAiqMZgd5Ch586JX6R
OGiNLJ2QqqxZHlsyy+aZ1cF1IPS1nYKZuOlohsqbubtZs0GP1JBBqQeZcG/7Xm8L
D7Re9xRsNVG0pHNWODyIQhSzN2Lmznm1TxBQBajvYg9qkCMpo8fGKZMDrPS+AUtl
1R9ThJVdDkX3Zi1ev6umef/ihJiIOEks3MFU3yx+B7REgkXMLOKz/i7nOBrZUrna
intt8B4DKBkZ1yNIQqqLhxZrh97/vCIo3jagPBTgu9360gpoIPvYc1BR99QwcaMe
TeRY7x28ingM02SfPiGYsLjjHpQPYNoeAbC9QyaXXStrW6cS5X62JLrdDOUDl1Ik
lB4XppOB0E+bzPByl32oZUAGAf0Xld61AAg/LqzUDXbdOUN0JOAEX3IhspWlXAxA
on7hUGFsX0A2yM6idOniD7frD5iLKBepmI28gfYWgug9gL+T6zID7/YjCl3Bftmw
xQOcmIZk4PA8tgGl+GCbpuhGdLqEplzieSkvcqB4JuDiDSN5OjA1uio8/yUtmtX7
h0fKbwhwWBCXmRCAHtAsWsTQiRD/gcksl0IV7ly3FmD8r8Vq/NcBMIFYYxWWJYbS
G1h3SHuocct+60Qkez2yZ+g9rBelZtZsR3Jlyxbfs9xf9igX/XIu42t+i9ED4KQ9
3rXmcpzqZbKkV2ef0RTrIY4Lp8PAa9KyRiv3tzVz/tVwjcv914NR5uMwVyYVvHkx
SeurGo5CxRmwkJ9X7b0aKakGs2LQ/f+Aik/MgqmNGxn3HH7MJKQ4HoZf7swGNoN+
oYdeC+Kfz92Nlq7pVlXbcBj9kc7ySPpWfrYNPGggN7s2URgNeJWai99X/bsn2npv
9OfQ6a5xkw/YfJQWq1SLMiAvnWb3ZeRN+BHjOY9/1YO1Kga3Du7o9HJ2TDEWiIaJ
mGWZ9JMRMxTc7mnuaXLr6iLhHDT1raGR5/dmQVA5gb/7knxyWQ5GevIbikC+i0i6
3P3YPs+5ZP7zLyrXxXaV6s9TViI13Qhvo9X6nzIUAfLMx//fBPcwk3um4GlM0pi3
5c58g4n1t310bifw7s5w3LVWEsurB3cCPZ6imKB80A33bNvJjgZoKPlovkLmoAas
6anSjYJLn+tuInZQ/wO96ZIFGOG6TavzmxKtHQ+LuGLHqhO4oHmgm26h46pqqkrU
qEoR5c+JxTcQjYUgJCBFjBQcJRJVlZiy46IW9k0kKxxTxHeD8N4UzqBTJ4a28Pj7
FHFZBr5j1T9VkvY27PQR8eLaHc0yaEQxs+DNUT3EQsYhS6Soj2JJ80mOUmIuRlg5
CzQY3iv+n9o7Zo9LaH9vRzrbxZ87avirRsVw42pHXp8VYNXDzXUDVs9XpZVUTsoC
qII1QO1GlvsqFEmvNUJhMZ8shkGiPtEY+fOetHYomTlPm6boHUBs2dj14V1m8i1J
90iBTFllXTWyVNYJIbj9si5nUp+wS4mx88qqZ6UVDggqGNnexNH3W0JIASyvTrxd
k+6EZJiN3jW1BpA6Z2yy9nzRzKnVoWUt12g/QQ/oJ8xkMxRiYvj3tMSB34YmnCam
JkyRuq8Z+OB6lL/LGs9YEAnLymBKbGVhswg/4G7WVSFejKnk/axuW3eGHLryl1KY
DK5AeTu5m3c4qFbZiHc8kauA+DVVB0PI7AF7vJNMfbOhXEzDJ10TUfc9K33/j3Ch
3XyvDdfLlrHeSo6J47SVoLWiJRI9MP+cSY/dNKKImtgr8uwaQTMVFHuT5s6MP9Y9
ko0Er5mZmzHxLEus3EbmQNqqSJc0ZChusVaLYIUCo10q5nJRU1EAVHm7yywp0eX/
9p5CfEQxxTcunUgDggIvZqAQ1uGNQWAjfynJ4ne2CaAspTbhClS8AnQwx2cP/0Th
j+CdICFVM4my6T8RXAA3hpV3Wj8iNKD3VUdHlHdKZac4nIP4JKK3ADr1caBn7cim
F5Tmph6QbmxUbgU2jPjVkMWZ8FS6SknNArXkostIYLoalbdDyppU0P9vtHAZsyAV
tUrR93BmUhdUHbU0I0/uNlLBW1Mo/cgTFoNh7n/P+EcsSooA/DxAHQp8fKglSDXC
VQZQwnx2jK+hABYhiYnaoO2QMAoA7Afr5jTb1SaK2CiCPJBMUCMkDHhA16rWEl8V
jPpXxOFa6Lnn60H3i2y7hO+ADalYCBk45lExPtVdsBpcCMfg7BzOIEN9CWQZw2c6
R+ytII0oUQI6hwkgNpYyRCioP4eCghNAm8KLT5plxtihen6/OX0xgIPicOzQptUi
/YYEBRc+T887FG9nFosmuvwtnobumytyYdLEgAc/VJ3WBNN4J3dD///U0IvJhc+c
9uteNLHrVMqheZgDgrKdj6CHIv+zz0IcWhL1U6Or3rv4CKC0htxZTMx99bsdO/Cz
vSL89v57EZ1kBpa4hi/m5HR6yWD5evJTThb3jOwjLFf7LBmtbrrL/MZp9QllS4w/
C3Pywu6CorfvOotvQJfdLZWN/O9J1Nw5KNl6cDcv/N0OgsVSe2EJ7PJUSBTwSnCj
IMyAoCmVI4v2TKr9or5rqZEk6VjsZmiregFMB0PgmhSR683ODjFmX6PvdAcaSB97
BOHkIRFb2/JRb0D7BIshMqWV2fzcUBd299Sbu0uzmCI67coa5wIs4GNT2BVXftGJ
DrG8dF/SlEGDnsVIKAxQgIy/DxGW5kTiZq/nZM26jtB7tPBAO/8eJ37qzMUKpovZ
WyI4VcN0dspumjfZOGorgyROrmGFhtaVSJnZEjxQ5qnRzHHg+Mwhs7y0E3P436Ee
ACbeApIaA8DIFXYTQ+1h1AlOtT09nWSFZT/TiluYQZRy/kd4SZdrTQEbzb4PpTV6
y18/c4xwt1EgOAo+Vy8XA/vBqmCMWd2TCo9q7UCaacQLPO1ek5lTeGgxHrVdYS+v
`protect END_PROTECTED
