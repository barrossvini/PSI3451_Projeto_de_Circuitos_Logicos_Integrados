`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rcuz49ToQU0m8XAuEPp4XGE8wG5RF4Jg5Qkm1jrrDL8gqPEp3mTU/c/jIU6op1dS
20vlV0XVbcr3EUF7uYsJdLKYI64/UTSbGfOlkRnel43Yba3uSVcwl94w7mnzW3ea
5zwJLqNlzK+432tVd4nn14LLYcLjFW6ZgESjSQkHSNpNGmTCIrpnsIPArQxSki7k
G2OojQ4IWzh8rwoADdXBpHyzp6QzgYuRSfQ6t8sapOdZhlpfC0AXtr8niMMU/2An
Jdyo43AuuOEtT7Tm+5DL7uQhkQYVWODjhVTr8p6yXNU98RKk4dnvdD7x3guxSHRA
uolutTzuDtc7YFmHPdQbc4TK2qK4D1078KulX0FchfEKwO8KRnWJHgTqxIiVDu1G
qkoqma7oRzQsHrt3ylMksSndC2cM2/Kk05CmvF0zpytpykeG0NcADA/3YoMLiYIi
D2sh/u4iMbPiQO9Erm4FmvUgKOsY6FaFaJOla8m7adAXVGtlVUafnMEME9eSK1n1
A6taWF24NWwEVJUiIafO6ORArqsT31M+xb+rsCZFvpLEsaOFbr/zzARAPToER8gN
3aP1/f9hB1a8Dd+ePJ1awWge/sZZnLpI+qW/CTkpuThq5mw0QWONmglzjzJeJabQ
Tv94kcWBSuCbdDFRUnYyFj9Xc2wgW08w1FjCRCE56rg4tozqEJPCFoIrJKpHUYXg
BVD7PX1VVqQYl79dp7DiApcNTtKdK6G6glAob4mz/DFB1WFmfj1e0xjoh9E8kjNl
WitxtQa/Zn9Nynv7b+G6nE8KtqPAaZCFjoJHQHj7lzeTiK2A4eB6it0MP/lEfYf+
OwbGNTQZ2IxGiA73aeSUQBDpCTdMjeSjc007R8LPLLTtv3+OXd19SexmDQynIamq
Ml0ZQJvGCWdJ1G5qJG6ZSHCHzP6baYOogfWVkSaxJEF/yKfdqNrnHaFPSvme/GM7
35td7z9A413w6xzQY9vfz/7oYtoMwRMjTcVgGZ9cYh3nk5gNQkn33q+xT6ds0gIA
O49+GzB1UFR/beWXDEi+50DEP5sTf6v3ptqXZG49rMteATEu0knr9RbtithMSMRm
uQ2n3hLFyKqaFyGC4J79pqdJxZxoeW6L1QeFCzSi7iqG+2/RAdSb9OFnwHrCxxJB
+1CC8pg2JeKmfJj4DnYAIaQDuhy2fqEMhljBXfjP1CCDaT1Cgr5Ikg5Q4zSd0qSb
eFTi1aX1FVuF05Nb8uFnpZpGoUV3STKrebhKeprPFn8znfH0rlz2ofcw24a/HENg
tKPoE75lxF6/7ZWwqEBu8RGwqvaIDmpfSJJj6vFHsvVJ5/+ku9zdUqLqzLAQ4h8N
WUM4xJ8dZ27OGpnp15T+4+/JSJQHbNgYuLEhwV7wdd7TRFCPSPFc3XyrZgWxXg73
NT2lMwBREN9B4x2+Qipey+po0QfPg9dnxBHDUgv378AYcJwk9fueeDxbp7PNpcV+
mu2Ucnbcklzln0+cfF34tOAZ80rKRYdGAHCnNRgT5E1/uOJY7godOEB3iMSyi/dn
AX4FzGcoso3WuZhg6kdSOjYTdxU4pKMSM+YpMjrVfl+GbiTVTIPDWMg+6DAhVAaN
Rue0b3uid4IvgiU4QWk+U/LjhWLbgNfynBj6BzBj2HE/KJB73YznWmD5W/85U5Gz
c+2XOy+2W44aPqx5u+lJFkuPqNk7Vrh7AQ2eX0z1ia/2AEhcX7TL7Avio3EsTBIP
Yu/xTLYyarE3rs4TZdCBB6Pt2o/zMYT4Uwsv0oLXcVkJfwArAc2ykYI3VNpL8hVQ
XrOaoK3kwpAOa4MbCULsZhpyptMeU6P8dMKcM3V1qbqi7MqiaAxT64ClsYxMre6s
hbBQmojJjIRDj4ndKHTn+K7ayGlR+896lVovZjtzMY7o4W8fYSOqn/O0jw68CiaS
ibf/OLJBZJvJZ3U+u/8jFRN+aCfuADLe32xSQtHv0FiA2+iC5HZH8GhMtkv8giFh
9CWNDBGpbG5ybd4vRDLGvjPBgpuiAtGhjKuUFvmGh/y0rrx6LChBQ+DUR+ZURDQs
sA+BqrtZGWuSZjk+l2GHGGNp5y9HFmWEq3XN0im5rA0yL+gC2EAxmgQaC/4+7KlF
TWyb4ttvy7L5cp+II9+uRypzqO4j8v5lEGB6x7bh5A0Anst07nkdAOlTw0Q42hn8
RARBvdlKcaJqunmLpHEzeqoWbugjwZB87KlVyIgDSYR479auxukvP7CSwqez8mWs
b07N0FQ7oMwBlq/P7ZKiD8+Fs1CmiLeXqhCFNta84za5y1EiFoLGj0cJkyt9xubX
l3+6JHmjV1/PPoQ6Kq/mojq/064a/xyI0fAxi2zSaOlVntv2A/ixzExhgzvFcMwW
KVlUmwmDswayT4FKuM6UUO7qnw2OXqArYpQDtajf7BLI6XDAzHoWU8v15TqwmGAL
u1Mpffs3x8nZ5pAiJcUbDchkHr20jObZSg4uSxjpL/CfzXbwpXHblGWF8VzPReY/
49XyVY3rAtDMC+ouXm2wW2jX1u2w2bIlvlL9NSYSuZSD8hzGmGJpg4BaNxdNMft/
EQWOrg8NW/Sui5o5Vn9sD72xy7I0l0Z7GVdgGJW49NKIncGcW1ddgS2mPa5iMbdd
XDvcaM+YYkVRzJ5sk8MVQbNAmJwLqjR732POHYJNJz6SfM93uhV8zbb/xSGG7MU2
Ni+dY11+i639fMX7Tcyb7rnqb/5hjdj13alSctPhd46uywwbfvrirvnRkAEw4jbU
6L0CPvMO9csox9Dqc5vlvoBQbrrbEzk+BBPVp9vo9fP1TAp4j1qu/ClISAEr88tD
Ypbv4fkMvSmHyU39xngVg53rj35/+XgcbL3aWGSd+Xw0FgHpIMnTQTkhQL/APlu3
cVY6aKJz2Mn7tkni5biKVczQLuOpRFDCSii3IghQhCqlU0Ob9rf8HRWfBnftVN3k
mpne6lN3THVlV0ZKbzh1eQ9KHkP1NsFaKLwGYYy4OF9a7jkcKOZ28bRjDSSQUI+1
6tdR78erSC4mjb3i75+IGjpKYIkOtF5VmgX/tvrSRT9MoYqyePXHNhOLUeiQvDFO
/+UVsp8ETT7JEbuoDhUkeIE0OtNSIQiomSSIngq49FYDSyPq1YR4np5LeGOj6bAB
9EvVYpYhJlrF5PCDmHT3y4H69Y9CLO3dAzrSS/txrH1Uu1TfyeXSH3HicOsAs39u
f31KmvkczIv3Pd/5wdaoqcEBx/dcYLjBQNL+W2UBNclykItq7g9L2oYncUtmhU6l
x1j80mQPEak7mZyr0vL3zIvFDP2XQuZAWRIy5tYm783HVUCRy/DKaqP7UosMUPeO
oSdtXMwa3rRmXYbOCjO4uZ2juJ64+h3itIemczeSSX1Tu1RvJ3jyh5CWQVJUk4Qx
BoAqtbUkDG2k2PuJAY/8Iykxii+/LqUh4lkBfYQ8ZbUIKeVJ2e8VUt631jLw01Fg
2UvKl9TznhBgUJJUvHHbPOse94G2PrISO4qBYsQ4jleU+qndNxZzpuqRb0cOtAT7
bZp9BQTjx59ayL9mJhvFNvDDDpHX7cUKwUAs8nl1u/F1o6pl7tY7cA+GebuitsA3
GpyPWnaywQFUsurqvIIh2wolWNZl3Jo1NSdv1issOdg=
`protect END_PROTECTED
