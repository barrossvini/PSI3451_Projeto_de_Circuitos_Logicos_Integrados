`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q82JYdJOknB9AVLVDVUe8IlTKlsUGXYqRX7fbRU02WuNicv/r8UcZ4GrTKNNBYNa
uD75Gy7a69ADc2CYmOvO5Bwh9mNTojbLUUkQnsLL/YXcDraME/Qqh5nnzOY8VqWt
s5VEzvHpxEksNA7WIhGUFOet/0x2Y0k1YO02qUmfFospz4JmafC0obAzfJl84L7j
0V4QeUd0UWU+3oHu1SX9h3spZ0eGWXW5xZy1EnzMRGTVrfaWITKR9uBQRpHLwaTB
0vtMI117IbeQZjrPux1tfIDxARPVCZIR7xoz8EsVLhKMp9AlFLUMhNBKV++2J2BW
GXMCXQp4GCFwsTSXWO7377yhnB7DCCb7zVtp/sS0jws6b1/Y40hlMdiSKUon3sIj
MFl1lO5Iy57wlZ4jRY8JrdhPQZ/ya39FigvsJSvtGa+e/f1UUP/zdiKtvjAxh9G3
1MLao8CBkj71AW+rasIPzLGTjcpTfG8KJwA9XPJT/3tIw7pTQywJvR2hCQK/sWxB
+9BCd9MzyXU5JKwisHCnsGMzRzD7RzNnYRCOMJBt8QPtzox3DhoKnYhv1+s95DO1
eCJCiI39Gn9auHnJLfjvKNykh+8Tf/291T1sw+n/Ld6zg438vJHy8Ias2a9BNBQx
7NV65w5Gz7A1PjUNfmUqffMD6pZs3t3uPCjtuY8OwffM2PDoim41vuZazTk00GPP
j2pNOdXUkG3y5DH+/clCF61l5CiLoh5s9TgCJUPbIWM67wTfp9p3soREI1hOQFD6
hbHnO+UarrZ1oeN5LfCKX+RcBWmPngbomlJWdh0KJ64iuUb6YDdqyMv9DzEWD+9k
omfEYW9gldYDboABGBQy12o0LVfWPqctPeDRsJUrb4GKl2mwVIYnEPBH3Oztc/1+
8ENnn4kBf6rIQREv7ZXLQnx7xqxj6rBnGa2f2L9pYCuHeRz/8zryy4J+hn46cfcL
i9x0hHu9uJ7C+B0A5SEWVfh/vf1TPuz8JWHK9lLj6f6UXGWrjGGziYVfQR3o2NZ0
i3zOc+6nhgLVs8Z5O2FKap+pW3jTQS54TMr+Y3IGh3sR0VisYazK++ZAnC8+4O3r
8t2UBOmwDDFLmxbUryx6jrLNmVDFG1GjFhBU1NswtdXZynb2hQDSxQiD4rECJL9b
pgLRnlWwoy2sn0+piQt2+7n2z5/HCmzfz94nrtE2f3JTMK10msz1JCJOEiDciTAF
m1b0AmCYf2tSciB8awlDISsw9/N0x6bX1aVzR5lU50GzkmkC+VUA/8zW6mlF6H1X
`protect END_PROTECTED
