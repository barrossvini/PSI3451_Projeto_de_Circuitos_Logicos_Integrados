`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rJ5EyyBYPGiFmFmTDAPZ8FDjH3WYv/kgWlqu9Hu1oCwlqqgYbqalZqgwA+fQ+ifE
j+uMcizKrFcgnERsBXlXZeiMJVX4LQEn9S/tBVyeU5Bd2JaCx962/VnD2vUIGKho
t9EGYWGWkkU0crqPACo5HyfcbfxA86JqzZ2clhkZOAYrAfaLLq9lWIfI0GvYIzqq
3QPUwdvZIehLtlFWUwEckkKBAm1QksPODOv1Cxo1QUGsVxf4nMTaLUvte0z9ScgX
7vL436YRtTIVrjFkWxHX3KgZHewhLSEs7eM7rbi4FTmMwZ6stdg0z6kV4ny0OToO
DCKtKoo7Y9lVmoZfYiHzGwfAY/bstHKjZzA5wHw0ISaPPBtMZnhTuuBP1nYbUGS0
7AqPoVy8GUC/RQ4Zxvf5Gff6rCcgH3dqLfr1QRRQrzaW6RBCmewozDTyldqLf+rA
NJ7vpjxG64j3vECL4uZFO4CnbMqzMob0Qtvh5zf1Ey1ocDAGUPbS3DUTgEAnGoW8
`protect END_PROTECTED
