`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cLhTLCw7z8Rh19lY91hqgKLO9ZBn6U2K+baPowbcetHY+orJSklMPQ2spdz+G3ls
GQhMv4K0ETNxuZnKDZbxFmk2LWyil6fd+Yo6hpZLQA9/Ri72XRn38KwsWRDKCJsE
dGCpNk8zIWEm5uD7Btyo5PPGPAH9i2IhsuHIpp5jWfpVcUKZKIj6ui04yz4u+st9
oSmrGeNsg6j3Hq9jIeeinU1yDCl4azO4YCqKpJ0Nth+XSxtx2TfCv48yDnBtbBlC
MVj4p8DqTVgn0R2cC/hNSIlwm1xDnI6K1JvY0KsQV/qEJzJNeD1UM03bEoutGR7V
zUXu0NsDH/rleSI87ZSBEJbC+Tn/Z8NrNxChKOJZ6VTbq5tzBBflQC503PJa4N99
k9oAIaEqXRpI/QGxIdDoh9maVs3ptPYRM4w/CBiRPyltQA/k92zNQxJNuhCfvv1L
WeEmgyXgxHaFTq7N7odoEUUYOfHfSfAIl6wXSmIxH1cjX84Z8O/F9FI41rxJlhxJ
NMBb523r8aFr7ldAjbuFrEDZCaYleLcm2d1xDwaUxoGzL6pUoFUeP0Q1PbbbjE+c
q4FcJQUzNDK/3VBZCM+yVn9ID86XkHLOfxMg0GymIILp797wCkuX1UZeKGOai5OK
lbPmzXXDBr2TWkBl/9grZcwx/rIcBAoK+N+297jxVdPHFyEYNGRdEgp72K1jEhf3
WZLmInybyYbRi+SP3rxJ3Tpl0oOSPKAYR34TU3MqrRE03pvKUbfjyiiX2NAofT+h
W2WeFou2PlAxwxzsyw2MJiR2odq4XXVitv8wLWhV1U5pmH8+NRs4sNBJUKJindZA
xCiDzdS1M1Tcl9R3gHE3lkqNwfQhvuUIVNIvPeTbSXq6athaJiPPVKNxxk2sW7+o
4eBXbbzF/7xCz1pRGSYbEQEnti4wf2T2cIwmKsPMXSSbKM4rPSW1/hLQsIpW8b8y
J+Ks4I0UQhPBwxZbmm3ZjcnfMSRt+VUOxpwwuz2I5Ss75N210UJToJNPPoJMtBMh
U03NmMgzOt5CIQuRPIXbF/ToJSrT5VMsuc1OR2fV8jgXWq+TsSeRgSClMhPS/fbQ
7NIc3EB+devRWDQ5/GvA5MuPWvRfdt8SmsTEZ8meg0TP+MwNzwFTwI+GF1eQYUIx
RL2avJug1cZhglinxU8JBfCR1BxaMs8HbsVSNoTVq9FSoPVfBfhHWuNl0IR5Rro2
c6V4l/6mXJd+pQrJDuESKCTwm9IdUJI8aq5cK45ParuwyOvB8737TenePzsNpcOK
1evzEWcPCoxjEl7e2VaFCygZVoSl9kFjchc+q7kp24KQfvxs7rE0cc/vWldMRD2C
R2Y1FwdKGye2PYoQPX0yFSrJH+dRV/p2IU2DFQ5n5PY=
`protect END_PROTECTED
