`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CwsjaK45RWCAwTfW02PmafFA6FhTA1FBC8qo65NHwd7+QnPDgTmstkWg41sT/h63
qIR5EGAUbHR6PPppGPWnGqCJluxlhhCxJtXan16KkwgWH4FQ3eBZxHj8ho96ewKS
KdkH40Rcua8CPCpGTgsUUo8mWz+4/vDaRwISGOzXhcUao3mJMXvrw7bHnJ0IBQlW
xRBPxIcO3HfdCrZai1sKbFyjprk3MvUcq22dHoU5n9DWmefOj6XZLYRWKOdT7IRG
cYQr7iSfwi/DpFw4EChGjOxAPBr4JKeI2mrH+rwehLr8YDfqLpdNf9O5cHPbM1oT
16dWX8mzQwGIRi3df5Ypyc/1VfME5O/Dcp37hx97/L4ftzVRXmePMF9ZibIpIQ1S
Gh/RrJzgyoHP+7wdVl5ZKK9whnF+K/hU7eIe+H3lYh5UdK42YtGNNwo4g+QPcRvn
nZMuHfKHXY5dZ/XlL9EgvyZIpuhkyQ1VMpdXSKLGmFqZm44IaypUHSWminvEPdbq
UaHYBwKd4lLYwuVJfmAoabxmxq+LIiNXOPlJhTFfs0LjnSdb3hDjRT+BlL33SD5+
gnWQcUhU50EIicPLMJm3oNvG4ZyLXbtfwkuSR9lxP5x9EN9TO9eo9kDDsCpG/Wgy
tw5l0Ia8qU6ZiDALOW/9V0AwHqoaQPUd0PD85N3FZMCxvsNmf757T6BSF78JZ9zm
8++M3bOXq42jvc5wp+CxhAL6IR/4+/FXdI47W+qlgTJGVwrwKuoZyYFfmKRr1bcd
/V9XnqFGoZZW4rxylx1Yqd7/9gW4mHER36I1XtBIVHxFxe0Fhh2ZO5+ViDssiEBj
JtGWRmn1hk/rQsxN6a1LoAYCM8uLSGqrtAOO538xv1Cx9YRUgmBud8L9iTLE0Mpt
VU8f7GQKPsSwkAkhUp3dYkWGQeo2Nj16yPj8wBYXCgDdQe/tccRRQYx+UgusIx5r
eX88BCdTDSK3wapWPATMniwEHb8+n41ahR4+SW3Ff6W2f74+odiBhCDg7d3/ofdV
UhEYQFJpRImHdeKkI8OAAFPS6HeULo61551OjjFk70hHYS6uNJLJxvO6ZMFSmwsj
palobm93lGkiSbvuysSH/zPRayCEkMhNgMUZGHtHhGd9YMrS02dnqpWwLYF5t6Up
rGav77xIUo4DUHPOK1YM7gQnwp/zbe5ceucecMcDI2r0fiQ/J2Dh7njB1H6y3sEf
x7ZQ8KvBG8q9wExb82iNrEsOzfiqYCqrexGyeNXli9cpRsxwA3RnO0Km2T98+LDS
KoujC00rabRIS2FxuxPQbswfwn56fJt8EPlo/WLNVRECAOMOPMr6/W4Pe/9JtEKa
zT2WNbzFNWEXjCwJ+l/i3khNQbct+J4XCB6PL4EcCAt0JWMh4A6ziuhP5ubj6bgV
IeZ+emUTqzXZsNeozNd3PA==
`protect END_PROTECTED
