`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
elU1DwAlTVvBuHHch8EzJhB/JTTMLdsTYrihoFpY/E1xLEVjBJvwPLOeE7wBfFqk
bZYBy3A6ceucr2W8p0oPgiuoq7qrfaEjiqdXtSv3iVNUwg8VWPMT35b6uZ9IcwE5
J4xauuniMus1R9Rm1VxBsHPWg6LvFJFvSf91rpDXcpyDvk4Z2snpSlCfFGXScsiv
XBENcQmhly8HoS/IKrXhKuRb2GtRTd0LpV44E6RjZpbeBt66Ah9FWEn1u884Slgp
IIMOjBV6aSZureCwtFmUUOIw7DwGWfB2VCxsmeIpHE4tUCNUPxGcoCwQRz8nKaQz
XWcZdFsZieyVdGvNQKT+BU2EWn6cZP7F7iWq5VzTPFO70ZvYsUwBSoWl8uf7k2Xo
u0IaQNsI7sxupqMEFzrHoMxKmBF5aC8wDdobXvpjXvIKsYgVbLBJZnlYkGRjj6D5
YVkC2n6eVvugYFcZ1mJuAnQ97Hup4VGw0ufEUGzLmP8KGQMsBWe7IH9Sb2XAfVu+
0/8pT+EZy0CmZCLrZ5fSE4Ilt383/GnhalRF5uUvLfl2/p5D6ON8rPd3WwsZOhr5
EZnWCQ4aTe9ym6CeJQaOSZPOX2oaVMrpLTbnQbgBC49dUMuXtJE63t00Vg1rMWiG
WvCPqzA02n9aJ1BjCOrYL3kmAoRpaYelptVt9H3Y+C/s2Ws4ZU4tPRqnA1angdlb
ocVwrMnThW4AMCB2yTeLT2ikFv77GSaByS96Lpat/UOEJenGTVWTzZMmCHUXDaXX
e56ICU6eVP8GA5aa94iGwar/MLgdN8szk8iZWwIbOfJpCo8gKPyPVdm/VDCJx5rE
EywMRtZZOgj3+qNeB3JV7sUve3mfXxzwYm464Ao7TD11s4ivmlR+IjXr9GQQt/Fl
FYHbAzVB/7bYdCHCZmdgHQXS86WwaOxI1scgaizkuWMdtgHqr8igpCHI5nBYochk
Ft9L3Y4TGU1xIC612kMBlYSCqeV5BGKijN6gk5cPwkarks8R3JPdy15o1vTWUxVQ
Ia3FOtbsvlqbWJGpGbtQAt1FprWVncl+PpDg6XviEvSBQmUea1D6kp2+IAmw8Ivl
1xz1fC29BQWB/JFRgqdkXb3B7bUx4L8JxRbzQr4cKKEFK5/vztlIPV0jC0wV/Wv2
2+7LuI5eCENl2diRu4zUpcgQslGsKfEAzcn5ezBDQfeqTDtdTqDZzMggKbLAJFER
URoC+QzuTTJCscraSUMudUT+7P+RsYEx31bXU5/akXuPzwdPDqsDdYOSJgVlVe0G
afMp0JWoG1L+5lcWrTbHFZhu3+JYTzxyI+pK81F4/mxdQCZyADralPm+CJ4WfTTN
oS2+cbJfzlXGKyQ8ih91CbrOOd9i91wHPG26+pAshD4NO9I8EPnIUaMhxwfSi6Zh
TMkV0zTvuFrKpO0v+yLuaIYifx+Ehr6kL8RFCkSVXgJyrYcH3QwKwt4FFqKgefLk
`protect END_PROTECTED
