`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QFVVt07TZBftnYsfTSt3mVzctmX4OAm4Q07uVZvbYnOAu8apOf6HjuQ3OlsM5kC6
xAAU9smnqaLqYUs13b9Qg2LlkN7IBcw/rsDB+I6z4hloggf0TF9pJ22pTCjt1F+B
1DE6JmZBdsI/ZYefe3g+M90t86W9huH0iQkfACBcem1zM3dHk/+TrpYrCBSquIyp
uI29yw84dbYVBTWX3VMWh5lt5A0TEt0r4n+ISvRik106rJePNnSmUzADEpMiEg1k
BTEzC2QY6xiIkISDzmQTOITiFeI6pVP2L6xi3YrUQJfpOP/41Rpcnvuh2ur/u978
f+ODBwV/yO9aueJ6t7D9g8bKGoFJUKGYBf27oKtfbcTq0xRWgaEmjRocs3cSIZkr
wc6alTCkXhlJBgPBEsIMhB8s37Sw2HYJUsHSFHX+my6bpwWqUa6UEFGZOWccD0Jz
hmO5pE+UAzHM8GK7U9kEjQH6yF1YAmWdoPCVG4I7wNsNeHG+J8X5Rk9aIM9Ft5Vw
nt7y6MfZMD5kdf0MMrmJMMTJw/l3CgjTi6Av4n+jZEeecsnu3NjR9kuxAvUMWNaG
XGclFsoweaxCwmKXdlCfLp/NKWpdA2kIbllyfAHE5sC1e5CdBKbglFBImBo1i4xj
qCuR/ZhaDG9G/SSAuARODl5da4kQtJCffNKnh7XnQHqrVBSRBm2uJohN7b0ZXWb8
XuEkjy6eyHUzA6DgF4sc15vLIFLWJEjmKBPqUN6wqF5vBP75PkC2t7bUjEhNwWDL
n4Fj58F+lj2QIGC6MXsC7jUr1eePLJ3aWimni0DDYil8iQXOT4nQVjuwlzx74Aby
9uOiOYUwMcwLPRdgLV4+Qg==
`protect END_PROTECTED
