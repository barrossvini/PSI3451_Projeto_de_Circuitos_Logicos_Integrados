`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qywf+Rvqs8WDwxX3HxA+7LUs2fEIKc5KWBgzTq2AgOGEkjPfVU2MGLiyUNy+zBy3
V4yF2nZqR76hK4hO78L8ZME6Sx0swSGJzk+uzKMe7ifnxC9zAsGJoh8Pzll5lr7z
Iopey5BLIoepd8j9HIysX4ic4SyZGr7Lbp6AacsUIvYZClY6c/5C0GxBnDiWQqRY
RWeC1IpP1EwyCI7GISZ44KM21OEm0m465nI0yhi1N5tEjOUk85kd3cxDHmPnTQ3Z
udOKO95GsHI3qkrofdiZYczaQpdalLWUHbegPSwdeVziaC6Kj95CswNlSdkGsq3g
GNnJ3tHBvG8Gq+MAkAmMnfH4NKA8MhZtkEgaiff4X9A6AwuJZkhKuUh/LRzf4+Qk
CA4KLLbtd9xzkeNnHvOGuQsDKqrKIAHh9GiiiapuyH01xDsmEg7Nh5ACKiwsA8p6
rVQHpli/D94oAhdm6XLhZw==
`protect END_PROTECTED
