`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gj68hH6U5tDdz7k2XZe/E5pjvHS05y3kfsaxQPecbynwCp+tIhrhnJkZt5LkkK2Y
uv23i0I9gMI66QDKvUQ7aTHtUzZTWvyx1PvLU3Y9u+gCRR+w9gWJSWeFEF4o1Hmk
v3ZtY/ECpxWNYd5dxuXc+/cG6qZ3PvsLGYAbVdUdy5+mzJib3NuTpTrf9cARhdUD
s8NnK9ghtVwUZS9Kl0qwRBlpGwjwDFETfZb6JzsxmCD+dhCSaLRr5vEy65Qjbrn9
qfEVjtHEH99HOHNQDac3MKuUWbEyGgTG3+fvJOLZTiE9YUlN5ij4dOkGBdM/3+kc
KqghtI1LbD54PguwWbWejK6+8Xk/MXc9TKZz1R4CBjvmITnnWl8U2zpjxvM/15qU
7O3bPJaru77z8TH1XGrVTFSRFavz+SIrDfqbl/8lNa+9P2KOCk/mV6JFNhMyu/25
ATPknhJIP8EAF5E2dXtGv7dXzOVLExEqqsJlf7szDyc=
`protect END_PROTECTED
