`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKlSwc5oMeZiGHfZ3RP6snO2JhRIws39MVvusPloARZeixflnwUv4lFsSFl7Elyw
d8Qz0hrp7Np4EfwjQ/mLy+VuAQs+R97Vb1dIVwpXN5EzxyuRCT91TlrCk6972CWw
8lvE3iUjdRXfTvyQoriPVq0Huml6UlESBDGBVbSSogdZhXmBgacw9SSM7nJP8Otl
T0ttPDHSbNjxaaYLaguj9W7kBC6wW85T+aKI7LTtldMtnUjnTZOQAulT8aiNTd9d
OfFXIElcOKUrWhejKpGscMcKEEvNbqcbSzPLjAk3+pdslVuPnfz7ga7UAM++fRUj
naip7HVbnkdFIaVI5rukozQtN/x7GLAUfFkLYqRzisr5JOmliq6357tKlDhvHfgi
nkAimu5fN4YfBRcnTTrai5ft3pciIFLJOVZnyiPfbzatwK3Nii9p8G+K5dY2rdhh
FM/gPlKKEhr7Q0fUNyfLXJpUyNqC24OjYVO3pdEWrOlnqm7EIpJTFR3hGWQEGWM1
EPDHnOSNfq7NOwwvE83HtOResQryLeMACeoWZ6fh7pM64nGuF1AgNB+3eqZgSl9p
pzMc/IVcmjnzwc0TnaqXRvuoBYVe+xFu9CCfpTj0swN7E67B6Nj2+Hy7+0/A9L04
KEG3IAqFaxeOyRdjd1beBydrcG9puSl24dpY8NPaGcDQd5GTcl5AFzs44ISx4ym+
ggTow8VEVBJ8q/OMunlG1ziVAKeXhaNOQgfAyTPorNKJBhp2yZHxaCrGvtH1jAKz
yAkzUuGcO4XuHmj4mbHOJymKpIk4s3IFG0c1i+15PgfKLIfC3YuwDcF4Ys4LKUM7
4/IQ1BxwWl2VGhap+aUwsEfW65gCmdAYrAw9aInnR6B2qPedcC52Lopw+l0BHKHd
CP6hcZwW50W5d4svRXqBuVE1RYRNGZz8IphPdoAOYpLiXoIX1KaWKMhvUQIC4Z/f
AkapLi4/A3a3kbO5u4/PVynIlIbneQAGQI1PxLhp5MklA1mb4U6409QQegWLbeEa
Ew9bXlFKDvYKlKWQXCONYVdxnzAr7TI8QgMGBN0w+YEsaCp6cqW31xwhAsNrTA9F
Ow7foTAt9JZ2QIsR939cw9HzIJieFjP9/cScAD70JogaImWy718yc5tFppioB+Wb
Pde5rhZbH16j/DkoyxpLviMgC7xuu1EEtVo7r0o9q45KJ0e96J8qNo1k23GOG0VM
RuMoBcJW3FFczGROSfPKs+Fk9VKfhkxRzf/VeU0rj15GpiNpUkMMj6hOZR7Ab5if
fkB8GS+NVMkgTIhmZgj3OscdR8nFXWjrF5129LGvtsuhgFsHflnrts3TXJkwiTFL
GYOSbWxpgwpu571ZXrWhEC39G08bTG9lP4rHaxqw3q1/HMp4O+ZvxQFJtNmgXcFn
IWY0FEN55T6BwWvhZPmUns7jq2EF2chvhr7PxT2v+5q9rm3j7GQ5Vp2KQ//Oq9ZN
L+U5yRFC6qqdUvZi2GNZSE2a5dZbc580nXf5b9fL45cN5LvHRLX0JvHFwMooBkDb
fasYh2MNHy/fBKq8jVou/jVona/qBpV9zjptgZ0vANvwNZIiWaTHBmLckWtI/xAj
PjEkeCu9IPnhdy4Hq34KHFDx58C80PiyJAr4biwL5OPIYggNFn5SFOsGV8JhEEX8
ZmrvYtX5NdcuLO5zu9yLE3I3oieI0PddXHOlxIqxWikZemd5TAPulNiuSEy3OLVx
d7I7saWMSyQuuLbZWz0zub0gYGc3OqWMbUku69Lf61cl6laD9R9TIv6NeyNMMRPJ
IFKF12piclQIeZ3RqbpoWmAE7GZ1rz6F+V4LKll8omKS1i2OiKu5pqMdR4zd19y5
G3h0koKD++2KTm6km7kGQ2qehyO6wzEaUOaFDxyIPAbHJIljcOyh+MsKInXxRMNz
Sec9mUVndoPiKTSKyKDWIu5DpNzJz1PLKNG9UKBIcFKAiGQeHuErQDW/eKnjjJat
5TK3j7/wbyGa6Ls4Qzj5dUKNcHLlsm4WvOWe1UfRBqgsXna7TM3EMBCr2ffqvBV1
u+KHBz5F6Vtnfy9v8uPJAHuuKIfR6he65WKdYJzvbusDq0daEA7sUAMaH3iYK9tS
l+rJCso98RF1EcGHAM+Lk0gIJWf2lvYNh9YkVJCpD3clUTFcv8PmqbwSQLDK1Gu4
r/EsW4sfKd7fNv5BpDgHFvhO2oO3HwP6zt0078HMSecSEhaoYh8BjhrPbLWnmEGI
+qC+BmKyVmcJuSXsDZNr4hvditCov9dfw5C2KsZRGcQL0YdiNAmviCE6R00uBok+
QZdw4bLRvIrWVXG3/zC8g440LtIbqtEWyZgc//ouvc5fxaxFv8vwJRwDckMsDipg
wwQ4DrkR4v2JlaVG/+Sz9W97lhqdS1I8ss3WYXeLprbNq9BRiwmJW4Rj+Hq3zjWU
+AYfeLMVqHurw+PudtoiXcgtpfeHQKGloOyozi099hyQO00K/uijaWo4NtszsBPo
+eGCUvYOMzneLcYR+m5L1p5fjtmAywheFlBw7tgxGBaxODTE8gDr63dDXU66ZYQR
t8ten3Oi3gCKE/21++sVHTeNZ4dsU5QCZCS0pFxi+b9goorqyfW1TfCulL6H3xko
p+xCr6Kr99KL6+Gt9iYFwrfhm0rTYVwijolqIY5xFH7KdF4OBmRhSBWxMG7aLcDN
KgciMpEkKY1zuXWAolWE/4K6FKen7Q6CvEx2JzZdu8U4QXFcKXM9COkjBZrcSp3l
EUrHdHFGVG+d6ZFrxV7N17f1TPgqKCI8oGOQykvdJ5vhmqFlY6eZVBu5eELcFkOz
J8Hwid9OmGtKuJVnAzsoFjfcGbsAbsayM4mAgOI2fukArflOWpZVIJ4Yqq3clOML
PffoyTeLJspBexrCFY32XnNqUx97qkOKnuOcyaLAZTLcT8QlaMNE8b0XXGO3EGE2
nviAwDEwoU2f6xB1YFlxD8+iIKBCqEzzF/WZiJUvQRJIIiwBur1240YYoMX+c2Nn
57EVI0ZV9osh++pCUyU28PzCxlqII643MQZBYU6tIo0ZRr2O1highA0FamjxneCZ
oIIzeTS6uRNuJ0NoWVIdS7CaOdKOItgRCdOD37vK6j330/Ja93l7r2veqAZJmDnc
pvpUemQiUZJlPKfKw0ldHnNYKqkeaSzL4dpP2byNEEk3TcoNRMwosUx1r3vxqm8r
1mbNjpPta1mh82EfWYs80Dyz0Prmhga7JaiQuIACPHF1v9UeyG+KamzPkhLnPRRN
gn9B00a2cgCz0wM2ojPaRliVFgZMWXeqIAS7wWVi6joJE1b9FDD77lGA0uB1As+2
pS2JEiIBB0ZVlt9Mniu2znmfd3gLrgqzwxeesHR5Je6J3ZKgt8aco6n7jsZGbnPE
cklJusN3FyCVO2c0sKX63Av4ddYTshFh9rcsVI8O0ChIkmgmVY8Z4q6txEp8lFqO
MB7ZYbGsGW3ifP/rhXn6Zcnjme5H3x4BddzjaaeLiQsdmoNPW1fBD53bZDS+thXa
B9fp32amVgWL1kgWltYmndTeZC1vueqPqNyOKAwnIcft88PDHK28OqnJA4ok1VLm
Pl33aQBy8rzxXUKzLQEGLbiBSn2mb2RfBXOkbi7DZFTGdxAUHpM2TS+LYCjjcIRl
ysK8UK0CgZRlnxoIH9PbKCRl179ddfhBOG+60Kp066WmNmmfXSrKIZsIRYhRxqzL
Was6Z5rprW0LmkR8WkCOaTUQoSAj8JoZJFmvnZSZL5C1jIwg5eidWYNpCtk86Xz8
afH/01TMcqygYHY37zUtBEDHcXIWZ0M7ml6Z6d6XnQUDm38T25hibLTE3xIlS2vn
7J8k3DWlZffd7jhqjy3W634mUkeSdXUAjwSylKrxeYs2bBfXqqd65AIGqzrjkcTe
7Kbf/IWV1/dHb3JbgF1k9r9egkEj4y8skyCs2ClfxQF4KBOqskFz4/xdbC2CKt9w
06UNxuu3jqtRMm8zvVwkIc1Ia8Jw5o5F/lWX2KKu0Fnu4RtBnhzbZXSYn/znRVCy
aN3Oo2TrUGkuU3Fi4yP3lTcSf1Kofwp/xhYIt7dDHA0zfMse5CA7MkgFTSjoyVkA
LPRmER0PBVr3IJ8JKR3iY93nvDDa1WUAniWydU+S+6OlhJoEZEjGdYBESC4QzAPd
ZOcSYmRQ925gsxOsbRMx1PKsLZVHmBlOxzlRcdvdnIn6SOXqet8KW0tSG5Rkv1ON
bkvUPjyGVygOLqsPpvJ2kK1d3wpx3HPm+E+sX4rKir7k6pokIGq/N3GDdRNFuVqO
enOLB+2BpVQpAaW0L24Q9LFaMTO+fRqKYLGmtjnreE4YWNiRbimyFa5dmNFFIfkc
GTMXGA9JFiOLErhEq3RROL1m+BrvxJKm/OoIcCD8tnxqcWJXSfBl53ffxVBry2S5
7SI0Ie5arg4G7GIDpUe9z0h5sOXtL3PL9qo8AtRrjWXWWh01NgTC3BMj/tgcJwlw
h5lTUQXx/Y/WKAx5ZH6D+/gGNpX4c4MQlRfXkj5K6xxeRydAJURYmmkW2eDY7MEV
H0uWkzClxlSox1/GO61/jTirKVo0GK5+ZZbPa196jhG4oyPR4lCYPuxhRwArnfzX
a7ZRB4x/ts+mZYksWaOXgaMh0xXPCm9RoCpi7U5t1sm7OrZS9z/52Dh6J3UTVja+
1YlawyzZC2qNDYyYH3rXoNGZQ0bU65PfAJSsNzK3a0SHH8iKtKsMSOxe0YT1uFd2
o2JdFPx7QZJyIOFFMcSP6WhqEWqC7Je6WlOZERIM5y/+W66dra2jiU9QZMw0tu20
xLb8nvQPUieKVFVXHlTiGGZpQoyDUM8ejJepFfnCMheTtjYp0VwGdMYI/EHLUiXE
5SyhcUQYqIt2KBqbOwHZ7+5bOek0HwCPqw62hiGvAv3HhPYH0+wKtL7yTtC8JcZF
BFlkhO2GlH4vl60Pe5hW354zwJX0DSceqvldd+GLlZ5nAw0oSEzcMtqjxbh+pX/j
ePLczqsLpeey7wVHMhrF1CqDT0RgL+LsMfBbiiJXcket5oegMkdrrlHTxpbCmuht
Iw1Uuj1GY+NOubOpxNavyQe217Ag5AVLK+jLgimeNX+hp/ey6ZlsVOifWW7O9wxb
MSDQnL3o443/6g07DIwDPJ1I1PsdY3/4GgZ/ZZoi8CgDsNC+kV58fk5XA1bDShoF
purzQ6axj3KK8la8/CL8GSvarh1UAsRUA6Q71ml5NopTK09oi/NeubI2k3KJSqW/
vATwfDVcoqKgwKvxwqCJBpVf5Di8ZJl4sU+1GoCGGxqqBJIX/T07TbFJMJiS/Dvr
7za285KsmM0wTmhF63I5XyDDqxJJRI6Kew3FRIqraLAGE6LvSbsDg1MCQJjFPLRA
K13zQnMIS6njffTKj5eBYdRGETEHW7ODLPAfAM7IwM3uoUDy2NoAVqnG9aVuowR2
2UXt1RKPwN5HARJpwEa2cBz6rJcXTjLWYyBRG3+py6eYuvLhhRi+aeY4/IfQFr8e
wsGgpdXOpnCkrmb4YrY4A9/ZOJJs0byQSumQaLiYAsvip+Q4iLZL5ZDK7ImlVL2H
/ycX64DP3Q2XJPmHm6Rvku5OOh85VB+Tg/gbgnwQ9qogOcwBHRAZ9liqPZvmPrRs
vHiJczRHLsxaxpgbeuqYLBoPQIo9T7252s6M6uNaSS9tAFufASMlX0sabM9AfQLh
bFOiA24ZArsu6rNYsD9CyB2kXAC+a7JyNGl2OfiswoF27/m0/UWjNo4AJL5UMpE3
NQqbPA57nRvXT6hLRllMvorZu9r5/zCLYS3WO7iZQs2mHzbT0P9usPqjdN+eGoCm
dOclvmbB41RPVr6cIDryMRWWFu97oXL0ubhJvTfy1KjV3qlt9fhf152HiAnxdSjK
Hlx5ynsfTG6qFRhKhoJpFsZN8OUwFmxAVJZdNgjUaJ/BNTFrrFvRhHK0cRsbw/qe
f0o43tMgH6PPySbKkbSnLxcpp5hA51KIZZWnSUJgljlV9lFYS6WEnRTRUVFT5JiY
0h82KM2ogvaGFerQmXENz5zD5kne/wkpVM8Fmo2jzcXYSv9LpOwZIppPolQss925
hQ1HaNSWo8V1qBKs1YgBqCHjZOIBYhs/1RThNwuyiF3qrCPEFgHFxgzH+C0g8yaN
fkjOgj1QX+VOEBwU4GxYyfNqkurGaL4+w0ARYUzWPyYMqdjROdaXuR3VdDbZE0lA
a4wp6dHR0UotInnGjDTdYvzhC9F8jX72abnr2FLD0Sb3QB2/0s92xnzRgFEZXNO3
W701BpKEzQWFXF4ygL+Fonwe3bu+vypwpof+D6HOIUh7z8q6f/RSwnYUj/gMewD2
LVazMxBIF4ZXDjRm9QasMoyMXu+EbAB7+VyEie7Nfi3Zmk83/QZi3vriFIKoq/H2
L7LrjZfY8S0VjlzXwJ41YdIQvEiGuZ2b75P/whLKpfXGEva2xV0uPeo0BZN4DO1M
SDhRDCvvmz/glh4RXd7eCYOgZeYMTQ/W6RBdEOasWjRgjDDRZWTQ7FV9DQdsGGaZ
WlGu+yURaOgI9a9Sogp2Y8q0uR6WHBQy4fR3WDjclUMKFs0cC4HItVSgyvOLl6jW
nKJY4ib8Ht7fBcmSsQY3pVEPOs3VZ3fmXPQr2qtIVGXEvHt0rz6UHiklC9HBsPtd
2KJhDk+PiB+KG+sKwwmgHzXuwwQaJ137O0VpluDN5JBzNHDc4kTPYdHxfEMzIlXe
hY5xSBPjeULpcxfZSbpAgpgZPqYJecDxTfon1zp2C60=
`protect END_PROTECTED
