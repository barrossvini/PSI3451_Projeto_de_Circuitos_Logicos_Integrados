`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LXYsgn6TC+Hd/XxGys8U+w9k5WF3NsNVpQs5fi0FJ2OlIiohT7vduA3ExMYV3Tfp
6VUUNBcQ+D9OSP3TAYZRfoCGexoKDEZGnQfkAggre4jT+yWrG1lHsvkOX+ianI9N
CJpYWW0sTyImd1Y+pwgGsf66jyVmCdvYcgKFLXq7V4z5Ww3wQpvpF8E1nNdd7wSM
`protect END_PROTECTED
