`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IEbawcBFVwzpi3l6TpFfLG9mfq1WPNvk76qFmLQvw5iIac4OOciyUQm/XbSD/pTD
yHxrcBBi5pEvM73f27s6e7j//Q9YytTUpvEhBAA6Q6Br9YWsYFDSLNqmx56VGSRL
kiFDBbvQYtwQnC2AiG8acPXe+1voVHMLmzg1z3VQ5+0i1Dm59klarWBeQR2qoQs4
I5Bn4mLQJzMoYqk/Hgzu1uKdO6+NkfRghsASqMDXw4nF+KziTgJTMfqYQHqshcrK
HyxLJ7ohFH9NyiSKL8pDjs/RfA7+hzzbnBFCTP4kDgVG4J0GE2BjT9Zec4iQw1vo
vOYIyFJyfoOGg+Xqtgi+5Ee1UUUMHoOVRtrMibpUfeI9hosWyslYNHY6YNrFy+Q9
c0deu9aXw+TKcjqmwmz+m4P7wKTOPG93hX++IEP86Bn7AYgzb8tTko3VV5ytCoKB
jXAteAU8YCRCd2SYPW66xH2df8+G1MW/OStC+5FRIzzjnarlYKCnhANoCDKU8Bl/
mbBq+W7hxJho0N0MXKXfUCue/xMbfbdcc0ELKaBddPQcLh5KB+a7FH3bXU6ow7lh
k4wO937IL3vCHLfuZePuv9+uHJXMnOWtyedL7RsuTjYAB2Vy0nX7X9QR6aYeLiT9
iT9QAQPuJzG5dv0B5LKOaIl4WqEBceiHoQUAmrCyygMPIz8XXEUnOzGZ3G/4hF1X
QLhKGmW8Y1sPWbbDIWB9GUXmqUhPF+PF5Jq1JMaor6A7IFspx3AzPI1YH80EK6eO
+85mj6wkWtfJtZ3VU/GknA==
`protect END_PROTECTED
