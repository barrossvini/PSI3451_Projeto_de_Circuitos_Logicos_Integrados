`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bfmBuAbFC/ipF2T/TqBzmXYoPvnuBbENeduH1ZsTxoh6dUnv5rB3BQU42lEreO2Q
6l0AzdwIvIGq5CE6h1PnrscQzl2G2vUw8lhplQV1qXviZ1v9/VPMMPW+be98+jek
1xImU+SAAx3Kb4OuSOTyI0dnxKoCuKy672HLriMwsmSlRc9Uq2M76nPdUghImtTE
XqUQcv/3s1N7j14RElgd7VTrHjZ9FP1vyBauvtkL8Usen2oRu4Jd/wvRAUrBJkD/
zQ0YnkPuuK7+5c1Rdr/Wd04D0wMPFT9h27eQptFVJD+AkEUHslAgnmURuaRg3pLN
tJbX+4JySefzijyhHTrxhUynhXumEAB1i01Ed4qZLNk6VVkB2uLO1IUoWDWsg9ce
ETDfcbX0TatctnVzq9zSVz+5QSKWP3m/M7R/Of19MBtYFHv73Qf0Wbw/ZXr5WpqA
`protect END_PROTECTED
