`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SbHrVh1NPRRYAigV7d5b4ntPOIJyOpdIHhvilsYPjT8HQnVPDH9FPFJgJCRjB7na
AxwJGfK30fga1eUiPcTBMSvhVClIPJMA7uVwj8aoioe9bDHKk74l0gYMFsWL/dUL
FhZ9rOpLaVXvEWqL3XCiMHwKxXL/I7Ci0YjCM3Y5Zdp91OaLsv8KJI5fbo6LVpnP
y84KyBLzQEUXe82IHEem/DZT65REsplKsY/bFEAMwjLNaZQ/4SAk6Ss+ofM1EeGt
vohxoH9khc2PGFHW3MMxFZBO5QSIrWiaKh9bCdgcZj6kXPq9aQ2BDENeM/Uov30U
5hGkyRaeTih1Rjo570Tj1wzZOg7r/gWsTslmpHuMhhAqPWlJelb6NFUmaEf/iYi+
1oikUeUcogcihr2/x7sqP+89ZJe/WqnzZOLVo6dvLS/26K3BjEvSWvRIH28NTOI+
N98j1p3H2TuM20ZxbKMCJZzwJEuQ+F8TA1w/fjXT3msNHddgU6P3fcpz0PoXF7WX
jh8bsY1NRJ26BS6OsL+TtQ2xS5dC42uJkgTWXmlvoZuafPhStn/EtsUmOqtrfyRB
gbzdbO/k0GJXMoMz4omPv2DhQi1SleppywMbYKcBuUi9J4USHNO5EQaqND9TidYV
itSNWWZvejT/v3XuPaAUJ4wIQU0hSEUiL5dDN9egIYLq/LCizESSwMklg7ukN9TE
`protect END_PROTECTED
