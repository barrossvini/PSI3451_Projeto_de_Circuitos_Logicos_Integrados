`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RKOHI6sSEc9fAyJ5E6th3gcvAYaJdLienrRxCAw1vBcEIWrPh6im3Pb3IHUg1xj9
1v6pkxXBpfTjM2iGq50DVfsTKQ1jw7nI9u3HBtP9SygOvDyre1BiGuusI8Etfs8e
yUNdGa49WH3B6Th4SWqfAE1TIjAvuZI9w07V+WP7P3gkZQUqPSP9uo3wyvkC/v9z
xXAY2x1nfWMJ6wRoHnAGUURghPjqhEMZF24ht3O5r/lZrhpkn25Va2Udr5X0QdlI
T2P4H8bZypLxJW5qOTHVgYIzE1gk9FuzwmmRhoP/D4fGo+6BU8UDzNyW7fQtpn+C
2DKph4TowRGbzYJ3aWTQa6ttAED1iNNJ/ipoKx1gvHEHAIFndqdnrzqpJdcq6Sgc
wEnppkqNlGjPDCYIE9yyqLh1qLNO0AJ0SSPMCNm1uuzJ6wJtm3iJgUZQW61xO0R5
HLABiWFw3xGEQeeiNHYGS8w0gLDIcBs3W+JQM1EMyS1W0wccp2P3QWd5H0jR8Z57
SPd8cjn9fhh+wjjphM+0uRf2Dlz2okMz9u9nJEQ01JdEJilXr9sR/i4RJ2RUW/wO
eMuRttqXYUiOjVYsancBuTKK9bpt79p9yTAsjP9YqiVrsq9XGwiM7nyI7Q/xGkiU
vdJANOWOGeOTqinla3nP5gy1N4iKQ8WJuL+kUyH2H6tdOvlEwXODwdO7nhT0+DqY
YdplbBXiUNsZBVWRIfM4IXkSmrOV040+r5KtwyqdxuHfLH1+BXIkF2XIrBSJAN7n
2/x3iITVhztp95xApLGmEkQBtt71Y3J+H8g0Ky99Fy1iHxID14wJc8Xs0re0Ck3B
mRd+dj7/qwQpN5hcHjcwVZLRMk7glFiymokGEGOI7bEyYMKeiWFXyZNB3TU9iBop
/blH+n6XtqJhChM9pQlLLtkr/qSNxRFATeJRMUb1g0AHzW46zXlKnPLTDkza7wV4
pvIhx8qTYDt/UE+QgVFctBXe70agfKSDHTTTpsq7zhWfKTGoaiecRQp9AEj2eLqR
JxNWJA7GpTMosXznyKwqCiDLgHz3gE49jJtMM21Xm3VQF6++E+I/q8y7wyrVUJzg
yEIBVBLUlz5GjdqJTWC5ktovM96h6B2H5fdgyyLh16nZ3rogD3N2qW8IMBq1JgzV
x5q18fmWNk3GVaAJzn47R0uUEWZkuPUAMGWsQ/279ua2wZOH5aeWzi/kCEqbrvGr
fBhX6IG0o7EV2Xs+LRiQq0TOBdiObFMBfYffW4s5NYe48ELZVgb28F7PIlHTO9PH
MKOGgUTxAvtkwOAo8ZPBzmh2Ue/945Qp9zUtSPYRUDH1Icj1p5tgvgBcTfwVdspO
LTmGexgZfygDr1hiTVITGQmnMX6HJEdfUA+EUcgZh6o=
`protect END_PROTECTED
