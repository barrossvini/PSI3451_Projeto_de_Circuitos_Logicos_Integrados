`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkrtH/nTGQ48aYb76/+f5QUk6c/x7xJUv4+3fK9WM0xQ8Gv8BaNCqBCTvz2LRmPp
R6AdDCkww6IOaE3JXWZ4DfGKoWJObWUWpdsRf7s6X6rG9ymlVUxOTC1km0ohtOA9
cR2LYvoZbq8AnNBkiRlBDcyEThTeV5pkQ+WVSCTSrk8L4ssa3+zLoqvHwgN40P8l
I/TwpEDrHdFY4Rr7Z6WJmuAkNja579uGzKv2d8VT8NVI7w8Q3ES6yXF5/Pc7jIND
qnqY7+zZrJxEI2m+qQQVA+vmFC/lP7DiFlZiIu+qWByc7BBk8ks5Id24xWUtyc6u
KGGkfr6bprOV6r6k5GXtxX6ZXzdt97UrGZ0hqCfB/U9RMPpKa/+UjJfVjvxcwpsu
dsE0+Lw+cuMBpEH3PIBZiokHPfhu0YPC5LSekVaLvcw3mQNv8ajpYP5afoLPw/T8
bDG2FrAr1pip8R3sV2ey2wnLePW1SDMkoDk5gHplYza/mlU7YxMcyBpypK3p5Gxq
uIcT76ljKydjklNsELDSIQK/L8hNBpWzacuHnVGrlvZXCz5ye99V/UCQ9+hDuDhP
a79IVQtYCNBLM7KDcZWmIK/ch+O16Ps8CQzbzXL2y0zMAVezGVvk6qgAu30Sq6a2
Z3kP/AAGWCCJf1ZCoTEd1v881B3QZr+AIlaQwWA1/HNRBFyc+KVDzKehw6jypMRD
7DQm1Cjf7gokm1Wz44ZilrZYb0GVXgkUzS9nfxuae//Pmly3vi8QO0Xm7JhXd0vW
aLXVbGtQtweeB7do1EmiR3wPvJ/Dddwbg+jwYObY+JOr/T4Y10r9b/OGYNZ5KgOF
b9i6VwgY+upIZUsn9XLCcJUHNNpfkyqo7tmbamA5nK7q0ab3KYhWBy2J6MO3LQGQ
2rhetTxmCf7Orl2CPT+GEa2JTJIohJpf5ST/wmDFlXmNVqsAJnAYwk8eG8oXat9x
4Ae6bqf+adfFfW75g7LxZqQm+QU47FacuQX+JSehEEg8H+xJ4Yuht7xuny+tdcP+
+kcMn2GlCDgxzV3E0XPH2x/kKK68sW3ZBoxyRMbDhlLNyLsugFaeFOkCvq+YfTaU
xJYs2YkDChjiXymAaX2i0h8i4+3SDAptEnpH7G/3+8Y0TUNDRBApzjm2vfduL2ZO
bbu45vkRB4NUDurTAh34PG6c/fXJUtqhI18CA1CwK7l9C1fxJL1FuvFEuCkAYze+
THC+McIj5Y3SUEwG/bVJ7ULScmtRYfdlX+xm3MYY6CKXB25kG8skrTlp9co8MZq/
St3cf1EgSI5S4WLz32osWQoE87UbofVkbbxtEiP3ufU7SOqRK7Bn3yy3TK/4yFxS
EOLpDNGeob3ScynlJjwT+HNVh0oR723y2QldBi348DvjakSfAk8cKvhAqnOmatMp
IxMuul0zMsJQ6Omgpe6qUhpZ32RSEHhLPhQDo1/4Fip+sj23UfECeVsb46Qsg/uA
BWJNFD0r4fT/y6IEcVYw9CtEG3O0HlSWHdrQmc4sGJ+ZfP5p4X1eTxBIEuSltE4g
JuDknqraq6WUwFhsKVEdiIrABmPyuC+ZtzM1NwDMivjAGCzodG9Ayy+BpoXjYwB0
JCzlevbdEFab8Z7ZCuLxXrunA5I01lHMW0e7tpI93k+6vyp7p7GtBwmhfqDR7nL0
jSRO2mc0QXkX3loE5vx/Ffbdp8Imv8bEfLiSaug2TlDFBajHXBEn6KkI11mV6Aaj
Ob4xzbFvCZn8IGzZgndeNFVLos7cYuRDAaFNIvjoo4FpZaWguUcCp79KfYYhKpER
IbHC31/QqGZY38cclI1KJcTc+Zw19jbFZmXgIO7zSOsjj5izbMLkhM+RomaH90s1
ZO5eQF2x5B6cYZ5wzB7vejDwL3VYX4oiBAmCOq69o5yfds3ObsXhuXuF/59hPfG7
ja3mKAs9yX+fjy3LfXkSdFDV1DUMVzAcSqVvHx96S2d2nZow7IaNKxK3PUhiT9im
4p005L4yjBaRYH7WNnrrXSPvlMGCylpspW5G95v4sMlYHTg5wlje3+69SkOonhC2
iJlK5GDcAl6ZRwNiRgDWrx8oo7ICe8qM4DSVvZ5L5xryOuZBYeTzHVBFmJ+kvLEq
BARsHm/qgWVQL2BFbnvjRiQV0I2ZWHRApULmQv+fFU/ATy+EX7WAKx+StYVsN+7d
WqywUx+P4Fu523sspdxPjEeeBN6xMSclQGn9oXyG/Gx4SYjDvfBNppuBJcZPCXDJ
mx65Ljrbgr7BEI8iJ1aUhh78IL646zmoN0xxFM5PMq6MFIItvAEQbvEjnYH5BPax
OZMpB9pIZHeR6NjzbUShXoRMSKEiAYbsWP+s550gazJB6fDPpQaY++MevPleb8uS
u8gCAmd13iW1Is5NIDzIKMvmzQNiYHigz3W4Dj2WLBlmPqGwG9OkdPedFMiUfyM/
APfhSsj1UVq1SfUT1SLShLgIwqjBm4XBkywJH3DJuADiC6DJ46MAekLCpCDmQ/gz
WM8Y9Buoeof7+Yi9D6PQQzYRPm2BJVC7+TlWzO02sL0EdBRboFYhlk8B8YlLIxes
csI8SXHsKBbldd7UAFfJm2SdakE42wzwoDFzw+H2nwsdkMXRv7jcwgfr64PBxfB1
dL60EX3YtNKUC7rdwqG3yXCEodtmlKPhVGJAk0m1pTzQJWJaDeVHXNye0hBcMz3r
T5dyS6j4VRrdPMp5fkpadgKPyNTo+Wi965QM5anJAz+jN5V8gXgwP9nt+WY01ALU
nZ9IgujgUkPS90M+8VGI6ZVbA1bH0WxWhFaTtz7XAXkH7K7zSaRspAOv90F8ymnK
ZTNOwS/kIOwJ/IFy6oN2ZUhC3srg1pZVie9RTXAXxEl9dMLsp+yi7a51GR6/ebMh
Afioaz/eb7AuxYZyHdWr2U2ytnBPwLDXis3POk13U7tQWyU64Uzsdo3wiyUPF98Q
MAJttixRq7+Og4386tDmx/2OoyBvORobPpWjyUhLjbfD2jQCZQ95Szo/Z5HP3Kpy
YREqf0Nx7b06AmJGXTbb9UdBopO7gn3Z9zPTUhkWGD20ESVQVsf7sygsxm/iOdKL
2kV+0ABoeGJk01BI6oIV4D804oIxHQnfu6a5h5BKfJAezD1FMYIy474wYAkSI1/R
PI/O6AezcK8pNpB2JTZEBVMNkMowLLTnD1DzpgRtCabM6ut1z6oW39KiUltFmUF+
1aQ25TIoOcwTmENMhZIvJK9AK7UIuJdH8A5i+A8Tuo9lAHGh1l8ntCrzdj/KksM5
lKi9K5Q8B0gnz0MXDqqkCvONW7NbmPpjHThq6RBaf/w7gohB1t5bGCssoA9eHCg4
Tqh2KzonROWEinYvcCACdJH6WJjdtJ6Tdc2mE+Qx/Q2p+4EsD3II91IWgElY8UKd
btVXfkj5vfVXzMt417DQHQFkFFG96VbdS91WImyDlHZBumTMkDiDKO8grk8ermtZ
ht95PftMfp6LBclyqwnRMwfLOFHa/Zxeg0gI2R38OmwVfmVDOLM3dHo1ufal31hL
dLbskt18BwFcZ7+APRFFahSDgl8tseHoYJGWKLS7lYDM0GiVjOS1ZxVoct4toQ6r
WARqMb7ftRPI+m3udvmRCdZ+cbS2kXpmp0xZbmxYwH08L4k41wpGo1GCA+m7zOcA
Qq8+nlVtbxPaun0xgPH/9ZxBmBEbHW4CodtqFNFSAfKoO+yph/LDiH0OCAYAhbI5
VpwTl2iLoYfRgoIMFpCXQHks8FRirx0KHSope7J3uVAaS8uz0onjlqjVOq0F7dnC
d5M30IxsBAUpCBs2SxSYeWQ8L0EH6fFx4gW0C54B1MqWZbvVTzG0vZSGIOJNy0za
JHfqdL7rhiMogw/djqMLts7p7vrcc9zSHzHdnBpIrzE9VzQ/k2O6bekpzBPiZ5Nm
f/QOPoP0hwYJhiUDTLZMJ1rC2Ilj73iw/ZxIzbdBMIEKaLhp/x+UcPmlPle8AYVY
sQQyF5ibXOazPTLNJCzc22idMtL3wfkhDXRmoY34ork2acDANT8m5RSE43g3HBtv
9IsgHC889vSlxH7bwjNjK3yapmxfpRAwr/0qBUQlk2LQJNA70Jl2iPTUHVmlm8Df
DCGO8arBFKYTwpNe6/ou2tNYPcdG8Vm61iaiX24FCBdy5FiPWNFQvVTB/FW51Bkv
pXgekV7xA1z/ljmk6ZhqWUeTJXnH3HDWVCDzN+41bqGdBHlghH6rOBXXSMU3y3gb
7xdYdLEENC9i/NqpGO4SvcwYAuPBk5yYkVZ03EE3qcoNUsPD1MJzknGMhVutTtQC
VTqhua5r9UP5w03vlouKia4sijDzm6TtoWql4RChpbc/P4A+i9F88NFds0raDfAX
yCQCr2tyDuj7mICKgn4YKpEPl5FITkVglnk4/fmzY0sqzMbRKVs5OfcUxkfbcSUU
oIkt8MYw3g2+s8PjB5vXpfW/O4DvRbllh6JO7GAIm4HWEZDfTXKps1AKLtHX2iLu
/cAWz4PdHT8fFTNkNF9xQuCYhmJddabvvDSv8ooHB7c0OIWFqmECV9xftFRC80ZQ
ZYT9Z72EBxpjQCnuNbZJxV+6Kr2hWuVifCsf9j4iXDzZlo8rhMST0t+dF5+rfAIo
`protect END_PROTECTED
