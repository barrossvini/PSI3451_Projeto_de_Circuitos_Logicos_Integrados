`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t/Mpa/B69nnrLLgVPRUtwtYfW9DnuAMwyklwTGjUfK/SW3mNOTn9AKDKmmtt6Tbn
wyKUgcplnLJP9T8fUQ+rtFQK7WbuuVNgSFNCw4hbFGp3ah05RCEblPJkUnIJvlIm
ESveJarPhB4NqcVcKp3Md+XyKeMSj7SBRP3lRLxYw/k+odNiC/vDp8ThJUbtt0lv
ZnuCep3ZXihaRXNYPkx2m8S7UDOfX1jsemHcK6SNCCOwoEGbS0TaO6DRZCK6cSPt
S/4Lb7BGcIVZKpWwYQ4o94NXdCsJZrAlH4ni6pBlk02P9MqIBTx5pKETln3ZoOp9
2T5ebXS8S5+7g3LKZ+aWfXKVYRtSNVE6nfz5VlUCNagt5jp3wtvCU7HelyutmWwp
r+L3Wt72As2bHSTcFBTtXuda1En5PHq0olePMiggY+yL5qikW43pqVsgtq2U7jKi
ggXCu2+Kew3k5TXz+bKYI7U4Vz6T8GOHlGpAgIzhTJuTqz021LNcA/NF4S0I0i8s
ZpuCbTIdUQVkRWA3eq7Of95KEesEbjmIqMTIfMtMXDCu8CdzO/m4Qe/7QBMxl05S
MXAFd6HyM9f5lTeiYeZO0oCxjjU7mh9RXKtPLnveq4gzlps9EdXvC3eOyAy275dd
AmNIdKeT+jy2XcQb5CMIXBpix+PUgc/uoolm6ksDHZtMZyPolFFWap/sJY5X7+PG
`protect END_PROTECTED
