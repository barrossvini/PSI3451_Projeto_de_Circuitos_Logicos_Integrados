`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+/yJcs9sjqTbC/mie7m6UMEzet0gmLFUfnB2KKXIhfru/IyjgcAMfXeOEw0AqcS
6is3L5jF6iag3uY7u6YoV/4tqlDRIbA9XzVHusNrlmA5VVw4Mw20CImHPqtFiBxE
iHmbRWhifqFd8tPDdR90ClWtKoRemU3j15rJACU/igmvCYlUiDtzih2WtLsEeCNO
02Hi8Ljd3YDP3A+/fBuRXBgswc2zZV70RWYPrLYFsll48u/qCAqpQ9pO9soXrW98
fELS6+lLjSuVuw5ICphmhHK9DZmZMZjQMh5XQQ+KV72yw05ANETWrwVGX11PpuPD
ZAzpLGgToU1JNImp1DdiYsUNbaOPHBx3QgQW5HSpRtCx8lkBDqv2Qbsm3Br3nkpq
J4HByyYMuHSd9FFdRKCq/Tp4w6KS43ZfkGjzrpoJKmirkJkELm6kUorkspA5Zc9/
dd3+Xk3VXOev/AtupR6WLtE5qvQHpXNARARuqOUBP8bp7pqX+Z7+iT1+YdRboDg3
R45QXi08SdtNN6bZPvRlG+FlUUOCrBkrAHnSf+6Gj3c2ZfYhJM+rbI+4VT5wBhi3
Wq4JZop8gls1Zcf8CSE0xTJahtVVp75G6xRFYvzArcmCNypGqoRk1Hd0byxOOsYw
ZHnMSFpGVgkn4XndRPZIVG/ylWWXjQtmgZVj/Jbl/PuoWNX1AQbCEMnIN41vRmk/
sR9F3RVOHjsvNFny4FDhTZaGQ71KK8ZNIx5OyjbmYmjrSOfW5Ph2kMPfavvdM57R
0YsegawPkIeaM3oTdkrE6Pyo20jaH5Cwa99HAFFMZ9VqqstqWc+n/kktdmJKTU5y
tKsuKULBROBiUCDOj0cw/Yi13cSDqhJrAB6iQAIbJwrSNML0/4lWatlnIKfLmgY1
vDiFmEo9hb9/ccyPKvj1UVslCm3qnyVaSwps3vKeeADYAdBFyRSVdMTBdtdONd3p
oUy8kuE+8/c2JmUOyIHSGSweuc94iHeCWbSQE0bRMKe+mEsUoApSq8jn2AN9y5+R
SPwfQnGry9BWAOzjtBhjBmjJ1pY/jwgR4fW2vME3VygR6IV+auGPxYD97gbsHmgc
iNIov7joD94TfUPW/q3/60fpTi30ULoeorNZxLV56Xq74DYauWlkGzWbmcz5R2X3
PVU/qtclybOekWlEbDaNbZjZO4iMg1GpJFuZhb5Pd7tWXEC5U53IgjgVLubwDxms
O0eGa0dw4+ppdvWlDUcF9w92S3qWNcoTnH0XrPe73tdwNx0G7uGNTJDmoAexADAz
6bBycd324k8qzgaofmsVqiKCbcWfqBwuS4tKIgzm/evEQAbcfB2RGnA6u3mw4qvi
vMD19KskGykGH0aFxNXQg4YaOWkwabQU2Ax3LKik90r3CB4BQntasWtXA27u3yeS
GCTubQ+vvB1NXtex2nnGXFjYIBsDA8YLQ76jKJbkT/8FlEoPkvsDhxjTHUWkQ64n
fDuelxqIdNXq0aCgzhhHjSVw+fnaoE3RRvIykmVVVrEdZ5qkSFWrxw5lK0DMQ5KI
Gjb/BpweTkGNOTg7Nt0mQtnQP0yMIUetj1hxWJYE+HmNweUVGJz/lFfzQayXVzWX
r332kdZ3+PwI+zR1dx65JF8+wG059z3lYIZhondW1eKC0SV98RHFTkCt4hmhUPNh
XhjhOpBLQW0TngdxC15vXhj2s+V3Cit5uiU5fSV56vrnKYycX4v4C3I8vCXoR5Ht
w+O8W6Xp8RM4EZmMG7MECF8Q/KwzmP6JFpXF02qkM9+NOiKqmibtCIlPo4kjdHWv
FQnxDgiYaaI4KHBfVINc3RPQf+GMulHVJjkzInMMhHKWa7q0VgAGYboU3ChIVaoZ
zRnqiwucswDmwJE+8ZejYIdyat9t0SbcqGKoUKEPimW2UPIMLh7qJ6UNrNEPie3W
3XiG3oHU1jNfsra/SAiptU+YL3tJRtH76FaDw+16tfFs2sBRb40z0NzzEsuS5ser
i8XFELWMQ54764jyqQNxwzZB/t8i4IdAUSd4Hw8goLM8zrFpGF7UOHZNmCZWzT/y
xpaui988CuWGqi6LOGtsKLoIIs6Do04qrkNxxFK2O+BoHqJTPwe0nezBP3wq5oP4
A5rt5/3gI3/qgVu8mRlLFzsRTYmn0lCRZ253JddKjiflblQPobML/W2SAx9ypYaR
P0vXjUgYEE3D4/xKJKLqYuy1tW65LjfWwHIZF1FA2XiXE/mSOeLbXfNk6OJ82tfO
zUbreQJSbnojigOKaBTHyJBMTI/CxXwCfOJryzwoMmdgpx2wX3uSEp+pcaZsSLIN
BbDWJensFpqdjwziymyMrW47valzxpa+mKs4AcLEiSyGBDA0aPloU6hrv8scsKPt
TEm3WG4rCLoCl+GY87j38jhkS3LlWbpwrHPgpqtkKq3iNGynz9jXiOmEF5oVpUwA
hE0ponpWv7cZo+6QaUdQR0Tx1gWRNQTeP7f+rw8bHnSsZRiKLao2qlqqdKN5ODeG
/K7yPBEcWsj6QCvNCKR9vWHj7WTcrb6FgSIzPYKOAPvYS78L5lTJ5W8u9MlZ4H3O
1LMFItVw9qSwlTMuh63kbD0GVNZIIw6h8mg39M+HW2q13j95eLcRH8pIO5LgHCRz
CBymACzb/o1yEVtCNu2ORcoetPOiAywgeUmzACTBa025T4UE40GbHj7j7bmxlmDp
xnqBNhI4j/8lL9CxqyMoMfsy4S4WVe7DowR0FQBnYDmY95lTlplYAqS1wAJ2lsW/
HcIhbG4ZXU4n+nVZMXJ5bA==
`protect END_PROTECTED
