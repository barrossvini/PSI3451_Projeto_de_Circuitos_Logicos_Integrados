`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+4wrgDJUQSJ1sgNkAZBv5k32tFJFAu8f1s45YQppPKQ+BfJP1SzLcwEda0DivmKc
1ZvS6tJpTuLzozCR3T6TGGvTMnUQP/GaVMkVyYD8NM3ft3LDCCl4ZrHOeVn5nxdg
6rvwL92kxo3jKivcQK91grpmUMFoU9lqw+johogf3Z1Rl5qXByLpLEvjxvZaK69W
ls0IOM5cZOI8FA33qqtajPLQvo6lPGm2U+o3m2z/BbyAgw+T7QhfgLhfstVe5H6A
/eumG++SG5oi6YgmA1gfF1rcHg8UKlf6ZAF0shAqGr9zyGoriqk3kuXEo4NNdqzm
dE9wNwZZkyuDaTQhwDRk/Q4DSoLjVc18pMlTZzz49YQrGWy/4lxb3xDU+6K6VVFB
Frrleerkuq7nn41l/sXZJVl7xoQsj92kE2+bdI3JaSni0FkwnbasMnielXGJZvzJ
9i3RpoCIjRVdeBYDdEFZZxIqQJqE9/+gnakiJXBgcnpf6x1l76ssENRiT4L6DcE7
6oDhoLKN4Dd+U9iYN5GarkdaPTQP4QdmAiiy3GG8Ut4hXFFMRaE+tmb/6LX9HWXy
aR0VnxpKFNd/Z/l+xt36jSyd8Wk+nioqUQTp07VkYRofCKHG6vXhLJsjR5Cuj5oI
wvjkehZhWXofZzU3F8z4UNRKBX+m5CrQnRk2ikNYeg0bOk0ybCoN452QgdbtDuHL
qhlwR8EyzETxjloWaP1XUCO7I0j+YCUMwKVUkT+w+a5963HXYuk9jS/OiaQ/maWs
SST9U4WES4RKFX74cmgvVVTne/GMh3oyqnQVRO61dJ9FYoD4Np2sIHSo0YZkFxiT
2Vu2THm/+CDhD5jQdpI0QkEWZM+NA5/hL6d7LwfXClL0OawSvqwkqdbhtcNYZdX+
7uhDd2OiyyLE5mTEUU2QvuUsFnTbQ+VAndaP/hqnRcs7RS9wHQFi6oY1i7qJbd/w
qMXwkylSK0Uc9Z3RaJore5KWD/EyaSIR50zcmadHxdz2L/kSIfSXNX65QXbixOPG
IggM4nkfgnNZsDpKasBLrMCugHadddtHBb0hSOaF8QbH8AKN6FttUW9l41C7cENK
x7xCoY32SvBupBa2yjZnUDUGjSWHysnzF+nLstfZqXSBnlkF4hshkRm9FAhPyIkU
Ok1hGWflaOZwPbOz4iM7UdNGgmKyZti0kDYyOWJc/CxBLtuKCnwwRlVhiABTMR4T
j64+0L6HjbttbkVNbT53ibA3t0kWsP9w61M1O4acXvpKCS8y+l37cewrOQzSThIJ
PHDP9RyCExlujDtrkl1yUC/atBww0G0aPM0WlWJCQ2j3TdiJyWm7R69UQbNdFDza
aNrBJcNlwCbfALI5iHSqwKUr0BuuTpFARvO0sc9UsfF1toveKOveevyZJHSQeLiu
sVvlHF0KjsFKamI1AaxBedkRc87es+8M/qD4qHBTXW/A3A5gthNGfMaJjJ98vWxO
rM4CuVa2lQVTmcPJkXzTKi9QwP8MnJ/MxInF0q+5U8edeoQpSVgRmhHF1hqrq3lf
eog65YaYMLUgr+F27PI/Dp05v1iGL7CXYRKarHSyuYhK5rs8saDf7U9aWbPmImIc
TbixUVxYwFht/CfoOJIVqYm79vMcJUvHHhpi2k79H9rmVcfy8dq7BmXozGslRCdt
U2zH5zFr/W5DIJyIaZPyUBXND8JLjP1spGL+AmSKqsCdbK409yLhx0R2WzM/tfPa
0ytDeMGCSBjzKFznNyIR/9Vid2ttIrKrz8Sw3tAAnQWE3csOb9+9tA629u97uE5y
aJiILwODjSTuWuj8AnmO3hc1po1FWADNup0Br0Ixl7Ril+gZNtP+rLFym7IajL7r
g+2Xp1D4S7woZF5PS1/PCRjDLzDFC58IeF+GGxsrPtyQtAQbxaA+Q88O7N8w5UsY
hQNzWa/NNm1T+MURql1amHnsCd2z1zW7UXrhllHv35pY4glOMc4IYk1Rk2fWv6Yu
gdQBYotjoWVf+/D+BvBlmoZKCSg4XApTA+aWLnrJLGKPgAy8CKttoq8sl7HU3Ek5
I4mwgnZKVTLDmsziFmfwvnjGx269t4dAo4B6tn+5o67VFJoLC5soyOAs4YbbLyAo
VCWg3cgMBu2AwxrAuBvSWUSTKUTKYBUspl0Q9AjOESyTetea20HE493geijDGurY
DUL8yd8eXhkYyfm2/bj4wAjEEV3g0VYMFW1Y/4EJ6Yd4/N9rxbIdXJRgEdbeHR4p
PnfEkspso6mlEEJrz08xlpdVY771S7uTXAh2zI7pDa2ajiie8uLJHJCzekogfJEa
Lik9yBN1AVflXVjqByV1bUNGL+0v6DRVbvzNUszWqRFA5VcJ+dj5fmrQraKj0eKY
T2cblq7v+rZGuCd+I61g6A==
`protect END_PROTECTED
