`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vsfrMGfTTAuWW88lxxQudgkwTPdFmExKZsEyZ7xsezMaGtZUPQPNINuU5ZzA+lSw
VKPvbDTJWaPEY05UrgYvQ2jaSqRowVGlnoMbFYPkUmPUu2LL/POt49WvWrTdwGgQ
v1ee5tBhVw3ROho7/HMF4df7DT89p1/d3eKCPYRMelxOv7PB//fbwG/XrnyudHcO
+cEM2ZtDF+m2ZJHcMccdvutchiw5LmKT9EpXSRnpOZuxrUaAT1tG9bdcPZZqYzxH
39+WSudx7e3PPe736LcUkdGpryg5lh4TLvPGlm0IwXhViGkdAwVD+ErdMW8DC8Y8
+F82qqwOHdWUDor9OL7oY9xy9tKGnsq+Veymq9RhWcJ3dsgCTXUiOckr5TSJPpnc
QQvNtc6BDbX8lUgOUxpRUJqfaF8OFwoPcufFR6w0qIzx97Njr04IQSazPnegCw8k
V/Pj6cow/Wqmxq8O5osEFtrJuZhi0OFLPvYDK1NtrNI+yY36alOweoFWzghactIl
jKDyRUQoSVcEqgiawttLBnNK+2pdg3pgaQpma4cUzYLYvEQAPaD/gTjwjA5ayhXa
0hspsWrCuN0T22OVINEMdFULab5oYipr9OGJNK4vngY1QY3abYA8Ee7Vmu9Zr3eq
LOhH5K/VnBCu+K70dlbXVEjZOnpVIzEzCWCrIbIXqZoj0/Nz6BtXfNuHaxQ/uySE
gLMgZvN+pNCNQ2aOuCK2UD8hkgDQGV0nedC8qvrqWvcMFP4b/93cF5ijfahWWZgu
3OgT64y6MBI2phJ8nqWT4Y8CSRq5jmxR0nIlppytHVGx0ZmdixP+IqfsWLwktqbE
IzRkdCVW162V3G/8xcJY/NIfnVZNe9Y2+Kh6sxRpz3grSjl6RXGHRAaKRpt2vTVN
MCB+SZIr6fY+mips3g/SryJa++WI9t8NzKM2ncfj3KQ=
`protect END_PROTECTED
