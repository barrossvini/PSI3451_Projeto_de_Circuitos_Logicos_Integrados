`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l2gDQhlI3ucbw5NpG2euPDgTZ/B1KRSsrOPoS50W683+NYymiX+tHLgKL2b/5Yjb
ezTsHuH+y/hBvbeV0CLxVBlLdxWxHgMFg26eRlxETCpgnmBMw6aBouBWXbyQOzZ0
5SGVKovxuSsC4zvBa7We79Nlv1coML/ZwrVBX0+IG7l0XpPR2vxr5hqrAF2sms5L
hrjjpELX/r707Gau/e370i6OIjVVAi9tT9QZfYY4GOQuPjaO88lGlBxEdpwpdYBP
2uQScC2zBH45RTh8DDZnW8ZXpiFKSOiOil0jHb/pDedk2uqSaMxx8Y5b2krdcWP5
gX1C+pRT9PBIJw05vTNLx3mqG9LhH60qwBs2NwER/QdOgVB3PpINwAPB22dxATor
RsVXpe+PkOpgFPcdSQrQAvgNSWC//2UwjWygALkPqmfLGL7OaAwQ9XbT0w+zI3MJ
jG4l5IvDkVNyRPtzN2jhFjt1QuIOObi3+VZ+2lpvHtOxKMHe2D2iLPe9jcgKa8Mm
ZjHuFXOS6Zt1/5PRluCXjTLPiyisTd9gWhlKspzKeIx22VUgaLy/fUHgjWHarzlR
dbnrNiw3pvVRskyV7tkojec5uq1gRNoVUW4VAeJDVWosY96AEFguG7ESVu9dG3K6
/zgJJIwDEarshXSkOAyGhIY6tFCBerwywM/PvuoNZz1s/H4QH67d/fWnzegLeWZ3
DOTjPkq1/bRvWfchPwhN6woVqoZ2Cm4c33p/Il6rFyfY5uLJa8DBWILyAM3b3o5p
xD7Vm2CkYMO3SHvXKcnmJ7G1RfIyZ9O/SmqoFyE3K2vZramGa477g7LBwj7PV/pI
iuo+ZBPHFR1qjY/pl1yjsSiIyK5X91JkwVj+GHZlpy+vjHtO07yPz3y3nkSVESvn
YdNhlgPw9WMKEMgaUmfkadePs903luGf8xNj9sSHGOlXWAUSn8CSAnfs9HvOZUhm
0MxbtslDgjoetrF1nyKUxIm0yQa5/9MQjUgITA8JSH1KW3WK9VOol7i6LzkIUISK
QiajGo32t+ro5a4IaWzJ/s0cDlHEu7PJ5GAIp30YeTcHDSofB6VW/F3HYuwCulbh
qlHfptsONXsPWqB2IL5LtQRC2wlwE3efrCtYrfbBepWVLRDMFDkMCCkzayYmn9is
`protect END_PROTECTED
