`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Pq/x3Pmbz6D2l94YbmIa9Na30b36vIQbO32PdkWM4g8CLNXK6LEQq3dtm4veY9U
uKMPi2M7S4JbhtOoLBWYkPEtptWpxJzxZMiVMHiSNODdMpif7FoVnNIiUd1LF0g+
ER0dBKzTgrid1VCIB+HX0MnkB1wZkwu9LutC2p4fTNWn9qKmMrpZyEjDrJu8/ITN
I5EwfKJsRVUivGrodNVlXBawtWQ+VR2PtsvjI9QbA1nlRelFHhy+6iybI+9AxpGU
K1X0+HGLxpt/RaS61+x9T/4s/+TgX/T8oHJOJ4x1nbcEIbAqOZgsRbyCEx8YBWgm
CqylxOK6akyuelF89wNR4QEscB1cl8yPa8hBpfUGqmPMK+Mc2tvozp8sQV4Kjffm
LuEZ4byV6vfRH94R67Civq2ZEyXQLPHyLREA2wUSxopyyGnULz4HYkhglmnFSnoB
K2LZq+rHXZTrSc3PgZNdcRhDWu6qN4BymV+YY1ed87IbmXjaWp6VToW7Ktf/gnfT
kIoWpNKd5NsiAqZZbPeoHzjBG3p4bGVXNw0KUGcs4rE6RdAlYV1z8rvNPKusSGZn
WwFJLXnNSrP904iarKIBDwvsWk6Qeox003AvPbztO0iNyu/Td1rLypqTa9QPpRH3
SEekXbimG/dAyz26Ia+Kpv6LSGheNiDjB3jRIMuYWjx5UWBjBFex58s5RzKbWfH0
+k+o9+N9/wmzLvdomM+jdng1mUk+/s5By0ZZIzbRYWS+wshjnY7vZOZOjtiqxaqL
o/3D/3Wd+K4tVw5N4B8ZOF0Py5Iq06pcnROQV2b2EyMPYEaPe9WdYKFfCCkAL+ve
Tbydn6P5vlU+aNkKLCpmQ/cgUIYBUVeDUvOJePo+LCBnzxc92Xv2WgsNGmuOZS0D
v/hIERkdJlrUcClrbZxdK0fr+yVKnlM1tF5IPab+Y+xC/W/GEdj2LWPz/8jeWzmq
9L4KVNELsz7vtCvs1Y9/QXbzrPYNV+nVZMGtjXxU5aIABetkfEE++7594QXGF03p
akAmBUJz7/a2SFIBWWVKnEiGmK1kA8tHbHI4/GOqUoNYDmACJGFK0XkHsk9NDkXu
HZyhH//iItd835fcPw/aUhsu4lrI5EUGNpn7rrj22opUX3qYAr9qNCfZvYeA7fqz
ZyAgvuQ0FelmPcnjR8Ib1h+xeB3/i+Kct44qDEj62tvdx4LOx4WG9zrbv+Wih+2A
vokB3bGAURQCHHs1TLXOeZE1RY5MPecjhxHRbgWdQ8PvGlcWaxZUvrHvk9ks0Yw7
m19VrG27HzWUv2xRtN/xfpwbuLs48vHv9i9B9j+FDaPc3qyjW/l2SMvtpMB48An9
/JpDv0EK32aVkO6EGJhBB5R+2bGA5eYECt3kG/eXs4XjV99L+djtbt1jh0akAFos
rc/m58avOKUNpzzJv06J2h9E3wuamkC95PKt4M2Hcn1oc6u+Ncug4EJ8W2k+dPNf
p793w3dJGrvmG/JXKPnbi+g+CRTh7Zziq7Br0SEWzJwbzSvoJ+kcMY+b6OCXUbHF
RA0CeBCqlFNrvZXZmp1P6Y9NYg8hUFVxbqTk6r5rSfp3qnQ1XINKUPGB4rGH94y+
JsYFc5QLoACX5MSPSmycT7lTZXWsCFQELtxMYKxe6n/9l5ERPJi7fd+uoDnq6b6c
+WWpJlazXk/EXpOWVugMWaqGzeCtjU/L19GMMEhntxHGT/ijJfvtR88U6DZlobTp
HFXUR6BakfOX2H5iWmDIntwBVVL9z6eIme5KP1ETmUR0nKwNq+5WC87G19MRJLlO
GwzuwAaifd//75elnkfzBnYHvfwExs8N8azcZQrywTWw41g/NDShPTiXW2uistTt
LFg8cRkvfC5kgV1aLsZPpQ0qQUbY7O9ntUr4xE+N6AZLp/2rVvVdxtXrLs65Fv76
I/CewdlIKPm4ZRThggbJAwk5wZzPFzOCOTXuVXz3VBX0vLW+9IDMHs1t1tgCgJal
zCmnow9OZI2SbVAa1l+e2wPkxX1AsVCoBlIlqzqs9tdwd/US3QzlGfuWY/h1r1jy
vCmN7zD+mhkfKVKLUWglT1ahRdtuCNGC2j3eGdAqbd6Xgp+oh+Nt5X3k6Ni9ksSm
faSmKk5kuJ2CZfxF+dW7hAKqF2wF58frYkoD+0rIK1NFAEyHoO1RZP82d2N/Xv51
vcSrvls+mW8gA01ZgFqUIc63gGZvh5qDnUZOywSnRWHT/kejEB5U9kCKMSB/Cw2V
tfDs5tjqxrSn8dp03FKdqZOu0nBlkpjUgYZK3NPQdfLu0crmASaR9HQCNA2nNci3
lZ5KFKFW50wel2ZrPdzZHlsSRRQUCo0Tlo5V9k0pIMkFd6Zd80pJYJI25lT7Ji6w
etQsal4bPqRBYKqQT/BLW01lsHZod9h56zVfPLmFxUl5H/zJx78695g+VE85gKqi
ibbIC++pH1L4PWcHOk0g0iJngOwf3fKFjZOSO4BhtkpaxcH9y0PhAEDGbR0P+5Mz
gQ0Z/B8rUubOcZY5ITSFCKmKFKn3HHbyVmyBWS0nabQbC+WgU5XA/H/KueZjwFb9
q73BN80qCCbfNnO0d1GfjMFPumHSdaB4X8Eej6hH1SYxQLqwDDZigNcmb7MDfWty
ElUPOX7CtrjCZVDjsRSelYmvqAu3o4xZVYVAwCgqF/JaDJEuqwu54zfHckLbeki0
JlpcTEfGDYNrT6UqEBlZ7VCZHlC82yGZVKxEBsV9O3JgAJuM1brlnx4FOu5ymTJJ
kJZVZ/iScN1psfWcpDKdst+ny8QRSGylN0mtEsjlgy3kwcieaaHaKqK7/HP0K9FL
PD8DPQs/7gbm98Se09AVPQIJ1DORB0MvlZfZcMiaizecdNfFjs8KPd7R+5oOQTbL
t0Pyg10iD1VS9DOduDZmwrzsVFRriWquBMnXqhGCS3aCypNHqzswZ2rPpZ9MXO7n
lanpGr7rOy6dvpIT9HKThw3jyQYg8Yw0fdrbzv/qXF6kGU312Ujh9HyIqEaZFSul
6QZg00+RB/4jyaffPZl1p9OeLAjP/ZJGiGv/Au07fCJ9/n7G5V6bb8kIpFwbk+cn
D9W1sY6laMp6uGkZVk6t9DDVmXA4OW7W4qaq+TX7HSYti8fQFdGk0f1ZZfrZChGF
TvjHMzwbg3B2Ar2ZWh8SQeW2BvyhOmSk/c2y+OVjEKHLpeS1HQ+cHV6J1f/9LMBW
Ua5XiHGKlMNrtZ9AnlL5BJpVxLUJBF+m+38CMau0QijJHNFl+ZI8/NGIqn5DzuGO
kJdR919Jaf08QJPJMk82Ie+hc14W8Vg3Ojbqmn4HJ9ZLoukxo5yoSgT1XazMCuhN
I5ZEwVQ9QSdOLqD1ZJSerscWOF9d6mbSXp6f/LSG1Q1bxB0K6cP3h9fAco28BeXO
AbxJFkeOo/5XDHFlnCGCEuzf83iCQa9yN9CcrCPhS/7f8pAsYV4JLvoTqlJWfxyY
2u14PHbo3hjvs7XUgc5suwK9/gnlJO/OTtKMi6/4AuZvovphtFg0dOHt8r+4ub7r
JI+2hML7pRn6JpIvNx7dnhpbNhYxVyKuVD9gtSnQ/Bcu3Rd02H8DvMhoW37kQ9qn
UPjthfQnczmYOat/hj0vggXuez4pcpQrlJ+cnKeCrJkztWm4ns6oe7mD9Wwibzai
4VsZRt8c4LzQkUnHEehPyJam+CNGdS8St4AQrweqNY/XqD/B/qdiWIKirLGQBPJo
V/QAfnA44rhePscNDvGVlzwemRzKkDhRej/NxIWE9rde5+T1H6LCNfWRX737N8mN
RLSSIhv6PpBIvLg9HfF28YlU36BM2y6Y2SkorMPjT+5vgKoUghXnpvf++Ysi3QMq
QcHt2ozHKjZfgXxA2KAFTO2vBqoIYQyynTPV/tzvMmEOsk9hNo75xCqW5bhTawmN
xFEV8XezSjwORiRmlpBdLVor6OFSWZ/EvS0XZbWkbeHrHQFq/s0RPzdmBN9MtIx4
8xcD3tTkGiphRbtytjVNNBWl6ra3fzNGXHPpf81It8RHFrVf89MeiC8W1Pqa5szm
mULhHUUgacN3IUb/SAWd0B0OkYAhYlozqQv0/pnJl/med5+Ps5iXxO4zTG7hwAL1
TnJttbn0Jr0MYLjDyYTBuzP4WK1qW+KoHyviPPXw0lBQCaofBfF7mtNzowqP3Y6C
7yMx7VbeBeH/4KZAGVGdz6Mi2DFWxGz+J+kGMWtWwE/pW9pHfMjKNpEYFo0BLpAX
Z8vVG0QPhGYMEag8hCbhb1f4KdmAEIH7Ahd/7yBRwhKvIKO3v7RkzEOZ0UiyFEj/
6TfCw6SQgQfskH2J4iwfsCsCBFX9DtTF90PjjuHnoUrtkxLhGg3x6q5SBGrjc3wL
YV2TEG7Mlqqo+hksgov21guAgHDXj7TIPpUbHpihh9u8fhly8xpVEe9krm6gaR28
Ku0G+RUVSsGzAZ/zQoDqQdUircr6SQb/yZWUB7O96lQMfs6T2T3+2KNCz3FNTt2s
+66qJG/cdvzMMdA/75FxYDDkAlZYdhznXTsWv4sbtxNgM9WOpWU8kZ+ps0MmZ5G2
v10Gq+nuWpDIxz4HUpw/odMszERyn/C+0lxYNE2B2OFHhTPJuyxgDbXieIA4AH4/
68RivUOKjoSLXtiUd5BuMNdpRtN2ZSfRDLUDHMNar2VUdrh03coynJcz1OLTkA87
gAUpZGOOMtSb0g4BUKwEJl5Imrb/mWMMMbtSbIvW5wD+eFX19S2RHKEAKCFIaKz2
bn/9x3uv84HDAuJYO89LwDl2pdbGUg8JFR49YLlkJ1ZD7qZG4Qx2PBC588MXLOp/
K7IwrMvJzDOkEp3p8xyOycy53OpzKzIDY4aIQZD3+bkunXdZdQTjtAwkfJNbwld4
NTI7TJ+YGQDBIXT5TT1HL+jiOnnXqKXFttO2lreKXDrfMhclax/5RzzRXeuorFFu
2GZD4iiEY4Bt10YE2srzBOIRBLfMFL9h2BGSIyc0ygw=
`protect END_PROTECTED
