`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JIS+AOuSo8MUSVmtr3e/NZ3RBqL8dTbZfeOSjbhsTHHFgI4ZMS6rzLYSW22yZpiH
8qUc5mjGv6nBieLDJ37TAHXd/dWJVMEJ72v8HA+Iqn+OHcnNpfuo6St8qEM+SQeu
KdKOuSDhgmcRgF9D2a5UliEqHQB6CfCFVeauCuax9377q2uu7cyHjXfYj8o6QcH5
oO3J30/XalkoelHOq293Qo78ygUk48goxUESXJ0D3d1H6R3FV11g9YHqvpHOgq8g
FjZ3RBY7PGies1OjgJBn6R+fDS1nSI67Amojz/1L5vsHc4GmUkAqKhV+H0dYU7mE
r5MpG7etLMRPr36TjZREg/vH9KZ2YH6mHDBmM+siJnh7gzVaaTspMMF4ffydwTNn
hrRXnRnFNKNphsCsEEmkoAegh7lstZSygH3G8XFfLfXsasNNBWhvdyxKlVktQzGv
hVACdgePxINocOVY6r426L0ZaG5LWlK7XAoO+PmSBiKqOLdkaH+KPfWw/qlbabfb
+cSSJDtylNnupvqRvi8DuqCDtaklq99vd1QdHatilFEVVotAdamgbGUVAsEylv+T
kQB5fwZBS80+L74St+aXNN0DifrEo0rv2imATnFb5UNgAY2KW8IHWfAeSN0nksAA
p4Sf3D82VbkGAqVj0DpEeMBcpq1SC1rhhRj40WuPFCeF2SKM4KMOfE67JxVXQJsd
fAjPYt3Lv5tblNo8bCcyRcLztSUH0DJq+TG6FHQfNG21ACaAt4u2HlfA+5PiIcsk
CNbuFzp0Gyy8Eg6EFYDnR60eBpaAec5Q/qIRK15TXCzsuext2KkWwyn89WMq9dmz
hwmP6Vxajty02JrvSybVyyxkG9tbTiVzDHDg8oZHcgCIyDbOAu0gBbbDyaYqJHeT
Upi9Cnu9UST0R4gk85eo57VKnkTWKEnAHj/kBC9zJf9MfZn4wZaN4hamqfTyyXat
kaZ0ugDTFxsLuuGQBuI0R0DpYcRbnKoqeWiPn7cu69cMZFniysgeLUEb4V338hgF
lt9/f2XACx5EQYCT2N7C1iNB38AAIZ/b+kyZiXop9HYDBYy5aqPsEsxkyN/4gJTq
ReLDTwoBuldd9zUCacuQgyNLbpAIBKLT3tzcnXNiX0vBvsZ7yAkJOOQKUtH2HXMB
dEzL9o5fXagMtaAvcJP20ISb3iPPBS+FE+0WtQNfdOjaO9Zikat8uVcfp61h9Nsp
k0jXXc3X38bhnnUe0MIt65Wg3vA+m4jrm6dfJ+EyW/hCNTYYRF4ctzcfeZ5efZhq
gUwj45NQeiLK61xJ6K03L1vKjNiVjJrQllR7JwnjLoC7mBOq7m4ayImrl4fCyISG
UdLAKBEdrNbPIJHM7xegK3HAosgb1GBGNja22lWPeaN4yGA0Vyvp1iu9V1zE213L
zvfigIyaVn18VhWXiNBtoN8Pxrkwvpu8na/fbCtSF0yqpW8HSFIUZxQScG2dT4xB
S8JP1aiUHjtLGzWA2uJz7my4iNMld8NAFYn8v5mio+AfLG2Gd1eD/Dwws+Ng4wYL
VEtXBpJf7JLHmQVyBNOQO0Q0j24IBjL4YapVYstERQLS5AfuijjG63UdeF05T8Op
X0MCX5sS18X8wVg+YKjxh6DnZ8af4EaWs2uGTGdS35VVNKcogzt1SUX/bnhL65dF
1OvRl3CG5R+MTE9m5Nnw2IAHQQv+MZ7eZiidAk0+aO9mWq5VW4SVYuIpTSjEpKmj
3TAjLIH/EKt3V4un5YnwrvbmljIIFFa2Vy5GZs2aNCyzBuVrz59XBSU50i5iUSrC
H4Zla7F5LoaVzhM6/8BHcUxnF6ehAf5rpasBgYJmL5LbmHBNVj4h11BiFcayoDAy
cEMCa5CWJKp1zBv+Oj7WXP1C1Cws1dwhmht/qMeepb4VzOLLMXXrxKBaq1qdwIWN
pRDd60yua5Plxn3C2uGkwA==
`protect END_PROTECTED
