`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G/6wNngcsnwmY8vQo6cVg0mom2gk0UL5eOaO/mMlQru9dBOhNi8Kkbe8CSqfbnlX
Vh38/XhiwkKuBfS0PzywjPJglAyUWkEYIq/Aau9eC0jY6nuPhja5h750m2ID9xwK
/Cbe2QtZpA90WLko/s55CC6ju24nieCQC/lJaezUvdXLwIN5IB4Nt60o12RYDVc9
ACghUIpzsv6C2QDm/pfrq5914FwAcQyQpgGctr/q0/cyOZ5YkD3mnkPJDxhYT6Vz
AfBPMJ8gdF9zMgCztRMY+q8ySSDtHozYLmYcfTwdBqHntj+1NRiqFR/VpwlaVxXy
syVv3dXQBSxnT3YMg3RbMpVvoUvwNNmJklZlIuRFajnqy4Sn8rSE7toJ/c+VwE1R
FPlmsPa3hryrxBfDWAikblcXrEQYEYFNrZiSgOjQRzBhi5s6tq14gzYkFuTz0358
xoDYtwCkVw+smXCbq2pmyD7Kar7KbbL4qRBn6tFmokUKizUgSGJ7Eqbzr9zcwzTK
bQGhCkaFGlS4MIAbVxNMp2Ci1DxSerpBLre8NahTtDFl7AQf8Yv5u1V0s6UPb5zD
iW4NoVrRHDC2QXF+5rMhXM0xlZo1EiYhgkffzjnov0zYF1OVz5lSxPLTOy4Of+/P
HizaePK/yKngtHQzJQOgQuA0TDTmu3b/YzZ4RsE123rlbmymWjCPo+wDzxxG9S/s
0vWedr+EKSi6kAngw0k088t6sFY9EMAbyOeNeGAIFCAIr5YcaUkw94haU7f0nY40
RDvG5A3pMoyrdiAimMVWyho5wXEvwcpk57xJsUTh+zR2o9qMrW+RccVkNT0wvAnS
8am7sU6yw0GXv+a58jIJNr7DJIzTEM7j4i89H1UFXi8QWiB2bqGZ7vMhx3xe+6I5
en0d40t1EYmUFKHcrHzZdcn6wF6z4Rwe49BGmgTX6WBl7Srw885PS94GFWntABIH
+ZZTZiQHPZisRgZyb3Q69vYXh9VOwGPWenOwOT2YXbuW4ufzeelQUT5dc0/ZFGsM
MN8bKNW56PwS09NlgGZeqUAd+wRjBEzoKJVt86m8pAiblGxveqcrfzybH0RP8/6O
ueaMf0yhcGid5DZ71gHlfjCxpK1jRzxb7vOHCLUYowpYjsl1bC/e9Sue0GtHY69n
pX6NhzJs38wIJFVpeaniRztJJzxXDZLGod28AVWWKaB7iJJ7a9FF1ycktcmm5SI1
Nc+ycOhj8Nbpo/JZGnvP2GDSRthKpDSANwUPqCSbAGE=
`protect END_PROTECTED
