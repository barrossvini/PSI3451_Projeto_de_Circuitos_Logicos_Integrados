`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73s00NQjzIgI9+emhMeCaF23Rz6qpL6T7YsIpEdfutGUHEI7pt7U0iuSN79ywvln
LbVyckegLO3+4DO3pwN+ljow3OH5MM+7hjI2RmJApUTd8pVoVTjQ5gftPlc1eZ79
Z66bQ0UkPM1hGZoKw5RkPIFLm6s3vHNAEAVuOGXrRAfsJRK5TFpyiUYIKZp+Jj8t
AFhFayA/At+AWSq+PyLTytcm41i46emYmu8wOupELFS7CoFdyXj5+kuNmG+qfTDq
1XNRz/2E5KrMdJ5/7n/oG+qCAxHA5IWNi5r/eJ08gCSXBd5dl3mCmWlDwLlGXKI3
t1cYmBzeKTOixI47WPB8LbwwkGMYjfsvO7zVEZ5nq0ZlhhiYGyoRqk6WwTg3h0uh
tupLXK0oy9Il/HrUKYTfzIqiTPxweOzgNr/pHqYzGyXOpAxTlkHpM+B/ud5/bYAO
rEZ8fcg4Pq8cGZRLhezhhQsSIXbkhXwdO+uMO+8z9CIR+rUV7rgiIy7xMJ95Vzwv
33fwxT8CNW4U7v1Zbjsi/1fcZskEHxkC9Py3bwcSHH+zC1LDOEBnGNOpCsBDxazr
pMvpF22GcEuIRm4tvV2N3fru/4bRUqcBHhfRE6YluGLweIQdXMm7aihCpg6Rbk6+
+zaFZbFklWvM9TtZdKs8QiX1qT0mUL4EMUQpHdRMEiIhmJmPI2buQg0UNzBAEXCj
H+vcgmPY9EAlIsdql30em2yeDkajeJKwks13gdCYpPjganaszt53HwFPw/KRM6c8
E92Xdo4YJYUBPj3hCuZ6X/wa1mlYMOs9RleXHXS/3kVJbNg6KYNoGwXudXOAvQXT
zR8GEBXxb0WvqBCAa8MnylUt76+zWarvLAO6I1bn2KtOJZzlNvHYVCm35SbATJ37
Uff+kssJtsTnfDKAgznv7/xozz8BS1zWNsmgQCWz8q/jNEjNxOckumqXuezbGfil
Y8QSGNpI5Ofso9vZfofVeFvNfiudmsxAnB+JdmVspHW9lNc5dIwdBT+hQyfVbSe/
oVyi6TENlig2Vy2VRfKV2Mf2bid9xFUtiDX3Z2IAbCxEhNLsqZwhzpqb25tJBRp7
ROjZ1VSss/2tU7lkSHwcIrHL21Tm23wQMCy4U9UlxDn9so3m1xt10mxhBqlFZUg6
YctvSom2WxYtFxsJYdIAGKWAIEaToIUc9rjI5VA3YiTXSpcV1X4+zggiiPv0atk8
g0espJK6xwAmlYaLmJsjLu2RBV65JCoG5ZP+dK9c2FchF6BcARXIs6DEHhxhyuI/
FZl/g9YyD5N59BJYqbmc09TbTk68iBbZPzo35dD1j564dge0KncORRt8Pz0dZmvF
wnQpoiC0P0wdYdpiJeP3sWaud5BWJVQk5H+CWUa186B6H5NcRSEY55i/hYPee/Hu
7d0Cd8jhQhL5dZGWhjpGrqaYOo8drfdIgFd7Eo0m5f6/L1FKBmPhM9H1V0JY8+bw
g5tf5tHDZm/QiBtT5Ff19ZRohmDkOJVOuyZN62am8jd0TI/eg4w/Log/KqWlhwec
pbJlwtqE1tkDqtj4+GyFW2AxSqKCCfRcSHxrxFKu+sfh06j4/uRX0n+8+BLrACEU
bzIxcpT3O0w77YH0Yr3Z8g==
`protect END_PROTECTED
