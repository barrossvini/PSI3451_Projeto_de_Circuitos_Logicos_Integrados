`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eEeKWDdfeL7g2NhLGvDyzw9YShTrqqEVIbLrRTKW8k223FfQ1L7cChcJ6a7US6DI
DkjNkRM3Z3bfCSJQJ3YMQLLk4jyd7sY9IfzYVQmtbA+xjn3HbH6BjsoYFERBe+QX
ShVydCAcVf0NhxqScFD6//Pz5kLmKMiX+v/sPmtnhfAus4Qp0Z8k1jy29Qprr8qI
1a1/AQNm0Ce9Hz1TyZYSQOTiT1cRossY6RosL1vG8ctj1buQ32aGWPVkSEbgC0aO
TNAzaRXptpigLqybSfzBeo7NiZHOOF+U+61qX2M4tAkIVcDndNMI635uwvKi23iI
yZVYJ0hfUKB467fnPXcPKcl/FYkjPnBJtZF2wLhyfAz7jAe+qE1Lx+VtriX+jFSb
+y5A2MZQIMqbnsxmTU8O1P8WRmKK4a0JYJBQIh7E3eJL5l4Vr+wbgzyZ0aixxcyG
AgrVjx3Sd0rB5Kc8WRL+disBSUzgtiKE6XfW9VUo+S+jzYJN4LTR40kQ4UydkxYC
Jgx0C5LeiGG3YKjgrb3b6rRT97h2odDAHa39e4l8uPb2I26xkrWw8vWClJcuvkM1
wzU8kAAiXI/vWyjnLPGbc4SZPbsVz/wTJhz3vrnREluPFnStNdAaAZaxUW449QXP
bL9oEQXCLZOg9rKX/zo//KOaueut4kmI3Df+TR2j7BJtIbmvtLMftpKBaV7BmDlV
2Hzdy49oDXGyEPSbBd3GVogVT6hLYK8LyG6F1u9dKOU8RMw5yxWxQPkk+eB91xsF
Jvmheunce7q8YnTO7deBEm5sPoyvt66oEE1kiWEG1ohYh+jBycWs5ERX/eCzPP3a
rmgCzHHCkIn84ltQKQsFNgZvlwhQAquURCPxxteZhouwVa1QonHDsXlXr7heRvk3
LqITJ0rstESd/Pb9+iXLCe18neAw+ghOuJyTf5OOh7F+GtIOvu3nkZ57GrPjmTvY
zLHYpjSyq6gPYjqblXDXz5vVRCHjgcL5m0McvCb/epzT+Z3C5dsJfHpOsufdm9rS
9uyOMFDnVgayFDdkdPyO2cMb+Pes9QosOeWt/aTWDSoCUWCKdDEmjNfZQbB0mrKR
SvO0Pfcme/GyRl/7KzqstMRPaxQ80qz6jMNc9GqMUfbxWEnVRFp9PWmcbYuiUVQ9
/8AInjBtqUT/ExPZjzfjUZjDM37MyPlAmFC8W1Y820Tj0zBcWi0WxCSM9wMGeaZW
xpCeEHcJTTAuyQnV6mrzBKgkm9XeG7NShhOXaytAW7R6YJZCL9+TxVXq47SvWS/C
`protect END_PROTECTED
