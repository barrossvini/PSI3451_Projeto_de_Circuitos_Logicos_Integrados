`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XcsnJozcMKCqooRfWBVUGm1rFwYKRWz0pWeLT1UJR2XYYjfDqQi4jnj6dKdYf92w
nuH2vHoUKYaACiyq23RsD6sXQN+fkJftcJlIxNH8FkB8xbqoh47QIrNqCNN1q2wk
xzkzKScHvW4JOPctXqDMlp01XS71zAJX+xxranrL0SczhdmdYmeq80xEgRpt5718
eCDXJto1uHvmejB/uKvgZ/J61wI4Y1R7o0nhtIbJk41lBxkE/iTZdjBjRB9+dVbE
7KsYK4SIFgXedK8TpluiRggsHTTaytocNi8Ebi0EsByU8HYkKReW3sZE25yNj54S
Xbq6L52+n2r+v2I89LF/ZYYUWyIC9VHghRDVej89gTmZM3adP0jMXz7mrd7UOkDy
3B0FjI1vQYmhheoBL19BDpPfdIoaLl1i2CXoxOY0D9b3GSFIPQtoLF74FAYRrhud
Z1yNuStmlrMcN/V6Kpk23y5eInYc8KYWUFJl7ryv2ePQ4YyjonSbjpjAfxlKolvK
B1QJ8G5favwt4zfiiiwbYSnnlHi9v354iAJaXcHEri2dOL4wECv5BXTqZiV1U+ro
NlICc9MY96H3NMOkJlryoArBGhgh8ukc5B47a5xRVwvM3Y7qBvJCGW+25DPfH+1U
AI0EHIIuFxTquzCiVHekGPyFxyoXdrNUDPOvhTygi8Lij6Ky2U7hYtCP3zP2gxxT
iuFIrPJ8LbfmRQmtcBqJpPPwDPJ1JiT93oBaPY/1OmzBKaLCqLkdAjK+Ne/xBCiD
xL1LutlDtSPuA8cIu81JZ51E1sUDpOOG1kM1v+wS9sHcPQabyY3ATtRRC6nsNVpo
Ueh4J2jJn61hj0x6xCKfFVjYqMfbmEbkFuev52r+Lim48McTBG6O88oymISfye0Y
EbC+lThHUMi0cQAR+ilmLFM8rLspuvPYJDqERTlEfng+To6QqwQoKPwRKHRZjP30
POS1xTBURC83Qp/xhF35gmH8WoBS+71X2sgl8m4Jsqi2lWfcmLFHsVHJby0w+37m
0Np9l/Gqo4h5BOaXIbS4VcuOx8ayqHU6AAIuME5b47ISn2GWGXiPkTZfRX8vZWl6
Ed99SqWKqJLEE3cZhYNxKGh7sT90u7lvp971Y9h/jDne0erOnvydH2LFhaztFaoG
lqa7JOdVUuCcs4EGNdCF8pdrdOYMCe+C7cH2vKhamy77iGUuy3s832Ig/llDEJKi
IY9nPIzLz6h7wdlCB8yH6D1VFU3r4PfMvB4JGyl4QTrdEChXYjplikLzQB2sYMIL
elO41jMrmHzPS27UlcplNG9p7rT3fmHART2Yl1wE+/H1Lme5YkZkvlEH77hkxuXS
Dkqf029xCWmgM7bB9n7uXW5q7H7OaW0KxKjx7Et7p5EXxKVaECmzN1895hZqYdv0
4YgE9Y2h+1arB6YBjtvCmkOR0kqXHCmMZmUS/CQQZRCi+0UhDNXgbR6qUlstHect
qHl7oKSLVvDr+qvvlfIMa6bZr26zGShJGIGXG3zHsGFGjrNa/pQGeW8aTpRaI8tP
uFKEaGtUMCbxIWpJbIVwc16hyQNBYxom/XUyZtgo+ik+6QPM9VqPiVVDtzwZUbLm
NgYBKTla1zYH9ZsbCVj6fD+usMQPftaz1a5xpMkdTADtubkm6Cgw6V0Z/YsJJWyC
GlU9Q8kllDds3O4IWavmtkpjGYX/LOc4RlTvm6vzJUvLGmnvMIbRXhwYx3zBR0JL
3lDeL244AfZxbsNdTxMTNEBREt0BY3OjHT2KFibALrrx4NsFWyUPUKpxWlfHH+HH
DIGsLUK6LqOW7V4kOjkHTLmcbrJUn/WixZpRFjBkx6wiTSghA+zrqCb+cFTIPXpK
2G79ouyuFY+WL+pE1d/2hKAjfQw/2h8xk/I/W3/cGk78XYGOicQUB63ycue/2itc
YxU2ARwleVhf9TsENqXLhOfgzhS2MszOkDuNS66O+B7XvJppCiAuGU9bYyp/Td/R
3cpm76b9/cpaf53OqV3n9ZmvCaM/l+Ry5ezLaGidoxPQOkQm/XJre0XeVeBgoAa+
UqMBWYRQqKOmgFLcZ3H9g3zS1gRy62IJupijAGBpF/BcrFmoa9OIH+g/0hbDJbvT
DB84Pc3xjSm8s2jnM335W+pPaHFxRD5LR8Iq1GylM55STfMtbNpL2Y2dIuQ40Og3
PvmkXVHhrXNooBbAj7OsKE3KiwXFhUx0kslRi3gnPq7bfvHql/RWj/DpvjopsZkW
R/oF9FKDXh09WUBoJ72Fgjh7aR6Ii+dWm2Kig2Lm3VX6M98gKQ2Emom6fvQd0LHk
X5Le5iJRql5U8+Lh5QxoA3UeISFlK+s2dETheqzcv6I+EPNsry/XqPob8cQdxFyQ
1tb0ltwxrwmQJ+Rx+VlkhFOHOjqhBSSkfZZ5ovggHunTFow3p1+TQftZjz1KaMO8
OejP3SjRdlLUq42z/YOLt8zXYhE7Fnt72q+O0m7NnLnogaSZmA5QIDw4VaZBtEOc
VpsISnnggCTKDSKDdU2aV20n4/6E9F8sYyXp5sBmIsM=
`protect END_PROTECTED
