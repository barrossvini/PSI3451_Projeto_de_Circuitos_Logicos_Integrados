`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hxfWq25As4xKsfEQXtXaFEMXGMKyN3QucoVkJpZWnDkR93SBXGvCGDXUAbpKXxBk
uCIWdLP81Hv4PyMGxLcW+vjzQFTaCcpfhHRBelMUvl1i7YewSZm9W8BfKzqVN1XQ
++NulIQ15ZQ6xSJNIWau1o0KRpcbyIvoe0+VZTycRzTjAhxPhccOYmiDmWrZrkd7
OW0E38nGCRfDX1ACbCXz1TlP865hYaLSidevBOIVDv8JZ0t3v3ZddWGTFZ3i3Uei
7rGUZ42YGOSQg8E21UoEQiZ5VkeDheA+brY/6F50Rh2WbWVlbMa6kvIJE8blK+1a
/mi000CoczMxT6l3c21Tv4F9BPeznWu22SEUzQsqKE8Wpa2ExBNgG0OXE0TC3u2a
rIC7jUPw3KcLHdfPlKZ5Z3B3aD6B+IDw9Lfbu1vx+/yl2DF9cEp8kC9OwW5ak7Sy
D0cjPEZFFM09IkaPOo8GGyW/pcjd0hxsxGepfyki+lhrKBjaXHk+cdjj8BEe0Jdq
ES4G2lfMfoRxnPUvP4JMl6FqF/L8bDp9DWkrZpjWYFHRYPQ5T7PmJr4D8O64GFkR
S6YO3MX9w8LYiGsM0/WIahfN/LW0DIHdHLrJNt4MHxIThvsdNVdEVY07P3QeNODT
DH4+ftZ/aQjILym5qvRl5M+FVntbAOx4W/rV6b2le9oTBzppkhzIpLCUhX/2NFqZ
0Eo+LEa7o2cZZAbvfA470QSYS+1cfLb/axFiewsOx9Wrjy5zNKqGVtwJoW1JKUKq
PMZHuWbpuBnW6sQYP4dSd3enVtriCWKYMiCgTM9T6Y2vTuGBLZshUID3W8wZzFIf
fZcHuO8o3oP5G3aRJYMlaJC9jqFBChYMYtE0CfBd4yV5f1WjkEFAbdrazYODx8hL
`protect END_PROTECTED
