`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5tCDoW6jiZ2bnKgEgPJlrZqHDKWL8ydeyzPVgtwuQLqE7w9NIN9/cX/cObGSu1vo
vaP/Efn3vpIvXP6LC46yH9hv6rSnHTrtPzTu8xlkOZGIOt90qqV4xV/cKr6wWVJG
3ZmFXAJm58U8BG+kPE6T9TmYXOpOD5cb93huq/Er2CbuZEmZqQg/AiGt6QKmd/iV
`protect END_PROTECTED
