`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R8STBZZfitpFo7V9wgsGsiU3NC2H5x8x5Bwf0QLjVaAJErifaqgL/JvjDzljRRpa
Re7Hnt3TyFcsipzwaG0oUahaYJIQKZf9vIG7yQW/svA0TJ7Bw7HyWaIzjYTkpHNr
kNrsa/Z5AyEr085BJaOSMJ8AksSAR86pvzcUtGEmEnLJxjlxC/TjHmj7v7XkR+eA
AaTWGwoLFg3owrlvJetRQPzeWAHHjoF7Q2B3I2UsZnnijalr4Fny9rLpdeT2NQnD
+wPdWSz3WaXpXRolYLSJNiO3VJJoahqdPfD7ALi9t2PPq0tuEgic9HbucVLkBrcV
6v7+jfj187SkDKrJ69vF3v4v+FPDcWPrGh9RaPjSstXg8gFfvlWL2Jj7AzDmZIqT
V+y5uNQWbpc3FxP3swfC/s1ZW5fxTBrwubP9L+/DsxK5HZ9aZGbkRrsJMVhkTDe0
niQ09SSIp2H3Urz+6Zv4MIcxihWB/zYZ9K80SejxPrfDrwAxUiiPZnoTVKnJRrNK
MnOhoG9oJdcAQP8kMpMn1GvgRTljItBL7kH4vq6GlIMFdb0yhSO98bx7u1G2dDtx
K4C2u8uazO7WSw97fsVC7s1dBY4hYpTiOrZCh3q9NGuRnKKSEUMwf+6XEmasM/jU
oxOUS3j9S3DNITxhCx+P+akcJ9fctM1nQDIeuLWDWEYlKCh0dkvgNrK4x/DX9gv+
A5mQAT34wTLQr2Bi0LCX1op8GEUNLjlPQktj6FpemFb1IEptysiDB3ep9uDNgejz
XQ5fcXtLwJV0bfF4GC+ymLr21g9IqzMelzPovHqzhUCI2Evo23URCZheqTsHXlOx
GhLn4f8bFaDHxz3hOssb9T1lV7yZnuES6O//20wtUv50kxlLRrPJMbMR5t8sO5wC
iXDcmKkVhQkWWRrH4hhJlf/kA6KojOxZ76nLQ8UcFgfvomDB36z1Rz6vaeP85ABH
gtimAzP/69378l7LWovB0mp8WyXzqWNx0ZCqLKWmNILeCgNDr8jA1lkrzGiayT+W
a9iFrLuPD6PToFMH5No4nBvpJQbwCQdkdXtJbLOuho79JWBC+2IfrTyTr7fGedmO
p1sMZdWvX4PMOmcvtHAy+1/LrkyGd3maoY6GlbClqg7/kqzXLpX0ZpacRZQ7z1Kr
O0rtkAh8x/XLInRSeG8CfEBC1hJBrOgwUc0Mhp5ezVHb+82gaVxqAiMTbQgz8rk5
7c3ptGxos2oSBuH8IjWZwDQ6u0or2dBxqTEOgwzn8Hk=
`protect END_PROTECTED
