`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XtmLwMA5UDMjepu3L5L5HuqMLN8opFQUvTlfpGhWGwtoBUiXtVHD60B0Zfk9Ujz6
7vED44T18vhxVuNfWE+jDnpxQBSFA+x7Sw8zdWcX4FIO6w291QKIsZ8+0XE/1cc8
lOfZ0Vtb0kIdKF0iKLMyT2yw63RXVHcF0JoXAwYlDiDiD//R+KuXuZ55LAW2Fvhi
MQ+UzH4t78ejQDvq6fVpZOVsW6S+2Dw3dYzGR0MURTX7C+CmjqTKRtLoB2TDlZrY
nwhkEVqiTT0cGVnmizSbskDAhB8d7hhYVrsgRo4E41I1k2TVtVsuis4KvQfIIpVp
GFFmpOyPyrDm69yfk6ET6zflWl+WspFh2uV/yRJIic23Ggtmd45Q9W5bHu4eYia/
uj302rIrpTlkBN+7be3nEW7YFV4lCWVasYUfOJVq8M3NJH5SJpcPQrSbepf9B8I1
s6d4adfsuSyGXiCEd0brKm8G1RgylG18zalUh8o8aY+jscRffNJbuauWKREaO274
0MhBo8KGEpKLl6TL9AXF/zTm3r2HHmJpQ9ibT//sVorSGaiVLDeQbRBC8PnefdKr
hcuS3fgE++ZpgsyDjJ4ZRk2EbB9lV7XID73ZKxCmX6D5Z2GEDTaCPvz5BYhTpWfn
fsrApPXxH01Kr1VRcROVLEM3VYUP46Wqblh2KyTp9v8gKij6f1rdWyXrEypVSQB8
W6FCFDmcixUF37GrlBxg40ecUds2i7mRiUOQsiXT77YV/cxFDuKWI4tJpvNl5/tt
EIFAq80PPsBJ1udtsbOhBIs3DEwCKRcjJ96yh7KEpWJ0HbDSeLyqemvo2MHZ02Fo
myXPlZgenegvd5Lr4ZQiEPp2jJvYXoERUgjiAw6tiRIMU3d/FrppWrGX9JhXil92
Ua2e8Kcj/ZdZVn3CAjLh1IRd3jkEni2WpUCei0PPFXmRNjMdyefM6F/rDQEaRFAI
`protect END_PROTECTED
