`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RwGqgt5z/BoxzYTEgI+ZINTsHLUhlueyhYFC2sAvdTmrZx2YusUpyXDj0Zf+6v86
TfyDTVUxiEQ4Wkdg0uOBagUwyJfRg7neA29a2iM7YUpZTidDVmIxFSi5MLQPWxGJ
P7yi2NIuHYTZUpM4bv+9fPccSJ8kb1Nwo92qjii0v6vK3w5aMT5WH/UvYe38wWFe
IphBROwy36Ob5AkvZFw8wE89y58w/P0jb6Pjj6H7tvwmsJVDUzOUfKxWKsVtBnC9
H5XfBkQ1ATSu5RwmlQNJL0NCxlzQIWmkEf3DsBtDHpL80co5+NXTQTaQM+S2T8Lr
cGgkD3etXgS2ypFnb3x9zBAgkvEDCnuT2drc7Y0BlMhctOl9D7K/t9+lONoBcfyx
txb5TkN1lUVZXtv+xmnn83ymu1MOC9c5m5sruM+RA5p/eR3uQEsagMiPF16/R+Lm
KDjG/POH2lCr31EAwQOdDBe53EPbmQsZKcO97QFlGRKMpmOrp6ncKVmTXxbyIrGo
JKTxEbeanTtzU/x94r+m6ACEnt8cGqBAppMRVGSo2znQIVeDb1rXb3wEeXM3zho8
wjcPt4suL/hCofMRQfPYgG4EhjtwJs+z7oNcu40bw1iX3C8vB/XqLcDujJKa8KtS
KPmeSg7F7Po+W9UykPf1VB95Tdo/jc9mFOckP5Lh+N2C+bjkNQJ2b0Y1q7vy09OF
Y8UMnsprauArXTLYaeSpJDlWOoSztXXoWOhpVg2TAyuoInAgYn/VqivYmMsYFv83
kqzdudbLrQI+oLNFxLtZUqa7k6hYEj8MPgBIg444KJftCcSBZPdIUafanqSmRZnW
Y607KWifI1AQnjCSC8jnG7t3/jwgLLz0Rk7O3BwoTuBPsT5UfAaPWkEKvZZB3ZZO
OrgvOooDjcJNoYBTHIww8oxe2bW/gM8OQfKPrjWFIbUMrlJuATfuc7xW017+g9FL
CHGe6mBqZ58OjB/M5IVnA8YNFfXdFwalGQWIUxaVFNEcUItoyg+GZw3rz/RYMYGV
FrzjeOf8FfuaFZLJfG68d92q3I1RETnz1K6XU7/XZLgygLSxokNaYZQh5tf3phcj
0Fk/GfgblM2zgXBG4ZjOWmkDhUc2je23hrhnsg9fCb8emP6xFZ5kVf1yiisLCS3o
6inswly6pvj4ZkDUMuc8VPsrxCLvSoU19khsSHm0NOA4K2X4DI6XqPpcEab0fBZd
TSDEHv73MXn8GWfJQKJUKgS2p6RTFbISPNhKsp/9rj5P8UfUSRs4HXH2Ey3C73JF
COBl10FGrw4dy8JdTZGAA9UYlHgOFAfrH2nAwAU+2ChJtCInU+cgaMPOUDDnWuzG
xXdBJjgpxQP4FVE9TVglvHKyEL7XMN1IN2xh/+27jDOhpcY6rqOcaeZ2GpB76IrI
tC4A3BTixtbTb0O8dbGbeJVlLzvO1GZKjTBZpbgLm0ygy8asehn73BAUE12tapdq
UnHRY2nykCxbjj5QljcNSlCpLKv6V15N2rAY551xeBIqHdEy7+7+oPc62hpB66Ct
kmwNh0b4KGVMPdHdsLB0auefwuS+VrkWAheItjkiBDvls22swkLPufdlORZxKyky
myfbNm0R6cFM+CYS3//3dvO2nNovWagC0QfBsk2lAbzRW1o7sy1KZVCcOQA83F6m
KWOjQKUY/NzKnPi65EGAzyM9k3qSPcjupKNTc77boRiJLog1Qf7vrhxDlpcbIsIF
FiVlLvPeRkDvGaa+38cSH0Jhb4yQXbU12P4Y0q6Qyouyw0mpXZCPpTYYQ3Qdevvi
zkRZ0WW+bibS7KRB8pY5peKOt5UJuZoAgoz9JRXPZhZM/BlyTW70sarWZWXEXEBo
1RT0XzuZe5OqdJVNOWGYFzeitBxCs4bDSma1fz0CqcplpheLAwK4SZEIJUmq1gnb
Y2urGmIAHGVfWajRDhiVK54utWO1DJ3uLLKDD2MBpn721pv/Kq4SPPNsipEvGHGC
hGh+ttmBgv92VYct4Cp+Zo28JDUR+NwxKc19avE8xT2bClqfquFF8cATJm9n+4ON
nDOOo26d4y4Fx2H9d4ZaKkELIkXZV3vxCX5Yu9wpeYFNTmDdJJbCnlmADWDO3gWk
25NJq/0S28zJDoO2R+pWrfDzWICI3Cjtx7s5yuge3LMNXJyQqzsjoJIDL0QpJWFp
9LzJxk18u6pN/PcZoHAy03JMQ7K8OLvHY93sRCOhXR0IdqoSJUH32Z/Eyw8TP3n3
5pGhdgW5pyqVHOd0GKJsugDmN1GoKqngBb++U5PvZeD49Dnp8t8NLuBS8N+nQ3jI
QgogwyA08KClchlQbfQmLYzglGblos/xQPacv2NoeEaZMnbxjyGtmo7p+1ahLHk8
LfoY5q2QffyniSwW0UJjMgK/f2MkPBuLT5TPIbogpUlhRpAJ+or3DhhoLxbCV1yS
SaIqzTLOOxPm+rih0SARWsrXp/i8mplF0SbfS8OCSqzEHX/UST3qZGDjLl9odl2+
ud4OHLFaidP4R8M9TgP1LvsKbwJ+uRi/sFTulvED9O79FOKizDmtvp+F8vI6l7/L
BuTs+Yw1+3QSuo5Whdnpa0/qp0hNagpXCt/QG1+QHlXm3VfzntUaocPT+/vh+Sx+
CnclUkjAQal14oH1FCK8nNA2k1bgTgJQB2L4EU4zvsxo4gvvjQxFBGIuD1g4IZnY
RwmFmhKU3h9diBf4SbbabtyK/sribkMZUHl5q0LLPwXbdxFtXrKdDoGs5QjawKRG
knRQlH0mSO8/5pLPinLtcfbU1JmyZwc7YDMk6DAaNwj7CmZDgs+xV3w1xHbEhinO
KR4QrH7tknT1cxD9u78QyOb9x9s7D2cAdU8Bpf0LWl0FlVsMmdOe7QjI5qt22nI0
n4oc8InJIUTTDv2kC8IT+tshscJtpb/bpwubHLauRWdmrUNvbyFvlbyiztccUzcv
Bfu/Cgggy0kpS8BuLkRkMTuP7tMuNsUOhha3eRfopFgDEfhK80ns1ZyD7PUKro44
fJQWzEdUa6Cu2sO6KHpnlbSj7+9K7Ni8MyVi5cYwroWb48+DW/GhhrSrvOhb3DFu
KaZyFBKKwNdJsmpQttr87LVxELsejq810I0dxsSMpOXaEr9LyeBYH6iFNPOw+YBj
mRyjfzn1ZPLVzzi/44bsJlgTwSDDM2Uqir0n5zbccqvtq6OCOc5KGPzjzXvNboh8
vvzA5xBRSrd7s1X6Ak+tSJJA17bCu1Nu2eTUKFlNas2/hkDyi5+ahUjBW2MUn71S
NpP6sl+BjfM8leOil+5E8AsudWs50NxEb479AVK1+V9BXx+AJSgGfmomlguTZzvn
ThfH9yOiD8ZH7JLADMPVeSlHpqQsaLU2Aewie1kwQg4zybeQxPHFsddB27ABi/YZ
WA5Ck+lwxMsyeQ9lhTE90F4lIfFAbQFRYdWLHXGx9113zNyXjtPHe3I2oTMxRDZt
LWWC2wRU0/8stxe1+Owc8oS5HQBS2Fk9fSJ3aof7K3A+u+eJLKGLfcBQIBcUU+ao
acHiMWgtCjOlO/LJf51YhW9tyyf3jJT87wgYalRwjmturYNka5+7BqfJHNT7UQIW
cV2Ps68qOhIG2vLrcc4HdpgI2UJOvdtXD0DnU8HZH4MNzYLoRtOFSBu3en6sCnPO
YL4Oz5dwPOBurds6irrAdA==
`protect END_PROTECTED
