`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ENdVgH8eVRTfUj6OjXObrGzEwoMbk+Kcdnx1fY+Gx8DynwdMEaXill0nXJ33eSD
PQfw7pHzHCaFasxDr7bpMlniCfLK6MO9dQt1KmL8alIumxvaumCH5+I2NtECoik3
MlB4piWNFB1t7e3YOxFiOQmSRJ+Ml9HKcuS/GNHfi+aNCYT3hvK1SU+rJx0B7elx
goJNyF2cPRQcvMT+dOlwrJSGu8y/NYBYYmC9yFREjGSXQ7hPJp3VWzdw5QS/Y9bG
ykfsP6Nr4yMvfIZLHT74qvm1TkB6dijBK8Ig51n/box6KeD3SIVc3U1XV8+CdBWI
AIYQqj5EhRULARSYHRYMc6bkMD5dVaGSRnLHEQeLCmXDonyh8gb804Wh7F76sSEV
WoJjjIOrzU/RaxILNjHcyLW65YOvA2VgXZXSHbi6UUJUVzWOsHXWtN17mAg8cF83
jIABcR6Z4UcivRGuuw8miZnqZ6VGPq1NpIIPqZAne+bv7sA7MCul9aM3lgzmPBvy
bc2TVOblav9rHOT/MyYF5w6zsOy7TLjcjfHpVRQY3Aq4QOvRvTBzo5UD1umB91re
8H8WGD0bW+3sYgy4XdK11KgEbHxArgVmq/XY5/CBn3slJy1lF8ld9fre9R+ma6oQ
C9GzXRtZ0QuZEJPTSxm7BVEdJAo3vsoYEFqGJ5fFkNNwV+UEZ38xfbxEhxSE/WZi
YtbsA4MJB3ewOPnSjYJxPzWrzU951poVfLqNdcXYseDf4OE6I26e8BINCxu6jkZO
u/k8mliW5mniuVnf3LYoiTJQhKPjF+TQDVuItDQU4INlrmJrOZxDSK/HQqwdBUJx
HYLwBo6CIEiw6HL2MfTwFA==
`protect END_PROTECTED
