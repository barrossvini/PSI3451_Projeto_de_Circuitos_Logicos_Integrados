`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uA4Bng4txZTucHMPTKKAI+oXUjyOtNB0ob49+o5VoPFY2lvuKv3h+Ma+mrGjbFEX
lYEXlP8cEY0SmK6RQRhGAeRFDbpNWPi+Diz45M6C0CWZ9tyehL5jhEETXUcB1VJZ
Wcg7CZACh9n09lyAW8gjLAPNjZEmVg3vr3KT1vFr+4qWMF/j8qpYIRcNEXSGZx4x
u/tQqKr9TH2rdkrSQMPb0fBpsvj+F5QzHMJVqsQOXtFwszBj9mnHIx2zGy6ELDhT
C1YYSyyY6P36zY5YYpSdE8KdzkC+UjDSsXNwn6mjuQuWa52b1lTT7DPoOlSXTFey
KGMM1LjNlQb2YNKoAYDUCwnj7AsTGHFAnwClaeFvaTQYcovoLnNXTHx0yQikW9kU
HeStMK/mrw2a9C7byqAKXLxsJqpsP+3MiGw+SCrSv8XslmxVjAwsm9ID06zIMC8q
JjmKRfzgS7khvr5otPSdf4swvVoSdlgDSoJg9xvIBbA7Vi9sZJTY2KU/muNJ6CxX
A9LY4TtpW40l5OL2bD/Q+x3bNv5mFZQQel+WMYnWGzMA2q/ZhQKgfzr3x3/UCfGu
wPxIqmt+wElYrHdRuwuHyWaNlGZgMIfk73m1TnmMn5nRxJ+Lese5pQjEiNaOljLY
evhWd4fkRBed3b3EZeOH7owhT4fOCwz/0Tlns3rDYVJW39kFfnhfsr/mHCvPyrYo
4qtOumXo8FnUX/4E+TSoiLyLg0vl6QeyAAr63n01gOXDmxixnWZvgy4KwD0YCYNE
JaIRXbV+HX/9GXSoWxQUCOYljVWPyDDNhR3HKDBuskAoDmi0GimJToL35uWfzauB
CqI44UBmAmhNs+UwtEGMvKMvXOOGAAYG/DX2zAVYEx/ukUuIZpdMCSJu0DPxrQrY
jkvcVQvEpFH8L3u6mESQDYjiipf5GD+cY4ZUKrF90cG18niBRQQvJyM3JHyAEyQO
TnTcgytTSacExM0rdDUuh+y4ooc8iJyCaLiTUseO0XhwJQrkqnbrrtxRUENG6rPi
U99E21vLLWALI1dcR/USXzEUJlrOimznmIko1CjWjjRHXNRspU/qCuBMVIY6LPM2
/epEgcgs9ngrw6h+w2ap6aOwehavGp6F405TNlfhjrFsj8k04UnjMCL2K5dpV0nJ
MjqrN7ASu/bcD5BLLiaEJBWLplRHCGPIeV+a8iZPbSnfSYPjPqDGz8GVPmQUawMo
TIYu2OGtYyPdT8DAE6U2okXK2cAuFtVqLXAg887jeEXwRYPlRCG6Olim+Q5wuH1c
w2Wxz3d7kywcOEygiFEHj4+Q0kKQiioKaQcYrPtc1JjPqNLNh6qOps6jmbx3x0jX
lHEeFRtb3ovfWE27ddKXGRYQQstUepmA1YIWG//P7mhQOrXqeS2z8EGWgH5u/zRC
lFgU2rNV3zQVwh+Z4o+NfCGLae/ISfAcZgJIK4PJMrFgdaMVenqlPwBng0LfF5ZM
1LA+c9OgXlP8LSpHciy3vMb+Nyu+wpd9lg6T9m/cQXAwKy7J+aVII1/ZoSxhrB3h
QL6jVuHASgSpy/WBgbyWlNDq3VNmQbzXvhsO02JQsbA0W89bhhCYBjrRR67Qs1AP
HMS6N8KULJd+macOJz9GtMyw6YRbiiGXLAkA7Vk7IxhmbJVYtvE8ft2bickNsl0x
zdkIgto3UXTIsUdm96EBAHOzPfaHJ2U8R8aMJHkwZPZRvT4EVAMxObFtLzAZeKIg
ixS04wJED3CFgcPM2jHPcYzmcAsBjljttqTq6RgAU60ez2abdzW5iwfZJ1BNSIVg
2vgpgOsWxlkL7gcBoT704ZHQpltjNXMUR9smakOcMKX3DqJNL3AXYV4xj3pZrzlu
Tnch7Mi2ymJVNrnp2e2A3hKo70UOWKT6ypvmEfozXcVsNZp6H2Gof5t1xWOkvtL/
4WV2UwCHrIa6FppeWM+PHn61yVuqdnOsnXDBJylQMZluuTgd7vlWhdYgbLXDGxxb
+jutgiappfQCHQ827i6VaGvR/Z2cv3XhpIfR3rq0TpS2iIiHmKL8g13bTQMdt/hx
tdM17aXRDpo4X4rvU/LZuP2o9oy21mrGzXLAD/Qg57fpBAJGEfGlafIn1FKcjyX9
y+S/W09hFcQ/qbPBQ7a0f5V/rqVhjXEOlAGM7AZ3oTMB/rwwon86OhHNOoo8UHjA
iXNMNIUGzxZBvhR0vj5PmHIlai/pwSk9FPuUJRjMMxEeOUarkf8hGHtPUiU/atkS
7JSDc3DFJnrwZYXWmdH766zzLezcx2kqQzvuLNd6CQHF12dt7RGHl1GFiCZtYaef
oaJ+YhV6SqmnPEqUx6mUphaQlkHvEkZHpLGQw2KkLKNfxQ/lV43DmB587psTuKPN
zB+154BZM70Nm47Bp/RWN71pPa/PcqhdCm1Is0tfn1/vMuAf993MrCidZx/Wz1MO
mcZpC4b74YMLy5PSm5ZMYxJRRf76t8PKimBR8Cssq5bfUhx+mTDrVLHVcietbUKz
Ns+JDuW+MWHsSEaGTPkv1+9jYbd2fn3IcQfRVdJOGILjMdEzi2ES7tNf7zXDiAxo
jPoPwZX1WqS5pcSnuCFlKkAp0NnBVg9yOtZxs10MjcYnHier9oH6j1na6AWBdV81
tmlRyYu257/agTDxMHSlnr3/jRndsAWJm+dZJDZ99qe0XY2REzrzz8fmt78bDaZZ
IfEGiUjdIdfdkpYKEu9oTSKddPCQrRKY8OwwyWU4PvXi268XTPxsprq1wLWbS9ZL
tr42zS9ZqlpQq6XZkr/j8NC2jMIC5M40XD5te06BKV/6LEFpNw9Z8Yyc3mRDfiUE
rD5U/Ogx2gb0EGAh6eOEcSWB1PXzOVhtQiDqG7X54ollCrjrIwYvb5UxbWoO8Mln
m7gzTDVYXUfFentEVhYMN4+4w7t31zUiEhHd9yQtm75jujhjR/8rvO7Iu/4Sdgf/
aSC/Zcm2OuVnwkxu3klh+HcF+aVQ9rqhhPv3lz2GZs+Vs1IG/CUWBKcHe9vpqx/w
VpO6FLcylI5TIWrcA/JjhHAYJSr1U6PWNmVHDaSC1sebFP4ywXhIcFsI0leG7F+V
+kmDGG841Jm/dU3BH/rO+i4hlP87IAT+d0/fCliAnAPSH++u+ES71g4+BR4WhLKI
2Wi5x788um8OS7NoP1lBdgfqlTqYYOv1fP75JMFCSd61Fe4v6zLiMFGeSxUj6lML
NEJlQ8GML7/AxF4k79g4chl6ze92EUavwo9VooTtnHqGIWLy36b2kEwNVHq3RwBY
zJzC2hg7vfdPIfZ6BxAHa4VOMrWZTwbDvFa4BqMrEczYXRmTxvqlYCElZDeYwxGV
tlqdyeyA+rJ1vAneUYfRMSore3rXyXpmFLaYht5+9tOWRDTLE8Jq7c3xhK6dLjLm
YoNvkK5Xc/65rLiWSDUSLVoA7T91+6+zkH6JGtFwmL2AfYtO14hgnFHNZsG4LbW7
Wo97kSAwsqL0O19Ui/mn510rpLjgWatFEvXl0/BaCMClcKlR0lEyhpw2/q0UlU9/
oDuJIMbcMPTKUE39V2j3hKYQfsypNLjiddhAZl8SftVJk7SBbNbZsIQY/wsUjnim
gEjJjZ1473084sU1VJymv0B/8Gff53XijfLkjUbYUhXIaoUnX9fnx+LjarnpcNUP
SPoxZhdacU1E7gLJvFe75A9ttoU2Z9EKlb1qQ3NjgAxd41nu/kUM6mtaTL9DnqRc
I1KsP8JZewFj1AFKPXCZFQ==
`protect END_PROTECTED
