`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zPtWq4GJM4OCcpuy4oqv/Bz/C+dhryYCzP36oWuk/ZVYI2ymPzTVVTNrB5jeFyFR
qH/o4n88Vs6fO4KQbxBHKpbHr9FNdBP+KcFfWjUwRQZRtvSBdomX1Wr6vsOL3M92
/WXgnNsRm5FYkXNSvWq+QyChWCdeOjpNV0FsPLFKLtSPrAEi8ZXJrZ6tgBcfIRzl
FF67wCLb+B/d2sXYeI1f8ZKRWHcKBsTO24z/rhyjRGpYSQPCWHGNY9njigA+zpin
OH3iTSIPgwj3YZm9J0rIkVuK3eXJ72RSS/kdIpZnw2D99AzqwWAQS3uShHDRIQKZ
NpWRMTFfdqicaizMQcLiz3NfxsgH1y0VJ27RWOLVl99PDAmp5qxd/GC0hKVtByWD
ycoEDSp84rKLGgWs+BN1Df0gP58txzl7DQWMvJN2dnTQ3zA+OQYQ7eakf530F4Q+
RJDG4Sbk+Au6IZsTWSN1og==
`protect END_PROTECTED
