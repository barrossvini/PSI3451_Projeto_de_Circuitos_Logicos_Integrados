`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gX+25oGiSeW76VsdUa8PUogiEWTwsdzSp0T7g6xKNVIj6tnSqsaJ/D1JJg13VsPm
b01gknZB0F4ksCwviRnmEdvymT0KvUBucGywHLK703/a0B0NoyD2pIQSDkwLezPg
Gdf26G8F7Kpi3rrX4aj7uAcBuVh9fEcIJEQ/5Pc3vEL6ssnL6Ve59VfSVDMawTMg
1YDXcbH4GTXs2bR5qCVD++1BUBQpez3glwnfkPE1QAALDtxPeE5/vmyrISFceZMo
PhSKIGatsppPI10Pjo0bP2QMb0FYqHaFe3Drft/pdHrQPinc08hhEdnhWWcnVkYS
Gi3omwoIi9f6I+g4kfiTyGcEv6ePu2PSXhcaSe+rk0ERVImr7bbFtrNljYpvNX6j
`protect END_PROTECTED
