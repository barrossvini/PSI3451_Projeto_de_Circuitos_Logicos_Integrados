`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s5xdSASEWST91d8lGqfdfgIW+J6UtFQz11yIt4lejCdAtzzYa5qQ/nDk+afuwyeR
0ccIELdo6FdUWAknGsP49rqP2448hc/Wiv94zqWrQdhDCvs46yGbLkqb93z8XxSv
bploiCqIRzGqPs83rZ3TxNjDTP3c0m2A49UQWUVTU57XhO+lGljMQNtmOzHiIMC8
J7wytuguQPcqPgJY9k1nvAvauHGkAHDe7Bj99lf5Mwqg82p/svdo1xk+BGSi9J1I
z3nQUf2NP+PCdH1FNrh0OVuduNMlLA8JyIPKPc23yb5I7VNAW7DNPLPiT2WvmfuT
Sh0+2JLpIyu2pQQ81r0+3i84ff+YWRQ+i8ZpTy/rKJYS+QlkV6tMT3uDx7j6xBZh
17v1t0plDEUwwXxSY6eYtfDBkVwXlCWBosUN4qkyG34rm+h2jQq24vS+ue4GaDtM
e8cBpHyk1qHPqoai2H2JeAinYr+ueW9JOYyZnVY5SwXYP62LQayecfAWHBIG2T0A
U9j6buYyZbsRknw9PfIPz3DV9V3Lbm5YFgf49/MnTFEjNG3KwAsrbKQIC5PA8ITW
n4do/yWf4czuoi5912DwugdqQu67Oz3L8h+0Llw8xhHKcB68D89cHoV1j6ZBMuxX
n8ad4DkcRas+vcr4ANskPqsJZk4DJJ3vLfiWPA6RlvBFi9i3qtycfXSsPQ3+g37o
MdSm2FOxx2im1p8P1jjiMaq3wVQEeBp2waC6U+ETk4AHg3WEA+mclHKRofe7NaVD
4MEC75W3uT+/u1Xyc1tsDKyxz1PLDUk5XcLnrE62NwLOH/XEq1mEFsHXkCdl6Uyy
fU+sRTQqmP7RpvXXaxee/TEaSbdonGFTkTSNrFROqE3KCXJQlJZm+nBSb/UmNZ4F
YvkRmiw6RSYPgRwPMJMaEnWn/5L4A+j1yiHQXvrzGr6Qngvr2bC+mHHW2bR/lscu
rlJVPbDrwFqhXmsfWAIy5kWnqf6PEKSc6phbF8emIVzmMYftBQCGXogqv1451CCJ
mZvHQ1P4IcHp51Ll8bLh1RaBe34ux9oYRgadzSuXus74DHeIPfcCEHK7tN2IDptf
v1PYgYBDd6fBL5K164/0zGhSMyrP30FG8TF5f8PQwAUISjGBdz6UiBBSf3nl7CMa
aXBXvjHBeLg1ZzDNLcOFUr2Xxz200uQQXw+TjkqBccJVUwOCvRwmnJftUvb8cUsP
L7Gklb6gKn8rbgdFMU+bhXkS7/iYgG1lt3+eIfaM2f2NZbVyHPEkPL8pMfF+3PWg
NQqJHIC6G5IAJZsDk/3eZSkdJ4OSe4MxQF0poTPrljWJwcLf0LaruO6ma2dCajEf
niq+Lj5+hu0o1j1jZkfUg4bl3XIwiQPv4x5vQarkaaJ69DzSmiv0g/jd5SXin9LF
QYnVgbQl9t9Hb28aFkMJpEX3mm6qfrMaan+Fs/yWUkxX+1EiXLn71CCJS+BYi5fU
msQAalWqlk2gV8Pt4vA0AV58JWXuxGBQRdaJBoyVIFsHCt+erAFrJwELeHg48iAH
8CcIdZqWMUKZA8ZjEHO8Kf2hCq8Xw+Y/y8WwiCQOFnd8graWOp08i6BF33TJ1Iwz
y+CsPd9ZkQbnE3WWVdLzmMavarfG+LQnoiZ+jAT1LSRbtDb0q491M3ptdQw2VdpD
hAc7bO+rcMYiCL9l394MiKDy2V/MTC+RSe0CxpcYpQ3agUHp7tapRGqDAHMbiGmp
QPasiPtmZAQIQNji6xePXZoY7ZdqZBG1/aW2RgwzHHixc51rO5DzdZSn7VlwVZu8
03NrdVbCW8cBUEjnJZdKIGa1yO+j2xcj4twR+DXqrj/r5Rjvpoc/fmW+thA59R02
dkd3lJdz1+2aSlaRcFQ1+fZ0tccs0qTDFZKvlOtuzqLw+f0WTo8vHLtv6ilRgWvL
S+kVbycFx1c9yiolBqtwm/7rBjPpEK/LaqvyyTtlLMI2UOrP4BhDLWILVwLuYVZO
GrcsnKDteVjTXm5j+FPYDKnK3ftVmSpuKuqvYoo3+0bKGvJJW1G0m7ro81pkalTo
nhfX3XZC7KbjNx8EJXBoIBfRNdCDSQH188PSSWsDTXopeUC0s384oZ328TwPUni4
KppB8s7b8vbpUPpWuZ3TVnpPs9aRd9spVALg9eo4VPkij8aNMIkjxILziiTTrCuV
pCWuTyeCbgLY6hx0UB9jQ9CVjYr0wih/NJhr0gV/XK2Xjmi5pS2miRiTqMUmFgY2
06A46MrPrIZBb+bhpo0nD5mJuZLVCMp3PA8brRAJfTaJ8pNYYgi9H56k4Gfb5mPB
axv+PKqoastZgPI7uwlOqPivchn4WBH2mxUPhG9KZn8H0WdUOJlyc7GmOkM0YPCS
X26BK/y1IG/y/EFUiwJVUIXgRiKMgMH3TQUi58Od01SIsCajRKp7J4NzxdASmDr0
S8tdRo/3gaCBEbTQnPp9H1RwQ4pi/WVQ9fzwVCtJaRmLHGEAmLfhRv2Kgnv0pqyd
LTLZ+63V8cTs3ePFGycTDGXjZEZjCx9mTpYPqqlor1gB0GwFoO++7FL0/Q60oQCK
sSW/PwP5Z1OpCOVjFQEMhna3BIoAVhbt5kDJnYDGTxxfHb8kRZmZM96nVOW2qDhO
hVMKD6B3TwXTF7JYeYWbo+HphfsuuaKKmoFbQBv6Y9ZgjHfrOCHPKJYE3ctfbpKA
RWe0Auy8mGXiWjlWKSZnCLhMR72zY98lgJnoTaT8kOZl9/hUrn48/7l+tfUvC+G6
mbtsm08tw/peprCegH/VjeClZd//DbxJoFP6FWzxynwyCjItNsGEPYe+vTyUTGDR
hvCRNjlIMlGYMXBCneMLBGT99f774kACAL0m9nytV0uAmWabVb6OIWpVd+1SPoT4
6SQ7cCv8ZfRQ1UQTn9JsqHqP6107XtbZzREKD2zWxzO6YuFr0MFTn1XoCsC8PExn
LFUhog6LUwFe/2N1eEZJGU5b/3R2RGe6UnmenFOwRxEifZovAKB+wECqAJGGCD0X
0VIgfuiRmW0XTOLW8ZMxtsPKALIlAhBkjTkyKU0vhrD5NfwWQmGZMl/bA/U3V/Gz
AAr4KJBkPyydfOJvuu1SWR40+V9EzKcOhgQVM5wDmeZezdBPVcFgaYWyGi0F2A3j
IwCCSGNfNxIg/bAVP+NrNteFBbcs6fYDP5BsI28cqZkPbRdaOf5K7cOFBs6ITYot
clPk6V37YtEfemhMPxvgDXcjaVruqbz2uOvk7RPU9bqlR2H+KBTOIaZfd0U6Rkdz
6puUikHsxsvKqnSV4NC05q2mkHjawg13Se3I7ubxNz9+M7wMT0PVnlkTxBl/4U0v
FzOePTPaveicbLgMTJZpDa2UDaDnuUQHm0X42IX3lfkMLJPMOrRz1lpOMtcUxfox
Ef6TViaRk3N5Cz16RLDBIfpCxH9ZDloukvrI65yPSvxMJh2dBXbxmijWlLcadAg3
mw3SwoMXQQKYpIduMZo6WuTwkgHUMZuHjIdmUWZUd7oh7nX1yP+zF6Z7xWZGcS3M
yijwN17jINgK4Aakf2owVPWMMEQLt6anJAMfgJostbAAToVmIWrTqGE0DueBwLWp
W9JESfKupg9G98KKr1yW+Z5irai+iPVHqCohHzDPr7RX9nx9w0lRE9giQApUTymm
+aAXQIn5PYeOtzKv/WqIX2H1E5riWI+2NGLE12pDch4m0/TcNgpXzs8oA+cxQOE3
SMJGr89VSsuMM98mXWNRoQ==
`protect END_PROTECTED
