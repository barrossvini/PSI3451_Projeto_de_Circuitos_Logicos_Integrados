`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
li+6qkbwHic72/KRZNpL6X/hr+I9hfBK2qD39S3IPX8npOJJg9r+PE0A3T6sPEuw
LovT4jdYoIUrt50QO17LaceSAPQdGH7uGfUGjnd9qjjCSBbcYA9uv9eWaMBC8P0j
VSFPUSNA1HOpADS2AsxP5BbZu2iSx7n8zj6Zy3c//DvRmj+BeLm4LUwPMg6GIKNr
EpyE/ZEho+uKVhvwsL1CMeax7RQBiyB23lH8FEqJyvZeACKMz6OODNINZ38UOcaI
Ug2k2GI0zbxSeLxjtUjelno8pF6T7clMLE+4kCd1gVzD4l6CEx0KI68WaXAjYCRD
jfqy3oQGbXPbrixgD0JL+///B/Pdii7hrQWzTiW9dib+2Qyy93NUPMJ/jXvEjMia
FcXIMcnu8XorsLyP/ntPg2IRY8GSvFmOh5PbzDZChfCXXBFTu9+mOSb77gFpkUZY
OlaX7ig4mLa+7FrFZp7fExRpKjAPqqiy4tIY6JVIFSGylLvGulENISUH2WUgVN3b
qsvBh7kopy1jk2OPl3YKNeWrgHaz+7COKV1ll57c5dwcGJQuLXlSeFn9B80sZQhF
5G+keNP4TL0k4rk8yFv8y1/iP9iqWiJUVFwa9d3gkbJX4jRcQbW690OSJfNQYfbB
SMboyErWNhB/MH17VzunrUe8F5D/CU3IHSPMFIQrhFji7GOcM+P+S1D4J+6VsYbi
Z47rep5SC8JK1S4FpE4Bo7yBtZdAHciPA3o0NG7gpH45bveQ+qjgmsMEUPgRGgzL
zaoIQsveZOhwi2Jbkodw7pNOjEHlySz9D1UbbClBrVAEqV7WJHo1sBTri/M8+GnV
KwseHl/z8xjhtGdHCCCQe3TZ99uWXg+CLUrD4EAoZosBx/X67FRVfxeNuc6l5dnr
ZbroHVgH7v0/HvQ98LYtt21YqapXhC7PI744SQzFHFA3YhM5x1N/pyU0qUZqmD2h
BVt7PSK3O+dUoRI5ow71S4E1qp4syUCPVHXwOtkh4KfObwr3K9IVsyRKJqmC4UzH
ID7H4cc7380y5TTI1JXHSKCBR7ZTMaQn39Ge3vyhkGjcqozFHQKWEzWg0txRltmv
NYvOS7ym5ogP0UjdjCZArCTeSJ4pCLZd9LQMKrmZ8IK6phl2vLGCjs1267n5CxgU
HqFQLBM582AJo+58y6s9ImilN5OaqTitzQ8CKoMZMokfd6XgiHXR8ZQCZsJjRl+L
X9Vm2bF4CBHMXTQ/2/tA+qzUwcUwNudRuKsiOVcfGQsmJSz0gGjNvuzXIBdqXI4G
oUg9oURmdMbT6BRiGIUy178gipNPhxkA+lbM8u/yyEiGg55R+FKgOe4VSQBAdGCZ
0ofoGfr15LxG9jGH6ohmqm/gBSckB2w6yvYe0ZtkyJMj5JzlDI2BEG2hPSoMQavT
tdlon8AE/Q2MjoWqH978UGBVhLNgwFPFZTdclxj4u4xMDnkG1nFoSDD12PBDf2EA
0Ay+RNI0yr3TLSYgJdM8qzsMM0FfJxShOgq+OI9Zknf6gX8c9dU4aKGfFODHXwhj
Z/gSiL/HC5bYo/7ihyG6T1cdWzlGcRrpl2DdExm7CrfEP1CmGymHaFDSZtGn6T9y
OtdW+SurdlhdzffJx1OkVbNO1BAjSfVGFyc8GrKnGvew2sjj9wz5b7skHUrzBEM4
Erhb5vrAXQHrGj8izQNUYMJvLoijjFPgwqiFWBuaPowJ/qYPsqA1khGze39ta57V
Flv2tU7YrFvaBmy2KeO6B4s3yX/noRaaGOCXpMVUn/qaXFFSvKxTjBSziD2b+zfA
v1oJc0ni5w3YseVQrgmA4KQpdOQcLJC0r+Ey3GEa5/ubmabD81BTyeSOOSYs0Sjj
ZEv9Bq1qxRulx0rrHEih6LnlpY4aIXOj8B2dfVPNvhfjbrqJt2Y9kf867Zda+ywc
qtMSSuthH9aPqMCqc7Npak4iZxcVHw7SjykHcn0cbL5tvl8QamgWSK6w2JwnIxYY
OOK2KFodjLmiZ8X1VC8YCR1rbGZjFskn3Y2oaQnISBfcZjZa8WIy17EnOx1+Pcu5
l6SkFjydr+9NNKL/GxN9id7IGhy+r5pM3E3VWJnbFhdDM5U2qrA07p2R7gaFWgwQ
Kd62+sQcLO9gMtN97m+AIJuDTZUDAmDJOd7cS3xXzIkkZaQ/y3QpQNI4aeZTa6dd
I8naWfLXiXGiv+xnhYuJhj+06Qx34Cc9EYODW3T7gEr46lWElU8eJv0u4bju40og
Lt0NCZb09UojucR4zOKoyl1OUdb8wlO61jDAWUT2sjBsiw8eqP/Sy+gMTwmZUYQz
WgNCCBVthwLkK223TtKYbg9qwXRBDZGzJxPNLbS1+ChF3WNa3MaM+iD3wxPEM5gG
abuKzMWXdJmu8N0yjGilZkm8UizgJqgkiuHFuqIP7XGzW3q/XuwWqpwu2uuvg08e
+GiRYE4R84A2PL/b11soL4kKXa4gJD0+IvobBFBsdD8ZzEB5Ywc6YLiNx9+EkPj9
f6t/yHyP2El6nSPeXEmTsG3xZpxyksF1yvVsXQNunoN3TDMWQ+QQVJm4swCO33JM
c0Swk0l/UoyB16aRTOqRAU3kXJWskKFAIl0nvQSZmiuEqVbrqWxpyipvuCEglpA5
8gRF78dbFZEhjniAt8s7MPLTGSE31IZu014g59i3S+Am50VR9doGAhRqiUEWN1v7
OLJiBIXgsqR6MEo5Vmtk2sHq3HkD9nTIibL1QQGVuhct/1oK6mz8eoM1GaZjswMI
Pys12VOGVauEVOOiQS0sqnGXrbV2YOM1NZj2inkQcpLEPeZ9W52uV2WywYDQK4ws
qAEji/VJHXEElSJHz9eYlyy/MqKDpIdVlSGkLh/C8bCaT43g4UYRQfcHWYwC2Fqv
5yAH925w80Pb3ZTuL4e2GzcsrKqQ+26BVGR1vByTIbuuMnxQUxVG5soTaBk7jdpy
ksMHWkQ3up64iod1l8sYyZWdx1dQYk9oqrT/cj7Xx1Ud4ZjcsUgT8yiBjaoqeT5E
CVcVj/r6wq83EeoN1TJ6OA9JX7oG4aU5BTHTXda2fZV57JvfE3vsNhdZTDekajOF
b8wbAIV8SHwxALl4VEiQ56ANG6otJE2FPaDldunNVq1XStB7vJk7zXd/fwbboffW
8PS6pbNwuU7IqJhBV2DJWE1W1C/dsyfd2yJeE1HSQLqgSbfo7/Le12Owj/MtsvCh
ovHcLsqtjeMibwOjzKVxfHcBEfila6a33/fs8J7PxiUm84loHUmUapgFpkaWt0om
i7iIWv+XmhI1TjqzDFzg9/5K1ZLBvQKt84Y3xLFhoFOxbqrP5t0PgMn/0EZv/tmy
yYpGIUxiAWxbm20RV8uePQ==
`protect END_PROTECTED
