`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1z5wMOr+37FJuzQEWEaqCp9w4g+xXUzCdAgLN3GzizAeaInyMf/IBu+rY0nZS8m7
cjgI8jEZ8+sO0r0z3xd7DCp2xmuchwBaXI2IBjYhMV4+fpSKEWeP64w9oBpRWiHD
1DdRX3fi984nhR61XiMD/IATTT5hSSpW5fpEq1t8Lpow1HloZZkC5Tz1QXXY2r1g
WFXbDPlkBTh2rfRCXGtG3I86IMDLtgOySPWuQe8056G/LsE97YYMKhgQq0skPPrY
zgOUFmv4LEUQwSeDMV5BuJUEReiONMBCTOfCwbyisYmkO8HjcbKO780ZUW7HQoR3
q7yiK/FbRNCAa/d2nglk0bjOqfSQCChUbOzj5Fqu7UFsWElBD9/k1wp+busA6oa2
CYCEi1yvpfqNrMhPtgvxdTZzO1nRf643m0VPWJIg2wYeqUuwS5c5j4fp6DBHllUp
5g7FVOk0eFrfWb1QlO58GPOcE8iAsJ8AgsnjRpEgLPWs2bZYuIkFv6B5dKv23TWE
Kp46EnwH4tHXmLm0JPnLPkLlOa2PWWn04qZLh/FkDZsl/zxWMp2ySlHaHH099Qoz
UY2ajwnoNB0m9qjPWGlmSaDyybvkdyDDkUrgyUbESUWe2/S4thmK0jreDi0LhimE
/VySG40CoRjFXJKwydX2wIbW0VbDtc5qd4i/Txqj0YFsCDLRdpb5cBcc7HRdl/yq
YplmhmJ8nj4Iqjp/XN8zex5BtLYL35/SCzD0KbHUTc6yJqleXLf+tcLv7TWONhIQ
M161HDdMzQFf0tGDPs720sk5LUYjvbimT+aSDMEYaSiyWYj4SwxghegTfbGw4IwO
C9wM34RUQBvBoQ1ogp5+9zFXJ1cf6cZPunlHk69jwGsIzKSAE3l8GPTeDRkeDmCF
czRvihg2IbablPOWwDJicn+Qv1brkaDqwsrPmzLjib8fNUhP3SYUuqTZGmK9YZdm
R3b7a7B5Z5TQ7f+cfVv4hnIOlVgfP3cnqF1+Kc9LtUEPDG8fIBXpmxgfO8jPBUYo
nMIkl8Octtej1fFG8liWRBMkaUYZ01nHLwNHE7H5YDn77UWMDBGgwsO9+Wpb4Xqh
i0GoqwhKcU5QeSheRs2OJTjLFnlHUBufgAP3PKKv90V+ClilrPUR4h/FGmAttizG
RsAbJVyVBNO/E6jTrTp2D/UU/Gy5f2gxdcQgLPdE9/D98KfqSDAQ3ogSI1nHfMBB
HgEZ69z0c7J1Ku5M6yirroBbM9QfViv7D3ZMbZpWsCMWd5pq9ZpkJIYnRuBAYoD0
lFR2SJtMRmr6LYFYF1DTfZD6lIU7FWuY/rEGJB0/+ovdeqI18aaQrf/0XJCzvlFF
UjmGLkfgIlKvUeCqkFse9Ll5PpvCXu09hhPwx9VHGvzc1y+0BQxkstKYBnA9KsuQ
79NxfNos111JNF6ciB/fvk7bip9pbUONJxdx08YmSQ/DLd/IUGH55n5oji0m7tuo
Lq9XW3ptiR/dm0XxkJmLaOgh4kMg48aasTqQxLKH007tLVsRNsYPk6stjpft4JGR
UnNyNOUO872lkvSc4PrI+wkUD57xjixLvDeomdFDH9QAd6zLJSFrRAydluNZGTn4
btUnvO+Ovy3+LejPdjeX93acZwj1PNpBQT/S/heyedloPFAzgPwwy9nw2Wj61kSD
3S91aiMnIJ4cFtzXfiQnjZ7MU/hnCm/qNobjTvfETBb7TCEB/qZ5YXlpFuW1RDWa
lnp5/AGUGWYrzm7u7HMydHun2M/l6m9EumYHHFls8DR1nKZ/Y8OiqDHXfdjBjeED
O6vNIkG7iPmsv9myvSuu8Hm74eaVg6kEeeHXJTxcZkhdIsjk6NdMjsz9D1gzAGMp
VNhrH36JKOUZAKxFdBKWjs7Sy0T3xusiUd45SGca6fSl8NM2q6Gg+z8Si7JcmaRG
CYxbu3s7kTB9jEVrh68SOA==
`protect END_PROTECTED
