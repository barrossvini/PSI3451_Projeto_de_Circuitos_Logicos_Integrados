`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UvHKw3yT8YicjPc77LeJlN8PagF97r0zMolc4JU7xJqYbGge/AjuVDclelLDt0l5
zmXs5XPVf0ELm1t9aXRnFMUs5eI8YQBOA6TVNogmQGGBntXcL4SacymRnlnwuxoL
Jgs759yhogbZYEQTWiD/EkS9OEoSEsz/GDH9AMM5plos1rzCL+N3c7oM68QwlnpT
s/6Cq2CxpDxVgyo/L9ii2bxqVY0tLQPcNylhBeKv4OlLTDrrNtrMUtzFzQIgS+2e
Kjn3cabTnyeuk5bZPeymse0pj4JxzndhVHbXoeSgqzZpotuAqvS5RfLAxllgMzQV
5U2FkaQzJZnZKXYgWtecWIVegY3hXt7sCaDoMLSbaEAQ6TAPhyzMWM5LQ1Z8uqt/
/CqkBC7jkIsNTV7ZybJJdqF+5DRllgYygKq69BdIfaukkKOPgqBZOb/nfru+UHYi
fHPonIJo4yCySktYY0RGzDvVkoW+lXiruD/Eev0K4vhqXNkcCosEw7fkwODlD8wQ
DrR7PuTKq28HnxY0D/VgfctzGTay5iE4HnL8fJ7kUOsl8magVJX4B5ekRt18XU0c
uj8LbdCyqG1sByjKZV2aL5A02Dwey7Gif/2xGXu9bbBLc/pbR81Lm6JKkBX5uMiE
p87iU/5pkRHwqpOuLprykuAYxczzH9QWoYd2Ph3bCHgITU0/lK9cvLPb/q1J7tCT
c0NrWV5ZppEGgTzbEvUUUmip6fP4VbeIdJH87p01ikzgICqC7Jc6iziSKMAMi8Oa
HQmiQLxUdD/E7wo6KSPU3pOOzkNJVb5p280yDOPP9tQHdrrZ8DxU35b0GHc8OVhk
HPzfcfkCtXAXstXGSgIEzDXK+sqUcfcl63zu9DBs4y1FjusKi3sxaDvPB2bcXUOt
jZJLWzEfaQYAJLHq5u8UclGRQRm+gFC0BXfHGW3tP70ZOcsCei5RMwFGaXYPgoJb
y/jFTwuyMk9Dd27iRjILwhJP/iYjUfJ7yUPSAbNE4DCzqSj1ALR/yiFuiLNsEh5k
EsYMD0f/VqJznZBHZys4bJh8tJ92rRtENxZjho+7OjuANNA4dqIaAwX8V5MJLgkc
feuGGV4Ro2whvZiLt1Su6BfdOaiFih1n5BdfdvvYOqPU+h4I1EzKQwq7vclm1mNw
BWWW4Qpct4cBNMyU2v+JDtz4K4STD+x8kuOZWqITErAEV6egC8/Ug/2HIRxG/ZmX
r9xDM+Xs+tQPIJrGariMNw==
`protect END_PROTECTED
