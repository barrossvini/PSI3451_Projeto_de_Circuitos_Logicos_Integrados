`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZqkMZgGnL1ViSIuA9lY9N7x8dauezweI8zGrHOSliF1yg3ce+MbZp5AUf9Gm7He
DYD2HlmQ2ifvMDz1bdzs7HXnSjw7C23SMwe60MSZkWI28Uc1nTncxG8wVDpHLrHY
yMkN3W7LIK4Jkq93i3COrk668pBkE6KXE21EeUj+ALMGuR6qihQdqMYyLSnpqN0Z
NfE+8txjtX16SFINDC4A4Bwuzbw9vhsHNhbaqZME6s94IdjhO9a0uIqIkQwrSaMQ
IBBwt6uD2gc2Lo7Upj+H/tjZPGFyDJYSbKiXkqX+XfuZI8E+igksHMfOrPukztuN
pB4OkSuuUxJmX89tdbblqhdjBBzc2eyab4KzAd6aM7g9MwBHBkERXn92WWF7Qn4d
zFfBRCtHma7DAg+Gu9gyjEF2KDIZyFIcU60YL8PHzUTXlQcJxUW63r7mwAu8tR77
6Bf72E2zisGpaMRmm6ktHuFgsHMHQp5G1+iEDgMLStbkBGbFO4VeJ5WdJ3JUhW52
En/h87S+9xo9aJ4bMWlYuboU/DEll/lox6+2+7AGXC+4Mb9WuHD/ZzcBA8vkDjVs
XEs3rvOxaOFrskBJrxS9lGyVwbEl6+hftK6+6ZU4yrubz5WGOWlnflywUTR2t0Hi
CRHDcDhq3rBA3ZUB3+89766mhpUCVeh3BnLz5T34S04/ODHUrcK/j+EQZ5MpQaIu
/eVP07DAhm56oZ6aGHgiUHtB/ZJH84RZYX+mqnVn8zfIiNEr8p3GE2E4KBiowdte
zkFUNKnHH+cb6epwSCwyzpTAXTiBFydCsJ/UiX3eX8nQkQZ4lsPn/lmY729ebhPC
ZIUBytsnyMZoLTjc4WSA0nxaLC8CT60bXdINGRjYakDZbc1KcGIb80OTsAjQHPYG
MUx0e2rnqSYyTSAiPSN6OzROnB/GPLjypgIodCowIBLAOTEKEMaqnlYmb7MRmZbY
RiUW838uoNb1M7yNGT/l/69akvMZ7hUDBwkfg8QJ4UiWP4NQVKF7hSvUkKfUXSuT
ApQwtco6gs/5356hObd3I4geyFQALUfZW0633VpGkoShu648et0ZazFdeNRVzYmd
36yOgxlOFQ1e+ZKQZjCYc67LIz5kxmTxpk546/GQOb1HDDio/DAf6UQcFaZ4DI7t
HReCjNbBeTDkZhLjB6ac1suo+aPDFEuz83yQNa4Wots2PWdXV8/aIw4cEFTQxqDr
24u6JcyDQS7f4seAFVL9fB+RupY/i/os3LF7PqeoOMFP4kHOIs9TWfxwXDVtc2Gz
p2Uf7I4CRo/o57cHf4WEB4xVrUAjbRIpqVnF3Cxayh7EnPlmL843TJEnz1VziHnW
4ymjCv97NWKLMaFQJusnrgZnzRKV3kD+K5G0iz+1XXG1zac4DYJg2JWK5Ll4DuJs
VYaS5ZVJrqolvL1qrASvER/tReRXgozhYCsB1kYIytAP4UeHEQB9PPwQ9Ynvrx4B
oKNQ3q5qAU3v1V5twaNtxQ==
`protect END_PROTECTED
