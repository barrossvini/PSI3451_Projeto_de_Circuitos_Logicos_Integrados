`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KC7Mq7iLsm3rAyhs9UiG/ksR9wCa87fXqyjVr+IOow7U1sGzJMASGEOAAYYMrDMu
PsSfK0k/rIit1uZRhnoQM+/+wKASYQHDTMhecJilqN9y0HF+8Z9YC3qTfXK7+m/Q
lkVCvcGq7YfJMGWcpbtRK5NZN27uoRoFLG/YaCqfGNtvrQG8xCjxlAKKKd/vxWRw
TGiXjVUhATqoc0TV2pcE4VkaYyc3pbgiozYVjt1co2ECh2MQcScUggjiqdWKloDu
C130aagZN78fwPRPWwXFQb7wH2Enu/APKP4CFyrKfbgvXZZRYOfNwXvcsi287IPz
kzLmknsZtxDZ/0qtSbV8leMHWxtO5xVM6KaSrL6uwufpEu76hhyvNud9z8wDMVUf
iSOiKbqn7+JGXriICKVTJADLDXfU7h5TJ/jXfkfxToVniFJr3iRnRlFu+PRi8NST
GYojhCAN8G1IUgRvc0ULFJvW1mUXhVzgtoDzQwqP9MnVJsl6EmHzaYcRwBg/gRnq
8PZDt/ne8+hVHHv6gbG73042Pg/pUinsHR3AX71bLU3vMOpoiuIDXEP4o3LUG1qH
50bSRY+hfxb3U6Q0Z4bF1qu67wuEBd3FSNCcqrSG9VVWqiRvZuOHh0J0VZ/uH/Jq
NfUX0sRuCjRpVd/J/f0nKjrncZMMFg8CJD74snH5VQb4G5RvVJr2FMUc3xOBJ8U9
Ju5BcGc0BBXPyuKw66WWmr+m6KzhcE4szLzYEdPn+35BfXPDDRActrBK7ROrEsGC
5xlTHWXAeV0lE3v6sIhKeK/lLdgfu4OP3THG/VV2sZeNViMmVJf1sqrpFfP8Xsm1
zpWehuVxtRtH3HCnTLuhEGoa+hKVwDu7iASkMKMfkrj8lDcDpbRA7XijBOhzyGO3
ixieYjUhLSilKFtRK+UElrI+65CaEl1wzyrx5RF3m2iJ4DaP1sjacb6CyMUfQ01W
ZSy2BbEbAOT5EeabbO0tkBEFrF/lIJYzJVA8NIGyabbHQBXvSnLuv5E8Y1iCA8fO
d12HWdkOHiZvqE0eT1IusSdcx14h/aCwCBWjdWRjCrPbiDCOnKQ60FN/29fmnXqN
S0fqz75UXmtIIXq8ZxmhWNQHhPvCexisj/wR6Gam3k7UZglDg6hYp2YMop39dNUv
QXJ8ypDk6vWDU/zeA+aGP1x7kIF67mO9vO38PX+HYNW9mKmh5/nWkPLOx0IYP+z8
3RSwQe3HrgfHYXgkSSpqNwJjHZffoZ24V9SMzv7eLqp1c2MeDqp6vMlWV2FC/RA8
hja8w0GMPxyZAjEID1I6X3aDcx9YoqT32UD+262RLkNZ3KgJ44riNky6HmomFu8S
9gEl6ICcpgcXXhAjUWdTyAjztCkyvY1BV0XARnNHUectDPBqUfAh3r0XhJYMzD/8
9QAwLhad+tPkpE0/L91yqwdS25vtD5kxQu80Y61KqPo4mKIv39xwxWezeBkK0QZa
De+1NyAp8vfAUxmzYHhYDZgz4aQBgwE6YLyfnUfx+P3ygKdWEj7eHC3/kIlWocXD
slCiDzcujFytgSdaX5JuNnLM6gUyExuu/zqU9P8j0e4T12Q6cdkwDhYMbLJ8SZMH
VnbkjJ4shC6Wcwjs7V4C1bllLXQYBGueMXjwU9pOsDs=
`protect END_PROTECTED
