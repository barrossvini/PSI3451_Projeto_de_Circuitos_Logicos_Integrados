`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLWrpEAxfdMncogiD2G/rHfd1BhkEjfY3/ZpL15AUxHflyB2FbZaKRFbxRgbXa1k
x0IiJWx4YmrQ1ZQ+b0o9wVVIVUm90PvbVD8sPj9IO/YssPCatxyjBYSQ4oT3ro9/
b0u406DKnUnH4oKU7tYhqEMOnbP00+wM47RHzbFNE1gvF3A7rU0Onl5KKGI1AXBd
ja882mNO2Wguf+jcHU1rr3yibHj5trnu6BxZ7jITSiSJxIjKf0p7XcHq85eev4VM
+TbVMZENMpnmk3g93fvkR/glX8XnIDH15Ih3QFnaI3JcbDgofvCaoB8VU++uXN6E
G80qfKV4Nm4TJrzd8pYM3UqJstf9N6TDjQVmsvRqZQaApw4OIJQVamBgIAJzTVn3
QvYRQ+qKWF+km8ybW5h+QWy6dQ0APNakus8WwOhcJTNJ5FaI9hVUp64lAt+UumYl
jZoELza/Xq1UMi0J6CKPZA==
`protect END_PROTECTED
