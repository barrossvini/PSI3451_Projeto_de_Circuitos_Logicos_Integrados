`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6C5vAKRDnj/QVdlyENiWa27a8pacGyIM5AQgDrJAsDU/bgRCfJhqkATNIQmA5ppv
ZrZRiKvKTHSsno9jl3f4KJlV1EaXOEmKZmFLID3lar3o5Aw4UOY1dSTqZQFyQoLo
W8l9bhn32TSygRSf2u7bENYK4nBdxF7i9xCVENF1gCeEv3cubvo+07CBhebAKES0
3LltuNemNsQunGKn5DSH4vj4HtUJFiPwtuLiNHS9tBVhnv41RZu8a1PTKQ4oa03d
0Pp9PMkgLwF6pZfLmwmt+kJ4W7F/ehfAhv/BW5atZAKSosiVFDdv0jA2xKlmIjSW
WeZAeNqtreX5ml5VW5teLH/Xm3EEtdt5KsmRJt2nAAyhN4Ofy8HJu50ohAECeO0/
3qGurcEXIacyCMgITD63oLshQLuQkifSTkgIe8m7rNz1Qi7J0ayirjtt5QIUpADQ
w8CFiqqeLVaJXYLlYGKXcWuqBISlXJDJLKc+k4XiSDq1/6fkIKV9MXn2yVU8ADX/
7YUs6w/hIYrCOCRu/B5fAibM0FD9v+ptACf7EW+E7yl3vUVs0Xmr6s24DXQUczVN
OTyxLm6s1ZVoMs17q+GCug==
`protect END_PROTECTED
