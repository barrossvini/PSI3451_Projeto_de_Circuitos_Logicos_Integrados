`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
72nQ5Uv9kziYKTiKle3e0Y/MO170vKNHBPmClnR9S1SgKcjh8iRtAWtI6iFa9YUL
XlYNIH/KKbszgkumMAG5qXY/czagCJMtB7F99Bm7bguKkK+6hNUsSDYKY2kx0m4m
3Q20ahtyE/GI+0Evr29ju64Ot8LiPO+j64DqFqmOYgRVfBcZarPPG9/TwuFjBjsh
uQALLL7bgQFdcXcnbUCwKer8R1nBv8W/E55vsvmgrF26rYpayUcZXSLcDpD3f973
G+Cezgci+CyVF9cH461lzgRF9XN/gnWsPMa1tJXoWpdmFoYcGCFUYhAXx6ouOqNS
YbhZGbmMfEE/hSHLUBcNLTMx+3M/CQbRncZJawlfx/6Nh9KM42oaxkLHRVglo4Xs
EL5PN2CGsVDG9YFxL7OcAqeOpw7f0SJXdZfGXOtw3TyePpdTP2TtYeMiqAUWPYS9
jvGDMXAJJ7S3ch8DQShl7xqLOL9PutsxDlAD3hgi76K+UcDyPJu54Y3HW+S+1+dx
xn4r/AVZuxdtE1K3ODvJLc8LDb7OyBOjdApXMVZP5L85RvXUz+lNZgOZ7N1H7R6n
UvvQ/nriQOwqFpvZmL/N1iplQ9JpwhyrgIwpykuwqphLwm5QlOwPL80Ar03oiyvU
ArlFPYdWaenurwpAfevNgdBy0Zxx7V2hv61GIOx4izQCqKMVSCGy2LUgGsOFo09X
qzeQqSmGzskU5ytZE3TDYRc2EWjBLbK49F7rLOQMxHbu1CwFDNVkwmNY5jv1UoaB
91/x3pbK+nCOnVp3QVN91iX5vHKDSGrR1ZfJ06fXNmmVgahBCgRnKAHTYf0Bx708
VbTwJXIB9SyHJGtiMbxKltYjKnNMqD1oUHtN8Z5jwIpIybWFS86mTi1OQteIEEu+
ZzmU39E49Ipe87dvaCKeAyOckiqmsHzxcQS+I+joJCMo/pXWmVVsxehOYyIDSb8M
J2LDtMpX+Nmu+Q9emAMwe/Y22vcCJdK83sjeBrFF8t/Uu3XoRvuFRj1Yvt7jw7CW
oOShAW8l6YObAvoSZWF7lmQVbvMe+EW81Ezw1NVWN5nNONeXbmHjYRRQR6mKDxjL
tRqkFXRoi9HUGK6EGfV78wynwzi1wW8xoXpi4XtzOStjngR9zDBwrbv6FXGIMt1g
TWlkR8mURwMvOAKSPhy59aroOWQFHxcQayCsrunq0O/8Mu24GfNX73MlWBmYqQnV
r2SXjM/p2WcA8kyh9pHZtJIzlAf6SMKHarNdk1AEEHbf+/u9uveezFa8u/iYx9wO
Wpxsw2IPmlu8NvZyVebaDjyDIEWzqnSVuW4KzJUmfgGvAeYTyMolu8csTYG1mRuP
5qU34TBzxjCG0siEeXN4AEz3Hrj9UG1VEY1vp/3ml0v55deELg57n2jCAE0uJP9r
UJkkJtyAwjqy+E2qkaf8dYXUAoJBpQc9Ryw38lporHsCSY8F6qG3T+4fxMJLomY9
wyRRiFIioAHbBXE3NzirooQNdUp1H0CcJKlSjSaxyVjN9v7ZR7b0BVgyOev+DBvH
X69E7LfjWsGhF1M1ZYmB5w0yEz0Ro37pFP8DBwHUdYuLu31a7kWmq/I0dV+WLfhQ
OV95TpNgE/L9I5BCe/dR1uJTCGdUH+qF3co6/zV8vgIBu63tvzEZgSshkMLaeA4L
bZqCOk3SsHyL3AcA2eBLNi3dtY5Y9529y2K7qnJ8K5jlzjEY6lIGJYUjTqkXoQIN
RiHERYm7DJF/8PMjThmEUsHzlGTNlUeR+Tc9SVYC/keKf+2alNJFUt05Na3Y4fw1
17uJ+7pzW8014lVBo9TYE9ZZErFIBMe1ZJsfCH0rMlnxCwDAeZa6Be/LVLYp7iL6
l/hQXX+5rgWI5dVIM4TjtuSB7MSyCFSqgfoH7KFYmv2OZbQy0Lqrn4g8pkSiq7BW
Fw4+VLgLIFktr18XtqQjgm3XMvhy7V0B0+6xU+r3C/fBaSA4EhWm++xgcpJJ5x7+
k/lB1GgXh7dZDi8HucMIIZw1wCKOdyvSC5sdjTni/ItETb4rR5XbKs3kMzkdImWQ
sb52BXTTsJWLK4saYy8ezW4MjRP/RrddSlsNszoloXh14AYbTiQ/9WSS9r686fjy
WY5Sw+mAKUlOb8wRfiWXjWhpvrxInXlW9mTto9fNRRaiw2f92a1/MoA+PxgAYGcm
MrjCTodQ5uJTIdAVMRf7qehCdc9PpqT+3dcOkfkBwJj0S7hVUTj1AOTZNRYtMzab
2X5ZbfYLIELI4eFuXu6n821C2TFHqrjA6rNmw2TXWi3HeBnL4v98SbpxZCNN8SXk
LNbsTM77rhNnXrCjpsmx+6N70cU2bP6E3rQmj+SVy4dYbuy5bkYzCVqck2seo70s
PWwY9GRVuJtYIBRmsPN2zc/13sEtSBMBbFiJB1ArHAnjSITcvcbvFh+jVVoGlizu
OSc6A5cWFaw1jKECJ8/eo8F+nmWswHMJNigiHJFOv20Jr4dVJQsVl9n46tbQbDq6
6scOCGXKtO1xwoNqx26zgP6b3+GLH80f8INGca7mzetfYAsQKNFOAN57MSZVU7+0
SKRn5HEyY+n+owh0s3Ol7lj9+RBCpANMOh2jXkRMhKiipKq0cBYBE8YuG5dsmr7Y
EA+dOrTuL5Hp0GZ2mD5QK22ptJtPFjeeb819ZubCvlb8bdBoAO4c2W1Exzrz1kaC
m5QohYuYeznmL4aCQ7ps3w5c7pggLz0g9rlJZFHzEoravfMkkJHx5nzIJq9bFW60
S1C6qyoKPreV7GScNcDD2LTUcLpxHbLDOOgCdz/4An/0x5QRUOIKRBb3Ipv1T9lw
I23JmTRsePIx30vIcmAPdyX/cxOspuaIIP3aaP1HkZsx1Ua2mBzLOo/DkJTVCpTz
TTjmt6wM/tnrfuSRtKut+ZN1UaBBvN2WSHn5n8zWYtBEv+e1iMqOXDtpKKFcV8kO
XhUqI+lV8eTGorCSOHgrRPhU3XqWh/qX8SrAbvgIBR0cNRxNZVKiJqR95OOXlA92
N48Nd//LsYVCHPA6rC5mkeOJJ3+Dr8YXgAkL20Xf3ZZ2yk8J5aCw+vner26e5nPW
D9CshR5lvGkNcUBXMsUBmVlo2fnAZxti+qVpyu7IdCcFmaGwNPasZUrov1T1Mbug
rki6KNhseKRO+OjHOBsdglkXVMin5s/VYZ0VRYLJJHKdpkqYjUMnHQrqgujsp//4
JDlIx3zJBgo0mzYjDDyecQg1JdFKspiVXspTMHrv66pWIxjMVQGPjs7hP63PkYhu
RJ6wQBw7QdjPYgIHdlu9jpHqtKetxH17Ya8k+2KcwGejQQ3P56zDH6jQmIdBZMSS
EhKKBrjO3QainWY0qaG87R2OxtBcTQJf1WDzzg9uRx3DoIh1hvshhZVZ7v6Jz5eg
4PUP68/cubgvovaElpNBZ71Lo0BfeXbldbEGdnph6YJWq00wpZp3ITK2iPMgJM8o
uYQZ1EXKfdh384OQljIeENKS4PsckOTVHi2US7xQuU7NTcvNc3Y9PlejI9Kl2PrC
WwYP+xiFZULrc8CLndT5qZi5XurVUBr7r5AXzwuK8yXgKRgg93tdlH/68SbKWagr
igiBbi4OKfJedd9FF6xyB2MLVlzMXzC12hGhQ1SvFnzhJWn8Cg4fHazjVvY1sj6W
toNyLxXeFV7lZJnSwl97Ir41tJVGW/dG39BXMoPrUks9XrocODA5jIo/LHm++5zm
PQFshD6mgoAWxKhbnBQmixm07BcoW4Eo7pa1JxgQx4l+aiGacY6J+DoXazj4yVU3
pQS1YKh6TLuSG3lmXpNOBmAoSvAndzfKhk/jL5X0eyqIDWXR0yQgnzFk8dIoka4i
lX4SCgPH+j8EMxuH89GHRG1mGOnOyXFDEShmwbHA+hzmVD4IWIAdCwgjTB8YmRP2
F/Blae4V0ERdOcE4PgGQRy3I70oz4lTIJ3S4GRTpGuswIh53JQtZOZmhs13gEFKx
k1Y/rPPjLoycvyDlDPwVr+AOEsw/3h8dO8hxSpZWBb/VVhTedOUGCKER07+CYM4X
d6bUOm/opEbJqCu1Ym1PydAshG4gIVqx6Cf7hbiriXryenrFj0eDTllpamHwwVl9
s4ldEW+YAbgtn22GHp2qzVkfiDcTotLQcf4+5hnimgvb4p3+KwKsc8e2lenOezqD
et7sTVCMy20sGszYglz/QBHUn57ep9yk5UJJXgyAN2u5BSlxdVyRZWelzqn7XpnG
kgDCves1Imv7aAgiyLO1UXXL10EL32l3ljdUHwetvBc+RQRLNVBKJEebQ1f7vQxn
+U6MtcanZb1s/mflgK6qOvp4e16nbN5/aJMVwcvvf/6uRXUS5oDN5mfCi/3Tmcm6
iDiXtfNTiQXmP6Ngy6kqu36Ap21j0Oeh+TVCmnCd7zd75IMGktJJrSEv/TH9kZ4R
xhnC44yLDtGdOu3zfjYT8RoPAZfH4z9KJCQ5DLIWrZHmCZAFpcevnSsvG7mYjFbD
V2xkUIe6wUFWrV2iBnxbRZ7yTF44EeZQfwxdBkaN6czyjjKdxL99xWSuJBg4ldED
cMcO6jumuWFS2eU6RaXzqKvGh0cwTJojJiaksKVBkYIe5dnuYbOx+d032S0SXn1K
RVjSFYLFdhNr/5J2/TJHuOhi5j2OHie+1uhHhcSE/kHl8CuKijDoF5yxsXpyc/SJ
MHFFvQ+rvM5OtSHZV/KSB4tMJKj1nd0Y2qTO9JCC5htI2ZmPShPlJgVzM4LX5t9Q
E5cRS9o1VkGFymZXMEq2EfqpaVoJUWAMxWNC/CNZjBJdnKal5f0DwuMBjcwnPy7u
FDkbQ+bdbmc1bDaDvVqKiXukjIic0ospxJUTGan5jAeEGAtYv1PVdGuQRkQxaq29
z42R0s8cLaTgdW2gVrt93J/AchmLnxSH1v5FEdK+EwECYvY2YGVwduHHE7wh1RiT
HWYRZQi7mTWeUidSmaHaXdoa+tW/COwQHlhnySo3OvrgZ4h/Dx8lAa7Qr+vUq+M9
ssribzYQo2eiM49/98t/cPCPifsMvq/p9tYHZRcaygjqzMTG0kN1N/qsJ6Xf+zB4
V/1EUD8HrEKEiP3DATWcbCUpyzy29zIF9Pv2w3ifcwvs78ddHQYfsb8FSbLgR35k
yv4mwZn3Fno9OMHNopVUcQSGAigUgl/4FdLw49Jmn+uYPC0hpAqO5imsYusW252V
bHUz01qbXwmWgb9v5lmsyu1uCo0MxKH7H+bs+djTUGFkSZWequILpzfoeEmoWQWe
Z2zIWjnB51768aHBXP9gUgYtTeVWdToWzBNMjCak4067D6ViGMx0Bc4UMhUfkFXe
GIp2aalDt7BhsnfZz+0UFVuKv0/ksQBbNYyxxdbLd5AVmMfgGApR6b8hkldx0z7+
U+bLqa490yXrqo90hQyGXWymVJHP2lekdOKPPDcb9f0wxlzGhOnyPYxAuAAgkIij
l6khf670cjcCpAFFT8+ZaSdBsicDZKofztfJXbpEKJUrN7HeEAm8jxMA0LfzXVQC
T2GVSEhgnzABeN1iQpmKFUNHSTh6scZVg1xNSpZqVyJDoxSHHYUXuyHVFQwaJVkx
JONcjbeQf/B/MDOxcMKRi8N1D8zbWYupxpdAG8IbLh8n+3u+nLaBmanhpOEzOp6w
Fszpff5fKzbnc9Wv5ICUn2lqvLBY3spSNIVWAxH5YSC3AvbUacPICZgjfIeG+4Rd
Usy85CSDsuQiXXZBvRD4TJN5rrN6dybVS5nvBHy5mrMtwu+VdIsrxxVVf1kjbcSI
UTsgVeas65QGaKlPuuig6QW7nwPH8GywvwojdoyCPuDxVg2/c9+69c3IvGonpB7g
i21bRkShBNU6tanrTPodqZoLYOfqERdyDDATRTz8rOscoaCJ59YaCQxVdkUx1WiS
73DVwTdeGC5h4P/t62GahGSAP8NvG+gkXjm9ApdCzsEiyg/VvN6yAtXOCBdGl76E
t87klW/JN2c/n5kD/VjJSyk/PPbH9MlE9IzU2TRe7VbIa92h5uw/AX5/5QHGktDK
08Io5UvolsERjzYX0Uox1FkK65Msn/vkvxgaqXmM5+aM6aG3rReCKWGMbKZQAUaS
IyQhNxo+aJH9CaXS7LexUCcXvmQL4X4J07faMC/XpYLhOvC6iRn5bZw2VI7I9HnG
++JpoMQ0EjX9uljxpcwobbu/xYHlGVouBPLzk+02EBoOZ4sQKrzuQuKmXOY2Rwlk
yMZbV4T1AT7FC0xmVZpELFXn4A6IBBRGGuKj1qRVboBi24yQVRplYPhBMHcT6gpp
VBGAtLslBCMSkENwYYvkzBaKm6LNNYvySY4yGIXhTh+V5ei+PzUOo4LSiiWovBJq
bxtf8HqjYAtXKLJtWFH+N8Rg40WSTUbpe8VYsenHHIGX4Nsc7ws07GpfSI+CGcnZ
owvx8eJoiBdz8T45B7vXbhxjs8NVW2eF/o9WQCGS27wQWhXKGeWlotaL7RVmPB2F
aWmxjiitYR5OFaUuNemffjqBwxBuScEmYt527+zWQ/Zy8d9rJ1O9Rj+ccHjWmA5X
Ap1Bq/70r+qbsO2W/98fMuTNpro8rByiuWE8b5RW39MWWiTB+zUw0Zi07QVeUTiI
s2QBRyZi7CwPyiQPhMVeksm49uGLK6YzJlIHYByhSjNl5QZ26d+0mArPFJLNIeis
W5SWjX3PI/cAElkPIo2D+SemFtYKs+4PHiM/kJoRRcR6VuxwcpGcuEunNKeYN+jH
oYUYnJMw7vNo+zmRKUsLBQzs9gZf9rPCz89oO98XgYmVjlf55oyh+OMAd/DwOczQ
qt5oUI5YVbC3alCo4HOpGSOkZX1o7TWpCOki11H5aIGzwe7dxlnlruM+E01kaosp
BYX5lCTFviTmhKK9KUpPgunIZNHMiIy53jLYY1BJln1QK8j9XQl9xP5v20SfB7LV
1n6WEKOLW+NPUi3BayEhx0quQEGRpMbY7aWzTEZQGfVvqMsI30KIjaDo7Ma0a0ts
d+SE5F5Yy8sAIBXdd75v9gg3nHnHeL31ozuJ4BHcRoMWNuwdOjVU/2Xk6zenOM+6
WeKjoXh1PwP59gW8semxvSTXlH2p2B0KgGf+qrka5CQ+Kb6DwN1XmAxVqrtnslla
9Sxnps0OE12VlxfaiAlSRO5ui7w0ElaJjS6Ma5LYWGcqtlW4JKLW8X+IpqHSkKNC
pU1YLXO5YT9KSRbO/lSHm1glclXXwhA4QUh1QmKEgouJ6LM6Zene9nKA3tr9DxlY
C62hLeVoPLDBxi9BBn7iBSWh+edtM3RVYLuXTll12u+sbwTBwdQrOPAVmElr74+X
b70pD8wjrWX1QtPMEj6YkDz83j3mHRv1NOcELHKhlDpj2SXG51jDScFoQXqZsfnH
MoG3DJie63QhNR12wKpYOCmTS6RYNgIBTh4wA//sDhTCAbkU9IqX7bJ6UKdDjwcn
jO1Rh7iD+k7pvPE5/lL6SgO5dTqj14VwO5iNqe+lQtq/GNgNYF7s9+0ISN+gMSyg
nhKSvykQU8Uw5j9BX7vWemUUHTNVune1z9+ogHShf/6vvgteu5VpN53qjRAZnwTF
8Jgcg682DhV+l5CRiUSQ9RZsQuY71rfXPSs+SFUN+21fx1U5xG9IbZwCj/kPpSK7
5MZ6rjZ23/W4ZF7bUb7nLYv3WOkved274QhhPNz4gSo0H8S5KZ6gqLbi9qu4tkjT
aiBZHnQo3YkQ7D3s4boa4Zv+EYhjbWpM3YTidUlMizabW8NQx2mbTT8k9hyASALd
iI2Mw/ZKGPuYCls9Q1hU5WLZckxepYqO/ItUu4YrPvCw/jygH9Brni/QYPiNItb9
cfp+shAylrVEoF+n7HLgbaL1Nr1dEYUSTurVNyoOF8eEwAZld3zf9fmZSKGSU4SO
i2QCykB1m9LBbK4PKNbmrhWfSq3v7Oe44Y+BZxM/249IgwIr0bG1J2Z6R1swUKAC
5dFs84KyLvvAQs8/q7VfMv7IZbY1IxMInsuUKVN14l9o3f4PLcymeken6Mun1zqr
jREuc6LLmjCPz9e6YaKhTT5mY26XrgImeekC50XHdkiODWl5izaqrQZp3sbGFiHX
4FmP0kr7T37a488OH0eVakbvsYiLwqi4TL+woRxuW3bixaOXFTRHXf+49Qh4fM6w
VQPOuKw2biCKjf+evpTDOExZxvDMuSV14g/UAzW2OkEUwQjD0DnEdFulM2fTiSLK
G1/T7qrywGZL7cw/aAV7kzt6gPbumLktet6//azf9jQRx2w4R+MdqBGEvTR8YH15
4b0skShmSxG+y4jUUkdsPDn1D75UgZfm3faeDZFgAa+KFJJ3rYaJoDonODJIxEll
JzKAHvq4lW8HrGPZlL+Rz1ulT9bGq5JS+wO6s4m6yVtgIpGVWpF6tpbGB8Igc4kX
4+4Kpl+5ny//n3KCyalal6dbbA8isxxyJYmaO7LUBD9zmSh63Q61PUwVjDbEddum
qggV2atEqZpHbiUGvABS6CnXlAmCqunwUOPEBbIhnuVv7wwghJubF6xGIXWdwFHd
QEGxYNeKVWnUNNXsmwo39Rnj+mjGTjNozy11321cVCEEGn+sN0tDiKvejRNgZ7pU
vE92EjiLAFh3BCYLsY6Hx4pIy9/5pKn8VlyBd5dcsH3UdSlAmIx75tZFo3UDzzLf
eUsj7EBFOPtfDhu/MCAwYxjBx9mf2ChG8CNWLLMlQdbgiWo1TlTz07+ox55t0TgW
9bM9c5lzVK9tfuGJjlxQ4d5JPvkvWLMDIWY9msJ8Me2BcFkYHcTRueAR0cI2IYvy
5apSRFhtMW4ZEIRI9Hax7p2Pq5lNDGUGH18PgEouNxEAK8mBe58uvoA2glhGSMLi
4pOdIhVNs9s5EtLhqBLc7fEGYp4fmg6maMdHyeaCJoSRAMi+oFT1QPQIm+GSMfWg
Bq2QvBfMB/7wOo+P4IyFyTVk8nanf06j4hTRiBKJO2UkQ8BMqpaExTx1xkFqpkCr
Yc2tGNyZxznbEX1kbat1Rdyq8PVwncJx/ggDnVH6xSyVHTpXbDugLoRy6e+Qvn55
GUtx9JxLIXtNUCuz5b+v/62X1tdLQnDk0/BnLVTp/AgYvcpcvZnkx5q6PjUGK9al
i16BZS4lXjde8GDCL98G5n33HdLTraWsScNVRxUFWF62dYg4pUXlhn9d8HPPlSzc
fnExHOyMf8Hxlp1nsU0Y4en6mvFzHEc9feorg9/LHlAGpgpiylDmb1hoHpy2BOjl
OZEQnt5u4zvxIfJWnQHuruVVt6m6JP0trtOJKf7Tw/xpbm7rZJ8s66jw3MCLs833
+Y/UgTOGXSiaMSkM6UBRYST459//agv8s9LEUvCafWkmgw74lqSiYz9AZNNN7mSl
gxcUU/m/P/24Vb59F/+X9HK0s8YAW4KHFlJCCIpuoz8hvgn2MkacRZ4Y4s6U6wT5
F+TnXyIneav/zjt1dhcyYoZoXcqaNQSFNGKvlqNennao8eTNE65KFLCUrP4ZRVxh
wtVCucDMjrnTurPeghy8K3YoBW1eAmGFbwgJjwMiGLODnTugyP+vo+o5LfOr5ReC
FbGbUE2N9843eKfa+sZAVJ3i5pjyAfuXXKs/TQ3Ye4Vy/8FdGR7FVhZRLXaRRNU7
KrLtqqMwE2PQLghMhQbhJGFhzYG7bnJu0HpIvdUtmlrLGHG+lWSgF8JQdoHidKPh
LJBWK3ZzAO36d3rJN2fPvVsG+WL5QpHoaqODkgb0JM3gcbCTilxonhSimasuBW+M
31+EjojXAsCsopBKsW4+TTml20/IOxP7jFB5BtTqq6bwuRGrUKQBlx9p31I7kkNv
V112Ca8xNprndQStnO9gSo2QDhZURiBpi3jx73KXOTEYLdI0OcjFo3lcOBEXQrf1
MLkoUWtkIMZhV2zXdLrs5BUCHNYMXluTLDq8/6/EpY9TEVRuey3Tos6j55fCa7Vi
Qqlnj8GFLiIZszBJ2IlqJ4oO7qr3H34Oc7oikllPcIN8w3lw2PKokbvmE34uYNp+
bCLD765zNQCGWOxw2c1bWxQeyExhKcOnmV5r7UFmvxTZO4N9ZMKPPY7Gf4j2wcFM
RDPHqS7/LmPaZHVBQh95Ea/SDCrQb2Lvb6NvGHu8wlPn5femBExPaA3rFE7JQgC2
1V0GW3EOqRfmH6CK/ZKdMJls2aZRFFz0msYjMPiBX91lAO9GM37Z1z/7j3QZpPZN
K/lGpwCS1r4tRhEsz8fArcoa8GQ508nfE5aFaYb5EUxL5EQI4nkXyICYJgojKetF
Sok6ai4A5AFh84JlhYqXCJXAKOYFq3EBCP6MdEY8ypQBAmtXTKgseKcrr2qOMTjI
NjfY94vw0Zog7nxyDHkwOOD+Vx5y6i9RTrXQQaqQ0ZHUAa5sXrXO8hKzS8uYfXc8
ZUhJPTzHngwBMSFm0Y0Ggam1uipB4dM2hOClWZ50g7sT0E9EnbzWHlZqxSalufUR
3mHdONqbbZbZ3RcCJWg89HJj3klSos8X8U7TipxxN9/ffW6zOqGd+9I1GGr8uIWd
FweorxxLjBHfigwMLF61Ogm1PkY0T5r8WIZeU7+18dMCcKjDrcnDDljfom7U2Ek/
hPPrcTdi0Sl+6ZDSbQh0PORYlRMRqsCR9BVSxesOPLAKsfN4Vnn7lx8e4PuV59P+
Z0TVvgUSEanuMqw7Fnnda9izRpUvwnqZiVubu2poSfmFp//LLcs6+8zzvR8YCecB
93F1oouWx+JDTqpiYUh3Xufpl/5+iUvm3tjvPJ3WKDYpD2Jov5Uhd4vVbD31meWo
xxvINAOO407esOQFwcTqMb+tjkM7c/nZ7EmVGZIDAsSLz48bGMbPQhkNtn2zEaVG
rBg0VWfFmnXhDUkC4lo3ax/RUvNSt8fA63rIIkb6+31Vz5VTchdz7RkVIVru3gzX
i6uv9YOulv/7QHudZsgfCRG9RlEBCrTidtCwzPOJf3I=
`protect END_PROTECTED
