`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3L7ZN5l5uF0c7hx6ejAw5uaH1rnGd0cPLd3m8Fvey1Z2xx1Q+NeJEgW+6EVunovT
BGv6ZQqL02Lcrfwo1/BjvvNTw2jS1Whq+UaBNQcYaPmsrKOsAsSfyowSywn6NzVx
7Tr66h0/MgZ+ue8fj3XsuZ37CIUHBBj4w3iNozsHdTTdYtl6KjzkPpkx2kRGSjST
H53vJejjaEb8vuEoZK3vnw7WXh/QZRfOXlEMJ424JpM3icsd0KyzXu+9xl2Ca8pI
FfeE2U8+Qw38JTSQ94cfRmR9KxNuc8TRbEFXfvL1mSh0YN7M1RVGFD7+ui4ihpAn
HTFkY5peH5rC+xaU1FD4fHoN9Wm7xPoMp4Jyj9on1Wc3yxwgCnRr75gjjzVV4FLH
jH+m3XkBejwzErWGkPYt/oRKKaHyP7079gykGA/vamUDSQqMRncQgiuOKZsaUkSE
8uYp0gjbm1Y1sUrNPo7cC9+p2NZj3HTefcQiAwL+8wfffRYUhIT+SkCUtYQ+8x+b
lBL2D+Nwn/OlkNVBSTdthWJ7v1FCLOfa+11wpHpCxxkmPim1AjRuTh2E0JN0pTwZ
/jX9+Mr+GPq2PuxtyMp64F9i1umm/Fnyn6WDbbAbQJzXVlApXWT4t2YbdzyKSW2R
qjdNoUxkh0WHJ9yesHpvqy9n7ctFflkaulovWGnKTMsEbQupJvrwOeoVWvBFFxHv
iy+4P2EbeLX+D05tAcO1qBcFrgimCIN/OC7DWiBSD6QtpR3Of0wbYjNL90YRVwzD
QsKXuhhaduRbmaXS57WTVtEr0F+z80Y9xSmewDdoRpm8wKDLWm9V0xVCBVoowCUr
jUfzbOtaj9lanLoZ8e7iVam7Pju2vFgPYKnNyXQ0c5WCfchOT+c7bjAEzTQGYNJP
5pVX4FS/Qbr55LlJMLjGtkY2k0FB2CNpkSjMnKVHp/YrCNZoCsFzUnZ41Vdv4Ubz
Jiul5n0chyw8QXM9POaLn1dMALeVWKhGPeheD45f3qM5fzNcsQ0W5pxKFlLc4brn
rf1Tlh1SjptEoqWBlgmK0jo/VTkJecNZVR9/Y3DC4sJswW/o8s6JjS97aTwBHp6C
4cnDELd2zKyNkb56twhybVCWhfa4/xaE/F65LOtbqtfzoGx3i4hrp4f1VxEhK9Ww
diQc6kSqop42a1YNWSvnNVpxbL9nR+lX2pcx9eKc8c0ftMQWswYWYHmJ/L2hS4R1
dvM1mFXJQ4Yag5l+zoJ7tiOhsKvMXl0LuSymFQt6WPkyOZCKWYwqAtfLg41BVukq
DxVeTe50M1BSM3IztsWedreewi2EsDIOl4SMlU/Lq+kG079RgAEDB8jF1ycUlaHA
igGnRzo4X++Qve29j4z/CcwZWBK+gqi+93okDhMyA5eEj398azCzdhfn9VvDj9Bf
ritiStlU5+l7VBapOcz/ti9KnLDbwQp0a/Tc8cQnHr7+LxEuoXVSa9tV+37H7x6h
dZ6DmsLJHZ4ks2uekOwjufLUoNgWmcpzScNwdj14oNY=
`protect END_PROTECTED
