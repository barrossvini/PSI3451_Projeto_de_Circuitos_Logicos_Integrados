`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R+SDT+gpFR9mcostdGd0BE0DvUgV8TdIMFyH/96Bu6uWi933PP4ulygI1vwHl3Xe
qVCBNwtTXkdjNh6Z/5swHcGZAyldGOKW0LV1COgJSNsgPrV20P04Y7E14/G7YiCh
UEkmMXsKiaVzsWnKjcI+QKvl4EMmFO0WDIxprfaMcYsYQ6FSMSS7F+bX21/C4rfF
1BEksQcing2fVGP+QZr4gxbr+ehdWMc/pJxBYMwfQURcEU+W5amUHnIWiZ5w4uJh
/bfjc5Hqom7vbL2AtbH1VJqEL+8XsBU3hHe1FzyRkvw0S6pGyLiXWBHwfbaSucRH
tghAbD+ENxT5yISZJV4lwDj0zHmu6qioO3W7ROCJfni+f7lIEz39gCipT0FugC+F
MDvffI4OxC8iNX5UNrld4uo+qQgu0Ze/RDmo39VEkxMLDajofaVj89/IeGk7VK7B
X+CvKnoHD7vGM/0uAQW+yo1attSu+LsYoNE7G+pLERclvSfEl+XM3Zs9ibgYAn9H
8fH3JkkFuTveecLO1n8bJv67iElkriDRNSUR+JK9njJWeZa/XLqRcZK3gqtzT9SG
rf+EONU0E/l8oI+QG/9u2Pszf+QisGAs4SyBeODTmz44wrv93pN8fVEkmaigDJ1p
jGRcFM2Ev33aL0NlQQQWFigBoUqtcS5ExBALvAQAsyvXtMlWhOhWw9HQWwV9dm1P
mYe6jRZabZwyPQ3Cjz71P19Rcm1gawsRPz/Wq664QLC8ZfnaQB0rfdfdIZcHIQI5
ekuPU15NwwCRljpbfL4/ww==
`protect END_PROTECTED
