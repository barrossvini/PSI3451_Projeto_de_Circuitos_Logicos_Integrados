`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gVfuyLxb8XJ76FjFJfDaVh/daZ10TJp1oj0zWASVGOXw/tHw6PvwLlMIAY41/an0
uzK9dAIgNKz4TvtVY0H+YYSd+gXvYmWLmC8oXY6tOw/5eVcswo1F7FzWx0rKsbi0
ggovjITs6/20jmROumSQnJM7laYR20mg2wn9i2LxAYHbPyfuWiCNxbkwQ4bg4b/l
Cl5kF6mgetM/9/dZvro2EooyxhtH++gPzxx8CippB5mIZiN1qm+jsNUDLmQPNKT9
bRdnsRu3DIemrJE6MN+LpfuXsoN5k+/5C7j6izfokzbGthQWLaNqM6+iW6fDdms1
yHdEKs+om33+v3/X2/1NQ0uzDOV7O6PuYjrfP0cyJy7N3M899yEv01MfOTwXF1VP
uCIeLaqxUds3gkEntZvrar5PMaxyUr1ru16P+f3ZgNI+gg6DQEcO2qDJf7hHk6PG
B/wTtwHPzVSlvUdmccHPSNr3tSiScuG20CohfKfTPae2L8mcNGrPiHIgfHqN+ZAC
Oul6mPcUNXmgKspLnsbuE7ocOZwYlDUW1VXAAvnt2cDeYCtKMwAVyke9WQCuLM31
xgaQ0Xyd9QgvzKcLz9IBH65GF7SbHO1y9eTfwGbEJzU9ZnD8huwAerKdZzHeWHG8
yZrnQOAQqakc/MPYmGRbafdhRhdPKAPjT3jpTDUK/RGtmcxgxmiDnp0KsunoyvbH
X8XuQW8nvsECO620+pjiVxFEU65k8xXQSe5U7egmOWfDE3pkwdsfNtylwctb9GVj
HAi6kpvNImfQ3DeXLCPJkWAfBVaXGM8quM17kNlN0597cq4pAv7QODCxt/zW+rDm
XRNwPBYIZ1B1mgTv/YuQ1a2t7ogqlMbMXtykyoWMbazwIhXIcz+N04gCMsehL4hU
`protect END_PROTECTED
