`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qdlhAGAxFErxeNY/HR3oOQCBvETXc519XQgKzPx17nJ7QlxPw6aquCjloI0w/Ck4
57Wm9fl0PwS2xTv9nBhRRhjPdrBmceQ4dNE2UfaywOJjgjEf/l4CYn6ArYsQmycI
NGPg4YYiRw+Gg0t9ORlU589kL7/QzonAhXoqPP036O/ohnsFTRKe9efql+32yUmY
zMMYzKkIc+McmIbQAPxoQmeFZNct4VHso2ooavl8uMRuGFqXNbrqBkRvP7hVeaqk
xmig/kO2TA4D2PxUAGRfQ3rS+dOKCHII2vblDN1s4kj58Qqpt2/eT3ta3CcTYQJk
r7Mv9Sdonp+g3+R7WI9AnvKREyV+j93I77q3+DM/D6XuCuZsh5e079aHpn+Ox18a
OTQUydI9Xs5aKeJhBw11/Mb6G7Dc75RS9XTZHXc7FxPeAWSSbFsnK0SD3teZlfjH
2RgLTERWj4ej71hMYT12Tst7bwiuSTYUazXQHZPz6qhUMNcA0gBxjhVDG4THWNxj
5sadFnw97gAiawSOiDM2/eT+c8IsL/a64dewXHNniJe4qrmc5GvoZHmNePFpKdMk
AZS5Wm6l9nUHtND1AWvXWalg4joLZpRhKng6qW8m/R/hyNM7gMLRXC3Z+S0z45FM
TnXK7FwRMVryEqmkYNdvIwE7OpQSlFOZxK2D8/4m/DTI+7X/eKej08EilM5dJK1z
cca4xSGAviUpy9KpeFklWbB6bwLd5luinwR61XA0SesyxVuTMKEMCKIN8hWulYtV
VfW5SiWximTqSoXWg1YP2agNw58rU8vX638tyhNh4PpV6ERx3TeNbUbp19s9ZBEu
EEkHbHufIJMZpcN5qn112/0r2C9ul8hDQLL8kZU7QYqEJ4KONW1rXIfforYKyeyy
n2GmJJwGYWCw1B1SAa9lN1EwKHigts1tyAjY5/Z2XK3yCBZSYbHHOWfjQlwk8DIm
Lc0y6dyXj0mkibjR2WNfacJnJ8H4W9jEMvIv7n5zEEXU7AMFCcPXQsnWPyxvnFd/
I0cgL6G4bvpgOLOPJXZTOKvlQf09SMVVJLGuZrLprao6+eSY7YO3yHOyQW4OMq5p
Oo0fq9+4R+7/KGs+FREt6dnaZXNJTfjA+2Sb+uZqdDIGuAYVV4MQP/tv5Dxo0d+6
l2ahgaVvbWnUnRxR7CPIWIKckqPnLXh7Pw7PRnQ3xRJHbB09dLeQrW8G3rcU0yyI
Egp1ROfVf5+0WXP85HnTVW/j9a/wLbFbBXobL5wnHAIvgvVCno0xZCnBH9AoD4D3
B3DxytMELGcQ/BJdhXTT25z8kFtFlHdsYH9YtdooZcawWppzKbuBBsyO2S144DZi
74ZBF1wX41nUHdDfxxglU6FzD5lqhZcM/zozmaHvQsheQ4Oy9i0Ve1n//ERE8sIT
Htc8BZakYqE4TxAA9JwibStpzIXrSeIlOR9edbySijqHfzBqHX1vM3t1GluytCg+
STWlmmtRlMe3QfWScTo19kjLsf/S4eifBBObx06PDowYPZzGPq3x6fqKx+puWmVC
RbPnhxpfiDq/9+Jymet05vJ1sqqg5c6prjk1ibUkPI7G0KgwkN11ilJ5IJQ0fZI9
dtBTUymLIfOt5ig9Em9vvqr0c+KKu036TNjnCX+h1tpeehxgzlZkjcsQ4h9RVTP3
Nf62KSU74H4bSL+tIFd8DGp9s6f1kOMpYYla+53GUpT9AR6fOn+50KNl185IxvoA
Q89xgfAd9X/8INQyU+thscqjrD/maB6F3SIwXQANNJvVv6ZpajP/kLLG6iCMRLcc
gw78SzV5NK/YlYr+dLvodaRe4f5beLwWjMjrErrATUK6AJElWGMrJqB/uVn/aHuD
FyZr6L3mgAJOljGla52NjWQVzkPo24a+TJ1nErNaYWsSlvFt+Yib8F1dEgsYIcDN
TPx9GECgXgPRlYa5fWZDtAQJ7Jfg+VYUQWj9CZEdokKrv6McfRCWwFmqCMMF3XkF
TlDHnchuGLpOau8j87/FRhUthmQtG3Bn4AZSV0LXrn+KnRER3CmHFh0qtzLb1d8m
jcYZaK4EiP/E7C0MiA2AkRaCpgFlfRPMRWoT/NwLdZrVy0VVia4BZo0X3sj8qbpB
ej/vs4W9n3ZUSYlgxGIKo2vqZvL7QWEa7B7YfdsP+K6ycY0/foTHGJ7ECZ5DPJaM
ROOmiBE1ENgInFm40oysg5xGNksGcKBug8Vhiu33Ou+GNkejsUiquF14vZ6dviFq
nUFybTpYLUcOYMPlJV59ayqA3ndmp9itDpRblIqLBVpuPRgOTqw0pmL6/2DP+gFP
RyAydBQDCamxHorEDMVyFoPjb6NrGds5T/AwdUbhe4b9vzlQneQTtfi9jA77KAxm
ndVmRg3IIkrFAHZ1GsLlMZpxrQBibq7Hal0ES302Z/a0gAX8dh4Up8rQRraTg2h9
yuQZldhVHIfP3gkrFjR6AG2LzUo0QwAcsbEz6Y4DIqwvEy0+oNVOBH3hKcgYn7L0
NyJEMBiutWIvupi+zIZQ+GROAbmNty0GZbC56lmHdMxEzPO3sMnk8zVlhGZRdB+t
WA8jn6IPToGjY9innuDbu//FgRQCxx14ociEuqnjva6DtCcK14bPxGgoYnXUWbnq
tMJmkiEyNAa9eVmoajR721wcgBfQGcktZVJp/++ZWAqJv0C+WSxd8kMEMda6gs6r
OwDROB+4JnfPYAfIMwDWd0xnjCV56PMPXoy7FbeBuegImVtR7gukSBg/1m53mX13
UPeEbDzpIZd6nj6J5VN3Wr3F3k56os/Xuwxs+yx3KfSzJ8kFamAaeeUUTldvwJK8
bggocORyUVPYES6PUrTAApux6IgDf9PhjyLB/hsWeqNBDsBb1UzS9vgu7bm6/7OL
Z0yE2FMqCTSMYSpu8lfD49p3Qa3MglJMKyw/I0ICR/NzZxO9RlHYtcBVXbVXYt/m
/MKABP6beELliV0LPMzrbyHA09fS+jrHHSasHL9X9Fm6d9VVeAimVcPRS/IEt3wj
XjlAdwHxr8sqGd/CM+uIu7CLbjRvz77VtILGB+QXvFyh6D15ZpUtkb4lOCNtHk+m
v+p3UYDtB1WIkxqcL5neIZPoQ49wm4aHSn8SxGju8pW3n2mWs8YlydIpWajyO1sj
CxI7kwe4GDoZjj8GboJHRHMt6IDVUSfx4sIY2JfL+HrOByOJCBO0z9PBj9rh6xPm
SQUh3qJLZKcVmEqUkgMu2/PxFvwETva+BL8HHao0jol5YJ1rSXQuBLPktfLddhAz
lFMcYaZO/oQs+r4Ujxyc/6HAxhzy5h92DfDBl2xBUZvDEVhnmkyoOcUycl0g20Be
h5TnT7TD3QFCZdCXV9DzojkJs/c5WcKqRGPMAMjIo1xxQzb23FSKun1jorC6XxAl
4MLLd9XP5oOjsjttpPEtlx6FUybD2IkMaixI1uhAzB0i6HylPnqo8l62JAX01vpQ
55bjOcms3Dg6uMv0v+e8OBm28oafrkZku8k17Tld7XkYT7evUY6dAbapYYQhrFKq
x/MgBh7daHYOWhC1Ii5xLM6rc0vgDT3q0b+L5me742ZIXAgG+KXGYQlydqBWbJiQ
8VRrriqoAyU/1+riRfpeK4zfmHDy8nD+0gkNStKEbCjcZ+LZ64XY3uZSMUH1luqo
igfzzaWF65RP5QoTqoaqLAzIxa/PF8f46JNHOdgScbQ8339DUH4e9BmR7BYwU0tU
rtpSmQCnME7L8G//Qxfhmi2wx0lqz6sXLM+ZSv81/xlHwQ8HWdEAH7cJlWR1ngjm
qsOG6lceZqlazT/v14O37I5uNff81wvbBT31gXfkRjbcpHlzSSqEoqUNcZGZsT1G
xQTNCWMXhd6xOLg+jwBqeF2NAMUHbz9wGl5IYi2LxnMFB5kOnyI6K97is2g8Md0r
bhip3JprrOoPifEoi7HOXN9Ovt5yNlqhrlDxCnXhAbKdnDZK+9AkIAs1IWWb4ikJ
bljWiAaWAvW0l3l7rwkUSANaMqRMkQwRykiFk9hGGLAkX1kjAnfltlgpYUDSkChC
Ga/3bM/x0fWJoUqh7XU37QuwQUPW+dRbf4F6hq/8DNQmrIVMXjlv/i3KxBgK+E0+
g4mXuCKRf0z7gxmKNKvO6HX3NYy1wVjPrYNtT0xIBD4FXNsLtPXw3vdU2afXzxNN
COYWRYaW/1xlG/uoSYsTK01AjcQLH1D+lq7JSdu+FXEWd5HPMjpA3kUPkUTNBGq/
nloPpwxwzJ94aWyh0+HyivxtXccdJSUy6B3Yxpr5UfgFqpWftdqmZevxC0+yY+5l
EfIwziCLlVhbuQ5h3SAlA2WwlOLxxnHRizmv5p8jiOB/olPXldmjSWeyPFTntCCA
/0q5fRsbY32D+HJkh4ytaXYIYjXmufSz+nWFygnecLwBcdmnsL2gJCDFBQVdCnBE
512BRn7/s4zLXkuzo8+byzfEXoGcsq/p6p9vaTw1Zr7sjExMlHi3MqCLOdL0arFG
mrXwvLSQIC18bLl+FO4z5b76RO+e+JIrLHEqzGS+JczO5ijy+v9FIn4b7nDt8vkZ
zUl8u2AXao9xHyECg963VUDND7zP3my13jJ33bk4Dk9L5oMJPm7SVYGJOiHKii5s
jlaUbc5rm46PBo7OZ5Gq4BEhfThhYOxnxD2eUQDSL5NCTpxb15MYHn0bbZjyM2Fj
LhJuMovpXyLN79OCtmJqm1AAy+DZfqGDeBItBelmg8J52ySpMSL/QoBisjBf6Clx
azlFIdnqXiwBWalbS256F2f/tSVrbcOY940VMvRW3OhbJGnenzwGLo83PIJutTvz
CgS5U71tPohB4iKkSZilEJD5UAlhrXfBqyRapJ3CK+DoAP+QwiRzyP28Ahxfbasq
djRVGsVb642eBnQAsdL6Gk2o2MAAFpjtm2tJ0m6lbPIYPy3RMzkAPGoclQxmstfz
gKudmvA/W7FKl0j72X3kWDWYRMm5LTHL0porfh+f+IPo2Pumn0G4rdeFh+M49H/3
+JQE0dbZ0CNOG0TBuwzK1eto7187DjNoZTBrbSwgB8lQj+YpDTjLesjNy2UU6gr8
7QyzRS6xaYSJNwMm13frFWqMfncqDBADz8mGMAOs7X2LGuNinkgcp1Sieci5zXuN
uzH/MVuapOh1zYO/2qU1JYhvKkfqQhR90ua5sQiILP8pBsg0o2MHMkAnQACsI0MO
HqXlc2ktg5UpP20CY6AAN9pW+UKFCBF/m9zd9bzobDOLPkNkYI81kREloJgTgP+v
G76kt7g+nNfvG8/ANzGitiEQQHIGv7ZauSutvs/Xdo+D0rcx2saLdqZF9eUohPo/
SsjQ0Ud84WunT7DKm86CaKmyEwBqmVmSLs7iRNLeOS71XqKqAcfUHESOF+z6o0u7
5TkLTo7EkGj4l2f3LBwENVjjrgYnngSzJolpnPqiNKtXbb0yiHbIeIFby91A7PJb
uoGWs9UjbNk0/RJswk/VOz7a4B9QxLFddg4XoG+yhBHzbxjWw1XnE5+tETkNsCuU
kXLAXLrrqrSxZGu07/BK34B4+6lrvsrCct1FTS/tjY3MzYACzSjqJlmrAX96jlL3
FAm/x5CNXaAZ5e3R7Q25wOljAK1XObML6g/i1l6uJxfjOFs4rEAIUGrm6Lp9yhz2
IBRFxUG/lwkqO2nvi3bcJqV1MpTbFLBB1mepfirNCjyjHgOXdzKUKeY00qChirvS
PUPdzTPG0rL0dQaHg8Jw1dobMvHdJzKR+US0m8ojuFM8d0koYzqQ4tDJcOHDDnJg
LX+DT4iLcaDSL9rnN3+Mq51ot65vLHYXe0QW7DunTpC+SlxoroYYDn8RWVZiQZZ6
s+Mi+TBynzPKQvRguFHltiwVLMdcOdAsgqjr9PHnHT35Ond1EbZl3xXjjRZD1KBF
AzYz3LM/sC0bPvh6SbTDxioOUmCzXazcEHaYKgWNseZtRi2htbDf5rX8CDjom8AW
XbmXeH2tyTSbpysI/rMYwPOQwj1MOGDnwTLuHCMVG0lcpC92TFs6c5XKT98mcEG6
+ANXL5IokR74l75IGbHJgEHXPXnWFf7EHEAUAY7cMC5T/KEIgFRnzIuhh0MWCdyI
OtGtBqxnSiELx9BOoaPU72YG2Xc1BmUgh4s/UM9tlCgR5CPKvCyFbpRgFf0+cW+M
CKtcVMEYqdxmi5hFl//CU++LFlwRluHh06h5u0X1YDvfvCVZXuaxRM81Tpdyet+9
mROSY42EkgBVlfdyie0ooUcw7Go5+CLpAX3F2oN5ftNjYuUoL63dB7rIxxwFqd5S
L19kO7umRBHNsmBmjlRw22vC3efkaZIoFov9Flz3hQkUlHjhvEUt7KV/SNa4vUb3
5Z1H5uA+jxtPM3r2y81H4wq7Airhhhjw2v3kbLVsqQ7NOB51fHnOqXYWpx6D51AW
Ls0Bebf09cfowMkshiGUPQXfuWFF2lDXaptkWrKJYPyFUYORQUsis6RQGWxPP5/f
MPL8C9zy7kTVjjoQqwFnuAu/lokEwcPzOJXn/4hTatW/FMqTS/G99HxOgK00gClA
U9L0xUAjqxNwZG30xIkZZnIRxJjHeO+7IlNjhNxbSpOuGuv+1UshEw7fSgrHdw4m
OgnVMvluUN+xwwmL+Y4BISEYb9Tb1nayhuRQ+duo/QhXiViHzxlc5PRDZCfcbLKK
2teNNtXnEYdTVftgY/BF1fbfhAvYj2d2KbAsolAIR+EVqzALCJvnVtem2teDuYXp
oEaT+mgkbUeOyctpGCwwBNZMX10k07Eb+Nn/W7mbFzBamiIrK6F4Fu++lqHeKUpA
XvrYlMyDOhoSRkKJwouWW76lnK1/HZhklQb4McC+bKJK39tm0iDPcL8MrMdrNFR5
O+MKLUsGXbxZHUwO8sAbJqCnjARNNP0TwoTg3VWY0BBAK1v9n9pYmVJje4EWncEZ
jEbt29L+XFvMSVHQOrXF45Fa6XS1RhFfk7b6PAbuUXKpiiWop2P7YOAKRafbUToz
E715z5H7UyYsKirupE61Qczzk5I1Nq+OBUNKqIQyYqlgLEib3TU4wQAdvJn7mjWM
YOhyK80MqgduMvhFSEEotXJWl+Q4L6T9u7p21hgZpb9fgI78XrfVoIQH7Engbsb+
FasLQ04HMNuffcUg7RPVeWlqdTl79LxHo5baBXDtrB0i/vXfyBnHl1lnPu1KEy9N
Ij8rGEe4G46bK4CHRfL5HqQkloXxM2/lg88JvUomeYCLO8WhYFd8z9Fo52lWgGqP
VxS7gUFzRztrUk55wFnPH/DcKNC+H+03cKnIxj5mvsZlFNuZvCCrxRR45vnCkjm2
Dmp1gKLHQkeQIPb1PsYbO5IVcBZn0kxPACngyz/MFKYRkqN3nI4aPlhDuyiPGTiW
SqX5nQom48fmV+TSu0Xo88FlwSVrr8kZDmkeGRwqKG/ckemhVIKgMLKOUAGEW9Xx
Bn73xVbLnqKyzHliSyB6BeSU6sSFZGGE9AIr8rTMJBaT9BMkIEk+q1f3aWBu69tg
ZXBz3iYdx9ttSyzooBeJ41L+dz05wmMmwneCfKxjEIDLGR4BRLDf98P0NMvn+gW3
41ihLn4UhEDJf3JT4/Hk3sghSylsC/lb8jlIZWz5JO79Ad6QEQPthmNTMxynqqFS
YiyksBMBQTu5P9xhpH8I30/wfIDPWZ6tuY9FAg5R+rlLS93a3TMj4GCFOLT6DJUB
CbHo5OH/hisMT6ivYf0xYT/xoU+BYN21qN8iwZ33gO/wG9zJrSgif0f6UebkWOYl
s2148lqy6OpjBw8a9sPD8UxKsXHf4XZlkfGU7vxKNGLijVxUT5iskH6uexzXetan
SxCy+i9UmrwL4mDIdeUR7RqiiodOcppCt3t9MXY35G5I4eZBgVDtqJY8ZxNG5Md+
Jt411ugJEpuMTGwsa/odWDKya8HSlF181VKaku6pBu1gJ2hi1CdtmSTFcSdPIeIT
BFQ9ZiJt/kDfLnP5K/9ePaZ/BMlz4rn2Tbieg/S+JtpXtRAMA/L5CZKQQtayfk3R
Q97dItfc6NBT4GfsjYSm212792fDblt3Cjayil6vyvqzX6Qpe3Cz4g/WvKhhhh+E
LV0jS9xCqY7zdlTNPnOC58zhw94H8U0LtzGA3361tEf5u/WGGX+5kEvJ5QCUipXl
Vy4yW0kjUQ33gA78NyiN+AmSYNNB5fdk2b1WlgHj2n7KerPpjjmbK/pgrHCqjHOo
2y8a3FeRkm7TLMFZMFvajcYX6bxPgPakoFP+hPgBlnFgbSMnf4xtVrebci5I9tEi
Phke+Y1pHfhqQquqs1PtKA2mtEPytMGTty6O5glEqAUaq5zacj7XWyXrL+7dtDCh
5a1Un1nPe0v7k1DmkXFlD9pHxKuKviEhkT5IqvnLdQ2Ho7yzlBFESq/KCcia3bVW
kgit9THU8B6/wc8mj5A/dBvKTRCukzwgzYWTVMj1VkIsmTbE/EkXAckGt4q80aDp
VInFQk2Wpq7T6DvrbVrASX09qWmlD48EDiA3Gj29QTSIeOCMQmtnIhWC8DUt4NDf
DZb8U0FzHWlshPecotVAhpqyR11KEnE92O0kwePX3fwR2Gdlj4LO3VlYo9rKdWlw
dxclnc1SR1tPcH9AxYeczKgFvYOYphnJ0Hfsi1/rLDtSz0NU4aTtMu2a1CrfamsE
JHRjvzasQg1xhr/Bu9+dAOV+4HFwNyiCusbgho+HNSPPbTV4ZFcf+iFspJENQJJ1
w/mU+Mau0A+Aqy8XLA6TRStiR4KEAZTgyGk5J8zhCxHLBsLjnRXJxvSWb7UllebS
SNT5151VaqlRtlbfqDg5GMZM+oxHncyiZsE1LzzdoOD5qpVcpAkS+hEpEZ+yxj1f
vNWXKn40XI4jd1JoalB+3G1bJu38xADQcF3WM+myB4boaVHeBa4qMhBjS3M7QCzd
kxWuNrtU1fwqEHyvy4tJalE7/ogUxAa5/dq5WjH2i7H8Fyc0+HRaye3DZMXJcyG4
I9dnCz8vZm3qeqtCEd6fKud6qH5ina3sK9iZOcq4gCQp9cdtFVdmcioR3hJz8OBs
UIFXHn2p/Ly/PaDOXfwaVzy5n1k/YmkKmUiE2b/jekp5qanuv95TJxFAgcbC6Xo0
sNykdgYeT/M43DOMFFw3A7xnPgar/6WRkR/Qrq15Q7QGwBgpdCMuFSwMcpqmXLsr
jXmEFWXxyK8XWF5G6polcxHMof88RJzqB9YDPwUrtqGkGzHnxhgdk1WT6JutMS4U
q+f11fcM5Ct+NIwHqamhET8nPpEyCi9ieHEuSsD2uy8K30skbobm7VNCBt8p5xuk
nqyylXZ0j8l+K5WidnCRdoXlxXsTD5Sab4uCAp91m6AiyDtlXBKui7J3kPu7gk4Y
2DaKWItx/wqaWGFvlnio2BUw9yG/2qCQhykJfqDcGCAiE/53zntu+/EXqcBoOcRT
DAdG9kjhyIQmWqos5NvOBPMSm8KTBq3RgdfTdfn9dgLmZvwYXPt0nRxjRnyLdk/6
Df5sNIMTjnm/EGLRydNbyrFF54aM4BckwDrPv1SJXMaM9dMuYE2xCjgmqsIfL58T
b9SKKNChmN5chadrToyLQHe3QEu+7EcekDVcnDsWRA08CCMZi4dyQA2a6run5jTW
NiozI8L5pHQPcUwdOkW0q2vh3XKG0tBuASzIfViI6hwN/k7NgoPa5TtjeP8VXODU
DIQ9A0WACKc6fuc/jFs3fbAHVIkIxaDL0x9vWkrBe2EFJfsuxIxnLvblkMIS/t8r
njkmvNz2qDyZoNSN7Rg070yFrfr7435Z0sFBnRoClwC0yDPVH7JzSbcs9BRH9DvT
BDtKNIP36VwezjlgLvzx0LoxmCOylmb2atxqqa8xFh+vD68ko4/ca4hMJwMkhq1D
R6U3XR+iCrpv+kcesaj2mRJOILZl4fcOV/uAY4HovyyQ7il6vnNTQ2BPTGhQlb7p
n+aGk2jXXtM2Q5nsKFvtPPMla2qRUytORxM7PTc57dIqxSQlkU4uYM7g0VAYmWpF
XXk3Tlt8+vO/Dje1YJG/99I4GaCqqhU6w+yFC2dZnfxPg28j2Xxgqef8qsNv3jyb
lpcVzwA7bCt9mTsQoUoN3TbznzFB5GtMjDDlJMCEdq/FzJeyqMU8JO6YkMgp6wBp
ie94wU1sXBTzVXdXnIpjb3iYXiRJwaLRFmxW8gvQVq3Q11OMDewxBdCuhnvAvvcz
iVEnnd4x7R7kC6YmTinamw/D1EF8UPa4xUBCGqiQkLxB+GEShYcony35xVBIwOT1
zIasiNLQkBw6b8tpJktnf/Jrpg/B3DfPTJSKD55Q1NO8TS4t6ekcXGkvwOTq9NkI
zhnVPpY2PV+/hlSj7BtZKTjUCXvjUjVO5+2eEQSi6dIHlztIqfXB7i9gT5DptmRb
RePY4Vxj/PbeQPbruqI7JL7Xh2L9AnnDt9IwvwB3h7twjC8s4s0k7DNVHBJXbfSQ
7CK9l/53FFe/EJDpwWvfVZ43+MWgWIBVQK/X/GNukQOAMn+8/TepcwWsTdGtj5vI
/OOaXYM7GN0mzOImsMn/40jDdotxWxx4jgL2ODbQrRB9a1MxesuntwtuJK/4mY/2
2YLBegMd/miZfL+XHOhSO6YzsmhvMVVU4yj4YWRdAZWegO3T46xAZC8H19ZHID/U
RuRDUXo8NOhNB/3eXqLA1cJoEfMUZQSvkAyyTQNUnEcIO2uv7hNdEPY8ldKGfB+7
FfaERi2Rl2wpjrwbMhmslgaSi5AOShMQ5COs2e3Or38fTUv9TmyNYhsUkxO33hiz
QP4rmND7QhfmOmOcsP7Y9CLVjJZMq2jdjwSl/ksAqAN6j7Nwx4o2R3l25/lp0T00
hmdBneZReP/1MWlLHlM8L8VaRg7IR+eWWmmzIxUmAEbrA+nNZj95i3CSDwbx3gfa
qOKWCTtaEn6S43bTSvh+UEmAms1Scaj68IpPky/uYEIy/GYT94EN9SmT7hArYwe9
Urv1Wt//dXG2LTiYbpBBgeyo/qll/Qxfz3ZIHmfBR8Evu8EWtym/5puTXr/8VBji
zHc7AElm4vbwCeQaGiMOSzGT28oazLVvGYgsdtrAMD/3zAhp+eWmAAkXMlVqVQfU
kl2nnUjBn3dRc64skcCn8dzyVoefLCpfRut9WA6hxGZ8EeCFXiUms21+Z3TZHyjS
oIsy62e5s0fX+KzqXvg+sId8i0NBfRaKm5QAvbz4TZGdcREErKRzJgrDt6Kihx5w
OSJReeRr0BvEHUOx+B8w4Ne6Ezf2pSOC1LwbPuzfULUkOPqxFC3SZA5AfuIr5/k/
0udF6TjZXlxT/ubo0ClcGkrye1pkeBkgayq6qfqwowJVhEQ6PX/7GzCoPVeckkMA
nuVMD8FlonIr4LnvXfJT6ZOEQcNGUB7hsnB3IERq6KZWDszNJOIHBKc0adOCGRir
SZE2jUB9ezaEtlsNSA2e+Ex7JW90UrKcl3w/hXV0f5P4Zi3ju9lWIbfeTtsUt//f
v0WNek32c3W9ptOkHRS457j/KIzBbhIt+a5GNIabUvLaz2yaRgUrO0z8/y/zW8Bd
J74UFEHxlXYHfBv2n4wyyuMmcPcLpyKlxzfofSGK9io1mtSxZ6i65v7+JOS0yhGN
r/J4TM/uKs7m2hYkMlvWdQtqcszrX/frPtiAYj+wlzTjfmtzOkmUvwFb0+zdP8Ly
VW5U3zIroNSIGO9D4gIoKS6a2xvxsUkH3SHERZj63dI6ZPhrzED6XcDwVUUPgzXY
R/yo1GhmWhgIDJ2zzE789/jIpjusixjWHsMQUK/Jld/akhbSSV42v61TBUyzrdkB
6VC5rVa298B6RLPIgIiOPCH6GD0GbvFvO3BLX0SYXUGFtFVj84+lIqnaoKpqYNd/
8TUCagdYD2I3t1fz/ZxQENAjAuJVv4iJ40M6k+TM/qw2MTBrg+HuiNj7DTBCGEor
X/+0LAIyu+ygHyg2aEc7qr5cp1oLgZ8Qp2aC1/d9FVbv3bL6ZaSYtU9+StMa7Cm/
t4KrY8mLOGhQiKhxhFxUduvNAmT1jLj4BPhgWoj+rgOagYgminCAhOdzGAlqQzwT
dd3RIC30Mee+YV24vuaVDYl2l0EdObhV79w+Rt5CpwX9VOVtG67uqpm/jy96vrT0
P0MD810PCBbQ8Y/FJDsK4rGKB3yCo3Oek7Tv8r11R+mUqpT6x0/c/otBx9HRJBY1
Im6kn0ppexECAMQlaFwBXobIUlxyMagEMV8ee/G+uENsvT/0a014c/jAFDqpUze6
eLI35yGxYCF2/WAQ8S+LBdbYDjghnFpsuMwP8rSmTvJ61q8dLij59rdvPFUkzyTT
gdp0IWkhEfyTTTbAy90UjByip/uqMBrwdh3F7QPfpZVNT0ezYF+/nt9VixGOJvhI
KR5PBRMH7A2maRqn4dKvsdKZPa0G53IDlTEtfWVoj6oJ3Ye23XeWNUP95FpJRQxd
cOywz6XX5r6LU3Jr96kWgNjzqSWz0usB94SZbW5U+4BQcWMS7tLL+nw6UmCjdzpW
dtNviUfTXpLuqtWeYORcnRPltJjK7AlVZV1ZOwQWRPnQIYWWNLCJODxcD4vzscTZ
3P0JMPHGjFxo9ubPfX+0OykKuYzKn5RY5bnPVzFsEVubO19KmLxgLAS7NrWrFqmI
gi3+sn2xuvvhSDhux7N2dnHCTiZOtjgxZy8juov1U05bHu73274OPiEq6JEUEftn
ydRB2vG8DFo6hXCYhKpRCwPOfYsnj/bYlV6m2vk2fsUHcYV96c4IcQfcwWU1eIE7
iqCqmlDoVeq+NLYqjWV+JlH5lBhOvoh+M19uE+XwkY/ea5pWwwGL8tm9lf7S0iUS
D+n7Q1Qd3YLgphAkD8NwGaYbBsg10U6CVkc+nJS2wNnPrJkyGB94RsRZ5mO6Ew+E
mfODH4gF/zF4OVdd/Eguvz3cZCHRjhK5OG1qHrU0CBGfGBsNYD5cs5B/4nFcl3rY
BYnWdjisdTXpbMPXTjuOCgWxWs3ppmdQ0mAozVz9W5XR60ys8jeZPRlFW3NL5Qoa
ww/DJ+y6ht/5Sztfx454bi8M06+dj1bJ6D9wuxzZ5LwGFIUJrOgdBssoLa1kGFB/
Gd19N62SyMOaJfxwQemhFbmpNe+OWWdwAbfOU9dwRD+CRnamYle7KsIZoNh49tv4
XmYyDuGt5QsbEx5sTMaORA8Slu4wd7qeRcArl5hpA9M6LnWwKJcUhiNdUCBlHeqX
8Sbq181TvWWJ+WalzFWBW0/I6fI0gFEEkkT5FT2b8MISwtNsovvhZ+kyzqjqOyhB
y07idNHsvwKOTzTRA843YGX3BeP4gQDIx7aewrOBkIaYvOXhk6wgpGJHSKfvd/Hf
5WOurVs+PthZNqlDnTT6PO3s+TLKUD3CRNk947zCDNpat2OtOrpwYiTAtnDPt9Ka
Eh+XpXARNejQ+qXLND+KpqXBwRonc1DlW8zacShvQkwGDcTDr90cOl9qx0lmPk/W
mPs3SJe2LOcKXeH7ZSkPHtMcFlOu3w9yz/k/+MrXMACXrY5243l+CajgDDTjr70O
qK+ml80mzKTuNz6h+SRCXjo6kdtKa+vlGVTn93y93ot0fj12TT+5RgbnJMMWNRzz
9ivWnhPAlw8QbJvGlBRNTzHxwA1wlRZdlumUx/nx7teIUX+yYjbDTH0M2o5SH0Nd
4N2IrAjt7Fr6AR/XhRvlz5GH2ZQYzVjbntqr9CTnLg61qsE++ufsBV+zQ4mPiv3D
kdWBraR67MtuG9Bl0hcFsS7S7qC4uvaYl0BKbee121Xh0li7ZptKf/vjrh2KyJ6q
u3spoqHOMPyTgNzh90+Ss7R+ko5icLXVJEpBiWKLQ7GZ8wuSjnnbHv8hufl8M13h
HFvOXC/7he3Bk+wcQVtUtgD/cHxheuYsKcDkSbvJUNEq6PdzXtMOcvYiBB1/IkwT
0u9iE1Y1YMLzZOis5DOLQZMbPC4Z3yqgyb/YVi79MbM8yYh4XK0/TU06oPyJurkK
AnNraS+J7DlUoGe8fPY7u9hHkldolRQxJLaeve14KWL8GpvI7BeTzEkpM6tU5UWr
qNYmqLiiQMiPCOWYTYAcGhHcl4c/cg5x7cUo9devzUXI3jB37V7VMA0MwXZyk1Uw
l27EWRWRFnWzsOVnmB2HbRwRgtC9af/il9+eRQghakBHLcvxd4Ns05Qi6NLeebbG
h3cI/cc0UOKS1xCS/k/mrjY9xwTPAixqO6BHUjDqrb5l/SVoSS331ePZR8lalkrB
WbdQPGaLUWR4XTnm7kKsmpJ/fDXQX1xGwNij8TaQvnrWzUovOJT8nHCcxGZrkdng
+JU1yWSsli8lvenEcxZUqvQqYWdFQ3QSxlil2DeZKBUhByNABVYMcUJ0rKMUas6S
Vixp/NqYnDiavVurZuzIC0ulYhPqhndaj/m8fG3LVyP2unNriIJeCRUjAPlyFjjs
qkTbbg0bvFwVx9GbVLq6DeeYFDiXkeEUN11YS2ksngi/Feh67XfbDQADszs6SKDI
4SxP/vS8lfft0tim1eeiknaHA7RL5ouZNaz99Qm9TM/0WJFhlGcklWUJfLm9jwSE
SRSMUd1LHZTImCmw1TO00SVmlNmrQZrhs0NZnYpMMBHbjD+lKrM/EfEpM5pFQ4Qu
sITkhgYiED/n3ek6WeezHTxLjqlnNVPtSq26swllAsUtNtZFmfY1a4k6npQtpuvX
a0+EIiCJQRPVrH+QTAwvj6YhCmS4qDqk/fTO8hc6axx0faFTMCtbv8YaI3nucuYx
TWnDSKkhGAjmC1JDceBQAh3M0PEdImqi2VajSt9a8khsfLgLftzMJDpRkCZZ4LxM
heuybYsl5Loo6BQ/zd3FhxC23LdnE2bmoVxuP+BM+lQZmypoSvzozM9SdbEZWYFZ
hVEQ425eaC8luy9lTgzZRYtc+dKVp+dQagspwANvntgZAtBDDA3Ej+X5/izCT2pv
6HoMSVomu+aX7nIr6XCK6kQjiR/cPDcz+TpSqaRo3MotzoTgLsed2yu/lB6a+1ZH
hpPoGBDVPga0VznlFd91ofFqZk1+FZ73XstT/WNp3laaVFegpptDzyqKNIeTow0h
UmFCjLtZ1GNuglESXdX2MCn6ePWGreH8A8jfECGXJrDeqvhO+97ZUcn1KIRgy1EX
ESrclGV9/EoDyigLsqWp+W42kWrUGqzI1rIvLHL3eLNbLKZ4Xe/lJNuX4kuYIIHF
mUV+ajMvQ1U4nrLNaVlrx2PlbXUO/jEcM5IyuYvd1rdYzqu88pBC/MDGzCCM6Tca
H5zajPfxk5qS1dqx/WeE1sEux/lk9u6zj82uAnI/M0ST1LvjOhTIYC0hjyFXILob
J4IgV8TxSCNIKKWsuNR3nsT+8lsbN+lPNX6nAqFYcEzqFg31H3SwGXPBj79Qw8Bz
eG/QgGfJ/egAqWMeGvHdcJN0u4PZxPvXhKnxHvhZ00ufMg+iHq6QKktsUAPYhp66
p1z+VyYGbk3SjbuaacrLQYViKdn0DHJcXLH7i0IOVCU6ubgXtUewgO4hlLFOtpLm
r6hv0Bl4EvuK8h0/7yKZtKo8Irf1swg108aPdm5fdNje1tBAA4LJllA6poUQ2NCR
BoFLJygrlEuo6R7KVZ2KoXnHyldKVZthwxMvLwCwm7IAXhqzj9Y//J2JPhtvUsPl
vSuUZFNux69d+4wcEpBow/A13wT5jq8/t5Qq7OrVTNJMoLE491El7N9Ji4rjI14f
FjixV7ocblXlJnVWjLbb7fjD6wOivKLnEKU8u9XcLRx4ZWFaK6sIHBNsLj7HkokD
Fcziiheyw2fYopzLpvLYPI8JnsrIMs2LvGoElZWBMYaBi8FgIFTMjhl+SBmkytir
Eg5qKDk0VnvNaBmtkpzvi2vc5do+ifrzMzDEahcRa3ufMe5IAAaSwgVaFXVJXuR2
SB4wTzM03Pef1NANZe1KChseffU6obbTDEJ1gUnxvp1Ju5jZE6HReeiCIFBVLlLx
jNzpomcLPIA850lNXWfBteczpF0Y5eUlF+SzVWRklEljOuUhUX0jvQH/t15a71MW
I+1nss8vEaCPn3SYd/AwxGsiTAREMXWPei4zoIzphog82wEK8UshQe80ZY4WkDTu
zJq3acyzz9L+3IwJeWOIZG1q5tfAcW3e7VsIT+/UGSg3UyMfpdvZEmi48V6oKRMO
4PoqdsP4ZohEWIdsSac5Xz9HzkI0240Mo9Et6tjPjLHZOGPnarH4rCRlbINHAp21
3EpGFLj392+zxb2suYSzqaDBcKMaSBjDyY274iXo1qNqqd4/ZoCwZOydnF37xApu
OK3pQ1mFH8u7aMUPbXRuNywhja8Fq3rbLj/9oYxiWqghnLgpOsLJIimfAkyQCK+L
hRvAqrua2DnTTYWDYUoES9hgRv+wAgGAUR+PdTcEFR8qVI4hOWnF++n7z84GvvGT
CqR9enrJrSGG5+E8qedunW/1keyDmxK1suC8yESZcPaS/lwhlfrp93AhId1iQbBn
0zlOZOxvDFWTKUJTBdOQcJOBJ4xchoJgz/JtcnTu0wiSDWBgOsC7S4THouFvceGg
U9ViOPa0SW4+Jt1d4oy2MQr+BTMirB926/3X8F5XYzu5N5MBI65rp5+iR+8oukof
hMw82IEJaoFtzNyyRsSyq/3dCv4L3e/LwYcfY5t+uT6EhtLpZQiukAHHmFxb/u8O
Q2w1QQx3QLQbtk3sye0UxDZDRQvvfNALdkQwjo2OCiuEzUCXtO5g+85T+gMSo17l
Ub+2R27H4TTw3NjWGqnLB5zaEOmx3JRp0JqHY4Yl4Z+H4htk6Aa0oGAqFis5R+qO
PHS/CgaWu+EXLxOO4XicrP4IKlHzQvMxp74GYFwyuk7pM3D2YfMVv1x9ept8TE6g
G5BUwLZ2BoxLC6eAf+BN43HY2PcG1s4WQmU0FlaDqvqkru7hJVPNu8hZPzRWG06V
++NsqYT/Qt/kEwG0ZU/zYO8aEgIyUtvnlhPxvkuPcn7t9SK15hySAvshL/wLYGmo
1uvF5PPam18AK4hcf+Sakj4QW+rIl57Y+6mq/7y2RIpbFbkMCmkiVGC0MzCaKJ2+
L9Uf/sz0/rNWvhy5xETHVhclPIKTtcw7AUQfV77R5T/7TR770AWrXGs1MANVY6vx
MGfp1hj9/ZALLeuiB4BwSuMRCwIkE/gHTrtmZippv3YLB8ZvEK2N3T+8sY6fXvK7
HsnpDRrdevv0NNap0FtuVJvhJj6p4GMBVIQf6Aq8ZGbHZJul6A9NDBdxmvh4/eoH
5x8o4v2rceinXDutVVAWWiPSBjTpyoivF3ejZG8wKTfqM8h0HE2kkaihdo4srmab
hfzVr5O/8p5U2vJjFAxkDu971CsHHBcjH07uIl0Z/HRFDOtXiJxwlnJs6mXpO9h8
fIfF4FrHFE/YRu2UcWXPcgA2o74EPBNb+9Si7MUDVaDZl+eEADW2HkdZGoDAw8w4
/LKFT8tbxNdsBOwgerQurS09N/686a2jC1Go+GTR22FFS2EUpKA2hidPrxoa45Ph
0b+rbeo77A8QJh7oqaHVSP6/TO29eC6pzFBAt0U4HOMcvJxbxfIs8d4boqSQ6BcS
Mqahk+CUzO2G9aNy8zXZm5GpoWGa7Wx2i1mmUcnIIZOIiUFMvjPiIHU5cNC0MOnm
4crWmGrrt4C8Dk9+klePvnJVv7bkHKL9MqhNQoZXLvvboF/Jknb2Lh4u2U4h0btp
6Sf1+k6IKKkYtJ9r55CN4NE7WM40mmg13sAANsWPPxBWy+EHlwTXYJcK93Efx0AW
8fPfcJb/YtFqiNuig+e7RlEEKoX8JB9dn64SwKiEtEg8o7errYVmA3j0bxaQJgIS
mHPiGYXV4fENgz6LLpduZGSyqq5hoq/og//8uGuMJf1c6WYrUElxEp5KJnoromOm
5TVUY+GOFmx+6E29suDHjecZ8GJRqfLuMvVietO5mX+P6wD9MpsDgaUPN3srTJMD
CcqZVd0X8EJ+glhFb/SDfgUwUolH/Tw/+ZZWMvC1URR4l9xH0pnmcy7Q1Mwvmd7r
kR5upIo6MW7gPG/6mi3mXL+3G9GKSmVg2rkKzDnxHNBwei8fiTv9BYUkeNgRni1m
zAlKLFBugAgpJFDlLSMfZgD3BgaT0LVlS6dt6ufkDuxHhAj5VrgMJWTjVjlO5j6V
XaKMNB/Sz70RNVPXo63bUQbZZzI1sa9ldsI8a9EqwzXXbLLaTGXMTuKSaLXowY/C
7ZmLlXha8zh4kQ4iLlh0JmkFFUZXTPqSHEeDxPdDqRDS5PTHBik5Dz0OA+EfUd1l
NvIJ/Of/LLolnSDqCulrrJh0lYaYKWdc0hXaI4ACL/sEj14XBpKUB3Ov8ZOLE0bi
zmYc+xN7LqeGzWFUcf3Wev3PCloQzgtl5l/qjdA9tDTKrOogMDbd8FOqkTrs4mz9
ntIxWllcilzp1WjRUZYdjngczCj1TzF7Q/1O3ERWb1e0W2DnRBLWTeydGCNnW+Q8
OzewraEqpOfIBkHGWSA7xAV8WB+ACR9Ftls26mHTvtDzVyBBFayeO2ABlJsNZCCB
fAnzsCx11m0ykzzd86W6UwTlc+JrWl9J1RfhlKUPW+at5NSHjy/qRsP2rC/tfexQ
1hvyNhCYd2I00qJ1Q2XIvi+J9OBUwT7KyGVhOft2g5HrdKGxuAVJfBm3HMiM8fbA
3Xpx/3G6NXL7N8XcLiMHHuOwBA84DxpSDiUThYXWqxLlezuI59KugBzAmC6ENkkc
9kaFLUCgzkC1dCCpLp49SBPrRRMDj+G/fftpdneGKLXPRhc8KuwnGIgaUvSYG+ci
5T5XcIpkkZrRIecWQeR7qenjJL06C26BsIJbOiUUXLWFuqEIq5j+b+qkBLFSSBli
ThL2wP2XElqC7kwpFC5LWFZevjNavnYFWAORCHoIPzdQgT87Or/iklEGglCyNffG
U0yfZo+k+W+yDWD9UMskJLVFdhrUOH1f7OV/9G8KwxiwnBpGEydJtNFds+DGYM3N
kHl8a4nWvhJfgvbXfPNweL6eWCpEYFLLamrmNwR+pnM3jvlQMxwOlfMjq2qkKBXD
gCFGXJAVxVuXSMFA5SIJe8ZBsBeNu8+pUO1FtyCBKJoqMusucYNRdIV/ZcgTwQF+
xU9bIBu41uEKCShFfSr/uPfdwJ54Q+T8LIDld5mj1H8gOWb9D6QFdrBsFH6wDL5g
srYi4obp3wvSPvTc8PY8K4LY1JMalCcc1tJQ56gD8EzPa1/Rl7IYmM9d32EmlkJU
emXNktj7JLdIQEely/Wn8yxheOFnspkBAdwoPEU7FgPHVpSFO/Q++QkRNCDV26QU
lbWBMTWG+g53rSlvQozg3pKY4E/6ZKgeuuveFeNtOKOd6vv1m89JURiKFlcnQgeG
ziX5DC2pSiQb9/5XWQKaZr+K4zR9peHZ0jPulmi0pp8iDgw8cnL4yYwFCydK/snB
dJzXUc/ZSIMpLiszFqgkCTex3Jn6WFdhTi6GnIacCjZyMd93sZZahoRwz+eM2ZqF
EO+x8ouJ34yRS6oZbekLasb3WE21ED3faXES30nTbqajNCZs5bXpKu1GJRp2jkvt
RVjlG9BmPf+9AAeXPHoS9LG7mcvOedokvMQqilDczI9wWr5JOCjLRgSsyqxpJmNJ
kMn5H4qpGNRLQWJrMHdsH3pdt/arm7UHYNL7hBBOOsdW6VC8KjD8C0SaJqc/cnWK
75mqC2Wa4bBcQr/UHy7TBT88nvSH1KOnpjzzNW76Q04N9BSG3Z4fuSLnWlgDXYSO
K315P+WB2Cq7GQ42mnTg08M5i71gmkOAAR7nNpmEizpY4mdr2mnndQRINPqSbkPS
JTfl/hGB2kgWbr3UU+fkLNJ3VdRtnIIIkSvn9B2Nh7xSfP7vT9UMIkCjAIpu+RlZ
OWXukfq61Ogvame+jBX5Y4hWy07YEpcZkuV+sIcmz02w1eubjU3tpqfv2ejP3bZS
lNTGPiaoiG/6IxUAOIW6/lV+GRjYb4wVX7AWUZ6uUhE8PSZofVZ9coicZgfrYh9L
aBl2CxyCxF+ptav8LLiyrBASkZyS7IArSfDTdNBhlNqxH7jRK8JhvpjuoXbAQsIu
D1wsqYc9yHmPN5CdiLkwXgUbzzSx7BbXFqV7fDIIutmq7lwVpqrghxXuSN+TFrwQ
0s3Pasp+oTP08aDHeD1Bqp8fN996qU7m6/B8NG5oueSJl+fMYHeqE+PNES/UecV3
x/j+KAUt1KegQRbAMbPfFQzPsxBtr+rU+Acz9G2yRMcp4tMRrkZb1SEpqZ6CYJBr
DyZP7W3p567qmoXsstLwR4npZ61WzhwSgCW4agBdMcvWmc63hNuOrBkyW+ze/NZ8
0RkZQNv6JI4hPRrHwBpCv6ivYKH+bajiaLfyT6s8lbFBvYz4Aws9VKrEoljuFt3M
TSW+2sOTL9a9AtRnsVeJqhtdv66gl9+s0cWYFTfEIyvNvqGZRgQC56d42t1pAJqJ
KIdziR/3Gj1RtsD3JWVu2V/nOXJTy+6t0P781xqB/67U5/Eqcq5H3i5f/oFSjEag
Wt+DjYLOsekijW6hMX50MYGWSoaTIvWf1QKdVZ05n79gmYO01xInczur4keVKNFr
141C5rujj5aLEp/J2IzwoypRA7NMAM9/F9+c6mtDgXuFVxHXd/kExcQIOkApNn59
iWzeKWbVMPqdC56MeAPMyE1NX0fd2IthqDo8/c1+xZR1vYCvxGxUhCcAlQyq7K3D
cSwiGCKFhpTmc5HOZqj6SIK0It0viDHpNCPJg/iU/EGhONY7OaJ/FOxBajUz7qVD
YToYJLleucT0mEkFlhlwDRKO3MxlW6rMq5YRKMNjWS4OqL9wE+rktaPsG2tj5YiE
Z+2CfVzUHE2a37tpub1PMtziZfFF6Zv5yhCMiTzHa6gmBLEONH1jJQzby6qhIRQB
9wa+hcD1Wm8reZMvE4Dbtq99nMk2JxDwsDx+zJbdmvu7CoRHXf/GSaJQ3U6ekPxW
ZYEbQ4+zQpGzvavUMAhlyfmqDn6UbWsg/NUWi57XEfRxxNKinZndSrW5Bi9oNMqz
rp+mVqK5x6S0Odk4Xh5z6h4EkRfyCavCQyII3SQi4neJfUaxOYp2LwC1jQZDzUS6
MkfCXXT/HfnU4gkF44+ESMnVR+W3q7ega33C9zIY5C3/3AL1+sh0ROUfkWSz3nYU
3JVPoL57sAJ+pBiHNHqqFDf4IPLHoYr8ILT5iX7nbGJa78sREbHFEt0KxXBoZj5R
bfEO7zeGfxFmH2aBeO0upJOyR1yG8jf40k86D5zIM3+VMZNtoA5WSn5i7HswPcGo
G1luUc7rofIDflboha4Flyh0eW5SeW8kKmawPZVbpodU8uKi2QnCcPEt0S1lNm7S
SdZ9UJ5zQmNGInQIRMYIkYUJs5yX4BinWc+1wKVM/OPonwV6aZ0WVQH7tfU44yLF
D+eA2q6icGtT0ON6cjn5018AilHLZpvWVpkXKZaWYzVUxYMCpkz8QtTjAqxDZNea
ZYFZMpztRYDLqtVh2BFSJyc5YXKOa9dIuC/OW4CRfYknxt+5nsoqb6PeiSroD7Je
gDWxJtopLrCormSBomaF/dEog4EGiM2Df5nRl7po/gBzwRYRxhd6zeKlzHIfaNI+
Ati3bDkxS73JTcA61kn6KU9GyxsmYyiCuj7aUB/YwU0lHRJrQX8f8bN6PXSKyuP1
JpMf2eY9bEvzVCvZh57NkwMvIitNym7oANr/PGW1a9awfJ9nhd4gHAYYdigDF8pA
JaRdY5/BgGP8/iRQ1upwRM/iFdUyjBbgJkzj5udpY4G7Pgrar+BrJRN3GsCHwC6Y
e+PAdsiFHosjJ5B72LmJcTOgOKY2k6G8umd+fiRFrj7CBshPSO9tAAaz8yEEKfkp
n2Ylvd+DqMQaHT+UxIGP4Zjzye6zlsSrAcXSH8eV2iGl7/jhd0PDn40ZxDbF2UAY
6wi04MJGfVJfDghghieUZiKcV9IL28tcyVfDExNM5cKl29WtovlcNgmGy5DPbogS
FWIBaUdUqSDHTg2lx3t+tcrxaUEKrbCysINmRfPwGLDgcHSJLpbXuCuIUgxszPhO
BN4JiZVL5JHsTxVknOG1zSbdBIzMf1aCtvLUuK0xPy71a+WLEsH6sJn9BeAlcxVJ
4CBsJqOAXlN/dCDEJ8rHr9EBNNMr1W1+a7AAuI9sRtZlVoeWYoDmThfBuv2X110O
gCu8Ay6MyJc0VXIj3oo+yGtnjAZl10WuTphxEW7CUBGQ8SqA3CDVrjL956uxle2B
GHO+67ASUQMCdrgDuBcMnqoKXV0MjaCZvdrgUEdCCfGx/HZQeiZrJ4lc1UJemHKR
Mh1Z/bnCxCNCHvRywXAUMEgFswQZP8XU9BqV2QV0QvHF+iRn9nzEF0tner3pTSqo
KCktSEWM5bmv8c0OI0lWRQK2iJujbmAxAZW/zoGl3XuXYNZYKDvUFcChPAagyclY
fNCoBF0KnX+w7qpbh36n3qDF2Xgj3/88kC/V8VFF7Lblo/EG+gXh5CDo9bV3N33j
HWH9iEez/26C2Us7rlkf0KwECLGCNa/6easI0h9SDu4C8FqKACEakdfhUdcRCr4w
nBGrkzcuuPq8xYc+ru/oB2+q9vJLNe2HyGilufJjDwTsOHYIRIXZo46ECSRBpHRW
JKTIbvdA2jgWc5n6tTsNsZkVYB9Y8o9h28z0X7/SjDdXziqOBhv6auRuXHP++xpH
DYNiYY/tR6ZOnbLgCwz7CzpjXXS7X0vppuNqyCqQUeuAJAKWgn5ZVkGt5z3cudwo
Uo6en5y3FMEZLvhtiXdA6Xbln7SOQbbLNIqq8ut6dTLbDc4VZp+JvXKaKh0AiFc4
sDQ+W+mZnUYuFPP4kwGDbkvdLSuvQwj4kDp4Niai+KZFxCMy+9dFzMDhkAuSqdDc
rF2UO/0jq/gF9OgwJaSzE+Re3JqkzNcZIfK+0iBDBXSKYQnYuby5zpV0PKahVxRm
6kg7CmbTfI67F4ad+567K1tfdzrTaAOCu6wsClM/SGbpZq+vUS6l5Sht7at7d+lY
6S5lX2B8ueiqDAr0SbSDLpm47BACLmJPqLVmvrLvWW/9MzU7/gg3iHOA+OjQMNkz
GKfEp3eLlTOjX/OGbx7sP91fKzNzaZkITWYODrbDuK65CtvArxo7BXNIFxgKJ6lr
UMxRmTjHlapUx3meounDiStgYK5+NoPm7jMOmBOKwU6qY7mNzV8V+ceGtslUPx+N
YBo56DkvTDvJjL8BmFcXJoQ652BiTczafd68212eeG7D+w3nS84JT0att6u34RJT
xlj/26W4gzt5GL/W1SmjGKYV4/QURBcsbTThSGCqDi/tKlDOJ/F1OSW4/u6+2ABD
x8vCe1RD3WMr/gpoNtokTHMeRos5mooU3woXXDWXvMYc+4Kp6xHz9Iyb9c2dvNgz
STIZuJuRL5JZ/xUwXFsmxb7lqpmU68xwtO3UeMgv1i2YCHYiiNxZK5q31WthoFKW
07Wr0uJw1vWj07dUvw3uWptQhvPKr0sVLXlxXKxvXy8Gs3cxU05ymNxNBmzY9iug
ojzzsjsiZVZGcbIXjLv6Em3gkcibjKHoIfC9RWxochpuln567JBOjMfxWoOY/PuR
Y0GuvTNWgb79B7vp6Fn4IJG3FxIZhD7Zb/Uo6s1ctnTzUcffNbT/cN30LBLkxk6M
yNplkMNL6dXhbSp4gqTv+KGTRPoAUbdK0dWoEDThSnQJiPiS+5RaMp4DdUX2Rpvr
2xwm15yJnviIfzcKSQ5cd5sOETGbAXB1B3rOV5pWIz28pM3TbCKJ7aWt9Hyg5OUO
U/eRFEmQoEBJT+NiJf3e15K0XBqXDiLO53LT5KddVQrkcb+ic8Ka1pSK79ky2c0S
Ed4dKz+/TGSY7FyMRLJ54ksB/zuVTo1e4iO4d0uoxYdZSNFhXUVKSVqw4Dn3UHY6
fX/6dCuUdMLOZydpLxuJKeIVuZzlkAk1Iwi34IzW8D2LuBXfTK14CGuvFpdVxry/
/kmXnlU6c68GmlJAJVI9+Pix0ohK+0kN/k6VqhbLJj366rbejs2R9hTMVwarXI6H
RJESCOuxgtK0FAwDKqpsxvsCY8g9NxT4moiBj7Hzz2ZYrrK/8yg6eFSfGEHMUrqD
3hxU4trljBNtet/8CQqsSHjQC7SOjkapRi67BUx5KCME3lBChBvOOBTGVrp0Zj/h
4YvlU+3vwwhEwJvWAfC09jxcKMxRcOHRnr1sUN63KCeniXnlgetK7Tq4WwVI7aZc
W4VrNQWvEcI6B1IcwPfqfc6ncaZwrwbspFGz0sXt1KZmF06ClLfMJeUM9LODWuLO
C1r+5hczzbHyKTMHIa/fgQo9zfwUQoZCY4h/tG0CR0lAul/K+85uyLvZWPgRWE/P
2gweIhwU8w0INT8vVquGj4SkO4vlZIOwmxpxVg0p8jTva90DknCLztTiWQQvOcW5
+lANgsu9Qy+hTE3hfvcqKzkJZ/V4m0TNYofGqipdM3nwXdXURp39xj3h9b4rj8u/
SBYNJmo+9W9kIa8ENIaoFovJdXynoOThLgrYfgzg4bFyK3VoY7kUYOcdttfzLwJK
wblZw6z4TuqzaaaxfTGvcKGr0n3VvhW/bCDlq/51cVzLS0lt8XYPnmMs3coyU/Jc
n2aVL8XSV/pYhRyRf949RQIWLpSULID+tPwyiHD1pGzGTnlWxy3NNBW296n6Pei0
h/suiicVK4XmJKq0fhpA4jQOznosTsPgFbGVHigckJT7wJPl9MFESsuC2VaeFi0j
vFU6vgkLNeNwoZEkl54bFRuGMEPeKyEL6lWEstLlXSXzr8eyPWcrjxEKiZaLFO5w
BuDOZ6mpfXPYWCMF5nspgkpL9yuM1OvZ0iRe3Gz/mxTceZXuOG1saERzOTLnp10d
uSuNOLcVv/0xjYmyt5g54PSi4F5f2SCmrtEFnZD3WOhnRQcGOSvOPgX9fNUi+PCQ
AqBK9rbSFqiXflZ4D6FlOOMJifg9mQ5S7qqQGpx5EmiEaN6hkp6SgYOhcJIoPJcA
XPwQX9ONVuAJJMs7tAEhNd5nKLyBR4NIQfcGQqK//ffcYQ2OLmW/rPFLw5nhGBLo
X1TDBKi9OrTWyoWqsEbHU5pVMTfyzluh3ToWIDovvJuwXVgE9fd0PX5gmJtco3Tj
RC82YaSkPKvXnnRf6KB2CVMPdNEfwmqj268QP0v/pDwYPU6ceMnHOhDO76ORiJ1B
lNcQKp56yfOQr2kEt71mS9s+FkP6QXCTl6i2d7WKqZ2wSX1clySPhHk6UpInmmmZ
zQRYv1TvkTmCLDTGx4JOmAIgtISsTFjkZo6JTFfq0xRoUXfuv8WQWIcw6KGv+Z4m
KHsBU0s4k7/YnasWZ3F0R996MgaOwBCGBZi5Y+196wsPZSifUWajR9KHigeI5cT/
my5rdyGMSA0ze92cTr4Dc3+wfMfaXSA6NNLcWFfru9bvth+DOzZ0fogArmgGm3Zq
/qFBzEQdgFelQ/47NfjMPrZdOjewwRAgjZ5zdZ7Ikv7xnKOQe46vEaBVbJksMRdR
b9h/txFg5vh5/wmi8hFGSw8hGHqWpxL6bQlwKjo4goPAqJrhCGdp951SYL6mIcsZ
lX9e7Ox3KpYkOAZa+ySk+445THEUbjSI4v8PNaCuXWnMKTHYVWvhKOoa/6DJ/jHw
1NKgyrcpRWPHWakl48ir8QBfI5aQWqqmHo3+ZOMqvKrSIpqOdhJFi40rt/ZoimdM
n1KNO2dU8OrfKWCdm5esdOEEKl/ZmPlx/JmVNm0fMzckZxU4fqg9bSgL5r/9TB/Y
78SnlwZmBKJ8aTiJJ7ir/oXy7ZNk58D8VdJIARlgIpVjwKhrY44FScE9bhbY0Ggw
tvqd4s4e5UVcxlbD3QayejbdHZZVjo8KrB4m66eWaZZAf31SBjSx+9PcPXxhswY6
eoAHaWD3Ahl/cuCXom0Hecr1zVjxs6PflFA8nMxYcLMLlntH+GsZr2STXNsGpzEW
MxbU8kSvCj3kZPyxik9A+rae3Msrlv0DhuVIihzGTTxxwrT9No0Pg2HJyEehpxsL
QhqPJLZepeosZwWZRriSIxTRUWv6TmZ3OJ+R9r5MsabqrTtm2CSOtegnzRGz4lIT
3Z/kZD/fm4lpE6EQWqTaoGJ9qqBcBVsqofOfhQxdzlT0AJMrlt+RyAnrcIoTj5j4
yHVSbxN4dmwFZn7OSOaD7FmW/adwqiYyb+07JjnGE3L4cBKg88b3OnvhhcfnHTNn
Y9HAckXqdSFBAU+IF/UfVYfBbAV0p1D7dkdMUzMQwr1B1VFvMzDlqkbh/NLvbuWi
0b+jL4Q92W6H7SCjmGacnoMZfEiKgT7IAR/R+cr3eFgrMDdkmy1QV1uXeHfpGxN2
B+N8OPifU7zfyUsoBSiBfvgK7hvSJF5/028bW2fCUf/bJpIf0rdeUubVccNvGdat
HFTJYLaLWqFZG2O4prPlo4XgKGM1Gb2UJUsBUhDUUi6EpjY/w60LBTCfug+hTtmn
KiIKSQWN7VtPhZvX6BoJm0VUyIzSpzaG40pJ0mHcsD/CJnRcqIQ45z+8X9rU/ac8
f5QJ5bOBgWs9lm4ozhLaC4SUzCiRCRukOZR3+ZImhaUv5cdjOD5Mc2LDZdIa1/Ac
VM89SvpOyZR0YnPNAtDIoPcax4INxEI5wYIxAPm+xsI21XbiCXFJfoYb0uk7Uv/J
mHJdIRec1RwIXJcbBO9XRTGGMK1qreX0IeMfEM97mbiPgqDYt+CQSk+rEfna/4Jh
ywE2CR/Ulj9LB96bkMWz1ts52PAtMQzJC90/M8IhfNw+OJ2Wl1V68XUK9+CmpqDS
JnNT3ogr1/zugfDtDoZFwggJ5Yt/MV7a+vWO/BEk/7xbIZ2tMRkTfKDDktcxepaQ
EGOitlwGLRsWTq6+I7jSkkBlDnACZTwQYbHdFX8bsP545fLPez5aP15p4kKxGqEQ
5Dl4ht4HR7BvxOYA35Acv6t8pqdEIhQVVIYB6s4YHtQRs2ikRiqArDw+gqRYEy/c
TVqlknBDqIBDYl2fyOUSXPglxEqpXu/C1HzHGLN68ahw8EP94MehaVAiA5gBsxgJ
80vEQiNqkVKihQeyl4DRljc+jcIlwAfipbK2DwymAeABVUtube8/+mZmo9rOPF2B
L+RdgDUtdFV9K9YmX74Yi2z+ZwDMkDL+z+k1Tj1ul+mB8/d0YFaPEt99s6QNpUpa
Cv+eOr5Sb5UmYhsp9f7VhIUNpxV0cQhJsUcb/z6UfsgmoU95drCqenHh4I9NVj03
F6hzgzN3ILPjBdtyqi1xytzW6ItYe7MX+JsT+I9SoYRxYxNy0rx7nxeXUPA+8gOo
tWW1baB2I26WuCAhKbzYbQ5Req4iaenuKE/oEkXwvWLKa9eQ470XcHjVJvCJrPdt
EHNUvstMPxI3WhzrZNR6xsHKTbk5UUZFmS4RPCHCo0URzPz/AF6mRCG1OqlmFWLn
z5utSL/1cBDZvvlxOxY/Gr0qNSuMJ4JO2F/Ecue99Xvy4Rgrpf0iyXBsWoWdtZAn
2R3O22NtBP2ofgUAPU+91jFHsy0LcNDRXZKJI3tg6b+IaiA7GqkLsdR7tJDtAPCg
WmDcWORTyyOaCcF/JSET+8pTzoDEzJKOmE1nf1vjd1VlFu5YytdOlHMTtG9qvSCG
pkWCd+2up5+feURj/bV6V24mOZ0rawu0DCp0BjDgGdd/DWeVmHr03c4rlO4slxq5
a95M1V1aHAqzdRKsT2S8gzll8mOCa+N+ZaOTuIhud9tbuPqKjFzeOrXSras1xYJW
2a1CWfIZAQhA01e5j5B+wU1RVHMCWrTWdeyUS8k7fHnQKfeMJ8uTlJsK4pKEwhje
vBplobO0k5x4+wQP6IbBlXGHLdOuX7jXn943EArJ6pB72eyz0sPDOg6KIqN1mcbf
pig6cQvFqW1+jgAkq/eHXJ6MNRs2GvSaYYWFa86AOu4e01H6Kj7ZNFRFL6LRBsOj
FJIc8uZjj4IT7RrfO30cCTAK4eKWN7uZgudn4qfbNKg1aG3/J/QQqpCFEc+oedOq
/jvZPhP4OKySKlODkzG+63updTKrnNGXe1tayXwC96BLY5CmiS89MUUJmjJbAKCZ
rgH1gTz9mTmLabP978CUbSFpVWQEV1Em+xy/vKAYBkyTHBv+2q4FsIV8hrGESWzY
xmjuMBym+/bxbOB5eTrKKEIRsRQSYhxvWnwx3N9jvwbKcIOXkhaedqmBNwVFic2K
ofTdEjYh6pgcBEbbYkXuCVe+WgppRmnC2ZC6oojtye5+/LJARyd66U0J2pc9vRLU
t3UTXyzxYJNwt6kV9Tq72CxB+hY1WdoU1IwE1zNoSHQ+pKLMmMISEyn4iIhIXBFC
q5FPjf/stqOZOeZ/8li5nOAYL72tEvEUOM9YZy/3V1gPcBCV5ehMZUB0Efx+wBgw
NThdtJTJ9PerFy3AqhtIIQJ+9mHOZ/oghwG/6umGB/aY8lgOYgNOnbo4cYyhNgBg
TkRtV0nKYoxyuCsace18LX8oIRp8rxhsbBkMX5iqBV3Vh5CFe2hOZLYhCprLozud
9xv7m6UXlu5Z8aQwDDMKtuv72FSgh8tdcf7Y3Bp80+4Ntsd7X9+ITQRgdCoaO3uI
OOScnfNVAlaYEYl/+otD+bmFa6ndwaVGv6BrDZVVzihP8Kjq6hiFtux76KP5H7OH
1bOFEHHaRoL6KDR4AbzAMx6LYB/Gi4gYjOZDT4mgbVCqpx5QKjPIAFqMHdQuoC/s
v2Me7T3RR50KmH4isB3SGErRNyy0273pJo4uD4vB4W+MAVqxMltBk/2F4gHwCnR4
QBkUuzfUrUDmp7OVGTCxgvhWfa4ImSXQRwlhGgHdjDtby1CnwFVYLjFNnF09PPIE
3mewFhCflbrTL96SeWfKh5umFiUD/cQTP7s00mr6mjf9KeV3rxURhQLedyL82iPQ
Yo77aQolZvTagdeCFJropXEL4WbMMpSylrBNBYVDaiQIL+FkfZNNNOJzWqE2+maG
tkELeFiBp1f3TwnvPCDxe4jh5PU5W+d6JFIs+mhlpXe8H/WKPW4BxJveb5akpTjK
ZF507ZQ9tlZxt2zJaHNFJCOhq9dq6iVon7MKNCJkRIpkGCX/LS7T6epqfR3TqdGN
rS5+yxg0/2r0uYfhruhYrt/4T1m44fTEBJHqkUwQdTF/MdUhqZMiY4i1lPP1BIfk
HBzXKRr+XginLpX7/F35LVbny8o+IuHRSJi6r8h7AgtaN6ALk5Y6fImqVFvGqp8J
G/usPj4ZuO1NZ9UYOPqOfQhRAlorTOhHVuzpnvqsnwGdb1ij3qZqP5XyZ31S2aOP
FvJpXyyhWkSvt4xO8KniS38Q2+xLq88H7k0u3Zf9i4d8EKj9CztdJ+ASTQiA8QG+
/xkg1UuuJTNWDIoKZt8bPQV3Bi1qoi1dcegLpuDe3GXBSFH7QoQK1ymhionnBXQf
djTJLgJ9pOfm2kNfit8h98JhDfdkLae9GjVlZaniZEaSbNPaf+DtMYaLl2JyIdjE
3cHyjusaY9Lh9gb0a0vI4aoB/dPZdC9/OPjtkb3NfbQaU/X3Zps+9DOFwYmAI4lh
TrBIimJQEN2FaX27TeDDrlfV93qWNI/GceXyqxKcvjHC/1XjDNW93L1kTVZDdAb9
5IOFbqUAFl0LhACEUPL45N/GSv4VEBWYkTvMGnh9nb+ehZb5A2FSjjPCwjgo9cpb
bsqHRCjHAOHjcisLB5D1a2ThMWX5chIHTggUB6wYmUi68SGKr0rFcv3wGs3KTBSb
LziHjj4GzASkMdodLuR9LNC2Yk+BdiQftBfmy69aCh4ZYk0jJS5Qj22x9hVxXqyq
n1KIH2ZIQg3Jkp4pKFhDUv3zMS055R/wZo+3fXWrk5n2yr+P3rPv/C3vpbLBlxcE
AmWkvu6BasMCyDnHQmrD3GHGUH8Cknz8srII7bMy8gvbhDn1dk4nRx/EvTnhwFMD
5yILvxcIaAdflqYdR0Uxx/SKIdt42maJmxL0pf5ahxTipBsdOGU7x7ukFX+mVFQQ
Bd6Vxrn8NlauKYk6C510FIp9X14bZCyMEEHvNEv1eUZACAB4RWCbvhJF+KTx/ENc
0swo+T+gkm05TXNWsrTq5QsKTMFFM0x6Lp06NQ46QmItIAQrkchTnWMunKK2Xk3n
aZETNlVHcLeaa5ecnb86z23ASa7EEzc/xfElMX/LEq3kXhXhd7M6HZmja2G2viOt
SkQB61p7knZ1XarI93bfDMTGd42sRsWmvjiJA7PeW1r8bc68WEVogHorcHzUKIwL
LvzUF0xK727ccmaNEIZGa4vuTThQ0/Lg0O6j3UDzya91T692olc0kIU1B9R750ft
sRqdFAHTYrF7rd+yfXE4K8a4M8mf7tWPDcOUWcfLIsiLpIZGS+BQaNcfPGa/ib9S
L6irMx33NeW52oDFMU1DlPWQAaVlu2EW4dhOR60a3/TkR1vsg+aL9DZ+8BS4dsAV
vr9AzwHBLkxKCX3BB0Huq62jvzsgkFKnriTxKK8K1NIAK8ab9jYYmH9mWi2uyqvp
8wdbjrSutTh/cBsUyXsvFZlwtEc34xhp6a/lZ25/CKmeFQG2P4Ob4T++aXNJEXR/
bVeXsQzO/GITxfBvIk3FhquRuuNYc6odGPpCXANk3tnszS53ZkG1uzGTny8/4uUr
47eH5dqrCrRGaIo35Mdg41UeTw5ivDNa0Kt8945LrTr93trOobmb0MVa38hEu0z4
SI3RdLrCFSA7dvCRKn/JshxxTPk1ul81cyi+Aqzzezc3F8kfVQx243AUbmee4M+6
e9nuMIV4CLs+ZwXA1114fu+ZsET59aH7/g1v5QyhSaAxVVTfYHJ6T8sYk+lTVLOD
fZdq+wDG61xO7mmTE7s4SRsOytn7z8oUJItRgwebAFe0v2jacpHGMLZKHAinOPmr
StGKqrfTxxpQ4byXrYRjFybJSl0gUfFKHaDAOd7qbs/5WSi2DBd8xlfqaqxvYPxx
sn1rcnXHH+75onQkixZprl7YOJtnu+P7TN0W0tn2E5nOEYM4uEiWOeTVFe7OOEKf
gSMWI7Cl+o0QwVz7lKihC+XPX94YrU5QEldXNZUJkW6pKzMupDJVboKeoZwaKfiB
gtG5RDco+P5YP/uqG4V4d3U2WkyymnyBlIGk22O8zGneG/ire66vo7QLdKsFm61h
PsJyn6C7jAWwUAk7HkhEaPn7BBKRsdMiqsPQaoRNHlRkdpAzabVe0S4ZhiEd9kfq
52fGjBO9IziNzozrkIk6pstIA9fQ6HvgrKgJ3Tk4YyC7122u8RgidkmZkCwaJ5If
VONWO/w1p2rW4AxnU0tpIwP8cpNYmNjtMb9MzpfLPEPr0vI+0GBmvnq4fmIU/WCn
nJJ3cS9phxFdd61Jd4QqFE1flBMfnaTG2xp3hK5mpbEjzjg7qBveyaE87VdChSIR
oO3zwn8lv4jq4P9sfIFMweIWGNgj9Zgq6WpSWJTrCSgi64KQcLcOM+GE4RIlHJdB
sFdZ1vI02Ey5PeZN5zCSci1DGltXEAxWWN27ZOc8gMeXygttFma0WqDKJz+NP2ll
KUuyaPaayekr2AWBKq3PlFpXXkU2Eo24VqcNbDkOXi0/3uWiNQHXNWdLInd7A8vS
GhaITDTHpH3RVYRIhBhN7L+AqDYjN5HTdFnLx5y7i+/7sj+GXz6sYST1ZzR5rlc5
jJkxbDfmkKd3vQ/JMNv58abILOVozXOq15D7dm1vmEMLqJHgsALBsZSFeUwXYvwg
92l5lzywDFE0yTMWqXTfu52xyFVMR1DCjZflQ8HMUvUCgYh6v5CeVx53xTSU06TD
m5TU4/Ztjws4L1uWdwSHKgGR8wfZo10Z2ixlRQdMiJbkxiQLqDAfSHPh4Tc5EZfY
FzHDxmAbxj1esh6xxRAZXrD3ZBYV9PXTxGWbMnJA6DDk7FuHGUaVOjsACzyScrJx
cjIJItFBptdMfrG8ky2txTRZpm0i4QGTkUz+xvkZadDeRVFIv+kgUP80gzT3Coyt
OODo3Aj3XGHSKSwQvkl0+FL+hRem0EyfoikQYB0qTZZKh9oMmwyQ2iXfLoXmYG3a
tLuqUGEvOfdJxkWcF35O0xub3a490LofcrpxO3UefE1MtKwuFbD6YIZ73wpIqW9h
OY1GSGpUREHKL+RCrLVMD0vnRDeKrbvCVf7+670L2Rxqng07GN/Y0Czo4fMQHT0A
hiE/HD70HmuZ1Gv4EKNjIYMGXz53nIUCJAgy+dOTuL3rtZRZ1n/f5+iOHGp/B2Qz
jlJwLL0pXqH8LanA270fGsMU7ZFWaUmxViwNW03ME7dH2hEppr4SpKI3xQHjMX62
t/CXU8gcz8QTYF+uKwCOmS6cUFQbbcSZUhuIe2HhmUMgdOR+zN30xndPdZaylLAN
ZSbs3PMx+WNKpTRaXnRL2QufHehahbo5qaXK6ROdMB/GPGxOv9Gm9cOTkx436YFq
JU0OSCBbciqYds1QC8UbzEcFNkZ47c6aw+XTkVUSPeJ+WdK2zZtTieYyI0lu+eG/
48TU+k2h4fBH7QQZDLiDsTaVnxrZSJZeR2cyy45gkTV5JucjBjVzNQ+p4dHoq53v
Lxi3gBoqI1sIXC5GXBDzklOxfVNhgnin9y64uwQQGmdF0hJSQ/x+BZIO/pjXCgUt
Ln3E5quanHmE61+hJNWdlsvZKbP+U8DAQWS8cEOM5oDedutqYYmL6whEUjwT8WLa
NwonRWkYh9Q0rGJ5W4tP+EAHBpHt9FsKO0AI7Lt5TZAOhzWWMN1D08LOAauWM3u4
7/jFDFdRygt+XpU8D6SM1/2hqX5Xps47GTFNLeyimcAdHqcjDTRvMyIT9uISx11a
LZighaF2z9k5DgHCZBHgB4gVQoNCOdEazqjQMWbjLWrLqpPPvYZOpB8A9kLVbQ+u
YBKmGmpR1Kl+/gE9ZriX3cqhAt8lUyyWYQObUUMMazfjZ97oJAJgL4zZFDXEBjEq
+Mgym3uy/C+3SK78XtUUJ9dzRJ/+jxvWQSYGV+tmMV2rtak99jABqsPdXR+IQiFU
9Ax1vAe1yc0tpjEx53VMTQYYnJbq4Q+DS/TpdMSeFL9w3vt0dfZhCquOQQ8K7bhU
hDJoE9hugYiPydmy1ODyUaJY1A0Xl/1nFmqAfrgVuCnKWiBw5idkbAgLIIhMu+Vm
k3E1mcaqHMairmeFVvU4PWqU20IXay0rRzZDacZkR3fWdds4w6xQ7bJARH5TnC8T
BZUscS4G9Vtf5JwhD6rmTePEQuSk6H5szRBAId6XG8GqGDuN2nMIk0tNwDblXKu1
olJuU5FDYcAn5mYNJxNSkSLQZUQR7+/+U4INsvI9HwdJvEPae9cp1WHz+JL5diGY
8SJKmKF7w65zvLj0XQ6xJ2k0pfgJmyI51REn2vRrFdSJMHkkeDr9AeVJekg1PZtP
ziIS+BLn21t0kn1d1wdkRrOtjOLgHPU4X4ktyrZZpmZ/1WpmsM4p8ogOxUAGeozu
tWoVRDRTu0DIyehFxcqkWhAGNk7GhoNrLMfJiVXcNN3jAV35atdvOQEttSq2FXxu
dWSSDccMLK6HRbg0Ykne94V6xqOEptLci6wAnCy9J/Qp//S0/WsTRz9bExVgkA+/
5AQOrHmo430PL29GekiWD7IEJxtovTvEsXp4uTAb2WxXJ0TxhzEGjhNi1Oq+/ztP
mTdqZkseUcqSwq0p3qP0dhuuKjJ6tEtZWv/R84wEu+vLv/gKp5sdAiOd2hE67A+y
79e0qTKzJqehLR83Ls0TeHFl2tBcMQ1heD0tmIsfcHmCjh+2dkLGOydk0M/WxB9M
R3rf9an4Cen9O/b1lIuJVO71eqexvriQC3zL79hJd29LDmigjEb3ZxBJ3qLTQI5S
olk1Yi4P9+d9xpbqpeoBwZ8ZHWKJOFionaeoIhyFFyQ1NmTRrvMpVOEpHk/zEQME
CnHaUbk6/rRDQXCPTi6AxL/yvpLXi46+FK/zfy/r0FSyesheVNrGpXOq78y0Orpv
lpGMFsLhXZJx3A/FA+Ffa0GZ3IU7cmMgRz9gCAN1A2FRZRuxmLpJjyV3FErHSBnb
9PA1ak1HWeXp7iNQ8WA8sGl/5HL7o30eHO9+uyz1MUyY+/vDwsgdMrFfb5fA6KhA
KdANRIkKNOngBQvf+z57slUVWb3Cdh/bniHeK/vpJ1BVhT5pgdoDBrEKyIXluC41
O24j69T03kf/e3atZ1isPry3mQzylsmJ+yI3VRsInW/7b8K5jkANq5F0qQJr/hnY
zepmV9aIzi48ENEAGaQqFJ1y1/3wyPhPDCQy+yWoetNDogNv70HBvToI4T3x+lG2
asW6rjQ8EFRXvMQnx1kj54H/ahMKrpXKfQi5Cp9u6VqVxFiZSx2dQ/4robD80/co
Jn39Uf9oBIyeiJ9RO3hw378YfkE6Qy5gfKxTLJzeIe/0NhrSScchMXbsaI6e7dEA
bfF63VdehDhDKYC4swv5R1g6P8e+R+gEDS0nYSXGKfC512fjiQCuqjP6nlyBicdc
VJZrVi7TIWRuxSI4NTgrpeLV2FrhSq6pjq7XJimjmbOcRRCLnntjLwNg8cqnEe/m
tJhHZB0EDnzJ1tPachK0uAISrO6kf8S/4gmI7D3LPm7uMk94WNHUUKZqvmqugxdE
geINkXyjP8AreQ39rfbQ15XrZMPekJGrBMFJmpdy7HhznSgOcyguqooFyHmNLB2x
QeG4ZdUjgquIQFfrqF9DIInUyqsDPB/Td47B8yvVrrGtGDrvDZrvwNJygs83fjXm
pqLKNvIkl1NGWmiTh6jT/WgZ5RLtbGTBxSKNN0jiE7juVEoS+xoFS/1Jk9L+lDzZ
lNGfkUkD0yqsbhUvLgp49bDotb8NBTBsIPtqOZjN1ZveWkZi+0JX2FWrBJnGj84U
geusCPIhGYeTcuo3a8KyGSEy7XaNs3Aag5zvYzUBql9mQKOHrZimDeTCRPK6epSU
Cg1s4lcZoClgFB1gR5woOL5fxrbvP+SJcUlSFnXs5CgQikOWuA/dJhjhHs5/u1Fj
oIXuPeodhufv9j91gaJyVwOQ7YzDU3seigt7+bjgxo6sjUVR2l43/tGs5fx29eyd
d0m/LP2rqKNiEj7LwUEn+rA1JzdjQRF1wJxYcn0p4vPHtNZv1b9XPNaQer36+sfC
TRen9Voh3BZr84y2iKLHeAPnBwP7R5RZnTR9Ldgl8B1ClJZqP9nCaZTZHlTR9rfh
frImMnhBvvcJtcMnCZVwS/YAdh//6F9qikF7SlbFIm5AiepS8EVGGyl6SftbL3DR
29ImDy/O8DuSAKv1Sm4maXiqtqjrzt3Gs8spuiNQVvonRXbz/w+Q5FO6D8lFKrTe
0zRD1o2XKgaaQTJBPPIiS91ejS4ATKXGVTehoxigGMVIzLA47zqmuzPeNLinL5uc
ZXiZPvc8DCt3WRRq2A8LuWdO+2L1BjzYBHfXsClDJvC0BgQjozhLzDoFjHk1kiF5
xm0JVDI3UUmrsuSaaKN8UoFLObZGQozyqEwffjlxSAPpOWLvxrMAGTTCKaH3Tcgg
QruKeNmbeA1AeIm6S3DeUpcjjUGi2/xUzcPKojpyT5jb60vs/m2O/9wL9qgVtHwG
xVBEjLemH5b/8YGBDn/u4xtx17z16hGPEDkCXKkL8Tad710vWsF2C7V3E68M7A39
Q3KoqMph3VjEwK/sQ+wgYFRkIBaNwd9XI6aBbwkCZGxmYGJty1mxOi7p+CZA7Kpg
FE4n116PEnq0ggOlzLNXXCLiUiEUusPuowitKb9xXDAAYU/qs4a9H0fuFMLJ7NOZ
6ZK5JAyk9+LVIr4y4PF0m46WcL2om5GTlQYfvY0dPOivCM6IqURgNOhQ5RI/KXRl
HXfj9u9BGOxkxc5378QD4tItPktU2ZK+eKg/AEj2x9S+gyK8EvlEmyYBPMUxAoI3
ufUPgm/NohgfjhVL3vTQeDtjjsPDEU1BUz+Cju56xoX6fD9OMIMEiYdgWqeN1zy8
ZpB6tBGJZ3Hm8aCqF6bWWljwCwqPOtqxcix/TIFEdUOEAEKRJ/4nVk9b5gaKxL73
5RR9G5nsxe5vqcAMl9eTP9i9YIBkg3Lrw2uQYe5CPqOvGQ4XcrM4HHi5UM7rCfLG
BftmbGFb4YRV/q93lVLfPsf9XHpyeuvnhWUyPlDntW7VG8r/EpIOtRtHMgoddX+x
46YkIyezxL00pSQ5ZGEtmd872Xn62rOh+sPcjnX9psk5RkoWNI+SOPzasc2ZFBfA
SU/cNqMVwSDJP+3j7xyb/flUCwfZb44vT9DSi8OTRea7AWYxGLXYfxK12wZqVyJn
yKNTHAQLeHRuLkNeBKHtelWoFe/Bnrwyl/dz2ctRm5JGkZnjKIaoMQzQNsJDB++P
MAojOnCqgc4hOgGPX0yNIzSux62uz5srpEvOLTdY5/E6AGJNmEx00PoIIT545CN8
wHtdaWvRLgbhqt3CZylSg4FSYES1kuxe2yQHaUAOoTpOj3G9IKoVfwSNtPp8aIh+
8CYDP0NoOevCxnJcEO7VKjFOwFr/3/5sGMNkxutKJXMTTrNC6Rx0F5J9rfdvNMKv
uRMuECq683K7iPXZP9jEzR4bm6BtDnVeP9zb9lc06FXVTrGzB3w+dhoHfDHynv8R
GkZstBRcN41JcVefPZITH4rNeM4/N93whKVnfJ9NPgb8SkDIM3yLOsxMhgOB9KUZ
c0Uiz9raX0I45z2KTPY8XqK9EQxIywXmyuhxhToVVd/Y1rYuGATStyBnwCdC4H5e
//fZ989UMXGYxhcWj+P1YirnyS+XUC5wZr7URCKK/4oEr9ysaGNeK1sAgZUigXDv
EbZ1NP/RZGI5phwHuzBipIX0pcvXLY8fOQEylPmDKJClVry0alvVgibuw6eS4jGx
iXrfsrKIxqPyIWeIJxAZfXc5INblvXfuOmKt/UutsyjDIp6cmwjxOH4an5Vh0GqJ
j51gbjJAgCbo0l1P5e6Iyi/131RzmjTI5qJ8T/4iub/0pWwoEOCc5B3LJlXR+rcr
NScXT2cW9WG7GvH1nzpgepJ09hq/mR/lHBwsVjlHyh0m/Av4dimFq4BPz2UQyC33
oSkIQNNYSJ7MKPe6aLTU5lRrMG3c+yuzMlUk5QJj6Yxe0QJLM2bpKfsN6I8ihifd
a3qN1r5y6hphHpbz2ZWh650q8AcC8zgSTMdYnTV2NSf+C8LyzCH/eP/oNbL81zJ3
cqjKQTJKxIGufezi63u8U4vOwKit54z6+Ql9NljE7NIx2+7ghqTQ9tqo1OzZIFg6
/Dp7rfKI+IL/RFY/GSQW9lNK4AKGapdvFvrT+wdSo2xp7t6tq/BH6cVLBmfY0rna
QMxfSlt2x2lMl+/uR/Sdd/wMFm56V/AknUsuHCzF4yVr4AlF1BgIl+fqD3e4MHmG
WWo1f81Zkkv6HGaY4xKND5C2v/9702jOszPPIsIGB8wHI0mDefGP9AXbKSJ9Yu3t
to/KWHEJO06UBdZ2UqYnExbBq2uh08HLjhiaWu0GTh6K3yNzNXdIkF3Oq4DmNURs
dyOEoWsA2LMC3A6WrsZMJKNom5ZPVe9Irzv3isDAzsxt561Zozvf66qVXOSGGLvQ
6EFQ5DrOVCv+4egq8BXFL4amICbJC9IM1d4+FtYRrvqVAd69mA2WZN+0g4hp3ox5
PvHetF3P/zCa1HnJ6KBcOCkV1W283kDLdztq7Y1GtPyu8aeS0e1iEsxC5B+CJiO8
KkAslbNy5ZJvGeZMu1os7wzmVDNz0afTzWDLVPQqCY8T2KR17zCJEVy0rc/4pjSV
ttCMNd4DvYoa2YMKmFDM9MVb5EnymaAvZ/n2MjCcqt0wWa7DipHbO+I0Fx4JP7/t
aQWxvyImbG9cMdjqF/S5gvZgvQX21IiWgPsXs4lfd0FYvVU+UKKI48MqNmW/cvVa
KdHi/0mcTy4lV7AL16L8FsAZZqZaZ3vzMdnLU6hmZ2XlxnFyEFJ8EXISzxOGNgLi
fQx144xWXzikiwTFnuTyG062LbtcJKrNRdAnjpHYK8mz6YxknG7B2Aja61cOwoig
b2hwGpV1iGMT3DIAUENBRXWuAYAOJCZOql3vhJOVTZ4C/rLrc3EU3yswb91OWQM+
vlMBAzjoFtJMgzD4uycRkgY+tqRTaBN4W1OeJuGkqrbwVmLJKcWuAtf1ny12wbmt
NgyQlz1Sb6GHURTeYVN/+nTd3MFMj4mftajFt4k1erPGSRgtlNsMXLN9UFkhM+5G
EGz/+PSWwYcPSWI8SsB7SE4b98dht/tINrqlAyksGI45gsi6ZCs35RDRlopXJ8M9
OQYo3Zry+WTG5CmkCwtwAxdtE9u0iuYIXhNd9qkwpM17pK+WkzuT0BJEnvi6MZi+
d1Iw6eaAox3cRN7VOd+6H65YCEkTUKbtrQ8GLu6cmJLTf28pVimMonwMGF6VsKZQ
6YnCXZTWATDsS9/+JVGEoKRcHF/Dr9wnxhx/gTWogDHOomJJmhIYvPWE+2NZt1l/
wcGSHvPxNL/jTV5DPjAD79GJRvVyxsd5ySlPusSQR1jRm1PEOCvukuHxfZg5+McF
KN34A8xQ1TkEFnjFimKwUpZVWnEUfAyYiFYOFnuRkw+qeRApZB89qIJOsdFYyKzW
0FWu+aty/ERLbVXrfR+99Q3hWv7gg3g0KvMB9MXeOEl8uCOFjeW0inLusOeGnw3G
f4yJckPggRkuV6MXMrmCJuUzau1usWYW717cs0aYepfR+3z9ioGgJxgLvvoMtKYW
K/fVGIekncW9H8+3JP5SlxbLgd7U4tcvo5oV2G0Fhusxrga2fI4rjZtXR/HMLM3R
WPLzDbiV9IBuYKpGKOr4qn4n1nuoxMq95Qde6dgt+ud2j3tSBBT2jmfoUW30c4l/
2PvGby2oKJ+iCPoiPsvJqWhrgawaaq9vvb4prga+Wftsbl0vg3NgL5VjMaTToj8v
aA4/RWUk0C8iXtgXhGTT4S2wfQZsQ9nWMKwbuJDrMg7dKPyDmzH4FnERTSmAC7yd
b8L+jaPIPJR1rNBRKlk7NasVAzP8hu+ViMgSU8xn4pq55h5U/K5rr6jPjvzh9GLA
mwJH1MxByhgfcbzuYuTVDFC2T76sw+HiTXdcTL6KBPCRHt0RXlg3FUvjsE7aZHVd
QKwT58512tBNbmDpwJWJBHVbRiB6fBJZ0heOwMekTW+LWXiV+lyY4KyNooo1MPi0
XGKp6FascEezKE2N5yS2bgaShz6h2GWoRnkrPR91EGG/QU3kV5xiR7Y+DNZN0x1a
Jnwr9U4QZ2gd+ZwXq7wlPbAh1moGd3MiNL/mID+tFn6rvRLGWA9NXqfSQm/SgBaB
YQSLqtaTBOl3W4pIedzH77qEpB8aE77xttN7/TXhnaEmMVB5yA4egYGjsNr3BXpG
Dze/4wUNSC2xJyVJl+F617wOduUXEGmkiZydMYT19i8Z0dbkCM/LG7VmkQpjPO3h
8DT7FnCfpxdC64XQM+vvmHnZbFgEOSOjz0jBu3a/AFJDpvrB/c6r+lXywvfhrr1r
J/Luos+iHE7u2Sas1HXLXkocRXyEI/DXS2XKFQqPgz2FSxJ/9A9D5b6P+pFEEO3E
Jn9ollkv4O5vL2gLYor7Qq9I4lbr3+PrHBLJmpNEeLdbX80OhY/0Tp/mW0yKwkez
zfC869KEa1WWLw5+9C71T/XH+Eqo7bsSuk4GWe/iTxClWG+EfyvUQIDc9Cg7Ys1W
nAlm5fh+15hDM13SafTu8HbslCqTSMOqG5TbGw/ALMzB32QxBUNO3lEXFbDFn/yJ
C95BpT02gfEBgyiT/9XHv26EeX778YKJMrhLNaiNU+uJ0RI+c9RlimVWHFXZaH64
AGEC2xODgrFYjTHZZGCrdyNA8RvIRkExFREsgMGZkpcQ3SMeIuuSc3st5szo+CUD
WQIeaXC4QlPmv8ipw0y6NII8tyMW7nrfRXkKE/O5C5Xc5GS7mwlyUHMbnkdZw1y8
0cBJWDv4VAohCMD7ob4kU/g+KsuMWncNauemd4u8ERmzKFCtXevulrGsUHq4xf4v
p7cF63i+Mnoy0x9bqbTXQs4NV87m/0W6Aozv4ZVzEqjcJGAzT26HoFzeLoaF1qPB
23bdopg544in6wJLpAjx2BtNGaSerMLUMol1Cd2en1fXvOeGjdauzsTSIwk8lFV8
O8qbKlwIhiDuSQcOILjnAdu+Ji8Vr5vwVWNGX2g5B7Cz1OGp3U6nDa0eu+m1Yh2g
1CMlpadJZ53xCs7savNmkBphv2xcAVcsAtJG6iPqaueRGm5V1wDMbccUxOspZio4
cRL13LclHxr1VJQS5tdhMeSN7q0HHGca1WOPlBlEq7TpcrPa29ERwErC5OquLYLu
j8q3cw0maFOq53TbffM5e9XS3/8Y5lnQbGKGyHhcGm3Xo6m6L9aLIVUjnEkcR1VW
6m6SByEU1MCNgbfMRNgOWiVKyidsUKdW0xbw3IhdNUjcGltBD5WieyLnaFmUHG+R
StW9YuclT0ASm2RVe7l2IuCPSTYr1cLlHUtq2NMVhBrmtGjnKlaidCzsBSIXw5jk
t4XjZunmiCh/CH7SdNwdHiesiNg13Ipd4j4wifKaGQlSPxYw/EJ4nSwSrJinGjf/
k2TzkbnQK9hvnXxXZeren9z+5Xo5R/hr7tygo7OGHVP7WqRBemPvrBPhdVEcTz/j
+tMU10+URkLLJbJT4nY6M13v7BajloBl9pavhVy05ib3xGVMGO81vrlxJ5j7oChF
EM6G+Oz76EiiiGxfGq2BdlkqSO1ZB/saXZDTJOKHT1qLM/JQ3E/o6kzpZE6CzA52
aRjJJ/62lTdfRWuHzbwGctP3xVCmME5XPLsAgdECpLKhzQixKOzG91p3EhR+/RMt
rLCAN24SA02jZxK0nnJRhKkk9z5vv7EB5rlGRNbiiT1gvcSd7JyFmIBS45N05J6+
juWgS7YbBu2qR8XP9ezPrPl3vZfyf2H6aQUWFLYY+YJ4Je0n46q3IsidkQjz8q+M
a8Yr0or8/xpJzo+5JMDVyO1ZBTsctV82f662+8dduDp6jv4GH2xX7t83Q3uOsuAo
hJRsF1USgJ6CCIBcGWGmf3g+f8egXeorMf/Xk+QbANaOH6JZ/iwhWWugdKAUxWxu
EhACqhVKznzu3SXOVtkNg4dYiFnzJiMsQ1LWPANvn79OPqrZs6NRPkpg7sLr5JCN
KGkcoqI2a0uPO9M79V5NftbvWttFXrJnDqOHVjm//1bvGt0Eum0k+gE6xLVIzU+C
xmnuRRHPsCj2UVtJ2j107Rhm5fgqsWOR/+Udqdq1wgBt0PtcO2wNmcHvAPu/0i1/
zGUndrTNVdHHqFRKnCjga5xZ8vVXVG9uqRc3UxFA1aQUg1OBtV/9e5LN2I5ATBNB
x/0mm59vptcrg0RKA5Qrk1poqLOc8VA21xVkjehGeSEmIBCZG1ECw28ia8flMBQY
kqenllFd13p/GGd+gisDDmjJs4vvRJDdypSzqkUj1GXhF4Djmr+CzwGb1qlQRudu
PJRifbM1E2+Y/ZglR03s1DiFZVpyx5wAQVvgRZtfaoafOpRBv2ccS9olMJ3fSAXU
l88ETUooKyEdYgH1xpwM/EaQtvbMfgo0c/KWAhiGJbK5knrqYw5nS+LW6aUPRWmZ
466d4JkmeHE+YRvOEtDboqtzwGzgd81ZN+wad70gCh7lZNA0OWzAXJ4UihDW8YJY
olYVsT1ab7yrYWFisJkVZoCeGevmUzZll9jugVAEGqiciJ44/HBSOU3xdDbivVoY
zN3vX0tHlheLMExA5Ko1qQZbKAAP8ACRagQGoXddDno9PUwA725WhznGzb4Yc2wY
zqkgqDGq+mJYd6FRvuGgnRgS4044ocsYkzqgEHkv8Nsxoi4lubnuXIVEkvmmEGBu
pYUP/U/Q2LYvjhZvyz4yans47/xnh/K233o8qhpAOALJOz6Ol1EQzIzdFvGUOvIK
SXQPa/r6wTs8GFiWyFvywAHSnnn4zGzhTlKdQ1beuIczdwG3OOu/f6CX0QjpPngG
ciMBQh6EyGlF44vsQbm56MTKlAYfUi1g7PzX0qgLdVJ9Ny0K0sKe0I2JMpvxohQZ
m3CSYxAVcEMVDm05ejxJPKQMSRYVF1CbeFhAHIFe4Ooeyxq40cZ3VU61gL8rjn0h
Yk+9rCEDQUbAhSH+YTJx98fITl40J+JQse9zJfI87y7W2BKnhRS8f5MIHSv+zeH8
J6Ip9QODQrt9hBt2EYjB3N0V8VfUg929avFZTmu7X3wzRGy1uuaCKvuW+Vl4rEha
4qt5j8cg1+0/nMYiq2mCS1ltL/xTZmQvj+knlxdxo2W1WlI7CGtd2urGaWEqZJU7
LVisnDODyZSvmB+fEMwLkm4dH8NcFWTg4SBeVj2uSbzLsBYeoKcXH9W91lkftm2j
ByP4gzJE55qP6ScQ9kMvzNDf2fbA2aIqVn3wAZ+R4woRJmcYIIGSPHgwV+3aGcdv
ACPUxWvvXySNMutuUC1+IdSENlRQdJMPiunTOyLPoPxZPfOzLJu7hu0LiMwpb8Nc
G4tJHICB+uGleyKGzuMtwVRrbEF8fv4N63R/UMR4i3x5JZjwGDMUmokG77V/3ZKe
Mfdp4Z3nmGYEY9AGphoVx/q0gJR1CMEZjo+AeXwPkMLZ+E+kOfWyAwlNTMyV/sEz
uICsn0jBwOhea81muBpb9QBI1MWDs6wsXiQe9yqpPpsEjh6zQhc7kwdJnnh19nUk
cyD2JPJ33x7YdiyzuNS5Wiz6ZiSqBzT8gwpayKXW6wwkE6x/21PDWo9pxKM0bY9o
HVN4c8IkaOXivx7e0g+lLs8HHPDOVH/NGlDYPufkCHTmlwGzHiIH4Q2pTZKl/aZ1
FdKG9uVeciV9PiNhvf2LlxDJQRlfDWQvcAD0tOuzo+CQy5JtSVcPLLlHwYhnV0E8
Hd64Paw/OrBVxasqKUxaM/+tCTAPg9BZVbcNwrufYe0zcly5NS64p4EYNBw54+bJ
HVWJD0dM5A62oqXqtcEKpCqgJAbSv6K8QADfdBvHN7TPjop5/on+OmaehD3m6K/5
jos84tUTcYASdQIXc0eh4KI7yr1lb+om+OydYe9nKgDMRB/dGBNmn5QLQIcXwdPd
Y2En9/b/Dp/st99J9D1e44v5q5u9tYvEYDSWo7h5YvybRAY+mpODxDd2iBjupaYX
cQuiT0rtF9XmB+IhCYQNESmlu9P458co0ckwcln4+1pQTblYIwRnBjyHyJjhqpyn
oDySIMJR0TTl7Uvri177A8GokPsc7ZSghB+5KIihpV3YtAfmgEpcpHJPOsVw06z3
qIh1qQEgD0YKRnYPm0CNjbSWQsPUCje3jqdq9NpVv0ibfFOQz/1ztRMzfHfSOCkV
GDbBLpvRIQOhdD2vRHpdyxyqXFrKFvof6W7ZwUvvYg3zcFXSQo1e+MllgccbiOOy
xMmgd2d6eFznp2Yzx8SSddMjq86CNjAXRD9yAHCgIYHT2yHo8OjN+eJmXvotM6lO
LnPIHw81ZvfBEqgcL+XULbRdTHZcbaaUk0nGSc1aNrwanq0LpwwCeOJoLHwdx/wG
HQ2OnPIIw2W+VMVF+SVbGrFiZcULsQVeedh4zvgLURCdj213buklXVkAqdoNQTpI
uVFAjwmqLAFSPOsTHgbeKeKwFt0EI1vKp/4yQG2VuSYUDb80Siu74oPSBoINL4nS
CmWbzLxN1l2iXH2OknlBPkqN/80xcQT4UYP7emk/24pJYh+AGQFzRygs7grMfyHf
QnhabVmaeRURUL5oSK+oPCl8jOVRE8S5P5wArUzZugi+ziMc4dhtMHFAoTI9xa9/
hj7mQpvcR3I7SkPFfRyt8aWJVnRgE8WsOIuiqQcyK7GbT2xXdYjpTvfABbG3Ouq6
W1m+KWHdz4uudr4+SE2y1KW7lhPAAVpwE1Mwq8mR7S2cq83WvIo2ruk6K4Ov+ac7
9PIAXHCE9C2fI5sXkx+bQoV9cb3dBLPp4LszgZ0MxqhcanbQF3DbE06QRZQhwzZH
R7vPDlsLFb027JpyTnUWOO3ebaoS0Z2mLEOXMpy49OTfv1N5PTpVRNafa2IVqbDa
J19N6N01GFG5NVfPxUh10KNAULE3BXlzUMnRNLhRQD7uVJAipemZ89CFBL6pCElH
+wIZeY4LazU1dieCdzX+2gmlFLxuH8U3dja8FcmEdf2WDQ2eVnLT5uywZupOsXyE
FzPHO6CK6GIPDeR7MHjyhYVGmjWD1yT1tpNKwiybe6YZ8wWqDWvlBi/nRTfyLlHk
mxdNHzYS/y//Wx++87zg4ccwGS3J+ZSLlXo+pvJ35fpbQyPoGGDUY3See7UW5gxQ
9BWDgi1Cj80m71uW7Gpzs4J16Xx+6YEw14ktAyCNvAtd6DaawWEo/CKv8VBGAyQt
29nlTy24JJzR5R/xq1xE0COCR5TA5PlCOWNINpDVe7k3hpZCsGQbVXfZ4BMYKaEA
DD53RIHoSZ6rf1e8vlY1a/PY1MWHx3Athwip795PuuEuzkBcwc73IuqrSExnG4f3
/GZLoNkbvYkADplxcP4dgfmj6zGKIxPIcGIwRCMELjbTgs+bjT/8XOouf32IwNA7
s6KCVlajwLXBooeXONU5CWxrV01lguAFQZwNAL99IQGGUdPBb8JvKuT5wZz0683y
tvxz/jFo/j28/XKq2ZpV/kEWOONaOvRCIJS9MDa/7q9qQs5dqOi366xUnA41UfVg
DoOxSvFStAJqM5eZx0YMvqsETBR6mJryAZeowt8wRxaSrE+BjWQM2BJeDU3y0VSi
UdH+MfKMZjVdcfaDY9cPbI8nsH6sWTj+f7gORdNXzGYLpZiWTuAUdlmEW2zE206M
frBJpVSyr5pNDQV3HlNq2DqoTfx7jjwMVuoK8ccFQ9C9KtFrBhPXE/swiW7iudqY
TOcsVyiT9KKfaTKRwLpzE01mnnBHal6vWmIEZGbPS5CNhsFrPeoGUGgZaDelzL7M
KJOQXGPVG+H+6aa542mX1gtA9vO8UreEtw8SkkzTqPt7HapgZ9+JXhVDA525qoK8
Olr2rmVOVeHKM+Z7oqlMXeP0XmiKD3HLq8vhLq8AvSypPTxNAbfOhg6kfvdeHTSY
BCo/IAyRBwaqElF+LY46ldzmQl9RAZ0pPAi78wwTzOJD7gVGcCGeZToVhN5H79O4
ZfZhHNNgYuhyRktVrMz0Whi66OA4Xi+q7c7AmJK7+eUPzS8ek6ckArkBm1m6KT8v
rkSbWqvnwxw/sLW3qNkFsUksBgSHl7XM9wjJzkJD9N+zKr32eXlOPKKOb6FZm0r/
4LFcY3JQD3saFvX7UzqjQ/BY2Bz7bhaZkYRmQz4GfCb5ZJn16FkHNQSSvTB6VuEE
KnJ2sy6vy9e01iqZOoHzJGscwKjxMrzw/9evUkUgmGk/3iJl6eHpu6t+EXP8ZucT
4jah3XukIwQPYGwoEE6yYJrO/74fItEvp6WM882bxr+FS81ggAXQb8b+r8vJ35R8
yZLCFrgD1dP8D+cRGR5LB0gkYGT0w9Ug3+XJIzMemCnhT5GV/3MkIrfpKngXPx4A
TgRc3s7I7e4a+4Tsv5B6oErYRyLWL0DskN4LWOQzYVlX2A0w1MQPa/xBZO/5eM64
1nMPkHrBGO7jSEST+nFoz8F801FvXtqHZKUaACL/mBa9rg7XLbxFpccFVfLfClEa
k1t2FcrA9+Ofp9y8jJVIYXPZBlqbUI5ms23Vut5UKxuFiFHDVrhknJDjbv3AFPza
y/3e4t5PFHehGH3zWi5XfQ9KjBPRmHhvuyOWKFGQNyWiWE1Npn68MR3724HpHcaR
KryVYcxa58b82CtCvUxHwLBlVQXhiTithhMe+YTkGjXvOgIctMRGUDfT1pfascwx
ygD0YDKFrPqK5xudZBcUG+4jYgRAAnadOtudhZG0EksZgW1JeoeGWeYWydYQg/Bh
2g0BGcBi1hAdpBHqJxDCfDI6Tj2rgDgO8dDW3vhGY/s3SOcb7TAgCLHMAJHHa4pf
8wRNKSy6Op4mh7ZrkLMo9a/IGh9KLC6kaODqFB5Njq+2KBHf84vnzDuMYACypxM3
9+4nz9sVBIT+mWycvmMBznm8LpC/mQhZ+yFtrPCPftPitp3EQj4Pi5qdw2ZnS5AH
qVutpKQNaqI5fNdmpNCU0w7q3QRQ8Qhi78ZQ81Zjv8+bmZWO50b/uxkjIp90zXdP
nO4JQLHRvleoW7y/WBjInLvPF8KP+Y5EVS8k6vN+zODpGK1QW2SqdMwPT9yFyWrr
WcuzejseajBDwpTDDdFIbCdNPrVQr1TCWyc4nbhmrLfTww+x4VfSy+pyq4Aht1qz
xV0EUBlPbA0t/Vun5rOLIRPYXabKpytyaLgpFnV1/4H45ln0V9+YcVTCw9lAWMJB
WW55Vrg6myr5mkg6rXvCmsQVbaqW3WJ9tMmupKwaXm84fVEhnBrlDlyryEa1aM8i
yIbEAAjm1U+putSeHP4q98M1GmJygN2B7xqtXzje05TEFcwyc7tTzkYQvzcm/O6a
nSfLc/dB0z6amik8qj3Z4hp7yg6bvk/xUptejbrVOT7R2nq17IP3EMoJIKZpsGvj
RCSvHnEttQISZOKkLK9uWsSu/FE2WKB+rVVrBR7MafUv8Zh0r2aoEbr32ZMkG7hL
lvy3wX1utDKbs5V0P6Fff/oUO4UP2r8SCBtmLUnky4zW575LJlUjp5UbFrzScgXG
Xf7EnNx+jNioclRe5B9HodJv3l6rervKqxto/bSoOqF429CYqveQJGEiXV3JvuLa
rlV5U890Ut82UJHeoiO9M59ZIXe3V+xHvK5CIu7S4vYbRIH87YN/LNPMZTEQfvfr
/sVbZ0of3cqfcamYmZJWbMjXZsCjaYjd9SU2QXKMtTT8wokBRNWMgCxgwp3I+sTP
KonPfOMlIhsAi5Ep1buZiIkDYXWW5w51CqYKSXNeTjMgxIb39/LfSFufDLYROBvk
IFvXavYKCNwLO7UiD7G6dRvimVlYkcvjn3rEOtmTiYbD641G8p1cVROuas1rSp0S
3YLuercqRiBn+IGQV8Fdnt7wZzTdr2HGBrohNkZul/C0irU7FwjuavQDIrWafOuw
S0h3I7TTLERWbznv+CMl3aiT7WD8sdxsshDMi13PbnUTevyx/q7RYJM53adZhbQU
6AH6QaPw8ZLsPCzdhGd1ZIOCMUupLngFBA3Iqc6fxiNPPpzQetFKaLP79Xmovi5h
zb+xW1XIlsZIzy9Jts0oofH/iiQRw5YUw/rKtBsRDJcH/FZrxfk5OkRplk6wgAng
vsy42miGExtGLjt6jM32NfX0y2UdCsYdj/A9n3/BQXri6i+ZJSs3wYuvJE+IB2Bq
cvtrCPaM2/fYPdTW1LhEwy0Xhemd5aEN+lh49LP6zEntvyLuCAwCjkRfNVYsm1gp
nZqd1FnqWFaBBL79qvVOdzedBLzkIFDhh0ggFzVOUrIybeGQW8Zt+H9zia6S++5v
tGUOq/SDQ1yLXrSTX5x5BiFkPP8YNfqbWYv7T2Lu9tSwIgOOJQJ99+d/7BH+Tj70
V4Tv0bWdafB8lnADvTA51oNKuYV/7RJVR9QVKoLNdLg+dG4QjcDaXC7vGAGromLj
Jnh3umz+e0aHmnwiBxAN/anzroajtCimdCG05xf7ZG9F6y1GSasBsiqOoW0/3jd6
3G903rLU98H8xqCe8qrvjUltQJrknrLRc5626qJh09+NDVbTMZEJtjehnu8ha4FN
pwKwMKz6BoHrNQ/MMi54pOzGfD0vjGqyfYB7BmWNFyCinJUeQX6hpsnH7163CDrS
9T/Ak3qxinh7YotWINTlxhM8DPKOFhsgWez3LbcYHL0YFwZiiPhpy0G5ygXBrna1
cb8FmEqYBq3AuqbRnyjtX2+GkXBtL+2KEpGex9qdj8AqDg2yUWp5bUr7lG2HeO/O
rXGJag5RwQ3oWa6PJ/YPfnRtCeFYFxizSxHbhm/WpOD2bvkOG15UMtOdMOmsPmWc
mKbtjBoFKpc7DdbWyuTHhqZGgB9hS5UxmPpcfwt5ew8RnZrzej7TBYL+3wO9w0pu
9tA41ykMLJLqxPrVQuN1cd8ULSlY/Zrn5RwZbX1pDA5DVsMgjKiJV7PaX85K6N6a
lExZd4ZFEnsZ0u6fFhke0MvkFZdkaVlfWdQRaqO679R6RUdO/UDrmjUfn2BCt53t
Kw/o6z9GDXwANxaOTZw9sTwkK/Y4SPYRtguBvRIh9GBCvuG6xuyz2s59+Vr8bsjy
zoguf2pYnZkuIYRCDjg+5nB8F6gaMpU70CR5pyIs+bLDlmzqL2N7JvcYkEnnlGsv
QNvZndvFO39s3FoqSA6IDSoG/rCLjy8fVm3WmIPC98BqdNnoiX7f1XPM+nTGk9Mg
g7qZ7ttDVIs1NZ92cld0yr7HR8EIswDF2WVE/cM0PSx2w/2GRNGdz45CEScQ5cKK
7fDUFj+/xdxMXJLB1V4wYVkUD++cyjIwDiC1LEoJznoL6ksDQrzgY5hskPE8ohZS
rZcuSPm2pr6/BkAhSB5HptePl3VUmEfPgyiL53/XIfFwdAShOahzzvGEJt8JKI7r
SbNjgpQoW0EWfuOp5KrDm985RVzLuDFA2EnCYWhixChLKR2U1euMv+n/Xu3ssbBW
m9gNSn91xdUNnp6dZ+52K1e2RP5M919yVutuTPOeNFt9I9BD6VWLMv1+1vc5HY1J
O99rE/O5O/bBg9k4OBgcqNC1ynCdTiM3POIABxGRrMjU7Ykb96Pgied0L/5L+m2Z
MILLfVD5g6ehFdd0BP5f7oTO6dpzxKtoR7Nj8WxlZ7fe7KFvV40e5HJFR6hzXpgx
S9xv3YlJJia119KVKdP5/cswQV0P/WED/83LyEoipEJRM2PkewVZ393scQzfyfO3
7rog6zAGzNMH8IEJNNhdFY5+eGOXGkFRFpeD8hFwtD+kdmgZyZDISPIL7Y1Xq3Xt
jdWHMq9XHhgkAPspUDXvVnZV3M4Wrbgy7DT74VS0VUhpMZi6JdmO+6gfxvpFhczp
pt1twFGHTaRLDnr+WfCnePWk5IvKlFZYGEX9J5KLKmKlsIlo1uzdxz1uhu2DvwF9
9YTgUPTvpXMBeTyxDoUOpp+sSMFvoSYG7mp4lZ0v1jlSmgjSM29X3RD32IulxoOH
8Etn8hDUaNZuP/px/5Z7JfCgoi28mEzf4uO+8KfqeXE3InwOVGKt/arzgEebz3sX
JeC8rN0R1ZlKLoRecmCMzwJuFxgONjETIifo7H0nIPyuXoBEFr98OGvWKAba9nCJ
6N6pViCsPJXRExuBUABCyxAgqQ43oUqJECReJQgwzt1rQ+hL4p4zcNeGlQUVZAFQ
kjW5YBgAIFqkt6Wo706gww5Pz9DHgX9ZaA97CrnMq0hvICPYw06wfQmADKN5D4FI
0wOH4ZgqHiHt9cB+wmwnMTzRExfGwRYdwxm1e5d/r1eLWdUwZ3T+KHzWruET9oxL
9J5hzyW7niUZb0Szbu8uNojEHN1yqfbfADn2VhXTORJESS48sDN6jIGWRuPJpFcX
c/pXDzSiG2S/M6BP60+c+dErYvrj0M7qeA3+f2tu5qqUSxlVgXOFr4IuFBQwYL/k
ULJX1SErqRAU/v56aJIVpxbRjJ+fxx44q8cHz5WsuJEvg72xQ7HTsr595camKMfd
Xk4JbH1zhjwvkSshuP+smpVenFKKJ24XzffgxagygDyjqsVaFewv48KdL2h+iayd
tUMSMeqM8JuCgPcxBHn4gnZoNnVx2FDY7fkf701mcTQJ0gOsRZWvUV+1t5T66n9g
selYu6TK1Y52pM7JQqwEmRvx/NG+DOe6mZnFkZCuANYe8r6q3P/in2maqS+PDSjG
oJx5jjDf3j8R1Dwb7PngTu6kFchyVS2zuLoDgW7aYD3YFisjrylKQv01kpnFX8p+
kHpMwzTsbLq6Lz+jjgLo45PfT7r7mmSGZwp9JXlpMU8SqJxlWZUdVMetl4FHpLkx
DapTkOEotZsCUY4rYb9a7yOjro/eIgQz/ZkR5wHlmamHoMbrntrnhGkEwt0Y1F+Y
tL7+f0N7fu8jFqahhJ8JDljFb3OZVp0fldp0T1R6/FjZ0rdGjoaZI3ES/7Fy7DRd
ipHifHH+PhzB5ZXZTH4Ufdo4igs4VWlzuogn/7PNS8G8hI3lx+AOmKEo0eAlfmp/
r0PoTOLaemet2w54eYlilG8nZxddZbAUYeYTd+yihBV2IAvv47NLQ427vGnIYKPh
dSQpAKWW9de2i5E/dEco5o3la5r9Wd/VBE1TUFEJCSSYY2bJ0T57lt5ZBC3t3Nhe
NfoggS2L/z9h6lMWTYzV9rK3vdk3I4G2wlxFyU8wUK0/FIJH13fyn2zBKIyKwEe0
bJAOFAqO/cP6Df5o5ggOwvHOKlqbb1DRcSKOVCOLBSZLfa+8uZPXoRs9fe+O+fHG
ArVMuhcEwfn32iC/jk4Oo8gYdy5dt/qhmKyl6hcGAobVgyClf91FQ1GFUgbMsWQ3
OuCb5zFly6D19m+AmAARGkPs5GY/GGN/gKWlS6hNo8mAZ22EsqalK43L7FJaGEwT
vJ5O81g7iEe5YyEhKYJ3eJrv9OByJymat1UvjKrxiGgn9tefoFK/QZNFLTMCGoKk
yJ5JSTcH9Q2D4R5wF0VOYls05KDW6w2YuuAShObjKJOm148baRfjylHb5W23HSv+
aompZFCJLZnQJmBu6vz2ocYRK4Z6dqWf3JCoIGE9Y7VAiTzKNyzxnKb46/Sbx097
Q9Fz3EyEvoBE0mfEFBvw7KV5tuaNmt5/Tw3s4ceXF78JJ2Ko4tkKo+GpFHo+5tvE
H027m8Zgjc73Dov5J5al0LU2rWdb3l8BRVtm9oK4DYAGytRwQEEOhCDUaGieYzy/
AJEhIu87BrGEp5C5bVXNxFjc1dkKdb2ZlRJ2IdWBK1LnqwfF+4NfDuDHAjAlObPi
dMUUSOjbr8fyGfyERGrzn++ankyzBg1nGhoSEWR+LC71tUGqqLjjOWqd7iqeeDWb
1dCZuvDxOXIH5abBPs+I5yjJsZyu/uqokJgjMaVTi/mC/+xUSvsZZ08myFdP9c6U
v6lfiQ22xq3VIyXpE7iQL9H/SMSTLuxGihRCoxcBPDBtuOxTj7M83w692G+HUMZY
gL3YLr/z45bQFysSSu0gFekxc8ORqvtLGzdskPmADDFxToTbpxvyerT+T0pDaMJP
Wx11NobZCWNB8Ou3fo8oRDg9auCrOVAqHIa9aECfUM2Vz4rTua5mpaDb8pHQ9k2O
dq35s3UxmX8SuZpdNaekvEBbBVsSJz6wWksZJZ9XSSZjL0fv1HNsR0onCWkjOnLr
mAK8JpM6POs5gRbrNuc0kO1bLhPvQrqDmdoc2PYLBPEmworXpPDyT2fhvNKsaghH
imaeVEXSmnCSraVYlbvx9jY3HWDtbQmYlRJu+HF1rrLCFeTzbU6Gifj746Pn2Ltf
UvMnaU1uGcGsv52sCbfetaVCic43OqoHBNa7ldegcnWeD/njtqtpUysNum91sW4x
0X4kl8RuTs2mWguu9UUo0zb4p4H7nUzcf+XLPZdRNDK3ow4fwiBCAnTPs36X4SxS
ayyb4TqLbKp66T87DncfKHq5CVG0zz5hP9g90UW0/Jwhg9ERCxUrrd9I39++Q8V/
IXmlnH5NuE6eesi+ziGDM6WdoJ0AaSXNxKDkCGklDMsGsUrtNpsWs32hZ/vzTTrR
Nl++Y63oxsDxmWiZpaedGouVj1tHV8eID7y4Cb7sTzT3bkgOWTqV75G/zCcLzN2j
mS5q3j6JI2MI7RPEVF+97a/Hv84pg9ITMTszo8jf91zaDpXp+3l8pAaJA6TEBjXb
dCRaTgN2TK+rdW6ZTRF3/a6Mu+0IwJCgSUDKvzP5glXXQsHdyKiyIya3nk2yKam3
qSlNSQzXGJXKzJbylokEQiUkFfzSEdklotjwc4yvHgFe7c0vwUk2axQ+DCVgmAve
1Vx+HcBKmLVb8g7JG1UBwOei1LYARr4wVIKGPBCElkjJCNO6munOoXEhZfeLHaSI
OKiUCjn/NzQ2DnvbxQfaWoMjY20EVae7g9wl6tfxqbV8WW3lEFA8ixnN3w7ngpP3
GCjMtw0sifAjCwmpoYo+LN7dBbaGhzAt7vHFqK16AkQFyHHzMoKj4xqRa9R6tzDs
DlkijGHHATLsk3peNQ/BJHAP/nkbKZ0gtx7lzddmoAJQDQLk4I7Fl1ZjiasrGyGl
kLPjKACn3hQYd7WQdoKIwGaV5wsAlQe2EaCn4O9ceYhKoXwUOnunHBpalBo1FHvb
JOmkpElhbuBFItGUGgV6aH4DFUwtquzhjAi922Ixffc8SUQ7fV4/0JT5s2sg+WcI
/Z11BjqpdfuG9G9Kt1rmr/UXyB2EpCd6yQVkeWZKpvFQgSJephOlH6kCAd+gbxsR
ZerPFCsvUIn/F9n52/VJZ0fTE/jRDdDH30wIabSGc4vnsZURWCYeXKgKET80Iprz
yTVOqoE1Ua9ukvMGrC6Dd0hHWS0Ao2fm8EHoOeMmjkVpo86BQ8DxaJJObICz8kVc
qkxlWbAFPSlQZPHbAUCrLM9Nhl2iilKsQLx/RyWFkSq30jkUwx0Ay2Ad2FAyFCN6
FXsc/jwcMaytBf4LLNaru3GGzxVoQ4EpFnvxrsgspJVrx7BMLtCKDS5x2Lnk08Gd
hHmgmrAgpNDaF71npZAyAbzlB8rN5kC7JtusxIipsQxFo3n4cBR1WsyyhYHUsFmw
4JKg4BnIABlydebPtJ9BYOUhiRGqVcbhOsTP3MT/YKVCha0tzNjguXtv2XyrmHH7
7gh5Biwd2eyClH50iytov8Rl+6KG3MMo8qv9bBgFiSiVcR6WH7L2O81nVBsFxiUW
SnlLt2sO6zDg+3ORpO2GKLdVOPseaXE+AY39YXzo6PP/sbWFDzJd8xAZIHV1E2Jt
VyaOmMCsrJLXdcUhMGGzXI+6l+wItOHX3FwkcxTxYoO1IYvt1FzUi/FzekFJZw/q
o0Pl8S3Jg84bkfKUkuRVlOZruPkQ58Cy8LhT8UznH747I6/EoSuIx2coQxIIhwej
PNBMkAJKVNXO2nP/5pXY8G9pja54AYsR5e/6MThTahjI/rhJX5hh9b65t5ZgaE4M
9IUGkKtyW0ASB99fhNCyWnERWAmJSHtMO+FF4ZjmTladVFbkvkAal3FJiGeqc2HI
mZ8nIJmlmka0O30KKXyhZ/GLyc+3QWhI0Rcfk+cpC/ADH4/Zm+RgVoejSAyKtOYs
O8wJxu4IlaWxcsQSjY+NzG518TtDBQKh0dgebXdSkgHWnBpXqq6uSqEsSalEpTUJ
SNfP59meUzhvNglqkmRypNnhCMwfzlXZSJJNju9H9paPffZByQn5j9o0+64F3KLJ
bWyV92/5qSjnDY0xz2w2WsFcwonbBLciVP7KIXViOIY4xsLl5hxAU+6PR/gwrOLr
RDGqimVqbH+7keM9Vw40u0XFQ3MAPTFdL+gOtU0KBUD0lL+GC+JzbHqTr4+v8tKD
SNGEnYzJL+7jiMPtFZMESBqUtdAFAISLCDPvV966jJqll6fg58FH55PJ3lvERV0Z
rsNmRER79Xpgwr7aMoD4S3c1gCSTHc1Ovw/8zgsouA7rbUNOKcWGR/uH+Psram4S
Dzrs6m1IxT8FCDjrVRpAQO1KV5LHZWEGCEx0+iFEurOvfA/MuNLLYsHAmAQIMv16
vpCR6vwI9FDHMcgdiUcllUus1KOPMlRwx1L/upA0pjut/x+ihmqUeN/F4FZoVT3p
EneUQ8bSGlJzobpzYteZ+jq/4r7GXivPaqp1jqcAABTivf0ZgCBECbfPQuAzd2di
gQphHu/n8ivYylo5oJ6mKkH3rUS1s0d9L3re5Wmgna9rzHgexUnWCxnNOEu8LCOL
7Im7k+MHDs0eQzkylQEl1VyRUJLgsJszoNaKvVBJz8+/bO/qp3haLb0f4FRhF0AJ
5juJkGwgl6vi86d1Vry4Yn/sMhwV0CXkLngDOC6Yjp2CoImIL6+K/7AX9CdDL7eQ
Qluvtwvrc1uqpi/rR6bBlezQvqTa31c47jZ8r7Wa8pYWkGI5FWlWDDKj3MVsy6cy
4w40UC41MK0AWPM5rY+CRFvTsBCPvTfJ5KeM8Keq+9SB4VdydA4O/aXEzYN9IIsP
2ib4WANO09CQwTfEiwnsIIq6r8/K41bLXtit5yLfyGh7UCWsag0Wod4Uns6la2OE
w39+PwikxXzMOe0jTro/EVstqPHTIGYfjth5SSs8jdBYP9wnW3uoYNlQTIiSQJ+a
uJxI/JZLs26PbIGWt0Kl00JKFwLRdafdw9u5ih+C2xeY74E8bvLWowOtLuEFb0BV
cO55p+JGUOs7B1IKH9c8Jft0XZ2Uit4CJ+RMSg9EhqGiPCU9h9Ag/+u7Jnrut5iv
rVbH4zpOeGmGjxY8Af58hUspy9v/4OQRosH1WSjeHWi5n2dt3YykEL3T8FT6OroN
xeS+/gHaBqwPYqJ40Sk8ofoaIdR/KF3S7Q+NSQXVueDjwgfzq0FS4mhTkm97qh2x
uDMFF7xm6mHc/deGj3eMjTYMilqHNj5myBEBiGhtrVPsbq0wjJi0maSoufwAFJiW
tEFuBJr1obrKt2oh/LNdZKRjqHrJwRK+OncIVJsNWmwh6iXzr0lJPdUOSNPcYvWH
GEyOqzMlibGcxS0FNCcbZ44tmJ3IDfs0v3J0UBiS6etn0s0eWhwlC9GNKWULYUGW
ZleYhhYYF9sH6B1m7sHDGbmuSw8RtACc34hd8QjEFCYB5glpl0xdc0SHsGKwNUj/
bUlBpP7X2aOXTSeOavj6BMFpbbb+DkqQYAhrV0Bf+2e+rCZZDfa5A7OedqTIcZig
kC4Ns2Rd3GANWdIZq8zcN9wyFsT/VmwlB66NJW3csqF/wZOThJ4lD3fJ/0u5KEV1
QHzLFJWsABK5dB7dyBbPsqVjHSOcCojF/H60iMd7ubwG9BYBXaPmDp+5YETrJ5Ue
SEEgfPTIBI/4ZbyVsIfg/XoqPJ63AQ1gdO8CkB/KsV5gtIDK8uUdSJUSs3g8GhTQ
smaABTd0fWu/6tRUT+7wEmKDR2qU0KkI0w/F7rZKoTQ1ia4C0wBaOehfB4yO7qKO
C5wshhikHBqGBHeuyIptd8DCH3PmvWAeexLJRU/IPPuhtJ4UCBBjXeomD3lGC2Bp
iXmHXktoy+1joZap+nOEGR5OHS32oOV4ChE7jJNnqOU5PhyXTVlD19BDDsPSoyLw
cwk78bferuxAy21n7eB4vkSCWms8HYSzLrT80ALVIn8kSSTMe59VJeDR6V3g504P
YEtbdcDi73llnIVK3lWaGihr+pPG+FFOR3BnP+1iEb2FCN7TEJPO+Px5PR7uaMzc
JQLmEiBIAuWSxe4nw5X0gpzlzOFd8Ql1jpgCQhWrf41WS9jDUvDy74HHXZkr7xyd
kaHQ+myDP3c73/tWh6AGDZS7chiDdwIOy+14MV1k6SZ23DLkcyLEbmInRNUtd0MY
0D5k/faCpEVWlWQFX6I3c4mylkhfdUt66ZEIawFuq1G0BWUODLp1E+lqv560BVvT
CJwFMmMtdyLzX6pbS1z2WGcC1eCdZX0TYoO/+YOxTfgjaoZmnxdI7eZ3w94zSc2j
PlWH8LV/DqS5MfSJaENVjWij2HPS8tt40LLir9sTeYJUTGiMK5vRwdSrvXSg3qye
7ZggbRmUdzziC8FRRb2xUfoRd3ooipb/WrPmY/jNYMM5ZMbYcbKLJzM5jUpAe7sB
hFF4Kc9s51W5Xq/LS9Fl3Z5XdhhMAMd26L9ufU4KvMc9MKZQOw1V62mBUjx9cI8W
3mIYZoPIyThPv1l7/KQtx0jOXdobYn1E0XKOyrblwW05IhW+3biDRuq77ZvwIdz8
47sUhlmCF/MB8L0Lv9UIqOcmcUaWNibTLnhZAPtBKiWIpHijKBAT5lzvOVMN/Q+U
IJV//XFjmg8gTklr7/NF7cTt/yNSW6yL10AAnFIKW1F5KrZYKtA0qs7rGycGXqq4
xUDgQOaunEEiW01xMeKOcf++BL3NOKvX6K1It8uYI0YCi5cGwM53INU8PJKB6q6O
AP6BNUzi8Dtwyrh6Td8D0Lfqh4vuRg2Xnsb4eaW9UEn2mkQdOtnfisG5nbutgjCm
mGx/GGPadPB911ryYVSgTEzPyrS0AnawRsJ5bqUIuPW/HsQd3efd1+joXKjHd8YB
TqYbq/bPG8Iix4WgHD0dQJxpab1E7YDOShmV3vXFIr5JnTEGkRtpSugjytcwI9Ri
PEiL0Pq2Miwm+uBGoPblFb8zaCNh00yFxY4MTcrugpfhOvlWZJ+xaGt3ZTYFGIYb
2GkcRTne1VaocFncgwuqi4b+jCTp+X7Tlhm9VV5d42fo/tKt/TEcrm07Q+GDZX1F
EZKXI5kW/W+OACRVdwDpJud5PspprYqSb5/8sQ+UPJJcFdfsqYarlLGujGWspfUm
EnxURr9/5Y5otvgxCoxfM0SfvYJoXsGcHFrYhaW6s06B8wrvLkVDbTZY4J/OnmlF
6/JkGEXMSXnOcm3apNb7lAa1aybNt6T5P2PzrL6Al6cn3cIHZbDymz25kdG0G6J1
u1/fzMAe9wBoJ7acEQe1N6wUh8T06Vu/KdXabCaIK/vz9/x+ne8wWsV6lZx+IDxf
jQgQNjzRwNoW/9cDXwNiQoWu80lanIVeWswcC4FswCCwvCE9w1kxvDKEXt6OhYc2
TXZsA311Y1cn8+nwvwG4lSiCD9TWe3+LRjEnvD+D/eofPq/5CxSifAtiDexP0PPk
P037v0li+g/0jALhH7vFWGp0Dw/yLLBS9+HR8WKfXTbebhQ3jIaZ6mzYsqq+5Kj3
V1+iWu+ipNc3dE9itJ6Yj+TLRmsW2GrvO1K4YNCDSRdPFqpjQ0wbKnTMmjzVxNyS
zWk8iMQjEVRCC5uWzP1GWmIE7IBiaG8mqPHIuTOwdCDoD1rybbqCrvKbIK6JOq0L
pKfpA4v4O5r3hOW8oAhFRSVHrPIJOqjbJ0TgnTOkM50AXasMH4JfasoiTb8pbYAt
7y3yvXcyQyWPYg7jZKUtbgKsO13ZWwc5TLoCq7sdK/yr8/eyQICx3pnn7JTNc4QK
XLj5y4efy+Fibbk6+rOiQfXd1zhs8Fsz5grIn646oxYOlOJF31boA86uxQ1eCdjD
1uUYljpjTZvL/3uatDVs70Bm/fdK8sVtpv8nwaCM9im7wDyjxEMYx6Vg8QRgY+nf
ppg7ZnAtHfVkf89QaRmJqpBlM5y2u2CVBHjCgh8AmgX79MoTMhqb43KzY25mj4/L
QqP+S+Og2v38bC1e9WnsafuJXbJBz/pb1bnIqBEEMwLV8Rs9TXLlSB030dDniONH
9i2Kc3A2g588L6Z7EJg00iq3aizRAC7+08IrW2nEIxpB1bFfQhkipJOQl1omRJ9R
/Jezbv2e6TEhOcrAOnvBdFGB68DPq/rS/531uJUh08inIai/+Kj57mj1ytCW3GIE
4kxp2dN+p/pcGhx7qDKQvsQ/UJzMthopiArwrDrCtWtJxeqRJDWCIpMcIYRVCoTi
XDF8I+ykEf6XTHZiayTumReGWcpf4eNrQXjozQd6rY4WinsAfwPiP+BB+KOSfSS7
5C4VYeU6SnGZen58UB8nO0AMRAxNdiIFx04a2gHladMnce18QH54W7aH03+yNPkO
5xYPfgO71REK/mT3rfzi3UjF4X5VuM6xaGYv5qyuWCmwKlKj7REQfx8C7nS4+Xjv
9SDfVPyOiBpob4yRUi0P29lEPRgDTpYBTUXN0mhT0xY5m/ifTvS03BckgoCalUKB
dcftuDjG3yBcBG1z4XOq2koXP91cs+O48i5HejfJwQaP/z1ADk6NXaNLJjekF9N5
ztWCAIKc7H039JbOsaHugiFi9poq/Rlt1sg1tPsPx5FbdyAU8VHaJuhNKaCJ/0WW
P9n4WOk/rAWfErax66xzIkPA6/w/on5UDu4BRkg6IZb/lL2fiTK9lAq32s2GQfWa
WStk4KfoJY0MrKAEcFhBxTCkNuxOTA7Zh3MT0K9qUtFeFNUKhC203YBs+dfw1f3Y
HitYqAaZ/Ax++SFpo6eAh6y7E9TV0T82EqwOhIKcJmEUkRB5+r03+OQF2bLIR7kK
MI8yQz9q9PwQswZENDGidFCq+McluOmo8ovac89tqNfnfsrWK2Rd75RcxeSA67pq
1Z8AjKvp6065n5Sxk4Xok1xp/A3VTi2FMkKU29Zrb/6KOO0Xjxm0LSO2R9MVKD4z
Vitl0uJfVgsEez6XgrpxISyC+KaV89JqlhjkosQYrgjrE+IDHzzBoFVuGFKr/Ehr
LgRSs9QV4PHVBPkpz6+zVEP7XdjiEAbMuI0o3t5D6KGBSORD7RI37wWu7yLvI6rZ
QY5v9EFgGoEmKKmBvwWofswCmxbC89UyxKsvr4naSLY0Bkf+EOO9MkKowFfQveGc
45h2zeWv8ENE2M5GXbq4BwxukCEDQUQ0e9rkERIEA29w7jOPwuK3E1oZBFvnpEnU
O8h8DWnhpePrCxbY9IM4E0Q2jhab4tpHyXOpCSb8dfizSyVbZfHF2upoeK75s8qy
PhsodBbjsNi42kjEvfpKRopG1/5e1uDnF/QhZSGC3vFs5UoKK3x46EvAa/nVnnqY
FDH2luJLq0uqZGYTGr1EoJWqloNCdiTIW2qViOxx0kAaIdU8ni6oSbvDje8W6SK7
ciIzTDOqwxuAWZ+uChLSFC448JZPHQQCeoHsJ1gO/LfjI6cuLlqt2olD5ns0SqWW
Unbm0UTKtRj/G2gZwuV9trIsSMsf8zwHu9AaKGck7mJvqotiFZc6VbeRFRQc30TL
v/X/q/dINymgPITF6z1eQ3xFEzESMJHMgVOpVkFBja8T1bznfLLltvTPPusvrjkz
WqJ7eLVX7U75fJhACDp8ETTfLKtjgyXrEVTx3LTDiG2bd/HOhjBDefLcxnR6uhBY
Z1sRnktqDIruPp3kTlpZM0cj6trsuqF4qPnfH+yqtcBjBi34+nD39Uek65+gQzRM
8wdFxTFe5uOBB1Wf9VZYez7v5L2qpKtMu6P9pZjvQB/18ECr4sMi9UUMpoh7c4hA
dA/e92squ10plMKJXpREowuNq3Q09m3l5chI84JVd+DVChe+ixAqkowEfGreDfjG
/DdC9dkIRi9xL5HsSxjcvHjVu/W2sbhb6GYXz+/dOBPUY3Br0LKXELhA2+MkFnJn
3Yovc9lj2dwG3j+fCU0wfTHN36FtPrQ2MpOYE2CWpQHmw1ua++h+du/vJRPgegPw
BnZgkUkxNMJ9SQfDXXd5BoUcD0QnMuUVLoD8tat3esQkWccZyTK/10RPH04F7IVf
EAPka44Lnaa80RjIqesnppgzEzZERgJ6k0pTPCsakry3X08BTIhRuyVfDyWyBia+
241TMjx2DQ89JMcryliHY5xkeyiW9K/TXy/W7wkOJiLCtfNIIz9w9hIkvtJW58Js
hZG7tzENFG00ne0TJ74hY6+1UHyQBio15r657oRxnUoFuudZMNucwiVtsnOtUDLh
pm/ocpcaU3F/kKl5efmmKengu5Hal8B4lcJkWNXkZ9RK9SUv0g5mkx5xvfF0vzNF
z71DUNH1v4I8hedrEeWtNtVhpISQPrJ1EmYJgRyiCCTNAl8qEGq8xVGAG+lk2EBn
YldcFLX007fgGCnkao/cFoi9uqBrplbsLOUfdVLsevOuTz36eWC7BMnCmPmdxaO6
Eow1HV3rtGMAQDVarF2B6D18Vq1/vV8LSF/cY0gqKFWVfovFA6Zppmu4xMZmiTL1
yRhjpyX3aP7Vw/i0X4KIi/OGMzIp9nWD+1JAXWeJQAxfAstB/ocai1bg2SFLczaf
jgGZlwWBcDKQaWYZhN4Lq3RGldHIa4bZVuX+LbJS1YgTCmCrz47KA/UrGnhiY6I7
LN2RBFI68bXCtPB17xXvKHkKawAWClsqvqMmOL3KW3gr2RP/7adb1lDf+MnQFRe6
fdaST29e3ZlBgxWKnYeCH4bwy3WmWYb9n/EwHaWxeGt/KmXAeXIQ7lwa4sfvFBQZ
+Z4JJOtMSUcQrxBz3xh+2bbH8Uy0Ps0u104O+UKD14RzWW23og9Ohnk1c4zJbWvU
R2u6qSYDH15c1f/kqCZGdqn03yMCebH5VUyAEN1XuHH874zSZJszlNZbslPboWma
NoPaoa1cCgWILd2daefF0dIxkMJ5cQlB4n6HDEt+Ttv8V1+pWJ9O927lBuYdJjrb
ULgePMbStZ5xcSnBBo6QY5K26xk1jOa5YaOZrcnefHyJtFbB74+jggJrGzzDsiKa
AwPj4piqk81BuQ9/FX3Gn/ZsBzJr9D0YNcKZxQ19JitdpQfanW6S+IMjIPAG3rsP
VkyAmpajFVINhZFnCGbIHwL6gVvs//ZxqJbReO13Cqjlgo3sE7k+QZ8ma8l89XGA
ZdG0MRDecp8//0nox2gEc0p/4WEHWLepLkneq/5JFR5QwEOEasiqKTJpPYzIupD3
xnfWomycoCqZpNf6CCudsuvPf2RQvsgdROWhas/OdW4vz6akpxGdZqf4dojUtC55
M9FQqPVDcF10OzAYF/V5DBbP7TLChwR5CtlE/2U+x+Py8oAHqiLmUMQlBrbS8umR
SAEr24FBNVd+XsM0PgoZfpNwisFLcKBsffWD0krWu4rLvs7v33hsPMwcusPj7lej
Mxt6I7Qfi8gIoHp7R9xYReF3dfDK5rUpG+a7DbEA+Py2/wIvEP1hHWHwp1H3yM6A
X2YLXKHczIO5AVa6gFXy94qa7tLtcfVIb+nAzHEfP38Q6pgHm6PapunJmLDevKpY
rxDVJTWH/R7+Y27gvKLT2PPyuQDGKN+/rqvaRxpwFjbNsEDD0K1zqBo9eiFw8eY1
1PEO8NrFUFFFqIUWVg+84ZZHvMLgEyqYUeDQhO+UVHy3VSjgx/OGg+4KoHodaAsC
aMHhfs+6IpO8Me5qVdyvYnk7HEaAUsf2QgAHY0X/Et/F1HemJ9oLJ/dOasTvBibA
NjHKOcN0IX2fkc1sA32zCUyD+eY0ta+REFc9qt15MMny7lOzLH4jgMxrng8mOHwf
pKXrzO+IOpOgT39IDaxHiZwWnn5H6r/DWvX//oisAUcRYfHPdEyZzeMHXucgfI+h
zL2VYrffp0pRjteGMIDTWqILLyb3uB/uEmRY1Ok/bDthFxi1a37zcmA3ACaJ+4Bm
uYB8OQ8Kphw52bN9atSzdv7pG6/gLedWp1BEyzGk8/WOkTTdrUmJ9Xhvs4Qah1Ap
OlgioqZNMKKINMfa2m8WOnKOhnhvGiOmcKBOIyZbS/rwDyvOL1YZ82AMiFeVtMbG
hArMpyxZmwrsmVqzugXAP94n2lef1atUZUWlGpNBIbWNqSCVpnFBXYJrm3vP4vVE
ZCJaW9f/NunBHrEiwruEv+cg6wtbcVSkci+3oRJntIBw8JDmLpUo5zyRPoQs9uuF
iyXo50+X+r4W81z83TAnrzkm14ueu6E4uCXZ4+tCA5ub/r2Eo4WExdY5d62VFm63
xGyOJtQcVjOgDVTZhbbtViwyhOdi9ufDPPUn+grkRAkDF+3Qtl7CuKVbmHRkggej
brWuV2NyybCoAqJ6hiYIcOsnaG7jYPCYwhPCmy7+NiW3R9ClWV34WO3d0TNoIJSx
OkrrvApG49q7b2nyfJj9cmEXM4QlSnBA5bgINijAI8HPTlOP7cpOxTEYbYADJR61
ImQsE25PigOD0dCmskQYV3OqUAI8fUXWewezZ1TL0fEkydQVlkkGXpIZuhucL3cg
pnCyz9xCN5Pnnwb0jvPzzoqLZ0TiGgNhNAkJTu+SFJoetg28QNvcAkgkFdNYktb1
S0lQlnoPlK02ljQohRdTypsG3+/LMd5TO3xG/UxaTZs12TyYjQkReC5E2C5fyJZF
Ke8+ApjktcTvJJXl5x5UXCy8H1pbihdzA6Qxd3tRP37pMaViCW7ktiTC7MryWdMa
MnktpnnvT6CaR6ZhGv9t63iaN+EXDbTYDB+K1vmWOSFAy6YUEfHpkoepYuGnkYF8
rbLMk9vljGHJh1/UfG8NnOcRTmJ640x+fmesKI+BoK3kisVtbGpMJxjYnMas1e71
FUXtOvZyvQhqhhH7uLeT0een0BBYfNo/gPjt0LRywfyisJGCZF3hNA7oXyEx1aVc
ILsOPGvN84RdDmReHDRk1DlSS3TuRTK+yQwZgAZLmVAADVCIZKydEVWl9Q6NsCDJ
fd4DmpWwNQuWUcDXgBS/LCt7XXke8gBgmlxPPZmJcwrWUQiSspeBhNqVLKsloTM0
SVXSj/LSyen+xo8YaQU/61ehYkukoWqgL5lyZp6fX00LFKFGNtNxIX/hCEiICdDl
+hel4HV6lVg04CVvZHQqwFqxM+KYFNusPKh+U35j0Rc0eM494HbvJYEL/YHIQClQ
4EM697I18e1VGBHRHy7bITnDD1KGXxaeSj1wO//vz3vhCMCDSAeRwg2Dpo5941xB
GTMLE4gvh6+ZBT0ULURTah8XnZM4HLjRZQHem0dnFpdLnLU42WVhfmasmhjXs8Wb
TNBx4lWHAC/7GMGwCkiqNjBtRH5bsshoPaXjKFKiZlNpGENPoUq6nCOcKKQUklU2
saPryqBDDLop2ERG99miHfJii2vACT6+NIKWGLgU9GovmZjNUSjW/O9R399rXilq
7X8UxVXkelH12skYFv5naH8fenLuTjDinAInzVG6AErSnmuhWmgLMCYhQPXQ8Riy
DBMCT4iFr1pXFQZSgh2ZmNRxTRfAVaQvn56uWxgquogOb92eAYxdIfma4367URx4
ZFl87NG3jyIk3a4J5zMUkvFqaGBTM5aJbZYYk1am2QsrZjggoWsCoNuAO2uZlY2q
DWpxioTcaPyywGTzasQXnkmKZVCbistXOkZcRfTKGBXGdTY/hwSJoAfeOVnfQidg
YWYzWd1CcQ9h7FU2/NueFoh08HUzFyILROBj+o42EWgS0EcYsGAiQXusFevx/WCk
dilps0y/tWWBOal1vu+0RYNw/OK4CT3pvMg0JtY3Jx3NRrZ2XwOjST65EKNbPGdl
VTfWkFhI/WKbqqs7tsbtfIa0V36H+OwDwbvVyO8OOWmTdVQQRc9uIVHaeuorpGvm
/jsWS7Pu8R8hVMdPbzzlH0KQkSEZR+kCY/mVVvN0oNvIg9B+1jYgMtt9ObAOnyX5
vjtbyW9F+2dzUMuN1KnV2I02rH6+5FLjY39DIcBrJ99LbVbA7RLz+YAWm89uFLKM
6JvmoEM4Lxu7TMs6dILXm/RZkOXdDJa1nTkWs8dw3XMhDJ16sKDexQVK6Jw2uFtL
FDT9Fsj2XyJVpS4egypeY+Ufq11aC2LhsXCkQv8ISeCl3RIVnbVwmYpPYpkjTMqs
pWKENwL5l1OEEenzZwpS4uf0xhzMojmtZu3fMVpnfSWPcF18z9K9aiQTRFsTAkN0
Bn6nRkfUXIsOJPwOWQL4iuAl4ZOFdGKgJnF6sPt7rfYS1DuNR5Z63Pe2f5/k0w1+
wY9FDP2dCN9GPdk32njMyyaap+/fmD2xxtRKFB/1UyvJzuiOlfEY70GmxvvTLn+h
jO8ho2LMklh6H5LEEexeHzhLsZmwARS/OpJM1zxFE4n9Jrh9FeCC2Bv2JVggMkjD
7PcXFrG79xTP8zcySpmGXNkVRiCW602vOn/PBPl6NCdflssLlmij6NE+LIdvEhzY
zvTmFhVLdUEK8Om991xX0aW0764LUs/nGiZ22qsGpAN0zW1JiXK9I5S7Bwq/elwl
KFg5FnC0qogqyK6IMbnHtDjor6R65tMTbdRUFm21aq3AU6/gRafCt6eKK/ny8CJ4
X4g3FF9LcnAtP7rKYk66ljEs2A4SU2rYZ5kZ/zO/o78CDlRAkRYl+02++WMKj+lm
lzJazH4KXxWiQY22ze23Oxjw/bHP9oMDhpUxvTban6yVGevYyCLZbJVublk3Zzow
jgzToBMsfYEohJtKEAHkngzo2O7D7Lf/4B+iELT9g0CqNpWAs7EUJR7J9cYLx9OV
yyBpx1vjCWEe3BYLckgr4Kceq0bUlr/WXnxBvSslxHomAcJMjvUaVB0soGzjoTEs
GPRNXi/583rystdvAR7lfopO4ztnZD5GSzHEqFexp0imuhvSJDUlySCwsibYcBo0
qhyIRie3MjuhQipqLtDYTpbSNId8gJoaPPl7cLJq32c0onng5hZbUmbIW1LHdBd7
ZTrf+L5CvJv8fosse57wRcHl4xS8QcbN6p6bm+NySnVD8iIMGro5QTRdGypebXTd
Hie0FtJMa8QCaHD5q0mowWhQeJ1oDxyzbjWk53D1LR2mKxlhEglnyAR4akt6In/P
JmfQoETuMRoVkeD9Qj95ko4tbSGI9mrEZmMUnXSH3jaeiMFcP/7CF9NnHN/DKh8a
70keuVlH0UZ99RFnjhKMLuUpBTtkqrz2yePGnIf2lMc4zuOIQwbQEsbzeEOq/pHY
L06pfQGfyAB5PYnoskL851k1R85RXfsYuwy5kZwMCsyRYqvMB9lAAPNT1BYT3mYa
UvXBGWsZTjuY4MqTXFihVwj2FptiI75YGQsCJMSQ3N5CCjwg1Z6fUto8z9my+JuA
eScb+w59YI7umudHRUXIWueR+GhWM2ygI7vJ+N/u+7IIBp4z683Ik/sq205dtjwC
A0X63TMeOq+rXftWFi12zguoEcZcAXGgZ2Wdjh5hS1i/On3Nms3cKNwXNJ45zQbS
1BOKznj6gHJt8qPxKjPjxcyw8+ExsLeosuUsOUTkw5KxnbBzOwk0N24npGVemQNC
jLLwoAMjAUGgxmyrbjGGTXELbVqyfdmLuDN6OLskRkjrNbyyDbvmICeiwbsR5uGz
a1m0uXH2Z5rTpIxxlXAoKPmgjxMd3384ejR6w+eltYYaXJcq8kN1VqPm3xh9wWjn
dTtZ5sz9bJdwLvAe78Rx1jm2ntcjc/pYlTn81HRHwfiBqJrkGV/Qjb39M0vOzdO/
5eYgzihXXMqx/jw1He8PrfeAdHqTT0VWZRrpNWhya0guhO1A3vrcsNlf0JmxKKGv
o6wHn6BIi1UN+MP9zB62y/jyw4PIKnZGc8Hslvg/7l8ivDqRjdPYxkJb+ru5BfnF
xpUngBooV0hnLp52+/pKGPqNkMR0JE7Eqi6TDyc2ZAiGlRWxtDvlVb9DXt6lUFHC
nFhElkeCMLnvmHbTQGxYrLjRRWJfhZAPeoLPP51MHqA85VuzMxDXuXWIF3VD+FTH
IqZSAB1IQ9e9rD5Ks9pbfsYcnbNEs+FrWo41WxbI9FrPGS3XvyI4NNZsCwFawGZ1
T9zFsaBTz0iFiUmXcHX/aXReGEhFvGZ8RiyQWHYwJILkL3xVlcDWMr8CEbhg0xIE
MtPh41lWXq6wWagWqZL4R4FTYCxGHxaQXL2F1VEUtFqofEOop8qIrAqWIeAujZpE
I3HjselSGw1Y9CLxcJka3D6KqtCufPRZfoCeOP+XGoF5iC7Hv5F4jWMHSnRA9EBu
ecSmt1ErMAXLEvzQQCTZuMLhdxeYUo9mljHJtV9smZKlQREgHHkHaI6IoncSi+4J
V+Bf5RPxR7fMa+o65RASq8iL7QMskSopdrGuzfOeUGiSYhZ/D6RZYwUOiy0f9sYd
NFuyneWcXwHHrIraQiPKehplEajvfghVgf1oVGCVIsO8pXU+xqn8MdP3FfLgopJZ
8dJBcL077Am/uGZZZRA4z/BYD7rIXsclORJ5FJwGLTTXzyKHFmbYrgYegl4i6IAh
4fB9sFFBYHlBJPSB7SNZFmFoSDLMv2/NCVU20JVBty2x7bcZbVVWAXJuCYNK1GlB
vSP/mUniP0jn/l/QCrSAITEABeQ+3Cbz3+6EGuZ4kIgMGdQ8VjQaeLRssN8JaAAN
ufU/64YHiQTuRo3DSCT9pXk7wre1jEYSo73ZZsfzywQhu6HvvReD95wJbdQIaMXX
vJhYtA7Qz3oHaStH9Xe4BVPRHBej4oM+LLEcwIOGeCF5+zvawsphYRtYNa7UeZoq
dDaHgNnnj9xRGQPPqhlodV2LUBmyojdMsjhuUrRtNxWHZsxWeDr+T0SKlj6lFK8j
Oqb6bUt1w5JBPv8qpwCdz/fkWGVwZ1WbfS1It+H8YSfOsSwYSpBYchItA9RKps2K
6Fuh7iZcBO7m7jePqCvV6l15eg3KJaTvxS7rx2Iy5CGnrP6fB/a2XC5U9cTXjFMM
ynuq7rN1OYiRpkg3MCfnCL9TTWb3yksPaUjPFfPzbKcTYEw1G2zZyx7pvS1+TW1r
1c6RXTvhOt23nnsn6cFf+XV2np/d92D/WG4HDBYth0gIuCTgtH6E/EMPx6qoreqL
iU3M2fn3/l/U4dug5aIBK6ZH9hb11qBT+IyVUs9YGKSYN/42ZQ4f3eG0GuY6j8s6
D1LA/xB5bR8AGR8e1GRFwlzrSQ8ZBagWCaOHfMJAhBY6lM/PkWdj9JjPRNAM0MAB
WB+Is2FNT6KDU4EK5aESFI1HV76kshmJWPWV/CEcECCoUnoWmW9bTqfvTdMpN0QG
ziqQdlDpPTeowmurSlFo+cTtfPDUg4LLSqaKd8fengfuMEjsB7nibosUhoPtHRaK
ac2LZdHqiFToHlN+n50kn/sQDgPqA9aOqA3ev+iKH5hpk/dtPFO14vgKmJaIhouM
FzlS9RVxatwZTaZo5T13qG6sgVH+GvQJ83UI5pcqSoLyGBcE4EuHo+OYo0lhTNaY
9LTGZ23yLc89IIrSzmZSOZUxxc4Yt8NTVUt2oti+WCV2IPDdjOKOqJOhXWiqxHSx
WDnj6is82mpDDJmLSzF6GKKdBqcq3uuWg7yr997v5OfZbq/5q4mZ4gVxYQ289pOc
Fbq08T9a/Elb3XrFvUv3WJPeynybsfc+12xckpsShZ18qx1cbzh4huPwRxVW5kgj
GJckr5hikBB4kouwybkum371fq3zp9Vlg3QraxtxUG1gvTzbCUwJ02G6dbYGh5Ck
7fb58Fo9fUgrCAey/9oA8wiB7Ib/b3y/5mrxvdYUF6F9xPQIRv9AwGBHlxIDnUkV
1SI3lJoH2Hf3NSMa57hn1Nmdk0vo3DKQwSNsUtBgJ5lODLk8Y65FzNBKLiBApUMq
s4xJ4JFdqXoAy66H/qteh4RgvZ29SOgusYplyAovhNyfsJ7jwJLtx5bIaFhtu4lZ
w+D+NHX+MGvvePDlA9VaVT1ddsgKoMjuzSqsEieW+irFqq6FXsMXeTvFngbervP9
caMErMNBZ/58C/PdfJ7WNrEpsWNQT9hIv/CeNh4wJdA/4BhU15larlUgDLGlYLNO
nOPOR8UbOAfXBtNC9LGpY802JQkFwMsTFeemszxIQSJuTsKN0ppDpBQ9dr829+bG
UkfaE+4wNuZ+RiHok8wkhyo5iUq9AFJ35XfhFkvUtOpWEm6Hmk3hAjkJOZ7pPpPN
8MEWySYgOmzuc8Ya3CnDzrXQhMw17VyTBFLc8m8HLeYlUqiXqkUpLuJ7GDE5xO5u
dC49Oq2ojM2naEML4nD2yAO4b2iTHBayjZkSSdHmGmJdF6uxrFo++KrvQdom+dph
Zq++p3aKzrZX0d0Dz2pnWxP2P5WqQU6FUt9PZIxYyeDtG0Zk69D3l4jicmbFDJlZ
DPIJ4Cvw4S18qemDbW5a+ltcCUBK7GngdMrd5UsxzE+NOyvtATbeINZ4zE8/cCcA
AHCjfoYVp9bjj2ztMHwIt1etvArwfkZc3vxs/85fJ2C5D18eTv5V1COkVfNsbV6E
9h2WO26QedsshzrefNnejiRwdNA8j+Rweqqxx0CS5X9LKE0rpj7/9UMlftsx0YiK
b4ZuB3dZd5W+9clPxoiT8wUWAutg3gVx2ZNKkvJELR8qzsZUS5rIb/rxqxKIeF3U
OK3uMjGYaBHPjJF7lzL+jl8AsLRUrUqkEE24gi+gO1fbKRl2xmwz3RDSuLVbD8t2
xM9L2BPiCmNtVUb2hnec6DyD5B9KHRBrSv3f2x3cYhyLotkui1qodADP4crVYEdg
CiLPbD+MuUexqWCJ5F4cXgmXwKrLN4QELzb8c1peG9L9jCKA/aqsdgogprzeG3hE
Zhk9nBCSG45c+60hyoGq6KBH87N6iJM3aQE7O+kYRkjukPpTTqnlXNXl/Qtq9BBJ
GqMVimv0OODD2hlAJvmPGAKCtuBQpKR/618J8cVDbf2xO+dayLiZAyaqS40XFJm1
gxWoTNcymwB75etOyyoZjChM0aUvRnNk8TiPh9a7tgpb4dpZHuMOzziK5vpq/mBp
0q5QQp8P6PzXYuagnJidXBAQWE1AIf4VUBEbNpcTMXz3sE9A4D4Bza7oXfIKEnoS
ZWDO/TwKHllcVvV8nfhWb/cFrmwdeSPu1rNlylWc1AUzl7aP3G8usZDeReMSJaIj
rGxRFUj0GTO4IkZjENvl781hqC+pAbVUOqMS1DXLo+lp6yPHPUKXHZa4PPQWkPpU
aoRSdebnWHQ7eSe8o4UdZHNStxY+Ld+a3xudCQ+wR3rifihA0bLUyiSm2aSt5tel
6Y+mkt0mJtjlGBOT0vGAidoXZoKbeckDSxsv1HZ6GPrCPJoVVBzhQ5fQS1D7kxoT
vNT9QBv0k+ZVSEBirz+2KPxiYLLDBYSl25KZpMmfWPluu2zFN/nz0McL7wWnqSN2
LZ7/L+tp23PyMsDW8soZPizz4bEjd+Fmeq3wYnRS4PVeH5Vu4e1CIU6gYrKyBDk9
cQDJe0REAoXm7yDYKxtmCbcpEcNH+71+1Sp0nPTCRjR9GLzCZ8cjd2VHXAEeYNcE
LJDGtFAJbBdzZHKF3Zd3KBWe5Rl4caTUzCyANcp+LwIv2dx6Fv5uSlpndbIqRlJc
honVWD/+4hLgq5xTzoHDMid+DxpjVF9fM+TkzvQzqyEk9Q0VkyjdKFnaOTG8Rynd
1NanDs19H362b0w4o2eVWz6E0uX8tqQU0vsITHx4kzoO7GjDHDmCMfzL23GtiZnm
cKymlktu9d9WnZJ2K5XqmzAA3RSo0XgMr3a28JCQURpw/Kj5SJDJ7a5Stw1Lyzbj
mL5+86sT5my0ote48qRrRuZLB92fza8CwqjJVHofpOu2S/ta4Jn5HbnkzrTkkPsy
j5Nx9Z0yMv6J9xnz+qD6dyhjHTKaPatO4KAsfpkqGlg3AZPL23Tyeco6NcHhjLua
jY3Rb54kklgmh8G9yy3az86UsTahteGmezTKF0a+HD1EvTutuBzjn0vDlWWmkveD
Soo9E3YJuxwX/YNj7C2H6S4y9hQq5+Oj24zq0ULuUKglt2I90CcTnvg+nGn6dH7u
j03MKVZR1+CHkMAk2P8BkPmyAJRcYk4oY5fSyst80GSQUvQ8AE3RKj0rJYwYtGVM
YKiN55ku+/026py7MKpfKLf37aY47U/5fwptGzD3fhYcix21Hl7dtkDw7boHnL7N
a3kCZ1p08qWolYA0+qrTYnWiC2Aq0SgdWAB+hZ8nBFB28CCfsgNfflmq6HUnGqio
4F/fugmhzSF6g6r7NwKRyEV/lS+z87k8cIK90uaICnYbmDhO7kMgENIuAcF0XUWC
tetYTmel29h9JgUcXif3oxeuA86PabS36OIYJrsO+lVuByTMJcxPw0ZO8xg7tzeH
S8ZjCFh7tbb1seeYE3TClVQ6jU3PtJRDlV4XZRcLXQpkLzW0ghZXYv+nuiH8ynPR
L9ANSi7Jp4w8jy4oTQ6w4g1J+BwrXQPIzSxxnlb7f+0PCANcsE8DyWVf6akGzHWX
InvFvkD7oKod10uMpL1x/H6UtlvHuFZvOeEcBawr8o32pMz8Pwtj14qmpaPO6Jd5
WcLFxiB3SeJZBKHu0OdqxCYyvjSFpfWZVQS9WDor2Pw4wf9KRrSty1vDl/QX38jr
Ghz9u97hKyd6n5TEVqtnfW7WDCYNJ9kBhUamwwSMVbOOv5iO8AFlVNawavyGaJaX
+pnFNi9cpIfYMudJEr3YbyNNhlUVrCVoN/Isbh+NRGeJ2ckPgSZc8S+4MYHoN2UM
aXBSj8zcmrPJAg2W3APVC3hmP/gKP4LMys6yjoW+7Q3NqiSj79blep1LWMceNJMc
rv/YU7YCT/ZSG8O14LqojP7JiZ4TUwmwsmVXvxq7zXJOrFOzDrJd/6PT1aCZ0TCd
NmbMDrwTp3D7XrrBlxUUS3yX4Tim7rr5k9fCS/sGvk6QYXZSETW8R2qAw/fecFVI
6FrWqcaA4lK7dZOZKiNIbmzq1NktXx6yWIujwBlkg6zkXTmINIXpUS/R4gSbTD2s
yYUno48cGMLwMBn3f/hIC+7wTalGTsyYgDCF22zTSKn5MfOkh8+2nbe9X18qo67m
qsAV/+ZZ6dy5JVYOyywiOov4Yytci4IEm/LLbjX/fXmf0coGFzn0a/4pdhiRTDOL
f+fXEIRwnv0gWspInXtKEIeDC0ORYLV9+Zzx4rhR8mim7Oxqb8Wbgy1amZcSrqcz
cLy1kFq8cN7EDArOitX2jE/Y4ACDNFtzgIwrTwvvN/jRqR0Z+2UgIZZDffMk5Gsd
AcmW8hrcfE4MihIok0c6gxnyEJ/+nQbQgxNhcRkRsxDp7Bytn0MbMoGnr8zEOp8d
uy15FNulWIgjgz/n19N/1FPzZT7vH/AiP06uAQnQjo8pDZj1PyRXg2ASa/4ZglcY
hkfEBBx1M4TY4VBQS7aKEc2hLu1eA/S0UO+gPt4D+qtOzKBJAIr4KocluD6UDaCX
uqSvJdtDKy0eP3jKrIVjkUMz6NONl31nb2QsI0ONbYAYYM3P4xFzlx2A9eKbm9IA
0EBAiQ09Hg/aHtMjRECofqGhnd3JN4sfTRaV+sL9UYbzlhosUQ4OIImp5kQdgXht
d2m54BVs8c1DBZZH1PuHrmoKlyMMIRm4NP4i33mKH8l3ctCsqeec/igEOzeRWllC
+wmqS7s8ZeuAedq+78nJs7MN+A+U0PppvbEdhLNxVvMzXWGrwPIUWR5TxWTwqw38
7Z1rsIS29P14MBpdZn22MNz/d+XQK8IRaqZ9G6Gt4iQ8hETxxi/IuBXPdllH+MAG
8L0YtzWR2OYpxhJ+Zs1vZbnSlYLNn3OgVYL0OUThpisHoefLbn3OLhdy6n6Jw6ak
/XyB4sgvetTQZFrhkZs+S78N9Av11fnpKY/xhJEVOpypVzI6BX6mjBUTIxYDJUQW
jisTkLPewl6diFzlXmcNZmzX35o/ai/70Wc8NbSIynRqDnhyKNKVMNnQFHCKVKx7
bVfBBrIe1UVDKzR+PvYLcdR5T/Gzg2xMOwyRHuJm9WHMXcRLF/Vb6OFTCHvFGobD
CME/raE3jQmkiQosrgnRh4WvaOL5kI5/369Ledfgt99GShbHnO6M1BljJWYBM6pm
h+3kOu15YHpA9wWsEYbFJmQrdMLrBuAMFnoI3RP4B3qQIq0huZHjGEG0YrgjnerJ
Fmtkz4KTyMy6vycoy8XrYX22fPqChpPVDLVpsl+L1Mkv60NSAN2hdkYW5N9szmVy
otXAO/5Keh/y2D4oSC1MV74TK8dLiK3wdsLqDfO9A+vxX8MKzOPeQgWKbiB7UTpz
vyKZnzovIo9daHI8IeakJTfq/d8oIsSngkbvgD8dIpttmoQ5GqtF3KhIOVi4zN6h
0gra0M7wr1IUZ2P8eqpz+GLBB8iHAPLoxjDkzUiK8T9qQG4+/r15ZKdHctmDmORB
sl92/XtWLoq0fHMFtyFQiiu1Ff0Hx6EiCAyYYDI+UPgnnFVt/47YNBtLn3wtIadJ
iYULg/FO8dKWMCY3uUmaAx/XmlTYrkJVFu9BJfBeB6Fs9bf6HKllFPDCvFYomUEw
r+SfuKfGbyCgZGqg7eGTNLp+xiGhPjWJOrp34e9+aqKMMq0M4/5kIekeL/fGLZBF
KYTxCTuAkbZ9JKZKYVtmcRiHeyXqIfV+ns5h9zor+fgJ/ajCrL9j4YEQ3EzRtEt6
886aMXmBv+n/q7tqje+SaQ+szlBHJtXM6zD/QJ1gClCyULJ4ozPhhsvT2ip1QZeV
UndBmAoFNwrzw/vMDCw1jAH2vp9+mg2ql7HBrqvzkeoLRL9u6IPpKkpxEIODLBru
CAGpI7r6ixiu/QsIi4AEw7Tv8BWSnHPlQWfSi2UgEL4tS+sRZYM1o/VervkzxPhB
i3qSfr6Wd3fpWQ1mOiC//mvLRb5bdRyBEDbcrFxH40um3CvHZK/wViXgm6cU8lbS
2KE3fc0bnJmkTjlPXjzpjzgeProV+uI8xZ3ZLNg+7iMOtcr3Omy/H9xLaWjMjDZQ
SrYKoulrIXgLFF7L4MDluCR94anCIvl4PJqpvtxXr21JXkcZHcFaeywIkBUt9BMg
giErR3/hAFAdCDq7+LTNl5cvf+KHI9G3EitH4/7F/l5vPA8hlcSf7nTNa7dm3Fme
fYJHUF+cE1nNMn8K/g5/aWB0xcMcf3eEe7ldgm6ipj1a+RA5w8IpkjXC9j8WjWuc
6TXWq055GB2wOXt61zh0+uEs2k02VMiNsHsounqNNml6aMrl21DeZ93hPUg0lzrv
/9XTgJJjSmLBpQvXWoXUPKOfvHkfPwNA9S+jvYYBNjA6lcwItFx7Ee0T3XBdEnTm
gcdurfVp7lVgneuWA5oehaB1nzpqwQkKQXsBnG5P7BaGNpj56XxM/CxYBOZ59KRM
TRWqp1AtgwHNOzMa5VvLHujNBC7OeZMXscKvznLZ5pinmpGS9m8Ksrlemk78+/Kg
USUU8bocDcRjq5xSHFy2U07LWnHNyBtiXwvHnDSgZQy3f+5+RkIsXmzyd1Jrb+FB
q2ErRyw5lXFdCu/cbhz1UPFBH6cvXZL0ZTAFWoE1WZjS4Ne6Vt3KrnCOkbUmFK5P
JSnHrCyBbnJz/2FoxgALRSy1uy35sH2t/RhJFS6RjPHU7v9FAVWofGHyqJECEN9/
BxVhmDdCSG6Ngrh/EbRQA2/5lImmN0DdsAhjUbzYXgt5FmluRmK3IsV2ZpoI3wPR
S/zYZ/iqrBgJN5t5JDzEom56Tn5XSOMfzjbBloR0ZkeNKr7B51lTuagRyNfKE4mO
nNAshWjdpnOqLOtR5Sfq7NQSpLi/OyZojR01l/NE7C52YYfrIWgyls0xANBOcSOR
skK19bUnfWAhtQvARL5toG3JpfULpOkgxDLvaP5Hf51Vlgc00hmck6oWlOfA0vTV
x7INK+wCO8zonZannaUo04YFlUfTZ+PGt/BFrAyzbG/ZRlYNQcCNFn1pJJFcJ4hm
WkOOXcaP9FPjlWW2W+ZY+tf3pcdOzwHhInKQtqwOVfbLXQO1V3rJOcpimj/xYGby
ayFlyrKys72+XEg5GQAvBpfoX+s7Nxj4pD7heNTWlVB3eFOfLpQrS2MSlNHiEcBd
DKE+Y8XnOQ5RygCZMz5KB/7SsNNP6fVLF2jhXjKM8vLVmlklrBsFFaNl85Z0e8OU
wQm1V5cfCxhZkWczghAtB2/kMy+K/8dpEiu2mZksvDqMu6/Qoxf5PXGoZBsZwCqJ
rukJTmOY5qfv6xzuggAL6Bzb/JVcOILzWH85fMopzjAc19fz82M16+/qItN/54nx
XGfvCCY2W9jSr98dXwmlNrsV5V45maP6Y6RD0MvmH44ekvcy1gbcqpQHAdgnBBbY
E6pkKUPUvV4SQsuCuwR6ODmkDhzQid7+kibJJhucpNKQEi9sZI5yzxkuIqD6gATn
WinzchOypBjRxw909QMfJPWVeSfUgxngMSmYsW/ckhPNz34LEGSzHPXyD4hPcuC5
RP5hs/Gsxs0ZpedhLQjl/GcynFdPdVnm2/QcHQtLdLKqZMmhP6WoWnzvIZtzg+T6
F1VDpxwXhtGKjt18F+357Nv6HR4zbwKUByD/+Vzfg7rhmDG6RB3E1cL+V91GB76Z
7kK6NvoaVuaLUsYCBzzK2bJKCdJ45VCPZn9Q9qcfarOewhh2m3tk7yPrk2RK/pSb
e+z6t0Ha8loPOaL8UZ/ipw9AC2Sds6At2vsPkXS/DWqCpxBU5Aw3LLI/1HC6fFS/
1sJJqHn008KiOUQgaQXGFDrBqXvKxiqkWrtJBwPzK2R9fKyFlrVyGU3UoIzQ9BzD
i448fWNhRz9BLoYIe4awt8/zKhyjz3HGA05KUr0VEYSJR4sOSLrbsPL0/VGrJcQn
ZQB7JeoB2zO7nDAQ9fhessnzCUu+51vAAtTL+/gqcpu7LLR88P42pKsl43gx0667
jWvDUaQKINm8qjDEsazpE8CzFy2+fecQzzBuGhm22cSq3S0vDT+UcLcuGJSS6fle
u9m6oFe8tHH21eJ3Rwueol4gGIhy1uGs8dsGCGExyGD0v1SZp+ThKcc3AOfMlohK
Eq4t6h7Qn7zh36OVGf+Uortc7u1lntRuuN1j18AQgfUjrHBDPL09+wB3SwT91jLj
SO4WY0q7IUa3Nr+H0ZusrDssohtoye5bH5BNVEFXcp1bVpi+tMARsukiqu5Rml6U
hWThigoKryQjydJJTWGiXM+9AG4FH2stUzQIvs7jxv0rEbqxeA6Z8oOgK4qo7pDW
vHVnZv24odpBM8wsLuKPUdoXBD9gERR77+Yhk2qi3IXjV1L+v/fRR6aCrpZ4p9w5
pUy96PiNIgAZT48DTw0zUPV6UmgXyuUdxrsU3yZSU+ZKhTiN5us13aliSO/+sVlz
F1na//eDCCXp51ady1qaUmmS+/wznzRmWwMEhggEJDFN+H0twlPpDtjQWjDKZsUI
IsBLoRawYhcKAxpknDCcjnaOM0VSvJBQWPcFmnbUoBu1r/V76j73o0SFIQLmHx9R
kY79M8mUZQ4yOC/uH68P4RR9Ri4pq/0e8ayj72Sz6MSBc+B0huzxZ3OhJpoLJ0Gp
488KzRue8odax06FX5XirYI8uhQz2kPuJmBcIf8ACmxLpmczwhxDg/IllJx799pX
yGF06n07bno7uAVw8XZ8tccwEUziL8nW3fE+kbyiauHDJ6cQFI8r4M8wDvX3H/1c
lh8nhLK4kxmnjmW7IIAlQ/h4R+kpeXZ33BjUtxxlEmMeTdBaat0Hr7dYMtJ0T70m
JBQNEo/tr43hcu6COl6Ai/Iwqn9gOK2y+YQsOjQOpW52vBLH/SdF5loeczmWMFV9
lYi45ROfq/Kaps0180juRRnag2xElKBXHLouC5NtL6jAYGQsKlLWSrqFwYn4m5Kj
7+NvbXwHonpud116iaqyATt8R9U9wmsxKuOlsGcrreIYEDvw4qQQZPuJH0jBC68P
TTwqlziI7c/kZnhVYstprMjTZS8iIfO8c58W79MpCyHVcdiPoQ4xsf3hFuIS08Ha
2F0D6alWerA1K+UBiAhh9ho4iy66dQiTlrd5/J1jkTn0qghQsHiZweNwrbwckq8U
bcNghdXQ67/z1CbxZcORuXNOJRohN6XOrZB2cnKCjP5fvmPL62gsSb90pxT0xqH8
mqnqsspCY7LPrWzU1uO0pCar1dGCRzJOmtxKZiQ79q57s7e+uqVR07jYbpUBgP9M
+eyfUa6J455W5RLk1aIT+zTO4Jf4r2mj9Zn5vKwyxcnOIvP8szViraYAjllt7NcR
/Lii488OPrhmr7YhkAZ2EbROrXUxKwJSdZKUyYK9FnAD326sNS+ELwdArt63f6TT
rRZoZLFHpHCe5fBUKDYQ4Xt9/dJQMY/yCXI7FGUTIKQfsrQRsZSgsviqOGGjqOhF
fpzESK+xJ9dbMlTwptG7tm+tF5L2GkujR747I4FKfgEaY2qD9sqHWNCyipQ6Dpxw
l3Em7wTY7zYTgP3Jfv9A48m8P7rxxDL9ZUHadxwAypeeQ4R3wHbBgMDmGLPeSBGY
AGMRSIDQUA9S1X0VyPzCt/MLDwzUql+W+rI2lvnncyOxdFKtxU2op8kOCSMyhXRn
8f5VskltPfoWgjYUFWp9PkU1tJjeIcqwcR514/YoOg0UIG7W1noOCgiU1R09HaBY
mf6uAyVVoa7hPUO1eoAHgoerPw3RRyM/8EQmqKVNdPNwUtzYd2gv/G1KPqBciFI9
BniLyQbup3gK5d5lQBcWiVCMyq4JR6FF4H2FzKi2flv3ROI8X8fRAu01tictNV5z
kvACbf8I12L6Ye3tW/F699pjkrGnNXpVeOHGAnwFLPcCio/hrSAIomhTrD5IMb2T
HPkgHhvl716eObhyGmOmmvl4sbs8n1bJfpYmtMbm+8f12Xe93npXwt/3CFjCLLvV
cJAUsU6ARqDfDyD0K5hQ/i3UR/J05pOo4sJLQyqaw/fZEgLuiVtyToP20WA/Jt3G
G2rhKWsPhtErLsStINH0XOBMJSvhH8Vf4QgY75P07IVv0bvP08rQ8f0r9XUesNKk
4JZIJAFAcDMcPukA2V3tbqQda3w/ut7/ZiRmxuJsGWNqAjKabCHax3jFcJH68gRD
lXMwZT1Ar7u8+Ih9hKdw9gBy8GZ7G6kLVt0A+MJgL721LlNGvMnif0VFJD+6GJR2
QLG0yM/HwV5ubjIWoItvBrTNNr2BE8jYiHLeCDYyvch1tIry+Xx3K2/x3vSEBE38
tKYg36efkL5wgH0mPmDF+IHamqYk4wCFy5w81B0lnwHswMKdpjHZ9KHOQR9TaeW/
sZmS+H71E2jPqG1vl5dBf5rL51xNmR8ZcvseWEU433fdEZJAQC5vNv2/yAXM1TZV
3diRJ2QB1ydx5aVxcqCIj+3WCsG+nZ6tLpxPmQJBkONQqJwVTF4HX/+IQs5iqwC4
rsDvThWk8TFDPVxnZKvwjSH/jf9jPsdRiC+VeaGF/G8o1RtKmQfFGnETICux+bzF
juJwD1eF+UM/U1E/oIUNAM29q3lmt3RKpLQHtdbNtPBYT0QIX2tT6H7/1npRm0Jg
v8GyPtZitxIE2YlsZZ5yOoINLWn0agmxjNth3uJOmrMz1/3MF6SdxdGIC8yNM3IP
Cydoe9ucpbe0PA4/sB7H5Ml+JPQKApiCzDFhkdtGKhtXTDoJ31Q1a3YqpAmdDPAh
68PnODF0OKBA72OtbbfPl4y5lPKRviz9091QLJq+h8N9eIRBAPLXjy2013xV6E59
4Wkj0wUpS5l3xlvIGHbalcvlsdcXPtjbsrjOs5tyJVIcFUQ2104o9gzKTr9JQuqv
QKw3R4ns1WFY0K7v1JPYYAate15EWvBGDL2O7aejEeurPOmJhJXAXW6+jQQDiitd
aXteSXLDb+SZh+gqvkpBAOWnIckqXxPDDbQHNvybCVkBE2iwdqnxrPpi0T2yTG9A
WrVrCnbJPWG5bDblkEMa3hJVUh6PRj03bPeCF8iYqTiKPwJqAV11YEUV+b6ubkJy
WFQPChpmC58rmykM2pB4MIXR+glJXGXjoTHqYzryZnOGVDIIy2leAefV5zh5fbVa
k/9NfIXz/lpfLW6RGPOgEviE9A9ecF8IlYI+OjqaZbmbc0tYWXzu2RlKoDweg7HT
3iGUJaWw/MQvbRX9FhxnvIGhC6u3Yw/fVdxO1kfmcsHuINXX+H62KBevwyj/r6aV
awuHDEUqcjedq09DIpaLwG7L0U7sHmyavxEGrmX6/4c1pYjNzZ0f1rS0XggsMPvu
rQbNvfErDIsEuF/Tl1rhTmTK47YpfV+FSRvL9NmI2jrf17iWs4aB1xVstxyWjJKP
+CQocbl8AomjPi02bBCQj/mCRtvbYYTheDVP9D2FGDDHw3yrhQ+FutlF6qB50ZI6
/QHNOv0eYcBmlkfvonbzJU2+Hp6knJH+hwCp2xcmxnhFGaVtqV8FtleD8kpBqsnr
/zVXkq0IvdbTisuSNGZvuiOjIsWImSwSCWkYwk9SIunpaOJajp+OufRB8e3dNF7X
4hX3dkc/82LgL5zmtcHs9qPaexUXz/ZJk+NCQ+8nIqeGQ5OLak57GHwwDL884ZYA
CC5vTwJFCSCC7DN0EolFzicZbkyFzcxqJsLiAvuEOH76ES+Wqhknw5oi7NGX6oc1
H+f5zz5WQrBWZrGmpr9CeZNCPUURjrQg+lr4f/MvkXkn3P1drdW0bpKp7tUW3LZ6
iSG9R7VLv7ogB12elSyc4WGTstVpdeteqUM5PA1eDgO3EjwTcJLm9TsQ/oaFwhb7
2RMmJVN55Cwvv4FHmYWmjuhehdudU9phHJIGcpWcilwgewXxgc1vPUl7MZqtoNx3
zsPOrEH0E3mwZTAgoui0RZODn2JrxBNhDBKlfjISOkz+F2VJur5PmKPpGFys85RV
ofkeHMD1LphtngEtZ9drAkGTPcqt+79Mn3LmgDSBgZTsbM1eZIQifw2XNJ8jRs7t
lzo1N6NzrMxr7bLg18cxM3t0LE+b1OdtYRRK7z8A31BILsNMgqq4xWxjX2nOKUWL
P8sMNLJ/y/EkEqvcMUwCZFDQdYtUIHazG9AXKSfd1flap9CYalw6cUeRRF5BTday
NaA+zsPv8JTgjMNmvw3E+CXCZZV5cAjUKCL3BXsyVXJbV5dGThIknR06MoCNLTWl
ys1n9DYSp8bE0GIXPhsQ7Bwwr7JcwJTuU+UHx8G/ksBbaWah65vCnZNHVvzvRLGV
gXJeEN++tddI/bC0SabPdL9FBPn2Fj0bwvXmpqMPFLjGTrpjMcV3nNUQAkb5y7W/
zyxWyB7b/kjctqXEf1yfK7Mh4eVv8CqI4E4CtYVQdv07KnI74Ams/Nkr/4kmNSNK
iUGWrkDwB+XHFRntodQZm41iyOAJLTd+H0dN+jGuba4Nwg7LglHjaLfVC3N2KyBX
O9R4jA6SFue7xsbdVrUpRVSk8tgpP/J1SDnnhNdvdKh0BrlZYCXj18SCc0yTKj1A
Ye0p0sZCOLrZuVkldD/lL+Sr8rC6LmE//aBX9edZwqtaC0js5VJP7vzPaNVrLCyh
ZRTEH6lOGfDL8InaS59UWe4sil+c24bP22nBjOXHJS1l51Sbc4f1DiiefHphbWsP
Y1wHBxKQzObM1nDiTBfO8FbO6YWZNpiOwmlWrc1eOD/UREecKKtcY1MlRkuwpbOT
9vTrg2RLpFtWsyBRnTm4Re1KZVb6bzZme7gniYSbDf8DsS5EL2YfJEGghzUd6OjK
SgLrpssodZCowdJOPLV6halUZyXJjc4RtY51fIGkx7ktgdmb03o3Wu8PBTt1yzrz
ThtpFifgcNLQslHfcBgZPSUGAR+wMvTNtC8JQKWTQX/iHh+Q3i/vrRGAVvMmhXRh
p/oGKkWJ28fLU3/VERlv7QK2Ypg0GFTR2Jfu6Q+i/BMSqRZf17NlXhkcX1aP3k+p
TxIE7UHDAIpkPGK4UWY6ABfE9hFmNdUrftOdYThtJ94armhLUpqtXC+yuogSq11T
gIYQYSRHZMe6jxj8TZ9izT7YFMcIIooj3BVEI7LBV9G6XOwsVAjnhOFs86N2NA11
aAAmSiFlYioFXKexR5DGiNBrwptbQigyQPFc+6tXLjo0/5Y2F3LCp3SNvYMvsJru
3gajvWR5dWKKkxsv5q4yBuCwVXKLAQJspYQ6pRpYc+W2W3SHzhFslhhCuzTYuyvY
DI3RwlBBNbF06s4xC4vQKjLmxAvl+IGovSnzlWhY9GvFmVc5ZqOOr+qWWutyFQui
RnhmYsdWoHZWPZ1JOQrvtJfWN2GaDKnCGDOLeJzYzbzePrv/Yj9sS0VjkX87EmvY
r7cmusqJIFoAwwCtggw9OpAUbvaY1Tl+KU4ML7jgwsU9vykU40V8OqP1IkF1spis
R29sUlD3N+Gc6kPOlWGyfgpooqw3Vb53Pk7fdexHinhgnkLi+dZLceE7jv2WtTwQ
MMWESvo7mUw+5PC1nbvA/dpj906KcVhWrg+5+Tr3+kzXf2QMpaw9gDN8nHioV61X
pIN8ErHyxHFdEpsF0axae1PYQGOD4/bxAZryrWQsRObJvYPUaChq00agiQoUi5A5
cf7UvZhJsYBuzXcL8/HG0BS0lXrHc8+79iuG+jwrNagXFxzZP/+4eotlAhiSGr7u
GpUpUybfyCxQTgUKPg0FxlKny4V9eUrwrs6gcEIrPb5zn0qQ7Ql2IWBpgE0ytnWA
gfqq+NGpgrE74CuTrGDEVSukUNL+4PzLiCZtaVPnJDCNQ6Nh84bx8tbyVuueZ/Fm
284CkWlH+cUNdgbfpofr4zCDY9YI1bDX5rPSJTd7/WucXJ7vakKea1W34wnfEbkp
zzU5dilvLmlvoIv+xfrxouzvZsEDT6zeLKT65OaHRpTkyMfvUBMAB5PI2bPP4Xrj
eD6p7JI/jwtr//i2U5LErAAGRti/Kl6xb42xhJGbC4ECELpqvaSWs2Jp3+l27jhe
ovh7pXNGxjeUBWGwzc8Q2FY8lNjPXldzf+v7dXmLXQ3cTL5jureWX+rWzmuyvg8D
YTKmyQOu5UQNx/I1eWj580wa9qetu+4VAxnihPS6RIzy5YyjbmtcaWUDnlhmW25O
mq+QdBzvZc08YO1fuWipXk649kzrYWE8uzu0rWPW6HwXbTxu3bJTkVHWmT57nY+v
TIlxDrt5PHA/Zac1ydYy94lZj6suwTYJcWtfEBtQ8TpvlFZMSYNpypiFe84DlC9b
D3ggiAmY6qOYo6Oaqg/bnPzIC+5U1bvbm+Yb4HOsewdt1aTWZL55xqF0cwSdoNE1
rjjXV21dL+EJJY/aNud3HcyQhu0iqQ7OOx7WkehS+chGzRLHDLsr+sLZJVT+E8Zs
guJ7rRvxt0B8Zcs/frakduprYDVFHT9fG3LAwrpD+EXjjxqe+/sQSZ//RVmrqumo
n5CZUu71BwqLl3dyuCPdFnxxBsAbbBJl/30BvN6RE7NfoI67PbZZ8WhdbEmcFCjM
R46XWV6yMl50qWOjJkhxQGD38Ko/5TxmqLHHKd9MMg4ybCZziHZ2Rpd6qhHzMeOA
WWq9lg2TZAu55Omt7mQKEpL5AAc+Fm7jIie6vEYc2d1aNfF81kvzXsHEw+aZJV+v
ykeMMGVPkhYFeS8FRXh7sgPMlhgO3hYt243lbtbze7tQEGfcJLeyt7oEJ5cgvyQj
iY0Wv88FkFBg2l2mB2KYOch2bvrt44vjUmQK0w30Vryv06Dnth/eyYYHEYPCj/GP
hCah59/geOhm6B+lT6UnK0pw5NqnoIh1Zi3s9p6u2l8YS2qYsJVmlIn/GafbgEp5
qs9u6QmyhJi/g83YfKjsIgsjBO4R3YEIfwwoKPanorMBST1jHhf1EVbAGwLknSUz
/7+3GAEp81RiIbPQruUdokgko8nUj65PpSh6VLooG1onimw8JaKjg/nfZvjc5XMM
qEey7oxCt/Sj4NnvkZz+Z1SxebfMoR/52b35XwRXqykGyfMwJa9LlYV+LAAJsnJB
zW7q95Rt+6uo7V+GlwyqQDuoTK1sUtytZ09gilZIXflykMqSvRpPyIPorDnhSZeU
ZqbsUsmGNbV5rcZnYL0QFEPa+XzRhEUdQqhMMK0en+82EX0rGcupg6Q1bExDd/aq
FtTvGCFrlluuIsIsUSjNLyimlL3P94+xRvEGrKVNQjnG0oal6lUig+H59kAnKvZQ
PJyV60ZmjV5DhpnQyx08HtTotryZJsDndscAhbaLbDoj+MQKwDG+6Q3kxS8LOUm0
pH3lr3aZSgSnd1isXy1FqMNGeJ4WshUwdET1k4ZoPV50EI3Wp/Q7cpM8vVTOcnCg
/BWyQXLUJ8F58k3NAazfbUlPMOWNhHGUFUXAPbAPPRw9/C8EW7EzFTUnvIzgiRrk
KofDEqJHJ0KJ0ieJoszV7aqiuMMvIzF6TTW0jsrYYEiMEXD9Lxd6UmrUMvZCC23i
2CDv2akTJpSsBqKFt52ZaFkhkmvvmDMCQoJYuqESUAmY+ooHg9JgTOJYTG4B9WBs
xMPul0pjRkapa/o1plNiZeAojZSOE/42qYXUQxYE36dWNBh4x5icGqcjCbKwAP0z
hs6u2mPZMeVWHP51Sy28X00YALrsviEGcMVfrmtETAoMKnIY+FrhcizzNwIKfBrF
N1FQxCQKx2jXo/anRo541zB18ZaSetPeKJxtKbuL8PJU36MOhPk3u1FeGXvf+gHE
h8L3BrVkze6r3GDjYXidxqHegvORhM+xz0nXW2DznSK0gb+stbTz3nmuS/N5itXI
iwekekS1x841yylJSahjvENgSSWpP3cJB/uHh/XXCqJOK8dmZpKFlTuW3DSLTgL8
k1OzisUxzVCMizLPue72PIoLH11uluEBT+BYEVOkm55Aqz56Dq/c06KelErgY/vz
5A8i0vwJQr9lHALHTfBsIG8A3xej6XCvUWhjqZWfmICF3CKIlsDHrv5KxPsxjnHj
MauC8ezBiZbsPDfCYgOKPCDsSW+g/oWDKxKUrTGYamlu64sOZu+jGTiiK8zBSNPX
5tFuyx2cvv4CUEChlrj1Mcrm4iGZ4apKbQxMLMZR/lQS3HQJCRuVgsAzv7+X0Els
spZXPz66jkfkzHFYs/e+0ujQMFcPJTR4AVFiuO9mU4ePQ1Hihi+vV+p42x+L0Yu8
/fjRnrpoDd0lGWAhtzBM4EXLki7puUWEg6NGeUnjfsp07Mguuri5CFw4QUt+6W1o
ZeYrvINzcniDSSRoQl7n86NPzwxSq2LJXtN6uUkP0o6qV57IqaBAG8Odsvb8Q8lS
qoXnWcZNHGATJGlttPn2RtJE9J1kyZmNWb7jyWbWfIgPM5HPtHple+Bln8GkiUNi
rnF/cSdhyJ1ZQ0JEN35gbYHkM0/7vDNzrCFyR7AqSlGaAlz/dfOnGBwomhE8znO5
0Y3miSFVTT/hlz6xwR5gYqyky0LOAYgQ2iPmfL6sUNm2G3VpNBdw/cW4+/JdBENc
bo2ud8XAy+nzOwouEVWUzR/uath95Ib/6Re6tlypNWU+4ixakjvhSgGSg+fSrgNK
90Z3HEuscdCCbXqwV75Qhdk8Jlh2Fpad8W1N3jqJm4Q/W8yX87tBhiWnZrNEskmF
SDy99WQ1T1tVdwO5XnSYcWLJYRuT/4rGJi4ZbMVEKQCWQYPIzBhb759CxxOVTdud
T7z8I+bPM45ozXMeNj9BelNkHfMoi5x4qfZYrQpLm78LqC2uyrx1d704jfOes5Hd
r18rEHtPPg5fGNyz4tPiP+c5jqzoHQwPqlQwtI7cYr+PxpedYb/15szJrQknugQq
2MW1abkSRlGp6cAjo38mjQ7SVqR2OBuaaFKUD4KvD/qA4PiDrgTvOUc7pfw79ban
+RXhs1ZKsY6azEkv8AIaat7bhLPbGtmlvVYRmfP+5rhmS9Zlo4Vr5S69rlFgqvDh
/rkVTDrcDeF4AFjcv/7hJEWkFOwiImDJxVJAW2ilCvhX+DG1XpjAlqFnNGvXy7uU
lan9mlnwmDJ3jHSXzGGF83GFrSznOa+FSxfJFnv5wWsHoq9xGMPUbDETQ0ClADHC
DzUao10SxtELM8mjE+yCxX16LogaQrOE2mGMcO4ObV2k9Hjz1po5xHxJBjebJZxl
PMYGgcQp3/KbOhFxdFcpEwIF+3rP6cehmGj+9qNeyRUhUrjjYlJVWRJ0kI8Px/wK
PZ78y74+adVICTx70scp3VBh+JVz2UpPCl+S9qaGwwKXHtuvrZrGdCiMHDizpJEP
skEodHDxYVgctkjAN36ZToz81ecLkrRxpTX0Oo6n+594Q7GoeiP2R3s/D5BZEw8g
0iXCbuvR00Voi5tFj9+TVQJQgIHEbuc5XzC2iWEhVI45t454aMt2idXChSO7n7/t
1koYbMuHAnjlshkq/OHECIv6Biq901+QGMTG2sUWsMjDNYXhCVc7l+i1jLvzpEkK
WY9f4JDV7523rjn399rMgXmjeRgRdTjxQ8kVn8xeN6in0sR8woGjZxGIczDC9FMj
QhqzK24f5JFtOVKrZ9mY4pUQtIAz+l3A8UC6Lp+BASXz5/YRIgpHLbZdpqIBC8ty
AAEpPvZ4SsCMrLK3Xs/oJtJt7LCYbkwHZcTZCfDOQSLFx5BBew6+rOt/Po8KKm9U
WJi2aGqyEfb5EQDeQx0+RXedUNNeIYfHbJ+rjVvVdfJQRXfsBU86G/csgrNv815B
oL60GNVrW4U8ubIHOB241jbtYSCfnaYp5Dfa2ZWx0fCubvukmnfeY+xzn95wo7fd
tyoejr634HAyr24DAcg9sBmrLsBZN90RxS0tVfyxiNOdK5nGr36DI4xRJJXras0R
mF4zgKfwwVhG49qh04uRyeeV5e2VVBbSDi5V+B1uoA3/q4ud6E1IdOQywevCpg3V
W6XRFb+WkqYd4k0hqSVRPanLcRUm5Ckqsx2G8rMB4r2GTPE6w0XVcSJwrkt8iFuk
er0OUz3l1PsDz7nxMaMWxi2gHinbdXvF1gjHpyoM5z6c8+LswhEivUdYZI2UnUQL
j8NekNGKju6LlexBXUJAoXCd9nai30yixo7yJtoys/s9YdcRyiJhasxtdptW75bc
aKFoBD/imq4CaKC8PinLvFGVwrLVjcSKTE9dfAVD4949Q3tm72oxh6kt16dGXV+U
4USfARJjNjAIkOPYWiRhIAF0mFT/DXNtjSTVbJOecriEpcZQI8w3cLvQuxjX5Qtg
bIRpPXNl6G6gCtNmPTkxbY+6qo/1aCcSC0rOKWtUIeyRD7/LxWeWKxR8cTPMEZm2
aX+jvbKpplnrhPnIrdzdeF+3q8TolpYY29LifVIPdai8LMh21Ht2P6Vm0sN31YLz
9nBVvgdfUY7rLLA2hbQIjqakJX+p/26nDKi8VX8DqWxFwqOQ3b5eBRBSsJjr+19J
8TJDuVnrANH9ohngUkasI/IOY2B0W3faK+Zvguy15RyXJi7QJ2WuTpTv7IO64FPD
Y39MH8px4w9/BkQQtTdkAsxDAw6Q75V1iVNpnhAe1EG1Jj+NV6IRads4Zo/0lfJI
lWUkgVNoS801F49iudx3+HejjuIxIsaEMsLcHshVShIEfY6HRLnl5ZCbW3KSYBFt
eVQOkZPmOCxAHZ1+vMTlayRyHaVdoSRTtGttO2sc3Kl3qTmnFNa8ZxCOOhXCZwqg
ATrcBbBH14E0/2W6xKR7/8DkFBVDnqyF/0ZHBSGdHMUbvZpjl8IogbPm3b0gWxKv
A/bM1fUrK8vsUbtKffom6CHo46kkO9cGyN9i8YZhsEsG6MGdB4DtIN2fXryEPaL/
YEtRsHO99ogylgu+ngC1/aVBL++3pP31nJtCWgVIxB+iWpsfbybLEHhILjIBnwmJ
e0DVdEalvXESQ9RfjBjzUpNUxO9WtwYCg79G4oBNJUqgf7QWmMaoSa4XKUCxCcXW
/F+2P9MMpMohYRpcMeK4LXBh5Y2VezwytZU5zmqhU+t5XAsDVQBcFVpnpUztKejm
uXdo3LTfiN3Dx4iraEK5Ix39t9zRemNhxNvuIcAG8Y2mSAjFyiByhVW+gehKT+QT
R+lpzzZSaT/1KqNOemYXo02+SOxaiMdyiRoIuUqMep9rgVFhU21ebJGVSgxctj2x
Ot3jIGRG9Tvu6HPzgdR7upcuF7mmcJ6eRHwrzHlhucRJcmwnM4MM8hiTV1sVWR8q
Kgfz2vxip8k54TAczJtDqhgVjXXk25sid/EdIo7VckG/+VUJ5TXBrkovw660uSP+
x/B2mVGS0/UnUdtDS/vSCZQ/H9ez0Ti+sGtXGFFAeEbWX8ALy+g8ocnqKiMAs7Fn
ugeWfI2qK7bl5wH8ez0qFMA7bQDyqREpwrRnvzLDxHY8eWIbwP3NAPABG+C7dRqb
wdiqdDND425xouI28uISQl7uDdsQl8Tce7HZYl/ZTlfsGSERSDbBuketVwPAJYg+
UZYMDgOTkU6QgLmoSCEQz2/7oSxq+LPiAfixojyTrVOJzWxpFbXDHkcxdC1lYDk5
9RySxdxg5hktoLndahit/vTwaNDLiYgPxmRleYDJWYva+5S8heKxMN4DvSBoAERC
Y4xPUDf88wTyTAYtcwURcz8RezE/jOXyUuU+T81LW6eYrdZzmztsOY9OwdTaR0kx
tGFFA3gX6cGNL4rzw0Sde46I+e0P5dktdLyPS65raaGHqvlsEK6Vvg9Zw+t2W3x6
AVqZ2Z16YPxFRzonmG7HJ/gu38f8g3qjfJU2cENpgrkEd2x51hcuZXngRpPnSMBq
laI1v3Oy7IAozOFK5XpRZLtCt2pwu0yx0Y5DeGtrvn4MrcvnlSJMcTHqtqAtu1tJ
D1Vbchrmqc/cI5Bi5yolpb4xk4YiRSrvYMQPBsvq924pYuxQJ35Aj1a/AAGpzmT/
aZjrp0FIL2qZ7ALD0yynJrOAJkjWx6LOf3uxtwSgb0SEGJBWOnyPxWc4kCRs/K/3
L7fnj81wQ111lPelzZJkoRRGO5oT7uNUf101cT+ydXgpS8k/GuYCs9U3DCSfZ58q
ydnSUMwvYAbMDSS/4ngaa3RFHjuIHCGHog2jQZj2IXEnH+hxq2kUEy3JLi7dmnEi
4/4G/bscPKxUeKlEH/dpXGZ9cdyDoqVQcgi7qJCGy08b3xKKA8YQJtaYmjZyrnPi
/YcOBu/n3vauAEAH7mxBqXZGfV19UXbRU3ExWFbia6TV5dPl/y4ABXCY98bczm3f
Mj8NBzrGj8/ORnMQFMeMQspUZgYfMfbVsw7ZwpCxN9tyeVKZUod5v5uiXg7Zsjl0
ceSOI485D6quNmhXaYo4XZ5T/ajDDDUWzBxCjuBsQxM8IxjCHVQDVFTzE/xECqj7
UYxHWWLvLs3F7l9Xn7FfqBNvBsh2WMJzV4cQ5lvnL6CmLGK+RxBdrUBzUui1B2Rg
S4RC7Ysg5FDsK2mF69seezihiqegGvi7OcOQJbihFKoPWOw1QSaXWrgVUTsJfEFB
cg5ETkWTCxva4lDqtEw0yOxEqgJfBGVMqFuPhrDVeEMJvU3OPpswYbQfXph5Qh/e
O39lDQ4Y+ujNbrxk+hmMTVkahQqKAJ6A5/Efdj8Zd/ygWdv4PHLVGqUKfr/XzPUn
DgrecAvwiv80BXyQ/vwUP8m80Xn4rTONynDdqEQz+RSWGcfBr1+4B0QKWf5r7OZH
MzNghgjviBGfefLfuEmh0qrUHspoB1BwWM3SUfpoxHALeTk5qxjcB1Lv3ZpkfItf
Y4muHLpg1NfoQ2i92WxNy+EzcBUntwKJKhOKjebEUY6f2wPEIygQTQYRNEWQsP2E
gF8DmrNnsA4Y/glp43WU73tjFcZf5ALIXDTwI3u7YAvs2xPoiIZ1h+d6KPsfS+4W
INbWxL5dKp8TRgoPTNwziM+mOz0l09SeWxBpJkt3nDyUGyYgCDh/+k2zlOOhXphb
xhk4M10fVSDfWG6uVsthFMRHhMX69DxgMvrGJPwlKSzpGeNrP53M3lV8yMoZauqO
6R1sYuWvGc5A79J+YpS8QRFjWww50KlEV4L7mcRMO461ZFITii0iEiGYuRuB/5eb
qcynA8TQHf8q+O3I5HCAwWNnZ9NM50WefYmJDuywpLEvUxaOBvYhzvqD0riB4lDQ
tTqSkgRCrKUoaHyuPtrI2UhdNmTZ946WnNml9AYbpmC41L3Hole4lpKL4mw4FFTa
jBFZhaQ2ioowAKCikSdJ5/IPXXv99iufLsebBkCfV+UDPcWmr0dcTT9RGKRKHOgH
4ejE6NYV518jdgL/HmB6jnCv3llVIlZ/q379GUFq+ZyIkMpfrm3sGaI9YFkJ4WBU
l26jfcDpKo4nYY99XkfUsbGfZ0AMFrOU4HFmk5BFewldaKvkRf5DrK9/i9xFQFWT
MNAaTKKWybjOZ9PehaSxZ4dECpNijBp7Tf7ujZwP4jj1JHlEbqPDu28QpivFQ2Zn
GIznUsDt2iQclfaP4HuvUVVVYO7tRbuCy0L1nLp0Rlvjzk5MRmdErsTGkbQFI2Vm
jibRkhv38M68KRhpScJXFGQIBkk9YGabdgc+I3YDE6P62KG0neBCOsLDi3O/5Cbl
97tjgRr7y0gc1JpjUISqY+pgGPf7J/Ss16scU50ozn11iJWNDrgrPqHAqHQjSBlH
7gPLWdaSwo2WBlk5T2Xxv7618I7UAbOoPqfqJ5ozm8mEGYpvnwItqXnrGk8cjdBx
t2msHwnHZa4H8lOIQ9js9g0xl2Sq92Oz1m6YCufWJFAy3UC2SxABOgy5SuKuW9MG
qD8p/rIBX324IaZThvxFKegXVikHV0Wa3dLky/OF3+KPp1hz2nI2Lw5VAlXrf2IV
Oa8GQteOE88VNtpsiA7+ISThoCj74YzEE5m2E/vsBCChpOKbLrLRkfECRgXYUkQP
WNLmj0p0Ht3XprsJzDCsY5etSw2cEsqIAM4bqfVRw7XqXOZ7dLe4h6gCRLK1UVlh
NxDXWa1QZI0sJOZKIr8srHWbGSH+jR6T5nV1n2KzOlNbVGndOdjzK8HHw7sKtFDa
qIbgdUtIxBAkYDUmkRR0UJbBILY3EhOQl5QuKuxEYazAjz0pQlR/LSRb+WDsuBXg
4vVrNZf0QMeX292HTSYB+rPEh98+q+szW32s0aIiimB7dQ+LJwj71/4svdql+Oj4
17YCw0864KCcE3jA6Poxheowe8Pjrfb4/KaVzlQtPx22BTIZ7WIHn7jszWvGybZ3
6vepN2qu1i9+K8skApS5vHvpsN8AJtwFJqjHPo7tjFUpf4UVqyHr3GRjjKc4S95N
EflASPZ1ERrgTEXgw1ZaM0yUTUPgwFAz1Jc1gvKnft65fA93tks1lDCwIcRrdR0p
YW9GUcXaeW58MM3H2SFE17ptA3PbUpDaJwK1cFMLab29twEgewcoIkiyM7RMhdkN
XwT+LmyBnp0KfWcd9boum3ONKp+JqCG4qTPh+lI+rzyPFCsqEdNgps2bfBdKS57v
8cRVRo0WOBilE177eChPHJGh4G8yUMqOsx9DXXzASDRpZSBePj2b355YlRwyVeT+
xnYPzTql4KB8HWj2JANzra25sK6QcDlW/VKewrs7j00Fk1YsDOmwaiHyGh74YgPW
afsXPo6uw8xs64wK2n5pDfff+lumCF1JNhBZQJbzfXgQOtMqlQPy8A1Rm7ZtAdAg
s1lTfcrfv+PGWloDvAJUCzjIxMR2oTNEImeHElgZJiSktjWTzkHaU9cA7nL8YgJ+
zH9d6DPZUi8hJPOffFoqWQeYMmbQvXsiuyoL5YtmjXJEgGBM3SHJoRzpGPvJv59e
GNyzjqR1r8iUlM1p7eWlHzGplLPjdTsGjRvUSRNGWcfqVnYfGadeP8kZSLmGT3yK
e3j2oP9mwwrPSQNSUVtjJ1UF7coIomBzTwbM2BH165agCAcQuibzh7Ovi3vH2e9w
rYlvBsTaVdeJRycvlEtwGjzaV8N921xxnPCKhMWmgjIRPe2g6t+isCj/flVq4c8t
dsPaYackWd9/pPwvr63WPoQBbAYAysRADvLW7mg5vU+zmJbpCjtCQjdwj3DCVhzJ
YrU1RSuQJCY7vJEgItWNrjKKyrxSI+32YlxsNK3obGyCMbtsCgrZO+C1Kd0NbXjC
nWjIngVkjprhGldA1fJO7rRyvwMCDwGtyADWqzDdk04CCIF0iLA0W3pLUA6/vp39
nTiFESfs4KDH49M+Ntu1vLuBWnLeHrEBv/NoQztoHUVnz781QNMM/fHVxCug2WPM
KxjIRvYHDYkANV+WnKJLW6PKh+HoJLBNhnSZJCmCwWdcji2vap9unVyahd0Z3zeI
HyZcnftUDWKT7nVKX+t7jJK8WQvKw5biR/hj8FdIXa/jThn3NFMZAcj63+zJSsal
aXAu8GTstOh5RHRI1i6U0ZKnOvqTrY0MqtTSKkXftb+Kx24GzS6LUuK8KfORsqIc
E1dk38/cmajhtbkczg5ecCm7rPYC+ABxi2eChsjLNhxquewTRYaIq1CdWHoMQjUW
26SYowYeRjKQSkYnos/Wc4qSvDzBRiN5AlkgCp+Xvs2jw3zDuiJgujUcwF9xMMyR
PsDUNQrGPoCHq6muMp8r8keZWOcEblYC0aDtVXxd9OBB95EujicZ/bhDZCWXIkzw
CIKe3/qmtxHDHyY0ODUwo+qt2rl8Z6H4Abwd+uVbzZCTX5OgWiKhffzjLOjG0yi4
C0ROhZvtdDgc5AhXYlQy1mF4OH2hNG3BcwEIHQ/DpZhQEKUfVJFpNoI9SaCkDry2
wISdmXnTaxFPRadKs0UEzi8L5bD67k4KbLpbdtFwpEKpiMC/OKvCl7AywXrcBKI1
VrMW055DchofVXYEFTRb4ySK7Iz/avCMKhwOlhiZZEJTZaIUOe05t4MOcXdnCkTP
Uv0/DrFAJBAcfrq2gFr9FAMdhlDPPz2GfGV5n+mghaIeLnBt74a9+WJW0TKVp0xL
7r4Ww226b/ECb6DsaGXSQEMIChjVmSOg4OzCuSsduYrucaNgSzUrZN404+pZ6uDu
kHAS43dIqM4HRasGo+TvZVaVvm+bFHHeGeA/QIH5u5Cj3x8ATJJ6y41IIsBe82a8
nbVIWMtSgPN4vD6IT7R5XacL633eAcV1pvad28mgTkUFLOyYXsVFOUH+v05w8VBI
aGoXvC2p/VgZbNbjSncfqBrH0SMrpo2NvOI96pTqXLIXlUoEam3w3VG/Jw00TwFH
aokDLPyHKZvof2w3TSvH16WQLHPf0odROn2sFxHRvb77MyCKYXrI+3N0YqHkJj6s
agjJ1/7TeNwKmYvwWkydVPkxNEmLzXgMuqxyKeAqsi7wyR2xCBpL55O4rtOBr1qA
rAjLleKvJepyq8R6VtItmPMJTNusVSxWjWAuMD8N1Z93aYhPQc3EbNreBvIFsVS7
AYo7zfXVg8egYQq8z5+DFo6hih6hRyDp3rDzzRX1l354qx6oMfBo0Cti/0FN1e2Z
oyyU3kJoxxsF0wEEpOh2mwBDOZwS6H/JvOVO7ijvr1TGLQMOA5Qp6QH5guLo5Xqo
M6+ja1VGdXDSr0lioykcPWom5MDXfQx2ew/anegPaJ2xq3mm1uX78oh8ekpdV9lk
eOI/sNBh1GfPx/j+6qBGZ3cn0tPTGQcpRv2ZuJ2qNEeqto3Mkdsru+17YoYPhZ+Y
FjRDzHt6+oqdfssfVdBX/WZwoH0k7sFkJ05dZSXZPCkNEQOUnHkIFaB7hprSVRN+
dIjfHDae/FINmTvMBxCRgmNsTH4ZJJhpnNC2MmMl28GUK01cs7ewtlJDzsFZOWU8
yh+xiLKNUOowPRAQAcBCN2a2/790RT+lGOsUjM/GBTHShuDiFaqkgQY2aK+Oh4rs
wjqoV4Y8vyF2w8w6pQ8DA8/Wa8ToFjSOCnzKOHqOU1DWHr/mjhUa9Phalawv3ZJ9
R67x+O3TVvedNpTl87AtgY9AFiMo0fNfxFkmUTtHhPJNQTam71alhDFW7WNXdlfu
3tQQFhtRenEsCjfdaInl68l8xCi39W9v8dBE6VqMInrkvFZZ6i4gz28sf7hmolHQ
9aXqXN8KsCEP9AVAy1LlHbtNGM00kVrCTU29gyftzpZ2dp1Uk+51PauR+Hack4j4
GtvSByfG62rRF02gMCtBJkcramTVA/KdIIVWaIOSiUnyD8q2qwQaD8/ElBIzuW/J
PebVFWQqLFBf1Ff7xijAOrFUJI8nBEiDaw2OVGQko7G8gXuCFSI7x3vWQEOxQ+0G
S5cjAnaPOvmEreo2y8asgp9arWHVuK8XGiYjmWdlM9/KsGjYXmK59wSldsMjtbCa
4+5OFgaGaocMFNJpvlbea20f9OGlSRHibgm+aXBgX90qhl5XXKySvSHPG7dm+1cI
ibRIGbBmSc4a5sE+64DTvLc6Hq4usbBb0srUzmM7ClLgD3mvC7hh4Ky//3EFTb+V
G6XJEaAi4ck6P9NjuXFqaMFk77pZK3d8Us2ktMbSkYioFwgPstQovgfcwBw85kB1
zZk0CgJsYDuYqR+gB5s3Hxasbiz6WP1bJxYZML8Tcs5QufaqqSt7QIFT60lXdBTJ
iZ3GNM/DyJkO8eUhtkKvb9uBTSomwZNWe6wPZGTzTjHikQPrdPYO8JiF/SlsQ50t
e1G/DFn3lMTzyquEIQ12FUULoEX0lmrdF8+fggJK9pyIIGGTAwL/afVRX7uVCVT+
UO3zOYxxqnG9Iz7gFwFtts8D52m3XYFWzCv2vA9MlstjSn9JBY93BZngIWG0atwt
aQZet2QcK65dFtrmfLKZT2SMH9Bz5EtAtTICJJt9WW0PPbngg5ZmnJxQqOq7Ywtn
ouyiuO7+3erG69LDChdHcyw3wXnRIrmqw+M4Lk0OkRpgcHVBv8xW3gt0So8cL0ON
j9xnLoAQvdogpin8O08JTJKX4Aqws+hv/X9CKnoJOu11CnSDwIeZRx5J/SWkUqcd
I3NYWERWUmfrrHeYVI2YNvRb2S9/9GfYCtM8m90RTrlSVEnoK8mAyzWZVx5bDa8M
EbvnAYeYmKSaAUamkAG8EF0qmHJvPxQOoFaPy4iA/5dyBIQks3QAwEstNk4UYLIz
5HJfdMqjJeEXKd1Vw1huZoLwAHlpbfJeE3vZUvJzVXntoTpJwef31Qzs1sHxcQX0
107kadqvM61idbjmCWgyvQQG27lCu4aOG02L1nT256Pf+ujoV7TfjeifD46uQ3WL
NsHhK1qlPN6a2cqYrgTy/YKryajC+h43xsguQyqVbdaWEibst3YE6o3GFH56FAK0
/WxhgqJVmO9r/oE9tps3tuaygjTbXAm54p0N9tEnjKaishn60eEkuq7ea01B/eUR
2zAJU5Qsprj6F9YMqkvgE7urDWpL1Hx0drH6RZ5FdQoEkW7AgncHNTkyZl3ZNFZD
3dFybxF1av1wtw8SEY2CqKIdYVREhkStI7Q2rRwgA2J5D4NWqi5yUwp9BMJgpbs/
iIRfoPrM1VGnFrWYEdlGydVdAbOyHY/TrKKQmaPCbKKSN/G0vUIxopBZV2umfcSB
OIuhC6bzPGi8AQ3/Z+LrOfMktyKcXL/FT+FOj6IHSnrfobRHpEWbj12XLUrkxvEf
EWYEvHHvqsSPRFJHp0n7AcHUMpBCwPDtrH02a5sclxBj9GoZUp2hEvYs1PFNV9y8
Ds79b4ik1i3imBJrZaKmCuvq2BQg31S0WRepy6m2NV37SjIy59q9w49TX/J2gQ7C
2sI3hI9KA3+oyPPKDGIV+nlnBK2X7uxInsDp/9/nAThOoxszukYpy3FHH2qtnYZx
SRiYUAPEIPR8PnCyZBM2aYev2dhBsm0dqNfAFHxek4LbtyRE7o2v2MDEVS8sgZd6
ecQiOA+3Kr0XDPf2nW1111nsnA6zM6ta+Z6XNROuxqeihC2mylO0pnFx8ONfFMxG
47oJhatsVLTDjQLG0xOS0ceLxTxoD/sQ/WR0bbehG1bQZtyJRK0RdkTvoLcwvAFw
tZ9Q+c6OITBuywTMWHR5jyP/9oyVeHxEKMxm/tpz6vKuNvRo63xxxDt7hbl2epMT
xsr+tGV1Z4+abHUIfZcCvZ/y0Ljq04pfoZ/r4wz8A1eVlEnhJx1447mmoJhqMjhd
iiFTejzO0UxWDGKD7VdZShc+Ho1/JdF6HmQdA2E7UZSNszoKCjwc8Dluzv5F9s1h
lBU4xZ8ccmWoUXDlH2tTyw3kfaX6yBO6XhBu0ukllwushliXsK4Bnr3dDhl/JiNF
RrNQlvuszKJ0AHO9YetHWPDVium5QUbFPE2YVQ55U8thnTm3m9Lhz8wwV+kN/juo
1hidSRPJoNZCo6QaKujIdebNqIdurw3e7jmsR14p3oWVdk9HGrYUfZMv1zpqy6di
3bv7K0beUUwilZfoLQIyvEpYvul41WoUH/80pkXYhnQDM4SwcUuFlBGhrKS/vVXG
3u0xzrXCmPiNp3dhhsiNeIQjnSBRkA8qLxxZzfoFZTif++phihb00ii1gVxBE85B
aiYXNIGSdaJyEbCDe8S/bx2J1aAzjvx5dPMB1cTzW4oJTsexwMmVNC+hDIbp8Pme
D9xcFxrdG92YdXq3WNo7nedjLU+Ahh5f9LtDP/mugzZS2n3YY/J6Uvrg07A3VGOa
tMeQu98201On7GZy6mWwdu4s1t1WyL7QcMbN8YFXn4b/SOTTgGJnir3JnDOaEDO4
2vIidtZcOVoGPFsGSsHaKvv42+HsRfgcCngcw+m+6zBqjEVVgV0XLhRU6b0NgPLw
bVVJy15iImS6GWzmXvZyiSPq/nDycDuXA+GFPGipx5HOLGy3b3PDC/yPkkYuA8dg
swqnYn0NqmHyd6gMX+k0IUc0LYzuGJA49AnxyeUAhQG4nXA3jYBMc5XLS+nvs+OB
T/S2RgGHatcBaWs1ru/SUnySPItkZgGmr2HWdRvIRAMrMa+JLGVig6TqvFJOdC9A
cAMSMSNWk6O4irUlMqcPkwxg+3jE1ecBj67kFFhg4vRUsQ76MMAhoQD+xbAks/oH
R9YmCDFzbrMMp4P1ugKxa1HLqYHIYhBOOz4RmlTsMI3nldhZ2Iv+aSWBI1idzklZ
1K7+adgRU/GMvispTnXpmIbYqqE22DDxTVOAH1wL3p2rSqxVZZbubFTbWKsX0/bi
YMSYQNBHKbTBWbV15Cq7+KIZzTHCJ6QroHhqOPz6Vnok3CJZTsqaElF26L+U0Ie5
nKscHegh0DFWlqX363SaQz85ozz6rjIJWQa7lqB+/aOFcRLMuLzYt/V+++wKr2zr
iJaJUSnZven925DhWkcVw9BrBYBXV1nqj8/15wVfb97kj5IGjsxPwF4meOvu6fW8
85DbHYijxWkHDmPIIHp5yf2uQ/gjz/uXnBDOGwWuXQp9VVxxDDQnqOAGRrPSF26L
HoBtxhNi4NbCSbwiUlirlXTE9dKnqmVLi1BizbfxhtdnjYrhIPqJlS4JAbTvrWlb
WFl+QNjRCe0KtG4rH8/ARq7/4DK9P1bIu7zOQz7EmY/r3KGMnNRHe8w9nAHQDYM/
meoP2X7b3m9D1A8CEIZQqBtMCrw47hXTgKlZSx02xlxeQsIphAZW3IZmnvpOu19C
9BVNf0BK1S2+slHrgPkQHrQ2P6wpJIIHoDmQDaGc3Rq4EKn8S3pLUnbGtpovQdu9
E9oywA63KAgCWvTllIyqaBTPQTuysasppvSll/3KAEMWey3Ea/nww1qyA7zsy+Rj
mLat8I49m/tKVRbTYYYwvBUpAl0PIRB60snl4dv0rzUmOnZOah+8H7G5+Nyjsf4k
xPY5lqa4FJpmlEtx2/5tWczgQrNKoOAHA4IbvdBIktmmNDD3O682KlO+Zzt3Qofw
s5Jww0i+NdX3L0oPLwgv4sjeCHLo0NPr7E6VOB1NYtELMEbkUwp+dxXcE5ihwW4S
qpilEpKXavmROqIZzM8q7VyjLM9/3GykzxfgAPnDRGdvuQ9xjnMDwpY6LpiTk1Mb
PGTk49Ain5IRtMpEW3/Mxx+7NzKIQumpPG2tfajjjt/MtZLHYcMUYnct0tPdAucj
823KMkD2JptAZNykl1k/lI2nC14ibvEbWjfAKpaEJwj6FpwKYy42Lugp2P/E5dvV
46a7Ub7pF7m6xTHwhbCV7U0yeMrgA7Q8V4Sj5g6qMpkSMxV7TjQW0TJLuV5TnhCM
Ub6fwuKm+TsduE8o9xMA1fcgXi6Vg3XDSgsm3YYEP41c6gB05IbMplKgKKvmR4kH
LqUJdjAWU119/D/dCWG8lqHB+mg7Iqu0cPCWFeJPaKnLzKBWHbOiqPiHPfxlDKd8
jm618/L0JI6G7KH0tSA4jImplyWdTYz3+FjD7KCi+8GUN/e4cX+MxpTayPphQTF8
ApNw6iF109TwBU3fEpGfIRqfdaNEuzxqIJQAbe3Pw9UFChklDmlkqEqfgG2FFEMb
ltjtGaOZY4DxZMgCNns/8Rs2Cd7gcimyS9iJYwwmDuWpnfqUBx1l6+mMy1qhtBvW
nXpjS6y/LoZa/rtOQq1gupvDER/kQ/y6pc0U7geHw4vuzq3NaIBrcJ1k5bvKyUub
gnwec467xdX6ZXpt9DSJstApH79rn4SV5Wiv1xA2X/SVam9zWLzEv3qmwqcqRKUS
BM1z/gwf2RAVvuyUOUPsUZjJ+RhZ7veTZpjz1A9jm1Xcu0FsP8ay2DUJHdjeTjLk
cuYh/uDFPzHv6788JmqmcQ8zDuS2ACCruJhJP4OP92eRDdc9lyA/k2iSXv2V+FFl
Vxwb9zYng0ViNQMrqyWpsMVXrUddP/JgVyiyqmfNm3zmIoZn4c4uj0OGSgnmjtOb
REdPWRbMwC84jFOXmp2Ni8dfzpUT88kroU65UGl0CNczI3L8LF0b8YCsYXhECb+l
ROhfIVhAyVlIkYt7sa47RrVjT0n8Muxl97FHnishi9KHlCMoaxWPslshzCvi4Fbh
BqiDbD4geFWV+sB68jrflbLtJ0zX4hU/rOci4oKAbjD4Z+td0Vd/YbzlfP7nslvj
VQJtuJea61wiS8K4kaBbBsrqwhPVA8WZKzxjmkTmgvBjAgtYnxBY8hlVG7mA94So
cHU5j7MFCIolz8hi5lTL/NaaCW3m0gVnKIKCW7Jq09isL1zIvokgorXcRcDf6YND
cS+RxF2vT7HuTQspMKdIBB/Ea7c4Trijp5QH7oKT25+RlWUWxl3ZrV61UAol1AjD
3a8yWqOmQ9FCwrZdo3deHwvJmA/q7BObCKrahC0BoJq2YGeyahbpfqUVs84S+/VU
BM2eo/xdefdQRROgbQ+Itjs9Pj0pqL+5ijn8xArrpqELbKW7U514j1dnDGwiJ8RT
3Ts6/sqI/XE2WxEg0h3KS8gYdCMQmiJ93Ju19+akNXnM9g0oeUOAwuZp9FwBnEdt
2zZUTM4t07xbi55Jn1b+VFWSauJt2bH7Xzf0oAGLh8b0Mu8hiDNwlJdbBdg/fA1h
Ae95kWDDaZ20ybEAD47GkUn1yfwzQclsKEdS7d9UV7cbwzS4pvkvPqJVjF81Jkx2
+j0ZNJsY2wBe+snXm70E5vLdcv+r4RjTh5lu0nIIHZOdA8sWbrG5+l7T7JRn8jmc
69v3Mb/+SH55+nY2MHwH8SJZUKvQ71aq9U7goyT9Ar1v9p31emMMzbKCnZ+NVKiM
NBDUwfhsgv9Kfs+qFT2JFKZ5Jpy75Vs/3iWIpF1E7ELo88XpQvy2GmDINg3DChFc
93cudvRaSTqN/279+q3EDgrxlgp/pDN+fwjEh+tyoQYXHwB0OSorDcFbSo5alxpg
ZlJAKnvvFI/mCtrCH7eMZcN7sHDBb3Qv4BZeDQLMXGPIf0yvK3e09ePrH41gFEEq
5E82QbvCa+oT9+nzYck4qD3yN68C9xxfymuXv/Sb2rxTjAyn10laUhSdpzZjxV7S
900LRjM3MmervHi0+/pcM0Fq5zzp+yl54VMT3wGUBJHUDf3pIMRussSDxv8jPuMm
T/Z0qewQcaQLq9ceMpesokjuQH4kgJt1ynxXjRShqljfXHzw8ix+CY3we3ryfICI
X0mUkxR4C9zeWOUZwWbeIQzm58E8lqCUjJ3+H5qRczzYRrrQpPNE8geVAWwoXrR+
9TsFlBDVGAJobvN6NRnJFRkSET9FnpFbuKxYFyo+wPd/cAZkXLbMnoqXrEag3y49
WWBYltwwNPjZdSYTVYog6UOHfVEE6LAOz0FYS+T8zAsVSuyLpPjCb8pONp47/7EO
QZXW23lI4A+rrvdaFxmJb4vpMTIAHEbp5dLmVUgI+b5mej21Svk4oh5kAC/2zseo
W8QmgsonxPismuDtlzMwLDb/gfFcOU4dglMaqOiWh4AW+uougRLNp4NGTck0I9JJ
9rtbrbnEb7BY5LepNh7jg5svQEdoOMD4wKkWvtE3iyyxZtWdLb8tHvcHaa/7HTMa
NUR2WE0hms9A4hNb8sOGw/ghWI/oII3pBsm37uhPytoyr9fA6TMlCavGcYfArgoA
SoqW1iTqTeYKqHvUNTCvAVWAGMI/rxAnq6uLJUWyJ0A8USPyqyYiJkpxhiL3Xhrw
3/8HRNxOf0K2iho3dv9vHBEQRHEMOR+ZLEyMYlT5Bu2OdwmR5+PWy/VNur+T+7IK
K+MP7c2VfTKDyJnqaqATtWjtCFW8xPY/zmqRRFrHf9XTdkzwbHv5h78tLxrOZZLE
XGw+loFeWJUUHYai7UMZUZintzKViE5izoCA4DzNRPJSY45kpJQ21PLKcxsrr6LI
winieNTih3A/YJxbN5kuvrFBE5f14lqwxPRe5UeoQP7qVdX6kSUBcgPXavC0OmI2
GgeZ/zr9mzXrp2Lpg6xcA0HgOYI4jmc/weAUmNbv1OBH/c3a/4wrHM/OQXcF4ux4
nhXPEhFLGEoq6PIHgknHd7/rKYEg1+/ZORgjgV276a2bXkEh6T5wUoCPi0kYz9aL
+RU1mHAKd17RaDX3PtlBFfTjas0PHIG4Hnd6k73GgFiZMULMx0baHWhXNeCasUCP
u9p3RLQLMpo398+Eyt7sobgwmzxkkzy19d7lU65q9QCnZuMsnuFHHzMWv+bw5rZ3
07wGZ+ZXaxts7uYYZV1WlgTbhj6O1jxpCaY9RQtrMLMfb+GmHzVPt13b2hmTAifD
4fZewd2FjWV5oC+z1uDc+jk6KzuZps+pja7hzwlLDGShGZN/FJLbg4Mg4UGyxCTB
kUNkI6hoddkQB9wHnYqxx8IxxhJS+eJiFVew6x6e3xTCHSfYVx/xuPskJpIrh0Iy
FEG5WE0hNuEeXvCPvb4efazjLzEvOb8fkKJTBHPkrwHR8RSKpj/EAOfxUwnkvybs
vQtgEH40bzwLHwGDDponiBjH3XqhNVHnKO9SAEexzU0hGSFuSmO4o0egCf1pHOEp
Rm4/A9iZ1BgRQ5tMGGWwlxOVFCXSErs3+j8X2kf7JyWx3W31HGJgEYB3wuuiRJHd
xSE2bgKDaGRXdGS8Lp3pmrMB/Bah7hf0Pa+9aZlOb0j6CBcPljlYyuypIdv8hjVY
F6YVEYpqRvOTtmHQsp3r12dmeZSuRGvwyRsOtXZFbvRVvj9HLUbVdVcknYglSZPW
0GCCRTcCIwvOOjsYLRG0sgMkv5f14qkEKP5BHqw8PFXXu8T1XHZB2t1ThUtCa4OE
pw/PKc/yXYb5s+OjdxiTt5UUMBanTC+ARrQXOgdM4E8uyS0NBcMyL6DFHzgwGEZo
2YRkQ8qnlFtQMsZc/CG4g7j4GXJbJDh4KhHCL/PJNFHhscrS//JEaVm8V0aZWhQe
fPB90mWhiLdiDQxhKd/leSFiwSCAnxHimhePNTm86DSHeTgLv6kjukqA3cza2xpX
0kld8NdsMEzV0MrwLC/QqkrIv9HEPkLehPWV58aQhylCvR+c1it4YfyqrQUMO1a4
83kGL22ZyzZQiib+YlK7KFHeyAu4GBdgGf8qbsNQBzSdt5ol22zZWjmQRC12sfo6
MgoPnRML9TvX+IlC1nxlKo3A3/HoQy5V7IKLRexiQx0l51fZ6S71CakSANKF9YhF
ZsSgNtjle1L/XS+62KJxfxrMHZSbSTLmuyRGpxUr4Oc53e+sECR367ANWFeLsWgJ
PrDqdRAtTdPGE1T0oszWJWl2IU9qGP9zZwD4WdmFycqUkJgipsRu7ANZ+B4gceGp
LH1Z5hUEqPdfElrYNn8/Fjxx6j3DfqVhyFg8xsHwUXw8Bg9PM+44UFq8N3XIs6h6
/FScwKWic/jVNhFX73MGS0p95+XusM1tfPY6hwY1AQFntqSGzXdyd6JpZDkvgCyn
p/fhEaLAct5SCJSdu3gZSFgoQt6DHrtSFqqLdVuYT3S8EG/N6sZtWF1ePzIUlRn8
zXqazN+48MjpCI4+4hTr4irpaUjZPGofpmNZtnf21knhe1CUINGNOReUN30pYvt5
7PIhhyY3AmLkd0KtuI1AVTJhQWp9rvNSrH27yO/ugpKlemSclS8ZRwXj9Gv+oBqs
NafPNsKDL8kVJDuaa3ie6HYaGxfIQGagd7Z7X9QlDB/kCBZFTqU6brvUOH8+kymY
R/EjxMgRKMZXIeHMvQAUS6+3OCMBfqGcyTxYt3mFd0viMmwCRPXTMg3G9kzyHPpl
8wy61sCtFuCGUUbjs9m+QiNjLV/FjqZfGkpFpTPCjyBgDeCtAXm9ra1vhmN/TQcE
QCR2OCcBa+pNMmy6J69+4l59AaNO/KYLMVuIBZOz9EN+AYx0MRGlAz7O6KzZJzF7
GEP5HUwAL5UGBOvw88CNuTxEZi21ATJ8cu8spwEjh7BbrNOtn9WQLmtfwduSQpyj
AAbcXg74GZzosEKkkHxVpfRxmwlEFz6o8W7xtCu42cjxOgRHi/fZqPrY83m8wx4n
4ywUmeQVvfiNTEkHPFpXId7fCyzw/rQHZnJIKqoifnFcvwyZBo+jr/jXZsVMDB7L
b5uKqDM0fjeT/2G8ytCmJzYUznQIqLe7DUXXwP/LYuq8WKpFPjqRFp81LUZlsDxU
L2XW5rrBedpAxoUj71rEax9k/5V8R0d6D7qhf1HGjcewCCdFaY+a9aiKi9mHnCZF
2vBSLdOmX1rOU5AgOMEhJbcZXascJ7fULTIZO970aLthUIoGPW8ab3KNG+lt0gEq
5tNLYSAFDQrhiFs9cTY1V12FOH99BgF1uI/piC8ZZTIRIrJqOz/A5k2IA1wl7gs9
4CmPIoJxIH/ubcrl7o2raQGmsF2HyTivOxKUwq+9m2ugYgVBwDSjksH+dM4l+ypx
8LxKDlhRgqHeiMyYJxnedt6ckUlbqBosYukNiSq7ragBXB3LaojLe/7NObUO/Yc8
tua+vTIKcnryhZctq5TjO3HGQ69YLjrjJg48r0CSgz3qEJp0xzl4+YA0azeNYGtj
TKexuI38PPzbao62NUOah3ElZ/fDEI0EDf0QmPvpx4U/mvtES/s+dO/z9054TscP
J4+sh8DoE2ACCgFA4uSiSVfsCoYyhMfuh37bs9wqHkUUNqIoT5zx/HCeuz9OrAo0
3Q2oUWJq9ipjhDAmBzJFg6hBHIi0Zc1m5aQoMKkC3mOKBVJWabeAjM0XN6895RUa
R4XaaMP9J/jwLnuHrj+tJSsZpSgmQgiDvJKnBmm3aLEU/2YA/xU5+VddPO16ht7T
eBK0sjJXT1aSw7ElfAeswsu3Z7jj4/PIk/6b9cmoWBvAjKWrpvglByDV+JDw3ho0
iP5fR98Af/g1+JtEi1jM6WQj20O7TTYzgBIXLMjxZmB3wfWfsClY5SrPU1IS3KDS
mZxBz93qQCtraqfTw+gmGUikW7s6KkDnQ3gabWG5/88TJZquDCYWBj1x9w63j/W/
Sl9vjxYAUy1TwGKNE5Mvf+8FYBU4wu60yI4ou2FnCg7rM3DvLagS3LC3JsUNAmWt
g2v42b/idXuclk4bZvtsGWi1H1XllDhKGtOCUKUG6c28Hm0zOUmKu15EPHud+YT9
VF9IHsW5imxwH8sfAO627yAN8UBtKfbGjsj9y2ddQFw775Mqnb6Rv+5ZrltJKY8y
nUlxBja8KdFxEcYo8MfWrse31WDlwc3V/UqtZo780vpbqn5Dr9km3/uOb6ZCMUsU
sA2q/fv0vqh5bYT01U4F2lYBA8u789MySkDHglUO/H5LMSxhKluwK24m8odXics5
Q3KO3a2F7boMbs4K//24mbQimT0EHHlQcsK2jmmJ0jCR3anIkOqqDPqtEI12T0Yp
Clb48tsbGKsn3K+o4KbuLmr6k6hHGP40zGyhE0C+K0Gc601XOMbWHKaPjhEMKbld
pwiidUSD67FVxg4QjRA7zHqvNLaXkJcGM6AfFo1iBm4tHlf1hTwjFc//YhlJ4aly
1oV1DeLmxG/42zEWY9oLVuRVe7QBMHpFNi8AXhadjfEgYrfBTZbzqzIAiL7bnLPy
t8EsUifViS1gTTTkJVqmQMZzgAvO5YRz/p0ZcRKOytukJ6NlTAjMDK8sPH8zXutp
gQFj0cUeSVd8vYW7JO1vxdAgijb1Avw4owhWFYXMrGuhMftApuHYOMgJH+hAbPEb
1TsZDl0H5ar63/dnthT1Cnu7lG0472AsO6My0VtQ2eJHAjr8pkzoc2cZ2WjBPyoK
VzwpXUFrTJSzBa2ywbfxGMD42k6KNMyJy3PUkxP7DS4XeGwlihYiJteaHlA4c++k
wUFm2HnYjXA8ozi526Cv+0WgOC0dKk0FqVkdgABs9Hdx6YsRue28ATK3cLIINvhd
peiBBPfUoodYoh0snRu02VgejE3ywNbgAkBOltMKaHa0Bmx8r3VXavfdXiv5fdfY
gtUCP9yGqhCrsUNlmgsYWj7tkQsY7wj6UHPNU7H44TYqeiB63sqCl8/TQBRwFWv8
4STYhuuQlrgedjLjFg/33r0vmuNCBncmLzfCQqkxcQttz0ueuqcysEIXMP+fd4Ou
lOXWVxw87jItOGarLv54qZKIU0JKARQes14F+41Hc40O2sRre6ymj7ed1hMpvNv5
yG+a7Z4vYiDa3ajfj1ClziSAKWqjdHoP1RzpIzdim7nm0FqlmwMZmW9qSyjrGD7T
TGfghFc2ozmcexmPGNJWSI2/Xpiq0g3sGoJazUNzhDPEtE2fEgMNEjwuhD6U2yM+
bg6HX5l8XC28rrCDLfewzKdNXUG3XPn+8n2TwX839+Af62NPa3P5U/pIYpb1MFMp
iECAudsOKXBS6qHWUyu3PE8cn5kc/OiqZmqdYEyyPw4HhtEgEhFlsg4Ka5oaYtDA
rceWHN4UtUltWJRXjEs1XtluBY/Vyfl77ScTwLsoP7j/bxIvgeUZVFKqorXoHON9
PYIZeUQa7twCeikYuNYclu816BSluQxIDnPbjlbP5SI2QQRS3m60lO6fctVkGAoN
/uSpifBcgIvn1CkhKug+VNkEzyYwFazz1a/XJTDmaPCNVoRgiXB05zobenLIfzQZ
aViP8p1/QQlQcqYrp+LzcEt9FAbIfWxFFEdMUtXpb1CIvile/rbps9yMAzbAlg9i
kPMCfsTwhl3i33/LgyzCcxan6zaxxW5CwLFF6dG9fmZZB19zQUs9Rizt+f/5K7yT
95TAg1mXnkRtV0tR66EcnnZzw2RBXLW8PibxPwu4YO9uDNezw72fXNGZ7MXJhdiA
wap8cInl3I8g/yjIVFLaJWITtpfc6PPxvfDAli/YlLOghYXiSXzbvGv/DqsmwHsm
hGx+B6cbOuDammDvuLcayh0EINgaaWbw/BMiEh/EYu6G9eULQRY3GLXp4JMnczgz
XAJL5jCD51jYpdb2ik7v4kkrhBRSUQ0Rn9mRsg3XKTWls8lFyI9VwHQSm/jtISRw
eWvKFCdTr4c2KDz095SnUZdgV2b1gEd3Yq9tg7uqV0fZYyu0tU0BggsCzkI2zSzG
C9OZsWkosAFrXOqMpOcPNDv1gRR68XwNnCr5Szhzs5rUf6+Wv154Hamzb+3g+rTT
csTRzQXsPqf4DKSo2jfNtbts31qbidjxrDPDGEWwhWTxAsa1J77/cYdTTk/rA3f9
m+uWZIrAfecn7LOlaxwzW2vvAGmxn0CIHjYRdlO8hwYvTOVowV62OrpnsvjrzSHE
jLpf8iGwXp3vk2clFnrry2n18+CYD9+txdz4xBhGSggtea3MPf1ztv0YGg1BVksW
gjPuelX6Jz/pdFWOxSaJlsK3GiSPmtTAOlJM39je2Y8sPToLkJ4Xa0GekBiYDzqm
7oIvgSuEBF23RmLChloiJdwcpwmnkRGnqDX/M9Kr2ikQyQGizvS9uPTDvZI5srla
0sftWWlsd7qjnMTj1BELcnKL9kABd37Ba4hSZ3MPRYt9Nhct1Sll1N9rEvSBTqov
8GU4dzblr6vy/6Zve51Ns3uPt3ApKmv2J/ZJzHa6PvOxbfRCb8R8tDZxCLQEjUYz
R4xZA3kfN0/abjlGxy5Q+/q80xbwvBhrA35pGJVXW0pkNabU/Dsk+q0MUTdsIbUN
+KJCo/e2fjSBGZM6kqrdNItiC9FZaOy0lNeOlPna+GchVK6Th4nQbFq/CYTIVP8N
ozGItFU+M/b/LLM5AMsBj8CnwkIXsTfpL7KwLdObQPSJwRjEcXNSkc4/CEEXITxg
hwhkoVd3wBVXucZbDPCUzpO8h2r4G97IOOlMAWKXaDcBdOEOShhx6U5ejHMIP0JS
8fmHtyWLh7vGtpZ3ZAKB9yfrCtCuXE3rz/9yEMyLFUWdTU/yot2zV0abh8xGrcQ5
Abapm9upQCMMO8/UJS79DU0JzKEFvcC0cdnpA/NBV7AFD4CViUJyLX6SAyMPmCWS
svrN087G2qxWcuzaYr9RxVtwgnP8Uz56iEttNBnykTc2GyAZjGbZdHvG++oQKOKH
8AFOqIARWxt9TrZjsWuJ+kJ21Govcw2eGwUOWspBO2AldXZZcynapNzFumgAFVWK
BZIuQ5ZuUp1CKAgVm5VzmP2eawZn6rNOzuBetrdVdBu68lR1Z3tQSF+/8QCQSnFb
mDKiWOjvie5YOlVhQKQFxOfNDQXeBz0sQ/hyH85Wx1mU3Fk/CxUeA1XH61SdSdnL
znoeCXaD/WAYJiL4emmcunrcQ9UqEksSbk9VwyuiKpxPOGmODxaNbREQkYb73oHI
HF9g4yuYC1lVq74ewlJVtwMd/8c7clcLN+udhzqbjmc07hFU/cGR17eO0AeeVQKq
Brt1Riz6KzDAN38ni46OrO3EVEPva8GchHP/sI6nVHtXP/g/wPK4qjarw8qWahmV
6Kdtd5yER2k7IevjxUoE9Ciq1XhwQZAQWuIwmIJKXHggHvsSDr/0VuFWaN7eaKyo
0EzYBAqurKO7XbdmIhZUwJGeYYUZ3kCTRYiBonMxitH4A0B6F67eEOdy1EcqS7W4
NUqDurBNAFLLEaK7xrMzMzTYKIhxZK1AIOrc2Ngt+h7VH1acqQ4Qijv75WW3kCWB
mZwE/ErR7gHmrJ4rjRMCUND6b/zQuqhIP28W1X5GTJY2Is+e9UbVhReCFvy3NVD7
CcgGarJAVOrXsftY7i+1mZitOhG1QB0Dn//cIZlFL34XdnHjBGMeq32WawQkEB25
T5ycBQUoY+c1Zl20NaJ8NuGGnBYS7SiZK+OJlM7ZSz0LWb3JtScD9ZPi+2oWXMrA
tmzwWkyRcJVaIlvwj9+Riv7fhv0z0riZLxMr0TDIKexliKyZiDrQbVb0RPKclPxg
9NBAckLBS/3GwCHjKIJhk7D5fKhX3o1T9lDZS7+0t2llgIpeOwMP+0PZ3ipmIzPX
OPCXW8vvGnVCb1wGKCjf1KEHwRM4UVMvPEArRzHhRDDR9h4oRDOtz1y+z8dFPQ3C
9EPxekOoxyrnRvbVDt9pomkPhWXKdR3MeZLcknQJjifKUWOHc6yJxabxv2VJMOSe
ZzY4Epgs4jICVX6KRG11eFiY/bxsYPMgvuYIKwhutg/hRAlXY7JYwTFa00CE5LgD
yqw853TUkOmOCBf3G3sHG1Qq0a0icu4R36Ojyl8rJYr8lCIVLy27b3eUsL/ZKknx
qssKRTRW80Pw+PN5BKP6wX7FvSquS8n/gjSmkA3Sq9RGjyPIX50VxymM8+Iy1Jh0
bODqN3B2uhUMlKWnvymRRvnYntwN+cNy4RQdNBontcr6glCa0iZX/28C0oCTzIk9
TJMdsNrESuA+2l4T7Xzs8Ac4i4qoQWu1NpaotNO3S/QUhy68/NLiv0DtEUcTH4Pr
MFMncM9w38G7KNdz63VhSTCQW07guWW2DuhkGe5iSMd83F48ZQVChIBHuFJ75pTS
fw7ppRBqH/V8e2cAMu+Trqvfyfu6vYuYIFEmGZr7rX9kvn2494hWHdXvGNuYtyHf
rmts05uAWuKnVO02OUgu8OxGMZZK7okVt8LMwm8sykZjGzDda7ozJQreL6XFgIuW
y6Uv3eZkUf2TvEVPi7SfsY+51pAmbJ38fsMKpj2N0zeU5YmG+7TFN/CoOnnZ8CqL
YiUrsX0+NDjcFKO5RGU1NlBtQBtCN7hAJymGXu3Yn8nG0k00/kX+zyVt7SQRoa8s
hLewMgancO1etVlaaz3eQrBg9+nUK19fpy5rz+vpaHXBNCBOMDM+VbtWtsFFpzEe
J463CiRTgBQIGqyW7JsGqngB6B5zZ2yi7y0vL2qseNIh1yqPz2zAl8D2xCvl9LpM
hUot2Mi86LbCT7eXq8pIIfhll3g4AewFpTfzD96daYlNkjgey9Rt6/WT0ily8lXu
wlIXctqwTNXf5790szsQU8Ji2Md82Vdk1i/oofJRFKoMypBjBBKfVcOk13ub43ZX
0t2OEgrHKMcvWFtoomtrCR4Wkw5TzzBYY284xuJH/oS9OHTp/+fRwK4vPcDp8Pss
uBiP8TCqzbRkaFIHM5o4gXdZD02lhfsAvK3mjynulodIgTF3FypvYKhsRPjeQ/ye
CKR6BaCwmxzVsmNOx09BH8auX4RTga2lo5ClQnnxh2qnfd3Ho8Snj4eXKhVpMiq+
Ez44nYlp0WBJ7GHAeFTAiGVkeC8AHhV6KZTncmPK56fyrShdk7Ef2qWqYOnLyxM6
AjM7Ytr4snFmDmsO7Gu062nVZ3Z7b/6vaC5QILCTqWokDTpcGtVSOdzHa+WnGAVM
Gy3rGsse9281VlDqVQjuLmVYM3SF3rBSviWbZ0JDiv56xRmnaGxGWmucUVKlC6c2
k1J/w2cXtY7GbgaoEY1NIKpGEUjQyBjB42KnlYPopPSnq21Gs/E8P6ocjtQQJTTC
9TDlfwj6+vpbcdVmuGNtCqZPnGZDpuKKR5Z9Dlb355hvLK0R1PbwT6Hb+n5JnMMh
mTMjaCvOD5D7VE+TedjELbCy+TUpMkinubQZF086SEy1gU1kheoanA0zg+eWhWr4
wpi3+22oAPoupxtvbtGn/E9fBzCo9hDNkoAQ/lnG2yHvuZg6EzeiovsFPA2wP1M9
QCUZvC+A4gfpx9Tdc/Jz27GgEUE7I7xQQ0UpCTgihroK4kQtbTHPnj4HEfg80N0s
yaLbWKWRixjJuSa+a8NEronF2zUkZwt4fdAJsnqsGTVALkNP5omFxb78r0E5xv3j
WdSHkRWFhI5VBnwAQqDb1HsVXpdVbTK/btkgAHvQPmLRhg62GAP7PbOd7VySZemY
7ZmzNWtf5eg6hT8zxKeu7EboCv7d/zfRLJ9LbT6Qf8MFnuCNA6HwTS37q9tQx8cu
uw66roeHclNlpnxIcoj4oyizIG0hnqVdZNq/Scee69MnmGEOaXXzYueueiXxUZ8E
zWAJQ9mxIIeLv3Je0VF+/topNH92+STZlOCQSphI62/nyvhfJC699X2JqrwQJ/qi
fbl+7rUU4hOR5sstVuUVnWOCz/vGWhiV8ffaJKiLZ05cs+NG0vIrIW9Wy2tEKkqW
rT4gmCL2cz9nLGQ1OOfPNtSpb85cI2PMZvAMj5wRcob7QqBXbLFtVZzXK1ieitTU
Bbz9qQubM5mRMUfAD7Xjw/YOrhI+SpcS7YwzLz1eVbpC06O9KmT5LlbrawoGhMrM
Q3fYo8NWPP7wkL8SeT8PD1Hpy60AAzD7t7rL2+La1/nVtO9bPmBRWzjHH9FjdriG
iRabKt7jApNwa5WSq6QsTr5r4mqrFkp54mWGZlnpqPOOR0NwlinkzwKPAw8flsA0
3Q3R22yjUullNa52sfssfv6F1+l6VcE4sEL+wY96U/cXOPvUM+AtAeupoE9k9a3f
xhv7PJxv/jmYOsszlAn2g3g4WyG90qL9e9GR/d6zzUPRZ22zE73k17HPR8xT1Ono
TRX+zCzas3X8ymP6T7V/t/R4up43X1Xlq7kJi2Rp/0w5y2rBoaWpHLCnNzX/Hk7s
b1jD+boz6GLblHmRfIgL2EPbvwhkMSitYEyhGOMnBJtDLMmL281hfn3GL6GMY5yW
Cn7QecVY7AGr/5grelOCuufD9ikS9s6kABKna/1w0LGk2dghIE6sGBwi8ewMK0Kf
EP+nsqO6a5eYehF9OGc2AyCchqiy9DcPMZCx4tebe8H7JioiWOWM7Nb/Z0lfAVMJ
5njdtyqTCu3BFws6qpek/7ZJIeTxtIqqY7fr8CfHUKQpi1+MAV+Mi3BAnIXY0epp
JWZjImm4kti9IHjveaxSg9c8av110jI3WQo4Hx2mX5K/iBcyNECv6M/x3bWOr3gy
5BVxrOZuRl280YJ9LAKhkVOcp8j1AtHf2iIGlUsgqcR3za4t8uRaTMWrrSmm0Hmn
ea0+J4q+0UBrXu4GID5ZF/h9nVCTbmD+YrDUgpOWNAJ0McNaNUojKTt4p4fNyXrf
YWrIsug2JeG2qu26/62ivm//S3rpfk2cW9dBPgrbsoPMgujCWt4Jaxub9dMEZUR1
/775gjjoWpQiDEfhYBdmNvjbMIzMng45SMIhqueUaLaJ2/EaLnUFj03WcKjbWdaf
/pXjaSvNdWXD4UvvJFVczKF8eefWJRWqdq/ruU2FWahyKjM8zzEim4ijeYlJ9clj
5gKNFN5kUFliDsTHrOtwBJ6d6sP10bRrCD3Wx6wyhHeOB5YhO1eeDrX5rVD5NZSy
spnWSkEuewrrp8L7Zjswwh+qzbbYv3A7w53f3Y5/VbReTFPfrV96ZHybbnjmhbZj
0u6bi0nag7JwILLPoVImexklJc2OvSJrwgZVkjI5LWxvOBeMNuQ/rvVKT7i2KFjo
rK8McpSEWSd7AuT9zE8guuu8BOiizJt8CZP1G8Jkxhe+yi4nw8gzZqiweF+XonaM
K4xHt838JCBtlA8NTdXNc4efrZjtRIaF9+GVd01m555ZPMTIHs6QwzaRvgZ3EUV6
KauD/xwBx13cYvcgcRsp/mCOD8CuYteBzBYPNZpM/62ul8m+aSoVSIjN57YU42BW
HWN5E1fbpWOZE82TtGeo7ll3r0cmFj9MCb4K6quHw3s9oLH0IBgv4zm+N1PLeGGV
YsZgz4EiHyN+oEGoHy04Ph3C+QmiyqbHhF/wWf4kby60zyMUSfzLG23fazAzXdXP
BT/K8TnkwLYloZRfnZ6aVB0JPTjWgp2Oz+LoJJFDNLOr3eCgW8fk1gBfrPVp4TRR
E/4JCXQuG1OO4j1jtG+dbn1esMdjLY/fc3SSGyXpNaPYdR0BCWJQVXfl1mj6y7Vu
7YfnEluPFQQdQY5Bm42k0VMj/SADgGXS4y+QII92qATrCFtxPxBrUS/hBJ2uujQF
BC5edEaypnjnsmKGdgjNSfNOiXBz6KmVcGueuQza2QMU/g6JoCg9zhWriGAj9VKm
9VlGqALrqBtbJ4qyorbFCzxurCPB++Tqz31i+tL5HuFpib2vpQf62nklZNi66H8o
kU6LoPVlLHnORPuUTZwUucApI3U/0fXvcIsFsAj3XBNzTXWD9IAgSGquTLcDz9W8
PEZCX9VR8F4/RwRneoWeThD7NuOIoS3QQi8ArVzq0QnVMhtc3JEcMg3w81YgbJFq
jIIfHTIXWw8EgjC5KzrkH+fP3aZJw8AfP0ljizmnAXGDfgqSpMNxAMaBh/S4qwKD
SsfE0IBsDycNafOQyY7vU5brGL5aEnNVroQarDP9WN7OEWS+9qVKhIpR0BZ3cZBF
WiQ3df9SnM9a4kymY5t7rzT0wJI5w/JCX8FfjyLPo9PV7q/dky2RrNaVMD4XD/tV
BTTkEiFbEr9m3vU2sXxSsc0/tepEntroZA8t6hyNCVaO7EXQMLr/LlslM/bplO1D
zBo/bhvXCBp4ncjH1qvj9N1rCrPcu3jhGj2yBWGePmK3r0irLr/dYeQ/9FS3MJ3S
e+VKHBhmgaQ+gRRTOoLz8P+mS59fWn6C3Z98z/+qKOvE2IpAqvmaSnOFkbQn/Ege
Gu6ZMYyktFGMVDvbKKpc/kwrIpqPAN072g0LUdDSGNGsaHJyrM1vyEAl6w4IeQkb
lrndxRwVqrWumNK8xtZXnYxx0kv/zlLg2SDBm7nn01XdSJhpt8zp6XuokgZDwq+X
She/GNZu9zD///yPxXb+7/7dJanNmwtfpBAZlD+UYxhNu+FGmOjHSHHnz4ssbext
qmcEbewfx7anBYfsAyhsKM+P7/oVFb5/dLdoo30gpZ7CQztxZK1SCb7wYiyclUVy
NiO+uh1TJx3Tfe6W2V8OIaSCBpw0g6yHp0VMMV96D1tvX8P/awtwrizUWNm/9zcm
O1vGunxgZlmLbYvqP2RHG72Z1IJilQ6undVo5qYnT94Okm/cOkpogznZ1Pn8DLCz
tM6QWgGTVLK6nUdYCJ1nt0nBfWQwZn2m1OCv9JDg3LM5VFqgyAMtiY8mu4XAkl4l
9ehrsBx1H+uq8tyLQ65cVsK+qrOu83Ti0J2TAYCTr3PSEkzYBAnAXDJOCg6cVdgd
T4DqhH7SAOLpQp81HLKqE8C79iqNyPPDjAZKBzAo5Z8P4uHd9HRJRxS0BGud+ZcF
6+FPJJKrD7rAKRwrAOAeTYQT14XgdQJnjJlgbXHw8m4FfqEZggyzE2WsVG2ooS3e
XgHx3ap4e93l/GzlqPifse1c3b9jnaEhU+vy+Dn2R7mCc7b/uD70NzH7VaXOrtXX
HcLTOumD2KWYXM+J1PboEjKV/Ix0WYWkuA4EFpDQddvQlZVi90uTgsis99i8SwNZ
N7Oex3s70N2SGT/qYJSXb6Zl968gry4M/CCPEUMmFpgySYMW0mgCst/9fwAdWk4G
kOLnlHgA36RJr9wezE1/AMnBefPfSZn2r+mVBBrUNU8vLnM0n712JwSSASQZnbTE
eo4TRWwVx22JGrxRvMoQLguzDit7V0WXTGAJdcsB2D7oDQm0pWOjN6MvZwN2u14s
4WH5erdzp4v35Va2IszVn09ys7BKBqcBltE6WOrUsWAbvSIyrxJyzCYMjB6hFPxt
tuqqhGWnhO34j60rjt0Zoy9nbYjjDlkZPVyeJopigfbYN1ouWCbaxW3Xk2uTVh7z
zIMfNwJ7yl9eC1OoWHytPptvFzQevimDduGbBurRM2ot3kFAPvwimHujGIj0u41u
ehXQtn17PIyK1Les21IIk0AghadfYFHhTEb6XuWA50zOUp3hBLImkoXy3inKIR3s
7VSZchSQll/HcJjjGxBcOPopPPooYMmNW7hAEVFasbHXlTCzSqO6ajo/AFR18ryP
PfzgiTuM6wxr/BOt/bTPijKahPVRsxV8y9R72XY5UoptUkCSv4LDT+t/3cL1yjMD
Pfxpyslybo9I2EvXcYtuoKQCjijf3uzRH56FKnxNfnWNfNmidsMaSeHxu/la/hrE
a3q7Y50L1k8kFhQtpL1CSOrJxAeop/W8EIpw4J2vRRWyBVEIfI17y/P+fD+I6f/C
MCLrdHd9JBuNw4fbfR3ozwN/EpDN+hXE4IEtcT8qzoDj7X+l4ZbkJL2hguhJlY6R
AAgF3DcGuYRRU1xRX0pFjSkAAKvQXAFQyT/8xyou3qxw4QobMWVdJoEldOmEdC5o
KNa9lg5E2HaapwnCrcqkMt7aF+sK5mZRyPNKYmTu1+fGLJTOzshUoaCvgDaFNG/G
nMdi9qD48Lat9+abYSKEpOlKfsA+1uLoP49fgFQZg5uNuWQ90D/vkoJ2rvLED/BI
8fmOHzzORjJRhGik6Sf2jKWhRT9P7/dyvZftMgSMtuTD0Ckum8NwnopYY59IjbP+
Ep2fwUJAUgpreU+Z6ETut0OwAi4x+VRUPB/T0NKVZuw9uaOzERG1saWYgEfLVwKG
94l8ASpKR8b8RGxYHYsVp9sWKOgZqABvn1CxSJSZg30Fltvz6IdYEkkHzMwhB9F4
s6UB4Pr1Y4SubLup0zDlvWn+TTJEUUt5J8dh+TY6f3GA7881+2LkVi32Qazkcntq
LrgNpXKEZ1LKXcNtOQGGFNjrgdLz2jH5ck14ADMvQDWiVNb45Vn0RFh2pXD885b+
kt06NVI44AhqrOUqTNRvHgufDAStVzpfhqgVQZoXYef72j5ov9SdasCJD14QNvPV
mhvxuaWyrSNstRvseeD7PU0ejEW6e9JXXHqQZsNpW+StGCRBUh7E5cx1NKFK8YPe
rdIEqhbmuQJp3b+zVDe1u+SCHij/kZ+8j6VUb/m7JSK67PEllHYJDszpB5SlX2R+
yY5DomCmBVRy4Y6cQh05p/MWRJxDtQBdhLQr72RCsXF7es4fEyxwn0bPlVslJvfY
2UNTPymCaj5OsbVSD29ae8EGKu3g8OptTT5k7gYHTQvqMqQge7qpi56uPTdhzcid
8OLQ5Y89wVRK0RBclhAmqpe4SPfmCf+uq+92gednQ2gvo0XHupw5nHcM/cr2gj0P
+jhx8TZ4+2aoIIsFrBdZXS/mp3IpUyc9oE2xfRwAAt36PIyvFimcCNCzNxXZKcJF
Z/TqXz6xFyHhl0C88VaFywX4bRukMhe+V/RUqZpKtsjmApP5wU7uAzcszLjkVHZm
37CXYbQq4T9WfHwgnxQ1DVjc0squ2jYr6sNP1NMSpVeJz/8yv3fVxKLVVpR7n8Sj
gdQOGUQ3Jlb44hwk+P42gb/dITumNNt0zO6ggjW67nW+0yjNZ+l7qDOEswfePow2
ZyS6TLwmbkrEvd01etm+zK9pa6zPEll1bKtUVQD3RgboYqu02hg4W3Bq3s3iGqC1
4lrdzU8xIpRxMxAa4i4kLVAMwW6jGNqM87+FC8nOYMnABvmZpzS5n5kE9vUcPubj
TKPX9LtQW2SaSlxvifumGkFHYmQQ6ULa/fVfK2MA5sA4XgylDRa/CQDn6Wi7jmjZ
JZc1Rf06DmJW87G15T5P/M1OnfO3BH/PRC6KdYbwHJtg+a/ihXJj9aojlSkdGdT2
r959JueEh8JG7BI9AkWOZ9h6qYZ6lfDmGlpZjDgn71+df0dVUUFSAJXwvUVjoYdA
mmM/C+3Cu+QfiXuE14IEv7PGASbrfTbYtP2YNpGoyg0lhFy5hEMX8MaM8LpkUoEU
YAqSgCpzB2ruJIczUsq1WJt9ySGYmPAolI1wM8yLVrmTaM22UrIZpL2SOfX2Qkdl
mrOU0iwdb7aUmhRRdZKNb29k4eaCo12ctM6aYylIAbRSAnqOl5mpMt4JT6uK45XD
f4dHJ3xmkclwALsFnr3NJl0bIHHLGp87ywzhGiaRRLrJ2F/NBMou97LMaGtZGqqa
EeXf6zpbBLS5giw5zdXAk6BtxUQ/LRpWjEBnpsffbe5t9WgOAA3u3dy9d5vRDcn/
b6Ai+OzOM4k2v1LYRlD8w3eEYo70nEXggWpH9Hq36b9PtpOZaskdrEJS7keqRQU7
GZXr9W267a0i05b5CJ6+Gm/zLqMfVax48rePl16f+nkoFBSWkseOBECUesAC/vIt
JMUphp0roIMppIU9EE/LTkhSbjwWlesuwR4eD3lOqOVjwcnfEqGiX0NiFrkBc0G0
Gg7s26k/uXzXEdhAu/9UYDBOWQJzbQtNOMygKh5Ni3FdSTL5JDTevGarXi+/f7l8
c3Mcg4ptBRZxSbVuPT+q798L0pbEiJCR3iDkpQdb8zDux6DgM6YuBzQoXZYIt0TZ
c97gSmaaoKe1dHZpLuD6nAokyyeGYFlFWu7EXnd8WMSEJ5Fn1fA8Ex0k6CwjM1kp
g3lazcy6xwg64Z3dmgZYDPzPCVpLIL/nnACW++97Vbyl3gREezLqnaOvJmf2CMDn
oSepQURns+2i4sOycP/r856ux71zQcODtxW9VJDztjSI3D5QyUDOz/PodciMkrT+
FxpRRSEJOQLY+DZUG8jdnguyCU3Z6oKQYxWCr6HLqy5rhWTB6rRFKeT9sN5j9Trc
TRzf3cYFQbUit6lfhVtjGXlAjJ858oDffWsdy/okTxIicW7ObCIJ4iNH4uwE8G1u
T9XptYh51JkBewspjl3LXBdL3Jn0nywo242KrFw6ZfMhBTQKQ4CmgCepLUX5H0Xp
zRvhOAhmNFqzkfqqIfHhGOIv/FtQE//B34BojGOBwOWhxfdjKZYc7xWHZRzIgKMd
QjNXKDq8zPRzon8/KDIpGe6V8awird9qx83s3o7NhLX3sPyRPQ3HV1gX7wk8vfGL
CPh31aQNjqeFVEiQSLIClVMTHBH/RjKpO0goZ6h2bnZKZuFnMYSWyXIhOef+gOA/
R2pg5gJVN61EhaeFOB/hgwcsQUXNvznp0I79soWLAHSfdIrPfatQyrC/94CUo0LQ
nGnFFRqGFge40tAfrXl4FV5nDRH4qoH4WjRKQQh0kJjYCG152ns7xb7U48W+yb0N
p/VuSmqGbY7jYSXULeDgzrIe/IlxW7aKzP01h715MLOYCVqjjR0iunXQ7GcX3mAi
Q07Sd2NybMESeqvaD9T0NDD6C3mn+5g9tSNQuSKWyfzL1qf7j5Z7QOdj3nzTDY6Y
jweLPdO47C2kcu2N2GnXzz/yKrwqxt1G6ZN1X3zgLLQoQF64I0wfPbLaLhWZWsmK
13Z0owwGxEp7Fxu/MQCK4rB8zd3GScfr232t56m7owLH69rOePb6hTwSSSnMbpZl
MKL1ypZ8GV+2C7AzpPObdKg8DFna+TFUaARCtXu7RjiMmDUa3VPzRYcHe7cyG5Hc
4aBQjaeD0f9FfhiqL37rL+jaIOxsZBwSsXub91Icm+GzyBjzULHkysU6Virdozuw
zSX2ubzi3Vj1sH01iyLZ69FcsIbHeCwZgKN9ct4rgtJ+gxe/FC0q1Ow8RLuxMVBk
JgwPL7+1Tk9t6ilUqZIvZdIkhrHCyQ13nf3eYslhOGP6njxBFqsd8eZuZ3TkQKrh
vrG/9LcOyv4MOnXASeupgM2e/dqChR5Uh4B6c1hduWTwD/Swju5DFewESKbZe2Q4
Z4aMz+auZyl+cs1TS4saUWSpS6ecMFIa9Pto+JywRI/3gZ2tDTq24RHblT67BK1C
Y4mXKdKOMklZw2WfiQ8DO5Ome+V1F/F4MvO0hiTre3XTXqm8xr67IQsxqDsxjnYs
ItBNC+6NrZ4FuBrJC2+ddrDcaLemv1IxU1vCs+87u95/02xPSPXMbMfiFcxt/fqU
PwpM6WXiLCDUp/xeqx4PlJ62DnzxZxg4cbD70/8uxYkRdYPgz26fNN9dRMd2cLpG
AqadkxpMxkIYoyIS0f8Lrg1EgupmDPaj2Ycew/PBrrmD8++2IPuDczY2hGmkWw/u
2/cMgc4LIgzWiw1W8r6+N0l/Q7Gddvy43l/rJHp2EWi1k+hXQ5iXTandw6CAH142
k2h1+NvwjMlbltc5IuhSPjsUejbMV6rfRNB8K4o9xdVpnwQuj2sBSW8IF2QZ55gW
EXZOOUk1fK//GYQ8sP8T0ZU2yXyfl8mDO5ffcEAIi2WrABefqQwyz9EGpuh4E2UB
v5MCB8BjqJz5YGF4P7Jr9VBvg35FOWFlgfd+o0nrQIkPiHSCBvC6ZG+SRj3oewR5
/ZqkKhCmFZdbROsD8wd5xQFTq5A+EYMIdkHS4q4biLRO4zBekNdLq2uEF3VLngop
r4TF/fWeNiKavtJRd3f+bLCMpIA3dY8fJc/gSOdf2G3hIVJU9xwQG9bj2X97y60p
8hS+QD/cCZQmjstlPS12YJ9/rCHDRQIV/vySAsGJpTCvWkQasv29OsXWrtakfO8l
vMTEm2eDKgtSogJCN6xwGA3+yEf/xAIwBOlRiFB+oOKDhi4hYoVeBboBCsVfEsAm
3hcVgCchzEUpgDZ3EFOPRu8a5gHzoYjaW54ZZHUlEJVrNDt2R9PQwpb7Djn0cgBl
EdXSiXxc/mrxYk/faog2RnB/Sm0Zpq7oLqclzuzgqSBZ+I9kCW1hsz1eCJmu86II
99TXLzg8NZd4FRrU0iqSS2Q9kGDu+kY7essrb+MwclFspDJ3S+0aLUSkTGFkYDE/
G6y1S0bnMiLSIIlVjFoTvdmDs4x1sFmJ6n8lVAoOJypN2un2VoZz+AUYg00iGGC0
mq3HnQ24cQRGgEsu33KVFbOHiJNLKV0hDMQVj1J2U/qBS3Pkwo9VKxnU9wLyxgPN
W9ZeWg2K9ICNvtJWiuTrhOrYoujWCCXmBXfo3ZOc5e8O9RMkT9tVSpm+in0PAy2u
imNIzWosPvQkHVZSTSOGgewhFlEARly1cp1EE8t4PWk/fbWLwt1W2CHXRQDFMWMi
0xVdRcu08PxPW4mq2HKLw/nGQSIKJYzEkAuFdbaHN+hhMhnIqU7+m4Nb1y1WSVSN
03x9CsMyZrkDoN9IF7axyJLBPnQ0nXVI4U9uumk8XfdHexnlhoj1Ic2uQb58YvG4
eY+jv8esMPkI+AO81I2TZjKdY1KCMWpRleZNglj/wKgNJI6wlqd/mjJIGnQrdeFS
yFzHkzfYmgxwON3umTFjFl516jhTr/VRZmYEQkNiIgsiKIzcql5xKDRBh1ySKjs5
nPCebJT6adlgU9NWBZrfU1lKBWHRQwjTjkN2gCSmzcWXqVLPJrG/yqVM6ufH69YJ
Ca3X4r3ShxqhT2yAVD2Mau1ZsOOhHN9u/zgOJb2+9V7gVNu3iQHtDuMjorwROwXi
ykynJHzhdzymyEiNp/Nupfnf7mlSkLYiPZqWUQyNRV4xMBCI/NROHsDsXel92Nb+
5tGX+m4P5pcnY9Wd2KTXNiuReG8pyNl2g9c025FNfjbFPqC/coN+3TZtY0Dr6Q+Z
dtJVDsTw45EpkdTqbaYH6iFMyrp1SAXxP9D3IuR0LxSswTrwE77xanXGD+h6JzNk
Aid/8s9Rmh8FGeQvRpuyx+9lHJbrA6al7mjN1HaWq8wXeg5fOMBPSv5C4BJCah/k
hgIyrU1SRSSfsJ+AeHZmCJ4kQStwO68OGtAaVXJSeFZNjGwfwDvLHTq3esgK+dLY
6WIiI+9XScMp5whOY1IbGSSRUmVJSVYrAC3MNoqaEvRtU3lGsC6eXxEHd1mB9euX
1BkkxsuoZx1m8854YyqRCx/uFrbfwXAG8ts0jvMriELYXLG4qT1DLFe47kdn8oOj
NVlZvUJpA3xfde6hsfJdmj88I5vOXOmljQ2dFgwqJ68LBeQhO0ywJYLmfGvdwBRB
na1GvW00dMHajkWv1PPxlL9LW5vxMV+AYF806KZD+r2stRD+xXTYlecGwt48Qv8L
sE6WDYDMOWBc7RvZ+fuj+0PhL/3QfpMyYte5/9q11f43TCX5oB2uF7kEY7+JiMU8
fbDp3Vrs6gsVD3pOv9gWBPJGqW/kVxAScwh1RB1GoaD1sns1yZi5C25YKuxmyASC
dSMZDMF+ka1NVRfEk8cMHkHr0xbjb3lj8e9sW1Pif9iVFrvJoIdvFnQrLGD3WzeA
hk3SPlF/T1o/O6AmWMzm4PCZllbR57Hb0Xp7n6h2/AM8+Ve8HYI5yT5Kz+L4KfQv
/hwacC532oBxliHtjri9YrSICNWpNs06GSMjGEJenFpE0MU5iv1FGJYzrEFxurna
hb/T3Zqn5pUFgwkJ7n1SSQVoF5RnBk9OxijSEljyWeOaZ9Hhc5JrFxp66gZSt1ta
7HLEQ8HEPK89zirUHmtTCkXDNsjKd3QDFyh4lZAQNl1L0GpGCfxb214u98g27lcv
rnH+yhQAx4iMGLbPaDX7mOVq048y7rULZcvUs3rNIh5H3L+cEpbdc1mddG22Asn7
cxf2Incw8FAMAPe5daHMWKLQ9xlifPRV9mkxpAuJ1MACWme/KAimraQD8CS9RveM
QYmwVOdQgA86RsjQlAwhAlNG/dopg5ViGlIW4RCh+3EoTKGGLlyocU+fO9lg767c
J+MBbE6jPv58aHcKWf3ZnpXJJPaeGqQy4Der/VXMBJKn2/XUBln3cDqvE2J7Dgow
UIdTPFVK6yL3sl3Gvl4uackyW+Xq15r+vB1uEYrgptkcqDajV0ysVAmiRnvUHqN6
h0FYtZZzMscZx5GoNpYyuToa7TeoFyxI8g7elZNZD4h/94cnFhoqWIuFOV3dI3TV
LvnnpGx/uZpMhmXPUoyYk1UJc6A+01jQTEb2PqIpF3Zg6lXguHc6/aP9O23dePf/
fQDfFL7uabmRLTiRXDlHhu4pnyD8WVd0IVjrFFYD5+EfMoMjdMIqvNiIhhTMSgc1
BINB36yrAkdte44/DTGRQvui/gWssxHgkSx0mFu5f6TZRI1TP/9oQBu+/ZV5tzqK
+gkRrzmxF6B/zYff0b4ueKJF9XfaXns1Y1R+SXZV85E2WbgGHVl6S1f/hSsQq8J0
p+KIdOEds6GynVuYIYcwAsmfcoqa+1wSMjRiI+14hXwA5HNRIba6ws/WG9e998WK
ky+sL1ooB5fKMqlj0vJAEwDeTP8LLGF/XUJgbuJDmrYmetd84vmxLGOdhtLbrQ7I
wTuso/w1XHz/XGxl0pooPVCnDWeTgqFaS/ymXhfqIY3/DrFBLf/5KJWqjRpzv/Pv
KX9KKhloRN+WIouEiNQWLlSQpMf9G/yVvQZde2pRSmd5fCwhdci04v+jgAw/Tamm
0XImM/BFqkUaY7XTGdzlNmR8kqfW+755us+gEPEvXcwrCwNjlT7IO9PNjAM+8/m5
y8c57VPLVel66C84va0BYUAVCnn++0uyr26ZWt85tTbw1pA+KOZPo5AioFPsWoso
C//4WMFu6X/en0j2T/34+6kc+mXLbV/gMpKcg4BNgVvdg5UsoH2W+wDgTqSexz3z
2kJhJXKZJuW/Nth+pRI9GX/8KOLhjx0122KhwMj6IlLlGkQwvpV8NbU+KOxLBCLG
BRaiuxHeYLBR7mvfaCcBMgGgm6mVOfsAToCik6Vxfj3p2pJlAINoma4I1ikBgTLQ
hQplkGPhClcQ4oZjmAZ/ygBMUbhH0HE5bIu30dadUx3W7as3u0fs1aGWhRudmTcG
f4dANFPAFzgn8+VeEAPVT7d3C5bBqcRQPH6S7YOyzToGAHOHTVNlYPvnJoOIRGjx
bRtz4j86NiUBxlT4aGz7e/FJlleFDtiNE/i3mKRUzN1PL0y+tY0/pp3cFyKrb5Ro
W8wSqMpG0jQyhisRGu3DWHjEZkeNrIApifTIDCENbpIJLKsUJvR2fsI762YZT0QA
Wz3Q1jHdI+GvBnAiEX/SqzQ1baZC0rb6YZucN5JRxzV1WaF/67S0K0xiXotR8jD6
Cn27DxS3BgiGe73BJAUuxg17hREySaz6Rtv8APQlwdZ7BK6zqxD3kriFtYNFh3zz
cgpocM1ImoQTPG3CUqwNOtGWVk1Qjh0/q6J0et1nGmSX7OrKidJ3TM5kAkjOGs1o
w0IJEc4fjo8qJARm/NjKLG3YFTxblNh92wBnmDXOMe5yOT7U0vvE3gMuuLt1ptZQ
58F4NiQ1sYtdDyL1di0jfNPPBjRMJgYtoSv7bSFPFoE5nV83SS+N4MqPAn9meDJX
U4PVBZjHsk2jlu/iTI4iC0IYZnEDBPwPok2BFkeh5DWbrDcB0yFadob4eEc2s8+f
wtUOfNX8N//l8KoHTWHzTVqBuc5gzz2/r8gkmczwFqwAR9oz+zW1ZTH9B8nUijId
lhy1kjrkelZXxyh/RgKGNV6A1Y6QyFh6a8PDPJgesDMgADjzJh9PXRW6fGIZYjyo
wZTG0TZUHuhaUNdenEi+WP3405cWH8rONC+YlxGcKwVRPdMDVY1EdKAuOd/WcSNX
N2DhU7ZrdUUHEFuGWUFajgqWf7Jv9WiZdq/G+v3J+DT2OEk0rXvKS9Gvcj2KrJtK
kSn50AK4JZKwv+SuyZ4GYhG/ompaEI+wizIEfQSqvJY/WyyvGw3PTCTFv41/FLnl
MChMDdzRPfoH0gd09lKmyQHSaU6J+DGLgm24VN6RfaiagvoftXODlbUHlQifQPnj
NVwbX/UzdfyzrzdnoyQ7K2zrq5sneMMbuxZmflDdsb84Mrnz+ccNnI/4BNsM3rPf
juFCnUk7m4N6AOl8UgT+naul4mit+RObmjzrexSpP6S/8aoK2L+yNPO1+EcdXs88
yjys4QZ3iSwOKdh2VajjBpTHf9rMEIO0lAirH5Bv3XdL3aWxi1jg3Fc4/5xgJX8W
1gYHeekwL4tQqdVZhi45bI3vDM+n9cD+hHwWTfagwfhMO4PD0uFLCckqGLiEBZpA
8V+Je0GOs+mWc+UzmV51bDbhioKoT2SCYjbOesVYv8X6p27/SaTeM5qZvxle/65C
Zn/n295/2ZH3fjvX2Rty45LOltJd6rVkdXsuBJjtrUJEBNtRjy3lnZY7ZLydQUOZ
QM+DB+mtOqh7Oc8lj3ZOExro4DVjLPPzT5M9VEcte05Xn6GK++JA7kl6Zi8HGoZO
Lkhyk6KEApTeGP8ivSp4aXJzcGyWVjaOLoOO7MifGGeRq7sl7N7WoEnqmrXc+H2j
4sbQPUyfNrDsVCFQ6TJNlJFnKqISXSwB62gb0jMz7T2iFgG4iyu3jyylgPDLuJYN
TKuqpVnmiS2SvfM3MzQ+nT72OSgAGJuyZ/UcgKFqtBLnuYTBZCFE59PslKhRE33W
ySFOLFO4CdeErfv50NTAgBfI52RD3H33F86rEBj0DvjULu8wOdEWEyILiC/8rGMJ
9kjlIuqP1lSFwk1NJKNfHPwkelH7zMzxPGsGp0fsbXpaii5A3wphGuNGvFIH5AdN
780crFFdh4Mn9fMhS7NqrXK9NQxG6jdyJQMDN2YUnbgyX/3s4kRpbJlulCTexAfO
ySRaNMpVTtAPEhPJWEv5GU6gtplKUBCPLSFtuuKNNAu9fjm8hQvLUFrVGUiGDnQF
bWUGOtcyCiXY8wzzC8ie2bRIulFgynpLF1lx6dfzjIPEsQdIviX/a/NQWzKFi6tv
dWhE5hkOuWfdx/5868rhrbTCnDaDxIN3Q7N3B+iOKO91DbgbKGRdJwdfOrQu/KGA
Hdt8bsqtHuDUmpE7rR4tG3HTdd0AGMJDWtTY2sGozLXwIiR2DqkREkJntyOFfM5h
Ow53fvTqbHKKj8F2TbpFmf8MQsHsgo0hKcuKVmpz2NI7T1NhYPi3cLWXHG1O5rbw
F1vXySxM1w4nyWHThl6clE4FN6PozHja4R/a82RUdVMVFBMwiMoGtl3qKuIRiE76
4wYFObrpbtnPcqTuVgyYn6XJgpD0Xu3iUyHTae1Yt82mLA4eo9EQtGau17mR0+Ne
KbURYVMuCPm9qPes0n87y36K5dwHDZCBOtHycmlQKuIR+NBf9Tjzs2O073STLYQj
0S5u9RAic/ScCqiYKCXXSlaIDLecWecGrNrNz/xO9pxp6kxufJaSSTxNlBO0cuNA
m5OC4cgVjVKIyZ1W4UfMQYN/g14f9AVYaRKNWX4Nvz0jmzOvJ/+jMCdPfZJlX4Qi
9XtYKL/ZYbrhPeeyGS9nUxOdWsxFv82PV4Ck5tjOEIdC+mzNlN4+1vB8ceVaT1P/
BBTak6KmiLtrfBgsNbFg29thHqd8W/o7kcnysuqqPlPd727JDEuDIuYAzepTSUGW
zN5WGb1KApB9R4GlsyWi2OUZMij/wAEEpIvdHRa7MM4xomqb02/EEuUGC2A9Odxk
xwyln3/BiF+9ZaX9qi1JNuveeQlUfvaLuTdqqEPq8ZPrx5G/587fgHW273rxYMTS
7AiVllHz8KWoR6GNdDNVCu3d3WYcExI8BVfloipGkNqKQbJJG8AGNONty40+ix2v
nOpmxXUnYcx6MrLZighIm+V/s7AIxoNm+Se/iZ31O8c72Y9JTHmwdpMWCQQ3k4+h
XDW8EqZypl+ZFyyBlakNB1lL9wNkQa8Y5B0WV1sLCq7ZOM7vD3QbqnbJUULrUdOC
jt5bQ0Vdgz8W+7paNNjvCQwuthKuX4yAhF4sO/ZpxMykGdh8RKjPkHhlFJQaKEn5
4FKF9ow8GywxiqN/rnMzUJuxrv04NuMUtxUScb51jcjO94j8cXd71nNY2oioKP7+
4JnyqGujVwYl9yhoL1YMBNP5C0yghO68K9VhhQPFjOQgv6SJlaGgFSVnOjflPHZw
tg+oVPdsGzv+lAn1X50ZZ/POeXNVIy6ff2zToa8/6DcJ0/di9ZTSGOTj/hcIjPPk
6MLfWj4kvw72xFehB3rsUAlOXwW0VmDhr0UiCtllIzYjOsdh6A3wAS1bUsnC3dLQ
V/CIib2it2TnPd0m9enLJdw20Qq1c9T68s1Sf2UF8IaZXEYZH21AH2P898ci/IYo
UqHh/nv+MyEeX5/fvUzaQ9jKZlljsMaTOh65vnsuq10u18ECB0lF3NSlYBe3kpRs
dlOABhpAK8FUO44FMabvgImyJx76MyRXtFagijrqkePFaKcGt/1WD8vfRrljurEw
8ephC4v28I+1KlIt4dtF+u3PjB9EM1Iziu6879a726TwAJMb2y2ujp1S1+K60zUn
6VIf038G8NvUiGApFh3cAAD5PV92JOKEQOW3aj5TLltCxslPDZ/nGrN+hEkG7h0W
69wdkxvZ4LiPQwovYpkN2nNu1QhyOF/kGb7Y3VEFbIhzkWYOaXhgujrlO/kkqXhJ
GPdJfsdx56M+jY8Uvuy2BkgLDfV1nwrJZFe7eNZjPLSVorej4an/r51NwMY/d/bf
2HVQmBk2tWYNnlxizPiJ+YWM+LnMLr3u/hTkypUftAcn14hf8/vgPkxNfd0E85UB
35BLlm6hWMFI7ZarfMgZ89sq+unQLU28xsce4eGgHfLlYRgKoXGp0yl0Qmc1KHnk
gXHH4dHtIPr/U0MrHKWlnPAPL1Q0sBwcTy6sNL8k6zUgBXdnIBzvb1f8SXA9Iur6
8abJsbVZjJMe9dwidYLbPGwzHIvOzvKzNlN7RCYC5+A6FLdNTttU+OjfLmqhRPaX
P9bGn334lAY+ZiYi1JI1CZ/ZG0SdXYy3FUiF38Sn/2YBRAWKmwo/N1DYH52RoYrF
WhcWPXWvWpQtpEqX45kGi1Thsh1FjwFPiPx9+Troq8c3oGH3HKg1JfHY/mPoqytb
B4k0OU/YVqoiqddwi1W5b7UxlyBmB0DNprZqPxbiuoy/eLL5EoqrUhD0Ltaco6f9
WBNW73eYomJAViUfmioxNYmXEShWbnvM1VLAgLgIQmjm3DBVY8sI0aruuUdon4l0
kDQ4fVKmuTBTPEMaRxYQBX/ZQp/NwPV87j0eO5W2jXErq2KImJWR2OECZGu+hFro
MHXLqLUEe7zE9BT5vIz1Rag4cG8EzJWi5mvhrCKLFVEUg388T0bFsvlmrjhka+1I
DYqhUuiSO1qN6pNq0CiX+67hDKNlREzPpDkFDCeEXMj/dS8h/lqzlzHbcusExjPZ
+xwH027aXM/YDdjQRKgw+1ts9ij7SttUcodpSIqKZVwcXOTQyLvyV5s6RbtJwL2d
bfroMHCZ33/716mkYGVecjAaAdsGIT8Svtn8iizdoGI4rgC4ka5M44oSIfZGsDJV
j9KmeYvttC1vd1ueo/1233BC9T5Nr8oYPQqfl+5mAcbnUar/OF6xBCB1gfc4Zixx
8ysxUL61J0MjydMO5fLsSG3ZelVqM0u5x7Tqt1iA8n8EC5ydXVXxMU0+RcH/8DwD
G3mT05po3FWYYE1QpqfDRQvDAIvtxqIOiB5Rirdwk7aZXgCGg8iAoakKW2D/9JVQ
ItIHlwW3D846+yfVf3S+jqvMWlLjQw6rCc+s4qMaNaFu4y0eGPWjgZFeHUCvSS9Y
Lt2hGjoz8xTE8GtSoKEERxn3ORDyA8FfoQeFBMg0GPOxh4clZXpRoanX/snAHfsw
KxK6XtHc8ps4Crm9qJwHkPJGUk6EX5uLcxFD/bO4+NuLM3a6kEqVT5+gl9vWzONn
bK0/0K2MGP7XtBJm1j1bxNPQBkmRi86y0/9jdCQ4Ymen0G5WmIgdj21hz6Fptt3+
jg8mSAYNFAp1PxWOuBM1pYGghoiPycpK+hk6DoMie4exmd+3qgpisnaDm0EkORZ2
iS7CgvtSR/XGlQe7F7ba5nPDOdbTYjO+VD77d7ovD8vGdKhTwPwG+hOEEX6DBRfe
uLr7GdjfsKg5Nqcmh1vdrms2xwiMbtfQygNIySd9ezTgm1a/VUXe6N3D2T7Fu110
FFgH6acKrO7+jquGK8DtDL4zM/IVkBXT3dwC4mMbqVl0uAhc2SE908KWI65UE2qE
IHuL77Oyehvw7ghf2sOHuLSMO7ANa7zmPO6DIEW6opQxRRLodXBibgn+o/LRBusX
Dw54QYF1WE3DjNTE9ZhSONvhFCqjfJu5y2hqk4kWv83p4mVYyO+14iu17uRumqX9
jKmlVoArBOvQUN2tnm/tgUTWR3tnMdrnJvoJbdgmXCQJODQTIlukhgddaTdQHMgv
znTg8i3vzvRNYXUOdwJYADeW5kC6u3H1XRL9tWhqUsMZzLP9J6+xSz9RgKjIdl/M
XIZKEA4ifqp7mSYGaOz8vuAzy7MXxCWOhemLwkbKrnaF1UeuHjgFeoa9sjonfc+1
OS27APXh//bIxXm+Dhu6t3JBsB1dotgX8DP7A2zURiwOe7TA/RfYQE/2pqroSgGi
A6vgHPulRa6pWFSqbhmKpmGtBFK3gpMpdrDbNQ7J+adhOXQZGoP5tQNLFGKAhmo/
HrbXcRTj/shLZBi4SnOZ/7WgnP1eLMfVpJcCUNgGRnaA6rlJg4ss+TYZTkj0MQpk
lv4MEMpw+L5mhU82MWjNUlZcXeLoOz9mmCr7lB9KdrpF5PzVDrNdDDa+mXVSO2ld
gpEbm9cdzLpoHsa76WIbQ1aPBKivKXA04pkGqi1XcEA5WnbPn+2Ojc8CmB5M5lcd
BZAxTjUlB25iDmb1dL8auKuHz1HClaWvMmPGNRwP+i4ls23qpR9RWwLfLqns3Ibv
LSENFvdgXUomWPi2s8Ep/QWx85DHZ+2L0zqS57XZxda3c1T9T9xoajVQ/xd1xiUC
qYtkSOFugeSHU4qvn7ggs/CoS9u/HAwcJdCryrkmSDZo/baLdf/CKZiC+mISN8ZF
6cA2d56DPE2j88huBHJjo/oltojTPuuwHvGrSdScd3tulMf0zXWkjEkUMyBsoD96
nf1dTk45+HWz/renCRjRC2MDrGIrLgXLKicpzhx2quFxGiSBLQzTJZDmZwE/DkZN
aqGznyvskkb5qCmA4JlelGlyYblNb6okGIRjqiZ6atvnQ0fFCNifbR6Drj/s6Tfl
NvfJXOqB/C31zFysp2oC3j+V6TH7Ey/t4zbZyCKdFICl5lK9dQrkd9DtZB8zpdfQ
+65qsFFtsYNh5jOF2j7PhCc3yWst/tlIKN5FoRo1KLToYAKkxTbAvvxB9tsa1KVu
TM+Hr7woIeeJysmqyFospK2X8owTEffrE5jKN6ExD+fA0TsOvZ6u0fuX+91osSmZ
Cs987b+4gm8cmCn5190tuEdOAW/h9sLLmDDOM71AQ/PAUrb8pQnETGwV/axx1lrC
nbdpJopZKpYf3cJ74+9i9szcSQPOrlN/WyFqpQDSduUQ9s1XR+pVam2fHLwCVcZr
F+YYN9uj/OPbPFDAh4EeNgqQfKeiCOG0hM3GsoJ9G3itFW9r6l36ce3gSlNKGqsW
KWXYHvdW8rN7zjQQVFpy99xuo//GcfQ1mJymmT/AT0gbesZRb2cXh04IfA9ieiPA
G90x6dS0j9kratxDbcmadnijx9XrzFG1zqdiL2mqLyvtFwvimQVTIBhF04/Dj/W9
eCd6vnL2evED9V+6Jy8xMcBrxf0cOon4LGWtwTkhM2kufwjW1F//tjHc5BFzgJD8
9hNXBmZz3sx2doZbVTsdmyhlOggwufUIe+iYPp/iH51D6KCdgaDbjXQQlNZQD5Iz
vPWX50RgXvY+jyEYW+aaKWUdfIwC4VN+2lZsa8nOeaqdJ/4MxEr0oLUl50vkOd+F
oOsWFlbffmG/heYmBd/UABm7ZdrPPNT3ymwBzj/n05iyYY6kDrIItMxBA//ErTR4
kZJw3B6VS1DoPRUkpEV48oRvDOzq/cqB1rAGrZWEQjh+qQCDvwIsgEV9/aHM+QJv
mBlSVqNKxuPTy1ny2gZ9+s+UjqjSbnd5SuYuimJX62fatTO9aVGOAHVQrNvvk8f8
kxAOv3hiqqxEVQ77CuIfeXCDDdF5717qy/5zDt9FHgstw8Qyzf4+J+HiaukPKmtJ
feRLL7ybMS5HRePwH48HwDOH5CDOdYGUA46PBn2PiP3HQmax1+Y0ZgoQskdQ4cfB
p+sPN7C2iDIvF4avj4HH1sOlfk/YNM4x7gWvaaN1pMVFWGcn6dY4HEUTfMSiwuRx
7DBjJv0MlpcpBDkiKJH32IZ5iOeTqTtT2MeV0HdpoRG57j8YI27Dkyv+n4ngGziK
BnH7L/8JjXKyKdjid8h8EWzIDrRx8Z5daWs61s7wQLT51bE7thmmLH1Z3G85iVpY
5vdwEGe68BSwiAP9kELnsXY+JiGYSiW688rHjDfzPPNB2Ag/d+OJFDOsHHCXlBv4
hlx97mPdER1UPFVzG2H7GpD9oTIhJG+GAEqloUA1V46gZysK1LLCfDIa5opSC52t
cgazHz8a2iOGlxeEpmmagpPG3CNf1L6UMkhlLw48VpkyZJMg2M6iXswLEkVaKj0D
6kIL1zIEWIYyaVwxQJceV+PAAcD2dveXI9nIUuIfhvbA3iq5FzPlbzi9qYhYfpHR
j13bTgp/kyfsm7COqcDTlFO4ZMtYUauWrDz2ApLvOdfynwc8Owh245sxYpJw+xZE
wV0Gw7JiyyVccJs1KbCmuvHNbDYt5rcWACaVLtSPkK6PkGKCbztRchXuiUWateWE
9JdxRe97G1mScZOrlzW/vFQa7jW9vVaLVWhzBDJ0bXbCqjaBvxW46bzJYVreShvx
z9Xmlc7FqcIHCVBWIPipHpKo2EeZBEZCd04VzcuD+VwNwEQKO9Ruw+hPZOwFsirr
3KDJpiKD/hNuXeWM2rGmfuyM+Sujx/79SblRoJVPV/6DqAXljYRuzSTmFtDY4YzJ
vlvMrWoQU6ZtLVduT5TnlcbCjp65vEjYjhXWsnEGbrUi12cfvbYKgHzSaSN+EQ7z
Vsre5pmeEyH/DRzG7yPx1Xc9lrlutqCM8KLmV+WzSMN3A4ChpVo+YjrQhVpNl+AM
lyt9BJtBudt8G4XUaF737NNzdlOmD/5MwBiZ/RKkA/e0xEXNlY7zXp7wIDa5+AhH
kGqCG2MSOZBx3VrbW9LVPFRlqIKTbt3wHy+W+X5Ed4GuXtbjMEjr9c8OxQMPL7sD
W9+tzmXTI5ugnB4mWzPA7MKRZ+RpHL2bLe4SInmLmd4rohd3Q2V7JewZI6VLgZ7N
M0mNBwcMXss+VpE0f0EnXx45z77V6UPROjO9wuW3k1Fp0imtsp7yk7P89L3XGiLq
80caSGEn5772cVdFsQza8iVEZyHddk+z/eut7V8DGc5xnaUxfDBEDCHLYvRgCSuM
tN0zjQZprQl51cyol53TdV+VkTWDqhwRmWjs7ss7j4KJvg27lNo1gvfExWysd9fD
2RXQkzZni/3C/UVudAgHSECjopbXL1qa3LHMjG77m5Yde7VRj1sqDtgFxdu0dLZZ
qcPa4U3TrmkaMY6ueRvSCnSG2a0fbWYVGoeMGB726pEOZ4YW80MMhnXu6CYa9Kgz
1yVoPAbRKmeDfD9FuAZaooc8kklZ0dCOiumfFCegTj1WH8lXSzWgiC9BkIw2sD2L
8NgqzeFlxMb1SV/dNj0u7WY6xkICVaOO+s86wViP8WM3KGuRWZsenTS393W7/PEO
4CbEVZawSlqE/3r8qcZgnxHY0gxxHamD3VimAoyBU5DY9Wx8xrxBNDXNPGLg0PO1
sbjuQVcSfdx81BvoDqqh7t3vIzF+iuB/o1XLiCcKcTekb7isMpyUn5mCt56YZrCf
gWxbQkf7d43xyAOYPSlHpNr9Uur6ZteFBFA+GVGoM8i+/bQ6dGJN/Z10YsbV5Msn
4NGTmQfW4FBuVHDUTx2bTGhwlX/t36DpROINFDD0tI55gXJtqJAi+1I4+Hx6gFS/
zchMTU5f5K4SVhmIaWuPcPBYNU65sboWQjy3qYpEA6YZRPr9Wui5SEVCqSuCeM5M
F5cVhg/cwrCIfkVO3PT7DAh6G3Pmw/TSibnzyl3LA117NbTvH4mG29M2pWo5HtQ1
8Ipa6axryWGYo7RjkScJwY5iifDyLxCugJ5vwEQ7NmFeYt+QBqQUM1xkzEcBNlTQ
B/jGonCTF8rTjMd7AH4r7jdeubsvQf1ijF2YtvzT0xtHFsE5YByMv4pBuN0FtSH4
AdlZCOkbIp8HqG8DrEFT2q4LQJ+s+CqeQsTlo/MhMwkg150lnAjKktJFnjpfGQxS
mdMgsqo7UrIRY2prAdVTty2A/HUxfh+6+0g0DK6ABsEtJulqtmHjKNQT01UbmJYL
sG2a6qdwco+yeeFPTt/A4ZPdV6xFiPzOOfZPwPby/C1jljHV78kXNrIChab7lRTD
c7owW8gwtKoYBTfi1wcXE8vtY/1lFFzK8SxZ3s+yU2BnNBoDqeKDNL6/d6ZPGHQh
7483f0UMvpGg9o2ZcQsDZo6S7uosZlNyADOhywLQil1I+AFc3qTvlvIdA4CaoaGw
9nCeP9vT/QIqk4fVNPDXoxGX2LQoP5MKpCSViD47bY2Pg3+OKRvj4jteeL1uC0lj
zS5KH1ibKP5qmeEgtrzlBijR9pbYMjQgF2VorvZaeidbT92d9pThStdnn2wkj9/o
ytvr+e+42A1ZPWdTf209jgHKC1GrVYaX/OW6lgrlpX1pNqnU1r9ronmX/iuZEiwp
cjELClJWYRNBtHdpWvYOU2D2nB2rvW61hcpsgsm5GIoPyhME8B0SA9z1Kdmukvxq
rkqHPf7TxlHRwMeTNTCu4/QSodvSE4d1EQN36R4RsfutdgtuzGIysNGotH8mIuOr
XNC0WG1gEQH6vKJC4Knz9x9GCJEpfvM8/RmhXHHHXtDJEyoDnoOy1uiOPmWu274k
zIeTVIgZhv33jY7ixfTRlyaYG2+yDbujLWIGrjaAdTaUw6CeH2DSrfNpcggp33Be
pTIDNRRZVmCbcWiznVPNlz+WCmzRuxHZmDVpMEw/OovXGY94fKh1rAkFZZZZjCNp
8B8cJ0XuMojjD2+86nedc32s6Q5QyAC8Zkw7mRrydgvW90VRo0PzAFcgxD44fIW3
vnQOSo7dMrtfBMYUJvIq5IswhI5LuJiwk+KDTBMsiKs+rzckO+2uv0Uw9VvXlK/L
Pe7Zvp++jHfxG2V7rgmp2qGN5vwH/jmuWIh8NTIGcyOyd/ICw8iFamUbqr5WRHRZ
876BHInuG2XTrvlif+6S2zE2kYvs5fu8eVcivpQVmBPn0lsEXvS2AwYNOnUf8iOx
e3EsxFakF9ftayJFp5kLwG/XaLknO9wwugkwh2RkPLiQqVEloXjI/qA+CSI+BpRn
Azxjr0qJCEuEhlI49yDCfWuSMTvnSi4/fZuahx/0fRmMuovq65q9Q5jguFt6GA/g
PChCirxX+jmsa3hxRl9rxAdez3JPckVsANiAGXXmLHiWjG2g6dJtoxacOyswBx1U
zWcZtfE3NNEqg2uN1KLVtznRDtD7y7YWJ97T01lz4rVgkuaR8JtUcbPElhkVvgud
iTmw3UzmJmVAHarx+jN0A7K9uLMIxyZFJ/gRf8Vzhdde/FOBeRQxSb70q258FCMJ
gf0BzwoAcmEuxXJTNP81TRhZRZHQKyLxPsV0L9QBSHNOE2/jppPow8bt/Z9j2/Mi
KQYYxebGSgI01V1KQ4/ixk/HJahtUIxZN5MpM/euMAEoYREVS0f+i3tfJy75khmr
I1D3u32HsEepRqLnqM/8A13amkvt941q1VaLtLv6r5vss2pqeG1bgGp05m0IYraX
Mya1+Y/qca+KxZCGLYhGLVzGc2QNJRJz8LOYJQ7z9y7lGCkC9Xk//0pdeg65az04
sM7eskzOduMa7BLmbuNVR1wRqoAkACLaKzzE9bVXFAe35JN2qA5ueTOqz8PkSME9
HG47zXVtcbvEGD9vn1te30n6zsdHAToLvhUtBWbS3ws/gB/cDO5ctXcbypYtnC67
DqgCyqklCEL9P2AXXIbTriAfwcXSrkIwg3Yts55UUF50wv8xWrNr1ZmCktSamg3s
1W3ySpxqFNqMcqMNFEgSPW33TEv3IFeIojV/C4SOQHwtScP+ENNkbAN3RuhFj423
f1YTj0n36SZBo7fg5h0NbjHtcBIRGOPgv9Ua2EYFeS0vAPgK7OBfLi4K1tMhq9+W
7XFFyeVX0IbX0vgzZGUNh7+69vvbA/r6hmCL5Hsjxrd7jeKK3xcliF+vib/H6VWK
2UuK5cW+IlEjQdhCe21Xl2Wx7YI2Ng1C3S1cvNv5irR9Z3AcgCDAVhKPLfU+lFnv
ts5HW5RyZNywjME3nT99oaUOVZO9YUQoSSUNDtX0uBqBNG9zQIS7Fe2hDsGKBSy/
lhGDHMSXW0M1b39lJVBSwbzM28/hKN3GMhuTcU1wiBoxN+nZMToePuhBLj81cU6W
pR6LI3qlct7fpnlEhvuhJTpx4Sxq7gNvftuvP2NOYGqhYdKgnAB+ZI6QittMnWlK
Ran0y6oII5MCHRkplscnGFA7Q4aTw6Fg1LEP+DQU81dw0RXuy4QuxDoHMTznDk2/
12xCtS6dLt2E6IlWEDBYKuOy9d/NOArDKYsIZ/BVXllW05SqTLa+DNluM5AXwR+e
dTFw1RiFDA3cTNw6vaGF097I/xXlgK46CFG1QMUjk5dfmwux6T/kZFh1dmt77RQi
5RMS+OLrgdwnemkfOitzSzOdDEXnSv013qD3vfScBBxAH1rS67gEh4yTS8aNC0Jh
qQG8TvhFqIJVSp+FQ6P3h7OXCMN5B/N8MwXWepJjmVUQKHxmhlyljBaPeNrxB488
2PxnPRNilVDnBLpTCVPSqwLC2mI3yGUz3Z0F39X6/ElOiqKoZvcqynyukIaXgdxm
redbDbyGog9wgSEAFxC2Gq4pp1S00+LsMMxE9mkHsYFuGCPT1L4uep2ZGEXR9YKZ
G3ukFdb/LnT9ZXXlu2MxjEEpk7f/zoUJl3woKMe6BoxW8kuzpPjaro8FJdav6KiM
dNoS3cEbzd4eCj3zf/ay5axu/lxvlWEyopL4vj0FOPzOyEu3Cw+Oz804snQ+ZNSk
Whx3KIaZeOD5FAzyX1HT8Pph5K+JhTL8EzjN2+xMLk7R40t+/Ayg0IMNKvSvKZd1
p6WJGqoWDunSJ8zLsU9+x3BXO4t8WWZCHB1Ag0A7r9TL7KvAWqMZ3GmnVj4zhfcM
rNbMyWznwV01eaFZuiHd5Vtv66mL0kiWJGVky0L2UWldH1mBFwnjm87QF4kvw3cc
vnqwyMraeMVsj94doCMpJUrDxqAm1DRpLJWjszRRP1x8B+g8VBzZ0hLK/2UPZxxr
RlNfEqk3ZqZguFrMCxkoyBJB70oz4FMsXva+Sw9R6plQdSzpvcbY3WMI43J0N2yI
vSNmDz7SRGm5TR96rcVMKzwbhBb4MgBaVUqx4DayAzxqsS8S+bhEUtko5WsDAIA/
PhylQc+/SwBnfMxtZ0HNCT5QbowS+NbrIOH5BfB0SH2fju2E/3sG45HWCj3//NBA
qCEdWULsQ2DeTlZ1L7q36XivfmmzPr41g3PyucMSaBA0bwHxg9oXXSKY6hYlIDnj
dlRNj5ckIto11pfkhcWX/OOr/+3xM2XwWIPwtjXb/GjoP6dn0uUbm9lmAPlQOb4r
LneK7fYVmKxDW6VnkkvXFpyckSSJavGTMWPtiuToX16b5YqJ6PZpVidwj1pj2tqh
m1HLv8Qa9WuClFDVIHGO/0rYGWFSRCAbI72L7IrDbfsnjwR33EMqJ6qDO83XsF70
g53TnNALBWUBLOxnTkKZfk9h39qhtaqY4XyjTTrKuRjNKe7J8rXNmadKK0/bDBxa
ve9CF3Yeb2VLvG3XCSAIwDGKzE66SWFk0fjC8ogBgqRVHASsl1VJoxzIVuohe99d
3rWc9ni3e7BJgqcZT11f8+k2lHfdX9bl1gtnk6Ju2LcvB52W2uxosoVXAVHNf2re
K6z8u/t9Acx7GIyxqCOT4Nqrp35YuJNxyGRDztSyOXs+PRNyaQu5+g9RXa8x0K8s
Gl2FRFECgz4vEiqYb1giKl/RN3rvQpptZw8PwtBHUAO3B3IG3PwK/dhRIAq2O0lf
PyMVRYoQFmdKurdQes5BCvFMBPpPyAkPEzMr37I7iaSrBgA50wfxXdLT2Fcc1ZAl
9D6RywyxIw1pdLOEufGrzU2aztpHjmj3/DSvzxWP22tZT6G+2YE/c0FvCo0wqdhl
zR2Gc3C9HX5usq/DTHGGrJ7aEpSC5Sso8VgBu9DybKCoPlrt7XMwvP2hsmUFJJLX
/aMGedrlDR3Zrtt2QxvFciS1cbvOI/OOHTeA7SM2Z2oUcZ7ZethDXF5B5XqQi05n
Ws8RTan2cFcTCi73BD25wNIoiOb6gSxzYKpyNdTBCrxqFeRalDeg3apvVjeHCK27
92JoO70YLXbP5cjVvTHbtxBrL52kuFw+tTxrdoUq5Igp91jakct57gSokYR6UJlv
e51k2z3iPTD/pDrvwVagiNe0xDT6+CMIx7+BbSa+44bH43mOZk0BASY0hcM/L19s
AP5bupTMI774M4BioXW58hGrZsNpcwRE5ke8TupE81RAuxEL/LoMmhnOmZObDaGV
SCOhDmUpqWef7D1PEPRgpbQYn9HIaWaytE34RKd/BZ+7S3SqguSdKbd+KMmHrIk+
3mxKZGGXth3zfNIg4J8Quh8AqjMh8K7wyOYVQPAtPiU56KsuZeuQwf4soPOiGmKt
yIMKA368VK+0Y1kKFpngxqt73FqfciC141uFUtCaNxkK7/0y9PF5Sj88fcMN2/9H
DUkCFwJsTEHcaMR73JhVJL1uQhs1tpszSJSGI4Z3DNm1bMx+YerAe5X0/48P79/p
cnf7CiA7GNXPTYvsgd/uFexgKDDJTRp/AkkU2HCTzSLR8kNCcV2652OKzJhIbUJB
HrIQvMaV2zPMgIf9gZrU7pYTC52ITIFnePDCGadAqTgcOIU+OtJiUfdErlG+zKug
5M8e9BwU9FwtoVTrwF3Oe3l9v2Fn4wC5uVzcqcXwbw6kITKBo7TlWiepriEFNINS
brqF2mM1ei3xUDt7f0ue0Q263Sj6vqPYK9OkRTJoKO89u8OCch4MO9QtaLBqFkbH
IenbMS8TsJT8wOzeRa1/5uFQXG0+7lh0M1U+F2lsGl6UJBITyVFs7cuKQKFXz6vZ
Zkx/6RvB93iJtEiblFvVdhICQEI/JwLAG6XPnLhHKSslO/eMfWTAFSzcrlyetONh
eUoWNbCW463t5l9TqyuEKmp9iMSBwd8oYA+QWGFObwcWrZEbVx1KJfUE3+/0aIQs
8wDRtirG3AWd50yYY+FAGqZUUqplADexw8fGUGvaqSZfmuhjjwX8luX6VkBU4Rkk
LGqIVqxcl3u5r9hXtjdfxF9Ao3HIZnmQqrvvzoZtuQPNSxN0rqLtCNyVmuQ60gnn
MsSLIZrCQuSu+pqoKFgg4cBDFDEi919jpE+h9wrTlwhoUFcd/N/AtWvns99pvFFq
DrxbfB+qk8IvxOYBe9asfX+8WfhKtVI2cOrcv7rR8RKWZw9mez4pOZhHXVQwUX1q
cxcYWfjd/amcLvYaAqDpWrRi/4QjU/fa2StHi1gcBUXlOmaQHxwCVinvCqFR2mSo
qwzXlHgUta5J7bRjuNRi6YZpVaKU78NRD+pW6AjF/Fa2lXUgX7XH+JocUUy3vP53
jgPEDCsi/TZL3eJinL/GvINloD5+9PTIosvCUcTj0qI1STefnD2ttg+aq6408Xye
NTAVRwvcaRbxQcTzy7FEET9ZGOVHGWy4yU0nHT1Lh9Rtu1stCq1/jDECClMzLgae
8xebl+lJ+gksxsqKqFXfufDcxEgi8fFFra9apSAE60ekMUUy03VxKvVu97UJKL1u
XY9dDH0nGDuFGeh4cTB6nZ7bk8IEVQ8pDCav+1LmRP3UhRgOxchlYP16DGaq65QA
CDUp3AgF3kpb08MkK0o1rEBFWdy4XOxe99LFoSoP1KOFEklxi8f/3R8kFtAn2u3Y
tENfyeFlTdoUBvsNI5QZwR+VBoQ2rbWVZKMR89Hg4q/ylg3gUloIOg/6FBYkiWuP
Gfq0lackvF+FtEVcVD/UwYPBrBT0rNSAzsDa9U3Q74xcGIVOVGn99isjF+yuJmcB
cCCu8yRHQeG/OVPLT7wagH7Zn5/Mkd8Xoj0wqzF9NO+P5KlcHu50236RXwm9Imvt
HGqjH3MbsUW+HUrP7whIgd95lQHoY3kvdLU9EcNtPpadhPdAOE4U0AmwyLAYUe6x
bcFEF57i2PBcGgXTBBPcm99MKlYWNrqbJXk0AHyiSckc/DK4iNdOHLtYB3uQSUHH
CcVvKr5mW6mqO0ruyS353d03dBa0JA8Ojf2RmIkQD+g1sw0iWVa4olpusa+mYARd
oDNDdMDHCNTpbEcB/jhlsDRQvy57KJ1rrNQ1gusaJt/R2RBr8hQwLJj1eXnRrywq
FkmuSeE41k93NNAEuVcn86m1lJcXiYWbeANYRy0YJvRZUDm87UuXVcnCMGXB+4Eo
g2zhyW61cWFAgT1YGk9aRdpZ9xia9/0LGYL/jEUKX5apVivwOmU2+QZQ+7t3Su4q
7+OVkcqp70jYxl91RoffqzntqYKk8HHIRwCdNqLNf/AAUBX9mJ/4/qRWxcvKeJQy
UKyrmctyNS99Yo/xo1c5xf9UnySd5Q7b6jRHW7gvWazdepT1Na33RWif2Ai3NqU+
vNUyq4w7uMJkdrTiCzvbFbX11SC+79caXufLJxazyLRk+slAZOK3UGZi2Bmr90if
oHnOfnfOSQWI6A0rDb/BHRFdF1e390beVdxFPTp31dIBI5+pPFMzCIru3HIINoPH
zVvJzTKA49yAnvgrekbLo54aEALw+NfdbD+ZBwyGoyFO7ipic3EGPCfLKMuO8EkV
wSX8vF8iPkPeLsD1lI/97Prsm43RbgGUn0sWgobJ9tp3ke/XJwmrFmpdD9muocmK
yymZAbXdqhlvNnKtIpbYp5vVnEC8TYKeifPjECZGrz83rZij0RPzNNTerslVnYHu
qPeRuFjV64hKYAEda1YkJ5Axn0VGv0OR3NDLkIh4FqYRyNrI5DfeluOdfUjY3lPF
qshIyD63NSbB8M8NSdUQejk/XFq5Ywyt0YwHvGMzA2yht+k8T5FdZDFWckpYswrH
+Y4ZVjiG5VkHwBa2r6fxisn7luF0tQ1BLzY1uk10lwouE3h89dp6HuY8GyxcDAyO
muH3fTWSNUBgKZD9AoAJMddCMe/bazdxlebvHUpNdVPvLjTApxoZOhLrn/v+ZrZx
WrrAao6TLWfSuYv7g2jVh31cX0zbWZ3eoqjLe5MvGsefsvvMpUHW2DYyAudwGiSu
5AaxgaibcmzITDopiIiBuAgOSR56abPBGxWshx7evZ0LqvraFbPswPj+p1J7XnNp
K28ikLdtPt0yjmsE0zCn9yl/jVpCF3vDNvcnqQHSeA3KUXs/neLBpmTRNcayGN59
bt+94jYagcyGVv30zDgDLqO649JB0oXo/mAYALzSa1x5z08z+FrWES8sR0EACSIs
59h8JhO1S9tulCXZCM8EBoCkCkJFBL+uZXo3bluwroF2ZLV5sDsolvAe+QWGUQbA
w3lmNGK4LV764bA/bY2j2327QpRPE5LrOslZscBPjndzn5qsLoIfZnXVtflNZ25Y
RIQbnz3+coXB8tWCtbYANKUb/rs5gL+9pEW8S1AtRxaEReqMILa3r/CF0K8b4uco
tkQoJ5iujNnyyhJP7VJIRLZlD5I1a/4b8HS4APd7vWDY/5vZguCxgbdD8Y4+PrGl
uELYnerqtOQPc0OaTfCMU2/oAtOP6jUCg/Dw3mObn3M0r5ByeibkhT2FXehRb+Su
TwRBObtszxhQHyy8YQa2/PYyKsYfn9lppcl6vpljAjSY754Is8hJxY610yN4nca+
2Gjx+nPib2vR/hY/FT8whb9GkEX3K1p2KlLVNxJoY+ZbtvKIhyPIHtuDL69NlyMa
BF3oU1ZOUnSXo404UHK+DBPtrvzgWB1Frp3bmqTBqa5Ug0UyNqCqrIlDd/xdEeuR
cXAYeQN6AFFZGt0E8D6aXRLZrA8uOQlluV3INqt76dWuhIhNIq8t0Ci01PE5LffQ
LcCsJVGyHNBFr0i1L3Xf21SObVkNfT1fd3nmzndM4gL+4+bhE4CZvZvfkz/x7EuP
9H2mIGGRj8W3YLiRHCEB4rsRmJaXTW8RWFZTK5kpZkMZmTkiqeDkK94OJx6E8Y9U
i+jjrNd0GQfqO4uwC/F88/9VD4mPajudvutKn2uGBUKLBW5i3z50vJK8pTeD1HcT
x5DOke2lgrnPpVHEMXeSGyCEBbu1dJR0yBgrqXSA8HP2XQ8ylvjribE9ceKP0MQx
h0YLhTLHtdfX5ndphCgpdzU/HHt+n9uaW9xREAUluQru38O3HWQ0G252CDP1CRsQ
NzoIPK0GWspsoDESgK/hjjawgeAI5nZg/yn7bxxqb8Q/BNOsxVB59E5sou5QI9Im
iFO6rujw+TudywnuVRtrqfWkLQQHh62uvmeMdWfjjH2QYsn+qV5JZZHvZTTouo/b
nzyDyL9aHcZkFllwrxe0yhWeX2rTfUZYfblhaOI1NuUWhv+ZYfciwndB9parzXNl
aFRPnhXsXXjq7cCLRf0AywKXbud5sqPI6QXpUis3FG+d0DpEmjoUFk+6pqwJwq8m
BA1tpigujUUMp4Pg2UzMR4maKwThJC+kKPvXhVPmudd1HAeveM9uc/S0E6w0WMpW
/0YYbKAHnEJRgHmaWGVjVmS40on1Kw4Z4jpTvJbUgd4zPrBAOxWYhDZLVTdvvTwo
rtHHrd/RUCHZegnvCMjz5VJ6dsWRYIu6B294P224nNE/OaEq1Ha9cj+RxCx/eSnj
124gWFPcScC4E4LM6m1Fci++c5Reh8o3jkDzW/RhFR3z9/p5W6UhA0Q90cagrK4p
AQ4MPG7KO8cHil/egmRBnAGYRIHchSdVtbvgMuOTRf/wgAdUouOgDisCP9oahupc
/+eVz4dsTf32KnIE58INK8pj046nFwJaiOlvxKykIIsd7GsLe0RsU8+KK9Ivqomz
2Ly+tcFTFnaMiOs3aci79beQ+TlDjoijkzLm25N0wHaponY59e++zzC8wsNKQ3xH
SKR7lizk7bMzepZ3EqwduyfVq+lXywQ5IcTIT/Myjt0l8XPK202tcHmtoSRJ5iPr
tMSMhA8D6wuAMo1xEKTW8QwJxS9AnluRNdC7hEwi61pcJpZ8oDT90ltvhv+P1MSw
Zv5RUI+bRZ3wDwxEOqbqeRETdB/BzDrsvB3AXR0ZWtzOLczA7xo3Hy0Yhxf8CLUY
F88KkffEhp2Mqsiyvp1bD2gkIVrqxFGZb4/rUF4fVSa0X6E1T8SsiHa1agEh7zgF
GsSuhqHcZ3hooGuU+M9uTwUI4DSBJDVXnVXihedL6IRDLXAyq3eb2P1ulY9c5v9Y
KIozF+xluXcRlgq+SwVaszkJpTQlTeA3xY2d/IXxCtPGPW/7/epdwkl/UxSx+c7H
9uD2w+JRO+PUdSjCRfhzQz+phuNGqLI4SDA4dTXTVXZqK0fDEsyCQiIXeZpGF6+R
BiUJHiWaqesCwC3qn9qnrPVk7nzLmKZRor80x6LDJ3J9pZUhesV0b/msi/1j4tAe
Kaq6KlOXO0Be6qSK1WwLZ4dNtcU59fK66v7KUtb3iDtGzw7X5OtmczC+BdRyEPgG
0W39J8dr0iDt2Lr52RUEhXtlZ6an993PG6kqUHupu69RbeM9SnwxWL5Gp4qstjof
3NF25EDXXikGn0sED6gi9i5nFo/LgJdpaNXniy/HQZjN3BfnWfpJSjrHDaiE3ulA
L5kl19uKdAN3HJ31+RUTurZoEYgCAadWECK2kfmxHHHS2blJmCudSOL79NkEbamP
4TlqaUKCxJ1cFVoJknLb+FO+sO4GRqKOpRD8F+xGRaggP5R+7Txr8i0Vr+REWG20
TydwPUlHCMbhgrB3IAmNxiGUk5UL0lsF7p3G+ZJR/f9Kt6X5zsmez7PpenSFdelf
3gvxhqDIFTfprDufIlRBHoWW3Tp821tMMlTl+6QMHAgziDsFYHvuvKDnh3QyEYDK
2g9vq7D7zdegT2E/eY3EKf/XR9FVn7DBqeFMuNIar8Z3lPr0vM7NKI/EXKg8L63g
GLRZth7CNyPFeuO1pT1b6xW8Yi74k44t/hWOXZ3HVaSQjcuuHvHvvnIQ971/Q4nM
4+KQoqWV4EuUYogn7Asx/Smaz6DERa3PtSvJE18K/SIAFaRl5mA96YXHHLyyl53/
oFyERGbFlpYO+G6hDX3JubwHTUKiG/+a2qBd97RSYa2XBHmupYcPRh81VBL7eEYt
XIWFu8e10WZq0hKg4h58qojjEo4ezXVI5LcfBUquiWBqJASt6HW14xXuaJZDy+Fo
wLD6wCnAEA0LnbFgsFEzNgcqzqTb2sj7tZKAPqu5vGfACOFjKmkEHfxUOBv0bl+J
KK2y8PAc7M20jiZhlMSS5MpyLxrD715AhbDXkZV8MdB/McFJcFNxvzl2krmXOyi9
AM0ddVH6vMTtRb6bFS4ophp8BhuUvHZb6YVlmxOSi82tT14yAX71onBMuNWm/H91
ZFL6CBblAS1Vnj0+pmPvYRKaE8BPlhwU6zioGHi+1ncfmfeJ/KMlCeYOReZ+HMOR
/LijggAcoXkzdEK0n+6CLe9klMqx6UjhNmJ25TclhRhWV5ZdDpm5OlvoY86ZSTga
+bfgoBKI/3742Ki+TCMMoQWcdK7tkFuPKmqL93g9TJt89weHVqJ2IidnhlGMTD9x
R1YSrw7UBpjvQj0HLxi3rvh36B5F77novNvDkpmHz3LOKwc9fAIxc13xS/jRSXEX
/8aEhfnfMxgZBhvrQ3HGcqHyvgSgZP3AvJGm+3EE48j6b/QIfgiaCmtq9Gt4ib95
RLUj/liL+DDypU9h9u9RHVlL25eeDxVo8fZNICCNLW+cHFiB7NRJroZKh8Ju2ZQ/
ZPb9ou8OwD8WRzRYOpTw0zks5wJuX33nBy8xL7qiH5fFf1qyC3tXbEskPS4gfJoL
yVWTCzZsUL5xWxaW5wFB2cZFn8Kh+KtYKzHjYTMNcNGnV/WgnYQ1hFfWGZyTXIlv
sEQqh/TEl8g3fp+sGp1YT9MAhSFIc8mGW0/CL5ZmSKuW41S98glDIgvC/RxStBlP
NlA/I0xYQuBlEA5iQ/S9qJLykykHZAtzGdUnMkIvDt+OQUjtQ23YAvNu8MNnrYvw
R6b1BcvMIMsnZCTAuLtQUA1TB+hZGMSLXKxV7E0FFi3EV1KIuIarlD/NMtQMbldi
+FcZhmODjx3Dz7ehV8h4W4HMcbYjVMX5aI+HtE7SOBHtrz//WBtnz+PC0NeEQlBe
XWs9eoL9abvOsCCXd+Flc1a+i2oyBbk5hpMVemlXXLx+nTcXIRI8GZolYSGGaumZ
UyystUc9LyzKQo3mFbbzC1fUwQbsPDNUDq7JAw8gRHYj0d1XQgg/yYoEqWMDfUvu
SJQCzNphuT3DdNnsAjH6JOhy16JDbWqCQg0YZbLVmxmAXi/JDJxHrJFJUbIaE8Uu
ubx0q1cTFRru2Q5XYLKWI2pOqNa8zVtO4EqVsJn0W9OGdW0dDOjhtsYkrjWiWx5g
uKEu0YGT5azwOI0zcELA3L1+QUQ8MjOvuhf1f8E12r/a+6gJVnZFBLm5RHG3yi80
klwZ13ISrhHFFm0St7wsKlCmMMwEoo08/Un0b6PYa8gPmEe+5UwGp2Z5e0ng2kzK
IH+M0r6pj5pjkvN+UxPQ64Mcw4Qa97w6Zn9AMr0AQT9/EujpF3JdhOrsvqVZlCYg
r1T6ZoQawRKrRh9YiahQXVHVW66JbDbIFnByetjfVOYHSqfO2usPUhjYI9zR0hJF
73MkvZoIIXPLyJaTw9iGW8My8MvR39SKf2tKuVU8RNLp4uJZZM/0zMvYog1LXAQt
rjxmjW/qa978kg71j0Od8Ei6yNbffl7jbyXddpq+N73p9ZloadiI8k5gJC7Pu0za
ziu7/zIW5U22PmXZChBMUq7ZaIp7HMX6YVfzKx5wyaEsgkC8JrOahpfOiTSwwuKE
otGzABlIx78OOiqhS9k+0rHanTDPe5uDANGKhIjDQktJPJCgkN4rac5scyUmk5p9
Fi7wmC0ZKGvrm0SYbrodqCTAt7vkdsi2oQxVXhhVR1skZ+EAiICAIvkqBr9Wobb3
XZpf+Oa5FS+Jx9k1a2x62uhwlPgLRoAtxIP4gqn57tOGAaAHkkDuhdE7NSaU5F/7
gVmLmCrdHQwsbsc7YCDOWexPcZ0waQQndcPO2k8tBANPlapWIbpjlC4g0FyrJCVJ
TJNLQQZW2IVmxodc6ljgroAbrH9w5BvHd762HbCyzc+ZCFKWrun3dz/5NfrD6V12
Gns+527tLD6F5Xkv/0f6TwNy6AUytPddDqWWG4r1OFJ5/4J0XSvplAlIJykFmTIC
3ebHdaLYWmZGoE6IyoMjym3seHw58qz7q54fEmBsnowRnq2M72LUqdErnWVtKmQT
TTPE5ZLkyVFXCU5VF8wELeeXrK8KxMyRpFrVlMBJZ8CraIdbz8w7MbkttWaDWvN5
kN+Oy79Pl/3vn819PFcznSHBfZyQ4wmQ4nB3qVS1LuYoKlcvEPLdJRxO6LmR8aOO
bKMQ/LiQXOQuL6+NEYHO0R4hvnt8dqwEkhqYgOG7xLZXlB/ajP1/oiJmC1uApFQd
mtIZ3Yp4QxGASRZ/tQLsj1iL9JVECLyHHmVf0ZGpf5CCL2JJ88Wq6GkoTVup4Uc2
sbHiYaaIveATRvuhjAFKB+DrcCRzWM27eOj0e5iTKGKVgZTri9JPfrAgh6yrWQ4H
+ck6NgzoBk87T1wrWBcVZ6CvKNyaapg5fiJ3axFaMyPuGEFXil+t2CzTrTPxWmSh
FGjU8rxaRpSBzloIOYKn6ciHCFuL6juQ0J8YWajVIRETyoVUNsbYvkLbwT/8Iqyz
SzZj/ztG+EegGpji3c2nYYg8NOQbXOnQI27qfrJwb0Dm/xJIIyNmC33s4R5CPl0H
/kGO2PJlHbtmzEKPsa49RI9rGZC9kqvvn3WietmA92ez5/mgbfYz8WAjjAtqPNjd
zUf5Wso0xF3vhbpwYdgXbCHU8tR+er8rmaZUDH0Bkh/+53beOdfsllnZZwEiEZGy
6xfm1KaHYSBDDFqDKGg+IMmFrhBVP8bkJIWV2dt5CzBFaVNT3FCyCrfBq5rsfwrY
AsLUmO2KXtSmAUhj3rCvF4313CAkApi4T+ctpJNKve8tXJBeXGAbjyRxBPU+Znhd
tHEn27WzsGMcU/b9kbGhEHmcyAvj5WWbgZ+NhcFCV5wLD9PW0kFZqiHU2i6FG4tP
gbQe8tHPWov1kqxI5MgqpjFybK+X8k1Dyl0ZHRwxdDyRJpvuXjdThppozo5B2x7o
yfhoSH3axUbtl6zMG2BkqUgZ6N+cZqcvUWorrO/zKZAriNhWCKvbfZKlkmOxtkmL
fKXAYO394C62HM8RtUGbEnJdyEZZhWbneSWpBX3cfXc8NRWPcoz0Yi6NMJz9FiTX
zYFICMvvS53TAatFmhbaKYMo1jc4zz9FvqDoqlIgSldDfpQMRWgMT8F+ii9OEG0/
Iapimfb7CIdQc8n6jgLPPcugDzpikk6HjWmhUrqmr+xMieg+C7sBdsQRk6WlB9zX
XuPJGGDwTeG1zIJyi6PR5gX5oHGosuvmu4dovXFRlOefndLB5MGpN9xZXkmI6g+0
mRzxPEev9ECYKHjlEB95SsWxf9LtpydylW46/suozBmjIQbjtSqWmmhg17oL40UO
09nk0mINvADAiC1dStQy2DRMbOnQF/Km4PuRF+MS+OIOAB3xLaYF7cT+ePZBe6o0
qzggI+Gm6zCtEnJb4s7Ut/yL0AYlJ4e1ki+nI/FxrIu756dBe+68bYU+x7DeuT/T
72ulanl0ph1hzyvVRTSfSAtD7qx0qS7f6aj95DiZz761t0Dp7jc3XK0hFr5/8y9/
Kg+W8GCNTs+qF3d6yz+0Nzw0qJ7H+xA4yMTLQeCwB38v6OP8waNpOrQC5C3QccT5
8xj6Aq0ltny6Bx0jnvDNo++UyooQouxyVgmaEQ4MmQ8PsQe6HXh46wK+80RosWqR
wAC9snnw9RA9xpU7ERJYog1ki5PJALGbrV1uhRsCOvIdbaVDBBemVQodWM6Ba83Q
vH2sG5IR2/f343maLjdGhPLwLNU5J7KPpdMYqQG+q9fSVfWJIjEQE6ellawMKPF8
yg1fp3mMMzrUySJjsZBwPzIAOP2+BIV9taVph+5KV8vh64po+24KbprHzitdMlzu
ulxZRxY+cErH8fMXv8TGtwuGAecp3jTDwU08Od38i5VP5FTEqIvuYZFdwKsi2b5y
QnpSwYHH89AqGQy3AFNzvBWszfc/Wv/Lr6mOR53tDazg+zuA98QXf/glkCvv1x6e
cuBR7nL2DTITIjdsswX2z6oql9H7c0ayF/6zTbZ/+46k23awqKX/qJtNWgKVDcu/
2NXqrEwbV64CxWMObsKN9W980BXs8IqWtjIOhui5WGpObG8p3yRPsPvYZfzSjBJ2
Q940eTl+4//HgKsFj6Sw9qyEbaNpIv1D1a39DqGzzS/CpGWGJXLf05BvsvV3RdUo
J4O+Cv6mP3EELqZKAXVGoAGT0E4ABLYIuClawXsqor1+DnUEb5X5BfiSuvUZi0tV
whIPheDR04c3L/hT0IcWeADPN/SmIoeyLU0o5Vi+dnvTwPnfWG+LSCsZrJjIW8pJ
wIX8U23ScG74XGKn3AlBk6AYFnisq3WIGJE6IWtzqLiiE0LkY6pn4cfF8Jj1u7F4
R0/Idux5dNu62CHHeEW+MfxkTJDRTUsNa2QxvKls95XBx2gIpF4WsFkJa4ei7VL8
/+pr8TE+0r8XoI8/XXcFkB/QuLqElN7LIdoDTlNGTBvHlceDJAWdNyN6+Bpgqj/1
iOJ2tNk2b5UUJxxOhSqTwfnmZtm3poHgWpvgtTUYbhubPJwFJwZrUYPXz8fYtP2T
huaZYrh4jO6++9ruCd+Y0B/8/hYDgbb0RQ9yam2HdnX9tXIOocXKLdjKFCisw88p
bL9hjuQxbPkaPShluvjBKgP9mxAo4kmeJHG9u9GWnGnvuOjXLyB9xcC18qdeqHQe
gt8prazmEAN2wTEXxNftJpaMh6WJJzXHRYOgCIjlo74MO3h3LqzyiM8IAtuxMzmo
KK83B+CZc4pJUvrsMGmexFeX0ZW+bnZZNmxOJizfsoUSeYciTootKa+fOWx7bLCb
xQlkqmciCX0ZqCfDJDjFtpnxcMzPpITV9yQ8Z+lfP9UZoK4QizaWx9KoF67DR9tt
omZC67hkAwQckTbS6xhBvrJz6bfGfeVt3TLczoFzgjiB9QbQqpV4o1ZTbM44BAQW
gflZt1oO/HlQF9YvyT4dMQ0ccZoUVZj2xN1cfvf4ML2GmOKvqJ2m4o4AA2a4fOsY
0ooib4VXa77RQWLydzNZF2GTdBUPQ7eBjgE/tZvrHFxf9al7hsJEqT/aCxH+ofz9
LVJDdNEei43GQkuT2SJ2tnHQNoOWzxgUxk3lFvrUHbjSfzdS9GDCenQ75dbglvlw
ztlL7/6sj8mAehbSa07bCPztBUDOvgJ9gnizPP60TTmfa2qPdOerMakB/X5yzU45
6U4X6DhEJ1X+CC8P7g4sZBhf3GwaMTX7S023Q4E+nuWQhxgy8o8ibavJFc39yTNM
RK5hscUhvDKr+9qGWcv3KHj+fvEbo2X2lKp7SNLhZI3ZBX+LBxzGvSF8pRe7yH+f
LJlks3+P4qA/AxpSzyBjZbK2yaZzTkWUfeYWg3ntnFWzaQ2kB/C8Am/ulp6KqDLl
4DPdwMFCLzIsmfCoZKCE0z4nhB/iKVWwn29pKsgXeughfjtQHXVRXw5Dk3AT0+8c
irVNlmv7c/EU24Ydk9owepFEPngbsKvUk9wl/Trb9FY5djJtS55HljxjXZlxyjXP
KXLkjq4elz3Npo62NbUvptJCUlN5jIlliZQ3xxg29yOzzyO1teKujlrvYCKxSENb
cOxDfcV4N3HbL+WtotEc8fjdk8GUddIYpBsLxASTmfwRzJuAzQc5yMBUkyQrVP7o
0xxw1zBcj24/Ria9NlQnObZu+p0Nc508XC8Pzb/3VfOYp4KCcrVt6YhgKfacknlO
zUOv/klRb3L6+lh1JSUZjj6ZJaz9uykD/fwItbrukeclugAx1AVJ4tzV/XIjSTyJ
AOd7NBnsvPa7SSURN8nzQwZ7xh7XTYduraY8z4xLwZEVEfu5bHhhx4+g+dmVqJzx
2KhU7EgEE3nq7GTdWk9kmqNgK0mccbn1iWau/e6M1xDE5Gn78BBGYUYRyr+yKKOo
CgjEqnUlnOTew9f3YuGeezSLE8oKH4lPmgdXSqT2+U3dqdJwOlkMe1Yk2Jp2kSq1
UymzwK3SSXQiY/pn4JNOgooLYL9GVXN6wFgVtTwpzRXVbCZxiNJlyvLEWRj4tYN/
mIbWQ14jp8XILKfRkp/s6X10iCVHQyb35WWxh4kdL2mDrHUB+qJCBY5Y6L5Dfc5x
Za3shNvutaAV2/FbspAsc19aqjtRKLGQrsLEjhanenr61vSkWG7wLVOT3nrZ5PMf
CbJhj4kzvH0POHao7ZL2epSZNlSZ5i1eAeL0qCXlbF2vMUt8fpAJLnfxPlCko9vD
k+DcEavHTAEAhKv6o5KGSVb5BWQIAiP3GbyOMKvm9Tk4Li3ALC9o6EgcISX4qyCS
lUhoIOkf2VJC+J4RDJpyJwlzDqi0BSQ9fw+NqeoR5k9o+ykjTHzv2zxaMq/PDJpD
w+4a5QnT9kDEXGScBGpeGx/ncUEsdDj8kyH1bCHtaOwG5GaAOuU2d7XVRPIUfrCZ
MytTPw/6aytORAp6hQ65XgwcuDCDBOjbxzxEfk1FfOCedlkLPERGH+nXS381RVqk
MpzlYWdJl7mrr+8GvuCmLM3lHYbkKhqM/eh3/aeIegvBUemxGIFckHwvkOij2rtK
EBzNnfeL63k7FFwUplSjUpb6ne9FjZ2k5twLgjd86jcx88u75cSVoJ9NdH/NhCIZ
8gax3/QKTuQBYwM6LeEQTk2wos2z71teFAGkMaiER4FsFZ/RBjTmJhrNj2ow1Dcm
Nchx7Vu5MKSnbD8AkZzXz7s9i0YxbmCTRKZlYx+7+HqHDOTH3oTPFF87WGlGuVwB
M+RCAhyYsEOdTdxtYvTJHm+v3x2bDOzzMWDSNrqrUPQXqCurUAzWiHCTunFPGGUg
PRf/KwG/OJcrtIfdT/eKD2LnJZ0erw0v+vaJw95S/LsFJ2DuKZlTXFsSizIfanY4
ewqPbsOzMlCwvwNAvsws8cSB/Z3w2VbmgayzNcwJnYS+6twz+0zhT4WFcrxXRdTu
V2w03la3INEfdVr0ZeSG/WUcvj5hcuN1fM2m5T3UpjhhazaOkeUrrMebGjFJ3pg3
Uo+0lJg2TwYF2iiGnzsMPFlF1O2lZcPPr30CsxEN/sYDm9Ucmn3VA/PuJ3K+cELq
ph8A1mTrRdv09t5LMkDxqgxEU7ingv29fMnFtctPzjnub/0ks8MQNfgtT2bwAeym
MkJqbNkI+KmzRhzpbVKYJZIOwPxhFT7R6JzF5xUd2Wl/ktmPGtFNF5deOmDWue7T
Vzi6k1918Yxpj1uzYxGnQtQ0gL3lJ4gqG3+VjgKzkAKddkmhj4+AOOcwfv+qbjzn
qKw7LbVraaAo0MEc7UXwpqXo5mxYzfYmtWqk0C6Plz87posLbR/j3umLpa5t3UQu
TCeRoj6Ll9HCpKLaQJVk3y8bv9uU7msU36sM39l3H48b5YLzhv1q6OvtikbdGzQz
SJR/MPErNPPAaRN9y2xousvNvVPOf/6XSQkZ63GPPBctXg8S9UZBmfh4/8B6SNR5
gQRS4crHFUFz5Bt6W0+8uWNIr+waGgcSDToNW56ECtrg6iOYsgdkj0xVTcqCvRQn
nwIvF3Y62Y45jdWmI3JfXuhHRyHl5nJLQS/ug/eJ36MxVsckwPLGQ4HGn64R3Ecm
mL01KCGUD9jVih0Qmt7zGzkBAF5djFEtULrHqasTmxLgZelxyS6b9UivPqaekkqh
ZnJuP3Saw90AkG4PADasR7BrxTg4HE3/oVtYdU5HqGHDEw612mC1joVh5N3ojaXA
GsEaAz6k+RUFDPCuhB5Rjow/MQTI5BPVQCIBNLL9ENDBlUzVdwytJdscT9lpBidW
Wz0oS7urWZei65PPKBZvrhDY2d5htIuIp7LuMHZEeuMTWK9qAcgLe/fOdPZ+FwvY
WVuYRYzRJcfaWwW/bIRCuapM+Y/omSfnaqJ2uxopH4Ur8joGqoUNEsBgtY3PuAOU
r2JxbEMTOfnm/F5kY+tzilAebWBZ3Z/DDwIqR4tRdaTHcG6gtFO5kCY9HLpWmgSv
FFIED0r7N9ptzBKsG4zklTfY2LPikt6vDdtm6NIHRMRMsLnlJ9Y2/m40GyVtmdyU
luxsQtCNF8ki3WtnqN4E/W63xtZyS5QAEKrqFaUUhLeDfl6yzE90wmo0iIQYMuof
McOGCuPSJr+DK5ywDAJDqiomYSDRNtrnJDYKLvkKmRrCuHKbYJTr1/gayfNfTgHu
C7+Xu9K7lEpMVwBWFh26R4OqPKWm5oBftZFKdnm6a6AADpIpywcSYwSdOBsXp3W2
eLYgNJTdCBVEjtMIQBIJIRDpdma50bSiq91zcrszTU1limIY6+v9Pkl30Ou85QKH
prnxBZLP2JRzOhoECbAsRtXXVKHs+DCDDlDyIqfnMqGaFLZxAbzHq4zHG75Z24zC
zbb5+DZXLBq6psORwgbxbjvnERP7dtYSy4W9tGWwOPhiCqtMyr4+NgPLzczkKqZk
HognbCpmANWj7g8aW9K05SlVPAlvNTMdNhyDPqOIKxuYjE1zMFDZcAOFbB1PhjcK
+maFje+eyEkZmkCssgQDxOdvq9uIJQYJ8q7UkSlzfYB5689IGSx46FXoHz1fHHMu
20OiEjGO+YrmFuNDXvY1EOqhfGBpXWIGUoUF5UaInqt85qT+qTAO8Lu/5TsvvlUv
3Dw3rAofGEer6faPVboaMvH+WTn+Y/qtrmyCINmdNFE9MG+kRjhKBlkdjkgAIe7x
a8ncVXjgIp9Wp0X9qXq0HrViheSC7HOwkVELQTuzb7uyTxifRI1JzLRbvFXSPM2S
+IJzK2McVnY0U6KXFwLbz1JQgDRsFZwcdneuuYmViwgJ6CRTZ7PRSC180fJ7aytU
locoExeNuflR2mTFTN2wK20tAQqSYE/GldCd/5MYrH9X4C+UtAIxLoTpc76M7yXV
Nhx9R0qWnSMCXZPYGGPq2z0a00CrZgkudfkRaQLK9M3CMa6SlVTn6ovHoaJqYPsf
BrHy7N1WbS2JlOo0WN0pPbnxnEfD7jUoNkTUD1uWqTucJAZiiQtHCNEqFasemCUQ
JecvXMfu/qvY69DSnyPo/5iurR1IeQvoEysEecwnlJJCDyYRxfgOzacMbGT1xhJW
ivnuTF83N173YVi8yItBJ/3x+GQbZoY1iuqFJMu96vo3/uYX3QR1PpzATsSfoTer
cYjklV5GYisU5C4ZpjxgohGqKoQreVjQr7I9rr2HElWJYKiC9oFcYYrAi9zU1mUv
VVUaM+Yt9YD0ZwfLm9bZKmRKdkUQruEzxR0WlW5AJDTVLL/ARWYCMlv6qGOxFvJf
qwPDxc9BjFePn/70WdW8wcPqlTgUyZN2RERR+r6yQqurCCuMfRPOmYBPpQVWB0o2
5ZwBZy9epxhdo34+TN7snVvskaqZc6G2YnL2bBPSLYo97tXyhqHt78OJ+IPlxmGs
wsqFUbNBeLecMBzFZNj8ras41PmvEJNafYg69WP3ZUSzS3W8iQaUjK/+ZjeYUAuE
wwJWAvdYCyoRZtiC7wzATky3plL3LAkVXCAQdG8j94hS+Rs6AaUy+6Z0F2SVCUvr
PPBvGfD5jMfjVA5QC8+XIJWJpJmH/sYDfRVRjhUPNzamh75ZEwA4Xlps93p27+JL
ReBjTS4y7BChNw9b2ZYWB9441VHV090a0zwCnYriZ4RQ413agXkSUBmzPk77E3bN
M0z+Ek9Y+W5Gw68VE1UEgFhH3OD7WLlLxQwkOOuI5V/o+EdK9EwCXTICdmHLgYzC
FeuEiJBdhQXH3SXMH2ybC7aO1PUC8XMNhAaVa40tg9llHhA6M7hE4FINcvwobsT/
isSGVNzZkhBCvrDK55NI18dGxaS/vps+VNjPWaeecpRP4o2AalQUQSS1Al099evM
s3/tvt7AIsxCUb/cMEwhF0kugS35b8LFXZaw6dk46ol5ZdzUka6FOcYxaZTjtgtI
ZGTtNcqn2N3CEvANVCigAhGsS4yYmVCrtCtH0+Z9ZFkEsM34ATnjpNR+oLJYxqaV
cWogalVkCZ5Hi+/Ae1QisdOJc/P/L5nOz+ijgxROUSQxl886XOtx7ZKXVNJ7sNzX
CyT68EbBycfbVH4aI6e/7q51z4552R2uAafC1pbfPk2x6fhtKZNcBEvHCnmK7Pi+
kilQKZ0h+k8M5jGTWijbz8xoFFZGqFn+ZhQHwdQ4RB9UPWnvAZH6OKZQH/Jx3NFv
3bp4oDhOdmJ2LUNeUdTj28V+m6HnFYokNUZd53NoF8ES8OyJiezaNBoqpQVGSAAM
9Nvz2ZaBHmVm4O3G/UoIFU4i7ujtM14P9l/cJz2rwjKRuvfhQ21jZHmxzKzffJuk
GZA5mBtjEWmopvJFJM4A2XqOc+8seROUJPIVrwnKTcBlo6HFQg81Ep6I1AFU0O8H
mhIefQWk2AvyxtjTA1/a0Z7RNi5B5pxVH41XVUyWYCS71nKz4j4eSrZ9NwswdEiF
+zrs5E8T9KtCXrdlESpcanBhh2jSN3Dc4aoO/JVldYkXXM4kD8J61v5RdH/+p1AG
mouvDF8rOovYvg6TK4w5zJg5WD4b3I8LIcWJ11QFQcYRJh7t8QOhLOv70Jf75tL3
TTj3ADVZhrejIdZVZSKZX7js6LAVFWFGBjagGNICIaomPhTHSljLcnLA2hP/92q6
5K0WJnfgjkq/C/4ut8r7vmmL8pbmYKapBnzWZvjKNDAad3hTVt+ZbAP3nJ1xdkQJ
7Gv4lnQSCsvFc89bd6poOnP2RTUHg9NNmE62B8titazVeDWLppHv2/d5Bl1GH7mc
BpzmTE+sKhfUrQ2AbTJr8p+GkL2jWL1ldwq3j0AwGTx1HzecuM/DHiqtN8XD8cQ5
SYRTzR6h7pBGcgi1y2IMeJ+4+Qe1TVZMd6kjdD9dyvIG5Xc6WxIbzfTqJ4I1gVUn
iTnk17bJnNxDHp35+sO26pcBrt2TmVl4tpDVViiuYfo94G6F++OV97cotWZs55m0
7NRKGCoOgaHCixy+wv4OYwxnEgjKS6+jKfPwp6MD7lebM108A4Iq79JkPwaUdHWb
6s+yu702vuaWqnphUr2HqT/2YLtkGhKbR8lbho/8HvH9nGm7qhA2OSbbdbsMyF91
+lHUfR/DqwModtEUuJJEsO9e5UpPjTU5eJ5/XaR5DD7Fai59QW2wCkp1RxhobIfK
59ovYwIeYFdwqEaKopDCHa3qM3usZq+k7eR/M3XjZ0sSqLUmHiV5jwLvLwwoqguO
G2cU8KOqgmJCNZrJkMo5UnXcUI/tZRCY/uS12ipcy4V3Vmz6Ik5+NEhrL132KZtu
Zw89t3AZcpqxzKARBva4azDZWEM7A0vEzry+y6epIsBDd0xds5wUhetTHGKUpNTX
FRGmo9cqsCD8YMGxZIUoZ1NrWGMNamjl7MDA1I4L9XQLZ9bb0mrt9eoOLWvhV6GE
oo/Wk6RZEXtZm9anI7m0u8UxMOYH4qc1AsFz1jp6x2ygifb9DDCUdF40sBVHzX8F
huItFFB3mO/gHAXWA3WlENul+zFblEnhbThDcxehyBmyhdima3d8KXuRDw8CEg8i
1E96YsSy0VSP93jGvHwQ5jHWCsqTP1+No077gDG+nmsEhasfOWyqM68LK+JFcjRq
BsOL+kI1+9qGRufW5RgDqFCdkzA54sJG9IoBapJkTDHYgbGKWXYCKFk7ROzMFF8H
ExoaxSlpK0LKnWcHR99mqrZU0eWJUB4Ng24Y8lNvS6aWtzgQL6CYaYRZz5on3vgb
5NWkFHpLyu938pJLL6YNcV1vR5OzxAK6jQ+dUIoQFHyNNMCGMqsq3c3rlRggk1CZ
2z8Taqdon7nK8XVccimfB/7CijA5SYzyU20j/Kzvv7GIY0iMCsBviLmKG+m4KYYO
C8UVVwSXeT95WN+WQ+M0ELKdmqIr15nsd3ziKhl+Hz3pmysLpRL6bvKqn4pZ+h/a
0sXTiyHDlHr/ex+4tmruAtEXrv1ammlJUUzYw8lJHk1MLrP2j06lqYz687V+Tezq
18K/iHDnjuUdAzkUgqdVh9S1h9xwYSCSiPJrWNXxsmKIcKBmVtHz5CF2j6VNMNFp
Gg7RXO6Hp35d9daexmMDUXshFwfCNb7QS2OPA7B8Q12wPFs0DNJO2rhX9M8LTkdh
p+kFUpOZ8QJwvcVH6Q7C1n+DR2TLe1qhAYz3OeQteSdQeR8QdcwLWRczmvIrRL0W
ahI1WOLvk5tHxoZ66LnRiI1h431hTYSq4unaVkHRGYLRw8+zhSPJNeX3+k9Z3mR2
ClSNHh5LNy2xFWULQ4HjZ4FKIkYsyiin0J0hXUP8Nc4QhPi7jvokAUJpYTtuFOF+
6vIGldDPdP08ugqORLJeAf7yIsAc4UCLu+jZJj/IqY3uBzOCplIqk/JNOeqzsZ7T
g2JAvJox9t45VhIEiLSjOoDYasz+inQUaf4Xv+SXR462ZrW3PQxG21SqDfn05cIS
8PcB92++qARX3gpWvhG92ah/q7NZ1HssDRiwBW7Sal+8T6GYsDiL1gP4Gt3DNSnv
dd/IXK48GoApbmANiFO/RviK4sdIJ7Z5zlmcsUrUgrGRuf9uNaa20Y2VCxoRPEI2
TNrU8QN19HyW9WThyXDWmXoV7ibasSjGg1MvrlpFjOZXBwcjT6Ht6Oq1djTZBEqA
o7F/Zm7llF9HOE2MORjH0Gqn18fo6PZ0twH2lYmo/EpXJ3WFMCtCl6QvV1UqJxvr
HgsZQqdquL8VEsYjfnPcKlXzZS5QWppfEng3QzfEa0QZD9ndTcewRrLisu+r6GhJ
sZaksJNy2vJTXAJODyJtX6M9Ebw62kgyxc29hhK5lOBMihFGYLHUt2/lheNg1lhV
KbyyzkcHkrzbVWDawBLRugSEiZlEiRm3yAdmLQofP2PuhZ2brpGO+JafnzWQxspB
kKS03ANaG1kYJXsvHGU3AdOaQK8Z1hKTe9i701LUr1YSrWywf2NBIABtEKzXuxbe
cmaUSNXgBdz8XtNM0lDXQG5NALtJJFx0qEIy7i83IW6NA7IzTkS6FT+mGlCwPAJS
c82B4FEGY1PiRuz8ZfS5Jqx6kENftDdm/Ts2J28ayY4U7Nm3MzRHH3TwkTRfVqtP
EhXDzCb+qx4MjvoRnz5xlCL/A25Da4VBL863MpS+7G6Jtre1i8b42iF2R2zAmGW8
Lt8RWUzwAd6cDdKSiar3J93LIEBB2XpVSTqhvSu4u2zPIrqtPXcF2+IVm1sXE2ri
Z+z+itWZIi2mpscTuVRr+OdZA4tQmGsGSCEE7RQmRF4jM7QpSkucCfKAL5P8m7ym
np8AdRX1BP7xrCUkkoy4+pA55hsXcVgJh3AYoEBnWZ7U+nAR1i1DeZBW+W54+Pt/
2gaHSoi8/XK0UKECoTFph+iqIkoKi27mvqszbAgqn48HjNEGwQrZn+IJbsEqIINE
6vNjVrZaSDoqp3QCJxaTZ1c+S1RS4K2rPre2fa2vtlZFrjTbS+gfq3VMu4E0SFmF
QcBAee4MDV7CBm9xhLiQTJ+fCXlOiA0etr96JenUOqEBOjZOUadKA6GvOxkutL+g
9uv3PPnIC0QtXs4vMPzCTv8Z8bl8bmNAPeOlrgXxOuiiamUQS59r6faJadz9L1F8
82BjKmfWwpcGwSqo157kmLG/HOrF7Zb5+tSiUA9WEvi8ht8RE1ChD0Z8g3ArO+Ho
pgYDN0qw8Ia/DFe6nddK9X/OMDLRe2FZI4QfQGWLiV82yE+FL3iHtQRkD8KhVW1d
gXdLVYiFWgNrUW4P+aJ8FIuF71ysy0eCWkN7nAMHWsfhw8ezdvbYvE0HEtRCH4/F
CfGd29spsj/KHwhORolQQpahm26O6rulCviskuw1FMJVG0NzpSjeHaa1AWkuALT6
tWkhHGP9wyPp6vR6MBIWJW8eWNczMy89inaNqjINyt780unU2ParUq+bJdfQuaOw
2XxDln60cw6AEtRUEhIhWX5a2heNIldzn/Ylc8drPDKnD1F5VW+xa0zhr4Y9I3JN
YG32oXNfLiusZtU198tE9yxDv5ZLgNBdFnGJrjdYL82bw9QiV1GY/UUemaX7KuIc
J4I7r0QTYeER5o8mO1GO2A5VxnjAFmh7CrY6bjvbMsJJ4Df4Xb3nE6wTASfyeDbK
nfRPPDQK2Vi1yGeyJisuVvVVfNffjGnBY5HPxxXoFF/ug56tVsVYRN2u0kOK9HaU
XNL/tKOp6G/LNv3snJ77R93ffWeSGgh5LXft/LhC6bSII1qIkGS/LEVoxOX6uanV
XIEmrIyjc2t5V0cDKGYdjEWxhLROWDCDN5DnPFFocwwi/GGRrugZpn45tPK9RuJk
rHT7QmPDmTSHMlegd2HRSQobl9OO08qtv6F0Py9ip69mGhtmubQZ66+4LfwUlH02
YhGlCsF7azmsSAS1Nx1bN6BFM2jc20i6A+Vd9T94Tpn8niUFe98oVBIpNl2lWDMS
FhVYsIvddrP2D/HMHD/L/v51xiK7PGay7fp2ddywz9l+fp9jC1gXTttmn0jsevi2
6RwI++VyRt7b0kKQElgpBMXIFexcqLHhCUXKpxdJCbgwQfWhm2ao/0FW7b5nLb/L
EGL2ANWYF5Ycih2eAGpP4IRtqpg8vnN2myZnQpgYTZk3JMgCT2ngg93d0Zij1lbl
JKVu3K51QgKWDzXAQLBKwwBf/wymthnUuU3ML7PCC/NSL6c8Tq+j40TtspoiP5t4
uQZTj68wjWKMmdh1rxyDvzeh9HcdzVNOslxos7nqaTuJ3HXryoxfdy6PmiEvuRMM
1Wip3n9jCeiAhKmguxATtaVrP30MyvZyZgu1DzwVf3ciJt1ypiBSyytcLob1hDhR
04zLMzEEj1UYbQ/psDhtIT6zdvz7KlNMvSNwQJHpFTz/XSjDc/9hs/P+Iklm04EF
u+5n4kQLCkzSaIp32BsSNPEgb2b2BsyK1tqSLXWBqGMNpIsvpeNpTssSLl8344C+
IrBascT/gCr1KwF7xF8UDShkbPuM+DHVUpsFpCpIb3kvPHtYKwZA6sjoYWAOe9jk
6gdu6Bz2jgUTmzOmlG6BVYO1ffSBBk2aMgTx6vWlF6VC6P3lIdyHoYoV8JIuVSD2
Iv6AwBqm/p3zuVr6dx8sW9jbc8MKpxUX8VopY+fJlhGoNmB9Y0LB7zekvEwtN7Ep
62d+LsMe/RegZ3YflDR7nDsWTBjmxYcloWBvrD4IUDk6k3WLBy36R46XZ7jFHXKV
lDEEkCUyJ1Jx0KUK/Pxk9SaAsScHsznbJ8XF1Dh94UykeQi8VgWUa6Jpbsl7IrgG
nWdiHgyh9KZkjGhEUCfh3ncsym2ZtT7goyhEBaTnpPDbBQanVwy6QEQ7TVfko6OA
tMpkAf/U5H4xcYJevjsTtdm06SZb4I97fCJknoRzAwLWraif+bLkr3+KmO9ISwne
oV1Vmu074aH5KtXVneIZ1fyz1aX+mMNm29p6h2Bd9VJkuo00N9CjG5/RD4o4l5sc
g66V4FyOIUlEbf1C9xOKNrZBudJ/yKyhoOSUe4jyD8euHTFH0xPXaRD8c/r5Zree
0c4prK/tX/wLGrjl8byEOwdw4iUISmtCNiHW4+VUWWIUEpCcnBpJDZmfEAbumUJ8
eP2gIE9sdTQUSRnq/5FFBoFcvTp6+aJj1WHI0dmOAkVss8HoHwh0Fdfj48KO1P8v
2KpLFyIhV/q069t5GvC7QV4tAv0Xv6vrmv/rk5tHmTwUSaSilxQXUaJsgrVn5MIE
ZpXqRFCq6FgctNRLw8uv3yMhW+cNtPpZ/rICwlhkvFOCxveFhh5uEMCdr8vO1dYH
YNJQaeCHi2Q/6ZZ2vW6Qn17YImzqGNvqhvnfrL6SKxQnhqERcNk94imrJ3+q2dnP
13qLtKLuaGRWQgt8xvGCYb0CGqYAbfifZU62SuyaRUtRIPPJose48pQDSl/uLUM4
T+5Xra863oZIymlM6qzpsc82ghXCD+nBBTJm61pO3lKrOUFlYIHHhGstm3WosajB
Mpd4lmm/xncI5BiMw5rMQw5E1N+KLdAZW3wJfCAzkXInnr/hyLDXKW03iPpL/5uy
WXu3wYUOkw6JBjD7Pt042ACGiASSEd1k6tO8dRwevjy/0nK2AjJBot1ovDp1+xVU
u9tJ0YgkLubPFxCM55hFLKJ3hBRnfhIXJNwS8AMMf2TT1t0e+rNxa/CH6tgbZRlP
1wuD4zVS0IchOCIdcU5vkgGv4ZJCj9KYcMPXoJ/1IMmIHlPBx6XV/tNQTChyZWTg
SxQYkWL5hsL7eMAkYCmWhuNQrIVlvk7pGLjOFsxhLTqOvVX+1TbywPKf6qGNj48I
kGty+OWIHaDUs+Kar8qSk2CIKAKlXT59iilUJh9POoQI1iqXAhc6QAh3DUWfTrnB
e5jGpYCUc+x1Ueik4cfOISMS77Gd9c1ARznXPPQ8gO06soGylI3rDQOfcA38rp+a
zpCeyJvEM24+KVUzscyi1pRMyZZ9OTJcbl4QgsYP/NWQooC+vDwQS7JTKKBS9fbf
vTcZ7+ocmBWY+bEjg/2Ca62e0RJ8KnzdrnF0jh3cBHyJIPy8/xTMLOqvWrGjt5ya
5aLt+4wYmWzKvnSWejXYtjwvqJxk8JcqVRpEtMh/d22u3hBqdjtRqzerxba3wCRB
MwwilvLqs6OtcJuGfDiHy2+hOsIossi6irbMwyU1Vz6HvdIa1xgl6MwxMaenKH2p
KS1H+ckyih3Vy1wEftVEJcDG2pO68OfqL6GxMXTbhRJNDZqnYuJuWj0vRkXiT0yV
oH2pjCh+xSjpa/Hk6g3sO3lGeCV2XXdwyZRLw+qAeWWnhU88j63xLmtLQQZ9Yjjy
I5qMvxkfwdg4g9y4F4+fPaLwEnBIhtGeD3f2G1wvhKwQh/gtmx712XNnf/8AeGFn
kHimBLtz9Xna0N8qAk8mE68xzSvaEZjcqr3AN7SiT36HkVsbV2sTEXKx9hu4jir4
mI0jygiao0AaoydBH181uN8yf+QSHFJjfTuoB0taCk2gz+9hKM0sOfWXfgoOQZYG
q2i/6Fkq/hjdynwgy5VioXdC1DhC8XYeBzh4WwRRJ+rGkrLm5egO/fo8jlpKR8fV
JDtAlo0LNt3Fop1cTCuDvklAk4aafPKmodOA9Yatk+/U8ukVrK5q8CTGkrJRF618
+ul9L3SYbMquwCeJjiXanNmIbj/9xuPJwHQ3ny9c8LsJce46jOGu07SbkTyz15yY
xC3bRaGVIPt3UKEX9GawO+UGizcAAlb7FjrgodPMlOKKO3PC8eGv1ZlWxMKNvXoG
BRyUHII4/PrvzncMe5l3GQhp6tHOhCXrP4+oHZEQXTCiEG/d6g3qTO/F/tbgkX+c
0KSyPM1DrlZzIlVWV5rMeIbvrnROdTK3zAckWG+AK2DzqdM5QkGBej6ayfyZOdVx
qeUo9ho56t0QGTpuTauKdNu8Bs40a63uAqeVtM4UuWlGanspAP1IYsnj+z5NcFGW
2YztpJeAnj9rB/vEkd/Zke7oKkPYxcbl3KLusFF3Suh9gKfISiNFU3YOz7XscLy7
m/DbRrf5SwyhGw3EDxtPNSEUHJGUokBDGXKaqbk3p+h+W9g91gJuKdgNj6QcKuuJ
fC2fGmvgogSdMEw6S4xDxLYw3L2pE4sVE2b1vmxyVwhrz+8SBXMKkFw9LhRCCEpv
iWOLWL9k+1I2nO/Lbcc2ADfHc0U632tTqOTuQJKh1ESHbN5wMHRJnzkcE1bD6YFX
2SHR6Ojoy4hT8K5dz9wFw1zAKqIwV99y2tCT8Pzj9d+EjfaS4pzyMolpLC8hUaRY
iacF5cAQYlEiacygtemdMGrBZ3lNmGxV7ooSkHu8+n44S3p3/q+12pX9HtWDDZY/
+GXp4YvIaQYCTqdOrDyE0jVDd/Wczv6aSvjWLWpmWSmwLhnMH1GK+hckcQxiWwxq
drtW4/HC8UR00RruhtYVa1gfL1SjcBMWD6zDMEflBWWgPgjSnpvvg7J9z+FfR6tA
7xZ2BAu5th3Ofj9gHVo646h+JSEVNNaZYt2rnGB9Q281avOh2ykbj5rUF7MhuZGH
J+ykje0XyLWoDArQAbgpMFeYnSKhSVCYYiF1gi5WAEl9AUOnvVlsfdEqcKexuyit
7cOitRKPH1JVEsXkOlpTeAH5Bm/EQT1GVBPuhYzYtXXSdwpHyO+WZSQqiyXQJZjb
uexnSTr926NYqZ6JgRoreuhQTeHs0c0tPZZm1UelAgk15T7h+ILz3c72J5SZPmth
owhbYoys0xq6UHNLHi7u9AqRmWG51ZVGSRQwJS2m0+zt6GbRxMDXmsoKVpe3tWXg
jT5dFAj71tzRG7aGOhcsqJrRkMgNcvi0mvzShhJ0ds9R2eQBeuHminwBaEQjRJx6
t9kqsrSgVOOhQ3+X9UuJlDXB+iGy+U6maD2x3qB4v6kR1gIJiK3fY0LZBdKplOUj
dnMsBdX0iRZlQ9NhfzlaPTATEgaySkQP4Ee43w8G5jV9GUGspokJSs0wNqjmVTxy
NMEswULB0RwIj0CW5a+pYRJbUIrh5BBcuE+OD/Jrj9GcPBqIqbh9QO4HgbqEf5RS
HegLdRHDR7w1bNl7QZL/FjFrVvVWI7RAQvohPNLQ8FeXIQsd5iscmt5QC5tzOMkF
1Y5bU2chzy4canfdEAkFFTTLbbqK1Bj3MXB84+TGDSVO/R3CmPe6zRCU3EiLj5UX
tJGISf1TWSft2Fgx/yhH4iuunkBG7Knv9giqlyU5OFPa51bcK6xq4YPVz/IsfAvo
IzPQnjHz7oCy5OIkecPjZYGPadxfDJ5AIIJmFSMCVGx/Ax/eJ59KBHSKz0uD+Hhv
vv5YZ558VNnpo/eeWmkWJ9egMFL6B31SgKPefY1D7DT1SWiewC0j8xaEO5VA0dIu
7fbOE242Eil0cxwxkQa/lju/AI5EvvMzcuLrAqKoVgo65ClSgEcxafqByfdrqAtR
8VTooExzhVvd6q2skuMLYhUVuPSg3Rq9M+8Bmrvgw0ai4hwwPOizO0a1Rbsho3TR
Dta1/Fr3URXE/ZtHJ8BrCHqVpovs6ot0AfibyCcHWzv58TKzD9b87hSH21lMqVeh
kYwkT3q08WTxgnBNLs7RmcnkyDH5LT2JKjZavIQfPDM1k0BcwlNGnua7ddGRdVVS
FtcBneDspCCf+A0PS3khaFEn0kb+Q844lT9QpUwa96pnSySiWREtrrbS6w3vQb6I
7TYdqUi+xnW2O0VrvKzc6G5svHWfEw0z7k3ovw2IALqjD987JfPpfJGBrsdYo4TR
Dn3duWdmeWzr+7ZMJaxuU33YHRR48UEpZ7VTbNk1fcuLeDPy13jvtRoF0C4AD7Hb
YMZPU/wvEPAuKFDibp/NXrMdrWLTXaYQSSsWVIFDkfxyu73ugYNvPitr5RXYqYg0
pCCEViTQV7ttUf3koyv8tevDdWW0jx8w+4JtrnXbkUOYUvBrfbJNq1v/MjV2cwFX
ilWgMFTHT11F0FOo8qCqdB7mpamGs6ozZcjFmFWS1r14Po4AzsJZGBvkI7wT15FI
o5zAD3zh94/uhF3klg5rcY+4RoqFQrZmsDz6EO4TOHkjvKM0+gE7lXkG4V3Cl9Ev
95EyZgVIL+r1O5GgkeaskMXn+EJvqDk877cUPKSZsGaDxF4eBElBzE4vIWy84UwC
kjw9QR4auDgpM51HHgz5paBmmMc+rvuEV6wDBjwZ/gvafT+TDm2BBhym64p3YuXR
XILo5z0FDFnOmWisnFMg39UBYPdlFen23+BsWTdGJIOC5E8Aqlu9X9UfRMmx4K44
Vm6Ptnf7gLu/KUO/cOj2MeU3/gMeH21kuBx9umf+nuTO/aLUsfPaw8iZ+rJWkkwz
PklxLVADzk60eCQ09JK8FBr38DTEDzWnbE54/r7EMJEkXok6/euq5fBFqELnN2xk
X+scaqWEfSm93vNeXFJeGkVXNfP9MAolbIsyOLmxrw1vh0jJ0KqQY4bBJf36dPEk
/rkQpAQjwoARGqwX/CmW7RBd8mFvEQxEraGh4gc/HGc2a0y0RgSY3KlR6nYIKakA
6oqVHCm6CZ2slJE0outXkpMA0ocBSXKoENw/rPZZpHsHDx1U5zPYieArZjNRvKy+
HkF7nFvERMaoya3HvMbGHKYwzIIs3pCaOnX3U6AaZLzdvWQV4AU1Y257SgdvMASz
u3VMaFUdAieqEQquNMwze1/Ii3vjty9DMNaUfueSDeP2ORqMskt1Z8Qq0J0I9dds
KHtI3D3COAT4gOWpeMtcZdMDzeR07Ccbx5ZNTMmppw6p8fqLdFoTA4alHjtp5YN5
1SLWozcF4xWQyekR3rI2jfkZBe86BZOoC/oMYgzkvLfaX5txey68nXmvenfphUaf
K2bf6NImm34hfz3b8YcQwOEYgrLu2aBhloctITq8LoDFYWBjs48UgldXLnc98Jyl
ecx6Q4NRAAqnIccRVWecKSq0AdUW9b/USCF6eowa6H9JjVo72leUYhMOQIHJNQW5
I7/cYTwOLqwHafZk6pnslwPN06Weh1BqDZ63g+7Hb6OizrZgRlULe5AAyXV/Xj77
f+6JZLB3/+WqyvJ3x4jjuar+joxa0Fi1NkzPhpILM9FFjDrjmpuQhQv2GE3vi45Q
rgybPLdL4UtdPTohjSGIMtbZuxLoTxKc1+W59Df7BuM2DmncNzLZzpmDLkb9IE9a
56pLalfUBV5pTl/D5rp01E5kYFT1jkGQC2TPfiDi8IUI9rwRsKtRhO5py3nvpnk7
IOM6+8iDzTumXm8bUuRV6CN+zaeBqDKY+YbPIhIkRbB2BCZDttIrNgIVzrozB0QC
V+aEluVgzDygU5NNMCD2Rz/l+8oPsd6XdMpKtgMnklCpj/0FPRjLXYUPxErUNU1X
+D9BKEEaLbDksthaVVRXigViG30hnD4dnqZkfyMn+TCBdF8u+zQ2UqazvACNim3n
xDmGAmIEjivRouYELZDoVQK1LuTkdLJ8xN6aXaH89BjjT6N8sCJOCBv4BQ9fA6qo
EmLj7ZlNJ4CgW7HNjpwopkjoFOV9tbQnxEF8M/InAiOVZwoPty2YRxAx2YALkpY3
LzjfTbU29p1dF+Prrl9i1ml30CI+EGqAxkkga8hDPnKKUbDjfk6zFy+umJ5mfZc9
UQB2hqfzCvz0Zl4xREKfXzNvbfhtdrc2Yg/Ygs1DLu0qiCQFVX4Q3+5ecthWkTdk
yd4Z/qKWxI6imk2p2U7XSHsY3KumwklWMERXuJHupBaVBXm8Q+4mW8QcI9mCvSPq
kHZ44/n6JtBZSrtJ+aCbjLivfSvbdBd4dbLnZVbNCnPOA5fW7b3n/O13CSMyckrE
De2pjIGaRA6s5jr5KlunyiNDSIqruDQN7Lq9iifrz4nQYajO1kN+MsQ4PlSdN4H8
D7kPxxb8dfAgBqaYlrLxMc/E3rFzpI1zhpAt+zkhy8U+UyW9dORgYmG0kTiZRiPw
0c2HSXJhXBWHaZQ0lPPQvNBnQ1GbrksuBnBsIiOLE6k+jGpEcL6Kl8FOgge9VTij
bSG8ix8mGvVMx0u23s3wVCRw6g6PF7GB0znTCT/j1TV2kb5Is1qN4jgwJ+cDFdES
kieAmKqrO8d7VCuqHrjb2Ki7Zc7uH39Ql5PsoITFfN1ziKResDSS/Iorduy53lPa
/fShuq5nIbCQ/5JopsFpadD7dh6L/kI8mfr4HwVkQJCB5kcXXVbGiPWu6RiOWd9I
ojoHB1SXYGZ/rge8U6rWLcrJLXAmookDM7N+dbKPyU5lLGeh3Mp1Rf+nZZPoMVyp
YdJypNP8hQGlspOwYSlVTN06sMRQ3nSoA2xJudOx4r8Dsz3H5leMsUD/vu0ljhTy
bAXY/Mh4coG7rNv7QlaoGsaGzRWRa6ylaDKoD+h68VfhGxSupb3eOe9JlwkcsoUi
gi+tejg62J/cdckKlX6DXeNtpNWlNJGP+SUpq06MQqVXcFxToI7nJu0m8sXcU4Qb
IPNOm3wmK94me6Y2Hatjfd6QYpZzC9T1+L6WUcdG0BHT0dfpPbdW/Ctk1ZvFY4Cj
pUEQe18iVKGhjMrI2tN+OSweamkAYHw50eUEn9cAYiJyrOSAlbchWP6CSrnII6o6
SqP/gDZ65RpT5s+RTJ4b1zNHr2eeJVCwI75M7lw3FT5ks/MO0nXtxR+qktPowc+O
mTRkXMG7STMckCcoZPvsn5PbLI3bNFjm2wNqkDBaJc+vOssYsAoUSzE+sv+RZ9Ja
mNmf27giy5BRcZ5Xmc4gaIqzNAP0n1+IJB8pAepEPYzlzNK4TOEBYiXDa9T0WbyM
BZAqB/ADobWgVS74IW/GGRv32xyD6EOfCy7RAnVyQ+L6Ee9S1S951Taro12DQtTt
XiMscf9q9yj8PZ205RDC5PqRMA+50TGJJ62DVPrPq+fkxx+/OhV8T26H5B0v5jzs
zZb/Wy+eWma1kao6kiBXrIJakgQhWuKMvODpCYxWudZAmgIYNyRP/bp3pWYc8p7t
biQqZrPR8sDsQ82/lRJekNTSPljGYcFe805OFZ3jbK/bDS14nsoH+ZEWQdzQnUtH
WHZ2KS8doBSS0dK1bkI6qmKKZPCDiKVcuPTM9z/h+dXTyUAQPYYb7GJ8WnrMpnWw
ix+XHE/arfuJuYeC4xRc2IwBcz3DygS3SoA4RySO4nj+5KVbv+uqWjDH3M8aKLmb
FyeePpCW7gTZkK8HyJ18bycu2bS4MXspl5GvAIStoHQeZFkIGzRHTWR6QsNEQW76
uwTyhxrURuJn19jthJ7ZJrs5bg+7Xm1uWxPd92EeyCrCYO38CX57OKxjLYIiEr1u
eH+TBHLdJLUZCx+rUdbL3W3HHJazIWiESM8SGpbix0cPuT2jVcAeaGg12YbhO00E
SZLXJYHilViXIDsQEsy7ZouMSc4Bfdl19K16hv73Dwx967A50oobZOWQaVgDrNny
tjd0m05zW5l33j7ZMv2Hd438L6EIozZzNYP8CqXK3dhPpza6Z6xTB7/i4w+Jhxkq
MbC0ExhCN+sxMDrdfyfFGC9v4cMCqpMg1Sbe2AOVWaZpq6MQ73NAeZwLd9BRZuJH
GYHqrmYI8uAcHBG5MW5w9eAx39bLq3nLbsqjwgLBXMJUotJwtiv7Ge1GiSh4JeFs
9xJWz+ufUgRNHEsJqbUSD7mrKldIEO+zhL3V4Gi1l+hr2qz5L6I2Seed5ZpM7+sl
XD3wrz6adMdC71zsQFrMZ9+5+7HkCx5J/jGpJU3i+EYp9iVOANpUQXcVbR7+h67K
Ra6AF/TrL2cYIcFvqEQv9sqp3lVl6wDh5D7qCE/pJBGE616XxAH/3mk7sJmaV/Wq
xRrOJhooTPOLOonTAgolsyuo9J0lT9jghzrinx9MEkS5Td8PeCmiaZLaE8oxEGIH
8bqmsKP1wXcgahW/AQH7TynY1hpKXeLR5Eno8+zFw/LaD/5oXXOYna81wONHr50I
ynBaWia8EH/I25rGqAdp/f1aLc6oqIa/iAfuIx05j9Ky7FL9JsVGIDo4xBGGq56P
b7kplexPyNF4USG6hE6jIWCaWjRqM3DRN4kBek7jSJ7cquufd6oaxfq0LHXASiCP
Qta0sJ/CzSD3+qWGgEugeR1x8hIPrPzxOyPANL1IZyplLfuJhoo9j7QU9H6PJaax
RP7l5FPJrbUJI92TiNu4OWK03JTXu2j4gI7v0vA9GUGIRbVmBWWBRIpHahNzdHb5
xug0dXaaSDYDqht9bnfEC8nygV9vESTDx6j8A81bX3AWCG4pF55Hx8/wPLAjEOtc
8TuQadwJdBe1zYUqIWEUQMA/8pVoxvfebsbBAdTJ6XBPatQCXhnHiQDW9olx0pJd
kciEqhtRHMOz+TPA6HpGLrTxVoNOPi8NeW5BDgcug+XDRsKsMYqve31ZsM8g4Z5r
ehA+2ngLpODR2493xJRRLWa5CTzBeUUV7KHZ6d00w8t56dwvoLhbdc29q0DN3olM
hL92JS0JGpo67wacbX/cKMYfyoRKmX/M6w5AF9SDqxsWLORAcXVd9/mlvpgK/J3F
sw5XfBDq1cangfv8YY+IP3All35s/Q0H5/eP4U42wIkh5da2+QxThUOPi8a1zEgU
ey864sbCf5aJKhk1hJktjxt2RypUSlRlHC3b6gzUKQho2b8kAqncMNpSD2sU18YJ
LBBWEWEawSQ4dOpdAq4zwtP7v25yacOHRp1rM60VM1cfWIEVhEjsiMvvq/i8T3/+
Omnsru1JUWHpe++SUYO74NQBIVPODiga3O/NcnTa+NvC/QGBhSNibJZOpsfL+PX+
EE37sq5kI5h/ZuHsoBDnC2X3EYnf+aGkYfITK5186KYFKZRI4Up3nupr5CFdduKZ
wdlQPojmjd28nOXzzmI8ilWKVUZ0TmMYbWv+/Eo3GWn8+5Z9Bojl2kDukUFCA5ax
Wzjj1tSbxezLtYsReE47AeeqUVW5HLWrPKHoWSQ6E4gNeQ/xTfNS6zvkOFMH+EJC
3ozaOBZqTCacpw+Cj2nbWchPc7f7WerY7uWUVtrva1g4+gpdyTRjIOM0cH9v7Net
FonCbERoWohQMO4axmevzRVIPEINETBJzyKeSRfICgAEoiSGmA4bilum49GgN5gj
YgQ9gRiHqLa7/9maKbKKgjtJw+BSaMevBQ6T8Ybrz694Epa6rCadmtjHQXlgwpuT
wCM9BQHzuVl94qHSg5eb1YZD2E6UTogP5DkgthWezsE7UN9uR+EM+LANs+kCsOYC
wBqPy0De6aZzolwBNqmqKf/1sIXTba8WKTfZa/PHGGyPAvC9X57ToL7+UhrfJWY3
Ck6Qqg/tZRuVXn90YwH4LWsaggI96g2ToNb7d6lylLNmrRw0JLCGPMowVswTsG7u
ztLbNa9udFeuduA4OxkYrGPEbGSD7YqD6V09wwW4QxRp/vZ/7L5X+qLO7HO87z+s
Thi9uqTYFEoyb4f0fqyzojY2f5ITLZpn7hglVbpu6nKCB07U+n0oXIBgiCoJg5n6
ce8MKVvChomxWe0/gG5+Fu3JzMtO1duv17qwcJHK7ZHpAgq66K+ke/kkM980fECk
6NzKFLA5V3mLxXXU9V+uxn4va+3KpzNk3S1RYdghOErenE8zu4Hq82WfMwOHsN58
bCV+bHN/AcjhzMcLOhm7M9Tzj8tisOAYOYhi1N7G3+NMECuaSEM1WUSw7Oa2z9ag
5RrG/SstwknFqv8WRlL4Q5K3bqdwNyqguqeTdWG/bPn2jV4JOic03u85FwS7HxgZ
gdV7sjrLBb2MyljWUzbWgCVOKzAlZ/9YCaVzY5C+8wMBJTJhHOa5r35G6TE3ChEy
T9tLBamc5qQN5fyQJrTTl0cZUQPrITczjCCxqpEqDoooCZN0R2QyYun4KGuw92Of
3tlqWsnSimVn7T47bsxiDAR2T9Z4ostMnc1vYOl913bDi/xvQFHIgXeF+Ut7Xzy4
5YQYHJDG+ivL7CynilJZ3fW0/1gUlC92lrm0BbLr2zCuim3xMMx/YwqDwKaKQ/Sc
IwM6Jx5Qbe1IL1v68ycnAr8p19Dqv4tPsQlC5DdFmr/sxFJIojngzb/FSNSj8uKd
eeOGva2D0QEthsNMQF/y76SUm2alntsGZ177OSwcTgXZCVUQ7zUGXW3wj2g1ONkF
OV5pUofN7VBAjRCUpDTarNc6+oOrsqu5sE98Jf9bACM3Ae97i6S2EwW1p9cu2UeI
jPOJqj7Pa3dlg/p3pu+pdaQ1tRG6dT+cyL/bdJQUzX9NjF6q3Wg80TqcdgtswuWE
atsWgTHtzL1tGGjnxhtENA990UkRFOMhvI3QDeXO0B38VC6iXYTCSsJQB5gz/crB
hcHPbi/RDoCztcrKPmvkYun5llt/C0sAhDuAakJCxG8BDBATqA8YsTkUubxIIPYU
yD9d81qvez4gV/LIwKMaaiS8Aosvn9TUtHR3zg95q1JBK/695+gIDnOmU0tp1y6u
qELOZ1izu1EnDzMWDzPuVQRbaeKipavxMLMZgR8Qa3dGBgUdree0pVA4D5U5X82a
6pxSC5//Q7v1Et7URYi1EkF+W9ixkNV7r2TnllUxdA3NjLAuG0RuEpdyrPBjBs3d
rcqsiqxXDogF0ia8F8rLuzIw4MKe1iMiJ9AqLlN4z+7P6SCJ/RKXqmeTEeVU3aNs
xbjbRQKeYn8AsnKYDhaXlLnp+DiHI0aPHUCcRGcc3d87cmLL63OFmsGa9tDeXuFo
rtcPsOPwtquNMwcWsLFe6CtfT9gpTpnE+g8jFOK1iWjNnvEU0asK6GY86g0JzfW8
c4Ymjq0PIwLwlsJDo8shuo9JmLzxxb5Jt/mmcPaxoEn0FzXRdPqX6V1ea0gs9pRj
v2oUimnbwAWGTlEJiISjAAzHBfkz7I17oDWtl9uuZrWzVRfvKxnA/W9/4vN+ufzq
mlRizL/QrYBNI+36vAkUOWqpPR74pLBvBEGKs86JBvWOkTTRarW2/RfnZ4qY7ted
8xRc7m4oNv7svKClxIB8INXGRcpfaFKycvHsFiXFJxS1834uWi/nsG5Sx+dQmk8C
tc6vmXOjt1sA/tKbo930fefon47rTMa9MU+pXRfNE4ZFYLKNfQGsQ6g8M/dgFy2f
gi2aPyexdm58XV8sHjXQ28KmKEJ86BZx+xgFb27dstxxKrxFvkfjmCRCq91XRdS7
BY1YxzCyjRodKhR3xlMAH+JAO/pj19qYrxSxltiKpzaEbAgxvJS/Fq32Ym+uI/gO
puyQ/OBc8HnZ9zzPHI7refwZPLXUhYSroaEyq19azPiduWq8S6y2MXb57EzrVUZk
G5nRNzQIQGZBv3Uk8x0gN7nJk31kwVdSWAkm4nWvV20fe+CrxtHB3XTdxvOks7VV
DsxRzLz1ERZ4jdqPQyEJSVDHEmpxwTdSeeOE6fSNNAJP0CV1GkOWiSG/tANd3Wnf
jXfphTnFrPVkv6hfWhNwIoGZQlghfygHvz+hp9HXqM+LfymhKkW13TTqM8SU33Gp
ql5edU1NxXgyNG9OW12AQJPMXrxyWokLYaYQfgNtPqcrh/shwjimcWRiGWZ64mRR
GQoQdiFNBUxKzj2iu+tmZmjnqW92fEo1pf/U0iInOqIFxfGveyZFkOnrdwpGxzs4
Unn3YpHgyl0FvFPirNBw1LOwx5vNVAOqZqGcPAWXxRuICSjRHkOarwzv0wGZDFVB
2Ke0Gb62MPeB8q0omFSqdzuBQ5QsPWpcmVSitLbrTyscvndzpXSFrmLP8zCBG/W7
3zVZxStJt/F4Iitc/+WNdButu+7T+V+GqDHunvOPO8ouBzXKcLeIDrdzziCCPkDo
rGYFi0xfIMT6Ic7fWuKSdIFPtGirZ8r7mQiSZahrV2KIPjIk1PfMeRREcKdTy43B
IJh9h0/N2+dAgJFuhvSYY2W04+1471i1AcdlnmNcTeVWMoYUSi72Uk2H787gNzZ3
E8WAGhb34n5yOYP+fmKNKrP2DU0WksHWSFW4DX4q7BHWmZeo5cE4Hx5/v6HFd4Dm
8VLwRT7ohrxxPKijjbIMAgwxAXb6OQdRgyai/yNVfZyfAjVGS+aG7+2xdZ8UJzTr
SfoMiUm2KOJ2es9hj9CPJ13kgR96rdLtjBZa4FlDWCHfZyKdwXratdJR8RZmqSg4
F+Lp10uOeLrAu7VBLy+DTaNrD4GMBLrxp/WrMvQf2O9pArXMg+reUuyK2+oc8+oe
GbbYoCYxoVmK4o99PzaJDpMVlqoVXx6YbtpNiy/Kpf5JyJv42JFE1JULFNBn+ax2
0FRUB01Aj/Eju5yrZU2E6qIPx9e8tx+R9/ZEuLkBGfwiyJzP1DZ8GMBhhUWrOFUB
5LmdXftTMZypKfP0OV76za1Repqla3gtylutaXc6aaXdhCIga9tE66gq+hOUsV5X
FDdchBEqqc9KsjkhlgnDQcS8mTyt9BzrDABpmqS11kejarHJtnJVfJQ/4ej0TM+C
7mboXky0KG47psUsG2qRKulW8YDfM1/uRDV2f0XDNsR/dB7sP03828FD9RRK1/VF
oJsB7Q+BqfSerK+kjJgHgK7SdeUczNdLMUcaQAcMYB68rieMe+1jhjK5++ErLHme
gDrKfVIWWCy+iMd2t/FhfyQNxhAUPQyVRCoJb/cps1aQ91KZxoLNw/pGwczIYc+2
ihtxY+pLDWwJhrtmbNaZ7lNetHo57kBN3LiahwmHgeN1VUbF9b+u5JyWwM0pl7ol
9+i5c2WIbc23QBTqUzwWrf1RsJpkSw/27QWCzni6aFHHn+6o5D6bOZZ8IBUIQmyf
PfdtB2GyECdHdSxXjE/a+BdIx5UTpR5YHxImqIa2OxyD4XInyR8nto9za0ITSu0J
+h8+V0qYN2RM0UO3i6Cuy4CkXnNd34GHrYQ0UW30j26sqBfhN80ss1BUvqIAZ7UA
3KmOJ2XPFa6fm7JYp4x0aj45Qs0OqQOQ4Kp2YlA1wepDgP8mT24Ki+dQ3hOScDRL
tuY6ztyDm2ENP8fmTZn1W2Uyu4BKjPh98PPYm8Ga8HlIMwyeKlIgXm4sx3p2lvSk
OpHfF8cErtPwlekL45T5OLq1tdEYFy/H5YfUws4N6hJ4GsoLNNgGg4dRe6fepJim
UKhBkKMIc9hb8YQ9tIMrBTYxnAKqJr6cfi70Psnnjm7WgqtqMCOQjg0lLyqwIs1V
KWzyW8kPgOuRXD47b7AAS45LXF3maUbodbb1yprXrgXyBRjrlgqOz7Hjj0EYQhk3
pN0u53lb+LOrix/ppSYEceceNdsLy7LY2QwDxEFwNwJcjD773gMHSlkjes/E2b6t
rTHzbhMiLVt2UQn2UsKLSTG5C+UddxTdrRvEfPbNCLgNoxvMI8gYYRbtxfdKjuHg
P+HsHKpI7Bv8VxJSwX0wk5NGCWtO8EloN8IkhpNPjmqziXQ29+U0pb84+8ZcRHDo
stEO3H7RZxLomlYHA5Jg7xVoGsXfLz9AMtGd2hcY/GEZiMpOI3DeI6O68SzCWb+U
VxGZaUpNt22YgVuwH2Jos8nJo0cpUfoXfUijrGw/lJSx4v7PJHJDFBU0/0wwpuFt
QxnQqKYGhupFBP8kuD2E801km5lLlQjyUEuOAzG1bpKkOtzRISdkEQN3kynF+0r2
vPxhCU0aymA3UbnxLRK/+FZniOeM1iv0QyyMWkG1A9n1Ysm9G0o9VNYB8CWd+0UR
Y6dek/ihtA+buJILsRSJ516BY3xxAlKOqX7KIVikGOpKhdpRib3PeBirUkz/ClJ6
OGxYY7tCH+cOXRDe3b+JOIcYQ0dRgFILu66++ODh3hPUhvrdApIdHZHd864FoIF+
pvNcjvIuhKRsIZZrS/FRthUZnnkFtftAR0Oyp6TR0gQRk1BYIZV9v0aGPRl1/U3W
xyH3ro2s9ust77HjvpK2Dcw2+9WJTJj5OUS1GoDuCezBMvJIv534qQXCa3K8DWcQ
xiPcxQqNKXB+3wmp5ubLBdtbO0hD4rR+fwJPRiprfR2Mdr+y8I+OAC0rD4O3/7LO
XWBZ84giYXqWdl81evgF9V5G80CIherTUIm+Zg3tKR7ygFWWBSwg2y+QRxBJGESw
5FDQlo984W+ndvnApnHPJXjI7S0HtXIr5PocMflcJxD28GUKC3I05x7/WKm+ztWU
+CBL1DfS+3XbE8pjG55F+nvvQNmmqdbqbkMmM2zu5x8VgjlebJqIs7lIxGWzNDPU
iYE9RHegu06GJVEdouz0HjcW3U3/68ubHCR4L7GV/P/7DO/TaLsYz5ZuHi58P90y
9S+N8OXiOgAMLXB6juN8YyWb1sk0QEWXtD12MY7iVYujwF/TNTFD765meOgJWsL6
1r79N34Cm+VHQk/oMk8UfChM4ZTL4ZFCJ8GbWbeFEejtftvf8FHucmOBymx1/NO9
i8nJvKUxSn0WtvZ1urNTDmcz15c+axkLIy1N5/DkuxBgfT2ltOdUMT0IsfTsH64f
h9lw3IhC7V/b0wEi+ZptpEgkyz2i1YJAGk6Esmy1vt1wbBWHQLNEjzZU5hQnmici
6p+QHLCvWEhc8QzQOGkdMaI/lDP3p4MvFK5bTbJzVj0knVSwdDsTxmC9gZD+p0Rj
ILVbvxV+gBDq5wK+mkmfdLdR+wIk/eCN42UBf3F9k7lMzISDmi8+beALOUUY06ph
CeCHdsC0FTuSGP+KZ0wzn7I7y4mMQUxzU80Hadv82s6LJ+IJgQOhRmTRkRFagAjH
keFt2bfSjbsTU/zvcZoGhzs4dyBvV2c2ZjGa5M3BUgLGdjkjzO0jocu8yCRsP9YF
ldsKkvf6/7SvNfvym67kdZRW2hKsM5Az46syFtM+9V7f8pcBNuTJCS7lxoEhat9L
jYtGMXjqqmuXrN+T/JaLEMxq0ZVbxSN1Hm2jIijERSqVOwh4rA+QGEq+9eGZyAhx
6RNQdVf9BTEwd4PRxuxz0yjZPKqEkefvbWQGgPVULYq/Tah9VYsHOiARRH4YuWZu
TQXeBLWYgJHSHZ8WVwQdtUe9DLVK7VRcxRzTPkD/7SoVsO/BdsllzgE6DFktCTVW
4ixE8z9/vrkqX3TVA/vtrgKxoejhqXhSqfbh5vQAUzF35Rz7kuu0FREyMf/bsdts
TJ84T98dLHhI52GohBKebmpEm1xmOxO8YxUaJliiAcEQPQvN+Cs8NoCjHhnSeSLz
9ppQ6Ago5d64crPS6yoXe2Hk4bHdkO0UeTxG91fvPUg9eIQkk3hGg3IMogz5XdP+
61Q2YBL6cQab+DgFZWtQet2DI32vs6dvlxxeMg/qMrFVSJCs0lHwgC8QGv19PMS+
k+OE+a8iy0u96zhLNqoZbm/9eJTzA60nur5moLE3E5rhpq6l4mZssALYsfZQE0i9
a/CWRShJOPztSSdqx9MXawlwTozUDJ2Kw4nIr/hiXMtx81+qx1V8yRO+MV4yTHcb
J49JhJhaPD2zbQ5YWHQT3ByYZ4frENIcHLB4Zh8iEFcbwecnYRNfsKkQBWUPqR3q
4jZ1Yb9Uv6ADa/aGl25YNY0Hxih+BcVAzlxRHA5FIBSGcu+tZuEVDTL1H/H1RykY
TxH9OfxzU1fuvTt3e2EnrrC6J1/6gK2jdtiBv02kqqa/eULdfGhiPua/Kdx3h5t4
cY3P1/heyEt3oxtVv/gf1nr93mOlcJ8R2y/Hqgz8n7hC/7XO0v6oxMw8Xb8gSudf
OZYGTBaMmBhMWpYjwcGuIE2sK/jhfIiK4JHLkpcjRaahnbviDBG8o+2DA3/Is/v7
MWiPb3s2BZFf8C3OqV30hyy9n4oLt/cOtHwiyUiQ4nGxii+uCQWfLdl56pVAjAzp
uWOuapadeOKQNBcmobnhenJ6VGR7qRXIrrhzg4rVY9pOhqxRFt1wXvpL37z5SWk1
1C72yimcuZ2nGweXTgdqiFbU67/aAfC9nCnLbLiTSPGFZrvAaWXD/4qHogtEYd8v
E6NVq7eMChEFMXTG65J1GVSdA3DNuQoGfa35+Nl/krRC+5UH3Pxd3EV9y0GOBieX
VTthcuya0I8FnBJEncH9LLkI/QWqvYvkADLVHY7ni2ApQqrRMl6lVfMVWB+YvlAu
XGB96kAKq9yTroxErdVnd0v3plLlxI2M6cy3/upvbXjQslZacxcTJwmb62XQYXKr
t02EkuLo8u9NcHzC7w+2rnlj+L5x/nBJTCYJpdOaqEPHpPSLU14GfsWHwzxqFMxc
F9vPN8ZygJPvQ9aVSwh5pwDOp1GpsiY04AwF4YDPJe9Q+Y27L/WmHv2r8KgZOtqA
GoISVFZkjUYPXNM12eRA97xLKj53k+UlAPAGGXC2jYTddKYkL4djBfCpHGgpppSS
RiU3jqoKKT9q6GkIMXMpxifJ4CNLj3R+JoNnPZ4zpYuJvUyhzifpjztLP/vvRN4r
O22n75kLtSKSeZ03F3iDcxOBWgASlIZOoSEg68/2VEnmVKNg3nToB0XndpdlxDKK
DKDNaoi/5vWuumfh+FSuB+GVO+WFynRcegj/AERL70zatrZZBNp7x7Zr3sKQYfk/
Zd8pbOvFYuYM3zJUi7sZdtToepzgalyOJ8I1PFIXRu3cR0B3rU1A0g07a1nAIb/y
/4afongxgttbbjGSFOiou6zdGJ33xwRZPIVWtgpvwv7Xa8vghya0tHHMxe9sgv3a
wVhAd/P+QySseLz0agQGz6jap8eCFiPJ4pLAQrV+vRV4XC3Sf5FZV78Xm1Vqz0xa
OHvP849d4X2MwTWVzhzVNLEMOEMY5PNrIaL3s+ZiGowUGQ+ZoWFNakxmMVPPHR9L
MznLfLMmSSoKaFB26MJ2oMAiyR/aJY/eldQWvgk73Q0lhmwPV4+IOPDswcTthsdP
7+RYHish0cWmV/6jyjrmWyk0FISuzq3T2p9xxDU85n2MB9prmJ/6Q2N183xSz75k
2N4JMVPcQRixgcqqknCUmxO/YVqv5CP+YvM6MB1RGGej0df1JLlI5xnwVD4xSz/o
Y8oSgk9FEdb3qY8ff0/u2sLBU/uIiUg4Xpa3ZW84bZ3upLERApivbffYPXH/Alk1
czuaH6ofp40O/5zoKSNmxF5rIOPbMBGGDmGVYzyn84C6XMm9l1mpLzjvqKUP+5Ss
o1tSfEotKvCUcdSp91jKwPvd+I/+rtXry5N78lxENRtHRAPyYy485ZdPPMiy08w8
1xw/0wQpXVAd0Qe/+lWY2n0MF9S5w2WGxuFjBXY5Co9ZIp4lJH3kBF5TXnTDlSRg
9V+bzk2N0gx2zXnwl9polURBoq0afHCzdbI/uWtGEgp1O25NAleB0GHlFkqgizse
pubFmZ6QFt03SWXg/Ufj1/oazQJqTwdPphrF1MKI24tzpqQvYLU5v3N0kAbfDWCZ
eB48olFrIvuEE7oFLucrNq3FSDRFPmZp96sgxL/k9zePWOfm4BEHniE6LCLzDiXA
lG+0RFmoVhFfDftym4qOE0Mu7ULsMb7sy7MBjUnnjlQy3NtLFvh63fh413TRu8nj
m7RS/RIfMIsmvfHbZr4zFC3tIHpAygYkNqyDzJJscRCSd+IOq9YG5AtxlXv/Nyuw
2ZXkK4f0LW04kB+amtRlSb0IecGppzvS+p0BXT4Q6G1kr8fSFGdYGPRzTqWTwrmC
d7aQujkQLs4ewuARKLHiFCwMGCeNhehpadXCI1fKG7zW+0bcCe2BqGZJHtOryW4F
BrJPZl6tCA3vwFcuzL1MlirqpRBt2y57xtAXmhllAOO6dAKjvYPn+3WTmh1rhoSd
vrp7kVsNGSzVrqTk9b0JmTR7J54j55Oy2B3pNEbpyLuJBU+yeNRFaOrpWPib0poD
vGFYoHefKBogJEsoVOxplBNXrjVMjhoaZQGn/FCXo844DacT+ud7vzTvDALoKUvy
CG1WbrPi2JH/vrChNQ2OdSssdF4evkLJY5qZFc2XUfmFvVUXUBbyGcAKiC4afrBx
dRI7a3N4fPT3fSbDNflySWeQxevxESXVsX4M9MuxqVaMDX2TGtX1zm6lYcvV3QsA
UVc2VGVen21j9B1n4f/4CceDy2G1coArPVrkUzrKlJKv5zh/tbH1hsgRkHxrX+TD
G6cOQgiC6IAGGBHXL49Mg7Ckpi/8LiSyd/HagqcNX6HVDtrjo6R421AaTZevpWET
68iOAyzUwbVBKfZAJPY8mCvOgcuRrSqLmfHHvHZUfMmXsnVvda1HmIMgFFTzjPse
XUMlDJqBrboM3qd+CgdITeieAQIDcy+g1XevoNC5sH9V68nucjGrHot83E5GRBuy
fc61clgLptEZJebBS90flpI939hsUbOxIIDeY2HVUHMVonGjGNADgwzmBurAwU50
Q3TJRwhbfJ5b7reFDyc1x5MIz0JBhNKUWTbMQR67zfsklEJrQaB6P3IRNGl68h8e
wTdWdTBBIg6iZcr8KYr8IPsEMQa+tM5gGVMARp2tHe6lFlpzAi5r+Az3MR7PoZ9J
/3FYEABkyzY4B7nNZr79E3aC4lQlbyYYBk/sBe7JP9GWADrwP4GBVXC0+q9rQWz9
5ptg4jlLo+mZrMjc24KQRYKUTUWxo9nUMjwbnkZnjeJmtyDaI5Z2HZ6+0JlU74Qb
YmKdx7ZsKUxrPKQUODcq8raLvzfs4hZihIZOIvi0WLkL4dZXjvio16+UyWRJxhsg
/79VtOdTNYrrbzoidtw2uZUIuPbvQxGJ3djHNmf8OJeb14rCXk8urU0ye1ETYUoV
dhXXoKmBDux3KzlSU2Ey9afqCzuHYhrfvBELTLPVMHrwqjteW3o3nnTt6Xp820kG
DTWTZhgXyLHTWvbAQnC3brdHWDfN7pUGjsoukrx+X+CyFIGNQunEmsF0bMboKbXj
+mhbHnacjwpl34Y7bWLglrfeIb+Rahu2Ub8R8w0yZuC7tmlZ5lGdfr5/mERbJvuQ
hFect6BYtVcdITA7C2HDhSsaJCVFRTUUSvqcapV+fABkyepNWiYLBhSwDD5JM6P4
+gGILc/eGgDectTPDIQk4QJrLHA/18kEu6FgprAnqKKU512/oPCPCjUKDdD/BtL0
34Dgy00dNnJdOIB5EdCIrYYTQHVV7NUAThSV1F8XQ+9Ock+Txe6RIBivc8hYp5v1
4jQC2rgaxEf7JwOBNE5M/kBtFVVXnyNFgqkdQlW6R5aMZFhFIjD1czyd4qf5jrNM
L79aAZpEIR1nKDhJ+Q6gWlwbz6ssbGu3AHlPvKIMxp5IDgi3sLB4EdfeBYlALq7D
8ZUlhaHVbksMhJpPIrhFl1HGZPgpikdKu5Sz1RZI7gGGbdc81HDxbcYLVaEWlHB4
Z3P3/mmSeMeJuWa0CiyG0e7wdrQvhjpfUCzbt2HIp2MsWbweHZEkbO7i8kAMwjC+
sEzTmZcS8j/2Y7Ql5lTwroQrGoj1LRsgbh6jDvqZ43hKY312tjpwZ+CIfQMx7Prs
U5UYRO1ivImyor0eYzKqIGdAjCBmwVSX/CYj1a/94OIjHsMiFY4e0mZa0SJYZehK
A0g9lTBJGxzyf+DKsueSLmZBxhWQhY5cfAoRd9eXYke/MgMjZSO+rVlyzCg+1VZW
5Ty38/mEoALZGpOKeyGCegbO2OpJRjO9a96LpiaavxLNdXKQgfLynKCyHshLSdIq
DmvrWIn3SYJWmgRsrT34SvT1Wo2KA3SrNlk6KSOhIlSYKb1A3BJuNNvwM0mol7wI
vqqOqhEIBX8q0IlfaqCwshirxgPTV/GYEzp3fDus3TM/NZVTh8/N6EG6Mf5Bz+n2
gIiTTFHnPTwgol+XwbxKTZCcxp7q4MpzOg/Et0rWiBFdLCfE5Kf9jpifcWP0NoSC
QDHJik2vZAtSZyoLA7LnMWYw5Tacp4FunMe8w3ORN1HHz6Qi4WUNL/A6dK0tmEmq
bLpSs44JouNV7XITapiBPOefma7YkvTFSbEOJXioUkSKmhTB3Sy+7EoqkIT0aS+T
F2YAJdFXaT3NgEQJQ2YwuwrDhctIK67BF66pVDhB61+sF6E5rGULJAdQ0MdQrURr
ruoEu6cIfxGEbTKEPUtgvCk9PVRsloDRq5ItpLmpSvcQ5F5erx77pAtKZYK6qVrJ
HP/zNNaPslpiFXFEYVHqeHJ4cxBmJllaWlRn1bATJmhICmTz6vQKBY77B6f+kBym
m8MRHuUIiQLCK4AMVox0DSclo93TyPKFgqL4iaR5Bn6qs1uyVs/BkI5l3JND05u7
DhJlMdvxprxNgKrU5E7PasC3+LLjJKqCbXoFolnPq/CWrWNyKTvJZT2VurkXrvlY
bQPnED0Hxjl+meUyfzTM5zvoE/Uf65MbOeUxiFx1QPlgcpJwz9BZs/AsgBHYesmi
h7/b9U8Z5s5eaPBQD0MOc8y54ElT/vphdlphHwEsfBts+YyCQtRw2AXq6DXveLYu
Eo/wj1iVMF+fNRgeFvgdMcEHC0bRfpxjfrxV8q4ahUtqp26fNBHqqsqUg8uiKYi8
y5BzZJLHfvT8YfuWAuEb9+ifjocJ6cWm7qX5503U5/r/EMbjUw8Ew2k7jHu9ZaXr
bhwNxi53BVRCPHceG2Txjiwx04sT2PgWwugCYxdDMTpCyBZgOWJJ56ykVDjZgDEJ
e3+PE7htk72QCDDHgIS4W5l9/YkrE73DqHWwGYUxyurid7irlAJ/LO0b49Lw2Jqy
HnGOO2nRc/wZTS9HVP9KdPgQXHQFkpbAPnnDBYMxHWDCQqYGEgluJ7yAyrAZeF7K
RJ642eJK0WoDuHcESb4QiUxY1mQY6mtER4ElhKpre8JT0PXz6oJv7I9JSuApF05t
Dy5xvshN65+qzM4nG1By0WSdRc078FtEeC10meSQd2QjVUdIeLokYWt6V+vLF32/
dUozysgSUiyv4ZOOj8g5pcCuQzp/fLIBYyYHjx41fNxkBmHTIPmR2NVVAqip9iPL
5uV0i7a7GHH3sSm4NruYBrhHfQGtolmKpW+mDGC0sC4XRVd6KbSwCdwR5Rti37lp
QCPmOI1Jv+2u4BocZbXBR7n02VP++B3fQ4NTtcaJi8d1eNfYh9BhwxoxEWPrhpr9
bRuoaAHAQCiYA6ofM/KWJx9k4HPdB8Tb3RPL3cqVQbMLN3Dr0ZDSOGEoXrSjF7Fq
q3yeupw3bm/C92QaM4gyTfr6DhRFXnUo9id/Go9L0Hb4V+JmCrRY/DKwIMSmN4yt
cNzHPIyt9JZpHeGMFkRSUjdWEiAV9JuICiZLshzUugKpc+/TrLb92goGsFbKAJVO
6+L2S2uqX7JuGmpjhY9pH12EDsyl66YiF2HJfKmmn0mlxhPy2b22h5FvJC668EzV
mz3Wt5BFbKG+iV1+9LSs/oMFqgx+Wf+Jj65p+NrfoMACGmgtfICgNemO9hlIL7uB
0L3DFUqxHCszlsaiBoAwlPUME1+lC+1xjhIWvFY3PmWt7aCUOp62ItFANumJmjAF
awf4/q2+5ilkxrlRX4dEViEOfB8PLN2oHU41HLiJrSvAEdDazJb47pft4i0856va
6k7vicf17H/ghnbAZW5I1DmH9cw3MeP27biKn8AueYHQPQ9diLAW5SbMaMRlJbsv
VfLzX02zD81PhgTJyLhpYtpEAnnNZPLQT4IB8PTDG1Znw4rNJRsaK4kmIuskI2a4
yC3ykMIvnjnANIEP3heeny6DwWv5TXqanF7QXMIODDP7B9Thh/MkufFoJiJfiCVh
29nKfKzY+NXKnQR7DHPQ7yT5re/+UzxNLfH8PYq/e5jPP3pL2cdrAl6hS3RTfVFj
WQQnm+45c527FHPIJnQ6ChWwrDhKhWl6oMzoQL60PCWMoJigTyycm3GZgee0xaA/
evsfH9jR6YX3p6vTpU6pHf/BZHtYCMXW9D+6rH4O/kJYXiA4xX5MCAgmMU7AtdHz
F2fgtO+cSZ02+pvv8k+qa1oPPOOIMLuc0vHCaoP+pp/fZ3VrEiTcU53bsfCoKswB
ftwUHVblqSjXiljiZCYKsj9CLTn36r6RJLPYXIErCdBCAJGzlCOmUlMLaHrPgwLh
d7beNO45uOvvGLtFwOkYDFBp59i/EZ45GPHANNIUCjYWnc8YEf4tiZf/xngsvFwN
YgMxksN3vIFv/jnA4kKMMFhfV66WW0Qb1XNJJjSLKfU6SoZjq+wF8AigEUaZKfnq
S6wH8hmZgzeiANXiJu4wCNebDWKMNI+1TuW7OLWniBEzu/DEcD2F43k0nMQ8obLW
CL/zNfVdryeuCsN7zV0QsfkedU5N8uXiiAxJFEmiKYyjdsmNKRr37u1Uv8HPoKZz
5KcblmAjd0x3i37AXLvNSPUCWinLWEQIHMupjU4NIUKV4ecQ9GAoTFMcConTciQK
W9Tu6iu8/s3ktxTekrr+AUjV+RMFRs699IrSriot8Uc1QfxD88kDa0EQCdSIumlU
s+LpX0qLXaTXzttFBRTP1zh4Sbuwr6G/aVBnHw+etZ5rKasUGlvjCZ2feJAaNK+L
vu7hmNBMmLdjvRc/XkAfagUsYY3Tw398qOCa9jj1KA8yoUk1iFXZIhHSEtqwlHMY
XZckeeXsJZ1UgDg86sPOmiCkkUvYjfrO7bpqCCgwYo0gQrPlsZgfyhxAy9AeBkes
DhyWDw1pWjRuu5SMkC5txn3lEfdasRimOmLzYTUYCp2SFoKBqs6yMnIGta9k1K7J
Tl/v2AMVN60VpS76G0UoOgP7Ne99hDyPWEcbPp6CzInmaumEZDAOnRpyk2R9aLH6
7Km0vMlBGNvtKsvTwDUD5JKsblPMwFCxlkvZcnolzZs3gCf2CV+bG5rH9/VC3FH5
/cVVBzXichaFuctdqSsOFSJwTHjVklPQSyI7eVO2SC23dTJCmL03mWlSe835L9ll
p51E2guSMGPj8srV4WwRmgUv1pYX8OBwLsl6TmZBn2NAAGcwBeH1Q1tbvocfstq9
z3n/nJ8SKWmTgx2JP5dY+yRKiODNsXCgX+w265GurP6Ay6KN8EQZz3zM5ptBOTVR
yhaC3rWtIEKRo/4BTw6jhXuNbxXyy0Gw4RR+1NLuWQv23jv0LrITvUCoFJoUXaRP
5HLmz9LjgIbsKBwH7yA3lGE8jeqmN1xNzKtBl69Be+se761fFqTbSEZk2jHWoni0
szFUfTfD0Eb/ImbY/tihpTFAkXSmYNHuw9S5/bO7YiW6UaAFUP2Xs/hM7R/G2Jpe
gZNheNGY/eHWHcx04JholR5plUTjcFeBNBVY3r32v5IC4sRTwOBjJw3anz5+E97c
6Sjz2OhmCEqbYEb7QsdAWIy38i5W5IfQUF/9NZvpDOWr4u9NiCK9At0bwRmecHNG
kFvRHOauhcp5qW8W6/mT3vHqinjxh19Ga045YENfzhWPNboEamX7euyxJ+D+G3Sn
dApSHZwviQ8PA7sofbcnuhhA40/klmYPMKhChYIjsrHCvPoO9n+fOoDZrC0Vm443
aa7IGU+bdYm3/Jb8ts0tqG7ySpYWAJM0WTQE9QBbKtF3OGAYZSfg+prBfNKbwUts
qXDzvZ4jXeIyWBwLIyqXdDZnBaQv4lWoHGSqG+RQC6zeYTYhXxMLEFsnRaK9mgq2
I28Dm9pHjrohiZBFy29uEoj274KL6vz3c2v0WL6IUEhNU1AZ9+ybm/S5ZHd1s0Bu
8GehV7BMMU03d03rkwsQNLAmiDt4bh7wlTB1CpwDWhY/uEQO7rh8KzPw4AKhL/U2
H1Hz3t1oRZkRy1QSkADbcV8jTTcHLIHOeB8PKiWw84wCL4eL0ktxY7kUHiu9AmFa
+iLGyhoM/mpPSQyMK1TLzc4zL57iKLyBhwpk6mE5KO5vzmi7nqi8A1W62mYfQf1c
EjGxDXYqG8/CFo98u+6u3rx1+xFNbS37EBFt8oB9/8KSV6NeN3emdlam/9+at3qY
r5M7u5K09LJH/Qv7z9m7+TL5fRB+kffYlcIdNqKNZCaYW4mbSuoZ3wcQfcH2CmK2
K6klEh45yEImuEUJ5AkJyYFTLuVdhR+WcwXE/+s7l45fQqip2mlewWi+x8y9uizl
wvkphEZYxWxphTkQLwS/xA5f6/m+U59vAN6t4S6YDjPiYr4IxVTyERrBb6F5yvs4
l/QofYJ0crrbcz8IhdG1h9FHsHZbWMB+YHUFlnrQGM/+G3Nut5E5OVN0jmQT2oN3
zyJTcuEs5/TtN0oNvHA3+onvrX+0aFWI5o0SWSF2DeqSGmkJfyYNd+p4wkLNA5Mc
LMV8gNk8lk6fVfuXiKKHhT8KlvrTVWbLdCt3RdswFZkMkR9dw0nvE0pA7bc/WEnG
0Rfxvc+PNo3lzEprHTMiWV+GqwB0+7fjVbf0WNkG8ERDxUECM0+jN++Vlrq9lBcb
DSKvK+o8pcyD+V0JMjcH1V/OXi5/sEbN4pcVOSBO/43RUIdV8e5YrdXcgwYuiDPX
QLkzw6SNS0OMCyAscIhcR1ZWMWS3+XZuOx3GclwShDJWWwfXyoa4f6Zo/Mja38wp
PSdXXPb7soliRK3yP7W3mPW9zzNbSB2RE/0YbBoUlVOvdJcCVuc31bvkY1PlJ/SM
4Aq/Nz7FP/SKgegpUr50UXN+gzaG/vDz+Y78KmRUHfoWNBveeUSJwlvDU/GIsIWm
s8laysDLD/oQmS/2zs3J/y6U2yEV5GMxpB5MR7BCHgL4WbuH9WOi4wEMS4okstQH
pHySp6ROqBllCylFn2v2+VHhbR097d4zFz/ZTv5z9fgX5Vqe8NrKdOdexG4uNn2t
DF930/SUjYwfllLgMWqdjUynU44PNATIUVzE5bkosR36+EOAt4BiweTPJEbrJSs9
IPleUy+WllqYOzfT0z9J7H/FVnanzHgISn+w3V3RIGnCdtrZ+Y3NIsZ7YCjBTIv2
mZwyUSqaTfXU+wRg32BbqalMdfVp88n+cjwUsEtVTuQv2ZpKB6gj8drhsHTyq/yP
w38QAVWH3otMhIhvIpf/AYghc6UVAx72ptkdvpfZxa5aQq2wAaNw83mSHTpXzRXU
5/O0ITwS+n6Y0a7IW0bHt/NEvzxbaUARlq7LJl/dYN94rpRUEVy0y+3Wju/7Kzcq
nIEj9UOCTJa5XCStaDgWDgxuSOC9JVJewIvVT1Na1ftA44Cfw10dU0Q79ikjyfs1
wnetyrNO9y8cXcTRsw5i0EJzvjETX0JyCIjAwkxZUXdVyhBr6cFok/0gvrSjNQKg
R8pSQlHdzMB/Q8XysIMIGxUok8OXLvjX72tqkikZeDHNSTKcTZUWV2BV7QDdfEEq
UBqFKqDIL7gXEK3/gcoiQ2pandUsJQHiXdCi3sB+7fCFx9rr7vJQxuCH4dzpfBn8
K25oW/Z1K4mA/2w6un+DxWKBF8ewT4EDGAXxerCpy+38JJPiD+2++uDo2kyrBI+R
gMAh2P9c7Yrzqoqp0E/Ppb/C/EsNYmDSm2nJI8AzfpwndXoR2K4LKrt8NQD0u1Iw
YCLyTM+vJB4v1zl7AWDMpzR8XaDBGVu+BMKlsCFhiDHfNvB7yTc/ywlH7Ffh/5dV
/tBC2RGLwN9bwNeKKP4yMdIxGVJlL+i9AJRjz3npuASpHvH/AcN1zxkKGzw0GEab
NV7nbtD0EyNF8j86f0PqDKN8ypDpqMz3qdQppJG22fcWsNKmxrEtxTfiLf97q202
tBoZyhC5DMl7alkyYbByv2ClHply8KH3cqq2oQHKBm1EX0rEAW2q6DyS0AMcN05G
j8AAHInD+JcjKWvAArk8s6kZXrIiNkACT4yRo7lLiJG7rxVe48Uxst1zPJnrQOl3
vStZFXtXK5/SsDs54S2tfCGpgnU+L+hXe7CCy1mQ7pT2V6hvyVPPvagy7KwMvcK0
PA7fkdFgEKVXbhtc9CCyq/p6DSKxjUy1L31iWgQo8lg4kYqfEbd8dILKymCaBs8f
qHmiqBqYQNQea6G0ZAWh3Nyf7vgrwvLGYpNzhtL6aLV9/x0nzbrXaq9FC6De0kMx
ceZA0Bbfqe5PLH7CiAIXiKq2dzqmfZtq1seVmG0rsFwmYkRnhycXdZvgs2dxlJPV
sxh2W4egSFvCEE3flC8oIb9ewzRWvAGXv+0vFUJKkJfulDaW7O0TJNprCvnGvmtw
jdsSXw6scRyIcNPCydWysoCXJ+Nc9c2EEEf/mV2BqAFWMl7/wmveaDAUGuZ1moi9
S/1pPwKIWRS3gVxhvmksDyzqf3kKRM7u/RYBBYxDXolFgJpvklTFhiGNzTaBCKdr
rldbQm88Gh6HbgGIsC8ZJqt/TGWhyoXIawRnMZ2ahtRwkPa6+MjbslxlAGzwbaNx
fYTavnUbMZ2dTCBxfX8VunTyq8pC17RNJErhzEFjyBRy1EWImlquNOzLCa7DJOGi
uYK1/uVv+nqkFQMxprm8UHUlPXK9wUCNO0xfR3AjiWYb3SfxdXYxQRZyhLxhY3k3
X+JeiDgWK9FjJOYJTRqrBILoXO/1fQimAVC/ImlnfhTH/KFF31ztMJ/Z7dg+nR60
5v9kUdhqrVeTRwBJjoi1yReD45ZzI6Egp/cfFJzdjaVwFT58BNaihbVBHpt0S76V
ZLZyHFKh6pG9JbZytFuYQZpB0ovfpjwqVF71XhqnjpiM+foP0WrBB7PV1BGVGnT1
x12ueKjnoOmLyhq8nxYuhUNgVabwTPhrqkLfiACpAqW8N9XQSb51UtOtoGQpyrOp
5NmwZH1G5RuWwyOvESHmoSg01h5fXMIIY/kVj2yReSVtgdE17cn1iCqbPFbDpKTD
WFi52hApN+cSPP8Ihyq9a7DViSmIlYOL4ej9569WhoLloqvxfkPJ84g1OChQpEQD
ThG44BNBDGXCUy3x1U0dY4XjKQMzscwtQiJ4KF2roHlCd53MErtx6I6IdOOgFZMu
OlJ5v4eMGJkOUh/YCDZq7sN4ARAOndmymW5bbmLMATK7qlypI24YLj8yG4sGE8gl
7cXiLJX702UPhXWMZfc1+l9GYBM3IdUao6tVPACclWpwRf1AKmdxGuzYVJdaVP98
rwn1ZCFc3d1ct0+2fKKvl/7N4kR0jlTGY+t4ObgpI4HWxL4LSaDOSOvwHy9Il3/2
65FmO8q6zolPuzXnbpuI5Z9eqeSCliwmrQCzvjcM+pIRr6+G8g5pKGZ7ySajXxXj
orbRUhOUXxFxCCZUn5YrjjTGQNRkb52dUvWSqMxVezWPP+iaHmcE7DMcOgSBlZ2P
iS/aNEhOcg7VgEObFl1RZ/T1aGTh74etklvAVjPmHTsKhryWTQ2XEr/7f2mEFCZ8
mWqNs9hGaVywx77sEdei/PEutV0pYBAfxWeLuRwO35gNXVOvrMdlJ5gEAySQyhmG
NPL0waQBTcx88qlZHVMxmXCazgLhWHMVvJR3cxsHaTuoemeEP64snAv5xOQ9pE6I
rVFALqyMGlJ7AQjGQeXJcVq2mzt9ZIqQkFyxWBQn2FXkuhvCSRWrmiPfwod6MECH
mHyQQ/zATh5uzng858YMwWkSZiyjcH/4vkHKVldjT+kwKbl+EDxVPCzl6YYM2UQO
x4DZ7962e6l/q+SAbDkCMFuGUtaThOcAcxeKw7Wnzl2BAuSG9MhYg7U26kujEDiv
iYEYo0iJ9nS+qhP/DYIDasqgb7C5Nidyga5hmCrDtP89aQM4L+a6ii6vf2urB/yC
I7JjjWRczh4XwpXQ+iT+b+osFygDl3BGvD0kWeMeHPZu2Lly0VXITSd1P6ROEKNE
AX0kNJhy4/BKswmcH3xLoj3d9ObBQjh0gIgyH2Ge+hYaYgHJMtcElAxXXeS8Bq0b
yBeHgowpaNfNF1PoOlBFFXzQWeobq6T23vEYmwiKqXdO73Ii7TrpTvG1j71+J3q5
+HgXCz2ngKl9ceNLXt7nyXzuaprLrcBtMf+j3UyEf/NSYp6tzlz8XSzfPUWTgb3U
f6NVPOlyTbChg9lUqvPQnhPsK1kVcl9UIUaSZIAflAOz9C9Yxj1pwq1yKJSloWTL
FUHCbV/DVEGlJf4cKBfFXcdn39exHk9lSKZlMGYHmyjd37inRgicNZpC5eH4YHNI
Q3ghch8elpm1c9fTupNYDMXt9MXRNQ1rBtyQ5D5QW3vJfEHw36MGQszbRb2MHQmO
RepTspIeZlKwSIjRR0Q52RHHnZ354TV5Rvrm/okykgfy0e1K0Z/HfcnzOpENF+Ux
Nwe8lPnouFas0oqHKnUFBJM0IahJQwRKCyWK6GCobp5n7td01cjKLYaOIWw2kMmg
j/j9R17SXKQabcNdkrUyGVycYP+ZeHJX77k/7Tw14xIobqJdvEdBKdHnKDpjebXe
/AlORLg6EZXJOxgGCOVF6zcQcZ4l4+GmH6J+rZ2CNKOKlvQ6ayPkvIpXPmEtdi+y
OGiIKolxDeZLKp4TWDuYd2sW4oRKMAvt4WVoc8iQWhrHKL73mmh4F3NrlL14UplQ
VT0UcQLHgEbOdHisdApVLR/8loGCofjX9lPoVuefX6/F279WKFhMKm+yLfrGEETi
a/xgX5dUBUQPp7FXee+f/jjBQKGs3qGBiPthMqxQMaW7LGMKNSOH6hP0/ZTNExri
i4JxoLXLx7g8MMMuwq0ohbq/JOQQMYw9f6Qp95A/LnkzQll75g+EbIzHK+fyaxNn
myPlUMJ0nSZvvHotBqQ1LPrmUAIoRMK7dlzhtjzHefPjAYDfFHn9zWG1lGAAXqEF
XgjX9KLtLJq48dFcf2eKPzjuIokjYt56BHs54s7DG/aKT85Mj8FluFzfwGxFdDa1
OcJXB9bWyPz5XZh6EI9xxO+Oryr7A2UzSWBsdO7jTAu5HXNbsoGXsuR7mVRfi30U
Tpd0pMnuUNt+p5nrp+Ue47ExgtCWwZ/Hkxll/2dducIcOcLOa9O5YV1BHy50uhH0
owZEhAIrAVbtXyeZy+E2Hi24qo4cQRKNMjJzsnSdfAoAKAgK7cHM+WgzTCPFAAyj
VnfutS5fnT2olq+lRTHbrWWD6d1Pw4lqgsxTKKLnrwudzBrovYScl02tZigFWMoD
FaQwW6pdw1RsxNhN3awWAY13EicLMtmTb6xkpSKZwWAkaRq8K9JD/8AGe1XjdLrb
qwuL3WIkC7shE1VnYAkOL+8cvYu/C9algIS7UglR7Dyhubcos2CDLYrtsmz3fMU4
tgKtEfEdntydXJIHUujf5HXNonRvcWgUllDMEXMTMloOrQsiUF1E/1qa0tzzssME
vUgdwfIokb+FAmh7s5twdyWcCWMnQThtpe7U1s2S9cRiegDahTHzjZNMRHKTsIel
Jh0OXf0metxdTnhm0Ao7LYSx899YJk0O7VeT16h1hXNciMzQZ2HWkYl1OUjx8hZ1
0Nq+DYXrXFHP+yZuOQrXDFT2vR+PBPujbCnPDtvHUpxWqldQF7Kv7F2Il+oyTtnm
TOO/m6FwpD0dL36nkGx+X8OhFC34T/ATBq3FhcTe8sTc+5Ncu89wUDVpCjh1FV70
RS9bax/bjNpbyAps4aiSktlNOGLwTTB59cchbDCEO9763U5hPphN9RQDrSaa4d9B
fkARwR61udj0pq9mzo0qsmq0wiU2cUzZvX7m0h8pYVFt41r6GrH8Z/hxW39H87rN
g+B5Vw7DsU0aD/7ma7aEmE1zoSjdi/tP+gbMDb5DH366QNO1TBfIDAUIFdx7aVwQ
VBk0u9fVCWC4baBfc50n6iXvbG0zNzFlCH7Pw/sM/Yz06PCLk2prvif9Bfe1Pbkn
cL4DAI6Q8GPG0ZadEFRUPwjiISIxffI71wiNCqW8wZ7qFURTGjyGYXrzFPREn+47
f4bkgNA64TweWdWrSVmyfiCFb4vVe44ZhBIDxDNnjdHUQk2wgMjDcRN6vqhf0BVT
VdKqT3YvwR6CqKqkkJaQA1japlpHUJdZdnts3p61oykaUtDHQZ7iI+PIWr3Ykf9P
U7l/490j3R9WkCNypInj/1N7VnZg8h4XT/2yWOBjqN/9q6qru/EQTWfGZ2Qbpqvx
XJIiopExnZrL1i5jCe+uHZw6dIWPf5ENk5rKmkexNmaS3zSmSmOyTg52TRzhrBv4
4XhkNBFlUXJftO/GboUWFLNmqgS4DT8wblJ7Xz90yRG1w50g4Y+6jJ/buY+/hLsO
MCd3KNQ2o3Q1Gzb2nz1l+jXAuLLii7crZ8JpvNL0CkmhEWnRFr9rGbd1v/TQHInV
D2AlfI1H4XQVneYeSHbxqh/eR8OxMDsoxEXBQwILINL87dl8RHtXUbMNV+iTvJ4s
H0iZrSRi1eWFLOYv+u5CVuNResZfhf5hfXxJLObak71BTRJPhv5mJunjOGLmVy+j
KcaN9MY2waxbeDqAO62SaGp3Bq1c1It96RxHefdEXbB4nr/n8k7Pb+P4zhAjfBOz
TpfeflWX4hs3lPOYl25lbcoIcwWtx3QizDs7akiCYV4us3jhyvx/9RY2Chljg1rE
3XZEVg2JiyEX41PLjCHX3OkydksBf7V7ds+rEHs1TWOytHWVJqmq+xq+Ly+orGli
2bQXDZ1N3jd4tZ8voUm2gL6iwdzMB4l9DYEf0D6AJdHfcp9Gu9LU59DqwQSkEwaP
n7xiCDP1KlSa7VBPqjDA+CxfqNVeuE1K0dm+iK47x/27zLEL23imARMGaTDEFX2n
dBJC3eKfbDl+EMzqCxafvWoliopLbV/MtJSYSNrXYVs3G5OTyeduIj+82xBPmXx2
/b2iR5PoJlVbMGJ5ucNS3vuGmGZ5ykaI6mTuqSmzzRKhD54sAuDzcmnJ5Chlc5lH
CLmEkPvvFlxn91azWGV5Y48hhTB6B6lI3VcgBugR65/szd1LlT9HH83eVkSkC735
9i7ovdSLuY6P3oXOHCZxtAdK+m8MVlVuDy2JblhhVFv1WIhcBE9aHrnfpLrO/dYQ
BgY5Wtbiy0Glsyq7XOk2SlGhHYeirPucMp09zyLb1I6uqtp603Qvl1RJ/OewpjBk
lXPNQcyJ4bnDPlI4OlN2oKipeAb3B+CHsazZTPacu9y0IXpbEyIcMqi6zlplM03b
w8GL0Gx0azUqNTBOK8sIgKf/+UcK4Z0FKGp0Bhx3Sw+koOuuFMAcx4m1R+cyWkqm
sZOzJNRNPf6IHalAJ8o9oTzMFqULEb6Bbxzn+ZoO01rM9hP1jOAIMcslGYO545Wp
meRfHKTHGBwvc1A+YYnJqrqXEi5fk0pvearXACouuPGd0sqzbk4FHUkiQvdy4JQi
/PDGNUT+Qm1NQzgooyndn9IrhlketGgsuIcJcLqrXV9BnB58zXKfHzKlelaTuuq9
/4VsnQBi/WirWnS65WWns9ffBIE5lCZ1iTdbTsXk5jPkKNtHtOLaNrwVOKKRLvFA
367ftQQYCF7mdRRlTlXvWqtkvr7qbgDL9d9407XzEE5H+oUfgJ22o2LIKX72V/jy
hZjYzeNRoV8EKHSID9XN7YnPaVoWlPUDNLSMEl7EFmF06d/EU136zY8nSvTpCBC7
ne3iu8TZXtI78t4HlphdiusaFmXbOzKpgtrWw1tL86dirN7nDT/uQKFaMP9tRiwT
SqBT8gtMGlvMrHR+Z8dXRpPBIyemnrkjC+vmUhGf0AeqvOr8FpyQ0cyDaDqVx2FR
bAgoqHIAUlXiclfhle/Se7ecKbwG61aLscJ17cAbFC5HmGJzAlwumdXa60a5eWPh
jKftmy9Eej0oqdqi58l4ZgCWVuVbiOTRS3PjG7x3WxBs3CNAKXtFho+Meu53+SAd
uxz6uPP4OGbBhA79H+ASxzRkEkfU6T6L2D/qaYSyDKQw9mVW8iqT2JAgwu9qm1DA
Fc4jsL2+QDKSjUAypM2/S4bz7CeGQrY4LXpy6p1GihfztRRGtvu3zeEvV8IGCcRR
8RU46OAuvl2BbfXK8xrSo6PsTPCxvpv5+eRLxvzwOOHUf3uK5VHwpKZQCJuxbUwg
zO4T2OkqX/TX4eyM63l2Nsq8AN6No+Q58ode5DaWlAVkJWazCYTeIU2Jpzlxzkj6
DgPLqonOWdTwK85CUprWtdeFcccJvzLt5n4Hp6/UAW+m9wHtWX3flqdnGlb+nz5J
BCLwJqyxDvr2/UiS56z9j7OMhnE7y68/RvLrXz0cb318/zp1lmmuBQo14ZcQLwjK
r3X/fNapbiRqAqPAnkSYHuRDj6eTsd5c2P+Y/DnlKeqeuas4mhikT4+bBuk/ANNf
ji7+t5RUiCwhXxSlutSwrhmwlb4VmpERZVbEiu4tyUH0D3SQsHXDFw7KsC3V6GX4
XG2i+mXcoJtjipdwWuWP+ycBn9nLW/BaC3JjUrib3oVLe1lHB3KcvuZC6eSKxGHx
mOkumK3vMYMIkiZgxWHork7D1bJaDjEoEkNmVwE+kRjCq6Ni/EVUGVUT9VAh/8Jf
qQFUxrSZnHm1zxKL7zLmAAYdp+x9Qn/pYLthldbpd05Wvchf4hTlW//plu/zdyze
GQ8LdAbDJ17boX1qHaLNCX7/QAfkkRp2nGEIzkp+f20t255M2E4C7iQBb7klFpg2
XzLrmza6TpFBaXVG1Ggw2mGqICjAwAXW+ZPUV7oKlCsT3C92nHcV0ZkrdMisyTge
ew/lOzZPZbJGMo24tES0Erx1XtQY9Vf5q+zn3bR9f/i1aLfuHWDSU9tKEniup1Lx
iW8kR/CnY+PWTYk3SMIKScCmsBURP6gnsbWWbjcumfoSqGKRxODkwAneSCyoYTIT
2i6xLaOnIgNj0YlO6EcmVjBcA4txcKmjo/66Txg91A9KB3Sjczq2qFlRwuKewqBa
tsh08op27UWU0uL83q+Evc+vuqi3HdBD5yyb5KQinmZOOxdUaUfZ//x/Dfr0UJJV
LJ6FmszEHT1GJq7dhXo/zmspHAthmpeGuWD4o1/krZLf9a//xTyD9ZAQUwnR2UoS
EWf+rAPsJwGuehLlR61Iu6+5f7t+doJ8jHjuyN2VEYqURTk3+vgQUcH6omCw/eDk
RC+TjLZ61nAsCueDUljrT6s9uFvowL+eAs5US2aQ7gzpeNn9lTVW51WktsJJNmo6
g4Ushm+fo7fzb1Hr+sYSXnOyGnTpE1YKJ0Oy0wSzxKbKNS58nY45x+rL2uvN/0RC
iFHmWNKXU734tlgDm+PKgC9OPV0FDf9aVMdbPMf+KR/nR+35/9dCab8acASxIMkz
7syFGerkV7oNpGXHTD4h6Hkmasd2y6JIWvN+CavUL4x+vvMq+v3j55HThynUmj93
ffN3wZ3T0lhVqVElYx42bF1BX9RnbsEbxyNb46/7Ld+ZMS87K9RQLmXleBcFYp3P
RqVR4d4jzdIr+ZGlIkzM+hZysa3irtqq3zc+pDBnfGbgjbtJEaGUwXuI5vXNPzUF
T/PJT0NICzWjCv+DA4rywRCxBNjYYHo7A+B/SyUzutEkQXkZ6H5GGVLcK3IV3rM6
UpJG1dPLEMXGdtB/UXQnrlYh6CHt7xrzROTbdiinBv3CIdyIMEitfUwuQR8dGze9
jGDOZvbTHqdCzSvg2pcobWoh0Zi9uKFqjlruQCfhqPNP31XS5/0Nm1G7cwwjpfpO
7e9dZepOFjcfQS38bU76OZgmo4FT6Y08L8UYHNIBCjs=
`protect END_PROTECTED
