`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1dmYN3A4Bo8IjDAPU5crS9p96iWb/quM8J+as2M+0+MpWehDEdQB19ym6zVbXGW/
G+ccgO3OgD7Zb6Xi3tpokcZ9rOEE2FToZADqiSN12kmr8euYCo5dTYSkcnQwTMzp
OCWBhlu/npfNNcyTN3fv+1fBk3Wt4+rcZnvUFqAYpHZnlsuVMYzKxuwgDJJoI9+m
BRXYgIvtxvAF9wZn1zViFngmIRs7oKmVZXq0VSm0n6U1iwBWA7S30eoCG8ODXh0d
Tp1Knzv3njoPIDhySL44lRXG3CInvocyl5BQLtpkqRI4wXuHoCbAV2oYs1B31JSE
+r5WDLFg2MbEAA9RSo/MPgBJhyiVwUomMa9Z/BTeh4yd08qqq+dGdU6ZpGPdn/f2
N6kaGpFyVi4Ck2vb5o5FSCNkPkHQFoM2YBTWkv1HbTVRtK/VIGOGRwIHWjQC9TsG
+M8HRflEw5tnnST71wwdOiWE8ydKaf9IpNBymW7ueoseUgcNh+LryJqaQ7IuYrCO
Ea6f4kgercegg5bDmXl2bVBheiD1JJTrbmBN6CzuQDxXoblr36qGWQvxuq+SdHJC
mgl6/Kd/cw6Z9A5nP7r7IP0cxqV+DQVLwRbbo2eCTSoPr97YNp4rKSypwEMK5pqN
vjZszBi4fk/wYd9xK244I3JimWjyqIEQrOwxFndOorJGZixiK/kJiy4VbXgtVZdV
TuKFqy9Zct7/9Cz/eee+dIzVMnP9stdSJ61ae+f+Z/sNOSLimwlmHgoQsdyq/PQk
6/4Y/RpqIWrEXiKABAHibG9jXo9bf31S3zV5/uyxGP5lzThxqQC0nV6cJNIPJBHd
jtqSX6pWW19ZMMHQMLLGjEyBb+i7FCH4D8z5Vxiy47rciNtozi81zfGFxXkcLM2E
TU0g0YMmy3tnZPKfCtGDNp1TnG96HqfDEtOjKGPpKgYLeXkvR5pV2qRfghav1ycF
iwxC3wTze0UqZIiskZAqqBiGbRtoQTpM42G1WiXZeinzn7/VRUxn0jPkKG4GcwyG
mGLofls17x31PxCJ88OUTIuawp6/F1N5jjp9GvVuBkV1NilAMLMMd6Mr/cZ/Nfxc
VaAcjFqjDRe82i0DOJmlLaVxSJ6aDMXjR7zAIb0ob8gXlJn5AkEIbPUXG2OCJZR5
O1QgTkpmbIiK41+sQ+ICfD2rzRIT3KdmialbCfXawNMScmwyYz2MSZO2vJhpZ8od
WRzShxRh1J52CmrvWTEm4Dq5Jjahj7yhKAa+aEL4LrZIudmskq5nrDWG25wSDfFf
lvupl0ErMWONEV7wNphQY8MrdUNjxalwxuSpmBCdz0Yzx5rdYxAs524x+ZcYAeqm
QHAS0RjdKIl7UOsviLhY+Kos3LX9bkXkQ/xoam6KonRYVcxmbw3Kgfk6lSXGnbMx
h3f8CHGex+KFIewBo0PL+0L/fWE3pXwwNrwmLe/1WqcOXodyv7cLk6XyuupQcXQq
hs4NIJLJ6dD9YJPTk68xqZ9Vb01QSOXHDBygHyStaVnEOTj8GPgsIiBWlEbxcSyV
0+w/caFs/qeyNHi+t6PLIJc6T8qFUF5gTdUygGWZDSmcoueyJF14tPxGnhqZ0rRG
Hwk/ZV/c8zCn9u6wGAZnDr12MqLCl3L6pK7weXl92toYqwvKOm9XwMhiBpOhAgga
HeqAQZSER8vIz5lfrAD8FpUWO+5Fedizni9Ta4S6DaVhGt/wBMgM6aJrAlONjNHA
hqvoC4fmND227AU4wy643Xjkaj1kXlU4UJmlWAZm35hHThMobwtYITsiWFD9Sv+2
bcSXs0Qr5N9C+/6hRU2Pmmmel4T8aGDYSTV4QBspMTFFR3uWMwXBY+BVgziiJ2iW
FsKzrrHHnik+1ES4iRihOrTu5Fp1xFbxKds8zXr6vfqneZiUQOnNz9ReDirCbLSV
JfSrRQ7/bICYTkCj/M9tFLFB6sM79ufbESGbfKWWwzgm8QNWBBARLXBjJPcnN6hP
YOx9cEoj+O7wpYQzZJXVJ7ivNLbiob24L0jxAS/69XbtXapndCF6GXew25CVJm4Q
31aERgU57wMV5rscDANPF/g7d/rBpLUs27mhzaxgF5pjDCneGslCIsCl+QFQ5BcQ
v38kcjx0eyJri915GS9MbX0ylpQ6T0OmECUMn/auv6Seff7hXcuANmCJ6YxwCH/8
RZMjWaZqcc9K98TzmkGNhokAUaW27T6Ih9/zAwNn54Fwz2ai91R2WcALUMt8sLs9
cv6NLdsUx/JB322yts3ZeFaTBqkNeQLJwbX9jbUrQtGnskZaR0QgQYpNX+ruoA4a
l662pXr27iY2L4xbeqolya+dYYuw/MnLiLnKficrNAsQ/Ii9816dO71fkcavrCM7
YWpfJXIArOn5cqTY85erCXsAmRXMMo+EymBqQKNwpBmzE7JvFe8MMaRhN/vM5+o7
/eKklDDIvbXbe3hV8Hpmh4/bQQHyU6DosB+K76KoV96tkxTDUUmueyuCKD9lgC1a
S38Xo8xU5Iit08xN+E0OiyNf+SjgDO4+XU8OWku3JlvzDcZUZSuH/B3a2lAIPbai
cVVOLPKPun3D7atuA0rYp2EkLtU8GScVd2pqXd2yd6mea/TD3tfOTOEgqK8/AsJr
mGYqrfR7AWzzADlzAA3JjVTtYGmzNNrdg93dKVkxXgGbSEZ0LJwDKXJgi7DcoZz5
lvyzMojIzhc56TKSMrYpK/7y1o5A8GISMYWQZAH542xV2IVVLSN7S73QeBWcKW5P
`protect END_PROTECTED
