`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GAD7i/kg3FL1KsW1uKeb/QVNK4TNqEqzCN0klwUnEpV9DwUk106OQxC0ht3fzvu/
IflUaoyAyBxWOtkndeIWRyP/jwET2IKWKnHhKz7xt+SMDoWCiKP7Xj+4UL0p+BQg
BvA+mx9AGkZ49apjkwAwJVMbiGkV+rqzG4QVsDScTQ4/8cSqPoderepDMeyFZNsv
KEqKQMcKkC6XGcFQXi8y9MX8k5IdA/VEExmgjfXV/eCB9TH6iz9L63V287qiKLyh
beqgesJzxdJR7FtawQNJe2b7wj4APzxVjlC+ASVL/m9Z38BPmeNw7zE4OyWUH/Ro
Vn8S+7wRvZ5oXkS8EGF9bzbaFAjcfxixnZOAC1PD6ase9aKdLDWU13RkfHZLU3Q0
YMRlkGPSi7eNmCBy6cCDI0BsNlS6HNCvNGNKTl4qkc/jZPaUs0M4ddWweCM2ZEad
bhJfXStKLRs2JOJviHGm12VbUKL4lIxDlqPd2gwqtBVm5CrS4IXrY5lMBBehgVvu
7FSWmRHjIfvyh2ta7APSjSTZBpMvpFOqlWRJyKXl2/EOOm1o/4JFJh1F93ok8gIC
zUMW4LlIaA1qG+naNfNf7cLn1eg7TFEvZgFsC6Hs4seLmzXx6aXp1owvSej8g4/0
YBP4rkGQ2nbTFtfYqvan4yzbB3DAq1H9w1TfNF+ksOdxA8QMNw5DTzOsDl3x2cU/
ma5FWXlP/+hGHKEquwjzpJBxe403Q9v6be5skXuZv1XyZ5VNyxo7n5fUkRS5xE0C
bSN0MoK1Oc0n1s1t0vLG0WwKwREHghzilCX9Zbe3qiGJNnjGqlwmyuV2l2xmzou6
5YI3GqW0t6SBbyz7RLWVQk95jF9Fdwb1ZOk2Mpr00U0S9unGkJgTOXXHSgz3iAi/
`protect END_PROTECTED
