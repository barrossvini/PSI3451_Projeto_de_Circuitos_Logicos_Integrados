`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PRXfsikxffR+FbFwJKo2ovCIxPCMscPMtZfR6RzyxhBB3qR5dv29M5riBRSvzk/r
e7ap4n+8B3jFeHnFd2K/YBpzs9aNWdJFu5cqJwmFYgUyhvJ6jWPK9Yl43ZoNUs4N
Yu5DlVlm0Hd3ied4SfEWHYTflUJ2WbhHVHFlIoSgdUPTGYRGLMnJ4SVJOtwfl2tI
jOW/rL00A9RRbiuVJdvB8i7wEWbW/KQef4eAzSqKjIYkdIBQYgb7qm7QQegdPQfR
/ombuQ6Y0Ij7SXENjUrDSbcIBNsbQtW/aXHLlbXTGwGU3cpf6rToEHrs2tSL+aIY
h2tz7iVSi5ySodSahKDehk83g2/h7lazSUNjhN84pdiKHzcyHvYXVHEYsSNxQmyD
FdVKsTL2nAjtInm0eu9z0ZM2VFdmp/ppStmbe5ljUlVBZviHPDsSSDqlU6jz5P+c
W/g2W/3mYT8w5xCNxctQMYDgo3490PSkmsHk5OAjfrqoeaGl7kNSpHZu4Oh7wOT6
EpAGYMr4ytjiG9W1DlKsPiRZe+r1EPm6+eInwjQ+afOt4kTL0mtnAr1p8l1kgaov
W1svBD+aXwdcQHR4xLo1IQ==
`protect END_PROTECTED
