`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aSmgN2rlqIwBYI5Q7+lNEEwZLtuyPgpQTabOMGo6VQc9FQM+/sGAOR7cBq3AcUYq
YTV+UqikMB+OIKW+3zIbUWgBHMUuzcIgBdGw9AFqhZBNWenIZY0IdjwxQlSf61h4
4k/EelkjfI4p0W4hiIRAQPTJk1zfpamtz0hFf1aanuNBFMhWRX2psAqaZInw2lz7
jFzqb8mTT2PnCRsCBaOQPNE/8fOKwipTtqbP4lEruDlwBH8CHLtR/X5XlRkl9pwE
CngGB/tzRvAO1n4hvjHhgztacc3KOiGS2OBg700RTCEDR3gI/l2cJrJ1f0k3R8hj
NiVJA3TCQPR/mrLY8Y0UVPEY91nPSmsI4dskVP8E4yUR3pRYB9uuiBrExTpADoEC
`protect END_PROTECTED
