`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ni2KqKAVknRd+SpRjyt/vybaos0OCLfd3Wu3jj+pP0e86mt2EDaGWgrxeGf0uSaJ
Q1E8xrfATD+dFOS0itM9YI0GlMof+Q8WbpclgCegzqBYmMbDCjwOiEPSHNdd0z/+
+jTitFO3EizesKl9PqXWI1ta8s2rVNZE/0Huw3meRS5e7W0NcNxBYrlkBoyxCjSY
3eI/ER+5dk8MrDuTpdzDcUI+y6fWrp5OYG2P4V9Z1MZxDbjLpaFFA32c7+3kRFxQ
atOxRoQnzC55kebsWpASVJMR8hmUS7niGiuBV3UHwfbMGyBhu6qWjstbJZaaz+qB
/X+RphoSDurRoUc33YpNQSSRhPx7tBXM2SVNnZNlGRKICsy1Owx4bUzh5H7mn1Vy
NEjb7rsGYkBF/x6bdhvjZCUY80mQf44wGbp3CWjWkwmzYAr//mqoeuCBZFtKQgLQ
YKcumKY2XfXs2Mw+JODV7dfBvJ0Ur+eyl9ik6OAa8NP4ZJ/QEythKEPFy6wPE4tp
LLB3BL6odTkQFEEUxAuDK9COvoxkrv5zINy/y1RUW6M=
`protect END_PROTECTED
