`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9VAFIoHApy3RIMPf0bzixkIlU/ZPfaV1IV2ogQzqZ64bZTe6oXTZHREJ+JCZk78e
qxHDwiFfDFuZRPJw32c1QQWxhVz7FQuNrMcUKn4XqUOd7ZOeNoLZKLJS9nQTgjNl
hEKNoDnVPNWPGfjKcghsEY5jUeEYVrdd1imKDDZojstIlZw1AHr/AJPGSkWGQw9o
mLRkwAOvL/cytBz99wy8AH4xxL5A6Hm3eqNyI7y7U1JsLeUcfyMVoNydPRofDExi
UuWDLYwfqvx++HCS2wcLCcDDPCRSipmkjfCpyElz8wCtXQgJnMW9vjaiQGUeDgfm
kxSMDHwnlAvMOlf3RiTe6ttIDyl155dVYGnQjRHX2KavWWZBYotP4bOM+MsOy5xN
qX0ZMQD1i1y/7+lOTDDu++t+LftofMO0YKGZ/6AmKqYlE3eAGTwuE5qiu2Rp2qhl
6vUYJ+P079YELEc4TSu2mq17R2Jdz2+jH4YMd40p2v/0NurkznwLJ/SvePrIDFXv
A75jebLsUKM2PxUQuXTHRH+gPxbUSM7tLSHU9wVX1WHIsR11T2j10/5KGhJHxskN
6GW9/2IVMV9oSMu8/QMr/z4KGcKoYCShjaaFCT9fbIoDUK6/W0M7uB/1KlPKZ06j
En4EOosC0a2ushDllYDWZ7TobG/GsvNXcCdPBeRMAHLqLAfEjr7wRl6LVFCz2y9n
`protect END_PROTECTED
