`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BQTaQtzfBiVHwHv/vh0rMmDQGy35MAz6+SsZXPlz+6FZunuq70UMErL3BFBRk7Qa
hj7dytzpNc50ItGOxXIoV/ToMN6hN7Ra+WBIp/5fJtkkSVRbiNT5ndJ3S4UYkTji
SzREH+rXV9HXD2zBGiqwYmKsUbFc9CTuzUTbfTv3AoCseAMioVdDhX6lKTYgdYZp
`protect END_PROTECTED
