`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l561ZVnlcqjeauBInm5DEjgIBn+VXogAy6StgpD/1FO0Qr/wLJ9El9A+eWRTMtzX
FzJ4anRoAb9wTjM0wv/hK3ktNrBEb9Bjbsxlq0TQdeePQo1Fqmzta/0Bx7J3HvIh
FqY6OFmfvhM4CqKFnfdp9q8zwLXbLvtBN5wiY6FORzfo6/kYHGrHW3622f2eL/eC
yv0klxk7mJJiQPmkVJL/4IQ6Wp25Mm0fkhRCRvHDSC/t1rQ4ase2oGjoMtrk5SXA
X9LMrwBGPEsM8NDBqzojaL+Bci5gMjZI+6RYBg1n/oc80le/n0/HlWLTGQBxoL8N
ReOfYuU/dqFVqVzWRWMPNPVZtVwhsArSW2Zz6HT+H8NKBgtJeJGOnQfY4AwHOxm8
XCWsn/hcJQ10XpV+ScBq5+z6kEsJrur8ZSGhX2M7vRFfIwfig/PszF726lAAEHPn
qxcLJBjUBkQsTlnSq5Y466C7/+6ehCfmW+9eYQsa4pM7cXYQshzo22sCRaF77qsW
PB1qM/VmM9rYeRlDs6lr8Ha0ztLcPmQrYwZzUrq85O8uwVcI9yb6CXEYVs8zXSgb
pJuKh4ov7UcbpnmhFP4UmTEi9UtSiZNtXpHbgCbmfEyS2MkL1PQxXjMN/d0POciZ
h33EdDjmhcmBGNraWuRNF98ZAEIWPd3L6jr0c6h6aEww0rtIiG2QWW23Pm4sprA4
RqvmPfx0/E9VEpm8SEd/KFV3lXKQvAtIoWsTGtisMeSqQFuuW5YbeRve8+tcBhAA
B9gbDEbrRcZBBf6djv6atH2JlY92GYxTY+qcH87rpcuNr8rOvmmC0mBxq26BfByq
qpP21uYM3YTSvKgZrjPyJy+6ThMVNnPgpMk0oUTixE2UKrDzsCyeMx1hwTgaDMk0
jO+qpI6mtzBcuFjXAO7xyDLeMR6eFWNk8DSRW7sikdY0m3Oszdn1bWImeCXBKYK9
roh0Kx5y55oW403bzoC1PFicCFMPntehtiBUJcaZ00SV7lzn3evX+t0t4jU106Ar
aA46okEC2od3v3dwB5NBspWR4NSfXLB0qqHr82wyQJ5ncafGzbkTd8jAWsDg452b
+BSLGK+DWTdFYP4+DNRe7DEcyqoNZkqLElotRZCGs+M1oVPAlxK6YZLKorBjZnWH
pPm24nkIXsJgEbppreys64JNANQ70TVTITz7BUFjtEEsTz5jR7mGaD4MPQFwrSOY
AScZOBONVDQR8wSpAmNOcZSovjJJNJeO7xfdvpYdHX/XJnaawD+uqgaCoS65W0AX
pmwAQH734g470PxKU3M54CDxmb/PCFf7kYp7LMCAC8SANXfScoDVhVP23yu0H2Hy
CfLw7AEeTQKzcte34BO1N0XSE5+MvPB5KmlLNFc9E8ZzX8SUtPdloULNT1FGjnaG
IM2BZ+W1dlhL13CxFE6LFNJbv1YfVxvCzyk/GzKICBjbnDHk0z5pBcfnIzCcXkN4
wBmvrq4IBsX0MeOKGaWfhN5XoSyc1GmOEWQV5zN5A6USIeDWHdgnfA+L1VDYvjlc
LUjdTjRQkGWg501EjN8JJ8rufCxCSvHaLkdP4Lxu8zHvpWWRiEXBbaHRiKIWtlYm
V7UPOVFNT/FYSXsV6RQtZ2w5kMqwM98irur9K47ZB91MruPBtUZkNuvI8NC68ptz
45pZPpK/KjDISYQ/OY7KuQp5cZrFvRhiKGwSPdV6fM7AMVnESStDn3PUg+JcEVNK
kjxCTrxedutAck1K4+JQwk6BGVgMoXMcEWmTju77H+hORCOn0sjSbG54K+k0cEn7
yoqOuvkIyfgY7jwOeIUCmPLn4yp09wSFEtwP0pszc4+IJMrK4mpGj3/4jAGxmPtW
Kp0Y5ANmOo0Q/VQDk6/iayvRU0ae1n5Tf9A9nWqwn6kaVvBf2Hl5EGAGLjgsNnsL
ZUryq2ImEZ6BiVoJXE7MttlEq+PHjnrsv4iviQCV4gL25Nzb1lawtiXMWxt4ivrn
C8r4HwFLRGiHNUfy3BQBFZ8SZDMIrju2r3a3USmK2cdBZNhtvxBW3IkHzojM7LYA
oiv9FAZTZd4jgunVBtyvf6tfhvUaSO0nLS4sKs/SPjZlbvz91eVGgTtLkr1Ku7zL
uK7Lb5qESJ5NoEHwgt4PQP+dwtbk1wr2DX9tozGNlt7um8XAk6rd6H+I1Y2HJJqS
FMQOXcwrfli0Lki+3UEzJ8OOK9ExSupiejB7hdNAF9tcfwBmwdqatzzTSKfLb+uv
pzWQBNoW6dlny2pokw0BHp56/ywLFrz3I5oFzQQJ+ve4sEnACK/nz2SlF1d9zlym
ZT/Rko1d3Y7Z9Epfuuensomgk2IV1+pV4Uhnt4P5CLQm+ZExRC1hiXUMRQO9CsBJ
aDhvxi9MZcjdwBgBfAZkSW+8Vx/M34q7pCjcSm1iQk2jyKotwhCvrB1+x0Yg6yvD
yU520rWJdJfarE1tn+aG6Ht4vmxNPlEwmSj/KohsP2XIpXYN4bsbuyZMLA1H/Jbi
2b4ipzCB435LIGTLWtj4NtRhCii6QU4sOdFOWzvT8UkKtc4Mw7ASrLqR+NOYXnKu
3H8SoVUOcJ4DfCh25WreQwQiYz7kqiz3wdmAEm+qCRKBYKufPYjUkJ+o/5emQxI6
uKultv+N7nidkBUjwBVE7bGJ6mVaIkIIybmtUG/ptMEgJ7G1sJxG/W7ftFnBnqgq
ClZxp1NO47SLsfSupWCzbTFA13vGpxwNcQBBcEnvRW36ZeRoOJKiDx2skGJEoKof
qw2vnUB04SdZdrEgVs3cbx8fx2nIpiDfFC9s0vpO1GnVoleqRx3Mmdsj+WtFVrIa
1qbzvp69cf9RFI+g2sZPQYDB5wzG8oyhmWKldjaFLTaTB9xTFuuVneoN6Oqf6HKp
6Q3GuSsBK/SqQTkr66oJQGrvK//2MQN3OvEJk/vst9RHHBYs3tAV6Cl/1pw53R3H
Lg6JhYE1JBDpeTG2cirpFJqe5t44lSI4zqPNnS/jWgIV8dHqh7s+FYjkrl+G//We
TmlMhjvoNjIKGXJNgGvEP18Hew8Bq/SVHEBQA2idgJRiW7VjPfrjovf7C/qmcIRh
mW4XLMYxRy+mpKQ1pwCvt27ejtuiQb535JbE7zHsmgFKlD1wDcjzOz7q8K+0Bf7R
qCPvhSmlO5IdGqnUDpmV5KmVkSzT2iIeBQs/G4Lf9rEC9LErtnsXoxwRGQ8Wg+EG
sS0B1ccz3QoLqFfbbhE5bfIBRDQM2XFsZc/GwPxWywJD6MI9MAwxSVeWRigqgz2v
0NTXAJl6XezhNxnDczDciq7qSKbkRNkFrpw6qZ9YjQPwLuLkw/kbGlBH4yp9hkKU
SZdTKCilJE8vCEG+GSYLSy+0yd8dftQT442B4NYK4eSOq7ZO16oTVNQeae/hSYeH
APFBJOIxzfyDw64UVYOS8eZpARPyC886K63HE/+1vNG3dCq7LQxcbdv+5M5VKQ45
otiLeTtI5Y7pIHZt/KOpGkTspMBKdKaxDLYumWSWPChFOdAUx3PtGcXWvOmXBePh
6LLr4tcdOlCpC7W1rEYvSNabgR/Sfe0f3VW6rVaF0vPWRsE6w2hwmSoyR6sE4lxz
qngLgAOrylaGBXBlWL0z0nkxTy9FBZcq4hEnPLAHGmzPLT3W9vUQ+FMfvCyYFt3a
wJDsiVcWBSQ6S7kP7t3BNT9Ua89q7VRmPRnwqWEwQUMRvcB2NZGsNxW0lRdjeiYa
0uHtMHgaohA/tMFBwuaUzGh9P5mNHHjfgaFNracPhJIMb0Vg4Tj1QwWwK6XhRswz
plD3Pt1o65E8zWEt8CXqEZTgWi1t3upPb/8vDZ87+yWl5wrQTqFeOM6xunqkcZtN
Wppqv7+O1JvMHPLZBtYgInk0ixQ3XZ9uxCh7Nu3w3ORp0zjE6b93cnLrAvKv8xfn
1+UhmIbX3MROU7GAs0SxCKWjap5DTVGrP52GQjY7oHQ1xqsZmUW9ZF6i2w6zlDJU
QPfYCDp5Wd4NfJaLhEaEquv9+VirsKIcOQFC45pwN16vF32gKfa2sdeiLtTVqeWc
AYMoC7sCamXUP7sQ/YUJvyxZkTRqzSUNmkQ02eVTAiRpXAke0nhHPmmeIAqlpHDv
6bnn4QuVU09yaNsV3j/Nnzz3jJAYViz4redFqky28iDJ2QvsB8TLQqk65biPgJwy
CmpwvCT7Kk2fOBbvaUzvHMN7s7wGkBavd7C2TuAV7iAqrHRHpvg09KpAgnriXl+q
haCzajTcOYD2gfizP7MSv+UMjbO1eIubDTKXTi3oIzxQbv5Xb99n3f9mR7AHPdDd
ldLirprjBlRPRqow5D9nRoCbg+xemJNFwMsX+x2ZVqmNjYBBm9qxGmwsZ8YoWOYm
1bTidrioueIv/7XOPdYFgWO/0YbqfUGXGnGm3I2ymz54ofeW/gUVnJevK1BcAGTf
J/P0gZfycngZ8Iua5oUKslbRzl+jkFmXnf1A0y2RD00mTZCdHWuxCX/HNy5g3vSv
ETgOrJjleue+esyx7G4cJh6xSMUH0zViZMEj7PFJIWVYN19KyhR76RlgWGv9h7hT
9EayQoxCgKAnG6/i9T7Spn+o647mhBZvMZoV/QCDa9tx3DSs4CXFSztfLyWUD2Ek
++Nd0uYPl6lr1AvvnUzzm276hR3Aa/W3ZXoV/FRei74zEwSagT4lSnrVqZEzrTij
l85g2w8NlOpYD2CLdPaxbCa4XGHPMW+XGgaoCUKmKWP3KyAc7BjAi3JxPcoH3GoV
zLwjfsj0XWXK4iRee+67x57c9YD+8McTB/K2F4UqBXnIpQj/I6t66uLrhuKc1QUU
miz+0+wElRZ8e9wRXHDzrryegvqqQNcPtbgNg4WB2m54WIGSYWhhPX0uV7ECW75Z
fTfwpMDPegQRN6Zkhl9pKvYOKdRgWJWr5s08zBfwtYfWpu7HsZnv0I1ZLgNBZEkq
v6bBOtrVS1CaTdwDgqplXHDviwcVpXzJHN733+7i01ToBgti3IYsdn9LZ4J9On3A
uPO4sCwvTLHLXozkUZh+ufITPheJ+x5GX7VqD9LYWN5tmX0kozruFwj+LurF43eY
h18M7NAR2up5Y/RQpSb1QcdvfFUDDzEsOlOBYjPkDBBM2GH2fCqN4Zms/YgcMk93
TGw7ZRVOclu/G1A5RU16RBFVQ5hpkaXVjVo0I8O2l1Zf5juOzmw/H8bgSCPL3+1c
ZjA9K2I6PVB6WAFgNETSduuHy1fbf3LSAYxUFGMTvhxG0j3aas2cZ49oE06QxYBZ
SHH/XnFz1sV/ZEqs/MnBZDmhw9DunuN1x2SulG329rWokSyLJiV8DvgQ9ojj6NKt
HBAfo33mUPM7hGzrwtiYP7EdXvMOIFhZ4DsUpD9DuxvGWtxR5vqs6v07IeiLPrLw
S9mq6GDNqMI2wbqh7WE50Hp39l/sCGx5O9trt0DwIApb43TY2DAfDNxQow2t/afP
C7+dvm3PzotCqA97Et+BX2MzXKglK5fROZQj2UbeXOi0NM2kZOS0uxl71teDLnKc
yeRbi+HKRDb7J1JtfYlNNOkz51UNArK7AjfsdZfXSFGa8hYWkuSBwW6esaSJW3y2
6ArQ3gzaM01XH/iK0NAKPST6MiFQoZQ0gm0mMKweBYOJwopEhVQm0YFSD5M21N/F
ZKuPHfUY4clGU7H394+wJ2ozZtPrLg5uuuJeftZOr/ZviN2azcg7dNBvbyuFo4Vh
bxg95dAv4PNj9YVf3+xHA8hYobeeAPrqtqw2GzWbGd/bLYmusWLcEY6wLrutfu9l
g+0aB0ShxEOOlgS50zRTnbLUcrKocRxD02MlaLnQ9bySTHBB8uHSjBsYFot9Gt4i
P8I5Rli6KoBsrcybf0Km/84S7m9w2iSITYPgR5gf4hPdk7P0L0oVNFQ7zm+zNgPU
QM7ETQGAE+EL8oJi5lmFgnwdKQzLPbImG2aW6RO2yX33uHyl6FSOfTPkcaslzzHn
7BqHRXCftHffbgYbnOKSjMqRNgXYSmd1f/+klVEwtvle5eG48O7as6DHgIRK+sqy
lmTBLaESfnL7Qn5TcpLR8bX/YMo3KKTgTYqsNpuEAChie2OrPgps48Aq6H2eyW6G
fhiHZ8kxupDB60GpRxxHmNpVxWLhEB6YYCIJ1YQQY7cuWZzjFkjZrolZ9EbKrJWG
Xile8ZvxrtUd7XB2gh7mO/7TT/MwDyb2/Hp0h5sP2eVaA55/J61TdgGTQbwPfO21
dSJ5mbML/S+ldGaN/ni/8l7p+P1qyVfsjxWw65DMyEnaHnzVMW26o109jyXiuPnY
TRKWDkXWeVBky4eoO6OGBh+FcJYGHXTSE6WcB7+TE3X0NiZI96X33ME2xkN2N24a
NvIqlESfj7UUsaPZ+awp4za3mI+/hMMLRajR5r63WAAFILzVcg1SGWHmxHJA324T
ISL4MXQalhUH3XQ/J0f5rIALk/STS0BfV7323R9/4x7gSoz3CUv83/xjKKGMRjrR
lc+gOVMXIA5OEL+jt096ydTbB+nCFUFfpomjEwDAYKglmCVigYFBbPLIsiwgcLWg
JoZe1slR8q4TMhggxAuQEDkwZ78h32/aGzBFWxRTvJP+vfpfvXd6Ipg5Ppxt98pU
6CVJQui38RLk1mc/ECQ7wuf/UTYCW2yEFyE8168XfIMx9BKpi6WP0mF99DLlMVBL
i4kfOOc0zLc+lKw7IAyOZWfyTw3AMvuU7cTFtxf0RozBFtvMq2K7a8LgRcPADsC7
/JDEWPQG9WCEPi6lxIed/s5v82T69VW9l6E2XAinL2ElLKkp2R9BrzN+W4KtI1I1
qWe93QPc8Pq9HVkPsMKKlSLggoE1oHhrZzwtQwIQrtV3aWk3AXLUuU2N/q1DD1Po
+ggEoY6AZK3wg8gsLtO5I9UwuJAL9SXOMDy+tIrnw/hA9EuGpRxEIdCKgX1BckJq
KyZcL/lSDe80AlrjP38EKh4fZhjr2amXKdNCz1r9nYBYKCO43SMrqBgb+C8xVpNO
sDcVej/I4o/EkQ2vl7d00K+pb4XmD2WXBjbqo16v3j691ZuPwadQJdxR3fyi861C
i3GLIp0K7fI1v+oM4g5OL0Q8JChD5/v9eW++giOAnqC+IFd5vpoB3Qe9EGF6clpo
Gvaeis4Bob3JCv9AuhUuDgybARlmduGVtnKHwZGIdUXZ2DNuC8zeNCqbgOC+hYRF
RpcvEF6cwzDPWB2jIkxqB9hbpeuXtFxdQ11iN5dH/rksS1ocVEKWLcCvvzKCfjOk
Rx4Fg4J16gneupoAtw5XPE6LaKCefn+xt/Be9Sa+LLUTe29GSbRPN71BJxhNuJyh
3loy2mxQvyygb6p862OOBZEqlx9G+ryq8wV6xTx+mM0lM5aKBmzDC07X4HATJvBZ
4WudaO5Wbqy86L3zEm+VksyIBeHSWD/IimLUv0xA/HNEBhueihUqtoXf6LRd+xfm
JVrJYdgizhRxLYDxmOYfhooTbgTAT+asPLVANVKj6zBvNJv+C/m9oeVtgJaot9Fn
mDWuf9EJvk18LTE+62w1FfolhFAzZbWmn3d17uIkgAHR3W3LhkMYb4WDJYmyaVQK
2+EnbOwUEHYyenRbfYOhoxGImN/18TjaCpAgyL5SAO3Aq39+JMdTqS6eagpPFx+i
e4DC39SWWB4Le0uc+ir6mM2rPfyXkCpL2WIxEHQtspKPTajS19dD0DTvocwDQL3Z
S21Yvy1k66dywnShUbutz610OG3hjDnZfKPQQ9pnAWSpL5WU7ynv+7tV4Wo8KY1S
1prTK+sS0b97QtqnF53bEE50TPX9jDLE62hxwl7Kc0e+Yd7C353E6NS8sd9EceFF
zsOMIm3TgDFsLo9OOtr+j+22kR4n+VmxnfOllz6kNELpoEkGmB1+GnlRkxPwlkLj
+JcRfU6mZi1QRlwBNUCRG/hAZBVALuVL8HHhvg/Pg5YYp81IzVaoKNgk+ABhEzfz
EOcX4sZEmcVgMhPqky28H50D2++liGlYEbemE7PlS8qSzgQVXARFPtQ6xIzbDL7H
f75Br2gR+bKuBtC7zffGlAvifC5JXj4Lou75CtUZ8FIHVLJaoO0bf5wDAXgQgYno
i1X8IDX2gN8va4ZXe1pkxFqyMiygRN/JcT9DbqqMNmV6cZRZkc+TFvTSOGdov1DD
eeK86oKQqr5D79ZeclWyPaNeHYGWpRxyegoFdpsvsnQ3qM1YCIkzERtsQnwZeSYz
/aICJpHhZM+6g/WK67lBzfy0AMioHfRPR+A1cwmgjZ7BDwYQahxe6ZHFVYTbIEJ+
5I4EeH8kDsaHP4Rall092Ddr1IRYi7mMCONmUBBU2JVJgpWZ+1e9Xcew5gERsST7
m6EkQFxoJ59TMyYee2vFrcXULB3k7U8MPkSIQyow4KTbkQCwEmc+WEH9RqXaDomh
j5HfOXZjfkcYUMvq0hhehAQG04G73GPeXyPcxhNzNx46tXY5QZibJdBpoo6Vwlqg
9SM/vGUg/73f+p5+wR/0tHzxV/5TwHKR0lTFp8tGIYZVfsewfqMAIXZ97v6CwRjq
HNfV98I4rgApKTSJ2YcMmwYwkwOBLQSaqJGQYPTG2zsiqOKZnAuD2mCapy1RkyuC
QRlIq5buS/Uj+SnImrGcUCB63burg4LqTEYNpWOcEoq5DuLApETF8GbyYv/ggpbM
mk9V6O5iKdpfwJ6Ty6k5NZwLO0il1NQqNGeMxvdFtm1fcwFX8C+LD3ZcHZzGPNec
Zd5O/5jrh7kJRZihdiIcGxBlXJ9Jq4HG/QoRpUog6b5k770znPajamUHvHQEQzVU
7/tGxKEIFVuRHus+ub7CvNg0+k39uXQJ+8G52GCf+5hnRBm7MtDW4ASzm9sFyArP
L/RJTKs55gP1ZJSvWp98BOoHtPMXrkUulcjx2SKImhjzxLbtSLRjQbfnQ33vx30+
bOGiJtxmbW1Rt4z6l/9oLB9W1tJT3oJSvLfshbdY/uy4uN3viikRknjuPe5nNhZE
YiKA+Qr8N3YW3OebgyH/Np54HQLdx9nQgSIAIKG3nRXNBZ4VhnZLHj3/wNosacZZ
QF0+VnP8i9yqj1zajjad9k1uE9FAe/9GhKG+3Q0Wf7vcdqN249j45m5G7f2RlMn8
tfSgY8f57JOTcD4+b0WMtSfVZhSYMF720u3aOUuWJzKVReGTAhYPU8ttXrzrYq1N
Xj2e2CZWnm5HUkE1AmKzudOWew3uxuTtplU++VLlyMQRc0vzfPzbP2DlJwySrQoI
vlTh9gatXAH57MRbWoJgMmSKvLbMzL6Vwya5Gmlhs34oLjzOrFO50bPVyo98+h+i
4jmO+O0yIcnTlShfjk+S+eiOLGBlgBjdvez6+wsI8WEHPyD+4/NBSDGk6IKr08TQ
s2fFfsi3uFHVVWVeejAKmSQyUumdG+bzzx6wcwYAAOTAO0et82ORjogvr2I4AyYI
Wmw18G8aB7XEDcu9Mv2ml8W+elF5sThGf2Aqgh5XYSJtNpRxoIU0oxGXNlzhsjIN
PhFGa97ToLwaR4AIeqpPdsqFbyaOVomXTaOIPtK4TB8ycr9MFMlrs528FGf4oge6
Cp17j3+6/uctAUyAQXDGxxSMOzt++QtC5CwDsVb80xGn+H1WzwNC3YIioXPTaDTy
RIEsWzYGV5kP8UrdAYivepr2yeD21StmNkSXaCNCWpbRf0gZ+FOCq7ToqSdktlGv
w6avrVrQICdUyJNyyaty6xiSMq/QGL+BbgbAmTS0JD9n7Bqfmb2o6cZ58iOe2wrQ
VwulQ+tgLZyeoxWj0FrslanWSowEJnkiy7TW/DD2qaMLnz2bFVM5OWxEyleehobJ
lSkYdRWYGxu+yDiSC2tglN0VVzGktmi/B+1ZVZpgJB/f2iFm4vj6kIlWQ2nCsvhA
/3Obzzwyt15S12J3qKzLCiIK9ghJzqQ8nDcCXBeNuGyh5npN2PPA9DZm+g35w+WV
raodcPxjAAUQsV6d1E6CpoVfZnGM4Y9qiFEaqoejdQ6VXTTLtPWn6YwXgmDxx7Up
nHGvh3ZO2NhFUHYrjRZRR6eSi3CGlD5bLXfR4htv1IUBE/7yp45aiaKPCsol2HxD
HjVzXwsT+dUjzhPI4ycpo/QMa8iv0C0hiWIVJEGZE3d2ajVWs3f62+oA1RaO4xBs
s9IZxYE4RyqNrdk+QdN7IjcjvHK3469d8GNn8F3jGtokDoPzaBeYVSoY9CSZA2BY
kcqUV+wn8pBgvz3XEOpYUSFeLD3AZVUv7C70WpLGc7o/Wv8jAzqSlLba756IUPg7
f0hcPysKDF9JN42Jus44nJcJZ+qwJ24FSqAfqgW9PwhbF+1aO7NKWNdHg9R7pFM+
MpzjC1dVIseXGw/1+HibxcZVVGf6RWOCN5Lj8hHSkM9SJ24XkaxRAaPqtkTnHshT
Xhr46gugG4ps8juWeWNm48HkzrUdgobhILZ2+o1QTA2DUJZTpzB5Z1qlMawskdJb
0gb27oyluLjzG4SbidyWI3BnFMdzGKk0fhIAZ2sMCOeHcP5YlW+R3EBMfCRHHvJD
Vv1TbpXaXWQGGrWz1OQ7SwbL8ooYWzNtPQiuVCVGCh6xCSuBLE1rrbQL41J9V38+
xHFvl6hnp2PUpYFWdWOKqi0YZ2TxsOmUye0vxQTPZi2sZxb48n0flmEj7VewCgRZ
QteaTRuOZmwUX/xjTq8bd9gmehcVQx8PL+b5lt7rsGYf6nH4EKJ+lmYOyUf4WKi4
VHMh0YOIoB7eSz/b1EbeHJLxhFOCuQAQJ9XFruL7XqjOtppWR8Oa+Jum1qN4nqJr
7QsAoB/AWBaKj/bAax1PNmZIu3gcr8nc7nlYM11nhwXJRuoG62D6TKpp2MX1zuV2
7fproOUgROljk3whpCqYuNxFV9/5TKrX7lDPUoECzKwiciL4QxCoCYezJzYDw78l
bhnqQo1pzW8+QkDr+mvmuZqey2tKVjd6GFze7r5OW8IlDmHSR2MgjmMlG55Cz1wd
YIu1l9I0aVrQE9YKlMGDp++FRY6P2N2n51TI8oEF/wmS61rGc4vVHfAC+egarFPT
JXaANUEI0vWLg2S0tBDfkF2RN2HWao1WLpTXeM6NkDsoqJUtFTKvAxOYMy2HhPHq
52muwDMsJsIlMQGgcR6dvUTPN2ZwIKzhqcfePLTN+o6SOYYfNmBqqu0Lhy1OHBkC
tjJpwsNrbTEasPLsuHtNZvmID9bJuDzKc34t4CS4rAaWUdQYnXHHQuEbaJRYXbM0
oL80Q+WfgRT3Ua8tBbKguyib9qoApZeiFky0QJdIMMU3Wq4Em0SIz+W1ts2tYkCJ
oM8XxOMRs5d7DcSOILPlOc23em2PhCRjM/GS5F1b1KLEgOGENJ7Jr2WJhdE/2/fM
1iQsNPpUz6yg6ZRuKMD1/quwAb3+3C1z8Nr337D5lGztL86yOlyJUCVyd28f51nk
/qjZ40aoJKZSRrsW9PExz40pfwjN4Ltta3KrapZp7oeH2/qL/bJx2fn7s1Mfpu0e
tLmWTa0Y59zQ5NdsbMuZJtysXMtfWuPz6TdnTIGWwA4J0lU1tMDyDn71d4FY69qW
J99tO7kFshqdahjJfb2ucrEc2ejH1ff2sD0oKds020aFBXikW2drfbyzeyuMRi9k
LyHJ5TV4UUhNwTgiyMH+htLZ3MRYdMSa7DkqB6BS7CRH2t9G5lmIeA2IO9czvT8F
iIZDfkxRVHY0m4QCBlBhzQtvF/mnJEbR9c0r60pmM6TlxmY9dXRbl+n8tUYGlCrk
oE25C9K7PJYPEfzIwCvfGCHhjXO02vbq5IMdZv4G14aqW/3B47LImehtMTk3DPLY
5d9eJ0SfZqn1h3hkFePgv/R/bjJda4EMoQNqADBvkPOBqYnxnsKCObwT8jFw1nkw
L7Yn5vr65RJB5WsrmCP4trwo+rmDWEo/6UdgLTxx6AY8+/jG5MmEKx64GRGhOifP
T6XwoEGB95tmxfJstKFLfOR/o2bhSoWeGLqpzdRdnXL74tnLcstqjWPtq6vFKwY/
/FBcWAHRfxY9BEHvBd/uQzyz7HzSKuaW5CR/Cif+I6QC/WL8K8JKGfTzDY9Qtopa
dHQE+R4nnrENluHiqDzrgMrf9vdvRmk1c6KhFQZAM8je29LpjYhx2w5qXMaOpM0z
01cCNvasS3A/1XjXSJ8heuTCxh4ZnQ8PElc45qSICRr+UdAKCOPrfn4Xt/AlESht
KppOaUUJ8BNI0safZZlqKYxNqWKqTsQyIlC2EqXE2qp8I5sNVJq/roxEfwiGz7+T
QbxomFN+uZhaGDXuH00JUASmeA4qr4gyu7F//dyWb5uASUfLo2CFwvyO7tcuxKUR
9DfXM7w92DtqULOep5jAh1GO9XuVCVAER7cRS73JRyJcGQQq20PZybrANDlv7wCX
Hco1vSgy7zXajJOuTUi0Fq6Pmnq8Xvn/PxNaZsLKbeE5Vei+OG29QxsKdoJUvZfR
Mpoz+0VdxNpUX9JsNCQdpZ1H/RpHkPU7gANsCbu3OORSBzGl4eSVzM0FXQZoDbaP
9pWPgNJKrcrFAMVdrhruU4VNIS81g28Vb1ay5eBiAP0HIR14uEfAsp6oH/R6FM9u
pMSgMp0qb97NMj40NUD7f0ghw3JqKpf1BH7Ih3VwhbqrP38rh0X5QeKGDhb+5evc
Jj9fZmvxJMecjWaQJOpgneDESH8MNcCVEFETO3p6Z5M7JpakhqVMVuDQzz8Ljmdl
s+TuifajJnF9TRc0a15kQWdbr5z3IoK+eKmmCHuFwbV9wEg3AJTUwf3/Ptx89EG6
5GRlLsvlxYlxGWtm/gyWSToTNpD57wG66iDASBOKQssjQxnLQShUjJbcQFwlZ6ya
bAUUPPhtTuOHlvg0hZUdZLbCAP7qyytP/Qm3Od4jGbszz37Xj22TFBD/i+ZcGANl
Mo235mYerJfaAGVyFop+pdA57KOCrub952jNf5S+VjsR0/LSqB441ocNyvNs/lFJ
F8W9NFO+DYNev+b+H06dX1yjwX4F9wv1FOPIkwcZL5iERTNlE942mFiLZgzFtPVb
KSQjaJT8B8Vt1eNVjlL7+zkOW/9P781rqlq5ytClXxLYtnqHflU9/biW9xFdcCIy
OPqvzMZZciSE8HRdQCubP6RV7ggAQWeC9EMGMAZHXeJ3HhXVbY3luk/yScmRpYgs
EaCrpSvOvGpSfAfMSvU3zMlSYM/PXnzgmrip/KfH0R1K5yDkFMxxm1ZgUIG4xzg/
Eb399XE1QOggJhrvMx8l2LXHHv0ee5/6hQHwQcGfE8HHLs/BW+yZpB7SwTa+chpU
1Wr3nJPjikJFiApLqnnNVbPoWsvUdsCUnfJvJBbqbPAwfpUxCyb7o0M9+1sOJ0IZ
/xJBP2hvaAN/B+K53wBVCw==
`protect END_PROTECTED
