`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7mmemPPuZt6gUwpjRYqic5RNyC7WL8jDy2oIXvMBzjQ3tynRnZ1JT4T9iLIq7pxD
MNkvt0fGeit4+lYwL4Lwi4O5JwkCtOYB8tZfpOXWIubDXFYXft6iE2WNKSTqNtsr
IAZXfGFdEdNg46sNPkKJsWdGtWUyAe2gR66PtPLb76Q7DNt/wFKv+toA4LchNrfr
Nyx1hekdji05GZ3O5n50dJnjDUiRyU6RMQQlTn3btQ8SmxvTWn7LmErY8VK1J68R
FmUQwDQ5fsvn3rxEiNnPW4pOsjACaEEVHAxulpJqQBXI4d3Kktvza0Mz8ciLOGL/
5rXh4D/ypH8QkOi98X/YbOnT+r5HBPqtdZh2CqBZy55K0YU/dr/bnTj7tUHYKLvp
K4N975ALsivNBaMMRj/6kfXt9d3RBTfv02WVyhzJRf6JkMzDyoTxBBzlh64jb3Tc
KaRpn/+E9EoJTXbaJPldA4QLEYDhKd5g2KUIF0YzSpFHZe+we5L5iF4BwIDusaB9
nY9ppugjKIkW4jpKMO035JiwpVXB+wReIhv+GWSImUY5dKTEjycmhzhZrEmVnROt
5bE60TpKxLUNyqIILtk5lxCkNFqH166cPVZaGE/fdjy5bOtJCjjE66pUt0/xdpHt
PrsU+TF69/a8+4jIYv1sO38zPL2nt17t2C9A3ZGlJxwW3yf77n2cuz+5E2bfBgZe
Y41HOXlZncBc4FcgB4eRxEu67yzCiqcxR8oITLPTx6eZA8BrW1LGgW6jfUFv6Dfd
2mUY6S09w2yYt2ynB8pexvzOggVn5rjeaq1/V5xRyI21wmDVmDjbRCFVHlSPYI+E
2WAw1P+rW5PRwLOAYnvRzPRgcT6uTeLolqBsYP1nN8ioguna4KMTHRXPSRvLCsVZ
k6WZz0pDxn4oYVpV1A04Su68aqNhMj/plok5zHA1BeQ4EQfjhVZnOayrZxfZzD0V
b4vhoTDFiz7XmCrm/dujwqlRuCEA4vgwwnJBx//rB0lWB5fBxZvvhlMGdroPDI2i
JzXq6nlUCBZ5DiJ7LXBD1zVKsdnzVnNjV8sghho/lAKLwIK+t5BvBvzlG+A6z+9m
pt5N807AiBdimW2AxQImCZJm/N0fJJZduiOpf1rPqpgq8yxiPhIzOZfFRFiH3ap/
FK0my3PbYpykjurSRFSUNvO+2xniRFcci0glhbr9cqk9tI1BlFq2wqqO0C9U2F4O
TCp0DVsYQRD/UAhVAhUVMKTPB8DBH3SRkNunvDXaU8xME9w7HI1t13NVBRRqocvp
HsoLxyc6Q+kyVszyB1GKSb0syphyrHhW+91CP46o6JU6PJJk0LH4rvyuRpJ5hwvD
gDY9of6EsbzF+fhh0gY41cKYuC9LsYF6PoQ9xnbjrTK6hhosV2KWka+vQ3wJM0qm
BXI9WYnVqDujuBeDXUoAJ4fxYRQOey3OuWoQY/HKkufCKBE3AEc5VT1fPL0Ih0Qu
oNpaj6bNciEAHUJcWG0RvDxohtH7N0Eu65oT6Ynb6rDrnxMnOwEg5R+YeuDr425S
TGr0h2SRoRguQWiTbG2Sb7R8NJChUrD4N+bvW5fNWM7DhCZNGhdGCbTfRkdz4rWN
CPTGcW64fiTSN5RUL2p0QGJxyBicwhhU5lCb/zFdtkKIucWQDolvo1AJ75XaFFrJ
VMtBB73vpuKl7gOP+PWctXWDGf80KR7P2eIHMOIfEwaJNyvgRXvLCRMlDWMS/1xC
8FtbQ89gvatrD+0R+O1m5U/tfEluW2HnAu7M1ujor1llf72f1pR7oTvdtLm6+zY0
jggFiq3IBpl8GIGX1DP5Pigu34wqHDlpZZ0S/M4XYW9qtoZ6X6h7oCde4+iQNOcg
uG6Qq1zHDCAutwyTliBebPKf64nyaQit+RtndKn1Urs8mzvHv0fShVdfCzFtKnl2
5l/9b9nEDoITUNnbP90vE6QdNna18C0jJgLLyAm/QJntymlC6edfK1k0L3eSJtqK
L9cnT+ztlVV1IHufxNjw9dTxfiLpk+AqI9Y3tpIPFRl0Ke83vYmM4GU5laD7QCYg
+W2QLxIul9fS5BtlNDBrZZN+PYpPBptMUqU0G4+Yibhe5aMcLfYbfLgeY1zdFDiy
3eRHboW6OU/cZh4f0C1j2M3anFjgsyrQ50I/ffrfeUnFtgNYsFzEyH1kd+Xyz5/Q
kOOHmE8sPTAzRheFyw6/g778aj6wg3Me1uoEiZ4SE4fO29wOoBbBCZ/IeOCuj5Xs
H51hExOMvkRzxzmmLH/wAsIDw/i1tM/5OHh0hXEh2B9pr3a4Uvmmt1F+gZ35d59i
cbXup/xYpNGJLNVz3pkPnRGI6kzRE/puJpnjzRPY/u2zx1JmvhCNHXKWR1lenprG
yMJLzgN5Dhj+eoK9g1fBmF/WGF6Vt65STQpcAamTLmDR9eYzmoi0TdyzEh5+co2b
zP2XRAKqvybCz3/udnNDfICrgrpFCyBUe0DrD6K3Nlpbjd8k0QEv9ym0JeAnr6C9
DBrklSHvzbzyVwzTdlhSfA==
`protect END_PROTECTED
