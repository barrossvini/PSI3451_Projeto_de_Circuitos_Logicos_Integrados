`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UJvKljedil5uEfdiQAQbfG0RN7YvuZa4XenrbcfHBK1X75VuxB0UGYwixBvnFMoi
hmTmTkbsY0cIxmORoVjpf8wQvgsRO0ScM8fVV8tQRDT9SEwP/bg07H32Pl542bTG
VgifgdWoRRxFXlpSqtdBGY7u+wi3PEMVESBB7pLk34x8B7HMesx2dS9hbA56z1YU
g0w1GtacHhKqWGJX1Q+N7Q==
`protect END_PROTECTED
