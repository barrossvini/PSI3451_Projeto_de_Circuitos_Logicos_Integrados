`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L1mmPf8KJBqUVHsUOWYJzJgd46tESf7xlBuWlw1pkVmlT+Mx6qZv2CR9BuMj4gC+
tPaGSLsA40X6QthRn1WIV3eMNKO2W+HUQ8xBh1zCuXVycSMcN4Gz/80SQDpjJlOR
aEVrgaBEi8xITB1x/O8sifN/1MKY2RGd0OSTE2Cd/fYpZ83sIKLJO92O72OzxheV
09l8pZ1lbLFDJSAATMZgJTwgThoPzmwC62Ezy1mZpI2PkUL5j2SCC/90T3KVyKCo
t02aKaYvgv/R5V6qetokBXwHl9HWQDhgoUqopUeJ5VNxRWevxSsZZZNLuvrIvJAW
Thzk/MHkt/ppPD6/qc9G7nsgA6gBekzbpKfU9SaGljwqvhXfVFtajrTVOge7MvxK
MZiFmJO81VHw49j5mAMwZpWqOu+ZDqCCGcsVe0BMVgs79uDwN4BsgdAK0KsHHwzV
5MQslOxN2l8YUSP8gOD25AETNUDP/W5piUhqykqXku9HP6V84jJSG/YjCl3yg+Hj
93HXIWAiemW8aGs5GXDzskLayOnsHZiVLDKGycRUC3fjO3TPgprHTRUqIm8Dcwx5
RuJn0nvm8BWMorVzfjx73ZFCMIjGPjq4ccxNwsUFajXXCksYLP0OgoRCBhkx9wSu
BRYWL2mlqHhntHMyEarsGpHDIaoeiuufKSiOSBtxPIJ55yFXpMPhVUVGDHMX4vKZ
5AhV/m3GeI9sEbDRGFLXeFo8YUzIwYisGjjjml+Vb6eaWESW+8b5q4+dQ9bOMbt4
C3BXuEDy2l/056DQXr7WLEeyDKznEAhUEzUX1VTmKy+XcQKj6dliI8AXkaKJDwuM
qWhnXukjPjQvfMtFA74gvfrNia/Kz0E/yGtCc++ndHs3g9j3jjGxbWO9L36JLjSL
6RkSDqTvljjITF4Q0PHedFZ5wt/kg19TUv+3Wi8L9KTgm1ZAAFZJDEddyiG3TRZn
q6auccbk3jM9mGQzN0LXoLs3PYwrha68Na2l9fbf66F7Lc39mGYi++BianvlteMJ
iX4XIGrASeOmVOVhtt9U+s+55rr+iSgoMYn2/cytWS6CIQtZ6EDgD8V7U+Y6alHw
8Do3GQvAFx0pF/D/Li2aJ/eCiR9nY7ZdNWuVvimKjXqzKp6psTyOfjLyvAzi9bPE
WKS6cyCBwZiROF81Taxi8VdLGYyBKqoz0L0VAMOgDEvFDhlacoDhy4rjj8W39Gt9
W06hNf7p0vwd+2Sw2o/PYx5cBF49Ln/iZg7AAuwXzI+JS4PbS2j2gNlt8Xrw1yYr
DLqqN6SfvpOcty/JCpIhH+Rju3nCybHsackBmbCwesjLKL1SybwD+ZJJuMJ2dwTZ
N/hxSCd22e1cfquzGj0FdFUgPAc/xhr/5PaTdlK39rniHQwAlhZj0/ZfPmWlol6w
WHktsouyiopeWwqerSTIBOiDIltYusXnxbkZvn1JKS9+bJIFy+tgM1GgOBZXFuuv
`protect END_PROTECTED
