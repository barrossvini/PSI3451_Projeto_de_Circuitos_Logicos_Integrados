`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2/h8si8Ky9s4VOotNwTNBT9+VDb/ih+4flDevAPXpeZTt0DjiwUbghSCYxxjK5aA
rqiZlM6pgn0mWWC0WiIiEpYXXkJxQgKumTX8HCegLx9V1n5x35DTy/2ITgx8HrLi
pR5rm4oyTTVyFQOwulVYtCBvuIlLdjc45rPODdxE6AFIywfy8E9Oxtm+iE49ABb7
lMeIg9tkvEP6yNzM0XEw0v2AsyLRhj7Ga/IBPFtNQh1T5qWJOVCWXxL74izfj3oz
jZrv7WOW9lYF9CmOICEBV3hELebSglS7pKfdUWORmzoHPg0NSQjXxXQNMVbk6Vkw
Ka8A3h6Z40S4tUF0JoCLlQoVHSz0bPjaN1dgg5fhotqc2tSYppaWZp6+UXgLT7JV
Q2VydiZ3fLV6st33z2oPBsE14l5W1huIlotIxt0+dWJZBwXZ3QECflOJb0zjmgin
ynqYNSYDCvK2j79DYRzWGq3Ow4lsEaSvWL2PO40dmX+37nYRHRwa9Tcf9DqtQNCV
R+AE7YfA9KYAaHckVruKaLd2Oq3Oz9p9Gx69iu9dun/a5lSHen7wCP8KeBTlt+Gj
sJwCTBtWCL1WWQjnnI+zZHZqVpfDGldfT2BGlWEgeLkA1z+8uv9mAoEd/ULEt+Bo
txS3ui0O5sEzRjEAmkJVab+iUHXJ25tNCCAIeRDpBnNCdVd2J8gWLBcZjzXFQrCd
xo5wkYq5gEcj7VC56AYdYWGJ3RRPSQegCxKgkrbr7/sOsRau3HlAhviktebFhn7X
zd5EqHNiY/uPPJQLJDqRz5NR+8bzcSPodHjxfjcFSDelSLWYbUFKTwB5jVBKpUxp
ajIjIniZaE8JwB3BRi4vfOy+PaHI7RscynOXvfE3AP0gFGidd9OMp0HEbs82XV1G
`protect END_PROTECTED
