`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNJBxq7lMVMmaSFCdGMlBBoa7arwmHba0mBOHJweRkIKeZf6AAofWXhsQwPqKJX/
iPjOSuCgIfpdcXp/YFiEw58wSqu8nDzCgh/TQhRRWg73ZLkyvmn/CX3VNoXJfaOK
LHdnS9RO+2iYfQCzhXQM8senga7rtpe3WOKWxi/vcD1kv0duxQpEi40zAp/NrB9S
WalX4jpDF6x0RtkxidrQIlkcjBjpt97bSbdBrsGAqjDyhUjGKK98DIqP/TDILEF5
Vairm5tol9yydfOCpI73u+gCr2CMq+rOItgnqbkQxA2MEJjjErkSwIskleQpE935
/1SFD+QEG0AEzX7ynt7rVo5sg0ieMW5a6LP2mjnBWH3173TJrLGhaGJimoiPDuEG
TWfZh6FQnFYr1smjFvm4hQ==
`protect END_PROTECTED
