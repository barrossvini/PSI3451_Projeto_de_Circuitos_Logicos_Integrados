`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aei9AkEvlK2475Gqo7g4faQSlNk25dlZOa+t/RJQ7nRThGx70P9VC0Af7TxhxEGq
bVOaxxwffZcSOl+ndUhi3Ni9IJTkBi8EvEqhVz3gGl3OQqWetrYtQ4XbGePhCAJ3
pdheiqnQ7ka0ZVzXbBoA1Xav2X91bTpYaB/IArqehwQ/Cp5ZQ+UnwUgbuMT883hb
ETTs+djCAfSRDSCrg5039lORff0zMjvcNpjKXZkHPVUS8XmQJXV9p+0VEBFGBrCR
NWWG61afsgJb3N6Nw5uE2p3HetFwqXV98rtI027TFGZBkHVfUvKUXWS8RpOkdMX3
MsjOiHHXKcZhtGzOQEEykkB7xr3UnSRVJVzjzt7zlxJK2U5h4myrMUsf7ndg8Fbb
rmVtwKa8G0IGKEttIh9y3vggJq3PD1EVrvZAKvnL3u1z0EM4bkZ9euVhANnfbgmV
ooc+pfsXeVxqFsT4XDmkz5F8IhwxS/iR6v1ThpRy3dEemhhQidjgVGV7a7l0hePP
NT8jH+howqy5vRrGMNk/7vA/0ogirvI0UBYGwlhh+SrUlikpiu5ibu5V9XZWxTVa
3BxpXlvHuTJuzPZmDoNiy2f/CHAnpyi/2FNQsWS+j73pXqy82t/s/tiDDwmzpLGm
MLVulZqrzPX9/ZqMijlSMXdYYmDhns0285+sLSurcUszd8BcYt6NKkJ3fX+pP1B1
qyzap6vZR9Cy0XlTnsSlbGXH8i4+jw5zLsnjA4aIQAcE5faDXfXODJVfewGvQqKj
TfJ1WM+WVKjdQ/fp8Wfharx3aXs3SeEE/YFGS5Bs/RPq0IXBU0i5V8ZLtgc2NOYC
ZTFj8SMM/q8xccgU4WB77glDSzyhCjtD2D57PrNjuwHaKGClYS5AF3iAZdrUF06Q
y7+0VqLhKUv0gXpGkhl0mNzOWbWfA9m7kB7/GW5RxQs=
`protect END_PROTECTED
