`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cA4C0FLITnzBqxYDJC8MiiAGHWChu9i9B0DuUZW1YE3azFrJKp6DMILoJhg+D4Zj
s09/HJpWMPGiCba67KhdDxgzh3Sc8eJgqKz8URrb5JMl2NyezbTrV0oXzMKAX1o5
QvNimD5EZ6DWIPOlQu4lltyf1g24SJ8ZuL4ZIJY8zKiOYu1Am+xV/HmE+L9o10Xa
o8IgqugV60N+lOmNAx2gl5PxvxsI/EXTbIr2rvUZubs69fhfkrB5FggqPrOA3a4Y
JUSJapOsQpZlaDXs9Xg3iuo7O1iEkedDnECBY55MGMSX6OeGnyIGhz1X3/aHPi3K
asm779DH/84ZHe1a9RZyCuNqj8NOVsRwi4WqVXeVKr8MHi6jqOKiASPkc1uWos9c
ovvwGc8mKR22RwP1fubRcpxhiNiBUBg81uwHgWteCMUzSYQxp+0oC0sOM3telluh
OdxfK4okCM8MJ/V5spiqghX6UvubJsZsgJiDhodyHkH/6qU1S40c50QZT4S2thq9
svDS3RxBRO/VxHMgeKYiecJBbjog4w7W7klEUgQ1JBzhzmMGAeYncSBQeQr/raU+
uVpK8CCoh32I+FFRS+70LdIQPcr40zWLAViOPe2k5d+kUghPorVjdw1FEW+RH7TJ
r3vDsdB1UFJ2RafIkgIareNTfJbrASSRf1eleTe/gOlnp/kFOCgQ/6ENfHiUpoAW
tMizGI7fr10W9qrP764lnULKzo7X9a/Gkimb7jXNQkBbDZIV8zLJXDYCrbAvcxdq
+ZfjcaICgVhV54UM1OlKpGNYXf9Vb/fjNW41Ya8VN7fRxVMlcDNWdHk7aPB8FkGR
5zdXEucY2xco2KtSy/FMSa37JkegKQ6I3iEmVByEwToLvQUz85K8SMvneLkF+Bzw
5X3gV98BZQWQSjWF+jK41lzMuou5aw2s73rgGvutMgXWdvgkiAuLzFFtT033oyNg
yUyNqawUPuWehf9gv56qr48mUrFR2HX4sTAzUfb+D0z5tiF1ygmEDMQ1NTwmnoD5
eeYhLZeuPVdfeIAr7f9F2/QWjQte4q0NArwwQHn19X8+Eorjb9gt1lFL/liK2z1I
FiROG6vSWRFQlspOf/w0hdjTcBooAJb1cLNzHQ8zW4d8dpbwWnVCq1cPNtHH0bzB
fRfXizKAmXZXIUF4J8Bp4qclOXJEL4FlMfoTG4c9r36b8cS2pBnm20rHlSzLltWm
XJD6gdCgruiiPMRLX2qc9LnnEuQTpGfdMaBTKl6RPCYJ/mSYMjLEe+ywgMRYU4Zi
mwfh+3ri9VkWaEoxBQtiu0r5oMDiyvUyTeIYIq64Uar/zaFhNfd1+e7pa+6TeBv8
aU/PWFKIMqxGwkMmh7/8/l8XbWz6Dd2q0Aj3zDgBsa4My8YOJID7ym/2tQipisAb
qv5uDFUC+R2rZUAfZjn/JlopbMlWBYiOSSwkBrkbLBh6lYELObvlooW3Tr4CmfQO
vrZ1oA3seUDxIOxJjePe/Eq+MExIQEWUS9xuSRd/M5gEYG79p12DYts1a4ua4bGL
MyPye1h+WVwqkV6aiRX9TC5zq5/iXstpT9CTPbTDN856A7vqDPsPj4dt3vm3uP5Q
QePu/CfZcv60pTXDr2lZPbW/9qnO7FEphOeAhU7Z59B7PGPX9H79lEFpPawOJxVF
ASBl1eZ34lP7Ey/BWzIdiR4GVxlZrmMkr7zABeKRbE6e/4egnQdZRcx+3iCs+7Fu
Hm4H/MJ2IlNy0SBV3XZEVOVkL/i5zNKCRotrn7GwIElLn6NOKgIo84MrwIS2hoUB
`protect END_PROTECTED
