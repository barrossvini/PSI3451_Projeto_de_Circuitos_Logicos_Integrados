`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ifwz+/vI9i6XC+VU4B2NB9wLDYT1g9cesRQ8rasjJPXdYbUYKLhok2sGgIQilkLB
ZPq9DeuoMRbObKLTA3oEhJ5w+9i8Oy1cu9F7Cm3OcX2H8fK4JpsIk6cyl3j6R6Iy
gI19voInr2Y5qvUDVcec6LSKUXX/mGgtBwzQTTlA0qdqpR2qnxWxOSEZgUKCFgul
F1BVo+ZPiOpdTGVSA82aAkd30ria5NG+tNbEUlZTZ0B5HEQ4ortTnuqrzWntzV0/
7UnbrrblSxAu9WLe1BQ8S0v25NzUqdKWs5Zn+SUjmmiJ6XmHJtDs6ar3ZDGz6B3g
eSUMLQ3gbeYqR4RKv8rChPMM2GJ0HRJwFUisEANLptjQCZAHVzLsCZUOzWK1Vesz
K25xsFhJvXZ5B+Y/X+GvKsJsbV2NpwX1DXZl4cJymIOjkFLefqMh1NuNYclEfA1L
ckReGOCtg/Owcrf4J+nUfxwMiXRfyfOQAQxfzsNiTERFGfuhhpgGpn1wfSCN0Xmt
LKkK+eMu5GGFe94jhcNyvAy4qMRvT3XJA1yn2KKAhnKRgWggwtK57BazjnT+YcwT
eEQEPYuHV3hbomxw/kdr244+u8ta6AdGCty7gIOXGcpSiok3QqSeOWn8k7ez1lUc
8pn5wl25ZEeJeMAa/99pohQc1XuXHrYVuSlT55D3m76sk71N8pDFLsK/5jqCJZqs
lXevwl1BRTFP7gMyX1W8ni69C25VWZOsm7lUThb6ay/VDaA+vubwM7s7YykV8jo0
/NCrv19vkGyOP8D1CRmiqlZcf78HOKqbTS1SoF1Ll7v/A4GnJ/56pHs7qzrAUzFI
WuYql5pvSGAMaZ2OZcsPeYTfBjT8E/EgTkXQHvL4Gfxb/t90cs05Q6ecZmm1txXm
hFXqngUi7oXVD2msgaUzy5uFA1MSftdqwwMosEK9lGfwkGsRbA+nomYVl+OR9fgI
aHGeiUOSxHorrWVOIoYrjKtAGsYSxvQYVyJEpBy6qERCXnrz3FzFYcEn6wMEPMTE
WDZQpRafZnSJBaM2sGRKYfMgApugLLGAPPuBpmaeSuzcnnWA2EbXKk6zUOv+fZky
s3V2Mhoa4zUG5uFSn+/puqp2FeBYbOXCsTLd0xLHNIC59621sOXZNpIGxz6Y5VzT
dOak7eigU0IlDZYhGmQeV68VssNcLif5Hioab7QmKwgdoT1VwJV913ND8lcmuob4
SKUjjtJ7esSowyZ9362o/sTLTcFd2uBL4UbDnl9GoiPhLQLswoKQmUSTiTV9JKu6
xQI3APhsIryWa7X9X2i2AL6hqBeePrs6S/AsK1XmypLnKmlRHi+R7/+3B47nIM2r
hzpzotl573Ri9O+qfMbNPKJiF+gEbEsQllf01dWaBZKONAP1IFKn3CDVK08XTYBB
DIzg23enW+Gs2SgEPiEj8xR2y6TGM1cpTEgxhG+zXdvNRzPdbUhznUY7OFwa+Xt3
x+NdhFyRzoVXaHOi6HUcBQ2yQuxGQGy6reWza/Sdk4p0z6Dp6V8FQgD4DZM/UW05
t4sW5bYWIipl522skhc0Mb3NES9YrvJRNrAhX6CTQyKTBKxIzXxSbUQRSV77cK/a
UyzoSqGidHMxJfDPWaqUadA83KvrcqlZbkYp72i+0JKOtoKnSC5ADXg3shODb2ZG
hXCEVA/knUNKaPhEC3LOR+5oVo03TuGGHibOhlIVXag38PB9QBjJWMNy2J+iDpx9
4tAgficunkhnMkfp1RCgXYU22w8kbLQSTWyxXbBdOM51YFJ1zE8KPAiA3GuWgJ70
gyCmEYlXay+g9rHC4jWa5G57WTV0NsWzD40d5gH23GkrViGCtziB1WQEi59iFJnD
h+/ObU8iEIFZzIDRJB08AQbNQfDmh0JzfyG6Okntf9bRMIFqU43/J/tNibgeSUeP
yNbuBG5eHFg/MSedt/40JsEmyABdR84fEyN6pCW96tozJAIk/fHfG2L8RBw6Jxsh
ZqZlj0LgtDBXwexNjs0jWLD5J9at86oh4s+osUU1ub0HeSHbTE6YAzHFtvjB092B
VndAv3zOf20Rm19KBkNTZnTUGXicF7DHny9XsQf0PwzH9h0z4Z3/de6h5KBhQnY9
Mb0nq82md+WdXn1o9i9RE4ZeeeN0gpR383TP1xFnu9AcIXqPmDSnAlPR357VHzJQ
zBykZ9Kv3B3syqcvGqNBYdnVIRWy4syBvREJ+wup3FaMfJTGW0igF/elISWl5tVq
B+mbk/2h2E8OMP1Q0u/k0mwfyNu8GxtwzFEzzvs9QFZtPjxrCK/lQyJdH3LULC/+
9Yht27vvYapTtNniqrGZwWOWDOWcWfxbnKstLdXLN+XKJmZ8X89DhN4f/TKFnKNF
3VJ2X4GAiKFp04/lLiEGA1s7lGYvLwxz0pYHfD+L6xANoSCglrUMDe9Sb3Gx4/1o
JtVq5q3WMINr9XLlsfpDX7yVg4LrqmWQX1mIaq+V6DljabdcZiZdItKfYiWqKgES
2nuJtoiCPJYiFX++4jQC82/QRQqBK84NKzyNl29EWH/9cEkVjY1tJ02CY4nWFan/
9NOTwIQDFjCuZRIALco8vpqlOBHdZU1ZFXlA1PMuTcQXjrZ0J8c8ghi4KxinqhnK
P5dW5SDKbZDWJTT5sEYgsi1Z0TkHZwkX3150XFI8jcENxTQzpGVi4snYDcLMrTrS
4jtAzj1ZVLxToxXTdwHfWQ2ulKOhQr9lJeXTD35aE22njbgA/+5JEgZpP7KICSvY
kKZQNLHOIqvpPN+/x3HFi4kz2hKRAR07HH0NFemeSzBexs5QxWw/GgRZzzP1wYHb
u3y0CN76CktI+4o0n14zC5SmdJW1qjJ/5KJhpRUrXf6M6sXjYRmLjWL+8sVDulmC
izcRCASh/dl5AkR5WbRf2D+Azp9Gt5Veb1JZKdQAAxbkf3yENi2uMKayIFP3F3/3
6FYT7lwRJq+fd2OUIOj3Wp7ZziNenTicNlbDifLro6kZjc5M41TjzUPbbhce4EQa
n2/NkG+j84KF3Uvv4p6qM7roqhgts7HjR4E9iLw6lak8tsPOgSeyLmoNeg1QQO0J
+cKqmeLhRKMkeE1DZ8NqQqf/d+xfAgDAqMfqBfc0QKH9sNZWEimVa7ejmQRTEFPK
XKw1BcouE6RuhlbgsYGC8COGNWmR/duHV4c3ko97y4bUyjhBB7rr0b2AzxMcVkf7
eGFzTxaNbDSEwne+X2oCrbbsvdez8c0roGtPuwSUiBUibBU8uAqVUFrvjvKqz1qF
icQxIbeZR2QiRLAmQoOGvq2nELfnNamvFAdTUGfdfGU1isVzMis1xq80WdfKnb4G
S3UkdjQHPi7hRugms03jpIWNn/pk3TJP6bzziqlYknZv1pAmJn/vWeO/t7Q0fuF4
5ny3qmE9QJpyQ4reCnuErEOhh0QQF7YtMvj0jCKW6Gy3Zpih27aqA9gv0IZgCYs2
wD7Fi6oSew9Gs8XfHWLf5st22fxlPp/rHWu87bLz9v1j8yV6OcGFdl4uYmJ0KrlR
jh7gIxJkDNpIJnq63YE+pqOwxLOqcJMSOp1vJHnKx7MvrIWlqpetVzbaeqwRZWy1
46lcmsPETPDVa1/rO7eShv3A8jKAhXwYY5lGeDfH9sYB9E70QVOPFAPu/umrrCu1
OdjC84O2/Dp63PYuuFgA3hx88FsF8NKE1FpeY+M3kPdwx4ebjjeOOgDP+5Ov1rZ6
BziFEHtsbbt96OqnLXzIRiZDeB3R9D1E8+b+R9PP8tDSplarTU0upDvI7JBfM1Nb
WEap+lMTq8bl0jYPb991hX6nn6S5vgFTzbnHpF/0L12ZX1Q5iWBPHbQmiuUydFN0
583Zbtw5GsgoGJUmf7AVRJTp/ExTjb6XhwhLNpH9ee/MlcCRnGQB9Xxggl3oGSR3
dfJF68TvTzMXB+79iq0IwwdoFAbajWozXhdW77NIl428guozmcHuFh/uRgW3ZRZm
SXaItUj8CS6Wo/CbbisVG/KCu82pbS/RyrK9Cu0KSxgaUyQMeEjGuy3InXON1B8c
aaKEs7Om20JD1aY/Duyx7hy8RKBd/50NkZOIqoRB3AohUI5oCsitt3nrIjr2mfvo
/tn07EqSirZ0FqhHbxH73TxeUhmn3rZ0ebKY/rbfYGOQ5KZD/Pl6q89jCMBfTtsE
6ZnXypjiXlo5jZpwdLgrlsHxnjF+UnHmDYGVhAX1B5bERuFudu/9YYb4MKbroQQT
dhnr9sDa4qzUjcld6CQC8QsRoYWKemlO2bkUPoNqMWepKMMP7gmcgHAh0y7IJDj+
bx8VXO0pSbMXS+fIFkogVvbpBKM5rYM/XD85tApQO56wyfd6zeuF0WzpNW9Z7awC
zmqnzaOc8y0T6jel+KSnq+cIGnxgubrLojFonTDWjiZWWwZMW+nHsaTyUZ/tMKry
FY4Mdsi8vn/v/kKpWC6/uZBvn+sveURR/T0vYGPhkq2S0VTRIYHaVhQb47vWoBeS
l1SXYX3p1jvhI07ZjDjU6/GBGaevoX3ey8G+0YWp0VRIxunfvQqMAnqVxl88j79a
EH5hjItehNbLY4niJgcQdCWR2wdqTdtLvjtib61VUSbas0D4JIOGLxNIquGH8Bz2
aJ4ZKbXrVkB50AHyEFYtMAxwcdx0D6UfnxRBNLynklNHhX50lxHVg6OwlHGLGFyG
cjT/NVC2hsn9pmnbwv6RayuRCSJe31pHqJRp9gaAWM+3uiQMvl1KwEp3ajHCvw4x
K7sb25BM27Pb9x7iVUSA5QU2UVn1VBCeGngvNLQecBtdwixsG/h2QsV7FllzG4LX
pm4UWT2mi5Wof0Z9JT1BIHFi0VlXcy/y8VqiDzIlJP7/9sYiFCKCsbK7E56poZpb
uoDhePUkJcf9a7f5IWJvZqRIrrYEznnbQUBlwsCVlojAMezOsWhgJqwtC6+XEYTD
+KaQEMt+FbUqh8L4RVpWV5cGji9/cZxgAefhWLK+451I39DOsuy+LpOqMcPNRwKK
x3KYeMeiPjLEScfU0NVivv+vfAXAcLH/7sVL5P+wf0Hmw2Q8twp2TKjfxYFipYuL
mNFKoLEJJ/lVSxlP14ZrVP8xUDWwCiTo9EMNuGvCm/+2dB80EXplSeLyUshRGNLo
GufmDNqTmMoAccNWneELuwUC/PaqAddVz8bNggGlZse/jdXsCtwjDgbx+pwcz6bu
QvranWi1dtielWY+7atQCDD5Qi3Dn7S6x5yaxNHeOVsKZaOGPmTporS6u2Y7CN5r
vBssUYU+mjB2aLLGou3QFs+WuR2TgYG1QjcpkjkwjmZ3I5MAbj2mJBDPiQOxu1Y4
cz/sIuwsg7/Y/8/aftkU2mjQV7nPj9pAnKEs4Rkcf1JUTq1fWdwNxgHL6LLoIvi1
2CKT1pawYgTJjurEyV0+g8wdFX0ew2doxDcIDPLd1wy7v4KZkc5iUFG/ExkfeNkL
RJ5OM1tA14SyY4gFV6j2BgQMMr2fs+NN8etAiTTxueV5RGxbmSDv6JY3GRPJqPQc
1nIQPF5jehWu/apNJiCjBhNTPL+YfS5ZTsbXdt3yxbU3RQgJiyap5ifT/YIOD74G
zrNaqwL1QE96Ghb4wh8zILBiJq1pTI8aXzjCyJgWwy8b/2x/uQVRNMtsG1NzG7ay
nLJ+TkJhTnfsutAQpIO2dnhvGe/xgzGpwRZ45ml8jg9E70co9ZEYuBMPVLjUQI9J
ZWoxlCuDJt08K+LwEI79mIxf83hX6jpKoF8JGZi3hDz9wqIF0Np7LFFI3BdOpaWQ
PK7xCQtkuR58F0IqopyU944NrL1OoH2D4IVIhOQMqDdmGeTNVM5Jqr8f3kJMtoeY
1IRLnDyx27VG+TZcAaDJYKEp4qHE+We0aaK+YTvm9RrEWoWK/rtZn/Or1oQRaakD
qCC25V+xNmNLqkiomunmlT/wOF6ybIviMlZGKaM9CQWRrHxLajm9Mk+xc0F0WffS
w6R9wDIMIV5f4QwsCdKDc+GUcqpjMt3DOl1qmxKxzA8IGvDiLuCwZ1qQ0yaGW9m8
7YDbQNfnJu48olx6S7DwkO2+XzJHIfcVz2UHqIBgAJv7NC6eG/hTUAmCsszf+8Qa
FtxBS9MpYdMWNiuSacUsul91uA3+H3LxbsguKGs845Fg+x8H+uJP30j+9lGNKBT3
q2cPDFKuef643f6c8ICDkKuHblPRQlIo9lN9QqwYC2At9sX26rZ5up4WsdXRw+Hd
dBgNv7jpaOCx+bcFJTjhHIHMTZasxg0+/k42eFcz8+hgkoN1p7b5fjZ3akEMFimK
IySe7qYrvRGuRTuuW64qq+QMQGjX8vVaGQ2M+ceGUbT97VzApeUo1+rEhB2zHFS+
rbbrCxiXvxEz/V8MvgjdYeo1f0B2H0+Xmvee7wIoyn3uQT0UHz/B3Pqw0g/UcLZx
COGlwHsz+9jrs1AyvnK2RpMjRF0IEL7/gd1eAe25GeeaF+mt7ckF1BSiBzrvb3xa
q7Nxf9JGCGR8bLPCPxwAhk/upCev151uilI0yv4nMcxIxdERbpgxHgBvFCvxufeh
HME0/QquPdnIBFrWqCRrArY5sH10iOEvavGTxy6lNle2mNoAKvgjbrP5cTv7yR0U
TEeGlXjpkcrid9MyKRzs39Pvv5LIsBq7ordVCGMlQNPkNI4lVdxpZHoIfHfJUvhb
z9QChuA05XJviwDsL3ACAHeE2uPwYiR7JmAr04LZW8UWIEAg7QdQEuRH+CsvCct8
rxJOHNyPqNzWxZDbq9y0XlxuDEFuTn8lfmfBIIrH/dWOg4RgnZ6x47U1c5OGcyie
yfHMxKvY6wy9e56/0saAuAO/neXfY/o3NsvIA96s5266qtH1Fq+yLnjzBsbdrzcL
ZLTOXuhhfE2rx0hATS3YFuTV84LgJyIQfNAaJmGGjGq0Q+WzD08O3WnpVfaS3HMH
pnCBfHAVk2T5GRMmbihy6qDS+ujvq+a3g3x+vq1ZXYoNk7WStA8Rd0PmdzGtig98
z5ldCnFCGFxd3RiZ140ojtXpygj3+TGXSNONClShWJm79/XXe8NPYsKT8aMpCxWt
D88jCMw7evPpIbE5DAcQMsyCnyCWBUi830y9egqbJVW0+CERWqREgRR0g/bow3UT
juhil3fhgDgI86JwqZyVik48h7+5blMzu660a3OjRQLiZQnxLL6HACvJ3pLab4Sh
6jzHq5frF4lzDmYf92luvUcy+QGWCIpHNDeKol22n9M4RjQNQpmQZJB834LUoAeM
3mAqh6NqvfQLHb2Iy/gouwYTBjUgYd6UkRZrV3cli12saCt1f2z+bnL3hxGDoMRW
xNVnFn0zsAvdNayi0MxBy3LqNmpIUfX0bbolcRPLfq8mD7LytmRED442wiP5X4+v
7t8CTB4mxlJConqNzAzgb516qhplACFUeOPTOxJAt28+8xQ/BbNfi/9BhSv97xlC
DemNb4XIWPZ8lsyHPkjSNCph3NQtS/VyWgKcjk7dQO3v2o+U4UUJ2qhccP0r6uin
GLIFfAzGmxuHspJdWZ0+vRVR9Qc9qT5VWxzdImR+qPg7uR5Z+g++ay7S0qv5q8VZ
x6kJDcg4zve5b7qLq2kGchqOEyr5HN//6Mya5GPq0f1VHHqF2wXNuX30JywD4fDQ
doSTPNrRwVOjCZ5RGJD/xsDXYygcuaqePgLgVRhpEwv4fc3IjqitN/Evj/WIAcmC
Ra4GuUV9nmDBWBR0nwRQlVlTLNlKnNMwx87uxiPTzKKEj1SV2WLdZYuWV4A+52+j
vSeMh69DK/hCF6hpVLOi5e2U6RG92ZvGeX+XumjWXMmqbwJ/L4fzHvqYc8DiaFtE
of9XpdJIKkJNzaLUX+cuBwrahze3M2I8dI1jpwNEi38wD9ApzRGyyAHssdBNpp/M
gpWbT5osbUHrxSQOlsEOAfG9ccjydThEOdEgxO2uVMeOtmQbVTQ+ZHaIplxGFa+L
0oscJ+TxlSVu8TDW1bhr8nqeWJt1a/5sv3/yb9n1YItAGwAkzu5y4ifskAtj8gTG
BZuze0thNpwloEgfWr0qlOMYMzK0F/px3oN75aXnBarsHcRHxMJzxguRsERqGggh
a9+UJeKoUZgnOSu4//LH6YJupTQM/cOqrs6kVNn16UdF+GEEqGMAku2ZWE8tlXXC
5FqdgMW/Si1hHL7UsfP2Vz1jJec3jEzHXMKb0ueRl+CLovGcjgeznztJO+7Xo6+A
KJNodfxNbGQgWKVrCLNM2eElv1kzdmlrtucr/pYOy2fWbUaEMDsHYmwvV6KzA0zS
Cdgsaz0mqqE0vczDf4vQI04ZTp7rnuEIys68Ynx10/oNdrDZeQ5931o1l+VLJSaB
bO3jWW0UuEBPz1nGLC+83vGaiLQTvR0iuzbYuyYNKpu3VmbRFfx5VijFTpHwO5ds
dF4o6yitSxaZUq2zaka4iabNNbZjztGo+Tefev7xvvo6GzAZ9srBe043dQmr0Bll
cptftFhynUeikKZofoRekxZkSmGpynK2SDPiujpIAzWKFCF/7dRDwXjaj3SVXQbP
nIRqtYZDTloWlZIqyBtlXAUFoBZE41LdWD7E+0tMA29qlEfvadQYhRhARkdP5vuP
2rsY6JafrZAcfOUwdkG3gOwrjN73WlolfZCvEV1aZRr4pafsARf3FYRWyKlG+zJw
BRW9DxfH7LecDVQ/YtxN3WnuuxyB3fxQHEbtLzXjRHI3ai3ig/UBsLGAeZR9OhZF
IYL9pFbnV7bUzPPQIWC2vNUDP0QaRfJKMFEvlp5/C+H7KP2MNwJHZ1WeSX29YbI3
MaxHkpn0dng4kNRQiV7IXb6YPxuKiEcDLFRu80oGqLU54ee3yUN/h0mI6H7PQQi6
14SJg8UplZxP5D9sMyWCWsZr8N3ePOUjUAxD0hoH5ih98qssRhzst7cXFvYZ26iC
Uyk7dbmdLxzTlkB5sJzOPcg7mOtEh+yNoR9fXLbXlJQtLKS4Caq4bn2HmhhitIpT
9flxH+dm5ClY+4Ptk6mIfpmpMM1KEHakm+MLb2jQhCrB386/78vf1AJZtzwJmSkI
oqBl8iBRWhV6x+y/e29ZYwldB8TZ8vtKltRDrmFLIAG2xXI5LPNB0o52UPkhgbXl
g/nJ8BE4FcyeJ1V3LzreeJG90qqJmzRqfNKT3rDDfHR18fdr9Oq7E6HVRVjNLRC1
OM18n4vi7YPrrTBZVCzUSnnyUz74FsJ1CJp6lfsol+88XyuNdP0uOpzD9aDIH6L8
EHoGiyK8ypM8GJKMoDy+Z1O7cNv/8owjVUG66fCjn1RGAtLjo8fuuG/sg6HQm4Nk
yPnHgCkP+XEcYNP71sJYg7LjyrmcPBT3WDJdWbdeD8MMfe6g/fKRx7D36P/YDkrd
CS1y+7VybriEFFsA4Zb8uMPMb8/7G/0RGNvbPUxFi7OlTgqkWTPfPv9BpWoWoVkM
1xxmsgCF5SC7qR/Ey86ugKw8Mkj8eqCyJal25Pvr3ijj8EDz/FXzdoFLYyAWEzw5
c24wyeAe1MferId0ddDehVU9ViJHNokcACjAfYgOe0MLbNklSlVsptip7gxT6jCY
e3Z3VEhUjece6XwvZXcHHOFsuuOLf4a1qqB8ptCq53GYRDm8UQJZOIujys1q+gbQ
hK9sfL1Pf5+ICbOqEXE9zVQD40nkiZb33WEJmbxa7Lzg9+KhXoeOURKHdYbLueNQ
4Csprrc6LgZMJxsc8ECKfAnzCNnDV3gNjFh8cSu0cE/Wi2tcuAd7lLgN+Gzpujrx
4uykf3/O8E44krgNaOGffWKC9zhbmzRGpHTAs3RqyAMmO+qfztEyze89qIY4yLGC
DjZHL2zGIMB4lDfcyR+nGw4n9daL8ysLQpZIlorfOYIKCWkw4ukxy4sazGyA4Rjc
R3iarS7CuB7XlVF2/JqNUAU4ngvwghb85L0zWBOHh3T2CFEskWs9htBIlBxsMfOY
fU2yOHD2X6MkSB4QxZ654Y/wvJ46GhowfSgXqkimkqBhvZGS6dH//gFLnM/4kSdN
SKjWXIhyf21GTOXZ1+4dW7g5KJeftSfHkt1AwsMMgHNzGKyC+2KI009E9R/ppVq2
q0YgywrqyTg2zgEPFBgIXA/w4sLI/b/dxecNhW5lcAyNKYJewwigXfnZ4xQDNYic
1EC4V+lKkIo6vFCtEYD1GBWHhQf3qA1AY9H4qIWBsG8EdcIGKUS0vPVecRU/9bhf
rchIbbY6VCGAKTz6ANCNivrUvvtP/iAfDzXWNDvWUU2RLu1ENg6qQiQ627e/849K
350/Ay/aufCvLlrHNASnacH2TU026/CtXNt8+MmnkyZjuO6TcX7NoYE7yRSX8BeC
jTFZxMofWHo4CutUccIY9UEFqc1TVee8CYoI3lfKINgbjecAm0edxqKVTHodfKLV
zOrDDcSUqQid5vQhfdeUjgd7eKxl286K5Jlv3R+rSN9TnK4xp2HWfGT3Ev4iayuB
kcrKU7uWL50hIDwL59OsQdiit56VdfkPsPjfklJ1KUID0WRYbmsRCK9Cyu518UpP
Tq3rv7L16VVafFMSYaZGt4s9bdgDyEG7N6tGlXN2s2ztWr75DQMw92466Yn9Rvbn
GKrXwRKRrCubv119mUi1qpRurgktd1/eeccj9q2hfXTVJQ2dV62ZWRn9dBTh300v
ZXFPvhBZ9f5pIQZ4lcqly9THWoqKSQskrVrd84bvW0MJe45ci3eG0oDqglFVhtCw
P+BHJDaO8LP1tyKqrAF28AhmGPr2D34N8WXL/nnpz7Gwq4aMcWw6nzjk6JPZfaJk
0rNymOMwBZ6BXS0P9rvx22dhkKK4Mj7B4HbkyQssvyIfoWyQj5OVzSxQNy2SEZCL
JPt2BAM2Sy+5E11gAfzA0+lyfgXlNRT3Sm15Uad7vEk=
`protect END_PROTECTED
