`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LEKBL8wREDPmhLvk9pbnc5hcEU0HTcEaRBndkxBU9Tpill8n/FfED3McN7IVBuWm
V7NbZpDH2r401Mr0SEe/td+1LtefythS+FPT5cx8RJIg2bvYbq7+u/qY0Tz7GTbd
7OXIG48byQ6cz1aH5WqSxzXzEQdcH9i4xBYcIA9b7TJrMTO7SEQfWSjSgGTOX0jY
MXCz3DyBnE6fXp495hetaNt/5U7u5nBFVE+TRc6/ASYe6irGAUhNvFZQ5SEs2Up2
SrQ26lPWX4d+wyw0RsWbXWO1BAfMpGEOF2BZSG147wc2qsj3pdYizAalhTMSlnAl
HP9lYBS7bWdUHgcvJXV5PXOWBf7r+B/A0QrKzwKOezSQiFk/s58WJ8LMvT9QFbMr
rgYlxdHp3XYE/LdN5Aq35sE42HoKSxdGEcc4LZe/h8pJ4sa79TcmE5nSDEJaxHSX
xS6PqNKwlh3YkfHxZkvSMO/asGC21sEw/KyvDKVdHM+T/fziVYWa0JdSiWNnIgeo
RwKuzuhvAQ554ax+yvvOt6fODUUO0eAhJ6HJiF8itWWkZzSgVuSgB302XW0q1Qp4
0i/Dv8YBTk5hYhHpTWX6yaZuZANr7GoX7EVQ7T2PARVGQVc3OUlYMREnhZlFAdTK
BgROhHGgXnDAOk/+1gAfBCUCGMA5/SekxZ3bf1ag9ktEQW9nlkPnJQfIAuVXnEBZ
wXytxDjaBSDIj1H6Q58yo1kTuy84aCcOLL4CCIV1BUwTaMDXd6t3tspkUfNFmdlx
tTmuTyz26KtzplEcd9K4qmgC67a7p5tYP/VVj47RK7EF7KOYmr4hjV9shZuvp5E6
bZ0iSC3KpPvQoXaHT/f9ITZH0jSgpWOH9CzuNCz/wyqlVsIrNfFRy//c4ujDWyaQ
l2nG+EzkJCw9QTq6BhlV9K9cgReolYMpHk9SVc2fouHhUwUsIBEA+pULZn4E6VVF
cwZWTzELtLtGXzrAXW35oFXNviWYXsoMNPY2cwQhHl5KSIsFmAriAc284vk4/rE3
V8PC2aUj6/wUzuVhw0U0Le3Kmk84uBnZNidW8QkcZYmHebvgZjZu+pTX/uwXrJEq
0ZVABZcA1VjlygOP7DI0n5mngX0PSqdpAoBnO2y3//kO5qH3T2frD2oSNsk9qI1b
WpbAv4RlBlLAwP9ujJqlaST705IqwMGjat1tgO291YbuzP9yLuZ6jybVt5ej3LXW
qy14uY6drzDw6kggwhCjTIaOGUlC2sEiUnICshmEr1eDPTm4qbsq8Rw6y02ROkSe
pnUhgSLdCV70+D0g21rXLVO13rZtXodInqUkgB85i29veE6Y6LMJazGBrcr9NOhh
4k24YD3WPYgBgFSzevmcy95aqDMlyTKllYRgXQhimRlCCyW3WuV1dgoEwB+HQcAL
Sl3WDMdCqZescCYbIj4k7Y56BtksGdWGON/Or+wGfSDJObiaEpmQbaVDWkjdhSs/
RGq+csEQDV56UKRO0vqVINRdU2P7ej6Z2Xb0pJNel5GgZSLf0dfnH9Bx+um994Ym
EQN+ZTPQgKf32xH6h/82L7ELqx+7eNjv6s1alJ75npZ8yPcLWr4Po7weOVwq9nTM
DOvCkByO9z6puYkHNjWoWiRLEkvEujt9xeyDd9tCwc8Lv+EE0QpqzzXQL7RD1M8c
mCRITisAw9v6I4duaCx4H18htqrh8IBtMIhZeJamp7/z2Ek2ovOUFcD3I3YIZoNl
cztJ/tdArUWbeh7rnwxg2Vg3DmhyOq2YqkVaqaoYxahIGCJ5430NIV9D7IpDipYm
L07Kq2zuoRTYIScTDD67MdnZMu0x8IFfTEY6dyb0CTLdnh+uV9hbImouFtWFNBVA
ewC/17Gk/ZL3VTlxUlCCMKOncBrldysXJG5jGVWWF8kf87b9Ovd0eEeIAjBuKMJn
RYi2Hpc19WV5PU9rwgW6cwh49Tjd7C+4AdKvT5N87R5V1aN8FBYsLCGYgX/JrZIi
VK1p2BTw4gQRZ67P9RRE5LDMwyFxP3om8R9jJLU1umNv/klHgvkDc0IjnA7PrQwi
lgfrP5zSHcrt7fpXcQwBWmzYyASnvI/1LRuqThleudZexMzoMMfWc5Srs1Dn+29j
oN4w3741fIvjcSAG3ydT6SjMmX3EiWV3KtsEPjj+jriKcXBiCgD73MQ0Z/DP+XMM
ytmNlR8MfdHwLE+wWWsd92VlJrS+QnhZd4epTF85CjqFNC37cGRJjI2McDVYNtoN
FrA/aD/mLgROw8TbHx/rqPgcdZWEGYq+YKIAbZrFZ+hV9AbiuypWADj1NZpirfLs
HVVib5eQx4X9wiP8DNS+a9JDDxK8GwOgpVB4GLdFYlNYh8vLuZ4AMDK7zKgx277u
fcWGtRrv1190TPtPvNNIo0AW/onY98uoaa5JqWMrdf4P+57yWp1xxp/vT8qzbl/s
dhsuTxMk2fFa3qJ736PMnpa23hT5aKOWadYfT0mZ1ts67kIrVcxlXbqeE6FOJ0re
bU/EhOLBjNNRQcSAH3CO0Q+HbJS240CW0Fj37S+IRlvCfPeHlzk8vUNehrsd/XJJ
H9LcnglZRK88mI6YscRV869jEz8++kGkONHXINLp4XRWTe4sEdLHSQ1s23ClAEpN
ipGF8CBO1lb6zRzKMM8ydqp8Y5HnLCKM8IKHTxJo0i0CWeon8wWQykT0s/G++oQf
YGjClgL7MGMuYxcl1joHvoYGVydp9cj3hf7U8DAn75Z1uG8GVG90E2hNiVKbgUJY
i5K/hS9svyrdOsPWOr9lpwwfgn2C69R8NxfsD2haOZYvtcTE4A1hDlWlYILqW+Yz
/MKEk0otkZXUwnPQqIJjnWMAydcVF3bcJHua8h5v6eNS7xgE4lHNpNp5c9QKDv1s
OGxiNmUZNLWtp71ABh8lFRb8pHp5HCf30/UPEgZYfto7ts+aDpmOI1o/ReJipp7Q
qNlnqwBos98b/aFpKc7e8/l42tuf2a8cSuAQZb8B/cQ6cu0Uf+d4gz37eG1UlExF
zY7nNiD78gHb4tcbCAkioplYanvDfWoY7hj08PGn3NDb5PGltxT3O/87uHYqlfpQ
Dw8oQh8fpmnpdCrT7bz/1EPmORp5hha7W1IUAsRepzp74uOBfjBHrq7PZ/LuZAqk
fmTRsX07m8YcJLCY+gLHp0FHh5EdUMZTpI8W3wmUKc3E+8awHnwpKFrC2TQO4R5R
MuzXwgb3PSdj3QAMs6zODml/C1zxAKp/pIi60ZjvAJ84aQlkgfZ4DlecEwHfKhuG
rvRlrP3I2YXkB2oNvST1frlaH1cl+JvnWKR3H10E3HoFzPSjBev2PZicKSlERRqx
kWerfWXaaAi10yPjBug5izy1eR93nRRs/HbkEkxaxNjoJV/ZGRB2Gh/t8uidxqst
KnrLOGfBaIlyUbqITiiK9dgmJb0HTiW1KhX51tGBBaTX85UiiwYld5r9O9F9NwTP
bxwYB07EmMp6R3zDexJ4oYrrInqY86Lc6nIweeQNbM3bpRjCbKkCLRq6dCXthjXk
b7qPI0+YWvfjM0aZKLcinlEyVYassrd5wCryDhe5MOukUEju0EClNg4Nl7feML5e
KaWxOAqGeGfzAHOQXe81MwDO+XGLtoQ0Hyxyk4luCKN4tycXDTTsIk7qxgrJqd4B
TKARSRebZneAL1dtDWfASah88hgSSOqfLQi8oPOS3qUd1CjbX0eE1p/gjfu98pf2
fRKyOlSHXGbBvReE+jZORyfGUfrNprZ9fY4USRT5lniEr4U1SRyMD/x1l7CbncHK
V5ziy0hYZFh2STJkQ20aWGmPYN1JaBy42vBgiXE/5LV5YCEZ+XoFINjRnNkfhssC
ENcUm4x6Mi0r+aXBM4Y9WTm9+LNdaUFzG19CfOQ7yCmCuFlZqzrYKSvWQO0r2lUi
YTnhf/CpSnUyBKdWLxCChbGU97Y8Ntnb/ARUmscGOAHi5TBRjYdQ8dwa+3ApsapY
pjYBziXG9F+lYsDHd1dB46VVwbchVGuRC2ZmCah2z9K5AlkKCKmAxRceMxHl3ntU
hANtO1NxzIdS5HrRWkUnmxjsZWRXHXB+FbSMTmRNHyvARKaRlC2D2jpzKT/CHVTC
LzpQufrgP6jM+FVqJQe1641f204LfkEINDIHh+PisD8GZF6GgWgR/v+U/WiZLmHI
7/Gwnxspndrc8qVQA3chOjnpGu/1Z/zXdrmSMIQkG4ThuER8/FRdDzLltgr2AYHZ
LUr4yGES12dZnLRJ6zAtGruNx5FCfi+dhrOCFD5tztX06dR0QKC/r0pbHzPsE/qO
DWMJ5aMa7z+XGjgb3LK+AoqQMi2giB/duwTtuS2p6P+9dhkXrYMZCPANf23/AVAQ
K0P0mmIcchvYLPbUF2mc2o6Trg4bAe+CJC9RqmcZOvaiKey/sDLkXa8FZmib2ApY
klPNlIKBHEzwhUSjEekGbnqlg1K0PBVfAzurVIO/OA0EELsClzbTrEDrdjYX9bVj
3YuIKLJ2katBWZALasYFyrjYDlqHH0us11jEqKXQPtNIpV1G+uByS7aEmOqAIwLs
kG2NhR3RkUdqoqqXQDBb/tZgiO42U8mdZUeLPVaHhp9PBhYvDpaOe2px+x+hpRQB
8mDf3XpUDOA2XMxDSMQIBpkfrW9cPA2k9BRpnk/OlBYZUtkdgVv8eJul8yyjBNVg
8i0OmWg+4owMy/FKVmM+xxVKu7IROIvEcBIdpNekEMyYhRSaNwhjc/jNMcZ787Sm
64JmVwir92ZIuHLkT0topCujs1SbSBY/1nXCyMTJt0M10MdcHjP4KR7ZBqGbuxpK
HdL44IcZVGq6KR41UDgCZt22wksGWHYMho0TPEH8fQEhN7biInLf4YGH9iobceCu
eNI2jb2q+APSy8cHIezDYgY151A5K4DLmXI/lWz5wwQpvLFQrpY10OxXjHairVOa
zdduFvwo4+tOkh9LJWot1qbVdNUWJ6G8sHEuU/AzB8+pigXO9c+HBSb91aqW3mUW
Ajy/BbFp7UmTBAfVQ1FWT5dWD2JuYnWUlEMqOe8LtlrIjtBEOIzmhRV8OX62hNox
XwqDhaUWDo4IlzI3o50rgi8+dEJNC10zGZSdcgvRoBLAUiXYF3lHQzhlbWM65hzM
jZC7RD52W9qA6l1vWaOdlT0f2Njb9rqrtdfvRcJ/IGITu1xuC/HoKG/ktIvFZcjp
q4QOviKqfXZ8kerSyIsT93Kjw+We3JVS3Pn9x9XD+Sx6Dd2UxOnQavPMKhlS2UU+
2Lg/+a0ZDqZ2iMYW/0gcjwaBKDEjKswYMge8zdSSbyUVtrl3aiD75vy1YjDdjNzs
PqwU95YsJVwmKR9W/IwqPmYErinOZ9QYXMiIDNJ+X4B6yxZG5mp7TL7jagPWjZ42
YtsFpH0XFURlmhJPeIjqxpxr0ZPcy6GHatNxSL9cvo2APTfsfXlec5aOs70JT15L
urBga+ZUQNeD+6ZqFAZ4UzUJHSGMeL+0qxwWMh6U1YoAYLEuEhoDcWlTXxAmNgTE
Th7hvoG21pOXJT/3b7vz3UETrwndwGssb0LjJHXgLHkbCBHzdknGljDOfLCvYe+P
JeJmB+DJN6LPVp12OxoMZxwv9UVYXT6zimeu+PsADJK1FRbxMgiRy044PNtXyvfq
op6U4fTxEVYhIqlNj7qHdWSvRT/I6A6MnqXz1B13l3tyFMYCZwWoKINUcXO5ucpi
Nmi/z000jL6QHdmM1UeLQ82+7bywCehj17jJUkxcUkRk4+g3dItmiusnN0UqEAB5
z0L0S3dWB1BfG5PpntA2SHHJEGE4HYRKzpnqZpKCh4jmKtTS/gzCJKyX2/IXh/k0
/5XT6Y+LDaPJ/j6T5FyQS8XhXPHXE6MkXbh8/rXSEXOpIAGGJrkAhUOUD8q38x4B
NQwPZw4F+44l6UbQIu7lWyeiifWmGacHz0WCj+eOw6zFfGd3o7tyGR30WM4Jc9Vd
ZD5MKu6+BYqxmJpMGaPU2qInQ95VwsjhTMnPPavJx6btClzPfhcT9ia9F3qCSpaU
cCyp0q454Rzgca4IgoYVxkurM+9Yl3dmlTPHJTdvMipuU+XrnrtOVihBFSn7YzP+
eyB7tkOEWnn3DO9Sk3tvp2W2w63d0gGuT7yeeea58tA7cTrQcr/BxCiPJj+l6l1h
ySDPwirPwawD+EvpnyjjM2ORZyFI/DX27R66/q6DvOZcKcMlGkNF3/R/rDOwt8By
ekYz7sUbgHHE6G0ew1qZVhvJ6hW8ztz6vIyKXchIMfIm+zjmkyxGxq5SjSEdQkRr
KmlkbNz0GLlPE/U22HtT3BAefRYeGC6pcDMiKQ25FsZKtThOVZO5T24muG5H01wj
YMChbLrluoFEj0hfGGjTnq+1N7MQZ4Z+ce49sTuM05nAn8hTQ3VGIw19fC/TaFz1
S+190gdWRrcPLWD4ySWBygRfZIfPcfNc2DHY9xsnfCDRSWiDKHqTbEt1LYd9REMn
vsvdJk1rAfXRxIaQdptN229XFmYY4GklKjXMh7Aveo8cCCshd+wNL6FUASTlenq5
hUaACt8Vf1qyEp8qmPZnwSQF0SpGzuFnUlJ1WF9iZv9StDkpFw1WwAdeuxqtoui2
tzEqUUXw+qH8laSDfJj4pqiBjMe5U/fRTlVbpmCOjiKDuHVWSxRmD1Repfgv7d2A
bbW2mapj5X7+0jk7msgbpgBFBxwyu/TNGN6oJVgPWhWD/UV0C7PTEnoMMSouGkh9
Zmz21Go277TpnCqFM/GSNN5EIvqSrTHVzyh6Y6Il+3R1OSn65YrEuDvgklF8WsZF
gSsRh9lRV0SsSOO8XR1rGwqaurWJFoShe4UvD9473SRhyW+VNt9J+KjCxIuqobJH
4jYtdW8FIgZfc0O1HYh7SCHP9VGUf08ow1w3WECPusbxYDivxFFYOG9+YrvuWf81
ZiYgNbiLgGRVtBa12C00PzygxycYjsJA8PWQ4/Zdq/Aavs0krpZzk90buJvAeoXB
otyznihcypWreg54zOC3soYzfIgJ20UUX/gJf/52X/axkW4SPjtJ79o8K8JBVV84
IHQStnY3U/JUzBLfgC11RhIgvzzbc88C6hKYp1G2uFVsKR7KTOTp6BZ+Sf5j6ZtI
pCXjNAyFnYaenkDT0RUjGeN130ROTitoDdYL9WenFcBvkMrAnzAeUiMGsxsA6rqS
Q4bJS+FDrQUQFOHXIPyofcJbXGw+EpYfR9oqV752sn2rwFNMqVohL49imc9A540s
wmFS+xPGTl6vaJDNK6JKcs5zvnv+5AdQ9fy5Ogj17X5JDqGDl8QAGrZ08s0gabUp
JdgNeYR1G6+QAE/3TJa2VFO8WQwi4SxiWiqz3stgn4cFLIzbPMgVeYeZ39DYLrQ4
IDXqHZ07oodK5QxgbrYnlYVSLYqLVw1erAs3bxav9eosIBAcSYr2JDOW3msXeuI0
zUj61oA9qFo5ugMNjhyUlSgGhUhi5TLxRsPoH92r3t6QMg/T/m4iJC9jz0krTxSW
E/iD0ziC+7MEsRMnmA/4DltA1Dfn8FUbO24GWL99UNvzrKDiCi26ELgo9jW6vhVz
y5mk4lFIj8yqzoqx+Ix1pGsulWnZDRFANIFkf6Em0JZ7NDaT52mAuqnj2SaqD0Xd
Aha3/OTNXbfis+U+xL1PkwLUSaSKdN3V3+SxAlMEMwE20KgGoM4GbCBi6G9gjyKr
GfEs+ELcseXLAwCCS+ahMskpcc0xr9J4Aa5X38jv/BqZjZ/9l7Ck33u3fFimXgkv
e40XivCnbqbAW5v7xwq1Ot29QcPAkVFGiF+b568r2BgKHPGhgXYAiGfgS9BERmNh
ZmKhxEMs/adZFVZz4VX7xXkd3msbfTTE37RL2KyIXbxgbDPKci4Mxz6jgQDRW15Q
80rhcocWOlKfkZNATU6gG0XXJI3YxSR9N+v0cboegJtWIY1CLJJETAO7pS1yX2Pf
T0XxRsnbjGSezMc93kI9F4SJY0wF0wADcjafE+aQ/O6xPQpwEBOiTdeKVpHzffp/
t7uEi3ttTxWnxFuusMZTDI/7fDtw3q6oWZPIpfqZ72NIbdLae2KP6h959HOOvmdv
WvZjmk+DIPaEMCToRDUT2ABRWmXqB/fT/1t3QyGEx9EMv3Aw0YhPqiWgfKCKIy95
bzlFmn3VSg3qtaZyAJ8Kz9aBilJgZe+65qj0S5L3joGLVq14IsbFQpTtDDq7lFL1
D6y3vA6R6cw4y72iPjMmL0tkE9CnoFeTaU5Ad6rdGYe0LU/yhVTngvrAHG/SW01C
qQ1YSmTOqn9qUbNRIFsZzGEMcpHcwPqmGBNMIwBCN8CQ/pH9YXpIbdRXnxfhNxeC
p8YvF4SgWpo/iUDKtepun6QYn177yo1eBDfRtHIbLP3EmMAaU4XlhJ6N2vPAUphx
EWHReqfQZZMyN/0BmNnAppbwIF9YvaVq6eYaLD7OIlcnKkleowhwvjRY5csU6XY6
y35A7jLb5PzfgjJP5NCTaV1v+2fhsk5mYXFxQh/fqQkOlKovLMY+5I+LSnbAuc4Z
IhzUCMk1yj59B1f2HfhKDsG9MgoNviTB6NLVoWv6ftf6/F5gysdPiNejlYq98WeO
O7fjDttvfRCpeTmi7tvVbhogVA+yLz6XWWDWjytHS9jqGNGp0Mxt6BZeCDhX/fmP
KpWqjjEYRezBBPaTbeDDmFgNc7QCUbhLcz8WSWM0684ldECSqQ5lpDwnxkclhxJF
QWUOWfX30FEXEaS0O/4p7M92W7gvelsBPuRHcio3ZoqCC1ICeJL0CBBDRGZn4HHw
nsrNSRoQchuV7GgefOG0GpgfwjKXLc1HMpGIZhvxZusEapN+I5D2lCC64xzZ6wgV
CVN3dnkM+SNu9U6ksrb8S72qIRJ25i5mwAVjSk7HJCFhnzu976Ty76ykHGqipjoZ
oi9ENeWMwnyL1M74TuPP3tykNF7ZjkOhWZItjMYrmyvLrfOxGMFCjxZROywlEUCA
xzVk90zIj7bKUcLFHGLAfMlGi3IAjqL0gPPvmfMgkRo9TLgeUK5rVKvZ7UgCIIZd
JVcb4NO+CX811/j5bc3gTYcUkEre51f0ctj++Ldktf/CviQZy+xeWE66itDnVyyY
fAFCfY7p5gakPSSZ6+jI7l1Equh7B1qRkDVoJrZDd0cMpGEcY80Y6gYJgTK9mnNg
vO14u0rgL9Qk4WM9UvLQ52iazU0AOuOluwjORf/k5odhuxNyXtMxhcl+iWLzp5mB
S1ORYde2HrwEr8LXbh6TK3TZPrwcFx7x8fJ3Wd9S6OimcAaGou/2WtJWNJ/atyji
oVqkposjIY7i2+0zL5d+wFn8sKmE4kDnNA8OqLnwXDTgTaQR4nw41xmqctWXA8M7
CUqSvG3nR3FWTyZ/WqdyCN+VO+w5SKAmidObIVVXYRIXvXVtj7cig0Si+GyuRoFJ
SvX5/MjUcpmIX9VNh7hseCAXxx9SEdkJK8ku1756F5nznedapwL1769uYvLl/IsB
W5I8yruwie4QYGMsn5hIu+anG1WXe+3im6yn3519+8NIlDSLLQ/RehWw+EWB12Za
/Yoy6Dz27c3Enr5HMUtU9bj1cO7hkWJg8cpwCT5p0u/0LcBjE1ysIB+3GRwDorM3
1OJzDtMenSI/W6vZdlxg6UsNNWNYmtukGUjLmbSB/Mv3Q0kyOrv+GKlxc9lwYPDW
KPvNjhhkyn4BpqBD5itR8V4F8nQFS+vX5akBXtVSjviC6iITOb3vHVUBZUAzE7AB
nWUlehtfc0okWDjDUbdFAX0BTJQyl29r/ZLY+hZ2mT5tOr07ZsIpXGcmDJZpIAK7
590lwBfB3HkSJ3hNil/C+PK3+5wH80mLOnCNjCcCaAdnAZrzzCo051/K19DkCwB+
WJTWuzZXFYf5JWMVWu0C1nBymZ2Ydm6Jz2NkOxgZuJwNOLyqwtady0YtFXrf1GEe
HRKYVDaarIb0/M0Yvd8VYLtzJCk3D78SWY7fSsTeO+JV7DpLXi0kHHHH4Dq2KAFU
FlMuBETf15c+Jht8obZiu08K9agH4IP9X27kdAtitwSuZQvLqnoXZQC0Kbcwjd7h
iazECof/ZS0tNrn0LIPeLZNwMKkScLJvdlbPGfHBsvWbGD8ka0IXHLmPsUz8ZkGI
wh1eTw/lkwIyLdujILAGkrzgn7rbdiUVLpUlM0BjMl7gZomr03v9O8bZoFnJsJU7
MeM7yne1nA+KOrAC2WdH/ECQp6o2kl2mbU690/8NCS14hWp8Rud9EaQkd2UK6bhL
ZMyQBD8XmusjoFP84uh322z067aaYEgqS4lWixkFbLlcO0QAT5T89O3p4uvy0ZXs
4OVcv76XWHX1Mc+u+xCg5QCsqbp6mMVsCgOysNG+qerdPyQzHgc9sSh3uwahIp7z
omHo/Wq+eZqNmMdluPJk+kUoNeS80fjJBWQ8ZWnZUUWZgrDA1q5wPU6A/rqZ1rVI
hTImxLaOLOrSN0kGs+mRJRmm7ZSs7ccgSriVd36kYYVjfYaeANsBrhKgCLktIDac
fxmamBTjjGm7vZT/CgpabLmvqh2kPtEI0qT3A0jaVYcI23BWaLYSNiIepvC6vJ04
v0vuWF9nHF7I9ul7jowwDkSPSND1GFsAPF+yV/m67ItT7J1OfTVEtuxo5DNeoDWd
Hz1ZmoYHdopbytFwj8lyK+mfM1ZL/0HfnN8TqYN2wCfCApHUbDSFdK3Aef3Q9BBW
BPJTQmrY2FTtl0mFsf3/ZjFyCBAHq1TcAofnJaaqJB7As1W65pFtD6Cj+8IcOP8S
VhSUrXF/9NYIXFfgWAEs0izCrGYcYMbXA/queTqXFHdQP7XGC/2yyW3tXkaBwzDQ
OoD+h1G6x6iwoCt96BbdhPtELtBB7SPIiih50XIXb5MfZmCjP4bQ9GZYhbpR266H
pZQ30yM5DfgtSijM1afdNjK/W+0wHpllaSn0cCUzfKmohOavJ6I8I1Dym8meAXa1
lT+NmCRsJtV4PeMU0NmxrU3IS3rAWdck83VHKfzA44yJ1rSTn2FE46BL2bBxGn45
un4g3fki/0/5IdfyAHnL+BAWcmQsMvjnhRfjIxoTbm32IQyskS3302Wvp+M7/cdZ
w7SSSk2HRvS3WTL7maiRm/gns7wX3Op2+03DJ9xa5y3w4TMwk0Ouu2tLFKd7lBOe
3Jnmk3QHtId9f0FUFK6kANQmNlJriuIMZ2uGUJF5QvLemNtqLwlTMIvX73ZcT6oq
pr5nu59bveMvTxuPCZe3EwhTAKPQ3jFn/TmAIJmTbl7nVU49k3PaZczmtndPGhnb
cOYURaI1SLuYBGSD/kGo3tUh2it+LvBmitoBaUvEqGCd+3KZUGnLlL6Vp6e1cEz+
O+EXHQgiS4IgGWrlBdUsAxU1UTnGc4OZNN7wobIiXRhy8ibaip7TtG2FQnvdl3UY
6gm3djU+6SHwwI9UvESjcIoplomqWBcN66oftHY7oJV6WxNb/Hi3pvMCbbbbIfX/
FubMOt1bItAKzfyyRjh8QQcPxxntsaliX8XDEFib4APSNv6wVP0oRs6oSFu+D10H
A23bQS8Fy9eumx8tChBGf6RTjfKOWsPY5lc+5NSGK+4wxUUas/ZkmVCwfaomA/Xi
0ELIm/r+b3pzMiSEYjPjcZhxo2T2Wk2CYDj1h0Tfh4rZ5e4uq48cU/1VFYlHtzOb
JXC1DOehAHXgLNvwm7rQFaTZlzCSsI/aJY5EOkdxWCC2XF9XIQMDVfEn4W9yQhBD
UDaxth9k4KiJXrorRrBkSgCLCTjjbK2ECHnxVXb7vQVSMWPZDavy9hSjiTnoIAZd
5nos5WPKhCEiGLyxJYY0QXv8vzWXe13tffS+W7blnuODJ8r6BJAOllOa7OXk8FPW
8vq+ECSc2ZS07ySi21DgaHwN3bguE1KQEaYb8LjO+iBO6PZntwEfsUo5PmgpQWPu
7luoRDcMcNVQyILGEqMqCnm2WnBgcJzbq0HhR9db0GuqGfQxmArKove3xKU0U/1M
FRoRdCQoY+kzbUCrOxceaHSSuU+QuVy8nfQl4jlHfCeDr7dKxrKywWCequul7coN
p+WS6HciNKwaP37NErwY0Hpa951kRaxwyaU/FZ9zGdu91D0DKR8atSPGPR0a38Cp
AoMu0oHshlY7u+vPBQnMSHiz6mqqL5YFMl0PboLrOpMwuGfMnlHNpir0o8xMNrr6
PJcX3YQd3eT6zwQmxOOu3XQpGhSsxyrV9iQM9Zi5Ho3s7OkmjfAvEIsr37F+gTY6
npgveYj292SXzYaecYpJerW7fwOx2WHBiFFkezfvwonzHq2jCHvZP8sINE0FCiaq
+pOmrWlWiNXmD5ntbzlXbaWKI5DJ4cwUEWWP6ok+WQRAXNVgO+S67wBzuzwG14Do
1mn6p9354itAh/L2zmpboYU2QJvycY5O3OuUkbzcDPr742HheLtkk+5o1DJ48ua9
1z9AcFPfksUck3Ji5lhO2HrU29VqZLk6/sJGs3AG0oIUY7Mt/j8ZU3iBJBm4tMyj
4giybSINq3njMN/G8Jz9ivDxCgh16o9bQ6uS0dQ1ykw=
`protect END_PROTECTED
