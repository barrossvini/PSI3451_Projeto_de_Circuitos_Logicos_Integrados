`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WqNWqDcGqR+8ZOkZsbJDcyjHl3mtYK84lhKLEGZL1pVltFfPlLgyoeNJXa97yqQz
cNjcCmosdcoQYEgWQOKZbY8MwRestzvFByLq7UwiZHiGA2G2xP6veShVCP/p7hmP
0ZgXbUDlPrrBx9Jv99UBCIxp6KeLa0nmJpkkVY57vqy8scrFi/iGPBsci70UeIi0
slBAhoNCNXCT6Mi63sJEpn9Vqxzua4v9u66zLYCY8p/5FaQDSqPbFwi16csoVMln
OlVXDn3BC+NTPpKg9H4XdUjYRaKrnnbKmEucykiTxM5+cZdNbyaeAmBpTC7j4na8
woGdZCPR5bhDgPqx8qAsUvyrjajAzyladiSQrFNC4qJh4v6j/25OGber2pznYi53
Mp4lph7UZpGgg05UgoYp4pVOdWzi2rc/X8yo6199huYTkjYXuPDh5FPQ3Ct1jdcr
DZqz9sx/cYtpF1DrkOZdy3bzXghHA0A2cNne5VpKj/9apEKcVbvhmADjAD28Weqi
KTHH/uEd8+OnPPWjZ/y6sR5E3DbXn3Ohdkam8V3nV7ArSM4M4C8BuylzoSa+0/Q9
1DlqjJQbl20auZ5KJ6ituXLJPQPmApPnxd8IQ0nXNkTn6vk0zxdZtaqm5LCASf8q
2fF6t99fQQSfumamywhE+i7Fdng8Un0rRYCUqkHIqLWbToMKKs9Em9UIw6v1XXBs
CsPjz83jzKKIuISWhzBh//5wPPyxByEPINg7TDBtn+6Vz5DFkEukttOGawoi2Ptf
oPEYAtQrp6vSSNe6sqRn3JM72ZtaGMWNRQdMX/v2V2CBHtTN95/In04s0qcd7Z6+
Kf69BeiSdFVpppDJCo8zTCbU+y23Ia04hYiu8+LAvAgT7potT4SxxBgcS9iE3cZY
NqoWlf9U4I1/8c28vSknPd58FsdLcQaNjX/fzY8/N2VjMh6TCZHY+R/0JtQMnmJV
7haw9Nh4PqXKkcEJpa/SDM3sw1rLfLapZwAgVyxuezB/a3GXXQZWTcR5KvilIIOA
FiK5C2NBycJ3paQ8TxMSWCUaUdGWo5k6C7YWDcb9Q3U1MjZpbrkG6Tw3Gwvk80Gc
kGCqOIKjXCNtuOZF22juhFWXXh7aXln+z63zZQMqms5b1TpHGodFGDIKC3FOdJQ2
tRb+LQQv7ivdUpTRp3nj21Rw6kCjuPwwZi6RHBRg+cgjfv8+vMd+53uKNEDCYaZ0
c8kt4Am0ozGx0m3vEb7WQafwH+CDTlXMpTyMCHCF3wa0nMEXhUUe1ZTbHLznCunx
WNHmR+OXRcPnXlLZnZ71q1LDLoeFCObqeU0dYKkhFTHuXab10gIYH41KnPyRcBMy
T+ctTim9JZXfG7evLzbJ2VcbeRmzJymE4EQamBjg3hoBDfrB/67nG1e02qM1kIOX
6F6PfQjW85cCd+ea8JDNH9ZgOh+dSTK9RvclaIxsGFToDa1Oy4JEuGrntFqTP1lY
hjng4w+O3vJGSG5tBSN08p/XC8oKza+SQTM17djRgwt6fLop7Ys0dbGT/qfqTTHj
KdgQC+mv3G0vYvHKKNyKtjs8I0g2f/U4WhJUwE+Tfsrf96WLdM5wqkdRGhkcuqJq
TcO/acfDW8GhslQ+Apqn5M0RMIXE4T0YNNZ85dbJsgiYI2kLWZmZSDtZawJWMiBe
jeFkM9XoQNVfGHFklAC+jTjniA7TLBoZkwYJcpISoHM4B+KPiPlEgbnzg5O15p78
VNWkGYn3eJuhMrm3EtxAGOGyUFvwfyWM2ss37hwIvMh62w0dvupADI69hUykaVUz
gYoWQ3o0lhT6TCOuwZARhfXrzI6XTreyb+jWPvwPyGAETv5fhmiG/GgroEelXS26
WLU09OCiz9ETYn2I3+6RWxdQ5xq4J9oXMlq5pYnjckqorxaKaiVzz22KzflpJEdP
hDNMLwxOqN2ywPkUqU+skGoutBg8h+Emew7fEi1bVs4G2jiGDwcrOT4OsFo6m3QP
VxOf0hxZdGDmDoVLO9SwgPLO4KBcFT32gigLoMLIFlLVg2ovFREHwB6TLOgnMWqO
CjG6H8oHRowR/JWPmpPt18EmWnFZU3ktned4blIelEIvWemqsH58jg8SpUI/bVRf
hThTYjmie3p4qRVmB9WtXIaqpdWZSDa6TBZ2Dhz1mUa8GX/bcEcI0klro+Cj3b+x
7NLplYKwOTakFMy2WsoNQJZWkzVpc6vyDnvJwKeIsz5ZBxSxe6aqSv4kGwpSa2CL
rFf5UAsgNGNn9v/Cg6emr2l9VmGvY7w87Sp71YUegvijVTzpAMybM/1hX9aG0HxR
dn8YvS7PE+XlFSUm6LFMLXek3VJPc3PlSq5IUUpnNT5zTgaN4ZLwjgXYceIWBJYr
EEid5TvZ2OwX6Zrd21vvzoWO/iwfxeVqkSHieIzp0e+O4nghUWa3x6TTNlQMQiQv
EItrinPnrPtm0ySB0Ek4BS7rhyFflPhTxSDq4EhMbl5WZKSMXdCmGPeqIOGKvBIt
QJyF9JmbmP1RYabcS0Y3E/s2UIXm4UhHxjqywhiRp/1jeLwsG3ml25yyQ/q/3FYI
nnW2Ol9boCHyptDOLu9sh6HZmHdZxedvXc7Y6SWScZqlvdfpWHJ17QSYtx36Q+MF
pBap+5jrjvS3z2WvgEw/zsklB2RBqM66qiKPa63hsSe2r6bcGmwrhnjk1mhvf4QS
c+sEYR9RUCl/FYcIV7tKcMLwXCSofOkFVXVXYLPZ00SI+jp7MgBc3mYl8GmeySPb
6QLdjCVsDv9ZFl7tyfdDiferxP/JcipSQUfgWQ2n75R2dJ0VEFWAiBhd6hGZrA1t
5X9r4yCYQ+SQGhjXxjhh+PtjY2E8ns+7ENaGArWSHkYcbTM6cbSXnUFdg9pb8BFW
ChN/syzHAx+Lb4TtbvNwYeTmHn/PLZ6qLFLKrM+IH68+3EPkprdQBzRmGBqivHOY
FRukJCJAtBPxp0Sfpc3K2SXC952xrpL/O6iwW/OaJw9hF1g5Lqx622cO84qA/eUV
99rJv8hR7kWiu+91pKs0IW9AVbU77I9bcB1VFNuAz8HFDqxDCd3jRx1BWOEVOEcT
KPAYsBKA9C2yYagXkiRkWQrF/LT/uCBJS4P5JPjrqf9UupLm0YVzodnQglK9MX3i
n+ULbl10x3Kq/ZiJA8tLWYi7Tohw0ys1m1ADCTourvQqV9v/KvRuOjKG1MlFo38r
5meQv0VsoyOfUe8OPjyjzoibane2VOLT9U5jazb+TvNgkof5pG1NkadtiZMQu2Ab
ilhWNr63Y9InIu3/xXQGFV0DB78anBxzQa93OIv2xB6BNasUICUGeZaX1+I7E6W7
BI0YL01a52rQoMpiRFtxnIHrstFcXAhQ1i4x8UB07iBwflqlSIyQLWV/mCA1g3Ud
Z4Kt8K3HyZDfY3yRTU9KYM8JxGI92zgZkc6H0cm5WhwepPpX2wkdkFg8kjmREOAe
El0YGx3I61OaXFaglTlcyJKtF9N6rij3EK9jbk+eU8z62RpttmseSPNBBf0B6yVQ
pJwMQ4RjIMM0gxjJX8PWdIkYgLGv349RLmEVDne1zGoUd10nHGorZbRjQ3NKIKJu
ZHzpc0H9ktOLKIXNzHqtNywHpYIVsAgc4UT5tDuOBnoK7G6k5U2r6pLonTShrzUb
xho6UWo/X9FuBmc7G+EJwFVZKQhOFQPAZdg3mwbi5VSies3q3SiZQKYFYbv3ntEL
bgtt41wV4n4kua9cX5+uR16588d+d7ySxDgCTp06N82iddA+J9e3JF19gucwtkw4
YNKvn3n6wObQGLhSj2M+i1+AEN2SYJj79wtX+jyFY7IlwGuLMVvpFPceIae0efDz
nBllQUKFlLzRaAWFEqfU20i2nV4ESYEaUotDidkR8U2v5qa2IqNrRyISTU0Pl8Qs
evnBci/HXEEDldtt1DnIn8zhHc3/he4I43jL7l8xVAnnfkzLF59/mc0FIyDSdy6R
i/BiahQMswk8p1h3JufbOh+Im1+iSqIyD59pKnfzA5V3wqSAOEq5pXAzIggh6NAq
eXBJ/CXDQ8nwimWC0Ig0v5YcMfk9rDx6y/46O70+CFd9ttkof4Aq2V1OWscG9+10
0liwSF1BrGwmHSw36eF0sDBDYt+4TrnlCCT4490st8bZLiCbO0i6flTENnkwrHbd
nf2lV78ZmUt3q/U98jEZjli1szCCdT3eimuNw+nvcoM0sCTOdpDWubBhVYPVAIGL
X6tNSdWA+8T4T/ig1CvHa7NGgL6NFQmobbqYCNqKt8iHlT4UEg7YPeb8S/Sd2/3H
qbJ2kNiP46s1Md5CTJoR1rJGZcIyyIpEr/GMNyVsd3WFK1pw0ZNMznbwTUkN/LwP
tWJ6R/Aa48ZwEu1YTSVf+Mgc3LtLfuVphe3Y+4uqohd+NKG8oxzSwiemI6tbH2PD
Ho1OQVJX3lYpANki1wEKNLrISQUedDKuaoRXsdbt6BLYcPyqhaxaXHFbuGwTYjSB
EjzY3k9qHhKhDo9U8NAVUOk/uSxOZ35wTWda6At7yxtyzhXr4NH2VMsiwPD/6zRt
4rvyXKeo+gsg8o0B02Ev2UHx9HDPwi8saEqEm+644YzXWFopPEHoM6LyQBvRgfnM
lOCN6NQgZhefMzDRT0aiZJuOV5FU/I2rAN3ikZQhhpRolYUYUR80Wi/x5y5Lk6eH
rSfCG1XKjwGso/rsvVnVO2QWtyUN9Ml3Our5OKJGvIMIJbABD86nJLkbsvCNkf+y
Kf4jBAfqcviReWoJvmxVUuw067DCyLgQ2fCmbY+FTHEjOTp9ISZvdT2kdO7EweqC
8ogEFZU6ebNfi0iwzKPudmp3bRXHlbEgEtmOEIzXmn3lEG1CZV2vQ/bqnzMl/X21
btNDqLFkQe6mZi/dgPL76gFpX6weP4R0fLfkcOdwNp/4/KVPAWIO6uQHoRGniDgu
AXx9Nhq39mjvZuG67Er5/OwurtsnhLpTfXrDcXp1Qr4x0fb/3JK22fbT3aw5yBxi
EuQtUsrHe/U0k+iLW6bkEH5go22oH01Bp8xRdKHYwWvWbGqL/ErP9gl9tnuTaX4Z
MHuvTjC9mckh9ip8E3YQqBAhRLVloRK35nEqrWDoyVdFuAKWQL6HxksBBCqZRkEo
Z+4/akEh+Ax53y29C0mB6pEK25PItvqjTyl9XeHsMiSLwBuAYSngRJJEy9Thf/Cx
5mWauHNWvPMdgLBX7uKf6DVR3Rf6TS4dlhnrTHcL/7UJIgVLAXGRsT1VWQTzjYiD
nQNNbCSUhRBbRw5P+rGhYZDRBvRbUvpAcr/VxldvRjRkatRxfL5QC5ep2PZTqVaB
nLEQ0jWvNkrjbypTna/18Oqb+jzBOCHxkT75SWewovTZCc+ynU4TQ0D39sP8DfkK
UOdQDdK7P1J0U85GQp/uhi58be4hxuJwTFEwVmk8JFIX178A1aiemLvKBCN5Y9Ki
E3HHkHR1AMcnWR0HQ+R43h4lBtp6/Z7MAm8KGakSi6549O182PcRxznQW3zY2Yzl
DaNIJZfslqzWei04unInQJEeNj3ZTysRt0jnd6wmYyP8JLAWClNp9lTx8psyEbTa
g65E1/Sm1qbTglVDI0kZOtTKbSz76n0MKqj75Owctined+pG68xSuHacM51kJ1NE
MPzRjyzoHnmJmkmDdoxVISvXTcOvu6d6ofYZyjB6JihVVsRvHdZLHEErUY6C5Mqk
yj1kyQxzcZwHlKQjhG55NshQXeeeMe5gFxNfRehFV/16ZSYphtwuWIhz5oUEvib0
+K7bb5Si2u6oI9iOuaN+3rfVvNuvzevhpluQoNV6O+92csxgwfQymcaehjakdD31
PuuwQbhyfBa61qemf8LBFYMHu/u6OsJsWzAfYy0djKY=
`protect END_PROTECTED
