`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ChG593FTA0CIbU8uf4NYgZAuJtiB9yv964/dEFdrXxEny4QaYgpSGD+3vfLdAxyx
1afY2twpbtJ1VktybzVx1QWChF5Pm+1kppgMcm6nWNtQUDE5686jWBTeH7BvTTAK
sYybIlQ7XW6J9mHMfeLfE/fbJ2cg/cqOUya8Zrt18fq1x5gvyOh4cpgOwJ2qFdjv
1rdIQteOlaZ5m7y6qfhilu7Xe8D7P2n3cly91fjFqqyhO0cDTrmZQIKe4M8f7G4d
62wOlIsTTy/tZ/72UWfL9aGoumGJ6niZxE9dKNh52w/8b+nwzpaL2czYSMkbw5kv
DYkSWsYpJw6Hx31jBVQsF2HScGzcSodTav16p2tECze1QUlTcMCgF6tskBkltvQp
IeIyQb5erTXuglBqhmP50V7ZHgsv/fD8a91tTPk7hF5VqjzO0zPeKQYWoZagE4fu
MStsU0ej2huG9SleX1v82Qze3AkwiptetYL5e5UJw6iFELH7YDPdCsVLWlcToIF6
ZGXtZ7VbDA/5Ssvkmu8jZZb0EKvGjQL8aoeapwHC24y+WGRfqtnvAmYI7LIgkPFo
ZuaRv5IHsshAhMjHM+tJNY0GN6a3Kko+DoBrYkgKbu1+33K3wc76Suk1EExs9bOB
3HAOVHTyehVjfuwcDO/NJgL0rAZL5RRBXAqJnPf6XCYmEPGjEzw//v3r4es2y8Zf
Yl9Ns8dgjysK82aajQ9HdV2r+/dWDtWo38Ja6FlyH+CpVWZRGtfiUSW+LeTDnU1V
2YWOJRtWeNnJTAoV9bMPIXF73Dd4casSKjoD/0Aw7/NgeP/n+KaMcbZ5k0xZI5ga
bXmQhf6MVKv3QpsQKJiNhvVTBYa2sUs4ujCfmohga215JZN1jTbr+i+A7mSZYisG
Hcxo3cCsvhm4C0lxMmeEeIArP9ofim6nQblwM8UHlkjKmsLUK9CCBaFmoxHbIhbR
uO6ed7dn54ivENPQemxqZ1Jh33TPhmRIg1E1ypuYlI83dV3Fs3efBXUc8u4r8rDy
rmR4B2xcDqdSTEbdFTYuD5Q4YOOFCdEYIE53CZXY7BfHKs8tbA9b3Qh+RDhp9TyN
4ntSoXB9SLaLw4pKkUCyca04Q8Xj9Fx7Zzo08uFTDrcHrqogSyPewXRZsqQnSjxB
020JQdJ/1I/DutWJjYHKia7HNIHFatXIPTQGuwtfVvtPETx++Y0wB/tvUKbrJ3l7
+lGHGjqrX3C1cCMtjt2rgGuSOr+9nGfPJCn0/iF1PXXdhIZavgl3FUFyMWWoiAja
nQ0iAZlp3E56TpllQZwHdw8pO+IVtkekC16iP1umepQErKOrGx6LXOhCNwVon0Cm
uqclKmO65INfYHytF0Hjh5/eLuz459ETNv2LfIvOu/Bc0QthYllD880ND7kIWBKU
V/zNZBDC6x7Sk4PotwRy9NhZO3UYOst8NSL0y/06dXjhfSGeUp6kjYLScj2apMxS
VwqhXrta9aNqOcmdB38du6LGGUOeOBvryjkl2Licyu3tMFOQ/OodAAG/m1q98fkT
Z+M4TTT88aVW5Ydwp0iBllmREaD0KPofhERLAIXq0PRLFyt/OsRYWwgj2ivHl/Gv
PxRjVBZzBzWHRlkaQxt7Fp8307CAKXF2zXrUcDBpReWIk2lJStIfstV4+SRgazW3
Oe8llkiCxOpjk7tfnvBgdSMFbnhnnsK88lOEzqErGW4pnBOv81o3BzO9bBMwTOnd
QDu5waWhLPBBJbMLPhLWGH3AGZmT6IQSo8zMLQFaaO/PEVTSR+lxIvX7yy2SySXy
5hO3yHXnX5EDAn9pKo9AvhGKqz+6fW6DSfnK7Qkg1xMk46MoR6TnWrBP9Oa9BM0m
Lhw4zPpIfPA3pnuQ5T2NwgxSI9saNe9PDpzApPj+6BfG3d7kkec/oHHTB4CcVm/5
hcdCbgVELoqlBxHyJe6grJMu9Q+/ku7ujzbjBr9WtVqnVT4j0ZTnxXHTjvYJs9qc
qxqYvVrgnFf6mokAo3dqZXrTWU9HbCSdfl3z7poz6+NQwhd2kUMPQv42wvL+m0et
Ji5ifpWVlND9rdh3sHf0nqtQKXbUA3Ehqmlkddn6ZcttXP2mI+oMHqr8cWe5pCmf
p1gQYAHgmB2qKCjkp4irIl33liv/TABaRtznGtAM4OSVwWxkFlbRr2gdTY9fv09S
d03YCCYNHG6/Y9WTH4rZ/hWjVDFTlahUjmKOE8TnNOdNLWYFbEi4HdSJWvigJUwS
DswDvFkP1bEgDgvkhB75RsEiw7sDVqJkf9PD2HccIr3H1LING0fKVrDQUwoFCHQn
f/yYter9TylHB7yBB7LIjkFG0fzz5Wvex4i05EeLPrwPGxQdKwyoHNHGTFYYPoPE
rBW7298jMFOcbL3zAVYY9qcRwv3b9MzreQSky3GqeXeLxctjtV9Q26Mzj86jTyL4
rSZ3f53zgFd5FF12Vw6wq2NpT2zFZDYA0CZagCXbTO7WxmOubdELgE5dmBiWjhj3
hth4vcJzcufRrHEb4CtO+aXth9dphx0AH0N4yrwiMBmpRDDANm26hJ4dj0r+8JX4
fHaZ64M4fHW5dbdtxb6fRojszXf/k+MtYl31/HTLHdzuPFbJ2RXX/qM9lMp8YmGp
Y+gXVxhgkMceD/a9h7i0+5yiAmXy/ak/f36Ez85s+nBzhsj8/OLG1KGmLC1PPNl3
UbTqmcyJs7z13iqxl4Jcs6pzcP6uaUY0YadX6NyDmbrdSvEuB9DDtj7Pm4H1jAAa
kUV8E9AxKwXnpKTUzV1m0eq5Uq2x41IHkXrxh38UDDa1OcCDp+Or0IGWMB+Y1z1f
EB5htHQsBGummTILhngNA7v76O3mSWzs5/2+/jVOGWcOtpraNsT0V9I62ekiN+iH
GwU/PhWk/gzPkC/xsw36ZaV3GYfa7hH8Wt/dgPqWXzWyTNdVP5DJ/6EwvLXbS/g8
sJi7drP/u1RCu4IxFHPEaXaPn0gdZGECWth8sk9+ZFd7rSuDykytJ7XcIA9Qn5jD
mMU7oPgWN868ki74SxENZCRLkwI7PnbDCsaKtLZp6FBy0mfxZ6BVdkrZOGHUeu1R
O1fGEvhdgQvyZclSPbOheV6v5e5y26EL8eTtZkiy063YyTnxY+xe/TY0KMqeZz6V
f4g3/+v/hxH+ipAC7PCwC56CpuqEV/9WuuH3GOePsVU6MFWcvY8+7fV6vOMJa81s
603GngydwyGNk1fQ3gfKlDn51b333Qyk2ZOH17Uq2pOjDLm94xIbPiAKFEVRQxt/
YPoTqOfXw7ve1jTg+OvNqCdRyABQ1RQ+UWzyipgRFt0QwuRZxc73MrtDIRgQUOsY
Cr6hEC5gFNd2t2NmX7iyL1R0nG9387VF18zcOZJp6OVGBeWeLqdGUQ0r+u2Ev8LF
yVqh54Mqy7CnsL4o6qDvmFRQkelbhYLJNOVnEQB89ddjeSWF65qFXCw1q9wsmaIv
24jqSe1vJWP+AIqLeEJ1rq9Khlx9rMUyy06hCYEvHl4Zs5y7R3hS+qKOx72joL3S
GL2COlwPkOMJZ9a10816hgOnex4fXt/FqMUlCRlxeJxnhclOGA9AEGPPz6TNdP7P
c9tYwBIQiL3zZn32RjW7o/CQTRrzUjtbw/uMvZvU99+DRXbSxqddBrv9fXbvKZlp
aBuqtsiMMslBLmqV6TiMA+mYbLkRCqwmBrVu8WSi/bcEWc+jbP006nJos3ht5wRC
Ys5VTtILxdqimVTfIqEqrPpAsF0faYNREzr8DsjrZJ1MpSQHcon/SThANFQ8HQVu
rF3HMHw2uDFonOePPAUbo/376jSSogQZXxkhb0YC3T4rh3iNE/E+b7i/BbeAd8I4
+MFjhDOuU1CBzDG3f7jjk362W2Rgbd8yjH+F8mS22jfBuAatXJDsZ/DtsLDGQKZb
2FYv3Na5uWV6POWuDEyamg0+D7gwBaYYSkebURCQJGDjQOvIK9YqYg65A4W2Rp04
Hu27FdPTCfloIDybFulOHQ3SdRwIOw6gohDjwOPIJu5nQRxcUJFfmkU486Fld5Qh
61vgXanCc5aQOtM3UfmHNxYuwe56b9NegcGx78rpGvJkdQiqm6HKikNWtsYVzSbZ
UOdROtRFceV2SP+pmSH9rRCghM0pO2nyIovehRA9tGN1q4X3VmyVJVeHxpjgGORj
7s0dkK+3CBJMLjWISNJxM/KPTGGd4lSC4+3hSR8YKU+/dKBxwitZMYzZNYQdPSvu
bxiD01e/7OB4q4TKVv/Hcl0uTRgz0k4fKv/Obq5irs5yQWKUxWbwPrblSqgLqj6s
W5j2nivS34xu8sIpVk+ZGOUOtEZCo3iDPn4hB/vH40JvgrGeSIxFHrhONLdoYfWn
UYa7RTtQD2xSt77EZribO2n8/89tfR+w9zVH7zHjm7l4cHX8/aCQwtddvp7eU8tj
VVSBd5yXcLVvywGqlIeChRXTtMZIunR9wdBF6EBDz0WRG9oKMkw6tasQJ6aleXTu
OIdXmPn66fmAGmrS9r8xRN2h/z08XuncssEDEoQD9ajC9tYqL62S1WQ8/92Zidc+
QsLlk80iGZQrE5lvBGVJpfAlN4zacMYg3gdthE+uG7u5lJT5FrpSkGSYcVg2XmsX
yaKu1wCsJccJtCcu635aE4KLDP/g8XzRDilw6lQqiwV+YOjSux3BCee5HjSuaQx+
bbv2OvDIoLjFUzpEnlZbwnkHLbwLFAZ437Fwg8ZGYptUXoc+McV9h2w5+AkM9j98
JNgPsO/TRQ2/JAKcYVOsPK982WseACd2HWN/rl22oqQHTPCmIwOItSBfdYGlSEGY
/WTCVxqyFMOpprXHBEpblKSoW5ZPv5kblmKH3z/q8PpRJVDBXjm1I77ykS4jAIRZ
KJ0w9NVcnIcHv5Qk7kb8KiJWY3iizi5etBP9reKQ/gv99Mmz5CfdVs3qiX6UktNV
//uIwpPguuyKLTFY/7NdYgz+VhGZLwx7XnagDClF7bAuM8oh6I2MbMRm+74NQkoo
UBOU045TvPd3N7BwCWgQZ4GZWtBupD7Qk2hSFE9p87fi6gFEyYRSOjjwP/JXQxFy
HKRFObmcb5xtt7uPi0uCnFPTSXiFjGvBk/g2VVJz9khMCfMfE6LjFuq/1TxIjxxZ
2DwfCT35RqW54EPgO1GcrlLTPRbUAvL0xPLRLPsixBO5vEad2bFbV2BxhQh9t/b7
sM9gvGOeQMYsjGB8O6RtvD+401pPqrTV4y2G47ECBaNlipBIoefg4E76k5rM3uuH
BkuzyxovhRDnWCEhsTBQ7jSfrVA1PJvxajCr1QSHIRNuAlz0+tCYglQi9w3z3mPm
Eaa4/s6a4Gr+s+4NJViYsqq/6lU6/adXtPM1kE3JFN1lMwZcMQF1kSPXHQ5LZzIE
jxe+NRvansdpTfGGSZurWOwXWVMJ/r1W0DxgRvyVjuhMfC6YJvKD9c1oRyvKmaVd
KYx6W7/Uo9BUEtJiFqaAh6MFH53m1m/ye/bANeYjwHVch/WIJEKMYwJxKFoXE5bg
lR6ctvmYZC1Q55ALzkHXSN+E6qSv5jfAMVdXFd9U9vyzsmuD7P+pEe60Hni+eyGB
OtQiUvXuAG5njcMGR7N/wKBkNdN7HsCv5AtqiUmvI64BdN01hq8RSo9hbvzgFVlL
XseJ3wRY7WnwahizNYKpVRcOr6MZHxafAoiYxiuM4YsDe3mWG25qVtYUQuJRu2db
xetL4b/96ue2xkQ5/XeBHYU0Z3D0vAWuOaFTB8eZkaVgOGKGfzVKn5gmBD5AqivZ
JfFBep9FTL9M3lGEOgvcXe7sRQExbfiLlLmy8gbamsCG042Usvrn0FEUDgrnicQn
LsO25kyRsQjwJcdg2ve62IFyZ9D68g/YLdC6p/vTTkTzhyXqa/bwR/MQxYxPkQvi
cb97iPILGSH3TBZufCLEA5/B62STq6iLULvhVkdjLY8ljUu9UJj/SEavNthEFpcr
rFyRo8atJuuvDHKQkXSeQHBH+Wx6cUOst/eJytIMEOGlbuqRfw1910qwGjDFo6DM
ymKYltOEt2K635FW98dXaRVvOQ0kvzq013NqQ3BTYWJrS7OUic4+ylyI9wA/gOY2
9YX8F17+wbDNseB7bptKUexUCotGohlSp532ipKlJjEai88oJcnIh340oXlIxnov
jsRZPg1Yx5MLPfaLLFVxfdBqBSS77DXaWdcP94KmNi2u0xgXSZlGRtUa7b+Pkcsb
xgRJjsEH9I6bxqJ2qn1X4X7AGJwpLopoS6Km7AZT7z4qq+lU0QsCunip0rn/+Q40
d6YNysRMb6WpufouwuDKMvzPSe0ZAyOIchT9NItKEsFcS1PZ8esv+rOXKtR3PL0V
5gqw9jX/+MCxGsvX/f5ETlFvOvvgdxViEdXkTGIHIsP8cIN0cXQyejvcf4rgikxV
2QOsmhn01BuGRyarqj9ui3xDhT/uxz6zEmZN3M4aQDyNQO9v0n6rV5NkPKJqj4qU
gli5i35IkFuvDzzp0W0rtASnmJ4QfhaYIEu/PWJ7UbpA7VtU7khSGWdK6ARWFG/i
TQnzgr3R/nL6w9ZIGaewJ6HAEXbWAcAeUg3ceFpJLtyvs+qTHPr/kChYEu2xc021
gRlxDdLQGWXP1Hd/nRHTO0z4hIGP4DEDfrRENd+9XvllgB5kQFFuSkzAJOjweYTP
tHSIvrd9CKcSdeDXOL5g2koNQEVYc8F4agfGx7Vtxg+fvPAxVa8QNvmPfjCUWvQj
yulGs0IMQ4QhhhKjXEBIEOz5ArlTSXckgQPZAhgqiTVG7LVg5gNzqCMbec/Gf3G5
9KfGypOgFQ4LZVIDq2UH0ERMCOPh79npYw+aVi/CADWl4aDkNQ55GuNI2+BiCJXU
RN6pjDiAgnKIzDFW6rAZoXIV+utlLmmkpTlZApZ2ePkyBu6J74pfZJQN42NX+o1m
Adu/+vu1I1tWRE2D6y79UgTHUq5YmUbOScGQooOa5mzwbQ3yPnL8mJKWNYeSfZVi
i6dKUjKvMXNB3X4ZH6FZk1ivuXBsrqXQG/5AdZLlOeoCaM7NvEQAwnvGFVlmrh7D
/+2CTVQ+8/VqugMWkEh+e6kizotHFuuzFuTsfw1tLj+ey7KTLax+Q6JZvipTMFjZ
9cYnHpAwvN88DUgjBsEq5eAhTQHGDldR5LP2ulC2ZsOX73iAy2X08vQh1X2TUIPB
k4A9NJG4qJn1crSaE+10xOGTns4KswPfLRSsg+7Nzo650xaIqFALKWb9zYc5tUC1
k4bnv2Nxx8+zL1yLiRovJJBgfMnEpdEiz8fUBkhexF7ep/F1DVAAaIHAw3Eh3DCH
wxa3SoEdIIVPhE4HwRIgQApZiMWVFA9Ynp3zbcSbnj4FamH0iNl46c6cnMKL0kjW
fx+X41ZgM2kN/FMcm5TY9HttoPaMDnf91BHG7kY7gmIJlTMpzKb378f6Tpgs3pp3
zTyDYzS/tXFjnXX9VizGWD54AVrjWvAeSgV3y52+4xhqEiHlfzkgn7swNtb213hV
JVihOdSpVhV57o10q0K3Ra8FURYe1dJoOtPPFGExOTHyp0cQzhMEfuwyp5iSAyHX
K/sEhuYLKk8wqg+CgTAGUY/XKNVI2hjOll9R72gGCbsHq3g/R6HQ7pqDzAdFslnr
aEXAuI/mIqnHPk3FOP3Nu+KFMDTLe/ktPzR/Y+IthL622AKamxBuMh7RUpNk7zV3
uFpEGnMkNqhg9P/FxlY+GEiGz4RMJP0O0Bf74jHeAV2uA1O77WmZaDeoaHzVKduz
5VSxaIe11sV8nYFZxX5m+hWq+ZeQXntSbURMqMZrDF4SlbfV5ASo1n4jUn6Ymmlw
cr2R1/UMno3G8Eh99LOZeKqmvfHEZtP6Ah87poou+qWgL8/g3uK4e4gi5vtV3G5f
7s6j1k6JutPoKpOGOzVGXwiJRxOEMnSUnZgFOAKcsJn0Zm44bGybPsUD0JL/4tRg
+4wd+2ct+AYtwm/yVVDsYAy+YrGDcAwjkYXTEtvm4nz56rduOVCEy0vqH4pmDrnF
lMoM5LDOWt8uI1idqDi7RhSCqaI1c/m5NhZL6wZRBcG3ann5odYbFKZk/iWRLZVT
4gCaNnzxg1ABkJT5lyM0XsDndzexecGVRj/5ytdYjUff4hU6VkThR4JjcMdgJ/xt
0lUzzH1yuRt51536M/LCFaIOYKdh3CRcEMGdq2nYpto9HnwTxkDKCVbkmMirn1Ww
rfr8HsoYtRgyUnwAu++ZnbakRfJY1Q3wXhBrMoLNTbCKwtZ6si4EtoURtukQ2+nb
zZEjlgaP2N3ka6Yw53+9tFd85WBPZ6l5nhOeDHtVBB+dNg/6+PP4zXa8sn/ABEeB
P6y+SdNEM/z0rKbOvaFEKaMQLm7Mg1E9CgRfCRvSRHIXwfO1KqRaAxKAwZjUrQKh
0bZ6UkcyEQgAR1xzDa6Hs6FDIBwD7Le87RFwFI2ZEcBvs4t/3hT6uc6T8PGveQSE
yofPlaVs39Z5IwQK3HeTTxRkHMMhGto36zrjk9e3IAyTwsqnIyoe6CgNgsScZTa4
OzeAhXS3WVCa2QpR+d/ck21W+Z/iqeFZEqfQqr6LVA3SOYwQvcVC8vlisbzpUq4V
9YrpQPVwwXc7ApGXqHg3+bNnKGr4KYDmGS3WOu956Doaxbq2zqhi7XSZK8HAveVQ
OD50Ixyb44PpWc54pnebotZZum3tVk5Hs7cSMifKsddE48If8jeebsLFTlQaIZGx
8KrTkEtdSSdvZI1v/26BnRNQxo2irruJEuItDUCxr0F4Yay1Pz7J46yfogWOHRCZ
5+axQcufkBzq6cSpP5Bggr6fyBqcJLpr39LdGIQDgxTUSR3eYG0Hj/PIDsz91XdR
7oPcj7xCIXSKgTSIvl+mtczeK7HhnOonrjPZq8jXKYmFETQikMdCW+HhHPEbmVS1
HWFvQ/JPsF/ipNGQjkeBf3nZY/Y/r/ERKnE6Sly5VFvDIgOCbq4Oa1J0x5npM6Pl
4Eu+kGhOjF2k7XUCoWVYeQD3r3BSb2gly/Vq/caUz7YBxQrLTp7Zga8gvDaoRKah
UxGyoIOgGpPFiSaQlUJV1kC+6s6HnAk9xSvxGMnH0WutHIoXs2qlOaVPWk3I1y1h
oWfD0zFGsW4vv1/TOBGguUWo5EgcgfrODi8Z0UKNexjgU7y84x3R/YZN+PJ2zFnq
afwjCLtD3f24bkkKJcDLtvbEOmzpGWwFL/6blcjbmDWSPfJZIL5sw+g73CrL3HWC
t/dAs0tIIyC7JVTQ77wIKcC3EI0o34TmEV4Ud94/v2SFffjI7aA61iyNewtKC4Lu
CyOrvEktymAwi5vm9GA8Y8Ev7iaZwU9WRDqXMkxSKdPEOU6YhpJu7bz6xNKnd2fY
bo8geldWp5/El0ikS3/TIoVs0bDJZ6QJ4lKxY8TTVTWh4P/62tKVw5ruYJXK39b6
F2/4yp/IEmufOrGLybt12XoAxbPJ/WDlNBPMpxMmhJHknIH/bogwTbCFYD9jYcJn
ccNBfDnY36XuXFYgOI12QrdjJwUZbkf4LUPUysAq9rl2ghEiTEbpSsNhRQBHPsVl
fP71wrCskjIR/3HriQAz2K2H6kcQIyKEq/SHhr3oiAtiT6IXvBRqQGlq3hQgl7rh
557+taGgtufj6HwqHZRGICyzRSO9D/NP//L2uojXWBVadnHAQYTjeyUMgCUuFbU2
hfWqhMo3nzDhNdaHstUvJ2C+mP7YEENweJY3m43cryuEnnfl69XPX+pHwrCb62U/
IIpnM07LsgC60gsQYeQM9KiD4Z/RfulHLo4mTdtXvL8U9a/m6jCOX6u6r9jxa2ft
67phVtMcwV9qvemQAyd7lsJ9Fk1WXhZvKeLooOfLNKw1u8m+QJauJyqqYVbcbU3j
el0pOxyBxAkKKUuBppGCs5ozlssZL/C8K1V/K3KsFioQGYEez3JK0xeu0eFIowzY
Z7kekSg3CTrcm3ONtMRSKPpHMeHSypsOXyENynAAKExmFbxEuFdbyCOxps9m+C6J
pg6vst9vZB9xCGOVsZE6rTcYIsPMVOuqSuP666bmPOLCsHLZV2zfts4taOcPbfJf
wmSdpHr+bML9VHyhsyQk7qtW6DuTEvJvPnMIXFvo5zRWzDl528DnBRmG/EeWY3uU
9rAR4F3NW9Ifn1plUtG8ZN3L9+nmqm1JM1qrq7KRPoFJUODcH7fE7fL0dWZWXwgM
1yrUJyaRkDY551VfnVcIt4lxblhkgVlpjeAvDzmkwZnc7nGI9FVI7zPN3ITlSCC+
bIfpZ8yF1QtmqI57HV/hP3tOTTpupAfX+zlolr6XFh4lkymvjCglx/6J+FNZCmYY
PTo8uC8ivKWlx/pjSkUS1cxXKMRz9v421ZmytFk1WVfcnsu3sQILc6WZiLHmC9FS
2Xb/tUgK4XLUBazLtSUicSDKrgEG2wSzxwvMw5GqxDqhkdudhiiXV1P/U+rOdpw0
wNKIQAER4iiA+P5PEQTeg5I6qEmGwksIRhMtzGdhJxeUigkasTMeQr1XhMALP8GA
O9qy1kvevvy9SB9hpusZnQ==
`protect END_PROTECTED
