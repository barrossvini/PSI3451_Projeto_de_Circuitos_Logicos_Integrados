`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F7tf+nH0pM9pNTuO429W9VLf5dzD2/rk/oCzrgc4gOTgeYZiGX9w2M84NtAG3GMp
zzTVpY1ey3L9Wiilu9xpgXEPRQw8agf9j5TQA5MFIqFr5g4D0zhJz6FfnXOprmWx
B6Cifdx0IQ9LQppGWIH84M2bYb5OsqgLayjdFCAJ4/c/ffM8zIjwI2wMNiUrTvDw
YhO5yBwApJMswTvHmnxQZHUaSrFDIjyHWpMRAGXiPPbDFbRX+1pWDRlO3rjge322
q0DDXVU+jVOqrT6wuXFvE6CXcIlw1KIizBWLqJG0zo6go0VVy+MyVwOzAyUEQMQi
N/rVwTAu6arVJa4OxW5woiJd2YHUrOxnV8QIvPyJAQQJjiNh78OM1KI4p+7x2ihW
1eDx8AiVCM/vLHOWS8nWHKG1ry+28zRvhtdo46QXkYH8RC+6QBk5ww2Z7yOX/C7y
W35uWghKPwAncSVPxQG+a0zQ6iasCYLqiyHuC9s9UdZyvKoNUP9s3liEVaHndqsr
BnhSCTmPi5JT6FvSgyICNdh+lP6qCKIeg5a0YeczxNHTFrXDjcwSmyWr1ETcQO2M
sq8c4Ompd4yikKS19fBBTkihDlUUGJrbsAseFITpkvid6e8ojEBU/XDdgtjfT7Z2
UZU4BcSvkN18cHGU38zh2SGPMOMUMuR2fv2roPH1RPBTFMRlaRe0QKDkonSJuhiW
FnPzwV7TUyuau63WcEq8P9BobLPRTj7L5FJ1dD2hbfTQDXNydpz6H1/kM0uHSxHM
tE0rfid5Wl+8kibXIqjqvsK6g2TQ/JHHRCBDBX1jSiBHZDr1TOJs0J7vcMcSCPPr
Ph9xEhM7SxtMT5hw+3E5PTTzZ+MHosZJMPWYbwZ4cHMEszuvjrLYmSEEypxvf97F
3hf+Uv3IQY8HqLPNHOoZKorsfN3ufzazIplb6w5ZKlzP/3oQqE5juDosxJhbYknQ
AHntyiQNcfLsB6foqlxDDP/ETjVDcVkmpLA16UVCOAzgIA8Z3i/1BGjjWm8HPeNq
jePGZCWKQHjvmMMIobcNePSDN5Cf/W8rJySkpQ9GRuPIMkXcbj8SkMCOx4Lpaxl9
KBxW8718a7+ikZnOi/hcQ13CpQqRzReFLoKmmNL+hH1BT5RmdDbbtejsmatxULod
62NyjX8jaCJg9dtGd3c3PPhptAtfQNsW/HFo4W+85SZDzZTEmw1yt5DFtzkrbTfh
k8OcxLnrVSIkM0dq0kv0dFc2iLYahvvF8bcn3g4eBZQci7qF+eHCreeoJZ4X0Ero
/Jxux2M9B8shmegAy9SD1m9obEAvD0ZAoZPD/A1wWg2IqWwXErkSwT7BuiqRrkS4
vHJ92rHPAPZpdXmv4RZGKP8/p9VOcx5YFO/qKGEPJJR9aeG0zi92yD9Zd+9g1yaM
W+MY/ZH50vNmWCKoraG3SRmVfENxcnmk9mo57XsWuDp1/WSTAaRidkJnZPIOTbAw
nGe+HsgJriyiGNuCK/t/stcR18p1mrcEdFWaZ3pEmq+0JEdCUfirlbNhMGu71zJ/
Sa2QupX0LOK94TpCjGIoAxISpoqR/xRsQbRYlxZHJXVDCb5UTr+xL4Sfy8fvPhWp
sD+z55dpujtf4FG1XNQ6uaZGF5AVtTc7KJSOCL556YyEZIKyVHnr7jDSWIrmx7d8
fQ3z0kPbLxtjmmZg8J4+NyOKAFB6fDzoEg0+61Wbl4nGifJLFje9NI0eHCfQjIVm
XMuUbNaLmVpooP/nr0MrZHwMklTv3ZJCTaQhY9ltkdGTr6B9sT4P0EktWJJmRm75
LBJupxtrDhyAzQgo+dQGRS+kTcS43kkC72oOH4A+qVrS6iZAKlz2Lry3g8DSjFdf
hEwfhiUt8aTEJXO0x2NnhOdj0OEkfDndy6EoZ4pPI9LHE/0UrahY3odTCi2hLSM8
tms7+uxW16B64WOLry6HXiWaDmtWgMXyaQW52DtBHSBccll8sQXKSxi6BicQaoXv
j+u1ic/tMCjm/55Q/3vaoV7cZHkydjhU9xwGysqrh7BRTFu31pSiEUWD2NVUw0CN
eYl+FcDt+odqdaTt4K95+85oheMN1QoFScrCoWg/ooLaJNNSHMxvrlQhRHi5HgyU
ToF0ukMkBbEAjbhV/Rv1D/qMW09HK8Ec0e8DkwUnyoY1KlfJCkiQMBQIWf09qRUF
zRiO1pq6qX3qt153DQS3VSFV6lE9JTz4xD51+rBE7CXgQDfYybSaE9QHmqCA6inV
B3rxjAZU42FgG6CUm7U8DZKxRfLvDw/UtUsPvuG9WCg8IPHZLgEtsiGHJ+gG3+so
cf9+s/j90tRXoFPS9wAqdJppPGoDXPDVnrS34lg0UpXfAwnMqFJbUHia1wpqnLNt
k8eknDPDdmDaqXJMJuy3eG9dcQCwHrfM+kAX0PSIp1X9pD3HcU7aVwqDVfr6pA67
+zvaD6F3j8JAtRDwh71s4c4D/+C6Ib8fS5fEwnXitxYa72dnwYl++YsM0Er1Sfbf
Nn60pkeZQXDZqD8UViOgJttwlQ11EVMcs4wPphd+sXvgKMTN3pTEM8P4Ryu4wSGy
x1/5APjWHtXwPyxBFqTSqUP+d9Zuh9qR4hModBxVW1S3uXJ/n5IcHEjXCtIxs1Uo
4TCbsoZFvTEocDIdry3tBiwLh4qcjROWVRAJJWHAgdCmMOrTQi4opEOYvKsqU+yy
EZm/PkEqfZqur08+9jufFJmozQ7GObuYpc20fixF6p7SNwFVeqhnFI1wPV6CmWCU
OlmGubzf7FKxuQtXopaxCSXfzpkZQ+IZKqVCEr5tfys1f94qo78YKoL/S7qSYebF
xPlcoAshskljecGol2jyO4u6M25YwF1v7HlyfnodZrVfjOO4mwkSidWpAVhAj2Dq
K3vBHEwsNnNSA4GwbtzmUu9Wo+ECxCPM+KNYx+X4tecPHcOZErLldxYzCnJNuaMu
6AoClsodzA8PWPJKDfbAr8vIAj052v5Y6urMV/rPjyD05r8GsS0Enc6XIFXTU1qH
nP+2cScgCegQLomgRzh8q9vayt5josEjga9kj6aRJuj2owNCTLVDuHyvbGwgZWtQ
rIWfiaNMevxlQDr6j2c7V2hhcoRVsKN9upGt7x6eT25ZvpCRU4dB2OENlwUt6XfF
/W3ar/Dn5mHQbU3YLRQVJtcPs0eEtTOjdBXWPzMblt2yKpYLdfjVAfkkN0R5ciqQ
/zriX41yf34lKWyBUwm36WewSZToI0o6bMA/ZHyT5VxNieIH3un7sGUfG7aZAfZk
0BAhrIj7sQK+efw/PBlmskp8ASQBxpWJqVEPdKu8y4TX0a+OyAEDvFXVtKNdSsUD
3tM8SlvSGxRHdEVQLseKLyHDwY56RS/sXyG8Y06H9/CIL1F5HGlg6OdWFiNtxSS9
p9R1ngmRtcGwBy35BHXLqyoZFwKeZd/7Qz9k7fKOg2K6mNYD6dH/KEDb8MW4ZESO
mdZULC7N78DlbkL5CBHIhnYixj1OIXClHotpwOczDHtrYDSW14WNJOLCB4YgqimY
8FRmETjkWaG2OnaizXNa5TSs6DdNvMu74d+BppEjQKQERPuKHoZPmJnHet5hPLMl
zGAtMa1/1pmCd3gLRgmVCKu9Ts64AL6Djw2wqs/b/c1uc+0YUaENCVGp81Wmz5/N
/38UyqRhCJWVqJpniKwi5Vs5tA75f3FxzKm5eZ0nNWF3WPAUjGS0Aoklbbp8COY4
xngXfgld4LF1J5ivmNng3JMoCtCaQ8EXyA5U6YHZMQ1dd4Z1tTLbB9q3qwdaRLg+
/wcHT7rZJyGKx1oJymw++dr7T8EmzNhSpKt6sJYbAR/SB0p8lVm5NqEkTgkM77et
WxSpBeQQ7YV4zBmeR1zXrAgB8j7zthvBj9i/V5byJ0E4QSLRNubuyZnBXshS8VCY
d1SAQydNAO/f8QsP/pzeopFurmL0PhqhEM2NH8F3F/wxS3uEJdfcBVCtR0SfBbvL
p9VRZg+wUop2jjUhoCGeidFLZsFrvDZGAVgR0AUPOiXHoRW4gFwlnKKPtG2TEvGM
+w/w80SAqDAg4alB7R+AAM/TrYoph6ZKUf8qontsPHijEUk4L7Xyfg/qH43Vuv/3
LbvERC0zabAFVU+vRDh+sifwxPvhhyhVv7lUi7oq/0Beif1JCmeBDSNIRw0HSvVd
uxKMo+aLh6RdR/Jxn1ku6kD9aNrxTv42MX4dUT3IjvomYcXxlxQxgYnl0ozKKX9f
CFymWL5Xfh+xFqcbybsqR58U/55C7IivGpzXU15JjqbbLJ1XtdGGMhVcmEBahecx
eXs1iUzmdhzd1G5LYH8HaoBQMTpx2F4It+g2hhmwcOXhOeE7y+dIc2oRk4sOTVea
hI2DDE+Ogd40VSdW56NwAaLQ/rxrALLDq5gY3tO50fuIKMBuHNlOkSTsYRqKGTqh
sY4qedGpNFFYSUgWc2gY0/YdsNHegPg82QQGuhYzLTEHh+yAZUo0wpkVdTZ7ZgF7
F0ws4f0fY5Zmh4S+GJ8BrNIMi9MA3pszH1q38SldQWzqnX6Nefm4X5HZLiXWlqgM
oHTDHNdeNXzcB2ugRiMc9PBlyi08wB3INSup3S8XjwGql5Dxr972r5eslwyDaabC
rwa2Yf42JtNa5UFaBj6/ECQ0FCxT/MxePxfCGbrMUhJWocS01Oppe5OA3bv+ZUXv
Jx+mB5WdI0wzySlckHF8UlGS2wgDLCtQSDrWjJermzEbB51QVFj2v0bb4dZMshIR
jg23ovCLGLz0rkhmwsXBW8R+sd2A/E/9xpnRYyEi43GObgGMigVbK2mDqvmrzHn/
dgNN9+VfpVrWD3sV21iDt+JOu+M977PrpUbz+gZbmOMD1jUVQUeFoukvCV2PJQpD
EDXHtIH6qraBVvDTETRR+qs106lNiPBhdAgLtcEmHcr/NFdfnrjHtl74ADVc4VYT
0ISCSabH/Uorr3iNFnp46iQCVr707ivY8FXVJT093pOxnxfcYx6DIN1Lr6rwEBFl
bCdMK0KROrzCw8MYDgsgyy823ooH1xVcwHXUlXihKlYLc5odKvNg3ykFs6Du/CYf
q2/KE1EpldP0yN/Z1SSjQVfQxRLm21tMMx7/5QLpn0B4lSkPODzf67GjhRf+JH21
uHdCLUGSMwBTCHLipQFRNQ8NICNxVcF1bT/P6yEzeofFGTjCsmtgEc+dTMMrRowZ
FezaHLXjSIdEkxd6QV59wU5o6Hu7gYRMDCJG0kfnLLadf2GDAddppMiYp3fdLrlK
zwBTTGORagVQMzYqoYYzGaWWa5rJa1+B+eWLf0YWzoWO5BI6ZcH1ebOF90qO46yb
JdkiDK4flSXhy9PoMzpkBtenMiqZ+Cpj92URre/NZdTDiVAP5X/vGGYN6t/dGLId
ZGqMRg4kSmKB8bgGvFFSLN9jqplwY1JPLxAxR6Yilg/SUvDYBbEm9C14O/bSjLya
YW216OCj8n4+NLKTD6cjnfYlF2lMQCePWGRQVh4avDuOWUXGLJhbWhpyjrCL6coZ
6xpPAgcFnMrYMdJFQNvXRQSEytZqOiNCZvEZX4KJu9X/ZOu9+ATcvEd7jZybQ3Bt
DiC0s34TqtBDD63q2BABb6LW1jbWlHZnk+wR5cYLm+sEyAPLJCz6vQnfJYhvbOwL
UUY31onWQVrVwGzJZuG5lPHLpzEquh2aQ2uIRPL0/r+DyWm0YeHNu1oZfsJqkn/J
XhHqG+fVSQ2dF/xrkhzV8657aljw33ohY/CQawQffVh40k6xzURaFo9QY2HKWBu5
v19UioWUTScx3sx6TcccBrV+3Crar6V5iwvPmPWeJKncwk6iY8Hlzt2EcL5NyV0y
XAwznRXK5Mb2oseJS39lAFrgtan+dGo0ha0pdY/bRikTAcd55hKUiVhl9swgYnNG
g/PdYWFg/bJb9NQboELJrYz2CGCOEHzRKoU6i91Wz3UDoTMg+MNKoygJGr84eaew
liIximU/Fuk13TEyjgdoMvXJbjKdDo6r8njI/W91PjwvQLg6O02m2G340izX6vUs
3AGJ3YwhB/NGQp+ceJAV2521Iwg0fuhdNW6+sDMEUUvCHncbikXfgQpGox070F95
z1/R4M1jCR2QQNZ1KKRE4c2YAsEShBNkAS01lyD1bQJ6Yd8qF4p/bq8Ih8T2DQy2
dHl9ytUnxkXmx0sMmD0zSE8SCsdTnzzBFbQodfIu3FNHZYDjoXRMYxJ93b1ooO2s
zyZJqsLKflskk9syv1H7yJJh0ES3rygdAWJIWgSzrHz4+jh8YpgMzXOXWvnJl47b
5ul1SmUfZ4doKnQMZLLHzpRS++YKUmzmhuo7szO4qgXNmgjl+Zp5z2+JJYGV3wYF
QBFy/D6pgF9TofYDt61knu89G8m4uaNJOXqRjWTbqfMy0FxUmgZKyTsw/DgPhLMD
jMjP4CjexrO5awQcFvn5fL0ifla4PDHJYT4fxo5D4A/GSsPjNwYSxYAXaH78xrCJ
dXxBXVKrEMulJW49W39uGZt6IslDSSyiE91Ex1YSzVxS8pjBHl0bfbawbHA2bUBv
D2A+s4/WInTt7XCWj3AJgC28DBjdQdheL88I3oVf9vhFVLK5lhKo/mpOGfOYy+aN
u6fpFfgiJCUXgwn/At38pgBi6C0ilHObocnpS5lSxYVDxTK5JSHvHulO2UPgzSWU
qjocCoYvlcY22Ee1uWVN5ngC4Ul38wYddU3r7hkKQWCQZIFu4rSK9bXokxPjuFKb
QJs0yENQI7HRvOh4NL51y3WZhYHpqZtlY6MegVeVKLmHaKMmfI6qpIa92dnm90o7
O3mzzh2V6pUBu9EgXMRgfjZFWwUCYS/QKRoImlQph0yeKx+GkpEZ23PtGdarJktC
XZyNUNrdwe4ya3rCRdNSyFHvs1Z/lGbMRiGSE/D4U1mGhxCKJDzekB/7n21oZh56
SBIVuFrykUjUo3YF7UpfxH+/CkH/BB8dpObQwin7QMz362gOftBBVX263tFrZq0H
8POuoTq+gcQWVvyhnMZpHmQ9Dvh0njn5DiaOuvSUh2uokjfqDJGphY2HsIOf/c4r
lXNHGdL5OGICTrl0i3HHdDeGIBMzHZYGfUZ491JaUFdy2mICeAJp99nb6wIkbIIp
ktcfuhTXSZO16HXwrnuPqRFDl6BM0t/QtTt0IRPKkRx3IAbLgPt6QoI4oHKiELzm
nkVCh7gWXLt7JVNscLQ14unEqsgTA4FzVh13S0a54i/dMSE4X9mXeOubP5WrmaZq
vItcXBuCPiPF8NbPFKnT/2DlOEZVLqmi+GzgkF/5/BqP9hvmNvOzEpYT5kjJByvd
7puLiHnl1iXoCVxc3MM94iQFNQ+Y6Bcdvsk1UVGn0Z+4MxqZeYoCs9H0re/xhUTx
/3A8lvDAe0eRf0bXMxq27nlWQGx3xSiWZNHe+4RH57tkfeyjgoAq/QXhdvnMbrLD
Qi1a/7/EzJbn937RHrErNRn2q6Jgy6Rhd5D4zEyLhiKLqHudNHqIKYwAMYGEKcgT
B7p9MuPqG0vXcVxSGJxn+sg/X29X8j4A5ZO9baqHwoMT5vHKUnj3HZWtv70tYIuk
KMgZAOSDmVogKKwK1UTu+Zk/J61a4N4pXjdXSg8E85/RYlzOLEmPl07Fi1wLLz6z
aG2yEgJA0wVdR9vNLLagzaxXNeog3hvBiPhJ8/GO0jw0D++iwzWP6kVa21GXCIeu
A65PYrH6qrQjRFicvxLDYe8kywtcldgEF12+c338O2QASVtgS4E3lpfKTadTpW1l
6k95Vd73supPmjW7uxgO0lP9emKpoEOc6l7ju7JhqhOPO5EtZ1ytaVjjk0sjRNGg
mhwD3YGQt7QpbHyJhYSgl1eXN10pf6E3tm4bfk0JGNqA5pDp38YWMjaZ5Y/26Xzk
vL0bcgWZbilDzBtpPVq2/1H5GggiTB5hLr4CxngOX73cPFYq1qwMof/h8/XJv5JT
5+lekZOXqNy6m4OcSAG5FCaceg9cdPE/uxSyflt/7cfp2RtHmzc1piK3U4etaNUP
H+JuV9FaCsCx+bEJIisiEjtHIPNDTYqiH7cLCBhEjMqcg7Y3TB8PoD783i85qefa
ax+uuYoD+ywOkcoLfc0xUbf0ynfYU9UNfsJkhltdZg6fWkqXUcve5pTymOHh5Dgz
XlhNthr4erg/pLP/sgD+UR8xEOvESGhgniBuiLlD+4QC/Mb/HDywlYqc1lzrKkjK
JVNFPQh9qJhpt+bbM0QPW8peJNzVwfppGElXJtqiIdiGtd6DbaXzNGfZGHh5rBKB
PDmjD7eQjo8vITz/RDW6UvXlFDEDgTAZhYNvFv0PxytC+o2Td7kLxaq6Fu5ygAts
eJZ1SWu/I2EKoNoi/SHAwyiJ1cVkPXgUm4Le4fsiqB84TDuVt6y3NWRxXb2rbpzv
Wpc5kkWNAdyFeYxk0GiM+PU+Yru3eTqh20FWZARInzyjrfwAl+nax2sK5JpzNAMB
SY/m5b9fnPVgdEgWx5mL1QImakWSL/whssRz5ai7w9CHpjxJaLW2AspXss032eU7
N+5mCstyT0gad2TC61HMo2xQ7YtWEykwiUuU9282D8wxqQmEbY6eV0ihTq220VI4
5wxfcyMTJl+6IrENv20uudK9pkzVNvwccWUpjvx18v/35GxpXTyzFxy51CqRqPsf
H52vCdxSF0H+eJStPNtA+6filLdUI9UJhxy9iVRoh7Q2MiEtdukN/831sobpkjHO
jzXV7USbKnrIaXYu4mZjj51aOE35/ZTeXt46SQLMcguGL2KRxPeMePPEnaslM1kW
c4rbsaPjdx/zRTDxEBSAcc/bX6HxB6js242ZAWd74eKU2vkO6YoWLI1MaASLaGke
aRGfPwCOH5nAGebHs5++8gFpzn//eLbbk5ae4bjwno08dExkF91IJj9hvCwlu8Xf
CyU3O2z+ek7EBx08wII8OrViR9e8g1Serpq113SFQlkLLNrQrZNXEVuviLGLXsi9
+nJ2QvwXbD77McrkKdWBDsNyt+2+PxPHPeCFg7Y374yOLn9+u/kIPLALQz2PiQEA
BjKGQMnA7l7TZuIjcit1sS3S/uulCInJBDZXAoBeBa0AcFdsRUG9N7FoGcWwZpRI
bEUd6NLQx4eXCvcscXlhjb7GWDn9wR93xD+RcqSeZOo21tmgOGLah67b06G+6Wrc
OdWKC5LLBI9DNbhxrPQ9BVgY7D6wrjI5tjMwCSiM5ruAFAbwGtbirISip6T2dPES
lkW8dX92D8/ui3y+49LfSbJH7h+IuZSYVTWW9LpGcLE99tOsTsgVnjw/K5aSg4+2
MJ4fqRmHh/Bc0p9kHUqziyBYZLd8d9UVUXpnJHH3FzVQBSfHJD0eePTcWZ+u9bjM
HhSKxDBUOqX23yFnywNZAfipXzREagKGIEK3cjAIEK+Wo1UbGzm8TUHL7/d6+ATx
JYQOhl4wcu2BywA4WxWCts6JtQYzI+uG9c7jl85uJz/7dQPXg5lgH1rGPmek+VFc
16K4+ehu1JSGkrMsRKjdt6/1t/Umk4o8GQslAOW+5T9kHm0wQM4Vsz1+j5J/QbdU
ut3AZ/j4Bh/75JqED1MfOjjOOljg+hVw0/4Pdcl7OXzW1qYdjRiGgPeJpCjwpb5Q
gzffoAxPcawtPlHkxs9zwfBdFyIZNSN+PO24WH209J+ikhfVZv9yrPy6mErJ134q
xeIj5sU60T6az8t29xut3y7M5o8vManWSYDcUuOYj+hnyrzP4Im229gvXIuUevug
7GlCKx11qpJ0CGhTzD0Ua11T8sTCm39RY2ZuCFzZS7dvxKoWOXnIXvdEu9xFIWuA
pXZODBNobwsMdpNNcLNUi5onuP+JysaDCVz9zoeApuXkl17XBdc7x3XswFdA8yjJ
dk0PyvS2ELJLjcVx46ZBxdg249H1IzOS9RrGRXxhzJYmNtnGmYtxHNEHMMqkBjfx
pyWrbsXAF1T1bHBdZdbKW8Shx+azPqZn7wpbCJUlCaD0SSB6bNNFx8CI72ayxrhN
X4ynEQl/vVwF0NH7RxMyEXyfVlvWMZsBfo80javiIJfPcRyvY3WCs8axhdiqhKZW
NSuzwSGsY2t5qUBUBDtOaE4ZX5fWBvOpZ+2xtGxuCddvShJMkeEqR/f9LVvJejlu
i6+vTM8fV4c+y1x8bW7iM7Om35WavYDuf1SBn+yLwjWcxrA3DzV/kghgtG4MZLE7
Xvz+qcBX9ARThKwZ4lD8TIIC4gme/kw13QbPq0b1VNnJ1jPPDuDXFhppNOrbuNpV
BTTDFTV96LXiL1Tj1iPJIR33bEao9VSKzRE16IUnRIJuDFOtnr53LkZC4WIbrAsS
e7akhOl7oWEkpuRF4co31/qE+yObBLKUaP4rF4Ke6SKLVACGyubRxQq0R7wBaNMu
yXKXDE1G3YaH3DL8UsHC5m6duZKNaMm42oEaTt1t06vtRqj2oAqvhafvCv4qbEQ9
1XAf+FXJOWBxkoWTs4uJlRWTnkEkwADzNXn2yxRvtn1yGsdBkrsRvobz2z0lTWUh
3E+6lw2licB1fM3qRrmGf2nGPkNhcRPNvy1P4J6t0Za+0pQLvMSVwSve9AEKstC9
CCbW3rz70aqAOm+k8WkXm0Lm2djstUJMc9UAmlFBhHbDqbJ5psPp/nXmeDKl+5kj
HO/0tt7zVPrCXMY/q4RVJbGFQWKySnWJ9NMd89gsIWn5VSC6U6u8EFQKmulPABH6
vMCRVux3zI6vZkmM3DLQRru85N20l3OzWRU/Wq0uPQSaFcwE7p0TLdJ0htmLyXbH
Khk/Cktqd8xiueZifBKXDqzcSJWxvE8z9EvM8ywm4P4U/TKHjv+9TALjYhrDyXK8
hBXDNGBtRKWKmE2rJwz2AJad9eugxsHL3YlJ9S+LAnZmDY5qckPrlQtUOehJxUOU
kAeo6iNj6KdxINa1ZnY7z0xMr0BjjMWtKWG3zhEkBRjVrAQBvI8wmzUXMoi2VpFr
7AHXKkYb5Lo2dG5hDjO/7EfvBgPXW8ZP7hKEl15qkILzdaMqNl3YK897xyUSbviX
rzYGVSuwrrvhvPDbF4dLD6rFYAOcaClI0h4/Q0iuplcDQCsoJkumbRvyJepBQTF9
9BR0HiP7pZHeIh6CgMWaKqTDrZFcwfDvmflubnqvJYyYYSesEKjVUaKnQbGJe9dT
VxzKd5EP4hD5DXgQJJthqGbqJAQhUZE9jI+t18T0R+l49mGumcjM1f8F5fYT8m80
/6x8+axWEIlJiGErA3FU6tvZtmGD3trhA3wWWQikbsp07/xIRJLJT1agN9PPn767
JWfMOFSa+ZEp/l5YsXkUD36FhmFaw5+aXs2/sfizbdjfkVz7o/8CQH52vVR5GPJY
5AOJPnRE+8TgrYP9Am54AY+oQMR/aXlmsSgXMUlLPDXAx89eLgOSbhyXD6U8ORQ4
od/KXJAwNF0i/Ycmd0RIK2L9CvB/gFt0a+6BLtPcaDzyIe5u7MXDbxzD6B6h3d0q
hxAenlFUPzsAdYDh1aCmdqcOH1WkxPS2qMsStgCsebNQgehW+s4xqbCCT0mBB4f5
2Fy51oPJRFw0RgMU6sFkg9e1hwxddrKLdGCAt15UPb7YD+cdwpWvgkfkH/3zt2OR
HhZgfhXyl43KDQU6iNvIiwYPS3hvvPhccBxPX7oK+XDuj+LahClcN/Sw8Ng9lor1
R8YBB26j9eu6KInoXD9GqxMmMKYq+5jZU0AtNotGjkhSlcASiaaGEqTeArYiH+6d
eEw23Ac/Tay+kTCTxNN+DATE4yqd2tadw78Lwe3vjL5Tjl8OcUbi6DfnBC9pBXLC
AtBG/ANj5RASA7kpRffTUjy8bowd0zO+L6pg1a9EtFhLw1O2YA7NPxDwRRpiCanv
hR13lkuWWOGeSZf58lL6tN4Hdto+mFw20JX0Sfm0HrH1ORdKtBRWubXL8wFqYSYg
4Nmu4aq3uKZcACZAUVwuOV04YNlGM70ukFxnKli8xzasQ3+QnVevl7uFTIkuoCOX
TaLSi5nHAjN6V/mqpPuo7CKPAObQad8JeI64Tkp4JuxxWcA2R+cKpKMgrJ1Btimq
usluQpkBa1ATdIM4Ty98BVKJb0dV8b8vxSb4p+bhFBo9FFBtgA8IwK+wiN7+ZW1I
JkjxtrbvkjxMxOF3Aq6miKjMgBVRrsqAprsZqYSxzLfmpJQgzg2Z19lgIht/WFtl
Z32PT21uty4caHEj4XtG/IYUWLSTHsqKe7zcaKW155l+JwOtoTPk5SNQd6ZutdBd
GZ4OIMDKTikknT0n7jg2Peaax+J6YnB9PEPdDtrhcuz2DqH/KSJU9Xvl9TXtJZxq
qnYL8I+KRIAyUzB8A9QkUHuS9qh9Z7BUPr9r9hPNx3an46TjkTVuoHpUnnREKsWk
70A8l0VnZ56nDt/8/UNCp5b1Bth3AWKIsw9+AuOSfspFOBrbTxKXTzEYVjOlDi/8
bYKUU8VrAlsMdf9M8r0Jt0gzxxY8tvPPna7Z1igIMcAaTmsdps85vNMblzlez8UE
b4fOXIsNkXRLfXudUBAus4otRE8UXXOd7dAMztUdJCWl5aJFmL8l+rC4Zu7sNVxM
dmw2oDEhTEbQr8ErQ5cG5Z6ZCWpJWTQUZxVx7Pmd7Mzd/MA9qT5744EoEn9NvohD
0/9WHXZmS93Qw084QvavpyuLhyePry6BuRdhtqzYyV/Vl787Ain5BSedTVp/mX9t
etOKEgHspjNhrIfhPT/TXmirrwFsPItA0La2e098PhkvE7flLKMPcsoB5mvSzuaC
u1dOca7qHoFRrxKsvgd2OJLUZuqLW6Wiku/jSSoxQT69ekFmTwgx04/VSXA0h9by
cop6jVuz6XHcmh80h5bfKN9+Wd30XEYiMqkX/VSIj+d2C+YDF2EcuHLdUYF+sVM2
E5sJp8kTD+k6ZjmLxAwQeztzJLHhvLhqQQ2AXnQWIvNetbqdVD3uSc5mxc6tCoCC
KdGDCwqcw8FX9rqiWEzDrV1dMIQ0oQvt86S8109araChRlYdb+9Uuy7jez+OSzIo
1yNQPdM2KfYJa3ia8xeKgwcgSjhCQZtUNV0z0+TTTbBNOBigWVQboch0RW+vAENZ
Na1a3bDnRYH6ksnH/gqhBR/JDK9pXz5e45nYNx9wt0k6uXKrUybt8bq8YiaBvsiS
HgVukyTsu91HBbcrKOqpGbZYTG923wExPbaW2xji1frgUWFiZYfQ2TkLV9femEet
SrWPEzvgHClN+UIX4Nl5SnUPznlCUZ5VnIBUWfBJn0xdyXjOqXvEoPdLbf+BTaix
3xXIlmBJ+NtAJ+VpMInk2DW8O6iNskHxdTithvVCyCUtCQirqjRBJhGOJi5aFqwm
ZLyr1DEat/zXeSvmQile7khhIBLUzi+5N6r5e/H4At6lt3MI7Errt6Ol7tzXEXos
L97lmBskz1Y1YG4Ya2N52hqR1ZnfuKxOTglETYyEHkz02eMv5LQn5llapipg62nb
C0Ti0sLD80P50p3ZoKeljZdk0BnR7TRNLV1KLg9aqf/U74utjw+4VJ9ECBr1TU2N
OAf0nGnmIOxeXdFyrcrifChCx+raIgwTU3+AUb1XZ+22uvPoCjuW0pfldZYxtpdK
LkL3Yz/kCjBFZD432WRq81n//dPRbW4l2cjyAnouRdfnsgYyLFOdrKdx00JO0HsZ
jnlrGz+8SpGTkCuk8OcTJ78AxUq8v7OeoTeiVTuYAgNNFaSlbO7C11t3JEu3u0x4
mo/v8/jge6fU3daCARhaw7i55Etvl+vnWJ78jAgECYIZEhQsV3gPrLTN5Lolc4V7
mRsGB/49rmAi20rN/Mi3Xhi30nr2+DHiufg8pdYZNlD5OlFiVsbm6sfX1GFYiyoT
4YrW1UtfooEHsvfVb+JmNLrAufXqPFOpM2syJsMAjyNwu6UXD+xWPBkRgvsPD1lL
biQ/0UjzyE5YLlfNwj/s7QmO9vo88AM9ATn4XDp1yVzAhdCdXgLMDtynk9W7qX/E
6zzOYrk1su0sp9/2ROQHgQ/9Ib7z0ap8eWLGV0oZ6Hw9aPLB1wF15fVA+h//6rLy
e14Tv3N8DL+Z3SqTYZKFe3OrP06xO5hrtKHHFRUH+/XaaZHCmfgivJQ7lnJ+TVce
tEzubA3Ngr4FD/stgSgigU6phbz+ZiK09wipbXhhwBll6H97cVU/3KnBvJ2/fGLu
LMbl0Kpl+VfVu2BsxZFNZnUmZ62H2efFTq5KJnzxqun12nMUn1arYe1x1+dB+K4i
5UiJZD/H0ghp6n/pkRyi4EEGCbvDn+gac0DPLtRy6WvtgHBSkaJBRYHzi9gbW3y8
BlyWNFqzgnB94qhpvouYiPSbSpD01QkxuCNCY3xxQjkSZAeaQmt5BnWwQUyf15cQ
6OOWko32LwcFNQh/FlNZTMPoMfPvDyP4UPzJ87Z2Z0aX5TXkaK9DJ5gM5AAYyIvy
rD/r0nhlXX3qonx5DQqkH9MeyX+fMRcWWcQ8oqAxHedYExVBVqVml/OTrTNnGCsn
JPFSB86/kZxHk8gtmJO7ZfrXzmQnNrKKht94YxfSyCatFQwNLITzxrLxplIEux37
+oKzZHeENMaYKWea5o4LuHUalvIsCqqXiPlZday4WTgrOvTzgFupI219RkmtdWSM
1As8lYSbUUIJTcOAo3Vi8RZHLozmm24omm44gv9PV+1AdqHkSjlBRdn9zoRe5veX
DT0KgDYal4Ch9SCmUMGwsGxtmMFzt0LLPVFoh/16c4Wm8SwAuGHZDQHb/RXhNh7s
TS2xDJHGRiGkh+WRzx69L+GHmyimAzyC87NguzJX9hzg00ndI9HReMa+swCECsjZ
eCt/WIMgOvimQXoxxhQIBsZc15Kgg693yjGEsRRE6aiwbAXhZRAih+IzjyB2rabp
7udaD9Hubg2LEqzgn5uEhke53//G5/X6bRgIVo8KvBAE8xtsHhtl2suAwb93nd17
VuYVGAneQI+fOvmFHr9FiI+F0BsytBDONmuvsmwTt+dRVNzLHSb3aHJTKtwRypMo
MBy+U7sl+H9Il1hcPzCWe8G3LON7cV0LQrCs9WvTNcYIn77TZ1zwIxw/kHobwFc3
aksnRMiMcBcYUZ32tmqXGnyYW9EmaCIQrytHoQA7MepIpG524hdxxaQY41IXYf/R
TyymVaoE8SgxBa5/Da7aPHk0NqqtmYzg+BJmKa/m13IQOtepU2kNv6W1T/Q6NkLt
aGYwtExxLR3B6W7U1hVQziaSgLMuQAdkNHGL/lWfjtRxQoyQyDJTU5iIurMYMFgJ
Tm6clbaJGQFLnqp1uiAtdY6P+KfKxx00srwnpYDVZEVj2+yN8R78/pEpLLW4Wc+M
aFCcqWabn3+GSB3LneITs9RiI1hVhCdSzVSqgrl5SKkyuMRxblK37fUfqe79Lmj0
oqJs4Sbab2PePgGfZzU50ziuwlFGvb6VYfyiFVvYbyh7IyvNjQARjEBBk9SQwfvv
q7e0BhJQ/8xxODc1tcqA3orogQC/xsNkdD1pa7SLdrgcmI0cpIpPD6msHhZ8WYJp
x8MkcTptRgQFiCQaTdYhHUKgjpdMG8TsSRx5BEk0CED3ijvh4lr4xWUpoGwkrW/l
AVpq5G90PpjFxPLZOaXu40qUmKNWJGrwfX9sFRF2ITOy/dPjQV112Ic6iQRucGTt
7E9TmLTtrc2UvzOVsoQwULFTisYndRvdDdaoajSx+7sM/DBEfHRHSkfst7hMKor7
w1EDpY3LKr2AXiDfhucoKd2Tv2VUF9F8L1r8xawzCusqvR+URLxwNUrXaukj4dFM
hyUyQNY1G4OZki5EYuiNKBCOhqwrXRlknj8w8eIDZpco8ibNKyZc0eaJxWolC6fv
AV0j9ZXeagopNo1NHmV4e77u+n5+bmSIoxzuW5giKN6chD4Cjm1cyOTHpm0yP2f+
kj3lX4EEsiCWU7CgX9Vzlvnxl9m+bq7CNms21TI9fBW0X+tjvK2W+cD6UZ4J4E2L
3WHUWwMxIAkXB5ZswQIJqIcTH7QStu48oniEscV2zQ0ohZBEi5XzCNCT8j+YWV3l
Rxd3MGyOGnrT7miSZXffLhgbGicLNnDKHXKHQf+I8lIhVXlEkO/KFdLq+lFTEOBd
00D0/G6n4Kjqp/AZROcPP7NDAak0d0N2xEbeQ8CqnHdTAtyIu+mb7hZ9x1STfnDE
j4kWyGitfFTw5MlyXWwAn7AdQsugtCk/SS7VDnEjtXrPR7o1KvclSXLcnMgKs1ad
uL1JvZMQszlDynYpiRXXZ5XHr73n7Jtn31MyVNohTwKHLzdQEp0Ut/7oE0YOZuSQ
D5DDkQX4561G86xept01k6yjHhlSDkfSSvUbL0/X3eW1T/Vr7WXfFNr1k3RGg/vt
Cd0mHyMmJfdU4ndtBX3YJongZT0j7nYs3wFSSPiodvgsYxEJNQ0ZeUjvo9iXDesA
QI+8Y5u0sGNsG/c1APWNB9ZjU4sP3Y2LFi4gPaFLpputAQyZyhQTof96iXnHWO2w
+VG2FiidCLP7kzto78Hnm/T5ZvlhKzKyZP5WvvX6j7RDKbYPHpSflzkE368BGF7X
tBnykNZudj0LyXTRA+4y5giUTCruoVtKYSsY1d2hQ1zMpjBrneXz5WubeZdW/qq2
hBpV8vqhYuUTWat360d4zLxtGkdnrlVCCQiTqKqRz06NGxHRZAgcwM7Kbfwz5jAS
UFbXDwDnGmKfmR2ZrYfijLflsEJuFf5S2Uf5soxrZ+UEFSS0v+fDDUECkGuB2t8D
TyL/B9E9X1nH9P60HlNR+p5JHA589BqZMJ6Spfm2qilQlDC/m1jiNxuBJTmVi5JJ
aGA0c2j/1KWgysJt7bB9yTkWLz0/yQNij1gtByVLLsHX0n/j6yX0r2rCNR4vZYFc
UgbXqPbu0Gfa0vo6HZxw0riGWZNGt17yLQJ/EyZDXzadRxT9ap1meDZhVP/RPGsK
DxhwVuYOF4pL5Z3sy+Insbre0NBAL/BuZUqCPSEZgTdtTDEwNUyUWvkwiWFMYRk8
I9VG5MNbYvp9y8egCbYyM3J5ZC08AKx1y+x+kDmRri+2FaLvjcGWp4ivFCguv3fM
VqQtzAnk/beMMc6AD1MX0VsftPYyl4m/SyMbUg7XhzrBe3g+aZT+exxFIDJL/KwG
/zij4NPIAbpMBn2P64kmEtVLHPKrD8mR3DO6qFL9p2F9C6G1N0RdyNlUK5bPv2Ta
wEkhjkz94gb3rPPs+k14CpUpvgVmfrk3/psa1wX+Q4RF4pTUlaNCqoeGef1HYxz6
8Mf3PmqoBTxW0CKbLuRKqGrP1s6ymOFEteJWlUAA48lXn3Okiw/9TNY8d8ILwNyG
PnzcFwE5edpfTiRUqxsEzQSTmLTDf66dYxHWeqIAh9nqJiWLw3/4qN7hg3QASYJN
lT5i7UREckwVy5zuiK5DzvjQQ+mgcjV0+LMRmJN/Ig7FdtlflJe7Oz8s0Y8xtjTj
b6qaxs95yg4L7LMsQpvYXn079s1rl+S+9L8ctOhJz+eBHq7B3VauNcXRonzwzL9O
HB/VQodgqg0/XpV9dx4r5lGOaZzJLM84i63Yg2+uh/qXT0/77GsPpTNWN6GCOyXM
2t07T/YUqkUgFtDRb9yIq767cdJYiTmDqWN6bf5OskBE3WrpQ50KYO/dZm86kwvC
Oc2djjQoh/9Da1aYXNeXz9VMg1cUCkl/YXTd2AwncKlC/Toy1nOoG7o4+MOdPSas
NQxbJX3t5eoXnPU+47cyNG7HSue8jdpxI2cblFaJ0xHVDcayNlBV7dRCwoorQxWS
JWIDtnPY4pcNLVlzrjQg/9BNEtGW6WiXmnJ+h2/vtRwNz/EtKRN/14ZgwE5AKikX
rWdQVXWdWmb6875nplUGvwyItORewoSEKrA0AH3ZgFWgmVgmFcPmp+DUcrudvup0
0DnxtwxKxh/uTvsj8/SQKZVtRaLz+R5W5cR7ga7iu7jNZCthR0if1OsvEtNZ0aLA
xVn5NIreYk31zVKdSyZmtM3pFJKRZpkMf9INqFM1DWShTLHF04Niv6njiulP94bm
eGHNr6LEhR2iDrKXsTcAxkuEhBtJSUKzI0SbAZKV0YRzaLql40l3CRYox7/teg8G
nAqzpLITk6VNZwo8ZxrSmx3OWc/1ziqCP+gvAAs2JPSkCwUdGFhtLT6VXkrRa8ZF
Oyo9sMoWaPDWCAAzAsLUZsbCAzaj4DgmhbmKZwQMKmiqdzLX6WNCz0U6TNqcVjT+
PQ3qdwCzc5mC2rtET3fktx3VYvPqDnZhun0ireeqdoptCXhCfvxsF8qWgAu7Jo1f
yOb4GdvsbowVsBNvoMQt7z4HtiDN7qPbjzdJf94F9g9FFSyiPUvyuhKxsmjBsbWx
M5qOgO6sLFROyhRZibZ3XT2TV4iYZzQii1RXXsd0hRQQoyJF10xaHdNHCzHazLnX
TbR6fauebtgG+BixnvTKd1S8FyGi2EPLL7h/nah193wycJMKeU0HaTXefrvZ+LZg
VlFWaH85EoqFfftH9k59uTQS6B5pZdIZQsqTOsj/UuJvdlcVds3g5Av1xgUWoJSz
6QAfQ6KJlXVnIMkS+eAOKI3TZreX8x/tVFQVHXoj0uUgrEb2ZgMbzNkuN/Cdpj6H
xgcKisa3bUfhT9B1z/Ip5vpgnFPcI4ZKsgQ+74lPTp1po60EqfVnmEGUr10DVFA4
72J5X4cYfWv328LYivAHdM8QUjujAVf2ce3L/320V88I+hJWxjRP3A3zoPsIYrKC
j7nlq3QCmCXU+BC7dHsA4nuG0DmQqsAL3eMNrkokc8a/hK+yPNM1ehZNakhJ/A0L
NQlLLwyZ4dr3AjlOu1MNO5osy2JcSwmEfKVbUOA6eWknFj41rJpW677dJai5MJM2
mdd0uB/Y14LAXCTDXv3RkJZW/BhdwdDQ+NccKQWnYreUxEmNCxv78kLjCVV0+YJq
uu6njyVfbhJ4XHXl4ysvI0zbFHJqmBrPKIMQwNE0vf/vB0wLSRcX938tHNE9Myq9
kcxNN1HQPLamW5rPAy2vgYW64kiLaaMbcsVuD+3zQ011gBG6Tfm4QwwRyGAy2VzF
QXLTlaAOdkmxwNoJX0GVM6OURKLxXG+2ydkqT0C8YyNtDdGx/fbwDdcMdX7eFtTQ
G41s7AE6RxNHWBYAuiIY+wzSRPjDhL/be5s8EyFPlBN3F2yob5R9q/RbOBmqp8o7
jb4gAAFfxOPooKoq4chgtg/8KQiM8FjkoOse+kgikUnnPFPciwXXonMnKUyMKGoA
wzZWfuOU2ztfu43zBYMw/U73f4ocS9suWLS44Tldl/uuhfoc81KcgVp/NmS9pxB8
di30m7sXdKEqX9MsMDxPcfh4PJris6Ukx2hP1ReLBc7CVBfzFO2enrZ59C4UoxlV
D1BUBbmkB+l5WZf0Byh4VTUD4by4dWhXWFplO3tMctNuiw9BHZ0ictraJs19pJg8
4gPBzS12Q0InK3Gpce4DeeowF8LZsTlChRQbkQLEQHZnXPIFDNNZ2S3SeMczbf5I
9+t0QCRVH/256gKEt186ddBslzTxigGVAsnLBd2zThrWzEfsUsvEYF08WZCqmMKB
2y6q6opbZ23pzzAJnHiVBko3/2CaDnGhPHqKRwu/83WZnQEPz48MRwjKKBJGwb4i
UhhxzeW1M2AdhCSSn7wprlO6XcZ6cRrZ10eIXkgp10cvd8yIxHl8ggdae2GEpZbY
hLRJNv7HPuXPlQexvY2FAY09VMb3JLKpxPxhJuguvs7NhuSmYENP3RVMk1sa71bB
qP1NTX/EUwGx44IUc8G/ETNDmffsXVjVX3h4uZKcv71PA2MxWK7bXPu/AtvzDlwE
Xn3Z+U9S3stE2ZvdckeRe7L7TF2ugoQggBsa2hV3uCuC+BWYkPJ17O+os9bHPFvY
V5BNNxIxKqt2huPQUpfETZHjZfNh8kNlNApgJ6wK/ahPTq3YKf4as1SBBZa4+Hb2
jrLYDqap9yP97JPq7TEhL/MHNQ3d9Z+c6Q79W20OpfPviOtKzvISEv/z/HH2pcT0
nUK4hpCPDIIuWuGnMQtl7TL16oqWkxPF+T2HT728cgB9CaVWtdH56yYRirzgHqqT
nG6bEbeD9un7b3UbY8Z4NZi/4H6on8rN9VeZg4fZ98ZT3ZyBPa6DsyQ06U8d8s8L
157NoNz9ZfWjKGk2/NC5zq4QJ1xZpwFk8XKVOQiaVhTYziIXiAGCCYw7N5iq6dzv
+BYhI11VGd3svc4Ek+NL3u24bh5myib8lKXRpwGRIZXMULNRFXZETFwDf0+j/iFn
EZBQah20ImZA3E7Nt88/sg15MhK5/qGWw3fAa7S02x1DM1/eczea4MsaZUpaX/ft
Lr9xNmy0QGL8TKAulfBihNfY/jSFjl9Ap2xXZArBYpSqpP9TQ9zOwnr1iosoZBiv
TEXejUX/0uMcAtDPAqx1pEzjrsD6LfyP0Dzb/TZATNl6HiRZ1Y5fj8XCxceBrc4V
uUpr7csm+XfGYogHZHSXpqLpNO1kO4ob5NM1kzqqp1ML2PoAXwWaVGghrvLTReUv
kAZoeRpKnTgTkCj0cBE48+ImlRHDI5Qu0Xzc+TlC0vGj+g96qkbtRhP0bVUvc2iW
5q/qBHLqn6/HeC0nm7kB9VPz4rXEG0wCgfBOfTM5WIsmnc218DjUAftZ2VGa5lJG
U5U0Nqi9Jn3b3OT0iWKYtFtiPsZeIhz0sMOCqv0+a7UAo1Bqq2G3MLmoPPGF+aWY
+DpcEKOQlHWXcgNSo72+icuHt/utSVexVBmas/aHZ9Zf8sGULrw93AxJEBQK3r0l
wsPy+mLQyHxLvgp/HFkbZqdbH+WYbaydHBIw1LllGZ24eW573JOZMHILLiRrQDFy
XRhIpROnWyymwL1It5SQI3MvfCYjfV1dxZYlRM/AmVAq1muJK8vW2lolPnABsOzA
7SzyT3YEdHzts+1juIg4aAQ3g7rTedbTwMrnydByv/14uOOYJiouni4lMX2CLZzb
b/CPVfh9sXB4vZ1UrnBAIrlKwj42x/asT/2JqyTmNqTtQnjZatmSVZ5357QHZkqv
e7zOrbwL0Ltjqlc6j2gNMNs6eHj0IH/euXsM5a3XO/4FAYw/uuCQMBOpqmwQ5FLd
Rz05FZOjcFqzqn7+25scx6sjN8Rx6elJoSIsuQTZRgDiOPj5PlTgQ8wLdvP3PUpr
iJ9E4zWywAJct84JjcJJkBJ9Qzy3yfJBcwpSFqjDD+Fb6BH3LuDGUwquJtojpsUB
I7rfeaBdZMp5eGbHGa2qer3bGvunVbJ2eUWEv0n7xnw2hhq1ptuMYBC8k5eZnGxC
RNcRvqZP4zXNsptfAD8FrwrTg4eV0cx3FJrR2CailcU0a0n2H+GjenQpZeRKqDZY
vCVMUBWihGGaiL0M+4mKZ4DChXT6VvU4XbktzSfmWHL7np3YSqgO+IRKOOS+8Lgn
QgMIzShoF/S455ms7O1sXhL7wwPFdE+9y+JzqqPUSv2Xqc7ISbl+Qwlvp0MUVKcm
qgBVuJeOZIG3O5Wb8mEgjKRciznGqByG9Fw+WWiyL6GFhc8Y5P36WN6/Ih56S4GW
exF0cwcMhugUahRorvmw4bpwhIq+oN2UkvRNfiYQ+hLrfKQzz4YUNU9pIBA4l/fv
edbIMlrwbU3JBk8+rb58vM3zdTEUGh8D6mu29kHaApQ9jsXVZtoXgZCzPpnOp25H
mrKSnac3NdmwWiDwwgvNedcY/8HbDTlFAHLUonmPW6ooGoweRZgdcCuI7kfCtyXM
/NHMb94vgoCnbc+PCUyf2bMTUt9R1clM1lBs+pu2Rk7Nd8/F0laXGH6K9MT6ecvf
lz7xQ11Jrk0lPfzgrCp6poIrJw8PhmhEyiEGLOEdnGBOcEMjzQ5qffFVaPSkTmF2
Z7VcMs8aHFsHm+AdfzQPuNXSn7AmRuy4Pc6a/tKKCy4NI9av4Ewl/GOXO0SV75AJ
RqBeTqCJlRL+MNG/BCGJW1KryQ5697ZfiRXi8AUrkH3z7AiijHcyAotMKIyAbGYq
mcZz6FDyR4Cfe0f7//3ylUCvvvHxqo5HfB9IQDWEk6u7CPISTzmoAuZ/eOWQuwlh
jR88r2o1jDGVfbEvm/cgTRJtyJ9qM+6aqyvd1AcC8jJ2E9HD8OhlftIGmKSeqBEf
vxTErTBl1MS8u0OlDy+wr/CPW+uIT9tZgg+F5MWCpcFpc0A3yOv5PyB4aXYVt2GU
aLbXfHqCZhbSOUk/ntiZwYXt7RBZ3oWiJC1kOaYkqcizKMMr5oXyjYhiHWpqJ9z/
c/+0zGXtMJhhld360dc8K3lVSitGEh6elpx2UsetexQX0mQv6Ya1/MnpV6DvmzRw
FhxqEPrqWq4jU7ly4Rs0TnHtczQYnPIILnzyXmXcTPXGkZm9MVHtPvxBBkxf1chx
cdV43XIx3YyJfsArM6arN5FQmtTGZTQmt09wz7aLLTGO1ewh+sXUMsguyebXMRws
2wME76KbzK436+EOfF3uSyZ2mmlQWHUFBr8cgojbL2wgX+z/LFiNqHlKATozjJ2V
vwS6vEZF/fSock937lxv66FkOPw4o2o/nMuAQSjcJR49XyZYFrsU+4Mz3Pj2ywO1
ddvmoQV64+OHMyPOg5JQIRhszQZ87myzHx0HeRfqp+GKb5rcEMddeF86Ecl9gaFz
8JRb9njqfCAImXiADTSJY/m1evwvScNHgqCJCHECTFcL9nykrWLz3HMnyBLhf1a2
aAHad0VprYboSNfHK18LY7IRdQY+rP1rSUbs6zzvIaYNYAL+Kgt9sSb/JDVBRNdK
cQpNvlpPipBORUwSBZg6EbD7ixGuXq/7GlO7AuV2YNItfx6/G++GI1wL3XVk+/LN
8osxf89wU0uwtXsV091rP2avx3eElaG10jj3lmcvqRS71IRCUHlBT5GRDoAt7T3l
d8dZAXB7QnyawrpIn/WR2pIqr+W5TR/LhMe3hMBtP9jswja6kHdm6/fRu2onotlf
hipWv5u86/+3/BlIxpHUr45DCEea8lqnPIGoXGiO1Di+Dr6IRcZmZgro368NV5GO
N1ybv85XFNOptNBD1HCMqzbyNMagJrbHzk0sIf6hhqEq82+40vyWk9Y3JZ9oqUq2
Ek9GqA9MBEzXZnrlXEIM9lNZ7ImAemlRwru9CMPLUH4MrkJwbjDRPXk+I+VI+w2S
JEUfIGCYofXoZqQHMDOiWevPiK4BEAM1vdwCODcENuBPdbHSkSsjrr4Te2mxUNgM
7wYWMeDNOC3IB+1p6noj+pD10z1Wnr9Xp9+hjiuYwSmHYldUiWynnc/uviUwN6zH
Fi4rlGwhvOEIpW9RKXef3ou5VYfOKeJUOMdUtDspp8bn8hPIM5b7UXVaniRpGUv4
VhmnIlpi9UQbNiAtmNC8zgJOUdE4T9C0MrZUcZkWf1lYk1v93zsqhU+4pMBaVaPS
SBFoA1O0Uc1rbwDCQzkkF1vyBkUNFXKPVqtrkzAmfQv0apc8VtD2pvWiBpsXvm9K
YTpbb+BeGPZfOkTKskv5BYKm6thFMakgZTeMilGoIIUpzAVdLp09N7wscSr3HuTg
n8uThBRkvmJQ6Jw+7BLHMFpMlSGdMyhiHy8c6VjuCFiQDUTSu47jgacImjdMf+Dq
RNI6zG5Q5pD/Dmx0GRJ4QA8vdDeDjRe5Dtrz1F89Z5m53KTQzrMxf6lpi2uxcSgX
opi+1uLxPYCGuvoSs2aN15d1pS4nuWlVkcpiBc6/7el0B1M9f4Dkmrlz6aguGnQj
DS5vXCTU7ATqFkB6WoWTV5EF1qJdDd+vXNInyskQiHDGgpo51B7xv1IRLvUc5KcC
fSJKaFXvNBZ2t2MhNqoJncjwkZujOa5qHgSiVIzVDBrf7WjxKisCs058UFdL3EGn
wvde3JhLvWaZqnxI0qJ+8wMPPAmfl8/xurx4I+3Wj3C4cMgA0QxJs1So3NpzlvsO
ubLAFsYo9OZNZ+wg9lmujelnqu1MU4I9Kc1sJKPN+yw5VnxxgVC3FCsMuAAX3q1h
KnI1S6ecuXPT4SZPK4NJjI1dksg2obD7CsHxWKk+Q3LiL312HQHWmLMgS0dfrx2Z
WMMaDHkWluEHK7CVtszjaAlntU/tQ0dR/qyGp8z9lQn4s4gnKVd68fbenYkrdoih
ij82zNqR98dr9AIG0fhTcJWEAtYoXTR3Tr6yz8+FBrYZ3asXC3blTD080wMp4SFr
KVkP5dGxGJdhwaxB6ZW7FULbZUsa03fc9M5tLpMvcyyTTHeCFe3QVFQkA48+LJmZ
g9wp00S044Ud8IoRpAi1lrPo24B/uObqWRHh4hqQmzQtweYb1qHBXg8exDTPEJNT
lmFwD7r1bFBR9Z4TGgC+GEUSOjGTIwkRO2EifbJObSxG6s8pgLDX1tVjgoiC9e3N
zOa3pi4yHxNdXY4SRDUzIyPLo9TT+CsqIK2o0CFuj0fvDSxARtAvlZ/30DlVGC95
3M0hU57Ebn97kinpEyXKkMHDhtZ+1zONao24XIl+hXcpZdcoNddCpum4dNz96iDf
Ymtw7l7vStjxSZHbBIinZ3U9re3CazH8m4EBVWW/syE8sc+JziuVukixn/qIx2RX
u6fzDzEsdD3fc2MqJ2IxI9eP1rbiMKNaXasSbFLcdgziW+xNCN8IZv+3q7YTuL8z
e94mEXwqKwUtVvcxgbpx8AnP9gT0FlbesQAGOS1kZLmNLBfofn/eupPGqAEAPR9K
UXE1bvYVDdUQHpxuYq4wH4MbxINjuCYS/1MIW7o4HIS0gMfJVY4c4npQw8eJ/EKi
cjrvRwEXRJOulfzNQzwUUfZNFUx8ENxGVF/xa2xLTh1PyLHtzKzmDT5cNOZibUWf
RGKb7KyexeWk6q6gsMTlVlemRXZ+BWEQH6G3FwyF2s/faAuYBpK0FbOANSN7skLJ
mrdsXL/BkwT2FeOi44UF3qcLKZyDxqx6hHaYnnyjtmzLG/EWcH9b2+xRJdbJ8yGS
7BtH9JFxORB/GjWhO2f7FBO9obulTo2O65ODZahQReTS7opoi3TNjg4ulR2/YdF3
sonvcFCwYWSG2ZDO3DSMZfoJiWuEvoU0bk5BLVuunRmscsnknVQ5adiPw3ZjwlsI
yn2/c2Tt9GdBSpm3SeTaZTgethVSwveV0X7DHqZA1Ok7YBGwEHz+SamEsHh4/snx
MEdJUkSJPpooUoEIFh0D+OX9j5jyRYOyJP1s1W7dgO20g2/FbYoMsP0y6im7FHl4
W3Iqa0ZWfqHfW59l+BeEOKcNdnijRfp0y6qV7B0Clw/qtgx1pgq6WhLYrn+LGeAV
OlC+mgU412p0aiQJXRlUtQWgg6UiLTWo0D8owF7IXP92VtsY0nrwknGJ43LTqTn0
VD7Me+OD0S8+xaeMM0QfNNQF84ln59tG1slgE/eyWqYApO+lxXppDdP9dVMjPC2l
eNiOGPjrOaOM+GIOI4u/DacF0K9BinPgDbbWRnaO7iRXzEwUDEvutkLyO1k4D7UR
caEVsKyk8Q3ggV+EGOe1E415kSPpMZhRxvpBItbRcFXkBcnb6B1wI+hc0ECxwd4+
82oRChBVf0bxVYy8sqtNCMoma+hS9XxswV0gn/fVyryVmXCq/i/wRv93gTpsn+p1
nKzPFO+KWxvS7vBA2SOASg/0168PEOABb71oss5tnVwiMnCprRNekop7qrq/ey+L
GZajXvKIkaHfuSp3BB5wq3/Sub+sdScl+X5xwH/SkCyiSzUf99MjdUzvdOAHYUxx
JfrWuW1Pcv/gKvydXp1uSEQQ/YFfISBfCz9XsC4z9p/M0ExYOKZtRooCjoFWCZAV
QEv/7KbVcO4nHEpbiXtJfY9IaMs9kilePnSpymZqgsbJyhZcgHGgGlx1rujv0AO/
MgfeAtawnr1zQ5382gYgPsYHMh0v0XwKon6gGmGIHr4+svBGzeugTXpWZQ86OzpI
RlanOa8xt/Z5mj3asAYTAViXgMnhaeqXV7ctLB+c+Y6ubzL7kJHmIvei6MKE4BSE
MyfoD5jvAB+7xn8HDV62vR+elVgoqR0wi+h9YKjk83ewvyAgN3swqb6v5JZwO6cT
1mUFymej/nwbGBoOd7aOKI/i5edrjGwtt47PaEeQUAfo9o3NYphLI5zvR1N02nbJ
BtbXMuiitHTMteHFk/JiUtdcFP6CkTg7lNSV2BmjIz3qJE+QxdwvWfzQeLOkShx4
xMt1iIdtN7DUDOL3qmYQTv7D2KB0eIfe0zLbKnurnIz9rjdqhsCAUfK3PoOYCk18
Hw4nA0MQd3uttG3StsoCLHjASvhRz0yWxfmdl7yZvd4lNYS2UTvTUe+jv8r7FNb4
XtvjDzi0N7B8o9TyBc9b4d4hfeez9a8YUnN6sXM1T+UyIPhgsygE9IbnPyuebAq0
b/W9VT+o8tNElnTKOrprv4/KaS5LCxYTz3qzOdNOtur9imVutpIaFRoyjOpcFY3Z
KxnRufE9/T0bz83LwbK/Home882qCTMe+pThR78kImSVzPAQ2jgiIrXm4yPjxZV7
o/v+KiQnYp6uljN58IpKam9Xfx8BltJ2uHIatGAPO248zxUMopfvAxzfPMUQ56Nu
UU0VsIGlEu/5vwfFfzYZiBFsM8Z/5Sm5FEsLrTPGks0/ZNtrcHQBuxf1Y9Lb3Kk8
5MXo625v6M0NF880ioIWy23jZXnYC6/ggHofRuHYKmJ00InW9Apq025OTWRn4lWQ
Mb19H4DOiVHX7hCFKrLhzQdXwS3fRxjGOIqbpR011y6RUHOkoYRyt9LmcdkisFxp
fSRX1aIQxRpXJ2p40GuY2+w057p87wtLtw4IK/fOiZYcMFZBRXTfIEpUdgyN+SGR
uMGPMeeUfrivD2nzBSifvJatf2FSBIkLJC+gzsZRWMnxZwYyMJQoO96iM9bHt12+
YizqezMXyKLZIy2yhLCcHZ3NpmLVArl+megGCarEoaxAZmN726xPUXBreUt9m7Mt
yzxjx3KBx9OryRq62dxaGSf+9PDkF1beDU7Xe24upUePKoxRvvo6uWscdujz2QZv
QdtvFMLdZTMdQGbWu5KVmZWu338IP5a6tL0/aZ7WLOeIb5/aZveOZFEwRFwVPHci
HNYYprWx0tWvg6qutKGH3Gx1klF50nC04qgCU89XMqEpLipvU4PUPgUhNCANMHTs
6U+ccCZ/ylzmDnsIxFx6znJmjjaQf6b+b2kJZ2EMhmtcDouBoxknhuaSpc50xaBG
BIMzWt1ymkGF9g2iFCdU/KU8oQxF0601isCJg/rP+zUEYCyLXh/dGUwPsr41KKQt
Ykwu5f2WxjLM/+dshc4Yy5fnUbiq7t77uZ9cmJFUZ9a47AqEIdtTuNnB70sNd0La
CmWpQiwIs8lieyYW9d7WfuqjOBVfLKZbZ9LRTn9jriRrN4HePw5TNgjl/hrxvma9
lDPw6Ijzb9Cs04v8k6jvI/zv9kgL8BosXH6j6+kYdsGvwlGxwY7YuFZ5PC8tBUMv
Ekcz2RcRVB5UiGwroPR/sAZ/sXjrLcUB5YewuA+cP5VOAvIsiMgZm9qtRSR5tero
nddGaOEorahD8P8z+ael/vq5PgeXzGflP1TWOPzhyEcUuEW+mJmHYCAZ2ffVkzGQ
xAebQhGqKNVmRT6/XLx4apYWLxB17IWIXj08MVb4WVuTfaJq6AdWx1NS6wuCcjQG
r9/57vgGD5zAt9k1z4Qhcf09gEqjyPaa1vhi7j3RhuUsZAbILLPOU16qdzQDIYHp
R6tIjHooex3pNU7GClLTe4Jc/NKs0Gm+wr14O9RLTk7u8t4M5C/tIkg97lVTaPzb
ZsryKGsS7S3k/fztk3olKXkgGIm4E1jI6jhub4tIaT+dLjpevXeN3sieFMZxZGCd
rFRLJQS5SB57obEj6bC96ncScxSAuUL3irs3DnpaeNyZnNzMQ2EHfFgMVy3Ci1sk
qrV0hB0mF7Fk50wKY81podt8npDGjxTlQNbL7+CPW8HcM/fqxngO9b4UFZePKSU5
rlHXjDPGqoGjijNtuhPoeTTiUqEIBcxYqQg2AZLU1oVpp/d5br4kCx7QJq/eM2SH
FUYn9z3IuJmJA+cL1BWZ5N4qykirNfVS+qf1qO7bcYF25Ioz7pRpkXdmGmq/Wnol
CnnRhg6cN4+yxgtDZC12bkoS6m83Qb+As+IAyNYafk/7VNSMs5YZPYgAF5HWZRqJ
jXs+QqZj8nBIVYTIHcewjR/HQVnsnwjxg3jah3jYZQGVEiLwNAjXpXD2pN9AkOkv
OyR2VwZTQ7aTOScNjY+mOOpWSVj9n6jnpnhld5IATwEW7B2Adk4Cjbn/PMhaAybO
2vg9XgzN6C6nX85tPQxRUlFkHgtG9aJKOvFm3Pz9QV6JHn98AtjVNzMNWiFny4PY
a8Uuahd2YoJPG4eFimITjrzek1U/+ydEZtFvPJ8V+IC3Q5VnYO+mL0gi3BILijUE
epM3uP8LwbVGm/i1fJkFiG9TSBX/EsukHYO0gtR/Kl7c+20bSLarEL1DE822E9xZ
zWOFKP1TQCm/ojHzYVHOclnzN6OUVKN0V1BZqTo8GyZ6s9O3kQ6RHo8k3iIu/WCt
R4dlUs1x+w7is4wn1oPFizjHDXyowEgC9oLh6+3yB7H8eoA8yzBrV3R5QA+ujE0a
nHSKBj3iblXHExR492dWnkokRpWlD1VwV/HA+k5w+H8UoJ2x8W3QIKyKlabT5I8t
VPhsdfLOXI2u824PoG5O41NsgeCilXhkTHiARRZgKvKDdBvJn9fgPXlOtnONUh6p
jXhNMfB8RrrlV4SzKaSPu1Nc3YPbY0yJHp+YFHDdg+t3A03i6saIAKZuEx9d9BxM
FpW9SE3TfPHe6qrAQYUVl6mG99Pp7eb31Ed0DL4Ri18TPByJtPXPzVnr5YtyUoaD
QzZQTVA++rqnd4qRUeE4m4zcdTlqyTy6a/55h3HDV7Hcz43AKbMCxu3Fp0camhxI
MTIZKFvyBQu7U2SXs24yFQiLr3SbUQ2CtZkM6h6ie/vvWX4NK2e/Emc++bspxmG1
4nHZl6IhBi+l00aEuPnZC3xkvADMmqdYvJXwthfobJq+4wlmkQcOjcHcV+lExU7u
cEwghLv7poKuYVS61QS2aEMCOR+FQAFdCoad9xida+bM6UoO9teqBd2JeqHb9OuF
2t3GDitSr0vLIWBqmGvlzhyjg9S0yj3vk4pkWFvjdZaP/KgDoTp40Xds5Z0B4mJg
dilvhiZp3egtxfyN6OjiHsLFoX8s41lWGOyRD2T3sNlUwW6mHtBaGjWno1vMpTMM
qrWfR5dOM2wH3ZBPW0Lzpbg5S5cgkSL5Y2mRtzU4TT3aSuzXmAjpBx93xc7IZ91z
MizaZcpEloMqOY+b5K3tIWKwghD6UTylYaccp2M5G1FHqI8eznnSHJRc/W2z0/fh
E26sa9hK6UXRzDEikd2MOB1Wu4g/mawkXbSlQvo2e4ZuyL5P6vKcLR7Lnvn1vDIx
W0gXSPEHZE1cZWPoi+oqNOQHenyBRepnL8LC+iD6ivYpvIkmw1v0AgndNQmzDpAD
H3YSmJD07rJLH67BqDK2i+Znd0aMcz4fGYFpOHxG2Y/o6wYSeVQZEDn9H98FVXUJ
7azbIKozLwnKVctBntUZj//1QpwvYurIhl36ctCvquuE7fWD/CeCiyPEBEL8N8ni
OdvNFpdVo6Hw8ThK45reX1Ol3XkIoXwgmlAOAwFL7OegiKodYTuZfeljbS6krOnn
5W+5zhv271df1RQKVmvdqh9H4tfLF5TnTN4Yodtz3RpDKfu6yNwktBit2+2sv5N0
P2RJi9YWsuDOnGVFfLu9pHEZC2tsX2IHC7FwCqimbMnPdX6DjsnQ2VfL654WXtVW
HFGarPpe6apGCDbK8VoXXMIvtwEUr/mm+xCkPof6nyrCzM/QOBwt4J9CKodw7YUK
R+nwG7FdnqqRuOrNLiaQAgRa6wHgxtA+5nW12L1s0hIB+V+7cPUN0xVOPgyVLo2z
n/nW5fdZn1VYILz6mVN9hHrpoWO7b0REbuzJtWP0NiSP9US9GBTNxMPyOfK7UhCz
79lS1YBwYMV4WoA9zbnwskzYP58+c+sw1EmJ1/A22yH4DaxhpOux4uFimNmPmeRB
NNDmbrhR1t2VPZ3Tf1MBzXjQtWdM+wL2hH4fqwYIDqwh2NQOsd1Gg/DCl4JTqkSj
W4/NnaM/Hrv6XiuvpAe6IDtrg7TacNX35SzOeSSmYL80C8/aoAc1ScMBZL2NjoJr
6XLGlWDkDitAJ6Lr7tGG2fjKvTKnF1q2gG9AVcfwkG2qsPHkIjWdQ374u7mOYo0f
yUKL4bj7wRRj4nUfnZpJypZ+qinBf5h4fQ0cXi82PXgZrQ+m4kVxmsIdI1NUL3BL
U/xprhSBRgSR9wCD2Aml+8318ld4LOU6+ybqOXDwCWtiLxZcJtIIk4RdlI+85K8v
VrmR7JNYsl/z8ZsTOHAbEi4izSj9jpBiRSEwDZ6jRvpotc57RiqBIPU6W8VmpsF3
QhJPFMjv9fjVG2iCXAqgXVOu1wsbrL63qqImZwaSICSHtNykaR80aAUnvZPWSiRl
QcMP9rKcSK4ndxnfAQBxdx2/KG40zd5/MighxbkjG9EJcaHZvm2wUQo1hEoOF7hJ
aLhbTTiafjhGw3gb+wPgoRzn+lUZ+98v7vUYsS9h5ly9gckRlJ78yqdTs0ghBmz3
1/SfMNCNc7unKd3+SkkXXsMvvo8vVc0/IOL2OQawZmXdJu/HJH9G4FkHZxyemS5y
0PGdUqx0ELz3xTGTOeaqsntBlUNFdyH8iqn3Jq+XkDEIMipoBLV+9oPk8QqKdP93
bFNa9bMkvXpVEnwWrTy3/701hb2LdQp2CY5NGNo2/T5bAjurtSa6tIfkYMEyL6wi
7Vr62S5o/r+dH1QYOwfOTimLpt/oV+WJ/qU6orLzmatHW8s5zorc4hO6FVkxf+eh
3WQHgj0HXgxnhZBjbXITg0s3W8FRo4CtVFPVC96jtAFDzfQIZKWd+Dkabg/oIptT
lKxO74stgS9nbFdpYioXKXJi6LrSyBieLQrIgOHn931oFeoIYTg0g2ko6aCu9R3P
7TvxvaKRnZuWJN/W1cwEZRMey3IfseqLjQfP7FPTI3Fh9pOG3/ACf+APeYycRM+/
rUAALEs8/bbTXX4+9sC8Bk7w0b5QGu/N0rtx7Pp0XM5SOvLxmgLPcKB7d2+8Sy/C
9UIjzPxHfWmJ9AHwSM1JqAu/j03sVZO9XYAq7T3/WkoWP5bmDMm3JmXx0qORlvas
ylc9cv/cD6CQUkbaiP4lQ9hdrfl0icynmllJKq63rgD8PzLiSWawCO+XTToRiRaI
s2MM4qeqhudBlvpjSSxxdB2dMWCCGcR06pDXEPunG4lF1cIaFs4QtlqqRK2sBFzr
V/RwU3l7+tuDq6bCR7bx7OARJOEGO4ITVZ/O5pmHrfDmIyLnCqbJyQ+VK8OH1X1I
tVXF6aNZt8YEaZ7pFKHISwgoVlSpraudDuF/4pInsT8qK93lfhytTjfD3OnOesB3
GU/7uT9bilonjaHyfeZQ5E6sUz7qCOmbSmbhPu8mmswV/L+vwpLnQ6XgjYV+2Tdl
wVw1jHXvbH0eoN900RShN6D9c/xGt5+ue2igVWlmejNx/plEbNLmfJ2ZmxW5+f1z
p8t8OnhaPIO5uVhvyhGf2YKZ7b+cs+e9xEn8IPikdws7J7A8e6MbkPLHQjAJCaA0
h6zAXREYgSj16+/V1sCoVDWN7ToYgUXuo81LjiJ0qdZz+CoCiS03U7J5/hy8AYBs
N0CJYFJ+JCHbWq4GE4/cTaWkWVG/apeASjTuOLtdzmR+AhOTI+7P1YNHxoO+aqa2
lHDg2+/jkHvJasOXD96/Jzt7rAietYhCfoi4Zmq8gvt2o7eSDCXdi2PkY/VR4kMQ
dE6P0LN7UgfbSnMRrPajH34NB3iPIirUKaz0u8XTYpZnGyGOC+++fsjSJEsYiuu8
ZfRkxNFMes4nrTdlN/SAbp8oT/urHpzVaGVjDdy4oQZpxuCFIl798+nWSBfKO9uw
SpF9OofKMtyfmNOV1ANWShACD30TtYDTV8/h00fViKQqiVxCXc08nWvQjO/Ol2AT
huDyJm0vqIZv1ErOOAZpMlONICggKy/J6yuV6QVRNoEexLO/iVZz0aq/Eq9McssJ
De7AqeUj4cPfcEm593bpavpu2hTZxsiqi/2FogT6i8VUIJk56s4wkrLEUrQIB7gl
lhQLpO7H9eI2CRqqGygo7LTcwruiwwjy3IEs5FyGOcxJBfML0yCB3M/ELYf+ijcR
kKbJSzYICdMctoZM95kMwEzM6FDq2b722wzvljjUhAhEGqaxacjG2vO/lZGkLvfp
GOyyKAGbmCWUAzt2hZwoM/zXddHtvtwUIVd6LHpWbh1R3ximriYkdeQLxNfLVzHW
FyzpEV+FC48yOP82KwN/YF4e1xDHufoaE98+sFAE06OGHDcMvXFGmPu0df+rN1HA
SFmCfp7bh930mh2VRDr4SY29WiFqDvC/AHFbs9LjKyXn7fE2YjOGfsxQLq1f5NUx
/zwDGw5YejSqTg79MBM1EP6ybqpkE/l/olic4RTw9qTbwm+Dtk0yrb7o/3LxQwXd
KcukxGtaWb+t4eZxLfSbCWeBPGxlkN8WxIiG10WnxK5RswBiKx6/9DcExTzBTqoA
NUIH4YZp+55Q0D/VuXDlNymEvhtBlOqxeEH4lH0acQnIAgmdxVtZOFQxxR944342
6qn/EiNO/mP0EoQqwfacnVZ5+9MIXB5kpFunIERrl3/kuDhmMdxHftdC94EQyRb4
AgZzeWcX3y2MY1PDTkzolvhptfO9xVn0q5Xbm2f+SY6TROPfKu06IJOVTbYgAr87
Xmhd4ZpsVBJ1SrfUIUxuWMPAaohDgRLx+aFRe4QO+wmMjQLB/cKSSSRerm4i6kE5
i8LnvgwPgc8qrsBlkMHYlGVTBAGbidg48eXsVNbbk4MKXYpbKoUTtyLId97J6958
WyhVEkHE9hTB9NEnoUPok4azzwdsUm6jG0kfND55d0aqEhNFchpX5q36DI6xpVro
MvpyJyopB32WS51d5KZl7hLNkbLRColuo7ZnNHq+lgIBJyya/uoji4KoqrSMICye
BjaSs9XfjVccX6v8g2EZpiWZgZvmxH7g3i/4Pn+BzAkZ/4DzoNwGh5xypuDKgYy+
0NklqS3PBJgWGkze1puC0HX8X5SCX08ZZBObEpjAPKgYzrGwhvHcuF9B86BpRePE
G+1jXucoYmSg1NEN4B8EHMj8SWctSUAmqm22pFSUQnKErPMy8o/z9VAGU6bX6WYP
S263iJMZp10WYJ+a+QowHTgeFhr5Rd+XYo2jlT4Iv1JwizSoLvGa5Xkd0MT1wT/P
xG4yL3Zm3+MEd9Z1w2TCfmkDnfeP7NsXN+Fv0PqVse/DXa1yr+fGTsbnqSxr0xuC
pJXdC3CFPzIWjJ8f3awLQ62uR6Z696AUjVtzJuXFNh/RPVdnVPy66LGUUnvyvzLg
W6ZRqj1DXha6eB1KQ43BqVzDzSCBav6GaAGYG+gH45iNQS1+s06Gto5x3IopeB5q
LTK99SJVW7MR5DAGB+eYLUxG/hrUN7HxaFCtIyZs3X1mTIBKx9xF10JpMejJbBlJ
LujU4joo5toCW1eK7/hO93FgGzufokZ4YMOP5qe3kN5n91w6aN+uVScjcFilbIGD
oiy183iK3uvdxuLQ0jlfLAS7Y2ARSM73TjjAt2fDSoFNY1i2xkPXstuyqhFFN3Dl
JjHJGBZCEd8Q+k5m3NyVqe29O/RnQ9L4tJkPieansa7cjYuYJNTvhrjUjeABIY/j
jG9v5EK8g8eVcohcEjWYuLs35bQEkDqJmxRL6LXmxBVHQ1vdvNFCcgTXCK0Mv7D+
oREpb6e9PWFBOJtrp+koDVdVqvrEIO1kjTY0SABlqJknoxtoIyrJltptSK9O1HG6
Wz8ZTssJq5C8mmgkYc3CojaLX6P+qwWL5sYB5Hj5Pr8HDB/d4YLHaqj84MyR++Mq
K78YoQYcAS2ERcDLJvR8+Tv1jdCKDV6D/KbzfJ2WO5teJaxsV1jHY3B2vhDmIG1v
R+7DEoF0T2wW1ZzDkEL4OzajdKJyulE7uuQq+Avn6S+Dkp/P4WerFzOsJivcKkTG
uo9rGXYqiVAqeBuy8leOJefV9ez54qqIromneQl/WRMmBp8K0bW9ThHeAkT0XpoO
1rVrNI5WF4GpZyvnx9Q1jv36r589BFoZsZfFguLtCQNO7gUNNTYhQfGL48NF8Qov
2zmKdUoj38dmoe0Bf6mmFnNs1X7f/O5X7hNxd7Knm+X1T4Mx7K6Jq0Y4v4dfb2hi
e4gcEzdGtSeb9B84Hqk0VMP9WEHnqobshEx1E8DVCUZF+x+nwgIDh5TG7s6rU00U
RwSJ8e1EeYquMNSKSwf0EAeuSUsLDgcGrr1Kz3Q+G1dHqUA5at99LPn7XKB9YtWV
gaD4vsAoyuG1T3TcxrXg+4VeZx3Do4vCaH5eVOw3yT7tdjlznIreqBarVYcCxduf
t1ZA+imdHmRKdvxW/HbmwRuOQKywA9JDOybZ4zr5SVV1YbB+RuqFod4I7uPp4lSy
0aaNWXTOWSJrmacINhEeE2BSXrufOiFSZuWTc4unylE5f1a+LRo83Ro1+4r+x6rp
lfT+1RvrFARVsVWEuGrPkgecXXjSUupJxLEM6otmGA9A4QYnHFcJXVr++q3I9FnV
jCA95GnCtiUlL/3N9ihigmYGk7a8jlD9tarbH89Ca8IDRAhpyhq2T1XfpGyL9mUd
7a/7K9Jiyhl2y3HkiNF3ty0mXAZn9RGXLMYWGLbmwREuywYLVT3N/1e48i1zmrOs
QLRe4V0hXTLWbgIkVZ6h8DxlhEQPnaNMZE5y2xv20Fc36x6fo8LGCiCS5E50nDmm
Ixa2ZsYgNAR9BDt1rL5e3qVAHooG7EuqHIbWi2BiM6mPIcuKCMhsCnlTzJPQti5m
JrfqH6JAePHhCSlYX88EGKW8/6IU6OB51oqw8ON9rokBtwSknRM0OUiSWccOiw+s
pggdqoVC3u6nxCrAKadAwS+xEBLsS39VnEyW/b7EK+fsE5QgExe00oi33zoSqv7J
izUsgySV2a2QOysO6n5+ISm0ijaW2TKGm5AprrOlQq7hk2KtQBq2LE8q+SrQOJxc
EVXOlHEOZm7YHsQHXEkw6oxZnpMn/+cyEn/I+6Rb4MZVLffRIi2I5mMRP4n7Mpgr
4JbLmEEE7UhuPTgBVns9qoIobRuBNgC1Hn9UJlV2HxjxW1fgG1O5Ov4/7CbBxttf
HHlRDbOXqB+1USJJBIu2AGGjhmT73sVE7UhfpcCngzVapEaLcnU8WjN8w3p0ykus
fZIIhWrkcls5wADV8btRTRiFa1JZdNYTsO0LXPmSmOBIIbv36qyvpwvvU8JN/OKC
zdQPhlc/w5spDg9YrJMAMOeM8HtyPOiyPPaSDovNnjNgbXOXiPo8e8JLNYpLE4JS
9DJYRcAdpaBAKJhlKOZ6LPDNMjps1Mv4WnLO5/b2cZxW3RtNpaMecOIUu9DI6gJ9
W4D9OpNamCgiLeCJ65lyZxluvIEF4SmXFxnLiMlSQSjTQFB4bjEHLbKZwBEXHrJT
fL2ZdOLxFDnIuxxiNcQxo75jbyDNFokVwXSGF5p/2t4dTxDdiRx23NICP+6peKAP
nPsVSTB0DHlP4bDYLuAUA/hhw0TKkuwFMjy6TP5K4lo4pRz+LBZ/6oShuAKmkQVI
sp8AuPba3dOEDZD6x+V7V9kXOvAMEgnQEv96QpVATy81jID9aOPWUdHzRVr12Qmh
buDKVpH2WUsemJKnG+j1dpasBHJMcqupXnxbBXdANlvwxR0/EZ8BeN4jLGo/a1Xk
RvBrTXy2DTq+pS8h2TJZCZUz3f6BK+NKt8n52DJj+ksqa6vs0xqqUTcdXEnWGUR+
xDDSaLrhbNwW9vnA+PVfxa29ADY4HSeDNpvzlEX7uZMQmDhDN/ErLi914icFtvKX
iX9kZxz1NGv/lw/3FnAk+oteTLOCm/8Nb/OVSJvgi5UVn3go9XeAxJauk8VqmnAG
cVS24dHR8p2Lv0Q+iRp7Y1LFQ6muD/A+qMUHrFCntJTTq+4bS65HxnDNiBPqLHmI
NrWx2zlKlqkP9s9HgGi11aZpnkCOM1h08elNpndoMZbZ2K0Dpx/0aDEosAvLg0yK
twhnEdP/WbHYrjfaaQvWwY18hwTaquHG/1VTCGc/4IibOK2a3Qrttz7ja/0vmPtU
hePVovHMWTQJK0t29TJh5hH1OTmBDRkCRh5cOhqxA9rTkN+KepPGCJNKYd0Kp4Mi
jmpaeeoQUjeGRjpSyUYqpL5zzaYN+dpLCPZmfITdc/+RwG7oYLHDzKJ1dK1krnsr
SUYJW6oOVu069nBhv7gc306o8nI7WV1b/j8uaWD4D2U8xNfBnJFoO3q751b3I66Q
UWo7gUjFp29zWr7jJ8ov/JmgTDZsSe7H+TLKHeOUoRQCK4t7MPKSlT9QHB5QXLbK
1neH4ienVnrL0mOKf741uDtV6zuGqSmIql0KfaV/msysupgwEAZaszM1OS6A3GKw
7mkLz1DdvgdOTA77xwxIapmnCJ6N81U97wgMwuxLSWmNe4JTv5x62gpuu3FuLjds
bqD5KH00IrunBDXXcqeeIwNOoOSF6Fjo9TQXN3mHbOWXmV8thDdZbNI51EQ2Km4T
zWptWjBEdjYek65yCH/e5v43n/yl7X5RdYl3/26XSBHgQS0JcKuPTUuUJXxPWvvr
F1gXyHCR63JL5/cB6GB7DrWjUbcDZUTPbl4JgcgQNElYA2k7EncfuIgPWt0JZpWT
VkgRj/znA4xMDFPe26E0NNwi6JX3amA65PFqw4mhZocgvKBbDu+mnrwbPfNrmxE5
YI8veB1GujstrVddh/9kPT86A8EwqsiVKhA+VxKs9XHJDSTX8V+92IT2zD//XOHv
ZbCvMHN1BYOYjQo1HVKPCVQ0SMY5pbaGPfsFal3Ecl78N+sPUH9bCxq6d0wcYSJH
PWZTSi/V+ewILEZWomMPH1yq4iccUyhExDCkNl2E6bDN7+jJUtPrwcVBmKIu6ouD
v2GMQ+r7lUW1OKcszFNmankMYW8Vmg9VACuuDvWisMO2zlbq0GyoQ/EGIgCr4LIg
zQmRCRNDclZFey/NRv74JddFU99jwPFfCaTT6Zi0kH9pvaxHWWcgKpd9IpV2kIOo
EkWWxyfwSY7+aNHTw8mfFVeFLm6A2VUnqV1fv5n9ziTEkajDA9biLCFqEgwKI1nE
lAiAyI0/0fZTS2SeQhrT/3kBUHyxtLI0/jxapikMojpNuapxlMgIILPhn15FxOzx
A4GbvpCl6Y4q0tB77gkkBB3rDdqEXc8oBa6HMPTL3G83ViIPdg9ef1ZWOMH0StO3
wpDeQWfbQmHQoSgcnxkSbWKaFmdZ2VFc9vv5E51bENIZRlPjoXx8GRYt+VD05jVH
cXPQtrrwNHXOO72R60OwyaDqfO/4QL2PLSNPwjDwsl7KHMozj0T3mU6cGN1zpDN6
blcgMwLPkPwqCWINat+ryctSgTDArYLN2a+3RRmPwQIHsj54Yrwvzniur6jtzC7x
akxm11JrlVRxSAiiYj9X8YTDVS2YkWdAY9NQ3QS6HMYI4u+eX5A308tk0tty14yV
ZkLg7PLQ26f4/e27kFQiHc6VHLfwv/BZrUFBwJBduGGp+IkqFTM0G3O4xcN6lj9A
c6uEypWyISFi/9HfPcbTCdaSFg2+4G6LMOAHsf6P09hSqWDs+o+IddGU3GBiyj9q
vNevsC5akcSe6zhXSZnt09uDTLHMB7ax0u+GIa1oMhEKbxeUS8FQwXYgVCLjw0Ni
v1+3SSy2ZBwuIrnNnjZaircIMRs1NQ8q85tB2upxfe3cFxeJq/2DFR41I+Aiz5pX
0tMSqpt2XsrdWXpR//5V76H4G/RN6e+hvhKCOdw/F2yXVxre72ssxfBKb+ZDik+s
PezjeyGABtrtTy7TG9tQt9wVlqol8K0awYG6Rm/cahM8CTjT26GRYczAGDnX5hLc
d9MMnDB2gskh0IbPWEJ04QtewHEfqI3rdf3qssONGRaKrbO2NZ8mxMFsUhslHKF5
rQnr8LLUILB2c0Z3GEhUd3ls4gVKKRXh25ZFxOpbfi2eDnqtpJRhkXNrMKuBD/SJ
NjUiY30lYBI9oG5fO7RbvmJWH94TUZ37lEPAB0vankTWb3qtQaZXWOjs9UKkHMls
1fBx9O0itPLcm2d1l19Fu0CI/nX6N/BwzUivtFUQgDL20RvuoOb7BEvLBA29TnFy
FLUgEHQ7xkfTBCToAI8C+LvHBQh1BN73nizui90PYuxcl+BvvAdLOwyOYe64a5Pb
5wD25vKwwgdol8hPMNUtw1DKk583SriPhShD72OBKfa7OZRJOkNk3VwdJakLbYSL
pXHQWV0wGiVltd4v2SidralfknYXHrzhf0pqyEuSMLEOibvwWfppq3hndlA911so
1gYxkWRa1UI355cyRqbfCvacpSmvhf445k3a9IGsyX7Jmhaqm3w5cTuAzuVfjGae
dknME42khX8kGOhEFjnXL6UCVlmmw2fsydF5RIu0exSpoqfQXjSn48zz9YfxZ/ZL
wueOBCHMCANe0Mxg+C1IlVpHPLoUL2zReVJ0lcwm8McBy55LUTkuwWYrqL/W/9/c
DsE+zoqHoU9++bbUPSJu/tC8cmH8p/gwZNYNHHPOpZ7/OADlv+kicGoFC2x6/Vks
XshBmTdRriRMO9akWh/72AlccLCIC+jFjXpvdfG9wJRSUT3QiMcHr3fkuvHXRvXs
K+J/vSp+AS56nOdSS1B2yOdAmuf4e/DjtbpJ+/7cHBO6LhFPiZfj0PvC3+K5D6Eb
SnpibekuJtnqzxwJU48EpfxPkdDvy1rs+lNMxDGDt1ypCX3sASRyxCh0225t7dRF
8D3LlxCaIC2woW2o2CXxmUb3n5EqWHcIwmyBkye/VhBz371XtAS9cSeiRARgiX8G
ziKMizx/3W+yYMFTEMS1H6XjFRNb+HY6aHN+v3ifnZPjcC0qQuM0SJnpB3QxQkUH
3m3EXG+9se+FA+2oQTvEjmJzcQmftjD4osazEZFqNmpxd4YenCY4D7nxeLtBrZw4
xXDUzRbs4MEDpmtA7BivLZj+/9h7HzHcezyW+wQ7s+9vuDMRpOTBUlMQcR/CYiR0
45rsDDgFDKazV3Nfc7rgrAUQKjPmTi8/5FpzauwWfr7L5BWOGuUqzNI+ih/xwEAc
krbtrequJrjwGkrIeJuEOczwZJMmgapicG/td8XqiNd46A7vH4Q98UPar6mGGTt9
7EUwJkT65wWS25QIPyeT2p9i6oDRjg0R3yuMB1A15UU4V2wAuV+MEeIMCEqfvGDF
OPaf8fHss30RQXpzhXSRajMa1pqNBwjmMbQ5hLh517YtsXpNp5FlT0LiA+DcG+R6
YSwr1SDtjlPRUWM/RkAujHApS/WezeJTyBPE9ZjfmCW2za96HAkm8tbNm1NlCvSa
a0W9k2O/q68QEZsDGYN7SauNTlATbU0a+sjupsYnuDh6DqVnY9OvuHqdy+9oqJxr
PKkPIlrazpQ0HaKSgbbyXMZ2L8tssPguV9RVK63YVjIBa6Hkdgfu5plA/9g0dIT8
5CCPIWadNf13WE6XW3NoF/iQWzIOPNkoBhEfkR4aG4OSJ3e8gx2CiP3jmJdABGfl
5sJ5G7b6NdZjviQJMLv0uRTfUS/YnUO2YQ8nh7FNqMEyaybLuMn9CwhLMCBB8YZL
wjP6OKM7bAL2+vca8D0408jxrnbP+verhu6u8VOAOFjdA5M66e0VOq5QlMP43Emz
Nw5lGDx6Jlzi9pDBwNJ8x6GEBb1ySzXvJWEHCOC2mExPXuwf0bFOqTdRTwx/dEs+
5yaizAIAzPt8slVJgKoGvuK7wZiJsCMlH7xYfeUdeczLcNDSVJEo9ty+ollq1u5B
JG1bSI4bSf4Hfc6rWhqplsEV5y2WfdFJRFrMg1uxHtKjYqGa3ZybAJTU//EGDgHQ
COuCAVcXLUBSp6NQBq9doiU1VfSvnVlO5QPvGZNMNT+S2NAqUtuk036OZXGdJ056
oldzLPwBGaPKJeke6mvltI4wwnPh6eEgv+mlEE1lD0Q0RJEhQIP0S0VP12/b7lum
7P86gkBV3GCEaInrjU4z7C67ceH/Qq/WmTCWTnY98J/eeGTRZn1quXpDdK7nHq5k
5pRVm/U3mgps6E6FM0AxleZxGHe/mTOAAJd21epMc2LijBfoWKag8Av8rHx0JHHn
ctu5kSFVdB2iGncN50fwkdpLq8++rQ3voVrCUuecjARIfv7BMantyGChFbXSmEsT
T3i9pW0F8iJmcYGl+5UMjnJW1f4vbnzFdFgtGwBv85z/QznstQy8A4PSxz4oCZzs
GxG0EyTnemU7y5dM8Mgbo9rPm8n94jHMFT87pYzbrsAEM6e5lCKmR3zk7GtnWz/N
/mkFqRmL793qn+75KUBmMt68F9aaBZPO7skPhf6uCLLRyGVcdvBfgUmIPeLgVKuX
5sWxb2yd55+xwWl8+LkzSO4DJuM/IuwLrSopEhr4PRwKy2XJaNTAZdvt3UNP9Nax
d81RzM9kSzP4hEs7sjBXoDmnCsnG3G2aewAWqeVeDMqn8yTrfaA5Yv2lO947GI1b
L2HEE2M0zWdDsovASFx19V5g7gQeG2SZl4P37Tf+LBahcwV81HLX+y8kdzDX+s5A
1CB3240UqVr8tbPVQ3xv700hItVII3gnciMmEd8bQfWze08FNJOCtSVrCDzhhAOJ
2jcL0dLB/JcEnhtK5oRB+2+zVod1bu9/4ZN09wr2WZBD1EaJIHiUNK+rfMAsrZwo
7MtCe2wOjulgDRwsWhsPrK7hVg22aqGlsO+QKJqhjkMVit54sR6d/S71qwOdj/52
KDgKb6CUCVYfTcd7xqrUSdXwDCWl80fl7qxI+gxfLjR9exk0L5vP70/A1Y5EpFsy
L7PQxiGa0Abpd9txqWgLAxjMa0cixv00zu7tK7G6s86XUZfxwkioVzM3P4z6fTb9
3kMnDY4kW2SlEbZa83Sr90wVpzeX6/G+IfRWabOF5GfSnzKjBIukV88Zn6O5CgaE
En6NH0PDJTW0zYRDYzD8v8k7/UyzNZxdr8QBzKmNxLNWmM8ujv01Rw7c+gL/7WaD
VnM7sPffPRy57fG0kjKU6z1sqt8+FmALWU0nt5pi4ffmB11Rxi+AOt7rgXtAe1tt
5EY+1XQUV8PrVZqbsj/JwyAE1ncbl3aCk8VaAIQ3EEMB22fCHlb9vQVXmf7Z6wAm
Q0bw4ZWINwMfVJ5luTlghG3cIeAscxVKx4EN1w3SlT52xBBFtLSMW5jcJYLD5Yin
XVpsopgejIMe4IYSTjlJuzs+1MACSFwnFn/K6WiGbvfytPYgp+tv19XvwAvZyWVg
qrjSdr6TrhldJI16RgxrXfx4BZR2MRKOK355IjHFaVFrNrbs9IJuf201xC99vY/L
AwbrYXidRFNszewkADABCA+g1IBxyvZ8CF0+FqQB9d7VjkokV+HcBY07l36rrQuC
Ql0Y8F9LIWmC5lf3fOlKQw9byKGsBdkjDBf2JEpdimwbOeLqLNQOU3nrAJcH6OrL
Su9HHbtX1m1+4zqbUI7EA0fSTKXqpziedkX6BY4bULZvb4XUqQQl4sq0lkhJMAfR
P1qFwOYC/kDevhy7ByBytwhxaNMsRohauOd3K2MUIO6Khkq5tjxgWSpAU6kwyV6O
iqELBeoQ8gaWNbK4tnzFm7ddZ7gRhfOmVcluujt1R7tGmNmEq2tOn3fap734zbZh
c1oVFmcJv4l5PHpe9XycSxVMdSq34nZ1Csd2UoqaWq9j4uziLQ7MKOw7UnmN8IgG
MwH1yjhhZ8weFdiP5ZviEajVk8ZOD5lM5TgkM5z0NcEnIYhZ0ahhsKyo8FgdZGiU
mbB09ZjE5LWn8DJjY6bSLlsVpVfHVV7hpas/w1VFcPh4gjYKzRy1zP+cCI7VLJVO
M1k0g9dEOFDO35ovk8v+Ea21fSEE9afb8FATc6J8rKCSOhrChqI1HKrwGtoYwaer
bGHW7YJIegkqeH/6G+zh1ek0Tu+S67NgE8yF1gKzFJb4QBx7KTIqJaKemzh5dj3M
309T0OhrH3ZxYEkc507+C4VrIXarFnuRpwcHUEKJEg36sV3kI9vbpt6qRIl1/CXm
TWtlARhaxqevzTw6maUu+Wxdu2MvwgAtd633Xr77L1A5qbWbF+H8oqj5+s7QF0p1
9KuO3iYpRVroyKWJwIr/irztAifxwBNeC1LKMZ7HN9oV7zMIyQ7TTibGNSV7Lsh1
+9V6imBTvSm3Qtc3a6g7vRg5/vZYeaGsj3cZum478HLJyY/wd3TPlK1HzLLP/uGG
QPaQw6XMDzLW/3ZdPZixVzlHO0zpOF+EMD5co4rco02ahH8var1tUGKu++C3O4sX
1ySa9Uh/3d2MmWWaG3x3NFziJ3e0aEriUQ7bdRjxyYKAx3EO/Jsvobp+JQwPlQ3C
uRzscItF9DoznW0M1NQbKT02E/Cit8R+29jcLzwIibfAryQrWkq7qtqDKD8Qn5nV
tVWEOebKGj6aC01k1P4NVRIKWdg1tsFZGuv7U1vB4TZSWwWrvLkaC1EHd5x3KZm2
hKPZc5t7ZW1Dyo+XgqeshvPYcZT6aTWwMbJGIbF+W5IbKBaEj8zY3fMywsYrLX5C
t57AiE4mKHADVsq+hbVd1dteUGATilH+OgW5kHa7k0/PHt7T7X+sGRhDQcmgdseC
dv1ALZSTFxEDAGuhG1GP48Dqu3sBJ99kuSPRa5Tn1uzDRIHLTko8BP3zW1FP6QdG
TPpecUmoWRIIZ0zNs8gw0OCr7IV8Zxx0XUeYkF1pWchY1aiHddjQTzJ2iOTzkVVC
zssH+mAaH2wg0HyVk6CPEuKRY8fAnSkc3TqDuO506qc/7KvyPVsy9wXlt6VT7m6i
TBWEQCN+qEVhIlKhE49Yaxxq41jT0O/zdFwTJgYtjOjziPI/sUrHJ+DcUNQO7ibB
ohjqu+1bP7tARq7RJKi5zRk2s4hepWfM1/iJGUAn1GW/OnoJK5r5FBFi8g3Ppjre
yGMFH5oQVEBHheS0iB92fKdc1/xkv1YRZPUcVgGFklayqmrZ15//HnERX9E01FQQ
7TxsdLnqTfanQJrQwD34zVkBDVrixVRJqbw1wOKncOOKLyl1fWEEbfz3HT4JQUjp
ms8s0E7W/SZfq2mX7nfNiNjaY0BhR612Xa0T3yzgxEVApqyq0IVrB0kggkZO9Xs0
nikjDjgjQHsJQ67cFnguxHbeNHU5JH9kPwLb4XzmKgji9hyrq+INEBlpQ5baY8oY
VZo9tcvVuIFDNwxEAD3ht6Lgk0U0Al96VSfsPnYgTGl5uI16XBylyBbRfT2rrgN8
2hx4WAZ5BrdcKHMC2P87PpjHBEZnk2x13hptRuHMTcEEmK2JT35xEyp2NooS6I0N
IyoIgISUVi/Y+vp4cpK31Auml7csou0EiKz50A6XYjEGTqkxm4k7x2Lgnw0rMrDU
u+shyGeD5dQ1+z12xDU3y2nmj/fvciK1tMNFQDAfWmLRY4ATIKCvu7WDG0dzxe3x
nKRJthEUHe1lbu8sDzhhX8kwlvnzL///60dF7SY1Vck7bxcXkenUvTYYkH1sB7He
uT+xLy/ezdnGKCCCNX8yA1QatVkkv2kV3Vyygobiu1dtywOiY39SHj/JJztG/asb
WbV1Qho3TW2ZrxEZHa98aSHMYDygIzPGiKOHqCMX40+yBKo88Ck4sLjUF9ekhh+D
ZtrMa7KYjdorX7rcEmLuptZSPtpekdxctJjiACsFXLNwO0jMyx195glBP7hjDyBI
zsVul0+Gbuy9ZWIqE5V4vCFre9QwoUIxhehGm92EYKMjSYyR3a6gHEIl9EqtbFBf
IhVS71eltUN2Px0GtxEvvf8tVfvStyDPsXalV6uMTKuhVk+sR3T+n5zUjav1N9bC
dYS5ctKSZ3T7uah6SCBiqnAQ2L6boqN+KDj4od1AVJJ/Yss9Kem6xhlAZdMSwW6S
hBujZ3wBeaeNt6HqFSmu5dOY+P27cICISJCr34apG6CwK9Wk9BjE8fiVQsSq2SGh
rlt2Ep9THM44IBCTZz4Y4imVT1lpXp20RG0TElMmudSfvLgpJov+Djhu7GCGP7AI
SgFGM9ZIzui7Zynuv6/O7BxPoZWXDafACsQZxyr4RrKofqSrmf52NE1dsyOux8pV
4Gb+NCahnByteyQDJtOqyduH+I16uvdh49d4OpAjM0vAAZgON7T0SkJ+mNelsoLG
ewRmlj23NQI5MwdI4D12zMa9yd3QC02oQestVtjrTFo3bvRvV6qeQGBuqkAV7xhQ
p+eectM/HOtca5T0nRmw/abhwtvEdDfLN6i2IgBhVY/OBt1Qu2z6bApQyYhbSsE8
CQNHXBsI6AOCVKy2fh2zq+o7pTGYCyjm9BeOD1z1cTuiNIjSAaHJPTmDgA80PsLw
SclbFKx62ogfIqHx5LAPQ9Do7HgFx5ZynnlUlWp90YPnbU6GLyCoYAxHcqDSr93O
D8kRaE3HxSdmIepeXQ5TKupZOITEQYEUcwPbkHxeT2GVGCejslC/Bw13rvneR9LU
B6pmvMgplTnSff6SHj8l9SHwkocH1BT39PpBH8A1UkbqxLoEbCv1z4g8U9R+A36t
Ri3ipyHsi/st9IwvF10Jmd+GLW5RAbGl8ZrlN4PyfoOcMl6CMs4si/FZautDqrh0
vD6oob8B0zU3hqZfHbi5hP0mDoQi6FiyT+4/1gljbOsK5QyrwX6EssL0w2jJBfZb
DTj9EaeZ2vR9eN/dOlV3TfVT0cU/V1wmkHgkn59zeqz/g3Hwy1cFrZZjauTewsj0
01f0vpIsebObAXQ8RyEwnJnf0qO8BKPSOMJbWF0wICutwNDCSLZ/j3ebWtXIrFdY
CzgJOoUm9vJpCGfdzwMr0aD3pLNq3embXud8rXUsIjqVD4ccys6wPSG9GMMSc8fa
5A1/TyZ07qW0FFYZ6HeaoDbKpGWqNJOF/7e/Gj2irWtSTQssw559b02s3ipVAR9/
6Se9Z9CnNKDQrBMnw69TlmBBGw3AzODU0p8+bW4NzrJXYNRIPI64Brqzh/KvdQbE
AbYA0hOSgfEUzL6PW8I5hpk0ZGTKcdY6YiYdAzP+yGfsOwOyHLb3Fg1ELpw1Gbax
LQk4NfcrNMIDjUhRyjugMcx/ol2O3h2xtqWj7boBX8hju9ZO/SvdTUe6gxLyBm9J
/eXOM8yIWuHlrsagbS9rZ4Jhs9cWzVUKEXnA89YjTxD4uVoho4QEuMvB+o2Zcxs/
INp47wSTtgYHd1gF+CZV/qd4ppiBvVu2+d8eYDBo+KObGqp3Eh6sMjaO6Doukszj
UrbuZMdiw/CrqvRvvI/4tgSgqqFjEVJkZOfnNn0JZujMHmjgiebhsZqCez9yfkbA
66BWyj4RDBkYP1KbLIUv6NXnvW8YK+7btNqHqg+XhMoy06ZEpfogcoXWtu5bE78r
qYw4VNh8mrhEpLDhuHj6WHCBfMYEhU75wt8+V23PKh1ku3ttDAEU0ltYFrDdkNpr
DuQNfdreOVvw7QZXSnx+Qv3bHyEezf/oGeSISY5YjJ6AEQ+SJf9kknKM+RxYVEmB
ycLLU9Y2gjOr6wmoh2+lFow+vdXt+cMNmIeZHQIs7Ra0Rp/TFRU47cRRmHSmny7I
cSHKp12skcNe/yAFBFO3ZsJEyQyJWDtoBUzos6YxF0C2zm+v5/9WRc+9pFVdrnWt
YdE7aKFSMxg7fckHCJ+Ix4NgSqkNbSyLZ0mu2aheLQ8MVx2QWnCazGrCm24Tj8KR
stBr5uGdEjf2aXiS1PjXUgve2ERA/MeBPDL9a85DAydSnQ2l8tvnHlKJoHOmetYZ
KWukhDtSJH0FPH5fDIcn6hz1/BI80fZKq7fL/0aIbsOyMNA6OMmDhMFLFZF+DL8s
+wNIYkGdwZixWOBXeG7HOIrWelWoS1qVY+wi2Gp31/3ARO95AP1YP+OTTz+U6ZAY
3sEfXcRL9mzPY9B0Wc2SFLOAgh/xV6AK3bsWyq2//AD4czevMEx889jjrGNWzzhn
aRf2MiZ1Oh9aTPx1i8xErk2AFM7mByhl0tStIjB8IVS/EfQJBX13B2Eqj85uSIeR
K1GeVl/v4g3Bq8iYP7+e3s6/dzYPLoki2l+5ItFHcYbJJL68t1WYOM8kcwhxbFZf
0t/z5bsoKiGrsn02qMzQ006xDjq4UWHyvce8i8L3at4lSBtc4OW6aZzoVthX4VS2
KseVBh9uMdFdavlhLbU/jT/fDsVI83d5DlAX2eyYTPBxv8xHUI/SGvZejYIw7+jC
qWuRzuGuAWg4Mk6Np5fFm/HqUM2mb9hHxriz5YHfKAiAiIDDoJNzYoW3YeJDEoSh
YRpGExYeMuxUjw4YItF3OzTS9CSLkMyWPI6xxcz2FwumbR588RSXs7jGaHlkhePs
v41nOkJrZ2On3GLejZnIDo8kBEzSNj0DKbiSNeDtiLB3bPsTmpFX3M6LVAtt3xQG
DcDnw8UU6ZN5NPMjU3f3hgSVYbn+1ML38hP7l7vSRMa6KKGxIql70u4V2rCb4ZpC
z3dr8+UzOioWqNKqMXS7fLb9F1hhIAhJ5SqYgthgSksipotbYDZJBII5Iiu8hHiS
4j++I+4EE+qTKqN8fFLMOZX//0Jst2P0E1PQrEKQ8bOpiFoYwQRsv1YFWedU+KIq
V9VMF2ImYVNrGGpx0UCXJteFSD9ZiFtxgqaWVg1S5bvz7dFMeDCaBKh/8k8Pf7zq
uN/dSwZaTnSN4N/ZjTcdz+PMUNqDpJ59X4wtts0rVCEIoZgdOTYJqWJ/g/W2KUyY
6eGjEbGHvWURJJ1NgaXPUQnD9tCdjmXbyhOE9mkwyVSnsQhDpLWNm7kJSKoB+EKT
vfhDy4M5v8UM8dMsjVAJaH5YzWwJM0pCeXfuxLBS5uc3ELXMLdcGaiasCCNVhgmt
Ni5jUkftHKxUmeb/1SOqDhl8iaXiZRkUdiaEusaHti6+26YSNJ6CF8oVSf2DbrQw
N/mKibimIWjjgDiV7ausnP2ttp/iX9eivT7cETAphvMZcyvRJyY1wVjblMOOi4Mm
PFCb1miUtWYHlbuTGQI1OQEM7ZdtL1OZ0Gp6JcqZIKrA3aXdObpB31W8FZX+565X
1guudCtBgCPXBgwNkuMX1cxGRlhC9WfjSC+/x+y3ZJsYv96O/Bl9TMBrv1QA/fAy
aym2M8A5T4f0ezo+lmrYbt9JyfGl3M/JL3CIcl0DFrGcHUYM/2Uq7hCmz/r6RGAv
SyPUjKU7thbsdaAkXmzF6s0ljWI/tAy2zGVSdtrIE2ZpqOkbTAvPLByJI0PBoL+/
HMyGstX6hDpM/UEIpHzYcZTY613zdZOx0/6Op3Uu1C1BmgccJTtX0onF207Pb3Zv
ST4Q9UcgRpQ61wAcO5jb96RZUnkqnc9vhdbepZQW6S31OO/8kbkaktNyrXzRPmQ0
DiyffkRL22A1meUOKf7/Q5hLZ7CEC32LbuOtgRO44m+FaBWSGRynd05sMblOt4t7
4vlW6sg4Qr8flKmXHmKocDpHOpZlRwc3+fcyjLYeZq9PrW5H2JcfiJ6eaLwbILUE
B9S/Mk6uyThjA5h+JNTkhdSFVOKSAXcDYkwlJIP09DUAR/FhljRpgDPeCmOhPtWV
UEherINk1MIjmI53UdPoWHmZuDgucoQaijDLN5fw/GnFZwnIbL31APqdocwFhioI
8i5ieEUM8GwaRyZwJaWYSicEsmP6DA7KOUE+EI4g3yq+y02ZsxKAwY/BUMukDKV8
/T93gRHqJzM7ygWXpRwjF6hSN28ItFS0DvHyVH1EkmCKlJEEga/BfkBODXFy4TRv
RnnaBG30aBFvZOHx6b0NiXr9QgTCd6ZV9bn4/e0b22J9ILGPNsceS5tpyWYkagJq
5uE+rCrzzXdDxHyXjZS76WBnHDr0vcjcAbi5BIj6NVoHIGbaWrKxdZLHAPQcKxQD
fprPJgOK/2yvpxau3RVL9jagUpcZbHddob5ttAZb8Xd80FhZN6IhsYvMep+4sFBH
HNpEOPEnMsSddrPrtjB5iuozuEFQ5pwjPxGDfXV4JrDQ/dEJsGkZEPfpHloGc2L+
jwr2Q1lc3ESnjsPZIXmsXZ10fLLhQIUvtSEXUjkAYavHIIXd7AP/E0+6atCiuxT3
oDo/ChmYz5jn7/GvfLI63y+DNMlQMjs+DgS0kf8+ZefJMp01Z23qtc3g4poVM90V
aMCYIgVhH2vHvamTwddliA1qtK/Eb+vD+Fxye34cvU1XcdiG1CPsW6Fzb31dycX5
j8gdw79iWcjnTZxfat5u87y668prnSk3l/0WTH8lxSQvlMfo9Ci9SJr8LpQq7qIe
bl/3Mj3tVkrCLLgdc5fAAkGJIEbrB2Dtt2p04A1u+QRuUwjjvNEfkgFLcVbVal5W
Npg/tCgHPg8WmbTEXF/IriYbXoGjs9GRQNb+aFWC10fG7iSZswHz/ieJTs+6u53m
dHc9dr8rKRPLIcg5H4hutGzC+OowGhkehP2u8avKpVwXx3ZpJzAPnQVHY3RiTbU9
vLP0DlLBGDeA8GDpkLBbGyH0E3V1azHGVCqjhIh6Oylnqnaqt/GZd4YmjcAXlCOH
2vtxJKgeEfIuyltsatfujMICs4ScSnTwzUyTbEPVAhUYPwHuX9QMeoaXWRQ6L4Tn
P87bDiNAiX3iNB36W7mz0OQ4iP2lOMZ+j3xxs+/MVrUfAmfr0btYiKlLBBQP9bIU
QuKLon+uk13BjgAsnUA0buJCWddOeDq1CYpwC0FT+nfTvl9GlCZjhozZ2cIm2se9
dgXESPmsnO6PN05udElzC2ZPNln3IydfwQ1Zv1dhhuIxVn3FGOKBNC5WgRHlv4yL
KdlAPlnb47MOAukINv2BP6qx+ixE8va8skvVHLbV1Im6laW2BdDSFTNQMOZ/b/UW
T8xPLCVYPYUEztR3GRv1wBIngeQCLd7MFTtxWeE0BUPQ22msxZ33JSi/cTwkzZHm
RTDKhy3VAmVEmUYIUNqLja+rF+/EWobLtqNr09DIuXBobNPBkScIYIzQyWdYxzQ0
q1xZv/0JcXt6ntr5LRgm3Rqap4cdTsuGfyL/GQpE+tBbnEkylV4MQ9GgFAuZTBOX
/tnB25KvnZJ0NMD0WLF+myWE+zNy6eW3GJdd71EZva2Kp1QnQt/LfkDE2fTRL6gd
RLavjBnHlwlgvkEr8v9Oa9WpBvBUySzyAYXAjRw2jV3tabVVliGuNFzCODsIHUxJ
IqVaIUFUCKsGX3bYNjfWIaLVWJcaeQdRG979F7Usn/7P5OrP4tqqEgPQkFoRMNI6
5cX3Dy3KtBqraxMx+mTJaRXGdBSb/GaPMIozZDtjweyMAUFLZol+uC03buRPhO2U
Wtumy26oWuzqpsID6HKE00RMHlour5K+nzLUNgTGZPiUFeZFYqioqKINDqFh1KzC
HcodMw/udOKwGXjs/aXm+TJAhypdAyhRFtgBkkM0J3BJ64DGayyQfjmnYBvkwiu0
W70bs3TO9iJ5Mn+VSLgsHfbIoQWjAo3symBiPBES5BYE7QZg0IOUL0niwXiHTmU7
74n+Kc1oi+oM8j0BjFhrdum2J1CcaH8j05KN5ECCvBGZzUZuip9lx2z/DzjA6d5V
V2P0WIqiQ/X4BhirYqNX+nSxhB1RPMd3DIkK0vKoYwEJXpVvzGJnmG691pjglVdd
aCJw4ZfJ0r835XoS74500+TFXhrWqeqIMsz44qtZIEvi/C3GQRa7o+fB+AdWShpg
mGyE1fObljl99xBq+JwBmkTC+WhmQHA8t9UWlsNUSqTGjsSyrgpQ68Akx6W9MGd1
wFMMG/tbdRRyvl4TtQbfsNQ/lrKuslHVmPgbP5w/2YCXDYPn+ZKOxhDvAHhOEuaN
C0frCN2Rfcl60Xy+OdP1M/+07xJrus1ry/OBgZf6AOaxk2fyQ13I13BF7j+B025J
b+zwaVLswrKAzkiZYSV5av7JQ4s6U647HtS7k4Ihbq8RrEgFg0FiCxRkXpJHuauy
9LA6idmvpGqvo2kJIL0BKomdr4ZZgyxbC0E2aAgaBD++tXU8uIoyj/pqVZ2mQAHC
rDD+DiqW5EnphbqTXP3usF+gyRiAEhaSAy6VZgxxP4ZcCfuy347F0esyNAmn95TM
fHxGSot7UWQKQrVRBK0Jo2Dh7WQKFPE4Txco8dWypjD912DriDZ1H3baVlhoxT9E
vUp4AtKlfMC/uDdz1R0ZzA75omaNpan0y+4zCPooUtyuPjFuT3a2/0jprrp5f8/J
Gf7FGCW9qhBOUS3Uou9LL7HQGld7G5AfnMGWg73FfuGOOPVOWHjpvTtXsIAFPuTL
DaheDuH71j1E3Gn5hp6fqrTuZwg03dnPOwCr+etob0OEeHBR7O2imGpfToxpFeUV
p66kYZxaD/NtUv+L/tmAZ49LBifT4KSAmFJ73TfuZBERW8EnUeLoYNzOAT0G4J0R
r5ryV/ruiR20LvNHBjnVojXYkpER8EMKHp39ehyMgjWqJE5NXPLHhoMQA/p/fYcA
RyJEz/Dh1ev9ia5aoBijbZgnO3VgCUyFPuElLKQIv6coVURMqVNgHD2acMxRSEqY
qkx/0i0pq9GfWWgB6+MVlJ/hnsQpCnO7CovLYU9dtRa3WqgOik0OpXM+ynjma/V5
WIb/I2gibxt5+CzjdhewPDjNuzGRxpUzK5JlVE1sJPquobU3Y9fn++u6OaSrtAVg
3qxwmuxnF2UfXBA9waMbizsx7Ow0Qz3/uvGeZtFsBBRXdd4WagPWuVf97Z0w8Prz
yc0q157Bwy7cl1gb6E2QPjovRZ3j53esqb04WXM28DlGO/lYV5FDRd4i9vOq1Sib
bHDkrdPAKa5edP1tAbrmXaMtO0rNskcez/ox1iYZpQN2mTKAoIDVQCykdIzhH6th
i85pYG6rMO3vvV80loTgPwNgVsppdpEI2631Ny0rVFwaqmAGNzHT3P5VmoH2VgCq
GUaYsvPdt3GWeKqMDXluEubY5hsQON4XRnjmW26q/gLKhf7DDwiFMPJNVwxf3Nkr
qcuDGmF09vXSe4xfyMuQ0GG95SgEDiqIxdjWfdWyVE8osXiCdXjXunXPOccZuoHM
0G3OmGEStM0pEP7GVFNdW1iDBUhUDcSkLQjM9LjtjNLW1L6eMbDiSaoTIX5N8lb+
PVhi5J0z31CkDyLNiPoUur2g1RSaKGbFUWaUdH8av5zRlGvTbebtrLswMJrXfGYH
115C63V9/8ihBmgg1cPuPTgC6Qg8cihyypBeuQY2UABB0B5osUTj/92tBwgQ0t5H
q33h6AvGgbXpYgfXvAhawNALV+JaKKjAx5AidmelVOtdktU/7S1d2JTntaUtZkGV
1m20rqmd/2JIY2cbHIMOT80c7CUv1+alhFUS9ki/Q5ZHl6VNjEQHj2WHfWqGlN18
YezM7PTfrAmRytmH/UhvCBXQe+8KyNHD1JB3mF0BJ+dJZTz9cWeAJr8Gpa10Ldoi
ySwl9ykyc3a1Dp28r7OBWEeJSXzFgFVuNFXOcG1hGgUkzP8xrmftCOyuXIw+kmY1
CE68iZjoKc2kp9/YatNBSvKayYuIDOCsfNPCgUoJElCvcWNfC61LLsM+LSe9iIAW
gb3LI8MgynGTfvs86pnltd0eMNB64Ylo7BfInsrUM//lV2tuv95172HdtcQDCoLa
k7Il5i+DBSO2ryUjADgMOcQqVvzbsPJeD3GmW3PqN3ymhob86Cwq71tWxQW5wfXN
FbyB5H/g5BDdgl5yU7M+5vmbRACUSQ/7xKPm/RxII8Iiyjvcvba9dQeqgsOFd1DQ
9EsLLMYVk0QLWGkGIuopUaNjnaw50GegKZv/Bck8qERHKaGEBzqg5CRA7yt4az9R
U+XV3bbPrsI0EYxwwNrYk4E/rH7mo1rdk6twE4I5R1Ty7CDxei+Va0ns0wKkIpMb
ykS23cWbgwphl2yMZ/XO2CTFXJeznAaz8VvE+3/L41M2VO1cblch0cqf70rQhVWu
OI24W0CFXFNFGgwgE+ErjMNo2/5gbgTFT+HyeT4KgMFmWPG8PMSbCf3NzHy2/fv/
qqvYTQJKZmkk+RtlVVxZlkreYt0gk2bEjQ7AUiHMz6YLv4I7CEHAa+pOMGDkh0Vt
/qS8WeQoNHD5TDK1ug28Yx82RAnolAM0A4npaUynTs7/Sy0/xiACcSaYwCV1ciim
Xf9krvPRJD4Wd8kzGhfCHpXRnQNFep+9MwXnI94EAm/I1V1Ndf/UbuBoBrEjU1eQ
dsHxwpmiYz6Xf7W4RU2YoEzIwE96iEmeg63clgGEwxtuEV5vk1EI5RXSp40+d5Qa
akkfV0PXeGYHpyIVTytnxPwUsB5VaN74nP+Gf2yJOnJyazTAUQFvIs8fQQrdk+2P
79+Cbo0Xbk1yxG1pP6v+IZ75cWwZRnP9e/PD4BeSDK5TJZ9OZiS0es7C1X9ackAt
fcybxT7KhFliGKtTZq3zaca3dRQa6X1hHLRD9dmqK/PNuuT+rnwHsPq8BSyYaFnN
5Bzo86U0E8J4uJ1ZLFYza/3NG5DgTjkM3s8Ck5RB4kWqDZd778fOIMO+ZwLZDfuI
rQNerroyRm3KdkwAMIXSBvSMn05HkJPFC1mDlatXVlnRBZpERoNmb84h6CN8Zz+I
IWI2H2TU5qhkumREcewUmftczLvGc2d+WTJHtFhsy0DIGyA7j/OHQv0ELbQ79DY2
vD7G894hiRTOPbI7PZBeTN6apprBXwtJmZKdG756xL5bcxqVqfW0ojTETTuJtVeI
VUPJYRYfYeHhvqQ+p54PptK84Z2gFWb1ThO+Xwftye5qeZJTa4LGoOqlKPmgTbzZ
7NJdZZqAQu/OYjPkaCkxbILEzN8rBzhK0zEzhi0KoVBT5/6FZ3kdglFXG5DvGgyJ
S9CYN9lpftkG/XzgGyujlhCubdbKYG0sRJjvoxMIfLX+IXYrRO1yUF2hbpF/EbRq
3g/CcwIepjCsYoqAOwZBQjCNztzPSvKG+ztlQYYjyxjCmgS/+yHdJtLeHjZvVGLG
GR/lZ+QxFRWvccseZXjijCET7E0mZzPPSYiflzYt4slpLRIkPAjYCzxMhTsgVkNj
CCJj68layAtpSpZ/VcakVe8LSBdRVZXkU4K2UhyYx7DTzM6Zkv07QkE1O+0316ne
YAcYllZ7PFhafuB2IbtXKDf0ybw2If+Eqcy9kIznOCEcqPzX8bDPCdcJtwl99HVJ
bpIy8fnhveQTULOniHZI8f+wl/Ao5cSqzXqjrN5005G3fel31mdPX6wUM8Cfo6OJ
3dTL7rAbTCHLUxKUBLdZv1/jLYWxeTy4H+aM6P5SN1a7DCnHyiNmqIdcj/J7Xihp
KaWr0viRGNUNG+u9SndID8+6tGcQdr9x2tZuWVMK5j3VlDkf3qmJCkAO1T8YF/0I
xlHSzdEZRPDePkXbpv+qAl808bMjnnWzG/akR/TckWirhAHitBAAj8tKJszlZID5
XNBg5niiOOS4vIZVGsFI7UMFp2quzeFQ+lJe+BaAvl72dmBT26tj3PIJ9WejlRoq
1j9Ry6Lk6QMyusxzraER0HPuMtqVbGipYUpNsva/TlklzmYwcu3HYJ2So4/XXvgr
iH2JPeVBoG+l0cLk75p1dZ6xE1sfGxN3hReJYlOiTVTJDVJ9y7hI3Y1uYbC0pi7I
JCfmGWn7H5WuAGjCe82H7ty1ozeB+jfBLsE8gF5Zg8ikgww+qUZ5620zvgEZONcO
wT4JQBJwO5SVWZQ5WLGQp9zSqsJQSNVF3tnS787uZ8Lv3fO2GNc9vY1ixXNIkomW
H46CQARaK0Q2au5YyTj8tQ90PJhlbqvNo4zgBF4RlXx6y4fyOwsWIRFBMKveL253
MBqDJWh1+u6D3H3QOYrDblxEpB3iSSHdDgDEKZcSr0EZLvYO5K4pSb3AOQwvfFpP
JTHlGPpEK5H5f/oB/chiKAIir/QXpHLIpINhlmGlWdjmBG0RETNIqNlInmt4+Jg8
fn+Y5TVzw1ZjBqPkuyvtQeAcZOLVGRUUAvErr1mWKoLj9HwLqPdg5EI3uhTOrhyt
r7UwW0QqeiCPOa/xqh6BguHviyb50ueKHj7gCDXv55/KE8oNSTtXheNV7+tZmMzn
O5tYirKhzwn+AeyCmfBaL0GDlxWFNEf/qPGaFcRtNB08lc4Enso3vVvlktlQGrje
B3cVZ4jEufEil0MiwADa3mV09AocGnHkNecKsI93JoXKLunHRZ9YWO7TcpjkXNYI
cM+XQRM9FB8oA8SCkSH3CL9epVO+a9/04N0FaBZqVLRUMXr7nRuYgqb9mD4vRIUZ
5zc5aMCDD3DgRDDLqPEd/+njeGxO4gnpPdvITAnHeCNhJX4VQbXkrDuMVG0aF6Cy
+YFaLZ6pSjRjVun7A+7tLA/g/G4j+V1297ZS4jQ65lQRu2SyNicqZi60k3qLVOsN
idkxSd50zb0STbbQBPGh2Z4NWNEPaes5Jzs4Gy2A8RmYWaJ8p2mb53u3mx219PFr
KrSlISkPIwV2ZRzCQtfMAw18pcVyyv57NhZkk0qXTdOuR82s3xNpQIFX6xgQhwe/
mnj9nrS5okZaEDYXfEYW49Gh2OrfLMUh67BnooyExWKOuHoNGAYXeanNbGa15/QH
srzuXvy3x1/avsQEsKqS//cVfC71YcF5n+2FjKd5aXRB09NXy18q2xM+v5UFgykf
uD9mx6XGSX4BP2UxkmVlQaBQ2Vr1z7kQrWK8mI10argwVev+4yY+ueg3MbBaHa6Q
P5+7LEv7majstGMDMikjfJ0Cn2AxXo703l8MsyOInMJ2UKn+KQpUOL78ZWL6jLsF
8c8K4GxKmDRHT9bJTKNgF8Jul1kJP/AkhwHO+pC+TsWEBTIPB0GSJsA3PgjAZlg0
oIcnsmNijBrKz1ch3pKcFs8ss0L3e937KFOXlzc3/u51YCWrXDWkf9dLo0rQ6wTf
TqhAv7EGoVrNQ3ogFC3zqOWXMoT4GUCOzi8JQsh8FyHobvE7GrjnmIzjPhU6rlad
kXG6AXqH/Y+jj8SkQAzKfloUIOyNXi0PWJuStARxO2njykBnBykLZOLGDvMsxKi3
tEJVb0CB6C3/d+cUDAwRZbLFKgzq6rsMZQ7v1cn0pYCCI39+CXlfm9GUQZ3P7mf3
RRBEoT0H49UARnpH1lr15vCV+Uf6lLqgX3ZreGXHXwUajvpIIF0/Le+SqaRuqh2h
WQmNNWssZw/9Q4LqctAxINsW+aX1oOwiLy64gBL+N3u9pWAs5vTiLwxGsRwQjWH/
uIkkDk6JwJTvcH6r2g6/zCBs5qu8Yf1TDeD/9P8joMrF8U6eTQsQjnkSzfGFf/Cg
cPo6MiWrVVFBHkoSDvOT72vqDsBYqs45pJdHAGgs1yyJk+Qv7ANnTAm0HcjsSnvd
LZXISRDTpUh/lpVTDPRrmgnZ0seaSyH+6fKdBYqyGcbfPhU2AB2aPefNxiJfivS9
EVIlYLGAUXXxoFmFPQyNaR9JMBig4kyAveYTn+vNtcgwN5YonQzPG7Pn9nehVgyW
cRDN0oidTIZOEupX56AekV4tNoUh4HIW7XCc5XWYwfjtX4VOEWiyroFGHgON9MsV
CHS4xLWoPUzJyO84reS8a1u6Dc45fjZhDDqXXimwNdOsmuD2SlLnojfdmiDBEVi6
B9QAeDpHODNx4FHPVjolF+slCHw5IuR7wYcsNupdPw6kDp1J17IwxDcyUvpdOf4n
3K3JxwZExqAD2UBKL8uSs9UmatpgPtJlqSZBHHg8Nkugkeno2k1ROltzLxMKGaJx
B1w5q6J3MpNpmH8pjb4qQZFXYv/MTEEYHrkVzhlWQcEIDXn8FkUIGBwNk1MuWXNu
LfdBr0pMpsliU+KsIYfsj7YjPgNgxtQl9tAxqMG1QiElCi8lRqxQJqtDvjw7kjOv
q0R7/O/ibdRxfc7qBVMGBI4CDymiTEAlbd4KVcjU2SSiVAkF4siDLTyZFqBZAYh6
oQy3CBJzeb7d4GXFZECIMMdUksQnZVDu7C+nhYRjgqF3nxkj/eyHt6/E4H4tCB+F
mlIpldPlY6g70u/ArplmeMSaPK8/B/9kx+n/qDUdn424hD/hy9yIp1gIryfMpSqo
2LlnO/9BG3y+4aQFy+n7LrgtZWd9+48x9xG2kHgjWtWG+dOYjyM+e5MYmAbMX4eC
RhR4r6wfZs7j+4P7oZxWraAAFkVeug3/YlLeIRIU07v8+CDqbLe9OcKWaP/mKSHZ
kyFdr+MIBhD3fh3wDASSpYc4pTJpavEpPx01kiotMp1vRbRBwweZW4zcnkIABZ7e
UuSVEG7u9aohkP9foYZOivfMuN5UaBlj3qFaGchsEvSMYpI3PI9ldtCKXa1LLyG6
fJ8VYjDeNQwfjMmUS/KM/R3IJqp8SlbTAaT8kTtWDf7iYA2nditiiXvO9LwB1Vnr
pZKQwNlopyDPQTqZLIOvRRi8o1LS8ZKxf5xWN36SFBdF8TDWX0A48daM1Xk3HoN8
hDyOPgBpKLmYI3iIRb2p3dBODGOlxo2fug8Us3xlAO9HUxM+C57645R4gjDIixZl
U13dnW9vqsg6r8RDde7b3ZAI5CFsE42gtZ67qFBWUxJYxLCwDljEv3jZlPalMmWH
YmVdd0yHhMSY2lktveKVvKoRpEjiUjjcUlWDLvi6V+R0guPvGPhqRjKRGxKnsoVl
rTNkhifkzK5NsWBSfXKMJs9qpCPLk1G0JX2YDBeZ1/cNZHQ/Xi5ic6sk9FUOclH+
P6UNdnJ9mLMascfSKxGWcHTmDJD38RFevRAwBcTw3okkARXqrJmNrX9T6jNBJiQr
/+7+2a127LUbHqJkxalhD3h/radyxXmECFGCGF8TQVNILbhAuxnF2fmzeJg34j4C
rdN4PUrhAQlnwdiXdIk3WhS4ugo9liaH6960XZxDtn7/OBannyjLA9B3V7cXmHVV
8Fj70EiyZKLjyndVHr10YwgguC+9l/hFKe3iVmSfACyibQZPr6cSdpqsfgr0OKwM
VZScRqVyR+34FR2l9DKm/GPSn9BNSGFSePdFKlB1U46F1HcX/rQb3yNe0aGWPOTh
P0okyANrjDllecUFlzO5qhCs1NpZ/hQuA0vovLz4cXtUJSOwbFDfuQ7e2oVbehSs
kYG8yyEZTfm6eNQcVTqWBOpz0puqycn8Amy+MDpm/duHcM0xELPLh9MiStchxe/6
eFFEM5dMCIT7Vw6QxFpdXmv51ws9o4xt36Siys6WG4CsJDUDhsDVKb7fLfoYhanu
ZbiTFdYl1Sdn0NNoPy6tbFRDCFuLszUXk+EQeU79FtXAonqdG9m/vsDGFHa7kpdn
PYYYiSQ52zyvxLGRkEzs21hLYnIi5B+Tmii5eujYggRl3k8X/nVW+dk+FZMrbwL6
fYGi5HPzIbu8ushy5e18shUsyEZkpm/yTcBCrsh/+tzvlCO2ZK22TpW/2mfCA1RK
bQH10jXMh0B6gBwk9bU1BW9XjCKtw62Oo3712jsJJh7d8qZcHRGM4TeEwpsCJ21U
qO/mvfGcMyc0vjWq/ahOd85xwe9tB4VKzN6zm5DbCRGZyEJahHtC4XVpnXd8PGHc
p63toN9RxNPyZRR4LHYZ/VH8TjWmPX8HhSVq8uxDjcmhh3WUSW0P2armZq2V9VsC
mK2XJL+qpDWCac26RlfTurOIfdA7ezwP8qlvLrkMbOEm23cKRQcpP1FmksJgnM1/
h/CgTMVpZKzwzXzre6FJN7Irop5gIu7WKkl4qxgiHNbtfk1v0D8p30T05Kl3ubNP
/UsCUEK9vFSbL2D0CVInuqIArIm7HemaSi8lu1ZEy8z+y+pv91a73UACWynj7Md+
eJMxe1gx3ZXuA8WcRmM+AE7LWSLfrJzdc7woifAxDmejF0stl0CYSbYqU0WmYi/8
GI7hmJoni8CrvKophNadIF9WaHsEVdpZJvcUw20LLAR2615HennvuAat83AZzuCd
14yjFt84Yhx2Pwzm0xKghfBOciOhxDCsck4u+EiMBSx5QdYzolBQw21ip149sVTG
S36JgDZJTwQ+rU7AJ+9s34+NPAiCYN4DnTCW0yycCfVZLgy9KopebS6Y2j5aYb3k
1sm2zLmiTJuQsuqt39u/IB22Oi8LERn5WxjNzrbtuBo6GbkNMBxPhHinuRObEgM7
/G6YmWiSObsFvBlqa3Kfrqv15eqgOaC2+bdb0cX9FhjQCU/30QhOiWfKY2h3W5Ko
ZL2E12KytGhDNI6fpCmiEdbW5oN1T+pYgSrvGNs3w2bh3ZEek5U2hgf4uz1LHaCI
QANIq0ddLynzoQqO4JzvuwAIW/iTFKkuM4bZTF9cDheSAu7sU5boJAA5SE/WscRb
O2kv+koeImp5KAUNwWE0TZ79kw5lLANOOgHLDcxK5DFqKQRNbidMPkyg/IO86TCy
93WLX/Z5uyEQju/L2jaAyaI8bYi/OYDtSY7y1lcZ5n9xRt6OAqAxhwrcLaiaW2AX
RvS13Z2yOnQ7JgBb29s9/LeBKdtuKAb/Vn3FbiMww/WFf8E9a2ziwHHQnP6lRH64
zuLzr40boPjocro3VLxmZ/QYuiI0a3HZpCyevJDrKECpiyELyBH0Rm+ne7+QjlS4
cCDQw2Bze4hGKOAhVYNVqfO0Edf0vBnuj2kMsRNkvD/mgH1zmkZji/arODL2VnNB
PUkGsm07PsCKE7hOFCbvPtDuK2PAZNKYXyRpm6HLSehm+XdHfQI06glufud3fX0V
SgU3ImlO8CPteDhkyGQf5PJ957M9B8NGGcAsSTZqETUfTJ/fdiYvVAVC/8xuHfif
t0XRCbiun5+txzf27PCvKmtd/sKuZYB0315zPLOu0Ax1lLZje+kxqygbaTj3jPHA
R4mdIKK+Y/H0Tprvw+9lJ30VQFFzIB967D6hZ8qCDe5WZ9qsPwVIaGcQJIBjmn+a
5kja6LwOyU0w3U3VNL4JlEgJ41vb6qOPpRLDvnglhwmJZLlEagIosAIai5ucZdm0
rh8f4xQSCkNFJbhL7yq3sJ2jbqXuqacpneNEYNCEV61quVKKE5S+qO8QfBKFIL8z
QgjXlJEEhEP4GqercHcLjwE2GGgVsWpLpCrnvBXKiXkZV5PwMaXjgbtk0tpY2SbS
QdTWM4xKLJdUTFZ2mIQwHDkN9sjyQ5r4AEakxVFdu8Byy3EfNcEweV7XWAZykETy
7GqhSWhljmzvy1nShZiwphn7LrN0ouBQYLVlIMzZaCch6R+J4okao2Whr62eDj4J
YZqTF/3W1DUYmHToSjG4/SwpumYhHGSY7SKRPdI25/Fujvbkmtt6Id3PXPz1Prp4
71JYAOa5k7Mruq5E/LXtFiOUh9l9Q44adjdmjdx5KCmgh13p5Ll0ng62RlQq11tL
j5Hry0uHUEQU4NiFMteSkLeiVX+NYzERhC/DW9inidtfoy6H//CpPlFCxtyMo4ZV
YzL8Lu+7EvEuRYct37xpvlf4R64Mb9L4gMs0lF5xTF2qp8UneGBuRx31XpsecnuR
H8l4xyJwHcnnFNYoCD1WWUIUWHsFFK4lku3eKuq9RKOyF5Jx2j9GlvItZv3eXyF4
x8baCXvc9bcRRaLul1jyBdjsbf6+4odBx2n68XINr9IdKwvbR1+mPVpJp5AAB7DJ
VBCssgXpytPVUfx7M3tc7p0gVBZol/oV9hZjyIjtdXDiN7ciBpQ5yGb37NuntOM3
j+i9olKxlfKgdpUE0m1Pa6C0TXpisW2dohzD1qnBCWFkgH1LnjHhVkhqdPRQSXlZ
bhW8819e0Vtkrm/RrKYcOVo+oQNPUiDvHo3bSWItDFrfFXAH6Aw9laIslNAXnHgS
BZloTgL9pf0zH8IA68TEewrJTi7WwTZasjyVC0ldi6Lbr/V6UkhR0vawd83eZkpS
KgJNZaYGZV6s/GqpcyS8D6zDsCUMpj1Nk+awxc39i/rUuWVfjVFxv0uq0L/LuC1C
DMreLwXcndM9ba/334ultURKTI8kk3QkYACbBRKHSQLhoWdgBCgrsZot81HhaVQ6
k2GURvfXCUrcKCqWIBIk+Y61CKOQTg+LyxGv1HaOlKLr4bz1oP5xp+wV92L6wDd5
S1HwJ3XU/4jeHYIZwRBSOKq1pjeJmGREMJRQABhQuAolH/ZQtaVonNDz0CzEnM7p
iNm7r9qeNrHfTGwFmveUQhvWpIyPqOjEVXg7NXQv7qmRZ2Q8Ia9LOvBSZC8k7tpy
j4v/9U6pLsjKXmahSAF7L9/1//GIvsqTw1D4lS+hRSf1Ju293dToDNkr05QeWyIn
DizNzZCUho+Nh1/ftgJ6L1YtFVqBHRGOgV86DxTO0JczjboJEkDFMXAasmtdINlg
a0Udz83TUKbO631v78pnM1w+rogzwW/lah/KgvcdRmxlJ1mk15D8Hnr6qULHg2dI
dD8xLHMhx/Fi06KRxhmnEnER/l8MlTo3ENxKLK3/FrOTXtYYkQAPcRNBDGrzZHm3
Uet9LKcMeKJuUEN9l96EErbQ0pAvILTwEL1XQbm1PuK3tjSIXsXWI0sQ3Lr/wgdY
got9d2kGHTGr9sy3Rjrwifg1jbgyQYRGFkGzpTEHMEb0liBQ/OajM0+apECLRTKF
T1npXCP4AuyM7bCvh3xseVzRpdW+wdxu2ieHxDO/Wa2iCKHzHu6rfgbunQFZGjwa
S5vbysdHsjb4fiZGuKXQfwjlETNs2rDJbLFgon/rqzfOu/I3e2o9e+7Rn74ZXG3b
JkkxuS8VSBOYNzbZ8BROnJM1sNztjjJ9x709GStTIg01RS9KVMBmmxxNVy5e1f8r
dNhMnTUJvCtAYR2EwqDlffXuzf4uzadXrWU9nD3qwfZnT0/ZGnUksGd+nhINtSMC
iH7tNzpq/Tz5bN9Q8rdr7r4pQc4sajwRhvXqC03mmOI9jvjm0lSnyU1Z4JZCYf9U
HD4HcoMvRBNaZhRhpEAZpb/BwEaP+KGrRRZPPIvkyk6xJj8XHALKkZFGw3nm7uex
Z3dL82m+zGh7sWk2sbWuss8KMwF7fkTM0gl1ra6oM0Anhfuzn+viFwvDRH1jvb41
0qe6wsFuETrzr6sr82AsxQHGVVziQdJ4JtThK1Pn9g9hIW+ERgoZIGh09q1UDaCg
iXg5ERcBtCj5Qdmf3hQFsY7rGQnqce5ZlzYpzrp0rG6vQ94XhCdkYsZ98QbNl8bB
yV/UNvHpDdmLByeULRNmTZHqWH+sbORb56wnUw67qEylsL8mHBdymAEaU9MY56ee
mCSywgQKjc/F7GK8B9go1ZZe94m+2zYYmS5r9GS4W0+0GHmVznps5PhHhlAXe/8p
LnAz68uvqOcx42EuJkIOH4+BEskNB+yfXYERK+/IB/R1FQnqvtfQa9qk9TW/ERR0
NMAUFH2lh+pQEIjIM56YorjP2srk7a4oPM1pRJhEy+Lf2vs3lFsEV8vY84eZaZWA
b2jMyICjnhFYWfnpCpwWGgFjLNPm95vldF8/rKJwJs+N1RGVCyE1VdaxZ1Kn+IUd
+besJjOn0E3KOlOMwhd0ZaxjEuD8hZyklLYeRtFUhvlXFyMuFNFG8+JViwyM4clq
hPZqBZaClfviSOUmk9vs3vpFuJAlODzxolda0hc6TM5z4kdWIMai0kVykhKsRjqS
bLm9N/cjlsHbXKWyGF1prptJg+z3xaD/pI+YOxV3PX4dtNCPIYuu++2TXz58cKtu
TFgpcJ/VhzhrkYcTA6N0uZuThTKaAyCTrB+M3FnAmltc0oaeYOF1JzFgDFg9JJJs
t0AGsk2ARJnWDHTWASnlbfqYxsVLIx+7rJNL7TCfDU6M6Ecjn4p8r20VhzqwDUSZ
qoN/PfT+EvT/YMpzYhE3kpjUgg21sEs36a+oycly8TUeOAiDUTvEtb2SUjr+R9f8
EuT7lOt/zAn+dZbBNl+S9Rk2G7xXdmshj/BNzMTyT0ksEzqH8l/IpKk/OIsy6iMz
L6DFm51kzg1Xe2s0xpTBw7uhjnFbS4fLJ8DeMPDb3wrJsJRMANoFK9Kj662OXmY+
lAlZD/PyC5qAhpCZnGlDx5k8m2C21UJo9GFEkAgrm5isADGqZRqM3rA4lPnqsve1
Rqc0WPg9GNwlXeejIoYgKX7h4zNkmWqPVm8F7oWKFNv7R07z0WEJFmEiq/MCMAa1
Kyn2fP3pA10CrNDXIPpLDK9gTn26rHf1tHTovRCFNLAdJA0Q/kwKR2slrDuiIEDU
/CRpEu7Fq4ZqH7WFiOKp/rgII/+a9bGhBrlGgCBNy2JqXOxqL6S8I0LJsqyzMT8c
Ml3wM3LHRKRi4Z72zM0Xs9rmh0rW6q8uuVpUvFRvpSEBfXsC+WdQNEnCkaCY1dZG
cn4ljqSxG9dkTxnweUyUpKedFBKAHKb+XRbWv9iG6JbcZZrV+TeehFE9h+cbd6bi
UklW5GKuQEp1W1o7zwqSyY0HrQ9lJYEhrTwv9YeHVNAkww+LoOxo8wmCqtN4CajN
A4k1R9vMcqc1P3Qlip8xMYpAMmYR4Z5M86nAW9KryOvN63xlqCdMMObuB3FHGhp/
3a7F6qY6TrUO2UV6VJE1A50SkFO0oXW3C4kEvfowwrEydsfR/+qzy+HDNBrof6z1
c6mWVu45jXj313+ROMjsHmabZiTEg8rKqOdQmdnv+kPRBs4wgpz7BLrMQqoIH1bP
8IctYu9RhTQBRXyu+V35NzpuE4qDNzOK7pT/vuRGA9jfj4Fp2GG5Gtszgj+UczOI
npHZUy90YPJKZJEXBus58BxSlHeXS/stoiGDTUPcczBzAaviGDe1/eNaHiBhdEh1
iiAm4yiqNzCm6kJW/EgyLdKk3e3wCSJDHJ1M2nstWQKQ8UTkk2k2ruZx1Xoa0KEs
5Dx1ha89UspTOpAc2xeA8FUaR2fieaWRvS2CHuBvOLWCVCJ665TnO9P1AUggefk5
zONN3XfSbDn0PY6WeG7FsntKoyVC5ADaRs60xDbG2Pik7XnhMqJmou91SqKZe1aV
zKNA69JkoeMBBThjslRTkmfbYFXqg3v0Ftdj8dCDmM90fU2TU3Zc7t9iSMZo9qsI
seVIiFTIkEG4pRYkW+tLArXh1ECJ+/qu0uvnhDdFJ2Ic6ngCXFVsFsKaEgunHue1
+rV0J5czQ0e+IN/9qU6DYvtmCcCTt25BUaFvYGdYWY74qcYbWTdMl7gW3EfKQMOJ
D9BKyhihbMxPchwRKfihe3cwX+D+1mPu2+Y5JrR6r6m6Vs4qc2W3LYrpgBQicP99
dMffdMc156aF6rLg+BKNL0Ea5fHZH8c4BvOBeLAA94ln5gnY5YsExRVrvGDfg+q+
sEdM2jXRzfNxJD2hYEMWGQD3UzewnqHrVUWYQN/1/1oCq4iwzwzalViWlRh9XCXy
Cn2ePQYN3piYTqQdYo3zA4iYFiV9kNuA1NIOwLpSkkVqEcm1PRym9RnQR4OxqBnZ
oiM7TvADkXGHTsJp0pp6oCtfex/4jv7hBTNHncGhau0awVp8iekVTEKWyW085tEQ
hYQ59NjFImKahmdxu/tfQcwosCWSnxA2cMj+YaaZBLwN3+86ZKT89NQAegKtuQTU
AEJ9rZWJyjOCuXjv2AQVZ0Bpj3Hwk/vw07uC75RyRV2OZ9vKJRJP5P941IXxIiwK
5GOtu0UEjPW4v5K0+HhfiTPrScQ/L+qi75HOjnquRwluFlj7q6jUzYAhR87iEcrB
SsK2JYVkoGy6Qdr7kGDgNr09ObIPL+esCzVBeR/Iokn67PwNo9x+VigVF+T/z7MJ
cYgfu3WQ3wTQAPPOgrhRdfF53/4jVCpZZJg0qITdJSbDRxyXjfhGcOLzYx+CsLsu
wULi+iCYGT6L+dxx9il8eIgg7I1ZE1ArR0W322d0BjVG8wnlLyAaDGCRiQp6X1/4
M6xna8qKlNI+DYq751pgCXb+G9+kqNE4uIH+z+5hBr9NvORfMlizHLe9EGGptDvp
MnXYMVkVM7Zux1j5sUokvMdiYw+RjqZjVXw0a9XTplDhCI50nVYlOUO4lm/8pDhd
heXKtJKSss3OG/68FQuEGlReYt9DFxDhqT0vn0ZiLm3CiDYU3Q7I5WThZJc9Kle3
mWVYyL7aPNdvwXRcxgEyDEruEVedXro0k8zqfm3biGP6OtYP4UZXaAUg3Kymckv/
qtyQnpe9yeL1abgiie/yQEbronMiFPZfIDynvwbi2wC69ZZmz5L5RxgxCZGdfMdR
F2Wp1iMFON0m0/hp1KOsfL+4uGPdqybTlP0E4/m7vAEdMHJ6BRpwoyn1/lOKxoEi
m4uetBrhJEPIRy8BV/J5YgpGkpG9cG0x1aKtweYjcf8khKVTH0eNXfP3UEUBvPwI
xK2FFn0GqAvbwJX7nCxMeindA/A/wzQmx09IHfcKRaXzO0hqDB8ZcQQVW7yEnw6O
70uHkvglIsYzUBbO/+Nolzo8fflhEqU3YYQhSSjPfFWHLfVqz9CrzbYghfu/6n+N
YPjef2+7Zh0es6+IQBRlstwUwlRYYDtgWD0SgnvGb5TsHjKEAJfGd79qhulWC02K
TEyIDg/tFqsETMmhpBUZLcWjdclCSny53AQXHzc5dcWMXy/Mld9PNkjtwo7CNcsj
mbl7MZ0eF0FxMjHFG1A6jRHlDFq2VZycnfMswzyQorMzvsciHSo88TFWhn3SnyM6
EOyrXv4XLW0sYDM1sIM6BUlHQ6xr1h+J8fIfi/bjUeeqpVHURuS0B0MjL6LJnn68
pTBofElKeLT/x6Kl/mVaFEjuzH/BXi/nl67+7JvQ7y3IZNyVMaNC6Sopht/LeakC
WkGFVTUszslf3n3ysmV7kJQdIOn4AOJK3t+27kzesajz5/sXpsa7pyEgvxjtInhy
seCsTN/FIPwUUzmjfp9lQgQ82GEfJ/rAriiu2AQS3p9RcbGu+a51pzHGJy2bxtmR
FBDKyg9FYYQndseNCYFO8Zsd3kPsMVLIE1OFABs8j+EeEI7yFWIn8kKmF7eX0YDD
KZm9LoIs8MkORTR7l9gnYB/J/iR1skkmc4kunvcWNiEFOcVK+EKsRtw8Gcz7mCM3
E9m0z9OHIcURpX4AGDL5IXpZSKfEp3dYSySfQTbgoBhsKdUTA4vx0MPh4qMSFzN2
GLhUqWNgSAdTJyFJ3eRRU2OH84yAWrLfN24s7bSQoH7SQlz6Ffe4X8sXrb4n2Ai4
dy88XNaSC7g8iUwpWCW1JAvDQi6tEwSre23FnN3Rylh5hDQK/H4qmXRJav/pb6iH
ZgeBXdnj8hLlYvfpVsKZ58Xpmr+ScmCqiMzxfX7klzwOPR0wVq+vGAys4DGDJRrn
DR2pM1NPQ6l3Hg0bXQJQ3BGMmnv8gi7GAoTydzNMspTcSMpWN92vCgF4LMMbb0TT
o6Lgah81OBrWxoqPM44JSLXSQzJ1eef+fOA7nUyfdNoRTgG/MhZq59TTzrni+GOY
D2YOoqUmvU3egsq0S/3JlS+t6eNf1+sQORkCRbSst0A87YvmrFD/2937+sXq30TK
oeuVHxotxKo7Sq1QqC6gPxUXvAeB7cdl2ZQpUWeJwx0e4LODm0G4GsDcA37YTi5C
Aq+Um8vYW/VvqBkDp5NBlyIx+TlObNOcop5kcIUjljn1EMoIYrxnFkO5e+PmU/03
ihxZW6FFTEL2sJWqkHnMLKusmystSYa4BGPWolnEQ0MpAJesHI4EIYyYQN+m8GvT
fbGyUwDv0vqdx6Al2FvrC5EaofJ0TCn9PPWXXTAqBCEWJm/KuhhdfqvacEHK5frr
1f6k8b6k8445P4Qp+nsqrD5UzMgtpaXqVGkp8NhEpdPutQKPccVPioFgNKDwY0WC
mWapocZ4my/CYDRJkHrngwWrvDZDgANJM5qRqH0gvOw4KFlMOto6YBaL9vdPsbdV
OFQVLZU0mm5Kindfrt6IjH8C6IWcx80q0OJ/c/ouLJ3QB7TJKRDYzSARA9IaVjNo
oR4Q/gByCm8JSq+syr2wlOpd5b71Buj3xbKmigAUrGAhxWhQb29XleO8mLcYTkOb
Bxdf25qelnSn3Uac00eyYhzM5S90XP16QBk6L9VhL5V9/iy7dezZ9yYcyn8M7XxU
0MjoIWcrxsTl637Ws9c2HOV7pIEUqQFK+REoB3VgVVV0ADueo2P1ZOug8vU/ZQHT
nEyT8cehWoOC3iHeKYECr7P2/r0LJm4P9PCTtXIGCsYORYLzJYObe+k3O2gxrKA6
IFkmLX67M8DUauD8N/zll60qBACNzQZXMrumOpSwdmYbcp40jamjMDbHSjPG3s1+
hIKu4Pwv0a/bq5n7PgHaBwUYbdTZBm1KYTgnXcRCyNPYfBRy8AEym/h5FW2UrAZ8
e669YvkxbR4dMp7blXye+ftTQzTzIKV5g8De6P3IDxGIrXw3hPms7Dkae+NfJlzr
Oj0pim9oHbiKWf9L5ssUSlquChzqXYpbw4DRTwxrpzgm0MZfldqel78Ri6GW5ybj
yhjA75pzDR/0mSShLObIpZdp1fcgNp2hmtx6ZS39c13o0XnWF5CMi0U+UPHRmB5m
TpvYLtn3kKYwq3rpZqv70hM/9fcs0twXiRfx9hJTJALOAYBT4jhvUN7t5r5mCUvO
svT9L+JAFtvmrIckWite67cKZrVkQLBkUA3ZKSr9C4epytB+3uSwXg799CSnATTZ
BmKeQ6ogsRHEJ9ckMRQ+Z6d/nYll1TywGc2xKdty+6If20S8JcGiRSxM2D4dsx5d
ElapMT0P1Ux4tbPHAAgT8cXSgVX1BeeyT1NNjoe9j907Gp1GtRWE1Pa0xb+9eZT1
asyFjGlR4ECDoM52goHHXjhAwBpRB7cvMHyskKVoQnD7XPfb/lXjC8ssGBDnBMbr
rtU6Yp2r5YMGYPtl9c+2Xoq8zNbo5FKF2td0pJ3iVaWSpNssTrmPlvJIDnmUGQbQ
eTR1stWkFkosA2Civ+72WNm1062hLu1jh8BpqpuTBFjSa07+ACs2PW2dO4RmzQ0L
rHgLFapRhvhnDy4ErD4jG0AbgY71DJ3E16EYwPyJVMQN6ynBy9q4nirhEsVVFQXd
Kz9Z+g+/zWTRSrFf9RLg/shZN+FHHv7VqYhISsIRCcPJgnOyZJ9s5Flqjch94p6d
ARta5Nx61ETcmlTpaTtsZC7bZ0phPhBSNSex2YK7rOp+gm96eY5uyXUpLE6xMLwE
WrIiABOaGy6IsJxawdB6Ttv3NryvI+zjjNHAxMwlvJ2J46avRvyZGR6WuUXPyP9L
ZnvjLuNJwcrduZONl8LHPaDbj2xv+HUJYGMcMLgfrYUOyIUmgYoQZprGDh4N/Wu7
Ew86i0YAyEQ3qeRM50UXDso8ME9P5PzuqmPpP5BU+0k13P5OQ0F+6G59hk8XqoeD
mIKee97r4zdtSaRr2k4Gr5dL8mTRdALuy6kAnuYaxoDolZZtmI/Z99XC2BEaSBzU
u+Nx4973WHAGNJEG7Le566kAINntapnqaqVVQtGeEA/1VboHPZG6+LvRNEVJbMk9
Fd2ItJTXTAWSoJdY79+ElhJePc5FTLA/FNnFHhTfY/UszYMlymmcrErTJGZOHvQZ
VakeOd9ZdTMdRJRX3HJn85bezSfJ4wS7F7qFQc9Gm9VczYZriZwL7JVK9CZ+5ATI
kLW44nX8rN+IeK2LjJ7WAW8iPAkeJPyLW3l3R6J5EvcMtxwAlfE8Vh6wTwTJVQ4p
FYKxm6xHrO5rJG/kek7y052QMvfMqm6NRaixWGffZyNxbpElE9ROVMiyORcHllFY
A0rP6ICPON4psyQ+rUpf39tKnWkpaIQb8gCpeyy2rClpZ/eLtVnF5H91spuHeO9D
UYPhYHuyJs5wlwQXHeaScQpm0T7hHmKeGALPKk6V+U4+BYY6XG9cN9zvi/GStOMC
GC/ozJIC1ntRuGMxPC/ICNahhZ9mAO3/12qmVY6pQdZCnxVFaXgDSsvKCX2nPbma
ML9lTNL7ssFJi4l42nD+BKV2QtZYYjhxkRtyhZAJWTQsEo+AATdn1U7ExqIUdidL
FEjLqKMwjrHeim9mmVZeigeSNWuYmI5jdA0zodn6DG4RDSeKhrpcdvQU3Q7s2KLI
v6Cps3wf3RRv5xi7bp2zLXU/7bL4eeAVrI9bnDa5OEmt6/fE14ga8oLGRalBgBOz
GXxoVvh17CaIqWN/xG5dRMsD7JcWoF9nMtvPXxZReHnxlQSem6I9KYzuI2MNLtZA
c1A+bMX5AXzyy2LAtr+SttMoUnbcHteIOUamMvyD3dXp5nsOFHEmTbrVdc/8o3eb
/H55U9E2RYGIA/hzWlK/Ag/vFKKBBGDlTPd8MfXcO/jl0FbMNIMOtj80yJaDWI/G
RKzg7jGFj7u65GCX4GKLCLSYQ8xNTB5PjkRff9NtvOm1RGfspLAySYQXMtCGVTPi
LgRjgKgR3sybSNlnpGs9sF6jhvX2A9h2MQYvvQz9f/8gMuwJjgNa+wYD8MgJBQ+X
wDTO5QcdTxzL1EjfQeBrIcZH6Bs++VubTID7y0sdNbPXgqUPntqkqEtKibBv4uto
jsXJ7X1YoC9x+CdRNjvqY9DdCSK7Y713aICm//KK2TeUYydzBgL1jhGWKFrvlEFv
8T+i2adwO6Iq3xZf9CQITsWac4FVZL6PHtQxxNo5iOV1K98ECYmW2FOSUx1hXHLE
k/VLA1GK7SWd9BrjJUeak8mpxubb4Xs8aaumYo/Qlt8xqzpot/jefARMiLvdFom0
H15a8LTX2ES4tYA/3OnUdB1b9QaSps2FTF4VEZ2wzYsxxDMhHn0wv61QL7USZnHx
IFUfIBflLy7qE/R3GXURaKqyJVBsYVRKYZOUtppDqfl395149e9niGVemF/PQ+4y
4c1skTfFr4wP5cMZbaviTvY2FBDzpqLejSloDuL9fmDjhUNaViqZ5P6/jWA2/vEy
uY5hbrA9QCgUiPib8m8BLaidDIZZa66LsO0ScXkTV60sqCVxDenbaRQkO2HL8XbT
vSdDvg8EVSPVhjPE1gtgtHRxTSwHRyrABNY6GH6OXwwLgs9e8zZxzbUEor1iSwNg
jm4bBtdBDyAzGMkI+G+w9OF5AEzb2cEMSZuyXmXXAitluhfvuVqNXlP5wLQm34bJ
sv42JfPEJLuhP48wxgXcBQGYTD8BfUHKxj30lWORLiA9DBeS+NzEd3U1MiEK09P/
G3WCYwgX+3+4qH2XFFQKBd1dnO03PpfW2eEIqC93a40CRnhWU7bjjMrxe6ozfUbY
fTjXx1ivXfe+uRmS1f2xhw1TE72KJaA1yDx+pvWc0r3aBcPfRXFMNk3zvhpeIVwL
gs+xFuO0A3SdRomffpPnoRb85aR7DwpT+8hNkAwXRBun7Pev5ES/7CW9XcI+ATM/
UzYgAwyfAOO30lzjZW/et0ZRfFPcm8wp3633iL3CbZ92TSCrSqOfWbzmiE+IMvkS
YKcLTJVpcPueUUxqUm0dBSJru4ZVTFU63mkDP+R71WZDHXzOXLst61BojTYMTs0r
jgHgB1ycIwwsdjD99nAwxtR/cQNNL9QOO5CgAhvT0dKBuoTEYTujFECCOeQGDB+r
sT6Sq2TOsZXstW8Yrzm8RyNbifubwRqanFYfu/+2YKofUhazKISjg6SCkbr5mAgs
XQUdDzV46RnM6JAC374SE+muQ7+Sj2xCqAXl5qIyc0/+cNa1c9yUU7mBAtA6PGhK
JuS0BBjCEI7VtZbW4Yyjpr/E9W7BLO8i6odyU0wYOGx8MmdQ918Hb0bAaCmy/CqH
o3fuLrS0kd7SqoFxkBt8z23v4Nni5rux7tPGqNV7XnAMrqSBAmdyEEJPFl8sZ0gb
CwqPLOz1eYM1Dq4Ds9tiw4pF2+7dBzwjZN409BYXbmyZz3oMn/L3rdWgU+K8Xkg0
Og8Z7V7Glj5SSDlwavVsHmEkwMNf9I3IF7QOkVNKCBSAi/Gbq9OEFuvmOb6wIxUW
eu5DqoLlb8Ya/p4jsIP7OxY6xXyCF1B0ActuPg1BNTa3qmqJInOet02c3Ys2Jkkh
MFvjDsQrrZBHE6O29NGbWGQMAaw+j3SE6f0rYtDqgIgLDvj08/+c86ZJOSbFopt9
IjoI7QQlHZg22mk+TMl0coZcNm/Wch/CGzcdEzxXeqYmpxw75dT9AfZLFN49E62G
RjI5tmwJKSU5oRi0MdZZccfKBFcm7H4jeZmMCT1osNtS6ZAkrZJa6pEYrknk/B9+
2ybVkJgEl3hAgwmuWO4nEw84nbpRCIUHUCpDfojQ+HhGATSE5rC8sCPgSuwsRmMz
RRqfowLxBOldq+nXex6mwGbiNr8DQNhfjCJNgzI+2Sg7Y9SZQqVfnreXV8O/rxvX
jfiMshwo/DisUOJ8Ai7U3Sp6bfLoPxpCGp5T3jDHqN0RClN6JL+tYAYPOMgwUlLW
XxajOhLYHPG5rBAN8k2NSWWOWs7gMGq2rg1qCfMjWzNYySfO62F+MqVB1MI1JUO2
NmAM01kUGPMDbSPm038K9QIXrRTv8fF24q0i0ktECHvnkGRXUhrPK1kxtDMrllcI
LhJcUC2kE2/f5MiqhN+4/FFHv8jq/UIVpg95Qbt8W3igrXpaqWH4H+yv86xtAWaR
srez6rCklt7z18VvXja/kObp+Z5PUnRexbRrOVcRtlm+XBeLUCohjW+25ZaS7ay3
Dy7hLAN6gV/6YK5ri7mzLDUeFfOOhh/kCh3ViJHjFEIhvpppTI5FlVOIBsf67GWB
Iscdb+/1xk0YNOYdRm1FDUMNw4qpD/2a6s4X9Bl+v8u8nvPZhqkd8vkC5B86Ddw1
TluMiUI0wVvMbnKIW+K2bw5Gs9EHYrK/eqi149pxQuwu2Sjg9CQ/J5CSZbimLnBw
zSUIJz6b/K6NEDG1sDlzcVRlMHTY/Ec6IRSzeYHHz7YusmBJHo+gMvvGz8xyLlBz
hR4ZSjABo2hXFBvF052KT6txasl3umtXnNwLb3NNCLVNvT6PZgBbBo4pXPauz2dU
0T4/n8AWb7Hw3lZVCbxoUkm/a9YL9weDyIA1EunIfXf3ZRqVpkUx8nYvXcbE2bFJ
mkzC3HeIFw2G6FGu+HUNPzmqdFWtodjo5WnmkMBPfAuEFzr/BG+AyLcC1ALtjZss
RZTRFsv7Ysd3TY0RAOqIsoEuU+N7FfUvqZQcUXGAVZseCRi2bNw/k59V/DVU+HX/
97Gc8okhEJCt7LeGYcBdD7dw3OPXCLtlRJXgpHBAeiZVbljkJIo7qXdm6HxLzWde
4yTfhSC9I9r/zYRebv7M9bu0TUXUgHAzRk5mlkhBI3mXHTVazcbeKRw0UwKFzyrU
Rh1y2ACwxIztSxY1+QwSp4kWIQIXlyoLSoOuF4RBAwL/cB4SipZCqF7Aro98x135
PoIDb7yjnthChg72yY3xCr/F3OGNqixX/2BVNkIbqNlYmq1yxhxr/bROoMH6cBc9
ypmbaRvRvMbVJIgMe28j5uBc+EiFryd3L0rO+Pvx8ZCHZfoilE5x7+v513hOUZiF
3I41WdV3orykVrYmpVblr6Qli9HhjyiX72WOCCFAnx0LCXI2kbuPF1Ippjzt55W+
gyyEl3aniDgRehbOPIpY5qDkfyCCU9LPP9G4hvGVvSvFUvsdSOhCYIp+ZE6vZTx7
rfQoNALE0W9Skccj7S7/TMQ1BOsLZU/WQe6vv/4BXhDKjo3iA8XJQhMhOjiFFB2W
jyqLCR3+QwLWRhPq9cYo72e4wr+pKkRkL7gO+aJyG8ceA59D3ttgX6Nm5xFhRcpk
wRFloaUml/oJYC2HMu27vr83fkmKGGgurMbnHGSfHOanof7Bt0E9mNUe+Qbb+Pgr
Fg6bet79+i6DeO6s7+NLQ/6dk8esVJ68tSrSo9aMVvgE1nBzJvkne/GyN/TI0+or
BFz2tg7/gRA4S4/cX98tEx17ZRTMAzYsdtdQq6G9Za9Rcv2QPFZgnr0ste55hcN9
/IySsGa/8D16ox6/f5JnMWrS257L8Lr+075bP32rL8aFgBeHgy5t7upQJq6Fd5Rb
zyxEmsB76QdT6j9p0nk141mTxbMf96WGGEb5iVKfXJF6pQXs9JfU84TCFc+lW6Yk
X0SxH3JMJSzmPQEVRGvmXinvFO/fo8qEHdsXVppQLUsR2PKhYCCUHUVyRDTsO/n8
BaaQ40hmL3P6QgSK6Y6hk0bfhzE/gfONO0n4YBFp0hFKpVnqIiFmNCqwHwCfw19A
vuX/0uysWD1i+mLojn/CyG0I2kXcVP9oS+/O8J3xmoXggSNlw0YgLmN0vskrF049
LFpZPV0U1WNqZs4tg9ro2kUiRdIN0oJQDmZSu7ePq4JHUdCU5SF0j5SeDZhvU1S9
jzl0R2MXIeBegcMC+37eivaQFcwBRB1x93B7GlCmAYJD34tftHCisQxSoXpWAS1r
R4bRPNHAAjV/ntkRgPw57zGTpyj5zqh1XP1FyHdzCPoR3G43jdiSN+um8tIGlSHV
qI26ufbPUSgSfUqmF8FlEEMbDDoWquxhizC/X1DOd8O8ZNktj/9TGy/kpDGZusJA
7Dlhgrily2wjmh1Ma2ZYKFrPxMkJ08JsAPrDrXJ4FvmJJo4BWZVhSt0DeuMtRs97
c4Wp+BA9ljxb6EKapN1l91HTTMO2HNIGzSQZoKoypkkQYUU3pnNnwNG28PwkLleV
jDOlB+Lb2e0gsxurrjzQ5w8yem+IP2B265NHn1s7+WNFofoQgLfuHnA9WOOJh2Ob
97TWCegHZyyco+slLTZmTZ9E3RLlvFgwj0FxjpZaexLxBUjX9efajNl9jJNMhFsO
cKcBG171BYn/y21Iq2i0QUH4xCi8dSk75TkgayA0Ma/4lzbsWr8hR9PnC5bP+pnT
80LLhWvgjMKd/cyyV5VL0tOC8goN2y8iFGNnLJIHOi33dEBipNoknQByFHuM5Pur
d2rjSglLFOM+eijzB5dUJCS6Aes5QgntleWerLBk30ZJHi1X/6mupcQJr49lhU65
KfsWXEw/nu9ZSRDGtLFgUc9KFGLkD4oCgsMD9NCFJeBWGKm0vhpTchHMXsvaWr4k
8V1z3w8IqVhtMm03TpSLirPG+Ol+NqZ8p93IjQ0HLRyLqGRru4mXVLdsbB9OihUX
RdeaA8h54mib5rWejpIlkq6fmVkG/+ANqIVZLGZ0PCIUPWiuACRFXMDy3etqP62z
sViOIG1svuMftSPTt5KN9np1sDB3bLALtvNvlPxj6lJtIuPIKzohGtgBDpHEnLrB
oK7cFZayrI7j+ZW9w1BcPwr3UzqiJvFL6XaUJ10xGEJhl5Eo5G4/bsnDm03V/SwD
JExvSj1+iXnqwcwwNTc4HAyeVxLbQf7gpmng2nvbIdVUWGlrnqkGJX5QucBmALjv
51pyAUavAyQ1chqC7utXBgGfDxfYb72OEsoJ07DETv+86J8DMn0kxV9VkNMg6AXT
w6awqGlQ+gDQY/78+FuZzBTJhZzSiugYULKo0I7q8ALKqYAlvVI2FGnXsezVxgZS
r+YEiNjSdar1QMo7WALH/XPidUhhZgGN6m9FGrKu2ZfanXxbqjdhpJ+qi2Z0nNEk
Lmd8GuaVUf+w43G3jmzrZC8ZjbnmZ/laGXKyhHfpoxF9yclXDs9SQGjru+FzqkGy
xoAdM16EuOXv6Xyn9rSG1YyFaKGwvZysQP9IeHchCwK1jJnWge7w4Z283cLvBB5c
kJl/XMp8/bp8rmYuLbtrv6FIoFiH61xlT2vPA4t7z1uLlX9ak2+pXIbgCDzq0uM6
SJqDPqHnjx2R5JocBLhKx5kxV06BzWMcd4YX7v6heb0CnSZmSG572wR4lya6BgYQ
eYCuw6mCLpkQKV4LDyYonsdDSf646ZYODnZNhFIfopLKFKgHLJ5KicSqPlBcwt9y
Yjm2sR7LMQ2sQ8pvQEiQPO1WSBWSPCah707oAi+ehfd4GCMVCsxbiJcRqNWGYX7D
XEpL86Px0Pj5ltU6INxRQM5b5Ynz7yiqc1+mzHIevbfOM2/IhKdIwEhKYUrOCQPn
jMfZtnrgsYrYh64FHO6TYIbFlCZbHOzXcItFY6LDyZeaBFmpc44PxlcLZhzOzzUF
SFxFpMKG8QbGD7q+lPCGuih24LjVFXoTODYCVDyqfXq1k2aYpQ/zEq2BoF2Vhcsh
7mKjenBuVg2F2VRWSvslpIiZqh6xSNiLP2ORS94DHsNpjJRa81+s7KRpk0Edc4eR
jy+X7VbxTLnprpfsyS5jXsT+d3GlnWBjwAk9Oo8cmIYkmBU8N+PtA5wNVjtlN0gQ
gaN6BRZmPS8d60cCtXRQWc/MQMOeZRMoHLyMQvWo9VIcjWJqdjfKO7qClOh+aIIl
tLaclvVGEt+AAalDtIdcE2JjBns/gp7JtbbxKBc7cFSUniy2yCbJdfMTk8hXDXiO
mkb3qFK6M1pH3kwRUKtskU32PWHOQTVKsu4d99XlUGz0213oDeyP8hrXJkySa7wF
HiXRAtdELebC1lCals5H+QBkxxF9j22cQzKBG90oxuGQd5faigGPmSdI9va2tt5F
Pq4LDIy6GGzp3V9+iAESDFnR0p2BFRAREsXGlfjGLfXYC7M6xJiwXA/AWdPSn6E2
4iHsZ/XDR+BEs/QOejLuWuw+Dg7saG0AY5sIUEliuv3e9GzTOQYChM5K0vxMlmZv
RbImoGpDiQui8TGh1fSxCt63MGKkdLnlcChkCMe5pxR01uP+9rsLsdOt8dK03kWm
MFDIIXtWTy1erYpUKuZOE3ryVH302jUWFaQ4NkEMyFKOn6ISjOVJJ2G7LejqHhtb
riP0Tvfjq7FoQUBr3h/UMqcyDyIVGRI/cjlW8ZlV5mYSj+wh6JzP60+F7Z7rc8CW
J9WA3DmDea9rIJXSlDCnNp6cotlLJ3Z1k4UCk8rBX/DI653eSkyiALv7ri3NoIJr
qBiJV7c1E7OTHS8kY/bq2vqJwTdo8ieq2lhe+nJjubgONXgHw5F3Wna6GHJyovMG
+6inIJkv19sMKXU3jIGGzznZO6+biFm9I2swFcGEKEQ3hgJ1FxSSZ4HpO5AfZq1W
huObBV/0QVZODJPmU1bSosucR/SzxP4/vRBi2Wfhq8h+AIpSv+P1rKBsvlMa7A6D
YRaPF9PufcLN6wBCEqGm7HZNLVGgGAMhaB0peryShVtfxMBcKY+rxnyhnmy7km/v
g6ZKYWJorfUGufVZ1AEZxPpW9xfCBWtTFNHJTrmDkh+ME/Jc21eL15OJXJxgDwdT
3lbEEwg6Zclbr77uCzlHu4x7M2lHmmV2Q5rHUG2GvO+QIoOrSqDlk15kVuNAOdxu
CQ50irGu7KK3GAUW9bXBPRS9A/3mvV28Hr1wkRfiHc0z+h+Fw4ULZE9WjwXAQrJC
YsEwD9OodseXZHuNq1Q+krpLaM/zJrgTrIoIfrDZZqi3aMXcvx+EGXSHuplOY7qv
+PdDYRbSbmvm8vQ/0/jrLcj14C5Aq6l7DDxosY2N2w+AGaLrFBth7zqKrzySI1l0
0LVD1fP29vBkOZ7lo6pIOOY+w2gqjdm6lIoxPMCDEd1x+lZm7G0KGZk0tbVElW0q
bEf+DeeU4I9Ee2SdaUn+1kdtxhChSJWak7FaxBpFgBd0U4kDbhhq4goh2FlcrfNU
+z8iS48mq/6YdmzUmH1RIIVfrGI9Z7D3NCNAzpeNpOa+LFM51a3IylPVnAdhFNrk
t+yN2mggrtobg+CYnnacqr+EQhJy5w1Z3zVQeKwD2R+U5xpAzTAaDZ0VzWLr2peW
Mype+LNBfOpcJDVDrfUgODTmUmz1DZuj9sVU7g6QsmBv3VcDOQ8aGcXrHXYu9twm
UHrL4BYVoelWzAbjharsWd7nFq+1Y/TVNwwx4w3Du9EeNsMmVtVx93N7NC2FL6tK
PKpGISzHXP5LpupkA/KaOVioSQEFgTN8VWfABzld7MZ/2Az/GejZZLA7Okdq3bx3
6sLWpMKxnn6ePVS2O+nWDv08shtygumJiX9iuU/BjT1EtF75ibkblFm8i0L1ewqr
Bq31X8kmdCWBuQoMG4fpdVoM+mfbdqq4s4ptZXwO58/2UZB5nahs0F6dsz+0igHM
U7xmA6KuqyOB9AnFXX+O/tNaadUoq3izwqvR0tlZH8BHkJXI1/IMoIyVk2/WqC0O
+CSRMRi89YQHv43j2P+wyVQPea1A9W3vcPpwvMJHl4IUZYa7xKUSUwPGKNBesbLY
OKdOUEH7v9j4wpo3tJ/vO0Gk01ObP/ojW2ja3dGeESi2zciQfdiRmKrei3QVBtn/
V57xeJybR869tIF4MXJN6sB5L1uR+h25MAdfTLdcyhukNmwSk+0nmrif3dfnrVS6
qS07SIbjJLSOt4gN8iJw+SfB94kWpeguklmqmfRcfTl0laG4o1QoeOJdvhMIa+7N
TfBOCQfJNeF9H5MRzZJpQBjYcWgfI+IAAsn+o+N3/xee0NnlKc8GbMh8quDXmxnM
8WOYdDtSshbYyEUMS5Ro2YtdAcsQCXCJkXifDv5/Ag1F2UHTxpF4lRJpA/uHvQOs
53oVkhh+PYf3y3YTGiaayxkuTBmEcNUgGdGnDHxmUIOYB9stbTbRdKQuoTRge3yQ
yUNDDIjKIoalX/V/YsdvAaEWl6Z7jfnffSBYy3Ag39HkhlMtuBszu2gmYscxCub9
aGGxVy7fs9mW4vUtZ/5drVXzc0w0ADgVKdqi66Al5g0+jldw7eOfdhr5k6EZcJMp
QDP0l07jRsuhCfJfyzcfOx2a9+r/V4IQaxTgOLuG/Cm7vZHlXu/0GmQXGqP8FmDr
sOIpsgi37FJ9oHY/5Bo+vpHFq8ghRLxjeRGhb/yBaFrne383cS3g0LBrI3HS8kFF
nDkzwIlQqPSQhkUcOXFVI7tya6NeOKrW2CSdsViO0ekFA4M0GkRBLEeySwLOgjTC
P7HSeTZjndnyMbL3MBrGsTPTAoeTkeUSpikqTTw9HE9eWUhsngo4GHYucd/uvy9E
RIoTC0+rOCW+h4ANvs7BXXx8OGDp33M3XTf3uiaSCLxY99MfUuIvDT1ktXAd0GS1
XAMgCbVGc/asGZIIeiC9S4FlPO/DURkiXWY391YB3TG58rCnCEEyz7hG2lLVaIl/
htdwlN/aPxc1KnMFIkj1xmT4/w3/ESIHBZqc74tnLVqbVUro0DBgVAWkbvhCqC0u
j3NjxPq3K0S6ayjv1GRoFKki8Nh0Tf6WjAj84KBF7856Tifik4/E46rCS+eFfRYo
w+PxjgH/yzRlcvZCutBMMFprG00ObHvLjsOvJnKzICGV8RC/Z9WFMV4C2QcKaEy2
z0ORgqq5Vu/VMTQwN2IhMQXthMhp46uNKnJYxN246x7BcCX2+ToNsvaYwo4jzEE+
hkDmuVFl7InEi/6hDKQO8ZIuGd2/ucAkI4/73OLUGQBnDel98ZJXKtRH/nFmORp9
Biv+vQK9R9z1FF1kAuyq4LtGSdqn5uf5YQmQ7iDwHNqXJQSl90eYf5RrS3G0o6F9
PndhZC+I9M0/hT4KzchYl6xsGMMm1bWw1eJyVj+S3w9TfIGqTfmNYBewyGUDuDiv
WysCHkJWvbi3NZuQ+U0dosjXSi8i5m3OIi2L7iLpia2Y+m4BmBEjr/Hq+FasFrrt
k9joqeeLoxei0MAg7y+9pAD1FhDqIVfe7x/2Vl3YQvCZM+rpCZSJjruy5qpjzooM
1Mc/w7sEb+AsosG8MB84BZ3CLocMEIN2jHVtjK5sfBaFjERuiZF/sVpZNWYts1FC
K2VELuVkd6Cecg8/jJejiBGBCKXVGigYMErQmf9/aT1XHVSMRN6aEhqH/QXzSppO
b3hSqVOnH4prM8HZA46NcIn0bBqlavWZq/1YASjRk1o0EsFFfwhV+2478CdmgXR9
f8oLEfL6sZA1LjfMuvjPYwaVqrkPWGVAH5N38LiuCQ8pkV9cZN2fHgQmMz4VVA6H
pX9uPV2qHCQ1ceps3jnhxg2QsX90hVpnWIOPI9BgWPLOnDlnPuVZj8yrfIjoUhZR
icJxT/3d+Lf154SUhNZcS8XgrcRE4EcZnntgSYm1zgYBeV4pL5nMps8snAuf0Bps
L+jlvPjUPYfphL8zFJKBbeh3se/X+A2aX6Os75k8DVGjetiIqKASC3CN03gzikAu
KsB2WCLFK9hZuC8DcjKbD/mJwVN8Ah393N1keHQMl70evs4XDVR2G+bdt6ex/ydk
hFNMH4pcFfSW9DvIDTB7pnzeqdT92GbeF+aWEjIjUqiy5soRhXDxwQrQYl9Zykzb
J3+B/HFES1GSJ0ovpAX56sq/BoUMYP0Ml8CzBjSjVRMUxhU+Q6C901WjbXSiwcIu
UedVKyeNDeAuE6Xo3G06n8LjomC+YJ2PzS69O70M5jeQ1bYWvMZ30tRhRFx/5CAt
PMBXq5QMbbH0g3qImKCX2Je58D1oWco+1I2/hBzzJH5TurcweT23te8BalgYxazm
WtbPuT3eh5ii6+ALfvZq+M+BI2BX3ITPD6b5EzRbkPEb/PNGNqRmspnqqsOfHUWv
6n1nXtkxPgmEhE9qj3T6y9DFq/ufcYkPNw6kNPHnqoPH4t0Xvk84RvPYgZ/fgwth
Lopdp+/8MaBb8pwPNd5GJqT/1AIDUJofMCIV46MTXdGSMWkHx5reXMXFiTcnlWiu
uKxPFf8M10CTq8KqLxnX9fc3Pz3lZRzOguW7Z3iQS1KL1nEAyANMyW1RQ4EPoGiA
xlZbiyrH0g1jw3+t8IdaJum55c+hi9Re5KFYln1sb0ktj7QQB3fmsT5rRjeEplZv
ReQWbe8iMKWXSkszwMWESFHDNnMjiOkYZCIxRtJr8ArX/iAoXdD97zPLZOZSt8ms
ayhSt7VWoleaNG218V8tRmHWaPqVIx+y1+ux791Tr2PogWeaX+SAxjjjigyoETHx
nNNSeoxtP81/C8vTIJXazWtcLoujUEMq5y2KN6iUsrR2EOmrgpK+GJkKrOd0Xatk
ojYz088g/uYmhM7Njp5VnUsGKyc2F3z9nPqSFAaJcTSzGtTclJPHWzYzPYzYhvgd
/gR0tTdaB1ZA9udHmsSPMlKNoI19k1l1tHjsYMoOrzRZkQovEFEk7zw/fckGVPVt
WOBchv1aKy6Od+ZyaivlyYo2hPbk4cSgSq2zLli8gN3o5+N3cGNms+poIy2E7JG8
z2+Q4sbjz9M4skukAozyKOEoSLFGKVIQBoybFeW2gmAHU4BQeJymgY6x65NpB9Ta
5na9YeYb7dQpiOqVK85tROjiPBI0X9wisZpJmwzZ9nRK7vAKjb8cpUc3KaSwzzg0
+j2lHIERqBco8i5aI7qK+9j1pWYpN+lfDvD3bQ4x81yQaUqvgdtXW2moxYvQLMy5
hXhNZsIPB2an7Q1/YHYC5IhZakMVJ4HgfMJirsQZpTNMqJajsBIH/RZM1Mb59z2E
Sj79hMYCyiLijPHeOfoDWesLzGzBsNfAtctcP3fvVigAiMrb6ITrAYwZAk7la8hI
ocoW+PPo1Gw9xigx9q1buAIYeQwrxw3ThBCYiPavls4NWDKM91dL5jiIztNBpcs4
1FBkZfQS9knXWYjinFfcfa7tMitdsZTgrEWodr2fGvibs+kG1W1pVmRy/4ZgHZ1S
yRZx4AYuo6Sq1ISeHCGjmW5PbCX26RZut+gp4ltvb4m3I9uDFguwRqnMEZOvU/as
f1DKqS25F+5O84Z9V7Jp3hIQpkoeadqvbWf0x6JsfVxk5Y/joPPBEc2R91hvMp5c
EsQwrLqBiB0+HwUIIFtJ7+SdTUSP935fja+FODK70PJX1Kh7i39nV8B7SvTgbD8O
Uqc7zExIxbXDYq/U+OP2H15EBwB9cUQcJyNbVCT2clf6+0C4xsvfSoSubN6QDjR6
QgDIgBd+89H+TWkXyRj2NMS+thEsONYQ2i+OoKEKta8Y3RHmj96Ihl1YjfKwdFOG
rfYstL37L/JyMS9wDZtHIy7HET/LCsH5SFBVeBNvWqfnCkuynU5b37D30N4z33Uy
CbxLyA5yT0v4fEioQndFu+rieMg2vwcwe3z568b1q0CH0rJkZGKrqONzcD8pZuLZ
hBf3LssYaBYQ3xRIlJX0nhWGw+iIv+bQ696R1TuEJbEtHPGM66m1tsNEP83/H3/c
/U+HSf9nQ9kv4NNeVle/z/WvfPE8lrIJ5XC5PBxY4eKD63mecz3u82aGxXs/PV0p
EFvcJMMnqiehLCuzOAGOOGEd+ZWqDN10NJe8ZfeupAqSfQfIrWRcq/7MXj4BaQKR
pBN62a+dCR5gNy2wkGMy3A2aQ1xcmw+fDXlF34qIA+xQ1jhgvGxoGBrkzgk3C+WQ
fC2UrYRlFAUYbmm666JhB22IQE3POEYs5b8gzck0M5+TY9FIK93/nZrrb3+pzYsd
5c0fD2gYYGqOuKlDmzXL/rhMN78+NqiuJ/jBbJchmXQVkk7qGdbojbwDzGKNcTrg
vfCxEsWEyrkzPKYebQHE3oXnZosoU+f9TQMbxmtd5VM/QwBqQiiuLMtyxAYN9ujH
4eU2quUSWUOcIAiMDKtCWfcbGEnjPRf5D6l4Ax+Lvf+0u5ut5V7OO/wqJ3MQWtkZ
n8qN3TPkFbOlPYQH9o5YY3fql3agOXGdJIz9+lf+pDoj0HHVz7G1Vkm2PB5Pgy4+
Z3zxAy9nyKIJt0fs3Itr9R12slUfs7QtLsmLPgC0e0qL5GHlEy8tB+0Pn0GYdAj4
1giT/6kcMSJ6UG+/7M66oBAffN6nSKWyou1IhzMhGjOst/ZeEi3uYrSQbCHMdWon
KEZ6RBIVDRQgSrVOCwqlk+hSf26icvGzGZx9gHx3l/sZZ4mebNQvJEzcOMAsqbsq
tmDsF5laAXih+UoH/EplUBsDBhyCLuKo9UPZwP8o3XZm6qGzRdGeJzem1g1o+MxS
p+KvI5Xy5IlaEsFgMF8aNaGJQ4Uvqv6/8PoxWgJR2sKMZX7iO0iIMVUHidj7DcjH
18UeL+GGGcdqla9D2CyMyhggCmJZAyECY68LCs2KdScgRmQnr+SHh7Jw9HDU5U1W
Zw6ylW/0YmCUBRNuUYiHo6dRQqyR2A538s/ILLnWX1hoDPHk4zM7qMj5e9U4l+BF
uExsCvKmbQlMN6N/+3kcWJ594c4izVEcbYmszyrTtTWcTaVjYwCt/LnjAknXAyCH
kwTiLSycwbYtqM075RwUP6pkFwBl+EfTY+HNRk6eJs7awMb/BeX4L+G1ipO1rF2h
xPvBmbI/U4ixfChpSIzs6XzMf+QTIaYUM0cdhPAqWjirgU9J6fjKIOu/S5xsnLwz
Ccv4CbvEdKI+souaaMcOIa6sX3UV/Rv8SwMSKjeu693KGgvdA4VLg039OHGYHK7E
eMMUmSus2mPCUT6QYEsbt4rWfsRGYP/zydtkBRawIeDdzEBcsVrHtlRsDI6i+7dL
fRbkOpqNpKfhh5U2yAe1Ue7erVrrBVIy3trTXQ6RpwUamg2JnFmLl4k/VQEtvCsn
gZ5pq1+Wql9WJCKWidy6UUi3tOB0VLOg3KHSTbDvTBWFGQk6f6DHIpr2QKcHQntF
Lq6/0pRJBz50QoETNWKMjFQ3d+lwCytq01oNUfw5Gs81GV0GgyxaU/pz7Y3upygp
gQ1Rjtlk79IQRSoxdFCHk/6EnXz3pYtjaI7pBl8rwG+S6YnsSILiY2bG00F7yWIk
qZ8kcV2nJwwO4uRvL3jfNrBKiXodnB+m94wyVxRi6sh6sbddpLcLYAYWFf6UrrUB
OtAz0pF+pD5m+tM7TMHONn+gMl8dWy83xStFgDeXRQ2Kqb2tNlENxfHwy6S091Td
tS2y+GS5S7LJMPR7gmTkbNWOXJbT75n1LioZ0EF4rsyi+uYduc5glWB+hCOAmGvx
KIJ4c/um502ZDbQDj3ny4wWr6wDoSyN5Cwanjth54WrBO41cFKzhLHW0rqokcS29
5gmh6gYiABuiONnyjgbZ5aZFKSHK3MAFqarSm7R3BcExb97iB8Fi6nfder2U1BZX
sW1ksIQyOwOstAMfXxkXHQwNPtvc9pSPzCkcIPpVTeOfsgtd6fyoNsOuCK39Le8w
J0a9Tfz5eqn0l/g8O88ML+sVF54tUhkJwjQSjbiUMkGzC0ES3Cyq/Mk8F+J7cO4I
OFwlnIdFzr8L3ZbbFgV8AUfH5jMVF88Z9vhwcqpjJq5vGvdoX3cUoVQEcgGgZqaU
ze1V6P7uvb76wUwT2v7NH7mcfw/2JFFyI90dh4m/RA75SKxno6j4kZriVEFpKH+4
gD2XYpmlSyyj+1LqJZV4rAbE/22c7uDRMg/a5xDUoyT2z6DgfhDOIRIjlsAvheDS
knSH17iYdZG1iwdk9MZEg3KTiws8eilTJLwf3OOoqbnf+R7v/acbLXMIPk2EEqEw
ZNw++IFsgxpTxsGI6pzY3nT3Hkxi0aVWcmhsrZ5cn1s0EEJYYWycoLrKLg6jyaH9
w3hxardPf2rnhKRKlLVKPlcHslu0tFN+O82pl+4bwpvOOisg/PsHxybgDeekRiQ7
QYOpAHEWZEVEhzA1VR+RRLef1EWCAXm91Q2czOBAr+jBG79K4nbslYvh6fl7ZEFx
/UJeGNq/jp5BDvED8GaAXquAh6LaIizYCNEhUIbiwQMkxEqEMrrRb0OhSc6U0grR
5f2BPRnxbobcXqj0XLfgKpWjBi7RyZWKF75JgePaNhfO/yFAB/fUmTZFLU+AK0JN
N2GYRj24mAS2rzV/bZwpk8uyPKeglCuZDifyAcUDkUvyKc3/7m4LaQSc5FfKTwOG
yU0SQocepLySkeAVi8sOT6U0GMo54x4xZDkH1s6BXDVPiQxuxqUxGOrt5z3hYeGb
9VW1GWwgoxujvyLXh29xK33Ftk9F20QbInGZcppYTPWGcmoTtt3U/xs0SRdvqbKl
dzmiy58Mr63+1r48dH652UT5+8cF6QU2FbpbvwfuLrH7Ic7CzyTVi3r7XUk3ssur
R1VNC68nFph4c5JZlZCVYvbEYjfT45VVpS56ktsZ7FpT0HPyTVIcDViZQEXunglz
Sh5qmO54pRMbxrVhN3VOYdFb1+evYLkZbu/hVOX+IEe1gYl8NKSudCTm5wc1DTe/
xUCD8jtIW7BSMR+e4ViPQ7IpV9BgtiIe8Wsv+a62ZSAzR2vYiQFm+LTyKQ6VxRDz
1u+AMykunF10a3w+I335WzdjRddCJ08kvnSQnJESQAE4wMLNjSMrFv5yL6JyVLkn
6BZuY6f/1apl/+n1qYoVBm0QxVy74OF4prMf+tezOaYCscwgIdgUPDBDEBxVjnkd
+PMyNXqM59q2IahiL88IkkHS5/zsfSjsJFso+nVlGPN86SDF8LpJeDRfk8xRVxT1
0Jl/LuV9Ns+GjTCpecZnpOfwbjXBO8yt4BpFMshVL+wXt5rFImALQ7m6fciK0tC1
BuA+NjHVuguPfrp9iK1e4H1TE6i9aGhOsHQ2R0EnnVVhfp0mwc48ltksSkw0Utpy
H+y1hYN+fs4emph3R/oT2+k/duqUUZ+Efq7VHVIk4TeRxXXOLvN3mChREGMCHueH
MMFTY66zuJ4AGRoqM/eTG7s6kBCQ/KM8VQbtOcwyTAQxtuidsHnR5eEZKqWDh/jc
PdN2MN9SVLRQg5tYmioXeeKXv4afuxiK0gOjQl4vJsu9eAP2SUdm9pVjtx4sym4z
Ktf6PU/W46FbEUyMYQtdvJ/75ywOqiMzkn94QNdykE0efA3UCUINAVwFw0INE4ri
VGI0QaVNP8KCshxwVm0iaRcneMdtToVURCuPBVirFvrlYR7VWII3LZX4NNOV9J/+
YeCVrUmOWF9TpMvN1JfwsUxbY+/RqWy7XOicw8IxlJEKI4W0B7xbehg8yuuFHDXZ
mjxvjzt/DftF5xepjC+Xf9Q50r37gqgtdk6/lUNAsobxxUmO8LbVRO+9SLb7E9Ax
mI5WCFk00b6GsR9i+DV6aud3LjjRGJYWkA6MQf2CJe/PvBAyN35O3we5ddUTW4Bu
PvNol4DKnR7EakDQJdwcJnPWC1GTbIX5Kjha/jIhk6lKRhWaVfBO+A06Kxd1LBaY
qYH4aGrh+Ca1ZAl7nub6FZQwugjMCNcW9JUc+z1YnsvYfRBxsXJG0bbtZUn5N0TQ
N2DUZhX7xXGF1BjO27jvYDdSQmzIPNXingh/m4Brm2yuIXIkjhjJig7/KVYrAgHH
sbbNfZKf1jZaw7ZIVO+IaMrzmuHbx6OFAM9wfj5ND1VG9zWJ3P7WJ8LkPJ6QArQL
dyPkrdjJEjYtMbB6HuhSWsMAfpw9buzwGoOMhOJbzWl9wRry1uVL3vRres9VoXzf
N4ROuucUqQZP7eoUgUDp9yvJAPbJ/YxwYbXQBc9Fl1s5splZ68eLLSFNpAnfHGGz
MAh3q3YuLX+l6sJqlVY6AMOsLWIdtNtgpeZMI3YpZtTvpPEAYStqg6IXxl0pcZ9U
Y/ZHTlHb7xF9EIQAI4/zFB8LxB3KFcKz9En1/GkGuxk1CBYn3L8bYsXzQKd1hQgB
GECnPmKbkZioaNG9xgKSHrVkHGeuNjNo99qh19Ogg2u/1YNFdUTACKucBx3iiiWz
WralmiFj3DKlgy1GyC0QTJ3WXWdIxfYQA/lRFI4fAqQzshCSkex7KyF1EBt4ZsUo
dzLAOkZYPXINkZADDrCk4XM10KnMGYSStl+6015Q3UQhN4TmoxB2hOhQ3niGnJHJ
Mp1wI+0ODF9HLh8umlPSzWbxTuv9sls5dVcirEqj1444Yfb/t7HLnKt8jb1wZBaM
3KZA1bayoUG025FNXHNcs8jbo/vwQItFdcX2+4iGpblslQKuFv3czuGFePg4lTG0
LL1EyQwssW5CYgGt8tqONPJf3qcmsztLgBVa5l0DFmY3MJm1kK50W+hkQWElqoEz
1Zm++BRGv2Y27i+kg3mxBW/VQAI1nDe/ucuaEDnxxnYh5NX3Lvwthd3EVUtSDErQ
b4zEjRh/zIsCyBJef0num+CIO72rGmZJ00/fKpNlW810ODGlinHO3tVXVTdwJqKR
I6SrgOf5DFJUC43JRPfsWwj7SZdiuBq8PVYwNesbe7l5D3eUEXJZLUJUTUsbg9Iw
x7OYaoZ6RpuQ9kjZLeruWL+Ap5N9mbpbntQO63hRQlMMhL6fcbrBVBHBduJHEvXm
WrNODqFnHY+alrRlWwhIiehGXxknqJ1kj9UPFs6iMGtD4gJ0GKUZO0rJjMzILXH5
K3gV6jnJFK4/ASV28oKhRNIz0fQ0wMy4VCd9rp4X8khqVibGPzwjGfVnxK7UJU0H
y4kESImR4IXNXHlCRK37QydJtg6Lv5TCZm8xhQD/Ie7je91D0+aZsGc3FBRIAbTX
oq/Ls4CrX/LiCHPlK3BEK/jTg+fslRIgzbK0nQK3w7LRFMgJDge0ytrXiwSP7bl8
m66Zi9silpCSCV2j08PjYx97PDnI7DgG42raGEf8vM23P9y67ZWv9smY4sJNriLA
Ku1RYVb05ZMlWhO3zOHyjeyrPdjquvXym4nFKbRtufaG+eWQ58JHtiSFGiw9AZIh
cWpsK5Y4SOijkBW/vQ9v7YHtEpee01LuuXY3nIWeoCk9ZK1tteTaih31CAmv9U/D
4MFsmQWzAfAigMOiamKQRxFLX2uJ13ZMhQyqbDamZ0qYvPBpm/rmu6+lNeJWSY2U
TtzHBWu5cmW5quh1CJ2MYPYcQ4yV/QxfFJenvqQYpa4ywC+0FNCnnHdR0FQLHqQB
sohnRFeFYnC2nJBsZhssY0jsI3XkYJLQEdiP+EFBA4dV+9aiEbwpIf/mrZ2xSnXO
ZUxlagm2O9zyEbrboe1wwHW6WALJIJtGfUodoUpmQ+bz9JTc8cqEbVjwAwXZcmCE
148lwZcZJ5ST5FDt4CXIF1mVzyz++4olZScP4VuodWega1sclvRqoqpg9gxRRrzn
MycxkS+s55HoAQUA0N8fZi1eqNJy6KgGe/3hmufh6MNtPhvv/TJF7d8VFjQcX+y3
BjPL690p7Eq8EqM50tqkBNLsc+FROZN+ExBvzHt44zSoirIvWteon1MiOGsYyB1U
WXPpGAQ4NmQbuM39kGUMikC4z4OW/zAt1sRBC+ay3Xqxhx5U0gniP0eGsnohEsLP
Mj2TszzLzca/scBoOXXOcE58mugAzKuoF3G2JF0GS2B13LsrwemnQuwX7Q91flmx
AQ8YkmrJ5FQWa6j1BI3381cHbfw8zF1BMwScyZrvCOQy3lA8I561JgM6UBL8ELFC
j+xA9aPtZY1JTpLvqfkmzUxrZSnfxIdVEUKvL+IhnG2TOnFunq0++oONjeuBrfAZ
c2lh1Djycdq4FU4gW34KKPm2S67yOr9zXVChGfwCU1cG2fhYYYQbt04bx2SWj498
N/kOLqHQxHWWzbdLGy74ZccIioEL+hryV/eod0SifWkpr1rUi6zRpeC8mWuEJin4
Lc5l/mCAxFWQdTKuMwXLa7L7TkqYiTl59ZfJZhejVEmU7AALI3L9Y+AePDrH8HFS
S4UpaJUkF9ZnuViFlwoPJ9/ihH3ncQiQfw1BKs/yZsxAGTFEDPzNS3Kx/FlJMGvW
GZg9ZBTxAjSfrWoS4Yh0E/eZwK/NZmMP/GCoKv09SfQmZGLNYNL3YKSza+ZPKtui
RQZRQYg1o8csRzcpy4EF4Vi07sihXOs/OUqrO1W+jDzxzSYK7CuOV84r+XyL+S1O
hXim+X3TnrlPOjbaRHqG+3XsinlZaXaAabdutjbITcWGaJge5laBIGdDu9SPXGe+
laFj/mLb/B6FT58fRYoruyXGaz/l9Cmqp7CGBbdSM+2uP/gv0S+6fdTeVmU3zcax
PYUaVx4pD1Wt71KLC7R775OD2bOzG9hbua4BFVMrQVhOFFRYF/2kMITlwu2ZC4m+
jcFPo6MrDfG+XYrd+n+bBlFdHAenLjnX3dEJhGRHV/3OzzJOTCrK5ap0vwUaRu7N
OwIyf9X/OT3mrjv2AMqMJl65/gTmqGBXPVYQPPf8/T3q03bayQAfriZ6zpxKPZDp
9qgJcAw67VVIMKOF8OW/IPsk/7oBuARsX0zJoFWPE85fu3TYlxA84RYSPrWlKKbF
dVo1Pu+Iaiw2aLHK0gL9u+wO2e7GNhwZg0A6sqthhRqBf4qOIkgLcy6oyuQlDefK
ZsNeODDybNqUDmwPzcoTPlHN2ReKfGdfPeY8pZd+1tdf6qlET1a/HlZu3qPAiT9D
E7WKUo98nQa/vpPwzWEMsoRvXLHSvrMcMqF2msbP9jPH2Cogy+R+GEcJWJRoO8+5
ty7r1n8S+5y0Erh59ZP5afMS2EgE7oPHS7VE+rsUYAKeT+cMm/SVlJOU8GccInzL
Z8jJLNqBNYpQXaTeSVQxVy2XOj5g3/2qHvTklSCprBpNEsubIKxF9QfZd8TmqDMm
+NIsj8PfH9OBPBM4iqsrVEm4dPx9M9fcMRJZwzOrtjC5NEs5CFl9cNEZZm15YPhz
HGhHmX7lS77XhZE7F4zkj9EF3/hnT88Z4J/u+m3i1wQZRW8YMuNQHVCO5aq/dawm
a76B0V//PgTsLdjCww3mw8Bw/LyPyK2zmK2dZm5YIDsDIDF+3ezL9KCcVWM9DdBF
y27WmWsy3y0xDelRxYAKym4Vy9WdGQL4bu+LVlZKBS72cKYSrbIfvubytRaR36lU
NoS0wL56LcksqHyza8gTEPvQhqr+7T9xJtq0l5JcfWtVEyYsuzQTe2toQGqjHsEw
KDk3ooa4lN3fsTR55x5JP64PtmcoZVC/FMCfmumwxKoyR47YnEyG/X3JZEBctoYa
A7LOHpjyA5mDlk7E2FKvp01RJJ0QC3bMmRhqV9p4AOBIyFnbi5hl3z3lCeBU/iJd
Riy8+zWZy5BTbnoFMfZBecnagexCAIuCMn706A+dkFyWKbmkPDuzZM1acvo2cyRI
HPUtiLDkreSolR33djSSocCzshEW54WKR8RuDbMrT/RoUt7n4VDLMnOby7og62Id
U3zzOoGDLAYxANxpsgSdYZ1hSdHTFUN2oPUN+s+nMx0TAXl6xFwHlmqPAeejwwmP
aN9k13f5oUSGg2ajelbFAN2yU4g8lH42mmUdK53vhD9Jb8YgV5mQUYsX1al8OF1H
FfXA1HCXdomZ6Ox0WpgPdDgT/nzkrTv/eMgxQVXGlQ9/ISZ9jlWfyUAJO1bzu+iw
lN5dTpfbjRIvuFN3lM3JRt/xjwOlXQwzpR2QdcuuzAC0jUn1BAq722nT0ofadEu/
lgq+DdYsqHBtGL+HekdaylNO5VcplUOgW6SHBGwjncgDg0L6K7fPGm2HFpUxAxcY
gcC02bU1e3EpcwQPTFOB2YnP2WBDsSYtLnc7R91DANtfYkMGj/jTILPoVGOsvJUg
rVhsbSvyhYCeXGQP5eARp1G5ayrLaEj2SFAHjKo5tPuKB7DYYHx9KYZ2g24GQ0Vn
boSqdttnPcoIySHWZiMl7Ml80bkAK/WLHq9nELsZ2T8SJUs2ONDaJ0OLcEEhpwzs
1qU9RMbNxoaK/Ac7Hizc/aj3VeKr+RDhPGKRdMzMMb8+xXI+Bm4OmxLF4vBY2SAL
VZlFb1HaA6/c4lV1hU7b/DBbPi31LmUj8OtoIpx6RtjaIn+tvm0/MsP9sC0cG+6S
PtK25SmeGSOL+Tf2mB/F6eoFIYomsESH28RWz5csiywOrWI/b9UUWUVSkYa91NVU
CnROjITCerdLNJCJDq5mX5p6HSWY/4YnPOfCt0JxEXEYA+dPaWJ1fyOJaLVjVf2q
qoSUCKC6wX9uOj+73FF9qRzdfPX8rkoxgAFQo8tNsHdGZ1Pt3XxRfAsm3vD5MTzF
8GWcIWpS+NP90ObibHtdssl55sKqtIJPnsZN9II2DoIYwbLVcR655542gqKnF5Jy
qEpWy+0pkfO8/2DWHV7WWGcZbS1CyENU7LmfwCa2KbsmTfAJ5UJxs5A34MU5lSLo
17y5ponS5oaG31/UTrrHvWP8m6eGa6TPnIXJK7HUF6310+bbS7X/aQrY+8vdftZB
KwndjwoMMhQhgeox7e1qH6DQeznPPOqswrc2yDvoUNZ0ONBKUGJxFHJAa5rePHR4
EV/1jwM41hJ0gJ90HCW9SPsCyuhwoBDL346qsbXR5fZRSnmpdHKAo9Nxk/SD9S2o
2T0YRXI4jJJ3P/dHTzJ8eP4A+bGO8yBjs/7IdB+CJa4wdlQMQOj4simq0+M9lTDj
AYbpPIm8e9oIMkGpGssg6jqfIplX3iyl0eWt92WiHAMjVEjP20sGsb9xaMFJSOiY
+L5LWOn6FsvOioGK/yhM2nrIIvTNhfm2IGC6nQtL/Lhro0j8FIa1v1HEmgiyGQbO
+x7lgLDF/IYzy0NrC2MsF06zBme8R/A8xIdAqxxOCb8Pr0V3EDGEuvZF+wVhF6dU
dtnD2dztay+AS081jERPenm1+TgtsrcWcEq+W8eduJb93+gigHZRoOkJfr8Fa3sm
ED4M1X+7ISe8irEDWWDli8p/i/tfE5hqpXllgZ9bg9Gn3ILeQoe4uRFbQCUb5Hgy
LwwdhMj7/eWnDOlPDoEeE1GMZHCCDlVoVui0ojhycl9eMQSPwN0yXhkQEirl5rZ/
mFTgWJ6SFxIIEuETCasJ7oP/cae9CqPE7SYrYcGaxg8qHN/TX+RDggPpqpAbwEbf
fA5Nuzc7oZQIxrJp+L2NFVGhmSFxR2fpsLaaOL/WVpb7VVmY99VESSjEYw0M3bv6
h/mSBBJAfXAObq5Ek2XBW0/OF/9HaQqFeROqcqVSy/1ShGYqeakLzMUaFZ0sLITw
zvyQ9c95+lbRHUst7893zfF8kM95o133mZbL/Z1VwkPr5oJSgGo0oujx3XTLN5SU
tMxEnPPza8YI8AQcWBSfOKMUZvt2vlpuZKNF5dDSdR7r6JSbyjpJFhDAuiMno7IZ
+feruJDWO084SaLRZAbGJGB0pob302HBIbaUiV9T5JJtL7AgFo0modCXnwG6Yhqo
tRXSRbiOgfDo8R8gZAKTVUTIxwgvbAES1TluNfym4GQgQHqRpJLC8lORUEGK4mS0
T3pwgfKtF48/hJ/JfMTQBIRLIWj+YkcVqK8HatpD+NE3oR0Ibl0eAgBa4+3r0UdY
BkmAfoiPa4tTsFQ3aWFT0Q1TGuQ3A9BTOWu6sQ92z/SHaNfuwTqvS6Rv+NnuwiWG
Ku4KrNc3GCQfHKgSnhhGZJ8xKdYPOszm2vUAAeibqhk0R7LxaK4bWOsDiYPTgzir
+vgOHmphj8yqRkQEjRyRs2CAs1nYtQACKA2hUOSV8tC/FU0Af2PXCpfZAFtxZn2B
zIgfnQ3GlFYxkC3d+TY0MVrNGHEl53bayauB0p3aSqssGYqDrXlAHGKIzaoo2v4b
4mLV+7JhF6sCM5dYIWYMeGNVIsB7YP9eCbA9FT+uulKE0htOKcp+UNzfVUImdV5m
mWbdCnRri0ca/cxzt1tQFdudYHHXoCvBGt5ziMuTI56Xsm1GjtZo0Q5NeGXjN2Iv
s2FUG4WkXq5O+7AQ+acA7hf6k1eaVcnSK90hyIxyYHm6KDYEtyI11JNOUljPmwX1
2dbBl+4bEISGjjLnyPfLnJ19kzfvIKgok2WeZ+sqtgC5oGXWW/kKXWZWmDKAc6lY
UIBf/KVaCC/PvImfabm71fXe9QDwmwZcnwUPa0ou1eAHvRF8WTxkjGFmZGEXWEdY
M3ky1S/W6JVmeTH32N9DG4OBh2WTHyQVcZSPKYUBDtEyj55WO3XjrDR3nHPWJBnG
pKRpxGbvDO26H5E/FwbKyfCtUCGg7qHR0d3o4sASQObAj2H+WGgS11W0+YSi3JJ4
nLYUGdD6e0ikv3mTAC/205sZnSsU2YFS4RQtutmKfIiEbHNFxTWaTffo6tgZa+8u
qsB/aZh1MssXE0Ha4TU+r1fvTSpY7QZ5B7qFhiLNSRLj1AgBsViIf2acROLEfYHe
gba+Nd6NAOlwWcsEQRZsgaTXGac5wdB0nr5EigK20yAllSEDHILhWULDouwCuVJh
/kcxnc3i9efpIcej/yyST9O6Kig7OQqGsW6ZmCyMCGUBvDl5CbQZF12Pl/3NJOXU
igU0wwOhORSIQRUuK1CCI1WsxWv7B3DXxVpa+p2i9VIxiPzJFlFOVXPVdtvvLzEp
aEg/LmaWhsAXM8XF1w11C43LXFSkL7owaBVxypymoXQhGrv6rkVrIgf7dHE3rHe/
imrQTpVCUbU5GJbN/BZms3bJ6CYc1VOLXufP0vtTjZ+4GuK1ZZ5UxDPaL8ceCkA6
Gv78vYDlLgVjxAiWoaO/AaTYA5FZIfdeUJcWGw71BxFECZYvue6Kij9dQemp2xYU
ox5d4G75gH8PWlCV7TCnod6ImDS0vvKKoodFg8aeyroIc8h2e3VkE2lnKGS/TlaL
WgOEOTsjFuhhbhGkT7BUd7RKp/R/Gq6xV7l7d04Z1oOh0vCh5eKk7gyzZ0imJ5ar
2cq+F3nLv219B1n0mQwG40uyrowvRIs4mAA9PFgntPW+zyIyoLew5SYwPFniGZyL
+uUc3EAdWDAciOiHjCImBmWrdd9/KhX/GygMdnQ1yNt4Uug8YULNq2xpc0A0sTPf
w8YYquM/xyKDuNuqWDQqoRESf+jalTjHLh6rJ/vsfxnILKFjXUgWepgKjLqHz3lu
qVRCOmUwx6r4ayq2uIHnjXJh5fCKEoo/eN9SqQva1P9YkCZihdmLi4JmRp8OVQHM
W1YehNC26KJaATVHmR/ukVRwOWczs4EUN3llZGSbRiyMcjh4OTbah243rRdzQg4t
Y8i7pVbU1TMmHmLlXidckVryTvG5rUyUpgbbI8y6orDXqtSch3xDhR4W0HyEX3Ct
XsADYo/89Xaw0S9BIkJsLetqFUR0IV6GCNQpRnxMCpdg3gkVt9lywwshzOCrTh2X
vAlgWezB+d5xqdXR/2eIdD+mX3OkZ16RLVrwSdhpkfLs7UPD6tCbbPzOvS6qRPcQ
kRqo9wuS9TTFYpXSYnV6hJ37adnwoB2bOBuL7EAygogrAsxbP5xcXBKfzGKr6MBZ
/7VBWcswgrHaQrE3Ds+ACMd3Z3akxJ6EZ/Tn1shVZdgb7iVRqK44GXoIKMckYbt7
p1PFazWT1MS2Bg4KW5OZd+rq7M+nOrFU2I1R6A8Rpf9RVFeGDqs2P/qNsPV1lxHm
VmCBurakFPc1mN1D+chxL8T0LLiIH1hSdavDPWahAKgtBaQHzh0pS6BjPIIgNsE5
E75dTxjYdMDEfFWy15tlfQws6D/9cOLFzeVHo/D3ZEqeCfXegb+U7O0bcUJtY/hv
kI9LoRBy5UBApqHQrDU/r6HQsuYgU5X894Rk6ql18a8AiJsQyBYkBJMVzBiT5PU2
0DWNPDEFBC+pUhliWq6ll6Bv4gvIhB7msIKMAZLhbteFwlO2OFL92uZbX9Yy4M+w
qwOJsAIoRqi7DcGf5o6zfP7Rb6Gu7rm80Rv165nOQJbcMYNyJqq5iC+37dwhleNb
Bov1hMim0b+oIFnTL8ux97Fqzqs+/U6AHqO1IxwyaFP+rpwlsWpaq2F3vb+g/8iO
C2LwSQkKFtp4YVBKywN3RsoT4F5kKzDsvwTA+FLkdjNGtGdbiqZ7VgQ/HkcTOxpR
rEGm76ZfucWAW+RJU7n4lUrSrEE2aSJtaiMOcjcGkhKSzKNRfAT2wPwFjlep/zWP
mqTira3p+1FZ8z8z2YfV2nVofYmDY5mn/WRjO8WpWlzH4EuT+vXpd7i315aHgoom
TkGsik5lNGvAlwiyrZnfaIDqOF73iG2utaLqbQrUlEMzl5qo/DrKZC4OkGxbn1p8
l5nZ85FpaWbXZ3aSzRljM5Qwg77AYqh8pVnJ6oj5maIKpUSzjoSXhvve0GnEbPTW
Jj0FNjHJne7gzeb7DD/A2huj3iuXuhEmR/AY3d0x0PxbULYEnH26hmp2qMT6qgrK
vQwLTlUP7t5M8CrVlx9RduNSI36OWwJ9plsY2vlQaJDdyw+zWhA+YnwFyAryIso4
ho2D3hdILbsYP6XTZYwZXrytWV3IORxAkHF/zTfzdbyeVZJej7BxKwyhuadKz9OX
66YfLAJ86blbD59q0HDmTdJPkA0S5+25L6RvTct2+HL8TKn1Wjx1dm0YZNaQvgcU
2THwDBuDOJcnMwG+k9QmczvpAfbm6Hlt9CJxC+K/SLqT/AZ+NSUxeeV6mO4hFIzE
LIN/tbRX+jdW0RjHh64iq6A/kOpfQNd3ZKuO1z3R7/O6G3TJgAzN5nG6C6ZfVLJm
qbKIy6vevCVuNQTQmWyAt5L9xuAfWiZy90SvQwrs49157v7Q9PCsAU00N/l5Xy80
RJNxBS/bC4a8rJDS2BQAr1gF7cVkKWCqjWXcWX2Uvzhra/V854T6ICapn3AOwo5P
WqnZnAvUv/ohpjonw+2Be6NzUJ+F9SR8+jbJPhsD+Zh7vswpdpeLem3MnvrWRvP3
QG38f8R3apFu2ICg8M8qlkDq11ZzP91eJdJKImtGjmAdrnDRpt/N7lHKPb8HNiEx
uNpVet07gZQSzcHoQbtEuHkzPrvnG/bwNQ6RNyfSTKm2k71RUPqzAZhBdNQ65JF4
fcPkAES01egk+OzGcsfnAZpohhWzqSSLYhXxr03xk1aqCb5YIDba9scCGdrkCc3l
qBzLAOOeBgozfaax36TGoxdAwsTGHhHhtFpeIF339svBReTmc1jeQWI7swxBO9vM
5sbrkmsRYbmrpgIjojEgKPm1gqlV4xlXIH5Xh/dVtrkPrtyhyWQvL0rlopWLdtDL
Ljk7AyH4Po9goZc3RWdtzJVi6n0sfr1UxfQRDq5KFt9jopShhKsSjU83HINrDFyb
CVdroE+K76nMHU7+s3Reok7HZb15nM8Sf2KVtzUs1n8EOl92Q6IBw22XmlIBTNAH
wrf6N0rpJKImC4FVwxL+bmmVNzspC4yy5ihi3qCkF9x0TqRpqM+/VL8zmgfk9sUW
mkyRqWYFUIDgSQRn+YcQVCz1L5HQst/4MtUTT2iIvR7FBYh4AqGx+oQe7uzVtea8
`protect END_PROTECTED
