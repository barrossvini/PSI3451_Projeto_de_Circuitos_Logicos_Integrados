`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0lwlorsh6vypvA7R3NQR5Jjq0zL1AvQMBIfKX60T6Fv2uaVOU+nXFSUrER4a7rrP
/NQYsulXB4eNHElyaaG/lmWuwy1HRXDXYYSj1kgUo11sydn758AmUAmoblgaIBs0
JwJzbQUd3vnp+MWZoBCMZ2O9OD+d/OWZ04ABmWOXoj/nR+cdFRMQi0X1XdVPHrtD
sADutCQXob6WpfyinCHuWbTGApS6c10EdC15lAjy0f5BUTwgsQB6S7beAJU76a+4
9gAMg5i1pdFMJKuk5/S3m0MIUvNTziccZUgjdFJbVoJeKRO6cdKXXn7Kc4bMVjyD
8L5J2CwNy4dt8SWWYY6ozbVDc/rnzehkf24QAWiwKVV9lr2Dix+2Co24mvyJnHgt
WXaPEbV21s4csqA2S1uoKcoOD0t3pobtDt+O8WWVyy+aH5I+8tg5qsPRm/veYZof
weR1/fPISwEyMz7C4SjDLs9MjXrD4mobQ2PDYhMDwXJGcwtgEyID0IbMWpswlfSy
/e8BCeZcjJWCBwv8gBJhv7bK5dL9WrS8+RYrWG+I9ZoewNWByNarbiJ/2iKvkcmq
cS1BdYlkrS7lDIYHZjNHKvCaRcWYrx1ZPNgznZUnLNE=
`protect END_PROTECTED
