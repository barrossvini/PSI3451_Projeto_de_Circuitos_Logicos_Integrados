`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axjHOvmwg9y82aiw2MLskeYtBSL1P7uyJvsYEZ9Pv38SrpnZbs86o5hqSfc5BO8r
1o2NjXL6wbyB1/aaevzgENt/7z5EkE86mNx3idd5TmR/yOEAovkPAjJa41j2Ro3x
ELAcPEfp7czvMkDJhul1h63dThLg2km1yk7txjT3bK7aqbclLqBXBsog0moj13f8
ULcCR+sqrZX37uGCbgzf7J5phySGkBA1VZf6bBZMTKwIrThcsCvcpWXNzhb6o6pH
VhpD0LnJshQdWQO/jcJpgxrnlJQoVysYkTevHtwLvEJiZ1YFz1L6qtcuoIE94v5D
MSq1/azhrUzY80e8Yeac9eDhEuD6l20Ni0MXWp7OjhoqlR6BQNh8bVz2r2O2hkG3
uGpooTUFMsbIRBFrhZr8X1p2er1mIWrASuzukzHRl/q37qAb4sjycxa1KX1nrsIa
u80wPOjt0ZVeavnpLuJv5vu4Jy1JSe2xow+UjXdA8QH3KuuFX8DCoDSi01F9bR6t
afL1pVML+qHExGtElQLF/kgWzb2IE/q0kGHU6pgRrt7/9gClqFTdH58bMIybLk63
EMHNNVL/ZMAs2tOFEeQDhp7SC2mG+vOlpPDzzD+t9dvS+Z7oH64SMJmqAYxYKHdA
4buCpkmOVnKBFK4K/caEeD8eM/qSIi88i6mq/NI2EMmx5FyidaRiKCJyCBZoqkxo
j2uD1w8YVfx4UbRTHJ33Q0K0IEZv8cc2AsP1XDhOogTgeE0pRtIbX1+MVg12oTXK
/uzsx8/Chxg+RvUbyy+pW29B7mwkBi5GZ5GUOSbWsYeETV4BN+rZuxFYjk4FP93Z
nq1ggppgFoKLM0hBgf3VOQ==
`protect END_PROTECTED
