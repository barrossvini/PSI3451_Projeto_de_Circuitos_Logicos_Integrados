`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0iJ12GtD1iPAZylrxvt8XuZvnjUNJ/EYZM9RjpqFEuIDdpXwnrSIW3D3GAYUcOAq
AVA1PfSWsdL6AHQP/LOFVr9av1JdJKG0uWKKOm3ZQ1fYCpOaMizvqKnVA93980JS
hvjwMorSjKgOpcL0xPT64vacwh53YovzLq3YdVtTXI7iSqxjQLJ9eY3MOV6ZDQbe
YlU3gqi5qAIyW2pmBnVYWuBB2XEg2zMVVHI3J5AiN9N9acoEUF/T7Ud8jSdpn/qJ
hVILZzlQ0/DxfdjeZWactxkHpuZVwCHV46TVQFR3NUQq7709gFa9f/SMnCGi3GGv
txn+ljBs8sz1V0oBOREMjRA7f3NjW3Fcp1NusZpn3oWJWsKpe+eKuqZc2U8p4Ch/
yu8KqvFR7beRRJh+4VTv4AHGe35k8Vu60q43qkFBI2m4XOtJg135Zw0R3gc+h+5d
C4bkw7RXIjF/2GLqqzm0gS/mFNgW8wLIfeiWycHTisz+5gLmiMQKZpWt6oAMKqMF
kxfQpB+jeCPv++pU1OKA3bZ0R47oYjAZLqpdfii1bOgSpy2JdUIBRSREYquV7c1a
JD7QTefwAtwztPigZJ2xmcmJKodD36uRsYetfg4z4aWFTnD1CDAJTLwpfsRf2Ltq
F1xd0dvkNN3PGQuaKVj0ZkKPD3taVqCZ97+IxvF8vV8S56gsFaXPCkcm0c3hRgqg
1n86ojQQeQ7wnc5Z5RMmdc/J1pjQsVcnhoVH4wuch+0WFlp8g2Kjs9QSOniRJC2j
6jZleXkAKZ9zndz4gWyie8ANsjZvJGM1K51eJJ2Ja7Ny5mkk9shtH37fW4DnDUIS
fbtjGSV1Dp1KFBh/tnIwbKiTrBQRGuUHmsUfwIgN3AwqSUTOEQSDn4mmUVRQAeVS
8UL3vkzM5TsvTNJIFpgj1CaIoCKuHEqA/RewHdKe9e1WjMX3CNr2MH8dxAZDzlln
iBaPkqn/gjydqof0kf72N6v/241ODq2WZOfImMb1cat8zENxIDkZE5EnQtqyslC2
1NOxh3AHXfr1FxTGxqX03n9eS76FRxDVepJvaiuaCzWLcBF1SMyNP6f+ULnWJqhT
hoBt8eCzgXGlaEL7AocB2m2+yUbhblKxy+m5ONUFbnYQeFwS9a5ljiy/ApkJRTm5
Vl2jw6dI8NhBx3sFxyUFg7NUxBXWxWvU18onrbIcl+KFHQXdKm0QyPzHoIEI932E
T3+WbwXHwMvvll0CBQT+vk1oiGKkGckUU2HYkeelj7KpRj6jFiQQsMX9CVqrtg5C
2cWY26RIR/7i8kot9haN3n6PVtR4k6yqyL7fLT1lVeLGrVwCrg9VOM1LXmnc10BN
8PKNfAuPGYS6kGRrjm+RcHdUJJYuLnGHsLP3DXeSR5UEGbJDdSeV8ArdsGALY+My
PTNmk0+w4/NCi40aml6+HR6+2CfmGh5NrcuG5+x7Q/Ltirgj7TWd2Gl6CNOtzYjb
9unYPXkVhRSHnXdJ5VrSBUknrwZ89cSnV3vlldoLr87SZhjuEgUDAoC2evGQ2Ll3
oZtRvABa17oKJX4XKJAEBBOrM4XErT+3D4pxGCJiM4B0DFX1TD4OzH6dyqiAT0Om
`protect END_PROTECTED
