`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9WNsQGPRdtQ43RUY5CZg4ery3w9scuUMJzpfho6lJIX/OXK2GHJA6JdmC7+Swjsc
K0LTMq0wDUOGXk3Ce5rXPO2LhIPzfj3W363qQ1RGKV6ef1TqyMq/VqovnCyUNb8v
6cUeLfEs7xJrIgtuLn8+nBCxBqmr5BoYEzLTYVps3ooRslcy2TsARZcChdCvSuKQ
SiRoD+peOPr87RqWctXAP+PduSCsZzz9P9YUsrTFFwu4uGktJkqGTT8aVZ8vVGKA
k5yIIai4QoblHxVJ4hgazY5RtjVnsqniBLyI8aoSqTqMGyWQKIE6ubY9QZTgkBcB
GcM3odXyIAYtjMvr73w7gt+U86str/vBnhb6u+uKNl3MKp5Rx4TWV94KicoQLJCT
C8160Kfy2lfnb0wm9RF3e2xS/8guL8mFr5vZdAkXEnAuT3ODuIsFfi6dHnBFQy/H
emCD4hlzS+vfaYd68O8/fwNVYSv8dilN0s46+T1C3UNq5ogxWqqIEhdaDpdJYuAV
HE7FptxVfRM7uB/Guvb4BZVM8ET0kHG+DNIVJ6qTaIxZ/VEU5GFfMfnxXDeEz632
2KN5N9TfBLDcIfArumLWSBPW9txsIzx4+IX4+7j/TSndHBnBWFCbJt4avxK3kXyb
hS8M7kQiNqFVTbVb65jQIXJxHRxBvSOyrSSdt7z7djy/lxouWVdWwLoxwlal8w6Y
da6NyZshuusCnoEPzAjVhFRf+3HPbQ9VzruuPmyO/mc=
`protect END_PROTECTED
