`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LzsEFnIVJdyLAxHzzTdH0GAN1gtvc9d0gPrdzx1Ai6dxTLlpdQizocxbmnHtjvSk
Dckd2akW0Kxkzx52BrBj8ZUAjpkOqvvWZOLxh/Gl+xpWNG4JMPHjX58p9O7RG0C9
QA5S0tio4z90nVyRr62AQuDIDRIPrHW0risD7ZlXpgCKB/n3cl7VX9PTMNY49l3d
Nmc8AAcZXs51UMKvFGir012jyUWibG7btmB51h+ku0PKONfhuYdL34GdGbiZIGgy
NAY06jF8pErrccoORoxq4MMaqsaLa1nBYADtiw3+gILACvj5k92rMpGee9/8mdVS
oeoQVG5faTXQDklDusHR7nxvRWqh2K3KSQf29wjfI891pqVm5V5e/s15o0o+RVv2
QXitLkaw128IlBH41/DV89PoKD2hzxrflmO/3FnGIvczA8+U/+dZ8Qlvztvo+T9U
eqKY+5g39WkNyLij0jrOVZboJIu95BJMGgkLGcjn7yQKknzGgKI2ArqDNg8I0eFi
qj50Rr3FOsNGCDWzZHPm/w/xVB3jVDvm4x0g2Wq04jgJM+CyfBws57EoS6CZH4b+
vmMzr6lIDtqjcuVr39bWCksXjFLwwYAvs2pdDeVl5DlFgP33pAl/Y6SpPDmjqM4r
RbeCKvTkuufKD1Vxo9dqhzvXZ+1ZgjbzzSlwPIG5x7wP+jwW3IyEuwQ7/c3hr5mL
s3GLkI2FI6a9jExfc1oyNHNWsn9SOKlJFabAJbojU1H3z9NZrGzthCs3OtV5TM4c
br5YdSECrRg5o1WLTUy2RyMZHpQu6BThuoRb5S6LdigwARmUX1nHmdpOfuc2UhQ/
JdxGBWIHU7RTebCjJqCBaRa5Luhp2DsRR54cre/EbOCCU30fOyhHjTwXy4f6qN+i
skW7QE4mGPIRcBbHW2pTQTdZmyBsFQeXaNUn/FMU7DQy42YDbOguR5CeDqSr2k0r
M9ZSQhzA8vDkP8q2o5jTRZynYMT7qN3YQhO6fr3M3JWVU1tx4RP+LMV/hfy58YCP
3E4I7CZ/JBK8VDh/B0O4gfSeylYCLwuSi1yT/0FhZ0EKgOH9ab4nyZJkokXw+3Up
hEqA1d26n+/TRd/atXJfHOxT1eo6X83ej67R9LCWvISWj6XozpfDcQt9J/IaTuXF
dBgJpqVmtu9b0nuX2vrv6mw885KcfQ8FAsuQSnefMa9AzKbr27XbXRiqztm340TU
hSstH1IqtSRTjf476Z2p5E0g66X0sZU+DhPfLBfdaFl0GG2fZf5wqzhGpBIjCcJ/
TicFSGF9maOZ+DfeJnHIhHqXNtgArxPEzeeSafpQCgzKeV7c4qQy3ZL+P5hXv2tO
BwIdUbf/pPCFgjLTe/WStfGwFrzV+kLRLHlVEEZApwH1TSugSu2NQHE6/Uvj/Zum
q0iWfDvfTROEPupijmOVafafU3k3t5alBps6gPlDr/VR9piTXUwrb6T7kxHgr3Mi
jp/e2M2R4DzYZFFGyyzu3a9zLClONbRpHozOzqIFbna6dwYBrYjSazgL7AhttgO+
nf1GMN4LZu9DzRy8hZpnys3wnXelgSjaKNd7m7h5NZTeBta2iBopeOYN/xS0ktJv
BMo6766JCTPAkKCJkPCQ+ucYX3u7pvL9+Ziur4+wTE4cTfE+JtOnfiVkiqo076zf
2gfvXgy1sbNBDJEIdbO3P5fVU3sJpv52T741vTuXh6jSnz6P3iIIQy0LZ27/2/sH
kb79bOVdUUR6ghTdvcZwQDqA5yvmNcTGuo5fGqzWGWPADxx9ntk/ln4ji6hfzTkt
pVXBOn98nviMg0nOEr5Zu9LNL3Ij64ZjVfGE4F356s1lc0QUyvf7Z8CAw9rte1J8
LffglXP006Z0FNJeZxSSkyjaMSq13rNQpc7cRUDGsU8pGlvHnlQbJLQcp4cerCC8
SoZWayY0mywKqpUk18SSoqL3gIoouKG3cT8dFe1b3Fi80yxqdnniD71BpwFs+VJD
GubS7ZcIQETyK+7yOfaGdLkMdKLBzkNqShdW481+khUz27nGkZT8cFBZMqN78bd3
S+Yr1NoWjs8odZiHuKudbK7DHSXAW/07WYkPhPEqwJt2oIruYJtJQxguheGbeVGL
mBYxK7NdUnMW0mPXSZi3u9A3mMlZC1vWYSXKCA7Upw2+LQYbjLRU553m0C46A4wH
H9RsthXk06Kgne9FYLOURcoW3tI/lqr4pf/2uZ3InIQ3+wcN5VUGCIv3rtp1Cn7g
M91Q8HeRp7PdSr0UFEJqKnn3kNAfdiDf/DFtprqrwYTz6UHcYZl7dTiQD0UrtrOl
xOjtx9hoPUbHmAc9tOWePjnFkLExCnp5aIFx3O46RpBypiFqTURXiAH6J6cbbRdf
sFDFSq65iyP80txRjgzBrD4EFdFJ9x/XNPl1DcRvWUQTrJCyVFXpVzGRGIk0tghs
SomEXlekezVWnzjNOfD0h8ZWV96tZeftyDoentQKG6D6/JDdG9SYw5E5K/lJf+ds
9c29kL17gJzkFeIBcs2ifiSKaECchJxEVpyQQY13eDtHfHpfdYs8VR8tu+6+X/Pv
fask+fkcXKq2itqP3wiuFPE+sRXhFEWLAkT0wPzTx50jUVDZuHplzswBAEWBvhRi
7cWTU7Kt9ebGkCWcwGKYYFxVQjXi0ZlaJ3kfUcEWFAue05MLNJeTYZHlrt2wOKJD
rfLeEr8BTwfDkGmnwwbvj34oj9ihJQQh3/Jv88UFBg9lMSzxYsgM5xxIGKkV+5x2
Dk+NPnDMoiYz8QozKz8HGwcixxfVtsbNBixkcttKA9zkc3wfG7urO/varbE0KbAZ
yRfmqEutTV4R4aVi02wndjHWS33kXSl7cvYbCI8ecjS31ARgL733T7TYbv1bg1yy
Gy7Z0jBshriTUUmUsKdlW3NjYfi8X815X1l+yIM9JC2Su3wXfr6PUv4opQx7L30o
KjBYOaNtLdMSBp/v6RT3JDYmSQHdkXd3XvXZqUZoZgzwebZ1jZuF1SFlah+AzEFg
HonWESnj1MBfJ123wmIcx0G33HA41nUNRedMXRpiFksQn1UIhOTONlNeEMIUqF2s
2ykkpjph4P3lM9IFBfLfI81u51U8mJgr0e3JZs8s5/vgLp2qevjxUKMC8Uhv3oSe
NkgqYFCLCwXGT9s0RmU8TxpFalNhYKd4HFpIK4255RspGHv3nYYn2SIVE9nP8zYs
iaWWxBx68Ipt6mT3j86NL2iTG7lSCo8xhNw/PTIBsdA7nocrcUR+5L7zEiTLw4Pp
+WTh9yZYMtdRq3fwjUvbCxKLXI/oCVPIE3H/lzCCP0XAMUIKshUUMLiTw9zG5MBN
5nWRi5ivWISbNgHq+u2dQ+GqcLpCRyhtpinyzJdIgGvVKqTH4b/C41MliKK921mI
kalYCbv6I2ocB5mCuBYwiLmnkQXbcF4DEcQZaa5pK0H/7DdhUDJt5n6lz7/0/UD6
6Ubs7TIIs3MZqiP3LyICWi2UFgfNUbh4vWq2ttu/h9zsrTxvVpw1TLPoceHKmkPF
sHT+kIblP9Dxkl2/lUAFhRR/Did65mJPZcemDrOstDKPobREbdBwHXo5Hu13m+z1
m0oZl6oDtU5krzFuxECd+nALtXlDpx17cmvIQFpDcEXzLjq3OBVHiUZTPHvatXOX
7WN5XziF9jIu8LRlN+4Nrte8VmfFFYypDJLcu0fgtyVKlkS+TobWrlTYTdFmV/Kb
q6JwQzfnCuWTukDCynogteTiUpYGAY8582Mr98dJL35FSml5eKCk1j1A6EmPP60z
MoWBc2j1YV/qq7kF9CYWpTqW/cKE1tH7UzGG58vdBLcMShiUQ9td375UiCtJE+n7
oimgKOIw2GgK0N5qKc/bYJeHorarjvPRCuOz+Eg2pBjKgj+2o5QYeKRl6CTj9GOG
iYwFHXXmuq1oWScIG9LUI7GGAo//E1HaM0YM3kAGotP7hJzCsWXfrXZmaUUG5Ngk
VKyDG1MzMsD+CojChBN9EdkFq1Sm3eo5CQUkn54yPNrFHymZu73IACXP0iPi1rFs
DSSGOHbH+EfZ9WHx9FYysUI9Nkds/6KqvK8WLvjICLj/jbF8DRloiCrsgjPSCHWp
DZeSZQzqThp7yzACdYode8blC1qHsEUlmbx/Jm5QODz9d+2MfdzoHbfXSMn8dKOr
LL1BNa7a/+um3K1v1ks1aR7WQf1I9Kb8ZZDpazvMlMDiJcY/S9z8lSC8kKtaV4KZ
s3I7vZofouQCcK/HdkhX6MjPO9AnJkJivQzP+s0FwiXUwOuL0mXlh689G6TBDuoL
oaiu840mHvyj30QBXXcj42vAQgdTFCGGcUPUbFQHmTpxUmsXZdXIsh/H9+ETHaYk
90cyqsXPXIuGLzlnEOMCf2mBUqeLpKvDJFp1n/dfKZAH8TlzvKpuhCFXSZKZ3zY2
ZRFrl2aZxeasJpyTkLHqKnJl6yQUqBtlJKGN75i7/UvnHhIMPeypFrsZYkqU4scy
Or0hpnFkUI26JA3SeXQNlcmv8WZW8cabOP7VTtiuNDxCgpNDs9qHWk3SjQ/s9cLV
RD0B3y4uONZwfYcMx/byHUMNE9nuZSQ9HrmD/3YcA6mPRXAUwAQ12D1bQH2K7Rmp
EAJZ3GNlxLnJ6mEWGE4683593lSZUkHA92SXUc5xiQiQqJJa5eLF3fHTsqkZg6/+
oJkchHfsQqh6FV4e8MyM4zYWhPdqsY4R3BK+NnSwAaxhy7sQJskGIrd00lkrfRFE
lcsnxLqxSid0el1/ey8X6ZE89Idwb+DWutzgYvydAt7cybEo4qkzDLTTALiZnRwP
ZQdcz7pxdk0mxBY4UQKF7gqAPyGMGT2cxzkIbNwga8I7KffwNQEZZv+7dxe0rFtW
2erGF36eujtCX7/jUHI/OR05MllxNwGMbc8lZ1519LDPwB8WwaFHjyvt+9RHdT3+
Zi3AB+of9JWtALPYS8aMtJVgSrssaDzkXorGQiB7LFtDMfYeO7vF5Rcvrgd1Xo9T
9k9CrpCy9pDsO5o0AZZtENOb0nBFD22CDTGmTWKjt6Xhodyuv+SRS+zygGxo5I1J
F4ICoz5uk4+dchyLdrX2dZRHAqbmCzGSDIVZn8ihuVp2fuu9W/IcQq8IZSGllADT
SOa1Gg1/WyggOQWM2kBeIab1pj489IlcUVUYCwrUN8OQxCu8PODh9FctOe+Qb30E
TC+xpi2VQkU0tQ8Y40DvoYwkQVMqd947O8rtrSrCPZ5nVzIfuT+IcWZyF/jSR8iX
aAcUWFuOClNy3531cdj+a5eTWYQEacGAeBKCuJns67JbIUHuBxo/GK1ZWS8cl7Pm
owrG9ZWueMoLZGCVyZ23mbGOyRogGt4gCofG6CMgzDs6w+pTuZG0SBfWuubmniUP
+iq0xilIjFhT63rIZkXt0l2pP/64MAoRhnu+P0deIs+P4isMp3Lm/935NUMgsBD5
dCZd3thR37YUqBvWU1JinpJM2BUDimo2X5T+rF88gBkFDNcXbO2+oMoFYPh6BaO2
wh7W9PJebSKqp4NTMytXp9QQgOIsLrreRiG2mGp7DtB5TaLl1tzlXQVEzeNWLwef
amA0k6qOXWbDrwS0clXq4k1HaJqW+Gs2iDLeZU/Yv0aCVugPRkVDcCNIrz+NN6iD
E//KAJmPxqE0VqQ9KPGw3Jn4WbPtZUrgPY4cpdLq+WpFayo8hTK7CFU/yWT2iAnN
eRMhcrmUNBG4NGRgwKHEEehi4UFZXbupNLEzTXHTff5IRJwLdx+hvnNN+kyk4CxP
g7W2s8gajf1Az/ffI22blMuEM/yc/MMco6CJ84DFL50w1a0mXFXj8dOdaXnHt0dQ
qW5YzloaDjOgZVwXgTN1nKWUgEabzoC/z8V+uUdYVOYOb1sBcQ6Su8Wq0IpYxtqQ
AMqxAAs9zBzZWphrzwy3X3DzskK9nRRxoRTry1QCFQ9jIpSt9CX7mTjlWdbar/eN
qe+Fe2O9KQmr+0hCxS1Dep+yPuHLkSM/fg33U09oTtdBfUo6LPLBwk+sJprRoVtn
Zio/Qn0BeATThT+gotRyWWLQ2VIFsP8iQDGenGTSD7ix5IyHzQXw7peYQhOSLNRv
2vBh6J/m+Qy7hFa8w4sf263dAJRkGFxPnusAlRWZ11nzwFIyQbhZCd7TMf1yfJEP
jqSo5qsKXlqRcazX07LHMo0ykHhZV2GzzYKEx1LFAYPqRyDQPH3Qn5gHDuAHDKGk
8Twd1wh40mEEG/IysohSxprv33gCXmXR5Lv1DBYKmcmG1IqF6ke39fVdrPHm3+Np
5nsfeNJe+ZhmbZKS2Dw7Ic3QXjuJsHE83ZxeS73dpsAGGTJvV4Ijw7ohJ5HxpyAX
MJk8y88irqFYFU4KA4wowIOXBRiWyGXM/ZrZRH8IJGO/4qcTQDobuxQVxDPK7Jh4
qL8sTk7K8dDTjvcB0AY4oaTDBQk1SD+Ba1v/hq9zy/tUEptjPtIaNsOMo1EQ71pL
U87UuuIA7B4JYfE0uRTbUAFzabKzdmIcruei1A65qR00o8XPtn3jt7UiTXLKlQ1W
f8zztQExhBWUMrMYgtfQfHG0tWv+FVSMv7RFj2N1Lk4cGfbNCUbQLNPYnks064pm
BLz3JEkOGxRvuU9wWsLf4/qXhzagd+QV0K5AE/bT+tdOJC5qLMiHrukFOCsif156
Uezkid925odcGyPMCJ68irVW8KuooHc0dWEXo36ykUi/mf6nZhW+K+t0EC78Ug1P
GPiqXtjUxj0cWFYKmDiCwK9eZa3YirNC4LSzy2FY7Lt5o8QDHp5MPXqHuqCLCyFl
gaHAdyto750+6Tv9F1bSHQHeIGOqtREWXAQHqhs1GEERDJPlnGDLF996aNpFLeLQ
NHHbZKlxY5LBoknewBZPtc1Rl64RqFBC+De+5FAyktN+BV1HhnCR9xWpNQO4rFqf
VlLh+MWneCZyc9+OH3H0+8jUAA2gJyAWttIDxwBUWWLOfKHbGhc+UdRrTt/dFAbJ
OZHzrKOEI8upfg46m/wuEduKmYOOU7a2O5QrJ9sro6UvPfIAYRC+EITL18szwGA0
vOytntllhMa5lK9hZtnbO53ONEHPBQUBmTH0VYpjYecsP1sB5Z7HQNqbl8LPDniZ
48mCbbUqVzadUBmIXUpdbeWT5eHGbL2th9FMZjJr06Kw1iY2ewaYCWyF3lVXW41l
uwCssLe5OAPMbA6+BfZCt5M5lwJwM9YvrktZ7mNeFNx0PgoSrGECxkL2JaAj5aTk
BstfkVLfXsj4BM8GoydSHTuKwW4Azw2+Agm0e23AzK0P6MDSvZci+Dn1DFaoq2T1
wubYtgMfLhRzP4WKJEexagXJ2TGHM0FfP7hGhxjDAPCFb4/nD8HmITfx3aTR9f1n
8IAumpl1phfWr2uxr8F4eMPZr6YoQhVL/Fdznw2fps71I9D684WW+oxp+hRtsKrS
MVjn0GNcJYEPih0GvxTT5USu+JNJYQLg/QnU8DXb+BvyGBcotHETwg8PiunfolgW
x94XCLqMGESMj9rdJabH/neZ45zOy1lwPNHTAZ81FXcrfPNa3H1EVOlNI/vYQ22l
Zpcx2vOwTL5CHLRT25ooo1g5bAevYSbbVT5/s0rR5ykd4kCflqMxOnPygDt0jbmI
t2by5176Ez2klrm1c8Z1T587ObOBI1eit7Bjbd2cf3R2lyzuIrovKXFLaym2itF8
8p3MJE26Uv3pKFme5l5Qhvrt8HOWWC9Gbv4U+j43DOrjgCEJoRQv8+64Z3SWT9Qw
HbVjfPRd9rBqWXorqjCSTRQJzVCS7DM7mbWmj7wELo5jQPDXxgnDjDVr/7tyqxIJ
OCWQWnjjc1O8jZ03Hi2tt+G98Cd7n304lRzdf6EnjTG6BxEs6HXgcfehAFEpK5je
BrZTcpjlJtrQihiUxEQZq8CPSTfZ6R6+qb4txwjTQumtUCGn7v3VEugt1CfOpfPg
dIvkM3Rx9fCevchQFAgDhQT3mlzVtV/Y1cpmFjblEqrSkEx/gOKO4RhX6QljSO3n
62Box08HPv308YTqfd2WfMfIofTxdD7+3hmL8Zeg7V+PdJm2zroihHsi5MtTk5a9
kRD78HJ86Tx+Rln0+j6PrFoaXX7cQdHgA0x+hrAi95PhRv2Q+l/HPsjY20RlQbkn
ghsbOWDFbcZh8D/5kkiNZr+ctqa/urXtnGZ1K1BzHPJ/QS4Bq1XRswTNKumSo33n
WG/9WW3ai+qMFOkGYx2BrE7OXpOKkTC+gWFwxaZvIM8t/xsmLz2g/a96LisFbOmg
bdWq/R78dTEXm9HpXTuDWJ1UJHmGppc9IJV+C9i0j1w3xGb1STi8IWAODRs1nb3l
UifM+lbwLc8zwIpcI6aNou9dCEPJAX8jRRwfmMW53FThCCS7iJAHYyt6re25TUvz
JHiXkG1hg6id+XqgYc7oqF5xA9qe1OMIuZIW+vNfGTsjOpxvt0L1L4VYeXKJhCXN
cDvVTEu0WfXmbnGI39QG+Bq1O3Nnbh4bTlM6UDqc0BwxrDIGmYErtRGoFrbM+gDH
aSjtNiQKfu4tnPMHzWy5+eLhaEIl7CACvXcUicyl96w8vcGr1VPsQBbzAXgBtacC
BCwiqDNOxKLIn2Tf2XefB6hMTgfek3dLy42i57ZodI7Vq76JeDHIklZIXZ43Hr3Y
e+hf8hqBdswBGASajQUIacZCQQLJPjs9iMEUsEmBR64UX0L7+OWi3F31L8yyof97
PyR0U+wsu9CdSnIn4jppEk9j27rc9KRL3oUZ6QpKxWVnWl5tusaRZI4PH+Ol6wD/
V3LZiyLehjgof14I0bk9u2A6ncJ0JyRhh/CdA4o3SW6T+fjiILgar+GJkOw01S2d
b0c1r9YLhWSoA3te+r0H9oEncgqTF0wJYCXKYxQa5BdfTymxMYz72EUw8MMB15lW
Ml/EVs8egI8pfYrP7DAT4fgaaWXVX1yI2ixEkRHliDfJxRbNJFIoDKcjFnDVHtFg
jFRCBSSch/hVKrZgHeABDcxP+yAscTRfMY1cBpwXOEaPX+9BJZvF2p+76n6MjbBX
P5njtCWyrXFndhU8AuYl2Us2RrLhq25xJykhLwcKiB8ehrb0Ac1ntnq/QFyLDnZL
D1Nm6OI3KuspsWPMa/Bkn83MXvl11kqq8SXa0fC+Xbl3Ia+U74Dl+0uTwBV6FwPi
n+BQIbsUnpXxKJA2z4Gun3E4H0yikf4Sbm8IepY84cZl93YIbLTFM6STRia9FCpb
Z1sfCXChlQBY2ZVj0Jkkz6TyhLp+k+sCg6qVFN260RyJ1oikCFnIdbYuhWQ+hDan
LFivoWy/SejJLvbk5GzV4CLJa6R/ihmhbH49C4AmEj5XH3FemcShHJa++iMkRmfN
Dlki2SeeFbZS8fX2MHFBcQi5P17vl0fSD8i8QC1xBkzYDslC+6g9Qm8QruZ5Wb3S
Sfih7lrUy1698CJHNg3fdWxhfQeNYa9knQ3itqUzdiKhaU7xZATsuJtjn9CDxkPv
4AYdpte9y1pceEY6lFxWOeAd3oL4AxCJEKz2TJTFI4pp3SUPsP+LLIv2mJsbyQjF
v/yKjx/RwVF/i3gd0oonbRmFj65nxzs77CgshEBJHPw/0vBGSPa3vbXDwOHOOhzv
JaeOrU0h4T84OylV6TJvoWzIAjznz1RTeG9jR6hzh1zoRZqYQ+kS+MwtTiCX72P8
WGV7oz275nT/ngyjxENsTrs05wiioCiF4nfXE1G1+5Qr2onqMdt5aPQGQCb2CG2L
SwxzpN31zgR/xl0ay/xd30+H172A6h9vvG7CCQVtDwTugincGvgLLp2FLXpVgpK6
mpdJwmv5vpbcnPWFP2hV2rzG4QSQRqRta44KnHwFGcibKL4jfEtJNX/pdYKlMP3z
pKsfO0fCujBkm2Fz/7+PA6kiXBSUN0ZqK/mhyObp6OVnhbtfMSP6/9N0GKY30lzc
teVmBZAet/AB0bMBL7G2jFV9JGpj9OIdB6bFhbmQqvYy0pfRlT6Xg0SYIciT+43E
hVCznAHbp9+f3qWe/CBFas5LucTxkZORQccyhLf8AhRLXg3QmghM9rhpG2pnGQWc
Lc4PVezg1vo+9vv8a2Tc8GCpFywALrJqzGWBxdAKhGH6Kg5HfoBB4qk8AP3MLwGg
yKUr41evNZLhWs1pKme3xZjxem+/P1WiGWWiLvrcq2s3ftAQW7B+QWY+8VitWqA/
59PbU68nO1reHNSVqHtEZbIB4VePHHTsx/UXA7YybLHIA8SwGeTNatuji1FYLU9Y
JxYQf7WRsFWgRxNvVFx8nSEWe5E0Z+gkBKuLdp9sD6l2A8tkGjoGhos+ertORCey
HseozLa6r0gXiAGxMxW+5REPQFxy+Nu4GXFCXsby5jtGMgLKzF2ShbKUGEOWPhqW
7rK9B1YepZxqiQMrTaggHnPOVrN1l+gj8m5NXY2sY7SG3Jto8nmek5D/aRIywQV/
7W6uybBhau4UXsD+97OIM1kvl+Duqm/d8f/p71O2SwsKRoi5Uj6enjXEpv+sXFDt
o98vhWjz0A7HU25Wt5pdPIjHZdnGw4/XHBxpoIkw1nViWumTThXtjR1sSfvVpHjI
EgNL9bpkyIib5JFNeyLndizNkBin6z74m7p21CkJ0wIqBoHbJWgCf9a2xx9jMt5o
1Id73cM0VmZYIocsrX7/joiK8H7L4IWQv6HaQpnT8BbkzekoR2zz/2IwKQrhU1rf
3+Z0NS1gPIiR/krbJGVM3llVVl8MY3CMdYoAZfAt78fvWhbeBhT+sIAp3w9xsU0c
Od5Smh778qS4nqTVNmvfaYbr3Qs6dY0sl9G58Vw9AlW//DGJGBT8W/Z2lmG8Xosc
tr8rkp1UdVkLT1/QJmCrOjNn6rR1iMrZMNMWwM8BiOYVqaf1Olez6SsKy7cjMKjg
UIb53NnSIO+gHee0Kgm6nGGDdmZLbNOpx76bsMyD79lywMclJR9lZTTIpXH1cfQO
vC4lujBM/vyFGMK5+SfaKrAxJ1uYZIEaEypppxdlf81ULNFCsHezIJFxmfDB7ejm
LSF/sgJN3gRMJ4TmhnkCI2re+/z/d3+KXsmm+ubEN6HGt2tVf6vVoOl35yw+RaPM
J0roVTHCJc4tZxsHN2KOKI/kPvdyPr4sbVy4hhJacOIiMLgkwpfcSm+v+J3dhM4v
XELVFnaFik6f2+NndPERKk7v87U1eEdsB2f2zDiCWAN0i5AUhm8z58LphXfOK1Yr
WBGG1ngp6okCj5WS8qp1dcMNaJ2JKO8UmRsmKXA2DnnLwqeqU1pZDwKagGnPmnxa
eQfby6o7sbR/Y1tqS3dlLn3BPjlSNfp424Aqv6Ttt4OZkxdggUaw2cj8Gj95ydyP
fpHV2o2IdZUFweCJOGqCRkYWkfjIG+X+pl2tQeppX01EkTqF0Q31siaK6F10K9ze
hrSWkpbnPBbjQwXy+WU0ybolVGS1J2dUZpesKWPKVsMpxf+wh8lWdJ9XPn9luoiG
LhbX5GTs+nJfB7znWMh3trZr+hIrsFg7MrkQtv3qeC7h9nII15j2zI+cLENRbEOT
ZxsUcfJ6ss9Q+717khy5Z0ALUcvAM9teSpS0nVmv8LslpZaYtZ8duk49DbfPQMTr
pLWGqBwL+0SPexcxb0wR5XLtjm0W8Xu/i/E4REoMPuRjAxT8IsBr2rdU4CR4+WRW
/nJ/kS3UqjwE192F0z630MzhAOJ58uPZOuEhWxUNh/QKr5LA23hsKldjiTT95rfr
9eqO39a0/hEZvpr24NFe1ymjqpv5tMhy6PJ7VhcP3NvVhTuDzA6IrbY1EoTvyKM4
HDD7g8OIzTU6xHKvALIQqaGusRkDUaCY/JXu8ctPscDYZKpi5oEm1GzYkfZRvt7A
Tz+lPv3LWLt+txt6Hil9gXzh8H9w77RaN/h5FTFEEgSdwuuYrxNyJkMeVdukQ6TR
CudvUzY8PgQPHZkN6+JgLm1kpa/KFls0JGAzhWwDaOt1rnKgBR6vvpY/wAUvRKtB
bMlngPW8XVmRsbvXwF3qVwwyv4PzzuaTN1TiCOes5uNpMak0jMBDe8Qm6Ev0Q+bG
Kw1LeaGF3zb000o1qzm7I5KpcF6P6KsGt2wCqqRHXGlE2RENlyOnGoDJi3uEwtot
31rtCRENSKyldIDyFRYHhB3YOIfRDltpMeE780eBQ6VbwnPNbHPxh6aJNE/BDmZr
0SiiytJbLE8b4l/u95TIPyZbUYXNMusyshaEL95FY3OueISuOpf9pwH4uFIM9G2q
Mql+xzdE0i88NruCzDVuoLPORcg9EEYp0U+xyAIHj5+ci3GHV5d5WtyqGarWyPgG
fTkzo2bocjTr1DT+FKnkQtUeMtaQni5MZCSIHOiAHLB7eBAmGSxETWmyO/r7CYY3
7+oOtqKyFBNxfZHkj0ZsJUJEJu6auxCbOyzQj8pn3XXjCUYcrm+iaIpG/sc39hoH
gKpy6T+SvprTVMC+8M4wD0CmtDCkOeUCGBlQvuHPrh8VPtcdHvNoQba1Huk9tZ3v
nwSeLZ9IXqGyjvHDPUiD1Wu0bSCEuPdJCh8VYVoZisB8WmxqMmg2OFoZAbM7NNTF
3/9vwUNp/SP96q/l/6bD1U8/RM3lMvYnWBHje7DwTWM0GEwnnC9fQ14246+QHaUc
VJqyQ0bZUSgMWqxSgUEU2P0lEt+u5qfjiTSgGahS/JrHFeIUH4e+oKkx26vrM1AB
RKBTc5IbbG5Uu3TMAPJG9VLXibaxyLk0ci7Ma3CWn1gAF6TX0hVfj2QwRElPLHQZ
COnnlExgbp/ISTbDVSmC1D/9psCVuBSeEGBMoJCFv75A2+rkNAqZ4HoWVYoaCI4h
obFknN2DzaSFbrQkcGUefFVB5EHSwFai4kTySk+1cHfwArwdgPdCeeW9gm1XQ7sc
ZAvWIFPtN/gEW8TosrAKoBVYP99AjQYzDIIFiynda4gQ/ahWBqldW7mFrYC+0rTV
gg8ZODjWM4YMogKcB1yADuySY2o7EmtNwj4Y0SIoFVPjLusMUlnCNNgTLx9kbWPl
zeOvQUS5DMeP6jJ0q/PmPw8imQd3YkSamKTunNLMFHJB+VFEaEwJHOT8BXXuISOS
KB6/wFBXWYvu/4wna5U5rgQeS79HICF+xtiN7VV8D8b7yVp9JNHDhN6iLObUJYYF
GIjXX+SMkSmyggvpfT9TXKUk200UDRTvWjt0o9qiQZcsVMyYnqVtPoVGYUNAmhJN
NpWhAQQktK8hcgCZMWgFiGSYJ4iuSjDxIBSfL6OaGAXuI4UfnU4vjMumt0WyoTn3
WWXPIZALDpoUYYAh52GVvCLWBf93RBor8Rg27gQtqLIvH8LwFKElo2+oDouUE5yI
+Oedun3wfhbjZGRmTx9OZRW/Z0saDxkSkxw0wtSrSKuQt4871BNF/Q+c5o7epn26
26rMrJJ00+kk6b2CTlmDSrLDBJ47kgraHG+sR+Q/i/9QnrjpQafQ88DHvCoaClee
W8wJFQuvyr7nL5wVvQWF/EoBjnirRzXlfIzT24vU0pDls2Lr34y7acz4P33VYaO9
EY6CJk59yVD0CYkWXGfSWfWBCuxEgcOHtdGIiYWyCfIrwFQz6VJpL3pJY4BMucYz
zObYFHlEhEMUdIFrx53ogWXYfSwgD0MwYjsdjxabZpT6AH43AiEJyQ3ICoVGrQax
OfUSu82oED8AKohUr5jdo3xIgyWisPmTyxLNN8QPhpU2+Vh1g10TK4rU3nOWSXDH
l8sGDKvevMB7YnaR02aJLtT4JR7Lyz6+xMcjRYZMj4p6zq3KazPTDdp2c4iyvzU6
0yFz81wG30j8LCccJeZ1bDeH9oZm5BvW7IFkWiSU4h8gnQaJewD67x1LyVgWrOEa
vM8oAS4mZVzce4H6+ZOCGZ3z3UWdNGhdRPktnhhN6A5EQNLYA3kZPSNLvX0k7q2Y
geWnBbdY6t4xe1tD5FWffS9G53Q3cOJOsNLGksmUpRR72sE8+2N6qAlMVQpllXZ7
QEdsdp1YGAUIt6ftr1CMTCVwkU2d7DJHT4fzXK52zwMQ8VIb2ZDHE4J5U3iapKm1
yV0/ULOVIygDU1Yo4I77IbV1EpbCGtS+QfAPZB9cvAUTIadpXHUWNDoiTk1s+bBh
frBhVYHZa7SoS/+140nV8FH6Z4I9aq5gwjDr568u+zwWqLEfOL/TbpcjvPC8LqcB
68VDXEmIbX12oFZAeZKef0bpi56nzLbUlghcMSWIb6CLDR0sF5c2P1GmrfxowX3X
KiSfJqwaNLltbw2fLGUq2duzE3Nbp/8sYAT6xGzV+5SNPeZpifIHHnBwFewj3Tgk
g5eRP7UlxbGjEOInVWflPPbu6n4aZV9b+1rFaCVvkThU8msVfrMvdkwHnExaahw1
xoONN78G/wDB4Go+jd1BjvhB6mr2TMOTK8ePxcWC1fiFh4vNujhtJY71ec4z7hsH
YQJmvradcIjrBwafHL0O8Wm5vvi6Mo9ywULxeHmCr5NwFZrF8/Bmx+3iPglZDyKb
ic9aTCh6GhFG3BxeJT9J8bAIAwTvCeYzBXhaMWlMuYaZWMVPD1QuXQFVmdxBeqs3
A6cEuaH/U6w+w1Av340bJ1KuYeoTAMvSC+80r4XDqZjjnN9rWQZY1sCasGkYXZSL
TRK7wE6DjuQ6jed5i5RibOZE8iItX/q1wlUPAXXraXelLGlBR/0B8GF5H3d8BKD9
5z1SHL/gXWsDbaCWTwUG19rbb1Yp/0o9n9LQy7YFIRSU+tSHax4XM+2MFs1Ww9pM
9IAPpc0sXkuLFR532V0RrAGUYxDHSs2EP9BKpRvBeP3H0JBkBvBcVgQLdTKEvfzi
ahtHBqooiGZhtzr8yEApkAJd+8QAX3SBzQ7tSd0VNyAmuFXxwkMJRI2nknsHqWXP
XfH0dhy7sujv95aYr64sU6f4aIG902R3/Vq1qyg/p8etMaMEU1eVRzBEv+y8jvli
peTmqDgGJS4b2xnFK/XCqogJ+aVskcvP13fPFFlp5/zLv8ZeHMHdAwEv8alSK6l3
QSJiXf6YoBy0xqR2m/UUUW2EjbOBaoDIzRrVBcwQXzcbYEWtTEEA3I8290Wvn+Rf
Jl0s/0RekCj64ZLs2ZLYTe0mz1G97UAt8ChviCPsnJPbWbWCl7EYpzE5T7h4LpCD
bwm8i+y/mtmFNN1QsS637JID6UhSpflx+6XxBx2P127dhLVmgbzw9NzBbv/8IJSi
F6inwH92Ol26OycSftYON05QBWrBXCmEaArhpop1mZhJ6S1AaAqND/kYCJZt/WNH
+di7+MscSVzX5cA0ejHe1bPjK4isPucUBrmHfy1GvBNDigPT9mrOlG9QE3QRemt1
MgTdz6q/AjZr4Y42qAKivkNZda+RBG72unthYjA+i/YH4lGvcLfJbB2PwlCPGfFz
JzBxYJ27vA1sL6RQzcxWyBzYXR9+r3lfSSbCiRHnFmzrQGs6ZPhbFGerxgAPCYwW
kWG+mxJd9zZXony2hs4gJ8nM9VsV76kl8z+Z97NP4YUMcDot7GzuAmxze9YDDYHT
vSGgEndPU7GA1WP0IIQRebcv/D8yw6nxFUXhoGqM+lEGsX7O80+6H9rpAtDUohIW
z5VZSXLMUhOmm1TUgy133+NJJ8YEtsn5IV2VFPNQy/FnxVjPmJIZE3Au2Jv/N0Ys
OliEZE84gbDliq5/1imk7VnQXUmmTxy2aQeX92Sd+R+McNgIHXK/5pckYtRz2DUf
PXEibe8rjVVKlCVOUkr4qNHGD9anosyOn+MmJUbzAC2w1nwWAHH1fZhCu5byP8tE
F+TWLm855zyyZnOuj+nAnKyra69VuQLWpGE3Vh3BkzntutYfgduCCfU2BereeXe7
WDxhPNAhJoAHJXvw0V6cua7uOto3s0EqS4Cg1YuLofj9CjxDCdkinxWvz3N9TF4c
7hiCMop8rliiMEXrzW1TBQIdNPOTrxKAZPhpVOZu/DBwr4Mu6FOEmz8wb8jdrnIe
+wOAqhIdawSJkyRa4yQG/ver0Pkup5vZnMEO+wutYU7DKvszMSxdV82105TPxdLi
fbiVdW0XQLWcu62HdSq/i52loHj2fKoupZXcyOxYfDoQqBtuCyK7BPoXf4IbrM8x
kVbE/TqTVzpghGf/Yf5hjSlRIjdhwGzadX2CKV3L8zBjitse58404pkeeEQu/7CD
aHb9fiwH2kM74JoIVq9P8J+BcQIWQRKHpG4dikqhIbtonCC9dTDbyRovcRScREs6
+kc+Gb4VFKib/k+9MF1weiEBIg8NPoQ6YWgcuYnZxBWFnWHZ8UA0+sj5R+VO3Yin
D5BgzJCwR8aGuwM8X964lnc1HY/ndcm8tYUJmCK0GTLNNfk42zkF+P54gC/QC3b4
WuuNHWKRQGU+4UUCtbLRNiF8dxwZ4ANXyMMwhpLIhDxrtBjrtBgd/CSo18yD5W6V
kALrGmMTh8HARADqpwj8BEUPnQY4bkZenYr2HuXjuDc5/NFxRNcJCw6mNetdoS9V
UaTciywvrjOWPoZ04UgoOXiBpvfwdLNJR5HSDbnBbWwO7Yy/PzXmjm8yRSp7AE8t
riOuhBv+11q2oQdIUlA9mrOzPzmOwNrs8ytsoka8NJyjjw7J+oEoS6eSAENZk6Dx
Ik62fnybWGJBzopSgfv7bT1uVReI5gZ2WpSuJ99apCxZMPLveBa6cJ/syDVlSKP9
yYuwitBSM22hRY3M4gqxzS4WQyh09KVTrwUnt5JLpgGjOgToZTjG6bRcCt/7/u+8
O4CfkjecLDUZvJHIZ9VgqsW1nt2u9lHcD78uxGEgyhSNSRkImeXr0ey2E+BhphhJ
2Yb7oQM8fTZnkxNy2IE+XS8TAOIUm8bYdMXvuC44XVdGIZe+4Pl54R2qbqIVGFMF
DK9VX4at3BOu7NhNXgXr3KbU416w2NZqiLBcfkTD4Xk6CYbCR1g8W0soXy1gDODq
U59gWYuSiN05HuzBOzprwWTCJk7HnBfTaXsxW24d8D9PoOH2RseqyKBIQgTg0MlQ
uKgl/ibcLoIdHAgccvxhMwrKm5PeRAHoc6dziG3rE+L5W7ag30T+/RzvWtQaB+Nv
QEkWxOrn9H4rZvo4RqjGnU/14mrmtgmT2qbEnkPI6AQRAmgOIalTzrIVMMj73Ubn
rCUJtPxxKa6BIXyt+oaApwJBbalE1t8P6NRD/yojv1dRmQrjZgvdwf0kWxT6v8ED
ut8Us4LIsRyga0iVeBtJM1vjO/y/8mGsECJkQDOiXLAK9vIKyaCMVfMG/EovOjGD
0XU4PVexUaAzL06gxzRYgeJR2E61lngbaOd7xABB1okjTuwPz6BAlieS/dtsmD4s
0WugE/Hi4KG7d5pMyq1c9qkuKVD8kiCR2ymt8hXvgxDnB+sKT7jgRFP5XaELeiX+
0oc41FahYGZRIvyMD2xqMcB9CUXpNqq+LrKmkySvLK6Emaf9fwXj5M5BXFmRt2xk
T+4myWnUpiita+7Xc+K17Xz94valE8d+52hhwgtom/1Jbnwo1ePMC6U+/iXVgG+y
+oU5KHgqWh6cBrdPAw+Pyu/4KGB2vYmyjQXg3cj4l+UPpHgmwMCF+wXYRSgLCCBX
wsO2+SM/GQ2tjYTEFisMXHixg2X+g8AIZDzmGg7JC0YcJEw9bbtjEkgk5Me4gua9
plTPwfpfjlFncyA+1Pl/fSLaxEhpEm2Hvbbt0Tp9oB/ULQfyS80LPhGRI8fbO1DA
FQV3qJ3WwLu0VwWaw7JoAbffDuEUvjdFbIoDE2z87Ai/D2umfU9d+9NROb3SJase
iviHXi5zkHhBeob+hZEZLhiBrCZmPYlByOFOZ9RDJkifsM/HSlrxYG5K6lc8LCNm
By+L5BQlvhwPwUdgRiFZHMgqpFDqJEYH/GrMZgYf6P+c+u0ef24QMJCOAMMVDR5v
6A1r90zxysTsKPn1gsx0cOMxFyi3KMilUk//sRpmqzBw67SJA7zULt3lJCBDcvds
6fUi1EhAkfrI7fbYQyNf4dKd3zt4zYKf7aFpXINejZ90FyR7fhWIX2Hgki8VwAkv
bn92YvGGqb4kmebEPo1iWZeJ7mi9M1N/0v6LQHz28Rqit2r6qtSvFkZm6pB/k1eG
DEiBuY1KgrPjXdpsB3hHYctSCgC8Djki2GzOFg5kcCunfIR5H0jBtJR6q8GRbOmS
1onZIDmxgm4qiVmgV3nY7rG/NDjXCOLWBMDfBdWcYLIBd7ZRIf1gOgXXEOuy7ShU
dgksplzMJLIELy22VTLWhO25DMtBOS4WF/618smrIvx/WjLf3+dDXFZbVVEJiMcu
Eqe7JZn5u/4rnbiXuc4aPRrIW4BckBlQJST4KHFXShfZa69+FoDvqDAMOklTBVKA
+yl4z8MmCrq5zY59gT01z7L1Dr+WDErXHUVqOMC2bJPEtsnwH+PQF++kb3DpN2SJ
KhZl4FIfeqXTx025Q0ZtgcRX9HulbMhvo2kUmV6VXM6Dnu+sg7tICrOrc0OzL9z+
nMnq2OMaMDUsfeg1ddq7IdY25GUOSPwGA+Qm2gGX+qZ8XJQqYRVWvGa6qT3M1AWs
vTDQGxlgo21ELGa7Iag8+rZTdX8OrCURjal6IgcroIRmDdiWmzwGA3JDVJMHz+IY
It1/1ZubssCjWm+gL8ZpAhgG3ddRToAJEpU46WBqOntj7oNfOb0nbWYlfcfVCKXW
hNR7+Rg6ELVXOJ0f5RPNQvU7Zneu9hpI1MVm/IJyudRrSURVVt+e02rvOR7g6zw1
fTEdH/4JA8NIDthCQe7/nIxWFlBqc/Algfdc2PUlfjHJJSXL8FdcT+ep6hG9AXXu
d+qHJmFACBzWAVwlN8h4mi/5hQ7A2edbhsqVATXoupyAeQ+C+9nO99ja25Cu/eSj
pFCGf1+goa+xBKOvOWFhH2it8b88qVi+9h1zduYtqdJSdiq/5N2q6JTDjCAGPkKv
9UmcNAIF5E+mgwpLdlQRnCQQfRQGsppqFllU8CQcp6fzTPXQ7da0CI3sXuscM0k6
U+kUk1CvsR5t9fY1/dMzwEQIy4QNrIomd2Hl3wnxjbSUP1LN4o5A1MeVwAv+aL++
QbRN4kONjga7Yzd46GQZH9wujiPV8PUdcjaioXK9h/uZPf/R37ebVci3AoBigxWV
h/2tXZ0rRmlJZ7eaONTPPTeG5jqH9NmqvSHD+4VVG7M2yhAet86cw8NwaTSZW75q
d60UjhO2Quh53sLSMgai9ciPK98SkV7+o2kqMbwWgdn+kXxzOcg6G2pr5L+Zh92F
2rNrP1CTXcGjN+QyNFyiIftD0fu7MbTBkiTIQMSJ5xrqhF0G1i0M51l15RTPk6jq
RNyUClOE0VKNsUshw1oikmdJ/24C8+QlgGbr/6PC3ryHHkMmcSpErRGuauq0twtN
Z1gYEW7iinvsPc8MILFn7g63l3c2bjT06IUlPuI76diZ+N4eln61HQp5DOD+h5Tz
kkkTaDtT2W5nYRi/hZ50TCr8EheMfSVCCBoWcs9my71u22Mum7yP+001HiO4J3Sw
8qjJFpfXefAnJly3yLyJMtEd4DrrUbGkXBqDMwwDNKxUJ97N4NnZEwQxqGLVUWK4
MrjOouDPlGvMCCYROuGlsO3U9jwQF0fulQnPCYvedOQRn+nFTTjkYUNrkjgmAddG
Z98fY+99VfK4iXI1DDC77eC0vJeOmutNIZLS1yCoEA32qR64v4jIrRkVzP8wb8LQ
3Hi9+losqYihu8rR1ll539DxBqerq3ACjow3zRjQ88C+r+le9/SqSmzALXLannKY
RObUon9oAws0gz5CGl13ygES2phczPKtW3jAxiY3wAnlh+6MWgvuCAhS9DGbDHO2
gObIoqfhiwL4jn16JhOoU1QZgzLEP6zVANqwbH6SA97FIQYsTEG7JQEofi3MxbAh
a56dp7hFKLsI4Hg+8NlyqowJcKviFSWjV0gP0kY6jNW1bmMpVJacoz0C3sE93eUe
p1hjQbsPWMLD7auXadJ73uPqDpRxCzx/8f+2glAAnHGH6COAvLEQ9aZquVnwi+8B
+xwmzQz8n3pV2IQ0JulyD9pvlZ14rFIEbXG6ZmXopk8E7UPnj1myIxxJX7YDKagX
JQKwrSGRbhtkW1pIGl/JgrKp+kKw+lHFUeutNl1lom/M3IkZYh9KneZ2yIRyZ60t
LcnlT09Rw1bzWH1DwaSoVnsD3WfOM7+0hW+p3/GvJywn7G0CvLZMW6WA5wfO8Q6t
unBLJ0z7Vj6Lqlcrb3PoEs9jtdpKgFeGt+2mqs3MpP6y+M9x/HtCc9+Com0VS5ZV
ptcw4EwnjWXzWm5uLcyuTlC1RVmMjp+sf3vlrROJG59U0zMwYfpTjPmhlSst9+Li
5kozVAghX1KxCfkFoRfOoTtN4Wrc2xyFnbb+shQmYVC6bIrauGlvoRDv31rbl5/p
f8+B3oUIXBHWN6gmBbnk1pmUnftMQkpkEwca9CqQLJPbNThez1GPA/Gm7sy+GfeR
YbWAvoC79FOLh3/zK0+RZbh7zTpWyIpCQnxh2/KQNLtLCmHgPbPhmVQjQqMe4SEZ
wegjNycfgt18EIliAmVgVCgmEgEMr2bcjP4z8Vzi335dILJ5snlIuSMemR/+lNoj
a8jsXa0MWa0zENFQTVlIkQCfggrRFnga9tPZKoUNaIRduEHwBMUEQKqEXPeS2Bvz
oxpZ8+2v/QVDw8+BsXA07fWh8z73quzKJ9NJqAqS1xUgfeEqxq76pDanf8frZ6Cs
7FckhW+D2OvzgnQGrRdCPOeMedXGekAi3sPI10roswvLMyfMmp0HTUZxAZyCewm1
O7RJ57GWPOKAZsTPOCMxqcGDJVabEG4dzSY38b8X37tb8VTGG7FxD94BYKztgkB/
huYTs5Hp3/vwl/tNQHrUrShIwsp/CL24F9xZA4hRMLClKNMRuoBBK+NqN8Qfvd13
2ozDRSUW6MsI23Bcl+RVtDakWyUgd8PTV+NF6HtLc8pWJi1X5QgbfpxGl1DsCl/1
II1Yb1s/LPZ27diwdnR1yyQI2p+K1FUsXZ9ksNbPYlZgIT8a7R8CuFZeLMDmc1Io
VluNyW3bpBx9hjnG1kSWs7o9BGzdJWKNU0Hw//yAIYONY3mXBdW092/40vSx2pe4
w/Pu/fI+yFNgynbRvZDiXXzs+6Ch60pZjY4GyaZF2x+zCdmujGAxkEaIygxr+Cb4
zFRpqip16QHsGuiVM/m0stDX+C31iMVS8Xf/aGPc7L+pIzvi0ZobFu1YwR6RUMvr
uwV7WMGQQgjKRlXC0y8x465pZUwAHjgdI/3XVDEw6XwnR7BcNPfTT+nGTlQ+h7IR
siLrws9WdDJ57/kL3u7Rvq9JYbVrtdAdOdTK1toFE0xUPvDb5rsV6vRIGXNeVYQm
T37XsK9Y5Hw5v0mxRHp429DcS5RdfWQ4uQPHJqQfzyBp3Mv3hWZGt+p6zyOYCp2l
rFLxzrIXWPaHQJ9klnWhR6VbifqBmHYQfVeeVh66kFuJq5JfcG4HoOkIbR23hLfC
Z0yLk9hB2COqKKPnSMtBIazzxJHWl28G02ls0QzB8/7botlBwCLlwZF+UNESo+xu
Erbkv8NUUZTQF7SmLh1zGiBNN/ft5PfH4qgLQ/gRJv+qSWofsF+1Xvx1HphoCuP6
zTlxKkGmX/NOfkxhb82b9UqSrMdpiYH5or5qfNqlVELxb5ufL6RN9P5uljE0ncbj
EIfbkUFsGiEgSh8PuZZpd0ezM5ma/8uD+q/NPZ1oeGsmP7cRQHvb9sqNObkbxFgi
jjxBOcHH0la+LzJvhUm/g3HRWm8g2dE2IxOd5U1hMkUctBsbapplweeNXE538mq8
hUMIBDO6JBat8JzNs/lvbaL8ZkcRHalEV2V9YuEXhJdEvs+ZjgCLiZdZ3j4xVek+
QJ/R5ODV34zlOueKd1eXiHXJPeQO3r2znnk1+pk/A84i9O81ciDX9pCSB7Kbb3xi
zZ5MMfNbzud6v1umpFi9oPaddMktR9HBRiJcFLm8j0T0EQLhXpwvWAIhJDPPrP48
PPK/I2MHupjCHVakqndoMrCKiRE00tC75raL1mM+8AWrf577unVf7cW883Z9aYqT
SAenPrBj3hI8c1UMf5vbXTA9uEdEPG3zo8xGTF+30/u1uLEbo9rU1/wUyhHCOrvC
Z0N1QqZ04PqbVtq+soFID7WVLWytReUD7a/3YiKrvLIsRHaCBpUfsovW3GmipZ5O
uyrLGPnIJy0FDAA3qc1t+ahDUJj1Sn76kX9ZI8ALOdxPQJndoffrjiiVLrQg+xVD
wi4Lf39k6cQ4JxTpr3DnWwvZuIq7r3Jc899TT2gJnHWYM9PfpLjfL2YzZqzFY8Jp
7fwcn/2wDPfbIU/wiVZQx7Yyadsd1kwfeD03EWilILzy3uWURiNnkQhD7guQQmxd
o22WlljpaUxq+LdHFpvrgcXdkWIevzB9zLj+Nyfpj7EYP+xplhubQ8t7X+/KJzqN
rxHtwOCa0cv6XfXtU5z0C6k+KJ926q92kKAdrFOBP4HOQNVgwPi3m4L51qv1wEOV
uwcnAPigKgdA5nFFqUIUOfJNf6XCLTj6U3EQj0yOCCAFQZBACaey3Mquct+NU2v0
/K2cNWbR0PXX0TSBtUtytYN3SiIFxWkWoftnY7kYv6OioJUzmA34vnAgnBTwW9fa
p2q1zCUCThdjwmiQ5/aRLXPhWDVLNhdwE5PXQ/oICVus35eAMIiCjTVNAnP1/ts/
GZ2LKLdtfMLwt2oZihyr0pNRW66Uqdq3MyOilYVGMwZpuilnHjvlPYHip/NXpmei
Zhw/f3pu3yED6otJEfdJLOz/KjeJqKAwZ0N862RIPLtR4lhCjJaOyknql3Z++TO2
tUqlgAUmVmt3GmRF7JtLoOuusp2758ic4cfGsZmr0HIaLrxCUDb0k/oC7OjTccxz
aIqN6tljhJ6gdUPmogHfjUZMoZbXr65W0Z2fwwNUhYgVWcCpdBb3dbbLSWXy9kww
xcEONk1rw5WuyGqZi255I3tbBXMvGSsE/kgeO32lUIiXrS1u0HH/A/xzEqaw4VVF
re+Bfs48Q2tKXABKWBy4c8uG521/6rEOLQBkknEc8IYNQeOM5zbYsyd5EDVqQSlA
n5Rjd7xk90TbwoavtkEWKtQY/CBsFBolMajAhbYKrsmcRKolcYyNVQpw1aC5TKYz
tPV8raWCcABQ7rUfMNob0Z6cj46b8gOFp1DJEpR/7L9Q3tdgXteYoMZB12WCho1G
6PX0URBGeDEHdn1peOyoxJU/SWPDC1QpyKrjYTVef+sdv+PR7kT7Pa9LW+fmlQ2O
hT6sTO5Xc6/v9TTnJAUsL9lRMkWQIG+YPNmUsN217yw6rCJaMJvPSHXqhnrrkVpw
0Eo8P57NQuyhb5IfFIxy/c7L8eIc29kWW/ih2mjp/WGPzUWXWEk/OAcrG7XlbwrH
bYwykhCk0EATDsWrSBVyaxF1UtcSmZSVum5yg+JPsQ1dIu8NhvcFlCvuOQEku1+g
Y/JuD6ZZ4QiUpoN5hsWULC0DiNSuxu2luHDdt4n8a4iLCGWwZImt/Z2/EZHhbvs4
AL6iHX1w5rhermRO0+atgxgaT2F2pWvuVGCGR+CGek2pUT1wk9g91N+qkEOu2ajj
p8HpJLCAch6ak5dOWoEeQsA8wqTJ1oJlHGpWoXliObqu78DyM3B3W+D+DwWwX9py
h+EGe3cKVtMDfMKuwVKTDe1/W01Dv9BsmR5wX3DHeGb6chEl8KSHgV9f2j1yArsB
RAW/AkKuV5KV82LqDjJ9bDKCPeU0X9TEJN7oUSb9HhlU8UBqncmVGoM6tR+o1OKD
0H2kd7kyAdnPkw/FDvt+LcS2QLGq5sdZrLyr4btlGXWOWgU7yjw7AmaKBgxN7U8n
4/NnTXstNCi4ixU3aQoRFs66eEN3HZqPuO1T5l4B7Dr7ZdnjT/a9zWpMU3qMbyF1
RCjM0fm5r8xEoekd55FsJQavgWVtQmWVbUvM8mnH9XO+sKoxw2EPVutYMW/GUKpK
Mer1RHt66/KqEHk9QprBJa5wloKkaJWdvsb/bi3fLFQaQlc9rfS1+ypyVJgZN/rm
CnjhfYo2wp6q8EiGXi2SM9SC5BCdv8orLMbSqMRAPmMNKyigDnP7JhuhdOkxXKKL
XgKbP3Z5RW10hyTBCK4ExDsUrwc8hK6DcBpYeJoBmZY25pdyL1MMJjEQqk7+X+8a
Kwa+BhUdpIAPdHoYuPxxVflYRl1U183xS/oRhi5RMNXtkbNnIrKqnlkLwdO63Yi2
CuzThhyXM08IO1aTXh5jOm+qIlNEFPwsuar7Glm1AZ25LUSFS70NTWQN9bd+eD+g
lTn8QkcOuj3mfkNKl5va2F1BCfcYzS6posISQiGqQCStdmGw2EENN9kYmhoRfZrj
bpeo1j1y5uTm3oUkNwcoJCw+BNPHsi8R37XJtKNtVXKviwox0ojD3wzHvJgYtD9S
H0ZJYil14D9ncu2ooB7FLhhxo2+0B7oCUs+qmk/K5bT1OzhE2xpYtdlEOH1ua0xe
NXKKBC32Ciy17QqPmmiHp5+Lb0NUFeg5Lgx7vPgaS8z9kN2qKWO0r/CT8tFyRm+N
x+Sx0aymiCYgwOviRkC44QyRHq+W21FB0VRX21y+CZAbX+a5XQ9jPIh89FqWO9QA
IC420u8HqrGODH/WwhbvYD5grM0IJrlOVdtPUBcRPuR8AUs8MmWVxw9Tp+6bnBDC
g2XrHdf525QE21FGmpQgVQB0cPtg3wJD5OEaCbVI/BpKWYgcmHHs+r52S5cpIMHs
Z6MZ6ShfSavGcdYjG4yP9q4VmJ0cIX0IXQkWUwCyt+XxlMag8Ro00lhbZJFkaRQq
9U7M0JuJYAfFp53+jijgY1iGflpLbEAbTKC9Dk3k0aWRmiGrthwkqBVE5kGJUMiY
pHVmd4m93TkfZEd5rCIy3i1CaPNOTqs+mOMIRFBRpyi9plhI4QzYrILUq+OwQige
lifm3gN3j7lrNI/VZwWzcbOqm3PGlXLlKpleidF3zBVk/dCOPA62kdfU+AUDQsUb
iQ7gXUY2WZNxOfe4hOovP0wIYTo4n2oXnx493OHo8M8adkAadz8yaFTnoglLDHNS
aHEly69UZYcUwusewYsusb+r68BCiixfOCQonSBfP+vWBdsMITejdhSsEQA9DIAY
gU/QoL79ugGK1sMxxqA6JYenuDe5wLEdg8mH2k3HISPkIUHZ3fJ8DrQnMzZOBrtc
Z96Vho77eEOlgVQyxyC9oxLOu6K5i37SCKLXRYN2gfxXF9whrU6rUBA5bdQNr1wg
rfjXcIfGYyRVKtsemxLuGVRCIBdoqxxiZrgkY0jUJ1WGScIkzRJYfY2LSn1cA5bQ
eLhynqdkhE9BgvhPo1AYpOVqdC+z736Bz7j1gK0YYVlgB6BOvl/E4iK9oids5eUe
3YntWfsEHw3RmWIqSsT9X1EtOu4PqehOHDaCrMUlYDxRm161qsw3zNlnG3mYhbnt
druHPgwNIGgroMfBOg+J5SsImC5CQcD0ZdTpWA2WEpk/MGZx8cRxx4K0HnKRw8kP
qex4ZywtgZJi/53UwPblzG76SCT9tL+fNasKcnymUhHa/pJ787vP9VKB+qxh428T
GtoMcX6UML+FH87DSGnSMWIW8Rx5deg7MnhwtfdaDP0n2GGewsPCbwl91u9koeIN
0CqqRoptt3+6P+Xdb2fHvKInFVIHA6VIPZZ6N8JDUqCqL32elT2jskHQngXTvKd4
OnmFQh6MLgjWJG3cTVf7K3m9Is0IuB6O5DoyepOaIFB8K4ZTy+x1O6ulaLo+NB/i
vVaR//3WhFr/f8NKBO5ZZEElHq1NJo1BZGK4J0W6DU55kwzzeKTUPMjvx4l0aaJV
f3McqDBh5L0y62ceKKYGmVbFff8nUdi3N7piJfZpfld++IpiVIe6saqOS0ADfOYq
4WMRcvFb0YC6+wQ8vYQ+/lUuNRXaDso6zNWmIJZsNI/ZoKkFy4Fy7F8VOHNtgBiO
i2hZXTu7zyZOj3xdYhGdqPDzXFzgldzmKhBV+HXy3Juh1lwRTiXKk62U3b5ypEkS
mn22GhKrdv0Lbe4RbWCxpcxJYBmiph4I9Rknjv5Y9APsyGXEHJhsnXKNbPIJID3M
GIrB5SDkb1RDyCR8zCGrT5AHOqttICr8+Ldl9E1+I5Pn2RZA+/d4Bl5E8LQwMU1d
xC+uGUColikgYEOvCv2xmgpsk1JTYWU/+uTpuNT/8HYfMXLhtoRo/B/cwMnwbdoZ
OI4aBNnWDTfYu6RT544s8LEyA5IT1LpdMl7QbLrMC6AtZVWi+pk7yzyontzJDMhw
9+FqewZ4BHDqQ4KVKHCPavYFHk0Q7X/qYY68z/rmDDcJ9G4+9DUrRmbOqyBw0wOC
T/WcBUv0Q7lPVOS2cy7ickmnS7Azmv1Jtju3pnmlQ37klG36vB/mDDvVShrha6gl
gCkXcOGdgpdXxKvvTrp1eQgakpozE+vbgRb+OTO/MuhsgO1/osbnIU5G7C00EsMh
gVLRLakZDqCw4MwdSv0nWeCYhupLQ+68mOhUIlSIYFleEtNWCay1kT58isgdI1E8
KfpjeLTFNVzFslmlulM1UEA/fActRF4Kyl6ouwPV70hLPZCeKBML7+DZSFvfrr91
V3aUAZXf65h+xSBrMLv8WsZFVbYJ8GcLRD8d2oxHByxZf85UqOvnCDeqK8JMA9m9
4F2DQix5N5QSwf1y3M82dp5qWcsA2IVuTO0aabDgodK+/XjpGcao8G+8jcxp5tHJ
W1gYvPlb3hJj17XjW8Ke6CFAM3tQaytpwu/NPAxMRxLfZXeO0D/KgZ5wRzp1ExN2
EImyH3tDOZaElhB8zn/OV4qMU57jGpvMHbiSetRWOd+QIVEjoEwYs4+uR4e6w/GA
zRpBbwdp/sYCdxudcV+02IgzwbFvql0gMbGs77YS/prlJMNKt+u4PX5c+WDjQ4p3
T9J7lg4QC+fIHiqgfKYQsAqnNc2PT0cMPt272VzhoYbZ5Dn6QquyvGhyxxochYPS
fVz89AoL4W7aUO5eUALKhdRWq5k484efm9Kw3K2MnS6LbdfwvZigbakP203MpqTI
FsW/J7LdJ8eIxRGOibZdF5Ee5JLrwNLZP+JUB2H0KnbmPY2Dw79uFBSqJDxSNLf0
tRdquGovqxB3kNxWUrjvtFjS6mrs/dPHK1O2n7wCNk6AuDJCeFVtijxPxuUa1iR4
1cGUzebU3MEannRvwak1btCPdL7DZ9ddeEhK0BynbBtTC4FAW1BwPvZjVgKhFJnN
eiCq5R/edg1u3OChEOiA4+pcjecYMTo+T552MHnJCdrJDVP1hxCH7tUKXqTR+7LI
FR1jBizuz7IJ0QlfJVyeY2nk3jtR8AVS5X1PQ2A8D+I316+7aU/2J5HIOhlK3aZt
yMomooIpg6wrET8ll+lBYdyGv4I1n6B46gnbkmuz3SDg6cQNXw7K+ObI8GC9M5bI
rRH6mZsWusaDCmmzXTs5AZ7NDM7TKpGU4UJFOEuX0mrRK6OHnYUsYi2oPzJcE96r
OPatxDDTYXj8pSPvRSbX0mWUoPZlA6R4ASasZvISw18AuAKRt4cqGTYhoOrZi3Lb
a0dXYBV2yhdyLViN8Z1uSN0jdwKIVVOP+ojelql4EUq9jG2NNpdTiX3UWxRsU3LW
sivEIJk9zlEgUjTcNv4pxnnGnAIUFBfCe+JTnBaXRxnv3kYaMY0aySufDSpm0pXi
14xCj6xxOuzN65dhyFM1pWEYorcwDQGYfFhvjpMdNufT78o+LGVbHkXSr1JTFhVA
+DK2ivRKnyBXYkgciL6ZWqE88RQ7llB5NfJDRziDQ7GE5jUxwxomeKNegF4868XI
t+1ZN8aoH+m0Ba10twfE1RHXa9GdGftlDEYfTFSa2CnaVYNEI+poDlOBOp29ifjY
zUJdaD+zuP82HCQALX0KCwLEo2npNo7mMPyaamCZaHe/2tTPvFAAmjLq8QLKALEW
HHLVYiKFZoafJ7Q/lN0drzaT/CRUD+ZVnqRsiXGC3brps6TP6xUstS6dLkn36UJY
MiQzooma4rS2bxaWZB6PcnJDg7Y4imqrCEMZzTvFOk8pe0c3Myd9uIuPVGsbv37f
n4wY+sVEUdHFt3TfQ/6MTBVMZWCrhgsqppoMGFkKVz31q7106swatsFNHhMntQfx
EPdIlmgTReW2/OceD1CiKY5fs3eAswCpE15ZihvNak0DX/ZJAUV6cxXHazX+rPwr
Ra76k+7QVUbs9k2fEMGN9dL3cjSxqj+A9X7yw23sQGuqCJgX/bS2RkP1c293Upzm
CS/CF7cy230QJV5C6C2pvYT8Gh4x4jEN9Qeu5FBTscsgVh1rNI7XWkAatLLRX6Qw
vY7woMjLorp8Q61XYBFvkfzjvmmby2QGWdTjpmqFqw9vguqcSava696Zk+/24P8T
RhuqVeo96e+7em+qu1qI7WjZx8YQikJO76Feki4I7/tnmIivyBBZ0T9aDV1vjSq6
MljFOP5Z6OUJ4zl+MXDU3Gf1bBTEDM/hBFj1KAMmsSAxykpSKU3LRUVYBdsa3Y5P
7137DSu+5u3xK5BC1ZgQaR3IO4rH4YYi0SKZ+tEEJOjdZidKlVq5IwFDNdNeVYCK
iEhAPdUjcKRyOJDirMnaZGyNS27787gVkan8RdXzhpPoSjQ0gQJ3stOWy37L+yrb
IPoEb9DZX1KrWbqtVHikBoY19eB6DYbK7MLCqBZ4ZGIuCvyblhJpJk+mD24W1gO9
OlD4hPlChrx5JbsYLZyTGrLk/8L+O7S2VlmYlf4MuzRqalHLVis89uIO/wtbReqZ
fwFlg7m7+1lYVgIEdS5IOGML2g+iEGFcd+euyv+IePQfp6QkmWKk9VIZSnHsBKbP
KDfM8gwshaGlBqhd5Ipy9CUj3iaGIeO+rwt41T7oq5g2ro1ftdHXECJ7VRX4JmHu
bJQ6d18W+33fxdv7cMUNM/XFwdvvSx9izVRvLsxqJEM4Qs0S0YOOPIR2SbERRO3+
W/IvC0KGlITHB+NhWTW183m11PgPtxWAz59e7b/K72uttvyOPCjF1q1zN7xqoBxr
Smn7m+G7wnl5Vy/dhtR0iZBRqy2iOrPJj2URuyK8jzp5fHfLqsSP/Ht9MfJ+ue3N
NqlUgShS/gJswd/x3MycXz57DuFzrTwpWnE10l2yrMXcjhOJIxR3e6mlE+5467HD
vhFUsPTKl1gqlRm7Rsp5E8F4y2b+uVW3uviIIjo0mg42HSwkWHJJT6Kt/J8fIkvd
kJReoE+GuAUtsttJPXwODPeON+rknvTEH2XzjmT9KBB/HNodyLt0/qql3VsiNCXM
zn7e7GBz1igAIifHqMeJiYr2tYQzhqfTqm55Rwh6zRNOgbMD05UEdZVsM/Tdc7zP
LnRnR//3BC9TJc24j6A2B+l3gZkK2cV8faPg53oJZZ+AL/yWxhlaHD7cDAAyBSl8
gqQrgxYC84eInXz7GWdMCgLoAEtyD/ph/1nblP3zA5vTF3omDGlkF7gUKzrP8gPh
mkMnTOPgBDxW9oM5DCQEI0/5cOIOJOQMw5IBIOl58OpBL4zNsXgbkskx3LNGqm6+
65gKTxTQisCp0d+Mw9fq0TBsXz+dRJv15M4kFJKHX9ydVIg+nNYblYxe8IsTmua+
1u+ialV5AIxtf1yCMfT+Bf9wtk38EH2iYyQiE/u2mqTh6brzslt3wrOpANthXiEL
vUtJ5O0CJrVqgsO2yBNkfHJ3/FI7eC6qrA7u0xsydtfLr4qMlZQ+obPxl+pDQJHd
DweX5S19DuFJA8M8seRoZzImcuGmup9upm1wvVM684ut+ZThZLaXTEPDBdLBOi2a
Im5MzyPC++pXMH5fkYMDK+/JseK+AYEkFRuArAQZnhWY/+DIz2eIqfoNt3ktRONv
Nwo4YV+/+jIyHiM1g4tZ5ZjaGm1FgwIC52uFZM5YdbjRn4b5qHAm0KEvBRMpD2WO
5eq3lewhQ2VMlE2h2N5gfrvqFVMAZNCsvloxoFZC2SqZzxVUW7SrxRIXeYfqjbRW
uPKnDzDeD745xmx0a9Hr0uVMJ542cqvYED7gLyLB8Eb//RQZjJNy6W5yNkn9P4Vg
dZris3Dm8Zn4EjCUN0Axa+IFK7VU4llbFKlmvorYQYdbI0j0J4rh1YFVFSdctYFU
gbPkn929ujJ+L6S7v9lvlMgu5dTPftQ8/obziEq8hFPO58+ymVw+vvZsy62chYYQ
J3uRn2w6hmHDLI0YDlr/HWaSatOdrqNc4mJRsMtolK5LrKjCwIxEVqEYh3ATz3z+
5n9IwI9U0Ttleiiog7lu4IymMl+T49Mg7HLhFcKTvmP0W3X2pfXHYaY9AtxscDwI
efpW4umTpFTU05tuAjMKpb0VOhEiO06wQf7RAAXUwlwSzsAQ5hoTNyeg6uXVJuK9
qCME5EFg6hyHYOJck/vVx7smLgRHUs8+BN8bH2JS9feIad9AJ0xtLv52bRW8RjhX
MrrZ+LT+pCtPJ15Uxo1Q7mlZbBy5JPqv6zg2Rzn9m7MJSXyBHJSxykA+VjcjgiG4
/84m35pvfyOa+Pubb6sE1HLvB1nHLNQPugs8su/K2rDGLcBBfM1xIRuOB72BKE/H
Do8ghJ81uQwusm4iexTW0LhP0uyAD2hCgJj80llGwZV+ODYi5ptELXN/BUzjyOwj
EApuEKZKtA3m9Kyg8Np2hSvm17eBK4ty2J3LahIuqxErP0i8Q8vvxt2h8DPRXGIQ
gKKIzx/gOFI6PRpVEmGnnHG+H4EsvarbyF3LLvgYP4HG96iTv61DEA71mZ4q6JLk
/Y90xLxICUb6E3/UdoOSx54IKIrqderHIvbSswDNyVjp+Mo5jOia+GWO37Lcj1oA
bH/yM6FS/ZBaXjxqMrXmWe87+TLm9qRrVMlVG4WOtZgG6L+oIrVy6/Zkk/p2LC8u
wRyPiv1dLT5LEpS1WxZUhdcvwp0HG6ucc/IGZ6uWg3H3vnI5ZN+hrfNC4ZGRO/9o
wcSo61dLkrhbqS+dIGyMCHBDeqMdtfPdi3bbLcbJJLGHCxnvrMxTymDU+MM6P7oE
DbpPQqVQ/b2LD1jlpknimCLbLg818DQyixD8XxyP85ZW9hpxewjyjB/IerDo2zX5
cq7R1d/LCDiTN0V6o+fK4HxlQmsTxzfN5KbIx1UHRpl5GCJdwxAhT65DxLsFtsBh
tbJNFiecwroZXEemBYYTcfW/ZBQMLxiTFP81YA49NflH0s9CARUGHcKHaQ4n+e7i
bXiqPT9d5Q9lEVhFnQ3/vlUo6/LJjU3FvK/UeGMaB3+2filgYZG72SFS6SfYnord
QbgCJvomrIfU+YSUd3d8vt5+9nJ8H1YsvfA+fLkTGO6Fj4w+fkp13dVePb6qVVd8
d4jLfKzIalV/DDX384r2IeAlDYmb2OAyJjddFZiKaOxlFKjLnBWkex4vVQxxE9ry
ayP6bRJDJcZH4VOvEmhmhdGw3kZUONneSgOIFj5HLEamV52V+i22tv6RLG8YZGSr
WPq0niJch7T17LCIxqwpDk3PCi1X2N5L4XU89bxvw//yqFp1uOhKGgrzf/tU6576
hE4pwshVK85fT+gDQr+WeowpbzyhF/fqxynZYYEx3R10k8HaPLiEQRH1vkOnBeTF
Btv1Iqttkjw8LdPnzdWPpjeFwgtCEYL5FOZfHgFk84F2j4d3Chtw4rOINXATfVoE
vzYp5ZeJX7e+UYKy0oYSbqUwmqF6HBictgm04qbrcuG/cXQX5BZxIA1Q9EKHuma7
nrGsfMu66vA1cOcF1A61VrLk/QKk3mQjTzx+AsFXGhik9Ae4rxkBWa/S52m3daKj
Xs9BwGFp6xSn94/ohyja7Sg5dVf2F5qfBM0Q1zVIMjKShRlLLMJxAbtK4cyScg9/
t8Qv9olEA34gQgCCaIgkkt1mOmEsJ8cPboPMkurmR5R1VQ9a5MppDuDgGt548JF4
q9JHwAMHdL1K9qoAqPRVvNywJ8e9ZDZwCn+gDckgSpY2ex7jqI5xO5GHwbIbKYHV
ieD/OnjXAtkLrhGw2Y68OYFyRp73lhC3au1ZwBTY8DGXkPgKxYflpwHYNuZgdX11
psrCnAC1sJpTWzUBwDJGs71qlWdxjm6EnVaANPQzMGboM5gt5qhyPvX2LoWFpe7B
cl688MQYm3qvbO61Yv8h5B9fTKTRUbS3+lNz4qLhx+RD++BEW+EW8iNa4YTHzF/x
uvL75XiVNYJzhZo/EZU+D3+PGnwI8vj/H2YYrCsdLOr+7rP2Kop92ToUvPYBHPlw
BNbELxgZHl+zFwLO2qo3UHIuyK3i5WyZYLfUJH96/Jeyfzvt0wRrLvYcJ4xJsWyP
YXBW/bMBTTtEG1UFgr34tXwCevgTDb3XykR0FsRkbJUaUm6gCaRz9Czkd1dXN+Zl
qf6BT4lDSjnbKFmet+vG33nDr5w7/O6oOvy2u/QVqoeRaQ+/rjTSljweCdvPByv7
VelPwAnU7LWRsZjRMifXjABN6Co7Dj1JtMAt9kytL6M6qRPtAIibYKJO4H88lLWI
cFxTsG58mTtThlqbEwH1GLHjUqHtU5RwITIkVSw0JzOTWgSSZQU8BI7jkrKq1C1V
vp0FTmcJUyaZhS5gM8c1WXZIaTVKa711kYB62MQeY5SDhDSTcuLfS5SYePu2ctwp
E2DNWRh0Wwr9GnmAxM8tHDAKRoPYYG6UT8hY5lJV8httZvEU8IQVQjHNMs5JsxrO
f8NLGtNZnowB4FiiltnRq80eopjjBVhlt9XQ+0xP7n+cZmmWnB91cD40NYG4Uumw
DLPy6bhA9aSx1EoJYY6g2nbIpXfMElxif72kItfVORCt7OQrwUN/SU90+pEFCIIR
KXBHJwsPEawaF0QGsCf+GEY4n0ZtJJLSSQtJ1N8Btqem/2j2+v+6jEnjYesQDGIO
MwOOh5YOiy4GLchGc/lhzBcszcfuJU9ilVkTvcQhvEYeqRgOCn1P6VvOspV0w/od
EXm7RjoHgeRN8odEL5PLanD1JM/DENy6sV4h+4cpu04fztwh5izwL3GoN53aFGX5
ssSV/01pl1jEpX4610zKT5+Mbb2jmtklYZlbCrS0pDoKJoY95rt0sA8AtpWOcGi3
SK/QUISo8Ntm66tqD2+EFOuIi3mSfjO/vdMp02aIypuYCA7Xbr5FnvaJt0X0WTQt
HTT1wl78/DKFNtCNybS518Y4a3Y07xzJRqENp4mRahbtNIPZIvQTad8Ps/jIk/NZ
1LWdZVEBGQfoyw5I7hv9yM9oqWFin3kRhcqE3hsI2D5OKkEf+tvQnzF+AGuvrA/c
fuw7glGjboCo7/EmV0HMXFP/a4fE6HJyc12uuhxGvzBaLy4cPgQI1soa2WT6wbO4
N45ZstyPTlIUJW+3164RojiZLhO/n43CcMMIdLboAL6Z1xC7J482ydRp3LGWbxzo
y6D4KMuY4o8U27Z0Ff93VdCxUvabNqefzYDQ8rKeo49N0oarByhoxx5gHDUVifUW
7MUBQq6lGuJBLqiaLYtrRUeOxmx2j0J5OMqeQAX7F5NmoSgx4On1ywzEIVSmwVEC
FSLVqSqIUJBaVieVLSB6fZU5LRYm1e0DtIqyS570YcVPB1p+ULSX71X4/dEspPO2
SCFRzkEqRPKll3FixXnnj6XQjHZw1H+BooMsdFWq9GeToi8vSjkQUbYp2LT2LTm6
L3gpSJq3617IUci875idwrEgzno6Jlpqrld0X70KJrNNBF4lUWVn6cekUi35LTaN
tL0E7lEJdtej3qS9VXI7vvWc9Z1J5K455rBmqxpae1C+lDwJueBE9Zjp13A6UH5d
7y5NvHyuKiD85YEqg0q3cIfQ9fOvT0F6XH/j/W6riiXpHjCtZSD6nToHo4v7/eyx
wt4KUXKUN5MrTtLvAEVB/MYlTC8l5suHsKeb7y2d88er/69EjRNcS12Wt6fofU9X
2ZfetUyW2N9HrwCSFaoUDJnUf2/p5mwPkGzAvcnw/qxmEHC/pubwvrHO4P6ugSnt
jJLninTZImWAtpfg7NxHwdJ7gmY4YCTixRCgpZjXz143M0eaIAiX40sdb6nqcmB8
HWlbkGIrDP0aXaZzrpd10fzu5HBiB1A8g+QdIFCJUR28MKajodbCycBB6MNkoohj
lVuPp0x3G2aZzwYABOg4T1qoGYuaLRlxi/M4aeoyz2pVE7QakQSlGFhSGB4+ia/t
RAYY4D3tzPBm4JGaJrFsN3GmhbKjeFjYlxXN7CQP4i5fsgeWh5SFLTAqSXDLIZi4
TBy0AfqqelqQL5/W1dDiG9dAV8vKYDkDL8ZutHPWIbpl7qy6nsfgVVD7jJ51zG7i
Ha6CLG1vDCcwrEY0gM/vHG6Yc9Tnz5/3m8bYWFqk3D+xtf7Z7VFLUWnkut6SZ53T
rnBavLGtpTXYvVEko1Kcdq+M32zhSDAOjrXEOAmVwByuJzmcmmRs27dmY2RGReip
/pkjZG9HFJQUok+Jw8yHkuEA7gERvvO/+2XAIYoo3auSnUHz9WyLG8/PBoQwq23H
GCoSXWtnwRsd8swlxFdNfoLejz4z1hJfJAi4rjSeyl8NqBWxlWAYOy8G0BVp6FQA
azNdTxKmzyWxM0TL3q4s0hj9hskMeeDeHS6n/CgBcrTD9/71DQ2uBv7h8REAZlpJ
+MbPkUAw5kMWoMLJUWhIBEMGfmqd36YIa9kFdTJlb44h1aDjeLUDxltrGMgEtvF0
WLf1w5NVuowsaSx2lXDdNiEYseqAVvxVeLmcws1hsvd+w7JJfBTlV9i91/LzqbnZ
D/gt2P9zk9/iRc9sJsphqaWMO0gJ6f2am4zhDKXH5IOCF2DlZmb3TcYr/ClHf5lW
yirwSqg8v/9QjrytX2Gh2M9+da0SuWfOrYpUGO7Rn7qRRLxkD0kSfcZZJpjzeGSz
UDaAGKsKdRBbsXuiGZ6tWcd8bqxtYyKjew9pxVIiZpOehxoXdsJqiNDpW4ZImO0T
g26hz85Y8LsreKXz6GUYnBz2CWeLorlWvjfL4q5jPQs9ui8GSMUVsKCrOdpqa/be
lBff0ZSl783ISVyyN1CdjPUcNDFA1n9lVZ4iWIS5gK8cw6NENOv00Qo+8zeH656Z
E4EXVl1knG07vlPGwU1471wh4jY5Ed48Fvjcasu8988iuqHabepwM7sApF3ouyfR
ikf6onFubeZk6X2F/5daV1g6Ccw+C6OzCA39YTNKfAb9FjVypQFWWKcS3rOIB175
VtXaB0+X6KQgIM3UUn/0qMThq/5X+CuF8/ydgTdSQ+/bUH6n37St5K+eckNX2VbA
BRFZ2rpuCdzG0EsQS4+sDweUs5jtqp4NrZctQeDGEez53ocfm6P2MMbMLnaH9KtE
bSfUxkqRe51AyPS8a1UqkY9J1r0wgBogmkxE/fdQejK83bb5RXKvGYtZloJHtSEf
l7m8iAAYd/ZyuP5bn/2bUuivmw7jU+abWYjSc+fSrm4PM886fh8v5c59ckv5SKE1
84CRVQlkWL7MU096A4hgP1v9bQZRyuJOGzMvi0pQVj6w/Tpt8A9TKyji9TdVUQvc
IM28r4jEQFR+x22/JTywHXiQiRGGB0SMgIyv5CjHo60a/K+v5ZddqlpPA3Ox59+R
8tpEatffaAUg4NCAaNCMgRUG6RfngDYrB9XuA7ZdbrYWFI8RrTZxDPaeGEooMvZC
/MschAtRZdG/hkGzAP5u0uWsJg6eTQMetgLiTMfOJXkH/CKcH7/mlqCvg0Fu0rU+
dr36d+VEh3oDStWKnC2ecHzFISjAaMwuzVVL3FZocaJ++mU2a7Ns2H+pZBdm00s9
COkKvnbJidiJmrKQ4u8Y4B4yI+GIy+etfV43Tjz38Vxs3RDQVXW98SXERTVnbWfZ
qxi3VWNiNXLoBY1Aq70Ms6RT8S3aDgHa7nMXCYeYWpATL2ov//0Isa776dl9Vuvt
VbbwVvzoi9NY6UuyqnCbDcrlC5oh+rxOLzT7dbk/myN9TMuvwfENCINkYEZJVgVp
5Ef7ibtpJg+pNCSwi+8FFpMP2BqBjI4R7+O9sfR7Ik3PspW5Hxilrd9LCelbJMJz
Xyl8QgBrWSWXVgb8UptOkLVj3TnJ1ERYDllogiodeVqPp407cJONDBc8zAp3HZK9
enNOZ6rA4IVY7pU6l4RoLE3xp2CWWx3lBAdT0J5OUjqhD9tY4fjMKV1OQxoj74/J
1ZOve4Ar3UQqoCOTa5Uh9Kp6jm1IELbS/H/sGySgRYiiKl0Rqg9lDNgVYyf4uV67
xgW9DgXDycmtc7IpDgvuMkqAQuSo/tAJTX10DuMYl0H1hdC/uXdS7FYQSOTXXVXf
x4fToXqthIxbwNLovDPolHa9lN4P1uHIo49p2VlU5z9X+LdH0s2prqA/n0Jwp28f
53x/1DhlH9MhpNQxR0i8+2Vdm0XHbdc0RoON8PvHN1tHXjxHkrG0WNcCTmazdY1p
K2lFq5Ef4ZrwQcWml4MFavIOHxgFlUFksARPUJ11F3fqSSs0OLEoYPyNmSWsN16x
doWh85fNUfEeAr6j8fNBZ4iU8CxiCI4pjfP4m5Id7n33uGH2rSS1q9eQujXIwFXm
w8Jxk1DCBlLNsxu2kTPRQYbvpJBytDwnOIBOjxRdZHEDpZYPiIAfh5n6e8/KMf5/
dfRRBdYP5MA49N9/Yrkv7+QyUXQYe1QaZ3Lkqax6cjRmqMi4SOJ0EFa7SsMQ/duJ
QVRyVRkc7SOeO8pLa/VOejeFhvtG0y6wGJY9D0j2J3vGUw3gLcu+t+OozKD2gw0G
qBg8BaTP42Rs4gWuJI8PnwQBNk7mwLEXmwYo23XcQj9IkJ7MxdVWtM3jHJdGiAy1
lCuXB2Aiy9ceoAPLwhWOlJvax5DmCv5Fapj8L7+vlMiJ0urtiCLUzadSN/vPSll+
aIG9xZSSNasYwLLc7RTx4bPqVkROoj3RAvsNUxHMYtLS8VcuNiCEZC+lzqvv0P4s
yOdVSktpD1lJaOJ411WEL8MbFPg0znuFDJqfrM9wxT0rzwYc1GC18Uk/kHMeN1CF
7SFOeLCDYUns0OEX8SsRbtu4jZB4wOFXWuc90Soj+azD5X9X+4aQwSe8H8REtXtp
RM7HfJToOuyWq5x5qZVolxcnUaajGajtp9hXPZprh2aYpu+LwNADmEW5IJAuXmSM
djxCDA6tI6jC9Py3JwNAShGs0UhRAIHDITuo4aEf9BlCqpF+c+BP5aYOG1ZH2XW4
oZvnqLCNTw/BGqUubWCUZQf4rWxijsN6GLcZWf0KwINQeWcKK3JoyhO2vA5sUt9e
+0zmU+mQunK7sXVuS5gc282h2GHvtCdz6QVTJRQOUBvhjKV9BFecDCUEDtzeC0Ao
TnUfwHOXv/PP34gIXP6Ic1x0hJ/BExPWnSiOAkU5a3Dcjaqzy6TXCMvkuo/09dO5
e7iQPuThWOgYD51ihPp4c6wULpcxhPDK+eKZywkrxRv2uJF8ZDcNXusaLZE6MZYh
RDGp+jzQ1goIKOj6OpOyJ/vTTAyZZgv5T46eV92Dxvrpy7CkEbUvEDqL/7kQww85
Nr624c7d844CbvBCSaEIh10WsCV1f1DRGtlPqPXf6jer/fhhhCbQLw//R3GEJYh0
Lf8iwzO3dGAY0zgfUC8Slq8pTonU4cSAqYQEFmNvKwU0DuIHDgH+SILzH174LjIw
ScoBbYd4Evpz3VphBrkMB77LzofSYc3Lk/KVL2vXcizrf8j72M+rdEqSFxoXpWpi
K0u4xE4CgrqiGQ9R7fNtxgG1704vmATpn/n9Snv3O9R+2hvXPhIK/iv40nyDX4XR
UK1xNRFqyGJkrFrh8DRaPd3jHzaglZf+wt7nV/r7dAiF+O/vCPBE23/Ir4q9/jPk
HRtCyteG5apRnL+Dd6X2OS8PTs+4GaoTaSmjYAaL4PVXrSRDhzbrW00mFYBye0J8
sowh9AnGvjYc6rjNLZTZ/RdVbLxX/xNbOjCskQ9pSfhFMkvBqG5KeVVkDaAR/HOz
7IJVxdpbdbq6QidAOfdx+qxr70IsZaAYj/7oSYgJlFVFk00Bc4P0D5nr2ee25Fsx
AaUBkhZB8xVX9mA5w2iKIomIYBGh7aVPXJZ//u3lZyGalmjSSpv83y6sK6eDWoE8
o0ldnoGTB0oK9+V4n64GNWYc34dldj9/o6lrZe4ciaNXApcoeTf5azeW1ejU423V
62DMZZ22ax19FxUv2M2UM/FqnjZ9N8rk2OQy6DNmuNXlTxr/WkW7PgFiZcFF9XIQ
FTquVtrGSZ132aQyd3PMfb6xqfKI2RzU/nKD8j1TzBJyAuF+H36FI5PqZi7Pl9O7
XkhA8ACJeYrMF85jC21/W/a+uJcpTpltfpLdGD6pzeYWQ2KTRT7cyZRDUeK7TRsb
iOuym6MbAHqUJnsmla2Ot4KeOIBFko+9rkk2P6UrvNBYSNI1kKMLNpP8Hi/uVm6P
F3OwOlMWtnybNXUBN19AsXOkYRQ43sJBVyqgQNq1meEPCtzyKlIm3LRzAYPhrddc
RvUfmrPRSznyWqwmtE89A1G7HZTqVC27C9zBeTObhuPT8tfFNvWdgprjd/JlpE17
pGluPVCh2GAIQU8GpaX7UWQFUYS9R3UcRie7L9nksQjNpYji7VbkLxhm1gg4yieA
cttR/daXlhPA1KFO+bAuKsRkamg4GXDMKiDMCM7epwuAcF67n5JRuU9l0SfFleja
5CxPYI78km8UuPMN+YGzOipyvI6TDfWLDJzG3ubQ4ZrSftRbPMdNB0yx9+zJhp7T
w64d5n8r2Oe9HJRdTLM1O2oBxWMaSFZNKO8WsL8s1XganQzPxa/PtuUZ1pKuGRrf
HstnhzsBd4B0nFdC0hd9gp9XR8avQq9Eku+K0UxmRMJad3d7ZaPTyuTFwQP7qLsP
+wL9VbXaQDz/U7oS6EorcOLxCFSRR8hvJv2it42xfY3Pyls/zGUc+UaQ3G9cJfVe
XbraJ9UhRfHrElAfiZVSedD3fbmbhSJH7k6jtM8LRAem6CaadIPJPoTkzl6+WwcU
kYx2YOCEC+2v4gEf7wCZhV5QCGnb5thZprO3fFij2/azM3aAa7zW7FPqQ69bmL5c
TazSyanyH142XH8NGrGe7YEwtjFATBezs3hKwUZC90h4h20MiwvoORedF427tzYT
kwDbb5O2KtePGOOpniEGeWFQ+ufXlNf1mQ5l3FpdG5/g2aCCLiy9QmjrJO93hRhT
vUEJwQQoSuRKDrcsSJDdmycBQ7b621KyHz5dF2mMZAsR0pUGtE5mKXsidMIkvwIQ
OuQxUoDbsFWabGSflZPRsS9KUQM0Bf5DdmvzH6xieVwIoz7cTuhlyAlPZa5Twcmj
vqK9geFwOinHG4Yu0Km4qXS7UekOSMhBYCMQCsXcilgWaRRZCDXSmfWTYlR6rxQ/
JoqmUSBooPOsFL+gTeQiT9aLvepiixc8K05EZAmCRBLkAHKGehcZ5RBGuIn/IPZF
kGrYaN/tvPIbF3Xi0kETymEAF896pH4MFxqsSi7/Kx7njRmHFPUShRztNKGTw4qx
8/gDaaItHoybnCssZlW5BOsfq/FKpuyPPT4Xa17uKyO7QufrMasYuds28jCOOs//
douC7t4GhRU+u1mjgVudGpjM1+TKOvr3YQIlNjyOh+72dB0S3SWYFSPzM8Fsz2KA
/O2vE2Cme8ftnnafy3vGKJKly4b0mMGenU550O9oWB4QwLAq450L/eOr5BjFxNLv
EXhyE8EQVGb5YRhw1URj/GVIQxun6ypEW0btDhQEuGYuM5ZgMJxOUmxwXqvoZi5+
MnHBxdVT246PPYxnreWb6aWRuaUx9BxDcddFx832cPyUDnEEm054ounriw6HPgBL
n8W7fsE5QbVTNzsVPq20VPKDs6+lxZGIVu/P+nW7du+gGG5iMx5dvMNXl3wb66TZ
keZ2ecVkfrxURtoqiqpWNUMqSwTw6UiK4hppekGrdcMk7Cc4FlWeMTUnQKgNav5B
8oZSGAyrYHmuggQwHKU4vUwUybl6/T/vRdHnDooRmi15q5Bae9Hqo27zqbA6n4IH
NfwhLTUHj84NwEVCpuIIHwCwJrUd/hgBMS23krSE2/3jrUKy8pOjIf/QX1qwZpqg
zrhUFSrJ5hKEowd9zcW60ckTHagSlgxFId2prUHrQBFOtb7WzAKlOhxasdClkFA0
hLhq899cd45sqbcZYCSu+GK2yuVH6CxI8u2xkKjDljBPS4Zi0c9CLFTivJox2x3A
p7f579zY60cyT5Z0rB8Bg6CA95xS3vWm877nfD6LaRoPDXsrCACL/WfK289Yg5Gg
h7A3EhqpotKMCVMOMjHPqu2YFIvS9J51qtENTUh5uPV0jxp9Hy3cfbX4FN6FYwwj
E1to6bDIqTX22dryIpslyFUF5I7rYx/4m8ytmZBgxHv24fMvGFvMXztgj3CnTOB6
cShYpoAnln/WU03nFAW3tk0dQ9seTJ8TZ2IqJ0b9FTv8NljaHWn1dWKaiUmXfMck
FhoTi+RGtQq5rOdu2s8iFPSG53LkO1y1LqQFJQw6dMnIUp7D6LfNmFDRwEdt+xX4
f/1jvYFTOTQo1/cSVbH0GIhqkrtvE32IgG1pwSUDPrp+0VuFwyfHwIqQVu9O+CfP
2taTdLEDiMcl4Ss3mUVL4uiA4pr6GKIrLsbEsl7+JAamXbYFPU8YOXPid9AEDHnG
U3u9Rlsgb2PhOpB8vzsb0op5r6m+HLIoMizeYdsOdxVB5okWPMyCfGow0BQ9NBP/
YNsOvO4boEvVScS2w9BQmdQ4v8loz/fs7+jt8TrvlhHSQbYIsqlsIVwSpz+nA9TJ
4s/75HbkQk0Pk0y1SaX9MZhCgekYbvI6nyIH2dMOw8kHtBrB9kzkLsLvaBm/gvdB
0NRH6Kso1p2eLGXbN2/VN1/j9GXaPy8U4GiD7m3cgB873QuU/kps0mHIQKdlUSpm
P8vkLjXT4f99d7o9nW9PpeQVmmMPIRT2xqLv1SPwE6yrPq08xoMsvYnXcQ7LQMoB
43s7qAe+8y4YnoMp5zDX4mJS05ZYD7D5klJ7RZybsrBDYnIJaAzZGMlsGDWQU+Ud
fvY4g98LaiP7J/vBHUqBzm7Qs7/Cy+YJMI5DWGnwA+cHOoOb1G5/7wwAvxLaLZs9
PC8Hr9gtVRhItencC3P0RlVD2ZzHlCvUL9bDecz3IfADAa7Cq+FrO71AfuBw8Zdm
cne4WeQj6/VDasivwRgKvOzdH8XljeNZbZv24SJP4qJympc73+bqvhlKbwvqwNss
mbVHl/vjsBeVN49z8IvpXJcqSyANDz3tfdpiXeILnhN/TrWqU5Gr7D2WzuOTR3GA
QgK5T45A37BX+ZksBMrxZ+68CTtNPoJ4Uh/Pr+Vpia2LqA/MtzJOQ+BlWZiGgiZs
CG5sp3ZRztst+OULoPRrVhI0APeTus0BxYq7L8pirF/2s+Mz7EI5hOk77JKIi1fF
GG+KBuo4rJM2Er4A3AEdSjuSz6qU7eZGolB345qDN9aw/akjIyu+I/DeUNMFAsIL
qKYtR+1NPtuRL1BVfbAz1KDJ3u8+0TxLFSWxK5vBXKX/piQXXgfd+T/m5fihLhqV
Kso1rJMo1X7jj60RGpwkbWQtN0pbpCC7A81PjbVCLWTpui4lzI7dmxcbMWJT6RFY
n0rnOfv5y38dLU9dd9tzmOFo9SKv20Q+dnS2w2jCEJrjUL/UkEn5zqLDs2EVbZ2z
cLmqUqSujJwaOW2lC1p1JPf/8T6GJc9PIwRB27F0yfNMfFmDzRP9LjjjProQS91N
JgQ+i5O7ryYPvEQ+L+RjoKh6P9alg6lmNPcx85sCfGXlz4poLFYrH37syChqKlH+
XJSfVCgFQEjerqje0zvn3k5Je7hPnxlM+uNMpBhdu/00uWAkhopNOAU7e9Ze7cqa
0vwQVxbvE/37OeNmCQM9LIscOjBJvkHkOgnMS4kCAoXLBRMOQdZgEof7WG/duS6z
FJrOsYRQ4mgzbjMbnFzl/gS51MNIuq+skkEkW3XrfyHBIHGgmNzVefMWfYZjBfMB
Cct+eXqBQNN/bPnxX6zRd+qrwMqTmeOWBO+2GtfyNjJpEm1z2xuPRuVl+hikUCMw
SRLg74DI+aEP1+44m/vFjiSizIzvYlMn7VOcO+NdjiwxarfZpc4Xz4KqRjcuJ0dZ
HJ+ijlNoxVfP8miNk+4ic6uUt9CYnVmtw9mUczu2qSSpXYeEvBk56AVaSsFKTwV3
tp3IBiHk+C1k20MDV9QCYi9TUykBRZ4iPkFYJzzzQEt69chgZNNAckiavdlrt7UO
pLOsNtXmu28uLEilyiS/57b8EYt1Ko5gNj86tyLA3ki9jzVi4HLiPUyQ01/erlfo
zyG+3/LjeOLs/gESEaYL1AxOxfOB5onmXGacGtmPqhyzhm3F5hPl6/s3vzkRWGxD
I14O3vev1tHPUjD1sCCPmiRj7T5P9PCtBX+avkIOrWTRbRf9Gs3Du327QENIuRdR
yrqDgk915ZSCYYkQmusMm41TtufnOEzv6ic9kmSGXiMZ/zi/EkzoVcoWhXY/uONL
utdk+vmUJDgHt+S+uXqzaz9JF1XuE5W2FspZhJU9dKBjMq6yH8p8BXhVQKAXOfoW
U8j5sS9ltCDGdr7jMLOM94iZwS6qSF8HVzLZODwAUQXfhvNs24S359w+mjrDYh7K
BHPCPDUQTp3Oic81A5kMUkcS7ftu3NcXeh9u0Pr8pAdQuKgoptx9DGWK3GTB73jj
9vv6IijxYi8Ax+J+UfapqimfzvC7g98/JMJsNuBtu4jL6oz0BnXvQFYJwEjHW13U
rwc+6ET/Du/c1yyHLjq0vXQZdE87DCBddjHTZwX86ZpzWWJUt8gip+HyAbSPbnP5
oxJ/zYTgVbXyp4izehwv1i3HaLu4+Sel2qUKOxCVhjOhJrkvmPGKHmQqYNNgX1GR
go64W8zc7WH7Ue4vJmUGB406e1JsHFlYXRVnxKZtFglyxRrvnGq9fxkpYixJq3EV
uEncvNY19LajgMBrUIgFg5/iQdQN+3GMwLeXCZUqsDwn9Ui9VqEYn4+DP3aVMUd6
CajzcCyKu8yZpr/+W2AJu0prgaw3FApa3acVeFuyU2EMGPOdZ1Q+G5dCrqZ4TZno
4UzebvZdmesQE3Ejt6etq3GXtX2+zHyNFpTXuBfYuoPAKa+t09g+StTQ3QBELene
CpApj7OsI09WAMjSTJ+qqj1VtGSnFkLqPSsN9M0N+vrLvuRb1VTWXp7uAQmyKVP+
d01ZoOuX+YJwps9fEyCxG+QYlWqwdQCOwty5Jr6BQtUc2ai3vFMUJkZjNPMI7Go1
EcO8ars1kE6t5q0av62CXsKnagFgkNjY+IprQ+ulrUUSniV2KGNB9q70oBaQQdkE
qTNbNk+LG7+tR8gb1P/janRmnNjW8NjPHLfepGekHEe6oUPCt5JYcCWwuoLQl4n2
F/VYuO/jEwoOKP3T382csriLbrxI0vgoaVTWG1yXX4/R2L5TOMuEDRnJEU71IHJ8
WQPm5zkMzN7MHAoPJ2IbU7FvaDDB92S1KK3+HAUpdfzriTP8AsCSc4d6WelTpYI4
jT8akHy/vWtWvbZvW7zaTSchjqwPOEmu1HPw/lXXRdCvZFTUUATyW7CbEh7ZAkUY
mPCYgQnrMplTj0yf7eT7eFMuLxx0Wveop3+1/NDBsWXoS/ppKX//BjI3yapTiK+m
AJwlXTV418Acxev1WWw86vRaSJCvkecQu4cMOX65ZrcrDKH5ofk/hmOhdLfRSJ+J
UrJHxvagwwoL1CRGPn7bb1LaXL26Fau0f5H6T9c0T5D02YPaJeFfKGW9669udiER
nXhyuBpi53Qhmlo2Rb58wUOAEKoNC6s+2EPzKnaQxLrlRVmolyhNnNGf19XFR1Xs
bjVHGZCPy2vWEdJFFx8xZAYQEZ7Hfc2qbboe1bJ2XRhC1DtvId3rhp9aBeMzIu1L
+E8XlxptxH8/kuwT6jY54NbFb+gWaA1vXts0Q53yzc5mF2Dqgfeow0gJVMuFGiYv
Hqi/8XRa3ct73K90rd59jHR/892ULwasSFa2ZDFbdrXCckNXuJXau79dCrIKPgD4
lqm8KrfTJTcRE/Lb+lYV0fWhUXFdK+ksT4ywMborXTWqUkEhl0CDlavgp6IrOgXP
9H/O+7wqWmlABBjxO2hZTb/GqqUZWnKp+pum7XdhiS1NCRqB3sFppE8VwqvZNGfm
J0Ie6y7I86k71JInPkC8sU62fkDMDYRr9zJp/Ttf5hF5L4xnY3etpe6Y6u1fsh8U
zKX2cSlsB/OBKxM6ILu9NkyWMvdF5Xfztg06H0KucJ+6Dj7Rm6R/8qw1KzHBVJ9m
CmzGNHMdhFvUJXBdb/maQL6q7BrUqKcx1eNBy4c4OScrRdW8JjNQSVp1fF0/89YL
BWVKU1NBGGmB7HzWK7Mfnzb4cfs38ZkZgDx6f7AwKRGCmnePtv3kGwP+zoaWlxLM
oAwyHw1eEy31jGnrvUqWWXj+06G4f9t534ussD5G318nfSMnAUy7+c60qXArPLNa
KHwc+QPhNLZ/sXo1vFvsegSK69KzRJxEi9AtRpiRHqEhQUU9V03i5FjATLRJj1F/
l8s11npk8toxAgsXTn8Q+o9O4CyQ945S7Oio5JXpoE7ZkmhnTfmwTLTauStuboxF
eD7G/CzbRq5aB4vbR/cEOzwVMZSHYR5v+uAclhvHty1JbfQViMWKUOhEhYdeYa12
HkIP0eie5tSF6I9haWSBbm0yaAefQkrBBUvcgUZvBjY5fnmH0p8Vki5K/qi941Te
0Ek1FnkMA7AllffLAjKUVkhypAbhZdBza8Wd3azXuvUUVYOnH/x5iDGzIi7S0RGs
4oCfMoal63fVHl6ig76wlnXwJ02JjnRXMHLbRwkVWUCTJfbCDU6ixm7WzaeSTziy
t0FlXdUhLbFVQ+A+BzWxw9wXDtOab3Jg0QGc78XMhgTvYlaQF3/QSTQpnblSXceq
xo75Fzp0+6zIB9BXAUUTI9Me/EctoaVjYDUJT87NG3cgSomwqavbCxb6m5UoPyiE
bBdG+qMh42BvZuE2HeN5y+eoNy3xJIFJ6pS1VZaen9bj0w1zExCK4kVqsQQZT0dC
mxcsum5bn06xN5hIfdjZrCaczpzLqbehqVrpirNQUa02piqy/a6jhGx6hF/IdZhm
QSED4l0wVHRh48fmSEf0acsxO7JdeJQvFegof4vunQuRYko8/7Ef1AyTvcaa1PUV
nImeGGO6WFQyQvAyMQ8P1cmmx1vJchdZZsGFxr3/vDL5qTKw3Ih79Z4rzWGvYagk
uD2FNMmUrjCJUBuQFUZmj4yGdwZ8GUZPzlnJDMaDKEovy+ghmI3Rjg95gB0XSYI9
qM5PdNlHULvdgLXZm0tZxrtj8Hw+hypxNoh9K8s7hn5BkdSkQemFH7em4WS6/0Gm
odiRZ4ZCWdDq+5qok0GMDnCLQY4EV4W1uHLVZ4N7Cqea1B6he4EXhytTXPdf+b6b
RVxWt0XmyLtW4UV0vz28TU4ULSKgCOIgvC+sx8ilCPzdtvc4vvoEQ9NSbiM1/+8A
pr/N/Lxe7iVhZu5iARZ0W7ZfGLOzHsB1ExKmjL4+SpXSXQWFjUvVhv09TigDaRQr
gwVPu+iRkstvK9ipykN6g5r9ZLhMLwkWPEJaILYNEeek0/bBoFAg4T7Wj+7YYHYO
OyzcvSMiEiQO3Xh/qd5Bo2kpFHjlNQ5O9VkmqP35IXgKZFwLyupuAtOvxNcswom7
gLxS1OkaFSFEQWNmXlaOKZ3VmxiXVWsG81IxgN9Axz2xQFilEx18NgEpLjc5/MPU
ohlp2ddV376deGdn/hvmXYFfzS2ZU3gIzl4Bgc8luC6uKaLN0T0Eo3j2X0yA8VVP
iWkzifJXSiP9JbDLwMdRg8eF66sp8DIavqhmGtIE4ZpoonqKI+72kP0buTiNdwPg
8KkcK1SCBPacinl1XKduXy3VWB2wjPcEhsw5rbc+ILa3waJRSX4dQoKMO748IbIV
dIzLVEFEZ3NCD+o5ugCWGhyfquWPJsVVsFkQDe2HYMysFCaxkDQ8VBBLN0FdFQ85
rcl3GLTOxJG61puh6DOl53JlKGgdY6NqAtOHbnSToEigsTz0f94eQzXRn3DVBiEx
BgKorFeb2tFO2s9BDVGCBzyOvvOZvVRfy+AzPwGnR+FcTP4bee4WgSZpm9u62RuK
hHmj+wA7/sqejxCdYcOtCCEuyCitsP22FVZHakCFRPKnqZw9ooNMMnnIEO4w8aG6
5UVlwt4wJGcguNLIB/cAjcB5lmpCk0T9YBqnYV/w1751i6g4864w3tta8R8p3oB9
RZqhAmupFgwAenMJ5bbt/sr0XlQ6XkSU5LOUamP/TJiUIvFMm0js7oDb2VcbS88k
ZpiYxjmE1MeSEqg2CN985Y8c2PGxB6Lg2rENHeJ19pRGzpzl0llboyQpwcQb4Q6v
CRAayr2wCxmDXZiOraOY6P1wZjGfssQWmV4FlUfbPGZF6l8VfWuATx6qxsBS/29w
ZLDwkcgNA8aGMBSJeNQgBjfu6gsqLKS2lhZE4LFbw7b+5o+CefLRjDIkzqbn91du
WfiJdTnNH+RMwcvTUU2dVHrqW8q5IVub5SH7obhUwLtdHfNCj90X+6lRKts8+q+Z
w2tGUvy1AclyP7YKub6cqHvVqGV11JBW3RIiczTVZazTSeEjjdrrtFxn+VsOWHaR
XPYK8kxB8rwEqZrW+fHEd6yKSu0LZrWHcMr8/xIehCGDzEZaxlIeqepqHi9JfYVc
49mIQwqm+EETvPFresFIH/ZdsLAaOYFshRCdXr96h3kSGTt9vUN//8EZO5QMsH9n
YHwaAIDAj9Q1qlroRUtNdIu5nh5apuoEnhan7nhHfFrKE/3Faznt0WIiYHv87May
4YcphubidKmGO68O8sXLqr3QKQ02OEDUnLmYVX8jZFO+HNZk4n+waxDrbryrwNMg
7Dn1ffN7DblSwNXlJwdGc7la1RPDkuhADYTZrGxIoKthdZzsazLpE0oHyp7R2C4m
2aU3qiva19GEvCMqXFSQ7mUi+WAwoRBcATcnBKtsh68zvj4YJxZOhZVzyAxIC1Vb
Ir7AJrjNrgADY2DL2dXEgkbgRzImdvJQhA0No17OTMsGivHBPYjRWuY7Sv0/q7Jz
v9cgLPRiTwnIRHiL0SfMB0m8M/pQD0407EX4VNYSp5Ea9V6ADBG5XBGfKbQ9vQsa
07B4b2anmaPnuX9q8dyYhcoq0BAn8Zmcs4FbmoNtEZhetKNi4uFeP7/sqKnKgNDc
jtPvXv+6TaeYm4Mxsmkjx82ZJsn8nkJXcRGQ/xUjvsrAp17irxGoS+Yv20z2BshE
J8SXS0u/Kkqc7tzpsf3vpPE9SBp5dbMcoSNf0Xwb+jFoyIb+WqBZlEhgNc6SU6bU
KjbBenqZqCI9tbA2lTFj3NuVUIn8clr9TrId66Md9XAnDNL3OP2xAYU9JYtN9sNz
6IF7eb79stjOifYOWaabqUiDbCf7+cewbdTdyaFc5L8ZE74znDsDSWsZLUgQ+G0W
str8Ud7891W0Ged+6h2b12grG5QyGuVrdymkvbdnkYxK3K8BaOFKVDSau+9JVW6+
MZbSNpUpoMln9HF/ezEAOAa208UMr4kyPZ+uteSooATcmMmF90Rzh55afAk4AoIF
GrEQrCaZId8uY7TfiDTuY3LtTCjRqboS4jADV/x9Wx+kL4ef3dQcLqVPhnBTN8zs
39XjWNiBN31r8OZIau2/13QdzKZEa5C7+uulMNPEe7CaJcGH8jEUOfqpiPZs94HV
+D+cA+oCjefkmEAp4fNqV/kesnl63WrLC7wj/O9XXb7KbDri9CJeUQB36ySw/yzk
YrC7BursawDKELGY9Gfxn5is1v0XsYBBr5I9rV/5G/nuMSnuWoqasSddKtSmBJjg
vftamdejgaYZRJ3+k5S9/8rWHQG9uC5cpvhA+tqnlYjh9WCZG4naOtUQogGGV6NZ
lEt0svlKOkhdI6pSla4buhR9h4nhSkOK1NncpzPcGBZM6lTT60E/XbK0h0zFuAQX
pgwBrfSb1g0SW4E3Q28Qm9maOIRIZ1EPCH9P1dVo8Yx1US6JzeT/Qp5OgYVyKRp2
12wq54RiWJi3wLewiKYUw44XSoumGpphTdM6xiEeCuLfTVj8ntetVmqKdvTNTZzO
mnLDlCWRONIN4+qR+AUkvUcBgTuNpImFoKneIj1VOArKn/WHvx+XODX+OInWE83r
hZSVgTxT4OKOHYHYBmb02R9nzupwvCA6nB2y3EY//PPOJ1jVeikY7pntkfqGglkP
fhUO0r8ty5uEW86loCX/NObz7346PSAii+EhEoLdSJrOnAIyp/9FtqDkXCaKwW65
1TutIYqrJA+CRT/cq5GE8a/UFeoi/LYIPP7sXzAIqNym+cnWkO6m5fMKAH3V1bnh
eY80VkqceOnMG2Hj9RB3eutD+NEy4TeNPVgZX9L7mbQ+TiAiIUk/oXNHA0W6wcjF
uJzh1EsOZkwxBh+d09cw17TR427gqtjOZy4NFg2nl8PXONaY/QDzB4XkII5LMIOV
sOh/qa3TxYTXSygZ4wXTgbU6igdfghwUQUbflAUemoGYQgzxi/JWntgaW1S6m36j
ih+aqd9vWdqTvOg5NT/9/avMbMNm/xi6KTKvUdMd2tPaLLrqZzuZbHFIkYLCEKC6
1iLV7PZ1tC87/E23OYk89PlC0S7WIEObGU6FCYCLC9fSXPuS1giiMOBQ0ZVWqPmS
Yk3t2Al5z7W/0GUCMI6zsG93j8FLP7Rx8u6AWh2WhWY9zBYskXxpvdpWez+NfLB6
+AuagYVKGmQyKBNW2EuqW+P2i+I0deK4rRWOY64+KbvcJRgbBIH2jJ7X7M1oOBqM
ZrkJEdrZTUwTSRBHGCAOw9PdPDsycRXZBdfC5ycCoK1gXme6lsWz3u7xmQ1GxVTA
LTJoHMrMyEDCNgXMGTpZQyWySw9xWFrZgHuPGZxvVKfPk773z5g78CEfQPljSYFe
rjpE8HnQb9xObvaK5djPosaqDboV3JQ/ZsoAWsiKqckzQ3dfdEHtoZIHQkukpiHR
szMHri0ity4sYiiUTduuy0OpNgrCImYGgmKIIiISZNlVTTFn4Iig1DAIx9yWpXn8
MsFlREDYRXtUmvFyh2P/9aZ32O2G6K1IteE+L1LitcasZT1BW/0PgERZ6/W/msek
Wf3oa5+8j36giHimUljHX8QmmxZozFu7jkkd9hRQQVP6K06G9w8I2WW3jfm4AMS7
8QnmthMJv3Fr3ZWep00i0OPOnG0qt0Z92lJxq1HWQRLtTKQmJdAoNlmM0I7XV0hT
eGkUvF0DRqPrJiTDPBUe1FvN9OwR5qJ3gY/1CX4uWMmp3imIVSxgwG9bzzV27mdE
aHQNRUNjZUczPMPNkXeqhETDaUKdyjATPBnYcIciUCFXIofQ5CEOZG4EZGZv0IN6
igzBwyaoY676Scs0uQKJau5yY49Vk/pxm+z3ntAE30BiipePZ5uyeAaP2qBhFn8e
FGHUhb9E/Q67mWiwugqPQvE2NvhjVoMjWxA9yPvv0nKwFDn1b1rDbv+Eax5P9PjN
ntmTQjW/0c7VoRcmqFahVDjL7B31FSy47HTSvau69EPoO1fPO2sgtUMn+J8gSYm9
6M9PBuMDymWiIg+2yEyYbToAkuiBTIzeTSciuSLwX5xeKYnt4KM3Hhwmscq9n1Xd
SSTSlwa8er6fObp67oPdsw00cEOvPBFhDTyuRLBdTvYitjns/vzcGxXuJAxYSZSH
sJZORsutAK9d/5naFrQXGB/Hhj3+6O5LBeHq1UguOPQ67kaJL1ExKDNnkskHtn5U
zp6OA3qPnAi/VJ4JU3sXEIxeDrtGZ4+HXWPjV2ip6FMmHxxdsND08CY4KmXUF5CR
n4a3leEH8HC+MTBe4HeJH8IyFOpMbNttxv3Is0YcR3n52xfFRNghgUXhmmJpc0MR
Jc2E0bXxcPHAt+W4AyCgXN85CcILtzdBsiJq+RFu/Ym34CcFtxSfgWsw1QfiILzz
15nj+irrLo4RXJp/Pt41yGASeTz4e6+jlq60d3fM6vN0Pq4UAm7FfGbjGV1RNngB
9hDeieKVH3uTOkuZzc78XGevvmJMCDWR8F79Wl/r5BVSgMz3aAW48KQQ1nVvWW35
Ow8o5PbBDok3s8uFS0P3C8OGB2yJJbEq+3c0d0ypqJbTu3HCNcet1UxqClpnB62m
zCx/tY17t/qtQT5OvRk4AELDFZfq557sr+PWNzexcOdXich81G4aggS5L4W+UTf1
WjHVBCDljXeRS5186anpYq/SqesCgzbSpQmJu8J4owbKvyH/G8ZSPQpG0H3eYrqN
/OnJkstJhGDXMp+pJVWP9f4mldGbC2JaRYkMU0gasGbc6+DRc9ACx5C1ScTn+FWI
`protect END_PROTECTED
