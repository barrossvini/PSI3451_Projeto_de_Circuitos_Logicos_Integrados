`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9/9OtAnhCQs+pNH77CcH9uTh/6TySyDoD5eIFEJT4RDM2P4qeXYcPRq65DwwA11f
Ypo94kgDJ5XVf5V2/R+K94SSe5GIDFcem6V7Xg1g7fJXPIDvtUPgVZf2dhIifaL9
+hPKXryeKQPlmKYqyODEDbXigAWcFTcMfK+ngxQbgYJyUy/WU9UuiqtGQLv7iVhg
DG0dL/DXK75/IIefVF29KZBxoDbUDav3FK8E9nLsTpcnLnhFRz9wCLcxcQRqc4CM
x0JeyHTkaXyHFU37N97T65OaC819IMeoCfLvOcRz4UMIcQt5agJcpDXtPQB+FNG9
cmSPCJzfZef75u37T+95HkbNvoaFCmlhqHtcSuoMEE5dJyDBeIn0EJOL6ARusm6d
JKCzyugPYHVBI9O9dN0BNhwbpWAzI1qfJgujZjGJOkQ9cmCgGiiv/VoNW9vZjUMe
kbCIsjOqCXZx011t6lGev98tPEWDGdl3eYMlTlmuGNsTiEy2nxzJCSSO4vusUZ/k
KScNXXU5GuU6nHNli4w17FjyVWEqfJ36Opj5PB7yl/g+QxbWJL/CPiwctzPJ2WLx
ZUooVMzHEn4xsAYfs8ZmdJ/+NgKPc4kIDXT/bSAmjQg6V37YxGZFbPer4YR57EMp
UvjFpBw0YfasD5nSMtqiLlp36c2Ciwp7lX4ylFREld5f6BiZ3EWODVyJANXpUGSV
hmIhgXoy6jcKsNefhx2sFyG08qLuZZcZSkQsE6kzzXT4v3odToMe864vBXHQI86m
dSysDixF4tKarV5Ebgxa7FnlbIonjzXe5UgwHV1nGZzoQC3KXOOHi0ulXTF0IByd
41qLdkj+GmuiT8XtD5AF77SP/9c5Flh40/U4OSkirJfxstdlB7qrrfsQP8Fs3Uhn
+2jxPQGfarnBOiKzVPiOvUVpLir1uIACXGkDj2CawKydz1Qe07JiCT9ufBJRPFD3
NVvUp1w1ItCYMXGg4qhO3WZqjHx8WJujzgnDDcjW6gPNOJGbbskDwrJdaQ+Ssygj
GS85QC35+THuBH+6heaCsrvBbu4u8XILs5iNguCJCdfeY6xasSMGJUU+69MNSq2K
D3C3M1kQWqiVJBKmJtc9Tecx4uMkjxbw24nc1qvpsXY6OpLmRhtmWH+JKo3Js1mf
y1grI9fhmD/bIy+B/BXTnVLb0aeTLrCKZNEYC0nKEQPE892wHwK/i3SOVlbX7K4v
BdLAysJF97485QmM2/0ZLoFnSl1Ba3efrntfKfHQkDyDFade5L9/p1QdR/YuwirS
ETzHJXZ6dP7HU+O6uV4X1SQrLgrh9bzCwMiFT0rwy4jpF+4kOjtqaNkOSyczw+W6
i0g7uAIahCliBl3fSo5NjVEyuwnYs6AVDvXG+PG7FGhFDZPlh7H2o/EYr6dOzRfg
dFA59HiwKtyTTZOZcLyJsOkasCW7fEbDpZ+XstjRVnSCS+BLYlFxKDL5wKFgIGK4
Nnsm0aKl13sIPxdlr6PKLq0pV8kUX800d4jA4oeehhiZ5kLS7MUMEzDdb1osxIqm
MdbvUDDx12oip9pIEeTjYC2tluED4XGqLgHsuKFRY/uuIckXFmtsN6Fp/MLFT3ny
v/ymaWP7/5EQwmerA9SjwsnHcS5PFvbNxu9xYUVkTuwkFhkPDw95qt0YSIwnLdpV
yYL+hOt/VyBUTqVvlEQGkeiOEitkUJQ/xAS8p3QzJLxxBdK5bT6SCj5y5qaOkwY9
3pHCSJWpa2PFCg5aeL//0lGmz4fgJnupukgOC/eiMS9NJFAjESUf1fGWDf6Fl53l
Jy0XccLcqTTMQdPdGWh3x7BDG6IzldvmZJWX+/W9r7WXQurPcHolFJOxtgm5j2to
/1mJjWVv1KYzrJ7GnwAzlRkIENB4Yzkq5e8aPf3BcPANIC1YOdzMiqnVmidGXOR9
3AnEg3YX32kTC49HESHdm6r3MUSNOUj5zv+wdINsFGlTVJV8rnlhoGUoSETbv3PP
YR0ohofYWSElP1TK8+ISKrVJQ50ciR5m6f9npYx5zBJb0V5TmFBygS9eIXHUBETS
43MJb08yndqMI+yKrD8Lv1pzwUu2egyudC1tMjKITHf8MaKNWb16nhH5EXtQFyoN
dBMVwRb/Tq/7rWHznII4ESrxE0p2Z0pBBAMG8GO+EPEYGjYBKtjVApCDCJLlyZjQ
qRL7AlxDKefPA9eV4cZrMgsmKvu7Wzm08TNoVw0jbzTdafXSoRet600AcCbDONw/
KOHCGpp3bWd3Yb3lLfD84SCNFhCsUGPGQSRxw/1q3wdSExj4CZizDE81E9qB+CUE
tfNz6YWd9c9zYryGIfQpHKhdxbpx6c+nIREZaG3fdF9YFd/GmmYFgZ+QnR5dYCXL
CUzN7bNfgGoJ8fUz/S05HqZbo7w9FuNJcYgYyNLVQJgETQ9ilj6Fa55ashFncqzJ
TmBCNcrcmjvGJ+jHzGXkQRRn2xspv3Lrfkegpx0bYIDbsUQFCaEyRutUSAD2GxjK
yPoqItUh8ritbj/hY1Xbz/SQyXqjV6KjT7Mc5Di7h8aEM7PjlFbs4cV3xdX50DWS
Uoi+4Wjt/VCALjiAu1c332mVPwqEBeZfSuIEc0fFCb9HCJxGSpMzZso0CPUPXJ2q
Px2jIRgP2cLg8cINWUuI2A6qwRrwzTVEpNLIvd1V4MT+HD3nsbrkmEPycA1FneaC
zi/GlAoegn0+xFOnIvlJouCeijYJu6RRtuHC4zm5rfmAOyYGRArwEc2uPY8OVE/L
6HXPaZlI38Xa+Ts0n3I5GfUDAW5UP/M3N9bkoWZCG8iloyXNtWxpJRvB1R71TNRu
YGKtP6UPmozb7LK6hk9kR7UDWrOMtRkEMJvxIqjBW7DwOLwp2OPb9cwFgtLlfcFN
7651/RL8UiR/fblQ7NezSX/IodvmErhwfNSXqOIqd5g5MGWbyNym77J1dcsLqPIB
twwnUC59t4snrEFzTNeUgazb6/05FJdhiCbrCmqvg48FuWH45sDpuRDOwZQZA4i+
iRlpuvZa8c7S57FdQXoMZuhKMxHZ9gxTPCZqXHIQUKEyFQActgBTY0TDHVs9PFwL
mQYkEaeY8v5iQmKLyon1/bH/rWk0IhqjXLMpDO95TVZlHHhDj91YDmTeA4w8cXYH
j4/30MFshUjtbc/Tx6GzM2nED2nhSnxELItdxIoLgrMrClblefFcDumjrXGxQD5s
nJK30sy/Lmo2JayV4PsZrZVoVxWBwu89CrS1+1dZpFQKRo44JbqvrqfJxHCpCnKV
8w9sUfyAopMPIbrsOJmUtjJLsA91agDABG1CHKsmMPA1lcJAHbniywDIwSbCvn3z
+38QKBxOJ/wtLjLYaLmCdMcAsoekikWqXmHsTl1bxkki4Am1HwqtdVqRUzvV6DNN
wyJCTMTyHLSZLh0E6Vx5lRC/y997+X1bd707qPU8sgKnEpQO6bNIKfY0FrvhFQSh
jPLhAIFIZG2XuwFOBLuzIr9heIVo4ledizgJwr1/gsAU01PUTkE8SOE1Cxdvx25g
BGB9yIOnPzdD4ypEYBPq26oVmev7H4ftDqAi9r9m1pz2u9dLIphw2DMlw+9jMm4s
/XOA/AmlmOxYCbYkcjkM+aIrpMYQ7m90E+0WWKBq7DHi1Zg2JqbS6GeKw1fwbnCx
hv32G9OLjcrZM1VnSBsQ0KldsgZhOfz2XN1+0zmj9E/ZCDXYPwixtEocC0HerEZG
MzcnIoFJ9Kp+Sp+gwmLdofh7XF3q/5GgKAv235A2V4oKUP6LH/+USkPcin+c6KZ4
/7L9jsWvMuPnXUWRWXzGuefsOPKSiaDwKdwdIT7S68SMTvs7IpIR4B2qKsChz/Pl
Im6ZU2MoP2l81cvmgj5IYSNlvhpcxZzh8bZ7nyEEFIP6RO9k7fBfY1WSwB+QH1AY
6zmdUpDdwL+XFkTI0UcTcg7PFVfqS1I6uEjUN8PHl7rCeGkbpZKxTH2NSwi3oSVP
Jiv/RciosjEC8zMUpppLE0mvDd5NS3yylTk9y8fMw/hNjAZM+lzS83n4GeIeLb7C
c11nBeY8zCwvoLbH5MMUunRXPtrEWiicKoqeTU+8/CIJKUoS/siXdg42gpiwZGec
nrp1hwzE8GFMBc2fAO9dw8UtWroi8pLINib4l1qgN4o9bjwJty2vnn+dF7P2avTf
SaMk1Lh1TxRAeBHLyfX9HyTRD9X6+uVIuZlUy0xEQiy9EjA/MLexfLlL27RhlM3q
AeC6gicIRQ7mk/3EnlaUH4S5+jKcJKMw/j0dEg5zJVIjM9YikBbkaOWqpImtPlRP
mPgrmLwW5e4awhEde33wT3adZcPxM1SKMJ0COXy0p0s0r23bCTzJqNkHn30KsFju
RbMZynn/A/BzzJxT8oNJKqwmyaPgcc99yYuzLayy0NGYJEAmTozXQn8jff5A5fWl
3SCESOZ+9cqvuymgmhBJd+wN/flxQ1kU+5AfR83rg2wnP8ejG6fns0SXvCUZSHae
8+pmn1Y7Rkp6l/ilP1l2LMIfFT18SQN1HcCbfGBkEbddBpkA3+HiBtGuVMZVZOAB
TAdQA/aZJA7W22krx5IS1str3Hqtoh0TWGUe76t2lkcoUjkgIUpXDYWxKCAMxDJt
hLm4MG05WOzS5rsAfYKH+2Y2vDfYTXZM2UW6EIfrsRj1l0xUhz/mrJDtGfDvD/Tp
yozMaLDjrCZ79RoK2nM+ZPZcZI8wdTyhF8nLTWYJULvx2N6BDYfmfxAeF1HpemJo
Ky4quLValnlmYwspbCxMQ6MZg6TLeWHYBr++i4OG+Dm9FwzE+APkS3WWsHOAE1du
R98d0wbyhn9hDuEFDToKSVLzJiO+heBtXJM5wvrHEH5MKa8J3kJGxuFzaDSLXSul
Aa6gl7Q5JS7B/2+7BIk83J+HJXa74I/K2VvPwK7IqhWmRaPpTbADUP84Bz3kHSJW
+dRDDyBWgfw+rcWOwvCgfg8c/L7HICc74tca2gtAPhtpdSgCoa9747SVVr4G6UUd
kEfKd8i0b4CaBr/QSrG4gF9gB6RE94m2QNTecA+wl1FFZ8Coekuy4s1dfFHoD2QZ
VBP3eZRUUGYgJ2McmlpnhRftG5YGmHUB/mnKRg/x7nsTGhhIY0j+7VgX/Q1pZR8N
sKucj+s1QxxoL5vOm8QCHmwDPjQtWn38oHA1k56lZRf39shSHRxJ5THPbK9wyCuM
Q65IvuugUH2Af/Xx34MQHwJaj9HmeM+F+gnnyadG28OUnjjYL1Obx9j9jMmxB6+g
Vk7m4riDKQ/t4PSgsXSoQbJVDmkD2/6JSwXlZ11r2DiK41Zk+OiK4UrPqHfc/MxP
eeY46gKX8ep6oCApGF2g1jY8ToaiajG3CuB4irMTgPezllsH1HaRueKNLCUOCW9Y
zacFYAK4cd+wWGBe9OPDtXttds7yfR9V8OCJQs6uXVmNEr77TmduXdQniEsYrpzp
CEbtflK4tN5BsvGotbnOH0whLWAQNVVaOhXOzd52bJGKCdJowgipKPZIa3SvirAj
T4rx/Ezt18e69YsLJxl3n/yGdtdaDlXwket+3nUV2jhgGfbY7o9d/MOHrOsgwBlG
XfMhr7oFZ42gr/GAUpsvnBmMnunfa7q9QxpSjDBTHlWiid9w8dQcA9Vtx+fmwNWq
y+X3Jy3L49qCW5Quk3zkJO5ZqIRKk9KJAxWiYdKDafc246t//jKcgVUCh4v2Nc+W
Snq5kiu53zM+fbyFoAD8gwRxOHijtP3YXrtcajfsB4+8RY1Qk9IN/W+WEp47fjUg
a4T8scISOcljBoGiughBOr1o/8JNUEwD+L3KDMKGkxK1HCPy4NQnF/MfR0gDW+6m
6Wm0JMhIBeRTiopqsNDZGYK8Cvgo14j4KMLVGbzwpoD1PdGJDVcEYZvkgZE09Gaa
dOkMqnLEfJvQLr4FlqdcBxvhjkd394X8WWyV+jL1H/mcQrVpywsZpS7tJprKDetr
L6ZZ3Oit1NF/iaovxx3HVzPLOagf91AfBKkw5JUSJypv+cz+AgzJFz01bQ38PKSl
pQJZW/wr9bcBRNGtGH7dnw21OHMQDGBPbJp8Vu811GIe6vYsTLntwtbxMZMXrVHE
bvqJ+boDcAEXmpoNs3TgJu/45qLYlthwTLFDzMDRU+0vN0RUSF1ofs8Oo3Ei8O3H
/7M7cACyYftcifvsZmR4V5aGOa2tgUwu5hU0UxSb2Hd7ZTUDlh89XVXHgyEt0kfw
HQlf95yRI7ovM9tZBb9AkZM3ZPWHwo7fljud+h/mi4qGTX8Sms29jCYEiGc0q78o
1I4I2ruJXdzNqbckZcjwUv38iTNMQFTj5n7jsQxWg1o5kTVd9m21Vt5mcAeBHYcB
ybGeOixERDZZ13tfgf+q1k/FVSTwZDLpc92KVQNbCQ8LBIKwmBuza6s/bh57nYU6
iPzgrGi6Y5nrzchKopgS0oxLx67KZV7xIK52mKqLXAibl+4TkAJXTlPUdDoM9GDd
4p0YYYUKgLDCyqOqRiRFr5UP/XJ0jcinURwMYx1SB/fOcxrWCRs9h8qFicGcnwqK
N8xL3fIYop+p9djC9U+NHG/fBYSbCMPYeFiZaDVgwjqOjCM5LMahr0RMJIvocU3I
T7B/VkC4FsrphCZ1U4L91rsuF9R1tXJ2jx5QnwWWFxNkFg/lCvbpHCrQzwVxFpgW
qZExZaOMVjqOv9rPE2Gw5OdUUrqT0MwBThNtM+BdIFXtml8/iY4qnSlW/qtwK+rZ
TPl7XiNeI83BHhLfHVxqw/qQsSSHefmiamwm+4qL+LLXwe/BqCxuPhw7lAc2Qbmc
UA+JTiAR2G9GjyzWFLno76gNzSazgl5LHCjKShKeDpDQyG4XEwrxAw+Ke1d++eKj
LigJfXFnkHuxSzaWMnmn6hehqf9xyDMEKjsBXd+Prm7SHVFrsrYylPElT2CFKs4z
PiZLYYwkMtw2dzPNVanjm61WXqbr/pdR3hDy5A7oNmT1TB9aSzEvnrWSiV9agbhv
/wwb5MNb95vo/4LtwnxauaDgXubBNDLDsAnab9dih+k1Vs7aU3EYpX6QapyyQ1q4
4AEnGNNMAuiWP/ShtjquCIPoys3XHizjXWO/rMOCwWq7zW7gQcH/MEVt9MjAE5Nj
gKHpKIUKSyF3A3+jgRpKHSfiHX7uLbYg3sKhMB6hPEwJKt8bL1d4qEKWO0InQ1w7
myMKflbAJwt/8IllgUvK6byNQX5JUIiGxCTkAJInC69UqOD/H9ia9HquFFzJ5Cjj
wm6s6YLHDIa205JYpc6mWLL+9rmjw3rRpJI2ZRj/wmU=
`protect END_PROTECTED
