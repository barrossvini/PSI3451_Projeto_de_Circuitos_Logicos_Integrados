`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uzzJVJf0FQeQEsCUL2hyPtDLZPn5yFDo/VGOjhTNWurgzMecg7IRTxnTi0sIp1Me
YsGNGIQdstsKBDPsF3qYGhwBiriKwllyzMBJ8ivTt8rhxIB6EZa7b3TxJbpBvj+F
HpA5wyTkd9BLQnLZKMyhZWJjJEtdIxzZHNt6yiPKJMJLtoUhvRezEpDrM1GGBuDe
xZXiMlmYWG7GWxAsNMig/fPvesCBD86kxdbdce4GKO/efaOawfb3j/lrbw0tVsgk
BLzzYj8AXq3GPm3+Y4tLbldozmFJ0kHRmzIYwX1hZ/gUU9CmZH1e/0PtK/VavTfa
B2M0N+aGOjYkrbkgVmfpon/hH0roPGWFQNndYYUC4+fvE3Z/zNs/xYMNjRTxHm6V
qC4KeudSl4BxTUH14q9Cij4pfV8sB0/Um/0+dL+sZjY3CSbyqAbeYp0mKtw4LEsa
whjJzJA204t/j4SROczhU7e5euZ2BwtoHnUW3c+VdUxpljjLZDGOTeO7wmj1UA2t
lz1BMgHdFJt6r/e3H+INiyUvkIc5JAF/hlZrxSKVKkpsdw7liPOFNUWM/hAY61Zk
0V9K9h6kq45IAIs0T57jy8wFdW/e5HvR9IKQ8iCkpushhsRgFVfRSlIVYLcFf2jm
vjQbSVf4rdQxUbu9XDCJeMetz9VnrfQfuGPXcl/COjrJe5/Ldri2a0uf2woeVIBn
0pvvzWDGrczkXDec8p3LUfhiH8fQcLWx0U6dP+L8MP6TK6N0Db3qHB93388XLzV2
2g1Rwe/QMQ5nprSmvQScH9PpwXc0KqjxG7uH5CSz6gJPmF9BgrSeNaEuoyC4jVut
eOMq6U+A51b0SsHXUoZ6TFhCVlEOnRmpYkQ9I2GEDadRpjRcIJqqOW15cdG/CnV6
shJiuCsn1qsX6jt+POMfHlr+xLGobMSmTVqR3Qszg3JuNQLeSf0APmLBHTP+TT6v
YVRbyBszIQzQciYZlvQxMlS9iDq89iNx6KvSrA2vi8HfmySs9Ay8nhWx84nu7xgk
2Hvau+lf0DiZhU+OvBPO/xJgYPccG0hAI3lFk9/8agfTRUm7OrdKCgs6ayP83Om7
RkQt7hPVZQ1MPX/+uThBLE8OQFFRU3RN03e4eMJgxotDkYcoXHTqT8mTR1Own4V6
+CG4EGVBxm2g/0hPAJff5Qj0Gq8S+oL0rG/mcyL//laxcQsHQhT0ojAQCAusZ5V5
SSHVUhIWxGl+LjS/DgmQvY4m0yOu00MHo3oY2YiSBKkwdnaf2v5fHLqDji3uOrZo
SJdzZem6Zlobtvu/0VJ2FN3TS0C5XcCkD4l3QOgXhI8p3iSTy/ifuggs5iG7dSVJ
3/OOlLZL911Hnv1pK7oGowAoKwbHRVAO1TmhgglJWGZxMNwvkOS+N8jrybnGnLtP
ueiKS1uaozu+pAg3YJh+wkrUelnQ/bERfbwFK9hP/9Z7BUw7aJkcpDnkSaZkVTLT
/d3aa2BNxN3X0WFPgTN42miW0QT5yPab4DpEopBc6iSofAEc4QDg8IM3pnNDVAee
7dQtNDr9Tw/N8hm4ZLmNUm9cfBdZ345C/P2LUVfi+MA+4oWcVhBQk/cwqAQkgpva
5gMPI9uaLG/0dndUIll1O8GbmByC3xy+KISCKW02dw/u7Ha16vDtSyVSXx3pOBDt
/qS3dAEZXtzfKMuUQ8beI5m4PpfkbVTvZG6ao88b0g4lYeyFVb6TTBG/WR2rB9AF
33uAAHt7DS2AAuQRD0GUHVe68/zptiGj6WNXiF1bOX2GxrEVfFovs1zxDdATCUBK
NQBphOUuVf83AmoERuyqgjgj66MNu+TBT8m6HRq+ENfggE6A87X3xpa/dX5am9uK
BINsHqCDc002a4/OOM8Gr/6Ma6DYxdbCf9mgH+tfnVYg8cxnFYVx16xALwR28lc9
70V/TRK+xf2GSQwZCby31tDOn1TRX6s0koBGc+viurY+d4DD/HfotrxtB/TWCfoH
WbdTkrBsNfToTP63YOCfJyXU2LvpI6kB6KLdJSbUGUxqNFPIn2kbNox1TDPlgCq/
cXr5vbeV+bWX4DK0XFaKjgFrX7hoV/dNl8GryIef+bRy65lk0/Pi3VRADeuWXasD
B2NgUDG2g1oCw3hl2h46vaXRbZmx44jzCKnlZiDGHZBfiAX/GVKAyC0oQLaAYhgF
aWIPwYLVMq9rpCScwjCryA/a9r78F4KrZyvJc+4yiuQdEAaFXqMBYi3S3S8S3k74
p//9Rk9lSTKeHy73yBdJ617yoMmt/AIcYMa0jaRYM6JivcTWDKw6Kfqg2NeFMfCe
jBkvqC97bSnCEy/d+5ZVZgAXtunZkoPitcRWrFPxjjooiv6H0vc3etTF/4Hsx7++
k2HYepQFUYJ4bwn4/qhEPvIgZmfFl0SImxkUHDUyHoBb/49GRhmVxGvbrXUepFWj
nFxpy0e7YoTNE1+GPHzwPEWeTnDG+A1uQCl9xohdK9qnnhD+rR9qE6SpgVaLY4SH
LOjbDjQXj0c3C2wyYR5IboohE9/VnBy/12qhH7vOgxeQjRvVapy/ub5lx0tihia8
kmx494uGzP0dNhUFOz1bue2C5IalSlC1ZwbSlcJ1wfrsKWwHunLj10aAMFDEK+yS
NMqHUaOAoZd5chaRZyvSo8HswUv7mbYTQ6qJvTkIdsr2iT8W4b3QKS9fx4nkZ6QI
DB4htLSAP3mWstgJH703O2ZU7/UdaDh5r3v5RiobztV7P2pyts6efTf2qarI/Hq2
tEa+HzV1ouvfih9zJGkdgdjsIzuTsrlNLDvJ2g8+ihJ0bFUYGjrrhQS4n2bbh1hy
gw+Qa7blZZZw8vnK4elTkUGwO9BqpiD/DMl/DtecOLMHu1HT0rAUvvSeUBIyHc/i
FHdLWM/1G+u3Fh8/J8vwx3Z3K2a6W9wM+S/0yuxhvZABOs8vqy0I7ni8dSYEBSD0
6ncvTCoIew2rDHxNS/VAFUnjNXr/h7XrXXRmLOHNmaU+97fGgsH3cgBL5QMSc3P9
ELM/RlmvdN1FBTQE4NR+1DB+9CN2Sl2SDH9qPHkDtcXDqxos62j4o1605hIOzG7B
UEATCwlrMblEQtr7gmTdPc6lrDSSGNmPP/wXKAD1wL8png7FUSdoq7w3yagixdI1
PkjFbcA4MX7D9YP0KWauGQgVTLt7KMse/YggBx8FuztMq3y7CIx3/h3lUY380f77
GizLnE5fa72ZCsCPViyfTnHv+HO+rAlTjvNg6CZfK6+7Biwq19tMISHLWAvaWXZ3
yUI6kvvPTNal9p2Ih0vHHpivo9oEO+o5Zc544/XK294jPD41YBU2hp352tjINYPR
YPR3azF4r1v0khMOpN0B7Pm6icCvlwPvc2IDdWSjrvF0FSlQDEB1O7Yp+SUCZZ8e
LH8R25Ovb+kS3uc6ECQjOSpw0qWZGs4lPgpAO4/Di764rF44mJMFifU5p2B+d4sP
So16WsOUofQcuMNj1YP1un39rq8k+bRtPMn1LqdeAbuwXfgfON5iM1+wNlQLU4XV
01DasY/oguveJNDVM4ybyOV3artLwGUS++LHuu278E++jIPNE/C9FasZyMEuXcOA
vKdu+aYBMRSIIIDU0Zp7JnI0SKCT0nT94EwiG5IXYGxOssZwp/MmgfuTqMKfLiRU
h4kVLTYGD151g2RYPTg6/7NwrE2GUBzFa3LndMGg0Sc8WBq31jhjH9XSj9X04o2+
59OaXzLOlZ1oRA6SHLx35slHbLI+x396E79o1jtoTruFDvB5PvvlQ5cmrlmw97GI
icPXpvIDSsiIuschPBJ1ytca74TrwlcvJo584QUSEc0CXBMqx2b1BW7UPkhrC98v
TZGhjGS6NWINbgwLfwWZtWjEomgAo3GTtpGIjylKEYsCjN03qSS6PzeZdVabvOL4
PtWNQcqhmvARWszbDjeEB07NfVr5UbnwuEXZAG5Ekk9KYY7gPwdZWHooC55cCIpa
/bbn5vRWCCyE+h9UsUzxWh1KIUs0mHGEjOc3ifXOZC4e23vSXzNtWByhip7iMACv
TfqvUlODM7rxKvFLQE4N9pib3LVIZHR/yBKmGreL9XvN1yl7gZZesGV31rjA3imo
cMNjsaY9jKoRRvzgXiYeeVUfU0LXO4QMrEj9yE0ebZ3mCEziWkGuRGOiWZnMr/4B
D+2NCGdFtQKK8L98pvl1JYGbB8Xl1XlxaCyD0cRvi90x9Jq++qF+Rt4l8a+r6Zzi
QqDGRtqHkCDaXG4ToWIq96E1pjdmbfePs78ki3unA+adG0G4Sir7IRC8ilODopSD
Nt60zoiQzlHBtQGuhQuyLFbNOkI+sylsd+5XA+XAXhW3ZQbDA3wm2enTm8RDgmWP
Dippu37zx/l49P5Loal2yCyv0l8MMwZnThT20+wdB/U=
`protect END_PROTECTED
