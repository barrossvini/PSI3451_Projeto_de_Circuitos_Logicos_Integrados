`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YSViNfuVbANRcQ1/U7j45/Ij2SVu0RrebTMleuAbAbzenSDrp4zWdSb2EkOEHZjw
m0+moJTMA86oK4TzzdDL/lGzgE0GSXOHLchNOXxkmepzL+e9cFaTaMzxBYtATqpU
Cs0Ce+q4Us9lTXKFy5BFqlvM+U0BN0q2r+hXJ/9uKCoRiAeilIRWQmlNEfSXZaJd
pY0Ad5JegCe9WRDNDziEGBjuB0NHmS9u/DSHSR8oCG/PwDrypAlXWbSlSZSDKmzJ
OK+QBXaW8KCZSB4nbEYgrP3onJyU6DHjE8MxHLgfuyn/jmdWDGypYdeEYeYLW7Hw
g8R5WRYiepe5EZDTXjPqw02Bb0igU04+yD2yRgel4ebEVxBfJ8W8H6SwJ3XSShUb
NnFNCbmx4U4mmhUs55FtX4MI7NCwagd4xiex6qNSH9unlaADa2miwBSdNsmA+tDl
db4vV5GEet19lhK+LTPM/EqDWGZsEnEkM+YAIcN9UKHI/7erbt33n99AJ99TjAEE
KnJ+Hb/fPCdPjCd7PQM7y/e66vGCSqWf75h9k7SdDnAATnA4dMSJfcRY1cwT19t3
bphmmqLshS0kampU1p0R8P//jKMnX+CHls0SQvMcNDt+ss7I6jWrSbxnSX35OCaL
AtbOSM7kjEl7TrXZDVGTNrU00FyxPGNB3WuafsVRtSL5VP1yBn4lx0pe5DU4ixDK
Xyi0Xg4fsKRWx/+3Q/4Xwhu67OQoqHnpzlsR70tttcjhtiwFc+dY/PhLAQByIECB
vwKXvX8l0lph00+MT2kOkbEPGDqfW1I1iFpgY1CTVySD3QjcGAEQYu0du8TsX6xo
CYJsQQu0dVXk4F14Fk/FmtUAMs43fzd2aQU2FYansqjcycd7OGbZnbTsEPgaasoC
NRlTFQiVnzKNbjL52k4LOYS64vIKrBAYunNtcTWhBvLV5PSu8bz5TrAnLPWfieh0
W2bup/xGy6Atzh/unm3vZrOVE5gDd4Ol5y4ZBR3kOJtbJ3VLE8D7TGsoXMWvWRMt
S1aC2BnpupDzYuMwcrD1qnLT/9G0J0GB1zy75Syr2MewfPq9HVyMXd5KE6wUrjDS
wl82pdffdug8JolPlnp53VsCKtc7hmEaqwdMC/vNDJdUhZsV+zjXjGsdG3X0PewF
QdJC+yeGRkvBBBGTkd1Hz2Vfl2Sl9x5QsjnWGVOFpalvlqcEJ9j1faZpvC1QE0H0
EUAsXAM43ZXylQ9V/7iHkvtp6J870NpXCvISlEFBdzouKpkt/6XNJM1pHlQVf0NB
DA7W3F9gFgL4XlLchKO0DC5tZ0CmdeHQo+SLaM1Q1cC61dMWyb7agqVVMJ4GZ5aa
Y7mtD6mxNRc6nve02TjDBNu8LYW/1Ot5C5YANE3WgEL+9/kK7RKUXg8T0JtxC8PU
usAmMz3Qovk/DYInGdKRr55ri3JRkeistXzy8f7sX4Ew2bMtTMGY7JMqp5fGD1kX
sqB1ozGAbl6VlijnGBTxhDghrZfWYWPGK3fWE2G0MeJjnDUd8YsI38RghqFwAp6C
N6sbGcma+wKWraWEhoX04R+5+hyPNfRZu7w5BbAMdMmDKlwjdUQ0bGlSnwjJbg7c
Rq3Sm4I+NIDptkqPZRljTk4Mh1Pi/dLgvG4gCFBjb+nWRyBOQmLyCLViEWgkWtXA
Bt9dtZqpdCMTanmzLcIbLU1HB7vGARfww7LtVBF1R/WuQx4PqfCCgfCLdI5wv4Yy
QwS7ehpmVl/5vlTqerze8rt/wfoAq3lFdt3bQceDe0n/dFXUmKscg/N0gzRYVrTR
TnaaYFen6cWlOY8VwCEwF777rsdLACKFmuOorjeFPWXAkm0TubJSoLHGJHU2YgoT
B0OcI36InOg2PbPjXXC5j0c387y9qXz2UGzo9AeuQap2aL7nUbLKh9bDEn2gY9MY
w8oTwadUHJwM/+JmlNFmiQktCFrfTyZMX2JcIEBKaGHgpgCrexZ7webDWQBvBa7S
S0GXZ53GsdilnIiHHQaDWL0RREy/92V9xmxer4SQQxtj/VeWNlnwWMj79sWRtefR
HOrmyZH0DAeBiRbO9+Xe3Xd0FgN8YBWHMXuP5ngfiQrV1gZOBnLtJrihF/ihUigM
eb+xQRQ2iWKJi4NirvVun0Rl78FPQwSpofrw60cf4t9TEc13tor8gx34ojxF6gVm
R8VHP69naAp10qRXyySA+itZsDu7XNfvXOoE5lO9NDbXN/du4+oRxNCr5oHnenme
6FEkgbPnH15r7Nv0Zg8Svpaz/8O3t7nRk5uGA+p49ZSN6fklPbkY78Bjvo0ggIGW
sbwd5taiQi01u5qWZ0/NenFTAwIODQa+fDGq/TDk3qXOWgVms/0wDtDt1klNIHTl
gY0qlKSXqhcJAJD/wKPSQXEFhPfU8muD24OsSZX3vEr3J516PiTnq+ZoIldsoKOL
8cnGBuD5YA5H8Qt9o7ZkhQIry56N2MUyMXo+LCUSrjqOgxl23x8eCsxfWoGjQIZ+
S2J7//3Rbl86JXs9vPX1cI9jtRFi2rftVihWPGsoYPAqYbxbTEdDZfS/Q0WAmb/E
8k66oSGPHw6zn2xik5RLNuK2mZG3BzUqGi09JxQM8mnC419WGLrAXpsKSdwBVOuH
yz9nDwSrinTX7ACUZdnoNu2uPQbq8HP1gRNh2NgG9eK8IsEIZbCCekC2BWd1MD70
4uvYq06Beeay3uWTAxw50G4JABAZ1kfbHbr6CUcgeMBAgcLNj1E5Pir5Ssb5RU7/
/0R6xXaTTqO4+BdSgK2DWe7MVEy0dQub+vy/ar+1j+pVZdhH9cwXMBcTDn+3ZQZE
TYJrD6smd7JsoFVnI2Vds4iKHPs0XkFrSGEyL9neFSZ+Mp0t0ANv3+hJZIhdGOSh
FaoBJe2adMv67ma0YqxI30H2p1GuB/aRyjn/D85ahO//2MOwNSWRramWBT5mvL7o
y8MgU+uwAFKHXVjKyHoi8wIwUydjAFLo4PsXdvrrxNKrTIYCjVmCTuHjEB/zd1a0
UBeIIyTCxggkuJ34mY6+l0cb9HSNeG6CuaXKearOgLADNfOJKotW7Ice4b8+Jynv
PGPE6fMqFhhPx8hdNWNRZ9p6JFLn9/eGwHJDIneyqeT+zzjXEZoA9OnWk439P9dO
dETUxueSFw0fJmnedwx2IcL00vJxp/lYQcDqIB8a+N8zPgDKn6PK8xA63cOjZ0ZA
vrxlyE/bqw3x2Is5dzqc5YIEzBo/QhlwJv8PUH27Y4lqQ9z+8WQScjaBoXPiG2hz
DtYiR07qmRkoWm0FnaFPAdDg2TopdrzDBh2uzvww4gs+C4vyBkIRWkaXEK/Dt10h
Pr77kflQEmCIwhHTmBHLoEV2dgFtXRX14PvTiUhjkx8XHri+mlyEJhZKlmNmptsr
wGZoh5pocDPQUtORbtyvIYddhmEsp48PJOfI8TUWIDvGM4yv8Y0UzTHOF00u7tod
f2BnPN73Rl30Uqur7Nwyy0MMyLYVFac66OflpktDdjJITF6waCq09U0+hd5GfdZk
1DbHgdAiW/E81acvGAxw01uysfm/R4IHETm0zLG85z1hzngb9Y9q3ep2Kh2tClMn
ZYcWTJRTYLB8/4C5oC5mHl3Ru+xMIfwdNai4ODEWrt94ewxRbLb5eubHNSIrucW5
ajbAPd0dIEQ6+hpaZ7ksInzikY0szBxdhwEG/4XtwKexu3QSlj5qHeaqtpRUmq1W
p2uFvvVF7sPKxyBvQL78Zg==
`protect END_PROTECTED
