`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
veJxCgdWxQ0j6bFykzm4rWXS3RUHuFDVfhll5hnQH4lD40V5gGx8Nzu8kgw6peKn
5o7R2YO003F8K9+5MC2hzBdVH0UmpxVFjyNgmhdcND6jHQXKtYX+KYkbmZJLFhFG
wbXfM2cmFCEZCN+5UijAUN50H3ex4hWYJDXrN0qDXacob74ZUn4vwWjgYtd/g0Oz
m1asCmArNXS/y6cQohizgxKgnKvwiAbmB00NfQlHbzHdbVdAUBw4JZNqg2zcarPU
bH8seaePhJL2gRrVBKqrBh64LjMdK7lNuCWw9Uw3/nD9SuMUw2JH34yF03uxdEbB
FLxIa22tHqoScVFPsS/jU8lXhY7oRzEkGNY7BPpV5ewVEsdPV/iM9YpPUZs54Zjg
ar/KWmvXzcBqzV+03BhA+C/6uU+hXLyTevwZCNe9PtsbCNEZmjLDZFJ2C6+WKAR9
Wk+6+ZePTbwdfAgSTDAmvASHXfz//ZTCtDmwICSP+shVixRwbaqmXi+MW7MaoZEj
uXRE54ZBLZJQMDT+sn7Nlv0izdgwq9PsMWngYBIfq7g6ayV0t7IZNyz5cuouLnNa
edHS1B4YtDYOKualm4bEJYUUOAZcFWgCnR+ygBxpDZq/3ruuuJ68USVI425EHrUI
r2A/pS9OuX9gdSWSgbElsq6NGp4EsMNPXWR+wEg7jyeTUsUcVLBwe22Yn4VVKeBA
PivjzGIfrPgSK7hL/Bjuzkxm5kYatdaHCJZ/X1GEfWrzjaK9BdH6kBdY+opMzk4e
5SKqfvDtrN+AlWDfATbYbGCdU+yWyu/Mvm7k23rmN0GJACHhaWnHHHZxXkopgLEy
s7GEd2JzQ4OU/k7NvJimZR1SuVcCqiH2pdinEeX1QDrnEE9agsQAxwjxpGOX3UUr
7f4Qxddptrswa6SB/u5BBaJHVPR9e07+dR5p3YRKBaoPgSIlVA16rF+r2gzex6Qa
rdZx0CmZYe7fo2tfRwKpTWSBPpv9RRP8r1Jk2a02Esqhf5IIV1l3RRfYIoy1yxA5
WcjFSZJL1PaNzCVG/iY4kb5uUkO1N7+lYv1v3TtPG5eo4wY46Gh8c3mBzoBixdpP
79mIl24jDPOQc/UUx/MizsJO0IR1xP4SZN7hum/g88gswHDyiV2LAF6PWuR/h853
qxFuff43L6EBjTF9tIwnOgzZNq+9O43GgjVpQn0QYYd/jXyIdOa5ak17+NEw8xPy
RBQxgPewFwtywLx0WCEYE/TqUp18eiYg4bIercQElan5w2YlabPThiN2SzJULYLA
2rvD7TFxozKUqpgouTtif0LhQQYuBSLxOuVwUkK/gp8JQyc1c8/D7uJxb4pw/LAd
RaPtXHbSmfQeyTbfdy6ATHGdx6yLNORa9NcaicehvmfBV6XKEOlOB92l5Zu2Yq1Z
S+rLcfkU9l33as21SKuOVA==
`protect END_PROTECTED
