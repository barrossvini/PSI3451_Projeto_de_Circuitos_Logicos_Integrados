`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vzqq0JHAw1No3gbI6b6MWD5y2SSsiEAACkglMlSTckREmJpX4hiwZd1ax7ozonmX
Ywi/PWYiOb002LeFXBvsCPcQCza4Wvx2Ve6yJQf3QUGXU3tIntHm8WqId6IeO0i7
G0jZ2BnpgzXF927zNKjwqV1KeiYti7eKe5XVVgZxLGY2tf5p/UDMqHj++wVAfv65
dD+nWkK/ILgjRb5dG8AE1LywzoRQ4EfB/0YrnRo6Dpp3rpfFWgtFtobytPXh9NId
Uv6A1NDbpw0Kh/MEiXdFyZjCudgvzyrm6n6BFg60F8io5AiQ9S8sZC2Bm3A3nkqR
LWjnzNqxN2sCn9LpfHdKd54kVi7KXi+qYs6GN26HVGuKl9w+JYAcbw236QUG5QVr
Gdyk+jF0/gE2X1bJDw0RYDc/Dq0AK/3LAA/IEe2BysBOFWpc+QToDrX/xm7vUbMx
h5UNLYLTQIaIuY1PKs6GshXNB9zSCvYxPTfqgQAjft53uqZxOkhC6fpskDyTRH87
NxXJoLODJH8O5MyOa34pXR44IkVgNmqHyPrQ2wlga2gcUhY3sZWdrSxLjRFg9+NU
djiqGFPMqOATQPyAPFs1lsBnG9yBRYC2WS5SzZT1USHmZHTBkoTTVLxOL/lOAjMh
3UFOUUl8A993ZkhXPDMg2R0b3FWbzKmhVAfKpt8JsGsU8xrslcoSDPJMbzfvejFS
+WjjN7VPKa9GfzbHsK0CGVqgE4OTHiC0vsrB7HlyM8kZUAyM+Dlhy8+M6Z9pPkeQ
hDm43A5zLugA3DU5fLsUXUU2fSu/451rbeisjDHYTZCpOP9lqvLAmZ5E3gzBj708
XjOGYgkpD1haQdM8ReGOXGx8yqc+LzGe0XGRNkdk1+Ae5b2lXhg1vraW0BE4ZqZz
yM79+7kLMG3uDbTshIb0QhPFsiOnYWR2C9Qg3DUFXPMlwJIDD9wCa9JyOW998SIG
eVzX8/avoRsbawbZFS0dFshS8Bw0EfNJqYxyoXrYHQRiKcXJjTBDu/BlGYZ4vwtF
DUmmspJSg5ywaIpDdXzMj2f3f596tGmTVF6k0FTyhylCK7MC1NCXjvh7F5xbSbm8
LOojZ/vSUjGwLUCMGiyT1MmqD81k9/d7HUq0xUmj3Hj+7j+4RmfeSC8Et45paDL1
jmjcJBPpthyh5QSTcNkm/WX22eYKnmuMdb+yRbgFayET0DNQOX1j/+CZdlZpul4h
jZoTI+/QOtVe1NGZtTfzdG8oii6uJ2IuS5R5ib2O5xqpF+Je8E8LU6tKE6ZcjJ0Y
mY+d0qTX1+g7L0s0grJOT+qTRe4aIZ48+wG+Ubp3EbYJrFwQJ6BXREJIzKE9np9E
EPRSLiFycDkr7UL4TdUJoNMwoLKKRREBZNWQbZLfu706fO/O7HvfrJuqWW6c6MTD
Y3Q2ZblR1fiKEdqtds4yyL/JEFE5UpJ2aBqdO7NXjKgjOixRbGj3QskhQGQqUVnZ
uygrXmhmkhQF594tq9ox0csCNG+m3Dgzefvgiy+Ma19gQbOw42q/pEAT3OCDVkXd
iisIRnhfPIhoa0OBzXX/pA==
`protect END_PROTECTED
