`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4YtYA5G1HUG0rWcXFTS3wl6GaOjGwD+t1Y1UF8ZmUN8m+P2gDkz1GDOkPBEXVSmM
xihqMOL2Ot4JMok+TmDYJ2TVsEErekrW+UlNdCxA0zbc5d+sWGTrYgaj67wwSkCG
2rg8E7t1/B4sFEFV7Ve0z0j/GsoJM69ePKzCY7Qhb4KH2mJJmnvYB9Y1Q0ubC8uQ
iAD+G3O6AqeGJONAnZixmsztrHxucu6spR/WuOTnIfYvkGSYXgt5gQjCpN/+Vuus
w0LAgR2szrOgZ7zovAdJ8R9h/dE+MfSfmv3rT9B1tF4K5CjlHANj8I2xN5JtlfEn
hdBzvVRoVmaPiknVlMpFQQOo218dIrdMCX12vzgcuhGTG13vCCP5xJsuHIu6Hr8n
+S67KwNIWYvl6Av+fTH/vad2SK4w7keU04e4vAiBCrIQlpG4wySiZ4VCD7xgG03K
kpW2kH/WIYsPxg0jqY/ZzCb4kJngDVZlu8H3PoxbyOCD5CuQSAnCu+vmygOB0pEI
y7BQPp0tOSxmhvQh64vYKaau2r8pIeGR6mgjyCk7Igm54lSppQjLTGR/QedPFmj3
J9eU9+J+mDcYFVOuv5WAJQIOK2PMEIjxz7UpfQTXyrwRAgH+9b/pKobXpO3KbJ5A
eiRFMD/osTbYYdAnejjWnFqJEjhjpu27LK2DfO/aVagnvI1uE6MOCxSz6nbry47B
XvlT/RYcaf28rpsT90OHrnz6xm/nfWZ5SpYpkTHXu30Miv341WwQAJqXGOII1YWt
cRl8aFE8R4tl3hALpSuFw90Um3XrBITWVnPvBhQGLHrSC9509RJFCIKRP3i+0lz9
IhiomBQWB8Y81LUm2TOChm+0/b+JKEMlbdpezwZeOJdvRGIIlUWf8WSPpTn9VGsJ
Qz3/bdHAa6nNNrvza488quoVgR80o96EbK0NcoEIMoVgAWYP/vEabO98tYKszv1+
KB0pB0OslayPhd+GU2af4oCX6gR+6CO8/WdIZh2dqgQ9iOChWsocmCiZC9xEQwdY
c6juM5ZxjGAOzCPjzyKZKgghYtwM4AmxTHa/LVmjUSKeTR/Np/8y24LZ9qjhTL98
sK1//T5wyrfGNyrbs6IMRFnfYf87HaN3pcHoaMykmJjQWko6GqeGoSv2Qv+/Iy0y
vgGEUoLscYqYEqwvHCDqOUdHLugvz5C5jqy56V80Illl26T8RSClhAUirAiLkOuv
ijQIhG7WJunrJC1TukEXZdgzlmBy3lpI6KDdJjxqqnaUqDDk3ViQC/wHt1SEmb43
s872VDgTwtlD11VlusW59j646ARQ4DmcaQuiyTs9f5akqCfg/IHBgOP4TxPhhdzT
bUyEO1m9yETjcSyQKeir58nZhmkZE7hkr+tpV+8dd9smoLVXiENsEeMXtfgcGx0I
9w9ksID+LMcjz4Vmf/ksBiJzvAnIUyVLahvfbRxrqCjEnwLEFDwSNrsi8Vo/E5Y8
YB3miw3RVqNqtpp6PhuykqIO2x0lSOKZgESPi2RdI8gI2QPwD/lxEmf+yNARo4e3
/x9dJjlpnsj9bESSgBhuOk2axttdTDoTbW1zy4M3dHAc3E3hjmGizadVirWLizhx
9CIgEmhmcMSXyxD5xCCbUlpwdo1t/eduQJ5O3pQ3VGidEg3uxzVI76LgNbMNaeBQ
IpYJTc3Mt6OWYXIElRiWM66WhFwC5JgbgV3k35eo8AQpCuVDqw4m9EmjoJeMgrc7
+6rmPpoCY8BXNWVy1ywAHBQ02EdUsWm70M/P8Sf7GXAdb/rENdFxCvm5wu87Qcxh
zq6j4du1jNNl4XJiz1+lrlDA7+87tQiRQ0656Rhcc5YibJJAMe8XuWa9vQJ2WZ5e
4wzioORJDOgvbBxPCHdQ0FEj8a04Z+oSCRwSSA/RwbSrzhcKfkeUz17F4IuYTYN0
Zdp0RXS+Wjg5w5hoEXYAqHx19B2lsA+5SeroXHyyBofxAkOef6DeP7mpntKb8ZGj
R6jkHx2biMglylPTuRabQ2mkA7uyWc+ChwLQv367NvHdaxocl5n/ha6Hxj2IcP9H
7cItqmAPX5MYF4xlYDBHtcBy+2y9yd/dUt143Wve9apuT1Y7VMG5wAV7EAJO1shO
9q2j15xX9aFqbElUbnWMVI5pA6NHZYpF4ZJiJDCsEDhwpfa0PJyzXDjcsD+Dxea5
EaoIHwOqTpHQa9kMVbHhFKtaooK6VzKSZ66zJ82FABh/dlyh0C6Pv3a/gmcEbGxq
hUaftY+jVHwjgK4oX+KasUfXe6yZftu2bQ5SnyKXPjXIqTk34NW266LtxoB5VRNP
OdJBDcY7L6ZJCrmCDWywaFiS4g5vO6lqzi0sSKO21ud4cqt3OY5amXv7rR9zFKGc
3dvjDXbZUiJ2zH6DJs6k9TexyuhsnwKpliV6pxR4W5jDb7NraV1rKRSj09Nqfk4f
iNJfJrthTBAMcWjctnkW3EXHyCVdUvqBydXXdjPqw7v1+LYj5P9p70UsGZxgYTt/
vrJalaU6y4aKl8KA9lk2J+NVV9CDO5wUs7dCGnkB4WSwwu7IPiziyJJPhtuhhe8C
kELj8AuFqvxlrbVBkmGNjv8BXtGv++fW4RWIs07nTxHwzX1TsO/Wne+6kSSpz1ge
tpUIJdOmyPtMbNZA21dfkg0jRoWhp1DCuC3gd7D9+mGwnNyttdlIFcRFYgosrzoo
RgkrzIxxZjbrOGw3H5z6z9rUoJPleITXwxPB9g5AET1+rbuvtv3ytBZvo65eMCPq
TBoqHAeuCyQFPoqJKaeJPOX2cKzSmUwMRWJd37NsTsXmOOfnQrwJfAUINnhjew62
+xVt9FthgNK6aY+BAA/KzzplUyqYVl2+iw5dVCANYgUg+E4yAQY2x1DvgGZ25iR/
fzbi/Zb9arUgCXzrlOY60xfwOfUvWzTvmGVEbsCS31M4K5YBYGGxR6hGlky1cqGm
Ev+Te6LiSCSAYjzmeG1RXtMRct1qiL9fh9sCwnx8NxfB3wXeVUurQfhxpYI3LN8+
y4pxVU+PTLt6HXZOq0SOAX9PyVaJFq2oA58hVjWcUqsN0IrZ3dnoM6IWtDSFuBb9
hl0s7AzqhZrzbvLHM0i1Gyon86RQobBimkdXq7IXlJSz50RrWUizvJJjacfZ7aEk
q7QuupIJL9uw0Td+KXsrFCOgvz9qas54jI991GIvox/KWX0lTh7+YG51sDuVsQcW
sFeMZtyOxXjSa4zNTnJ1XNC14c3OjepXCb2YuvB6MDfvoiMoUdEKv1TscBJi/8Bl
xrHyGj/KnzwEX/yg0cX8x8BHsVM92v67PVvIJ9dyYNTcVDpbbHBkN6Jg+gtFMxOF
m9s75v16nmyPVCSs/+jKhqNOXaHMPe8pEFS9eQlffdmeQOOeDrpVQMwubix+ILxP
OpoHGDwimjfw6hnl2QHXdfrt/t34q/VxE2HAAql0MedjhOTCCU4T1WuphQPDGWoH
nsD0mvQ64ETIIH8YPrH/ctVn4D0IvCDsm228CjzDZQhr/r0HFAvNoipyCrJEO4cC
sdJ4h8/ObQFSKAh5jCq9net/lgevhgyciDkirlikMQmxEiFotsGY1a2wLwt8oMwu
V1CzURWfA15zx+JqBNRmn/EmkBqScs379pvhey5hpoVJCAYM2sQgffTVoEU9Gdag
XWaWXwBShXnyDizOwJgEpjFiZQ5FNiwE8aMZdz/MvyEqs0y9WUKBYnjLtJ9rW7hf
9G2diNk7SDkBHOTjNnPCYPfGexohMFgk9uy6oHpHeBXcDSqAlIF9Ibom7nruV4C3
Pov9d9sM3UU1hcHkJqSlrz7bfpXyWdE6afUWYmy4oQdPGdsvQrwkOr+T9FxfZDNy
n5fHqkQZ4lorDfo6wWIRheCCk0B2Ccu6caDO+p1/zqOkctPRhimen2H0en2fFOc/
J9o5NmVv+zw/vr4kfwahiT0AFPvh6cFHJXamPYqQgkSQiIlDaGFjY+dOElUqRs5L
gvSRIOkWIYhDHZif9ptQC716fKXN8HQ/3OQDmBc/ewdkIgqRKjfvifrFkLzU6248
XHQ9M0Jxix9NcAYMh47+LlAt0S+h2ELasX6TCB+VGqfJwDB1dnUEuaKvt6jhIDjt
IsZV+e7mKSkAV2u3t7tn5JmwHZAaRrmSEP91MTXSaLsDBEcB1PzxR3H7U3Wq0r0C
JEnTYEnIEH14hgU0HJ1iwsyU16fFar3GITCmeWVDl4e4AnwORhOcpwvkrmh/Hjwa
6lPV/EC35ZO2gHU3gVjfKFfC7E+Jo7U+Btpb/8mZPpQhF40TgFstMkubhfizJTqh
GqQt8CIoLG//tnk6loMZ9NBgXdciQcrHKT8C5EFYJcgw0Bt131SIqdFhiF5RzKhF
jEcpoeG/2+NWE7vjhcOvKhmhAVXXUTLu5IOhLW7na/1i/KMayk+VBcqR+g7lmzfN
5mzJ+pf+y+drFVzcL/9md+qZAZ/gwTVgnc2fmpdbW74jKvdDNcVWRE1FBZsamwRX
WQaq4uhNhxaUNAOOdUjbmpyLinUNfIlJ/aLRDQIAeUHIZH5K6HEe1J9nKA/+orYb
I6hCp9szz+ezWThP+nDuRFi4rsbOBkYJVT3Vyz0rHsk2E1Z3KUxDqC2wu0gPZVY0
5WZmva/InIiTAwcwwkdokfkXARWYMoA1v5Mbmg8jbmnGo5kN9cSMkhmVfyi/wb0r
2nJ/tJFoALfabPCnDi+4G4GEVJsdgPeZDQltQEIsz8GMYA6nMjbFa8TZNjH63hN8
CDa1fi2N2u/aLsW2QlfCodzchJTBVeAz22OYTODqhPVdiCAbLnGul8Q5pgbZzPoc
2g4x+LcQsJAvl3zAKdXjb1J3d3juC1iXQaeiMeGIlx2ZPLkRUi54UFulTmpxpLmW
W9iivM+l3Yk4PIcQ0PYyRv+OjLgx91VhYTOx7O2gtn/9MrqB7SoGKvTrFHDa0q+u
g1JB/KQBz2mw7O6cYTXPU4b2g3YSo8jTYIgE7oagU2694l60dbe/41avl77p4RdE
2dSdvjHLcopkBJDR5Tl35ucIEWZesl6joO5mZb0bIl4fquQCL723iSMewPj1sCwn
xFQvMkMotdZuvMLEapCkcWm7TqZ4XsRNX7Gx5exmihMExPXpFwr/Mmffb3PHfKFY
78QLjULrG4So9ZWp6VP65y6avA1sjfMJBikNHTAKKTMgAfnzdEtkJIpWIkpqK26+
NSpxWPF23PzjKL4kCqa0qUrcD3VuF2dwSo9fZ2RBx6yDgbqoTvE8OeQHHUQhmQ8/
UuNiMbuoGzjDMauu9Mo9MjuMlG/iaVXw3Ys9gD3mWafvYL+JkmwCZBNIdIVB8xaU
abRULab+uxk87PqnGQDYKMYELWBULFw6bLR6fiQ5rx785qQCmaMZqCNP3qq3K4nK
MjXFB5EOQz2dVD66u2I0yJaL0zaSxLFU9/BbHPc1Z2hurtEue/vLmE0sRtIfx0uj
HvVSXCdUn/mTitVj4VM/SjNqgKvUoGeVTPlSfIRRu5rsvBVpgjars2/Icb7ns22q
RSKDzRjqkZStZUhsUL1+A1cRpfC8bL3jCDwgff9sG2YbYznlz7qs91mrqIdqnuHr
G7jqPGSOw0F7nHoBpjMGNgNokGOhhDDgCGUJnAFPBk9tRgNAUfkh1S2MNWu8kv7P
XUx9T+UWf4D3B3lTfg5p1ZFlVvoXSUhVmkasJxZlsbRrKkgwY+A27PAOau8OPqpm
AkYud008Y5/d7tJYVi/0ZjQQJKrfo7pZ34RnesBrNbwUmIDOD2uysTgRlQsesPVn
5AqjmttikMLg/gfLAxOgI2zyRndulypSJ6OEHzprzyStLxZGlBzwLCOopsZ/U0LZ
LhYKW8rFWIlHR4ejh/68eAqtGpeoGxFuwyjm67Uaq72sIJ1cnfSghO7tscj9vNXf
BPftzViigG9HqtGUt6zRGGKK+uio6i8RKGiv+LgKXAO9IiVFEtQtK9fjDWnExg6N
DVdzyOjeLmNGdeOMGK8/BdCItIGLUI6dPnWUj+n2mCQlQ7VbMQKlZEFxV/pMSMxA
EKgw0HgsddWla0B/W8AKa7OHuJNwSfodi56sgY/VmziiTkkQlbtZUBGD03nlRNI5
pIK2kvRzy1np/y2Q5dLCKzNkXsPMp1fKymiAxG0xsTMUYcBTalboZLBoRbI1o11X
kIFhdijvqpreDfNzWNdSWoL2zoUAWRgMAABp2xufh62hg6nvkCRkbKg5rPf3jxRu
c5jv/adTB58EwEAvMZwwkmQowQl1Djj54AuR1xRfEI/X6WuJ2SGgqeM301prrg9t
WJjcICSMPSU0mJC5Egm/Pa2mBn+3WNA70HfoUQTWJKYFEm+5YCXyJkWsN1+cEFev
96nzGFABFw39DtKYSRgIo7B1NW6v+k3WFsEajINM/NV2P7MoYk8J080DLoNfl3lq
YCocYC7QbQ9DBh3aKqVXAiKhxL+C5OsVd3ioD6Z46wU8jbMx8o9RDED+GnZCrgu9
6Qdx6tBCWUW8kIdrrhdqW+77DPlFCl38df7tILKVBICzCT74HUuH/yVknhSiDUPi
wa+MEOxSprz7L5XHXp043EWWiOUDARiRqeiH/Q4imnDXpX91hKMWskTW5pdHEkhn
VXOR99osxtGHxwc+j7utiCAB/ZK8yTAV3GOhup/FmTZXvOIVZIglvoQUXt/ubm7Y
pcSTgqaTCMJGYt+f4532gvRbRgHNMut0Zm59Xxe3isSZKgak5n/Znis4PbGNyk6D
BH7bYwI/0jNfh6vUN/d5/V1KAOPLxSeBrO+Xuo3vsNag/VRNGQowWo3KxyByQCki
rp/0v4N4/LBzh5dT1lKlx9Aj0aC7u0LA1iYWws0X9N68ZmTOrt+ZRbW4wemJdA4F
m7HvK/MTqLVPG3AyHbugmzLoSemVJ96IMxypzSxkDxCN0Gw/JkNptfnn0xHvTmxb
H9mmH6WVu1ddkuvxioLXoNjjjGdHRdM+TVTl7cASL/AU5XRc9B8tc0w9CJU8JXKk
LVq8QWjm8ANF0MiM1+OpJqohDvgVfbdGt6kswC9bil8pIWTNbv6t8fgvdnA76DGb
rw3hX9FhIb0Lo0a7eCJedo6xxgkfg2rPPqrrXxo9UQGo/lQhLzFS9Rl+JV6BG+xV
7iMJkzRjiHO1gp06ZDJzhFFhxR7hSdZeJxhaNJy5spfAVH/1EWve2ZKiywxPod/i
S9kgiMHrqU0NTBxRgkGgQ+ayReCYhT9hQxc5MoLxNq73S9YGqQOdZ/vfB3CSjSQj
xTsRxZRzWSZxWHEnUO5bvean2Ii1oPgCL+GG4lp086WL8iQ6uZI3Ln1vwqkv4bLc
mzawAw44M6DA8tv3fVQF65Yls623YzIXTG0ojY8fjnbBlZfGd5Z6kSdstc0AGfpl
pmona5EA1DR3C4Ieldb2MEtDOi/vgk7YGtf5SGrTLcPptOaFfW2HsY5hG4n31q9+
iW/wMvdQwBxmmF05ja2lNDNFayGufv3CIjp6/f5VR1/9lCgWVmh3GV29xVIt9unK
dqS1ByRcb0KOIPC+R9JUs6JNEhQm4TRBL0g2UVRiX6EhK2+5qXUvMn61aUFWsGjB
QGVSo9XwdX4f3xUoVfeEJpbHYwnQ51KK3w4n2C9rJ5y/twaQs45KJIvxCCUdL3Fe
WFkszscwQ5ov7DIEXZZhdWoa6DnFQ4RJh8SRX8iOBdf+o21qK7+Vv6RhXLL++Xwe
WIA8tvNEM0SWSkTcahu5mSuK4e4S5k8z58AHxBjSZw6oHhJhsh5xHiDrOEGiBGMB
wH1DH8+WBXd4dWJW0ovJDhlzbZZobXUwopX30d7B5ueSp3q/QiEwHbvFzyI24blq
JVZKDH20rUK/l7GYjC3P/ajAeRympSatFmfkz+n5242yUhU4e60PoAiLn6EhydZh
RzzAcCYjc6sdQeffu1iLZ4eqeVM9igD3OO4wOvZbLJYiDdzTmYzpb/ByGqYHu2VA
i4ezVMklg3fcrqENQYnrDUl6iI8A9TFz4/4aRyCe+ISnJDxx1rJhbqoODw5T4mAl
iqw8cvdEZdZr+2DK0I8fAvpoajBzc8NykqN+q0YwJ+IAne5Oe+gnQvqsWvEbGi04
2KFzpHqe+7lpZIDkvsLgY3Ufl4dXcdeHHRcQCVzCgugn6ONvahzUHlPzgpw4hhqb
cd8RBq/YJTLgUF4gBNka3gVVCjryICScxArJmyFvpCehLs5fmDhYUKpXAHCVHUjA
KltcyHmUEsjPFyaffsVLoVvJbHKgycIpY0JqPnJDYyaPhICBBtTTsRYRp6Xqjavu
12wYbuKi6ZZQPZMcSeO4+UalHWpJ1qzMYS3XqdMdtLgTcUG+R2x7jixIqxdOw8aI
IP+/edVpXydWrOViAoK35LYTW5IJO9BDiEI2XaZ5Vpig+kztoRT50LC53tjrJWFl
l73m2t+uMMggE7yWEA13BnI73kZ3svpsYGXGzFrPBs0=
`protect END_PROTECTED
