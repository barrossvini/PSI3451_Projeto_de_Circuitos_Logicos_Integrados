`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2TAH1TlhXAvECmOXT7AAdsn3aUVy5B0ga8d2HTh1AfKn1aAF/BanS/6NLVqX797a
gSSghmmU4JX8Qjb3v1bNBNdNFoCwOh1GENiLCSN9B3Pi2qmDdLFCHwRv1MVi2AzM
oDQKhlQarxOr37O5ah/ckBcXFDoXy0qdij7FvzKj2imfFTi+nR1gR0srjhyzrYia
DnbR7URjcrJXSc8PilBrKuiPZ/LEKSV/nfPf+iZ1jTIyHv1EYzpLIiaC0Fzbhrnr
/oECqE+drMUjttU+wu4K17ezFxZRdqSZoF9Ye4m8pNJa1zMWA5QLZdrk6umuphe2
i2148heA9JPJ4yTotzl6hzGfw9DIQDd2VdXvb3RWUpYgHSU80G6NqytrVGvuFfJO
+RtBqoHFhrpOOcCYHjMUbYW4fv8UeTsWnFVlQ9QhVQ89uIwElSBVluj+WC+di8dr
agnp6CSE1dF+aCIxRigpWGLX4Kydje1czVpKM0J9IrzWMousGppx4oXBFrhiIH9e
C9Wq6UP6reeGsMy0lT530Z39A+MQ5AvOtvf0EzgXpgnonbwiVDYLccyOVxNQ8/gW
QI2lDsRExSvAWFiILsuM3rKYoyKviuL662dO58pmyqfAPKJHhSVKAquXhvD7P6RE
3pLOokuWBC9fvzRrIQGTwkzSoxqnskfYOvpQ8tVrS2vg5Las1SUzp2UuUKCChdzU
vs77Klvb1/2auieeqEowm8goZmHovsf004+Lb7oIKpm2T6yZQYmmZNZMOJQUiBzD
rs26aEmRmoy59DnJzPKBcv+J4wokimOKHwl4o5hlMXw1FRwnaOmsdxq1LigJZ+j4
dm0g6OAFiWSep1EomgE92Gpa80GkUC3hhdMwzQR7i1ev0bKqkilbbXM1CNGW5uW/
0XxwrU30P359NsFqNpAD0/aDopkt11BRHAbFgRTpBT1K+B9ZQMwNASb2v7RWSYjN
zU3Irv/97EdVmuH3BLL6yMqYUEMKuO20CpMm00WC6NKCZU50Mf1qnERe1eu3UdC8
5Ym9oG+LCEe6y8Qou6MAfb/RiwtFL2zqR9/z1lkR6CBte3kxt5HtJvA9MfP1CEra
FsjYT75+GdcVjzOZdwj4Tqm8JtJ/j+RUCcUAjKQ1NhXOHIuII190F8cn/fhd9/Mo
JmCBN8ReRYsh2YRkV9ijU5lnoCHUNwHzTwjzJgFSkYp7U2fjsp+UC1JqTsCVknCK
t5sWnBV4E6V0ZLjLxrL5DGUg0muJRhgcgB2/cfgQLfo94ecuzJojdEizQFypciiC
`protect END_PROTECTED
