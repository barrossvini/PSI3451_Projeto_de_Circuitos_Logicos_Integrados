`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oGTVdKBfpcyRF7A9ckNKMJyTaN4BxvbIII2j6fCaAaQ4fkcpYViGY0XvYhNOIIUh
DMHW8GyhqRIbLIAjayDDEoroBNo1CprcJtdIgsBvY1tDNsW1wOCtMU17banYspAJ
cgGX/P5NB8vy420QJXPH6PQDD/c34KLIT2EI1aNC4R6ZU4Z2ohXhYmAJKJ6qGDVJ
L89kLBx7n/bHOBOsk1ahdDYm8QDvvkz07eYdLgq16PMAonZoNdpkAKqpcN8J3ZUM
10zlisa6uajX47kKXgb5yGHj+DahDpi9g4AqDP41uz7QmmHdFLnBBCUVWCrEboNS
hSrExZbvhkus7KshvSC8pYKIR8ZvpldHaGy4c0J+Z/tHuZwAUyMth9ELf6jl/3qA
LRMi3kLMcU7VrsnbAK2YKsqK3Tpjoge9eWjqdHGQEh9SOWXbSrnNE1t7FYYD5ipC
C4N7RQ/NJHEryn+hf7JQTuK4uQGqE4lGE21UJh0zolqF/+JgLXAKsK/2YLG/c6tG
u1G3ha5vm02lUFWBcffwTDokDmJlsgjMI9yqbcDQj2XQeQSvL4oLr2ZYjEkrNhJd
vvycoSqNFsu+urjadMvxz4qjtgKi6CTK96DgoM2Z04AGYf7v8ijUXG+I7KMg2LOp
D3bpzjbKpj6kh6EoMfqN1+2eD2LIjR31b/igldZWHOSGO0lmsXY3SBTWCZSwe4Cr
3IGGARTJuHj/dZHHUlx9fWcRMvJeTfU0cNFO1J1qlIwbAxU25w8LFs+rA3QEuPb0
eavlC1Hiw4/AC1pAwY7/7um0WsuYpbue2jJeuu7WVg0EiutnWEiEpRO1Rw7X9LXb
8qqAME6Jvz1LfMxqElYAQYxHUcDLB8OyZoszQ9z+CodPBdKpfanmoi1G96NLuz8x
`protect END_PROTECTED
