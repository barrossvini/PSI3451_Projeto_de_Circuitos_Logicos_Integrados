`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oloOUNed/n8f8TViu6RJXxK0W4OwcPfsb84GUlQzPeIJsM6+xKT9Lty2yB96sKVM
8X5AOALf9qz41hyS9N06jYhumUkiIvw/WBVrm+vBiZ7Cnr4mhef6hykMiUEsRPsx
vhgj+0m9tHprtdeGaUEiuyjNp6eAkHB1q7IqHUNo39m9TVDB0JrS9bwkQ8HEDpf/
glJVV6rvnAIJByP8D3OQLviqx5EHLmy5HMAwHXiMAOicjSGB1vsd0X4EqgQi1rNs
WAQbqsQnUlDmgipFXmqqTRtE69b9mOPBsuIV3WP2p6tL0m1f3/ePQyTAhTGnD3cI
nOfpY5mkzPCDKfsZRkI86TnVWWTy8lGFpLmyxiKTflp0+tyPTBupeplhS/2kjd2P
sZWuhj2l5lMwmXlo9u2Rq0PwT2BPEqMOtTA9mOHuL+QnWpz96DWnXRqF+vVzwEkd
zoRRfy2k6KCVrRMf7Rid81umdzM8pfkwg30MsWPZjGfhJtpBYDlonBtDHC0tDnlt
l3Vj9h0GikXdClME0W+/ReftHb5E4UCFodYKZIanGN/Alj0HLw4LslgLLASV00v3
9UHZVNPcsPcLavr1Okjoj1UwH7gr1k0hg65che6DZVQRTWrXETr0KdkmMfYJ7uPE
t23NRF/mi5YgC2xHlM/1yiTWZIXxhUzzmkvKT5Lp9eNdnSMNCrPfeF3F86hZ0FeU
IVn0VmA6X7fTXW67z6GvgTLBBN5QFcpyw6cxKgtB2Z5Y0nkSIzQj18ilzF7WQdYf
zLP3kQ+l92XqYSm8Jd1G1aM9z+lj7rk3fn9jsaVppYbb6sU2b+eqCFrRafEF5LGs
Fw6zXPSdUgzVucVS5s7tnz2AqU+sVHAAq3KIHs/lv9mJVcjnCqJYW0ILfd4lWS1P
HHpq81q9GDy2sb0p2LoAM0b/qszOSvgfKDsGgo1ztBww7AR28OCJE1W1hooDH50w
/IuLGR1BeacGwbmRhnupLGVAI15CWBBppQn93eLjKcvaCuB1Ap1ICVb2p8EYTyso
XU6lb7i7GXwRJBrPXS1Qtw3D/OUyjweRwkAgRIOF4P6c9CG3WH8s2jIbe6JG9C/W
f49vKWy9GmnjHswpRxPicZJj6QeNf4G9Is0hBd8/Tqt7h4+PABCLXvzabbJX8fQ9
a/tlhTQ4jxusf6uf3evNG2IcRAbX1grUJ7M7tDtKsoaNm/It09a+jhx+mgsq6hNI
nMDmxavm4hgcVhMiTe9bNrnXp10Q2acUTWNXDWOIokV7W7u9BG3cHcggVkLEJ8Gh
+EU91SZPfjTywvm9Od283s8JNslNhtRyNwb7L6i+D0IqjeAjUoBldf2rfL8U08Vi
EOs70btCcAPJLf16hg+QqQ6wPzKfGG+gNvCSDsgsgz8YfE7Vng0fRA3sylwJMc+D
sIp0S2N1ax84OETJJfnsZn8O8K/u9S5UQwErDY26EMh6nGZ02lp/rQlPYW2JgXg3
RqV+An45rLV5A5SipC85zu1ZRUy2Y9ifj9IvzOdUwm7WxhlHqbvlU7WYqyZyz6Mm
ujw986wLRfjQtXQqkRBqXHWnD/Z/31OwGxh2vpiR6Pq7W3ZS8CBuAznfyuuk6vBw
dD+NSKDRjZkOY4SXw3uvDhJUzdOnlop/wY+12fu3Z3OSVcGyqGUD4HZMbq4LaZsz
a8pKfTXghkTTLKFZu4Ua12BvhRnQBzmIED9uA/MLLFU47poqmwzK4YYP5gcFN9O+
WesgX3s+vNchNmf39iHSzZSEldOXG0BH20Jjb6DiqvbXaVEOJb3n5Fm/NaCh5o/Q
JslYBaZ7MtLw64uw34ZugpK+mQyHYvucBPspHF5uL4mpidJwktS/jberX3RK1q4U
Y3HSUeiKTEbdOGNeU+L1aokNCRjW6fsP3sslypt0jmCTxIkOKuTB2h3r+c4eLGN2
BLZoAFFXCGdQSP8fRJDctbr1OqLUvhfUE91LHDmYYwvNjmEAh7UUP8QBJSri0Ybe
yZ595/qeOWjvQDtEB/onhdhACPQOZn9ugAc/PprRglrc+x8qESjDaJG2ZcFZVWO+
2whs4HQZzju4ndwDy6zvagcDQmpvBxGQsJ9LZwBMGXBuTX+k+oV8fgMYIx+W5Kcp
q3s4wCjrQpo/L/2AOEa34uEmwOs2mnlNFNvQ4k4Hmrh86ygGKvUyQCyS14eYZRa6
xPlvqYe/vY9lg29POBm13+ozSuxybegW0tjumqYeezoRbnxHEXerfCJyotsy7A+F
/M4jAnqmTB4/L9N+Sz4yKAU/NOQ9ZTEBWDhR5kcW4YRAgrS/Qbb3SyAwCT6NYrEn
yfH2blmupgghVyX3AYC3aYEz6gT7Py8pt1K6dzXS2eAi+CaUV+UG/JyWod/XDN6G
U10eqgMe+RVJA2uQYaMKp2WcY7S+3O1RnjPs4ne7WyBJknY/pDmZQcVktMXLPE4e
+nPDUdyXSPtZUNYb897sIl01l3Pe8gicNJ19UgKFcMkKZUpbOVQged1+i8U9Ygoz
2PqUV4SK6TKL9swe8Ku0RuvQsgWBsYi3zct00FfFHbEWsUjFrbzxC/V7xBbA/V2L
4R2JdEIbAP9S6pD6/J5fICFLRR82Ic5w/RikbiVxdNjyVyuo8lWBLs6Dp0TqN5JR
ITRjF3hGF6tDpSpMCZbwGe6JEjvlJeYWniUXlPDc9W9YCxJq4q5Ybahvv1fMjnwn
91fDN4C32L3HZlB+uai3Wbn3LAPhKAVIWxhnLZOB6P8Pi3Kergs3EV0YyfzkXkgR
Y9Pw5ly2JB3t+BwyXRoCPLe4kKu/qznEKb3x7snIyHXlQBGFd2M7a2zWg2LiplkW
jbC6aWwGeQXaGAHf89MKQGMiuBAmRk/C7BIV0xqZAApYMnCW0jS/xRbZSMGO7zr9
lVrDGuTtIk65CeWetkrXHI2hzkq+Ok3UgLduwb3PJwBYyE7lPHUEPSEQRucaWDHT
FBiomz0ExkldBRIg8YBWpjAWgkEtOaeAq3DHAGC8BagdIh5Mr7jm4XZE8Ma8rIEJ
06jcr3jU1NlLvIHbiIvLzHkqWksC0ZcXpiuu4UtUPIJL+BP/zQz/zLX3qXGm4cXq
+UYM45PHejUB+kFFy/vpqc5nDHUTDW60MIN56k0B1hn/2vvNkKkxb4Vk5tix1+iE
+iUuXo/HbTyboJmWFMpBNYqNY8N/GHvd3h34VkjbRarSVDowUPZ/YlwDnGfFBA9t
aYgKc79I4T4g7A6NZ01cdcP7FNo5fX3c7NQ4sTs1kMgLFwYiaqzV//ZzXf77SwF2
a6Ee+0MBrQpwM1i9tbfngeZURTVUGSxHcFBL/72V/CD+TCFk5CgZa1k63KmhlY59
cV0ouDLI7TI190i0Hr63fEYDZb3/bidaYAG26HbzB2UtU/x/c717e1J02wdD1eTS
FlAhn06SVsgT1Mtyr4h8j02LPsXcRF1ttll/UVnSlmD2+ZctovPind0atgETA+P0
+31D8+49Qf/iZ1hmmYp+7W38K6ajKAqp2iXQdSWmj9HeaVBobf+WpTX0XAGbahwV
lrcBnYCxM3HLVVANpmOsm7EMTKNRL9mulJvzeo/NOncZhmwr/IQ74uIkU4wecOGH
Kl3k0ydgquPxl53OsKRkXbfOAzLaKMVKx7nVz/bf4KmRwY7u7USyX/yA4ClD2Ihj
qjff6H/4a1BVAohVxDXnTH3aQjM96QgRxUQxnN74avw90k0QNSCQ454DvmY7HOjU
g5myqw2osjh6LPsqyNM9teDScsNHMCKBpjrceO8/5BNLThqOtCYimh2UNIQZcySz
ZJaOsMgacubO09q+8V1jW3XiWBEGAZZjD9cokneLv6A8jLPbJyIyYmxBqMt0BVLY
+LMYYpAaq9lid8ZjvgGpi7YrE3Hn2IKqAOimwNivphRTbq4fCgi25A+Orahls9+G
2/aHaIAxQeOgI4yh6FUDPq21DUc+1Ldq3LlvHYPtQlhty61kAjeKTd1bQSXFOLez
TY9nvOu4fM4z9zyjd0FNMlN8cpXSCyQ97s/+zWAyEAgo0ooZt8PL2Jxp8934hbdR
1fWePR3ySgGVh1NVc8lPWb9QHe9PIAZ72tLbYw3JCR4a8wzUKQHR6XJ6clhaPwhu
PVXr8Vt0w+sBhQsWptKeX9wxRGJH/s2zi0Oh7OpwzCeIhPUBJclXoR0MiqExHiI8
o+H0QIA/jWQLu4BhypOhzvSjxuEMDTkcBCnAnbmoyZknxwRz3TyQxPmIyLMVsuz+
i8MDo4qXQlKly6P5z04MuvFwh+vNwWOIiF1Kq2q3+GrxkkU9y1j1V0gTcpFwMPEz
k8faq9MEEexPw0NzwpCAMF7MR17sGnWq3PF8D21Nm/Ay2SJ5vkabUkTmhD252d0h
A+js40qIxQbwIA8vBe+7EiIBanjyOeGCmlbwLau3c66JhvmtKuaC9WJi2hE2UKuk
XKg1QGVW08GPiTT/aMc0eJAq3xRKpNiorDWZ6/R26hCdQZ0TsAZ5GKpClAYVrASm
oiM31dEKUkEJAFSjUJwM4xR6O6J05rueDGHIJvFpVu0K/X4qST6QhiB+Nf2D5PF5
PeN92rqyf7hnDGjUnJJM/kYatysUplPJIGc4rJL3OnV+bM4lbgamYcAiadHYrmXe
6rsge2aOd8Ua2FA++uf7hogjbYWcFFLvz565W1tGEiFRNjpi6KqzG9GqPeBauR6h
TIyW6M6lua7tE6SGeUmdYIxZ0jPgnLTxKNdU414e2WCK1vti0b/I2Yy+dpGsQnqN
3wXRlprOfcjzLKPclAbYFzuq0S0kRXwDBMK4QfTke4tnj2Dd2uwGLQyZTU/4ClEp
/zMEFEkrA+hd/y0naxeMJXRLgF2njCJN1B5WnibltqDqEzV6z/vyiHhhv+9tKM2J
bzQc9bJiE9GNzT0G7jY/rNSJZrAeY/jnKoieWszWLy1LsXDVuYJk5wxDHTQVlrYQ
IOPDr5oM4AVcuqJasJBVrJev+kjuR5KHxXHNlk7ns7cdUZzZRmhg9lbKeE0eUGad
DbEIjKmsew7GSgAgLlARdVPATfChRHkhQJzmPy1j89HTg/raahVPoYH3DaISIhdH
5FD5VMM66msdMhv7wTvbmM1n9ilTehTGBRtfFAQal+l41pwyDHwRD6hq9CuWoEHn
ACG16vbisqtSFzYyW0Fjx0K7gJScRr8XXFC1Gp6nXo6g+OWpv5CXEJ872IWd5bdl
utys8BFvxPhLPmUJOHLZ0kCvMXb/OQVbxmSGQYUwrDA8GrUy2GW0xciVP1hSyPiy
z4WEE0KTp4jTE7Hn4Xk1M1IAv0ObQV12UJzqssTTGT2PgxMUn3/0Fq7X2B60xvie
eSIFzgAM1oVOl6GCu3nqXnsvNYnO8+bybwCkpWzYfctf+aqU+1rsD+xAVZymK09S
vTGI+ZkGhoI98eEinhu1RNAVF2IdT78VEM1Mpsojx34XNi/6soFJLKSr4jFdxxp3
XVjSjpsXOfWVsLTV7gG7teo2IeJFWjw5YX9ZYkNB6gdwxIgaaC3Vh1I+j6S0FUWe
75klPmDgtE4TGZE2ZbXDb88gWXrI2qLkA/5d1H85wQJY0Q787KIJl4fVi+qGFctH
a/RuAAPPy63EkGeWr90XP+4zH4caCtJ71apBTBLaXNuoxWL+L4wcdTg4r6mNPbgc
uoi6sQTyaJY2abMH7Vq8VYeCyEwRIXPGPrfRYXVG9nIHvvl24NAjXOKfaGC3Qe/t
YPEaUOJByJvaHBDv+oZiabWpuGNNFgES4gNx8JsfXHssb+xJRf2FVmosbj0qhPPU
ztqiSr5sbmTzc2E/fzg1n4nACBMHOwhUMwvkZWg2fp5s3306ndkd8VGXhI2GwpRR
1eBhJbYU/dCw1W5YA9a9uxizD/oz1niuBAua1Aohl043z+iFUtc5sI2Zo6mnZQm3
9HDnAnquesiX8/JpyFv8bZOoQ4neGTw9sbSuT7wD39iKOHK4BfriLUt60Ggn/1Li
xPbuVQi1GR58ZPOf6K7HNBw6A2SGh6P9XxVEFv7GcQtWNqvhHMCi+OcGdk9Q0ojb
kPtLnro+evX90YYKcJkawltr6jsM1P4GHHxiSO1Xb+IrkN9nz4VJJfOGrAx3dLgQ
MSSOO1A0FjzHrjiLdS4GwbG5SUP6nLCY1VCwqs2J00hCuzqAq3PUirVxZUdBst3o
L8gC/sdZRT/VWG/2dnWsfgoz48gMzah2X+Yi3i6SfMnyLZ2oDrwXfXbNkJeWf679
a84HT+IS9otN5pHb+9NE87G7J/17nHeW4crGcC4a+88l9L7x7ledsb5uPx+Dlvuw
jW0BVMCjyyVGFcSxjmuVb5FV2MqMpulDS4DAix/fy4yPOxxtf2r7YZQJdapkR+KJ
6bt4tN6Kxbk2H+y9BEg58KDnTOLnEgr5jJlBj7nbwPtzPHuaswwri+15cInEerT/
RLPrQSOJNLd5MIpfhRjEhV26NZcA+OFD5ks6F37ddSnBdhKwYf3lpFm8RwuO+DQE
IoLzkOi3gjdGyg0KBF7Uk+l70OC2alCKTSHrN836y8UAAXPB+y/7VhhB9eQoBK4/
ZUI8CSSF2C2SbVoiZpZNrpTPpZgpPtBUoAW4QIs5wvuIrNH8shDcyKM0KZp+2rMC
Lw7ghwI7qGuWtzTU+6YeJSnpAKqmwKj4J0+oXPkE3Yv9lfN/9tuoCPHp5OSKX6wM
OGvP3pwawbUstKQnELAPqQqZTtsylJ1lufIS7QjQg497oEH8/oLNgqea4jpD7tqd
V+SzQEHB+7LjoedZaM7j2EXpCL1Nf9PkUWbFBzQZbaqye470Sg0sBsnRLLqvs1+2
EwNr/c8uOlVD5OMCVMvZajuWrtpyLyS4UJVSNS/mvEdGd1r2rdfsPxH9POn4GeO0
Tw3NezHcClv/WwgrDlB5a7J/u22k+F8lAj20bCLtsOClbV2cEFn866pLzJKQiP1v
iXju2v2nuHyOfNxVa23riNBC1cFMuxAo/Owh3te5dO4c0J0vAemHfCsGu9id4muZ
7GAqoNzwouxWtgfn5XXZrPAHQCzBKTNqVLcSPqLHL37aSdVczBtpUTZ+gblGtwpV
2lE3yMHUiptHvXw0AVgC1ASDChYgCJVxIi+PeoSimvYPa/b76sZ4wDJFmRtkh6cF
rzMBqA7hYCOa0TW3yBbidIJph0VwEn6H1n8MP8PEiDsgNmSvwY111DO+vJMSjb9Y
TEGaPLrFPNzqXoGZEELfZXUEnwBKfAsGmg+bf5ftpszKH9AmSFbfLqFHD7+Mb/2r
VHMb+Tw9a8nK5jmusvjTko7nV0itq43BByfWgLm97A9csDrPO0gksoPhSs5Heid6
+u2/B2jGic3I2vojS9SZRbYVP7EZmYM6yXTv5GijfsSxFlygJpfujbrLMiLCJALD
v011cufIo2Da/ZujWUOCXRkHrYjmvQV1u/HR/dLpL+pmcVBQuQowda+r9OmShllf
TP3LA8f2Xk2TAG+M/UfaVav/sBfTx6v0lbDIuU1da/mKoTgX8HGp1iDD1bC25Q13
nHZdCL4vJaLVByQIkgeqjCScXydDGIPu8iCwdVR7zazYWLGFa3NV9JsdsbNmEZ/9
qS6z0Z5zTGOtzFvzoZkq13gUGBSAjaj/rhoeJ6uqyC7zyWiV2rj4Uk2/k0nEAKTK
X/bqyGN0ujvQgSs1fkA53/ID+qYbdgFDDMuu4c3y4BG1iJhcX7u6/z7GafeVKFX5
jrDSqkHUpDWeSNGBhSJVPzpncDT+t9+Feb246N2Q9QKT/fm52d2yLFQDWN0V8o8X
7yy28t9bCNCoiEKmnFlaLK/Cwc/EjlwpQbCZfKW5LR5xnoRCLuIeTt8spEqNt9kO
Q42vEptC1sW+WJINxpE1OeWSFuxB6yBwsvSbRRtzKYbKe4UnPgUlR1awYzd6bI/5
Ap9JxarwrEvyd/JX2Q4or/0m5Xfn347ul7pv/kM56SpmaVpEnOzDkTTAf1nLTJ+r
NcWCGJXYKPjEqmcAIurdHrI1nJbfSyAslyCKSbf4fgCpA+mnubGDWCKwTE54BaCh
9X2OvokZpseJ/t9SJ2qZYBlcl6A9B0JRj7NuVHm7ie48i6A9OOuxJPFlXuSsPxnj
hyOMK5eigu8wJyWTmpCq/2Anu1xTrLfNnkjVXB4E9S0ZPNLgm31Ook71L+gcAjwY
Mga+SG86aGL92QuaPqocrfKEAq/nODkJBOdQ/E2rx23tKra+IJYkJODFXjx6q52z
gvcOahQnTKzUBV8YVp8LG+L2ectAxHZVVaEyWzOZ/AUskWKYPwzibr4D+gTyFoPc
TeMRMkxKg5ryyCiWqwfVyK8MRRrrg4GDmuWDOhlZPHxVfk+2hfjwugIvQsKQO/Pd
BaX/bJOVmzHGKjKyTg7rMOfh2EeUVPM1Cvetf5kzSdZVfZSMM/XU5pyupD+1L+/a
ZdB9/EhxgkhY1kARlOWfgf5gsivystEmyLXTrHpXG6iGirsacFN65HSbB2qEM9Yx
p6DYFHJEb7tMimbIRiabgKzBqUV1ws8HNrDg8c1IcoOoJWWGqx00DjFUfvD1/vpl
Zlvnxw9qjY2DQwuVXrd4o+KdouQ/qoiHBm1ohMbMv0t0g4pcbYQvH860axJ5O8dP
UuFUKgAb8+JQUJt66H9TeBjcaBQSHEIGo9wr9q15LafH6rBgEmtOHV1qPPf7cDfr
9AYoIRHxKQyIbLtmkCmTwgldL5kMI4s8p33mVzui3psPsgG/50Ghi8cav7JS0GrH
VjENPwbF93Pa/9dIWkj4HBb+Kl0tv46t64iDfwZqaOpmPcgfczJX993ecBNucNpW
D+sYe674a+ReoBNqD79HOwB7hwHV3O17IQsQRaI5CyOBT2vQ30F9trk/K9etTcoV
JrIA707AU7fUO1vIsAMkaWgthV3aofN+/fZ7BlsKCtRSwHwi01O7jqYjb4JzdggO
CEmUNptfNGou3eOZD2ma7w/IrCDHizMHqmKTG7+//WoaXILEJmMj8ZNfP8zeTgqE
var6PuQlrq9gQpbAAwRrA9+RQAnSaHBpGS6vKVWn04gAnxyxxRu2ekwFR7H4/jkC
ol6f9vACaePdYNMFAn+Kcd2GWkmX9KkIEpsDcNFAvtm7fT7At5moqK8TPVrtLPid
8w8ouPllUvM7UAb53yqyD856aWwGcP69+tdOV0fVg3lLovfPUpEiA7Qzb1tKJ+5t
SFhdiaNodG3opgs6s+I/0dADNUsqxL9KikLxiBBpuqNdA20fUdRYoF4ML0WC7f4f
RlnUgjZbqTWcPvXPY51MxWRMHSzBFrjMEotWR19/pNyJqrDP0Wbl07K83u48HDqM
YXw4CzPEK9WnNjMmW1fcdEGrWBh3YRnR5r5o//3QHlNuTRJwkLYfd1FW852qJ9e+
1ot6cwAT4t5vVGnT+u1BNwcFo7feL0ylFZU18zL4RoaHIo7SJ/4rSrt+q4OXcbR8
CxWJ+vX2j1/8J9s6YWBlA6BeglJ8cXqGf5OOh952Eol0JKLHCLULXkvMuzK56jE9
bFvuspDr1dyI1eUFUuEbyAjFZs9Fq8bDvw2badixC2JKoCCWNFDByqc5CBqDORpx
anXsI4SGnSBac9znd1h9AzeHkKUiMYB/wdL+V4zjFdiyYUNlJIkWDKd1LuWw7by9
HtgmKCOzl+bNq/hsqtGuSUfsAMIF7SXli7BkXl2asXBPOzlAkRxZQUQFDILFt3qZ
JIueiCVYgv63lw3eUsTZQZIpJCMs3OZVnaHkgmqzRf7kPILpnoJgOUSv8odAnE/d
wF36J7hVLkLicJvs3ctTSwhfA7TH6kLTW5ykcwmT6qLaH3KeDQ4vhncrVGafNJj/
N8VRcFirstvMeRD5wZ2mlkkezo2agxvKMo0MH8NZBaYyDo6i6QWbkcwHwERSACIl
ObM1j1P88q0huixt8MfzagzHDE2gFJjLuymW1g9IGthAftNa0tXVfRnKFii8fCeY
hwMVTx0vvbloMPy0CPRF8gqGVXQMUElrIJsrWbtd1DNcPnVsneJK1e3Gt5weNwp8
XWqnpgsFMUF5FwxSsQscFWZ18YlfWcjmTovdJ7PkgVfEDkKDqVj2CuS39FOPszbU
DvpfUL1vsY2cGXYxAD5RPWBS0IT3TcH7oLnKJv9toLP21WMKlCwkRJ2WJqkZO7Nb
8W/zkvXLsgnizNOQsNt2esQrJFjs4EZxJrQGFFiKQ1ebO8VR7kbBsF/ivgNXAZB6
eZ4v8NfjTD/I/CckHKkPGMAg30ig2Utf3q3pqc5yYd10SEkbbCRIP8hgOecs//gK
rpm424Tf4oGkPXXoDQv2YK1aoIYvl+Pt97D4n6eezt8ehRxh/SAtA0UjySGFyUz3
NnUBRMhh+v2Q9avTXd2G5Ef0S3qdFTNFtLvTFJaz8t1LPTpKNAUNvvfl1JeSx221
OkWaWwmATllVv4sY8QdPG/au+MB9Iu+7Ign31bL7UAukhtS868CCZZIAvrIIPqH1
6lyCDXmS6QJHL4dXcjXEoWbpZKoQjTABSGN73EqjzvQHV3I93tDQfuyHMe4dZ6tN
N6tZAK+KIUtxpqtXDGMcnaL+10ElbRH5m1NBmdMhAjw1B2L1KQiUWUBBfo4bHk3+
ywCQ2sutQVYkBM0hRFbp681z7CofzQ5DMsd6nspIsnc8E4riS1bdk7asHPUYbFBO
OaBIYI9etEVOiX7JT/LjwC0MiVKOvZpNXM8pPCf2tpOuCTIkN3boSsp+XwfY2PV6
vGHAIuLQXmDvyJu37KW3YmAcc7uEKdZnkBjSV62Ox6RgWnHED70yLY7KLqtEarLt
cEptfCcOTNdWEejN1viwlrPaPciSmyfNJy2uIFwd4cnv7PSA6yXFIyv4VGS/CZO/
QjRMQf3K/yg2zYv9a1vNXN0q7QHd9KzQnSYB7JINebd0K7cQsHKLx4eRqaNxBFOO
I25Xa3mQhaoNCfPJn4kdP8mNmX1BDGIWsG4pOU2DgGYVNjgNPk+4oIx2IrKpmvFM
bLCfuwraDhHz2LMFowxjrxaeCwfiq2UT2zQqOMktaian53j0Op2tNR3xmIt0yX8I
9KeOwdfGI5NW5l1f5liPUSxvQJZ66In5kVSt8jukrVfXT14R1hYDn7Mi2GIpBfZN
HNt4bo9NWpF0QSnBFcjBc+9goplXjW4RxBhtVZ3/uhPXSOX6ccq03BzpV3YVNjco
CiYBOeYGxziOTGNDAQCR5pj00ammB3sd8IZ3Ypm2dxjsXR5rvtzwfoQu2PyQRMTC
Z+Xs990Rdw5ViCIOaXaKkpsStY6VO+fK6fHKSL8zWxgtK9eLlKG+IAtZMjvaHDXU
RLTz0caNXlPzOv/2q0DkqmUF5pZFbCbluajHl+krvDYAfrLbzKK8fnqDOOxOn9yK
4i5Q5UYfRZntXxPl+z5M+8NryztpNoaeQZxp74RAC00Hv43MzNOecrh/+o9jWhi1
PB27tc5CO87LVTWzv73qxjNe40mLX1g7/pDtS48JvhGN6b9M5lE/Q7Y3h6RxnLYZ
hQy/3NzdR35ru24a/OqVWTBwo+SrJ64i1wo/PFri9AAYk3H4w3cg9PWKKTX7pWwi
x7xLd1hTc30rnXNbUGHreU0/xGyMcYkxM8sucvJL4FW5/ihnAxo8grfcSHuyDXT3
nXzz4vXLs9ZONS88dA6M5p6oeaqZM+nrzZmoP9Y/EnW6XP6Ae9eT2OO+hR32R/Q2
hBWe4SvQ3p80L7y4eWR517+OMq4GJOs3I4e4zax1VZ4TiEmdbckDePt/4mHVbTpQ
Y4OfA43i5YqMDrF5sdq8ZIlNuzbD62mY6pSzQGxqjX6ZoKhX1CZ4RTWwWaVKJqoL
+Qz8f8SICO3k0D3CmvMa7YWL39jrLKta+yh9WOedcBAaXFXJFi7ZVJjuaz6sDGV3
UWMoMYlXWV+vqNOWKFjs4DZDUBLRd+POf6HwCYyqT1G3eGjQmNfKxeuJOEI6lLU1
zoDLgNo4058kc+lx7pKI3EiLdvNCHLMq1WdUrOlHXjHUSwwJgWjH4SRCvQ7aAgHL
6sgelM0h1PWvTorxzIiBhiS6KJQrMsI2RGJPKN3Xt5V6ZzfgF0Qmpx6Do2Xdfyhh
6nwIlikFVuxfJMzExJoklaOadiUM1I2JH6hOg2ilvm5N8baTc4Q9pQjMMlgx3GH2
PBH1OMaLw+U/I29P+qW6+eTzr+SU5naHqJeMYaF/SJcE0MXoO/FXxDIWpGMRdabU
HDdhitzs7skTyuCTEwcha4kqSYX2TJcRBlQqvLMmFDf0J9voNErDCh38lDmx3pl/
s73IfTpm/dIaF2vskCU/cIonPgbZEYCf58xXJIG7ODlk4JdxRcSznuwYqE9gMylW
K5KWAEV966Yo4cyTfvi+kFtgAdOa9uayeaPBCxnhxy1yOoPLHsnTwTdsMu+DndXb
VxHy9MO80rk39th+QyTQ3V/Rb9sTmPYwnp9MbftxZ+LcoDjvksN4VSWOUgDMiAYj
PjuIlMK0iY0pj7nVH0yJgvOrjdbrsVbYL2GDj/g4jy0i3bIjfq2oOwU8B8baTbd2
snxN+RrkXkXRF2DVx+UEvmukSmaAATcJSlGSdp09lHkxNzvNJGWNeh+JWVM4TqDi
BmLQChT0c3ysM/1ilo/voLMEuraCAtMRVnE7jLITrB9VAVyPJe+MQW5SeaNSxewy
IdgksEPzgL1dG4w5d4SCe6PsQf/kJ/QFswkTZzFV+AH936JZIjtIzbRG+be/lfK5
JyI5LZPKW+SBgALe55kOz7ayxovcISeugYiU62gE8F5ri4PsVvGS/ofuZNym4OJ3
yzIWwos8CpgI2X4UxcQbKyOh2aHMXHctqOXsG2GfOZ0v5gKCFKVCONNLGHBk2P5C
kpFjaXJvMwkwAkZ3TkO2UG6pmuSjOz1rstteKNmczkbOlnExAXeOWOeQfU9qKRKE
+r6JkZmtn+IoCcp0CQ8ym9JfRgBhaPsC1TL/P8W1Rn9mHNJ4rBy725LAJrR2L6VE
F46fVLiaev9LaaJr3F0aFRJ8GpCGg5+eVp6GnpmY8MJj2jskFAnhWOLJYvLKh1lC
MU/bT2d9dGifmef3+VIJYMehvyKWk8eD86kOfwtEr66y0l0zWrlvaCOVCYpya2uP
x+QeAJrje2AV1lBKlLidkPvGfKuV8dFmsT4sZhIfDW1YoBtukNaDn6mfjcH44spU
064tUpvC5VqN6AvcmBjxVcZ3V1JTBFKpxA5JPmi8EMf+wAy1v7DNo91BUk/BKidI
HfubOUlYUcDeVLfxAER4c+wUPI47PopltfNoC7smkdE=
`protect END_PROTECTED
