`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yb1OBvIl5M/dg1k1rU+hDT0ywsiGdEy4nV5PCng/z5SjNO1oY/yIB6/LU2EuRKqP
JJu8B56Eh4OvbbHonuQO9VEJwXD2lC5ZeEl8q7MZs38WGlg4N49DI8whaPubR3ht
s8NImaQKnTmdDZWXHYCQjkTSmwGd7Wh6wzB9NF40A9mkXOlTN9Y9IkwJ2Gk6RwNC
2P6cuJwVLK/DaSNRITzylEE43p98Bz7e0725wOqRJDgXuIli9p1ePcur8c/HkJT3
CJd/VZnZQoENf0JFBMsDbgUGem/TCuxrQjvx2AQ6WGUMaHrTbjtcpBU/W7ADSQGz
hNyTyqWXuyZS78ViNkVcdY9nk8Etox01dZruf2eHZ8hO1EZeDe4ZCJFYKYDPDAfv
1gPJZhIN8iFm1uf8vePhsyu8b0jrwOrPvv0Oh1LNwqlZ2FbIlJe8W+PpKLYXTwAc
Rmiia2vD+GZBoXdfNnN/4Rj239WL9f5vKY95J9uFNIoN8+tbjFKLFgVz3XEnwPE5
0UrID+bF3lAKkpdd+lZUuafopP2uEvUexAA/68eUdkVvNDGlVH9hN2tO+RivdITr
ytUrqoR3NWhKSElCp6Z0V0Ey8Y3hqIBko504FVfOfwsHJVe+lJMpbjV/LbZUUUSa
GEJQzmc8o9Ms/TLT2cfZ54raVu80+P8lT3mXnQ6kZA66NoGKj3cot3HDaKEaYYEX
V6C6MCRmsUBcdNS5Ar5wMU44jCyqvGVTUBwwlbr/iberfwwRVhnXNfgcsuplqjB1
F/Aox3lfNp0lzSj0DhEtnJhySbXA6rvS6ScCz2KjMbd0RdiHcaMMxq/ghN9pV0ZB
NxdhviG7qHohCiMgfU9U00l3KA0lp2dSaDKiB2xvZtgmrt7wMmjSEleNc1mv/x0S
R4HerI1jY+krV4Sl3EcfcpLpwby6IyGcItKP40QYmyiypYf6UqWItY1KDFezLXey
FhfAt3py9BKKpk8JLAr96Nv5ihny9kQkCtp8r+sab/flMqFljuhtOBqYK6SeRTFL
ITNF/zqGnX4ZAyQlkjVzU6TgX9dKIxR9J43hq8q4s3CjfhTIMB6bG+0V0wxZg8G9
ug+7B9b8bXv3i/BzakSt7Se4/KHmJ14IUhs7/sYa3ZX5MY4jIRJ8FxT3kT57RKMs
9EQr4Tn1sWWbZALTlfTk4V3n1KagAew0CZresgN3y0mos8YMOJCVCSor3RMXojyh
yUE+rsyxpFMYfJQKaRkWU4t+soPQzZ41BzXxPvTk2FxNIeplji6h5596dRI84XGR
OG6XxVjVAd7CdXBQA13Cw3VRyOxD0HCLd5kn3SmjuELhIQ4+z9PwkVMp69oi6+YP
f6w9W2m5076WSqy6AzjNQCBzC6dgI+6KQv5G31Y0UyYqMbvqZTJ55vkf+jXE9oLn
Hg3kjkiUiUj8eZWcz+xtpwfUk1KimndYLGxIUAXs1xBIwadwi8NiOgdzZ8Iw+Fw4
DKcysWLDRsOTeZO+o2/4kS2zMN0A/00OIanuZUqikHUw/2RCGCgumfytSkc4NcH5
LsDrFrS9kb+qehx3XWVeBorBH8cC/63oZxZojgOoNkPVAJgiV943M25J8OStsL0z
2uAXyhQeGBYMK+bi7V8RWWRGxGtUUSZ80EFRothbNeki7yUfM0sCbhK8Mrldeexy
ArXyIWsNhxkY9IPF7bbbRubzdIyQz1dOGSRRko1aH/T0ijMa83K/dMBH1bqHGJWn
02RAvSNXSt1IADDd2frApe0vko8ZXmaEkkwNtMTKVrYzzcKQQIZ0rnbC2j3tW0H5
lXXd2GiZznnUZMClNgyPp2YfEoJH3nJqAip0gujI8H7d8iTkzaqt+s0Cx32SestA
1/A/iTBGVIVxtxmN2m03vumZRvYGXelkARImzXH+xeVOr/E+U9T7Q5AyzXkq4rcN
octB6eg8AgvtRU9Bsz8jeNqQypl2OR2A4JFx6nQeh+DIo0WxUQIqCFgBa0lkWiSL
ntgoAnBBVlKk48/fNOfj0SgpoJ4fIeZACfHJ7mZcQWiAwAzPgdam0HAff6N8r0G9
fEwYJLk2xFlUv3vH7qffaI6dTuJ3j7ZgfuNKCPAlAWBRi9vrGBwKQp7KoPhaELwU
l1gmzqmaYrbRWf8KY+h4CYRrlunNE0+EhZIh4QrHFS4kgjnqPWjBjXR26tXuOOJW
vsrwFbM1lfU3FOjFomMZzOJi03mwQSzHGbBkGOnb58Tw3slPkcrhDuC/6UxtEiZj
wwMoPlmYz/D0yj1geLwScaxL++aMgS1ipBwmAKpM/4KbyipqJMqfKfO3h3Ifvgxj
vvAzoh/Y5F4cPDDCGLPBlrbrgh0nOmfMbHYhFNX4lbFmgNCY4GFxFb4QqzkUvIpl
`protect END_PROTECTED
