`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GyqogqLnPsgkTpvpfxrYLsij9LEr5mi+/M7mPET71Jds63rR7L5COFvqkMJSNzxQ
kNWoQBmvlK5XnibrzTVmnttFmKzALpEwhA06/MwaR75BToJlGF97ExFAxIlLyOvO
HQbEHHN/YIlAnHRxb/YEKssdc03G0HPtNt3bP3MUxnh/0u9oOO1ptLIZ6PsVpcok
qqudbzRSdky6rqQ3kolMDdBH7K8cRE/KUlv9XXbMtTaL6KxFslUjGiSl6Be90mJ4
7zNG+h1qK2/WsgXuAUy/0xInmzJuYwDAbMH0HR/gMcdeTtOyXTPgfBO+mapvx7d7
qP1pZDmNswq8FKkdxyWG8x4TFxu/jtYNaNskMeY75PDBzv43ZYO8iqegnIx4Oxrq
Ht6WX7qR9ZqhhJNxMgTAf87FLFpD92n+3FPiH2iuRtjvVKY2HDro71XJ7EE6LjGF
Qg3J7JwNGgBh0ByKZUMeDSLqyYmDiDbrTnM7rXdRQUsCQcRMKROXozNufNOWrfVa
NCPftU09DnT7gLdry22cJXZskzN1Bl/3vgitrbCGTWEfIyUnNozWwCjDp3YF3BWo
0jSa2Z5ApKBL0gIgfxmnayZcCf6X/5umyRtBgvDqSYsvZzbbEL4wECABeK/1zPIj
K7rSK2lyaJ3b1kOPw/vAhTayxIO/I3NncH+BgNICAkiYMtUFAIjONP2xbZzNoKZJ
mIw1VSfHYZ5cHb9+EnE10v5c4v1vuGmSRv6D3seq39wvk2lrdoG4U+mDbJ8wmQ21
vp3RHt8mgjAF5tgkjw8nRs7yGqweSkwcekI4LjCHZ8o+f8zUx/a9SV1Zo4yoLyeu
VDpOcldc1yDmyYbT7Eq1l6yYtOCTu6Eg8F1dHPAjm+us8Kn9i69kH85T7P5cbVv+
BesdwdO57gDwGru3Hf1Xdvf/X5u/3hl7NX8s8Xm18dP84i+JtAzVfSD7T/sfYGTt
iNGiFV/Ztpt8NB2TaaENnMEGTbbByhnboN31AF4mzTf+OO8K10VpHOCeMeGewNLd
TbWT1Apwd7BHBEDok0YetX1QwyqIDqaeiB2DzeX4M0eY90mYdEn3zR3lfsMfQIDO
tsVCErwA9wIERuPRNIsEeUXse5UNYx6mws/cHqigXmM4Ky/6PGwXKBT4odHaZZ/5
OppCyQYmHiXiN7nk2qBFhkLJ94HcPE6c5jAb/svg2tg/iEk96WObyMc17+pfe6vZ
4wv6QyMmesPQQM9abTckVLW1KtsBQTKwiJuRs4/J+9sOQc/2aGZvo+5bS6LEjAVJ
+EIgjK5ROEMPwCeTRwt2BkbUh+eJ7jOgcP1ZLgjNWqhpez8XWOzvyQxzM5082Z/i
aKyJ6O9c/tbKUZA5xZCZ6xyXckUOGehQpbwVLwHuR8fI4f0mQCnKqQErLY6GuCen
eIXzOpDkxuDcYN7vWTd0eJfj2Hwo6heFxR9srT2knFrqkNL450b2Vr5CHOQ007l4
8lf7H9faTyVY/M5ivF+YcXgLa+dqW1sDn5xoaZHkbDQW80pM2tzUpPepp0xpA8xV
OuiSEYGp01Y3fjCYQio5Vw==
`protect END_PROTECTED
