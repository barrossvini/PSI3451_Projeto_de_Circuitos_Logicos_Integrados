`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XX6+AKDuA/gAzkvqsty1StVnIFudJBdBwL5GLwZX9Onr4uzyS9vaROaAGOChjCVb
NVeZBifV453f4NkVGsH7WGGJJGtU12x5ZsdhM6HUa2wyd7InboON5izJ88eMesMj
r53HvaO93MSkXikg6ATrJR314sXXIzfOxPzWGPFLe3KX9CTM0YuZwtVMgxUdbupd
L2FmhO2XvCT5gAgadaDNQb8aO65y2xqr6XQEcwyBXqhBRsquDwYf95qqVUAHm9S9
GJuRiRHBRu9cIUhb3s7yJrLF76GGx2wAWeYLurdHn/EQDY83Z9Vt3UaEgYLMkKBU
nfZPpaE1UITsnTIs/Tkvs+qRrxpMda+h7WUj+TJH+L5z8ug5wCjjjK6jqGC8em9Q
dfmWBlG8mUN9eVfvK+8/R1ipdXWGx8+WQaBbS+o0nKL0GJMPFKKTwxhdr24D0Ffh
6FTilS5DOzHqhgR4mystDOf1Q13sty6fjSLXlq/OBsIi+QB4TkOPvRH9MpaHmvFp
2egJxEnI7oJ7iwRZS7RVPApzkjBg2XN/kWyX6dV2XUOwQHKcTX2a0BR0pjcYcNkM
oS5kUZ2vcgxPiQVpM6z8U/oiwypyuvh49Q1ZSP0Yx9EN6EGLkDoiP7Z8qc9SeR09
fDZReV8oE3yEC8/EU1Dbli5t7QxCBSqHb0xBvLXzqZtEFI77S4BWldcDqV2HXgLO
Zc6KVNAc3nlAhplV6IiY/A8w/qk1D40H8pdkjV4brOobgqVUq3thgH12ixiq1q/b
Fj5uZ8atJ92+tn1sBzwQfjijGQJrMYgMFe9QyeTbdYpM5KoUUsmfb/HTpWaEKjBW
TllCbzA9NVrEpNK44rAPvvVG2PAjMAxVMkFE9JRtSbiuCmew/9SJ/a/nWZq2A1gu
ELM2Jig1A/Ism5L6RGZ1PcGjRD6ThTExNPuAS815XP0viLdzj5ouKmw0yLiv1Qh6
9qvM1QdR42ttZIGlzMesoIB6VNqw2LGEBu2MV3Kka2PB9N0t40Cyxsbea1X/tQoF
XK2hSk9NGJjGzjme1eNqr69RtjhDjiX3isqP2t3qjrvxTUmgQYMjveVvmvKzK/jQ
xXTbtWOKJ66OoQRD+V71f0IHcZghaKQeYPS7eKNLF+BfXKCDS6La288oAZxmXpAr
x82Xo7CPmsjlLUMDbOjtlVAfvcHSr2x+U6G23i5Tt4aXHxuVV32qPkedK4AF39Qt
d53BLIHzIkn6pcAvGde0r/poqHw0yrx6ye/JTH1iJE1ofe7rRRsTWKsruTdbXw9R
`protect END_PROTECTED
