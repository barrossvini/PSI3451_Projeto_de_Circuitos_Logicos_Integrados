`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ooe3xhWSQgKFwXNuwZZqGAv2HHd6DaclZQZljZo4nsq5yVlopIiE7W84EwV95R3s
lBfrd0u+oHvXz0AZqXoZZ57JnLf1zdHlrl1jWDopqXZgaufufqn8Y3W7uCx1PxOn
q9DfEvDpeH2LZT1Gf7T3LkfE09oaPbHSvnNTVxiY/NHkIzvqFRItsuk6T6/LcwzV
aYJLDlyWGakyV8yeKKoSW0s6Wylyk6W6XP9BpE238dPifWVEvJqfKXmtLiA7Ipgd
aLJrjRM/e+Q2qASrhsS+bjL74TzLTTpz3F2d3t0GREByl3mX6OerDbtpoj1dqx8u
H8yKoDqFwcNChoXgU7oDNUHe1ZnL50+jlGvtFCHIqJsQ0QXAQ8oHABvge57kOym9
+vylaaYkEQo3xU2ibM6PUseI72KQSTjm2DZcCv3JyR+hgOUnfj5I7ao/mvxCGySY
GHy2bu+mwrkDoceekzEyKlEsPAWYsnj1PmvK6kRFkMOTHNpV0vriBfOCrqbSxVUc
Z7SlfkkpN6BeS/AYMjKaJHIzsgjSDlNgyY/m/fRsp7769lQ7bE0TLRm8vkLWGDKv
p5hUn/aWEoxezKbOHasunlaPE+XKqoeo9+vUY59OGvE7vQP4iLuoDXDMoykzfj7R
ctkN17xooVvHFewUG8MdOyuFAc54pZlxh+iTWbjh+Mv6IIjoXLFDtC9sUBfOmW0F
MQV223g4tRce7UBBZtVnGvMrBYk0FbrJUqWPpCJAoAZ9ztUyRrFOLJakByBxYVJS
GGbEvGVadltJj1/27SRIDLBGZPnGU9MGp2PDNHctKdVD+YkXRCsKpqvv90R4B0XW
OIeyNNiommbIbTSnkn/6vV912Y9A55rmcraLUQHAgVXg3fBUOF0MCtg5AJibjsCT
+Zq2WjChOrGP71rsNYpczVRerHjOssBydajrtlPDFY4=
`protect END_PROTECTED
