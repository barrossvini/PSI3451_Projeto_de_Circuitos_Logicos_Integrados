`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EpnUjMvQpycL83NtsDwg8UN4OrnDEhg6XDqXFVwYWD2Rr6UcQAi84qYIYFpz0fxG
5djefVn8XvsMZpzm+t7e2Uy0rAHmIUyNZTYIA4PtB/onBkcpGpSvcJcYXg0ufouQ
oUa1qlnEpi2S5rrXRAHHNlKL5bXUQxnG+PC+VnDz2YpLCv6K5u5kIb+wDc25VuVl
ZyQlk+oy1CFzpo6Dx7gmDuumyABRpxuy3t0ZjC1/imz+ym+g3B4TthoWsk07QSRQ
QBdhAEn5/Iu2ua28Rc+uv622lAUcOw4QbCx1mpv93tWlZiYTvrL8svb5mdhzyCSD
MBMBjjQ3SA4PtXyXlj1oqX5vn8nwVui6YzuNSkVw2uyxyDKnf7bHMdArJgu3caqC
Xp6M0dQek8dvL3xeLO8xmeNZHqXLCKq06d3hkYc9A19lBc0rBDqnp4ZLJt9KXKng
nLlJJ9byxwz/wILNzBFutiTsOD18+QuxIpU0R6zaNFg=
`protect END_PROTECTED
