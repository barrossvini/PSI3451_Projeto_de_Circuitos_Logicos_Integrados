`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3YUXb0zhv9Y1m1dzufSXSKOX2gfTVjjfsfN2CAaCaNN3uPFDvATLvpFLnTR8X705
FUcC/91tkyvXx5cTQWKfD28vX8p75Qy5nBK04ckCDlYxIUKpmp1I0MTmfOUG83ft
v8qhWgsIJwUxh9I04dTgr3xmF97X3vI0v1rS7ILvMyfSXVxMOSFRjAGt7EImjGgK
xY/VTmfJrbyXKUvKIxLItm2QIfR3qhvPF7YXkJYPt5NNczCWvb75L/XVXcGQ6Fef
ipV5UZukifjQnHiHRUJXel4gkqQrdPv+RPl2ghrBwfQjSutsYKzzzpOU3NcPFKdr
WMR12fW9scxZIaSdN0q9u0GbOyzvuj30cD6yah6ZcO0OlE4syM9wI2LNpURpmPEM
plSFd39wCnXBNZjuheiVOlfespJySKiKjv6EwHLvrhM8OqTIH3l1ZebpR/z/gYhT
pU7vp2eh12nyKPwC5mDs/XvQLX8AnpNFT5KOZR8R8r6y2tpJilIXbTNzBdV+SiBd
9zDlHCPxNghT86EbnXmPNLl/J27/vm0aEExyLJutz5CpgXeaU1pp3t61erBO+cWO
L0G3dw+imSjb7an9NQpjdi2O1mehnpJwLsfHkQM0a4/xUwdXnKywRNOKb0bqlz25
53+sUb8i2s3aJHKfaH+ZSoYTmQKP8BmTktPfURC0/6thqmNm5AAgjSweJAUdQkIu
KsmO+fuZG0LQ+o7epicaw4biEfEKUFPKYKYAKI1bgaSY1zWMO8HrqhvzsQqwJOeQ
KE9ZNfB9TCwIzImy3sxL8yWnXFwU/+zSCsWVQaiYMPPa+sUtzFHjNQsatEisKQYk
OTsritzzsSuoz8ZJpmD1KVo/yXhls/dDJjJL5jhULFO0YDMn4S+V8A/bKtgrQblI
B/6Z1LWVrWiT1rpFpZ9ioj4XogxQG6GwleoXPzn/QhZO1r0agUUlt5hI+Zdjt416
ZmqWCeKkd0xfCOwPrrZE3SkW13OSRcmIsLDRr+aWVm9HG3HiA+6hnJ46YwXulUfL
WK1tJZ3MPsKo6JRZnX/HizzYkYrJLWFyCGmo8tGFbS8JKwzsJWtE2gFC0aPlJU0N
BQhUlpfepmoOA5uwPsE+StQoUqqQ54qsVGpoP65yKFDkHWOHSJt+03z+DEkWCvna
pFQhl2qP8Y4kGDQWFGeYq63mu1qu0L1k0IORoxAwy4kHDRvEWf5HHvP8DjxUPShe
TsLdRbEexUirunNQKcB4w3t86AN/txWKayrIUWI/MjJS/p9jeYFBwhRmifB7fw4c
vCgcRPTwAfHK7xNemtOr9sq5KmOZk7tpZTfyGK22LryLbh6J4mKOaUGPj77eSkyK
6fv27H+xvFz2MsrUMIsu9qLeaj6IIDMxEWt/Bmb9fJdmok8dt+Kbm+9V2x420LXa
OSUnPWHbvijbYrgUvrMPlviSq0KiRvHd5pI8YIbMu7saijizkxgpGUWiAPkrYFI2
eX4jkPQiHcygesDzfSZQeoKqysVxnHOPgzgAjug9xgp6h/kfYfGoTOsMc2GKd+dF
MNc1nKmh03AUxH7EFZNTQ3vnoNM5XQJOkUcfwEhGeCB60qNVlYI7/FPyq1PPBfxt
SSRzSpmV1/UZtmtqStpxN/NF7+c/wmzv3TTneGe1rQ1Mo/HGICH5NwZqMsoucz0a
xQA+AW2BG1OUnqJKrJFs8EikX0rGF5GKf1tkzkwwzDTpvpRuurY8LLsd6OnsMLRl
wASgpB0gy6OjQ/qIEsH5scBRME76bwlWcUY9dT+7A9nDPJUwq6E3Q9/Yi8llIo4h
LPs0xrhwE0sk7klNTbCP34ZxeswkQPS98DW2agsylpHAxDFb7tlJgajT9lBv9+xk
uic+lB93FbEZwIoDNsOWGoJqIkXD2bINR/RzTterzRfGA/f4tz80s4i0CaRX7enb
DcFby7xXDpLePANvDxz4cAprlyukabzcRHmCeJkjsKP3neLEAztLhs9kbEF1PkE2
qIT7PnUadog7mXblepjHaSeISwJ6AKnEN83mqKbazs9DMxBBCvcplVis8am2R0Fb
Bn9hiY46BaciPoli2bGCZDcGY0bPx2lfqE1k3RB20VeN3HsZEtyFCZhyfLjcNT5P
NwXl8H3YGvmwXTtjW1aIXFqq6HExQuTXRxebiijxmQ+9fRvC0acApBeuRW9tU+O1
TXa3b1DnWdpDjSxGv1OQnJKJ3j+I/FRIrnzGFH/gkDiYjYVGihRThlcs1KY9wwu8
BfVbRha6yZlKh5fxKkjU0iaL1sPPAhT48n86sl9MSbr+fx7G/FEB5RBARF1F+mbH
CyJFa5Jy1ZMRuESGC3CAkbFIB3wKai84UBLDFNxBgqrwYJbw7hX4+B1tDvBvzlTg
OZF1NxCIvR/ah9g2KGfCuiKsynAoT7U6BQoUNmahWv1XDnaTkLRvWgo3AvgaISpx
ni4NAkF0/39bxfDHUfK3UEZKvylmDyXGlKtUMOp8xnY9fR3h0VNsBrc++pDdMpd0
L1tvp1PnXE5y49cacffKehsnW1KDEL5hdCuDh9/tjc+4/RjoJss12we+1mGJ7lBj
0Mo6yvqKzFLQ9VqjUH3nn/qjP+oeIvQ0S0XET52dxESqC296XaSCs+p5Qk5CJFA9
nchq99Y7VM9qcfo2VeX+AhluKTImFy1v/4t1yfQ0UBSp/HJmMeaGnaDgkatngNCb
c+INa6DOhWXeXfWIgT5di9ovUmPNh3SaUglv4t+Wv/Jc14B2UaoAQbvMbGhkIK0F
x0YpHbGjrTNQ3N6zFGUo8y6qbj8rnMchGIaUtL9bc439FTCVhHnt5wz2psHuKVBS
6KX5fq/rmk8nUuW4o/OHpS8PCl+iwTdiBht0xkuSR6JB4NKwSPY/EC7UUn68lnJR
PLEAvJCRWTliH4NI9REoznhOfRtffXx2nQKNIwENqTXssnZ47pTS/07KK5mzeSH/
8WZr9mRqWREmcKfzyoccHMr+4YGf4fiWm+t5pFY8wtgy299x3eqlvJHGNjMoWMzS
FNt7M41AYHel1JBQ46ssQdSYJMQqVC1UubSAJs/7u6VaifxEiNkMNET71HBjs7+6
yKqa9VbZe+OGfEpUJ0XeZhGsw1NIxOp9PfbVvcLWo6+M+UO2vXxRwPI49akw8c65
PViK6KYoaHrKnJTEiNRtA9otbJjJybX+sj6W233CwbykA1FlpJ4JrgJ0dXUMXoOS
i02x1NXAIR4Qt1oL5QpXQ0KRulclrsiaO4lYXNJaAkgHj+AptEzNk3Nu1Bl/i4rO
JhVT4Gi1AIoRFfJupkbSvKjscGtRiWII8P2rb+GKYD0sHROyw6CGX9PIUVYat2hB
q70Kwi4nXoXKdTOnHQzywvg+Yi8mX2FWlo1WsDQQI17qejKiVD/8EtDRh6tE/0Z4
AkI8esIzZK2wwMe1WMn0E+Z7Xt/xJ+A9ugFkitmyyLUiA8M07H2jBFZhvs96wQW6
DC9kAnbqm4X8h8cLkUg+6v+B8/Brb8hBolV99WV3oVpVqRZwqomr2q6h1T4aKAzu
oERLFlAOEtENq7Ysq1uhgsmGwxTiLjT0NziDdCX2kIVb0uNrl6WZguFqMqc9n6h1
p5nmVxvjhkTkYBew/DoARdcaKBff7DNpCB2ENkxBwlr8HBZjIjOuwlaF/jvN6JKA
2Z1lSg6ibwmMH4S4BiXfGpB25rUpsFqgXJ7mQW1WW23ejRfzdY84SIUE8VZ5VUQb
/vK588/GEauPB2zWmSbzbxdl50FSKWzunQIIS9IIXJFTc/XbwTZwMkfIrvPA/BNp
cYZdh3MK5UL1Ud8TTGB5YP6VLHG9mRYGS9FpE9vCkzRDGIqlBgFAvkpOnQMD4ru6
iqN7Zmrq8u04XsmS7jGM4jqZuKssAO95WHNCohUQ0dMzUwvQFvoa55vTe7PcfctO
eu/7rtqKZLDxM/ehghYpZiz6+cZeU8l3Tf/y11lJF1gjPbiCP3+XLi2VWmDDShUJ
tOimVf+HVuizhXPs0TK924BdCo714ob6BN5+1AConrUUN5zAQbI3k0el+PHDN85H
F2K6+Kz442Btu1RPTY54nffRJp+QBHmksg+uoOkbQE09rJT9NLJ4oBqx7tTHqME9
eH4x6plmQmrfrsU4fTMkgVNsaf7Xa5PFfibCpTkwI5U/Ll621B3wDVbFIpF6kumK
xvtOg5c2vTjvnWkxySzfft8DdNMAGHgeupl60c9VQx6k3V8WaIpM9/z+X6/6k3KB
d3kbIlpc6wWQWSJpQWrYX4RMqrHyEmFXAd7Oj+YRmBNQ6iB+AYGP32ehYME/DWME
1GZNMov0p+E8IcApQ9ihUcS4uQMq3MfXP6MEZlmgB4MB1c4j5eZicH1bF4vWyl4K
maWmk/6Y1IcOTB3IjJv5m/qVyydeSaRQMv3K2wgQEFWf7kxvio7i/Je5yuVNmQk1
9HJGRbAaDxb4189ZU4l05OpCxa2zX1XIYO6e10UNChMzYBc0Y68iqQ0xMqwC5O+c
9o1wq6Ue22iyywLnRfDQEni9oUJIohEpXio5oAPExJfjXFqD9j5KKj2b062yd9hv
PeSZdG8fBsDnSJcgsH4t4FgFlOm/a/O8bG2UdGugtqiQpLjBQjFV9MXwfZAxMMAW
+QWLhIRHshzoksrc/a5QNOXdgyx6ruMEJbyQ20G1QNPW8Zy2NEXmuco0xLFQ4lLI
vV8frklP2kUnIdyJYYwMN37e2rD3o0SYynlz+u++uZz0DXxzIluRilwo7nC4uNbi
bO0v0h3T6b7EvJoAIaBUg1zHaqqCPjuNxkT1c2Od9eDVdoOoZO92rXifVkFFK5bQ
M1O/fOAg7LmGIj75sQH8fxliYzSXMbg+5p8S4/yjUVY97E55bacoXKnGgJm5TU26
kS3jQ/H/T5QODO2c7RoLdN0hcEqFP/jJXYdXZi7v7E6iH4QpNdlXt+1mtBrWyIQ/
yFpmfjgM1D0arvOxFCBHGhQNntPkWdPckRR3yEX1zeMzLDtgtMg74CbvBOuOXgbL
gyaYDUOtOi/tYQ5Du+8T/Ohh1eD6iS+ciaRyhjMEOsLOzuIltq46r/O3VVe+GmIW
odTwMGWZ0tDt5TRmOcnImtlzpWGVG6OO6eHzqqxQEKaSzq0DZx6IDZc1qsEG2U7B
3Eacd9Q9ApnodzFSV6T+eZXd8mYG2w5nxwj+7S8JU6kcvBKqRVXtkRbzFqSwHNK+
A9klze5rK3xHvJLJuQtWWROvrvj7eF5T75JDCcMEd3is8Q+KnlJrIqwpw3gyVyQj
yAvTpZwMQMevezuaadIbFxGEe6MowX4LgmxBnFHPaU7hiQjQtAcLw3Eu5Gj7+Kih
yuHzeTI+Gi53fsJrLOUPYF8sxuQATjUXgdNtmVic/1Fj8/YKUJOfRqW3yhLaa0Vl
ohb2we5D+uPUlI7/X1xhJDnQpOxV39a+gBA6UJODSFff/3MsOqZtVjCYTexbJeRh
ZyY4/aQQUfmLqP1NMlyNveITu7lpjXsF4gSp2aO0xWW+tE1mVKLp6xqjZki38Ld2
UGLnq6bQllHGsugyC+wCyeTwErM2DnVLgS5d5xRjbun3jfEJcHLP6nqgtD8+7nqe
lBhf051pLZ/ZShu0i+rNr3+KGXl9ihj1IY5UVp+b2CdQAYS+KSEjbfVHC2fhGsX9
UMHwD7+iOcXKjB2oG5nNkPY6s0qna1ko7a5wk7XlNS3o77Ka+WIkfCvAnZ0HpCOE
tFeD1zMFIvXC3KdXaQWBYJkcT61i5tKozuKAhYoWsdKVBMQ/sQoE4gDvFbCkvV1+
fLpBXfvU+6nk7O5Rd090YbZruYC/CWfShBcL/8mdGZRm3LhlqeFU4JvL9f73DHD8
RQg5kudHkVYbErGnSZfNdqIexbWU81KfHwo2pM76Dz3qwudDSBSXHes85XWifiWI
UhxkzNoc0x39EpQev65hMngCE9jGzBhOQhUjxuzwey1UhSYmAVAWXBZg7eHMqngY
zTCPnGkrlugygRG9v3b6zAf3jUhWFm7r0PQFRsumvIdm1Svtt1USgUl4l976DF4n
WjoY8/P//pySaIQ4nyzm/GLSedXKT2AmUjoKB969Z0AtwmuB7iL8BZy0a6g7Q9Bm
nfc+zB00o0VViagr9Q7vlxW2vErpLVf1rGCkpwtTLeyJGFpzv2sS7dFSxWO6rcst
M4il+CCCGikyFPSPZSlPpPA9XwvtydXrn9hifuCnqZidbl2s7+JlkCqA9aDKYEEc
oe+Sbg/FbCNc4yaMrDXog59HNAoTfaGc8UoDiwAhCfzKNAbTcwmXFsQ7FrpdkqQ6
rkfWdq/X183x8U9aQ4Naj/6LZ1VW125hzXAZnfXwlRrZwlBvPkggzoVowLoT4gbi
csE+gEKvmpLtdTOAYBPFHUoPpdDddZot1WrKFFUsMrjD6MsbXWfycJ3rNkZop0jN
aru+pnFTco7KJ4CBOh8KPEeBPaMX9XDSI3VWHAKammy4v2nU2BwtEqZ54boqTC2h
DTX61WoBe4eFzr33hJuTPSpnXuSqPBlU1PFTwfCHQjUuI4qR5ZES1/DJl/MlfTC/
raiIGDRuUbOV4xeXcat+eULEiF7K4+iyJuLKLz/z9QvsIe8SqNr/1vPePftCEnqJ
DF34327g0/hw2Wlugd9+2kT/FDlqF0XA2cxXH+8+LEELDYrwr1I0f4FG1Ypnr6Sf
8zFRjkGP9M5s2vzJBNmNkb7pwd5oDx+shoZEO03y9P2zWu0bfFll2Qa1Gxl1EGF5
rEigFAxqvipCLrZaZbaKFeVWVxAjSazGXLWSqNAF016VcgGAWhNL2wYdduWL0Qwx
OImm6rej56d9CuBQurr3tn3JpqWQHgDkW6LR7o0zXDV6wImYpLQfh+uT9q1kjWqi
ANgo9qP9kiR8pgHDIr+v8cbEY0tH8W93U94Ce3mPc8TvaPcurHpzNd4nN6+Ch1E8
shMmnBaEyMxKQ5FaaEoMRp8uco19HVyR5OGIuigHZTF52y/p052ewozTbkEcMUzu
AHUDmrn/tP3fzdR+PXCzVi58gf+Dc49rJ5xKd6UZje3M11VRLGszWmer8Rd4Yjnj
uaKDeo9UEEsxAq9JApqq93E326B4XRSw5XMlfc30YVC0LUdilpj9sEwPu4f0ZSEc
x78ztvhJ6fpoeODo3kM/wrN8vtNcM8ZogKBp9+KeZ4NyPBFOhr2eORMoRnUNBZqw
ZMLKwNhUCw4qQBEW8i+4lZrlfvMM4VwAoaEkwOeSuOVWXHeSjqOQYR2l7IpArAiJ
HvWn6OGBoVofP7/rpvf8l13aMeMwm65AZ6bJIybr/SvreLuS7uqQsce6OE8szsSX
R/W9ZyH9RXrvrtkkf+Jmaki3p+vMupyOND7ku26Pnrrn2kIo/0YoNSFub6jcYkHi
GbSXY6l9MNtnD4FgfILcZQZq+lt65dHYtdJDaDBzZphA5DO5igejmiFBRXDbSRrE
N+5fgFeHR7cP4OMNouULNN4pPaeR6+XFZFuDsvxzSTLRIUv4n7Wd5yAeXPOWQwBc
CLYzL0XcuDu8e8lgs6VxgLcbGmWnW8Tq0Vfy5cIoD6tjDhrsY2bE/QPNMSj4ZjWp
JxAgAi1ZPbXNDMFZdwq9zR2T3k53Wuqp2tftn0wulfo0SkCqtgtbFo6WgGx+FMoZ
+u55Ca9IqCWBDTxrhII0FD1H9d6swlz4xTyS9a2ElJ7cUoV/U8SZbKarO/J3CNVm
f5TpTbQDDTVHxOjpQZp1FgBQpX5EO7lhNvLNvu3RzKlJpH33Lz67uK17F+NuR/9U
aEcFMj2m6HOctSHN/0HBPA47NfN7e1ud3yC9FpzZsHrgG63fkeYYmo3lNqy98jlK
t6A8HlzWmkUO4SbTFpNi+5NNLzFfaSTLhRwkVZIZ+FXyPe7RATeXTttFgdAfafxC
GeKswmC7eIdYFqaaeU14+F1KJ7kSkssZS115AhHIC4b7eUv/zUIHoRj0pr3OQkGx
uWopHn0+pddW0z2mNsmzJvUoMshlnSBNLiae7IM0skJ+xTtaxptc8ti8QDujtEFF
+lJEZELVuCEnIs7gv7D8IFHXoJgitqjjz1KzJFJ/CX513GKEa/cvhLtvMR7yEmfV
oYYh2eLPBm+eVOPN4PvCO+eh0JAaJj2suf94btToqKcWKO1nZtHxjrvwh2j9VsMo
W+nKwd5TmAmOvjTAIWy3Vl1aijA9z4pw76JiS33sUCJtlFEE+GpILx++Dd+7Ptpy
HhJHnhwSMWhgEiJd6LSzcEvQ64sWORFfETgK378lwQgDrYEHuVAqVfvJgcX+EhLL
miMXECTSnmVL3sPlB/NUefX4tQU7Irxgniq77WISrhUAg0ICS/N9z4hSStsDiqSe
CsdblzsAKOBDODexVN7ringrLWWtw7rdF8DCmxCkYhLEXIpmIWKiqGKMJE//J8BQ
ESmAx8VqisFv+JYOVn/vi6XsiL72w6fjChv6FYwJgMV7wVHc94hAAdRZ0cq0eUV7
iEE+5kDHAcaeizUXiZ4wuyGVM/KeNJasjlXhvf4vH+bXU52ZQu58ybaSej+X0gVq
9oslT889N2PPiil4jyJ7twXQCZuG8kUcuGTDnGQESyJwsZf6ZLq1F50Z9hpfr/DF
/Znd+ngK4C5Ubwd6P8in17VQOuPIFucv6DWZJwT3r0TybSuOqP/p/oU7KSyAGzLM
Ri4IjPcLW+lA+dlC71wAGCdAvT4zd7nOZIuxPkUluz/a4cNimm24GORbjHRB6RPl
BxqNBvq7tJQj1C7BYwPgS7+ui5YU3KCnMiNN+S6MoPSyUKvC9L7L+GJYWNun54Hd
xyHA7W0MvhJ1v8LLSZ/4OQfX1shyagFimTMZMaTPOcvTDv3YRuuzN8+D3m4MTtw+
BZWAaUwMtN9FW3KfEi01rN9wFN+lbAmvzYDEjIZHhgsICNZQmW1ahm9cjt/dWHpc
u86UThrEolAjkkQw+Nl7CAdelM9fAxnA8/XrxTt5e6pMU8xADDNT4g3ghMFMQ3Jr
Qk8iwjhENTo/dafIqiOEQixxrdLRgO1dOzsGVV7duV/WLo859bTV6+aSV1xZRkBK
2jP6jVEQnTiJC9DJcl1o5ZF6Wk2J1k+HRkDNPOvGpLGA7OD2fkqY/wQs/daTWd/w
Jx2MbAisB7Ko2Pvv5rOMpXas9f/UX0xioScLu71K6b/m7clsOycL5mpkFNd+rkcV
YRTqLPIZ5rTLap61irgnANC6b1CDtPM1iW3XqirLyE9lkoG+kjcTyoTe/qx8zXow
1YJtqlDdrCNco9EUGCrRWm1dNDIlkJ1nqec9bPIaPRfVLvsMxxuIApthit50b/73
ibB+kS0glEloBjn7uPTGd/03OgYfYhAwsLT7ViArLbBo6I4RXJLx7ivHyOYgmdrt
awFiM8/YKk5wbx+Wt6vtlZqPJYrR1ZJW77rETqGbAQajiNF9anbulZhzzwFmxfsH
QAUlQY8Bjmi+yFT2DNIeYdjAe/vl72X9U7cUxQr9ecPlIevn2cUkV6J2MYmTDYiL
d6iQWS80Oqv+j+kJeObuDvRbT2hJZpVhDnaAihkWJQrWWnU8vvPaNrAqWAATN38M
67MXqD2z9xYfCgFqIuXapzhpb8cIQl821jy6c7tNydbPMGMPZSKmpcPs+YeCA9iK
4+tNyrcppJiqc9AUPTZ5r5ilErUCx87cTDTsG6Fn0pyCkbnJPMGBWpgk24B87p19
QY5HKXjQBzjKXMRdEOAf8Te6IOPUl7jq2kCEF3lHyT9PiT6ZegbZmcPuQg8WPLuq
1ccyxVR4rKGUOw5mYYtoORDpH83R/NvQayWf0VZd8juBpGyDIvdckSBbjAkTQFOn
HDst3zeygRJXucn/YmnvCNLEay0kF05ovSRWj5jPtvVC7YHbO+TKQrH6m/f2mXD5
b9sMIHFKTn5WWPlthe8akoxSQIdY5Wo2Isp016NUDmEVs0KJOdZO1SK9fh8h50fO
t/x/WBeRcJmv1Il5GRHAZWWV3G/VPf7jTgsnoHVC4YYLbH/JfB9w++mRG1d9Ao+/
MhyDiKik5C7pCrP4rvrb7W0g2SzHTx+3wECNReua3+3GnvOXxg4eL4SNsvjFAiU7
twKStePF0qIHs+nbcXMjYow66YMmkc4IoV7Tox+NX52udNaJ0QqKVlFN/BhMiIZV
BcnOtZ+7/SX+fkK9hsjvkC0zdRjIZPdqxmDJz0jcia41whrihQpDVTbINgs1is6P
rVpNajgzuMOvl3uejkYMRQj7UKvs6hFDd0phIb5QbJebaEfTPT8gW7zNvw5BcvAt
6B00/yUJIINUtUZC4YoYTGWLg3GDIqtJpwQLeB9rXPTPzmsXVV7s/tpq3GCGORTv
v+2NQ12Ip08/84oNBmnjCjoaZzcSaQ2HeitgOyHZNgJnEN9NJ6NJyNzJqZiIQwfr
RANNlsYPtrWr9HlXY9f/LeCCPUmCrjBGO3nU3IiPEw0Bbv+Yesxx6MskH0qyLYTM
or3Q11oxS7vKkZte7ED/5Q1l/4Kd/H9FDjGiDNhmdilNPnN3lACPjlMTcOk7zG2N
2kvU4F9pvSZkPPSNgv722OyxhL8OjVCtKtYABUCi64Zc5oZDrsbYRjbNSwjmVrt2
Us5WxkY/mZrRkPi6/L3jHOl4fwwZyZHDaaU7EeWvHHyJ14aECrh7aFZ1mj7KV+X1
U6+2B9bxHTJA4Ade4E7bCyfwpwyat0/qWOx+bWEQL+XZINCaXnN+N48952MF92T6
uKXniMf5YWY2Ucm9kAXxf2ploCzq2f5PhZ5NcGT6SdNx6tUmAxhPNb9ZMco/Ddg8
ukMCFNp2exOcpnPN2W/aCFzw6Yl/7j4dKcVJlfgnOSsvtu/7dvOQE+QscxaO0E84
MTM4uam/ldzYV+5sSjusJpCG2LiTWgKagCHzBx9lWRM3IrBsQGB4W9yejRWzS3vR
rN6rJyEUxKaAO9LsS+hgsW/bXaSQ75Wl9S3pbQn5CDEep74l0hTgOlqpebnqNuZw
RQZjKHVHfG5ak9FtY3yErIUjwz8Iqdv4McQI5obhylgmPKbc/sBnVRKXR3KVvyTf
2UaDZEX1nJsnT9Zrvtrn+/JzGvOTX2rt9+dbpZvp04mTewA+/KZMNaSnIIcWO14x
zd7N5Pthe4b9iXZtzCFiFj38YctqYYzTV9H3QgXgW4JnmNxh/3gCPjgOCGRwaSQ3
nynPUMozq0HlAcExYAbu1BQhkPFqo0qMBqi/9uWGmw4WYqcCCS9TdSoM0wkQZ8mj
kbtyjWLt5bdPZijdnIEJ1/jqbC/NQ0khE24I8km/Pakjy9kQG7HrKM8F/+BZTt+U
ieMy/rsd2vgh1np98tqArc6BY/vAQP0ad4ggKG/LC0PfS8aeYn19z1KLBmyOpBFL
1x0Dq8MI9RRopZn2YC8GGjZbgjEAKT0GRi99VwL4lAFaaW8mH0gy8mi7QM9iNMJm
5XD1y6/eQFbSDSjkiBtLP4X4A1jnrDUpB6GM3gtV7WiAkz56qHouRR/lkaskLwS5
AELvJ5Bxo7qqwlQlnYMaWuTWGy1xeZ1Bwf9asf5wp+KliF2/J9W/gaSbbqLamP/h
2d/GkG2sz2Ry2MRGdbMQTYkfAaLmh9ArbZw3s828GJKomWHMwE8qoedmpbs31G5/
lq+TpQ0AznAxMHdoT+xe3vLgjrlaOKbcnYbbFrNtkI35Y1AHURz9NKkshKroWUeE
KvK7v/pDwrPkaQ8qqHGF3FExc2fphwlFvPlPZJTyKznV4hD7aCC830CHWpqUlf6x
03XG9MVLRm2Qok9z0lYaf70z22jLm0DQ7mLIbdexKFVLwwDZcCyGBFvHmpxRsy3c
FpkB8MXtei6KA5z+5kax5toY9HIVZETHdMgp6W2thxAnPUKGaw718e8NRbaNoU+l
Qm/CQCOy+F2PIzxOyF6wCcZDnYHS7i3iFrCerNJ4eOyZeYdSgjl83sboTnVN3WYB
ZTmNrVbYBR0vj5jWCE2Umwg6bbVHjvmzUZZvtuZNB0/enWXW9nmBK9uFzpSZjJaD
50I2JqE0ydGxwazjc9Uj45McMPnkEB+IleSfyfJzdvJBeD1xfbE+1pADMxVDSFpi
TfjNJu7iclX+k45scEibGGucu4s7hovInO4zjj/TcDUMYf2kbAQBM53l73ocQE2C
yyPAFpWdavRQzjvyZ2tPcwuggNSm0iooTxGrUTHjj3QKHlTjf+35RqI2rsaYNMx/
1pML9cn0g+iRz7U+1yW/1CbAgjqxkRvsMGX8HefuLwAGadExmDxXGZQjolvB6ppR
Q2aQA31nosDgteWW1bHg0K9G3texX53f/XIFNo3TCvEZLsywnc0NtIjKbp6x1Rqf
TuDJdZR8Uo8Qk8rEeWZieQqTImcm3tv3ferf/Ls2mqkSPmXyqkf9TzbQ3vWgC/oF
RXTv7DQUvpbRTL7pxIFsincB1SGJ2IG7tOl95AlQqw93KS1AEgRvsdfg7yohoszL
Ck9Ay5d1ObFnxPO1cdeYLI2hb2Vd553bxE2cd5DY4Wj8dO/5V8me10Zizhne7ChG
6SffVoDirEkVtQytPXSbC9kTnU8ratKFSHFF4rLfLk9TUH/c2teSSNz6i+qD1IP/
lF3+N26eaMfocuzvl6hhoGJ2+IT3jw7+DG9d3ad/iIgDiZGUZykCTMyxJIbq83oH
mUnGpxzmPRf1ImSQsQ3ka29DUaMq4XoBo8O3rDJxcgj2vOZIsbyu3ccXVr7eo/Q8
mlwo6IEgKaU4zs92BF9g6i9kt6b8ju/DhJvmkp1DIlsNcWXqlX1/Ky/75eV2DpxH
6zfPjQvtCewLLE5AON4H3pAW8+czCgx12v2+urlknYuojnVivQweTKgmBSr+4F+c
wUyPa/DC5mMXwlk4/Oxq9sWpnxwoMbP39zQMnSHlFefoPrpvbaGzR8fz4yMajVsC
VAaL0Zscs5UioN3pos2EBJ4ETtm2la9L1GsM+9cng8Qv0bE5txgeL7e808cPeftq
jSk4S3egMDGYyN61oGkqloD0w3HpFPS+34EvKUKAycG/r1JUH0Ozyd7XASOFLU4f
Jf2u/m7lJ4Wm2N7cKXbxwudUBHpnCAP1/8PwxFy7VlDJfi1jonA/SLQcfGLFxGiV
y2pkX+vnPCrl9VmKmVx1Op1YryJDG3ZzVEzoqze3dmCpFa2V1V/15i45J6UuFBt/
3JFU4rWewOeyLtMKDqqqdQfIzlwFvYf+fd2oQwrpxJopqSf8O2jRoD2cHnRE5EaN
ogG1FDwr/vrDtqPECkP3zdPCiQkbJStQfaIvr12qP5lUvqdEMFk2lq/IweC8FUFL
iExjwLlYndT+6wa/EJZVEIn4UD0uyAHzkZkPvgSrnvMSQQXTfviX9Whq5/sO479Y
2HmuuE6zClGumc6LoSHDqacEbBe3F4P5sDCIlpaihY2XjHlopEOmgpf2X7g+Ee1h
V+9R4AxPDy1mY+v+vugm2fZKVby6GaHOz4SSDK8B7lqqsBD8VRsbk3bvw4MM4r+Q
yGZaWirrvrPKC+2QHc5FkAlJbSNJLND6WQmYyP8SR1nIeNjmTD+cXOWjx5uyGF/i
FLgJD5BPJmy4E2gHWDvLvMVwWOocUCKVIF4YCb7YjYVQPerBdAaCfm4ct0iMoEvq
eHiuMsfsMVKB/kR4UGGsIykjYIi3TSIfw6THq1ZeELvbTIpJx7pquJBIHB6Vxl1w
kBTVfh74hTEn2IdhHhEqEb3Byx97e4VMgrK8G6F/DeFPXQeneOgw71J+6sYzrg6D
vl92vCYuCX0KL5TTF/A4MdmzzFB3vtvlK97TRgv1b5AHVZuelvCP/0GEiD3EnKjX
jr5mlrIk1ljfm1WNoHk9Nh3fdkszpyPy8HIWsi+IbiyTdYTuBEwUg3ZH1GGlyAyF
X8+L6e6FmK+LYz+x++r2Tfn8eZeWJqEsfrraY4RTsITiJbWbvzPprMyxxqmbHSP1
MRGRILNbJEryV1ql1GGnqqhBkxxg3hJMlpcwZHM4L0XSgJlNv+ehJuW0Q2O/7foT
B8xuorq6OAvNnsX8FqFGw2vLNVz2o1DKUl5NHHdQDDJgF3bpSheJWt6NJBmXEXsG
XY/YWYvyher+ovkbmxGVDfxzT1kQprl9UMAIQoxJWlitxjPpjdtry+dXtGRKpl8K
T8aCx7m+0Wf2wjytaRWpID1Atd5cavpV6yztvZ3yDsMZyr+ilUnillOY2VrlGGqh
jlKdsB7JO9yZ+p4RuzlkUTCTliRDIvho1rlLGHj5axHuUJjOeGX/PD7LZUiypBrF
ZeNCBhKfXp+dn2/9O3KP9BbvuHnyeDP+c9e5NU04cJZbMQPM4+Y1NzJzBIwYa2vJ
kgHeXQG9DDAUjll6hkyv9jncCrgfTUxHEFoyQe3EY1B3WAgqzWf024gtsG3ASARJ
JXzGts7qc/Z2WJfVswD2xQK+93VuiZLYgJO/sCn4Ib5x/rvgCIyalr2+f+nFiEP3
MXWCWyU7EjmtqOrxVqqO9x1FHGLZnpSKoxTbFazKPThqC/ePG9V3HElYSSR+wpFT
W2NX9IG7Ud2lzZBt/iEwx3blPWP5tBB1Ex2BO7mwnKmO9zcnLg0sh7eBpQvFyutr
M/SJ9UZpfZ8Zl/xrhSUBFhsYiwjJd6QxN8YvDBdutIV+aDqIUAnW4ueRix0gUUYH
1t7hpRrVUpaIWR3WboOT/urd1lKINkYq9+lS7RLuMyyvVYg857VUTL6HFtn3toL5
FBNWBng2a7y2bsHU/786dZBW9ny6KhgZv506pGSfl2wD6tQDO6PY2bNR5V9gS52T
alZC3swfXG640fhYeY76KB8pTylcsTwO8IWcgOro/q6nxIxMmQzaz4ulLOU6StIe
YkIxLgFJhwl8lYbwzhP1X9qKuZOXPAqwOS6eoxjTHV/MnmQkh8earRmhTT4Ud/3N
u9cn4R79wwAyj62efD9nMvA3cv8Jax3CppaqDE0thw+/rrQp/qN3zHTjj1e2GpfH
Wx05H4IUbHuonKL0cTOhNZ7NHwuXl2Xluf2bu7rvSCx1qlGdUt99bFmNPLTzTnuH
fhcE26Oi6HZ6uQ8b4ibEgcZbQKNX1hQc+rbQJ5Hab+sQ2kq1O42BPIj75V9lX3kF
6IQyQpwEcK8shkK9UsqAloEPeDJ85FwaQ+xbYta9dUpCrtjX7/g+GXo/VzR6QFMC
7Cd3jvRQyNCafrqFBz2SeFXXSnyER0h///6k6kaIjYMSIrfmYjeleQewZA09pqcL
/+dQaJe5unKbaUYjjVRys0vuDWK+c8KnR+IyuAmtGzbAFcp9XeofmNwzjNU5t3rT
EvujGyRnXi5w/pxOpMCDxo6xvRnekaEjW6uqJX1QHX3DMzzHKwfZpmUtwqGjyfYR
jwQijsfQYYyGagAh7N4FnonTUB/8g7i7iWZL81LcL6xCjoZNbcS2+W7dl1hbUTXn
3knrRrZVyVxcJNKp6WYjRi1KsMRxPXoMRH8VidmUoJlcUj1L2UmGOS65M6YFUtR4
VwVkP7N5rnaZnMe7RZZcZzK33DFTH56lSoxnMD/lv/5WZcOd6wYyrTCQa5p1N2ar
xe6nA4nGLj6umLVX2FbhiovfLcnXc1nTJWbW5TtSrttq/EGusWtYnRg+UybRq9Ud
Q6/ljYF4ArVolvCNOlP54kUmsKMvsNWyR9Nh2J0PCHH6mf8Y7a+prAmMFTHZfp96
EpMfGmXOzABFPVQsn1MnmAnIntE1eo7Y5b7sJ9utSin2RmWQutSboHR8nQH+MLmk
62rgT0taYt9/Ibwq1qLJkaGRXs+FXznVTy0fLIgsjf1rNBLHHQ3G3igjBm+9ZUqN
B+0X3oK2pkLt2/0ZI06cptipTXYYXz7OpExZ86ZYjHioyVDiYs5bbcSDGE19fo+D
kB+JWxR/85qMRtiJYSQ+Bw6VvhrZwhwxDOLmBo0RE7nsm9eiM2QVuCPv3AZB0bkT
3bpojbYaj0KwtnKG9g5oghz7eNx/qtJMW4YFPM+Jrh4FUc1AI+7+V2TPQYpy9cnU
bhSaFiTXXptqBl00dJh+XoP3jH9zZFsdESuE/NIIcGCzCWQ8cbhN+ofNnaXgJ/vB
8MZElW+J8bZ25rLs1wrFENXMarLDASa6oYJkz4LNKoQCfPKYmf/VD4argPKCzGWs
UyTuELe7yE14xm3c+cUbYaiD9K+m71jTarG1yG1fH4q8kMvCnV9sk1p9iLTea9l6
99OF6LauPYWrACE8jUSea31dHANCDIJnbjt0o6y2dsqxnMe2993THMHrwzHM9tOz
OMv5jbaMRVplyoetLMIyF7Ej8WQwqigi0fcaaEx739cJHGmaW6RcXwwjSlpf3FAN
koD4PWtI5eT+TfY/R9C84DT981hGQ7E/5ImFhx9wBBrNJRL3fOsmpJE5d6IllYJv
7JIXOEhKM/WWGgr/NFeM2kNrCAmpcG46msQ3QrSHtd1lP7+fijrQvbA9pwOInnVt
fE35yDKMv2kKWkELDJ4B0xSwfGSNPTEEaUBZpixqqRdHP78KFQpI1797WoYNhrkv
ILzmqYZBolTPiHPPQew9OUhgVWSrMW5mzReRtJLKRSpOJ++2SEAC5FFoofZeUp6U
BE/fGTo17XZicMTFBpsDsyJIDmJBDG19I4Ynm+v8rE/dy3bbfTPOJhN5ue/MczMm
tsnVQHnazJcFYoWRwVauLSmkvRFSoFlKDTyizT1DHurJfM1QTNu8+GSl5LouEWXc
yWSzEHdEi2pgis9BT/RIGm5lWGZ0W7+psq7nZwJrOnRfoFc6da5FixI3rx7Bv8YI
04ZPOyy10Om0hy4sagxIPApdO8hMAYkLWuRSaI2kjsaJEwDlQVHQNSxfKK2oY+XK
OzMZmbz7kWuR/zu+pNuGq06vOxnpFXtEdNKqM0Y1yGN98VcqbjBpPp/F4qux5pVP
E07VX29tbtx7CP8VmCqvgc0YX5Q/lIuGoMxrMdUHwLxDRiwNP6Wtgm5wFtZRRjXD
R4z059Rvcb/Sn++AtYndnbTwbckbzbZ6srBPl2sC4jV6FX7ONgB+AXfJJ50/MpZq
XHojPjGoLASmBT1yuN99vYJHnkwBxmqSwR1495xCIzh40sVu0qXb0IqPtoruvdpH
lj+42Ewdf7E4Cz5vOotyJLgtPFS5SSpfoaBnydp4y4f1W1YrW4RWS8b9NcgoeRNe
BHg2S563Zn2NQM5gqKN5iZuWjW6muLQL2VlZG5e6PJ3XDoQzZC7rugS6QJ/JKxCa
+6XEZYP77EwbdH1ZfqyS5Y24dD30bmri6kud7hsQGT0u1+fsrcQsKEIcrgA1MjEB
x7ekuQJJ7yOjRRLg5/kabn5U+M7/pIi2pvFVUmWQRpSaJZMzwfD6MweTFWyDZpKg
4LIVjcnaQIg3MjMujzye/vb6XwMtO2qK4RqzSYR1ulYA8jmjbPKNIxRG3OQPPNkw
VDDlWcGfnzlS66xckNyWf/HOiQ+d1YNQCEXEYCL8xH8JZH4wMLBcmnSDBDSiUZ6F
xyTgWblTUSKEUMijVyJ9f11kLCSYG/Ho+pjAdK4XJwSb1n/f10G2wbVjsnWee5IZ
pdb2XEq58LgyG2divdXl/AUOQ0rAeePfl9cmGJiC5K1YHcn7aycFhysBncywQMa1
YBcT79cJy/huoPeCnMHeUilot/c8gQq8cHvusVWg7sYOdxabQDFH2vx1hjEKw550
Vo8CowohTETR9eglyUuzCy4JXv+zb9lrqq2ylCh3fMN1lsI6MI0ozipPI7khvSzk
wpQzjjFw07VXnpMz5iU1E6/J/Wl1dgMUIDAbF+D8CwBDck9EFhM8HhO77G15UcEj
vGgiVYeoSqeDIaiXoxgrzD0U0VdbQ4M3VWjRDJxPtTx7T19SGB9R+JzBVpNf0G4g
UszJ7wzQ1z1eADIZprmN1pGenqGCdNh2u3jq3hXdS7aip//lMACPkxZtGxlHtfse
Qh2Ef63NlaT5LMugbBrcP54dCzP+Bwxh+ox90UoL4S0NZwdCMmWqNNmNBjaNOO+F
n9bJcJ9iqmJjsMqZ9P7J5OSVZe5eldj938pnM2ug4ZwPddu0k2SxdZB8qEkasqur
psLsB4+CKxz0FudGScAVPk5qzD3kaSxzsHqhdm4y/AaS1LU7Cja155WLz/VJRmAM
n2q4sPPJNp75YkOyhCKA5lz3phQXXSm6o3u6d3RI3VsUZkR6pbYRE2z11bFKmfw3
pVZy68XZsizXG/Q6nE1R6XTn3kmDdjTc+ziAZCaKPKv1WO7PMd0PlZhFMohIOwjI
fbeFlqB0j+zNE+EvdCDwsB7FNksgOIQXoQXEZxL4XozOycsikejXQmXFIvNbOQmY
38ClaP3AYGZcdBnRcCUKKKBudmioZrekwMFBHMKRa8OCbvQeTizWAML1ekSRkM48
HZxnf1jRl4FQln30fOZruF0MRAU9fUhpADoxAI1CZQOxpfOOFOcRpEvanuCAyVeo
eJ1zYlEMw2nItelro2LS9wgmWVO0EZ0Csi31VOFTqi/oF+DgXyfj5+VnDnpFXjEV
+2DKEvzDKOi0RdT9EVqeueBb8decMDd3RJC/J5r3LlMDxiDSxYQKWmmkKkhHEWgH
eLzsxyzLIGZt2IynVM/37+3+c6xJw0oE5HJyyXot7T2Vv/nrZWuvUtB8YQ9sNlKZ
ll/bYlXMmLRHUT/Vot8LAXaZJe5zQnCJLbJnIIVetZT0uYGKtZcdR8O5/xAspaca
7vfY6NE68+jRn35p+8E7Lr935ONdms2KPYSHIvAeqrbxfbMZaWggdS32UagOCf/U
q6dW4z5jCPPB8PWaFk/OzO22MXaZmj++w/Au9Wr8x2L4HVWZMfWNfLs08V6l1cyt
wXIFRIHOqYyE/c1r304eovH5VWeFHyzoMQkuILbFn7MhI2XrO7n+u1PGJEHzODp3
wJfZF8rzx+2HIVnyGRPb6YHfb9BvpOQ4em7c2lWCKmQmX8KnObtyyDPHeoj7Qj7M
GKHX+akouKqEXdFsA4MyvoWj7G0JcAGXEV7J6V6HvV9XP8Kdn5GGfVvABxN2GejD
dJXrZO7sAZRy7eF9ZK+ZbhCvks1xra9Suhb3p23nL6iKZKifwrG8pUw/SxX0F7Xv
qM7l5oLKM5+IZI58PkMaBY40f+rQzMNAQu/aAb5CCSeveWBRS2iq16gNrY+7c+YB
T9DWokwXF5HuguhBsjLHcsDRhECFztJcLkpB7YREhRUMDOTDkjB2ah3pNjPgp4QF
VL0ZFU82l+rlWst+Ym9B95lD9JEMqe+acg2Ndy/UQXAFUDyifTl0ZtAxVxQMh8xk
8d9F2v5t/cy2ye3yAGZ8Sx2IB0BSAzjfeSXe49z9Vs3ZRfxrS9BpwqP4Sy9yp91B
dAu25/0WLADvvsXoOaDVm0IN2uUng4/+kGudRPowhWNdnzdZenfNyMpmNkzU8/TI
6DIfPi+8J8CnezN4RM4X3T9nUcmWBrjGRXH8PZgNn8swvRJmI2JxgMG/kALQTUMU
E7jqiDqii5sz3mDK/tbPVS26U5pKYroESuV4Ov0l5fVtlpxfoP9muC1q2ke2KTUI
ZvcuSL3a03AAktK4oTq7EJbotmyyz7xNHetpZLjGY9P7GUaHa6xHFIglqSPvJqMB
iC9HyPZpeT+sR/gZ/X9e4S/LVHdV2QNJbiF5AcT/j2+QdoJiVgVXF3Bi7dMUGq7I
2QXSIhaWINS3Skty1janB1/c+yos3GLmSmnMSZf6sdWGOVcgjH/4WUC4BuMduGng
ecIx0zt1SKhOysm0s46bYNTq6FlKn+f5j/xQib3tqfpXHXoEQs4nnKnHQ1yxRMrY
2sNGz4+CNmk+enUjSF4neTWd6xlXx+4fo4zbhH4ZaCNZqhEsEiRNNiM46nO7fzrr
TN6A5Km+vtN7ouWRYAJhjp4VPaUVJIREn/NtulyqXPOKyp4ae2wsRNgkPN/6Z860
YrekFJ2oqOgUpaN79AuFmYH2t0e/Fn5f7jumt27nWS8mSoeXAHwP9YI6hGqvHucx
D8XJ3A4NhSQFTRZGnnkq1TTUiblWkjNvLdH4qzYy3JcVtTpVMoj8vnXe4yXeANLd
bEi0R0Iu7Cz2HE+PZNW35YQcOQEG033xcW9M6IhfUN0Au248YXajY588LlaYOi38
OLvsvDxlvGwc/nV0gz62iRevD7NxiQ1J+UyFXORFuFJHQma6iYUIaLo9PDTz8Rc1
Z8V9qv/qk3cAjyKEHYaLyR5EmvSR2Zw8aYXbqrZLd/UwKzv+klg+ztjZVGPKa7zu
uw1L6liehHUONO5+iNqEQR09ggbLf6aKnt0GyfjIm9wFh4U1vtP8H3uGDpMLx3EX
/k12zwGqdQJZtAoTpk3s/FmxLttikra7aO697YaOehj10nSKNoZXOGyItFMNlnnr
DZs4OTXhYoNsQsjfT4SQ9MNOc61wpeQwqChNz1tMzzrgWwYWA5bdWFL9pztrt9FZ
9nVrrvFGxZXJX9Z5BIU8V3zOcFH4CapPVhP8moYOUBfCuhKvy6EZo+luuGD37Ome
TcZoI4AfxWeUr6s5jPp//x3OxsedM/Y3NoJ+FQu4uuZrWnXTeKtF8d8sA7fzdRfr
n0cEQAaXDFLFOV8vxCjK7Kp1ImeiH+aDN9JeVnRuUPPOmyyof8eIa294xE2HEYCe
Csp0KdkVYVINy+J0gEfZ8Nz7rTLhGj7BNRO+o/LlyfM2oZrXlY0EGo2CSLuj6j5k
FWebpRVoGJVD8IcfIbzX6dsymCTGMTVGIC47LPoupe2jwOGP7DCe//fFJTHYK5Q/
dJFdi7jFSPAxvJ7cr3/9BNTA02ctLIcUQT6OW6205yYKGtorTLoZcf6rI0p06I/A
qclJBDVMhlxXYdLgte2SCOPsVD9v8NEYBY5+I46H4UInAZdEdDrjYBaUR6TRXhdJ
lbD7Z6BrPm32tQ3apQX6KPA/AgzdHPl5m2CnIY2cBmrBunh2yAOP3Ykw0rJNBrib
2wPMl8vG9l3GDZa6WeVZaitYl+2oLCTKLk8XdmFtwc9psfr7gkWL0IugdoPHfw8X
YOyYRsl9QUbHyLuYYlFDmHIjAH0SI0N5uBVsSd8tXLGSI+WPSvn7kwh+A2hn/rKD
DuzXakdo18UZNmNIIg0MH9iLj0z7RipspDh3GiZ6/pFtNSUVog283ptWh7f0aIYA
AUn0MGNpBhaJJ1ojJ3KMMbQsx4A2liF5iVx0R5/ZOxncqhTRLmZwW/igd3odFjbe
9+Iz1h2NM9p/JIk9lUiJ6BOitW0fi3uAeZLZllmvZgmII0C1IqkIqZhk/Fc08VT3
4+H2Fnljhid9J7JDlL6e/DzEkjNeGgMo6xZGe8kmbv5uvpAxqLnbBj+LDWvYoQbM
p56fi2E64pRLwnKzTLTm620LQHU4ah85L24eX1XTETHXqqsy9ky5vNJISdbC7LjK
U8WYhX8MHuDIrmecofmbSdbxJNHZbzOCOTz3OG72XEecTafxC3z5OVEqvP21ZrY0
76uQ13K/BB3Xvr2sEnp/renBVP362RRmqMNkhCHL38gS7MeNkDaiYkMAQCWFhpAJ
OZ3xqhF+1S96E22JuX6anH5ylJUdtlFim5lDAaI+eKeXHavqOGaNQcTH2Rk0xQY7
NODCx2wOAuLuoL3gbfyenpjW/Mnk1aRVrI6lapvlmVf32wS8vmyDxCoYeVqAKdwn
55pxZyfQTReAR7hCgOauHRPa5sgZnnQJVAnJQa43CenzHcNchgyrFtDXgq3P9DcP
S9QGKQ/+mOjGCynUkDaCuJEHesQ9CQ9Rsot8221wMyWsqnUoud6KaVQpBo7FTADf
CtNeevenCIYSjiws1y3BTKCoBgljXDvrdNxRjgNP0t51t8y1ann+0ipF9gNByF3J
uLspuu6wvo1JfbIYuesL0kycPhACgJkTTeFh/FExGXCxvVALmUceGbZmUQz3PVaG
c+NdTERaEO0sPILYsc1ffxkf5HG+ic4nQgjNaRb66bkj4MkQaxzUinMP7zDxkJuW
9vSi5OTuMISS2t94kSkR4g6mIU+QCP7mdqMMO/s4sWesPs9KpTrWyfruSbo7inTv
CEBAUlno+KwEBROPVcbKaG1MvTJL1/yUaObZu0h7AVFYGNkhgm7eDWT1d6MBarep
EvXaYGhS1cAhPXiA5QNNAGABBoJ1jNSBX5EGI1T7pKbj0/czYca36I4H0w4GofIR
CrXBm54CcsbthJ5R0VVJTbF/n0NF8VB0bElqKuVCl+yLRQqLbvl+wMwCWshczg6W
Lt0l8La1Vr/vMEZ+0oVHRZYfBhWZK6SVPLBxWtjiVTlNcEiTM4V4664+IS0kJIOS
RgFLBdFKWzriVYGYAXiTS2vTBeuQP7dCUy/KDCthDRigArlLTcRpwFB4lhZ33n8m
VDulfCsgblvSK9iHTrh5ZQ6tKTkJKVaCuMdxTj9QZQbkBFoY1m6eZEDn627EY6Qw
+We1kQz7iB88HyoKb28MYiW4jryS2E3grFL7cMS0YmKJTVypRNfd/jpM0kaTaGo6
9oR8bP+5ohngd/8a/Y2OaSDjCIZ42+N/Sm0aSUiGBb4NpjgufCUsISSAY2LoZJ7Q
9Bquxw5/p6sZX/qGJ1oS/XgDUlp1tWzxeSywQ29RuO0lC1hCf0rdND+y76FgUwcq
6ffJeI+0fD4B3p6eZGDaqzBFsxutW+C+8vK9Y1VJCArhOc8WHDh5aDTse0tQDcfb
nq/iR/FcK/UaDPEV2iZX7+bUdqM5oiEzC/uo9BCDvNLf5CQPtrYQmQSIwfREUuZE
pmfuwpA+NHg1Xx0L9iq0M1C7UnYK9CBd1xG2Ciwqj3Qn10+4k0NhEZJPJvqcoRuC
O2olT8wHg5nSjh6B9sRQSZ/AnU3lFO6xEPC3S7dY1vH3lwnwaD1ov1bWlw1y++k/
GvBOCmKo9ghwd2wPVk6PE+8Ryq25R/X7DCmgpgCiicrBXZBIKivYmDOOhiC/3cFC
ySoq4TT5P/1cBkE/hKUfAXmaRvHL1MgngIxcKIOwCkmt8s/8ZrU8pPvsrjTuNqiJ
q+cdyBUxSkh6a+mkjMXqPJEANe8rZHeC7dmEus9a1wZXb5sJiraKup1Kl38ugg1F
WxViVFOIp4KagWFDbWIu/P/CdJU3VRRPiWRfDNiFZtMxscOZoAULcOTzxA8g5RKM
TTsSI/Vl6WHdMts2IijLsivVFvHDMFrAIsUXolaplOYrKvuSMLsmNS6gvqrmupQr
UZ3IslWK8FSQpR7b42A3yXa/FfZiv0zeSVtEE2U/DeKXyvv3xK4Df5ICdrMcDBi2
V+DhzJFnSxpRVH1SmL8ySGEqwAfsOeM2v35/J+ZB3lcucj7MTVGjZpDOySkSna0N
aqSGeD5Ql4JM71wlNYuBHO4ugayq4jhkSDdRcCb6pvOO8SIUHT3esdOqiC6cgP41
Oxh830VtW4QOoZkhuAY5fnkheUI29IrDTX4ZrL1qJnAqEe8EFhZZROjzASLuAC48
Y1HNruwfU1OmfUoK5G+dM+xyJ/ISG+DWmmCpyLLzpBMy41tgnXLhJRRFZllKlq6S
Y9pOYW9mqQKWkKEJPnM8LKFf7qPPO4+cwuxCKw8bNGLz3gkOdoUy/V8hFXqegyJM
Mpy8LpVkabTguuGcfsJxr8TyHIv+/nOsSWquv8mzgwnFVbMkcds01gvDio80j6k2
OOkO7o+WghapnF9qkEjujyC+Rxjvq5Q8NEEP92cbEPme2RpS5kyrHF2ybhqTqJhp
79GMV3JIY0W+DPt1ndWFKtLJIriubZd1mTZcf4qZpPFQjVxqUQSIHEsLlQY1epts
0LyN6/98XSHeGZKnJSUC9pwi1klm0l0LLYR+vP5DPDXBCRNdwgS9Uqapeeqylyhy
QdXaEKoN+1YE17UBLhg8BJdlj+HcMfZBqMnDBFVcrZVdR3qWQCFTFgA5LNwm6IXM
IZ7c4QpsXIfvaQkOkWbqdMXWRbrVSgVFe+IZZYqrBGEAANfDnZxNr7DbAhbfg5MQ
8XMHMYXcMDjA/gBHdsUKkmmDXu+hv8ak0NglzsbrzlVlmiPg8NsOFhd3GUNxpxTN
rDIfyD5oC4dEoHWyeLubfTlwwfxnExUJaY+a3DNrb4B/SgXJmhWEcmwMiFpBF76n
+KpcPEkdebsXi9VVghyTpC9dYFsolGjoK7BIWY9nyLl//ktgu4/uWVHvZDbUkYJY
6wiY6pUnd0s1CAYCeQfKGiSG1oxo0HCc0DkMJOeJsqKy0mjBJglnX0awhVeoJNYZ
a9ZZiNhjN1ZgA0IeswBVZEd0pboOrW+mID9CAYa5ThhKe+pZxbTGeSqdIx+crCeF
u+ZVfvg8HG4Q5B9n7Uu3Etq++liJR4itiV1CPI8ADXazztmpmV6XbC7WQZTVeJcv
+QgR/N5BVk/35MxeLT8q/THVAtuAz2iMqRega3Y04AtPUAla4AswTVKFfyEIzdI0
mpM+WxlmKM9LsfMs9EfIHLMM02GysxnnS9tip538oLMrqJB9d5n2o5zFc5CJu8GS
t6iOid70fTrdo4o12Ee7e+e9ZzZCAPsaVB767GEF9B9uS/JoQtm6nPYAV74YQMSl
jtXnyDPU6wxyvVTcDkhwfvEqJXAm0Nd5Rc/vwerJte9DV3b9EH1F/Uwm6hG388ol
s06VxKGNT96XkKtAWyXnyQemkRBR7a7NpNHJoyCKNoPHcinjDMQ5lZ4symF+JROs
fAyjnJ+iaz2O0dpOUoNts6+wMPXlQ1gEK8SAIDF0h3rhGcY/CQ/IIUN+EVFMD2x5
df1aj9Lzpxeq0Yikdr1mybrOUCu0nMA542Sh+t/3yi5mCv/AZqWNpH/RqAk1CgVw
+EJe5by22uk0MW7f1YVD48sXUzC7EW/FfnhNRT9mFH4cQm9rF3Q/SdwmoE3tApZ2
koKTeBuAK1ajdJdDpvEc2FAlDz/RGrT+iWfxwmS6fxhUhcs488vxlsGPz20QF+Vf
h5Rpt6grXMW2Mi6KBGivDkSdcZ061iiCHumww9m7Ck3uWEqGiToIAvSnueVVOXpF
gk/yFVjiWRUOnAHIypaVwoqx3gk2nwvQEAdjb54gRRRwSTxBT/SPtmnppMYqSYZ5
YENsNdg+39GbstsSNH14Q+6hK2PDh10rwzmKaTPwSikJ9+VcuCLd+sKktNCrv0PY
MV/it/o24gxRS0lGs43Ra6+yDUc9cAyfS9jg3lU0YSS/wg6nggWuJDpPoC0isOfk
RcRsT9j8/KlJ2bNf7aXQ5pQinl6cWgV3+ZJp7+OYymRPIY6AMR+RYUamRsCA4EF/
KmDK+9Xozil/6xC1vOCsSDAZL42QcUSuX0OCYyrzZVvmpK/9jovonRWhEkp2NtP0
/gS7lZeaXTCla6g7JPxHMzgIrY2tmO7nOlmKz8avgnZRARUt8b3vHm/v4+wHj4O4
0KY94hlaJhnP5zkqjH5wxBsC1t6gmatPrcxhw6gptyLr3QRV7cyKnbCl3Jlzf7ce
PEVvj/3oEF2iLXRH7b50LOctFyC2oJUjt2z1IuGRGqf3WLJ+rtwEa759Zv9jSiZ4
E3yvmKexxSFbmZAbqy9Dy4avWzyFF4a/5jlLTpc9AhxTfWgqUISDPNEukjR+gQPA
KClGH6cM2B/hDgSz/du/nQS1fjnY6duugEj15KlC+xpKp79oa/JY//lMKNt41oIl
bGb85LXD0ohuiebWWk6ldMRrhxlxomPMplwpwIdWNpopwXyZ4Hg/sph7g4Tm8xAs
lycDHpqEZJ35hWsCO+05rcbuPEbTvkjKImzW0rh51C4KkBXG0Odl6scIWGb4QM8E
uj70x/8Lm/906iLHI9e6kVC6vWzH3IflihebFkqPdyUuJywFOW8rVQIlNQ4BXYXZ
fPHkRrJfXvnc59sKNi1x3AnOXtN9nNGoW1KAq9Ude1qrxsw4D7/daJaHmxjiQrdd
X68HOiKu6y9+jMlKsCbwyaeUUWZW/pMV4Qo+Tmlp0p9Epcw81e86xL55WKYloAoh
7BAcMxzx+e467kViMb6rzR223+8r2xQRP3a/8wuTzlrTr7FrycuAPgoo7QHdRQ/R
rGpI2VrGlPI0FXOnCNO5EBVvAMBe2sbs9O/s18+/3vKMwlNXIG71f72dsgurFt8D
4U6u46HsKa5blLfu+QEIvelGErpALumSEXAk8GszNW7ssUI+tAQPzhRS7JsZ6g0L
orfY5ZdwBHGe43bUGDRv8ZxU7TaAjsNgTrBub8QrNJpEpv73GY0M+aHNGLheoREA
b4K71CS69Pe4MMdqLYnz5cAxS7dhzLSdgM+2B4aGDcR43+4qs7IGPYkZR4Uipbz4
qpQ1cG74qF2vPaw1O/FC6LWtYwANSuH7uovdh034Tpk8OjGkQkdAf3N42SSn2GLb
k39BVZOHkmr4vnmE5p1M9EKDiSKqAfam6D4AAKncP1acA6p8SC4RVL5dsivMUGSO
n37JNzkWUd6lA+aLCU+LC2QFsYe0XBnHGKiCrXwlAVhxYFmTdpWHp2EwPtHTwfgg
JAV7zUVUqs9zxOSWfR3hNMktZ8EirBf2UPXiRfd+qMHU1q3MUYKVG9xipp4B3qtn
w2+PKPXUD/GXsw2zOc9Ha5K7m9C5AoAS7hcuTmtLlCs7HyiQ03lpjW//Ol06Zske
Be0KZXwJnYb4eYmirrxHVjAKCSmQM/vt7tWg+IUPc8tMwIAk5qCb6lkXHlo/QY6A
GZ1DqxyF333Y4Sq67kw22xaYs59ikQ+RckJrkm0JxxfdR3CAJc4BZqSvuu1a8IMY
+3XJgjXBur3qbuF2E2OShOnUwcEJhftT24DqDogVAFAUTDoe0E53nE0thUWVSpTm
paDJhyivLz+3Eg0bVki1tbuJRpfY7KfKvka7aZOPXuqRZz0bJPEwDZbZFbSLQHUu
Riy+ilUPO42ikzv4gL/bQjDCavsOXPss9WbzoMUPPzbEcS1PXRBMOv7J/qfkYMwM
t/ZjrxXXpKmb+O4p/mIgoRad9+GcMzZ63mkpQKdTWviJecGESfHrSWpIG+ZQKu5x
6pj6IrRGsT9C+crnqxsl8obhMSzJn4kONrLJnZxGGWf353D3923yl8ZqkrQDDr+x
e85jrGf6GNDc6pUQz6J77hZIcl7oIX3b+kvl90Rf/tXHnbBfyZTk1fTm+tcvu4yL
gox/v1BACKURW6jHBfncNxa/OuEIfUPvE0UqAsaSyY3cFGO8EW2tGYPhSR4MRhka
jTERb/EB20jwtXZrYj5EzEvdmzsDZn4OubnoHl7UYwNx3HhGaN9dnDEHCnG2rofe
9xQdqSYtPfW6bJrDIESRmuooDUWFRmNwnWWxPPDFecgJjmsN1YGb7qECyXbRnua7
ETC26RiUvGFEcBqOs4ocMEsYwMDNAsIFDCsPrBPPpF6ExbzqhbLN/lpEyC84zZMg
MMnrV1BHDz9V316HYg+qg7WX1lIyn8W6WOCyJCdKYUddj8OwvjCKYqYVBUQGUfcP
l+po1Ql9lE4Xg2DBj7XfRKuFLU73/1ktsY+CKyymQjS+YGFf/fzjLnOxHpmNsi3f
89ulnt60AtTITM3MTtYvwK/aUlWxnDwcCyh4q+t/OpdQIBtkK42zACGLWcgMsvtT
4QrcFAn4bGY3pCepD4zaFOb5TavjKsYH3enARXfnNl5F9NlY2lJiTecf8BQFObDF
QFmbQCjv5dyzOhbAYVcdRXskR6JVtdeGdRsya9l2ihQ7riWa6QL73IO4TmGKSTeA
eLwYhTVx3sD+wvmz5elfISEGl0uD4KbmHPDGuLuB9WFKm33KIzT0IWZ/ukTYHT/U
KdmQaINzWSKCFqSLtOQNBf1DrnypXbgOyFV0x8fdPCe+7gW3ZvpGsYwCzRqtwNKb
n+QEab1rK8mGLd/dZIq36IZj0B7J2em5u/BTyfbx6pug/6fP/7XX45q4tk1NWEKe
JLSmGA5/u8bQ9M7MI3dF7B+mDQfD34q5PcDKEonDmlQmp1MsW6e+MVN2ZsNg+Y/X
Dbb+zqOt+Ui+/BfzLcM8mRG46zGrSEav6UlYRz6D2BcCUhtx5wc/8Hhbq6wz4s4b
E065278cUlEtp5KuPyO9c887MpCoiSuf8ya4PPo8DR37X6lli3S2Hu1aHywc/Yfk
x0TRdrHb/81Y4b/sZJLtOvhyzgLJQ/WHTnG6ijOag9thlb4LehkGxVe1XHXgw6zV
NwC/c+uVu3wvIumymRWvsXdnuUITOyEH6u9N4Z+i9RkoAKT38VvzryHbuk6IIaK4
+4GIZ4+mn9EPmRE+nSrg33DuAglNHvmlzqigqm7f++TpyqExH1ON3lDekSH3Eam6
NnCLCuwEIey3O2xZhQDTZ7W4D5Yupx2Sc0Gmk79Qn+soam4u+Bcax9d8QGp1yiHz
LC2S1tAdRUZMHCeM5sYcvlmbdsMAUi5rjy5wX8MRq/dU5VjmLJ8ykInPqYyZM5HK
OYbD3PpwmUQVGnNegleEoGr0jlNgUtQQfB3wutR28DcLmELZADsuVf5FK7JTiA74
FfVScfnZmCWZB71kqYzIYQpGpTTng4pvjQq4JETHFdIqcYZF3ZDjrhxPQNgG07ud
jXvpB2uwrJeonJS8i6umXRRSDAVVpNI3xcCK7V3hfEAEpouDGoqwVqGlILx72f5N
SQnL5Tp17lKNoz+kkiTcZgj31+yOU+4V4vcQtAIl1iWy3DzyxkNndjUjZ0+0krK3
+RlGTpItSJtjYko2EAI8omhO8Pt9B+aACCU3ij12hsEuQx6g0g8dQ/INJV32yoxF
Jkv3JU2/ap4us9y/B3f6vNx6Yu7Yc3Yn+V0iREfIMBenIzRgHNralhZzGC/05IsO
6MIZ/DmlTCRPGoDPxZGP+OPPF5uCaUWNicmm2E8EQsM5Ku7IBFwIMTW/L1fOhKI4
+LFi62zs2owU4gvRRWt5J7muyNgiDwjYR96cCsd2PTSnfjqunHr2LrUKy9o1SZmF
K22E5lIul5UqQBtkY1LYMUdsLb/3T0NBJYwO+Zge2BsDbzjq0SuAWVMLk4wUG7Is
ylyJTKdoQ0pv/djqE/2cinDNz855E4B+ZkBIyWCU0D3A9Csn5ScOl2CS5QOdA5l9
PWkicLzpjNEo7sfx9ygcM1L8jqWRdiYtUX3NA3aXnMX0HlXgF4JTg9hsgJVMkkNd
5f7flV8BuqOtiQlUQ249H/fRLRFJ09UdNBlbdnX9eT1AgAAjxu6ARLJaezdOgtuf
TsBG39/n6BgnSquFzSiqDWd1rXVUNquAQZXU54achdA+uXNCnWVJJtki9Z3eLwYV
c558p0/n/Hj53OWTrxJH2PWnyhQy+xEqDSA5DDgE7TGifdZ3g1nsYtd3UsoE72BV
WgVV/tZbhRmbsjYESKTUETwC+/iIfK5T1uZ6T4iC80jof+lL74AoLOr30JojpGwx
SM0nlyW6cZOicTLx2KQ5DZ7IpjMkHayjEgbcGricOzZm+9DhynAZuXpGjisj2TXs
Zkk3IGMmOASnATgWjLA/OK1VIx2CeYEi4yV6DbWNEkeOc5HZ2vBIxzAury51xmi+
Z/7jHoVJNS6EpXVzZERrD7H1gfdXcjpECnY/6NsW//HEv+u+gGAeUcvTLu5Y9f+3
wpKaDnm9u24+4S4fxoNrlodbakf7z7i84RCVMkOGAEIeTFroiUecz3OCfHPEQnBh
qIw5HI8jWW1+vJFBtwXmKAoiud2fOLgN0/nQ37J6g92JJvWYSz9Ctdd2Jmx5AflR
9rBPMw7h55Oj7Z5fqnonnTSW95Jwxwnxj5E1OaUTFvpeLGe6eqxj4ITJ9EBZbJuR
HetBPpTSgVkIAu+zXPjzs6kD5JkD4B2d43tRYXV8tJ1xHeUhAJV57Zlj4B977Brj
ofBviQDK6V9NmitdTEdn18iwPiQOSx5IBlTieQnxWxHJY87Nv3X2MnZqYyKGJI3/
vO0wLKwSZmdft7ttOAwJc8HzliDaVCc1tdpMMJtbiwkAqw+0Mu2NO1dCGtqp4Cxh
fa2gnTgnQGJSRLBz7Ei85Gnk9Yj0sCIQdXuO4E85RXpXNbNJLvBGZJ+SXTkAsHhD
UMvMD8SLTkSsX2IFr5teUgCLyKm+UoE90swPXyh2CG5naPeSfCMbUWb8JU9I1Sia
Qmh0WYk/bK2/QaL26LKW5/QO9K9Hm803TYJlHzvtjItUeZEdIDN3e25OPMdnKSz8
f/bosX5uzopMhsMx5Zchdcrh77E9PUkdjacsLtnT3VjTF3/YyddmEnkVhY/xI7cS
tBy1DSYCoooBFM1aS4G4E3k+kO9ifD3epThA5gRfeV0B6U/FzbsOteLqPQZHQVjD
3DjV/92vJfLz9/iuc5bS4LvS0NVzr0je3+0Cbd6aOSIhjzJw9nqFPpguD21XPnQZ
VVeQI7MhfZYKhaMPlz34+8XEUDmUtMsdw2EUR68uhpnCBTYCZdZSTOGRafGcWGrT
qYnN32zghLt5vyjr0DADqVLGDUwYyz52+KLbX1/mUeEEvMnQDmZY9gkEi20wdBDm
RzZrIgt/tLvCDY8lxrd/WMNFS5NCZoXc7X8hiXdNtHeb3Kc9QlCnRQony8rgb8sv
YTRQ4hGJvILtzbjwgPKAueZanZLYugZxYdklqchGeqqANMIAuAcW+i8qhCXBStSn
NsPhjXyAACOUwlyYoNRJXQwoI6KUFqT2qNOZEmI12jBTM9BCnXYpIq5To9wguXxE
jXZwrLgzBt5FqHSgktHesxUHwwZowpKLFR1nNzF7Ju9q5W3dVBPqkpnLaYfTTVl8
zTZYj3n7V4gW//wLIlOGGRqWmX1UL2xo6QH9uB8WUzTUiZBTVVoSg8UfRIfXSvAA
YQuO3mGqV7IvGcOLY4esFo2AZD1kdRAqPEQ1tFP6CWCgNcjMJd6fCkugB7XzBlEd
3KYFY6qIwyjtvkt5S6ZxwDan6p1HeTHn980BS+YiTSVNoOkUXPj+77tjz/1Bbn89
H45FG6zQlanFdAlEV5iY/kH2UewoY6cUaPQ0lYef2piRZf+fwXEaQpTPqwemi6Y5
WJlKhVx7A/6FU1K40Dx3us0Yqgj9mKyPwrBg1eHq1XkSTOqmYcYGT3MVj/md1cBp
9pQxyrG68l3wcZYLx9SFAB9XNoW/fJKzRdrtcv3g+tXvMe058ClWS6wOMUn4Jqsf
fyjTMfIBxoFwSE9YDYh/nt1L58BBXS1jQi2hE4+JxYAWuM65MYzCDc6yltZCiPfY
NzyivNpIL7ghMsAP/b/ORDR15+6DflksfLrDmwZaxY9JH0SCIcP78uD6JLFOw+Wy
CDEjZ/gJsY5yDaCLYGrlnNjQwr0rj4+H0lpmT/tZ1h+mJVrpbff0XhkAJRLdX5jQ
cvmWcwNQM3XntBIB3iuO4fcABSFu8GqIodxfNs4czNK7hIfLR3AljA0TeD8C36Vm
AvgIdKz76cDZYLQ6TwoDalNQouEX3q9A7ZJ9gTBme7GuPyxamzdsngOjxCR1YORU
gF6XP12/aPX3UahR+yi9pAtwz6y7H7v9HI+90r6Lqj4Vsc9TkooXRhIfagn4BK/f
jVdtIr5q1nCgFa/fJwMD8WIAdkM+I07VyhS3+xpJphP2+Du7xO2M2X70RW4SLJKP
bpuT3k8SduX73SOP3zVCl1zDjDa98umtAIR5MdiAAv4Dk1TYBkDPI7naft9xUECl
t/P+x+O0xEvmFcdyWarD6yBHMIT9ByuQQLJIZrdHUT2z6TxatBtrR+QHMf3bv/5i
sO91wL29/QpN+vaoFU0UsceGDqUXj/TBsj0ahQW6792aQDfGRwZSU0WyeBM9Ffz7
hSxPmHGRirZhxbQHRs3DFKV2JL+OotXhmyfTGkYutN91u0OCfWJV3/gFlOGUq5GW
Eah7rVfRQA+TsTldkIAuH98lRQMU5G7NhKx5yAHhkskYnCes1XZ+6ua/NqkMKumv
dzId4WrYddo/Dq01blz35vBZy6jpMqdn9Q+8HFxsVYQe/YnAx727MVayKl1RSYVs
lv9+Q2d6rGFNVi69gZSbRexEAr5ZaTuZsVcIh6QXhn2KShYiwSgWl5FCNrCSZvvQ
rgZo2uh5IeIndLBMTzuJYA8VyipaJAiLyQRXPXv/sjl2kgy++CUazjI6GGsplHpS
DNa3QZiSRzUoowq6okB2AmtvC1duv5aO+tZYUBJYSqZWntlHV/6Gmz5gBuwMezBI
8WBxjwnXuQZeSoimxaNPxnFspBC5xh1twavnDkl41n/TKkxkrBMi4+OJ38d0gZ9z
XKpsKH25XXntYgLUyHV3RpVSsfch1qnS4uWF5Va3F+SL6cuKh4tH+LTKg8scp3JY
DuZC5t46BBFDv7LkU9PLT2JUylWcT4D3eG1Y7uppp6ehomxqWRgFu57w1sSmXt6m
GZ+dnJnPaZeUjDa8vSGsiMvA7jz4+OgwmBDxwnVxfhhovcfhSN+RvR6/Jv4wSvWU
tSmSLZ3v3kH7j1W98AHjUQnheoy+/SkKlRu5GwyGQebjKx89ejPxBnxFU66Dt9Pc
4JqIMXUxkSu9Qur2krPj692PhVLmlFrmTMlGWJbsXgH5fYz4s4B4yZANY60n3N2a
cgRQP6hqBc1Qw8UYbERLg3TwPqJqXuh01bh8giDRwj9YLW+oWGtgv6QZmZskxXzb
zPw8KMLeY8fOHeEhMHTh9u/gt31TgazTK3yuaOHIaRpb44chHwzOxodFnadwJq8l
ZxuoGeKDuYcyGqDzpb+XL/EpoUbM5IImxby6TOx/GvoRt82daIbSECK1t58+WU/I
6VBzjbdnGjlOtvUDAKkCODz2uanAOsci5bvHzknP58q6TNE9gmLZ74xYCB47KVQt
OFumHZF+0k8vVTYNs/Y+kBplfoGM5k+SerzdTOez9L1lINAJcQTOofIeDCzSV4Be
dYNeYTtMyQjxJfPSfFMOVNkucVzftJeffmBYuBDTFd/zBoyktXaWh6axziM5OQfF
Q1DvJcwSb3B/FbsgZIMTdEKBbP98mWq9uL+Vnbt5nZEKLnrhYSlXbjqLmkVK0PMw
LUwbg/4XZMeKL2xYv7JyefzOtpgIwlkx6gX61phVytv9jDaBfiL19yD2Yu0wWEb+
A3RYUOUv1cHGNZ1BKQR2tpO+QS7/Doy15to7m9P5jUnfoFyfoNOoLMD/o4fnteDG
DkI3SguOfSvWFob9hG/W+P6/t7E/f4qFqWuSL9aaoQuxCHFNvcUK7QoXyjwu0n0A
TUu3TvFyR1KXGhnVlwHhrQgQjblpx9DhEQelFWF1k+o75F3EITBrVwVaihLx3feh
tc4RoylY9Mxv+3hsHJb0bdG1LEggxMc+eCfc4bf0rbYqDYi0LKxDNWCcUbDo5Ans
frFDk0i17rOjL2jzVi7AFWYq8W4MMknWz6CBMgLbbN8AIdjVam4h9O45DCdq/ttB
LRHAMRBpQCqgO7HaQhM6lX4LgDpywc4ns3WfFbtlUbVBsjqwszUqgMo/+D+zKtmQ
8tGL9qiEdkmcFgCr0uVjXzIUXTPq5QHYyzVB5H/RPFC23pDeW5O0xRg5em1fiX4C
UbRGN/VkYWNEIo45jv7pdIuoMfW6OKHjGqtqnE90oAiROUQYFaQj68ZlFNohIeqR
VOQHMIdKzypFWThqZqog8IUhN54HNGbUUeVBnrJKJKkWQFyKo4HcUyaCZWIg3Puq
AHnod1ZR79bbcy6acvDL7X3jsRCf40e8nn/JcLyWEUg1Vz3l0X73Echw0kabF2Oq
UChZXmZ5b6YELU4YnjFfphMCgLRbvlOnEgWS9zS52U3BC52tjrLDtmGJEPoKYM4+
dS8SC14jefUtIsfGdrwobUh8nBQG3IFIh5cRpamw2Np3nhpgt2xlNYmGnAV83xtz
Of0u2N68nUPK1Vb4o/d5TRuf0pmH4aN7hDMl+GH7fx6uiXeDjajfa0lWoDEhW30j
xTI/iPPXXY2U+Juv74sBZzGxUalFHt1QXLUUgkakqtyy6NU+6WRvF4wGCVDh9Azb
RTrZX3/P1kkBGfOzMrggY/xryxLsydeaASmr5mylm1nK4HTv0/YHch4VV9Vw/ARY
I0EUk64dVYhP1tGIV2ag8cH07yWU9z4ipsjN5SMN0GeR1cXA6TcDj3qRUDCAKOMz
xLHdONNdf6urf3sT2buaWpnQYwqpTVjYLmaQ7CzzwwcDWLYPd6LEXdA8fjE6WNvp
I6zgQqx98mE2H0mYNQW7x6xKjOG6+pa2xhH/L0SiJ7EYI4+3AYyWz3hZrHZysbkT
sCSywmc9jhW2FQr6JwLGsYscw/hcs741EWByQbRpINetL6adYEnY42xMi1/+BpmP
do9+v410rR62VA+iqsu7TOm3cPeCp3vdzJcrOQJb36L3/jTGo7IGPrUGRf3GGEaS
Wxpx54UmPa5IhT6pvRkh0nrYM3YB+JuPelNRqfv7jnoXM4x+d4TIu3z6vAhmc2ba
JN54T40u02MMKwX+DaamCCWpJN9E5GRkxCyLbzCiD5qSJIh52VK9KET6nT7yk/JI
KAU9Y6d5s3silnOFRU6SKQfRaf7KJp0RmgG1nt/nXt4Id12aC+l3yWhttiyVUuNl
g1Y84j400WBekfLunu6SGiNXsA6mrKSUE5rL9Eh1ecqOdmXwyRDe1BOyl2F1PmMM
4Z8d+MARFtFgQadQl2k0fYiXq0rJXsPp39cgmUwVOhmFrLxZW9tRk0k0iKlzxwyQ
qR22G89Dfhv1vmPBbnyMXn/RXIse+r5rIXvuyl0yAvfSiEuZgwZc/P59vTwShwJY
uxPsRSm9rK9aun2F//3EVqyWwB/fLmG18UUi348+jLTE48nCIkVVza0je3Xy6Gx3
HNkl3ldnsH1ijx5MUKNArXiYlrPoHb8elg7ywslhhR6huVrVgH/TCtljDBxR56xo
Eoa6s4g5FcmhbgC+HF9fa8oYtbhjp5mGWlUpE3ll3C0mszuuxS0u8tBWYNRbBFPE
yGTGT/1uG3qmPjf+BapkGunJYE+RpV3L9pkyj99nyqiq08Ap//b5cFMlc9Cd/0Ev
lFNTtaMxMVh10nct9TtvyF6nwQKfyOyRkqzt9lqWHhf4zLD/Ov4DOm9xNf0nbc1c
WGZr6j36tHZ5G3jDVsABdOXn/xxmAwNRmE14o0+NlcSAm0EI+4sLv1VC9I2+oG80
A7BFSSFNAddbq1bsFvOKW1+7BQGdbDfMQedjB50weqA4PlPyyQ8+NT+yT0hkHNd0
gYajjxXBfV2QxrpOvp9B37VM+bOS+xZscmz2dhLTNy5uj077xHxgv9kRZXeFU6sg
PXaeCjiLJwOAO/AF5iyPPyKnytb07m/zKe47ONYiUzlkGW1ZqDAgL5aQfJfg/iH2
6uWxeFSZcxfJ5HA70Feqvb7lgKdfwLTshrx7y06s6iwF3B9FNM5a+AFZkKWGzm5l
czKI30cgUlY8kFWKJ3eMi4XVnGH3lphsgBISn1BvWMNH9Ea3ZWqHBquFsFHsWta8
ybV2EWI5BtP7WNalgbNBTFkkBXvkETuW9+a9EyK/nk60sJKBVQsCA9Bn2yB6CxDh
7PlPxQtbtj+6cwhnbx4+Vp0oR84QCLKsYJCBEjUB+HXGvL5OK35HiFkg7qfqHoS7
WSPSN+DcN3vilQHVhL3DC4K0M2c2fJb9CMG+XN5VY3wOOecE8PECOzi71gX4PoDX
gSIcxO3dlPgn6X2UkV9C4CiNp6Vn5WwP47BnMDs+tapkBjlf1NSC1QsBcYJG05kt
y593iR5AlDGL4G0KHF4s+BIPr2lBCj11YPdEoTbdtEhDlPg3f1F+u3UxoAV/JEfk
ADlhkQ6BnMZofQndNfvJYeGbk7Ot5UlbubLH5i79Hvx7OfKE3mNq4OzZQ5F0t4kL
yCECKRxAB4RvdPHzDQdiCVrnpd5G1ic+LS0LEnCkudMts56YZu+ZtrwhzMeYPESl
mVV3jFOB9XBLBeMwJ8xLKSIcUbguG8cPF3/TZuTFIsDjBtXhY30vrFAiWzHObqwW
buFk9ui4kDFN8VJT7EDvg5t/OuWI9ZH0QUuqecCHLd+JZQtbElbxnCuBBb2oCL+X
KLrurYQCDKETHmw9B0RrUyZlK9rVKhOlnxhz/g+qGB+dicIThf5Ort09vVALnKEv
Nl+pGL+lApLTFmqbGOx0dQSy3LpB3O5NJqC73TYao7GoTL5KHAXzc6Hz+6WtW8nT
t2CVh2ymwzT96TNCW9l32IGBc+OcNQGTedQNqCLrpJplv0wLMV5BPO40GioGsFAQ
+GS+VCItM2U9VAu5FAq5amLs0q9JhZDBkPp6+Fu3wz6dWzRF4B/KmiDJ97OANBqh
Y7ryyzsV8llCu2gEWsT8emI46d4VGAb+hwPBKK7KeCrZmkW5w6gYsfmxEcWDO7VB
AWoaQdzVzMmcE8Yz4VBJq+2RunYwm/BeQeChUJMH1oFtg+20VAueJSdQo94qsl7Y
RBegtUe9IkREEHlK9G0TZ/dCYcWy+kFK0WHlm7Ku+tZmLJys6z/wFVAF69/utKTM
1xD4TBwPc/Qq80ex3P0tfGUxa/2cTTS6ETbnIgD+UP07r7AtY5nRoDppsxhueunH
7KPlwxqv2fsGS6IATGDzYoQ1bCDxYhey60Km17+s3URjR8EOWpNnT2JCVSjJMPsI
3T3QVHFzfhjv58Q0NDvbiZT5UzvWUFUVBesrqsSMw4rNbyjNpAGzJmeYJoXb04ec
IABTHSRS89e/CNrmOk/K+TnuQH6/I03Ski0QvfG4eszd/Zo1JMVdBK+VUA0WYDvs
y9hKufa9PYkD3HUcT/AyuXF17AJkYpxBhSIa7y6SY18eoG/6Rjce0C/3th8r7uVf
44AoMcIP9R619lMCv9T0MDFSlHCUb58yiSIPzMVUNzVAZK7aBJ29UElQ+xEho0dQ
TWmKLiXC390l+YCXsR9/L8Gw8s58cXfOPHsScooFHoCuGROdfJqskcw250Ahb4i8
40d51oVhwKuLkxXo54fM91ewoq8JLZB9MlFbDtlsxzqLa1UUIMnvOgZEKS8Njxis
PliPqS8apslIIHwZ4gYSlE1+JhVh/43hyUyCyBKOwKxECLhuF+8yV9i1UGrVW180
gj6Mabs7SfW+K/tdSkJTBMViFQcn+ELiZmExW6bEpEHB3/YS5MIbfeLbVtzOhD7Y
iI+7wdO4+pU8I35Le62jLa3F2hr42nAzhSmtzwZDxk7tWuFGnNx9Tr7k6fTzdkW+
zGSB0JihJk+QQ3VKab/oabUnIvKqjVUz6kpgnMG4VGNVSpWPwOG4B8zDSNAC/mY5
DsPSSVkOh/tOUzvjhe8E7f7W2M9nw4LNi+03qpUp3/f471OvVjm+XaRDOHPlH2IK
EzUa7qqxmZubIKrwhMqllWr9v+A/Bz3lW19xjNiiD7Kqxp8VDp4mS2FynZezzAx8
VFjXZgjWBOSAHI+yxl5t5DevpwinSTTYudlfTQeLVEM7KGgW+2mfh67Vt4wKKBiM
oElm5DhXGQwVsDm8V4Vky/JXiMfK28KMUCwUUwT0Ig/8ZeOgHk78pk8Pk517kAyB
DXczgzG6TOzEedQJxsKSzA+1wynDM8wQauj58eDRKbBywE9Zlr2ceeA9VL53+K6X
wSjcT6NtIS6RA8U0NDivizWF91ftyb/6xDnxN8x0Qo6/BChJ46aV/zdjz/Y7rG2B
Kmi9VqVWY1dm+WK3j+rSYWk5NXRacPQHHl4GvUCCZsf+4kMdNgeASWVGPgjxycKu
6RkzaPNlUkuOKxyyPva43c+tYBgIadaCj9ca9AB39XdtVg+RGijhzhOE9ttCqnFh
oXa8/93VAoy9BKN39gBPJ/94Zzeac3UsNwqsFIOUVUEakAdg6bcvHfCws/j5xPf4
OFCoO06ql0SFP1e6sYxfhwx2q4xe5DDocVPd5OYrJov+EDCo+MujWMUGNmCTPjtw
K8JkEZci0r1elislAYTwtv3xK1jdK4aGCpvzadkeQkqEOwqhhicZEs5O5pIx347q
eYzhi+9LsVHPprEPNSsjxJdRu8DigX1f6YInZaJo0YxDIkUgoat/t8EP/EjHUaTh
mwEuZD66HG2MULPQhA4andsFwxsaRs2hTN0rauAJ1G6fdDyKA7JB90+x6S4byVxj
0URRHRusmZ18bXXzjSxKGGnyQXWwi1/xzVPotJlfgTPqocpLQ5cv6hOAEmvmcOFt
UY9sqlCFp0r5sJ/RaUJZF1noUymAKHfw8lD1EL5EBwQKI8A6TlmJnOGASUHGnO5Y
vZ9vV4eijF0eUF+aUjfyE4PpfQ8zUp9Yc8YaVJoEtnCt/lQkP62xjxP/T3YgrYHP
HecdH+GLPdYx0+Xywt2BW4SiVDZmhQz7jeLRm81Y0RkYqEs6aOjBv5X65Q3bquTN
pm6GxkUYaY9Hu+Gx4r3Y+XF8zyl5f+VU23OHAfVHZLBku02g4GaLQLGNhbHjH7CN
63OUXTSwa6I/IP8jWOYiZdFwmqiDkotKpT2XwL3/QcKu01tilCTdHY5ptcPMNJ1H
apl+JJfoBVt5OG92YDYJgUyzQtm3f0MBv3vheqSAz5QvGUZTs3lnGEc8nudk9lDA
Hf7635Ued4uZNnQJOwPy4CQPu7kX3u5huk+3PwgDQoLCKiv1IacyMrOhFci9u6VW
6HtGt5rz8b3GRVW4yCf0uTWMxXzjXRAQzFVniYfg3kzYIaN+uuC+2PjgxNy3yBLv
Hrj+GYirQmeQNj+9NOlIGAJ3UJufyiFboi1Hk6eV9tcaF5da8AP8D24ArCJvTTQj
XKfWHWy6dUhPwOo7/LgsDJ3qyMl8Ofe9vO10LutleLpAH+uo3OhNkyzscDaC3TDy
vDqkv3dy320AEunwoEluIPVj6VnYWjZlG+JIW2CjFFgimtdJN5sy3R+qT5JTRtm3
dIwUyNIJ7fRythxOYGFH5ZQBf7r/O4xAy3Tx7E7nLqqrPKX8Ua1vlyu9cZD08UzT
Y/KW3xpy4UML6MRDo42icBBpCfaxC/Uj8n3zKOV4KB6aQzqWx/bPkZ4yNz24jhV6
GmYsem39a/mA+76/vXTXdhrcyQcTsiHpP1s2i8EsNfGoV5gl6CR+4mfWk++fXqrn
aIhg2y2kBUhDrT0YzF92/sR/GlcZgp5GMM2gLrpO66a1rfG5FjES8UvdOYpBA8Xt
NVGpTh5kOV/z8N5eSDfcBuA8ivTOKTc1v5tsVIWDD1JK6ULAbSzkKkWMIytQyBNm
wqVzFO2vCPCucWvtc5QLNeDePAXNfxTeVKda/qdIW1kEGHb436SQOIGRKCXx1iB/
VF5mAM1aVgHSGCnm8StzFI13oCYTkZOzzh9cIGY9o2zpvKSdY7vqqlL8zrj3dvwv
Z+7eBr/kQU0ksxwLOUUs5mUrWgOI/Sy9Nt1oDBe4kxVsNuJst61GOGNe3ZeICU5h
irt5l9W8LvHo3Oi3aSHS/DWGo8gbvBdG6OkezwqLPLW68ttgszaqe9HTNARqYJAL
40ZxfwmECg3mOJxQ+6WAH1mHkJTi1eoAg0mzxQT9Yep38Zc831SClVeT7Csof0j4
GPIhZJPIz1nwRSACmj1pFskoIb/NEITu9NUGbwoa4I8ssDdcPECtcUE8ohicf7Du
42lhuPAz/yYL7g+MD6QshTIdGR8A9unwuB13ZxmUffCoGs4kLXcxJ7YFKqxJo6u9
Po+ej4GyoiQXgKuoPQTvfAdnTfMePKHJgrq5xcMQ+er/M3RTOkrWtZnLqUzARgts
+Espc6pYciSA6ysghlJpjHF3/a8yBFMMfL/0KShzk4bpjJKhumzV9aL56LcLyT4Y
SNfWhchxylaIt3vFnnBTZc/iEkKgaqtJ6P6rUGfj8Bb1FYZxWAQTDAwEnedsq66h
024kvQADrLmD5FWQ3IEiV8Ox+X3JbIJ2+krx4/9jh35AKgOA05Wiym2ZMVQ8X0q4
LKU/1Qi50DYBwx5AgdCwK1So1x73hfh1GwrAe9UsYznYyxcNqH5FYAmYOFWgmqi8
n9Y+Y2DrXh0X/QzrGyOoEDoMU5LeSg8dNrgyTZm6wfQ7731eXBzOSbSbt+IPoviP
NVxx/piaKdh4S9j/eOs/NpFUAMky4ebMMisdAcUGUX/r9cBhPuf3+JWXwbZvnhGA
FY7qilQTHajrAHNhmq9sV7itREuchLweDIAcejhFSiOLaK3oAD+5eNnJ8J4vySj4
7xMiImdz72Incmhn2N40LB5L9XGt5kafrGiZfTOtzGLDq7L4n9X1KwGMc2q2+rur
nRvawL9/G4H1S68ayER9vT1A15+oSOZ5zx+uBqU7h5eh+5wgnhiaVxEnya1+7T3d
sU2kLHa9HifhEFa0T/3JxuSFd+ucqqgdcfpUbFTrDuMilYh+A3/WUwNhLZNR45ir
TO+LOssbOnpj8yyquBF4MUQHP3HdZ6TAH8Ve8WWyQZQlxftGmvddZMOPxnhDve9D
yhUv+30ct3TCS9ruOu1OxwWCQPbJRepRnR1FxpSGFBK0I0GU08z5mHpDwaQbKouH
eMmOmXHNVnKfmnrrwgF3MsKSWD6NGj9saJUliU38s631GxM/6Hh/4w7BEAZXKFOa
NgqXaRphJQfrNdziSxhet1yYpS/A6r1Am4ITfGYUz505eQWdiodpiGUgZl2tHFhX
ctzE+JZ4uiO+RNbKBfDrEQ0Hd8R/PjAuhlxZ21vOhP3p/Sv8QXnbB5w7wJE1yy6W
dE1JONLulIG5tON4TfWcvjIXWQslDOEQE761an1KIKEKfSja2y1hW/nAgE0wbD9H
1GK4ayBszddFrddCrkpYOLgWDHNKueanRLvz0GNPjygVv0VeQ++ruiTGUhpjusKl
C2EArhE3bDGa1F9ZnqrPHePebbDbqOd+YmPSZEboXOy0FK/pUgAcqlkJhrz7SmY3
4dDKp2we8xBas0is9P2jsXevjpbAt4sw+wC1j+hwNIkfEI1yrRvPDXBfS43Ra+2Y
iQL/caNcxPW7a+msGyZR0SLo2zM6VBDc6VqE4G9zCtwRQSFwlZ7QLEBQ2GLGvzUh
wk/A0k1VlfZLLmqO+35TOjJIItyti9/crI0lY/pi21eqyt1ZNbZmCUJgLUJx3ESh
UEaNhMb7LzKNrEb4pYkIhuFHTtQMbls8SxtgbNHbBSPzV5XJa+ddSBMD+TmkTji7
b94ECL9R1cX/IHfhGljJ3hHKCG5MwV0/E20B4xoPrcdmGlijS5j97rsP5DBgGc99
tlsyfUY4L3jt0w1bIGqnJ7JWdut/Y33vPjwMEgtqsM/4TnnQBBE8C6a9lnBUz/Pp
eRQERRAmAWy9Oy8PsTq/o+RASV9dGM3J7/BR2M8tBLNZlg9sSXztMokz6MGtnoHW
O6iBA63hLKHoEZPYCOit214TNMl8eE6r7ZdTGOk+44U7FTQWiP/wE2NHQagc7Awc
yNrfJw+0L4Q5YZ2w0pp9l4JICFBzdsCezZZiNE/PkWKTPhyl7iTWKbcOaFn1HfEt
JbqvUIHJKQZU0lskJwRxHnCuIx8YM14Bzbxr85IPYpadEjQp9i7OQ0YS1Dg/cWZZ
6ELpcjEXoKY8IX/+fDcZqaLdpi52wTrht8DzwIMwCYdm3VYbwU7em4uoiFMgQ+vn
trt+Su8Z7Y6+kuNSPAOg6jARFVElRpjrJVhSRlKJx+Vpg2EqQQpdjy+6Udn7oehv
PoJZ5ZbKClNXGE7BKUNjJaHTqD6Y0GpNZrDyI0DLg0FS+vZAH2fmmsKzW3BxlTrd
T+eUHPBUQNjmlRa9wf+4Foso22qPu+S4Udb68Rn9KdLXz/CbOzU6Gl+Ke2B6OfdP
1z/2eZ59X2SAe4/0d1QsETuoj7Bii2oykCho6MdmuvjpCkIyUNnhQQobb/6yfNpf
eTSfGUny7aBfe/csDBNPNjVSZfMwA0dHXaAwxNDCqsZuwjfLEX6O102HVOAcWNou
+CsGOX4jAylu4zDO/LcBt38Kx5HyzvYzWfENd43q7yKIjzIPwY9hfdeme1R1yYuD
5lyZkxFSlyiBSs91CrEOBq8D2fJcyKWJ94Hp9tVA/YiqNyIgzJgwG6i/Dfx+X47G
brznTKJEkBJ5a6+nNGRi/9XPXF3IaCZJbAR4sGSntLDyl9ok3R2HDZ01AKmzVRvb
U2rLZkUrV2BTM/sV/LerZjhRMiqG/a41hAa6pWxMFgUrkqpy5Jvvr2MMIxeLlRyz
PxlTT5oZxaIcEkgdzctscc1xA8KW8KitFWeu/gA4KnoPjFBf13eEUXB0WBCFjp+D
fzBIHoggWONX3U92aaEMuWKVUo2FckohjXSJ3r9mfVtQrS+YvFDEiQMyasgb9Quz
CmzDviNmdideYQY4hE10n8DHqeG/iSO5Hl3eUo8AtlUu6BS4UZd88nivIlxj5FW7
7z2JYcTOxMhrMhajWstz5eHMQV5SKgBXSeiJntimWSMUznsGyt/fIVl92fT3qvtr
nw9btmV0QTcdidFXRepmL5eP1l9NU5UkKr1ft5HD2HrVi1/8ZCcZsAl7U0xLQL30
fg1tnvhPmylLp2pGxW1EKGvPvvM4Br4KR/5vIt9synkpjvUaaHLqlvpGEvZB85Yr
Xay9KFWLOMKskoSVBmv/d4ll1OdUKsmnl/vdDqWiQ0B0nxrbkjI7fnaGzaQ8xze0
8LA/gBw4vJg8fDa4IISb3RUWwNsZqU7k0xFqnLfWI/1wDYJhktWWlXtizGa4BpxJ
fI0cE9HQyPGCjmV4wft8ZoSd2iYL/lql2is7LJexeTM0rzigulv42MzpSMAM7X/O
zzUpk25JwXVf2D3/UTRFrNF27xwUKTbAWjwlI5T9pOK9DkaLgdCQr1kxiGNToWx9
eR9awYxLlv0yjJEOWX4b+KKvubSD5OY8R76YSEFu4zk0imeKC27St+Qn+k7YE/mM
7VTKpsssUQkSkSPAq/Fu/eNfC99fHUIgBIchc/H3taZfGhdCGXj4lkrTn3Z9dMj2
jVjYBbTHrLfDgVe0mSzOhsUT7ZiEXzP23ag+9HpCW6qebexQfAS6x2eJc0xOSEBS
zZYvclS2VHViQB8gl3zxavYoE64og0FN1Ghwms7Vx2HI9QDCr7g7KSuq147b3bAB
jYDY+Pa9FkTIgtvq04/gjpBuHs/oTNC3YRcMusC0gyoXbZ9jAWaD5adl3hYvDFBj
gk+bhWXnQ1sJ6fqeSK+5k5MdOP+/EXLBMwsbJSOJi0+LKhvHtCkgBX9vByNvBTW+
uYy0vIxzyQ1dEFsbc1PBU94m3eeB4agRdCJTZuwLe4oB+B/0yMtXIRYltwWJSo9Y
jnb0y7g7JgHMhtuX1sOjK9HeASWZ/HUy6INpMQN9BP4teY/sF0aXx7DhpWh04O8V
S3ABE2izq+AWeJeXU477qJlSh6SGAOQSY6CtZq5JItDZu98JmRqCQIWPRPM2xocu
N5AF/AEBRwK8GDkXaj2m+2pZ1/jGuPsIBk7OnVQOkGJcefsuhXhUi4jLfyqFW44i
2wwaP7qej1aezi2lEK6+eSwbJ+FIiPUZUdlcVv6ed8s/ZoW28Tzvl8MriSJ/xRKb
lrpAadDzAFvpuhpfdJuhqCxC1c5CaweFS02JVMBPwx36wXDTbrjbNocoBd5kn9a8
XYg7pN6LUFLbNpnqDlXgnhCYUNkr1FXNy6U7IiCEU2yJTlEXoDoijzY2VofD5HRb
fOjOGul5/IkJoG7re8ao5EfLhnW2ADotrK4asj4cnnr2tEXO16oWLM98OEv6ypv5
4X15nZO0H9RzlM0q4O0Q4chRthvpyRMkTlOhlKMmxIPUzh3MWSK3T0YNi3Nh8sP5
1B81ycRGtPAXlGjVldgHHnEDw/rmCEa1dZ8ck3fLuM/uMJTLj+rwWnoIyVLtn9PJ
eg+hZBIyJOg1ksbrCqgz91Kaxnh6uCdQC+ui24RbbPhv/xmbGH+oJfRDhv/W07cB
9HORSiqn4sJK7V6RFmHUSunHJgKLWN/KWOmDdZzx++Q5sZrhoMYbIgdifNG9YYId
3VhhrWNjIiJ8nhptfGy+Vf7pCiYXKWad/fLQNwQwsAOqhNW+1CzdlrgZFAwG/VK2
3CBrLvzLdSlQCM/COm/Lbobjsc3rFziZeBDH/iafTTpobFzoj5RwCfKq0Rm87xfc
FRNtNmyA1quu1iF0IHoCJDFNS+eOE3zisgCyIh9d8GidH3wrVP69xzH7ZXcMMesW
r+gbrWSnY98s3ul98i3F4qJJ+kbOnEQh5Wr6Aemo/+4+Tk2FCtMKh2c2QaOYlAXj
JDHishYBq60iY3ZwBXN3aD3gWSBnVqab+aCTZ734rv3iViz1/Kn24rd2BKigO/pN
DNIf11I9CbDNLVOVHKityVUOpa2hR6Q+napUTZt6IdthP6ycvBS+zZLFY/1xrHVe
D6cy216TYKelNzbalvqvj91F95qSXvZ16PWdRirGyHESHOnmZW0NggWZ+PitaYZn
kYI0rCA/UV43gEPnISV3fkC7en/k2L498qsSUoCGgBMSfo8MkWykDSqiBfijuOZZ
XDkNyDQTpRmvRyBAZlZw5hKvFBck4DiB1H7XtAw7m8gH0A1sWB1y8qFtwJKH178c
PSdfVUI4ZQR29ztJ/3vxPBziweTv77v1vjMkT5hcdxBdvsmVpxCMLkrh3KFkjwI4
RzW0u8E46vqfE7y+dWkwQ0owYoizmJG7lwMm7XxhiLi9+Pout4x+oBPptFZPO182
Ry8KHlE04m0/q4MDtpuvPSczbNJU0Eku3MbV6v/d8mnwEWqrIvImiq6za4fBbxkE
9KHUNt22vN4RU/PUhn17ZZPueh97JM/NS4i7etzgL1D0SDJvQb5Yk2fD4PDq+3xg
RFN7r++5cG8mxE7pFv8+wN0aDZtQW9I6F0BKr0IOPIxI8p01LblAsPlqKdVlOVBy
I4gHq7TuqdytKun1kdNzpdW0VkDK93isYZHNBxFAaDdHEZCdkPC0Z+2rb0zdE76U
MTO5v7tElQVx04SUYDbI3DNh0/hXlPJUO25xYuq3Dclg0f5FV3MwssiDuXplBit1
zQ3+6YjkflxdYPZmI73KSb5VzSsPEQAaFczH26e1ZFwTRPAwwxRLv81YF/gJmrgI
3yKv63QLeTxgWe/j+Qhpvuy34froz+DwJTYRAa5nJIaF+qUrLKpjkJPlKRBhnfeO
uC6RPln/7+vQt/e5agWcNwD9C0+/PXGbVlQF2d1JIEaJEy+3ieMNfKkY2lciU9eg
kegxSukPo4nntjlXoF3Z4iKSC9s44Q+nw8WoYmuDvL/lp9j/Y6Y6ioFmAG2x7n35
G18mzFF9njb0HfI+bZIZ4Qj2Df9CI+p2+7L6PRsyPYqOTjNwyKqOVK0LMgmAVMiY
OwJ00r0/DkGBCahuAWr3Tf5AsvTVNfCa+vl70GPND5aU/5+DNijQm4tQLOTTULtA
QI9rtVrYWZFoN7Vmn51CkhzuhEVviYRATGAt1HZ5M23giVV/biriKGmxYgl2ufo4
GLccUc2HBuKBfnHQU5vvvtg0HmGOlN/IXgQUO8NPidJgeBmXVaulMld52Af5yscQ
ac6YaNUcOaP9Y1GKQJpllknnO4XhxKz9inF0odqyOPZwxFF83o6VSfG0YZtyVRB8
Bpxb0Stw8GFGUtcdzNeOCwcKW6xao123Q3MxEOqNdjkj3HtFL9XLIo2te+WjksaV
08MdX56xTP4bP2EryzhZdESHkPIq78tci2eA7zxnwMCgjOjkbqfZ4psLXc+yFINE
EKyaSkYCo7gXowbpITF/xPlCABzKiQgwzsHgO1H/wuKhUKaU4TkuDIjkvFOo+Kxp
FnMeeq2lBAWWdcWNhlX3jrnfaBvmJ5/pIy7sy96u2JylKU4qLpvjWi17lszq5otu
JcHMK1crOXhDEgd1CwHUUbd3rZiwo8DL7TpTbxNsk2E6r0Bmi0qgbLAZa1K30JK/
f4vLbYoD0sHNSC2pyiyvE3wjL44RYrwYLJYcfnTSoWZBRmUVn3iKC3qjGetOQJAn
z7RGv9feDZOKgeFKjb9b7b7xD5h4Oj1lz9ykCRjcsC3GZi0BsbW2gCrfTbD/u9es
sOp6CcQqwWpF+zEyWpQw1RCbzgprCwY1NWLtFZFQl5uTMVRGHJ+aPWKcZukwFjdO
1eiyuxcprnZQlLSmQpDA5ixmhzRpN2L4igW3e98ZpRmwXLJj9geyCN1ieILbm01K
D52/wEDWTn8qZkNy/nBgmClsv+P//jCJZz4M5LMEQQG6PQuRwGHQRfYqz3tWd4a4
IYWwILh9dqqa9mG82g+UBv4AvuOPG7ZXlcouKSOy0lPgmKgsu1Gc0hb98RP9EfRy
bgOPSxGTGVaxJaUxBKe0HDgEw3OVnXWb5A5LYf209VFct91CFybWCffdSMAFd8Kd
pf4T/Q+3zhkg0KLbm8jA9OQaFfNEKp+DP89Smnttx4tXca2BR+0oYyEeVNU4nbQK
frO6GOzuO7JLXr4/Qa4kPPJKtKulMDw9tYcN0X4KNbmNMjSVJMCP5PkIFJOkbCg6
wcYGecbMrviSXdq4RteWNZiPbp6ZG82UsJxV3vtiSGb+XhyBC6KUunWjLGOhL3TI
gSQK/Yc2Ne8nEoczBXPMeBwVJpQxh7w4p9vYhU5ZgPpgT4gdJ3AOB802pJ7TbqgX
WAD3wv7UqW/OukGBBBiFi1WiHZNv1fE0ePV1FQjNMYD/4TyOCan9KKOuJv3/g5iI
xExp8T6swHsw5lUlC2FVKU8HRUMvv4aKgB/t9e8U7gh6dGoyxzZA8Qfb6bMSguxf
pAeiXz4wvJC9DrS6DLZfluX6N/yLYErli8yg5egZXnYelTgWEAazjRPfv6IMNOvh
T479G6Mf/3EMVPlSUDmag+R2kbsF4lLvvEx16LfgNiKyCGh+8yHnEqnQCweESi3M
cDGTsN6LxzDwgHk4fSqPul21tRhgvuTLYmxSbbdy9dTFfZ3dz0N1PAxuerP2vMj/
5xkUIylD+D2slyj6mUw9+q346Fpp3YBE327H/sS4TMi4ZUcFDIX0GGtscQnpbV90
9fqxdDu9wW3R06+/RTmNZh9tZFZY0eelghnsO0+aVmjMV5SSQpY+tom7A4leUdRE
2kcpBwNequtCoPUo2Xxi0OyfHO0dShmnqPYyk3BQGog9T1mFrMnDENDtDtravJRW
eYSROA4FOeFz05lYYQ6ckc13R+kzfjuLjgviw5wGgUG/9kMBu2YiqFkwy2+9w05f
xijt9rippSzhJ+i87iybZzkWIcWHNRyjDMFv5SAT5tEdHGcIrpWboEM/t+rHULjQ
N164t8FYfY1rcTqXmUGj6GHjOgmVOQxqQF3D94Mb038YsJ7qpYiiSj7JLqkw2ON9
+qtwJw0o26ECpT0546ZAfKiftMvMc9sEKw9m4meZVvzaQfwafCY6mQSeV5CiemxW
4dDCuiTgUl33+MrDIrObaI+qn4VgpuZqpMsK/6Z65A6okv8FN+GaXccLO0GJsfX9
wbyed0OSyYCxpV8dMWz1UYqQVizRWamX5OHETYfLC91vHzID94a94tjfp9uQKnqt
A4M7b6DIo7KeeFlJZOqW31CuokOZsvExFq2EDcYlGOgkvdmM0xTU5Z0tqJipkTO6
DTPXGa9tf2Ro1+gcNAtmjdzZaroUE9B6Y6X/kdfLllTn36mlK7YZH1LEar019+/O
sW7BrKsz6oZV0YMCpmBANee6gXSufqCDDNQX7MM+5wbLrGqQQhkQlVFtshtPxEwu
eZcyX/kWHD3QaxyVYOrz0NhvslzsiTHSMgHn1RtUaXMdfIV96nca69rA9ElXEe2a
v1OvTfD7RW6AlLEXJvHXfdYpDFR2UOUKWx/1tKjKvIemycIULhB3GxVEBOuex6pQ
8ZScQNOwdG1OCBoLN8LwezO9wtI0YuaguEuIzMe8vp6gfIZbue2JM3N2dhl07Dz8
uFxRT7GNWE2u2z8cLxsrby8sS9QTOnL71pk0XcAL5NpSyepplgVVevh5Zd+9uPB1
CPkKa4+40IxI5hbN9IoCEejjRS7ycB4eufLZrueZRXGuGRGWGBXfY5POOPhMvKA/
C1ILFE4BlhaqYMpqqqQBLUy+/b81pXcJiKGwu6DOeycMR0TdneqicbgJOtpfPq1W
DGs8QTXX19jZumsU6l5oS8dX5+W6jv6M5D1NNBAt2G/TWjVsGwMiM6byymMGPDOS
+ruFeeCvuxZQRu9UBmuQq7yIIrIej/3aOJKQfb5T2nknUButWadgVIZMoA73NCJY
vglTzOBxz+0cgI6LxTOSIqP8SDPdU9YoF+O4Ybiei0v5D7vBQcvwO4u+Y4nWhZBm
e0F9I4FEirgbF3oFvMgNGjgU8lbijGWSvK/kp/Ns5FuyVqJJ9fNUQWhCwMknknjJ
8nGgbBJbP5dzi+1wBS1HJLjIgLGAkj19cRZXFZkuMls2327Oy2ZZOt0BLa65Gd6b
LEuK3K3dNZjOsM6fTb3VvzZojjxRpYKNR7x11gsk4UhhUubDnyc6HT6QBj+Egt/m
lkUT2S5jD61BBBnJoun3k/k59L7MYuOR6fH0fpRb0E14GxmLqyEnVGUUFyQBuxlj
uMcQ40JlRc25/i7K1lwidyvIsm/i5itd1lUYDg7wUmTJx/nKQ0izXon7gS2cvHHX
nVUWMGgZrP6hwvtM5oqW875vgtgUXS0fidFm914CObEkTgmrbZ8WQaYn7UCxRqN1
40g4F94EQgOUpwFLhYcr5HYwH5O1zlVB6Oh9uTMjGQcw1jwSk8WrNwVIRXoucO2B
Yb6U6sD+kLY/2kZYTlKeBxZnFp9XhoRnYnrwuvahvP4sbIIE+GnAjW4yV2FBwBVl
SBJGqKQ02iEYpuavbHSB3xl6z4Bi/rCt+l1nrixiC8IZSmlqu4J56XZ16Mu3f4UC
pGepIrGVHanaBFWuHNGL6+TEYIRGM3USBfcqLfCUq4my15bLJsRhYTcTK5q/09eG
D/FbLETO4bUIUD2a41GGbUexA3U6JnoAMZBRATpMitzHe4gs7/MxvhqH7Ibazfv9
yhhetLvyjFL53PQyXfKG+PRiRfHf3N6K76C38ltZystY3UNuC1UudSZB7IuPMpYl
DDObfNji6NKFQR3SauBigXnRu3GLkW5UKicDZnRfhTGG/mAIndwFm0wy8gpgWKvp
yl4h5020fVbwfHr04r6j6cytq52eJANbXqcm/kbeB2mdPq82pEYJhQdm8/gJhp7q
6hLP9F0W3zKsiV/QoG4dj0ADDTy1lm0koeoSzuCd5FDWI73vb57MeZOxJTxjBOcW
dh5EAn/7QP7H6KoStZ18IWeAd6dbvvRgL5TxYsDe+fonNyihvQq2gk6x0gQGXx+k
D53o5j0sc/Lr0XZyr+QIIFJc34n0MqENUZDQircqmjz5QzymR7EBJXJH5c7Vuul2
XuXLB5CedBAFlZiClWApkz1/MjIEDgyxzE7EVdCZh/N7V/4zO4CFtPXFigq0mFYe
SbcQo0x5LRUyxbhs9zVziFgp4y2ZjCZwWeooexU7GyMkkacw5JPLSDNz846UKwZ3
zMRvwlHeJTxjKsNhmjvV9iSxcMlHty8CX0do1T7jo+H7Uq+MSuvCcInDkv9m00iA
zvAQXKdYKn5L9jo7VWUkSWOP13Zl03pPCiwziz8RhaM4+FPOROKx95w35m5L9jw4
w2tg3mum5eH3VQhk9jftlYc3uOWF5quuXD4tS1i1u7c7wLlbpwlRxYYjnpOpDJHC
yaHLLDHUKCxScVNTEkUs+ueR1PHpWBfwKKrd0eBjQoGjzxpqqsI+nQXV2aNbOD7W
UNanjxJy9A4NsE1nVEltu/uLFu6SAz5ze6iWwacFS0iB5RLSoXTEieNvrTRD2xcg
l4EzQA62bTr79OvId7MOGhDuh0jHNw42/qhYYnPt8F8JlJKMheWRmBcKXWYRbi5C
SNAjFyM8b8rShKbr/0pJQ16PzivAOH2BtceWmf9vmV6RadEzFJue7GLqB0OP7+KW
BcGiJXCHpWWxtm0onJaJXGGFwn7t6VDEVXfesmjREK2aHqIXFAy+TYcWbJgYHJyy
Z3lsxsgx2CplwJhKKjVyfLLdQK9DqbKja/ecp6kL8VTJGfrWwOtQ04Q6v3yz8BKe
GyXuag5ob0rzO/sn7FcQNi4Vdbd1Gduf12yrVRoYUuSlgS7wmZUfsuIeWlnB4KU8
EsNfbA2CL6yT6SN3ca9caxcRlxTielnlgfkI8/YpWyDPbfky9tLpyph1n+9bYf+t
/OHL2n9lBasLYr9jOcEt55cccT7dHkQ4ktn4VG0MMFgvwNUJ99XOBlPBaSXHFxM9
RgHar5ztPFH8Hp0hGlVsDiIqM8NXORT6IPHqiDzy4Yex50jdqzocLAEAVEywzRr+
VgMBp1BtfW4uuKVf5WQM7xsoWgh6088XHIGXfHv3rsgnyoJnx925TigE6mhUOETz
M7R/PGVcbKoarJP69tfqBiZ2W7IUtgYAS3V7Y3lWnGhFxFuN5H5MYjK3ZHDyeAth
rySfHtBxa1xc0XLqV2zek9IVyiOf0/Tno1U9aDcm/JxjYuwhgwogZWoneEijoSct
fPKHQ9XUz37V3rYPIWKBdeTD+ZXzWIklZx32t+ZZHq4gevESOxvlgBPfgMJgx4/5
d2QtWkeVU3L9Vd4DgEFtjGgXCitqDpoJ6ImrkKX0xpvsIJve1Zens/UKhHftcjVl
/qoINBfeLzQsHFac6+RKyw9/psv89bWN7YDUmakjaPaExJIAMKYyu82AO3QuuJRH
Z3IklT98k/5iSBW3EJ2iZ6sJ3YooIr6kzoG3gjqbCysO6fiZXg9lTQghz2czi4JL
2ysaePPqsRKd6OUR5CO0d6jT3u5IMX1JK00ThXFI7hEjiOYJ0rOwkguWR5iuqD68
4TH2N2O/CzBEDvT4UgHUNPtLFyUi42ypeWpMTRrf82sVZCD5j4RrIUZGbrikx/O1
MHhDQaFNQ1/cG1uZe5tx3fffa/ntWWVV7TxblmEk3Estq8n+CNJQrjbfHbPMAbzN
FZ/2hFp2PpU5tZUxz90OhWhrySV+sqwH93trNdZgLjQM2dlkfLNYtREUs8HqCPvz
PdG93BVWRcHBzPzd1iATV8iXvMZh3US5Myakmte2y5TLhdXR0u2Q5R6qAJaiez9x
AcyX+HHF4+ur9/hO2FddPlJP/hFSSnpmTuy2DwMVARrJWOAwbdSM3mETYaflLNo2
GcxhHGYzFCXAD2jdHF4DETgOIYqb+2cwN8u0A/yc0L2IKlkX4Ua5YLRI6DOalJoO
9josJb2teyDVklSRYzlwiGH8hlB+nkINxHL7aLL+4P0tzVf4TNYdDFTS7u7AHb6R
M+AbJIQH83kcBj40ycYjd60gqLMvtSnXFQh9Cjzte54gxtowyZsi6mbLsafZMQqu
myIYSw1bjB7mOP75OhKDz/9AocZ+KgKpOc0TKJhx8pP01oxLCquyIoVjj5LAMUcp
e+scJa8Zary2vtc7oYKXRQs2OOHKYLt9xxKUz5+1yJZZJnzHm6+Onzo3m9bgGwL1
gV2PTP1hbyNIuZ8un8giaMc09k+uBf6dlhy/eCaV22gVGCv0JfxxiFG1WpR5MnK/
COBvtgc/9SlHXk9evypUh9cyTbJQj2uocJ9N/XhpL874Tps5kSc+nqactokqJuQg
oJkhmBINQTErejxfnG5Bs95UKoupHVDwSkzalTjmFgNzn2c53y3jO7ZVFs15Tmtm
0RmbpHWKxKNootNcAEslCDewTqgryMhyyM6UfzGQEDpcM1m9AqyMkWrf918wNPIY
GFMfAuFjv6ooYHkjUyYieGj2+8FD2wGHQXhGSlb7EW7S3tVrW6zDf0OJYUg3bhuA
2yCEMHY7G8hMYb4GyzRHKO7+2x8ip5zK/5rJwPW7/9E32HvkNlOK9oihUROUk2Iw
1y1VbKW03RWv9SV68dgtWi9Z0GIGRraDpRUYQsxOJRAKiq4Udfuzr23AwCzPfnyk
TOnKoNulT1mAikCeEi6iMsUDHBc/qW8xodLPQF+kYaUYxcPiXJByShCkYPGfq1fb
N+OT0+EuDv4ScUxj0rGq06Dmw5w0VJmXNCP5m0wLz1LEk2VuapUJ1gyw2PbhuBVd
zfkMmFckGslvA4NA7AUhdKMa24dxbZ8950kAcnuEEiGs1ty0IT19WZCnF9lQpuNs
xCpssBeiIGo4NYHrZYCKMpn9VhYOt+K9uWxcvSwWNPbHf74mFRwvpYzj99uDvAiB
gRy6xq2djGLuFK7k4Kje3xUDj7AUj15FgX/GBhGH63bzk9RjSYnQkkS13XHfse8p
lVlirpifsu/Msj96vVMSL6Q9xpMW4u557FstT0YjFyJ4iPfGXVlLmC3KYc8pPvgh
Sj9ZaGp7lPj/qeTY0x4IwAxEuuJE0stko/gtsQfqKixyKr1QzBcvO4ijJ4gp3nq6
WHOJrCLCWPOIzDsFwitjX7Gjyeq6c1sn3fJtBVZbHeXT4tHnfOh2YprjhH5O5Ceh
q08R4WfDjGuvcAQ0xi1O2rqHc9VQyOMKVf2nH9JieQF9yGakO9I71I87JSQ3FREo
N0hbvBfTryj0spTnIye9bDEn95oy8XuUUB7l62rpK7zddcxeHekiRZREsYuOzhup
XUGdThae0Loh8l+slP63T7UZM83Jz9Y0zaoFuzA4MjcJY7Rra60l9H7tzTbIjs4S
HiZy+2dXKO8vgBqA9WT6cxp8/KzzJf6Tc9ezcH8JCfr7YwMRG3g+MoKW5Q5EhHh2
KZ8k+Nk1kAyINmHMVZhhHXBmW+MMsCJ/W4er1TY8y54nlq8FfEGhdoSBuC9fZIXi
7HXiZHlX+mYBYAfsFrPOEQhqPxusbwZOXpP5825Tn1xQBzM/mDz51CrFKI5OM+FX
HNRMltXW7ItyD5TDkD/l6wFEPcbpqYywHCkfwnzIii+E+mr+1QkWKsqz7mL9WZA8
WogkTVVycJMcSsmwvdP9uDIEokjn7s2ZventlyR0aa11Fz0Zh/9EhiuJfVtKcXFi
xyAFlI4Rl14xwo7eQb4AUf53e0b/0gU+2PkidT+owuyhEgrZ37lfEEe880JGOzkL
3bTgrLH/VzL28NgC9rOVJNIg+AXGaa568RVjIHwRUeiVbKj0SA2OMjcLRsb7okfa
4dCEjKMfRMdXGgt6qirOq2UD4aHSuw36XZvUkBfTJavJVgXx7e9lKjdUQIDUnoKA
E4C2VfvgQrAKqhULAwDu7Bjs4gDz38VOmAnNFbOObjgjTHK98u474w4uv9Mhs9lD
2mN4IpXFtYyauJ3joMs9hwmvkpkFQr2TKqIN+NhzOe7jjcJ8tgRK02XMgLPRW7NP
FvPqL03eWff49VPw/25BQezLnS1WfgkY0l1MP61deEN40BiKQ/sG/3/FrmDBw0ZC
lI/PDxSCj0h6KKfKRaa07Rp03fj+LArKM8WZdklg3ExzWYTyaUkQEyk70t1curan
M7KWTtuSnBs1wgRfY61xtt+IxO05RKyGc6JSPYAG8J3KvCTdMeyow6Va1aJEbKlI
dLDUCL1UCCobqZBiYWNBg3477ZqW1MUH4lBQj2hpB37NGa0yNyOO2ialPNoAjwBP
shWpcJgHaBYAg/igjDKnzin86hfEYnL3361T3trh0Kezhc5fikTdGsxBJRkbkZK8
N2XOCh0Wdv1uuoPuCl/mvnb/nTN/X9lIHtytYMM581Px2kfAHNuq/V08kPCxEgc5
RU828hqwbRkoyu8jMZ0vh+IR3WTJpddFzTPf68K4gqCk4Nv4WqVr0m14Ku+KLKkX
j1+xHXj4ofz8B2ezft1xbL/FkG/CbgyxzsekZzMuaeAX45mUQaJVc2BS8Ci503WN
sZEwCK1p7WqhA1yYMXxANh0m1qCTBJFreBZyRvi+36BFwjy1sJnuB2xrgTtcBEmt
GjHs2eMhpGBiqLl5m25UjJEfCcfpjlkGFnF2DhT5BL8Uf1teVqKM48cW0ewAIEE4
81WBclayXSWQ0cDjTz7q2Uqs4dNN53KjdxFLR4xTT97Yz4BHxV+OjO+E3KEBYBO/
3wuv0eCB2TO8CrWOy5qMwEdbpTcNu8As2v5tt6FgSD/73B9mfbQqrYnzV4TMNlHl
PQb9gC5xaP3fQKwiDHYqCTixC6CyDEvXEszjoeVmyqGxM5gDjZ0r1s26BUZUqlIR
DfOtoTflzrgqd3xFILRO2HS9fCw6pJ3MBPUty5FmM0vcOn/liFV0kb2q05iqtmT6
D/A86VzLoIBPDkhFAOmYOOSx4w9c0igBC5GpNyekwUzfEQPjfjrhEGA3VG1wG4pe
kmHQthKaEBD/aJSJlkFL7IsFaVzuSS/Ea/mq+6VKtL1zSCG5cUL6UciDyelBGLc1
QoizTI+jlpMDujy99gnTFbBXs7XqzAkQ2NmK/0GnaqgaMGVK3yaVaei2c2NHsaXS
MNAwuqbCgLL8bm9ptjjufnPLaWbVGI9e3/ri48v5s/Qe5/zkS4MaDqPz4Qc9xIOv
mv14F0CeNdNpIcuJGSac+3LxrMDjgMZGIruX+kqGPKYDfuRgMcPlNioF3f/nsl+U
sbi6siKcTvuazJM5fPscZCj9RVqt9eXaE0S3UZqjKuY/Fzl40gEF7qxbIig7J4Ji
w2ardqtwTPozI21LPh2m3a47/rMW8DVXKBHywtGXbj7wz0Z4RxDbhS12yI+tvRXA
HDeegNjdiJ/cyhN9t3wTUjAaWzmNTFfRC5ngDuRJGhx4zTnPCAxZ0CjVAbv+UaMU
E9Y7s8gJbSe4i5AhUa8yrPVKjhK2Dt2kRb6WFHxURBHdJI0EnDUz+TXo9hXAPXYE
RMqu/Da1UxIdG96wAO2xlCoKWj0ySxlKn3Z3yJuL6Zwh5E6SXCIvUwesGTAf9Qmy
0F3XelM+ZwLUixP+BV9zaUmqe5SYHYV65bH23ji94xzJqKrEv3+MsasiLntSb55V
W+GM4c2eV6kKvDHxZXLbKoL+pcprVC2ft9WluM1XXyKHxP6ZWYGCPzaLjd8H2jL9
J9YrjoDBsFCwTIsyEJddoJ4dXKsPXAmxQ3BCpUx38KEQRfBU3zkSwZN9wHtbA0CK
mklYRISAgNkg/DVwkh5PP1mgwqid5B+UYo9Nawf7YesAz24O61ktZJrxjDYqL5jr
XlppgrXqnSr5E7vjIX/Zf11xOfWoopCm6tYdLyouG42rklKstxE5+Y8O3ennnit6
fQIxBULXcXti8GGO1d3vzGi6qMutv1cdaF1c5J6AAExdRYEerFUQ+iX07wNmpucm
38h2VU4vnOUEeo8Toy5C5nQmLW8wHeNkGCciYZIHvywbEx6RBDAgSDSSPRM5Ely4
lZQR4iLI66wp0ZbcuEFOZfZySS1YjTVJ1oeBK4El7zxqgbbRkjIA2C/sTtRuEN5O
3ejU1QQJgLZBkvY4h3x8tu6Sohi0gTXOz1Nmq8e/B0/8UpWbKHanlXp9ndUk5r9z
iQgm8iLzeyAfQdo6/C33FaeRv8R5LH8+Od5QYJMiMi8+K6nWOoJ43pvTpmxqHN0O
FeQvCylFMro/tKDSfpLjSnL0/pqbQGZoiyx6ZA8EcR4N9YB9/rfsuSmqGOumWIQd
g053CMDM3figFZjZwngD7W6qV+d8WTvs1P95q5NTPgtiN7clhljuhrNdcxKxPAI3
t8r/bqb4PsdqgjT83/dEgm3JmiGCJE11k7YSE7Ab+xedmUgwUxYvgc1+128S8T8I
WHDpHI66ItgtCpdGnu+D5yCGoJl6nUlySPd8Mc9uxFp+r1jWPPgVI4JaFfgkPYpS
5zMCNwD/tMnX3kq5WzBR4H3+cwOgeKV+dJ3R0et7MrtinGW23y0VMosd9lkTIA0O
8BHHl515Um9Ilt7sLPfn6cAa29m07aJpdEbEFGR2D6TcfflmOWG8d6pojp5C+ljD
OR0Mm3aAE5D8aYlRLMd6R+3oss/qmrAU4lh6wp4L4MRZeNoLwuNnCHGZUXdADOhs
xC6ffHIMgURWA96CnY6XjkySGIpaUT1iNQKWV4fOf6edreLAoWvQwXDs+Qrhrxa3
T2yHrejpVjfIMyijRwyLKdsXrgWiAu1twtnXKSCfOm2Tgf5NlhPxyFtoV6i2nfMo
2yQ58bl6fvwgOMeLS706rZA2T8nngRyv42DP2kgypigTA4BgJudqvttnNn4+I3bs
JfIrq5phONOJEvRO3CzzWqNyxNIVEnhgyVjEvokhA684ZUoL+3SGSt4U0lOAdEO9
06oPy1VxcLAEztESDq1XslRWqB1e27+vcYY2AfV6TKd6shfITFHsuZpXwNA0BPuq
JRhVBL45PbNNUYtlaJaTfqZreroqtGFllXDEh2T94tf5fjX75M1zx3bOKTiucJsP
KsMrn6YTbhnwuC6ixVG4zr8k3DqfLilSWDwFdvmY6UhjEdRkm4ZOxDa7Eh1bpx1d
1JFDjR2YLA1z7IZsROTNc9E5n4jUbRzkN+X7Q2Xg4vU+0q/DyJzNyObRUGPc+qiP
8+dVEiei/ONqbxvangt0skI0dcjReUSbkrtnt/yz0VdbzQ8/wBilUSOWagHVYFDX
o1D9ANZ/Z2NnpPHOs9YhfVzj30oMHvo8oVHTabhRS6ZCCd48auxsl5b+wfOmAxDl
bKSzku6yuCcsPXC0WBWjgqoHpa5rGHKKmhWnX/KckMu25aprUDxQlKk+itVgJT25
KPufMEpvTnwK5B3IdkGGcV4aCGVDxDq7nZmGhPX2fN7KYHIYVfDONQ6qXXT6maaQ
7IZW+MRL4Yh2Dcr8Tvyx4bbiym8NhE7VeAmvNVj5OI9BfV1RpVzH/tejqx/1/FnJ
mzzz8HrN1/5ScIvNXSoXPSh+KvKJpUNKXrEKDn6geBHz5r0H7/QKryvEC9ZS4bnL
p6HQCh8zKWx5duRFye0gB+MOUhyRR0g9mgQcctjzv4rimRiBWh3LATp90hCYqPf7
jNOKTLEl0wQ4FKaNdflX/Hga65qWzY9vS3ataA0MzhX/V/MEnkChY2ijJ08fVFgP
UStS77dkUL68i72rxOs+wTkP/J85d6ihwYFaYdOqIog6/NUsIbOxWhLn82Uv43WK
baz9embpLCo8oxZyzDngCEtJuDtrV1m0NpQNb5oOe32hcg7TbwH6iCkWYMbmmPmU
3BpRQFWehHZ5YjzwYM0gmmzS+xopHnEPzCytXRQptpcmcC+ruJpiTg2XADUledGG
4ItxxhIv7nQnLVFRpnfsVscxP8WU3GJhVEyzSNlJOtUK9sxOlotn1L5M4QEjriyz
PRHoUHZG4qfd1VifGwGM74nkoIX2dNZQjBv+ERt2VgEOEIbymFl43ZvAjM+xbsHa
hKb2fwaSbRhKieg7lsKh4tjEG3V29zIdj20xiraHb8o2t+kX1CPPApjZf5KOyKtw
IrCb03Jda10UtyeaT4K6mNXuN3g+yJMoqzeYorv2ROzX2yiMfp/F2OK9X+qfwRVY
8mevl66o1B/TqNHdUZBF1bxlpTDaQoDEk4YlwlaNyz7LtI7matsW2vc3n32DA5bd
AlMgwAAjS1IFdGJCbQphDnQM96x0/DsnUTnose6p3dy0GzbH52NF6zZtoKulLTvC
1XPPByeiO/K9aXYPI/WjNTqkAcMqzNK3AD4a6AYioCwbfZCo3upDBlGcI9yPNIv3
iJdvSRK72v0X1WbDp5pnWZLtkKFGynU2YJYTYoaK5n6mARr4uQg/cTNWJv662xDV
ixricSJ7oSZFHDveHJcePpaZwcOsf2a66LRTmzDdkCE7SF1pkxEb1/+dqnHOw8DV
BPOdHW/d3bIE8dS8EE6X7Bp5xy31yC7VWJxftNUeCZH34QX5svWi9mI+duehQBM5
TFHKEJuib9MsbV0vc5551yKvnSumQ/Kit8MDL+hQZFJ69OxhgUUbRzNEtiG1yUmd
bpaSwBXTCvjXCGKXT12POJpGBIw4/VmkgnZvijTGlbHyh8FqM6+pOca4IUB1Gas0
Y/KKm3VQ4yE/d18MgSM1VrbgVSTSGr5nNwVeP1+yUIDFMHeMsaUh0J7vsMrQIXu4
jNXrgi2Cv0+Tkr0cpi3iMXoUymONG1Thz8904KkRd8Vgu3zpS2aUrkw/TO6t3tsY
Ysz1yDMqlC1ZCLa4rN1Dyitv6PmrAIRO3c6LrI/QxzZ+uAniQ1yx0DQ0HdTxU3SL
LYh0YKdt3JLDX4wP9izDNVWkf/O/CNswQM4MXjCmMU2ZfBssrcfijRUd+75aMmdk
s/LyYMRZhgeZzceSzfEcoDvZHQ+EiO8QsiptKMwa4f6lp/KO+Ney8D6AN4AuNmiL
IwD9jyChC/Tnp0K2QwxprEThLm+arAfwznTAv2DUROmYSRBNBz5ovgOJtXZAXb05
5IKCRri3ecv47DxJyXkiMmuxIqLvNYmv17RdtGVrwQHS9qV2p0yMD1c68a+5lI3H
Da4Yi3m7YEd2dRgZkHQmD/oYEg03o7GffCtDX9GY0Nfhe32CkspTEq8LlFkBv2n9
KNYD1xF8yGZcJO6QjkLGdXWsl8WjWyTKFScOW6kyQ6qahBT6ocgL14zd5Dj53QTx
d4F0NwCoqfeKCA87jpXMPTXeqNx0N8HKpwQssLy5zGDWTrmXZSynfgyzUsl4XsSS
PRU8D7ZAQs1+BGYpHszcCz85hp+FNEP8Fqlc5Rll7lumjIweHq29/bchrnPnFxlo
d4vRvFxgsGM1AWQaYTWkLyvJWvEb+ESud861natxzruSWAn8NUUpbZmoAAfBNhOJ
bHvYgzx7uSM5vgEF8nKwk5xPHW9JtOvhq5YqJ7Ts3YrqJXPfDPUCHJp3OMeKKvIU
etctau/01azAFxrNsK53aqfQpE5lhajxMgfKbY6s7pAV4xGs3Bsr1lyoa+KvVk7x
GUVp7iKf8fNRK21IQkPaRdgHTJV6XExKoYgKw4djIHicIMwRgsEViY588XelSY9Y
x1GXsCc/YIXlGc/Kqsv/Go0xUMzBgvLrgbxMIO6GMe1ozgP1QvXAJJUjwCqHZPbp
LimkMdgjCfN6ZioaLp0e+rjrwe5RVSaPiR/U1U5sRyt0wu0wKJnT8ZxdtcPD7uQj
sMCGzvfO4QjmPqJcakRjjoLph7iE0m9cKNZc/bxORWzAX6HeUwBfmChPPtIpR/oO
eO9AGHRKMcl9x1dHOowI/gyr2Ow0/BATAyvbjGsuxyzSH/GA8qKC/lcFPqPA9APS
WH7cEj/bbusIbokGtTOFutBR0L3w63lyXxDbnnh3Pkbq5ih4xZk0Y8TmOtRr6Qxe
lvgD3vaOrZxlLCBzUGnagvQpNZeWug1xEEMZjEsec307o8M03n5OCmCrN8bNF5VJ
demQ4l7WxpbxLAdwWH5Uj4SwOZD5yKalFFIoHzH5Qx/KA6F/2XImKfCncANoW0Lb
yDpSnLn7eI4I5UG+zjhnUSTrs9O0c+DgQGqArC4b9/lj8qBYLaanvNNHLDafFl73
S9IXSnn2Aai1uh6e7idZWVwD4HFSkaqTomw1tJz7J6IhRpxHuooTN35qlNLNsK8U
Lhn2fYppM7rTWzeG0unhUZy8oVTvrZhIQPXeVIxf4T0+EhbV1pVSGUPkzYrQU6MS
Ks6Xu/F1t3ndK3xQ0KZ2CpT8+Gun6PRdcQZ8a/XkbqNTfDsELBvWu3D3afGkorPt
b5ODievcX29NXS9z6HNOFbhSZTIa2A7WOf5HYajnhMPdtcorgBlGNvr1eqmoj7iT
GZ0Sdg3YtdLeDdz1+OYcC0X3lqirQ5WmTYQmocXuwVooopLIzOkzKU7bkyIwppLf
glWWwvKcKlXVlOWiMwIVulA4Sf/4w/QlDinK6Lsnh4NTlOji6orfZTuhnFPM+1Cs
L/PD7PB2Bbr2bz7CYbd1v5Y0J+7kKXDUHDFfeG1rkTGaJzNGj9hWpzG+yGNZ1pdX
YRUCvxCmYo88M8IZ46SMPep7PpOjlfCEy2ia+r2tHb9sCJLtPounlSim+3Jfk9Mh
/N9MSpI51yj/IXAsTurzy9hAnoUXimYiqtZq4A67pObBlEJdDJNSiSTwfO8vT9bb
Jmhsh3Bx3dKd+a6a0ba1k2OrrAMWVBQjX4SONBn/FDDuG+ldjvrV/90frXvlnKU0
4hVH/IoqglqXgXbwOHdufEejdU2/nirW+z0TJfBeq02Opn6SUsodw4CKNGxtpltQ
aJnNNh4YuLHJWHQ54EgQqM6zUxqf09fOMNS9issyA+A6yswmUV5EzkmZh3FCwo3r
xuI9WOi9G1UxIQg1aCtzdTwY2xVPsXVrHJR+OgNhExJNKzy+iJLp+2Cd+FPLjgGH
MklJGIcPi94LP9+ZylJRRO6b38F+UhNVXFu2DuY492+uQrTqgTBMw376jiSSp1qC
Zht/Z1MznHY6lPFk8UpLUM3P7vX2FMqFixgm2tH/EztKMEn75TLcLiZBr6WPmyuR
Et4BANkOrXgKDOi7lkLDHMXmAWkMEvlHUK89ycvpdv1V0YUIJhriSoEAffEHh+TU
YTTmO93415lQoH3K+nI0XohzHpZ9hSPKIU+3UiwnFsimqP5krbB5MqqnOeTgjdKO
noYtViUBDulIfdBrOzv2Q0zrVM24sfk3JhqUB2cDyOk+56+VUm2/ExpUftQdcLEt
G4Xas50MIVD9t3hxgF/HHto1U1QvU4A/YAC/KZ9gzlh6wMuV8bnQGGCb1ivKED5b
JH8Imody3uPcRXAkK/8TDbKGv8e7GgmbwYIWFGKQhI3bibjgTF6D1JGZ7/KxQhBc
RQn2Bbktm4teBtFh2tQBIhoCZElBhN0IiZCriw6sNH7R+ouwVU7QDj73P3r7Np5v
Bn5bDH8kDnJK8zQjyjxlEGM9haoQ2HON3eqpI4KadWpeXGFkfHHFqbGDk+uzJy6B
8M4O57tS5OxtNDY7bOwbpUjTIp3m0MSnk8N/UhUJZBNilqWp5FTV2Cyzuz8p+Uuf
apKgCqfhyLY0SaBh7PPq/NCVKiXMoG0BefWLM3Sd1cXUaVnGv/2YqbvdEbJAfJAp
PVMOVVrnBiL+YmrvV54J/WXPVaXr+XjNGFyFQgKSN1iQeYzwCBWtU+VrcAWIS9w0
UTbEKzx8Tux5SipMT4tfBHhOEf3JRkzTXizJRlDxnrNmsGbp1NBww85M2p/kU3Lo
l1ISrrqEtb6/3QDbMpef//rPEu5PbwwyhCVSJ8Yk39SpXy9mQLbg6iNXBUmOjfNz
qs3szE1SWLmWGmv34/yNWsthFrbItPDuGb7LoDt0YZ8d1l6tWXzthbRDixffcuX/
ojfHeL5BBljp4/NKGXqme17rlIBd4PmbYrC2kkbeWSPN71cPaZT0U8L/lq+Sjyew
KWD9R8epqxOsXo549Z/si+OcXOskToNww539LwPSqSatULpnq83v7u1b3TvUMlpk
eropA5Zk5bV0iHBv8uXMv/jw54TqAb49jF/VltgFZwwLHQ61av04JgognEnjUaba
fVVvKe9FfLXZ6mo8WmJ/CG8pefO5kq6aPxgwg5Bo/lKGy99Rl9SFrqt76rEpEp8e
T+SExS5R/JLKj1Cf6Excg6EG8Wiig5plEaOL76ZU+tQ7HyDM5Xx8y60wu+5rMrYz
gtkcmIpIe57oJAxQHfgQHzNqzWjgK1QL9TiVeCDQgeodpouxvU7y6SF7CC/3FaRk
2KD9Gk51/eq9jv53KYe87ZbS7llgLRZlI8LJWeshrMa3hJjcjTtN7y5wmR1W5DEe
Z8olR5iQx2qO7wAe0qjY0Y/noswMG6NFN7DmeoKjGTI3BRzDj8D6XnvtIMbz0ESS
67sjnAM+8u4/Hcqx4Fygd7oHw3cojD4jF3EEJV0x7xOdID9KFPTf7d/dv+CNdOnD
yB9zPtaO/vtUYbXAnDMOmttdCJ531uxfMnbqSZ5ZCsP1NlifnZpxIM3tiNjH7tTh
Ws1sOwjVjCeBvUG5vG6Dk0kVPcwhMFXvRd2OSbNvI0Z7diOzofavIuSVtCy3KUBY
BQfbElM7R5hLzcKWd74fRJ1aaNoMP+zYEwoy9Iij+AQlr5NNWhohOwGqWvyjEW6e
Jg+wV8GkHmvOffuxta9RLATx6ZeyIoa/iRjmucPiH/MLCi3nMqatYrDfuy9dwbUv
7+ehrJlZWr09VGKbUFxb15wIktTI0ixEbxSqERE7s6VeVjITiCiTqfjymBQm0KNg
TEOTtOIkxbDKfSNFO0hfgC7tzkOrynSMeFtyXEYx5WTU2p710bdMURBam6MSadSP
UCsa92aQR2dXOVzCQXYCKvHVuMVBdwyvQynorxHb8FbbO7CEZ50RHNEc8RXGRF6M
nyaAffqaosCNks5ZjRB9OdVmY/Uw5BdZFVUSC0pw4yTN/yxI1OooZRoDIzR1BbM+
MQWpqtnyW5X6AqDedolzZyMeqoMS92wPCLQqGYApVgD0zQ9Nvg3OUK9SIgw3hrkA
c9z5vyuSZNCPEaU4vGAQtyZPNMWcrcJv9f+0QowHHQgS0B+/MVrhyQvLlY/ESUXl
0jN20+jtWfCTCjGtRvDduf1EaWrdLyGyMi1qiuJQF0odic6pv7vl5NhQ4D+pDvbO
zc9yXASqRD94rCDv0JxzJSZF63sQRX6gpkstyeZCU4Jk2eVUmTWKjoGf3da6Uewq
reYUIO8qxMsqwLAaGtfXZMrsRKQO2rb0nzci/fjdVBG97m1ALJNioqseAUzuk6Jj
xez2wkP4f/Xg08p3P9ecv1yMCRBCfFZxAksc9FGFhvs7dhoJAalgGZ2FUJtkqSJx
vR8iiT4yXAcnXfICPrHIBQt01vJ0gl09VV4foUn2c280bPX1nFJWTobJgvqFd1Az
YqolBZnIcV8CUHkHHDocakCX92v2vwwgJPmhGQjKJlA5Qkfk4ClOVpNTinF88wdr
c6lfHYbv8CW35M2Na5vYBikLI1TADI0GZSSpDEnx/RsYCrAyfRrfI49PEghesTLt
jQwYtcU0nZaANaDA62/K8hRvXk8jejAgCm9+IdeCUcM8V3ifAmBpDbxNFJasev0K
mzbhTiW/SHVv1XvsjL/TdYG49goVoK5GzU80Akf67RLk3cbYGEn+Udeb6aVqg3Vi
JIZT2+f40+trpm/8bceI/SSaaVJMJ7JI/wp7ewZ1uPHWlinA0GOBqPWFurXMf6kP
8YQIEfR0C9WkvKXKS82eQAXJf3xKtbXCX6r6hQ4r1rfSomXmab1R93CdDXCLAfmw
+S/vNJHldx32+ouRG6tCJ6zoVboM/AMcgggxR2M3LZsjOXT9ByQUrrayiw41OIuO
wXl+8iK5lrPQ41h1zejMbuLvSfhij3xqXjb13Y8IhsndqRgwIDYJKAyMbJyX1aoy
Lt/5uUMIxLWOiguvAfdbwdhBS76Tu7o044ishilDycUe0PCIzVr3utWdvPaHOz+V
ydvf64eUocAAqrWQ2zjqZym3NMvYoM/MCZwwwsSmlE5ypmQqembWJQY3Tdlvo4GV
041NP5sBtramSuSxxuIAyK2cIBhbsXJFXrRWHh/jhTESX2O75liY1VaKMT5f3qzP
tQZphzeknj5erurT1SUgtaahTfxJ6IUJmVWg3rccUT4KVWNjXmDa2/9/p/oT2z+0
Zx+zcflPTCAZ/MWKS52FUSPcdmYGmP5gtwCmEMNGLwjFPMkmIw30gvQ9pRVjsuNO
ODIzMoZrgDW6wyhOkqzUKmeJU/25fvK2c7SteS/a/uDW4WhiGogA9/JdhqBc8Kmy
SblA4v3oI+yXbuSBLtPBAQzP+FFZX1U0KNvXzBzVoS7a9Ygp6Yz8xc6z8Ogll0NN
ahz7t3tNalhBMOzPxXdPam4BuYyZICkv/2P+xUL8/oNmxDNeksfqhXF4z4nsvM0l
7mVDnAwHWcto4qwNwlc6WkfKm3ypXFYAk8rTa/XNVaT1JD41X3k9vimh4i2rr4+m
w7sNIxyUseiOGhgCSMdvxEcPnN8eVhucuw2IXtTVUFoHZsmdPOsrQFsVaMA5x3iT
Ux/oVKoOXSXhRMlagAJP2Uuii9wfNK6N4M7glS0wS8+Q9WQLiVfPaquipnb6f+SB
xcVnv5x719hQY+o5CatxX2MX1bRKhX92XXo1HJB1liPIj39V+PJ6VQiK59pmd/Dm
tYeSD3CbFeeR/8VvA4tZ4Y3B0QG0LwzFOK2jYQE2VwiGz9l/6J3UQ4wba8uhxPbX
+wcbVycYK5wIYTMxSC4BJDdvtCGw9PhC1OrHNYDS6TZJjcHAax2w2RdS5/B76JkI
qLZRKS8MuLaeJfo2WS5jv4aoi1smmJcjf8XSnE9gO3r0Vtnmyu4DuqFavM8K5cxd
yjkJYSKSNsOA3h4qlupe+M+T59gck6hOs/CZxxsPce4MmvkgnFIY1AvCD4h/I6uW
rwG3OXY29e0VvLCc+v4GZNEe7h/msfMejY4bhiTHyOanck0bUaGjpaHGEYAPjqT0
JxaE1J8q08V5uRoHI9wb8A4KKIkqBYio2E6SLvT6jxsSQYRgcUPTeNyRCSI4slJu
tpSHNxvKpuSHs1O+KT+EHk8oQWCFY2BWdOGM3FAy1shXaYEDDEci6if5u8+gPgt1
gk/Z2rEonoQgW55t8rBAnNQF/EEFgNmagQNTyoVbyIHxZEHQm6Mr430b7HFNF737
8I9rpZU65wd1SiH8SpiJI91KK/RHWRTKddWl6YiEXg2Nnr9VMgvy5TAeShSBbC+1
p1i9aue2k3J/4rwEyyukFPg7+sgKuW2Apxt3CHmlorPLjfknYC5iCmSLKy6jtC9z
mxW3hSKdwiNo986tbsbNYfgZe7JrjS45p628weBZgTGbB83rKKiCCNdG9X2TBbqe
rJ26qcmtRIhoLuHoGM9tt0VJl4b6N1kXwyHZ6WOwmC0n8XUJZoniMv+cIrhm7CrF
Fg0hrKQfI65GdsZWZTbxCNzRhGo9ttKfoyU/kUIrlCJIw0+QIlEOwlt8uCuVyC7C
amcOXbFQK58CjXad0lwpFhhtA8dbp1AqZj524GJcbEFSPtgAf2jv+d6uMoYsbqFI
zS+QWeyA7cmea5wsq/cbZlHxfEe6J7jvA5l06arw8qvPj7NNQtsmM6acdxsnbpbX
FKyQPpRLQ2vYPmAHtft3YpYGG6ZSjnL1EzQb3lu6AupsdVvHmFqxeEHQQVBVlXn6
9Np7xx1Vddv2xMJmkXi71BJFVOe9O2AJ7PatteBwMHC32qohKj1Rixa3/zSCUSDO
2vDZzROOz2Bb0nGJnQtwmKsGq3R4gOQsJ52c6dUTEVUm56/xgVscotZ3J5j+cBqG
jN2liyv6+kX7GRaGVAPRNdrEGdaV1kh8uev/+Ga8a4VSOllEc0g+oY1EPW0iqcba
jCL0OkrMK7XUGK4zs5kV2hCYc54i2jA3vq5DRxBPrZIUUYUBCIT113273Ys6HBdN
0dyIAAsaMRVOWHHrgvydQ0AYsbgjHuZgTGoyv0Fn7OuykvCvBaoIY0ocYYRyGBE2
DJKQfiRBk4M45n4AtIbBE15U3/HUzGOdlsyVorqdz27Q8J66hoENg8MBmp3Y3gLF
uGvaMxdJ4lXgM6pTLCeWzTbuI+rDszv80lzsk7bxUm7lu10NzVEGK1rlVB/sINo9
oqDMSf2IQKK6Iftbq1KeSP3xrOfafxNzVFqg1MepZtOWAMLHurGkcGRurF9MxQGr
VaWTrDG+pTQYCZ2cY3WhmOlnTetKOM3UYMjln6GvBe6krV9MuX3xA5THwQylukaz
PPMSjrX3gWhHWgBtToEADS1059OzVYZDWbnv2w+FQkIx4twhPvptMJPz8ufNy6fA
uqEI0dW0KgdaxzKFEoJZML4zhev8aJuN0r1IUVhF5wx3lgebk2zLUhae5im5E+Pu
XbwmSCivjOrCxBE2JZ5C4eY/T6AJoJTpaORsfdqU7mSQDidYwfaGT9XJ4tk94JFB
0A6bSMTRj4YvQyBrWJrOHlgcsddZxaN0XWOuVur7CtzVcyfrOcwOrRet2hLVCsM0
Hw4qXffn5jlN4sJP+0fzACOUP44hY39fr/ED/4xKfT5Tyjqn2QeIZ3S3pjPqj0R/
dspbhBQpnGyqZPYwZQYzhxu08n8njRT7QfW6eusqqiZajthNq4+Uopor66T/eE83
FoeM2947/q0xX617RmiVXVYHHAH2n9nSvQz+DB5WlLAxH8KrK4Zh0DqyiOPJ02rU
IM2pZ8jWwP9DQ+z0NQSOzA2w/qJUoPKx2BlyEyCINd6B1NHU8flT5BVArXonSl0G
Y19pEow0y2lF3pa7e1/99LaXxbYWixw2a9BoPi+ZGeqrE/TGvDIGDbmKT7OO6Zy+
6hPdshUqQ+MpZxg9Qm+EDNdna4e2shbNh7C4KyTyOeMiSl8tk61aztfqIQh4ET/I
sD0YMKYc6EXTYCKxPw1RTBilJYKqtlxMofkNOot4HupK/JKbbA7VrYb0E+pqA6Vm
0yhtet038njpTDkzp1TSOKzVj6p4zUYXPMmv1lpeg/cwF509iFZ0DOovwKmVcAP+
tFFPHIbON2Q6t/zEv7DjGKXoiRl/JHLyhntuPzGcbnd4/AvizOQ/JBCfgNhEnV6W
BCJNoFMWRpckP2kdtV7WSDGNYoz+TyJBMZmrE+GF2m80n6JTNmE6Y5nEzfzraK0B
R1uI0+JDs7KsWlKw0KLwuzjkWwzekL3j7VKGZ3KgKUjFvQMnzF+gQgGI6pZmCxbm
TmCnH43C0viIhP4x4Oh/YZyAF01tGa6wwlLPk7A2RJwQ+hMgJK/11n4J+Gv7D+oS
iBaI/HsIhShBKcewgBcjxT7bARkqfwOrnZP5Wyg13TnEvnhqURPck/PQEdyw6kCE
JBfmYMLp7EIMPjwVX0mgZUn32d/1XCPMNA5JAICzgLa95XeawDfyBBdufSUewqiI
9lUQIdSYbLbicnrkE/7qGyNI26RPYRbPKGO48qRw3eJK17UEnZxO2fC57zM53zpj
QzrR43kp65FXH7Ugdmo0FP7Og99X9f2FWuzvPlv0Hcb/OIT7kQVEY+vNvuN6kWmx
0GcH4oKndIGelDeGtPPvywKNNjOAjErtT6VLiXnZ0odzVmLP5IvYDxaRGFBfSF1E
OYJWqcS3ucR6pPhWz8zIZiM29clOPR8PNuhjNZb0LHa7TSot5i1xzBew7xIfiU9V
XYm7YH0jMwjjjma6BFgSHVo2jv0Qxrou2HtU3OwWzrgRCtB1/alZXrdCBsEVmZF1
L1S76+yKR1A7u6jnUo2/5oRDbh13LYoNmEYHcg7XAZnk4UWR7R7yi7tlN6eTc1Zs
yEu0Ic58Lr2RaEKPQzpCBqADlWEdc/4lVcYV2SzKBiU+LHPDm1mTvs/qr/59HbH1
ZDIvHUfTXQ2ZwdUaWCH9L5I2L+jy3QSyex8qcsJ0LkOpseJpCWWpihK/JZA1e9lK
iuPt5e0TMY2piPN6hKdUlzXtAss9OjCBpHKiyh1tyTKqSefXz7JrpQWYyTnP/TVY
nhDLsFN2UkZMB/ZhbzicKWKAmuaL/2naB1q0l+gvfZQL55rMsHvHRDGnfTBN9Q2I
rQJnyIhAGGWEpTD2gp6wFx1G3LDMMEHWFzLN322h79+9fCjgZlkNHYKgZh4Th3u5
koOoKcSBGTVJSjcgzdH48nA0WtOsmD/FTeWudSPVXrpUVWqzb+XFxlJCbixgguOD
vczAoCJedPzAjgIoCcsuWhkC7zUqN2cn//FNKMaF91pjQUqAnbs7qZyZmkIgnVIv
SknGWz8epvJh//sXzfEEXZGhYxS6Hq9wu9G8r04QBRxviAq2Y62hMhQqrvms409m
JatxD70wl28AjvaOUMtrAmTTGKGsE2tbbmHYwAYi51yUn30kp1Ka7ZJaijKs92er
OzFWijKUPB7f937Zo0ZKOv6jvtFa6xr37CHLUol/F59MiyCGnVsjEhnsaQzUONDa
23+iOAGCJpAA5HT3rokDPGPDMS7GFqT9qT8Uw+PCpMXyB/ZkdDohQJXmmmYuuX9U
N75JjJ9tS8FR073qPlElWhvQ07GnujT0KCuoOB8AJwNNzhYJfSdd27PpxRQzIN3r
pUy8y3YcZuFCBwr9Q1IESKm9XER//qLXpZ7NA9eD5CKCHpOIHF4V50TvUqDByzIe
tnHW2sp4Q70EuV1BJncf1e1875+HBYxpZFnLHA/mHgyCPH1+fcwJj0Rjqu6xiSRi
FhekXzk5gb1cZePaVhG2q6QZT5fKkV9Qgx/Ej0EoGddj4BQrWkgPgtI4qgsS8Ivu
pLmUQrvPm7hpAuCmwzkjIlAkwEc8UH13lq4w/S+3bQ3wdVJ8MhKodyXty2uMiXyY
V0D6EpxyoXzE3VbRMOcWn0eLC38Jdp5DbxkYbJboTwb5C/6EDRgT1g6giQYsBDoP
GZWj2z8ph94hvlcssuF3uBj2nO51bBMZXtARkmaTMk29k8bhIkHwdbyNthxE7gXK
GKLX2RNoOxx+Vmyv7WBKpcO2SxJ5aiKiRxo4F5nxSIs1kxvduYmKCpgIUEoTaJVS
zNEKjS9zYCRr43Dt7famBz9UiVbo6WFq7/mR/w8nBof0YXqqaUvJkwa7skx6KBsG
6YdhR7uOu0K2msfklo/mRuVES3pB4sjRvSyYBT8fAfwkY4vCGKCYxtjMN+Lc85Xf
yND9f/oKxKMyI7dwgRYpZrE3JXKn8Wc6Wg3XDUOoL3GrR9bbvrdr4r7YPaRRioY9
98oY+3UQnMq70PneufMudrF6gxjn2sQkTK/3/HBAKM5dNh885MvdeBnG60YgfZhr
/svf0qkWmiKSrCrogN9U5UUDM2t3Gq2BcjhAriPB3idqQkM/5GKOFzQDYNAkaBhk
CY/KInfgQK3/OT3cFKFQJ5yfdeMA60lXjCLS3m84AJrbAXZ7v2DgyLZ4g3oMWRnn
8bnrUDZAP6OZrj8wcXSE2AupqKEbnbjmflgDGu6rlML9xqBqZV+G7MoNi28zwcQQ
CehGJcXFZ00P3soiatqudfu4kz5g0/arr7EHO6OiCa4zUXuSGytt+nqUU30nqcZT
I7z1IKWgwl40QSS/BICrV8JTfBPpxw/aBIO40ATXVeIIUukbDgvknhbER43+c2ia
VPVFkmOh9/Zche75f0gqh9AulIvD6kmOZZ1V5ajX27wjvxjJScIyIhXmeryopUAH
JG2MDyX1KGIZ0fxQWW9ODMKGNTJ28IVby2gY3jTTpi8vRWjW7gv17LbS7/8e5zIM
7r9IB8pWAAQWRKaOObX6Zz9BQyXFWZLnF8Bsu/Pm/kTHNs/fnJeINc/sEgmo/tXe
zCqPevFP7RtJthP+In+Sii+PIdDF+ZLv/ufWPIKZs2gAa9FmyIVhk0nzOy8yaaFf
7vMBXR5xF4zFwMYWf4oWoUBJ8Z7sMgwSg3gRmZ9OmYsgPK4sLI6cBY032DpyBQsh
zXoWXjyfppypzwEQHCKNp56Kbl0QxHqbbTpeAan4kMiCIizuLVu4hSLT1v4fvdqq
Rr+Db5/UxpPa2Dgyf3UJFo/RbaMsVUr8ZGJ/1xN8vwDIMrH56AdS4YE6WaTH7GoL
3mnw7BOwzx3OahqwoZbVrK1vT0g8iEHdkCsPxqaLSblFs/5MNliH4cJ90a9UiMRj
9on1NqXHHflDqHUyg/J478k62kzkVMsqViVluzdMyGGFECqf83z/0ovgooiYbxOd
xbnGOZLrcKPbWWzlIob02yJ/xqUatr0c80BEwu+vV1C/Lkr1qxU/8AOoH9qfag7W
i5BKsNibmHc1SutXG4CveGZaYSNELzXB8WrVs/eJZk0XdchZV3oaD4dNnPgQiYtg
6Od3AFGEcDyU8SvrtCfla4zcUTQ3judZOrg4OgpeqZQeEZ9jVpP/F4ax6sRmJ2Ga
MnJGQishVSaiC+yoEQjfVcaohtP59i1tHv1ScsWDaz4hmZzFZ+AUzeUQIkNCvzBw
nWRDy1pDeFyX+iITfQRLvtP7zE728EI096T+G2+aiLWPO15PGTimAGKRyp6U03vS
zgkjvR3yZITosgh8ppE+Eb4gtufzp4ihlJ3CI5ip4p14dic1u20g3mwHpzvom40X
A8E3FwlaC0Zohk6/agZPR/gg9vKnnUIoFb24dhFx4FHoTFIAX76CRM+cpEEVlF+s
KhwhaEUczogXpkRsLOwgMJQqmjxrpILMBeQm8z/RHpR79Mw9nHUY6uDxhRlwiHoB
2nivdZ3a8f3aelaije8EWtfHWTpj8axP2lPifITgXseKBXgf4n9vZBPGSuso2gA3
7QoRZbkWP3uHZ6WpDqPzwwEPCG3BFCS5KaSg4GhQUOlYLRUAYhQDJS2NcUsEhT48
J0wHKmCqxNxgB9SntipjzlsA317/HMXs7F+ZCRHgaAI3gYOM+vLxVWb4+y1+7YnN
uuZ4S6VGDDXcnBEXNW/8sYavTQorWLKLI/zvaYpo3NXc1AHbtT6JhdPGHTnS1PmD
CAs1zRP3mJBhw/C+kb55n7FBF/WypnYicb6JD5eXbSMvZHpu80jhjPZ+/pVjTEkK
i3F2YsXPqfHylryYm5PD4ow/xjHjZtfXYR9MPIYMRLHJHmZxWJ53BBza0cz4Xt4V
Qgtysx1B7nrsNfYbp/C0Wg3ZUO40HD3tdsdUt3mYESlJ3ye/gxaph0PUsBJ+F6Gr
gHx6r7BogQ9rB1s15Lss7T4ZddI7daa2FZkorQSE94cYO/1dUXORj7QTCEZJeERD
P8v2NgVIcEdRCq30kBkTGQnKhy0EX72Iqo1WyAYlseQJ8yntp2HhfUONOu0cdzxO
TJ0T8t0z1y1pzKJYDCcJgsSGXm2FQg1tJKnyaqPUgNuUuNIjTKxV8gPrI6YFhleg
4w+843kMPtMl6WCTV7WZz8qEQ5afq2A9vMNunLuxpR1P5IRToTNpoRr2iXGe3Hko
jhVoHUFVUBI+RuE4v6f65DQnFqrWPKE7lu476POM0yAaQ2vo2sAdG6jOJQzW1xBr
DFpayq0xD5x2Mwt3ZL8Gxj6wq5aA011LE52ljzQpKiE3iqcEDuTp7dmJdEdpvpM/
7wZ6L07DJNmazONKOnG/AoHLfh3QTjGQ37tQZFIimBX2iESIQ3p4TuQMXrA400vN
oRlSNbLgp20sKSoYNXiPMKxacyaP1OdQfOQaXXOf3+B2El1yOaNFssRvn2lteCrw
V0aidSL4HYpsZHZr8bFFpZ1Axd938fb6FeIbwmcP2QwOTEEzZhfZQLVu4OzQsQUa
2kSaPAfMKHwbRMQI7vV1c4AdKuuufGdYp2uIR0rJAGcE4M3tgwQIVPbTVGM0+nH+
Sr9juGmzCDAJJTEDBtLf9I9/meHStQ8iExrq24pua20MVlW3wWBAv+9v6rPviGsp
kEd4f3wxWEPJXpghyigWkKltKWQSIMfbc0CbKckO/4hil7sly5BvIVNv5fsB/m5e
ezTaHVnLKp1rKpWh8LytmSNxHQjLmD9F98mLX/+2k9sJ+2AgAmF+eu3hbh8gSFFr
6PtKFDzDpzq+cEK7Y/hy+lWKwUfFlBTxcEf1vga3cHzeabFJulaDGOp8zIjsO43j
jG26FHbgYcetnjs5mE98ioHGyvcHmP1hMBnDWPJaGJXebJU+0yqA0MxpdtXqAUXd
7SBQVlaVIvlugoLHYPcLahL2eo6vyHUWdIqhh6T38tRLvlr+XX2GklOVcbgDbk7r
8ha0giEHyR2somrR0+Hk+10eTQO9Ch9EabKPpgw+1q+7vazT8c22Y+aL6+BczG0X
gmVi5UJf5thFGcptnknUH9ikjtkdBnwUQF/ZOBytJR1fFUciyP+Op5hNUXCqdXtW
GnCwaYnqNc2MKS4wVfawKIKT+pOgq9LC78QNR28YMdrecmqEM4UR0TYLLSVkzXYa
+HdUfzS90Xanzupi3t0zVFx9dZy1WireRgTo3etlaP3+CzyubR0QFQ2Z5TGHzh1B
Wm4FhlPON12p6F5WbWSArnCRSGxktYvnvPKYhQ7Cpul9capH64oJ4w4Kmv1GmMxF
bWdC+aOZ8HdhUhLpeDnmRrJgf1NEI5pRstmog7XgICAU/YzcgPw9UcmQz9L3Qhdl
fvrox7qaSjRx+ZF2j58eXBm9GOXhFcQZzeqO6StiMyBhYiVvemRDyUQ5MdW0+21k
iTTwGg21HDidKXIB0+rG2rLT4DQyGmcLe2muLpUdV7YzZFR0Y09lJWTRCOojx9rs
kiZizBJzaHoksfI4r4pTYaFNC5tNLxi48JXmr/0lRivtTBDkF97zwVLCiUANb5Fk
d/pfSjvkLeUAVBKzZWkVlHM7agCfwX6s7opqP9DsaQFd68aS/hJ0JNRp0ktkN3W8
xG2RaRTtdbGgaSPlViv7zxNk8SauABwt5WhG9+2dCufwzoMnqTvsnoVIaS5l3+W1
Sg/xpK8NFq3guQTMl7hJZU4w1348NUZbF8K1DuTF9QTdcGnaZBh8yfzUCbvfTiKa
tj22K2krwN/elLWZrG6s05FMOdpzU/GkMzMOlKoe/kW8xYOZ5q0ilv1dLQatjpyY
A1YP1laWdiPhjvCwZxmKCG31hNsh2YSwNR4QYpHhMeN3fZ9ozZBfY3fGQOKArLP8
7F6Z/Xguqbdr6OcHCbQfvzoc30f9Yh2dDqyZMqH/hGmWYNTzLeK/UdSsbDz+cGHS
E6G75cmF5Bq8M50k76pqrB3x+D7KShb6AcBLEEWPOGw9zLfeBYXY0K8pUJ111eZj
DiTjEDbjDnmFipqx1XE8htX40p+6j6Tiq3rBPYoLffsvuQy7WoOsxMChiRagw0tj
UJVe5HU3RjRyAuonOuPei9Rzus8v1QHWG3CFtcpa26NJahz3E5zB4X5uZb+jqkRP
yklgAQJznvf853/aZJXNqqCCTJ9wAmuxV/zSvQ8D8lxn1PjUVIS1GSlTuQHSa8Kn
r2+Q2tJNjWYwDjjr+SYRXbXXAI6j8AZ8zthrQ/Kl52umfAQ8Bf/Du9An/a5l8uLn
WtO7taU4l/zFlERMlK8i4l9+2HsBldZYEYwsd7/+Z1glJXlILljgbSY8L9QOr6iP
/nnLeNBa/KfjBrEi3tl/kdDpw0incAY52a9dWCZDcjo8QXQAOmMcNLO9QhLrd2qj
M3quIpMxKLhAbGx4Huiyd0LuthX7OcJsjgCABWqltCnRUPOuBB87YvrTz/0fXR8Q
uLFUJYIJxzouRRXNGo1dMH6tG2zVwn2qedgavXleCr8U8TV/8Nex0R+w7ILfq1Zd
Gj8ypp9TnETGpA5cj7TL7les5bXdRI+ayugaixprfxyqHFxsT+snjHDbC+Co9Xtl
k3TKNuSGKk2c/tDF7pPydodN1vUyfoVdxIAFcHgxtwcLkPpuUSCgs4xl67a18y3r
lhWmMt+ZvyehE9D3ugYuY/WeF++QrpwhFo1PMkcpkz6rw5qc7idw0VTbuRkZMKPD
74W71UqOaDtiOoc8KboNuwu61M57/Hb6J+bxU0WxDHwbZiuQWWK034O9CbnDYzFA
XCz7C8rQXv762Uwwfuieg1xchOmXW3uID2k4onbPQ5VoGYC4P4sjIq5SUphpuTQW
+oLwnhBi+69fSdb53NVe0jr58aAjtNw8t9+YWYts06IJHcgUnTASdkqpgjvMlKYw
tundme2WntuP+aLMTlPdNiqmmjgWOwfXfpiL6Dsiv4RRtbVu2B52EfCbIgTh0Owg
UsA7D1tFwhHdnLeJncCrNkDtasrBAS033Ej9fFCltpavNOh3i6wakjC2rNM+pkUN
k3Fg7KyGtVyWH/yXfXWo7QtWPgGJ5DwnHC/sSlRV7/IXWctWu5meBKrVPs1NplNx
A2BHertHTRVVK3dlba2Lnq0iPHmkM0W+zNvjkFF/J0mKi2r2M4urvqVIG2T/ytQl
4il2KpcUv1eA37sEkirExjcK+nf09qGvTdtCnWajZEyY3D3iis0rkUlpnEdKpgqP
95k0O+45e6uV7o9icC7C+LIAiX9znantpywluPScG7btG5pUaTDuuWyj9zT+dUQB
HQip9mQIrsh2MRR9CrbIs0VLfzVjoY40A/cJgQg4zqdA/FmD1hbwdGZ+MWNihTJQ
AM1Nxnfycx8kpa2kdrPxxr7VarVZi4uSLWCao71lzqq7UBGw7tJttzDeJ1T24p6O
q22J435t17rNJVCA9+g0VaR2PulQkCySeUp+oXejYAme9DQihtl5bYMufyWC76is
0mUEuQObYIGVNzBujJJ/PoCfh+TS9yJ7sJ/8XKiyXEXfPreivlOztjBA+xENu34C
fjTobffi6fGTzyLze63A82MYsDDlN+3e9Kp+npUsAipsQvQ2UpdP9EDoNY940VLH
hUNHDhylHjZiW8VAj9JrehY4kjEJ3TxE+kgKhbo9za5PbLwp9wn5N5xGnHUSgOZL
D2CbknznXis8kMlh4fq17m+7mjpna5dYfzdRkVZH5NoXZLNW39rypb6020+YnK2g
WVgdHenqeW0dY+hBHXWQRzU87ONbORtrrbRxwm8ROGGKxuV5l+dYq59j7mgne2JP
3dEXOq++UAJNJDOTR25Nxa1tcqielB9ebE16QRKBZds1IqfRU7+EC2yfSSbWtAMV
U1YY46lzoJfhFLp8QO8iu5bpNSpgvkM5b3V8qqBlF8J4k7MgSatvGeM07xRv2ilx
vt/jhuZ6P/4aBhIoI/roVQJM7vHEotgomdt+auHLtrPcZ0R7l6JjRsN+Bvd8bfOY
nOmHWYzDxa8z/fqFEVauv1hPNE2JVWIEsyq6WpxnfQ0loSE6sfmGhTZKcQk12hco
e/9fC2u2dZ7O+HtN622T4r/xAnACk2SDfZS+scLxto8N7tOdR/eACUpb2fNJVr6e
e3wabts1gdDXIN6W+fStkxUxe/6i7ZRh9QyyPNujDEKkyHrHwUrB7Gct03bYDWAG
VJ/kOeOz8FbnmLexmC80H81ObBZpGwFQl3t15tNBVpM2gtVHeOSMzs0qhUR0oUHl
h4U/O+PtAVAjjX371PJeW9m8MGj4EMYwvj+34s3F5cKAynUCOw/tPAODn4nv/hsX
BJc7qZObmOdlJ0nOEtTsuwPWGeG4oxvzhThrv1BMrR0bGiUrRLsEmg4GbrDAqgDU
+mPSaM3YF1c7caeJCjLFzOKskQlJLj2SjmteV0B6t0AcBka7dTkmVN3SiGbDV1tW
ooKYfyGRWbEl32K4D3quRf4ivcO1dJdl1sIvNoUoB/RurFj6gLd2vmf7n4WI6SeJ
xOp81MR8eWvWRaLBiKUigv+RF2XTphHJ8rjEixPUvKPLctyt3atXJy0EjutNeyOI
YaLIXlwp9sEInR21TRyu9Lno3wFGOZJDXbxAgr2rJdjl/UCs7lDlbGnl8qVHd5m3
frTuAQD9N54lsJmGY2F9MYAktvm/K8iQnEGB3HLW+FgBYHu+yWBLJ/cLXIm/+3y9
fCIMN4YTFTuaz3fS1tnq/UuEbbSBXzncBNf/UEN+zwTm2s3OpPuBMub00aJXtm0I
RhuScfljUk20ytJrCz55xvXhrYkCzgX39EIhHnwfIsqPU9vlKfM7YWoN+2sYfDTu
Wj83W1u1V+mc2CDKOB1nKhqm0xk8U8TrYYJuCssSdmYjwKf56F1XRzvuvV7RbZ7T
bxPhiIq1W8RF9CLUsJmbRnn73n/RRjN7/FqNwV6aPuic+lqNrwtZCCM8DotqdNWj
URoxlgtHQw6+UIgNCT79zK8jZ6jOQQog6oxlVzC6X1VKVQnkJAwFL2rlLGkYMBf3
gI/jImITl5ql3Kn/KCEaPDN43p3mc1GbANoGhSCZlG5cdLMJpTnltkwAKiIhusVU
ftKi0rUWIUbHg13ENDh5L4j8fjRwNbuJCI04N45uSE/2IQgizz20uChHYiB1oHc8
6US4EXKfOCW3e5ctMXrnYmhle316kh6xnLifSowLERAsWfH4bv4MUHWKjISUIN6c
ASvv9LUazVxUS3jbbPfC9UDnhjXCRYOh/desBylDGKlh5pHfuYB8gxWNhppp0jgt
FTHT8HXb2yeAo3xv87DC3ywmQ7Zd9aaZMDA4UofSyivIhoLXyFapW2xC15GJbdW1
2t5KQKJQBRP1qncxNVnKeUJfzgmj+QPR+Z1/vnWEXJbysh5XjVKnebw/v6bdb2Wy
qD8bbBodskVH5CN7Ol+2bA9ji40LlQGbsww7dliyFi1gQiFngAMNxfrMgqnD8NjN
rKKE0hmtSG81O7YxEutTaDLw9e9Yr3iM2QeSbI2ciyCrfbWvDHMn+qSKTkLIaOuV
lyOxTtYEqi6CQZtWFkjCtay6+WUQ8kAGL/4lQb62CTXmizQmZgh7IIVf7VAZj+/U
CRGfusz8yrmMj83gtOMbHFhxmkMqZ6Ykfx2N2xZ+5nb2aKIhsZOJppeMq2CsYYr2
/40MDWO72fAli+a5cVBwTQggevlmQG0hUKwRfiIO8Dq2UQ5UcU6pdTrRq/wbItkh
r3r8f3D5XR+jMkhLJbMy2tRvfmPnZ+SXTncq8ykh7Uczotp9Em9TR9dhx+oEv04F
leOuYpNmXG36o7mbkzmWynvVuwf7z6EDn5uc2vDbsQR/naxwMrGZ++aRS7XqrIr6
9TMhkBDJxq+02hrsFfPfi1tQ3NcLVQjdGDwGaZBmYTOmd539i35tHtADv+szbdQM
Ocz4lAorGIfG4PM8bfQuwqWetkNuc2fUxxzJtv60qbKWKKnEXfSQcWc2KxZ9jy4L
ct4kYTEYAxlV3KzQcjtTZQpU/UffxX6KMr11WTgYBVdu8RpZBwp0ecv/14BSzCOo
Pgnkq8zXje79KptDM4RES2BeIRBcQFDsSVjCWkM/RKWEyShBx8PPGVX586EhJkdN
U9E9UMTlRLpyVYZjEJLDGT2xMjL0py2bco0ncG6fWPcvVfFsaK+6J+N7dz6FSIf5
NlkGzJxUj8N7BTwx1xQHAI1FSKBhX0t/9FVC4ywaDn2xSQ3lZ/UUDLs4X5HJJVan
oIJSGmjf8lvy406bI3baRvOzwKDQ+zmq28BdHokFz/XOtcNinRIdiBeUlEf/tHSA
pdMjtkQ0fIo86DjU7wGNC4nupW/YDvBWK3iLFwLDgSutVjgaFDz3Vtygi3O7cqNg
sUD9WRrvOX6PcuYm9AisYWKbRqD2n+h2tTbBD7hqsaYn0lDUjitjmeDA4h9DUYTM
DoSzxpIRkj/f07fzt61ZGAenCoZZzePWIvQh7pzxe7iy2rCD1iyVeY1N7wGljkHR
4Be64QrYZdX67wjtQv0WACcYnYXhg4IS6qWi70aMeaGCR4EC5GRM5uHPLEcZzTkh
ILgrenFKIT0fQPypVfdWZ5XZFxYX724hvRDy2+s2jb968eo1/+bMDnzp2v5ZO9AK
xmcHGMzUHUeBLwxQBnrkmScKEGm2Yw1sFtdfIsfnK/RyvtguogJZaUiM9Z1Qxi0r
qI5aznQoqUvT7GLJ5jW6WoIKzrkTCVaqodKZIkFBw0/IA6pHxQ6oK9vaUHiO3H0u
ev1vKUp27VhuYrVlIkDnaO3t/oFW0483iaJCZ0g1V5mNZcyX6Z7cyGVIUhc4Mi2K
iyvGKf4UfhAdLbPhmRozaF+0wCxsCMBv06X6OS+JLZOjvt+mRcip7++P9K90Zxv0
66is8/5zIIh/u9k5HUkVohKc4QtG4MJ9qZuvTiJ6U408CSGnDGiHGFGa6MkwcOlZ
ykQBYOJzE1FS9eE2aFzryaZn8BADVnpOiJR7kX+cyJxDxJRWByN7DObgg7J3douL
QTCbhGSU6buPnnWJpfvVGKbDKDCSw34AMhDqiQorJDDpA50LsgX5FO0SQ63lYOOw
GdfmjMzYzUOFzSBH2bEBjozvkeV199kym35MlVMNNb+rvPwzkTOD3jBVu+hebyEh
CBA8Z6G3qmv8nKFU2Wz135DM9oJPbfM3+ByN62vZtZKZZ6v87gnlHVpF6lAL5odd
zYnvI6NShfe77zBUX77Z0MltMVoAUlALpsJW03deO5xjGFimkjc28/Ao9579O6yK
uKqRrAon0tSDZc8xMjXDuk8VnsQxP91PPuO/AiD0eeQ4acns7YfY7NgIfFrp5Tc4
hODfGSEJAMG9Cdm8uLko4MhiINI0u3RNwTJ/0Noz10edn6xbGykXe0ucAe5grCJo
OphU0CsTzXeHvdpeKCP5CtCJmY7dadX/ycx8Da8V1QWs7LEuTsQMfwGRxwJN3drC
kETHI6VRtIx8a1jtJE6w/AWjIu7k3MRAABAGRkK+x8OaYF7m5D+Ny4X1LeQeNxOf
RmahiHFPaiI2e7GeZ2HTYKzHhPCOZPEWTzIi0c6SdlBg/vnGPuORyzBsCpqqz66D
x7lI393yniC1pwQ9ZQb4cl3ejC4ajJcZRP0O46cy1GWgd5EojgBhgYOKMnKIZ9Kc
OdYuClhOhrWeoDFG6x397xaZJ9767VLyy5ZiJarvDf+27453pe3stFBkabyGhA9y
OeSbZb5hjR5BTfliEUVOpZ+Ae8pgRDVFy3GP/rBQLqbAEAbDkCaIOqQa4ENypnsU
0KySr3DvEMwBCnbqvYgFw1V1nnNrbaUnivu3uBD6D9gshsWsnP2sLvWBZte0OJ+B
artK2ZS7G8GXH7NnQXD3vtWVNHYlqQXaXDOtnY6xjBLEs02U7sXCX1PmxkVu7rTL
TN0WIQfI07HwXGkqrFJ/oNjOSrMIcZQNqxFCeWJ2W5oj3mxB/0g1kX/pyyIsHNu0
IWFFv7rb/LrBHCG305/yPKTo9hbrPeLHJ/hDMCDyNthFjYN0qmQOYpoT+J7CgVnq
Qdx4qk8fxJbVnYpnsEgjdbABZSLPtOzqgVlr0R2fJYwXY6AYwd7yWMPp0m3P2SLE
ywxIKV/Ub79pUDWojEgVzLmf5dFU8/ClI0BvsMIE7H/Qt4X2+Yxxqd5tffjlviH+
UbTyQaYbWrrPkNJIRiqVlILJe0EwLNwCPmZCvseQhG+VzZXtpYN0vSTSV9SzGkRx
ObRvuR7jwjipVxrZbZCluilQRn2lw+qbwZQ/1XPgVep3hS0tjDGSVM4D8fMlM6E7
DmEqRebsjl46IIvC3IicoBCUp+MFQ+VaEFGUCTAU/XuCc13B+aO1a6mz7BampU24
HkJH87KhJ043UFtaMXQSy7hy2SnAEysBy49zjJcTFhOSCKI2tfjJceO4+XXLkTMp
E3N2mOGHpBpQ+xxjG0luxYDiK4TVWbRit4fWX3Ujm62xSgMbIcRs0AnjujPvtPKg
kBEFxFHAGDqxzTSTLSnd0Us6Jl+5CnD/F5xxL07bLi+u1YQVQ9TV7IgA1Cqg8SVC
+QF90LiA1k23IohUOYqIzcs3f6YCRdAUwkfRGmZqPqOHpveEePxGn3KlVEPVIkzq
u7gaVCeWe3j1gct1qbMGLJtCnQH8LCrYmEXeSowvonO7G+TLs+FYplwlz+CIIajF
cvZtT86sxX5gXIKeiCQFto92yTe+Kh6LsDm0SpRfj3NTYKdPx04VF3FUC3NqgejG
ozlFZW2yKTt03LEWJ/NBPEmy46GmN7NEx4vQVu2tbisDbWhVix8V3Q9IleNmeDHQ
eNTQ2aE8A+y7ZZrUwtO2KesBPD6i/ea15RRtA100B5PyrWkbyexAH3s7zCtSWrb6
KlkSa20TuCG67nbo8byNfwA7Rl8PWcrXabxA9Bz4Jw7FTc9gvH5lftggiVdaZSum
zu7S3R/dythecAGjNEUVNTUGKzcULnCotfi49mrtQVsP97IpThbX82espsCvK8/f
gOhZLlHCWh2V00v+WOq8nRHOdJvLEJ5Vu9nFmbtXy7NxipC7Kx7b/XDDUAJcBqlG
IVfFQBHhQ+U4KimeJoMRn+dPlsyfdavALrw4B6SVDyKxquP3dMXAFDwsKbALpSlh
gI+nhlYifIkvjOBtNmng61GEJQWBYzAWjOXlCFzB3PLRx5UiuMZ7tLjitT776MyF
zLUUdBKI2jzcV6U4nKTY0vq7VK1Pbq2CsQjC5EGVJgVRxmkRD90913V65a9ssMc2
UPpyUcezxlGYZ8N/UdT3S86+8oZmewe4wgb3fLsDh0isAvN7UO8O9Humqxze5iKg
A6vIfo/YsVFz/LNXgigyFj+d2xEJJ8S/U/H+6DbnK6SmqwgVVUBa51Zluo5+1t8G
K5VFwcgCPcFf8pWixmkl0fcPaLikobSl31WPVwb/F2gZOGkVRX1pxj0kY3ryYUJT
lmPpbVen4ZmRl+V7dUuMhSf4xFyToFijez1zN2Bfy1h8WaNnqylh5M4BDsOGdV3E
Oof1MEcmXhb6ZoMzhoip8VuCaHRbRG8cjZpI0u6LCQ6Q9lxKImp98VKq1WEdgp05
7YJd5PJaugbj5CK8eEKJnWqRBywglUIAaHiQNhpCfOmYx2uBzwTBesNpgxRaJfZk
x8bcVYDk11ezA5bsTDdlEJvmml5gOjf4SOtaNOseYs7N3o22oQFsuwgp9RQerkS0
L40xMSHMpGCpBGCt+yIp9SsJgbPLw70mX00Q8kk6AJKm+47ne8Cyvvl/Ugmy8IEv
XBZl6s1KLo03hA3Iw5z5n7nLNb+hx9OF0bUgEz2KY5vhMlYavLE7Jm9ajDHLywiI
RK91PvzoH3OUSeqeko6IGheAOIipqMZonClYX0STaEsDnzAfKY+sDGnrLT9y/xPL
2Z+N5eYCkdxFwcZdnS8kOeKbvZel9NuMVPeHhThEPDSHcVynxJxyb5VupF4Ah6Ch
kHiBO7JgQSjU5hSEmpzJyT1mewE33q9iZO1zMuiFnMPGtu+AaPNb195OVWkvcSXO
nTrMwe6YFUrH1eGQO4GTItltY/foob8aY4PATakIitINBN/zLdVzOwozntVg+dKS
gwzAkTpm+IC9VcHK/b0wHqRG/0T/hsF6MkhNAsrzl5Z9R5h27GDUSREcgJJOBI9c
+TcODd9B1yoJlp7RFY3YhnUWr6c+W2RGu48MbGRhE8ygoFuvANO1T8B7vHczbwd4
2mycycqgirHuswnBY7v+u85GMK7qEK7Z7nFZ/TNQWdpYc48/lAGDdj4P4g6M8/nR
MSfDxbMpvwiIA2q/z6tNOgJVubMS0lSrWH9lRxWEP6Xt+WK5KnNe7GNsTzH112+4
sVXtMAhb+HS9T3brX0Dt5jDeWvRk9XZMQo3Mq1MIkl0zB77VdkG1mLuj3GEAxcRR
vmM4zS7i6qeRUqXcoLBlUzuQ0WgHAyKouCc7Y1a7FeWF+PL/sv6FTumxKJCk1RJv
FxBJe2G2whv92QfA+oQ0CP9K6X28jOMy/0i+fSQ/CoPEKyVsDURlCfQwaY+P0LeR
0mO4zyh0CN6/MtCf3Xoe3Z6X74gHMRCF4nXhGlH6IYUJ4hsj1UtCg1OW3nK9Y8cv
E1NJXnDI7t8zq4EZHbeVvIeY6DOsN02JA8E8na9wxWzNuLlkpzYXos2fL7odmTxP
rZXZ5U6ZYORkiRITUSdWlEoXXcYTGeBiTaJxDIPj2pks96yYUzyzpE5cj0Oha4Yy
RL1TU7W/J1VYCENwe4NLH0bdo/Dkby+0vX0mrZl6amQsHEEHQFBOA/+PdGNWSHUH
DBkx3t5iQjI4Vbg4RKSHF7cp7gLaOl94PLSN/UiFca67ihaCJRglhd76z2KnaS28
OK1OA77dK+rbcxNDAxhcgMiVpdIjmgZhe1M9LtU+nXQXDLR01UNXLcirWYxfDBov
SQYAf6VpGK1DPI0gY6bcqmPXKgih3d1sKgexKmXabbU8Q7XB1naYmPvUCqnSLTbh
PZ6RMDyXoXixfO9ItgnoiPXT3HZYwAEd5c7wFmIOhvaAFIsVZKwzliCCWd2yI5HZ
j82SkLCJJxDJ+2P9LHRP6mBnKcn1D7O1zR80gNlMhBU61RbBZ01E6OwP2DSHI7G5
bHhvFR8lnBxDXOgCsOyPYkzpzYLHMYyIFDc2zKIkPmfLvolooOU0d9y+55TN5Vns
x8WV0FnmjkFeIwfT5YPKcQ7CR7NHZuvI2VH9py9C8GAd8wP3S4EEcpbIjXo7Z2BU
rIpia3SyYjEOEexmj3jJPa8IEw8cV7G48cN6/PhwugJowZu2/q2xeERx7OAUQr3W
ZeG7BgwnMKdxK5O7eQcWMydS/vClGqhH+8hACO9UlRpA/73lLE2BBFAMKEV+IqrY
hX9VRcdAMl8mlaE31dT67iTMvGth9a6wLhF9L4C3b4iPJkk2kUc1729VaF+U5/V8
hPbYSYFPeT+PXiJNmW858ccpNiEwDzHYvKd4m4EDi55AfEQhepAY9yzEoKg27gm8
F5C8eHiUSRdiKOgg90lyrPf5w5PHJpOjLed+mhusoYu1Bb6xgBhNIQ9ZjU7L1VBI
Y412ioGeJz39lRYpBQy89Mc8Dso6C4/XjwRqzmBsLgYn+IAR3iu8CVWX9qDY0wAU
KUyysntQkp6+fvIX7OR8LPRhSYUGioj51H6dpDwX4zmgqcO1EmKG0Ar1uJYrrZ4f
g7C0/hKVwzl58YrLczrQfxTk6puaMzIN6xG5UjsSgoVa7oTi0NkrmLe9FJWU2Wph
nAL5LzmPEiXq/yw6N5XMYAXVLaXRLstQKMf7JOlYARGGtX8GHRXgOtHshE7ysyjV
FCmVU30/ze/gKD63gYQppGNlA6+PZG9QU7LZyawBfh9iLWpZyDutrnwTqz0ss1Rg
RFglSQy16OQh7iqm2zHTFOYqIBAlChDRl565GhWc7/uVTmWTXZ8dNkcdp8vMVzQd
+ctwqsonNE2vORKz/Fj5X24kIPM9G3xic3kQXwqi+n3j06eHxvV5fH+vf/Stg5/W
pamE95E6NdUq9/pNg7CqqRE5kGcmiErEmzjZUDFP8QeEoQl/QZunuJvzt+qeXmyd
6RUbzHk1HMwfKhyX9g0BWWXF03c+AUplIFkP4fYTYSmIt8oMeYMe4zT/8rINOviS
EiPB0qLa8u9fWSIa4BTtWgRGZ2s2c9fCaajvwcOTgQW1XFr6o7H+ExdlcHRECt89
0tixZNBYLcTch9aa6Gv2s1gICXLc0jbHV7CceGlf8UTIZAR78LsQ4usvWCq4ZbSj
4tyejfYto+4ttsc9axDYR/qedRAgR7O754xasIo5pvyZxJzNfEkuHcLvFg63F/Zh
EISZQqIB+cybVpTCZi8MbZoCdeGlXYZvSuN7tn8l2I+vhMmEnBPs6BGhiq/Wsm1p
yN0RXyULVU8XUPvjN09WwjGDVX7gREdXYiinVNNj/MLUcMSfnGIGWcsYTkJ66+DQ
LmQO8dq6bpQym7SacFvpq44APGym2CuYWCZCQXfHmtT1sK8x1K/+uUB3pe7BJ8O6
+Vl39XuCJm+XcR0YdtQIK/1ClUFkwtBU1KM6C1b9V+Y9pYWMbITEmFUGW1vjPrEM
S4MxWfuEbRoOYEdhmSjwvervPn1WBDUBfl/1HvMSnRNliCcCJ7MMgbtHzLZAHxm/
U28a8to5sCxhBp6SMnnbPXjwFMmwis+XmytKFfn0UagtawwAydNw7WegoKdpJefZ
1Agh5fARADNOSqN+5VDqzhHhFY8idNUQcWlnK94jC71u7TAcL//dKTzD0zUxG5l4
q0g67si8k3ontmF4jf3jxmFc1baPVAB2H4EsxE+MfQykQU31kE9+AhLA0/QSBWW2
sIes4ae9glUQAXaS2z2JlNyUVq68292dsbixW5Sebi+tnci+1lCjzP3rcyXZLsqe
DmFNHm+gh3IPt1xOUEM+CSoCK+VnX9J1sJIhU2srDc/+VTu0l3nZ0OdYA2ZwjdiP
HN4N9lQV18KgIRGyhnXmZNDA7kh2MOUdH+u63519OWnxSVl4X8nYXHpBs/E9rojo
To1MNJI0BM5T7bK6ptC1Y2py16BA4eVvDsa1CmVDA6PhNuEzHd0Knbu92r7zQe+G
lekkDTvV80rvCmPZrgpL47Nd0xWb1A8zVNwwohh99rLn+X0DEq6+M5DHuBHCTn9q
nuPdUx587UevT1BnbVPtZ8AXdNwjreQWpMnynrfXIXVFGwCuYi+/vwbenkEcJCOg
YbOEs48CQNF3IcQggwoZ21m5wqGCBCUikOw9oJpsqmp1LN+GgBN/lFVogDvhC2Yv
fWtuJTZFasn4EoNipEogX64q7QwFgZyc5Tgwdf8GIU5+VaWIIAM3aRQSpfqc/1rn
uA6pCEbIDOgZw59PsekjBxvToBeAmu3PzZDGZk/Yp/cO/1vemp1w45rWcaOJuGCI
E/JgP+xethyG/FtEVdrg+7iKEs1OSqb+jlqhfJrsN6qbGi8dUtmh5lhrfE5MmOx3
LUyNpIp+MjB37cS5tkFa4lso0c73sL5ttMzLDa29XBsbr+/FPzsAXledLz913BFz
e9Fr+xhG1jw7uw9lEv7ZEvP7pWOjReNtyvDe5HYh1AHEWIBffQD2+W8e49+Ul1mr
CLoCU6m73EnJvzBqcnUilu3KKG2U1pVE+EnX8pEdYgO/TFH7BAobUUx2wxn9vPlt
VSeo1mibz0iBDBzFecRYj1aMcTBKkuKESn9DumKkhE32imDg5q+YN6ArsehBQpDW
+BZSqktzqDVllvfChuSaWrCDUF8PX5oI/Fk3hHxZpLnqAgrojwLddsHTjYxABiqR
JguddHuXRXQN9i7te7YR4LL0UPQv/y0q/1ebchqcARKDGQSK/HPlhhm2m4FWXdjv
yOjIhyGFKMAXDiIKkScevQqmLb4wHnpAUO11MxqnXwhorcYrSk1oYauCLiUqgdmN
XD04BaZyvB4t+QtWplyAQycnPoxVA0e5VaDohVCtarkaqPgfikEmSWJrre6dD8FH
Nop2gnwVFZshPeMMbwKXy+YEOPSASNlqhKtc7IrUJbH5l51/9WfycnmFlX58RkT9
N0To3XTi+MI4dl2gE8l7jKORYBCctrFX/xWrz6zuJ0rg6mj1TqbUtWCx4Elu+M5U
Zyxcqc1bj5Sl+sXiq8itD0GrQ6HlDbJ2sip2NbdKMSQRB37HCM8sZRNgAv+t5TH8
zY7KiAQfzWbwrSs3MwunDf1l2IHoPWJVVLkjt4cM//J/Ps1n2eI5Hu32pbQlrkSv
hIMROVZeYJ9HPGg7b8k51ee431GTvmRTdLd0IQpJ4zlP1UJ0USzFAeqajC8M3K3m
LsdnY07O6gBQX7rltpN6OBqWA9PIcLAkJQOzbw2RVVv5zw4HHUnImPcmmwi/2M/T
H6ysTirMXtq6Q6F/hTf5PIpIuBzmg55Hgp8l1P4Zg9m3SuA9MwM+0f05VbLR6YYr
7Ge4/hLIrw7C2IIcxh0yOH56gqVVzihYd/2xD9iqISz6qDnav4sgZaxFyfx8FM8U
RvVW701xdqLX7gB71HaijuqS2/aYbk47zBQMTNUkW9J6CID3kaiKSOemtyPPnas0
rwAUcw523Y66WD8hORlWRG4bUlhYQNKmocP19FzfsINHC4g1TC4hpwzVg82FIRse
xnxSQ9vn+5Z1Rc5P6Nanjf2cUArZVbUU2LfmoNMIJgPnVOXZFQkP6qAAo8pH6zty
H/OpYz+FQyKL7dqHfJLkHyxDXaUZ02Gq2vTe5mSG1AxPlAD2D43vIvGZM+rLyTx0
7nfS3Hoo5exOln9Q2cM0bbj+O+IDJJ8ofFmbudieqDzYHTCHX8EUUEbvBdmLWmBW
r6Bt87Jf0Cgc168XHT8IHq7j9tZMwlcs+jQt6LL0aT4QOkSSfJxOiqyhnbGdgvkj
+KOC3cOhBBGSHheuCXIC7h2y9oXV3od9rHbeaojfcJONuUCJR3s46deEDK0ePobF
CzPLis3oC7Z4Egl10bXUVQJDyFcsVfdNZ9f/J2g4IJ/AqcmApzoFFT8TbczXg8TG
R8IXaZ3hQRo9YlpvtLsADPJItStlUbkAR9h8XZRKcCY+Wq8JNaBrVwJQppqQDtGB
TyWG0SEqdZHP41W50ZiHQ5KQT85nIl92QlLlSmskK5QdN/bDJKvV6AmzFpVveMSF
O1WWgv/EU/aFPFlfERdkF4AdV+Fpd+PLPkUsM/mMSkwWcgwn1I/1qK4AvvyS9nzF
MbI81qmLGqsBnf3uzR1wGSFFVtxHkWarMHYfEwVgbrU73cgjzYGtRZuEZBFsQyQ2
VE1+QZSRDYoYfvxN1ahB4Mch9aM5oOLRetUp97ASeAPwr2Efzk4bQ5XbZhXaQALx
KUEeLPtZ+OWbaPwVENjjnpak+qavO2i10aBHDJZAdke+WS7K+aM2/ijcTzYlyKDA
sRYy0VgJg4yYJmi/T6o1zhSYydSNS2qFe4+vydB/lNdCtU/vVFuS9VzK3ZviEjWT
MQAF3Ol2OgllAtdMYRoGiGgeFe3dEo1zRHqILIlu8OosuMDZKAL9odUe69BJQEoK
h+NmiWXXUo5gFApLnKtJ4NB+LKqF4hEjypQ8VNmKGeakzqiq7QdviWVo8EdIhCdr
UPEYFd0s+tsT+8rKLmaUf2OL1ePSRS7F+xOwHKqa35xhxcOnzR3gr+Qa+UJmYEwf
anhvlhxV2ImLSkUv2o7o1tuB1WlYow35wQwmj4pi/doEGxgKJO8oYqQyJxf+cDvH
nwSx3eEArkl/OcdUgtPtTqydkJ1xhM2aboTav/AZkMQ4J9WKuNzwyy5tIjL7nR5f
IiQD0my2h7FeNZB/WMcRiFgnpiRMJzYbJvuId1lw7E+di2Id1aOvS/5Dt6K2fBID
QlJkSyUESEuTKgGe3tkN1Gl7niQKbAP2iB7ejAo/vrSEjE7hIhVkMA3TgTh9E7Kh
X8MB3Iq6z70wacMDl9b+OWKimJYRdpsGSU+dQ1vd0qLbEUzTyU9YlhQP52YXMVtr
KAvKc7B6k3Qa0sYledXiRnpk8ZomnIvDi8zs3/E80i/ZJO9diQaHVUbP1BqjljMZ
RlmHYYBUPlC000jeJob0c4hi//F57/xmipkCZSqIPrAAdtZFLAW5QrFqaNaD1aYQ
oQ/r8VYXEkM7UVoSAIy0yhkt/kOddByXhYncvzc6Dx7dValpTxFVenFf7HaVBL1Q
wnaZ7sNyhHPPIGZMwhzmHjk+w6ERb+nlaCmsu8dlsoeAeMaE94iQimvFN6k5kKpo
0G0CHom9s71Fgpy8LNRJ0AmcNh2E3dT6+w0QYkj9ay0jDLltBUiQNSrCLmLu5Kgd
RcFHUZcV5ufH656BOf7fyO4Igt/Pm7NMIHYsjDdvvAXMfctAtAS/SgjipxmdI+SP
CkzKvXEE3MnwSnMYurX8segh2RkEfVc/45ZulFH2yBKqEogWlAH38J0eXCT5wo54
0eo+ht1FpLihkGp7P7xVdIWzcZpBB4im4o6G6RCGF10ewrGK/mrrrnJWSejIYeSW
tMHLsk2w5gJd9Yxs/9eSF1nV0LML6Z3zDVWMjnPSUkItf8d9E9NUWo2gCk/CF0j8
NMwt556ThAxBb8ENwKReXZnWgslG+cWcCqipk4ZfJNMQPiG4xHYUx+b1nogezNK6
D1O48zJALPochXPYK6sb9xgX4haVDxlFCVVf14xMAwIz3nt80mCFr0NVOJmnMiB2
KZt9cFwLm8iWyCLSh2yxnHkA3GjXONLdRvsn/RV3N+KJvYi05SLnMt3VAoSZTIKZ
esTnSe6+8RJIkNE7P9cqwNbZJpa8NEyj0HRIPNO1T/CCO0jBPcizr0dTF7EfqSQj
SxjMn3wP0wFT5rHu0QTGOvuAfHxKwRgHcKbloX7qQsxm7lDrOD2dOdMS4eM+AXUX
absPWMoZU0D1GmK3UY5o/i0hBdQ5zpjRlZfQNsXOqNfFVs/O3nyQYrikLYXf3PaA
m0iflPTlah6lrAW8eLUgRPaSV/M8FzNv5MfASJ/SCJ4CqmqcZcJwonqNw8kVSsX5
/MvNKn7mQOzRyXZSofhxUGBLhTNENOWCbLStiNyKJ6wQgUAcMcmIC47oYkrtO6V7
zBfAx2oEZNR1hkJgUoOjdzlEsT+Cizc3UH5N6Mbm99GFt7SzFQfsYtzEQmC5paMw
5YBwnWI7lr6eKbEBREciBF/pZtPxt2E6qeR59ZQHaX1AOZZLR0AUi/7vZmmSvYev
DQS25jCGf4HPnVOBhTDcBdExwJ5/9BFycnrKFjZfHqTENV9oow4r8///HoKHHKnl
H0VPDIM6NJc6M+/XA7HH7O/H9G6DN+3HwgktSS/0Ga56YGnkhERSaKXmKEDbkXdr
bbHDPObtr4ZMhtS3Zl5Do4XnAVus/LWtp3N7Ekf9qbjVm1Rx2yLR5/3mHy22rG2K
MxEgl9WKNJI4EYaIlsYzDmqIwkH9X+dMJ5HAEAfhEUaWH3WavKqC4GEJQOmvch3Z
04EozNDWLA1QgePL63hTaYSCZPw8tdKLevhX18HujBtCVW3A/6n3ddyJFf8Kb84T
m7ehhYL5Rs1ig0WsM05xV5dFMEZWqKw4dgtBp340DJfh2yPFoIheFnKfl1pBEfAc
EKhotQrtCda12bmV34jX5DATYckBxiNi42OX28QN+BhiXZS3nordhH+5IVNTf9M8
H6Pzqf3RRSv1J5zar2MdaD03B3ruQ1gTNGFwYbQsiHd/Bx7J41z7hlVEjJkUoJNp
j0ugJIoQpba21XgTdVy4zCkHaQQD6sZanA4/T2TpasGaeteKrqXIrnkFzRDyRxMN
DHtzKiFYJSX/Qxc4HqwEdQ8UWzf8GK0ayxe25EmRRrhVRGvC4rf0tXicIdandkXg
+sXxpt9lJJ6ed8f3732yW1i5HPoJ5rZQY/5L1AVQXT0ipYAQGum4pX5VD9tLiDgQ
AcbyIDDBOgxRPRG2TbwWZZhxHAVTXESeKpGzug9JqwwrqbcU8qMtri1aiSYnV8fI
YyldsQI1GWwLzAYPHPtu8ds/E05B/2Smat+sdZN6ror+aIFUF7tjJZmvhsXKJFgn
tAPVNNWCRcdLPDWvNpSmQSMKNcOpj7FUedTmqynGIihpKQOcguhzsdambWwxo/XN
VkjaOPrrfzWQ3iC/VZqwr8ubx2jZZWYaM6FQLq2JBLJn77BrGc4GZrE27G7nkI5S
CZ+yWPLH2c8UWzpop3MrYgjwo+S+s39ObtLA38mgMWRZuiMLjHR9D9ZqkA28Zri2
O5QGqjhWIUR+ZNoBRe543Dn+mO0R6iUQlD8dPkQWYTpALzmrUUvbuFNStmOUOQ/O
F1bN7M/qqCSY4YM5Watobc+JJogngf+Tfu9pBlPJ3s96f8F1rxdIhN0NeLvvjy0Q
+UDWL2k663tsE2ltaqsilKzGB/xVssiM7lAEgm7RHTLts1FyR9O7K5hT6oql5ej+
KjRyT91Y13oFknFNtZ3QvAn6TUF55bVcM9pWH6X+0vlkg2pnbZ48ouHImZ0yfajM
uuTjgCag/YWPWiOOr0FeNH+nFoD9NhPi/LFdP98YhHmB8foxjyJOkTcNjkO2Mn9Y
tECm43NjvZH2U1uojFnv6lG/yUfHgdWaQ38QAlbfnOxw8G/bd/iWd7pCH1NZphFe
V50YetSDZqLiEXqfZE4QiAzWVnzoMp6UCG4lSAG46vtTuLW+xZ22B/n89U6kDcvg
Kh/lNBmVc5jpZBahgfcuaa4vbfESEI/sMLM7crW+7cJzfpUgJiIiRG6q6qvDSsZP
O/5RND3fe9KZAefHCtvXWJyKBbud6Q/BBua4BVg8Zw48FYUbCAKK9v3Q60QQZO5P
eiZWBQvRN2gpm9Yi8KlcBzlV0mwpsJwkyyvM443ne8xJAWTGMaIcbQbWe7kTwgOp
ksiE9hFcxbB5cAdOM2enlGYEby9hr+96M0qkKVdCluR+RekyJikO3QnNIeF1y7fg
o7Z5H2aEwN4WoSSkz99HYBMm7wI9BG5oEwDShrnFzHFnxjN7UNEc+tu0b9sqXJhs
E27fgeBUv6wvg18dStN/0L1SRC8CPWeGy76r49P/UvEB4JMX5A9S7ZgPc5D5WCGI
4PMkcB1Fm4VUUgMHLHpR7TqQlztVxCkfKExPAxlf9yqdeIWO5vV7mMOawjjSlgLz
VX2JxF0LISNmuh2whYJBKBWEeTbaO9AQny13c5Vg0A3S2+YNltswVDFaBiioU0eg
GJVrZlomYAxTQS/Kv3vzUOFrdtHVUZLggTsA6yeEPIqb8YAlbns0AtrJDPKNnjRA
CYa3r5LfiqraCUWhKcFBqhQhERbIWs0shvwBqksjLCbU6V5+oJJVSw2qVZcLoq0w
r3eMR5yzymn8N3BNgfiveejOXJg6FhfLmHaahwlaKqnVbi4JfvyNSm0h05shkYBS
0aihzlzDpfeZNvfJqxlS8FmkIcxIeSnKtn0cipng10E6xOwYcBqg8yzOkEN/bOCz
cxqUxwtWXDlcNSpsTbqn1Ivpof9LQPHx/1MI39Ttk2ea/6jWVWei1eRO5lmqvtOf
FKnzdKF55ez9NKeOXY6PpaM1Cw92Ur5nBlsXEjOBVjTW2w+zk/KIMt2q4ZAaXUT5
/oN/8Pb4eQ4c0jQIUZugW+SvPaFX6LuTDUrCObNE57fE71tjiQ3qldTajPRllPgK
jdPWiQUdFNTuly0y0QVXaQhQPSDNY0NWIVCzQ79VRoA9UumIlyLjWZuoz3QJcNzJ
ka81vC17P1J95yiwfWyLEgSVukvQtYIbeWSzSaU5i7sRqZnYhxNeLle02NFAJ2k5
WXYnU1mKvRcB1vhR/Xzq6pQn+qg1rp7U5NMHBSJ9GfA1eaXpePdZirPYvUA01Sgm
o3au5ekKPnDx8PgBfCo5VUB6gtSdjnAEgOCxiBi7W4Pm/p6G595BSkKf+a1B9482
FyJFX0rTMOHOzBYt701ByNBP9TSdWFFaUI55IXYYqu+1CCqUtpG8MKJQpS/z27/K
VLWRcuMCscdFVw93ssHhvqR0gH2CEzJrOJyWSXX7pnt0pxmZwIxdjMXsFSsLnb2C
kd1fbbKzMgmk10q2H3fu8NbiSie6zqL152+BINqzh/Pq8aCCXgm+wxZUUvmHclaE
e32kdcM/WXoaEDqX0qw03miOnQ52fQO9sBGRRC3NOuxnAtDAeTp9ySN2Z9Tysydh
rT9WsrX2VIfUArMtj8wudtSLYZNknKTywKNUmhOlwvYu7TmK/9eo13d9EOy8J9ES
sJ7sTrdbG/yn40NiTOgVLx+j0FrDWCUMjHTTWcFZlrwCDOa9A1IG92wxgdLR3RFt
j+akCcS5D+d31HaB5tVN35yfg97jKpjnSF53YU05oaS1qqO+lrAIhN3GNCKfx4+M
QMWndt5Np/7exBg+DZ0Q5uGGbbqN0Doi+q6bBEe3PZv2s6HoB3O28uMZgaw80gkk
AtFuy+gTuNcsQeKY0oM9Tn3MhH91bkHBBiuXY+qspe4DwW/C108KatAGdH/h91WI
JFeCIfcJDnzS2ZpXwlAeRtc4xZ+ti+3xLet6kDxjfTq340o+dBx6V5I7a1/IQPho
MJUc/Dy99wLl/0snnefZ4PqlyUWA5CeIxvCsuFQtfnw92ATsnB3rPUdZfkOEeXbR
2E0zfHD8HKJ2JeDEpmqt9QwnuYyVXZdZqjzwSOK8z3z+XCDSYvGTjmGaYxL39MWS
Q64xBhPpRnYeOxMAT01xGoHFR1Jvt7jiJTDGFyNK4rAzn6TYA+3w2tb4+Z8KlBGQ
073hmWU8J2A+fTk8Nj5u1QE5brzM9Q23IiXxsNuULRdw7SPBKiJwXZXz9nYc32hk
q01EQq+zuL/2nrbsF5k22AohTCx2WnHlCEPa1/TuVD8Ua+SC/ir4vD2ijUIhhsji
Y6iGmnsS/uMSeHwjUaoJmRiaw7e4so4Wad4uzBWwmhgaCTofT1eqXgOIv7YGSMA8
08O23LzifINgxajzA3xLb5oFTv5BL5ly17kePSjZusfG7ZDa/DCyMsE6jrhSKwGe
5c9vDz+oQe7P1W9n9q/jygPVwVGeTgmCf0+GmvBFMV1nIlDCAgZFd4xzjv66Dp8v
4JEUK9LHxdlfvuBqlqbbEFkmO3pJTgAMu2bjDvttOAzvQYfw/sYpDwLPDraAemYX
SHsR//niuDVKNS+idas3aHsQ3hYf2zDIQQ5SXsq7q91JSdPuudItiWRYkv9D77W8
ggS+I9yHJCZtB6W+b703GssbiGR5maUpi2/9Jv/1KCD73shRBTOd0iFP2e3Bduaq
B627OJ5k4xfl/Xkj1MzMqInrhJQ0DmfpaLpmLMwIPXoCMOMPsLgPWl748dG4IxLj
tiXZ69tfDbf4LGegcBsNIiVkDYD5U0GAlCJaa+hWe3nZEr4nd+5IkOVM0hbcrL/+
AaRfC1oUlPSHdSpbTriAJGUHOYs9df2zA2FY80HR93Oy6AWsMK/PgR6lcgfu14Mj
j4WedhqqHyEKaDnJbH3kYTJgSZzMqJasLJHCV7TsFBwDhAmlLxArAk1UbP0AQcA8
TlJGSGXQ6fGsOG1+CpUMIhczz9tCtrM8k6KI5WqS6bE9vwd0Zbb0iZbeMUQTXibw
InB2pNV/yeZgHGEJT7H81nTvwAHaXldOLBoM6gaF2VixBtmT7rKKC3DVKk65ZwIi
aTBoRpzz3ECTLa1u/Gg0HOfXBXOw3PActNbuP5KdZFd8LNKn9RQlwlIui7gubLmx
mWOGzP/efcF2a3g8bNQjNu5Y7TfPLCK7ysoU2T3lzgGdKWHLxdt+RYGP8Ixh+QJ2
b4LJbuZmB6m2TQRd3Vcx65w/4zvVvM2xL0aDEmPkKJUMF7L3hckS2bD7NLJiFE8D
pDezPcibsVM23y3GWif4FaNJ5DHB4oFwRGKYDVhK66ur0VKl0AiywuWbl5oDnpxt
1kOHYtc/PW6NJjKH8Jv4ulTSvS3J/GHqOFwXBxzw/KuubX+3UPYMVMGoUUYpXSEj
utjWnxuc/TruhKPyDiXlPC6BIP4Bd8ttE53Ey0g5ihBM3xICax6fyVwwr+lLL7uN
zwr/nROZoZM11m4DPLBcbA6Dvtjv3OhAREcfRArLN/9u5SpxvQZe3fpwIn6iR686
3wdq0pRrNYjSbgSmo65PXhKL2jEEfbR8dW1xduwLkgVxuZ0hTNnsRrn493aHgVdv
r8GbR18sCCg0wdWemMUOHe7KSSekeNxVlovcw7bAFDYM4fcjb9OF2Y0yNySQ0rQt
eOwRxmLbZGtl5/6TOGE4+bw7y1lpI4S21bNnMFCyeZnu7EkSCBH/vrePl4u9ieb4
iuiGLdxefNXAXqG6PsGO9nNVO54NIbE4YfzurSXTpyRsCBgeMRB9pMWvsx7NnC1k
LcI8uMr1qOVANP8kRc+Gf/4SJ1Uy7ltkq8kJ+Cy2Xqr9vFbK+vWjICA+XeQ9jJbw
hKUrPNXbmeCaf5LAt5/++o1/9I9AKskem+EQ780kPvlc2MiCP2R5eM3aIOTUWctZ
6ui5fBFkBDKWZhUXD/0NEGb1WIiIiunauORGhmfjPRQSkScisnIRfydQtlzjGjhY
toeiOSx3QzBcATr5ylD3Zp99xt87YNE+yyx8Z5RjUy1+AyeWpyS4iNQU2U4TE9e5
APTYCMhSl0FVnIQqNuZB0wskOzBvGlBBDcP00KGJjJ1MLuGWN/vP+66xep+gC6b2
+TpRKx1IZAhn+hKHdqrXLLB9hL5spNsEYZnPoO/jdVVOWD1XoVNscOmOcTaKy+Is
nzou391UTuX6lt/VdF6F7i1wBHbUc8dkeDgOcZi0O5hDkxdKmuLcvOmWOB+tDL78
jNy6hFANXwL+BDgxO4LCUsnFPKc5l1DnnbLMB974rZVYl2+t2vMFxrOesPfuiEl8
OnBYtolHRwg1DmYFFR0NGev5j3KbeQb4B7a6fCc71OnmfI3RMqFS2fRMjmelC8F7
KIXNmrS55JFzjAE7rT9wAnBvlqcDNN2pHNJVEojhF4BkBGnGYWgfY2jiV/AdUoDA
iR+OcBvJjIEpYHoedPrcMMBEo8cbQiZG4QJEUVdKcbEjkpT6hU6wq+BUDzw3RXHS
IGyfExuPSqWVHQey04abnH99pgfMrMwQNgbiFeWOQf8HnEprLS1GJLyu9CrsN+s8
FcJe1Jzf8ntkSqvGzE1H5E8k7tREknhNJWvczKsXkm9PK0uWyw5tEQlk+lh2PQNo
bo2WGjZhq1Amiz0vDaSy9cNKzpkcdwlBFNt1/jMODXCIM8wTJdESRULmDQxIlFxH
Qcka5/NnUvSIaRjbiYbdcZEx0q5W36Q923sbI8tIKrA2E7Tc7+42uTGnDrVVL+OT
Mc1Bjv4IPe0bdQ+etZtskTOc6rpfgVklzjIX7MzqK+PWQaAkOmyLEofjlwc9/c9a
t1yoVsF2csz9AXaQpAGZtM4uQD8+1kgsOvamwE0QO2qKVvSJNb58ieIXjCBvjhh0
G9YZB6XiCY9Ic7Qu1/BBG/QbiJJ8rKdeNNIIykXQa60+3HI3Jhi8IMg/emFjKoYV
OPKVhWW/rzbbENOAdXShhgXx1wB+6yHheag0LMBsqB7GBFoLD2fNQe3peIPEVYPL
f2sfcPGDjun30S3+5SgB+meFSU9QbElJ+AJRn8AahCuL+BHzylhHOQsoduus7COd
vQ+sIR3ghBZCI/qJPsK8DX5Im0VFt1hW9Gm5bFgAaGr4z4XD0OxkhI69IICoEPdc
doZ/PMibX983bG86Ysa8zqiRVBPip5ySZNhKFRHANXypxjG5EB3WaTf+Yaus8GNF
IEsabw0GdlTnABRizWNwZqA7s2GVO4S+U47eV//Stgf4b52QaWWCBEkMKrh7BSDV
hCalNL/gDk7VaXZME53U6ewBhLKiDJ6daFBZqRFHecUGWqC0lXei5Q4V+5uy63ol
vqH0fZmI3Mv05py1BOxvqg3RbIEToJ3mzIXCI2zq2SSLebmSAsutKWxOzIFHHB7L
ppwLTkIHk+9oRWnLyB+WE2Ilox52iSwS1TsV02pMMFvjiY7e1bGoA5WeKtVf+tsu
ejzcbG4eu0Pv+3X0Vs8lmt3bzdS0U9QEnezkYGvjnSn+IO8+bIePOAxW+Da0oJtb
pbiFFeRd0RpvUZO7zNBzap/VH1Rk5pZwur/yma5ZIJH8WbxiYodfnz2ecthLoZ0S
fxWodDEQgSSmio/0ydJKU2qq5TgX79FbD3yNFnyf25cjTxH9r/5RLUpYbFwDaT4n
e35V4XG6CyWDxslkaQ5XqEG3MtOBxuUiu3pS1ElxFpkc14B5lZhWCcVgG21jkLK6
yAFzbny77mynOaZOdmyEM2r1FXblXh58ybV+XRMERN7QNFxvLdkQ9jLfpBam7Ds5
zZo4sucSg7/vurvkBvhT/8Yjk1c+TQT2Uxd8Czrty1jhrjYZx35iieHV9k3r7tJX
JoNkVcS839RG7BwNsGpGu4KcvPKu5klS2TrhzPsOZr1PlaxYJeoNbcdqO4f3+313
Dpw62+gz6tb9Pty+mwK596eEhmTvseY4/qMoaOoVJ9lNGXezjxr4mKAZGKdCwU5p
QNVuWdGvNY2xgUf1hN9Sbkzc1AMcj6Mx/DkJJzENneAxbC88U1+dsSS0BhjV1zzW
wmPpCQMc81kspCle3+yb5P0QiPFihyzKVDa80DtR3B3Geuh3MxLq2fe0GEmMb+tn
fnU0rWo3U0B88aiaxeIppqrlqAxiKP5A4+Nt9BU06SvfDZk54xuWjUprg6m8kRma
v6635tfA2uTRrsETDTin2DGhDLLHY2rfdPsOq1358jeb5LqrVi2zQ9K3zUQmB/v4
ZYavmNicJX6d1JaRW7QkrBLysBL21IEkQ8vNVei4KdBWG4mMWt7kXo+3tTB65quG
uO1PlbxNmnHaUkJjOg4PCDswMUoZKjiTkThIlUcDSc3oblJrEjFuC03sA4IlQznQ
94qkNTstqpVzw6n+PdCDYXMYunAIqxTwGcPSD2yC/6ds86d9A4h/3BdzRNSOLj7N
xJ7ztF34UDOFtHFJldyojdcrra34+lFyEAhsf4Nf0cB3lClcNz7BSWxKWIcpJkn1
eHixulLsUkt4JnQGW40xGGjWS2i+hGtR/BA5nVSLzdG0i7mgcgtHP63aPZ31erm8
/26DLmBxURAV8sl1jYuJAP3SPxgkUP3+5vtxpM613HolxKgYM9OleAiff+yehFna
oBY9I3Pnw8Q1AwhmfvwTfBKnl+yiNnpOU5fTWgAjoaiLdV/E2fCPXWQupAPlQTVx
zBfqkX1gKwWft6KPUQUX7kCw4rqQXceGIf4RoW6FlG4Ht5EvAwiC73X6sX8dBGfW
ChM3dz14cwAjewOyif3ByJw7InZig+GC9yf6BmMGcdk/bEMbINMjwKGRGnMVAwzV
BDHr5gqe6uMmJ3oH+1HAq5u96oEDmFt15wZBEaZj365yacwZUWHsXeyDNMgmm5MT
TFLjI27aTSsZGZxCN44JFiJjOtYCLCdjDYIoJmOFuscNSbpLuoAc75Ym1JmuK2qf
eIHpLPtkmiabG5JqaruCdZx09HNi4IZukLXCqIag4RjXbNo0o4CStNDbebSTt112
wQE5vVNGiEySvqhSx5KXN/tRz6Ykc953ECBvLHPGXPd4AIX4znepZWBCO2cfXRZS
7VQWgml56EP7kCruZoIW81j5KgV/scXf2bQSAE6i0IDzSOQhvSoqVOTDh19fy6rL
S7r0LScXFQitUYu/Ow1pTgCe1pAsjjfiHur9oUn7MprPntDf5xqq2BcIMUpNERMQ
mxjHky+zZ2mGXng9UNQnQHQmnlR3BpO26hF4xtF751/1ZehhWkuwtWb3NbpsS/VL
AdMhbdWyfHF5G74lr6jxuPXbeylF7Ce+y/tjtQJNtxFfrGqyfvu9pzG/77EIB+nr
gZlN9fYcKmdzig4EjcQys1TZeMVTiWB5DQXGJvzPKLIplj7900pbixbUU/PCzcHN
UAHa6myf0Z0cfZ1IljWm7g8wTRz6lfeMbCNBDFcObw3QsAkh2BcqBUok84AAosrE
4E+2owzLjZu0Hu+gioG/Ku3eMuNYJzX1+XQ7tgG8wQgYkicUhemB3brwLyt5hxHO
QIVaBIAVC9zHNiCdS73KR1fmvOoKgrV5yk6g0DOdwsoa5HANHd4XOwl5A1h96C/X
WgItrhc7kIK6oD65wcz/XiWgBWoXSqp9pX8eTwz8aNVmjK00rRkNtS4fBAt5hgR/
LAY7GQTOktDuBqFHP3Y03IXfHOySV32clH5mDo5nf04wucVSqmrcNStTBcit4Aj9
ZPnrwMnGedrJO7ElG/iwzjfTu6Qv6VQV+/QX8xaqA+T5zYvoZ7YoUpPRWsVXUv5W
LTcSQZ1NOu1cq5MedqY6kP1Pv4eRsEA3R+6qMeRWv/zpab1oSiFgxXh+NVU76iyi
djuuBBr+ffAplMFsNesEqIEK7KoG4qH1LUZtJ/c8QEFdKacUOnQRmr+hiaHhXBw4
pxseOIUioYBSUG8Mc2Yxz08Nlf2hh8ZnT+55/cM7Prfq/e71F3O3wG9Pbliawt06
VrokDVw3QZH8BOolI9F8eL2LPQR9Laa3Pyi6vKJZdQxXkd0LFFA3ZR0HTy43RhpF
6N4nYXlbN2bxaEJSkNdPnIO1gyfpvIWmpwXg4adYfcfBr4dEcfQdoUJsfuPgu0Vi
2+0yFvi6dvRYrK2L3U1EfCEjG+N2xWrd+SqJz4YwCfVe0DXXbXLvfiKk6Ps4+++s
uWGUY+ms5+BLkn6sOBj+zZupw4w2ASXItjqJuxUjtTZuuoJZvugngKqHig5DR1bU
5jCBugP/GfeYJGzcYLpBzEfj2xS1/E6snHWRErQ22kfLQj0b/Xwdk9AKfgsAA9wu
PDCeLTj4LqmjDCkz8aFPlQQ5yUO0/VIE3dqk/sDFeRvWqIvp9bXG7inQwDcyBuSN
Q5axs+lYFoCcDJ95BKapmSHR9+wYfdI1/TS9n/6J5mwvvO6hLBBUnhuboiuBbJyp
PYY7KUUsj98AHpMSfumZB6s6VAgNLNfXIzF1D0hjphxYuN+HiWWq4aKTkXI/EPty
zaUClqX25C4Gd44pivHgqN7qg83D0PbuX9I6M+FWmViGCVz8wxaG67QGlS9F1umh
zLqbG0rMMGqzumKkge0HTeFa0f1YFMo8uwYp5rniuzHTct4JZvykxmOy7Y7Sj5bE
E8WIn3GBquw94TJnaOze2twmYtaGIapHR/GVGq+/F/xnfBQq05X5b9oVayhxyEsn
TA8pCfCrFl+AsRHHgx7/Yfe4tXM5AE4LNhDWZ7fiu3NrVtHWSWrq9rqlSvVfCdk2
Z1K3jVk7kvMz/8/DGv9oxjCiQdL47kzLHJRScNKG3vngoxcRlJu7vBFlEUJgoWQj
lUT07IIN14oH9ZfgF9JDl1URj5jBhTIzSuUvSQ+Yw/wINthx+B7qByPY0yF+ap8F
tyF1TDKXsxN4umCE4R2B9oLVV/2T1G3niMA/yxWQwFcHNd0TcC3WBsSGiu2JGi64
JN9Rz15oQmjY+vrx0L6wyM9nFGTRi22BnW06LjXMc7ZyzEpTNDItWQfO7w3ysjC7
1zacC0XULBrx8vKNsT7/y/r1e/fKZ/pYoR9sRpPLhnmNAA7V6Kf+qSf1DDV9b/OI
4KbJ2mwAiI1skdoNALeFWOywUDCw6pQ97xNFwRqZHrZXfrAyNBIbOahWPmYND6Y2
LyYTA1keP1p420K6pe0jBtvQzwoRgRN3XyyB45ineJFd7UQFZCzIzNXXioLuPRa8
z1W51Rq8Jrk9MHR4t4zZO4yMUQ3gBoWDjK5BqKMAlIh8dVFAa3iVN0HaEzzYtCD5
jyKe0paXRm22v1HIuqkTXqZQCZdJS6YeAURKzzVFVhjBMbi+m7tzhGhkKPxBSe8h
N7Wy+5kCqOB2BuoNWs0LgltYGoSFZjBeZRFvxX6pzJ03VSoicH/VJLxNoprUzZSC
UWbNcWAROIaVLMQ9zV404s77882CcyF50ErhEXOHyWekcgvZVzW4PzHtM1srjcC5
wOP9vXiolppNZDRAxN+Atuk309yzhGFBQGXaX0Q9i+SLM02yaz0vgL+dKUFBXRSP
8KD3QgYdWZqjsR6jG7p35tttyC0VQnbNgxuJD5TfHqFmO0G90MIqR3wEg8OlNAGw
eR6GHuiAUp0KVEhYiJAUko5HQgeSvNCBTC1z9gTbi7O0SDc85rbldjqmOmnQtMKp
0IK2gdysxwZzuLWHL0CH+CsxKL6xEXF6VVBnkFUBPBPLw7yavx9Dyy+LL8sB3v7I
mGdLIc0d72mjQ8Ix624kWbD3ZyyUKbNwz9w+aveWj/Wp48qtvFzYFi+TlXqunzKJ
GUvTZNXeLo9tOFlzTR+y3Fv5EWXqzpM4zqTQUTGWIgFHXEp+DfxNlaRKzC8Cqfb+
6T0tw5gzJnECdBlC9gLNs7lYo+ZJeqJK71W5TXDm+8o5pmhnVVdeowRYpIje3M9j
C6IhLpoKdP1WjXQzfCamS4nfeL0h32mrbwVA0bwsGA1K4hCntn8loSgZtLow5pNP
QlzZNDFwhNjFfH7P28SZ3MKvmkqGTs//1ulxzzRg+4lqTSZIunYHMhz8xSa3NI03
R2h8WU2YutcZB5SM7tRpmOxbmAvS0jycZudgkyqRddL3tpAfDgOe1MEI4TpVglwY
Vm22SrMXAKwrsoI3cEmDbAPrbAX6GG1xVfW1jYG/808+zBYfnUnVV1t8bjpNpSCK
ok3AmQQSXXMnPLEgrSg9tybBzTduaygI0LnQIISz+lYSFQoO0LTBAB8V9JaVAjym
6OU7tBeKsNTs+Az2IHYYDA91qBunSqWmQHMp9uKS/gyG0197EZWzcYPwijQxMap9
BYZ4hbeVviMF+vFIKG+kLG9pLmFt7YgHkS72hViV+OnmwUHLGw0hMPUhItPD5n5h
E4cfFTGaHhTjuv/cX16Soj7hyXA8c1nkhYUnl7wmewIaqMsUn6+vgJrRCaz8kutE
bmTkJvDfyXYZSNshFZ2+dK6zlKyjyLFlyixefvYajeORDGaz5uKR14O38L0LCkAc
CVwni0ogDzHAsk1T5wZXmb87uMFzFfhqjY71eF8x7y4+wFmDf4OUTIIy3tX2TZxz
fat+a9Ns86aAGLQPt71mKTBVvwJ/iLt3OfdcNoU67KmDMYM72tKIfsPM4gKZ2wnG
8Or3v0XD8k9CQeUGe37LLNqe4QtRURoRS5KQ1AEXopJ5CbAhOWxxHuOF1Xfh3MJR
dzgmfo9AFGK9cdo7jhah40Rt8sLJnNMlD+hzIzA6xqNIKXMNE+XVea4D0stBrFbA
1Jx+LgP++VBFYL4q3Issp9fKQ+iwiiHKHNF18cktQcI3OBb0DbttiNHNl6gJPDii
3F02RnnYNWvOa0K9kvx8KJoKD0S7R7pL59guT2ff5+lj3+A43/RSHRvOGze46VVZ
3kQlfO8rXVgJMM9RU8S01fuSFsf8o7i1B+f6qWoAk+E4EuXS4Q2MkHGGokrfBdRo
R1+NjNdRvI/IwhJ45axOcKXRVEkb9hkUX6+7EAF+UnLx+iOGhe+ETws9+0kQYeo5
giVkVtmooYAp4BpM7L0X0xbRrBKJQMAV98wk6OfMgdq+JrhOHIe09Ps2MkaOy52q
AZ3r7ER57LBvI2PARMpStN9Uogm3hA/hbJiZ3GejWyWAKv2yxoqNsU7hPBa5EwVW
aCIKiD2t1USvkx1n0KqpWPGhLJyfpkscFc3C7S9Mei3odwuuBCw8q0kAdMBlRyGq
ETNuBzE0sveFtFt05NfKkb1MOFas1rop25d+bRRDyMo7NHVz7lqPxVXo4MhmqSPz
V6ePICiiP6hzM8ANAihiyHyL/qZwWJaiiDc7Kjl2KJ3OC5FigycN2sq0vZ5zvFAC
QkwUaxzDZ3/XQPXnw8dmNou7aGAxpiOamFV1fzEZiv4VK5VgR+7PKt03aWzIu3WU
Ey+Ix/lpAnIx10sjbuHNAeMJ8PP8KWFoW5/A1VUK8myirRkahpCDaEJbA3nRMRvz
sCx+Ks0lH2x5GSWpYUwexBCdwKAWW7XY5S3qV8GVThlPjgy7SIAZ1dsb5tuAEdW9
iuxEHCvenqN8UaMvGlIHHy4bgNDDQ1h0i9NWslh70xwEMIAPP0Kb7VtgHQ1C6ePY
6s3hBP2wVDG6uTAT4zQOt5nV/sYgmGlSHkjuHt5uGM3NP/LpbfaEg26z1TRwRMyX
zpWnmCdNsTwM2x9tLeH9D6qdf9ClB5qiHVNK63FTogo0v101IlBUsZ8JgrdmpwWO
H67Txsj22opaN+u21CMHjcSQTy0jx2pm1aewf8wMS8VYUBUwoLKSzGp6WE+0iyLZ
dQUupKLzZzjru9J68dcBICzAtoieHs8cmUsyJVd9h4gObC9H85G5t0QxsRGJ4vvo
DUE7VdSIVW4DyWW3RT+Vr+04z1McnAvWTc+9Q/b8IsNJw2eeFEAzN4SevTgexYjz
GixHMXbvlFip87+vHChoG2BJ789k+XLWVia9CP0zx3Re8uE2NNsKBBY0JTvnDDa9
aNTNCqfnZBQWfJqHIYi+yg77URO0SjF47I95z32W8nGV+F5aTaIx3YYU/MSjT/eC
EsC5fKIGgTr9ObUv68hmikIJkzsNSG01ZZW5DmIG8hsFUHhsuhnXCcb+y14mofaP
bkb2sw9eNQOHjrLlBNEWlAiKO+LcOfo3TA6J7qNkrxEL78Gyy+WaUIFzNYBv+Tdf
UHNW1iSzTZ1k0mHDinffy1rUMzxnCgPRY8d/S2UkT5JVXz4pTfHJvcFVc24zhBtr
yxFjSGAb7SQ7tKhTdfLDo6SGKQks5Ox9rJJGO8FJjWQ0i9A2aNBRlrTKKYye8P0D
Br8L0nW0BCEVKdoCIrly0jzVP+N5zL0MJPLSaB5RI8QghTHQRSFrexWuUX2AHSpw
1dixR2ECKxssj0c4WeuDyWA6NaOb0G48McE420a1kaOQmzkVPgx3XXWY3ste34uY
ibhu2aytlwBTDpjUuXgmMUQD0rUsU70pZ2Dsnybr+rjfiXSHFKliuZj5zw+Iv5t8
D0DblILQXgmgx5cI5AS8Wzgm+sbKcrLN3yk60DI4Yo5ZAVE6TlHomyiRLcQwXVGy
6XYMz+h9pxNhZ0jacCFHFbWj1JHIfypoovZipLXVyU+OoqbYxfFtRXVx8ZwUhUFr
OieCAGgkRJpf6j5bTm5hPLzEGsTyLXRGMTRME6mCp2aoA6ATa8c2jCNegz8lcvXz
q+vwShCg4tjMUE3qLXerYvQTH7Kxe6EbDb6y8XkcjT/AuAR+NU2rH5CLH5NLtfDQ
hL6jCZ/DZp6LRmXVJMo2m1/Q4nZY+53IR8HumpPhWXitY8IdJXMk6gXGuCumcKfF
s1DJ1Vnj7h9zdxVvuGkD1uag0/mhAsurZhAkyKFFgwQC4C9QqSkXI7lTyclYLTl/
NTp+2WStFjAVevC13aEt60NnYoiNjeV9Ti2QXLnekrccm+qParqbUHwxxbfU7gIb
OOrRUw+d8sWw0IEkTyHADkNZrUWe92Ca3KnXCopKqahsbPn8LTmw/6wneEOY0UPl
bRgfwvGI7Gf8qXqqDU90fwDR1pcSAdJFA+LNnSoGk+e+1kAzE0gyM76PQW/v6E/W
f2jUKD+wJqRuRmALb7MVrJ7piZgDPhgUot8n/1Mg51uPaxPW/gNPedgVistp8XP6
z2OnB4GlyE93+cNG3XCeHO+MCK178IMLac+zYFRKgLHdDuvZcGJeKxi8NbDM/Fe2
nOwI6Kp28TjG2RD/ie1S/05soFxU+nskwcPhn58FyaY4kMC+YT3c5wVBp+QM1FN9
4GEj1+pehEjInNSecqFO//QU1P/mOXe6JL/lWGxHxNf9do7HyoRGWHJCLGSXRdHw
0h991QWY6MTnHVmnHesKlTKssY90glVKaH4Qz8ihObontxQSVgUPuhgu8BVW1wAU
vny4MLGXk2JCKj7/4vj8igCQHrNasYG9WSAUCYHfX8zlOPc54XYpC6kGqsvDni9s
J9QVDnf0WQX4wOYTqtuZ3C/WsDqPKD3vE+/oUKcpwrwccZc/tWihS+m2sppYi1GA
5ZzmMQRXqD5mTmIMROCzkxWjzH7RZiyuGnk/6EQqqX2hLYqVtsSnj05ULDEmRQeg
RR4g0zWch0TFY2ZaS3ehjy9fTwfIiOq3caOMZZ+WkR1xvI1qfXL2BBpnbrpxbW9o
Kz7g0gdumLI0tYijmw/8+EdMRdc7Sm9a1mPp8HTPJc4Qeg1SITnV2mAVEpJNehn3
mo1aIxaYnv81d0OqZcJpEyS/6PjfygtdIW0qtxeVswzEFCVfNIPQG4LO+dmOLyng
Nce2tYy8xX6iGVP8wQFZrAM6RipiUf3Bwsi1QJxk68p6u9ZpoSHhDxzHdIrbrliC
1vm9donFfJwSJguPtPmmEE7juxKsj4Pdauk4OnB+shddrnOGivNzChWLENzHeIab
QxE0OVnOOpVXC1bOuxuqSeoII13XWEMG7EkJpKr/BsTM+SMcoxtvYRXz/Er6y4lc
XIaW1hHqKgXHJkRuJiPhPUYk3yF51kajVcF2GoMgx1oVlZ8Jg3NzMS3TZEClQqAX
Ey+dg5RErxVXuJvUBq3JLgYzcfuy2kikmSxwbkxahFqHLku6rqOCcdjnsyBuriMg
SAO/gi44uk/i5KqWzPU+p4NBUI9UK8EL9JpOmOLbXabs7a887HqW0mp2ME/M+T6u
JhQq570TnFD9pgtQzSVlAXXysso/o0EihEcEQS5Ih0fFQ3gRmdvgooz9xYuXLmpC
GxAbZYntP/+3/nvFjM6ycBrxLLDmYYGV29L5gAQpKBZj02lalkUGWBcNgHWTIL/B
YHmouYFBRhrR37I/PLhVBkVS9U5Y8G66CQxKuKOqDl2/83Hn0AmV2iHR3QqPhevG
mV4XO9h+aMPYUtfWAKsZ4wuHXub/qLb9vN8kqzyKc9644r7FUyoAojNYBHyk8w9g
rvclvPcOcZt3ljz2pOMA0nd9q7ATz21ye1h32H8zMUV5ffsFJVeMljhL5ISS8X+F
tv8pA7Lra7HzkyBEIdJMG/gfHqdAZLdF8WSYYDP80fmKgpvoNJ8U1bDBKcqlhCSf
aKketIrWtB+KXxfR3LFnj72PyNnMoE/0cN9temnsPzryhp8rLGWRBBbzsdgBdPEU
3CSEX8DciqR6FQK9ob8xs0dHT+z5bUgEcd3uQBoAUisZ49tJ++sLc8tv2Zh6/Uty
K1zexdlwNYVDK6X9ShRnHzfEi/6EUJgAWrNfjOHAA/mOWfkVKi1IA+PBuZCd1/sE
Vhv4lvbcWiG54ybpRgmgiEBmP2w00Bnda8tH2HXqSMkmEjrWiTErhiaUheAHFqZq
KPZ+f4+gGZCoobgiKyhEqu0iVE+dXNORhWMRVYuMsQHRgCddACmnN7UuIYqfJVis
TkkjmCOzsUICaCpkSD898bpIbQDO3Dc9AQtN3650fATbsT/STy1TscWqS8uy0J2l
qzycjYTojM9CNQOBXOw65MfhV9GMvDmuA/eOpBx0n0+2IsHh+FRf8JgSjccTTplX
FVNhnB23k7FzALEWPqF95UFJ+gx4kTDBqtRYnakMSpo+IrKD7422nHVyWXkD2Qv2
e/MPZQhU7b8UKJtSuOqZFi0wx4kkxZR8Wm4ZjIyoDDc4fJsSY+Luf08nQBSivNT/
FMbA6cIpD4KqtYSmXm1phQFE2yyiGa89EovdoMJ9Pje6dk7chpTH3wpEa5mUyJS9
U5UXy/bJNCXq3aVmeW8aKzCIWR5pBt++9Nrtcu5aH0ZdyhZaq63kwW+sHybpDJWg
jbMk3AP6MgefoP8pT88F6nRrGZETOcHeO0BtlCf9MTifL1TY/BziGOGLgo2xYeS9
fmY9/MDycLHAWQklTySz9aMhSNX7ZCUtrAYiDdWIHrzQvY+PvBl2p3cnwMDNFFQK
2BkG8qE/2sBy4qejZS4CDpyfYgmApWjOcWXamHuZ3Z3+7wsNVUDiEUpAd8WJ+ZvV
qLWxB/JW2fQaFz76S7urXNWchcxDzCMZzv6c3L8gMboGTlKvjrqf08VF9AwfZoEf
Pg7QD5As/APXZo/hwwBFUcNNcs3f4boPKeW61AGu0enqF7CSmK4P3qoror0lUeEc
BuOTtOLAYxWjjONPyKorNX81eGUvgsDIKCpDQuupSxKl3Bx0sBYBkkopG1mALQX/
tBPtSUkHyyhxyZd+v5kpGq0Ue/gXTLNpz7qiuv8rvyO1gfxida8tpVXxbf/mKfnF
L53RMcmK6/cJ9ryRJcmQ0nVngpfoj4U1xLkcaEFrnl5d9DNiu2dHtpwvLGL8QPIF
BoGoBqhMgDfe/328W4ahk/ebU9BRLjhPRfc6bEq2U0XxJGHXLp1sxujBFK1XvgIP
dp9u5uPKiFbRtyBKQ2p9Q2VMJlA7rS8kAVsn6l4oYsLje+0aA8HlYHe60k3p2gxW
SfG3qh9B1Kd4zXIjPJt1oKeX0AeXRAroJfPgFSGGaYczpcRusTsYSsfSSZPN/KQO
ARWmtRu4CHd1i5Ok3zsIkZMt0smjeQmIpfHW7cNORi2y6dgqs/5A3dOVEo9rXJ18
MkgUn2jtnvFkefKPUPJ9hrOPUVbsKSyDvBODmXHCJyM6/JiE5NOMeUID9Yg5PgIs
WZNvF0DX69LyFecDtFAtwEpSXFG3MGR5+33AZHyhT9elCnGsgvy2DIlp6172Uika
ErbLTM3g12ZRmL8Nm2IJ+4OnBaDUQbE5+XHOfKGBaX9q+7vQ65mQdfUMzTJKKcKB
gt5s/jalrdDEPTzhSvScnhdHixK+6y2qDhsvH9og15G/kW5EBkMubmLnpZp1vHnX
JHFnwPpKJJZ1KEBClnVfXRPIxCUe/RgxvzjZiXC6550x79vo2MI7BFlPeUjN+1rd
gfCHQurg1hNs9o+kG2PUywb+Z41Ck6Dva+NOGmEx5bmhhaxyTCyMHzlvn3cDCt1F
F35ldo/N0qh9ue5hTsgG7uWtR9mYpZoKYqaHot+XpDBY5EsLEcdX0R7hEwqa+ahH
Tb0SNb4w6/Y4ceCNeL5EUMN9ReFTQGKB5fZ2MBln7y/Kk+J0TEfRs1Q0Vd/RYb3G
ZKDinxLPlN8d+RpNpXNqdD9lXhi+o8S/93DYmkEFW7CYtlaz1I5OYKvGHLe/gH7x
F1FLhlHk9ZS+EYmCcaw6QL0NP6q9fanSYVrVzpEvXNpMNCBsTzXyT6MtaViuYoL0
3tw8guYjGPobxRsihuiqpogdyRy8m9oNQmZquyFRs0Pt2QamEsVJiYv76ZhKNL/K
ir8in2lp4SJq3cm0Z7msfnzT7N5tNcdKUCfvTV6uMVnJF7j85+zbSVGLdo/1889X
LJnz4Hel4p6IimGqQCLNrlEasqMxP8GdFf3VeCrjq54vmXej+9lL+/KRRv3BRBT2
klL+u1IemoIozbwyQ6lE/Kat7CjN2MQT6MdvtmVOsvl+Jn+Tz1AlyiZaxYT3fyTy
9d7PDW1U9Qk6QMm9BHF4KmCizNCXMsZ9isV4n66yNdpXcZYJhFB8KZr+A/eXFUeX
Pvwu3dka8c7GKHwU5MqHQyszHZwlTVH4BthRcDKmLhtSLgMJH6IC9HhxrjGw62dC
mozwQ/8354P2Cq1bHfkqB0QQowX4RzUUTCnRO3yWHb10vJ1Nl0XS3Ae/4Mj7OKnv
1D1AH8w6RdKQuYeiWIx4LyS0fUeS1JS39NZUufvOhPsC4VYmb/anYUWyIH5UYbB+
mhc4OsGNAJjNhEvWquoKwojCZ5Gc8z8ItLNZnJ0o+/1KBF3b5/qtB4dJIJm8+SFR
xTW3cU0Kq8cWZ2wAzkJ4Sl8AwI4c2h+bV2a9UXe4so1IboA8amiVg7v7iYH3m5s5
o3qCgcJV6UUDKzOeY/3hH3FELigGS2jG/HnCZBkXffc0udOrz0wqAiaSqStFu+XE
UpXpxmkWBhE3ka/kPvOYov1Z/9ISYW+qPUC+b9IaLtPqdy4cPUF8uD6BnfT6IgJq
JRWxhpUWoOWxNMkouLLzYty66bW2zsFV7656p3hLplgky4KDfz2dhX87NYqvmFjC
ZqDIwQ4kuoFQDd4E0S3fFmyWhn0ns6RtpZV2iLv1c/yzLgBf9fCZt4wWUlDa0VC4
aQz5lul2kwcXn+DKoqh9JmhvfTrto8Gdd3/v/GTQkfKlZ4D2z78L5NMTD0M9e15z
NLAUhvCMNG46RIYjv/BHl2HE5mytnu940IMueiqn88pTaRQ8jbyXtusgQ1Q7EVvE
DnpMcorGV2BaYUBB+iRBg+j7JoUKAFpyBgpbpJ2rXmyBJx+HmvZUNbd2atzyCD/R
EJppFKr5/5WhsCfj2GqVU9UUXhsoYyOlDwZ9THqFyDZRqSjecmLpj9gRQU12AcqV
3TIZ2vGl17Fp4hcD674yepgBKRwQtnRwdSQ7SAMrsjLjSYHNNmJ8fxZq5BxxNaWD
GNEtNpJjuyKtPHLBzGX16coOtc50HA5W+5AkdZy3bTrzb21G4EREj5Tt9V9fN5nX
PsQsPL0GzPh9qNA7+zTLSQJaKoe4aJ8pYLL46PGZ3fz8FUhlgpAoW74Ka8PltVkD
X44n9KA6xbI12xwSeoQgZZ8CWIOYzwr2zAwPxaSg4zDYKhWzqFicmXdwhpucnytN
SMTOm8FMvbFXpNYE4I7EJB21v0+5Jd0YYm/36lRGjOU4fqSUyqLuH8LkoCkxJ5qI
hdrz6skJdOPQfN2QoDzyhtWx21QkUS7T8pMYA0UEg4jjGGWNuHER5mtfz2VAwfJp
NYOnUwsL+PR1VLzi8nPFjIZAII//+GZUR0GcCrow7M2laVTJteHtFzYtWZkVekn7
9N/lGzthct1J1faaQl4IoPppj/Dxh0o2KW/hvfSyp7W3H9pZbCffq1Z1Dk44PcbF
s0rd9Zyh6aPCta/zQOsFZQ9ZJZFY7pMT4N9e7k6oB4VJNT6OOaubtLFY0tdCq7b0
HvA4/8vZfzuSWBJG6f8MVmbfxjHta7ITVRXYnURVqoSNL47gi5CqJVZmOa7B0G8F
Sr1ym0LLN+Y/Rn9U7LBW5HARUeZtULPyUX+IIH/1r2BlKdM3CSQTIDqzHK0lxjAG
MtgMBLjKWOLiHLVMLxq274WcrdtuJfgH6a5X3kPuq72IBB/9MUISWGKiSeGKc5o5
RRgn4tVdOK7nNPHSB5IcHpyEc6w5P7+dczTGGCz2IL2MTMddxXFXBBE5i3pSz2Ih
0hq7eiP/Rz+HQVo5w7kah/J2OnNk+CESQWD5gNCMCq/rfyRNzbkjrYMeEx0If7LS
bNeHIEaXoDhT0sCbWyi/KJGDxm1PCHfbl4RL9y1xAoDwU9IsDdy9OaqGVI8DJDqw
ygxS9lVOZ0qwUUAbDsh4v3llps9Xi86MpXOKxnScN71E0HPzyiuVQUO/Z5yWAXAQ
zc3iTXxQHVSzsv5y5jG614f1ynyd2FsqZZjUhrihnKMI/16cNc7b0swvDxkcnjYG
LA+IAo0zun7s5do6/W5wXXrIuNFnXoKevHnjLB1lwgqZRY+NeYfuhocfBK1XWr1k
hH4MIX+BXa6aoiMZpo7ISCjqRSJl6x1E35r3FcJjQU9SSuo5VtyKKo9BVXNfc7P/
U4Oy29fEAR+wNCFbRExzPXAazOT0WgA5AttpEquQjvbuzusLVtYlz8E9ClipGm4q
bVwLUjrxbCIRApB3u9ApwKmuG+NV2At4+vMhJnHUT4vxCcSWyvkPK20gqSKJ4HoV
jIU24Fy//01phH8+iED5x6UaMpHH/12/E30DySMwwgPV/I4EkE/W4/KRLMEWXsFc
Cz8oeZos5hnyoKgLu1ELzg1ryPfexg8c5OVR6ilzIGdibHsoOAvlJV0Q9H0A8tPb
SPnrgRmo5nkx4hRkSBEfjrRvE6QzJ78wHzY2M0NQwx5WgWnHtQ+vyLxmUUDlP+qo
Ak5zN6/gIgT/KkvYdeRtzW4mbxFLXpeJ1wEBcxU1jXjKxflZCR94Jwepyhrfy56V
t20VqMx+JJuL7caKHLSBKVUtNxdmFpgyDYK2NGnCiBxUyWZaS+q31h5//n5G79TS
OgWfkerCHEJpREOfNb+//s8kfsommyRy9J1siar0fo8SRvrB9eijhZ597nwQ7e1n
LmUzMgUidODMyMbpcYWUYpxUThHAk6+4bKSirzWCv1S3aqUYGwVnMjo5xk9qON0T
eymKse+A6Bf07QM+0qN5vHP2Be9QpRoeVRTmAc6NoNqrlnZZ3/ZDK4HAUpMUe6aW
I2cuL22qTA7CboHYO9ZuUnvF5NpNcABpWjiOEMHHfsXVZ2v4KC7rW0k0iJDy+2oh
GzJ5QW4sYMAieFkPoeVZ01thPA7XIx9XkF6fNh9TcVB/pNrXD0XMpmQJ1IgcAgSv
blwjXiMScLlEY9FijBnu2LI9GxNjrMMUjaWIP+WWy8TJL6UqLLmhQNGqyCZJ9Ly5
IjEXhIgH5/42EzrKXqXwAPrO2VVLb2NmMdC7xPAF2Naf53CC7KNM1rYT+evSy+G0
kcEetZ4tfVoy7urkpvvxjUxMGoIsff9m/i0FWh9+gVAuHZ9E0WXTGDvK3cbg7YXz
62YWDmnmTDaakVDdkEhJacjqvnGG+McdcqVP2BHFVk1h5ZfVe+Glq0aYBd3OlmZR
ennhpkFsj3MsYUriCRVLsJxKkAur6vnG00YC1qhRBr+1s8mmi68jGUJxm4Dwkhz/
FpYCW7Q+yxOsGFlRPeQhAZDM8/fO0kL/qY6lamuUnU7sR30pB/Krk4fkMhsXydRl
no4Ae3jnoR9jRwlxBoMHGCVABDlkesRki/4gPD+JfNjfRhhpJfE79zK3vHRodV5h
nQwVt3fledTsdlJsKFL06jfhv7NN3feoZpGvmlnKnDrRat012wqqHXmWhZlBlddh
bJcCpX9Z1udIQHZKawlU88TIOjIlS48zSH2fNjZeYvGoxDEQgf/8DRGB25rBTb62
jD1tLnmbr463ih3nrb6zs6maMhb4FzolzwzcNv7qscg4GSQpWAObzDirLuz61hG+
kEZqNkBslZ5jETXqAhm8pcwQufUrD7cOPGASO4rNkoRfORIIfaBBtQqqRR9pgW4b
TRuk/bSX5bub8soKLcNCJ3qQrjMXQXSPF78Ni/bVXuPq5bZ2bbZV7p8/nm2QU1T/
WF1CbA4CkwxaxhBrtNBNaQC9JuQSc2byQBuRFxiL53gR1d76DJVXh3C4xgJGBo19
56JWvT0t3eyPsNA/p8wZIKscF5vxmYHwA+7mnBv74DKNIbc/hfWe5iVxQfOJ4o5X
wn+BT8ropNhgU7wkYAPs/EWed6mZBPY0W7nOq9P4YDPbbPzpY3FbLBbumsN1T6mx
SgC3gm9FHE4n6HaS8z+6rn5/BTADiVzXms2dk2wj+gvoZ78TPhbIzuVGQf5Xardz
+walDBq7Muu+oY0/NqQ//sFir7ceN8Rp0Q8BbTtueonBgnojgVhrB7+n2gg0tj7i
cl4bwKPCF41nWd/JV9M0cwKuu8BAOROW4psCIWh2rErXuvjWevRqfH7R313vRXxg
4q+yxECeRUIxWprEww8FKuVX2/ywPXzvWPqfvfVCYXM1kPbrIwS11vy+GMb5WIQu
o89kxgIvMryvnpP4QhdEj7aJ+D1i1IKA8NQcG1+CafTWovxDfFQT/VzzRiN94c+W
q7eNta2WOxqCTpjf40R+EiN4kkXXBhLNKlHdC4B/mtEvv85EuKgBUyuXMtWliCSZ
wgJsIoqA/ygOq4FFa90LTgXUVLs+mHnDCclF1S9qeq0jxv6D50HxNHQ9FcjZzfJ6
Z0ADZW8E7/M/EJ0ZEtHGifK0MhqbZIrGfiK/HohBO09qbLnHYkW/Q/NVV6/Z66cg
kPQN6uy+AR4KYE2b+3KQFNExVXbKR9dGXfeuOAiM6+61EPRYg4Npl8ZJWT24ad50
qkw7VMnUwD0owBQEszpB5yjgOK4DFQemzWvbtVXjh0gcc5OfrXYB7+H++kJHTOg9
g63r8Zqi/IK2ljoTf00/MjpjOqz2WvnM8Vica5d6znslrw3zhrQ1gJjPJX1Zcj2V
8+yOdptb+m6sY6gzw3B5REhk5GXYBk2bXF/+LX26ookeKWsVUcL6cAAsIYw8ZRlw
2m28c4RxDj9qTGtr2TSMNECl1iqVORMeAs5MJoGtzox/k3959y+ccGWa+F61ZlEm
/pP9PVg9G/iZ5oPHKIGlec0urRfn7Ou3FWoSlQ+6yKN1FeqQlSPdPPcm9EeC9bwd
zwU2n28QgD5v7Zhu/3blEmZXIczc6oS1AcGyU+dvlO6fsptinknK+CNne7zuEfL3
3LchsjB0lN/OOsJ9foFogwgwtvrbdLR5CGdhYxNEsetukxjtYrVWFDbgRaC4YxPq
ReAOKEWTMgxaqcDoB+DFLYZAUxScMZ3pPNKuqzSclAYjTpwYCj3qbRKXtPp7bi7P
9k6HiGruK3hBW6zZJXehfi76MKWc5tt2KLnrMRhUG1woehWqMHapXSEY4vZo8CRP
5edvK6bHYmOQnezBPWlXgVpXLaCbIixYr5aHLTGZT/aR8g4VAHDsbNF72o9Zmpc9
gEwPjAAH4uKn7ZohjBgJvYe/a7LdoaM4SQJBrQJGgYXUuhZfcnc9iqhgdlsVmNTY
pCnlJBRXg00c6roNzcOfa9a49K7C1kLS+RxB/aWX1GXsDI6mafbJVnDwzA+ryeMK
+d+1ElrkNy3Bx8gi1b9914FJkpVEyUZoi4Yu3CByia1gQWUqIJztvD6ROw/WlWT5
6wnu+aYxsSKWi22TNFZtMNd2/wyHx+KGStZJ4JSxBjlIC56HyPZ3FNY5SIIxJRER
4P+3m6fQl6LNTQHTLGdLanDNuLNYHjHzBYdxe9bDdw90kuEzRXLTVL1z/n9Tn+so
d+0QcXyFXsyMtU9Jvfhz3BUA+DVZcwsm42xKtPgzzs8osjoK3lGZVB9vZUxVuLAZ
B8Y3xp45NV+pyF+dKk+h4ffmG1KdykFKcw+hX3dvuYBhKLowIBOA6hWA4AV+ymiR
ULxaWnzgPrChGfLINEBzGTgpJZ66SWRG83YeOejD2yCFmndV4gvSFSMFslOfab/r
tyqQLQCZVA5fbMLpI11N48etYLH0oRzosTWhTDI+drgAG+dGDMnMIgVi4VwDgKsM
TWK2B3vts7GDz69qNJGkuJUqm5aaTWJVg4x+hynmreyjk4tNbC6p2Z41XcpgNo0s
JkdBa09RDsieDBP7SyiWs9xhjsgkOrYT+bwSnN5x0kdttpwmI5ft07xITJ69d1a7
vaG+eySA2hMSC0gpjEZ+O56SN5O4MeWvPlxQ45bOI+ZYrxOvMkP/ee1ULs+Yt08Q
m4vXA10ouLXC2K3whp8JK7zaLnhC09ZthUACJ3iJRmC0UR5fYHfd7MUMzpdm6qkW
GMIQQ6z5wDfhGSLacymkyHrdZcqOx4Y5NXo5urkXvkXjBGI8/wZRUPBij6+qiwhI
3y6v0oNWmqJ+kuiibQ6LyG9piUZIQeNHaaH4r22Jt0kEL/sHdflYbybvr25MHT0d
HKS3PkSrwduRPpUB1gZ6Unnb1Q6GSGnveOBS+3g1WoBQzgN20AKOHoYcwMOhavRg
CRF166DUbx4ReR+ufFNRHqYL6Vb6ZWDdireqLLPbsceSKkAo478ASC6/yC4/xt3O
hAFRGH2MZw9RACJK2tmVC9fxEoBnRuVTeddTDK0vD8JKlIhg9pFaZOqGJtJ3mcLP
DF+ZKGbHDELs/o2VeKVql80mN/x1h8IvQJ8n5OQv8hL20y9ph8YULJ8xnbnneEUy
6A+tFqSRbvcoDY8mkmTJgQFSwnZza/awfn9ivumA7FsKPv0AyJ4CoKirInx5JS4f
6nvN4Y5nOwfK0MZSTFDpLgj5/dqXfghMJjd0UmkmvWn8Z7/Uk2DxxT20ZwWudCk3
kWnqZqecYqNW9r8jhrXVGLbZpN0kFJnPtVEaPHUIO/QMMOmm6qUP7jxdOkBxvX27
+yCuLt7Fvdpfy1qu7eM8Y9hBMVK0LaPJEkIV9d3mcXbo8LUKMizsQYXxCwXG6nBr
VdjEARGuwlhWxIXvXLHKa6166IRxNpdekQUmkPNvbFBF9CeCmdPuBVIvfKbzmOFT
IL5OP8LB0aiMnqgDJe1peNWgXjf+XwF4UvFEQ7vT05xLEQ0/1yHuP3h/q7vREDUx
HA+PUiTxIEfVHk6eoC3vdEMmEoqGaF4LX3gDM7gdUwGD0/TW4D6Qfty+J/xT9kCv
IE9ME1v/fgn2QyRpGx71NoTeIgC38tLV9yE8PO7S0fz/3mzCkj9/eudYRy4ZQiZt
mm2tRbjSy5xmhDVqGYAWaOJxUO8yIEZoIAE7aJ6Rg8ZDP8GfVgXQmHGnLWLdncq8
AxT/j2ow621MbfT3FfFoxj6Q53YU3E3sOqNlV7Uhc2mbGc29GBNYMsBTsnZviTE0
HTM5PZbhOxL5ZF3xk1ZrBVmntOoxfydIlEys8IV5wAAsEUegXiWcK5Hth35sKN0L
osAO8sprvPsc1UfJ7ZuavzAmXE69oL2S4yiTilXtG7avAj0nJYFAw5wjjQQM3xP4
o6Tveil0R29NFRYkmC6IvgDv1aVzRkP5qz6tjPi4p0j4pIXth0xcd0NEaoVLGkwm
JKsS0bTD/TgtcQFsfkXZ+72i9Y9tFtwfh5q9NZ+Xg/1ZmFscSxzrI+93zezwGqT3
XLiD/JIa4JIX942LrwdIiNw0XmFyboX/qbBZ191aN+4rgFt6c8q6gLarKwVfTXOf
/I/yYM0ylo/1Ci56wPDw8JkDiJntpKzbd1Gte3Hrr9mvOa7R2be8qnICZC+zcFsF
vlxy7hupHWfqpEMGYKzjY3HOpOSkNoieztKFm71dAQ7XKB2cSQcyK40wkMcVtri0
QgabMmeF1ushTGPxjBUFwjWVKF8OREsTvkdBBXLPmImcQoNxxV6mpja/dDx/5PBI
g+l2nBpDHhFSeumRF/1vJF7/j+C3npbxqmEA+Gf0jPUg1NI5sIJweiNCx6WCUTV6
ZxrBwZeQHpAhtCLBoTUqpuYOt+efqPubsHz7KVJFpRbMtnPwA3AsmSzOEIpwqPui
7uYWdo/ao0Ch+9zIyFnmy5afnN1n1CP1Wz8eYY3MM6Nny3/OiMbJbdwdimMnEytL
OibLZFNdcP+MPTjeKv8ZWDTTSZjLr3xkAwZ+OpCsXGWyXLwlGAWGeG/MgqGO6Yjk
u8G32TnsVYmChEDzOOnvOBUatzumJoAf+V7zt0pLLmFXka/O4Hw2+TD98IpTAzQI
7DNPjXGCOvxZkqMcv3dKRiSl1A8A1zaHA4zyXdkQ4a5Xz6qISX/lHb6jl/w0Goz8
GSLsF6O4REvWqx1I78BqKpbgdCO9S6HLHfq7YmYEEeMcoFi8HY4VjuEVpD0IoRVJ
CjNNc1epBq3Y8fRjZDtEeoz/j0LySaYG8Vu1X+eYKHrYvWkFLJuBjbskVsA5MaT6
phoAIN9zLo935F+ULyyWbXG0ofhSsBn+7LD/8H0exKZ7DEE7j8qZvPWtoVstjd6f
Lc+lh6SXIvRJ9te52DHQS4b3mG1/3boVo103Uo6JB6E8aiLjaSFhD0oNT3ZHZIEM
tv/8cDxepe0ybmkpPyx8aUXTaZxyCaUXKZhOVlL2YEGFN8ng8h2gCQ8TmG7KBubW
QmA+R8RCgDPx5yGGUh8h5szMcQrrb26O8gsP/H0DGlu35xcjYO56cAl7gyGehta3
UaGOpYFCl3acW0PEnulS0a9UnCYClvlgzrLaE7SaTTdnZSihvpJ8OKhDzwcDHFnO
NMuEyYHoIkQ1+jdS9UkxZVRZz7dCjr8hSjlRokB14X+3Lq0jECnPJYQaNrtWGZSb
njbHc57E+LKvp2z8xLCMhGeA3guamQqK7utlM5Un88O/g0EYcCz2kDRmegj7+5D7
CsmE3JlYbQqYMFosqouoYgGfFfkya13XK1oq4dYy8kuDZLS7xFv3ngEI5+3pS5Ry
J8MS6TE8zbhWWaeExCUTUSCYNLguMUKIpNcNwXY7o/EjdZvuAjgPJ9IcBwi9NsiS
ww3jGjOHIgKKn5z3jtpYvm17AyIbW0TC4ePhAprYH0lHNisNYMmsHk1korIb0dC0
xXllIGqxz0E5VkhgEFKV83110Cxus+edABdk8JsYFWjqAUoPmLRDn62meRtJQuGt
0pGxZneDyOnpFCncZQxRW5i5ZM24mLaQgIYVPys+azNjUGBPaFf5et949pAjE7li
9z1Qux7EdpLlRtswjxeLhvIVM11eLghxkZpRrsX5q6Rm6dOKOq4247x4VeoabxDU
LGvTKoAp+B4z/Zm4iYQNe3Lt7PNHgnxXMxZW9SL+jYxYUtPrEIgqPg/BJiRYXWum
i6jGO/Hw2ZzALucN1zh8/cFuvol0fUxcwlv3arIqv9uJv4iUN099Pl2I9Fx+o+LV
ANdu9+DlQAxlXKCBk5kQoy7peWr6CCa/jT5JTG9KXHMn5NO4cFwqer28PbA0hMy8
tSj0zMSMfF4yVULlJY5rI3dFsLoDWPc+sHhdct2JAL6sJaBNoNj6qiWuTxCBttvB
WRCAxtVy80nv4c7eGyE9Pkzu0j0MOPDDsKE+8w4osqW7JEFLUSGrTn3CT4pUKV0j
Gps9AFOuweQ23H0n6KL9x0sis4u/vGCg/Jf0OXiuK1oFD58vfvKQ1bYOQbDchUBQ
Z14+b18ha+p27PiQ8qpTRxEBRJ6Ve3CaPhuc8ws5HNWvBUxxPz8FnvZyzttDVYW3
1dEIHizfpuJ9DbXMUXsRQ16Ha+FWeYo1kQifDyfo3+1QHksNbtzlNPZo5PLm1P/3
lEYjg1/96o+rvmXmfxiUNsF/ZXHr3leqRa+QX9dj8M4diDvU0gWDvWgWmRGeVpDf
OwDCj5EMQROZffj4ikkfCycVJ6nNjevzQWSy5NkxaFK5PYAkVKWAsBtKNCzOL8+i
oBJnOEhgmWQSIVh/QmrSLgndB32FXjsL0xr7nPT40p6YG0Q03CEbHaikUfHx9mJP
Qd2AJDLuSGWPCTK43zUJQQMwaiNMSjgonTR0fnCmT3D3nG2EF9rv8N9j0f19fros
mDt6elqqesg4l2TlTKSCGj30fditBbohhP0dCU4NohQ9wYjGusomVhTobykFm5Bm
HXTumZJbBWvAjXoe32+6fM+rhIDvIouEPupAnu9c/0YaFTGBEgHHbO4WRMO0B9qQ
ulTQsBZGtXdAMAzDD4csUPIfVOsRn6pnXYSY7nIDZ+IyvnEnje80/SgfOcj8qp45
t0L+tmdF+C8LmaEPIxw735aPRHHs1ZJGYBrsMTKWEXmDQqAVZHR1HDQf+mQooOV+
gMdLclMZnLHiIPHLKnAFiK2AimcrENqWoEX72b3gMtgJgf6PRWO9UmPxOA2UWu4/
vT9PiFQZzzObt1x/AX3/h0zebVoP6L/aAi0/3MQhsB+9dnGuURaxhAAFe/fMB6sa
H/RU/GZzqXIavqWwgsW3EWqkNDaZyRY3/14f6wmngCGTg6u97w+yScTuJyK28azS
E1YFKxR6SlF7rpO0lJKWfBSxw1PfZ5JyUDTaNi3VhXGLyXlKvr0jogRxMHZzkpee
Z8gALMP6IBCfA55gsjGB0GfqNxGQnnB1Ah6hdhCHc7PH2T+P6dduOVpF80L85QlK
nrB4RyYO44MuqrdN0qEIAze52E/GyUHUJ/o4nCAQretrvaMbR3IoyfsZoK76RZ7Y
DugBSQ2B+ivw3MGK8sTCUM83rmdossbowF/9M3hX9CyPq/YRsh+6jVHbH14thEGX
tB4cAIL2nc8xfIfXsePqUajxyVYLIl0xiQh94yDGz8eS3KEnrGruVcX4v+SAUnl7
JAo5AesNtkXb2O1TNU3QmyimP8BHYcm8OXXzLyPXotB080t7PPbeHUiGW6/M+ea6
de5MXxQb58xFB5V6MBdfo7u5iA9+c2szcXpOCH0wTJ7L6c0gPev8PgXsDhWRzC3m
u7txiN6M7QNOFVcbH2AEdVG9MI8CeJDC00Q9P5LTB72y98AoiauQ/EjOA9kfMK0Y
0L3wrKaY/v6c0GL/NEgnXOArpKefnbVEBtaL04VVbWWRXUJYC4C1484E9VSJDGSN
OSDXndXW99uAZdCnZDmFbtVyhq1Ub4JtBwmjEGCVQ1SXnx//0typUuZ9bz4pfMkN
b/+f9v+8Dd3ihHzIek25Z9yFlmJpIqmRFSOJ1zBki4v+lzC4lskS94kOuFB13WkU
iKxhsk3ENK6VfKQsXWuRTPkUe697wFbL5e1XO9Lbaz1o7+9xbZAn9jVjwaYnEpEK
WitdJ0OQ3v39D7SxhtwJyCetGBu6nWsGml5rfiAJuTQS0i/64p+IvFpbx4DVdLAL
rWvymtX0m45bDJixJmLOAKZ8GmdENi+yPb5BfFQveyaHRd52JvJ9SlLCL3ugWWEv
y+b7Ho1UI72sgQ1ad46xltapBPmIXOotQqSSVDt4GgAHvDZVDyDPbHj2M2b/FMUD
HAVdueeUhF8wQA40cqOeXiMGux6KtcQt0KZSRIAGn2pghnE8BeDSZ26MnE6UGRNH
mLBy2vfvOD4m9/eGhrgzEM3xn36ua/uDfFdV/E1uXmcWXRRYx3SLD5C0a+XUESnX
d2Ka7HeI4Bd1mT4ss1pQGNeeUH40U27b5nyuZiFFkaCTWdZssncONb3nTLUCf4zr
XyYEvhnenG6obd40EJb7Gz0OFYy18+G5rxU7YASYsKuLaeUxZ2+HgrADL8RKiprO
JmbU3TWsiGYEmIczxYMIa9gIneBeb1I1D/UcloqgFOeTKzYhb54IxkF2MDXXRNqg
LcDNkz/3Th4iowoD/5lUj3EtYO2d+ZQc3Z0+ZzT1k9GpS3CV6TN+haXxnuhE3/ht
ZmhcmTCuowwy72BQygirYhYbS46JZCKBHyPnW8m5Kzuxm5T9jx4fQybr9qG3JHzK
lnzuN9ko4tFaVULql3vbajeBFvRAVpgV0eLlkNtjezj/1TxupC54TCx54bxJAfvi
y+QGLGGtyaL9rnrDBM3z+7SSIqD1CvT9qJGqe/CMtCDhyQcNh1ZyFtdSrZUO16N5
6bJssMrlstwnL3cARUJdn1VFkef8mxlc0IPHDeqQIRQrQLZKGbyaqw/FGcgycFx6
fpG9D7ayMz1vRcPgVWGauTyfjYr3uMMEfP4mwWeiehfcWGCLuoh68GmZyJ2GymeF
W8ba5bN9Tv7fH5XejB5ZGMxsinWPmTf3Mbz23Jbs5yku8NDO3nAIOWBU4zLBRgl0
83hFC6MXTl94lvd4RvhBvtTYLlxaxdoXZ7kmShkqjT81kFdCtmDh8Afthgumalr2
m797x1a+hxC2HC6N5fVK3zEqnHnhVffcgPgaY6TVo01rFdmo6AfZ5QTRW7MdXC3L
vStuP7xoroJVn/riIQbeKi1m45ASzbfEUM2TXlR8mUQpbdCEdx1/p1/seS9wZSTi
GF/Xp5fWhkXz/hchtJ6HlYuYruT5MJq9pnY5IeZFioY1KTel2S4H7cfTcBSGAtQ6
TtxbOXkWxK+MJYU60urm9GK89phOpefYggHEUuWtClXovL7JoE9i0CE2LdtL878N
LSCGAaZACJjPYVpxS5lt0vhrPFmcBZDPQrcA4iXWfPioxVtgMESQZgUvPWqdfzGZ
q1w0tpKpVn5/u8VjE+/QketjJXCx5mvO6g/FesvnBA/BiRChVj0nU4qduyLX4nxu
FVIzVqvQxr5FTesm8UZrQYQNRE9KCPyWq19ZDcR/OMtidSDMpeaITcDB5z0ifqkB
pr+2mlfzgqO04Gn0IALy1saHJCgGnzUeMbWpynJoqSOauYabKR4WsJd5Hiy7idu0
QltjaKni3mJparqYKaLhDTWW+5fhdA1U1xSriiO5Qxf22lrMn5ZGADxBfEpK0BRS
kNJltzBX27lp+g1IhxYCU5mVvFfPq1hb14uH0IRloYZnXTSSiOq+wwIz1btUQDQ5
kjp30OiKsLzPeA0jLyK7TYv2/6Akc2nTw/WZISBkgKHUrTDRxFNZtd0+XSij3GQU
Ju43i3ywakxsav4S8lbwhXfUEAh6iyqhkFg2pkY1t+xs9E7zXVoGzNnhv4bGiSCx
tZK7qyJZOjPjUA+j1rkOGHz0k2vSLmz14cML2yZlklZlGiqacBfMU8HE0wijuvht
5xkstuRQ/0ddUBycK26DN9J+3i3TpHiUqQCOhmjjxI7MJaPuBfK9Lq/bb59XFCt0
lEk1NgfYWIxcy3Y2jQeiFNrP/wQGffJamgyGFYMxdZ9IvQF8OJyy1CqFwZYcSnrW
fUzP1q5CAVRnml1y/QDhWftstrIxVZx2hL8pppk2StQBCfXb9lcht4hvN91DraSh
A/LbINWFvsiSsqxdnC61M6hjZ8aN0umD15QkUyeD8IRyyTJBaAlxCotwgt2K463q
RXoQwefL06agHgzQsZ2UcnYN0yekcA3JZoLn+iRy9qtCXoFpWHy8kH6rGlAOeRtA
PhZKFCEZh+rR8nE0Z1LHWP8Am6OGdYpME0J7JmGjj8ortTodVMFT4aQ0pCzG7MjR
ueWZOYoKcIJhqFA9DRe3iJ3m+9NFML0oz2drf5UfW6YF8kqs5OsQzmC+DoiLaG9z
0MDdgmRVm5GSlPeNVZT4GE4m0dhZOa3Wj4ynVBBARIxT57zyg/syzkHeQLjnVPfJ
pwox0UsO0586jxM5uJD0Op7LGXRzVva8s7zDKenunvcU9n88EXOetA5CTUBF7Sop
GXBFpu3DNf4rxAAQ42XpCff7ddWCHVShNScW06dyjYmR8vkKVcgaDvDSNw61csg7
hjXMX7QmrpmVciU6xSAFzWetvgbjVZTQlnghbtf46ofDV3ZUUIfO1paHJYE60l84
yYMuZK5USgeJYX1C9YfgDmsXTBRMKoDGIvQNqg4mMjh+GCeAPfcsi6va6Zb4MWEI
8Qo92xssuGKYU7a6ZiSrgiC3K4hQYy3zkcHEhmPRHIYHXAthJbrKfCGwK0I0OTno
MyTJbcsxIpGffIxwSc0mhxSW5GIyuRlSkAs20bOxUGF3XN3Qj1Y8ymTzBOX9XSgz
bxkq2z2I0uY+cllZ+H8PvrGtv4xJP+rI7v50FYzpR0Uc4dFuUqorvLPG/koDaqJ/
ZUH7A5tRpQzt35eu3CHwhuw4F+T+VmxsfS+SNPAAUlmFQBM4KdyDqMiSUGTK4p2A
2hIlNAMxh5mw4PjWb8wEWq1CzvwtNUN/WoSe+rwBVQns755qMl3RUNfbCyBkCECC
DhyLqZdVbO2k6GrNbJICjb5CKA2ps2X2/R97jtvjTETCNcipGgyZNNPxgwvEu1DY
FpjojFeVRRfLYTAzleD6G+JoGrgBuZKYOLrlwfRbECPoPnWrHUSob0h+z6FShUyg
GqbHjxNm+udwQSGusFGXPWIz8AnXYGqFDGOApWK6AFyfUKHr8U10z6p5A9H8lVSB
veLX18W8kRqwsCp006fhjm3IqRjcPwLmkNUUDFAKn0i132NW53UNaNBBEvPW3VKL
tqcd5VS4NPYCUqUy+r/OpBLie7WHBjawAUi0zlrB3fbsO1WsQr87f/87dDkwjqQc
WzVVHUgj7IzaC+1+TessH0HRJ+KfXLAUXs+2q+jDo4GAw66rlxsHOWtL6b1f6tSY
lmTfdnIWPFrzPr6nTR7YaOZ14poj9Ctx03m0kgiu5ax+OqHjC+qEo88RgV8nPLWi
LV6nmRbhCqlO2ButeOakUn/L/+a3S9ImzO+7TGNV0sy1PYyc8BHxPs8Ws/e515Jd
tePp0HTYhmAWRDdS3r7YZ2fS9JIT9CrF459Wxie6aJ2qh1fk2R5K2iQNgjJQ535J
UDtPZORnTPkX7o/6+2gShbL3/iGqPTjgoJcESPhMdljyBy6RjbkA1PEACleTyTkq
/D2aNJCY+fEx+ZV1W/i4P+hVayCzSMK053JOCURfvtbQ7Y+wpnAtCovsdR2xt4Yl
w+vA/0defmHItcSrejSJDVegHuLPui+7l0oPnZvMWjyBc+E6h1zhv5BP4TK/wYlx
+Icabub7ZsFnsxNYV7M6LbhLlnYV1oVHIqcg4ePkub/mavyH3Cx3uU4GOUI9WuVY
lxpWM47VXYppHU5a9c+OcvcBNrRm+lYPiw+09bG64jQRsPtVxDaG9jTs8IbFDg67
3UxYHqwPNdIekgE4mPmHLJvRjs+/T7D8WZasgK6qDzHIQEcuuwU1B4pa9yiaFjoo
vWkwHkwLzNCgW+JbMXTJyJywjadtXlN212aMJD6Yrde3162lNmrKvQSl+W6QTp52
lFTgiAVTRwCItoxCd/RwWzRsTuVq88G8h57swB0L5j1aggwLYe8Uk4MGlRtPNAfz
51nURJ3XZP/jjBY22GfqsJRAJ4h2YZbAyJQGObXHeVqBjLj6Pw0tJHs8QCV01wVk
H1CmiGLUEHqRvJBbHb/c6OO11Ivswlt98WdqqQxL23b3G6ZzuNteGd67N9XJ9CQ0
fonqYhhYEGC9D5oY+Mq2exOgN5M3VMCCoHr7UmT5WR9yk8slJK9bEI3gzdDke7h3
Noxv0O6SGhmv71gnXkhmHCCMXKddLT1U5mlYRPnyWdxtrT9N5RcseUkR8uDqj2z2
swfg06179Enjl1zqOJoyJ10S63wxgm8BUTWYO/+uFWtgufBhMbh8arFtSoSYPZzw
IKmIiZF92m/6S85iAMTmTtS/3lylUySxkSeAW36oxMPEj9O13w1LHw5nfTVY2UMm
e38mrmSEp+azsqlSOO/e/Mo3FK9Hl9wDULC3c9GsgymGMQ5csC8oWXWCau2suvC/
cmKb1siwiymXF+Kzz2NmbR7Zsqc3nb3v9olky1d8gvPY75L5nKbvs4G43LKWNR2D
eqfjiPc2xJPbDaDQSiblMye+Qz6r0RIpJ2HSMqqAyQj9KOEjuuAk4sCIDHWJytEo
EgterAgZNhNPoyUhwi4Aq5dK0ocmRig1+KG0To/nWO/ebAqGDEXY79RhXE19EcOv
GIO5DKayYhnTzDg6Od7OQwH6/rMoqBNM6HaTZtv7SA1nV7C5ODaCFzQLIyT4dqK9
0m/cULvaoTLNGXNIvAFKa/kbiug/qpUP+AA/Vu4Ylgmk6b8pDf9Dkhqa/QauNCD3
5A/OI6sjiWMV3VfypcIJrGmrLA7RiGkeH+dflmPD6zhGtLZG76tbV0nxULV3tR0G
j03HfQ4Ift4THpmorapu6wW4BwoLkOQCdcve1yLv8y75icnIIySxc5Vub6+bfmHg
96iD7D/KZIVX67PfuBSJ+Uw1VVzmJeZeIQ8fLw3lw19UpIr7RKs/BNHR5KqSZuGb
jeaVTNToI5F+2BcumzADBIrG0W5xfvtJSsp5Gl+mM5ZrNaZxNRdHr1K3E65rEMPS
+8nXwVFwDXy0r0w1Ms+ADUA4mCm4HPsMuyO/vuUmkzphQL9NuJ2yGOvdseeQemJ6
paTJb7Gses4YmyLqXjWcsnJKePAr6vF3Lq0fpO/Ga2NP/1e8D6smsKQPXKapKvB0
P9ivg6LHsQ+drNefWc2ATB79tZ3y1a7xv4DusuHer5JaP4mGp/NW6bFDTrd+rU2V
6sqQ2hleGl8ysUMho48HQ0MIVABKILiI8K7ReH0Lwut1oLXBlSYxsqa18+zlTYVV
f+CTYZX/5X5JNzn/4vwIZTJqstyFGW2k9Wk9d7vQJzFgxDQZVAyzzlxdFtbLps06
EYobKDfUKuxCkfVdFVE9HpytEQVL/Yh81oJkUA87s/mUanAoKesllWTtbbrLqHUO
8pJmop3wm8IjHrDZ2MO1in0TjoZYB6vXCK38nUZ/53qsl+J/ice1eK/fms7Na79s
gAsVeQjux/mrB0mNP8HDLbZ1invs0kty3ivuPigyNsKvH7KQOTuk8tU86YL8rh5C
pYd3k8TP5/7Zu6MR9I2hsKMQL7rPx+Kjsf9d+2EKlRFwZcZC19+1ymg7vf9moB72
tDDKYLXT8jkNrsRQdTzOrFzFwexyNgqCjnlppOV1FO3nHsnE+N2hpEw0gq/9iJXz
EUD+3NfmrTyfmA2kVTKDFWntIwdTXrGUNvZiKs/+GoTUFV2Tbcl5IsXP2S6zkeHc
kpZCWapXFZN9w97qSpx69hWgjN1o5sQqwQIHQICMARWYvyCozGQ14Rrwd3pyLBX0
90PTr4L739fEPGV3DvakxTMAQTalHDylfAwbOMBsCeQf3X5SL06f6Mfd9V3QS8bo
CGXiikU9X4of7ka+/LuGqOhYvnXtCW0QfacFw/XXvMy2pIkV7VkMFfkVXVVUNmO/
kaPVQvcFxr1kbMK7bdcSZnjvN+/5+W9pYNK3UuX/FA8okhSP+j2XIXICYBSJSdCm
zSb2OFLbd5S1ryEpseFyReacW6MRidWoulTaD+Q3Z84Yiptv/qKEEn1Sp161Sc8M
TGrzrdvf+5RTWCLWGbOtExZN9JeJy3nQGa18wM5492LMSpqrRsHWp5qC+A6I5FxU
Gco/1eP1D11exGyM+hLvOe4r72H4GAw3FJ+vuTDwwOh6OwsGXu1IbNiR0dZfGXEJ
JpUTRKkXQuicg37gh7uMUXe1zrqzq8lPBCNcjDW9pLPiCfAw1H+/aPG/N390IDQD
lP6lniaDdWWB2LByhxoXgzDx8cl52yxSat39TSh06Z+kC6Lo5x7U/22tyZyRNzX5
eB8HnzIRBQtCfD0lrJY6+NVCvdSFE5YA6KQ8F3Icg2cSlNWe/wyQOXylq9r3kKyA
ugC1li8CyvGArXwsknwwryW1SbTUve0YMZUiKu7CeyDZgMUeCxyb51q2WZx+Tr1r
Tx7qD288jQB9OWCvsWQ5rKht1E3QVqg6Z7RHecME7UF1Xg1ycwuIzIW6uVv6DNC6
tIYB73EY/x3RGMfr2TCtaMrRyCplvEvXVtqWASZCWOGJv41Jkim7BxGlq09MMtuh
OF/lKhByLc8gUBew37eXnhZJ7qxwMYmyhVc1ViX5Fy5bp4ziUk2kdj3+0ALIdQHw
6wuJ5DluLS/3efAc2DTnTyZqLZLDLH5YHfvFgRyJxkH6RVnAtJ086ax7jwXlRaf+
uJYIsHp7lBnZtZBSolYqDC58AZkxsS74G0P17PWXfNZUqnD2ACZhCfGwkcA97NDM
usdZ3u9R4WbbQOFN5UApFsfyuxuL6EU01NvAb6mQVtzF1tCCljaatdmnlAjKl10J
8eE2Fvo2j1IM7XLOZcVU31R/UHiFXsY9DSGqgBJt+YWwrLIHibw3pM2VUNRIhKuB
eYe+gBd6vaLbOICXJ0jwgFwzNmK91Awc9B1OgmgSFDv1qvH3huMk2W/qYQZXNgkx
R9WHBoMAGSYCryCI5PrfuaTF/GM25NYTtnTlmYQ2+bzNXuodZHPQAyoGJdD/NrgD
pTI6hxoK2godfThanmGtGLhnz460zzwnXhhUhpc9qC7qNxVo/lVCLJ2ZehPFM8W1
yqjyMNXpW8jLV1OM60jqvM7kht+S71ooCbYRg4gLHmjf3d1gsJTLolFWSiRGLUT9
5ahtRRf8oGU64hIgIztWVlAVoMagUKtql4jEsXRy4+Kcbppw+49fbiz6lkEoPE7N
/kuooQG9AEmAm3xoYNxu84U1t3t/W507aW5JCO/VTRhbmOnWGTyRnVDFRKDGAiFW
L2TsLJQjRb7sJYm7rlwwwu36DxVvDrQUezwfstZcMW8VIDlrX0/Xw8gtaxgY4DQZ
DB7psFtAupC/mW8blnfK2jm1GDHgkhGMmh1TRNQSeN8W6tnxNJ1g/wgG/taSc/Yp
501quBFVhDp7eX2hpuXM86jgpfh4kt3gfgj+Zmgxi1gIJhwpGUidDA03mcjtldT5
2YReDW84cf7DBv+BnNgslK0CXvpr42UF2om877MaatIwBR+zzVthWFDdeIQj0qdG
46wl9cq0bNPCyyUtMk8hM1okHrEEKsn1Dy6ZXifLRBwTX7KgnijMWtj7SuP6GrGb
3y7ZO7eEd/OZAndZG6wXQRP1YXBPXM/NCqtoh+AX7ioKsM3kJJngenbfml0qYM0d
F7tZkT4+cf9UWPDzCV+ggAVnjjFh/IECHFxuNmGtanXfWUCKAvMFib2kKyGFcjP1
UpRdM0WhFgbFTgjHFEnziQbKzthD6/Wb+VAl9hnh1GGR3KcgZZYVMJRPtITr3OGM
Nkp4+USEtQWVxnTqMUbGYQ1xNbV5V5jBaNgNENcTBpEbA/o9bYW1VuEGW6O/Tr17
HiQl2cqwCbQz+uo8wxQr8lSuB1pb+DvHcRqydfoW3BbrlzP2KJAVelQG4UFEBVdw
KMTZZYCRgAfhAAzKijiCvxH7GsE+kM98zbjo3sN80MEoYEl6tkGgq3ndrFqCR84t
R64vhgpBrUJbv4qDWFhKxeArlkpXlf+jhq5DH4A9ZSnXvlbJlbDvu252MsQAPt63
kZeL/a939eYl+bsGNLhWEUNeZj3IpMXBOcEb/h+1FFE0BOkAL3w8weUqTeD40/e9
VMRuu8MKUP1D1QX2E64B6ooC7lqzmDpzcGJjNCHchYYUSx8OM1uL7OurppoZRCxs
RGK1rFLWH9xwX3cQ82K6AoaffRUkbeYv8CMmaZ8xyaLoPXz5UfnDUoyjvUCd5pyQ
de5sBbusAQantD220KVKmvwzKs76XGgsPPGTp3j4PS/Bu7jf+w4LNGsZed/Oditp
mhCY9ubdCy7tw64pg3dPcClmcb3Fa373Ff3WDdtEivJHZZq7uLFKLzoU8aS8ZmHE
8/UWJLtt2f8QB2tZ0ayVMKsZIKtPcOqQupk2yT8h/1aoD2wc0T/LQVGqeVN9AI/+
9hSudmcZX+klozy3Z7cxnDIlU7P8DIRlp573YOpMD3b/RbexaZFhYsHAXsq6lYYZ
fNx8Y3nwi7o8OZxYb3+hgD0NEe6L0duXPVuhiTNZc7aGjefogK/sOpxqEvCrnxR+
TJWOggrv4LI05sKtNaVKmcNnjQSnuFv/uigm6/irK9+QyZ31/faR1E1n8S2AA0J9
ljr4y/djjfmfGU2i+J8XCY9NmL27whk/vgAjm+/1vJH/ABSHb6pKXxyEFq3jtD1R
MDUWX9DreezqJINJkj/eHvONFkfR75WnG23XEgET8WRgSHDxLIcitx3iXVAxHlxW
YdERhGmsJJnu711QHp7oKZK1B8fKV0uL1oK/b10pOR9yUF5y9DXkyrEozKTtW6cm
YAo3phSUedSIm6GfU74wo8pAxRjGBVsZA2P6GDWVZEj1eH3JHd6BdmONiSHgkoQZ
sQnOgctSljJXPnh0XnqmVbwbg4xrdv2cpsrH5yJcEywuOo9WFhEm4QkjkoFqkU1P
RgY6sPP0RV+6eahyvJWKQ4Nzv2c10zGPvVbjps1vhzIFqMH3zuiimgq2gW8++nlV
n2wQHkIjfTCNsjUhqM3j7daBU0WIHqABuZ/MDWI1TUstRPoAf6KswTT61zW2CzBV
VYGTKzm//j5zVufAQp+ItEHC/ZwKqY6+eW/uJzjSAz9G4e8TW5LvOmGaQxrNFryq
nXizjvqU9mP+8BzQEfT6cFnvAErb29KJH/4HOB049WSmE957bts2jXdVbok2WM1Y
haPpxcoC0Q09urCzCiJZ0hYrH7iyLQTa6P9AcoX//Yaq/wdOB6o0EP65Waf1eDS4
23L1LO9mRdrESk8qfUErsWzeruPlmzOchkq3S0T9lFiZ3P/wuBBqvJluFfFiLyze
PI0VmWDXUr34cwmxe7JFscn2OZjaw5ons/TVDOapy3e4EdyP3a3vP6TcGeb5jalF
zFKwYHD4xCelFjByA6DEdbFMtMoOWtx4tfH87IH6kSR/mGpTO1/vY4KIWsin19yO
6ayYGX9mEAq5xaOLVedl7TpKp+14o1bOaxSXQB6OlvybxhMdvo5OG1EthgCLbgzk
+PoxbMEg7Rt+v/Smn0v/FJIYm3Rtw9bRo3xIon/I4ZCloUiGddHiOl7tfg9zKfyo
7OnirAh2F9fVOhkteyQF+dyTxCYkozZBZsclSnz7ngUiH6btwZ8+omKgV7+LjkBh
8md5orKTXir7VuVxuIyTgB8K0EzkZ1D8N87sDK+Nj/yPl16SAq0nIXl/tGLpfOXu
F2+BSTCk/PZYKzZ3pHJ9S6JlOnzOH3brt5zISE1yMRGHxFxIRmau5thaouVxYbcx
S0mSU2ijU4uH17iO9mUKDFsQ1+M8VRjFErDKTuanJXcQ5ud6yw7SqxEFglFdK1d/
LD+a7KXLck5yzg6d3BGnZhUhcFgvm4Sa+qPBMsFoo2iu4JhBG49GHeN34JT6KWcY
BaZL8WPNiUPJAtpgBYhGzPP+XSSdapya44iWIj90n9pxpu5tIAO9RZNI3HlxCV3Y
FN0+JuVkYj5ApN6vq3Ui42Wh8P4Tx3hZAh/c8UkaWNwNlatUhS6ZK1LnbuVbihSm
H48OlZO131t/PZ1vOBZOImY6dMPmo+SxdFY7nV7dmwwisBOx90GeaC7PAMSsnLvX
WX55sATmnRm9YPv23yg/9wsq43YDcSL7aZY5J8SY9PKKbeFNiRS06UEpnO9fBK1h
uiXHYzRdDKRQRqXTPA0I9MLMhJTQui3bX1OwwFK9o2Syhg9v3LWZ7fdyFlwTw+lG
UAk6wZ4LIvVtzC5GwAiqVbsptncKS8I6hRzMmHCtmcd3nF95GN/WOPjXKH8+u7aT
62+IuAIaGpgRq2lQhA4SoPAZBV3L9ACNeWzgjB67ln8nb7tOeuFS2/WV5lg3EsOX
whVyk9yGBbZzZkHtfZk4Z/LKqyQxXDm9zo3kpCgsWWYu9zcYX3U4+4h8m5D4duzM
vgUE1QcDHPGdnI3PJr9AKi/Fu7PoOJ0GXdPPHcIfBdBPlfnyjNNzspcZsg56MAEm
qfc2xsKVK1HdX301u1yTrXf0USzgjWitRJge9UwxWCwffHTGo8MseKwcfpK2qA0y
/y09PHrCEODl/739ka9dveHZVRZiVsIEZC0Ic+swg5m4Ph1duvDBMDpL2M0Xi6ZU
2u/He5scUo/5EsouGg0YqlcRsBRuGDpdN4xXHQa+EbWDNPY8JcpPdZLI8PHUauJJ
gXkWjLrnlfozQxGPsf3rMmJci2m/BguziDFCLXQZxF6VlLdcQf6m9dYq7i1YF40T
y34xqBYkTMZoDq5CYkRPE7fC9D1QF35GxJ8XNiB9eYoxf1wSV5Tqp5UQoigzoyAp
lZ9fbkFIKRPzc5sGX0RzEbkUJFhk2bsLmjvpSwBgFxhGl6+4hdCl2rAvkXdGi3Bz
4fxvAPCIhvTH1szGiU+3CsRvwDlqpnH3GSEc5ET0Q5BVrxZTNmvXJS9dCL/iVWsb
GLVGmat+2m0iy8HmbAF/PZcTyb9XtO9J2aVRDiyqH6wxfjKUSX1UcP6fbFbtyhOZ
jx4h/PFug1ww4knIQsf8QjeJAuUcYUMs9qtYknSXetRLFpMTO6YIxuPyrDPF3t5J
ExKDdwksAnyzEtEb/Fe0fQOf/tA6cYqdvaTiBc0o8bllYOF/5aNGf907io7iv8en
i4cHDMHp6+9tesApCLaF3ESPvzCVUQzFSIj4S70/yHePiKKtBU0qryGT3ocmwVfO
c0Z1ATj4EQPsl2WikXb+uRWpK8sMde4XQcQD0e5UwL1s40R0mxTrA6hOkt41twis
IyAN3O3JYM4S//N6ckihOZMi1fSxfPdKBhBUr5S5fBauauyzvCJCrf9s1gHDvZn5
4oKDtq3aNh4Gie7zsF0pZRcnPllseWgxf4Xy3riL39OL7gES8Eq2vLZv2zyFcVVc
vPsuRvBXZ25Hp5qMryc1pk1NVWwWPHYxTcLp+YvfVPzLtuQN43nAdfmllmLH6VAz
Ry6JtCBYnjnv5BRYHtM8eD4fIRbRb/nkJdAYsLUu5GYLqrdXOgVbR1v4KA88EYP2
vUPo6uzADAJ+t0RwgFCZq6nP3pj4gEXI8P3WdBVBSKpeEAfzZppbH9TqCBSIVq86
Il0siveMrF1PIdNa5Ssp59mlta92ozVrtU4oH+IgcxGwrTkzTHhJ2d5cNeD2A7un
Ra5qY42/k/litaDgEw7+TkPtQBJ4o9988Nta1Mrw2eT2Vd5TxXZXNrTwXI21kS4a
idFF2wD7pKkImQtXnxYNuuwSsDm+5EXqBZSIxVkcKeds3sUhDbawIF21eHxzmInE
2fIxMSlx94IpQp2L5fMtLNfJ+zX0nXJwRtsrdCO2LpgGXDuI0WgQbIfJGRs+DbCs
fpTdx/KtS09eNNcT5y7uBwUzu43uVvErf1iTZDp0NwdA++k0EAQ7b0fqoJBWUpEZ
7QqeC0QVAdeGOPh4cev2CS7RsrbtJ8wBjHuFI83SGVMYNCbKniqcDfoRa5S8s0iR
VTTXi6U1KmxmXGqm1VkfsOrEjqDssRZrR7lTrIEVlCUk7so7kzZCQuTRf7WIC7dt
BzLsNrWXETIIdTfnGJTu45oZBCSrdGfj+G0w2B0rAsGWB/frQw0Y5QtTLtyd4HFW
yeZc/oT+0StobkiDfH80k3Ig40Vk+/xQRJia14GpsCXaATiqJm+wUGj3fCy9vN/m
WmBQ/hnbsGT4cAh6+S1xkM9uo1HY6dxV5RO6+lXVIBIXqO4c/7klC+TKCJqOLPlA
3G5WWBhhKVNywbh/2/UR7nUrj07XBduDJKaLKkwo9DA9SLv34ICt2t2iFcjABXx0
PM3xUuRPTsrsr+2ufnGYvPxEMsbwdXqsmsmU5m9zVl3Wt5z6GSvRdijU1qR+OMyK
GK0X789uglbRlzY1VFFcZkB8K425RbgtYUlMPL7ArMgvUKeC+Ksxjl+Kik9UKFGX
bYOPP30b/OQ9CrT/ErvUyk+Tnq2B7jIVSD+8aAZOKeZuG7y+Pe18vo8qQGtI/wkG
NyR/zEiwNSdGvWigPETW+x2IMG0sI/+XmX/qKlJSvMJCkXyBDmP5Nv90EbIG1bbN
5CaJsOHRONywoDsv+xUf9q320ge040DV+wwTM4WKFT3A4ioLrNhiYKuDCIvRmeJw
GNJ0fFLkQ/X5nYS898awfIO1bGys1XJXS5ryz9RnJS++Ivbjbb3mjwGYZWJxpfwx
dRn6Iw14BCNZJgGMD7LXXzLJNT817PKQpkIXtL+wuHTErz+gvYTd3+8UpYK/C7P2
B97l7DVz4cZEJC+3UFXpjrP9/O8Vu3TorAfe79Uz6mRTn0+AQoXzeCTzU98J82KA
7UwG2uUfGp58CHUbgUKOrpECEjClbxSBNl+QN64ZWXYU+bgMX+MYODXEe6mHSCpg
IsMOA69yy2lW0PwYjqFIXXDER6kd6myxvdI8hWi73cSe803f8vyDy+YS3iwXwTr8
ZTA8Xjm9GY3d2RpcVtZMwbCvwT/aquau4zlRy3r7TEJsO+5K6yQKVS0QSvuW41qf
UF2pFFDm3r8XfgxgsAPHoEJyHSyRgfOXeYLUa3Ykmumur7tf+kLtJtVsgFwBkj7t
CMLm+MKmAWrxGnaOWMxF4WruSv0pfMtwGEhc/XPD+YVfR6w59Xd4pHy/TmvFfm87
03vqaU25L65tdJaMtFxOySVGFrrMIFxCz2h1upHeBQxqVAPkStzf9V5dL6R5gZel
L+Cu+7SwkNoj4ItJGuDziRgVvWrS2+iLMkXDlc8zP8KDKaXcBPnc0Yi14VfRQHxf
aAYi63A5FEZ8XXkien9Z+reAkE9GmuzBEyp3Tyx1SZhpShpAGw9tBP4DXicTqwTM
KMWMZzm/BWs9StNUNWnVpjFaux3cyuaK+RHzCz7EwEo4ycg8U97RDlRYCCqsCEoA
qIpgu9GRbGMwJz3dJFtdDccaHBANe+lAgl6mrdCGr+F+QsPPr0OCVOIwHytLfZ0p
WackMJechyccrYRK96Nwna8Tqxb11qqvIaVUX/5LIsxvc+Mr6cmd5Hs3YNyN/ezh
4MYCrYJYm4c1+SusWpPLujzuYzQwlE6Rn9aHEJ52iVSeI47KvsEhTWVUZnOlk6xF
j5vP24qZt7PgrZH5xzr4TE8tlXJpaj2kSNpxxj9XItnq8lxK1VCpyzAcl9cZ4vUP
VkXcRbDKwmG85fia9/xyJ6ERKTRlaAI/5MwtnPdihTpiWCeTlto2rhxZUeFGnRH0
QAKHDDrxUdI64ijr9cgb/UOvRNXxrA5THKRVv1kzjronOWqLnYZJ8StqOAxXodoK
LSLMHMzNqeENZAKztlLp+UDdZ3AaWY689zU4ag3d8vzL1u4Imn6TpSjQPw9IoSzF
wUgWAxdwSjwpPMNRE5R8xdGeCYl9oEMItY0gAnnSpKa+QgDrji8/4fA4cPPKOMUf
oZRyE4Q02F/OdAcIZPETA9FPREu/C4c82eg8MpfeFmBfQeBoHLcOIufb2a5JFf6s
GSTDK+es6nBfnVkTiw87GD9wGaATIXcvfevPCyJXrAslvWrZ90qsbb6iSgj76gsq
frD/y+rHHPBJDkZpU1WKN2IvY+JLeoXk8l0LzDaQqt6llsVnUBJtv9Ll8tiDVSva
M9qD1oglRkuin7xT/pc3bDihRa9p+/Jx1hqJq2gmpRNHelh3NSPcgf8QVFEM/azB
v4ZTnqVv/Dp+cjqygMoO5c+V7SJC0LIiXDfLJYb8Hfs68YYtAN61UuGP5K8ovBcF
sluHbELFjugAlwnDjvuKHZ1OCNGETclo2rJlVNfRHQGmg3QGbeD+TEvrUQnGXdAT
eXDqqvWdc4O7VNZ7My5cej4rRhsavrIK1HAI2ECEybrebjcGwumwQEGYAeSwQAA4
lVNPFGqS0SE0eGK4L4lJrSVy+BMbKic7Rx9xJP9qNvQnEwMzNuYCRi6Ic5zR8Gka
nrDhVWJTXQfsdFpVVyVreo5kdx+Unoia2j1oQvu81p4kqfYyx8hEk4dhhhpLJkdw
AGXOMOxrH7xXHrTasBcFROVllsozsf4XpW6mxQJCoSaSB3OO3eRgu7I2RWaNMWv2
uqDA3haOp6vjRWqZ9FFGz+eZlD2hzvI4jH9TV68O4qK83J4YCm1p6u8KpYmsQn/L
Z4R+veFtqehdRckyrP/uK3lcELV2PSJXw5p98twrZyC4RxNv9C7pOBbiAFn/OvFU
T5UKJWwH7U2Z0z4Hp8knOuL4tG7q4AqneeFoCsfvl19IV+myDtA4KSr2CBYQ90qI
t+mci/VnAil9t6oXwwjUuQ1kAJuP+XwL8u2it07fly5Z7Ck5MEc7t/iTU1KCw4kI
NTpFXHWNd6IG5x/88T2sKApcS1rQ1ZZhRKjKefZ4G60hnZK4qknLsikKdhgiobZV
9qy+Vl7tBZF72Lsep9bJFckFqisWhyWt8BAnMKUb2AcqLpr5SD8Kg2bdpuddqRvc
zYDpfueUqUDb1W8x36rVj5STOWGG1DzL8KXEQaZzDE1BNuYLo+uNv3Rf7Mp6Sjjh
L4FKr5w7QIcYXtGRhL+L8+K/u2O55g6izl3ZirCIh6sULAAcQDvjSL93GGBvXeM2
VhEKUiBpzchhDZoaJgLcKk+iQI2Qi5orQqWwk93M5bBxC0asDD9PaMveN4Xi3UmY
/Roljz1FgZkBNmf7HwkDT0vdgN2Nur/WMY+jSZiXldL7PYcEAgZUHa1EYFNpfF7V
TDLD7q94nX8aMY/A9F0rXGKSvmVH6KKRvE1Os0bemn438j5iz1T/r6UH/XleEdFv
0HvKLt3uHqrzQC6yHb+3jQ/flbA3hvzX7rEocys9FSXps7dHUXYqiubT9H9y73sU
piVh2i/jPhcMiNn5TjFUFL0kronApRrvsqghSJsRvkEqDHdpxuq77+9sQURWuFIM
1ycz+R1tYTC7NS+3dzfWXkb7bRZoKlA4ru9nH3tXOIiV1d4sLCpTFfnIfvTzFCmi
Dpryg/jE+pB3sjnriih48qUtdHwMF87gn0oMjVVQSE82oC47YUkvx6KdnHCErGsE
sJZVA2MpN59GQmNJkaERZpfqvWgmChF5yuZzPLCZ1ZgjQ+DNFWWVAsftSQ7zUMG+
9vvq5FygIQ8wlZxK5ABd/MbOZVuxhq5Zyg2V4O3ELP/mi9QglchN39C7asUEYfWx
yNDe/8vi6u8DbeLcEssaSUuZoLjwj2ojguOpYwdHsB2lzkvtgq5gqtcoj5WGN98H
jDLEBF7yRmc+d/8y0DBWQWFWqxbFj7rYXFnTh7dcXL58RaiVGIV1+sI2dTlQPwKB
8jFNfpfPfIkOna8gQ4yE443f4UcB+toKB61wgBMq9axnnibDYk32eGZ9JpQZGpPj
wJID6ROWgZzA7SVwSZH4PFW8P1y56vLdGfiZ22J3sZYgJXOSqbWC6qIEjPKrvNWR
EifpmIjs/rnPCoOWNUAAGXLUvYGjBWWxnjTwyBwJZUk79mtJyqjAbLxD4ZbJGE+K
xOkl8cd8r1QOj+zMSvtNvUasq7od5ca+EikXbLvLPGd9gslJEIqPHmyE1s/MgUpU
WSfIlDA8p8GLfyie/vtyI8VnHe2TdmkZC7aXTJ+/0qly7dOVILSVPT/tifcUo1+b
LqoVkLOZCBWfi5VN6Dc7g+E/mjC6LSRhyWrF6SLbTcnFrOmBu69hxwqGvn3E0QqR
NaxXU6oQJKK7RjPQORARwW8uvjn9foWxncVHQ7iufAzynFNbYm/WuWGvkTS5OkSF
sUuxny4B9ZslraUNDdFD0X79Tq0Q63otV819aRfUd8jNjHSdfUAT/dqOpvAEwB9k
KhGzNZj+C5FmpnZEHywUtJPXmL0IFzsisPwYSn7b+/tuaAUs8iwyBa4xFEcfVkW/
hNXA11uztc7j0cZyPhT9J6BlH4sBZ2rveQPGZjte45ijBk4g3bu6RksEUUEg03V3
j9qIZlwrr8rqrZILv6zaP7ShiopS+Qqb9jNWYLZbqDiTokjMOilMCpqgaw3I0JUn
ncTNq4zuFdBPS2lWe7CCzw9MICJ4+oZC00Vt+HDsMVlre/Tu93wfuzGvKkB+uRlb
R0Q6GmTN81oLZrBxQv+/wlzuYTVxUPB/wcE0AFnqzgei9Fha8HZSKcpc7dSMAsgd
X6eCMBljdtRdfWg75ETNb5drGfpLoJSynK47Pr2qoOgEHuou+7pfMrs9JPYB5A38
4HP9KjQn2KpgAQUN/rhM4nEsZ0laWgMjV2kDyzBm1Z1pVNydD5+f4K9wtrh1l3m4
cpV9MH1GuabaUSiylEjtwwUYZPT5nL4TohtRCKn99+OEMrbxgStWRQJD0Cye0+8K
ExLnyGVrv+HEu1cuw2BwcYNHjhEU+ePEplgEPyJEybxcRaIi+/P0MiDDG95pfjZn
xtaSbPCW9ms+6j2sITAsT4f6b/5FdCgBzBWUvXdPA4cJHSUUrGwqK4qa1SzT91Co
RAqLweH+bzATa/qs1diYPaIlc6ybtyG1Q+S8iH8YgOiXVMdW7CkaUKkzcaabCBSv
U3Uu22ogJWA6U/bIWsneZMJKvbIxCFYP1M/WeFtazfBz4UTrO6penfx9IPBot58y
+KRxusZj0I3TNh04E8xwCEl1g93ZiZ5yyu5QA9MJ93HEwBZw17f5pNbxOWppzigS
WLBh7XNUEuI73OPTYnaAA1QY/7b65ezFFuNtgCSht5KcrpUxPZeoac83t43iM12x
d1UNBK09Ezht/SiSuL66XFWGJh11qgIJiFXFMZ7ztLJdaPqdgqpA4SbRJb0dxPsu
nqlkClFNxId4GyEosy8PmxRpz50Wk0/BCZnTo9MVEHjV/Mz1m0oV6QZ3mDXV1xSQ
xAUpP67n8xMtUlbeYKEoR/BUKkeFbV/MbT5jfIzJ/kQmVYiNSfsCP5hfHIhTUZKD
MIgWZotbl2qMUDnmFHXTAYrqGEeGc/dihMmeOVAw1M/o2M9iLT9ip6bXAGTPymSC
i7VGl8nzfarVBi3CzUjA3dAh62TGG5wXq3SWMBfXgB4x8SQLeg6XVYumyXUk7wpQ
bz0dmhTnMzZI3679i/yEOuGeTzgO7bMDFWlsOKoCWHzX2bnhVQHqPMc+tIGme85Q
fxqh0ZKt1BRLQcArSd6W4sG+N9TJ46sMOw7A12ytmQzzqqIrs7l7/z6p1ZHWps/p
JDdriWQdO29zj3FJxmQCCLq/pJgDjqal0Ju140rMbIeBWpUsJKYh4n7F85pOXp3N
HsnOBTacfyPEcyPiN8Z8flB0OvGZvv6wb9N/lvfxI8odccxLaAggM/WtG8qwbUAp
S4VrNZrAMjNs7hDAQMOGMpTdduFiIJOMf1++MFk/uGuwBBsEB9/dLav2VhWRjh6e
KSbWFmDihBk/PXtA1yY1Enzj74dXWw0IZdbf30O26CMy1IpGvcm8Xq4QtV16GCd3
8nfck84CwTHgb8CLQNvme92MpnMNoFHKgUni0JEMoGSs3zplhciKq8abQHbvfxqS
3q92wp13ADt293uhWhvu2SSluo1RJYRLHzEyUL5NqWGP2XDA1fWV/kN0Z08zDi28
8QT8q13rK2L1FKPlrRX8BxW1B/jQc1fChjflAx9HQidspPeFyFmYqiui8XbpaAj9
ZmVcghcP3G02HwVu3AkoaTNLw8cRHiOHe+N9WC/ToBz/VWUnhZng2oW1TyrOdEfp
OARFZOI1O6d4oftM/Jr+7h8z5sEI9RMF++r9xJ/kcE+lVZOQmPmdBc+OA3iCpzlq
6cxBIxCpi/+vACT/9Mr3uOQhSi5/F5KrwIlK8bb3ySo7PWMycRnSh83h7RYBr2ms
lP5xZMe70dMfggkDAbTzTX/OdSOEKbFiae1w4XVj083lMqKIDt7vhtXZQd+cpCg3
whpYTsviNvNW2NhOpVwmDE/kUVPjwK00xe/IvQuwrUJSByDd2dIviyJPFpC1Q1fa
++gHP4CpQfI5LeA+9HNl3765UsziMENAdmHYCYzQv/u5+m4/AbTY0ilwu790cwXl
BLoNMS78doUWU3Zw/W/6aSVhw6cmedDQPB1usc+Ukg75JKV8iobcrh4xxZEbt4w1
e4TRAjmXxW6CkertTkYwbOu7D7fAXP6DNi4GVBZ2iPKI7wsxHIctcpW3dH4XwIv/
R5AhJYpGrajlqyEAhqLVIxJox7BfOCp4R1hewcmPaKw+8kDy+HT/mteH82dRn9D5
qSE2Z5tO10Wgn1+/miG3Eq/chi8f+EnauzGdI1jKjhV4jPM01SHzLP3gZLhMm2sg
yGz1te4hmNVrZZk4m5uoJVxgtP+gvJJU2b01zZV4BJervQwxxxgi5shEErHc5lOY
gsLQhtBMFOsnwSiT9oi0dQBUFYYTJxlP12c7ZzQI/FNuzSX0q7YwK+K9qqMSAvPc
gGFxuH73aTUO0jRSTNvI13frohmrGcoBBiGk+hGeF3LQjHsVGLCOz2CLS5pIwMX3
3Fnp0hL9TgjRjp3uVGwZPfigLKSY/ejI+tcVM+1Ka+NX0/Qd4ChRuM/i8C0/n2oM
qXM+daz/Jbm2DzSi0nMhzC+/1EOqUzbIMXgcN/y9yfef0eGM67dZeCQU2U0Bieu7
KE8BqTXQPgnzSbL0JfoPmCo0sY0Yr6J2r4aBViykSZijU7oRgiut0HRSBYQvl3RQ
zu81RFFGl6w485rsKEwcn+giUSQ+CNQ52a5ycHHli1Y+ahO09fx1YJxe4/fEEz0x
Sz4ta8GM6XnhinqWgCv4VmOcjObEMw6zU+3SMCKnTLYDaa775rI58lRF6Y8lpd+b
OhIiBeYak2wcbvdu+cCyv7JfVpCwBGuLejj/tGVlb6qw5O7xdStnmLYWHjq+oJBP
Ps9zYgNp84rvpxuTLqR5hMivKMmFH3ona58MAqacJ2GoUA1DYY0SithiOOX1yrt8
o22jZU5VVWKk0kXaOE7WNn+rDPV0FaHD09+dNpguKx9V87R0K4JyGSauIebciwdE
afmbNg06eEqO4uFmC6WixCo3oL32+dLF1leQzSagTTzBFi/+cieDYdQXLKc57JWf
HBdTKluzCSf98aCk+DdIdaK54jFLwqsoDTKbI7a96sIb4ZtC1U3rawN8lZrWlMqw
UcAXakB4zcf1l4tCTaefHFeEoVrQEj2oqnYREkfV3GIivfcexy5gFKUVWEcua7JK
actlVQyhP+YObazmspMwBKup5JOZhkrNeyYMfqfx10tWo1ZINHoMJE6chTPEuQcz
LjrAagFd9pubaj1fI73q3n90AwS1NREQZUsgNsXAJQQzTecy41mPunY48/sK1+4D
5m+1Mjkq+SleInDSkZnyUgYHyI6Tus7VU6ayzJ0WJ/xm7iv6V/+TtBirSwMh4KnM
h7AoZPNICzOofbgI7y2GV7fFBJn0aqbSODbx5cIwYz/FEXPszj7GQPV/nwLM7MKO
/6Pt4viRfKYAy5MKlotTZsc4MBOrORNe6K+89hoB2qmT+pTbKiYlVGKE12o10Kzq
6OwKdraaW6JxRvwOsR8nCp++yT+cQWbY/U5HC7gA5i70hF6WXZRJaerUAbyzooXJ
k2EfFgZa71AxAVZksegEnLTYrDEkiF5eGhEl6RZ7vA1hlyPmc9CNWrlqQkA/kPBi
ocbGfYvU7M2d26760N3T65aBTKP3cvSYYAvV3cqscpUpoZLROqn5Vjm1TRd72nkr
wry8j5XmG30tld5EM7v/IqPY60evxILcMGnpCf9IbSvNHYqaeZncnlVOeqzP9nFg
DvSxmVfnhXpa8+8ehxvKK6A5burVIU5n60xOub/14u0OR4uyP06xjIE7xDHQuY6a
SErq4zv8GNQijN32ruaN86hTgrRVFg9QG52p1OKHxqa4FO9rMRtpYDSWdKBfa53M
VtkuxGXM94yG+N1TGuHr6CKctkjGGiKin0QbfJkOEMCj6qNy6bb8csjrnzoaTftd
XboR1TUTfTE24TUoohIP+16LFKRbSIxm3C7AtccjT9dgCkFoDn5gWN11UggzPYd1
9euKXK4p/fmi4pHZSEW0ixrVQ0gIFSXIdtUAjOtTd1VjnVVUJNHPMX2/bX0nZJ2X
0iwyhX3UeXOYrSIl61VF1VriR0jj7FfDy37JNW0LbChsLdXYnnysxPELl22Wsnlz
Nla7KUoAQ/VfPTQGCqHIxx9X90g1s3Upgg67hpEjw7eqWfXvaIIzNkQfyWXZKJE4
8ewF2VYMuJVBw75zN3T0BAoVqJ5cfM9Aihpe+xbC3rO2Ew79uXAuwo9hzZ4Gr3Vb
/Me3TsSHKRA/OFiWy0/KhGHg39yRsrMFxi2OEgDOeWZ4T8QLQeIoVustVDhm3Mgd
5oKxU+6p9/cCuWZKLowmEIU0lAQGYm+4NNP3pi24IFPFi8ZgvMJw/fMMzP4H9bAA
/RCJajm6q17cZR+ceigyULtMqDmDqTeGp3qWncxHaLqVpchQRkZPdXUaFeHLOC+H
J35bORMJ6eQUYx8Dsz8coQF37l+tmGD16KmxMK1BR8FckrKuhyfqh4kGHVtBSiT5
5mxPrYvzudZH1fptUDdC5cflUO15Wvw9h2OlNF2ZKEn/ioU79cleiTj6huzojnqZ
zMs0P3De7CopDv/O+3O58RkAr3SliCn85T69YLpV6gR6A1RS6VF8JobIoKN9/uQm
jPqt7OPzeuDPsz43K2en0TSSSfW61na/pVIOZDvX4yQ7etUK2etddLEbcxGidB3J
p3jB7/AyYLFc/TPqgyaxjdw/TmtlzpH0tSzDJChrxj+IfQyY10BZpcOGWItPBIoB
ieJ93jj3kIazEeNrcFIJdrrRGldzWJbfEWdkUfDxs1KwH20xatMLZLxnk04xMJlk
vptNta2WDGBO23zLRNkqq3RLhjUTfCSux6TISwqLOMMk7Nxy4HcM2YMfL5dRcxYf
v8Tz0kI7EylX6PMlcUdAtaLR+4KXALgOYxsCfz4bF5qh1MTYWc/91KvShRzf7b+W
9TR8HEQKLI/y5do3cB+XkZq6Eh5uXIDeZ/umKkPcbywl9CaVIFTo3ppHAP6Rm1Hs
Uusxx3sDu4XOXbX0H82D4cVCEJo/jrt8GYQRyaGf0L11XPcYUmXL26zoStE2O3AS
egAfphfkSgAba0YVFpdFbGeVDVy6gOVEsQGG3ZuLo23s/BcZ/zpAUdUHRxNnB5Nf
zkHYP5A2OhbfZSAFEyK61+fTDDm9DTE/a0EBh71k68NN9RnB6Juhs4lmk+pozZPU
mhLxHKivBaKHYeB+I5wXjurJjy+G2yfMf8OFjOXeC1rXacHpTNSpnq+sskoEfFvb
r76rX/avtcSaIlDnJp9cL76gQ2nywT1DeZvqW4oMKNbml6jvyIRo3atBIiOT369M
iZx4Cl7nvWdxphxYa0xEdiM1QDhuEXMdCjKCQKRuvrX/WQO2SWdd2J7XFgtu7AY4
jaG+16L6H/sC5w83KkYesFlqNNhD0mXyKYwNeADqEXq8Gxy6VXzipSR27rktRfxW
ocoOJIbMxbq72xhCoul2xpFdv8UnQ/8/BYzq77muuYkg4j2Kpr9rQ2hTahGEIKj+
WBsGme3qEO5jODnYiG0h9vVZcV5HO3UzAq8k2P5jc2SVZ2tpfTVfe9CKFVCJH/ig
DsCCQOi7JxBRnd+U5eQ4dW90KH/iC1/t+zUfMes/EAeWczA0N8ZuqoY5ILCUSYkD
+N9eRq4nFF3093ezIXjodoTx+fBxvV0BES0NwXzCk50N8ZderLq4Un8i2qwoaQc+
dQoLuO+S+CvbQSOloryXHi3LBRY9nArRMV20vpE5CcjrOt1fkpQhVc4WurEVlA4F
r9YZRgnhU/GoLBmWvEhId3JYsX6ga9/bNDQ7q8QCf10naB2Q/F8xwwXy0uK9azNt
c5KqUCdoznpo7ZzrfDKiIDdZdFGyYYD0sy5k+NVhhfrjK0FqujNcMyLDsAIf3cIj
NjsT7j9P3N6bZckek/ZEfEP76KQabadv1EaCmNiA+Mv0oReE2WxgMW8Py/CUZoLH
FIEThvva7SY8OA2OFQ5ODObVEWPZAt8973BpjTAHvDVZwY7UMcPZ/eUccvvIjPQW
sbRoTnkrWs0yR/okTgoOSDLWNJKzthH5UsaevCAemTVFn7fksZaQPdJGytlX/82U
BWdYqv4feuRMBDJawsYYdrqJwd36KV7rX93bFBlmLP5f+tJgm5TGW1ga+IcIrMOr
y/HNkfPx0xkhIPEJ0JGotD10gXYcNzVl5Aj02kwQHFf0UuTqqmaIyaUrMV2iKvCx
vkit143amA26UAqE/sSzwGwdnQiIFGSPz5Jz5kg3JoOjdRj0raGhq3qLhlbM97G9
d8kllnS/NCe8cfRlfmIxXLoaT/y5Rbb5AFGJfXtSS5ZICugqSyWScOMbf4774SVj
B3s7LQMuYqh8S3eGrLX0OX56791zQ5udeuqlcs4tb1dQl0YtF9pAt/cUPYNxtnxX
yMXsDQFe/agS5wqCAdYsI5obYBsGh5rQrA/XaEGldCFcYacIq+gtSbjStQyV2ePZ
6Oip6qO1tI3A9w6bTUeJr3GNwH7ZOcA9NA4sdRK+jLJGBC2agkWCm0RDj5VYC37c
cO9p2qJicwDzZy49i3kl7syjzHsh3ZMEHcZwvom3RzHgF9IQV9GfDV92VPM4GEWb
Bv23YkYG/kDhpG4zUpu6IzlcR5rXwtglP5sMpgbjDEp9y/bf0QUQtFt4Pg7X/Efx
CITCms/6/wQdTwUcn8z3rnlqICrZ2V06qN5AiyYUYM5TLvmMKNAN4dV8MClYvd9m
dgvu3ucVtYbhbVEpI4BP8pFStMB6A3AnosTSoRoVDUWaNO7jQv/ljGCDcjNTrFiO
K+AJS/q0SBBYdkd+MCYWexurXQqutTA+n+8etrHjsmf0PDdskIX4wLmHmZG4warT
x/e1IbaxYBEfwQPaQZYDCQJ0FRTVD7lRMzj1gZJEDSt3KntcSxINLDJQKjfCBNJo
A67EgtveLdSDdw3K9AmOgBaqHxLbSh/PhPbcaubip5BtTOvX83W2aI2myByARiCu
IumzPZy2NemTGCN1mFB2F+BjCE+z/kOPwk+SwxVdVByjm6BrCTaLSobMfeDChnKT
hswv4XeTRIJt/thIXKSZLCK1RL9MSP2aucpRJtu4W+YqvlRgv5hcTaFUssZHxkTy
qQsvhJCZv5m0B0vprX56EUnETSybHTjDUhKAKsIzttFVhOQtiGn5GI1b136jlGue
l9oFAVRQ0+IYMR4SrlxskCzR0DWzf2pRIuo7qi2pPD7U+KzdmHqQUDgBIO3fk6ia
am4NphVCxf2mIkBu2bfzdVAmJaj5C7/D8LkvyE/xUILWPjw0b7L09xFOp17sikQn
I7hP8DutO3bs2l1JzltuYBN0KyeDy6WMoRIvx3YX101fF2ScY5VOqKFidin5Op2F
8njxxbrOSuQ8k8JK6X5ywt9z/ueRbnt/l9pGXbWnZ/R78ompccM97xTvRafDu/HG
eK6w7ATXjqv8DmP5l22FcTBfJk5yRxdzIDxhs4ib2RzJHG6ww8KIBgej5G7DJoI8
KtLTt498umvk3GtDMN9mdjEnxl4GpMf8tE7OAyxzLFXnX1jzdjUDrd5sSq42tULb
wmh3VF841Z3k40azNSVWRob/LCgDkla/7U4mWM8USHz9eX+RNCa/vgfdMq/3o3vb
g7AfRLKgmIHvwfUaonMx562u4d3NLri4gA12W+fJkCfEBcnRV1yTFmS+AW8EOOup
/5K9cGcAtvb4rLXODEbDayDdrHj3Od01NKZL4T6oIF3QjjYldmJFlakfiUWWpvWZ
9vC5DXQ2mtdY+dM0pF92NUkmeHdCUl+xjxACCoUG3BqEqdSW8dJW3Ma+jBqRQ+wK
mwXCFXr2stktFHhIBYB8i+Z2VVEnIH6EJj9K28yZ1OhE8tM2liEZ4jphqNIhCH5Q
rN+FQll544XCtQz7dJVC17pxh4EFSR8V3CaKRtZ+qBKKjd4ekhBlwByykTmcF+ZE
6DFECNa10sszl0x16sJpDKGZ1sDEPQLLOXKixMlPDBaZALlGAND2guXrN/OrTcg6
ATft+aWJHb4+AsvLFUE1EnHRRY9/J7lW8bpIGbGYxcczx4vwuh9EvPhEQvV2zu8m
QnduTtQeMzT5FL0NQybjOsYWYIoeL5n7YkhvQLmCGUir8b81Fcmt2xykrKHD8vAP
3CQo0x8yXKcu1cm5Pnnq3tHtO1iM2VEtvpf9OmROzqnfchsUj4eBq7xe1OltyQUX
TixHZnw94j5ukzr/0VWQM9xHvGynpO/gB2aQv5WIyhlX1n2pbZZ5DyBlb2pGy8wO
YyA3ILzDbxiwj+U+kC8ejnsTZWBrJ/O9uCeaPOFvzMKLXGezCmQENDZAjVGBWmZy
8cKABLqS61XVrQ76VAb6a87neW0OM8/ZRTuoGqHWgw0ZBDyvbyW+edY3AaHB/Pd5
VlIgpo0ZCK+1Ucb+nDWbw6SZXPSfP0/19HEn49iPMpByKxE9s6HrFK5Plp6ZUt04
b7YGajQrNf9olT/zl2GvsTyivIgomOqV+tYdynEx6CZOtV0PJX+BrWc0PJDqAGi2
uQ1RjqdQAXMihPSDgtJbczAEs2wfsVvqI3R9+i7H1LOu6r9BOuc7KSm/t4WsS4Kt
f5ICxKFtG3M4Ma1TFB8IyTAWkU/+xtrMZ4QlwKFw+KG9ezufbaG9ZRVkkjYMRnnc
caie6DscUF8+jq66fpspj7xwvSRhK+27kJjyZWl8cJ3nwzEGo3MD7FgZx4yk+VsX
4YCaU2A4rlObBcc0d/9rmnC8d8tMYObzDEAlxIXT3bFIaWBL01ahvKmHyHuRycap
XBEySSw5zinZ0OPQc1W47qzftJnSqFuP/aSN4LETjwPrfBTnikKt0dhvQPPUzqo9
0YgoL+513h8jEcL2hn+u+jHv+YzLV3GWwmptZpTIYP5XxytvxF20TYmYWdY6UEny
/3TVziup8qbPX+EEE8QI9Vd1YcHBsXfd2Zx4zYaouUkHJhMs/XdXjC/46Oj6jQKQ
4ucXgmkQ62p0/zONR3vCKOp6tUYvF4NeYDOREciSSTOXZxIElBsQoyInRinqdOPM
5g3RCB+SFOI00R2owMsthQ68msMFuVaO5h2A397lbHz6PX4H3JQs7wK5BGVMBxxa
0Ov7OJ8rtBQT3Ksxtg1z5aYxpWA0hPbFh3LgcZ+3vjPaXzpau1E/P1xn+lDDvnIe
fY8fqwIO1rctIgGWs74gs02Mm8atlEZX98EftrRhiI1zovSrLs1W3m2LXvDTyu2j
ZRBiHB+BK+4dEFnKHISl+dVg2vpxSkM8Qni3eS86Uqo+6LxJ/QikX04URWXsslet
Ivax6Xd3KueLZXFGc/5BYcweM3J48eZ29QMbqhbkQPS1D7ivhDd1oAxIeGl635Uh
QobUsRf4ZXax7/phYns6RZDXE02VFYChLk7n9WvKzMMnGgKhd33eGLbz55fsj/og
Ekj0Oiqy9xZhozOMTC4TQyuUNjeAZF1zd84czXQdoVBkl3hacCuU15sw+PO/HBgU
sDOThLPKZsDGNWUoRhp7z3YZgrdC4iFM5I9xIqJOMVFOvMuBWqqdoITOWlkd1q+H
B0s8bJztMHlISQD2nCagiHLuCv8zoB3VtFO//CXBxhE7jedjiRiZ/j/VHzK3ngGY
YW4gdWwScaPLc9xWN4HY6GSrAsIQizmEVsDid4Rqql3QtlC3sJ7xRAz1A/UfdX8f
IbqN6FC7zlgxXjvyQJj0c0zhx+kA87m79FDaCJf2mL0kTQ1zKqPsYjhzxMB6evxs
cj080Nu+5NBiM2WZMsYp6bCTZwq9QFm86Krr3QVuGIAsT/YbG9qDGqHe1OdgWJE3
NCWIw2z3hdxl98aagXcBOxD+znoWYVCtloRWhtmLjIUl698nppSRzQT+RYN8UJYp
SK3s3tUpIz5BdnAfYmD+cpjszRfu7wNP6hS4kqUM+mI5KoiMz04MRjDGY18yBv8o
pMg4whapzrWSqwqxhMc//3AwHRy3e1pXs5+CymmhDFnvHh1Dlc1a6GAEM0mfy/Sn
gAdm9ratYHLc6JRlx8W3XrwBhYDh0mmTK7XVyCVWqnLok8avMWdrENZW8MbLkpmY
n6xl8PUWyarEDa1jtNDi9XF8OcKPn+Zdyz64HUgupAMNNJDNOPuG2posnW05no04
cS5qouYAlks+D7Gj/sOvxld0Y9iJdtKqjqSAw0mvPM5L2kVipgrRv18U2RDMo+C7
/m7s2gbHgNT7yrO2YQn5vWbSkfmIYAPgV8Mzs4jWMpG1UGJjx3ElYfWGu4eu8VNr
fzKBt6lV5Xp0MfWMJ6enS1d4VNJ+IYodWhXk1luAS/fWPb+Y8Q3nwsdwSeOde58H
25ycQlh1JV7kCg0wKOrq+FC932Ain3dN9iyiZbuM9Y5pBNzQWajN0Zw3Mr+0NyCW
wi2D8OAXr25yem76AqXaHpWckv5/LcLxpuuwjEgDF0hn8mQi/SM16uy6tsjO7c0R
g0Aj/bJiYWGK8OVYPUdSt3SlJvob6VTCTBGLQEUL63Z6gJvnNCNRmCTvOZoHTcgj
mKTzGL4ZZeP2ZaJHLsvQLLrlU5z7WDQvy6imOoimAsLCPmzKv7h9mxl3K1nSRfnC
K3M30K+NKo4fOvRUdyfv1lWb6VOIAfhLMFkI6pJi/IVSe5Gk7u4nqaPwenxnbQxx
0hhwJa5pxg9sitVoP+DLu2eiXUjtDAAOUyOOUhQlWHQP6XV0DBqMskjYFGzusvFh
BC+N9NXjWWWfqmwH93NnIicJMQ8ee1oHBda1Et5bVi8ej9Rx+LIlC7M6bjRJXeW3
bESVP0ux+O+2Vf5zVxeQJJB/KdrN+K+Zmfsnly81dX3HO1nNMheCeztEy1MkL4rc
r+jxRT0OZZ3C1k4hBLDJrwfCFLFV2+3K4LT4vKf5WF3Y7Hsc1sxJ5TdvyLaVyb4U
efaj0PVZI0o18acqFSseSqpqAZ9tYNBJdMZRynESIDdWGmU0Ku5D14ssn+f6UhRW
VW3YcS4eznyhnPNeCwZVzm5qAV53HC3FE3ZgKPInNPpQwdb41Z4KodCzuGrBs+yC
NaegsjD9d9IfhZD87l1N+r/coqWoQdbJO09GCBKce7f1sBPfCcCmZUuuzwdWuTCA
jSbbkXiQI9nVmQTfAq2qMhcX+Nr+yp7tcvD3ERfIEO7FcALjGXgCyvGPjDSkVDSc
1X6yBE3lhO3YakFzyH3rNv5Fu+Qi6W1VFXBPCJgnzwUs0LUMfsBLfmmBvKpVrXD4
9TD1mzGuujFpPYMuW15ktbcZAhlW4k/UBlCp8y2rpSc9Q/Mf1opPYFgVNmmcrEv/
yEyp1+irx9zWjFHEvS+xxZfU6J8Whd+QiV1lBWwA27LUnXrmn7Rg4a4g3mNUCbXw
zDYYDPqhrCt+YhRiyl05Iwzjona70SC/1wGUg1WKjQolLV8aG0ITmyvJbMEO+KS2
oHAyQX32k8bNb+n8vMEU7EdpB9vkmB8DRA/LdG+M5FOaJlOcABwbowYzHitnI58o
faYD3X9xBMEwfKiYlR4jPVjbJQmJZdngCvNEARI71WwCzDAU4iwvP7xh3LFKojDe
RxRmHe6SIWEJ4a4Mb1nsg6zsdZNCq8r5fIisj77+E4KKAi8yhucJz0seUIxtzLIY
fGOxJjquEGvGRVFto0tRNC1ANbQHQ0iNUmodk6U4kjXVRIxyEHueQKo3kQpH/+gL
cbHTJ06sH+K87jmHOJuGQ/VgtkuU1zenLhc0YXeH4+plB59Rq+dsLUkOhflBlU8M
0B+/zCoDrY7dkb0efte5sQej53KpiDVDtZuJeRPTDZzIwYLqrnB3CysVnuxSKDh2
Zrh7TrYuX0gAZABpBKep3wV6+wSDWEIkY6Cu6lIh0yzMkpKYhHFtbX6YdMBek0+C
B7ISwU2LKXXim0aYyYpDZ3e9OIbRM3s/xXT99M+dyvDWB4dyafFxlqLP5YCFBtNt
tiKOozt0oyjboHJ0FydVfdPaQXAXPInaFM/ozG2uG5WX9+QHCIQ69ka1aRpTaMGT
ZCHWoArAfhr+nXNyCbU2/0X+z+Pn5Riq1I/1dkRANDrlxMTMIjPxbYFY9y/cVZ4e
2C4CiFF4EYy+0Jts+DD3tAIpAMQL5snuaTKe0qrK0v7SnzOJKTwM4SsSgzv7IjSM
+oFL5TjQ/eevQBYKNvZaEmkeUT2OQUksWAhOQIw+Rd4UX238LLm1jjDiu81wWsAt
4/bZGYyRcub+OAqmSbTdOkB9ndlyW+oIwHaiR+VewFFD3MZ5/7fULjFN2s4xyw3n
L4ZVhL5MPznIuOFAYhVFLkCMQkbg2xY2Lm4lidHI/aCiPCmDB8dSNj88HPWJiPCg
414R/PXHJ2jt/XvDpKxZUzsREvXw+n/n1isw1wssaO9k6fS1H0jgZ7RPuAMazN6y
OeKmhB/QPWpnHavdtoop98VjzISPL7hFpr6uTpwoCXXgsNpFjBtlTde+SdWT7dY+
CoshMLRNfyyXu5eerAt/Fu8QoZl90Da7FMIG/rmvJ8eAgiciKb2RWIQcb/7UPFGR
NJ2l4jJDhxQRa3v8i10/GYyOJ/079BUMOykJcgRW9a2pn9ogS+22Mu1bFZHJf2wo
3ZN3CVoJA9b3fX4iBZgm41DpeTkvZxNJMoJ1YegQ9l99RjO4qMFhJvWS2sYZAsLC
VSYrQKN6klgOvRjgzacLHpsm8cF8tUf6E4ey0HJBb/C6rjCYaGxi0selpAVbGfof
heQraM3BqTJ5i3iFzl2q/Jqjb8j0wIkHTsWTvMED7S2Wb8zeU00NdpYWKmGrKunZ
KfzXQgG80SKi52kRAyPWreEOkHI1x6rAo5NrtEjnmOegVhDWLteOCQS88itaNqkB
39Ym6cRBZd7uycq6N3CprdJm6u/CASNlJJKhOOkcJIQm8PD/q2kwAf+hz+qqi0HW
+n86WaTzV4cq2KFr11VnsGPMK8vLLjtjPvRfTEIUWTROQgp+RST21U2RE0P9iqBP
EuL5V+AlknMh70IYUCvDpaYpyERx7sBdHtMqTZJc27cDcDugGKh+CyhE1CJrdnzj
4Jzffm0wBnh5ugqc2hWNEhpB2M5UVsEYFmv/mEN+zSQ0wiCRrwGeY1zW21waJNeT
3raUQdvaZ0kPpqVU+CpdDvQ3+pJTd29VRlyGRhNWUxn50EsnPY0sPDnrIJKRKixT
f6D+rroUfgvRQIbwMWheZLvwgXXA/cZuQw5RiUHBVUE8sChwSJqUnQlUfrdMUf3K
nTLFl1M0pcfdXX/M83mGMZc/TWNIMTZESZ6mE0HPdU/eGUpK0Pjee4IE2LnBW2aE
81Cn+qT7+Q2lRbuUOPPOMC81Y0ljX+9bMlFfQQPYLCq7jkcvAMORdrpLBPylqOhf
FstWnxgXWPwLg5bLgym6DbpWCtW+RrkTNKtpPo4RDqSEjNa2oweuxv5yeFZZ2nO2
jJ23KR0S+UX9VcFa+UG1SP26Cpx05F8B+pXm34KrFEcmvRjFJ6dmEprwYPrybfJ9
kspG8dYdEIRiSodctTyn3x8tvQOZ/J1zTli0PHMTB0a68VFtSqK6aZGhMZ2sr6bx
B+6U4uyAyp2veCTU3xl30Je78fxBT2/UeDVipRIh8q8NMfovNBS6vRajugc9yD6D
pmHpanHjKeBkfBzj3i01Foala5yN1SKVNem8IhVeQbrDmbOXqANjH28yVSfr1KBQ
etVWwXkeA9aB4f6bTklfdxqivL2zujE963PiSPigcDTK3sTylKFfgT2cmPfsemMm
vyeBJQRFFljUVi30DNC0kCEzbsFaSlLsW8UBJFenbar/GGNmQugVj72JKJ2wqwnx
lqqKzqbhk2IZ5HITknnQsPnAugEx50eWNwxS/r1Ee/3xlXW9jlJ5RfdNOfN9zE/g
d+MAnjZ5v6lolLCpCPYuJCAglM6DhlUSuyxF2fjnmJE+fxbJsPkEzXwnl3jfbtqE
W2a33lgxiZiUfwkuaT6/dM79HGd6dT0BHCBSZUoyxIcTqGZSujuJfhggxgmJGVwL
4anP2Jd81xIq2QO3IT+DBTETXvs8nbyo3bPwhkAPSq00cr/biXYtFvFKvivbDJx2
WKanQKbTxaFzkbecFywz0FDMpE0G6bLcCfhHjyTayTnoyb1IdaGzWNn2A4l0cs8+
rGDNdIxVxus6hkCRUBM1bB17XSkohcJifCi7qIre770gv9rkd5AMmJ6Le+guOafL
UkqHPWcWzG1PuWIYqrLsPCMvlQCA7rKQsAbkV9rIKqXFf+yDbxb8PlHMyy+C3fiL
42EbMKmZ2YJPKr7KsraNyR6qHXQk/X645zcPIMqnBCClK7N2qt7YvCzDKovo8PD/
XHDNy+umome76Y3VrIUNvQH8S+1y0EJrj9s0aS3f7/GqUP/wsZAteWsSKdpaUW9u
htKKLf5t7ElpKwyCiU0SSLYWr495wt8Hb83Uhckqevfmf0bCBnpLYqC9iZgekvRV
LKEdQgGLp+IKlU7ydrkH/L3OdPiuTngy7AgO6qDdi0tjsee0i8xD7nFl+6zunmI7
bbfp6JYmFXvUizpBMLfaTNVzsxYaiHqMhqP/YfTdDJchvWUMqWPd0czdAzqy4KGu
531yms0kuoS+4rZGhMWbT/53TnrwA/NiOCLx2VALqJVA6d5amQurrDxUl5Q2gx3N
1UTliZQHX4sGymIlnEXQJ/yQK/dkp4Tne+0UhYwQ2biZQQmZuC3eiPmUQYG9zoP4
x182EdDJbjFmz4GFavVsYPK5kIdr0AyaKAPgc5B85VgVGtdt/Lbw3BUuot9qgPIS
MH1JBo3PoNQtDM48X6Y22CSjfzEhOaKvKKkveh04DLTVExXcfS5Rv31Dn1JqJK4k
hHsaz/lVZBQwUgfiLMoU4t92rFGTUGn6a7OAiZlJWHGjk7QFlWkmBUx+KJ9THG5w
H8VhnLqbAK+p9hCo/5xrZXu7epdGLDFBjBJSCXnILtA8MlLrpAOSb+J0oBeTsv2k
aM7J+jyXtayo9uSK0+VX1JldEfGyfz78tK45ABgkWjbFKrbK1Qx4Jf8qrthO+BJu
prL8ypjJ/NRs6kSZ/tqhab1U3VtWEeVGgvjFenSyDs3bKZP856+gCXdOvyx5BIAf
9fAUJFBn1aY6BCMDqJJ3yZWs7/z78aDjP1wxqNE9QWRddjdqt4bwbIqAE+um+iSw
4qIsb+pHqM/EC2ia660/nr/TebyMT97IkEeIgmyCJhHumhibLLLvigZETQfqZTOb
dPb+dIO8IxthFQiv4l6z3Q3JqIMS9Jsa55IUTcuL1eC8aygREu4V28gUg9IZbxbD
TaL2mXaKk15OEu5BrFUC1wOY0QKLK1+fVHblOhZYWlHlHvclyhE5Awa7ROXUn2fN
ZSYlnRwkRrxcP3zM57ZwXK3e8VojxoXcRQpLv5EJYIl/6Gr8QaMqv9xm0MXYcXv/
cIkX+YyW0E3scNiioBdf4sBDMJZea3llAy/lY3vNGuXfw8P/eGW9Pw8/uMoYZtex
FYlsUrBjra8nPXhl9qLba35aNdPvNwNcpGZivUfs4hEn5gPXOuSv+DN7UtwN26p6
/JsRp+gPYZWbwcKzXoZNhsEXjBRE7LUMmCqSTdpUigdoMRsQOqxqEKoTukd6UA+0
9pLvS4z3BNmyZ93cGsnUIF6EHYTaGXlPGXiyOjWbIKtxDRNNpNVfG2mIDrY6I+rm
TyH+ITEBdJmVFm/lVPMCbxk6N9D0mJc1NtK4xvaT0FhBjSC2htQlG+Eh3sOf3yIB
EVD7mAHt/O+W1YGMkX+hKitbAWKHD7wxDDO69FHM5t7mTtx1+i3opKXPFPpIXBkm
CwIbHJy3l+5NVbOH+HzmrIHDiTHxNVtiyjLN+ac/MOPDpShqWY+JTwbjSu0ooaV4
Usl9uQhE2buHJPzFGO73QV5RkigaSKLaS1E4r4O7L1lyzJt6unYukFfE99OnUR/m
HFsJqwJ5Dc3GIBhRgDYD+Lt0Cd5KQL/8jRmQHudsEDEz85igj9ACZFDlcuVV48ax
gn1MoJihrEHki5K+HjMrTGSggyutniKPGYH7DK9qNJgGi0s+Me+xOTW038twKq7q
9HFXZ+dKXXc4wIjYgKQKXzA/mJZ5a4VEVWKyG9e2yswiN4L3FZQ5LwvD7o0ZCdUc
RmvERlLot4PgyRVtrLjEQchIj7oYqhOEXd+54c1Me8NtWaoWJB75gvPLhR+3wAlr
FdsWp2eUH9T5lobsKCSFzjq/Y5P9jMiWd6+zhJPTMsZpEx7EjCXHP0XpxaSSfUaB
uOM/JP8LmMVeZt2MZQSOnC3OZZW9ZpmIck3w98ucEbR5zXiixpKXuiOrHQY/bkVr
/oG93fPUDHo1P//zE5ifsgr/6FIF51eTB5W6vaFgGXvl54UtMTRWNQZU9xrmJzIk
eTl87AsHdstmnKq7hQmMsMBapEvA+9nJCLJRfuclZ0s/DnFZwtUOqWKSpYAMLag8
DgNmMANrLeR1NWmzet3GYDzxBmcE0rwNPu6S15UeDezm0lJJ0kYXCpP12UVmd3ar
HMS/M9HM6v8IvMft1GMQsOdUMfXXhn3OnTuL3zUglnfpH9zCWfhmcTW0TBmDKqmc
MV7/53cnTZLVjI1g5bLolggfUH2lqce0m29YN9AzXCzknHV+TixMAwosLbPeWMT8
qcvnwpA/Xxd2ABOGwX7riKLH8lSBlnbvYYE/LOrWOHX9KZ81A/8mYIqSJEsYx5Fo
prtHaO6/LUdeESJDh4dS3AywQ0ms17HMen8okhi/fhX04RwHs6PWE/dYnz7ZjR/X
IcKgd8s+oycdOYPdRuXhpHQLmAvzfbyWM9lH1C+8bYnP0C9oC7Xq7WbijZSr3+jS
LZQRern33YSc1FDk7QzvqD4/7siDGfc9ueCxk4/2CbHWwSQK+diX07W4eqp5LCxC
pl76iIvD5e87WfuFf4UErJ5PCAAou713WpVdoiilegOm3fUMdRO4MVqGrUJu0D3g
nl/VUQrZAWVvUN3AFAEMqtOgfP8pWE1D/aV/hDtsN/a7a/Zo4tMk+wOOm0HC7azE
//fz25pbxFTxHa/Ro4jkkbXF7G/2aFWuVmemnie9Gur6QCjXTgmPIeTMzUrzDWmv
NzO8sF96CLNBdarLS0/AhFO/AtfmUdEzsJ+PU0dCjuKqbE8R7LYTFq6xXD8Z7d+Z
ceuO4QBC4e0U0cOELaMZuA8FwBvPYzQ+BHS4p14vjEU+wPuzUVva9liZyhbnx0L5
8GHxZ/OAOPlsW0ZXc4jMcMgeBYUGoT4Q8S5i1pvHR1PdT7KiJeyKN+pMen/ytZyE
9m9JosUpP8hwRBtXDr97bEVc44y/743TqlUDvgGYhYY=
`protect END_PROTECTED
