`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jsXW/Z9KM+0IhbVtqE2mJJDWQRYw0XL0ky0zfQvhQSzoOj1XlulsC4oSsHZiYxgQ
Ty7nqBBM8j2ve2CpkzOY28Ic28PuBuNj2vlUUJDGvz0t7PTZP+BcOb6lnQaCX8HN
Lmb2P/fSajvPjVKXImflxux+E/SQYcMMNh68tFKBYLJEiy7SO76ihnE2woaNXFfD
7OfqGHMpPODcguq7/0r+3zoOJDzzUzuxti/Qpjmh/WIZ/gKVl8XB5ZKpw8xnfMXu
pv8L4N/6IsLot0qAy3JHWPkzCInUuRkd/O6tIpiZ0NLUn9E1pRhqjIaPQ54sgeUm
KYbRZsl50wt57X6Tqt7G8mG194AJ6vhMWGLZZf1IkwJUHLjwgR0p1L164EtPdn+g
Fpfk1nIPT6pNfyvVth45K8eh9U74studkAVmgGud2Kt4dtiYvFLD57NMA4nwNxLB
23ya9fDPmov9XUB3I11WIfZb/A1VGmJGAkYUJ30fF+ww4acbZl+E5Rw1IBQ9wi1p
7IanPCIYItH6vDPE2vtY5OUIEMWzNKMvTAIJs0ixiMRd4l70YT2Y7LYn/Ct0s6HT
0MT74gvJCT3AO6UfieLYLXETx1IOjrwLdhI88qPWJoawO8nK+L04cnviCGuMIE8U
uRr+kvVUC4y2Q7wtG6bOp/oWPSXjqspj2yTTKYcrtaBzjK0TNuq6Ia0YQ9VG1icz
+E9my7FYFaGBXH1sZJHqfOH1Q/40Fd7dpy1rFcRFFwJvzwEt2XP9LUcjHoB0UVDm
BT33qAH7YPatWfmJed0GsLV5/aqltI1rJxOMmM8Z92gpBwPOqC7w+KgJhNjLAo51
bTpAj0+XzOKsyTv8KuJe1BDojO9L/oUnMQUUu0XmRNs8AoIwKrzAoGLJKVYbHBC9
OXfiQFjcd2ysW8Pb6eQxBYVUc8TSid2NEzysBlzOu1qXbzps32aNC1PZAcFi1Gmb
sYf2vOaK5a6nez5u/AAtmlEG6xHf3efLhcV8+1gn9/jMnWlJmhe8GwA1gQwHjum3
TlAgWoXygs4k1jf5XRx9rIkeBtnjeXtHqARS5UrPoisrxiNWoh8fhtkU1IL7ioXZ
ww7irLMeR8B2ksW8wBQbQ9PM7APj7yVr7pSuGUd903Daq2RRUY7LbCoxmyaH8epw
6a2w0F8z6jov20H7VS1y6wcdBWJgtwyAHPdILFNgc0TZT54hQDhccXB8chPU6eNb
hHGL3KxId7wI5voD3M8Z6/hB9EbnqflrYqDlJYbwxgjmdy4BotAEgqFKijmnZnl7
9FfuAW3lEYVVXHFPptCp3Jjm5qr4wMA6y17tJh24Uz6U1RZl6oAMaAdZvVis025y
QIii4J3bR87GH7o21qPdhN3bJEBEBSvUnOID0f3oi0KU2EP9V2gmM0I8VbYgFEqW
TrFfhetdcGi0YpPCgPLhqkjkI4jXgkUal6czeJH+O9jMGf2YBRzxmLKpQuSpce7n
4w6TrB4ZwU3znUp+nKhBlKscyGIVAw7sq2/eDdbjf8cRpYY9JKkjbZTvN7gYJWge
WO6zzbOZAm1hgGas9CuhAbbr5b/BiH6kEznfPpEwU3RKccta5Lpb7O4wceTpPo86
JhgnsJUjkrUEEPn5MDAqMchr0vW+ZkuaJW0Agoo85HE7OYarzF4XjvLvN17fMInI
m5cwXwcgK1nQGnhJasbOQF7K8JNsZ0nAGbbfvUB97tQSE9BS6lsxG08i4N82jAKK
arvSAqza+qutvB4BAwbpi3FaH9SY5/c0GW7CINmcASEUqQuDb1oEHRJTgcQsfLR6
1xz7UQengDEFIJejKFJEyQD+qlKrUzJ4Qw/CvPl0Qx0br06hMeBZXvcpOYXhdgNc
NxMiqKOw1Uz5o01qJH78ejhbEGFvaIrenuVxKfCWNXmnQ/OCQwZnFeZXOxpj1tTR
a3on3jTBJd/RebkKw4OitMeuK15kO4nwv55phOhv/F9zVIsaLRLl1/NxbkHBWhYK
luS3yL0NlyYlZUHECZP5608ItpwWAVkUBYriE8VVKGKoy0oeq8AdtFPPjgUmDnPg
Ftvebxm/e+NIIBL2ZvMrr5kiPs10mr3g+msauegX+hy7/aLxj/kJc/KjD3c+5Ujz
BnMF94cCXRA0wFxIJ1B7VemFxaHd0TzQpkIUFbfb9Z8Uw1RzaF1xRwd8Y4VRCs02
HCNgSiztZpdqV88s3F8NcL9YUPiTqKCxlKP6whcHMtnNu2gRUOLpkckWTQcpHiNJ
YpYjoeK+M5v1pheAeFwLb+adwO4mt13Fuja7RnieS0w1i9Nowem0fUkDYG9RkAHf
QDnQ/HXgTpAVm3jEAdJFDAqyq9v0K3zogrbj/QiyYs9cwIlAtG0OnCqULqwh/C7z
HgVw0+71UalKY4EVP6S4jc8kA97iz6bPIsYqlc8jedwRbFvRpekcKEo55xb4IVz8
7tH5wLGq5gC6wC+fQRHt6jR21yI4S6svLzWrAlOWVgYQBdUkWA46hUW7zNpRq2q7
JxP87m0Fg5fiLor1yihLfZSmzRhwRJHsG9dTeY76y3zY73pbWY/gdazD1rV8nOlb
AlEnbf99qcP1t02Qi5Yqm6AfhtTUEmbUZoXwonHXxreli1xmXmiNDJ9ZyUcw+5AZ
vy+UbEUJdG2pGLdGIbN+Lw3LF9+uqJnJ/YPyCra1raC+YQWL1nHN/vK6Kh+OhtCY
6pWwbDzFtj+O0voPpd5xnjhsgl8Ypw9UL6AUMwQBw/y2dOFwshrYjgNcu3qPXqTi
ovtZzbY98MYcKMH89aoRaemvvPWoekEpt6yAHykh6sVPZ8F2uDIVxu3ZlpjPSacW
J46AgGj0AE1Sp0PKxOty3V4B+JJWlPAl1HHs/AMz0AaIi4hsWNxlWxELy21Ktzm4
K4KVF8A+jbXaBKLYUDG8BGbKNhppSAjhbEjaqegMFfzkLhrtDB2SheZLRqiTz6Jc
lb7ZvKF44MD5AFY2PXt9ckCcmyzMfw93+HEicM+plP7wjjgfCocgN3b2NXQ+wI/q
vLC/OKE01/PLsz0JLhwJxaWtSXj4ihgKFWy231B6iqazIw+VqQfvhrBvwXcHJQf1
Lkp9/ECYLM1HjN+VkhCdmaRpdFL+P7VIoPZPMyU4FuPY6NInb2Y4x+OFI6oj6QE8
ep+Vs7uCB17+l5Y9GJY4PWQPbeWQkq8CNdOiHdtOmXwuvSJhXO9dCOnbdVkVWogk
4uyAzOy21wUJXnMqhrvavxN5JS4F1lEXvfs2rVak4aEGvsq35ymv7mdTJ3ReHu+0
YMeN0A+9VO/u/+Uxz6MfBSsDDNzTLSu7afWJqreTzeUfcX7V5tmmgDMT7e2am3a7
yZ7e8NNfyywpVL3WqUUeOiIq3c78pkVUuiS//MZSgZ2b5Xj562/CfUt57KrF4BUY
ehy56AFaEuw2c9ntgTf0J5s1IgFstJO3Wt/VWGhI5j3FrN/OMpXYCpFdEjAmXGnV
aRnzw+z3ny1S+R2TXL8foEHmTMTQKiLPRj0WPZy3GZgIq9YA+iVFFMtQqo/W782p
ql8YiKbSu7eI8ORm7IwmiHNLWhXL9wtK47rLEG9jd7TBCw2DZjkfxtT+Gk9IYxbo
+78Xz8xnA1QBZ2Qtdw9DcegQdZr3TGy+0kR9h8OnmE3EwpyVWeh78QuQi6cwMkTX
eDeUEDZL4tMttjGHVcbjqkiwpGZ45TdSA+Binl6Lq2HHsy8jElsfJe4U28zfEh+s
0cTT0ci+dzvIl//w/2O5SQ==
`protect END_PROTECTED
