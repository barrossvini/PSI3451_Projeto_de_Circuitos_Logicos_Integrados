`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CeiXJUTXryOvqhEPPZ1ZaLNdRymig8BL54g2oE6mQTWvSDAYvdyHe1136suS6zkS
4hDl44QrWZoRht1wwg7AycxjNjw4gTmdFyxPmV0vPRFEJAASCtmgWBTKghKcG1kn
7GEn2PUMXhIi9j3GvIbt3s0b8ZqsbwjcGR/ILdddVe0hZlbeTDnuBsyLNHct4nvJ
d+whw9wT3W0qVQLqfkU5616OOt5NSwjnhEznLTQfn2dCBlicTRmg9u5mZso9TID1
Z/y/KaGI3VpwTIUIjGe8h6IAOQlro6ubCtGy/ACaQhGeRZpR0cB2QcpT5Ptkwj+W
iDp300T4i4v1pUCEYtNY49xnhKPRYMlU2v4cUDMvVsS8NghPfGIkJTPeyQmMrN0i
CazpDZ0bROMJ9zGwQ4i4qwc66KJrMCmCilps563GrQI=
`protect END_PROTECTED
