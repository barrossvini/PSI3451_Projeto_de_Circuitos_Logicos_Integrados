`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qbO5Ab0nJYfIuH3+ULIT2b7MiirhyTuH8zQ5uo4PWZwzw5gFjcRA7kDlsLV/lVmP
gSioLZHXtHivQHvDV52LoM6KWg3szY6m9zL0msq1Kmr+8jAKFPaJraalSvXqoVmg
kkG8bD8+Y7C1R3jfu/tamPaTsgui7jTQ569yt59ImdOlyH+/Y0XJv9we1Y73GFiN
bEJOesdEki428himKj3Agnd9ksdA2J6gz6E2sCviPqUEhgs7Gl1wdp8GWVjA/Vtq
Q979t05OMPjqa4LnrYutoYmnLc8JII6cwnnjt60vtRnLBJXU2c5JTtlLCcVPZAmg
Pr6wpTz8vDPpOdfe7ccQ4x2Zb2eDpS9ZSHnRqFXHITVzclP7Ys7JTclwTDg2HRiT
U6a73PmSbyBcRwG5QI5ICKFa6qppmrfu7cjjgGzm1QqzQvIREJ/8nh9Rv/dH4Xm+
40OqPDd32MbnTkkpdTslhDJdJaSE+SE/Vi4vZ8BqyME+x8zzpqAJri0UivNWCJKA
YvFM3Smdk74LG9fv1Iu+9eUqIz/MIMMoEejWp5JSKA7+uHz/aCkkP/6pDXkt5wF1
kwLeJt8WcKdLwmtGOPIyDcrtcURBo3kQ6JVeYPOZSlfG9H+mj9+blkh1GuQ+KRCD
Sbv89e1UgwQMYBbdXHSeeJA3BavWKS7NqNxuJ67lT8fCZtZ9esGqGL0KV9YSi0vc
B7YYWEOZYkl/5BMfRIUcBcvog7yEUQrnpce2Rzw/C4FeI7TsZmrhzLXNhefn2v/N
6XtXTpzIlwrVCjyGzGckWVw5R1tOSg80Wf1nOvsTB05TZADxnFw59YyR9HE8F8sT
mFrTAm/msphkG3xrQtZEXwIP1CqiX1Hg+Qj6ysKYAjMaFFzmX1pNbhb6mcRHlgIP
QyhoWWUOF7kyOUplbnX/Q7Y1LhRp4w+5SuKcr6aRlvMiHQo0iViL/KVGe7v28ZU0
b2YrAiC4IlG81Y7+hm/cisrPIbwuDNiDJ9C4csRsC3kWKCEaYHCFYikufBE6RiTL
K2NFmlYWTcCpy03lNySxg7G7QdUeGI8t4/uRQtC5MAuupCZLDf0+z7m1QsTRQl9w
TmL14INmm421PDoJ1vw2DelcXw9rjFBnz1W93FANzAqlmVXDOEBQ1PnXIJ0vdDTP
qtQAw6vhkOQbKnnXj0/Pi+MPcmLGw7gLf+8MelxBenpfSD0bjzjKEMs9SgfDmT7F
4sx45lEs1c4LlxAV7rM4nn5HBIb/DYW1rYawoiRoCfItx1412XOm91vbJrCidfZs
kuH45h2LHQEzROfLta1vmPgCxMipeORJsAS9kSYkWWm15o8KNRfPJ1G2xw1/J9SE
9CKrfKbhpwmBotr/WvwJlj9nPty9ZR3Q8UaPhXEVxp+BZLAbxw7xfBEkL4b3VM0i
kEiIiq5ZVaGsT/6wXCTiyTyfmoi52Ou9QEAWqKjSxc0fP3MvTE3DvNpqbwSI/apZ
lB4V3zW1FUvD8qMCTS9GIzBJIP/YB6OkD0vkAWsP4a56x3eEI9OlG9Cd/PS4eLeM
z6jxDu4LSTXnUX5r/Z3aTPTReotLze4NigKMcXqglJxZSkl6Y17/jMtOu9gaej8K
FnhRtpEdtchJld5UuCNXCPMIpqNnFPZZkIgm9I/FbZfDEW9PpOWV3Pkxb0tuWyAN
E2sZSlkg1Zv7LgX5dwLA+9OuwkNyXNob5gLzTT5b85T5oq/Y+1Rbko+4wxWYVYmz
dcOSfL/ljqCLFFjb1u5ah1rL3+EvpJxAdQKdpbkgOQd0pfgzybZFptPgo9qfWEJD
qgFg1R1voTsl22x5U4S0UwZCFrZz8v/deiBxkx3ZXXxhUt5JC1oLosqNlATuvH/q
2pvmP6W2lS1IMfjGfGFC8bfSG0cwTkP/8Odp3q7GY2UFvxexohUIpgkp0R8m9n50
AiAcl/kHeGdzMBHhaauDpY3vliiBcJhb+eClIx9nK3at7kAGfZfqGKIjL4l2A/FQ
7W4VsrdyrVyDdkD+WknMYteGC7k8nxjIRSv8yzCr2Q3RsWMoQHWWdh55UdHHKh2z
YENWVvkArnO94z1WxYBiCCsNtCixHAak/ok0BygfhOz8SLHpfhWHTYh2QMzHrNyh
0KECdnGyoHWPPoIBULLmM0fcMe9kSswnj9wW8sshzL/ZoBbQ3ERyQWn3WafmfJi5
GJyDd9PTz+il/l5RBAXqqcG0F1L15Ve96fiePnrsNKPF/dlhjLBYPInGtIoGnwQ2
5870xJ75CgvHF0iFFmHEjufaieHzOq3csvmKYdAf3AAK3t4qQuk3FChcnu+PrqLA
RF5cmAveQg6U4t09jx+4R4SWF3Ypb40WGFS5OSmkeigCkCrx/IsF2xstOPfUOYXO
s8nuI9fc+ngLOBkzScCdbem3YsBoNuTc5Ivy+TYjkhM+7qgHv4HO2x0w5onAQOqP
j1gkLJAa3AmxbTHf+UMZYb0S1WsAJ1j/JsrKv/PIvcLZOG/C68ejcmTJ9aEX8IdU
wayJ1j/bGFudQn1d89ILSIEYkiRDDeL6yx1e/p7ftM0jjrCVYBwrPxZAjVxA4Up+
c0m1cXBQVvmv0XPiaOvUqvmlJbLlVe5UygwV4/v/C2WaenWMT1K0vAuXKEMG6+Fg
oEv86CgYLiyn77FChj9+6fp+ZegOKEvPS6hNc+I2ZLwSlav4DLaujFRYdDOMnQZN
47zxcBnfGmJ1kwisat1ebrPCFiQA9cvXxuaRfvh1xHj8kTOz5e1T4djYOtEXFAo1
O71QsF/CV53jPpPnVexYk1AUmUDhqBkg7blFRGeHfqEU0Fi/Q3QNcoQv97LqbSKj
BWSm/VBDTLV7CHm/kwGdiyM0h0XRb2NdZqQvO7Zi8z+H1CnUwEYj/1THPMe3XgwZ
rqkksetTav+9qau+07ThTHd0K64SIS36EWIVhir+be3U04tdNP9x+KZLAmGlmBdD
iSdg+H+0eemxwWPqsUYNQ0K6LgqNrFjYBDsICWrwL6fInUJvElcDWVsOm34Mbiiw
hClOk7tl+m8Q2/HanTdOLFD57IfoNhxJN2pleUU4NGqYH0jDoEygZ3b/vhsZXU8N
rLqJYFgxx3cH5Z8BOcAvwA+tJ8udupd/1SoSUmxcD+No+yAM4Z/TD5SrgJ0e7NYQ
YxLkkEXfdlWVOvDNKUMBO85w4fd5yTok0XtYWwf+wkQRlEzSC7d8QTW1ohHw5fc5
roIXdehPgLThTJz7lGltQD24pb1qvExrNltB/wVyJjTAf7TJ8uT6bC61xHYt7TvA
ya+O3EyRNr/sRe/cLRxBkoLf0bCrX4hs8WFq/RD7dxZBV6A3BDGV3bsDX4TJsBPu
q+kf9NjghgJ4t6/utZoKttF71H+hUGss7NXplJNeedzXN5lmyiVXVKDPHMHqUyXo
tZhnDQonuges2VlbMViLdpUG6B+61IF1U7Khjh7H58a5o9Jj9gCYpPqDREoGvhHe
YjHbu92BJKRSVfGfIw2S8jLRFBqhHr7OjOMcCpyOatUDS8sE+Hv5Cb9T8LbnZqWT
p8seVhN9pp+Gsa2UoiCx0NkrlqbS/1M3uzj+PpNwcevmCMFEN7aUrFJAys85lbdT
2Aa7eFlb2qGjia71mg1Bw6HveItp7txHRNCzGynUdK7PnlpDP/fp5YIQiu1hT7+1
sOZPV7R//7xJVJ1494cX4TIzukqyyGoCmckSA8xMfa28XcEqMPyoqEAbH+jxrfnu
F4rpa3ZBsw1PwD4B8FGvyQZiHb4UzyeGYJMDw0kmoddYR8aHj08c1I+sY/9s1vP3
AWwXX086eUv26i3bLdzSDUu1WndrXbzZGkQ61KhCWvrXMBg5f05zC/VCAz+XMDIw
1XHkqqGQNcSfwv6BeDm66LThYRLjn5PLy7O0NiCnA0daIohS5Q7+2KQFfc1+iOz3
qooiTLQMpb2ycA8kj4X8HV8XGf1m0JS7igacnweqdeMfKnU2zFNqjDTSz3mcTb/y
vLawmGlBAX4tuiMiuuKkSteo9G8IdQ7m0I8HKojIy9nWe72Fng2bbyuQYVz1Jlej
hg7oXM2uZuQdFXwog+kdEmxuSOEIlgQn2A7uEZFqjAikpIhG1PTyum24uEwjnfAi
36iZhRk/rW1yGuXsvr2TbgdEPkiiXzzAr6xM6o3qCHK45V3BGhQTXSxcARu0zkcp
kuI7jhg5ODny5QqJZctIbFFPGDPMQ0UlNYfKccL6BH0Spk2sIonQM26FSn7PqVwi
7MjrCBzfPfyJeL42DgLyOF0TktfU3c+VAguXj1eUGGBaGBMDWIx/Qo/zRYqgK266
LFpGGH4eMCKqAhNtVwhy9ecS/Zac2wIHafyw8r3MnjZ+gPrg5W0yRzkSXzBY9e1Y
jZ3Zr7NtQRyIXVLaKMHQM8PmbTYnIFdkyN1FECkipRVCTFREq+onE7crM/2TMHo4
gFoNKTO7hKDbw7F/yfWuplvmoG5zABs4aUPzHFJ+axyZCirDPQuY8HAap77hfNrp
4wlgX9kQCai13CtdPs/rfvjJmy/yHM/I6U17GXlDupqN/11A79ODqxi1dSWv3Bfp
xA86oVJ54gA1PRbsuCrycDW94lvnLrcjQlqcPKfFzNbjXRiyRBylEQGi1O0gaksj
jTHSCLSdG+ZxVHQWnBcUkoqZlfQH49BNzyzI9pdcH8ydldJ9jPFbFZnuTgSUjMwL
9IxNj270QbroQD/9QZzfbWzBrH3fc70X2oJCUhs+opxU+v1+gRErgTwGzJJK7Dma
Po6lAaWv7n5grnhS3Be+1wsV1iNmvGawQKttn6rZET+tlNFSxXEYsc3swkVnKvdY
L7e12rLdUh5Sl4bCCnJuVKlAd08/QyED7LKL7MWMaeGVywU7fyfdZBvwheLkWWlo
JMIMZ1Ykf4IFEpHjR3nkBmQCkMxr6mwzn1GgOsBdndtp2491nc3C5m//7NYHTxBe
Q30lVtrnPI4rI5kdHhJdRRwJ8jzRygTC+mcMU03C7UGFmnUPPd/H0w035l1p+oop
wXIqnbItgRuHmO0xHHe5KafT0+JpuQsr4Vx5tW7S3JIVQGdUpZmo9xQUQAUDsWK6
BpagUw1k3LcrjduLNckzR1LjHITyKS7pxQLQ6QbMDcu1pxV6mEAY0PU4lhuBaSmq
0TBkq7b23uXCx5QG+wMx8QEfCGV9DASLwzIYhkWvvQY0EZf6RGBAiTVqZ25UEYdC
loKFdq3BvmqcnztRJpzCxKOm6XzdUKj9D3lAEWgayoJSM0CkUzBERWS6sdpT5av8
INNNcpueE6wLbNz/F81s/ZV/5eCnNXulzMtRfwbfNYOTL+Utiq5Ld2G0Hy01gnfW
xD+V2epJLkYC13LcsvXQaQGgDfXnX6VWk4eCvamQDzZr/DcldNWw1JakSBwtYx3o
jOVEt34ibk1QGhhLowLzV6G6bYsZNkTb6onNmkgYWUOU7DPK+ByEbDE3hdVkE2EP
WawrspmzEDVpHnjQr6vgG/4rwzzrdzVdz/+ohFUYsykuIP588B+hYwzXef/ZqBDl
+TMCxS6ZP2Auw9XUNNNGenLYpDslMnDrmlOSmS5TWQ0NVwy2JTqPBCXAbenYTWUg
iwZH1bPx/n/4gZbmJDjhOoUpe0nWA5NsIqRUmQB0ARDMH8QDkjbewDTv6ShOLWZj
jrAi7i0hnSGnXm/uewZRJSVp7xme7jDM1iEeI4XA9GrqV3GDjKHM1yIKDXQ1E57n
ESvpTXPo4MpUniecK2GaR6nBm35kn2HYsf3W7wfDoLz6uwW4yaSpMEtD7FAj57QW
rCgB3Asal0i69f44jDt+eAcHqJm4j828n5cSqk9N8FsE8E6aEntCfrm/NFsbZQOZ
a8Jgs86aQDpfNs8w5p0ySwoKiTqkYU2sQygrZy5Ss3s=
`protect END_PROTECTED
