`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PrPOHv17qfpdTZyaEXZfmmMOb9nio1dnQFJJlpK4FwUTDMTYX+pngE+FDhmRcqiY
foTlo69qSTnjZ8aX/tV0NgsY4gYM51c6WD9f9gDKjKrQLPDm/Jq0eBYzO2SnEQC3
J0ZtYnhQkK/5bUoIbNmV6rij/L5/8TlAHhSVyx8qEGxJsukmCwgjlm509NqZa+fe
QV+A+gVUcmEtKBPNBSNuJ+1PhsG+UW40Hzk+Vtf98/3SdOXVX+E1QmFDOfbFGeTD
pnSu6jtrWjw5xX03WZy7zQcUqDnkfp1UI0FPXdGy03/d53I9MjU+Gbfb7GAHl8oo
UnpNj9D/YotxxvKBZ0ow+PBjvP8fRm+27gl8NY0b9hEQUzeLZCSZmLKOiqujrbNI
wV+0pwfRktD3NXC+UZgjoRv0+/JWU74gGt05VmnM9koci2I1KwMhDBCrvo9OzT5M
DDWIwpj68Zj6mXraos3iNjYJwVV/LBpWw/GlPjguDflsAPWjGNsYxMsX5K9kxDWr
SRZHMJYlFX/onteNnPS+L71L69YbAA+iA4ONtwkqel+siIgD7TBN663X8brxnU5P
`protect END_PROTECTED
