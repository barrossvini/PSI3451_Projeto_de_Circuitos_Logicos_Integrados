`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M4cJ5b4hTTUXQ7koqj101rLJ2jXOcUimEnyfr+rLOfTofz7ouaq21WVDB5g0ANuk
fwjKDk5S+1sAdDsMvbzLK/vGBBZyjulOSiR2kj7Q/+6sD7sK+FR1DHqde6R32OZN
kNrpo42z/EMCxhPsJIQlmWAmMJsZaLW+JLoXRnDz9TmIna4UFMy3hezskg9molsT
4517N5TFw2F14zIJI2Qfafh11YvH/60mAzPLgUGCdPlbv4zrUwLZwVWwfRVCPZEK
xKhFsGfCkW50EcHEEITEJQNYfdlXdtb9mbeGkNIwzrX1uNGA08qI4Jj+1zxOV+CO
7fLgXnOjmWDWkbozqbbrErsyWbJgzp6mpzItF6twstRidgdHSl7+z3yQpN5i52Oj
ypKe6Bmyb8nqUGviofLfmh1Ps1rlsy9xzlsXE/JNYsq+szX+U4LnVe5uIR8WyoKs
zwDh5HyP/Al5GC/QxQ8u1u93LpZaUPONr85Hj6LpB41jMkzqrXJSE8utZ7spwI5D
Etiz+98NPkJN7fiyudrZsCx6xLzzeE+Qm6q9aZQ49GCujE6lcY/Vd3GpCyKqNsI9
bQuRzjJpdo7lIGBAO0YbNPFi23M/ec+glL6LKdd8EvvX9mtMLOnUpb6Mubj5gJN8
tmK23Pv64lWeRpSvB6GO893jwI8WWPHqomkcGU1HEPw2CGzu+Q4ZioLUIRh3sYzC
umwzbu0RU0wt8cXhuINwRFmYTH5WDFw1P33R5n8m1oI5MO+T2zULIY5Rzc/QiwqI
HKA/HeY0G4v9GO8csOmylKsfptuiPaL0KfpaU5ZSQQjFrbC6G2SNRbWVcfR3csBR
Xm+Uy+kQiN1QnXGhzUcX6FlQbrpQIE/s4VuAxN1rqtM/VLZiMWjXfa7uVSyao1eP
TX395bdHVLk9gllpnw1FgopjAOPeFgEzj2aBlUvArX+6tB3J/lS5u93oiXrN0WEE
q8OlsCkrLboo7ePP/RwQam/QNR3EtZXG5cmnH94tz4aNI7rM8jw7u0xNAqn+MZqH
f25WoF5JC8Dv85tDFZExDFsqmOZI8YDWQkYzJkZnKGCxSW8s1vcDf7PkRPQPEByU
4mZ2UhddoFJIgEGpvk5okHOm4Ymqdx0SsHnD6V6w0vPzPZxZKbljIsUPPgb+NYjr
2n0C4kyUpOmppB5vnlGjSjQY2RkiyiQl8SlEsjQwCjs+V+dT0lzPAoIoznRdEI3M
y2XOlve6i8o6cbx0xqDNoPKNplktd6uuzGqDqZ/H/NRYlzIZq2hjp8itlNIt7BS3
q7rjq2QGcSRKi737N8OJuFKGJgL65T1bhTTVxcTd1hZZATYaHp0w/9XeBvVTRXay
0NV8Kyhn4LEZWwiGIjN9eyndYTWNrU13imzzldsmBoKW3JbzDb3T4ehizkQ5Sdfz
yazfoZw3Erc6pTaombmpbTgXl4UMPYMOHU7B8GmNmwI0DpLL6FT6A7ikA5A7Ytt3
wmGvZnFfk4WqGjU4mNYTnthHD79TmCz6KLEVA9Ljv2FUA3dDw8LFBZwcaYJGZwtX
oMmx3FPgEdS+X5B9MQQ0d3Yr6l4uKsBcckErdm/JZe4YayZU8IHxJLFDRDChPimS
ladces+9FRZfGCdBUHy4/yw47YGt+JQdGiUdwbsvQKNWh0cNV1+eCuZglsZB4EA2
pZSKuRGhgu52qL2cPnvIz+7igbiuGSD5CUpJo1Lph9uza1QwEB1qlfLCCFSmXC27
QwJ8o9EMvAN+M/Myc0lrFEx8BO+7bKjCfEMWweFe0zPrXu2n7Hu5K4qn/Shs9EXV
ucDL7PNfpD5KQBgCzp6zpaJAGL1l3eLsev9t/+yfAxMbpuP/25p6QXVOxA37jQrI
NHkuIKuyBkn4dyu4PFzR1N0xsiLPDYPfKOHLL/rfoqvJwBTdRJr8HwqfgQPpVsrA
iGA8pVz0k2Zf54edDsVz7EBKAgjtVcEF7Ij6g+YnQmeZfsVSViZx21Cl3bMIs20I
rmOWPGE17SNPvMtunG3bs/lKNYuTm7Az5LVkoBV2hekRCXUyGVj9rtHAM6cV4Sg2
9slqnqlaH5POxLiZP2U3pS//T9TGQfPUOwTFQxFq2Iv7nRKrdiczmANUlLWhCLJm
iI5foywd1SnLle7OI9T03oHAtpPBJBNFzfuTFYjd5JeNOwCtQczJqw3rFJ/5gCWP
SM09iqtbL3J0V8HICTn1haqfM3qWafauEorw4GtSeqw=
`protect END_PROTECTED
