`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
776E6hZbq9j1n17iUp/DQTubiXpuva8LN32oPu420ASFQBynB+IUf7D1VXB/dWZK
RxTgXl6yDgsVulkvRtyHNZdPxrQtSKnsCRRVn36H2WUxTnOwosmllad2tq0fk75E
cj/Yiroua8/8jXWDVWQONBKV8CuY0hE8Kf8vFCNiB1XjCBKgGIBLNbKHQtb8FJG5
VwqGWeQSdUJ+eGZQ/mi0/v6ufN0QJ4lwm174vw7YVR9N3BOiHK+SVvda65pAm4T9
5S5WfPxdmdu6QEG0TndPqEptm1cToPuMFP979/SCW3ASDvrqHuGtEqXkBZw9aWVD
hweaMCkQu8rYfl2DSQlzfjJ/r9tPJTUPylCGXo7vdFukGyFYzy5W533Xf6FLl4WW
vKSXlhSFgdm6MynjPsoyZYZGL5YCunhKkPyhgoHhxOEdxtFhpeT4YQK6+z8ukCZ0
9a3uGdYcD1ZaZBql+zE2nE5WPedTYsneEZXzKmGjb3jbRJCuM0scyNYjADJfagoK
a8AKmFhQn5LJ0/iBwvrB2w==
`protect END_PROTECTED
