`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vs3rSjK02vlq1/qrtHh2WR7Hto38EQ0tnCzsJoY8roij8Qjpbd4ckrlhDknSAuvs
QTsDHQdB6xnAoCGCahx6WmisYhRpl/eX/1nLm4YMbZRn6PWvpJDSF/hvNv99bvkf
6rbm5q/Sz/jJwGrPfwQax3xOtZtYqekOSe9dzLaWXEG+E8wrmcuTyJBn/Qt1Kk9G
d06ed8HWpCiJRXZYdk1IYfjdP5QTOmaJnIjuXy29pnabp01121AllbL3lRNa7ryy
yP+niIQqk6zsHtY6rCS1TdzPNwMlyN4L+u6bvkJjilZe3XfP/HHhUiVfr2emU5Tv
4ymQseovMxtefaOI8P6NAmqTNZe/f0axBCXmloBqbCQpD8EoTLcdHquxBsp0gou7
CgAb5c3gAy0Lrn89tJ0oK9+Ef5IZw/1HOvCdUeBp7toHQbCbHoXDUCffwGFifSE0
QYNOtHafZRz1JH1y8ncrxZRa9R8d6b/X75OjZZ2T8V14PBJO9hrTjAMhk8XfEmwd
YvZK5uR/sVBY+uKoDirSZ+pRA/LU7apqwvFV8jzw+fBx2qG/pjDe6brQRO54VcqZ
BFUZgbfnmqKCHJn+zu8q3gAMRpmsAmVLYIf8UqfK5hUZrhGEXEE43XUPfoqWqbu1
QS9d0hDOEsYtuWZV6Zrr2T577q2ndC0ORBFavAz3hloUEQVZHgyvuxYbkm9odt1z
cJqYmhaU4P2n9Zf7C47IlqyJu6NxFuTkrQfaS9f8nt5hKfvO6ENt6L1BAZycLR/3
u9iywku9eq2BteKGOzT9qIen/eVaDy0qHZO05mrBeaaxPsXF6S4ZbkZtS9xEdJR7
P6VvzH09YgNFxZ8yQ7wKsz+kME5Ctby1du6klp/cYeOazN90egwCdboy9QznW4Ue
pMWN0akWjqMHzJ9E0QZQLEJOHhatCM1ush4jr+E/JMHmZqH963JRGVMf1jor9H9b
wE88hrLVDYUytlq3z4WcAKDbn/pdK0dLJQi7aBFg7b9ys1yujU8vpoDciwpjpD+6
9oDYGr86oNZwj57TiZDrS0Z8it3CiKIfPlwy/uS9g4g=
`protect END_PROTECTED
