`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OkR64Hu1qHXt2KIMNDA3KPhz8z1exgG1PN0pIgvH6QSuHAfMJX/C5whKPf8lWxEX
6CSZLMu9EPxNOX0oO9wuo1tMxqyw8tYjUfm+izKkdZ/c0a188ikJlNj7jabt3zew
rlX/xDWAfVvLRXG1obN4FTk2zWbT1oWcbLnvbkPm8UjWkmxOBnpZWFsxm3Maw6WM
h8FIbbcF5k0/RPP/VrgLSjeJKx9o+/4tvsaO6uqjICOPuri/aR5lb7THVQnYFlWw
evWMCJYDmmZ4NaPksnPw41srFmJhid339t9I+OeoChVQUh5tMFnVuDi4nn6lwGCH
uCqAoqKvPF06+hSOJwcMOdAEyL7NdaH3ODPylNccmZQu7wxoPvtfE531y8P3NtVk
WOPw7HjXfps+547zPU/t3lPu5RAWKiFUGQYZ3ReLt/PM4nXa2gML24Qt0Fw+tYl8
cAr06eZbIlYNc4glvEzaG5aA3ia2T2r0DNbG1KsNCl3lAXCgi5jLmpErk3GFtMNu
BVm7rEvjSsz4bYg1OPE5a/hV1P9RyLrTzJLXSOH/ui5gDRxbA62dWFVLkd9UJT7t
0rQrzwWHa/BTE+sbKXO7Dw==
`protect END_PROTECTED
