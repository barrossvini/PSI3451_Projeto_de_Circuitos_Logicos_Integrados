`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hihVeXhqTEDMeDhgqlEw7yhxyVsRhjg/o5Xa3mHJ4j8X+ZSE1q14LKkMcrfCULLe
fZT5wndcF+expqUraZRu49C4aiIqCFqE8T3GNEZMHDso97HW2qDXjOMM/V7emFCz
4mk/5Hlq/1HE0uGN7+QjAvIWk3km9Sctv5ZQctoPGwk7upjxum+pimbzfQeKl7Am
e+k+JE6ekI6j8TJ+lryYAY/gS/i0X1mOrWQW1MZK8MSlNBvsoADGg/Y6CbdHdwMu
CWVr5TAA9N76++aiUqnAgGpTh1UOrh7CUhnWcVBTXpWqOVUp0259awvrtDvfh7dF
RzIUiz+7OBp0R5dEsfPd4wKKCFg82GE5b98joT+NMojs8YFBngLy1xZO0CSxEIZA
1rhinILSBc44xtASlXjxEMddUvxCOTwRUDLA94BWP6yHe4qlkVMKbiPZcdZh44jT
1Pm+4X7Ak6c1F5v08SIcUq6/TuezvNistEVB3kMs8dBws8RGjCZxVYXdSWAeOazY
WrhW3m0UiP0NFojg1Qi+LpaHUPJDd5/Aatw0zxLLB2KHY71fLAEBwV9JDq+TjP6/
mm4uwkvZuVhEwHCinVIgGDNWZf6JYekkKzuY6Jil/ScPeLJjaQM2+TW6raHgDCa2
MKMHaKakRx6+XAVNseMEKxiCRISTs/pvgC5zX/dZO2i03vMPgaAETQb7uztbD2xj
9i60ZKIdtQS+TyIw8MDGRN/86g77tpN9fpoLQmIG/E+3EpcWTX3teE88Y6Km/2qX
IszJ7UndgOcAfoHlf5f/w3IBGIzRKw4Xcj48gj9J7K1AJZ1be2utIqU7VgQUjdb+
Lk9bO41IhgvmUG4lBcyrWEBooCyPwQbI62tYkrILabhyPF/aCX07E3D5RqVVESZI
9LOF3vHv+wjgW1Ce7uBoC6EEMpELyT4L+SkWdVWzHAE4WzU1tvMBV15sK1roOYj7
ls1+uPgT0cD3x/LPYX9vhR+XygR3M7ZmJ1Jx5htW1xbVn88x6ecwFUh5VG/8Q8Kx
kDYB9SZWO7cicxSYzXLsvl1yAbHzvAAUWxgBmQS06coqj3Cb5kjrbYrpUcE5Tf6t
3S1flCw5AAJO1XFIwQ3btaNx0zA5YvXZagGXwB4i17ytn4evIVzceCSOdncdBfsf
iDlFKpn3OA01IH78THZDU7aV0nJopYi0vCSyPpX4TrQlXhuaeVl7taUHsulM/a3w
9ZwGMVeSQyNCmbIr314XloT44rFVeGLg124DIvDcJ6KAA1R9nsR8WHgtGxuBMM/a
/QunvUALG0PxNCjBoy6sc/yuJ+yZfLr9cC3lhffryFBqhcHV3fnu2zATa7V9av4r
KPv5HdWFBcO8AjphlRBc5F/caCe7spGN0f08SNBauUVn5iQHmORmj24Nv/bhKB2z
Qtmf90AZBENPY+6BJSH//LFdnMbfOluxvyklSeF/z1al1ScYHDTTL+fSIhD2Odgy
eap5WHRDTTxk+U+98R9xJT+++NqcVtGApI8F2Ogci1beweSOTc30dG9av7aNtEMr
IUgfU4ErlR2sSHvUqK8LqCbxXd4SYzllVtkf1OwLpvruYbNDFJLkAdaqyAOiOwgJ
jhU3e5JnrWQ1lOoKiFrtwDb7ly1Hx6+ExKnT7SPBxtDy2dTM+YBaLtXCMM/u58t8
hjsvqWZEcWYejuRfwNaU62u1IlHGLgqEKpwmBaWIFgtiuGF/I6SVxcckl2cq0J3v
QhtxTXK5SlpIL02BKjr0JbkDVYcZHu52SRRX8zqQ9hv7JOTiPyiqkC67NwretUg/
5pBDQn8q3CFtF52EqMtSmRMZ358Tzhh9iYn8fsRTzrHdgcVckjvJ3d1jvRGe0uvI
5azvuIBGK0/bcmnGOxiMtlnc8SAk3IWTAW2j1hS+hmYYm9oBxVbC9SdKvxA2mPHa
3tV5jzGf8yBe15qLnAwrz49+sdCUWkwqSR/Mz+tjuFrFykKgcqAQ/P6Iigd6RYQt
u0xML/nc8FHuzjIDRGjfRv5rFAq7rtq7EbSg2KzjlvO7Rh7OGtqRk66xaUcMg+cN
5vqh1amu64x37HUVsd74kIYely6CHU7/bSNf5cdKTj3nSV0jH3afrG9pfK+abHPW
J6bk85lGMqfWN9UmxzXFbQ/+DIfI2CVZbJ47nYvVL10L6+ezp/9wfyyx5ZxZUL1y
bQgvzxYIaDhiYaDS/AohJRXxk7UUbMZN4/txNwW+rdR/b49hh71DtVdmsKg4wfdp
rC5Uq+A/SJxk9jH7/6C0FYefxynSCjQZWR1DbuiR5m84AaRr2e0vXdsUuqmPqGiW
2zJFmRs4fSNaXCiIc2F9dXJ1G4Ecwl85cOCqcFwjMam0VE4SXikTUiXVrrAsJllj
s7vqMWWmN0T9C1BNd+InY8z/hTp/TW+umJ8/b8ogFYVHnwWOeRXTuRpnWFnJqaX7
C8u5khFk5Gwev/GSzIZyaLUzcUQAPCSiTsDm6D9Qv8gS2h6F3jC+35rBNQVsAzl4
k6di3rwIqu4h2nNHnEISgSpLv1HUjFI0RndSksxEirYaNed11WvgVkqfcaU80221
qDpPMUXHr5g60PnWexTL+zvnO+1jVnQ3OJ13ns5CU5oncaaSJPKzl7ZhoV91HWi6
PbCYLLcnKyQFx0ZnIXxZs+ON60KYZNQuRc/X55moLzlrH+wqJHC/CtB5ohPvAZiN
tbvPcEFYH6Es3i63QZcxO60yruYNackbpGQ4iBF9nrbfEp1J1O3ZdtXZHOfRrF7v
iqgnWh1fmrdYpy80/pWYehxYamKBeve1uEGaiziWyO/YlndJfp1FCpQ0MOSMmYQJ
hHvQnuh6eeiDEpQ/lD/zR0m7Po/WpBRgMharAzjeLwqgHatm2S/q+gX+mI18Ephr
O4gz9dBNIT0MJcFGomxta04V0i0+KVYpY/Tt8thcRGdQTbxZ5QIMzjyWHNtSuAiI
o4qUeEaa7boDQO1NEt8kaQgbvWZiGCmoViVlk2UYgZStDOu8OtBU/glN0F16gcMd
R4In6v9JV+vEbFTNPF6USd0edDpjUDWhYIeth2HruU3QaLbbTnVLYU1jyXaZIbaB
ZWDnr1WKw9ypT7U+R/mi2Rbxde2H7KRnn9sAKPSa8TT00sCjzDNAYmlnFSaGDzvl
PVw2HfuKAI/MyiCjtCU2uU/UYRHeDB5pACUZhfRpyujevtIVrjPSSGlmLdi4K0yE
IVyB4Q/Meayv6lYhavJRnczP8c+WiVeMQ6YOO9o/VvkerypNPvhu8yhAIZjJDrp1
tFbgPy805X9JcIq5tBfGxdeRD6c9ZE9/m0ujJOB+1qTnvMbFAeEL6Za0YcdFkIWN
7ay3IJyg/Hvjvzw2KmMfd20PpSOdIuik2YOtoeCYk4Xpvm6MXtka+P2K4WMOAix4
viICnUxEbADhO0zvsRuPxbJDDAuN5GKYEAZ4fhTqEplHervSUeQ6VKoFOEk1NM5I
pvXQGJc+4A/Bt8c4cBEuMmVZjlApTkoSZk8VS+cprLxU3esaU5qidmTbGxwspSey
YYp37dB0hbHLQTTDekaDN8Awraz9l4WZOj9U4KDo8ruEn5xev0Ah2pJhpQqHnUd+
vGAQB5qaucWzGg+c3TdpOKu+Kt/8DOnQ6xBaSoCQROZ0XL3a9Eq+jUWXu1H57L0h
jMloIedpRCR37uM/tM5TOu4HLjoeRqvH4qQkEe+QbY4LJLfETp512wjjBaO7VZ2Z
kbJUEYpbBb8f7MKseLUFyYeeoU6i3ajyCP3KHSxkrkG5g1XoutpqJz6m1tLXMAAF
BG8iRf8z06qhPvs7gfP5GcUc1ibsfmgxZ3lxrddwYSqFnzVaJ9/No9knAmRdAP1C
Gn2/UeAyTeuBLIX5C30csT6Z6HBGGRSUkCgoGg//UHNYMXB3GWrgppeRyHWnJx7C
Ms4l9i4j2NQ3/SxbND2tWA8By3on/3oY96cWesLeWO6O4+7icy48zIG3dEklDRmG
zqpheS1tFr9gbGdikUHRRnV6cFVqCfux4pHHLbD4avV3+NIE7jNgT95Ke5YtFuX4
pb5Zmlzk58xrcF6MKTcMP6eHeiH4Uu3NrbZCM8B8DdvBsfcbm7ZFtut79Bc3aEvo
Y8F5YpcIQgzzA+FWWlDUy5N3xCpJvSU8/l7QEtZ/9Jglfi5ZA3TehpGkju3MYoth
MEmq33Ap3503sy6UhbJhFYRQq9H7Z87i/8LU4Hn/33yE81AicjBe8eywJmAzKoJB
ZOZ/gUTwRTWGR4/yypdckI3fQEGFzsIWOnes3wq1cFj+xXRdWB9MsCFCrxnGp/IO
idEQq0Ul0cUHgPcwCiCPkWRy05W+3fK9YxlEhmyjR9iLXIx193RvF6fqgzhnPq6e
QvYWu9V5l+RSGHixRTaeueLfFawJyzaw75xAeMsKHINMNzx0NPx8c9erCSVHWXuS
Lw6CtQ791nUo577ksanox7lkCrKZ/EuiWJoxZn1tbe/2nLXz2EO2ugqrXu2irmgK
4lwTk1ZRuNKBMJ4NMn4F0ijpSnhCVsUmaMf5brbpG2lOQSfpxjxjED6VjCU3quR0
x4dfhGHUCP+jLg3gGxMYwo7lZjRwRkd50dKi1O00gLKa31tMbdpO9u8KRth8Ci40
CK8U0sthygon/TZuKhu7DGj9D2Q/GO3e5o5r/+t6Hm9dRJ+grZ58+4P1kYgzuEKQ
yhAeXODqx8rCO01Wnaz/tAx7p0qtFu+ogr4iRXPFZD3FvH1qNsxGOSOiuYBcKne8
bq8RgidH+LjY51VN9PI7mUSaeq3MLTmJ9NNrVjTbBbIput50UV1zVab4l27lzLTi
dUd9iQ9tVnls6VWXShgU1c8qP5usAxOnEWzZt+C+WvkZkmpEEtx6WRwRbhLNloXT
twg2IMgKJearo4PyMUjJ/UVhKg59B5Dlx+gJocP64mqnYBZd1toqS0LGZ5AZ+GH1
hwIqF3U3wkWkBqWjbPn8p7udNO9/SijwzxiOKRAJDk+IgR4gSJMl/VGB4U6UZ7U+
phcz50I1NbLyfcLdZkTzASkVReiwOuGvuvlDaCrdqWzKMyjO4pEFAU2fZTW7XKAR
qdACX1W6ttQlyshHvign7WbM2RwtoOdt7PSS7wbTMIB3GB4l4jMWsXvdtHH4X9cH
12W7a3O7QnIC0DuKG2q6dRa2Ioo76jFEcIjJVDc9dv06p1fzYkF+m1b++XcGvuWo
ax8t3gpBl5Vs9NyVB/jt5130FPlHhh6id39d5ak+dALLpVPGr+q93qZAd2hb4o3v
2scXA8mCjwSPrHSpDfn47RNmqsaW+I2pXVpLoXyYuGJZ6V92MjenJLZRpkQ3Ppkv
9dQVicFq2JkS4ExK8VgLQ3SM+c8s8Cj0AshlxUztZhUTzMRW+3VH8najWevbvupl
JRfNaHpa3mFrA7YWvJggVzRF06m8gMa3zqNR6iWHONw90wz94Z/y/u66y93f2XM2
E6DVgueFG+B66ErNHEuiHftfOX8Pk3k9FUog9gXq3T1JFZGdhf5iSny9tVo65dm7
c4JzIXEPtrB/WAU00S/9Mov4suzeVukMSRDTK4WGucdnRKDtMzyMA8G/X5kslpBr
Qp9+HHFE7eul+Et9q3LS+iiX6KaCsCcgHDyfIT6h6pfOl6VtuXDaUGJOBR117png
MbRycupT4yeP50E4iF/a4P4MEolx3dYNjI4DO59RAvvVeectv0HIOF4rWKRzb8kd
ANt3UxfLlDEWIg07R4/mCY+f4EA6Fy+Z3T9wWkV43J1NNuVeTk/pI2XM1dnH0g1l
aUhzciH4zGd2doiKG7Vki57F69CKLr/U6GO15G1XVosCAuYkxsFo4M5fJSCfBqvq
AYiHCe8/a5Z2us5GpkSBd14DOlmNzRH6a2G7f4swhaxIKdFn6bKGO9EkcoVjg+jJ
HkQPOBJ5AUdSlBGSUZYkqY05a7VfVdpb2CydcHYPwTk984qhvsEj0Tc51MhJoJYX
9EFETdHWpy0gDyR+tb2ajvTom61BCt5wf1aiKawULLA=
`protect END_PROTECTED
