`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q0S1eoZhOwhYITPiJnkSaqTRyy2RXFBdYrwQymp29I4pXzTmwYJOqbwfYBAzkJEq
iaqyPPgPWsrhdNwlelNPYOE198JN/h493dHPydeOj1d+hccedwjn6Pvw05SH66RG
9RtiWI55mTP29v744SBhKlN6YJ86iFU/Q4K/HAxJV2RVHLSXpTFVBab2o2AXEFSh
MlFHjHZOp7TvVtn7Fa3QdLdBq2o2tcacm2iS/zG9F82uBuSNyf0y00+OKdv+P0Zs
NPCtz6y/zO6AZAem/MVuOe0QUO55/xC2cQd1USO/aUHkiWYrkG+gKmLP9BTdcfgT
72lcJDGnZNv15b9y+qnIDY6LzDiUzxTukXSHgqDCsgyWsSiJeWE9R4Bk4q7T1Ync
Is6mL1uG6UKQSIq83ZWFxzu1Bua/0CXek27036xwB9QaLsBJmpCOEnBvqE0a5NsC
PJHp03mANn17IuSaj7lHtLfzJOLscazTyD6P6x9UkO8mAjkmEjIG/J5jeuclysQ+
pMvXVRKMf0PmWitNpOq88LMwPIiqhwD/Qhr5RPteg01azVVqo8yOZVro5E543u8m
Z1dFc+wj36vs3fzk/naTCTXU8+V28Zt+g2wMxwY90LJtF6dDgg77YSrCnVgArxDF
muboaEUWp3GTynCtb/3UDGwDC0G5ycAxkipoWiCbeDzL5JiEt5dWCuSM8Tote9To
aQ0YmPD/mJeHxgIejXvcImZ3rUfk4tRUKm5Wo6L/lVWfC/jAA0h6nZfdV9n6PvIW
iqtU82D2809dbg9XGQPcn5u2tnOMFoDMQmznJvhoMPHofVjdwG9EXIfsmsozp9gU
KLzztyIrTwukBqTnKufIIzdGl8VZQ+pbxDAkDtIcbbLC+cZt7BUleAwDkoZGl6Dq
jpE/08SNgwgLiACIfBsQuEgG0GzZch/6RZajjBMwxoxCtLdyefSbizz+gDZsRQGB
NFBjbnFeSUDuhpgqohjfQ5iOdmp4kLLYsXOPrgz5X6FluggK/cP5JB5NqHP3kDwM
4bhyYDaw6ggfp3LjbRdNQc3Ila3V6y8M60vSqzY+cUhB0tZz6NSYVAy3w0DpwmpR
Yzuf5AAB5WH+ij1FScRur3ltjTnOsFDU7KVUbvkbEX9WOIJxYUAuNoFJFXIVLkNf
DCsywDMKJi4qNWOTZNypezW1pshAioXR8nZ621/OS31nqAIccSK8OPUvmzdS2EQK
kU8OY0OgniZvIuWY3s+bD+xQR3ozXamjzz+CpDPg6oP90+Nd8lP8faQ6QZ2QjzUV
65LNhjTZ6wYxoSZZIJaCEaThPh+ZO7npUzHEEfvhtT0kp7guRBgMxquS0GURBj/h
jhXW7HsFsxmU2fJV/VF/SbujKFyI0nagFz0KqYu6f2yXbEVVRqWtdEg6mSTYBSic
+uh3EVE1DQWGN6TW1pEz9F1V1oBRZgZC+uFHTghpPb/8+R2+98szpRS2SHfUBFae
f0YgfuOMLMhSjdT34NjhHIW0F16mjqUUn6ZwWKnm8Wq6Fjqbgqv/U+wObI3Pnc96
pXYj9LocA4XnLXttnddPddVTXUYkUzVhzxHaiam8ZYE00VRUw74W1nE9b2VzSVk0
rB2Hd8Oca5vT8y3vMjRZZj1yPhh8kNr92jQYZ98rQUn6tT0sFd9BANvrybsPHV2e
b76Z0cPFTckBBa9WoAtt8V9EuxVEASW/YeM+A85PSfA+9Rn6DQT74DSlkneSIWqQ
vbC9MuM5a/oDXHsklBdH2A5MZIp0xUZrqPgpqWTNZhX64QISy7BB/fvNPFJQHa5x
i+Jg82uhkUeyUfAWf05QR0s8yIQ3aoo5CFbvGQR1WscPCGCc8NqNQIFCtRKbj/7Z
zAUbcyRnL7yWNu4/scFdeZCQkA1Ahpa4QwG0iYLfv412eb91ZgXbu1WRsHPvqQJ9
CiQBB3za8+6jJeHZBcPWLOM8eXSM1CyvqjYBbGGG8h7WndtDGZmIWyE1WHo02/mo
FiyRbpG92JZtywISATGWZ6Wd+lgMPoOcfBKLn8TUHLqJh7N+PZtFlMNgZz+j0dEA
ZKRzvDZLGw2WKK1RTUjgwFzMTgrFaxiMTxVY7+WnBbkyUAsx+ObtlbPjBM8ZmgFZ
0uZRV/VFrYuw56IEFHDNbK3dvn1r0yRRSWRaF6JzbnMWm13d5Bgjb5ewXR2/W3qz
Ai0h9emzfD2FCyrdo7UUOX7qDeCFohZaybTNWPiHqlTqbWZwqZSLxia4OQqfvu80
10XPtzKCQ3W37oyGDQzQ6CrQj65kSybC5G6LyeGT6biwWRYdWXvTfA9dlG/K3ejn
pu3EjMM5zKcThdWA08utXpMZo1Mmd+lz9o06BoB8Jw4E6fY8EuBJIuBlz7dqnRsp
xe9d9hjTVIcTWU98zqQPOne82nmq050Hx1ASp9do34x80WK9wNmK5F7yyUu5DH2O
E5G53W7u53zHc+PGyOF8dIpr6g5jmimi+8gH5G+EBf6PfrmVwXFWTadzpMDd33SX
XIoMF7ja7hoMLf3cycLW17qgo9adx4uCFv2vKC1uyQ+INLP9Gqvn76V2qU4//FSN
4+07to8yQOWTp5exOr6gjBmQm3wnaXJHzzFgBGQx1o4tH+SLg+ptp5oPyju1gmGz
qEyf8zWladdusw4XLYKB+hIiTYVHZUPwNsQ8ZepfMqrAjciGDIOEvuBKjrVOpyIE
UPtZoHYYL1OoyeavVnIk8sFxJ1IFiX84nBdO64faThiLIBjS/tckIILBpQfqdbEK
P6ECuEBu9YV8uQOr3iCuitFfAPEF6WZBRWGI/HGsTTjzjaySgl+fEefkK4M/NDve
mpIqiqIhe6SbsiaxSegAMUJpeOKd/RSg2Kf/4wCbgavsZoUARfsCko95dUZazP3o
qcZbBgk1dubaO67ZLKR/dQhxRPcr0HSrnWS8jLpQVu8ITsRA+yAmKBEp7YxoaoPl
WNPWrcVXbKpNUo7ZOqc341lhm3YJWyNU+13znfouvCwDj1pM++bLUFrgwdBIQO7D
azJWfkmSFp5nbmIR2MLZKw5smf/XXMnMZXESTAeH9xIEB91OrmWyAkbXjKToxbQo
r412C5GcL+cuXfjPA72X1kPFOSaVoxVLjicNo9/ho+pl5PT27lIgICuKAaPsYNkg
O2AwwITmmXTgcS0sl2vjeJP35WJ0/HO8qLRs43F+/ENh3q4V72gwpL34FVDtzWAH
FbENWKlQFumBx2a94gthaMOAW1zhhQvqISu7J/raWKIanSKHLW3fa8ev1Aq/A7Wx
khxlNBpgtef/KzzW+fZYGfJgpjfnU5EriFV+PE+y5ywFGf4rYQ4wENj7FGTJqvxd
rfHfurML2fHkPjTbTmutEt9g3AfpXzhd39HR7AaIRFhLaWGfbaY14rb1jf7nfoSH
nyA6EOceTm9ljLfmf1x4JsXWQa1QkPgqBfLgpi51uWAPWPBQeV2W1yzBa2fVteNL
AiWcDo69pXdMzFVlqLEnWbA6JX1UPMso1Z76QA/V7vt+2kPbxonOBFmindYSdLoJ
CatBaYXE07dNOZWJ1INu0YW5ad+ibKji2QehNrvWeLiAs13Rkfh3hCX9opOI9cD4
djo+OHJ3eJKaoB2AGYdmzk1fVJJ7K/vLnQMKk5yt7oX7QnlfvdgoisOQpdUnZysN
1k9mccS3quM4DT1YBUIboriFBtjzROZ3JHLTfLp9USUx8yGu+N5bJ8BtY8W0yEwn
9mzas8R+bFZtCIqxdFEF0oqblqvbuy+8lwhc/qD/G796ygygcNhP8jBASyBxBMc/
0iNI/SW2gGuVby6s0K5jm5TtC3jI9+9yvb650gNIm0cthkqgGgBLFd2tF9taexAI
rZ7rBmJQ7UW21uuwiEAUm9rKzqBZi1rfPCKReE00cpggX0eRzG/8nwbqTMoKDNjC
qXrScwwDJ51TqJ3KaCNXSWHODF7uHixstiv3QCx47zjKzF9USH1CzOsjLVpNK2Ha
OAPxUw5JayN21bHluRdlnn7Y8xLC6orkfosEOkA0lJG+kxUjqi/Qx9Upv3p/UgMo
vdEj5AymhaMLq1UDDjEqzhnokL8vvGTHZGJQPGKiZCBjVMRGGXtOyl4wx/cKz6Ga
HYPDmuBkJhnysTlqmFkGtq2+XlSCn0eFxxAyPqj2YPXYJWevnxVb7jSQAiVSCHkq
ScO/J1L+BakqaoeDwCXuUrMKnYMV+rFDQBVGLrggDs+by65xTqz7AmvziMdAVwm0
f0ABKh9yZ5lAnDCMFJxCMq21TRAa8IclKxW5UtA+XgmpUZNOHb7owo0C5fOp3rcl
2h2bPdg1JH7TsyGYQ5EqSjyM4ij3croQenN8SLr2E8kQYH+9TfJd9dN0f1CSJ6/O
6IHXKehiZOEqGFiJretPyB9zimIbtEf2lg0BE5hXllOvV7MBygVNQpLE5FO9fFHk
bJS/qxfR2jKHdjxpZDfVbos2wxmlYrI/0La8wxWljsl2I2yuE39tv5aFeYh8W4Nl
45QYp6CVAep5JLyhGakFpYgGXc6mdXzvkDn5QMcKjOdlSzKs2sYeGukD0ZF2gsD/
CvlD5S9DABZSzSL3oP/T1XMdZ/EYWuZ6UWxi4cNDv+qybarvPvahq1xaJElbS4/3
covSergp5CVRrJ1XePD+NEJDMndGma8DdUH+eMfdmaI2h7QquRO4ahQbWEgakZlS
g34VtOjTJofrgpQ8dNaujqRHpaVeYENnJ5GJZzvboldcfruYCiHJCkNDv26W98lB
P5wthgcfxYITs4zNWpNY5oQTHholiRiVIrjhOjrP2OQMI3p3T8gVmq5n8kOsPFO8
Yad5jyzncneiu0qervmZHDjrrn2NuHj40Kz6hqnjBvYrk0oswvuayNs9gaIH0PG8
DyHn8qn74k2g3clNGdPEpIDP2nbXga9YhBTXn9tMPqAwZdmdjM9e5jCxsRc1GKLH
ScPozno3MhMg0Fh3FKhMzYu9cWAv+KoVvxqfYxG5fPb4Oa4k3lwzmtDg7l6C4h1y
/+evwaEP9KFdWCvnQdtglDJq2wudRF0JItJ4qpeNPJqZcbu6z/uGajlR/N0c0rTt
eADAEWbU0OfXcoQfAGLcsVHHJ3qYMnPU+E7o+ZRoVxAYk82PgFdVVF96m6Vg5ZXz
B2SHoY4jxP9w4KGFJUBGPuRnnOsMvz98Cuy65wjkHSZRhGIpWFYvAhYJKRTQ8/qI
scoEH3Y9sBPc4uAXrsJjpi3mbz7HbPhzeYCbs4DjCeJJrg0YcAoMdPwPiMcjbis/
6L22nxgjQWfvHYnOntThhkmFgtzVypzPRxz1CQ2J8p9meXYMZI39qQLlW7kuDsjX
nmrhx8Ig2hp2uM/PAr/6+5Ah4TqmlytBDqMHtg6iTKIJ6mxyoMut7RMbbCohid8c
zoZq9WdhexY2KYrhy2kPSMgXxlo+QrWRHQh/nWCHY362/wCaDsDU82J/e2J68Tsm
dUa5kttt/bisZSSPYpPaLK7xbNAZH5mNO3KNh3fqqqVtDT4NsvcACtE4pe1UVGzE
8gBVAxzSlrpE2YtOJ9lI1/vEbrs343hCmQ5Vq0RmAQyJs2nOH/o/4fO1SXYWvzYe
iSbHdeCrxPd6EgexDHgMk0LMeytYIaCBGBxLxJ26o9j0zQ//VEM3XUzN/1Pv5zaX
HiUgmKjV2QgNGYpmOigoKjBt262LacmGd3D27syKa5i5ByYawe8/0Z0ImdAwjLY/
7Xzr6A5UUcIyoQAj3Ykf6LVdcCRgwlzTQcuwkqHGYSbmgwLf2jpO4176pdZuJLUM
tIIlw7hS1gD23bQ8Q0mbE3vVe9MUpj3V51lT23IS1ylPpfr4e6mQ5QFGVwUFr25a
gNAITz6d4PhgqfD9UQtX2V5dD0RxyDH1y/uyd5O6Qn7fo924BCjX//tjAOyDU5rl
VKOslmtuS2bskWn0MqBrs+WFQ64lfJifPja1ansnFZ80YD9I3P78NVA1/u/AWwhj
IdhCQV/+toMfxDa6juaO1ERzt+FGLZro7+KeDjTMyFzQhz8nu+MM9DhhzYHIqM3f
oFo5iajkAmeKhCCY5wu12HR+HAvCYUpmjkhfmb5XE/qId9AwNPCYITRZDBShVhIr
7pC/AjfgNYzm2jHgPEyNWqpH3tiQuzi2F7BAYqhbfTfxjY0IJWXXzAJdfhELkC7/
EdD8j07f/M16+8OjPv2lI8qRqYg9F2PuIJ1IiQSiaOWbOPDb5FfSMqLhNWX6P8ur
AXMkFvKERBO3ESRGA6vmAJAla8lYJPlHR5e2vIwbxUDjKCgRDrokdnH0UGIZOoc5
kYILQZS7Vqc4NVt45YzDQrULffGZVP+3v1TpNCDdwIg/6FUBMNQpufT5PeD1IbyQ
ltFV9L/fROZ1nCY4ar+wiNQE9e8ai3epodlda+lG42JcVUv8kgUEhPO/9Ev623lv
4ngpbQcDZhp765U0JHS3rV2rYfV3BybtKdh+EGBKMSDoPzA62dSaF5mWQwiJTUdb
JbHBr7XE8Sw2uiWlp36jL7Hrutd/S+g19gGlTeQmajw2LVHArB6e/C2+h5rhhu+7
03EA0GoYh1kC8v7uk/lPeB7wJEYbmNY1LBax5M9pE5ZDnsq1/8MMIvJi6v0pikH2
BfR0QMRbjfmGmZn3gav8VyBLR/OCZdlQdoYcRIUH+Np8I+W/0MZY/zkeqZDRs2Iy
x4Qvf7wnva7elVNoOUVbGXWD+lqYi2HJFvZRe5FsO/I2t3JVVFQEa+DR9NUMCaNW
yDW4RkhDKqku4/WBrOZqjcAcMnS+oboUMlf+Rwyo5bZ3QbGO+DovKFISpujRPIv3
E6WTwKaE9evbk1KJARkci5AzakLDaGRkesPHb+VsGk018n4/Vl02lUAJWSCuDWv7
aTEE/D5xiSZ5dUKZ+57zQ0gpW9VucLgTgPZmkNCTdi5E3Vko8/odHq8GD+pQUC46
ZrXFsPxGeoR18+KG7pbPZJBU4/uhlvTjaG3fLGFb6TPuTTNVj7nOk+wAiKF5hDUU
XiPwmmMLgmeiqk3x3YIqy1czivX+LZPG8GEpFbMRwiNjmHxv6z1fWd8kUKt8+hWg
MgwuXt6YBDRT62c3MLLouHUN0DLlVUGCqu4drr1Csx2KdvvX7ukFAA6Vz9/E5jvW
daJrt407WbGUFBzXTv5dp/NRXuwPfOzxuCpxLqlCuk3QIncsfog0UpNeVUB7aTOh
4sc1FBRMrfhLVELiawmP0hwSEo3Qn/Dhay5hjfsnlLpvIdTQBHhOEDvV6cPi3r4D
wpYkXbH8UVUZJ7GIupm2IxLKvGCQPHh2SVQ8sMiYrU+LwZYOcaTrlPqs/93UAlTS
LxBl1ReB7MyWWp1bXMga6CwhV5EET7GwJhKgXW1IoTv44ioRIQ68d+RwzUli6RfT
IHMpYgFy4tCfkX7wrVwJwXo3UIf07TQmEWJ4lGzkUFfA9otStNi8gTVr0HrLOa2z
VwbUHauYQ8NwZqyubck6Olj6RaGiNc/9vrjU8NnhFyzfAR7pP20phGghhsmUpfUj
re1WN1NPDM9C/TNi38Zkwe4QFMPij4k0ZtxOYNrPC3lLSQqXlgDk/R3jVHfC1vYj
AyjUJTBqwp6LB7DAM9OmrhcnJuvqTft2NSu+NrlYDwuyjj8Fo32x/jModpQGgUdd
YyttRLdJKj2At0nVEj+M2pyYu9cZORfw/22leCIzhpiKWbwEiE1Nhi3jvrZXhQHp
+MVyIjXrqCYMZCpu+k+cPWNxFak8ZM5p5nR4kK7swl2ZvorqfvE67KcGds5IiD+o
aL2SeTLSyNqEUSaxWAZVIfZn3Xgccv9kvFNS04gsljWvTK3GvIbnqFB7cNQssJqd
IO3raDPKkB3vVDjY9gl6rnMnrSk4p03rZFXfvML19xsBAgmN9R6Ae+5hTzgri7HT
I3yFMBNYfxjZ4SL3UEf41D1VpkXqB6yI73xw5ybilO4jI6Iq70x7ONpTJVtxmwKI
2nCtE5KO6nnz5OxIBYfK9Bg6uILxEwkVhl/ZjbjQiyxcEUX5Shl2slZgY0HwQ17t
djz14J3dExwsUGmKWjLR7xTnWyY+OhfY9jOKjs5N0buYzRz7FndQdBNCI/gjXbVi
AZ6h1X6K4aYSYEoSG7ioDAPwN9hiB6XsQs2npDS0otN7spBXZ4Ihhav0Ammv/1lL
X0UHivj4L1L2MXrl8W2RUP6ERAjdOfdlcNSbqKB8AxHqcVSc/XwBtxLwTxppgTQ2
u+/4ADgdNA7gRjtC77NfETCoQafxxS6ZgAvWGNNdzmrWFRgxhnj3O9w+HENUNpZE
9SmL11tnyqnWMXCc6AhJsZO+mmYEk+KIZmlPfbCNWf/3ltL3h7+5XN9CFE2CdC8r
Br7YF/r/1HNLc1q6tw/x3R2uU5P/x7C8yGn2IdXn3kBzW3hKmWskKjajbio1ZyaC
WyAuDOjWeq3jUxSY4dXeic3oAd1ID4km9OYdCnPm0n1opwpz3dmhg2+7a+1thpwT
sY72x+HwPr9UKDDClJEwYpH1uTcaCt+DQT7u8IUwvC4kDrQ+lHhm1pSkqtbtn4AZ
MpFfuVT7pCshG2RvfcewHlPihUjv69R6QQU6wL7KLvkPNskn3poxe830GvYTDvW6
L4mBfMjkRh8V6RSaHj7eO9XmRukSIguj+ewPOPddYNOrQer/aTMXZDkz2a89H9Pi
V0dxU8cu+8H8dKe+1yxrMi67Sn0Hz6sfp+KSlFY0LjsJsC1kWJTa6N5ax76ifjKT
U080qS+UWIJdKYSWpB/3hRACS0K1w9f16JUYD5fK2ieas/8L0fcVt+ut+YTJl48o
KjXaIdvxYYws8fXTNoBWCWERA5qgjcGC+R96/bHswDwscmdYQfY5j+FEIfaFwG9q
F8/CgvQP7wkFknkMHEmYG2DJHyFqkOzVatFtK60fVVrFDuXAa9DOtml5ACEEHntS
reAWd3VXQxN/MidIVm0OYfxUoneQFEw0P9P9myJ7olUkFPRz6NRtaq1HkT6aQdhW
deddTUFdwVfkWzfgCM6In/oI54xSxX9jZxpifprH1riPmaAbz+xzSk8/oLWmz/kj
3kS0CxqC7MXTrv+VCo5QaiDImEEcp2Clj4WirWWSh5/7GD9nngKdiKFqceTVnmPs
59xbGjGZQNwnSNHLTyzl9k3vSoy8SrJeD8plDtk0kYhzBlVBRhqp3m8jw8fXxRT4
7vFcUq0oDDy0Qh7zBORtVarihkXsU8B/FaKWRgCZKedHP26kftti8uOwQiMZimlz
uAgbXHY1mafXcUwlFs8A5bfpebskrUn69EAzI8B14CaLEsYVasca/4TY45gm1MWW
70U8USMVOOWkYDg18kaL1PE5aQ9iyIK/AsBrlpwrVTvOKMd8//WQoSK66b7G4uFU
6cnYJeO6ftOYOGkVYYPMK6DHQS8G3M+PkB60wMwyiS7POxmruLK3Np9fOHvyq48e
rBJhuwLSzYfvSEYalP9YzE//AImKtu9zor8ajWcCPbDWFep9ctyY85XswXqXigpC
q75VCsoxrT1nWGH3xQ06OlrbJBatBEN/8nPR37kgZie5Lq58Odx/icCbE+xV/Kv+
LtHzq8KysRvIf4YEUOlsfXk/XN3ftStmdjZ1DalPn4tTsUTQiaFzFr7UYp45EoG5
I+RNZ5F1fnq1oDCewfDtzl/iKnnqF9HtEFYHhxPSkr3J/QhQ79NvSdWdvLL3N6sI
KFEfysLHgZKKO0Pw9vRozOmIdN3retGdybC+mnbCbWSqzRJOJUyA4sOzfszmtfh0
mXPuW19vt1CI4KpUGJJkgT2SjvvZFiK2vzGkwrN9zfzSbyCqKyps6eDvKSVwQUJ4
nbI0UQMwztMbLBkjeK5tocHRd6rayy8ocuqX6J4is36MiPW2UV6tgNuvKFtjarF8
1aRZw81hnYR09otbp8LEnHHdpZul5x6KootcP4zsxlA8Cijk1kwDIZjesuIP8nk9
+pkOeh7bxaD3gxe3lGBsPDD2UroW1aPhVu0cJfDFK7laubSuHTCzr1t6wL2UOIct
i7UXbASZ2s7nWP4y6kuL+U30UwozIdraNrHTfxEocSqnHnI4omhRBtmhVx0h+QbK
Vj0MjztWsOfYcpMjVcZ9L4U9Wzx4/TjzWj5+9ztIOda+zTNNzvMO1zt4ZKo+Hmp8
xxYb4tEW+l2oReIpe2oItiz2MEMQLhDh4/qMrIZzDgT4KqBPw6vxQf+DUUS8915B
882YzYvAT1QOsJnRl2JUGBnsZPqc/mSsitf0c55Kn6F/cgYRPRQOamZuRNgSu7E1
ZfFLIdOBapvlVoaGT47d9WsXhechyF3CJBlznzdXBhy988+p0QQ/pnCpZ5S0sUVU
XBv1+Jr+qoPepae30QMdX/f324OYfAk/1fq0Nt+y5rjAqOLIYUYxcPggvLBBztbM
OIZrFngN6uywRroQtfqf3qfMjvAWATdFY8ANaWCLGMTGJ2aw/pbYQ02zAO0ExHzi
/w6Qmsu4soadr8ChvAmgCehgV/2KCsB7XkkBsmLEwNBxADWRttUcrOwP27WRmPLS
Zh3nzO/epWsa8M72GglprMfjKq8eh5BL2EkEEM0cEjgMVid3O9wksUm0EMvL5fmd
7OiUtO7BEKvLGH7WWvZQJz+AHN4giblWItkGWR2ZRQcQ5lxXoKp7J0A+RJkDkkdv
PYbQa8cA0dBhfQNtocZioVNYj4ahRZmNrGZBS+Ets1yC1kCJNiMjiVXQ5/Y7CsBS
IpXL+MsyLCi2Pqko7vdFGZpNBmGeQzai1rcZfoi9svemg9z6qayGadkBHhYsd+VE
qiz30gvWVWXv2VXQtvCpEyGMinmuh2tNIkrU9lYCBwtg0KC7a4BGUGP0SkuhtbPG
kSso33uAlZAMQNnYyBWjITJ9S724JGAvl058XoVYKHOByhEpWOWGYj05wpU7Jl/h
vpN9WIVh30ajGwpBQ0W2cAnj5EGChSuqEdJt+7PaYUGROfSlv0AAPzjEkl7Vu+h0
FL77Cux3xWDpkcLiK+hvSJ+E+rC+tv5RsugwFzLCq+JaiCLIcRmdk23Ll4XZF0t2
wdLylU2M3eSsFn0R1YDoZYS4qVOFSCNOB4ovmCTt88kLJ3f2yC+LKNusDzm7pTS7
ibshFFYzRAkdkJBXetn32L+0QQhx1Qv6ra4dGp0/tbhrrhzu0Np/B5l/CN33cGrK
kTm0pvtn+H7/JcmN8zGBavcMsQQ59l1/ph/6IGFuzautQzQ7UAP3GQOqfIxQMUSp
a9XtH6nHCbNmUDgeIar7Z+PpKVgNAjCslabS+6p8Q7yJDICmOsrpS5JaJtZkzIgI
6R++vypULLKPzagfTFjTQxu+9w6uEzXU3Ebc/CQ7c2N/vxZFi9IIyY8m0kLvngyw
7jWW9khxanM019ybgNe1LWKUBsl3Lyychvi7vWJm8ACJ9jOZVYjuuEgwg9h9M/FU
27lNbcOiIeWW5QgmbXAXcdG4DgPDaEn6n35lc1lnf2TqV+CSTWYAGA0gNnrzzI1T
WtAbc7USFXBvuaAcGIjd/Uq9gPjuv91cY9mOuWkUz0O+hkKZHuECFIH0i5i5+YtF
N8KntqbXriIp3xO2UNx0h+ZVM2hjy0IThXrNiZGigx7EiJSnXTvBxCixEdU7HbcV
cRg3O5CrC04SZTcXdhR8AlG0bTpaytwN9t9JkpYNWs3uCZCmuzAbt4K011vnAD9H
mYpodhtyhEnIGt61I9gR7+rAwoNzW8eAut1iEje084BIfn4Knzvajw5jBpW7WziD
MaUG7z1oug5SIkX9C/6H5Gy5JA0qig+D5ZuOYzKcx92FpALS7oMO+os+SEl6ON22
yAdf8huxqArQOFjYWHkWF3a0cORfe080RBcbxaRfuY5ZfZxHdlbQ3Zipn0P89ndF
yiqqOFwM9k6cCVAD+BRGl6/WxNriP/elHrqgHdFhHRhuYNIQsNgHghWuK+H0yN7t
kanLEG0NTyKG26nEuCbfRjlIdJweGxTiXoHSlh2BOOQ76nbUADDOzx8BwtAGMwYb
MYwNbRLUbxM2hcsi9d9ZJ/Yoy1ASQYWZJmwlEa6m+3G1ZC8IFEfrCNVv0mZHxF+i
OjdVsq3yeN/hBjWla3JVaLXT0Bt3gV8tmW5qCqa8cU0/VvKSlQw8DrgHvisPDIpJ
jKfQY7vjWkxpPCvIWsxdbwbx55TijCQY05CVa0wTaQqVN0YvapecmXu/oetL1Rsy
H/vPqB5ca2Kk0bvakiV3FsIG1DKjyidZTkJrvk1LBhJDQEq+JaKZ8Cf7ejJSRHqw
hyHDXSXTv81FJjd8UtfTAfYuzUaqr5Fp2AF8ydyOHQhgiLJTKJHgPFWHtWNjgAwP
NreSsRJsh9GzAuDHipJpz9/muuNsHIEt5XOKL6PLv3uNhpz55Op16bkoAwvT7J3x
mq0TRqTiqbUN8ErO8g4huesqb7E6Akk2KJZpfgR6149qKZFIJvHLx6j9spEWvy5o
dEUXaJPPMCHDNwKF2fYtx9tLj2Nq8lwso5yVIJ/alEBPCi2LnYbc9us+Tj6wtH4s
XwHDwu7LGoA+tdiKdj3LVRLFbv8rCKby8mK5rDWtmu6kd3xGb1Q3ebDv20jxPnLA
RtWyLntqvc4OJv2C304/F8Rrrw/I9TQiUoER2MjuvJJXtJLpX2xK4N8ZteCCr5YN
iAIXlLNUZPf44jnTxLuMO0zPcRxllo1m9BT/N+uaJBtxlPHUL/xAzQCJpIrUFdg2
vo/UCsj33Mucw5BJqMAG/eCyLIz72y2612qv9spibN5eUnVjsDph6b5QhPN4IOIe
7/CwMuCbNwvqBWc52+IgqTBIon4vM/ruO3/XWDaudvGlB1+02mcuMk4Xm/bOgj0P
rdAc4lElslGkti5O9O37//Tk1iCd6pc5YqxVwl7NLC2t/oaZZz7LXB7JbCHIguoI
CoNcoG/UdSAn/HdoZzsx5WrHM6UGPpYLOZkknBEIHQQCJL+sc0JaTLOp2xlCzyFt
kZfFqqT+MszHIC5cyAKkirzXBHSwWK0q00ALWHg17I4XMZFEN5l8RnY1dOaPHnIn
og+8D3bglaFpw0dMq4AB06opIlEvalFPFhCgjHxVLHNICXMmUSdmVtYxDoGFuuIY
9AF0lsWlNoVmjsMay4z2TmZv0nglqAtMz7u16MH6mIZ2V1rPun8/Fp9DSyGG0gWq
AP0RUZiTiCptDmrQFvSpjpZ8zwbpGqE1rcLs1F6xpCqZ7O7rIYN3CvFIb5DSvK7z
SthW91ViVLTjv/t/iTqqeuY0SQS1yU1FMi+tMt55pXqc6SQb5VZObUgCEkvNFDuO
RzIVlgPiQu5Lh6bAsKZgg/8BLNdNok/v42piwdCZ8skPKzOWif/nZiOUVvbaDvs1
5ldj17zkfYSjAkx/KQWC7Oe0lsn7hzCYxjL0Hlc3HIl01rkz1nxJBYoWZeKJS6Nm
7zw00BsrzR+ESoMNuCrW5a7k7Y0ai6yg6t9Mvr0UiMPbhHdMCd1CDg+Up9PKUQ+t
ZVTSf+OMXdZTDS/vMwHbhjyshJliXOiQ/uTxWJ+U6v+abdA1Me7NXLkyXLOwy10k
OElUK8tWLNVd3ghGjgmrdXI7/uQtyZWEmdk90JOevWKu67vH2qxRjgVGf5eXV3ll
//t1ydWJj1uBXpsdmNR+lbVkobKK0bapNy3lBb1uSL/tZlFqJg4EQvjfoSCqDSS6
nbrmegfEFqwHugeBydfbLTTN5JpLmR6Q/xfnieU7c3dyao5OmPGMTZf3CywSa7IP
ePnB3hdsKrjJsPxfKWNgLMk4tlxB/dF4TeuRPMU8Be4MFiPpSQWIGS/1C3dOcM7n
f2AgetTEmBW6YxQgPLbRyJiNBzH3VS+asbnP6Qpm4tIrNBkBQGg6/RF3XM9zbjaa
yr4L4HMYNcERky50BzRqv5qKmoU2yYyS2fcyGS4QaUKKD69ZP/GIcoFTF7gFdatR
pwKpRo54Rcq1URtq4BCPCHuIsFAnY9O0q57q1MClx8AIVhANa7GBDaZQ7GjrnP0I
B+MuPqAO2eyprQHxBkYt/rqENtWpFqU6rOC+HNfefpeEiXxU4MX27IuP1+L8Dtkc
rULNtZflSyxLY0YPPyqPeCKzz4fgGnhToAzh0BBNRm8r2Wk4BPtlsuOQWKnhiEly
XTZ1lNDE2OWulK3Ob/xOeuiiuNx7aBlvEYk73MqOdNrGMvTopQIjvfOCgsW9YFle
HiZuxk/Mw9z2jpb0ENv9Us2gJUCteXCuD5uCagGIw3dkb23YpB3O3954p2zpubFt
tD/Qs0A4bbgh+n3X1gwesgYpaLLAKWb8N0UorXseIWsz5HMUqJnubzlfXJ3DukjB
9OrW3ae7zqAbdjGJpwNZKdN6y3GMtsZ5gbHDDNVzd0WEeuYmO0/zH9ET/fhXRUY2
OP21M1Kv9Dq3kdJUjC2hraJ3TEGUkZycNKLfiv0gi1uAeeX0Kfdn8wj2SHhQnaGm
y3vfL0eS8OA9jCf5txcBmBFSVZZrtogZdS9pbWAckskPNzyjCyprOBgObLHSN/3p
8WjWCEU5I2R2VpbkKBM1DjYekvVGbV9ocYsbVJpF3dS8uCkHsZWJmjc8abY3JRTh
NMlm3wIYePI0g7Y0D1hXt9vk0WbmsQKr1weCfnMMJSj+ztbryDeSrOxFozt5stoT
0B6rEoLOdv3brBuUj91obqOVjMPfHl+o8UD/XEVfdBf93kpnKSRnIyJs+TdDFNYJ
ejw7HnQFsFuxNKRYqWFwyIC/MAxEeMKOdMetkmqm916QYGZ+qtZ0cx+V585PEkl1
XH8ejvBVfOuuUl2pvdeNy83ISzyQxkLmoa6mSPoMG/al0+zot1vU7cnKlIh/xzZg
iNecAiAuVaL9F8vHrnYHMjLNLnUX9kBz8XOzkE1Qtw5n4RbzjsibcUxk8aZeociZ
P32mYyN2cYbPwseoY7ZFZBMZXoQVRpnFEuMStf2OcdZqVQkgRkofShl+NeFonlaE
4XnJuqKcQDz+5IlJmjsv+ZO1sUPvwh5Tluwdx+9hqkJ38yoDzGi5Ja6TbPznKhoN
qR85/210wFa+QFLHMQsC0bLNqSM3i6wvqVPaJQmGlEp34OXspIQOUimqCVk3jPvk
pjTy5X6W8KNiFMRv57oBTfe6DEhlW3N3f9q+QkkPKuQ/qZ25rXZ5uqHvetJoTJKZ
gUzde99MDckoL8LtKukGrV2NGG9jJAvdKhvf+BTkPNMT/7tgQAKQeCKboAbUXmvP
6UIDVEz0n7FVE4tQPt1FfrkglxAiya6SFE9rlMQ6hLmQJwIzkSZYP5qNPm8U+VET
tFl4z01wnSiIWpMQf18rJjJJTORo7V5i3rBVFPN+gakX2lHJNmV5P7YYYhXXS6rB
H6chhKQzNoTaa7oLRuBFC9dw2amtaAcBBD7dPdVZmeV/k3bzD/g8YXFI2dKSStvP
xyOu7UmRKkjRDsPnHHde5CvBnpTEDrkoZ4C43i8/J5t3KWe2gcnh8T0phEBV0Qbk
kYFCrvxW/fvPkTdMlvFLksc3Y23ulp+jjGUgpxuDITKbDa0PU6Z6NmuaGv17Cl5Z
fijYRqS/t/mBpxF5go1gKDVSzUiQ/2El5J9lMP2fpF/MaKemnVLjjt4g0ztmPp8c
7f875iOplS1hi+OVjfEHj6lLycXQc3+d8xUyP7Q95kI6k00qGHPe+d/nXBUFduqm
LglZ3uw0NDPRitRvlN7FUPvPPkiIzH3WotFQ3U34P74CPovyW7FRq3KtYaJ/zXD4
HKbPyG2RsijCqIbPIkP4zVnUlG47PzFPdSp6dFJKm3jyen5fmrH/RdEDi9EUqyQK
NoGkgMIDCwbXDtiQSgOALE9E0laq4R1TjIvH76L2NgMEfLpjmGeGo/hRSyafCgm6
XC9/SQ9SGPEq9wIzp5MR85KTUZkQtDTPYEqeOY9YobVTsyvTqsJZduJUglYPX2QR
1hSDGh/syVKUGTWtOXB1uCM2WNlkbPdm7y8Z33hc3IP4eXtqsAECkTgYMhAB6gIa
mjcozybu1lZZ/oF2x1GXTmCsUrZejZh7Su+6PR6oQyEwnZw/h7hEXfJFRzQHJEy9
mF2TkwXEJ+wYT9G6dm5rty4vxEmy5IPICznOtUZveuUmNxa7KQCavVSISjO6rjeP
Cp0jZ8+dUXxeOJuiMsabCztMhlDZgN9EBHQFJmFQ00k4mdYGaMkv4YHPhHkI7AE/
Wzz2Fo7GKgXthpMfm94waDp+Ga5GYC15I1J+hhiteHRWhgHXTvg1sSjPIor/EWEC
dR/s1M2u+1SS5ATgvuBk8zOPV/HieUYi6HJkeyvq6P+K7hAwhqbzuS1sCnhfM4Gw
gnLgBtZv63z1EzJdr0RnNXNWK7YtWPGKs6k1KeeVCzb63++U1hOISz1qcjiKNuOw
oiOgSN6noPdu2LOIVI8m/qonOOmaNi5MGN6VkhZJfoOndGhpxgrO79z3ioZQ2hfV
vtUYuFit2pMZyjU6eKgJbWkTJgQhr3YU95EXtfu0p1RJbBhzkO/Py1vTiaWNTN/+
quK/MQ1sTIAdZOD0ErAHVYy2Bz8F/3yB4AneZlNoHxnyU8rL7icmIUYymYVPpEgW
73F6WAMLgfH5gmGKg71869Gdw62QlSvPtO0cZwBrW3NsNvbcpBUEm+xClTmvgDjM
5772y08wpzDHHcnKtFlwNI4kDpE0xqbtqBZAtBFRa1BHV8OQ42SniLuUsQ+aMYvR
k/HsRzBrLN71aKbGpGkLiMGOAzuOWV0GkGTPNjdw6s2+1JK0cqg8CDChonBhitIk
LyknaqhYmfkFTeKjeHchUehrVKKyX4+BEDSsdHckGr32WUNHOw55x3CKTbzzWLa8
8eu7IYyAN33AUYWmMdNvcB3StsIKXIqpvi8wyrshpkdnbGdP/aAwlUDa/Rr4yP8b
Ef5fD6o5wL6aKwJdV/5Vu1TBAU8wi4JEeOdux+/Oqb43KrWjG0LH+yc7CT3vsgre
xwfOwLqU6iFmr3Cdxpa06seRqOuO54cSu94sYGUVq5MZVTxGlKKkfpx+NEAN08PA
Ok2jvPAdKd6XX58eqCgUGI3XAfZ6DpxiLXxAgP6Dt+3kmwHEfjjDuV1kksThBJVu
q/hsj8rSwYjJjXYubD3mATz5ehnIS4CtJ/44QDCCMQhIdqu1CB77T7AM247EwnjS
z3UCIjFF76k9UTMLfkegpVnJmUgfWk6fwy9P6fFhaHniqrgoyXw6Ye5fVzzF847f
E1ljS84P5y4pNhXznpDou7Z8T14npupdv+e64kEPvohGcFRQthjYt2gLx3Sw2o5a
IhR79A5S5LSxkT/fFEk64VoaimN/BB8lk4jJzLxAjW6QwNVaSAegly+rJklvsFKW
MFusm3jph3GWgVX1kkRiO6NsGptR2o912DLrHuSy8OaabBKe86RSUlvcvYrcU82t
ZMCbrQZD64SWhx/TVp7TGlUMD9fUDcu1cWAlgCgs1b2iXoG74donhpeXtIyRYPz3
OanAifSfgvK9NFdNJWdOQFu1ekjx9f5ewEiB25dUDf+0FYepX/1dAZ2aqKEkXWus
39tGL9YdSJqQ7yf/IEzoKZFFBjPndEcpu0C6nsRP1cOfuqKGnAWuh1bJHWGacpkH
B5gp8cDMA53WtRDoYCRnmCrFR/asVoki0fuvQssHKGLsE4kuHlBgMwQrdFYZb3BK
GqoVPMfChp+ATq8k+UTLs4xKlticB65FsC8u8hYgVM17CjiHnhYA7wn23h8LSHun
AfdbXE8CchJCrzi1lVeVKqG9YdcOglbXuVJ9mXBFhdcX79XUBoLihtQXd84r5Wsy
9Rtkt9CZh0g9JxuITMLN5u4EsL6gLNvuOuTi/KzC3on1nO6PjfLqDX7vew+s/Uwj
OAhuLSztHDNPfTa7ixPW7ceY3tbipnNLRnWL71eslnzwq1ugNGIljsuCS7WsCmRc
AvV0RnbCe5OKTBqkVZtjMjYiVn2i2I1tc0kGbPxyZeQVZ9Fn1mPRAluCDEMuuq3l
fkMeeqhXXtchLRK/uGHQIKmnCIg3PctbHnEtSyE67ubs6t2I/OF1Cmut+ykOSLUQ
u8Ugsaa2Hg3zQ05bmHz1W03qOUFdXlijtJ+73ksK3JHXK0mte7EucwJjCwKdWqan
2J/MWK0THNnGTAMK5FeWRJELeGF37qw03ZP+2bEPfuw4b7FqOyNDvYsrFb/YFrz2
vNEFCuY/38CZ7L+PrrZyJVvkNnewZD9WzuGUKHeUBce3ueexoLfzjrqi8Go1Dhl6
vu4LPQpQ2rSoehTA5rCZ9nH3dXWjb39e2D67Qtjpn+pho14nZ5fS5G9FOcL511Z/
jNSzs/5o9XHvTYo1RqdvlRwDhT05ORMOPmJZhpfJDK/Ryt9wFlFbS3hc2uqx96Fl
ea1am0u00tClrVYcuudGePpRAxnVDrl9U8PPwWvsndBamXP6RktEghWSYtsjynYt
lBEJ9ja4clhVF0hC81P1ajgMlcisjPhOuUqVcF0N85TzwV0s7sQWHcx5+gDdaXRz
+HPH9VZ1vZuQGtli624XqC39qoGyhqQ2BQcRZX8rCruTvpTXqWKTq9SlH1MdYxF5
TjKfzX9QueLft9dn9nayLHizDkzK1mDp0+b/Sn5X8PE3TzTz+YWKXiwWvFrvn85P
A3z13XobRhpl/EvMW15O7mTYQ3iulPzxCmCgZzNWQn8CFeT8omuhE2QwflM3LkN3
feAVsgu1clTuPHMwzjziD0Z6A67lGgY+pk1JwBrkBGxNpaBjpZ8jLZZ/7+/SM6PV
2ZGDZLSUJ7bNsBmJmOorr1pNrVYd9RbZ7IeRd9gW5rNmJX2u3mhsU7USRX8zhvn2
UfBkL7vHKBM89pQaZdFv34G4lvXUQnk6VBrxXFyynuW/eDyjUTSh9zMzLYhpC5e0
lrvjpf+3HTkcp2S477A5tsRJsp37HX4hTQy7S9ID7ut1ToBC8JHj9NfsmLBSXuBF
kmPdM1EYcI9DitBh3ahSf5Eeo/FwX5jsqNKOYJXrzy4qbR/5mPZYAw9ytRS/aEd9
53B/Rd6BMrrpiLkVtyD3hPdOHs9oDs0TETPHSqbZ8UMoK2QsybnMmpx3zoYm//mi
YGGK7q3w+TktKFv349fnGSRG00eF1wW5ktLk+9Gir7BSmOenq3WvWVogOXoP3wC1
GHDXGT9ah1FTksuXlIOdVKo9AaxeVY7wW92avB98b2Wn7FIM+lc84wxoyvZJiy+F
iD9VB6wM0CDPQgUoAfdDOnGzLncKiRBY1cNBggk5yMdFW6WK1tLNsh7a1zXpw2Yw
zrTMJxyYMI56CjcsXBrE8S2YXSiamHXjikiwElxZmYjWg3dsZMA2itS90b3B08TB
SNiOihkUCaKL+iK5D3UrWiuRyR3oP80DQwzOrbFgLnY5eYkfgOZhToXX9qUqWhGv
3vW4m5LbcY+zg2nMo/zHcHTx6T5O/SMwNOKsNvkpKr7uWhl6moXakdfNl3K+arHI
8dMxrsKHHwMU3PxfFWDX+Tj1wtAmg/brevv1bx6V1OQYdgZ02onpuEW+B2dxQydJ
+dHhwQIWv8Qp/dby+dr805QD4/mB4hFPX+/WQfC9+kQ37r8d899NC8rs22N+YEip
9Vcn5iqym4IgOftX1A6WY+EoCq0O0u5Uj/gObyD62OPhWWVPQDMDRsfsVYd8LqQs
hIHdbAmqsQDdMu7vVnzS5iebmuABpaHn+AuPlrhcAIy8OvB20SovvI/qA+H42RdG
QjUKchdNaUEA1FYu7DtKkR9RRmu/JfcC+rvqQkMPjhQX7LpDufZ/Vgtp8U6FZ/Sf
1SDQ5vlrOOu5T6aBx28Gggg0slMOVmEbD55eyQsKcW8Sg9TzpFVFj5M258PLj5iQ
OCbL4C9SEgIJz61KDOgKt7TPwV2YqniJD/JJK8PHtwL/u07F76EK4yodQriIfw+Y
Z2oMWhPLDQbOnEFgYIFpe/Qf7o1ExZ0ZhNhfYFlqmBqClj+Xqli8ej1K9FhE6kAs
e+lJlRXui+tr1+ZkkPy074XgMzEyRLxvxJOKcipoPNq+aJ8lSYKtsNxH0Qff+xxD
bxRjuwO9Fjy7Z4qIoI4dBEa6MxwtwTW88N3n151Elo3hX0I9ZnZ7NGRSi4McQFsK
NtR0tm32zS2o8KK4M/74k2Jz9ZTmvWdMpbtKjKM4usBc/eLB8E++Xqvm7cyYmPT2
upuRsbgyLZRicca40fdVBiQrIG7ikc6pekVs0QuxW/WbFA5wfEUJym50deszkW/m
1gTdLSzmGYO/BxA80RIHM0QPPlUzS+30A9DZaR07jdFmMsKnhO60AtyL6V89oS9l
eBUUFp5wcDqKyGfr0wxRYZp14oK3EEF+3Syk9qIgnwSEy/w4GJvUTNQ1q1NCzTU4
2tw25Fgy9hAFTlJctb5GgVS0CM4wx4CssVUYrAXTXBtr6NAAqZlvbqaqrdAMlXsU
0CAgU5Q9rqY0YoWesvVa1jWUOjq+cQ/0yG+LECa4kbkFWnfkJbr+Cv4bQfcuVW9T
W636F0OjIRMhqdSea9VoFBnfIxkaKxqjFzlBsZuR32y/QOcNkuFJ6csv3N1AIDqL
mTKggShRvG0VmG4UIi5cgD0ZWPCk2CXFV1+d6mbgbzT/0fJxszvbaQeI1jbSudBJ
hGpPoxgXaHtf3bs3/SY9bQJxwGsC8ziJMlnxCbLc43uQkgkwIIAweEMCkN6OjbSp
7sRtrnDWtVNUbBVWwgQ3wamzgaGIOTbXdrYqU+gw+dagr1wOI8mU/XlFbD66z4Xf
sq6Tm0QW3MZisK9pU5EtlxdvpecvgW7f/a/dWafg3NYOfEk+v0+Uei0tMZQ8LFqP
0rzaI21gSfzfpYjTE8MlCZftkb7k0pOW/gBcTd/jVGpnSK3QqSMKyWCIvn5iHXdR
Fpg2WR4Io3nSMj9+A832Vkb8CqH9GDfZ6735nXgnRW2fdQ/mKBwI/TwW8CO8k65H
ffBfnZLN3PPfHKdn/G1KrhpEmr5+VcXejXJml9YcKNedvlew2gWJpvcaexqXcHTz
N/bDsuZBqDA2J1sTajaXfhc4LaXKkFrPdW/yLOO3EpXkVsGMgxh3277E5lRxol3V
qc4lBx/yV+fs7RzkBQ5n9aViDuqfwqekvb0UwUd7Yy74Wk6bJF4GHRQ+PqWhNJad
AqExNHakLgLisGAuXHC9XnAfR4U2qHPg0tQPb2UPGUY99CQEOJ54GxgqE+SFs9Q5
lrUcCJD1xSlWvO7QR2FLIx1D5oqoiN3VxkJVPw1H7FNILzVCC4TR+nzzKfytAsBY
l37v1hsOgoP/f6CUjmwsd1uyvIS5DyBUoQpcldkBR05qcM7dBcd6kRMM65mwYL6y
YTD4CqwsnAy0TOczd5MQ5kso9yBnzlpyad0lyDy5uVgafDtrgBn6IcsWaTdhbGa3
MrjF5O3pgFAb6x5deaJ2wDY+9KF3ATd/e8ZSDdC3HXsJvmqNMb9Iq20IVERpa8Yb
og61r58zohv1dwyyf9IEuVjUpApB/y8W6oei/6hPpMsFCrEkC4tYl21JrXj6ljhK
5Jhb2AM96De0LsWwvg6nAFyQbCVTnaM1p+MCEImVR7EyqVfgqyS1g4ka92Y8Woro
QI/7UZR5bi2r51coYk2z4R4YrYkgA66/km+uJuuDDwxx3kToPphYUSVWvFb/bpex
0/CNI9Qr9abroyaisKdWqlSFuHkjBv8dhL7rHkSxqN/GU0M8golcyprfSlkxHjRO
qxRpqy+2XGe1K2No1mHSeXA5M/gO7P3An40ZizBWvAl3MKtPlYmwDJ0ASHtCUf97
aFKMYu+F3BCVihfp6Mwd5Bau+mjCCClkDvG8E0hCxmKSz8oQudBtRE1gAPhMqa8F
CZPkHKz9/DKO3GcGT7RQQXY0U2X9ck9Yn8qSuadBFo1c10TaSpTKC42J4y49IGfm
WTBGkvLzSrUnAs3Hm9hdf6XknJyQE5WF3TljgXtHOnBllJRByak69n9gppZ5t2f2
JMbDtukts8cTkVTxeRm0zjquNtYFH1Xi8SoRaZVOGyVqgSunhpEcooGuLvFxl6VM
TyNe5+jZIgBgMSwDGoKydaq1AeqfNZqzMGZqG7lrFkOMJ4MxVTKO7xeXbq1+sGGU
SmeT879f0AiriuXAXE0RweSGt6TlFu3VkHeL6yDP71iT2UgWP89mwLCoMclsIyxq
tVHJwqoagRoc+f3/51bP5Yo9JQdi6UO9n50ppbomYYG7xxXj9t5SnbXDMtWDUOES
wACTF8aXlGKaTnZ3lpRIHibaURKYb3Rp+SZcra6R6bOGwqYTiCdUc6TsZiQETJTx
9lbx+ITb4QAzCzpns1BvZoN8mcDUBvk1fSmhnx1dMo5bext+oXhbqm68RqsC4sKD
VAuSShEyGx0h+3fJCRh24N7PceMcsPpKlr7hClHPuJp3DAFxohK4o6m6jd5m1oNC
ZVpDWTZ8jzk5ML97srH0d62WdZMnHrM8ETXwhH4ZQACIgTPfUx6w5x3EpPv9bgVi
YP1ZlKI8H7odoNXC54t6chH8/XL+xK3N8D5Cgypm7pmwGHV0PV7tQfyU3ih2uygV
0JhqNdYNXL4N5UnCPHZ6fxRdwP2s/lEEAIk/+2ezrJJBcTlTHRHZjEPyhQbcAo/B
VkNHuGb5uMcD4ZmLiS+OqILtU43s/jmTgSkmf5AxECNKo1m2ESgz+x+gU4Y1FiM2
qd5vMaxdShv3jQmwOPJXSB0vT9NUdURpOjpcFhGbLDw9+SJWXFr8WTlVt1Htf7AP
GF3DTFJZnOjB7J5xCfSd8AoJRSHFmZhjm8MIUm044PnSLFBsPXIXfoiEXwRy0Qc9
wyHe/wkW2f8fFP3pV4ZWx+Jp+7yM+AVjFia514jcUU84e3bvJXiLADzYvcXbM1Dl
jwIU5hhOh97aQ5EZeed9GzMdXO07E0UjhHvhXtXinfKWppqWVLG0TrNf9fHPnD6Y
g1QFxnW6hjCYPPIVo9tV/FZmhj3AujTOHELS7i8Phf+dqAs48Gwam5z6mz3paAKa
ylvr+Tfs59/ajy37tQuD1zfVHWRvRF1pwN1rMsApT9wltRtZ7F5ayFzXdkC4y+Oz
WwVwfmHUUQXhalwzAaql+4Y01v+CljVb49nCrKCk5zjGpLYPWePNnc6mXAVp7esS
pgye1DVQf8WPbVk66eHC3T0XTmVlz0mT5js3/TgJpKFqBNsaJUt7X6WXRkPBsRAC
nsGSfC2NE87cyrkbTFAdu9Qe1Q/1e0NCsMVhovg9QPUqn219hzPC45/504I3DNdH
Nzyj0e46lEFji8LDefNkD0HqHen5Zlwbek6PcRat52mmmhuw5LvGCjwLJ8/j+58c
iWoxw0tWjiG6ry5FBSXJ2CPYS/gzHAn7NiGKon5JSmVBi+KcmVsglhP57cauWp7y
H5sMRlMWl5WUiXDm9dFuq0nkNh6F2fUhUat6IyF5NcmsG543EWMZsUH9djHnP1Oz
EpvKK2nq1GVhJ2s44yRAAa1hWzfm6Vik/pfhj6S+6fUNh8PCaRxWC1Pbo0JM+g5X
SB9758wOEqSHt92L8I370bamDKXrFE1GpX5/9nsMyo0w+8Ga80b0wtyQAvPJ/q99
fURzj6iBXGAZFbycByhWULvMJYgFLtt5rRpuSh1my5tx6vY5FkaJr1PQd4ekPxF7
+3jTCawqRLf/kTo3/cpK0o4eENW5zDli/KGVyOoJHrTQuMzkXfvD3z4RvuriHJpe
j/vCZQsCoZH0qlTcLBDVXQUBxgwtgiPqF8aXCd2pOztrUdE4wbXcdL213IfUkt94
dIEsI0W/yXEr173tZ5FC7BtvG9u7zv4CH3s7SdWcAEPEZAb0H5seXgIJZioUWwsj
g4IPMb0qszvGMpvNmeg2FEW8gWvb3a4rSxTJskmGW48DD0bF6ax1px9EAI3hQNmo
WQUgMmY285gJRSeZQFxNBD1jYoUtLWsB4ISoyC/DhwttuKfUEFsqej+H3IzIrDUO
FUQoHoIdvG7legkMJFapd/wW9btbcvyBc7zPco6FfbX9ved5ULrMUJtTX9heyQg3
IY82ZJplCc3SAWXrUiL8VDf47GhF8qcflwaUNgHVr25EZV8QO/RYNrjTMry3uEV9
LmlntKH6G4uNxFljYLz1aJFvmkbY8OpZm90d/NPdMSX/ovaPxRSoQOVH6z5hrluX
P4LGGya0kdgYH9HmHpVzGGSXjHGMLI4EykwAHe5O90TktkcfUFJvk1TXeqVfZbE9
g2vjDjhb9eer4NTlcqo+1+mFPrwxOTGHULd3L9aZOBuX7siRitSQsUAlz1vePnAX
IPZGOaTL+6TVsbjlvJD3K3VwvK0Qbc1bkE3X/Rvd4JP90luYUFWAAONAapbCkiaM
FJuNu+y8k585Jki60lYKDr3Rt9SlYt0CRbGhjtTH2qlCQod8KflsRtAtPj36aS7K
ObAx01FzYHY/Sfn7L8gEqUlK+hMcBmjDeZvbA5yqmz9+HCBKsPqkv8OEGK746pBP
rKm6JIvIgqQKs69fBGSZjqfDb+xDJh5sWlmHYaia5a9vEkqZqfndvNTlYIKVEs3r
yx/Fl+etSX8nYDZra+jbR5Q5Oh1sabKDHw1VwCyfSP/FFgZ4Um8LqZxc161RF4Uo
mPwfRa7zedlUV2brqpwuo+Ds/+kIHQPp9aehxirbInb4jn+2CtS4CYrWrn3CLZuP
ujO3vWg7J3m+liL7mrnd4Mjo+JMXrtHlpTI2kL3QGJqX2nr7V7fQcWzA2uadK+PP
ysa0kODeNvvE5FpLJEHTD9TQUi3hF8t4ZpLsBHves31Z5hEWbIEZOkUXjckcLJRF
/Dkj6Yvi/sNBFKU9SXUaGe3xBKCImhiOCU1wBi9b3vnnvb7HCM/WGQzOgFzjNXHo
U0+NGhVH5xQuO8qKiNdSx9hkTnS+DJTn1etrQqpLimVe3YzHl3gxg/NWvo3nRjcJ
o8+gR/duqIH+bPZQoLnHhGQcExWjqmgm2lPE+Fbt2tWugbo1ZGlWhqmFZmyDRtPW
rWV6hOW4NxAewyCTb6J0+IaMSonkfUQzb8Pp1WES6FtLW7XCQY/T2lHiZFcWACk+
73G5e+l2PLii5m3ZsCFi48bJ6nFr7cxO+ynR+KqAeAQTEaHPoSXXo1iTREhpJN1j
uBWLgfkaLS+J6TlS+L0lCOZdRi7QfJEMiorJxemwqSmq357wzZCXyqo7uMdIkuVB
T8gmmCP4HYv5iq816HpKnLssYkibqnmPvpa2xU+O7WJHOSiggSKiWxLKVNJVx9m1
Z98joIg2naZfTvIiuAUjgY23umOSHl1z+Wyp8flHwvGJZTu3KB9S9FlAT+EjgHkM
lUMqpZJKj+CWS39+E5PqvclL7CSfMbEuA91R+efv5Ksl1Jcad/IqcBhdm3oaY/8c
iAszIWQZ0B/MzyW0hoGwaXkfsJBEcsqruf8fyUvtcpLky2HMKnTQZZcoCWFpKJ/4
ZmDe9kE4G5P8t32FslZNG7NHIJ1pr8vz2ShI2xjq/uNVBbCFlrS2kFCPAGc0i/M3
Ydol/KqHIphggc6bNaWmudhPh56FDfcdCoernOguk54tVLEsTPSWg9CXBeMKpa9y
BIDMA58aLrqFDUQ1OXiyBYaS8O4D6LvYktHdh8Hpw46DBrBVinnDoeu8/hQLmcYl
wwA6vXr+RHCLm/ruh11EzxnTuVBjBD2SZoyb3y9bbxoGLr7plwyfLr0feRja1e/R
hr3GVOaLpJOcHfq5PyBrdQqL6mmp0D0+VsIBlF+/xRYVj3kl25KQAKqq6uLsHQiH
k95Flbhh9YLCyzey4XOywV5IHAnDbROORX/D7XMueKzeUmohadJ6X88zrL6NWIUe
PUdSkjZbyyu+3UtHlUUHiBvbrYonRjSaWEh3HoA4RxqDboJMo+P8C/IWxxCnHN9C
0SaUnZ6LX2BMvEhuI9RRFjKONNv646hLAl1VwLdpnMTWW9/V3rhPs68l3DWaa7i0
MHISPgYFNln0z+UjM+Ev8tjbv2Ga8p5NV4e1mPkKRoCdhnTDzAZzJ0Ol06pGlLyb
ok9IMFa1VhlbusVs6BUOUBgXlHXHUSqL+qEG7aCayG+poraPVc26cNput/938RVr
JyXqSRnsNZYEk15LFrrzr35P5nFwA/lN4bZX4o9+wbF4FNmHeLRiOpBsutEhoJFG
mjjn658JGxbkmcfjWyto6bP38ZzqWOmfD2RyRiPA3tHXM9aoQzYdl97pz9AUlHlf
pJrOnhrHlqHUhME4Yqmj7NaUcZrcr6ZSUjVXs/diwhtpvb3kPHBcbLZ+LdGrHkMV
TXuCBUFDqhDdUu6dVHG95cNl5XRWmsA9FM9EH9bbcqoFZ1aybjR3ZcThGOvb5Clc
rzujIV0cnrHPQh8CnyKm1jmNpfOSUz6x5l7m0iHuH52gCdqidhfKQQvlMWyuE1AA
0CEMoWpmBBwI+H6Q1oZOtEG3tULZibmP8V/AalWt9k438KuXINhABd3xOWRyAOw2
4FCnvOlL49UmUf2xepuEocrhDGhXO6+kMslXCmdvA1dPKLbCeya7X7WMLcorQMZ5
IYW4gqy/AdUADdFeUYPecL8yrMnQ7Matj9iY1s4iHizBDRGJbi+8tc4PbEzHQ9QX
n8pQfW9pDOk2HpSHtQbHeKtbIZR7rNd5CvcrwrHn9a4z1pguS/g2JrdmevLFbZVR
qwWzYCQ18Nh/1M2nHPE9SOu2h84MfNxqnoYvaDSBDldQvd3e06HTgJdmZ1Atkvkc
d/6rDhty8QPAkccKWyobxNJ5SHiEkiXuD7eQlIZpjJA9E09ONueNiHj9z3cp+Iqd
attn1jnxBvdreNbrwNp8WmHu8VKWYMJTUzhCtpJ/XgHGPAhPCh0LE6w2xCJtUOdm
ylGPXThZOS3stGQ1cwxPonE1yCJSAcEz1B8IYJcbTIkvRhCgw3BiKXzY8SA1O6DE
pcgIT6q+Id0wnx1YSjmwMBtxSM1gOEsvaYr/Q8HpbN3FPFIlWqFe+H0Pj0N3Q7wA
ABHOW4JAhrXcFJeUimONsKfRoBEUsUclsXIYqao/u0fD/TP7C4yc2zw+d6hWBsRY
EZCQSq2tWrJ2CjbrE9G+KEKobrnoGPiCVsiPNBAg8SgE7KtxAzpXhv6/tV/BoLWt
MLY2wPLBlGOc6Qhsg6p37zvtIJgNJ5cTSk/7Qh9j4EbIQgTVB1GNWTLTbIZ+vv1j
/5En5a5lIFXRPE3LZOrz6yHqv/+udS43lTs62rKEiayzqGjcFEL5Woj+OMUmr8o4
eulTPKETiO8/L8kwgyo8X544bKcFtjtTCOcpiEpPrkH48ybzzCpIMFmTjtcYt3p5
SfW3jI1GxGgVuGQMRY0xmtw8Zn8MYFjywmHp7cG4698TfMkVd5KPx2U2kEHMiRsg
2hYrVn3bjGtuanP6DDxov6odckOA63v0poZJK2W54HaxGN95QEKfq/tbXS5+AqVU
X25d1vOdZUA8SlnIWbUckNlfKsORln9KQ8TvxOtrK4WpEnEORpiqVX0hwBwzmlkL
B56wa2C1IjJveCB3PU9UcOs1BW9DO8S68t+xwQCovzezYGFv3Kmiuu3Uqa0lJgKk
q/GpFSVlu5zhrLryJi/ad1BVltTeY/qUyLIbOxPsTa1eCHF3V9XT0eo2sm4owSLV
rdCqbGsYcz04znnpMvy6Kk7xUNamGaSXezfJmbJc8litnyln8NDqJ/4GASIddeLN
hX9MM46Py1sa7Gn4LlyWqYTiGdyW7qjSOa5ZZBJJ6mKyJIY58rKVjwQhxk5XKtvX
mFX3bBMVoDZlBT7Q5qDBn1pegpJELEjFVzVeiPxVtZp0dtjVd/FwyJwOo5d69J0l
bCbifcF+jbqctbc9ajQCxX4bf34DoeoXuf+L0WP5d/WCGHbO7r5cCStfOJ4VGIB0
NShe5PYvAgmYbIVvurjrBplUQXlGsuT+QjBAFclSBVZB9dFW1aqd8exABTp95mhS
HyeRmeG+mlpHRriNlaGXw+sD1jWVrI76hEPwNnCnP0hVhcp6HrGYnAl4HH070EVX
4mS/709IriRFaqAhn+ZkCAMN1BycwrNBeR1qCUmYj9BiacnhdYFoe/dcXifmHHE7
P9gp9azbLiLXRKbvJqtsn01oWGqYmn7kIptfyBSYI3YE3bNrb03uxZvQ5bROamsn
Mm6/6mw8zHkomeqouqxzdYv1V1AHq67DxVtyohDIP5keLgfbBSL8+zbjlqyOgTJG
w/Q1pSRFUTVLrgRJxSOQip2lXZsWBsQ7Sc8lqD+HHN2m50xsjtI7yzrejLty9JeL
SqGwif8alVlNhAE1z4QYk4mQY/cm++LRSB9MwZV2ZMm9gzBVvPyjV153JQ9jBUGf
ekwSjqGn7TFSvh17Ojtu0jG8JXGyCPSKCU04Rl88gEbjRoCrAfv8ru782xiipj6t
v7+rmQAVKysZpE+yACalwOm2YHQ+GFTxI2Z5DN8Qp9z0S7ABPiZ8WDEVJmfriqsE
mIZOXjZAHCnSZf8RFBKFXeZO/cLis3BKgcFBUZMC5wd8ST+U1lf8K0SopevnQd1W
ZMN3MGmVSf/FMLawUN30n6ivUEP1Xp/Cc8LAb9lS523cWFvjVAGcPMJ/1iYvueO5
VwMlQq/axGvmm/Pevulf2C2f27KxPHggSbnmwoWhC07MvlbI5AtA94eN864KWv8k
36ZhNm00qumddDUFCr7EDm9vynY5OQ7NskxSKWb+ufttpMdyOjMacEGULCp0Jf9X
aYcf1WeO/s1OzyZFbntVhQTwwC1EfXAMETjTbk5mdNbMoHoYaAssEOigQD6Ab/Qb
xPLGWQlg6XEWgpQmC822HPWJ3lFFbggPbCViUT0koX0/tLh/zT598Utjpwl2exuj
ZMRKPanvkBpZViW2tSaid4lHnNcKSIHTxA/ZmwahZMbAWlVhIZ5QJrxRUhM3FC+D
34gj1+jrBHBcM+x4YmBajo+eqPqQ1spooLwOanGDBTBhmNY7p80xqa4+qdfEYwsF
VgFsIcuLWA3ARJs6iowcHS6VB/6Ru+ANoFqt0YVgHwBBre5aAwI6XFB3XuyQ4kGX
tT7Ihw7K6z1TXbCYImEudZ9nCZCHqhKYwxJt8j/ylYlBiQF3nzJHYcdc5E68wFBI
fQBre/ZBSIx7KoMPJO9xstaKuapvmjXgGShA/gZIQ6dcMqv8KJ6gNmRiwJyFoyxj
9nct2QcVrX/XFfOUI22ULgNR+A7Hsc/HSueLS5aEWis0SJbqKK4j1dLN/e3SVlSl
eP91q5UpFoZSlYfNgYRxb8dLT1xTRGN/d3nG/Vq8m6pp0c4QHmJwdc3i38aG8PYP
qG8vR8ZFHp9ipJ8BNHJzJl2FxFpnzcM+DoMMuggmKMGpVd8W51gD/NtAvebK0xvx
jVWSQQvHXBXOkXbD8b+q+cXUKQNUewImTH+tzcNKxr2l6QXq0HA6hHZbJXZ7Ao/3
sheSSQfb1sxjHn8/zchfSAo3LB0SeMLbWVBsMQsuX6jQN10GwpCRNs5UGY4ugAmi
aU2ZIQnC5r5wgsSHpn5IiMt8Z8ifXMx6F6/WjGNrGdnhxYal96CqmBPfQ9d+z1g0
82HVzp8K0JCdiEs2m24cLc69AYOxv9XMp5psieS+ObfPhOe+MDQpxNvv2g7UqpNc
P4SOFR62wW+mcc+iCA42V2yOwU8TXtEffiUl7oqzBQQwUxHYu4rbUtv+UrPDHY3f
/PCdItGvqK9XkFDi3LWT/kw3f9MwFSbr8YA9F8dw3pF08JOWOwAzGCWRQ4Z4f0qi
H9TowC761ZwCEUkMV4lUyJgAkdvx1ZaUXuTWcSJx0CILCXv4n5vrwa0CgkyECrpG
AFfHn3alZi8QlGO+FChIU3ECeXqLCwUwTvC66+Tay5CtEo262gZu01Wi91LtniTh
EVxPTZTO3Gqke/fk5NQO1MeLDOKNPKoQmF2JnLLLxO/yLE/vxWpC1JubZjjbERso
hQrM73iraYMoTQuFNHX7lubttY8971HOpVAj6KWoJ8s7APpBB7dRMCcJd5eEBCDJ
0lss9B+zwHIpFBV9M9Ov/Ft33VMXB096HSHXMrT5D+bTkhUdHLCEnNvqFSeJG+Yq
lceovBcilzeoLAotKfEOigBN7dPvEyUZFlDymvDt9FiZoQxMQCxO9Qa5N3P/P8zq
8Z9rr0IaBX3Tqg394Ov5PjeOKD8IjRVZZuVofU3qfCOaVLHPfcVEakUQr7F6mxDK
Eqq3Tx4oJ1pKT5V5a2VSCdtT60HL+//GcJrH+mNLSnoLexy5TtPtV2oSJ5J4pyFG
a6XsMa6ob4klBWnTo05xhcF0+UsWbd1xqpH/b5cFIe+j/dLg36Jatnai7v2jF03w
BlRIDDGcADUUUuZz4H78XJ3A7hBas9uq0pVkWU1+R6MjCiLwmOCYQJgaHi1KAL2d
o7WIINL1YuXNc1Wl4U5Vn9fzheGBbIcVXWaKd+oiJP20Ua8NGJmGF/VI74gFodxG
tangtXi5b3kp3y7N7BD1AdVbwIWlbWrQ6pvjIdozcp3ChjQL0pt03naviG1wnVdg
x9x+jHdegOKPHHMZ1KL3Ate46S8CppyNQRJaSZXTTpHztfo4uTkSIMai5jw1wPZ+
Gff3+MYT2q0E0qCr2V41T+pNiWAGgK1XhuNfCzhYrYcudC+fyVLLGV6MakwBieUt
4IdEJ//bHVcV96LGizfwILdwIThDSsYp7YIS6SV4oiqwYiCCq4kigFlippvGsHcT
/cXzoEprIa6wPuhKub/NY59b668shBLRHP837N4v2jgWysjomupBCaVaHUkNV7oJ
cuuUzXOYHrEw+61ic4bP2ws/mpU9ESX3lg/Hwcf4IsTt7mkQsBpy2ONpznALInMB
FusiLa5lLxPMoFvmY6VjCV6EhpVBxur8VvOpi32uA4ZbGgA06JsIGGA0rQNIDHIK
/qoS0vlV7ODcJZhcfa/KNDEUWSQx0ONJ/ioR6tnZnwbECByVBDm44wuD7Sf5TD5x
Ipuut4pDh6VuVI/wkZt1NYWZYSmYVr0aKWngsCFHksISBPUGWs8GcKd2r+F/Hzaq
CliFzNTMl8+IcD8aK2oJFqi6mBphCnFuk7nwpUiTCf9H32hUTgOmNq12KsaCVqv6
iNEATA71K2wiwplzBAeDZUAHzuZiSMEojUc/1BogxduDBuNwtpb6AJMGLNLOgk1E
H2/LxYElHww2HTyUwAXecGX6AlFwXlpI4HA/BMhsjM7s2M8RmKNjy20eoNyxLPGo
A+nVz7LKdrbdpNJcIcbwmkPIARLPxYMNEm1op+O31fzEPRU1Ru5fzngVyy2HfYgV
gRMIoi9tlNLKDwNP47oh+hccofQ5fEekVo6kCIC05qKl66fYJEgVqNelBSWP9bhA
xMYzvEBUnrDWiFGDTYB8fJwVuUaGQVbOYZckuqcRgRHg68x2kTy0neon6eHbJzh+
Po+HIgYKEUcnazH99/iAZFHsPMm6JzaVvXJsI4w/3zuX4v6DbHCkCMSxhYf5++N5
ZPGHL8Mx6o1MRNwoBF1BdCTVW1qqBFE8pHrqGEdSXm2lOnvsuVWvvE6vJt/llZTI
qjlzThF1Ji0etOxLvY6c3404CjE9JatHhsMkFXJ3wJIea3DhZESy0kXXvTxMWgR/
ILSr8RmfotDulbEpo0zuijkx96Ng0Jog91vAYOQ5jjzkqSqCIQcSUqLv286I6cqM
OU4IaMEY/qtcQxAoM/0wZw5w+kVsCpnUEZmSwKBRmuFtbEHlRHlqp8mxiijpyA/a
q/+JsKk81kmo+2bBGAtYdRZLvDNWRzRhlIF77YDElhFegwcx30OMg2Kj3YU+sg/m
gs9bDXum8y28rA2yyuiDw9g29/jUbJfuzh2I4jt0+OxAVqAV3slE1d10KskOg72/
+Ob9J3EQKGersn4e8jgoSKIfF447Zg1xiNwVyF4qQBNrTcCZLJF+RH9Lzvjzy1jD
GDf3TD2i8WAH6im5tsk7OnYm8OY4BHXZv/XjWswnRkHqjfkrEcVPR10+B/nTzrh5
MDiydrB8pSfPL5c03NEQDlAxABFGvHrENZRgDzRCRZjhYyRaIh8HFh66zQDu8Mvd
VCvOQBnMkLdkPAgCJm6gWrwbx0qzuZ0M914ueZWutIpb25hnZFaGjnbOZLo8Qrie
tk6oAsK+RAcpMKF42gJ/4ldpZUTLzt3o8hKVsO3/xCS+GlZdJ+6zq7CfojdnogmZ
I6S23qBg5AEPxwKkSLNLRKsTVN6IbyjvJrRanUYQZd16f+2/n9emWH6Y2n+mgFiL
M1DxIRvwwFERwzV8BArkfFm1DYJJdg60LnsKavLIhb2QGCDWxeIZ3F3mEHXRR8H/
Ic9jWUOjuAzueOGbd+g30yi07VY99YSRETcJWaIC0K/7SMjgD4gYg1gBp3jqN86s
Gvlzf6NskSvSgxDJkOfOXRX0FEHBIfclGOXqPLTurwMsKqjMzd8yYttSu2sR30p1
WUW6RB0/RdrIfd2yeJI2v4/umNjFTD6mebHVx7y4k/PRHgalHpkds3Kxjms46S2O
HlLviA+JNJeubxiXyRRzNZfdR3ewe+DO0yI0zpGTQgotAb+73OTPqlpsNmPw4ARL
InthxQ5qNjZipXhx7VAx5brX/3qDY5XIx4oksiZnInyxASGhzkgi2m9VM2evDyZl
AByE+hMOb7ywmXdCxEV1UxDYgfcCCIkJFchsk6fqfcHSp6lH/+3pk7s+uEGeTa9v
Ko2ebNCbbkMQZmKaPzrCuhpoMLKZzf5GvjNPEb9iTpMt8YycSGWrkRx4vZxVw3P4
hFZ2RSPaYkKi3g6ZLJ/WX6ABsKup+gvnF4ikOckN6gzykYXnvG7TjXwlc25UJyFt
boHNaY4p6a2nNJwbXkUdElZx0jphLoVAEfjgQWj9AAAtkCO2Hw3kD0rXRn3PRqyZ
XcpbGKS30plaO8AZ50HQGF06TdLsvs1o9mjPSo8WMPCWqtbAEr5r9Qu1Lgltm1Sw
+9ZUwn9kVFpJMz1T0hjuTi3XT+2oTymBtg/kiuch8yrTVD1/sNJFk7ulMmtFfyuO
cIGcQXNWfGlyDiW0QnK/eBHLtZ1VEwyzKzIoNTjYvTxPdconUAdogYPhhiKyZdpz
4p59HUVDlnfNE7/wicTqerFriJx2c+xOcrZqArr4B1PLPSC/QLQiz+dk0Yp3uH8P
RJWZRqZ36Mw9vKeZgmu28DPHgdLj/f4ejTmEixmaowkjmrBR3xBxG3IUc4TB5IFB
pz5z+483K1CMMatpMrXCIuGuPDrr9LGStmI39PZI2fqZko3iccjb22dBfGVAL1VT
QTRwZUgCESzqKeW/o/tzb3eP59LYKvKPSa+yxy7kAI7u/C8//gGwXN4eO8Oh0N2M
IJQ58ro4zZWDiRahCZPBVlQU7xa2ADzVj4i8l/K91Afnw/1m4GKcier8mq4e3j8W
w1MKdlNSw2dWLibGv8E0D86xqUQ5iizpDemzLYjinGa7qOgmFR/URZjEz12Lujwu
QT3yGzMsbnWYx0kCB/SVIqTmd/nokyUxvWDmKcP2A0NFz2tPWQNlqYw6UTVxf4U+
OIW0vOjSyTuNLhwfH1HnBM+blQyF/784hSFSGydbDh6M3fmDBaaVKSAFffl9+t+g
0+FP4o1jUtZ9VmEPKdaw46qOpFagAlgGl/Ez7ycE082Ix/HqGq5Al25RqtAElEVc
/LBRFbHPo9q1j0yLhXy9fYqF5AweRI9sg7aG5Q1YRwDxxUv2AFSWdwKXaXdGHL6p
yisZKMCe4z4dBi9wC2Nm5P9SI42/2T2NO+p4j+IftQC6f737mPfrmzFXDLVK9xzH
W6mvYODLSjpV8XzYbjdzbZTjI9dabHneFxAez8gbdTyMydCXaziWEk1iX1D+jujB
1pUCULl6AOtF2NbCM9CWM+JL80SkzvcmRYklpfpNxELkuxNnaaRYkM4i2qQsq68x
HJpxKTdko2rNXakYYI8SW4vZrh7negRZJqdSrgDvOyTAKz4VHvK1V/X/mZx/azEL
lJXy4t7ADX5B6v2BTeNcE4YbMvpO5WH5VXJGBxGb98NZDNsJmTVjzXmSJIEogVQJ
s29z6SG9Zx/BhsmkQsIyaITdU2ideaI0FwdkohpWxSbgTMy18ekPZo5Gk71cxs+F
y4ICnXj/HJIklEGIjEP7ArzbH8pHESe1h/ES/IPM6JBhpAmw6Rm/1xUvX2TYb2rB
/b4BinhCwAda9cZxvM5VTJe1azBLRRd9oMVTId4+NXPr0qHC6+ywAQvMWJdWq6ep
6rR0x3hCXUkM6tBZHLqkP9i/YE37t8iSiJAURLReV5Me6bEiDnU3z3tfmnKtoGmW
gXB5PtXHoytP5LPKyBgC09rTnJUtVnWCCsnA8O0/kQbfqmvYkPySaCBHViMc/LIL
OTggaJOh11jGJ3eHJUj+RAnRw0lVjRhW82gjmiHbot206RR8p38juUthIsXzIHar
jBYIP2YADZJ47mMnujcYzuaYEvdm+FvZQP/s2+9Z8ucShixBERMGDRTZH6ejC0Po
+0uCgQq/SOldaiLypjkzzmMnJtHroNTlnufGJO1Dv49g3eEdF16qAmTP+2xCLc54
E2j0kYKVNrzGFRILLU1sGXu6llv+mFGIOVsATz+tSdWnETc3KV6E6oXGKkHOWJxY
jW4mnJC2UMYwWdp+I6BE8w6UA0Od4/FTHPnNaC/zjgbvW2xaVp4NGOtp1N6BMiXi
HrS+VJq2ahT4R+5m2Z0T82+7z2szrwXNpzTZY4qd4LaOaAo/DFw5cEBpcCRj7kmY
yL2JMKsLnLW6DsOaba2IyPZPwnVkp5DYZboW5rzFAe0qV2LfQtgdzOdqfdYxa3de
XltLKf7ucpKlUznEwN5r3X6hu2G4V0x6WTyC6JYtUl47rxqfwrO5VNATCc4Py6lA
aDlCihLaTUrzKa9QxcCORttEOSs8oUk6OaH6Lqrx6v0nMeLTd283cpvXleav9pRd
Qqj4VjNfb6ZJ8XeOhstmMez1iKVBfrWgbxsTZzIS9Bif1vrgLHE/XKEjPrFj2t1J
M5encoOa09AfG+Cskbej72EGnIDgbk9BQchf+lWE/k7030LRRznimL3Z1Wml2bN1
p7FP8jY0O3rOReNXonOUjgLoV6v+lxd8zjaahyCOwkR5hINlb9g3eysSUTssV8kR
dIGUCn95TU0I+dW3kZWOkmlCb3UwEHcvo3XTxTgMeYs1YoeN9qXEJTMjgD78NYgQ
En2+EIwrFl6SO9lhoY4hYjSUkbIilV4ylDruWM0N6P2dMnaov/cx4suJr8oOxCNf
9ol3H9PDJu674zgIog+/tSdgxIaweFvVPltp4ZWT/8G0lq4IIx4/Oc4+kg79bvZN
mkAo5jXYhSChGfiL5no7mBPD2RG/EpW3kfEXOXmyEIUIxKsVAcuNKdzgM1201sTl
SM0FGWWbKVag/vH9nIMG/XH0ObarsU+hqtmmkD8xp88LCWaWwy1F9Z1McSP13UBR
ioGm8A6TJNXRhmx4ebGwfs1WezQKOsSNjIasx989Urbq2cNgjY+FcoDXheL+wLDa
oLRf8b3Xl2vw+m7/4FnegPPjNlfIyDH1LleSxY8E8lFf9mfWAIsIrxxuQA1W/AFh
0TclpZGiqBYILGF4HDQqAYKZv4S13iO9Cq6AuBKxACFJdUKiS//BXcT3gjEIPB8O
mtyVyvGTAgKP0sU/W5DE2gWfa69NmCTs+ZPE5BAqrTke0KXmZGQX3l5MhW/fjDZW
ypHhueGu02RkqVbv/qJhMURvftROLwBAx/lUoTf+ZBxEQPFLwdqDbkm8vMA335iW
Fv/D+xXdMYZw4TAe/RrEIsg6oj1eADx/ND7AYyHLZHNEcUVn4vpcPr0btTsKftmW
TIggaGPrpfP56xN7LYTxetZPJhOliLUShek/3jJs0bYn4pLpT3nYUYSRxc2a8IHK
Bq/MJCcdFhl+dA7g4dT6FQ4YLT+d0g/r3nzYrrro5VrYFlRvA3xEnFibKYglYt4Q
rYzXR7pyC94z4+wbAByQY3+gNkCias4b7laXnVW8uyW45ymREj0IErDza2C9Lvdl
113LL/Oy4TzvIJ22tpcAe7Ch/p6E8FLlvvLwSF4Xwsl9SBm0KzbYAioeAk7FhMMp
6tlU+D8DPwMUVmgtZCI5iai/V/ZcjHh7sBr/Z7iOUDGAW7+LjyHkpWhUezio1mKG
TJc6ear8njWYQNZ/aHqvcZEd4aVkBxL8ntRvdCxY3a8o+rDtWCK5BC1ZVvCHs6i2
hTs7v8FCRx8xAd3PNPF6WdLgMtHwJOXrjNOkgtDC+f4AV6YMGKd0zOKKgpzssmTI
epP7zXO92P8UT1E7zqMUNqaxtfGNjyncJ+sRg//XXdnUXXK9grTpdpjvurj41Z/e
BCZU0MHfDqXPHFbR3YXZqIEsiPaMnQTrkMznm6jMuyoQItBEBqO6QoFga5iyJuUH
lLWhTODzB2PgsNxMwDl3Hr0aC7xLH2+tQ86e6q9kCWTPPe+/xOFYXifB29J4wMlX
fg57nSVx8uA1wZk9d3mGpqQnnsZZ9NQfFNgkzH38gvy1TI2EK8zsmEtwCHnvb/4Q
yVwfxER1oenEitb2eSMvFx2USM5B1YF9XjTUANYrxVkaOmvWpO90G0ZYOSFOFZy3
okymvfVpa2ygT8GKU0406GLeuNVfD4U5fNHmrlOa7kBKlPdRh586KTBbMgUe3ADS
BxT+l69d6wai4aOWPHxi8YI/ez2z9Lo/p/1vlVBD71UDnK91oG/2retE0ouDcWOq
d7uxJOriugDv41eT9Z2rZ17WEfBRMUR5MSk9834ttp1W3GyXhAry3Ek+h2Z3o25i
BM5cGb9sJrCrOXYAcJI7u/cQ1t0UtQr3xrPy1ElqnhPKd5B3F6ZjzE+ywnZNWZQ9
aZIF7vm99N+iaCQASjqh7MxUr1Ubc7ajawBFXCB+yNroj4mPynmPj6nFQ0EULJaa
NZMh/obt/r+3WVXnQvdEQDf6gSiWtZeHMCZGJ32hBF9/jTPFY5u8Cnc5xR9gKxgQ
VYXECAF8EY+vgKegtWxmVgRvbtGZ9GekRl/PowLEIUD2WDP+1yWckFojdGCzXNPZ
M7cwgQTbcPKO8I7l0aNB0TMjmtAYozRq2WLeB0okEOfOtlwsnPB+jlpg16aNWpOQ
dmn4ezrsnc3/o8MZcrhbvh4XRcVSDiETDIwf0iW1jn3VyaLuwJQjmquI5DLRjfVg
ENJXX/V3aayLq6ROL2cN8XRPiaF8LI/nvSQ4hO8YAV6HGv5x019PEIqcJTp47H7I
1bPOqmFiK/CsNvfiPsoT/B1efZbpWEg+9kQMXruIpu5Xg0BmMWNpw6/CDCnJ+KTJ
Gyk47seM5wGAC+qgpwg5xU3I9LRetaRSrzDRYWu+2HqZyzJOY4NrdA/zU71+QGrC
fzq7/xEv+hvjzCZr4xhVcnVHFx8J1bGhode1YtlTsu/IXzmWQmSTz3zO0KxoSZnd
5a7T4LRbBZgtz6idB5N8GuNQb+R7ChYQ8bF/wO1278vlcrZdz2p+fZ77yYxP0XUP
WTH4eoVfBResOcX/Qy8U2o6N0keZ26GOa6qfF5s6fW7Joe21CZVuMTFsd2x0Anuq
Zl3iIMm5TetbQz6jHZPDbcxsSdXpOKBNGpHGb6XtALBp2zeIhHnpjYuXIJJFnHdj
lCt9gXi+WmvYP8iHHWtjeVAbqWwLbsUSGlzFalAijIlzI8Yb0GQ5ln2tzRQfLgyZ
BWNEg3D2MjiXXElECAL5dVddah69DhWTOzwxojlUVsf3cSQrBOonc44Ad12YJh41
5zwfm4nIwMUjjndSbS76jyNS5gW+rRI1SPSVmh2jaafwXv7Tw5Olr33J4xEd6IF1
Sz1FrUhdFePfNGtabWT4WHAtfQc6HCy9eeKyUWE2zvyavU8RnNC6epN62fOgJYMg
gLvrAYAeblCZrVx0vG2vIoJ12xnWdVdU6QNJZRNNlYVequlhUtttaFWawEOdAzJf
KP7K0eO86sZvux9ZHwKjysDuJqEZZQl8G3TEGg8JAaKDCXIR+n5XKTtgw5RkthfK
hTiiewmDdX03CH4JT1KDqLk9ySv5+GoP1b7w/j5w1qswRQTt+xLvwEQcVqTHUOED
VckF2TI6vt0sHE9S9sd4WirLXNzxJpP2c8yiR3st/q/SMlLlNNen6/ZIopq3OGwV
TIuMUlvswRNLF2HpCnWtEwHWa69j8zRJ8zkkSpsBZ0Epz7qZw2uezLBuBT8r5nUJ
t+IS2IcRE/rzrVQk2b+uJTlLkxPYrv/faRkX6czwtENH146BKFQC3Nj3O4/41156
U8F0JfW8OEaZIsPFVRhggL1CFCmy91l8GZCd84/m4wx84VemwD22bvvSxO+orqcE
CxOz8tvTIiRWdSVsRUQoZwzm6XPDPoEPfrMPxUiJJBYfxGOpAAe/r44AHh8qxkQo
DjlMCt2LYJgYe3slq35uVOgTjqioy9/ecgmvUtkB7nqEz3l7T1BdovXH9exzW3I2
YNPTVfzC8yMRvWkZ/V840VBLAPmeGtTjer5BMRKxcL/QYY10HSYBz1xJA04d2ULT
57w1NyHPBc1M7btGPtR9DhvV7/N4rgRJ5Dj3sgMxnLDqufoZL1knFNk3ayFq0VWD
6O36GnInAT+w2dLoOsG1xYuM4pNg6CGl4NLmeoEEwVN2HaxangkVNmFou61lN7mX
BmV62Q8cEko4hNgzviVZbBTuHu6e9yWgkMfsfw9KRI69VfhTSanBdywv39axAse0
OYWScba2G7nSfOjjaReqW720pmj/3YI4h/BKkwePc6rIRRW+M5T5K3SDnfArh6A2
A2wRtQA2apD8hA7U8JsiMEWw/9VX45jx5nnXN356n4reoC7AOESWatq4fO99OJyH
CEawpBBjDwsFow15pJRWIzX8NF4bYR94/Qa8A0wKE4ZXd4d19jZi/OM3MDIMlfrA
e1ur+JzAozFc2V60JMtu0M8siq+nglvtG8Ftem5YkbuM6naiNgOeTrkOQiQK2zzz
sZkyFCaOU2bJtLfu1akYpywcvcV0+XWCgUkODHkVKWGrWl3oEEGgl5ipF4+NLwqn
rZ5pPAHOp8YNxiinrUjxH7/465kGuX3sZOMHAMAVZn6QZKaMYxVPgyHe1s549Cwd
6PeunDzHJ9RpocumwJmiPdKaB/yIE1V1g6qH4DPNQENG3HGixxx0oIupNxP4Ppw7
h5kgskt+WrXQiSfcRVw41SCoLqVpeN1VMUPr3MWc6ahQlrs1anSe/f3kr3R9wWRz
gpmdxE3xpSvo+VwEpkOz7ZjN+1vqrZfVDm+/op9kozGuuBqMxwucIz4lOEgENluX
1Fo5t7PPrvxj8Nces14XC4OD2L7He3q9oOY9l5WHUvNkAJUQuMSdMHG2WxzpmaLU
9fJFmbGz9Tff0h97DamwzOzc/YNwss4LhQ0NfhSoKUEaKCIeHeudjkuN/0G/8YSQ
dsLfsa6fWhBmbVYs9FHk05ut+zznGaUGA2e4OrOsHr5nKy1JQWh6aFWIW26EinO8
Vx1w4+kYhVwtQR1Eef86Oj+MDqUFC3rGuX7KNJf1YYSqKIYsVADUI7eBsYmyB+WX
As3lmo608pKs54lzQBYvSYTSWCcHjmjyKyYRSvHVB/YVtdQptoEn42P7/YJec9f0
e5ImoIFx1Fwj+xZqkj7eYoQUUibgoiCMn0tTHLV5TXunL077k3OYfPvow4BuUbjR
3cJKNzkNPusDSs+fXXu9M7jHTN/6Q594LtupopOsNLX1fJaf599esdny/qVysojn
tWT/WdFmpQgmDkpEgYbO61r3FUR/EO1bX8YNcvtDSmHCyP1S2HXlYtgYXHdn8ylv
lKI91qsq5wYpBSUuVsHwCM02R6IIjRZTDzcihIOa7V9Qq4QqegHS4vYLVlIdMazM
aEB1c8EuM/5uCLEaCCF3MDF6eU4LUiIZEJpgC1Pvp0mimAUwF+rDHHn60GrxWKZ5
xRbhHppSUPoya7zKoCdh6NUeKeca1otDBBiijkaO7d5QKY8mhA2ha4D3yrHCD7vj
2exIUm6AeGH53JxoWTrE7SkQ7jZG3r580Wdn98a/7/fPutFgCTXOmhDIYZp1oHRg
OpZG7HAu/u5xPrMH4Mffb+GrItpgkQuV6X3zIAyc8QMlxfdeRLw58XbhGLgNZ3qF
zoLDYq3zR5NWJ46BtgeLKUXgwRqOopGdK0ruFgngZMyVyFqWX4dU6OtnlYkhJ33D
RSF/21o6nm/+fjAhbXpe4Q2q49WBifFhUpL6qb9k/7DUbziXriaV8paT8QN1ap5b
BQ19/4gmFJSGgZzaBZajycdx9+Dw0Ykrc9l3Vy6zwlQhAobMqVtvXGNDw7nF1cMI
bJBKeIJsj1RbaEyKoAKENX2SeiuT5i3028Sw5pwTNieLRMdeVj3K3rQQ/icotn/p
2azlrltIgcX+3UJbQsXaAROP9lgZFs1Ft1dqpHCfnuyF6mHME6Te14a+K3mLWX8X
TDMKyLG+LLEncZaViVLYVJ1eACj5vP5dDrJv0HJ0I44qqMCGiPqXJqcljcIE2q1p
zML6c4Ffq8CjyZWhWBq3tZNxVzRiQoJgeq1824c8rj292uAZAuOvrmDQcSMKk8VA
bYucdw0DzPdaqnXmN1/K28MJkIu8Fv17eIetqfPQ746e1+qDlOPkyIzzsTtSE4+W
R/Tw27M6dpZVSWExKVD6g+1VQwq8EQ453TLkMOyzmL1KqsH/OfWCLZJVaM6vRF+J
aCvxkrax6Eqpv5ak7RIfJ3kYWAjzx5s4hJtDaf/ylm2hLpOPUV6ni7QdxRlO5dGR
iHVpe6THNLr9QkIuH0e1NcDISUP6mrvHHN+8yyn2/veqpkSWTdPEDBVPaK0AsOlJ
V/wbGFfw7qAHxLy44mLjzyv0fgX9nANBSA0zt9ZPOef7n7RBBJL33+U689kcBER3
yMf30BJGgNXP+kU9zS503Nm6Jx9I8K1O10Y+s781KmT9bmQQJzbxtTY6uznGSr+R
sD83unXKvflvYWmjZrf9Tqwu2B/sUdSmwjGzXrWsrk3jZDMQY1cbnsd7vwHds2qn
bxoiaTBAAI19xOcze8T7fnwFFdo/30aRZwfG0frVo0WkKuRMZZPw1j5VdQrFapzr
cCliX02jCa50hCM9354efk8h1f8HTlveTUtWi/vPaLzw9AB+VbJHhg9J/4gDXVs8
VlMPWbMkAtbj2HvFpGkBGODlh3pLfFMuHk2Luosip5eEcjk2I8kJetMMfvi7ozMS
8A2zzsNnsOyLlK9yEmoCPnJ8YxWTw+0GrXdMDACaaRD3WHW17YKAgKIvPVN/Llo5
derztISl8ucaUJYQ3vGAxbTrYPCo4+bGgHI8OjAFPowExPm6LdI9d0N2L7/nwNQr
/PEbxrptl+Q3EWZR2gWOnI4dUJmUG7tfyStGR/odxT2xarEB7gfTmaxhjcn+7cdd
I7CkAbTtDH+ynrP+NA/rwGR6MVeLvfWh9xXZcyPq4qDy09q9SI1Nr+Vak5g9QDR8
epQeUFV1jWyFhPsqP3g7YpnZhtmFT3oj+VTifZEpMUv4uoCpF8VXfn6AKiVJE4/x
iCOc/+RXphtivqoBjJl7hhZD20ce+VPPz8V61rvUSRCRnpWbj51WhS5g92SWAnMs
TDM+7BZC0an6c7FdwKAQQTLbi2SCWcry3ZnAqhCvM8uBWRfB42Pt3w/LKZUgdZ1A
CFkAN6jcYKmv0pqtw0nWveD1U77QUr6Irrh/35l2HLeJ2grEtSpzKk2V589bwKgT
kFuHOFuLjTw4qS7dffcV3c5yCGGyGc3S1RRcptgqJiYkgM+dnH3rXuOcRjJOZZ4p
EfVuybE+V/sojt4GclQyBwIdxDclr6eVnxntm6hHrX8PrZIWiuvSQrDooYGQlhhe
mCqSkNC3RT6rBLgEQZGI071xScgAynTKHLr3h1l0Ppy8cM6x0gZRQ6NoJKb/o7Yv
UbNzZ98n+gOW/sEj53vnKKU/ZAy+vtfIn7x8rgqzx4+r52MauTaLzhaJXOP1VJZy
avMfSQlALMRboTzrUBbwn+QZhcguXNBSnLgLcdbNlpyREXmPUrJKX8yzsu77FLLB
gHK7BppCC1LENtziwYXtAvsPjjKM+FcSdu3/KXkZcT+CX3Rb2Bfk6oQ/QP6/iaG4
BdHi/pcI/FKUhuOFxnmDu5xDeOnWeoXkqxg/CMRqmuJYxwJE+WpYkP/l9EGzQJi9
tl6h/D+OHfVw+VUjdxJS6wqRmL7l+0UsDELENYnQuOPnVBQYw30Kq9KsK5h88l3u
AmqgBy+Js5lvOTukj/ylK4YvLWkU9i++E3cziPrhzSRKknxuiL8ObRGqjCnnL2iS
F1iFy53y/Z/yK8TVqORUUztLRXss+FfqG/Eqz8D3Q4JjyTuC7rFP2qlbtQGZ1rMz
lsLuDcL7o1op9+eb1g2B/z0NilSX2brFrN+JFYb6ImawrIviLl6/wt9RONhjOnJz
7V291TEmjOdltZLWZF95UfA5f2K3eWPYsCsps3xxXJuC5QOHrHFX1v7j8hFbwLOG
LUen0dcdB1tauq6oaQxQgx2B26jjlnVEdUr8ej6cK5d1HmDMT0Bb98oLUlr4jPuF
8KQnxhrXyZCj2u7fBvfDYAaRTnHFGm6wkffwiXWcOHmLpTTVhABNA6SEd4RTzpGm
WiHfjCYpDRIFRb9ph+Qs8wn4rtUer3x0Z6B5/WigDrMD2BK/UgMusmSIeDPkpCZ6
HoU9lPw6m7jRHE11Cn0+cZN/3QM5EmpZHVVU9w3GiVDmqAQNlC601DDigliv3o/s
HOJT9GgMcM5c8yVLwkJGhaWA4Xr7kulYVrxRsQDcBWfOBUAey4JzX8JRmQeAUlRz
z66gmx401XyI1F05dxPy3g1JgWAk2shGNkPccwUrFt6/pOoLmVUlwoSCF7j2FwXh
2nFugCGwxVm4K7nWDxaTVV21D8Aann/Ixaj+iGzjsdJQuZ+vtYMVyQKvoEcKSoMm
hI9iEBzkRGwR1T1KyvKRy1JntMOceqYYiXt7mGRfaEOmWe+3rw5m7H4IEB7/cdgO
+PUu3vZNLZ/clyg4nTGj4BCk5mHwclsXFNSJAHK8qBqwN7FrusAinshkUWm5hrah
tqfrVEH7WBu+ANYjaLMT8rwQLHp1ektQTx3sjZnloM7XsBJ4o+Ip/II3Z/IxkI+a
KPVmxJRLYCtUBZzGKkCN28DkM3nnAK/WrQxQJWJNXhA9a0A4vXR/Q2SRCq5FUuPP
yACrmd0mLg+WWTUzNkKXbus9wV9xAY7kSEyOyo6zTkNlVRKYjOckOBKN9TwF9nQn
OW4jRNQL3Rjbu4keXVNSLWwZyG++oVDYiykCj04n1OcJ9e6k+cspeTg0bMvv+Dyr
hRxfL8pTj/+nB9xxw4Bi0qQNb4ra+dmZjEOFagntnWB8QbQ1pYXmlTofnWsL2gfe
U6sLSwFWS1wMpaR9MPYwdvwSdXEMNBpBsSgDBdYHN9BpK77I5hIoxEq4Byj7/ZHp
u8sr55chmVZ5GGlX910JsLXTskkXelQMK53yeurlT72hJFH50IKPQwJLxY6gj2HV
ZlLyfIcU/ic5+EL7AK6t88KBnOQchMR6bRCf1Zlsbv+zZJD/eK0gb1q53Ksb4NQV
Lolf8CVgKWj3nbIyF3zJptpy7kCsWFcEjDljjuo94gFIJX80W4BaiRNftpf9DThX
Kb/ToB0L6YY2X1T2nsyEitT2IMAv9NElpRlkSP2U4Oj2jOH5rEslJlvfunlT2BRo
smndBHpK6Z8kk3yEE+MDOTfisbuFOsWtolQXrRHhAyM51jKWNHGc7OxH2QPUef39
tiOgXbAZYgGwtYQ0kSvk6QcH88im12QS4/RJd2cS0nFJ/S+vr6XzkR6pAf2smUnx
wgQYOHZmzYQn23Y2zSxcX/Pjatu8/CcRKf32DrwE6kUsdYyA1qbl1yedXYXtANbh
5PoJsVORq4aQbahA2JBcQCIwylANfvpwjz7lTVhIx53in0Ma3+FjUDG4CWAA0Vg7
fxFuncUy8UT1xiEfj917ItN+V6Y0K8oMooT6FAnR2xQeHHdR3fpqtZ7vVA22r8lP
LRF+CWButLjMLMoAAGwF1Cicdk92A+MGva9nQs2H4MMMhP3KMxc0EYlT/HJyt82x
o7eyDvN3BtyWV89G/iGcvvI+OsMb4dmB5I8lA5p2f+7MdJ8yhxqopkPeeZFU+aE+
jX/VgJPuXUQ4lrl93lNQ/iAPoSk+ekIMHN6+iIkhSUWEYdfiABDd9ZPYMCyfjogs
BHmWdv0ADhWVMtwuA42Pn/dgQZ3I6cQlmE2dx2XvPqyq9dqkTR9OSWURTXSb2Osk
7v7z0kz+EnWL5/yK8eWEYVOa7edR8gi9k+Gincur/a8gvPDAlMhkBZ0LrIQ4FFEg
MxMbOR0xOhnjKzaidvvTzlC5J0st6SkDXE3qpUVlUdMvmM4AGpKGjgfwVCUEbCLH
M+ksFW2Q8Rh3tMsgmTUB4x6T4NuoIt71x8tGK+QkDLXSKuwgRbVavjeBfpqa3CnV
/Gp/Euqvnlb2zQv0bTe88tv5J+u5QfgY1Xnh7kHcTmLzAmNu49AUqDiiCtwFmWsv
IW9JMp4slRi4+LhQA8jmS91nQChEnIJObHTzmQHGRk2OzbwNBVGXAqMyT4njI6pf
+B1J4+o7WjYvHlLBzrm2q36DHR8ZwQDPt+YbNEYOvRPyczAzAzN/tmG66Pj8rHpT
LwEdQNdlEpi35L2nvkH6YRNsB4j7zAQgc3z8c/0Ty9/ypY++/0jFXNDubQdRla/o
232kCHhfWrDvXXX4jti7BGZPNsP56t0o9+wLd+VEYWD1YreeOaKU4ea1MMQPueBX
9HfiYzoXLnE1L/l5hVRk6nL/NTzfDAJsoxGGHhxCX40kjYGYH+tIVT0+kC9FYsdF
oe1grExWZl76JviESlsUPOx4y4WxQ/bqVm2G/WGrTVeBcuV+UQda2sMtHmpOqHTH
DRGlHBwvlYIBUk8ML8GjIwXGLtY62RUN8StIm8zDDWDeciSgrQBcTnWFlNwSPqLL
/flWAkQ/3uSvXlA3R3QQSx9kYQXnWqOpfnCvY9GrI37siEXOs/wGdnRBSdZ6mQro
h0UP7t6079zJ655U6HdJ8LeSeXXpPvHZwNXQY4zMMHdxeTWkfu1gYePIwI9XI+R/
2bvRUK8VtLuq2ugWanUFXEw8eBzfvXyx4EnS5MgPvSaxJQRO9D1CWhVlJ9SN1niS
MnJdOO7LZyFN6KZ4lvXjW1HmrcZ/bBC8fgWllyJO0HeJw3l4Wb5Lmj3TePvMH6Rq
SkosWl0VZkpLH9+M+OASbJfXY+CzVXVWJ5kYyzMl6lXHQ1/P548NNUwfg+yIAN2M
vuPYZ4vM5Lpv6DBD+qx2o1hNSRxd9KjW1pnwVb2/L7GbhTjsMixQWggA+jZqWUWV
Q8jHQCnmaR2mCMzYrtvJXx5iM/GMKmGYy1lTIMXAToIHKxVgi7cZ2lB2fVNQsG2T
DboKH1ONCoagTjA/k3GiLSBqFZj/9zN7SeWhtoaqkvZGIoDYenYfy08TPfbOFOFO
x/8Ldk0m6xQSjloEQ+ZjvXoYpfyXPAEd6iJBw6yAWW25N1Cr2GO/t0fRSal1a1l7
FrkuFogg07sXjjOlIa0dJGR8iOqLq3kh4Ct/llwr9GqNiQWwubDtL9FyEuR/nAwr
C2Pk2wtbEo2H2o+NUTZc+1g6RgNOSicSdFf2Djqt6kx5hClvQFyMUmJORSsSahP6
zXi++4MKPT6lpja9nF0n8vYbkH+WFQEs4puX6/vJmluAT7TaFuipJKzmDM7ldtwp
odyb4YTTZmnmsFiAE2MR6s/+7HJZ7mDe7XE8dxkP5FqD6RxMTlW9B3RNLxI5Prvr
Sc5edxA+M8IJRoxaUhhwPxuyGac7t5EPAkH2QJAxZBGefToqvZBH6B8XQ/URHd6Q
GZMiW8MwdlHz5D1Jjm+7bCuS77IzsZX33a4qiFSDkbhRKOBv9hcXOG9XzuzVIkIh
wIAcBgOr9aTH6sUSlmbf8bl+ORn3ezonOxueFAYNvJOCmzJnj6R3ndSTRc74Nemb
0vx4FvWmVENtm48Cf6D7cvbHNgubfMjBH0pZOya1HeFApFAWqDe+O067D38waJ+0
DDlQparNCIJBZNQTt0zEgLcH97xrGFXqHpXOHGCwxILMfZagZkhXfW+l3nhdecr+
wUV/cF1/11alYrSfOkHmX2Mb1niV+nJz4Vr4fS5r+KG5VsT8X4N1U1AuDSgWy1BL
9xvGkQLdnLEqEzaeUq+5DSJM2k6TIJcPzzVnD6VI39YHFjCX5qzzrwv9fBQ+tPvl
bKBaepYj76RTI+fxjT44VaPJoSjVAKj6mXIAK6YPcT40bqxIolxl+k+c+A5YKflq
3J1wP5SegjZFvLMnOtAmMfUJqcnYTP6HdJJRtz4FcmTZEWMfckvWq6xoNpNFfiFo
tijJJVx2bteqCVj2ORWUSK5uxqvHsloEVYkrUNKbsuwyn5d9y86y7RKgcKj5yMD2
S0F2yLhC2sW3rkVEoUkYAtrHGougsBu2rLmT/a3X9dwqd6XvGCwQ4QO9bj41g4vU
QJQFP5qisaog83FldvviPzCOza8md7t4OF0n7NzQi6gsMGbjyNZMp6ICoR0z9eAR
ftbl5EqJoFVTJlxZyJMjtVW7Q3neaCegg4YrPWW0PxOkq+kXdEWUJqvaOguNxlXt
Nrv7Hu5k27Vd6qUvoi7wB5ciqlWXHvrKfo+OwK2tdjJVeFJTjDCrJfQceK95V0P4
pT2Oo8ZNOIHUgVkCza5VLWi5GhG8FBGAR889CofOeRz1rcCflrb4fgZ4xg6Y39UI
suGDsItVC+WR+ZO6HSPf5VPdO3JDeqU1pk+Fa5+3dyZsUuMf/8Rx1dZfvbF4rMLq
MdkVPFQHZP/lrQ5ytUOpMZj78h/oia8r461bOnZSyL86ddLC49BhnDqxfLwah+N3
MdzvLsSIY6vp2pNSndl4kBU9iuaJRQtDhgUjXAWrDfMnu4V6o/ehwQMG7/YQJzuO
reUiCd9EMQRdxCSIEeXyiufoDjow1lGoC7JjCS9sH7Q8qA0l3pGdGZ7dBKlA79hj
NWBaxbh2pOREHZfDMc4mKa3eIo5wT5qf55zPps/8XaeTake1WUkvSXUHv1hu+/hT
ax9KJ4PdN3tpnBqWNUom6FBSWDJSS7gz23ypf25ZxftDy0bCtadKHmrL5Pd/5G7W
9cN9Po2lj+0oebj+rBFwnQCjgy7IunERZtbsPX4dRiDFCgw3H/m29gxY1uq9tvYG
LPc8QJDmiMj62yqAjk6aG2vZC+Pq/jAK8rSrJSM5iklz77bqPStfxaCsYfZx+/96
FXvDb6gD1HF/vrrizojooZ309k5c+RS3VNFuDO92MrWxRhG6QpLN6GigU4L3Uvxw
1BmzwtX4XcQfdcS7sc4/gkZs7xDg6QDkcASRaZdwILv4l8P+DnSzhDAKo1kevtx0
9Ajk1Zkgh7k9GGCDF0+0T7qZvBCnUkYYjg86yLuklj/NPirhuz/nKqPN+/Q1qdsp
RI2t9hZ5U5IrdvPMknmp/XoygQs0QQ9nRC1N6ljZL8BD0rYL0ohRHCaqMHPp3yVA
M0Ek1f4R64ziA3PbvoAOJ6haea8TmJ0bWUL4v60FiJinjLGjAUMEM6MmsHlcZhuo
0E4x6q8Q6lKAPuM5JxHTF0hIU24BQgIE0pLYeTsrVzDWfTskCgS9hVrM3zdVFdXb
/aMNDx5hQHYOvIpnKyeSkwk9cqEsiJdTNWjDRy2+74qFHblWHVrmCyH0/Qe0zoUU
4Vt+SiB/FPCxtZCE9V2FHKRsqT30780XKLrDpmxJjFxeSGbuaAaC2MR+Q/eb1F76
+8awNUuVRRubcLi4DbhZS85V1xaWJCasVyLpj3DOwBLC5XTnJd09AnL4tpjo6ssR
hdKpINfJW8YLU06YPoUrkzaFhrHUEkYy6NUDSucRl2+akI2rkgF10rCR26nFJyEd
VZVb9OwJHDb5/EAQO+PH8ZRE7jllWNlJNCbqKQhpo+xLqGi5bMOtzDHCv+0QNw8n
Za1FaHoVshGcyR6gOAjhRoykRLSVQY850d4VlBYLhOuAHYK1M2QRcuiEx/oOx9LN
6BfHU1G3vszYvdjy7AcGOes615tNp9WP4Bp8WPYLJC4EwIjLHwD4z+oaLHv8ffDu
bYIiTr/6eOnrBbJL/0ZuuvzOQyyh4FKb597DGcsZGjzkCHqyPigta2fVc/3qfsG0
zxpN2DlTn1+K9av15aIJbkriNhG2eKG84V3t03zyGrGUe56WNZbtDIBsD/1o69ag
Fjyt2M4deeUdZwMHhlyjFK7xlTWZqlcdCbiPvXFZQDnhUiNlFsmgaphjscndvNpT
cFyMKTK0EO7/9GObb7hULZI9R2Ta9rH9IOUZlsNqRuVoOL+83HIO/1MA8EfiULDI
6+MlNA8If/NXeprYmAHuKRG/CKFFTPmTzS0fe/680u6F8HMbmDCh3noeysHKPd1q
hNB3/pBZQ3yfv8foZfi+qu78cX8zROvXT+GB4pEaOgdgi69voXkHousdP2ubLHS0
xBBRga9nUOBxLlO89EUM0E9X49JYyHDGlsf7gwaOboH7zRct1TosWtiKWGsd6ahw
EzHsV8hXsLBgMcKtAH9u+N6AUHQAZ0NkQ4kx1M9SYGqQGlu9SfHWsq0OraLSKHYD
2byljocLDiVSbH3ble9LL371JcXocLKHA8ePlSUPXsJBTb1IY59hEcRaLT3vIm+K
ttt3+Q3pjgMVWYn273SuZqRbs+5pSqSgWn5Is3Yy0mgfwlm+ZWA1qJ3dERZcJL3J
7QD0lQZHIzUu4hc0VynUAlOglwMHMR0WkLuKewxBt81ZGy17755nvqMm2Bq9em8Q
0dqlykyX4BzCK57HYI9sXOB2fHIi2iWVcM59gOsh87AlWk7IWmu+6aj4b7WzR8du
ef6aYkQZMy4hbBFSVCswLebITsJs1vaMqHGeHyPCizhfCyPYo6CNFoXqFORTmBBp
s2zVLAcYUKqDhWcL1eaOON8iuGjiZhUfrLE6BGL9tPWYaG5nuv/1K5dcWBKWL8wr
igbC74+3/yPsleK6ZsKGHyGkCm4HyqYfZRNVBeLsT9H1vJPmVYEinUFZSV0Du+yW
T+X8bDDdDQXtvMS5dydDjvqUUCH2i9PDyXVnu2K2Cri0RGVY8kerMlcmzKIqfVFk
3xgf1HwljS+KNppSjrNKwrZTQapK3b3OoiVQJm+OfUlUWQ4dnd2v23prsoDSYj5K
vk1nlAUi1bSFe86w1ifn3JrJiGkXuCIBrz/hcwXH9m6YMRdzYv7MED1B+49jHWVD
022w/72Z4prE6srgZ3dsOiCe6ZHXkYWsOJnAAewD3cDSfXuwAPBimIWdmOcfLgLW
iOwkSDsqCS6UhfX4Lgxjpu3UQ4Do2QBJ/yUNl4HrMzvnXQvv+L0uG+Twuaf2emWL
YmWCyHJDWXlyvKWg1Kgs9XkHgW2U1PCfvQsIT+OtAuhSbxivKmV3zhQF6+CY6MlE
DPttlfBsUjnei4nZ8gWMoecY+ss1UEzp+HUkSrPj5VGhtHwn18ghbBsMMIgyyTfU
Ar2/lpEa/2nAk9SW4XjN8vrTKAQaDmQnaZZA6SHdgXsRxoQs9taQqBluY8SYt0lL
+hzGvxphLaZtrO2ICz0zUnH49FQIMqN26HCQ6VTvVbl6CAEQR3fYCylWm3irNE3P
QY2nKPm0mBfcPoRjEv+gq1GxNjMVesPYI9N6Fwo5YGHtLmzB6D0aiAd0W/PTCgmm
30KgemL+hjneO7zYYsVhJfC/6Sp1NEGPPaFzkil/QTS3IiIoJfaiam5nDeF/dqju
SMwJ+LOj36+EiLOe37SDjtX4AEf8x+ynDeTGs/iF7Hrtigjl1cd7gMA7RmfH0WGe
VOUwv9zst012yJ83tQEEgC0fQxJlMHvDxjcZqVtBQFgQWuT5S6tIkJjLznXmew4p
LWZW7flsQxMrhPwVIpYbFjJ09ZrXCEkbv+z/Vo4zOgUawJSI+yRMTWBnJRMrTNAS
HuXYjV1tc3LOXZwH87xFrH4omX5rRSBDCtagfKIC7FnMA3kgTRJ/D32oZpdgX+0+
f4/at0fpixVU0ZaiCVLC0FSNhZmMZjvpO0SXTyC5O9Mjns/58mWORuPOko4jf2mE
vudAQEmN83e8XuDV/50ybSSK5agvvaxOh4nxiTnEWsT73s8iUxbKdOglRi4Xwle/
81HMhHLxV1J82tsJfEYG75+me4Npt4q+tPQo5ynNRKpzSe4wD4NDsBwjUkBd5265
QOQQF04OEF5Q6l69ums9A1IHRXfpBOWt40M/oPT/xOVCeQYuGPTeZh67esrfCQP/
6S64JH7XjdnsRYx5Fu/Zib7g2rNRLc+rYglp9ocPrMABkZ0Izhr4QFJl7Rn29SZ+
6jykQEhmt8p6wwAVuIP4rAnEqKXOIsfg6uzEhAI9ofQDJfJurIqhon0gSG6NayoR
lShT4Sx9E451Q9V5IoLRg17dRhHEDlenhC/Se9WOLwzUZcbHjQ9D7/FPgXADYcIE
jonONHAaiOIhHyLMh1ERfdF9N+dUTjN4i9xD81NLoZiev9aDbVUBO6/cKZxX13JY
Z7rmjnS6i/8bJqqJ8LmQuPkXkyz4DC5ZfCINxG8YCEwZc4uWQafvdsOj0ao9club
tNcMO84octYe80VAaGaL7V13JlDKBHZzUTBydQTFIvG9uLAzjAtXLUd9Wm0OokV0
HzvW+t1u3kywPDGvaX4q9IWfcX1zmsoYACNG0pFzGGhIchAjL0GJQ4OaxhtgMVRr
SeUDqwS9SStOTLxvPjU5/R2e2tZnHCrtaOYvoqEo8VzyUkU4Y/kZ41GkfuXUAh/O
QIahsuVWeCVMuhPpZFuzlQrw2HvSinNS5IEQGJonVXX4YygrZnd6zvai/uJDvV0d
tUxKnoLy0mZB9LTOG4x1+tMPkvpUD0nf5ziIilr54JBoyI2XJkxN3YAkoQ/pJe4A
Y6rsBe1R6QC5YAV1wLyfzsqAAXnqpXDJzlWdS8HNMorDQK8Xb3c1gS++6su9AUKE
lGXDBf6AE+PQ9ikzfFnfjXJWLtCCnK/PFuH9gIMsivJgqum2XYVPgXP+MgQvBa8C
1hpX26n9rZutZqqoBLU2R1pZIOm9iv88NMTePFYk9CxD9rI78cU+qGEbLJMzcTz5
sYEjIsbLFlI4ei/y2AJZ3RZFHMHH3csSBrZoqDhzgblpANLONxddQTkMquIYUCG1
xtw2jLFVjtj1rreHSgkhmzTNcGGxSqLrMrYrwSBAvTDhKIOLPk5ssSiAKBrTIpXJ
Llpks4Zbnfmv5MlSqmzv3P5CiEv3DTRnVJHW2jr4tnnT0n7lwKfXNFSOwLMtAwJ2
Md1Hel6c8tF9jSLZY1w9mouh3XMjiS9xPP1G9IyTCL2HSo8q/wtL1gFcBzsTQW8T
hvYGnlongtzmlaimEiE+MaDH/A6dvrc98ci/yP/f/NqNZypD4LtrKr1mGwY2ZN2F
BYKMoa+cev+wS2aI/3qRaODv+C967Ar1Nh3jCevZsGbJCYkglGKvhjG0Jh3rri/v
F8AspNENpMVluHUwnE32+qMvPxqnv+6+wGz3yfvmT7iYle8+YllqU3pAigdRMeSf
dLSzQt96gYqv5xPwX+32Ulcvac8QQI+UesOh9hIJKfwbAdLQzOIl6UB99wTK2MnI
AVjIdra9ej93T5v+chM6b+z8xgD2OZprDMVzNzVTlCbAnHA6o4V1ZkHWmRd4jU/P
OP5qAkjTOPVzLR04DSxGY5IR0bGrfnfdcF1tCX89kpt0ubtQGrvv61Ugt8sZDZP3
HriWY/O8iYUoCi1EHuQ5rOZwSHWWztQvsa2o93/n8LdDhdgFRmL7VV3Gg3yEIWd6
Cj2bAZTLVsiXd/jvHsY6q25S1PVwxdQjYVKH1JW70avXuLIIGLxkLO4VU6BFY5yR
vmgBAYvblqid58o/jQMiLwwVPCqt6MpUBnQRLFAr/Hu0IxpTCbClyA6KFut4D/Bf
lPOOP/dLR+o7ZK8vGHV2qYSZPEVS0Jcs+eOpfbfEBzTTu6f7B6S4uVCl4GRieg5b
jl2Fnj9LO50kVn59Q3R1ehOrD1OfXpmVAHN3CP6TKg4hYbRVplxs71LXQc7TmYYJ
wqDGLMqRGq7Z3hj1BEwzJHGERIO0xKayvquDqzRHdRh5Mt7P13aDxP3ImaEhYjHH
+q8T09IX80lWH1ZH7LLPs689hc4y4OD6XFQ9VouyclAsNd6yTplcUAbMVzjsHih+
/36qVyGC5K26GGh28MlYdJibzhVsb4RPekRFElbJKDiNrpq3l5wE39PJ2dESnTu8
GPi1aeM/fghkDwSP6jlne5xMEQkOy7m9QM+u9bA+inn7X2aFpb652WPVkBw9PMzQ
IEZ0Z78s+aST+Mr7DQqfzhzYqyf/J9wcsVYsdsvgvT56BbxArwQv5swgW7sDB++a
dtPJFYsV2lofnS8rV3xhUIsKhoD/4yqid0uMzF1tIezXj4ve/Pzp7XotaaVCzFjA
MzKWh9lw3w8VHr6PhCWFTHGZ2vjWzBiSnLspYSNkGTaCBB8aCWsNMydAsQ7DuLfL
5u3ZUQ0XMAjf3JzxphJCC8iQvzLKH0vwke4tM89Ed6VqLhfrect1IoOXBQoErUw3
fK2Vt8EbrseS9LvPs+j0LzHb8fwXmBXKkZu3sxQi84EZ8vtK8oFpK4E9Mxe2msZ/
xg4zUkFoGtFpe/u0dBAi3S6X5+sHBWDgGrDuTMHHpTr388IpoETdCz/JvoJaD9Vj
uXQKleoITXOM9I626iSMr2DKwNv1Nvybt5Q7O5lL837ArS3SaqSLS/UQqYPr1Jom
+PCR7XH79g/Ddbzh2wDl2PIsigsi3hkDHBjowysfXnM+qgTrj+nx8mwPccUC/AXa
COddOCJmWeQFLbtX/X4ZWrPpfzIQoyMsVpAoxZedqIVYdr1dq4o3VEv0XCbYdUYF
xmrinkxLRqLydgyvcKFZ0GZKkkQ9S9ioAU0D2IWh7esW//Vso74EngXHwa+z8pz2
6Q1BntIkhz1FM+bdRikQAE7DmPZ7FnIy4qOX9Uie3XYXu91vIFTeUJsLE+aXubbS
adxAevga5oVkfHt8/j0DTUe4Dn3T/ePX9FoFyW43zLqtmAvfAXgOuPQPGh0WTa/U
UFTh6dm+sBEecggIBNOfKGE38978lsoNSTqv54POyd6qHwXlkZBtEQxoEAld39Tp
Z/bF2re4eaP2yBO4Xnj8b6JcjyTyNbSrPYhnxhqcO77U02iRbjTLFTq7F0h99wwZ
lsR8qNm65kIKrpcaI0Bmwc1ObtK5zmqu64uXOtQFxVMGE4zKOfHJesy/7Hcwa1rA
CIq37bnCTr3i/VPJhKWJCN04fNMLJuFl2b/J8Q4d8l/qIyYd4pgHBHeuQ3GsXdUB
Pyu6B617RvuSF/TUC8wXEP3cq3fqqNSTodCtGBX34QQGiVjqkEN45PbnSJmHuR9J
ylQ8B7g4GWiQPOa/wy8oVAOONUtWi2nNLEOymKCuDDI47tFfxaiZk2tnqiX31+62
ou02YB/ywow8Xd0oMWWp6vVpYFKuzCJtC0Q4clEyoKwTCBIpZIJCuQF+RlpWgMSk
VNZd319Xf0cmCUsN+Y9Td2zoSnztjV6IT8zlqxF1P6o2ttplmM/8HCardvpg3Asd
QYiVk6mF26yVTWGxkwiWdsYUFO/VLcdojBSHS1zKnFsKfhqSYkjQOtE6++HghJP6
iy1OxVjp8a7nEu3WcHq9x/IFuGKmFtbd7HY36ac1xmFAJt8caoN/gdhusCzjA0bM
On5LbJnPz+3gMOmzPhyDceyfbLDajrg7G4RCgmRpoR9W1Q5jk5aOX8brj+Gr9Utd
QF1g5l8v8ndMUZvUgZq8q6zQ3Ow+183B0aupU/MKLVozjY0k08lXP6UF1xSqImmp
lfCQK6QtEjMWd6AQ3kxgD7tOEmI2l8jG9aBo71JMGNdEs83MVezoqKSBVgrcp6dU
HiKpyAXFMJnpOs/9sSoCjeHHfFAqBhhoubzvv5qyiZPALyNL7Yrmel2KuAPzH9UW
eBm3rRYRkyVgRoUVa5bLYcBgoLupFVwu/T4Qg+77kpe2NO2v2nQX5QtIDng121is
Tzsuv2ROmA3Wwb/bDVmugD2eqV9jxua/8nCtjpbSjKAqRhCEMacz3Y+1H/T6IUx4
4/i8zZOv5jIR61V8y/eDbZ7K/G22HE2NSC8p7IDyTiL22RW7f72UfAIBYKJTXana
bxffzdNXziGOzTUqMg71dPdKgu8wjHTuo4b3z7wMlVsD3Slxp/bHjW7CB8tiQ8Jl
KsU9Lh/gq07JN0/gWywFS5xExIFumAOgpKS4UsOZ79MKKGzb0xKEyxV/eYgGX8lL
IJMP4PXleyGOVdKwB/3zhcMBcf9bktPzNKH40FxSSgYhdk9Knbguc9eT3vSen0ox
sNGB01DcMKm78cUPbNpp0KqCGBpZu9K8tm+wurdZ8ZkbFswKZQQMSzukQZjgxjDx
qD7/QRaLRyhcXiMaHwhvoxNHrK0LV/Z4KsvPcquUmy/VccQJpK9OWpDw5BO/JB27
AkAma05SsautP3TjzzsnHkhmBkcAZWPlIsoB5fHpMHEOd8ErXUT2UddtUxkCidmv
kRfhDDl7/AfpFDR7Q+FaoyWn2lCGtMvywFPrTjwNtiCluJhbZL9yD69UftqCHhDS
3UoKl8jW/SzVjLg3U88X0WoB9oy/saKjn6txju7ULyU2iO/EjG7MYvsMJ8/lNqpi
mF0EIaJ7Te1eXJ5vcZgxGrCKsKXtzA7AJVI14gN72KGxQj0megyj2Y/yOiWP+MRW
13JK0TU5pgUm5a3ffouth0M6hEf32jbY3Ln4i6tbLZf+sT1gvbKwHl/hL7dI2Tce
1U1VoS88XKGHuC1L7kbDaPIgXoL4JEO1suUO8dL43bqjghaIoX2f8zWABaQBtJpg
t6OC8kQ8lnbiaeMtLxDOnrvdNGk0webETi0M9E9Z2KADdSFBjV1Qspcy0tsK/Nhq
NpghE8pIn3OID5r7mEhLqY+u4AWAVrOs+ZsI6l5+5907DQgAqU25+GqwIoW//4kd
jf4QOM1r0NP06a1E0NeFnx8BI2bX+1mqkIi1Wx0A39NBn4yT1eQy33j9l1Aw3no/
Mu5wWMueRgpbgemk30V7pD1qYhK2PyiRYALM0gh4eScqTyq8PrHV2urAmAi29UTK
UtSo6WRDjGE5RfEXvqjXreuFAOBVpAmZc/FZU+ALTl97wQTNk47wKatNnXI81MmX
ZVpk06Xiq3NsmzRXVtxkkWUYT/xqgTnn9wlTJaYDJL8UHAg24MP3SWrg5cgQZBgm
eG9qY4iZkAEr7lpADqh3RZDbuKcuy0Oz/Q9/K74D1hhY5BsKkLFJGeLGYk3lWlsh
1d2OuB9dASDM2YKDBMvUhSiykHuYeI5fgvXdGNXTTkIgzriV8VXAvxTfZn01zXur
fiJYaGpp5RohI4Hda7xTkMozAFGOISmXIDDfJvJIxGJllWbCsIE5W2ppjkiHN0RI
Epk0SinveZ7ucTg4Q1PQtu+FFlRCFsXLl1U9svVo0op+lbnepyKM374k8S45jD5O
Uzh/d2oFAjKdujmASTungh6vrBjcZipGj4j9lHjfJiP1cmIjA/jd4EhtjBLi7qIk
HEIHebxKu5uU+V89fw4UcQpEZyd7tzSY379TcTtj/Cxe0aOpHbmh2WoGkFgfYoi8
XseuFaDl7WBu4bfq/6oFf6RlBqfjVg8dZDz9kxOIvh5/S5T65ImQJt+ZCxvAXjFc
rhfwndu/gHvn64JqGe3ELpouYsI1Xyx7errOGbpbhWfZdebdOiRQOGaKvfaNUqZ4
NZzMR6J2hWfsm3xOsYS9TJdAIeESNsgVMVmgeWc1aXpEscjcZ1QDumZiabYozH4W
fn/TtO0S8CLsQVGTCwN5NSXsYvEcp/06gC3S2GTncaIVCa09A8inxfTLstEH8wkw
E8I9ndLHdYcDPu3aBPn7Ko6c9GgnVkKhlTatVH0pfzOrcN8PuUshkIJaotiLjCRn
jTu+9jclWZ8PneRS6HW5HBjK891atHY5I9Eh2mjSrlp5AKHDZ4XbAx00OfOxxh4q
hKT0iWluG7vfchB2YsjUQX0Z290i3CkYZew4/B+gzY4REQVqQW+Q43aHz8KhPnzK
6EgxsFZ/8c+EykLKq7skFZWDDbJecyN0CMtldRaTXVGJJP2JZ9bsJjr8I231Bh2o
281sxQdge1nDDn/J7eCs07RBnpAXjkSDc6ysRp/v+tn6jFUwOTmM1zsXbh9Cr1cE
k+bNpCF3uK4lYoqWKUc8g0OdY/vQ2RbzaAr8SbM0vvynf/XNOuKFRXnOuS2nyFhc
duDTveAi4m4ITl/DHyF/37uPJJQ54dXCX2FJyPjat6+ptdA8PJb+AMgHrG6GFQOI
Ktob1E7ftco0XQAR6v2UuuqS5ofYhycEU4IcTAI6XdPYuHLltxZjmexxEz8LHqQI
keWgMZEbhL2DEdR2Zi/1/DXotq0b4QaO5hw97kk3pc05JOZcapodVgk28/p1ky+E
JGyd734/C/dgnBRPdKSeVpFjOBuXZt4M7xbIqezWto1w19eIiKcbkEiBcMHEa5rN
AysxP1KOm/bTEUFnzy0bapt5qEY4XXpD7n+FparrLVkbJHiZxb0aaG3fJi+KuNZJ
kSXFjrmUhl34NuAGWDqNgMg6SO8wBeYyTG3vsRwRpMRClERNMG76x4Hyxk/N82yT
1hD9iUgUL96G/cdVYz3G2ezZw7nvZt3IU+WIzPk/R9HCEp/3Y43Pn6I62S5XTB6q
ufpuCMxqka/y2RDboR9ZDcisPzT8romcLFw7Y5bjcultXB3hQ5jXIFnVbFiIqN+K
3edh0w7fNN+hC1TI1LzdAuv9O6mcjInjEPOJO9LuFlO9IXcrrHiAeWK7sk5+KUHk
tP+e94BBoIp84WhfOljOZAZdQrymIqGxn6DdWDqXMAaX1U4LLLbf5AOEzq0kURFk
Zopg9o6LyiiC+rGcpHL240GWPTkvr74bSLKXllj0jUlDWZ3H6N19bGO1Wx7ET4kF
Y3gPCL13i5yzTa34d+W1eiTBHvZJXc1GJQ/2P8ls7k0Vr6KPgQwQKOaYuZCKKvkS
cuA3mys1nBqcQJPAoM9KJZb31qDr498UsYRnvEl1CoA/9swf8X36d/gJRLiMG78X
LAHbJ4MvJrHwVfvSAwyMgOYN55me4HxOLdw12Dtf62zY2nFdatXE44Y1RFFjqed7
oMN6Xg/mt0fChoNOdvjOojGqPQzvZjpmuQlrSgOGGqpzV080tIC4vUpYnBwbgVy1
ZdpFLZZDO8ZXl2OuDO6vXdyuEWcWR2GMbq2Ddf4u2jMi2xu+nDE64nynWmhTeTDg
gUoTnn2op/9yl8XWuZBxkybGFcerJ1w+fCjdAbgr0aYDbKu07WW+JRZRXh0EtNps
HU7SeaTno843nfzk2bttcQFqVlhWOIXqT6xm+HepETdnbFrGZ3oNHPN7tj+sMUV/
r3MGZkxF1+DJsiuW9hvkVmc6PC3qwIPi4ODWPACmw3EtNoKF79/JOpAtae+ftPXy
+dOFfAy2lr+FMa1gwiuacO+qcVVec+xYwj/bD10cAyDiHGjNHetIXhv7R7/D7Ilr
UNXXcY1qLV5Gjayd4rjrL4UCo+Cpcxw+BVwl2Evwo0BKC9w95yC83Z72SI1KlgYl
oItWJH0X3c2jisIKY36yl8Gd+4yTKhdRdiJ7SjQ9N7GM/meMw0PiFfFZG+vvBUL3
bH65OuO6dUMlRpBWkNEgkxFVscgiBKQ9MEn9rZ4iQWcRRlHCAOw7h6Mq519Btzuu
DQYWr0nik+c80ZrMTRnQjnYM7BYvcjxDVNf6O5IMMQYedDDrlsjzWo2AhoIRicwC
FGdy8dZv3z04UyyR555P8DagwCR85uLY+n0Kuk0AGgPnEKtRHtlIgv6l6s2UN/3v
wA8HLTo4T9DjbkIn8MnwW7UPPEIxgduRditGjy35WeVREU2YGgitZKKkArNfgNlo
g7Fn4QvUzVXTmhox/MeIZzEEdz3qpNfiVTItVchDntbkVClARWv4E5PIztMsGbVq
3Uh20EJHhrUNJSO78WxGHaUtSvG3lBrnoksBZnxPXbPJZy73tQUjNg1En+AQ051j
GsoMqC0ZwDVRGbEtw7BsFiV/peYyfCapfEi9wny9LY9LMPIIW7c747Ny5Xatxiip
pSdgZyoyGkbpDsIXqCsHYlmJe8n7EjGdUnFk254HporwOW+a4aMLcPZc3CtMe5za
K91ELA1IiUwPU4X9iqbFzen0v6VBGZd7jHdWE4NHWXOzwcO2XCpubz64jzfHiij1
GmptG6KPAFbXSQdAqdJGezt7+p3ORMcPEu9qleInL3WNJCapHHqDGZD7uTFY6e0X
/K/PtKv4TAE478uk8g2sH56TLGmFG9bBV1FeP1yZnWAM2poTpYc/Vrr4sPI1rU+/
6k5qjUMNuEi4Ifxw5F395mdVlIKVOuW0Oo0/RyESv8zvnx2k6BgxjnrGaq5VWpCw
UkaAjVu1QMQ8e8Kx86hzhuEtiY74zicAqXZxHu0aW6EJ8KpvnR/ZVL5mxyOKogAO
y9ZCpFSY79mIJok7fVIspcLqYpW/WmiSHWB0o/S4Vq2uXBSI5NZEeVZN6VkSrxzj
kNvpbbNoeUeC08/7uRPgkSnYdhRQaptnKuSM72d0we2gwl9XStMoOguHqCtMuWc2
tYTDxnIv/pAJQz1YriNjdzNIsuwMwcMBEf/ifoqIGFidJIp4VPfp8B8eV76qVkID
YVhHqBN6juwu8THL7KK+DrGTO9dWADAcs4cs4EoJofUBsKSdEN+sG0rATk+VlnOU
7VA7m7TnN13FqvsIDqAqCC9taqggKyyfxEWqz/4PQiEQIvHsellTDIllQfMIboYG
Y5A9IX1MAhDWHD4+VDaUGmZZJiDYvzS1id3jV3KunCICln9QsP3+fd5fm6UYja3K
8ohyjBTseBAMZfpGJkMkGyDeSS3ROrr+LIOsF6yc5wtR+DbDYObN+yHbhkwk1RFh
csddyR8hfjoiQ8ht/ni36Ftp4M2RjjtqofAR4Rtl2z9j0beAD/FM5fAUfj7eaYR+
75KpYga1R5DXypyy0DjIMuO/Hp+KylmyBPrPiE8nF0gAK8cDpW2aD/5Uu9vn1Ak1
qVqQ0RVeO+/dOXequcK/LzjJcyc2nrf+nTIVL7BegO/9NGv/KMTOQiyFwoGUFQyy
MBlWCdlTiR7R/7Td0jgNsNS0vablkDTwARVeOvpmxS3kYdeCkKV4+6OJ/s8o943A
rigqxTSgEfVMvPdF0pdTHpewk+psxQCVQjMzSrIjWOh/zaNAvJOR/SNxQ0db18+9
FifgRBJTSXzky7CWOIZpyXxAzo1pNZKrKy9XbG8XAoaod1OrnfSojc0QRlMrqRAV
BrYUZqf8IkCvgMuSaXlYaD2N9uNQ+QMlBwb3D7qp56lwiEcFKUxEXjRuhBlcVCBy
d9plnM77XCdIN8coX2L8+W6+vSQ3CMYJOpr6ha6G2GLKb1Fv8/9hzM7nf/vrY94x
nVLqfqukvFw4pr4/nfDq/3r/no+7WyXKt2ZguBpDKLqhWAJKv4Ai8zUvHdEjboH3
3fbS7iRs8tENHxLK47xdloYR0PSHmW+dHJNLCicFGCfS1CfFCchL5PAeh6POHfyN
coHYHRt3ZMCYx2EiJV+yhycVwfnFYjQgvuExOGBJPfCr9WOeLE47/AcCBawBIVWp
kb9RyXOw9pn/DD4cemIt1wgZe6hWJFpXviQ1tmGtAcBErq82zUgDZEKjzG1JT/91
+W8SK1jpshoePTCzB+nVvHTYbogIltkQSYNIjkwCu9PLbRaEQkbQaW+8XxCOko1C
q8JYBxQalbL53WYe+UuoCTUiscLo+VulDvybW9hUptqXTrbU5qMn4CTJaZaOolFf
S0aagrOsU90AFqBlL8RbZdKhkFxTG464posX3zLpjBToSuv7tRw3aJ1uKNpo4TEC
onqYyfBlJQ2Wsyu26C9PxJaiiMhRh+/3ygbpJi8Ymme7r8N95G6OFhj7HS5ZZO/p
Pzqxa8HUrbPkfX2tF+xHgH33Ra0TzdeEWpKeft5KCl0elxgzsbtz8XuItj/GG2Xg
tXzEsgB15Yer5j5RbP/hX8wuU0D7QrOX6BLyYoKQw3tFiDuu1FPvaNeNWv0sP1+t
3i0S4Bzobe3cy6J3DVH3Gd0v8W+7NoMX0RDIXLTeLibkmREQ+4H7p7OT2MxXtz3n
9dR9hD1POQheN8UYH/EkZhzjIneobDe1zSrKGKRUOrxFgeCzEu/Zv9ZUNI93sN4N
x2HMalWWLqqYBYxVdX1Vw9Mk2O2dzlj7n45dSnIXOvjitGKxSkoOXX8dMOAysnab
jsipxtOtkOT7xHfoLxiWIm14/9UCazLLcYs+oi9im+0Vs9BApUGSzlbC+n3+9SEr
7EB34QGsYyyiQHuoClnWIk9W21XXi4UrFODuQ4M6fz4wySQE9BUbCDvuOsGcXSoE
krkEg/yaD/qITI4Uy37KuhSydOAyF13I9nemEkTbXpAd1cBGRGYHH/IQPTVsqWBM
shHM/HaQIyC7F7cYS2of2gmhqjjEIObWvSiBPoW2hH22s55WzmY7vfA4SQdqXCBf
clu5Oa/+gl4ZgMRSBx/v4Tg/e0nrOgbOf5aWBG8NH6escCNrgTDqibS0l6fLPEXz
mzMgrLZ+5qHVHcLA2ut0zkGszd+2hk955Vu496w3MC/xA9MKNxReZjet7vPzkPmU
bJFmC0VpgM8S85H9j9pNIskZY4HHsW2H/8uMlvGrPR0cX1WY4+S39e8Eb/hsliBU
3uIjAr17z/YgZGWTJIK3k65vE2/Ren3/4Fg2FN9FZMJWbKr3ZhLrCPAXFc8l/wCZ
uIRV7zPWPcfXi8OxM7cgTPds2JMyW1OduxV+mY+be2vlqKZVQqhyDLcG6/xDNlyd
OzMeTmIjT4HlC8i6Otqrc9s/UUNfRF3zx7ePhxVFgsiAyV+xXNnH+HynRhqX6+FT
gkus2UhvRlXujReu+LIHTL7m+P2oQ7Ds8D4Qlw0pisTuhtfCFXn/aVSo/+G6rb/0
kusjUh8AK1ZbyJOkkrsEealBNhElfoKjrnWk0nrflsnhKHcXOyrNJwUGRuwKMmpX
9hHEdxlLwAfLthKdqFGkOqBjCQDbkAUg6JuqotKNma1w8eAHAixEt2t/9iXGEIkD
S2WHTOsM/gofqtRoOIzDz2VPd6AS854ra6xQ2weHkqDlFXq8qHWXp3sfJ9/5CyYe
htn5qTMiROyHRxlRCYaKILgNOzYsqnR8pcXr8SdIUvOAbBj3dGf2eqHflxPnbF4N
y6ems2U2tWPLkgDcNp0hQ4Lyw2AALI4f5b1DSkj2f5DurpvaYHaZgpKrrHUm0TCm
BxkAgP7zwmZBxWsr1HU9o23AsMhlJ9LHLqb61k8FrBdua16iHCisXwe78GCVhF05
BGqlm40XWox0nIV+Mib/1J0sBVOOi/pbDGLKGE0DDP6/3A4oSZxzPherrc0lVH5u
RtkTa7evx0eBe/k8r4zsH5TLfB04yKbdO+M32n/wKVuWZTkMP6J6YCCiWmqxLRbF
kYtjSsDljLncHDrUZOHpvzjDwPFOV7WqhjnZV2soUflNw2ZXOseMXSMlvy5P/TzI
N3K9ARiiI1AYkLyShsTpMuRJg0rQ8yXg1OtZSbTsLAAVu5/XgwLLj/XmaMlkjGN4
0EPMDLUPcVsUX4XZAlNRYetHacyUN/Rz67Yjw1310g2YvO2+KTmNCDQzjLBoU5VY
IIS58j5rfvfVamRkA2Oya1fkt7UlRt6GcDvh3EOhhKOJ4Y1x07Dve4CVuxfU5g+I
wIT5Hrkdx7NH0t5DfXuC4n8cZ082Qxp2aN/vZwIuBsDV/R3CbOLbgLrH2hsXAAoL
R7docmdtjQ2l6tqBnvv7/7CR+MjXtvODez23N54atzRqpbraRIUoVdJh22f8Dl8q
hNbD5PRAQOSfUT6Ay8F0SBm+en5vzJPiWp80j7GPgJWTsfnPyRrO8A7NAmj3rktJ
D2tgxHR7lXZ8AndY7uEQFtZROjVM8QdHpV49ONKfH9Wor3Xk4GiVRvr4+onUdRN7
wLz6nYLtrhiy8q8PpoX5hkRAWm4IlFkcQorz4HaZbqNtKSz8q51ZNHEn4+Cf+fKp
tV6tei1TIDODwHmHNNWCMnw9AZbhrekHs2zXq/TvvvEXnepzf60JuUcPrbruPS5H
tnCXZmvmNEvtYPsXhvbOWLrr4n5AVFormm26Pr/T2/9U9sd5zuwuFr2nw9aRJDv8
lw3LRnuOqxyFFjJQxcvwAq5qrCyI4jzIUBZAt+dDu318c+AIKbneASqqg8ZGOlmP
enLVKlgEP+w3uY/C8zHhjKceYdN+fjw7hyxevDbIS9M1W9hCSdVbfGpV2y0CJ8OD
pzUpaELASneqxI6M/saaX/yzjiq8tuOPhRDEaFdU0rB6KpyNxVUbo8GwXz5BkI9N
nW37PbyoxRvpKTYaSbPbXYknLoF08m2CzxXOvBQy5dFKLI/ceoKGKhNc3vvj8IRw
H/KH6Z6ojdC1eizyzx+PPBI3dQrs2vrL5gefDK3PfENpNHmp4S1r4LQYxK4AmonS
EeA8Q75bIelZwA0pr/syaq9l3eQFrgAHASUf1PzPVnnAUClhNI8VXJgXU2LuIUJN
wGn0kKCI9teJbrKJjCB0GU4JO6R6fKEAKdWkfpKaN97FBQ2FqpMtoZRvftwShC/B
LdiSTSW4RjzSBInkke4BrzceNrkaBF5CTRV9tzPiiWX7VRQq4Nz6h560MZg1C48C
pV+3PGuPqXpYMBbF35vVqX1m0IV/OIoSoONK62o6t0EApoZz39eNOKoSQJpU/5AQ
UDYnqFfW/uDk/MBsmJLSjL0AtSVvxCzTCIsTwcob9iqj97bgIEPWmx68OaTjpxdG
KeATofysE1L8L3YMFF4ZnuGv2xjb9Wwc5Q7QlCy8Wx5AmyfqhVKt6B4BK1cxNztM
Kj8/mGjpU11SiRuFHTYDUY1oQO9Ky7Oo2KSyxfjtx+sPLbaBLnlj28qTT0UAk1gX
ZQvwEFuDM6yCKLkNUw5IB+tOKWMs6uWmPrD3Q1uNMWhMLND+SIWcwubakXPQ3X51
fFEqWh7pzCz6rS/KKnEU+EHW1mqbg+lltY3jzc8/YeGg+ksHnKmZ/5WMWVfPVOzK
6gdJPPmD3qn6fdhCoQ9e4PrSOsuN/Fotgqsm44seO7/YpWyXk9XhkJDB7F6aCFO3
SlJIRglFcD7mDsYcbAdWD2S/7qYLYPvcUln+GZjzIr6pL23elW5hGov30BhHoOLx
K8uxhwNrbmjAfQ1cnNFHuVVIoqEznX63nco/mSvTXntUzmxh4JiLXcIEyBRkBHrJ
tvOit99+M5iDyrp4/TSGyGYjAXt/h3SXYcKSB01Auo8LeWlyoJ9495cgQ34AclJ4
vhjof6k2uN4GFGa9DbOAEh9frcO1g41CI/uEnxD34nWECfCN6Cz/igdMKZ/nE8bt
KCQc85N4c663Noy8mkndIvmSieRFuC2BNm/jEOmSxOX6lKV93odQ4RwAcy5AlGnI
QJ9IYRo2rm6g6KNq5Ohhl+CBpwt1I4whssgDq1hIQ0DhXyGPk95BRDOgwBiGQprp
o3Sw3K8+hwPILEbagvOamfOjpKtZdPOwZD1B/KcBN2gaeY/I1GED2V3i0agW1tgG
zYW0Xp+EuoaPXZZr/YZz44XLMGQwjrBqRlhczP6kDEbozYl9sIMIxiPL8yhPvY+h
gJeyJg7br6L9KvyYP2iQur81L/MTJpfACiBZCfReNn6sOQFnmv89tO5s6gvkbhKW
LSsBJuRFijdlBR3LogaH/Rt4Bdhan+xaDWYL6LicAkCq6/aIDgX2WaaHFTNURzOQ
vm1NNd2nTG5rpeSrdSfrHSVYg63b0Y8iXW7P8ICBZaln//HFrS3n2/vi5FTMgrrJ
gbHbfm1yqJEvGXIc6+YEpShYEzas2JI6pS8yPyPZLoEyVN6K7pfIABOqbjnAhAYr
FyQXWpDyCpcWnhLMBnNgCRia3pFWXos/RwEew+X1HHnDZqxYLncL0rAQL+7sXTgM
nCe3Sndqcb7L2DfNVRff0QfjM/StxfBw0mH8LcqxrKAYDzd/Wtxn6Wzp2/oCvPl6
3Oh6l9vkbjAHDcDCRvOuyNRnwMc2vyV0XcMS+y6I8uNbdbbF7RqovJbEkfjuMiDU
NY+5sw5I6XrNL7tg9+CzUTYRbFD1Y3hFBX/oIcgDO0z9rzodwC9ZldK89qMdFLaz
rbpTnTc9tQNPMbLWRleRGLCs3U6qZxD+MX5O8qxLjperat6UaQ+mOKAMEGmkYvAq
tg+A4+IxCJi/OHtJLjQ/J+xIkNqWQ3/LTvuG4aNHkP427Ds51drB8reyQoH5UVOd
oe8V4G8TjjvYeNkBvpjDzOKxv8A7lUxrih/96F0+ubVcyBYugACO2dbmoaguqwIK
TLPwNzMi3RfYVi/VRtt3q46F672TXlShqmYaysCR4YJfloflqT0ifJjhAvf8eZiK
xlhCsjgLkHkzZ1nzkq/ngwhsxVO5hXWFi6rHxKRHfDbAyX2LEDQ0rpoxi4aIBmxC
vrCjqBcgM82HA9PPPzLFWfqxW2hhA4F9o8zidXlFiWRvaX1llxYj27dXCita+OEC
8MRK92jiD+hvI07Xw/j8chmYIu5MZcPVUh4ovftNAXE5nVJyYc5p5WkSlQky+A3z
yE+Oh4dfS48XSzgazS3OfGHEAKBEZTkrvioO+FdXcTfAgn1KDD11csWcSzQ6CH4q
Yi+0iTKNsrGnEXZIvlg0kdWkHqZ/VciP+FhCRvTTUdlb+QV463BJeZ0FAJDEx8hY
xqPoFw5N4lAFUv/s6GlpFZMf6nq6fhc0x5lYs5LkNBjqbYtq5mr/o/xcIji8pUQL
HoJ3EKpmQC9B8WlEeQs+99sjlSBQdFBdsVFu1Zf4+7hYABwCfxywWPDdt6LNCXzT
mTWVZKO+eRxuP6kb8RZWmc+tdCgzM4tQoz+eoyn3cvjzV+ksdXoT1F1ugMkP3bNY
/6TrK2rlyBG7JaMNEey6d4mVegVmh2wg5mK9WXC2Zl7wX/I9Ox6IwXeobuEpDjws
eUtbu+M0dP+xrE1Ht0kDa1A0jO6P6seMRT7ljHZLerfttFSHga+qtmh0yN+kyWlv
iHFXxzMT6QHRR5pzeF/WA8mDVOvrGrZfxOnM6HM3o5QGB6hdsWLDuuaqv69Zu9Hj
x8oekRH8NPU5gn70HZ3L5yDIFnwtroJu3LHCa/uhsK9w/B6F0BMGNpCAxTzU0PU/
KljzZRgm/50zAVrgDhcQ/LDjCvESHWxgOtkNkIfB5dCwe0fqRiT/AENEi7Rxwg96
jIQouMBzy1+oGdrR1K5s/HZizeL9tGUwWbH2N4aYoLj9YSHlwKurOZ8+gXT+WbKP
HSNqoSGhiq/NElSY7eVBFVPcNadexxkVy6JS73kcN3FdVCRJg/R1mpMUTAJe25La
zw5wC7xg0v7oDaA26Ru2wdQHloQSekNDF4ODsH/RR+SuigUc/io/MaHXjH30Qd+h
eibFlV01+PO61JUyNlmLjAA4Fk4uk7B744Tifd5UZX39HLHZ7+UfFN/55xPzk1K3
JgYciHCkIOt4n48CBkEH2BiAAqtQRYJ/AdHTaYaj15FpW03PBfghoAcQvkaiK2vy
B9v4qmRCoSn7NQLpoei/Ck5bg1tI6leUr/iVcRryeUWBoRh/hiBIymlsb+ZuoeWk
BIo7I48v/uN1bbzqmum2T3kNOUCnpUv/MKHL5NUPgEVFzl9nZWy/1JLuBorcxjGf
wQNIYrh/suYFB+NUq5aZiQWxcUdszlU39F669yZK/uCczTcTmer//hX4ctl0E1kx
cxCVtq1XWJ7Xx8XbrfNhjw5ecceffWLVbYKZkNQJLHdB5iRqw8lpcu7h/18Qtyks
NbF5YNA21akSFFvY2KlYGAFz7TyB4dTTKPA0GCusENQ1VRXyu1jz1pAGaT7dQAb4
/lv2R5Cg7CcKGrPox6DtBA06idnwuN7ZNJaiAdqBU7FfSj0CY0zh1i/jTxh7qXVw
BtOTYc7ByfgcKwy5MysqZWMSpL8taOZqH4QofteF5eaNp7yQXPMZ4DyV349RDxJ0
u+a/nuLSio8SP+Z9TCZbo0PYFVqQTnMttOBeMRPJlSfcE5EVtE8iuQz7e8/l41Hg
64csbAiz2CbwKGXcwk8fSa+hBfIV6Rokq58yLZZq/TKBMv7+tKInCQoEKr4MuPov
HS2sWOJlyw8yDGp9u38Xld7g7WvLP6gSJhjNkdwcy7Q6IbRqqBJfoNKY5Pz+Dpi8
AIgbTKborPqvaMCrjvKQh2oLPfm7eavuX59RbGcYqlV5kCxgFOJJxgFACee+14k6
91i67USRAVz/RrnUYjtlwdCoz67RK0SqG7FiPuLSjPrAjMXx3Tzn8UoQ+s/aqhRZ
rnTe6XLeqz89OclrfGRpwJGX953tt7Rv+x62AmUs6GENPgsSzKsU4PjvB7n6lkma
bhOxCYvaMpGlrNFpZHbqsmg5DGWcSWWpmzgKoy+aZbomAMoGtKYzCH9yxySXiGeD
yieptGBr4YL+YlfhpQmhpmt5AryUzZo3mLO3KyPRyyuelKEZqHLtmCx0hXOrsfhh
QMptqybfm6clcB9FkBTYiayCcxXvZxg64WD38/etvNuG7SPnUS+En3pnEIWLYTCL
JnvCYbdAlZSu4uiuLrBkAHN+Tsh4jcxMctsJebasBUWMzJxp1KAxvwZXqLRDaigM
8CVaIam/eG3fLxcy4auc2fpf+juoi0G02twkjDj5bXE1in+gjVCqUhgxpzhRG8n4
Hb87rY2stkG1JfKUfisq/NuEmzCChG9zVTA6emV80OLp/gLurfO+918Bvs+kduje
ZizAAZdnq4Wi6Wdvu+hbOfyAg43/WMUjWxi1IaaT+U9IBb5Cgn5E9Vunclko2zqw
RMnP8yuelbKoEOD3Jr5O7qLP42WsIuhyOQwCfj/uZt3OhkUBbpE3vx1d1af+hsXI
5wDCPg7TC8InWQkNF7gYhRtWKQZNC2tT9EMyjCIF/oVCfMU/DudSX0CVn+o4zsoE
pCThR9vIN8CXkxTNcMOQSWyTTJD2TtupoScPtEpYJyw/29UOPUhA8HJwfLzjJoNY
U06FK8R5ltVRXNYBq//L3FPGyPzskiZzkmoNKb3Rq/TUf9AQZE7ajyr9Ollf6pVI
We2xS+hxbCKVKmAJcENTib2kJsGEbdvC39jkyljMCRE9Mzq/t7/TgxsFRGZB5s83
PRl5MmDu5dBIB0oGbX/u3Ps9cNzADTgtNnM4uYPvUNgnorrINq6Cer5UA5k8v6jS
KCXwBEz6gCujweNPAsQJc9MSrzMHP0zZ/F4YgD0AXYt0oQq+uKDqUItya4AzpTHo
zNn6DAH5fw0CEEfWQ8dEqNPaZ6Kw0co78deZs8zaFQNNWM8EIfhvy5P47oevqj6n
AkQNGmzKMq+OCTHlgM9AilJ3yinXPM9kLnHfZh7Q4GtjGfbFxw02NN750b0wsZHo
nM647j7Q731VbQgbqX66KO7cWx+9ZNNERCyipWuJNCZCR6hCi7aL5ASSaZVYIi1a
6DkAFCG/s3tgp5IkQPhXc3ozbU9YPMUMfWESVPNvNCuf4enuvhMBpJS+VIhAyk/p
mo6bP49EOZZnBovYCWt0hXUQYGEsuTVl4n+69ILor7b090HhDwawvtrTpVvkz+kZ
ITK+N0uNIeuDngP7p9Z3JiypWktk85kHOzW+IvhRf1nc37UMxV1b3w0Y0ZFy8UMn
dkIh0XXDqI3ZmVAwZ8bRh7FwuxRIz4J11+IbOjvuzT5lGTtmqjeeRvNKS1Blcr5n
B3LJUieiPNdw7IALyGmG0tMX942Cg/Y4EYboMub2Sv2A4OeyN1TJF9zPmn2nXL5s
aOIv92lMkq+0m6LEENhOqZeViUIo+298x+eNgf/QdG14YIuH8KhMIUZQ8+IoTp7A
PE95lqWR3E4vzD1tzU0orAWZACsIHiXdmyH8ZAfOAiSwweHy9RLkHGYIB9mA4Ott
BnP1Wm9AT9dFzZNnHhF5f9t9ebWojV26JNOUmjRCFHtCd0EsLP/NwQj8UtUDbap2
LHejR8sNZ3NvHYARLJ15MRRpomfreE33LHKS2KpclkB7Mi9V+oCMNYLXCZXpFYuG
NkcafnKFYrNSPVIrYQW5RHCqdHKha074TJLN8FrvlIjArdfpQI051TzyU92jDY25
bRFBe1tWLIYB+VrjhkG4p/7EggBHMpt7Z6BlqiUVzdDpQwaE+/CFVS7pPz9VZK0C
8x51qb7MCQxKyPJEGxOKDqa1pjEyY8JQUAbrnUXskRAReF7stFukTENyYdAubct+
GnxMcnvTMISx0UTnItWhXR2y/7pwUZiN2vuKsdKgYsuK4u/CzURc5aG6MfFwV5Tm
JTRCYL3PaFVB1jlVd4DXP2P7yOhUA08B+JidMGAn0dy7Kp35tC1i6o51vjGOWu8y
XCTIIz/dyVZ1dk9XB5bA1rFN0kNtenvu682Y2HkT10OndyaKscrqgKm5kQe4+zXz
AD9kyfSCs9jGGLlAcMMDXEYYJ/HxhgsLjO4WqsHUD34A6iv1tIRcRFagYh2g7bor
f86m8uqcQ/SIKpSrLuaqnyNEqo75IghObMDeEUKii+fUmRQ6M0F+WCrLqoJ9Ly9x
7TPJT8U0a/zmDaYQvUyd3XWD0rDSuTiXStb2U8OmrI0VPpBkRyPipQoIbqPjOY9z
GZeBUOOAXn3vyzWfjqKRcadY3jA2dkgI6hgy+zXa/SeF+my0TOmq+JfVf5aqo6Jq
A6mDYAUYczsopJRvNNVCY8ruTQqAYhMw2eIlay5ZpUIIjAn34CxxCYKj1slLx5gq
u2rt244ertv7md9DvPRpjw1XFsD/ALtnJy2ASJr0hCNW7mpuj2StAjf1JGd91Nk5
+u7/kk9QmeKkGq9XOzPMMwlFfOw8B1vZ3cRM9SXkxVsWwHnkr5ckzD00g7+fK8Qp
L4kRcwOBrMsR+u7iFNsof2V5TxEMBCLNJh9MCMXfYXlAoYf7SpL/QoDupf7pl2sN
rbcn7FGudvhmXgxQiZFoI0CJZnxyvKSjJxEQQn9x4kBjU7Her7aKjgDRwvEVbSjR
lx/R1IlIv0K/K8cOMus2DQrn88X7ZyzR66BUyqi7ybxUBvge105KJ9O3yKo+Nl6r
GASrwGV8RqZCtlhCOI8KO8QeguPJH2hk6oyYX4r4sUvzscytrs2WrGTfBb3Ziy44
ebQHFqXJLU6K2CtdhCXyVFC+dbl4o7szhX45TV4a5NboZYJaFrK8EUGu+MAzzgmS
QsCsm5le7G96o96QFASc952gNU+Qg4rLRBiHFhRJtaDq4odlaiM4ubot/L/baO8x
B6KXqb8ZkDqFvDiGTtGwb78jW/i1R11Ghb/HG4qt6EyHtcSP8TGE00+gginGjidJ
aIkgvpjYVb/7BVOAOtwM1UoLluz/ExFYe2fnm/FpMCWQTWxZVw4SWa+zUgXG+Cl3
ULF5OE2gRQhW829AYttA0q/wMHKW/zkf4jDqUEqJ73qipBmhvHchZoUWuCds0Qub
w+nbhyGmMLmDoWNDJm6DyMrVbeBIeW2PENWNNyHIOr0WLvRp/5R8GEcgLBQfYkz8
FQtNkhOOA061dVim4RqAhe1MAn+SgD0Ua1mKVD37OP4qKHftA+npxhfP5JcNNbqL
FNx9ZEtq74v+BXWK3B2lhdal5oi2ydaAt+AY+f0dUd6r1JQl5oI3DxKczNJZE/5i
BqTxd3e6HhtclA+yLD2YFXVCApJctmA1mBgupUhrA3Wxj1fawxAQ3I8X185+NnZl
xRpcltmqEqCLAH8QS4TZN5XoY/lmEBpoorAlkHp2jiLdKWa23liOXBv+UXJPftX+
biCgPQi9xVsmTJCgKpHF1hPu8Qicx9/fdFLN1x+8zhCmTDcRZMaUsKnLqO9VlVrU
/YQg7S9sHzZqs2QusIX9SNHrQtmpHSRwZxsEuiTpKg62uNqf2SydwpXMFZqLeZKq
KLOn9ybCkjHH7iSl0WBcBsAQcNZTPcc/yngcqMp/o2QrGMVf2hSTanSiSOR65CrM
icMlyIYEpUqt4WJep9Usck75cV4W0tg3hG6znLofYuXWVQOwFMwjEflyi7vKnqM1
lPusGGFKAHLWBK9oI5BnI8xvTi9sDa5hc0Zh+qU6iGnn5DUbMGOjnyKvQgimjMqr
7OZMBECS6IW+fa9fZxvmI3PGpLhXwA1Ot4Q9uphTS62+7BOMi7OBLYflA3ZI6H65
2D2arB4PZYXnwsK6+uqv1cX+uVYM7usgu+CB2BGg++vuxqydCiyCYGKRaj+exyBY
hTVUV+y4THL0NiVjsYP7oNkgY+DxBFG40QbwM/xAJYXl+yifpzfM+nLw6CQRTRqa
2YCkDEVaDRG3MHYoKT+NetubS3YwpUnC9LZiH9j9Jar9EZ7R6kzYDm+kYmn4lDTW
xvXmNbGdFkSff/qSXJ9gAlIRhq9ZRPHyhgzWq+OJ6J9AdcuvigKF+53+VjXO5Dnd
x1wZ4QqEsaRaxb2talheOcBhhHQV79VpypWL1tXMzezkyNETWW/xVc4KNmzFNOtN
z3erWKI4l0k7HKzz7TaJ4wnLeZlWDakgoP8BsbKpzOUjG/s8ciM++wO/pHUeveQY
8EYH07Apw1xEcfMpa66klLjXcU5BwBaGnWYk11PJ086EPt3YwJmeL+Q64NVK7gRV
SSW6DaO8zg4fVFg/1RekSPkDf/1jajsvs5FLr9OcY+15BPC0BUyqH+4S+LI01FvM
6aZu/EcPeR5/SRR/9OY4ZANe44f6tL2Vv5toQXKTIcNS5z7+7rctipwVowbuwG+G
afoppaJa0yZFCvb7YqTKZ0XSL9atLykFtoFmeFYykfumG5FkGRGq9qLZmAcP8QTM
Yk1hAU5LFM8Te0kehC2bedVA6avg53VOnEh42Li6plYk1x+XC215wCtKly4Xs/18
tIwqXwIZOhwN49NoJZzJd3Gtr8gt63ldS257xqCxNolBmaWwcyUXUjmKCgz30vSC
80vPIuIyicHxRzWWbIvn+Ld2aDghRttUcfUcGj2wfCfkDWTuculQSPMmSR3qCXxX
JZDOOnrmdSNRt2ktmYGLSzxxqK/1cybAeDR7ZsL9MjHjD+nWH1zOlsMPLDkQw6Rz
UuEbYdQBlibXxkto9svWl2MeefjIBaK6zYQ9qt7NCjIPdDZMeiFk6aLGIMGEFZ2B
KGuIOqvHEqwa4X7B7AjQLxAxP6ysWb8bEhV+jnFDfFEknIlHb+sXphVwKSp2KE6C
qtWeyNI4OD6pCQOX6qnRRxCLbcwFqBd+PLSMusEJBiYXF7schjOd6pbO5JJEjfo9
GY2uCYpdjjgIO4P4cORMkUTmYGAu/6bcM1Nj2xCakHDZnYr6Ehs54OINodzRNtnI
XUEMI5ZsESobBhuRTH5k2/3qUXg30quIpYjD19Wjrf3mlBFhzmg8njfiC6/BA+mn
1oyE0+SLDwyf0reeQP7dl943CblrhmG1FoHhFa6E6X6UoTV+gchMdzFYCTJw3tI+
vVrLo0Zw58Dz3AqfpseL0IbxcT+jeckUhSrWsjXX8PZEu4Fv/GC5bjsYl0fOcf8J
Fc1lsnzgMuOGF+tz9nEdpB0qwFkg9H7ddDoySygvUbKvsFzfnC6TbZ4i7N4LH18w
x/nMxA41Xgy/nEFTMRT0XEpSaAziTPoxaSX51dZKPo1DVCO5j5SLNgjPwOkni53Q
OMm9+xc5vHUsyLXmcskDvQtRm/wYCbcjJQKeQRuaCdKQEoC93Ffauu7RwCD1KZ4Y
+40Cj46ytjJP6kRSLSFMGscEEJUVtllg/hAWDGUxnd+y8gWVn/hJYLaPRLzItdh6
R1xydRMMb8soYC4yCgU/kTSdoiX1+JVj1iTAdJIuBIQCDHzCb7GM+ZfNLBSXRLgg
z/SmbNpLpvUvB/P4eAqk9iMAQosMCMKoX3Erg6VEnBmp0tiNPIVGCOGg4orLRn3r
ySKb3uaGBK/1/sf5Dr+4yUf0wX9W8M4auCe3FKwjac2BVBzsG9Fb+B07TLeopBua
EPzbzddhhoKbk9VtBTtyx2hYkXEeK/tRk2Mvw/wukzSXAjDMQt2+T3cuHTIFYvY3
z2bcfmvoNE5emMY75fNhv9YUkaNqLjWvFrmZuRwSQQgLExP/gTVptiwuGisic+R7
Bn3IA33gqypiddpn5t6+BxHZ4xG9JlzeTy6Kr+tDHnASsH4OKo/bI8QzrDF9X/dL
2926sHuiau5HxAx4jOOpELqdDRcMnoYVLv0SDi+0WJCIJ3HJJT1kTGEQRwCVmpl9
J0t7Mi/nFb6EiK5n7+5Trb2rmaLFavFSiVnZvg+fYnAMZdAE/SZZbyXVGlNP5zqe
+BcPGq/XDKlp43oFYLDwc76EB/jez1kc9Gbsfb/FLe7p5OUzY55sp1S2dlaSwdMY
k+Z89R02mGUYpzXf5LETTUCCKbGZ66C6qk8v9lwMFMbnR0SW82xuvTX3HWoO2hgS
Kd8Sy0d97vAHz5iMNd/MzWcOhGrTrzVetyUiyIMyc2AMmIEc0n7NSOJoL2QaTACb
pnhO7jS7lep/rPWemrpVfjzaW22dmMXdFlEZ/1Kei8Xn7w6i7IRR+JH76OOIV5hY
10xncGtTdkplmsL1CP6UO0Wo1TgPErs/P7qfI1snjchJiinoxlDUFFErsvPaSA3y
EcxEzPNEZcA5WAILJzANHbIlkOm72HZ4FPytmzqvPtqmeHX+ytUaaoZlYGnH6Hu/
N7Hb5lB2xeOfzJycFfKY1Elvx28WLJLdmAqP5MZxEwjZ5M6Wj6jGDjwBavsLj+ph
BNwDHnV1zKluhPfo5KmkoAXaP7eygKnWi9fNzfRd5X9RhQ3GEzu1TZ20IfBJYVuw
Bt4IthjpSXNU3CeD/EB5H4MSKoq75VEXGsHM1nMwbDV6jd5Kwmb7OtM6YFNELyIV
zhMkrDHkJQOWWCTW1ZLyugPFDs/dyZiCiKdZj0rLuo636LmylGL/PvIyhyDJe3/+
GVCc7pzrHtMmCcT6sTlEJIK6IUMxjKgMqMoXphJhmrG1/R6O5gtv3GJp6PC39x//
mU+0KNP9CKZaGzx9wF2W6WeLoBoMDWjT0MyHHsVW778hvD06fzSRHE0cG6MsHwfe
cW46nMlR14MK2yqNePY8VuWELeOrsv1Gwbn5aK0euQMxqrwpbK8teCbF99BkUuIu
xzej0HtXXdv4j5kDzkE29XA7SgcRy0fBHn6B0hVjvHxLQfm8f0AOr56Vy8+1Vt1n
QoB+TC3vqqFXkPctvw1NsLharfDaaxzTj0sU/ORGKfqvJwpkkOj7n68v3E1/AWTF
n8tEJT0ZcOPhqTKgaItAucJtDPLEqeXKJx7KWXX39ogqWv71AjMgP00YY13D4v7z
O/h+dLfL1Y7zMieGkiL1NdyJ2WgfWDgmxmWPPYm8vJ6jPZOWoeDmovgZfajGk0Ml
x7vytpSta2gUOXUjZb3oV4TboN/JPdWoIOK2EZlJybR/0QzuB2nXZRAYVJRgy3Fk
to0cOiLdlzVQblgz5vnwbpfQipTmC8Yma3k4WInpN/JvglmyeTIlkIEnwqvBZgVA
dtmFQ9IoAsuMY4jCqRv+oblCgWIVOyWBZeIfuUbTxqZM1rwrgWilv4cHbmADpM59
S/DDhQgX2lZ3Z2O+lm00ygOIIQrfI9/RrjbiV7YfAeOpaL2eJeTb8caqC4D7jroz
joQlHdWGufSjwCMUbuCX0Pmko5SPfEneRBgkfvxIdoU16UOPA6iW7tTzkG/+pnbX
NbkGkevAYr6NieAUNLZ+eLCYP8VTqcqN6+m68q9sdhooAKlNqZH5bWOgg48ESWgN
W1IK/eflbzCzDG2OI2kxu7fML3oUA8EyE8LDU5GKPtmvSkzyuIMqPtgDQXKpW5Bl
UHMMiR4r++Fe2toqEXFPGd/aCwu3u9PKVPeuQzEH1QsrQUid69ycd2J5tmA7/Wf+
2a1s+m3ePIEU7n2GmHoZffNm4mFDdTAQu6dQvX8EflZcSYWjR5/RZpN4RIHBLBJp
q+MBqyMqgRPxwwiZ60fftttBjrzOZCxDqirwfGavalaZ0Jo8e5zGgYEv6Uzm4aEj
X9JXUeCzi5/6vyJNZKcpxFkQgAB9E9zQMmc4j8mvNX2xPBCtuFRCjhH7lA6ABFiO
SW9wNFkc9wFiswD5aDiPyQclZob1NxnUyPw2h5dY7rsMrmY0QcImWLXBUksSnu6L
VXYgOo5BLkC82GHr/quLlNBbgDY3sKwxS+KXGI6CQwVywXU4phCxKIVBB6XRhMaR
AT9vgu1w0yDBaXVkQN/XYpzjOai4f9j+bi0uE4K00LPcLrBpJU+7CDejxzRNNi+L
T+20Mk4zBnti6aYEdejFW6LkPRozSDB805wIMSxkCsaB3asWcdc3MmurGZfqRkdQ
T3qQhZ8RIAkxNI1AanfZPqJMdS1CzcDX8iuZaVE7mlEy2VE7G+lOwRS5mP1B7jAK
Cni/4Q1+nVbxjDLg4rxxcF5f+0E+pL/g8x4Hkqt7O+se70uTxdjiVORpUD+aJtN5
ZdkME+sduAN21jKmwA3qCYIulrDr2hQsANL4L5P4TWIfB7uFIr5cs5awQo4jDRBV
O2bjC/aIy+2MSSZUnrkgJZXul8hJdewqJ178NJdDYtxey26pjlfwmsEwBIi+Fdq2
Hv1AFgVZUfx/R1LewX0QS46WhZWdfedtZ7eslYfEw/AD9qwU84RS+806qKQYFUgc
qwzBt+Q10SFvEcnFsFK+twHFvQU1bxGF4QT7X0VjS9dFgNgAOzDzEIrWFmJqep8Z
Ba29eWNB3tuTt80qBVC6n4Xnc1E7Gu2nE1u/HFPXDU2XZOPN47JfVgDTyiW1icgT
1c+zVXBv4xB5OplUEQ8szBmQzoymwNxk+teHF7ReMa0TK5d5xhATJ+uH5hsH5Iok
uLaIsiUsi4+vWUfR93wkWoXKAA8oe+pDsfQa37seI5EK05ZZnvKBoilrs20INQaC
cVL+TDYglsML6BbwE1NebwspExy9aVvF6LEJwncpZW6uqp/I/czJgAudU2XZv8bG
Ze1QKgokA7WUtcx0xGnBRZZL5sOchacRoiC2Xd+Z7sgxlvVVBmvtSxPiKUahNdAg
KLhTwGHCDInwZnzdllxjWcQjcaKKvIRTS8t/J3zyIfd4rqdOMEtVx4d5RB6KcSgp
JLZULYg18HOne5TbNbT4sHIRf9lwXY7wVy4yUORSKDEv6aTi54BtbqYna+1QQ/be
+lOKB1o/OltyNrOAJ03ni9Q6JXFjsPUQl/jADjiD8Cd/fznBJU4xZ8bKgH83o2bg
xX6Hhg/Th+Jg8sBPQV2pF8puCm9dQ5gxosqTsN2fGLRkSXGcPHkyfJTG6fRfNNsT
c71HJAdyw2J8WnQW76AkWmkrLgN/ay134HWqV/hyJywH3pOTivUMhSWw3q5sH3x2
bpcbRF1dCWMaBIM6ZMbA/tqisb1Bp0+wpJIXyz1dELayp2PgbgtcoHZAu4NdD4RF
veoHuWKj7StqL7V2xJIEPK3NSOGAzuVSL2d2dtwzUxiYHOT12r1pGVnY5zojI9Ul
Tbnzs3t8E6RLQf6BXZWHtfyenZxQqjmXh8eH4jzSLIvyHvw3iBIqyFeckd+BAYKn
RUw2nimt3DN7FzM4daOSjel/Kf+XzJY/GRTvoBqIDsPxIwVCkLVs4XW3zdr14Wnh
QGf+m1e4b7CRDznl01PyJ3KY3pbOdtsKWesFcFhyTQ0dWJSpyPr65qCRbWsvpUzD
5tIC49yn0E77ggYWEkDYvP0h01zWQ5liANKKynUMFaDCWjPxzHkZC4rv/FAYp4sS
BTNHKVydD7aUvWDzcq3xawZRhhmmwfApcJ0yz/rCGme2UXP8BSHYsL/lkv0K4E+T
VUV0vrJcfJgI5GTCEGN3GKIjoF3BuieHRHF2C0kq4AP1tYVix7s5M6dhbVMff/yC
ZS3OCgpnoE2H51XHZPfW7R8nHCNDvyX3m5h5bBZKQyp0M9nyAbONbD3bNReD7qre
U7AQD4M8vfCH8riSHdfhbp5pLBPzN1sDZZBC4yFtRvT7xDlE80HfBW2PQ41LrVP4
UG4UNN8TLSmuYmD76Z4qEq9ieqkeNWE6lGbsgtJ6QU17Ocjdp4FU/gzOMQR3og6z
e+VSGOrB/ERzzaDxcuLrqL02wk+S2oNYsySFoAHknC3Lhi6auekI/mRlEHC5ol4h
RSlTJBTqDzRkASYxNwU5PthnQfQ3kR8Pbkdr7w57COf1ISoIIR8mhN58PVkjt8Hh
X3VVpFe17dmIwa+cOIHyYRl4ZVtPIo0WJyUC6gjXKermKPPQGDDsODgOSDg5ncXK
Nf9VHjh477PGe3p5FrEjwx3AwzWkcdv53HPOQXbGFtU1njg4PtoASGuXpYcYNj7R
lRFwiJ2vz0cItv39NYnDWXU6Tcv3KrmRBFSFNBHQdwgNDuc2votHAA7+DOX9S7rl
bKJ4ZNZOqkOg7I3SwqEya64k46CK4d6442H6SEqx3w/hcyAB7d7LhQjMBMaiUp45
BhYbTG5u0cQfi+my3edDkpeZMuumuj2JkhphD2IQ9jObOsP36nIerwTqpNRyfzrH
3+9quNwkc5IGQ5MRZ/BRq+zmPLbNhzOLn1kI0CHqKM++/9yFckCnC2Icwxki5d0g
TEi8eUvouNZOztkoMNeZjKzNcWUvuf54NqPmf/vI4YgvHtlLsSQc5IqdIQl3ycLI
JSLod7GJ/Uy9ENzO8CHMGf9DNXa7LGWI9/61StUewOOtDlKne8Mm4B0jqs3WmnOt
OBIArGsm7UfvUczNPRUFcqR8RXb0UXD+rlobuPfDEwAXQmcvu5myP543Lh2Xiaad
IxH3PA29G3paBJpIQfDgjaZz5Dz/HT4VdrsS+fhpmtC6xtgAW4/cvtRgp2QkU0Gg
rBobjl3JOWewudZahXeyVuT+H/9JCRGRyQDuKAjdXhSiT6l8/t91LWNT48/ag9A1
Ti2MQQ5BKAB+AVoBXCvgGdFDTNAjD45ZsOtBcij9zatYC2i4S93ChRMTtXil6bj4
mGRzEVDL/2hT6OGFBpdoxz5n2zZ/Ry8Zvny0Cu+Kd1zN3yUuFL5tR6A/vNe52QwY
2czSS9GU4TEoflTWm8sjRzxZymoZMDSXJWw1+8/GnRGM+nzK2EecyhU3WJ4JfUFy
kSShSCrLhLb/ysEcdlAnOv5pDeAI6JAi3cfJj06g65580cQnSeSopb3O228qn/Dt
e1QH2savt6GQGrPhaz6MabBkV7zdJhArvo1wEgIJzRIFLzUfeTTfKi7YCACZj18d
y0TbHOjMvpTpTfbCFj0gf8iRWbIoXLMfGvtvohqxmgeshnwjH2HA6CDDvDFFKmvx
X/E4aJbxQnB/6/8xOwRoGDR6rdmDKTlD4KPGWPu5YXRmnVWeWuY93wUX3JtG3k3y
V1T5hYTDNk3SBvgqzGWBNe73TeQGKiLuZnjzdj4mEqM+3F7jbBzQG6MSqR2kOczf
f5dNBVZILZTjPvcIo/K0LFlYch8CzbsbtR2idswcSNzktErNesk/ibhCeoqNScfu
g4QhS+xyQBubceK6Wm2P8pU8x62ip7J3JenYui/8l+T63VBGKVVh70CYK0uVxIis
srdmsgyXIpfghMK17Q4cPkmzObJ5YPeu+jrRpltP588k3FmCtabQFGbhE/2qvFyL
wq7D2WDugfxBy8pYs9uRJ7C8trujXG/m1XjSVjr8LHeg7zQkDnVN9m2jB2zFUktZ
TU3Y8HZo5TkI3OQ/aBixzr9iW3UanyawnPYGZx4GV2Q3O6IRUJtWWygT+YLutBjW
iv8MwaEazJn8Ui8aMwlvAc4Wn0b4q9Ly53wCdHMLpNd0GFU8sHOJzIIj96zYJDPs
it42NV5EsTzVZJRxoQubo+d1xO3ZRHN0jKnqzHZtbXB7nebWomiO3a9qzKnp5rCy
+ub/tQL0kv5tO4WKMLRetyw1PZiJ1qBcyLZ+15GtKvLQPTmofBa/NYOklK/aV5NB
Dgu9Cq4wH9Cisc/Uux3vQvCqib7WhS/KfpDnEx5mB8dgunpjNPwGglGk7MW8Mg3F
/pIfN3oh7HdurYRPojPjd1TAl3NPCUPkaDM7r5zQRweJjCh8CDNcsqfk8OFg+u7n
LuBpclmUDfrgIkG3uKRp8fHSlhvIgcilCCLbHeF54lSzYBRIg83alvWn0QYI+BjO
cuJn29DCDMMDsJhTM+MqYtC0/mS6oyLpXTOIff4t0wgWUC6NNJIQ0KswjV51WWak
8BtMRNJPo3EPUCNjXYeC2ceJBy+UaPHR6X2tt1djOzuPqjgGOAb5MRV5j60OKe36
cf2Mr/mYYmaVXOfB/kHtaUaEiOVPvaS8+gMhpOwtle+9A4GFM9sltPxmE4oxOXbY
kOPZykYJ9ylNqUHYSK+Y2Ry19azXXQx0lYD9CzHIrdO1i0gX6NwaBn4cqS6nPRn4
jTrvz4JXNjGtjmARSb40zUNX3vJlYBnv3i6ZmuyC9zoIpuO11BRhjILYblkSMGQx
HgdSorRb6eufT9Tarx3qwjalPYqicBkIO94o0+ub2WZAdlimbMvwdFuEoBvtqHxj
CYIqodGEaIpEs69Tmeyekzu+cOVu5EmcUYHS1SVko67+Bmka8A5WsDWHjPWynXFk
yTlqGSUhXdkauA8MryTCgRKhBZkoDzQyBl4VWiXatbWzFWBfprtHaisPaftaJ39A
iI5FcN9K9iJ4WIunKT9vcUlNtTDqEHtAby415SlMdOPUoyPBtAxEExnFsIyb1qhI
5rP/fA3bBwueNMoxnSaM9DeMuYZjpwHIzZuI4i4kA3P/DrhCbVpa9Y0hJaKdI+qz
cClT6LaJHY7p7xZmXATyPy5pgiHL9g7F7EujwOVFfrxX3HnZFOpan2LefmPkCCOa
n2osqzlqhCHRaE7FoDGVFracGEO4Jm21ONkOzJfbkCx8nnHgKclm5XG3NcGzqtLj
xllBXIsLuX9KbjpZeyL3iH2nmwSdFDGd21/fGFkoW3vzq5EEQZe9VGO10yV/WUEL
Dp8g2y5pclzWC/KzGI6wJAN6Hf++28iKkrcVGRfqG9kF2hjUgoemOfCLFhm7qVaw
tcXADrRf36lo6rtX8gVNIa95VkMAEfWljPkkAyD/vOe4lBZMBxWoVHeqdmho6QzN
6FMD/SY7gFSeAnXgJsUDq8EoPapM4LV2/G0fBPtJWwEbrwON7HdTY4yVAm7korq2
i8WnImhIljDN0M+S/1xjQFRk4NeaNUGeZMP3a6JbPNnW/FH2mKBoB2dw8t1CtCV7
IntN+CjPzPNDGEftV+h/bWgI1h3/Myhavyz6KLGfpxmyKXqhgnQH0ow74/d+vaWn
tEpeP3L1VuHkG5XlIfQ9rGrpPHpFLZSCexyS6x9DVoTmWF2LHUV4J8wtLpWQ0pPT
wQo1X4RlQHDx0sodEOSa6cXoAmOcmvll20PPIwotEnpDVRLF6b2qy9fcj62xih1i
IPtSmXJZlo2U5ZVwxbyXrx0SjaRqQSBUyquWfs4MA2/3nLvlzDXdjxRFZBvUTm2w
auwRB4PF9XHO2cPQg1/hLe/JazpQsR3ZeLv9k/LJlGzYc7ISqByLV7gey5T0/EtW
GXqVRIouxNNMKl1cUJMhseKR1J9/T2GEVVUhIIG0WRhF/rUtG+T0fcaHdwSswrSl
E1gogZvifg9TLfCZZoZ0asLG5JwXsda6nRWcHj4UtG7PIwMG8PVgu87QOKtqCMe3
WuIGnZb9z6kyldHTuPXFB6C9VtSoQQ5Gz6mVEPj7YI+dVi+LdKNYkMKM+nsKcbLq
agOpchbpsDoXwW1JhDolOVymCyJKNhGsIGYPzuosZ8WwT7cyoUYTGRysTO328d7G
W/C+9uoYbo2adZbIk40WKv3WWlH+cDwm1Ji43yIEiBHn2mGzw7bBSyfMybjyAf5S
VL+3pue3CUbR394fgANHkiJ1UZf3mc6il+PSqecSWb609SClaN1abH7rOk2Krl7D
VGxDkLaD7fGPWQQfpID4vT3TVdAytcX/g3dsUSMMRAOlXH/8tQ6SPK4Qxqoy7qQb
fwRyOlRp5dywxLlAV5DP7/XnKf6gjUXvw8b/8NLYz5esm2Os5is2w54Vjij4GohZ
XsTQ4ZCghGd4IHmLSBNMoFlcgHRJivHdo4JLncq9ckX3bdazEA7FoYj3H2upPUdd
bKhTB4gpAM8AqCi1FauwbglsR0JYtREp7LZzFSJbZmWBmE1hlLWr/9spfn3Vhbom
xxGy+H3viOJE4IQBJgRZ2ntNXQKCIKjxqJDQ+ordcb1PGuGggWS17EcxbjEw+qsT
Y7UPtqPpX4NO+yMVpW3IacMwSvHXePT6dbeZF138wWINg6vBVHQeK79GYMl8Jdyq
cLFYYNVRhIMnCfM2i8mFYhMjLMwG0VwB7vuxq70dU9JFlXQ1RPPMOCj0P+XNQSwD
gYTAVHY4TrsMI2IizudlEyZ++SGOpr/AZFW/VyzUWOH8lN8ALTIrRL5bAUCA2CfV
mCzozvf6pRBQoCNoN4aCLBKTFPBAJ7WwBFi3IZ1ow3pE03rv6NoJaylr3R2hxgUm
8N9NMKeOg4Di+Qk+FFnEVYqZd+DrpThkVh0KfUSWVL2QoPkJLVpvPJ6cGxYqqO4c
831T7ojd66Z1WXHZ9t448Uw8eSvAb3TGl2AuQbiZ0y9rrrRVithlaEYWivTQ5TCw
tUIje3VU+isd+uHVpO8G+E7Fzdj1+FN9bBM8+CGMZWK2h5eLpxOw+IJpXYd7Wb9B
Q8SgZKsXDY5/9k9zp12Em4zLnDckYHCzp2cQkjlPri/kpXULp7/CAT6WomnDJJlO
N2kaFH4C1rJ2V2tLWJEvFEtsLkA1lwwMIcSnt9Ocxv5sKrqjaX0DhOFY4VVO/Vux
lxL264b2iMCsy9VfYm7M0cA9ooAxJd5xRouNVUYfSRIk+7H8u/61x8GBEqbBGJRL
zY4jd4hUYDgsVHtqPcz2zkFTcJg5VGrHKQHFMwiVmO7BHm0Yqd9Op0U23hESPifh
Iofh107CZagQc6EKuB0gQ9dBAd2UvouYfTqG8oqR/PHsRRgec2vbdNkIilvFLyyc
abnYsHS1Gjd768azvYjFY3ZBr85uMEgaOKfParkE8p9qd5+KFqNuOXRF+DiO0onY
DIHQbGy4+JpAT1MWLTmfcvlhOVv+wjnZGyXFyq9mtJ4ZSUz8ThuLNk6mxYzHAGN0
fjsdx8kwL5SmjXfR5PHgPbf6nhTIsQr9VXI1TLcBHoyx8ZEpLNnYH0YXCDfIdE7m
sQwOSI9EmBwyzBowJhMjkXtEf4FyIKyFOBLbdonGqImmUarDHD9gK4/m36T6nqAw
t+27uzjpxhTzOiUhnWlNe+3HOgtf7p7WWIdVO9Zern0JNXBVyrbdVSqEZua5zGDz
ElDvINLvT7IkHVotd5pcEmBEmyskDw6vq+Avh7eVPVuwOwFWX18nRqlYO8QKdbTc
9Iad9qUdge89eww7X+l251zBI3lEz0QdgkupQ3xPQcMSRb45HBn5K0Gd4kIDd5JL
FQ6ldVjJQ3DpAzrrwIitGGGerzCLrUDx/EcfknaFrCORM93hYnBqsedfrCFk0aqA
wUNFk82b95F/T7O3YFh4sYidTgRHeIJkR9F8DDu3xBOWLQp/pUi8D0CTNHUEGqXe
Dc9A/hBOZxrvEQnge8cxRinReb1uTaNrfXh58NSXIUrlbJ+eXGtSDN8yHgVTTTfa
3/MR4ak2GJarl2L26ppExWufuZFnCIb50O+7YdXKHlI8LXksu5RN1UMiltczOkB0
UL5uYUGL/PwOkQJO2PvusucdC0wyi0rpUwFioycWCLa3PB2Ha+hq/Lh7FMcPKALX
ZKH9tH+ZH+ekp6TxKLvG8DUAfuTWJDLTsw2ExlPEXdu+2cf58HpJNYSU67Lb8N60
mmKS2KPq345a6CwlbqdwTdnVOFZkU9OYWRVx2eTxXITNHyqKskEqrHQi2ynebd8e
YCM5A3SD179gV7uIcveK9Wp9V/yzuYBoDgG+sbWBQd1Un73G4yQq2wIxFxh+QDlb
5/TPyQrl1RvX7zaMEHoi1ghobfCb+bl6JZ1UGHB2dtgH4cbzSSgrhxUnDNBqm/SD
8Q6NpqjO04m2yyaCwDmHpp1u0jAxls0m0TceJ2h3b5HAexnYIm6M8FbgSaB8a7fR
iGOAuQK4UabhG6vVMuP7mqJFQnBeyi/s7x31cMq67t23LU+y1v/ysIdARHrzDDNL
2pskBWCQ8dVJlFstFmLldA4gd+28FklnTiwwD1Bipc23ttEPr+iSTcr8AecFfPHU
i+Neq9TiHJgT5IGqpCKa0ChehChJvvT0XTcFiAMiMPIJt2lN5NK13VN5BhW3a2Vx
5rQBgVH7c26OrVbBtRE42MK1y/BApvThzzKoFyleFwwy5bPZ4EuW9cOYnwm2vefB
o+Qo2+j6Eb7sWdsDlxDTH4Zz+YzxKZTaVwKARU7aRpO2EN00NyMx8aqBc9xldlJ7
Rwkw3lHjkEPmEFZZ3nkEJyNtDFskG7/MJHbfEO4mwIkudEU4qyERY6Nb6ovug15/
n/+2lqDSEjcUFP4d4veqBNc4IbtdjbPE/qG+GhdpvnNI25s6fXUudLoFS6RJRG8i
DK1aM+40i1v+6XKsTNb6dBeZpQGCNTlhzk8/5M3hKMzGq3n7Eh49vX966ZidUm1Z
HU21w2ZSMD1tRMoKmp4U6px4ZyiaKu5bD6sLgo1E8dk8JEETZ3L9+2d/fN/jaH6d
tvX1aic/XsccwXMe9sTTz+8W7JpitbVAJsOyKXFbcZM7Q+iBrOsfR/5e+uEdEcWK
Y8srJIJ+Bu2C05yHsARC8tAT0GycmeyRS3+tKEvO8wWaDoexl3jv0iTmY14fbppp
wUm6tDctLnoZSmeSkciCqwrYRMUE+F4x0TawNvobvg/A34pw9Q9xS+lolVdRS3nl
RgcjAvBNt5r0VQbVpgxVAUIBf0AFPpaFYZRCRMHYgjbFpc+4FRSxt+/uMYOQv6wz
lPITHqadC9cGKheFbsGP0fwb+DyY8XAMNDen4mg0iOLpXO6z/KGEiTNnrQ2FYOMt
vj/OEnW2rbmeXEyapnulCHqFTMkQ8UA24S2yX+VlM7Pcth+p84EHciru/JY0zSOY
N0hLPMh/TyvN/mjbPT21HjfXV7q9QN7OJSKxx0Lg6KVVs9ch7zXA0Dag67YRZD9c
MVKGLiI7MkGarXy5x8zvQkt/sp/ysaD/NoR0ycuOO0IZV++uyiScss3mSDcU9yvD
KEg9YCm+N/ZIP1QRFvfcWHd5TL3+DpijS/KiCIn73gfF2tTU8xRGGqRXAww2Ri3a
K1BmvWtGizEWLfmhV0LcL2MUrkmg9mQwfspsR1KuvuFF7LJIKR5Xe5iu7VhNzgE4
QQisgFyMn7zsProD43nMr0TTt6+qYeEBsQlojsbejSBDCZTTZ1aov+PVFPtfJHCI
4IXgAcSeAm/20S1zU234qgbUmCQtobRHCfg45S8dAb9ofldUGbzQ8fjyflBucrU6
1f+8lCbC9E1CT8B8fHUZcMktbPSbMlPtjDXX3FwEosAirFJaJVEuBQLiipywAv2H
Nd3HnTuDSfjVoQ/Ecuw5UfSl1X8ICoy7T/c2Ys+v3HuL1Y3HJSQKVf4QehbpdG3O
+APtk0JlDia11wi0+g9HF3gs7xZh4tHqH+VjckEhnNhL2JTsF82u6FM+sLEQKJ/E
G3XjWOjzg5MKgwnzJ7koChQ8nNr4VPKf+G5mGYmEBXRHtOpTDHi/87169h3jPEzP
spLBjPQwYtJkVDxPLLV4wSBV7RE53ag4+uKPZqNg7izDLA88nnlGmaZk3tFMYes/
+vLzhosLb5X+nCh/RQraXAUvbRRWi1UlLHPHu4GYvBNlGuU0Ke4tuLl5V3q84J3u
QjTDALcLpkWSZe6gJ5pxOy6mnnuIrVPOo4GLrzn8UgeqPuJSDG/UwMn+9GC/Rtn7
PaYOFfgVEAHrziMN0CV5WjpUuK4LIZuXsQwELCHEGHTx9oejxpGKQyPp8HeNa0/b
5TCYk0tCQ+QGAQjOETqVeTiR3RCiyurxu8jugHuUUc20EJSMLvyk1YvOrVrw+kq/
wFdIqMtrmX0T3WmX4BInxNFoT/LiPRDm6iSu53DvH+arxQcvh9KOznw5gmpWUl+S
SKzyqYkYt4bm1GWkCmvBvxid7IlQMJl7TNL6b6/XNE+2zOLJ+7JaKoHoboWeK407
XnrpV6gYA5RGItUC48h88VerzV5f52pxIIpPBnVauBvhNwTu55/3tG/mRbxaVIya
K6XLJU1ONIE+5BFWLQuiI7inb7G3mZYCPUMGJUzil2HFwr2KAGeiHg/cqWnfc3bN
kyO7s+IJ6xEhTo/ssECeRtNIhbiCBhniT5v7WhB40yRPhXekLIHdftsToKM9xugQ
OWTEs5s/TrcFkjKjF2ZSKtIqd7CPvy5Fyp34lyPAlbv15+hl9ME3a6Yo1SsAjaRj
4SmFiZAz0mEqn4uuHT6Ox4pxhyzjhJA6i+nmBeyhKdFkp6+hxjqHpsE06TIKfhIk
0T90IuI8sQqAdEx/0QUCpQm6vRRQsrrZibA5KkTwvNFqESW11Fkx+TDvVgL4M0oJ
jG9LzhNKhg3NQngBl455RKd0c0JWeN6Pf5wZT6Gqfcj27jENkQHChi6xVsViba8D
Zx10E9d3YKSBflCghKHinWi0gYF43CohDfz/nKZU7NGVf/l8NZNlLNyJuwG86K8f
O+fLney2N/tkYnHhEH43WAtZkfOBag5LyxrNQQzPoKip/+n7p48IoKfJqPW8u75C
dwrMTJfQtT1JOvdC+WfGF+7MmKOgr5SolRNLotwiIKbx7WRMBxQGhz0Abrx6sDNb
w5/zA4ueQ/0U8l7H6yYXPoOBHJ8laMXEqMNwid7hbOJ0lZQpzkDvC/XrN/99j+1B
LmBpfs7wzEAFXfny3jC2Quo1FbIK87a+n6QTZ6uEqOAh/f05y0VydvNaseCfH4j7
8sgtk/VI50qeA5RMErAprPzmH4ikJkpDJR5D7/+IxqHCO3xMyf9Wa490xJT5Mkg6
2jyd52XzyVv8Af6+3JSLNCVbTfM09Ho7QD3C2FNqHB0z4li2tPg40u88RxEMQifV
QpxtJHKNy7IRA6onmAt+rZmAwTKWC5pqXgTrKfySYxyVt125NKiIuZExGrygqzqB
ntRRKplf43o/oAOC2cIyDhQwqt0KGLxv1jZATsxRWpDKpN+cq0hOMrOFvtOG7vrT
ZIGUn07KaUZVZ8Iw1KybpY+uvhlSFr+42N8enKjuyzNjUEmO1efnGorgMvcisuXa
z19eQ5tniV/taPL0Dzk5hPMwaqGTzPAWapMn/ZzwhyHd+hIvHPhD7Pv/0RKRBALJ
+ihDJN6JPS3WMqOfexDp0U0irYCG1T4BS3mSymCpsxhME6mLXbpeJhMJrL5tEjPR
r0k2QBr0xssvESoHlHYBpSbj2K8HntwtX9qfGQ5Aa06omPdPuDOG+hvMstGsiYRD
9ib14m7YsL7pAroDdBNnq6TUguBYu7M88lj47SjVfWw5Rp1sCR+72NQIG1YSzLZH
4zm7PQ4Gu9JpIAp5xTMcWrIi2mA3Ru4SNqAUkw0fztNXppZMQ6ZJ03dwz/N0otUQ
+LEgW0TTLMH3+gncN018X+oU/4odCc+1clAFWfVZT/kfDo8ethKgrXwFZ1LpEu5o
8BHdUA//NQMgjSkB0Y6brEM4+4Te+9Dv3YxsFHUTnswB8FQLJ6GRUDHJh8Kv7FnK
UXr+h6Wz0x8NrObKGPMV1KD0uRRhHM3svipVVWElUzCh3JGdfEkn0ZHsdMRADz9u
ZhNszlSQFF3s+t4D1o6fC6DJAqvP9dZTH5ATPTrpcDDJD/NVPsaRhxD6R0herKa3
/HgXTV4bmLeaj2PzoDSnwlfqHeAkFifqqn707KgnWudgXTKJ4z0ZaiAoAxrJ1PWu
LY18JLqqtuAM8iSYjoXMgNjjtpIiyjP3wcMNiXQcymth0Fgd6aVFliLTDffoe+8Z
pbMWAS1hxnemLCySaZrTf8crWyGWtVjRgghynfcyJ5Ra0t36eApikqr0owatHzFW
pNMF0pCEpxDX3uidY9ln2DxkRIZNHKftA4rXzZBtnGhTrM1kpfw334S3uJLwbi8m
ClwrpNPW4UgnB/9guO7J9YJ+23he5jR8U72sO6RpI0MjKEP7Zs/TjeepNexay+6Q
rY0tNmf55X40bH/0YLBG3RG7GcbovqsZZtHevU1i+FGUj2v4MPVc+cisII2o324B
sKO31mspehCMsuFHlvOPUJg7K1pP0P5rrEYoWrPl41lDoO1LLoKr4RT+BXlijvfI
VulBfxQIYqHTrQYwiMBmMMumDfajsqQVYZs61BzQBrW6sueufnNxERQ+UJJ5IQnP
qbXB8EVD6t5OjPq1GMLZGjoJe+ePi974gZLEo8UG0Fpr7tTdWRaQbyK8SYq0kAfl
AVLWPfb30OmpPWIWXJhdJy5kCQfakYMnHZli2p4mE4Msc2xYQM0l+L9qU+LKRub1
wBlO33vjnNPwDJPk1+2d2q7JB4zClwaoSTgfSJHJ9xpmp7/Ez17HOv5HB80A7kqG
DWR0/OZnq/e2GJzUCLNFFFFkPjbI2nkghgLgJGKYAfNm7ssaepgGLKgToibXoyRI
R3FjpIsLZYfrIApmUg9F4NoV3VA0TjwXRblWeS0qkbJbkA4a9inlYjSiXlVJ9ZgT
8FJ68BgQh3y4ATEJwKJU+2ePCUnUDkc//+ZOh9Ic6e/UFn71lzs3MTaq0bonYv3p
wWteVMhRSFeFmFlB3MxG4tjwWR6GCu24345/HS2jsqk1SxBnr9pdRAHSbiUvtlrB
dAODHDm6hQi33sxKlnG6SADMu0PJGHKBXz2/D4O5noZBA7dMjze5DzK+GzHP0b9n
VQAU9zzJYcO21OFMURGChJOr22Aea9QeL5WOOsq/suU5kvDrPzndNAXXeOBmsyRK
lpz6M8rSiR2/j2eO/zeXgVOc6CSK0XwfisHwYeEPyxrpHyd0XYdCiU1RCJhUT3n2
NmCVlN52TVm+BoVg1cbV03kdk6uI+7QFm12fHQGWOCOrkVb0NfcxC+gi3odoYBvn
KpYClP3C17gIoenUuh+hDSp4C3w2Pzfcs0DO2sbqtO4nu2yWjzTXSZCPQyGvzNhc
o7s1xTcEZ8uOnAzMzsmPQb0qnBUUlA1tdxMZDbofMTcmihPSJ5HojqTrBuZOMuvI
Jv95ZHa8u53UukwrpQPE6GrvYyubh7N7nqNk46pcGmrLw1NlIYguqP9ZosXvT6Hj
+L0KKOTVBVNQ0C+Ja1nkcuJjYb56zOUM3rH8hz50hv/u27F+dnvS6gf9kHZav+gs
vjZzl5XaGJE18K9ACC1Sz3gamzrErp6mw2XG8nKp44wus4dxfEsft0Kdtklm9zhk
0m4Rs/ZYvqevaSqTcwbwKe4VqbF5WUuMsL9LcQTgS/xL91iHmfxjxifvjuGS62nx
5b0KCQow56XNECfEEyrllH8KRynviS6nEZLX+iFPJj9RpaeMk75/dMDrdsJPwh17
pCSVhm9mWT3JZ947QrPDboxNktft1q/8BtxbanbF+CFgb1vkmWxEAYvnT0K6/z86
AwfUbgr3nq3LfDr4QX69JbxTqzV0sEaFDvv4nb2RMVf7Hox6Uo2CqLvoHuPxEEQa
KUepEVvtk7gjEdtwsmrwaZvchJjjHCv8It9qaY1Ce8J7Z5bc9ifSlWudy93hXZCh
XguztI94rXKxtVnhFDd1LlvfLnQu9gWF9Y4W6lJGXSkipVyOGIJTPAVhLwsdHd/d
p+THg+ayRodqcnt1/LoTwxJKAqAg+SQoQbg2baquTa4At/kRdZftgHEpya+3vxd5
p4kGFDewWPtpY/+x2EO+oVsPc12SWbd1L0JsbBrkD1EimTpTm1EB+bmsCVEpiND4
LaJr4NNMv5hdPC3WV8h81XOwJXhjx6gcDrWKakNbBbS46eUylhwW5Hd15Ytx0hB4
3cOvGV6DIVlUMUU6AxBtO6rxFYwrTUxf7i7YUmou1pysO/oymnIPSZ01PvMa6jRj
tTIiIiz8iwSDtskDaQI4tepgSdKBwukh5IspDtlPGkqLE+sQBEkpNGGEmTg/WDHX
tXGEG0xzDhkwpCXOgYFiTnRC49dEPYRy6JlBB+YjFgDIoobBv6Nc3/cIvO+lbrJd
g6qAdhyd1sT5FyQx3kMtWTon6DHR+110XMbSkRSPvvak+ne+uXYQu0gaS3R76gA0
kYSJUaCt3io2ESLqRzJ3DvwlxLHUeNJPzB405YrsRAhqiyLipkpcdcRwgULtL6q7
4LGERK2SnBLEbNOT+cNYt6y6C2azsyvAzbOz8YtmI2TzjvGSYjzFQoFLZGC3CxsN
9WsVlal0n/BehDWrtMRg1VyoYh5o0k2FTcclfqfOjNwDMVs8MaNq2TLsSENrmjSH
GRajqaDc+F6yak1gMgOtHw/cRCS5pvGZx5ReyEePdsywvLWJ2ENAtFQJ3/os7mna
aNOmn8Okh2o8Gp74/6A0no6AttN37XoSmEJrTgAnqvMDDRhXvhLv4W1RTHO4qvWW
WEIUwqZODF/XJ9zgyNFdRhqGB4sQSoulqPJC8W/RlI069mxe8HyuJLMCX2SRrtVT
AHFPsmFrgz0FYbAIKa2W1g9fyexi8CqMLwbWHAm4x7Pt+RSiXBsBt5fC6dJ8b4GR
eQhCPlhJDYAAPQxOdMYpZwIMOkUrXPxddBTEcYQHA3jBZznssVCgnqqP6M+gd7tg
FGVx3Za5eYMkBRqCMvFli9kwxuABxnXDuZyNE6ZNy0cx4OZVoTjl76AUIW03zawK
qtPrg7YYFrqJsCjGzc0vdOezqKEjaCkduh6yUT1P1p/ZcDUKFqEWX33nri1CrsQA
vkwLTP9gt7Z4KVhwPRerf5g5hAJu01Z4jUqGzkSrkMmKyPDy3jneCC4FbP/hNFr4
dPz7u5S0A4g9ESEkoAoOZGtbA099jgbLzMIZrDeuMoyRyMqGhhkRhoRVw6qdDAc1
fb7kUUayeLfkPr7rMyW0zonz/Hwd053ty7gSIPen01kAWPZy2+UNjzIXC4rsKV9T
4sOnd+CXn+0Sfczn/52cXdzOlusIHQXnDZRLPXy+Q9isFD1dD9iYjXIP+qM+Nnns
JSLo2KrPfcBnkJeQhZwV6ymWNNRNbEhEfFUEtVoyt8RMppGaqkLRVMfzX1Q5CJVx
Bzm8a9vSwvofOAzvrP3jr6IVoGups3QCteyldT6idnl7CG4audN8ZxAZGX8FgI1S
mvweUgt8cLFjCmfzpdky6Za5S0ZbTnpqp4HwQyU/Lh+WfXDxTcdjaQPeahIC7/nW
ClkSQ+7Xz5riF57fQKuq5OUgK3CDxymU02/BRTjHL8rGEh1VSAQg/ZfeKPbmkgZw
dNGGpMi38S9fkANVR4NGl1D/KlWhCsTohsf4OWulzVWTY2I9uV2E/3ePWKJM4Pkr
cUig4nDNpNeFhOk2j4VJ/2pm1hHAiR7WjHbLHhXZdIF7BOPOxJQVEm1xILuDH62q
QZGQuYfIT+2q5++yeeUKs+2qEaYRNEHxGHiz5pojd2H7uupraqRJUl9SP43cP+1f
egt5HrZNcBhFyZK/KORK2uhnjFtGCPdfQiBsV/jfkcKx5xIpw/xypa/VJLnXdX3T
/ylhR1c0GeuwI3+/QQcfiBwWKSgNoj2+Wz+9WOFMMxH4Gk4dXgmUwRbwKLAVzB+O
cnjCaFBrFVsFoHTtv4c31Jl+aFBKXRBbeEQA/oRVOpkaIKCJ1hKmdCzU6U7ZBdYl
U/5wrbyztpTfmH5mYg7+7Qfg88HuEXFN0/B1jqiLI4+5XsQBn6/D7HJ8UzGUNzUb
xsFCNb7lTwAWUEqhLe+VWkfvwp7MtrRM5Lm4gJxOKzaagM2ePEhyf7jvPxvMn6g1
bnMQ1njt+SjjWhjR0hAADg38lftj9oVzTM84OL3QYWtwh192p7qLvXCZbsg0VWH0
WZ20z+n0uRqVGMpTcqAzpHdSVraAtBPPMmFbuB7ZXPo/hKamwLQo7eu8jD4w8mpF
Q9m12MBXyQpz41wxNWBNmhbyZBsWyWcHrzLQ+rrdVHaepdO6bqHeM7zOr9GTn1UH
lpeDEggd7qt1ZWmkUhiFfDF9iMgiHqhuz8FNEAe+LSgys9hf/FrX2MgqAGI0/Lae
nvhyFkA0R+tukzVPQCTrFOuSkSm4+ixMbcy0e2PHI0S2QQV2pxkBDjMaNK/KpvsP
EGJid6jj69eEvWbSwU+/27aDzQca2PzEh2jklJyK5qX4rjRdVE8LJ3WE/gGnn3kk
e6TxRpUaU3Q2pP3nTFCIAcGGtpPh6drkGypjmIwN2xsPEXsriuKEA/k9+RO0FaPl
xYlJ473fTqAjuMeLq3S4Uy+RghQ7FG5siDmyOLZ0STlAuO3T8aMz2bqhtdNzALQt
xFCR2tOjL14e509r53Px+JByt+5ZMdpXLr9RCCL6GH5kC0ngAhCVznWSta7FSqnp
88QtDDEpsGBcf/hqOSbbNp4LZ5xsLIeqI48ykgRhCrk1Chop0t+mR3RcQWifanuB
UOL7/m28vzOhn1tRFGYRtavxmg8OnePkntnPByxrmA0vFVGQsvELirn2KyUZkwHn
vScd+LrkvvFKeXb8aUh5NMCjcnvzsLfvfEGTUeq8osnE+JY/+b8H69jjmzs+k+vB
czWsnqObnPS7ZmpCVKg3KE3PZlvYUZqwhEdJMxPjN7LyGMMg16dkGRxG3e43t1ff
trgobj7z/nE+kWwAj0l5wkAgabtwrj3BND2tBD6w2G3caOmhLAuZxNcaPdUHwByd
wOthTqLPL2bZzv30pUQ87/xQiF+WY+hiNaygiqRwca+cjXaMl1ljRkYrL9S6qTpL
pph/Nnbl3oboWFWwOI9dx16moCUO5A6nwl9Sqegl3OPEYkguDMichHhYLH8oXoUQ
RLGxVtWwceVRFZG6xNReQaDukQ/LKTwIuXJIV4hzISP3RHI81FsS9VUz5YKOWvc+
u5SKuIp+u2aQiDEWY2+9YbxA3sAD9MJcnKHglqTRFP5EdPYNJ/6vf5SJaix2uUsV
RfhwNPv0ZgVJIBdMYD/5gTuJ+41DgvG2BqGk3Cp0mp0Y8vrGGa7fMsIA4LHqMJvs
0PQzO5rQbLHqyfyMwe3YzgPRtKq39IPZXyWHFHay35NdYf1/cLjr6S76qiJchwr/
LQpjWIax9Vlyw18098fyQoxHveluIYGqlB/loYLlltHQzxtbyFl/Yy9noZKLejVi
4IndHDEr8uI/p1FOXmfp8nhVAF/q3Zj3MSi1vL6fCp9EvyCz10NO1C77UddCih6J
ScbQNW9+owETO2n3t747QKIdmBev9ZuAKCNab41tM7ocIHkpIPmJd7vUOJ57EsOx
SYYKI8wRs/aPyBa6BpItRGapIIPFbBiaO/jOeuiNsq459phLwlAL0Pk1KkJoxCMt
jEJj6NnJ0OaBhTDXzkBTMTzihKiS6SFBksCmoZVpKBd17u7XB3fT4CpJoSfjdmeP
I2AsMZXsi3hkQI0Ru2Y2zZm1m7b3NkDgNykon8yN+GHhgWs6UrnHyfulWIMdfjPg
0b8Gm+tActhbu7MW6W7lmBoKZyW8C55WU5sy++DU0KHtLNdekYrWr8TLFlzc0nQ/
w2bDGQjSVFnVriPKljSoQ0gQ5OxsIw9k7byDJEU/jP1U7NQHboDN3ZgLQHJ8HCvc
vG/M8gtiTKQpCuhUr33Uojj96mS+cBwZcqp3vcYVzkWr5v/yHZcL7xtPOCSp/bJU
gm2DvCjp7GCpfJYEDyFOvXB39YnBAPinEN863doDShzMrm7zNXvDAOdru4e1pBdU
LEry+M9rd/SuFYn8UvUKO/JfXJVyQgEZcnocILBRaVZt30xSDyVxoOeD+tjiG6Xx
dHyEERcLQG6OcwuzJ00cCLHYIO1k8ikuzJbm202lmUMt/srMg2LfGjoRe1htxAxO
1g2fScpyeCYZPMiibXg06M7oyfnpFmA70L+hkVCfT91V5mkbHoVGOpJ3hbVuYU+D
qDTS560Fq0mlZZ6Ki5ixYGOMUwEK7YlUVEW0v7L4oEj65bQXJ9sjm2iUZzCeW7Ah
pqbvEzuacqIrE54WmCWOWCMeDBiF6/9uSAj9XsmvxkKoRzJl53IPfwQpmE9GGrrM
yjOMaxzeiMs26tdNvFiDNbgCatAswN6EsQTwxKOknXCEYKT8+moOECWg5WuL6Ffc
sqs0MQGT65QeZs3VIWbakQo3x9isqSQLYWd1ATRig5/Nr6MoRW1sJ+C4oeVC7+Rp
ZdL1m+Eqm2yMwXziTG+j7s+lOfP6KfhFxMCB6wAb6tvi8AQNJHp6eH1xXAIFVUvG
I9Y9QK0xcUfy3EcttWyheu7rd1FAy1u8nimIVFqchSz++EAokv7heLSht6CXcc23
Toj/6I6KgthKXxgDpkDX8WOJnaKL5JKKMQAvgN+5nK1o2myKIBHUI/1Wqb3llCWp
NGpYtaLsb1PX0fKjqqjQj8XnMWnj3bo4zlmB/XV74v0qQJoyC133CBWjECX/gn0m
hAldQdYLE98yZd41zA3VQu1SGfWNNE3T6FgKzcUOyFqfd/vwZxOsae9uCBIaTEHd
hqZ9MDsPpnFDbEAyv9iEU5Ieq4R233efHS45G7sCJedArmsiqEAfmyRQzJSeM+sM
f1mzT+octksPCwA8ORaB+runN4Cbc7/8KS6Jz9vT0yF/Cmse7+p6HU7mEQIuQpiy
ZOSX9tSZI5SplEJ4qOE7NeeAaPGJuxBzQvXbHmLHzRgbPToBlFBusicqda5uHQKL
uVCzhdWmAsxRC051lqCHvjsbEUTUwkLwzxKw1YtbgpO8j5A/+gPO11O4yigCiA6D
jOQSLuZbzm42mwFZJTahJZqY0VuNAHlHp4rOfd9Sgk/Kqf9IKDatxjsxDTLMZJYh
tOU9UasJttWSFzxgPJjSHjURpJP2aDstBW5OBkQqb/km988xMaHLiWdQjY0LyAWZ
fpppmKFEa2Bgnog298J2ZGrhoEydH8BHCadBVqRmiHEASe2Lyq8bcODKZbwDq49L
a+qIhqDU9/4ciipph2uKp2r+ecOgWe52SFTf74MvNNwuXbAMsqJtaP0DltwFfGYf
AX64M3U+yuKtkG/kyEbdP2jrroZ3Lc1q8BEZtWwU1Z0dMg762oCsHrojn2bMw6fU
/5LPXPqYiuK3PrP6yiSmQuYjAxOHCTeh36gF8Kimnf2LyW9Zw/NSV316gw6U+FX3
LqUVQ+pYyvgoh11rC0m9bZKmqtQFLjO//M/8Bkgi80Mve3bd0IaXrF81ImIG89Db
9QPvjAXBUtKreoBzFY9TDRjNT+xnUzc3u+5NjDNPaGdGvVKCZSDpwq8jj0uQN3U1
cGEqRWw9efrX/4p4Bx7W0ZYWXwJeBWe+BGPkLzSZ1sHixL/oPDUC+e1JP30nmvWk
v7qUvOoNx1wK/RPZLO3Zq63O/DziHQhzIQn96+rmSBL79P7lhlcfNi/+HRpH/aQ3
cTUxoRSFGhxYmefVVPnUebMgOhq8CKBQbtJtddyY36KisxR9QJU7bolVxnGn4T2t
7HVUZ8NRKvU1Iqujst38v6bUCzAdp2GYf1hc+qtOy+ZAxUPYsCsge00IMptJmoku
A0VY3YD0IhX/Dk9QXqKvC4rZD2qKkjIqwcszyXY1TwjEi/TeLL99/waW8ZyZax+3
rc4+RJLmucUVMgpu1KF1Nf2bX1vYt+kTrGbIyTb5Mm+V1QSqdc76UlDu/CY1AjSD
aTPLHWbdbh/lfNmD484Z0SuV0fKMP1ztVvFcruvQX0pdMEv0cq5VE/Bv4lJC/GTy
HaNQeY8rYV466lglxidJU0ll3373lT8beUpiuNHF4Y2Rk5HP6zRjXFUvzp+WJs3i
`protect END_PROTECTED
