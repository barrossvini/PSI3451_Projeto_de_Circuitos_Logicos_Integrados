`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uIv75ZBQeLawEJ6/rstLfSrdNQ0KA4Yqta1bChAm0QdcTjWeX7SsZ45VXFDcmz9f
IqEL2j6JeafU9JlXnLG2+OBHY5OQwlq5cpAWoRNtlEdnuSUzFF04GRRr2Zs7f4og
Djw1YTUaw/gL5G1SoFJGadIkdE/gp1eJP/ut3tFPsfFBTZeuVIzQcSBSN1XtfJ7M
WJVGI1oFKj2fbvvp5lRuTXc7giUs5FVnsMBAE3mgzUZyxvUKZRNLu/CXuOwnRQBb
zLRrKV84nG0B5RALfEEqzIoDggNKb2ijeW74KViQH5/xG4iypq2Af2PBCCfCpCza
H/SvgFk9EIAiDmgMvS/Uca2dbbFEjYj+DfQDx3dmn+Yld/9Y2DxNdtQt15MwKg+I
J7Jc0GNSXqz12pk1iWlJQ4CVlpJJohCviJOumJgu1smd4xgpoCpwSExrb4ica7Pk
fUKE7ByTAsx9zHMhM0r2NcIkxFm18rQeH6/Z/vwMp4DT/RdJGodrPwlqhLboaJJe
39Jf6r7gvJn0Kw9ONaA1kHqf9uS9F4v83Hcil4w89ltChjzi2J6KzECP+q0Xco05
2bDoxkQD4rIOtWENxezG0gtwpNuDcC1k2C8/SRG19hHvpgZ+DDnd0oBa1NExc6gE
rB/7SrWbh+kwfG+mm3cpLqzxhEyg51/fU5bpZTv3tsbjyZ7YsNWgpgpKpeZkf49i
FLfM+qx68HjrGSvFsFSJDIDna9gnq9dUoOTtvfY2foHou6EN6JuNYoh3umaeUV5G
qr3jifMH+pLamHgVXsTEZg==
`protect END_PROTECTED
