`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L2PKXqv7bK02S/ud6AKwMlcxkb6bAgOQNJBjqzabNe74p2R7CjDGYujNu8/jkA/q
izX1v8pr/W/cmWlwKpoZ4Vdg6iTZ9tItxdod3pkA7+dtb/mY/eP8SiLkMZaTthwu
I2Do44bxSqPC4lirmnI7B7zXEkYiOMO1FeRejC/XjiAXYywV7rj5C9hiRymXtKC3
tYL7dg5Tbu9G0VUpbXPEm4LtxVBPK4ufFekwGyWOlHmtaR5acK3CZeITz1THp7u1
E9h7rRA4wxa4m4xF5xhyf3huW4pm4nBO8goXaEzS0h8dtBzsE/ZYcarr7HUO1zSs
Q9I1sR5wbm0oYAzNQRNpF0Ya/21863Xl4TDWvqIdzApzuAx3F17e48h4MwmuNf02
vj87i+5CzRY1+KrPb6uB2PIZ7G7K8LG6SazBRFTp7mtFGpiPplQb+VYPAfYWnAs6
Z4YEV/pRy/DzyAxVbjAX3GSD+/S2Wsw265uhgkgtRUnFG/WLfXv/7n/XJeMaKNvp
fKA91iYWM9xWhQAfOM1YZh3S2aI6LUAcW8RRTUAJaNybG9X5oAryvRAcAZUk4CTg
1lwIhr8pkd8yi4JuVhrMHvZQ2z8bVd4EfPP+DafhnThxTQ/tnNt/vtTffOCo8xNY
LYvN9Z2zai9TJfbP9rVY41b3o0fQdxGfs5AtiNPi4GyVHt8v+Ic7VfHQH/RA0h/z
H7k+/sb1BlQE49kwQxvGFWDJ4BrRtk4uoOh7TbNaFVCYX32LORK5/D+iFt5/VTo5
H6G27lbSWlB3/1AYqNIdLO0/8g6qjjme+K3hFoZ4vGtK1O8iTWd9hQQjP85G50UU
qcp7h1ThvId4o+aFJk0++P94cswrs1vKwZpRXjtzpy/RFIz+VZvFPdFzK4TUVofL
8xaawYTinMEbqKT7X2Q+/yi9dl0eXbVU3UJlx4E8nCc1Uz7ZE7/x0w88iOJ4rQnJ
ZqYjXwOVgUMThwdKxXRO9rptOdTpj18vNee6/GdxkqqINgC3cgMqGifoxj7BBT3L
xH0e3fsqyWCzFx8w3PEUbd9yChIYNSoww2lMLGZpAsE5W1Ednqj66gV9hJODucUW
SMIdGPFyQhHlqohk1Q7dwAqQ9ACpomY6PNzclXoj0KYHRwIP8YrAqAAiSOpo70M/
5V94+05LmZhPBZm39uwV+trWJ5DUTowXM3/+yUaMnDFYUHrR8NF2hZrZs25cfxpw
Af11UkG7CTNGJTGxB9SZS7R1v6AOS7QiGG02NlN4+SJ8S3SjiAfi7mI12khzhce3
voOXiQ+/PMEEEVjkd7UoNdeq2MwnKFckxfbYJHyhiQvcKbUG1ViNiQTglyqI89+U
Sc5d8Ri1ZUM5m4zz2cwz9ZdxddeylBZD3Va3PFs2zP3ntcS3Andva2gc6JZkQI/G
CQX+MpNEOU67JPafFLCe+tWnmVTOf4D9TwIkwHpbbTGcdyDVvz699/oDQtpO6+ZK
Xadt5rOLtcFYpKIZpVYOlQ==
`protect END_PROTECTED
