`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w4jXj65aYqLm753ulWuRaPZTNQg8AiKcTJSItzC/AIlu6vJGII37HfxQgFnKr12k
VpNqvG3dfK/k1pv+mU/2CxO1Et3KeuBnW2h5T2ftFZ4YwgDje7QLTqGFgckJ+Lrt
qYtnstxSuhoWDsanGHJn8D4MhtsbP/w3MXtwcbhhkXCitdKV1zAfjojPDZzQbtgu
IILHNQSnYTqLTyXUF82uzbcTBI6+t7/YJTn30qQIWck0TQVO6vCNk5HrVLLi83/f
N7WzcdtkI0R8TZNysQByNPgIr29cAfvZOLTlz0Nt7QM0QMxq4GkzsdseA7UEu1+h
QcQ6olLXRBhdOGg18AENXBzshZdYEWA+J5dlUxGIRJ6HiwVa4czJ7D95g3R+1DHd
tF5029I3/FVm/ngTaYzfH+zsxwgpEUvyE64Ny+ZLU3YOlL8q15hm3tHEe0bUAYXl
Xt6LYUgZUT7x+/r4Vc8HueNRCtJi7Ae6ZWzKFyrIKS2A8vs2XO+5e7NCtyNx9Qat
pjRl36bTxNOzmAKQGov3sHKxQVVqYAE8JDaH3+gKKFc3w1lRio0FbyoDlPjexlPz
BjeG0asR777LMYxmrsjJI68Vio8ivQBJ8xXmDsDi3PJWEpqIicgpyg9IrLIUynvv
M7BZpCe1F6pxn58EWHe+XyV+TNTaEXDwzDReL4JJPm1apEd4BoZWj4G6lodtUQJL
6hWP0GGHsge+6QiDrmDXO0ZzOLUSB85EEuC2Q8KQJpBvwwe9CdBiSnbJgpPs8HWN
NIu2QKceemVMr1SLImZJG1fwY1yEq1qdU9ZVAjVOHGhWIADupZ/jnZ3UrsfVGZcw
OEkhnVI4lhoup9zwvcCyhoKXeHDc9vSlRjF6Z28El88UiJNuqeO5xF+8/cKaKj8v
HRpXA3CRFL0G/96uhumIadK+R+iMuVWa9z4v25zCJ3D5VmmwN7kHpOXAp7xX5V1e
fXeEoQTuwTgpuilB9bHFS8V2MSd/IYIwwCaSY1i2Ce9WlBMLLYh3Z6x8yl2kVOBD
4P8HZNUIJJ70FtvUrLom2em0eQG/WEm9g45nC2X+YQLP3IY/HaivsSKG+ASq9yQJ
+NW0xsdkDFxFVtek0nkgVFCMo05uI8Tq9GOMr1edXLzrtbLReQHtWswKFgB88K8B
fKjI9amVNmibeWjgX/QmitWxnb5H2DzvzShxBeauJnj3nd5LiA/gwz1ng4vHlrZm
/L7iaEc/+Rq+sqAbTMve5SlTIFb2m8JTugMEmgdtob0JZqzFXiwMQ4RQ9u19v4EO
vaEcnU4WPDvILRUsBI+oumeembSJ/cC34DMA9zPkj79PG5StmNDUTV0Z2mdhkhcB
bd8FLfAz+nDA/TDNl1jDP0gB/nvjnEiMi2/vKhyovCGK+LK1ldSRHETBj98t6Rpo
9h2tVZcQcRG2Neo6pZL+4z2PzxUIgBtA8wAAm6DfP8TuYb+QtXgjDf8c1/J81qZK
/kKR5ssxCvIOd5pskE7PGHLhsu5TgrrlRKfnmgfTuIQXppzRLdpMy9r7ju+Wlzbm
cA6NH1mFEGeV7+OBACjrEnEKglFMSgmYxC7rSBn6/bknty/lQhg2jLbgAVURAWWm
kA86vo+VmVPAJT8TYCr0B639cl3sOImrafG4yzAvvmy8tfm8w1mIddq1YKLZe/NK
JpRaqzZJhZzDI/bqbVqSUkPFTu/xyRsU8qIjxD9LaIbgw2UK0Jt2mckx6sNdIsvQ
Hwh6pGDEPIQvzF9HJhTTDNtI42alrB6d41iFUtnpPThAxC3sHjZ5LXoQvXXbasq6
okZU46go4Ztbtio9y4RY9SjSDNiBrQvf6aapRToJNWzCqw2cnd79UkidvwuqvptM
49qRBM+x9LtECbBmt0FjVhA1zesmr37ry+SfGLvmy9fNsP9DE1jDbMbXbVuam1mf
ODVkOPv07E3TUpNcHdTDRIyMqFY96U3J/DA9AEQuQ86toUaaNw+z5DXep1C2zHJK
2mbsxkgy8Y/Su1re5eEZVQcf0sn4k2MOSH4HOSVdhJHHRHaFGDHUdSeeYTq+PKXl
d8+qtjkdXCDe2sW/Igx3ZU5V1Gsc/ZiEMyGxp0n0d1SQpmY2HvWhcoUGioEky7gq
oy9yfXKIKos3hipCbvis5Fqp4Ihn95NjUQhzbIZYTrMefnhImYqDqsKyImCktVMB
hxUepLHfamnq0/AbfDzeYetIdGumIgfrHCAY1BjKX5cYDUXmCqKs9W16xyrrkkQN
bAuNA4CmXREh9j8fBjXMAUBYGLlQa9zY7wXSMTBptYZFWPfsSfNCdv0WCLIm5V5z
1dFI1UUj7jhQSmYAPxEt+K7YtazkU4orwbSjAM6dTQpcF/5eF5INktQj+Q2PhlHQ
HK1qwvGyc2U2ODHSizpdwzsVTAonPcgrDcKMDvNCjE3O6CXYXEAlUrp2DpqGIEtS
jki1jEN8xoypYOdJ1P3rrCSOfs8GzielIGtaNlwEsWLQsOXnbWJCkBqwAckV6cCc
e6MFBfqY7ef2XdigDsbm7yISEIK+sjEEXgrTF0jdUI5SBOir0KYZisAeZGuMAvyF
kVtnI8PBjZiq7tmFcsC+vplAdr2KSuvOGdA/b4EY7G3rculawZUArkaiMPviBtvT
ed8/oYsyyXDdk9z7AnVVROfT4DPRVponaptbZWxSrvm2W2I0a86eSd6W/4RaSA8J
RZVbHGBWrh3/MeJU0xzGFumzaZKz/MhoTG+9DVLzWvR5PEbO5Pu5o3Qcc84co+dj
m2B7y8LuPybqddq9IksKLsRCK1YR4IbASmTiv00grx3K/ruE2YhTcKGHJsWBNoDv
pBcA6TgTbrsBUnLcKlhSfKjzSHvOOktjEtHc8cVJLmDTsIKcGRIDjpdIj168LMwZ
gC31WF+csUg+AfH5L4wmIVnYQNTiAkF35PhrWIpel7qBDXJmhpXd8GgR4SFRI2eZ
oADXfOPEEaGJm0uO/RAkYpxeAD4asO7ZQM5FZ7k1YPiwCDpfUIpc66VVYuXvuOx0
Jw+Su1Dmfp8wnlIgjSMPvxnHdXsRVoSKhuz2/rtutgZu1+zvUh4OPEcOqb+fxCsj
3khPlCgswV4Gz6fsYR1wM5hcHzExLuIE/zf4DX6C5yLpwAsNwi2ic1KR+/tGjEoc
CbOEC2KtfLuAN4owkzXbE16DTywsEcsv/jt5LNBP7DgrWDFvExSavEljrUXvI/J7
dX3ETVgJ+7Fq/9TlePRD9Z+eAtIMdhWGkR1QzRnwecyrg7vgSm9qUDW/KzhdAdMC
eFlSjwOPdGWPci2+0bOV9SC+83tEaLw+G0I6XSuSY3AdPJlUv8/XcPORu6uGSUaG
X3jzW77PTLYhi409QuRsER3yDmPclMCKBHXuqg/ZPFJPpy1AdcGmilME0Fzzi7/D
CHVAshh/l+aaiDKjvczQg4zXr2WBv1/10F3Gxs+jwXkcz6+hH/UD8MXRCloZC19C
9T0bA8xlukDAorNBj8DB/2o+rvUifLbadVW0piL+9m/NZiPe++kKqM7OG2yp/4Vk
86l962nvDM7q3TNrC9n5Jxm1j5b1r4mnXDdw8wBinuuKefCE4fuPEOh36JEkIvYI
p0UjdfmwWR9g1k4wBoJ7VZDBnkbLwrePL0hfySurtc00BwOT1c8y02idgXWymy6V
6VvHmdCP/c9+31ELyAl2DPvfthOWDEIRJeS++WnvvinzPhO3yYRlK8ueF+ehw31+
GO08GKJ+Hsqwzeo5ykTz5x//g4Vr8tzp6P0jhySKr5vYNKPYAY6e5IoNhsD6FRRn
kaRGNQ4H3QxeMwn30JhJDqf+aY7cRp2vSb4kzTuj6nRy+GGXnSi8RwpCSLaB6UYP
XxVg5B8vk3nowfJwLveSYzWEyEn//hqNInJv5ejWe4U4NhNcFIR1bNnmWPfx4HDr
20Ka/YG2g8XNKECL9lLoemhHfGbVduux2+56ZeUkzanOglB8x90ROqVyrCEkvA7y
2UDJJwrTZFepN/TrgObGYNXHD0CTPtx9PC6OR8ZFYY7wUi2y0JUWXBcNnJWpg+By
uiotVdti5H04HAS8jC/UoOBawZ2tpMC1OAJIWWnQXiBMyykq1cIg8mPvUZ4s8bux
+WeQ1Ry7/62CefZvlipoYaFenawTVEjHoyCt6F5DLfdzIRQ2tfCj1aJquri6fn4h
gdMdK+/edwS5q2LVaH3V8+FH2yJv+rCHJOEhDZbfPtFmjp5RIDj7dCpzNUY1Q8zn
+S10XLJgBwOSuMeQ3xauTmgrIH90//GV0vPfKCqqmZqbki6yxb7UkUgNkjnbhhbF
KloHThe0ErzyCezmHDB+it9lspxTImWOYkzfPnbz9CZLj9gG25Jjqt+mfGW24dui
xkj8NcbDFClLDs6dXqDrfUP9kWpdt3Qxn5X4nm/OXS0FMwXEyhBKabpr9vhL3pOJ
0PSXsTfK6WehvPRvYaSD1VMdYBQJe443h7HQHFhF3K1ogbZqa2z5XHlBlIz2d1qW
oNfBj2dqtXSYXokqB7AIaUlkSIHA3P6n8SQF8Yb8bt45p/+nKCIXppL8V9E0XScm
JiU/ybL95pxYpM5T77mK0e1iBTrw67ZqgNktStS+zsU8od0T/x9XbCyAUgdO9bcY
upm8vFbm9AyA7890IB5ijkhK7/a/wOEHFO0fxVfcoFbKTWrEbtE+3o/hkGCSkfCA
m/aRO00LeA5wAH69Oc7eKyWPDooq6eMKBXamhJ3fWHHW0TEi0KqAe2L5AV8WD969
6B0BCfmTLLfsyoxDZePv9NjWLwEEDtGkgHSdfcROKPqmRr2jDels5xH3Q0FZFjJv
pMENjoV/o1In2Hrv4MCuXTCp5dhHjQ9JXMt02ZYzrZorJOxP6G1Z2YmpK9AVLgWX
AA0szygkWQBm2m5boP1gFIpgIyRitaM5mEpu/fUaKfigJShGm65YdTZKa55CfXya
/wLxn8vUTUjiN7Ul8F7WIc0q6N81oaHY/VolxnhKzBrrL21ciuwrKGjeKNyL5Crr
RaR0f2/y51Xr0vW9WfuKoG+hNZu/v/ZIt8lpiDGyLIZutM4wQrT09BXEQGv4zcUK
e9PdKjn1u3F4tHpuERxhqG3+87VZdrur8Qrq7YtyxlIbSnxiUqL26adkub7l0wSh
aEL4DVB3gctx3lZl2L9MmHEC+uCNyFT7GD4tP9UCfxIBmhrMRw5IxtlsIJP+miNX
ogVT02GTxWRqqOAS2SeY5Iksp0ddvzZDuBdEtXm24GX/oreGDMccRqHJHuqxomC6
o30z6iG6LFIQGNqDmYYJaAhX+QEDiT+8hb4ZeuBWCzhFaeIWj6NDqUT33IfaSYDj
MS8373wJ60PFkrRlwyE0euKropAtnxh+AI/JwPdljgg0mtpqF4B/VRHrR9r3U2J4
LzdT5/9R/ArO7EfrADK8pPEGaS+f91Nc5o9wgT1kYxVcSeXk6qKMO+nra/eb6jfS
vGP/o0e/x2RdgCX2RlDqiR0qXKPHCkzmQgTVadUZRCui0HZ6xFl5RpaP5hy1f1Tt
gDiL51VSRVNbB3vf23sWGz7V4hVrleWEnAnx5GdPB8aniP7n2sDhsmTQyB3UTZrW
xklqppj1bFIL/P2BkvjxXXlMC0JmjLlJpuW6fnc62DRepvIp/rvtMqvp2Uu8z3hW
r+9HYafpPV1sHiWXXRQdszLu9iLdtcTd/L3nuwzvCLQt+Insv/kKmPFu1Akntfed
b/tWLobaCDjTXGtTKWM2fBY0VSkbB7sZbs2kgvSF2+1BZ5b91ohXmB3iGQv3C2yv
BSH7JrhGco6mmnTcI7zylrmChUViJQmulHvO1e3vA8jzSrNhIO8uR03n5qWzq+he
E5x7+HiQf9gc+hmcQufE/5xaCOvpKlhoLU+chnnHGB+Gc2CXqrT2tPsmovGzglEx
HsnGp/UZes1OMeKq9k2D16drOsByTagqsazw6mMmHejQLIA24n8UbzJsXRtXNHdQ
id/7KUWc84XYx1m4FlzScglWO6e1S9HtUP0qjKtklyk42d1aEG3uVwfM7dI5V1Vb
S577+u9gxJHdPbOw/RWwGGrTdnJnTruIOwanwiMXEcZwNE4WdhgA+o3twwb5Ze0x
MyiY/ViZy8n2ITF7Jn72Xw24l7APDNQc8ZbfFUv6sbVH0Xya/Y2Lpn4alUlRxTD+
HrnMpIkM8LeVqPBq88wqUtp9AOJ3EYdz4K6oAewmi4H+P3i+9V81snvL36ojZSSc
g6nAe60Xyg2Nj7sns0OozMyjnO5OOV1cp9cgz8FrDSPoK9B9TKTfApLjR7cp16Zo
YdLMdBI+8w0tylNvqjDbLPiwOaSYmEQZ0X9IZyiHwws1/ijDerBdHFu4P1NeEGND
6/ddg69d3R59HvO5EB0msSXgnqnsDypS52xllGAsE1bhML09PinK1kr6EEr+dCQm
DR0sOxJz8NY8MdOvtvga+Nx9E8S62LPCOcnEHpOGozK7wtVizqKUKDShoVMcC5BT
GOlg92ECrUQRcrFuc/xTWRKR6ij19wyRZ3HNIINiMQEdfp24v91o0uZdgmmYmVJ0
c1PeI9xQEXpxP+1ewFiZ76yoqLNxk6ErOWDxHzTrT826puG0q+Eehcn9mYFleKjU
YS6EeIa/z26B3wNHGsQ7WGf9Q3EFqQ2aegY8CIs0E3K9xTTn7qCbzjPTyZ3ql1Ji
NJAqalQzVFLNJBKmB+OGI9wCsVgE0f2r/9FF8wjM7z8du/zBN8eLVfvHGIvpPm2S
rkla6qSVGdsgsW7HDS6XTRlC/SM0PJI8OULTO2vAw2mS8Rlb2yLdgEQq104627tI
elzK8z8kUgB1lyyy9mzcmEFFv9pU/CYeLYea58DwtUxepVi9hCyd+2trQUxJ35HF
MhmnX1QiFbC6MsBbK9sEY6rZ27OZwhLGx5I9Q3uxRrCplVWt55xmCUQzPo+I8/ZA
2dZ77/Er9vKeuoo9WxDQ5buxEEmY6GpTRuSM8euQmlXAqAPYFkLgIjhhmM22Je24
bAsN/COHp48yJz9tZRG9OGAJWFv7X37tM58ejTKqJD9GJRVdO+XURF0qYZI+Sa6C
vc9iAbl5RZDj7/ooQPpRT53GBDEnt2frO0eL397DL/2LsEhqpBma2qQmR7zDYtsY
zOLKjuwqQ/pI6MPY0z69b8Wy6KKlKH+5xHOumKQqV5K9o0yhS7EAumLhqLLYINAo
jCf+CxUtlJ1Ym/3P/kLJpypyb4193iHUrgB3HaMV/wkIz7M3juZExlK1tYpJQnte
QMHeOrRwo/VU4s32T8Og3QYcwtKvhh/n2AK9vdb2JBHJ4S/apAhUxgZPy20pJq+O
5WxD+gOyu2PtxSZJO8kQ+T50pu9RXc1CwbYjhyoSRO1Q+5jerLGUg6/lphY9xZbp
9dDtqKxqDrvPZZbgjI6gXesC4pTG63D/42z1u349DwfAd5etTjaoeEAo4Tip9SrH
BPs9n80XjwDRe1brPbDq7eNDweOdohGHXoyWJBT3D3PANIu/7z9YUyfQcurNMuVw
DiK/d3XVipmELvjdFCm0sWs+qC4Pe1LiHgHO9SCskVfPUvlEvprCijwhDR47BYbt
4pe6nNCl31vu46fCNMos+smqqXhcGOZ4bXDqAj0sgapys0pEuIydKtPrVwuUBlKA
qBs81eUmGG2q0O6AuB3RjBUwXO/XjKxsJ5zp26rXsfp+S3/GVV4RAjLohfCSPX1E
OnIEJ6f/Y+e457Mssz81MrhEKsbPvM8x8lprouOudI45TluvW3rTWbo1wMP+GnN5
6c4Q+NxJtx0KQv6Z/1V0hO4nmmTJuN3ZAHbwPiQr57SyU/1HjG8OPyCtEgqAJMFU
BCRJr/4ixFfMeLXQrttCEmhbgvAGLQYESi3YcbA3AROEIYflQSls3X0oFNAxzaZe
YVBSm6QpagaJ2aIxgJyOd2wvTVnS6tBnq0UeWczs7tA9WwI4i1pbPTaASCL9jlAm
UrBuS5bQ6WegLOGiLyEUy7oejRPmJnAiG7jDlHQx7fmQYdtkzZXXANrHmhJ42GMZ
GdT3iQCefN265OBL0B7RcGdaCeyViewxuKUBaBE8iU51/gx8e1jDMRoMWycazuxg
/yEJ/C+1f9IUu6MhRRBYpQkfZRDxyATRBNRTMuW9WQyE1dfeRWrcqjAGGCON+A1J
oU/G5SM78Iw9bo8s+3FllJTKSnZ7fy/tG5QKzYkUn178Ke2S4EOyCGEcYH9PsIJY
K42hulRhRJ807KI9nbsDFR8ZeNUef1MBKg7iNb/Co2upAqsGoe7Q39D6fMfTUbF0
mm+QWvNNgMt94DPhi7zkLBqzCSA9sO3hBJBGkqEI7rOsMi70IOGVjDe+AMCyRCAN
KKrN4v5byun5IcHHQleKVY/xZpOkt5Q4iU7eiLsv3wqA+H4ZiZk0HHRg3Whaqxtd
2jz2X1o5AY2UmUVVmPpMGd7EzXsvuSt3cf8GI1pGT9qrRYsUYHYIU8t3Ua7F2+C2
sXpUHC57FhOdV0oqTNulD7Q1bZc+usDfoaDrQayL8eExKdT2cWT+0EhOw19t1opM
l7fIUxXmYgQUi3XRSwhupthJp/nBkjyT/KFSPKN1+vRmPGD4BhtNnV9+zkj/ZJ45
LUKN7boxd0YbDJiRwyqXN0I19p1yO0sHxE4Ucd1VJKEVJJUJwypFb2Y6Gz68nteg
QFXUwkfH+zf59GEFzpAku2Vbrfxf/vx7pOYn8NbkBZ56u/3ruWSf6umtGEJ3uPI8
YbLlBMPAJ8c6jedqIGj5n5BIvTx6097OphOIJNFfUoG0cRePn3HlToRQmNonCt6o
DAO7JLXo2IvHe3paMaBS//Gfv83VzbsCl08i7a49DgKi+053SjOdHW+OHsBZ0jvZ
blNEWpSzlV36Ae2zjG78FZ0cOAXLR5n3C/63HsE6cyIfPjMyjzTmwztlBdcBy2/G
HJSgfnHwkXTEHzcfcqFJAz1ED8jiiPdeUwBaM9fINezodXLFfeknHC3mqYKsAOH4
6/fIzoWlYNL2xtwzipMp3dWpdCS5A8lxzFGp9rfKckYKtg8vAzCNOS2PU0SOZi8C
k5mU/39xa9mjF5ON5ufa7oJ3yYZsb4Uh7sPpY6eiCLnsvhyDVQwpKyxMagcq4qjU
voK8GuopMcVP+rg3epobH31WQ1HS5BpWL7tJk0jMa7KDcv4JkW0EXVsQaw6zvCIh
1+vQHOahFZYXYNbUccGPuQMx9mTObK7kCgflrKMOih9yg6p5SFZWx8W781h2TCqQ
SORJm+/A9YerIMVZdFam7tiJl3XW2nCOIptLChC1pVb1mFgF18OZZZ6NkWOBIiio
7E2OEyJoMMQf2RCRvOAycZk8ocR3AgkZRmnRWQ1FMCd+NYpeknrOebRX4Kik9HhK
RwMrUgNG7++V8hF1EUaJnrVe0lnw/5XXn0nv5Slqf3SLuegSk2ss1jX2cdm1BegL
kyz/SY++Yi/poyWKIDHE3a4WzI3YCUdAxpcHRqCg+q+MBqyCUbCJKm0Gky9vpklk
9VQ+kTmY4v3XdSYzb+jdIFUPn+gf54jY/K4NiP9THHtTEfE3ES/X7QuoJtCN7B+6
kNxet5VygEeSbWdnTjiSz3sEL8xoRbVGAgRSz1C6qRw9rrkFAPGCGlTlm7IF0gSC
sJ0iA2mQAv6zoz1EpH3AsipBeH16KpmrvvmhEd5qY4MoD/FRdWUlmd3vFvN3x2ul
3PYTDZJIHhXvE2zivjD14ghCN+mcrWw92IV9LPXNJwVrRrgiURxiOYBAdJuY628h
LHYXpZGD4iL5CGnG8KEigX7WLLAgs/Jf7NjP6el/lqmmCrcqYDDsqVWVHSRcXq+4
eaTDjov7GneC4gYnRtKDs4/voEYiaJim3gfNcNHHSxa1t8cbq2p43qB5d+7UpHTp
cCcf7S2/n0uxqL71msb4IycCRbnroG5F+iU0EOwrVCI4pP3EGy4M5VwvqoTfsFwD
ktWyAKnAcKOOGjRUBjGxR8YuQYg/7poOLCWCGqu+i3NDZFgz7hy1DoKm/DF8Buuo
QQAuNmVkLx+v5Irr5WCy/zXslMfvy0wCDarzXh75VVPjzACfK7Sdrkd+mdGVI9f8
IsoBlSXGa3xK46K9mA9QNI43tTxsalq4mZkAtiJqrUkw72NSggE1SA3Dt6wW9myx
pPa98VdqB6l6R8CCs5JjkRHtDHk5rUUEXG6m7FU4CSyGEnkOp/krmQlgwzddtmiR
gA7yc1g+d1MtRSSpufAFXDY/+xNCr8ZZLgLX7Q5+LSwndT7a/BdNBGP0VZHP32OM
vBeYbBMbt9WKFuxyB+1s4yY/Q99J2d0txMINsvUV02g3FSojpnRByxtu2vmXmhC6
M93LXPW8WPLmnsPNjYEKnrFrVXcJy9BTqmpaId65dMoppdK8yR9ccDhJsVd5yGm9
U6PgQP8ftEypa1JpGj+tNaO/d98dT5SrYX4EqLa1XSUG7SuXQqR/L0kDTj6Gl9ao
ofTfFc44YPOInS9bydPUggqnSew0jElZ1o6THUS8+mOdR/9O7W6rd+9vsYbYgRFi
s7y+UuTxpBTqUkNOkiProgQFOnjTmy0BweWJMl41qCIPedmhM+dwhz1vRL+E0inL
XQyPIa1Zp56wKH9OenLIDqbjXzqOK5RQ6+Dmvj0stXqIEL4TxvFnHdnTSIHNy5JH
yGZvATw6L+WmwKbalBx9SiM9dllG4+uCFYFTaTFp8de4C+tIi5e6U1YZwuLjmXXZ
3AVan3dhjhRoh0zwrwOr3vY0PpsQ1KZzmRcBSgAZfjmCTjDlsnJuhjA2pIuXZxI9
EvvWo9FvpnXgEHRJmA12vPu4pxpdxgXsZ+Sn1AV9ioCct+/E8NFo01HLpwNyky1n
DQEOhYUXJ+JvdKGKLhdJsRWfkVb2QDB64WRGl08R/2sZq1yXckNTkqS2s/ILARnw
o4VOTlkNgodpw5VcfKhTi23aZnLIajwKv22olwW4Gm1alvtnrLF2O7PeyFosqxw1
97CJUomDpRrQVfNJK3b49QCaUK/pbZhGeXN6bCajOlNwoKdfMFj8Oed24DtXNfAJ
BL91X3mnjCFgBkVYNi0OwOx/d6Im+GauYVZ1FS7ovX/bVPvU19xeNqxPSiuPX51X
vwUIfxU88GSIAp72iR9uV5iCQdmd3/S8gYkTKOEBUwNzZdosXlVfuuxmZpoLp5Ny
D7FzMbbUO+6lS06QB6MV/isx6CZpLymupg9gTYwx8Ml4SUXzIw97hLh3X4QnumUF
UQaOr8/iHsAmemeOduD5lryDQP3eit1JtmwQUQhDfkrfj/9x1H5QPirVgLvJPQO7
3eVOgHJsdI6DoFbbLfo1pQqvlHpfyxG3EEbimmpmYlzX0adW1URzee59EkNYADsN
rpj95efkQwJ/P5KDXtQkwGKxG01tywS2UdlxvqxeZgt8HE08pkdmKYCBtyID/fry
7G2LFOxAsxkJc9JPdUjEbUNAi72eFzWnGFdCGIKzZsDciF/U8AvCIytR745RrJqW
RdMC/4j/MewMkaF63pAj+cA3U8OJxSgiTI5z6HjOLPHoaeWwb/tf3+2CTG6tIGvm
MlMfhEn3qsgwmJ65N1D6lyw0D4uve/8ifNrhpEpG7PRW7TC7Tr9x6bSs7y6SV/ou
Z7S54Q/vZRgiRLnDzrMfcbEE6jtbU6D56tQ7EqIFhyskYADl3Y4beX/RwmWxls2m
2g1aLoFeTHvjbmZsly50fbl5aFnmot5wRu273oMSuhqTIugfWaHnaEM5epK/EDgp
OzxKCYP7Ch4+Q7ipdvp5N36ypGbkeGzPlbOzJOO06I4gizFxvRwu0aPR8cYXetcN
tiL6vvbF6G6Vro8HYKMkCR6cGSRsA5MOf1uhyQYkSzYDLdwyfvD3DwbX7MRBhpwW
QQsNXfylHMMtYjdEyJG6QPKo/4MaJdgXckTvArNNN+0sfR9s+wATWwuT/PLk4m62
FkqRXkTKDWOrupj9hY0dgYAfBHmBL1hDXJUzGtEohEJOaIRKxrOY5ltQTwhQ9eug
SfCZLU8p3ZGUDt0Muzu5cqSS4o+u96pF1yRMCVrsLzLLqhLlh85vW+AbR6SO/099
AFLWa0TIUXI2gff55eG0TQV1g3NsI2UIk8izl86BJIcLlMwO90YJUkSzr0NQGmhq
FIBinHSu54yn5LusSiMrhM9rMsgGOpPRXW1VjsW3zuD4RqTzb9vvS1/gjhZT7mYH
4WduGjVB3Z763t6OEQXqKZrKJz1pYSm36/8yStD/eKSlVxLFXwcooMcOJXX9nP7G
DQKDh7AFkcBKwF8MkvcKVHbSnxcP3I4Mp9HuqB00BUfrvXFPoaJXVaMfTUKwiWd7
JCFvo/cbQQJ+IXXRIrkKJuoQ6T34hndlgnEHoMUnYfQiUbpE/NuwRTNfd2YLuWf9
Ur5X5scK9jVl2GZ9ncQoyDIb4+FFIvKFa9zVIghCHVJ+xgWZdR55ebwWcGJdGtso
Z2Mzxwc3BDVAErkXhW8bWk7hZVuoeKH+czRuhRTkmy3xFzwZiZh5Z1HkT6JVklZZ
zSCHj8mRWdR+XRT6yk6Qjpmv2OsSRJbbLR+bgPXZY4hQM8z46ETfFzCY9JV6rYDm
fWoiqSafbJEg1flRVz32GGA3gSPMFstKhLzb0xjXz1Od7QX2y6T4eK1s3llFj6Fv
WWmsH1OnfIJ7UVI6MTdCBnc67X6lKLDa9Yh873WD3vqV5CQtIozsrnexz534rf5A
h7kflnkiOqaouZMZoVvn/EiIUmRGrP9lzE8Y70OLQ1bWJHcoJAuABhVUtqw2dLOY
chJ3GtsvYl6jytia9CEVsZ8ngh98phDy0n9MXP18rZmKQWjpr4ric6+j9pplrUxq
TC9/CG4OSkm1rpRlG9xwMNayR7Mepfk60De0Dir3I92///3wIXP4EGyT6TTHSaKA
RGJSDaM3rzdyGyXYh6oWJReu6k803zxaWFgMyjRVDF+JvSXHdFK1gl5nQSN3Khrv
oCrmxyiAO8LCFVrYepInjWIKiu/Lp7grRceXoz94SCX2wDet9h845TO+1Ds7UFZr
h9H2PsazmscsvsvWbOToESXS8YbH9b4ArJZqY8mQilComckMslytBAy4cJM+hURT
DoE/6cWtOLtI41HMoUQiYeyNw9+ROnFSS+21K02jJ3unm+na5Eldu/ykq/anYrqZ
wSTG9A7gUD+iAAcbXh6xXbTHJXlI6+XdqnBYMmpVQYJkA3xIVilmOK63wjy9KonF
yphBpoV77G52V76KDImY6ovINQ7RLIHUrkCHZdGvad/obnA/vxlv+l7PAzY3D6Lr
QG3OQ8XAJYtX915B5eiyIIpDKk0k3sfCavrKnONa8Z9UrMhfuCDazU4cYdD/JIUt
QqifU/dO70iwtqITWM3828lUmKTj/b+tqVh0Y3vp4Hd3jYFyL76Q7BRaVceW35yd
TzvtH9++fU+wd1kHVKRmjzZHSnBCP9R78LPirnTXpXIELMAwiGHbOXCZPOQNy2a9
CVDI52aXyvgZBEusrA87jy0P8MNv1snGBMX0pFyaBsSQFiGur7ssPR0p4PymNBOX
sdEBmRyRMz6Zm+fe236JvtNqKFH/xOjm4U+QWwt12nLmc45FqQ7rQEalIi32IAsq
IdsacERrPttcFm/yO/NYuAVcdkxLvg2tgvoxLl/8IXKFGkIo45Q4U5BWbHVUXiWZ
2VwdxNIStWV2qUzLk8giODCuJkVEk16Uotav1sRk8XLzDJtosqHLaKyencbFhVOf
/ZDnKxJZ/Ss/cmTc4oIBiwxMM0clLf+V6K9DW5kgw1NbjGkaG7b1PXAUcgjcOgp5
cNli8MgA7HpiX0V/kmDhuJtPI5Shy9n6A63UadpNyIO1iP8Bx82NyKJJAtcW0fCj
x0Hw+K+IMLCjDb2RazrxEhrbkpGWBGATt2H72lV+GJm3PctYDpjKhJWd6s0GhZ/R
frAFUxqnuZznsE92Qahfe81dD6Ad3W/KobVw342k2TT31HjAiTBCsMK4mw+0CtYZ
ohA5tdEz5L7QYAvDa9awNJ/PDQjTd+Z9jyxg+Z7SchuW9w5z38vgmotGF48DPLZD
btM/796w6mXGlSUm2Ycl+6S1U2jHgPMRFVVq89lLI2gl/CeprF2JD3Wy/rTAkw4u
+Ch2Bw8/ncKO+oWaSgiClTq+aQyBSOMW0rkXjAwiOGga4wTda5ls1qtUrITQsbXF
AJH2hbVPHSq4bvHBNg1wM2zA2rLrMQ3engsF+02cl0tx9QsWWUXR47F9hez49yNv
vISSsqOYQnFpCxTon1n+byuKMEEdA+4LQzRnkNgMz5UbthnJSyM0Ju4wGQw1BMws
nP0Rmfsox+ZEYugtujLDBelhwB0KtuXVWT9SR2Tc2nzbxGeqJK0cQ+vTaVtNgjBg
6DHqqoDLeYIzWeG2Za93qccTtZqWLIyOuPQp05cUwNccT8UAyMcNLdpC5u28AMrR
fkmb6bA8gSimrKHrkdWqc1cau5IVKtydBVBy/KFQVxKirZ0B7X3IadERBvrmzSuk
1acoqilKAGfWWg2Uf7Pfy6IuUsV3yYa9Jj42VlxIlmFwVJ0PPOYH1MND4dLF1J61
EDcd52f4ZCFT2/0p2lk5lWfoCMM5c4W2Nmg6Um4Uw+htAJjgUenApiE+s5ow4Nvb
yxHN1BkZKr6Pjoh5YHB9DFK7OBQmm191KK+li5b1pGluLL7NbEf4yQ7JnBgW00Jd
nLJjiAkGpXXWxL1azJvePbyzg8W/AJ6zvKNzW8C8aAd3JcxeL565ucIqgA0fFXDW
22i5Shx/ZmZAPB2k16CLLfHHAKgYA/9vLj4855A3rox23/AsBRpFq6w/alJOw5uf
bssgw1lqBQtHXRsK7NPPAHU7BRXgRqW585Zd8E//fdmttczWRRDZ6jYBvZgzdIqJ
SzDOexvPiWxC852MzJQThjPM2zIcyexSAHzFtXL+/ZoVWBfZhn2pIk5lgsC0B6Tb
M0j5ISIo4c3R+NIWTJDXSpa/lz+WaqiIqH9Fbkr18R0tkm7aytOHh1ZTlvh/gwSz
qzBzvzNPA6B0a1V8EuqG3NKMiNjbKHZp63pNYUMlLOYzRmYLMDPOdcI89p2+xFUM
fX7d6iuQin2IzCEjiTbXzZ+XHEvWi36/VpwUhydYatBrAnI2N057igeQjXPtvEJf
y3Dh/RdQ7zmJfdcEroX16ozyQHazl7KFjoOkc4Go4g+jQVCXsD5A1lYGhxakoEuj
0jPdpYnrz53XOwG6wVGirigjvAimzzy+TgjptGemAGprTWB9RZEozHP5mSlu1gpn
6zxhaKWeoK7LMemQd10TUUZxO4pzJxeaQ44mjH/eh1pNNZdjbhp+ok6ng4x4427F
a4NGLfpwtvw4C0RA6UAJan1ffIz0jGOWg9pAOw0Z+BmqxU4+5QMCpxNeeJk1xY5N
2FdxW/PzpobBkOs8a7M6XE3V1Gmcma1GU+6ZXCrrVwDfv8IA4J2dV7flZnO56peu
9kk/VcQhSGsjNZZqtXKakR+YS9C59vraJuDRUJqwIMIOFPEfBmCgmv4jc9BsVc8W
77X3Z4zRpm2BmQbCFDGcX9RVARt43536KVUoovP2sI0v2sxUbL6xldEP7yvyBQZL
Njf0I7Fqlz68NVtT5Kd7s04TLyLRlmOKvoEvAo5uu8jtI02EAM3FMmD8vi1jhRso
8lHV84Lcy80gqh3JnXXVZI5Hns6e44KXhlea4nngzQbTLtvMHLwD/aj56Q6vfJ9S
ZoDgiQSbyWkTw/XDa3xE9YlCDyStLZL0CKmOlTgBCxAE8FG0Gj9zvhFONg8tNwVi
cs/gF0GMGW0gMPiyV5ozA56Bx+4aNL59C+8V6JcSKXJyeCiihQXl9kmOAMRLE1Os
ycERUUd3hq4MVQT4sSJ5BTRCGCSxVdx7zte/dtNlYO43jRy3KHOSb/5QwDtWqXng
7nctshdXnMD41pWxB+7CQTPajx484I3691jBnHy7mXHq/KtU3CN5MnUE/1uIxM+R
7gb9rPfC7hL8dyI7luxY6XYQbuahjbd5F9NY4sR78wG0XvwnOtUVXYzX13UaCDMX
gd6ee34SIPw8o89b95YZ8W/YadLLyZuOqdSoEl7NN9ue37s7y5bAzmCzmabq7VZw
BPDK8L7dkVh8h3/73gvKiWn/OsoTuumgy4xUw7qhxiTf+vhk5ybARbNSenJwRkNn
Y27YThki6iD2jQhh3KYsoIoDaVDNdsU4BoHZoIJFCzx3DOu2Ih8XmMlqD+TtwSoV
R/WCzAsSqsOnavVIV3UmRBEcZhT8Rg6hE1yRAFzwNZCN046hkb2ULk/7KTsGfOQi
IZmJ4goyUyBi/sczIYclb0ZYYpQRAGsUqelW5aUBYUqLf6yOqLgs+0yVZmWiDVOm
bkkoo7oQd2DTQRxjs2kd9uGu6FtTb7jL1KXOZUYEmiPb8z6Dyb4vpYIBV4xNnOPF
SS/FHQhv59sQGgrYV6Tvo6e6K1vE83hlHcv6K5wrF5ejLVD9B/5vDCPOBGl33EH2
aCUt3tH3OF0Kyiq6A3rHpbBWG4p6eV82J6WMrr9dDsrb5sU+3BfIrwKegb9DIkhQ
zzVherLUdMbmMYgpHdg4dWsFhJ9p9e5tfpOFmQtvLxjKepVrK0dSoBvu1FeGNbRO
kM7zUK959ojw3CUT7EsRZ27j44TdyjPihUlqokparWuEI5HWyzHkqt2THPaHsOD5
VVxImjxG0zSJpFpSen8qI6I8JWLyuyrpl9ZsI8sTsFCMIlc7Z7EsAMsrgrbHAmPH
B5948VevoVXfKqqPkF3ehnEOlPS8QRRgJzHFy1QO0F+vh6czcdSI2pRcp0km7u76
kOMpzlcuAGozo8VdNN+GvMHpjxg3Bgs9jtXe24QC2P3goMspzkcjniknm9mIrmVP
VEymzcvmGljh09LdNCINiNkUGQ/w3LofFpcm8N+6e1DFmxRvl58q2D3fPWW9gbCe
Bd+5YjaxO1w6GUGZpzRnAy1uVrRKMv5X89oyztYeDqJLhlvo/A76NHiOU9ClBVVd
e4cgrUVbK7N8ygBP1EbqTtstEGdkAcozL3560tIRe/JWIiCeqYb0via5Q4GA8cHZ
SUCOXaNU3/kjjEMqQ/cs6cAVmPhFNczUm08yqNUOYKSs3aardBXiQ+sv6qF6sB0h
xhrFOsJytg3a/sl2k8Wfd0zujxp+QSHXZbtbsdTXJ2Od5LAtFR6KnHHwxiIJ7SVo
fe08YHTXIY9nzr5YMjDG2+8oohLM+sDHREFg+t7brwWY3SMZOKUAO6wQ3Z58yGkW
JO5admHgTxfXJVEdvrPemYO9hCvoqO2Aia3K7kAN18WTyd4168KcvslJHGR0epyD
yEl0BfD7EHOcwJnKF0r6x8+mDp9yK66AHNEosWjwuT5zwmtbuscaD0hwR3D8RvqW
hca9CAr+klZ7D6vulkNJrrYeyWUVkwh4JuDKZzLRFZgV3riK+1LFWrUYkvscT3zH
k0cDGhbdmMZWRNCCXo+dkezbA5csjMvtfHDS9mdFaT6T+KFnJJ2AF9jbygiVrEVs
vvnRHf6r1Uzt7OPYo6ByOz0I3H6sDDGRwSBEIwMKkCjnz0rPOEzn71bQLjvdqAN5
qodXKR53IovQyl4EZJBm+zG7lKGuqRK1rshdIMLbsHxQMFhT8ooHatIzpUz77g0X
CShBok8THfx0KPGldvtHVEq7oRgjeKErZL5R6Op44yZ0MRIZ9arC35ZPxZndK0b+
3WEHg07vdb9ncc8xkhOAN1Mt/QO361tJZMcxmBmE48Eym9xJEnN7pfHWFms0lNhy
njv8Mjc8WV2RzCDc/dS5vuBTNs3ZbStaUq7zvDFxaS08vRKoaCE+Qy6EuhwVy7QG
U6ClPJdr3dSHcjDctIG3Ztan2IbLIEdi6YbXo4/amOq9/GPgk/wR905p+zMqlZZj
NPFGPKylggm3ojKHfEE5sLEMb3dL9tn67KhuVi5W2sxETVpRj/JkgLuj2ZJg9/2i
H+VTF7R2AuWbc4M/DwPZw+8yWYrSsXvwKbBN4za3Mo58pOzPUjVGSN/Y09SsWZPQ
sou6s0N6Y+4yFmBYXlpYz5sxSsyN7ubsOL0ediNbm5ijbTNYQHwHjhjIdx/aXSz4
w0Qn9ACJ8gcKMtNXFCpuDjaiKJkK0FhfXcFeA2r/pgE5cDa2b4mTkjnHOkUe4lXa
+NXk/0cS/8UsnK9hrsUpDsymI0BhCMQVCwx5xLy0U9pZevSQSJAbHzPeg2xz0pgG
Uz+jIj3bxzodHm1zRVPyn0oBf+SImftUUPZMjvyvwirY7l2aZmASLKNo0NQkGj9h
t2fiizokbOim/0twD5gtQk+F9bW9q+tUFUE2VYwc8zuPDhCQ4mHqf7IkKgqpi2O7
PUW9FaUiAQvQpldBLou4bsi9clodAMOuB0dKOP+jSqCZmBrXVcLMpo5YlJ/fEQe3
0wySnVjkvNEDqQEOfsuiweai1kK8HIK+KdVeWOfs2qkka+W4rNnE0xa/UTZHO8UF
YgXpXeamGhVLdnwqf6Zi87AuWlxFyQeyNrg2yXQyFkiTa6bU3m9h9XDdyJeCsN4T
cq2p5ik0zyZ4VfIeA/0LHlma34U7hZB7adgxVh09XAQUl40fkkDPpvwvXK+blm78
6Uckfneh4wEZjQ2FesAdICL6ceW8d0GdSI8mpr9ZpshNs8zgO6VH2VFGYuEXZo2T
Zo+S44L1Oag/6yM6qcpZCU/qQVlMTubIkxXCKTKMcIiMwVH564gAjut/d/N0Z0fE
toc3e73Lw702UebR8e+wQke4timWavlzf9zhPqP3zODQLusVz8O+sx948S4zhPWm
kU/VZV5dgQZ59LVzV/a8VJHkOlTouA8ZSXlk8PGw8N6mU9uFjQbkVUP4VTqJbZxH
2ROCZ9r/5cGs6u3do27vHinE6ABULox0h4Iw9+U3EZkHSRnDhycKq0daUoOMLnLF
DF22s5PAA04ync7tVPO/Gfs3qWAxBG7kQKgyykvNGZq/xTcySOrglFuBQmF3Cj6q
wH0mdCkyIL4/XOHxmCARfy4+6TgBAlv59sFXX2jLaLEI32/Vzg1lRllJr9KoWvNl
WVkJ202dyc14Q/E5anNmsvY3hLQlin9Z6Y+J2jnrqPuwEVEAmNl7PQmtIBoNdD1p
tf/diI5/YHLV6FBCRSS92AJOIQqHth4nFkbdD0h8VPIcWVIKTJFEaPH0STK4SzL1
IyNxlKIqzTJrFc4WiJslAR98x7ELx9kGGssEG7SCIUUgOCnhzCKpClDsXATx0O9s
LvyIbJuo04znRnnC61uar+GEusYAByF3JzaSTeSoU8hM6aB3zXqU9fAvUt6d4NH2
eCn33Zf1hV6DIa6zeNKre+fJyxjbjR5O51fzWW3700wvYZ+z8QJ13kVhwp0EfnTU
KAEdjZdqw1vfXLBa4cmcnqZoMYrcXCVokBPA7nY87QA42YHSwc9/yRnYwbUXFh0b
Ts1Zg3NrZC1v3/3LIpOm3rvKPbHC3Xtp3lpcYW2RjH9KtdXjaU1V62/G2TRvUK1E
7mfYj4UHVnywokQAKWRlnDZAqeD9vT9G8l/smO7CZ0RMuhRJHrKHGP/Dn1vaCx2h
Mb3OBMyzHOjqCaDcOgL88Kg9bX6py7buLt85hLquyf0NSv3vKVJOkEqQQeyHcLn0
N35YlJpCE/wKl8CYLgppN89kltA3r85d+356vZ14DxWPCCDjB/wFbltXmq13rpHW
twyuC9bqNmACUhbLCYYCb8h9HwbvdnsmmK6E+5SnzqnhIVaRIornhtW3N9FNtz3r
WbbSbfU7HXv01LJRdm1bkQcaiHpzTubHdMYSWKo5aa3vHoc/ReUlYJg3DVpikXnP
HHSQk4oCo1UtIXlP9tdTu0BJpdGn28D15ngX4HMuRNUwoo2mqsmG3lVJRdzfRwju
/UHE2SOALKupQpbBEQNLHyJnZ6ZIdRoMdk4rfqvQZTcSXkvNrE2XnD3UxFuXUUmL
vLSLAB3881TIaVhcVPMVonAC4n4ZM3wGogxVRFb4iu0qTcjURVrDEh68G9S/3woG
PljmV2Y15uWi5byUGGmGRa4TbY/mk3hlH3uWXxT/vktdOBYUHKDKazF8gQd6qjF9
qvzPbG7jS/rKt8WDU+QMuti0/jUY08sBMzYaG1KxVAFpgG0ec++4XZRCJ5WpoLXz
0qe1wlbSY0pQTh9QLFBdEWsUinpMzKiK57Xz8NIlte9JLILFvqPzKq8YxTpvrTJC
KBmHh9AJSY+R5JytplU9oKQDl2k7yhP/ofjwNLBusEb4R0NbGVi8w6cDLu6Famph
GZckeGsLMLvgmB9hEPbTVlniegAQerdVFjFl1+aFsb0D8PNmJwTItPdCn5fvfGUZ
nm1dK0i4HJIMwSSt+LbiTFdvqkqF2wMh+2vRXoyjrwX3blnpAGMYYSrlm5rFfJ8b
61rEd5m5u+orHBttUIajRjPyCE4AY69JxNGwh+T3X4e4ARu8A7TqhZgcxr8yI1+t
NIcHiXVsHx9aP+1EadlTF/aHYiwYxV4eJoyBv+DaSSrrImDqN4y2BHu0yfuzDTPv
lW/M9Md/TDo6rytvGxsPUbUfMUPQQNd8zGg7NlzTY3YU2mE45Mfv9z9eAgxMAWBD
kg52r1L2BqaBkDlUtrAadt2duJHY+WZPOiof9WE2uv0f0GWbkTAyT+Dx0g0MhSvD
GZ7brhaZsIZIjBDcbuGhaVrZhD1gkIMmsYiiOS51ojtmCZdbImk741J2ZiH+FUFZ
QPAFm+6gyLKeq/nupbyUWh4wx5RxBcMvqMw31RD2MiPnNH7sMdg5s6j6l8gS8moP
lO7kggafeMBsfRAF+R9e7NU1IQ2wcPbzZiwxYitrmxLim3J0P8Ixf2S61vMwMrjg
WvlumPC2DzrB+2D4hgiyj+OYofuZeRdHWwZxmkFZkKyWevhuQTB8qD6dFYu4U4lu
JFP9m5GPWtp19WkN6pbOR7zcOumdo654JvkXvsURNbbvQuvM6gCb6COMrWVeHssl
brk0CYeM2fU9DcjqllO2p8DyzCAViRVG+BkKtPD97ePZPzwybxPdxoTv4DX2UEss
xhclRXSJ8ljlq9zO2l0n2SYnBqjsSPN7VWbVok08rfcSycZHGTyQFj7756IKrn5o
qIrdAPwoQezeS6JTG9KGh0fRFguL8+ymLUvqT6LXG29vYilofEhrF+PskX43vBIV
tsjkKrvQycBHcH4B9/Gx03/a70JCDECmtD1ZmO/+TTs19JlV2vkC2FH/TKvNTfWj
1nEDh3n+yNzqDn229D0+nfyDz5p3Zw++3feBFYVUta1axHvAXyrhXOhrHqNfLm2t
zdGGiL2AYjdhVtcS7CALoRh+p0r0sNMZxvfd+eyBuFmSBYBd/Z//joLQicv2oN+T
4C15dzthY2cfN0SSVRqcmGOWzLgxGh3KxtOWIISSasIiJ6w8GFlQnPZ0CTbjl6JX
eNBKT07rPaFKkz9I4x5iCggNPr0aEehzSq3wpMvWqFtBkEXO2QpUusninDg49di0
0Etzznb1DKNYAzQH9PygB5933+MhjGI5Tcge2Irdb4hJd6OwHjzpWxGLANGrDbjF
NV/7BRZFHZjYuGxScq/MBADqEdUXvJpgKT3qjbfX89Y2QoBO/jtcyqdpfI+QCD3E
IqBHNl+5j7Gw7RMDNFdrP+ILjSvfU00poIDHbfO/Nd38z7MVKYrBVyG+8ffeGyfj
4CGLXRCBuRqbn1YtmwfQASdzvr0gn07Q2kpm1aWSItmRClU4HUf/Zbc6D+W5vBlx
BUeH3+06Y95CttO22wqGzmNq1jV9w2gpU6ob3o95/R6xPBHcxL1UOqxd93ycqyWu
M86nPI00hL3A6e+vm9nEbMiA+pSDCxWKpoxgltTvFQ6QqZIHN41JskxGh/9WNVRN
kMVnr6kI9BJHmCeIFJmSBKIENALgybl0FN2Hbal3P8MPUFtQ4kQwRs9/aHPVhzLS
3J3z3QvILrmMZVwqIIU9sBCB7HD/8gIt//enmkSnR1SW9oKjegMIXntPD6XkMLkW
FIfh9dNBMB54gY4I+n8V+VYBWGDBBzEhcJkR7NrtpVLzlur7UJa2Z8CEGIE4pJO3
z115ICz1JXOoMqLZZXhWYDX3Q1CzC6mtcbIXkblPmvqrK8U5ShvhFmXzyBXLx9zn
kZbC1PDefpBAxm9Pv943KaNL6xxlz5y3JPBSjnlp35aTunutcSnQyaWxOxwff6Yf
kwLOK+/64v6ZRbuiNMR4ZJ0zyfoZg8rJ8/96LNxoWG4grvWyLwxwZ8ngHhNOgzhV
CYEAtUVDsNVZ2GXi1NRkOqIP/Jc9LVKc4ow+u3PgJnomRFRAgOFh6EDhQKRY7Y5z
g3SFLplPTGgxwm+JavdI61ekXag9OQ4i/ed+MQL8i7ME0mc4WOZcpQXYIdqips7k
41ZqJmrN04gat91WkuJCsaZTAvKw03+fLmv4z59eNvDiaKf5dDbE/i2s6bfsbLTa
312r+pmrzFZw7T7MzzXyV6G3f0FD/udncGS2zNYpYFngi7HugTBUhdOmwpKKBqLC
T2PnR3SrFbpvWb86JL+mhCX1ciWf+zvrnopbzMsjnkJS/7HEpwFc8nVhVyCDiqJb
nxxX2maqzubUJjGXQFhoefLAblsAqzgjkI0uRTAX8DUG/OEr5GQMAGgdG+hshcUE
yjhI/3VAPvxkI8CqSJJh6APhn4nCeT8+GAvrQmiS2ZnlUmQsuFd+Oogb7aRLtLVm
vTM6h0YDxS9fUitY84bPabNKbDQ+pTdWf4aVhI1Vh2hIFi66D+Pn6cv0SOytWeUD
kfw/5iGGFo4/EIwjulfQyB+/x4T695N5XwNNBN4ptATrR5nARJsWt6BweRuNi9N/
47H3zezGYMYn4y5XAFXL3G+sEqhHEkBAu9va+JCr6luow0K060P+kmdLCox4PHwj
NbVCr53Q0JP/JHcF3A+3IfNdxYoH7bUL8UOh1o63M2dRG91CZQsZ8elAeOj3Lgym
Desh1H0ju9mRNpfTfClS5Bq8kD+zzDa0tHqwsl5z+mSsQ1DkylOnVowafbLEg7v7
qpZCWAS+p/wm7hPZErbWQb6+Eu2iUUK19IIz5ZlZ9Rfu1o26PO2dZnZFLHxPT6Nt
QuiRDQSgRaWX9tjGE+tJQcrxVGsUnSYO3SnF4HKMrOPVzk+Fzp8QkxGSNW2kdd+I
YVj4jmJ8ocFYtSsqw7eBFpL5//KIXRvkun64/eM+H/JeIGirU5mZX1w5D6FsV63j
sx/pMPF/Nv0RHITTOBaAtmyAimhUfcI3AaPpHi5Nl/7Z1W9Nyc4qXHLbw+ei3elf
RF8Rq1UVcL/7plDveKjnGwmz0RvZzFmVBbFYd3oYlmD24a0iM8vD2XnoSwoHpnPY
go3XGpdCr4Qdv0XRCNJcdGCrjkBWhGYO+kwF/SodNi9c3WhdaZJaxCdj/HRQvv7L
7Mr7KQzOtl/jR2b1IZBOE2J1wV2A3MlBuFPxpVcQNo3+fs5ZZRW0p2nC4m2F9ffs
u8F0rQA5VDeXsgwO9c6atrjU0gesR9qnbtNmDfrlWVPS46DRyN0r7ioi0/9TH3DJ
ZmPktDEYmNVaX4FOIWfbjxEVaFf3gZrvLW64xFQjqho1DW7ODIvR1LesYhNu0IOs
inYeMoxsiD6WXmsdJ+88Tz/Nav7OgL9jA1QQp+5bJTVFNBsQ2XVXpfc890ODfV9K
SeQnZWEnY3Q9roq4+AobwRXMO0fjOjNyN9bh+teobg6qZ1obvNNrymmBHXZ7g59h
AD2IU2R3v5FnfarTuCzHZgrwWksU54w1Fj8/X4T3YrbJM/zj2G9pgGeuRUkbgqw9
d6C6+k05+rlVn4AHmXfJuqNRMb1HY/UE8TjsEud5w+VHb+mev/YsX+9+ueby5o4t
Gx7FdVdnf1XMW6l5EweVUg70gKQkHQolxEwrm7S+tXLrIGoNKv0FB7UsmImKXzHz
cx76lQvoo0XgAEqvNzu+vYvk1bxz1InmGU7guLR6GsOw7gEhKhzfiKF2hKe7hhsQ
RJwlEhrs8OJDIqGh3q78QgmdyFcfNIa3R3o2sqDka+JCpdXcdvQlexJlusAZBwu+
is9NWcDT4IcGqDrSdEisLSEAbsoCJThbtsbkmBqzA1HrOHZODK37ing1mBRTABHj
/I/HUoqRXbQVXyeOdmnOzcSsFSZL5UUL6YZ6oSOaAUBye0Ce8HImH8lcjnHMjutD
L/4fduIUhRoUZsqBIR8D8P7Rdv4Q24p48h/rs4SHAKbdgBCGZiEhIT8q6h45rRU7
1h+mzVqjl3ugZPJpsuC6DUvxgIhAqLvl6OkvqHjHajzyQO8f9cSZONPcojabtUKE
/77u4UWGrgKiqqKANmdil3YHkB3ZCKC7EVvRNw9dY9hgntkpGTD1+fUq68gIjCoT
fmbCTMEU0zZoqHdxyJeGPXUvbcgAI1e0Ppz16bMxoVh07xfyp5vHL+9G1dcwGdRW
5vJDie3KSiV4gXdvenvUNBAlXwQKclkvpH729bA1dQZJeW/5TgjP3iTaPMoTUUcR
ttp/aFYI7gKQ33jyh9Bt+uvH85Fm84ocUDAWgfIQ3WurtzW4HQFJwzfpDxCNXSPg
9CesM/mY455iZXAwz58aJ8ED5IPE+7MiyjPXlcbn7VIZiG7RJZB4t3RAUumWnjxO
g1xu8+9K2qKHsfQegnRFRTAYJHPDFyOmLV505v4RWEvmMspe+SvsNHNjEwaheQyD
Kv+my/RiiNVAfE5GmuoDzzR+1MVPMTpKP0ktnpvycrvp1J9ZDdjFzivN+peF53Vt
gfqa4uAQgV6pblT+c5IL4k/4RVZ7mCmr9GzLCiCy/ULXtOlm+OI5dqv22EdF2SZT
rt/ma3qd3KAK/4qWA9koz8JyEs/ck4YaOMP/JPY9aB4MKkabeE0TZ976zsP91BFf
qNeM9pLahtwcNo+SVm12FRHM1wFqJHseW5NjxJHuXDQtL0U3+IKe2IlIQUNyvsEa
shltnjLyjeVJUqNCWnRjMjGN6MKb18DGWVBNrmfUMCf4fnXhM7dxLAiiA0hbNhUu
1zNc/GO5ATL4NLN1TKGaVTY3LFw8KxBrI6qvjSHqbQz/hp6YJWIXV2kotHi+RHa+
Sp8vJ4ij9MGiWlV8tPG4ddnJo+e1ILbSEaXtHK0Hkld3wbCfM4ziRMaoqzsgclPE
5Ax7L5O/8/dNpQKvfPVuvmrxuo8QguaUqE1cbaaj5VYSOAOXMztVnKznO2YHceeE
RSOxjWd5Ew3xHurqirDvgidNm0tb8LHeGIVL13iaOkpfZ1Qrp/xdibFkg+GecDdF
sUYRpK0snDA4mI0HkTk1bIi5oSSoYPa2hkwyaTSyo80vWjMXoST/jykI7pa60EGR
4yrJYsjDHqGP1u34QYlY3E3OsNHNoY7XsceG7n7z04KpcrcZUYMys3rNVy5h2OfV
2FnlSjkLzz0MnMIgAPIbqa7xIh/gEhNWl6kaG6L+SMbdWZD+41UyOFdGX2gMQK7J
a5s4GOPGW8B33SfCfArifU6mbwgKGMpKtBnlTyUhWN5YPDTrTVyauf4KImEy9/CG
mCVKmxbcvAChbjxZlP27CQP+aYpU1jbs7OyxLBD3kdaHNfpV19ZZo7sA/gdKipDI
xSONZaLlCLb+bE/iof3nL7mmG4LzAKbuW44n1k9riG0kQOwQbfnXc5f0jxGK4Xuz
zs83bdoBDu7Q8QbadcEjHjmnlse7ZNmX2AUa+/ZgY7YQXaCkMeIuo2NNwXukC4e+
xtLe6Mq7ZHZiW+F693QxisL+Ulwir6g5+Wd9WjDSt0bEZcFqlQqilfFFQi/Pfwa5
glMpnX5rOYtC+6AbHS93JiuSz5yETBOk+evARDMAhpJgJ+K+WKzZ/BER6s8baDj7
hwrjR9KT2ZDFiEhBpw/dYRClSSJxl3V4IjvEZjz8CKbi2ItR6Z+GUQ+wjLVVtyW1
gAwh9RAwaJxLCwy/pm8XRbb2VikMjTX1Xxb6LefaP60Z1OoQsBWw6rVLp7k2J7Hj
fuqcErsQElqaqfqlrGCuK3Kh8yRbsil7R1buS+sL6yekxBiPV2MMhS7jPKeLgk6g
E+663TV9+isWX3QgIoKXNkJOHKcg6BVMVJ5XAmyOBUZRvKTFMIArXBPatZEAKBzE
VNEXVZTqSf/C8NPp4NT9KRhgN3egCEi7MU6wBcV815hCAVQjivGqZhN2AAgHI2ck
mAyqRmSEUlb16KnTyu1fCPqynu0xq0ufD4yXyQX3hClWJkBR+4e/bISlpSSm6H+f
81+/EXpfBVJHw+mb9c2eKuc+ddGVWgxlXvXkyFO/w3+hgW4kvYvSHQIQqrVmvVfR
BoE1bppmyN+BlJgZQXlSZCHBHrF/4jgb+UNcYfcobhPHPYHK6rvif6gMUXHm78RK
2BjSwj5b3QFzKEANsXC0wqEsBc4rXBJRuYVeS9370lW/x8ruKLRULj8XJyUTvf8G
0Qe+44bhwT5Ph/Sn+IzMUikZP3JCT0NGjbDGFOUmmw3JYDfsRUmOpd95zh7Ne0xe
uELVxYyNjErGQZBuK6PXvWgg4gKiOpKAm2rO5QwCbTDuI51zazMKmU/PPJhi7Pz1
l9xa8t4mHrKLsiueEpMEWGYLwfphJlnurl5nSFGakWuxi+c05NV4LQ9S4yRJ+nwt
B26suPoSYFKOTGzXPAtJVJoUe9AjEDHk34FsoPRLe2ZH40yODoRiWNZMb8Nv8toS
ZATR47tFOmFRBfFu5vIu58I1pG0qLsWdcSnJJUMA0Z0nMBX0iu39rY53h73ZCJWF
+SksVvQEi2fWud2rzc7UPVPgSBUIIQD7mbzNQfuj0Dzj8pBwZd4tik9MB2VABNtp
XQulWEx83nbgTR6hknBbDFxsVjLY1+Lg3O//sz9KtthRu/H4nexd3LWftPgpkjzJ
Y6gEsu0q0fdex0uxUH67NQI6wwJMIWWKaIDmfTNAsi6a2NVnG5BA0XKysp8j1C8k
sqEXT4lTsCvnquwBlR69PA8Fyqh54UdUNrVIqjHG1XiAG4ljTcBTXvqdndnjEtfU
5Secpuzt+Vw3PtteHNA+QPbAQK4rwEZRNAQ8bBS2q1RuHPH6ewO7UdqjaqFakXgZ
3IMKLZDCYHhL5X2FgIEtrOOFtG53AGFjDv1Ugn8b056PBSLlzEGELaDptipBVAts
tgqG84FSEF00lG2/YjRjNT5AZB55DX6nRSUxir4cGwBB9OejR13rFb/PDIJe+zhB
UDIeqxG0o3LdrbJ999oFiQZcLNmy3YFIMbbS483nACR9ccnS/nuVEfQDIYRb8SMx
MaA399uIKpN6edNitIJD/DiKSmzM/SzFuQF5k0otuF8aLvyeR19MJJhgPbH0GWrO
znfsNrthA5mVtxG2ZRb199qUGuFfszEXXGTl5xjakjVL7HhQGne8+a7gikNYIG9Z
bVw9T8Xvm8oa39IUPkFVylAfMaVdFwGlYSbr6NOqqe/JBPnYkdGWB0YrMJaNhXXP
bOEc7bf+U3lFdxFrqx5iwS3ShXIlUOaHXJRdFL37i2k/0z7gvmkuT2j0fm8xmrUL
3mApyPWtmKNaL3fW4lnv0wvcksj2b/gZm3dFyLbYckrOg2nIVb+DCWLhICOmW/iZ
GrzuU1S7zPuWXB1L3THLyw/niMLxcxtusOOLRzld5EP8EbdySUtYwF7lD0Lu4KCZ
NJ6dChaNXgArnuCJkThYIuK8YagEuxq7D2+8MHxEdmUbHvjie5LlXwz1F8aIYPXD
v6Qf9jHErDoTFwJdGNQ8YsVGZEmwrbRGYnOdyWWKeZBZiAIw1eSdhUorNnyRXx1T
IIw+OytucJBMbu3K8cWWwo16LstNFfGNkggVwOzEWacJvsJ4oalXSks9BogYNVI5
+KopAWzUMobSP9CtXX4HqEJ205oycGLiNPK+oj73QP/vmGIp3HjrTHl4nZ/zidGw
oIIaQzpiqLkQ59c/ylbn4RQ1WJt0/8w0cpyXKe/Gi/TCpxBqaFwxQti+JEHJYbqQ
ZteBIB3Xcy8kpdFlpqEkvvOU/aq46bclJxz7xjjHG7c1sUydiF6LPlWD5lo3yoye
VwoL0ZiSdu596kSpHjtYuSj+BkNl7KFy+heDXrEYOr2/HyxI4G8cc15dmcxiUheo
y3+QBhobRJzgnZtWE/UGw498MlCl2+M7fdsr8hr7b8wbeZe2Ly/TxKVWXHsgLC6/
l/Su530DY+DX6QKB/rh96J7xJRKKchYSAyMz5eEbv927EasDOEkTzufyfKqbIDev
GIHh/S2bwN4QwK1jRr50Gx9IZKSvKIRze53NSuyUasZkKvDAGBj52+NbkSk/1XqM
d8D5aARs7dPO2VCApR8alI6/gfSAVTyQhIyGTKfXbPCa+Fn/uWrtfANmNM/lSi0w
Hq9MGJ9YdtC3COELkqk7hNhhVWlUJI2Sce5uWqOC9fSFAiPlALZ/rQcOlH+/3lvN
dKaKQcEiAPY6zH/0kMA2CD+kc0phxeuGyhPCKFDorrsdQzS6noUfxDDLdA3Jj+ba
fgGGAbK6h14+3siM6orG6Nxcyij+CS7emwi5JTFvRI5nIeGsR9dpB21wJUCjj+vf
C4RmYk/GnX6ycyYHXr7eHFwgcHCSGy09ziJXNxRQCHB6DZc5RFsCRzFNqA/n3suT
/Cwra/a5bAp+v44G7FcwHDLOng8GRQyO7dEXLAglE5Z5UmDI3O2cbfvui+izEqIX
NjT0zOrMQZjuiebLco5UVU/7nF6dVB1svpJaJUNm0BfPjadGHhzsieQqyeFA9SjC
v9FpcvMzZY0167+qpGAwB3XeGy/nJZ4/StPJeuKw5jLUfT1t7wCqUFdc5VHz07LF
683dnI5a4Q4KCv+ghnj5lIRGQ1yKkRsNvD98tJpKbmJsSF3gK2538g0wAaNWV0WD
4+edE0gUgncTMHxGzXhM+uW6MJuFUqcks0u2E1eKV+tVIMuzeggJXrZ0Nn/OjmkB
uMcu2tN5Yl3Lhf9L03Pbl2xN1pNPVO2+TD4D3AMOyr6Ni8VQnLMnNKzqDf4IMwOh
I6I7xNFHmbE9CtNUCt+KoYHJVfGSUsvkjc2LIuUOB5Fzf5aT2kzQ4ONps0C61Lc3
VGc1nsc36rs1bue+RGrLhKZksqtB+C75GHkK1xjuBhKN1BAJIzNXPbgmQjFSwnlQ
gy7Wr1HoKFCadxYLbCzs1takMKWhEEfSkzqrP9PJL/PCthjVmkXWL4pUHX06ERSo
aqiBXrDwz6S+wWRrveSwP4+/qWp5qJjoMG2cYMzUQa03PmROsSrur3kKkcg7KDpM
kuvH470m13lyNTY4MDHF+xTwnnaDYkfAiC+H4kAO01VkILyQD91s5thk6LfUT4rD
LneDyOVsQwIxm7JqMSOJT7TvX8DpfVz4oH78hZM2ROCPvOGhvuRqlu/PnRFtTcxf
WZZMKZwKdH+OA3ehYvz3R+FC42ff1hS94oHmb7bW6/L1Wz8giGwGWzPGqOn3xf7N
m6Iz2LR7LmxBMFU5EJ6kvhkR9+q/zKs9a5354AUHRbRpqepSjm26pKMwnHTIWOlh
oygiTdr5ta+NEFwY9jh/09FyyQs0Kggs1Gl61N+nhno76rwDeNfbDWDmciiiWBEA
Gi4GLD0KTwmj1kHEROb7n2KJtqv3zxwaSqckTcQnFfau5ibi+L9WS5WHKU1vBl8P
Ff/0JYq4cwIMB515brdsrQjfOwQ1SQTSUFk0vjpVac63qyboFb3xecx0Li5DRPOm
5BIjYWEIlhuKgu7ZBDC2qqmNm234evO07gqkLicG7vC+inP652Vlir6tWU9c4xPK
oOHKvP/X8hXk2O9r7bEqhbMgbP9z9vLdY/ChgzOfZmagTMK5+PVCpHmoyJD7aEGZ
LjFf4/OK1x/RncUXinD8sk++rIDnfBXrfqgfyNgZeTutCcdddag3nPmnMvYeqB1Y
iApRkiiiZj3Zr8ACSJQCx6DPdBbPGFsfC3SMPjDg0x9sQn9Cl830djnT5wAjMRn5
EZI9BnjhpuhQY0Ybrxgplrf+uH+7s5RrAQR8P4/C0Ezct/eHjPEzsHY89nrhqwu7
Q6J9oez/dQYxUWys8fH8+7kYFEcvAgPrsss7z8m5jc1T42qXNdiJjGsgzujj3Oo7
MvjZQAlZ74Wwoqvx8LtbZ0XQxl2GB68A1bEFEulNfBTysIYpC/bejbdzkQI+h+bL
Y3xHb0sVzfRvAohXRrgQCRpyqr29vIj6bFLTgvLof8YXKC4z4u+/iAr/AX1WomJU
OaXPp51zqsqSM+essmRpccsxS2VJgnLyg2nyW2MqqfSVSK8uXVtjSqpNfhg0iQXx
QSu0H4hWZIc557dZjvL0Id+CiUrzv6WT7jOtkxVIgr/GH7pEUPhpbvUlurVehOda
ZyPeeAtobq+xTHYAPXJKaYrJhzJ7QSIAMssQsuWiLSLq65U0Js01sdudsAe85N1B
nx4jAHrBdV1S9z0fq4tpCqYrzVrSOxYXL1qSpR3WDBy4+5aeUrOazdPhBueSSgSW
rvT6efbCQEBf04lv1LY2HqMUjAC8RB455zYOzVTVICpMbm5ZbkGQmesZNlkf5yUd
ERp9mWlwMyYz+RX/0ZuTGlqhqJuZ4VBqCVZTQRndTV2uyLgDYgUFl6Px7yRmCuCf
WwTUoV4sLRO3oqy3abokYnp0zt2snkVABssUW4hL/g6N0aOhqP5h2KDYr7XFMtdv
HVVMn9EWwGb72DDdGu9GdtlmWwjSl9IxDGtNoVzBnhtCXdAzjwWCK7/6ik0n7yHH
3QqCJEZtzO1piw7eBeLxl/INbZqXUkrW4FuPQOPCBLrPvMa6Ph0XrbbwcWLTWzZK
HX2E30i7JieN1XGuxQ3EuybNopUzMzPQswJNAbVeeSMSeEOHmzMEabhI6VNIgIrT
EXkkgzURllOK0qOyj2mr0eg5/sHgt0GTkU/7ze9CxffQmGynq+Dz9e8ZqBwFdjw3
6cw8fI+HJbDHk59J5QHnwkwm6P0nzd9HoceUVRUuE2uy/xwi+gAzFq7SZwr760tZ
8xHiYoVH6hcX8FYT/+sDcyKsejDPVwsYw4viVEHbdnRFsA0+NTGPxGniCVGhQKwQ
Ks/W4rIa5c7MhBgqwgUGlSDINrSMVyrA1hh5NoA38Zd2a7Gxrh7IQpZa7yAY8nyc
mbqT8lB28hEHdZ1t+bwyLflnsClwSDK/2rghcqu3oNHDaLP99oJKv1ToQCUsPgjU
CJEcCRiFT60iO/Ivt78YxfkMsCSt+sPV7DFwf7HFnut+ucG+4K2pn++Zqb3ea/lN
GV0o0kZLWFMUR6o/R1DiKg2H5sICl+Nv0DSFprmEKzgLj4kzzG25CFnHFm8ON7IF
vRcu04/kX7wYS/eTBeXbJ3iVXcu9YSpi9P7oB07KEkRQDyYFC7t0hz6fh75jeyny
fXJXgIamYR00tNZWf1RKRj6FhJ7TAbW7baLbZ21ufUnT35ctXRSUD4QlbNKOSaXA
hnlBM+0u4/YMRibznaLei1Smy0BwQSLQU2VcfscbIj83Uu1PKD2LTd/smUqpqYty
wNYuFdrkoVat+DLJsV2VWcIxdxiNiCyH9/eRqQMn/me8nSS0DJTO60T1glceBlpq
VYzrMsutiR1OIgnLcI3M3teZyPoe9/AW35E/+F+kiWiE2JXi8sAl0IeByS28x446
4gwQ+R8xtdMdKcdiHdMJAQcyWMg0E6iihTD6zng4eUK9OBjV9o2qliB7tUUecF/i
FaFDvjqmqDdBmOL0+FNy+/QwVTLa0Hthol4IIaTzh8lIEsuNK7OgPCyhI+w75SML
W1jk026fNCvA4tiqKpkk5Uynpt2DVqhvxKSo+2QXdsG7iynjdgPaIlzqfUwFdgTc
evsKfijGkwq4NjPyL2PLdF8hmYFEBbeJiGrGztkdtnWyRB+aOvoPAtQF1ssSDapW
Hpsw7xZHEpPkrmOTWAtTiJZ/ZRr6IMJ5hnaX1p2J8fyO/37+eRmX+Ge+Tg+4Httu
3TH81053l2brBcW5gH0mAIW4e9Lx0VY7yawrcqo0fhpdtGcgJ9O9MWlkzbH3OV0O
2/X5Ce1H5cpTyiGbmH+rfxvta9b0R0r2XqrnpbTlHzBO3jbcOpkkKNo6tSTDcHwE
kkfyuzb/6w6s0wai4xlfn3dNHJQuuSG9/ckgUKjUqnzNBX/EPaKPzVosZawjvXti
7URP3Q54Y32L3KVES9iqfzro+whj/QXLBXELtZhCs9NzCCduM9zIdb9X/P31PZSG
w70ZdPb92RszZaAO0rhvOcrDLF1v4SanqA4esdGMoazMldwXIYZv0/0do16IYAov
qmfcgbLa13lerwBnBB4dy32YFPtLOxu6/JJHkNLVSyadqDbNYOaRa1Spn01qyIp/
APYgXbpR632YQlmHOwavBlszS9P28LyDBCyYq5gsXeM4igGQUgsGWeGart+qgrSz
8eRIHcB39kUBgADzf8TneUm+pjo0vearO3upBu8skdwAIfmMhSuSphW1N3z+WubP
PKsQYExk8aLX5WGGTeQlWQ/s6Um0GCzymIYNu+8duX2QGo67X9GKn65ANcR2Elj1
2mN8TDKynR+t9RPkt1njjNOlrSzqDAcjPzfVVdDlKrsK+COsk/7uY41SWdsNAlQh
7ZIxh5Ea1muJF2ZmQXCZVoM63HZpRUIBZGxMtetpkqufMcnKxWm0Xj7Ed1eBeuFO
wPLiTFieTpB7wS2rxxjHd2jIi4XwjAez9oPprKnu5nrx0BkyfwX0oHFJRlxxFGRS
srs69IN3hrF49ta8t6Q7Yq3+QswmTBnQo37YNRr0aSUnB47mWFwiAMPKpzhhZVvk
6TGSvxQxPXcPiPY6etJ56gde+eM53vzj4SAFSOKlhpor5cJtIR1XGr0zZHhtxn3x
MxqbSJIxGwMoZY28SAWUpDhrgGy+oPAnjekglRX1dDlU6vgAwssQZbKKe9elwQ67
CkeV6D7uMtsZAllMpfdyCwd1DzkEXW7zKuPyBKYamIOAaer/wV8d15jdn0TWhIGq
0k2+sKwgo8DHbNyKxsZWt4xt0YGExBsp3OMEx8VqE4nK/PpVb8PLunkAiPuzCqSp
ZJ55e8cpe5LkcR90fwOZ3rVPWAc4qa1SsWfbcVIR+R1DJtcWB9mu7OJDIrkcRQSI
J36Wl+1pe3RcEMHHAq01qFJoMBICpVE01h//nicLfhbP3zEns3z4uiq9DFkf28An
/2CGnvgjRBYvE3vSYOnqBIx5xX3w9CV0AoIod+cuWxaOMA9l34YugbSs+MGCkgiD
4BLwSde5oAHoj20llsMsCALIWigBifOqYURzQKCkU0AmUcLfyIV0/v4W6UONW29b
N3QmALlUeIN6WmHpfX/l/tRbMAyUFrvjQbopiwPphFyrKUX1PShHXkRSy6DtWgMR
oBhSfyH85qFOkBlB9Yz7H5J70TUadbeeYU+aUlR8YctEc1w48RxzJqidd7oX9S7x
1NQM86azIwhm2EwVrU1AglXtrdyXIyry7GZ0OekCeE3ZnNOkejXkx2lxCQJGpoHk
Qo//2Z/oPqQlsvr2ePEkeLhkkt9JcFFbBkCURkpnQ65f36ypCoFDhFVrZiXhe0CW
W1W0XTSNGot60LxN7M6Bq1ocJvzKkcRRnCL9NXMsecY3md+jHDOttGbr3bAlUEg0
ymrXTIIOi0dIsNS/iPsmFIwB+PY9lC5CCqIswpI7YhgufTgPRcndh/DHpdrioPn5
h4NjsBmPzSaXlsOKHr7YT+HyhNYdueZm+0wr8Fawj04JAZjy2IJU26QL1KgK5VJH
Lx1dkG/DW5o59zhpukcvcLPZNaIX972s63FWIHWZf58S9gJkNElLJxZBBRdnU4Ij
VDF2hefEc0dj65AMtUYcBg+mlz8gYzbJfRkUCTog1M/obyzZj+d9hisSexyuIPtv
MTCO3dZs867ZltfYpjXKwePzBLMVYA/ykpPN5jpUJr9BnVEbi0JFponBdAhL8JHp
W27twarJAnjORnTvvBlOd1SMCtg7ks6AQPpQXMQqPA+ZvIu5GSfczxdhlhm5LEir
QBVEqNT0NzLRLlyjq/x6ktbttn+zCCk15zN+gTlQzXOA1Ndsooih4WGsA+8WOCum
a5J+L2OP9gK3WVWiBHp63BfSNRjB+p+j/WYn49AcVzWWJb4fc5OA9Pc/MZWZGWn/
mMb8GcmfKbjyDdEhgURXm0fQj1PQeU3UpchvJMpg/PvKYHZgQtW4CNWOsd5j/b/A
SD2DJKRLN8IMuHuAc6ArULBZxgsgsQfMcrRIBqb/o5x16RYNSCfob62Er6fjLDwV
T6PAQT2ZE5EHWOe4NFNqtfpVGajiTZRH/krzNP42OYtPIUtesWykRf1wwb9L7KNb
nveBJRSRUYqvGrAoKak7/DhwYt0NNSJfBs08+PPkjOirw3o3Rb0dp4OwwMjoLdjo
ptgqSwyVITBo6xTuzAzD5AQRdXiHJyM1x0S/nzYKpdUZygigRJTEF4IYskgcY39V
0s+MP1ZjewHNo5HQtxHOYpRXtQCK4IYSNcwq9+Mr5cIXpbqyTKNDDrY4J3JjKe27
QatpZFmN4CgZQyWURnjMCvYLoCVcNP8Uf5KVWctHS020vC2FwjDaJQkDi2iO+3h1
o9xS00f59bDoa96WQduaiGsidMI9ER7EbJjlntd20cOqpDAwHb081vS0ubEAuOTw
7YusWMcCdg4Y1qScdqCWZc47XbVUqtCkaBuwbnRFAa/2qFShY/GQmYM/ei1PP04d
SlyaNG0XCsEdOyX+arCKrm8LMONvVSMShEakPNJy3qOopnQkdDmi6lj0J3QC+fqk
o4YhcIEfHYFlYA2jP9LaJS4U3g0SpuOrMSUb0mzJOm/zhsnHle9C2qkGj4mvu5kY
oLHQVP8Z+Dzc8kY6T15WQHW40yVmZAGALsMyWjcZSiHPE06GUOPqpZ0DuLh5o43f
2QFuDBEbRrkWvA8bpfqUb5osC1YPssa032CbTfL9oObO5+qeSEsrC2o0SnxS+tQD
rIlMVh0WEh/P7evNJM4/2SmU07T7+sKPXD7/Sbkm0I5aS9iZjCH1fx4f/+mBTlbo
nMuPJDIg78AckzRYhnebmRn18Ts8uOfaQyq2a7I5r/V+C1/5jz0Q0BOV/UQ796XN
tl8Srts8JB+kw8GCTqLy1b8BiHv61dJyKEF2X80Lc7QIUadPSidJH90v8tP5FXLD
WlgchzW0h/OErJA65GNKmVSnY+s8aKBsy9dPU10sgpRcC0I2rZOch6hf1TLFji9v
lKD9FAfpX32VOc1KUqnK234+ZlAqXdkhlepTPryRwOIovyGxqo0G+CceYCK447Nb
euvJcruNRKhrIGCObu1y2ZFQY8jgLwNTpHlkR+rJgucYEUQG1EYwck+pFshNFUj0
ODcn0ZyQBgBpRtqQ4bbTePe3C5ItvNnxnwu0AUgoQyN4tCnXpgfsJlL7yz66ep3N
DTn4pINQIkhi6C/SN1BG3kiadPeLkKxBRsfTaiZ+/w57bvylzvLkjSvihbrMukIh
2FQLQKBLEXxaBZjq6H+cgenZSTY7bah7mMQyMXyzB7k2NYW6j1p/ZS/jOyb8eSGa
GfgfEdSwyDhHizRkRdfIs6VP+ipV9oDRwQCeSoUDvOyoP5V9SuvC3KVKyYL4eTje
7L5esRFw8/wBYbls29XbwYYRUiJ9BovBd/I76usWB1ncMuZjuidk0nS1rsOmC5Iw
ZY34aZzyH3GU1JU9XroRk63D9a5tWeSN+JHoPsjkw1uR7syGxE8lGvVJw0kedwnc
p52nARi7ya97e0mKkqsPYk32a6jvmVyOVaLkRuoDCUxRUX4Qp5nhn2ZDaHdm49QP
Figk1PcrNQTNM7EjCdFuj2A9Y/fqyizp7jOQeHXlNa7SVIcwoKycOyMSEEHlsDIt
HfsGBrbRN06yd0Fxpu97r9DYncMUGNppMVfwEf/hpBo/4THIUNXIbkpn0m2HUhpf
D7DPJZImyeFgwsG4IaClgmuKDRF9G6vIWW0i6MceatHAnzOpDEo5weQBtOPo9xtY
Y4DRdEySXc4DUTXtCyyg2DLJyVm0d4/SWXG21ueVYJ+bW609OLcNBe3moNdynwv/
6Wer+cUhm/+xhFiB1Hkf23R/Us26KjoSFwKNbaiTPWTA+eF3g05Plf4Sz6UGJoP0
QbBmHgQMuP4CTei/KqKrvSgQFnEFmS7aIU7EjXkSzQYo01WuzNA9pwz3OFqFWNiw
IZHUauuF+fllVpoSzoTdrgsCqLmLbcOyHgXZnGwadps0kOsoNjNqrzQfVGfkY6al
YJDPxEMMM9rSACvlFa282RQYrUINF4LEgXkDgBE6EUxWUrAs7/W2ueohTtI3dVAq
UzQonLNWuOaFS3DdLBK6ZiJD9Ho9+rNjDl293ZdAn0DZfFisS0mUAM3aHrGWFqb7
F7j7t7oYe69oCxLsKVHFonE49ufLoqjhE78jaKb0gJyhVQc7EE0/ZgZxcSvDAh1V
BeC7Fac9Fgsj5NxMepfPKjn1jdnw6Uen7NbK16h2nUfPjMu9L9k/zvU5vd26WTB8
KI4rmyL9S/RiB0IYLU3Y66UYXQf0bCqJ4rDOPu0YEUfTV7yupCw3ym9fFUbsJUmH
Yqgrngqrd1npW0VBTF0eI8x3WXoqKCdRg+ntrnw7+NivLSGQ3PytZ8aIgiSM43mi
qVdoKj+6HXm1IKlKCCQ2ub+Jj2dlsN/vdizns019V4i92CwbPoi1CI1vGzkxjzzK
JE0LdhPUAjKtOYk//2LpDrUHjDe1Z8gRipLwgIv2THC1TxR8961UaVMW50QRUp03
uIChYqhfyPcFdM8T+hMYAd+KrOibH56TkBSM1Auze4Z7yCimQ+PNa980HhK3ghUF
cXVmo/IPMle5rwniiGaVKCpRulCobezIyn/iLJ8Bvb9tUpH1xDI7cOHHbinSQKyF
FYI4zOuoBuisp3XywhrPI26hV1W14wwETUWS4M0eZT4UzhlYm9CsMzlEGf9ZTghJ
sqbYzZAVE64dc/dH/xydhhLgjANHDXoz8+FZcj/h4JuoCzrkVrX0dmRAejyzQjo1
aEipGOtvUjqhRCwT5ORjvbyWMUMFoP+WptiA1nnj7b92aTm5HG+OPisevHtESRHf
HUcwqlcFe0TG4mxuum6JAECdwFpEcEvhd8yiGZUBASWlrmm4GPO4qoALiYj9sZsp
D8M3cVmCDeZ0k8/HYEAcEqgF1ZA8VgTj3P8FY8JxkO7v8zCgG6Wq5wg9SA6wazYQ
K6qMXlxsNn1ct1nzoAPR169LyWa9Mc/tXiUbqWoxfHzDZPzH9Lrdb++0886o/Hi8
9OIIrZJV62mPFE7h/uVmcX8L3MJzijmHAxWyf0rWP4FaVLrhfYMRZN2EQisXIJrP
Vc490jYwiVfBFpCjdEzgpvt0uSc4RI4I3E/Y4Ah8UDdWPN7mCTb3WqRRiQ3YU3pp
5qO2d96df2GYmmU/1Fo7bmaMBD1cQHW7hjnc9nBK25bpDmc+dVEncNb7JRmtN2EI
ulTqCG5bfGYJXvymi4KTgm3TJpgHOrH5Nk7QUcQG6nYwkVlJ+E4Ychq7oP2fXMrT
mQFPVBQiAArBppTX4wOuO3x0ii1fFjYgvZ/vK8eYKwmTcccBXmxFD1xtLTv9h8v9
BGs1j8V3q97pn1cXKE/mtjM7yrJSmHeKYW7vogLT/oQL8WjwUkRO6mLSuquyivM/
N8FyuB5qWlfqUKMmT1rI/a9P3U3G0QV4WpCDOq+HFzfs/17/0zAh/0pqxauIszJF
vUa/isPFbKtOEi6Xu4S4AEfJy4VNrrP8Yqs9akh7/2rCjIPQL76jNDaQqDUzyAPV
z7jgznl59552vp2CdEvjt54gpuzbrAmMZloFPg/srjbvEmgnzJ+f8pot4LKWkRy/
kyTZGWXDTFUW6m37vAR1GjMA4zJkjAWJ0SbUPgzchukYqf9thHW866ia8RvjM1vY
F2xef0mbB3XtK+3rOB/e83dfHdvAtx3HTNm2M7/afL7EeV6rkBLPGMpA9CdQlv17
0Y+N9X2FBmLvyNEPTNKTSDvzbnSTlIcEG8oZLdT/7YUggp2wJdJslLcKJFDXDfoB
ubU+Lnx6bqEaU8tJRQ0zEcX4WbdRobDLw2uNqK1smeuXips3+esULkwVI4kVhHjg
aHUhk2ohaXF6VvGilujLyfYAqQOf7WZnkLAO+ENPerKQZ8kMzqf6WwsfXm1YHj62
c9jUxEtxsXd2/BonAvnLOccKhPx062y6CzZ+dWsVjHstmSgwpGTvyjXkoPGDLDR1
K7yuZFdg10rxOnmgF9npNvxG/dJQNaeuzCCgZ6Se64mgHLMlfGK35W7kY6V/82rZ
u9LPxw5hm7ZU6ZWlV0yKoWdhhKKm4RjDacKrZyWAzd+7NIs3Pay3nyNBEFzORIRd
m8aSK04JAH3CbGmhI+kDo5/LFEVmBWmGRse8c7Lxe7mR5SBEBEi5L9MObdAR5ScE
2/3YyFjoNi2vu6QYX6b7GwaO7UfjMRyiWo8hG3u6u3HWPRfJyaUgA7ZqDXiol2Ru
5W+7s7ayp0sgntkIT50fBa22kukWNQpK2GDWWd0rq/U4VLocEoLVFyQZhIwc7+UF
SccTKuaKWl7/d0XmXdaLctWPkM09lKvA/t1vtM2LUvDn9PV7za1jgmAJSbaDpDMT
CKQD9CG/zD/ablS2BW1qpcksSuvguUTrJHW6JJ9PmHFlgx3z2noWhOAOjjS+UWD0
8EqbkgglmDI54qulSQjXfGKGHmhMGZj4CwdOfToToWZ5facmxrHaM5NtSBx66TF0
DxVWwnAOqrfsLnk7YRP4Res4YQreUctIl9P4xybUiBedSzWxKnkus1w6itNguW6L
+K9Ggtn0I2Nk+4sQ4Wk6JVb8aLKS3IHi0EacV4tyrilzsBzXNcp1kqMTQd/6bGwv
7AiKeW/MuylQcTs2rZA5Rbcffpi3u0yTXfMfcG3pz9zUtQvBKm6o1Ds2ugeOwckt
h5BZaMosaFfQ6xaZQy5lNHRJ59VD/+REoJtHi+K4/G0pttuz81PKHw10bh0WvkFr
EU5xRoVYpP+ngtRy6T5oKhvwmwCpVLiW5/oyWGUKBWyi/8Edzca9AbsC0rXSkxxS
/G+qFVD67fetAcL3y+F6J3em61FbdkbRLKqWL7hBSjk3+BUCL7HktcM9MazxS0kW
IZ/VPx86I4a7/1x0V+7jt+ISbRmvsZpOaGyZ4mOkMAhrnh8hAtShcBdAIJDRCQ4f
WqyEsiDx3fhDO+ufOjGGlVbk60kMuZNcHSVfKowvulEVlQ6UWsBQ8ja9bgGYPYOF
NT6sIyHylGo6TM2eehUUfgpBOTdXUBzZQSf30hl5fPGaXzmssXLjLiLOn9VWLMl3
plNSCUu+gfQ1kYLauJ0uj57kK19PbavOi98f3/q/KeQ8ds1PL/+Cqs9nsO/V0akA
h/vsrD8LVbB6fyGJlpLSNVLc9NgaTL67/ZK6UZKeybtJOx2n70iNAKe7ZcaxTVnC
NRWpsML8KvWW++bETlniFXFBz9zIUGmycpc4B2cqogt65P4RUpOGF9yczHMWUxps
M9SSz7pENZ/Wm2FEWuLKU1GXZwl1wFEaRehpGNtzEc8XFE6YosMwKk2Zr3eJYw9z
DVlfvVsUZaQtVMchaIbYhsPSUjI69qFfGKr4ehn2cScNuOf6mqEnUXC69IaRutNz
jTsruemXUFMLfX3cH/0rNDOUdCqirJ79ix8l32brQKeGeb33S/nhS2onJdZamrDn
AEn8FlOhEetM6ODK3dBt/eaz8HS3Lq+fq6yN+5LJJrfqsLihW5NJ29+wjoeK/HBv
dCPN8mXeJUhfj+LD/fA9Lni/om8w6NDtah0eMtexc/8w4K/D+8cqZPR6HpH+uATr
4XdSS3KCF/nk0XUy4xgltjtwM33y+Nc2CnXV+m6Gm2M4uoktCoramyZ9ir8VFZpS
IkGvkpJkV7DY8+X7GKHTbwLdMnD319gCD5bK909pKvD16tVF1k7131tnsrvCTvR4
YWAL4deujENTVQHasQD4X7CMHEQeqRlbb7sRHN1FDDujaelB/ZBs5ewMg1P4cav8
5/RVHXH/7+STG/L/zdMFCgWaNviPvK+wlwFqZ+WrehK656sWqjcYdgO0UzIAzXEz
AWEZ755MfKSf0Pmkn/0gyMkKIE4OLJM3ig0tV1IC0ML9TreISqSPKRVGEbv+Md5/
Rk/gg2vf8vGtxpJxLD9FVxeDPN2a/Bb9/jovYJ/iqCU9R59Bn1kt7Xv+YW26/kr0
4n84Yvpc3N7eENVFAlp0cE61i+kTYc0G602ykH6E0R9IPFmgj5YXZWE8hg5+ev9T
19C1xeyeCZocJvvA/pj8DfZMY0CELPeE0s93+oVlw1WeDUtPMgKcsR8VGO092f5y
OUb9wIU7cVU0nQ9CDJlCk3zCzOWMI6jNIjbKOcDsaslZ/yZ7G5a4EMn97uFi99Sf
Awxex6NnJdDEQ1VFLcMXG4B5NGhtBLPVNiD2dZMYjYWbcR1jP1685sLVM8JAgsRT
2JVcduEgbGO2L6ur6EUcq5EITpx84C0NXMejp8iCIkE9eKg/1FKAWW9DsPEDovAr
eAfsG4TGYrM/sWy2Mt8WyZPefSriBjYH+7QxjR7lNz3iwy3rCx3+CW6Op1zOxcK7
01kMQasCOdNOOpOtvxLtC7Yber928C1X89gy5pFOAVhcaB2AbcGJw0hQRdTnT/5u
L4zxOQO2d1Xbxaw/vQAhTET8RSIhoF/QCP3BMu/IrKeYjsw3RGLq2y4Aqx9xdss7
hk5fXKxgtVKhLyrcaJY4q9kZE/Dbb6rmmo8/XsxIffvG8E+DSam82cJnApLmZ5Og
Z6DTR+CXAIrJmtkFxg0sDxOHyEQE+uHBVM57UnlUYWCp8ep4ubvghG7figRPwPH1
hkl7+w2BZX6JDLD9vRJ8y0Xe3scPsMcEgWJzW85lkrGvJfdJJ42eUzURe4oQ/Mzj
ZfMXm1Ro+o7Y30CFFwZAx/cHFYZn0KUIdUIHsWHMscwHDw4G2Q78740gTEOIHD3q
39rdMWaZF7EHsbWtiKdS6uEYmN6Nqw/vQAwdPez0syxrhPX3r7N40KbIKLBlOf5i
+QkmQFRYLKRApjMkTyL9o3OT22tjlTKRP0+XzEtdm6UZQtH6jDAS9nFEH9Jgesjk
YRsyPTYHF0J62N1Er6iioqloXZ/5epoBpRK/2YFdUioTom1pFt9nDOJ7q8PRyZ/4
ceGMQfupXMilvOElsRuaDejJbzjWNXTU/edD61G/7ivdxzWXNokT//06n7/fmXB1
Bj5JjHHpqzdQr9WfRh2i3Af1eO5jPrTFCKPZ5YC5zHIzrHc8KTHXi4O0vzJRrvtv
D3RGkjfHwHyVXh3CG8U3eWPnrRHEBozfEdmft+nxcP2JsR0Jk/4hfpB/IWD9jqsI
N6Zf4uj7pz0X67zKAY/GIcW4MD8iJClO8W4WZyIcwAPqtRoGXw83Cgfn+Tqoth5/
tZpf8NwlsnWmRSF5NQQdUd/3/rxDX9wvGsGuCN5K903sgwFkCpW/AeE46+JRjMQm
h77AWj+jb84hS7JkuKD+Fn6A9SlGAbHCf3piUaeFsSuBEA7N/LeWtUJOi1k6vy4O
+ZIsah/6UZclGS2IzVo7ct1bONpzvwUdYdZldAUTccSgabrB8WQAn2kW7sEQgPw/
A5v7RiBhMQDrDztDgtgp8knGSqMQ4a63fcPdZbDR9bLHzBd/e2SzsV/15VTcrPV/
uoQesJrRJxVIilBCE+TH6eFaYmRwHKYQ3rK5IiWvWHs/oFoVPrJ4mkWSL6SRVt/D
3Ewbw36Juq78/yGzB/VB2M15koU+1GdGgHdUGR9RKiRqCwlPNbnrowNvWM0wiVic
QVoAH0Z1ZAqCtKSHxuEv6+T7L2gQbd4OFI4TEbFaTeiXGZ1AsQC5cxOzwQWtVgCu
82kutSdEkmWdqwhS3gNehghTJr2wvEpdSkd3PZJoQ6otgDVLszs9t6a4AoMBX12S
i5h1eKYYJie3kR5C1P0a51HIWvv2tldbwxpvdmeOcY1Fel4QPh0b/GkGYGvkIpxv
fZyhhZcYGw4g5987Gg68v8phIygT6rE8U3yywIe2Q2zTcmLijK54zeUR7HCkFHbj
Ws5Nwfk7Dzt30Ca1rCPuNYrWiJj7E+cLz4p70NGQdi1Cr1SsNvxdXGjlnBj8abEX
yxTMgZeiMO7HybA10/ZKJAwyZCcgkhcnA9CqbK4OsiTTKNX3MLuSUoQkSW/ObEEp
H1IiTVdIfwzuBxK8W9eKqMdhQUNjE0qkr7zwTC+0BtDntsRmuW96Kg9IhX9YAiGM
eACLwSUpZmcJmVy/qt4gJnOidAcbXRwczDD1Tx0AyrkQBm11F6Ila8vfpC7MoUDq
kNJVwpV+ryk+aKUFby7cLRBSTUz3I88rsqXkGZjJvEIJgpSF0j3q9dxueHOSFsfR
fRVppqk4tDg62KVwxMYIPg3on4NV+EDpDGnA96cy+67+ZvVYlkAO9lmPD0Q3ea9y
ZsSn+Y5h03SD2+HNxXJ/f+Lh/4fpKHgbyEd2UrOqJUSETnaQYa2b0OkhR0N7rBXK
cpsKKYnWxpvmwEHLe3/ffcv7d6q1W2PKTqhWZ8V6E18STSPbb+1zjX42RkB0QlDt
4ATGw8hqpEWw5HIvcaRxsLpwt24ZD0ux+8c9rgqLYJx2ew0IK/SxOodzZ1JG7zwQ
guNN0bO1qFsVrBRw17ck+T9O9FkwEP8vzyN/2kv6trytjI9dQqG0XznAISp9w5K2
zAjsWrObgjKMIiA5DquNdqYyg39Ne8yRgLqwLAEeeELognNrUPQpAo17qInmrGxJ
uTXcUYiADoRkOkY30Ga6f8v9BKlcJhd3Q7aVukYReY31N5Wne5F+7gyazzpzGp9i
6Ci1gaMOVX356Gfys+jigO81ZzB7C9VsrMy1HfVKMXQKEGnVcxd691ccXbfpO3HA
7oG7yd3BsrwVv3MLvbfmCW6YEXkeJi79zFX/ebwBSZDqpzIuY0y6hRAGq8b2V+DT
sSPt5w23b9xV69xr7le7thv8lDMfH+2/g4MF3uROc9hTd6AGTteN6KnesjM3Yahf
+z9mcFoz8cPqRP2nq4cicC9Wfi8Z7VjILNMim4kDjV8JGap6jQ8iPXyJdaZBn9Va
WOadYp0gnMuaFxGGl3LwnlBkhAeV9rY+sxLt1RKX5cBa7+/BNybqnkPcVLVAFAMu
OycFf1x7ke9p4XLeuHAw32SD5Funkjn1ORytKjecUda5AMP6RJWhi8LmKTu18+f1
ktJJkrR+eB9kvFEitbo3acZjxQ/CGkWrAdtabgBKvZXfjIGCODKXK5+bk4CFWk+o
FmMLLMN2rUh2mRzcmbiqG9aknYufsThq1lTnsDI1l5nHQ7mE7fbO2hxb4THYj0k8
Va0MbtfkTPWMCYoaULQ0ehZrZgJhazF3XlAT34S4h8VzdrX275QZsx7Ql449oRCo
i3RoP51UFv1RLCFCrcNZqD1QhzisxhDJz8QilLPavcAmYHhKOozV+NQF+p/+bFrl
5UZlV5/Xfnrd7E6cQFjU6OjyvS5KVmHUzHcMYTxcrwcVXZIPwOY6O17Vh6NO6D12
coM+MYJPcJhS75RQEO5AtwpUin5n+8GB00/Ro1XzQJlOqW+YF3lzyWIV5EpxbKcl
rQBQaTHYSg8e5IiRwP7CuQWQ8o6UI6VqHDLjleRquJgqwQlePI+0+N4STqC5NyP8
adNl8J3ixs2bJNHdsaWel5J6C0PEnlquwEIvuu/XFkmo2oRvNZBCNzNSOeb0xc2x
n+faRDH7wh6HzDoFhZB/EY8j7rHrYrHt0MTdD+ZcMGrVzbsgmmdZrfukz4+/VgEE
fIynyJsXSP0Wm1GCu6FM7G93uDdFHB6NZUaQX5NJvby5tP+WxIs+Iye6eYnuCfP0
TB6lbisssceLh4T8H6rq1JqQr3jeCb8XamSAJn+PPiaNl6oTrSOtr0UN26vKbLGt
trLJk50RH+dt9RBDZwyusDlSF26K04wCtwkQs1PGMqy89Yg+bQyU3uYrCr/vA3V7
qGd5c9FMqC1tuMG5bvL1+RNRMW9LVJrIATzz8EYGgu33CEF0cjjzrKtSX2/h/hS0
4vjOVrUGOrDJwA5rgHH5fRl7gPDIg5DvrYfGPxpy+OcxHxsXv1gL/jayKsPhdXEk
fGGIDfTMwM9UFAK6rLGky4B3VXClUP3VTI0lj6ib5WZe3Vtyg3blaFnC8xdaTvum
Qioklj2KFwROfMtj0sl4HrtSCRhYDm7FjJeHvAZtYTKRMl5UPGZlwONedCt10dlU
UozZLgX2u70vPmanKkTpFGqkFmWto+WPULhUkbhoolw7g/Cv/VMhyo6ztwPsAjrJ
2pFTHYBqu8m/F4jVT57e0cOUegyhQGAKjlLh/iOc2xsNdgnS9YM5VEF3eAL5B1qw
g7sp1QEDKXL6nWOzIty0XzR99aITLLrzqOcJCYP5cniOEzd+4E+GkqYNCTlsUsaN
rx55rnRboYq5MCmZC1ovq/W2cTmKVYAn9ztOvfmncLC/ypKn2inaL9MlIwPX0ZpF
DALmnevtuzbOucUbBhn3k96ITBFTosEgeJikYRIS+jVJYVORiLroOkUbX9kH1kcf
XeFQdMVr/LgnugoL5c1CYHcUwpaKa5+ISDVn8DS8Yku26NylSc2dANWtmIFkrKbz
+vf76yINehYne72IRLV1neL0iJu5dwoApuyqVFs095aK8g5Z69yFTNlHIaCteg8E
k9yrlUQwMcuUFMMnzPQErol9m5NIGe9q+cLQ4wmWXquALfD7KqkyLQ3iJmRjA8Qv
6kNyu1dEQmu1Vk2JfF7fIMrnDgB3s3O1y5Q8uyCoIE3BlVAL8H2ShRVKI688SzY9
KZXFSCklVEUG6pp2UbK2i28caa/Cvu0vH/+F//oJKGZWOqMysL9u3OR4unX2/3Qa
iailwTVJzrN1khcQgtbPHLkhnti9SuE6oE6iravfR4OzN5mOtneLflDEjRq0iipz
JBN3iBStSGyQpmf26QQPsJcVNyOK7/Eb8LA3bvnFBLx7F0sNF6He3Je5FKF+TU3S
0yemWpjndcwzh1xs6MocVYjR4Og/KGamUTex4Q4qJnCD+iNw7XsadoFR8K1KIsbM
cb2SVc+INMRXKriga9p+MftZV93V6EfEMtmzlOeS9HH6BaYeABhU/BRWsWkBVI99
N61JM5t9gQEfP4SMlsvH7CABnInRMibe+NYJjCDCEyTad4L7qS6x9OC+zbuw1Ejm
Hs2rGnwbup1Lqo9PHKV7nkCeSnhktIR9LOazrz0o/qJwJ7PtxJoOL9E5xx0jTeZm
sGBkgEAc38MrDVxRvTGhhdBQJ5QB0ivzhyBf3XV6Tbz1D8RU9M4kHsvgxUzwAHB3
8UWJkf36LvmyzAkwT7n6v/YfFTxIkPAaa+UxrlkswZafgIGQ+cd70WwRypqg3zq9
edZf3SHgxit8WMJblldnF5+o/cpRv3fAy5QgxVBERjkGzd3kxnWa3e0kBJV1ajT3
paskX3GgbZpBZD5XZ44N2I73Q2XvWkPnBvlYDDMAsiVsfkeoFDU4RmWxdRMwaSaM
A7GgCWjOQOutsFgBGUws2yBfvPfumJM8sKnJmJBzRUu328xvFuxiofs3V7Sxus/4
0Q5tpL3pC9EXli2abIY1TRFyQZLk6ULGC4zF6U9zE4AixnfdDkyyjiPn+u2mu5x0
v/4DvWDSliq2KH6OXdtTB6nmOcnJZ2djhgTQDfI/ZlNzt1+ihgWProNOG6AUWfYP
WRRPI4xMZQjoflQwQimzUkSasZy+pjIshL88nxMf26H5xBWE0pnFo1UehOh4qV5C
xbV1ZOuLYNaND5VUk/EJQSsR6sUocKtb0ad/9ORnZbsBvNyT6iqb38TSt6C+tr0U
uW7O4X+jjFPgIOf1noOxWrnt6bH1y9XlFBqqKtFkedx/SKKBGMoXSrF5PuJ0AZ4n
cnrYoTyQxkPuuyQidWY/Px0KCkaIejWvQWKQJCtvnJVGAmScZ8ApTuGwtKIXiDnp
kkH5VSnLfkvapybG9orqYz0zZ8invbLam8V7zSmCLYuynAdJyzssaofGn5Te6g1D
BUSLIIlH53Pap+JN+o0NLlPnayt8/K77wFrFHDdpaup/AP/38hV9S9INIfJPCaQV
3EuAO3Fcvv6CL9nafwZNzm33EqRn8KbwFWG8C5w7476UxMpcgujfHf8VZyIhN8kp
PJBPPqlI7x17xwLumbXuvSALAjxmKWzuUnV1SEFRPQw51ltjZPbAlMU2bpXTKrcP
L6jLn4MRQMYOg7MI/D1cRNaHS93sgUemQHJ7EU0j82Orn03hnyrzrbsQqY1fXpQh
RVLuO0/eQdrtvt+7nwyF2XfYmIG4pGbvdbnDd4UgWZj8zVacRb24Tw7JmvJj1bjs
1joAKGCRUQ5rb1zp1ejCttWSiH+CY4ESXbC/lcVxGb2c3nJSqo5IpeDNGRj+oiEO
NKn1jEtS6GuJ8qN36h354l8feofyA6MfP7NlEK0B6WhMF20cd0l9e1r/TIfKvezI
O0wuuAP38gg+bvEzpgHSFI+AtwUnSrBhQa2Nt6HMmvG5kXzHsWNnyfLXp9ddmeGU
dEQalq0Xj3egMzGO0DWxXHT8cLTQ4sAYInAWyZUqeEpGn7LyYnJ0WiUl2mkQ+Z9+
acmtyc8FfgMYUvQgki7JIo5j8C0jprrspTKOfLAIUClGGSlXRUOSUia/e+EyrV0j
+xJ3daUNExNsjs9aWys1HLeBqF5YM9DnZxRno22IsRNumspYPIuKCGEb0xCmtYKg
8OycjxgwOnJlipd7E0nGxMv0HJgVHq4mC3QiIgUWhD9ET5KxLx9vZuR4JrmyFrV/
UMt+K22w5jrIpjQGLXCzYRxlCy8ms8+FmoUqi7xX4UEYgM+56PLkg+YPJ8XHOGKS
ZTKtYYBqFPj9TIRD3pNqSKbv7wP6ftZdi20x4eOcoaiZnZycpwx6YmIicVLi+GlN
aGTGuLok5wPQauSTM8wKAeoTJuM0LoF5qOI3E1KamVPmzOwcGGErsvEfR4jiTvd0
u0j6mstNb88VvVPIDwOxcpa/kYL4ymrd/gZu9ODpbXQ5EdOIkorASwJP7cpTsfls
U7zxds/LslDQBYnkIGbBjKMNrUO7+APVhMaLZMoEEy182FA2/wkfeC2H+v7e2U97
G7AQpHmJENjvp3LEt27/UELCDT7OH8xytsJXAVxnmJgXFcWDFcG7QmCPFv+OhOkH
GjasldKQVkFht+BTYOCxXpfp59hySRrXhT1OdaMUrwHgipmXebSTRHgzvJcC9mjZ
+P0Mt/SWf1OUSfM7/EQkqAm7JSHMwIRn9chMBqyQM37lB8dMnf9KrelxrvC64xKt
zAOhJP7ehGZq1VViDv39LqqiZ//TmV05zl+xIQbGs6LoPLDdrl2tnXUO80vzZvKx
srZn/weiLEHYxMlsCrIYoxwQYwp6qr3sqUtmr8wUWoRbDOU3VLXKAwhxFD1qwO9A
e+6xSXOLYh8Pf9hhRZveS7Nz7IRKrgj8LcpYRvMz3y8JFXK1iOENoOXLQ2b5Mo1d
iFkZTL27avlHhlOzccThG2Jz6BIkiayqrQ/hxQ01Bn1qHkoipU7EHlsKLS2xyfS+
v+wXvaebAPiDYSUQZ8o+8at2KiVO2oE0f9RiiXlg+fcSn9wTLGWT9HYFmRmF6Ky/
6CmXYrncw2WHgsr92ZULnKbsZgh/e5hsk6YkW5n8PHh2w8VGCXXgN7/g7xC03s9l
FPPq3uDxOJX4ikQcaX46jxeymaxbvkS5ZcNa+jDP0JvAhZa42Weu2mS7g5ebiNrh
313MlEYE9u7UusQDKLOxQkipb4nuiTZYoqR3P/03bkUldMPUTslvv9KgQXp8FztW
XOj6GiV35qQaPVYA5q/O+XvZ7m9USXnLpU6poXf1nXtkPXZzUpYH5HhbZvOYaLQZ
T9JZBhivDRyRK086bZ39vEVMWvAUADKfpTX4yZ8yRUDPfoGCKETNF2WfTqivpo3s
svXaX7aE870MxVj2WINxepjfBZF0fq9npFWmUdivBcBMoLzrDyCj6dlJqCyVXumq
R2RjujDFExSYG6DMqVDp3MY5a8jApja7x4hHD1fMyrlFPQyzkDz727vx2e63EJsy
K1W4RLuwgf0SQrWONj0oYZ+xk1Q+Qhl7vc3729qR3JWeet5+kNtKqUnDOtvtT24q
CfEkUnJBOlvc+UO7QmAlW7HIGrW/cBdPrQ+hJDWmdP0BnmxwjnNUIqJdllFl+xWb
QR61IV+bJM8R5HzOvxOTzHCG1yJXQD99WeQns66AlYEDnw9XnypbQiC6yzFDeQMx
RavQ9jp1UqjRsi6aMygglK+ad2ZWVnv4WMXGmDk4c5gvli+mbZyG5sWyofo83EGj
Peer9SJTWyKtrxDD/x23DQn2463FbXEUBW0B5LEQnSW4Oet6pfUTcESNBjO074bk
lAENdkPyVMXNfqdajBD3dUicOzGRuzN4aqiCQYa4IuBzmDkwBZOS2qNyTO7oteDw
DR3DoiM/OeQkffmsNNK5V/cA9FDNkNqaNirCpn/1oiNzmwCQDvQ1ps0bZbDMn5lw
Q32YRG1GytaRO0bp7xpLbaswfcAgvlH7Y6A20+JvKmP2K9MkzCBgkYXuBhclXYE/
SLFrdLUuncwd28AXQCAgpHpvjoda5bDjLZozPWyUQz1OQiFFUYhjIZEdCn8eehvk
vvaVlQuVWzlKFWbW9nqnAsS3PgJZkQyyr1Utk1oMtLf2tYI44hQJIldhOK6JiXCj
WAns882uO/j31F0l1eyowjLT3B0j2Rd5V8NZLB4DuUzddkNtOWt4bcaag3xlLbof
4ang2REclH9sjLVzF34YTdLpyE+zhapDkdLqJDLsm//oH+cksGJ9zcngC8BiK5wK
aVzbfT+Z1SPvTZVUsOtz3z0k1LQ1Zejf2GazpC4e1qszRoiGngfzPseCLNTKXorm
sxcydNKJdIdBjJ+Ug5BLgXumhSef98zIU3HzA9RVO1GL+rCS87BYPvvVRSMWNviy
aJr4ehnmWUJpZvbriZGnbrK0fU1wZxAywKfbKCn238hs6Xm7FMVSEF68vW8hgeEh
+xxqMDMVFEr8tY4R39/8M9rbi7EVsR5ntumdD8jXTIMH+UhbdB9LpqUTNWr+67C7
uHK6K7E/WTPNuXRC0qSmAI6fVkBK0FvjEp7P8MTNnJApr15S6xOqw3oZ2ShHVIcM
hwOiPZY0QCYD4NcEh1GMV56aYN+M1ZDWC70J90mqybpiqmTj0ZKKUlnqcyD7zflq
PnsnoqICfDP6Ma50kdCnb/dM4UWzAMSPDbrvP/2afcoedVQXVvtPbPbv5gxsVb/4
1yzqmhflcHiquAQXXoMhXG7MtamNp9MefVde5ycnkM6S6RnUqBEdNqAH8YmDPik4
IuzlofzxwSewQaBtvBiy1MlDNS7miY4reml9ZLiPynNKzYqSszkxrEwZBrBsCzGP
5Tbsgs4Ggc0P6ghi1I5Y8XFQg7sjk0ixaKP/XYxKVsBNh5oVW7J4aNNSugcqbFEp
PoODVWgIqbi5W0ppvwl7DQLEQ8sU7dRBdjL2Ye4Nm6xmesNOYcGMxPjscqrk7Azc
WCSrgfL6yWyzUVfb0pRozTv3MeZSWXiaLJYfeKKv5Q0oNMiwgmhPtYrPekZGCLVS
LdLmx6tVuBTxgWffO3aTWRXJ5BUgA5wShsQpbwfUd5lK7WmVgkZZtCjmo7ordGh1
XafShDurUXSMV8kCIjazqoHTFy0deaWYp4IR7lq1o7dlRFgGXmvuLRgD3ME64OrG
jHvSo5RtS6M+CHwDDDbOowY0Pdvt/teGQdm6WMHjknDogJmLKxTBJ4cMYBWoBH1f
8OBdbYV5L/FL/RjdsRcXjcDfwMVZ3db4cTr0aAJXDk3zESSsLc7XgAgxcyvsLqwZ
+SmTcGEtpVA6tHMcD6YDNJYd9wxG3nDpSBgLWxV3R15jQj76b1Rv3k01aoAkztoR
C0L7Zd/0gjSHIhvZgL/msxPXLdWtmPZKf/VVUm8aNZE89whLeQRnrvXrGIPL3K5x
xWyjDjfnrRgPmM9DUgJcsYMAgRIamEfWV1z1xaOQof6e/uh5xmgPzSOrgZ/iAric
irDM6eRwKAKuLo4sYSlrl7vVqoWD6r9WInfGP1UuVTYlmaWhmXk7jW6cb/iCSgli
WFiM4yCJVgfF9slbSGAO+0WuigwkEO0nZH7x50gavigMUeeHMygCq18OmsulfHEq
x86i9wa71NU7a5DGiqcNwvB+mX1Z9QoeNYDttHj7ZM5bwYY29BeHWyK+6ZidTxoy
PPy4t2/6q2ypYs7SC2DQkOy7ehq3yfzqemhAdEJ9KAH6U93aEC0pCaD4BKkWAH71
RjTQCzoj/jcQPhM6/2JMluVadhkPvR+Hkgsf1d6JdpToxo0KfTMvrkhvmyRmohDC
lMRwtJz1SHr1Y4h8M1VCrwpmXy1Ev3SAwAOu5Ea+Ih0x+vq7kpZX07i30lQo2ydn
CSRxXky7m6XkSLu8W0v8CZ8jksbvpG7WpujJHtgdzoZ6+ZUY/4MB15Vms0FfoyOf
519l2Fk2aHUiptEB7qBu5upqvddafEtIRhEp+nZvzsyAXIwXv3Fn3nBwN8ZBtab+
vQonDpur3KNng3+4LH4cuLxrkXDLaBPWnay9n7Si/aTH2752GZ4/kKSaMa28CWKW
NxJcixTs7eJ6ZkFAil8bl7YB5ZXxPq0PczZ8rBpsmxxdpxIKqVi2TSwKzlOtTy3+
jDdJ3YGi1LBpdcGy1Ak4HbQ25BjE2fW9G0cFgcsfG1/zi2wbD6Zhx1Uqk0PQpd7l
d2nS29HXQQxj43o7CUr3FTv6UPKPWtLRbO+qMcVpARNqkaLRgvvI9ysQvj4sUlHB
nhKkCP4yzg/apmiGKZqA05+v12hN631mkKstlMm+5/53wWl61Wj7JUYJ5Mpd2w4i
MWD2awsrVTvB8vTBSkGuvZbqV+4XLz71BWsqnyDxveiWbi95mUhS+JDpeaHsj/ou
flJqI0Mwwv/R/AwmFcJrPuwNQH1ZrFvYQyuXuz1iP66hrCTX3RhzEvEHjgDACUE0
E3IA0fDJAIOyyQu7TT5Se6E11deNX9m+thmUxySWK0BQ8nzvJyHaGyi9Czmk2Fjl
RcpMrVDwC11Jhmba9qxY2XkTuDwASaXAHQlkaDQwkRnnVWDS9PyXyh2z2xCXc/P2
w0swZ0r3nUscDrUVITp+YoQDfHPBNqvIt4ATGwoQeEj3pOGOsA+GILMtrIwKNsIl
XI4wD2wGa0Hbt2pIzRYPyCmkyjlFwbGF1Q8zJfsPpMTFmme5wFeqnExrWl3JjyPe
P0eAVnXeQqTW0lfZVzUNEONb9hlyr8YIgGMygWpX8BHcPTbuP1XPDDmCtq6UMTR6
fHlzzEjpeVf6XUn+VquR79o7pPbgT29MgdE9kF/+9Zs5bd7a+TcCwM3dtT+gIHNr
p6EbMq+soBstD5ff3lW693WBD12quuk2TPkXYps47vX9Mzw7tWfxMpAmJOjZXV3j
ECFU6jMnvfomif3x+V/Y9IGv2ugp9BcMzoudEx8/IKSj1heZjR4ZIFm4yyGzCveU
2ar9DYeWya++8GnjT4nSH+elJZx1/72jgRkkkxP3cBOxhrt37MP7a8Hl2m8GnX7B
eTphcmmxdDaMQml/dOCVAoC/TbQPiY/oDFhjwdKxhNnk3yj2rDh3MhP11DhsA4pE
lvZjF9pF6f6h3oBo/a61hIFAjQ6O4JAL30LLShHu8Af3k28vRU+zyP+bFU2RFP9G
teGaiA5/3v6IVAilDqzyyzkUoji6S4Gpzlw5adbA1fJk/z9XEaPvE0Dk9ltFfS9+
H4oTd91om/3Cn+ONDONIDSUt7x5OsTUGWyInwFf2B9jyUzKyoo6obOkd9r6dXDQC
9KkkLBusn/hHCYw9dKc27R+dIg+634WluW69kz3i0XYYcoPn1CSdz1fIahpNXXW9
moxjaqplgR2Ry4ZoKtaS0VDUpGMATkmJaw3xfXODfKpQ3rSrTTVyrrRcWPWgOwAW
CjHOf0UxhR+INSQQemuOCT7Vx9/beGu2eVrK5wwcwu1N1emDyZIhTi0RBsmpGu3R
ygpWJ9OpyJiD4kET0WUD9wJVRDearLyj7XCRJk4R08V0Dya0vvkkDacId9iS9HVj
hMliAqkWrhcdsp91WQW5grr5pwLJJTCYiyNjE6rm2MRd9VobviBoipJh77KPe4ze
DYRSCdSfsT29jVyqDhVwZQq4ulS5FSKS5Lm/u+lE0c+9xskTb1Qx5l0GYQFwwOQU
WSUr4ArPj9JVrmztipjZPl2B6fwZpIVog/ZiMi0dBP6PD+zZjawJv0xeUzovHBoP
C7TvHCWVtcjK1IOyt2ImxlKhU6n04zBdgRNs5Gd/Pn3+Ldfoi4I/a7vU4pqg7sY+
tg176J7deDi5Ep9Mz4IvA8w9C3w9LA1by/QztLjTA2xHJDg9lNLAabh1z7X397uk
1FTpV1KJVX721u4sISQX6MSYzrw1CEfkgoXiA2QeNm2RUGxBHybsAF0PVbZXqQgX
Hu4FPoYfdi9C+yVD2BLEWcilZaWk6jhTTsneCOG4/bFt+rvWVO/HhTn709HAsMin
grJoPz6Q+6u/p7bAi8yIF4tkEQpDbtFLhzCtFWtwRxBIWGFjKViq3UX73KHCFOie
w0exk3ff58016dS7Ggw6UkhGRQNylVAyDeIo6uGtX1HTF2JT0d445+xmMAPH1SIa
iyF7HAQmixp2+RO599NF7PZExostIsWLhDGyy3hco9YRCjjRWJidQD1ZU2r3z1A4
v+c7J9/i5sDtYprD3b1TOqgS8pIlXCZE2grrqNvAvioyVblKhVXOKuU/MO7QBoNz
AxNCAo49X2w534kEk+JUeKMzEevEe31qGoTguJ+iK2CQv4XxF/F6uEvRD16V19kp
BH2xSo2W1R4bOknKSVhWtVpIrczbqxgVjoBwahZg/7dr0crJD+sOa5h7RrfCSKef
PE1mmQMG6SH3/Em9z/IxtXmInCZh7/WGh52fjFhbl6aGVhM+9afySwiUBezu/Bnz
eceZjjfhRWoQHCFxG24a6NNEL4TO83LyWMz08ADMlkhmoSNpfTIeDy+XjAnmrVHh
j4r0MJXB8KAlHtgBEmGjiOiqsnDTDIvzrh6vyENZjD8qW+FMwP1DSqUNZe9hoHrR
N0daeBt7W9KDsBDJIoDZNjrX4vbeE5ezle8lKT43LkmeYm/4ansKTA8M2jTPKI/P
O1s6KRSHra1OluUSpNczVCL86ciuHw0BWtJU83zj55uUlrCfDqFDj47g82TK+uIJ
wYMkN44ovi7/o0hHFXzckIISh1Lgw0pJVYQX5gsm4qDMn280EaNX5J5OWxFM4vHJ
7jbaJ10YVfLoe1tkoM+H3yGqrel/FNS5rEivERrkBJAhd63iGsBLNQCij8Xbd+Jt
pUIWReqCu4sp+qicbGkM1ikebhWxl1DsoWHsIAxpisDuB/3vaZMX9eGuL1cW4bf8
vaj7TyTHfhxYxMiL95uMqlj+z3job2FFr1ZnnE8qpoX6u4nlDaOoBt7FoDHVuAuq
azF4CvQWqW3wZJx+sa0pMLGqhMS6M34rujsEibKCH4ieYYS0r46/KZguPxJsecZH
tbs8cojWvoGkdWZGDoThuxSjW6JBwbCY89/jEwjmpRqW5h5YeBuI7kq6OjkukgL8
smXr0QGTx9exZmYrsF63HOWAsTS5zU1Vlptw+utNGZWV2DYvGpvBcgQKsLUF8Mgh
gm+OiQFn85dFASXsKWG5U+tWUE7w+11BXYYxhaIjWastulYo9JZh1z9dRZ51MuqG
OqOTWZoUl+YvXHISUusYkm+h0qcUR2qkMrDW87ID1U2SotGmrfvq2stwtiTCRGFw
a0r17ZB18BsACpmeiyd/ALPy9NyOr9efpO9JmpsZ1tkONY+dk33+psKBMGuUtxX2
bbBAila+d20JzFxWD9TAkpCp31qHap35+ZTQ8KHW6IzLdbUVwOx3hc8xe8H94ZDm
B79Pl/3Ey/+3d4/qonAanck5HlaXicJ7UTPV01dt24qficbYURUd29/WnO5UVddR
H012wqxslvKZ8XuZeKEIsk5Imn+JjJYHx8OKxPUIJ9PnzgwaHH8NH8IBaNvXPog9
alGcc6tve2S1hV8akCbf4jf4GlCCCaonBHRxRPl53cWOQjntn5G961/t9Ib0FHkx
KUtXtqOsS8FDpJ43YfhIwEw7nEL6zO9RD3PsVsjm4y9vkICfYt6TwSQZQXDmGfwo
DiFx/I1lyCJHEzZG4ciQr2v3R8foU1v/Qkhj9T+OTN7ndCxhoNQBp+nK7Nrhl9RQ
6v7TxJB6PaHusfUixD9L4mswDLEuinRoSI4WZrzrQSYwAaAKmLmwdaohB/hy+5bS
wU+bVMGb595EkNczc7Avm1gj2xoF3d0CqeOb5Bg680yPwSLVW88ouWqgFhcVLpro
HmNEj5SDgmZMouA/C4a1AdLSeDKic9w+vpvCnsqi1MoUDa/tFQAFsi3kg2sZonVZ
SKhOdB6jv9x18tmZY043mgn9uyPEw+C164+7QIyWz0SiEe426j8p16fr4IOjAk7Q
l81YgmzprdX6jIyw2KgQ19l7xD229otwSWBFwW6mR9zZZTyRAc2ecW0tYLHWfAuJ
uSNURULnGdMMLEzvmKIZAEMaAkcnnV+Gp4z1GRU+hGdyb1wEAqexyz9sdIqS1uTh
f30TK6I/w2zDXAZ65zrDkiJlp3kHomtID5RMY8/ueubs8GIrD+XwmPEov30yypLc
b243R8fLZyiI7EipSg6IuZe5KzYbDpXC1mWRBf6BynpRrK0IqyNFf9wfW6XvGuUe
/r3SR/MjyWeoRpJJd1yr69KmRkd4ivn8DHsO8U3IGuRR63ieBtdJSNRMl3zj1Xk0
leXKmDZeLjAA33gGVkzqrJdfSaIomWnNsKKp//tlglPq59liMIuYY8w/IrMLZSuU
3UhI61NTdLKHI1D5ONVynGc8LzkcjzmlgC8MaYVlwVPBrQ18J3jZQuoNju82sr2T
86gwz3Nzurred+Jm829272z76DjvFsTDuyrE39+nFEYsJUw1eFw70hGQsIjet1b2
1C7ySYV8ubTLx0q3brxD05S1z8lboAl/x5MxXrF8NW6NLLqsfDbMD2QzlyRNs2ti
o2iGlF5KegGI5EvQSIEkfHSnGakTqGPUtGSMhQqA5/J9sANGODz9HovkYdcId7Fx
nvqvdVDPkF+5fYAwzgsgXACpcnzmmCPdi/DuV7+4nuqqlIvMFHWlZ5H2eIA50zCA
4xYWai3cYy9Zo8mhw/ARALeE9z1Iu1w8IPv0iEPqZ2aFdRbNJJprjl+4HYfBxfbE
3RrFkX934iekw6ZZN2o25tpQf6Fi4YtNLGl7XgRViliT3c9bNyGVb3Cy4UGXTySB
FQs7YyLxegHTEX7STB9qW5Foml6/5ckiELJvEzQ2Yd/n0DrtDAIEjqA0hNNkF7Yw
IhwyCNwrLncu8erJ28FeH9MEZRbdfHubExyGxNyUmDJ3c8pY3H0WASiyIjN6fA1A
SXMnDK44aKI4ePWOOpVGPEcgIQStFcTMqGSpNn77HQptXXqvaSPOLJbGmztHsqrm
1A1dYecLi+wqRN+CWITIjR8LSwLgL2iEWpjY75Z0PeMWtxrDcidnRml785eAvveN
mRJmTI/I1pqNPUvli5HNgNwDg6unnHp9Kk43U0cTpYxQ+1B6Ac9wNcccV0176mtm
NRNdPZUAE0fKogtK9+DxXv+amuzX/reyzdc/LELnAcWFvg6sznmre7L0YaB1/2+L
oCPDQMjPVo+qXUda1iKEJXK6V8IQK8ojig4kLnTyV/HTbiZnQbOFtWcTR7mKT3xZ
v3gAhw9543bkCaQ6UkDoKvyfPOzHnIF7r+MmzAR7y3fkl+yayfdEpBm089vevOR/
z1gkPB2YGRkR8/PCoO9KtFdPqoz6c1ZZTxSrinAto+9uZRyWwPuNb9vEELIW/I5V
sMlwZpWDIKA9jKjoL4NN/AU9pPH9qj2bDRsiEaU51oQE3fJnu/cte/7BVpGF/+8W
9stBPslnNqANNBEJq+Sd07eBAe7wSZqUDu2H73P2WBxGBCA50osnfLQzZJdMDHVR
yTJLGCcNBGNqP8szoM7Gqq6HKWL4+GF8NUbLZKTA3WMtjNMn8To2hssOJq4x3oDZ
ep+XMBqegmM/n/5TYPcXTO0Ut5Smw9MHJ7NCeCnXElKE9GvxW4ltk3J7PqbdkVQo
7AgkBKyR3V1oDKCfBgxmVbQ8u4h00X9HMfgD+7ivQ3jHgK41VaFVOEV1yNBPsSls
/+D9jiQdVbqlmYtEk4jmKXQcJtY0DJCg/zd02josYPARm5PiVWK5ZHUrU8I3SDcI
8hG0Mb0ULEKZvLqn+V6d795TEqTNfZTXdiSBsujcb1HzP7IsKXcPthZLd8WTBpIo
uI4Y09SGUcHQXX92dsQ0V9jcZkO3eDHnQXBb6a1CqGImzkJ2JvTHQFSi2iGxM4+r
5aAUS7Tje9JMyP9XC3ZW3LRtue9zezZ3UdXxlkDcy895FrUsJhQq2SUkH0q34gfC
G1FAybQfY9VQPV+0u4JuWId9lnSC8I+VgV9AOEkthwwxNPgtPghlmFJAvhHIv7Pm
iibszMX3qSIOvRW0yTKmpVkWuqZzkqIPYAPfZV2kASorGCWF3cS88afdzx+GP12X
51mpgVRrFZ/bXZJfGB/2zvJMWdXVxKLRLt18EG4ljYy81VJp5OlxFH1tGeb4svTz
7SEWXGiKcmDLabiKUy7dpyucf31LbzKHpHQvQx/VhRelXrtK8XgSj9pjSZxvGQ38
u8nLxYEBWyCX94XR8AGSM0kddXCB9lXXZkWLd/yzX7WPwhdET5iBPwph5qihbpY6
o/fOU7Rmbsku/8BoGlnfKbB/QKiWdJZB+TBUE4qHoCrAke2/cnXnFZLh6zKiY5sT
CZzpTTeaNvq4Nq3ZGDDR1CMK3noma5kBKV3EJI2Z+RSRIzNRZHNYbR9F+0xqnYhq
UD1pJ4vGV/ntplaCvbLHv9IMOggBe1hYX3hCvraCL+0DiKpAvnnZ2ss4iehgPgLq
3A1Id1MWRJySJmFcoJRfgqgLh0OngVdcyRcDHnG/MoKoSRiHH+l/bYu4OwbyXfhF
CTpOmTiLnqA+xPOtmhtxiHYWT2yK/1yMA8VvvEGsZlKCRIv6nStDhHD85AXLVfod
A2iOb39HZ+577lY6NCsJl36/Oadmg66HbtNT2a4DLBdkxDAp3PiuKDs0YhmDmTy2
VX6wh3+TMyLq6gJTugGphxNWaxB3d6YbKeGUzqud920ujjqa4VA06FlEryh5HdAm
ra6DbyL3tzuzI819FK/ux5CwHYbENy3bBtEEg0pi7eabSVanyMbSsj+kw2uzMMzC
/iF7CGA3+441LEmj2YWQbauEs0wBRxQg3Upi2hCVlVn1td7WUAZ+DAUgCxeJWGGa
ucqBSzd0y3u3g3mZqEU9QIt9k1+zc4KbPVlw9BZUscSbP0geiGmvCdh6A1wzo/4P
WRbDU1W2J1K+Z7lz3ecctkrsTvoilhTyQCZtbIV5WAKCuJGLELoMNolQQu1hYTnW
8MDFZGiEhVOKXbvKZpCqzWdQG79Ht44HkMscJjVc8FV0dRE6p6a8dShORwJ27a/h
xIG748C781TEKxHM2us919FCbjXZdCAkqc+Locip962yXbOL1VBCmMSKp/A5Wd8C
ctAq8m0BksRUBBejiOzrTOJ0wAoc9xowkhVSfsfnEUMBJ1HhTpxFLOogYCpSHUuk
m79tAT/UFlN+ZsCdpwwXW8nYeo8em9JhP+SnQagYtQv+nI1w/EPfks/Iu4ZGjIiA
Kf3PiHUJFiI00MroIGYJDmvpp7YjE8CA4hBa/tbwT3iqNwsPdbzjumuTrFmJ8AYe
n6Rj0RJnqpRg5pPsv7937NukrpmeHULGGyTa45zUrzTrIc8QXnZfTw7QzZdB2fdR
1iToyKqtACPXdTQngKV1OyRjenqrmkthu1zO2j9bg0Tof+Vcufzdey1nbnGImHE6
CclZ4DEp590/lwjqIf6xdQUbSKEOjo/r8UG+Z7QTZjl51tsOkZDm0e6L6KJESEVU
wwwg8dcnpD4AePArK4lfjg/NLe9MCSKVE5aCDfd0/DXkToOXVwRbF5iFl8yx9NPq
iwNVOyNoRoEly2uCkXo0F7oFu+IKK9j6KDrT2JT/bU+VhnvHIK53rA/trVCbvKUB
OBnyGaqdKRuCf1IgbaMYHevQ7SFej47E23OlJF6tanmCLV0JEaeX5qOp2kMhfhFZ
XbHljLUAXU8gt28p+H8JT7o5b1SvVoaHhGDJ7FW6uEr/69sWBIAlI+Yv1qh8qTYn
06bn0yo7g1lBRHiBY6oJr/9gxw03sKCQjYyhL/G/pq7rDIXYVyuY2lhE5U7BPVIi
5pjwiGY+aDEhv+oQdCl8SYi0rIseDz08RT4dDSKa8IgEgggGTzfjISuVGKBzyPxL
ZsqqoCKPExoo24DYlD9JPF3Fg4Vkdlg3IKG4lkXM0EuYJE7j4L6Il+GBYJwmgqb2
hW0D9+oNM6yX8QQQRQZBFeho0sCVMTUAtta/6Y3ZkjqCZ+D5x8gdhkrDiDy5D2uJ
a3EsdZQe0+DI8+Cz7aElmJHxn1AXnPGJXGkfcgeXHCFooIInQHSHG+ypBGMN4Ntq
898Hy9FZX15I8t6rzzuV6AiEbYO/bjKK3XFJiakbx99GqIxp86jkTq4p77iIUuD9
9RhArliy5uzjxAsywYWhiZRzF52kySN3Z1h0o0Zvnwg51KHgr+7cx/ed+TDgWMB0
Nb38/F71rMcl9znnbpHAHcWw6DXZjcvLmClnIxqc8nVMkzPN/BKIm9iyNUh8da5Z
zmKXPxlcPDfGt91nL0CtcsY4FydxgAipT4QRI4DTtCh11iGtLF6dIC5MzxtNZtqe
w1UbKbebYYFOpNI4ZbTPcchCBoxFUhIK431l+PvFCTqWhJ1EyiKh1kZgXyhtAV7u
doMZUO+Ov/1MZUhHUtSyNnbzBu6jvlpJyf2Lk74aXJPXuHtSNJvLM3VuNblbeoLN
tC+7BU9LxcKcLQbyHnRjI3L254oPHdZsDpXzzXTeHN5xFLiEpffFQKz+y+3PBSC5
x7/CjmIhLP+XJPSP7YaLsN51X99hl1JL3g68ZKGh6pQzfEzilV5c7owvQbpPJgv0
DIDLi5hYkDzdNVJTiZhgi7t6J7X8wB/o4WtmtPHs+rw28WQkktjaugKXPGDpZ8Vd
y/lER5EAGDqHF6qGVaPTrK+JgHor3u9F/R8X/OU9H7RUJMD+qiZSjk37jxQM1U+k
iCG4stJX+PgQ/65FW3+4a3A9gezOTJVb3OWYahXnPav/eYGfCJj7/SdtgK1eRSiK
jPxZWRz7PnOEIrkELUpkPkHYEqqKtYCjci4ZqOI1WMxBud7WVFHsmkLfo5j8hSsP
RmL5UJBCAJcNp+lSmUhVx6b3HOkzbv5K9MTol4nVq34j9OhjkP3u+EI2S6JfMO3p
xxlbWOGNaPHUzDTZitTWS3ArUrrbF2SiMGiHgfag9OEZIKZxs7gF56/AzqgoCUZa
cw0+D92QrF+BeMlz3GpHXYtrfMulGQR/Fik+/iuJc5693JLJwGV6eF+F7rckyHQ4
X1+8ad7BGIlqbfTJtOhH2LTKMXbIPJKsLnj5opBOPYjkQkYAgDQbT1uIjal/Iz6N
tqgRCh4IvNlp6/tZm1/pv8FpSpx4iNNJ0Yj31/xtzzyhUPAOp250DrWY1QVj+1jL
pg9ucBVF1eOxgevvJbXAKxY31kEVWyhBZms+mKvQ5GmQiEDkGBFceiWzKSPFgOI+
eRnJJWGUoGTRj9O53S2KttYA6fMIugcjJI9bVGLZFNe+xp8YCNNzAWwjLQ5josmc
+wl1oY53xBy+txXfZmognQ8YJDAAIwDT0r071kSTXMHdYH9aQuPP+7A6Q2TwrvkQ
OaVdPefqbvGoManitP7UNJVSH8IQl9ecii9HdY7gRhXp9aI/bQkq/BHsEVzh69kd
IIYATyPXFeUldLDzvvh79usizANTwA0RC3/JXKaJpLQER+TezLTeRHPX04G6PAb6
6hNBEA5ogYM4VTb75FcaM4c8A3ZrPvJH5W9rt76lfQYrBZGwgNhgyy9Dzkoi922E
1INhNafjfF4tLMW5J7XYiw+9kzzJzLYwSuHlsvl5toOFu3GMkwfMBjIYzW6oamGK
pWri1pMCTtp8z/Htd/1iN1PBwWFihtDVqDS0tHZS3cnYdMBRoLRtT3us3y6+wlWD
ROZ3uR8qqqCVoprgC/C0wdTvJXhFyXlITzzTUczgtDDL0crnZXmKeIL87MiR2K1Y
8okCAUTRYS/cnYsY5Pv6R9FiIY8G12jcLDlG11zGAj1L+u9DAIeeZaRR+w/klWXg
HsqziRIk1QpndzLRr1TV1UCB+VyVSPEiNEYMiHrf01K/bPvEm8DdY4mCWR/h5H3O
6D3cPCc4rTvGjD6iXNHlvjTQRIFn/yW7dZQgNSdj76XtqPzVXswas8Bx470ATMIj
HkTwtxnSLTRDebEeUtNlEOVDMnEPy6onY9gCYWhNdCnyCYs3pgEoTxxaEosJRDxf
hjXfUrk9ee53hXeSXOzwTBSz+PRiTzQ2RCvJJXtY8wg7PJi0y2QLPDlTwenftBUg
e6snXezhqay9XZd2BUW1301RZ+dd8RFEXUFoEfOeVQNg9nnxT4IC1yUcev2xR8hf
ikgR0JBaZmkJ17MZGZBZvubD6z+TJ3QUPGGJHkde5azOtCRvigZtxHDCz62UHkr2
xCv0tDg03lA7HuhSngr+xSyf0LpquiYaRRsezCDgM7eqS6HGoi+64apSjFimAbGc
jUa784ViCcgZl7zDgz6ImWtCMO9kegx0fRmv+FiXhopmBkA1p5LzB8PdEcxXTwiC
GQLKIjO5SgSvlgsqw+KhVo9iRmmXFgwhoW8eM10oBfclWC8UJgE1CDiWBuQDG5dB
p/H9vJIpiIswv+9KDGu3P9qLtOSifCOeKTdPemcuNgBhAeHON20ThpMSov/CeoWb
1zFa8IM64ZJH88OEn/xWpTmiH32okjot0707Mq7T4E3NAH2gJ1egjq3Ez8md7Jnm
4ce9bsikJM+Qv3ebrNT/802VIsa5hz19hdSmtNIOdDPxT8WT+t4jac1YwaSmZrJR
/Qn1v8DG/e/qr2FFTZwxr+LtoL95+yJT9pCFLBHYeP43jQeMffkzkcFlGqWAFK/2
IxlarNMJmoyzxxaD28Wg4OwtD9oQ1dF+Q1pA+46LTemZD6lupUt0iwE60uwFtlUf
gJfxTz3RgEWAE2Q0Yjr6DK6VA0xeWkAkjzRRMEXR7cIzGRJCuK1jd9DdRAIl/Biq
OLlt/LkO1wLcWeYP9JeDkc0E1fGzn6/Od5HmyJe97VE3B5hBw9ygh36S6nkunkfN
ax4Nk7bc8U69//0f7ocmLf9itxXmsGKw+gCp4Z4l84SJa1jg02t+VBr2ys9FuKpY
31HGYSXx3LtT/pRR8Q0B6hM7NVZGlloY6W0IDdhHJXPS6GjD80O1CRVxek00UALa
TziEUwh50k1R4pfMPiPIfCZLdqUrQNEneU/JkGRP7EZHaEF2yTK8uIBlYz+UCa7U
SuSR0nMr76gQD/O6ZuQjOVSVvoA//Wt99zqphnIGAQlkVM+Y5WiDsdtXFGLqlnEu
O2X3R28AS9/FX38EzU5eJ3vosrYnF2RVYB3pBx1J8Q302Hpdeg8zMO1lUe44I6qH
E3Z79v2cWfIsbMRggKP0ujD0Pi/ycjA8KK+t2WCpF4076BPhC5Upej26sa/XdORf
Fvue8o5EFZSNUw/Pea9dQvQxRiU16Xw1mZRJqwpuCACcs5m+axdsESW0tm4D2RWe
GpWWbDcvZqSGqt9pjCeJRwOY+RfHPwISnc4NDO7mKMpU3/MZoxD1+4roXvDlNpDd
pF7LcJdpBYe2NlGwb+PlN+PPv7raqMk69w3/zyK2DFiZwESxdQDo3zG3Pm1yh+jd
Kh9mRV/qT6boElXS1ZNt4RCbVAZ+q7RwzQSrKaL/AkhoUZwIp4S8INKUD7xSUNvA
RwEWJwQ7JkYfWSHcdyAMH2NozSKMRJ9v+JMI4hC5RRk1G1b3LzFBs44Pjlqpods+
SVhOn1ZFWXlMj3IEYNDx7w1KkB+QTkViS0E3mXS+qhYqngsN5AbFfPLYMXgCfzxQ
BXO5UK5VzTfWLY6bjmBdw6A3YN2dUkXVQDu1tIJZpRpKGz94E1xP7wS+nISi8Z39
7cV2TFz/IP16wkOpbuHwH3IZXf7Q/LHjhP9WZrhR08M4i6ozoCQYILGpOx8WfyrX
BIikuYBBl7POPEaBPUbSgDHkPIKv/NaV1yPog/6/KQeBCl+sLMLtHPiWQsoVo51p
TH7vR+vJqayEiSsufJxfoMXbsMK0rFITju4+spKwXnP8CKWz2wKAwko9nfVDi63D
qnAGqQ3e2H57sQfgY3c6Hx+0fS6N0+r4IsQJonHkO2/EhpQLA/VUlpKZzFbzU2Rq
RW5/2FxsV3Qd5gYW07BBNU58Ma4vd9b0H+Qq88V8mljF8Ze4TaJdhwJufC5RdAMF
kKReYapm2wA0D8zlC/ra++Eysanj90Mdx+l5zrkeY+nnjsfiDasoDb6+dKVmqL3S
OoBer0XWBlPzscMjMD+QhVEl3Yl5HVL+kaOOAydX82RdUoHdo8LiwpNJVAQ6j0dt
5EcxZulZxl6el1WuR4ocPSVjsercG62zb2woerHqlDp0b4nyazQc9wQerwjcX0RK
bSACo8b+6Xtk87wZwSdUcjxSArfJngF5q9tqK5JQIMryZcORQa4rpcLrsdBGCplv
k8Jg8TK2UhyWksbHJay1AgQlsSvk6t4Gz/4XxrhmT/Bp27ws1bZQphXSUp+KRno1
BjTBtOUKTm6raTOVfALqqVycurkNqxzTEkgnB3gAABqqy7iNgZC2ecrMn4Xf0QE5
oCK9+OYfQb5TtAP4YnEKRJpOz3BZ0a/jCfsfpBsxs6Rt/JjB0Y5/niMtSSD0cOw9
GDyu82CCYpMS6rX+pOwCRKAOQSvbaR858s2WVpVUkbXR3SeAUzvcoqcbsZf6fSeh
DVuTFOENxtz0QPYW0iLDFlZcLXXK/RvRNcdaL5Q9v8UaVr/BiL2ciCZvdKxClbs7
KELjb/67wIc62nd2KC44i0hV/lrMhX4PFSb4riyNEXk4j5aoYRFKZ2p3aLYWDojz
KXpEMuw/V3sS8p257dv4cnb84ah2OyP4usHR4UP341vccDT6wruRq/geo8ia9J3K
6kgMflqnMCCVLChcmm13U64HaA1IOGL2jDPq27zeeh8an46iYTzRHmLNAVllzLUZ
DUE9jIVa0mgonJmIjbrFPXMuhDc+EnDQEQeTJ6qAIKPKkUJolT5D2LqrVNVLeV43
CZET2XZTJd2yUbnnkIk7GCgXx2/7PcTznjWrOTur/DaPRoT+v8owiyfp1tW6VkAv
mLX+uhJ9hhF82fj+dESZROaPru/1E/Z/x2CY8weGt+QdDRmf4Of1y2Cs8MzwmSFp
PC+aY/v9js6byrlexWIKaj0TdBkWRyE35IW0Mh0Wxvv++vfU5T1Fx4CBiS5Dd/IZ
5NX4OMrU/nEguhli0OTU3EdUIFceH5/LX3fZb1Tu6VO5pLAAhGFQA+6zOVZliWAD
3nXPaBTzaHT7oyZ+nfCO8MkByr03IwNXdRBiRA9cUrjsCL+1F2MgiE1IqpFQwBPj
KiSzRkAZEHJSFWI9VT3FOw9DH+G27CBS3WbydxE+SrgSneXWL+sSL00TkgsmPDYc
t/uo2T6fhm7DxIWUly5jB2nPbaaNnhd++1EBi+W6JoQnO2/p9y2wE8kXXGphGItU
Asm28ZqqXA/VFOTqU3RnU+2+OeUCnUKFmavRB8YmqCoaRrgdev899L27H0fjCK8+
TCmpOl4enzOxlvglYNnvUYvTe5y8eiLAE35/iwimmk1pSyrV1d8BJlluKetuDRD1
16oRhVOZ1y2CWzuEbJUqUcc6yDyHxuz/vPSR0nHKAH6SmG3Cb2U4m08xoQD1icZ5
7h3L0ZAXCDCvtFuIueSMNfQEAO0usgsJ/MrRuHwsEVd21jtoNE6r9Rt/fshqK4Yi
kWaNIjZZAJXfODRBAOPaKc/bRJ2Z5MT/6VzVVbN8m4j6hDF5vsrf2TT4wSSaeOJw
7Ke316s82/qTx5mfvzTqZbkNtF/W0US8wk8pK/3dOMACVb0q8UbeT2zZs143o9u4
HF1AOy1D75SEiip9S3GE6Aq865X8ExfxnCguIne8pdI8T85H/ZdGZZjov86xZm70
rprJUJlzN2fXf1ndA84wWsINV1xiq8xfjV+zLoapOOCx0tuE20EWCAqJfqqrAMHy
cFTctfD7SyVjzDFsBQR4kuHtOjVKNE7+6GvdP/S70245hip3QobP+xKJRwDjzxxS
IMONa8kY08DygUqeYbtPoUCRmghAdvVoEpIkGTGH9Xtc4hlOYmJyzJYprOp2BSar
0bmcHmtxihFYrNysQO9hrWd+44rsx3e2qhp6QpL1UjF4I2CF+cRUsobXUkFWHDFe
L/vdcJJLC9ZkddYtrLBBgxEXOkBYupIsVZ1/nXOhOdFHxdiuhnBZljagJOEgQKcU
7wT6AsoAdfEWcxGae4bfg/lb3Hs1B+vFiTdGo5IJtsgL8U7h4SMU4kzp+FPbdwor
WncFlKyFK6zWlu70+AnnXWw+ML/gm99FNFrrJ6spVJzxs5ZzyFPOalYxuavIXVUv
nH8aVaH7B7/MHUlJnr7y2+FYmQvBRgsyelR+u4lzt8ew5rDTwGVxVB0P4C7XsB6K
qy1Oa/veO19R4WdS8NZ7caQ1KBqNIVrY1QBfKjUmuW6+rUTHq46LyIKMVcPgAMRk
fufOe918puuBkrvCkHp0iChG5aWxbb3YcZp3WwKv8ld2vaMu1iWDj+tn5VGPBS4x
q0jb6Supgv2HB6n+FznE9nx4S6nNa/ZAzG3JMBp/9PWxTZC4jQbDfwQIrnz+XCGt
y00YLlrDV0Am9R2L8DHzTrX8sT2GIBtHX/25VA5BvOvdv6fsupM54r4dQkHAk9aJ
WKCaFDjY/hwMLqLyH2/i+XJVSqyQpekbSnijScnfDDyBDWATnQogf4fX8VafkhfZ
uXshajX9Y+M5HOVXyb7o0IRbX0jdK5RGh3qUs30OcFWezG7u7vm8IwQ+/pPwA2W6
nTsYvaZ304OkRX7SGmumX9jDyB3TVoKctHnM0MSbYSRxrzNbYFKFL62MPnlMRmeY
Ch2+QTf5NFJuZ1D1ryrB0iB7SAoTtxDobz9z2sAlR+TuZtlGTDvDMaVgmKywVsVl
1+GLygx+FiIgSzfaQRPxMYKf3el+s6Iy0lY0wLAT7KPCIUEpfA+UDwEOAbWS3xzq
VfkUUzSdsUp83Cyf2OWth+JKR0LxU5p0a4UH40Hzg2or9cAVwjBkGIW/vnOr7sYK
+H6CHS9+5wnEm3BWoDMEoco4TXOrMv8fv1A0T8CUPOjSo9FYDDnBinWeb/WoXnny
fSWNkC3/dNZZKXvLelqPHbE865khoMNFY5SoBVh6LLqK230pmKLK4vSjrXFBvcbB
RK2pdRcL/uQjDoforkcEQbNudSYiyzliO3FEwRfOLi00lOiVeUmRub7MFGFi7SPY
5Nr50+0yPLQzaNYHS2wgCHR/4wdlOM4O8AYuP0nf7nNLMhOcp3yIhXWqzc67SswX
e4tcBTZMyJ+KrFsyf/dfBud8nbgjw68lp6iRQC3EqGQibNX7LGz13qFHYQCJNjo8
PIGaqHgPJ4pg2LP6ziZacbu3LEkKPlTYUuVVeqahwkExZLTGMf9fbFEpr14pwySx
GRiYgqol/PybnacFkkW2ejg36dyub+yBYqCSB1M7WBaspdpPxda5p7gclOiwG5Kl
HTMuoPt9u26s1DVftQ6iIfrZ2weSBgtWq21r0gsifDaGVrctUb1unBsT11HdiDmh
6+vCn+zrPmNQOt/dfN8SsqKCJ3BG1yK9wG1AJqvsS1XzCpwKUFCWTdWdGSuZz0wE
46DGxZCKeulCHRbAu4G4jOOQakAlNs2p59wwc81rekonj222cRqohG8J9Nk0Fjyp
Vb1iR+c8iRq1/69JYUCx9qzXgC/f2g4DLWRxMIqXbJblgK6FSdteWBW95lAr+YtJ
+cWxT6z8w7B54mnmo1xD+zYywDQVgvN9/mXG2XVBLmcS4Tepqa2RtgRrqz1/lA4O
P2yJ0lVuelNP/G4LJm6ZDWisffPhUClG47BWVFFIvdmLw4GqK0Epa2I4ndx7/92Z
PtzI9CXJsd0/nuAivlrMLVMQA8jUt0whAXbMRcm9eyPRq2bHKb+HBfHZn5N+cLi4
IYy5Z5M7sn/IluEHB25X7JOhg0RqnRqbNqfxUplbaSsZnCJ6LUzJdqCENFvcdWJ8
u3lKsTz6Ld4NdoAnMH26daFO6nWkxi2+lFOOw+TQf9YKkUqd3NeoR/ZsWVj40UdU
mTiWPufphKEVMJKsl/RUY0oSicGhdZKcG+eSrJw/rM5xJU+uWid2fexo2hV5ErgK
AMSs36Ifi5c5gjVyUXbqxBxCEbqGvABphM/XJYEu1sknyZD5YKEaEKyooYgO3ROq
KjQJmHENQ89KAOeyHcZLDTKDGNNFErmFn5ikRu2e3CMgYI5g3rS3HcimuITm8vvS
/UfVIqgbnJ2jrA+GcpvDNJlwk1mGPrN7X4bSj68bCnGBVYEdy1IoBMUM7psVy0F/
Q3zf1+HIOrhCgebhRkRhoSSznhIaPbt+AVTr7BsAOUWCSJR9Uo4ZePdiV1IxKU1P
q7ggo3qOxwI2VaFvuuleY87ftB0K7alnqQ4HUV6BzhLXMmnDS1rEIpvyIXvQy57x
ZvCCycBIA5k/SYnSphZK7MBozIHl73KxDA2ZzddcR4M2o6kqjQqYyVIws1IYraBP
inwT2d+TVNPYbMzLqGYJ7Bv6gEpjyq0UD+mWqEeB5SwCXHwg5W1wjpYXlBsJd3hx
LLrtMQKgnMe2Gtgjd0BAa9oXhdGLxB986tbolpbamWh9RyzlILFg9ngW+kv8czs/
YDtKCDgzzFqS68nksDRnvwJxXOoceS0whRxUAuTMcDojsQrqq64kG1rigIhCPg7s
AukAGR6Q+ogbkesJ0e+v0sZDmWCDkuKqz8pCP4QHvFeLAZwNyFv9u++i+l2D+AKA
7nMiuvPg5hMb47czL6IWzB23ggPP1FOYrPFR79Y5w5Mm6VXNzOyNSHl7TilN1pTB
XowdU7cdyYbpyf9DtEtXMgswDvBbCWX2hfiMVNZkimMpbzsUuPRAz1GmBalo1azY
QICVaIb/9GMQEyVBjcDu6/6HiiCbmUxdRmACafWYZUyl0jyxxNEoZ1xMIDevR7Vu
z+v6ye8lCZZpYQKqFByGiAMMhVTKs8wjll+6ldnbJ70C+VXkEvJIB1OaY5KnbkMQ
XL9JC0BJ/MyoEQW+V1eU9MPIIpjYm3BbtpW4EsU8CIxzo6SOKElGH9rcGtMfLiHZ
MlD0xun0uYGDZFSZImW+SUcKhmkM6gaTLUtRmjvo8HinnYnZz2Ki7xEqQe7g6Zdr
k7mr/b2RmM13ujRXRw5joYPaGpdoDKUIhS1ZyhL40UivcrlBZehQ/DLC4/dB+lvf
BVuaqoPzF+U9nM1V8z33eLt+YvKgdcNn6Mqekj9Mq6zOIO9Fj36oqVCMFVnY/9ua
ZqhPSGE88xbYNzkZMnWPp3KP0Oz6I6xOASaeWFDcwfqKytKb8Z6XRdhhJCZsV+io
usNDFqN40NIVazjKWNIWyCu7XXGQfGLdNIYNyEuUNyi1gJqA6S11ycSLMPcdURag
dvRZ7aqV3/Q+o17yqwRkeqyRv5zBP1IA/Zems6gziQCdMo0/ZMdcblNI0CiKeGJA
HqoB8mdTVdFXAdmS1Ec0y0UH5SQUCj+fC04gMz+FiNKqKNnSDkXnjQJP/xaBiC/C
xQvWeEpKB1f60HPLCvv8oL9TrRN2ry6YJHX5kL3bKrr6dMaKVjGefai3d7JTEbp0
UGuvNSRFUL9+TEcNprJ6fwS5BQuGf9Dm5XrnUtCwa7lMprMF3zc1RdYHu3sj9SWN
EzAMtMCBBi69quDOnDEe82ruhwUfqhScEGYcdeKQ9gD6SVLuRYO6ynF4ITqIxgO6
Ey7sW+LYPCcFBUu3vVhSUPSM/YPGYMrlaMNoxudowvGO5zHaOOxKThuN3yrbVWBY
G3dvxpJ13OpCsj2k0CV6lwMNpRBgd0Wm5ISWW3G7ZmMrER5zSC7FJKBM/vt29UsH
ly47E9h/jpmVdR1a4xkc30NMs1W0FYbc6WwKDsSQumiVse/B56jme9OQ1ohqOuei
wOheIMxZLbxTdzdiCM4/aibscun9FPVv7dsCYze/tQSSGB95GLl1pB0usCRAosQ6
Q9rIB3q24FXeK7c/3kLNL+51O23dIva/MfQWC09r/dsEV7Ywv6jv8546RjYZ3HAy
jwzDjlmSfrm+/b1siKn4rtbnN8Bdi3fjGkDPN8O7Y4kiDF2LfZHCVCznL+GbKUq0
5zANqf30CSdWoRSAd/CK4oZ+YLZtA5GqybaIeicCzxA97CGCnOwUxz9/fHL1qVW5
+9SRQBnSWJrsSQmLDdahO9j8CnCPpBDZ6Rm0ZTtRdeUNRmrMAwNtt9xvPs/m4trI
Wj8ZXkDlV6T2mRRsmOXE3YhZrqnnGzs1n+KIxzoOHuL+vTs0WmVSCS/bD5SIvn7J
F9pAFq213Ek4zFSIlSrYBgTYN7neaM9Bk7EBhxr/S/Cgr1yo9nf+S1Okw7xIrfsc
wlMY96X/PqDLb4Bnmzextz3bDdS+3IfhHP5h/nU+0iUxUk8yuhYmaKGRLbLWHcXY
2GVtZkNdmqm07JAPz9lLa4nGI79Sr6GOUekpBe4Zm1KMgTOBQqSBleWQNmd7YGQq
w7alaKPYorzJpAXtmKy7uicPqjNSeLIluCca4n5cUzJiR/Y5pDpk/4V/XS1i7qB5
mTIUKkklcVaB0BBwX7iSKx2RXxoBQmdSEtvzCDu7HIb/gn3zknwYUR3G6MY/m5o6
GkPNjMUM0P+OHHdzJ/w91MTx3ohojRiYywAdnPIiEeh33IRvtDVJUNThKulRx2xJ
xIvMT3PnK8U6svMBI6kEnyICyBopa6/qeqmFXHOjjUd5Rm40LKX9wGC70czbly4A
O/lCb5cN+YSUptRPr9WvnIRe0u/LeZ76E2b2cWNBV/TdZxjz5nJTKVI/ylkXTzEq
1zOxBF6pma4+q7vHYBzTYfpHPW5+Qn6Kki6/QTl3Xp4H1tR9eqlaB9neMlYcxw7N
3Ce+izkgFfZw8sDwPqhERzRMxNNzuv28lccOcsKKgODMLpew8s1JLmpwlIT/BJKd
5knyjRpkrHmdBlOeSwiZS3yYGeFh24o9SgL6Zc29Za0+lrtRqf+50yC8OT8OKK56
EtRNXqQGHaZ4M0Wujn0fdymjhHnwm1vWDe4F6jaUreKnGWAVs46l4Wn/YOOUt2yP
1Lv4ipd0EZRnhG6n0d7KZnehw6Adfjbfb2vg4E4LFD6R8uCxeP0X35I8brdY8SZf
QN82MGvZHWPlYu8UJfBcwoc5A1+GLApET9p0q2r0Ydrmrp+Q6obGEx5qt/chqSH9
R28pdyhBKOFaaf5TRoU+9FA0hxaUifiGlp++qJhe6q+WTfpAo6NN13phNeIBtY0v
QZ1ZlyMPrkgINANUoXsyoqjpXArjxSju0tE2Iw7F9ucspUo77AiJ9NRa7NPOLIW1
k57p/ijxqGpbUuc39+L2oSxxUnPMA0PjV5hh4ZORq7nNKb0D4m1EGI59Xp6OaRKa
PDAmVTB5eTe6IZZw+tICGK40W0pKBb7/HvuJ1TN5yrzihOPDAgW3KYmnkOb2fYaV
In8dQGcNqKW+ynQ6/moK6JpcBjU5aptBrq9ZFNqQB2Ms+75rnkUDt5sEKyTZNyk3
kXMsVU35n/y3LlPxHZqkMLAGO9QWOAWaAic87Ft/nwjBRhOrzI62e9KVuJxHkBBk
LcpaRmMYgFkl/iL2koH6AJMUpmWkteSbSdzy4BNn/TpeKnjESrLXsvrTZf7KZLUf
Hcajg9GADDXiDeRSUbJNzAsy1K0OUZBhj723xE5ASKR0T1fj9q3Al4z9O6wj71GL
LOcBvEmEZCBTY2QVmqWJAjYW5wO+ctNTvc+bhmiuLxoqYVflBAh+ddY+LFhuVIeA
yk4n+RCtr6RLGQvnbdS6Lph9fQDPNpEwgbxQPi0zdykGrrB97owYvjJzNYghCkGB
ZYIeAmvClIVZBoIsdfbIEo82QLn8i5cmxQ1KjmSRYFkl2lDXl+WpOR61oXZuKRiX
xxQBDgGT1DYHjxa/+dr8JsoDaMGF7JcTiNBGSzEheodHKIPmXw9owRP69ru8acWk
V6pMR35uzQsC+f63SO+qHcWa5OsOvEMXVge0NCBOTlAZS7ELEpZUXvPONtTKdqU1
7KihPO8+VBFxx16rD06p/HfKOFgAi1Nshrg6v831Ll4+mz0+taM3CxDbum66KGTG
iYHdMqknPqLAYWpfkvhDGXDldQVIQ3w+DKDZe7zWeDXa7E09Fj3AAO+0NgOSZQ/D
nje9gcDuAr5Op6i5TpvNRe7BdRo9LwGkm/qC1yRfy04e/ZTU5iZusIgMT6ie99zl
QvczwLa9yokvuxjUE+3Uw7xpGQj3CD5bsMPpMzmlysyFh8Uj6OIeUKuv3+xRHQF1
TPblAYdzrJx++mnPKXYW8di4IH5Mf4lnKZfWxVXbinNN5/f7+0UA6FmxWYnU+heV
O1I/0r+sUlK5utHqS8mv07B7PmQchdOx1rNfCqiiKcZxl1SXyfNZIVZqYUZFNTOW
Mmfw9HgeVP+W5QMwYhgpDERgZI5tunNpEQn0jh+9yq4AU0i51o8Zy5lpSDi8w26N
A+DPtDWn22PtcgLZIcYE2/266HEYkblmivmsAOlgruMdiUMnkxUN50kBRqArwVZ/
AMNEQStEQPKX/Jr9d2MGizyMcLcLNO4PoCkxXnSAjdsY7y8779Ut9i1HEi3HssLs
n9JfrvR9dfWqUq3zf+STScPu67MQBuvsoD6U1TR1DSV4xaAFCBy3stkK1e88StiT
u5vB8u7Hr2nnkFlZ0jdq698KepPnF1BlbO+xXwnmJOCIVMPMJ3e5U3m3VAZJd6Fx
Ips6pkqnVQ23SYRZPm3VVaLNBHs8i8viH1r3054XpqK3v6TwgspHN61zDzQw4wf0
OVpce3TZ7542+saO3rvymA9wf/jw+MNzJJxs+tInrkrDLy1yxwjXRtqxhZhedoGo
DAxvtOVLfyjU/2JpTKtkwHWuYZ+rV+oDBdGyfE8hUjEKDT03lr8+IrEO+MHQVZ1x
sj9BKns7ZKPjyT3LeLrsnYbr78byiNrGZ5L0yUbvdUPfRIiARa5sE4lbKoKBUXfs
fPP6KFt/adpv0DyWgu4oAF+QW0i3Xj1xoj8+8QHbvWEU4sSh9IeAOKLuV9yqXKxP
tJL+rLUSfbBZzdlBuhm5yD0joevpwHYAWpCPPV9kaCFewuTPJ3FNbbkTsY34yiR+
a0WmG4s6rMVjSUvYuDZ04t+Qy80Z1mGswIu9Tt0/EXRxEM2KnPlmsdWjsUQ1gR14
Vis2/HMaE5nFJJnYQJdR04XWqeF5r53e67XiSMXWaOdYBydaVV2xUR2ma/SyOteJ
37dHkwkZMjfLJto9eBU3UHR5mqTlw1ePumr4ZbKyXArLQq2E36D45qGs3o6Z7WAW
XHybDG/3ZjqdvGrPo4F6q17duS6u7ZqTeFeghd6nM+lX5hhUCEJhQ6HmF7Czc74v
TCHqNgsgcI9p+wx0XxFXIz/mxIKzS4vN1A4slWvRgDSFg7P/gfyxq/Prcu4Q1cFh
y0dPCUR+E/16Xpx7CgDhoDALbD/Xsmve850U2HJKVpm0aR5nqBf89HGZImz3b7Ko
F3Z96XeZMaJbjukSQnHVTG9JDSAZ9DMGQu5Acx2Wzy7EUTgOoXtbVQ7SfdyAZXf5
BnVFoDM3Vtkh5Lq6dYj1orYwQdG8jlN1qeEYL24tbFSCmy/tgOMqEcJLMV6HTINS
+XrkRoDUOBJSSlZrMLHRMRZ5GYgWHZNa+tOpkjiiUesJ9a12TsyEaqZ2TzfbP22B
Ef0OY1Wl0WwfgsKLw5zfbbn1x/SuxXB3bs+NcI4WP1S+h/ExXrP63OoizZB2sI2R
fiHIYm/Ds0vxl00mok/xXplmVtZqbqdsQI6o9NrHdfnFElnWfWSf5Wxw0WvlCLWe
q8orlOPzZ8n5jhYpp8dngmoyA5ujJuNsYWRyg7hHQMomF2N4Ylg7o72gLwBxEPAb
aOrmd391fXJdsdR09PQTQgMkPFaZv3Y426WEFASIIuYoKEpP9swJef1FR1RFxoIV
niDaGJWB+yy9g0ByBo9kL6PknbPBYg/GwgJOw+03xcGX0pzZLMw4BsAIiG3Zc2FU
O6J9+4lkjvl26Z6VQneoI6XKb9ZubXrQlBi2BdOQVmR6trcUxXfj+ndDarAEOUfd
8um5mX7KSZUAqe18WuUZx5JQoT7of2cI7IPtqGe2m8vxBzRGEmrnqpClC+quztr+
PxCKirpyVno7B3FPRZSxsfanxZ7XCZeuh+wqVwYSgUGBIb0xCsY7R9CQsTx4cmiP
Z1NdJtDb3CixhjVSoRsEtkUjmAjLgvXngupWbOlz3gbqMMHViPdfRpUORc7Cs7Z/
Cn42CdfnqRQkd44Mj7FK1rKdr/ufsJAqCUMATvfbHYFyXqGY1ISoLiWWzv4kCJIa
wRPRG4lHOS7jvDGasAVw4R/ZEQt+ny2xKSvOJQXY2Foul8FZD4kwtTToYEG515Rm
DVkCNFOtTDL7qkF1A+NYgxPvw3WP4oFI2wrrL9reoh0kavtpiao8G1lGNMgnm185
ru+FS76JDtUMREiRSklWcarsipGRNxpuyKAmzb8WtEmHYbfOQjo0iR3QIdvKFOYR
zdpuwduhmDDHyM8EXCkPcX8+XeVpqdTVwJWrSrNNHRb94QobJJoMJk3ohIV2VTB8
643v1J7P6HpsZN6NvRR8FickROE0pYtJ/QVw44mJhhXesAsp8CIjbwArLcRLYZaa
WFO70ahnNUoENVcHETPVkSPCl/WBkXoXJPUnDDH5fabYUJK0pL7rGuPX2h/oUz4j
44rEmWAyTi9qiu0By4rbGXNgze0Lq5PgGxgQV8Zq0jo27nkCscAnor7vlqiCcSA8
4YerQ/9ngxmb5E5VvA+pVc2lN6UbrPt1Szvuk/VB3yADGibmTfyd3+hAp8bNfa23
/esJTee6za41faxFCoNQu2yn/YOZilqHFFrjpwYzrjq4HPMbKEEOiPwb8361SnrI
uanO2Ok/yrj5TLTlWB6N8SKMicK5NlvvIqZjZsefnXjyfYh7qXAAouxoIWVaFHGz
pVZyrjc+XcFHtZwq/Lt4TTyi58kLaywxOHoVTkBsZ2Mh7kDwixzUpkY2ZELSr9yw
loHi1HQkr+LVgZFeX9aGv33g39Kvg3/ZYdwIV+7Ezob0DbBB7fuHzw+DUEm89Ly7
dOISgy4eDCSRELQb6+6C7/USLL509fVZ0hzGUGsTtBkn4tDac/qJfKDRIRvY733z
4E69FVFBePWMkreB3DWcMTSyhLXwTOBqVAV6l9jq/Ns=
`protect END_PROTECTED
