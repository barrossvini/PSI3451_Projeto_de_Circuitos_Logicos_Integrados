`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9x/0+a2X+lb2DWruAt8v3MZLrHUrbd1EiQK5zbeM9Gy1kKY61dq2mLdpDuNOqcXe
IlZLH2jOfVTHt+LylN/Hcx3oswFbCPyAXTA/GbKQld2qmI32kqDT2XLwLaKLRF5e
viuQzdcDLUcsml12iKxCIEIdyyunp8cqCa0rtN5U1z3m21M5O5kz2VpxXRMriA9o
y6C9T1K4P8FZcAZC495zO0r7ZXnzu4rcJ9r88cH0Hoi6AHwGyWkdxYhtyVA7I7if
tJ/IfekFHzCN5WFqp8ktFlrD1cK4XnPk5zr0WxZ/CPfRLdDlI9oT6AhOiWJdGsGn
uUWY+2Xd4cCvmCQQHbKSTorxeiY4zbW8eET5GrBtz4/w2TGfre/fkLAomsIZ24e5
CrXka8/tujTS2zwEVtZf+EzH1dwHZwDYzXB1lUSkHnrtz6609GWAVNAryGkwLqET
Oy9bcxjkoU82v43rT2U21a1iytl4jOA6Mtt3skYGujS/Y0nRk5pWR+xkMlipidZC
HkLzqt6+YiyyXxT7ydWYajL5gzXx/gC1HS22UlJQ4+jh5wKmCIQjPJLvnWB+gTAs
d+/hnw+/MQ2kT+fd0yycZSKV3DwFhlgsO3PkphhxV94B7XArimqWOU/wGiFXDuPh
HOHMMsMD3o5/io+4tXETXmuHJ1HDSH6geXNWqTPgUlndkehtGokrJnpDjkiDqJXj
qdhFmIbtxQSd4WXfyzVOzPhPgW3HFvpzqepHwAgnQCFqF3QBUGryusYJP+6O3fsF
YePeTwnJJzb0NYGm2PFPishsUXUlc6ncDwARFS/OUJMGZT/KuLONYlXRi3zScGl/
alUXpy0uOBcjQjMUrRN/niU80eJ8rQr81+bh+5dyT98aErxHKYw9WzdzEKk5fF48
k8iX3YhEOlIgAzBLxHapuK2P6Hhovv8KUfliPIZJwiZ+WFN+Y4lt0+KhdxRIVqIR
L+ZB7J+/CorqTOOJyPKrId6aNvna1cXV4XGjiLXU8VbW/fa3hDD1zL1ZNgpSW9q0
nwej1gOBr/QweT+xp1ha3TVr6ZaG4CNt76aozDHAzZsrwe8UZyeUHlHinvkb58cN
r21iYSWNPjtx0kEBfv9zvL8Q37kjJ8md2aAD4On02jFmi3bH24D54l/A3R7Zjg+9
rzcD8OIDuC+nLWf0FY24Fv+/TmTyaMPWw8f9jTVrTIUnXQgCBzKkO3J128WLo4GZ
2HT7UdkJTPy/d63aRaKU+tTSepWHhAtOOH3RL+HTFjTr8tLsXp6p0XIlnPhOgWF1
BzR2wTnyQNJM54V9fm5F0uJYkP3hwKUjnGYbJV7tXKwQzCvGAX6YWn9LMM6RnJFD
CtTTl9zFfPt60zK7HqiAp4GEBmDATev5tf8EGKOdMDyW5q33Mr3Syhl/Xz91h3eW
ZfqMWu9bTznpl1ad3beDL5iM7oDstavEdmMRANnz40bpyikKCd0cQIYjFFtFTTzo
Y1VmTjz2geBDGo9j13/thTPEiDEBJnmVzE+fflyp9v2qiI+gnqHV3tQsgVl5PkUN
21pTjW6uK8/VJgAT64OmUclZdcVYHDLGcC71j0X4/p4h/Z70/TPbK+JrW32Wdfsy
NVQ6SKvIL8VqzKNjiMPXgnYQvEP0pjF+M7Dafs0dB8dYqmjWQ2dBistsFbsdK8fa
LS+O8YjtaySFAXXrgrhRpFchxBKf2aa6K8CIQ7ARm0tXyS360HZuXephPfCpEN/3
CufIPk0ZdSCOcsIIejy17ejfxqiUqOodYIZITz22KLOanpCwPUfv6nDT6jN4ujrT
Fb0EC/LlubPgm0lSC/kLIfS0MtXEurBZbcLRsaSV5e4Eg7shHA29SN+sUICtp8Zx
euHgaRkJPpW3HjPisHIM7eN6XbYKbD5R1d/OlyPiDmioq0wqAZ28hP/K0RMlloMw
dlXYntxvFyrvzBt6FMohztcXBjalKPksyGfTgEGlOB6p+q0RNrkBeOIEEORUt7ly
SmVPGsplmGmnVDkbGiXz4LdiNb3vhxkFVNNLP4dVzuvSbSo9+ko+WbY3P7jXmcR9
ZChrYjfXDEcZfd1l3PLnfvPsTBU3uazQaNIT3mPs+gl8J5+2NWOin2fjNoT3DFPn
X+JBBd6Jx9yN2NBcPDGO2fbPQdSVqFniO+WovW4MTc9o/Y5Pik+o5edhzJSva9Wu
IRD2Q7ZcAX0LvEubW1n2pX0O7u2MUjyGiC3HhOd6j0LOaXHv7Z63fQXUURqFlpV2
+TE8VUefbgE6CtNulrLu+ajtvjZNm0sGlSqe4MJ6bWfnV/QsZgkCPEDlc7dJlk+r
/oYKq1xnZxhPmuDuMdm4JLanE+ukdzvdiFSCX/6jUAcYnysVGpCxlR2NyrvjDvLA
xFs5oN93PU2AotHXiHU92xtgGSjYUvc1tLtb3Hvw2ZJxJ6Pemxg0uWV0Z75ExyeQ
GZ9whUfKw8tz/el0zncEVBgYIRpFZ6u4Z11DC9vRSlf2T9cWbMT+jZ/9noEH+Ip3
SgVMdB5z8/8BZOw3j65Lm6rvRlOCsfYwuRCZ3ve/KsSIB1GVsk1WRQhDq1SxF3ja
vKr7KqgruoVHTFz18ojdXm5aWk5wtfeEQn4VRuV8iJGnz0lD0dZKE3ZcYAJ4fCX0
LGZ++PMqReQBE/1WOW/ZsuyKe0lnohU68bkgpNTZJVZNP8WnoZ+689Ds+YwLKvQu
wJ+LUT/pIe0nRH98W1kJGDhxP2TCy9poEnLtZDNCA3FbKRY0r6JpAavcIxtM7tvD
W34zMLc8qQdLFiYk3+lD/CLlqYOH5AGeqTLoLKkwrOjdifPQY2g52jSW7VZR8UM0
0wRwwNoopAElPkhQwhaj3yevFk30nvPASnjYwAHT8GUc4ZYVSfa1JbYWxzL+zr+n
fuhLbb7J3Rt3k8Mp9pWQUaLwDYXI/dqJJKz5gseRcbvZXHOU4UTAIe6al+pmoPNg
yL2l+X999A4uqG/znkVvbXmqHIEm0M0YELl4iqs8pPJTO7JYT0kwmTUKHaMCXq/j
1uO6ah/i9Id9ktEyLk3Gk9jqB/AedfUlw0sgeLfpgERHFaJIM6pvKMEuh2Jm0NKK
WIs6KmMPuRRBAD0Lznv8zyJu5X9N7I89k/Xy8tWIDtf+oHtoIbE2vSeiiLjahPF8
am7WyiTAzp8gw7KusO6XgQivI2e1VQqLgabbjZxWwZjS0XWMb7w8JJuCvfbB2VfX
I+uJoLoqGn4b1c/plgciqn4m0KJdWTMO9SMrD8yHrAHAsYogafYT6a+pdiz/jZWY
oc3c1HnsfwbHZVO8VlJZms+yODrzLN2CEA+E1FuXw6RfatrH4ZwmDc3Ud8ulttbq
ETednYkiG+poS9Kknyrxmhu7Kyk9xh+o+uMZXDz+P0h9h4vde3Ti/uJlCFKWNWqQ
QvRVRoA3l30jXJKt0TqonA6jYIAPogBlUWq1cg15nf6PYGBTsAMsMXWfiq9rC73W
+rxD3zwJRSM+/OjCFmbnsBt4buLwypkkG/e49WZnaN8krt10mJLcUBXmL8VHT/JB
7iNfdIHfow+AVAtHQobvpPrm8BV0UkIQEN6YIhzVEm0s6LGlA1/oEenvlP0Lg2XY
5SHDSy3GQNxc3n3U9IX8rCqj0N+fPyslDF2ElIiJJ+m0NJY8ebJgJyLAWDMe6EhF
vtg04n3Qdati0HFqCdcWLA5OUSjkuRP7xh+4yQIOdkRPZscG1LtT9dPB5t4QA1GL
7Nr/yqjYRglQGrhBCelRkcQF4YSvAYhzCTI3YhiDKy5y/F1aUWGtIcFih9mu7gxT
dDzDkb1Wwq29cEbtW7444EyYhh7Xs8XWMwRaa1cSn6ZOHLIsTTezTRbMMEQ6P6+C
foBXZB339cch9mel9V+bedpPHN1mWEdT690rylS6/AZfPgYK8KVZ00d4mNCUPpdC
hmOVDJ4e9OYbS0vzkoIvjvIvA1x0Jh2T5K6b9qgruucWjWa81mcriSHBY1N3TZ7z
g/WlE1dkUVTWMkFEtap5Ta3oVgN4FUmI4hJRshg5HkC5QporZMpb6yHOMBPIR2p2
YMfyAdnZoYCZrKPYAmYfwNXws/VV5KCjXR+ew3aVZ/txCKAQ4FtzmLXaOb+7CBpi
+mkEzhWSAtrnycZJVoG/H3L6sB8/AdHE++PhLfzcZtseisW3tX9es/NjqiwkKBNr
49d9vyi87EpZLAwWK7+xa0VVFUgPxDastkMvgs2NUcytvrIIZYjjFudME/JttAgy
3XRixpn3IOPFG+FfIYEr/MeBXlOapI/qSLaYwSIJMgyOSaDAA2JbZVTWy7d89Ygy
hdofMdiwH0gYWQLa3xa2zHCGdJpqGrOyeq9Oxh94taCuqZ+H5qgqB52SvyaY9fbW
zutrqTFtllGAMTc6xmVIy8tFPYVcw6jrCD4mw1X/QbOJyTfRdDCCl5O4eZrsami9
9oOVX2RMVY/pE+tA5CDn4N+CHgbNLgmtZzT/O38Hl9xXUeKnidFRyOTXvG6dHnk6
cSPv5pY4B8Y9vGLKehcBfF/BUTCgo62F3tswSfSrPEXy0t8EUprWtjhp1gpvwGm9
ROpYeR7XKHMmh42Zz8gMB/oCkIQJv4AiuOhb8Mrbiu+t0gfWkae2tGhl9vUuHmgU
k+vpkflg0mm74QZWDac92IZLuWPpZDnxzI+9YKKWY0MEh4eMfOAE3yAEK3VzWIsG
t0DHTpVOWRE6PycQqCD2WnKncfCBhEywmePF1IYLDTv2wd4ZUcuiodqh53VIqA1C
b64oxVvJIIlBEafHtxqgUCJ2uw9lRTI0xoFwAROCQNyeoT10aoXPyHu7Ri+gy1eJ
bFBjMG+fdXKiP823Y8ndUCXFZZt2z07xoSJ02cBfABOi+dSrHq0sEC4f7pAHe+7G
yiK5rWlZjZhznFUqtbp1Kvzdc5frmT5DZythek5qBBtyI5fl96B3X7S+ZvHCDxwo
CWqD2ZISJ8V6Qyx6YYcYjYtpu2b8NYS8yiHvjXG5JM4C/xQ/DEMwa1N2dBM2DLe+
khrK4v6yOp+EIP2lXOGQqrNcykDzu41Ju9mpPII2ti+bhyg6HZLkKkWw44GQ8Xms
p0XEXvuz62JV4SIfRNPy7EIIL8CoF9q7dXhYxpQGFsVao6OL6GnZVUu0MIgDGJh5
JpA2dcHkc/cpDXycq7Rj9IUIB2NaNLu5sYrVqFI8DyUU3sxOXTVNF2tOq68Wksnk
y6ikYqeE7DY4H+lOcQ6c0s/JTpHT7xZPSatJxLyLRJ/2jHUipbUNixwaJxhwVyPb
c5OriXjCsCrsubRvyhYsnrE7HxeqLfpja5YKG9xAd/5Ujx1pZvUxy0su1ps41hii
YEAANiXSeiQEgc7wbHtmKMfkjjrhKmBn8kBmE2RKpUWjiof3Hwd/FXBfl8Ou9aUy
kmXJ5ZrZJJxmfG3OmE1gKsL/GU/Vw1ND6RNkGSfYsyt4IiRBmTfOPK3bLb9fokXK
eRP7liUvrXZl/YEpOGqVl4liO2PZKo9HdZJL/R26mFlJ3Ee/lFyQX5yyeSEAwlYR
xvYjft/qbPuXCpiQJBTbcJ9vt9Rjre3xumuMBwILUXIehjfS+zy9BrLGOk73Zy/7
y/cRPqSSYgB2hOfYrmMmtqt8HbD7TIvFO6QJKB2gSf6PXV3zG+53uPK0/C7LQHhj
B/UhtvEFn1offg70lY9VsIGfQBAc0Z9FhixqHSNMeZThm5ioXQcrYcJ6GDaoAc+k
GhGUAVbLf4J8mJ0uSoKNLKFOGhm69iw0khOa88D9FwfrMTnnTNc2pcvVW4qNYreh
vpcemwtjmZeE7u9KdN0h9XRLWedDPtFOPJ9nsb4bZxHOpnBPjL88kXcfw59RUWa6
KgfWmnIPGPZY9ghiS0b4CZ5St8vve0qxlzANucT4IJTO0yZrbfnh4HQxQFtcO2jB
zWkt2f5PATagx+nk4/85pxXF1wxWdf9e5dB2w5j24if+2h32XGnXOzgxQ0m5fXMD
tEd2qzPaW3O0uy9vMu4KxA92uWsng6dq6a6VaOGaqUJNx6KFmksoZhKnus9Ebufy
LIdMmr3p5R5jaacqIR2LNMsMvwfXH+Cpka4UVbWSZG/mSJY0fh6Fa8k4iIoe1Nw/
uxMd9pb3GPDbfh4S+owOQmy/acr7JwZBGR7GqHrge4xuQ1wrLwHwcA2p/jM4VVN7
nI8H3riQJBe157Guemj+R0fCGYfYQ1aSjrMoaH75xnazKECtOiI7UOUS1vIXMtqz
fsr5IP1JLzqHPsYF1kujCiYflQwOUuZLl6st3dW9bnqJ3EymkXvzMoG2BAXUD+ag
OoPLiCSUJC4TMs74hbQhk5KYeEd5ZsVE9I/fkwRvVSktNT4Jx843uqmvBkDp3srZ
5PxZiZS8i24rq8Do9YdhQUId4JsdsvVmaHJc5mAPH4+jHd/jeIK1Q2rkgcplUWJ4
VChEDs5R85gPf+HJEzY+W//UnjPelmqZ0LVdhjV6eQveX2n5J4pXw0wZ7pmgrSPw
uMpIKS+WH9MKVnr4DpA8KrDq+PW55fB0kEEVTf22l86IsPPCkAUcieLkZyGdlw1i
LBSMu3TGDRrsJ763mtikkjUkzWDnmFffaIeJjcvnqyk9nyAPA5OA10pexdT44KL0
rajeeY5CIlROw47qv3RRcvxcD/z85eFMY8UwU4GMuVjavWg18BBNbvtFHVhQ+KCn
1rO7PDGoeTYIPhj82qfgrgXFb+DzU4sqJxFwX0oiZRZYCElF8JGoqFJ7zn4sXtig
tCXm733Ie4Rctuw9bMw5od/YFofptBoRt9lSeLAuIFKtGtq/NUXJ+ivrv2dlirvM
FqsoC1eYCl31YkdYvvYlRT8iuNeAjxoazrMlnRebjihdoi4xUxhKSz9oebbfH+8d
x2oD8yeeVGs/tQz14Rqn5ve2COgi24MV0kjk6OM3cir3BHWn1pvk/8V2rVPvB+J7
TUYJ9g/kMa2XdpKbmuH/1c52pyYxVR1T6zDnvLIMoc+P6+/XuvjaXp4y3fL2JNcG
sxm58SDfQqTgrwFRPSt/0Xr116cDYWvXn3pMj+4WiC/5BXon6QNfkJBaUPrt9Vun
8o5ouRWAejq8305Vs4wo+SZY+kJoGW2CazMrl76sQC5/LGKG+L2rVg1pQL+pt4MI
gRYjcwO/GIINgKZGetxrmYgxbhmD/WohKQp5keFBH85cthYFfn8TFpYvGV0FQIyE
zLQOw4rY0RXd2GgwQuH5ulzbr3oIHSILYKJiSoK+0k94ym5/CGSnk3bSsz94jY93
KFidXJmpIC9RKnOiEnRFdch2hT4i4+GIYFw7BeXXfRwoBQNRGMx3TAnwaDJCqoJ6
h1Ewl9m+oaNlItUD7Uyv1jyUtmhLWfXgTS17Xkbjeq62VyssKqK5zw01o0mUoAmS
AREF0595xpmGgmG771GKWNUrYAskGpyvO5yFdnaINtsrceVqZhbHkz5rBEs+a8eL
mAUVhZBXq9mGR/Jk675w67XYEWfT8MirXlbtc3mJC9hX4WoIhCbY/R6tkJ0silc6
6ChmmFLNjBml6Xgej6pyct+xsa/eSQmRGkEhz6Dx5lAYMvAgAQSXPlHvdWJz972G
UGCUr3Vjbl4Qu1LhXjiDxwlSrE+kwnHHeUQSGlVjti212fFxtWF8X15zRScHwcoF
LlhqQzYE8TeRrpK89qGEVMSZ1jACHBHEE8PLm466iNRQPQcxuCkdaoAApukAL3xH
N8XDBt+0SQLx02MpnHrOwm+GL+qSTsgNZ6gJMJ76QvUtr2roSRtF/qM1lKVy6tkm
N4G2t8ILnbUrHdVj6pAWtTTAXJpe0MAgnvquMO9+ykBIl7OsWtuHwlAqS8TTmVL5
nZ2geQ23Z1rwypuTt4DupchKa1NMU3rhwuYGeq49LRN08ZyoG+znJQykyx706/3B
RXg+q7TbyGMlYEGxAuW7b9Sqc479qCsyWkiG+YxRuFoH7bUuSQJLHfYR333GLlMR
hlNyQV/9TwOMqCUygKDbH6ebQ3rXfpjvoZuosfRUAskKuKs41j97z5EXpUpR0brg
A0Bwhr94WSV4ONbrzsCc6VI/6yjF8KordT8E5umgfDgw2VyvEi9JLudu1xeBJF1N
8qdK/FraV2BFJYyrKIv42EPHRW3Ixe1UR5IhfH6jueduD982a/cEWbkRhZNiJtin
86HN+8DJk41UAAfnB7KFoixlul6J/ljYTUQzHm2pKjp4d2JwjenvInulNlSkHIlE
V/3rGVNIk8sESe8uiC0XjVQiyhDfg9XihO786SoTL4hNBBK7ojXVbgc1nbG0JVIl
4B2qrpAANpHdUtEmBfDnPCMR9wqcMOyddesvy7cn5ZbC6hqBDKZlTzuYa3d2UMl5
leeiwugv20fSgfHQEdlyPhhNzJT6ZFmlOM3xz2dXJlw61FIop056r1PMlUUAW7DS
7yax4cPfciHjWM1QD0dRrhoC/3CZaYTeyJX+d6eoke4xuneIsNdf8g63/tOgnA/1
uwmqkQZ839jyLaGlArN5UvUELu0vEtknDXslIA/Yr7VpSXXZkl+F/qGi6MZTCDcn
Oyk548DkDWN6YFVss84eoauueYD/xyWJNZRw8n/p92RP+ViifmLgy94ey2TW1yxY
uJbKRr85AAtB8Qb0MJIK/TF3WV1TuqH1bMZq4Jfc7v/Sb+mimWH8HceqH7pEG2s8
jepmtXpRT23F0i2E5EcDC4UsY7+iaVrUcckB0wNNXhrzD4wczyocUedb94M6W+DW
BSqo+6w3/JjdhmBjHbaK2wQWUJVmnaK1JTC4kZiHzap2ixxnVE1penqmcepbqVBy
YO9W9MY2y+/vzdeL3WfoDy0OZBcSruNF/dcqhCzUQTh2Pcm2wtY0/bY1KSwlf8l/
xxhTRTWDwoSekHIsZ1puItAu45k4pZz5jotS2ywLzyaLig1ibzkl6fTyY7Lgtbmc
msSkB7eHC+VJs1m0qaYOsZEGyaE6PzQH1aku7H6ZoiNM5SMD/vLlcO1mkji640au
8v11SV42hckT0+ZjoJk8UQFbwF5J0YsPFulJj6R0eo9cNENffic6PF5K7kdA8bWy
YCONbeWmuNdRzWMa5+ip7YYBzkUnW6JITVDgYg9hcQSdQqn3ubL7CAdO82kP4TXQ
ErBBzwcLSgB1HjlfkooBboUxG3gKWMGIDvjCwFCCnqpveVdR96Ug6DYHKYLrAGHw
C0hAWwgNNo2hWwjFKiTV7pWFPCz2Kfrxueh81oo5TtAF3vwa4oCYg2q2MrplPJik
AJ0QMizPqqjY9X3Odu+TwX1NfjNmhlpniKzUhqUqwPqpm5IAy1qcXXCadZ78gB1Z
77r8lpKj48zpE9LzhBGS2Ktzb1tqAnjMOem1mkUB3jTnRh1nU/l/rhNNMdPypB5z
ds1iCbvzpNqL2hAP6ibZvw6fuqRUmB9eHnXyt/BA98byBIRQy4TS+ddtFSefPOGZ
My7XbDka/aN+1x3kWD83zRiuG7wBzsFbfQZXCi3K5kzzyAUpKGZnzS9WrCyMaJx5
dzx4SEaViEJEsDeL7bOhPHm2zr7m5CHBVkxCQEqTaPuIqzJCTF3slN4E7AMjNnJm
PoXpnZpR+wM9uedRND44bL16rFxfquHmYz7w6YIE4hTmWmhZRdWlcGK0yTyr/9g4
/w+TDURbC4qOxLiFL5INzcEDevLSWl5Q//bEZRA4KatCvCyWERU4fNT/G+g3fBde
IiDO9llX30BeutmN6NkyOg8DPdXgB8X7iQVS5DUppO63oDzsXq8kFlK2bBgFsPtr
Ly+L1VW3Y3FO1rHAKl5dWYgowa8qcMKeThpnYAFzgjQuuEyG8Adhvj03DaQucnxz
0dlTKNWMGKzNTv9xct42oCmUzPpvIpMG3eUYV704oHtED19SWwR+wyu0Gc8qcDTd
VwZwlv+OwBMvDkyLAQIuk2Td9dss+JM781zrg1tKwH7wrMKRQcFjAPr0Kx38PVnw
R8nq9klvrz1aurObdOoOJpJg3HUZ5h/WHbtGcss4O239hPW39DpUs8gDiN5rZP2m
2wFQSlnoeBAHSE/foQxq45Bm08Z6T56iJE+pHVs1m2fluGuV0Hm6hM2VOKmzLKch
Fkbad22OmVxUCMjFUw/ZTUIFCSyfWQ1N35QzdgcRhCp1MHp9K/6GXHMg7w/0BzAW
PIJM0vZQmdRfIYQstsh1j7sJgB9HlPxMDrkVlUDC7OzqHXnB2yvWrBOpBD4uEnma
L8K4VxL11STFZg/H8ilk0rd7510FfTP6IQ1ZWaGr3rZwxMVswGpGNVk5bkJKBM2Q
bZ5+3d5Ixuoa9chzW2yqA0T6rxkiNrSzw+Lq/gbagGVKOWiupx6C2e8TwPxNb0lw
dg5fkPqrS7HkRqKbsN0mSMdkFxycakx3+xZl6dOfOs3K0xlC8FH5/RCg59CfW8h6
uuI1HKUVJUTFZVyO2ShPAXpNPJFX43ZX1jciirFRt5dgZ5WxGECVm31FWtM14TDx
Ww/hS5MJg8XmxbALWZO9BKD8vpWE/t3PBsnhbWFrXaH62jFv6CJSlQZH9I1WFQ3R
T1cN1AFKkQEhrUqsVKXo+5qY2WiADTOAhhWMUJv7al3c/W+RZpott+xeqlCIekai
8AfqoOVMSBC5x9UZZXkwXq08oGpt017TIo8gG3KVwu9Lncw1FxcUoOnDLMKPkYRl
9j6+ptMPbTfjPxeoHiAD9hXVt2wEb36pHIqisBxEXpjXKhIea/4NkjqQNGeOe0N4
c3x3pPTscc768LC1OQ1VvaBgZ0SAFx88A4CQOSb4VS7VEIQQjg3PAlC+/GJ69yl6
a8c0KazyOMjuqrGLZsvL4HVFeeuyQQo6FFAyH8N3KvCRu0nJc474K4MynBBOzUJE
UWyBO1Hng3IwBhThj6jfhGop9jSIO4WIyu/dxduysFX8Sh2NSCGmqn67Fw2P5iNp
MMhwFoV8ZJ+ZZSSWKO2AYeY66Wjtbg5zJJOA/9erwH7zMVEmdHUt3eNFYYyPs/dR
3+FsP8IliCc24i57y7IIsN8o8WrPXyf02iLDnoodl/H2iGrEf/mJ1WphjCVqx/QV
nq0RA6MN05ZkTuIEJfPhHlN+WHFvlnpJ+pr5AJalh8XBFM1KSqYig7Kws+7T39PJ
14CWhlWlZCGmnJIpTgneO+SWgSGdjKnsZjV3DhHcVWxdql0yFNDhyJGT7qotZMVw
O+jZ0QThGH9vxizA9hrdP8MoqJvXiuw+ZBttkYwxjlrnaXSzagDiPA/hHWlrhfQw
mw4J3Wm/dDtGitWXXuCf4HXlU+cjrbD0ngHuPbTmETYuGoZ8mUz2xgY3TwKT1r+S
TgjAjo6uq7rEriU7LQdLODLLZ/G8q+ETB2lsWWzdzfp3VAKjvO+xU/xtF9kxkUmQ
qRGkctBnXdGDC8if+Tlo32eZirWi4ftTAy+bdkjvr3/7K1tVO5DkeUk14qPg+vFB
yzSsYXgkaNbe+FFnS0eEdh6hdqslc7Ig1lRXGm4Rm4JJBrnBYnnxI/++Hfiwz99y
BhlbjlW0/eZoG50rt0Q8L7fbzKCwMb6GdMGcEIXevtDp4Y0Mp3Z9TsMQxu3dznZK
b/gU4c617HtIvA8LkNmzWJRATxltaqGoSEw453I7z4WujbhqQtHYIVT9BX8/cDD1
/Gm1AWU25D1+2bQerju0lkPy33tla6HAkwPN7UN5Ld4mggt1u68GoiFVuOe+gGDC
9nQrEEapjJIur9Nv6eWNYR1/KPNb3NfJiDvxNtmqIJyV8oWpDPWTbq/tZD7QAUEZ
4v09mUQektnhLemuY8eZ/DTz86vMNinV2WcRhYbhLpojQnLTnvKBjcjNDFpPj8zW
LcK+RGXIgAV2xXry+cM4ohTIBOsnUn/ia1DP3xEBH8QmWWWAOeMfbwaG5NNu2Ei8
yn3NtNIL/ZmlaRjZ62+9MOX0E2dW3Y/AA+IrsCLgLfpjnBnqFZiAw3+mjlmM3XM9
JnppeI11EbFsYvEaf4EV7pVerDH2DbXC8d9yGKdyeWzSKBbKZSsbcHK1+5H6FPn9
z267YN7WlQyLNTcqxsuiKbfTNUSSTJt3mrR+akd3jBgG3YxMtEiPkqNhxq8nqGD7
Ca8rNJi6JN73CBEHrt+H4sACS5Hx3UTYFETVBP3ruBscU//zkD/GPbuSKJ3e6jHG
RLtjPNk2W9fhxxytTXI3rryyYjY2xy8wcMn3hhKzcT3AqRuSSJdQnHPN/WORYLoU
igfO7Iezt+MHcoxAIUec6jc1roLER0TGkTFOVHiAEj5hg14cHJEUPKYKKUo+eAup
U5uZFzoR54KRk+VGRqMM6kbhKy6FjbJxRgh9sYGqe/Ggc4b/CoiwW/zbecQHwIzd
N1CrePL4g5czYKYBAhaWm2BzILXncdjV6+2Ne3xRXLAXuxFH5lh1nZhWDxJ2IAzC
x2w2QDC5Eq6Ft8uAVFt30ZnEFyaT80jUukYUvPCQupQiJn+8z4SemSlebUBV6fLX
nSWkwIQ0JSG7O/hS4CGKTJy/ZbJVO3yvCKbyub9+C0hK2uxkEqHDXK/qGxEMRfip
LpL/icRRiG4cZxk5iQgSFpA4UoPmz6cE4i5+/QSEqaaGIXmGuHhcTLKLxEsWhjHM
kyt8Htriq5JXGcfisJF+Cw4uzuAtJW2OURC/L619o7HJVSc7fBGV3mBvh3XnOSgM
riJk8TeHZnRZp1VJTseNaUZAmsxJBxhl/weFK9OrRjZGFzJSchjfmEYkOO841YKK
USxSma4e4KmFB6XuMGE3zbvpsTPOcS3w+iXiCex8Z2qjYfJPmKit2VonTJRFdDp4
gl6LH6PaeBRp9Hxx5PFKhTGnwhaJYoavAm3QDFabidlzqu3KscanhBgvCmX0ABDq
87/sqzG1HUAqLPZEHCsMeuyNthPTyablV6/23zTtTsiknj4MZ/cVNASPEeZCHzX1
F2Ap2IHedJpE8u7qcqhyfVFzandYPzCGjKcG2xfs0T4ev20i70ct+cP8HLL9dNgQ
sJNykgew2USekx1/2R/dk7htFQnjpyUOR5mZbTSoZplOZxtoXbyGqs3mhzQ5puIH
4EOeLNoFto7suO0Y0F+RI+OJn7myFeXNiCYyR6Ljxs2hUBHSZJfu3aLcXZHlIGs+
+zJg8E47Wzf8jGkeKO1lpOblo4HwQbSJhLIpDwCklidF+fngde20tjsKobYeEA5m
H8RFM8B8tzZMCGKn494mrYKcAwXke9HlH37dh5nh6OC1XOb6HMtMKdeQ+OdiSBCa
rr6BhFSmFCX5rBAOhr3CAkhANYXgLYS8osS4Pa8BWaVBxYipxYx2CAu0pSTrt6KG
6mU7q39J7D1Ia/13NBc/fHc6SBof4ejNdR2pYWqdl5Q+NfNpUShdM17bHzuK3HJR
yS4yOWt54L7/+7arspGIYxd0KsuXL3nLUVHu0M0xocVxyIhnVBvax7kZAGoTswtZ
VHRIvNO85ovJlo9bsv8JjvBFKEFWIGUWfxNwLeRq+DReWB+OfdOxtJic8VO5dKPH
TMpxQl0qPoneVSiSMkNQKFgOwj1p6IIG3wNazwkn6y+uVLmXkiXmJgXcbSeXld7C
Ia/3uvhsYQzqBpW3sAYVZ+Zi9gAYeEpajRTZEI28b6hxG6xrMMLJ7xyeOYrvONhw
BF+GlmNZGMYVCH2zcFg5OoIBH74EwD4H4w8fZDXXor3Gjjq1WfgcJLCIwzwkNSrE
j28dwQKw7TnNEw58QaQWG3JG4Zs71JuyAxnle41UMamyAtdrG5nuFsAkstbUwdL1
8Y6M5VqZzHTlvRnTclDVXHJYTirkeh1m3MAeP3zv6O+r6hygoiosL1EhCKQRCRYa
s1Kb+EqD0Cp0pPR93pwAGus4cw4X71To+CZEfrmysq0P4ul44VFGUOnM8BDhIVsY
b7ZeHY9gnKAGUL05E2zAUgvuh/gaLd0slqu6SO7RpCaP88i6k+QLUbOZRpGVniiP
yzt4JpmMFCdTqwQajbi/CXfl4F5+ESco1czQ4lNvEShOCVX+TXTEEbfJIDsDaKNm
nIYshS7iNBgef+fbvefX+UYi/Yyj3PuMAOkqHDx9mAcVBerabOvmUz1k2y+12HSc
qbz/eztJgBYsJDA8VBRr8kKFEcUlr1WgR3LNBW4NwkEbjImi0s5VyI67ZW1aDFEl
+vzFpmezzIO4CPTJNyBhzA0bOiDWemMJr5/XqTyzg3E+1pG0muJAnuWew3jdus06
5Pm1Cv+Is2fTVuAbJ9tp9tv6pILPwpta8LBfBAHqd04zdYNY6BQ3r19Te97h/BvF
k8Gea9alZIPE7H8hJivKRAQsEO63M3+a99EhBbqsw2Y29GZ3LWdziFVwRW4I8C4W
j74X7oTISf2ivefIjg+vZj/f6QS+1AC/UAQ8z3EsO5Fda5URpcuMTue70uGk2Y0l
Ws5A3huWcGqjxn1XNfe0VZs12bX4pu/MDdsQ6LzVxms/uucZilbPYFtowOWGHrQn
KEOm+W5spnYFN1P/fMKdfrqFBLjN1LLh5kbxAJGYoAtr5zEHZ+E7aICigE4zjp6E
mmIrOsiK1gvS+dD7/nF53KMio48DXLYii/j43qbwnywzHThhhcXJ/dD9MGsTrZkq
HPyOs8VsDCdXRIh77mNVu3tJouuXC4TTIHhRzIL8CVZc+7Nr8RJ0uKGYInfIQvvf
4vMuObTWNYpcmYQZhn0C0V8uC42gtQkO8XzVbwz/DeclPR5QebBrR8VSHdQr76VP
Ge+RB7XqljBWgaQIsHy4Sp8vHtb3fbHjQyt6eGRXoG3yXTFt3mbkeIIqqBHAtgeT
IAQr+gWVGi9w38haCRfI/xohMEhFMHSp9doY+X/0BEoL6VeEd/4y60HkzVUoxCLU
DR3AuhFnzzpc1lnuZTKmjtcaGRMYqp93TV8FgBughb1LlR8XZXNMH++k+Yb7W4Da
xYGOXxH2KmxJLrcRBaCTDZRTvWl9qBlH/dLPdgwirXMOBVCEnPXnc+jKsDDmjmxc
Hngl9e7Y+hIJFzU/SZ9TkuUkkNKe72tAHTP5sQC4zUkZN3G89hzrG22hXOjnTN39
PCasp8EiNh6RcQPkTv80Iue8lAGjxngDX++FHeJbRV9QNGw5o8CQidfSNRaHhg/A
X1BVS0loeBzJoiwQBMszNbg2D6i5VQOU0Dtqf70hbEGIqnGlfN219DxZXcMjGAFf
pJaUG1zZuWkd8dc1/lmjEzR9wBTKG2pjMwcN2yNVOM0H+/G1aFdzQM+ppL1gUT5v
4APJ/O8Ci5O+nbCDwdVqgwJxnGu/E96HVpPFMGOlM295ScBnimxcAjkzgiZ+22bt
pBFHJJqQ4NgPKpXJoTiSx9FtZOrnA1CeULC1AqfoVY8BwQ7dZF/zjZ2sTRzlmcuw
arLN6nEMTNdqDrTpRV1opBnjTbkWF2ZjpJNkaaC0PlOhrGANQ6ptg/cmGvNJcQC+
6k8Nic2+9KUrHhFx7V2jLKhjdN6x0alMFdm0GsR4abIgA8GMAIT1PCMxo+ah/i2c
FNM8DhD/A9JIJPuBfRlhr+q/PMlxBRnHRet8wxl/O81LgvzJfEcWgLJC6uVvwuKA
nin5ej390KmgvAVl4+hOej97u2mAZY9DVaVZltzTauOuzEHUZOwGvBhmTEY6IuHs
IZonk2vFw190usvJv37XxBk2/cxPbp2TR8gM1jpXb5Savr+V/1k+DmCml+nDAPaP
j6ijtN8aH2+27ks4gUG6iyaPwg52mnXSZ13okdl6CId7d0MmmV8+sf6qanIGPa0i
LGOaG2PyeooIag9wWTZYoCFDC/zvBYE+aWZ/hIQ2VvR+vBnHezNyL8A4TJB8AcwJ
4QqWyQR0nJJf/HCNGVe0Td1NofbVR1dcLYYBpBw/Uti3kRe7Ifx3D9xW4ucG3aka
eiivZc2oSjHgvTkWHPIljJmbAYb9mlZ6dlilmlkIUhPBWDK1Ae2uWiWdJELMxQ3e
Ezzdv+Sut+uvjAxs/6NG/F3nEfcVGMmmBSEBvijCs9hNTUxzu1T/QxoQixes/MWE
F8h+PbZhd2L1HfprE1ikwTi2/l6APF+Y0YQH5rSbIObzHRLa6hDM9yRFLsRvzoXC
JRE4x5rT2CR0ctIhOTFCMAkLWHsGEJBY1+LAwhBRqjB+9tfWb3YTfvuYKKReRR2Q
0byyFrR/ccvRXd5qXTw53dxCQju4r8swIfBz6IZ22iRE6CKgin05c+UbzcA0ViKw
z1qudfZBhMO60FDaFxK3VTDy76ooRqhjDPc2JnaPqWEOEH1wF0oPV1gw7vMiKHq8
MsYVzkhgiwekR2EIX1QK5yAzzURA3RczHgYzJ1ZQm3QqziRxbjUhQI8A0E0fX+Dj
N00sj6qtPFOT59SW9LfSoP5vRiayR5I10DlNB76VVH8zltA2wvJSOGHJd1OrakTU
Miaohgo2xvTm63Xp6MhY1iMWs4ZRkED+a9qEeanlvvio5d+xJ/R0Un1ifXFI1t5d
5PvnrRXwoHbTw+t/gyobAwuz+qb9md1+pL36p7J3F6mgE3x2Ufq01sWK705We/fs
9zAzY93MEp9kUNX+0IJJkaeOX7w+NsPxe4LxG3ILJB2iwTLvkUizPXRd1e1uP81b
DNNUToUX52DIBOKkuiSMgYyPe0x7qivc0Ns6H0CEztfinghWBX9UlmwPeH2a79o/
/hkuAzOR2e7i1k5TJCsi9m7tdKWPYoqe2Rg0m2mHh9HYHRkH6rXT5zHd5CxyKcwp
0D9b497Y8D2qoD9EJHuxWr14AxIexHoOy4mISKmbZFPNRUVrTHehLtrUx+8nKhRB
d+ukMDZM8l+y3LBHen/z14kwnPoZHVAfO2cZDpGZllh9WuWrvXJLsGz+gBJX+cpY
s2IkxmSCxsv/9vy0YtYCPKUu7sJ2AIhvMTjBCid0liq83HdUlG5rbLqTP16jjhBf
GHMbw/gehrnJpXWc0OR653PvJGIFfk2mhVIlHcL/5/ACQXkWWdzsYoWNO1HonG+L
rxxLiL1dpEOKwr2qGxcz/KFg6YJMpRK+Pazwocp2V6INCFrAzwe/r4uIemNugQSy
+wYJRWMgqtq3jvy12CwzstiOatc4Z1nlme4+kSgSFJsPjnk3eKvRQAFfpw6IaYD9
8cpQg6b4PWe/8gKkPHemNgJB2XdfTpoir3CuLgCE5rMm1AF/6oU4TAzrRFqQ2Zhf
1EfkLsPdYHWYiMdJ17cI4Sk3mw2VntIvg35KW7x0VeXZn44DsrZodRr5gDQ3/Vv2
sBmL35Gfc/ZewGSks1xn+4R7O0T3fxKaqNd25vq3BwOh+qx7zp0JBp3srPbz6s/7
fCnkKtH19lSPs+3GGbUV/LKwtzcxolv/k7kZ/hJ1cPcox/WMA1toqadOpk6tsa7Y
lsQeHGpe7M+EMvO3owsKQ7WvE8Jy/4bw3eyLcKVmiZbuZcVD3rQrW1q9fNIaPAEO
DCOHGFpRd8K6Y/2mQ9Xlu9Z49aWPLxWjs4Erwqgs6q0D4ep3ILVqnXMfBdSuDFxX
gHN2N8gtzH92N1w+zpDeIEIfqlrr35wVKs/wFvaiJQ0ggWQ64HcKnTivKVzmGROd
XTwlpiyzdoijtgkjO3i53zfFBKRTWhe3MXhVBzTpo5rrtz3pj/pk6uJ1OgZmbs+U
dTqh9P5YaLieoJLZA5EYY7tfWUE64qAZxGg1zAyBZzjm2nh7uubyyAEMVqHgk18r
Z/K7eNllmSTa1Ybg1txDfnmk+e/2Wtp5w7zCQqCMb107RP+RZpiX4/OlXx2BSjGF
vFkl7izfQpyVEsh5WEcngPLbOAYYWgAwqSjsYJeZw2LRsuhxamePf1AxvMsBU9zF
/zgl7a9k09KBGT921QsMFii0QH/9Bexq3iYvRlUESfHj/+m8VwQqkiIaFWOdPcIZ
SQlAa+s/x7KhWEYR91XrkDEgIhaNP6binD4WG0rKBpRhYkKCdKg1Z56UV80pn5ig
UX9KGUWeShBfZqjL6S47MLyHUkMvFxUUl+lo+2zmQBW5bTBPwvDA5H37lP9nFUeY
h1JjimiM5b5jsoQjn/CVWkMkmeMKz6z6MaHtX9FC/imfwY1rV4yCQ8ayKT5wu6OW
5HltawEOoaB/mz6z9i7udBa1K7HktY/d79xW+KxvnrxBf09bYgMH6u09yGxwCPz7
Xrh4FCGigZwFnYEf/ti035WLr8YGmWt186YfsvnW/Kapl5GWkfRSyp8QeWlG3tId
5IYEhK0piRhWJQ8On+ST0NinGts2Ip1jV/2g67lx5nETAlcHwSst6IE3M0gEt1PK
egfXxJZ9LMvUoKu/6BNix0rLFfGXDWGb/ttA9Wen+xjgFAlFoZPOSuFxHHWfTuKE
P+NTAxAxlqxIa/ZkftxKJQHdvCEArqSkv38Uwxsix9RI+wiGsSIOO1dmNasWkbme
XVQ0wsg8Is/M17Dh50njCKdh1I1sg46Qju2FZ0zq9rjD+WGNza9247mDO2fVMqC9
XOOXX2M9JL/B1HvEh7pObyppBQQbiVmO6SfmoTMDvQKTiHXifoCbYonfuhRGz6JX
KoaJOEBVHF5347Qc6btcZtsTl5RBl9rQ0jvW+DzrYVo8wCavDnqYR2hLM7u/nCA1
ceekfWL9j6OXIuIumhVWNQacK2lMcRpDGwUL7Ux6GU3RljW50J6uJiL0Ec0tzEl9
RJeLuKVYUhl7GGOfvK3HunHCEfrCAPiLdTTmvktYy+pIZwlemkP3K53GwDFzgv5h
JGmtvzBQntT9M8zZSFWt0g3Mi7EgZKVIZBVviCkCORMkEvTxXXggEitrmK5uZor1
jATFlWbModMYhob27xkeeLDJfFVipWuWlMD516qeAIFr0OTlW5mgJV+yAxtO1ZOY
7enzxohQVSTnKx0MLr3tK1MJxY2JHjGuHc9mA6tLUeMhFAfPQ+j6Q80gxE88RR6Z
4GkBjfZb6xEdAlrbZZKkfFxYR/ckmJdKwnaSeMo0c9rG+vudr5KXgaT6xAkg07xq
xG4kto673cKGw3fU1vsH9XMBeX/qA5L4ShFnlssnlSY4kXshXqJst42moAAI7+ZM
Ds0uTurTPP7HWtjS14dsmLqXjJgQ+UkvQX+lotNgP/JEwzDMbC2uU3Rnl/0l9hdZ
CLZhfSAih66h1ei60qbs2q6kYO/qPp+phtP49GSyG2zYR3HLSk9b9M3d1HLCrGOu
hlgcFKTiCQg9b7rWBGSRp4OgLG6KJExf4Xlm/vk690OgUjKo717Lq88rghuwVZaC
6PcHcdnh4aYkmhzFskj2sN3xvw7nYoaoGbG6y1KDwDLZV2K/4Bq4wqviTflqxafx
2hLcNe6vKmppWpz6OU1qXpD8ddTSD0ZYpB17AYHvwp1XUiyvWXR/ouCQdpKNeatd
xqRo98qAOB8uTNHZpy9VtxhkBYHxO2p/bew1V7Ig9Vj9VofLAXux48gukZBP3uzL
H5QdeE2Mtdg3i7w3TX7VH65vSF+doHT44luOoQubu0AzXADtuSFIX1J8ZjXW3GgU
FHmOyh5pszr9QpLpszUDiI138PyUL8p2eNE8wJdLHGbskMjBs3Oo8poOq4cgkEOQ
n8byQnQLlUNVwCG8+jCjp/ccd3Rre/sBqJKELcUyyaPD5lvghDVlNp95fugAe0U/
/IyZsyk4jDJdjHn6BegtfN241DmC1dl0B8jU4yS5MJZeWo7U8TUrqd00wnKwaenR
nRPMm20lpIaUMljAcVWkWewz8NK517QZlC1iDmN8WOppOSm2rHkm2JnPvSZDwbG9
8bktl0PS9Nt11XzTSPc723v/4n+jKSZa1rvIixEa1MdXASo+Uq5ydb7EqekWOF4N
/rSryFWncAB5mj5WZo69FgYJYfGVHsVlJ71BUOlLq1Szl/o+qvj2s/TV8B6jfXF2
JEhO0JwTfqWk9ce02cB6jot613DyqgZchgfjSnKzBUinyDtQ5N4UmMP9oC371izc
pRyCkoovbPso4jQSgUHlcAASUDdJXz+5LQGk04l/etYBQPCIVp3etzq+//yIm5bx
c/4WDrtgkagJXW67N2noJxoEgEvWLEKDnEsuTTr1wZyVu/Sl0mg9VHpvTlDs787l
EXwBZZklQD0kjaxV3EeWmlz4XRtpH6MiMhyn91NIcO1zXe3ROxn84QUzVdJVNu3a
XBJeMJ30z6+xywhl0p6f5p8Q2feBTAtJxLtc0dMXHA38EFtH5NAIvS8x5658bzMx
9daDa+xADN3AfZ4wEmJ5PIVc+42m0ZerHNt48msZYWZLWgHCIGN9NzfiV6H9YZBR
Ztavtc+TqYlDGelCyWoX1EfrXtyiPk4VpwSckpcVejhXx3QnWuVTLVdulo0Q7Agc
P4ibuDeZhLFZEnt/zCxwfV218bHtHzWT2dNqD55ECqd1ivZKYroPKn2F9MQJ7Wkm
fcbq6DgtfDdnA0aZnl48/jWzWR5t8sXDbEr/qPoZltO1jOxLzv0Sdn1cNEKQV4Mb
tvruFcwAbtWj2taSpH8dOox/di1DBpCV1uGwSQ1rQeRcqUjV+WXt+5RCfOL7ZrOA
1TTxPeLW6C7npUeb/RUTARVb/JuhnHASuK7ZhgQ12wKNbjFpDDnHmGRBi335BxnC
D4YkvvLea94WMPp0y2NpnLA5Fj8RCxpX9dg7MgPgRGZKM2e6mdNClfwsJHC5g6MN
yeiPnGz/Y2c6sXgX0fwje2rlrZEdylP1kdrSKMrSxQbo48CJcWacnmYXiHZukIs3
xks8uHfxfrXM85iFS8tUbF7xrPtUekAyJhpwyYlc3XBfaktJ7tQ/t74ndLF9u3SN
8cshqd0X6G6mj4zex5Bl23kml4tfC20DojgkT8oMa/gKrBhOktYySniBXeMwChiK
0wZjcieyYVvFdqldv9Uyff8W/+xGZqZo3s7uO4MvtHqp5ikI1HVhtez6cyaGChJi
WqG0y/AU4lSxdEAWl9UQ++OQUw2VdLkIechHsn5nY7EFBpneAA/mCoLe/hIznMDG
fZqu2c4W+Q4Nsaz5niQZqXYtZ2piAe/u49LwwVAsqGAvb4gyMlWXwk3XP4SFUqQP
VImRxDUUJ1QyObwE5soHltXK6p7eJ9isCXv2oWrNTe38ltC9yYBzV/CjWPybIuUI
ekz9kszuyjE3ozCg9ZuzCBOQe516tg9mO4JmN1CrNfqRvtQPLpaGEvAMzQ/w6wrJ
RlS5qeaJg/yMZBIujbQSyyxBDxoWW2ORJEzZPhDPsI9p9SQRqTLnksPEcyiiTLC3
LU+0I7N1i+EzT8yTUrPhDSvl+8XjSFAbGIP/osj2wC7LWH4bXqA0r4aOYPqGRXKE
nxl6EWGxNp3stZlQhYYgkRIGq2uu+rJk/Ap4BvGOtuNOysxH+RHrqMZ9PwVK7hJA
jHD7M1AK7mpmnlU48xv0flLerlF6rojzAlV0QqN5CclPs+gmjiaTW5Et4ryXlHgw
avlHXoiu68JEURGAy2C3l1Lod61VrD2BA1EGepyX5ltJXL7p7UwKXZz2Dat9/jqF
IlOIcu/U4VKqXRvoRqFsppmJ7rypdP4a0z3Y17pD+zKHt4xulA3fRFJIxGVI78+E
FnZsLgfoULuQz8Lgc1pVJc3h0Oxrl9EHdNaq0/ZJDjqP+TXT1RI14VKefurXD5sU
bkXqY2s745VVg/6Sg0TEisEhMv0pTA1Mdib5SO48L47WvqyBsQ5u03t2wbyuDdoh
xX6e2KfJ+Be7flI19UEh3Q3kHEknmA/l6r8YTGKXMIYXo7cOZObZ5pZfqLSkQwla
P8rm+CJULkVUtFypqTHd0B/p/2UhW2+M7Vuz2KDT5c9oaSPn2oha8VkEUurNfiZo
5i4hUljfCz5v/qoeErBHqvlF3oF/QgS04KZ5dPys3EUiVt+IsUqOiJjqI974CG+f
VPeT+dHaKiR+HnbkFrZONbScUNWyyO9OhiQbsrJlef8wjoTl5l3HiVGwpCcc5xYS
/pRGjw5N0wPgmBHZ/NZx2K+CQHAZrInV0oo/0yD7BU8mfe5nnD7lpvWc/EzAv6y6
YolY5O2Ziy4kP4jgsPaW5AOtMQIqJmQ00xZ9K6+VVkgnsu7LvilK3JN60CwvUqMF
TwmzmQTkKPJHji9bP2Alf6OSoBPuyyF7evkhtuxsgXX+5QUCe5Bfyoki6SS5krdP
NY05KpvjO2oTfnIB0bAsPnIeFv/tuzhB1Wm40k5P3dSZ+DUakAEdO2cHxHLBmg9Z
A7IriZTuHJcUP5c9thRPC/GIcvQcOiE3jwnVSWidAVT/LqeOgaOYhY8Y1oLX+VLT
+6IO//WzAulIiuimc2lRpaQZGtPkQ49Xd+B+EbuRUpMOOyjUuy/nMufT6AwVrM9a
VpmPWvhXD2gMpW1I8t6GS+H1fxXzwevpe7pAE6T3zKb0w1SBe10CrTwAQ4g42wG1
/GhB0yHs02V2pI+pDqUFNQ==
`protect END_PROTECTED
