`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DXZWFmWPnanJKf2qD6+1Q55H1AhJ/f6t5JdheZpbiw1aJASoZplLMIhEANXjYCkl
IeZ6VxqGJAETYax1Qhj8kUDQHjP5LXKLEFmIX9/9Vg/VOdRSlKRygkX+y1iLrdy4
H+srN+wZMdCPNpEVRgJ+twUVr60tohVWAk+0mpHz01zlRMNSaUJYbVVwvtIKDsVe
DhSwR5oHlu2mTxQ/EzlRMOtAixq9Umk6YpPCyAZFwr6ecaypf3SDAqEBsHJV8Np6
iqcnuvaFuTjVqhNSNIACXrROpkbtPWs3Qjjsb5khzlp9yyW879R30cPbgvKi2t3K
n3DqxPw3VjjvchMzCY6+/2bOnjqKXBNUKNEdlJYwd7GjZqXbwR/riSW0cuYGBziM
tyCSjx5wJpaOdghpvZPOvvXZ3EAeusd+k9RLpAaWBg7GMK/B/RHx/Kc8mESkMx98
yjAX1deM+EP7xbe6mJ9MxCpd8IKHu+xY94XnQVeICDu9L5ddhHVyHNu2rUce137n
l0leEVoBWjspFvZOvU3m9AcfV6kTUWiLAjfL6XP4GNcmjJKtaAGSE1XLxpGlUBwo
j+Tt0Nmy1y7YFxKelvUsg4S6iOOv8dWWIrJz0bogJMGkXwrzumMluD0G56UBsBZL
Op1JMZ9mYlpVX+AoHcwVI0lag0DQGfWqUVSAw9aNSNTrUm7Grx8W+NBPPo2ZxRVW
R7N37uAmqxfYtepRnkZMkw75+pXxXdN0gtm1/RIzTg4W2RSXHrNhM/Xj0VK/k4mk
Ocd/qxx8+UUa4RY9R9WLrxkh9/7gW01ZFkB5orclz9aoLHje+HkNaee9qHN7XQGy
hgH+Fp0rUVhv4IZVII9T6nSE324VaQQo0CQf3hEWhYoOCLHQSfS8PlbB+EtDbSMO
i97BkXWVjctO+oIFV23U9bXM+dfNg0d/FuZ6uziX8wAeBsJfU1S4/frnoIO3CNUI
o71ac4GahIcxAzn5a9F3T2YSrpiTLLvQLUDRLcvW9R6jjIH1HUFQQTA9XY9CTpp+
tAvqBzgW/xJHqMubUGZaHsg3FIOFFOzB/9Q0UxY1LpfkXWve240TO96HmuvrISnD
J87oGb9YSRFtjmia2EbyRICvw9/Z2SVdxjkJQgwM3hJ7/ircIygYEeSM5on9V8eG
qqbMNCwvBEnyFUiH0KNQfE23c4aQFZjZnozjJVPmdZJjx96IOdvjZwvhg3BImxl/
y2u/jSMiHqP/UwKpAjYZXrQnXaLDEOfmT3GmwM5SJpViv2BAkS5ASmRy7bH4j37a
n0vJ5CM/Jy9F5I48Wkd4npvbzVT7OIdvZDKcW/L3XP+KGU4WqRq7RaAcroDL11fv
kA9V4QNsJz4kHAP7wG80LGNC4vcCXu99ISnniFyAjQZYCW4FNrCQZDZ650fbBlzj
jIgGfwQRn8hslgUbw3m2YVDo8O8+ROoMLWU5ROKMiwiP7Elb2drezNr7eALI8xSp
a5oSFPNa/9npfzuhgEU30WbajW3+Q8LGPW4f+BW7y27gKGTjcF+NBCEt1kILZrmo
tWDXP+8xHpuruXIETnTbzIrllGOM0M57dII5LBNaYl6Uh6EIIAmqiUNknxDVV3C+
xI7a9Q2UG9kyCY1UZh4o2NDMnHXBPLUWwbD7/xoYU+APe3KGOqsuCK1GBTa00NoX
bkwkfg5mXAY+aB5/2W9xHNN/sQ3p4FcjLsB/RTWWdqA6XGnOMp6ByPgSLw39xGji
EK3LrQYksCt1NLVrDCsKT/K4QfQHzPQfPMYryShSS2CbwLV2Z9AuQH0+8tNX8knd
femKm8wbQDVxebJVxVNjjMhx5f4ADP6f9TsjPW4JdSnCmZZUxzSwQK3jbBz36oMS
oQVyfQPvc2zPdOLbRdLKO4OoBuyfCw/KjWarlFNsrJn3nVHaSqn7NSl1mC1e4zJ/
gk4bpFY4r3OapZl6qz9oKkRvt6w7o3Mrwqo2gw8l2eAhm27cCyB5B7EgBBHR9M3d
9mJuH1WB6S5+lQoZE+V2/TvJ5pAKSP7y36Dg6zzymPTioOPbqYFukuYH8/r3ToD6
aS2FmjnBMNww8kfZbMGcXGeNSHmrUgUUoNr7jhaLz/6b2UeptZAiAR06hUiLwtNd
VjvYTZhMWiyMz5NT11/i+dEoQu0r7bDVHf7IsaGyysN6A63SigwoUoF8d2kJhhba
5EFP36BFM4FC5/EDBvdj4RT2R9i/YnBn7FKrM9T4yCXIhk1F5O3OiLssLIkyKoKV
EqfaOfneD0nce7zevTnHQj9V8sntak8+Tk+JSLLnuYFFBtUEgM3HfeI1J968vHb/
wWXWVsSVGeIUtCGuwXhiVO8vDApSIsjKEneZrzbF2WINQh6nATlYlyzrJKC3f0vX
Vld4wJG7bosfrL3Daf2oQDU0TsBTX9nn1Vm5MhNNGVgZyVhAMyswb9dR3CdM5n/g
obwzIsVwLeTaW2W+/SR5B2ce6zXq0gXUicfbu3irBvrMJIf0tb4+bpnOW5KRnG6s
OxAPnC6LMWrYhh0GBxg2BvJWfbjcobMgWN3HijjPRYPRRsfiEpLAqVLxnFnXg1mH
seAXhWotsXMbOn7co//xXf0VpCv7h3DzQ9+ylTqS1xjYe5dfOjbaj56Yin46WHLY
5CeSAs/glOE7mkgOhaZOTjNXd4G2b2PFtrxPK5nvIakaIiF6wOc+9K1Zsr8JhQMb
hqSBQQcBZungkoydghYVD5iKFB17HSjwm4e3IJqTOOjFOAit2K4FAt3h1/GQha1G
YO8Xh48BhILuVytfFflTnoYPTzAPpQnxs5VyhVsPWrmF9/mjmlkEKGE+8GRLweD1
fQQVmNS3XbiJ/7LBSKBUNOZI2DMcfWYTgPFvt6YMfRmR+SuvTlgstWRoPWwh56L9
4yz9BDzBW6dC/XJPLHRF8IKvVVEpC8F3xVZ5fcQ0pMkMMWxpGTO6voRVTM/H1wA9
R/xi46UKk5Wr9SI1K1AS6jBoYEJ8WNr8u36GoGZwZrEydFNLtyYcTu3+JLPD3KHO
DRu8+ZbvFl364sXDzcPNPnPWNxcWWkhcHn5iO8DhViTkmI2+/M2S/oWeVRQnA6Z/
FRaYumDraGdoosLN17REQC2hfZ9RRB6/77D+PuGeVIVsyjrtsnxYImPoloC9FD0A
AGHxDkp87I8WSlg1XyowAOWscg3uNjoFc9B+0MXZKdUQeOPAZOW4sp7wFgCnIAr9
iVPyKudMqQYxcZDYltHckXxIPUqVkdaFXYHzFEkr+VqZocRJYhkjX68z0W6XpvX6
v5+vK2e9GBBsrEXkcJVJTXKkC51OYWdQkAflTtoktxIucMF336tKmVT9vttIBlH1
Xy4cWDUjYm885PKmHzwW6fX46q0VhdgJjQ7qlh2YnGgP/JhG3o6h3K2wy2Bqhvm/
YwmX9ReVv58z7zBp//K0IbuNSw2VijsjGuTxmJQkSKQFVrCveNfjbVbJNcG7jJmY
OGSxSl5/9G+Y0bo7KHryKg1kwO//OEQYcmnnQpvxUMYjmDiu5jdgvlIaLsoN//HW
tMrP00UsPoPgAQhvsts0gEDmylYYXuamP9I9QcZkgN+ffm9SX7FZzrrd0zqh/v0d
jcCWjqTI9BnC0V7r7YnEU+UsfiJu2EPQpZ14ThvCDSgRWcoovxNcDJamtrGrIYMO
`protect END_PROTECTED
