`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GA+J3yyUPvFLEIqhET5iQT4T6WANdpP5G7W0yj5gYvZ6TGNt6zDDXdFdj53K2Vjk
ydLDr+a3Iusait88ng9GzOCWxvc8Q2gA5l/O2cTkAZcXdo8C1Xh6L9/YXTmsgPYc
m1TtfgkymnIhFzLAMVbEcM1mpk9wHSYwAr1jmkHXHm58rN9QlQLvIAoHmfnccwDb
fYS1NkJUWgFugbuJfkJib5hOJ+oHOgG4mIIJgQOrxPlMfj57QVXzHr7r/xfyAdCB
lIGmIaCowE3MOblCIqDeFENO9kvcItxUm8atMRfTa49Zb+ZrIVmdPfWImk9ZEY9b
sb0pXY/ibgCCDapBXWylfMmLWEQFrzFSSbnMY9t9mqvGseMI9sPpl58TOtu6wzJr
P9x2GDoSPppRF1FDRobfBpEE6faAE7w9pDmCRz6Ip8r0L9H7wgvJiqOlMOu7hx+I
TI9KR1k7ccLn4IvMvemFbM5dxzBFUze2zLt9TL7Yix+VVk5jfpsfDRIG+h2UzY1r
z4OsnVjv5nZKt27zb7xLMRvf+dL/WV4yqMl/8xSCvtdDTqus7dyPHnF7BhZUG412
pEW24L/l+hsfawRinPzWHH2HdEgXjuS1bR1PO/q4k/CG2F+Yf+4yBWlOD78A/4Xi
Z9z4rCs6zXBfyQslfYq08Bb1FfEfoJhGTLJjGKNQ+jR5B0+7YxqYKpGkk/qMvUZf
0WVZJuOJ8qbZy8wZ9JoaBiM3IG22Pd657sWQXa/L8DWj9uCnvuWyL8ajOrSOLBQK
+/xX+R019SCcfsLjeyPRyVDHMfv+1YAM2cBVpZ4kEf7WzmajZIabDFgOkn0W0pWJ
EAShCKQeUW+PAPdq0A9o0vXnVTP3V4rerjBPbX+4ohIWCS5OUzyILg7EhYg1euKZ
YB74/ea5qiLqnuN5qOwICoipg4tgzNtCIaeh1KnHto8CHEaJHgxTakg+37wLQoQG
RFyn84N/DeTupjc9peSpmanTk9AeTJLBk9EBzxM4rn42bmDgNgNpoc8nlBkFLFSO
g+NvFtKgyPKVh/b+saPruYauWl8KC87F+PZKkTYGuUN1wDFfU6BMx919l845ypVU
8i+CJeTpxWt/ACeOZa7hSb6KGhgyRZO5OKfZp7j+dVUmof2oG9ENgXTW0O6ZJOuo
d+n0fcAVOFsD1ND0k9s8QDUcgCGycuue2k2YQS2ctgefwa3FI5axyPLOuRtc3n7S
`protect END_PROTECTED
