`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aFSWVvE5wRV7Idta7Ddo6nh8YrogJooLAH6g2WPF5EcaJoKggKagtUTCHj4xG4lO
W7IINUhCVnW8FdNrCdOAATwV6xbw1Jc4LjALNBLUnc9omDMd8E3awLNoqiAEiCmG
UrtGSaAGOLwFcPjHcj+TLtRu277PEcSXEqKRf9hOgThFmrWfgt42WwZtXqDe+x56
b7rkAIWON29L+Akp8a7J/5wnYc1jsMoJ4MkB8GnZ3c3M+9Vy4YNJ1t6RIUzQ2WCa
M38AI9Y+V6NWwQK3TxYzDkGlC9Qi3+K8JK/JhgR9OdXGnw9oKVW1SrDJTvnKzWe+
8DIIfGHIpUNfnvkBPJQNwqQLmAQ5NgORja2XVMw0AlujXfpql4mvlNTRU+L3XBWe
QaKhcmBG2Jk3eQkTOv/Shmoq4UVQaYhE4bBDWtdbOld2KAjY3WE/OpxfsrW4F4Sh
DAxD4XXXjjv8XfTsS5uhbOy2pSa++LvBnCJ+4iGHCPTEKav5ZHpfFilLeWQZV4iY
rya2dtWiXWWPx8BSEfvsDwiaVveAvZl8AlS7BeSN6rAUKitKDM32OG+meUf0My1l
CkjUaSuWWUfUqjgzNUTNcem6eNxjhjzEfIRKy+LlG2LEcIPovQd3/D1JFKymwdNX
/kou/bV3hlio7spDr6geMIoHUTqf4+feo5I6HlY2GsHPvcuybCv3cPpE6lOWfWtZ
tpRbT0EoIGSVnuF67WUUW0MXjZGMbmTs8pS7nxBnjSS0mFwCCuvw5A9YL2ZjCrrW
ASibziT56JVuOU0NVEfL9JU4sXlBoasn+c4Pal5z+axrltUyf1Uuws3DSj55Nq0K
ik8peB00k3Xt1mJEFUTCjNapVvnpNeRwLk1IZB7fGo8Pu/9NR9GkiM6J7reFQxQ/
NyooulrV6AfARYdxjx2nWsg9N450lpQA7V/7K3YUzXzk2S+FlZI9F37pzh+intOG
eqV25KpxvU9HDI/Fg+VWH4WegOfZtaucDVcM/ueR8FEta6d4tsxC5L4c7EM7PwpM
fzgkKwpv4v66NopxyR9o0ySnx8HXBfQR2+qqFXthhZl/Sa3P5szkHY/eRWUdtP/n
9ujsyWjRlm4cPHigeVa3Oo7dnmnH3s5NS4CPk8mchmhAPH09DzjW7/u+CvRrk8Ik
G3Ue9LufMG5GNveWpAdZhGxolApVkTX9xyoaTsHkq+BPGFpUWcx0DK9auiVgVn1U
Vi2JMInvneZZHRuY6VuxKZTKaxy4zWqB/xU/S8yiUswq16kfA0Zb5lDkQPaXiiqL
TPwaMTYzD+IpdE8eif6qYzWvDKCcqIc2nRxrYrHMgUwEZxHBM2y2FJs0LHSOCJSX
slq1aP5SiqYKcVMyGN3V9u982pAys6NdivxKLOgSKcDV+Umm/eo1wm2ymKLLeAE6
xiQTXvHoBTlSwuRNYXSD2BZDNIgO6qXEQ0sUQcHEwkEHygQZArK20rDyeSLXdIT6
psveSRh/oc9dxd4mIY0M2+PEgD8uy8uuZy7a4TBH4dp6V10c1H1rF+RV9fXq2lc2
feo7GPSjp2v08iJU58PvQvv112JWkqE/77DwIFdhpEwGnmVoj/uqKBdIMQlefhBC
IutNUFH5eYCHJ9Uz8VaOrswGuYgs9N/vOJRnWP/2QuG15PHpA5sTAtXtzuNxvN/n
KX/Ex7UU3/is9C8+c8Mr2mJA4MrBo1058ab/Qb7zTDSh1AyVUPfzyKiz/T7ZPNBq
6jlTG7vo1bzsEjqXZeEwwJMFspQDKImhhxo3iqYG2BlFOi/UMmL6YxN4mLwW/ZQy
px1yaQK4YFFd3zrwefbshkCDShXpdYYPJ6dIOLn3wlbuFyXLM7tzmOpb4bB4sKYu
6v8Dlyv15dXXSS3Vfp0HK4fenR0c3vU+yjdY9wdP5YdZSoaiTwU2Cz93XZCWzyqz
rvZB/+8xBp+yesQao2fC/BwJHox6z5ZNXNf9MUUWYTBbo75BzbAoyiyb63KMGKrR
dtH6U15iIj81YdkNaWzH+4QiCfUngNU6446lFJabXlnmAc++a8Au1OsBtGOq34a0
U0+R7L8GxdBkEpz8NhY6ReTbUelMfWP4Un413SPz/lQtTWJZw2OoDIKkhJR3wwLz
LnDekRNknFayCAd0cXlI2Y114Z0J+H0xPzXmpA36o6KsH9VTDbG+Pg5Yb4ow3Nkb
B7Kp9jnkW/zfUufBK9gklsACMzZO9tytTYeFEojUcoaLa2tfU1U2WSas72jYGj+a
cPHl8w+j1bjaAarmeyJqjOMWk6TfAA4Mia/uIrlrBehNT/nLuB88JoHoKee6wWBa
x8hhlInjY9lVKK2doQPOOqFduqVyWtgGK6PE57nGI1N34NLbSmN28zf+SBF/tTqG
E5ofPFzougPQ5jyw3HcbM2LQiVp+NAyUkOzT3MvU7NKkz7EgFDDx3ESrMx1BqPJ3
TpLtUQ2Sm+NYFz4H+bJJ4Xms0JF/EYlxn+pZiDjRh1BZl1qDUuaD5WSl9sroHLs1
FHVGj7kFkOkTsbh/uVESzETwWeHqm0S3S359TtiygtJ7A+SEMjtG+sku7OT81a61
eAZhw29X9Ub0AmSwtgFwz6dFqo9NFbcu7KyNyju24gFxzkGsHl1h5QxitoP2EBPw
CgdKtD2XqfZvcYoxgkcfm5/r0QtEIRdShcL96D4oSegkFaDDUl7EVBVTlxvUN0L3
agjgrLxI8QxPj0rGQ7cIgOvXWI1hk6qUCQRsJVNhI7iw6gjFszUotic7MDiRuUza
nOnzvmjsMdS6sfC7TbN2nqoYEbj/Vd5ykEBH6ZMk2ZvPv2IDNzYER2xzBmpfW/KV
x0QBg2WGW+t4OOXNWsbDN66VO5I40HQL8mgc2si7vCybV3EhtFICvJ3un2jT1yZ2
IojaE41YborywCPwHJFWOXJFYOMiBI3vb5eVDxlSpzCHh0eQGRspJ1rfFGhol85w
56Oa6vG8eNqcDVQY6btNjT593VmWa6LhVr3Uwh8setoRYCjSVXCx8HaBFViW6PdI
/S7H/tkrO+HYcOTgK3PryPzjFZJYUrx8gT6KEzdgcxoSzSpTvESyMTbyC50CyjVY
26bpO5vB8TpE5ncmF9Bj0EToH3naLFutaey4U3DwssY7GfbFXfmCiaf564yXZu2D
QCeUVTSwg0qPuVC0A9CwBWo6WZPiCMvJi/f4aHhBbWQ0JGGe9m3cceOCwcpiRTtI
zqRvSV4Pm7Z2XtpErB8SrKVtt8L4PScwUIoehyO0upEKJy6ATEoKy7jw/kQ1OZb6
ezbib4QJiUcb3ULxsSnGWXlnkBwfsA3TI0NVs3JKKrrIz+P+14YOg0/y5mDUkzQY
ZTj4Bpupq4fB/ObX14eJ125vZDykukMVm8g8qB8PpcRe6dT6WqmyD9iSfO0dUuSZ
BWGebK+dI+xNknik9Qp99d6pY0hR6th5nloM1mD3FOjTVEBisH5e3jRVbgCvAlIi
2P+2UMq3RRz10/sp152RDce4bRDjnMBtpZP83PuxDhRN8hOGIenP43wzIwxp+ket
hjvpltFBfo6JqQxDrBVF16jmF1dO3JFH+q0IXtDvDfCtjYDqo1bw5H6WK0cW5/8K
HF0fBEa1cTpI3eboaEtoi/uYTphaVIzltfXN6lI4pZaecW4ZpDeCp4v5MA67rOiX
pQoexXSZY/nitwIhhjv3y33UH9mHl9LPNSws3VGIY9LzMFo0HNSS3zGepiKwZtA0
JE7JCLiFmDQHUMv+b9uZ2pIGsyL+TXVLRuo8eFMSmFAgIkJwlGiWBB1CSklHQqQ4
cMMHqUNn8jKi8R0N2WuEqItnF2CMgGH1QaiCCG3MB28OaJD9l8VeT6U0qa3tnHRT
o4M3vDeAPCtPAtt4KwN1mdyvk37LZKcW4z0BMMKjIs2vv0/OV8eVIcIFh8ag7rst
h86QyhT6q60C3/jpD1mW5pEcPCzTRGFzm/zEtnfkXa44v2WIUV9u37e+WH3mrjex
xh23kIVsvyECGOu65q9r1a2Yoh6GYHTnukGrdBiXH/k=
`protect END_PROTECTED
