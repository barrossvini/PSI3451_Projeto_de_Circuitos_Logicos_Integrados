`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UEQLdpldUXeruQ4SwRFwvQ+X75tG6SnaHZ5TtGtvXQyuhhJ0NNV6RnX/KWHMxLxL
7mV9exDVsxctoIMwegGp2jgL7UaOKYqW1e8je5dWZNYjSTJ3Ild7XrHVUmddHPCz
e7t2H3j3UGOIRQSHClZNmcixHE1muoM5Hn1yuzSUjCfdoC2NMgsA3DOk2ot/kwAZ
fyTSdkiZG2DkTllcqn6H8+0MsDWq8JI1OAQMxaE1lXNo5d7Oru0KGp4nxJ7rqb5X
vvFo+fmzIS5XjK6m2JxgwqVBU58VpZBnVwkV/MAPLUp+oyBWglaKX87M0I+QJl/Y
8Wc6yvy+hS6sLFaEBz7NN9K/bXCuHjHeJjWSZ/734ayZE5gmeEP0cbUSRdH4GxAu
++guCa+/KeyDSxLRAwTzIXNaQhm1qXGDUUxnd130MJgaKRj4ytAklK93CIvkB2K4
0V6cfAaMcC7YGIG2I0mGyPlE4/8gaKviMqmrZp1geeMw6OO0k1EpQHMVs6TTByqF
0YTxxbADgdvwFLcE0Und/BGs7gRXZJfNon2paEDaP+ca3kF6sfY9ezpkLiHxDgGP
7L+RMQP0FuR/08lbZqqBxNkYsvZOHXCl0XIFG7+GgBiDTR1/lBiBAfR4GHOlvn5u
P3viR9yDUjambhN7ONBqe4qxg8FBqzYkXCe7I7wsWPqux4q4Zy4O8HwKxGcXFh71
rtirf908Ph+Sayyd7KM1Rqm8nWjK0seWt7z30eWCRM7TD9EaMnCtuXe2wBZnCr3T
pCPfctFqdtnmUXwIj4N9RgJxwGj7+PTn64c1ooXogyzq2nwHiypM3JAWIt2GXMr+
70JDs5TEVEd4lp57Ym7BZH6mEDIaILZUgQhSp+eK9dexLuaPcORFBfIrFxbxrlTH
orPIfo/hLpeg0JxLK+1KgdZo5zlnT3sb0TuyEsAPXt9KWqIBNx5FbQ2Ent6aa1z1
HO3toceO48yQfYht3UurlWP0X/Q4HLEW4tjHTcJwZK6HMNXkZN600HWzbMCILesj
qrcn5ChEMD7VqkneSc+1ALP2jL1x82YgLk/MB32UBD+kOpiGjkYckf7931JZD7qw
JrtnXTrdidoXs1KshH0dtrgbZ/8Vl07DiZRTHfXpM9NPBexbW0jJKNHUNflRZ5b1
i56L4KVbyGiSFqcK0dbLi0MmAaP3Ql4hutGCGPZJOCSAIlikHCOn8oMn1EV0MgRG
6G8G5kUFth0l48s/1uXK7zhtuZgvOKSeLjM3LwLr+16NEmjUIfxHialqltzeRerh
PX3qFnqgl2BrnebSZmAdI9clLdbQzm8WR10C4S/aSZC1iFQYFh8/lmZZKZFpG2rk
Tn3ewUMnNDXh81rwdKt7o5kQaS7iaxFEcIyAGe7FbHP+Z2G3/osUWSHtD4pZunAh
xKkDJ9uKNHF+E4YnkheYZhbNqGME3441jlFpQU+KjjLP62eELv7u9xi1fOq6tXlr
aChSy0gKCd4FQt9Hg664MaHw5QSGTGzrAMfCBwOXwmbvWJ5YuymkYSTe5+IZYdA3
QwRJGiYqcPHa+96+ryHjmpZseZFsiw/j8OpU84huTEZX0yMMLhiAlx1OsMud+wxt
TibCzy3OSoG3guzj99vn7VRg19TDyyQSrSypuwn3P4SKajjsU/zwhjRLv8UxQT1i
s6zvkVdfv+Tvzwd2rNGTn7s091pP3ZwfHu3Zm7rAyqUKt4Rt7A2IGtx5YERnCMM+
czz2CmykQss3eEto4qMDFCoQNPdwc9HuBICx5NKhRFrqY6KUL/TKtttu/5fOTt1Z
a7A/0NjAYm+yjHOg+qEWJhCT8iqkPj5IO+NHvUQRAkYWomNbsl1CphBWdo1GYptB
VvfeoWFqUmM9whWhKazIWJVapQ+Tr2CIDzKIw4oLYWw7gQobD/OMTLvGb7LrcRD3
vznU7Nny4pIIaTD3V++tYUhXhK21qaw8q38KrGAleM7bWZVrP58QsVx6CgHRVkMj
chhmCHwH5Qi5tUEye/SO/lLYdQimid0N8I4W2VA1XaR3HUkQ77zU1/cYHOY3O7cu
b6+hVDr9Lx6P3drMa010rrLgfmK3n33H9AS2hi+C8cjmJ5p0JN9znuUuFwSlcDJ/
81Jo8Qf901YC/djBFwCmgb0ahhCHwXm3ASXaV8IarcQRS858PH7Ih0PLfFe42wsN
VuDRl+QX5HEUhl3j05N5SSNj9gs1GOwip2AVIj0IOnY+LTmezijW3Oy6/QI8QluW
0RegHtL19OipNjMxuuTkhRYi05T4iWauvruXRGa9XaMWXPpLE2caf+Q+9oyqgRdG
uKfNmavRPaAjaHSxHuVpEdhSQST2P7jURUc6hNjlFLAlFwMCy0EA1VgIvIc7ofSl
nIBo7RnT67aHDgadJ36aSkWO5xz8mIVvkveMm03Dz7iMG9cf0WLO0B2yQ/e7saYR
MFMp7x3BWbfHuTaZIrKnKsH/P5w33Gg2Wzi+JItS5gwMnelD808P1syX1HmVzSEV
IC//9e6qI4vBm7ZAme/Skhu9ZwyaKeJLHjMZkgHa77lDw8yOEk4I2c21CG8e94Co
pBykLMWuY8bWonFuz04ATPbyCuLVXKXrHazsTjlrO1HDYXxYMMZLfeI1QkFTpsFx
KwdTvrAwQ1wOdLI7+mB5BXBsmUeFK0AOcWw9G6MExkvI/t1q34/q+WbEFEHIRXWm
8ntqRWam8oE9z4BdYndwr/2cNwpxgTY3BYwdfVAMgdPXdO76pQXWhyXe436fPlPl
BcJIKBsrUPNUCB1bvztB0Q7b7JRtYDbE/61TN046Bg5JDOBXCP3Etgg+OeQw1sTG
n7S2pleN0eOFiq3y8TdPoJ7Va/XEoSq/8oYiIaWDbHfjLHBv6YynPCOmRmY25PRu
PgDjcl/pA4uD3cDSz80zW8YVZPzFfpNRnGPD2J0YxGuD6CIiA1ztb+/w/DuMk3WS
nQy4xKLLWRwARfyCfIUeMVyt2X/0R3R4BBJptsIwcJcECj3T9eLs688pVNz8m1+s
bzPrem/1dwcFQo1c36Nt9pLJPXX34MCYKur11Dv/mjh5Si0GIbSSnxuDFPuE3cms
nenjOndefp1OOTRFp27Dygb1JaKk4jjys2GorAItANpr+CyrntBqLywUKW7Di1xX
nZ49cJ1PrwtIJi3r8dgU1e7w0ad5IYt/A8koyvCAXhcCXgooEDCQm/9KoTji7giR
24h9MQUhRmKxWPKDC5TapRu28HHUHZFKeJS0IJn+Ou8kuRgagTlZLWcy+qRbdtp0
RyHFWJRYFABkyVFVoiITDTWpSbetIFCJhlR0iJDxZTFmPumSjG4/CyLyKWGoo60y
W1sd/hBeCThZzqkWQBCfS/d8hZaLurDsH4ZUmn2iHeGfd801kFEH2OMNGsGhhz+V
JTtkdHzSI/2kf5qg8T5p6R6ZDxoeOGz8pDRN2tZKCi+OOj3vnG1Q/0VyqrYbQzPU
bkt4kUEySHjMgVBw+fw4WDEXQetuymPjGOnR5+JkSdiTghf0C82QCTpeNf5K6dcN
7AgXJWtMJX5KF49iuEDktGbb9syKvK+K3cugiczeQhPJ7UbEneBFZ77ZGT+IUQZO
edpPGwmUmVJvqjPNlve4jIpRrF9mDrwJjmDtARUS9QFijXaO5mnyIvmLzfOjlyqX
1JktyTLShS6938dD47y15hI2IEM4KwhxrPUu90C5qfYAEb/NrzcFOibAcsGT/MEo
hkpRojNcxHnqjbLkjirT5Km78A5OQPKX6prkJEZaUtfulk4DPgjA6qzb55pgkGWM
/ekPl/zhtRUpCemOQqsZrrnDsNO8cZm9tvtOjbjUmNn9kqAhkAeAYnBzvROg4mQ6
t4kKIkXhUERvn4JVJj6vnxkfc7Spi9iZV4y5d9bX/0rukl+Sz03AyTj0XwR9NYrS
BVBPB7fN1/c/9mDX8KGYMB2rR9NdlXJhvjycpr//uotj6X4K6DQO9e8tzeHMu5yT
HVQNp4JirjQyhV7YC4ekXsGLoCDzjdoo3ynd8pyD4vihSP5u1YPbh579lx0TPNb2
Lm3Aqni/LWi3uqKKM5l5mCSA+jzLyOzYGbS0dgVYAHSfP9oBG0z0rZqJcATA+lwR
14bvN8MvApmfLCGDsFeqb6VijukcU+nrFCQXUCkczfRlW8G1V0bgQAkeAhOiah0W
GqvIO4AeP++f4wC/1kWjhgu2q5jHBM4ZYh1NSOx9FgMfz1xH6ofnMUbMsSNucGYK
3BF72Ma/iczDImP3VY3dkVpibUhYLEPulLLp/Qki3GDiMV5eWt+ilDOPWTLv9AZ4
2fKUYYY3ChWxydCxD6BL1xSE2xDBVYqLl77x6qBtYYhLiEN5uelSA0T2KXWtXt/I
PxJln35oMOEMuDdYYxqlmRzIGSFUgyPjA2GTkY82dJ4u/c5gslPoIlmHZKJtkkPN
+S/cBLhmCj2Ro5RVxrGq3Je+CDq3D4QAZHv8BfPmBUucen2SLtJf/IV7TnqKRCM0
dbOJYtFClcv57w5uPPCJl0i0xe+GduXXYiA1trnTb6welPKPJzueGxOcC12/V38B
8nh1usRIEXLABhe+8eQ8jzx+ho/HGnbY0RG4JgzhdyPTySrJzmRd2W/BvNaR70W+
ItgDAz/cZ7PlPVaSACggjsgJbDD5G7JFaDnBMX65yrjsivvP6Vm2wGiNU0QAmhCV
Sm85QBsxQCLiTeRSJPhYzZcXNHAdINVyp7KhDlPFDAEmtRPOTbMjb2M4wd+oiumt
YjHMN6AnlU2lWEAf+N0+34RZk4YBi3fIwL7jZnXGA6H33tRegS8lk2WAWT9z1VP0
iKJjcOXZko0gLBriTxN2oyQXm6rQgMGPNsatq6qQnxFwx4x+6o0CwLpEujJLv+7V
YFrG1YAZRG2owuzD21HNcMGgNwpCc4uqj2CffuLsCZvWby83/0QUuZ89+4dcd/pT
F6pzq6eKHDhMsy4sS+TApXrsFVcaCP0fDczadl7nWrLKyvd+EzuOFJie8gqw/gR5
/H1Lx94LHsW0kylxRxSgQvJLsYE5HhNAofo7jqXKRpwMqWFbc1dozWdP7Kj1b4VG
3d6P9VLHCrD4UGLnuPGK3OnBLc1dzA1OTZuwyi3l52UIE5ZfVyNIHB+eAiPvNLdV
MvWeW1oMzUEOSEYaMK8EkpbOLrdUV8mHWXnvKcTYAI//fZbimign/f0mURGS+8BO
5QG1wl088+ssxHJhIS+N7Nxy2KtOlMY4Zr0luG1rxFEC6YuqkNHqfou4jxDtwrjc
GIKfK2fjhIUu7Yfg+PRSKYbHMRLHQNgkRNtP6INnClp0O0dz2M66qPcOEAFXbLaU
e0/dRfe7o/Jdlp0pofkKgMQnmlSHzP8ePjxqV4BovEFFeuIX2s7Cl+ag7nTeRRWJ
AJ3KHLqM0oVjkNrLPYVVfENLthAkOYW9cliL36Wy00/VTh6a1Zqs/xSErCUSmIH2
VZHphBbwhZgWf9TR/VM3A+O7mOerRNa6qSq1/8F4jkT2Y+4yb7NlV8Exnul7oYe1
grQa6bRM5nRL2PAUD80dNYOP5qPs00oqrGXjkNfnbG+Vu38j725Va++lRakL5H6n
weSuEHh7a0ObhdOSocn7N+YoABPwzTHGNpwG0AWekOdGj0/J6c8q8V01gqam0DbB
YWnK0yKWipVIGnVqXPt3yUmAzZ1BPi3b30GzTnumvOtx7e3KAD37A+sBp8UfzI5R
7b0jo0FAyck7u/1z88orObnfosIglBwbpn3QJjKuexSTotNsJVqBgpYcZ6iH4df2
GAMvfyIYf00y0/dLUi+gt73/fv3FkgtkfA3JydZ7Oid+KqZaisG4Nv49KmW1DJw5
b91UI7EnNj8PKMvYq1Yvmdc+y8yW2ymgQbe+Xc4thG+GXB7Ppv8Cz4yRB0chnjkW
gYAriVw8PwVUQPluISa4S7ktS88VmzLMN/9PCmWhTcC5gzwRsGCpVqx41AAQFbeY
T+TvQnlDcNboFjMF4T+nYtH9r12bYi/2622IIPngGGQ=
`protect END_PROTECTED
