`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BNxH/1aOpFzNUQIPbElTPYvqUJT8BEqQuLwRmXPDncGfYahZ1dOQPkAybSNyGKKL
NpvSTLGgeDRZ545aSrY2k3zNmTweHwEEKH+g5Pjop/FchztBI2zpjf+AuZInhmqS
YZegGuiK4Iz9BI2/iOJeZSu5+Oz1mGnnLj2NLIsCa3O3uAeH8n01ZVKf9sK3WQeb
xScn8/IsThy69eoOsJN1Dhps6YhxjMvtMDZdHgHaTE7HwJx3NYe4p6mCVqNcntsi
jB7k6SGsgvGeISqhnS6+/kEQBnF2s7iZDuJF1CJkGdDdjowjJl+qS4r93JW4M91y
LX3NhO9gSH86/xHvP9zatM5G6Y3g7kd48ZJpijpvKsZu0vY2GkYae5nuBUS3P8D4
LtjvaEjffJV5DaWRALUuDMfBmm+3qU86dFy1BQNXNKcRktkJ2EgciguZ1AW2o3rx
LsfI8Q1c/zwasz+XNeu0nW8PMwJVND/yuv/NentvqxfmpvL4lu9Tvk1CeQLsSf82
kNZJY0x13u3SFe7XdRWFrPRnzhisedaWb8GQraJTIonA/vr97/cuJglda63My3zZ
qtKIlOyivyvZw3LE9udZZLW5ky5XSt3J9JIUoFpcYtiUYvwY3ml+5yB2RgOEzk45
0Okqf8yq4f8gAGGjbd+2642hVCVr8msuLwN+2+x/f0Qg/SItfjUWmZSaSI5zhWII
kjIGZVtbvelnakHUdsudS5/y5tEDIxEh+dvMNqlr3Kud3f7Q502OntDvKZkHrM21
QcgSCYaH42lvalqo0F5wz+lIM0qxYPFs+m4I4dcvQt2YsWYScvYWUWFIR7rfjNhJ
`protect END_PROTECTED
