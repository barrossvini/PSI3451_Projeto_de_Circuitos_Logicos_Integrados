`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+WqH7MnPd/uqlIZFt+9+SNHCm//LGQlwNyc3E1mcOIuYa8GMUY/CevQjfnEAjN3Q
7CnSugOulQudA5yyPNulyUBBeiIrtqJHwKSYBacsCbjrJTkty52uPKodmo9X+CHP
7IaIR51QSBX8ShsbDG6brfxFkmiq0MQ8saPsBwCdFdlmheleHW8o98gR5LvKsisM
m4jnEdQAjFOLehkbegsnEOK9X9e8OboMkZ78RfxMsdYdn/8OmhEPNadkFo6ThuFf
ekhH35INo6PdYnQYDvvMEPDG6OyXFQfcR4mC1Onak1ipFJbMX9bBQS2ic+vNEc+R
3GT0muGZWScCdHzrvyjLlXGkF+FsAG+LKCyqRSA8wyWfuUvyVngGxV29u6ufj9po
OXAxd5dltP7AqwDirhvIJlp/vhNliGa3jdbDnHvopz7b1f6H1viDLA5J/9et99Sr
h8nWfhycxPUopqGqiJN8l3q21UIWQVUifOm/R2fbxCOe5+plxAAtQrFTur+dkvmc
k5/1o9PhLJupSSYUIi2E25+NqSK3YQ4hzMh75t2TzeIw0ZYzjOfeDqfm3Qn7n4fd
LJj1Ek9FrXodVsVhLXnIBzaeuABfhjDnEzBDyhuwwYiQsknDHO00Ii/h8svl/2rW
Bgfx0XtQD1UuabOktL/Spz6onp2WW6ZzqGs9edn/7fEliB9FJ8Wc5NrD1yfOqvKC
cmRRb9zZghAVvx5lGQlQcbpl25Ry15DV+R8yl5kRVMBjJZecjdRuBOEZWXfjT/vj
AMBZPQszk65T07fHnBYXCFhR+BZPgN+4Ca+dznQQdPtM4f/nbi2iMrssfepk7LMr
Dd/2pzE5VfizMiGA0FlqDxHGF2AiPYCkEEufi5ruwHQavRySobQJEZRPQ0oyiBl8
d1x77NxtG4zVH3TvVnCqIpaYRj7CWRi1nlkkptylzL5XC1XNifwo0YLI+JyjgF1k
yrw4B1NZieEOu+1qyRMPdRt1QYtZ6Sqjxy4yeFNpv4HwYz0O37F1CwKlFhzfXg03
FYfyDEcCZlBZen1INLUSqSJzaIx5zu8AFTBo3ajkwQzwVuxWhisWcN4h1fJNAYlr
6AUmiKUaexr8azoUKMp9ONhBG8tH23U7Df9LceHQInJK+MQWeMaYq+qM9U+/ftXS
d0HkaYb5QCHMhSzMaFrY7Qqy3uefRLEB035zQGhNG8HPr3ZPji0zK4Lf0d+pQ5xe
/tYBXzWyRgq9+ndW1ApmoB/DLo8iFYptpVnL6VrY5G4Wu5rjpHcfHnUOYjmqnLVR
/p7llqhs6nFEAEHmQh/7bY8Z8ixq/XRbOxLQ3v/MR4SukUNP0wWDjC4HDD1M9BTM
T4IkuQNweXSYTxmVr5ao041uJ0u/MGFnlKjxJEHpgE2mWmJh+Vb35NAwcydl3co8
H4kPoGXTRtpdc1aGNgFm319OQ7oCtvHkWNsQbJwh+HEbaHjSBJZeT2oq3hH8+C1d
c00r8wTG1B2lzCaggyUOGp5m7baRc8VwhjjgOF+xCmbCmTj0JXCHCskumLcwSNY6
xpAdU4RXlngMHeqRE+bR7sD0RzxsVTq0z2F3zHvLO8EBCzH6nAbyU52OIvKqdSN9
53Fm18p6j/a4X+YfbEhORzEMJMtrLkMa73hhyR1/DX77ZssZm5m71UCvtASg6yA1
zz/80sI8tlpveonsYg1NqSqd9SuGHUeuEEOKbIUEJCG6BS+DDoMY5YOoYoUeP0kI
UFF6HGsIMubRC+8EYlX9ehiIP1+2gf1sh7Uo4IQnJ+yN08/o2s5Zm0IDOLY8Wb5q
40u4w4tyBsJpDHEcoEV6FFMNgGueDzFT8YHjihDgRikoEpf9hQmsXBi3dABeK35m
7o8Aj/SQO6kQAWvJEgIuJWvqxoGvAMkfumr/mdNfN2fSZpsGPvjvzjbhUngjLlac
mDZtjmDJtULiFCPvQ2QqRDOPIZA+NAT+51IUgrKI3B2l3vToq0fOrsbX4+VC/GhH
YSxEAXa2xHa0FHnadDQCytejfAtquptCgRGIMz0lD1Gx1R8yZu5ei8N2hQ0JIYPk
gfn+Dlc80i6S7CL1FLl2Wroa056z8b+wIo1ufHL56H5NxnokmId97ty8o51OO5HQ
94q7Op7IWIblLVbq9nueZNUhJE9I1F1/uceAzxg43K7QlEo30jqpMI99dUPdyskZ
yhoT+eykw1euLihsSvczqmbLL3bb8J+BzTVqGNNKITBjkalVO2wz0npyhsO0owtZ
L8BcKZUjdJg28/PvOzLluTUMbDxRpm7mQjavpgzat+FQYS9a/vLltKqQpQYdaT1s
ExtEl1Cj9oLllWmc69xIZKAIkwzKm52yiIPATXlkPYofNVxIiFTMzf9gENVUwsko
yl0vQ6V37TgeIObfMoA1lpgr8Agtai0ExatPVdGHVVTpTCPfzcj3+4SgRiz1LgEY
0yIHv844+Zm9AYbzKNABHaM+3brLVV6CzrCjiBf4J1jACudda4DutTtqWdlquJIi
bIWTnHdaTOLI9lD4X/srmQfWn2hPGi7phqtxffwhyYnyLHqlGEACRVkxbFDO63Kl
FxNWfV5gmodDOXFL8EM0dzS+r8sskzNp4i8gwbZ0ooAh0D97w24bHbG2nWw9DeZt
IcyosbjnTtgRFsaAj2z1RrZLxGMfkBG++VKjKKSwU9gJKqLM8C4U5NwgFnMVTV83
+0APWVXdRGLIlqJCvq6sgvyD6X2rHpfBZwan0h9/qpiGr4E2X4D1pCNk1UdrA+NO
ymZUEtO6d81CkR4nWshPwZ3s/K++5WqZekSkXfO+HEpu+fh6HPrjxwkpWHduVGr6
rR5jryKR0hm8ia19Q2FT15lY6h707BhKW7fD5sn2DKsyxPT9ozlKDPnRxzNbQwx0
3SLn8hsYSAKY6HbQvspzMp9x+4XWKjSUdsIPRVPfpd8ycgYnHgU/uetEletwSafj
NjJqj4KLIr75UnBbMfC+xmMgrQFWoF4y2OCpotOsKYvp/d9byN9PHNCFOaTwxp/P
WjvLQ6cI3E8DsQaYHbFJ8WQVM5xJJ0Ow2EKaHZLwEtauyGFCWaI8bNdrI7uPCMiC
eOe/3qd1oCSElpoS09HR5Q08rWekUOv6Cw0945ibzi6PNQvTk6mKGPBNrPtIEyyf
k2zoKx6FT3pXF3bq3gmDGLhhpMR0YZ+aXsai4GkSjtQrOkSOVw0ctrJv6l8jAXfG
CknJtwvM1xsKbFz5lzIFW3E1p0AsFZzMAEdpGghDksDxjMRko5I+gArx+6TNr5jG
wOai69sJqRZwPecRrV3zoZVhLv0yvSGvyOOpu5geOQBAR/sXYjfAp8joJ2fSY+bj
nWs6NYS78GIH30tuzBD2FTri5H4QoS9LhjWBL+wlhv6zmhkK73yP8Zn384UbStA/
Fo5NyUAywBkJ0HBW3TrXDOqlcSqtqW0O94xztRxOqqKAD40RFfaupXTTf56wWozK
3CvTctjTrk+dfi5kF/wkrmrrBgtkbITrUs8N9yGCEzG7gmlOyN2WCTjYry6+HHzV
AXSpRYCpfqAeGJj1VOixbZAYa1nO0ikuw/DS6dnOdUWgSdDmIgxfT/Bz+7w2vEvy
I+Ly0TKFZ1r1ua01El3gXqNG+ELTxhAo9LpJcP1ZAttovFrrFp6u4kuuvkR0hZ+J
cE1yTINJY0/QwVI+bUCjodc+GqsK8p5Vd9iK8A/EGzqxn/1oP6IWh8vZCEJyyGy7
aK8K19lZadPnL66aGJyLKVN2sOBzY1PASNI61zofJTin0YzevFVD7rKrFFfDXpdQ
0vhaHymyxgCorn97eZg6Xu5SqN1bh0wEyom384ulWIsnZstnuW6l202BQYmoi1AP
0ZrdpO7pRUmC6y/QxgJiGQ2/Lh3qRBh5ZXhEQXvpzXj72o7zq9PYf2qOVLCdCp+l
myIeo0R+WWYi3Tpx6oqbLgrvh8RTXgU0ZjHjvqD+FisXbLbX9sZvK7/fTy/fzHgo
/djt65LkdbbUV+hpoHFIpDOpemgKmGkKqmKnO3XQ71hS6zvbk5T+HArQnMZ5uZeb
NuX9wm0bBEthCJNeifJ46AeTUjl58esttNRL/rXGJYLSBLBxAI5UdGTnXmRMJA0K
D8IJ+/GXtQa91077eYl+AuyjdjBbDzgdNyA2KHS46Ox2yBIOGkfISwFAzLBVyR+A
6hZUrS2qFoeW3XhgBHzSGtF0Scbce0zr8ogUMEswxIC+jfV4cwqHelK3/GWitQcF
+KfUa6W86RWBMDP8CPlJMKuHEZEyg//rEJIITIQ+MUZ+3SqCOTLrKMVNmZvCasym
ZDNGQaIZGMYJx9pW1k/86bIywy2XLC19nR+32REkFPP8CGRKn/qBWn4hYoJByz+G
jyvSqb9u/xnuZFzqmE1R1BiWFgemg7vuiJR8enyy62sum9oXSlwcKmkfuRPJOB1V
k6jrtD8nCrKCWp8FvmxiJiCc3gwqHoUotbf6Xa6Z1FG0rOZGxcClCx8lAu66ODG5
Mv3coPasjIeQzL027oQL5f5cE4AbdS/+Mv48EdexSZ9bMOP3H/3iv06RGd67LKYv
K66Nsj+XwOtiSd4dfBwg3/RsbvIWMExZoTYgoz0xy2Ozc7l4J6Hqru7rz+exIWmw
aiMqw4vo4nBF2QzJkg8UICizDVfRqPd4zQDTHZgl+YJ0KfJ7QsfTSbiTTnUlfQdp
vh1VhWbvhBw8trDuF07vEMAZWI+9T5/xiIb3Rf9M9MfOcNkbvZJzoTYzTqY3nFZh
CQkmgKez5ITPZmA93maRqcFCwCq8f1KtwtjtFMk0WU4VvpPonLhn8+TqBu6WNKwV
qcEA5N/zM3JpLrZZV0VFN4hS8TIhbuiJTHb46fCoMPf9h21aIkVjBYqJfVa+qgvK
zTvjvB+3a0Xyrq3ByM6a5YnwKzYqq2ektOtYuHKXM2jmbv4QAF/GsBg/ky+96MPm
fn0e9lYTTtWLtcX8xAdB6Y0AM44bVtnpmNIDAzz5y9Cs+dnS2c5zbDMIfsQp1BtR
azrNoRYyJEtaDZH7EasFRnIt8+X0JN64IjUcs0Ps7nHpRDfQx51vun1awVQFJVte
o/AuXh3SVwTAwMuD5L/pSHXGwwDjgjnKPqHK+t8qA46tkSq7pCuOC54153fyyN4V
pdd4urwPH9+/OxAQIlnwOl509vRGn/9uO8sThBDVdSibwhVMkLr7mwD5gTu/rpWc
Gh+bEwFvaaQwZjDlxA2rbtCw9TS+PIY6EVAhhQu03PzOnpzTve3mZewuylaYFkuK
CDGkdsdKXLrEM1NzeXD2cLW4GKr9oCDOH6PC1yJotA2paS7mL3sUzrd1BX2Oblws
jf8KkwvYrxlFXRtR2+KKM0DHJiBKKccuAPF9XXzhjCOzmkEQ7kjysfn+stm3+lJj
l/djO+9DnR8vqgbl/Ay8zD4IWFRoR3IdM+nb4ugpbPA2rEdl9xDvKQcK/3R5RN9M
4m5P7r8qu6PZ9xDF/jvuChey9RNzv+z6jFrQHwXREmykbyFUcMZ232z+4EQmKG3R
tjyq+fTybT4/56PfHdjr+YMeYvPSc8xxUSqIjAM1lXTensbiR+ydMhTNUlR+DWNQ
9yJmv6nxKEIwYfXwGse2qxCVI+Ze7T3qRoE4tY6OWtzpTLT6kLs4bX9DYiDOP5++
WQk2MCaLgzdv3aFYQHQSYqPu+3omtwmp78m+/d4pQnS5TRyMcAZsfZV0B94kQ9eV
ggN3A1Mp0ki9cQSk+CDUeHrteSkloFAOdaWd1PWWoQqKrMTKOFrhEiRIZcvWZYPL
AvXX8kekWcESRICvZtYf9yzGZp9mnx6zPJEqh3B204SwtlcV4iBlKMyJvqcrNhLw
Al2SeqJ2cGD3r5Qbr5Vdx1rK0ZM9JH5dULS2i6KWZa5fZs0hiAFiVy2n9jgI2jad
wrhMBMnxwImEWyXRIR6nYALPZg/KZAs2EOMx6DuAyc1mP+ia4+hFqXlpOr5RelTJ
ew0UvVYXuUh+dJLFkdRqymz1oqqCXJ1SKcAuSLiliUSoUyZxJCKFuThTATgxROt1
wdpK6sM+2Q4eoo0nBzNWh27Qg498nFEUEJ/nfi9i/IttSCTj4bVTq6A1DZOVmLrm
0oVn510uXLNcgagdm7DUYQ8qLjc9FWQTOs2042Al9UD8PB9utXJAFF/d1PYWou3Q
MZBd71CXL2fS+WYLhZgsvGA0gJ5ayOq2cdFvEDZzDjjeS7QhyVfuwMw2ZArhMGaN
m7v2jljQ3GXWuK7faVDLxkQOSHYxzidslSRAkqi1HIYJbM9FwjwUZrShP1YyvQSg
F4gq514axNtwJmYCpdm24Gux0MwN6stZkT6vclcyQwxRyTAmWFzJ3t0LOsGzOH1E
lwaeAhRiDnVkquCGnkLC95y1+2uVOktAxdyW6aalN9CePm8Fda4QVV7zXPbMVlHQ
VQpgdQTIhWHCSsc+am02uTORxTqDkftUVl5kGM7ODIlkcNJ0+r2M4Gp30jIjv3/I
on5LjD/LtrGj/SMYVqlE59qEeSJK75PYQwgnfUH1g++xCP+CZbYCK+Q+KfLW3hKG
HlC54M74Ohpv8CKBDawzJ0GFJYCEUzASxtq3LOTTIl0cgdz4193FiWY4gyu66aVr
FNuYZU78AIfhRa7IXA9QxBI2pDSmwraZDZ+cwtyAti+UQNRA5jceVs8KG5ZoPJlI
bMudMF1/2l/VSvfXgQ3ZqluvY2htUoxrV0CXLcTAAeTBq/+Wy7kLy1qtZlfIw6F1
jUUaiJUgVoUfnTzS3ehCs6LK4cSMKfvEt/0WauXJPOYK6P9d+e9b4OTCYmRPygbT
uf8dIb2zpbAWKnzOm4UJXYWOz5yIc2zIg7EEFYvPGSPSGBO8QiP0eD0MwQtpDO19
NkWu/zo3VDa3gM07XqwXp0Aq2IVXSd6c7UU4OgDe9pi6l6j5P9FiUO/P1az5QKm9
3Zn7BOyydIk1/6P9f0/6PiEPSq5pIBnbD3tD2IhCheK34UFTYlkaboEKVEyf3zDH
OxDf4ibipPMtoTiCuP63wtUJ7DeeLLHPKpBAsBcphkOTTxhwcxdDQo8uwG/niQVs
flEI/RHJXI0hwsLhbYJqjMNs20v3VhuCvCVap5d/bRSHi6KQOkoCAOWhOWKyUn38
xFis7nE4AEpJZKKbkOGvypj1FPetEudkmunvoriUWNmvrZLcmGWro/3Moy1yusnp
H/mGDiE5kVWI9iS0DxK9O8Klxrbn2QxrqGUfSEW/u6YEVMTmjR2uv5GtCSsB2w4+
nhNGAwVD74B6agyd98r/dJKGoQ/kFNHECUx/GHvNdN2C1SPVfEokbrEWC09BDOO+
FMssEl/dqM636xrhZYke1liRWt6cn8+AKxW+VMcElhTDstv1FGOR92aTdtTUabRO
LMZBzGv0nbP+KiyK3Qg1nGedUjhWwWs7QKPTHynGyxrdzuIQ5Ese7J+zqh5V6gdA
jlEdFPZqYqkNhTWQNRNA0bkpFT/mh7iMLtrZgZelk3VealQsmSeLyuDW2zE2LVKf
ZMkan3ugie/9XoGSWVdKEznqo09InY1BV/lxwyDuWvTi+A9E5+0HzX/akrGBCgUN
o3G7TalKjpOpL4v3UGeVRZ5HfLpshYDtLor/23G2UNO2dmz+NB8sbEtHJrE1ofYp
uVrWwOqK7ztAa4nee06laB+lZFy2C+Hi9gI2adrJMlZKcHO7bpn+cqyfZ14HIv5p
7Y1ugGRyHp44RC6/WlPFs0PN+u0E02edAhb51s3I/SwNg/PCeHhBKqVFdijP619V
dNKyTgBRc9rwAhvzvWzcrM5gdmAoyq0wGMSeaZD4lYxdzUE1V5fZ3afjq34vdBhs
jkCtKFKcvqZ8ReArao2kNbfS8bS3UndUrh8smnYUbsH9POvjc6GKgOQTGECwVFuD
Ma3huoz8a9lqHfkilYOFBfg97z4xlc79ep12hSH5FlX7jatqYA821MO3mIMmXaWG
u74vqxW054UPLAtdHTx4xBvzejsDmHIy1Bk3seUhCWjzyUZepbJ2yjErIHsv1KRr
657ZvOvoIV3pO2c+jP0BlHg7OB8/gvWSo44lJHuYbQrboeXd4Zty/Gy8CgD5+5kB
e0vGFLhm0nzpZQ/4xNm4eWGy6TfUu1e36xvRXa1l/2UlXnH5G6AR2ifdvBq9Ngz7
t5Q8HjaKyDKTsuHsgYgMHIG0b6RhpAULxk93uW463Etw1meMca70UKrd09fndM2k
wDErgM85tKpajUHN+qNiK25napTiwy7k0XQAhxkLk483/NG0DtVxNcLXbB9kZdwi
rUtJnJGKfNZpUaz7FlBEv35Gwu0lm09gtnKXzJDFNTylhS7sANLIiVFeY82QRNrh
Ltqkon+H5tY3Igjh51YCXqYIH92MyE67G1ZFTpwEenUkjJDdHsjWFJehY7uW0LlN
/lcdyMObWraeWrJbum3stP2xiqvFlvpkIWp5CAqjtShj1uUshBbw1Qy926FXlAcK
kthDATrMI8E0hoNNqxmgxj4kA9PJWyA0qTLkcCg3B2AbYTpwTaOGB5GohJhJCBvV
uOpdKl4v0o00v7HL1E2Sw7gQkgALIWNL/+/iEkgNYO3ZyMEKDBXPHfHnrXFkD6Fj
GiOTB81+EPT1hVUY0S10ryyBrCMFFc/g1D4mLdx8Mj0r1peqTqthmifD14wOBdsp
M7wuYSDcPlV/xH++3ZIzxF7qX28J4/Oe16ADiIMhyNAqL8PUPkUclFOSesopsd2u
WKoIRkDV/bZ+gfTo9OlXkQiQjHMUM1I30hd4jMicnJzIP+6x+qbykcxP+zFvkGV1
mpANkR92/vz8a/B/0Ml6fjeUHfvWgfBfywk95q4NzgebGdArv2dmWqkjy6DsUCRk
MjwQYXbuj9CmspUmiiqTYTkB8JPcoBFx4cv6kXwohG8o8sJvTTu2Zf4svFU7hoX2
jbqTcVe8TPl1HpkM0g88+6J9+Z2f/ULFm78pL6BzdRMIsQw/FFk3cM4ssx10RBX9
5j0AoL/bKKRTuwPS4/4c9DkkCwclwneqTt/hjA6RJBfnJqjoJ9Ko5+1kUYWxQDv+
P1QOZ0INbTuvjGaOJ4smi/jf3UZ9BA4o4i/EMIwg5gxHjsAivE2H+mQh8Dd1PTTI
7MpfF/WaJdelZDBwSlrMlc9cJT0B8nt6wGLFs/Mql23tmr+z1mPhKVgFoO9/SBU9
tmCUT7OXnBgmhCfvFGq8Y4p5cPOngp4CgaS97ZlW3snTVniFBOaJA3JeWCJuEShp
NmjpOSvQ4hCOMNXIz9A9K/VFU2IAJVtacUPahW8Bkcsp8/2FafIBa5AMufX/M+I0
iSypMfghEUK3bapT1BrfTLRpMURNlzjbDBO43lXUOWNybrh5gzh92W2J0Zf4EvZr
pHOfgzqA58yfk9K9eSJ9026v0MHs5yo/H7t8f6RHPqaIyscEO0sLiWHD2qn+uR46
j7xlSJK81YW+1kyfG4OD/OZV0sN2r5+oZdupAkZwTUQmyZL8gpsNw7LNgy7qtV8z
ElE2NDk/spmLC3k//iCLn1/ZJnvZFNDY8UM5KzoNtDE/mqelE4uViJxnH8/56cyg
+V5D9h35FNTQRN7cE/coIfBL53CxGhBMzXMKH6K3XC6FMl+yjr5m/TBWRxmAhlv7
RCWaAxvBT8/pMWbuKllTjz5o2QKHPSsoldeGl4xlLeN5dNAf3HCLnnkNreS1IAEk
HPkEOXB2Doz7g1cmKwWYCMAUaGZEILxnYDziRYCd5b68NwkZff0whptB82l70eq5
UdOLc27xUi9VxfFxOetM0cJgbFdbv1PMWI8FcQFtgIMw+OXIL25zt2bgJXkDGyoF
uSO4heGrEycBLgDkQp5Hzxy+kuYbqUtdtJcNM5AVEmZ/BRYFo8YYdSGoBQEaONla
1anBPMEq1ls3gPhSHcJQ6fj0LzYI5tzyAVnq8n/kOYsF1k9on2V2uX56GyCvfRiT
uB0k5t6DsdNE+21N78KTYel6Bze2q8QpbIaeBkeFgjlenXeRLku+rSDpkjDXRhFF
shY1+/agR3RLgXibpbM6Qzc/wLBxbgBHup5trgbi9NrRODB0qFEtafNWoi+L0I0u
FJDlwUgoV6z0WLo/gPeW6lnFlPop1/zJYsjjP5Ie7wb9RiUUULH4sZBEa02BsaqW
eeuu5k/oey0dP23O4CnVDqKFP0JsBOrEHKpTKYTo9WYDHWf5wcT/bb9kVFGwiLNi
E0xJomi5LXjYeA1ehmzAjWQPSpyZxGM6Y5318eWv2NJtpvPu2d91sCHE337bQRwE
GxD1GFIVC4ss+6ve+HusJmnALesjx41C/nOhzf30fv9hkMbTnmeL7DODOAb4ZGoM
ieaeCdIpudUYG/xZJTFKy7VWU+ft6gRKtN/T1nPTNvPuWZaSIAlrY5ylhb/Gfkx2
Yi+oQMG+7QhNOCWwdm77mZJ9cD8nranbyYFQe4vxeB6fZkAAcyWNiZy4GMfmSdS8
W9PMIixytF69DL7iZ5Cvd1NO8q9Bfc8T0ECXXmjk19OzFiMSacZCA/jBJ/5UKalX
XQPM6/qyMvMnFWuz9Fm38jraKswTr+l7MYwlBf1M25blxtt6pnRZehXEGf6Gukwi
Cs+GWtVEmAgZCKKWYzefqmRuDtI55Ac0NjLKwj9BwOGl/bCUjP3ijJcpf9XydgP9
yA9BBJMT2fMqgt4+pKVUMcMZ6zDHOGb8879tNnZZKarR++8V1mzVHVNnn2zCUtI0
JbyN+TaiSeMySvgrLH1YhfNPRMcfEgXfN7NHJtKq/QjuaOnFCZiR+qyfN3lMlb5F
0CW6DT7ghfAOlnwOHEDoDJU/J9NZL6CpNsfZClSN0OC5eGiLz5LuQ5xl9IMb4Owc
J+lJCr/80mox0TAf1L/tLsOKCD7XtpRvXta1soXsbvSOQ9dhxifdDefjvdYSAQOf
Gk7u/kRkhQvbdmFznvp0dYiulFgqeJbxrR5cSX0Kl9qhzLUz16AiTEzUGWvEZrij
7xlpM9iLBdX/tJix3l8HDaYJ/8aGJ/PDayn8qXgtCsPhXWsJ7K7N9jBllmu6PqqU
k6R2Rn1xNg19+bQ0wd7L1YRLfRTfce/+Stp6VFmHoh7SN2idfql4XFQlDWeT8xxu
beWoSK3RvED3u9ToijsnBvpcS+2PkGqIOxhtuV8KkAKss2Kfveqth+5a/+PIxUIT
kEVifk8VEAfpnE0TBumK1EmVKYicz8qws2yfS3DBUm2Crlm1j83a3GWibziKcQTW
+wvXxrfsAa6bXlgXpBWkZFAZYryKrHYij3opkzlFRx9QoAMYlX62Subo8rDegcrY
tZyE1saP2L2d13SoDiyGGbiGs22SJeFYEIWJw3/kj0i3xo4IFn1/mdVUj/TNkc6T
afHS/NwQXQNvbPN8f4Sh9gQuzsvaJ6KT9h0Mx4TNTO4GQKyIFT4E0Kz8vx27+lBu
uoWcj6RUAvozT2aLqjxZ3HLIdWHUmOJJCc4ys0Yq4a/vuNtu60R1F7aqSFkKaH8d
3yDpNVw/ODUSoHeeahuHKLLij+JPVTRp4diXhKs04tcjjMbLMjPFKr8OxOJw+lZv
/k2WCx+W9ZgJgwe4xuYg1knUDlfNdfmwnqwRoWD7f7kaE+o3DWm3JVw7apqINRU0
xD2h/8mK8Li6nFjwq5bWSFMZNq/Vz8KTvSAn+dGawyCbpkmQDQkFgJiByu82tprQ
GqW5aOiVIlKTID9Vug4gVAwM8ixfp3sRR0/NG0G8EemIBsX4uIoU0DJ1tTMVNdmP
TSYjczMEHvfZg6+ygg5rS6JPI947ejcoDoWbAdxQHjPdm6HrfLsUKpvBZJSe1Rco
0tAtFpLPKNIhl243NFRuH9SmIBjqIC9sdmSvU4Q9Yyi9PGZ7ElFwWFrOwjF/AsoO
2F7xs6knk39DYMvnd0yZwUCdBRvCqrzBLDk2kRSbIVdrRsb1xJqYGalSp8DUCnZg
Eaj9rbyLO4xJ2r2DFZrP1WShcfYQYWXHYegNE6wfUBWaa9hc4HZMZqTWnK9WoTgF
5b40G3GLkQTUNITbG7wX6qQr72fuOQpqNC9cNz+kJxN3UIz5xtr3r6406caCRMll
tFv5hOPrnJLDansy/ySkcA/SW02nooP0Lkv7ytB8LcrMOScpCYN3NSZaD66mig9k
y0l5mcNB2zYGfmacQjdGR3YcpeaQt9lDMCCVi6eXueAj75VLLKKKqBXJIxMigCjY
DkeeP+8x9yHhZgH99xi8/fq79WUtxd+Ef32B2Ub7pkByrFequ/i2glIw1T5A6bvS
f1vqruKxfk9ayjkzJlz+FqkgSlL0s7tRK8G1rgvd8Y/m1sGtcMoRMaFY9+WmI6Ch
3A7Jpw01HE2BvHqfRnL1yyqvbyh9fdpU9SMWpQF1Dq2WAuchvl7SsND62dhVHhRD
Jy4dSTHPbINT50mOBoWsatUs1fdGF9uPtfWgu0OowKxPJR2UzWZFADMIO9MVWeMz
c/o25a7WMtN0uQ/Pr48IqXDBHadLOyoS20EM4K4E9zGklkAsBm7MK1wXE83HF5ts
aMYJazZSV3QV7xaFLiOBjPoXHnVExBdsNrsy9SgnZc7wrry+s1tu/299GKBdNite
KVdC3gQd4fLEqvAGt85azfDW8sLw/GNnuVXs9yUiuWYM42YJiFsOqXoEWg2t3wES
nIEkqvhB0zQ3mnQEl0G52c7sYR0mRRh2LnOKl4EG5/fzmnsWFNBOz9TREnMrVrMH
MuhHr9Wp1jrYyOoxi9b0bjJz79L/GyHqv7KZsSdA46uXT9D0BA74DXw4pTzLX3mh
uBZfF6NwORJOtQ4uCoq/U5/zQ9bsSN1lhny60qP3qnjIzQV4jLkhkSA6XNU2J4gH
GACEULz3Wl9z51VofiBvEUKeyaTIp6POxXelzWhQ2O+T/NAQXKwcTeGwmCIXr5GH
XroEAoyhE8rO3Qgm9uJzKnjHtOOxxNxhUbnT/ZFdOHH/u/2XO/rPILR9LEAR38WD
dzVFJfAGAnsdR95KQygfEplUJCMQF46CTz/1tqOxmsTXogVTLtNk9y/FWM6n4rLa
dStU28BK/nKkkDUBG7s8+SHeXfHfPV7BpOGijtWnl+pzeu9eVM68RtDcn1N9DWWk
MZkNCW9/JVqVOTP+FJs9LwpHmL3M7ks97hesXJaZtJhIPzmoBptZGy+cPz8gmg05
7/gAQxa5gFDE5PXtFKwj03N6lQwOO2cKrxqiBefud8OmWCwx1zblc0TN6TETg+Kp
pmbV/FaEwSwrPoyUJ3Q7nudDYZBO/mK3QtDvn5u5kC6FigT5uizy2xF5zwBzR3We
PD4vp3LNbpF51SABHh3G0h9tZfvEsCEAy5WDHNVJ1U40Tz+dCkoeDDOVtJJzpG9a
cJWDEej5zq6KZLzGl3+5TxnsPIzeEoB7waeIE2raB9Po3iF0cwzUlz03iyZ3Myjb
OfWAXE0rUp7oEiZVOKCHFvlRYoQRA4AZpImyVtXzo3EBi2w8i4psaVIrYWuvaqMD
QeicYlnJCSS6Wqta6w7z5yN3T4xUen+mEiyRgg0qJvjbzkxpu11uPio4/NUc5gji
MeUu3JXnhvu16H06drFlU2rCbBiWARDc/ljmxNiDg5vLkiww9GFY9J8jCRltZ53p
yppRUQjvAvKU06ISQBx+aX4rRkJVdO45wsqE3cJ7qhUbrLGWakx+L9bBX2R0Tf6K
0nOiBzXvdgauNm4zbM2/rsFcsWzDMxLQGfFvz2PBohMFC56Gf7p10lxo4HElWDMY
NYCwIqlH65BbGHL4LP5bnpJ5MQxbqiZTcX81R9lcd0fxiafpdIeNUccjWpIiXldE
vydpYtSqFQWW4SNtxEQ+jEgi+KdMECU+eJQ3Q+m0DP+oz/2p+tH3sC8tKzXPCPAm
iHG4D+yh5GFC19ZkFjJmc6mM3xlhQvTCtyv2T6ELn7EUWorTnckVd6qzyguj882I
6ZxYN85cq4F/kyptUGLDt8Qb6DohR9G3XJ5lTCwxXv+Yk7MXBVI3urD0h51oiY9j
JXfXn2ETOFjzP4doC9aJ75D0BhHseuEMXY55JqLCUNrwsR8nlFW7qyohU/1MGy5N
K56L5r+mcBlCzbmU576bs02ffwSixN/i/yMheOttmvox7C3VavBRlniVW9tGMNLn
9iw0ra+/ftddE/ia7nEkFMBaVznGnWAD9OoWGLOXslLCduCgRqF68f4mXDHqnGQV
v7lgHZnWsep+Zrc5FNYdcdKvr//locYiK15ac/KfWxcN3/4RrBQBih6h3Ik/qkX+
nzJrlWyNwtpZN9EhyzQZUQrHtTxy16o3ZKNKwOPI28irlQF0EjzdUXUXQbZJk1to
qNIbaTDH5/Ag/cz7WfjXUVu6B6zepGHzNWLU6jFiLt31Qhm9BYy06ti8s56bn4o9
IdQj5aIIxUaDx9bqf3W9LUPJSg/7L3Siqq1iZNkSjbvAdOCa0ro9XTdotzBtSVI2
KHF1/M6E7t2tcX6LQtSnHlEfrAMGGvJcT2pvRnaXG0k7zFr2ZR8qIlnXTm5BVibb
2je2IqBQ8xMEjqJcy/XaBO64Ybw2JasLHmaH1O8j+vRfAZ4p6Ua1q6WoL+zWfGHz
ZhlCCMySm+Y6drx4S/pGi3WLtlNRwvrE/4/ILZ26hJF14vE2HaNW+TkMq3Sn5Ikl
zuPpdx2NsgcQyfaa3gMul5Remc77OtOLEeM7jKDx8yvVZBmnHygfJrSvUAZKPdy4
mVQI8EMahffLZqDonSRL3FlN1UixtwyL5ArxiSfGdCx37AZYe/v4WJan+y3kYNjE
mStNzmTnQrxmisv4YXBvsXFNoo5/wEcM7O1v3V/18YvH3DPm4Zk0vjaDD8o4a7FT
vOJP+7ww2K6Xwzktv5zJi/9habMiTkwVlpyu9xK0VwF+iMw7VMQ1cuSf+Dvwx29K
cr1N1BDEu1P60sCt3GFVqaWSFVLUlppi+o3jup75SZMEzEZTbShqZW/up1HWXYo1
mE4+rW2St23g3O/KYfBIZf32/ASwIx2thhb5L7OCqlHPuddA91jqPzvHva6MdTMG
sUhaoaLuzQ0+EuACRVozu/GgEh8sD0fYCMwb7aOt00mmVkcKtiPmd3GbBr0hJaPL
XtAtCsAd7Ggw3O3fQywna9tPzXf7oQXXgFAN8sg1tZshr8Q9PhpldBaJH/6Sb534
0H7PFsUg+SxCOU5lLoRG/3oaRF0kgkeXpoaOjSSa19hLUeCXaMNxZJVvvEPpXt2n
JLgW0BNyVY7UpjP4Hj6+5mW0db0ntkyBUUoNfNU3xW3smsP/AprhX/c0yPQXGEf8
QcSdVwLaBMIncadYqH+EKz3WSV5JsucNQduri7xLPjwdYtDCI7RupRZMU1xaAmLk
O2tT+/R78f7iG9QFoEoag6ioJUXABYXpeRK3Q+fnOvPdJUDrjHm5oOsJ+xA/C26r
VrrXr9qQ4ejQUGXXQNCt0q8uZ6bF45vbdz/p675eP1xuufqSnEbXcwrL8xeuBOxZ
aj4eDs+MEzFOWOI4P4/5GIjucWRk3WRkj1Pt77rh3RdpsD2xeutei/YgVJ8cKx59
0H7akLLjhq58XjYvA5zyE1DJgX4u/30L1cJ1N8qUQpqGbVoECVfjfo21HXARgzFY
Jj37SZsBod0T1PviwgtyNlTDxgeMJTIGxigsFmznwXMg+/qwo0mS7IswdeXmEcDg
ZlCJOeuWvpa+/8/OiJhnAfrwnOoYiwgwlw5IWkHcBVhlo1UgFEy+jxkTc0Vjhudr
nurGWEsh9uyQxUNrX1cso/oMspHobT51DHyl11yolhE=
`protect END_PROTECTED
