`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SL+g/q0F5dU10qmRFF9gHhzE/K4UEpmZ0X85K8HF0NMZFUvlS9ohfgnWexahcJUl
oiMfirJ90SotiWNv/1jUS1Fl6RQgCK+48FOTnOJcBnoi/bJ/pCXqqOUXKxz+UqBO
u+GCLNSCFAqPQsCKQQ1ANkqm96P8BOa/ie960PDYKiD69fQvwX5fCulPZ4LMZHBS
QlA7nHEK9heP0vrvALyuGhu+Ulg5ND823aQDJVwaSU1wkVg6zXT6NjJZ5OedEt0b
rAplpiZGFfDcgbKRgr8A1RFawlvPqEpYe6rOpe6n8XwtCxM2u0AdvC7zi6TKitDI
3JsOBFdeIKfM9f3oeElTqq6QVmbG6i+Y9zTYLMMZZYOJWbcibHb58ooejbUgXCP8
ZV/rxg5kfYYpxZASF9K740W6q5UPQM3cuXHtxZZTkbYCQ7Radh0zP/12DBFTz/97
Zfiza/KSJdiRbQVg9zlTGlFmDhgzOZXmINbiQncVgVOsufBMptmEseWl8WzoUgZj
bVd9vX5FkbYmZbe/7TdlUKPd7fqt9ba2eW7Hy5k/JFanSRsQxW6HG5rzmqq8uJhR
BSNmcxhF049Fr8O0oK17feqfjwI+Zv0i+40v57KkdgXYxoEFh1+u4nUBhx337Bvw
Kwub40Rr5u8mvVmOll/9Et8cLFjsh/6cVyXSRr879NwSck728vicsFaClJ9HDVsO
2Jn8nMb62qC3g9CbVfViJNUbr4V+VqvtgHNkisyPZi4=
`protect END_PROTECTED
