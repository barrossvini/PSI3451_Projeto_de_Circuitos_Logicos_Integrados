`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EE9xLjDSPzSUgq8MoX6QgSRsCuVZ3SdZjJqUJaBnnRR87gdyGlpTqJI9TsBQXlQ+
LVjbJXdtsve5RV/wQEUSdfwgzuvdkqzQK36jZs+1PW58f8X6RpH7NCGxkLmXwzv8
S+OqAowQ4oQt7fgRgmCXlNqe72SxczT9LfwhoLgquK80kkQm364ECXjlLH4WbQNe
gBh2Vvy/UnqR26MdO+m2vQpx/j31ZQQ++NsGfowUej5f9xYH7wsJhTcmKzSzn8bk
+WdWHfjQqbJPSYhyw0YXlSEwO3FlxLMafxqeg61meaPq/ZM4RyE6tGfUQuz78zD3
nVsjnFdDO18MFdapTUyAYb2thUjI3+P+U9KF85Gh0RQkC1gOBptse+shPlcyPK5G
GQiU5ZNtUqjqZDecfMXgPVpaEO4izHPLH4bdFKT4v01KsSlfmipzB/dQXW7Umw1H
DD2RRUgtH19x0ctiVTgZtmlFiS9CSKv71arEgJjfOPXZ2rScFk1GYgn0sYGC9A7q
HGSDB9hjSBV1sMamA3qEzi9CyrNW7oijsKjeixphmVLC8Go/r17kySSWK3iPtQdL
QVpKfZEtN7p30z4hMoDC7mUOdKqd+fNq3ZUzsRJg6CFn0QX4Cyo6b4QqJNNghuZA
PGfR7jdoKMc4HWF6dIcrLTbCwjsBSlgkV6jKmBoP0vVeEu2q2iUUBuuZVlMbA2ZP
xT5M7ug6sDaFMFO11aXyzQNtvk2q0fxJOUF+Rmw9yapo+onWy37HLUjZLO88s0AF
luk/jNM71GVF+DJ2IrtAXPZSkuw0TE3B5i6Dp8Y4T49uLxcWrYdZZSU8rMTuvKr/
d2ijGw045xL2KaCu4xOy7zBA7mx6c6WyagBY+oIS5nCCSRhGd9bdPrjKvCn9bQp4
d4xnFJE2L28MMb5qwsJjMs87kYub3l9Gby096Q+LuLimVrmspqamnlpS2zQqmYQa
3lmUbINz+Jz3H9CvLFJYi/W6kPGs+4baoudZxmyAEOgiD78Mhw/LXH5obzosdXA/
ev2BLaWQZhriQie8ooCxLcsKP8V2LMnGVwOUiUteWRMCOfXThJJgS8vtcrm2fJ6b
s3RbeY7ved3nhG57MUA1LH30LMhnc2EesPhSIJ6WBUdwrunXEYyhtNJ58tA478tZ
A7FPFFEEGt0Woku+E/YZf8v/ds6PmsGxGl3AYwKVQt6xw6Dggx8TptEp5OcZ1mne
jEFIiwwdY4qHhDeO2wzy1aw76wbRivWSjWIcJqfwMF1u5+Tw9lvFER8cm1Fc9h9x
9Aaw2hW7HG5xzK9FVwkYs3wkU/9xKSTD4hDqUFMMR0nQCNNg173YHgkBih3T9jdj
A6VB7uZbEqeXVjLcBKDDb27SMNMlbQc5VI8XEthlRDoHD7acnlS6qHETvj8DJpXJ
FsRi27PCAdpT1ypXK5MKGw==
`protect END_PROTECTED
