`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H/HY2eo7Om1lXpJOLQsiqc3idL90586y3cD6fmgeGjXxRdrkJVr45O7rcj0ivTsq
f9TOaJ9dH+qppkSsPp/GRHTjXgXYq8qaF6BZvo2Ehvpusf1lCihSEFQGHRj6mDDy
LcjdrwjN5bMaWLgWq/BjSVCtygMkz/IUHeNX2CEZqRN8qH9rQXNSj3yp3ZQX+NnP
5AMmxS92O51Upapyr7Sk8e3dbqvGShwc5sdatGhbbWht+oIi1bm+L2FRB6/fLaIX
LvzMD+ifBaWvxv00k9tJyPNrYszSXDZEUS/LQ5D5owgtJXIeuTnvlBXBBv6X8WoO
7yEmxcWBKh41QsGENXfK4PtB+bWEQLpC4P53FDoEmzWnoDCbW+zeY1gmMHA3e4OI
NhFmolFIRioVAssUUsZpT4PCuXg6BqC+eHQWu9Ju8eqIGHF04IWmpjAenqDp40ui
pBNsdR3Cd6H2T34e1t84jghw8+46I1qArQtbhZw07xJECcKyDsDY/so0gKxnWfJN
tLFePARfay1L40mh+lgRY95b/NoqgvFDl3Enfn0tZzs5kXoqpkvNmWTSFB2qW2CN
TKDAws3aGYgmaa+0vigP7NZZ5OmcK6Ud3RMvcZ5A78DaDftjjMin1WE3w5gVPwwp
8/uK27BTxX8KZmJu6xkGjesUymAKTKS7xtE4eegfA19nAZCWZcMh8m6yFaAuExyZ
1biYGnDr5+OhL9j12n8vostN30Bs6RsPSjgZ8+BWUYilHkQKYsWd3S57ZTZ76aPc
NkgG5bt4ORTV4oeh/SJW15rZdralLUKtBreeDGzgeaM19nUborzfrFIVhzVINbvg
C/WlIHbKUE3aPddDkuX1A3KzYzhiynW1yodqE7ckm60vVE3EUXyOZhHfdQeNefCx
ggVew9edDYtEpPalEDj53tZUQM5uLCcgAq40ZtBuyeaaXbudnz9fQS7v2ywSR6++
XiSRpQExW1UhB8UTgbWIe9FnGEw91+6hVJMaRgQbjS7ydOI3YPxymxrvzEy1wm26
Ru4Yadi/6SG/zYnlplLxTMD8fOTh1jmqE5aH/q1ZqzBqhqKzg/7+FrDcoMeqsi66
WAQ50QtDq9xY8B34XanSEmmRqrkWwY3NKSZlNJAAWwrmG+5U5vW0Ya9lCI0WTWsj
gFIfXz2Do609NA4SCBOxciBWkefiwMS+oZGMSmMgNy2pgZvCsQ7ZwxpEMTfcc9Jh
jIjIllYP/hqXWVdFnkLiZJrp5SXHfYa2IhmelsbwJcA=
`protect END_PROTECTED
