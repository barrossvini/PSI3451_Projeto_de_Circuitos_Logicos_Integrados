`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FmZTlwdfU3yKjEVb3DpMVvQL2lk8ACVdsAxu1Q22F0YrERCXhhnjJZJTyuU/lPU0
BqZFCzDWUjhqw+zqbxb5nIWPaujRLmFU1gGwKlELEwnSPOgY8dnzUBMRLUXG1ZoW
3ZO3z1DfwfEewaqTecK33xNwZARUGTcxbXcWdkY2Ns56InKS48xHOpTFBXXBw0i4
nFdoSxZ38O8wqwZltFx1V/PB36gMTDEz67LdVe1W8amyMdbsEF2m2vXauvCLm5wK
mJScANawwIp+q7hnyymxOJNijaH+G2CzL01pA9vGn1iVbjsG2kTsnazmzfYoA88j
AYF5ZJ/A68KIlyJdKoJpFIKp0xGi7TUt8UmrrBawqBT1AErgen3GrHtTME8QrdA5
sSomvEV0gkbfA7Y0Y3bRJK3a6ppaCGJdKNvF9tZALOCcufoqC+RPFPS9k7FSIKKa
ubF2SECJJD/0ICxv9A29vyDwg38MjJK1+ESrzEQP+2QXAvgR+GpjB5seshslVkYB
O5/qjGvtvyLeDxuHj20pWTEFx9Q+6KWfPRWEs6NujofBOQ8ylI//qYaKo1mRJzYN
RUtlWpqBPAWkasDjnyVHxq11jGjNAC4ZNMPsmxrXbsm14Jh/Qrwsq0TMB9zscNZH
vVZDHGuPbIh+NWPP7FhL/Z6XHWWAMKBvrLAYOgbL6YFPL7K+Hy0iilgzSwa+M2Eh
7aaKfBYA2Gn9oqPg6VWwMP6fCX1zEAhq4e1TGDGzoXrQ2DqmFb1e5q4xEoYg0OP+
40s0SNRbwm6Tc67LKoupqN9Xs45n8mf5MaXfKvdHrMdqpFq5YNXoAg3W/bwA1dOn
vNM/Ws9Xk1NlDG8DYcA7Sv76a7HpmHiIhZTxLXTITbPXKrZtFQdcbUXzwYDIAmRu
sIa8QTadn66Q6fiCuaQQ294QvBTyhw+hkyEZEahyGtMJCOvks7KPJo6zouv9X/+N
SZ8BQ34KdtP8MnkTl46niCX51NYF3A3p1BQBQt4wF1Pg2k/ovZn44UAp+lAqLHB3
OeR2k0cyElki6sDJO0l0J6zsrN8OFghcPwvfH5g80rxoUb6en46B2X94jTzO0p7y
t+TLmB4XStN9nInMmkekUYO+Fg2p0kbfz6DCmBMg1Is0IEbhrUtF0VMTabXxE61r
gNE74Xz+n2vrlAbFoGJyYK4J//w5DmFIeD3ZwtO1BkT4mwcK6Lo3wdN7lwjxAXw/
G8BOsekU5yxhgmlbUDPUjEz/eOxQpGr31jmmT6deGBesIcyQrHVGYxvhkb4xvnQT
+WJJjxS6zrg6YuEovnQ1Q+IaYHmAFnFPdQ3ajDvalyzZCD9cuEADjznrItb+YJJI
9dq+xPIuXmfqueqZtmjWS7A6FLfC38MkZVn5s4qpMm5N0TSz2bs3KqbEA73VZJYx
Wwcc9o0R3VW1qk+Rd1kE4bjfYYjhiRk9Nlx7LUDci1tJmsILpIhFyJL7j9LZauHv
L8HuEv0iZR3O5JNEpOO3SXnOy9oWRIUWBjOA3Y5Q0o8MIJ7ABKhxKPaI4m8JpNdP
CaaEqhIAzh078jGJ6q1mm+ZexMUDK+O2qGPedIoHVqu3/vMsQyfloA6XjB9mhfF8
mHb8Kj2F017q/MFaa+/nt3GqiquHA+EJEGTnKxEUUaGk2cG3GJLne9cNclYhga1+
iBfsaGSam4j0rVuKF33aeYS6cxQSEpty64F46XEfEfZbrXzfz7vcJSUBO7M/a1pe
2fMq90rxtTb4wPuJQsjTNl253HNvfrmH6slZUxEofICXVff7XeEAtQleLXZaEgXn
2KcFelgloTLamKfsEAQgf+xsZOF5LqR2MQwJ+PJV0NrijqhQ+B6Dm++UKPv5lu+i
xk7omfjJpQAZ0OQXE9+a3o6EKLVWbEyi0B+f3RwNvens2yJdPDh2lNS0RqVxPzg1
xtIfCnFv31ya/ltyWuaPwhvVAinnkBf5lEm0tpGYw+C20JOgzhF2HVfX5W5jOvMC
PPphz2fdiE+1i+KBMg9noqUmsZtktgxA1Za7Tw3cOkrjvmhtiZ8EW9FCN4ur3Wo0
AGeuMIhSGLtEROkDrqIsDAmRv+JaOVJdL8MQBOqNEtZyPepqqa+vhCDWlKuSkpx7
Qho1759aPZ3J0NI275VGO/g3G8+slz14RCa1er44Qf9Kfu+M/IH3Bc9W5LJSq4lD
0CJEi7Q5vWn0K6Jfs4N1Od0RsfZ2mXTxiLxDkmNfRUwXM+1cSf1qboMny7yi4Xun
8Wn2SkSKc3hYJTjlZ3EAKp9R8q++qBfm7g+d4mwxria++OOhNyF4/x3ej6hXdjSL
Vc0yb66Df4n77st13Uodkb6o9YkH4mrv9kODuQ+aJpsvYFacar8dVKJhfbwWs8hS
36UrMwm84d35RWvVRYqnAwBC25xsVbX4z22FeWwXqumSvnSx8vN2si4v3QbLjpsQ
O6hPBgkqkcQpyFG/2VaTtPXlOkdS5DYH7GIeXNlmE39it6CvPK3S1YAhbJ/4JNpX
8cRFpNvGUBK2Dy4k3pISbTk4iU+1VD62/tBr8zS8+uSn41xOuwhnPYQilMXXtro8
zmVU2kiCsFaYEfJGrpToe4TKDV5VDXQr7VQkVlLY9S+sC1xpMUx9jbe9hCVWm+OZ
g/huAw3ul+gpRGa84/UWjrWn6LZVYY+O4k0zw1ZTbNJRQnJqVGDtBSu0z/+f+pDV
jH9xZ7D6z0bdIsugS2pVYN1yYuf9X6/kWVjSQiIsNzAeZVZbJbQuzV4c6ipyWuVP
umjepxfSA45rE80Oxdvj7BVmva0jBjJOY6nsefDNTPeXfQN+VFGW3NXOby+vlIf9
+vOjkv4pZGPE9w/QiguAm8gtrsx0GO1PjjOlzARGCo+yf3vsIh1cf/lC/lSB6X2A
olqq8vUQp5pr/VeKux+BJYeyypSMVrVjD2M4nf9q/AccjyBHd5H/v1lgTOBvRmhZ
wae2JVSYWO7OlXPDLOEI7XIgwJJiWhuNFsvIQ+PwRTFvQOMTnOg3cNVj44lDnWdd
RvGbXMHjp1ynhqSBMeYnPTpTRSXGcgY+f+I5173jGPkgqiGyRwZBJFQUa0Mt3VNe
+iTOBM11XCtpoJ6/dIioa+xT9UIRO1vugWNNW84xqYlfBPwFtLf1fjsthODLUoFM
8EImxb8zwm4xC1oEqijj1VEZh+cvgIeV2p5SBsRe/KSB+YBXxALW+VRmT63aktoX
fT9JYXKU0fVITX5hXEX6bkiJXkw/MXp6doccWrWKQykIUPzXrLXzQJslQEiOZ+0H
jltAoF/v6oBRsvVIDZMehvpHeB+r8XN4VOdc5mJWZrFf3Q09xUUZu/54FC1Xoxio
ozvii91QkEdPrWuMtrmSNPkrsHdAv+dDjgVq98+cLNeG6F5WC126o9DvS629DoYo
TR036PDmb63C72ZuwzouuiNqDStetFAdC2vgB2Ba80swaBLrp7HSWxfZZvvQqCzx
KGIw4g89vksh+qtjwLzx3LRIc7xbS4nDMB4WkJsmF6+r8Arjvh4jI5qKRqxvpnxJ
6LRiLUwXTJoyqbQbMLCsnXGdOfYJi3h46jmiqEMyccCgvm1eB/401YOiDiVfveza
qENGmmb+qrUYSlux2YB0ii0sPo2emTlV2xdAAKpKMXxxeziPQYotjRw3lfGWxtEg
ObP9Ak+uplOY7o6h2Yl3nWOAhBoodw3bTFOqFG4nwOWfPu7qYu8Et2tRWYwCaTUy
DYRuNhBz2hJ4hNYh03qQPCvlZWwT9myj3LJ7N3ld8Fzd04V1dRBOLDFVrRPCjr9E
77c+Q0GEGOLZALCzIFrao8r2iYFfnr7bYNSUDdZ45Gsjjb3RMNEUWtLyBG1zhZov
mzWkhAkpLdy6VMh/nW3dwO6QaIEaWAq2G2dyvxTKIHRVkrVDod5sTJNt3RuOWWTT
5awr3XayH/narMkLyhQzXeWkNnWXFnMu94owztamyVsrhWWEDuLDe00dl5LFEbcw
khR6rZXaFGVvF5bUAXw8pQMyqKrptDfw89tePPyKyNcVCcoZqblwkFGfNhfWzcP5
VexrxK7L7ZRASJRaIdBpkuZHZSEcAfFSpe0uYHVuKLWfUSjO0VP8JLphuThcAHvj
9L05wNvVvniDRJvFAHrfDGK10jbFZQZI3ZZ59oEy1Uc0aPRyAvoZ1G5ranbumR/N
F9EQuiKosHaHjEvwaSBLzGvcKSffhmCwu1PS3e+nmkniaHsnB5EwmrkLODdEkQFl
YcjiHGoOD24Wyh7PrEFCSOf7V7zEaYlZSkZfjBa1fCWTkWeP1RMH/gdHh0nUZ3z1
AXawMb8NhfZizRWUDdh+n5X19s0bg/kRcv4ShnfE8qfOqASMhvhpWbUKJZhXERpX
pakrHcXS3aHYJNaQLafxrRXzdKBsI6gqOzAY5LEwkAJbQXTe8AdMsxRw/bwpKYcG
w0F2QeOsuoHZ4/HVaX3aZ1dFkVz5o4bjElSqwGaTp/RV07L+qWav7tijRXqEeQZI
GZYZA3Sh3nLHupZEXNhicJWkxtRjKRWdTkBxGVEopocvB5AudPrqeWNQrR80NGw5
eJvr2QS7+n1jsf1g/h3hj/hzzicRIg2b21oTKBwTlqsEWyZS7Ka1rBtUxyfJldHQ
Z0mRp1SNMxWv8l+YkvbSgHf10jli5UdmhdlLNsu07nHSKI6ybrFamm2BBHHTlL7W
nFHKvZNgjsh/gdXdH0J+qi5kjonbe9X596rA+heGwM6NS79T3Cj7Y4T7LGzUi7ne
hflmfe7VSyOh52ysi9lRbdEk/d3UJRgTwKo69NhWkEgtvWzzrWQoKupZRwbMvxjY
k05coHlZGrTcRzgkxfb1+XCwyWeZdiWOWLNoI+OWHzciBiIO5KGHwgwExBeolIEM
ZyHYJA3zC6INbaj3i+Jx9vN0cAV7F59pvk12hGDCpFgyA28YUZSwAzE+/RK7ih/E
YnIUKB3ffnQ3dyfIY3+4UZl++NgzAJByMgZJk5/ViO7H624Mayr0VI22EoP+o+gM
iRoQUBOf1KNY2NKqcE6A22GG2lYpzSiJCp8OF6B79SEDBDwuLfe1YA/VNh4eN9MW
1PFxIKHVc63MBC7La8mNkPYtFn9wismxDVBLW9AR+GmsESB5hbIFA+yypX82fY1+
P8FS7ZsqRNJCgHVor+fmP6c4+zOobdJj/Nrptg6E51cHQ+4ZiIGb+isYW7BstTRR
IonrLu0GoYdygiXYYWafHITZL8kxhmvFD0gV2TwwftKj791Gphy37/pRbC2bCpYQ
9Rg0hKNDWEWlJxS0YsrfJ6ARGh9QBivV3eJOJeHs1Qmjnv200mYDyc8N0ynEULLl
ypSS1nuWdWRP6UqymoOIYrcpXdEHJXKH3Y7a84MwUrNgQY0vQERR50V8JpCiN9NZ
DfP5xgkidtT3Rx6yvmH1bzFfUV819rTrHMU4K3j0QsODlZZAYlp/EK6YsnJUpal/
ZVJevW/J5IKONWTd+/nilg2m9axGZ6Jf26G5V+Izc3FbnB4ztUBsQvayREmYqODT
OXLItzW+SLyC9eJni3frpGcuRCwb8BLTwXgj0kUJL7fhyPWM0nZ/0bbLyXUHKqOc
NYg1iSJ4gHbLWNvfJBrVoj/0zHlWUWhYKaN0eWPR/nYbElGmpjSK9lyyHkv8gnlw
159NQSC/TI/EO9flSArvdGwlNXPDqaHWOo2WLDE9zH/HpaGjSLCM8NoxcWhsRZjO
2yRlnIXlGqi5RDQCCcSGS/XEyfFrjRm2915MVxZltXjIqjjnGOuwDyy2gnA13GXP
zkh3uAVWjiru/xKutyU/fqxIWrwXueVYQs+req/rxFjC1LqBny+tIA2GE1t0aDAw
kdON4fPfHFBaS0R5/pcYT1iqYTwP/VTonTD6oD1DDqm7kRLTzVlV9wRRn6qa46/J
+zM3E8O9qH0cKk6Im3IvCoYFZkN/EQA9Lqz0yljHHCMc9SG9K7f498VO4yZaQAg/
ba95SAOYUcjTWtrG3Sb4g5fEsUxoNBkivttsgrZLkdM4Obxdvb68VAMrae2fcsJ/
Alz05Yzw8amKbaej77IJLX3895BtpJLVyMx7K+PsUL4fdxbTQkUYGTEpL4o4Qt0X
wKsOF9P1g0BG+Y6tuBqWsF58A+FSZgOYImArcVsEB5cfPKu6OVxwL0TMP7m3o3Mj
anqBJeiltmChhwoyq0/1y9/q6f+G7c87M3Qf+3Kqg1VpotsstX18nyGHwWhfy2uP
AxWv/suX/AWkO1EiVO7+gevbpF7BMjXUCMk2yUhUgo5KB+LfNJIyJ+kYHN9tKUnJ
yvwr7ghVzN+dyOQnZg5riMiZsH70PohzIcm5uXzEF73hggjTdONHav6XrpcSTX9Q
BNvOuJBed/6xMLjVkFycOwZqfQlBeN1VP7HcDNxUSPcDCytC+0EeqyyBf2Wile8z
mF+7C/wjU4YTFmFqXRFCqtdV8a3j1p/nOzSndYSDEMP8fTpEAhtJTUTDnOQenVH1
e2jmFJsQtggpIpqGaRQIob91Qcy2sobn6ImhT8t9Mb9YZdnirP9mrK8GIizDmCnN
4lUL6iEtiVDYIuGWnkbva7MtrBg1lI1LKL3ZkR9jdHacz1BNYbhniNnaXOSKam1o
QvX4YDrXLLB6HE0s9n3BAFIXCInRvjxW8lVK3YIRHTvDS73OmY8bUc96Ei8qwdfw
Zs2GxSFgGkA///9oqjJKtt/uwn+dCSOXqwGgyDlUPuvIOOjnkPP34CVKZrtomK2U
3FyLyDnGWwxZmV7O5ehsgi14TMEaYcqgEp7/ipjp/hFxsbHdaLMACf8xU7ZTuBr2
J3Cl90j7A6MsJlfq8EwNqiczb5ohvJzbTeqGw9yxzi+3lEtYiTUnhqhUggz+qoTi
QUtrY9AAVl61fJ4jc6o+umuiU5b4glPR/3grGB6SyP+xuilnmeDc86lpCHFONoVP
JNM+JjQAbdvtTu5X6Q3hCDMlpdbin4VvIcZSBSrXGxKQdeQopxZu8gp7igETHhzI
12AKB1qRSzDtcmE9tp3k+0MwGK3Rbvi7eMax1tga1bmKsaGAU03pHLs90QmGjzML
0xayu9obIVaaAt8UsebWRD60bW4YEROcnk9aeMjRJB64Rua25TGjTePlhHQwjS0c
oKBwFOXdwpby7DSKlfTueJjdRIGpxSaKagg3GvbQR7sNlQfR3w5ckr4rFsA5qOgZ
EpNGOfWPriG+1whVLFw8zaKudRWbsGTqzfojXqBRghA369q/MRPluquRAAYQ00tS
iW6zLu0kR9n/o8VHqUt6TidcxtH6ROSzjr5bkbE2/XkJBOJLZbtMTpVbh+1THxQ6
U8ad1qolQ7iVLg4WX3V65td5FZiOBMJGPRpzALmC+psfuAdkgJj1m3kQhSjnKcXL
pLI18Lr5eLP9vfflB+fp8naDkMjnSWeIaZvVOYc4X6GNN2LzgjL+KGe5lJnCi1Os
Y2I/Q814O+wzqkyHNS3rWsjyOEFdiab4dRGja5svlmcOvb4qMw9YgGyPlv8zfBbx
VMNUAwQ6ayPv0xBsR7nBtYaK4PY5qokQ/FfHFc7teTPa5qL4+lzxh3p+uEQwt9Ps
DrEbvS6Ose8ONhNNng79xUrajnfHHMR5kS/mPODnU10PS5/rzcFUU8otGAaVLzml
LWmmNSOhA5w36uvtp90cY2EbXqjUrD3sl6JEayVJyhXWP2biKBMFQ+Q3k6UejfIH
/8l06SUFdW8gkfdgiEfdKwERXdbGN/ubqTGCe1IczQxfAfFl1NZ84OTQXxDk03KA
J8Lq2abKNVVJeiIfh4zrr7+Un/70ctTNcAOJxhgFCfWSjenI6GVJ86ogr5v5sJ9G
5dtwCae7c4RIy0rq0thwpw8IC2ctWIqlyCxF/LXfCorIrusaUriPQlknVjUmj1F2
G9N3vheluq4nXOjlp7ssCdwYrgo6S5sZxBga8WCCuanfXktXdmZpNxRnRh9gSC/M
FpqkLdwj/OzzYeXeMkWV4pJ5NFJFTLupVp5/qqkRpKOENd4jRUJ9RFZBjYSG+iTt
F3HqWuK1uhyugiyrosICIURVEFVoj+rb3HQ5qi8CFIY+cK4vR7jvaQyJFilfwrpy
61Tsd0hkH+KrM6brSZgJvPhWNdrt2F4WT/UJxxTP9TeeGXUW2JBOo6fSkROBlvgo
8h/RkR+eIItIUTup0/NmPb6l1v3S+eW0hE8QUWfgVsDH4TaaI+LH+5EkgFTxStKK
Mf4KQheijnFyHkm0+e4ndBld79prx2HL/sIlJeFvLy0ypyVyKeZ8F9RgfsbTXGNl
ipHwGsmhsd0HsBFgyBEitmGaKjdrasHuz5m0PJE3jYX0kruhgkKgrp7m0GHfATcN
tMH4eP8wdh5IKYR2d0V8kr7lOnUEfQCyGB4paipO/g6ycSXeDuIZ7rWo+CEFZOIV
lpGI5osDQLlVHAlUh2HJBG3+cwJF61F9y2c7I14uQgstDRvsbzbhrD0lpyveylhl
tXES22m8pYldBogpKcBkv9SmgMVD74ZBlmnSJrlgwjVlYIdvAafzXfRGb8rcBiuB
RxuozMWNpXFGaDmt35ZOEabzGnJGaJU4z/pzpX/5lMUxUNPTMj4seZRru3rNxVU3
UHc32gmCReU2EE53V4JODQzx5PN6i1235c+zqtGbBPTUDNuVU14x/UMD53KM0Wo5
Lar0gEJFGwzzo1orHItmYGAF/AeNGoO8wVvATCDT0Mpb0FScYujiUeEN6MZaooAi
X81ZKtCJoQrKFlqUEvEjiuSB9B+3O2Trl/8z/6XYzOviZF4uUfw4PIF/QrlS6mq4
UVVaWhV4Rr9b/nOXzQ8p7ZnRERl5x1JyJvDXz/DEptLNj11k4RqbYWqc1umptP94
WMYnkBSDTh04mXCsxcxf42Ul6MR/d21OcklHsYXjqLb2lC3cLbxEEhCAapcy4Nhj
1rrblsthLgMpLjFOi72c6N/X3O89p3aUsonNydEENvWtdR/9Pu2YYFGQ2ACNOk5M
T1b8CgBMCYnPKILIGYl6VFJrGp+eXMiyjshfuSPmOd0NVZV0yTywRBk2sj41dNnG
5Qbdr3wtjoS23VR4DxepYGidhpYvkcQVZ5RSRcTqMP5FEvnHR1Fau8Bqp0SURvop
ne6tY8JlaQNas2NHJc79eocVVRkUW/HadtM9dTGVMdjMEzRytZcDFNg7XRnLVOa5
B8E7hYdhHfQgVsk/04zvHR1gF0msLvu5TOYBTxMkAor9uaoJlq+1eV9eyyG6/MKm
JJRnvWp0M/F3BrGXBlvRghMQaZiafTHFRdp4uFOHnWz6oXEj2Eghl4Xp6Ur9HpzM
QwpZQat8OeUbk8nnXz4KsMkxK3TEGpC4CNrEiA6HvwG/nHIUvrbdWxnkLQEQHnKp
uBZ2DubrmiekFS3XVP78shQP6Rn0kXI+aE/59mbQMVgF1+MTGD/lx87TX4P2ltxZ
jxqBCxVjm+88eyFicMP0yJ9m4Z1yCX8gc7tKBL2yPatdJiLmpS8labhB6y5x9Mqf
pD2g1GMC3aFRrFlQG5TA5UI8oF++IOdr1a1FZ+1/HKEhhjPtJOqZsWD41kFDJLG5
I90A6YtnbduQIEl1gKBlAacn7DR3uUAgrGiMlzfm4c7FRA0BOZP//V/R00e8I8ST
EztMSb9BqjNQa8BN2PGcNEyINRpspcO9km+x8IG52atmbgrqyjTqiT72el/ByR4F
koivfmMKHEuq4H/rnNpTU52qcvKH/ufsEfafQRj1CHFy/90HQ2goeNqkwP0v0lHk
87RteBI/Aqck+07DVDPI5f9GB6e4a4imnKczkIrHXhriSo0mSWYC+B3KBtOziKSd
rKy1ujcUVxL6TdBuwobxbWw6DHX6OR+/GMG0zVXhFM2mVN11sArRPbbh742PbH0A
2pcAtoDR/gc7LwbuapV1MJa0Z2LTMvsg0I455Q4AVaXFdue3DpLX1WEiWlI5meBl
JeafS+0JbofLvmrUkiCOeYvJqgvrLIDiiI6OIQgIxVQzQOwzEObzXQepV++qajBl
nyJJDDGrtyCVH5dhzpeatMC9s9VkHsIX0C0LvIHeRa4u9lf+NUZ5n5QrB4Qjwy77
phtmuKtxsBfb8cKVMirxpH1fxube3gxZ+HvC/Uf9aQnzS6hSO3JyDanx6i5Tocru
Ab6muHnpouAxfbIhtdP9HKXhcdEudP6f9ZD4zot20/Kq6thEyragu5UYrQmhHiyJ
UMIXIYSaUf1OhCzWdTHvPoA92ielKJRSJWrPO2wfphbpj0Kb+umXk5HJFytGtzeF
8Kz3x5MVfU7F8HYbjUWETyEa+YXwVyMbfELpNcRyY2OQiUWCxYivIjgUrWUeFLjR
7K87wstln57HNd0wAraDZeYvymWuI2CPkhDkShfqGS1Q8cjvWhdAt/B9kJmXRcF/
vCpnD0X7SWTBlkbTPj+VKUA7mDH39Ec5GTQFVkD4yw9eRBzqiQnsNPPjb6CZAvlB
VOhtup+USvEjZsuW0PJfEuIhDVuAHeSAMU3aZIBZIkres8M0KWiIe3vXqQAbpFFi
ZPGqUgVhInuWO0ei85/qxWMkwi9WlARTPTKJmzWPRVXePF3YyzJyppP849ttADnl
3mXs3FblzVNblJ/QYzYbBzFgDPojhl/If8QTaSFa9q8HrYfTjmZpemMQAyrERQyc
4siXwSJG6Pqb62qUZQpZp3i3GfSBuwSSlZNPl8pxzPHKuve/oa/nPp9Zki1LDcF1
gPofoy+eRLyEt/1NToe6CMjtJ8ccJHkLg47Wg3g7Cx0ix8/+RxmACVrjcwugKq0Z
UJwDTgZQl2o/GDC2skFBqxgWSf2/UmCMHtukgEHGBPbfL2/88uvs5fcSwN164HXc
mt0o93e71s81Yyjqi5YisWp/GdtA5tZZcPLTaTMuLf4+Cv9AHm83dOO1FFxOwdRm
vtlc0xH2ey16++R1fQuiCVufFXtnm8d56u3wuWzmUaGNYKYbEE17gehhqnIAfZWF
xMLbyLl9i+h/USLcoLr9hIBgdkxndUT9Zrs2oKi3O3/quKZE1cIQheGJhGIr5pe1
mo7tta7Cs12q/A+aSarN3nodlBvRczRCYOhssKjzo4VsDrHWUerEnR9HM/CLltsR
BUGYgzUSYo+kdWmcovyJrBl4ndOGOC8L1I9LNUyZ/sOnRZnJAsIKQic8JIVit5bm
yMlvfh7y2uzRUy0i3P2DWXFCg65dHvTwuK8cMm3woJ8nfPySodjW0S0e30damKGp
EM5Kk+XyBZ/nfn7CTLjs/u0duiEl1M0Shicm7/S/IDTvV8ZIva8kSwQtSG0OH6va
C9jxWB0w1dbII2E+MeRww6kF/VyZxqo2mXqFl5foV8YQ6+OX3Bb1a05MfsOK413a
DL9E79/gosPKC8G6sjNHNvkijJNyLCv+V7YJaUX/OEHfOJc+fc7de28+wKjY99xF
5F+FWmhg9Ng1Ex0qDlA6cDoMQ8ntrfGVZigE2RrxGbi34lVGrkh4AI7W7YPBeVak
hhhvKcO7OTGhUSIUnnhSX3TeaUwHyWb9Xl9xjhHSiTYEOxer+5xjtPgS5p2DscUY
cxwFWhH00Y1oJnjnRiywNVT7HndsrguHy8Oj2SGVNN2DMjHkqJnqP1T9HqLlTBPy
TSvD9pQUfMrX8iwfgIGR92RSpcI9byrMPRrCHBJYsu+I+5biAbp7L+MJy+/aaYJk
pVv4sbEpw+1fIjskCYjAiRln3aUJ9ztdjlRtG1yYFsk671uEVzbSWMcrL1ULo2dy
SFfZ7EdOjJTBYoTm5ftp9obYSkcvmz+h3I90Edmzv6Fu2hZly1u7HRxqxqc5oBn7
YJLsp5s3Htv4Rsz4GjYFiuAPovF0YYr+hkYM65XZznbEa8V+sL6o8W9o0wPUBoSo
gJFsrQltjaIa7hsmyx321iQskXSuimW80ImYHleIugWI28Li7CQ4NIdo1s8+FtdS
0fnj+bxHjUj0URBo/akG7UxlLG5gaP+DyIpU76B5gahLKZdpX2NWElPmCSZu362Y
waRkbUbiXLCSOMkXlIuLWl8f16PJySCW/9TF2cW517WyGC7j+Vauez3HbWoJX/Ky
srXooUVF79zM/xuLdmbqeVmOR0FT+vqO64l8pbLNH7pK0H6ZCWkjAPEjsEiCRg+7
PAMcdHkFpT+UoFrWtmj0HkE4fjCWbNFvawYFwuArc0V8QlKWcquxk4pxnpm22TJb
Dlfb/VwELfIFPcu3INkPavv9OjpGh1mOzgDScuRyj6wHks8jSkqVqwLO0MysAkbY
iZw+TQXL/CxtMUpeo3jBLbfQHlWn2pXr0lYOQEfN+TJ1CnMOa67DlAbVx4x16LVi
1ocKLGm0foIE6e9pGwXi4xjSzauZZjJvpWd4BeTC8872gLw8YZL3IinR2torAo0k
0ZKW8ww43WbtWCHrbhwuSzIj8l4ETHCmmvAqTVxkIhsCz3J/NRL54fBhFSLZww/t
SgTC/mjr8J++Lx0YXBhXcz9yo6QaYTAQ/LkJX/3M2eh483jyHZ2qNiMA7Nyiq9LO
zWW+LVPYsyt0Xc17Sy/JBVri7ufIVgYwjbylgd/TPQr0AhHETkLSz2JhX2gmTuFX
lOWqH8E0wjVJLbLqAhne8kLHOaRkeBfIUWy/LezxQnqiA1MZ4dFHJKT0R17iLbUE
6Nq0dd0UBmijkn2zC1lHb0fT+Mzo/56/Dk0YsOVWLKCSuQy+lhN/31kgN4yUuqHi
kVUJnWN5GuVERfAgNYqHP2ylA7P104RlICWOGyumT2XrE7kIWHPA2nd5o1xro+fN
BMKrl3zhfbP0zXyXhRoIO3B2kQe8+jMZ9Zjk5PtZBtGx5OiJfIFrAUUeJDzSJd2+
bbxrgbFjRSaFhcyuYC6XKalPtD+jg+J8QwrToqdh9mvRvnwZiYtakXAAZ9lpCZpc
/m9h+OTQxkOG4ejBm7T6xOg1N2citrFDmUV8gNtpQGmQEN3RtyhRs+abfjIaPpC3
ttchDWWSmfxJ3ffV057ENqHXcYGVXFRDUsqMgpjg8iOik9fbyZJG4O+Ozpxpgt1W
2j4sUIJznw6x82dlqkNnDOpQX0qNrO/1V/kGevBrkTompbVYsf9wlQdfhcbui6D9
JmPIFQFHRbQ8wOMZiy5oo/NycJMtbKKsd9VriMrdgxY5Ib30rKXUUSMbG4CgbY6p
JLViNB1eaaUmMfClXBOONwwHW5b5wgZj/ZF4DLZ5AB26HtxF10ktU1Jp+YrDCnvz
44wOPNisOPeK1Y270UgJBKfyql9cCxmQAusbprfE8g/XqlIEMriKhCBuIvJqZ/1y
BUMYimanbfb8Seeiom/69WGHRc+KyyUi4IdFxt8mDPGaMiuIYo3WwvnS+MADfGHA
6UYXJNoi2xOrzcktJbiqUeYsPCQ4U/XxUsBahKqeulw92kx55Td0diT1m8U9ISMV
apBkV6rPc8sQhZaVcfJFulam99t4h8AIa+dawm+Mu423cfH5nJZ9JhmPtknUXq1C
aGV2t1IV8IdP3xCkDgd+Ae6C2e7ouZeerP4NzffRrW6oKasg8vhZ+y3w/+wgbX7k
cgVmq3kwNsp/fo7G7pZibacNM6zofEJFREf1JKQeu0iTKx+Hq12ZKrtnD3H1lY/p
lW+KkdRwvz/TlPxImz9Jc4ukwT//G0Hw6sMxfPqKApcKCLr7cGTrxinsEZfRaySb
xZ9ZtTbSPhDaKYmfG5LZFbwAr+0H7mu7or9H1JRXgEDzVrGMJ7I8xQp8Vq2Id7NH
w3lTMSg6Wy1GQPi5Iyb2Nr8JoQgXIqZ1ZKJ++Q2hDgQvodigfAZ1r0I7dCRyRJdE
O/NNkFYC+8BhoXfGsj4QD8DHsKWQDj4GMyMY+Myhwjn3/etWAmsyiusz3zGZvFH0
YzXnyyI0lbC8wxgjMaKC2tOBcw2knUXg+fXjdMlJEpMtcm1BZd3RICb7Mb1keXpZ
1MsChtVasqGQ+lhfBd50tvTwo94ZJG+a928qz47paNHoqivc/W7CIBfnYWaQWBZi
CNChssR1PqwTKkH4SJ8lom1IHfiQSpPICMVIbiokYw7NHj2AJLKb8b9HYJh5hxIa
tQuYmCgCAP4gXQvCE0I55+e9FZTivv+Jty5Xs8khgV8KVOIbHkJGdgMUc7NhecUJ
rXfQtMhk8ztNxBqaV2zi3JqJKFIGw0vhb7Biq0Nn/cjC7+Kwer17TsnksyJ5w7FD
zl7k//VSI3F/wLIhoh3Rfu/kkkUEjqsoPlDjcx3W7GBeCOw/7ZDzGjREzfAYhZMa
taCMOWxXH0nVOCxTcVWkBcYj50+Tx2qTD6FwqKG37JNJRLSDwOm+6E0ZLkoPG/B8
KFIM6YYfAu2KYDj6mAtIQunXTWlj2mTudxy0TFie1oVXkQomXObG96sOTiT7S+lv
dOkhLcakWledmvmjldvCCGpxXlc4wGvW9pf9jcmmIiN+30MyGqea6uu85aoLX/X9
EDQnrw8i1bZnZTwvkLpESrF+B3thld9LzOumXTtvayQs6DCmsrkNo8h+7r4qT9W+
NFOd1nJ0MxK7RuQ3kMHjKbcFOAN2kvL7bj/3BrWVRKn2RPHI+JpNeXWAELVuyVkr
aAiUcCFanMDr+yW9ax9Ox1PlJXgqV6RZAo+hNYHbfI+L5K1F+9+ozYELbRXD7c2x
pSmqLgFkl0JswGS0SKsZlKya4IO2gpKAPssT/KtPHYOc8Oh2mhKHX5Twl9Y5jOyj
H1ZEx8Xk84gEGL+3wNQJ4RJujpwFjM0VndwZr8sDtZEcTKKg4UtTDjY7koHMa7lu
im6J5ZDuJm8qeN6D+eTCbn03+oTwbIkUDYnAs8VCyNZ+50J+A3uzHJa9BU8O6tv/
eOLbx9x95Un+FB3Y7vJNybA/Fc2hPtwciv9NyR7dNRLBcii85Z9JvcMdFXF6b6pk
55zsU5BUdX7UwYV1sl1jbxlrkILzPr2vEGLDZIpLKiBfY5bhEVBLxkURVWgeKqvs
ylmPLMuM6EHOY6fiU9eQgeh0O7OROq4TxtsqwHWM0IcTxPCnpfv+nKyxgaNcwjnq
dClp7pLfbWfzcC/AEmd+SaLOuOErtg43yH5zMTIlrBZfZYMtgVqDc4dfYlLESl4x
Jc2/t0MmBq/GKFzFgs7qyYl8kzjU9JknWX9TRo/3NCTH0Js22KFN63weFVykCcU8
T4a2VYvVdPdeMzzFebjaV2t51++kMVdAAMwplUZflryXP7m4rP4mfZJ926glhQNw
IL9zPPoTBXw3rugFfmZVnxTBT3bRMcE8In8OSVUoMSyDPSXJy0i5Xj2oR9QrGlsA
m78Y1bgtADBfoXgd9c+MBcIQvs+zMG7DvXPaYkFqHNML+MaCQxnGbVRoVa3DzodW
7KMl3zZOJKR6N8h/1neDZA7zB+GxzIao2PBR6G2NSzEJ2IwwKD3bKwsb4KVr9fGu
bcr2YGRUkuAzKJwpXOhjdkMeu1thuG4vyqoTzqrOgXK59wnYQ8ZhpbBZxzbgAw4h
VCWuredla3ApyaMjL2NAa2X54UYjaRUSUDlQV0cHTmCgXbA0f/Y17V/YF8sNIWGk
qZO3Uq/JBtMeJrkn5PbZtp9sXnGwSRwl3r83QxzzSJk=
`protect END_PROTECTED
