`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UUEWGwetD5MTRm8aACygni7zQutPmNyZCkZQjCkEd7C0zNEQ9RVZFwtx2zZJxvzV
boCtQFJ0eK1XQX+LtaQWfGYZZBEs+ffYG+5xzo8ygGrBAIxcfSzI6y8p5VIPNCLP
OuGM2/vnZAe8nOzIhGT9sGkGnstbo9FAQrwDyZEZ1uZ6mhy+X7qyu0pBhTPF7jfB
0A6CoTnnUCWEOflqz8AlT4ftIk/czn80mWtC4vDFvEaoiD/vbnBRR5d6B4J6mnIg
zo5FduEwXoQCQnUcAJGKvxKqH7hXk6q0+sFHZIiHGDDRryyOOTPK8PgNg7F2bxRg
QpLetiSrmzfKhX0b4AA5j8Qm8zsVhdzyPUo+ZScC59U8aEwqWyrtxfNwk7lUajO6
Uzwf10iFXA8182jOT7BOG/5aVpXdWW4zC4UeKNgbBW/4xH7ZyLIkz7wntxe6KEJR
5859UNXTpvxC/HVu75hOYf2unyOvYPvUw/1of0TFq+BvLAPcby3CIeV3FKvh1X3E
Q96ascrZGhEzE/Fxv/ZKcFz+iAuxUusi0dVKeE7duw9+hQtRNsgh2zfMj8Lop/cf
U4BNgOgnSiH8BkemVLPxiPOG7+E0zs7XO8bobaibsl6pPKJWH+4BRY90+rek8yOH
dHGaSkq/oNuJBu4De1I9IfxQtTlHQ79Ki9ufJnh3Rhg3ghhZhRhYry8A998wpUZx
rpDshgCCSuPgNheUavuxNDgTXVL6c1Nuk+FgZZTC0rcRnE8yRoDTBhwO+eVUqY7T
8qyMvLILgr5fXG0vBoxgfkxB642HSdP4pTZito1TEZb6RTCkY9jCjfxo0lHoDJkm
g6fY2eUYkPx9k4A3pPEnLwZzdOH2cv2tSRN8ZaTX9emvzYMNtXJAXWABYohZjBHE
pQACeqidmtqqoiqdOD8Guxq697dU31oN+Zg8VsB6USG9RgelU8dst/xqSq5iHoBK
Xes1Z93zPupmOv0Ak30OA2Zzm7EMnr3WM1DBpIEzozIXETgwx+wO6lEv63AmLjOW
zhXZnpBYo8L40XaiMkiQb+a0hHziLIDhidzKKHz0Xdk2wq6j5ljQSZKEdiaWlv0u
AHD3ghrSUwlqHWPYUhrRcvSuQ0ZIrEvqjOKLEtJyiFYBAAwSwaueAApTTAjy2XQz
ncyL7f0OCot2X+821r2VsO8swnnvq020tBpxVY5toBsHxoaBUYwhYNbfZGdku0OT
b90uPRUCRTp4rAnzC5TDgPf3BIcROn3cQtzW/qJmc1CqSHGOmVzOwsve7DZ7TJnc
fqZhV5V2uGpWDIMjdsFkDEyBzrV3UbFeVK7S4xULUXKq4dMKQJBfORnTzJshV2G4
NL+6FFswKx7XJ6kuVozrU8nco/Mo5pzU9u+IGr/3DX/fyH6c4TkXT90P9hSblMir
sjZIyx6aZKH7cQGLFALyTA0AopX3TEs/irv4Cel+gPmPivKAys2xBUvpDSfHVPxs
VMuu0p7R0RuWqnsx2mN67MB/38/jttHqojok77f4VhFPeGVNvgTt0VMzlP1uvERJ
jcmcqS/U0ZysnfQckjlxv+Sfy45pwnnj2uGT7nvcEcBof80HCJxmDvKFbI+AX0nd
3SlXDLx+iN9lCPSBFVVzwi8Ff/VYRem8qyrIYNdO7I29dIjpRPe4LkfPBR2Mo2pR
u7l3g1weQfORe7aTTwiRNYVoDIn3PEdcImahiiFyXjF/wHGk6ZiokUFed573avhu
OAZNI2vNf0MijXi6QyDWKz3PHTygtxsBfUgXC8jfHdHjj4/anEpA7CF1if7IeWVD
IG/SX9e8lVk3eo/MLIwphiKMZoqdye6MRBeGaKF5hJrwYvW9N8Yq4gwmhqeLX+cR
yh5TOETxDo744hcYJEP6DJ1JS9nLFX5EQ2ggHijW3BwtdbroOxNYQPqdf2E77UOu
J5jQ7Hg/pEBmYe5E1Hx8m3OZQjjK3TgQ/7BH+0WtIr9P54o+fnWr2jEjjYX2tRV+
2H0vS9nrsmwl6mPwa3STide78VCiLD8SF5KxS7ZvSOoxGyFUBLJAHlG06vVi57Hr
GUY2jFr6MQzbuKfMIxbQbKHSTtQwu9iABiWrwTW6aQeXJ/VMO9NCnBG4LPDYpgA7
sziQdW7dhFNIpq9DhL+IjmM+uzhnoi5H3IXWk5rhHnlD/591s3OryHiF8CW8MwyJ
sPpTsawWty6E3u+1P2f+IwntH9VaSaVjvrdNl+Bo6d413ix32e4k2IRvgiwZJszG
rR3Xb+0R/Zae+wJ+bryURdytrY2NRvFSi4xoLpWvejSBJvHri1Qhoif8xAOqMu8D
sHnfZFlJw2W/BFjwP2TgrEFOAW0NwnfWuUVSMecUA8fW+zt4KTuujq14p5GHt++l
UvFGtvL7uGR6tPYotKwC8REhet7fCTbArJqLpgbS60nSrP0g5nRkMvNstPTeidsy
Vufp4KoU7/XjuFEHRepYXhzN4rJ2mXCYIcVrBPLN4j/xd8yDHClogKltR+mfdPDV
EE2uq11vz23Ng+Zu2hHOwG2bd9DbqyRLWiKh6WMp0uKwBGKvwq6TX1Vwp6FfZqkZ
Mr3Gw2eX8zHv/zUm6+kw3Ss6ZTCxkGLXFsuX1Kigha3BOEJtMxB33mWUHsgVX111
y3RuJt2e/Zm8ng5Y8WSscG1ZIbbLEqkNmROKQVVjMDHlwuBITqng7m2Clc+NE8Ji
D/AIIimN64CpD/QicHzAP1ZIbfTkZYgW7O3/aFlzeaIxxPNaNFPIBu0Oy7bUQdAI
t406vgDk7Z7axFT//EVFEzneKNmedzifMmoUb/J1kVFPxu4yel75XXWWrG+0R+Ba
4yI9RSwUs6X0BhSc0blfEWSt2MNJSVylI82X1beDGKoMJx0RxtodH+u7t3uZZkFg
LmXEgRr38G22eUvIqFWQGMAHGoyy39Pd8tSBU40qupf78YNvTXgx5GRIcIim1T2q
3FhZJ45vEufhqgVScTqf2Oujyp88ynSXbpigvLYneOpWjjAW+sHn5TQOFDM6w79L
sf+qEoiLT5BESvSVzt/l7sBrNGmbn+PZBeZE0KbCQnB2XVjRRVL75oBtVhkR1DKL
Y+fiuibbfl/VMEK3EB2VBF84DbYcKHR2FNXoMA/GxWUPZG+igM1rZ6qZPnSXnUIr
Wv3MMfmuzy9nTfuBj/5rS0TJLKp6fFHX5ZD5RK8aHKzZ5ZGRKxfEDluM9DsUzmLj
IxIbU37EQeA0wMx5kmGVrFJ7Bj6Ig7BUIhP5NrLJlHI+a72RXPjV+HxOV52cVuV2
7lG0XTE6iR07ptC0HmY80iytOKPud9vtltfdXuzlNshPvOY9OoJQN13kk6c3igwz
3yBM2cFmx3tG7L/dsbz5CntocQU6eSfc4pv6RCNdqjKUvWfhbxCOTTAQyv0/hUQX
QAj1HaWjPWsFncCSSfSkbxPPXV2Rwj/nnezqw39ExBDKAbntSWMyAx8s+5Y3521C
asql+fCXhv4ODCvzWpzBc6Ht6hYGRlwsKIsl+en4Wvkw382WlL9BIaCxMVOCn2bV
K0noE1tpcxnzgCjqFxvEGi5UiQlfRdPeuwnqbVLWdIIZjS5CXP2j34pL5lXmsXo3
/DYel0zTQfj1iH3l84ibJoTqKUJYBdWly7TsSkTRaCuFBdxAQxr63a0rLysUI706
nnspo2UCD1bEpaXoloYUrjlCqtGCnX2tSNc0wD/mhKQAaZOZxJWrQRwlmNDK2l+D
Fxjvdx33BVlWC2WkrzndMMEau+p0OG8eYRJlO1brLyJ+/FoNqtVD7q71p4bD2lQ+
xxB6p2Hlqb06rBJ3v6rG3CHl+w9P8IdRRnINWespl5WyayHiJJ+9/sSHA1h/adBl
dBn7lo9RHxqMPommtguw4/soARSmd0hdetsJsA+x6M4pJoufND1BN2IYHjzyF8B/
3eh7ZeyrnP3HGWiODsjEVfGK3OA6N59GtFHS/MlaWR37dK4/thcHRwT8iZw0p9r3
VLKn4NGbhVfQIUe4+X0XmLVsda8JUAg8j/J6tAyiUNhSaFGKAS9MZmDfHaxzxms6
za0KCxCZE+ohWPVVOw6fcJFgFNXtgzcFGVnDFn9h5YTGGtrEdtyNCcxvtFY6QTLY
h/5TXZNrbhq6Dxf1E0Bt+L4DclOyXGPsPYHP2DbtRNjPQKBjZIP6BJHC9vrK5VG+
DJuFQx9XWhm7GZX+JRI4KPlocbsjQL6COItj8CUUalnxfsOf5F8JewFUx2n3p0pO
3UbGmCmuxJnr4OhQCPj/MZFWI4a1253/hvZjfVcJZdwuEtTrMVdj4o0hsvX1WPG9
ryUohpqJdJZ+Mcj/88ugN4VeWzRWV57akiU+4zGUAiVvp9gh8PfokVeRJKdcul7s
6aZ+u0fKS+/cVCNzVip8oAJEJ9BQuLNrDJMKw33f7+mptLyynsT0T9rMEEVS/UIx
2IV+UIRVuzyop8ipEehBEbtIz+SsvV8ZQ8ezRJk3u62oprEht2JmUm1h7bt9XUZQ
9tg9Babv78LXGMArpMSvVif9MwzpQhuYqpkratJ4JFW3D3xxuytR1rnJpHbgk980
YQ1GqmmtHMqKFgqxjbJZwsCM5aIfcHoK3WpZgiY6tn5+RpOGHMyiFbZ/e/qt7wOd
ZgwsFh3On2ru1oTyPsjinRwBlPBYKXPwoz5LMJz/5Vxmx5nNeznf0IBH6L9W4nOw
9hZUfNNFHESk2IaV8DFlTB7KveApdNOctU4SD95xNvGhZYTxbMQW4q1DA4K9nt4+
SP5VDlcpNSMxxJ4wdjfc0oaA0X2WAJcEOI2+3ac3RJMEn/8xX7MR+jnzx2eQ/d8q
XoDVjX4i0DdNNtEQ7pzzny6fQ1o4KAJtq9sTCePn1tjZgWZUq6c3CS8bEAtOb4Bx
SlOB4SsJ1kM0uxUgLVzhsO0tnL5CD6ofiL7QvIrwJZQOh8NMzW7Pa/aNyiXUDYwc
oW8CbycWlvNLo8E7RsUNmYJmGR39IYzVc6xVT3UfuGjkSnRYgwwyjSDCDwP65JAW
nvmSLmMWGIPpSqVCA1VJyoxXSAFymktvTdHI1Opkm50X8nYBD3VbdkGfrvDoH4Gy
/Cg/nK6M1So/rgKab9XBooKxqmN+ftIrgP/adGId5l7eiomVLrp5EmQODzGVoBr7
lNm6jBB8WKhe7tmTSeYw95v28kSkJnnkHI2yLLkbLDaq/lmjCJ51zsXte7nuHVI6
ho9jvhR9Lv8H76EpLk2FsEHrrP3FIQLdPTFo7j6ftIxDpyf/1/7vAiqKN7c3wk8S
jwmpms9+zntEAwvEkxeUsI1uHV1SM5ro2wivlGg6TR+6wVWiXNNIVJVFndcSzWJh
Sl26qmpwj9ufV0CNueGD/ytbEX4fsWKkvde3D+9qdXnLqw4szDZZcmqFg7XTQMWq
s4fbwJFFpVsp0slowLBXcRredX/L5bsF9JliFkrlVjr/ok3Nv5rR+FB0wd3u5HvC
AhFtlmQJ3eLBgud3m7ENBmgg/gfw894NBltcr7YlAfZiWWnzWvAbGu3iF1FeGlDl
ve+Amyiaxw1eTbcsyeLvbcsiiHN1lvTNIKcv5Qr0bN6pV1/tT8lIlq4NOJIHfp0O
foD15yryYbTm1e2eaRkLvDApvAlhd1Hr2viDyEUhMfKwzWrh/SM9A+oRStRyJXS+
KZXlQM8YxLmqR2fHWEKM6llBjiVVGQG/rqC5ThJ/fXJPbraSjbrGbbNFAz5J2PPg
qDTQ7gBmf5hvfSvxve12E2UFCndhMGpq1/3UQZaeWVvPiXec5BrilRhtcl93twX4
Ydhuzw2+mKQXCjh9HNXW3P7EdrUBb/duVfOGx+ahy/xWgxMGBQjow/RSJl9Pxu6g
d9PetOVHbN9S3+TOwzOiwNps/bJeKMRObLPfvKsQWZHnIRfNFKlKuQ9e0vcotR/u
AcWXoyIZvMdEmL+A/2XWByP5bUpsYcH5hFv//z7fFQ8zZzknNywQmDvTLKqTeTty
DoL7OS9504t7aPQwBj5BtbPAjmkPwBQyOBVsNpBBtGn6Acqi4PAoGRD7UiFA1GZu
a0a8T07N48HlgyZ1QLamri5iMrp0upxlAlAgIidhaUvG+cYaTcXdLUaYRZuwyU7c
sElotOseWwDdfbewNSzXkLHbcr7EanhVvDWjIW9P+KtEl2ilKNf6WXBfTabJaM8V
aCGVm7NIYipPzIMhElPV6pGsW2pX6bKL6PFwrpOcylwn+2R99klR+ZVtccdoPXhG
wDa4MGtvq1qp95+EELlIiYCoc+cJIJ4+5HhH4Hlm9ZoFhy9sQ2c2iSY17VQD0on9
Lh/OusTwzs6kQd2fKApRgovas/SR/fF4hrc5Tr2JGY9yoTP4YyW63eNJxKMf8JLS
3hyu/xxi68DOTrkK+/CKibO7AKByzWu3fdPp90WdjDkheVIGcaSwhmDcrhPR4Hjz
s7iZuCmGN0rZHjBp+f8PVEeJBYwzF6td1cjUFMC7/U0/8lxtbmwNA7XXy8yIjHHs
tfPLVLIf5i4SkAm16H1ArwUO9pW1TJq71fPfeoLNn+76uoSEVky7Ql0qQ4r6hCfM
DVQ9AUxlmdryuwtkJ5bx9guyqvcfh8mRmtWcEAgH1mbp9dPtN+w1+DE/ADDuFyzV
ENBQJ7OQtBrxGJd7FJnHGSwMrsVYLZqxiYcLRxAyC+MnAxwqlua10+yJjxEu2qPQ
E2PM8swrknbfKwwDYA+ZSKkP70nO4Zi+XQQNq/iAlkQ81EMNBOCbM00CK26acxpx
5ER3K5eT/pMNAab4K8mb95PgDmZ/pEZjm/maXzvxv+uy5G8UMXTSOCHBwvX9n0i/
L9xvzqULx0Z9Kk2TlVjPszJGGkdbCJC+INIWFXZmrEV0hQWpgVQ/kV6ie5afcXPa
X1Stko0sczCxmPgrZwT1eLPhLGzuXIEoofzJS4wiOyfiwYExfkoXK6Pnb+AHqmOA
Z1LZWMHIRfIi2WkHEe24ZYD2wU4GLMvt6GtAj2vRVkyVe1qZrFBonXSieUyBBvOw
C/9dPP1m2RRTV0BDEj+1OdDOSWq1oC1vH4TnNM2hg5dIbFtGD2JCoEvPnH4zJPXv
kb65yQbX7Eu8sJteKIdbjEz9dQhr7F6/CFqmL4Ke1FaBfbL654uKjIiYxYfjjdTv
j020t54ywYT4iR9gFAcYTNkHlWM53iIuHOJdm5isd7jpotXHYXYlqU/Zm/xjEQEf
kgRTxvWu1M138kdDi3C4OXIpjiN8Tl5bozD+Y2SUdFzYBYMFE3gge8KiQQ46mtF2
5oMEqzJdhWGKuGIZVGnIe3SyvBr1CXt4+fqCIu8c6yO4qvEKZ4Y33PqwML0I25eY
ZIEisaCohFT13BrM2kZkKQ==
`protect END_PROTECTED
