`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/sQSxpAuyV7iTjOaWVPUXn1mUKiMAHS/CBzmcTxBe7scYfqLFi6PJYf92ScJQbDS
a/bhFxak7NNqvY9oiW51st4eL3uSoIslP+AEWyABBoL5oMwCwc6JlLornwTb/vvX
YxzR8UtHmuIeBl3cHZRQTQmEo1CONERYmsHClmPu601Tvt/UaP1NH8/e1HyY4/7z
eRukdhunzVN0g1GrLZyY/z5iUHOPLey2FAXms2sIuSG7+LtwAvVZhzvvXlBp66Uu
IyYnESx01Tv65yh/79O9lyWVzRsVF+JVnfuvgL1bIzOqrph8qzoWymeNxHIqSElg
spo3v+jXqLl1bvOBaOHRNz68qt8q2KJtuH9UpcBqRxKzqRviPjJZbaJQSA37ZbNM
/yhPT+RrVjUqjD1ZTHmNWWqfsIjBHUu8QoFP6Z0IkwtUIr00/TjMammbzravgQfv
4lePSRFreS39eHEMAYVg9wC8MWsGDRDfwke/wKhk2f8m6y5uACqJXU1yH0pNrP7g
Q2UK7AhuZFGh7ROEp0sBzAeJ3pXKJZH5IdT7SSxzumRE0WXOHMkDHRAHtNzzxgt1
8AyJ0muHMVtbXv8qoBkDQbSsFQQo5QI4dMCW5YTU0WImFqGCjJQ0Yr8wfxEfO1Dw
WJ8iOAn/T3/P2jsyazSyks78phlhlUj9DyQxRfBkUpnGKvSdolWAmScNv9O2W25I
MqciwCB30FTmLOOq4ECzTVKElZOKAMkpwJ/PxSH5rKsh7Xkz3P6X3L7OtDmbO0sF
AZf6Bdh5X+Y7NYCk42KYJNjT9uLZo/Ezz3RlJ8fLkmW5BvSPWnIOKxX0K12c4Fo8
W4jfbeVErBWDvkOn+mKtVAxvNu9DHKlILfvUNg8Vdi1ZudZx2R6uwCGGkJmm/GSO
6FzVtm3oNvP+39ODpgyOuEE7wkttV5qvtGWL/Si4ImOCQQUfwGc5dsOe71wPATVW
iRM9ZeBYb2MjsoKvUbGZXkwjbL2kVQKXbr2pKaTU+eEFLgN/1Cb0Ev6KlGA30DAD
yOXYBPSFgrGDny+A8CEtUPGgIyo1bDkr218qvxsg+9TIZexmCF36iis4QNnmds6O
yzWkdpZ6pQ84em8SmN9cTCUZcOj2hTVhHE+6W4u6o5BfV+R+1Vte2nC13Ygdbfsf
G5iC63OsthR2CrOs3rglmNFoLEtW/r21amvq6RUyQiOd17p96tOc6LPeKa8sQ4+I
VfN8cJ9lk/y06DtMJVzYn/ezITCbRyfULh7Bm4Tv8MTCaR81rasGHURv4+3XpBu3
pHNUTz13jc2mr86eZAHyAe5S4/jK3SqJzb+zx4XgSjP7SCXEm8i7Uis4mmS56j7e
yhva0WjJDdpcrjFmL9xLBoIvW49YV0x9Pjv8v5/3vKAIQmiz/Yq/Yfu3mP/NpD9e
5RWBLVF3IDxKgVIeme1HZXaDZVjUgeBnyWMV5A/Ces8LLqvYUho2KEaUGIp+i5qW
nVg+mB2JNN8zC//drEQN5LBlvyln2U+QgsASBq/m0nLAQBELNU5IkWuZQujc34nX
UZalEXEfdjNNfXVyq6iOucFb2sF1B7QWfwH8EXFHkXQxY8eTj3ARKiT8YaToSqyM
yowsNshYRvHZc3CJnDIegolsDQzf128ky23czMGn6pf181Wb94LzTGMkjARfzY4m
2RAQ18VeYBEi4rSSbKZmQHXSoiiwZo/1w3Elkuejsa1HNx0BOMxPA+JX8oBt4vFf
zdG7ruWQPmRCDsfAK1ZntwAt8X+8+VC/eiKvYdXQ4Iikkk74DO9DtIV2sDdq8Qdz
gyhklVab8FK+U9aFmHMCvyPEByCjQ9tvKAoTOhtz4N1l5x2X2oZlWU6AJb7XRRBo
r4yE3hXE9n67++Px1503Q3IsWgkMPH7x5yjzOO2M2Vx11jyNL7+ZwVSMaEThp4QI
CHrOUj8JlLvne6OJoMr41taug5phP8EvARzc2RRX7BvXIEP1/0/ASDmxKJnEpWjv
6whbcymySYwJ/tlWZFPDJp9oJbWPGInMzvVoTtL72eefaV974V+wUWXKMNcfC9mc
YR2AILNH5FCPFbF4ZO+1iQUMTEItKXq+deh6xA8/tGPX0EG8lrDI4guJlv05rV7C
7pXApWdEPKxcN7E9MYachi8cNRyKTgpM2k0it1zToGdUzI568jKkce6iFvQFGdo5
mEZiac63jxah+dl0abD0EWyn1KkL+6m/yiEJu69meOgV3hmfBe8ihIHekiLEpO+6
xXpDMAjhNc8s/70SpFiFLvdBILUm9yYbc/kqNScebcMGjORfPMdBx8zvZLuhQP8y
epQLP16jqIrKnyyoSv05QPpoIOhSNw+F/6LbQ3mEdnG7cFXVq2Fiqncyx+LzXsC8
bQ9XN4CneEwNDx7zyuwtJGByOarOREpS4ncBBNK4XB2ou/iD5vIekMB5Z2T/pu6G
cErBLxUr7VOnlLBmpXIHSy004fM0vR7GXHFSI+5x8o2XIc21+cNSqKColcSbPFB1
g3LMl0t/4TWhqdSSsPWC3N3ml5m4Etq+Vh66wzk04euehcz+gSjK2io7OHAxrY2y
nyYhL3hx2T29tAsz9hFcrpNYkvoyfz+V/NgSWKtKwARhUIJDgWGxdCS09cli/WLp
k669JPiI3KhhM5AXmJI1MaXSG6X1iOTDGsGPwDdpxE++CR+Vla5a6Kcik0PD+45E
3pooi9OmqnDyV3juUl0Nf9kJiAhIh8bLGe5ktQTq45rwerC4DU8RGRqbu8tfxyr6
kRt7FU5Xlmov6FDU4bpFjUbI4J0TMktas9vCpkaXYqpeicaEs6Qc/33LlZieIkI0
23ZltNCCzT1n0txiBIKLyzfm0DYvw1z3Wz++hmfJH+52ezssXtcw7Me/KVcxYTUd
S1lTlQmWdAvO5EajD4U3dpHaBWN9a2sXN498c5pgp+FZ7yNuRHnZEjRLO/yGqFT2
VRNYnk13B710K9LNOC+fwxoZDDXS3L+q+x3bzxo5jxHfCoKP1DktPLYqMkHh/VgO
ErgCB5DUlywD9TO3ZmSFUxGtAnjNs88RPZ9dBscL1AO6F5ufY7Rf75IRjx2cPlLi
ydy3DBWJX3rBh1zueKTK+H5k8DXyCDHgip37s0gmiMuidlJ0hza6OYGPi2Gw/1lp
GBtXMAJg5UK+l9cZJ8s47Yk+KEGddK/Jyhnmz/A0/vhsAIlz/SioVKdCM7JZluNS
Enhk60hN+yfdh1bTYjOIQ07Btic2oNMoLnRMqmp1/8sXgDorFtmVhsEUujMWFquw
wUHssmV46QrRDhXABe4dhFc6+Kyxg1B4/Hg5NH8QPznQm8ynYrj31UkoagNOJmWI
U1NOAXvqFNwVfuJGk+ESVDBvPY1CSl1RKZTkqkg8Q4m0OVfS+EwL2wKm0zcsA1A8
oghMh8gBYmoWUFZ8gTa/Mb17PG7r+DBfToo5RJDL/pUcsfRE8ucbguNLWyiev60z
FfxZYlfN6yP8EvL3cdmeayZ6x1SnpJelQ4eu1UDaIWrMg4wlFngd7P3wSUHwKBTi
6GVZ2upelvetMS5JT6UBeJdGvi4gzjEwZitDG4NQ5cPd+z7JLHsN0L43ScmTU9gm
r8pCXLPcWz79wjB+0O/ZSLQslpCOZK19D+vz2e7s6jopCvbNezN3VUQuoZiB7gHg
`protect END_PROTECTED
