`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/EUvsZBMJUMXF8chr3eKE8mTYxjEuhO5Q4is3BBJqYpdTEXWVt9vfN5jqhCQZYQ
UG21EmlBhK5dMX7Q+gG/X2aRtIdJ6qgAuOS0fY+hCZqnxzeO4iG4O4eHNIyCIqoa
PMINgNsKPdTC+6lL7NPbZQ38iXBlhf7tkrjjW4lk/s9R3sImLojuj5vydC9vgE9e
cx5KLJnLEO7LcANs7WDA0tFgXY3DCbblGcMPjomTXzNBmgUNAtYcwcjijeS4toUF
Dj5640l0n4Q95swwqkPK0Te/9D4Gp7KtVqsrHUkNO6HNsmAVqDe2zEAcNOZoTMzk
VYh0W+JqQ8HFy/PxS05cOVzYpdssFlx6qdlHkuUMROjvNw7vTH8cwY1afqccpFUb
vvYP/0b255CT4Jw5yyxFLDwl5GXCm74Of6tc1lJFA23YK7k+1pvNcGCHgb/H3/LW
gDdARQubOxAT1u1wFCp36Ix+0dbnASH8GnnPMSlJ9y6VqVHTMVJaY/Nccnh4TXhT
BFadAi+XT3dYwPHmmbtq5dzsCbROMStL51XaelT0UBTNbPK/7x1e8jGSzhfgueJz
NNDREiWr2J6wLdkbmyfcDdXhaxD9nD5j4aD5eIy1R0nGKFT7ZbDHZgCUOO2A6hw+
PdOw07ggbS/dHeRRKR3HB5s2u0ZdNzSsYEG1/k0ahZTnCxejy0Ag/bpoMR0UCLT4
5+Im3Rvmgf/skVEQqLWqtXxePvLC1zgQSc/LF8Bu914xnKMa2AFoAFikwiDRUVPx
UbFId7FqBRBlU3kpx6RjgbecxYWzXPf5CfYEepWiubQNidjDFNIiYcSmb9VEz84b
EU+ZAk9JNgghYfoFARI9WjRwEjEGbI5U0a10yktAc69nqfg1TOd7ULtetCdMTzmd
unW1BkCJacxXAiymM/YGvVJcmWjfP9Gaa0ZhAUb1LKBUp4ADdryhjuQVoi8OF0YD
4Axajwu3QTV3j5x81hlvM3QK+GFQOZf97SV8xjv0ZhaDDEmVFltD5KHP+P7vjsLZ
v5yqZ2c+dTxoRYNPxM6hty5zZhW0kbTlEDi+EIDJcejg6kg33Bi53DxeNacunIGW
TlyZ4zA+zuehqluofrxR3n8Mgs31MidWNzVsDOrkayPaXRKSQ186PpVxvq10FqOd
Xbtaud8uxtSlIWSnEFWDgRYx0QcsYPXBeu1mvYS+PH/RtKPYoRsOiR3bxjCFaREz
jV5BbnMuZ8tYxka3qBYcF95XWx2LbLuu0vPOErcmXi+CHRKIxAP1INXzjOxuwQRL
5xv50Z74cjfp0+1b01Ec45Xs6TQQQUICKq63jIVpxPIuEN4oc6NuZj/dSOOw5wx9
2wriqg/6LtY2BmH4Xz9Q9s1WMKfNkvi3auDx4ssUjg8wGz4KGVQZYr54tP0NLJ4c
j3BIyvvj9DArhq2e6kWY4LAxp8sW/5OAs6079Yc5KaWRGNkV0TDjODQY4/SEq4RF
SK6j3Py5YkzRQMysfnMjm3Q0Re/e0ovqQy3qoZ8edFH7tloBgf5LaPQg3GtkqK31
1rb3uToIckji3i5yWumQcB+lZAwTT9jYVa36twSPcm1VPBaEfo4sKDqcaA1s7Yum
lKkTEAhhZ0M7m/U0PqH10t2KoaxdOCytaICwTPeT2gkauoF7qkjIPV9rNXGsXEQ2
dWDEGq0w3ZHYIDlpauJqN1jIdqyEaBj3gTLxHNIyenFokFieH/JsUtOYSxlHxo+4
nmJpPU6xy43q5n8vPvRmDlXVLS9ny+blzAk7I1d4llVIDh1uXo5qHtCgw5oAPpdi
piOArTWSMlYz2XQEnpbqLx+0jckwtel2534h0z8l9OFQV2wqfBnGTV9cKcFaHHvQ
c/zDI3MOK6ZWHbfRNkBXnBy7MqrSgnoOxyOSvogGLVrxJRO8dYD3UohO52fwRksT
tjHHx521zMNJI2O4373GddfVhPDAJYyi+cVuZ7kCTIsgj44rncffmAmA2tRDcgBj
3K0lKhqOm14oGZYf7XFEiFQ0OkkeAFrQ/FZl6h4W6pmwz50Ai3msp1Use6X2zGeF
Alqh6i+fUg0pm6Te+OapgJdGzOL4xUhxTdaL7+xVIl+iVXQsAvxGA77ApMqWQVKc
49AtqH4xhvtcKlJcfQM7D4x3JmIJjjoGrICJvNoHSD7N6BAp1Rm5ZDRjrrOjwUkO
Sa/LLWGFFBdIKQcSpVoMNe818I6vZoxJZ6Id1mMFLcgX8z8K/lxOH2nCaAsWcKmX
pk1cGrPd6ypFuJCp4kksg4dlpQuthDo42v7xsUNE84lQKLSmz7cK3wfNGx7Q7wAO
WRqn0ODpf8SW1+nC2G6F789/7NNCEpFoeiqqymBlr3sLitNr2S+oQ9i9TcyhTf3N
vnAFnq9n54zNQ24YoZhTeGtEypsbxY9vvyUYqwhcivMEbs9crz55mNSDqhVi8DrZ
rA8SF/SHSLmB6ETbRXsSQMjySFfhXuFmaQU0z+O7X+xW5lmMkm+fmo0PhcYcxL/l
EN2QqHC1HXxbP/5b8Sic7J3JA2KjPBolUPhm0MT05i6XiV0v5WK7MgjBD5zI9fKu
geGC9J9fhbVvcd6C02nC3syOczKjvG+9HPk/4cf0e0fAeO9AiC499pWCrgLR6rCD
949JG94PdnQs4dpZuADIRUXlE8+0NN8wwg219lUBAAXnZjR8Rz3oTh8mCk/JUxWY
kl5TLpsFTtrw/P/BUnCxNCNKN32Y5mLyC1N62esO2zIbBonjQC0w2pAF61AfKl+z
g2mI0Yx1O2nPISbevuI4bnriV+GiZnb/7EqFpFfCuXEbnxQg8qSuwcQRzUpCxgDp
jHzcjAN/4I8ry9HrAIUkTBx7HdzRDv6VE0iDibmqoJiJOuqwYaO+ZfAj2tp3A4Qn
DJntUlhWPNyUxcgI+WrzdPh6S9I8YR6yE82HNt6W0nZmBXkBCkbK73jOsaeQRP7V
xs+785KUvZbxJBuYDp+FGMo8/iYbXGVdCTS8dUAHoHjI6KGLqy1XeN90HhpIc2EA
z+AkUgpO2sgHOGYk+gmW5TIF8CLoy5H85zDqiRl0+EXkUGr+zvBbNYfX+uUZS74x
JnzuyvRc0f7DS6Rbqu0mCvKnqDUVW5Zq1UvTbNL2i5+v//pjU5vIH6CHQ5LXNsYn
Kaf/YXM+3U+LNF6Nsyq+0YF/AI8q4Ubidpky9lCKTlsX5MfA7kotXjaGBxatoAKm
8mvDPKWcoO0SFaGN71KUc4B/d+ANRZY/L8ofo9QePkHDhls+HzoA+ADAs6UxFo/W
6G1QMIO8X1QxrATOh7FprSFdo+8dYDa6/j2wNPEmOxLpwEZKZsEu+y8nvV8HTrnM
MtKJE5tkESpOYVaEzN257DVOWR31S8BcyQb2P5YMxN4MC6NoI9E4FqPBc8edthLp
WQLcGKIQuFmyFPNNcZXLTOnMQEwuCdz468a0KBLeVSVEqVLsZNDtB0Uk4pPw3CRF
Rw5/c9smURgIzpm2Oa4hNBg0mPSBaF4hc7vQrr9oDAbSP5J2i4nQSKS8XjAOB2s/
gjPFCw4WHlTrpyNcw0Q+FRofijLaTMCyGSO0SKYl4wGC7VUDhcCTtj2QAggsDRUE
z1FlvyiL9gyZALhoysMM5wy/4oDtdcHX2F+7RNEmCfI0yZLC0SLQtKHgOp+ZDA0F
FRTnKYTGHDzWMe8EVM4RKG4rDEfksMSY2NkoNLqPeLCDCrgm6HhNOHKm+sKedwhP
CLHxGpnR10VivTWraUWzgF+x8H94mWrJPP0qlV+DOW5GNpRC1vdYHXjH6QgB1FCp
n0HehjE754v83QIO3/TIT58Pu1GNC0hHVzDhvuRmkUsiR7SvuwifG5OHWrLqsFia
YfhIWvuxe6M/OnGWOJKXcpPvAsVn+wximFqzdT6UtuZB7+7U2b2DwzbIWH6UHoYH
q2nwUXT4Nlj7wUVqJeqX/fv63pnDsT7rUUv4sbtGJ03Jq+vji59pWVGl8vOvk2Aq
o9CX0YHPC1a7EYIlpxR0My/8Ogq+LtJvkXNYqkzqp5GPcS98NJRpGj0mxBY4wfit
d4PfpsZMp/rOELJCVqkj/oWPBN/bKvrDQw4Llf7Sm9IaO3orjWBQHwDKaG9ugvkK
sy4ImdV/KQlMuCvWFr2G7jXdtUnQeCyAJE10Ht0c/5A9+oKvZV8PaHncbpKWxF0P
iDrBIlL8wI1tUlBbd2u+iRPRSfris1KYz7Noz0hyYDq8moQgvYNV1g2gHhfzAavx
0fzWaBHWxsyUUsicJ4fBI9jbGht+9W4n4jKFIFB8GF09CgxPsZ34VDfcppYa/Uk2
Hp8Exsr1jWS8MFQsWG7l1Eo2+Bt0Zhv98dnLWN6TNefS1q5khgx2kpyVgvnFjiCI
MCkPeKfjLMtHPd0pBLHY3d0UHWYLsHG1iuGlFAWA3EgLOqeTorKqVYFUv9tCvmtQ
aHz5h8iv4s/aj46eJcDHF0E1lm28WCgKl2/7q3mtJP3+eovWLk65D1ocK3Hb9sec
OLQYbC6k1r1twl4I2WkibSXTJ962oUplKSaaOKv/TOlqQsYrRqGB/Nek62qvEP0U
xG9CbhGgzVYOEcrkixpNqYxlUSu8nGt4/z/Xxv3ieCr7zt3mcECvkiZrJ9+/ZIEn
XfbZAqLixYohP8Pl2Z5/IKDhhMt7eWpXf8WEVOtG+76vqkitDTd9+nOD+MGs8bGg
XtG8SFbl0Zxnf2KUGwBZ0urJOaY6WgDao/utFI8v0oXK7gmBSLqZoEg87lMjEmtk
LoSad09MJjURL2vWBl1kSJpYtYF9X1UPIURtm4bCDSUy3sgj7RfAEfyrDpetA2PC
MEv0PbTG9UPP5enC5UpU75HAKufTOL0QXtVLXg1BpSgw3T6GSkH+Za+cJMZ83Vj2
EdY2S2fXnVS+EZ11d4FPi47nmXqk/UMX78A+5COEPgoHYKQaCZuZxED6Ak0CDWih
8n0yxLge5RayyPobZIqHQLC70MTU89PqMvlRUy0pToI9XTPP78YBEbv0/SoVeHRf
UbQaSpPRjEHDRVqisVSFcXMBe2Mvegjflbn/yWfzB+2EuDCTp6gPboW98JKfP6Nu
nKO2fDtind401FG4AEpJQdcCU6AeV25DfLYoRMQJQIrQ5cTM61lOGKLVT8kwfJro
CZED1yr0uGXolgFwvvkxiZoMSp1v4IGUNr2gML1Kioo38nOaOlHgD8ROTMcxphxA
+2fsbrJdn+RN987OwIclK8ZxR2qtx8XKrGCMxAmvSpQVva+Ch+hKUViAQApz05Cv
jIK6U/42ICSFHoE0y4G1ilmv9vFvjh4cuzey/HilFuXa5TBSg9Id7sCB6ofB8jRZ
8xI1a6V/MhMxQo/gA1Auyv48/fmYGkb/Qz99vangwcnTIJkCbS6/acdwopexI16n
3APZd1apAe+oEzS0R4qSTBXSR+P0wo+e2jAdeZjybJDyx6w7jRToDHFo5m4pdJb0
WyszHoxEQtEZm43Blj1XaeYHqqOoll1LAZSIZ8mNf53iK83s5CvXXGxGEXeT/y/F
p+eNONZvAZRlBeUppxuiELbkdVDzgwQ9M7iqsaDTDPLCalHZEUZReSLA46MBCXsb
L56P9o6ph8XbtBx9JpjL/lceCG9ZRvYOuXjN8iPSmY8vWwu2AvoBL/Jv69xQuA8B
hHb63WbJeCHp+maWo0kQ8iSMwWpfvP8Jg3HM0Lgp/YK0GD0BDpOrfI4HAOa3Cz34
vkKmbcKPK4m6MGrKf4XQ62VTd/wZLo281Rbr3hqzUHYEdXhcE8aF7RpZLQmgMmOt
Bi+nGZURchlS/V7YuAuv0EJ1BPvVSr6xinvwPJnV50u3rFQS43z4ZrtfEe1DJ7Jv
HLsn9sMUxzx7HJNtsqmyGM4r8XnISR6L0SCCGcPcWixjF4ETo4JbWmE2QEoVu+L1
y5j4ibahR+ElTGmCnTeN3zFTgiO83s5iBSnfIgPzah3NfTiRt2n+/AQ9mHax/orF
dw182WMEbZl+1dOOqEJZXnuf3Am9jh5wXndVmgKDZXX2jtvVL7FsQ+okfLQIv7vT
7f4YrhjN4HEr7YDgPHAOeLTiXlggv5OTKSYlyMx8Td+Q3XsMbyHiXTWZl+68EZCe
KsbHZWDi5NmYDh/v3L8hbrkIVwfqb1z15VZBgxDwiAoai1qx7xIaRxjwZSg+L+Sb
p2NgH/ccp+Xivnjha1CCD28mp0pOyCAAgHBRXANfKBWr5a8Gvakb10Vh8+/s5R8g
DUiYMTFBPBAp12GLm/OHt6sMlJbFNRdZIQX3LJL3+VHs/Tsug4QY2/UbnCVcMuKY
CcXBtwR1jDwa09pnCVDWoW321++GlGF+nmCD2zjFhhXp29mgthpHXU8igg9Bro7B
rFGclqrw/655OB/8zSNxvsqHu1qnKY/i10d3lf//0oz40X24/ZkmnDORvOiLmIvF
zmSk7B5WFpU9QYYLyulhTmadpLte2hPPo+olwrJk1mQJc9V4sEywgiah7sqBZQ6O
Ty6W9soAOb9FMYGzVvs9kDHCu4QWumudZumdXsHF9BU2kcXeduRW6obiOMPwfYaO
54QnMF7EXGKTBzPfKukXiTn433AcFa3j20cg1Lfggj21WBwD1XU3OCPnGohSfW9U
3DWgkI3rAB4AfOATMPQtstnT8ttaYsid+lcbWQP3CxQOTv3OMgaPwT2v28e2FsxG
f85ORolwM46wRSlrZrMpkQYOmrjKnuCcPhZoKjDI9ULISF319gk472QuHqAy001R
iZFOoRdaQWh7qMS7N35IxtQzvLG8eqqFVPMfaz5clx7m/cjzanxNoppWrUF0ex63
sGzkt3chky30W70g6UAUy+gEzfNNg0+JLjn+mDtiuD4Ona5E1xZ0bnOQVbwM1hTs
6CQY4XmVbIszijE4eMamparJYgNsbgmQr8eODw5f9pOaSvOdEjiz6Zb8znThrVfd
bDhj5rTrJYm8c9+1tRFLDcLvlwAQ8zIecm80uBT3s+0cAhKcH7EeIqIKcNnV16Fs
qC4IuU+/eRABF9dd4hizEHy0Wf1GcnFzL4ybYjMgxg37YsHoS064AuQVl3TncRgU
QESQwJsxNP21HlQeRBfVPwiGXWvB43I4wDCyCi3HGOvdXV+o1gLm+xQKZ7FoKNrZ
2SkkDmbK0vV9/A8xh4lQRz+0r5xrCV3B+R4zeLu9eZgROmK5pRnZ8qKBTGLoiT2y
dZwR+h64/b3LcEcv8H/dUjYxB3qja1jQeYDip0qVAHTJf0L7jfhaoEeq5Xnlx1JF
ttNvlH8CRcO8cUsjBKl4pRjsTayFYlLJHKYrkk29YVGo2veMD5IBPgyZPbqnnUBm
yUV3SxGWCYC2JGCbIbfaqdd5hXGYx1OCytKV44BDrID3Mq8csoSO1Lmzf2mmzhSH
PPcXtRzySNk1GnWVPj21KMBieM6vMEwSxjqLaCuoJDYcQ/8AnPy2RTx5TuFWMkhU
Sj6DDeefZJ7yqUAXB0J6YgYOfMpE0MI8QMPfVX0RFoaSVaR0xmsBFqGk3BK4bhwa
pfFWuw58YB1EzKJRsqlhIfFo4/9r0yCEfiOe9RGqFOPLGTgmdZ2xMTG49MDh9GRg
qwsZfYsPxtMHhwi51/OpfqwYc43JZ02Lvj2xUZM+7gJyvxFUBAfPNwhQd/7cqBbz
INpLqfOCP/SqF8oM+USKFrZp1twE8vTZI9fo8Ua2GBoqBBjte5p1ioBCUQZvtlJ4
O96w+umKsuwx3FFZld70fNpNfMiQ09Yd+Dydzrmu9FfThceyQnMi3bEiijDSgyuK
phLCHqaqzP/TkGJ3i/whoAkmKxY1qxXfYkJ04o2buCH6WCe9BUogKNnoNW5UEXQ2
eowr3zow4ELLZWycad87sJrZflt70oPPkJK5NxwKiiFD5bsaFgZ+Z7XP4kGWJFT5
fgK8dnIJ4DDacvJPepql6+3XS9BJF3OI99mqABI42T56BeyTbIA+TEDecTBbA63z
kiVMveUjW6SOvApnL/FJt+HVZ1lqCk8NCcX0WJqJ54kR7xZsDQrdYRZjgO/yrrwF
HA6gEnWD/Kyqx+YRuTE2wwylRWvkgDIZZTNzpNfnveJ1Mi44nmxEwv8I+CCAgQta
e51VMfh1yPxSpk1l7Ap6kRfeD5Ly3zgkenZio+Wj/dQvmt6h9TKhevwykUuMLt4n
Pzh/PXd6KP07D82yEQ60QPMBXcoho795qvTRQOf3uM6Z7pv3dHzIGDr/MnCObLpc
Kx0n+HxsJuyTQ2JH95fIHl5eAtsiA45b1wKVS4bDz7HcqdnBH98U9jEmFr2M9+2O
0xjXryivdqIQ6MXWCv69NYk45FqtkarBFa6BgMITbgLoWtrwwH2ItWkX8OqGvweS
cGldEXg8wd/2Bqo2cvAzhYb11f45phbeyRkWC+7vM1QkZDFwAmLoNhB8TDQi6A8n
48KZfj7p6q6V7jE3D8LQhZEFSgnOoCO7yWFRZk5g2thtgucmGU989wlO6tFUIKjo
+2QaMbdol0zFL4dWFTrw8fRmfQHgfb+tV3GqC38PZ++D9dZKiAzgktwko4Ge2bp/
rerSzmYKJiM15HH+2qFAgsWX+lhKV3gFAiF+dYE4WTmxwEFllZ9E9JuVwBoCTZkV
tZ2d/U6H5YXgWbGKB/A72w1UU/1GzMudxt1zECdbV6L4ATwun8O2jfX2gM6ezriX
YTN/ki+8kqKF94hVKUaBU396jMRhwzU1VzV90Ko5fnJ5pWcvokCHe3OLk85ly3BR
//j9ck1ga35ZwSue3S2G3J30s+A+bXW/9bvBhGUR1BOGAj0CEGJWblBbbwa9JKuQ
6DPtn1eOMsei40TBM4paq49tyaaIQ+1C0N64fttYvXGze/SABC0de8J9XgxkHPQK
GMZs2XAJxggFwheoarqw9X/Gd+krtB5TkzVJg1/gjtD4LTbJTWbJgftzq7LOm8xG
DTBoEsCbsKFqFskTLQcGfvW3kIMvxtXvfKpW80zzudolrdX7+tqIS9u+TMTJr0V4
vuP2lFvoifCK58yQj3uaUUskdlWZbCeJqQyHnkyT9oExdjzWb47iHObKwKNKTE6V
RrtrYZACPWDgZGmQfNqfQDgHBwm3h5dkSFjevUg/OK1yjMrEi5jwFQhCyrt/Ml0Y
3SHIzYyGzrXD3cAJsyKCZnZwGq7o8/biRrqMD5DllqV27QiqADAi2z5h1EgA/R+T
E+RZrwfIDfdx0py1o353h5isPIkXrTNUAtIItrOLQSeMrM9ZZrZZSBcumxt9VC/a
qymtkIueU66YMqynnF0nOT9H7+Eupo8fTzvELFWCRdo/PWz2/KrXiap/1alVUgh3
2/20Xfr7ePoWupbV220i2xwhwg7wqrY1kYX9XBM9EOcQqj+SP4WYN2Zrkwf0L3jg
v7xvzFzbWYAp6yIi/Aj8+4t/COMNPDOEGOSEfSL9S4OUEGxnE8PWUhYrjVKu3oRn
y4WQC4up5Al07F3tE08vsehtVy8+LCofGUj36eGh9MzF60oQnWTbPzU+QfhUWJk0
ZprkILWwIvrleL7kBaMSEKuKAfo0wSJ0Kz2FVLj7AaAyOBe1i2pdTrIrLKzzEbjt
xCHoj5YqxxHOORXmqmdTUXPSfuB8GRahAYX5KNfY2dQccesynuHtKiqp3fpgpg+w
BrpFN3y984U+/EWpGRmBynShApLrX+qiMrgrBp9R4INI8zgAZ3XEBkSPGxe3m8G0
i3mRTu7RrT7U2mthrIFH4qNV4MbVEYg2QXzkQMAB4ombMoy5USBLDDLMJzep0ZI4
f1tca3/gDhry62TYcBcVlgJBoTSPExMDd3ZdEssjuZ/4rNOgMjXC52P40PI9Iaqu
0NqIN6e3UzoA/aDlTv/3TQacKVKAYjwQJZQM6N+6slsJDWwTAbFYOoMl2Hi+Gj9t
03Ofz0NjxHJ3JuddMjIk17mr2sgMn6zp2kzA+04iYx4KCUOGFiub26WnXXk9dSw7
ew//zUl1WLxx7Wq7jS1BriWNwsnnBE5Bb1brd4qaFejbrvkav1TszEr9BfarvIT/
0C7t0JxvaA8yyRJcqOB7gimiGHaujXLOg8gWYdysTvyhkJyPjMHR8O9M8w0nDyjF
OUa3nwQ4gOAMmfxiHbx0MiVRut33BI0q0nW/8JjjJW5jYC98s9DhUo7Sk7Lw/tGJ
S04iZp4aaMPb0Zi5nPCiZsyNRCoXfFk2MP1cKV++z5CnYx5RVBc/VGzPxzjdr77E
ZSSTkGFILHh0dnFfGlIGmjGe9v+cb5UwZeCG+gGBy2ZL7Ux6PQMprnwVvk+12cij
B9vyvAaqNh3PNL7UhzYwz2U1pjAQi93NhEykmx6nAsFaojmQPbTM4TIauFAS6zCf
fP8ocj2eyyjqUXLTsw7mvVI2ikLKjE5/MLlxXrwHXTU3g+juu6sQgWZ4Rpqmvemx
4PdRZlcvKoV6vR7/lY3lb5dL2NtjrMet+GVPJMxdMCHVYk2Y8tYWbM/tPzagvfJ4
+29QYE7EbiGuEgi2OZSIFh776CuOldZnOOs7+2WmLnh/UdPRK3p7H0I5lIZHaT4a
MCybYCxNpAFkUXNew9bBVz3LbV9eFBFC3y7Ux181NBX4S5w7HhPjl+iWrlNvZfGT
ZzS924w/dviONR3UqObHXI79FRaqhIoexcQd1L2BDwQ7+JTHD18/KCEjqRuvS8w/
J7mGhh0JZJbaVGs+axqnDj1Itetr6/kdwRfUi4cDfFInrgR656A5GRA68aoZFViZ
eTJ9dloY4l+wkkh6Wc5Ys8dkh+Q761RL8YXaudvZwg78VSGr1W8RX3k2pRL3FhHa
HiIM64Rz6WgRthCdFDtRc0UO7cj/OhbxOycQRSZRhgj4mw27SJuQUVWXAMfmE1Es
+m6YA35K5GAY6/+BWNWGMJzfbtqom/qF95EBwtOBp0LBxqRFmiRr1i5NV6nq4Gir
9/W/FlYVldApQI54NYaTf5QwKt43mEmEC3fw17o5JRc6FMuI8Grv1GSSv8zkUAO4
vioSi90R+pzpk7ZJveF4ciIJRpjDuAmWuLqelIK9CfuqWtEQZJMglTOJbx5naNWW
0SSON9hHMi6gRsxQm2uzcfHSssOIvw17VfEucCL4LV4e9kbKwLoZzkvoLATLt6gT
+Td7uqHBXBRa0B2SF4n/1mmL8g+70RTCntOJ66FqsBFhmo/fJz932IeSoF/7owHx
dcLTjCleTNlj5Xe1oAgMNPhQJuSHVoBTyoJ214chqitzaMKHYmZyPIO8pt6foipY
sGXF244Zzc8DxIu6xbwJWfvuD1vu8Q4j7TfxWTDI1AaPqgmCaKf3WJQjHBBfaVAF
gwEQJF9grabn9alpYVoyO3tZ8kuuTbza89RIK8h5TgMJVR4y1MwFDaM6HV6KTh9v
RYuoObu4zMtdJ3gUUhl9CdRWALQue41MJbRIAtx+0FuhEvzSgj1pBPVcIuauKQwD
M1a1hKcbi7yvFjJ5rg04DGKXHNbtTB+34OawKbMsLK6TfglVuqObm7hIHTfFGkcA
pLweACgTG4yQiF6jKkbRR9SAxahzL8TReVFAGznlSkKTroG7YDvippCKytbuv0O3
HiJt+6EgVvECoJuIlo43r8JbpB75j61crFOrzqw79QP8MqF111FKeXlxJMD+F9yt
pTTsCFl2b+qs+txAHWNbKs+ndtTgZPGECTpVA3yXjdQI2v9DrBTGcBHwAd2bUYms
MUNcl2aiW8+dtg2u6znG9Y2geXNirbJsrpxKeRPbipa28Me53RBzn7fxwX4jPgqE
bobunvgZM88O01G95CGSlIp1Y6yXuCe3N2QxxU2bNUE0V//ylDxv2GKimgypCPsn
PyHM4WP3UOs6IvNf/m1HEPzxxfC9Huw9WJWz3TiYCDy7UPVqOZmm15NsJqMeB/+r
JbIwLCsIqpB+6ibi5gZG5Dl7o/4uKwZrSwzC/06OUwnjbS8t+tT4a5KMxm6/kEsm
K4d6PXZABLmrxD5APUzdlvpE3yaD//7XOEK0y4QTEcoxCwzvm5HpvuBQzPG2o5sU
QXOFFrWimNtR56Hhb+FSPBRwrOYX5Ed/9Bx88Ct4dfftu6vKz18SMxz8seiuLvEN
i4kNH+WZuq9NbHYn/DMbwOeGrriqQf9CONII53LGBw0Ig9tEAi3FnmrbXNLMGlpn
8XdYygrRpSM+9xysaxJ1Bo2obO5qJQse9+Ac7eGWLc0cxsH61NjO/avBIu4I6NR1
zgICxXzt53ZYP3tOw6sVzrORui75TApiI9bvHiwjMcSi3rWcIz/6ufi70YVxUN+d
syj5WqUM8MmqzhO/yikHGD/uTvzmLm85W6sbx5DrbwIN+S2bZXkRC29ls4GsMnv9
NR/Ry84nlEU6lpy21Mq5t366q8KSQmCT2ksL2dL1S4M89oIanMs8Cl9jIdOyO1ux
nl+OTs2q68TRqnj5ndSS4d00hm5PeMdUVBZ5wA1vHFGrq04qmolG+kNxbjalgkHN
q9qpwnNmA+Bdaw+kN2RCd+kVbXYGjrI/pqr0IAC3A0f1Q/PiIK5SwIjqW3KX2uUy
2P7JYW+Kknjbd5ee9X3x7+da4K/dj6QSM2VvTZjR28aso5Pr1+PikrczXqOq6ZbP
TZUQoGlOK6XrxLpJ/Ty5p0FN6tut8Mjop+PvMle33zg+1kMF6k5gyy8wqRnNWhIW
ZB8x9dW6bFjj5du+4xbueAB4Kg9lLLZyFHqP7WfjXg7+0sMPdYWkOW7oYk6FSgl0
S0In9DzMLoYQK4xg5khM2AuK2dzgaQNtrPUsVizjwNTEKF0Hq4By7AIPBTQdIROm
1PyGjOTfYZqX0uYayWBO6zJQ/e8fyRIsNdm5C88i9n0nhmCLint4YeFf+H8GEoqA
JDYnHjulBt50y2KuU1LD5NHXOdZe4lMOxTN6rmDn14uK0IJB5rhle8nRFNHqOVU0
hrVhUG6JHroBwNaPR05L+GslX7FlQbNvXMFSnu4K4JmEyhMUK12qqQwmddXW+gGQ
Xdud0X45djUf7eFDYnM+BgKKI2v3MYS7rXhBDcB656w/xxUaMH3CJN7Z0c9bTiZp
uQfA27qWQYrfeIQxqCGjypJa8E7V8vN9c8BGUi79BO+nN4Pv1YIDqquOf8clc4M1
IVtDQnuanhIrIpGNcWHB3lnYqF/0aZT6ouVQ1GgAWQOOSYqKYWwfmWvmuVRZCTsp
kTI+f9QlKXUrwHfnk0JQm5J0oWG9H5Vy16/YCwX42F6EgLHe7YtAnTQI2fDxa4NT
oyT6PyQZRDkHhdXR/nezT0GrF/jp9riXYRyWoemUdKRA+PSrOS23wSLwJWqMg7HY
abYp8SflJnL8+frv9iJ0z9t2H+YsHr5p1xBcuD4bQzHsCBN9Fb6FfvyITqd0nxke
PxNd3xj+LHBlveqy7wjcm+lefFyHK3kXH03nIxxmiMrFxzpm7An2SzI6KNVkjppx
ebEdAcHHEqNhuvigVrD7ypK6DKhH/KkzxZ9MyQj8iB6HCQX8WFqMYwRhhiX+MQts
yvA6Vrxl7RUMY74xukIx7jglW7rHGf3KAh1cH1dnz+07HEZRQUfhUbQvYcFhCEUx
OrBBD+cMNlgQu1WS25Lmew2nWtWgLBMXevDucN5GyhryE6XOeCA/W8CBC+fmtB/R
8nvG1BcoXVU1LzQgi46Bp6NcQnOnjF/usEFNPx3saxHY9NXSaasOud6z305qpbwD
8tp5totgBlQ5wcbWwceezSeXCDu/U/aGuhHLtTR+UcLK0Eb5EvyLmxw5HRQlB3j6
vJ4esQi2Jz6H9fsZq14/92iMmCjSjjPJyIHPoQqgm2BPBvQV0nhPUnlT3/o+R/tp
0fVMAkqEKjH/Mm27GfmWwEcEXLDLxR3jzyaSwAjpmkH3jaZ4ASK7Y0jNdPtVPsSF
wSZTg9GgbIqcl7TBwr/X6ZUAwmwdZgqQwy25Lc6JAhD2SwPTk5FMbbtrsJGixqso
4FAQq02d6W1bzxIYrxm9UjwnNShkxl1CX17dVl7/QPrMQ0uhaQMLohJA+JJmHjYW
XxHAHsI+gmzBjs4l/BPsyAkyMjaUxqIaRHlBlsXbxJlYLJsWgh1I+esD0R0KWaLJ
G2VNrH3xAKb7xgJAE1iDySBgHZ4QuF8NuZaU4G7JE/oA6Nyk06OuCdegCf5AaDdo
xQ9TRzn1wAnpKfRjmrQleGKYzSTjySJxa1OKQ5NnsRHaRGcpZYjkmHzIW/dyU+kp
u/UrUa9ctjasu8OIXLPWpuhayXYe3FZvVQoY7VBG660mpNK5ILfHaU7Xo6vIqM7h
yl7LybMW0Qp9MSGxkJpIxf9u3uK7by3jPvxHTfHgmqGuCJ9a5EnbjhEeih7Cj6KZ
wZ55BdYhlle1eEDgVTmstWYmnLEMew1Mrz2wandMbRW5ZYcX3/JyH3f6sRoyxE13
kv5IamUtxbZSdwASkkuHXHOWcss2rFccF9MBg5ZrbEfxpQTHldcldoxvf/6+ayXa
HIR+D11pTyvpOlPise991A26DrRKK1bD8jdl1kY/ARJ9oeZ5uBSoXXd0tksgVfOK
YWmkcnoeujH814kQfDcCYC7loQWSDxFIzpAUxp+/136splqXD95+oLHCl3IcHQ2W
A36orNQ30WouOvbfGk24VMJEB1WXY5h8o4rubnsWIyoRo9xYKVLEpcQbg7F9JLab
N2qYf9/O7vvSNJQzVlbMC1VL7hdkdYuI7ClxFS0zsrS9A36enPz4BJY7lpLYOoPQ
+ECMcI/2L/31ejR17F7eUQmHTV0XuYjrZt3toN4ChvWEbp8UlZbfXEJJUVhPnrBh
OvRgItPhvw6vvEnGIivuYEcoui0IHHvTbkGQzx5WTWXf4BIJ3gnm6TB0M3PXnvHa
G+c+Zo/eYT38gJebgjyzrST2XX/AJ4/s+KBi8G6itM2wj6kRaNCCpQJv7YGRhxUX
6qbcNOe4GzhgOBVpXxSIjOpY+e274GxTuCEj/nK7o314timVAEAN6QiiSvXVLkeL
zyKBQ+RSYR8GSypWE/ulwdSdgYc2BIWUCzDgorJ/MQ9lO85CKolU8Yfq0e3Wdqnz
cNP7bkU3MxKbCAXhbDljZQEDSBxbQf1L13mPeGyj34RW7zABolWVBY8401j3r8NP
GK8h79EkJcynseaFJqc54hmkuGko5vX8KVd0cVB1RZzW7HVfpqamRdE6O2mm41X8
RIQ0cTwUsmEsjQq5+qTfFr6K0iKDNyrmr+pz7AASpxBHT1ONedXdTER+pgXFixH2
4hrVbgDVIApHxPtu+8Y+j0URhzFCyWsGAf8ZKYOumeMsjPUwHOCC6EvP7cg0lruk
yDqoBpEbvFkmt64uiHLzJ6TnyDldNFyBx3yXwIvz7qO1Seq/Krfo4IKVb9Re4o2n
H+8DmIopzH6xzqASvypSfhlsFcfVtBDoODEGytxEHh+uYHQe0IFYdTM30sMk5oLW
ll6PPV2Fyqh7ref/8oCVl1HjU0OSPHriGNVwlF8RyIOPC+cXjlOHPaAD42+XLxys
iF13FM5h1BR3YuwPmKCL7Gh+ehA6xt27oceMzgnPWULy77tKm/Bwf4KzI8/b0dbW
GJ/DC4XdXadmh0o90zfE3PxPDfRA/S11rtbPuoFsbdyD2j+cYBlh/FWicxekXfBF
gm1fpIMBgC2ZrdbHm2XIxmwt3ZFDRoBOXBOLEpf6PJxwElVo6jYkrPhS3Q+ZzH3r
JIHxM1xs0zZk4hJJGQEqc7U6GtSrBVDhegxKvWp+BB1pg+NodNChKU4PJsJ4YczH
bh5k82m9NoQDABGezct80eunuKFU9fpJ1y1ptLYBgeTy22k32aAytN4eRwOsIeTB
OKBnWIWEXawtfNYx+jbp/GPivj9GXs3cvT0KSamGpu3PchGvlX84/RLmoUV0EhnX
oXedq4TRWzsN4GqMdzD1qnlpF1bJz7sRKz6KpvFO1Cos+BlEvyjHPlBhGlM8sIey
VrI65gakmgPxiMt1PZeRteZWBvo+eU1i46Amem9wYMjSiUGHnnA/dgrXonP1DGVZ
XGEF9ibae6QPtp5tZAahF+LwN53E/Y8E8TAiZY2Tvd2+x1+A7m9ERrErNGdUk/VN
ya+u3obaDKMIQs0oiWrex8F7ZraXcchDFDa2ZxWOkcaXm9DyIl70LXglFegjsxaw
IgBW7awngFcClarKfthka/DhOi9fESocX7hM9GSg0zcleLur2gHNxzkwxMVOTZkf
IFW1mDBO9DcE83qxbEKortSqN0EVmPU5yPTZla6VB5XBUb7e0iey1hYXmH0jB1H7
CXDjl+vYv5NN651JRD1nUNRmjRL09YINIIYnSTVWML9QeXKbDSNspGEn0vNlFTqU
R+jiCQS2j5tr9cfLZCMOejxc9jv9BIoxTwlBk9oAsC4Voqjsi1orr4KSakh6HDou
gEpXSupjs0xRjevclC+bvQkYo6eQxtRRX0TdLbO6VNH0n3ulrFYJp3FIVMnrEIS1
jupQpodEIx3DHGAXO/cQEc4QoHcrcrYD4vSyByysOuD5rnye5Y8tRHHWIuIcC9+0
rPgKZVvXg0654tk5yQ5MGumXYrO6ynERr/K3ZO6ean7wtomVysnWPxVRbEIVEvq8
iv3N5P2qzST5groXPnacXcu+xd1zwsHTshBVg93n6py5hmEBBrhyUjm8pfv7fLGb
h5SOIw+Oc8m+wNpcpeQsnDi4tKaj+8/ssW3fRv5aRCld/KtXkMT4zvIzefYqwgQr
i7gmht0ycrff5XHD/impV8M8hUdsAE6wYUPZmleOSpLD9hT6lYCdvuPA9aOYlVuk
ulGooRC3A9aEUzjnvn7H4tlYYS2dMgkz8R+lOD+rsIZZ82V6vT7kzBkdLrQOqc2N
1eQierbP+4NjRWuk/YXcAEcC6c8ETPn5bcUzC2k926qEh+xvJFolc7cY9yIkYd3L
cczuen4ynaZ2GDfT/9L1YNXLGKaR00F1vZwvMyBnY2y/PDRNjOiuL1cpJT+tRpSa
ctZax5Z1T5INjLwJ8d714HdR8N0nXvB2j4RFEvC6TTU7pUcUNhdWZ7DjvaMNvYo1
UmaxyhWGgk4rMUt0ldOxZlZKX3KaHyO3Mi6mR4DDKek+qX0BHsL050aarjoKTCr0
PkwRZyVm22mytYjHjpV/13kmTNjhcR6LHUuJTN1oC/rsCoK7bEWLL1GgmJDDEP47
vjiBgZ6RYG0zySf3+r36TTyZtS38pVmMcJP0NlzocxLmJIBjzaHs/NB1J2yHEo1y
mBxxftxIyY48CM2qZkYaPyPJHlDRha9UBoHErbiuqCgO4LP9WbV8rIWiLIkllgSf
RjFiJWgHPBK2wzx61RV0OZ4HK7aAHgSt+TGgJB95xzVrGoim8ii2YUZMJardAKv9
LYXxNWbx+yvIDIxJ+U8HIGwm5D7+nTdI6//fv5WyLznU35wR5PIeT/9l8Hjtts7o
bJz78KdOFadDGI8Ayd/Csa7HcGepgG7XVVdYE4yuo7FpQIneaJiWTFCXUmlVDVUI
jpHu3Oo8sAkh9uljEF4NvA1T/UwXg3af0Gmmtgwn8hHLbVbbBbGN/wdLw3yKV36b
quharBJQyMXCOrUMsdW0Galke036X5dw9SHz1bHLw7G4+AYW9JT/V87929RQZL8V
q3utkMc/HBjylwWRVyITAfBPk1DXtmG563JWmrB0kyxtXuc/4bIUk4wTr5vlrJML
bhhx8AfZWLYvPZD53AjpUfQC4vWjUennw3rIzQjYItln32AyIZ+vRyGNLiRBOpC0
JeDpKnJI5WZqJ2DGgDHY0j6RAcn4FFVEaTA+AySINqXg4VQHeoAjnD5fojXNh9WW
sFrRdlbR955LXopOIRS4KZHw6Px0Neexb0bdx6I+R34rndJT76rpqRuv+c49dq9o
4UML9UjjQnypqZe4UynhY/ysiM8a6JZXKN8XBbB6Le03YYZFPsAcGOeLvp4gYY1d
bNzuu1anRIpBgpY6PetOAS6sR2/ND+dJTXva6Aut3EcymL19EQQLlQfy8vZ5dwuz
0xj1Ch2SOt3NRHpS8GDuDC/AX30iToCu37K0U9YQUcQmiXSXRSlimA3fDNcut0MX
O+PrYEg/YAf882s6cx59fREwKSAmQPDI03BiZOQgz6pivgtHQZg5BO3wz8x9EBrE
eJ8cfG6EyzWIEfjEmPUQl3o1sXDvLb4HgEgn582hHQy2gjDyj36LiuJFBmCMvW/A
kFkS7mRy1TCZMgtJp1pK6Y1cdUdacS/RW9SHk8si3BeRxNLVOJq0XeK/LzAQeg8L
A3D0r90NM2KRH+ms9ITJ8WVVeMtlvbIwSUo7RE+eOml5WNJDuql/NKSSm2aBKgb3
ydDPpPFqY2wg+n2TBe/6Qy1KFixbYEqXuSn4YyM+izwJ8VbvNoxlgmrLb4UvVjZ/
LkiE7KQHKHs2c1yJZHUAkbu+ne+iZd47zh5OiSgC72+qu9lNKl2VsxBqRnCUuSdC
HiDGc6AleLgUK77hXMkE5M42AnYy+Mb7pFUgNQ7a0SYWRao8Q5C2z5S1rq77VRlS
3gwQhIGfIO436mkUT9dTG1hlxpf7lYEJNue12fCCYN6r7+z9MH6wbD5nH8jUOXK8
qSk6l0S6EZjtv28mhDyvsm+kg+WWoI7DFSSXAkq0JwlnTD5JTQjGj17nUB3+7QtE
tjcCQXUn1RNpe77JC62A3ESWXya4xVr8fZJOIBia1YYvJD4B7TCNL3s5R5xDp1Ke
GnLNCcCkGgXt3GKkzuXMboHCxQGdoEHvcCmXuNoQW5C4Yxuc0NQL9LnbA0fnfEO0
scN/K1dNBWH0diFBFVMF5fsRjAX88AhIHo5u1rDUCCC/I8NROTB+68TIIGgPTRfB
Xx87D0PIMtqe3pyefj4cMcxib+Z0sZ+NX1cIyCJx8/gURIbRHO1SVeopaxx0sd4I
GG8fVsqT5BH6cSUJNfdwnUB4c2ZlvK5fO4OkF4axX3yIQ3LnjwtOeg7LbJl1UCGU
3sYyCgl2rGGKfrPOdec/PznN3AdusgkIBjBjH1ZGIwX6bPxxtSZSEb0rwzKzEUOA
XGaeK6qACCLLFjdA7bTah4q78U/oIAscZPC58/HgeRxbUtPWYnGHDwc9R0iSDbs3
8SWywYzeV18d2RkuufXc0BpKOYjNKBvt/vNKz/i3+JMb8aHZExn6oaV0f8QQdkEo
2nd0HhNODmXnz39ZZn2TbOg/sBGMSTSVbkkHmPQ0XBkhs02r67ksjZrjBgUO0Nnm
eJA+fNr+sAw/ST56blPAjX8KCHwp8WK/iZzEONPL9ISJQDPbchC213phNJ+1mfM0
frP72JwS7XUend4E/GlGL3Win4s3f0N9H7DFb4KlW0lSYutdxdEfr6yf2Ui9rgTB
taVVRKiaKk4y76yX5FDrfpEeNB80xrrTcG8jRNpXcd6izFt+NXunFrPzeZfNlY0X
l0psDvNOcomstoinUWA0fpWD0gpI67lqLNffGndF7/lXTsrCyfrhwNGY9bECst2R
gjSjoD64LM3idGbNZvIk3kVS/bvXFZBON9btCj8kk2BWQAaDq7GVhs9+k2LnmvGE
igK39KzerCAcmKOm++fMiO6EnQBFhNHXimK7ex4lB8/5tEaenCwDjvNKUG7s16xl
x1KlXhLAZsZtjrtif1UwMjSChwGT43QtGZyo6pFVz6lj5ko6bwp+iySzxLCi+HB2
uAwsUHSqJWYdat2mDnRh41wi/qgBTg8iLe6JraipbXsOMjLNdoUvXGkw3fCk8jec
vgx9QH5p3kuHjR09IGdmhfDztPANcg5cbgetFKU8rfmdGX4Il5M6ff0sRM8LBZlF
KGPOP+bdSqaLN2eGlXFkvsTjgy8hTcgCCpXkp3QaYDymlx6s7haNLpkRNiZjcevG
9n4Zwz3As7jKV+a8ECLTDdUFn3/5xxFBDaZAceXzlJCdHmyeE7/pwooE3xST4wvi
e5/nJfEEPJBuRZJgZs826z6WgaVtxEwNiDNfr3b1X72VQQvfsCVQnTYPx48KShCB
NdPlOyLvX5lA3dFE0dsL+OYee74z200YibarUzpw64XQR6F6XPkeiiCObA6VXFUK
P9yiODRrwHz+AuMjdFfbV8iWsoeRRUXSveCOPLeoD5uR1jAqy0imanEpvw8KKjbc
Ysq7CNWIzaann1mDF46/8JHtRILgiwDArOB3xbwIQL9L3dihHb7E2EpSxqQqWQjC
EFhlTEr8V+wfhUXYl+AE1jySrp98rqNP4+LtOETBRwbh0DWabPQ9hF9n1HGsFyte
i1WVmw/NRiWfIlQsIrvDlSNz1b8liuCtQ6PHWYk9GfDf+K2htonXKg8cDHhgHmhd
dJ8ylQirG2z7ciMWLl2auFogicjiQsNb24XG3nnCJt5mJ26jI6bk2LhqQvaQhOga
KcGAVhHDyoW0t3KiobQ+Io2m5yWhezq+599+Z83/QiJd919GRVOzm59TS7gSh46B
1a738mSgzCFlKLQIgfp0RFswsu1hmoolIVBaQO6q4dL7z8qHeHXqrWTayFkIkdNE
ykSceJpAvreGH1XazFUwfotbxvj9STMeQk+uP01fQ5GNzvCDjuvhHd8a0pTJFwYw
yHXL3wrBUytEXjgvy9CQyRD8Qlj7JRPcLYZCS/bOt7KF+2dvf5ADprlb3JZSgQxK
LUBjegoqIb1vxs/nV30JQ+8YCWQzL39QiieDyBsnfVJoIDg+cvB7r8EfO9aUD9JZ
m1adjMHG2U3b4LrEShhYYpyKoj6bwOO7m/nhIPIFNf8DIYX6aLMp96pRwSEqoHCv
yhxmXMo3p17d3Ainn3jWb8BL8oCem+r2Lo8z9DEgsOu1tFZbkGhlUDU5yAkfoxEK
j8yfIOvIHbl2Dn6IvhQhi9jUWnDGd+wUDBhHj5+Xi3Ag0zSJ1NLZ0zs+TpK+4g/8
TtIELSQ5tSzz/2FJiQ5ft0rZM8B6Ryzi44yvYFeN5KgjrI8lMGiCT+bOZ+2oJWPr
JjCJwRXRKQUlYMcZ6+8kZVAbjECCZ/g5ZZvrk1grdkVXFDV78GHGsVr/s8lA9kVH
5Kl3I9gM3sI8pHC4NpdWXj8zZFVdpiyfVLmruSIivV79pGIKm3Mvxg83h/IA83Kg
8119p1RWaYzfZNdUNuissRe9i8eF9MgJSGoAWkmFl7Or4688KjKiFonqPi6x9C8w
eNqu2S/1Lpri86gTNKD15LC+nd0KZVtSjtRjR6ZCv1OdJyUOYcLXEy1USf4vAY/+
Dddm7S/x86la7LJ9bQ1B28HC4iasIxSvpo5djQX/SnktGcK0X4MLGwHrZ35H06XD
GzE8N67MGTvVU+87e4rrdXeWkmHKtHfSCto4IOvCbPa5I27ptEqwJOHYpF1oq2Sy
cZR+XNIHnTQ06i5j5u/Yg6NJTQGOVvqlSBHiWvsOufaD6j8dSqp8BWUL/BdGL0HP
mH9bNPdeg8XqcUWXzC54fDenjrVqToPCqB8F22ayZKeTqO7yJHcojqO1KxrIQs/n
6SWNyZaGIOge1MfwNMJ5G3wZmbC8+O5FyInZHbdir+skBCy1MXEHhKVZdQVGYtCf
exea0NVGEI6jjMsksTU0luuGSePLKVx9oTB7SKqRm8hSb26gu2y+tOB/Fd7b5ZaR
/Oz5AtFVJDPBtLGvGzQA7/uL0Ks7SCvCULD2s5AxxjJZg8jAaptXSvE2DWy+d+QI
d3ic8lyl/EqJxFFuW2C4ZMcjsp3DK71TbMjO7wHus6u08EBKcrtpX5iuL4I/FWWt
oEscsyD7+P84Hx8+Qtej5dpE8moSi4cxOP1BVNwWu7cJNYDI2zPF7AgoANJIj2Z/
0k6hldoPeSy6SsYNGyWvLD5CKQaOnDwUXeRy+o7xLcKRoeDu27flzV6PdiwmH9V4
leB36Kk3T1qEDYz04Xp7Z1grdk8im4zQwd0PRS2IzvDXiyQXN4TXmpIvLQkgyp0c
0F6/fCUObPxfpwG+xAcLNr2+Uz/a9vs0BEFUTT3Rw9CPoE+BHDuW7jz5LprG3K/V
7R41zJDfgB3QJxT6Mx7f5tbwnRHMnxH+qm6EymgU1a68RvVs6ujIoxBSASoex4Rb
tSH3Ybd6g5Rs/Y7kUWsmZJ6hwia8wW9BXalR756IZne2qee86ljNZVSsgbYppbtr
XotXifgvz3p6EuiGx9YWCTM/ASARzJAT3KhZ1QfUDbK0jpvndxQaJKROfVxv7uAG
+z1eyOJZM0PLK3WyZna4yBsYFMWfaCyVSduMbwYMMToPhLvdHvtE5WUXWlJA4PKW
i1/DdwAEusJKjcXXsxBt0VW1ZXWHVBdq0ohzKN9JKtee7rwYvTwl5o5Tz207BtSn
UDyD7erm+6qkfGy3FUwZqoLjsAal48/k54zlL6LYIbVbqb9S2CtrlGWU4ncVzO66
0G01SaDqIoIpFDSJmqMLmsa078Z4G+UXag1WBOXdKXQAHA7GOkTFyAXvXyYlopa1
5iHwrbteVmU+bszfqc2rdExg9tcb8RWes3IJeE0nJbYvmdvQuy4GzncRdtZak8Xu
gRhrM5/jrrRIl/fRRrrFX01ceDZuCHjY29nqzhBGrCZc7Cse+E5xOjTlNoaNfVaT
wK1zncIZnx7ZWxDpcRRLq2FJ7Bq9uTgUe6cshW7+AOiPnzKDCG/35bBao6CcDXHK
OPhu6hK57nXS8bmecSIzyZHCP6TVRYYieXdESljh69JyW0QlFHzxSJHEYHJxgjbU
aI5LoZo+/p8WR2BiYb1/HG96LuLH5tLUotGFEfgiIPSqwskvn7Ooii5cesl25Vms
BBynpfXW8XhEctjZguPEt//lMEoCDEE0BmIkE3HGziNgYJkgO2ciNTiyJjJPXNTG
DlIePEYNQPJuaRZ0Sa3MJOndjGI63Zw2emYAX/o6oDFVfZpAp0WX8qa/bI6zyj4V
VEOA3qj8a7Wwaga0d/fAeKJnKl1nknVFJyNd3MC2jdiEm/GaQ1ALGWyWeISaSsPg
olFL41KgskjveFo0gkLnVn9tTB7mucj6e3pDrbTShhiBrHqXN8VYROjcr+kzhezS
wEEKBd8tjXXnLts7R3bnIfgP8XmjEYUmJuhYHw8fNy6mEo/xYBA56rH6y798RiNL
+lO6BKsIBy7dH950QINS9VGqPk3mEZNvQ/MxFvFivMuiYv766/4wQmEhHqBSsYuQ
P7ruKWIxzS/xxYVAUyj7A1ovAnaw2+YPsnFBCIQWwCeshz90zFs6wlBFfH/D79it
9leYAXAyUSVN4kni/4wnYtyBeqjovV0477mO9FzYl+kFPisEzVRpZN/68E1subs2
bO4hheNVvTo+0Xzo0sZBjSGramxEF0FHy5zK6m0XbdkoqZAIVFtlbOmGg2MQUqrk
9szgpOFguaZFXlzqsjg6CBXcP/0Ll04s+sfIApPv2tgWXvOfjegnnIY3hpkJb3Vb
DSGXmn3LgnJrkr+KAMVr/Iy/KKcQc2nGMx40QqF8a1SyqqkJ+7Lddgj5mm9RQFx6
+dyUspyYNRfC2Ybt66kFu0pGBaCRY1RccYtFRapVfvwj2Mdm9ztsOIH+LQSffnap
tCRSpcnjmOAG31XNXYmivVblxGkDsOZ5yHM6HRWUzQo7u3ApvpHUYpO354o+w0hj
n6z3s78iHqfG5bvfWPr+YmzkUCB4A39f8cPG1Wryj5RSVlnHBJkzNSdqT2+JyPiO
ZTaBQd/B6LbtwltwatvLJzv4D7lTStudwzZWiJgAasxmK6gBqCfcdYxz9/r1UsIA
EbicH0dZjp86mxoSlVQbQo42RLysTSAx/yMrGQ9aObxEnEmNfViZg39GjX0sTSHX
eJjmlTRL3tLNt+fvRzVofiPk4y38+TKF5sd5DcBxWDiAMM80xOOp8OXxkHcJ4/Wy
nKBGTErRRKbQJYTveGKuUp3aX6bDAlFPvKsA/DNWLu0gc8lQ45FDBv/Hi2CF30P+
tHpvIb/bU4IYtf3xUu/E+o8hyRtb8YXAmtjCzWebO6Uk/M4Yud+NHgBhK5NmoJrv
owPqNwbOhO3uWkcANIu+A0zjJWjMdpdmdIcRrIKdR3QS+mkxwmqB8h9GZafWZA8Y
1FlMhlOzFXtgfdySVmoMEmCNzFUhH7pK+EllqPJZTUqhL9hR9mdMp8S0lBUcUwks
sxD3zR0D85y8wfqBsjSnyU6xTNpc3wQyiILXMr+0nyP+wjEO/G5A89to/5B7KoSj
T7wv4OToXzoZXpKuruO2pwbi7j7jCv6OyQmWfRdbLi6n1EHGrZ/ojWYylwxEsgBJ
IQDwud+OZgr56dZNf4PUGG/uOfhMBRvqlK1931pMVwrXVHx57f/5L+fGZVqSvpjh
8Gh1hq5gGS+VsgQc7upwKCRcWJt+uEzemlQTZ+w1Gn3D+OKbw7l7crqq5s9lg0m0
9Iswa9gWgtPPSwGdm3vhRZpsMb34jtucFdwZYDiOM2Haq3nIAnSO4uztGJKDTvIe
8MQdkTfcjgaSuT+stFcHOgEgJ/NymzBgVU/7LJIdGofhLJAkIGjcc5yMSUkxaK35
BLL53nK/QHOW5Uhl/p2hiQ41A82rbuMn8wA3/NjrsgfKEKhJdoRIiSynwLV5tbYF
q46UFHvlzqd4Vq8NtFx8IPgEMU86l2TmCnHiuiAhHE2avETjMaaE80pw3Z7yGfBo
4PSpUQnBQ4rcQaVTGCPoeKQsIFLsiy4DMA66pGpHWii4++J3Xo/pqWF+B94wd2df
qYTtuTA8J53fNUA4RtnuraETcaZB/Sdta78jAkGe/V8BQeAC92TPWvuKOx1MpZJ2
alaSW3lmlOS+VUWDCz0Vng1XDQhSOLLZmnXXk/EUMarvaWMexxhBQwG7B3l2WCtU
5ONhnQIrhQpMpk7dHnQz+G7Ytxekc+PF4dNFXgpY0nfRe+AE1B2qBcse0Acwbs8g
iYoi2cD6VvvVDydg0a3lV+7UpEBeAd3ZMfejoWK2KjiWkUlj8qIsQTFp9mZ/df48
rboYnox8aqAV0IfY9Ph8T0YFpOKH6oxCIc75ZCVwW670enZRA+STUYxQafd9nLFU
Kt/OHce9fze++cOpHmCemTbio9flbacxPYQ90XLIIFPx7dZKTbF/Bdw1YTnEWBg6
ECxxtplF3ZrWJzwyE+HZtS7TN1IVWav55HlGNRCwlXfPYbd0MleGGA9B9bcI5Ne1
4Moc91GVNmp3OoFGYW46xZuPPMpKCcjSo40zst4RASGgD4KMCW/KlEDduExj08sq
MSaabcE+PqLlhFTg9CbtOy9XmCazwJLRMjWSdvPDnGio0ujo/DJMnIwTZdlfEz+n
/W7OtJkO9lXxvfpLgNKj/ndOjyB4wGZbmY01R4aryAt1oa6DJmXwXDeQSKLIPWPR
7DSFs4rB5OaznfFKwPLQMxhMAZeIc5owqy6HZqUUgirShg/YiYnaxbclHsBOZCFw
vzTZJZH6W1R6WyaQgYFju5fBEwcYNz+0jGVX0vPLJOIwAnpuC4zDU+YO2SGQZ82o
lMcoqwwlJR8l6Rj1Rqaa75iZc8uqo1+9gZaAOavZ3l9QojrFado2h5ZlDoWoe924
TucAn5aPGgQ2Z9qNLuegZ2xIJDwsNF2GtxL8+z18ARgLZWa/91aJ0OrwWTnK2qyB
35cKJipQ8m9Hfbr27IObRlvlXdhvcBhGuvTE++Xg+Fep0MkvE+HG0NIfQWDHAMc3
EVq9Y9uX2MNYFGks/NKSMDnoy2/pvNm7b17Law2pjLmK1k+UECZ60gCNvJaBIZs6
fAzFvTsjT6PsS7eJoPW8rE8FRT3FO/Sz47ySk5yWrKbYMNintpL88wizkBfgGTvb
tXcy7F4UX3PErMBXEdfsBcYLJ1AwhU1jgqJLPnNgqBKqfi/2QLb1vWINuCCsn84r
TMdA79dTKj/1qESihdhle72F++kBjiH5i5i2S0aPxiBDeOs6q8DrRFpXJAXIxEhL
7wjUWW411NhGR42lzwTGG6CFp6Mo+Q1s7aDLhvP+bQHSRSZmA3cwKI2PbzT8Qu6V
/PKSivIMKpeuryJ88kC/2JP1Cc8LWIxts3GGLOdUk2/cczUjNT0pn3UkDcnAQ4ij
1IrjHdew+mdvp+uLA1HOqJr15M0DuXa9DUkRaQW+qdgoHalyUsxDOr6MgVqj8+fw
Sl/qh3Ehzqu/JIG9QACqBwhk7r34dlHVdMXOZn7yAYKP/G45ObfOoy7OvVsnWOFm
nvoL3TP1HagFrAwPGIfzGRw9pv4hk6ajcQv/Lo4fGRJ7h0vi4fL6jHwnStWJ+7gm
mUKtJLcdL3kWpIPk9Yu84ux7acFdjAn/EQlAppxkilRKwVRDNOaxMtGtfLIhgM1T
5BLgOpdzbsxpE6NhpSKX8tbSn+vrTnHlaaLG7MMIMoemmR081e+i4M6aGnmqlB4w
DMtp+W6s4+EVWa3JKA2jxQRX1JIfaq3ZFz+mKUB09m3ywpuFlveRWi5eQq8elP2I
djobadv5SrOfFP4FWXKh57xSsgtvdI8XtjwJEeL3ZxrY8bKDT3dnzeDALXprzuyt
Geg7tEOsovXLPLvs72JEfTnFtb+UetdpS85PTCjvxdzqCVfp42M2XqJNnZ7RJaIl
GBFPu9vLmedwuZBcSDm6Z/JGXsBD64Y1f2QePXz2GsI8IH2zgSKso9uYRk8D7bUP
wYfO/LNW+LH1500CGBuIkMtc8nIOVtFSs2iK7jGu329eeTT4guxKpY6/F0CM0iVg
Y9e9B3Ca2eyLiFpasrupKG+YB/WiQkRJ4AAyYTzrGUkJm0XvMQw1F7i8RWAWRvyq
bdBMlSGZzyjRHgZoLAi2V6Z9UQMKCbxEQd2TijvNgSF0w+8SDVM6HT//ZVUioHa/
WYAL09hqJNgmsenRi+KkqRFKW9eK6QqOfu7pxTfm1C+c75zMN8zkD29nt5mXpbc2
g+SLwQo+4u67ByGeikPTEcUv8fnBK8bax0yOeuJaZUXsBBCe8bYtm/suLhFn6UCg
E0UpQ0iUt+59b1stRsX+CctjR0BFmUrabAGuWNiwyUEf/7tJqpXOs4DIgQA6zOcb
LHJmtLEosqdh9WNrLbO+WYDmBR9um2bMy/i6BBgxoTwtmCcsOoc7zVdQ6gvyT8aP
+3aFZvdOq0zWYpQcaUVzKCZoWHLQI+bGZ2lQZJm+C2UfXKCFFdkemHLamHfkY3zT
1WlJRx9s+kD2Y31u8p6QgY5S+AO0D8yiejDx66hucNhbB/vncg/7ASFyfvC5X75W
v6a6+QmWmvEhTxN27FZfoyJfmheVIRc1AslGEvn3RIq24Nr08m9C4gHd4bCs+beS
oTFfezxTpn3MeAZGe50M2MbpEH2lQNabnWs5Qyl3T2K9nWBA4dqwzSqYqFUO1I9s
JIzA8N+svGoaGfHClgosi1ySNn9tHVcq16HpJziUUGvC/TmzkrtbYZkxKqUlJz0V
tPKUfgZPu8HyQaPfI3bhM9ytAE3NQ5/rpXJbLT8B5+t0ML1IqdU+rQr5vXCi9Z3y
v9pENif9Ue6e0CA0taVqV5TCxX/yVckFbn2snMNraA+ivGIEnhYt+VbC8YX0LrRX
K+oU9Of7a6Ay1ML7T6zvLlZT9Al8m3NXSo24PiLRL4Ve7+STrnlFrv9ndRb39cje
TGyJp7EYrOfYwpqA3R8JCRj1iOlsPuna1wnyxnWI1EdQfEQVyZIsZ4gOv4yBDIs7
dkpHgldHjnOOSI/Ex1cd0kpaEZPkH8piXZOaHf0U2zWk5Tam3sgB34y1hsD3fMBh
CK6Jgz7JHirD3LJJWIKZRAqRmzow3UuDomfqBgRo6mPEkmbmbxggBgwa2MY0sbVf
uyRu9bU4DfAQ+5Ks6rGOEs+W3cmh3jifNoPkmk3txXZ7fEkGyGVGj2IlJeP3svhQ
q1i1Xo601Or0+cxBa1+EaoifDMeAERdEgypf10GiEDvizUPvW3QjBpCLEP+Xbxya
NN6t8CxetVyWQ7oQaCRoTLu4gGekx3XoDLexKuZROxAiRLYJQehw+6rYFhcHPak/
vMP7+oUnafVk97rZ/s7ZJbZBykL8IoMxbJSj9pjuWiT+6wlblHQ5OEWZakKF7ISR
5pOHax+Du/JWyWSHP1pMuaXsDP14bz6hc1sNn8w6GfQh2XUXCNC6pdlKho+GmQTr
twK9H79JAWEKSscf1h1soC1rf+Q2ud+V0E/kvmTth4HWacVEjNMHaLfA76mGo3gI
jH9cu4qhgIANUX9nxLbwjpEQa+pdhCnUcdj4fKu4eddrnh6m9LI+EM3eKi4A81qC
syXMdA2iSdMW0qq49apnc5wbg7+MUo9qIIMcJBADizl43MlIXWZzbxiY0KrjTgXO
MRS0NsoeP/Ut7XnEwKVjwQ2UnyB4h8oUp1nxoOXrJTQvYDqvKf8OuT4Hre4CqQ39
kSWTZ/+Y9l0H3dx81PdtV+vR8vErp4SKAUBlK4PfTr8rk0NtsQCuAni6+ASBjm48
Uk5drna66xP98nlpyKF2EiYvOKDSushbFMogT3uwLHe609yOSPb2HUn9xN1esXc0
TeN/cziMCwUdm4RM7lZ8EzfcCtC3w809dDwOR5/VNIDMcke/9qRsS2knkOgUEtyj
eBLareJ1cAHgWGScMyEvuSpeCWi9Yd7scVR6Is1SzMI8QNmqiXwd6/h0SO6liVvF
nD8qYjyeK02cpaqUPsmsWB+mwUZXwM+ksAphco+hff4SaXO+OZ6Ae2+tNM6lV02x
i2dWsMgu+ILmKqb+EL6YqHIDiWkl2p5FabBulU1ODORt86ENkdpw1gF3BcdLSh8G
Do4fbpRYnNUdSIQCrvhumVffK9yLWxVJuTsDObGt8pxGNRyDsVr/r0VeDtCFCOLr
c8Dvs179OlW6f1e3K6kRMTsTyS0hGLY/yKzCX5Atxr+AGSTJzjebZ33d0S63BZE5
yPNF+50gubyxWtpxBd7hrjhU472pJOJAUA/xcjS2ixiHjn8XOUdMfZBng/MRKvY6
i7Bnr8Y479mFIYSRKVQGAXxlXtJe1yKus+AOa1aGaNRXl+iNHABenkhctzgDKz/w
HsE5zPmgYeKF0b5yyEpwE27mpNpZWbY9IwZVMQnLgEbdREwGVM8DfpQqUgXVT47+
vohJPZmCpH/rR/LKAtEK0bhUrkGfc/b/XGj+DLgbICow+ZQ/KfU/Q1TZeeH5oDV8
KmJ7UXHTVT9tMbkHiA/tg9+dMiaUvHi4uQzMPKzfEajJXssXboqPf4K89CZbdi4l
hhPgYlogz/CBjWY1mNZcGq+ccYFFBDGdlYjwbSt7wW2THY6hMYjQ0O3PHEOYRBY/
6YCdCMEbCJGLAsCHnB02vL/cmMRZfDeywutjabVyxrMs5ujF62nJW8Xdr5DnFfH5
qW0r34JMAWdOIL6KpOjKuOkLAS0JLB4ISMyYoheBPj3cDk2HfKEVVN4vtsbldrNU
qgpm+npGtIYig13ozQ0cVzW1r0WGiKKjif/qH56a+tC9KAmqkXXb92v+Ikb3ouVp
HCr4Zma20TBxNUGxknW3yc18tBb9SqtxcDFc8J+JrhFdk8rD/HZa6yIAFT9KVGck
Zuk/HHx0vwSi96qOGOaT3aTYPQor+GqgXLJ6EBVnGKzNwvmn4AkPgrFsERXAHLfH
X9ZSaR3PEvvZg7h8tYOckZfeg2KVK568TOtcTuqQ5oY4SYTOE0p0IjpymLRrczeN
Q9UJeCW5ADmoNyOdtzoH9Q5sP4PEFh+AbBI2ccjkfkG/H99G74STmy56xHmQ24GV
0PI7sWPt/qeGjqIjH9ZUYvUAiXcDEJ5fV6KDDUUTl5kaHSSt0DFcwqqMH4ycDQoi
h6MlTwNXYdKcs56USFuURlL+r/gi++SulqTbM7fY1NDQ4U6JSXuppEsbYmJ0it0Y
QqSZLuku+cyCv9NxJ4xRGqWJ1mQw/yfT8NtCA0IzKpOvRiJlA9f/fsQjXl9QLMmo
wKFLhP8ny05MYqI9Pi3krHhLEIpdGt5/PTykBATZPEeQX21F6HGgoXFUl38hY70k
Tyhm1dMEoIbmf8ibDPi5A8Si34kclVmzgdAO+1xAPvQTESLmJu2BoNACwfupwcp+
nmQif9Yu8fyYnnEmVW6su2R66OCPepOyHeyfDBgBmwYTTMgtOKp2wCpP3KA15KLS
aVhkZXK2R0rnLmW8/dnsNZlQi+Xy79KEeHsKj/88yOcoo3VjYJPel0pL1ZK55pGo
uSHMHC0xwBm85rKMtUtM1hfWY6wdGSpSf0rLIiBDp1wYivdpNmRhjndiCkAqWdIl
em9ShR9/8Pz04zhCWM7AoomL6OZtqXOw/vAgr4ZYBuMxbE2ieVkeSZftaCZjptMH
FOYU3OpvWgp4e1prAXMw/+oL6Hz2ETdrBQ/Tn0+EG1NLxldyPQ8xvaY5UpyujNYh
gL1K32vR7L/ZvypGVILKzrKDVbOLmW5lknYqiW9lYcgHJNS/lX6jjRGSHAoZfWjB
8XH82CIgCHj0rb25yaI51iJ54+X0D/f7ovPrDlPDJO8ao9DmSC/Lw0WsPmeviWVi
BWkx3UeV/udUYI6D8+TWDJ9e6e97V+y4rPMmy/q+vim+A93MqfjsbUzHNRRD9HCj
RIDnvyj6WhlqfJIsRG4XizixB2pDr4Xe7HTv1DnpiNk53ohieZSQ5eCIVq2TqJd9
IoKjbZG5vE1+AUmmVD5dZq4iEv60lBvRsvQdQHKk9NxokkACvcxnevLhPKO5TxNP
6QvGEK051zDN8dVJ5CFf+TEcujQzJw1MlSKfZRenlfNSnSySH6Slr0bq/uqnEPnK
FxAaJLUwoAGmRcqRI3qKZqhabrFuffRxtQ4QThWViwiBchffTFYzhv7+awPweNn9
QUSBbikGLPvkUzn7DqEzHLIvWc5t1rkBsXi489fyHhKreGks1WmvUs+UnxWRULNd
w+bgD/4K4RankrzTE7aaNMPI3ttDNtU+dy9AOC0jS/qNorgNGyq2Dx8oW0tMs6tg
DA8ilRt4Cuk0J9mNGHet3V3pjZAv9zINKgaATg4vSEVfBc8pdDzv3czBPilJJUvA
+7gkQa3VlWj9cZrC8szzSlFZ7p8ahtC9lzLMyHljS/UkSAOVUz0LrWYJGXIRC1Gx
sMbw6lSPMTWVf8/PK8H99yM7Mta3hltw/kKKJu09UYCbS3K1SqIQj77Q/R+pG9dA
3ubzBn337CV8x/xHRbASJnNeNW157Su9/DjyibjI2LNt7FfMMH9Nad49uh9wNXJZ
geh0dTib7ZMkvvozq8l9X3ug2DprIp+xClA93DmZpUZ3MixjZz949pBL/ApiDJ2A
zSVXsgGWBw55DbI1TQfhj6BBF4pV/bBmK0iDnIb2lfs1oR6lo+mPOfO1H8YOatyx
KgK9OaU7cAbvYcSTz5DJo3Behq/QZy1Jz+GPMfkIVTi4wchbbuuSF+1QvHUckM4V
Ds10bzNxFc+ipmgY4FAJITES/VC7ZqaNbB2m8pb/bR9i2x0iajlepgOmp/aKh6LR
a5CBQtQIPmayriwvmGzoWhSVeb23H3gFIazZGzlCfNAs0Dwx/qP6v8Bas6ymbhG3
A6cEFw2JaoJMNBnb9m3yWFYmqEKDGLr8o60UVWEPg8WiJ/BGF+kKbDV/K1dnYWBQ
rYBdGKaWqVdmLzU88IuQXh1czC0IsDBPAVs/sz4FVFcI3aea0YQ82I8Yu+vngpeF
GVeVR32w0StnbncnrVuoCPNtw8yBN96s7oQ7Vwu8hAqDyHvNnzC7ltAiK1V8EDgE
cotl2FgS3dpWN/8uA/g54NmoyLowsqjGDfns+MzY9KCFVDlC/9uKqMvE0Z5v75f2
EZkczSZVyf0ZZPzuqYac875mLqOLbLSTsHgqWVdPf13RcpEvN++aGqHWc3WnY3YQ
KImbpJ+OAR1BYFIXYGYYn6t7+KAqif9MJRQ+tYMu9CcFHcFpoEdrTh9Ia6qtfuuh
C+uvz1zz/uLFT2jkDaffK8twgZrhtgAHsWTd5UdL6Vx/b+/6UAfp0FMQbmI3gRhk
mGwVNmOnPNk7HX+6NFFSlPl/ra4Egn/h4EHmZk3Jh+BEsj+0NF8ox1IUNLMnEsTj
wNNDLRBodQ/MkYeNcEQnG8UMSRV84KwARG1TqFU79dq886wEKaW4kkedJI154pEd
ymUVTt4Vpulh5d3CFBCqxec7RZ6QCyqP7pLTREXkP1IAUvjP+N9DFPmTTQmrU8xb
Tmy7cgXaJZcLhoSZzveuu2z+9XqMPspXEh55T8nGBX0C7P9p2HUlpscURyI20t8h
GOyRx1vchWGOreLxA/H6BzHQCQw/7H3Rr2xD1tO7PT8D8/mECzu9TTkIX0NoZREj
UOTwt02o54WMW7FWgMw/iycY8O1+iHx7Gqjztk11veHX/1IKmn2yS6nas/eX9nE2
+5yXu0e6EuCvhutuHc07sSOQ3An2p0DYJfUDZGFEDtS9R7YUCLBzicuaFGh7FUa6
XOn9oBWEIn9Sd3T2H8HtmDthV+vVEKol2fhVcmmWP81lwC6/HSwTAR6x2ygk+y87
hZPxRtDA8yCgi4sCzKxIJbxTAI3km1pvRqrMJY/TlgLb8DAVT0rlgBGPhkgpUdQt
Y8FQW7HuukK8CsnqQCRZ/nb2OzdQpSHBQaL5fomRN/lj7PnSRfNx8dQ+RJoUYqlz
KkdObOBtjY/6vxdk7FUwIaMWh801BC8JYsjvB9Nl5RBT9+ARz9F5jot8SyFSfqi9
gRt8luMfgoQaLax2yTZ05BLnCuEMgbcjckCdZBmdtu45mttbuIEG1djWoOHjAdtc
OeyvOnGRFA8bh6h2Kk1U8UWKIQAirvB+t/2hW3IDTBPlXEa/4PJsfMT+Kb8Grr6z
Xbr2GDh/wnZ2e1yRlBV7a7U5L6FnGHF+wcKTBH98iXjUPDkx6B6vT1NOGgutyIVZ
P+vD7Twf1Q7UdBCz/W4hk6wTfbCGJTqGx6VYKgfesB5x6x1zp3Ef4fMbREwU9aaZ
V3vM8bZJYU6JUUrmC6WBhM9I6YqMrFf20UFRw3a9iE/TL/If81wIfrYIYd7GvXpj
G/u+/cLtWy7BVzFa+pV2N5aMxIXPUUyg84fZwh696rbfRCic76ljdVgsrhtBQCy/
/K264EfeQGGpK0sCfFU7v9js8JkSs9r28zhut0q9xEjp9WgcqOtUi5J8p6NE4h4l
S+FY6Kw5ZZnAuwHByzTYLqekhSncwK6yNeNXWMvGKVI7ddPqgQW0RhN1oGHUXrbk
kptD8aLtyuAnCPfRARrQwqY/VUvHCEuxVbtZdfj5x7BJh9NEZ1Aws2KtGPj8wTYp
Z1UHWoC2fffyhoGUyqBuEIs54wM3DgY2XQiuVRDMbYxvueezYlRHoReyQ4p44Sad
fjbaVnxsyUD7Vt71fzhaAQ3ka4pWo9MxVne1zgaMcH7cx6tjSpOK9seFXB8y8Wln
ZwTYjtduiW5skOdDh6ohInC+3uF+m9csi0izSng+LvfgZlb1ag7+1W5SNY/wagiX
fkkeUj048Olf7J+hr5etZOjp+Zg+FSWCnNlIXFXMdUUfOWAEopTWqMVL+bc/riTf
hralEnPrjZm/YejCPAy4UEzn6o3zimKjzHgLtT5VURTuD3CUFHrfMOnVJqtftG9/
xs/jXZ0q9GLmtQtCG57Rhbl022hbe2/NKUO7H0xuMRCi6aa4/z7XZgcQyCvGBYlX
iDojR5GO008Du57LtkJilNsvxIGJLjraGXFpk+OGWJSfZal4DrQ3oYa4OD7I2hVB
NoE06JRpmrWg0jrKCK2NYwIKVq0apdj5ETzGqnByTHQ8CNCmyBYvcyg5zbFglQrh
OkZJe6fHLNecubl/uJ0y/W4UvGREz0JLGj/IMHAqPvTg+yQGaaZA84uwiHT4ul5W
exx0oDAE0SSA2HRq3tvPiO6KNuSVIaFd+VDEpS7oiO8IxycIC8uzeWdyCwTWWlVC
Udj484DZrJ4r9EnpbUg0hwqTbiBu64Ud0TD5tp7/Wt/2MThITY1mU2jgGJrfb11c
rCJyKb9FDYDtS8G6Lf3CaJdEVx9HfErrIWfHzVAHZqkAH/7H36T+V385Ro5fQcY0
nyWd9/sQCAFGaHJg4/AcCMyL+lT8RxNGVVscrtz9Dpcwq1gBlF2+B8vpmAT07TDq
jOXiHI6hKUHaPhPgVOkm8HVQlpjsaoeb4SGHkKSU05ad7rYMEvaHLDEjH7nz81I/
tJXUXI5UAcveiT9RvgCXhbERrCtGcKi0BsyEtTZ+nnKKw/4cIHoVqmdu73ymLoX5
irS7y1pBb5HZcxm13eRQwcL5ZW+sb9xvgKY+EbP5I6KLZsRZk4u3SkhkQg8NfSS9
wy1LJfQpQ5MFcl86M3fBkUjc+ko0pCJxEUCtgSPdQK3VqUs1JWuzddlGFHV9ynjv
WYS3WC2qqcNU3TKg/j0UH7TtPLumlj1qPYUNChKWfHqvEiD7kesIWQHmJnc5kF4d
4N8121XPefZEcr6PkIbozTUy5hwLvoHLPi5TaABBo1UG1/9YpI3sdTu8Jw6SJP8c
+40JCVrkpP3uc/sno1hAgCUbeSv9jr6PGRec0RsmxTVmQPi5A76DdruPSG+lqYHZ
yo1YwKfGud/ZTII6Gi4rb+2xvZsJURUYS/SnX9KVwEl5BmBcJ/xKumEw/9BmTapM
+wC+FC4U/TaRoz0xR96a1fEtSYHvZ5r6oMKdl3/t4+A2JQir8xNKYkqXBF9X4K4V
yR0quZ9uqGtqH5WvEoLqoPWRqdLf641WLJewp7549i+m2yNkf1H5UGp55JGrlzvI
55AuYZw14fGA5RKN1hk+FvwS3JYt8UZ5gBx6cJlG5rhjEGHgcGGj+WEowIFslIVl
pPj5FtLHFqJ5C5/y/QQGfdoQgONV/PyD+pqI0hz2kgRj94fUoPqAaSAjNQJ6SKjr
EfW5D4dUaSUKTW3JOcMU/rML4cBFyVmO3ajwb5tUc+lGLuS0uDOliGCltwzuo1p2
6gFEvmPr9T6xJWyY8j4T9MWwiQTEP0nRAn0m6iUn7jwhALFtJ57dpLcn1woJ+W+V
eSQgwXl4Gc14IBW90j81te+OCWSpkmtGkc2JD881v+X1YlyFIFhCcSHee2NBtZ+Q
1dEGVqxZ8VQ7JnM3GJekGvJqWj1qXKPbMfcE33Tes5Y12MPHpq+pDjMF3dOI5r4+
B59N4xPwkJGxKlnDoKz6KXfH8duj3/oMdiCWUHvjtPKYWLgLKzifkYqFnODphhBR
MjNYUvVjX+asRREcAesa1ACir8u1QyoJoOdthGvyQhgH+QL/8uTwNi9xJrNIKHjJ
LxAlqeb74MlaeSiD8iv3Rr54Eavpu0ew2eQInedEfVyb3DPbZdsQVm5oNALqr9F/
tJBXLliboxYM1IADhmvKIH7EbSaSGBIDyjZCie1lHBJ8DlO8kAPWZ4+kd8q5lWqU
UC11drXobEzdFnLAHLMF0KeN5IDixdwzPFDNt1bQIn3S2TDoD16KPQMHYsenXDs+
zTVtoqyAKYjLNUZdYJODa/BDR7KkxvnqJgB9z0LqPp9o/xbG45zt2dNgKL/38MOQ
f2Oc2gXgm3LniDrXpILiu4T5bxnSVS/XWzCWAOZTtmocU9DNahgiZDQVEYk9rD+J
f6BRiDCUop2DtHbdgUTZipavfGXy8hiaGud5uASTa9jCDv+i0IssFbvROY6rN1Tz
lCSZBGRe4gRwDq5+DF95iJGXDV9x57kzuKm5U3S3Mf8QLOTtxkj5UP1E6b3VBYHs
YP5j6pMmyUhplnADcSIyO5oAU45/izXcpGPfy/iMv5EOpUqDuAMql9CZvimVBzZu
PM2cAyZ+2NtzSU1Utw2S4wMZRiNLiPIKO3L6TnOqHIe6rHspUYdF6XYEvdCqE285
v4DRMRxfpSXnG7PWkzIK7PYRAuOomzG/4Tc0wUwF0IcawtK/pd+64jnU99YMwep6
n47qU//8GS0+Rn/+clJbCG3+OlMgU5rZyn4sV+0K55wT6fO0zKSk2+zsSfEDp2+e
d29ZJL9S6QrQ8JT28oy0YPqKDWTPNNo7vp2BYElPi4siq2NmukUxgSS1VyJtrOyF
M1GOBPT/BqEk7syNmikclTnsLPpgMieNQoT2HD2qOAjOQ59XCTkGKU6fLStZHyG/
Oxg4qZAASyKrzoEB9ig9YSk6by8iMQRyFmWANjuM0tB6kM17VDee1QCXPxmGuctG
JIJsEMNtl7RWWvYQkiOyBrc951Ja+BAY2xsLEwbwTk/r3WeIGvg6bV8Hhf/ILk6a
5tsCy6m/y7IvYUMm2Gf13vSvWPnpArfIzhg/fSyrTaAw+AH+y70549loox1k2dtx
PGxVMayeYC0nMZVYFet6pCVZeBajzaMATlTM5yinEgFHjNHOktL8ah4aRihg0ISe
fWs+PrqwO00rsVL0iIkZtyDEHKXJRwO7WsKS+bLrvRyr1o45mDyPAKvcNwi9cuAZ
5P2a3Lcv52SWEnBfgj5UgPGlSE5TUTM8JDieiDEcL9rnfrBwPwaHaUarplyJQftz
Gp5yG2Tz+0rUOG69e2IRvecq8Qz19nzCepPBouSvTrawalT85cYuBZonNvcLazig
KMxfhX2GWdyyRv/A1BFpPNV/sJfXvzaheFcqIa4f2KzNoXXtMP0TZ2bjFj5BiNuw
+YOnrxLw6itS1Tx9P4X1QUNyjEFacXI0hhLxoD/GatGlUt8C9GxLeubjwcZQsnAU
SwjoTvSUhaoC84A/78+YRCd+SQNkW0E+dMFk3rFJ1UpL6L0KQds7C9do4sIZ9kqP
MYPXigo5CyfagTHm2U5nywfSwJ+YzANDmbDNjscfFc0FmSeQ6S1UWNNTeHfzHt6f
v+kTUtURQs852JJnDvaqyOExiJlGgyFb5WGFaFyr9MfJnqTfk7irM9tf/NW5AnFv
O6F0sOBCOK33mJNgmQf7W7S74dmfnBfkyeWrw0FLduo8FAZQSroc8t/Lv6Wa0ZzI
svO6xLG8JX7eHacKbk0jgSNzSTgBJDrclzZO8N8+F9Lyb7Vq+UuP8Phn/D71SqaI
W+ahLlqkhZRDEhp3uksZJ02wPZxWj+DnjLhQ4CFowFjH3+XYaH53OHOkzqrVkWHD
PpmyzqFk5q8Lxnf3nc9MSAjowu5qWwumHc+M9lTN9EYclAc7OS3V+9qN3S7yMhe0
oBtusHTDvQ4ba9Pi11XNzI96azHzAA0gYZZZbLOVo7sV9W5VLyEHRpBi/yzZnPIj
txrtVgpjhIyxRFnV/D2rExq8FIu7ZwNZc0PuH3N+C6/oZ8R9lZsupt1LZE0Y22hp
89apXg7HVplu0mFMr1/th0oehbUEzmseEpO/bP4zuvHRadTGoc5IBEMb0g5Dsa4P
XKlNV7z00+q5Nh1EeekoafM3GMVQMzmpudNRU0HXa76WR4gkeicJhYV3J+DHpLDi
rm0sxzC7IoEiaksiamxNZJ8wgu/rrlrbz8EB1gEvflM3x35m3IF0iV2K6mqxcEaJ
1DaSNj0D8K8uo/VueAPf5kwp1e+sBdHThcQnYpBachNGq4aKG2DGnJVBYVSsGMLC
RR81ZHj8BmtPikEjltx8lqOdojp7sD+sdEaGAnNtRo3CueuVV3qrvzN/dkCcS3ra
h4QnZPwBzNfZjgpV39fEhUYaQJYC3xI9SVXK7oNGsBTHmVHU8A324U2SxGO3KVFt
eTuYxY3CdGx016tnIhCDo9aogo+UTnY1WHL36yBVdPSz6qkQNKBEKMDkOuny1xg1
e5WWUS0IkBJ3U//OhU6yYfYgBc36c+nnIAL3RTO1Bxh8fwBsc/A5L+2kiT1Hk2df
MwpxEmC53c7czwV16M++EXA0G0aosoU+c9OMxTv9ZBm8sAVVENuVLmjjT4mOS+oA
AT6XCiT6U6/Qg5/37KwQ07TJKFdhuSRisQW71x5vDcZF8NJGrK1fGwY5Izpr57eB
GSiqPEw23hn3F85dFi18Yjt3YCJ84AHnbEQUVo6M8oy9yjNdR+WUJyhJaJVEr2pU
6A7Td1uGLV0sZfLGobK4rvsNOlal+nlVJSNhqyukH10sZonq/WzvGhGY9C6kMLlh
Zj0eff/WeRAQ4Ir4wIbNtuPF/H/3L9cqokXnaQguLhtS43rHptyPcNdOtADgsJUs
rGEgs7Jv9qcC6raFYXzCB+AQEDrWegWNzg6nfT5f715x/RJfpoUpH0s8kkYFdogh
U7Bi0k2NV43qClqEMv5JwCa8qna5zdBwde7JuIMBVlNNN13ZU9vD9Wh9ICHJCVL8
oiEVPFek8f2mRdHHx6aieoaUCxvgjOg4kCu2zPbnlcGPu/stuE8t53VAMbFPS3P/
XavnD9hJRFRUTrLVMjIg+xF8GoELl+/i+LB5rWd9RmtC1YcHg7Q1km8fpgDcvxO9
r+lxAWoQnFyYy4Heku9nqqWviQLHVIohJ3a2AwQBqYtQmeQ9HhQZCbwIzTM/3bfD
zaC3xFdhAlXaMbknJIomOqfUfSjoQpxiNM7OMI2WSnf/JMEh75e5LiJXrj3fOJqX
VnNbGj16wsvgA9jz6Ef3mxp/KM5rxmF0ni9a2utvW22GB0Euud+P0GstX1Jub9d8
IX8LEzNN4tep4nvBc3bjFqZBfPSDkcKwD338RU4DlTJz9ufJ4qnE0+f0lHl2TRsX
yGEcb/IxysJcerQov5VeBoRbhMBQOUHSIVkCNyWdPOPzcARVcZB9DyO/ih1GjW81
ZYc/1uK9vMxZXYtryQ+I/hHuNB+hoWHWmID8/AoS+b2N4otRn9BnYeNfchqm3vMT
fXiL9AR658WriakYJQHFPW9jcoCOC4HZItlGZ5d5qwtrSaubFBqyLxhTCsorZG8A
CpZRxkJf4m2OwewyQEplXGC2zK+QIAoowWam7crVhu7BkEc8hVE8gdOScX6roZ0e
BZuIpGg7r2dp/+S32lJE0oBeSKYCClViMbd9Ajxs8YQTe1axc+sKggldeDHd1E8E
yubY1Ogtoea0bx4BX8ZGFnRUXKcZtgwo/pFZ37ZLQUJI6kEhKjcaebTBnEALEkhB
XCe7VP1SsBigAZZEi4QqVAcQWg0+3EzMAcQ6qSf2roYIJxv0swEoQZXOI11NIfvs
2cITiadFoK5uKyvjOEbdchSW4UftPx7H2/u9HxfIPcACcGKNAqQdV4Zt/5Ew63EG
qq5Eg1CZNLTfTaVPyzxIrMiDCNmlILwKV6IzGA3qoNqIJoIvGRoY7aGCCWFbaXbr
uXE3lctzbsgn5SYehDBmps9ldzSf1jBvJicgzIbHdjZRwWHuTIObm/3DurVsT4ZB
t5NX7wW+/WWrEJJNaJnIpBAU3Dz3RZ/yebVVubmBmSE2KlVwP5OX2ocVZhHbt+zL
HYq61QQ5QlIq/uHJDEQjAAw+K/28wI2WtMT7GYfBD9PSlr0tWD8eHPv10efsvLsz
zGZu2jMAtkGjkMyRXhibpFVP7jcBy834ttRU3emr5Wunfu57m+P7iyFRfBsdG558
sTHKSuZnrhBa2eqqtOki8Ipb91ptOCixk/kCPK4/kC83t1MGRBkl5VRJbeKCuyDn
Zsw/3G9p2l9RIHg25JlGl8nUwB3PgC0+MnP7Xr+pFUm5AD7ajKOqzKIbtxUaEFvd
J06nszrVYeLKxNrw9amgPjCq3C1GIfL+gRhpnGCpUs5Kddq66S8Wzsh3w7ESH9/N
1am+adKe7neMX6yFQfwq4bz3b0w7DUYfEk2A5UmPz0dnA4ZntVmexFQ5v7MNUNBW
eJ5lA3foF55rqeHKyoYc9HGXwT8bRgh54R5NHdsByeTKHGXj6cXR3rXbYQqVn0iL
C/r3234Lt3P41XzOBdUZEJjmwUXIfMjl+povt5VI24h9643G6rX6R7zPjU/9P3l5
25VcZXAf1DY+pTstghpaPUtuDEDTpg28c5jnKd6pXMYncp17axSeGny5jZYPD2b3
fwaihZvQ+0/Ric/j7/PMszKdXCyEmoxTmlU/boMLx8QEEqfZ3qD2tx2rhmEsGyYZ
lYjelL3vDvanTQmanPg5DTmYajU2ngckVNG9NEiMoq8y7d24Vs4lCpqiyJHLEThI
x0BsaUfws/BsXnwrXvE3J2sLcaCS9K5hKGKzr9wHbpG5/w5jo5xGTDFdSjfo+tiU
O3ij0ED7Ipz10Nz9yJ5qGkqqvHFURnzIaDvovzQBFjADH7JhKngc/SgDO4z8r8g9
79YMXfGhmmrlmHr1N7KW3MUV1eXxwoFtvyy775R67WnEDXKXlCkqJRS8VlcQSWZM
bpmgzHsOMioFs3Sc6RC8dl+QBtBgrCR341c2zVzRFwHlhG4bcDueKc8Xa2fizWS1
zQObfawv9G+7zsExER6wcPXZdCD9yh3Eil5qO07ACHd75qwsEsLLtPi5uaRDqam/
rXMU8qi3Vedd7kVXsVj7B1ffiD9WMFajzZF5CDTd+dIM+wPaOjpjIALLOkLnw9rA
r0PY8DwyBgPE/vKsipVI2+GBPNvn+WYYqBK3QtKi4QF6G0iREKlwr++Et51pi8KX
01Nrxag30O19pce5gtOSugRrJZpA6FJJRidxHQiji73fdqUIM+NxIkjthvK7dkg9
a+1S+oAwf7kKhmiUB3xsw5CFKuPKoqp8kkPzQ1+edisi9NP/QEwmRB8c+vzPKlOe
0PypOnMxRqWRPjDu/5iAtFqikHdBnIMzTJGoE+Nr2PaiZ6B5cpiKC/liUjQoUwRO
JDjUjQsnLp2DrNnO7Krv02omVP17kSKs6MF5BOhj8yf50KcRyeb2k8Qw4kUxCAvn
Gm/h7tV5vnL2B+HVxFS+/Feo4k/urYe4RiPTkSd4BeIeboSMi3dCfa4mvg5hS62G
eetk8jY3EWPdzb1guN/rtWBOD82Z6RIlciMFHI04+YwOLMefOdVDJQjiRzS9wkIX
jgNEh70TQdwrh92lGHehxxAgnTEXbrEgg+HHCJf+oxqYduhwcdnnVEAi/V29S0KG
2LN5GB2HnddP4aCBc0EzN873RvBrw/9EkCEW5Cetek/DU5z5s8cibqksIJnw2z0i
DgI+a42xMxQ5bRK0hRLySG1gbN5f02s7iMnmdu01hLGpFHGRJK/CBAOw2qzDnG5k
LkjEKnsRRna20lPsPMJ2DGF0jmp8I1/SI55SqYINQPll4rFRW1QHRpjVr+m+2bxD
ZHb4QTAnTHIH1UeMIxPWkLrwowwH2St4Ywhcc1yMTKSAlcg3TJgfqef5g3NRkkLO
YpJDHWbnEII7Y6UXNkxAYlOGEFJYjRSyZJJxxEQnUw4HusHTUST/8SpAxt4zJsUI
0jRLmckedJs6oclhc82VL9leXcNHe0K+iYZVFrORXsgrSEELAxOyOPNmh3oQ2idL
ku8l+LPey3yYBa+iQ3B2hNczPGxhjznoASBtgRO7yCRXSn2AvLIKS0fCdTPfNb3n
khN0nlRfXM/pYniecLWVFmUB5gAe7a2kW4GRf0VFuO/dlyAyYJJNgLsn63HEuI+H
cFSaoub2R3fwlnUhS4uivzZscOhSZgPQUyVdMGxDoK08WmALY/CMcblF6vANNzdp
FcTiD2iDHQNZERKnyUdSYKDUIJdke5s4VLxN/k80burmnysgNQZHQE0KKAe+VpSO
wQ3ch45IQgGfUYnvQxfiiP5pB/l7xPSi+mu5h+kU6gbDrmh9RcFrZW5AQO6x5KKE
dUfd9FbBJLD7YCg7IULGDaR3mWXJYaEGOdr6r5iuDqqStwtKlxhtEJ/fgnICRCq+
9MZ4kifBGIuDmc4qp6ScGI+C52wtS9yHwej/tJfjp2c23X1JjO3JpGgHckuWAfeM
TuDZGmb8W7UVST0t07HK19hf5b4H7H5REt2BwHZdSS6pxGuOndWNPNoaOb1F0tNZ
lMBnApSMRbkYocofLfnMEMYPsxfV4Jj94Ubv/4Lcj9H4zkFn5yFpWpE4WmkZi+WU
hnLL8nVXzeJ6AkZpt4dDhtXMskteO2YJ09yHAw83WEVdzyKx5ZBEJS+lJKb3szuE
dyqs3/JY/6zFAAxiDn10AMUzXuxAKyPukMHFSHms2OhY+M7aqn0fFmx4hayl0rSf
m4Le6Fuk4padhL/jruXm1wHLaHaUqHPq481kCF2vd1uE0yUXKyVB5XrV46BqLMZK
OJepYwbA0Zbqy6bmkM5ZYlM3vnNLrX6gKAG3Fp+lUs5QUQZARFX811frgHVAHMei
irB0OJI/R1a/jKncm4d5BmKQC8oEFWl5uuzF+1aqd7C2ZMReU92fr4/wcAmtazz+
cnFykrlQnuIjmEM/XcnTxItU9yxwzCy1MDe9N1olwcxZlruytZwsdlEMonQLc4zY
3UA7exMgWsuZzxpsBXe7ae1ivn/+8AQFq1LByI1AV9zGCpaMMg6mNjXX74iKQdfz
UbApe+GQgSRvjTDhZ3IfecFLUi1y8lN4Spj52L2qxTc7Ezn5hxbuvg4sgNHqxusq
AawbPwn20wQPlFVOG9ky/IWDp0gcCF3xqu0O9eIIBx+Xs4gt3z7C2+oQCopsAXl4
+K/CqUM5XKqCioWJve0M3sNr9FXzcv01KDtYzgnoiAj+mPUMkzvy5fFqA/KArk/v
VBcGq4m8+8sFni65VxR7EbjaEcMDMqahqLBbhKuCqBtbhK4YNnlZcSyA6APRRgDI
l/Zk01vang+Re/HFLdUAN6U88aHvRiMGhwlVinbme1EzI6iN24GF44rDSKQj3ho8
kGK72CRkBZMmCbsFk6NSG/yagGS9RawVAWZNMu8SXeMBzKbiV7rHSN/r2RVeHubz
4I+cSmVdwEb6Ux0kqXCGgT5bUNr9gfhC+gUjX/HmpPd66DnbPD7i97HkWouQPsqt
fR8/jYfQeCYxEzRmPoOcYC0E6fOYR1zeaBjizpiMdHJnOwop3UQNLlQfqir0++Eq
B9WdORN9raCiktvcJFHi3x72oV04C39NMYxouvzKeN6GhStgqor709TlpFPm7Fs5
mqbofz++sEeILR6c8blZzcqBw+tJnOeZfAUnFpmth6k6zTpV1ZAR1d3B7BOzUMSE
WQnmWA1ELLCTndkg8dWNjLbxtwYZHw2iPMjK/DN0DvvZ+v7g/rj3ZxDyk9c+lGFo
97qWLTzzwBzBGAknW+tqZp+JUi64wbZvegzQdSwMf52SKnusLPF0xF4OKJpD4yGx
AlXLyDsQV1ZUOjPlghuMUsac/8ZAa4KoDKFkiz4voZAnu9XIKt4MrTvuw402jky3
iZuFBZ1RPnVCwBQNU94eugNCtegKzUGD/NuA2kW0/liuk6g/8kPIMGzWcEILtjYI
Hama7a5dGsRlCNzYad+UbNVZZKWLThNQhyKtFTjT8wO/P/JDzvSKNGeJm3JIluo7
uq22HfGsrIkafO294Y8MJMZWvwyt+gCB5OPjIsufPT8aWj3B3Dk5XESo+h9HupFB
SRyfnpTnvBoqBrevwx89+FRqRK8vqnYnOo8M4CArc14Riog7Vs8/BgIAjNn2urVV
seF2UinBgxlLPVD7WnPlPejBH3T0AFiuRb49OWcS7utGy+RLI3TqccEe47WIS1wM
7xILdXHsxosX5N66UuPL7+4Tn7UNPqTKmzPzN5JRt119EPcNZj/ckree/CvZNPev
RVEMNXH5TDO6wyZjwHLNUTnR3th/ixctmbgzoEuf+FL4LM0SFYfE4cAj5wE6f7Hd
ZGYXU1thwxbXDP6l1xISPGArpLXzNW8gmhgy1CI91ShPLLxiSN+HNPFbJ7AMIIuu
Ck/d/G5KiZAs4yQGPeYnv7lZBVzo6MJ+xuiUj9vFSWXplvUqJhfE8A5hs5Skib+8
PUEVBmviPxJ04mSaBDmprvyWBLKhbdnv1ghQf9/EQXsmtKCH5LmOGIGOdLZfr77P
Gk39EkdXNfU74YeQJv2mbFBcYB2bML6cVMXSVVwgbkMuE5dVWC4zjMSh6VSbPF97
SjjFNtK9zU0r3Nt8JTg/6H43Gso8Tq++ra+U60eocJfO4exSo5zq6xauLoe9phfP
iLhR0GTm0YcWBpMpV9pWmoC4MV1gZ7eIPmbOiXs6m7h7gm5qtwwiJjBQx0wGvulI
fkRRUemOBuGHfbdFY8s0A3qDEhy2zs1v9ym7wCr71ltA0iPCa9pUO9ngGvRAJvvq
zifMqs4P7rqLr7PNDNiGnGXo4ZMm/cjccaPgiUV+czrKBcwUWIGkHSy6u5IH98Gj
T4EQMwZHBEahmuRZjJA/9/65jw+4WW7QUwEam9qEER4dqhCplxDWUPn+5N2Rvnyo
LKHnrMwWsUvecM7BlADSHgm/LB4xe0tNulML9SaPoaFh7dvd1F9oPxCcYShHBKRn
l2OurAg+LTOsb7MuHVWP2LwETetynmLuNo2Rquuyd7x7wO2EZti/zcmQVCAc5F9Y
0WJunH6hPeOQ73vuMKXl1kLskIjKHnSg8dhEGV2/SwKrQ4aD1T/Vc6P2u89TQ2Qc
2kp8Hx2dC60OpXlZR2eh5xGlIgwy4ogMofJC0LsSpYywpMy7C/xghOiqDq4CMW0L
bDGGE5qhdEvDrUomNNX6JPoLZmvwrHN8XMCCLs3rwWSXWoYkB5dKB79Tl6AMuYNC
iSBYMkkCBPeMC1v+EMguTdtrQ/43M6KBm9GgqGffBo5AyxKIzFplMidcDSpVSgfR
3oWrEZIfElRxVtI6MWI7Bfv3cpYqKz892Cs1ODAmGQNBofZQgg7giH1gfeTk/FKl
H7Ixo1K7BCnR+xABixYJDp7JkJ44HkAkbD5SjtDd4rDLJq3vabuQa6QCQaXpE16A
Qh0affaFHhzEObKoC3qR+UF6AIGAgDDpguTrJu/83IbwUL3vKj3R8xTKqT8hLSY9
EF5eMfEZ43YtsQ2jsKlxn9Ha+IGo1z6tUSsjEXZZkaE7GfokDEEutVW3s/lDFE+6
VOPHC4FlRQjcYwoSvxQG/i7WDr1xdLt7MzJf54nWAuEld5teyg2bjWireDjjJ77u
ed5Y4HbjWhQC1HRb1RrDE7b4M5YOYzT91Ix2kvlrUOelRYaI8Ih5x1HAmiuxt08d
NtGLvVIz9n2pKwX4UlVbVmc5iYMO/+B2PEoNvFq5fpG9J07SbCXpMZk5qT0laSwV
xil8j/2S6slIQROSuNxpL9PiZ9wMcp+rff28oCxI6h1MrWhyeiPnknlPVM0XBE27
NXxWmyfq3/QQd5y00I9fIJBlr5irTYueM/RF1Bn8yTCt+CLHFP8tLNtc65mqTU1t
Fp2v3VOIVK9RN5r61nIkDNaxK102q59jFPc/6iLB4Uyp53z0E9IkfXcUCHhRQYwD
d7FmYNmj0hITempULoGIwdA3Q6Ec+KSTtl1VgV0xpLoWceuiBxuQegI6X4cL+7Rr
9iBXPlT+I+/KGh5PBF0Snw7qB3pKq0hdULYzbyekMapv/YOk9VaPSWsYA6zxYT58
ZPduo0hinzq3ujJtvrCPVrMi2DJmxywm7c06B9HzQ9LMiTvf9Lu3VppVXdvHOPSN
A8aF0lrRNl3THl/Rf/Q+XKl5l4bphjEf3aRtEoC7wTPAnLoNc8643SCaBxXOKKJl
9D5rzykGBqZQ+4jl/SPTAB/ZKahINiY11HJERgtisyx33i4oMPPo5LkRVEfZ5M5L
A7q+WQJUqOC+gOrUw1Woi4srLcZCRkXrxB/U0RRLvN21nw/NPxVWAbzTFYG6swHT
jF1yTd74PIEnWacyxGC09gH4Bf2jrOVdo4AESQ5hf29trsl7FtwaIRgh+4utIx1l
pliezBcNQ1a1E8+O1mNtIklHySVXqCzQUrUwlA22q7utuwFvNyu2iepkaV9h7Jb4
6ObEKM+XCz0c/sGpRpnuymj3OxJdkHCEc0ozRdWv384voCXm3KZnuKK7w0mCDCJ/
jQpd84aF9W9EZB+rjyQ5cSHCGrzgIgIXApDZ9mktkb1VvwpJIRo34hWzcNT1Wp8w
3Z4gYokUgSCyhkBGPPuVLgs1rEAXAiseHsEvb7j/z9YAg+BCbayQwhDDo9594K4x
iS7LfYDtt6AfcrsTC9fPFq9lMNkT9rxKCojyB7TO4dE4d91zlEqSJgCKMzbEmGz+
A/BvPvlQ2z+5qIp3Xp7kNT/XcF6HGJ9+/6rh5pVlTLnPih6bvEcSZe+njq9CM/Gs
/Chdac4ULJk9+wxioBUN9uU2ayBCb8wxB2n9N7AqlKYKoJScyfQwr8amw0Fp0UO2
9FIh+Kww3NwHObzLACQNTDMKq2ZnkXIDCRR7JvlLtS2+dFCt9sK2RRWeLFvWmrXU
rGMQr7bFi7oPvpP0WJ63RM6c1KZnraGtqpKYvwoNqgbyos65Uj6AeIBegnCr9Y5n
ZpSHXjdTWPdnf+zZHw+7dt62gRojW/B6Mt7fmutbPh+327I1JIj2ju1ZDIWYUrbR
PZhkPbd+/f6FCNQtlvBldVctoM6MqBqxoHVTpWoF2KCiYmh+894Od3Ilc2RSwOIN
sqpxntVcMeuX8IZP79MHXUuvkSzML+ulN986rS/I04vE1f9Jlz6IKBZf/HJNUBUT
0NuC6MXNg71d+ek6Moawc9sHRA1raaTyW/Cdq64TB0e+2o53sVPrqcoy+QJSKwti
4alujbJM7853/yHS9+Gqo1ntHAmZn9yiLKp7r2y0TgSX/znZLm4WxcF4Wkys7Gor
DnsbtmXTtz7tX65N+KQBczxZ5o733gv2dhgDyCgXH59/v/ADQqCa7T7C4JQA3bra
p8ho3RWkpo1koWOlntnCa0wFIb8EL+ITaK7Vl9tnYJosHG+r4N9OLTx+8q3vFYpp
edoz1IhZG4kx467xcMxbOm8Ka/ujfBwpXl/DKesViheLLV9TLURo+edFjC3DRHX/
ilQTpqirQKb4+j2f8cIoDLbKBz0NFZ7wQSts3kgaVSL1L4MIuFf7+kxiBUH9i7XJ
6IvwbV0dONl0nzMnX/G3e7QIPVlwK28kn0dxYAgNlNJ0CwAVHK70wACE3lGg54CW
tmWEHSseyR5zpd2dwa1dKDyKJR5pvFfnF2yD+v8Klz0t4CEFk6+28mwZyrfT8NmW
ypsC1CiGaTftRDCHFd55F4OcUeREOuweHVvanrE5xPdECdjPB13qd6hkWZ6gre6U
MdiMbC0ejkvG7Nm3ZOLC1DmbEPOea/h4j5j6K+L6I+hXDdeYvypVVMI+6Trg1jfZ
JNgMPSzSf7fQMH73ZlmzEVBygcc9LjGRBU4Bw5OYfcTW0gTskG7DQ2CIfD7sdiZt
wKu6zE2wyiCWO1UVmI3gJ5nzIhux1/rnURU3/7/vhwtEvcr3wL5anWro+GJ2te2s
WwvP5zv5gfI66XE4886mlfCuz1VVenUNCpRPUV413LSDe3XF1a5mHPDciLwBtHDg
PH/Qfl3J07lGXR18VauE4Bh44e+NZ5ftGS5mu/46NnD6f6c0WOTb2LA7mVKyulIr
bLihiP3Qe0WBFzvcLSU2h1qd2PErlzsiJv+HPy8VPUFD7HWCV8hiU75R0GaEwiLs
6vaeWYP/TKzkGzMAXt9IrkKHxg29lYxga3RFptRTbCkfCH5j5DvwrxyKyPB4hp+L
NtELbVYnd5G/Pw+kO7CeaJM2o2tnTkDpSZOSJ2fJoJIgSeM2h1WOBM9h5TTvXyzn
Mt9YgumeOXq9wU8Z9LCaFNHdtp1zS5ot9xf12lDSD2uhFwhZSGaZKSRkvO9AYiDo
bG9UgMOYw9McgBQLGFBmtCSPfSxjylHeaK02WcZJZGXUtfrUk/sprr9OcSwXCywJ
/4UQ0dFeQGQAd1UeTTtUaGP/mtBJ7oK1bYKVvCCux9FMglhIu12XZ/h9gZ24+6H5
JouOpq3qUnLHOzM/bpRHaBfQzMPYpCvn9NC52tyLNtzVi0lj6Pj7BbG1i+DFuql7
xQe8/XZusqZLxuDWRXvw3DLnQKNluwl4eunmNgBvoghYD+SCISHhTdZI9NoA6imM
3Olgp/Af5it/AfFLhxy0fOghQt2wrpnIu8ed+DCQ71pTOfqmfVbsiTRv+zwIfs3k
FYKaf9ydttvDCYzK4ALkE33Ss1k/70+PcZZcKc/QVpzpnfLwBhcSL8ITxBPoCq6v
JOkHyuREiwCPv/wcPUG4PeJro+GWgqO4wVp+sN0RTQM4sY0mrzoYkzgfWbqdfY9n
vLM8rJ+C+AoebroErIEry8C2sPuXX7aw6F9kUwxaw/8+51axPNqEjtD/nv5VPUws
TW+4TXXiblcoh/yY1fMEDEkTMbyk6I7tz7xaqOh2MWI5iyatC65tc7PZMSAgoOWw
GI/ve4ufSnX9O9KNI8d5CuUrqBucqApFLxLHz6EqxkGhYJBNQIHdKV3yn20/QgOH
YS+wVKDNDpyXKQbGELoRxqh9DcgswFKUskZDjV7dyeE2n/CheIbVJuQDaPw+SypK
lD1LI6cNf6B75ZQaKppmeUz9MrWc0vhqfA1MTspiztfSd/q8uofX7gLcaUHoAwYz
E0nhYLuUhub5MeCVASI3u5Cxrbl8CfJ7pu6s+joUoL3Okc8irpBtCesk2J21mO95
6JrmglgeYJsdbmN0dvY0rzzLsPCZpkS4t9F/SBWfBmvWHg7z1zbMwXR77t1U5qxj
7RC0pUCCnLUTMxCTvLwE3wEWrmgyCMMK2Y91+XBXbF7p5a5gHJyDjICDdCQga0rK
8dX6X5xrwAcxYBC1V/AZFMN76Aufd67hVWXTFdAITXzWjy4hsCY5CvGJ0FYD5gDF
XV+VUml6yz4sIjlUZQ6lByoDcRHtDgOL1zE6QiCnJ0WjzfQd+fwowasqYLM2AwxW
xEorHoqaNvH2IY+GZuWRGcvzZCJy82y6TuDnz0UYJCErrzLDxmSVRTO9PxvvdYdq
c2Im13G6Y1NvV7bTzpBBdIkyHT8LnGzpDUZfoiXLBymTp/Jo31866EYld+EWPZWW
TzBTuNQ6IBygOJ4foA35JGvy+57MR1wtpBvMoXuYCaFY+hYgYUanLibZlPKN4fvS
nrmkMLKwN4APviM01tSA/b/WzuwCkc1dMBOWka57NjSPwMhvVxN91GfX2leMgrAS
319MVwoWH4dKP0/Tn7vzOHiRC2z4C6GpNeIZYV+vDIJZw2bqCoY9M41OvdgzInd8
3kiZC7bUJvinFInjH7S8wJEIDEKxD//OJeQXBPpbj6mX507EzvSF6b/fV/pC0e8M
yuSePbEGwwkrIZ2h5Tdlw0/JTC4hDaI+2ceoLHJeKfMmtsryPASlLCUcDnWabBW5
4MoGAmawI0dx1R/2U/nE8B90R6REJojkiLrlNHuCHGHAzKW4RZMOmXz3FtzfoV3F
jpXJmHVyVF261MALpnfgPLSzyKT8Yh1N3X3Oh35yk2arL1UrR5+D8geJJay0t5f3
e2MmFol2jnREwKCMjlgMibat8ChhMn6LYhX9XoNRpEzh4/2ZmcTnPSCyAGwCm4Pv
0wOXNt2LDXk0Mu4zhBLbtL4ewvmzNsbNFSoqaFmnxPo6c9bMuEGnzTDmXFv/xk0F
djWMm+oSylcDQaIsa93AuEue+pKrg6tule7jAaRlHVCDXopaL3CE5sw/z1JvJj+C
4MPkcxPE2A9lJo5o1++YBYrvgGTC78msznMUrTrz2IrXfuRYoJcuWRK+anPZZ7S/
5u81aTNGpEXXWrGhC9nlaCleD/AOmCH8m7kVi41GvXYN1LhQD33bMBH65xxViz8C
1qsJKp7AC6Yp8e9eeTBgmFHpdEu4KOB5APBAMK+8sRGf3D7bxsnB6LWIlUQjRFJk
dO6k+PEIcz3vue9kzeJsEFLKIQmfd8zjqf6lqrOYDqLK1yOHpC7Gq5y4uHMvikfU
UTsEoIaaz0U4AfRs2xxfOugOx+PzQhQgYIC3xNXtBTwbn/c6eymbv7fSpFXdaTm1
ioo5RifTPpsTwmKjc4CM5VbKe9XzxFt2F5fd+m1JrvVT1VDMrGxIPJ3pdczQCEMC
J757rwfzW3OTzPWYBQEvz3M5P2c1ux/BNaC356VO6Mm1L0dzRL9iGIHeXBszRweW
5bbW1tv7xAUZ1O4MfQiDMTCooYdpiRHRU+t/RUaGu0BqkIVxiKI+IlQRmpSJ7Yuy
N5bzkl5dALjqDZ+cQufkHJhcYFW/f42MX3FEcq/6cV2DmaKrrk3W9+FGsOqBiQI2
RLSOGaO3YaBOVHz0sQ1bg16DNRJ4rg8ERY3Lt0eOzXW7C294kCaOeTE+U8Jgt+7s
+rolEast12FGFrPs/VJLTlp6G28gwHd3CC6iIhI9vM20ZALh2avKjPaUKSeOwPLk
TPcLHIhibOOlpjS4eZOLBDiRrvptQ2npR4fmrzs9u0nNQb7ydcpvrCDbbXpP6WWq
JR2lkEcdriEORwCwqV4qWHnIi3auCc27qsVMGjdExxdfMysmFiVrqyKnDMn7K1Md
G5ACTKjdA9y11i6vLXL2YjkOmhLUS/XwFTlY+or9xuJSH7zFZgJaz8MLXxA+U7LP
0TksOP6dSUFmPuWwfTNjItA9wWh6XDvn4EL4uDpdHGsrgvGWEg+2319CMCj0JRtZ
wZChzQ/9k0Sjt+DQTypAxoRTguUUyLTO9Cq591Vtpn/D4l9NsDZ7IbEeZhNjRWR0
3QL448Wvgdas88P+hDzqN3oGf/VvxGJK7WgIA3y2Ha/599emdINkuwUaaJS9g8B1
DHL7YRkLi2OYIZKeKpSB4fHdF9gTxqdLvfhQToPw//rENn7zkSXFs1IyFNe1Ui09
zlvu4nVTQymhSdH9TvqdDyNdSMF0Xqdunw1MkpCFioO820tWpLDLjrTLOo+Dhj4+
KylsjHkZsZ2xcQbz2zPzDoUf4Z70JPbS6LmB7sASnhIZk2hxvx4mfBK1p5xFuXDR
1C/Z7mkXw+cH1QNQs95IlfIgXt6Ag1gdT1p29pDuzP0D7TKgnwbyjDSMgC9iSdrz
sXqN5PGSnHSOIuzQLoTR5rOdG/w37sKqo9X2rXRuOP0nCSLWwBxNbPc/GMIjwq5J
NnsBnVJ778j52V7aqJTcT29dLZen9wjx5nSpdAm9yFP6L0vxRIYvZ9fVBsZ6cryW
kYTF4cu+w1kiWtYu06KIUi+kTa5FEO9ODB/Ej8l4FG7yXwnQ7AIGa3F8VWvmM30X
S1unMDQdneQJ3RK62PCEdvbZlzayVwvZYG6ebRkMl0sbZj5pzbptMy5nzKgmjp2B
S/WAcGJR8IWKS6N20Q6moJEt90nxWZghfyrOjupT5AR94dRiuPkRxKS+a2ciGZl2
KoDv7NUnWy9ZIOxQ7s3nAZUTQaYq0WmjTDZ1V+MyuSpUB/AKMKmN6oZWNo8qGAKR
PRz0zw9KZe1+goZuXPkwi8iVkGmwIP2OticOzKiruRlYZy1rN4QVNahEhCKv79Ch
NOuioae/nol01Svcssteo5Rc97nFtiLard91gOiZTCpFSaQ5uzgm/yOvCKORdA9n
wp+XWEvegi9ZSeK+8JiiZ9JQsRAw8TejS85VVKhqcZzI0lMNO0CgW1JaAY1ofCHK
7HBPOYnaAd+Su727BHog7ebxpxOXPNGnquUvnKOp0UNZes+Xc8GRTyWHcbZbPsjk
jKdgmRFJGWu+0c9YGtpgjsphtJjpq5pKviqrwilvqGbQ3uMWoMQZ4sS1c/X7QnRy
Xl/ih/QqfpH/+NkIjl+Sz4j5BJ1zQCNrQQD8yLwKBDW+Ud97s7fXq0KxMTrxT1EQ
wugty6QUR1aZC9kGL/7flX/RXVDD9VsncVeHNBM0cc2wOd8axAqJ3jrogvztQPeY
56exKRBh3Jta5Kx0uxZIuWIu0+26VW7UlTcSLu1dAfdWk1P8RUVFNL0XstHHf8IR
BkzbTQebJp9cbKp80hAxf//dzindXmyGPaG2Tt/K09QxNXq+nO/2obmCgkvEW2Sm
0lWKf4mur2w4gzBD7LVrNy8af03CK25y63ZYULYpyUcgQG5dO9qjQL85e8dmcQlf
zsUUMcAAOMdIHBULkkoMQD8Kjvwl2EJzMcq508G3Zz+rCjZT3hzfpg/TPTe033zs
UVco2AC7WuCywFvNJHI0QAMK3TDVs9OkDBL2NMJ4epl1ZruF90gakkgc0+KonWzM
l7pEVrFvl98LL83cEMhbb6R5Ycc+ZaaaRtupBE1hE7hxxGXd5WbR3XKEuFiJe9+3
Rbq54su6ZeP0TP54qcOlETzYBj8kp8NTYwsAv6COLPsDaUT8UVv1BFA0U2qD/kst
xWxsn1l4dZSLVrAaF7tPRTjGxgkpJNeRIplGVQ3ZLAA2B1fTK23/XKHp7AJ85nky
nq7fqlwrHqnfTAydvzozpwgUEoMLYtyuBCsgvLuApZ3JQGWDywZdh6+kiVwDhKex
X22K6JfDYlz6Tb3sEJM69AZG73EjJoFfGD1OCYmTZ5+Vb+cGjL0bC09LxwXiObUp
FrZoGSv2sZ8ZCOmu4ifkNM61Jpxq5WMvglJqOpkVzlvQkYRJoALT6eb6s1W3gMQm
wF/ax2pg6V1dq6GY6X+yp9CSJJgnWXguc8fM0M9c5Tu0+5Xufwkau0JAUigz8soA
CdYSWqaemRLGThkw5SONnoYyeq7J/i1uwZChs+SpPXvspC7Op2LtHJ1aHdjPXvXN
92ncd2zKNBUF9sN7X7nxoRzHNhS46ytE3+iiJpkJfrTdbohVXJZqBJqXpZoucKGa
0Xm8Sxsqrcse6/31HwrzEY5gFvNnQzXVpbp1F4rgk2Lgr0xBEeVtSI+RDRDj7equ
aVyeylKuIDtQ9A3jdCGKbT1nKhmUn/Q13FwTUpLikgKieQn9TRbvfHeBYvrQJXaU
MiDP7oDet8DdjPS2px5sOGRPzNGi/D+Gg708z65nqHbhUZ0k9IjEUusTXsPYXZX9
j/LoNCoGHKedQt0rXAQnv6C4ocv7vG47U0NFNXntl1fM/sBiVERHlUgCWN/MJO6C
0EQ3Xmhku2/1ggNqpenTvmKQyNiDpcfvxaBqDuOe3dN6BlR2UDmgKq0BPDsgLGuJ
VOOXh1OQTVC3o5Xf23NivSPIeNbbBOdp6G1ktS/+Wq4sazsKXbaidei3jXCUtCHT
rd6Pu+9gX5PG/pPZslIPHG+dLk0q/xuKpL9x1LOBCSw/lXtz7pVtDFKDsX1Um6ve
LeXTHRdGZ+muWdrXe2GH0MUKtQt5gG6POgHSQucnOsgBgYx6PqCI1F47pC9674sH
uF139chPd2dkPlLx/0i/Yg46XLt+0xk4+U8i0d5PJwX7BVSQfyMeUBN+XsfGNluY
gHxrgHhaJzmBjk5vWkssfKMBVT9tVCXKU4amDKE2Sbqq5/2uU5m39lt69JuT72wk
f6QhHWrtQ4hhMg1+n15BxUuz1yEHmNE796D3sNIv5E6E3Hn6UGCxVLmfw4LCAhQZ
FOxXChPfLixvdkasKnd0WBerQTUH+whvuUDzhDYXXgMiyxUapw191YTmpM25KU5i
9hL5xnQprHRFyXNkR7PBit6MFi4zVyaVweISHIzozoVUIHvGEAzx5ZEiwp+3vmxQ
1k4GBO5tiOnMGqZZ6NLT0hsXwtFeTueLzJxDRxf46OA1/QHYn8v1Ady0pmZMZPu+
rL9/LpCNJ2p3uqjKAnSJmRFzQix7dav4DZLaimJCxAqx3idSthaExCSXCjpo/f5o
piZvAPR76B5wYYOnO/59NYnEhPH/B0a3bFQQ+mvCSKAg1Kxnqfomn0vIiph2xufO
c5/jOkz8/RTSx/7pD3QaHXCmz4DkHLSrj+CdNbKsahwpG08NozIJhcV2MrBgH6Wa
fpTprqJuv9p6HQNKdC87hEUxwYeHfdvQFd0PzPNgv1w8hKM8hIlYvSsASeQ21QeQ
fNbyVHJoAB3YcCebQV2OfFV4vsLFI5nJx0mhtWt3KdfH7F2eB+2TDianW4/ZsG2i
7XYn7Od1MPyNrR3dVz/SRTxbhWrbacGgqfYFRWrc2gFVN+tCN70Bvsu+zbf42iDj
u19aSkg7qWIG9O6crG+dclLlFtVZJJAYoE7rgKlVwD0+qxGf0V/g2f0Kp0OHPIHO
ilEI0ItenUqMVFX6b3mjH9gvYS8NOva3Ux7+v8r1Syziic/ozDAYRxiNNozyE1ty
TQ8ebqy5tIXFyhFnRi09Hru+FMO8byDaa3XmdB2b5lcoekkll4LkF+8cZV3obm3o
l+4/Zktj3Lp9OwNFzfuIIEdxbf7B6mrzT+I8QdaFSob9dm/etUQZaqnDUu7hbTDJ
bIXuE8k97l094ufoealekiFGjRgXfJBsSqW5QGiCz4ok7pNtI6LAyZX+uTd1QHdc
0yDSGqyMJTukp/fBO/yR9bO4u29T7BtHk7lZzmnSIzmQkbOvZC9n5LM2EXI0eocV
C7FobXa8Gs/rPP0pOXtGYczyoWMzwMGaOFpM+Pt2obEfeaoVSbQFYm0IdI0S30/g
b15ALFHciiBp9CZOS2BGkFmj7ASJkKfkUq7UvMPlXD5Zwn8U9IxbFMCrRA9fxpUc
aH6shJARX2Wq0XluLd6auZSnVn7n1rOYcQwiPxBRCXSo8xWrmY2ktUl51aENb79c
wpP48BncEPTTvBAkW/uuAA96NkMSFfH5cAN0xa8SX0p2NrGKpIGcZIAkYCRxM0fw
oRSz1s6GVTgFAaKp+A1OaUfBOZKdcXLbzzYzoxH7W0DPHs6Ci17lLBYs29l//ySM
eI1OE2uHFRvwyhCoOJdqN+UpHaAGhFoXcdGCBQbBM6/LtpEAKVGGMs3y3MBocYzi
I8edKnU+ReCHcwXdq+9wtefw086aMijXxv4U6I+SgVz2h8pMytaZyCAdsFwFImGx
b3yFTF+hoJXkfGDwCrYkP7ObftAW3/5ytLHZDMGIBC7jQlJI+GZD7a2ZP9FDmp7b
56YQonIfORaN+EVpQz9mesTo6FPFnP5IUdiZWWvBRwX76w5JkLBQz3cbkUrjuIwr
3IQb4Is1/mGRiOZp8PG7skYWVQ81fslJloCePZgxfl1+OaJrFHz13flzele6bh5t
dKPGawPUbl2osiErPVc85f+TapfP2LYvk5gmMxxsb3inSxGvVv9mGh80kd7VvfFJ
KNiNYfM68XiF9yQhH9C6OpS0E9uNAnBOl5NloUqgOIBXElYEwGEg/0uejhYiykMT
h89oNrrjb3u3Bz09VYQ1A7JxHshNjV7zJHIsW2zGqW5nMCNZeMirg9xCQhTA0vJI
sZZ8zaDRZW7eSm/p6x7D+QOOjwxKqd+ZGzwbvgnSBx3JVjQKtwd+E5yQg/clmlbQ
twVHCQU3iB4XttsaT3Dle49niIktPPmvz+U2kQod4WA1aXrhgNy9TuCFPcR+t/DB
mFZMLMS3PhsK+u7yIl1YUry7mQBnrsSK42vGjLAJu2fpShioeo+ridq27fsMGpuy
BlLbazNf7cUy72teBhLQ+g+0yvddeKLStXwa/99bkLLKY7lxv07UaohpQalAJI5G
8qekj26jncujwM8xYji1yZmWMwwv/NqxEvODONDAtT0c46S22qEdteokwqdHcIcL
3jwh38IRkM8kn71coHQBoaCS4Ga5jiYUosQvUVOVGvz2Za72yvUmGf9GlbrZudDc
pH6rTNijTpSEYKUDU7EmaJE5/g5jb6sVF5kSbiY7+1O7iTr2csZvyPd48NjssOsn
f0mmXYFOa/aeTfmUFbPp4rBKjxHhhp/E/I30m9kr4NkrDnGuZSXQV3DRoeELKJto
9a+qrpZcQDqD1BdaaLrq+q+3MDeC+l8/3EXM3Eino6v7MNWON0BDbJApwD58dzgN
MJB0nYcV5nDt2XvlQGnAiYB6Xe4IfFqMQTnF5jCi0vxkKf67i65O/oYlVD60VIA/
jnSiQ3SnxzZx21i7DGs27iZpDvafce0pZfoEwVRu7LodbSG+052LABPOPrb51I29
rtDimXZiHyDON7KZvUpuTbTQmbNYtzy5FdtmuV/nSNn984A1v1RXbMpwPle1rQ+8
dEC/DyI/KoCW6vfjxtxWKtiSOIashJDJ2IxiER1nJYiAaY3IYPPyMeX4OFAZUfMg
zaDZ3o7mSppEMRWSeUKhir5rcN26j/a9Lzt1Bw04j5mSPh4VIw4hfTuEZMqXJd3S
bGC7cNyLig2s/3/3HKB7RERj3fCXW1f2n39OAnieZ44OCKrUN+ABnUOwrlvGDesD
isO4KELGc4ThdCMRKMN8ZK9aEycq36ovECY1A/QVul3DTbaSHQ5Wjclh4qY+fG3W
ip37QLeJZKtUZm2Hj1g+Lc8dmg53duiEeLFb+k45tk9Yja/XaKB5z6oR8kvDOs7d
nntD4uz9adoGa9TEhpr33mez8tzMNyhmbBt87iluYIx+hUrXt76T0of+qXcobPNm
RSEYEbMM0tWZTaqOE8l5AyeceOpfQS2tyjrsJ2BD4a/6aQMnR4viHSNRkFfkDYUs
GkpdloWVAmqGKhVrjkNERxF24SkEbA+aU29FZ2C9upZqYsXPbje7ab+ComMXj+Rn
YvZ6cU0YLZ7wfDd3uUBuh12BLIXvvjC6rNFg0LP0aP9J/nMh/j/o7EUW/9gJxjNQ
mI7jW0Czbd8wrVROlcXyy4y+keXDA5Pz91/jWJeTmqGqwMec7/u1bIC/9ST43LX2
GeeLyhvE86tirc0OqKLgIBFFvMNnV6Nrd0v5COteP6E+rMafWm8nqZxTkxq5haHd
W4waIorM9uYrZuvqMotOGYWgXyhGxW2IaVb+lKCMt/HS2jRHu4rbod+wMVbd4fYc
EvJbR+iw6KQiLhSpTwBmniBQWGEg9XnHFdoOuFjiTf8N6Zi//dG10/epRmgcj0QA
pMwUtXcFcMqVTMvUthYTBPmbAoVvqVa8spxMOb4Ujx6OPp0I8Jh2bSWq1O5SQPBc
c5OEqDHpxFLuhFdGB+PYZr2nZKEdSZsmItl+FjRZ3gOXbXbln0tUgCHYBupoR2y7
SwBQf9KDIKZ6FczXHpH/IMlgOkl4hJabzK6T+LE9xceXIm8/fL2vdkqjCU/3ofNh
IkbbqkvFMSGXtKXQ1qG34XO2uwto25i1aXgOxH/XLCMc+UpT6v0O9uztapmOg5Hu
3YkZYdMGJT5ox1QASLDK0btDWBiqSdgX0wMkkPz8+MZTOabgdKmEuUFN7VCfRhSK
McUjs/6A2+XYzEUE88HJrPvWKD09eULRb/buxoNBK24WU0b3YC93pfchCL5tB0BK
GPj7dTaOqX8Z+9UxCwIqVPoVAWUkK3gjeKheHRCHbw1g7egVBbbv5aaUUDHGGSpq
tSOo5b5lmZ4PPJvHUbuMgsOsKDwYgGkzIpkEzAJ3z9Eh0c56o+QzECaGF43UgysL
F9FRO0TxWDCjzsl8WRjvevaTAHMLrsm6BnglL4VepBEQkXhzJW+HcdH0S/H597HZ
TH964oTZIVbuORLMCOpbU9EglTptUvW8GARptUE+j6eAn61nR+kZ7nZZobGf04ll
TBNwDc+yMMb65UjYh+E+J5p/KbuGCQtlVobT+OyIe1QupylZhJpg39CZ12xV3Xrx
eCbqbTz38JvNE3oBU7g399bghHtKT/JlKbvMlpMeFk9D/dL9WvtuMEtjqycxkGGx
kWWD6jdDtDQKEKVv8YFfz7Osz4oVeR5pSJQ2xAzNDPQEOVtmdl72klXmGHwCHV9P
vDbPE7xzR6x72EwjzZaFreAiRAuaqXnX7vFSpMI/wFHclP/+qYLfEjQgr2dc7VaK
I79LipIFJoJGA/2hsaTzmq+GD1ORdimss8LxoZA8o1J2EEGNRN9iJVNUBTUKKuUg
AR3WKX0Kw8htttRcyO+EZC0nFMCw1RxQRPQ2cWLkMkXmpaNX3fMxdOtdItU+vmCC
C+bUtKD/vXgyheqBQ0NA//dh1dRVhrpJICQO4UWA9GqOS8a7wfedOzO9aIW4eVU+
m2sV0yaVDf32qE7uYzMW95bhuXf3w5XxN7ObdeMxuBGWhLfGnaBX/nZY1puP16b/
jgoYJlME+2WfrFuwVgHKZjhU8/1zSic5gOxKGURcbhumQVZiwAD/k0t4n0D0znnC
dKDUMhVeVY3140HNsyqvumx1ZR7UHa54qqXrkvO/egnJwTe0OJuR6ypqB8Urin8Z
UWpfxBkkSIemlCrzovruFivWlYRoIlYt372OyIMw2cyCCAfm4J6nutnIMtgz2eAE
2kjB+JAwc1GQtEt7BwrlYspTFjPT9jMDuL0RF/ddc9vAYodSW1UhZtINIypYiFhH
/uT2Bi2t7ntpkTr6FlqQthD8tVxgQQqU3cfwuXhyXt2QI8Nkl9vydSEjRF2yUwkM
3U+O6S7UU4jS7TJgjxgWeEKiSllddRTeeFhP3ba6Dr52/ucZwmgZVZeIpPy6uRN+
JRQ+f/p5jSDZmEpLllTz8ujyceXY1sV+JaCUOh0GDpzFnFP7w2t58X/ZWS1Thust
nHJz7WmO0zLSV4fIb+Mb1uUFOkdF9q/ZJDCYGbpQnJh2y6ux9aTVoSZnKFfYjP+x
shT04VecoqgJ03d0SajsOMl0e88j22rDao1EsIWFpWAU1cfiCOFhj1hEHD3IpvLb
ZDa98bg0jPIHy998GeegJ4hfocGnHYQGExpMs95xR0IWlvEqj0QNfS4JGaJg4rFe
lGy8osPh+EhYSoY1VT4Bj+vsbIvDrj9Rft1GCu3TBELchq0WMGlvCGbBBkEyVnOU
95nsFTYuQCT0IwW5Bh23roq1N5/MTeQXb/Fk6GwWZkV9Sncw7cOoaTDgyo4+9Y6P
+R4WYAiV//OY2q2Oxq1mjYaSFkeNgOPDZm4S+VDiVdl8kq0E8Oub5KI08jMCxft5
ABpO7MxCQfesTBgmxQ2ydebG/WqRj83zzVizM8AftgJyrwbyF+p2qpo3aPwuRxW0
Fs8xUmXQ/agVaBJ8rEQIctr1i/VzErRqc5pjmKoLl3QjOEQlbnk7qOidQuJEghMF
eX1RQseFRZHmPIoqRh0HyJvE2pU32cATJjeEBPt+gayMGVLTGwpisZq8BMr7mT1I
mLKRV+i5vEdGpWkXIdGFaVUe9ORf9919VRCA2kv0RedQsENV3Oumj1tu1hBxhcA9
9DzvQDrwRYerMuoJf/p5pVy7nzipgMCxJI6Q0ePpqf0SRUF/VigjOE6a/rfMEXRW
hInJfSyv11zQFQAkGage/zwfkn1RKnSN/E0rQ/HMc4Dw1Q99pd6GhSPEXfTPaxgr
RrPR2nKyUNluRkNhpsnVwyUv7BDRfhnZHtnlbPw4QHhJLLh/pxsckuepTeLbug4J
tQ0yR6cB0cnWD4iBR9tGp6APGsR2VjTbhu3OplD/285yRZUWI1gtIU8nVotqwDF1
kVZXHLTX8H0Ve5kwCvKvMZRK2+in68AvjOgJJHYOsJk3XuEJeBTuYhHR6OHQ13eX
sZjeAtMcKAIlNX32rY+62NQP1mrfiUaq+MQaeWLg0CY1+mQgBhn/RQ7RWkDkOx+T
luJITMlcb59fxN7fIIAE8WpYcFIg/dzEqiL2H1jmbvkQ/e8iiTNiEqIuV6nGOqSF
p/CNE72stI+dAJKhTfe1qyhh6Z068oEebzcZEgT6DmGRQW1m2KZ476ObNJ8nf60m
tFk3D0oGfWgQRP2yEB3ZOo8fvTn4ztmtnancXI+XziXYmMrgkVjYnpoxzpuxuTK1
bTRjeHfA4V7mArBho1NteJ+/yTxPfFV2Yv2TCF6vVXL/SbvIYlBwO5vAolyJ9vGS
WeFR36qjeBV3XsrrfKlfql2QLCsvn9sU/Wp0m0wE+QSxdvdZnHM3CmeGKIXSGjT9
7x+TRsh578PtcAAnOp0EgnzV6VxNHLcXQTaMcKiWif/wuziggAC36lpbIYDnwsGm
eTA8xZ2wQhhpV8NhX3s4oVVjmwZeTwjgM/0DLzDQXNLlZYNiBLbjLL3aDP7k5gco
epj4TE6Z42Vzby4vU0sAsY9+hxs7qO4Q8uSMrJ8DF06h30bd2olVdcCB8pE7IZIs
URX6ZBncGVpTLyfRAIMb/rmhIHixwCAMqqdK9YY16+7MvPDYgHe6a3oVgceouXPb
h3JdNUwQAr/MPy8psZDs2fdbF6AH0jSzwWp5bGkB7+KTG34vixEmYatcftlG/B0u
Vvwi8OGLqXx+tLBOCgQj0z7Wih+sBOY8fRpMx67LjEdS5+jrZ7tWIFbZRVI9epv0
SiJqKwDhl1a6Vd0enu7JxiezkMJooK2HocAtTBlME4kR6HkHngoxkCqPovj/mZd8
a4gTNWJlyA9+gXWCjuu8pquwiTKAZFn4SorA6FKaO920FSpakNBVjnPK7+qIqv6P
oNuNcUksQ5uhiSxxIrr0mkdUAhdGuKgeYGxS8dwgJuiDQN8Y6qrlhWbePp7q2wx5
Npfw3mBQiwhT2+3GohATAdrBycL1wLnpICHHHeKUNQXHYY9Cw5O4s1MdnN8dL4dO
daqvNucobgYjvGeyUZiZMp1KWMkSR0qAlz3/jBRFsvfciMYUIWBpZa5JzOnU39Ba
B0Eo/HMsVoIWcGCpVcR6wjyPQ7/pScfo5AYruXyDx2cvDsENGY5GnnITLxUPxadh
qXXfuVlMaCEj5yAmaZ3KMUmquLnke5b8bDBX6DCRvejFTiYG7FHInqvYtT4jG+2a
N6wcriTmq1gRpKcEwpwlgPuJL3DqYh4WAmL/3vVFzE/zKHhZinlYS9OG+RQIVBao
NgBLW45Lxv8ZdR6PbO5DPOkkD12ihFOCFZwsmxrGzy1/cahR5BGL44y4w5qA4B4y
ZCk+C5DIGP+lD89+7wCmbhOrq1N/3Rd52fIKI++RW3VBGgmUI1h22oOV4Uw6+TIG
YMp/c3vkHmm7sYEJ4zJJAFmTLgJqRxD8I6o2hQeSjkEeRwyEALg6g1VkC1moLibC
2nOpl5tiqg+wBDw58r0f940e+zvPpQwnWjFXkKrnH+DMB7zcB1uyxcxtf60lgK2E
JWi//9T4NKe1go58WWchQo8Xy3O7SEHAgaXvzQ1gesTpI15DjG4SeSkJ2Q5kmU/v
esC1f1lua59Ar87BfX0V1MH5aYvxdhBIWqcbptOoz+ITz4Z4gNzWpRMcFtaRm1YD
TZ49NFoLu8qlM+5oXvISRzL6j+HKhzmEPZ+cDx+7LFZBN/UquT3aLtDJDxepaZQV
PCPfype7iV665MDm283ONqC5sWcAibDMxmbEp3nHQ1BxWdmnIhKuQ685InX7gu94
a0QQXE8b/1WyHoSRTIGRmOWtD3OjahHgILaQxL1QKraVIMO5nKn+EK8cRd5ZNNcK
f2U28npkS9ag3wszuPjmCjD4NwM7y5g2hidKnVkbObKirXiITpQYXOd40IfIOLRZ
ZUp8oaHIqNzeHN2ge2fctJRZ0n3LeJ2bDZ5mPYuS8uZ28mTNf9mw+xL1VtzjFS2Z
WMC5uAVa87v1fKW5KX4aDVufAgYiYeDeNpxOlD7jR0Kin4ULRILJGrEpbuuQWLVQ
QfW503sI1eHGMaibZ1vf6m5nBov30FID7/MH5ogFrJwBiMBo4OzhzNHS671RsN1y
akMbQNQrPYo2jq8BaJmJw1xzE2wffo1gjdxwhITNp6YGnWdcUYe5eZHzz1l6ygGP
EedCKmnq7f3vV41agqwsbKmJuOoNmCcLU04vnn91qBZp3okFyejLzgCenOAnQKAd
qaJjcdY2VH/41ONiAJk8UeRn6Back67wgZajCt3UVWgm+6Sd0DOfaGFKpk9lwaD/
9WbQNA4CrQ0UP3/x+ZMo4YpTePDxQ+JaewA+tRqHXK5owcdoMcGXuVzQXeFhMQ7N
9fHUg13E6EznUUL7RWgFp3fBbga/nv0ZoEfcp6fo4DOJj61kn8A0WkFOmuZOJAmm
lsnLPsICr/r2HqNg/6l4hh+wCK5z/Y76JUnL/cKJXe4r7fgSLiKmhD1BzPgsDrTA
amMazNybrLyN182tRmNPqXZRYY+jyxklfc8BBYgING3XRB/HQrUoi5jRYx2cti8l
mMyQ/DSbtxTf4tkKEO5S21M4b3T++gfcm5phMRqzNzT0rKZYpb9Zo/Tbk20ybOFF
8JEtNiwPMfbpKAUveZnJSqQ3feHSZPOmWxr7R31tVVpeXEQbvC2apikLuCw9+ch2
CzJyZNiULVMR7RZyfvEa6gndCJVR5VR0QzkVIXWcQcFbL6yblGkBu7oZ43RYdI7c
/r0amL3JWJkcFVBp5Rir3OaRc4vcCZ/VMsfja/hWhhctDdbXn9snnEfiPq2qKrQg
tn/O0BtrajMIpIjPaCh1EqsLskg/NLU3MMtBdM8kGlQhURIpoF8URy9SQsD7oMPX
Mdg8D5gMOfGQsQX6eqJOkxminpWWGro6/CxvuGfvZqYEMm53AfMD5N+0qMgXy3v8
N1vSWBLBhIVJFC7yZaBY4oSGapnpaG4QtuvMIEeLf0R9ipuDNw0UOnslAJbdcWq5
0mY8pFQXlNjap2uULIWbDflokyC7s8ByTf9HqHvB8wKlyNZ5iZNcsCJ/KFAiyIPX
msC5tA4Kbg3qeqU3chD/RqM22rFMDNavUZmFtIKclhANyfu0DFaEFk+kp01tsVH2
1saiOHAxMu0F2uHl3rDz4W9C+MoLW1Met7F+PMWj0aKLymWm23/56ayyZmoHOtT2
DUeJQDzNEyr3IfZ5Nfx/aalKWAY+Qa2emvciyJQtQK3MX5hlzLOfd7+K/DBju0CX
vt9mvNn+6MrUsmtTJi0hhjTOGhnINvBarvGy8tNgf9YfrWSqYcGiahjhYK7E9YEj
zSy19uslHGxz5WCFy5vRCmm4Os6kSZ0rznvlDcHw7KUw2gQRGroFOxxlRVYcmlf7
p82+x5u7Zs5A8MXgxdIPbFnpNEqp62diI0Khr2ILvKBHGrjKH/YvHRQZFYM+0ld8
AlOIYqjlE8wW6I9Wi3nTdT0RbkfnwWyY4QlY99p91gBlLsp4kjkvo5JuAjRzFFBk
gxMgmqWfV8hKTzcoBfb3gtf2k30JP/p+vvrtBq4gl+TX1yi9HC3kSe7TwqMHTWR6
ijSOYOn70DRCjTjlnN4xHRUK+rhsFtCLV38UIh21pOGEyi5JJeJdh0OoxEH2WUQT
mz3ofg+FFIH7eVWcQTyrZ6bTCYCPbpXqmcTO/HkL0a95iV6ft80LbCLJzq17x9cP
KNZfJbzU113s4yEoCTUkIitiwoDTsh7EoBra6+vttC2HNqedCcsNFae0qhWw88qo
XbZgZXqlhvclrgeEsEQOThveXkR6sH4N32h3Tj2I81h0gu3bTa9dPyFC8y7cXzUu
eUcP1geW2XrwJ9kXod0dMYCRjnv8XJG2+3LlwMMYHdcn0dlU3K531ojbDhKugzy1
CpN0k+GD/GkoDJp5RTYbvdp1NL5SjjgyUre5z336UGkG1d3JS5OKSBX5VbLQFxRv
rhbkhKvehJ6mPp6JsF9Ue79i8U84v5LUyzFRqcqOXVAkvx40uPwT9wUZua9awxo3
ij1Zn2kemfTEKaCh+VNN5asrBVLSaW+jia7fj5H9UuNVWhknWhh1cXJeMrz/Mc6g
TEyLTyZn6LZetBLyCTC+La5Ei9CcFul8CkBRVLZ4xsO0Sw5v/0YVZZrLLZRLNT3+
sxsX40oRIM7dnwDgNMpYbFXKa0QEjdCBlEFK1Xe0JtoGgiTUCWzKE2tjtwswohIn
nPRVQIKcwh3O5zU9heVZh/cwHbkh7BdbBKkhLeaUjZHX28BhonSaHktZxi6sxTkT
AnAaBdDn52/U/Ev76Tg1uAqx3oMSBpDfUNs6Z/Uu25hpiBi4vaxFOl3TVYILSoj7
tuMD2UDFO9Vs4qTrTHyXY3wdIXP0lHLEQyki65OIe6Q9xFA7cO6J4TO+ju+CfyVK
1LPrDAoXrlkvhVsiroU3qiOfihyvLjqSee5aPlYJjXSbXpUuDpYz2jxxKcR+AwOz
RQSaBn/OeZhsyrqN2jgPHJVfce3BV7rtfwXQ5rH3ns5vjjEv1O2gFMM68y7k1880
bxPKGrcGJCaLqDIddBO0qpS/3mrEMVwVHd3l3JV8ysafCjF57Qc6CrqKPMIEfk0l
MOXrhsQLxu5X3BolSKLke/AdI3XJ0YBD7Cf449CoFdqdJ61LRAdSOfE4FcWU1H+b
R86PYnFqHRAVgnjjyzwc1rs5aJHR5ZvnrIlwyYPVUujXoBnhR+EEKpnrePsxEWkt
Dh7e0CkRq4hXjzpFlsVa6ow94mesQ1vtzRH8lmrXgxv5zOoS5cRyair9gtyAie5V
ImqvRxWaXW4ERC50ClJ5ql5U4GpyOJ3Eq/iPvTvkxpypfYutlX/Ps5jji6JbtlbR
QO/Q7el57ccRpyuzd01dinrmxS8+SVMcqkJTffFpDKDGnZIaUKCOJVQMED/sophK
J7cGPHOiJv4f/52F1iThMDnUPyZ7tEci5KUBlBFmyfAXa8i8e4wWpHQ2RrpWZXzl
ov+04CVj0WgjlzVSjAvEO0VCzHSnXD6OlLNrAw1M1AymZ3v0yXFUISTvchCm3BsJ
dc3cEh99D2CBvXOnAR1xUCUrLfmDZN7ztfyt82kpfU20h0DNiGuqWJBC6x3BzyyA
tMxlfMkTOXQ3KXqmhmtlGIQHeBtND1m1Q04gHMA74ixysWsHyubL2pizGvCJ1yTp
XucfiGK0g3DrhUlSciVE6yV23yc/AdBprEFQbq0xBLYzN7UtprKCG3mFBgP1pWTB
FEOvJRba8XvzKNZ1h5HPYHsQY6pUChybkK9g0FpKsSZn3P6Erj/ADnQzna78/Wjb
/3wz+G9+DqqnxmuXAWrEJ+xbwSlqz2PL+8U43jrUOM/XQZfqpoT1bJxci/BL34+6
ixAK8HGctdDWWEoUG5O106fp7rVxLFtidzxpYWfdVcLiUZCSWExEVHgZ2fEytbdl
YB9CsjXGBXtSunpGJzKVbS8XU6FHxdVGDFVMqJBNqfMH0LWFl+krceNy1Bzn9vib
3Furf+0JiDefvrC78YmwGn4ocCtmvW4a+HNZoOdYmKrqJNyxSCAytVFZd10OA0yA
9XyJZgZiid1jyuWnULaK7ABJv2PHpTrkxYhedqCgIHEzFqsgPL96zE3Vhh7T/+ph
7JsQMN/lUczZSMhe+wifXljqnLwhhbW/Ng7R5NIrznNyUWv4pLode6APurbbmzbA
5RjJFaFX92MYLXugI2mxpAtsGPbOOybko5EQ6CE1Z9s3AOLUohO9WJk9BiocQ8eH
bn3jQc9EsRjKO+JwbNgbgAFrxsnsy10Szz5Ak5+dt07ILxshdTkoLUg4twTlYJpT
Tfu/Ic7ICRXnQKWwM/IcaCr9hw/IEAwSYF80bB9jxGBBeB/aP9pmGq3kwLDgAJat
hKH7RRC3gDYXPot5QH48opCgYy9cx6/ESynibwb8z5tH8E9VpX2/Afq1xmcZ+ija
AsEkmgehCwVhWJWjoLTDmUDTL+wQSTZkVgQg+48CVTmI55tY2yYLNtKzmwyrkz8M
587rQlENPorJmNbQAYc+SGWSxEr6nNXWEuKduPuhg9ezDhQOYSkRlJIVuUbQCfAe
ZqlNTIw6dYEE4W/X9LuedDZRMWvYjDl2nkmWS0PwcPrjXQB8koimJmC9HJNc22/d
P4g2KMoxSC3zau8NE+dpSseQR+utM+4j6eYkQkfPwCIXUftwk34eKbwli8fhUwRx
f7QDbgXgPVG0ZVLzy6He/kR5h5P6eijOxVsBn7v2aZsER+3OnU8nOvW4JOAYFgni
4iJywMm3Z9nMfveX1FNE03RBV73tnfcMPAvzH8LMlcDi78bhwbjI9niCQcGInDwW
Vv5z8I/u0K6nhA5DNyfD4e5Zajz8JDwFTekLJNu8eSsm5S3z93BbzJPSwij3tRhs
vcDuR2WsZDO2VhNseT1zjkr1vLpikRnwJU1utmAw1YNNP4NMFUTXDnD0TWaQN0/H
IJnWAQkj5hziVxWz2PkLOU62DfX+q7l1rHBbmCMN1yINFw4Xkp3QkQkFztcD2wve
f9PRlpHGOZs8lRi2tz7C1rIc6dEief6oWMO0dNiyzHQrgF29lJ3xdgvA44c6hEaX
ppV59Vz9rn8GV+9yt0dMm/nh6/cJnyMDdLuRS4ZsUj692ZdX24QbRXiApgsHVNWr
GcG0prXGIPmX/D1SVP0AaNvA5Lh2VuIEc4zxm9OU5DeG5XbcYOsxpX//WWu00K1G
3ftBRvb315DlOTRkWyFB5/JmS3+cN2y69n5zFpAC9tqQ3srBMKOsxuvERrPTrnJC
ZmHeqZPsBrpbtw5SwYBNe3Mf2Y+QAgjIDmpDZJGkHdw5o/IlPndRpOc/LwJvqK6E
yz5MpJaCoqBtgtlaZWacnOuUraAljG8KN6lzgrA57yXmAo3hSHD325LbUAWiDMw8
cubOO5A+UbiVcVo6VtCDjUad1MuysJx54Ktc3cgG8C3CwOPtQASDB6bVEiZAkxn6
1MBaTFl6FbhEEeBTAkwJ3ZDVBaSiP/M5s5vtQklgBQcdwyw5s8cEs47iXS86Q1CH
+Tt7aWs/8tfvIJgQn8L2JPvYLOpXVw+aey2SuFd/+e+lIe8mOHr637RSyJ2eJ1hd
ZEjO+4rVjAh5+AmzBCctSpgU4Lg/x9fYrFowA14FbFbJqf5Z73c3s2ld5SyM19sY
HiLG57QOQDIR5dAiE6YfU9T8T+eLptjdTJgCFy5GHFPrY1JgsPFzWcjdHoizcCfO
3lfMsNZqWVZOQj+pSKimIwfsRTyweR1vPahmFQbw6eUaYrdg47nhAXIhZv5vvSmA
gs1IIp1xhEbTZepuoKM1e7yxw+OB0pzATiOtKNK1OkB7fec4j1/4bQLgLUbVqPO5
glzbctZTl2T9tNb/gl4TP5x1SQf/qBke8HrgiQxIH87peg4zrBkjoukbcL+JtZDz
gbyHvuZD/SKQO8jgwgiXgoHgXt1AJ7UReljsEmOq7ippGniqqqNT5fI5a386QaRm
O0YHggOPxLuU2Bv9QKej+CCdHvbpV/lNQUipY9QD8hEJ98Y0mCxMSCG78coehxje
GFLt5C0q51DkTzQSkw7PTd+cWxbZoWMXaQAlqmQ6JmS/EUFOUGrHbod9elCV5HsY
k3pwc8GKun7rUQM9j887nO98ECt1h8vnmxvd1UeGHCzaZyZe/a7lRRUp67r5e81R
PAQ7Aiid7YIfLl5zfHhdH0xC57jt935vpGmXB9OSUg5roxHQ2Dy5CF2O1celndTm
9BVFTP8cWwOMv8MpPPUe+laUAIz85PvswXrsjpt/E/sgiTnxChaLs0W8Z+RW0aD1
0xPInY5NJEqUKjOEpRCOBDyhbMnOi63ECugvfIAfe8/TgAl7xL6H09Cz7dcEU+He
s1VW7rCxJQhOaT5KYz+YYJzJjIzwwagsY7Hz7I264i6PT750OC9UJtD+Uz/9O/1D
Q45KQAp5vgu6KlGLsZSD24CCNn/0jlmjODmqnIJWswCY0h/cleWhn4tSpXabDqin
kmZibtFvVAE/zTB/pB0uNFCfzqAuX5texVnZdhU+tt/SNXMfsNORvPlFgvy6N5rZ
96wuvLnfw1H9iC2R6r2B9CU6LYgfRpH6oI2FquVXcYezU3b0KCJdkHcPbO0UQP0h
9FD9H1xCaxVb9Mjb6XdaXZNJoGN3vAxPU65O1AH+aROKBOM1SZWHHi5mTVMDs4FJ
NdV2jkOZzze+XVyqYcvw7A1kaVRgO7/G/BeX7CTt9kStpno4sq4tbkda0n12TjrT
FB+XDMGs0L1thX6Y5JiQijUqttIw9DAh2uE8HCGctAXifOqSVJdgXJwKzgqjKQoH
hOUTRuksM1g9Iy8QQowiPMJQ80GByeLYfX7soYVKJ7B9pWC6Hndhtj8jjxxS/HKs
3x+VCZ1UgeCEMBZ7TYeOYSFfYnxl3iBEX0xZ7C3Oi7Wju7qPDfQOAqJ9fwiftZ0x
jhjbByghC+XjtZW3Q6PsxF4+rJkIQEI9iwaR8cGJUSVTpfJz4mefBMbQiy2qFuYj
xzeSJuCk95iTnm1t2b1G8nmw/MZfTp2+4AptoZzLMPe3jsZ5XX3gkzm6c1ofzETn
SyBVc0ZNZ+ROgXn13r72hUiPSrFgCfdyefbFmPMrzZQxnD//u7Vtj2GHm1ws76Yw
reZ5/eFTAEXJd23tmjjKzyWD3lRNZLDuZzWfMIfaw5ShOPb8o6+as5553JUE6yw2
hBeG03KqoCfc2uxRdlHYMvpPFGEEfmENt3sq86WnpIHaQcVNhH9zhps69pQrMP9j
3mzJqTHkHuFlldhSmEHNOt1fZTQKTSaPfMMzPfC0H0d6czeYmxY1DKmm/qpnfDb/
D2FPC3mEGFw2I0HbvJ1XeSt1/ry1YopUJCiZIUGBsDM7h/JM3J31G8S99/sHc25A
3SD4/x3MkRA0H/ESKoOIMArW8AvTWFpDTrxTy7nEaOkrwJpf5pUfDv2RetI+0IYm
dewqydiustMY1iW6ZHw3zkYr0Dd+vfPdDvQcTT2OEjO87OF4zhwnwFaZOD5QPoCm
MEDaNtUX/kCLbyX7ZNKd3x35MQkHn21irKU+K15e6tsK9hoXejJ5ccinq282Byfy
bKEn0EelfnW+chXW7N5fOkEoMsCpgQSsghs838QJE3uIPUhJWlylQo1sQxohLdTe
wKjdNksThjt22DqC0DwJEyvTw4mOuspw27BqkiwYlKftijI+LdC+N5z1Iwem7Lff
cTzEQIPtWt3hpKHIeLOoNH3b3B8ajrZYyq9GXGDtFr+6FU0TdNc6QygK6CJ1NWVN
8KkpPtVaURhSfsSoUY2Dm/8aYOOwf7tXgfcnFqKpZvAqlSOArpF6yV6Y/iaBtKBp
LiEJfrkMt7zlmPiP7X7RjNjJ5vQlj5WdLSkARIj22X/OIJP3lBypbEU9yH3/0faA
/zOPm21DMBGyNoZRCdVNC/sm7BP39eD1QrE1bD4686ezWJsTmJTQ/4H0wcv5U65o
eTant9DQFRbkYY8rvh3YxUj4Wb4YbrMG+U+lWi6ki4cAoGVsruSaLSrx2VW5rxlB
2X2+aAZO5kiV87o4vgWBSnnwYXQCWYYQuFso9WEt+fKihRADyfpfXzdUPiGrif01
GS4BUwjPOh7u/0v+ITT1IGKotDxwQ+ic0Y1Kib13kGALX5th5Gu3ZmEFL5GtVoAK
odtPGdhNx6VlkEFid96zZqDAjbGDgN7NvBUNMzQYrcU1+lKgmDtZH6Jt5QdyxFyO
i2x9rsqfO3WkypO8oM527MiXbVPGXWZJZ55kEhuidmXnhMHP25YoWZk8vc9I/MdR
nA2zkhzEg9WDYib7Ei9EdFs/5YxXe46IC6xG07XcBTMPTSnulRC6ANZ2/B0iR1HF
c44v9t6gOMkW09jZjltLrrLWKiwzYC5TJtDxCuuaKSdV902vffni6VpEP2CesncE
opLXLSY03dCZdchCftWGyCwpePekpvw9XMljavRDl1TdmqrvBvJf2h8mAIdJ4XBF
J8qQxDJ3dnIR6aDpHGS1oFLPSp1sKQLNp1S/cJr4SBdiOnolDy6gus2n+5WfZvdL
YZ+S9HBlwkVI20f3tgT2+PqEcZAKpEVcEFwLeVoUlXihCErTlmT0Ei2WxIU422EH
DPSWbfxiiMllptqhEB4tj8683bjNhZp4ygFRc6DlFxKXY1LSmKsM9JIKfFOcroyg
VAphcKGiFbe+Pfyq0D3fakPyT/EH9jrVr4QlHBZgQ8yj4X6s8gniVEtoNSWQCXLs
yO+matgdpXpLuGniveZW2v41LoefsW1hX5QgIuii+YYcxQA+cfSRWTSTaIevK0dn
WMDnAPTRYqNAEpYKtsu4GifKkNcIA4l6h1cRTM7liYfO7zeDPFfe0Ki8+BqdSL9t
0ya5oXjLADgiku8hI+ZcQpmvQH7hrQ+xTUk6OOSxwWIDdlP6GIollrmtS5THErCR
SCL5VF4jSUJBuL1NSKyxFa4+DkKj3ZOY2EJp6jIq7LpVeq1CoJZfcv62kaw/TUNm
/RKgN3i9dLGz7DiimilUolaAz7rTIcLnpJPD7Du/9hlLC6651qh3YjUoh5f7110K
3VvajLs0WNpyf3SeaD9CEj+J0EeIijSgGkJNb0FyEIRF7a64CjdRvtcb2JCQ9U5q
ls32X/OhTQOSA+JyvmeTnYDLYi2Ogfc2ETJ65/PFLAoIc7EQ8/R93HNXW3UtEmEg
d7UfYRJXV0cSy6fExBMuCw5AUaV1N4+TwqkrNyYfxsBGzZikGg6vqddU1xEms9rC
arE0MjtOA42so8jg0nqRG+qjKFBDHGhUVkhgiAK/o6F0SHFYqkHy/dqd/liCph3K
7//fU6xZZNYh2Bzg0scWfp7CQzmU3eV/3zrYjzPmcI2YbQVjP5Zea9U5eOPCCxny
8QLn2qm89N8o5uHconIamks5nSndcnX7shynr95EN8RLBDpRsPuaiPEgTrhbbjv/
la0XcFgINYRi4vqcUGjYPUToYDEGz5e5K6ClX4CW+JBU77TZ6t5KWXBXit8MqI+x
x5xmFPHEoZgvfcqLmfOELvs/HNQY/vX35JwZbeG7lKgwOl1dkN40kwHaZtlLEjFS
YpMmZZk0ktjwoE9FLqSBq9+ghD5n+J7ra6QLiszwLgVjDIF8a4X/J2KMDabk088I
7qW24ExY1HwayG5aXDbINj51e+W2MyyD3TJiXW+yDS8+fIi1leZMc9VynOvpPNk/
ERadgz0v7CIMvgUVsB9eSlxO6DdvZFmFTxknOsNhdAQqkcHd4Mhp6rxBU5QwV0fh
MCxrCX18hlncqMYIAe0sFzrh4cUYO2Iv7REUkK5VpFGVVqVXMckBgH8susXyJeHB
WHrliurPcHqJGE3dC8Kn+mrtQiIMxHXJaGIqLUC7l9loniYCArYt4FhtAHZSdKqT
Et4T+iIBjk0MzwZ3bfyqUJjXQ9L2G1mTAa4qm0maiU0oi7mkg3dhQfZs5FY2c7HT
GhmgcnAoBeJFBumu0W2wLFbz84x8BioN6ra99txccHDv/a8kGDC4gEl4P2hMHlqI
SWEXecP/nAKVbTdapV0KM33QizdII3abv6zJrUmjEHj3Ugui+pz5q+zok1JNgmku
zw7jD8Lsb9IL8BL2xMVjJD+lxFkCj0nkG/gqzi5nllPlpzgoJyzW3UX1swwlGH8t
7PAbI1kkkI7FuHOYrsiMzIPefR32jHDmqnxXxzt8f5aZu1fPNa9ijlzymiZV2dgT
Fxxachfr3rr3YmmsKiQ2Mzoop9z5ziFAtN/O08++Lg/VQySGwZ2WCDmL4YPZUBa5
0TLz5dHFv/hiEA+R7hNwnFC1yqFQl7FPXpTaFz+pGQ90hGFfRy/OMkfbWYk5DaUJ
IbpCPd0cIKFlP0a93RdIrkwI2UJydNf7GxxOKTU8RUcpWT3odiH9xsCn4yH8q7i7
itFyr4p6N8hHX1DIs/e9apKUfk8kAuxeLnpf61JwJJXMZZsftAitAoZZ2PwJ6Cux
KRi6AvN88NYJtPNWJQUWrLDljMevV000RRw6oexUJDmcVYFlEy1dLKwR/7XhaFIh
GW/ijqhKVSUjbT5Px7pf8ej+fe5c4V+A1s23XxLVpp1W0K6HJljsGLpESdFwUgNV
YJyBHd/p3O7rvrkJepznMWsBGRWe/Q6pXuVtGLIB38xWoJc0jeHCjW5bMSjShEpb
ON0kk/tBi+pu7olTefmHbPh4J9HKpft7RXACBgyPbhN8qjPfM1GeHUqmKneocCrX
x57TCVPC9zzHEkMUBkxLnt+FBqcw3BVTv9YWZJmuuX4vx3oq7uNTIzJLgEAcCRLo
ukv6Ydk8iEQa3UqBfvTz3qGdv9jeWi3dugL2AflXj+jLTHANzzDBCzG75hU384nR
vmk6zDDtoXWNRuE335ewdj2/UMkjyI7JQGfS0NsbLH1XcRys77462NMb5nOyiuZs
e6qbYRVJK+JVh6otfE7IVQ0Yq5mrqWhhpzVwdqYn4HUMn1u7rOWz9rkUk5mdwi2k
zLYbJNmg6Pk5k3/hDhhmpoynCYgEAM/QQv1UO+UsNdPoVM1WHXguFVCzKrqyfAVL
qlNxK5Ym/IY7cD8/H631XCTjol1aWSVbFLFOUd+DqvTKXBgWGZTw5JtNSSQWxO/6
1mN8n8/TXEUAJzlXVaORwNsap7/KGZYzRPjqC+mfUowmpZIDGxTS7356IaaC8wd8
y0oD6b75TXmQxzSgbmE8t555Wtqogrk1zDM4tbMlfWPhEfA/zIlwJ4+D7jrRIF3n
dPoAtiBoaQLjpKEVtTMh/aOZIwZgnSQH94tsiBwrH7FvTUL9kkX5cx6OYRjZfFyw
FuNya5HN8OZRzAzHGsZYvjGqQ7q0sB6DoAY1olrYe6b3dE1/Q0s1gegj45XDryqv
ZVXmCFi0H2kjHPjaCYczHZR3bGxXiBWXFQTmKMSJOOxDrft46Sht57HP5U+8VNjT
nkVw00+G/+nYMjtljYdv/EQL85t0WUwza1ZcC63SCRAPAiyVBheThacetd+5BhWu
S8GIBwV/cPXWOw/yMhmN0TMg5O6dWY6qFcfTkeGyDDeRNivUkNLOt0B5iJt5lTJq
yVuSU76sbyqQ66kO44HKNdqtkoW0fBtlK2EeA1OfH6uVo7wwDZgsh0TbFTEbW3lm
LR9UOC6c5ylKbLVYgKXzJrGVWkrMA+G+V9eAsoXdjdDiic056Odn9s00JXz7eOm0
QgiefTaKUjP06ir39A4o9+/7IF/rOZhup1IpeG38GFbBjVnuHHDAthAjxvZZJScM
c+qZVqkWavxFAfNN7VdZ48Yzya3v2CccPxAJOopkbztvHQuYKTlL1o+b5s0IIyRG
kUxLKOHsfz4zB2bHMlCILYjhl1TkT6PkStGBaJA0f7qEqLA64AORtKqk+rdiStpT
PqiJx4PsW6GzxfVGcZMdJCAuZw+yWJs0MyqFGcVVcUpNtw8+/Th2c6B69jllLoTh
cWnvOjzOw8sNjA7f0D+PjV6NKb+1jy/nSVwI/pEI66sC1sE5DZ6CR/M6e05yZJwC
5ImfNQYB5xXXUpvOGkNaI5Z31xyxNnp9CcBtYVvFzPySJw0RmxWIcgpagg1aPLAo
a54JOLOKR38f77yTXSp68T8bl7kJBh1IX6UtqAJi4rKQ+zAQx2FojulIM285vdjD
t7YbV1E/rGxihT7LeOyeos+4kuZLg40N9qwOuvg6oBOylf7XzpUWE8aNOz8xf8Zv
YL8NU1irz6/TptSEoFY/8O6EE4ktbzOXlHMypFL75L2zhOz5tHSGoPd3lLp2sSDW
vWSFEiQ0PNOkOTfnLogXT+F6qNEQZ3owZ87YCm0H1uWsIYzKy1SDalY6Yb2OJzko
vc2gPCW1R34GLiNeK6ukvy8lx7WRmLzH42BKmqJGocnxVMTMwyaXx739S1dDNVen
vilHNy9T8b+s82TXLQAQWKuosETlk0cXsK/SYI6pPEWoeNj7/VFGd6Y3AuOiGwef
jz6HtrpepzB2+Z0i2l97d1CgsBGDSWi/G8PqxPMwf8/8ylJ/PSwCurxgEQFhyWWf
REIsS9foM76v54n4kVkYo2Om/W5T9dbE0aaogfmh4kCpOKZILXN6ME1pE5YC6s7Z
GIPnyd2H8zRgARlHZELE77H2jk4sumqqUVIp2SFTEqO1rwKZAkmoKwND0Hwi1gIs
xROwRt9HyA/GGXzE9/P8t4DJhJd7YM9pbQIVsXFFABPxTU0M6s6dk2ujmbO6u5m2
b2BJc2DEkVJx8QswjVtE1lh41tvs39lHYXgr5aHACSAiggwgrmH6G9H+YNr4cTHZ
iFnCvcIPA9Opvn1p3s0J2A7kxrY0VJgPnWIJatomDTmDXDgRAVoRupX0VaZzpqVr
LaRmwho8bZ+6+p6F650aUmv8ibxSnG3JDUVJsRU5zkHJ9WtTMC4cDdNltsW7YMNz
bn8j5wMJAUUUiGyOHa7+ZFFvkzQOJoxavRIr7njUlzHX/75Rd4hm8Xijneyz6jYi
c96aIw+cfqSH5QLZ0rqToqqORnZmZPpC4o3pwC59H8viZPVRLYnVoSiZ8Q71WNLX
oezcQ8pzC4kVzuZTvgVIXlOKgE3Cjpd2R/p4lvizJswEfSEQbiMQXRSHJfiPnAHG
pXUHHtzjCtGFgDlaHf3W9tVe5yRszc1Q2JeSNTD5u9xU53LyTFqVuhTHetEFMOGT
17ot8lSBXL2jMTsjmyy3pwZYA+0PkR0sLAlMC6GgMDQkR6gnGsOYAmPfU9mIG2bX
B5sLk94x8qRfW+vN4MJY5avJbu2m1i2JUp76NJJCx8ikjdPM2AdMqJ1tOe38basf
xBRHwJvzJx+97OSBdYsP7xymeq6YUpI2HGxuRaiE97vJHjNa1kKYDu3UikFev+PF
OP7KMycCgaja0QRF5GLtpjKC4I0kt2Hdvvd1GX5mYfozI7Ojo3maLLZWmQV9VTgR
5AVdeTFLuRAJPdNV/UT/5dMWvKLNDVib3+RWUykDNsjZBM3Jc9vQw0pZqqvSbh8M
BY894diEMuezNu19pOtMfE3Eoq1hW4qDpNTmJyxv3tUrM3IY+MPT+G/qmVBwFo+S
cxcpeB5iGa5rRXEsqE2jsGqLYXEE6MjftwNaPLHTuaIEo4qT2sW3Bc/l8Dp7KYBN
5SDxM+Aoea1kofXJnyXAinh3ncupffu+ELeecq1dXjfUd2+V1uC2TCbgjoOcVuhX
bZceRz5HjsAe/pSOuOw++ufRxi/E294pxP+ktRfmG0nRZoSsPYux34PePB+szMSB
ikDtGhlmZgEF+rspTt+/L7LiU3wzaedwrTYGm5Ogps0SrU6jimNnkvzvbxlZ/WXC
+bWRnDl1wGtjQ2mh7SFAkvEr/zldVFhF2QMK+QRR2abzVfUExgGoqlPvkmOrKS7Q
5yvj6gOGWbX8n/dgakoxg/AV1CY+otVS7CxY7z5B0lIC7bEcb1pqVsZUyGhLHIBF
Hp8bv2VDevypvzD+pP/g5Mx4L3uTy3qpe+sv5s3wQyD33h+pqKf1+3bzYiRXjORZ
DVFWytSFQN6MPR76OnLMjVV9NBDgPmNuIoNlcIYINGz12oH8crEBbFIOPHit41O5
VNVtpQJC/ZU6/bW5fJzeYeSsip7IlIPR9UCg506P0LpkYXOYGieV+vnMJ9zgT7gt
v8Zq02wdlMdJV2IG0lFuQk2LEo0t/Q29K3ElU2CKIBdGXsErZcuE9NMaW825QQM7
KsU/+upVg8OpGhBSoxK7+C0uFb+H+xPd24UcXhRi6Y1BhnCCFPh62pciFr9+UZFr
EyD80olkXQlxRbYxKeZuzDSjx1NXDObdHtkYBEPRFxzUvgUPNosYOa6/0xrt++lg
BW9hsP6gkRnRhRa4aKtivaJl6TFZl5Gre4FmleJ4i29Ck7sVeuApa1aMUr9wXmLM
t8WUC7HRITSe2LSthWDDEGYSM2faY0TVYlvk2sU/yJEH45cFrjfDL5tHPgaj2N1O
cPrGkE1iTEWnSaj9ZBQLjkmjxUNKTbH70FX77uYtmma1u/HbPEdYyECgmTXbjmhB
orSgBifrONobLZZxcHSf0JL9uGDsv5/J1zywmoSyT92m+vD+tnFHdKctBFO/rmqw
wfk0ibxyzd3Qx4moKDD7Sa4TFzeoTw7P9WNFCkp7JhST3/HO2ZWZOn3n03GUl9QA
zJkMw1iAoAxKcDKCTl2uht8qzfgo+9PLygYralX2v7clzp7ch9Sql/qgaW9KHwES
MqLvbrwkJbzprYEHNpSOyXHuMJM8btLXK4Oyv2nkrB0GUmumDFofKCA/QTSpYfIp
Ti0WbgOHjvrT2XYx/LoWgoySHlAxxt3qBe69iQDgMUvY4TxgbH/Aw5UlBUisYX16
SSIXmqDjl8rcdO7sYGH/tQlK0AUJa6m7PcjpNPQTlzMYxzb6/T/ZuuTmJXcUKJ2G
snFv3wNkmoarenGFofar59zkljMbrHtzgomwidNiuK0/v6UYjtwdTUOp5uTuqV5P
4I90oqWVdTTXM39/WN9L5yvY2hVm0GTsNKbiYTrDLcUQdBi0nsmSDNsMcDbeepMQ
r8WDJLS72IlXu6Gb+qX4tb6IbXDOYc4DnldvcPuz4LFpDKCYP/VoUazpcSsatmp3
aZveWaxRxCqgheP+af1vNPrLofozBkVIkqp66K9UP1j4xU5MRigsieAFQ0oAnlfA
MuAyC5GYlEnSBcZEAATixDaiptEHNrZvRNI3wmlZGoj7p6HJF8K6snNi5gxr0raG
UPqKo1mgTziWW6w4d+Cwd1Hl9HBP38e010wPo+2VjerX5vuPY4gPOY+Ili13/2J0
zesrizjXFz/ilOnvp52HMcx6Nt5lndqZVDE7VqmNUfJZj79zYutSCDg9wBv1VIgP
J1XD2zTrXvQ4mfDnG1ioAKw0hKEpK2Qjkq6iSGER+az9FQZA0suuPuyieGzmChNx
169P5cKswrEvWGhga391+ydgRpACTikb4xMb6HV9WfLklCqbMR+dVtElSejc+qyU
icBIn0/X6kmo0WfSouYXV+i+eRtymFTBUrYiEl2MzBZcFRTSVHnmpnDIM9Yyf6MI
40brzSodORj82v/5xkab0F+xdOeQwcH99M/sE6z+WhECc2wkQiEObhDBrnKqQna5
FR3Xtom5n3WBCS3pwRzxWxT70ygbTAltoHenU8s17HFQV9JQU97J47s92xfynNEE
180po9AOIzNpzL0du+xMmyo+H5pNz5WIorL9AKqqdalaJneSlfmEP4b8DQlEoqH5
yrlAXxnb5VawUzdibcP0z/U5H7sC/AzZ0jwv3aVLNqw7gMBgEsSYlrG7dEnhkAYk
M3l3NQrQiJIosbR9d2JftRWWwKEJt+ynsAweQI426Dch8w2OEkcFDGjtgtZhk5b/
PnX0tHHO/u1EfSXbIYArTJ8/YvygNjOCPXvzDnCYS66wzP7eEhyuYfWbL+Zr+QfT
JbPcjf1NJzBc1/KgKVojn4HWjE7Ks9KuA7p/9EH4VKVNppV6HDn/jj8HHaJ+Qv9y
lumUqWOxPip7/Rj6/ur6b7rWxP4wBg8rA4kKdOfFKtWX8HygK9L4cCpY8p/t2erX
qB3MJ2gpGHI69aXwINk7PrVTmeSXyFErUU+i+DO6R5SDDLQImX/L72Dl8CYCA/fl
lMUDEeNN5qVe02mF8NhN3u8C4qk2VRLpUGojunEMg6+knIeT3QGhAvxwKWypLpG6
Vklm4nFeW0FG43YCwtOvzXN/oY5A5/iX2Qxmy7eQt+o8CsDIm6eZbacCeZ6TEU5I
3Kn2D+HlG6ts3y89M+KecLK5YgifCx3BjjQIUE1kGsOrAh4juiN65bY6ZJYCfx9H
mle7BLfxtHiRWb6C34eKXrst9R5/KOCt7IMqThMb5mt18AiaW0NjmVS/gmG8i7+3
GdKV6KRzScHdZsLWluqUlCEXV5URnP/MszW8p4BCcfF6QxrbnoG1jy3P2f+/664b
K0B439aKnaG1nnSisZM4SQLYkkxblpugOXcegK6jj/hhk++zvvjqBGoGeF1jUO0I
Su53/o5zJHqRzqTaLvAgXzkdkUqDDSiXcwm/BbZWDFOMccEzYuOQD/DQdAWqSLdJ
Bc/zHyXlHA1Z7doSTTyKh+wSJP0HFrwot4fAC3phs8Z2gaKf2mG1rtztlZZ4a+rI
1EKQoTK/IZagQLKxD3Myos3IA4aS1EXBfjTiQdaxoCnmYVhxm0nRAYqHMFn9FqH2
Zc7Gs2MBBip3b0eB+OSyzC68gQBDXHxrGF7KnoClGWUJz3rG7aMxZmtyd9MqXG1i
UHMJGCcNG6bB/n1wejucMQLA5eOnYrZpEjXw3S+yxc27exyL8aOBP26Fnhkp+XyY
MiJb5HRpGhOy0mhVpHDse6ibPGaa55EWnYxadIjVa6BEHV33P9SnlNJZqmZD9xcs
cW1SEoDqXyPEkSEU9sx7unHpvhFPIBsh40tZqspXoN9Jyd1CUjtPx/9vPKuHl+36
Fc/peUpxODZ/N2dIbCMKfEODko967FMDWJq814X2DUbtkGv5d8W3JaE3UCNaPSs+
KcnE+R8wucv3/epmKcPFlXxB0E3wmFClQZ/mCxMyN3JJFW6QqRGnDnl9X7ysWhvk
4Olch47CMYZZW1Yl9QmKa3c5Z3rlaSFzCHAvtYT5bB7JJtKi/92kscFBwyX6ffu2
JK2iv83dOPjgvWjMTdY869cq2q4bdabm4PX/ablMfgZMys96kVRv14ZGBph9vXxx
eg2bMEhFayc7ASx+JKI2TSfHPb1TcLWJZRiSXzvPp/og4u1qCGsdCECwI0A4QoFz
9+bmz/YiI90Qz+6n4c6Gy+jrXeiHK2NO1VmFNkkgKkdSrRZZ2s96B+LwwuEy95E1
VLPAetCNXbFijxYvWQA7XzlgUxpKnplxx3EJB7cknA8mhyWF+ovaaxmSLNXPbe0r
PsneRevGb5qo3d3p+uncUClSbOmX7Uh68yZ81L1V+HRhSHR+nsVXUE/J/2LhzJNt
AyRtIrhp2fKpyUXEq70+fs7XBl84a9LB0+Ptxfw2jae6oldYJlUo/u8im991vXkn
1a2LeDQ2XCErwfAJZ/bugImyRSOW0m4g2y7b9IWss2mpq7b/19ObTMJBw3o/aiNz
FZApJ0kYykVjXxv7+Kj0Wtkf1sdvXCCjd1qywM5P+zSTP955FvSaAGVQu/TRhmPx
hL+sSDDNP+lmY22YJ8MzqHn5Crc8E6rHzc527e3nLOVmzARg0uLGCJK1V1WaWoT5
7XD0ebplWXCe/9izcmgZfQ1MzLDUYzIkfoVQHaWn3cODwsZ5biukQgEMagpiUxIq
OISIEOKMqoqw/Rwz5gn8CD+pR0zQy4+3M6ziyMIi9sKyzF3uZ8NeD8BbhjdPPoYc
rn21WdS12D/2FDrBDnEoFnnb8nlG/C9nzFCc5nN0BH8e7fqCLnVJNnI41RAskINE
m98qRLfE+CvK2ALFJPunbC+KBFP1m8hWFgwHUvTXptgEcwYi//BYPSo3+EdJYNCA
k5u/fAuTnSRKBDX1Yah//lt6wzO4lr1TbCEl5uS13nfs864jnrtXaom4etSPO1bE
/Ef9zvWg6QXL+M0hSpVXr46q9JLPBf7sCG+BArFs8MSP8K/PI175/Rq/HpQ/0ODv
45AAXajWcStHc3gXOFkpYizk4HoceHAYX9uHrHQjJBlodpXKSmF7Bs6kc0gNhVYN
jiOOtuyb2Z0uK1eRkzohlU5wFpeRydbxyHEZUlwBhzUqxDbPpTvTrTds2mlRwZ4P
OwufzSetq29mmW60bnjzqBC8yMAWVPj/xM9Bvi9juUwWrNu1vj+iWgnb+Almq+Mf
N37/QQyCe+op12w6eiB45cUFkksD4CJOK0/rUI1B8kO/thomllmWWSMrj2Q29ym8
yrscbdD8f0C0x8xyov1S521N8O0gkF1cmJDrn1bXDQkV1qadXwNuoXC1P76SVU8u
v7kYPtn8kDcUDnEaRdsq8XGUEFYMxf1vt5zn1s44X3rxk9jGie21WMBx2pk6q22V
S3scy4PtcfPOaCpMFhPsHHPHiknGep/7oWcX/TOMu1JUxhXfpitEdPmCpmLxATOC
mKq0I7I7vdpfPZ4KT8FDVmw5FAC6lp2LuHg/V2LN6d3+p7LZNSnL/fjrOWLIzj20
huKX0ji88npa120QTd4SKpVEVNGellkOuPB3vgVWgUU7yi+k/HpYnkt9OmiisT6a
fn9KenqYWaKKWwFnRFPziYYaKkf1I+Dv7uokdtZjsHW963lVt/vcT11vRH0EZaqJ
IJ9i/XoZQTtAaNi5UlVbqvUtR7OrcBPDlj4WeS1M6Y4T87vEJsKuB+gwpMi+aCv0
5WQ/YFQtGE9k7LT1T0cpHW/ong28dMzwk1++eJVasy6m46r1CftPAJFgt1Aog4cP
muGbcgZ1IbKb5Ue5NDMTUWgvEBpqg9oes980MDEv9C0mIWJZawz1Z0o4zNuhZsh6
yTEghUD54LJO0j9AZuRARFsd2pdmewvhBl0KLmjU1wuNhjJVzzeunSuoTg/Fbay2
vXRGsIyu+ZVxxQJ+D6a/FA4jfuyfJpsmCjyiKNtylILn1fQ4ZyfKD850h3DzFajE
I5vNtODMxZV8wlFduKlu2/Sn3zw0WXMjsOvdEMbzO1Ph3ZKTKEDp1ubv2rnYMvDv
tTvCuEHVRttESFX0yDPa0u81XOsZ/oN7gneGi2qFm6lVd0VnvKVItWeC5fIr6PJT
jgOWd/tkZA8HwbZMJPbxzZjrrWB+dkXwTPEUJ6AX3MdRAsrSmsvVNWQdx7VgrFOv
5ObJHtElvVQzU3Nqll4eFA9xdkkJ3EW6M5fbVFfG/wznCTjnIMxv7YgVb6cJ5/qi
UAgBYf0QFTdOtuq3xEjSCfbK5+vJ8Qt7iXPw9Uq9b/0FkeA0SRy+tCMbU1l/1Ibg
SKdmAG2PoQ6dRm8hQjxlSdNAeBlmvypvXyRPGHcCtkGk8Yezj5JUI4JyczmFLnU8
8qrUemhmuVqml4nD9/wu8FJ91UKHAYwuQOcHUFxrLp1LFimck2smCDxmYPCBBuwq
k3jwrYUAMq2RHygQX6gn3BRw5zSqzF8QtKHDugXdJHdDyOWhYyI1Ll1XFww77BQM
H/GRjg3/dULyMdMB9JtiNRycanmvTTvqnE+LQItTxAryEjWR7wl9/IkEh7QjEnXl
75HSA1pyWAEWdTStXkKcfM1/9h8856u7OFqMfmv/ZyG261kUZRkkVAf7vpazr8QG
Mp5bJ7zCB/foHoTjOxVvmBkpa66FUjnvBvcwf6ARjB4IDeTEclsHcX2bUigOZpen
s7XsOEZlf1RvTTZZQz2mhO1rsRu6e3Gu+DzqpGMtx+lYKJHsM7YCq36pZvuVevTp
IN+51vbxnEu2fV7K4+rOilvIu/AVZcQ9RWgSKipIhY4OhdFPY5GdtvyHkR2t/Nqh
Q7SOdftU4u/wrxkOIXSpK9p5pjvGi5b35lxpgwmdPB2ibd596qielKhKfLg45cOk
35wKcAeJ2P1y71UUCRr6UY4cHZxYQ6y/XO12wh5gx0RPcJB/eYv3o/KSqFlt/Eiu
6UZltgBh/yGDeU3wK74CkbVRskoU4UjEfDdzeoP1geUYbzwDKJFGEZWGim2Ac/0E
Vam57f4AN5ORcoKSx6HtiumL+uORhn0DzNYEdOERrR8Tqr3w5cebM7Lhv9hTBemn
+dtHiTZ3m8AfTWgnopQ3u+C5HkCkWG3Lt01C1lD5lRpfNQnEJ1bdP5n7gslMQDzq
iyHY8aqF/OUMQeIj8V3ZwZyypJ70xjHl2tt46Xi9+qxkte9i3Q5vwYt08rqDSUey
QCfEAWH0B2P9HyYlMC/r6AR8vK92DbF8Z/BCKcqUUke1OTV4tRRvq3895dpnRk3Q
MBJ6yOPFsoICslQPeSoWS+t9/zTzWW9jluqeZFPWRFmYK9tHotQyFcYKz0B8bwcw
gmSFSqOV3WQRHX+VJJOPPANfyE27KeJLJ4JWimjd97E0UGMD4BjUM9USUkXpEa02
J8l284kb9jwBiIN6zE35PQbf4COFjdW+ueBln3UtZ2puH91nQgHkG/7hA0jgbaHN
FDW1E3z9WnkK7OiCezKld9C4P7pqqwR/r5Yputgowx5b3Oj4WU1gP7Edm1RcvBa3
3DvwvOlAy9DvMgTcKYbdjCPCbGnRTCEhntmUYDy85HICaAKV708dOx9ZdHxiUSwS
yNQy+oSKkbr6moZZK6d+EQbwBWFZo0dX7civ73YVlK/sbuZdCv4PDw0QxkdVNBOX
hjQuIc+/LS7+uTN8FHhNGtTP3GxqdLpkwJM58AloA8VBKwVMbSVTcHlojTULhtAH
6qbaiUeAujyCtX5BxKITyozcWXPqpFn21UoRQEvxRX4UgbJVdNsQVWrl4QRr+Vif
Gebeg1fTq2sX0FSHh+a9GrLRu53oARbu/jOq1Av3PI+2FwU/bKxsXwAcKZWE9Wcu
Ao93YPlnZdnFMfU55l1u137EZposUR1i6aQ9sKORm7ffBu5ai67DhkK/BTr/+BQZ
pRPmBJU9H3v6KAkUIwZe8a6JbDtav8+WMS+zG/W3a/3KlLLlvHdH3yv3BC2bpaRK
YTjn5mPMeDvUJHfGE0zfVFPOBySha4oHAEhNUI0Q0uVnHSXWb3TVDYvL9OXszTkl
8qf/zCmvp3huqM2xKsgfa8ESbmCOdLIKTnFD91drLl2BwcOrxY66l1VCC+eisABn
ODeWFqAcu+yo8+pcRhHGgvrbGc6e5CcUfTvZIPDumvTSvGPOiIegKtyguqX9RCl/
KkpIJKsB2RSkyruSgiyB+IpwlYFRFt0QJEGB7IHSPSBZ2UHce3lR4szGZtvyTKck
PDPy483+u84URYptbyDZW3YVBhkxbNjZn9JjGvbwXDnEvfXtyBridkDXPJWgtR5R
PehudJBHyqwiEwsmsuFXqBawwNKw7LnFu+Y8bM64cD2w3Rb+5SIb4u21VpR5PYG6
yWRKP0FsFG1PGHlSaF2Vj3HNEG0+APDr0zVDpl1edRz3aec9ZEG+Wy30JuMJcrfz
IX5jrr9k4qPHWd/JPBL0+EardbrHYfzkmKeFWAjA9Os67O91jDJhKP8mU/9WFp0g
ehLUBxeqGqy0xJg32WhWKwbWLeU6b3mioIM2a++tInAORIoE0LRRdK4N+FiD5WAW
lxQQdIo68V/qCg57Qeiuf6fSiAvu9LNSjirpoVC93e1vw91kZZ+pmiM2B0/o7qp0
QUYrUb/GZqh6z0rc5H1k7QDNIVNHggEBBUlGMmzDYB8LwUdzfZibtkH22mZo6VdK
HcNclJVwxWOJldvOEHaWVKltaRbm2BS5jOmoBdmNwEOiLKZ8B/itrM0Ax4tveKsE
HLumKxwu9qhPz8JMCM4bQLMGbKiVJivnvfCuFoohjDmP4GRauZ1Ki621HSc/P9bF
KICYn4dDIxdnA1WL3RMyM5ZcclCJ0VQ5b9D5+U7QZH0dCNdHDlwWTpDHMCBn0yie
l44Cnuzog2lpxfcj4R7vPEnoWUxTX6VQkO8XXCYF49pdCPxsKKOb8Oypg9w/yEKk
jc0gttY0Y4qD2+GBblYq73MU2AtCaUMrKBvWB6furWB+NHBUqfZhpSncav90sah1
IxRA/1j/SOkZ4NvAXkLdXCNn5kWou1a6XJuly+os/8s56OkgjccPFMxRhfnyaYc5
kTEavGPsbEMIQsIWyzwfHJU7ZQOVBDlMwt5GwSI1vMjSIr/f0JLvx9x+EGoSWH5f
7XIGkJju1rgo+Vr0K3uz74eY4m3Qr03ZllXehB5+1C2vFL7Rb4x893ooaXmgdiG/
EJav5kN1XottghdBJzR9yZaQBz+goVn81QU0gbOsLsopGAvt7cq3yYkZqxNTVhVf
6yBGljR4SajI6m8+kosTyehdF5hrhBPHYNVDJLJkSjE5iLQjY6m6tvw8B7+K93mk
ERurzgJaRss+fS42OtkG4OZFORwLLmysDrKrwMXGcKZBg4RN4aSB7C2VfNQWnyBG
9cByG4+Eje5FvPtVO1bmeTI0Be1pgLbqjCqh30qkyXGtVFjCwQ1n4oAS/sfkM5bG
SgoUVaB7dhX9z86BB4T6lyw5rSLCTAHGptzXF+ikheDEFPInNSw64RQIiOIYo8BV
tW3bOzh6Nj0aZI5INkPDXwIQ9OYb07pzNTxPx863q83K1gk44wi1q1LohnlG4qzo
QCXFbHVXPKA3hBmKLgBB01sFgKnWtUQN2haTyCoGujl8C3mc0km8wZCWBIsxofzE
0+C+oOxiwhvq98MCZfvJeV/xpwEo+SDDiK5gEedOpBXm4ChmGv8ZiyMdWXzf2UzB
npu3LikhW2nWHvYeQHrRUCL0/9cMzmbzOn1ksWScCGRDTaVy21xxo1RJTbbFdpCK
5pkzv5BK5piHhcNkFOWktNqWcrFOjXRRVTygBJvOHQA7+vljrgM9Xek8Fwim02/K
Ql2tGceDuu3eAlDUHjiVuNUAnKP14qHb5XrXsuCbpFKpvvy5j/JD2tQXgueht5Ix
AJkdwvrYZvohyPY1E+kyHcz58KNUia44GCbO4znEroS+/PUHngQdJI+Kc28PrQC0
LkSaGxKCX2qWu8Bv4lMlp82K3mB2IatrLfXbv49ofqUSMhEouUjXtBbV5OzNTgwr
jN1S1XQMEZGL1IN0IlboRn7qkJnmJp5CBbRUxFrtEYkJRfCprliX2regatdfM4cT
QiUHGy8X7qNtTmdgMe1bWr6enUyhpiAitzZ8fjSjs3taXbACz2AV/8zXNryjTN7I
S5sAKAPaIfY/jiAUFQiqzEFGvz9xqrgrWCEW2D1X77MI25p3wnBfjTQk49td+2tT
7OM+JebzZTqotrQKCkvI2Y+cZWL82JvlOV7QnrMyoN078cCWKcj2Ihwc1YDcvrXW
rt3F4jytcjPiMPytUl7Bn8BToTSPmZhDQKOx/UNzAPh8RlZPNDT+CeRIl1op9myg
AR3FHEN8dWtMGUWs+dhCFVJKLTgo9vHBSiIbQKOZY1FXo5EcInpXI20eNLbLiplB
zdGLkgcSc90u/X1VHO5wPVaXjo9lI4zodvj6eXBOh/q2Qx/n5U/W663rUDlFdji0
FU6Lf+4WAShhoKGbtCEw8qD9dYrOboQEvpb6EOPP8ZVJ2FAmgYvLy30mGRUsI7I0
dVSK95pibZUF45Ytl0TUuWCUeBsCwvZivOzQhJQv3l4FUnnOq1NMH4VRmCK4n2/P
mmV0+GTUZdxBTSsMaNAQv4BUxRYVf0MroZotd9D87YF13LtpQmcsI8L3chQ8Omom
eHRvwzdRnpPHfn1swuv7wYOrSkQmAfKX/dnALE33gmYcRWjYhR6H5e/DW5h8Zt7w
A8QhH8PnESP0Z1GKdJAZjrpFrbol1z/WJDVVOtsg/IUnwtI14Q74r2DU//y7FIbl
BJPLNEEc43FR8ve47rBqAQ5nPUgz1EIZc+TU+gxuzemX96qHps5rVQxDNqRBtw2h
DfKTF9gwWKJ9yI+KzvrTlqLZ2cd7h9qe6QRHSItppN7/7h9YoNA4zT4lsetj6KdQ
4sQZKk+Fy/n4OospI1e49Eh6MDcedsMN2272OZbdaHv43KY3bpkeIFIM3Eho3K1t
LTwyve0h9ak89R4/fttdVVeQ/Ub9Ij5Hl7ohxW3zb2e5qGu5pVlBBPjCYPXnhJhP
/EMqispWtbL2ESqWUR+65fuAa3QnuvVjjjPWeasVoyV5AIv4EQTpzl0kgy6YLKZy
4acjq8Bu5CkZlfYIVZm/rf4y4bs6F/xWWl3eCe2aUrmy5xFUeb/Er3FFvHIVuz8a
Ilb7s7pOySxVVEeYTVt2eQKFJWiw8zBkMLU7PK4XUi+FpJkdLCDu9UVq1J7IIBWp
TWg+fx4G2Gk6bIf8xmBQLYIMJkQF+UmVo1j/0v/WBFHH3MJiXu+VLYxrkHJNAV2X
OhTpYEUSQS81mdtEDGvQJGqkrbpmXM+KNRThUglf8o8GuWudx/6Wshe9s11pL6BD
od276P7O0nmYX9XchRktxyvJ33lgYsIoyle079uJHiIATAt+uWSqa/BHjzYPNltK
RQYsXJpKXp/MqUo9HPI92CwMMOgpum3rNs34wdfHQkg25iZP8GPV5HpV9gzLnc1Y
nTLQ36s2dghxHvlUJEgjMAOcEzAMUWeWzgMu2ZdSPSj/mGESJYWejkfc/QmwB3lb
gT03uu/IGyaerZ6Uz/wyeT+ACkrhuKQzvLisU/9Y1hJOukgBS5IOpEs3x+HAUWII
pV0/IF6fqy6FzlzBnt3YfPtMUllze34DVoKf9sF9ElK1NVCtzx80cu3cuCPBpjoy
iq9VhlHKCNjkjxc8dYXbqiHmNBL5MMcrWJLSeALRm4gQd4A/qjWB9VseZrse4qjh
Eg8/R9WYeydYCR8szyOiYWapD2al2lpvZnXPvscQv7J6K3wOJ0+WbxXGLUlOVPUA
yJiPyoWaSyyGx3AnCaFjcs6WUqZ48oMFvK64kc7elZM9WzABN4XGiti5SBvD/gma
5jMnUBQuGr7C52W0HHjApU+5lga+ca32gCJi5IpPUMvVYNGJLT2akl7cdegjPzv1
ZAXPM8Ki28w1qI244T/UqbNFo0AtCuBGaMsKkT9eDgflvIHQCE3qGdJIndqlU/2g
JY3St8gTkp0cAyPV4e1DhWecWZahMZSHBj2M/HFBK1tWoJFGj3a4JCYMjKSagkr8
fxAMbdYG6CGzS8TZIim5oL5SvxUD4gXnBHpXHy8ILfRQO7K2ao0HN+otLH2NVeuE
a+0R8HeV8PCLjrvtwRUmYzYkSKRjKRm46xHhVA06PKQFLtW/w6acbtiZWsuTowdq
3EYd2oT05eon7uERGU0pS3FSpIl+IlcfO4TD2AGPDz0HNCMP92dT3tMbYXM24Rxe
Czz/fRYbvI3sl1KpMB9QwGjEA9suSZ6IHyEMNPohkwfTwr5Yo/pqcGSkUx4Fq72x
YkaxrYspSXaNX57NFeFBCYcIpj1ngBH8Hps94Gc/v4409wkz7dJYnmyZfFIqwQ6G
2dfaG8MjCfrjm/NsCh24iXyyi6nYFdhbIIGpAJWCgQ7sjWamn993o6EDNVOGZ4Vh
al6Pl5FwQ8Tq3YPTfBRqdynOatMLIesAw9F/S0uwlacHkq30GW0PRk9ET7OLGQvs
YZ0/XOEBX8pik9+il0e2+wryv6QlMB4GduPHIPRyHSzVdcqcc/TT4Jw2miz/cb14
802XN9ShFElfTRG6c9/Fv0OaVDbuPz8FJDUaDQeQP/JGTG1UOh/mvCDlr/EldVFZ
WFTJ1tNeYIbb9if0hOFfoWi3BlIjVb7FOQkvJuJAGWprC037f1nCNfQboeXb/+0z
x3yx6iS/bF291/OggoSqKiUAtGhvJ/Z4tA6/wMcDLPMS7y6VokDNdZnd8SnsZz++
iBiwamuFoZ4DWDdhSGNZI7ZrajwQW8fkDzqmE0l9ASKxnDhLU/nj1ASpC0BM4Pcw
/7wLJFGKEzDMdXBDHBOIlZ8vs+zzx74Inr3H7iuZWTx7OQDxcQU5vaifd4XNjAFZ
mJvEQnJgWnBVQcBqds+zJ2AKtkqKutQE0fa/QMTE8S4vY1GFAdAtBlY3xwVeHtEy
0pALus1Gzzo19w85XUfi58Y/Re/QI+wtv9bxXClzfPvaLNq+bnSY2fjGPTB4xJvh
AqMZxmR/28uxj5yTMC/7QEkS5WKVzdyBQaeIC3E6tTMRlWVA7wDqsVzHOW1Upi0J
xIoaoKjZdl8oyY9MQdMOmAtz33JVllg/jKOMLz+Th38nw0r7uZlK5EF+NXxWfgjl
BYyJ6xK188lvVHEbjYBd1nWXYcBLvPjR9rahs6Jz1AtSc+5hFaHom+/tM9Lo+yKx
rgi/hvI+VUYd1pxZa4kRxLcr3ZdierhGzDx1dV07NzeEZ75anPKb52zwXAUn9V0K
4tBbAJBXET0nvOkFLypvbVl6f5W/B3R0vVRs164mmWNnq96Qts7k4NOM2AO3Fqki
iVqppkHJJ6MKLjgcYIAx2Au+mXLWBJBxc/67wuJBCBHnplpYHnk3rkhIWy3BeO4F
HR0lhEWSTaf902Ft98RxxWdhsUU7i6ZaGnsr/I32zP48wiQZgdJgH78c3O7mnFHR
2ojpZTJqKq1R5Dw/tc4c3pAaYrn2ItbhXhRie/Ky3xjTigPcI/3TPteF1fy5h5xm
IW1SoOeTyjRvOQjF9jZM8TDpoM89x2kWd0dYJ9zmEi3yTNQpBgAFB3achO2eH3W6
ND7yylFY+OCKSTsYdJNIq3/7dAYXzGsFNSCcjCZAOyaQxV/vTWegDFT9dwO0oB7S
bflxQlTTlRHw3+TDiUEbE4ibctB6rcqkwhO6cLUi3hkq2To4ZWFQrCmbJ2wNmAAp
Q+T1d+G8Vnkd2YZZkmYJyjUrn11+FMWg2FIjUKq+p4+o80YsH0u+8iarCBeTFqsq
Mo5e8cpGkBmVe4dbzd6S30zBbIt40diejm5m0FXTRZip/BBEEWMbed0ZTGqy8SlI
EMXhjqCoyQiDarrzjKR5fNS0s17ZxYjBpMv4/Ke3rIq2pCNHOyfUjudt8/aRztlU
mrSaYKdQm98i+PebuEh4+U6h0qDVrCFEBq6g1kMV6rIyguyKeB9oJs+/k35Gc3oY
WytBoJESVF/P3FnMjkVXMXBe7hfgYq3jd/Y5DwyCUIYaQ8ZifF/I2Qwe/wPSvTlY
zrif+jura9ztRUy5j9IKuEqpyqyvRp3U7PWVddWr2SsOBN3xtujTAqY4o7fZHmpU
/uYXEcbEez8MwQToZXHhv95hd2t/zVcoHq19qDxKDsQI0sXuklEpcWCfmQtCDXsc
xM2DTtpT8Mxb+DWAt6r+4rKWIHI0pZ0l85Wa9393X8KgK6MY4js5NwMXuiAv2Q9E
vYyaTMBvTVuFTDGflF3LcJngQPGYxUj2EUaix26fQAuW0J1uWEErg+umQaduDXhE
jDJfwTztxMMNvGXFOAFgtlcyYLo/Lwq7vnfq8Y8bsHSRM9aBF52JFThKwVFvrgzV
0qzcBceoMEmkZR8bKu91rcT/YpQz/x8YpqVmaHdSTnSYigvGJrTnOgPcy2OTCU5Y
79gCLzBPMgMviBEw/7gJLoY1h+rtMUykMDsidmhGcJO8CuT4oR1tf4DmMGXireSl
hut6k36hbswbim4AK7X2OW+vedi4LZMr87Xb31Pj1upRmT+59tDdKXg3TeGNtFsy
4RJ9klcHj+fjUmB4zdMjNG1tu0rIjm2juwth2zW8DbLVq5XAoXGupnN9KqHfWJna
xRshv0mMfHU6NERRd9453XThAxRulAR5DUNILhmLos8dDUkI5FpG6ScdziVscVV1
ZWXxNhjOvf1aP50lMVZiBPkjnLDzCsu9d7FwrVbG2S1p+XFjMkGGKZx+gImg1g5B
Yja1bxeLu9wZy1G8k5s8MZmCqpQfX6uEFw/yAK+bRSixYITDLCGPfIIkA4M33NnR
hvt3unpS+2g4r95LsiaMfsIiIbudA0WHoyRfVE6FJ7PNpvgwPzKKahCs6yD9U6+S
hiBRaoq1vezHeVhQ+rtTw1cubSQ4+Zeh0XCFgnrdiCCIfk7CA32qJtikaMLYoSek
dh7pn6QVg6oqwRJEerp7TC53IIrxc84T48aMcioHhGKcYX1rjApmSORdaJK5rZas
Jy3gLASt0xiT/t1Jj3wGZd/sRtUvoihA9xPtWCDBH9WJsQXfHQIVmaOGOE4bGASJ
gZKNa+83aMfq4VMeFoJjvPJlBgunM+7L3oCWJsX+8pw4TCW9olKjY2C/HNBj0WgC
qlbVVIOSG5Suw6agHF/JdAZJsMFvt3aDtl/KhkP9ADGGsc4ontd9PUZ7zxESJTNf
KjrJjKUKBHsHZfytcw6IJyn9JwAe0I5IbK7dCEG4udEfypHR7sdb8MoabMb8yAl5
J99DvfeWQusDeLwISzEf4dumZv1ihAB3coFAoexLea2PInOCppLJx9o63igqtoRL
A/Xo/XBHG9iq7NaWdJd4cmf3iFR7S4vmEQ1j1v5jiPDhilwVgojHpmf7ARLuoSCD
tIDdRfzZbfZ93eq1FPnuWrhLKyPYLBL/Nb4sqHrlH4DPx7kfGtOS27RN5Lia1Lue
pvSSvEJsaBziv2GWpPuoLskHPB1b+noaS0W1xGJKzIf4kPN1wZmQIsDAMPaQfgj6
mnCnYoCAOqSLfL+oWn6eT2v61u6YNzQhdb8hrhxVvHyKb78D8Q0zqMVHRRfEiQx2
fP32EOUERq0LVOUXmncGUVFh6mOZIc64TgpKnVs6OvgHJ3pK1dSp2zc2ZanlDpmr
cQEeOjWzTw9Jft2skBYdmA8HlNeMThDK6OeG9V5XWScuyjYJH6tDeoYvjTUoVejX
WcznBwwMq3Op0efmjjvzk81m2ciorSgHRlwIQlK8jgdlPYDUVBAeX6JAtvWSxiom
OxVtV0IibjTxM/Q/xQhVW3GKetEbChvgplXCj2OWkT1FyxmNwPeSp4bMqrhZHehb
K/nQq6ez0Z9fVqp0eWligP3+E3AxR/r5zZvRU3xbzDIBxISyUgqEZDqOHPZmWuiR
V/sph2uBMh3VokzGoE17KU8FS0kN99prAhn/mcVG5dTDUH/gyyzD49NzuYRqM+xX
c7ZOY9uUHVkBYZl1yajkjcw0qpdKLFMzR2Pz9IVNK38zbJfWRvowdxWrwL7kbCit
zq3MbEa/s183R2sjUWbMO+gVUD836OEavc9AyRc9r7WcyY4kq7cDOYDS2zVJLrKJ
EhvMQ4ySU/OBC6BhQkO8uRexhUtCYDZkjLrktQt0clwJ0KItvgAs/yM4Ac6JwTl5
M2Y/pdVKVprSwqNsoLimaKz+UyWN7Va3pOqDjT/1GWRMsI6UKD6Em3QdYh8VEICy
3mJdYKgL1QrERu0nd/WBrySJHNTxlqYxisYNyuDIpEB7DWtXSjntqfQkczPghZtF
veUxJ/pJhwzd1kAPg6LwLxF4V8P2MNP36LvIjOKPndPn5lKf9+/DEknJWQ+iA+1M
4XREMcYg+kvYEB+SbnBZFKRcRUCzMl54iwIknKAN+VEBV7iQFDEurvJXHSQB8RSG
Jy8EQAIojsJCu/jBG7sxoAGp5w2X1TSuArSTjCwaK91BIBvBbCr+VT9zkLCAOgkM
7SLPxrHwhuK5qilJoPEdoldek9Dxq1GeEi2ozf1SlXsSIpXQMmNArvaeMrqPHkwN
NTT54rIXa/ly+fxDOnJhxJM06GoSqqVAPCjTbwVXikJ/5F060flqUgFItebXZ2WZ
slsFUnp+gIYzHXU2Z5FkylOuzHlEZHG/cjcTRNSHsfBZqyVgM/yQPnYLsJs46aDC
/QSBVCiSad4zTcufxt4YRBGeatkwuC9+Ksw3LWjibrLzEPr/jLA3gPkxtKw3Ipjj
dcZIYKxLNM2sjf3ghcnPselSFfWcNuX0JW82B7kgA/FxtnX+jO9nzKan5omuP/2i
oHC3SA9ip1oWu/e2/53fykvKW/VbcobM9zIi57E/YOvazEyeDR9osafyI855VDzT
S1Qv53kEvBwUehokree3GhqiTOp7WgOwpHO+4GJ+HbP4SM4m3x/N0eMmRzYsfRcO
uO9uVA/gLbTngO7zh+1bHKi6rEDTGmaBjWvkwLVDdCjyb5Af6Nzke8RORFkdHvSG
j4pPwO3ZevxeJG76npMVgt/j4XnHcOE9aMjuklvMVSieGm+kt0cedYlAQh3cI8PE
tgKKw3fhHeqUQya0u6zNtvBtjGn2qgnewLHsS877lp8eNSMIdb+2MMeUX0wtc8yF
4uRFefzKuzlrhqtOJ77QLjECPw4/b/T+scp61tHxKxmaUBw6FUABLHcVFQ6i2xra
koo+XOuPJ9haHy/VdXX53cF/PVlKqgKbSfZS9w0gtMxKYSSJcsW3ypp0xuxWu+FI
aWBNqDZ8FvF1rQpmqB+Gs0vLafZ+/0+k1HceXM7b++PEpfxjpJnNaNiGxA0XyO1o
UuagFN2EM+gx5Ys6zyJ51Cg5dRejFkQGpusDfd8LoJQRIS5IvF2dV8sS3UkSpbRU
PwxjnzpsIBNAdqwTIyBEhS49FqU4K2p1Y7RXlGAMBA+VyDj/zFnjfcddMKJtDF16
ci1snfOkRU5I06FpOpYQmkhVqje+1nL85ePXY8iQLLvA9liMHBO2f5BUKXovsDO8
SYpw5GGG/Beg0jZE9Ar7RslYqbNCxdYiKXI7dwhMirJWW0aWS2ao2zj1q02b1zzR
6xCSEvfyJT339xczoIOsj7y4jtfQZNJc6PFgxyzUanfNyXXQ66OBOFF/JRt0/sD3
C9olt9D1JYhey10lnVCoRGsu8Z88kNy4IkBmCAtDRIloLU8XY/Ew4xTOhJIthjaq
QGzSQpLYmLFHfgSFZzhjyK+T7Qp0iR2fVIumlGpOeCYCLYQAwk/EADpKSlT4tfHU
4cng4h/xNRwZML7XUlP4HCQKWnBCSnU6JGyWPEOfuxGrocilCk1jUWnLryNfLQbr
UQAdfTBFB12Zky/3/FG3SO8/FyCk1V9S4hx9XAWIAL/BNnbUDcFKXPO0q0kckgvv
MKCRA1B+kCtuVEQdQePfZjiWfP2eUhMS+t/7ieDo4HPT6QbgdY4PjlE4Z8QbtMl6
MuoCbNp9iPlTdEy+ezCTYlL68sGwwrCZuACY6TykOWQLnj7UhiZChivj8mv3i25B
SyH+eZnoGbQlTH10GNKveTTfKmCz81n3NmcH3nPw6VXqAAY1y5SZIyxPLPTNEydD
gHDp/927ncXiRBgtFCsPURFmKJwM2afxcynZRT1WFD6OqOqw9DDKdhDhqKcuLk8E
visYT+YoPGEmuWWdh8ORx3krgvevjiqKLMWgW1+LNrSHI23ailnlPQN9atrWBj3P
C917PpuHmHN6C6rvWc/ha6VhOFuv2AxwcVtlgAh/+aBYCcHbcgJW3hUGaIpxxEFY
x//dut6tKm83+AydMM1E1uFC6N43O8pg2UvdvraBMK3AMsOPaP6lxZnwbRuq7np5
WiNzZhzgv72zAFYzQ6QJsRcX/QcoBnzhu7dyit9+f43a5xszaMYPYe7cGfNlyT0B
xiDWmUgbn7IG9O3BJopAVHVeP3CEvaw5rMKTrOZrggkcFr/+P4greJE2KpWuZChx
/ErziCW52GV48My1Jl6poYZMPrUwpcNHtcmp+HU5gOMKyd5hf0JgzOM22sPgZWj3
Vv7eienzE+watLLIX0YJjqRmgWPlR8xdrZqxs47umlQ7EGEgiBLFulAJLIGISebH
h9wF0py/CJ77rd44/C1W3oRQCyIpaNB8g0meEXU+IRrscpV/2sCOqV7DkO8Nrngs
FF4quwLvQo2Lbu+DIqI4zIn+aBMIU/mXV8Lt/DodWzIzFZPPD8yQYCcmkS7kgCBb
6ovpx5cK5cbO5B+xwssCXNWX0ELDBysYTRhgPN7t+A9ZDCwfVTd29EqXZ4lncH+X
GQg9Aep2Z7SBqpuPpb1C5Jcz1SccVglhLLZoTa9eyLJgXRMm6wouyqfYc+tKS+BB
l8KTnUgRtUbibP7x4mMGJu38v/ivCQbh1uJmVJNFh2MQKFYm7nBIidGImwL8tiMP
0o9lt5sZTcS/oeWBC573Ln1LkmE7E/h3vlxMcQOyfMZkl5pxqrftPeRmkQYQIZrg
7JxzePG0VZEhnEso6TSZdunQEyjRkvKoo0DRyVOKx0TuGN2/n0wxTS07uOYMBPQo
UjwqT0pSNy3QEqXyvd6yO5yWhZ7YCdgLYtvwdejfkbJzmYa2tzDiJp3WTikVzMnB
BpS1I6/IG7ewUo2B2Tv4hxuuJ6Pu1KFqpib/mt4dxZbXT+oS+iPz+wTrlfQeMZnI
06/h+hT28UyF5mBEde6XB0aR/E6mMGHYB2R6dt1nvTYNyJ4N+SkvOekDbGaM21IF
mfLBhJmMbsIgXx0W/s7KJD35MQBb5lsCAPcCZA9zl4thoB5QkYbBBiP5VVrnn+Yp
lswIDMhFOp9Vu4zjQvKyE/zSjh6rtg4ropIPWJXt30KqfywgBOpSX99VX77kSfqI
Xm4kALIMo2UubHJSsAqSq80sEAKDMj/cO5sWVjpF3/S5l2PnhaTu4m9KmKCApH7E
zPa3R0AW7MJ5SufY2HFgFKn6HotU9gOzj+5uw5CoV07WNa9i2c1OpITMwRBCXnax
G1czWX4WGtn9F7z6qFKWY9By4BBvL7nvbjWz+RBC7rdsGDzwqdh+XnOMEZ1ehFi7
e29rXautLhZoyIu0NyelMhM6194xUYe3yg3cVQb8Nrrgi2jtLA1aAbAyZbvlXxOy
DFWZahoWc47zUEc83f/fzADxl6tdr15+gnBaIPCDNSZM6j/+hvXcnstsufvj0qEG
Zfh2MdDWTz0rVm4CgE4fmNbCmNrYBgPSqKm+Udxu1iCVv6ywGIC5ynjMk8AA3SJy
b90Ri7ZBflVyRdmuBdNQayPREy1VENapKtc+dcKiwpjzAQyfusJ2S5qugdTuTBYQ
tZ6M5IylFiJlZrk26pYYQGY/+VCW67rY9bWKPbHxGSU/Q/QQYuVZWiZAdkrdboXE
7hHkj5osupao99435uUo1CDNEW/PUK2hGSIucuOCmuAAusH3ojDFfSdj+TMdgb+g
8hXKZSXyajN2R3dlcd8PvbiJlmFFwQwg+KKiaIFZAwg4Fyx6ryLdyzIWbcU+Hz5m
BXGhDAq7dfSUSFUZCmbyZemM/DgygFisdj3rUq5s0tDrMcFl/bQqJXxo0cBjrnI+
yDL0NtQJaj9NChewBVPHXTT2gRZrkmU8BMHR+BIM6S3hsxWE6La5PBK9gOutvny8
UbB1UlmVcDnmJ2ZontH/iDuMl7+bWKERlvb0Vzv+Smc5qlMU8CHZ6G/fRtC6+o5L
0402YmwEtZulrVAtMHEHECu455C4t5sPbFwT/BCP0pY3QE0+4dBNCCMQKoLDZ2rn
`protect END_PROTECTED
