`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pM9ihJTXyG9tkVxiOpPp4V0om1m3PhOE3SNiW4wEzqugGx+iSgf6g7VBTf7njGTN
I5o6l6GFFGbH+AXqudFukqZ3ikxltBHISML0dmWcFlTnvZFONR+wVjO7Nnxp1XDl
L7qvUbdkT774P5YO7SNhrIoSWayQUsLihuL61M4zcMcW2K5F8bK36+OL6J0Jf1K5
048jibyR34fOKirMIReS+C2WzMLLwNS7jAwXqdKEuEo4UIwNUgg6xxXQ+boYDzfj
4QBnDtu1K1OiQYPAZvT+OwijM9PQksyBCourXWfkDRngaCfQpofjFK0Owv3bgPvQ
lmwOK/zybEbS5RyFRhplnJXjJqv/xntqNIJr5lEBk+1JmM9FX98sMdQ6T3P7TfDX
xM6UW1Fop4oAT7Pn8c4zbuUpl7N02rEYUWRLQZb+h6MnQLJjsFv0uZON+UHKXZ9/
pzqVIEPU7U3zcmkCfS+Orpa4HCZNRczsuejJmGk5uzIXUDgxudqbeOeiziHHm5ha
BvxyXKzeFyVISKhyFg5HVRPoeCXaP4vllVawb6PDVnouHYIBsk9KNS7BTHhmyD7z
yVWvDNQhuiuaXnC2OCu+C1cfLtXBSxKIc75nPU67nllFFic7iCXJdJsbNp3Ua9g2
pYOMCPPZXgdvdbLJpnyy30TL4QtRFJCXOUkkZKfUZNg1hZJJLcD7Qw0pubufsr/c
OnkbVPxBTTO5yiEfLnd5D9nYBnrVJiHUdZGRefmQTOL6FRdfMuHn0Tj4EZgoF8nC
aLREhnb1SH2WFv1OYtexQHWSHHIJVzpUjfwnsNVEjUgdfhkrspgviIXNL4WvYWac
Inm85ZnXMa7oEcQ5zbVmKLDICPZsetwZUfDrUJGf5Vd3RuYvrhHZeI8/IHwH/VWh
PcQcpfNhzyaAMKJYdCZXpb3xBL5wp1zf8iBfEYV5sGs63QtJjYRKV3DeEGqe3XqE
L5pqYLlTwAAlGzwyK1v9UrZL6TfRytOkgFAVXhFOzr7AF55JqwuxRHv9hUx5CpDe
chwIPzMwp2RCLo2R2S1oxyaZD6GSFukZNmiRumQqYHRIOd6SKzU/T2wNtjxFNT6c
EsyFrDtlcRGpJZSqg5feweahr8c/a/NKgNx09iRcST65BmI85q9H3k3Sinp2Afnn
OW6eBHrvxiz3kUi7SE6820OwrattMEH6qLwI5Q2CCTON33jNV/OXgbqcz8uDk2wE
fLwUPKzs3vT1kiIgpzQFSFI7VpddJcFLV//MOBzZ5Y6BzsJTeftnWS++juSj93ts
s/46qmL9C4yd78lZxtqugh2TUqj/eBPyCFAex/9zwk+dX6nuKKVMRMfKagl8/84j
zIwFk7b4d0QH+4BJemLOtBnYasDUng9ILrQUnzozW0Im1xLrq84UUXuJbYYQIDtH
ZMGsW0yr1LWtdNZGwrLajfHWzC37oXWv7xR5391b7boAEl0faqVAm3UuaV32kSMu
DiiKQTqQz91umLA5Gtm/LgkNcwY1+Gsrf2ceYOfsPoVgNCFYm+Z0FN/0AdqfAZ8T
Pcg9xcM9WQi9i9etsoW2kxe+FWIBUKK4jIN4MjS6TkMfGFoVwfS/8MDg05ubYyMK
N5Va/tVAmOefcjLv1AjaEKAuaw1QjF4aN8rQzp8qE3LxAMJxvbIY4uiIvIy0Iy1n
8sGkvMXJmNNJzLOsHWUh2K8R1w3EjhOobyH2lO4jploEZN54AF4bWoR16dDjOudy
ecn024bVuGLzLJuyYtEvAZCXyVvb9eEJwWoz5eEaFCl9DJz+z6YmVkgyWTljf/zK
wVKC0vKv80nojjrHndJb9/8aMm45HpKw4Kj+c/IA4ApDRhNzFfzu16/mHkXivhzW
FtnV76yyTq5A5eXmTwjY+/++2Cpq76Q6nkZfOknxbL0BTpuY5x7btJD+lerIa0C7
V3YAYRT/OAg4i9EAMcqilCnjLgtVrABIicu8Edo+Z97zBaXLASJm75/BMNwfcDL0
BSl6WIoc9soVh/ZI2a/4wDkw8CzaBXa8aeSGWMZrcDpwND0LPNN9ZWF/3Wd/cb2S
Asc3KKEMRNF9xz6/Ao5wcDUhwjuJjCBml9dHnBsdlM0Woh9gjcHiYmb9L2lAZWhP
9z9d7P2g1n9CGQa/meGg8XpuE1ixHfuXwYBnrFS5Z6ABmUzYvbcCVR72ewYlxJd3
LwlJ65E/+F/iXFnIgFYkTd+8o/zFiN5QpUH2jS35JkaStR1E2uJCovKydCDyXLxM
X3f07h2sOQ7CE8oimcFFIqcvmz+Aj08GrT7GJcs4tHLoYRmFSE4TnYbLvBnHphdX
XaWRJr/7aGRGCzqVgCSTIF2Zqn+uhi8JAjtuAwwgXkJSHeAuP2q9W8YyH7XP3snk
GI2oxGpouauTCJ0apmJX0VV38C8rt5PhvbNuV5Yn455OpZ72yjvlTeDqhaILg3b7
No+A3S2Kq97bncRO4P5ilRL6MC+qvnyHALwvoH+vHXdvnhXDObE6TNUD2wPVUTan
7Vrk/Q8ba0nEJN9FJFngvC4ioQgzvfOBNH5oOH6VVR667KZshIasmrso0TJ9sAnz
N8hf7vfZ7Cgab2bVHU5E1xU8KbL02uKJjCUrAMEnBirpFQfdgYUoXfGsz+p/75ix
aYXxjObVtcHrQksknyrxmA==
`protect END_PROTECTED
