`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
85ejNlkvW2vs5prevrNCdTmbe7bYG5D+fmiHeRLIchiNovp9iQb4FVYr5XO5K9fe
/CZebkCFfgbfmdkiD98g6E+SP62h9aQWOwz6PBGcYaib16E5UXvDxO3w6WYxjsYQ
RVuM18P/UGUIvX5wtSXXiGeTg0CuG7tinNYH2GVJwtlXWNBxjqN3PkHxiWabiw94
2VBlNZO/gEZYpOc237fqlegTDLcFH+WI+AiVMCsp6Xg8yRTsa99IHw0IzMhs4Icr
Rrt36wNHonYAe/GzahjRWIT6uQ8yvbJSvPtmUhOoQOXAoT4GAhYuXcRn+cBuV2Sr
avRYUEjQ8QzRTKdSYQiFdZ4E4ytqHEY93dZVWMpbto/wagwkFfKoXc1sITbRfqla
ADIgyeVe5F12Bt1MfK8FJkLvMfoBE+ZXlClR0B0FXmKZwIXzoe8KWZGE6MI0GUm6
UoZ18HzJO0PcQBOV/pbJ3LESxi6wlvh2gsY9SdKqYUZ6gn22NNoDzttvN/Lxgm2U
cn8nqZaknthCaGK7GY+JfckHLhKEioY1CvqELTr2hjbZP5Vez27Rp2aw7upyS8Jh
KYiz0PxRbFEb2Ds2AAh0oSybYydeHwQl2pYgx2JCNljqF3xVvQX2akC0DfGxvMBd
OZOjXIkxSkT2Fz04meY2t/qMDs6oANO3L/VmfnDlrEi75Azm84pN5ZRaULWhI+TT
wNnotWR9KCE2hlWP0HWK8aSkA7ATLhF0aHhpgSPsXrmTJogcKxXFKheYJTgfk/4f
ovdGg7Om7VUacl1LL1uaDwHV/3082uEUc7r5Yz0bgO7i/wnByagISnGm/bLs4FQQ
0cWQL6cOeAtb0TPXPCgJTZEyjfiVR0YQYtAugjfdc5JuCw8Euq1iFvbKxWSTgP6S
KMVu+3Il6e22sIAVcdj27NuRE+sh+ICPNunGvx1/zVM=
`protect END_PROTECTED
