`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjDQ5UmVPdHKhplnXtlzPDXN7IEjrA2ZrG0nor+/4FrAbNHTyWqZnNxW7rkZHKLq
nw7PmVT+zCwfaWboU9vW29PYlb26Bpl8Rg1oBDKP7Ik/VHgs1ugw33Fr1EX39s8q
SMoFKVpbwY2s75qhqVhplRTMHcAr4rDp2eu1cq4c9Mk3XIpujcQh9CUSFuM23PZ/
zeSSEM+lxu3dcOvDoddm7jvKBo4rEfuklnviHVVz21P28zUi6LXEuKh3SHjZs7wy
CND17Y2TWUQOUXQMVlvVG75f7iu/kzynHmr3TnPr2iH7OVnPv+2xEaHmJGgWTmsW
i1YLkO2nr87AT+yXyoxzSL0GUz4JYgSMXlyw5MEWdvrlo+ktNQE2UTQ767YYVeJe
VHAehHutWodsmnPtS45LfivLo5rLc9AoEkKOjijcRyTfRNCz2leB14Pe7AY2sYtZ
r2jkLHt3cqTX0HmqPiCLo5gR8hQHEAVf31PqpCvtV/6bFvil4d7MYVvoi+TyQKUX
2uVpbP5T0QfbmVhUMIXZSkkMlJLF6t1BldljC4ZbW+wTl2jWLYFwrlZWyaLf667w
4Wew4JUzUTN1KqMv19FpNqvrMSSIvD3HDQX6Exl90XDiv5QOsQsOsABzjMhTyqIE
G/cXqIlugiYUSgTYCSYEHBzA7YMJF6Vo94g5x7KH3Vdehte/wbq8FkD4CVsK4HLx
4Ku1Bs7+FGOuFFqH9gfrtrbYndaGV2PvhhonvGzZp6uHU2vbyi783s6e/rrfJ6Wm
+tqeCveCX9M9ajIRHnFTnNwIC4N8qIaMObWJg7CPjVjArzejg6dxQ5KTJagaekrV
nWA5KIm/9PxuHTmpiF2Nry/7tu7E1hNtaMJkr+oe9mrjCZt082Yd3n5g5+6VvLSC
c5ruHhrhK7OVkDkq8du+CTSUHiKEkrYlX4A0Js1GVA+lJZkQLf/I6O63CrIQ4P6L
/MbQpz0aYRnIkD+vthwjPjB5xIwthaKw8sUYYd4EJcQ/deMnGMM08QqdnmuvY2Bq
ubiiikmmudL6GbD+LQYGTHuy8I1Q1TrF5KY378631veoP7G8SixcnxeHGDOqLCJr
KKPj7NYNrX43qnyoHveup59VK5p0af9j0rC96jcgl6wcKZ6t1TwwMAOmUq4A8ZOx
+hg/Kpm401v6Tp+QHFXZN+qmnBJjR202Qk0j0aBJzu1l3zlBDL5y7DqvYL64kLoU
K9HTDdri/XaTa/S9TsN06D5upLe2Feeryo+GJVYFt/INJq8ScjrQCvXq45UezMBU
J9H2VwCvrCMD/2ABTgy+GcDAUOtlOY9D7eHNxdfw+BnvQ8UMDVrjddeLj+Zw0mbx
qj/RHnGLODahMh/iKVXR2y41m32Qt3/FbgzTq8wSZ6izFoicFHx/5qI47Dvifx61
Dz+S66BmZ3FUWS3ik/M8PjZxF2oPhhEL1zLc/7pT2MM=
`protect END_PROTECTED
