`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/tmLWm1kkkWsuBUOGJx9WT2UAJuGgXJ6yOU1s9EtEgXvI3K33RgZ42eUDAaNMwt1
Q7tZiTojZyygDXTHs3G+4/Gpi6QAc4ICeXFuwKYwHTRRiPj1hPpZoMHtb6wHPjfM
ydds15wSa1tZ5acx2zuuYSQUv7bzt2m0ob5mCTYAYfw9Wbo5y0TH6o2H3dWxXygK
6pGmgeWw8DVkDOwmsKOE19O2ziUvnQs3MpV7FEWpgV/QsXlX+Xbv2/Ur2uLOb+KI
h5jDrxSa+0cws0pL8QaUlp3IEJhQBXVSK/hEN1vBCkLQzjviT/HykHDCxFvpzf+N
0wB9XGhKw4nULnoayezlZSyHjtW/qrdjXJViBPe6pT5aCe9d8YK1wRVFqScHaa54
qqUHK297gp6792KgsUDOnP5yTvn/PQH1XmLjZmdcIFFpL5KDSJ6S4p8UA8Uue53s
1b/5NR7Rj8iEBURtkm216ca7whfxaz1jV00q6OG7Z4peFUKcoCae+t3l2cMJR+AZ
Ag9fD3AkkBVtMjkZDLZ8ZSQDW3yYqM6PXqFc4D2NSKynMWxM8PdGeyp1OnegdFvS
GJ1IeVTN0+YutzmGmf/njVmi/BJm+FlETs95Xnq5jR51OtsZTCuAWd687d3pq24R
BmZGBq9Q08UWfrnCmRCrigUBPQEXf23P8yJqGbzoykvmIRi3SRAhhMGBLRmxmexC
psz6wxi1BjxXtE6OqflCPLZa9CSyq72f+0fqgc70pn8=
`protect END_PROTECTED
