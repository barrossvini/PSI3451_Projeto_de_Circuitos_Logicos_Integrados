`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PU9ct9uBEAXipQqTfWMQ5WZtKRlguOgOrHObfnJWqJRGwzuLIYJqNbPMA74Fdq6V
y5a8gsIWX/pSMZvEWhm818BAMpIVoQIakn6SvCsIxtjXsOKW2YSVgilSTk3024PX
KWnVjocD940pnqENvk5yhTfMY/Rel9VwvXfM+i6ojm5uMMuvjRDzylEyMbgM6qsc
DNxAzHd8oGsgKPzjy83tau7l0NnmGfvqDCH0/itIdZp9D4CMo9qcxp/OhJg4gA5b
MimkLleWu6OJhUl4TgMEpck21Lxb/WGgPiP6/Xw8B5qzovh4XUjQmwmebBUG7Jda
bnezS64MrXIwO0AyUN2u4Z8V66uTuw7qkwUUYRbzuRZLuKYAto9/E/egluSpAcWd
l5tqws64k1QHWmWPeUD2Lh8EIXNeZ90viH7CbWfCFKvp5z6PQ7/sVM60ijS6kqUw
u4z6cGDvP/8mXMeLccsHiuAxQ6XZGArrHcurQsdN9kcSYnRuy1YLfIKhdFMkrjwR
slAoLitcF/AALrKqusuBUDRy9lvZ1sqDiX2PecnwtvzcDuQlBo2ycq98/nKxX7Ga
qHoaU/05OVBuAkxj32H8vASeEsgj1fkGEvFrCxFBF6d7NKUq0xkZ7FWx4X0iUQlQ
tKSg6wv8XfA0dNjJC6u561fd0q/aQA2Mq6/e31WlC+BPTsYVUi5ETslrOvAsJZjG
+wcfe1/1jcC36EUMtebEZIfBl2pkdKh4mjj9oK6ShvJkGmXVdwAhuUzZr+0qwicy
3a7GlFgUqzGBfengOLD2iZdQCnV80+Kq56zC4zb8mZg8eDwflse3V0xyO2Nh8p63
u2FeouVT7jnRqzp5J2Af+9osaTz961IPJRjGIow98Cwf7Y5PBnLL3QL92MbFT7RF
e31fU1ThcbkjoGAYCOkSx/uwBsLQ43djRvOZdPrtruJNwoNxt8u8qZbvAPNiy4tI
bOCltgNc113w11huc5Lw4vWNdBVavdCl6uaqgRTVuiJM+Oqnqz+OGLd1BWHHfE3q
4VpKuwBlN3Ze3k8jgHY0SSoaGvuUjJ+cFEwxbwWcl8IEvc7Gy0iX1H9RqN9KUb+l
GFSZxScI9d18fDQ1rXOfiXVQfKE2MxyOheWB8g12veWqwg3m/HiFyFubkgh3fiYQ
BMhjDQakuxp1aCCjmXnnFx1VC2AjnZ4dc7NpLf7VFeaj+ShuHBiYB/RCeICN9lOi
aVpVf27kBZ6Acw7Xm0srWjcKDinHF2WibIaT5Sy1/JrlYuNFiYoBhoVYhskarW2r
GTB7+C9oKPSISBbl8ojCcLQ+UpKgLccFWDpYCOPd6AQ6WRVTZpLvad+KZgRpM7ou
//RdB7TcZIRgm+P+DogrmQTvVIRgTB3VtsNqhjyhzbvJ1JNhp1CXTIl5SssMzqWq
lQhtdYI5/AcNe3VsaawlNiGZKrBoUenMpPXeKDdU6rD6zjBlBquEfuezoqnkr0v2
1b6Iu6tfqCi8/zktUMSLxYL73qvZDyIT3HX08GCBlXLNN0B3h+MCXJVB7gqYzqUV
p1HrW72U4DUbH97mYKnawHh7gyewZ7/iJiozk5ySeg6cDpepGW/HdurQ7UlHQW9t
fmxCTFNSeycaSLkJiayO92hnJigo8qXkLl06d4/piwm0T5xzFw2MesZqS27JFhF1
opCcWZjrni5zxU8LSCzJ3g==
`protect END_PROTECTED
