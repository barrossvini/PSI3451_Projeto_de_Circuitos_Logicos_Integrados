`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+7Mu3AdgE/A4iZEVaU9EOlfoVJWIPB/+q5q7Qt08jx7criZkAv7nwMMAfJgnbgfg
UdKUlsloQ5tvZjQuIrr79IYF2/1u0wBWTVZ3MtnXxk735RBGur0BNJpAN981R3sc
jrPFseq/9rqWr3cw+DcWHceUtEHPoqF/6qwIbx87wRLcYcomCkEYKu3Ya+GQSA00
pPUW+uc/59pQt4yY8CFNLa0oD6v+ufAC1GaThLWak/sQWIOzxJGpxsmsda/sX0ia
ahv/ildbI92WTG9N7vNByxHUCtKBDtlWMdlivH3iqHUyTtFyQ3hwfu3VoY6aXkua
6rB2KbzHXWByhjMb1OFJP7C373T3VeCzTeMpsu042kWXHa63TSWAYXUUcpqqIhTN
yCLDqa8308ZmScZU8OAOQJE5Mh/+ylXXsaPtoS2iamlBIK++4LQvRxLgFE66vu1J
XLZztVsWC5Ayt4KApW3IfHim3cZZkCdxnhoNL8rxM0LAQLefGHQE8wtqarFe+d8o
9RzJyWBcFWdesKYiR0M8inDVJ4GoYxJHaECUrbNSnAj6k9Yjoen9O9aQexvFFFIT
csH1BLQ/8jEA159+S8W5dgL8MD9+odpZyXos/nIWFzKLd9FTJM5WSMn8gpzqJbdi
COAmwOF3LF83/+p8JKvgHnaA4z5MZi+9hddqgRQkYceQ+cZU6f5ymAkxDkPvaFqT
eptRSwNGM1Zue+QSeAK1hUolCnGFlvpD3Yjr3DIJB/paCBDt0FLFZGxiBPlD6XBg
jF9F0+cqSVnLQuCVHb8VXDKcxfvmzTrA/0vGiI42E6K7gC2FgW8S1acKmoANRUXK
I/XjXM/2WOLmxW8d+p+164MdU/chf+8j8KUYyWQjmx+a+kMgODiMJWTK1F8NBF9y
+t+ZV+/P5gxHmG1rH5ui7N8umI9v9JzrCPybNR7yxzvI5ZRjWW664qIYfpzoDGch
2EPoqFvujnnu4tL0TEbWjWrQlzU1DPMGkNXNtOMuOecqlwWWs8MhokwoHo+RtVs9
EaqMZsk32CjfonNbGha8ybC1ejb+afPxrzTP9iLzs/gbSZn2c86klj1W16uHmHK3
6lNlt1+Hd31Y5wcspG4edVJZ/0L1u78lvjaQOHEPGtGX7xBhGqRsFmm0r7uu/VoP
NFJOW32LE2BEuPkfhVh5I1q/BLLhGZEdPLP/i4LPur1eCtjO1xjICDZAoEVjStrJ
s9Hf029gRPMyCKGfjYb45D431NePQz9mRECvbjRc7SUXl+3z7CUgkc8dXHjt23IL
`protect END_PROTECTED
