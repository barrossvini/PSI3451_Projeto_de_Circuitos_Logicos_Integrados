`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FXhGsIMBlkC8mqpPUULS3yOhnnI+Z/ZmHdhJDOYAQqUWImmr5XLPPQGrAU6hQ+Ux
D2uuIkHtULfoTt2tUbMTe+IMT0AJvp8UEBAp9J8QMEcc9fCpiieC7la76Kb324Q5
P4ceNce4QdsG94F15ozusqxlY+4omZ6NyJFdpGQNJhducgxR7goY9S+GHnr1POXo
8Mz9Neb+l3tHy6V+PfBqHhSUWz7XkZ+coRnlijabI42Z8vXdGuZAPb9UmGIbxlCB
doS/JVgIrrIS1b1lPaSWZ6nBpM/76oGg8FLUQ6Ez0aqA4IPInw3Y3LKchMYWxjCg
0tZg+BmZdO+DDiwVGxBvwNDs6KNL8wtka0Luds6EBgEzmWDfxk7n2F2ZERVPUdIj
fy/qGLiZSbxRlK4Lfq+dyjgAUfYmyhhnCsBF73af16Z126ixHA1cOdyP3dDTLGfd
QskIk1WCw3vfBdDpoax8dZaBCT0ABf2OLylnTpnxTEji1pXIx6hLrgMsOF7HT3fc
6KlmobV9IahqlqitKCjijVRRhFrVE0utYMYfVDXD1AUyQa31Kf/laqA7O5g8ywpj
ZvTqOnvhg07LqZwikLRpSAQRwOCsiZ0DoerkOLOIkzBysa74cRxv+OlYhGHB9KNP
GiZyfZD8/A0Yl/7UkZgUvVtj9uGNfTNaHdlhqtYYQZOV3Ak1gBiAwY4lzoINPeVD
Q4B6789JGEeWZOK+fFMlIpdyrlE6N2Etc0hbfGrDUYtwn+9PcEQGa6QaWoazJ1WR
4k5Ii0if+WFpV9zWgqJGRuBXMTQriE+7DKGu+UmVBf8dNmmtmdRoX3epRfd7xOT8
owwbvWQHbTdZvpOkpDCYdaom7YXnbR0QIuluyFBQKlh37rb0UXjZWtHHohHmAdFH
FbKXU3+KT3vPVV88+9tUDvPOM+dYZu9yICgCBdJ49jbOhVHyzxhsL2ipMFDyo8Rw
n6chwp+vrkEkXgELxLydUggJQJUvCKJgRYlBkAdsFJaSm5OiJCSZKGyV398p519G
7VRvOsc3sjHNG/CXrOiescntnD602c6HmLqBahoEYhax7E7sNUWiN21LygymRzOL
G+L7cLZ6QAFGhbpwN5NBisobHRBTuKVAl/pYb1HplKNDhAfboCTcWUY8jEbE6p71
qj6MeMJC52YqRqWBLtkgHUjadJvbg2mR6MHXy9GCbQCcnnBdlk6ZHj6RDJcQBZ+E
+ezkjxTCLhY9VLGfpLsLzEjfkBxzOz6XATj9pn4zKzbZ++lqPgPdgNNp8emugPW0
yAy44bSrAr2mf+vJ8Aig+17FhNE8UD89avkkSqm5Wyv66IP3CJKcSlJ3Sojf1Q9J
gHVfoAbtrGqRMcyf9YP3KLWogOysiXcbsph2FyBv5uR/2UHp+Iew8y0+PQX9cxXG
CBuR5O2/F8TD/++i9q4jCu3nmR2oNraa6Qwv58MB/VuJFPgR1q9LTFKLML9UUBGS
61jqYWsFmuPH0FXugzyDUcf0Re7clPx7A4dZQ7GD34Eaem8WFk48TQn+yJTdgyf1
sOVaTRzc0AOLEoDnAAEDD8yAYgogevxTW/NlPqA3iq2MHEgM0scL68SoNTe5i0an
5SaWLDwO16KKNoIQORjva7ENnasfD7FUEBjomUYmfNuvVEO65RozaK2gnczU5Kms
YjCfLRPmtUcIUVWIFY0rqWx+GTshT/6lC3x4vIFlOuQ3/yMghTg9xI91QH6DD68b
/4ZQL8nGnkOCF68v9cVASosJC17flWNLabWeeCfo7A4P78tcBAb4h1ALpBCY4JlS
`protect END_PROTECTED
