`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SigJXtmB1Z2zOW+l6ECXKf4YjAftCfuzhjEzGAJXHgvmj7Pw4oL4wsd8/5GextSw
zT5BU9g+bcUzeOpBsobfR69lLrsnDyt6CNMgZPnVBPJWopnboYvLUMreSFNt+s//
QeQWk4lVvvu7HpLBzDnnK0GM1O3LRy873mHY+kHarcGe0NNyBG8gqrxQkq0q8bWS
O63sWR+mYmbWkfZt7OCUfZR81tl2azXo53nY94civ0prD+3DcUwVgiNNeo2bK8jH
Y5h64hKrFRBzCWxqoGwf2/TdJto6nUMqMcca4Jqt/zHqCsJ/uxgplLOhKbV+MkhX
VQduqyEqAjmHZbrLZHWV5bg+d+Rgxb2zRVs/pdtB0+xAt5outFlALB/OCSXa6bFt
YzIEsTaalkVcCQFeWf7n3sth2VmmCdR+Ed1umuucG+pTcEGpGgUJR0X0IPNUFzVv
RWZw2qXU4J8lI1y64wbzGyHT0JNnR9J/4bTS2upZbxU=
`protect END_PROTECTED
