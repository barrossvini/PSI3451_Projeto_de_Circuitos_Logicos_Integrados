`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AXCT2dGKYWKevSsh2Fy6Y8r5YmUGi9/TpzQ96KasXThrcw9M/Kh7hSdF41g8OBy9
JjlojqOWPVc0QlFFAe7C4j8L2q/pmPwKNzP2tE/CKllDpAFuSxaiJVoQRFdsUQSC
6Xyf+3JtJUJUaGDvrHRnjKzaW9PVMehV/AA9lm2VwCK57VMvhy9t37UcQbakVyVh
UbOxvA+r7dX8vkAtJIPnWzNFF1vLTe5fMKcOCbwxx5G7fIMcyJwYRhPfHk2WEj6d
/KA3d0nn9B4wWMNoCiQxw7+TDjNJKBK9be/AcXbiWeFzBKYIadqvGjNYpRQMaM9X
HIk6NmIseiBhPLGoyIKwDuyzEj+LHHV5LZi6eTNRWR95c4wz5MazTo+LIFOZJePh
tVJbX6CfMU6ey1+5M5Q0e3eOUN5WjFuKahdoCxHKTrPfCZn5wHClSY+rtgbj+4nN
VLPEFSHp1w5NKZhYehgnf21i2IIia+kwdBw+yh6nLLlFgz73iQoc5JcbdXZPK8mp
oCM3Piah6cN5m+P2yyoRr20gRC4Ny4rOJKHEyDpvj6f6xD74S1PvE/kecUzbu9xe
f3rnDdG/u7AAyRk+LLnwdR5OHWvd8DljAmZq0RVXBAv2iBof+X2D1+Uy5jEYiT7L
wlLcGoF0zmJ3xG2+ulZCQwHMrmQUoWwBwE95ZMipHTZCX8NN+UiDFM0pveR4+LwT
hRwc4lNlgQPM2c9gU1woiKtLxuNHlpenUw55zmTwEmhuV3CpgbWbVi7a8Epv3pMC
vYERytdQIWyEw573qqyqZgQFxHJHygMnuqTLtVUujVuquPdbnUjL4IS+DPG6ibep
X7Ra9WfUWiR9oUeQK4pkSOS6+EtlA2CBhxNscNInUGcLRug4UuD3mtW/mDzF3QWN
EK7JsB2kXVUqCJxb++5DsU/+KCcgRB2jED4TOVvwilp2d8yIc6D54aiLbjgs7Qsu
7BMM6Gwz5KVnMzEOOZnkH4mdksR56tUamUQhVGVTRnbsrRWTBmAu0k9lAjUyIuMi
UDSMbbZbdETuwoGT/Y+8/WSEnjt+8neCCXzC6nfLt7BB+2Cibv5XanR3fZaFQs8c
epwz+Rl03fLaFGy4B+V64q7beloEFuMaPfxT1nZbYXPBGUHTIehAHDD9mvodMAoz
9uQCdS/GRsQ4e/BmtPTAgW4pE831WIDhdN4AlmGIm/4Yp+MZ5DSYGH3hLemeycaQ
by7eu0RqlDfANXAuUGQneKA55JU4nDStj2fiWyLiyG3Dz9HJaDco40Ux597+gAXM
ba+aZ8ZaZvdG/0UQCEucTOdNGE9Q36cOw3EDGcmQODadcSzHwsuDydPy+y2G/ak7
Cn7S5+4D7x/CBACpL3mBOMGR+XKFNS2JOlh6lZNl+0d89xaOod2M+7V7xsSLkCXH
bhp5TdaV6oz4PPM0s6yPJtI/rs1Uqe5r3a9n2T+n6yWetY6W3vXgU1Wv8ZL2hhlQ
HnXbmFBgyYY+/VWTAZzsYliJMv9tR7J+7Lwm4J6KlQn4qTuV42iXg3qUBZ45ti8V
//MR0fpHe6/taQ/iID3LbK936uqOPLd7MxNruVLSbA8/hdFU8xzRmMTW/V7Y09xm
fp+1Gtp92iBVv8mmHuu5XPihqFkIKpOcC9H9yXfzspAcyL0KvyasoYcvJi0uOs9r
4lc680mmyC2O7TXRbutvzYx+EOYJhAJIs5N8C77kWzYeLwcqlr8NcGr+vbx4aKa6
V9cXkmJ/uyvQz6u7Oc0b/ptctSCOzR/MvoqxCpuNDgSeZz9A+4l7+uqe0if6e/RT
1Co3eyr1ApczT4aZmO2cCiLSGwAbQiyf4b+lXB1nPHuvZZcQ8aCZemDrU1H6gntu
7Gyrq+qE1+Ff+zOnh05+0SGvHPzNx/pjn5Hl8ECO16HeJKMyWqBy3rNnJNudVLhe
/4CXZ/DmyE1Dv0zUT/I613gl0iW0V0rTuNKiFRdN1A4cK7EZAg4d8WKAS4mttLHN
YKo0IZROR5+dBpKNj7TUZgKGjdoH/Y1u3oz7cdQ5h8v9tbDNcRX7cQP1RD1Hjso/
DnpfT3vukdTY9DkTL8GDFWQAp8ei8nmiUVRYHN+Wyf3uvYWbFDG2NjVCeQB+COIj
VLK9DaAASpt1K3dvjPTt4enNr1uzIcj5En6IpwSwMtSKhRQkcmjBBdktKYZecKAG
mPRi7pZN+50XxDjVCB8EcxE2Dv7rqNzJhyX79otXQ5nXYM3IhV3yHOXbZU//IvM5
7HT5WBU6pzokqK8ER8TEdxqgMdvWgMCs4Sv2ojlqmdN3LT9HiKVtZFIrGm4rlKmg
++RcyMFLkZcSxkj0zdHRJtgCMwtho9PesJin3bwQ/ezJZoDp7kvN+TmYi+uY14/Z
jhzWitzngMJ5CP0YlEaXqrDaaxt5dRRy+gYmmjtc8yndhUgFozgEX03nzygw9eDv
NHdyEgKM+tB8JbAlarj1PlSsp6F9c4hFk5rCTEr3m0vIYgYhTHqJLZE9skfYgmFD
HsHfI/0fvzBJCc9L/cWcT4Q99+nEN9uVGrTztALNZzRks3nNkJtdM9L1MQ9BItFc
a+McNAzPG2h7EYHDWQ2RHgGkrG6wweLCVwoFYPvC1HOc7Sd86x3IE6rO/2YKaSWK
gGayBiloSh+s6eI3ih001a5IYyxb32Xbdbg++6aJwBiq8O/eNex+jWTYofjdMTTi
YHI2LP4hsCUDMq7gsqluwSYSFu5DlgQkpkFxyNVj70EdbNNcvutyj1hy4On37CNi
JFfjTPUj84L92UcuS4zptfypso+eaG4oUQjZ+4gI1ws54kwuDuOGs96peFvo52MA
DSmRSlULkO/DKUhhsnTOcDhWjA47yQ4c/n1kICGyTDNJ1ivrozlvd0dqCKUGVVd4
ouNQZ1NlanuzJdAZ6LBFkwvpM2coH2Xgt/fnpwwQhjFvyynDuuC80drQ0mgiFrat
Pdm/bOF8JUKPG0Li3BlWz8vnbyiP3ESeUmjliQDPSH0VupIsW+KR3kvbSczXR8/L
ernq6wWhqOH6B0Je2y99qt7WMSm8tnHJ76m73XNIYRC8Ea5mjFeIxdRtkknW0Jaj
9hEXWiGWdN794D4RFrp88uPpt3i9v4xBOXXXlHXNIF79BBHUC8bPjjOBG/u+arfo
NRL/lPtzXN+ISAadX8Vi2/S2Tjj3GJjbJg93xIlgeknpVFURXlsl/BigFzIbHw8U
4uzV4031WOZ6VAdpXciifBo+BOcNofndXZOM4jtHp/J/4qtMvzO5qvCrnjY0Choz
xjhNKIcGDCt9mh2MIai7+HFBZQCJ+f6HihS8JJx6YglMK7F0A3JQJtirsWg9IMXY
+XwmrdIgnp/K/2izbtmfaZ++qIgUmZCOiRKlymsFpuf6SlX0xwss4fLxIY/JzpVZ
b2d4N263BVzfOVDy6CzJkBx6/My4k09PdLVxDXt/7V5vEBJeGvF5URdUgaztYfin
T1Nuyjet9zBM6PrIuo1d9FCqqpniNkIFh+GrEv4lGLoz67lchtiHx7qaHPqxXxO/
JdkH8/fWk1g0T789wNmWG1CCX7rHvg8oviNiXNcqS7JHFUndM257LX4JW5LzkPOr
CYwJSs6b3bGi/UgyVfVghTFK+ocm3LWxmfglPCO2jPJWs0EELoCqOpjnqcnoTLEZ
4G9f0tsJj+ehozwwdYNjPoNEIq1d4n1vl/BkQX0Dls7UeTROQI99+A7y0yNYbwwG
X0eSeAFch6/C/8wgLgFabby3L8BxtA7tVaut9ae+r3PWPcWekRG+vVAT76Ebbytw
Ba3Zg478ncIrT4bZA9DsXffAkfsZLE4GyLnii6cxvV76vjbJaqUaPqN0r+yUQhXm
By0om7tUZWhWFGx/LYyhp7MbqOjXPJ7nJd+d/Pgwd2ngfnLzGQ51a+ofDBcQ+trN
qGfGgbAs19TsFUszGHQQDKQKyEKxqtpxZ/diTDtOOyTOyiXKI7JVzlpArI02CkuI
MFqNoJ7S1qvdlF/zaDa3vbIu3bfn1PEPVJLsBboH3itvyrKUoxSZvuY3FAcpVKeM
h7vInbYeX/t50d/NJXYe6b7I97CLCWeQQ5HWcv8klVyAixyzZJJdUe99qpO3YRJP
9zHaq9TPTNt2Ei1+pR0jLLdqQAadUToH+ME7Sz3tLZPd40NYzJHMW6GFaGs2gi9+
9V5D39F96HjsI6F6yAtTMCP2pE2bILlUwcSkQ8R2Fmcl8PMdyi+gn3dGxzwfnG9d
C8NiyR+ohBky5fFKh6gMIUl8NwKsyRhlYzl7mjCMwLTxgWSfULlwEalJRqQewV2h
tXH1jPBlY2AtvEPeuFwCcUFLivF/L9rUKPhQ51valw16uzzKlGV+KQCyLHhcwTVs
pcdcZvdzF3+aVvU8BJglV2VEqBcoHtxWSI4ZL4/aOKrDjJWPaKIECYaOckoI6SBr
Ps/6jaYzHfQlS6ARpG85bCm4LGXvdtox0te3nHhhAVUnip1XWVKZYxiAdgkiEHkR
OMd7AtkH8UDwGhqD818m7EnsxRCSg8iZbgSER+WdzUdgXRrmDCloxXdvq2kPmd9d
UzP0a0zPcF1sxbX3dBNG6YzZENkoKIMKZ2S1xv6sllGqTtP4eN+VnocCgPEIiUSO
ju12z0D7UtnHYfMleARqosalq/EJnrW1VRx5pUqBE6rUlaSNvOaFqw00sGPUwmPo
avp/H/C9GaOPyvSXsSreEX2CSNaw38rhh/Xf7IwYHZ8rz/To1xQwg6FXje0Xe9gJ
3ZsbPLJ7PGoL13PkCUWXvg2jB/OFJ/81DDs0nC/VrpmZSO8QsM7lxd9aijfKmN1g
T2CZ19d+4AJSvLx2M+uyt/SAS6TqTWSIkDd+Kz2UgeVXVKWZKusS0TAWCS7JIupE
pbX+5RuJf7aV+OwWHsiXI03/7JVw1JWq7+/nIQKb6IFr74ELK6gfveOPm1D33TMc
WeL9bxYkKo5a4mmxFlvZbGy1i42SFjcDG79Bch4DgYsxY/giTreu/kBOQbRqE3oV
ZMcndaki/qRiP262jyeYkuIoSYlYl/IHT29bDYcgw4qEeaQnbahpubCoN9g12nt0
4kViiTqJswdI6TkElboo0T7Qqanb/271OTm4vcFd/2FCMs0otVWACtn6vDvnwTEh
RYp+gqkEu8LM90Dtg9eDtNhtsFcapuUF3Phcn/0jWha2ODse4F5gWqllsGJWPggh
b9uq0maHDqfpQRQ8JACopTlGvWp0d48hCOxWoVo0Hmf4M5eACjyijHr5P87eb7vL
BL4LG3ZslwaxAvaDagABdknsCgQDQgydD3+kRf4iENELB+bWBE3eg8GzxqoNEWaC
oYwc57S+YHTT/S16fA46WzsQwkpjZWrP6UC8NoIP7MNjVFCrDSAtj2diXYT8x2Ak
5Kgdz0+9L1Agp7ZodOO1+iXyjdLrILyc7Yjph//l6YFRPr0cmzVQ9p8lhbnmAnRC
jO9bh34cvFRCYW9a+PVunfXzY+6BFWcIXQQrrWF6ZprnJ94D9PlYHSLJNA39YJIv
OXk9ECAWHZ3kSz5tokWN2WLHQ31E+hVBituKqmyrovtd12SD7ZwGocdeCx/AWFBJ
o6GdNIUpPZakpnucFysUFtkEV6V98iTL3ukoZORHd+GibLUpdNjNwklUP0Bol61/
dwz6QFDBhLQ1uog3zkWWR2vE9HOs2g1mXcL+bLA844Gx7/DRYQr8bqtiwlMCaMuG
zjnn07iC0/GQIi4AEY2LUu0re/Ww+RyB7PeyzLVkYCDULD/JShuI9JdagCQsDL/l
LMBWLL8J1pAT37vCOeieGPLEX3WpvbPmuWZrqF5KL4chSw/WijcwUkyiu2ywBEXn
Cwr1oXSsijQqhr6WUIfZq3JRTcxAe3oAmJsezctrS0aradqaciv0kOOxGmUueztH
rHnvHHhJOo0ZhHfXFZSROeEtfO24cGmBjLAa6MBhq6RghshlYCgyQSt2GHE9dqi+
4BCIMe0oNYZGMET1D9G/iwNc8EcRNzkYYklfMCBNZMja4ZPK9hxMB+4PLf418asx
gXKhX/dvbjhMMllfNb1qGhOPfFgpou7dyPjc4YAx+NGW1eNEkM8KH+F8ERPwjEvh
vT9cTJO/g+zklSm1YhA26lMzaejHtvoBMJIMtmiH3prU+2y1Rn4FbnOB1wtlomjN
JhFUWJ1abvPUWgPyPjgBlbqKoFhF6zRbiuec6w0keoPg69aZWzs4nmKfYvD7IpsJ
X5TKIVheOy4NjEMWX1LxgxyXcYMnfSoAHVjpOuordcNea7OZamb3MqCKhLIZm6ZQ
4ALuOwew37vLE0YyMMaHa48Rfdw+b2CUc2KWfjVLWlZ1crsxJqHd5CybvHK3OLIa
NtcpN/m6lw5dcvt9oJW5YNy/jvkBdMDyp6TedwEqqIQtviWdrCv4RRsbNE44jhwW
ljsE2/5Kh1n3CCw+CsA/1LO1gVlDE6Wwoz2g/qjNgWv0T0WvluKiZsG2Wjv5j7eu
tyHxRN1B3fUtOsdzuvQ3Fzkyw2sDFnuf39tS1NXZyNhIdmiDUCyBuIDX9d2OJ/rw
1ZRcXU8oyZebjMNl0O4KcSSgMEFPWtWgoiQrN+2eeK9vyTVHjar+eYgDjf9LeDiA
3/rH58kXaJg0GPijPiSrNU9ftjJfKAtbTnBHOhR8wC57UO6WF089ZqkXqClM+lln
lmbHWRJ5gl4SmgMrHBwckOehmfSCmM+u5hmQPuBYQ/hRYzEWjT+oiY5Cx2jt9ksk
3qwwT8EI4SbS6EubmGGu/M969FUyIy2TSj+ekE0wjA7ZAkSYYsW/l8DfeF3nzx8G
XBwh/r0IFt5o6G1nn3NhoXvC0P+mYORpi99rchxXVK20Wb3cJQYhVC3nuImQGoSD
mTS5ItZniuAeSxeUCtQV+iBvDVKVKxCjfHBvsNBrAuhhCNWWkdTMCGyGPSTXqMNi
sPQmWRYdZLRPrlrKFFW6Gz9qHT8P1Yo1aDF5wdmNOjywc0jfr64JAleNQoavEdyJ
MLhc945hR80WtHuIA6AeqDbVbO7q7Nb9uZsR77b1buh75vgqGB8K9u5IhC4f1Fmc
uK3O1ePtKw7JlorfrvokcIsrn3lDlcj59vePYwlLb/FT6UrEHZWXrnYNRPAUIXcm
oQ/5B8GChI8lEMzsUeOf71lq0EIAZWMvnSwhtdBM+pd3ppv4fGhFFVAyog3QpRck
O3gEuhbxSascqJGgX3FyAqXECJfAvJ79BJZO3q/Xy2/L6YnuExtoRgDbHJPBNOns
xz4j53TVvvhYC9ySbt1DYIDKbeOBbMF24CZGGv9gjOrz67Wmn5Xw5tGxXIZMVvPL
EFHTaviWM0j/PF9e53rrC4KmW3erJVuCLzVw6yj/aWbL9hNjo38fRmljQmkxueMB
FuG3NVjKCP2SUYyDnHKuSmPnCT+BY6QqMGwhni6ApShk2lZtqhMHTIENMFeywrwp
6ElaTtKWcnobdagpZnEP+H/pwWyqwheq+SaVLAQ1j1BJwYd8q5IREbO7U7Ym+GAm
QruQ21wSzgvKTwIrIvwsUgmvtscCbvRNgZRygKVoc+0rxdKjDsLD3Ap4RlvGtDzB
tN0C5NdFVY2AvLz93LOd/9ws5j3rJ0773KLgftXyQFM4ILB9n5Uv+xqSBfRjibh1
udVqwRgICHH7GekS/jkifOgErVAwrDjmcGKwmeLQgi/2xn5q5+2k9HgtF2iev+Bg
dhVrKhipZ05HcyVOHGzdtJG9d7SOQpmFA3Ghm25IwFaZ7F2713evpGpUoEhWpH9Q
1S20R/JhWqJPVTjhl3d6UBWENoQyZUXYz0oeoDP1kIxszhSz+fcGL5R1MCNLoKBO
WOqLmIU/UnB9Psd3jy73qEBAyIA2tdaQELsNgtaMjyMhVzNP8FVgjaoT2Doaj+5a
DPvgFftO4PkW2u8vPmjg6miAKtqXd3Ama9eYfDBJlFiMVoAwdsMB1RVYdi+I97gM
Rwm2JMIfEBdoM+UIwjP4ITLwjA8wqYTU+ZiNJ832XYlCpsszX6TMmGdTSHneaGEM
lPhSY+SEtfPckNSX2jm1nYUUQv4Qv+KGAJ6GYz9Rh/1EJYvKyWSFS9cLzjCYgOUn
39YuZx7OAM0t1H3acxbZiyBeVAgzHVdXgTQ9ePRtQWjEyah2msPiT/8ULLGEQ61t
LxzzDbV0xEQdGqFoC5+wZN9esRqw7IBJh1eprn7QreCudyTcGNX24NtqV4JcJ3+r
k498Md3B1AzvPWyD+L8OQBbs/m6/e34VwNrVUkLCzmwIrci386jJyHZq1ItNWlYf
1i56OVLE0HXBq/LmeST2jIO+L+53CvD1iok3auBHZt+nnKzFJuWEsNw+x8CyMLAW
3+uywkvq9Iskn123Op8yZqC03JWt/Svqb1UyUs6I8eTu930m6FoCVtkxCh4bM11K
XT9cHcs3v9jR+0OZNsxuskO+dO41kdGlRCFILfDkqkgozhCMYbtp452P62RHofz8
TbI5S7uJhgD3NiY3BQ8F88wRZQ1MKqakJClNl3wzB+PRfKYdr3T5nzwnfHr1aTzq
VLmLIvxNV84/x4YtZ97rMs30y0zEUvT7SgP+Dn22TAxnNWmhyLi1P66JZUE4mCGZ
3/V79XM8JFJZQVdoVGbBmIdYZQrMegFbhJ6PUSiHknP1ipaGaD+CIf2FHpsFhgUW
yZc/2mxUkUBQwL2QLXDqncOWs0CYZVPkP3bAALFJYTt9AjAx2nsiTegnNuIR3YRI
pwSyP8VD5DtRZrrI12do6CdAoMeJb/fee3eVxoMcXvSsA2RUkXJq5G3zI96bFWAb
QMZ45uTePxypYoqppKa4N20ohIp8qGFfDvGk5otDugXssd/+BYzWf4YNgQkoWcnu
1WK1Ai2C2BQ4dBzUF6rs5/62IArv/lQ2HhoqOPBOQlhhazNw4tcN+jEcZtEXNOqE
hb/CN0RMmRmqLhtCK2Kww0h6QQJfJGelQWQIdRpw7lgrQL3EN56cpeiZZM4L1/in
tIP41qatpxmowiy4uXBB72oOyZqL6l7b/MWx6RRxftbEhBvAEBuXfiwCZ0C4BnL3
1hYBKZ5+4qP87nLqTv+XQM5S/6fQgU+dWM7g4fsRezCuBoCZY4ISxTegsetag1/l
HvaKRjxApDXWztn/FvyvEpawkKJVsjpY8bd8mk/HzMnB46xZ3ARr23iengnDIeM1
m7r28EQnNSKP7GxGVTEHA+ZuCFgBTaVeh/bpnpQuG19M9HFoDNUQGjIxIX3xVSZx
6uqLUGdbKztfy1kJ1W9eUDJ3aeUwPRSRxUNSkcfHgQb3IehDSnkbrjvQaj2B/DCq
gSk2BR7qceY3AKdGHxXNp4k5kQDJR+ctW6XBkFfcNzJIuoE5E/l00q/bmvub2bGJ
yzieK0z+hDHydJqOFO/9fRmQk0z/7/Xoznn6gZ/3EdW/w3DxCQkn8Hzr616fol+J
ypXKEHXEqypEaoXdzgGCNxvJuQ0zGfxV/aO+srqvtIMqoFc8yJtD7Vgi4ZT3Xtdc
Uo78nQbvmwa4/idM39sYcYwt8V8A+0sxfje3QLbe3MF7LtpJk6EdKincDSk0NIdY
WtrdQty4OUZko1RYNvDihk/7QwD+xOhXKHNl3JEyLozwiMANK0GVDRt5GJ1AbEz1
JK4cvko8KOVVXz8ZF97Sv0unNgQLdEEuQJ7AX0Ucy+oG6Jywfhh9t5ytypXiw4JD
H58+DfiNlyH8YiqxP3zWwGf+DWy75La4NvBOaYM/ZyVU2u2aLIw+Z5tJmZZDv6nJ
7XgDPqGvBmBK4T01XQkA7n46lMFzz6t5BMFVqPTpNiaVEMc7UaorCsQVYm5iLwER
FrOOxrtFKF/G3X//yK2CGpk82gZ1okbsHWc/E7ouj2OxNq69qHIVjJRyGAsW9SAn
MiyIyZf6zWbvl3l3CyutOSfafuPC3NWASlNvDav9ObEqYPSPg/X98ZbVyKemZC5P
3EKTYb7EHfcp9aRV0j7cJVwK2dRU16+y2u1RZd9a42UWhmU4Nqvct+WqbnABiznv
i9enN78fk6XzoqNVkIadM/3NuZLPHg15SqC2BrcgvVtZKsvPm2lgK/E6iDNV9wSi
XHiBQYp9ylCoJt2yWG2HjwOrZXBqSX5kZO3XR/Noc8Vp1GKiIbO5WnJMfTEfwkG/
kk3UBaQ/IwVNYswt0HJFVhR2WB9KIhxXf6RyC7U6EU2r6+HIYEQWYx5Xn2ylsLB2
4aVLDqgpPCYQPsXHBwJOH7csrne05VkjKJvthXrs1WsWPAOPGwKJCrZqdRs0Jolz
D1zQtg1jB6SNJadG/WGYkDGHBDPOp4R/3BEkMghD0W0OdhDfPDPj7Pm+7M15P0sm
OBoKFPLee5a06AfymlHmQ4xn4+WRoqXG4zxM8b4ju5HmudfVvxSyNmNMVQt38EFq
PoSW9MGcVA84RVhHsIIaG+aWPdpXO6UT8xJGg4FCeCp5J3rIBTL0y+r+IVIvlYlI
1pfxL076oWhxFdbA2reopDKXY53I/lcLmFBmvjgUCPze1cHIapWa9VvhLxVQ2BX1
qtvxo2XeQRRFc07cLAjYrq04SytSzNz6fOGW/1mhFuJMpAcW272gRHaNzml5vUxs
sFSBwJstYYpnjQ9cHIs9uTEbww2S7yROtGrJRgApOvwXr+0tx+92j5uDF11SgIkt
JZUWrekYfmwuQgnR0TY42amQttCp0jm9hZlIGtXq8z8Hb4/69tcxwZlUf40hOT46
yZ+foBe6lE8HmNGmI+wupN3DUSoYPpTuZVoP0FMoH32sRU4logUR+uySn/K8k4VB
C/MPPVWyzM03Eurh1Gg8UyZuHJjATzdpIlgx3Vzfw0nJfUSm4KU5pKVg4yWWYhmQ
/7w1f/dr/n695CE0HIRcBH2PYFl7g/uuJCMzufJ6eB64pRvOtodbQBs5RtPMNU0T
q6qOptqzy/1LApphMVHZEW/aFjc3CinPQFzTkA4Ffg1RUzh39/X1erGvcpa3Gj86
VQ0D7J3MlW32OMc14dxdUaVLz33WZJq4C/9qlvJpK/KizjhUBFQXh7U0uCd62I+c
AFkJZwTmYuuPDlof6x7RU1kOZyrMuMz8/WHB+JfFvdWCRqOsDre9nYcx7Cz0QrCr
Hf2mSJQKrW0RA5iwymz4n4/fEGfVsU3gO2BPvP/W+TxGko5TSNryqaJQaGyyvfnI
ZXsVs6xxo9KK2taC9NkDEyJVYRhsAlM5l9GTHbgPVq0TCcI3xU5A12XBqAlQBhD/
4HWN+eefldfbg1WIQFYfsqk83rWTvuX6afy40/JlnoQFka3wKIcrDE6getn002Iw
paqluPg+77AJNM3J2ESdff6Kh4fRaomynOhOvz3d5x8NdlfUpxFIak/4qdpC1v73
Cyk7EgWNVWHJy8gvG2ABsCU1Xvqc7xohnkIIlGFtOvfQV1XG0Py+ndJJ2hoF0Nkz
kxOiTGhYdW/WRFDTiccGPsRPBbAo0g10HiL+WO5NsztjwI33HKm+6+b4VFEJXGB6
JzwafIp1Xipp5OrtBYAW5PJqpdBWGumda1QX9harw4KUg0N2k1Gb6nvAiCjyR9kz
z10Z8aKZS8ZOj3h/0KmnMv+sNIYTz/AsQuiVukqdAfJiCCWwy20J0UMikrcq/DTH
jA/lsh5MU033YOQr1KX6PWZ+g63PcsAWDHBKlzaP4YOyeaeHrluQ+syBMjoNDhdO
o2uMaljJtduk8kr6tntTjw2kjb7CGLCxWNKA33UyHyIseK7HzSETjL6miefcZTZZ
JhaiPy91+jGqy3NE52BgBCujH8bfRpVlaIlYdcu8ZjXLRRSFoDfknIhKit2nd9FX
v0rCpFvV7UG1oVYGqTRzoaMVrJxmfFc5himMiSIKvveAy0eTNrtD7UVwcYeiEkjG
PGXd2zBVbTJUICryVLbxHVoAfko4zl9IUcyqz/cSaPPblLBiCjzNHY/axvdWJlOt
TLoC0I5fCwbu/FC+k/QW0ZwJz1SInx/xlHgejYSFfHFTZAa8V4UmFwdbNTaQvCV7
uuUHlRtsEKX9La4sIHqfU8vXdI5sKhA+w7OplngnV3992WyS+vkRirxxjKTt90I3
5T3cvuim13kWAqwjWd7wvBRdwKZsa3j5uR0249T3PdxqQnCtrhvwqqkcaB0gOU5q
qyAShc6DCVdjKg3yWpiXptSY6mhsFlavuxeoeB8LYJB1qtH2srEWHKYRatUIXpI+
tWfHIEGW+VIRRYPwSMrS05Q2hRcNhzyVviSZWfpkfjdqDqM2fzu48zptsjm5Pfm/
H9mxyo8nmhZ2ZfI+aJmZ3/PR5VnqbbFzqEggQzn5g6cYrbPE15W1XFBGlW7ZvrDa
tdt3DKdPV+qjz7zoZHdrAfnBaTOpQ8RU9asT5J0o08RSsrHB7o4uc87UrheOAPgg
jITkRBa9UNF3A20aaeJcnfa16hv4xYeHsf8n9eDPYPLOen83ZrvIdluJZU/1JJOh
CrMUAIqe+cIIk9TNpp3FRRbbkcgdpx218SwxSFDrPPija+lvedC4+l41UjzL7nsz
R6+93d+OhT7lzAAVhQ3DRxB8oDtXjGxnkUiivJRFj77NrbBY6a8i83+Iw9hK6n1l
H3IgruECxPMeAfHS5liHJaq4mM5qF2ItNfSdSUqDe3Q39d9L+Oo+07Zfcz3gabiB
avpKPHPTJ8P4KrXU7NaiaNDblXbCUYirsaWhJd+ybAuLJ1XtDVcS/2KSQct2wqEm
5WSNYXfDC75+Da9el/RYJ1H+Wr8qq3bCvmOb56zbbisxR3GU+ytTVoIqmRlzb6SB
qKiQJAJIjE8ZWb7PEq49d1UVcZSrxF4ooui2F7GyuaayYo2YPf1wzmjm1zdiMe0l
OcjKnto6phMb4EnElHSRurBQ/wXJAgw1+pFn/tHxTsjkNOjUEPwHWPkXiADHlN5G
yscEyGbmtDXz/HRs0wUKM8LE9BFDrhjK+qdIRZgqvle9FBghdjvWGzba2ZiuZU27
4CyrWu5i7Ree+dk0edm7CHngZ4l65op7bZdiGFsFfyu+j8RO25KmGspKBAojPuw2
TMfePBkIzv00vbg++e9JRp+ZxqUtQiFuN/KDI86ZyYV8xstUcPRBobjznYC9abEP
kFnwi02VkGuxErGG+xafV1ugV84uGZyTFMwMOStyfqiSt8TH/YSb1U+exDuBW1L2
jO5mX5AWGi4gTwd6xs/GdgoYWuCdM9HR96gt49RF56o+sPmFRI9bh5I/0XPgwayT
qs3lAKPL3w2cGYShVbwLLObzVHjFSGbN5uAted/XI7SY/aVUBmYVEUc509LIsUD1
DABnPRz+6p8z1s8Q0fkcN3L254gR9I5v1PYNzayGcYqXZI1GNQZgYxw8qrDCCdBd
N6DTzSG3h97TWp2lJX/BEGesm3gPTlbO9lhAamgFZVT/JL6fxh5Nr2+RGKy1J8pJ
q0uAHPYHNsqxTszDglsrwyPZDbAn89FdWmJ1/mDNb2IEO3HuNaaayXCyffedBWzx
GfQclilDKTFxFYwoGNr963sfZtGHgpxWWPAmjPDxILTu/hgZEUm1zO/bWlWtLqWf
eotAIBJawIttIQKECGraDr+TXGyKaY4nQwu60qli0gPak+78PeY+YQxTY8BwW1Mq
pqUiK5fDBXclA78Y+4AnfbehPqvrV0cEBX8m84heV+ZYSjIbZ0LpaWi5qQnpI5zt
2UKxCbPvc/CeyB01ZvFq9FKDlJG7zscsgE5njcPpC3yPULUvKE2dbQP/WINJcat4
5z6jnUsR6giM5zDwzA9K0QwoIKQ9xJeX1YZWq8pHa7t9VzHzZrEZ1BjGaeXpdIB5
H4cZ/rJ2BMFGQYtdmFj8ApSYpd0U86MFQ8dXdKQXfzoFHF+UN7koIe8jJnsxKIkc
3p3HisTAKuJ5XUO0Q+L/IDXyUcDzvOW3kx+41j1sUNJZiNSJ5kYRIVR1ZV7hT7ou
KS7DUxYeHo4CnkRUuE1sWlRK6e/CNvnZ0IPFbZyvBZF5y2G2zl64r20YRxZ5cECc
McHOuwbZE5s2ShP91LTZ9X9V+VoEpArgJMv61fUS+tL89w8fAVIKKi55YJrXPiNs
5Dk6i80SFhbi0QZ6aRKL/3Ym3G0UYjuGtclgoifyRxVlR1006CBM00SzVkWpifrC
5lViGklD9k7bEB89okZfSw73LYTgPL5pDFRV4jUDPDFRkQNzYfSyPJuqLR/KlzOJ
CWYCR0BaeaVtcpCSVzrLeiKZlYFyaUhOv2T7sGyZRrAPu78ERAAQCgTm1s5GdeSA
eZu4K4eF+lrqtD3kFbGln6uPoGzQNWwJ0Q3U8RVHC90CzVGa5RKboHZEaQWax24Q
3dZwhCll3O3cmtOixQgKntVZCHprcSMMJ/zW3Hd9bOAzKvzyCJgTeFMcBisuxO2V
8XiHNaKWUvh2HLsJVgrC/EdqBmiRn9la9977NEoAUbSgk1Zjyh+yXXW9P+b2TD6m
JpSxfpvgrbiQRkGIPXHNKPyXEcZJda71fJwQ+JfixrCze5a2IgMfn6EJeligMAmX
yvF6SPFmDf7j6Xboj86bHxwhTOyLTIKQ8hVRFbukZTtbG6VIkw++dcAjcXmigeSC
CQpkxaCWpOMmnk/2cFFsAfaueMk6dseb7XT7vk6R9rV5YcpVUVs9umW2Ap0zbZ7X
kqx6nULBCTRQ6o6EjhFnBHjFerpMzn9cM52n691m69Z4Lod+4aSDLK4XosYHY0Zw
kHJwCJdt331b5co8Y7vpThM2p1F9PQPg1hU3pM7tHzZTW8HiJr5CYd/krPD7h1M7
INgxUsBqYfLY/gmKgkRylU/0nXQmPMGMYcXULHZjmzxg4JGvnqWsEz/XDpKob6sF
hQsaKNNVsvJmkVwdikbeskZnnHznDFWHhxKVtH+3ngIp1mr6TSatlo7qHFRTx7mY
QMqDJeu747i9dHUh+KnI9f8hH8cF0csMdztoX8dU6yPZyv2Cw1e1g7OrCfKBuLKL
i5FE1gF1MDDJqRKkKtVkIgiPychHfLDqfEtcMRypyp1s83/nCfMMuzCzHzQ60FCj
rMCoecZXWRbotQGvXDPMDCU24aVgeHdulum0vVbntYrKG8ng/hMwSpcaW4a9hZiZ
YyFu/THTO+ayifGi+0PYRyIM0W3G9EN6XUl4ubRwpx1VPvrJJwsFoE2ArTjLdYQH
ZcPm1ynCcYWj+bT+HivwD1xO78ZaEh5c70idw5DPYbph9d2JnP3qY65HxY5i/p11
c0oIGNzMggmxuy2HYUAjVBnuSexPOjuzQfslrAn+revken2OyFD7vcvhNTmncdkv
H10qr+OGzn3nqqs8K2/HLPi0I3of8IFXupkn7dyzj3kbq3PFj3L4CTIJ8sMgQXK/
bb3pK7MxDjSMT/d6tfw7FDxx7rY0tAWncm+23YNdBsBlxYCBNE+oP1hALFLHKMI+
6zNo7+YvZ9JalGE18TO2sj+FbTge4sZjL5ITJRAuotHhC/+pd6u9Zex04pegmIdi
KndByPEI5hbinbmPWabtnXD88eLVHiDkKLNYGTETDrnL6D1uAGT33CKrZN6k5O2Y
ltut0uukv01hs+0gB1xyoTIlkEn+wD0iI1AmZFZOuA8BO6rxuDiIWixaizbPi4fe
w31mDlJMGC+e1kYb60aqDxG7dvz+2MultdE0UUijU74GbAVN251YunBEurIHxfnK
Q63X54IeQ3ibcqRXSFoh1x+Jz/dJheMyvIGHXtfRmW7RLXSGD5dv6gV6Fndy4dzZ
ojkhA5ZyihSt7b3GohflxDK4+ckYNoBbN6kcv41f2Kf3u4pj7cG9cSVcAmXLnH0z
nFWJ8CTN7wCxxSrT8C7jEaiC3OZuee2UZ9CZ4/b5Z6PBKjjrWXHcZZj1Xl01ZUgj
Lfkp07jXs8NyvsVymX/uZemIiH3CVa5M/0ORZufNlFY3ob+OxxqofoFEnPs173G4
T34h7PHx47il2wFhamxKCrljV3FkXeEVF57hcVmb/muQPa1slV2oNbhhg81NZAkn
5CeG29Yr0Sqv+3W6Hp+EfzQOSK4WL65YkrZ+h9bjcMHlkfacSLeSIWipLPUpeLoz
MBBV5663lwor5L9QNSZoyr0YPhAx0qRjrjZ9SwUoIKnkXjhLnmedxOnrSHCX1A5O
IE6XMku6eCl41lLZ0l9utVfFJVyNHIM18hRBcxxqyZGkuiITaJ3+M5E6My2oYoD1
W5htWJZGGAOJLW+U2nNXg+jWG0bb4I5XQ+94fCNlKFyeotw2is9/Uw783KniuaQ3
dmsyc/CqUaEBUuxPE4HR/bDkx3saZiRd1vZeMy+AHZ5j3nh3GsR9isld4XnjpFHw
CtQYt2R9G8oWQz7hIKsFv0qMLp9/4F18dzMMFAXJM5qElqJx+9rAqMJA/1yRtOvb
tdkJwVn6Kh70FVxtdoqJU//OaqT+MvkjT2ZSSbIkVjq3E7skQ/7fXyUHzvdcpqL5
ePOfcELe7TYZGTZiK/lbWJIZdE70LQIfLnrwaoa6I/EkbSnPn1Wn5ZZ253CpWdgN
ExDqxtvxDp/k8+0xCbz0F7IDP7USYmp/Rb+OJDC3OlRecOHLc4bsxPtPZgwu7mbz
4wNLsIPVOx5jjg+74GShCenx2/akNK9lTvdsCkZiX0tGpbxIu9+8im1Fshb+lr+p
g8qqSg2pHeMkbugFPWMQyg1XnpUnQY885btVH2Ihw5L85tJxFb7OjLNfo+leanAe
PYEThp/YF4+PbOk4wP61Gb3NjGD+2zcTL8xPs9X3AjRdmiiiqvJC6pggY5TFpYxV
2Kw+RQ6ONcF9XsV8E1plbfXNxxxdZLFO57gC5F/wWDHJeGslW/3PXqbzu8zyRkAz
S9RkdKHq85yXbso0byciXq67m31+ojwXEnPUMFko6YjVHoV61qnMnEflqPkcstOs
+KeeytPepMlyjvR0ruWTEe8D4bfsI5pyUVUOQoJeLKsCQ1pzkaWlDuA96sGsRuNr
ixzJJkkFZOQx3dExbVbiYTOgShW/HJlnJDvOxfbM6UVuJ1BIrsFYJ4XNp8O7M0iP
283ttFh5wRzcw5rgEUmyPEArR6rcofVWj9rou17i1ahAHCMq6g3cVe/Pa3dFck84
e7jsBk9m0E1K2Q2RQ6bzLUew0uwHaotgoBFGmtQmPhbs00FczeBJJmpb5N8lwvtv
OslBph2NBXGqpKl1WyKP1Qb0Y30EKeGUQgQsXSsezPIjbOGhgcpAvdDAFD2lXPF7
xLkNxva/1LE4A9Yv4pLnJQxsbnijI+ckx0fYWCsAoq+68egpqTsyvM3S/X7tmJip
j1jAXNlfkO4xp7arlEFh+fTWc1n9yoeFbb+9ZOPN/G4dZZv+qcdA8DLgDUL1oBPo
hGa7GVZq+b3uGcFH7HPfdQOYdOHgGpj5p936TUG+2zogjStaGig4MpzUtAOTr/Sm
Pgvyw32EJdGh023HeOJ1Ea6cCNfHcg9+w/hgUspmxWJieVn4UVRBhIp/fDRJqbA/
c6zpw4nzSf4vxtcrEbp3W0EH1D1Udw9m4tkfSOzBMIo4+OqGPqcmU74rvuVaJNw3
3kNMGx/Eix3MufXgiq7kjHNjFqc4unLNGO8dMs0p6lNwxmLcB7Um2IASuN5zeqgD
2zir+4csP+tRBBVPMH5Tzy+/WIaOHdzStBmyKvgU1MhcmVvrxLagBkM5Je1eU1aR
71iV5u4Ts30q1Lt5iYPoKK+F9LEmv6kiRkmUuyHoys5JZg+ulNAmn5WtNxnHjRJt
8zYaBy0jP9uNfyr9pfDcBoNWlwLOS+M3EpdlF55YQr/TO3i896r10eGTe4fdg419
pZjuwLetq4APoZj213639/gVfjWqkZ3zzONgGCd0QnU9dgmmCyBCZXb1+QD+z/MP
V+NvVdIOkTwf1T4XLdJfQ7NBJaw2v4sTqrsIb+LHW2euN53mERb3dDdHPQDAuw03
78eqLpHv+zSGZUZ2r5O1sTb01HTHLKnZPmSM/agnqHKChbNGyvdpUDRIZEz7iH19
PYl7FpD+nnqGi7PwiCMM0JY9HF3BCu//UUvUnvUw0MrAYnYFp0wP/2i3ZUnhIoAI
V9QWA9xdc0xX0zERm9U+5Yg7f5D/bVbfavwpMxd6mmWiVjJf3b0TKA2UP3dy12j3
ytVAGesrIR8BR8aWGw7pil02k4KBZcRbl+KeutGeck4irwIYvW7NyVj5PRniIK+1
pxHu6GjIJ/A7TgR1IW2eh3NTk2ryWLa0xy0ZotCEBtrV02nlNGpiL4ObHlVw22Jh
63f8Z6g8SeLTMuXXECigz8um49nGOVAFIm/cGyfFPhjmak1sV97LmkYb5gCyNJIe
E0Ca/VIgVF7VDe8D3+3O7LqbPt6Bd5C/5oW0Eh53ghV4wj5hWvYpYpaOHDs19QWd
tRxPn/eanwwhGhFFc/3BLQW5dkS9vJZOGFmmPz9Bu5AmNd85lGHiGDmnXy8mtZPs
nnZaV5aNJXikm1vPmpKMwAPCld8ZOAUELWKr5hghcngfhEczlPF240orfZUsMKfe
N3D9T41VXPWqelL5/gINlrsHoUlBmhCBfGFRwtiplTNoeL7fsYS93E6kgCKKK7D4
BxmoxHOJgaRrNQXQwS45nxsNuGMmoxOFsBi3MtsRPnmQi5TLheiSLquC8ta39BKX
lnNWBZSPjGvq/Poh4VrrLHMtnhXRmtlFcNnx27CSWAVvvAiVKyUji7P/+P5bRU+y
YDzeUBtLam0ynJrDD4UsYZb853BI/APQyoG482DisQ32K6b/GNI1OvMDCg1+qqbT
Iv7xVds4xVNnYlv1esxd05Y400QOcSms6wDZrIO1gYGkPWUa6sqewBv98+xFa5Ep
M+IPAcY7uzphNN2aZXNR5BIjzjl+B53eNPTwCfL0anq5iUuo8ATGy4BMg6ljxYZ+
YQiRjJIdMIXjOAQf8dNvc0v3/57dNkw7QDPfRdxzzzfspm+hTVJH8bddMsCixe/7
5bjQ6jetAyxZPTrUtHKi8NrboRC+3zRXfR176xk8c8Hnn7U2mfCFLwxD1i+/McOd
P6JXE2UYgJPi9o8EieMu4lmLHf/EjcUfWV6BvTReePjGsRlRFP7QdhyOJUQMeo1e
zHcvuYM/o7n2JAbDWgxx/ZyjKWiGB+RVzO0nQsIUJNyouERT6v47u9ab7c+kvGp2
6TEJwIOjGcekC1qyXifZXRppAXBcVRjutQmcvubrXVKAZP3T6ndoioGTHMLiGvUv
0xqZzZR0RnsfJ1KFvapyMghUJHlSCIopDjV7dhd5nF30uIgf4x0ELQb40yS+LjBZ
wULN5C9uFQHh0Pn35VNBBJ53x5PAHUTh4yDRv1g3tXnu4IZVyUuA9/MVfiSWobdC
xuxxHXmTf6zR0ECbLUNTbXO3cDRW30GhJ90B9INSSOc9G3nHoou3deglctJV4c6F
BDhCnyRFmBnkbU4FSwi7xIO1cbuR6RwIW1Igh1+BTHCK2kVxmfFvr2PTh+l9UpPy
/LMKYCYXriv8Tjcz7+8gSVmA29r6/ZdCJktEjQd5BjWVBmiI2rbQviDkoifu8aDa
g8JVe9ayLU9CseJDQjKGn8QbZ+ZA4teX6+st2WW6qF2iIHcQxiFdS+5uZ/EAIvuX
oKvNT91NH/BnmyoyJ1RkNvovinJhXk4a2r4pAx0En/J/Z7kxfXx0LK73CFcE7TlU
GvNLng3HMI5zb8DhRRvfNbVN/sv2VWwKmqXdL8DgGr8W4eG6ISqW+yeRVtRAq8hp
n9LRNlm88UxdmdQ8YTWuxXRpRD9JLutp3Wf8E3sEUfo2KM7byyJaGHiXKVN8bYz5
93bVmZSEUuFAegA6FwM7wPiqubSyO8jLrKJRFFcds9Mp41Gg96BBjp6ctqd6H+Xa
jDF/dD3GX6Df56nlAzG3zW8wCD16mVGckbzgPn429BPSwDuCdQbuvI0YLwdqeBbf
9E6ZKkw5i5+sAe6UNSANtXUcIP/bU/EItoJZlpYplbtnv6BqKtnWHgzIfpbXswFO
PZIOtsytaZsROzuLC8K4c48pTgL2a4lI0peowZExFRkvJamNf5xEChPo0n3lx8wa
knC2qwl6LnhRUsAnnyTE2RP3g8mKLHgz6whSvzv3mCi2qGbgT0LQOQaSZQratNo3
FQvYTxzrfbbPNFosFMZY/gy5Rt7naANl3f+bciZvglfAopg8zq9G3S+ZaVEcRXiH
c5u91oa+QkhwnkLb71nIVm7FirV8mTHTv7A90U/m8ku//kQwPgKcRAFdIGAZm6NL
CX+G15OZW6wDy8NtJjUpcj24AtFKOvYw/exavQt9FLf4AbB3s9uFZLYsuMNLG3sM
/vac9DL574EpUuB2WEwPq3oU7HTNp3/8yVbIupmE6FOnk6uv/XveZRd4DEPaeaBz
kkKW9KUWoilA5n576HZc3g0Htr7y6b3DITwkb4c6D4TMWT45X3iGxVfdGY76lOe6
PeKe+eK5RvA0DlDIjVMwaXiTN/MO/BKNl5iAOKsvYkp8mIz04YArYbLWg3ZF36XO
H80CQ5UWNXMUOJ+v/mTmcazHzZ97mp/Nzj2kTL0HTOGPm4TX3h1V+kaLwIRa6qkn
2oxLe3EEP9wNsY6FIrF0dUBpxqJuAziyG0mNd5/0dngLf77PbtPXNLl/T2zl7Iq0
O1SFESl1KgafN+7nbN+sRSe8Cp3lvqm7SNUOgNpAgm9MZxij+5HnIRthxSGC4Qkd
Rvia/ESD38814pQc+/FSzCLMyjb97TyTED6/T8zTK+DwcEViBNWDxQFu8Iim8Oby
taQXkwTPiSVM3M26MXf02WvTrDIKyZQgddmqIGI1hFz2wmh3pLklc2Xao61c+JaL
KJRme4Fe1PcIduaA+Q7EpdAN5colvD/lEA0I9UqGZBHjy70hPspuRj+T0xWbk4Yb
boS1LYjI6oBzegz/2aQYyC/K/tqoQTAS8EgbDdvzsnlROeKF2Up8pD7aRXNdWxb/
0EiVx/fYxxAJVv1z5BnkK3lqcVrzPqH3JcxkrqKAUWFg3Udz2Ofgka4qPapo0czL
+UMkBN2V0mwv+dWz4Bmt2sM1iZhpvtZpcEkDsZ1sZDHaCJ+TlDUy0ZRtSngXecMD
wGDcNU4F+4gLaDFwVqVLkwkzmESGIEgM/3HUjUQvioGwjrhX6tVPZ+d/iHOLw/71
/gwBXx9mNUrBaOWwh9HMlmS0ox59qHWRY5rrbrEu4bnf7cn1xw8JhFQQsVVJ6w3j
28gmepBV/ruQZEeCC7ThjVr0yCuXwVGv6vORoYdUEsVyti4PzLgQDl7SYPAgY/Rz
f9Wt0Tx+/aHv+VymZp5fz9/Ahs5RZquWYgGZ+/itTXTN1dQQ8aDI7wO06EIohfZ7
fiz6TqjFjqBxQFnz/r1VM89/WVcTlxqTCYGJGLcFsf9j/MJo7MWgd0xrkqrKSXA7
OHzIpUSt0F0KQ9TYMymrx3wcVAZQ3NobRxGOwYRQRClOZOWc1SoaGKpfbR1466KT
Vg4jA+2i3a2D87XgdxfYfSuHL+YpPbiLOlu8+TyRsPvnMOqObkByPB3hG7dvMGpY
VCZggc7xrvl5rOGhfg+G4tQz3x1EiWQsr9eyl15fP96FebzYE2Xp8BeLWFFqrNtM
FkI8zSjMU4xUUDXXPtOnalRSYtjDiGxwqui4fXBt0Rzn4x0bB5dM9JqnYTnvUSQP
twpjLV5ZksMHSDCqx7jFKxojZSMccbpi6/KMUsKlZrZXgE0I2cS6qmwhwu2i023B
geB/P4xcXiKM2sDimm4u55u6N6mh7iCxzahUYjMOJ4RAR0pH7TIig5ZpXDCPXPyc
IhXdppq42AQQEsZL9e1RPItX0NxUyuVTUKJDIY+Sau6Sx3KLDRB7NkbF/F9Kb/Lm
TL+TQo8DJSICOktC1nIy06PJBWzZPia3ZHUHXMasLwBc65aRI6Olbjh7L8LIdty+
f3CgI1tfpwIbMCQ3Kh5qdI1sd2VwxEZH/e7/a/lLEV8bbm+TnL0nuQoO7k2hx5Kn
g6G7wM8yQuyaKBOuVEBXodvSp4ucaPNhHWZw8llqj79uZdsM901l7NsWyC2mh+wr
2Qc3BtqPgwlop0lLMh7VLsCl8ZmcCSNoNtpozEMVc/uUvUiVeMVEuTJtvtEE8YjT
PEUQxzokq6Mo6zZGX1DY+0LG/sNXg83nGapsifIqGaMy+ZeWHcuI8JwDAjGbdi3d
NthiSaapPkRZVIjSmaHgSd1PDx3cuHOcTTfdbQuIa8RA1Lm//uQjKtYfs+SdJHRy
lMN9GADalodXSLJyXsw0PCgoIlSjQGptatEfaILikRVMd+T1S+2h2PmqLO6lm7yX
ZEbOvyfm18kuN3/m3l1fsQQSqxs4tRG/dQNMXaV/v4c/spU3QTcpyTvxB44W1MOm
iT0WMiNYYpRCWoMSeiDnyBrEicd2T+CdnB/8KEkjDCunjzzpuGiEYk3CWif/n8sP
dxWBK24Z9tgmyzewLbPO2N2YasjgF7fU0q5A0PEOMA+f4zxoZ9T6ygA91ZcLlSNz
Oufznp5YuPZF5EoIH0QIikDXY/yc/njM3wtzUT15e4+Dvvpfu330jRPWKHfrSvkN
+qSql6TtFtQeSQBYfdTl7WDO5Vbppc9eCz+7BBc1vMk8/7oiHZTiMrEIDygt8L1y
D8lfXDlVCXwigdbw+1g2iBQpiM60P3S6PThGI839bvPIaq9mjRLXJPmlDH4F0Wh/
3lXuSo38CyxGsO07S3FJ2YQOTI118G5mzPGv+fXDl98nthRJlZur4gi/aT3a5Zgl
j02KFtJQZB7uDlF0cJf81iZyQ5AZRUeM9W7ekBMV4XxLsfSceWDDQyGLeSIpFh5n
tIDc3aE/EaEZPzivranxxZg4MuAXUgXpzjW288s7oxcE8cco3g7s/q0ZXLL3KsWF
2CEGxCjhr5WycCuFLUxUxcmtiGHbg2+r/iftrnBHJhedH7jWUlDjTyu+5cCPP7MO
MM/Qne5UJZhQphqckzr3Jl2BIwAE3PqmtZYHS4hHSlJxCUHanB+GD0kX8GpWZ85h
NChfis+D6hN+9kms/uZZP4MH/D422j4ViUAPIRqruLv5gnikLeWxC7rGKPmQugZv
GuxAE7/CyIPlbOb+MjJ3YqKiVVx2pqSx1wHuAryJzypBOAqtDMxZTqB/uZM27B6A
EMjwlKpr+0EReYJ4+hpEfVFy0C0DmpDFuNc4BQIWN5uziVv6FndX2/Y7yZL5ag1C
3MeBCkZDe2BUIOlNEvkeSNiIZx6Rfw5kATeXoLTmtseANaQfQ8pLkH6GvlUGutnG
X/TOWt+eriBHBQI7woa7NavAl2lABvJLLcdzUrff06ryNz4mPUEsAikjAus/pRmK
GFxXbAlOwggLuRejh1tCxySsJ8J4Qy8L5RfP0gZWHgG822Pn2sX1aie5TBQekNH7
BQIrS4c7O94yMc/u+TjoaP784WRNXt88EILd5Q7oyzEHcH0rzhbi4+QBETtjlDCn
1EN0f5q9mt4ngHc3tNhpAecsG3hQQEYFeS7YETdHxvfCMONnxf/0cAVb2syaFdXz
KdDEJ0Sl9dLjcsb7DjCKX4FF2U07brEhVw2fJHI8n9PBastN9LkAWW0HqViu9R9M
gl0CCwbPZbuy+GK1TFFsIPF6Yws3ZDEqAdQqTEi8SyxEOn8q3NykVHTG18vsMVef
7yrtqNiii+uOwE9V28YGycY8PVRuV47NgPszUjcxWdc+pPHDP9vbi7qUILnqGxLT
VY/3rgnEN2R4KWjVgDJuIpL8Eouf+SMn2YRZYqOlanTrXA+/svm3eBrCF04A9zI0
c4uOBCvqZgtT6oPcum8v+Ge0yMlmjMxh7XwEiB8zqmx+o/vJT0lACQmwMeQmnt9e
PbSacpB+u5NDizam3ipyj6ps6gH48hO4x0/+zLdVdb4L7lag9cf4YRYJC1PzmUN6
fRdYr7s/G0bb5J44CDGxUGqr48/d4Mc2a6u7bvOFR4sUEJILy8qIC+DCtAixWvJX
6XO+tBCJCYr2PwfisovGC6eYT9imSFUIzhSudu8kq92/BuIaonglNJ0q5BzqljJT
UHeEpKMYCfn4uU66lwaOncxGjyfEdH/pOmvrqFq+xChA1fv71vqBjUVwE7dZga9c
WToXSZ+WnyXqo1vnjO5SHQrzbnPM13m8XhtDJcrVkoSlX4aUn2gpmRcH4AXvLzwl
c4XRi4+peMbRjYbmd10kmZaJ8hw05LdpJpTKf57ivDKMWR/x/WQ243xvNVOHrfCW
8/J8bqptNKnMD4w+GB+KSgkBiuQVBzc/NmIA72mQfzd45lAMz38YEsjI9r5dUp7l
jgH+7RM5Xc/bOhkZ+rf80YaAnCxkzIOFFmYfbDAy2RvC/GG8phyZcQNCGjkvRVLT
MuFMl5ubm6qMDJeq+V4Zdymu1VQoI//0YKnUgqW9SX+9uFDlyxpyZTr4yEzVZW1M
gFYW4TitHMvo6NGFRJ4SS2sph5tHD94kaJPrGQjylXAUPCoj7QH4JdhHvgYgqjfB
gk6SU7xvQsDCMFmzYHZUOLILk7NwXOk3LR8ghHhOYSkmaaTTV14hSHWCQSfnLJSX
2rkoK19qwKK7FMkt3GIEt66uE0i7y6CQTXXNJDwMGgzi9aX3txDwNpjFaIOMA2Al
K1fZM3iSFeAq4nJwlDn0Glt04te3Abn44iJJuPpi58CN18YBp0djQbn45JQ1pWni
JUifRQeRlI0R2XCkXC28uTJILUCkG+j3DrznaGtbNGf0qncq3bUmGc/w5kUSRY1v
He6M+V/xgME6UmRZWf2Fbn5+7zIuGF6OhbSm5MF+0TE8iNEKshQ9ehrnfVMes8lj
5vcf4whJW8iPklNtRiANQCzIvwishmPVFdP0TFqvQsec1yDxiiRpQsO/88RCWOeq
eni5ySyeBwYvYB5Jkm4DCdTQWoxNEznYHXGZDl+U0NsCSLB1+QvPPK7o8WEfIAY4
ijH79IV3WCdxunLUeGMmGWGGZuCO/epU775dnLBH80zD8YDW2GF7p0uejQBI5sJI
ejY6i3Q9M46luKmvbgIleBvHZNLCaA6Idz1IziDemjElshpZF4f0oZ3sOhfP1urQ
VlAYiEsdZ5DDXEb3/BLkr1msyRX15mhw6SxGKWPWQvfdzhUKOsXtEvJQ/JIADbeS
Voiy2g9uzWy92yQLEYyVVePlxIr5OyxhZ/VZCmK1UG9b/zM0WxqTQMtbvXx4nPPU
oFcyliWJ9J7Pl7PadXuU0cm400MWT0Ht8bEl7jVvI7aNuJEWyzOJ4JGCTMLyaO46
1qY1DnHc2VM+YCZLbkm+5qIHHTM6vRchi1z5pUmELBXtuKxbk1rLo6xlyxSSyYuM
Eiay8Po7yTnB3y2cbTS/pDfwM1jxUpuWrEa+85V9LtOiJUegxAYnSRySTynkNgKv
+QT+e3yzWLgIIGJGDP8OiAFhrtFn7xuw5WsDoEEXCmgXBf2xkKJKPwEtj6KNsByF
LGa9JDC6dWoAIVumTz1dgmozDzVdtLDvnKAcJHUs4df5HA2U1JNVqvtZTKLZGU+r
0ghjjtxe2KCYOUM1VisWgzaqKjck4HX+CUZPNrzVBt3fZaSUrAdlg9P02YVwUmA8
J19GPGtB1Kd5sFCh/ZTlSl6mSa77sBZXQjS0DLW2oH44v8zpIuVxTY2DDo0Rc3V+
UVJnxOGlEmOXrIlmLMavNMzXIGp5gSD1GOMnJZYAdcr1I3J2w0N3D9DSS7U9Matq
7nR0TsTtKln3BMMFmnHM1R/BeczGDsCTVxcHwiaoaOBRNstXGLLXsZye/uSpP1Ec
TqkceuLv6sf7Ni8AzTqal3p1seeXVd1j9RAlH7pwlcNDp5eIagnjGsg0cBt5NnW4
bxg+RmLxqiLJBjnlVH1nXhrfMJ85KNl0+t/dn02xHhaCy/nTf95j5rVxbs+tNOJN
9bcIFHaFo0AaTxPZBAty5FYp8IZjH5HLObefKoHOKUaBwUF9prHBMTsxmcTmxqd9
ZLCMA/RVU+GjbdtDPfalv6+ebB4UnTFgtYx99gLlisR3VgtdrYTFxaTaLNXXQ3+Z
OBQ3TBWSPPPrG8chkrOP/60uuN4dWJGTOOq1ecHNUjIPGDAE8pLdXSWR0i12qWjp
IF/lh+g6j3Cr3TSpiJLQ0Fwbjwi+ItRMXFNLGTrND7TUY6mENXaT6syv0RFqLq99
VJ/leUFaOZRre/Lr4q8Db6tQZosvdbtj6Wi1RoiyRvvrrW1xBV8K77jp39FG9Lpk
y47RDycmVDY18rUyUItC3YmgQFDrUZnBF+wm974eyN7Pm1tcU6oMfIzDPQTcjL7D
FpSAW8E0UTXw2X01K4GDhNGhFLyGzhdVEOWjZm6MWWRYPezEmn+ghh+i+4IZputN
K9+2kilZkeiS/w9r6Des6FXtZJgephJ3QEcDnGX/bM93SfBD1fZYz8aRRBOpPXkw
O9ynrUVz7edcEehlN2950rCqNu/z/G7/Xv+indeAXGMA2pXfdW55A8Rluhhm7sVf
1adUwvZXB1YK6hRI/L1fLE3oS/7HxU6JVyricGiRFRyTbSxNnA4rY5sCCK9/Jgb0
xXjrSSFWHJF+i9KnYoHUFDa4DsbIb6mFEevCdJweQtUuKmrIczjQiGSkgCrP3WSw
YEAxi4siLowXBdnku5KyBmrsZDjslm1U+xDmLbbUZbu48aII/y2Op5MklPwV/VeC
FM90v5N6GYDMT9ccNpFzdOkmVeJ79SJB8+iI08TAbmDzkKqIcMqonqPOdQGswTMA
JJ4I+wa28IXVBxAbQG7KEBZmHFL74fAxeLIDlQaCPHK9DzSHUWi9NRXagWdhrHpa
Sh9spzGZMmhGC0xHLmRGQ2Enq/8LTGhM5HjQmHZFl+Q4zWPpD9iaIMT7gjj1bYIE
SLfPxNxGqh3tkrUzEVdiESaPmlNWehTCI6aTqKp/l6QtOI1NFRgWE4NCaO43YNic
jzl8dq4JG4FvnX44bfk7GnguEb6ENDbNQJKGYEJNFE6CrVFUq2x+Rf0yf6QZMgKY
+l8TUQOTEWxg+7R4GTXGIjL/WVDonESFzx1/NkC/M4RgXS70Pdfnal4pWpboev5B
8RUxyWLAFZqtKUfBRSB3n37mjoi2aA2LoorQSVa+to5n4qU8d8FKquHR3Qo4H92v
oKcmE1Vzs8Dw6BWv8W4fEMLNbRuqyqATaiZUaqn5UtqeR5O5fQW9jRn9tErXFwR4
7wp4xjAbzqRZFh/ePf+7ZkrIsJw2NwPKHRoo6OVvRTtXMfBDK/OZpC2/5hreR2ox
GBxVy2vHty0GQ5IkvBNHXOBIQeMkHaCGPSX9X7f9zfXl5/9EpRLN36I4HfKzDe7H
n477NzIdEGe955T1oefBlSWeSBFhwl7DrMhkP/eSXI/vyYsQFRrUiVSm0p/pIlf4
el4Vgqkyl7Jw0MRzSTl+M1Peq96iRp8elm6cz8jQgZugiNtV7+ffXWQ57KvsjCkW
ZRDz9onNiKin1YzhA1oC9+8LWYw5g6/2G4Z2qV5XnPOUD6/IegWPcRSzwgGo4vch
dLodN0xVVdtBG7eXv9155a1n0c6n+rWN0ryVxcNolDGYJEsH1Ctz/YelGFlAjuwg
YXq81pRhb7lL3sHZQesgI7/Wx80nCUKPaswFMAV8NenD+rIIIq6jSeqNL0OXo5TM
Vh7ARTY5aY++NRTfvd099J2jmVwiQX3zlYk61K8D4SrYb9l5Ry+qUT9ULhFtpRf7
t7dlj8MYYe4ThEAYNTw7ltKkvtfhAd87UIuB8deENvnNUxAThZ2da7xxpO6v0PLS
73xdNAZNm9nPpPbDL8H864X+GDaWVTUY5PaVXYR+i9jkDRM5pDgRl/Mk5ncjRafV
vgbnnyisFHonVNXIVSPdcct3oQFwmVSW2yE3p92n5iBmznga/3/FxJY2sV+SL/vf
n3IHa/Qy7lLp37VvamdIGttxWIYDMuOSUayF8kBArFCWBhZl5a6xk5iG8Vf+2hXc
zDZclHgygPfUUe9f5rhTe6szQ3SwVK1we/Hp+4o7Jm8tQTTdLyyu5B25/Eb7HZYX
coS0fJnw7+iva4fgQ40Ujp6yHLJJp05L1tV+ls4KGW/vDpd1hWK4wfTwKH7g3dsf
7akq1bb83/D+5peMPOcgK2edwrBhHSL/Y4csF1LAs09jEt9Tb9tFPbhkZVW6vDF6
bBDuQKw//LsTFrWoJUhkHqNd0ZOpdiDL+DGv3o7knKA8ahArDY46WnJf1HLfdUEc
xq3QKukc00ANpr75IrUUmdXbojFBa265JNLTVxSi2i+cqW0QJs0URRg3iIW4FUDh
Dkn3ZO9sZ+P7RA4PcyFNyPzoobmjsaMIKuGR0sVa86579e9cLjnZzSWuXMsoLGiQ
qrIc/u7szjYou/qsk+mmo7FWARPF7NiSD3OH3G6JoKv3PoZoI9VlTpmT58Mr1UaI
s89wEjpkYzXZn5zZ6b0uVcan8mcSkrTTqLOV6Tu7QN+zwjHDlzsqGaRLGV5IrPiY
nBpbs7k7qySIbIYJvpgviCz2nRBcnnwLU0IErUDoT4fjbyzacId3XkXatVEuu2CJ
zgxN9J+3qqZi4yocjfSOYH03To1dW3ZciY9CB3Z82Amrh1GygoFYc3feMAbDZSoZ
4pW4zqdd5pwZN9fM+QgM7xolDFSGmAYpZCB8rbSSS1Pvv6CNYRFIz3OrMXF+CL2Q
6YllBp4TTQGGNB8Qr/OJuYhiaEomXYIjAVXods8J8Ard90KK8gbiAV8URY9A5/Bd
HuPKoVf+Oex8mEzXdtXnwh78xaSrxWFBAFdtXs0oLz2GyrP/Swn7ViJM6crEI7Cu
TzMtJjLZhXrsYsXsvqWCkRkFy0EgWYgCEIUsZoh6CKvAXQki6/HcCpjA5Iupvh/N
0iSfsgrWperZ1edegOXo7URR0QojiqdURGWBKUhim+M+El9SwGY8EF/0PqN/y7b8
Il7xrPeH3WHb0FpQxWWBNSBYaZ0AWaTWpE523L6z+vKmdpVDrdMe/e8UGTrDFusH
CWRD+91Pr2AYjxYNw5/l5NkID81xHZFBafJuEmjBjw8BGYiJ065diTh3HUDgut76
5WakZb2VyFx3a2ND/LNJOsrb7mizUf+46OurIZmVKUWaV0whkNMDZSkOBqIQ/7fF
Ox+VXpyYs0XZwaSXOtbsp5VnnMLRx7KV+YSQ9lKwSy6XH1zclm83oa6VOp+piBaO
RFhZuLUxvgxP8LqAVZGfCLCeKj5Fw5ZPbYs8pk0DBwLE2E3NUJEWwE32vvg6+Jjy
kawf+v1j2N7F+PJQfgc+UUAw4pWoVV24RfYZyrl6efVY6g+9B0j2bel1Qm2oL2ev
Cv7TD0VyblSZjJWuCngCHDdu8QPjxCsjW4Zc6P93igQJX3ErNHnln9Bk5vqu2Wcg
y97ouqoOO+QvhzJe7DgOkqAiagnrRnaF8SZSguwJ5Pb1cE1R7Emy8/KuQiyjQ3+M
YuQQZcOOsAyGIjrFocWprOzOFIa/8nkaBM5d1kjnp2FKaIdR+RW3mPw78MTQITHy
GE4m24NJYxVvIszbUKFeyzDxGktYzkOLVovhbtPsNQGOs+dvhYLv7DXnn7WoKL01
NESC/So1czIjeD1I62unajeTCYpSbKVYH7YnKHodO/hjmUsu0WAJUBoY8644bZol
o2C/M6+RnnfhAu1WEQn2ijKVVQf5Ula59irknCqqwv6q+etgkaAJMOGjTq/fVDiR
yQc4zPfzWXbafdaZX2LejR3hB2GhWOY2r2iZxJDJf55QBpYHgmsIWmQl8MW8xisJ
aSaWR5n9U6ScySGC1zO8Ehhq2U1C7mdAjDMtF74ngf8rij/NBfnChELI1mhQQNkf
RQN/Bn5gT36qVdE8iR/2jSlsq5Rp88AMyV4qSnTNYUyy11UBLccfAS/HHSlJ0OUs
4uTL5GkzBQgLOhsYdlEUZVMEQoMuBtudBtlEwTb1mbKqdr9+iteXd80Qlz+knApR
4unmmLGpSoTB1R7PDYBEBF85xiac4xhJ+DI7ygO01/oal7IoGKfbShI2Aj4IapQD
rtqQwBhdaQDNYRsL7CVCqup/KFvTExSu/H0ashTx+0O9c4cGAWr8c/Wn9TG5nZKP
UGAW/mdEVze7Gng3pPIvRo4slo+fxmNb5j586/vHLLahvV/XZ5jjS/dzVcd/1g3a
UkB4QFejToU/AlL/qURHEyuwKkx+IwbXY3I7mN4uUbc31qhk04w0gIFsdv1DmuCh
BDAjdhonXoRMmdhS/iwBV6fZza1Pn9nUUjIlRAwy/fL2wbsaq5wktpFhEh5jU9+l
U15yMbjuezfM17qh2BQSWLD1TkyFzVfGvn9ZYnWYe+J6m8iPCYzhWzadUbqt7bd+
/606fP4XskHHdjfewafgjByF7y+hbZZriNzABdQCX2uqqsNZtB6L5TVrvMCUPGyS
3Z/hNEKKRxzK5XfZOXuHohoSrPFAf/I1x5/Wn/n3OrSTIAWezvwRz8mDPmdnsaqw
fhz/ZWmWt92E4gxiWn6kjKpfbhQGloseode+j1Zo5tvIf/Lrv2KGpz17I9UYUa5K
Wi2xks0pBBcnFr6+zr6CL19opyWnpJhrLYGcWZf+jIhUDaJ5IXxq/rnsGqtg/mqa
XY+03NNWgunIBBGBSssu8oJ2lxvk2+QxT7HhpittWPaVuiAHp7UEeXx8E7n8GK19
b6DcXAWZ1bi3+3MmEzcrKfMrbMkU4WQ+zRDGa359ZUXQYlgYco0n4CrGh0d2us5q
BVlx1LD7GdJg7J/EK0oe5EOcnDUvwWr1sj4uRl44VVTZoenNx4mYWJVVgtm45WM5
5hkkZs1CTNWWQdROk1+zr7GkA8ZzX2xHOV1bCGVAqWvWScwjhX047OhxTmrDvaAQ
NjWYs0PuX6GAF39KWQtV4gp6+cDMUbrvLrdope5rGGvXElOuRt127xomDQGdtubd
tnfE6cvI1DSroN2iJFEFiLVYP1gASpr6gGcbEY2fCh0YK6hOX1Qc0VOKGH/f8ZxB
n8kjEuzj7Oi1a1V4n10Faq3xXO1BsR/JaeJUTySwuA0PoIhY56PVwunFLk0/t0wu
Y0fwoVWOAs0TwlaEg4562C+OOsS3xyO3UqVWo7WL9+7aHLx+8Ro4mjC6R0FWdhZv
00t6z3kQMiCGnMAlff657GgDtpeOyo1wibIsEeh4w2mGaev1z4gZHOg+6Lfdu/Eo
Pe9XDxulJDjaLOA6kwAdlc7TdfCSSRBi4LgqmtvoIzSmdHPJCTWSUhZC6GdG049q
zowm/3ZJK943jlJf0BkVgqk9ka5gXTY2xhvJnMedXnsJAGtjzckOjQ2bbuLqiK0Z
mjzqPfZBR2xW2231vSAMMpEfova752YyghWKDLhTJGfKHVpkR6N+iChvLL9M9bXP
XW6McGC82d43zxllk9eE+GGBt1G8zug3W2Vb6EcApt5UYNgWGWDyxy3bclE8P35k
3EFmb02PAZFnTpDMdIVPickdaDoYX/6024i3fPw9K/dISS59hAqnQQSBP2hsKyWH
WW61G6nIraWx7pfx3WRyOTI2zQsRfZXxFXBZdeFS3YdJKVg7KpwmYlVkeKrgyi23
IE4Io8yzOjMfOi3RLKb1qLi9d/iEvqcnpejAPcY1zoQeRxv3TxHsWjEotZIUnzAh
ovdZQVIFBybo9fbjL1g02OuzzfZEzyV1wK2Sd6al0CXTAykcUr4OJfNmmT/xjWCb
ewZ2Z1dDoijpnaxZ4A5DKveMZ+4RX1T19rWvlR8h/q1xLxb0eSbyzn9vTnS3qmPj
hRsGk1+ZL1bKim+VP/EP4cJIIi/7lNf0K8R+BqVs9CnclXOSa8XmCLc3AVL1GCHJ
HD7M8wQdaiIrsa30F3K46hgcJQY4ld3Ns4XQnFrQoNCQu4bDgu7q+3wX8TW2E59V
hjEU/zTJjWT7NqU772jVSZqrCDg6cJcC2f3thDFN7ccoMQJJAiKSf3HqWSmTrCGZ
ve7lPIxSvlFs828X88IDXOSvfYeRsH2ksZ7M7aDqswwfkquuLLCb10kPi6zD0kNC
SyfVWJ1PldSNPt4mOUfx8wVCx5OFPq2fjBkK2fiu86aUzJx4ff9WU59ddWzyM0tD
727QDu31ZYJ0x4IxbKwO/8xvjL3Yt/kR0bqENXhUddWR13w5qlmyWBbYd0Hke0ms
aUFHfaL2IqVkaWcDvu3imuosvEgotDcAa3WQkcZklaReO6VdoNV1w9A0cmvEo+3J
s157GsA3A4twB1lIjjE8TA1X3poINtPZYMhTigfGmqBIrlIEyaz9XalNHGbuQzuv
ADQQR933dF/6qo8SKg4bdgGo6B119s9QUTwYjk6njpriGnjQiosEmAx+qeHWIsNe
MOsjwR08cv/eCPCNlXQcXjpurtXiW0Oa3a+L4e/P8+y4tQBFooMRSKyFh4S/GDrl
vZEHYGLQ/i2u1fdCymjc0jmkhUAYC5BB7vnuWDV0nuHglp17PZgfJk+Mq9hwKLbp
FVOX0/BVEnKQ/AxyGlLySAy1dvrhEhBr/99O9/9Sg3O9cmtC5gVy/ORWrExxVIIk
A20BibdlfdiRqHMIcmDT9Nwdf4jB4y9q/ooap8e0viJjCLMPkrrdD/k0gvLcwEqD
HE1eonusKbdQdo3btArwPtrSjmEu6Wqjtv0pTjTiTLv2rPoPEqJ+mzFv9KK65Vnh
f2tWMeb80Y/SQn/2dv/ZJC4KVMvVwVNNVayUSlYavBL1txo3x7L94WYE44+PdWRF
7cWRpYdHUKd5PJk9i4yEFmsCKc2JLVJvyVmL/DkFfke4WR/lOydK5/C8NmES7uN/
Zci8D6cNwWs8miDL83pgHnlVCnwi/x1QtMOztGpyJ3FKKn3kvMMi6dV5XvLCBB+r
hjbSktrkk+mQ8Q6UCDKgwusXB/M580ZFJxMh0iDT5oBK+yyJCjqOxw8+rFafL5Aa
UpEoQuWbi703dhhX0CVoLFHwiuUDKsXV5w6m8JgrFl3jBWpGjTLsqM+ycFjDhLYC
5FLc5HgnK5IZTQaf6AZyQL2kWIcXXgc/Ax44/2VAG5N190+uMqT6W5mkBHrbgO9s
NzPRAqaO20VaNKDu1ec0d8Ld3LdZ3LoKB2m4hhFzrqazho3uc88n1Gg8H5DyYux0
3dB11UzBflwICKkRf+l52HNHCKMW9C1KkBI4TTyr3dcBhjWQldfXyeQfYjcpLyxJ
YzVmSHq24zgoZuQZSSJBrnCprNIKcjzh2so2TzwMSWaQa987nxFdVjlezp76zv1c
VO+MFRPxKl3/ksSOcIyxCrTTVUHfAjl7WFQO7LdHtnPe+smGImu+BnnUupkFbLka
aWaj1JYOw0iV40Cf2dpEdDprYPLl6fUJX1iPIkZW9EMyH3S+Qx+GRH4qYrGOE/LW
qeUV1g1/g/dM+vtm+1pkXoPxfuvUvrPvBgoLJDQfKVEtlmXzwgcW05rxevi8Naa4
9gJi1tYMDoYeHWUAk6TxNrgLQpAm+CX3ocC6wppq321Z0+Kvwf2llfEqB7HLdYr0
WZBckyj2XG6HE3wDQ34X1VDZVQxWvT9Du2hnY8kjBUM3rU/KkUyv4g2B65P/CLbk
hc8uOXqa93MSjHHGkBbnD7COr6gMp2tmVlNyPTy8yBEPWiIU10rlj2z0MVI7CfUX
ZdJgH8i0gSjpA/0dn3SKIyDBKEQCYJ2MkuvZ7Ki6DNcbSF27AGUbXDLDMmgzGMgg
SAcGM1UXaspMeTRHK7rUt2RW/g9rz/cZsu3Fp6fEEQJw4qYCvrXdDw2vK+c9e6gz
VsLhyjbUQTDDAhZZWbPQGpiCP1oRrgRd/7ovhbsek3VwOfa8TvZ3SWrvxf0ITu6v
Ric+5o1mjFtQet8On+p1H/w4kqg+l/kW2Qg97/qPSKNeaFKJUsV64V61xrPxaBhu
zLFV+rlxwraib9za5M8Uh4xbwz+qHUG/cwBK1YH3gb5/2yGM5wlOz+Ab7ukCmnbN
sFTRzGB/fYV7AYSsuIisSvhMFG2EXbaV7dAsddn5w3JH5E+OpNn3hl4pIiTBiVdk
MO294ivjBY3Y17IRsqGgEU2QcpfCjDikrG6UtT14ew0rbjcscJbvVfwcpnDx7ICL
ifVvqKV3YBbnunxPXCoiA8j4Ncj1hpA1Oq/80+6IWchwlPVZ4mjaEUBq3nlgqyKG
dfoxl7sHPunhuMnhO9jBXuqmQ75OwMsU0oqwtwWSynp0QPs0/MdD8EYWqd6S0OPS
Ih4Gh81DQkiD+CiBiC/WWCc2qstjurZnILg5N39hV1Kg6YhQcIeBkTDbwEBeas/x
WHZmGWSNunyGPsYkgsO1YDxcmaNVO+eh/qmm3WhsrzBHd2Wdub/xfsMMGgy19Kp+
SUaOCC1TYVFMKMAX2PyMkFasMnELxR8XJZT615fWPFeDTuEW3+FV//OkO8ULLavM
fBsjc4GXLuO98WUCh29DIt3caUy6ix8QUIeYIEKIx92nKqFZfo/U15+HMxSlKamc
XdbwYhOrKqteiC0EAIbkjW1oJ3aaNQfPz8e0QrDOLXfXCG/4GX+NaSGflY4l1Trt
XpL7s4Oqxm7WTQMvxJkuFAaYh8JcflubGg1r35OWLAT8WYY1slSz/Je4eLb2OiWZ
+p1JF+5SyO+pBTgqpRyRqp0eEYL4cEabxd5zTx1QLfy7hHybW/86kv/Xpo/eNWRN
U37GcVyYiApMXNGdlrkjie2DVMucOnJNyr0XvE59+9xt40ea+sz8F4go0s6iVI4M
fU2Ni/O5wt2V0oGTuWjlx0Zvr8VIKDmC53En8deSG/aJRHcU4zdAEUB3F0MVGE8O
+WUIs1R5aJPw839tyj9PA+UauuZBhg5chlp0i6hSo2kRhWiH5NEdiwBTuCQ3g8oW
Kx9vKqjmdRPoQavRQQBenJc6uSYtAkqBpae05az7VW5zqiw/H5YLtTrldl9ntlQl
m4DsM3l/4qWafF778Wk2Zxgztznx7vF787OMKTG7A0S47U7QPPcBLw01ANfWqmew
NHQAnNASIeLj3xVCOOn7r/scb4GRCFUEc1D2ssvUO70c0A2hsAcAJqsWjmqrOVSW
pNQVHGttx0uWBTKoY8w1bA6s0FhFT0QPCEo2pR2GAYtHOeETTUMQfGcGBtfsL7ox
R2yBr/4WuAOrrMajNo1Ws4UIPhM10nzYMpWyva2WLF3WfiWBVp3DWgF0/stmXEOF
Z4SM8i0Lk4I9VJWNFgJPUHkWFPqvVND28pmVitH0GNoYcQJYVD+hWE0s96/5u9aq
aC+gyOldo2VMGzY/Bunncyxte0f1wUEE5WuqwSQbqZvovcot4rJSr2zwF98TQfzH
PZF9+HvNRwZhNGyZ9P5ghms/WID6D1HNqqyQy5JGTcRXwrbspzP43dMkS/e6KakS
RoxMS8UfNEEI73UxgMOr4sY81t2Xw55Upoao/kgGUjZQ+AhfX3CGgl0kT79Xu/mu
z+Sc5JCeHWxSW55QBkjYgjjq8YhTuR1D1nM/sfOBd1JbZMxM+IhEBfF90gKCt/Xj
u92+qn06vv5cwFIW/KyNPDV7egTrL10Blm1tmya01dTv50N2XHX1ETbCewVbczmH
HXqaqLYVSCqR79QZYM+VrNhlH73UEdQr+Z240vj2FU2/Ux1HBtngjt57rKD1tifg
RUvoGd7IgtfWj7pzVmpL8+aH/SZdKJVIrUK9je32xaA0Ctv9zWKGI3C60pVRtB5h
rQpJoTm0DUmenTbecJUHX/GNSxfTNNuMzwvw6sH2jj0+5CEYe3WKXCvYpXd7zBzC
eO31QpPuGITHEzCFrvJrnTYI5e8kS/z58j7nFFVyZXowYX6qsNmJyvXevTq1Hzxv
ePVRSNQaUKHQx7jMqWgZrc3xH7lxzqMlWcLRyasFDARxgxmz35xGrCBnHKaGymVM
mERuE9MXof0utxnY01XX0UbpxgPo4uOgJwRJZVlJlYisYgFuyw1zSYD9fOwNRPBV
GHD9OhGXVsToDUhSho2kTO/PghS/mItE2K8BSgpsoohS/IW0Sg//3DOfO7xUjAJx
HaGsIJnqsF6qunB9MR7VrWJZnVHm0uYflU0aRewVTU55umcZAHxKEHGpEh3jAvjK
fTeBt8IzXj3NSwXYK8EfJs1t1/sBik3dhWK7KtZM1w8/4TGdUJiYlgSzABm2T63V
tmOTyLx3KSqmWQrNRom71o3hTcoF5LB+39gVdwtdcSokCOjmTdhMnI+hRtUMsYF3
0V3D/1vPYErTd9yqwwGc9bSrsd5Tqb/l+Sr0UTadm1u1+/TywmsrfX92g+k9bzsU
sZqvKEHnOt9nb9dC7u3nxz4KsM2yfKsKtBImQPxTeDJ5X/KWM3h0jsW3F3rF0Q3V
xW5S/DeN3t5TGYjUZkoSjdq8+DB/jhki7IzHt+88zsjeN9tR30NaX3yfc2x3G3kI
Av2i9Daxrm2D+pjGA2mMS2uiO1OzBDrm8VYjutyBOMbL2HMooFqjBiPwXpAU1kfR
tt/6+3p6Y6tSzi376xAyGzqP+vXCObKhd8DR3PLrOtgOWQuvEaH5L0nDYq0sdZRo
lvZ8XOuohsCTxnB1nEHZDJlld0JpTE5Zr6jR+GnI50z4xQdCxznDri6x+6BHz4Bu
keHkZFbh7Gr3gPsjY0FhhCdjCol8B3cVJIxMBDF3XU3BfN8miog3hZpB/x+99zQ3
vMyB6pTN2OeolQImihX4pwApafZQQfD81KrwOGHUGsF5ILfCbqvr6CGcUDAEW2Tu
q49S07RroTAkUhsqdsKoE+c91y7s1CWD0/lq4BbEZMXn16ymjyGOzEyc6tU7ERp2
6JimDfjXuazPDBIC93i1MM59dpHO5xM5opHECEwRzCNusA3Yaf91r/bcu6Cks9w+
S7FOhlenLLHZJZdLUWa4UGEdFT3N67AeBHoFwPXhU7H6mAjD7prs3W4HtnHiD2Af
fq0mlfqCHg1fzfa0cYqTs5SYm1baN3ZS9jBg5QwnotJKnU7YaN5Lyy3Swmx0DAeq
fkVJR7E5R8XlI5z6fiWKhiNF4+gX2e+oGHQhgpcd8vczkBShcW9ZVdBSsv60eW/N
JFB1+wPL0OGP6bnX2TLQnHp7FbMvJvjOrzpwyTWXQQG7ApxxN6JR6Gpmey7EDl8/
Mnt6Y9t43c0K7c4v1COTHX4yO/5FSVXEBfgB188TKyzmfa6kzEnwRy7hKN50DwEN
Byz4ALJtiblCa9qOEmanK5JDrqe2DVMeuOmRM8c1z2+J4q3L50CIs7ZukVGplyto
uwKxIEdOIZcmabi4ZiYA5G2wQLHCZ1zklw1CrwE8UKqHeQbycK2jPUYro4wogAZi
MejvuPl/hHYXjejd+X2Z4NFetrCo0XLq8wY5FArnEUUx793TrXYMkpSckucmESRH
RSz8FDwE3qxoPYDM5DFAxgqWp26P+TguenaTVN0a7BBgYxBmZGySpdla46dOZUcB
NWSFdOxYgA5bunskFLqiRn+1kIrDUWyD/feKlNHJnKXtEN/uvZIveK5pmWFS3MYr
XHzggiZZOBoYIjqsXVlPGyuWwqBtESuuuAmasba5sCg4SYfKeE1vYNAfRla2b1Sz
mdHJBP6J6BOs9q9IYp02hvKJxs7led/vzhUp6q7GWSjT6j61JmkpCcTqS8eiEtLl
1bBk8mKU1DI3hJQFEk3jecjDj0KDaXQiUDdOz3s+Dw99C6+JyEdNe3Dsx/rzhHaK
XLlEJ+FoHRJzWwZwkapJSYkJNctWxkAqnbw4wTlLzJhlNi0n+o3cwMy+hvwXJeg1
iW4Y5LMfdDggPB3ep6WAVCUo7MAQGlmNbIfUlKXTTX/s1vYqX+6cdZw/sRntBdKF
XzlMMwPvYD+hA2LVYpJr2X1ze0ajXdlW6GPv3/lBc8rp/yjNGrGwr+3b3+cj5LL9
bTKSgxWsMrKzu7jeh/oTWW4GhuPrQUU2VLZPm/76hb10QHWXfqD08lZ0OvcdSnCD
HD1onGtaWvvIcTRTHQIpPZ9DTsF8rT0cJ4v08ms4Kqp1hh/ODQSArrzOaq8kS10u
tyvMBcDG57+pV9CXOle0wALAA6ckfzWgrIgGYA5sVX2ZzDsjZrApYDMD33SHhpqs
sZhBOh/1GsmHt48RubQjZGGlnSB9LnixwkdlnwbITNr55BSQFWNOg3FireyFIl7l
nO7obi7/Z9cNULETzsVUjdcKeZjCFcAeU4tWUhEtHTM97U/1TEkU5DqhzOEt8SdL
y3w0NIePML/qKoXVUKFhUFm+7wJWbvTSyEhfoB1YUdTnvNTIZOzBb4XWpTzg63cP
qheH11vWOTqf1krjP5/BB8diZgZFSR+YcZVXwVPOXfnS5CJO0DLHxoJrGjU9cWFv
XrT+hAVDB/ViYd0aSV+9t1bXxj2wGGHi9rfaw3ltFBi14TsRBSOUCVXhZGHhLLAe
ITIwej7cvSRU9gMzKE+jeLLt34iUrd6ZrvjLlMOYmWOp6rBBrNm4Gv8qFByqt7Bb
GkAWxVjh62lcwW0mwH3V/IMpR1ZiWkfbn69n4Rl2YtlLAwThsTpytruoMvC3B3EG
hmopk6qqRDUN5sFmduLR0JOfzYMlVnjN0CvmR02wmMAf0bmWC2j+K/eSHIx8f44v
6WRPe/Id6ZBu1F6J9IkTnp53EHpo2zICbWDZ356K/L2g6v/TJXziqPPqLmRVb9N3
c2+7RB7GmrR8I670TGHSWhxVT0PocGYo6omZQJz4m86WnWvrxEey4MitUSUrQ5dF
vbXR1joqmSRELVcN/62qv+wauXLb/c+K4R436XvPfYJdYA/1CYZ+jvKpyBDnou1Y
zBuXKpxEdXxdh2uG3mE4xJCgh0FdEipzle4RXafRl1oVhW9+bNCnRJsnsiRyGx3C
yow1KqC/9kTFL7BYJLXRAe+3LD0U6OEu9G/3OA4jDb2tz1IohkHgJJtaGx/TKlax
3rkzaDeSznwWZq9LgVJGPIpf9iYtnCPTk9O53awb0f3dEEWrVjAxtqFc+k6kyOB7
B848NFfbXSyYmNkiw4ZBeudFlqgTztdYIc07XGtjd1Ml0tBv9mJm9HIPtRBGifdu
aQqrDOk+lWUzCshP0xOe+dvJpU/4DjX0Yb031CixOHGuX0gMpwzh3rzMhvMonBc6
D9zBA4QKagUY2v8S8jOa4c37k5omCnBSL2mvjoMfg/zCVP8DreoVhk7Z3PCkcTNI
Et5Wd87am3W5uLrOiW+PVv8gCkLITKODflddnkHx5alNc4JelRMY4OnkyzB77Gcw
JKNkUXVV+LvMHMFst/QRoKLGMGQrWH/CfwoErYuEO5I/j9t15eAd96uZ52xD6ruZ
s+edMi6MXin16QjPXJ/Lh64/U3HT6bRcNDQ8M9PVC2d+gQ6Qru6KLOwsjXbpW6MI
QegUUt4wk/K1aJXAifcdrKbOQ1a/Z+8+COlAySpv4nTgnG9DcEwXThshvPmYv3WX
q57o7Qhpg2WWit2BpzrZWUFak6m02rXupGY3VmGAr+FnefrEsemIW1WALNePXcYc
/kCNawIEJvF7TZeagL3ft+f09heOT/ghiVN4pxV6ck1EVIhh2hMh9ZsLaV+gW0cC
UgMcORItabXEuKfCnRGpR9u7qDjEWKRRwWyZSw9yjFYXy/AChWw4z8CkmsJaBLwG
djmM4kCl6RWlbT4GvsrBRa318uFBIhXfxrASM9CoxDmS+oZ84ML+S4JLJTR1tHwa
`protect END_PROTECTED
