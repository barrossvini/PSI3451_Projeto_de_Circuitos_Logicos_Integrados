`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SS4yihYnXAzg1FIAh9JONc7NRkYIx4xZWcty8l/GUptZIgNSQd68r3EN29e3kFEV
Vhk2pVmT0euXUJhhMJfvKn151vGV+QLYfKTU1VrazPyeaKL0gfWCcbKowjoMEuMw
tKkNgNw5b5EfLD4F897oqB9gbJJqJnnSwKmx0eGhNIykZYA1QYeQTz9AwupIcovc
cquSBBuviT4DHXRbmUOC6uTYUwsKSkYQ6CrKRHFedvRbnvlGr30G+UOugi6tXod7
tj/PO8Nhy5RYNK6ZEqrBcRqy3dCwBSotD14ATI4XqNrhNmFkbHkmdk3grNFTGSF6
Wnq28WM7gRvd+R8R0IEn1wIpQmMijO21AVojg5tREoy171ingNzka2lKnrkrJyFS
Bp6/+yDP/I/0M+Z6O2ZBGFJHr5nxY/o63uumzJBwsEDPGX9nfk6zyFpGrZeCFpAh
ughhIjGZhMJpt7QKXrIbs/MtIpItVT3OvoobxnFVekSPVLdtl08cfS0LaVu6IZLk
aTCzwh8sOikYShdiZHvVZpQNtfp6dOIg6cg3EbMYNlAcsYpwatszC3TUX8Q1uwJ4
bXXS/BZa9T9/RxyeuyieqQwQES0AQ+vqwVU83seQVN7HIkAXZqO0FjNEMhBtyYB7
C7ucF7/FjAhcu5eOsasmqHevJGrGejKqXE+98+KKeM96yuxnK6dwQktjnnYwgGxk
rhB5KVjq9VKLEBNOHAS88+bUvRtabl/2QN4h7Ei+fuFBznn37g+OMH6MFvV2y6IN
Fey6xtMcATj+iZlmrbPYF8n7fdCe/5XXVE2RScUFYoLKUH58g7I9t/7cXXsVQzu9
hMXDN07qhh/JOkJ8upLLPMz8neg4Z4N5N7OF1sJog9SO1dRvDiCYpVyi7hi5wQ4U
AnxFkFUyajaynSH6/DgS/O0fTS8V3lrUAYv5uzhT5b6cygdMO3Wxz1eWesh/PR1R
U28YFdI38lJ6Kkr0NCHBOarkxyzAQHI9zqKAR8aS0HeSpdyKX8kKwIQvueYNzBwz
M2gerJJD/7TpBoADXCc5HWv/KPXGMW+5Niqh31lFaegz7RDGovzN6X9s5CgN29XV
GWiScYyiP4DX9Thfs76JeNOgv097KKtN4D07fdFHOAyTVco5CjUnK6j4H8MZQgwu
8V28D41G5df+64fmlyz46iePUF/8LEEehI72JuFyFLFs7HfjpkZsRtFRDvdF9uva
iySWQphk8p1nmOnt5lbeNVc07AYjDdQ0kpULsqU5nJ5C1Qd2w4uK+vDPoLegGlaR
0LRVyqdE/zydaMtun+M2A4PHSNnhPBM6YkaXRZ8WHvkRLKfbvK0HSvbqwVox3fEq
epj5AWbpsVqnCxPfwKaI8NiGUWsPknGdz+BTXUgYZYFMax+Dh/J2egXyEbSho9zI
PhTnxH0JMA9mc120VoCyXSTFIz4Bew+Ed9G8KS5wgbfZ9tw/hP5tHp5k9lI7uRXd
XmPYHff1XMU/xr65poOLy6lk4Py2BdsEjNSD8sJ6x3m9pId6lRR2elaeElysN3co
nDOWf8M9FWxNtZ+EONzTsA0K/yIz7m1Jm8EIjdOsV3T4SDrjzzUqOBf+LD2oWFAZ
srcKYg3rspHu+9eGEk/Z/Y8ygcw6PNgKK2HEKIPBULhLA7dRzgY8l9nXIWZ8AtHs
OlXno2B52F4bTwIiPHYe5WigI+xlvxBGVppfaPGplQ46GvfJjyl1EOejFl4dNDL0
38fNXvMmDymkwtl5U9s7mp+0AETpw1NREFXYNGn34SQ+gatOcPo8V1G86auqFyxP
W1qdYEB3Ie4nhJTf1MrIZ61afdtNayuCi4SJICR1VVK0VWNOBtFbo3GIklb0Kwl3
s13DwEZdVWwsd0sB1op9MA==
`protect END_PROTECTED
