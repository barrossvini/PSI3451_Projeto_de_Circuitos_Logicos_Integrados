`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/OCdJkwUkIG/jyLaMcqT+x1Es/6tWzQ6f4/KuIDr+mOD0wkZQ6RiuaLrZuu6RYdi
/aEFr2bRk6ifsgN+lsGX9OhFC3JjKOOuvll4+tdUukVLDWpvNrt6oto457mkrjPq
dwor9R6haW3mKwTB0MsLj9jV56a1zO1EfyJgV2d0ENFnYDr+B0fFHQ3fKJVaBCNN
grKZwxO7BLPIC7oLjB2fUrOYoZyjGkorRdwaAhZ1LaC1w/BBNQqfV6BeWzTcui+D
kGJI6PRne4Vo0lXGR8A9pWFMeTmJtv8pQm6In4ybJUpHpH50YwbMd3q98UoqXbkB
T1nZLHXEOBaazvWMWpHKDPzytI6YfCm/5BiRN3LkEGICuNR+IA0D8/FEJJr0KJYd
tAvk6fVz9bsUsdUlC5Pp0803oEMpt2ky+k5kHwTvalV43BR6YPQGFLwYxT1ZD/PT
rzMmKwR0w9+UzKKbk35EWghBtlB5t/BfD+sAYg4cSh5JVvpqxgN7AQF2R045cV23
vt3It1IdRCt3r6X1ZspHnFdGtwobq6dUJWwWnjk/MyIGOcWcLWx9THOh9uiOd1Ti
q/Vpx4RQN5JLGeGbfdXAwYvO4jS7VE5a1Lh0sp5g998+Tluax4cmdP6AB9t6J3fx
2+XfXFvIH0E8Lbaf+rvblsYkigkvNLVY4cGNda5Q2nuuZ4kJe3JV3e1AsPfiSv8Y
4sgPe1TdFP4TqFB2XqFSiE7C1tlT5W9C4zT4v0iZtBI=
`protect END_PROTECTED
