`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j/eQ58OZO2b3RpZsd+6hF+ETYIO+v2CWPhXlydxQiRG4ftYzjSa9bX7LggtFme9l
dTmG056eEVA1sglXbeCjylKVWKHmBqVaRbyBGEAYjdTZ1/D6vH7sRUIrL6u84GnI
X/hcrsOi4rk1qJp6H6wGGD5gXFQ1IcQvuLKESRmaLELmjRZRgGVzgCoQnqybA9ef
WciW3Dw77JBIouEp8zQykls5ANQcMfR58lOuJhSRsRcxqD9hRfYEzQVb+vqfIB2A
rHEPM8SAwSxwlKBecxu5B+ADKhErtMmcO2gjS4RHE3kXOz34faKXIZVWE5yiHffg
3c96MV+BgMUD03oD5aaerwnoOMhxUSuE5+20l0sj1HdKpTXhhKGRkREXaZlOzQul
9hdiXivb4tuLSvQ8qWAwdWsf/B2352pV9c6qZSxpqIP/W/JWJr9Zt5y02qaev4WW
wlU8x4WycOHzTlFM5qzT28B4ouYiJVg76s++ZRoAbzsY84WxHZrJXB3iTYBZKkg/
Qf+iQSPnUULjcMFUXnMcaz82jT5PU5WzflSiU01fpJOil2UxHtBW3SggWXQIuoeP
CIaBg80nfUFWJGaXg2adjQrUYL1505wncRvgeTfyGLlP1Ze5SmMGALHFU/Ur9Axi
l5sRysAYF+2Rdyu2nT1QZHv2uvFtjo5tH9Z6Keuageq37QRiIgLrYFHb0SOSVf6w
`protect END_PROTECTED
