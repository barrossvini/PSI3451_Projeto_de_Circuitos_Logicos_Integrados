`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ggnK56Vgt7mx1AWDzodzH6Jyznf8j609xikLwJpTCKKEZ0rWrd29UWgOQulRQif
eMPo1Hnd59DsfBF1sj9ob0PABZELB36+oM6cniEhCLHYp1A2v8zbXoEkX314ptUF
ct/MkvpEy9CEyh6e23gUtn7B+RNfFTeW1KtkUhwkBL8qf28y3cWkjMN6lMmmAV/b
l7RmEWy5Hbzxg3HL0sSzBMUstKwYTOcuC86FAeehQY+5QvMjwbTbforxdQKSlxxS
E3Rz3m31pU2nExzqrybynhNqw1VAlV16wMdaM8YcCZiMJ7/6tbTY86fXx0zE+NGn
SbVbPG9bi2WW304AOFZ432gRFUgqm0sdiu3rEQ8fWaqM8OcGtgcs4EEooGf+nwgX
BRhwWTsVJp21RZMVpIiJ/YfAqVPGaMbIBRnxoUl1jJP2ZRJjDz0Co68Ba0Kdc7nD
9sS0cMzw+k7nfNEhANxRs6MpH5Fj69gLWkeQoItVbR9IrpTFM3hRwTfqeVMKrNiY
Sh2gkUIrNqOBRRFNXgoOJO/7z329Y6fPODodSgT+ZouBrHNa+SDG9cDALfdY2U74
eYxsLDGyQ76pgSfy9d6fZMoj5wrDUK0yIvpS+W/tB0VvTAPwfVMpWmaeigzKYlnz
`protect END_PROTECTED
