`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q1TwrIPRBK+qNIqonQn/Mcz1NC0wxQo6xfp105U3AR5L3POsV2THOaySy9PmMYgm
K1r67NIkm6/p3yk6lPYKagzlMS9hWIZ2GXbjQLGHUDmSBkx7MzqBCPi81tOOJraC
vEwOZd9HJNpJWKM7x7n7OILuj/RWBmJlfApfrN3y6CW6hyJYfnOYi3aRhQZPiWBO
zfEuW3M6ThNK3lQG+xAAz3l82dG9My5Y+ryDRatUckgilHdUshQuqWQ5Krz+b6H8
QZ5TJbeR9BAB0O5wA7GS2AE47Snwe9CXXCcndC8LlUCm1OfYTX/ghHxHllGGgS0P
oW4M8hFL0XYKHlHIbKICYugdlruhYCt567xQcpHtjh5IMs14FvN0JxwofmjSUKeD
Hy2oqSKk4nWXCs3GpRkEbcA6v7ab5Gf8oZmWyrOTGOtrgc7LflpzaiAa5VADoEVJ
GCx2TNssjHM1fFDedZW7H+LPBYZ2w70nP+hEfgcwMbA+2M2zO9mY//4HJKg0KWmB
SrG+7gMTXBpTHw0pXzuTCtIctjhxABKvt+9Mdy1fu+kmZ5bscg9WJWRj/0N2jY5h
HCi5I4aUF5FJopRISn6TMYrq4Coylh1dOmtT0i/zf8ZZ1iCw2ZWoIJxQiEqx5AiT
0NWhcD+E8vmVmdRX3peJjmlkRX40GciaVqZoCAWHUAwOEAT6mwvDycDgcGq6gaHs
PEABHZv1Y1adoPqstzaBLFbH0dbbWd4dG9HMClyZX2M=
`protect END_PROTECTED
