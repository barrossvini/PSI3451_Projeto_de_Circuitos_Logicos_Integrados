`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+cUx+PwH5U9FaQcN7SeJbzvI1gNN8oe3GeApTSZAm+d6WcJmYHFm0yfC9hXaioT
mZlKVkYxiBk4SQVXeW+4l3gDrHoGSd8wGXyFNtVWdJMzQOIEqePjCmv6PlEvjzYo
I7QL1MoKv1t/eRFxGUfN2MB2sB7l+rw8wTOWtcI0MajSxzzZhnkghp3QXuSaudPD
9aR6wN+MZayW6THJaHT/jAHS+DM8bu0kA6xtjJOxe2EfCut5W7aKL7AHzOB+aEx0
eV5Q/j6bOp1xioyed3VPDTQtXtVPqIXQwdT4Ud2nNuR5wxFbg67p0hAb+VD4ZtTJ
twM0FLfxkhL3n25xqdqgibpYIwr0NL1M6FbNHuqdDYu3h1cirjOgaKtxfkt4ugt3
zJpuYouH8y//PEywGMD4C5ip9h/VcG8rMFJmynyrUg8D3+KWTaYaBeI0TDxWSI+V
jur16oWoXCyxLNHh1tdlJMUKcK22d/t/+LWCvCEPDSnsxXqSyTfKkK0wghKH/rLp
k8ZD58v1oNjND9UKFbtyMECi1eWMcvl/0ylJPUtN6M+jlXGqPpNmRHPoSZQi58HD
nBfwOOT82SbVQAApkUdOppAoxMBRramQ9/njBpGLVLJEDbzbuzpEc1P8IKuvpAt8
nLCnIjFYvy3uA9MacZVYaPnRzz8auL733dS2OkDjRMClki4bAoexa6WPTWxxO2Jq
qtf7ZwGAAbSmB0Z4OTj7fMOnXYv9+vWBmwVak/I7qnza8fRa2tp+iQUPhmyHHHTX
XevTtFhCYIJk1JOxpkMAqIJ9DQXEFCaevVNlBc4EIsr+QZ/KUprfMsjle01tItM5
axgjPKVvRx+/VW+o1mhpdwaNi2LvdpICiCLuxeaGCbZwaedeZCEPWHpJMtQ/JGow
BOp9jWrneW0AFMu5VDMMSbJ4Zf7+96uMEDjYXpl/6NWrFtR4b5igeMlwkxTM6j3n
wxsh/vImN1hh/6SFWq1Drh1SOloMH2bGCuFl35gTlLG4mA+iq4j6mV321yOIXoAf
kBhOI2xzosbRIGmr2csDqqfoQfq0Ib4EvjoczmBsHus8EAn68wfwQVOICDWA/mOm
tgnka7LlufSRciGqlQAq5JxqPljFHDzMAM9MhffkuPAD9LKvinQQ8BjPpK0x66rp
Y7BwqWcPZo02Cl/dnQvuiWbK0dy8B28GojWxkTgTwviKO5KWqGzxhqaLfVkk2m1B
1gD41vuoVWK+1d1hrCb19fbNDMz114jwAj6ONdNkqLZo+pSdkmClges9gys5U4Eu
3J1FIhmrGHYXwIUQC9IZzSfLdl3nTwxGbuwCetIAwfXOFM1Q9ZOVUxAMULRZ+Mq/
ANE88Za1IxxV3sGWWROr6f6omzLoSv91tfoH/Ehu+BZlXw4JbY5Wi7Xn6eou76H9
zpgLmMNUG+CYQ/iEc+VsJ4/YSqBxbtxbwxGk1EQ0xz755vWG/3G2jsTtbVaE5Wsc
o1sOGx4sJTf2PzE4pxl0M8bMTxPWvKfqHpNlbY2xiAD0nt3fcMlttm6TRBzYypty
bTJTdvCfrL3dgE7WB+6qotuV51VWXauYKLtPKe/YYLEX0NY8MtA38GTuV1kQgM4P
ZXyshAjP1beuy2Fe9LmpRiBDZ8L4LXDijRgdsTbTXtNK9cvNHBHeq4zF9AIzhIKQ
s8dgsLfVuYRDiCObJ2wbJ2ZjK+9AYWXReLjNyLd+2bY3wnPMNLj1DOpBPEneRDiH
Ex5MJ7KA4rPm4PRSgRQNOzq8G6rch5Y1/WFc8sayrj0xc38rZ5ekB1EklfjNKhtD
erkr7dEQALOUuvFj0SzPpfWrrz/C596GqQ4kTvEzWR5w6uEwlQDeaP6NegiEgvsC
YfX4lQ1J7/FY/22QS1ZAggFa0cUN6/8TpKr/1Kdws23ggli+ETX18UEwJSyCloTb
aHfDuhumIs2Rv1QL/CJmwZYQOnUtmV6o3Rw0Tmg/y61f5B79cUxcWfxtjI/J8d00
5r1T8WChgG4m91MRs/es908mQpc32vqOdZRvoq1yTMSNHqFvX5Een/AVai/vsDDr
jWM14RkeLt+u3qt7LJx5WzvNXswscRuipVE77qlnRHblzRvHIu4t6x8ZvN7vIyl5
3tFRpB+at2Hx3QwrNe6WMxASu1Wni3G+LHdmYjzS5etrZEl6NXsc4GU90y8vautZ
wIKDFUNnA8mlRN/Tv7PxQXAFi0AkeapoTQlcD0WbMLGQfPoV4x65t1Bx7DNZ1zCd
gUM3pOxQ4bSiCvzOwD7bFpgEpstHFfRb/xUP6gwdUzXIAlioWtKVvcnYNM9J2/A/
FRvsAz1lX9gp50RJcQyGBh4U64bHeEGhap4OAlzted/D+aT+eGtjTsOzMztXfP61
gor0mqAQIhfeBbNZMdTk+PHAWdd3YZA5RykUNGzyjHQdLjpeE8PQKC1BUigBrfwH
Z4qt0cMsSgeWqgo2hkMrRYE+5jTu9OqMqpCOxK/moD16frGDDSd5vnWMGPyDHD2s
d2ECstp3sYKxPTN38anIo4orgWfqW6eo2DJsyIOORDolbw2q3ExT9O7VGMX3r53T
FLVk8kQFnjhLHSkJyjHKnEyTbHR8eRM//ervuEIuLfv6Cxa69bTRrZaj7VVM4v3C
wzl5tFE3cgiJVo0qdfw+Vg4BNdEEpH6URmZwlYU4gcZ4VPB1fGlprnsNtAE4neL2
1KV3hwGAWl3GUVP+0Rpn3mS6k/qUvd+XWuMYws0WgUoikdEDr9VFYi7f9P5zjahC
GkWyeSMhKyxiFPiGzur4ZKKP2Bw6x2z8h3clnJ6mTGUS60UP83JDsVvvnMowqaP7
lkRzIj+a/3rFAKb8t/q77gEVH0/mt1zpnkraYuKg3Q6pqsPR1UYDcL9uE8eNUfhO
VhtDX9IhPD7WwWdippSOxX7N2RwRYFVuGYFZUpj3tz8di489flBZzwE+XsK9Pz/p
qwB9UGF7JpIbwpbrOKX3Ujw88o91cNEa1IxVkBQU+NNIN92JMMVa5WbdvwYTWUMF
C1fXnn4H8mgQm7F6Dkd++1M6dt00iZVJoYbKX1udsS9Ss4Dwq0UFJQl1nilkFOEu
+mpSEABjv2gtgRrt83qO11jrC/Gik9NDXVumrBbALFN7G/alDjtPoK8rDa6Aj2ax
RSI+m7/Mrc1xVaMpym2ggBPybJwo+fK994G/uC9u4dMjaOkavi9TKLzfTfrMCHO1
H0sWdlWdJ2zckSpQKsfC9f06ABmqJFeeNMt6qUDwh2itVGf9nagzsPWUAWkE4aGS
WGb4U1niyNDT/AjB1diLoU4Fd5pjq6EKtkijQwae9kchumZezu5tGpWhHOk6mlDV
HLfaIQEv+yarX0WN2bf64w==
`protect END_PROTECTED
