`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uGWIjMH1aHzQ4UaTpVpyB33ckD6x1x5Z8B1dHg5uunnNyrfAiLtcI9qpchPNHY5I
4rWzqRiVVi3UJI9k8un7WtUB8qG6QzRtY61hn6t1MhKLZ3MOfBiztgM2CwTpGI8F
y1c6MswE8OEJbsJdeqTIoPyCsdK90ACSO/04/+aiP316gbdWs4h7wH5UX/oOMZ8O
V9NOxyr8Ii1TrbN0cTlm0yfHHbz96BYdxC1Vxsse8PkAjyPyx+kFuLjD7H/WlReQ
fpiMZ22aqxto9HdW8G8TULE0GssWhRwrQ4wilydoYo8hobj93QbeDzVj3EdF52ZI
ra08H8yZSUlYZXNtsIAu+f7K0Be1YcpIP1ntxF+jq0ZwpfpguKre/pCBv3GC7duZ
Yf2BMPwKgh+foBIQAB8XBg6Zu9qk5+U93W60sG0ZEaahDVq5EX96Vprctxq2AdY5
DTc2vdqREuDlHG8L5ERjKgX5MBcylB2FzHTSC9+ufiXK+OWraC7NlYa89XUu1FsH
bBRbQGGgjfnr4dagGlsKbpsAjLVlMjKSNf7JkdpXgyc1DStHUriLspmY6ZVFYkkb
ZAp4JMB3ucy4lGGP0rfPxnC0Awy2yjId3XudJJ8R5/50Ovit7fZFItN1zT4/ZuzB
7TYvk0/thlQFrAm1eKJYf8jmNLlwSV0t6tya8JQ3+jC0dz2y1t/Q2LjjWPtyJxz7
gSMRck8sUKiPBTRB3RVpWaoahO3sf64NtK0dke/2VY1HVBsjrCHmRYP+cKi8m1lu
FAvuYIzKmGz9ZRUlE3/tqMM72BTrNoR7p5b6GgG9RKmSH98Uj46cWWR5n/eg/hGr
07TxQwhEqIt6/IvXOD3+KIMpvUGxKyC6tAvV56MrEMpPoxDyszxosLUuqAjOHpaM
nNXta3aRqe7d2JuP9h7xJIQHuanC84jdoSxoYN1qbW6Swqlt4q9rqAg+DsoJCRGa
lVi2mrkguOwWKSncob3HrfLVl2pF9TZgmxhDCK2HuLY1q+l2XNMxQD3UWuuoy2Ja
XInbEU0bMjRPKQ0PkTBA1OdRaZ4f2I939JLJJii9ioryCud0E5qJj0KPijNCHyZI
eTs6KZ/tedlBbwxrXx4H3Q==
`protect END_PROTECTED
