`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ae0dguwqwWjoxRJfKRZG3bSWNiGPM9aIMf+/ocxceBX1tYeKu5U2PIZogPo9dD6S
vXrTwzCLTLNNGBl/ayt3QKQZUGXux4WCq3xCtSIBpStgpl3gJKJntKLa4uDBiQhO
g7WjsM80eglTkQvvdWHXc7tddDFgAwNkeREEZz9zA0xovnKyqlOPM5kAhc3liqZm
HalIybZ9CDPSNH1nyK49y3TyJ1PLD+2aEySY5W6b3kBwCX56O/aqWt6so4Die3yy
6faNm6HAQmxP/Krh3rrHztLygRepzgyxyX5wMtW4F9ZasTXFFpRiw/uF1wqFRAlj
BENHaPaOYKrjsu/c+Kxh2Kz7f/XzEJHbXNaENQ8G1PhGXU1GKGKLVUZEeNYvFMXf
BFqyYi1/513uaMf7pLSLoLzV2OH73ZWJhfQpc/Poti9ctSXMngEaWhFDDUMI8qfG
yOQgR1lX7BgvBNX182BB1/g/z64R+jjbF9DymQnQdFMxocL4VLAOIgogOsX6E79k
ZmdWIGx1bBnOOfU55wOiqjwc7PWGAN/HaFQMcEKrcfRZXToFa3ao2TaSppUAGTtl
DS0TpE2kzgLTBLqD10WseHwJZZy7LEOkLvzud55yVQj3QPWurjgqpFdm4jE5xaz3
HdyLpQULN0fm1qaaZpIa4ZCjagsfr9J/tB17DemPmmJnFLJQg3tqtEhFo5Mjlqsn
n0J6v91HAIpuWau5VnRkOQ+2zy+6X9cQhGa9SA0s/Vi58tg/mkXtl1XwA4RBkSsc
hsNNCYJSNBTeYhjQEXffxkCi6jlWpl+jYAnSbk6tvJbBEOeqCENrsgNwP/1dd02H
eyDWnsEySX5nRopnzNm0szxx0L22+5nkh/hVaXV+1wmKpeQWBvVdO/wrNFfoLU6O
n5FF+fpcPtKu9mP9Swj2aP57K7U7PA3fRew/hr0XBQS8nqM29YmRx2Wq1AF/TYp3
`protect END_PROTECTED
