`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQzLnxeO5YKI5a6MLxNL05lCBugnH6ihWshCEvELmF5vu1Laa71POt8etU3KwPuU
CF6TDj8LPs74360jP/KJQDveGqLPjg+JQZimu+m+3b/VIKU+dk/l7MbslgVlkQsV
CUXdjg9LOE26g9X4BoitWFHwMe4xP89SXA9qHmewL7cdasEIJVeCRf9VwfPzuwP7
7ESdYQndIYsLD9eV7fG2xddPh4jLykKlAlU658DnbzOuDOqXxnnCHOm6Sh0zY0iA
PMEd6gjjCKSKrTW0vx3M5fUV3oopYgPCl27jd7w78ULTMJx3k2hlI5+pSHsaw4O1
mG3yHwoWpweQrboe9XSdKD45D0mDmGj73QoTuDROvjJ1Cirwfsy65wp3rdRoTb1p
tSgiLg7NVUtN2JTWuWmSmR0hm8tbH02Wk/UueZ27WovfSS+4UWjGgXU5EUamS/sm
KCeI3u/lcYU9zpEK3CI+U1UG8OsdfeOEykbVKBYP1nMfhNwELWRnHrIGtSnZw5zF
Nq9InFummk4gGPspbyYhs4K2nz5qw+k7DyPnibvbF9M+3Y9+abpb2TuqLdZZi7NV
zJ2zVgjSG+s96+2BQuH5gh/8UNQKIyDUEBWPks65BxxPkR/AK2KeDAbuJbn8rz+d
0YC/6Hfnv9Nv6Ki+HnvHKyqX9vtV2YE9Eqm5y7KQSTJATpBB7rGkAXt8iu1+FYK+
qDsuEa+oHJtj0px72K413UB46+hLxQdN0+STylqEJMCeO9fnNwiub3LNCkaYe53O
Tyb/UFKwXAdMXZybQ9jg81zJUpNlGFJjlUPmDRfU/us0dEaG1AlpBewAzUaTo6OK
L2fje47/3BOzJPYM8CJhCUfHcuAUyuwADuEqBAMhaKj41VbMlIanJgslVdWXAntf
wsFFwB5h8bdox16sqz+AeW6RFBqFDrD24SL7v8Rs675GwDXiRxZMqqqwka6FiW7v
8sznq/ePbcUIEoNKSFe5m8NDVM7kPmMIpBi8YLyiguhcGXbXoeKH874H6X13SCDb
I7vX4IG8++a6Q91K+RIltyiGZsoCJP2+GPsGH5o9rDSq3ggNeZHAOlAlrQqQfGwT
PvrK1NZ24cNTRHPPafJybpY/zihDMD7h/NOazB4lvLLeSoDnWUzP1gn7yjNVf0FD
Q++e0zRE+61RmN26ZcP2ASUQ+j3FLx2z/MD1ELa2Sv1PjcyyJxJPhS2dztXRffft
Cvvn0SlhCN6/quxn5izRE8S4s0xpjye2i8KFJhixzuEJhcjzLs3CcI63tHWCFfhP
PfnXS/eeOtVC26AB7OBq45s4X7LNvUwg2yQQfQIClmJiiZXEuOXF7/Z8wlzrKnrt
CD/OX6yXPh6BuG+ntWXblws6H6/a7jVjDHbGWZajko8h97b3aVWMiKIZx7tYvqEP
G3Gio71hhVMeaUJtBG3uIXb9Kw9JKlPS2zoaAbGQck6xWgddeqw6q773RBBnohwM
nPvdvTOWHdPzchovIuugqk/GgBP4uf6qFZLuUUYcs1dhj73PhoxV+ccXr+24Hy1T
IGPEEbkhKZS3qAO0tQRI4WDmBTrU/O9n3I0eUmqrqxtKUTNd7BAnu5AbWym+Zv5A
wPbk95lLsP1YVP1HbonDf96Xxe6n8XYAPQLLLw0IApNxH8Jjv4gMNdL7QbHaPUQt
zSKm9Dbhd9ziyDxQvVlIyOPIdyuneHyWp0ok4DUQXj64GK0oqnfMU0v489Nf0V7a
huQ2mBtYcQmwDF3Dk7YsI+RaprZWGAdStKe8dKeIgHCy53P/apSftUN43oIkUjPq
4/kw0+M8gGrSOl2bs25GeZno+pfF/SvKfOGrRdFK7uFz5K4gELGQM3Yl9pfnl4Xp
NSTkDjbo0JRbOY48pVuivGDH2BU0kYZNabCu1AGMy6+CIUyyHuDIepSWEjK6Ermm
DOVUOuQzYxmgC9WcO/CilLO4/XBvk9ZJn2GTzF78Q95Y6S54sPikuyqaut+mceYO
Lj1eg+MiADZedTgw08pd73nMG+1nLQia1Bz6uMFMTAIOKOis1nivB++UYyUIrOMY
mXowFu7ECL44/rrf6yAFPSafK6F1L+xUPoMVtDPBhaLkA/EZBxFl6GyBkoy1yp2j
iwI93zSEIntGLtV3y9oquAepPIxRJOaZAFcI6Y0crLLuckAXVE2CSZ1oGMsk3kkT
JRazr6hm4ZCKEioDlJ8XCqBYjntuERcpDgZiMGXLzxImQIcUSqdrd/7QEOYKjupN
8i5MRmPUXNevNPqnrSReEhqOV0xX8WbKTZQFd7oVZ0gkS5bohiaH9cYgLSzfuvGD
Ff3udy2WTdVReJdMooOfE/r5FP1J8HsAp4V9hj4q5n4el9Y7kSnWJ1L40S1pQP0q
FJRDOGyN4J70t+SBxyUVgejzzGjdkx7YfJcFEbvNHZNap/uVmSVzz1Al2NU5jssO
pT7df3yqZUBynFsFT1E6bMR55YtlpnQSFsmRbMSsQO4AzXE8QpQovaQ30q1BKcOY
r+cgO7FxvCmu1KA7Be3zPzGUgiKB6ZD3qm9CBH7GqkPumYNjTPBSSsViW66/JfSY
SxE3SR3u84nmWNc1z5+RPdufxuu/+pWY05dl5Anh4j82I/jX5Gv9SdPovRxu9FhR
uNhtBtRXmpPeDKvQO4dHfR72CsSJ4vdQ1Blo4Tw9JiSHqYNPazmBQBnGtCiXx1RO
m2ddvtEWKOvPpw05QGTeNUKoTnR4NnD8AZxM2FJIbh7lKNP9vIutVcQlUKtZ3+UK
w+UMPq6v51JM1vtR0cl84iKdzzYg1sISKmxw1MfjGXVmSWoV+wQZM9td2iTg1KvP
7uqB24xj+4ZsMoCD9UNtSKraItvzYJiqfsTLjV0UG09uSFeeRq7LubXqjsLLdY2m
1m8aepUDqQrhmBVkzZWHMN4oO/rnQ4f4gLrqMpS4rOpMnEv2LYhNyJP1LFE5rxAH
JyrABS/IJhWLSDeULDMuGhn+Ey0KEb6550PujRVYB1Bwm8fyuDg+QzZQrsaus8vi
ZG2k6Fv76VYXoJALHDpvnoRywB6ejYh1zP4aX0X6hOl7vrQIcVLDKT7VgJoDvzXL
h8qFlyYywfiFPsEma2pPuQJqW8Q0uHiwgLoAZ/tufz25VIbmpdqNDmBwFR48ZCGU
sVt00S66+XviW8y2fCnr/zFU5/aixPiw1kKQMeq1sG3FqUBtDonM4+3sTYj+eWt4
5adwKgecumovL7PQ3bwPE5VfHOnZzs2vzhkqauzEmM133w0/MyvJ4VBfl2cxB2j3
jNp/5jyvEHBk9dNQG9KlByiNsVfewcWUwrQspSrHjJY0kGpg2hd3wHDcBk4oUMjU
eeMH5tf8N0qtbLCpbSPF+FWwM0KVhTmQBlVbtMYj1yRbM2D59Pcef86wheCxEWUp
DgRPRDjP+pcWij65b8BMbthmWG/cptM3uBCKVrQT1oDvJJYM+K5LwXZalvTHd6vz
t/Mwe+1LugD5ofkRopRKoKNTo5FcuT1NQC+p+gkAdFjaXL/54rVE94txjwsBmaxf
7HF8mee4/MBlUeMHz2DPMOaxNVdpGyraHIyhJyjVSJyfZ0/SiNO9GLtN3sRexg6n
jxJEx/T63s6lknjp/dwExCcXjR9Ly14Q+RB2FX9y7MV4tSVvh3JGzcv8iMAjTohK
LO48IfqbqQxsDZUIrYsxgg==
`protect END_PROTECTED
