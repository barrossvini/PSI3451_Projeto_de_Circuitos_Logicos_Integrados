`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C8sxDHZl9q/1D/DErRehaTWn+l2t/trENR3q23rLXFkr+iOhue9yIJE9pv/OHGYL
SEOwcZwOhM7n/8bWPv3e1z7TpXnXnetrQf/j0iu+oNTSrRPaeWIvTx0kX0SzlMPj
tsFrc/HWPqyMjlWF/lQYiEwcn2BV14G8ejmz+S1ylA/RvU9zub9Nme4B4bn4/w4s
EeScHiXolEcizqrWphITl5Yo/v8oJpUAt43UPcmjnUuaS7Fd9VMX9cmmNrAyJIFb
/ud0CeDgNHwWqolzuIiUUwS5EuRhaXmgSTJWLrWXxa58h2PP/i650dDeFf7eYtnR
D9V7m6MXbCF7YAwgeJGAqN7tPhyX1KUJOldez46U70fv4plAN/v9+hbdJBBu5eYb
nZgW2hUO/FOrBqKb+j7DWj8G1JapbC8sunUHjB4o3maEPQAXM/NiK/jfpDEMbn5/
8xvSI5JD1+rBSfX2BVeeryvsG+5omqzwbL8Nr2W7U3Rr1C9ZN29AxqtM4TZn2wJj
abpXc8K53deWnTKoHImi+X1PMbe4cM1MKLCUb9Jl90vUCeGKSvmKejOhyrQDQ2SW
xLJbuK4Z7q5ql/IHgn1tPTR84DLTVoc2O1iZ3HdDxt2/3Fz+jlx90OajlUr+GDXs
GNsANeZ59HgbeXcsg96ZREIqRmJIyiSNgEB6dcGYrawN7T+Im7cHVSNy0sZHoZOi
3061/R4uAf37FHiN+aVBafhNRTjHmPisAsCCuLXAkTQOL5SAOzd6d//QSJLp2Ea7
R9PoW6BbAmVMpOAFaI4ZdGG33CrM26Wh/zrRrcOtH9vclq3itx93UhS52P565vVG
6Gh250WMk0hrjwBbtsCG9LgwIKc6G2TuYIC23q2clj3S2FPtc78zU5F0cjqHDVnd
VJDMj8bRgTU6eTOAYh4sMmLewgRVt/NAhA6kWdySOU0dSz38DU0HcmfncNVq2/m1
hbVrPh/HnAEBICOInqOh9VrZy39RKEie7cE9O9/s8mtq9xOJ+cWU+dHwMDL8cwGN
JyxWf7ejJIx588dhOFkzFF1whCXj63AprkpNkYTZpTrBpsn1MBT+HgUT4W7IrsHj
IWKTpyjv0HYh8pdtBKiTqBIBp+VD7evmY6vVjmhcfwhEOS89A02otIjXUmyEp4TM
l5E41MgWf0vfinJgngyIGlDk7ZCD0Eq0HSW+YeFdvIiexSjyRJhvar1R4dH7Zfoa
VrTk6UHdoPXd3q+LYnj7phPArVQolzF6EzRVGPuhmtwrHHufjnAwAWBeCSg2sKyC
ki+4KsV9E4fCSah/SwgNh92lgW4mjN7e+vsQ/+7MTkz0AmKOEkGWnsITw3li0PLt
zaMvg1CYoQa6VqZZD2N2/1FHAir3PwyAq1LyLLWbI1YF4ORhvVjOwTsWVdmkX22R
PO8IFBCLPbPWP5azseALtsMiUhcn6DNua+bPeir4kc3mplyUTBNRNl/zNyhyfGd3
I/r2FyZhEypPEwleJuPiploUUpBVUmeH95NVrrXJ+Q7UK41FK310RB61pnUfg9/O
mfUvXsOWrlJpZNyiqhyqdA6jhKWl7XMj/86vBRYleTgdV793AeAz5FideJ9qq6pk
5tWvTUbpn9QQ4NsuAALu1CptWiFPMqobE34RfWHi8hb/u8bjv3T4DmbJaxMo4k5B
Uhk5VwtmqOFtybeYdNkzTVaaXpl61bsJPkqCzuAOvpFJOAq0qDdAxbhCWfygHfPt
18DQFGKjpEFO/J/hMpB0Smuy3H1AXljL9RMO3fAws7RXkAGvHPA0RRkkMbaG0Oh/
4lW23V5vFlpNfdLwOI/4S9l8wl4kcnp4WxDSfI1A5bXMew0eBKmR2iw6PX7NICQb
CEdz6BozV9jdNw41KhaFC8CRV4X7HpYR/ogOZz5SJ34SE/0szSgdY936ralFzqcJ
zZcX5BDeYbcT6dQD0Ca7I+yeFHQQpUffYXJV2zvpGyX7jR6OHFO3QBvI4Wo988Ck
K9zn6XC+1hgCFJaqwOK4Eh0LzYrrbLgvUxQAJkGV4prswjYU6ZRbzRHxlwlQ3uPX
BFRAdWjDG4I26qd596jduG8M7Yd4ZqlmPg4DQgecyLO3MakAuvd7Mhh7desgvNAn
1mXW9UPT3MyMzICa5wjd9TGtiHW8TN0EbS1ypL6DwGOD03cm9+HTOBf27F/uW6e6
5iTerNFty6ACJz6BrMCJel5KuSl3TJYvfDsw+VLdr0w+pn2QtRcPssfpO9D21dOM
VRzjdNx5qqVHW78CFM9uvwSk2pLclFca/lz2dm/typa975p6P6K0MsyzFjtwC0Sg
o7FKbqpbPF3/Ba/ZkR+xMuEGOIi1Z0/pg5m3dqbDtdOCwLk6nlMGIuxVpfpJUKDa
ZjQiItQIlx9WRVNxYzEbLRXxZj64PN3FLSZC0mJEBp6rptT94Xpvhq8vvXYoxMlY
BN7DMmQLyF7OLAEiDoIEqsS+VZxJd/1Ks/9EFzjhNACkWBqUYDtCMuqIEVYz5I7c
MncmIeakg9fhDHaoObFlnqJK444VCWR0IIBhCQOBprIAi14ag2XT7wnpyebv1I0K
Y8QMl2rMlJK7xajHBeUHtanu0M1BEVFFtEKsJrS60R9p+fzhbFPa/oEnlfGO1nd+
9XXoXGBZl5dGqxlphqVapQOtNCn7T9UGABagMf7gvBi7gc3iRQJf2Cirj7Del90z
iuxtdbV1bydtxEnHb7RvY95+6DAZhhGS9rPjMoct7WF9iqJUipsaZMABPGtzszsg
`protect END_PROTECTED
