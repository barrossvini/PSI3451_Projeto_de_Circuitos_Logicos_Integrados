`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zJJGXPledrhPT8KkIJrzVy+NaIj32snXcEms7gwurQjFAM5B0Jvwmog0yMmOX87g
XW25vspf6qGpr8kliTo3mrhbb4bPy+kBFb2BS96cy1mtW3X1IAOT2YPxYUWQW01P
yB8GyiZ2X0gTTHlS0w15m1YytoXBpTqPlbuHVFKQuHkrFoQMySY0n7GlbKNBseih
RjXF2D+nl10A4NZeELe6Pq9wFJSJjys/EN+z6rVOHwufI1sC8RuOWDHNw0siyP7k
CyAFXOj/vWrpO4jxcNW9JRUFscwqfNrIiZnrqHwZbLgJWC9i6yaMXzskTzzX6Bcs
U8pV4xTcIb4JDa0dU2qdzhHtgojRPT5Rw/l4rGrSLPX7YH31Igz3gSxIUEt/Coiu
4E3kiaCOGkTkpteq1VJodrN/JwMJCqvb6L3In1G9Dc4=
`protect END_PROTECTED
