`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
revdpIFiosDnynm6Ew5HgrBanD+PuXC+hQlDwKl3KyxseMWWbYCZ4KdIRqT2pWHt
guRxQXkPnqgSSjRsixG9KznBurtkdCk8AAdSdd3TnTY1FDSP6Ixg6100EyVHOTlC
NThlAbDTi/PSTFuUqnZFsMfzPM3e0vs08YzRg+bBkPqWnMCfAnwBMJdkEfWTEyVc
wONxWUTEtnfhkmirS63LDyGfs9O5DlJCaiFEQQyA5KDe0uYGfpz96K9mIXZKObe+
V30JiRXzuVHyQxs2epSCGD0NQMsbx54LZqNr+mHbgGL0W0qkSTFbtYDxPHaulc25
DVOGhT+m88ZlyYiPVFv9SPRY9Q5gKH6qlxQkAPaEeroKO/BU9934aQpLYEC90kGT
NT4ZPxvylxebuWi7pxBrUNgtBtPGeMdPAPL5zh7ocldapHYw9v3U0Tz1NkgvHtWN
yGF/OmoA/IYhf500BagLxsNNp5oT9lyS4Hmzv+kb7w6lhc9HPa8U7ZMyhi8W9ZYH
+2AjBkSk1gFwmivj5W51q5cpOH1zttGRXV1J6Idj0FqvZBF0NbDrCVOuv64QZTll
CEZLcUHq34pz0Ls4WBXlurRW7k+1LamSUv30bJnrKkIoglmzsKVtNXE8eYDGz52G
fgBoL18WsfE6xoWAqsw42Obnv64nTJeiwV3Mh5xciQYsDRZaGfEzaWipD6rO1cjN
f9hPR1On4I0gVF+x2p5dNkhu6wQyymV+bRsXYMCGlcjLjHFUnPj2qfAZJ30wxZE4
zRQdRGgqGrI1qLjMxlxCt0jSr5cNX5WzRWWwcyRXtI4otoxaXVUnaan++TIHvx9v
Yh0o9iWwY/1C1Aqe2suuuy4TlAzaAzSUg/D8ufqOmFCBMKYF6biSGZdX1c5/O4QR
SvQMierRzMKu0YjlewJwKIRtnIDQ620JrHj9guvT0BVMfcE8avNfvL7TIXTeNafG
3vdWIhJT80Y5hNIVpEDJKqCHnePnFGQLtEBrag5fA9cfV+UDgAO3FHAABg/d7aUI
rXamPANaL2pMcDAaVFosckhHuvacWH45XEU3NQIy6UTj4npzAEon8C3XajTbLjXU
`protect END_PROTECTED
