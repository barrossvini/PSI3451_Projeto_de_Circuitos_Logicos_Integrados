`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tzQK5rc/s0LPrueca1JUeaGeY+g0SX/B9T3fl5FVtjrrIxs8eXvaa+FonlYfftel
RoxOySVjeuTenUiAmBERwfWuX09lvg58gAAt6fA+SW7GDpdX7/A2vIvze01FMjHu
m+/i6IIo/dIcWm1capwjDknnsWsbYns7d5CXlzwCjha5Ybo51nB8vTu8yivCvJub
0HrtPH1ZMHANUTfwYSZbBGbp8VsRUM77wM0jwAi+072QNewK1qWVVUStSEWOAk/C
vf7KfgbK6ykYaz+di51ADTkgl+MUivrlFgfGhn7icHZWhCcNULWuQMkfmOPEwhLM
jmcdD6yKEAcibNHuZdI6t9fQ2sRvy5L180lVV8LiUP+h0CxZIs0YnaQoDP/l/8FG
SPertnVu5T3pGpSQnH77eKk6Ea8yTTlnw1rhCSoA/boXyO+HELRYi+VFS3Sa1Wf8
7zyOOt1IbBqNddvzifyzPH1TWKlJ9gaMeGyoRRqbJBUtQXP4ZZEriVcneBOHabiY
cZqTeHhbTGtbNYlX/WRjeZpdaNEp/qmgA1tnRmKOP/rZDvBxG45LHF3rX8X92QYd
44FukE40QTLEcYTS1S3eZcWkJ3djWE0CY6MP94CySlKXEvw7Ny6ooRvOILkOjOrV
6aqXk4jMZIbeE6SKrRRzQOGohZWAsiFdGAwXpRa4qekP2zeq3mAYEDeBsMA/972N
Q8TcahFW2yEdMBCwx2TmTRg7FzJ6tVSllg9F8PV1day3ahtugEEru886A5r762n3
z99jWr0VVQ4ipUMCpaQTvZiMud8l/O40K1bAIM9muLd88WG5eU3LzPWvcsvOC9rU
0Ao49qxp4O7K31gghcjtsGa4UjvRy1baIsjHYR3QUp2speGaBOlty6J5PEBpGPVK
rUn3YdRWXbTL5UO+1jlgYP+h2qRS3xIf82DB7/SI22kVUdSd3eG8fjDMxDI/+R9H
SyN6MduyFvGiWN90rS4kV5nYf1GD/ayJspmR7NvSlFEPvUo7HlSi6bNAd3maBqqi
rjPnFpwOZpbCyPFR9g1FzQ+1VUTmr8abTUSYzay61fiJjMA9+L7F1tlnqGfU5g0f
fOExf/CcauIQBEACQNiPVEOp+yf3Nc+TNGgnyYMrP1C09onQXnlH7nbJt8woth2m
pFLk7qS/blw9QaR8JUsOyAH04X2iiGyYFpYMIkn9tAEtBopOefKNk2LPGSSby1Oe
Q+iCgR4ovSYNzbQ2rCUx8Pm4pG/DdLEcY94DUvcI0a9ch2yNXVInT25HILPg8RaD
IGNQnDBNCDaLXwVZuuIjJDQjpCTo5X9q/r0gBB2i/VY0eM5mKxoz32LvdMaORj7U
etCgtgtySUyCg2CxtcjixnhnIlOBmmu4MntrbOt1f/P3i9hg0WTPJPREIXFhTQg9
mmCDETLBeNHH1gAeUTZqD+7pqR6qpejUcpRSofRHranC/wTgfyI/D6TjjcVUyg1g
KTo4OwW2Enz8nS/yR492QrQK5kqBdt5kZvG/ejZw+bPTjohrvaFDHRz4gw04hViL
wEPPEG21j2jiyipTm8sqNao6yPIGsmJxeGdWZa0U8u4w75o28fb/Ckdn3HTeh8+K
vfIWcQq26IX25m5/4SY1V7axsVXG99C9E/aVXziowtoBA4+jjXQjyHTqkLjPY4nH
KJrVsSpjDonxjWLRYRZNNQuy96ZH1PverauVFSUaOMmT42eLNNP2MXEU4i8fjQ8f
ue/cbURpSTbh5Ke7jphFj2xBqJhlo0ud3K0GL5zVRck5D2+GO6v1c5LX/jIJKwma
GbQHySsyQ2oSCZ89FH4kBNMHANhBp22OylMuYKHbmFScGp7XUj393u+OpPXj9d63
+vbuaDfFZG+fGiCp2mPJt5zP3dYFcIZbe6AxXeiLa8k9zLr+o4aPpIWOJmo1pOKi
J+U4L3kxQNBdRxWOkk2dQsh2VZGlF3zhGRp5+z660gjcDYs1FHjVljdm5JK9Zzow
F/0PEJVHx/oIuJTf9au6jAAyBZKIGXELsfamgtK0lrxDTmRLTYl+QudbzAQw5Oka
qd+GykQ5hTV8EjAHxns7d58ErZSZoRgxQD8QUt1Sp7kNbeUnaykvZHH9kxsF9J6z
ikglTOlGWCMnB2Sm+UpuUVQuTKBkIoCVeRBfL6a6B7AUcaTlL2f4vKqpzBlqBUGL
O4iTghofWKj/WRFR8QsWwhOWyiq28rtnCZ5RxtB5lJ0rqZRyahQDDUgmWVW0KYDd
jnRkNDvhynrOwN7whpKWAOwPP0HetKPIRNZ0tf5RAWYFmxv1/A57v5ddgs2ixNuQ
JSIIFdlF2V8V6e9a1XhvlVAce+TSBTWats8nrPZz5DSsyMg4WmMl9tBKofh5dAxU
AlS0MlkA9cNaKzIJ4nrF85QE/2tuDe9g3Lq306Y+08Waqy35HIsb32LMRXla91jl
KPHDyP0K8oe2PZHr0zbRYLiF48W7EJzDpRFW8JODzJzogMTUegm4M1bnYWMooC4G
UJrjJ+ISltgP62swMlbFgnzyQIr5bumZ3MRr3UJfv7dOoCyeSh1mzmaqirhZierr
8MAVM2dh8ntQ0rjHgIr49W9bNTpA0fDBv4ZI7t/eCtBkk5ancFqKqrUDngSbSmPf
+vKLDifr+OdPGZnrpgI0RYPpX8QPwh5GVfg4HqE6QxuWebhymVKtg/0dYQjP73bp
n+fK9Kw8Oo6cqokFGp6DNsQKwuWpDgIu2a4vY8sbFOS6ifJORUrs5vwCtql7LAsq
aUC3oJEYw/XCuzPF5Avi080lvR7gGMN+pRtGdkzpQXcHtHTF5xWzcwBrZYvesdY5
6VNFj6QrK1xu1vOAT3+IbO/Z3BJRxjovJhSNHdeAkb8=
`protect END_PROTECTED
