`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wwxh6OpyngiybvmWe1QT6exP1u1DX0UqfNff6Z4gc1isN2NlWPae3a8YfH3S9n3z
Pk1V3usmpVkYMRIyqkvU94i8T34WZpzSavhmdedN6h5IYA3PY6S27Z00XmDjDoFk
OHoGUeoXcYAVB89Ck5jvcirv68dm8N2HSK3Nqlzbp1LZW7RzxgUrHayZrraonfxP
JyxFvQV3gw+CBJEbFNHUdyRbtiJSilTIMXw14Y8kbpF5DP40+FL5ZmSFRPQuLpEY
DesuR4/pRSYYrfJoDa6f7JMqXX3ByVkvWV4yUSe147g0tp6gb57/D3BO+GJRyw5q
+L6QVMfcb0EwkYaj7Sx0prbi1pWryeHsTpSFEb0WSdcX/wPCFnm2WtucXKZyAEVf
V+CP76HmXyEvcUDqTneOg3rO/LYAA8+DIVEQ6AHN8yrche2yKin39l0o3Qkc3Vl9
w9Rhw0pZBTXSv1fXovzeGFDRiPiQku7FppXjoD+VPHLttY8KT3T0HfehVI4t+4r2
YmOvDdMUfJRB/ZYsD8NyBcalWhfrk5RC0o0jCmD+WSsmHL2TLcQ6ntuBi0A+5cAA
4H2k8/R1cujXs4RNfxX+nLi2tDiYOZAL12B9OIQDhYg=
`protect END_PROTECTED
