`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8PcBetf1h8b3qSy9xVrqydSPIvhbJ+ff/3nKMQVh7446L1pVxizNbOMJTNeaCfsT
iiiFc4jUkepc7+jKg/7pPQ6tBs4n7HjqdKUtumnbYAp3wzvBXBZ2BrBspSaTBa1X
Lgm5puV3jUueHnCWizY0UzNSToh/rY/FIRdHLLS2N0eJeH4BOiOVXtwQ5ZXIcL97
zosXp8DSdvHzRwvk7058uGvDodwW+b7yy1rQQNePa1xbKdzI/yPPrroIGjglXWbo
Tc4cBFZs+lGXgkaQRYCy+2wXBnOfHhfXAiiumeM7zhrVTcAGmKx5wxzWB9N+eE6C
AU/3ffI3lmmThjR49IUqz14j13ZOZJo4Kf0pz0IAdiWkuYnXgHJ4fouLo9XoUDa2
hXGnKtvhWdu/VinwOeeMPPrR0VIvhAA/nkVSYY5jmdyp9jrfeBUQLwoTtTJ+w4ko
ev6O0md9KR0H3tmExHp3CQ==
`protect END_PROTECTED
