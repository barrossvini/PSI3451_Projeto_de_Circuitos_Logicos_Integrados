`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WJLd6utAVupjLQ27BTP8nMEqsTtSQDrAaewGJGX8eAQ2Dxu1rH5Lkoix1Ki+9odO
LhHelEQYqK4WK8pGDg5Wqmglw1icIagxcIHxBepYMLOZBq9a1ze5kSiCAQfyBlTL
q3WHlheO1R1FHKVRmDDgrylGOAdFb63+JEPXI0D07qvT3A4U+0F2U2sZgEulgOkK
QDU5MC7bWNHstUWj0jAnu1QPDWl+KX8DBsGGw8ZfHN+YoL29OStQakR5nLUp7MSI
E0i09hQEqbhovN2F0AdwtOCnQRtC6xXkNbs6rJBoLtCVXTTZx8MGzWA9tPcC3Job
nQw2ldJ3XtMfpnpK20nwRYQ4Kpa1BkOBiGDFA1iZqj9GhdvfDQ9g3j1eayL7lyNc
ljlCZxlDv/WaNnHps4UWU4RuJWmk/0+p1IzgRiyUktggCKeYUx9Y8cKit51Zp6bc
7Drh3n7tHMaInJkS14vLX3CW61QKMm3/iWqmzwwIbl8N8NGaTviB6EqUz+g+Cw3h
51J4kcu/4fsi2Nt0cQz2upqjpx0ql1kUvNJFq3REradjg5LrO7FB6QL5BGE9xI28
Qx2loLPZ4WRDGL/ZGSmK2bCaBMiR4SMRbTvVlYr3aLZmFAzqRgw0cR/j9PyAdfDi
IXJ4mT5IBJx+WYhYzn1cLdxuVGB3Qlcud9NUekCEX0678tFWgnLyozn1CMRDX0LP
bY3a1aP2nQa90hnyZZ4eUA==
`protect END_PROTECTED
