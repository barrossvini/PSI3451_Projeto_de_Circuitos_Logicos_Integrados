`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XmKPrAMDNIn/IsypjHOiIubZAsajvHxx4FqgqjNKAg1WQdDHIcaXZQ/A454FpGms
tI0wdbeken1p2BJio0kHyrMNP9mxZdpqOQp3nIfpq8KycGNJ9d/JB2h8xf+LHC5B
S7VFBSDp78pA6iPZ5Jtj1aXLmzTrUl1gw1hoXtagggPo/FhIdxYGsARNIsXJZjCI
1r5Y9RrePsga7O5wZGnQLeMLIQTcGSTzpT5WN4jVmeO69fzDVM6Ue3NiqQn0meZ7
Yv8oVH6s0pJ0un/hfB+PAvyYZlnfntpx5+mbuB2rHw3YOdaPncGhhp2u2rd8QoPW
57UyAl92veZa5tYe1JVgPlehICmY7Aju7AUC3xLoLnuTYP4CCvohus2H2NIqs5Ya
5LUm/bvJafewHMRd8NcioaNE2pkVFPAj18B6oitHkDaTpeHuAEalwH6mNzbGt21s
4L13rglYf8QLVa0Jv6nEb1r+EtsuK+qEOJKD+CxdGXUek6MShRGTtxLAmcqVwK2l
9Fjg1CT06dcPu+MmsRqx9NipLh8JixBoekP3jbs5v140rn9bENQ1GE8oZHN491w2
4xY08aH22XN4jSC3j4LHGezJJpAkqDx9ZBL/BZkT1iTnxAPx1hH2LUUOXtK5ubCQ
qqVKiaQyE1HOJTBYUzXTW6Vj6L1WGJw+vPi/qk5Gx/LtmJNLG79qrKkfIgIsCaFw
e1Jh+PBpC5oXMitkYcIbUGZkIhW6//PAxxreT3MzcsgIYrl+G+8S+HRRgfBX78DB
tUAXldfZ+hGel2Ei3bbtJ2A4LxPzIu8VMIefdx9yVWE2cl6Q/RdWKkN6z10ZIoF9
YrW9vlI9GH8lVUTy6MEm6V/dr6VKssdf8vn/L1+3UaCpF4T5PhNCWS+rnAQLRmQC
nXs57IhsE98Mn9x8rJ74Zh4J4J3M6Y5c0+7kUXkdzeeUX8YKaUSQBpE1YbvYkKeg
L3QxE0ttDvPrKfCIUtNVACbGQxWcpbF+mRfp+44KMd790NbpB87fkCH6o2ID1vaE
OenE93O837gcJqjLPyWjIyupthCy2D6vHmdZpIldbGwkPyZE+PJaIhcsB3FTUhhx
eFLNvYAtCq0ULVegC3/UJ3tKBFHeD/CBPFqgLVCKZyb06KbSR6drx5ekzjj/oXvn
ZWOFnUwWJHuzP/jPVulayXBDjw7BjvTqLMwM1ZvTjhUsqhU4ma7j/3yqzq7+9bx7
yXfeavDiZYA5jeomLbnnb5Z/CRVuQP/Yqb+veBx+BFcgVD1GFeVjcfj2kTxQA738
SejFB5UBXeIQpIZo1AalIXZc+KS6O768PORZYNcaXU3w/fMig12fY/TR3L9caimg
kUJs1/YuqPieVqm2iEfbjkUvXQO70pwXwcBgoc+m3qSxKyZsOCKPKwzXHRqRjjxp
bZp2YOyn7angV5meAkYt7V3oXJU51V2oKm4nkQLLGCneIXHdKvykom46P5trfxTg
IU94UhCR8VcySPacejbhQ+sMivitx0Umd51NAgLlZ/4KjIMzcaqq4dumzTl8DKgO
v7ES5YnhJZvkGaYOuCYww18/hCVDmK8EsYn1/8/ZvBnJ4Q3HAXILlw/1C4Srtiiw
ao0slZoqzEZfj72T1uiurJIAACnzfaNQQ4cFKwMk0gY0mN7zVf3b5v/nA879aU7/
n5h+njg+oHyB77KTyog9i88kfCssS00sGirEQFXczwF681GKLtR39SqEk+U75S90
bm4aBsyJPZBJulVoYzXfGi2xyPUuxSPdpVjHA4Nxdv11q/fI8dUlYw5W7l44HWoi
No7A4qmTnVxWZRvEzxmmw/FXMTlfUuOjNEs5FXAxe8NFrrEHcM685yio3+K48o8N
yApN28rw2KYwVlWQn8TbThg4xfqPSPjckkqnFQrCvT0xl+NglkU+QTiTnjD/MG4X
5UrYeYYYQkB6KbiB7jYy3k01LbmjRMa8ca8x0/Ih4jwmPi9bzPSUN3OwoiEfexY7
4RVRqKyLbFeDDRY2y2i8vbgzlnIBtvj8g4LUIZYjagcEZayt778T/u29D2kSywoN
UNevRWC5TCZaWW4Jatj5rfdzJs4Oi+lJ1p6Glr+UusymzlUGvj9cb23lXjGrCZP1
1mpzWhficP58FP/tdRpLJaXmtYlGJwHgVMZp3aEdTbHbMqtj/R7MtTYb4pcM9mN1
jeVmnHtRi4oDOlniYZ5W2gftDnmyKizR72nyuTqzcaTsSbnI9tKtkykls80mET6+
RgCEBCmo0G2kXUgQ4cMYWS7Ok9jIvpA0WvozGT5bylQl3ltqTEdYBolK7CrTppVr
lF/1qAINROPKCuRcZaZHupXpwf8zAXqn1tBRPwh4CYbFH61hQQxy2KlfnNK7D1Ms
ST6Ivr3a/+CYaHgTWvxRHO102U+V+N8YldGVjowTFBQSdb/kTafJAzbcPwuATsGb
MrWoH0ZXa20c8atsksJeD1lGwVIkqcE7JyyrU84V8CL/1XTVT+U1yo4oegfFMRvv
p94JbLVyVePth5gRhuuSuc64pGynwW/qnLy6NLapD3/+lkL+dSegtogOtZdxij7b
Wxo1A4s7yV/qz8Is8etzs5d1j1Z1DPpKhHfM4X8UbUmtcUTZl28BgbPdf4nAqNSd
tongyY2LC0jN0GC3eqgYCK+S4kihgDwWpAlI6l+ENQkFQ0sUzeeH6aj2u6RUqAVK
bCFy0g/yu4UARAkMEO7GG6BAOem7HHdWgnXuwS4HB3psjzoYImiVEbXoUWQinEl4
cZNuVJ5VnfjjM2Aa45DH6zX9GHsUY7mvYmaQb2XCsyDVNXCrGb/UycJ9d9lt3QFr
0xs4umwMOtR4/5TbU42dv+cs2RmrQjJyCdtd6tbCdR0Jb1NVG4qdAsF7H+vT9E6O
gUqqQ/+JUgkJqme3TzfXraJAy1XUEWvWi2USJsGqSaNpbpSr3EAgs+uR8WulHb2K
iMh4Xxn/fGp05GKKUfnzCkEoiUXTaDXUqhC0+2RpXGBguwzo483VGfNd/K/oABMt
X8W0VBzKruEnwLQQjacGgNJBq3QWekZIeB7r4B1AzEB4irV7Z+pguxO49MeuESbK
mQHzt6gPCP/ta85oeTQk5ZniF6gkSmb8GrEsk+lf5McdZLqSdBUlDalwS48V9ZLx
GOqo2JPIoGaOXad9ss9kJvGUxKrcNBJMKimtaKu7G0P6PCfeMGPHxzauEq5P+d5W
KmFMLSCAEg5Kvg+vK2WA/GrUbh9Kl3WL/ESEMuNTLQPMxmBbRCSC3W+fNnU4+rql
iwWFXVr3OYN3Vj+0m4Tw6jWGcQz2Zd6oBBGgrpOS8bEkyi5zICSqwIoOE/DfNQJ5
H/oPHX4JzCdmWSWmzagdFy3eLzIKoPG9/Ai9wkjWN49le+tFL5qPbT+QCNI66lAY
mboCYCj4hWNxFI1Amrn0dAZ5HjskP2FMBMWhAaM5Vs8StohSXdBGKOUVPq4hfef8
p6f40fq4Z8/8MJbQxQWaizXTQIufO0BTr6Tndnq55oO/ROXN+NnrLYjkDx6mUPhP
xDMH799rZlRAD0ijVPcZ+o7b4Ne4DsPvy1Ec/97Y6A/T9sb8d3utFdBEcJJYmkrJ
W8jhrl3rmsAyI9lVihy+C41rvHW+z+imb+P8Ee8VSGO72a53hpbkMQYMrSHbPyLH
O9m7XU/i4MI5/jDKoONGrz4YTksrA6Pz3wAeb7l7i7Sqjk/nKKXC4varxQaP7QF0
kEvDVC1lH/SK++1ctlDiz2D5uzQqO8gx/reDLUEX8/5cercdoghyhtzdUJMSYPv/
slp/6zVbG6/tvnSTj8t5cJ00D2bi3CGkqTZXpjNFjA9US2qB97rBpiq66x6GgGmJ
bh/DnfAjonfMGfG4gZGa3JQw0vc+Om2zeyvlggX7MP14rK7yRfD4Qwz8bMCy6fph
KrRx422RoYcIoMEg9PVnjJ5O2b/+YI6PRhjZcvS7ynBQykQiLVsBkndQqAT447lH
0pg6X73CtSN63vw1SgIpvzaG97b7D7O1Kxc2uAiFMqXAG/xJMI36a2P6zHZF4xLM
ESsQlI3LzlVVPbWOZwWz4u8AZq4LKhKFF/4vSTD0x7iBvEmT/BAMXD5EOl1KDnau
DbO6+6YHHV1aXYgChGLzQs5gUc1KN5rn5emNVgUBZg3+pRWHqPHx0E2KzCDoEkeN
AvvvSE57/RraIXgtxDUH5ARmJPjr8r+N6JwbDWEBKdyC13c7b4gwxmOPWCQqTRyT
ImJTdj7SltIOD7pfxcoRQ0vl+PQsn5jy3PTaOEHSFW8TcwxomhldASeL0XfpO2KE
bIyIXUB8t5mgPliuhVi1vpij2HIhVL4F3cpIjYokEQCW9nsnhoeSdLY51FuPAqih
8TBc7T+yS6ctBhz8O6hoU2nUZUYh4gOBwd/yLsYyd2fs4UgXd+4cP/yQKzI1iAjn
gJgwO0EClZXPJUs7k8ZJbDRUwJaek8Ixb+ZNANWufyZFducCOEKotjwf9/f2Qbe3
6awjvrjYkPGTSsL3aOLKJsJpPKDyFw94KjHWdX09pEBT0oik/m9eVjCc7lQlWmEz
NRQpllZp4P4yS/Z1f/h8U7WZ2bBkJwbyNQNWCWoC5m/KuVMQJmnbOm69WC9ecZqV
YZoI9Ke7LymTLhH1/wDgAzdbKCdii2SpaJ+g98Frm4ECk39HsBrlvhLXrLpIe2Nz
Vg7lCPY/nbi+6D8jfxJ98GXJQP18pCfPW4iAZhlYJa8mhEZC6xbaQbR+/pxt8FAj
ZpMnnfLiTbzRahQAXHGpIUGgVwdRJ2xiQgeUlX1U37B6+pq6h3rfBTHv1hLeCOoJ
cT8ZNhYVucNPtXorVh5No/8soGOwHDTJ8IxNYAzbdrCrhTOKAxLm6lAWuw8Lk7lD
btx4211WFMtsnieroMO1GWiy527ei4PSUlLdcXoh+JRJAmVxSVdGBRuNtwiygJXC
4UQDjiDzL1sC57U8NUnPIS0gZo9oOGFItpxOUPzC0DoDInkndwu6ple3N/dprA6s
sAquDqSUFn9QqwbbR4qphXAoAMzhgz9CFRbb7BwhHixPsaVzDHokGDG62ShVp/in
VHBkc1FCvGK6TrfRuoO/h/GZNcSLd47keYOkv0ufRWZ2PFn5zgUwYWOpyxASHOFG
BQeke+fBaldSYYB8mv2c2uE6qE2SUtiJTapMqkiyGBNFyliUORY4ufVbJI3unpqj
QnZwZoKT76ROSBjUcn/M+26CGYGf6IRFGo0GDfKvZXtmyjkLtMjvuzlt9lrQ7Gd0
NyqWnO3dL+jvLfA9W9I/buoXVijVlLpR6CNZXymhFi4PTZJk9VDzSb9gxN0Ws0dL
ayKBRFo6X7nWr6NL8cx3rybyeWM5B72tcCb6n0fcbmzkkk4Zp91HVeDwAXkvFi91
2s54Mca2OSF/qjfRt6SUWjgpM0p6I045KaBh6r8gyM7O4qK7q+tIVAT87R2ItL2y
LMGTpwCLiPjengBm9YE0GmaYa7TIAn1EsCLn6CnxNXTA92H1uu7qXkxw1FtLtPeT
QmoGcxYWkaScz21XTS5MzkhTPbdObGIk0EgQlFV+P7sTcVx4i7pUKa1p8NWJdkk1
o5Oz3szx2TzYhOFtflFK50p8zIzs4ZxhqMiXJdW+y8PaHp6ITd310CdZZI82Y7rx
+6uTt/o2zUa0oyjIYgq2Kg1CZCCVCfGdsLlRBxyCenC6XKssGp0ZoZBA/vDxW9N8
Wv8qNrZdaDDjRgooxab32yo4JbYpvBlC9y6rNgllYBfjjZ0eyRUQGWcKoAfHza60
yKDWY8sgCQMmb8ldqPrB4xxn5LdpWzLko2GFz8PZM2Daz30Atsy9ck2ZVamlaedj
tW2Mwy1Q+WtPPRSPvCSY0503BFMPfU0IWG2jzyOnRzv/RoLyFMoqB3/nEHJ4AMkb
tg7gzY8rNEi0UKRJrIpVtL6v19UpCBOUzcYWXT4wUKnhpSGES8L9mAfGqKlT1NHN
fDLzXye7MtVFhMOUg27bUBjeYCQFDm/pxyeKcjP5aZf1igXQixj9Qppvy3L9stWH
0PL5Lgi+9NY7bXx5ZN3QuvT6VWelXS7h2pbjp7MyoFdKTP9hYEwL5pVz6bTNtICl
KtCjaxaxM6XqMuXJ24cxDvLlLGJCgKaxcjxROKZsc0vkhMqToe40omZCvROprBuM
XVGj1qgi9+Cm4laC92s9LYoK3T46upu9mgjyTNw2xz4Z+WH+KhRxwLbZZMku06FF
Q5z4aaOd+iurG4G99I8D5G7MOQyuFLngfwDok0aqfRXuQQOfh63fqsn2vAFnCTVg
a4+yQjHlLc5bCmwmRO980xs9cvAyl8gN8i/CqtnoN+YN03VWCoyPsfKX8/2PwrUj
jhGlRdnrpZY4hBDdc2WYtvq6HVWHev2MVFNIV2xfc690sVjShmmvNWls1Tzi3ZFp
ugTXhpzJmogIUHknkMd0shb5lZpL+dfkkQS/+JAROaK9Z8s3F1Sl4DSbLwwb7cSi
nbxTRhUebaMmQMRP+2gjkt9bI34Fjv4Od7Aleddxys/IiEc/XDu++I1Asfl3DcfL
avYIWwCBfXCIogNvD4Wb1iBOkvqUQ0Olnz0AQrQaew7ZmAGBECxUB+nL7w6duVu8
ZKbxNb7iv3JctcMqs46jO1OxFKHh+1gIFmrOnkNztEQHeJLRM3aEmxV9RQDlOlzL
USn/LWyObeLtnpFVZzyn0X6iyuVDwP4vcPmC3sux58WynSLpaS7qi/LgC6iwI7hC
+7dM1mCPsf46L4axkd/7TIP99seRZxRTcPg4YDIbr/nOxAezuZDQcSjaTtkY2+l5
qWbLOK03P3wUx+RBi/U0XMHVUDGFy1llOvrAC4Q2jSCP2+uQHfs40fHYCERggyfW
YAa71GjDOvxE179f716QeMXQhkugpW1GEs7mhCvYzBGXJl7sonYl8b6CYedl/yrs
oSle/9ThpuNrk4FSar/Q2w9IszZWdA7VNPYkZH8E4tnQ18H+PvOjIH0/0Ho6H6ex
pthCg4MCL7Vxn6RmVm5KDI9Dq7xGXktoBs4wiWIy/RwqDRGs9Tcywr5LdsvwQfX7
we5QIeD61hrjeFI7Cj/7VN4wAnvSJf48T3GU3UrnBTRWosceUj8GmTDHWFIOHVD/
oN4FzLkdASjnZh5BqL/qgqXM80zFP3hPRYVmFOYnawJ+UnWII+z9iWYuru9eqzTq
h2GthBJyXgW9pJ5HJUXoxKfGPsmwbpbR+XofejOkhpfgETxud3zUq9IzONJcwXVV
WB33I09LrwCFfe3NK/Q6yxChkibLxAdT0Lh6s3AYPVOmUr7JcOostsEIoKrsIO/5
NbNYmm/fhcjbTEgE2jiR4vz2lg5xLnrj66BYQEnkGii0U1wkOzPyU38GUduJCG1J
Z70rGF2NZr6en0Kty9Ccq6BD6XfvEkKwVnKSvaziCOPSECzIaUXOUJva7ehPClPD
PJTFMYTPInX1axCvKAwuG3Ve5xLqMCkoox4Oz7b2Lg1XlZsDr5KqXkvPQ3oPok0S
k3/7bgdoHJ3fM6vcSSDjsZP3H5N68g0kOeNdskDEpFdPrW2RRzEbj9Cx517jBxTt
jUksmrIHddG4VDWherAzBq1jmX4lGxPAOHnk6fCJh7Dwh39txIQMOLOKcv446Uqf
4bDqnEo4T+b/EgJvtdb2LSjcfUFK0Al24IXXTxY4MMuPjCdxlJ1Gzudgtj27zNnN
lA27fTpnL/Uh4QkLMa+u2Ht/PukBap7XJoMe9zjUPGsFjZHJFumaFFhRd9p3QWzx
eIUhSzfEES+lpk/zthPmGZ7RUQ4H8RcCihIGnSV37XXEMLnInfOWduzFTU35hI1A
p5umwUMCjsv65camQPmRfJ6+6jV9JQiPfIfatSHiacbB/qaTEjnNvSB8440cBdvV
ExWsDqZonpUPxyOZlESWNyUxC6IBvRbJpJAXipMT+j41V3B78vYRNFm6kpBPaM2y
uf5TM3q+xqSoeZHI22QSiKWXztcY67IjW59EMyCLmYr1WnE1ZRKnNwVVnZm+sked
6cawQ7oegIlmHVgJflcO+mCIkBPUts5naaqhx1HQuOU9t0vusVG5Ijy59MUwoxek
HDC04PVgSMYgvYaaUvIqxchexrOrKuZ8+WWkUTDKfjBIDTDST8R3mJBnAUp8sYwA
VLGFJEWIS7txy4N4tDbNzURo33Br3zUECYev/A2yP97ic+xAAZ4NbQXMSEmd41DV
X0WPxHramg9DePwFgyVCs76CkWDBHw5fmESWh2N5PhQRrg2K9OsZMazYZw2TG/Zr
6msrH2t+gv/mBmWkmaOYuKUnI6En0UrIdpBm4fHl6y37w2YB6YY6EUziapBpHkoR
rnexZ21fyhfGV/zgOpKb8Eisac4Np/NFFLzPcJAA1uTmywsZtlluNIExr/joawdK
gdEHYXrrS44d+LMf4MJ19wRFt/EL6XQ6U1DmAKTR0ChzvuY92tOuyZiraj3XA66H
b4C3THWkk8A9Y00rxfr/ozM/3XnOVJtvk9m1coUh6A7Y1vKd+WBBetoQC6/YL5tl
QYLMjboY4VSSVagFQDpFFWlupvqIs9jIIZUqK8Rj6UYtHUcWOw/Ys5W4r8SXD38F
pm4RVYfqiqRh4kcKMEM9QXWLPvsPN9FABuLPj1kaG7Ufn2Pj53im53ZlAsQjQpwv
37SDCLHaozuDIZ5N3FSieR6mil0k8MOJrclEhfLXoS/cC6+5ZEbxtJ435RTES+Z+
+Zj7gePJQ0zKaQ5VB4yENmpAO2VgvbT/ESRwBEsaZceYLmjVTsO0jNefCHOiCBO+
bmii0898ixp73JkMRAWonVbh2F8wKfJnZ3vs1Qt04qmKBY4wc+e8tLr6u5tTH1cv
hdQhpVwY4+1OvAAqP9LCUnik5OBMB3mLuYQpD1EsPvrZ083JLoWKnHRTML4tzi5w
mwZfBoScPWp5RMyQojxGiJCXAiwD0JFC+LvbjDVL/1jCCRMGwfAQ8RI2f5mpOrhb
vfiM8H60l5+8zrHpuIFU8iUN+kIWz3mX5DpEab9h/1DZ6C6ZbCCTUjAF58By+Ozs
KooxCqrAa9pX4GxjPWBacvYGQGGnZdlQK0LmuQ/46q+kJcHcRW1W72q3TMsPVgcn
f+c9cuMrGDWeq/PNr8GznAlu5s9dwZkmzqiMh0dcx/SywTCAMg5gULT+Mie4T5tZ
dSD3dfOnxE9IE71URAYrOpYMVkvgPYGUlMopI5jJaUAW6j8teRGR1hswV5wjviSK
azVYgmXOEETgm9LVMQyoRcGQx7cKcCS8DNQ6bxpOKLU3cAZFZx6fy7S07C5BbkLP
iIrKCiquhK8OVAZwac7C35N0XTpoZLLe1lWEQbrLtf0F3GTDP+LbvC7ga+Nbf0XP
T/k9pt8y8pJBoY82XMBLgBxwdnS1teTy1s9h5UwEp2nCx3IZi2XeM28Y/BfN8QLZ
/I8rawZeDYl0ffjzr83ovOgTJTTjtJSEVwxI1mjR1FVsvGldzmRtEwOpYbRjeIjd
PZ7xiOCgXkIznGNY8D3CykNHKgsNZM3KpZZHjK4s0ipvBtMJtkp+M78v7Mmfv+eG
PQMjmMG7pGzjZS6lDLE0QdnB3tfBNDp61+9v001xlx5fN8aLyx4sEGcUxpg9AuqL
sEj5ClUFxXSgas9mR1t5uQwsw5Tr0F/hv1BluS344B7Z/Ani+H5dL6M0lCcVHzh8
7QbDxkUIxc7jhL4k8ZTD0/oEVh1Gas0iEFnSf8KwAYce5GWCDKcWYRDtZRPVWGO6
e/t/BpoVvuqHeTJNWctUZg7ZhtyalpXgiP4Witqi/lwT/3i6Z547RRaqcvzzaBc+
BDr44dihmVFSGxx5WRiUSCGPngwigkYH+QuGsVB8XmL11lAGPFOfZsR/Akv9TjYj
z6f1Q/lp0vlrBuM2aZcvs8S1uaV8DlDAWVWGL3+x9p36n0TXRIrDZJ+L0N6gnmr0
kMf9mZlWBsLc1Lynzzw8wCqRYoLCQyINj81Y32AfCTmz1Xc+VyvZxhVGya8w4002
WaR0yJuKhTg4ee0LDe0S2RI+wtw5hdkRmqHMXcguugWLaARn2arA2VxHGid50z7Z
Bymz0Nyoh0JE6c20Zd+/aqVYrSe4t0FqKAkQp23rBlNMsqbcsLpSVdpDgV1WHfNY
WnJiJfN7Warn7tlIAeleOziGLn+obkN//3YSLMlTMWJJUKi5GZPXt+77szpcRADi
R5JDfCCt/J7S+RYNgjS98UdnTCuczLZuzoK6ZFhFnel91pxIJDP4GAONGC8Opgs6
wtmnNh1CD3ajSCtgw/QOfd5N5lJW5MgPo/HfVc/iRuZUpoVQv8b7fMdQ/yoSlMNB
mhTJ6zN4rhtLmWJSAdo2TBhDeOfA44OAmw1vO3e+HcVBncUEdOU4b1BHqYYxCvyb
KhGh1gM/bbJ6cpBb9QAIBtp1QnRjWDqhV+eUdn79WplS6blIjCoG+m8K77VSeOan
muXvn2WA/y+GAHD++r2adxXknJDGasRNCV9urlSijybrXicg/4hhhUSI6tF0GY2a
8vhx2xvAlyLQ9Ev8gWbUqv1U6eQD/NL7U3NvL3kIuZ2WV/21y0odJVUp7NFKa1Mi
F29X6312UDMH/Xt5a9JRvYnq7hclSvllfsix7JPGxtTLYY71y+2as/+sA27g2xVO
lzpUp2tuq7LaO/8UdB3vFNTOknUId8l4x5aXnTQGZojo1rJTiBNT/DrCaml/QtgD
0uGDAbTxloh3I80U2OZ5q3B75/vctrKwOuIIWr4T2cx9ZCdiFA9D9y4t8RUYpf3X
nLp/2s59wkPUU8NlzUjNfVkgFcA7tHijNGCZrP6qxYC9FxEQN8tke5t+xGj1Utwm
mUg1qG6ma1by2xNriOBPmJ81e79gQ/2eE3vcTyZwIq7QrijwTlghaHqiSprUGQsy
44qYFmLhw+QdtQ0Rnm2DufSjFGQm+hQAlGS1tlZeDWowAtNLWTlqXFyfEsko3KBS
eTdA+tMya84JyZkeQnZ7VXFtK/uKHiW0DVZWnIes23OH1p04TTjkSXm7V1fsa9az
5OGHdif9rjjiBGM2m1oRBmGeZ3hoUtChPOnAFHgM8rYhLWrhKhC7eZNmyWi9IbAV
Ypv9/BVkmobHUYamW3iGUZTUvky68klkkDNH00gSy3m2VmVw2H4tW89TVvHin3ha
H5cfSSTmmzikEHi6fTZrcspOpGFt3MdCTVtoQLOj1vlM4iF9a8Xp42vXoYzrK/gf
1M//ymix90djuy+mnbd/N6ofYlfUIH0xId2pwngzpvTdUGi+YCu3J4muBOLr9n34
3Wc+lDfqjkQMlHpUzrhmIrZyw2ouQO28eje+eRiVNCBd2MLeCNPz4dH3VayPrGIt
fj69Z+fHtqgBPrJKTeHFljnP/5KTyaIqJrOIKzaAGbqtbBws97SlfEN+Vs9OaQkm
dTxYOszthw+/tMhNgu/jjHW2NoHSs+xkY4fJu+DjgyLE9K86u5HHcobETFnb9zyh
8CJeE4PrkaEi6UR1KvnWraEoDgTpdrG9iu6B1e4uMcM+BK6g+yfiSExKiOBNhJ29
2A/6QBrpY8ZfH9+xwTxxMB5W3kf/2j6EYJgrYXQA7tHJHyKpOPGNoo2b5sgaUiR5
syR36rId7E1HzhLex45k28EdUw2QgfPWtCeKQT5mswz+KCHopkzgqv33WPda10zR
p36J9BFj+X9bH4kDGlTfEcJDJK6pzJv0fYeTNTO/89NLvCZrAV4Wk+LRXSN9+R+0
B8dCQyQa7AlRUu3ZRLHpC11j+fm0BWmTNl+uGvnCUm+vIpbqh3yX9hTgdEuVzoDy
akLiMkWQYVtZ6avTGgDHgN7vQIJNSv5cJgJj7Q2drehcCuHQdhstcyPL5MKcR9lL
BFAnB6WUvBqBtJepk1RaSE0AtXoNjoqhA422ZDpTJcx2mqRH1Nx3i9tVaFR6pR8B
q4i+pbiF75lFlanNCfv/6JkpaNZDLb2G60pmkQBTQY8TrhpVKNR9NkV6x59q8QvO
izqgje/l/3jhOElhJZRs/n9ahviSIKBCLPHia/gTsnOzxrUDfvr/3XLPErbXA1Ey
5r6xnEV7S1bQQ3vLynLxTHsYOFtGPoWdBLhc2u5yj6RHpaLShuCE9InXTFdLWplO
NDYEWFT5B1NYzS3v4nw2YZ/Sx4cM0r/8f68n3ptGyt7wJ+7UaQS9+O/m54hvui+x
3kBxMzmIARooxqJ56QT7wSSYGy+h1eWthEpFBGL14O/FyXXAMTGzhLn+HdpjahQW
isoFH+KZ39GAUX2YsnpPR/932wC66OCHdUZN/eb8ZRWevqKo4mean8kTE8VcZoPs
4c+grqvHD8TH8FpdK/P1m9IRSneZxlfFcB0jNpwjUEYBuUgBBh+MPSJIAdsPORph
mz+Byd+JkdKddaqAXKfXxwin57FfUsltUrlC3aSUyWI51RaoGvGHJ53eSDdQzier
DyikHo/r491f88A5H3Hn1AJVG+NM40RDthE91OylCz/2tXVM5A2VCvEay1XtM4BQ
/1HdVplJFMl0lYMPHrTJyVJQWlVHj2b7I77qzl/UJ0/1cee6yh6STRXHToZg+p4s
IsLE8rQL9lJyB3hF/4/zDcwU1jBxyK7Ho7D9t/l5rL776KdLm+T4flzFRvoU/Xdo
JcfG+d7Rn7NHe5GbILYDibXYKnduHRf9POIeYKLH9FLry1MH4lgXJQw+BTaAdphA
FNjhe+McxcJCG1HL4kO0+crb3CRmd0BY3oTmc0h3BE6nkMBAQsB7CXCG/UrLU//O
LURCThsIYjDipvuikgCaGjylIJBh1n5GHOGxccfbHym8JYjFuL2ZXj+5G6RyJc1y
mpYoQr0r+TmWjQ3DFEljUaqZyaK/eNUHrmIrC2H9tS7n2n732K8r5Ig6QD19Q6KY
4l2+eQw6vI9jc5h+q70xTrTeZUYqv0j+mp7qeKBm5TZMO4WmmXqrmSC6vRHSoHJ7
yK7fh5CVswe6G25bzXb51pK4xTaMENxot0b8wu71CyfRo8Nl0ZJtHut3h5S8yZii
grRfsoBDaOnS83XnoaaFbmeAk/J2A7WYUhrZZpI9+0CH6O3/zC93CYes0D2fuiir
MRYFtQk6gMOBFpn7mhnxTyHrsBlEuLFtiE//vQlWhi4J3VuePEaMVMXYX7jbaz1F
/7ioPyymikcBOLHhwSaypF0tWNguyEgE5h82vFpdip7Nvqt0pwOy+nkXKx5VRetn
kKd74bU+hT0P+3d4Smbq7vNlmayyH1lPZjbY8Bs97dyGKpFFkh81YOk/EPZwDcHc
d7d8ZpCKwan5A8Z19tdHfYoNSJ4hSca0PrP58ZH77yJD/T6VqnOAfDqjHdaiflYl
FJBCR0IhlnhcMbKwRd09sw==
`protect END_PROTECTED
