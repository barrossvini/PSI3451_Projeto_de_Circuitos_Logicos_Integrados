`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g86FL4blg/VXA024jnzCjLvXXWsxYCpnG1/6cqEV05TJnRyLaJx1R2gA+7NGiAHF
IV2W4WdrxGFsxFrI7fWEEakN87c3UBeLAvOm1C46nW2QDwAFbB+yWFsrVXk83kY9
R5BV55he49mz0VdK0vyMHOhykIWPbqI1R8DLIHRVliGExYf22/nTxD2cAMYLIV0G
+5EkgibujWTnwahuvMwSErqmEmo+FJ9A8YrXylraMpPmCAGak/2TxFoHlyc+9cX6
6qdDAnYkisr1GeTB7mdt4nhPMRBzcL/jUXSN4bS5k0fREXF5iWiCi2sjdgxvNbDl
fg8e/UpiU0KiCenCumIhGsp/OZoty8ozOosJJImmcwgTqH/MbQBn3YDfKFd6ZFzp
I6eLzvcn+Fm7k6/M1xowOX+6NBW0xqQHKBfbb2TmaEgp7+qzgXL3y64XkDvpDiBW
FX1tuG4M+rxpuHsX7DWL9lVkFmCwlkG6x0K+b/6Bjm8DfEK4NUCgK7rwtG1CzO7Q
`protect END_PROTECTED
