`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X4dJY/nFXvD1ja7Dehp9uXMm9kM4dD2/oF4wGevBAWZX5D3HR1hB5wq29XvPt2Zz
qKu9LEKdKMDDZG3psYvGBv44Op0afRHpDVMCJtMOfrtwhU9uQjiRdV20U0/tWAzg
faXBei3Z5Q67CtTGSaN4+CdZG4crh7aGwRSxLzaJ2RA5b0v30By7Gk5dbVsZZgPk
qSxbpEaqLvSLnOx0cciIwrjFHwl5S7VJR/wQwNuQxnnX/rMd5w/hCuouYCMQzC+L
sWoGxLKebT878GF7LlDBzx8qYDNFBRJPUKbBtJfoTbZ0mSm2KD70X4XjMODW+7N5
uI+lu3GAjHNpeB8s1sdIosPWfsj/+VnHB1VUxusjxnte89AhsfZPQwVAGOz5HeQu
Y5oYIZLhVIQNcXYLaMdmgZXfWPHbVTDqzHSPHCWZj8Gi3hBefdbti8xRLVRjiGbh
p7zGhyCKmgK3sseqn2O/VRH7tZQU+H3Zn8ZdGFKwAXrPvrjsslg26HGQi5IxCzuA
5YZeKXVa3qDXyO6qpj03SmXrN8BCM9S6sXmqlD2v8OvO+p97kB4AN+BC4LLq2zxa
t4ySyP6aQ9XYnsXZXXmsWg5aUizell10gHA3j85BIIaK+osG7yGW7H6UaQZMh9LT
LNvU4y/ATfmlUnAkrIBUjdf7MGRyTHeM1T7xAf8E2zYouFNUNbDlRD4jrl9Inift
37l2b+uwyONi7CdsfDzx+fyg4tLzrR+5aQw1OtTyLWOx6Ql2RSsHVKLVgzRraYIj
1j21wmS6qV8Xg+IjGWphC2Sq8TyGGgg4SevoOgIYwBormT8uDiijPE73uPInF0+5
NPlsqRlOdm1nRe/E2DA/dETfIWhlSz17lmCHWDVOWWVjH2ViVUXkKmJUmNRXvz9k
hflSPc/VUxMZ0KcsjVFSt227lY5A+aIr7t3ZHN3g0j2/TVOjTwEBDU9FPne6DQ+i
lZGckAXQGGhF+cEZaJ5MQQp3sWaqR0jQ9BECPum7rAXVW0geTtNrjn31pIaNXiKn
cEpRcjoSycSGpkWlXPazDNNYXv50rzef1NKmc1epBQChY5dSsVcmiGHYxzb1Ic4D
I63duAlsLt9o9KcnVU3nOZgdKIz8WyO9seLJxFUycGb7M7z89NFQh6s+aTKucwzU
VlWbqi/DxaUyXHxAGMiUBGc78ww3AfP2fDcUfQaq37rULHbW0Q3EQMi+VGh/hUHg
u0n5WDAvBgWWxra16pvrTqwZQZrJMssMGBFD4BeHBBcsa74qLx0kJ1Z7j87r3v9q
63cvKurpgqokfe+UZYa+q4oW6lLa5ul34lxHPdLj0uEwzzJvajWmVF4pAIk2xh3Y
PNSMQkrfb0qZD76PEcEwsI3mDHVH6OoUMPcE2vRK8E0jTc4+McvLilHlE8t87Ito
eueQkyr7RNQX72KdFpTI1s0J1Ub+Edf/BHV6UE95Pikl/SD4myg3f/2mT+1KWppI
M68UblZ3twT4ezVAlw5OS1+T5OTe4IZD4KPJU40OYO7K0tPmNpfGpfijyDhGbcek
wZvhIjd0YriYcmzH4t49FQ1fo4QxpFYe+YiAEcVlGhTZVyx3v4eNEFNmnSf4vnDw
vx8eIOinrmvaAvidUoAZzqjS4n1kFCMMyG0L2csWijWTkO63G4ijncfczgPIwvgW
4IscmsyoQYwL7bhj/7sojmG3NHsHfsAdAILfqkTCq5V3JzyaSNTNRndjQTw9PDMW
zwcodkLx23kqlev/x5xzSmi5gLRcUpjnfrgRztq5nmo+TkajYFQIabinUa4zneMl
3eqrwxDW/sEZc4fg5g7ygaLWMQFFOoQFclnFh6gTv+PswfQZzuAw9gsExYewaM+v
DMZd2NDt/9t6YDLKY2KYJy5lzA7ajup3EaOfW3Dm9MsjIm5yaLtq2xjMpIuUsfET
47x0vByWxwXcB3kpM/TzQoIJJ7AvQjphWJMAdq3dbBovhF46BmxRZS1S69TjNylO
vj/haTUIy1BSCBnMgkf6ZjZv058CZEQ220XJev1eazKNqWCu0/uC844PgGkQC8TY
uFfPer7wTFxz+GzW61hexhHk1JtyLeY3zzhl2cjzMMImdzW4/F4PLL8JcA2T5GUP
lQFrPwtrc7dIUFe1P7AVAoodm8QXxjp8pj7fGN3eCl9q/rH0CnUrTpKEbMp6+1AG
vEwDBxtVjP4w5g72eAQtBK8K9qWt4dW0+HukjtfbOrw3igDW38U8Xh3WkMEp381k
RCwWtdvlH5zI+84/8NXpunW8vWod21gNhUVuJT5HhAy/Q23i5EV1+vSHyTArMIKy
3s/rYVVfpNntJkgJ8lBotLMvo9BQL8byXENoAOv06/3pPc637REK+91IBgsB0i/D
oSmif7e3xsmQAxQhZinaqQON6awp0dZ6DdwWPno6IyVucxtqp7Rhq9kbwEU7jwrv
9ecuCScDLrERTtupQUUQZFP34OMnYNcIl8CrKl24SWskyxQG41eovyI9ni1Sj+IC
QxGVDDTvtAqPIMnu/+yRQ6h1lWbuC7EyiLsXAYKJ1Zp2QlMTsN7M4TWmuBgyaGtI
TH131bjdGpGzOsB2bPz1R45cPmQRVfcD1G/wJ4JK/n4Rby9Nan4ajClHIcA1sg8B
ukDeWiAmDpr+InVfFW6ZoryHuX6b5PuQsyMExuLoRkyWXabFmCNoF3rAo+YhhRmN
xVKetOckF8Gkd21pqozBuevXt9tm9ENGi8oMkzJW1fK0WXJGo/+PWvU/LcBCJVBM
ZJ98zDpOkm+HjJFOAwmJkJP223e1FXHXJgEuCJKNXOPpy0aKzRAnKl7khOSWKwaS
COvew7X9BGhyx4aUqElFpTK6wm4NEx8HkaLePXL9AsUcGl9+hS91h4la95QJj6Bk
a5IhNX5FReRgRSv2WD6p7WKOtLpIeQnnK8WDMYFSY9rDNLSloi0fKkG8SmCkk3Bm
yX1qC2evzIbIjS9Pji+AHC4pai2YOMef0kwNlLFcVerbUM/UlT2Mk6PYUzWCRu6W
3qepNVJKMeDDfYDgUfiKah38D1jYI7XliDNCwFMWxXQ8LXigxSgyL6rHevkqBx5e
/bYJeAxIqCVOqRd0nAhZJND0jcpWw/weoODC26bm9u1fELbTPpLLN6XcPynGVRWs
danGqjCgI6Oz7y93KRxZSm3hnmsVYaSG+HXp6f19ZjuhnJPUyEg5dKLgDT5EfmXk
iiyfL7hrjR9Z1PFKOR6g3D+0i59X3Y6I08lXel9cLt2a1B5d8ZMvXglgCLEFxr6o
9L3QpgKlXUDwmLLugR3cBSNTtmVgYdy4DNliTFxgQQxq91boaNTB6afvIbV92jbQ
mlw9aXMAG5/RhIJWoppxTC0lyfW1FMkWV7Wr49NE7bUBjKzMBWb9l5+SAj8PYC8A
aFKMgwdm/8xuKvtsdqxqwIq+nkHKmh7xzl56Gg2WTrpPOAoWf38QIQRHAiziEA5H
qe52+Ke48rUWD+IUvrAhztIKrOJtqz87hVxnHAAmGBbwh1mGRhv5yb3acC1pJ1uK
ZlbgTgdXlb3VrQPEXPnR7NPcGgKzFJZJSY/kCjf0fbNchPJQWMO8fcnh8ycsnzuL
gqjF+jgv+bHRemdRH6CTpXFCCZh9qqRyVHyLKwMXvkw=
`protect END_PROTECTED
