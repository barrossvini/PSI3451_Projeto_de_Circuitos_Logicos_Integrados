`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5HU6fHNNuob7wqbtblQFvspbsBoMK7y4uKWL044xXECX8mpalJSymiWve5M18Bez
qPC/DtWBG0j2ILhez6gVGQlr6efsLxMIqkDrYlXnSIw+Txz7YUwjnEN/NTBsCrjm
8WzBcCzmg+At0Ro/P4/ot9eNTd+n2Uf1FLwLrregyeTISNort+0vR4SNBqf7rJNZ
LAcF2Jysg/opvOBx1zeiddovTG7ISQcp1+E09hq3kX5WGRkpTFCvKYKKX3SsTo2v
hoTavxufNL4KRfzMCBK+a0RKL26cMK+9OWY1gBBXiXIQsqqS0RPAAelTTGuGbWR4
6xIqCSkVjhqMtIUiHyGOZHw2+QVGw1YjzM4oDKWu5CYxobEjM6A1v0nRVIq0IQNS
LhAWOwHcPheNLxbSTjqMW997oUO3HpuI+qwAa1jhyifp7Hn3pMSwS4YGxlIXlc0m
lXX5KmqAvDbeHSwrKr7qCPukd6XNH/TWDwL7XSidKtFwnCW/9x1ta2iAfFCxc1gK
SxYofjiMEToPcAvBGNmW/kz/XPUxVOfTQEDzqfejX3zgj6m9I5o+7RoV6L7neVqJ
Z8MXKuTC0btXa3GtDwiZt2qYiGQOsenD+il+PIB6v8G12jLcO5YaEsDgH179wXZ3
L9iMInMjPnVuNdwkrY7wACzRUfpvPc3wgIe7OcV5jjWaeRWpFK+9f/UBsmEl0Xda
sSvoH2zWw5hZf9onT1VtQk82OfaY1EU22eK2DJSdo4shM8EugLfUhTwmpZcoWVgm
Kx4orX7pU6bm/6KcBVjdsDADtzObLkVevBc2oPXfJ1Sebg1PQPB6eFB4ZsmEsNSB
MR43PLIIsk1X/Fjiflxw525P6rw7T6rnS34fF7fUQQ4=
`protect END_PROTECTED
