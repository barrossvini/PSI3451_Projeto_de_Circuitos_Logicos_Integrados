`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cx7TdrDAgov4f8tJJYLFNLjz55Tz0C/Sipf1wf9vbe3jV+1TVC92S06kmULCsBTB
n8lhK7Isep+9IbkMGuVy6l+g446lkoet/e70+D8th2ZB7dwg7GZZK4VZu96nFjmu
aGdaMe/Lq/AV4vMRgXXZj4cCG0iD4kdEcDausO7K/luyyyUdODIHSq44DiNiRNm1
XswAHoHR8heOfu38Pf84+LLuTnWN4+WO8caAjU1eNZME19ckfRJdPtgOEAc/bURE
oBREyXUOqr+VDDplT3ryKx0E+exdDoT+WBaMDFUnYm/06+5IeNfAG73vIE1/HhZP
PMvkpAoUgKgzaxgm91PCNdP3YMgY+SxIpsLCBjo9GZKAdHmRCr1vzG88x4/9E2yG
G6qmxv1hKEmzE5R8sBkuHcVGMbhppYf63fZQa36xuuxHd6+SlFVi8lV1V6ycglgI
Wqh14eYlP77kryYkQxZMmlyyrIdR4EgEcO9xvihP+iE=
`protect END_PROTECTED
