`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vF1fL9O5mhLq1frY7tYJBkHy0H/Lsag6xQ9j1pdsvQXr2pq/BRcDynNKeDrJ/rHr
DE4PWek9l89BU5hkus6pYtJmKkmAUJAYVCvBgNiJzfR5Vxc2XaF+CBntmarwB8zy
qpfAYJ0zvnkLDgKNPdohhwEVC2MTsGePm9EKebY/N9a97Ct2dNy+3JK7iPusTHK1
xO28T98QICkcuN7fsB6ukaW7pRBNu2U7KbdaHuY3x+DHx7osARRN8AQ5gD6Tk/Wu
T3RmQmX1YiVZFdtuOUT0yX+fiyIuuqJWgfEIBnvQLIiZL/n3PPaZYdR5B4D4t0v5
itUMfIHHWBt3X8HP/H6yf00gzTLR9AVzp70byMq1hlMvODYm5r6rJzZlWaM2bYZu
1RVKSaC20owdapJGyo474cTmP+uiqU+eMDHSKjyY58FES+tb180WMilNNF1d2Ito
zyn6RzZw1MGN/lhriDhLAxhtkqn6p6vbTLeBfoagTsQSTB+beNc7NMduCZ8VTris
eLb8PbfLVQajDhQACgkM9TDRGBjHchVvgyQC1CnEIW+YGkJqEyFa5Opw+2Wxx9jE
/1vjkgOf+y6TRwwSNAHHv55pcB5S3B3TkcXWC+JP6HmuDrrq56fyEqlqO/ZvAGLp
UCZM/VnDnoek7qzBYgIPbByBi+3keYlBM8EXoHlhOJmQFnnlt3lGBn3vsOc2WM8Z
zqFDdppdACexdgQ/npG9dGt+F8vNlXGIzt8RV3zdHfza4fo28XQcn8MQLqcSeWyG
733+eT7iG4IOOlSEYeAK/ejJaxCF9kTZ3Ymia7cpoq/tD+g8xkh+xmEx74mRRnTz
kwotvhaTWijw5K6kPkoxTD2QwH7W89PhgZuvoaW2WuJR4gIS8PBisn61m1LNljKy
iqoNNr1BIL38XhMdDfzlyH+2ehXljXb1V13xbBzUcaPoW7/FFyFKG+ohV0jqZDcW
7AQkWmahdBr4hdzN7GiJ1TT7AwjLLziBkEy3LFKwK2G+w0JeWWTZjfEP7A66skxY
YMcjduwAxgl0ieVTUdIOK2t/RJs5av+irgaygKKSf/b0rE1lcpQBMpUbws/vizCw
BkPREb2YVH3HJr0SV3mE80RYo4c7qNXAshrjF8zmpmU/XgHMlLNP1XzihyDlnPom
OecU4iZc0EYTVjtURciJ25XfVElXiCcWqXwwnBLbQDHVIVS898yTyQTIjiSVFItc
exBd2SGDjuw4USd5EnO+TphB5Hb740qPogbTs5LhG3RYixKygPXbhPrVLfc0QUs0
zdK26/AMKvKJsQyh+pN9EFF2rxi1nHYsUiYBZQErv/NpN/IdZ5+DmaDPbHqMq5Km
t1cgpe3TSHnbumpLnFmoXkFcerlPv9j0ZP44ToZvSeRO3a7rvaSbFhqqRni6mcCU
5aNHjRbm94AiD/yrly72GpPD0083+MLzYCEdcU7DDWvNscJzpAbvRe1/RKkW4Qva
YqKHzVum13fH3EdsQT9udL903xECLQ2KBN2RFISxds3V5VfVCJ4/Ohsa08zVaFA8
35T+zKmbToaI8EoqWVusip91r73JlaPIqWzovi2rEDg1ExeRqfkfRXInRR6eAFmY
KBn8tGsOCeRbcVKlFnh1J8ZGgtMHsE5zT6WfRj9HXRD7st4r4R046NH2CyqnJbSz
AyR8RgNXK3Y0XaqZfh8uY5eRhKum4ItxDJUoDeFB3vD4aGpTMgp9mv59AKy/wOIt
GFF/LMMZnQZFxM/qBtb0qFTG4K4iJjBMlbFhAz+Zb9MwmLl7EOpfsqX0AX6d0Lhe
zBY2VRGHS0cLokreCm5T5skPnjZwbMMXwEeDwPvZSp5n6o94cain0XhMEjXt2S/m
3mZ49zt4E/klwJELpyszN4xBjvGU2AsKjK3hD+f6qMn9Mr2ZaWHQq0GjatZDorHj
FBzzuWg65Tf2E3GTvBUSW/LPV4/eJjc05LzGKDFRzvq96yAQlV95PY8nef2jXpgX
1v171XDCx7M4L1mSxDOhVN9FqKYQK/UF/1Z/x8yws200Xby3zRzasYtXXN6bkc6a
t+eJ45TC/irjP+Tmsh0tdVNmS6/xyuMN7mNscsCrW89k5r9/ecPQL38GIv2xxOca
XlMlJ9DvnmEKWJIzw9jFYv+7EOkCeGsQ7U21SWOyUFDasCNftRpp7MKUT+RT9lRe
b08MpYhw382eWtDxJ3opd7LwIbj08PIJKCAblfJC4izBPgE80nrep3OYOZvp8J0K
yFBBswBR7CIjMD0ZKx3f4Bi6XlAsgNUB2ZpDPQfH07b746VrxnK+Mbio4qIikNSE
P+HSarjQAhh7xN35sERwg9uRgKcvtKdHOwJOqn/Ln6atEBBHMAgWGRqnRMqKh/N6
jRFPmqB8VgA9DUIfsxgfN0c9QMWtxCdHmefem6pbayg2aiKw3sS5Q68VKsV6XfdP
HiEmN097qsIUBgrE7lgLhaukbWhUDGI7+TkNWkoaPpWXcDRMtmU2AFWuTY/W/png
kKnLcW1IhQIIO/F6HYBZt2A/E1RxYdrJvwevBAbvj2wVb5GK355FgIGbrMTEKKrj
bJF6NmLEnQmta54v9neII2GwDqgO4XIC2OlJWSL3EwLqMnq4Tev9Ch1J/Z9bykDv
K7rBw/fEaIxuKZTbpYFSHyaJtuk8zUdhugmYLochINA5CV08VtiSTZhKaVqYViqM
hlHNa1sWcO2zlOTP6UHLd5O/KDB7fPqwLb7yXTvaRyt2RGlRhWfV5Jmp+Q03vxQU
dWya9K10+GP9EWarObRq3VD3zZp80wPOxtTh7q8RXJZLOi/2bzAmqoClNA2dXJwk
V4vZq8d/zy2Kxl+CG19YaQKn5lJvwc6PQsoQkYO6dH89jflKYeRzDKjd4nvPAVUJ
CDMLBwu3gf224dgZiKqAgNn/GDfeOm3gfystLJgKbAszwvKYRW1ivyQjp/L1cJ4H
AP1esvd3PKGfxuRGWviGy56ttQe5MuQetYIIrTOO7aDBTPH/WQX2ljD4E+asT4yL
JN0+oNOGEPH5AhOnAg9oQ7lC5MZvRYkcZKCD64LwC5rybzo3t3NQ3m5H08vL8THQ
n4le++dEqjSvQYL5xgyb0eIZVCo6nGZRfiwAo651J7N3LlmYp/PDve33kmYEVViU
xqIHH0Q6gsbh3mrfJrJ4BdR5GM1RnvUAHwPh4e8/uCdCPbZ2GCmq6XaPTXZh1cIx
tDYyJEEt+nNdkELgn+Lq4kxV1QmBedLOkrHYC0REwvH6c+FGFgIStmTV2qfrG3VA
U2md+sodDwM8C+GNHV2eUjjqWo3edSS1xOWXZnQwtdlCBnOwncBK79FfVeh4H25H
WcrVi7NGsTBfdqKuoBDvWrLRMIbc8u4pRi1A29OcCNwVbHGyvgmb3smg22DdQRRu
0E/AThhbZcOjEMv4aU9hDNGSXdNtrFkHqI3Y3xYFTiYVvIJNeMIFNiVrOblq4bqN
W5QfZgPu1FbmRPXz3cZmwN73HR5CsI5+BEEMZ0aBDu/2zLCCgIzczVmLwa50vdYm
fQSfyO78K9eczObYIytPFct0wSSarRXUm2nFOgyO3X9KB/wiP+lMQc9GGsHpEW3q
sxVyF/b0O1EOrDY/HtS2QFItzpySDn0Wp5zg5I7H2BC6jwCPEPLeKCWgRlEEESDM
GKud7h55J4wvVQznBzh3NY4soYUiJEqva+W4YN6KaFMBzBUEDh/t/cPRV5SgdxBH
5EQyb3+z7N95c0Hgv6gEbEIOIhYDH1Jx+bwW+odMR9/L2+DfQskqd9Y8nBzhgJtN
nPwwVUfxssHa1IPelB93ptlJDzzysrOzhPI8Rno3/ewQTWEmB8E/kV9gzPGfT+CE
uxN1diyz9GK3eQQZ42+XyoH35REOWwqHPnk9+PoWIkcZtyrNOcdLdqXOF5kTyD5k
qqYgW+hwQpuOOTJVSV6SpX8wy/2c0DWpLk09aotNklJ4JlnsgsWkr2yxWI+Em7G5
95CZRHU2BzikShIZzc6g28VrS580gWj3JKeJqnsJWaQF3/77JMpCBvojEV49kX+v
pijmAH1/W6NP86sKbh6XHfnnSaCRs8pcPWIBXwzpZYt2qTrentGjcFJG5nAuFcx5
sbZqJcnPa6c98B7BFlGAJrYzJkHGNjUWZAy8gSB5h8QvcyJ2VxpvmjtUz8+m2iM3
DWeIoKIC514GszZ2QAiNQgSYx8nPo8nG2LnqiylAAB9OH/FS0AkpMQmU4ErM//kK
/xPJ3LCeq4uLEXszVdjHfzURp/wcGNG1T6n1gZWSnR5dMMyYB9R+vArNc40OuycL
xmA1HpilLzwmyP8nbe3dFGg3Xn8GdT2U/zMWql8FxJTZA/+6PyrmLVN+n4RJL6YX
Du1JMoj6O4RGnqdo8XZPyeQwyFbWogFjNKIW3QLgiYZt/EPgAgsoBiwqQUeAQdNu
PTReqL74AgIPooRl8aEumEg9SKDeyPVtmaF9dn76nnUz/qKmywSIbmZNIyQmcZ14
7lhNPLUjSGQI7toKz1LA/kQL172c2xv7CFbdElDEgZsa/mAfG5Mpgg7a99K2vr3/
B5Y/ixgECAU7YLKkf/f05BPO+L/QOQ7A85owynOEwSPBMC2UVxLEOO9YAFqQJvF5
tJnnYsQVoQTTvWHT3Ygm14W6TTEf2oUsolRVfzu2PA4SlstzqRhUn8PsCEyy83i8
GFyAvSN/4KvkHqgAv2APL8PqrWEOIhMvMA6VHJ5/LEye2nEcI/J3DAPMfDYq4UNP
HuN7W70UILIBV2qe2Cg61iY1QKWf8Dc9+A1JnAxIl8jUUE6EfifRgSPqThdEbaF9
aBbIoZI67kS1lIcY354oHS6rEJRcROoRJU4jr/gUcI3WGsZ6+cQnNQsrGbvHUuuW
I1Mkjr5S57xXwyaiyLCyVb5Er1xqIvPb+EXjFnquiHQbO4ANGMlRkbHUnTWjFPzf
NUESqBIILqdhus+tbE2xA9FFH8y8vjcqDN7sTF8mhmgi4eONoncUJAlOefIIszRu
gAUqwm9sd70IKW5dUSWomyRV11z9FCJvXt4a0wBSaRWu8fbMeVAGGSrUkL1GxTof
cj5lZeKxuRrszCWF3zM8pNtRXmuaCwbeo2rzuafXarGidFNLGgjwpBs8Zzzmc7VO
xpWrUHQr3TqfuNio4xdlLBO9QdmTXS+tczGRd+ZEcuwuBrZy8LS5A+m4Osix7F0p
VcBW0sDsRSbioQNXiCiexuXHNuT2B6eaHLm3NOHfD2cnizPTXT2C3qMMJTuVsBc+
xLy2X1vZcm1piwuff7jyya5lA8hQsXuu74Ioa9V8qeMW4Hy0woh6BRl8ILZ0+RRg
ou1Y8+NXFfb9AfyPXd5oErETbXVquJdXMm/iIDt53lWj51mBdyjWxn68sKKlhy7l
K1RQ1Z18t4IhPrCvszMUVlght6N5mpRd1MiBgkV7a9ln2WzySPudg8Po882r/dH/
/PJwjveQMF8xmDF3r2uIYf+wo+JQ/ls/VQfWXJlCYMBrkzVx6QzMKSKYClGhA48E
22cF0GHrOnMl8BmQSGe1pLt8fAUkSe5Pz9Kr9GBtkA7dW1wfKdADbmP0/mBED2lR
Lx8LGCtGuelrVXjhbJVVNergtK2g1AaEgyI1sqDzXmGR14UXVstCqGVw5Te0loAd
SubVSg4vikUo/fhdS8kde1Tfj48X1Z0vtxf8Spf3FoTBGty6350Nwc+nFNF+a5UB
VrMgq+RnYZRCjhpRQqwoLe7m5qlmzMtGImdkIQvQrebcr6jdx/0N6g+FKRbLp9D3
I/RrvVGQFSbe3ALA4i/AeYtZFsgOf6zNLja1qcstsicatPHPbVfeyYqsHASL581K
UsJvwhlq2RDaQSFU1r60OcEfN/wmjDKlegtNdtwfVpIsuUAnK436a76I6S1Xl7Af
nmskgX8lSAHsoHdm58a2JNeMLOwXTjgY8x9unvjLzExtpTmYBTZc/6tFcEcIiQrC
yJie3mkFMGJnAvLKfpF7ZfDgNFQoqECqfyXtIozhV0Xxw3jMN8W9FKrvEqTc0cFl
RoVRlxkaiuD7Ckcn4idvMv4aiV6ptrp6KTHCpuAV1zmljd4pMGFkhaOloimXiFlD
wsOIGAV1PgPFmvdZlJhqUYJFuUEJoj0EvYRm7l1TSUnQvLvQFdVNvmYjfsRG3utv
+laf921gCS5mLHS4O4dXcQU8u3yB7Dj/nDgpFJoS58xMRwCAAoFh+vRJS9b6dzZL
ByV1btMOGs84JaePZkHagG90gsxhnoP+1wIx1GdJp71hkpWmUB24S+5D5tHqP6yG
evz8RBsLUO9rOOEiCWmL/q1Bj2uVAQ87GyHidQksAzqpxEmQDjBYUxJZDRZnPspX
ZDZgVxecWiLahnpqo4CBZdi1n9qjjeXPueGJs9nLQHcwZBDNz20178gbvie7TKpk
HSJdTui3oEAstl8OsP7EYU3UHNSXB2J4v3d7DCFSL4b4b7K9AvOPInokMjUK4KOJ
cwKwh/RyALAzN94MsckctYpmzNyzEWS1Rkdg0P2rqsFT2tZEWexxNpZqVo+LVunU
O9jnLLS7aBS26/ZpFLn7c1ibsyM3lBXy0blQuKu6FN2sf61qWRLXT2WI5ZQpfl1g
z3fgZKbQV3VE8NJpj4cunfasKMy9NmIa4DAPsTB/Kx8wtdeap4jjmafmok4mfHB+
w2KNceZOB2IW59InZWPJDlnzvoiqU4atiGaF5gOeYDgb8VlNz8++kQWAn1vMYV/D
gw/g9XZs+dfOzGa4ie1oqNNxQy3BZzFNpNqVCUbLUXfny5NlJ9GTgg3x2LHNVVv7
BlAG64vIlekAxmCOro4Y9rAlUXEmM0gh3b9kop+kPV+9Q33WrCaGZed9LM4FWbAa
6a1UTNZl+T/mn7dF7GoEtqEH7sCnBYQ7CCD+05Y7tBGBuK7Cq0Z8afvod4Pnirlj
1/OrWFrwo3LhoYM/2pJOuZb29j3r0iQA0rJSLfNiEbKrDDXfj72fWqRyJc2vmDKM
shE6H/BqDq2I/TGIJ/47wy5dFRnXhQyqwAmXJGd8ryNuCWFS/s0NLXPEyjhlb8i1
Urd++zKRGF3LX8nOmBuX1Ld3fPPoQah184BVk5CHE9lIMIeS44D8bgGsu/MOKfaT
9pGFJSbY+/bsuRgDATIDC0dMLprOF0g4v2sNefCMPVxrbbEn907cZC7L4mGdky66
6sI4v0zAJKZp3y9JZswM3QBpKND3NjmlycxccvS7K84tot266TJHQE67W3oiByRZ
uSe7XXTzG4OiYX6fztUHV9k/w3oZU0/80BG/2akUJk7u0BXxqsS5DioXdeva2A1Q
xEcd1yJ5MW+YeoW7ewhumIdEFXbOTqipYHY7P60uiXQsQTyrdXg/IHAR1zZU2ozF
BUNcl5UFxwCNPEcH3Rs6aYIR8zL+gn7bqhupvO/b62jnaQbGiEFdgmrzxJQWFa29
uvjNeMgzJMcPkNnJfEWEMQXXSTv7eKh7wfX/6EeKv/8kZ6eiF403xHFNSRN9fien
KnW6eZl0eG7nBIpA9G1BMpw8fWSShIt1cWtr63qKOgNBIRoqILeUyvOotUGARAfx
H1MhLuNXXiT+kIUwfjVCBWAmfiq9wIGa854sNbtxeWLpMHFOPEbetNaKmpPtngKH
k5GLjyjCbLEmrAGrO42rGkziYVgK+wsxMVmnUpY4HoRU7LVKHwRWtRcAjfFMcUQq
64F2R/1/glshBouRCmU+DEOuTLWPNlrhZhpXwLlIoQFki9/L9GLuLLnWXQ/aWdUy
O4kVuEjykLjRCizvU5r3SqzEAkpam9pzI8gzDfNBErQyDVqs7i33mPKv1Xb8BOGu
MDRNDl6NBlktPhTDn4D1+w7fTyDT7yipuj+m7KJUq0ZrEeGtFucS398nqhOtTTHL
HMZ4RqBHCaFROTh1p0OFeAqYxztDbNQqVq6QZpXYdVBxzrRjqXeo4H9MVac3fISv
69WyDPgqpN7aKn9R57JY40J72gQAU2FoWRqszYqSw11ww8diMsc/GDvB/Nj7Lb+e
hJ+n43ge8+EW1JsfFsl7QTzqIy/bVcuP41VQk+RjtMjDdm4u3Sk7EXT+l1WDepbX
oRDCsgHcoGI/BWPyoqca/etGOc7/zchfBDxiC32jQMc7vVVglRJpmKVvSvA2MZTG
Qyv0o5oBdthCRJB5IX5ZzGmhUvJ/0Nlqp/GSYyy3UX3qhmsGLHcw8vJROdSYxW/J
Q7tuilw/bhEM79J2OnohWvyE7nGuLma+HM22j3kLsqavTiPPQV6DTCIayUre/acv
qSVwBSwjSm0ZL4cDbT1yrL9yA7f1ZH3SI7/DHPWuisccOhp1gMUkavN9dYmGbcHx
mVXMGAeORU/c7lF0OyWL74pFGVC7adAHa2hoZrYMkOnDIYKz6pB6eNWDL5gSpa3/
rQnh4ieqsjTzWi6WABlfpSKwytH2yqojMzTvbhR3t41DucGJssF37ybeJ5mzURcS
U+3RTpGAVoiSoNtQ6q4FdFzyMUUM5Ez77wEp1iq27vVEkBKkaazH1xx7V81Fd/zg
7RRUAg+y1j22yIceYU1Z2MvQm1v4vU+6NFBPqM//7cVVEhsCw6jDMs17FltxXpNe
G6G36c3B6QOxsqJqlNz8OkJ8erB2rTLtPVaLzW2ayul1todG30OmGOqw93vX3P4O
7iQMb7HWDA3Vb6K5x5dYzyMmuGunU3yma1O/jhwmsWstf7IBFI9BTihBd0Ro1pc5
JXzgp5AuvrfD12biyZR9c2qYiT4S2QpTWJC5QXCuI35u8KPHByUKw6Rnt8HPzfE8
9pEMfzTu08Barr6rL6J1eJFCH8u8EJ4ZEWqUXLjtnUdKCwTkNDOTljvFoyAMhlKi
UUmtwkQPv2l9vZEQZaCe76Rh1xpuCbE+TTz5NTjbz4SBPxdYFdXmp/tm/vULIhuo
7ydLof5Z5DpdmG6gYUt8nLzVfoRvMO7x6hLUMooq0st4h7gJNoCRVkZZy5iLkDru
iNuTgxPQnQFFfVambINMoSLFbEKS6zD5nPqFrL+DlU8IJtuEhfWuB7nQfZcLqLvq
IWYPRY7gWB5XmxvUCyP79Nd7bLeHxBQMY2/vlQRzTB3XGAIK0cCS/S/RWBpPKYxY
f46a1YLYY7G31JzpcBcEQnkbsa3tbNkVuPrbAR1ZsI6EAQjUsM91yWafZRLdX2BX
5mPg2ARNUtw01JlQWy5QBvFcA/fTKNkTo8XsdM58q0E/sGD4I02HV0/HTopBd9i4
wpYTZoGvRsZtX2YPBXIoGMhpXyziR7Nem3F3U7xHMJHdpkJvXQb5b+NziHR3Er8v
Cwu527GUnoLzjwKNlOuKywi9uxmMh+QSqS4xgvOlegx/2v7Zn/daz4XR6997km9E
h9Er9T9iyO/2eyk4zsA+78b7UvPxlD3e3geqzb4D0kwuylT8fVWud075NfhAqar/
0neOPxx2yaj2POP0YklQ6Jnh1hPh6Z5KhJNQmajShpfLm6MVOiQlw+7j9jIbtPuE
7EuA4JsMxuHZfekoHQ4jBqBkZ2kmHk6hGB2m/rYqQlJnwrmPVg9i1zc97e+EBTgP
prqRJzWU6GrcX9Kuj/iiQ/Yl0oh4u161H65WEaDyakiMXw2OMgPBrbxvwGuEMJnl
2ITIWSVY83cYH9L79Kgbna1WbUTveH+6yVKk+lbbHN0qa5T5Jpa9BqVFYupSTbDH
hRv1YLHii/wAIRjo7rPkVU/5nLSYoWncxvQ1WOOLVS9FrnajhR/WnrcBmIabGdCY
xFZ87Ymzr8ydCTNJaBBAd0fN4I4vfZxFj0nfyK+Q1vz24i7mR5UbNEqrDESgKOdP
7Z73gbdZ1WsBUsxzH/ymd1OgYefz+RiWpSCEccWyHickgNoHpP87BI2Ly7FTZ6Oh
PTQ+cZAbnpE4f4p5OYuyuLxaoGGamgWSaNfa3mW09mRSuS98+y3Su4XWMm6qXWaE
rNBS0ppsxL+JqGhi5rHRcY2dE3Pe1vDnk/oc7bM7Yqm3rOM1Bo84RlOuTHf8WwiN
Shdd34vw3h6B0fslupKTPGe1S5GOZ4xNUwN7C5xO3gyA5BzXnu9R/JzUP4WKSG0J
0+HV+M/NCTgXB0QHtjC8/cUJpGhmdi3nFbl05WvlA/34URvyv/jyyV+d5JpiGW3J
X2TJrnKSuk8NhvWuPKQbdk435+pSvwDnheFLUWRYS7o+78OVyShlINg0DoMsHOJP
rZb/+isOsOyq6WAZPEg1Es+SF84kMeWEHQhtdV+MiQwEiiu2XfEdXoFCtskS9YET
mfHkwWErV2MwTjOTK8jJMUe1XU/HTbXYZ/8yYh0t3F0zyEGUnGjPdeWg3msFf8rP
+N199t40JNc7YvrfSvlEEFB7RnFWPNI+CzXmnIimy7R9gQQElPFs95AqDN8jejAx
wUPT9WTyOuOmAfkG1rKrs9Ob0AcXH3P3Oe+t88XGWL+EbXzURaBHLVOnqEUeMZiZ
8Aj9fIrnp1DGCbF+/DQ5YnNYAgMr6t/lScG1q43WBLgMFt6wMPHnv78W0tbEhs+4
qhmaaaULRU6NKAjpdn6Joj1aXUrhMIBwRh86mcackGQoqscamWCumQ0RdRkty8pL
nmhaBm+sclQSc1MLfrlmMYUKuvi8wEBN0Ky65zVdL7weAhWwUO1I9nIiZFyS0Kt/
tzIxxf8gKp/juhdOrm25Zf7FnEQ6bY4+vVg1V7pVu1zlv7tN6XbXO7HgObvdwlpf
f0udoWYgbXZdt9XRxlnI+sBTTO25cXsMj9fAUO3PErhnXsRWJ1t3KVObH6xm3RA8
7TtDy+pUmuripq4HWoIgUj3o7BLnI8pV7WTu31MwMnr1dNk4SKgB5oroSbAMhMKL
oMOTMcEEnqHd9P/fQbqpBN+JSpD9xVRRlwqRg1yzchsgVUDawFJYdR/TRu4DRpru
uk8q0KdB8MQdp0lecQsyHAEja+wK7Vvcl75EiGsDOPFEfsD5oaZJAbxfcnx0S0Zf
i58N6EKVlCaMHkDZTaDLt1MuaUCAB5OVRM6FDAMVDr/GcPJoXh/JTdEz8BeP0xBy
/NXRH6UGnccCUgQgzWjkAka5DtmK5VFcfj48QOWNBiEwhiJPZ4woz3/dCbtku2Rw
rlygAwuVjDNY7NErM1nZ8MMu6yilauDjG0+U1B2c8/O9zZ2ReT8UZHb2Ci3UqjEm
eUXgM94HwQQe+HFvj2FiOtIhqYq0xR/vbk++5cndnxSfHwN6sjKxvMlBg4ADPKS5
UAT79J8Ux/S1CB6EKnOyTM8pZDXBJJ4iqiK/bKxGs17vH9fpMyc+5ZlBwWYbBcCM
TxLRqD5HEuh3eiKZ7VzHxl0mJuPNeZ+GgUrBw+w0cKGIJ1qY+xA236fYpYkE/sMD
qNuDmkdK8lAuG8ZMJU/+7+wG29bhU09MXrltgtgqtHuiXhU2pqf+5iQgI8xd+lQq
yxWyFm4U1C/mpYItDFN4NndIgN3ihBVn9/jSdKaUsqloCMJVtZWb1gkIrO3Ehhqv
BMnNgLNePzWarWfeP4BF2gy1yRWyIEtPnZfEMym5tVYliE6Av567lujunDIrtxZp
Q4my9kI7onxZ8WGBLQJPhOYoCbjYhb61CtGFu1HlyEZkly+n5YcZPZYGZWmTBk4j
udLs9/wnEMUnAOxf+aED7QQP/gqFHKC3QS7wkBtARE50Nhyd70hIjq0ZjF1OuEoo
fZkRObZtHiQ9bNB5D9cRmlNJ+NGG045Hkpct2E5ueEuL+X0MZAPvsF4ccYL0DhGj
2GUlSAQ90vbHBTIl2BUn3yrymJlcVvTQrs9cGThxO5cRKE7hpKWBQ1OlzjDun9VI
MN4+2cWgsCdk4GPRl0haffEuP6Gg5bJExKNXCgeAd+4i+g0rhOI91XTjFvoEIVgA
Y6khavlqNnqWvwTQKR11qFTrplbfc5+yL7JtJBpxxrAeDtle59Q/l39BOUtoBzje
MYsp0BG0Tgo0YnFfpWqnNIjt2qpLka3IxFON/GMriJ+A6Scj51R1XywIK6DHf0bo
IK0vULUdnBU+ROHnR3v78olLDp5uw9+pwZNyqqrVTJKJt6hr4GqWL4LGcYmA0DOQ
qRl4URPraIkqQPQt2zW+KvIpTww3aV6wQThX2FiEL+Pztot0V5VH9ZTOgqN/nb7D
i+1OCqYiXSVqtGCwR4HMgGelEYS52t2odo1QDPvAVIYpcpEPgecyJ+a4GqKiTksY
TCfNV5mgyy+0jtFPAle3PiNsaAl/nX2dV/5U03OujyZacQ1T2YWUTrvRZuE0YJL/
BNMsfRwk08V+AbfG9edNbyQOq0qrDJtO3lfungrdJ72fxgzDM2ajxdZT1BzhPzAh
jqqdYg57lVM44vXOP38cAZU5fSbYqZI6RPjg7TmPaXJrMAlDXXtmX7qGaQDp2V5C
dyCXokTvl7LiyfxQoyWg7VhOOmZ2FRDBh7X/qASzfJ1flEaZ6ZbqMbwbp0sNTfTL
G1jhmUesmvneWk519GmXtTxbmr36QLyPJMFmXpI7JGOJQpMZQIUYHOWH2RRc1pSz
bf0nT+dGJYOVmubV1TH5p/d5r2NYGu+CU7fEt6JcqNWxglZVbYys39A/SvTieYdF
fUPqoXvm7WXu6EzHj9jgWKPzaFotOsgLcSpOYqXVuswc7dU/3BPvwC6+QSVWnDDO
WpjgZSYgyfslU5nCjhUwl+m0pW9UCO5X/dc7wd8zjyenxkFusiQE8le0R2g9JMgf
UjLbKHWpSG6w6a9ZjIE9wViFdNa8sVrj0ETJsYOOcsyYMCfs1aHdB8lFe5q84jp/
BcWEmEYDPoa3rbLJ5fBdgBfA98sdEHG7rdoJD/YnmL/zGI0bnuW7X9j5GHpYi95y
jYhf2+dCFFm1CWxxfXRhQ0+kcP3k8Eb9Y95Hz1oK2nNPSGIa+EE8fsJY7ubv+eLW
we2O1zU1jeFxDyxZp5uh6xDx6xow+8PpmYKaYi6zQbO9h7/17m94nHy3g9hRbsc5
eH+Dog7395FNamnzg/WhFWcg6V3W0X8O7mX0iDc8gGarGOm2/CbS+NUECBJdDvWT
Z2dv1woyeP0ETeqg0OkRKMIT45eFkBv9GODHLLKi/Z+/0RfZiavm8cY8c3x3M7cv
3ayEPJRMwLHI6Iyagw61SMuRC4Vdta1H4zweQ8s/CJa5xsTp0MVmqQD9OjPCgz/9
5g+zCiZDwwTB+WWXFW5Ff8Z8rEubCV8+QXzEjmN+zQnY0bdamDWU1V3Yfn01ZRMT
JA0pARS9fyWIZCSHZvvVxE8CcxdVvSM2efymkQDSgdJUVY/E2jUkWbkY40KWFjZn
JcSPa2q7XZVCAFTe9ZjlfJHBN5HBaSNWiukMyh+22bkQ7g3dna3YRmq+Z6V22iw2
rQF2lqXvstTsyp/HxIr6JPZ6VTxmUm9oR8TEinsMqaBiTpi+ssPfTB9W9+rdVHY/
dJEv+Vjiy+rqMXgIJmfkPuCb6AuIuVwWA2Ii2HIr9IlRdJue4urjoxERBKr94ImP
jgI1oDEVhQUZPWjF8EU821dh6jM7i6ZRSVFFm4jrh9ODhpeRB8utRxGdw43ZbAVQ
7c1d9ap8lN8eMUJMfJcpmb00gLTQjvr8gPw0R34k2580vNTZIjWsfIGa+/vAmWyM
A+RchtvJnqVsQjDTTLRd7Rn0VfTjdEApU2SHudybYDKVD1P1GZ5uar8Hk+/sdX3v
Qng7BM+/1qeRNajyy9H9a26tXiTBVN67oPtFtHzCizGeZST9I2IhXiCPg7dxF5b9
orXEIDEu8DkicWwULYCZloI4Vp4WQsZxhkiSpZbsrt82kFnQSU7dbsUIz9KhONM9
MgcgrVsa80kvH6BnIp7+8kTa+eNvH1BibFkRbRIdUurADaY4KzXwbl9WJVKIzly8
y8llJM+g4bI/w7oYpy6sWcIiOAFCJTmG4d2UTiAepgQjjcdeQ4quLUEBD+BB9pca
OGmp02YXSBYt7glr/3B8d6DEnkudil3gEk9xgd/N6BnCYp2lViHbQvplVzG1zDMo
coAdZGyoNZsUG4Jyo3jQ6zoRpGBDn7AeGLLWT2g/9JlWXOobVpJvpQB1ApcMRIKd
cG7qz72A5Vycqg8HKaVufrEsGBa2WEFibs7qiI9lXANuxL1ZRV/F/huDmqjZ0RkR
B41j0oyZ+lu3unNiuuG1uBPRRPl6vZtwwuwOAJOUUekhKfJTVsMUUrEC3YOD0Zr6
jAX3H3Y+QL3gw7NjXpmNFpbWZ368IGNIyMYbRRy1imfFTN11HnOItQ0mavkYRbIA
4M1/52o046dQsAl3o+Ng4XkkC9YW0k88iRZ3eXdYI3rQkRVKycRDDIn1ajbsns+6
Lgu4e0Kc9eWI4jmYF91Mvrc+d61UNRWRhAwoL6uo0e6HVlm7XHL25Bsd45HGVZQd
3pFAuA1iL1vTZDdNYAfe3nh0678QV1p8/E7tnbRgFrFUFLD91D+TYLrjwtXrB2BL
ml4X6MyDTI6Ul+jLz7LVudVYKqMmgfgQOpb9LI9K0pvk423WzNaiCWvY6j5tleB3
dAHpgXwIU5vd95wBcBKr/KYTiBA4CqJ2B4Fa5lWlr703OaFPjKT/FGemgPu6pONl
E8AZ1c9xNkYelJSS75PWiIQe9aBXIyIwnOp21HSo1YY8omTLFmBspLFeCaw0bhqA
RJoN1NV/cG74ZprbgtUV8QkBCuyv5JV8K9SyBQoVZBCwvAimxDStdWN93YorJNPj
wjkL3dYH/RAxyKbZLZ2stqD6UV0gbkZh6U1OJVnHmjmA5UwbnhMAeC2M5ARCvFTR
whnqgvurncxUy39WsQCdeAmU9sHYBlHUsf5kJD+InqXA0Me5MiWtHfk4cmksz1lg
GZ/IPr1Y7FPuAdctzVxFpmlVYVPu6oXEwIbvb/eSjdasZFJvV68TZiLoDf4jAACp
eLQTNb1oysvUKpOj9eptdNh4lMw3atNC7lbkBAQS11YUblPIncLmXL+ls7RNytOw
owP6jVUNHcEaf818D6pfazsmb3czPhFwleegFbQOVI+Z7+Ji7S7zIvhu31u6wbT0
CsW1mW6UG7A/QKcICU4eDlHWjjl+m1LHiGruQL/HF4VbZnkebRC6JMNFCQhLJAn5
9Mn3hIZMP+2x66iyjmGaGUAPHLRwxbdXtDGxAd1IfVU+Pnwd1IzhAK/MsoWw99e2
xTSWuADhxSx/q9+AXEbFWwbYCJOUaaoDx/d84e4CoU3w23/zgnqVpLT+PbzfQVqw
o5KI1HOq79GJG5cyRJrLCV5i+tnLFOinl6MiQqUFkYeIxal+27yK8GU8lNGN+u20
v8n2fHkiJLPG5Ir25DxrPoxfYCWqrxd/wy+UDPFL+YdSx+cBW7MwIYMDiD6QLI15
5dSCQKjKkUc986h88jqsMhJFpsplLjGcB0AtPmNW650UJfFRXPEO5osNBH11zgpw
ogOqx0Ey4Et6xUUmbRcghSnB9xlDwv85e6BxJ8ZHI/iEtmFvyeVzPGabnOW7ioop
4n+tQagTmbbQi5MaQj/trcSwuY6ZvaCgHBWzurBe6jFNmrKwqlis9q/8J1P02t46
p8gZNhxfJ/sTZwl8wRu6B6YtWPDOjusuBZsN+6Zf67F993gbfgudO5JIuRfDZufW
YW09ZN8OpBv7xpH5jEf642hPSUD3DjYE6xJcKIcOakxfOanEjzIsRwht86hTP6mh
AwHevlxScufDRKwVv0VeFgmcxffbGoR6TYtWPYvO25rrCe89OKCQch3abZTuWay/
ONRhJVcyb9NENK5GC5/dDN/uEbrY4EwrH6J3sMXk0ikUvcFcpYy8+6dPBJOpGdI/
shtFEM4vWvo8KAQA0mkc5AnlnrxdH/tC5bkj+9Q/vHAL3W/6P/eayBIZPVQBFRU0
5U0W51ZB9Cnrb4J8u02bpJX8s8ScVBuOPuBXuX99g2wQZPWM0EbhlgAtv8s7xAP8
oFRuNxepdRinal7zBxqjssTatEfCKG++TRin8bsFMC2JScA0Mgx92GXEapKS9g4J
fg0YEzImdH1GTOnapoVtN7LUFcTgcy8HWtHmsSer5lPScJzjbg2WLqnZ89Iv/QnV
htpJxWco5NYiq41AGFwlwqg4nJikpux0uaDjT6sU2morCk89RnExqY4zUylgG8cu
qX3gNGaqKqxYEiqwReg3AKhiOs2d5udp3MTRgvWtwV//HNEi1UWUUMYDEreH8e/N
Hg1Q2JveKFMJykp23dYOmV96yZ50S22NIKjmXTzcREtrYX4l1r0LwUU+tYkSFmTI
5+aKhmNA9ui0pDxLvV6OOk2cDoLXZdbCo8lIIhj7BApVUOrbtfz79+Ct1UCvPHDy
WleMeZu3FI0De1uiwzfAU/QDefTcpLLkfauCKaUP3iEHrqsuRPQmfd/MEvEnCP1s
sVpdFPdkLGF3AQsGDzwfbcc2wFTQPF6tD34Cb0Gp1wcgoZC5hwYUMgdO04Qt2Im9
nHHfCma57gJ2En4BCVSusz0sKs83A+NifGX2ljrkoB6j7Su9ocRuoLUMoi7WWb8Q
LRXPSBuBfcPQs3k4CCsYheVr88rXkYiWvtXZ5LGfX9FF4sOW56uRw5XKHV7g6/Eg
gb+VTRst/M7s3Vy4rCjRP90aYeyWwlrkh84rid1/hfYdG84VfumBGl+bXfXOtb8s
B0+9WOIgXbe0E/vlWxWYCSNen89BnjVDoY16n+IUmk3wZ1RMb8tWKQBxUm36qqre
/P2da/d5dDFMeEdfKpKE9Axe3KJ4FkEyLezGv33wOFQP4SuTvM9JpaHqqfzg7v69
oeRKEPmnehCObln61t3lgzNM66oxvqTXCIO0gYXSa4mYcbXD1xQ4tCqOaUoMIkY8
eWccKp6NvzERe8BuQrOS8HZTbgg9R791DBwZoacgFG00ybgin4vu8Q+iBrRRiqp8
8D6fMa4thOffuj0pbiy4fYEDTfB59KAycKM6qSLlNrP6uoITclSYs6OuPETHPPb/
aoZHVCIsbYVWuT2gWmLzNqHyX/Uc+UtvOFovnuOx7bPkoKKxWdd5k/PqT0ymd7k8
xk/Y1Df7Iz8NUiJk4wPNgX4npJBiNiAUg+iHy36PDSITm0d0bQGPKvAyFdcNGX/Q
06lu6ExypKyGJAd6HghK/kBteNzAZsKL8ruyGhfXmvPQ0BcaAfa1soze4qpa5HmH
mUTOeucmgatsyKPSEt08pHZh8RmREUQgqksZin4JPEKA22NtjOgnyhGmDYtBFEB/
qnOV7cbkjXZeI41+N7Hb6seWyildKqzszHy630xgmwV0w/aOB8W7lUyui5xhV4KO
9PCTBsWK9eWs+5R3nbq7Y9Sd4MjmxZPck3rra0TWncBxUzL8sG+mt9EViqwgJDsW
XYL7XlR0FIC2nfsNCC9XPWGJ1Iqe4wchj8jhDFIo7WwhEEBAWYU0HdnnaNuRIasB
01FpYYvotM3G0/bH8E0lr1Q49AYwhRq9nw4HbppahmOm/DYVnVjvy7Kq44mOTDiD
klnT8xGTW4vZnFjUXgm60snybMmjsNWHgnuqQ/OEDAluMy2ZNnBt4GQvDsqTBT7a
lqq8FlMbpJb299tuC6Cj/vo5Jh14m2fkriRK4bsPGW0UONit6o086r4GT9Ej6UBi
hjn9U2mNZtiardY1WUoNmrU8698AzonytsGIHYAbcpdif7MhAeOYVF5K52YyqjbW
P8tDNDdj/o9+wBpfyMGBnkl9OoXrTkPxBYGzLMuid92ZM4oq6sbi0Ns316Jtvi1/
DSN7RpbRxaDKMEmGiNp9AfDVsLT0MoPR5uNg4gFKxgjAikSfS9Gq+pPTmZDIapO5
N+NU5Sanaowe/H/Nq2fWW9V9AcwoBAf+PRdp160W4R49x/yvqOeP7w3t8SH7Bwqh
cZ30KoEuAUpw2NibH9IXLJgsLY3V3fP7cSBhnxc45yqrXRbm2rXWVov++LeVOhT9
s41kw1jlRIxJw+K+/QCZ8EN4VDSGdAV4rxGHcrfg30OC9co2DQ5+ir3fLuV4iT6R
WU9IvzSxlP0XwIBhN0jonDa9c1cQZ/h/YPZcVIQK9mw5f6cmgk6nOuYQ86SHMGo4
MqXYGe7A3mmT6wJV2XoSbOKJlR3ZKspFz+Wr6l/km+URgMEjsuoX+mMI4JbQLnQ2
2NyVVpgQb11as/pbShPqo1xbiNHjpEdFiFb23VevdpbdFFTZ4Qh0wLMO0Emq7Ont
mpdOG9ZhYt33eg9T3FR5kAMO325RBkfSh1OQCPGjEKaAUmbJTZxnvrhay0im7t+e
6k1jqTAk1/t33mHvHtYJ19FV5aJyYnCdUq5j6h+5xoz5VUB3oOfBWQ7fwZg5EBJT
N8UYJR1Oq86GtFLPm/G8QEIx5dyAjK20fpY50NnhStWZuJ74piBLYVx7VQOfXkhp
7vRNSxu5J5DBH/iRD9P4sCWNc75Hh5tIVRCu8XGl5Kj6PB6Pgr1PBLkP6w6UBO91
sh+h6S5WnydU2N/XzpZa3cm+5eDe28KB1Zsc+d1LxJeJ8PlWpPMa34GA4XvFTjni
5x96e0Az+2keCn9rYGg6WVGRt+4EBb8iLT0Wr+1qnfsVZ3rvc1v5QcLQzz5vhzZ/
UWJin605py8xTyclMPJcLr2I1rul5Sbiwq6lFS7gEUoHysDppx8DuqI9JvLsvKf3
yMRnbi0yMutCVeNvogJaTMK/Hs/FWebhMk2bwM29epB9RlUGfKqz7hCbpSi6NcX0
Q3whigRxsguHsnLRtmXG18Jw8AyArvqvDCCkjlkwuJl5pq9shGg8Cuxsfz1fsSbe
2jJp0gyqofmpWNWtnQsW4/1GsNsXpRN96PnTrQLiV1Tj5lG7DgSPf4LcfXsxmAlF
cWPmP3LjFKQXPqXVxe733KILR6nlT/3tSBrC3a4Z2i+QGoOoqeScfBrOeynGrCpg
Y54Uiv+FVNNSWY0KoXOsP+XKmoGKrHZzQa7cDj/Mlezm9mGOuHIPdRG7RV6KKJmz
W5SsUkVCzQpen58UbMnVpn6mMrSXJVM5ORWem8Ldww66d8WzzkQ4shsRJ5Kk6T1w
rbLgCNOWhQeHjBxSGe9RmMRw+0/IFIa4q9MmrQ4lgne4dE4H2KOsc764tRVCs3eb
s2H3YfCYU10wWMT/i5zkojte9dtfckvCw08Bq8aBw6QxgzlyuwxnlbxqoMx0byNc
snsHtdBDHdg84O0rx667jr6ylZETyyXhN2tZnreXOdvej0qSTdpKG7LbidbnYdZ0
SqvFepIq/wllpu5r7sR6pvrZuL3zPzmPBnhYYon8j2WqXCevSEwEwBDrlbTdyPwz
Qnggmwdzip2r9xVzmTDYQVNLIMTvajiXrHUo+elWiP3WUjCLwG5AajoLjSgIGMiu
Gd5FmsVF3b6+m9OdsfxfUuGhfzmBx2WpAZrxI8kxfk0w2UM+iYsGQPVgwedTHyi4
mSddpQ8QsJo/YLD0NRKpUXlafiX651clbeoWPlCoA4d8e6QMpljkytFBidjlsTOu
TEj8KhiVc/n8BC6SRK3ag09mxDfH+oRNEPicWlmvYqNu2vCQu0Wu1uKqZ/tmug7d
ebCNgbde3246AxIWOly0vnZBKztCwRJCUeICGqAHZDpi5mEz3jfV09MJaJL1IeZG
ybuTOYAPNsPRcfYGBqOAFKWnVqNUBu5P3VnCv5xC67VKtg0jzBvAtX+akctvU1wL
Mtfe08fSxhwzXA9/nr6jH8HnTWo/1mfKIfILZSsbnJFERI44MUwBd3/9XI0eTCBf
IGPQ73XdBn3DHizkaN9KhY00pYRo9529nps93q0rNvulL1bXIAW/fcdNLRs3IiGE
7Y/YNEYh5KnFZnaOXBaoch7OZVBruEBGoOalJKpgPfGSq2bSAYRVVAh88ae2nz0O
Fgfz/X5ThslGj2N3L7N1NPGIGpALbeW71z4PADOeRgBXt5CkHCMnBFHYQonNVf8/
dZUH8rYxQHNC+lCjaHzsV6pKtGycdsbrzSyynpo7nZGE1fxrlz2XIE+RGiSjIJXz
eGKNEt3yR/5rsqd8UfUktteppIUpAqDCSyCoh0j6JfdphnBNNNIdH31EYRKCdGG7
x5DQ47ms3uRn+YUXIHZpotO/IDHA8cAxS5A9/5bLjcFLLhpa2yLW3AD8x9ZiSSmL
9B4iCmmREhAnfblot4jj9z2AFm706uAGCvc1qFeFsqYhArYiIHDYFKWeBeh/qvJD
+bIEa1iB0yA897EkrE+Hp2MmxzTczH4fB/663twefP+SuhHo3ycLEMtZHL+ZsGiR
fFbXPMKLKx58ifSFw2Tpg+kCs2mhUckl9BWsKkdWXbI1inBpuEkYJ1eocH6KrHHu
5CcnR63m//rZgv6teA2i43Eo6iTF0eSz0oEWfOjPUsf88XOO/z0aF1hOolRqkmFG
yBq5COJKUx/kxAhPEBDYKqpeHSkRLqtu2ZKd6W+bMl4Ou4vtFmvG6OPghFxwSYIe
yBFXaI+EYUpp2gi5ZCpEqwajqFwGZZmbtJp9vrSJ6tNIo1RuIaP0jR092HGLRYTl
YDDr7c26TjyOuI3PoXvNG44SL3GRfa59O7wDwMyK0CqVmsm3PISe4UbFB45gxPZI
4Piw4X0hgLFQSgKo2OYUmEkuBPHZJ2zlUveYfZHBdnVV9XeK2oIav7Nz911V2HJB
6KoSyOpcoI+7Cl9v+/YXY1VVCUjZIWADms/YsFgm+C3piLrf+3dA+TOzAaRWbBQi
BHktJc2+4GhZkptZ3NdMzd51BEtHhlQXIhF+95bW9CmRYEef86Z8ALk+r/MtgQcF
7+8GSH1EogLOomV6as/HLvOAzOTOAEQx9BQYbrQ/FeOIPtvoxN68qDaiD2upmiX3
6iimL6dlbNaGrPaRflnSMHT4HaC0VTz2xwfGLX5dLPxRyiseN+cZF1E9PXrDnXhb
t72GCjF/BkZ9waoIrYCkKbZ7GkBLzpoxmR6V4ftwKk+mFehlrmx2lxWFod5FWnBc
kQAx5JDnFsaJot2xT3AYs+KDgbs08Iont8M8SM2WYDsddjYpomHbFTUJdBRC1abf
ZNMU65chWEioQJqaLslcoZu77tlzD7IVhTPD0ioQOaCxqegaOUqgwSf1URFI052E
e3/Vh3Pusi5z5f5JTMGrFYSPxWdCKw0Rex/0FZrHXcW+6HSMlqX01YiwItscYUiO
kCv98QycOvWmuyhjJz/HqwafytX4MQVxzx24bttz8W+wqlCx1S07kDnUW/DopaTT
2kdB8Y/0G0xRtZG6lohrD4MpD00pYcgZ0RU9qNHFlWk7IYkBjvuRBMKSudikflx0
oE6LoXUaSrBeQlEKT+V0B/f1K9QQTbvsHrO+YyUSoNrZnS7fZv0MFEJLv+gYqJr1
aJB3Wrc9yraBSecVTuU0/ISQB0McG0kJ169AtX5pl+zEffhvXNkJxbJSRjU9oALn
/zdEQYmQyKdkEOYXTxMc5w2D4cgHTNLmE/YbHbMWPlQm/7MYHqnZpxGhQC+X4CLP
MFmgy0lzktNTNKYsJpR2ELcwsoCF82ntvjmHqIFC6ndQTFzX/bEY1n/Udc4MYpY5
YmhAdyzA4xlIDiAMNhXcj68l2V+eA75fENMWB2ed4idf/b0lPAFOYOf8Ph8RdmEH
gdm888edBFkW5qh/l5Tmn/hlNwibVja2YaxfDYPHKRJ8wNt3+V9CJRK1bDgkglwk
RFE/MokkL4msvYXBfy7yT1JP2dUzVkb7TfB+D7lJt4s7Osk+mG94IunFm1IMOdGn
QAmir6rcjh119S62cNmLYKJlx2NM3q01k3Moqz0vfDhMF9AdScftehyuReH7N8Bg
8bUwCz836aOUzwqWQue+P9a7GKfLEz5JEK5/GOFaEuTRNkmKiezKluXbbeHM5JxZ
+zz7Th0mMK2cMlk6veYPDI0bLFiqA9aTA2ewT0k0X6uUhnt1vx5UJ5o5nVV/2fc0
c+DP8KXo9fkDDiwewMLZQ6aheYfhNFa4XbOPes03Dv1fyHph6ypJCmKTGTreGSCE
nCUh2JRuUqxWKxYBY20da2zBEIKqtgMJ8BuMGukPj1zjkpUSZd1/a/tD00nvszSw
ji5qUlrFsq3XOyuZNppWWKHs89zV7aYJ5Ysgs3zVADzBNJRg2HUOFJIuoZ2ioc2d
fe+dN90Lb6PMCaMpujDpX+jB7sH9hwZtKEDngRvEouUStCk+Iz7B1FRN52zI+SlZ
xjVP93muvj1C65+pYqCAO2VRPqovLxrgZ97XKLTGqz6DpmhfzLeKq3oZ8Ja1/jOu
MGDWrERw+wvnEFS24CN6/mf0NIKyGyp1/2GqTBTcp0Gb4KqjjEMEQw3tQwI64UWQ
ICYwaK7esM9IOX4pQvedl5ATWpJGgSqbLHI2UioCXqZourDy6sOi3F0+f2wdiaHt
yJjJfTqvPK2kz7P3fqgw4BaH6LcMg+f/0KO4P6cD99xGE6Vng4vA/4nX7O6pv66S
1u2P9Q6dYqVFmVETpl0cudqDUcdE25RzKcmgDf9EuupkYwPMsi/rmWaGgIu305zu
zuDQ6/Un/nuu1bOSa5lbJiOVZ99A5g2Qu75RBelUCVXiimRurOcP+miUREGglezB
bzf6uZbiCUpHC0Nvrfxg/txwLuvumqn87wovVIG+IdBwCo0ainvNpGz8sKYzxpnl
cHjPfGOpL/TbkUbOF/VXQWWGR36OHc0cq71I4K7uYYHbDKZBzBtfErHUfdv8Fv5x
+0OyPlS0YUvDOeToImW/dEcPOEzHgbm7ZqiNeyUnctDfK/2FqQHcR8fLWNDZmtVC
0X8G8Lsl2t2I3/Zm4Gyou8CLjB9Bo584LUbHrcL+n5t61jhJ/UXNfsAfUYQPfdHR
CWcpcEmDC3Ne16f1S+QbZVY8kKvtw95IYesx4vH+bMNEXSENFxUeF9wCKN9L4Nuu
fVSktNMrfjcl7SRHkCtW40HKTalzhbh4XxUsNsABkwiWRgjCI80oepyWc1pz5381
S/FqSMe0eL1yh5dPU3vZNrjx0zD27LSYZB/Z5CUE+1kuSE2FQt8kxoEQwUU9bpxC
iHHiZGGuOnSf3BMTe/pW74/4WfdYRE9jMO/DcO2w+9Pw3jpPn3HHThVN96VPWwWx
BsniYmXNWdZJ4jkdykT4C4t3z50cobiw5e42qBUm6ikBLIhc/i3ZfGw7nqFdvBN0
N2T1/82wU4+ZNDQTIDridjUtsogZ11s2E1OMaSvhWvNRiOCFWdXEdNOT1tHpFvQ+
A91p0f/IHaYo3Q1y7AT73FRwsEw2HWkVXm/G8mSIMt/blZmbjfQ4BVBo1o+iC2Qd
7BlA7uWdlrhG6zb25NtysDxM2mazQtF2tDYq7Y7yugIIRERl7BQAQwPMUU7Rfl8Q
Tr5ki1sJkPabgHJ1RtBTC2H8gXflYWqF6Ww3O2NPLW3WD8VzF6h9QWZJraHYSQBi
FFyzfrNF5UJnRVXRpJ9Q/Xr3EtYLxU/fo5oCyjF7WZ6vDXD4iyNTHnJjTqee7uQI
uLFstYv/0iEdCG1v1zMbPkBNAwGsxVzjfFHjtocDGuW1qsnXAcvB1I8NoykX1aMq
7gWMeYnPuZyNdd86XPV452d9QC7XEp89YGtTErbEYh4I94lh/p8nqhj8E8mR6IqW
jS9Pe2K1405dEUKzxLqcVzQRIermuOHY4niNfiHvQMIrkkYwxk8zxYM2S1WbJyj5
YSu5o+cbeMActDboRfrkWy9MRueV9TbT8CaW1JkmqM5Cb37bEm810dr3pCfb7HtB
snVv1NrhIDO0dJDHDe3yxtJq4BkcPDE1LHuu/VsFFgWE0WrXBbxUnPypFZFt+gDv
9mDRzjrann/DN3FX34owbB55lfjHH55XiQuwRnuNvK+APgZzHcWYrTJcIXeaToFW
vyj5D0kT+z9rHQRMJU4xGwKA7tR//g6jPTEF5fGNRIMm1PmtvMzoVUApD/24sLzp
8jX3UvANJUaFyluvJRIPYtKj1ntmTP+x+oSZAXxxiyfdaOYJ3DmsFEfz8QE+n37R
nPsybEfKqOvo+JtoMXV8OJHNeDYX1lm4m3Pzk2UGrPjt+lm3Io68/dxN3BSPtuSL
18s9VDo6DeJRkdrd6p9tJg4IlUJ43tYKcNj0/sTdQL9rIBgha7ZIJ+LHuph9F77m
wfjwZ61wLkhxfSFzWjvFBPYjxc4JIMZfy+fqIz4GJYZkYVckR/ZPtpeOkHJoBa1H
2APuyauo9dUEayKpOamOsf+x49J4loUGpGUhYGjY47CK3n1wSm7FogIL1drCfvo7
vqKI9t/eGUwZqIKCoVVQ+dh9jMFBXi2zQFa80xiM0CJv3Tsp9uaU5GZmH3hIvbq5
Z7NRdhX9ywtt2HcglO/37gnim1fjSuwJ5NYu4PJTwWbA6peS9jrX5HIwf2lBMkcS
ykbDrgtHaC+sw4UVAPF6d3wIoHdfUf0DuKlNgAn8apXHHenql9STuPk+nvLQJioh
FIsq4gLAiZCLCZU3VPnvEkouBRHRTYQmfLhFYCeG3vWnbme/NmV0d3cOY06zpnPo
dBYhD80ScI9tRH3VglUYLMbMjvGJJPqlLq4oy2PPBdLNt4cXF6kvsOoPfn+5+xs2
UT5n9DFkjZLFbOI46OxUQJP1NQNGWqlxPEP7ftOb3PfupGFpgd51txtYedZI8Sen
7OFEXIH3Uk53v3zGkXxztzljGJfQXFG1axLyrEOudv+nVF+bHIfVsHQFlWRQXxwY
nzScCKqP6WMVtcPyWOSiR1XSKlJKJy1r5/v0+tNug1uQ4sF6UEBLRDxn8xUN0eHm
wUHNl5+B4yzrYlsuQdWTgbjFRUzkikDQaeq5f1UqxxFJut6rTvopGpM8foX5ehU0
978VqUV6foOs90CNT3fa2QY3bhnWFQJWusySeMB6tJ2tTyC5in45nnew3dmNyGN5
3DnbIX/qEffG6l3TZjAljyigJG1F3l5LWMALdLO5zR2QgB5Lcrtv5WgcPHwrAJ32
l/L7lGr4/izkBrudTnB+cgA0dVyzzwZsc+hKDCZEikRLF79dtBuqGjr+NPYhZ/vV
FziuFaxbQMvHbwW0bWD+KMOah25lP/nJVi9BvoB/XXcew32R6qYCN8wqFpplSWIO
sElyJcLigGjlAVb1erttDazi520EM3006+uu52i8I0K0WM5rk89WO4nCh+UsWcxL
Rbbm8LrOjS7A9eINdbghbUuclDBvRPisQPQikH2aDtYvADC9xeaSJ1u7POLevCI5
92x/zSzj6J6P9XxV/32pu4MCSyNSRSd1Z6+UCP9BXtAISkurNuK9ezf2Rty7ZkOL
rTZp1PRkOJxU+gOOtrZ6Zcd79so1eAkoYPDBYso/CGaeyE+yeg3EfY9dsDYIH+ny
a1mX1TslxShOmMpdSQwDu3UXjnDzU7IoPqzgCVDZGimzdA12Cyl3aJutnz1zQpkQ
lTDCU6CAgys/E85lFsSPmBmFZ7oon/ySXPcbeceLG9IHW1ejWEoy+qx6qtRn2B7N
OlmQFS8/BhbGQHfqVTorfLL9QB+NwyEcUvRB6Kn4Sg0tg5+10Zbmm1Uhhqqv9Uq/
btO1ZB65lKpFXwG2s+jWbwzaMcM8eF/C3zzJt7kj7uCcfVfpNpOP0tQsqYulY3yi
aRGnn7ld49T0IxRWZ2Qprx3NG5DbK5iYyexdLt89HUbZpeVnt5HkCVYk+OxIdV8M
TiB85X6grSPTRyuCI5dZ2BLVsP9E1m0CxJpqjJm8DsxvZ0BnLSB7g2y5leu0LFeo
HKiWAjbB1alFI8VtRmTSZo022ihIzrukJcHk4IyvLpCeLbRjpjOa5Puxu7lAibb1
JyMQtzDrLTTRUTviWIYyY+lqQx3VKRHMaD79cDtchuy8e8ybVSxF3bRKWi0i3Ub7
GK5uQz+QJU+rSAPT1MAM5nqycl6CZ4aLs6On8Mz5iVWMkUFNCb1Nfk9naVosriKU
wwmqsZI6LwW1d5hZW4rHE9AIsRBHGfx+uT+9dXxPQIfUgnpTofJepAd5Kb8G2bpP
ht8G5EKAa1IXDdMLuekK9SHrxIJEdkp0xOXJLQQ57wKHxnK76THzSOhTi3GoQYV0
VyiyZchsnnW83I0IwVVV8JPibanAJR3czpo22jTxLm8KAmNiv/ko01VeWS3FHOhp
JhCMwioDCi24mC2r60xB7k8Rvlj9/Zjx1cC1MGgRP5okbnYExlocd7ZER8Tyx/BR
vbgIvqZX5ObjIWyo/udta43ibvCZz1fVbRk+3zUFm9o8LEyCvYOqwQoh3+4Xbo/Y
VZx030dzQ6i2PTgKfpl0JH0lg+gFvv49dNWLHgPdOwxfZw+MOqKQZF3PW6QvxWau
p+0x195XmAQliN9pgVE8rDRgJ3xqBkqnORBV6xgUJmOXGmZNFRU8VnqNuUrVu/iA
t8rxfpa6TCJVRvH///sNcHK4nqWX+ak7Xw/g5B/O8eBgQrCc6FhRGgNMt6SAx7OQ
LCUXohFizimGE3VFjydQKP9v1L0RvHM50H53UXGW3guTy3UZ7FDkL5m7/d1dBbec
khzCMkwfqHfTU/74Mlb2kf/mt1lvQjvWB3ygbyguNsTFrUpObPcTciDgoOV5SAYX
+/NVrisDGqwntXXeSiwZFDlAxcTp6Z2vTmfQKAt7qC4GrcHQ3Tn2uEjjKCW6iSKP
M+ZM3uuKGefZ0Vs98VVk0nOIH9LHF2+DIo2CiiJ+kxd2mHT40DKynLWvSIZjpvhA
HbIDTOoSAJzyzziK2zK44QFiz+pJYZzAM4wu7OIsDh1MAfPLww8AEW0gJzjfDVxR
o/S6ihkqb+TdKhrWHrSAQ8XnMoPE5AqgI3yqYha+7mKKbQ6ibK5XsdhRAV7cIaQe
NeXUTWX2L8SChJzrlO+WLpTxJJH8EWDUxz3+uUrvlV3jRv1NS92gcPIoxr2QxCkr
K+0PxNmu4XA9bqCIAc7iutbAxJBrw/LVYweSMfWEP0E+Q7RoeagwyWa4x2mg8HYE
EeSALqPibI+lDIM7R3EYjYcOdUTooNqO5j1Ly6Xxb891gmoWXbvtmJGO82aMjHsg
lzGdhrodzv9ruy1amfgBSSf2EJpBxGenmnQjKba+7PHUeFcFiLPNdb9P8pOb4Hym
qU0sQlzAWSQvhvg7fZMpi5DJF8PLhz11Sj1j/frQE2DOZDm5hykUC8LP0+QHgFLv
rBLTN0xd0+b0OqE3acEcekEfjevh3WNCJ2iRGmwZOyGEn6oAgVyCfz72rZI9cYsN
qy4Y7y3LB2ZThrnW3rvHzWJibIlqzJdaAbnMe6pWIEjdp+f4XlFVFISp/nKsEbaL
EDgjTVPpvLGRCzkBNMMPptUHegttQpH2MtQiQqZ2onVSulj0p0Ld6Puv++0yvf2Q
hICFYJZ90MTMwXRwAUU/T41OqhxLUh1eoke3fsYQ6fEQJKknM+CZf14w16N3pISb
QKDWSk67WTZi6xMPqNwdAgXCstXcd4wMftpI9EdrFfElFD0HXD8+gFVDxWvsVh7Z
hbBDl4m5aFHuFhB4mlASPb/QTex/pELCNgocu19vthnYIeBmawiwYyeMORjhSuii
iccQXRdHjx5Qen55C5rWr2L6eswC4OE9nbJv1pBJ0quVGfkHH5jxOi22RScv80GI
m3m2gR7pLpGwHKz5q+1L45SabJ96XFOcWEIiVl1e8zr5zx6uFtD2JuGps4sj2+IT
o4CNpGBSISXPVP3e/3VPBhNtirEgv+LTiuGh3EEJzUpT9kVLwX9HHkb5v9P5FhFa
RsYyTzhs/b3swo/vLw+7E42fGUdkd0Vf/UZl2BGTwBiTve68+IJI/cfClUHbdxAt
BMb/bBQ8Gn9LDLr7w2Cdrvgf0PK41XqlY8+M4A6E+S9kodNxxyZeVhh1ys/n7ZiS
RKNBL9QSjgk7vCna1V/wykz0Npk+koG5AqJPY11A8JI846tEj1YXh5EKyOtzl7wg
AouZh1NR6Ws2J8YotNNz48ISxkmdhgk6huwh16+pjJI0OHSWA89L8ZTMzUKoxENu
EA0iJvt3f2MVDRC5957WHaWzaDuf5nQs3kRml/f/f0jZglqkW3KHuOGgTQtEW9ge
DC1CrGa1EM0fszoZEr/tPK+1oCAWmh3FVB3fM5M66+l+EKLjZ+HXJdi8QzWxE9Le
5IIF78JmcDFSSo4n6IOOgLiqGeFX3Yb+7Ifls6R0NLz8USGSi7Dk8yPtVxSev6vU
alzm9jSgRpNJ9mq/ctS47yyvkO6Zh+d08NyNJ4s0cdPm7JOR96iU3A9knwf93XjH
FMlNrNIydwu4Ub3OjlInYuQCFCsC+OJFPUHAKV7+hpCg7qBgUfPgTYPs5tnC6O2n
+C0ysTTvnRCOG2VEudV6KyHoqhBRfP3BRkpdhqb/nwESb763xcEJKtMK17XVzBFt
nKkN51rJL88q23BjljUM9EFbAv9vgmt4jbdmv+TrQvuPa0ANLLB12f8jZLENNi+G
wgGLEvP07qlD0DHQtS9kkkuFbSavfTto2yeHn214RW+lh8BnF/ejmK+mtrSYE2hf
XF5grtuCWAIhcmDLzMtZpIGExJdZwbjcfHpa9m6sTghT3nTZZXiy0kWpegeLN5ED
r8LX7T8ILRFz8R/ae23f4c7xyP7sa/EFIRygwr6ns/HlqXALAzOQCY8tUn7a6vqp
B35QTgkViAl9VYecvLzmNto3sC1hr+ZHstB2wlzwwkBdEh0PlR13w8JY4T8D5HYs
twWxiJSbcsfenOVK4T4o7QSojq4Xn2OiNS7tZnuKQlLFkDGr2kTX0H8F5tcJJIiX
Y+HEC15PIbE7p50pN62+UxTYq/gL9iulJ1inFVn8AzwJaxp48/H2ojCubpKN0QOF
BfWnFn1a/MkDqZporG4BH/1tWvw5ni00e2EjxpUAVZCHlhPxmbmcWGJtyIoDq6+D
q19AUZXQMuRsHRQHnQ+PlNJKN5i3IjUFucTjQWXIFh+ulj6jLD+we9PZx2jFGjY5
9Vz7YfKA8nFspEJdfkzQ/Z+wkeripz30fhslQHW8F6Xo+CsRhiWDeQtsQQ570Bh9
DefZ4J9a8T0yUecA6ChzyLE8oVQZiIHFtLWYv3VhCGe0B7OqSRQwitXxOC88oSsb
J2Y8UNLFdlgtmFdAC9irF5hiC4JB57k1B0K6OcYTEXNi17DW2//id/gKq2Y7M/X0
BsnsgSsU1Ag++HwolF4LlLW6tpu8A+aKWs/1dZxdY38Naj+VSe0aXkKbYLKmoo3S
LyA1yIOnf4OJ+emB2/MWyeuBH8RU+QRMqZu/IrRvjQ4LNZVRpoud7dnYH4z5Ax3h
v9aR17V9ADZKZVBj0MNa6dsx6SG0nDGVHid9UU773hqnTu/XMuYziZLz6KaXEjrQ
7RXZKGf8qaK5Zp2trxrgU2FRxEQ2EU28rlJ2/H/fRgbcoA08Y8JjKPyk8jqbJjZg
wpYOnNVGUYmPs8rN7mO4jH6bd2FjSi23CSomCMYygL0egbBg9siUBKlXjONmDTl8
vIiX3DVitG229u+AHk3Kxo9oYtxPEX6bsSfUNwZWuMaW5U8prCFHcXab0Oaz/rBA
GuZ8zcqXhvjeOv/ZS6XHqG/orF/znajot/bt5NbpM4Naoiplxm6mavLVaSPaz1b1
PvtRxSYXvWl+KUHFCqhJgM6E51Q43YkW7VUdwepJVY8+sCGtM/cDb28vQjvSbgt0
mhu2p4PW0ZB0lL63EUjfOCbbyzqqbgIT84OEKqBu4Ki0CCqgpfti33voBxiXkv3u
wm1dvAXpMJ4lNC4GE4EORtob8SbT58n0eMMqlmTb/afn93s2+r8TGfBdoYm/xTVn
WsC546reJGtJgdvYM0AY44EoaEM9fDwEWkrFGrThczYkSMR1ziO8wXRkvCzajXPg
tpw+HrpmYUWbWu08rIIwBFXIBuJsIMWJ+s6DD3IpcCCotJjtzfG9uCskeEjZE/oK
lpulPP9w+mY4od64V/PS+WcxA1CwY/hVf1qIpSFBEk+TmSdvzXD+7eh4Qqo5sRdT
5vRYPy/7AwFTtSIiqsg2AlPgobntC9mdiw2EJrI/ryBuPISxe7rKLwHGpYJJswSJ
KO8fd9ArNEn5Luda7Uji/aNdKv8Gc0AQo83FRRObjIPu0L3kW73PnUvwBKpzBjXH
sFw5lUu8ZD4g7qo/xDG2wId+ppCtpijOQHjGASRFUhuZdVPA3xxX6XgT6e/KzfGB
Gj6dxbLrdi2g4Y8S3LXuM4ZZzM/56y7Jz9xQ6UHAN2QhQ6Kn1Rq86LrXXXpIe/yI
6W1qOgV99LwYr1xyX/pufITNHM+i+1zxclp7MwWatU/hkLZyIoNNYClKNx4kmrRP
/h/pWe5RMsJfvkmuRkqgyIVeXQFcTGJ/ENBzc7zxdm0tdTV/jzCDzM3ywH24EnYT
KLwrXn96PYYtSLlu1e/zNQ9DwTfmlZ9F7w+hkjvJeF3+KNrmRNxsO1I8y2ucZjZU
aom4Dt1YpvTIhpUY2vHHaa1aXsGlWhWsA5ahmOvkliDnMNgqB1XNh/YSXUvY66Xc
2hKPLa09yp56cS3unukoeNl10yCuaXSm9u3LFjP8IEpI2tdpVLIagSoEAMojh4Z0
sBydRGDanS0ra40epi+KlpOI/LaY5AM0u1uwVjY+P1cwFGZ33KjtDgpd+pda5PB1
FvH4ygeIUL1hznhKk33Am6vHMgHVikv6wFxU6Xe1Jc2ePNN1J10UHTVCpBurhGAr
EmOXVUG/SWzZnhLfeM3o9fnQ6+CaDxRcam6OmB2ZAIeRGDoh2l3v7WP7CqTMk2t/
gUE1tNWQ9RbcfB8Mv3sZlNAXrXm0wuZFMyPPkHjXnb3QtsHp625YRAOvUqY+2L6K
p/Tx6io+m1g52L02s1qIyyMSZ5P4Al3CR03qaOsT56HPHfWP3la55scyFo5VbY9Z
chME/8CWGbMZJIIPCsglwDphajJTC2e0F4is2aCNn/BRqCOxzmH9RjM9fMZvvnsG
7qgr+pRjdtODZieXt8egoi7C1tpB989U+CFQXHRpXvX+ZQ57wCGJ3EDPuKlF8UIY
2vA3CDM9G/QFWQE+fBoUi/0StQ3ZSi9n+1TsTTPqSoopDeNIHLqzjfwkcHphAOZo
RnlkB61B3hpQ0lIjf0EY8joIY8ZbVSNPXl/LuIAhX1zWuiBFMzV8KgbS2TE1lKJy
ViJ2yr+Xgrwt+4zseAjPplmAY2essy8wsUq1TsjX7+hPRamLgn947UzT9qBCD+gZ
7CbZRbZWjAaUzkQQxe6p9W2byGj0oZUbNtwGhsE5nNOyJfctC27CaHfiA2nt8UiD
kEkDS2YHMTYmmuvo8DsQA6o4GlLf3HR0D88gC+op75I/k57T5+W7tcM4won+jLvt
9TACPbrzMHcx5lNZ9U4SNrlnjODVHlbf+ZIujdlDL+freNpqulA2ezG4GeByjFC4
t7xdeC2V0zRaPNjAzk3tvy+33KXqKTMX38iPqhrs1KWqGmsxclCTIVeJKC+FDLl6
ZKvA6+msVal75bUtvCzSo0IDu5/l+AGoPQsPspS7Rng/8a6h3ERTgkH10SzSIt7K
3IGNKvs4sxVJbQmBBQyGw6dNiczFK8rGlol8w1azgopWu1OcO4ztsvm9hAeK50qi
o6bx0RgR7vNPdA7R5U6Pbz7kuK3xPf6kZrHXmx7GEyY16UvBisSc2Vp+1VLVgn+Z
eyQEcx186reLtit3DSQuk9ee3MQ3K3C2KTv4iqUe49/a9/uDOwRMOgRq0aPJjG+G
UtMEbiTFEx+OVIrQQSbN04cWfvc4FZwVnOba646h+H30J1z0hYCpdZGUZQJ5hNlX
nvS1qiqRsBbL64ZF/siXib88M9IWlU0YfY2mmYleMwNsGHIbRDGVczptH5IonhAb
S0bEPS93PloTULGFC3GsmvkGsRQUmWQbS8mK+dh0vV3jUmyG39wdqcKxb6cVD/Os
06Jf+ehavd9Q50OZF8B8kGErbYaKGk7SoKs9zp/CBU21/d7wmQpXOptjKDwad+BJ
O7X4P1PA1HOUzSQwjjHlckvUG0TE3QAcPHm5Y2kAbwGvc4t+m5A70+YiZMoKXxve
P2SzPQfs7hC3h+OAskXZJNvg6Lp3n7w3Z94sSIbGvaJ5MyPLrXCQcGzm/LZYnBC8
CKmMVY2QaSDhENKZh85hPEHcNorOPOJQWpDF5J6y2c4k3SF5drMCZ8xh5pJimwLX
VDyxACo3igPp33hpz+Dzq7iMtXVy12iMCU+HVgqo3elYG9HD1KK0AYp+bGI6eZAH
yIOnLadr/eebyoXAb/gAFeWAKsQ7v7f2x29qXZeTWoxQmKejPUMu3TYQ6aB+Uw7S
2Fv9JkQDYSvYpSSIeJFQmqSwtXc5iIgSQT47VJHmiPvQDHKjMpqDnmJgs9koAy3N
mAJfK1EjxRkRQG9QhW4ejd++ZrMMcWOmAKDb+ohwT2DuXayfREJTund6KHztpp7E
jkV/inziBEtAvSdqzDLIHlQipjpNvgBGCuzDs6SKRCwojSG/Qz8aX2Vmu2Vf8OQU
3p730v6cg8ehX+36Bd8xJYtcHLsJ0vJ0eA5EkgcOn7p6dhlVkhJkAhGql2SiCNEY
xorrEFdcXhD1QZiOZjIWtGdwGGRsFVzC+F9Qv7Pa74BstVvp+SydZHnzZgmtvZG4
vm9uC9bRv7EJFDphJ+H5ccManIkiYqwPT62yVzaoYLKS4Oys2sZgQOA1B29+29o3
wHkyaWercAFYqRtkgOzjrSfBs29ZdS6/QKb7EXquZ6OxyLT6/vGzb+hqw89HbAy/
Qwcb7W7x06wn4055F6ZM5hads2vY/Js/n6jwqg/Pbn2UAtwIbEYahPVqB4cWPA2f
H4l661D1Gkjb/ab6Rik1ZcQkeQs/66BlhsSwWMkctlK8q/F4hYwo2SCzocq7L2BP
eGRydC96JSJAVyFPTUD3Y/ffOLu0Dwe2XFsNXgt7MDq0iDI1FRUFbh0rHlz6A8Iw
2QcoM+Pe8DUObmaibMoN8BS6BdXREVWL9FOwY/lw81yQxHTg7fYgAkg3KTQFp6lw
hIg/aEBkTHtYHmTitgfLMM4dP/hBcW2sZF1xPbS/cazazJ+5h0sIMTV0T1o+5CXH
aktzgA0PWTXDjfmpG175UwYy1E0MxRM/hQDkk32fSRxeFUQZjiAWWguwxtA0xnZT
HWLRAZqT16EZYxfjE797kRWopDtdGMdXkHCHiWT+tcMsAgNVhoRdyPwYbTM9a2Pw
6i4yVn2KtWa7oGmUksFX+kq4kJgF1MJRlXfGWxlHJPwKDQLWSZmI2iqN7CqdulgI
dZuHXwVrBC6AE8NX8rtM01OZmSZoukLTVldklLLTLyQ/bO+7Re3pmLgFRAiTUcw+
dC3vBMYrI30ml+q3xAaORLqShXPd0cTWPfo7N1dkr3+gvxx2GDjrRk8B+9wCMaue
IivfGPSSPoCNNq9mOWfxF+TyOauwPnnAuYxdgYfRfVaDH+aOah8+vTdCCKK/+yTu
WtU2oqw7O2whTeE5GG8zN98ODdzcoD+QR5NTpgKpV7745fP9VFaY7vIs69Y4EOTk
4thKiZULGecKxz9mmYyXiHQ6AB+s25rmjLl75DOrOKCGyZ8/XtLkC95sA+tVnZD0
/PIN/Vroa7p0u3nxGTagetLecgLoLvYjcB5Na25l6aMcmY11emkYba/0XuRXK0dV
r0BTLwBqCEEgF3ry1aar8dAkl5R8wkP2JQewwO1kPfCgKWauchBAgTATO855zklJ
fTkFmwAjrhlniEHDdtTLuD0hr4T8rfORNf2dEN7kw0Af4hNbrb5pslbNp9ubsk8B
OsfpfWviRyE9IxwZlHMvAxQB2JPt/NOAqPuS3dJQ73MNjuaaJq/fg7WANTEscNhD
t+1u54qBCNGQjYTvzWJWSpZG1EtkENeljnIozrphbrM2GZ4qnwDTJTto2wzpOX+m
MLPq2sKSpgVe/1/XOSlLyNOP5BmSCX3fl0j9HVwIhJcbczQhtCZYT8HAyE0TO2Ow
b+gsvRwu3pgWgpAhMFGGxhYhLvg3UnN8lEJLA/Pvr9U/KXPIDC1tBZZVIvAf+F1P
fB63NVHtnXJS8USqcgd87BYYQd9e0aBL7Rz4CShxBA1+522wYlzUveTZU8Hxfaz4
Jr/Kp3h5Sh5x0p6FkEytNEgWMdAD0fK5TJeThqfpZtlbpqDuBIUmjXFlW/l06pbN
TNTogeYhcwGJW5zeYWj6Tt6MvGBEmKUfnSXt9VzzhNzXxaPsO9wGZznhGU+KMH8D
lHcMFMWxfGDeyw4WnofzwLK8GjOb+6KehCPGjK+42BAm+rnzVbpSe6eLvOpWt4AA
BHSiFhYGnvFFNbFGNGy6IrkRFpZahSVedIWMCsBmagstXSbRqrzH/6VeikRdJA0P
k76teTrvY3HlULfTiakVK0wBKbLjShKjLJc0ut3CyTOcm+i8DnkqeEPJMJQA4KAZ
wwG1e46gkSHtD+xqukIbN4ykWQvfI/MRer0q0xVLwuSHeRyXfgdlDVJbjmuWYNk7
EsvCJMWDTS4Q5LptnqA7OV7RmpoSrWnnhndBlhBotkCzTP+/4xHNvO79NUXwb3IC
/7e49z/+bRWjl1ZW6rAMvvsTWkTGYyuwNMPCvYuAV+gYS5IWmV0B5jcrunxSZzBY
y/H2ewB8FcrrRn9VpeTecV8W02XCnY/5h+Zwo2uWBFJdy9NAe4z9YPeJtWwjRSU1
o9ZY2coTITQ+yhCBXiB5Fnw1jizSjThNn8TQHOSI7QMdt+tAtNoS7Sl0EFXRuums
SSE9+TQ6JrEpst2QuUX+LtdV6dPLJKlG61ia00dcX5KIY2KmDsXS2Qtpa5Yf71I7
sO9qopNxjwYiSQHXEMgh2EdhoQBTjocTQqcclMaHuyRqQyvPQexAavKe+wDd6dxr
J/FwaKumjrticQaY/rZJl8rkHjOACe3U7SaG7oa3O9YM15kuJvGes82k7SX/f7I5
mNN5obRVcdn6f6r7A1xghVjKopXk42V5NYsZryefagIQ02fVGyNZkRZlQ4taUl0f
iY5EhQs2tx8UbYZEcSJx13g2NyVbx3BgJskG9p1A8DM48i8bgDXXUYFgQo9TE2p8
S9ySfESHGFlDHwbQsKI8LQ/nHJFxctj5rKjh6TJ0bYLTElqVnI7Dr2tLsQpp1meU
S9ykGUFm+euPESYAtE63HzzFgVX9lmLKKYI4r8CHH6pHqS1IsRMpqHkWHnpqoF+6
rhpbFeMbEXf/iybnGxnvRN+R4PQCy/GcDtnMz9pW6awEIbEVVsUjvLeaOHdT5lUl
V6azhyGndHuxXrJuoZ+f25H2M0uWwOlmWOy0WuoZiURZDwOPw1i4/oBVxn0CSX1d
R2dgw4lHX5gXpAFjKrrm1NfEobqUrOCLm8VlLilg05mOQGttxPKJvmGoA9HMVWGL
z86hmnFrWMKzJ1ejFMq97p1355ji8d5rzNN4+yEowsjnhFG7b5OjUf4Wfp1ayFT4
Jl0vknJiN1CbMzjWf9T1E0ZQsXWPrWdUyw9Qm4jloPMfFr291EhN4Are3lu3NN69
CoJCrnuLYblhufpzWjuv8thRX2LYaLiRvR1kmKcGp1+Dly9yoRIfTTZkzW/jVp39
+1SXkZ3dIVYQ/3TVhpfckWvpH8fR4jNW9dK5b0HVdvrvx+hJZrdW1K10VC5Ywdri
6eTzt5HojSFD7vLtdmf8STqNfkNIIkTiqRHDqER8/rl96l52c4pJseuGkf+ftrcb
2ogugkUpuWG67rG6DJ6YdmJWBxyVSBjXZWb5ztSIn9EK0Hbq6GP7qZP8LxBsOsXU
ZxfOfsSEcoJaC//KbmBImv/CtJ44gXbBUlARIzOogYeaIwtJpn+DZJ4CIkvVKPr2
ajHbJ8pQgO/e2B37Eav0eUXKuwm/Tmjx0Zjar4Dfgd4H0neWLt1HlfW1Vg7hJ2Ma
2/KcNmxN9xckmBkP10IJnI4wmQgXUMFuXIEgCN/8tCLjUMVzudZFBm/oew7WgN7/
eSZUE48ZLoW52ES0J1b/Jptq1LmkQiMemDPDIjbQcgRpnkwGZNoDMClLZ/bU6N++
OphyiEl7cb3ebK+Kz3dWkrFkOeA4U9zehIrJPilmaxtucusQKLGZcRIhK9KzpIJ0
b0Kevt9QT/YBhL6Mp59UOPKY+TvVIfDnGgoqEYcPD4OsykBjVEhbGT2/NQX/isjF
gLPPgOOcrik8MTuLahsOQ/DbXF2zjCF6gUePDTEW1EIWyPgoEO9RsBKCSa8pPnws
zb+lw2JQDLyKqJPJhGgctje45L6EKk+KVCuWGZwXwC2OWTBXUD9gNPtMsXyikwJi
YlXyOJzxiXsfqJAKGVE40g78xI6SeMrXNy8GLjGW5TF8E9MduUBDDkiWnZ4m8dc/
6XE4ujArIDOyZHHlZF2Awi4CxoAicuVS7K6xM9GdHy0ED7cFI0EDjP3yYPe/c3E2
6PqzUOzosiHCVjrVVn6uxI5fZk+JxNkGhZ4gxuZH8KDco7mlS4txhxuB9u5gte7z
+wKbJRTH7DeI63+Wck6jSvZRfNpApLLzi8d2ltfAVUscEaUXH+R5FUR71fGZ2T24
FJhtea9rj3SFH6431gFZ3XpGEjP+TyFm+v9hvk3ipla07pQ+HjCV2MJKWC8hWYzE
VM8ZWdJ1jR2QRvDk6jM1usCou7A+xkXgDqSj33dCZV7wHl9mVRMxYJHMycHcsROl
yRECHVrczP18VDXQs5sspMNGTh/HdF38H+5hckhvaDjAoRTOGSoHQRmjuAUexXJS
bA9IEhIkgA8iCoaH97couW9MXFwq5lpA2Gz86BlqEwTp2Vg0erFCExLQ3vmwqcsk
/OeJnBj9qY8zyMrQRc4VNY5pNCf2w3SE3HlJkV33sTJFdIcGYJopmIy8x6PHQt6o
H95Rgj5CNto3f60JCdhmY3o4LER9pI7ekylhR3yiOr1NBVLGARibcIha7s5Ggs6A
4ikHT4dCxF67U1UbwR9+Nt2GB81M7PuS2fFqupkg99d8zlhyljdluR9SWgjkUqCM
O1t5OPwvwAOINxlMTp3td4qanGmkMFoezt0jFHduJEKezHVZ+JrUIzvXHuNrPySH
A0Mmz/gY9n4nDgNaxUNrt+2eQhuMLFRt1aFWxFh0NgOYDZyNNOtwmCBG+FaK9+lH
iN7BGeDwOMrZKUnLH/x36jgvOnjtLwkV9kuQSLdsPCL1dP8bkNZyj1HTMfR2wHr6
/Zdd6DJzzVi4yF4QwHbiIBnTPda4jVRCpy6sAXWuLX6ZwGDhJDeMUSHXM6vFHxb4
it0HjJlvbuW/BEwzi5RHEnkiS3OwYU83E0cI1pBh7VQUoDevx40j842ADKDeO0qZ
+KV8LdXjHX3BC9eNg8KeRPWUJCEAw1UsrPv5B1hfGuSVKwJ1VXvSelJ+r2fKsVV/
btPHMjBlGtTHJmXNSwLaysyLM8x5CY2wOXflzv29/QMEFF4OCG4sEUtH4+OkjFDi
7Lk3XYQ2znkz3qd6LnnJjacPqN+ANq+CgiSxd5TqOXUCBj0mN9pFBBAtDDS1v34E
PXaAcRV3mM9Qlc0RzZv3dHvjAlMm0GzXmJhRTpnIia5xGUV37KfrVBjbz0CEXINp
pnmlC7uLKdemFu51VyElZTV7d2jfNAbl58P89w998VsHBsizcOwvvYIbnAWrQ5rK
NMrb9P7niE8omxHoYSir6KGFfuSlhjRhGltASFE3pId0JzHsnoeMOnkzdWkFvvKF
pZnirlBePbzjKXvAHsDajickyIP2YTmMYu1ocFmXBXDZ5rCmp9hhZgRgcVluQzhW
qMKC22qF519nwBWTFCT4lD0m1DYQ1adzRYxptfOaRwR7xthA+PUI3puBKqOjiIcm
RyfajtSH656g+3tulMQdt7QeSMyXRerb7WB3S/OleKJUbnb0OzKm86ByXOzOj5ES
sfZiM/KIcsp40GXfEvapNvP4VZimdr/k9EyfM2rDMrA1sKlIg6ue0PTGdcZbYtJu
ytK6HLCZ2P1Ik3vf0QLASpx44mxGGEyYEzKz/vdK6Q6ArG7bQFV2Dlhi4syotXNL
YkKx3JDbhuUJldL8oKs88TQt/6S/A7tcX1LrWN22yPYDBk95sRdgAnPbJstH58ZR
lGojhjGsl5sRlgQcODyd0WHB5ruayPSuIY5+wNlqmJ/qWiSz/BPCz/KuWeJrF3h4
jp1XKMwF8gr+7u0ObH2K+SComDNiCRxc+tOxKn7kjja89nL8lwgwcpZ5cKFg5wr8
M6/LDmNkWyiXn+KtAua4qHPoKKM6jEbI8KtlhecljqOerEqfTawU/Oa8Mpq8MbcC
sIHjQ/cgVbKp/bsvs1s/QCvU3FthLqjYY+mKobHJj+3fUkcPXkqh7a4QBir+jKNu
187aFHP8sC/wuvHJjmkPLDd+sFhnpcvVv9N3PKbQldFlXnK5f/XPUikmSoF1rZht
pY3FEYEyDck5/8fYb2ON5Eg6YW7Tcx7tIWhA2B/FpXq1Fu0MXzCn6de1vOZVhtsM
Hls0w0yNr4NiqEKrYkX/m/Gkt8Y4KZLeWDfDJzFsF93gOfEtNV+EcESnvQeCfYRc
OPlLEaoYkcZz4WErf0xlMuJ4gDfnPbGN24Kp2wv7fxBtVMyTTo8RBI+PUY4t/1z3
WXmLWJFwJiEJPUtOnwz/PkB2jC2luKncLAF6TJo5MPC+93Mgb5LZCGDRWFtWN8oe
hK4q23P/vP+5/9yvXmunyY3wqDYl8uwzdNFFd3AZcrkrykxOh1fHiKgc0/rIfA6Q
iZ2QT74cIlWNWKIpQ/b/JkVUz/YzjSoc1pZGx4MbJAwkI7D0SJ4MS4uYX2bFCXQr
KDHgl5DJsXS3dOGkS8/O0dG5rbESHTds1PtDUW0rAHujUKxs2dRASsACQY1VePhh
bN0YIlj26RRkFxGhpqAVrUGPrRQrh+xnL18h8Ar2WjvtRLMLi8/j5GRP5foUwf+U
yWBx5jl9Ra97I1bkfZzVjJJEy5hwfokcVzHhkTryyTk4PHG2CsHxJk5+toSXIM0Y
8wwN5Esj7Uk1Ik1C/8a7MPldZJN/B+oM+TpdzukLstKCbNUzoyMfooNhYbwIRUL0
Am77fXJrWE7z/ETSrSRrGMpvvbND4taYYtrPLIP/6ut+OfdWULoG/ZzVoqpYpAGw
EJM8D7Wk+q9ShR8j4Q1Fv8w6Da3jws6ygFyzBJZSoEcwW52tgUQi3U7Ic10C1WvI
mXdOX1ZwmbXrcGejTIwBEKdhEkJXPjBoeNzYkXH7nmJIbEDjuILJfNX2EQBi0GcD
gy9Bx28cFXQ3MiasnC/HJ7XOaDODNWI/kx+6SJVSGX1csJs8aHkB7g+7Y7j43T0f
VU+zjuyhb+RDgjdC5D6nNBCrywWVLzEOCI4nejzyt2eSsE7mszx5g5CD7AMVVg2D
VuoGlP93gpdJkx91823RiATAAAOgDefsQz9o3VFC/njEw0/e3UFA2VVMIkJrUhLs
y9VR4APTx8V4IMX4OfHcgb8j432P4Ag/l3AmdFvaJ8yuHzruqDBEp3L3IYUy6LJ+
2PxyByj4UFdxSURo5+9hEbQowmgNUEqHYWa46NevjFlv+JAK25/Lg/7qlaXBLe4f
seXNQyah9rblMHloC5Dl92mUldjoganzRvgIVqBHsaGAXc55IuWg0gXxZC6c1QFW
OzogDI+3awv8NJnbOCFT0X/Y6zOvWYSGQal17uUVDNSq9KMxk9aNuknfRln0bPJD
1zuWkILWAz8pwtIrQran3gfYxFR/XQb/9QlHzL1YviZufJ4sGhRua/a3tndElw/6
yukYR+51qMxA1zqatRt1l1yTCv9TwjoOufqpTgY/lNS9f4NWltyWbcKQtuOjhTk1
5VGaXTfGLGzPcn1Z167NLS4sLc0o6BIeJeIHHWxu35O6Jo8dKixyOjteHIGyzNJI
LAD5eIDrBDy+DEArj5FvFQ5KRRHh3vJf6SpSiScI/YCTv9QpCrxq7BVa/sdXzsAt
Kem+jACOjvxWCt+bOD/NbYvgDHc9sF1y6RXaijYxUhbzEZJOERvMRoTIOFshgZ/F
hlSLrd/qPhf4SANAb+eKr77Gb/HBmP/uK1CiBQZHvpQgS389h63uarvg3cMhVK1i
jhSDch12S0d4mWXmopiyqo6/l4m8Euabb2aqhwg/uVwMVOD6pxQx2zqnYqHlJ0t1
d7rA+koHzFVIz1PcdoLuwyswJ02tg//QI6E22P+9YbCoiaigaBlZ1KFW82f45zd8
h8aZS5uqYNOaMwd1xtj6y7uPVmWORSH0G1yZz8mplFAdY3BWbNspAJJz/lO43czE
yyw6WinrH/Mi5ISwkawS7pNNQtcz3YCuNhaFv1l7EGxzNYygLstbcvPhYOrXNYVq
TvbQoZFkMkmBOr1r1dZcB1au2FzUxexMOjpWJLIuAYKf2Zw4e01gWs6mh6g8v1ie
nfyEPKdqtKLg+1SqdHkd6e1XZJUyZLHxO4mvyelTaJwpLF9OWzpYFzJx/hH5iPc6
0Xt6T0mTCsX9Bi6SVRWsUWsmdbZqaZDH8ow1DFlBVbOFGgMRZwo0/KIp/dmLQD6t
PCf9B7HkBe9337IlL6PCXA/MHuGjWD4KqkXBc37ylwaU+2hUuUDlNh0UD2kVjhtY
6BAjmHKT8H/utICNoWdbIyXqRkYtLwgf/YXfTa5hYayc6g20ZnLVcZhtb9EjRWkn
r+mJEwCUBmD+TO0O/P8MpMdSBnpISOmQ51YisTgIFQdyxXgf2GIC+8NGvNUJotUP
hjftnZ6BhRvV4pjHAe5Q3mKSYZXqGx8f6bRlJfHQg9w6ZF9iuGAwCAe6Rd5vAp5E
dk+gdbFlv004/bhgZfYCOX8PkgLA+VXR8jVGuWMXaLrqwN08uugg4GE6BjDEeTKr
akO3NeP281saLmHPVcnolmcA0pByDPXAN7NcIppG3ZlbeOj3jpJ7YlGVTtKBkUYR
9jYGbWIzu0S172IHTdoruJKVPNgrCWHMTMKFRLSIf9YaKnbCH6lE4pmtgdG3kORH
IgELYMB7DcHM14rh12THrdbo0MJ8hyaWV+gEcpQn2OnUyGWLvUE/gid1tyEQH7Ow
K/7TvLPWXq8rxG8xnlLCAhEY3EgRnHgnacgo1uX7vdq/4pzdLwi7n10CE7xshC3u
XSMv4rCwv4HMehZZqik/VhEhexBlxsXyGLV/jxJDCB4RgqOIYIttNDhkZzx/9ydD
5rgUBu/NfdydoxyKqA8dFlS3omDi5R6UTsAHhpuIxMzCVfLM3IiY2oV5N2os8Pbe
7iKIj1/IeLGLIhc/AKCEA/cb8y1ZhoSBWXUTC9FX8Qzx38gCZocpOsmzVOzGstcO
MOOcjg0cVMIyJF0YVJg5kVraA1kPg2yQSP8jN8+EyzFILw0TeSa3dSGFWMviC0/S
ghfzcWeeltjS1RHrwwv4QsbSqeIXkWlLpf7VLpUYkfJf7AcVFXmwBhmNFzx7aE7Q
uxeO7Xnw+tZ9SQIp3LWufrp2dAqOHiKyA8LrrAFmzu+TdN71xSmJcla8A7sOnIWc
SQdwPE2wZhFxRFHLpIkqrG0L66z3urtk2eUXH8JzqOTiUzEStmasADt6qwuG6ki1
/aYNbv2ouVfRvQytVc8IPZqV9OwWLGQcgJYUWjpSuNeTQQA6WngcOIL3YcQFwatm
KM6dhigZ78xJsy73PE7FByHHALwpH7c3yEnqgtvOD1kujAFNDPxKnOFPfFVOyA6T
9bdeR5amdsb+0Lmj9vpmtaC7r7Uhnuq7tm/SkrtZIM1gq+bgrmLTBDsyIhNT3kWQ
RztxmU+p49eih53a8RB3NaizFgM0jZlooVDV0HKhz5ufaoqTvkiNoC9uWlFK/pwg
MoxU1K1DzEEJE89Ft/0g7OO1kG8p+TLWa7k64lmpiv20zyXOqW61I6cEeFULWQif
u1pN5EI46Sigx6OwA3bcdmobnyca3T0a8LndOGYatQ6H2Dw7+mUAF71NqhJHwdz6
b6FNkYE4R24XrhPPxIakGOwSKwGQqMLd7IbZ9oJlhyAE6a2HhuXqqCwkZQpHEyV7
PULEE3g91x3rXUskZUISMKeF4f/PaK2sNzcGgulyxV0DHa7qaf93BQ6gqg6I+Vau
6udZ5UYnDFgvDb0bhy21VPZQkMM0sEc+Cv3bFXumNklQlRb4z1q0ay96HC99WTdZ
x1eUPfejFkaw9NtxoNtPY8O0XSQm1dFpngUUmbT3XHbncwj1g5BGYTZ9v7vY8OrU
3Vi3npsniovYwAPQQ7NVv2YAAZhHpqGtLyJyTzDSVo7U0+igYN4NRYLTZTnC3fsF
UhNczw7kzdgYIyfCDogwh07NH54AfZBgd0Ue/8oICrU5uP53wA+zzJXwk9tGnTav
B2BjWpwSHa1fGegtfKu+7mw2mygee4cLt25AEyDp71uqRxojg+r62Wc/YRA+yTID
iRxjzy6JYNLHx9ETVy1Mf+6v1NcEnSpz27O8VoNVdUhdc3Co410+uulV9J7F+j1U
KPu6EoyHgvoRuPBnOvypSxe1GwDZ+Dv/jfeG6TOu8ceBJwKqQN98W2FF+b05+zxn
MW/Cyh+6EE/P34fET+sXWifbOnbCPCqt/Nh6TBw5C4olPNabhljHFWFzVShu8u0z
sh+ZtOSz8TrBfilpTqZLxIN5dp++yIpo1pFMUx6U/BIqSqCsaPuFP8OWTPpvWFCY
9DbYNonRQSI5WaiYKZ5BgPohcK7k3rbpfpgKbw8SpXEx8Dcwc0Mm/s/Oe59zUUuZ
ph5xc/iFGZb/Z93xTaoKjML254lwTXSwsBRoiZ94FnIJx7jaLbNxvZiN5ydRR0gQ
dSGiXgYoggRULtYKpkvAnnFeHplxj3SHWOGneiGcF0ReveotLR2NECO869/wmuD9
rd8wNXwpBgG26HN1E2rfPfFDw8rKpLtV/lWD/4UhWcwCQ6hP+YdSCitLOIbsF6UC
ZyQBeBVmfp4JiAfMMGyNc4EL0mhoTg33Y2Tb0PBnPcdDEx847ixjbHPzPIAs+kvK
bcgaDMSFT8AK4BuXlBM/HmscEZGXAT4eaaPP9WO6k+fR1UQCe1+Ghcj/rUSEOj6v
S/UpcGleKQHJMqwIJ2GJAQiJJ6B+y/IKGk4Ort/naXJAIezcmM0q9+AsKicBbZak
iymjon1nnsWje1xUMhyYOwn2zkYRLccAs62rBawYuOXjZqpNCboTX63B5saw5iLM
WirFMBHisLESYt5+Tf5T4IHFreRB1uB93klGee9lvLXvZNcBHtseC0OxvZDeucKL
nPCuZsoLJLtnUU2aeatuw9XKPihEMPukeToE466zyuRLER8C5VWQCZi5aOU2FDa6
FyVofVJSi8QXoJqZHTt8Fv+9iUuSLvkH3qsHUAWOpJdHP7aAYetbE8oaqAkXUUSd
cEhjHK/l/WxELpLv6CkewhXI4sCZN97FkNMvmlSVO4XgujSggIFj3aXKfqmEZfHO
zJYsKqDF7sdPNBgBODJx6QF8rJLQOtZySgpf0Sy5gtU4Pasuwn2BkuzrlqMGja2q
fIFITwl0rNiZ6tlOG5lld7YV3rqLLealC27w4VCEgMwzwKsYR0biVL+OQ1RWevKb
rOP3+q6wp6+9Qtul67i+UJ6Y/aDNV3u+gvisShDZOGQZkYxe7nDP5cp+REZnexOr
vVm9w8s+pB4SKusZCtaVITZao25wBYvNQDp5H3KMDieil+gOxHovspDIHWx19g+L
/By6ZWKb4c1aPT22VYRL1tDbooKqNx/oBprqYY0T+6JXfYCT8ARkMLsjr6uUu1mv
VKMAcdhRSgY5YtMJ+IR4IYkl81voGbMvUWTE99BiwayLrZLz90dxjzgBtX4Y0lwR
X13TRWy9JLd7P1Fisxj4pjLSxzITZLxtqwwz91D4/71/SPn/4xAGd9W2d3H86DjG
6u9Hd07ZKYDURj9nYz6ZI6/66QeC3XNEg/vwNsJz3kHtyo+IUEN6jYiFysJebkYL
jDqJelPy3bd/+VdBDrxPrNNnyJSwcP9peBKjEUWiS3UbnKasSVgR3yy0XoL1CqZ4
zROamwSaf2OkRhFVZGHeNRaZBNHY6wbLhlsm3FMn1FQfpsLlYwf8vTYXo6TC2/K0
yn+pCacqviaDNxxY+CliCaoH52iGnQVQPJTBCoiKBVaX8wwouk1dymRvPWL6iGKX
2ttTptildugMHLx56TaUs7o97oNL7Qsa/47sJwMwCEeZrErI/X1NPz5wVe+nNM/g
JAP3zfjU6bmwk3qbj0ALJtZJwCxvL8DrwmWHPjUMsq7CNBMtHzSnhQlEW6VHmgJL
3QPTi9NsP6srYu5/G5SidtgawAMFc9QzTos6axKE0ai0fk8U+nH/FBsG4YWJMTf5
qe2t7WWVUs4H8DgjtqczDMV/DVpOFAxsbR4HPiwPWGzj+8QlvZOCLDaT452UgUv+
2ivV9YEreyYbfbHeCASBKdxx2xEzn0ZYBcha5IsdzL8/a/Q1a9GDJ4FyFBB+twr4
BLAwKMqHx5JZX4/IZGz00jlkEXQcq6cFWnBHFuUYkXAHJOerdOdTF6DWMBAMkyLe
LVtAR9yrNMcDI9fA6bpENdbtfM0Htas8PEUZbw7SEsqOjNKIRrfmtCTBw/3/rLO2
mwLiNcStY3q3ZJZhTCJz/gymvXr19XknUtPIt8NX6u6azLsk8tMhfjuwj4MRLHdZ
D99ySD3VnC+qs69vKHZ3EdH28J8m2VBZK/lbP+OBIGL879yEsgwdgWQBCz54pqQv
0LNTRLsXi/AwXetKeLyWJr+CwItD+SvGSoHxxJPSjiyd7BwIr5y3OAG4qvy1i0lI
o9SI2fMUHwzYBZkM+fajpPuwLZun9SSygOwMlFTyOLpYCHFoTU9udhoLNERvRMcs
1AoJ3EHD3C6nuDFa0lt/hMlL44sKns9VU2fctz6Oy68jGwOYoi3CzIgQG3vJloWn
gz5/8C6DR7W7aIT7JRcfzXRCk2Vl22c+gowyLQq+XaCgW815J8cRUKhxkrwsDGie
CO9vsQ37CnSqYtSfSqmuppyuYNbejV1tL9pxzpiBOXDeOMuW7+e83pu5rcnjB3jA
qEUM4BFz9e1YfWNj9yL5DXHyrGhKSl+9+aagFlJuBEIkiA/4o+eBAk2wjgp1yVcs
D4eafNJVWCV7f1EHWi1hYOg96gdI4yWxCri4alwG/P8v3lLFtY8hCkX2G2G2Zoix
F271ZF2IJFg3L7y1wVYDHxio0y87q6rMzq33eKvjPxZQVTEeVnT7rsTlSSw/xB7R
/FWTsy1MRGRbtJ/p6MBXPZ4XkS164Uo+ci5Jsx+K5qtaqn+4DtQIkQxDXFb6v+m8
YcAa1UEIAgGjhQNiusfh/FVtHXK8BzGGaYVrV1MDRujUnPiax3QODrRZLjME76CX
P1r00qa3UMTLWx6SIoOZJomcnrjpJndIVu57IIq8K8LZlKIc7zjZUj43tE2yBpTa
nOBVMk/G4z9yq/TJLRA/Htx5EOmC8xOVsAqWz4bYWGYBdbDYW5usNV5fbszDXLnR
3uNfNl/jm9PoCpAsSC2K1CnX8bMpGGSp3xXAxkuJv2OWcCzb6Lxz98xsX9QN9DmK
+kmEZOOxiBfugbW53DnTXdso2CztcNWrwI1Q9r+AAuNjF0Yy/MvLKeWINBrODaOk
p6jikRPeWKY+PKcM1SnmTWtj2QMXYitxn9G7u5eUkeAjZTtDY7uhv6IrOpAIb+vz
vlhAvNXVwu+OLDZbzLweKHlxt5eVMlv0eb9lh+8BosrXX0N0RDX4Z5CL4mMdebs/
lDjx7cuIWOsxsTdVRrmoCwcNSXfUp7BcpMMNU1+t6n4FGjIgNaqMpkBkbx4jeU7/
sE5wN1SL+pLMWq4/OGTIcp5tCAVSytZqB4BgZR9SscKnI2g6MWXKt6cDMT4bqntd
qV094UoGuc3Q6+rCiitGUghFF4ZBU5qDpma35jYVuFbyxnzUluouhLLXR691+0UL
/rJupHyGTyEIYl7AQr+PmcveLTkqxcJ1/vcOgpFoL+3AaqQwdyHYQ/Mo4hGz4XrG
X1Xurri+IPlekbv1gV9HBv+tYnbyhfan553iHirNEhG3ZKSneEJ+6db8ua5j0vR7
55wOcv9f+prqKptzipAc2QgIk46unHz3k85sgdm1XJSX6D/td+pDkre0WoSLY/MY
Om9kM7MkmlHtxlHs6sSh/4JrG4jUNv+DebNSpFVj7twLDD42j1fx5IzKFr4PnsI1
XFBMP1KcA3o+a1LasTlwDH03TP0+/3Wtjk8Is7F5TDHp7N7NG+aj+YoC8D54jJX7
45AnjJJ9uLV9jkZeMN/I7WEbgmSdNu2+gFZi1/WJHcaK/+dmG8LATeaQOwjhwtJq
lrvaIl48kf35k2oN8L0IaqD2NmEFf4yb4ll6j3aLKPpI9r7uu3T8KcMSMnW6VylG
Cjx44zKRe/AvUAVRO7MbKLpIHzgW65B1RSfVoVkUu2Bdy25alhRj+Np0okiCt7Vz
OxEWde49ouGaMToGn0jIivPscPH4jRwYi+VoSrqEbCUceV6A2okexzP8VYPVweju
brRAa7RIhXlN1cGB+GY+/n21NmOSY5EDudGkqqrL6yPJGkhYLh4tAynWnLKcGzae
gEiE430xO5oGDddTRzwWXo8ScHrKnz8FW4ORLHWxybm1P9WRuhsSww/wLpoFQaT7
mRBw3GGnsD1sieBZDYr44/ANC6gwqa79PPtEgBFqCT1JFj6FNLsHUX4pmjNTP1Kx
SOIyCihHG3k5EyOev/okH5Y8eXAiJkCBKWiRqRN+s0tPijcjcDL24Pt9YnZPH/lT
J1HKcGJh73uX6+0yXO6TOJ+QaqopnPAhCknMACsx0VYI3HIXds/oKO4ji/0JRFhX
JbeFZgQS2zsQW0IrMxPLEvj3Rlqwh2ZXr0Z40l8GM8Az/9dexaRi3TSA6Hwn8HnH
iL36Dq/10Jn9gjGEXRGmh458kS0W907+RzGvRgVd2IWBHBolUZ1Ob2DryuUU2T1a
Fc5DRuEiPbg2dJY3QFbRXv1WvHLiYirN45SoBLqpmyBcWNpU34cM7hDHXePVpD58
s79Eh3Hg/4rawbxoY0E7pFkmH5QeLtK5HPu+Fhnox//2QdxjoFR5/7WAd5+3SmlF
hs/TactzhJRBngUbrmKJTiD4zevO3BrotxIgw5cLsv9ev5shWimcP8p6nP7BtSPR
pkeHuN8Iw1PZwpMR3LfyTeILDhrghMkzQ7+YpqE4k77dvJSz9J6OD5fKlFS+VFze
kGWlBthy+xN0UaRiAIc868ZONp0z14nktlWB9RvK5p77cvlScT//pkPHPrmcVZv4
GWNxjnnHzZz124IOFqhRlkkbLB29NGein8yvJ5nCGBOZmtUn5l629RK8+/N7/akY
eKMoDN0SlfS/mxemzn4r9QWL/V++GYa0M2pX4EYuj+6TZNuszqWJ/aosqb8kILRt
+lb5hJnUNenie/g27MvQkLYR7+VRsS9CO0KMffMXcAto3WDyCDBR02cmLdQVYSnj
i9GP3RiUNv94i+eH4WC432NmdKFrUZXaQQvGKxIrTnM5VOCKJCDBA2ZSYxkQwX/N
3UO0BxYutHeYYPu6kCRy384rM1NtAkz0HxwhJo07VWR2Fy3moLC7pezDg+cTnubd
+APmVUmb/FDLmOJKBkn3xpQ7bMkzCA3gVoCErBzTL3WfumpQzA5DXCoIT5+BRz+D
bii+NH1axqgmYkXWJ8Zlpm3h4e65JmxhM5i6/ytTZHT7kEKdlLFsOqCmNBXs5a6x
4a7rBlbk6guhx+ESMy5JfAs+TEYhZdREk50TJS5ENr8Rh4NNlWwT/qIhXGQ2aWTG
P0V0ok198k1Eg4GjODCK8C+IzAUXbu7/O2MORJ/OuGUTa17A14dRbjb5Q9r8tpsC
HshnZ4QJBDW12IK3AXBYVpsqy+vQCypecte/bIhzmSofznBbtK9lxYLvbBAfgPvI
PZyovv+nPmE0yu057G15nHF+4xNKp5Bvhs9lJ05cm23KedrOnC/FLfztAvLVpSZb
QJJGlgF8rB2rssGHkHdwGi0jAig1oM6J+YXZODR6OYdHvXkgph44YEStMlq7KbtH
eO4Q389+Vy7gzScsNYjh0ZNDSUqgwNFHF6dg0YPQMw+N2ihGFX1hH9YUPMVaR0oy
SvzOU16d483tzyL4XJGS9rnQkDrhG4GFUxSzjq24UF4Jb3t9nECXS4g/DEdMSLHb
o3w1wvgpp7rE4nImrRPJoFAsCgLFGRoOrw1kVIX+DmoNsiwAYujrZbnvo07qJJNB
iP6PVfAECgulYjjBD1SVrXi9qIlC3zup9pDlOVbxFFlwK7ib6K+jOAiLFOYrmROA
M/aML5rbNYJbGFD8c5AO69mTL9q5G7ZAyX3QaLXym901uuMnDdo5Z3PZQ0CfPxcJ
x/xl2BM6MbuXNi18r8ZWJP/I7gvgBsXFb2MHwOvD80y/o7CEzlrEMB6t0MEjgng5
GtoqK2xqblbTEqT0V7iOmbF9J0ZHOPwYrq0cBIpVHdd/FhZcojow2yUSnc7XIb4B
DI7T8KTrX8I5Qwg047lVqIGnnd7OBSukZCx1M/AgPNsp31rYF0oTJ80b/TUqt5Yf
tXOXzslgi3efWnWaz5EhjkEAtlDErd9N2NR/JRMufResqW9j22EzwUNGyc27TBVe
O5EWD63ko2O2E+yr+QfiS1Dabz9JO/yA8OdP7Qt5X3aDAt8Fhg90xmGFU6LtFiUP
4BjSbQjQCtrHWdmpQy9JiqY2ADGDjFEJ7DUisuE07gJiYv1fKBE68gTVXqqxIDkM
uv3hwleoePnOwpuRSBOueFCtAl49GS9fxj8ZUbH+MTpGhJT3AZ21ZbiYmd4hJYBz
szR9KLPL00plX1MEcs+E1FRPVoKusiq8GFoNOCyI0SiAwFcSC2Wq5HazRvhjQf66
A09HLT/jP9BYgjAAmx9w06tnaikAC7UOapMN/O/dj6LaJf4oKHA5RztbdcMl/gEy
pp1U+z+0njG39GadxUVZ9ATHO0hNu5XunCAof1tDZqVh4MjCTx8iDAMiqLvcAbMT
Tv4+HUGapvATpcnYSvM9uLLvk3HceSJ0UV01UGpbZuyMLhwNT40dE/1ceew1K204
jR4eIexDPHxGjkQ7cId7zhSvAqbXnjMaljBlLzKYYiXMcoWKdoxA/3ny7zQAtIlT
tsClwh0ko1WU3onAmHudOkCcuaRJ6zrAWUy/6WCo5/wn5tS7E9pAjUfBWIIAZPf4
wdXKAHNOpHn1SI+fZq6MQq/lzLceAjxWK0O96dRqG/mvgdKWNmNBFz36SLSQJexT
3r3g0i5YxArcn2OWMlRftO2Aol0HN0oVCU6gaIBzYr82cyoQ9SjVnpniPPGVnZbC
pI9IJXRKRSuitxpyhxL0apQFfVdljI1PtpnhdUtml+TBy3LN6WZzExRInO38Uk+J
e8vkNIuPxx7d7xHvxVdb2B9IC4TSRCz+5DXLcCXKUx526ej2hTo7FQiE786tAz8B
eJBnptI2cLDqHWSD6cLcmWFSRJVhyB9O972PPAekOHIWmxSx8Map4jDzC1Q7rPHQ
OmGD2WE701gCZGusIOomBmjdKItczzUMfmqdovLfMmh3gkXbry9vXuwXTfW3mWh8
tnSp7xZCT8l1ilBmazUejy1gUwvV6TB0+Cl4691vu3o3dBYBpm9zwCYR139+hlEe
XT2Zlx8lmcGMk7Y98VL/e2FvscX0IZWHyKB5nEGT/9c2vHXhV9bwBG/9hSWSNkpk
drqr9x2mpirahYpLSXLvvNc7xS3cANqyzNLiYpyspr/MPNH7fs7iiZpbH6G/Sf24
XXZcVulCIJHGwIihWY8iMR2Jq1rrrOFZlV5FfJ4coaFFsz+U5Om0zUJ3bh7nHV6S
uG+E/JZQPFdwhg36zrddS2ML9szf2cJBS5tF48W0vrPfNLV0xG/fAmXT59rt8+vR
b9KQIflKyGJPCDslXzpv66TIXZHj46aPXFmZLS0hxo0D2ZJgI/zfwIVQ7zL2EiYv
y3caApLDhKGHy5v65FTaz7xiu46WB+KyCGXFRFKeYgfXYVG60lkNvCpGvMhU0Vkg
TFScLenSC45Pjk/wnRk1UCQIy/Ny1pZzTgqSL30lYgOJX0w16SDa6zuWM8BWWlgx
NWqkxAnzg2/gwww5t83XlicG9QRF1JL9Q88mOCRF9v729p6eNBB1DWnfUBwV4p1T
ULKMtuYbz+d6soz/tEN3rLda54o/HBA1F5F4SBkEAo8iFOqmdorvnB0DYCi1h5GZ
dAjwTxQEIfiJreL86sWUyQ/u9Fn2wDYcxpfHKhRhJqiRfRA9dsBKSiLPzn5IrolM
wVnwt7Pzf15hNEnnu4zJJhrmOy1kS3koPGaOuvMhqD+FgjeWPJV5JnwlLgk4HD8f
7HYaqqArunmMikuKZx4ZwgvKLIfEOqJl1sBg+7LgflwXSz5oyVnfjbU9/Mwd3Fj9
To7vxwHulPMfifHKkjc1zmxXd3+1Fem7UKV7xW9LNhHSKPwRkI8/Mp6pXUlvrKtR
Gavvb5euWEq7Ucux2sBJUJ6Qehphi6+wNcpBDb5k35Cb0W6ed/J67KlMUS/atYQ2
p73c6MOdVsvXWF8H69L2Yo7d/x4T/+YlKyaz/nI3aIL3hW67yYefFio0QKWUqPbe
qkJDNP5xi1x45GKRT/UC+YuR0C8jTuteSoyyI6fozBHOu/zSYodI+mS/vjdYWa3J
k4vhvvlyBc8IOXfIQiHwRHtWTQhqCa3qfp2TLzp3/M1XfO1nLIwgk5hsoLWLhD6Q
q1MwPCMBRK1GKLChaCxTdBElEhJDbAOxTAVuMbf6N4I6nK1ZmHePKrghrO4cKPE+
AK+rKyK0PoPrQPOdVxlkQAXh5qiQ/ydo4ZfRDowefhx85Ev3n6rCMk4VZuBsZNAK
02342j/GcRu0mkNIQDDfdgnuinVehBRyJ9aFyVa2mDmAwGFrFJOyAHyRXoSFXthf
Z7RwOan9/2lGeAa2UZGJyya823/eFtii/TyygRGj4Cy1kVrdaq+j6qnQsJeYezir
BfL6HM+HGxZMGonxk9nLpJbUNi+k4bjUIfYjuNZkJs4UVdnM4zCSrdljvsPqJa8/
vqyYAP939eRRcNUp1ZEjU9BGUz/bd5IVXladYK3lP9ZZxwlpXx19JwWGcPoMX1l2
pkV2SwMS9/ZmmxvVN6t3HlLvRiYqexJcDI+l+9kLUCzh4ry3+VUtg4VahmtjRMtV
JN87Rwq/T8RQ42at9LX2JH80GMGD8omxhdp0KTTCFAE6eFV309pbDmikAWAT5ujf
I7Q6dsgiXWH0v27lCxQG0M6YDOkNWryWIpel77KCr7alTTiQX945MgQzAzuQ2Po5
6SoFtxppmkZhzruUAgOwaZvaxjBzsIVQysreiCiq9MoLzo4VEL9GTaMQlxo/56mK
sVx4/0tSxXElLQV2RkRXDiVCX+E4dOgcqtMMQ2ItJJ43RjCZFxMbeHgFv0ohaPSX
sJm1jlkIX+MCRrVJJ+eXZyfSjzOW0gM0j/RkU9DZQHPMlNKqcuT0NBij3U9zEQ2O
m90KIhjAPQMPBI+pIGG2/fynjKrUIUS+2iUhQhw4MSPOOQ2Xlv1IkVHn9g01YFlu
F7sp5P2rVBA4VJGsZ6fn9iYdhSoDXGJD+ROjEdKevqD7fgc3PrL0IV+Y1NrFU9oK
ygi4zLm12HYbc2Pr85oczVBAVLHYFM47tiOll238stAtxkwMrN6wchTpfgjcQRN7
mvr0+kvvaL4z4+jxFDrdMEc6MHp8QAyIDALF40PhUDiOq/o/e2fLmXVLW9fjP/d/
pTlxnnuWNLas7/brFxPjIZrFYAziIZww4h0fKCb7qU/0QN9zftG3g2xoCh1UHy6s
PbtwtEXOSOweEg9wMaO7pZM0QirJmcpjXA2rQNOH0jG+kU4GtawLHBLOBIwAVNjf
AnUBlH7jQHcvDw9qZ13nHP2sc4bno9ZIYuWS3Wfdokmq/wnoafeGUjL6jMDAj5P+
uL3Chrezoa5tLMM93h56FY1IbaiRBIjRIDLo4S++0pY+62Ux3HCSlhAW58m7ESnz
LyJYKzVhtEpMjAchc9z4GK5wtOJqtMQJg5KT0Uf2e9EynslhOieibQewvvxuZyIz
RiqlICe/TSZm9QrszrNlX+lvSTSjoNO9i2UerG93Sy44H3rGku9RGwrfD2F2N8je
LdYgvQibEVie1t573dvXXwGnIexCsavYJWPKdgGdy8zhJKADJIRsGIxK/dw4Nvae
Csv19ksM76EW/o3AuL4lUQMVJc6xYnpqmASCt7tk2M3Oxu+d9F3f10O+NelqFag1
RnGJqDnoBK1hGFDrcs/rgPw9mfht71Nd9FiFgrpmBsojSQGFpK7/HcNFec55hN5+
ViyNSuO7jmsMgBXX0MO0MSLYRv6qMsE/vS9Z/o3ORlZ73GK76oXr1FBYbdONdv5k
LQ10xsrxBiBl+Tn2G5SdHE3AZzkO2Ol/EL3AuipTxCRlePnvwtQuQMRf1fLo5ccr
vEPmFLLBGESLgwVMOoyCXp3jKOmg70lbLkkDbXBzY107IjqsOUHFSbiyo9xV87s2
1vGmd2E0JyFTdAVdN+ikHhav0CNc68bTI5ytkPx+nFTaiqh37TJaFbYVO+ehtbg9
L9vU/4SdRan6/RrwZYTx5DxQvITOzcu6/mq38qnRuNX8EE/ftv+DYWkSwwU9aQvg
+B+rIU21G1J7J5tqJj9Z1gNqrLum213pCbhm6yVVdcMzUUyKJmlcDgRCdT6CLmcv
Q/8fr+qpNAqFhlI2PZST2WrtNbbcDpgAP64c0aTAwjfdNwxayqjstmDwSuzfp6vP
5C7P7aVc7BUFEXvTZr3Kx/jRru/QJpMb9Y9eTlmyiduMDDiSXzPlJSL2DSz88x12
tUmPjPQ0RJgQXL6BKOp7BQfwPL8g781VbkKOoudOlawpHiH4E6CH+N5018yx/z3K
ir4p1jULJtF0LZRk8lpEM1RuXOlycqsYkssAWWylIVIfgznPE0Ga6Fxg9kleyJgj
K6idyVUui2gQh2KC9wWKTHRLVQVeL8iNgShk7kDWgU8DyuoIUCbvjuYfEk8AT5fd
IfbO4L42zTaTo4VhRrbD2KsWVgB7J7ALd8XrZV+1Ub6lJAbGfzriqwS5iJxe7jg6
aCiAmCCLo4tu12SuSr2hCHh7pjPl+YM2e6O1957NXV3AliRqTLyLklgeDwf6bJhs
0DDIJK1cCUZZiWeOGlYTrO/WOhi5fDVTkbKn/Sn/VkvE4a4oJn2tPvzm5RFe0rI8
daFrzGcji6B1RqKPsoiLUfyWdZ2T2ZRS5lbdqZyHgAlsVCGJpmIdP8eWgoWPQrs+
EtPTEo/01WIAu4Lcy/WFYwuYpKGIKuqGQYak2fW+50pNEuuNgFqDIZlsn+8VCCI2
J+KTbgI5n9VQFdnrZzBw5MfUsKDcYFkRUerR9nP9JlixHHuqwuCglNImBcDEZOHO
nRj76gLa3hTbnO0vSPTpDjg/ZBuSVLGuO3EPQ7ybW2lKCib/2wm2roRMCLPpD/8W
ldHSB2lXEs3IGnuVoq15oLa+aJfTjMUWxlLDZN8S1mgHII6YAK5h0hKNlzEfjawV
TtH0nFEkBuf0by7L0HKh4/dTPiowS0ug7kQAk8UZoYzxVuCN18SzIilZkBd40DsP
gvqAqPfiR/ooqSN5kXo+COBzI7V3E/YWvW/Wfp8XOdmam0WxMPOksDac0c4Gi4KX
NaNe8NNmY/aeo5hSjY4LyUBdj5GKZI71zhFTrDqZbWuRgJFjdSLpjlVs+mnQZ0Dr
+Mhls0pVZPtCHNJL+QAVo6LXOtbEiYGwnr3avKzantNjF5oyHAUpqimK6eX23SgA
v6LitjL0RzjXBxyCGjtn0e1FE2AGr0PM7haTOJVEo2xMForVtgFaB4WAqVYBXLAx
k9LpFiwvEt7l/m77SL/hxUFy7gedX2cSJva00rzlRaBUadvDyegi2+j1012lZc+4
1mWJDeZLyjv1wOwJtt5o0biP9eTSG/FnsYFinq/JddVy8wTqcVwVsEJQW0dz0J37
8xmsh8TfQ48RUzB6/CIFGQRZk1f/fNfoU/NJkhNMYjgeDjV5uSV7G/GiIdGD3jjd
7WEh8X0w4RqbuoW2pBoUMRGkFzOUZQ6z/b0jGv1OeiSpNs07SBcNZNpglW22YHdW
Q2EzJotk8A3xL0a2u0yDnM87edslg9/+NoJAVlANFbUT8rpcFmbL7coYP8FDoeoP
80UPp6m16NQzYK5Kt0X3AnCJKBSQmq60gQp87RfKrXMATWHEXBFbyd0urS6eJkTh
wEaIWe6w+grntU4rn+R3mzYSTlJ1MsXxlfZNwAwWT6VKN6BHzNmzhIpHnxPGt54V
vTbyPjuBEJxyv3cWUZPhGCeUaPzqCBRTxkJfa0daeyV9lenjVlzvF30Lx6vaJXzC
g4jKv8tddYQ+1DHGxKqHiw2eOXmrNpgHAAoIB5XlHzQGm2esctLaMOSE+FPxkEtM
ijyG/gCHFrbaP9W5bOK6oVJdtEqa3P1yveY03fBv8Dp+0Dqjqs3NmohH2CkZak20
4umEpAnT0KoacKBGjpbK5AuZjB7SL6N2U3Xe/bUXysFKOo1K90b8ikgkCefU74Qo
RIT6kUW0fP6rtXh0n0PXXIfqLg0PNxOz24Q3jVDTOM7AT7egOlCC4ExFvtmR4dqq
viEeMb7m0lyfbzfJXQyWI9PmnxCWYgzxMmYAB2VCa1ylp3RUfZhseK++cJZkiDyu
Bf/65lI5iF7AhyiViRpmRuXKeNt2Rs7ZEZi2+lEhgrQu33DhsIgH/pKSsAqBw+03
TwBsh2Atc+wUhhlcntJRwjxsgWpO/NxM3i9rRhKnTyMXnlbTDDLXc3HGBkeABzBu
DhWXg9NvhXLYRZcnUecTIR8ZcsBUxsg+GvyXr6zNAvhkTYR7XqdJAzaMC68Z2WEj
2dYa3wcZhndQlJxn5RHjAIPMSnr0aYICH54HYVe+I3vShWcPvrHco8eMku1fhnFf
FZb/IFL0obxpNNYkbZJkRyx22EOpXIEnwYjPv3Am3pqbVvlmpPBJRu595MmxtJQS
3aXai4So+WGxVXXW176IQcWgCfz9AMfNxYxj9ifExGY/0pYrRbc+7QoWqwFqw1wC
xIWLi4Unl+rxgtNgvKQEQLqCj8saAnu1BhkpZZxkQSjwctSWyDNACvgosy8+ix64
s7CizyK0hED+wp/gmspEn4xpupvLjJXWmZV8f4R6JlFcRTWhoT1Moqj1546cwcW2
ggdzr/yaFbUkqZOGNnnLaXK5wWFIoG1pyUsLwAm5VZczP5pmgYHjdLKaM9A3zUZN
RuEyk9VYRGXZlRGnBlDhTDJe7IddnwmbS5GIjXAd9RbUszZQPa8lmy1Epq8JoyHv
tLQaBdkfDDZLriA+UqMtj/Lf7dQSkBq4YukIXuYCKWVjk382dz9oosrzN45+72TA
sXHjnUHwX5Kdysy4I5Qtgls0bdjhrW4w1l1EW0JoZ/D2b/roadUgwGb6HT8cL6ZJ
5gUnYhpyZO0zvvRKiwOFLGg/BWeZgulFXsmVxGgCCsXWXa2DY3nR0YX2N6DnSLU2
1/8mgaIJNkpck3fFOfiGscD79vP+IjcpIekDVU/ny9B2lScpyrJY4aFJfTK1gGQ4
/9paXZIzLWLuamXjSN8pD0NCFi8YvwzTVA+WJqRBL/u3Zm/dBhkUmMl9Set5QxwR
ma+tgBXYr8MC0f/r/SOINOSjWnhif9RYsihbjT37eHwXhbFSxLLSRfu26EtaxY2F
v4L1bECcFnc8f5H2ibcY1UWvkaforKSUkzPnfnA23rka4m8BnfGoPCeigO8z/3wQ
6vW+YAbm/DWjGxS4I0W0+KYkSH7fJSK6t7v5WlGs29MpK8Rhn1p2MreZYpo+FiNR
nImizjB02SWwEVcDSY6umX+osZ6SLerMGPf5zCMFtX2rQVsd4zPzWcVgKqOq13We
GGVplpvoivbYufcEUydTRyJc16oGo/nEmdewbMw9aSPWXchx11POtID55CurGKdm
P+vJjrRfiYxXtJc/N1+CtqTtjsRdVIK0Rjnxw7D5oi5kbe/fp/UMEAimLJSV15Cb
7htRTt93/02B2vscMjqA4vZJ37cn5iv0Ysod+ARFoGlR4PWtbfRS+D+kD5rEsrqc
yoVB8Po77Z1lIuNDnRyh5aLax8uZKO+wVtG3bel0ObQOUsyXaOjZXqysF6340U+/
Hojczpux577UVGehXupHxvcp9MHRUciUyx4nGeBCscQWo6zRBf2bv2VDGmhUItjH
Gsvm+fBkUWd6JR5SWmTZwL/GDOMhP8RrY+L65flAYv2h2uj9cgJyrVtvnShC70vk
4hy2pwqSrZhxsaQVELoqUm/fiDLuuRJM2H2AE0Bedde73BNtbJQIgABX3WXQCnfL
Szfpw1iCGov2eew2gctO96YLIL4aZRSUIpUTGiYlJ+k3Z6nO1J8jHsAwD4E1eoZz
1rbDoyvLmN9zHHCGQa4whessMWfEO4Pzv/Hmr2MPYJcK0fw+TWcLUkVxe1WM/wrf
zZqRq33ol1WfsiPsqF7PtJyAkbNqR0c0Uqh6cPG8MxuWil0fqSgHHWWKrv/n22Kr
enw3ZPe5hcVM0eZuLqZbPpc98ry5q0/6BzZWskqi+2iGoHwgVtg9Hv8HUiKqHOte
r1bMYHv/uV3EcpoGSsWKX8EDPWTtFrHGor+R7qR21mhBhOXAoLK80kY8ClmLKNoA
s4oRRrY8ORSYvd7zUquqaKGX9WVygt6A/3PshxccqyizKSLOROLdoB2aKbIQY9+M
/cLYQX8W0cFw59BZF+adBQ5WkhIH4np6HdUMkprJYdZRohuwbVT5jq7gTeuJkTIr
DO3EtuWdw/XhBWFpyCJPsBdEwg8jE6lvf5Zgb77gpHyvSoU5xeMagvqDnOmYBOEJ
lrLpPu5fu3XopuKeadtpiKqBuARyBRyFloq9zlib9619HW11nDFFVi5DvHXBEuVb
47Xam6l3jd23peHOT7HluR1PACtUcbAi/Tob21oq4AO/1e61FXPQLZK7nGtYFWVx
q5Rbnb5w7i29dLyy6z/Ab5buYMVID3WAOjaKX4ENU9y8fcFcfVxnksiL7PFwCc6k
QkZh/hJGVA8LgI+H2wAF7ahyzvNOU88H0RJruGDXsWz9FjZQmq1iWCL100b4lnc9
9l++0woEW9fMOFiYfvqgdOphQJ2RPOnGzM1l0VDEY8rA7iDRs63rJlc0nkfB+G7H
UEnLw/Q/L6AatjJaV74d6npvAUhQoE0W1iwsRdXjp7PaEokLPCdko7geQDgJWSE8
dmYpbp5zSqKsTl4MLW2nV1vkJx98MsEPSPE81yX+wsNsm2IaWPSlaPonP0D2iqWM
fbun9JYHMTu5tGIm4376jgaEXBkCuiPsxaPBQtC3rxcry6xnZDTbqRTGkLZrs/35
KGjTst3e5nrGtGc/LGZ4hZSUk4UpLXZHkoo5ikziQYPdhCHAvU1ffiDgV5c2vbgX
rgb3APR3wuVUOCLv2hjssao23s9olRoWC9S8RB394i41TMgdiXQ7WytIElreK7w8
Wk6oD9dXm3c7jkyF7KgOPmp2M6hJS5hMVPR84wrXRfTdqp/M7MpFbW3w48ER+1vM
yZv892EwMHKstqSN8V16KuSNjKruDDbn3ygkZZUtnCq8iNSIcHftXDe1X8YMW2EN
jfAykymtrpmgxys0z1tNGY3Di1MFy3urogExIIn5w9uogAYR8LBHR3biR2zxkSwu
ALdLxOL2NoomdbX27rrdB8VAc3BWduXPGtIVHDAQrXYymA/SCSZj3gJJxj/L9y/W
FX8dorXf8z2g/Y3Vid3KDdmlnInh0d5WkP53Q8TJDhf1zmRNKt+wgsl3tdoU/W8Q
NHpKgcVOHbUWqWqDnDl0Xx2cxsiqW5PUJuxe/1Tghf+vurZsTaSuROeR2Re2Le42
XwPz/pcNP/2xzCuRB6+nnZXAXfbOlURJFpTOKAAxefqxEpMt5iupa3EPqnvb6Mtn
Hb3BZNRUGOHnsK8YOQVpJRTr+84gLizRK4Y0F4aFMjPCfcXWQmYdKhdk/SxGi9p1
7GpTf05YQ9HeIjDx/ThTjYWGeHnYkg2JClOczHa5jlAb2oVv3hSYo5uwd8xC5BLE
GfzV9q6iavd7DEDBoB9pCy/XgYzx/PAy1MzqsS5cRHUWZEDN+5dIEh93lOmIcuq1
WGEP+fLiDHOk+g3sOr4r3bfH2MI+OJ7vjIwjTfGCkmmJ8/eVVqKcK7p2Nz3Lwmnl
qY+GoyUZ+lw7D55dazMg6jy52UTC/JbmG15cRgrpXhl/xbIXVS73OsQXemo7RLyO
4xMCrcZo6v0pPCVLtv9WL5mWJ9bSJpIzf0Wh7d7+iz2cQNNff2Rni2zeO3ICJ+TN
gbEhP3daDQlfncb6DxkgQ7IEt4FbNa8oJwZdPMXLCYCPrXIPUE60fN+935orKhx8
PYtZGOUst4J/rPJtzH1nBpKC11F7uX2EDaJyL2xWHjKRSM0p4rDa7w6mGpPkwtS+
WSBFXyi2ORZEW7Ry3nAp0srDRx8bK3w10KCGz5MOHpasv3M83WXKG6WbudQjsFmS
xej22OZEhBUfry0p/Bb49yzVRfZoeFWRF7ftD3Z8voCOnubPzZcspgaKLuh7VS+C
XC3/flK4j2E4Ar4XBLvFTje+cxnSYAkVL2NTESpzw5jOBktmQOyl/3y8YKxB9JpI
hgEl+OLzWZe5zxxVLO7BvPEt2AUwh6Kf8c+Dll3U/XFXZmKmcIfHax46aMaOGiEY
nOp3lbUkyTz9p64/A0cKGmTshyP75G3UW8k1Jo7a0aJcW25gpchUSBl+77R2GeWT
+G+LBV/mJI+0rE5bw2HSJI3rmyYpN7i/hNx0QVNQWHqFPfLgGtGf2ESEaKHOgDTI
4mmBRmJxQIex8patcSV2ROyp+0RemLcSlGyOWp+JquqDCCnwWC/YDXW2i6xqIIcE
DaKd2sJxIYB+QQCD2j2+wAqA50NoRaWbmXueJ/bJ7Xo6z98GIDrySWU7ww3badpo
jSNOo2tjbvsi/Dzm/vAVve3FSJjPHVtx4lXBkIcYCC7EAARV8skBEsHu7bz6cEST
dGI9mMfyDnQdxB0j1WuXvlF8CiiCtX5lEgtUwONLlMCnt3StbeEY0di1JjgzrnOh
2lZ6wImExyFxu0GDRV4r6tHpyr26EDMNVG2BScTaUn0fkLl53wkjN5+04Vc+9FuV
PeCjmcqE6d7JcvMNa23CzbL73NsdCvI3ikBj3dGJi+kWFLY7cjx4dk0rM1ZMobq+
MXgk6X8KQ6GAGTZfJgHkUnsWFsOqAptXk693gyBJiFFBbx3ROGUQdXWwM5BfsPXe
0DHO5Hq0ZbcosWkBQu0w+jUFf2aw+UlFzSo7guXCzxdOdqb1MfPkETrLO7/sl7+h
ngY92CNVd7Bci/u40cXd6/e+KsQgJJ5fch54+zX5HGZKO8LMPAqVthgNvVOpx998
cBsZqy6ymQg7ulkLaUS3wG/tRjkMZ+TJ+EMxrvQOYhiEN0Krm65JvWZWiM2OD2Qq
W6ypNyiDBdga16lg2HgQrL0DeveXeC9dYDgfV6j65eGTiVeqqq0FGqgA7xedc18C
WBhAPJYG7cTMVHZnRKkbRkwGlJL5f9rkk88uFZB3rMf0Z+C3TQtQLJwKa6RXYSng
PXVolppgAkR6ywfjoTuh6OVvAz2h3zXxrGg95vnrUVxUIbyTa/m4JXiNeTDxx70y
kjZA8oPXcZqgzT5ulLHYfKqtwQfYVj/03ZNPCq7TKlKipL4ea5qGhaEKbS8GIvP4
QduE8RUIzXlEu7ckMHT3RK3dDe0hqYjoGVsDQXo1U2n1twTonHQjWYTa5q7y1foU
dNwZJMn4Ktg9zz+IkuaTpFnXLEEiSXJeWvV42XVO7v5UXjz0NzHPrlwrcGhfoVF6
JzSSJ2untHaTF7L18FOJAKWEHeB0NJEp9LOm6xzBVsB0VjzBE/gowxkLjGbcQhDX
3Fy4NzFp7ojeYu78rZWgk4gyxQFh6qZXFuDdfyljOQyu1lYIq8QxwSwGvz7vsZpz
kB6CnE4biydVBwqh5nlDnghNTqF4tdLDoLZSQthC5/HfL54m/W0IODfZQDNGhF94
bCLbvHY8n0lTQXfzoyMX6xkR+6jjJLVVHkLhqCFvOfx15IJyCqJVE+VqH/fsuBlB
WKKT9XIkxl8ylluKVRv3p+OjOaLD2XetWwNqQLR7CTyULY3QqcFGC3LKdfi6QoyO
svoENCsnbGj6JZIjRmKuBOUiUXGh7DEgFxLX/qJdudwJUXr6hrAV9od2u5C0prmx
bt8Iygkl8lZebgIROwEdwYzv1asXjTgUpkoOSUaVOu1n60YpmooeNRySayKz0jgq
lusfO9kcRsM6pDz5Vqaogh8c2LveCfphtYADAVIBsxs0kZ8HplfJuyZSCnIQjt2o
U/IILel2RtOi1yoNKOrAGvXmBF5ovPwgFMo5Vdc8lPiCL6vpNslJFAlV/4YK/VA8
ckuJmKmvNDqTo4H6Gvk4gPW0MA9r8GubXDbbeaJnaftjpWUH5M2H788gjsel6DUd
v4zedhkcbOOBiEoW/ZbhX3ezmiMxJD6YlL1He8bf6ltdJfUQmMpLfIp3lTMIrwNc
cMWjpINMWNxVIIE9wH4wMhqYRofTlGdUrKHDQS09WCVead7a62XnEgZ4wNkLNRqq
/uJX+CqJjiv0S3nHCZBPZ9SsiDiFbcSCkddiStw6MwF1ZFCjdYlQNlIjWsfnPPkT
I+RqxpmqMV03Dt79XPxliU65bCJNui542V+WF+kb/PbRkdJ3sm3i/93sAwOkizIX
GuJw41bKlHQRMMPaTZCvtWXWiSmLxCe5W3/w8DLT3aVGgPt8bN1hdQsjgturNEoY
ioXuYgdrWIvUMjVTAwMY3zHSkO9TlvQbeLn5ZD/tPf7zpcgmCPaFmQUe6X6KlPu0
1hB6P3rxd/427agrVxGMYoVPGTCmjjZ8DiXMpEjdq5dQsE55Kpwjdpqv9HcgPS/Y
lX3xTunbeBvYovFZxiam9vcUd7FDxn03A5LHuW+yyCvOqTIMXVY+iDNdTuwhHTf7
WxAb/cK7Y2hg0IsAxhQMZeNwQrhejDNrymkhWv4/iO+iakRgOnDIuDcbQSRdf6YF
/trFf62F8q+oqH4Q7xMwsy0NVuus5Y5yvo9xj07jKIWlAEOnNafmxEsvluDIvdl9
4o7H+gx/UI4+3GpMDVIkS2+2mkFmsRlSoILDfXGMXpVah08DMitW1QKykQQj9ueE
A9/g3mpbGVhrR3f0+cTA9wuKUJAbQHVJoQnbco78cbJ6ZGhET5u2YDCZcYkyuv0l
uQCe+459kNGNowb/4KNvu8GGZtH1AsKcJ++6DxcDuBLbnD6x5z1ghjKfozDJySeq
OJ/XgforXBpg5qYRrdwth0l5+PgbJ4mo4u1pReEp1A6ZG6l5bg4Vh15L2CvEfL5i
45b2klGkfBI+eWodi6bOEQ0J29W6lyyns7HKQWoLazleYwTL7ucVPYfpq34ATPSU
IqMg/RiiH3MvMDPXPMZU/OXovA7vAVf/5npjVtLGdjPFFnvld+BaWg+PQOZMxeHU
cTd5BFNIUszguzAKAGUZG6XCiWaJbKY9JRIgTezKkSiuKx2MRH3YdQvRjsxS0pGX
XHPy0TfZcXmPO+Oo99lEFaE5gBYxsuDWO0nTIqrhOdf128SXvuz25aq0JaVjQei8
1Gq6dczf5IzKK2exiR98FsLZJ7Uu+3OLTBw5Hz4rWRiwCElsmyUX/pwndXVhbEJA
YIN4U+gm/6EFz7yf82Rrde/HQkx52q39Z4r+XpPiko+ZTZr18w28AT2DAZajSfSV
71G2VO2huQ5tjMlr+f40NuJloKQieVXnz8TgHMtbkRI6XVkqUsptn6hG6dOfL+fK
ymMsFqyAQt+cyRcd8ModpslFHMkXfCXU28HLQugMjPgjKudWABSKy/5PlZSqCDt1
9pAYKrtOgVB83INnBXbvemtIbjPrkZ+4/7sFYAoj2b3Fir4iSUHtXbcgHrm9/uQE
kixHiP3zfQ8JgHgwp7Ia1zkjX50N1rMT2OR0n0mVQHiIR98Mk9UDxHCCi2tupJjb
M3OuU4bgurD2FReRtv7gFH/HGBaXuSwwLwbH3wL9kxpNFRojvTfo77+3/uQdjwAO
hsjjkTDDIYxQkHZgrZ5m/nhEmOMZIoXpPNXkMG0xSHjmLBXNXbgOwuEWLSXCCBXI
nhDYxJlgw4k6UHlbiqhvU+lIXSmKRenYFTRAFfusCKlh83uaxaETQ9DZTHJBGO3s
W9oc/azH4eOs4XGTiBjb1pV5ZSLrTkY6v5Kg6vhWUyRI+AK996C2Nxp+drcWud2t
6EL6BdQd7/+mJlKVsWZ5Hoy2zZ7swYXVSQbwjs+iNZO2h0ZGHwvR88Z2tYpTEYW2
lnVDdHW4Ffp46tdVvUgx+CWcWUO6eqFHQsvU/2hvx2rl88Jko+fHQjN0KCvo0Emy
ZHMPavzHuEb0NWQ0THqsE1TV15BbWFhr8w8xzbcBg26op3T3SduZ0tcQuhiWfpt/
kPZTfvQrJoGXiPi2mo9N/B0Q0Wl4e7J7KvuZ4E2/7UK0k4eDYnX8I2LNBhSpmAqU
EyO538oNEnIb/HnmTYVaEH4s9+IobeisPlnopV6KiWZ8WXXzdmF+C9HWYhJCIjZP
vuzyJ65nwaoIyoPbBZXak2EbGXOrqHqfhxaW6Rs32tIK/unBmihrKz+whwm6P3LW
cIn3EPz+Ryy9ts6TDasrxUx0AFPmSlDYMzrPRoBnspwuwXQPHAXKkZqM1GuZ530P
u05LmjDAs+G4cb2X0Z+J2WtFYsLCmVI7hdTNvpZo8i4A0ySb3plK/4rdcbU8FzVf
dODiwUpBSYLYzsDpb8t2vhsaukvPDCwaUWdARHONwiADHvHWxhzevVnAnNjTd3Fz
D1E7FgHZ246V/Rfo/UMmKg3bBkjinOETVeBpIq0Nu/9MMwMVJZYleNz+lnKcoUfe
BSXsw0beTYPwWSmcxh/9Af2jtF/Mj0gnLiR8dfvS3cpMjpOmGS+wfsCU1LCGoSdh
WScgmEV0fO9kMv1T8/HKzzESiwvm4ghPPpjgac/CSAm7U4Jf8ABxIsC+m1T8+wk1
OPgCzhb5tq+7iAvrVeHGZVXI93JjtXWFi7PDEN4m085pyMcZ39D3NzQVStNCyJtn
rB3xO2FJbpS+Ln3mteihPFcEBsm9BSBZaoSDf3eJ5sM0B/AiSuoBcwfb5l6vbfTj
/jVPV5XPhviZZYhlevPywer3e0nRNscG+fNQ34ZX+ItN3xOzc5f1dQLz2pCrxR60
4wXkk58wsoqnPAD0rQSZQKgqMXHrGr565s+Gf1Q7W9E6CP8XuX9GvSaXdPtffCFA
PFXCLjkd5t/B0uSS2L3oaXCFBxISCQWfDhftO/GK4KwxByn4RSpj/NaH16kuxquu
dnUvFe4vAtPa5bKSCLblAb9qgJT6E7L4pMouGWtuIvfhpfK6Cmz/9zC6+1lsPjqt
fFhluc9p3Uk5J8ee7AVoTl6jC87Ftnmy01jnk+Lz3rqcP27YL9jZNHzo6tQCquhZ
Q8MA58dc/z8BYwbxNWgs5DB55tjco+sb8bwL/DezT2Gyo8ElJsbR2zqZK1KA2z1R
yVkqz3fMcFW8lUh6nqeu8HeOyAFeemL++c98yv4f2a8xKuqeZT6q+5ZBqQXHocGQ
H0KrCMLFO/3PFBC9BT8iUbqV7tiXHCyxD3NOeNoN3bOkmSjY7jlvhZjb6ERlF+F5
rz3pOHW2pC57PhNPBn4ris4P/eNxxBsBpjGO1htaVbA9ooQ8XsIrPtIrMAXTixVm
iNS4jK5hM7AB5/RBhuTJ2ZVfStOTcn9aEs5ZHe04Bf3XayhZBh4s32AN/rNyBmfo
YiscVBsM69lGWLDAPeY8fWoXPIh7ZN4XG0r90HJNoqCprw0DRH2/PycZoQT97Mld
nDH9QXXZqcCQqP/G8FY4Eo7wMsdKjie36a3oeJ0uVmAiQyUAFfggdfriWKkv7A7L
SHFBB15D0TqjT8dgOq3MxAHcE4SctcUMigBG51ySJ/BrDd7gdYw342X9S9tVgson
1yISZyCyntI4XRBF8AYqEupVMR1poegnrxWqzWpEdyotuwAuCaeSmbLB9hw298ej
4NEv4HmmRUIZQa2YKVW33FR8NfOb7Z+s8QozczyGSyIBMmg5MU4/lQaCp8qWKZKn
oSUA+UmN8am38n2H1KRNiPTrsc97+RDXUha41ZKf+/O0YHWokzVKeY+9oFQedPv9
PjTm8CB4niOOtIzo8dQLCE+AsYqu5vdmmyA7/+H75uI2zVytWKY1lmcLH0Ji+5Gp
kgdT2FlCmnLlP4xwUsZtrNF8xfb2ItvKTrmn/PKTwh4LxpIcIk6GL75HgfT2wIo/
wRJ6KVgX0uxgXg6yL3mZK75wXaAqITHiR5/1l4V4ic8ACV1votY88dk/9bphBIaC
z2hadv1FU7sNHTIyYPXReCLpunGC2fxyvisQZR05Ab6pl8NZSGca+VEaWrdvRmhp
WCW7I6RZ9328hwjMFdgnpuaELSOO2GAtEX8ww+WVrY1NpuNzxliyL1ejeAUReY7J
b6A31r2/cXu2t7S04hxV57L3N9ChZe/vfXD7KsNAZcr6Fn6SGb0WpcDD1l6ME5vZ
xh0eAkDkIoq2/JAhPU0DqNOgdzSAk+QpH1tF7Ll1LtBGlQ0vqTeNLuu9SUVgBB4o
813heZXpd0boAqlowjHSr90YijJNIMXB0+kucKBiU7McA/cajXab96PDHDpjSJf5
f3Xj9+WFiI0BXWuwI1yjygFWMjGMaGqJVY1H5R/2dYMPl1lqQvYE9q217uAoT9DD
B6kiujQcc0vA/YBwuRiioj6ogfDrIvZsYOkAxOfu69iq6ZYFqAyUVQCpzP0rOyP7
TNWR9xNsOoTYz3Jm82ONBgpeht7O+w/7dEmnu8ixs+YBYGI+I9jzGCEUbLznHmeV
mzQPUN9iU+ku1klNoZeUZEK+LXLx2G919trEaa8oi41W9VbRSdk/ibDYS/icFhvF
INKeMjDxVpJ2xqQKgD0qVDG05KhsJzgsPsZULDixCiM90uUImzoy/eglMgHCfRh5
7tqtjB4dYcK9nJn5nYnr6sUOT1U0of+M93sl1Itw/zT24YLsDnpC8eZmPbxD7hhS
nt1hYT2HGmYKUdthOpQqzK0Io2Aur4xrfMkxKrErt4ocBvv+7zYkfL0c4K5TNuiR
DJjkpNtpSjYBEMQdCTcgteGzQ1EamYlswjEpXExB/KzHPXqvE5bpgSDz2J81+Ana
h+gB/M6qjRk2J9fDmJvqxRats3yzbbpgk44dVx5uIOivZ1NCcNgmlndHb4rHZ3YK
zg4KLv5rU1TXLepyGSfMe1rRyKJzvcLxrI9eLt7uDiypv+I2RPK0LdgYyygtkQhF
1ndxirFKig18QmU6RsO5LjKK+nalDHHR/QQZNDxWolOqVxWCWwAiw9JfpXjBD+pq
t+SEHYCuS3MPUopFhsAKk6SnW9pIZXEGf5fLUlYHXgVA5U2vZPJLgwlvjLVt8LxI
OIk6/PkGk/WxGLxWpSFljGn2RPqNJPnjv7l646jdc68fOnYZl8gyfkpljt7APOga
sWzybxG7oA8Cl1JQhCVPiy9xONozftbOi3JsMtAYqr3zHHKvFxJGuAf0QRtspqpO
dJdcrBFC5xEG1l/KiqUBHfCuj2fDNqqhySJMaVwoyciHMFBqU6IKHMqZuMAfg+LO
wLv0DMbZ4Y/6Ae70l2TsRbfYbOiEi62kFiITLBcYr7w/ycAtXJTfWIx1aC+mPYGN
uySnFrjC/mpt4fduyiRVb6Xq6zw+WWd+1JOmU3a2a8F7gPS2PicWMaIvbcMv7pm4
B7BB8JFV+hoD/5Eq9RqhdECAQ5d2OiMjk9U9wq2sEyNA34O9ysOSGNBOyp+ssp6S
oV4XNrpGQti2OmB3WgK2HZVhp4iU1oknrf6SjL57tCMLSeqhRh5zCzPfhfwxKCaF
h8GUVSSnz3JKTcnIFNYDKVRu3fnwXQsoPOQ6u/7dUGI7n8X3DxTVa7rqTg+LHV9K
0QiMmzMqpTlmUpZ9EMqm+TKOvj6214gmKDUkJaIzXC/g19nVpa44Nx64E79MhK06
fkBmP6hQv+50LJ9RF2u7oXmXptQcVtTrZaCoFheASOkxIba4x3FVTpYh5PUDA0Rh
QltIhYhVFxui1soe19AAPMJ4va4RNmtLEND/j+kFtMM6/DUTCTpv4hj0OEvsBv78
GtnQ1op6hOVvzFWW/uxy0Q9RkHsJr2U2fwwXqeB8K0M/KeS6a6HSjI20gdFXNtR6
MiiksW+YWF4+i651yfYTw00yoVOp8KHRlC1ENTWA54gJfWQEvadL+H38rTcoUcA5
EQg1N9tHf1hppTumzCdCNnFg8PJsXAZ5sgyV+4kUZFnVEcNxe+CtR5N9mN1o/avd
GBna9Tlf1A7PQEk0TkT/H9PxHr1yl7tZslDzbHjYTqetX17HuJdZnF0GjnzCOUxg
69YHjHKi4GsbSCFChBarDgR2lSCYVdAa1lc/DHGkkw1hGPdHswNlZKC4wEhfczFw
3jCvDKbeUMV81UGQWrvEmHd4sHXaxYpBOGK382PkmPXyBGK/8FL1RDr1e7V9Yjju
UiJUUpfTLLp2BSnZuX/6dYFxC18J6TQOi/cLGt2dfH1ahqlEf5AZgPEpcIdn3cPm
s/QLMVFMmmE6/IQRSQTQtzg1p9vReNFWBXFwMS4ESYIqSVcQBQjn4vdae6rbmC+P
kc3x4e+JRRBAuR538zJQgJHI9w7EU5+BDrblJOheeWG9o1eumzjcSEjPaczVVzrY
Y9y95Sfs7iZ1ZLXZF0x8+7MU3CrfqPVgtEHA+mh3N8H99YO8WI0lso/2CH8XVXkQ
ztT53vY3WBEh/DtA7OTE7r1v1au8n9VozJknhkRDU58EA7iEDZPPkESoiDD9Cisq
2rC1tbpOi7FWFqIXvT2gZxcxyGNbXHBtK5Jici3DS/S+Y3cZGX/sPGHIIMApqEC0
LmkPSRc69Svc08s+A3aN5V4DTLEwp2m5++luShqFcYoyBBWH1D+vpP0TML6p4yPq
QUmGlLXh7ssE2ma+Sf8+tV+5Xcd1p2LCQXf9hEfYd38auOmZbPbnhj5UjpxAb+DP
NNcjIXJeeVyIelHDWRD4yaOVTcNOuRpY1lKn9Xh4C0zBtbNH9qYxJj4XFZAp8ni4
rueZqygBJAYjrvFYQjUJjpYm0/62V70NfnlWsoB3d4J372FfuYfeme3JUqzoIQed
sRXjBqXuODMaKXWWYUq06CYR0LOj5zQZQFKw73YQad9ohYmi5D4zIvHDoA3cdlLj
Ro8LLkWzqBiRUsQInRBP7aYeEpuA1N0v3vJHQz+Rw34VD6qXGVyR+n9ctEs0EJG9
7bFrElxYHLap1oECg7aUtz3WNa0KxUA2jpgToKGhS37G9SjgN1M8Q6hvJybIWhtL
w8g/WxbzkioJ3ooTYgct8yNf9s65HAeI78JjvB/0Q0id6KHA8WGIHvP9RosTrX+4
9xDxKimrez10ck6qaj0u9TwoBQCRaVHIE1GB1oAG5dclqjRGdkxqnBFAsJdhkGMP
259BtMSBKTDblw/gWLutigTZLPv6CUm/Z3/g7OqyjUcWB3Ch9bZsqPkHXR2/PESS
uq84sIKiFreVX2VX3RiS2Lw/YIlMJx5LfqcXte0huhtx9rwIvO2n7qCnEOOp/LgZ
fx90zkoHN7J2ihrz4pUJhABUHPmfvFG+i7lswofN+2xIFOgTD261EjVGU7K5mdAH
ih1jrRn5KByUKQFCf7DqKOH+sPhbOpWxoGtwfyIDfQNz7xjPuIwv0UvSfYb8GbqA
l0sNktYTb8hM9s/AADcrBw5O3MMp5zqSalvG7N+GmcgNOxF3DfwdjBMwrjku8N8T
q+iPCd8rnkwgxVX1w89gKOL6dx6pIzmd95gcK7oxMlZK+0mWP5YA5kja2dICm5n9
EWa1BQWuCWhVNr8utyikNsZtpl37+AZDjGwU+wQnQHlbAhB9x5fakqtLaTeWc5eT
41tl7N5AOGgIk3ATRKWjrLqLeCnvAYhUztGfepS/UuqdS3GcwdZsb6QHOqqfwTJE
GMInQX6dMTuAJVnfJWyWAlTOi3nZ9eg6T2R0Neo6sGWVnBULtv9k0b5VXapRSZq5
fIsM5mvo1+PRUIc1CaCcw7kzHhXMkganbYsQaVZQsPaxJbcWTyMPxdg28WbCGWci
+DyFx1a7H8e4pAHz58azH5gVL0xjNTISotetIBXSve6/THXK1/5ZXqz2y6+njJBh
kmyGnbnL8uA8F1EJuO+PZ1dkj9dK52ZYa6TYmPFhPZ6ptWSMR1QSNeLzmF2e4+Q4
90l4bzNgqYipfi4MgEMzpYbYmjzWLiNZ04qI4J97nfLvXtFx9Z6VN0jQxlXtaFNG
nIlVI5SBJd8IX1tJJ+iXKKxFDqnaDucMdF3C7lNMgJzVbq++jRXDWJrxebSATH6q
2XkRcK09DEiyuASBQdgcP2wJzRiMzubO6Y57+G2478TgSoSsaSYR0T0WWJ2fcNwT
toWijXR+yFdgwWKzqzX+Cw1F2x9l28KKnrhqakZ7AlrzhrfCIPfCPGFHY8tSLuSM
4kONutxBZcXbH9Arx8fGr8VixSomgrFfkKTj+X1Is/gSe7CFrPR1oCwguUjngfn5
dimugEGnVySvpgfqD+Cbx1ZiDweYv0+Jb5uly7JKjObNYPqCTWLCZkj4eHfj7Dj6
WJrISfBEl2oJ1fu9lWxyl5/tOOCG2A7dTM+D+la3/roqZeQ9BWzwOv65gPARdTpL
VyUYKaepobl6rwrVbUK/xHBe/rj0HBlOPitAo/dPGmAiS71xA093uvOeoGESki8f
VrdRgirwPHDXmFKe+vD6kAuGkHCxNYXhu+R0oAMrue+cPkPqGrAkY1spjkvu5RYJ
fJ8dG9WL2EX4+qUX8pHSCLSXkkFOs8GFwgHLoqcT0TwzzUugMZkTUpgmfgtBtWsS
9i3fudhc/KnKWU87cFck178uGgrR5zgRhPq9j+UWSbiwVY4Ut7TSZuFN/KdrSMZI
yEgetG0g5lvKHtQT8JHjuavMxHuxdo+b/AZuyvTdKEfz9S1bra5mfTfpbCGdNkvv
2hUfQ4jZZIvSSc2z0T0URteR6cCchcotFqbcqnheNX3bUz3kUiTImIrJTUnvzky3
lb89E7kHbothptKWAEoZs7ec/3KqSk9ft+VJ2kR6Y4fyMekRc6kJkWRLZoh503tt
m/HlLzBqjYb/wK0wvyZHHWYSFBW25VVNPQn77bFCR0OC2DYCwz5RwhYVD+iHzn4J
j+CnDUhUYWiE9/vdZdWNdeQq6ZoVYRFp15Cmy3NhJve9+AT04kUfnCoY6YvOMTbc
APR+4gfPfFbSXfuQGKBdhYWNls5Ve7w2kWr3xtrjJ0NfQoS0Ibt0K+K+QUjIs+tc
/yMDAFbQ1JPzG858acOJz3kWntS+GP9N82p5N1Qj/fAV8Gs41jAliL7WE+KWBlOU
rxamdFKdSe9hiIcpq9Npr6V4Kl4JDr6kUvCMOyEo6pL+LpI42SZLAKr0L2eqiw3M
pylK0BXhARRJVMeYV7rIqKIGZcN3RnW2YALQJerPjenLV4pUf0pPkg/DFowlgqWd
q+h65bZvtCLN4hbPtzV0XpAQMytAnkHl3bCuRsTtC8Oz0LTT7xUpC7NaDQToAMYq
q7ltcKPGRRe7KBukO9yQYWMk+G3utQxLbO13Fku+b5fdJwFk0o6RLs8cbBFecPm8
PUKLygmBBOvMjNqp7o5IXdDYXfro97FeC5iKgblcE70MdGMVUq8gmxKYWqzlH+Rg
DUXzcsIC6AcAaNj47PeBX29WEr96gbKbtj9b4L39mTw56CW58gN/15Zjs60viquB
h/MoCQLL2vBER8t3yQYMUmOqpnvkFY6eE4bh2ZRX4TeNnAkabFJaKnYzqNpVgKYI
IoG4j/Mk81L3SXmTOlQ03OqmzKLJ50Ir+i7nkT1HgeWBG1JgzoVjWF4U+x/7q5+u
S9T2I0SEeO/dIllkTxBiGC8CKqpVrPrP9PUkhgcHQmn9Y4RowlCEWJTF04aAKEWq
FWiTTMjSoSjePO4AIZjM6bdr2AUqaiy3aHZdsH78ttZnYalBQqBS0eRovYXn/u++
LVkMaq657So9Pc4QPeSOaTIE3zcj4nQW2rmgdOUmwHWbRgvpNylhaJRUib5PSNxx
oCPtAKYOECcHo6T6BqpQdtEf8ICODTvITk4KymSnRErflaqcetqMahhyTWKvEUwM
OrEn/EdBSECEfHxqHDigokjFrukdp22yFEr3vxeDpTnOexbmN3WOBCfvbrWMkdD7
t78DHopPlszJbKVX5OS7vsN8U8KSC78EvEoHF1+6V40w8KMpdtIj6aZJkKLj+W69
4yYD2dzY2EJ/Z/g+AMe/KxQYbCEe6MNSmtzpFLUMtiCcRAyIfOgWIxl24mal92Af
xj4o/+Ooc8acOb6lq9y0JOVWHO1+lqwkcLikTPKo3q6AQkf+mACd4JNEWTbeUFR9
QQsB6s6tteWWTeWbFK8qxuJCE18b0R6L7TUgt7aVKM2dwZvuYHK+ZgpotQzdMJr9
A7IZdC+uY/YIQC/AXN7R4XDM81gQlBOZ7u4FePJTt4CR8RBJp9kmh8BzvvzTHNPS
7cl8OJiw/niFiQ58w6gPDo7SC3GnQP1PEymVp+WAyzKZ68dXn8BGIdHJ5VRboPPo
S+pAGL+9xaIrDlAyVTAXJNj4ryO6lUYr7tvmDykKVAJS6QEKJTqrsVnVFVCpeo1t
BpoP0T6XsvRp8g0zwKDuZNtJI0A3N1vILLQmBw9x6RoGZNthUTsS8SBRHOlOuYqY
jd+vnqCYQX/2oEjeVHipvsgw/8cdraJiqBh+AqeV1PwtU3XxXFdBlru1da0JqR15
D7e9+JUl6ZEcdlRdovI4yMkekyoW8pOMFj8ooDZdbgsxt72J2iOR3hKFU6YNcBmc
5rjwHDpnvihvtASgl6lMW4piQSrvKdR7kQR0DmYpyEOwx20QIi1PbpiYA7qu5OQp
H22blZAWFLeWJ8l4NEMLo5rs4ev6c/S1nGv3tU1eBvv6vSHmHhvVJYwp4ic7sbac
3Mj27Wl3yTEqj8QqNp/2BaoQO/kS6WUluEIu+T6OoMQiu4j+SP8ruPk4XvPspOku
iK4PIjG5rZ4Bmj0Dy8ejQYI8Lh7mxXD0VREbKbhdOqrJUn//0fFvWZaR7gODN1E/
5i4PvIRFCLKTkAlJ3Es6AycTHKrvCV5M59xrrvAXlafLMr4/19tgomPlKTz6pEsK
Gptxup3wJ1+e3AIy37RLNHibEsFo7AZw1qbLAjWvyo2i2QB9R0fTe1xWgqmrELKM
0MeBAXu5s1lRzYzpPC5RKU8UBQl4jmCIg1bkknNuj5/DR72QycK3v5DzdrWMXSRE
AULE2B5eyN1WMc5svaH1X1z8fRnY6upzurbl7uJA2UH1F81ESfi2easTqXOvIwM6
gMKsl0oSTvqaUXfwNPaE/QsC232GEWrRaEFm3Jlp/JjZkXlKaCAblN5BxrPzMN2M
PM58NyJ5J9DzjSuUzCCmAjutvQxhMxW9hRCRRSofWivmXoDIZqIDeuAiiptk6oyj
SsGdtGe6i47fw4BtGi3pIFpRoYRqeA0txpxgoYx5CT6wuX6kJd8oPrDceSEiK1yF
dVNlvxmQK402nhalbNZtW9UNhyLPd10w5QSU/oPLyyaxytHSHmKYjdDQO2rcMLRO
3qX5Ir9Sg2rjClPO+jLYpP/2LfeHNY/EMQ5Oq13z9vx9Fayet7BDh1v37WJXn9zd
XZuiHlI/+FpxyF50R+yB/6i0XLj4Hv9K9zPVWG0cs71V8PXKbGR+IKkvXGSogd5q
PHn+AnAPFHkoJH83pNQagWbB+MnVfRXsCSbTjIvAkC1UzlcjIzOtk8xSkFcYdAF/
uanp2H7kYhoHKhMTiwc+7XZyS5LIkbiCprZRUglSIylT0W6oWbOitCfklFSehK0t
NLNpExlFRzo4keUWybhaJAUKFO/RzH5xH2Ig5NwS7GIeYFn/7DdDhEeWMRQGrDQs
qD0Mwm5A+vTb3zJUd/MCaG/GU3pR7V2YOH98JpGNpTNT0EVWU1kfHb1ZWUQAQlee
0CGSoh7RS76u5NdCXQQ8TqACRTtugq+67aCLF19whlIqm42Tj27ikP5SOwFfVdqw
DdFPPqDxjH1c8RLWqMf5ERKsdodhPNjxc2KSQGwAitrT8vSfOj3Q0/HmaNI2y/xA
z0x7HdWgBMTEBEihR2vmivDae39WhfGdYf9xRWas+FI6IMfX9sCX4Ffys0P+v6jd
Ts90h1fdiUvm22KIAONLYFjEfp01DZ5xQsp5ycW5h7WAKlz2gz+eYsD8SfqsAuJi
DoSZpQKd2qpS4jxIURdYmJgcU3j76NHYBCj5XhBoCNAetTA1hic06RB2YmnucF3P
SEte5SI83NMLqkCUbukNRxVisi9P0S5h+eaOYWv7+FNCbGpc9EoldcSrmoL5rSWV
fA73zc8GlXfBjJgpKL4uNp/CuhcK1CrzKmH2raUZdoQnhUsGkdelyage/ReaIbfK
wwqJsoWoSeFOPHn3ddJsE6W7iCc8Li+J1rmezVtItmEuspRqHi6HGDSFu8ohUij7
6Y5XkvGHSSb9AEfm35in4pHKUKIFmmEvDPmZekSoYTqqcs6DyFEjEGDm7kywtwVe
v1RodexXxpP1QdK1ETXP36xq2arVERXdRk3I0qhX87kzfA1vtoih0FWfr/w3AzXc
B+hMUntM99hMjHPv4pZFsal4h0h4L811XnbjZCf3lKMjuVHRRYfscbnv5U2XUudz
yzZ55wL56iZV/dpn0ZUW2ST9xFbvEOk5wgFaIRMMSeigdCQdW+4uXqA4xoLahUt6
/j6SGXRzfzg0MqclZArUwoK4IpQXpzrC+En4Xw49R9O0vjPf9JUO9siHGAijxR9m
T8ZUao8MxWmZqhATluRa12weXOPKwJKdk5PgpNVHdIU2NP/r1AGrFKQsG4JL3Gzh
x8XYEmohqLji5KtPs4Ew8vwtuF8XeSBOwjIagg/6gEXQm0EbbpvuLtkWi8kqW4zv
5cxbNtyO8mBKtDovDJUJJdBasDkXszPce5yckYygZnALWavaY53jafz9hMvXomo4
ws9cnJnxqH0vrOe3t6pJ3s0Lzuyk+E+DPM9KGldKzHqhbJoWlAWjiWldQ0EdPHHB
E2xmdLbz7bHKBxK4iDR68FbHu4LqA9c/UKW3N4IwHGDpArAjuK+W0YoOHH9DATkb
/jv9NILt2gPCQFy6KN2Lpf7oCTS9s0R05xMVRAuenlSN0hox68gs4fYoOe1bmMJi
LX4HJ/CrDH+TIokhCkBQe+NeW8cO/nszDTVSLaHblBRwHM9YZoT+AcFC9deC8M/P
BYmfJYEtS9odn/uZk/SNiVayYC8Y0VecgDWmkkZIxCf0Q3et6C7yXjLiIZzX86xM
/vAFmV0A1RJ6OLsI+EGYMWiKuXcismjBLO9HdjnpZizEEb30rfy0hR6jndBFZfQC
zwC9mQNzDRZJzCy3uzVmOg9AC7pUkGkaZhXu6bSFxxCsivMBd0GDWfKCBE92vpc5
O+ft/2YgyxGirlEt4SAIbMRS5mTZ1zSbJpm7blRD8PNPkFAxPG9dPMhtybcoZ8Q1
oTGOFILFt+kYVdZCvFpKpubZ8+CRuD4t0/Ruckife5C12CmFbGdMos+CWGcoZQ2c
QGwJMxsKi9VMjaQVX3ZyVVt+T3ZIxAaZ9MHFe7NVdAyomXaw4vldBVCSVa3ovDSX
oHtV+olOIu8DF6IT4K19U7reVLQjtM9aGk4vQkAle5gcnL3RIuiXTKkJaDgKIedd
601FgJM4TOUOQFDLyBy+3n+T2eDdQOZrMeRI+JO7Vio8N7/nBYPpLAfcJcrj0gZm
qqk7o5JJ4tavPIyZQCFQ0k/jZzkxf4on3E2CfoBMb8vBG75ZMHeer+Oa8trPQvc2
qGArpYnA/gCUlAJTbzMPQlPSDVrm5hUZoFl9gIe3kENLOdGu+JwGdoELkJv2Kb1J
1sqHN18YfvTRDLoq7DB/E742GgoMpffRmDR+GqAMHKpFJWwrU3JjrOqZZwoqaoGk
XZUPJolJN4yPm3Bshh3hfl76Fm7ou3wS28AIxqfJuFpSc+sgR05n7z0k7+Dl2uQI
R0ohihgAEVY54DtEiuq+RMfcFUgTxMTmfj4aeNOqlsS8XtifYW6WXSxdq6e8DSWJ
TPO4WGBliD9muLy2S4zZ7/aLNIyShHo6mLz5xPSwGA04iiU7FKnkfvnwGGeBUvno
hJpBazRVdGWh8LQHLjdhHDpZ1ynVNZFvdN7W6zBww+MN1ZkEeIsl1eR+dWmXMCGN
9GJGRZt94Ad9kf+y7uCA44aPqUoJFqFwOTW3QhMCUBb1ssyVxyWqqweqVV2IzjbW
6iz6vj5V7fwZmqhA3PTptO3nrVOtZ1NxaJ+7nyH8/aBToUfJH+oNxA0nwxG7VCSb
iVFgroxgDi2Xs0+xSepGcYxAOjCVtF9sqOIrTEM1HsPGyFxGJ4zXZF+/V7LehPDq
pufX6tWUXsdTq2Fach5Ozcnn9DJSnW+QJNFePmMJMz0SvGmboxWJnTa0wtLwhv61
G2kRcBxkhDFl0JzYsUl0to6TxxkHaklj+OC44q+InQfAOm906J3TF5VUfnEN3GUh
eao8z1t2RqrZJOaGep3mQ5EI6rt2kQy7CFy12ZQ8wr4nMbw1tQRuy43AQa2y518R
oe/+xbLDIH0+VdYKvRq4bhwOB0IR5pT6sPg6J9wApPfVpI96AkCrdAYZL8EcYaum
s4LdkyGsjWbVjPtTN7y1HqlD0YKbX/Q407dhwd7r9OiAczlo0R939VagN6JrLQiR
cvWQ5Ih7xUfJ67rDjRH2dXFOGdeu21QlCIdhPja/NEYTy8cQeBwR6D+7doDtzszX
8h2zGpawpZbJNOWdxF0s4Brz//JYSa+Uc+XfQH+oqog4pAKn3fSoUCHRtqYKkmhL
xd3ZQlBdJBjc1qHuJuNyGy2wX4muMHBWBA4OHJw4TQBJbMBcuqCUqyVYFB2YQLZ8
gkIiGFH90V67bN0Pg/tHqJ935lNHOKKRRnENz6NwHGg3aw+NOUbcXPVwyyu/GM/Q
Cn1hPmeTZPY3//SHI5/7jH1utucQVGh54+AYphfdU5Fjwdij9XbFzet8RYP+bMUm
maEHJjTSXJZTQQCnIqTFvhY9IkiJxHKOez2/bZVgybu/DGL0KhgNPZRarJdf6Wxu
dO2NRcIAi/biCwjk2geZ+OaeRiskqZJH50atbktNsUWNugBbSciIpGKZ/jPZ6Pv3
en1g45Nx7665mJX/fxhXktmRKNQCOme7287f0muubW2C0tA1c4+vbuzFd2hIkbWh
2s71Vk4Dh/RgV22YdQrRVi1G/0kMIsW/Lo+Inq00PA4mtikUs8HvIYL16cHYZaAl
vujJcMX6Kat/Hl8pvLiKZYRpcUOAzSrYxbPLVLllMX+0aThoru8gCFpRb0beXRGi
VHRcuHCniph8Vr2oorGiLp9qeppMTqHk4bi4S5t0+iL7efBbBQreeCBEGCN3FCqj
ygfWOqz1lxMq6IT8Aj9HidPZUI2OddfhLZlhc9FBwpv/P086zhB1EtmstnQqOZch
VQ/Kqe6aXELDKz5DO77XbmBuNKR44ezR9bHeGWYh0bJbrkvlA5ce3C+9gzrQlWaA
1NE5qks+cDIEk9HFsNfglthrU1xvR95/lwvieGvAE6PcpwdPHIg3/0rHvxBJoj1/
iMpD+gfOmzLlS0Y90UhdzBrbEJUif2/x9ogDCmFz14eLslkeAvUezg+sRqCrK913
0DPCSnD8GXAaa9p9unDZQdt+C10a+TbF7TI54+64reI+3r4aE8quXOk3AgBk4Yly
1nmwErOHbqN1g+RtRRQlM+3yjT/OudFmFRdB56Arss1uSQMIs7EefZxz1lj2Tif9
TI/33Lnw+FP1E5mIeC+rK2jOYxr15JrG3Drwnp9X6wDWsMNnVIOhqGC0nDlDXgrc
/qpbMAsDKkKxVWh0YC0xxxDXv+QU+ZScRdqjPk+SmGxcemrU3bZx0SDWYyye676a
o1FE2W6l9WEDrSwjyg46qgTuHduZ5R1Yjk85j6c+wbxsVSgMoAaC6PdcQ5vxdD2j
QokE9JFB2199sFhEf3m29LFLOJWmmnY6nrJve6DkecYDA5QcJmFh+l3xbf4sA54t
jmdSUi3Oq9xjhXXEdZOZR3n8vqrVNnGzzFatPSy9WEy584qPmHUgstHLofxzGGs2
CVS3VG7xHLwR4+8ZTmuuKe92k8S9B0crzL+HnL4YCDd8XUoPJe23vx3Au9JuZdEa
AOkSdZ4vY7tdOmH93LsOFEuysXRCh2IYCGkt/8N8ljFX/8KCdXribKQ0d/iVXlI4
C/xMdVXOx8iJ/gRZFSvI80kNUH77WgtqAwKzSFaq5+mV5/AhJrwB3CcDxFZjS4GY
IfGIlMAX15ii/7xiwoxCdGg827tZgslxsWtR3Ze0EX4AxgDwfDb6fzk6rVzKmage
unaZq7SQbN5Ymt+IBKe/JLli3HbrPYgWgS361AdmcTjww7wO+w+xkpIE3RXq+6re
cAsEoC6WSB755zCNVUVtNsF8slEwVJWhdKSOEEAaSOJhIHStS9gGneVthisgoszz
9G8gRdM6KVbK+wUko+WllCJZPNnVemLZnLlX+mUQA5hhYYQwsq+O8qBMo1kbkOav
RJMqpsH4AyyIdDIKRXz4qrtu60rEYAocIfij2SKnFqtcZ3kk3RkRGxplH+JPvK//
tBc4/aII6LnjM46P1RfpZA6CS8LtUe/VaNvE/LpywEPzYyyI4OL01ZXobdt4Sc2l
DX1xkq3TMP0SGh/aOrJXvF9m3aeMfL0/Yd06PAnEKIvRxhIg7hNVvpum0clSSbng
YVLwCQiEBiifsi7U8uket7kLcrJ+KrWj1Hktzq5B5Z7/wcqCPW89Dhpx7ioQEm4B
61YdDNCpqhHwpRJt+CHMl5SCpALMeQJDTCIjeUyGd4ff9mn2z1bxK8pg6bYKfyio
J84U45NXEe6t77kXEL43FtbQrlcNCg/IT7TbDijpphMdtrF8UvCB1WMJEtPemrmB
7V0dfY1Dork0Zt3UDZx1k6yjetwL/RqadRs5E/QluZXnz8HmzGLafWNJGsjI7yLu
SZxwRYFFJ00QJs8WEF5myNxAhtSqKcC4Uxs850hmJi20wyo0/nrkBAy4YINzYkuK
G+XY4XDg8+CX7Up8LBqvROldaO8ZZeFrk52WCf58fP5BVB8LYnF6hZQ5ivc1KETB
/8IJLbzlHV/334dioeVudjymQMPNd61YNeSwXYAHMCpU/5vz8mu5QW9WizwJNzxh
7ulPAkirxveu8IOm5GRQZ/uf6QWDuuGt/M3BBgG0C/spnz/YGVYSZIcTkuh7HCaV
6oAePtRuJd1A3EwKDZkCLFz2AtBvEwFPLrPgvuLRFPGldRaAfkEYhHHZvEOErhNb
zF7OzkWi4UgeNTqacGMvV8B29uQqTvIxNvi7Xl3E5Ksy+fq//UPU5YXrI96pDwYe
dB9mfuKjn2xbxjZMCoiZslGV3ErJM9JMe7/R6cxG/Dx4Qw/gaIEjxSQlng63ntz3
65b1uzt3MNElOPW33SjPGUdAcHdlaTKR3BzgjQOGTB6xa01Vkz4MaXDjUOAhvHyD
abT/XgsNcOncfFlXm5XpuX6m3OcHyS59rG+X7QoVLQKvKW8gPm2jWvf0p6ovh+jF
yOH4bnh+K3HBXhhBlMjaup7DajxQjnUTqOfE0sStZ8fJCzORCYTXbKKD2F/RebCZ
mjBFeHkG7VmNGUuw4rt+MNZMmA2hcf/OK01rSqfbLhE2gskmpyStv0rcyJzEZO2/
n0kgF+bL+scOIYjMTJvX9gQhhLCr8glM895vejB+dgpOstvJsgI1m+H8JwrOycSu
sLDldKxoQHFjRjY1rYQWpt90GDJx53xRgX7RdlygaMdDuQK677viPMOdn4UQ19q2
0n6SzWHQfC8sv3r5CzDKpZkU7p/86C6yZLVvup9iR63Mbd3E4N8FNlyb/GQmLdwR
RMc/NmEs6+LDiaaY1DPvvFCdxAfzwULLC+WG25x8Cdekw9l28JIH6K/tHbrs3TcN
G6+vnE6BLyXZlLjQ5gR9ttx/BkN4oR4CyLDg5Its82KO2tjXP3Iv7Pm4dvV/rHM8
fWyNrtOE+i/bi6E0Cru3TUjAvRr/mJ8y0d4+pgRKBZG8Wm7onfHcVs+jFqvQ7kzl
VJIdNyHu8yd0gQVGzr3r7XnWxiLx2I52cGCqRK6oHSeHiByQ02+20J/4EaA5J4J/
eXqZok2A4L0UUGOYI/kq5KF0ihqBXhE1YTRLM7U0EeC9uJnWnLwbECK7W+PWw86W
svORCM/d1O/byz4qwpsSzzV/fHAvxCXPVNbhcAMOL+yJlruc7ct788nZI+ZH0dWJ
VJNVKhNmtEupHrj0eGFvyR1zLZKd8sNZvRUFe6j9o+WUo91o+S0bLgj1TFX9hbrf
uvZbO79tsNZ+5sGsypcW3PTPR7V53/ONn8ATq8yH3ABi74lAlJZDlA9BdmcBrEUx
o2lJiy3AgMP4q8vcDaNu6NeKqxFgjYayBsEM52tU8Zzy0P2dRoGABtiN5cGN1OFo
1za6gz3kl2U9abndyOAjIUgFDeePUNTSuiMWJ2JGbazrniVSg7q7Ms1ALyg9B9TW
gXHAEC2/x/SDMCTpjCN4+wPxd21UKRec7qwgrWZ1gwRJGPi4ojB2dSzFHhXS4rPX
XKUhmFuK69+Ja0m40fHXlOWSTtrD/0WIB+EDmibSOkw+nCjEugRo+BNBpxYwcDlz
8I9KqljS6NpAPkgvie0I3RE/0artJqjRq8nKT6LQ+Wtt3hOGsh52P4lbMpb6ClzX
UO6YLLSF/6yGCQSOVzu931RPSs2/5lzskBbQMhwl7MqAlvKphIyYX0uM8RK9Sv2M
2g8ESdmctMbWBUKUgSvvl+5mMtK7zGWPSul3LQVbpyepQ3esB4rq1H82yaGfwSIV
i8ETlMFHv39ULwKeDP+IvtgFf9h209moB5akEqOKHPu9n62nXIBS4RV1YjITMDoG
epQeu1HQZUJxSSax0Lh7qKexOuPM2h4jEVme8WrEo3QqsxDr/U1zQ2jLKtNQ3D0n
r2y8ArnApbm4SYTnaqYl/kd8QL1D9Zw3aclP2vUc8nKT1fOur5FI1ly1EgpTXIAm
RQDRx42MATR04eDI6gT8gV/lWvxYYW9b64om2GnzyqY4IvSYwTwMJroEvGq/QnmY
iaVZTijUqZijQ/T/D6Q6Lq6gJkJ6TWr1JwpdFc1DnSsI2ity6fC8wYA82/F8EBWf
lDcC2XL2Txh360J9K7dJOU7KAWgYyzSQNpzEOv9uFBwlebw5+a4dWNldcpfIc78H
60eBcOQOMtHwSTxOUoNzfMsCEjryv8pab6DyAqddOMJIbJ+bxx6aI0Gmysusqv/9
Rhb44J2WCjeTtBdOoysStX8EDWfvygLSIFycUISZjKoNNP0WRUNcmjGHKM1s8TyC
965aiXMYqE5sz4U4DjuEITF5w0EpgQtpFay3EHdNZjrNtXTh7x9ngUSLrmapP7gE
qZU9mmbAF2SLZqradP/3nnAQ4HdUFFVJHuX3xdBwqq4mdO4mik8nUvgaM0mM+3dw
lCEgnNwoq+GRL4fnFANwJrEmSzFqR3s5fetrT6Xck5d4YZRAmFc/ZBW8Q4vvzKqF
z/9udLmmP1bg7Wl8SDi2bxGpxviEsMz9iP7ggJK/BKs56scbazp8uAZOfIGA2+S1
XCGd3/hQyFX275VQuk2+gieVuLJTOa/f7/BRoDVcjYBDC8iz7gJsdFA6TF0q98pO
NNoZYUXRQjksBoh45iZCQC5zHwxHaoicXJqe1atwwOBFkIy2JsOx6Ro7RlftWDkv
RylBDnldziBD8xGZA7byzwYgwMrgOOs307bSQUg1Pgreq8SlKgwiW31/+ZW4mNoM
160YN2GtcUughANgeYpZkGI86ztktBU1wI1606bX+xDPTaIZXFe5lk6p0SOXTYs/
dlMu5w+Mw2yo/M+8NykFwFzjYbvcmX4dCbnT1FqN1YDoMZvvHAzi4Cw8jCu+XfzZ
RN/8pzOQACgSmMlG3Be+duEED4lhH59b1BNsE3VAXGYCe4qJNlqirVqOWbERK++f
JMQf2E4F+a8UXnDAPVh1jtBAOUj7N04S1lhZPpmU0FYlrVNlJPCYAwfU92iDmtek
C7uM3ciYnAmznilQC0UN4NKJ5vwe+mlnpkGH2E2ORYSHGDwmowe8XF46byX7pshH
erhQXiUgNy5tzulXLoTuhwOIpFryJQE5CP4O6sDkfg95QCjmGbSNXiz+K6RUXM90
k3EkDaNoDeyvuyhCrDWlqK+NInfFar5dOXIfpxEwQDKBL8zOBpE7u/Ae4kF8Ezm7
jIegFhnHv7aCPMAcrh67BKaM51yJK7pqxejMf/LosvIcp3nip9iRzewRJpbD3ZO2
DDuNIT7uGt4IbnGtjfL5hLc1EGMPWC+NvcUmj4PF0YdCoilfYmqje/HJO2TXhmXb
RXhNMz1kxfOosRwa2l1DW5UFdVkyjKmAlkYMq4UhHk6u5DWpGVaZylvhWfg8fhUz
La2P0A55/Gtpyt826pD/vnvWB9CnWcVcDEI6ad7MimDOzlm5b7jVg71lsetkIF1E
dHyxVdDYXtfHq90gLjzSZxhqxH2auHoBSkiOGt6vdygrIO9BLD4nA9DnW8D7F1pq
QVKy8jVqMUdNT7u265cfGcy2yKBV5Y2H7pm9JCQ588WGTx/Pqyicma82jYv1+MfW
39pk13qJ3qCoVeQb4qmCI7Fsi1WiayRvYzAME2itt1uu440QfSYmirrKvEkiGvNx
2MQDB02QApyIanBlfzlI0umsatGC+yG6jXEq8Aw3vZnkdMUHsrOmpLHO2vvtiIvg
mZKEiASM8KmAFSbWSMvYrOEyEu1CbANDBNCJQquYv8Vs7FOn0UYCnLHTDOHBh7Al
Vtp30ldYgQd/OzUWn0EqT+9mjPS3OHibh7jLF8mfQe2W6Wr4yp5zT0JFeVKInDA3
He8LWjz/k/N8efmlEbS7YarDFteecB/L5OdJVLSkeFpqcF1fIw3aZrRYgYXBu/1l
RDDWKQ5Oa4zT5wYPZP4lvLoYJh9xPAKeBFtkMY21Aw8RFHHH7cD9o3SHNjR6Sdlx
/j3OoqTZFuLXZ/S6CxxiiIrTI0/eFrnVOdg3rvAr8lgh1z2HVCYyuNGST29I9wrr
N27zLmtTARkzoigS2FNvZFWCZPhdFUbApms5/Q20pjTJaBdZIr2b+kYONyY4+Mmi
kJZ6d2BJunWXsupnFSHoZMPW/9EX2B8kwEWbrwhIWbMA332jue+KCZhi/xA0VIoH
hRjipIca6mI9PMgZUNz7g+cvScjH2T93hLpgqWQyR493p20iZuXUIV+a+5f3Vcsc
b5JhJNWweJDayDi8j14U0mb6WhhuvDp41udDp5lnldO+rsaFDYTmRNaBMP/DHZ6a
cBiMsXpdDM6Jwo6gYb1mK/e6RROIZ23nOIS8iYuKLHHJx1UKzHAbaLj/QWo8DH9Z
YnoTQtP7wtiP+2WvwbcOrn0aE2KmkiI7tVczcElUuMTajPgE9MMQDrIv/SafNneN
+nAzIieqfkLCNS/eAm5MQUPr4spCSvxjKTR1ljHEbXu8EjWu339+WzcCvbz81YZK
obQ0Op1MPP7LPfl4KpLlGF+P8nxyIeeW5nYgjX/qq3uxfxoGMuGWKJyjTFx6fjIw
7DL9/WdwZYgIvVGHJsbxasLoi2qN2F2dwvW/4LeeGHTfU68GzrbiBau9rH/+VV0a
jQ53fc0Mim5lbl0L63UkvKygauUyKyLgh/fgf5tR7T0Jc28DQk7ZNOVbhao8isdM
mMWBOUWAV/pCmWxQCsJ16WFxL4AdexC6v21d+8UIsKnDc/b0uNBYX3NDBxsMO94B
iTXohwz1QkBAD2fQpQ0YkHlRgl8VSsCNbt6fCppiE586LExxJ3NqTgipXunGNDRQ
0Crl2JCM4mjp0LAyNGlZGs3GJxi+LcHezIkHe9q25xH+GwpZrDjtK/QEXbSLiZOG
9WLQGq21NuEH3bIJ7e5b0esFziyfB2JOdR/PYNgPfjMiR+7u9aPVGAqB/93Fyaz0
Iwy/RDQP19gbjFzouCex+uI5v7H6Imoc/vOHUYoY8oBdvooe1bayqGyIEXa6Cc4R
JDof4FEnTwZAHQ3bxLGoanxWTFjfCH0YJXo3TYsDv3LuuxJbnbtUvakflqpZPCE4
OEWle5nFfQ732KCwPSuFOMj81dqfxOjjO4qKc/aE7pM2Yj9D65mIey1ceYmCk/y6
RjiReqDdJrNKy0WV36kquHzCGdI/iPlrpTZTqn/myL04t1Kk5+R2b2iqExoqHl19
xdhNOr2NcmCm/tH98+diiJu8za7cYjNlJhbMC07VPSbjy+W4+D1xGhbpOy8esezG
q7JqCaN1+TaXHXZ0vZGd6kIxSnXpNxLS6JCIXbpsbcivgjRKKLBG7Fx8n1AubBly
Cuk0WAQdqM9qfTtwjMPBo91kM3E2hqirW5J+62ZQrxgFu78+x728OPSoR0tLZnUB
WMXyV/5koz253Vnew6qC47S5cubLCw7B4NR8n0OAsBn3ypsur3ZVYKpfl94hzVqv
VlN2rSUEvAygyIm3JEfy37450rJ3c0nTmgTl1oT5HBLr/ohKHxOgfDuV4iE5Eawp
9Uow5OXzzWWhlxImk3SV4eBfXx9Dl+KZeKheKm4FLhC3evNDxIoASffpX1tAq3G6
1cBnEwPirejFvWEVxTvoZQZ8jAT2ZnWR+cSgFfNvuWfg4OP0f/h7ZwWiOzDMZxkX
zUnlHmR9jiy35sd9YY/NxbJuGA2vR/FXp1FByFCXg71Z/jlbJmZq2/JlTKwmcHig
GvcEh1QhvmBoHRJSpAyKmye9BXnbMNc7msSI/MxJ6uGrVch4HmXi/Utd4psdpS68
yPeRKVjFmHSS4NmFteDlP44T7qn3n/raO/w6hPY+sIHVpm/VgdK07Fdq30Ks+T4B
jTA6pbx9eO8kpH8il66wNluQLy4CMG7NKXsNwRjzDrDbcaadqKCEoXYeWjHjI/+E
vPLBlONDFFs334fFaFKsUbhlsq/BJS93RWgpoaBc7tw3CCoODPQxgQ3TmMIXSrYG
syQRBJWHLDiX8iQL8svOtakgbpgOv/ps6cCPFh9mceDJGwdrihRIGxOI5cG0yOIB
j2Ul0kLz6ZfpJXil725Rp20z5TVN5eqtEbf9f2Jj2CznafdbvhPqqqJu5RvvI1X1
69wzIF2fvZJGiuJtYqN3ibxSKFISIJ8PbSJM6Wft+emeXI7YRYK6rU/0AutwdBXv
1+hYNUIlUf2Nufvj4RxVVi2bY4uIuNY4OZK7gmoDECSNi4PyO1gRNVXvtmuzbve0
vTm+rnh2h5yNp106P8nj3AGMB0r6OlC4Wu4rIXkI22jtUZ+kSvcLu9Rc3v4g48Uo
dl2P5sUItDE/yc6pkFKStjbSC0Uki0UatrjZiivASxSGJgegR5OP+fTfXYClA2Sa
xssuogokVpWb+/pge0v1OrhHciZdOSH3WlSgc3ts2Me2EzqxRhPdt4sivZDDQRjO
Mz8kIl4j6WDfJeUmDq7RIrQZMP2KngZnrQgiLxL9RXZsZ/jZx8JMfDirtCQzK9O3
WSmzOg4Kdlmz/FvMX3+lGOGRqCfzU5eOMRTa8m3QWZrGORiyYWYkBbWEun5XaTh7
rM/Uz/aWjpXrJirDy1jx2fRoVuHEQ+biQcQGBtcshJ0dIgqOILeoPQxGw4QN+oHG
xq3UUJqwj+PK2vuABxIrK8LGtHPqWSNnZfysHP4f5FQJtuQZo1bVOhEFTpGXOaO7
7t+jmzgIpPhBLy2J5+uKv0znPPt42v5fFkVaGYMnUXRJKlsScgN6uryOCbGLiO8i
jLsvnmWeADxzHdWIB/SkL0PN2PDEZjBFiJ20qnd8M/++DoNnAIEd5U8g+IYD5Zc7
d8jtzMq1hGLzaXo1NgVNu43L2IAe5HMk3IqdG8Wm33krfda4qNYmE45juK0kpwUv
QK8yoguZdNql9hMv2Jz9fOWdLGRoWPbkX5lDBIfVI9IQwWe6nBK3QUGvsaG9kx3I
TnMJd1rEOpKuaoSGWpDE+NBVI0lY5t5HyJMz1mUsNmF7MurxFqXqWL+N0YeHtHfg
AHTFKiSmmB84dre6rHtV9cU8UUKeNo+ZlaRe6h+fy8SsoMXLUWTt3QFzoA3/GtUi
/AaFwzYvzMJroY/QM1WtuV7lIZAvsGYawqjtcTuE+xbr+j2lUBI6tMbBWua8ASuX
3krj4FY1rkSbfHeZLH5E8CeRHlu9bq/QAXdVUas8mGt2e2mywnb1H+Lh/tfTIFDE
Mc8J7iOAY6vRuIjOT6/KAFL9q9R/ORnSOl5IssR3PwBLJWcwZlisEvELSqX8SwPS
CIS4MTNVmenqSv4+FLX353H7dKa2ZAB7OAT6naieet/i6297IYoRqWiSKvYyYtac
gRj7/lkPa/FqN1dpCRp4YePem0xDi/53jIau8DDmO9lgEMtHXOqqDh39+eKUBHn1
656VGMty6GeuPj3h5GuoKkFCpv+xJLZN7o54HZYfEyOWT+NXO28ZvP+IIiHc9NdM
+naxi2RFHs/K6TbusZ5ldffrh5c5FlDMgRn7iWI9Ste2tLF20IGNoGcpsAdLUKW3
TCw+7tZVpbil6U/gHPE3kqj/3v2t+O8+IM3S0fcRbyQ7KJ7Ole8BPbttwf7Q3fBQ
ChxMRUobXV289uVoGOXqoxK9iFMVotKENJRqAu/M+pM7olLJxbJh8jQ+NxT4krVi
dKDM5R58Xef35D4a3g3Caxf5PSke0msLUHKH+put0mzIC+VYOQnB5t/rHTt+TLmT
KhwPRhykfYzCLp4cRN6kTR/BM9IRS3sxIuJG0GLRLDCDRN5dBwDfKT/y2wBhZj4x
3rYRxMJ29MWie3IpWPkSqk2sYNkGrHwmYUy+UumSrFeeHP1VgPuy8srMKOdKY3XI
xmSoTvTrwmrO0PMiEKEqDnDCfJPnCNN5qwq7b5FBRRbxnXcC/44zTC3+s47U5I9T
fWT2b5NiA8yjp2RX0ZrUhg6zPHE1/E6Ot9clCPPyIQfpwhhuzjIqmeRN2YDRKrC5
4LeYi/anJXSrjy33L3f1JkyNi4gI+tgzOGKsuBXk5fY+G+IYsoK1R0p9+fGsuMXt
P8rKbdGWvuqoxQaaExkkaoYIpqdh+I2xW41I+3XBeX6nhKbPLNyILlKZjDVWfAkp
dXS3aZvv6O6URPOvx0r0uSG6ZqETyIDYFSRsI1ZQWnmfHYN5aX0zfVTmEE56GAEd
9b0mbt7Y6f4VaLz+3WcpG82yCMS/L+bNin1fI/hSzAkCLBHDg/zXZVqGqLxTdnGd
Jj6PbefIFcdWm1uIsaJYR3A+uPrmEdlf63oS80mTLWn1PJkOw83xl6W1U+p3Ko9T
J65a21v0rrtRiDpsQz78tu109tHCGK2G9lPMPMXJBzgDoOk6yDJPJ06p/WgPnkga
L443BIiwFmHrEtmV1rAcl63xSNCYaVYZw+QhwosZ847Nou9pvoPzYpzcqDCX/Mti
7zTT5cOAcpia6wysaGSLAK7r6/Bpy5Eee/mSm+U2lmoTCZAiKHlxxvxNILOi1z8H
rZz62Tm5uAN3H834HLJfSTEMl9hPxel2M0WcAIG70K5wpZiBBuuWhuD//TQK3J1O
/0jebklgQF8GRvSor5w5BX/7W1l5fdDWo6/eb+g9LSezgOSC8g95WezMEifraVDq
IuFkLmAgsPUQ8ugRoXvdc3lmiE04mPaVX5n+OC5e8lmvHh3QhSUKZvr/rNzVuGLq
gmpZXHq3EhSzHG9HJdeEtMNmafUZoyukm54Y8IncPYqd9XWv/OCqNMYcuOnpNFWf
i46M8WckOlpOLmftG/48xGKFTZFlkr32/v+C0oGtpfuzpoRl9Y+4fesJtlIso0nK
EK8WcwylyUx+Pzg1+EsIMGuyTPAJnUGt4oDv72z4QWSP/vJzj5OiN5Ji3A/gsRDK
4U8Opi+8ptSfQcppcQdm6jmmEl5Wx/qZ4ZDPv+v/kw6n26+Dzrymk4qaED/kBdyU
AaWGDxZDiYDzZbZ8FvXOdoDkaEHEw3WbW2kBdSgAa27bEUFTC9v6HSsZLYuyHHRQ
pXw2/CPEk7lp/AMXVKYEazwhA75k9a9dUWSameunSt/olXYzWzlK0q3QtWPMbbIc
wbKYmKNLrMRlG99xa2gQ4Q6RGCGjdC5ivfPe/WqbQzKohzMRfGw03lKtOCZVmnDQ
xrTppAyRvKf0n79Oa16suLqzNxxd+P7ZL4qHgWu/PzugAk7tb3vJXatZZwzG9kXy
Kz7zRNmJpXSnM6O+o7K7Gr7cpY8sLYVFoSSHKUSK9S/nkzX7//NUSLswA3ZxDAO+
O+pnuqlhh/SgB/wT1oMTC9R4pvP8WAJ4bSOR4NwMUPFrNd8s20icfCD61/oTjq/l
acmkKhEzU/RbcprTnsyouanXI8ZM9FDMuc2o1Z/wSprhwFpD6IEq1tZnhbmRvtvk
pCFfwEl8pYQkVaCWpADfINeqNvPj2czmyFugTNRTFe3jsaYIVOUPBs6gu7pQmlC5
Vr4DKz6IytrXFTtvoK1wffaxVr0J69UwrVAIOquuepdAClhYKROii6bJz35+XshG
6FSYIUAG+VHEQGEmUJc20P8NUyAmcXoVzJxkIHUZ8VAmocAalPD/Udw1U9nm0V4Y
0ZXMy7wfTLnVmoIDkvVz1XWG76mhQ0Zg7zY6kwRkru3wHfrwApZ7qZr8/1L9c5P1
PW5pGwmVeC8cOdx6ci5ZG7YTU/QTCX1qLW4srxAKnz7xLjNbM/Tlmt75r13RoGnZ
YDtJ3WanuLEE+0GMDHQF/azNZhiGcuiz8MTIRYG5BL9V6eeAJLMrK1AsJHv7ejQ0
XCYjjMbQhKNSycA+xPCBu04alAsNNuhHl6Eqha5itMyR7UIdkt8LmIuX9KDiLF4i
Aiat8oHG37OtbiDxaKYXVGfj4axP23YYodsZiazTHoPM3RcnaSaJ7RhAHhCmiy+S
4kA4UYHg/fKWW34R2qKhCN4TTU6KMyS9Fti4ji0RWQ/8JzCI0uerT/CLLqsmY9rB
kY3Pse0A9ON9nqu9yC3P4GmGJ+5ZslMIoOgGsw+f2zpDtgjYpIGcHi6r8nrEEe3w
PrGOBsQglNb1wW0fNGcG4yZF6SGcQA0zOHEfq7sbbUWLNBToZaYb+90E5lBcBGQe
SpBUTLOvf6dIO0Cif8xAjwtbAsdAGn4fIiMpwMpVt1mNP+zcfG7HrLINBM+Uvsgv
z9zCxlJ6jQ2h2VUOT/L7jJ2Ji9VxdZF/5zJFb+iuEAfYZ+EayqjuKy7i+5LQJQFy
lW917uAgWlJWleelaB8xnxxmSTng8MLlXKelYTf59eedKasMvt5yStvDywsDmRAV
ADPIs8pQUtqFBNy9zFCwx3SH/oF7fx5lGPojJD3lf8jhBvDdVQXXlNtaUOyokAV1
zFFjK3I65FLTO5hkcmIMdvRb73gaC0h53HY8ARreEyWdC9dHTDjt11tca0yNfD05
pemPeDA5qNAYDwsyy//RR2ljlXouhZFOJWbrHgTRKGpmlkydqRkpEQIjfeXiOE9H
BUvAkUm/6jXCGSHOMYI5WViLYWeTAcYFzT+06hxFPmCOG1H4tBzBps9qtI9HeIgr
J5d/fNsRoHx+h8zkT+THAEhmg7a9ECC3J8dOBqiBplVzYGtZSlzSebIdjsvo98Io
sQ9m9Eaok3ddlU/FQ2gH1UWf0x6xR1tJGQvaxYJThN2O+qN/ERE1+dlCxANJInAD
ytEcJw2MmIDjnI+tuaOqZrsPG9Jmim8jkUJAKK0W0jWk4mnDsiq5U+GFiAetd8Jv
Y0wDKlLpTZHl+IyvanbwdKUcttxcC2edwJPzV7wmfkB5TnEXNesd0TTA4Dkh8AIo
6n0mth8UzzzM7XVxllbRZDKr2gnXFvW5UBwTpbUR2gE0zf/lAsJuNWKqlMCGvslb
qFW8ssCExTH9q8sGgAsjdGY2zL5WlwqrU0fQG8TTr2iP00k+c9rGjGmMVdb+7CPZ
zeBb6mHdJHcyo3fxTcvM4IiAgIAbzlvyfibjLPZI3a8uEz6IIUSJoBJ8YFhqiQSs
nB7/6giKOhmEebffIsCGKT0PiyT/20MPn4kq6e2DXzL6vEvD7buUlmVDOTFKF0T7
2gm0Je2lDYJdlxgXwltYSTXPWmbY6HwXjlqU6Ltr8GcXvo52epBpg1/IUXAGgitW
46nyOEKZa9kbRy+dO5zM3FfFeUAC4cGZrGNlCszAxISCPyy3UOWVRqwUa2T8wY1M
5S3uqvDxuypfKgTwR2WTY0OeTbGIlSPc51Ak1m0+CnfzWYP6KBQ9yhGWv75mF61c
YBL85HwYWSMB2wis4JlIPP5bAVqcV958KicQc3vBylrq5atg3e2di/YZm/lI5ruX
SgyQAEged8zEc1eCoDwt9mgMv+XKHre/kV85SLf0T3ZyhbKHVwE4+LDOAG++p7Nn
Oe764hu4wGWJJirwRYC6QR0adhusjxvFE6rB4loSP50BsThk4t8lwHwLgmLPPBbs
MTWGfgAEdzg7s678yinVd265nUdsqdYzZ/AFKPWCi8eOENo3bXVnUuOe9+ubr27y
U8onu/7SZkA4DyMoQo3jY+uQiLgSQ8+zeHcTcSLc0oJLN1vqlDhEXldKFTfhAXHy
Nys10QzSj9a3guYQm4lVIbhLW8rdcPZPjUjDmLXGtTqStLBC94/fAHfcMiXcbzEE
ocWWL/wpWVpm4gQsll+9sHJwVgU7JNIwBftKZ1wQEhWuPUxjoh6x74qcG/bPrUli
N6K5sMaZ5GWftqsrXbr0MnJeyi8Q62P7PCzC/eUCM8X1FPYrumjqtns3wUqEVQkm
cWQaOGqW4vKsLmKpuInVDmLjYK0Gdjfykut3/sR+fJmhUXmQyC5pB3gUut3uEVZX
Ele1FEA0UuVpCiXu7ZxPv6fluckF4cwWr9hroFv6mSjL2t5LuuoLFlD3vo33nKer
8f6y5BfkdAqN+W4PfPVlle9mngTZ1HrqmrXKVI9asIeflMb1C2+ZWMpRseBB6mRe
zSBuOI+OIekeUak8p13slIRoFQzTQiUuSP3oRTi0MknYchHbQOLu/Xe2urdLXxWB
NWJdh0bu6BREHWWVm4XsCikecYMz3Ds85q8ngKCpAsc7Sluss1BovTxMTWVhdZgb
q5L4GlgKo/T0u4xiWmhlXLmnklxzfXIIePLnvoAb2bXP046QXSzgnomPAwe+BIwp
r9cMoSxagCjPQgJFIGsEnZtFLwSyD9l4IjqvJxsnJM/gadHRXNddCccrEuTWAnL9
OT0K/mMsTldGRKYpxLfb/WaOelqbko6Ob7VWd3IgJ6KG2L4ENA5Vdg4z+8PpBrnR
Bbjqgrt2bUpi/1yR7I+lS+SGj0FEciOokLxrzsJx/DgIDXFR8fmewsfXR+chs4Jo
CCD/6YBX2Pj/zPQIegfzr2oC8t8cd3Lu5vJCtYWeUZhxtqwZgVsoMUI/7cC73/67
NeYKKW6wea4JQfmS7rC7KvJ4ll29wHtQML9rg4oROkYNDnwXjicNbdIEdVfhnN8j
s1lk8C69s7iAUrkpSWord/jfy/8MaYZzojEiu+H5M6pFvMfAe/Tim2Wa24SF3OEd
zyzagn5XJqcRKjK5rj1PkcZjBEIzINgMNM0N2X6kqaXQxYUA2rM0ZBuOHh31imGf
lzhPGLTvoeo2psNfpJpez1vCHcS7WTRJZu8orYoepBNmVLhw6kQn/9CCXFx+peK+
UFrUjPMVYHKc/2jZq5VueDrSIWA8rnhcHNra0kDbLPjXKAQVh53MBj/T5XJVjbhQ
1iVSBskhXkPJ42VDoUN1M3hB8IQ5Xz+yc3sPgGP7YjB8jYHz3cInJIa1b+mZCyTr
6yLoT7eClPolLWhYWKwqQKmr8hTx7pD8xlOF8VYlvC8xHFWPrl+z4Oev4nenEcD8
TzEsOF27A6biDxkkCRXia6dgU8L84oENM+ywT+zyOFVAF7xcLxdrBm/gdw+HzkGP
lyRWY/P9LCZyQdDg8pqt+g2GRtRn3QbSEK4+qxpPvdvKL/8NdgBXjRHc3PaK25x2
YHjD+FSfdJyLmdoyhaRpYac7w28NszCewZ1oBDBy9k8mA06c/i9bIQewYHYtgMKs
YgI1zWeFqarQBt4Ly82e4qQhfD2TL2iKq9lYiZP28Ogai31SUJ+b+KGntlbcC2Kj
r0fv2MKYBGNivgjXMGVcozHgejMqZ0NxqHUUEnB8ndGpbfthjlNmf9TceBYz5bGh
vjvDD/JrAmiVZAUpUy+Ef1eFPUr4zKyCB2GGYSuaFeQPRWEKHyPzpEL3urw7kIQa
VK2F1K4DqhTJlW20o+u+n7K4ARr7hu4JId73zeZXNLuaJiwNE4ANtssV0XdHSK8i
hsV9+Zc9AQpC9nHDO/Knng68DYDrTbW5IETAiH97zRzU+wbMyxHCB/u2gAnROL1S
ngZF9qvmF2hSIF/TCr6mfAMbFZ2cN44ZuXIdlKaASRblhCBvggUPG7ws5xyw7YVY
IWr0K0GkNs1n4v3rm279qYxJ3nNcJ4PqDAFEPxgz4EcB5eBo2IWw3+QwTdNvY4F8
8pFVYe7JOxqQE2of5hhSM+aKsfIWkgyT7ZC6J3MYEHGXz3dxNoWZDiIbvcMp1J5q
7oYEij8OQp1IRXAjGlHupnSASnpQGX/H9xrMWOtg8tLSMEHbV4Fu1ZXgWHhk20wU
iw5MfWSvN/GWNy78EpgzKyDsjlVp1py6ll+caNR6Xq9SL6HnB9oF9NwUp5x/UAyp
DuCqXnYRqiMaPHoo286X30zk1m7W8/zyuPG0+NhwfqYEEag/DNljR9TZtsvi+64H
o2zF9LcQtrkXqZaC9cImramBV0JG/ii6HYMZ+vJtrg2Dh96kLPukoVPrs75exgnH
LlF0uMjofWiLiKTmkjjaAvPQBEUxJaRW04To38QbCpL6FFMQfaXZ+ta3bNCE1mmv
zEbRw6n1DQUjjocgv1RFW7ZyxjKNY3RRR+U8gwBgWe8JRsvLbF/26V0bqLsIm6xJ
QtDX+TodvlfTm+W59577mAUnrHaZE27+p4oTw3nFdqN3sQlzHZuolZrgpjxvUEak
gNfKmspMi5zw1XQxFzNEuM9z8/XvkZZF3UrO4sLHY+sDnJv4gPIAZ38wchCWXzTT
ykce9exmtM8SX0vngdA7Sb2GUoPDIpnmkEldsaJhIHpQvLcamQuda9s0xouqnI7V
nU0DLnKp3ca3tc2tK91OnHOcNqAxPmHGA/zoLkrjcVzuPLrKTo+LUih1VbR236VR
dFKrWOgDA4OUapA1sR9PHQou4GBKKzOPBB1DlzquH+kpbuN+QEk5sP4j/LWwF8zQ
iDGxwBIdLsrNiLtAonSZAhO05yCNoeX7ys/4n1CBl70gud3SHnsy/VaUPDaysWdI
oZONLd+wCX3hSsG/NbO2c9kR3Q0v8rTupDGJBWD6x9Sji3Mdvzg04fonNWkebz+X
4PN3maiF7011r0apdpwN5yBE6eW1FGjc41n2hI6Wy0qwqV0L1npGFth3/ECxBN9S
Dsb/KRjKfdr8dxhWUmzlT20byGTUZU/FE4Bqt7zC6wRjHVACAss8bu/VVrcFSgvv
AHSmZpyoa71KC8YM7k2dFlVNXHTqVdbmXsnlfg2mDZPOPSqbegTgJ0rEK4YfyNF6
Pht+TXu0kexxFjKJTIpSDyBLgUDmXb3LQnxU3kSiIUuT1k/doNKQSmCkVWpDWydV
7f54N+huxX7WBQqED//8QA4CLQlKqzE+HP3goCNhE5jD0+PuTeK2fvHpU7Cpqlc/
gd9nyvsA+JoJ8GBsk696zs6aMmuj4VaSelD+widsxuG3DQy0YsnqNoplBDMkQ7Hp
pJxtWNCIORCzdepwwvIPADGMMqb9PeykzxPTVPGusev4AnUawp0v7YLlP8Fm9ZHX
4ubcvpfAedFXJSxvgqv9IJlgg+fYv3rVAyAmHN9QmF/8dcPIIQXnnoieelPg6jmE
/nlnfvTfvtdiMthvQaWETRi9JF4KFdxQP3Aqed7sA5lwBmUqgNt521Ee2y0K/Tq3
VC/G9ijGUlM9i/9jdteh9gIJ0Lr9LN0Tsp6qrEL6Mt/IiDgfd9q7wWYkuKKHPMIz
qAYbhrpmPosHbeE5ZrT0BqbHESuEQo3pDGpT3gt7WaK4yKCJYdZaPqVbQm4j06eK
EYr54MH0rJ9BGxjA1kLQPPiy+9Z1PYh0aOYSoI3rObX+LL8muTh9QHkHLsLSvtfN
PFbIfYo6n5SJs/Ie98zJk86+4n+cYP+bXJ3K1cuR/gClO4pNezdbsrsPz60fncaz
zDB27BqX1CC3huhgHnU44J/3CunS7sSM63EeFgqnzQS1vTmmBZmHO7Wgr8+hwnCZ
UE6qYLPrkw/NRiY1JprzWL1gQpwLGrtjg1PahxQtY/FOjsnSxagVXjjKY9dqGwxO
PgQsCkM5Tk9BROobytdJXflZP6UWzbHNNC0L/3nIb1M3LByM9RdYbVU2u6Wqdlas
BoYtJezhrlpUG7PST4ZMq7dRSyaHZl3j1V83K6f/1bAgcvQdEz5W20ToQHkd4YLb
iCLf3CWENk8ZMgfkgyVcEqC0x78AmZc0akzukBRc1rtVkYki0S5VT67Rcp94bx9y
Wc3IaUPZUNhOS2WAc/qmJSq9lanR8BH0kkxnnrQTZGKAq//H6hmvtyIdMM87waBQ
cHEVLA7qRcxIwnPt07kcJmLIOKfJnqP3QtBYay4tK8GTCiKJ0xxGDPQdUQS+xKwn
jTvq962z9OG5GSAfu7HOcwQ+DpOJwF7Xx9mJutR6ZP0tcpgvcyFMXwVfsdgMjx36
Hu9QJRxdgGEyhkJER7cDNWgEyRFHuGaxoARf37kkz/o3iI5mjrrXJc2GLPHz02CH
rmWWsJuMXpcsQFT5DZJtOY79krFl2ftzWDrBowj12ljdaR3OaFVG/DsyT2CbkOLx
jnfZw+y2vWr6fBXneSvlKeGiwLEsTuT8wUKt5D16+RXrdED2OOw7BgniWaY7X9Ey
NxkV7KJCV2bFhtnfmdjubgeTrMotfJCwDzDtvHKlkRe7Ni4Q0oOOP/JPRVNJ4e51
plq/4uSUSgYdbji1q1p3hAYMiry930q8HW9C6UqeN+crTfeT3Oq+ha+du8dWP6Iw
GCZZL5T7wuwi+kMsxk2I8DmyREAjs26DC+GhtjHbN5hz/KilHQH1PeoLQbpSY1O6
rCfAfbQ5daEHTkHYmrVJjN3pxMCYAjP7HEqR0lYgj3/khqekMOj1eN3ue4oL63Ur
sfua9ZZRQjsdC7bCOUUj0IR9ndGVyTGN2L/D0WFrCWrLYL1bNiU7hNYkWD6czg+n
cPOllZavo/WedoNr+eQegHm15YRGevccQBQizofidscHgD3zzo7QhFKI/VnQ1zzf
cmU+spYqjXiBMAk1h8XA8vNm6zRJVJrWFMLdGHVSqISF2SKQ/+i0PifkYM4NOf6F
TZWH6TjjJgUZhgh+1rf1UnGfdENAhAGueyO7KirvllpTA9lVj/BCgw461zbAhBpK
jRs/vWhi2mHAvJhVISaQudjbd0pFTYOpm83lv6hU5RG2gsj6lRmD42aIpUt8v823
c0Wg46wgoOz5/nb5qtNLHBZbdX+/DrAoe/VOFuAr2KGwAM6Ax4pCfhaAyc11ath+
GZDRxi+49k6CYwj551JmkU58cbvmILPVsRE6isaJ/FFd65tZho2I3/Ns/U6fxrm/
UoZ3joHpZ4NwhQRs3K58rfcmBaNhY105ll40A6EcQliZKYVXfT1jEcm94a1PZTGi
rBnaGp3xpAt6zuGvHGbSUhUeaOtM+rTjoxeBod/ms14G8OOqnbvhm50SlLeU4UeH
e97G78zaZtz5NmTXWSdtACPhBEsYhvci3YEH91cBePrwjra6EgZjVxsZ7ADs0+cJ
hv9rUJA41i389+W2QhskI5zYhxct/KJso7I3YejHdXrMQjGPm1Id2od83X9yEpdP
jHqqGQ47fK5j9aaR/B8WxaFgCC/Vb3IqT+yOslKu4OFP/mUhYpd/T76HoxUCP2L9
7UyRzqo/1mKfM0bz6H3SmsH/6z6aknT2npR4cPHSVa51FtQYgbw4u3POmOdvOtIl
z4cCF7dS0RR1pL8Blxg9KREmWSfL5q3FrMONTlVQV9x2Uh5FytzSlH3DtBtqZIYk
gk7ZyOKUv+6w1HmY6ia90qrhKakzf9GzOuXncaxpYASVwPI4jyz3Y1S6qfSWsebC
Xd0cB/BJp3Txb+vawDuJHD0y16AxSAzno30EHElhlOO2vpKfcYwqXcelT3KrTGVe
NHiMElDirDUdfSI6Nhl+ua/i0ye+xZwuO8g1igaxN1EW+hmex3sgTivUndhB/49b
paYHZSuCVXDollPCPQaiFgr7TzjOu6Bsdd5GRavtF5We/eSlwORMpEU5wD923nDp
0Ts9XWQcSUVXbvuSgqGNPY0rujSvdpq1WNIzhFDV56JVoG+BjRie4UKv1g6s0oxh
ciCL0y4d3DVlnLs9sZUGG5OQvtVw3G2Jc5VcTZ2K5MTkPLdv8jENUksQQaCNnCNW
ZyyXJIoHnXM6qrf6uwenUrfMf4Xjf8ASp96xEXHo6jC8MIN8MhTE7GmrNaHxbwF8
OHEMTgz4IrfH3e1RZLFJfya+m9p8MTjA8rHLG9C228ElDCL6jvVhN50ow/RYfmMc
hYpfkWLzClWAJ1s8+AdyT5eK+VfPiHkYAjDfpZo1mxAtfkBEra+lnb5NI2MpH3Ki
JJOGTa0ZmASTzh4dWZf75PCZk/raYt8zBGF2XelzX5a6lui7bTCKyMDzIGB+W/vc
t6HDDUr61rioSOwILRBnrHkhye0K1WHj4vsoVz4pteHSylKGWLhOkzW23kqfvexN
wscgTlrUCKIdHOBESBNi/zO+tY52ekeiBaWh+BcSkL94siD16zDBXMKKDGif49dh
Ztkv19Z/YI3gpHqzERs6T0rQsvNkq4vi8fJ72THiP2jEEXgZPW20Q6o7mJNdrw7L
uwPsm1bZmzYDg9BGodJ7XpCOSPNlUoJwdOFNtMNUzXAybyciteYebdOgiImjNkU+
SEaam+sEPPf4t9x0ZJJ6SJNTaNPInuTgfK3sWNPwPlypz1907E64a0ojPQUq2r0I
EaGATcDWWVDzD4diSUuI3nhHsuYxsH1pFWj0U/KvF1/Yb6nMgHVC3sM8t6IKY+nu
T9IYdK0uRWoihdKuTT38Q2dA3gElv5M0RLtQiJdwvw00B0NUiLvsRqucsyCyB/5q
6NSmWEGH5inE8EnQFfWAMNxDvwx0qg0DXJhBNC/Pnog1VpZZmmEM7O3WOURoV2ec
n05168lKJBuIIQTesDmfUdOFjfSkczruLqvDVvbJwFBoJAfF5JawHjvXZbDD7sop
opDp0wJQB1j2JGOtzAjXFa3BGN+/RgOWa2Cjyga5dZgwlswP2lX4Xf959iCeE/1y
vXavTBiF54mcEUOi5awUUN+NIqFRSDDcfM13vIaJtYNLX+GrQHzPuFSCGqO6MwZK
AGsKnAoNoVS4OKCF4V4FtdEgUI1lqVro6UhGb6C+ZlshELjXz7RpWRB/i2OoPVPr
PNBMj9NSzZIEPwFmmgo97JIAkKocUAJnXysIO0ko9B7RtPKRaM2cZdnaGWl4ott9
GWPG7hWncxmRcE+Tslr7YrfrCvWeIT8zR3pvrMzyvZ7MrMHe3MKofYfl/2fbwisF
B46O3Ua/ygrXXhOh+blzLkoEqcsv8/2XiDuhR/aWboxt8VDo0sVMW5BG1K+JOCe6
yFfgqWp3t5SycsS0+QAMTTQNp2raVO4QEeyMXuoeaobkrSxA48ILvVLQt2pN8YYU
oMNKTIucYb/5sKGD9HbDklN47ZjMuJWIhvyEPvxZRiAno//Guax3KlM7KUfllZOd
W7FnnPQ1jbH8zZQjPYnTXneYQv/HRTOY3gJI/eaSJ2wS/cbHJnzD/tvXMuXfV63s
wWT8Slxk9xgoQIWCdv71PMm+0LwsWeZVkeFSeTnmNzvXFNbFMgWw/WjXWBxLC9hD
+nxWG7W74V/JYKhRC/4F6EMdSbox/Nsdo7K8W1JcJbx6NE6t7SvarXbz6qVer850
ZS6ESRGM1B5lqo0NzAsON1p8g98A/TeC+oAvSUWQppARG5OpICdiT56tthptLp/K
PG0QV51Js/0pPS4gvJoXk3o+B63WS37rtDuFn7VqL5F7NWrzFjEoNpRfGZv/yS9Q
cao9h0qNaUTXGQR+7spCWJ3sKL6tipEvS4Yrcj042mWHVBfGaTEY6k8+CBfLhb/T
f8rXwCCBDSAYj++UVWL61IYaIJKgJmaoejPhYP0+1dt1Smu+R9Wlorfh/ELmqBWm
eRZbvv6ztDlMxKTm5fDkHr00pGoVoTCqGJRUtkY2EeCiOc2fMB7EXJYvA1O5eHaE
JzH0Lsl4OlnMeDlP0rtICcCWf6dDj73098YZL2nMXG5axqACu0xtfyc3oQiFTO4H
vuix7wRy9eu8dEL9weAnuDVRFf1AXg8LqEzDlsngU5/hKIMW9wdQQPugdQcarZnz
PGsoBQI/ntx/mV1qrRi+2S1mTGQuoH85VAPAt9ymEuG1slWYxa0LbiGU7YFMvdoM
w9r6JkUkHocqO0i2NdEntHYKWH1dace6xer42fzD9DycJjuKi4Ggk/IAKTEq99T4
/km2sXar3hOUWiImmlkmx+QLMfElLq9cTTb47ztxsOmrLGvA2xrR8wC/laX/V8qx
xu8Xi8skzxopPJyM3Ka8bALxqoKMXdMVsQV5fxNPcLb+dWBgYrlZEFX6ViLcnP5b
8XlELqgAoyqb/thYS4VDX8CsDFD21Wvf04mppFdgPWSwHINd6lxSvspQ5AwS94Yz
QDtXTzZ/RhUQBWn6XGd6qURR/z94fHczFJmaERv8c9s2mc60mT0NgcsvvJsee/iG
jICCgwbUSJ8a8Nr0ouxVQmhvESfYwTxauh+s3yJpCOlCB+JYv4ARHBMKLCJC5H3G
emoZttnltTRPE/qB5b0zlGsJ21aN8cVaPAiAuLaUD98xNXC7b6hOVvgW4O7mfdsN
MZqmlrT86qHlXZUZT3oIFL8DoCm5+9NpKtOwY5QFqfq8GVzgj5SNQNytFdmIUUsx
2r3P4bbsjG6qTeegHx1kFvH+dUqSFG+pKUcn01w2O473COUMxlquRI61R5gNceHe
8R89bUkl80PTpFtkeK5wLwsz95ydRecmReYo7qWEzbx3q2fs/XEX9nksQXQ1wPzF
gqBFGFPfKwzLLcKVDMbTFjL+9iMXbmyJ4n8zXcdnhKcGniCGKxTcdHPkSuCtIT83
V+nQOJx0T7wfX4Xaw6ErCJOYSPAejBv9iopQWKHzQOaiq0XXTCU3I23lv+f4FBMD
txj7OQRW8xrjqJq1ZYG2doIY4Ke5utXZ1km8sw32UGzMu1qLMPhq4sn1P/8cK0dq
WJLW+wLIJ2kJphIm5CU2r+bT+LxtX1pAuwTKim3yIyGobWjj/peyrsl34uNyIlHl
/ZN8covWuPetHyOw1p7TFBuWwDpjSMlV4F+Q26KSEy1iam3APujnNbVvf9V72QMn
kHoCa1TEyEXKm2bH9ZTyHuvnXynqWK3XhvO3VLTOKPG+GjbgewP98SNaKxzfhRhj
myY5CX7TKt1UGHu5KV/lwzbEf0EUAJhZO91YRkhWjRkLhUzUw6JtTUkS5rtFpjWx
EXxdsSdylC46XQj4YAriklUaB7QUUB/YhtcXBtstER7WmxoxFmkzEzvw9DnlCgjF
6jA2hP+b6OIJnP1HmiXK27U/nMmdLvol9hTMiOtUveIWK8s9vSF7j2tnupWEpr7g
cgo/payKVbZHGy3AH03uSUujLXqonKP9fGo2ysmOvKkFCkHz7vMEMFEP7L5Oh1lk
avqItaD42IWmPVKaaucmLdZ9IYYUDklLMQXjnkV/Hx07RAZCTvv76v10LCUJGZW/
yNZopT0FBik6Di8rogoYtVKYvD38T5wIn1TxqR24NmV4UOgaZD6spoqNZ3McQWFn
3xhIVAZwaKmK3k3XRnrmjD9vldhTBrn3be1O+KdOCCbRkeirdGuxwKqWiWvkn+0t
MCSyp1yfjDvGfelP9WXYrixT4GHb7jvfgv3qXkY+IHqVxD/pFClW8zzh6nCWtBTJ
vNNG+/sx2E4ZjiPIgGKNSofODaUSdd+yBwgPSg0IAddRP7dlXGCQ8w6Qj6yLDUV+
XykUpORrVlimj/W0ExglksMq87qTnjkjSouQg/P09mrzh4Op3DHi8piLDlV2zXIm
rmtHyHFC/pYhN0/jD7tXs0nmygI5JPp6QD3HuS0dKd7ugu2d7N/slG5h1+of0Mpz
lk+pShDmOt9VFDLQ8CT0VxMfef1zX4bLBVsIQNmaVYB7R8gdMoUf4ubEVcqNuZ6W
3pgSy305Zp1MpTiI5I5mRUBlGJHSUuLFT74UtKvy1Q5LjUeqDJRPdAVFhzl7sQHQ
R+uWY6s/Jd0c5LpLpdMgbwDVb9tDQZecEOR0YOjmYS0WJBrXu4pdySBf1xG8GyH5
/SUaZ7a9CWioIX04yvrFvMIo4OyN9Z29u6gr7goOkEb8X8Y0ObDxBWfmKgcFX21k
E3YOHtI2Dg3hbxAdP8MfQlhIBQYjrHATOdCZHfZXSl74qnrD22ODCpHOFDwrs2aJ
VMXM1ireOId+efwluC/mRnD9XK4vTDgtUZKpnINi8V7Iga1W7VDxuj/h5lRvnIUD
esFX5Y25Rwx81xjDwieWEwoLlNhjD71rYMCyhPsbHR1O/U2TXL5rLR0z6C8/5EhR
FtFYusl3SYlQXMO9E1aM8RQfoJHWoOBmrYkhWgLLE8W1gaJEwg3kAN00qDuVeFMu
JaoSOV7pTdfQQjj4+h9aLUnxOHM2XJLSn0+nBXx9NqUCwUoOZ+xMqtOfu++UWCxR
ECfADP5flET3vLKU8eA1R5qBz4CEtsRk2r0mMjbpWGGZlrNL8oDhFPiT/LVTVb7O
+xR1vsaVxHe8f06vGN7KhanCqTtOTLa0+8UU/q8WCje4OpoOigGi+i5jL5lDe4l2
tLAp8QY9LL4yzHC4ELgqyQSLD+/1Wt8Pc+oupV8EbkUv7ZW0nTNQfd/QMdeWOJbB
Da6F0bOylUfvHvDfKGTxt673NiIR4viIWF9HFe4Hl0LALpG0XNdTUjYCf0ya/jfL
SLsTe9m3cvD87FBQEC3sKSFA0qRHdArVyhJB+Juco5bQ4wSPwgXw4GDXGUb2yaW3
Q4j7gFROUS+qIu7BQF+3K7ytCtfeb5/iHW69yFQcIAqH23c1XWeUr1jiocChuZ9p
S+a4RxnzS+IGbaiYqChgo+6snV+LQAFmImEZRpO06BMj8aC2mtfw1rLmnx/dRhld
wFIIcFQPC3xLA4EAQVy3bk6eqyZwIR6sA68AAzA2W89Yqp68AHr+Z6WLep6P18AR
A5tCgcF4MZ82TJwfWDT9zHB1CCUMQMriO0NmhUjgLcIK6qwj9qI0etyfkZ1BKweM
7N5Oav6BPy8PPpOcor3nPV6HPuRBud6DxcpD1j8k0g/uki2XX1vFg2LUDx6KtXDu
UkWioAt6b+LXp6evtcQSzAPxuOcUIY/laWhqMYw3X/RJFJ4Y4cFAQD8WLy8CHme0
cKD2jreQmpW3K4gXg/lb5dFsdh4G7e9ZHDA/ctUAjAxvxBh+YghLr6VfxSLVGgj1
jv33j+VMBUvD8gEQJNfsT1sQylGLiOh75r0fcgWOWVHQu2MK62RLj+0T9EUHuoPN
8bHFDmXyL+TnqsnbX2cAWQj4NsQs9cmBxxEw/omrog6n8p/HUChnAwGaGC+luCZz
nk15r1DSGv4ar7FXWQ2e31X0e98tv7DAHgI7NrTeCQqrPke2MdQ/UscYEctzOhqu
dGQMNrVDzK7DmjwK6SEpKvDPZbqJTMSEDGQprb+AeXGW6NqL9wVEQQ0Yq95sPd/g
ofyjK3Eo0duDq17NrFOg6smJfYQ/vMRdUvWIcaSjOQ5Iynfed1Y28CjvnYqtKZGR
Gi8p30rjCSPvRdkh6ZMvsjE1Dd3F5FT/OXSK4zaoHWpPvD7ZdAM0akDxa3VJ3hdU
e9Lo9RKS/v6hFoAlMo7e0W2JiHF2GdDnkOaSlfvQvRScz0cm5+hE+fsLommAGWHr
I6eVvhHFIyXCDWVa6RRPd09m2nm8xl21+S/8AxDTfO26p2v/9TtOh7HmuIfSh+7J
dy1rEeEqvniaY2QenAysRWO6f/xlYySfqA2eyRSLHefjVvA0QGxtv8leAS0zElOv
xGm5Lw9BIAwvF7phgC0DtIEZ5NskoyC+048ijC3puTUqYBdrOeLSvhDInwrVtMen
rKkpR/T+WOoAxBPMU76FdvpC7SnaZsmi5qN0YnF8mrZ3E2dQ340N7sy7lUzofe+l
6LTtYrdeaRDxGDAxSkTACBudnn5/cdgo0shMvFQAhGnNwNVlB1X3QJYQnfSWCIMk
UR6e+hhw+BynhJLpBouhVbeWiOJA+me7DxRLUavNSL34XaUHF74EHNqD3fqQlVeI
gfaFxYCp9Wnlmm7wu5jJxMZY5zC0kqRs2ixXXPOyPSgtDgcPMrosg3N/mR1u2bnL
NTtZOnyk+OQ3DkkBdJF+OhtrFDwmzNtI7ZlHhlkRkraPFnG2uBzpajcU4aKxkXHI
6gc7JA0UwDgYJ6Q5S4BznB9zclcwpofajAdDS0NwupEkgq/jmHEYU7gsLxxuZW+R
vCp2nSTPlq/bX/CV5aUTvNHT4AbpC4Cy+HGRDF+Rhlo0x4O+V3w41dLcKsfbJf7h
Lr6GIkzTwJwOB8A8tL0dd1SJ8CILwOsPXdSGWEGRLTVtHCdXmGejXz+YYK5PwQVW
gmpa1PKK6l6BRUcRn4ZqewNMcLm5SOFDrRe4kSH29eMDDxvErbuI+y8Z+MS1Y0t2
y/xDdKufZ3DJQXBDDlvAgKBR+0yRmbp9/ev5h/R0AOY7OR0tQbSoWvglAxueLStT
weCG1MshFtxsg26FNOKt2r1E1raj8T/SPz9E3H2+uXoW2EU90BkjMcMukkA7ICdz
ZltsFSj8l9FT/Hbj1t/G00kuC/Y3y74PqbMfn2AP1rlaphBklBFGD9hAluBGjxd8
1HwAJdze/OHZTjwi8Svfi4XkIeOLpFxTCHEGJk7BJ2K89xB4WB6h/sLP4UHahLbp
mQM7VNN8teCME/+4NsUtLD88Cl6mOf5EhIC/A8dTC/eR62STWoi19eFJ3DpUYZhD
XUBvvcCd7J0mknZRyT8cqnW45MoPTxMpxNV01w2KFsPOzACr1WV9PqEOxX6lk/F1
qZHIDFh2jnuXa85JWGeEL0y3eynV0TB/I9nvVhMUIbSVJRI1vwwnPJ0PNIZK0Fob
QyZhV0RJO7n9aNk0JUZLsvbmh59WrvbOHB8lIiUy15uHj+IdrDQlOj4zKTiejtVd
KkUL9IBUlKwvUv0zV+w6oGy25xkqmDE1DKa53GuAx9Gtt/onP+XIMFL6Lj/P8wCZ
WOyh1Nv+mWd6HsnprzMyLNtOpvlC7UH0NmnEIDqn/urZ7fGrua7L35nKStpNT8SX
ArN+NKlaNHkuoaj5lc7WZkGWlojPevLjaLCCPqI+CUYFHpDrf0i2HW8d9LmzLsTZ
uGl1UGoXXKVOumdJsxtskX/1Bh8K1jdF69Pnzvpg5NLyX94rRrFP+00rmJ29uBdf
oxKKfhH+4Dl3bqc5aG5CSsShf9aTw5zhAkTZJhbW+UOT/g++EAI0jLdDz3AY5UMJ
0tL09XWgEVTBuehD+gy82xhv1oFsAwsE09OJ13V4ayG61161r45C7J0M7Kbaqfx0
cVBGb6secLZW3oPvfVmzzyrNAlOQQc4mwgKXWqPRetgIVEH/Sh8cmPMqk8/f1k9b
itqNcLTwSZjY+k7DsR7fzB50A/pvw+SM+eMBIOplGSKxo4lQWBJQnJJfCpP+s65K
qW1rwaeTnHVdk/OXw3Pe+1lZaAUYy/nBzWyMMYQSmRIzN1e11zduSF3/jiBcTSpn
ImwPjcEyFHUOvLvvdT0Jsah5Rt52YDEiNdSNkoSUxHjkAVuRWjcFW9UIIh6/8LQU
KOo/1TulWgN30qE8DzNUA+6lUNu8jQlQ8YKQsg7yX0v8ZnUcwefye3noPrRAYRxg
32Kzv02AyKHittCnUA6uaKJd5vY+MWtzd44H8I7YxqEGAsjX93M2DBMzW7tiDJru
ob4SGX5FeWiO+GVgxBbn4ELY+1aKjo3b2QjLov8/lzWtVccbx3fCaveaGa43Ay8l
AoGycoF+AzbqZ3JF4HFJiagaJJvYKsQdbB+i5g+h5jwKJKC36JulCtn1ke5pFkDK
D83Kjjp7H6SWEYdieWXA3XpUd2VMHrUTU2FJoaeYpij8iSOIE9i0cWHi0TVQtqjv
QsAqWp33MAuVcwlNXPX8RJSSHkku5I+3AF8fySnScAFY05m5EbutN3zI1Qpej1LR
njukdyZeMqds5dA69VHCBfuP/Onfl52GpVKvgtWpe+mrdFiO6xfKoQ/tKkni8tkk
JYZ5n9B/H4FqsUSSulNT8qQmYRc9roxdzy0IbbSAXrgsLHFk/qhuj+2FPv2LPtl0
5UPLwUln08wGruoOZeR6+NixFsFscCvzD3tOQTEKJnT8ZF+PI6Vijpbpja3ExNuH
LYSUYOHbfrp8As7pHHe3dEfcV7nRz98o8QiCoAGO5+0a6MTZY1pPlYQIE3CIDeLx
hBeWHKMQmjUO0f64t+e9s4o5U11jkjGBN5qR6J9V9kbBE3syRm4RoCH9o+Ha8Map
G2/abyT9jeBq1CZbTXq2iXeuqrzSLvBT079zs5dEcMafZOSaSwmiDlCrXxwVh8tL
NN4720LD9zGwHkPv0bcaDD75NYwws8CugUuEjmJbKegm3FXj/y7Pih4jQsGK/KV1
kSct0QqS+5BRHcPpDFZPa9k05c+GmiFEXSHeSLh+iVlza1dEBeKmF8B9TeXGakA8
S/Othc9YS6YIURkgHDs+3mMy76yGjg7/bak48elcU46AFLLekMBNCzaIIcpzd34H
AejVlL5XuXXG5mLdx2Rn2MBSIHwm8MG092CvR8f8wvS9qOZCYOmMR/Pj3//jYWAm
TeKfvstWPBoknIXdtDTutodgVw8rBr2EQ1YKYB7Gb/tyrMum9UhsKJFTSCNZirm9
JZlqHJhL8a7VBWHwPp0DKNZQ++POCkg66uOYT9MND199l82HXjqfVFM4ZaTKEppU
VvGO5A0EsukLw7qJybqcw0uVkDHCHMWRBgLJfAISDx9HFz0+MxWl280gXc9E/kB0
otBMey1yBN7PftGFHY3HEBL/dLySsG/4hfDZ3nHNxBXZ2lECbz5X6W+zbcAQDoRH
Wwl/tnPmnt2VfozM1Al/uPqh/pNzfWqK82jOD3WEiZN6u9GWa7m4OlMFWrV8c98W
jNXlC5XdJlMKFydOky3rVm+Nvb3R4y/6TaAcVso8VocB3FLYrTP19yqAFS8dj637
mbLol8/Ee7g+/ist3/7tGtIbYNoQDAudb/HF7CYflRHsVp7tLlxC+nG705jvRexC
pOXvDU05ozTC32b4UIP5BPM5nNNOwlpBcy16a1vUge+I1L4PiLec3X27KG/qb7y3
JvQQVp8ENCUpM+Yoq25GChaeArgF605fxg0pPBAOiwUcaGZu9Sg57rVlV79lt0gx
WrU+SdPZZUY4iHXjiB6xr/9G5VUylzmYBV3mVtcp3K332K5KLWXdinkoeL2RcU1d
+ePEFv724bTSCrG3X49RUnE1m5GPgDKHPQTQZh9AFmutlb8HVVSB72KqwseVQ9q0
NlVXdJSVbMJwvCarjEV84KagE6TtqQ4UxPO1jbZr8EYmn/rA4kURdjLeGDTrQCol
W0GouxQi56GpuCy6X/n/WLUrIJfAHjNMAFiX7tLIXNTQm77AmY75rKN7WPuGmbqE
xNGCicrNQtl+7k/ePDG223HgvTzrHr5sQrv5NPjkcIWQlQ9AT/QS2rL91ILTo5QG
AgY/DtebgtJC8ZK/z/jxCkhnKveyr0NU3zBu9u0rShR1G9aTPSWC4MOcHcjq/oYq
84BgXNGZRoW8eL27wZvkpjIjgnUuyRLCs7BHjb7kEoNLye+T5ndnPVRm8boL3+Ns
cZquITDb5EWCFki/m3zXmbfbdSDQ4I1wonwPf+515Z2i59nmU+VsU3k8v0MEh+fQ
ZrR2IE8qDZLq8gY1rhsSXN5BSUPpXfePKacEnqgxiQ9os8yqL9kZyAxQO0j2quG3
S3rnqXM4ALKIsOj1fpcND2ammDVHkRD5jjFouuYHQsiGbX/C0iDrop15IRgfLykh
LKpI0MknhO2J4/peQVUQXTfAoAIRvDeCSPykMDG3VAciw3bFhivHhqXk6Wistn5p
EprgFSWbiCvRmOh0cN+KloBwLhISWVX5fUtQrLXSWn+dzoNdLLLZ4tbkoceYYBad
OMWNhgvjr4J5bbEKGYVrGyqo0xXZ8JpaHv2D3EZ+ezbXuh7eiG2gbfRDJKTQ8OcQ
h8bOvKYG8cVT5Yo+Qmqzufuub5eX3w5hscs+OVnWN/lSkb8E7eITccuYqNUIPuOH
D1B1llElq2I+Zg1bdhvVM1Vm4DsBjm5n2NMlvMz0oY7Lpsu0kJR7mzIgygTKCbCH
l7jfxCMaVh/7BwUVzBmM+qX/b8SlChRRfZikTDL1NtFkv6197shgjcJ6s7v/BJSw
EA6Cv17G9H/AlrbkeedjbdaxKoLwF+mmr8/qRzIxVX+VPgneBhOlcd4F/E3I5h5n
vkTpRFNqIqvk8enKU1FcLvisEvojC5w1Y84jZ+f6TCWCE00cVWIkLRZ3Czj1Y7Ma
om3tFtkL7wOFmdHJRW5VCtSCsnfSQv0PJ0g8azmy7pu5JpvWxqBcgBznUufKbYQo
T7KdbD/IbCdgWNYiTmBDmns3zb/4vmJlBkMo22FDfAdOd+QNXmZAnNMFNUWsm9EN
UHbY+LCbd1Q0wtWubg1YzLo+ibY+7ip24J5/ZHR2ZIvuomM4BEQ6vo84DMj/RdCk
XCnyt9GYIqDOxPvZYtz7g8oIOgVhk/Gk8dlhZEIRfCayz7BV5IdgMld1ptb4UVCO
W96lHq8wL4rhTaWN80VzFD8kmiDTZFOkmdZpy9CbN2/BCJGHJYj2PwHlXCNsrx4t
jUo0h5EeIdT2tIKbX6DNQp5yqpopnGqlZV1C0z2smXZs0iNkGNLUi8xqm+bWeCH3
G7X9QrL6sKt//Sjqunxik+eoMYuejD0vYoytB39q2P9KnEBXQrREctJICyG1nlPy
/YqwFvpXzA9fQRDvlbqy/wSpJdqWHz2A6qp6S64S2y0gfB2AbBy39f8xlSqrzwDV
svFt/u60u0Xj6CnZxJlc0P4vb1bI5p+8NrY9j8cBR4wgBu4PoV/0FUEwkabH+cES
V/xEx19aGAKxGTS7aD3qFHOjAK4M00vrRJWkMNcTXYLweJ1JGVcUG4IF1xfyVTmV
cnqe8k/c2njJw5p2CcAJ62yZx17P71EyW/aFShK3UdUKzfRyhshW4zzySRU92xhm
V11dL2xo3PnTQ3UDZgBeuayHWtp78HkRxybg0esV6X7eJQropxOPzN5pYaArj2TX
J7IIXm3KiaZL9zVP1XQ6yyUTiUW+Tii6vBfw3wb1hMjhLPJ2+bQzRbgLxG3QP1+L
rDos9aNwgC3kgtU1xhI1zbxdPSOBHt2Y26AQwQyP1pxQKFXy9jdMU4/0SlIO5nRV
lPiHUj+0n/qH40X93eXMQV8e98letmcWotE0icLdWxqj06PmFWCzPpy7XcZQ+KnC
nJweZqrjM+dUUTKv18qSCuWncofjfijtlr8R4MKVTAbFJfOWpWc2MXTlsKZ5cncx
WTfcmnxDoVuWaMzkBx6mwrKAYQKSlo2F5xpbvr0BcRoI6q+TEvbczjBeWRkVB9G+
C+D0k6MasYE7+sWl/uc6pRcocqu9TPtqP8eqxpkf5tONBJ3WbswFsYF2ObqLQWxT
t+506fkdOPiQoXWMBf1GTrgsUXEA8YmbJjdiTJCrlRfLy4QhhZMgwx927IsMsjEE
whEk7B4L6+YhzaxXnh66pDdsYSKp+u1xGffhgYIsqTrWiwkbBNyH5q++qnVmZMw6
BRElYMZKGWyN10v9Vv/BJEQCbzkSC09RWoyxD5aMshWEg+sCGBtCxp09Z+2e0npc
AWQ+G37K4SX9fmMCBh9c06SIl/TwsvuWjVeVe1jyrBihVzARpxK2zv5XixK+bXq8
o93AR29CvDkrjA9da8yEfZdZEcFbLJ2oOBdpG0nHa39eXqK6AC1KPZZ2eBv4dzzo
6TXTNXqjgQi/UBCx2P582XNSWgaSNbEgG/BB8D39xr5WutxxZkKlSIXTXZTRV84c
BaF2ep4In67elmr3bmjxMTy08Cd68EIzTiJ9qpwf0yGprY3Hes14KOU1kiuqj2ar
Acya1IR7ckzY8f+iR9oLg60Jn5TJ48g+FFxidyjiLsMK1Gx19YZrCGGaDEi812ss
AcqMHfgir1HqIy19bv0He3wd1Ic3esJYMfZEckrey5/R2sUFTGOlyKacfg9flK4H
afkLZy8fbIJJwLbJ1/6SrBbq5wjm7r/Yg5BYg6E4LXVov0zFheYcwRU/9wjawKyn
a5H6In2NEmqHnAORUECjsq0fOhxVRPiEFPoU1Gamreg/9fDPnqo93HW/GdfJ0ziP
G1mokC8HlOWPgjxmuvLKILChfWPZ1TXdbjALYujGRYcxK7kmtNJn+Bpu+Sw3CNKL
3I/AztcDDHD0OLNBUCywMYAGTBeNanEMcX90mMCPc9VBnzqqjPmyfkA2Ie8RwvD+
uzyOFtt/eUjoF3kdRmeO645HdAYZGkg/OTDZ3Zz+xbHj1u8pyAyFPHva97v3dbub
i9apqh1hw4qcx+EFjmxZDOvJy5CQy7dzkp01PuUntnDS4B28/ohMJCg9YIgEzKrY
krptfCu1t2qDJCAkhb3dLHwpl9cUL1DRtgxzMuAxvAGMFez1XO6dvwU7UrgCjH+J
Cr+fZWU/6cMenKDuJhh5vp98pUVC4Eead158/OjvN4Y+LCVWGv8sIl3B/YY8qjOi
SPOS3X3PV5IMeULNX7KRZfZIRHRnQTrXkTl/aLhdsLno+dR44puTUzPvkvW/T6GV
wRjf6F/7Ze0p3a+EaCtAgOrR7FI+KJ9/5X2+K/iUBiqz955m/jUlEd6dk3E2dBB+
fkgkgE+5lZ7h+bBtEDZJJeluRuiz6Sps7muFa+xfAwR0deQSR1snfpM6K4lsSSqD
rIeYeMnxLw7NXJZFPHzYQ2sS+M6UhV0Ea3FacOfddtvfC+E/koz/KOQekcLDbMW2
Ohuc/2gSndzCc36LrkFzO/J1X7GKPuFkxh+mnxVHZ3WrlqxWBIJ9kfI0tG+45FhR
ADWopvRqw8kwIzqaJV8UTRniktB3eLactjs9h28c2SguTIb0uT4NghiLoAeL7L/q
KDtGc52Fw8eiL07tqRS8wY4ZuA9Mo6jMusDgOwg6+DRfaOd6pbHLPx8mv+74/hfx
vkXA2ho7T1bCicv03m93NzbxeVgBD9j9SenyNNoR6nEH8miL53B2CGLWpTJKzr06
V6t3+CvM6XazT2T162n5wvDG0D0X2lyS+Vw7L7848JU0dN4+XiCR0eAKMbfDV+bk
goDe6Uqns9Eyd3uTLNssWSxFLF+mQIF+RFOQw3/7T96XvD33vIhCpl5/GNdaqt3a
vNNdglcO96WO5eOIaeWNAEpyxkT/A9UipB4mV7SrdtL4ZuZqxBuCMsaPT+4Xn0N+
bTqzjIR1+PH0lXLyueH04E/Rm3VK2NkLPnGeWtKS1MdT5hR9Mw8777DyV3ICGksY
m/x8m7nw6wNgNyB3/69LEIDjFTALAVxdgDPqadNO0ycQhnGqxLnvkKfDs2ZCvW8k
br6eTfbKhla1FGTrI1QAU2Yeoxfl+Vr3cqgXrdQS85aVqckgIrl4NX26NoTvbKSH
9ZJVa5QEWsrv2Mdn9iw1/925XlT1TkGD0pm4EA9ZC1AHku7tj0rVRtsh/WZHjjK9
CcB893PY4V8lQsV5Wx7w5J+pSaLQgBhPyylH2gZqC0OCtBH4ulXPeT+F8aCKFUIq
Bc1s/U1G3sIMPT0Sa1dMn0v43wIfIoeFbnGoYkKP87xDft3hVfkAEJOYEcYPNGf1
d/GtUeLB3X3vKBomD4eOYBWVILfarKdPeuypYOYf0pLioHYaQiS3eWldg1oLRPkC
2v6CPjfOXzDVznKpK6j/YWisj19JLqfXHmic/DjUsjVxsL5UO2vsBuruF9dv/H0y
R2PnFukli9mox78Mm36gLSQnyvAHKVpE+nQLBM2h44VOfWUaOHscg2heZUmp+D3/
63q1GrJL6VfocuHKg7Fzja0JAI4OxAcXKHSuwpJbgl3EwUkf0tjdR/BSR+cF7Bb0
J7sMYWMShOQf1Gde8ztY9TFL3jHU+epvigz4TQvhQMZ6cbdJhrhTkWEtqAW86dUy
ZlYDVluvrUv+KnXhBo8THpwu/FfL0V3yUVVEb/fOKo0s04kFgRG7u+ebQrJnOqbx
ainEu4UIrD02ZEOR637ET6sNDGGBdlYD8f2RxLu1D5i4qc0As08VD+YAA0RVzp7L
UQAXW1F2yWZY77BgS3pUuO018M17lG7GIVpcQNNb38nFbQwMo1KjZhQOtKgRbs+T
s00GLNBgrddhPGSSXvhd1z86SojoC8v6z2tberTCJbuW1OCOFgMfu9iZxVC9e3Sh
mcG4qLC39xlS4+11wRyQA4XmyUjbKX9+QQI03FiuVB9Tfvph68YT7DjC3H9BALFZ
sL84qSmMbjGy92BvENzDFeXBAS09rszgEylsUIviOZFrcwFCT1ukAeQSTgmcqv5c
0/g1P89YiTIPT3r9WS/taEbENGL74T0cYtt0oqGflc/T4Y5n2RNFXBDhH82XThQW
3GhjwGKhkJcXa8Cfm6a71x04HHLA2Psb5rlxyDK2x2YmsX2k0y+0+1QyhEWaZLVT
kpTISkSv1iDYVP/FGSbQJ+6YxzXBIfULA02uERUh0OfUQsYCueYQW+xv90AHKlNL
Rv+BENA8S7LpaxAfg6aA3iQ+BpPb7zkLKAqXTqhM/4RSxcYs9yyzRdp+sFRSYzPo
3mq9Mx9p0UtUWH4CeQgBxDPsSaqZCTYTrFng8MPRm9MB3NCuRFYu2bUgEQYURo4L
y7XQh1wBBChHQRJFVeyXcBVrMUcZuqta1AE4mjlI/KwU3CT7sRWgCD2pi47NSWko
JvT4VvjWL6vqoIdOd7iwCMcP0cfFZP7mibvVbhISSjfcrza6rHR1ifHGkZt9AXsR
j0NHbJhux2UuauV6gu9mk8f4S3nxGTkSr+MBUgegF/2FgAjm1w4btncXE3siL5xd
JNDiEkKFanLQnTmb4n0hCfFFklxIOs7+SMCv8jVG1ZTv17MZjEAiOyfJNaFE7xfY
kiGlQg5dLIvE5tG2jdQ6H2rmufQTstSvZPJvXlmJow2POCkj08lxO0IakwOVwL0G
8Lrvti5GTkN7xBnGM1JqrNR9mfBiuPxFBjhtz5tSQjuVc3EOPKlGQGZaSM0+q2Rp
9i5LiHosUTolYDCSxmkwwMX/VSnWor0GzH07LFrRyHtw8oHuzi+GBcKB1pOcEWuC
jnU8uCBpQvuB/dnHzXl5Lmo44ux7axGn1bLqx1Dzj64=
`protect END_PROTECTED
