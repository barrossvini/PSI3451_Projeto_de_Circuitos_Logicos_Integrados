`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjsT+Glej/0/SMd7ve6SKnE1SMB4Krl5w72qxWTOyelENboQl0TIkyy5hUzf+onA
g60mqq8uYv5HDo3xplzXY2oRhX8MwPqr4p7f8wk4tW1DAIaSh2TbG943645XFh17
xxH7eipHMrJKUIuCSeVvoVdR5nBgX88BlW1iMDxISB4a0SPF7hN8B6QpJaxiSxMz
twLmwS8tiDqtHHPJN8LkMu9IsVHr70qNQjZeT7X3BViIlL1T899/kOsrXeSYYXKH
108O3yDrbyhJqmZN+OI5+YmPg/72d5SPgOc71/2v3cq/K4jE63vCcvvIlTraRH6r
DP2+XAoLNNFO5M4vuX9Wy8D0zuRp1XraXNSzc1zllcsKlqxnBtSSakEZgtBif2bw
qNRZ7qW+n0ZWAB0CdQw5UBrZlpUURbLkUrfHeV8K1ZrDvcAZLBWA+SxIOvtZNiRo
S/uynOnuTeFGDs2J2QzzBcrXktxwbDz+U+DvFdsDCdQZJs4+b1wXMTYzj4kgjOLy
TjlUFlqwVisXM+kgpR7yuWj/qZtYaVt88dYfoe6QlePVE8hdEhSmc5E2Yc8kBlBi
v4jk8pw0mk15iROCgr62Rf8aeznP29F457enrFId+2zr87jYfTqKbQMJCn1inhu8
i0iIEjs0j4x9776deTcfwsPowXCa/sPWhdfe5rInUrK5myg3KCFAtmsdmmiV5ZTr
9IJdtNVS2QIjs7AB3KN1MYTZZKox3u1r9RlfpMlTUhAtv3FJJt8OuZ3lsFwowRrt
3/2ZP+luumejKZdEAEg+M/QxE4itbtk2R/GJCfyeOmmoc2ip9Uh8d5HrOBTkadFX
swOweWEStqOzGIXfvWuQNsiTZNYEq/yF/RQAKUVjdR2Gq4Urp5exfTHstEhKyJ/Z
4HZ2HvRYXPtooWaNZ4RSp3mlIG1drwM3a0iCtPGjHEtnYJbZl5krbNosSQza8z4m
H7fP/V94fNraJzHP1VRDJ3Wb2kirbqqvzGqO08JgpQ4ktNqL38fF+8buPBu/z8N1
esR81qk78YKzw5kW65eM65AvJM7oko2cAqyFC6FLeY+kKmqHcTpXLnP+Q4MWupqL
xXrhBI9VXw+ZflCwa4fIkkG9pg58SpfPQxVm0riAdyEAn2657NeJLok4XfdCMHd/
pIUM7F951fQb7Q/hV+5baLHAVnm92STfGbgquERpK8BOPnK5xNmLzvlDR2oQnD8r
DfF6cYkGxuj5WtrKkI7OPXiO9xwXKTLUBecLnYpiXP4QyZp5krkxCCQPjiBu0WWC
Mo9NxRylG1CvRU1OrVv89dLA523NBZ2OGhwaqXqdp+XYQjbahDuqgU/OU3CHUBc5
kGIm7AKTDh12xHx9vwyA1HcJEQtbKcYGMQ6dOMYN+ae4iaxjLOfKsakMkZY3snKZ
zpKpi8K79+4BJOsykFcKreM6OQxu0jd/pvPE5VHNrygszUitbjQxvTVcj3ilkSvV
lLNwvHHN4z9/eY9cNN50zzXlgmwVroDpues0cE9ZKDxm9p4470/Y4uKD8JA7lz3e
el9Xq9uO7o28BeglqdeyFaJLG6IenVJ/uky1JflC/bvlKUMMEH3odF9jmQqnRhBn
OSC1lyLlMpgyun/M84gLBnVkXEtt4TYrOcQue7Pm5Z/RUm4OtUx65SsiGp+5/F+l
6klRvsTFYLjsCw7FR9bsV/eGcrmNgJySds+LULfuvVCN02WwpBqj9y+AScwtGzCL
d981ZCYASEg7/b6HaM5W2N4B0v747VCqouE0wNpxGMMg5AQtNHmYPYMuT9ow+0L6
HyFhW2TETbdKvwcsxy/HGFBtLmtk/hl+ofMoSttIpnQbfvOEu2ESLOvPxOk9PXRU
kQHAc+awlkJVrGu+nHnmr537Wra0K+2BdttjKNq70yPlniuY30ZnP5e7+sfLGN8h
YkCmY+vCPa2Elp1vdGjzcPuERJifPcI6gqJqoPERQ7rd8R4QrtYsoUkrU0V17Cpc
yvfuJW1dTQPS+hAoU9l0u1MKrlO6U13+pmjEwijPz76xSmjmKOC8wLwJcegmC42R
raFfqXV9nn+oKp+q4g3avwCpRgkxvxbpN1J+UQbDeWd87GYXla0l0gTYGE0t0AJT
c8DztdpvUSunnuDIbV/E2+Wb4V5aBXoPGLbZqdeYztkJrS7WH2yJGMtLEPxGlpJX
lgveYG3OiGeA4rZR1AV411nKhPdYIt9JiBzMhoKOor1RJPBAh8PwOB38EggoUHnX
62A9O0Iu8YWNJr6NqEbsgHu0i+VK1e1beUatiXQiqP9bSHSx8OWjiiQ6zDzlXfmO
GR8JCUDEE1XGdO5f406pF0zIme0gXyJoHlkg4L0y8wBWsBNRfUBlGDh4YkYEJiz1
EqcT1WhEuNy9H8eGl1suaw==
`protect END_PROTECTED
