`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NyNdQc8JYJPRepv4Ls6PkMi6dU/28dvEWXiIPVeSNbJMRSHuo2XoejgH0yE81ZLr
Hs1cMjIYFjFD/YQY9VCSRxoLO9ilhC8BOXuzS4I+4xxL0Sgm0qHRt/a3aY2p3gtT
VlNsUKH+tHp00isp5BBqZQxEC2u8dmgPiFKrr1lxtPnVq42Y8FKA+0LyzpZmYa1P
w9HeHnk+xx3Jxe2Fz+a1I1O1C0eei5e8wZCdzxCy8bFzf5kkT3Q9/4mcpkAtlS/2
lm56XVwfGB8Q3bhseQVDltgdOcjmVEKAE+8iyBV8F3zeyp3892KpTN4nsy7HxAJb
fZwSyR11Xc3qL3INWx595KnxpVRFSfqFSSpjoeJlY3GBC80HeBqo9KV1/Btv3Rcg
rkXs8IfORCw43uKHMB6snY0pQUbbWjhQHcMGZ1KvoMcRUeAE0iSVP7L71ss25Oo+
VHctCHexp07rvzPf4bOcH+cQtU4emADbhpeEOw+BiiFyx1bvvhL7Ed7PubaGAqIQ
QD7Wkx6Mi1nX8hSJ5Frdz5jOCiYsALtmGd5lsN0iEvyQrBfYR5clyphlnyk7kJxq
FaCHRVcKXoFytKTgtt22Ry/hfrAqhPj8Zli2bT2xtW5DosTKIGZyx1wY8wOg1Wud
jxjw2q92UdiSpBocZecHhR1zgzUnjWgERo83amiWYLnITSvmJOvF0xV7JrXK6mBP
hwwUSMD+CMkdYHcgLThA4RFkVvOO50jRq/L9w1oMbV3h/JfZqlF0E3HHnuD116H9
wwJTILNZPIR9zeNP/pTnjPRRygyOgKY6Jhq5k9O50p1nALIBPN99Gip8UOO58mzG
KEU/LbDUpHz5S5011GkCfZKZrnrkkS4Bu0ZR30lL7KTfCnEMX6JJAAuHL8VHrVW7
licd2blSgX0uyCPN6vmrU5lSmMTGCm1gRiw/4qgYUD2G9deCs4ajyMBxFOXvLrY2
Dz/1Rx/7NsFedEEYPZxXlYun6iiH99cgeg2KORKK6nxbmJKH8o3KRSnlk6OQR/Kn
FbN901vUXw1icmZs4mxm4YouomVg8XsQGIDLN2fzmUZCmlgZ6FXU90twLDWf+6oi
oSaCpJHSK+La4gObTm3qOsDBzroFczw5TVvWb37vhibHDAD01EiE6qi5Eb1xdv1I
wohP6Q1e/t47M+IyHhM8pZI+S/E/biXKemU2R56g00PV3AIeOT/RM1MaoytxQSR1
Igm6d9n2ZcCG4PGHxwRaVAK9cH3ePtxJtlabQxh30vAbO68aIwYrztbrqjZRmLRm
kErqXQ7RAiFceuTEId/dNRuyvtqkY4sGeY/vy0ShI1VxNoh/5+ANHw8LEsPwBDln
3j86hu8GPlqdfvP/zE04X43DIKWj94ZCfvoOkI3ulvhA/6+8ouskRXxD+Q5r2aUm
yfQTz4roHILw17m20jYkzBml/b1HQlShvKNTbaDL7sbYP5j1v+AtAGwL7wBb/K0Q
3Kh8gxbuy8rYf+5EG32Um7GjNSBpsBT69Eg/pGiU3beAiU+fbsaoT6yoyiq2IVPW
y58dHAPyIiEi1rUCgZ7Xej61eZW9ICifpy5p5dJe+Lx8c/BnLjkSh9NB02b2OvOO
NIBrbEnDRTRC2o/A/wlsbONhRGnHm9gI0hn29dVypqnhftSwSmnKmbtuF6bcOkyp
DeBQWYx8w1uEnRU6VqEdmEUS+zaNtX9ec3KPi08i0F0=
`protect END_PROTECTED
