`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZQ66fb9llLMiOIhpDluSmvcAjDbeswT2AOZVWUeM5I4VVfmH2tGwzAjYTbiRbka
9VcpWRmAOwy0tSkGgpGM/nro6GjtZDm+jWDZ4EBOh9M3IpMS989oCKB+iQGmcLJO
WOU3jFh98CpHtDPid8+79g9FA0CNAJ/vU9pNwWHmX7uYmP9qhJj0pR+0uBca6OMr
jLybVsrqWSqE/TZ3d+eLy0iunFNfBPvwOOT0Z4fu3LKyrSpGMVjakrk+QdztrMI2
WxOWTg74VkXcbi1OFYEfL62Si3UoYzs+akvwiYNYm1z30Cox6vW67lFSGG06g5a0
Z3vyH/gaPDUaRoPkIJ1NN90ysh0p97QAVOQZWQRu06B008z5AbMzrTsd6SF1epkE
6p/MC91hmVYwR8pvFUP3kejUwSKw2XMFOi7j0U2qoFhjMoFUhFDNuucrQ43emEmx
g7YZVhuuwzlrl1aR1K2yWH6DfHeVLNawSk5hDxqRl/ieNfW5oyCzf3tvXsMqarxm
Wtr4OZ1fOVnWJkuuncWGb7KznQxr7ioLMtPJ0vXaDCRK5uKeN31QlW5q0e31x80y
uN2RLUbNeB7vzH7xbWRsOmng/1rjeogw2dSV1fsU8+Ml18KpmbCUlDW8h02E6es9
pEn3h+F8OtUT0y4GIVRXkQvBNFOL+s+lFiA6TaOQvuy1bGS8pUhEk/sK/vaNf08S
rhNWdtr9pOFhvOT0CFZZJaBhdXdsELJM81qOetuPl46U5xAOmK2AIYJ7HTPlcHeN
WmTM74L6jNYf8VfpHJGNnqBeCtpSyxd4hm4TA6o+epFYwvk3nxnMTihT7VR64HsZ
43UAqt3rn55qSBg3ccvS/4QyvfkBy4iyQCdFBCYll/bp8yQlF9RmwsMO9B+drKOA
V3+HRsX7zX8WH+rODe+/W0YSHEowkWmzbnjEIhCCCr8pWIh0D/LdeFfHFPN/XIav
vyO/u016ROEhN4RpMNTDikut3mftRPPzrvkm36UgEpBlEfAGher+Ky2vVTE3oCBg
411c08mkrEbnDvn8QR0db1r/tA6SleNVFesI4TUsrjdRD6VIM/9IEQh7PG2dnFs+
5Tt+Q3ISo3T6lca7zgu0RJn2XK1xPy6k9tCzPcG/6DQEOjeIwK1qfIufN+TQ3Izb
WlI4f62Mh12HSrJUimQDdGKKOlDNCBVaSY+Sgd+pYPlOEkGCWPy4DwNbaJUj4DFh
74gIqRfiyzfoKakoVUdf7ZXA/Nqr0rAp+DMw+WIV8xjHT+S1JXeny410GgwBt2uT
bOEnGpSzyt59vHhKw6GQLBpwV6JFqPqmp2XufAxzKKactLFuRZx3TOGs8pT9z1cE
3l+rM+9+MAKAJsZAOb7/Jr3sBjLJzjO01d7ZyDozDiISRu58zjachGKckNtr8ET9
yUDOsmsQlYYkt71Dp+cgmqAowgyR/O7lu1oOWj8+lxP6stBDEpL3SGEadDzAzKjd
m9/LepHiWFV6RDprwl5VpyhfsnAJkt3kIUjHELdoZAuh0FOjAab03xpI1Sy1e+lD
j1j+0yRFPhB7Gx/oUBtU8O/kVl0FHAgp55HjnQj4F0E12bh0GqyMfVwmNVcytQeP
ZJHpHph03sW/QOrsaFlwNMqG7BSTVs/GNQLiKHl8EGDfHBkx0bczR6HnjlRFUq5U
BlXrR2upfxybbRccyhkFQX8IBeJ/PuBLl7Hnty/edLvkoHVRKoJVvhF/8rdi2U37
TFbiKcjCE5CoY//5OoXAgpRVBSGTnjEzaoK75LlKfCpPhEyPgXaMRgoL/qZlMmLM
pYqWo25StzO5A3PfVzzx62rYIGiNwX2X8ISgOTaZrCiUit1PKd33r8Opl/qGQl9j
7j0UwP6+wumshCa6v03+lzQ9JfLFfduGCnMX8lo6pSVTdxTWw6SIOy15q/wM66e4
is+a/SwK64zc23qqUmVyRhCJbAuMrqFnYLlbCrq01h10vmpSCl+Sewp6CN/daHj+
trIH5t+F84GQvQb6QJ7uTL7bpi9iXixJAiqy75RcsWJ9rLqsgMIbZ/6aoUq1ErUj
MLMU8/e223tdp1X1MPS45WQy2rSzUfoMhAdqqDEtk7JnmZZoXbI1OLUwdcxVskKS
qh/mJmK6mH6oKbZhGKGJ9rTzuHCSnCeYo49DtVA9OjYrk7hvimbw5VwJT0vL+NMy
9AiXrGunQPcJfC5HxHIiGEwkpm9v269YUQPoojoLgF6vB0ksQ6BD30JDfEZFZD8a
e3YgQYxdCId+f4uJjMvhduCX31SA08J2T/ygHP48UmZ7eyYaqIKrl+Ee+jtOSci9
2vUDY/IWtRj27gZpxkvWz/6WoqVs/LcqZHe2KMYmuO4rZLCjldDxCRI1dhs5r8x3
x/h6+sfZWsCNmOnDln+kHoZnkKY7vAUb1mGesDrfFDAOA2mFg76R81/WEsyp14vu
zbkfd/HoOJdGVJE0EjBXC+mbNCpwo6M/dWRPzFb2ZWgRiYZ+s5DPj5misB6bJbN0
siz2DFmppl6j5rF3AUyTQkdb70f4L+zg5wvWDvWrJkFHO6mnntyvnrff6k1rmcKq
uy/2/YsqvDqfhN9NG/u7eebeuDWw+klVE3GjcOdGRjkUWW+2b5mpl90cxd/qTfHJ
vbYbH1AYwSyfkvmXrkD6/JsnIbnJrypsf5jlIyKwD6rJSui2b5y+gRJBEG7tBTby
5HazWYBQ3zWFqr2hTkIcZRgDwcF4dvh5bA5QUxTEPuA2KbDLwNvyF4Ma55Hefn2H
jzt0B5kNGsjFhKkQBMlVrek0OzLazc/NgO3LsSveHkHiR3yy3hIPXFzj6mP5s2Xm
6X3npP/DqvUlrsKirh3x1qhlX7XdlbdMTY7PgNjr23xWXz72la9QR/lk8+S9B71P
05ugQMJIPnkLhJoqP4euxJOzOIzpfr3Aoj9T6Xe4TIEalT/cFpdP7fte3FjlRmwd
vwhZ+7MMVnOxWELgLWI7OCZiFhSR4vWByW4+CQqh/qsLE6JqfVR3ssX4YR+I0D7+
WBzRyxOFKnL40lvGrYgRrGBeIekVHcQIpaqoFPNCN4lznpwgIXFCYzIMS5whhnpw
ahlN0N2+P3JZhZrBUffeE1H6OZVTs7U3CaGrJR/IXbRUwUt37dxhVW0a859QcQff
ENS96gKkj/eW7lfr2ClEJ6Lbh06C42TQlm/yBy7x76/r2GHwJRShXk41v6QiR/8Q
6Am/CCLYp37AKopSHEeStollJN/I46TQpIY2f3JcSJ1nawe2cIJB+D47bhFu2h6O
ENtfjZ62v39IgbTKWUyM5vX95U3yujp1emi4IvJ7NQGzirbAqRgvqqcT0bVHxLNI
yy+WPPfOHNRMDwkqN0DRIf1/b5q3H9zwWbY0c6fgkHFFam5Vu7xAcV1Sc4vNdEkM
fB2Do9RFotUXsM1huJlIVa2AkTku+sx0qUOilXFGQ1zv0cYsY5gPzBwUYIfB98Cg
gmR2c71NWIZwoYSOHxNrN0KH0SE13wYCdPJ9P/sFa8VsdgbKZQcCnDW66JL2L11+
JR4BvRrLcFSGvKQlFqxu5Q0+s9pP+p/sEWAL5JL25Cvn9lSekAphbDMn7PkT1X3H
rz2RVIF7sOZea+rw8NdD6fbY5xOvElpJOFdFCJP9seGuKpKWeqxvgwpqxec2WiEQ
qa6XstbL/Q2obxEtKeZWHd6iOc7z/b3yxGXIDjDrM/RCQ0W57/k8J8uRT58Pivyk
vIaFCJjlmiL6fU401MJ5k3Nuya6RbEzYeLH0o9Yow15Thy2Vp6ugpIkhnABljwHA
BP2hWGmSGvRBP3oZpnL0YM41PMlxJ2No7bFkKQGx5Buqm+J+F3p0HSnKCvzUN7BM
IGlCsvBcUOyiJqnPHiBRuEOS5TfB9TvhzUysWj3FFYmXVZlccHDLHGK9lvbZXHis
+z8FmN+bCvP5S6oeNk2jS8AWJKJ+YEWt2T5DywK329tJjU/b74AK16Sww2S+PG//
/Vu9KPAsSpsoYMLxG9Fg/uk1gLHvqrSN1XcVDDy1TT2nFBf5fdRDKS58KzQm8+2i
Z6/rRk1sHEiZFS5/zOSVsXZ80MsV+jabyt5UKT1+dX+aRp/EED4Gz6ABdSIVPQ0D
JJFi9ox4D+wjydu35d2OEo5AJbhXQhmyNudCy9oS8xyKlKSVPRrqVPx8pfL24z1P
1KHiA1L2Z3xuJHpu/YwyeYQ8pPaLs9F87o52LTXSvYyp4Zq17D6xA05Oal6R1uH8
78x8Wfl6ArrKNJxo8qrOrj+rQEz2JSAauyVIdoOgBniPGzy6wDl2VX/bMSbDh7yP
BG91Y3ryFp1eKgi2QRIa7tXgQjstmP92/Ng/OrR9tYQBVr+EKHCqYX13Ov5iT1zG
P+/ri6kXMYna010/ADq+4TyUHBSOfFQcdFpeVnKVxlL1rC+DygR294YXITiiUGIp
mhgC+YpRfNJAEW8/QSKw7Azg01iiCHAmzLwOODQ+mU9S4K9TS36SN8crdQ9MwgiK
+6gdbqRJQFnOCIGIOtEX5t3kj2OknR8/Oh8mymQNOvY4nE4WTVKzNkdgJ75nNvOm
NXMcVVPXs+4JBQF2CY3LVkZ5NXWKkQL6waYca2DgymeKL1c1hkzxGm3BjP+11yVy
dIEqfMFlU6JqEro0Y6zMdBsYNpu1EJ9vI8KGpFwe5lncRiFBkg77igOIIMzA4mnE
pz94xvp5UZWhQnrs13DtoZi9whDjPThbeq4CP7PGEL/CpjzO85t2S+lejOR/oU6l
cmrNiIx7xqzqxumxoD9Gg+lqLBFTWukA3CQIISR7ZA4aTPQCB8noGF6Zo2uxfraH
ojHpbGXaHaGXtylu+K16VHsu5dL/k0dCtipVWP4ti6xnOngMx0oPyAySDN2UVLst
umXWNfhAhmQrZAf3E31p6Yoob6+wPWtjyI/FcmwbfUunzwpxTUq2TiRiFz1k2olh
4oq/mOwLNTei7M7UhLk7PczPqQtscF/8GUU3j0jgg+ScD/PoHHmUzfGFi8TSRXHZ
qjjDr3cHjr65v3OG9DjO5tAPeLddQDaIrlazlkF/cHmTQ41b6ngM2KSi5lkmel4d
097ux9cu1Xhb/Zl2AvPbEAazBJqiz14J8QFLiFvaalYL+m0sFCs2r5dzAFieBcl1
yjqBPNXk+cIrZwSmKwdL0PphlneNLzv2ZlD1HUTQ9vN8w34vP4WQIea+8cM3LcN0
9HUipha4ZkkxyTAGAorjsOHB+oIcjqLhkJSG+UJjC4JLWfaelWF8LD+ZE4/xkAOE
2jvcP1NSYpbAWeadJGuTH3q4lXpnre0e2b8N/JdsVFKPY8P2gl7i522eW5FsMOjX
kV1UTbqFt70jh/ayhHK6aW8u4I3x2LCEXcU60PlDmE7DnXFu6uZgNjN1e0ixB997
8ps5/Xmpu4pyJY+s62KNtR2W7WLYHixxFRwCDXGxoQ1YcDj8kr1SMHQIFeOboksS
8N4Q0w9nl0ZXlAgBFTaZKTFFPHQwDZm9ah9SH2qpeSQ7gxz0uaMyLSdztKkaeftk
jMScs/cB25JVHbJpEpclL1Wj3kF+uO/kd2PbNBL6ZlBXwmgKp/Y0/4P1Jw0mcIiG
TDumB/O7amshvhB6pjS0w2V/4Mk78K1Rk0+wNlp0MXXRNm9Alb5di6O/yQwfhV5Z
/7hYRJbiQDxWeICJZKdfTA==
`protect END_PROTECTED
