`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0O/WawRGsPNFbjpxjdttAlbINvPgC+1MYl5xrrbVKMRtLj+mH3a0rLu9VO6SfV+A
kSQD+xk7UeuO+Qbd6KC3C1nrVqyOw4jG/MrUnp4iOpgKuhSb8+oQPs7O6CQa+Kdn
Xq0cFj1re0FovThLHOGDb7AJ9H8nb8Aq6Pzx4kMt96/SHmeco5PlY3mHtfjKh7+X
ylH4VsU/iLJcEyJWYoPfwB+LIdeflMXFv0cdh3ZPTQB5bT/AWQPbv4bec7SpqTVl
StF3C/Jx5zE3SjBDJOfZyR73Ob75cTcsrgceIxqjr+kf/pl3kKFEL0f3RJRKZA14
2hZYKhzA47hV2DH7y/ukQ+OLlzC6zthGtPYH0H3zINKvV0eqwUStP+m2Q4lMT5yd
Zkr7J1IUsuByMfWyZVzGtsnhW31au7A8wseeIlh65Cqm2eoDviB60K5NwSIB4zmp
WjnVUaImlLNeO0/DtJUojLLGEYr+hfASVk37+gQ5WUxLK6cib/6Gl2QaEJSNhpFY
juoPL+L3dSa4xaUSy5i9XR13xdq36l+O7PdH+W33tYM0VGhs5XGEAAo0JROwX4gR
CzrdTtz92i4AK5yiB9nByifLVHiZme+FPFTITmOOnzGbZQKZVhM4E8Q/vIE8b2JK
q4UnKJ99LTvuYYG6io3G25KOM4WcBHuQiKu4IHlDFq7FHJ2Xa1Go+sXWPC4amFW8
bxKJ3O8EZr5aatZu54XtDs94doR0R6Et8ux0eAstEuZ0qxGerjz8WsMx5Qy/tbin
2k8sUEkLenCmVGDGZWR03wcJpzGNA5YYC0uQch+HGNSQtvN8LSF31TwBMyBZTYE3
dvt/nyK29aA1cTXJhi0ROECR/igNnCzEdFKbwEl2bGf/JcqyoVQg/XGX0pJVSRa3
Lx2ZHw5SQ+2RX8YC8hJiLCRf+cYPfwVBnQKl0eLVr/NgmEVFjwpU+tsHml7y6IK/
KjPBywhBhY12su/Jov0nfFw0+EfSrjygW7+FHEaDuQLTEqQb4+bQU6tg9nolbfVJ
8wPzy80YYhcaFWScEAhFrQ9IocGKkKNMQ2nhbMUsVLVJuJYmo+t/2gC47uXVjFIY
QoutJ7Vxo/Oc64potL7eoinzwBtdgm0/aIc+E9DLq1/iZwleKlKklCWnjtt3kqPN
YPuLiJcQ+Mge0Tm5ExbwNHbmPye05I9RiTDdzxVy2cVlFMSjzvlu1XlrfA59v0Zz
/F5OpC8rblKwFoihxePC8i3kn+FcUwsU3J3F59j+g9NLSC8wpYqmpyG+1nW1fTvA
Ll4CFtMu8aRNaJDXAylDYs9RX5B19aExswXuaXJWgH1/50/PTZ+KYmVytVfRUTwq
zziQv4eEZItDn/ytu5aps46q6qna8v86QYZ4+Lwna6UHmAgV9N9NO4pmOPWXiabL
Cmc7esrjm3YoRmLj0bP7uKKfLhAAq9AXz+vR71xj81VUU/Pd3pF3S2EEGbhtZLos
HF5huyz2SMIK8D4ol4gb0LUVuyvLAKXL8nuf+ZKi7xrqTFAWZs5s0Fl5G7/SByjb
Uh+iIdUMbHptRnBzl91AEWTo6oOVOTA5w5N6noY8nmvy//u8P2SwYnnj5/mD+KnP
8B6plJijCbk8o6VyrjzLDTpQSvFVqBwRhCa9Hr6OjEFHWo7NDDVkT9nKSeclqDm0
f56chBIut/mXorMYzwDeEk2QcyJCLvIupMjC9EhCdVWSX4qCxqaiU3TW2TvRXk8Z
i015Q1ONz/wKrYxmtIsAz/QmvPlVPBiK/fHljtwbo+mFR8LuyXMvSHeGwzY2FV2N
L/ZYUDZ1NuEGeozVPdFCKeXWJ+3uruhbHq8zsLFocvN61h7uZS38pkD2vyR0M/TP
BudjJ3H/RgxUcvxAsf3Bsf/aUOP0GRsAp5hvcuMrTuR6jmBk34UcjJh1XBVWEGq8
xG7zaD94/uFFgJ3LiYjMNvrhIq6mucPVEo2gUiIxNTeK2wJknxCaXOqmHvho4Q0I
0NcaAUbRdvYCpftHIp/JJPHjZ9esS49OUqij/hPp+YR/lTTN6LU5Dr2BWVUi7vLB
/WGGnWVO/b2BrlnnqO+YO8RX8Umsx6uzSWeeZlwpkMBip8/gGufn4uVbEf7ZSx7W
9ANgNIuJTBWkhAJXEUffZ741c0pEJyD213losuI+NfOtxizBB1eL3b6hxJkWKTBE
ACoNJoqeJAGvoHTVEt/xndlP8NP8MwXXaDmo4Yitx3/r01yO6zZNSdvMITSccuXH
aOfXVssgt97n2cevoVPMIVz3CyAGCO68JtZV8cj82/gIFPTDaHebJqBv7IVKaE+j
DxY6YcwHhoJOaAJXv7yAZHYCFmvsIjpxFOyTU0i5UthNulMc1U0fnvkDugFvdGr/
s328+YmGAaly6OdtfvxH55IvLLL7htaCRZOnq+dUKzgNbx7yfecA2L/S8vmTl00A
ELeKUjrGiPP6kEk63GKWJpr7MiXQRqbjgyCR6ePjo65XxYttzm4dovHkYFz1v79d
dubuCr7zztckcqr4l8Yjeh+n85DHhdPRs4PEj9pCXhJpj6VtvQ3clJyaICfNKLgo
w6Lm2GI24fODQg6tFys1i3RsDPEHB9TuDCQYV1exf1BQU9lxWTeX/XiLDEcT92lZ
u8JufJoiTjEnAb9Lv4Yk+RATw2ol1WgdtXc09ycWVgT5rrXmtsY36HAZHuTfyxTl
N4J0ropjJCjLogAFnXWOl1YMRTihsmk807bXTedgHDTwyDlNZxQNZ2Glga2Ox+WW
fWMBDeRA5d5loWKvuhuf11xtfkDjwPVSQ7egMPKN/iZAEhtqQBuKT6/uuSwwxu/N
3CDktBDJwpFaVMrGjTIYMQq04hkfG9SM15KmI104ylSwZABxHQytBn0XeaLU8BLf
4W5MU7YmaTs5v/FJ/RD2Z5k+86lHcRC1AO4jlwjB0+8=
`protect END_PROTECTED
