`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkh44j1Tx5yNlwsItYuXngJxvPoG+WgEfl8lRtoZ5jE49QDBvhW0dLuIVXEcfRXf
8zooxVns4xoIlyldmeF0G/mx7QPffo2uCq+GAnTQWA56M7+yT2uv/63ZYw33L4OG
L8aCxOJs9AMHZ5zpIdM3jjAe3r0rYprrN3K186Idz8jdsfvQzXq3nK1l+DG55rjd
lYjx0/e4ehMPwqBVCrPHY8SZWiPM9wujYidTbdd9LTwiv+tqCDDTYxnTA3+VJau8
hn9zFWLjYu0udqvxSJEhFuAug1Z+Hwl3lxK38V986EiO5vqJPULmDdTahbwyV4j6
RhKT37ETaZfCQd/HTn/qHIe2T30cBbkhGkUgkQjSail0M3BSLPJOGqRNTDn0yHeo
xItvWCBkd5vDxEKsIw/s09DL9Ik1FXXxBkFgBZIMqzWrO0OYtC2xJVUWdRZdfNgs
d7KA30p7WFvkUXN3FVTcZazDAGbl1J5PA5blYZX+84SFbt7g+/eFcgwDkUBodm/h
RFKHN2QrV2AyHX6hec5YyLyZhaCrGK1fDs4gubc7oJ6Eu8HVngaWpDB/+bJ4X/43
sGsj+5dweb1+XFtL/3XIuoX1NSMoHsLFNn3ZsaXZsTMa1nQHfCkJV6QCw9ACbTx3
Cr1WVR5PbXZJTGmNa+4faFq2oxV2AoiBriGMK6/gFI5CiDyknk9CLvaJsp+75ma5
+oSN7gzOLFCMy5ibpliA2PDHcPmVBjHwzKqWL0uuam0JF5MP9L14s9+DrQQZfi0b
wrRw/MJibn8AHAreb5Jx36j8zzF+9TIjYS9c7Kf+uR3rzKlfoonhIq8cZMxLxoHv
zs9r/aXZ9W+IlAN9kk8pZJBQ5FxjBka2DV9kuNScWi1BJTaiw0beB3ldCNuJyVuG
fzjYINQYWpgxv6YkFzqynCOn5mHW7GYrnp5FxCQnNowcmvOmiA076JoQ6BjyRJZp
LO7aI0c2X8RLdTVNE7xry1UNchHZeJX/J1CoH2tPpvUgeOeoRHUgahtGRDn8fm6i
wjy0IiWuD9FAmFcjn5PNAv6SaiyGBCI64VKwYgtPg+clAG50uX3Xi/UxTGfNcZ6D
nC8FQNMDi8vGlfN9/IO9aM/GT+Esy4giHCDB+KQddEl1lksJO3pEMrupKjEmMMvW
L08K3L36aK/SQYJWLQKqhAYBVXta8K/RveB9qN/KSP/5tl0TYtQPQ1MkVE6oDpyy
tcyICTei0pP5oDG4T4v2H51Gfwm2+HtxKaywbT9y6FvVJwVneAyFy44RitG7nIN1
A7Yt1+dZWcy6hmvHOB7yyTtVwYGqPFx46d8vz4KIVFTSbolrNracYguHJNOCdj7q
vhZ38mQN09Gg1rmdY30/EPX+KCfYnuWHzMJbJDkFLeu7x/mS0fhT5fQelM4E4Qku
3HxG+1eCfT7+VgmQ+5FKAWP9AV2tXIYualgUICSzUEYX+ihdz2M0LvYEEJ82UWhE
Xh4G+sccHFGNTPKIkTchaFvfibu3eeRRuEaH1E6o2KQvLP8H8cI/PTtH0WKCxShP
5dx/eRNaYSHPDjouwj/44WF+TEQ8Ccvqhnz1l7z5TThHCjezbZeJTC0vkEV1p61i
fruFA7GnvE0zI99aE5L2I2anQeewsIuLpIAg93GuXVJkbo5DEQC7NPlWrUbqTguQ
e02jY5vr9RbzwHhlCJSSxhOUH2KgDkPBO1n9VrHIMlIoeBSatLwW2cqgXjsqYXsz
78FITJpkA0bEMomGvNVf9Hv/7EUOgRUA9GGFhnAxfUZKnMi2KxWHZbCoonPCgwoj
VergFQcwjajitIUCaB0CRFZfzW40EhiNtJ9gsDY0pVTgIkE1MzFfYvOOTrYJVu/9
E51cceetnMpXM/4HxYiV3jU2kf0+LHlA2YxtldMZFYcbdvD5cPNP4ycLAlvYx2A7
0b0GWMjynqnfylZRd5LQgll5PMTi4Fjq/9BnZyD46GrIKhCjtX0r5mkOAxdc8bck
bYo0OpV5QI6jQFqzjMvgcKBawv8xEHU84gLivJWOY8FFHPy9/Cv8ujREzV0h0hRR
vG+tHt2kqMd4wNN//M12a1FDiYszE70v8WFgx7W3g6+24J2mg/VGPMFj805lnIDR
yoc1t/lNWVgabI6Tgtwb751YPBjczMkY0cLT9br4NswScS8d4soEQaTe6QbOFf9e
MYvXFrV8vevvPpF4A1BBLZplyj/mnkT601wtQiNWBW0aayhLr7W599HWzcnBK/4I
2NWhgWZxlTK5vpAGcQ1Zp6VFAu4iztph2F9/LpuixFwxcxUu/2dB2vYqS6hXfdTx
G3uaN3a5UG1ueNp6qzg5DCOYR82R12ihZGLadHZ8yog/jA5Gmtw5aFVRpuPDmhRc
w7+BAghUdnGJd9p6SakISQKrnyuSiTJgbm1C1/xiSsu+VcxZyzuf+a7tHIZUVe6j
PsrGIvoC8M+T/0la6z+moELTb/ZtLY/z1NCM+DMKF3FjrPLrUJIYOT+fU89Wd4k6
1qEgn0OQsRIPQ4W573/fDn3SarN1sr11JE2CAL3OgX1NtJgsScbBAnEt3FSEQweH
rMRr9SosZ0++v1EhYkNr6lD6RXTBGn1MkFl412gMQIpokiPHoFAjgZ5JRJ80xu/D
VqihgDv6TQiA0N7J8J5gQQB2LULWCU4L63OvS4j1Z9C2QMfmlRTfo+b5sh/laWh4
Q1oPCCxg1iQTLE7dEZ/okNmh4FWWMSA7F6QacDbZGSb7IImHiTzN3FLRooPUN5CS
ti4zt57rxxWyeBX/Jd75vBr3XpixWIv+QY2ZwPFvg4X8yAR5wLo0UhM5Se5zgyVl
odBwWBU90ywqeJrHwqADIb6SRlrRA4UN8Di7D4Bzd5yuKwn3ymQ746AvChMFEl9G
D2CQ5zdFYPzM9G09Ttxx1Qs2tOb0JP89bglOja9tlygIm/efUH90p2Qm6l+Iu4Xi
V0he/SYAE1aiMe7PXfj7iF+1vonCom1jl+1XE9qa1Sj3Hbn8OIWzgJd2D2Mx8XIc
aM9eSox4QukiNYYN/pDRIh2fqCrRTVz0VgG+zhXBYw/ZGnYWzIaGJ6vGbl4rsnQQ
MABuz6T3yRJjzmafwt8RbKddd8t9ryKtg7FyQRFq8B2DRLfMjSthVARefxXZXy/C
nd76iwq4yPoLQq0dQ8ab/oQ58YwnW9XpfJcrkXJLphaE/671O7DvsjQd5q7E2Qoq
16RCPxd9Wyx14bJ1u8Woi9sTm36OGd9HXO4od6RAqQU85z5CnqzLgVZG3GpCTd+H
K+ELeg5YmoILSOK/a4cIGcT6LGiSDNjojJ+lvbnw30JjnbPxjtDKsKyWoNCgc6Gw
NyakYcAJGQ9XGdsRYwmxl7CdYOYdXLNH40TCTB69/ysYSfwG2RCHZyViJk8o7mAw
KYt2mnNe+WSTbKaIbzvLPW847e6ZMzWFNUzdF/2+dlp1zuIGDqdWhDgPtpTnlmCv
6ebvXwd0EXeZgBvnlwl0YUXelnzRd/qzrZu3YtNukjEPv2S8+L66xHpXoZrreEX9
7URW3rixqtLXIPGdzG6YxtnRs+aj6KOpm6KFXmI3o4i6/fQqWXwPwcoOqKdbjmvG
4Et8jigjf/sSi21Zu7LfqPluIOSZn2PRr+hcUgNwZdMfE5HlZC6jB/NzEL8b1ebG
+aAveT0QdbTPGpPE3acl1q6DuA3wxFA8YlHRjvtIpIdvn7nJWbI+wQStvw4KQ8F0
hvCARdTJrarH3Ta6BmDrLg==
`protect END_PROTECTED
