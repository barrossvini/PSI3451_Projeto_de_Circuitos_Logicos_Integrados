`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yDrMaNAgk4v092NvlhHCXGOzVaIJM7AMLZBMKMde6b3sMSnmYa35qXjttjuKwXy4
A9Rh9ppEEjC0xPqppDD4dT1UqroSqH50EryBVYLNLehyatJXa77MEUpf2IeJTjps
tbQ/b84kMZOZm5ZgKq1BH0bJVpYM7rPzFCSdeHhhbCKRA+pstJEzD/kw0NS3twBB
G0ZjBYtoH1GXUfBTkM3hotWkX6bPDZx/FnmscnUeqZfldZUDdIB8aRfrN+BFhRy7
2UsFnFuE8FddtKTCHqW90gk0ZAy8ychYZ4Z+hCYcxj63X20c/evaFwXLL+Fhz/0F
vzWDl0v9NKhB7s8HTJ4Mt8W4RT3OXfRGU4ZS9ihjPIpSqX7A4wtL6HyCKrW0hmo8
TwzPbpgp2bQU2X+JlCPcq7fIr/Qm2k5XGWZ5V6nj7uJPuHdXUNxRfhGgi+iCnJ0k
SVw7CwQN7WGgYezRsDm1qMIyPnJcSHFQVkFt3nahnp50KpHKS47Ud6NJJ1oiIrqY
KIXjkfcuBR5BuLf+mNQs9hAC0qOtqGUcNoOAj75R6wQ0wqfVgDXJ2BqXFpdwCtn9
fhpW2FE5CP6+IoY0oL6XO8A6u/44J0ACd17KQjskoJeQTUGLOkOq/9DeVPRP8pbH
8rYQxGkyD3tbrEn6BKBsEJVwTWxZcb8DFbEXAW8Sa4M+jgK3pmj1orpkmZyj7Ygo
I4tjho0jX6eZYvQ/AobGFrAOraZR6wLW1qQ9Zj/UVNc=
`protect END_PROTECTED
