`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L7h5S62iP2Z6iR2E00E9wvAVA9zDclloi3SKgGrqkpAIiJs0hg99ZXDBxMA8ihJA
Blk4KfO+sCkzuGHZgrfwAqUHtApq5fRz0oR9Wtt0Yf/FKRxAFme3wv/TRMNYIK9N
piJhcYMb+i9OzDsHFuawC4/IBDZSYA6Tngp4N+QktarTuEE8xcNTx/PgNYsCzp/S
yKhUKw41WO8HZxoG5d//zzGWI6EcOM2SlFgGo0do9kwSVidBTcTxEQA+lK9kdKys
BVE3eoInmBKi1r01g4DHZF+DR3MNx8a9/u7Csc8tmICF+qXdCF288JrMSCgZr5sm
bDzApS2HV82skmSemFnEXctmLtQ5TspPIsvfWmq/cz1Ux+OzjPk1jHqZVtc1SN6I
/Lbk5JdaCXqY2wMON2GV5IrigaO/CVTKDPZPgccbKPUpTw8iVW+/cTcGEPYYO0Ws
TyjWoY7DIvRiHryc68BZZCUREOdzzkSZMD3WwDDQBYqCtHQPygmxO4+Li18dLd09
miVQLlVo2ktassul199L6HwoF+t6aSTJXJeDC5rvAEGbWvr/CwQQF/VBDeDPM+qR
o9M5h5UXjzkXI6BXMuYzJo/K0jdPYJwnztoaS1JmAaknSoijL0JXGq5GkFj2qwf5
HuWKdC/InqOYIRoXBHa+pVtiB5zqHxELbW/fj2BcX3ncft+zr8pMu2aWFx2BnDns
elxo1HbiiS5wP9mA1uHPyBnFxYOk6dqN6kqFPAjYGVuZP+xL/5HX0ADKO5Pq32Ar
1Vz5YW+LoimXm4fLE9YnxroxurDgdimmegQyOoXGa0O/s7m+navj//P8hAFKBgbK
gqDwBmfVCavOVVVuUa4TEf4vyLS+iTkO8HdQirPjJ33WIRSJC0pt/7Xhrdx7pb6Q
Ky7tFcz0b8hEU+ojp3TqPreuSxJWt/Y0rtTpmTZnhQUt2cRZSFvgLTw//gLFCvNq
t9qRrT8V2vmoYd6HUqyq32gj0vomZcg+uYNzLDI/c1MQhVPA2L2iLKgpqoY4XSdj
MJ1qSlu4VgsVqmzrEEAEXJv89AmoeAyHZ8vJizBr5DTFMrb2XEfVkqTswdkC7Mdj
qlyMAen5GhVUbOjCzG5Ez4A60EQe0zZ/YBaUQlgZBDp1gvUK84AdZecPZP8NGJ3R
DoZSfPg0O1wCEanFeplyXWRa4C3wc4eAf2eLnrOzqGdNLCOhpzhQgtO63PSDMwv5
Ji2WouLKtUkWu6B0y19YG2hu/bU0pG4jUwVMdzukUBE16bR6bHDU3OmzuWlvPzaw
tcmwzfiKh9vt450+CdRlyIYPb6ton5xWNwkZoVvv6htc7mGIrW3je0ZhYXeoNFTw
bYdRAzBCYKNfoaL7HMz4OodO98CXi9Ltdg02MjEtzndyRrTSeueay852Jwtba1hw
hpO3VmAzVMzzh9t3laWgyah0ZjtAMZmhwDu4yvdKZhRfr4p4E7uSTUuB55avLeQP
`protect END_PROTECTED
