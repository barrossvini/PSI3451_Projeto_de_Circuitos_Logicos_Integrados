`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fko7djAPX8xfQu9OFljKvJIhg4A9i2Am1AfP7sxfks4Sm5OIB0ZD2RbdT8ttfPPM
ykLm3RTfTrS2ORaeoxlzhBbTv/GwfbO/YrY1VlimoI8P2wZzemfxhRdOydgGLueR
llTN0DWztfMXU5V2+DQqtCgPcc3s+1Eg6ESQUs/WoUKpQ1WpTofu6yd0FFGx4G5G
hEgKF8Hrv0/YVSP4KuZBpQWYklzblbFFhzxL/FbPgs77AL8V4TN1YCtHk9RGu9br
JUSU/SBsVCQ2EiwHxQXYSuRgo36UbDOls4yJ4KHbAzEMzp6i6tUNDZyaa70rsJS+
tvq/d2XKEVWXIRRmg0Lh6rvUcbhM/jUNKS754jJXhg8qTbp4H8hKdikRtyphCntc
8SlZr8BMyNYHSJAIBxwZUJiusn542wUdix3eDBSGr/bRs9DCxVZwY68aRzGZEPz3
hSG9Cb3yGUItsxwk8C78VOn8WErGBRldNFP1txA9j8/jsKBqB36FByLp+cEepsMO
eHwwSupeLKt8jjCHc5H5u26ofUjjKxrp/q9uQ3t/Q2yltvdpjZ8fqS9hKukdqEsm
zUreDxQZ+Tz87BSqebAd04MsE4DvyFCpXL5doq7Dn86KLcyP23OIi6wocXLhxjMq
w2Pm3t9ng11qvR2AiPsAOlx8oEaFXRgC0ug1hD2CpQaclY3RWHxO5q8GzsAJDou7
GUrBwFvVaah6B1Mr2zQZX8XE4/1EBiZnUCZhzdqJ7hAlTu34JuKdcGT+bsBNzSz+
oSWdCtzPJIg4fog3q5qRLukFbHJ0jyqTGx+NLVT2h/hYhSY+0m+J+mMTAopxHQxJ
/ghVQXi7osluA8FqDt6LlPWqOsEZ13huzzgM2iaorbU3MSro0EJRs6yr0i1bt0OB
ggyovkTE8DODsYkrS3Iubx8DXmXp79rnswoaWQZ7g1cZ0UcpxZdCAKjTSQ8fCDBe
kLm584Z+zqGquDzG0/e6x9aiOa0/ztQfxzM9MOUFRGnhBjmnOsaH628nfFVBfjmM
n4p5RYjU+joDZQh7gKn4FOOyPkyLNNjUM3DtHGjtLyu9x7cW4lJl/a+TJndT2wVo
ofVAAa59y3P6Z3PcPOrI9HdKgntfMtMm5dQFu8+y2ezGan5BD0AxY5MaccbkjWwJ
v1QJ5t/Gy2LmShT5s+cwKlqUlYIRhRI/+84JKpDUn1t5W6p7ARuDUk7tZQ6MR7+v
WOUuxvosXkKDHi7F0Qqg84iY44ai9hC2tE8Ztqt9zWg+SeSAkbz2ztKqdeOMrLDu
MYgUwBmqSYrxP28j3fvcNZ/aloCNHjaAMKlXX+qQ5ldlrnQisWCPQ5PeWddZvuc+
YPWbX5tk5gM336o+xc4//PZStwnnky1b/MlK8IDicF+BvqTdxLDCTO2/XMPtoQYV
QnF4gffKz8Tcuiu5gQ04dS6sMp7B/B+kZcozWapoh+ajYvZOpxop/yl2XkYeu5tT
olSk/FSWnwis3H0MW2wi3esh8SgXNjVCv+q+PzwGgrXm9i2y4NYMZPyNnVX4cbWe
UBYRTt2+c+mc0tyofEUZMwIDlo6acu88mFL7/Xcrk1IfdO36YyJk1uIxPdoHdZtO
xEjXdmzk2VYYeJTGPWSd1nwA7GPZvkAuJt/ZM4tPu+gKYRUZN09dPys4oGK37IH4
CQz3a61pM+j3XLtFyKPaCqP2uIH9KGLijGa/kdeKNJxlCerrS7/AkjghRdKk3MC+
0uaF9d7R9rwBdqUrQlUCxRh4UUEC+Rs/1b0mJwvFJ7bUpgmDOm8JljsHvrnj3XP8
Johtr5/76bnm+9RDXBVD9Y8CV4lCUP8S+MNqOC3k6BAtGcqF4lFp6mBXpoXNC5OS
iFQ74ZnV6pwjTNM5YH3nph6c8uM5tdkP7XehUD4PtT47jIcIjZ0IUTeJIxx3tksw
JZvXGbSQ122PxYrBFEQ/X8p6Pb7mEUcrCTEOMSVptoL2Rq15sZCV+YZxA3XTMKaK
hy5KISVo4lt5m/gKptXlLeqqNT55yENdre9/SAHsgLfr7yWicRTllFu8n0pqhdUJ
O6+ZgY+vK+Z8Gla9QVCXtW9Q2KfRb/IMhYuzcCF8o2m8JNVXgFT1Ng872dADuBP6
O9/yD6N2oDIJUsBOrJbTN5ZF/qcWxkcFdynMAJIlYcshw7f0I/lZFN3JYh+KJW7x
8gP5qDAFoxgVSWte1XqMwwVutti/D1v/Q44p0fHRq46j7ugzYmijrDdpHVtr+GKH
a6JrODRPlNP4zayWMPs4AVKaTJCzQxqq6yUr2KdS2W9IzZg5sIsCpIOR3+qaID8I
zWd2hih8qmgkFFN7OYrIZ4ihXt0yq+sQinZT3Ez0ayMgzMzWfCtwzmnn8nurG1Bx
+gMNeEhZYZtH+jxQmcb0RXiMGPC+qDlOUxGztbrpP+ZsW7+RxiJ2P/yEofpg3kBJ
`protect END_PROTECTED
