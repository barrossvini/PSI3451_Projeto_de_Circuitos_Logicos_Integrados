`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sr8eTV8ghkHWCMrbcY4bAR6/jYg55vcTswzYXYKUKLJ2bZ3dmeRjN9mjYQsrGca8
B3W41ZXtOiCEgbizaJDQN76olj5221u223hXdrRAlLyCH1Ebuo5pUt/Gi4PmJsX3
qhqg8VQif8hI8qanpSGjD6JYddp/DoDWcnlLu82ryUZ9DpGfnWiRNKj/JWLMeSke
FExLPE79dnly1jjIFKjjBKbE+Ce63OMDpeObzD3rj+Yjgl5cErRTevK+oGOc/LOW
KyLWmd4s66gx1Z+sbNrJjdth8EoO/VC6b7FLJ8KjF3cDtTMa9hGTh7aFbrBF23ev
DFw8lqk3rG0HJT1DbFKf7DqUqnqiZSxeYL+mDYOlmqRKRkJL9dtcmiu4GrBidzPG
W2KsEElrKp8eTT7ZLOhZ5W5c2dS7q0Qbx/5CSkeVwOo86Ibyy47k/VuDxhMU6WZA
e63AOtp59ftWJZhHp+36TsLkV0aUYnYrlwMH7fC6H9r5Gj9ihtCFoqdGfjNGy2uv
a+Zs+4MAkonaXHxzO8FOu7B64/uKqCZDFpnkqLwf4p7XtsOMq0WecgkKOVER1ri7
sW+vbJNAK+tLJI7ERLEryP8cv6/pppnMctOw/khJMVhsvIP1GBppLcxByouwyMSh
327ZRC9lJydy7QQXLuNxG9GjF1GF+80Zo29uYpOM1rm9USfpwEd3aTVTMA/dX9O3
UCHUqyVUhsxzUcj7/ix5FcS6CiSfOzNdx919jdduJcAugdyp1xADS3qytwg2FX9R
Rr6IEXYtQsPadmNw4p9Ijavfl2IZMTPrr3UGy6c+tiPhIbMzDMSD2TQLnfPiOOpP
Kskx0l4cizUYublRQyyeDo/Ab+P7mU3YD4GdrAiXeBZlt3zTs4Pno0sQ2u65+2Rf
40QxVsmG0daiwy6+1RCrH5F0Gz1z18RIpufV8W78kSlQir54c1loYlR6BWlSXup1
MvjlPYyiEXHHyzPynVes4NFZw5m4GXomc44XI4XxvxTqsdKrYazen6qmRB+DcSzd
3cbedFLOpXyldv3fqhBsb+xuJRR8p3A0dvgn/WldQ9ZBH5K1VaYBKj0OHGU8yxuj
dAd6jydc5d7p15uAgBwmXPNLYvUUGp+fEeJyjlTHMT/gfYVMzn85Mv/THhfpUm/x
64lr/Jvo0Yif29BNfvXfjkC6Zcny1fS/i5RNAc4hF1S9HD1aLYSNuzQetkSMNlb9
WZsP7dfMfDeXPbijCNHIsKjBgARroQdART6oLo6kf/Q4UVSuLzMKBvkM1F6dCzdu
VoPcRuIeD7oZhUJda1voY26z88auWgzVJkwBmxqlMGfBzqAXNGyWTUcVIQ4sgOD6
f3yJhKE3ia9799+eOLPFOjMacGV2YkarZMQP2Nz7mxsifldKNfw8/GVhf1rT2aJW
Wyvm63p2Kqn+I/qVPcDSTqIuDTIz6CCAjdBERKu6Ax+Z4yaHOSauAheWpZlzFGj9
ERRMr/Sisj1I0VbNy8BbuwGSnhTXo/bXkQUsBibOlKBPSiU7USCZR9OmnaEmd1l/
mg+A0cR1A6dlfW/Y1B8SbvdJjNCVeGQlyHcFiLNvbycO60AbjChu0aPffswOfyKe
TCJq3+R/7Wm76OyNllJON4QoKpqpRXJAuPsfAD0ogaiKGXQWXp0b0BILd5xv0ImP
jTXjVWEd54G9rIviseRamgjbufZXZR28PxTL6F/Z1N1qNyR2Bgz3pel+dQaSWqJ5
YLVNO9uJ7hpiaCE8WJtg7dpVazellqSPuyUqGI1LTNLGWuaYElD/PkPQPcD7GOpc
Uv7+escT+B/hK3V5zoAWOuX/R4P1cjnDDW5T87Apf5Hh2p3Qq9xu1ENPcyfkrobo
VmZSpUtAO7Dhdhel66i01Nns7F0Mdpg1PHUscuAN/oSgKjMgoUPAFCQoo9v8Ue78
zhOcegXp9ZiVlFCz0GfFxB5qj+2DqSIdeudFxz3Sb/nK6UQRb6lhEt9HyKx5LQIn
V0OveQV46+8/2vM2Q6ZSC+NtpCmhluEeIBZDFPvLJQK6MNq3hK9sn/KTQztFyuw+
qbT6dbeX4dTSBJ1c6xQZGPrxMvufZMw/WEr/aC8bGhBwcidZ5RvDL6/688e/lI2r
K0LAtnarG9ujTJ98JutEk92FBaIeD6WNqqKdVBmx/wlh/W+xIw2xOuSktz/GZidq
KK3oLrFDpSqHt9vk8rPGH16xUx2fyyIr6nu456M78rp3P/l0PfQiB5iig6CrvetJ
0khHy6lAK9EJyNfJV6sXhMD53VpuYMcuAeWLZl7S+GaJ9gQnP69ika3J27WA/LQ7
WCzL9gs9IwAAApWNHAtc5QHcuNvcEff+ytIBI7vDssjpK6phMUuvzRDSgS5FHszX
4Z7ES5wm4XBq61c0DJt2+6ZSGgTi2ADZnQPPKJ0VS4KoLASh2IhqEPntoxbcFoAA
r7+B4riprHfzRbisjogoLLgIKh+X7rNJTwPpLHGyQbO4MKPphtBsGVlPKR8r/JqX
ayMymevzkGg7mYkrQTk9iWSguUwlRbKqg1U8qRpBJmwxZosrP5FnT1+9kDZPcspM
Mjz1OFX4XMh9ckk/2devZVHSYPillKm1Rk69FZLEFpef3GWfCr6+3LK2tZPxl7ht
6nZa9UnrjwWYgY7dYIB+OFY1h+jrrrMHEuwxtOsPFAysTH6JsoRQsu2IBBVaFuOL
ccOd29VXlPJIdZ5TYxM+tiwEVxQoQYa5s6TALjTo/rNLbSERZrPSJK5NS5VkZFpG
MYGnbec73ZSJtX+w49T6UZzcsIWao7dbfJvzrPVvwZU1yLyscCpsPGXNcJZNc5Nt
XXfDd606HQQc1uJAYuKYL4TmwJhKTBOasLYQOx0MCR4RKv9qpd1T/pyIG9gcXZT1
KbbgWtcol9lzpJ3+ypPOyrYpD1jhooLKydDStiIhxNRKIUTL5oIXAV2LTyuZeKV6
OCzU3uxoMb5FDnBJQs7nCLkcXduAOTCUry5W75xKXWznybRR9y+/SSbyL2AX8oZS
wVeBJ+MDCInGsrR9kjjiFzHyrjbi/0fx2yjGrBLi3T3xs4ZrPunOlhgZGoMPAh79
s6I7ucd2XNHcchUDdmRBC71QXrSHOZ16irQGTmvgI562jWbQatY7kj6Sr4ns5Guf
44vIeLxwGEn4Bnttjmdqm2BFwgABPpCPTLJ3fjvGBFXv9LrK50ri+tFLJk1Iz7nU
Yllp8DYNgbY4K2chCQjpQTpu/STRrYksuPfw70PqpJrutyAeuXOIH1CcnrLhRlsL
DWOYkZ3yxQCOxJz1sKKzLZuWkyG8DAPyNDcgtsq5XdxVZ0D293TPYjWUQvycO4R9
Y09dEtwQ0GzxmEGs8GDAmyaaOKxEFKjR2JZ3AoHi3tR3suFo5U7ULR3SNuodtGE0
0DsAO0xFFW7Pl3C408RDWLlsX9A0p4gMaLlj8064pK5WBstyl8Vhamq9UxfRZtpz
+vrpLGDkLdYe6lD2CVgFOPG2kjzvEWdG7oZ7AHIFH6nm0MX7AGLzqO0DFpbJFjpa
Omefg9ESuXS6xoM55AfgfoTgiQoogDE9qnna7mG2ZqnrLl2rmsBvfnPyKN8bdAhj
NPhRastfmDumBk3XoK32/M6WWBsMJD9j79gbBfWAQXMzUFK/ugInZ9psBr5XJkK5
lQ0wnd4Xa4plU0SrPjhAtdzU8Dww6faUCgeQNRdK1XCnkn13CYOW24TNyTJ/AjVF
QrBmIe5BDFyqbuNstvWs4Q==
`protect END_PROTECTED
