`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V8PWWGroVIMt001H8uIcOcNPqZk6QfJDs8nEplpaZ0vipAWUKWQX7TQBYQ+Om8Tn
G2Y733F2bKwS9qg6uVOQ2Sxho15tmqgTy5EyINuMwYN71aHOEDJ01oRS4ILo/E37
a2159EmzkLUpZbEYAj6WKKeY9ler8EydH5NzHzL7TQhkHvYCvbMYD+Tp21oMiMLi
hebW7EkNrP7A5Lyl6IuwZ/bW7r7a2X4XRbVyw18r0t8N/+pGmH7+LYPHH0yWyEmo
8+942xVtZqJ1vuTBPwtCN4AWSzgxVI7Kjg1VGeAeo6cOfsS/WQeXXmyoTYgbmfdi
OY2A/BxgSrC//4IKM51LZfoFT6D8zfHKTUN3lbDTxT5MQKpjrnA+lsN289RKL1sg
xU6tIBqGvKM3C7wfhN2NlgMT9w1kq6tecfjRZJzoVWCcSFaF4hPqVZ6b1cyqwtgL
VQFHGICpUBdDDU/H9rlwd0+QRpWTknpFnZELXqQKs5XDqq+hKM67LQpo8PJhNFup
4h0c9lIMlB1T1kr6lg8aM1HEdV+pyn2hq+IuF62HiqjOA2pGXPEtFlpgKynWrylq
FXpNftz8yViGmUBYapDxjP5a+69PaKb5WorAJVQRaW3VuasA/AdCydAeltMsK0+j
igWxDkMgnS5ePLpfMDplYhdVUKOrIsax/FzhaIGzXAQ8EI/KQHQ71FYqK2giR4NT
HJhMqMCiXNJ50ICRtFyl29L1/ojnSHDKkBqZ7KiVhdo=
`protect END_PROTECTED
