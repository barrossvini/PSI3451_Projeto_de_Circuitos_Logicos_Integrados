`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x5ECy0aPira1FyUG5i13esVECq+ZACIWqAS4jdtjthzS2b7u9VF1RfNai9DnZLOW
90F5xNAI9zXAyLdHawYmBd6kavtkY7nOJgehwF8VzeUzI6z2Bh/Yn2Y2ogta1M5A
+NLWdQzY6BMNFbe7VjpTlw+7et5gsBQRTOk4Ono9wmbEwsyF4yXLpOGEqhmz5rOh
vsJXRu0fS3gMfazQbETOTegzD8tsIa6HPxvw2A1tcniV2gWSi/ndVkziz9S6f0D6
k2OGAcgSL19yzlfT5lJlf74UXjnomGj51XNkD5oFG5a+CPo3t+w6XaNcfBQeMXpR
Lvi/f4mrjpCfpHyO3L7tWMxfe+N4Ybwb+cYdfTgfE8DxUkd1aBbW9BGLemXTWfBV
g3WP/lA/FUUTOlrki1crFHe9i9XGNcLUK2UBnh5Hf/cV51ksovb4ohxqqXYjl4hl
v6EGC1yNArmfW7++zgzKiZlpARHPzD3sThHde2q93Fhgrb/nFxs4htdaviGPmSNP
0zw6n9R1RQGmgCvPRBZ6sj/e+xD3iWQ4lQPvB5xpJBbvrl7ziWr7onCN+P4jv4uN
k+sxlClmImlSPO5vYsiUtQ==
`protect END_PROTECTED
