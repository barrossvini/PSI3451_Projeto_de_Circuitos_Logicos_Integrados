`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N93b1bOfHgy+kRclymLoGrUJaIFpLgV/gEMTwqfSyPDBOsI1WViQIOKU5wX82b/1
u/fHicvXsB54acdljpE/8+kBrrhp7pJTr7qR7i5FlK1OcBRSS6IEPfts9jxhiPLi
BzXA6EF/W46Wy9XepWtbNrn8l9ANmmR7ULwu+J3AApFkivsPXtFW/yMLK5iCJOE6
FKRVl9PwcNRsx2ZSnT0HmKoLcc3ADFbyO+9QgNrFSA98QzDLHXHS9NR4TapieCJk
SW8qxkyt9ldjYr0vXLXMugrKXgf/Ee5XIUGKNyKpAFGinOb+GjiT7/5sy0EWRxKn
O9C/Sl1EpQciZfTwvWBE08XQg7ITPY984SSLO4QL8yLA//aFUPWQz+eUzzxqrvfB
n/vY3PnGyJ39Lzg7MAr42uuj5ycPAmbWR0Ll5mu1XkVjd48ZGBuIsynPSpqmyLSk
cm5o8qc+K4S0ywfyiJnCEsTV4e/vgRyajtwb61ZMxT7ouwcfCAT3EDHyA7HkddcG
cZ/PEh59gT71pX2JNT5KEfv/k8z/qkD+eVK7XFk9DOvPcLyhEh+RbfyMAkHvvi5d
POkR7du/iuX6+M4UPxxoO0c3BsiIoR9sNEt1IETNldOv3vVwZzhzsmlqIljJuymr
Qna+xNBR+TtgGJ0TjW0XVzZx9cq/0Kkmdjds9nAGNwZvpguPDvKi3MY+KbJ428OM
Te2w1qnVt2O4MmVCjCySBLy6uUO4JOyl8WjHz/C4lNchi4b9N/M5JM+4gTWHFzPY
zALCEbQRMcPJ3QW/dYEq1I/SuyX7TVCTysboHa4NPsRmBJBUsiPXc437X+OQmBk3
JGsRqACLMH6syMQyzME0VpznuxSesl/YV9+yUK/3glEeEciPauCwmq2V1yxAcVp1
d6PVuhUjQsaoG/6JuplIGVho9NgWtOSqioLEZJgfqEYSYgToHbGmhKQifcUcinOo
4nNGJjAJ86QP5etPy8+UT0tvJ4DsrDX3o7zANxMn6O8iPw3KkW+4h6IN2QGXCVLB
B+D32y3U6ojqcCwxklfbtX4Uso+aDbPUyaRVNRX5nuuKVKvK5xCwpoLGvUaZAskx
nwKlGgJMu6TE4jmNSrjGyMrqxvuF7RVfyKmsDEMIHlY1A+4ce8dSRdkOWfUHsNl3
raD3b+fFLh7qXVWGcg4OiEm2apKUwGAWilaIBVvUWeu1jOlZ8VePknqtfQpYak3+
a9mbFhfIO4YUJZ9Vw+eLMXJoyRXyS42uQttziyOhlop9Z+K+5CX/N8tR/rRf1I/H
gUhPt8juVX47OplqGMvGkVF8hnygT1vFFswAMSF8ZOVOY3q8cCMgOxMI5zKEFxE8
vXHxgJqpvSz41i8jlBMOe0dO4L63UCIVvJnN9WC8j6WhGkB9pa/Uka6TIYlB7bcG
kBiWppRQN55cmQx0w5aXcz9gsr+DMraUqAB45OqtEqlqL2vTkZ5pYMsHEJ0FbvUy
9/2zqwy0B0fpMDhh/MQ/tdVPF+I4EC7/x80WNadsGptUbAlxSx58BeTGIVTLzKen
WufqV7IdDmwbxu1HKuvgL/dlW6PsVHYnvx0LB9RQKBpW5aHJNQ1lVAjXUmdOvqFG
5ET2LoxBDJgSMiuLbf5qRdPk9MfpfNvZpgPvhDa5RMdH6zJA6G0l1Xdjx6n/0I1d
u1U5yXmNHykJyfWJ/LxkP8yToHESNrNyPA4RCGFKZ4ItNF1FMuEVKHSqSfUN0wXA
CvuCwxOv+UAwU9yUU2W6sZExBOfxoykT8448dMuJ1jO6X4mnnuE3aqnIh1MAKtxN
Ya+58tfUxOSPHEzQjC2lRENUjhJK41/q12GMMryUFBtsA4K7Ei2QMM3HVH7ksjOS
P+HNFJ2d4kZu8EuDys5paYtxmrO9VhQID2nHLvd7+1DRis+0ZJxJGSCtMShfD7DM
KvZe5TDYQjYwflV2NxQ7g9xZk1ajT5+VMi/vGcAqf4pd6APoU18wldkOuZ68nZ11
CvXfBbQj1YH1LV+sAy5MOcfIROHdLStK37HdynnkvwlXPHw4MXKFc8gxqnhja9QP
lnjZPebPbllL29uBjVXzgZwBxT8eDOGHTfPjWX+yhroizy/iciQaGDvqD/dFK4xj
FFczOYMT/s5VS7a1F3hSLdLzzH3g7TR3uS6AnV47DkgEMKtKAt+dCXpwHwm1fzQ+
dU8qSSQLdEe+JzS5QHk5QdxYjvrz1Fwt4kKyw6G3qrEFt+D/MgW+w8lBtSCKYH5l
bBGx1UiUYLho6GBPajcvU0M7iY/vFCZc1Eaxfx+CTHkkNDon1QZxY6NAmLX9T+om
HOIYHpDNklJJRkWuyC5c+O7xoPCvjHieZt5JG0+ofwSJGz21iaJWFcX/xQVJKDip
A/RIrLGOGQVCHDAHmn/YFZd2sV05uSYN1TgM/Th9wJ6jHF9XF2/EaIvurQainV0K
6IffKVB2CaEysrJ9fDs9I6PmgvGfegA9VUnsTdHVgSkTNKemRpXo/9WWT/1PAJwp
z5NM2BoyV+UvtB60aNfVioFBMtS5htOBFHhMbPJBkyPNcu75iF2QNo0HT4Bjq2Gf
BkGV41PZpjnCf1qQYFc1Q9hBgpzt8Q7InxCO2BWxVqjZ8qXuZRc8t80M+ov4xuxg
R7+JO0UGFzBgzN2sKOGuCPFWs6rfhmlZf0Eo5Dl5IJV3FO0Y1+YFdsA9rhh/nJS1
SB8ibH9GCP/SEZ9v7y+LuOqB3jNbwL+8lAzhec2svyNjn3csOd6je+wMTbOpN2/9
4uXcSFZ9OfyoPw7wMAE2Glmp04lpVUr7+UfD/mCKTvv/T0V/duXKDsMV7LnLhEou
inin5WJXRwZH329bSIuirlDoim44fYKxbXTq7CymPaxC/rD3jrh21kp3ZbogFfx2
1AfnuTzRZJqlbfeAUxdYMlIg/KToDfU3EsUgAaeXbqCaQR15U82Y5h5wxVFQ6ng1
WDSe+Oe0n2VLrlPHWWrT0CRpQ9xZlZvdq3bSrR+D7JqyIdN50Qvo8wvCLnFqwRPf
4OKXDQ/MGNmyw17dInssqdGV5wZIr02k8+jF1Bt4Ry5gAIEsQSZG5gY4HE/VUVQA
5h8RVfhwD3hPy+BdrIZIJvM5FZ3AwEVKQNIn+XfPxR5x48FKJtq5PNlgN4Tgw2Zk
G2HVMEtSPlPVhfoG0c9BWesB5BiQTMXdaUtwwsMQDngHViFUQLow7pNzQVJfDpmf
MWfQaYV0zmGSEYDDQ/vmTKSErRiugKUJTpppC2CRflSziYfZltLAyLy4+BBGvq/n
Gt8EArnIaL31gghUA0V8YhkuG7kAl8SF2LpExFCDenuBkyu1uG16zQWRWyzbixSa
VfY5iZ7jBj5gjvJD9fKSayA6xc5BTRCi6OxcYQJgWsJKIivNlSstrN27UGSZFPLP
S6Qy+TDCxrtRE6iAj6Pny/ilUZrti+50vBLxLvl9GqWn2IrVRQhKb+lidOi5vReZ
NSoUWtiLx/ffobmZgQX9RjTz93RtidK4sge8+k9R7DqR3FGUBiNrAsSiRhH9bYIV
vTGf90H3stvWTX6fe2Wj/y/R3IuVVjT/qNOYunfqlbW/HHELxBOVdng3ohBLv/nE
MnGd6aMiQN4XUQxNU6DT9plqA23RE4UZ11WHQoBHXjxHqUZThuXdbDNmoSctZW/r
NWVegWOxuJF5OI52+/thRXludDO9cdc01P+R8o2VyXfGWYdfXW+uvANzehQ/BY51
baVg7HOuklW8of8HTAK1dQ+HJvl32R7h2hyEL75TQwy+pQlz6NepJlTmvgOEDOsX
u+J/pjyOcYap3vmK7H5GFCsFu5hjr7F7TnO78fcwf6vUVWy6MRRSle7m0Cg4cy7G
QF4zNFhlGltVml/Ff8a6vg7YYvWqW2sN+fyCJ4W/oUUIDVEW27G0MMCaaLDNquM7
aCCvOlfcQ/6L61NtmBiDizcpmYrVEPA4eLEt7fvjCqsLoYdDCMjRC5SISN8FXOuR
HaOMqiCtH0sriYuW+wMu2xEVlAcszRmn1LorKUAdtjSpNxKztlGkf2TJsxTmRl6/
A+bTmqJCRizrF4ka/VOdTDfplUHyeod8FBWcnPAWDUapPKxKQ/g4iIHc12q36sCt
6TrmRUREX61kG1uxJhN+p5y4PLofweYDIcXMIitUXQJgb3i/EpoiogfGIdpe0ALu
+r9vO8ppzKre+anRFqgALFIL18BPwj5JeuFuThHdm0YBv3wzLPOGFjIWMX/SowQN
xeHudw/KgzZpF9GYl8TlDzH+5bdktr3QAe/Fbfwc5o3nZxImlgKDrhqvE2fxgijK
vVcj3dLX1iSG+vw6qkDPTK7NzBuKqoHD5sMLLzESYP5Jqt/fmYZGNn3lKWHSrheg
FNyUnqP9kVNZvgYlDib83ClzQp5qT7I7DjmL+Y+Amxsl3JLNE8mLG48nhDK6tWpy
3r10bIPSrEuHikABjtWQYeutNRsyFq5VtWGMlLaft4E4cDfnSXIE6RE5yFD6eS7q
//6w5BurUzTjgVTIl4xfUybnC/vJzPvN6CczY3iirJbgHHPnqaUGihBJZKR1t3AT
6T5RvwXUXHlo9Q7YPulMKjezndSFOG0dBPGNy5V0IR9Jkcr521+6M2RBpkNMXD5A
U/WhVksRWEsfkh+FFQ62yENGTtuiz+d8Lbhvi9eWiMnZ8AUEbrBhbAXbCMkGfMe+
9d9kWCw9l4nxbEl5FBXkWuhxajajvz4sRUoIjkXjHg+NcaZXObyg+HxXF+Hqe7Rk
wN2Q3yWu/AKf3Z3x6RGw0EATwuVzDoWlNpdpgOduELQTKKoKhiMQpTYcYqhElKEn
D5mqnERo/qoSVoSr5YgT8RTq/k4CQGFZf+MuvWi32YtgZFDGQAPXQ5Aduqt8V+NI
jl9Mvlq7RPbcx31LK3VRXnB2PZhupOraaRAFDMcQ1jt+MdXeWBE4oopLgB7Y6P8w
nhgTBS9wB38Gikgs///kN/nYCLXZHp+jGvAZGGyl7qXe3sWCOluokl5XgowaFU2P
8/nLWMcSKbo9HCu4zCM+dhOopLKwppARA2CD4Am85h2vdKKrtVpfR/DidEp3lYVQ
7YhruJUSsLw71ijxMmQY2/yAO8clW+FHTGS9npLQ6vhKQNjXZP9I/yCGVWsulee9
z+mZ18o7ydK7TjCFOntoCDo04m6pIp053sIjFYNS7fC4g7TYdwRRPujFc3blwyam
secoory0NnpPVdrRMUW9OpLxBGT8MqHhjfM/vipxyjNVVJiOnJW4PcDpQHpM4Hkj
PT8HlgY1twRpAawlFVZz6pq1DH65wp0EQn4o5g+olYzSniCVv0w3RLEuZj5AukBK
6oH/6tX/USzSMoaGNMFAI15PtL+94XQVnjLuKfdOadZKBeVdHfd8931sEazLN7Fu
q68z/QCQNCnuiFgC+CNTmH7sY8Ei5q9uO8Xg+1mBkQNi5tFYkwiMDtlE14mzyPJJ
CBl3xM+gl3iXFzmQNru2GwBVWGeCSvYvOOE2+XeqzXTKuKbMgLxp+b9cUdoaQi8L
tgNuC7Mvv47R7E3Lq0cfD3F/LQv/ccaR3OppnIRBu6nNCJMwChcX4wM8aQUO1XNI
BqbVHC7exrNKgC4NxyITcX2MoUzhzT21NnQSrSV4kKZ6Ijd/D96/3PV2GUmk0YNJ
QHYV2uZWs4HWZFS8A9a30uzXa/bTC8RzkUsXVy3qh9hbDRUn9IclevPAfBosZIDH
1HZqu7sS+QP6KjbBgpoQkLsJeUMmQEopRTmxx3MCPQlFHawMCLAit/N+ib0MQt0m
MvP0WPK1okCSr2s3aXk5iOV254H2UDGPVpbBZ9A0CUfwNB+blPj0kvmDzO7PK1Gy
rnG79mPz3cQXIqLelBLvtESBFKnoFYlczGz74x6IzsKsUZFaX9dO6MoUH0Y7wRmM
M+ykaAd+0jqjL0Pc6nn2WxuShdHRlSHOcIhg0SIDw6kj8q5fCCtFf9qSDxO+4WUk
CGr+oyIoVWLdGlQGesABCYxLT5NqI6QL690ZtlEtr96meHCcED5oRibrF7TMCd9R
YuZbKU+qb6sCbU3TWZ6V1QnvE/XMbNazxP+/FziAYcAqPYzUUczeTS6LJzcSlO5u
haMpr3LFVPaouyGRYyCGw3PaBUdq5kdI4xqcHfAoAM0gyeJvc+8yPH0D42nmHsza
DVtr+irxS4s+OSHcI/j9ws/ACYST7vW0HFc7IfTUW4aFd6IOFI5K+wbVOWvwkKcE
X035blsGEw1O7Zzt80JEUrCW8i+xAF9d7R5cLO2Q0CIN/OyZrtK6MrOzxLrNH8lE
beLsmToyEJjLBwONal0CDdPrVM60UzWrY40Zed7TMBT6Cwm94xSpnUJV249Bmbm8
jwgrZQpHLfCo1MUOFjOTxPmqtbVT/OduuvpQWxr5CXpqdAwPHxW5CasUrnVFA3sA
V0har+OE7LFm/F8uqhPiwo7y4NDKQkcw+2nmErqQ8UBsA2NM7vKq5N6tX9tRE9gR
W64aSmmd04ePFaqch4Nzm0oG+YduI3B3W43PvV/Ysi2PzvVFwhIzlYyA02xePC/p
iw8OovETymW37dqCl4z/LG13Lwr5KMtLry56UZK+L1ChwMJ/eAZ52W73CD3PJQkA
WYCOW8Uh5Aj6m7wRskH/FtAoPVLix3a4l3wsGGqDSmMobetltu9cnGsiiNdMGFwk
5H1l3ej7n07FvUfKS4T9jvYZz89xwNrPXXNb8fvUoBR2xaFMkwBMaSgRLK2fVyv0
KeLYKYIO/VTqHS+cBFV8eQ+bOECprRqdXINH0QgqNkibtvU6Y0v6Rg9dVNL9wJ+i
hKrZRolVuY7S6d1Uw3fHZdL2cmrDKtV5+vf7I91UGABugkARzjtZVVxkrCRarrru
k8FPMLMTS5rlIMhh/SQbU4xVrnqKWOmMeJWos0Nz5Fd4K452EfCxw+ziDyDx+JLM
2fSUbJyNo7tTfHMdXdWBH436U4xx7nyVc//8y8hr7ttp6PFyfLsLpZNLiaLBbCCM
lmEso4KOOeFFlaIuf+/jjmzVN9ZrvpT8nXO9cFXQmxEeOX0JfCXPL2PBa2nH7SkA
KVU2GWzjTF7g090ejR2t/sk0xwCedKtvWyvR9oLWNOrPU+JfVHLsDxKmQRKfPQhD
tww+WBK785ScyUU+NniByDi0p0pGHXiRButrmGI3pAkxLimNEkdmu6q8NC6ppkIc
xSLxj/5/q5coWhDh6ZgN8uB6gF76wSL5LLghicepGcHd91VGnwFkSEPGlYKNa6PJ
PzCZG6vjT9LB7kHgdTN7DxodiDCnCgW2Z9zLiKe2//mvYYpIQEW1PDJuQ44S6NHQ
IxN5Zpq5dlgkB1AnROKrpg==
`protect END_PROTECTED
