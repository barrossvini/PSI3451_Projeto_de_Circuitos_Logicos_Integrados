`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eL9tUU7kzj2Be5OM/XRJ+X0bLgicygI/F8ghor9PNxkeyagoAnzMYRiKW6TMgM1q
onTh2b0jk2RCMuyGYIlqNBnbHvSyoSJl2MmNYEcZY0q2oHIbITZ/Y30hfMOql95A
DZewH3HfycICG1u6JxIamyjy0sMAZQ2PVtYeUjdvpuLLxFhvmje3A416wRzgUGzQ
yfrq3vaBHlEWU4dhR5W3To8XxXgJ0cOmSyZGCSSfqc460FPSCXrCBLMI1tj85T7E
zTScBm20yoZf5l0iSPeRXHpDvbRhyfaLyvE658e+MQyoShewxVyXs33zwTh+OJnl
RplNOWaXOJ5Rh63MAp9VccidRVOIE1uJFy1/fflHrSZfgBgFMG4b2R6cxoBxuZdW
O3ZSH1tzRRJGPvr9ZZYkJWnqbMG2WaV0h8gnNT3t9Gc1AGmh5okiAYiEI2XEMx2U
cuirRvS2SpYA7V5cBOh2fCOew7sZrOC7f3hs9sZoT3TgHkRpUK5YyJlLMW7d3H91
jOcy8sqIODr2GYNEVsS/UyrZHyuRds5tNSmALSRIrw0wU5KKmZ7GdY/coVKBWw+B
cph7MrQEeChKIiz+x+FMNa41CuXRIkah47TYW+PtnHNpn8xQU0cwiBFI0XcwXmK6
i3clS43r0LT5X4im7r4Z/Adbt16DHOXdAQiSUbRgnzOMUtADGD4I/R+edfrtYw+t
nTymMJyIUAzamHMaKfsFrgPA+NGUTTiZ87ypv+CFLu3QXe3kA1PlPeVu2gl+n1Zn
uERD4wmSWfjA5+45qCYlCl/zw7E90Fr4qb2s/bd2Hd9JXFLjwzOnyX8avxiEW514
QFdaB8yItOR/RNZU5/xMSdkUTdh1rK8lJh12sSE/atDQoKTf98387GJh6C70BCno
BrOKXNL00cl/zzOle+rV0+M7Ry9NdP31K6lNR+LGD0zd7Ha8G1H9CnxObNuIFrHk
5OeO0Jg5mMul0o72lNndwe4qd/dSutgj3pRrUpXyjvxrUSkBGvT8EZyqo5uuYwuB
7QMtb3fa6o+FfvFw/Y9B25pIK6BYqbYCZwOOj5rZHyasyyTdxT/Fa9oM7IfehsSX
E0SDsrS9V0Wj4cYTpTk/UdDnAG7nyyXTt6pDL+SpvradQmMvbQP4fpEZrqJbQQIa
7FsZcIjtIfc3Q+BtFBbwk+4sTSUruUDNOumteqOaVP0H2QBcf8E4iSNxv/GmFalE
QD+7HkSr7H03T3KDlU7tXt+RJh2xUdNmVS/Q9nDsW17efbL2LpP7j9WLUqIN1dEp
VBendS31X/JSM0ZZ7lrJQhD2BNLkszleFEQ/uGQmujDJ6oWsjbmPvA0txFt2EZeL
rU6Lol8/Y+aB1GiQqFf4wRpUpMhXzn2k/vmvntHOyQH4WlsFRrSjJMM/MAC5Jpbf
RcqS8M6s0MOyyCfnyv8f/3Eu0hq6JyqqHmBNPy+xQDBv9pjCw0WCWF4T4UImEnT/
ZPpGBQMFSUHwWLQ3UKpkTIl3ZnmLnnWMH9di0P+4CLQmVuFBs+x5VRy4eeg3wYz6
sqzWSq9QYSc9pHulkxA1kMJx0KGxvZFUX45lJJ+WSca2Fz5c5X7EZzfPPVWVkekA
SXq9dcjrjs5mmoHF+yqzHRx87kcRn/ZNdiHg+z5FHPYW41oXfoXWPYpSqdWqciFZ
rnPag0AKGjW200f+iLMMYGX7jn2X6bNvsnjhObyX5rmUU5fDYXDYkHcVa+GJ+hcw
`protect END_PROTECTED
