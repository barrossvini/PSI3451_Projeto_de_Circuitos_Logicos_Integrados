`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S3Nx0VwD65diaa2o631NrLqBfVfypLtLMk/EqW82rNUYGHz9AKN3NH/hUXx5kDJ6
V+QEXHvNN9WPY+S3/fJyjupv2SkhyV9vsh6GcAl2jsBkQjfXZGjyMrdS2u4Mls3c
B7uk2KtWQK0U9/7+8ybX+GBcIzAZFzoYVoMruw5J5mv2P9A5oUaM8STSzysh+uan
iqECDBKJSslcueuY0pxLQ2MQv30ZkmbMgnYMe/B1MvOp2T4ZmJHwhFNqFCauLwhl
KUFUr6v9kgZc0/e2ZXC3+3aRvtOBI6HmRS+yT6xa1RZEq4cbPQqLeNNXVSEZGtTw
LaChi9WJc3Lv3no+wLAKbu2bGJYGRCMmAtumaNQGixTcWw47lid0Wy8WD5f/jIQ5
qgjQD1Lxw8ohW/cXV0KK/HfuA7q6euSbRHZx5RJ4gEsPeICqmlqfFCYQNST/0Lkv
LRfCZOwvDwrBYFI8I1U+uTuSI79CjyfbCckIWNZud070UC5Ic5S9PKGl/HZa51Ah
qa+gFxdM67Ldkv5ZQ/eiCFRo6xHsf+wfr50VYJb2tmlJPMz3zyuhEkh+KnZFGs/B
OlgntEdjZUxnfTg9+fQgdkBQLe09rPAVROywTbSgZl8UIVD/lx5FPxVsCbURdHEy
Q3oVN8/ubkEoOMjjN5rJjpASudjCpufJ1PyVeuxkmM9Z666ZHzkXI0v5n1gFt0tp
Zu4tIW2DNkXQDkDrv6rzz8ZHHKRHQ1iSfWSOBGZwXpzFfTLh5ASbxgxe25iT4qj2
9+7vMGX3zfNZxeQ+QNvV6srRwtt4ZcU7S2R8f1va3y+VDzzGwT5p6gvQTxrYKyJp
5e7ZQzO5KjFEfZtwK6HbNEA40bVDVTQoUlhYMemfdUVdZvfmMkU7FJtBVE+oG/KU
VKZ5Xp7VDXRbDVfcSBvNrU8QzFMRj2mEwpChzI/KngvFM0CZPkMYDbEQj8F/hYrT
J8EqcQNnX1dYA50oai9CjyN2rHS5NQKoPst6o57TvksvwR1IefqWvGwGJ6RZ6jYc
3dyly3/HeOi+f7cHqFBucv1wiq+1vuLUeQ3zg2SJKe4uZred3BArMCrdNe5ikbXg
nr7QKXQ5Eq3SyIocEq532BJGRmfwUhONAV3mVsGqA0Eq6tpSRD/lWL33sV2DtqW3
ivd6va2AaxDwgGBE8TghVApvmV5HKfSoxYgSS1rLPxvFwKvU2Pmdh503JQQSZ77F
Gn0Ro29E5hWJygotwsyousdOEkvGmG0HepLY+CdVds44rF+25xDCAJoZhzxMwK2e
g3YrWl8BdFf//e0Km4ra+WX507a/ld9URCNmjeKZEDca5SCz4aQ+P61D9+77bKmt
c1rpaPxb4hVyLzpL0l6v0BSZmhL2Sn5q54H3G/eQNFUGrmpmz7OshB1pkT95x8O6
rl9IpX+yXqoGHg9XVhIESfQk6bGM7YNbeN/2tDB2pgRxxE9utuFopTHB+t1K52uc
tfEGW0KSN2wCYhn1oS9PW91rNOtI/r9oKo9QM6Cgw5CYL1F11dKRhxYwrJ2IMS9K
Y8TwMVJfflbG1wTYDVIEAtv/ZYjRqp9db/DMgY7fO1FsEIFFTSoMjDrETaokfEWx
58OvoWLrN5fkzro7V8M6ph1jpsQC5ZN+cEAh/D1aRTglkYPumjn3ag00LbFQNv37
BDstVL5MSMWZigfLkiOMGtmlna4CtBGDEV4yA4F33UW3AfFbzcfz/U3ctneW8Mqq
j+H9pOlBKHOvmKqITHCBqGErhqOcvgtAJDl8k654CK1mZw3PnvAkpeZL5V353fB7
iaJCHrdhFY0oJU9ZilHYxIkdtsc4NIhjjWPSw+yeKDl7eGpkiuiXLqErQKnf60Zx
Ljubv+IrRVi6ZAAnIflKEzv5bsgdMCKzNLzQCEAc3ef6hfcj7qVrsFofQFvaaH2x
019J5S679GM1mc2Qc90idvzfOIVB2awmmHxrFFTxv79lWJURn2X7GLAlxcC6TEXT
BRExUOio6mJodPnCi+KdSws85B2JY2WwARPNWuRlN0B/6fW8ouQjyc6ZWV22biBr
C0s/h6E06DqTOn2cYUdQcVi2CJIw+he/wxc20w6QqtivP5lnE7kXICp7CEc2qYIL
0Fy+P0/LWMctxQY3cxHCv8KHpGbmwLsDmugkGClg4ChrtEDY26eEOP2P6uqoZ8yT
gZSw3k/OIW7CcWjU1Ivf+uZyNnObioZ86NhQZiVaGgQq7B4kGZhadd31/BA3Ny2z
4B2AyS4VQj1A0zsRBfAmdakOKuNluS/MYENePiDeZ4spMT+8GFkeG0YCkjaqMCao
VQJh+5QEru7zJmYON8OaJwjwMxCTow7uvKXyK3JEfCDzOWm6dA3OJKcFUuDXhC7M
BTUxHgWOr0PcHnvmI5ryeW3IfkvQa+Bm9oSRhqMQt2DPWNQDTeNnnVGv3f8btVKW
dO65m0FrlrrMhYSEyBA/tWEhKldZj9w27rDQLVag+6gj7l6N61i5gdAC55/CpCt3
gpBaMtinuFCeYpT776Mwy8VBJdppmJPRd8mh8IXr6liYBLWot+kFSTUjIYwqO5Nx
EyNbmCFXorlf9eol1N3AUSQT2xibSiMR76ANGpddvEAqQ91oOA2EF4ZZ60khu+Q5
+aYLFxsrB1B8WZNGlyhb8NCw1Ni1VCWl2uFVIoxLSQew7UfEUBnjEden07t1H+i5
DSorsXEaSXmNfXJYlIJYpOQafu2nqYwyMjs4/iflU2U3NKsXy8dNvHJclrVep7Xp
lTK56V46rnUJg5kodLRHsRRZIobTxkWl7Gk6D6f7hJW8VfzA13nAIADVjN2GBC76
P8GJ1b/O540mhBJdoUTrhEBlNebsju8eJuKk6e4t73IjQkOiYT8p8cz0hXOcIQJX
tH44FScrhMOUDdNiyg0qwZenWo7NA3vsR8Ljs7aP5u2+s9JFyyNg3QmvGsYSaYIa
hCATDO0v9xuQXQj1o45WzdBtm9PTvEDU37fD6/jtfSaKlSvRJPzi5y5wpwqmjx3/
02uwECvXlgD7gZpYO/3DC3i/YmJoRodIgfLrzxWh7/tI61oc/HmzL/LPbSBiGyni
5YgO4yS9MjE7Cr6x/tV/aybjlYQAz5kRuwfo1HddqQenFo+Mp0Svkpdd5yQqRu6C
mzc7phAzj6sY8qdGEh80QTQnVpdlDa+FS/GIzfpUIDCguVJE0zVNRmsHOEik03AZ
Q0Klb4u5J/Dw6bcmtLYP2okLQ95S19HC4fl51yzWF4kCcUeKruJ83+IleEv9o6r5
nJNhStYn4MOvtI47PWIqWg==
`protect END_PROTECTED
