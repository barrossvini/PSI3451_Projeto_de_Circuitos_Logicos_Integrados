`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mSyFob7cYH0pNStaDDow7rC5E0Ld6zOAj1IQ3/bKwUVOKfZ4Lxci0q/CGPonfKrw
LSHuC21CJ49q2KU5LziG7wQRK4JtCC6T2ZmXwWN0MeMoHWegeoifeOevePIrJzuf
qnocgeHHPuI5Vd0hzoTMQS5v/Cyl7IsI3yA2PxTYv5U9oC1xgTrrAJKZLHUvoReo
Odf/3msv8FCberKqhZi3/yWS0N+GGQouQMdLvrbG0Vg5iroVnJOEdoa0rs5OVse4
DZ9k0GhO7acEe7ZXX2SSd6p3dOJuOJ1tJcLmXlz7sDrqerV9vfjAd9VgGHRSevFz
spHJcXFP6NLd7Lfg/mJDvEucegTYPPUgmwRkDP0bJgHKaR18xPj6kYnLoRh/N7gB
sbrr/HI6OBfQs2noWUOHLCW2cUeB1qRXpQZ+gY01ehkv/k6ZSglphSGgJAVeYErN
1fAmy6Dn1N7kIeEJ/6xsxZM5jhuszUvH83eFCr11Aiuiw0NOB2gO0TPkbWIGxYGB
0YCcaI0qxdCiT+qmVM+xAgqVbkTYW+rit75TveE33lc7CG9xzMbDS0rZetFd2Dan
6hFgWiF3QExQp7G2Y7Es1ta5WR8xEqYk3yHuOGuWF6mh7gw+Gubor7Xo2+B99uYC
lL1x04GXQQ/52QPx32UEx9paiOXEdGOj487T111Oxj8MnkAxC1z2tjJe0MDVXRVH
aZL9kz/iBOg08EBUv0FgPUud2gZseaBfrIiEslmCSJh/FKxWzz6a5oP+9H6ls3Sz
LssZMlCswCsGVyVwSOWSp6OnZruZWU1eeMw0QGyG4Zc1y86qCr7q/UHsUNV3jjdY
A/gI4BZ2tNa8fgEnWUMPO4v+UlhKpEMaS0WbrtV1UwkKh2+wlFe+HSCb06crvmZd
iH4/u6WjvfJo4zPGoYeeqmfF2OrcKfq9Z4EWcE6rpLc11ZV73V2tmLs+TGNzKDh7
EC0Wl2wiDb02IupBXKi4L917eScMxzFqZJiGMUCid3SEY7LvYG0ztHsAV1Zlig5t
JDay8DWj7YX/0GCsWd0M6A==
`protect END_PROTECTED
