`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h27V79iMdGPSig4CazI+j4xGRGSXS4mg3nh7X9O1hwai0i3Q7PkgMMOUGLN/KCN7
yAeQA7AzmFOVP8a1TAe+/nyXeyJoidNLlCHn9XW1CYX7OKVCCP42YEvJUQnwACXm
DPsXhlyauU9DABQdd9KFqR0lmD/fU3BObXjh20J/UJJFrDjGRzCIcxAeIiZYxNbZ
t0tuj5OT9YKL9o+F1KTZczvWyvEDynV64lO8VtPcBX53Mzg8gZoRAaIhUVKULOP5
EqJbrVidrSHGxHmk19LilxKnQ0RlV9DlXfv/MGQMf1TMiUEEEKERrTNILq8dk+bg
kZvd+W0Ax0uobRog/nuUS55ObgLWqpg+qy8PmhC4pejNTDn3B0/9DxiyuDOl8R56
N1M3hFqbmwY4YEetetTs4tyKNSNTSQ+bgJELsDdoz0EMPSCCHHkWm42zrS2Ww8Hj
Rv3UinyXJKoIEju1do9FGE+PYuYic/i057/Yfnt0tvIav0u9H4VqOcuxKVfD12Jo
4GhkUhkgKNzioIXi8rxIw1W2xe1yfoGZEHxBes7lt5fo4yXdctJAhnf/+nV3Nz+l
ql+sMs5GoSv44Fqy+6UQH0ldLUSjV8QoBsxJUZ8O2U7/Eg5s7l0a9iPNDX7fCQf0
U1O0NK5ADY1zljCB8vmk+9u+6OkYkXedxDKmJxxLnVAMVDHptI5HamC7wLDkQP/J
2CHtRniKXDg5qpiL1ZUYYntNQxjvbR0eJUZtCJIdcSYRwpTyGX/NDfzU22GNKubz
UHoylFhKSRwjUBbnRBiiPqwGxx6TSOjp9LhjAqqT4jEFfGNqh663whNUUh9OEWzq
n2KoeWAcuZQ6bvT8C5sr+TfgkY+4f7/VVwj7dXpCgMqpN/B0Pr1dttpEZz7OQnlq
BoUHGWCvKNzUe2ald1aBZ/9ferbZLmRiUyoAidCDhQZGHwOCPk2OW7CQRnjO9CW2
vNWM+g5tE2HQQEsdisk2GGsHTz99lsb5e80fDy3JzwVJRwWdaSpyuVyCzbgUuRK0
myk3Lj3jSkJvXFd68x4kGvJ0h10S4SS3gofeX5h1xS5OggGq6f0HMVq60M3zLOwy
rmjpPP9Yc1pEZ8eNXeNLdvHbLWGte+RE+xdk2c2paTOQqzoFU3AamjgxcgQHj3mU
z1r3rknjY2bzLh6mMkI7i5eTzQPbu5xqaUmMbl2hyXdS4cHDaVP5gWRYWHfZxefi
o0j+trTTJ2WyXBc6gIUcX4342u0a/eltyU2wne1gL4Sb63oYwodj0+cdhmda412U
VDGAAGrx2GYx25ZlTYM0JgxMjhaRgmN2IABHxl3VbOSkZzDFqII8EMqz63tPvJJ7
2HcJfKlP4VcvSVv+bpufSVkYY65p+Phi0b8HWLFCYK3ALtKJlCAijcSf4nhC75T5
hiBGGHEvoJIWFYT7K/YVUQ28UCy+RjrjzzwK1djdO2Ntj03DRCkaqt060DNYXYt9
2oWacv/Yfj8UaHmwPbkkn1ipJF9nQWYWD2qfD39TLrRZ1OwObchv8HYOz8kbEafg
rXGrTREgePX8miv48aT6gR67TUqJYH0QLYFHkjeqbR9WITFYsfQYTMFHGD/MNS2q
uu3A5V4hpypLIqbHtdGmzJNwpa3vPB76P5kBzLRfIZHFY6DeCeqSdOsjPLW14bgL
sPkENougi4PspD829/7Oiz1ieUqLgm+pBSmUb/r3JUE9VP3NwiY5La5jtDpsrDBe
T4TXwsQHnt9BA0gWQsoauBoNkp2LX3Ou7u7KM7DKTkBpfEuQbiGZ3kSTqSMF2TuA
a1swppi0KrKevgzDaEGN4fnXUShmy0dreuZVfrGKCy9f18pgsN1gGYk43vRMbM3a
7ZA6l6xqVL6iewLlTJg9FAQiuB2O8cXAQP2C8OMZyThtpX+gkw3jAnqNJ3XZDXI7
tY1ZWcNuLqwSjp5mRuAYZrIYUJe8g4cNQFCyHHGw1PqSkU7fTPeeT5Me/0mvjNZ7
TuxY3D7GCFpkJ8aTUJTty/WpRE3JYJCHRdt+t0SCGZlUhhyEG8h4lG1gEAZNgQDw
8VKMMi9T84lo5kGIoI1ot8Wh6Pb5zXEJiyW4Pt/M3n5hMfic6hsUVmRRtfUyt+g3
vKuHEJMo0UM5L/1tanMQvIARFfqpoErwBJoil2SPW+MnGtChJyw7k6YkIdXGp+hT
QjNlRJHvBAVfgrM4R+lAvGjwp4jWu64gqlqdOM6jH9mJGLsolprPA+vF2wBimk4l
9wptngtdqHtNK3I4aVASXnGPYhVLUhQ3Fk7V3TImh7ttOyWJndPs0+G803XXlgWY
1rA14I3KOU0jlOgXkRgh+B5Mv08J4wsZoQnIklNa1UwDDjCQCY9Wpc2JvnZXipca
DzyHqW7UYePFOpupMciMmtz9aUXf9SuWLvLnebxxHfi9vsGhC4iGIbZ8at/jv3Ig
37gCf5+mHPzoH9ps5fA1X8xt1UqCjsE8Ev8CEOYwuGgOOHHUWZAVf+R2MR1iy8SG
ZRgyjAmSwObA+DMgwFMYEGL/KhJbRC2iwZnnASck3yjeInOJ37iJ6W/O2Mb4XBKk
aCTvDB19DuVgRo88jYNpVozeIV3jcs8KMCMT6fRvYEbvYOTbL4K7DQyDqfdz3sVK
pIWdNKSMrTfAW677xUyhjOhrBwwB83w/Ss2szNjWP/UO7QU04K2jLxTmRwFPIlkU
+Gkdi/jlOur+GZJrDKnNaimusdJyVxVGwRRuBUXBBtlP33gqEUzqUDgCYbFyyxhD
BhzhcLbDucSY78qxhW0lFecp75xNmtuQaBgTi05Xwlz5YQJ+mK4jgsRubgYT/ju7
4rYhc7iheiEyn2hK8hPNkPYA20BxwPvBlXEVa1UGJMzVzrrABMOU75TtgeaqD3gk
phAir7UMOvyAGZE+YHWXXVzO2GFfiwjsV1q8XLiCOclQ7DjD7JeiIg3n/g7/yGgL
yYHgL3M55u5Tkk+BMO82MxEIavj4xDcfhQ9AcGq1/RObhb6Mdm3bBH6Lm3CIRdQJ
MyEOCD96Ng+fvdALYqum4oWKI7FEMOcfT37NIp6IWzId69F6e4d2vyVWOgCa2O1o
I7XGYmKfseE043UN1YCST/KQrGwaZxiTiZTz9AXuuJdM6zSpxopWgF1G88EBQats
IedP/gEcxv6BxHxOruShdT3nf/rkjukVPTPH5TaWGZuRkXGhnplYxuYTp2v5jRMT
2Amqf7qUJFM113bRAGDRgNZ7j1ppnJPZvil2I5w+tNVcGQhK5+UaT/uIZ2+rvaTG
zOB5mGxsf1wHyHBO3p07J6UgDszD5o3lN6lAFC8ZNDgzZqAVotZVw9BgSHqOYnrC
SnIh9tG33t2q4UsAaBcA6HvMsC/tr/DIjMD2izM34BVBEPcFTDZKXiYjShQlQSdG
f1W0XKTIjRDFAEyNsvMjSSjiX+f6u5maa9Xu+GEAyxpdkQFPsyKbqSFwXuf9cdr0
CZyiKLhsXK7mvRgtLDUKm4GiRlj2Yk3U2DKaJJmeEZg15BRZzWCXs5V8NqQ4Scxl
wTUCFU3LJ9oLxsHkWjNYGn4BB0lVAS3yZWCBrLnBnYy7IgyXbC85WWE0S7tfPdCu
W5A/cmcZwhpnaWlbixGlBIqb9Fi+27LlYg9E1ReDIEYtAlqzo0lnCNX2wjnXrPmY
1CGcjtIzYT2VgDN0+wCpggZNu/fo2bTaAr/cglhPZWkZGYmV4WyB18GQIj52CS6X
KlO+7X5KqIfYtu6FWDJGh/HqYfMnZcdUWnOGHMs5NfT6KD1BA+zXkfxwKLCiLW98
78X96bIG83nHxqkE/kHHz5eRXEp+qkQHTm8bAkMZIjP1MGexJyD+YSTwXsYwQZa6
PQULv2uBhDLNyhqAj0/XxrVDKiuTG0ZJv+X2oufBNJvsHk5IRyY3buiDXR/5HyBy
W3o4GoK+edPtfa/SHma5+HvkSpM6tR8YvPeVD1xDhSzuc8L1nFqrsaq4tQygA7F0
2kdA4QVy2LPAdySjIz7IJalz62WIscNDrsExFt7UR4CiIBf8+Fq/d5MBchYTHNZe
tMOH/Uv+LzUWp0+Z4H4jKmSoj0GYIZAMQVPlHa/JDVxlYDFknFUxgivzv4PF0N+P
6XtEIsg6a6GLQRrzb2i9PTmYc1Gn51OWT9iavjo3tZQ0256SrO7Dq0zzq9XqbXET
ZcR72wthjHzBs8xfH08FXx4OPDfZGNpok57kdt5HHbutUWzs6XxvmJpLiYhaaByU
NxmLEsng8b4z/imaR1gDg6G1A4kKJj9drStRAcmLQWHHpjmElGJvRkSu3BXv+OVn
n4oFhOST6JQjE94J66aRtpGjrCzM/OZTeuAjEu0gmI838Yr9uXo19j7DDBlJlFMO
UbfLEVlOpVXNpLAdfLSJp3cA3goBaMWtOvQljZjjIw31Tn7oWgaJoIs8dbX4xWOu
VxHft7Z0MMWg7EpuZjBgOppqJaOXGICCj/PkPeQe7GYorlPT1LMa8yY4wD/Tt/KE
4PB3HmFkXgdpHnj7OUz7NDxEvRKnbsyEqw7VfRNmUny4VTRrjT8vOg2hLHJATQe7
Qx4sxW+toGnkp2E/34kXwTaXxu9H0NT+aajvHfdSEMQJPzGn8cpzZOVrU5uHk2yu
+0U1g8GZpYpi7bQ8AVZ2B00LzpfEOlhyhNhthSqHa8IKq3sIfK7jZKWdyN2G4fpv
1jGGduhK6hjMKvLCAqslEBl07/swi0D93U+3wbdWZZEbCKX3+KlPOi4QUT64iOxS
RWO7r5mxrYlJl9oW2UybDkpLMbSJSKXiObdmes+fPMmtLP7T2Wl+/QRNs62wHlbt
fm3slrAX7oWrPS4KzO0YUlObQfhhQQko56h6KmgvVeAHWT5bNv/SlbNGl3hrDsok
9Q4Hj6ocGof7LnVlWcxWZ/olV72FlqifGIyzVJizr7n/aZ+s+0o0tdgeFY/cCyRt
pPNXBIlOJXE0aSLYF1SE+j0U6FnNgi3H3inSranFeZvK7eCbLxdarjKBrPAVFZb2
Jf2Ny+snFcFm8HvUVyHH6TAmsALIMBwT+OYMWHIyFdvQQYxYZEmFBASY0HU8s3mf
99wJ0nTaf2NCw+XsKL19f5zUnxjeFtjhZ8YM+GtP1tLoRgXd4DsOwOHD4zf1dyk4
5xMq27DKkFQvH4obLLImISqapOuSqvJ8eYycK4E0/pqur8swxva1bC6K2vuGUiHE
PBW0XOzNMaF8nvh8vH7+94ZIZL5HksTdZoL9QyglysICJVt4SgDkhMq21w9A349E
FUI1OroMYevN8OlR41z1n9b6YMhp0LcDTAV6L5GWCwKslrEHgSExWbPg4zFk4P1/
WbLbNf5yuXXi/xk1vDINae8nyoERh3c9sWKjpydriBDVX02ROWE2IJ07TtqM9XsQ
qeYV9Eh5Zsl8rE2gWqg6aUEfpMgJFV04RwIbVp5/FUnxpUCBfDuB9QYgwnqgpPia
JVmPZRhTwKgSunS0k9w3V64wLUi1a6qrkv6vhXwjDQoMUncQfGIOd4UjKZyuQw+/
KJUSo6I2GxLIyvky6SUzCcL+dpjPVqN5KQmr6NIIvSknuiSKH/gqGSHHceEGSILR
7KiKYV42Qk/FLUU+hxFrOvEemuQ33+BwptrjBx8QMvbTwomaQjxifFVAj1Mh4/jl
poXZtDSA2YszroBsXR6HGxHeugwtZA3QiS5N6yNqRC3/2/6VI+YQtCrZRwYsrrUl
cEC9gwc93CHA6Iyo2+gf+w/Owjn+YKmciegU0O5xVj0q5nk2RPpemfuW42asdHza
Piu7KnFn1hEYtUHjOLXvdtm2u3ZkWa7PdYpYH1tOq1YAMUWc+4YrcgPEraq4PMBY
TtvAobD7swKpc0aB7IM3EQ83+n+s8Cy78jL+ujkiP3UHjwPWHTpJb7uyQ5Xy3UWA
JFFjwoCFnymBz3YXoWz3SdNSI1NizOnJ0aCynR3gFsNS9TAPxbcqhxvvRSJoIvur
sL93g65T497kirx7EonB4aocI2P4ZJedUbSMy7PO11EFkIJYi/6rBMfnzS0Jttaz
O5HkHq98zcDNlMf3GHfHutve9zRWWiJS4XdK8R682Ff+xiqxOtpjHda1g+3Ijwg/
z9IaDXpUGip4lb1dRNArMPdo7WH9lkpY2hfVEVDIHZtcDqH6veqfaG5bX8wLI9NW
Q9hHkJO4NtzTYNwN/BCV6vZENN9wj62xtHV/3+WxkD9oSH2YnzslGHItAeLmcAfB
X+wxTFDcd2z3kHVn4559+F5Ilv5wYLzTlC5xsIrDx5VXvjHoKhfzQ9UDTiG84V+F
7JTmPJjUU0mepCV/J0pekX1Omz5XrU7cNcEgIM2NQdPS6oBcahJrV/CLlGOAuULp
ykhC2OseeyauT369V1O8TKjyOrmJX1DYHBil3+lYlXLcqqkUZaSwMqvLwvNuNNQt
MpiO+tnogRm4ej+pwbpO3Ix0F3EcROsG3xXmKTjaBWUWgFiUwy0E5HEpZDn7sZWZ
paOhB8FY9suWN9QT0cEYGz9k87g22WBEh/I/cqo3xQHabF837b8mDjEQIlCymr37
8+sl0OQnj95GU5zZDAsoubv8fSakAeZ58QTX4H5Cmz4b1wsV8aq361jHuYSYI1Rj
wmOFI4WFu94GbmDBuJ0RrGN8HQC3/71w9h4wtFIYpoanJZeiZ6bSBr29ue+2akUr
L8wyoRCgQirAguoPXgGgz48qlSOLM7YS4qVpGR0QZdE5a3eYA30wvcY9tx8o5U07
5Hd2oPoM7V53n7MfgkRbAAwq/j9GCt3b4mttwBnQZRrny/Ixc7BrUaP1A20zi5E2
qQ7smWMif9vWaM7Kk9kuQONAt26nWRXn9JlUvk8jcblU7ZL1dpmn1TZ47Uj6Nb5F
n+XKTFBw+/hgBLDfVzW+aXfzqeJn0IwfkFFfXjXicNuJPq4gFzK6+uYay6HJAYki
J9aipnoNZ1Tq1jm31MwBcRTOB2i6d6qr/YOIio+3QhWOLrCOYy+f609Q7ITYctD6
yLYC+8acBJzQCtFWwYFF3rCEyEpWNA8xp8eWAfh3TxAfOBmWRzrtq2dOaXlpqpnR
vPohCFgg7kchHFQEvTRsEfwX2n83eMiitn3ILGSNhyojpBvNCsDs6ENsZhnbwdwo
huNmBUQwn5COnDVdYiPV3N5B6cjc5RFH4V3J0wzXZrweQHlWh+fRPGDFGNufJSo6
AOXCcUIuciy4Mymj4q4qbOB8sytnT1FYt1OP04bECko7PlR2D7urIjIG0LgchUnD
8x23gGscvbRE/QtsWw5wb3ksKoDETfa59/fMHfPgwkxmvV4bQtfAts+73MwbjzqG
3q5wwPEYJwdPyreQkivnXCVdqcTt8kAZM9+1UUDiuyPC04v/Ly6/OUqIra5SYUMq
vCJ/W/Ym+ITP/znWu6CGShS3LPdCh9Pmt2to2e3JgN5T+Q8CINDKPiGCXTIM1vLH
RhltBlNBndD76Sa19LaMw//+0CbY2I2B3O7jO8CKXG/almJTY2391TiSwcSp3JJn
zMjI2EX64L9pnW+NJLlbfAGNYEE6J0MaDjqR+e+8aBT7ZKE2tTl4NoRSpcS3cRp6
fITuPl34Fd9nbq4lNuWKo6CvEXraTNjYjgin0tBkP/k266oKc52A4ElQP7ISd1Tp
H2D6zhy6dUW06sfWRyR21xOvrScOBnytL6Gl3wUQeRI0jL4fQLOOnwF0UzrZeBhG
Ow+cwnG6pXoe3BhAY3Ln6xYNTuASEnGW4hmhJZYmpzmTOjsWJxgz9IWuNzrM5ZXQ
QrgXTu63XsErMJQ4jOVg8Paa1f74n9wXA1GRKGjqSvDPrWGh5v4cDG/9mLRULnYV
gJG1drPgL3OJQVMaRaxpVBLlcd5fLua8zOfurk1DLdR/CMOshcQXACsAz/KZOT+O
0q5bl/ecR5sNY8HTLUR9iA9jreh1NSO6+0C8FNiskmD7OyFGDZTAEnE4BcLsocA9
vTKJnGsJAbV2jYwuIy7QR5JsFRmaN/myRLjwyoJgkQLcm5/pGUlDNWyz8Hmj3zZ1
lIiSL7qTYXIKXEJ7rFf8Kechcg65xA9+vtKSqCJyADqXjwWyrXedaiMKqsBvviWy
KLXFB8B67fsjRy/JHg5mfgyo7xEsSSce1B12hbWz8Q2vji/VzC2bHty3IZ4OhsyO
4M7rHI+zYxPQq1SuO3WJWnEH7fT3l+hGYcCK8owX+XIU2KxJU4egUaO5bJS891Sm
eNohJQxGprHmLm9h2r5HDzVpQK1y1JENDx31axJfxrrhath7rn/DrqFruF4wawqe
kWZPLncT8usqfMvbxyDeoZ0z38olJjhZaXNInoLjt4e8aBGScUtxur7knM7IT1Jm
Yq9ay6DXPsZ01pIrqRJwGP17/DWfPhwJmv0YygIOgYS8VXzC0pcISEW5yUprTXZG
8jFlsq5Ok9LeSaUOh8VyTF13cGYRu9E89VHkkw+e8Mpt8Ij3pXN+nPhkU3pYbb55
vJVGNnPQpGPSWlgKpDBOtvkB5Z1GmFAVOa968/kZ5Dulr8M415bZ8rPT3meyA5ZH
09htF+gMHkT+PAhMOBMQsddYhqKYA3q9lStwo84zQZzT8pgjMN2MnPq8EWyeaIC9
n7dxPbvC+rj/JrFDum5AqUnoWKo+iFSdjKbaob9MGd+c4kDot5gGMpoBCAOJF/HN
R6D0jDLLTz7f09k/RujOaQdtylq4vogz6tlcU8cGlu0T/tv37x0M7EH4SU6T7AkZ
k+7giZWs4eH9G6VSH6bV8CwEThc2stcNFL4DFwRuriPJqixKSj040/citHLGJZ1t
MNf02MwCpAVtpYeC3tn9TK0i1MGVto0tjduiuRI75Tu4uHJ6FXAQ20ZguoFNE1bY
HlNnJZeSpNbV6qnxjAVyNUAa/KJMu7pQPFreYprWCaJNf5SlEUU6elBZj8EzXkOE
fW0Eohv7ZXXcKJZ//j/Aw24wf/Usi5gyMJdVKjbql7nMacnSXSawwITsOAkAsp+d
CbM4LJp7N3s0GZZ9KLS6cHvkBguxKpKR5593GX/8/adC0WQNmSulzl/2zt+tn55m
+aRXybngwPOUTSGNL/bKiCpve9TAgMlCkggVo0x079BcA6atd1YGnQNqnKPPGNk0
t0EBOvU1GUpIZPY5N5Pf0/KC+rvm1eS4Ln7ABOgOLQr5WXHFvW2y3Lj8CALJrRof
WIWlC9aPw5qEuzF9vc9cpoMirWheCR/eGcnid82MQgfUn6Hqk1bZs3N59cccgduh
JAWgaj9FNltPRvLlyBQnNCG9AsArjlmTixAFk8kYquMoWAABI1CejcxOQdsfQ7tV
0UUux+P5ezd9cCaKjQnoHYMNpzZ56Hy8J8ceVotqitrFnQ33aAO+rRBARtOW04RN
Hljs5Sb/JRWQt8Zxpyg8o9GqYI1vsMPX0mOz7Kk2UFxQa8ynohfWY8AgZl9nHRNQ
ez5wl6QjKIN0t8c9g755a05AdgSogKlcLLdWBkkESRycxhwppvor4ZPrUzeU7uae
OO66ggBOvboFiHJO7tXCJ/Kk1vu4m745Wy3ieAj5zGrAFY5LabGpbvMsrzdI7eZC
8qi2c8cIJJK+tQhdXQqSWeMbTqxkOXEkwqcYZHypO+vKbW/rvM3ZsmqA52UkeYXU
+GCFTscdz9nIFz/IYgE9Llsnr4pca+xj2I4xFomjBa2XoSwQEQVlK3afavzDjfXo
KBlBuxcrcS22uS7009VV0cuO+WigMl56xRoLrbnPvlYu4y1Nb0yPBhH98kW6xPvO
Ax2zqud05tOSPyTPPdjF1U63kmeZtnOUb+D1CWLRclRssArS+RtmrkCwLGj5DlXA
p1MrtoLVU1Sn1lFKzKduXCMUB6heC7W8su6N6662PSz/anK/jyp26hNebtH0dZP+
CGV/BStwluH0zWU78F1Udye6MALkMf/G4w95XAwKjHhc6G2AiKHhFGPo3DmddTRd
HV9pwRxvr+tZmvK9AyJzHy66zxcNtFefCOdkD1sq9hRt2fKJGeSxBj/Rd31G9qfD
Ifk6b4btuQQkI3iMpzGdJ6neFzx11iRo6a7byegeECecQDKfjDVlV36vzgTgUJHr
Y3dgFvUHFl0ynZIi77GZ02qIJJMS+HbXZPq0AkJKmcRgXomoSjjUOSF574CRnopO
CY2VsDRntneMBjrqVJaAJq+7YNzbGrgLdx35c6pH48ANWUM2xNj64m25PVLhnZz4
VTTge0ZcFSIH5skk7f2KFu4d1Fw29qbE0BXuTKDnOf9eZYUdDUQ6uUkv1c4FeP88
C7nV3e0XQDi4v5kKNBf9mVtGvpgEHfZTQPMVxom9r8tX5RTEnhZB48gU1enbdQVj
WVgjJ+HKBDThbq8a7TlDdPHInnEMdVw5OHzn/+LZQS6bWCu65lhYaR3OonV8xes0
uJZ3neT6qnHLbyyNVzu7fXqc8h240FT776LB9J8/2Qz3NPkLUjtYNCqY+KPsy/CA
qoVOSNdBBJ8RDsUu2VwQWFvM4tF4VvOMddk5eVKVXMkYjcZGYUDoRqZPf5Y6epVn
5qBOjHxbE6ZRiBncjN44lhcMyvpVPe57M6Csvei1pXWPFYOPiw3ov7i5aLCDMNFT
q0RvzLbB/gAFs1B6Ik7dgv3zJrFCJQ0kWimr41ihLY5PN/BQA7zNEoQ4MM3Na8OD
l9hZqQWrpLtYPmnzSMctXMKG8w4b5fvDCKAXvqq6aIG+SpLCEJbGh81HlszaRfGW
F3EtO8ExToQVKCLs9NY1iEjGhrniHMcT0aO8vGFGGzwpSBhGE42rDol1HWb5wQmk
a2qHqwp7VG/ElM399HJfqw9R9Ek7i3PysmL8YH1/husINnf8z9bpg6/QQAPQXcGX
9HlpSZeaXTTzC/2/Z+nEa984IWradNVZrF0CW56ra2IJWRgpv1hDzN7UaMSm5UO0
83vPocWQuxfw0JkbhfFfBbOi/dtjuty47GQsWfiL1aFZ1B5EM+1xddyXZ4AyJdzf
Zxyv6lCgogTBotP0sNdJalKDcikLvbB9RXU0K3xuTmSgpViC0dVO5cqtp0XRTAkb
a8CT/NquPIbEk9VMmhOtnoJBk22g6GEfyVZozzInMH/rCMjT9ML8DpVHednxnvN2
oMrpR/3AyVu3xeka6mNr+JRtAhEndum6cCn0PTqXOJNt6JCfxIywM1fawupPmIrc
XKgEY/GkVH2ArJgfk15m2OY6Zt6lwQgpueJZ92tWpvwN6ASzSQ1LBifT1SKE8z5d
b3UCROyKCwZg1WX7WKbVWxy7EX0U3SGYUNwwzNOkmztA2IaMP2imomGR+Co0ULSY
4NyuTX+avhJqIlPj3MGdKid/wLkqNIwFjyc5ENtwCj9vrhADg0fUO00IMvUEYFQ3
RGp0G2YV9vGZQhF54cZOh3nzZtvBQT+/gxOwSJKkHANQ1SnrQaYeTEG3Io1M0RVf
JKE8QPMzbxySYi2Me/oo3HGoXSLEV23p/RhoAC8fErwjmwydu4zgkpIwXx4oOyyQ
neagL0B2JYNQ8R+l+RsSDXGL1EDNse5PCyFx+UEf+C/UIMZPLDnFbJ1MBanr7Aae
I4slktrX0IzQWoa3FoTxIOXNWPclZ4qVQd5DkT/L2pV4scSk9EsfIRdzBfMlLR7k
bprZ2kCQxHZNi1yoY5ILtytvdkJb31CDqkWqI8rpkk5m50F6DcO8LOBo8/d1WU1P
arVCNVZJTUw275H/ag6NlLMRmpebDZ6Idtm8DafWemKUCzI4S8wISbhuv4qTWHex
EdEWj93HnJ5IpVlCCP6LMw/YeH6NoJIYT3nP7Xs5d/PhGuXuPs/rf5JMseD9Z2se
0HYCP/o6V0uLJ+8CL9GPv8YJsutK44Vnt5WLPjA6Z5w4LIe8iiGGyGR6Oyqyemmp
q2MKftil0QHaUkLt4QE2gK8YswnzhGUQwz6A771Xagqy95RyoO9G6KorTQtjpDJK
4MKjSijC3hI0/j7864H+Ovi/daL0tX3/yKjqGbAbBo02JySbDyKxmBHlEPn20oyX
ADcu30E7urftsyddoSN+iaHLaVMuoeSrbQAN976xrJy7Ih8Rr7SJDnxCDMzo9Guy
oicOoIVDraCn+B56hNd6sw/WTzuT6W6W8x2JCruYM3aez2inCqRs9lYWxvmefqTv
2skcbbDnni3u8W+N0wXsG6xisOYZs0sfuL+575ePKC+sF1gz8wM3ehmXtnD89CjH
l5eYuA2I0LNEld222nST+mTzGoxdzaIsPGVhHyivrjiYDz6zGipDAfwCdzgUTrXS
Mm2U+prVSYtyYC6l8UznsbTVGsJpebLFnV0Tk8ti2tX/mzqFBETGJGS/FfMPWhFB
ISFrsM4zKMl2iLV7ARNxF6qZhrcOC+EdrtRGt6QnxkpEGLsC/dnBl6EZnGr9QjCP
Gs3NTsuuW3jEPBaagXfLdT4XYtAZOz17cFK5qpRAGhMxG3Y+6KvJeziDJ1bIKyWj
7iXMzydU5D2sSeLul2LgOcspR6n6E7UZI0bWlWG/aQinA/N8fAP5sfFuZ9Y9z1AL
7FMH5/EWwk8IxSpsZXeXBQrZ3jaJhCsfEQG100nbZre8NyLk5n8gbOzUQclTDgiF
WP23ZuvKMn3cvCdX/Vsi1krmrX/QEH9r97pGjjfb5Jo1j8xLsOlv5qW3M2Kp26cH
vZLqrtC/ENKtYMSU1Lz4jDSOx9VOxfkVBe0kEYHudleAQeK3Y6VRjZpMoHtsgIvL
whp94h35E53tOAwhY9zuR/B77SbxZ9CBqwUZB0oMRLn1PjYzdnLTMz1bQ7SXWSYm
JNuLYfiNASHp3CRWlMdGeypNjyBKwL9lcR1kTkX8f9TCCH14NRzppgo6k7RqQwuG
NJmlg2lrawYj5L+cdu/vOOmb8QLySaAO914+ObTSfC/+y4eVLn3QT2dUhF+RsQGU
wXS42FgG1GEA9vDHDbz0lAO8kyPrKA7ld20pA/tLMIFfUXEzlqn8NxGQ+LM0ylRd
SpX7zTJLaPLCdKd1/6GivbvhY8+5Ci6XR2FNyS+cVT5cyQQg/s1wmYQ2Ds1S3TjP
q81a+kT771akvK8Ood1fNd65s6jg2bPP52rfXtSgKxsd+D0qKYzBI4i6HzJ2AwRR
v8f1dHgFwuLudPwe0cqsNxXPtSTxdGMqY3C+QZZxvSqDNBIl3t8GhEvEqtIodN9V
Zi9vd0BmY+49dX6oHfNJd2oZvsy3IFzqyq4X4aY5fQzoPdMYI9qCE1lTed8nTB3q
6x1/t0tmvILoRjz7u+YxGrVel+agPnCTo6wmfbA7/rIMkB4iFBNgqLDI0EOk994w
POhimu8O7YrG66Lc2A4nQFMiib46Y75Sy2OJbpgo4yoJuD+brEXEZimeeH9F04+2
juQCSYO/HjgGEvKVwQjxwXCeTm2gLefedlY9FWfE+IteXo0uyTdtCXsrm9yookIf
KmrLt5/u++4NI0qjNO4V0DKb0bKVuBQYY5COGxpoiCTnB6HAlad1FTyae01BMVds
sTOcGpQS66CAZPYMESBpnYEDVnbSSxpL4zYjVJUDrfUyLXYuvz0VYmQyrn9pzI6g
qnn/sejP6bt+1mHR5FZapgI+L0EbVwh6qcUlBS64Ho+itVgj1cr4v/w7zfwgoMD2
+6xZM3m2+MojiVmz5biuktjpFTJPYIqKRl91RFARUoQW+tgvmGjmn3Nr1/lmqhp1
+XkmdeKXziWzQuxqs+2Kn3/+nTm66uzlxT1LhDh4qtdILq9gNgbNt3UQmSp+IGOz
W3jlvdaBtAtHA+WZAS72+/kABQ2tmLOkavvxMbR0FcBDR9L6ZhfkGymRDgX/pz9u
trCbjYx73R6BbJ3QVjb9hs063pX7OxvQXYJiON1TZlPZBy2Ldt2bbcWFuQg9Fivf
4xN28bWKEaeTBN2YE+ogc5jsfYFguvBSrav+ewI3Mr2c6AuzaohhYLZ1L7byrluS
q2snDNxFwiqOCFj1VVLki/UH5IBOHplBFNM+SJlXTEBp1Pug4Ed5JlQS718pJY/U
TzfVuI/lOg6CtJ9CqgpT7xpEfzUlGGHjl64gXUFHC4sJcNpljZ56Ze8KIC4sLC8d
wYZtKB1hWKF3fNv4A6sXyU2oMfoFL3IXc+DpKxlqub8VHclLVHFiu1nFbsxFNH9K
K9P28apiFhlWx9J1RCBKw/bHnPMiUoTgF6P/FyO9/8Zuv8a7Yj6BVrmfQqxzzK6n
1BY3n0vktQv/efx6a0zeeJC8SWTk4toxEwvO2UzxQrJV5ioJpSfcTLHZZp+0PLdP
o8JEca3VCjyuBb8j6zIMH8H5Rz0T5A2DTd9+NIJCJMcNTZoknf0wvgIgAlrgD86W
+ctiREzDmUMHxxqNL+MU+orczNLiBzJIp3L16N3Ik0f998giGh3KtWoagdt3ND0+
ZqcwXeEID2bWtHo3p5GeNnaFYsO+FRqKTcb9NwfNVHa6pfIp384X8vLGFki/AP6g
50PBDScxmPPGSXfKNOFkrApmKpqJ/2SukKbDWFaajJiEG+IgE+zSs8j0W7hyLmoL
TiKU5LP/wgptYTezZlEOflq+xGgvDdhCTkPTq1ihTbWuPa/AiOUlMBSs7/pkfabk
985JtbInYiQ0QLFDiyVmdm3ESxl1RovTWE3WYVbg8qIoRVxm8htat5UBCEELWM6w
cVAx2uCRCqghvbYCGnb6vBvbNzRH5FPVVRuhrDsKbXRRfbyLX5uKI/rPFKqRDYQc
kfOu1rTjaNbu5u1VNBvHBvvwpI8zgkNUwGsN60HGjCnCn8NhsOKNJWe3mfAowYjh
vB950EGMMTe7KQnsb1XovCDVRo7XgKT/jfYWvnZfiv7U06O6cFlztzYgBCzxdjKK
27Smp3BM1FYDjQ4JXs3w9QDWASDUvMnA3ixjOZnBJ1A3a9x2QDz3bx2tCeJWElUR
1nIvYEq1HrvO7EuN47dlmL9WdsRmHiadiChuPLf79DeUuOI5g7+rJsJ2jWFOYx4G
y1+Skn7fcBa2YCdACMcq6SJEZOeHblCkszrtePrIoMNwFEzZ0sTRtR6IlY+6+W9d
Vts6/ch8acMC8b0n+nDFTyqJh7Sd1x37QMVPDxEk4sSup2SFir7wa4h8hZA7ADHD
RIIB/YSHsIJvxSkZwGsFfR/pelXkHOHyTpWqG+VhdKBDznHP41wNwQ9uXS12098w
mA0/DLj9keOc2J6as7nWxSJjzK3Cnaf6ho7sDF9WvVMWpiNwZK+h9EPtBTiNhVEj
2IRunzi1IHRtQAvNb5MnFaHEA0j+aD0bQQCkhJA5tG3BgpcAlbSksZ7jGz5ZY+oP
szrdES/XQyT7vViv/D8dsFpTA9zICEEyQS5ATdEimo9D8EsUnLIVwMZnu5sfq6PN
uwkKaJeqgw7V4aqyUsxOfjxtCdNsqOw4AUvB2zCzK77r9A6KF7gNkMXVsoT2wM0G
81Ut8y94w71rzJKUVEKiYUlWruHdPr6OR2zhMDQpe2ZSqWLf3rgdfn73QrUyGRzl
rYwfGKnDvCJtEgolns8/w/8A18X+PZQPELwnl0DwM+TrJDkGkSPglYdKhr/k60Hy
3I/Rpr4esUHDBM5aUyQZi4HVeuIq8dq4mUDpQP2DgUfUPKltWxjb6c4RohBHDusr
5NkJ6IDRAlYhX6ut4WmNC4r5rfdrRdBwZuMPmYrvwYpRb/lDu2AXgTAeDGiZdaSd
EMBC8mEKmJqqkOCxAj0kL82SNEbrbntnMMgamKZ7MyvyTcxnFr+LBp4Sl1hyIuJd
hEwpOPOFLWdU8nD8buu/dRghWYhDhizfqnYrJEVda89mnoYHa9gtw5SF56OButGZ
RPkhY6H6UMW9j+A2UpRoF2MWnUw6DER5MqSn+z8kTdoXnaikJsuJ4qORmTtt7VZN
kdgZiAlogseZ1FChlbxaoBY3GnnquC+UhE+qgd/VqJv/grJSFEsrIDodo3K3zUin
TbneewMxUDOWr45dC9x6AmF11peuh4grMh2Z4aCXmtwJuhtCRz+5KgGQ2fuJMdJ1
F0cd08M3HCHDy9V5FTW51R6rhLxSG5lf6OIrPBu4y41hmD47RJLlLKSzxmZSose/
TCDlMig0qNGZvuPJG3aeXhcLQf85gOd0znt/gNyGF7Jv76DxKhnTv10n5PRp5ftt
YC0NFXLDUwKUQ1okm/b7iOVfD8AMCtqBytD+ZvrTZoGY/t0/T2/uptmrkCdpbyyl
79VHkE6QwVH3Fsef/jMAIOCjHd/hkspCv8lZrLN3HYf9FX8G/aW9EL20pm6V1utX
FK9ZAyG5szfK+OjKt1oGrr7YXXlB4sFI6sSofXxmUYMlDuJDeTFWnFByxzz5Tqsr
RGVbGz6cjkEP42jInINDBT9gBcwIRLfI9/ipvzWWPP4ol6MUOeS0y/8YWCFcStFd
fciIaSoNL5OafWvuY2HbFDc1Bno66W9QnTx/73w7OzNakBwsfF7w8BiBENjk8zcR
FpEmpd/1AclnfzYDaSNq691pkhoIcml2AbZTpSUXqfwX3zpDG7LXoiW8QfEmqx8E
YRiGqc5aD2mCm9III3a4GFCBHME7LD6xBFnrHUp9qkO2ZBMY3Y+EER2CBv4Hlmli
ujkA0LrmslCrCibVhqUKWfjC9F3rCMO5QsI7RDT2ATyBvLbCDvWfkVxhYKUEpsA9
t/vIkdglWhsf+3ODsrimkf+vs57VHzrah1YQGM28ijkaseNTWb6uy90ujVO/uOTi
SmvD+F4XbI4IHvQpPegUNoyY0QskD7N6Y3DiGo1/IDs+Wr73qWWa/+6IGnkI0Eyt
R8aKC7C6vocSGkpIjyaUFQ/WnsOdZzEbmcubKFjVz/WpLfj50zY7TA8E9GruyO64
BEUchAqiVkfELy3nsvtKOQoW+hs9Ih+/1Cwlf3Ysr3OXyaA6ZzNKSIyktFl80B3L
JvhRQmJbkVMmlPT5xIsmC7zFpETmVDvbca4UQc+5LQczDFkTOf7aKi0jY3l+Wzhu
dD1k4qJCV8aUfvesUeZtEqiuhznvSP6h4tIGN8OcQotaIXELHCYqv+lVDo4/3pGR
Nx2sI3DBJiZ+gvUugKs4QFWKdQAbwmj0PkLax06GNw5jbzUjHsl0SsOVXrR+jMyo
zyaeTyc80N5eqebRh0T57+ogVFfUPyDIek7o0zkTL4yByClSxxuZ38GLtpniGmtD
JVKQNy3HLTCvQzWWBk5dLXHnLM4iLOeFFU3x3cPLEPEcQ7u6ZXRwt9yTkUo9fvIM
6T2YwVUImf0fX0mv6P4o1fDWyLYw+4Zpp9fP8mOM29SlB9MN1+5+ixmXwBh4bmwe
Zr1kLST4Thy66aubwq0ykTyZCu55iTln4o4EZKPzt8smq77CMixJYwI8/BvwRxmE
C/y2WsnUv5Y4TFbVNlCD5pQIxKEzY5Qqr7oURsBuJbFTdATOdGbqUwLAmVvwS21k
lGwOw0MS3zZDl0rJ65vi/gi6/Uq3YW9jaRQC0zhtGYpVeNq1aWMsOlzneYpB0nM3
KnPNNec+yBpKJw7hqbtahi/6DI9Y6Q1ZN9tvKbx2k6+trCr8uQMnBI6aSMukwYXb
pT6X6fdqI8xyE7Ao8ErXlmIWI15KKZYQC58Jv2C99A2rOkkksMVTOH1ef8I99AdE
RePbeoA1c2l0y7jglFrFkJkLSNKRxWXRVeLdNZ4ydSmXLNaJ9Yb76H77SuBYiH3J
FtP5CkzFwS9GS2wiBbtYV6W8mkoSZ378MyM+45U1AMqFoWuQzZC1CbgReKqS86bL
NQs/swss2Kei7y6kgF/95Djhpf+szEI3GfJrtgIf9JD0bDX1UBLsZjq7uJ07hbrz
5F5sd2XM5OUwmClq4bAV9Z/yBywApUUWNMJZP+GH8HkKDa6nEVAaJX/VxM8m5mPS
mRD+1FYHQ/V1SojSOd3hCO7VbaWEAKy3CO826Z41NE57Y8/oYCbezfTtuMWMON7Y
M/aPdtD7vGORaiFbWnQ2dXNN5dMx4LaZJlZTkC3ude4FNZtKEAV0VCdB/Cif3u4d
Nr7KkOWdE0R0W+I2AyxZudeWD0ZpmHZEIEyVeaI44CljwJ6Rzru7Amn89LVMlB1h
xpfJ0vflzmFbeHykFSlq0fUePAuAmSGVtE1Q6clysTha/cv2t+t2zfV2EBX8ksVY
OhEpGos05e5SkCLTF1Ab1WIKLZnMklFuOlecblGeeGI1akOUDj8q7tmoq1DjFKjC
wI3K6rAHTc/m13YHIhDjsjy7mhwtlj4yluWZRTqykAcPVAxtN1ya9YJ2k+W5G7IT
HYZfC/xHLbRPitL5JLWWMR+IFO8E+kmf8T6sphMG7dyxWc7JVGq2m5/kLYaSEFQW
nr3UuIQju65zbYeu0sodLDB1yPet7Ui30xCKlQCdcCO6nlFU9Mlqp6Yx+NPsIEVW
omMVRl1pXI4SVDkfwmbd1UgFF0wzdDRzBPLB+rdo75LQ86BdNAROVFaxOVsjvJA/
W/F4cZaixMwvF1oHVeBbCSoP0B+8FO7WsYlK1LrVcpnCRBqKc209Q0Cekg2fl5hJ
MTFbGwEYTvdruMhxWXHEEVdXx8BisgAT021V2Zz09NMcNdmskf2Np28MJL3rSNn9
+LgSV2ss7p5cKj4el3JrR90rWOJByYutPUXKfDLpK0XK0J2w8lcvoc3KNsv6j4RE
02HRTqV4ioYV7fNH5KAt2ubjYEryELe/pqLnMGr+rsjR/C6Md9vivb0kFumftfsE
zmJWjKcZpA60PK4X1V9SENpK165KqI1dpflceTZtMwdQjMm6gkXSk0npmc3q9C8L
8gpAY3GbrANoxugnpjke3DNCSdbAvfCuETc15KUdH6hstNgyi1CUENdlNXoMIpeN
pe5JWCkhLTpgYeOzEkY6w8iY/RJEIYHg7/ec2LTSlRXKqbuTxfaYjY2wFmZSvvf9
AosVbWoABozlTvDt6SbTK4fbNZ0pJbgSkwJOOP3wQcSJFTEywuGl60UPXJSSbyXs
2PRm/N8ITaRO8a7G9NCEit37oJlCumj0te1FfpeCkcsPl2quUViPKntXZci3EDch
9U5yf+aGh1OeRybvCLgPCBhRJrVlBcZiB8EeBDjMABDzxbRQz7hpnCFZO1HHhJ2/
8NNJz9J7N4v8qjLlQ/ZUvk/ve5MmOd/8SK1rIHzHI4nX/1KGsOLkuOPwxl9QRtyc
PWYb2GJ8dhy2e7HPvyP0KpE7cQ+Qs0uz+0KkKN73M4Ovt8D+t4SKZffLWm/E1SWa
0YJEgv6Dox8ScD5KFPPhDbeydAGAdTAJ2h1tLgnWI69uj6Dx7TaMopa0e+KUQVuB
xNScIrToVAavhH5LgUbh/28/t6l9oEGRmX1KJfyjZjv2H0xFuQN+68bD/CslUMWh
EHmtjmbkkUoEkC9VmVNvJH8BKU2gFhenN2/oaWRSAXLcx9WeHCgaBpm4QsGMk2pG
mEz6sp8J38uMQOa891mV4+fYxDDmIGQ2yK3d2BHwxYp8usu65seGxbco+zgMhYpn
S8lM4EneUxQ89CpQtXjQjloz8h7b8kxk3D70sXqczEi5b2SCV8hwA3UNhRj25GaL
pzr4Pxf1U0NLRInGDoVXrYtVJOzI+fWJzS7MW9R1Gi1jfCQAa51TsNIofuHOOg/S
7L50y/BGZqWNc8UMp+1giCY47+qf7YsSClb2TMqnRXKQTS4iOdvxDBkNvneTK4M+
6taUHXxgxpYb9X2lk85eAJ+mjG1IZqcfVjjWU35bVQzzzbTNYIfrz/Zdmfllx1U3
ySFs/QMYqT0XXbm5xFPRnpX522x0nSAZ/nrBbAlI/S0x4Ih0YZQgLcGOC+fRvdzH
Y3Xmx7LvCS/ix99MuDTwIWCGdkA69UmyJg4fNZef1lVnmXC0aXFR8CbEIWSZ/+2G
dJ/m1DL1XW6A+Rg0E7nehrtVyC825cnKA1+YoBN0gvNycbJuM55FQiCD4kUXz3sz
fS/XaU6TUUd10istF6cNZxU6dMK6jVWt9V0FzsEXvxUBC3FpPQRmQgF+YCm3uUyi
DZVbZMFxn/iGqlvfvtM48VfsuiqxVfCpiZ62C2YDa9xLb0lT6djoGxgUulY7kyaK
yYRGxFc25NgS/tKYrKg0MkHSCZJg2wzDgJng2IoKOagJWS2fwF7nI0gd7MRK9vH9
2YU9syT1B7uYnTTXbELav4kz/7MhrOHIjicclY4NL8PqiQQUl1S3hNCF5ZNXZDBx
QC7jJkst15QXWZ7d76AHlSCB75fJIMQ3kLHZypzdGb5fBm/NARrEGRB9ppA0CBii
hJi/TOHnbCrUP6n5m9qmOCs/0YFubQkljDruo2HonmgD9akPHxvQXxiOgzITZqVE
pCEg6M+h932Oo6b0KfhzJ28RhTqaHvywfcxQMV6J3V3ormFM4dd5Z1P0SOUUGawc
BgwQ3ziYyTZ0KcehNFTjyuFfm4SqnU3JkGCGo1MYrQg5eVRZ+M985CwKYx5XtEmq
FGax+NoWKuQcEkfitX5+0ALz95xAsIMuV3wO78yNdnHm3xNqidqVeVoGLibR5gtC
WkpT0tZJqdmbkt16jcTM1z7xB0eTkD/fo4yCqTzgicnhFHuDAx/DnaYjSB0JRD94
+y9BctkKMlNFxokKOr5IxG9xJ0NzmmZgz4Rge3LxTOxG8PPfqy8JTV6mNsaTxygF
A4p0EmhwvZ7ZQWPnoCuCj8QI8K4sOBkJm5BtF7arpRIkg63bnpT2IzXQ6Es1QUon
hRzQPsT3keAXWxmKMcDIC1HncKTC2zbpYYiT4Vfiv8/UM2fmeNJvjh0NID+Zy/oG
424Y3sjUhwIamWou3m63AwY1Uolwyq4tkK8v20XmiJsB7x54uujGOSzEyHEKPq2x
ky4Ccuc4X2ChjsgF4VlH4LE4LynUNL8vpDIsuBO9L5dPy4kw+YCG3F7v1knr3+Lc
BwubWGTNpi6L06EbzxiIMUHEFcvHw2JHWEVydNjABgzqYwh/osmY+3KF5HGxnbJy
s2IpGqrKudVIwaYTWJTRyKbqz8a3s/vxqQijfK6dlcpm41qUg2CAfSTo+auGworX
mUKWXzlULnVjdPt38j5AmBp8ERxHurul04RIPSGgnW2++/RN0xuyHIjHQIGFSmNN
vCDOD9WgE7aD9PlYNwjhXAtmA+Zu5Bkqz19vBAl9zOupmY2dXFlQSt4cRwdO0Lsb
4N/QnhsDMKCllqIkMtdqgqKAfhCVmMPPfKzdZ0co1C2ndy/bw7zDfxfhWovI2We9
9l301kKUnJTF2jQ4yxSnMn461NS3euOaMzJJOtEFyCbScLtDlULTqcZVZ9twFhmK
3s4D01gVQ4sACxdJdTwvJCgWoCtvqd/XX4rXhIRYI1DD4EBwYueLBgc0TifwmvQd
0xFoKT2rybKDbm8TNeEe5mzYw/DmSB7gqtwYst5ogdX+fgkVF7VQKaQTzdq3h7uu
PfTRWhwfBktT4CPFSJLie305kFw6yvZ0VGAPHSeiSH66Fn3CxBXhy5U++9oJCALe
fEeCCcLgNiApi5IrOw+ILCQaKpcEBi4WgF5RtC7fVqiKiklL4kUj5oqF1xkq9cyw
AMYkkLLuEDBCReH6Wg4RmDmo9SA4k2DzrFieJW8SpNhQeb8XwPsYcKhSAtSnz74U
L4/Vdwvp+XKGA5INjBcyW/YHvkvh8F1fkiswkZ3rC9ds6ny14FHm5o+DOgNmo5HR
xzUm5xERoedmByXx1EFtvMgdN2t4ypZ2wocsjR8viOdDoGy0JgUvN2fypLQAv74h
kQRiJGUgVUXzZjvzsP7PGrFWj667s4T48hvjd677t8ZuciVPKjRIlId3SL9rX15x
l3zZpg66/oVrGwH33owi/Wd5GqrGI0rW1RtQWQ/Lj+KNQdxhZxuca35j4u/BwVqF
VDyLhgituKVwjH5ZZjW11yVUZhMjFEA7WnCAz/3fdTP3UazKupU/ppyDT86mhz4V
3oYf5OuE1YUF2TJ0vRQy/TYCCcP3+N1FNkW1OMp9u2sj7i3eGc8NMuZuezl6E5OR
RBuktDiZm/atdsjKLxPdZdBQOv0gWfQ9l7yWk8KxxEVDHEMpVmCp2MvcEcP0dXt9
VvNNZIQ5y1QFfn0sT9D6sFjVyd20Y5sJHUOenwc04Hu3AnCjo+tqkToIrMh+peL8
vaGrXOqgdxqZD9om+BlZ7wHi4SvgzuZ9cA461fuX4usc/cqUDooHShmIfBGBzhRb
osqD54gqonx7kxl3lZIUj8GlscKx4k1NEf3i/0C8vJsOCPeHto1wmZg0vi1KLkOM
DcGOeQRzNm8jJv61imJk8DGUy9wzQj8bDWD8W7K2yAez/X9M/DsAXqolK9mmc9Af
OxXaR8EPfm8SAvRxiKYGFn3zSP7v67BrJ0bF4RlTuUVWk2rXRpZ3UgCP/RbKhZzJ
DwhD+iFwHgQYGTPoxr6LBARL25s5w/WnwWEtPyJloT8nWgZWNhZR6L2up7gV4+Bs
sB5dGNypy0r8t4r5sbqeaFIPW+9rLqkXRpleI3QoW+ZfkzjXLNdzTp9fzVjsigb+
pQVaLSH3RbIMqVs8IJxajMPd9jGI5pDcGEnFSZepZU2VWhCYjVRKHofNLF7nHiGp
HUjNS5pVKzT5h9+/zXKAYuPF4B0aMyxRsM7FR0Q0cIdY+rm3fOPqd6aUeYAeZXZr
3ZSqg/Zcncw6ON0zU9wecK2YgWj0MeuVgdReSj1swg/mSEZnmemM01j+QCQCz4yY
cHhUZwTruRnjKEiJZs/CenU1riPxInuq9sDOsxzYBXqvoBYvZViX6r+sdP/OeqWr
jY386BcRMNkzqGHoq5K8m5l4b8RgxOXQqZ0lSlQTR7L0uSv6gDD2VAaTn5Hy0ocK
PQgnIUzUiA3luPihuMAfUs/wMqIUHuqcKNcHuOQVTz76yf3nAUPepu4mJrx5PHGB
ZjPdOO1lK8xbtpC2KBI9PHbuFZlMFSLsMm7vZB92MVeJ6/9d3CnDApU77AKzcPRs
avBua/+xoJvWv4NHIK0dZ+EAO1Ymnq3EWLGEnwbg7yrIFYVE4wBo5YdIqwlwO3zA
eibB/yLzcI5pBenPfm7HfIJYynKGTuVcFct0Xakm6WDq3wJhgqJMoyrCT27i1/tw
zpxJz+4qSPjK2T02ObEJN6OteZyBcuCRlIJ7pf6NKIu6rV2sTJyVei/G6HHV70RN
Ia+N20uLMCadPxJ+dvlOeEB+DPs3YiVUtMHMISkEwV1YpcCPLY1eUlQRoSHMVVM5
4jmXz1cDWee6ngZtDpxHm4V0q11qggOsowCkFQ+4x6MtBw79exnnP7mr4mLB81cl
OQCSUUoemj0cXgU+i/FFe+LV6SWlfdwmKQFz1U6+aJ6w5M5pNofMqLMCYKEYApT/
1uWZpH1VxxxOOpfeU3WGHxqNsss3VW1PNdGCuDHWci33wkD0Aj82lynRb/75j+ZT
sUvfOkq/M46SGiGO80QSYRakQ1sSmdjl9RHGODmYJUiAgWjuPXHVgWuFszL0nKg/
aqiN+4rEhCfmhGI9W2AifVTw4xMWbaXbcE14lHVhaQ2uYX5OrTYf8Tqbc9lb8m7Q
34xfOEtq5q5IyvOnKtZY0iHQW6kYFV17WmlrEyAfufLDky3UelGNzOs+SwF64Fr9
Bp7sDy1sQK1xU3dKZWzdOCFlrqXJNXPpfUAG/jPjjmOfp/uyh2q24FSRNe6ZqwvS
wNpSW0xKs1X9dbkCvU79aEKce9Nzqvrc71+O1sQs9j0FuUzsBpcyTvokD5BgGG1O
000QYsv8hNwpLoXWon4SQmHdPhtBENdT4FemZQa5cwbcCyl4jOvf+D1zVH94vmle
IpT4uf1Sk4h1XsI/gdWeQHzAJQOTdeGjB/G9VJuTuCcG9yg/8a+6EN9CwZ7um+FT
6qkP2Cgg2uIFQvGNL3l2tRSfI+c/iXYITZgr5TreZbXfoAVKnUl6iKrkqyeZRQJB
B6BIDsujOmRZq1KDQrA27EsKHSGi8u7CAzgoW3VcnT3QyiA9X4XezdPPqrF27CMm
S6KL98fft4RkJzQwOSfLj7V9RtPLNJ9wQCF1rPopMK6WiJiGVfpESe/0bTW8wo8W
6SJC1lmKlgcXgI0HPG0h+tEKYm/7I/RmYAYsZ5sj/xgwPG8zayrhsYEXfC/+HI6g
D8amfs4p61FyAFCCHvWBKuEvxJH44D0WladLBla1cOOMSJI9bKDtMCH8cyiSBjRE
2Xn52MG+pI7Tr6vj9DjBvatoGyC45ijEqUWBWHAEKpcRPC9Q4rurvbZcjqMZAfZm
GjgVK9j/qMfvLE7RYkC6KdSi6Av42PtnUVDSwPHO1iBljjQHHzdfToUfFUFlTHYj
AGcnwby1z1c6zzlWTzYv1ZtzMDfCLa43sY8TD/ueuadKgJsY2szi8qsRVjoXq2Qm
GYEJMCNWwAq4zWKREjuWTKMFvO/AnMjBDxNB1pcDkSaoLbQq5EckVUSzy4tPft+8
0Jp4GfupvaiAYxVNyZWFuG6+M/V7iOnXtPSomHaiC+QFkTfxebotZCUnd497etHL
U9bsAdAcnkynrFSQWzpP/2tEf6T/qTk7E/YzVhNAp9VgPAcs3J/vX9V0XKlu1gtW
NEcq+qdpm/0iAZmwuhhGhhpBRlMcjuwvb5rdNbFTwhd0S1hNxfN5Y5Dz2wEXe/Hv
2Iws7CgZzRRVUt+ks8u23ZIKHOEdi6v8RLII8/l3WfINPaq+TtnVyuhiCxb+Hmz3
3Ed2mnZgfkR4OtM/wtQxwxIInfxDgXpZ2+4EDcprzVKpLIgZuF9E92Vj64mWeUit
0OB4N9PKGiJ+ZttXbDbhfEeR+HyeFRYBGLjDQlh4psRlf4ZcfLJ1Z9PQdWbocg3t
cfimIbWHl9Baddh9DAyURZ8e3cApY5yvMHMCTkzIkxjC+xJW1Wd93Nd0XNXjY1wo
VfijPo/fRYgAy8Iv1OiJOuxBIm4mVVG/kakNPF7nkM7WwFqNF8S9yTZeFxUVFjr9
PwWzUzvNAz74GnclfyBRsz/76dhPZ6hWsumAvmG1np8IbGU/DWeJj+y31r9LZSsn
4QE26wVOUrCIWJf2JN1TF5R/0ZBRhG79AlFW87DELRxp5uwNxjYe5OFPF2xK0bfC
siO1r1Ezv6JTFCBHXy4Wu90BNe/pwCx78uht5RjCbmJNCex7bJBKigwx0lGkaIb5
lou2t+gIizN98v3hjeCB/imbzfrVGC7BdQidvRGLAuFUvJBsnhuGoZzCa10n30ku
8knZiyBLf7VhJY5wj0lbu2OMWr1A9+uG1waatPNMNKWoY5rX/oI1fCtWQdrdLHul
o7QfisAd6rzZ4iPAtwsCw9pvJg4SmyHZ7dtouTrlSu4IKhmsvjhCvZ9WFRnai09n
PK3TulC0t4HL/0WR76bljJl5lCnRliYBcllsLbvOX/Z3fqgmT9pdqvZ5Jzk90sXE
FzT+lPLiGxL4JPvDdpEOiadJecmLdOOS189Lqyn45yOTWZQm60BuLwXt614duiCH
elhWqX6i39WikdKmmsAwO8LUSerznms0vafqTfZTD8QECBS7FXoXU1t1qWndZ5Vj
SUiJCaKWAe5oAUpYJU4CU/BhL+NVvgDBzOw2F5NXpuRjIhoNjHHFzpoLzKAMa9Zj
BGyDqDJvl0b++fCt97ThdG2WVN/eiYb51dPhG0Bnu0dj+iV489yJ/BiNwzHXw7Fa
M7xG9XuqEqdD7AZUpIEjIaDjZTgdBlTvu2xz65GyCtSOhC8z2+mzncUfr1jnnlKV
r1/Tn994+WHib9kUp6N+EFkFVfVZgImu+LUzSEEES4HGHqX2LDRN+LDHzPcSKoSg
/sXZVFt18E4VDcXDe6j1XXIXs7zvw5m80P6/h573Fl/gbVTk92F8IwQH96IJ5ym5
5BSJt6Va1c4NovtUEY7ysg2JxeP78fpOYqG4fyhzAkXMRKkKadsKwcqdiLwGpi03
ZuNY0LZ2ZRhYMoEx95P8KjxZL9BYkDCHiE7uyR0weQNJLEaO4u6CCWRBz+ikLnQq
PmB7qmTegQTWMk3RAT18GE2K4v3kjxATlqc/oGteMJ/sEjIeQJ1vuanAUjsg/9my
6b1PyjuI9zgs1uU5Xqbh88tqwBFPcQpcroB5zz/OZzG+TJfAzlCwMjkegjGB+xyY
QCQ/V3VJqUbgU4ZMAG5M7sXEgQQayvJcWrx1jDTqtV3Mh4neHlnmUpaEPemaKhCc
+Rx+OS4Ma3rZbfwFE0s6k9mSWHtlns7/BR/337N3PvazsmtPX+JTHBEXrqsrMR36
AlgpVBhKVWb2o8nH2i5kNyVCMOU1wiP6qinpiLYdbC+cDJPK1bZfcOUFiqO0v+Bv
gtrERH3PbvKOm1EcbFb7DRoi1SHPuCY10GNGpRGOka1dlCANIS2Qa9Rr7WPOpcIv
WZgy7I3aDhpDMwVoAmI2LPSmhX2eCNuV2+vRnz/IisI1hC4Sy0E9kPqPsrsM6G6f
6ICTogyhcd3zvGevoAHNoue1gG2nGJ23AKO1Q/ldGspWZrs+w5Sl1jZGkrCSJf/t
tLrbjijD4Tfhxqt6xghP47/yK3BLrPeOzpWqss1uRwFxjrjUdA9q80rLJ1uVSXmQ
SQiUeVujZ6ExqS5J8PVHNXyWYMZ7ItUvDxy197UKQmGOU0pM4udwr5KHDZS9+M4P
5lOeDErmU5RAdqX6Ec/01RXeJzBE88FXPKPEt5UDhdU7RLwWWrkqHv3QSPxn+MbL
qhwTTKhCLQ5nfqvrE2Fk5KOCkDoPOLRJ4dtyhN15c4wbWW7md0RyHVfAvabA73aW
wynpKnBFSQvicv/rUZ3jdaW0ZNgwBHvJI0UhB7T7+LN42dY0geWP5YppmC3YZCgu
JfnJ98RQIsWTElZkicHiyAgTzzdMw+nPCbdYynHRoEz1f8mESTSvfq/BTFleJpOr
C9+bQVXHHSWHY5qhbu4aK5cDxesmxIR4Cz1pS7ozez7tqVMsRa9B3TbeYFj/79GV
cX6YL/YSoxZoi9ydpxkBnPcS1Se1fm+NGYgE18/yLQTa+DRtmEVM67e9up9fP+nK
1AhosVI9uUlAVLZaiE3lx8IaxpYV1hNm5uQ1ZEMfF0US0friUj2G4PNHAr+Wd5cA
GmaEceeqk10D3iK61GHJazDkYVqJng52ptJ35Fp4Fk/lhaQkFcA2yun881IoRd65
cbJeJ3FGkk3cCry13Uzp/y04XTxwS/0HZXvWo7dslrRRivlvziTmz8yX8J0RO+Ss
gfgEdAQ+w6bjlzMnh6sTDnOVppejHoDIYgwSzeC7UTbk1EDDhu8RM9lHbozeJkKI
gml4Lm3Eolw8qDPAuvBfrCxhlphGfEl55XRXTUH8Fn8oD7ngGuuedFlCDBlj4LSR
v3GJfTQd1ziccuyTZLRULNIwTAuA9cEUPM0X9H6LC4ibfYTl2+QBchgZriVZoEOh
os96QmEe8yWSLJHk2ftkO8C6317fwby2gtOD04Mtgsm7AJggWxbvR/5WbDOk4OBC
q9pX1TCUt+kbCjxVfsxCXlXmEaEmK57EFlYsauyqqe6iWXWy+LfLRFkkcAxM6Fwd
z37zeu2hgN1jhhadYMYNhBrl3o5PJZkhHjdMRlCQpgFF/mm5gb1puRZq5rhALUh2
aBMoDGmfGtDuSym/+gZd22q6jwTRi1ojwZps5nYekXM4DsmhhpOJbGe9Y3rhM4tj
fBTYoX1v8Cyx970pGf5ERyF46oRfbZEdbjrE4EPMElQGjXSMV43CU7kGQV5zWY5M
5OsYPtwaXVoO7uK+Js48o37MD1zgQjZuyWwbSmguhRlkFj3i8fmCbPBsTVfWo4Dv
X07/cB8Om7d/RxHFYpd662xc3G3YSFUo7PlTOCGSHcDUBMVVHhA56/LJOxbkCtDN
b/Qidnfz9vuUJkk4ErUHuPlOlYnjYGAO1/osayjZDZokVCGtNFJjTtaon/rI343h
G/ixAWrt7XLnl1agjg/+Qo5dl69os2VAMmoPXQG3Koj+MzgcA5geXkOKSWvOQCZp
ZtUq43sSAGNTjed7M0hOa70KsqOKuBasMYdiMY58o8gbHFcWI2ht4lZiNbmK9mNj
4/jaBaxummTdO8Sw7lmL+dDxv+Y04Z9gmpE/VxeLChnNMvYuTkrPm6zKXlLJhZjw
23XY5DywcrvU9F6KbnUcpc6e+MAzct623G3a3d6/eBNzr+CN3EbwWlxsDEdaJ6AR
cIfbnwyoHIV6aIfZdYtntKnG2wsDWo4ZqOuxXzMZDoUmhoMH9uIhN+0UTC00P7WA
8COV8U7FzTvIJ6R1HFqh8rx4+TWsOcB3bJpBbE6r1b5neAuhAJnnhRFEQPwlMWMf
+35hPGqhcwa0qU24jBvN8qCk+RUXSgQvqKdeaId9UGvb7anAweUTSMzcuZYD3sos
0TY0mYj+ekxoOvXS9ASzHPZ13SE/nfkyvdHKqoLkusr+l/FK0ksijpMA6gCyi4iN
DwFwosH1uQ0jC17gM2yNZlOSHo1ljUkP4BZvW8GKDeNWIeInV7FCcDqPhits4OXZ
ULqfINTtwzbMG5K/7aKO5Y1W8Y52cXvekQeg4plUkZY99W8zx8kI2qGsuqGck8CS
f58m4VbNsm4OwpxkTNTgXQjWnmqNV8+ky8ul1HWqUaTUK+zSrNSfpLfHok0p6sye
JJSkZ34TLipb8swmonULKpJcULSjud9jaL/DF8UtDvfxyicBR5zbwu/P64f1fMzk
p6eA7A63TzzWvsW0p5TP+KcIUNxDYBUkfxfzxiMxR2xqo4RWJOmjDIAGc2qcoE+g
+hrAUuuDfifpieVyp7VfH+JIBFj4/hOfWPNRAhThAI3YunvcufT2+t9Ea9sdnmjb
JvzmGO8VW0r54Os7VqRoAdW9rkaqV9J+nul5kXdyl1cvNvzcUtV6msP7+xfmLcrQ
GL1wbodBLiQdlrzQhcyoBLiBha5xTT6PYOps6ZiObM257qKMN+3ZN+DSfTpz5Wnz
53LT4RapgEft+Vf3G8SJSC4riar94LFoIVxr3eUsTx0om20bRmIi5KYsaX7hWoOn
EhBIy+OFCwWtZLVlSGN60hMW8xgYk8xDCn18wj6DeNXIlB71asJ8bP7gJG8UuEdF
+gfrhNLPk+zhRHLfgPUrPVOtD2ug5VUryZDHg4CA/eCSlVwsEKfisYrbCl1GcbNG
Nf09bVBL8KyZw63eTi64tElHIm2CbeJTuqjWw8YpnQczzxmnEfTTR223Zyn5nsRS
uoWi/WgfLb+qmSwrR53N6pEUgFSTCjUTHHFARzWa+9Sdl0oA3OvN+sJi/2VvYgbD
h1TgqLm5oacoH/w40laMNw4Emunpek5PgnLdkx5f5oRbBQe55+09mnH1NU5gNiF/
3FOmIPq16LJ9rzqTj9luUY6Y5p2yUSVbbIRldz2HOiuNUwSv0FpVXoUwEIctl+RF
FUHGaxsH5pmdSkNkamVOpSipkfHJh0pbZ0ChDE5fZ3+dzclcYxaegprSShe6NQ9s
BOBVTCgpfoYXZpzPLz8ZaRP9CzAR6DF6S0zPy3rMeMQ5iiT7eLd3vcEdJ4p6TtNy
xl39myaHtc3oyl0huE8iQy1o5JR2Rg1kGqQu/5M6yWM8GmVxT1HrqVTcf72zHlxc
r5wjzGS/sNhVS/P8RNTsyeG+Lnjv5AYW+xTynjdGvM9KgqkhRreq/XCx3DrhDm/K
IXGomPwrDUAKm9f5JpVBUU14Pajn9VdhBsn+5SmloXYbXRwQfFc/0kfpq9BUJF4j
FHTM1awJD01XeAGCGf9DMimKesvSi/fP+bZOSBKcZ/pL30H2oW/BsE5W0plDUCxK
MDvE4C099dc3BoxaEJXPioUM0aG7sVQKT5Bo8vOKgvZkN91UEimE9vvHv5jBX96A
gULflV6qktX8MfCRYzfxZOspVt8Fo0wmObQ64hDnAa/UlWFG72EfjXNSF17KuZ1W
MRnUBkPObIGXKSsaqd/2l89FXCvLHLYB9DiMhEncysmS4OSDj2bgLmZUwD1kggGM
QLVLEpUA9l7EzvwHzdxvzJVsQTw6ejjs3jfZo75OJYPohrGhhC6ZyHFpsx/wdl3y
qrawGC+H9/RS+h2VJyrM51kVOAleH8ge6DheuQVru1E/WpmdzODfrbl8YExj9+Co
Ziyu+9YE87HHgnhC97VwlqkTfnCYFaOZQWD+N3fWjFj1J0tKa/3tci/rfo3YP0eP
KQjVapvLqh6u0APS59PHq4hMsYeixMOVoLrY4jLL+CfU+HKLzK3N7CVh/eeGWVDR
ZXTcjA8Iv51vNO0F32peh336hdO33fUCxn/t1LMd1D3tEYDDdh3zZWhq9znJZWon
5V6kyuxE4dcTWafaUtSB90CQEnm8cq+THpaW3SebAdR9XMKNRpJvYmzf9VsA6gZn
wiIvIkMEJ/d4B6uTJp/lz60g3/uglBwEptRa0yg0czw78wLA5R7qZodloyzbrge/
i7aQ4y71c0WvKsQPlku1+xei7gx8lHwgTXeq7m/JLji2ZNtWLdVHXGCCpa0f4V8C
+mLAzpsPemgiLNzwGmo3TD2fr0b2eYL5sv53DXSWdh80Nn4uDfzI3uTH/+JgsXNZ
GsdDkC/UTG98PRWGCC+CGuAfT4/H0ipmI4eSihUliphCrULqzNW6rUg3YUUY4hFs
nLyZD+05/IVgzyXINntUUI55U6YAeDiCBdD/LZbm41HIRvHxFiaFSXthsMX40Nye
Lv7cnz0rnwtLwKC/RQIxk/EjPl2CINQRk2IPtUlR9vKDaNlGOhCxYJhYUGyhoswb
MBcflM4u+H8u0ptBp/tUBpaYOrSQWHP9/LSsjdblEJINdmfdm4zOsh9V4iO+PHsz
wF8YGA81kI3/eKomXHsVc/GMFckA3iHZ700ManMTd9iRnbFp0vJKMVI97wC3QglQ
Q8qa5WOyXt7m4LzvQReU4MOC6Tj0UMi0sdGGCGDnww0kNjLttK2Y5Vlh3klEknyT
NrWgsVmF45wOrcE3Y+ob+fd27ypT/2M6VONIvOrheBqWBclfhBS3oVAYw7/9qDzM
FLmB7RuN3wikE0ehiRqKmNfi1ftuq4gY4qBsSs1QBOQ1NNHuF3qn3OXtUEaGWbQO
GFO2U8t0H2tDeTOoj8cLT7JUZkW56+XSV+vBcJSXejdeTZjN9LwGYUlUMPI4Zh+Q
lpN0MZF94H6MRk4dwiFjGVhe1fykYdxlUsReBIJnF+36SneGrxn2lDeYMPPlsrMd
SgWky2I1uKjTGcD8o8aI651Zum9ZxRTA9AqpDiR0irI5rdxsPSJ/W0n1Ns382x3i
h6nTpHtM4/AHsRfoKonvGLqs3w1e1CvD8F2o8PuCjdZ6JO3NmwV+iIaL6WiJf2Oj
QpE68c7ODpvSMWUGhIa5+PeDIICnv7sfUxNmJwYs1HcGFv4Ra9M6ZfMfdGT/U88Y
plZ/LxF0LUrIemEnGPWi6w8BSwiT/FsVvqjF8fcInPUqoYzCAf3/cgfSAdBS/kEk
PzRJBRSlxGJIqKOzEQsR//5jgp0I4KxqrfZdz0eJf4fpXiqwofJ1E93GxMsx3ZVl
TVZTEx9ivZJPEP09ROiYFj+8aMV7juRdehwy/y5SbwPhTXeK5LMEi2mNHvldfkBA
3VxwMwgYa3nc+/Iy4DYPKdJVwsXLKi1Catz2I180d42ex/LXuuXkxsWWSCrXsuAT
se37oLF3WR5vfDEB6NSTcYaJqJF0wYWc+CVJR0G5FEcnKOHbb0z8yyQTGFcYCUbf
/FPz0NgXxhI75i7NeKZoDJhtsdsh3s6QrhLfexRVJNmPfS3vpX7ypQN0xIkKijve
R2HfjPill9FmMOXsOCyXzyNhWUqIf8syVCxh4xe2c6hcYorKg3akJXsuzxhWmzna
y3r6wasf3wYTHSEBEy46/M853oGRthOYZhkqUuEITwhGvXhYoTSLR6r7rThpPZQM
boGXjpGzo3V+0BXeNN4HPIefAfWWTE5acpCShFgyjx/oijhcBqODWtZlmfvjwXWO
CZBFakrSA7EZ+n2VuysRZRhpytPg0yFxKjyE8ZOKVOP2lxYis3WWGRC2SIiTudkv
Fe4MU6jZioINfTYC4Y9d8XV7Nd+V/N3yyp4GZqbtjaKLkDLP2eNYsMy1U2cbQNWQ
rOn+mruAuqlQg/heG+RhdY5Zdi6t4gt0Y/cBCKcLsQbqw6nWBjV34VDcSsDCDhgZ
BunIgCBNHJAMR5P15PzpD1ww5CIf4wLcCFHDfiTHebvEIJ9RltLsJwL1AX1qOgoR
MLtshjA8DVmaG4HRpef7VIYPWy0x4rcBLe9guGBYosMHieKx/4tEXP50LtC/3kFo
n2JoLPais/NGdV5Z6jceRg656it24ZEXkei0Z2TwQQMPi9PbM+jdxREAIaTFuhrB
EuGlOCBnO2gHoCwXRuIQI7kWbnLg7Gnpgh8WBF41uUc8OAA+fhyKyiCCtpVcQkPp
kYe/QPNkMoqwg+Drz6ROvxgp0MW4DFhHfsWpwY9NQtoxmGHWY+SFdt4hOzZbcqx/
I5+B+ne3nBk/TB0QyDNfI5n5uAufIYdLbSv+/KtDamyge6QqXSoQbt9JTFGY4PJP
WTDnWvt2lftD3tVCxlZyTg6gjPwfgywCqlFWRT0m5Iybhau6MN+rpxK+Hn4MY8zP
hTlwDqHqiage3hv5Sb41WGrqpKaJj1vRB7UII1tzRlldBmmUIDntoKoV0KoSPsUD
cstY+Jd2JV/fwNWrJy2I41zzOAPqbvqU7q7DaEpcbHh2X8ymC3mduIoIZieWKwJ2
xi8RUiwVE0UecwdCIqt9fuH7IxXYx1zlM8AVezZ+P5dDBeXeIwtAllFRgfY5GAxb
3rfo2mFTSGIYsDPuhY6wuPE+rq1ZWOZWPfq3BFXLOnLUAXWHZaCLCGJr3ezCISr0
NOrpNc1P8WCn4rotg3r5UuQbIPvhs0WCaIrm7xucPF06C3x4st833H3KxMz09Fsp
G8Ios1nPiwWy+u9xTAziMi1iI4XUtox7jCBs7VMwh8/Fr1VJKjZUxc+CEfKZBokI
ALcnInN595KHKJIuSXK1UjymsvTbAjvwPvG7LwbVl+O2xWcG2YpCxo9Oz2amov3a
mTDpBHETdu33IWJgLnM8BrRLUo+mrKEc9i9AyGeUBqnxDN+5hwRyuJXmDyZpCM75
YUTHyI3O/Uv5KpyKvcmwcN9su8FCdLnSo0V6rqdqgmzKRK5OYRFKakzn8IBGsF3f
PpfOzBsP+24CTg8a3f/EfB8D2bIndosB7hZbN/jRfLlsTns3sRVO0GwFVyOiUstP
qi0AWUrqt0tPA8rlDJrgRg1UiC25BlQm/IyRMnkmPjDuabwt8G/mh2oRKFkcIFh/
R4AigJSvQFXBK8bC9Yb+JNk81ZcsleTnw7+1V2N1tO3WPU6fgtC5R8tKjshgPImt
M0Zq3NnaZCh6LdVNvbZhm6IVHHRLVGrCQDU5RVsP7MpCDeTu7lziZjjatS6+5//z
AacXN61fUNfUxHih8/07e4Tfxf4LZ5/Kk8u+ix30OMfxxSr8GjiNK5A/cY8dKL9L
z+xf4obI+DM6XZ4s2ei0w8rkr0Ce6/jcGs6eAB/3da8TJjq/8aKf4vfD292pnFPZ
ZMhDUpMT6MPknYUAlTh+qTWnPaKedodFObS1MsTQMwxl6Xfx774mi9IWsKzReX1I
fzBEeeW5neuGEW2rZxXG2NTt5JcGYX+OLPu3bF9T2VTT3FhbnvMxKus2Ood/BphH
yGvyV3SibDVPRMO9F7XIbz8YpUQVw+6PguijaFlztd3EOFlv9XINZhDP51Wvb2CC
hSk54J/8wnGtLdVq96EMQLiBZNLgHJj9n+BJa3HUGzu2hp8FnlW9+1VyzNMeD6uX
m3QZud6AYMPY1bWPpsr8MuFQxaHhrAngh8QJuAXiOyaLckz46NmiHLMM6RZ2BM1W
j6+it3NhwfmaqTTdI5N5fukOVtkj7DxfgCZgSvvNvGEJNEbcIF1XQqaSdAkpWM6Q
hU445r1l0FhIpc+vND74++ZxUNaksjcdjznyCZKVFHUl0oWgmmpWDf+h/p2NjlUc
ITPAmANli5xycN4v7NcsQD1eJWXGBUzjkTiIs7wBt6BohSnW1PCEJzT+nyUm/D1F
1PTYMF3EDMTFHS/+c7j0WkwV/U+n6KNia5AzqXQmSvHfpLwoeSvNcIzukiT8qwl6
dGEJywfagv8m/m/8IV2ee9/V31ic03/Z8xpVROl1oGiNMvwLy7Ws4bHeOlqCDssU
x7uFWArOR78z9ugXuBhPjX92gurSgmb81iGxbma7Xp2v/lNpmkPLOAibe8arsyK5
9dET86sGbJQVxC7F+1/PvEJlLQNXFr6jolH9tp6Rw01tB6WtUZr+cA4nDu0Gg5NR
kF4mK6JHCUkwOYc3pRDqpDkUbMxU51emc+Yir112vuGq2kSytRn+dXnNbh9gWEkr
a98LDn+nEeM5P1ZhLxZiK8p7GpHjVeuIc3H6YaRQr6R9U5csn0ZETtpL2FY3RKd1
ezT6pA9uuBohE/pNmBv+Tk7YyCbqxXgCOtPqgf4Rq6OgIev92fajbILiI1rL1EcN
9DFaHqnNbGqVMXI7bviN8PNVAWY4Oqgc0gtoo9vjwVkg8q6qC+Off2/R9ns5q8Y/
Ek3q0oN4qMjUzhlX1l8JvPxuB9RHictE6zkFVBFKTCyrhRJUMh+zdOwRn18PehrH
l6KX4MXHWmyEte3vT24bg4hGbxfq4f36YhoIiS/VJFyn4MjDeWCjhm2Uuu4I3pJq
77U7lZW3NM0/xZnZyPZY6cfcwwazi+LZK87uiEC+MvWyrvg/lOKcUqCRQ0rcJzqH
y2rAxJ56mvIRVYkZ1RxzCq5ir0r2GiHnyr8UM4AabPqxts3gj2ne0TMODclzEHCo
N/8ZhsDpBj8pBKDy1GuxG3vZF5SverfwM9xCUZbv4KHFjjA2LuI4QbugQFNodRNY
+p7A+OKLINzwtR3zF1h7QM7dmPY5ZsPPIuf7fXdVVUCOiyP9VrP6TACB2xPAHXsm
vD3/mLjY3yvAlMKqwSAH73sX9g3vdf+2xSGBvxMTZWC6cozFi+q4YflPIZ9j+tuJ
hzb4Ewl4V1cw8JWeyAzVIvMCGOT2vBENfdyUCQ64A0ZXdzEysqJnfpQoyj/PznrI
AoWWIP4x55hKTXSAl2P7BE1Ae6VQAxERF5YxWxBF4QBMwIKqB11E2m0H+tsOTXiX
ggxwG0iAa/1G1LpmGsvBa3CQKMVftQLR4MnGfK5w+zVqMNR2IWkni3qGVY5KTT3m
WNyBAP06sgIcWCtb5M29TQD0I8ZQG1hiJC1FVir6TIWwkLbDh+IQR6c0q2i1PhI0
+JaGeuhmVy9gXG9suT2/A3mE+fe0JkRMHtiSBdGjNUJHKAkQ9g6pXqLRnmGiSGWo
Fd8BiNFyZ4rcDNv/zLiTQPOQVD7d5Qg/y6sno/OLcRIKUw8bZGMoRICg6S8Ebox4
VREq8wlSj+io6SvGgodmj4/3RERCavW3pTW1HGX+Jc+AIKwyrkODMijFJirtBWZD
H5rxApGBJIJ3IMZXPpTQ81ePRdmUm2ug5PoF9u1DlmcY0AUktq/WeEwlI884s5sZ
g7XNgjC2ZX7WvpwEUzg2EjC05gLwSr4qaq2o4elZeWBtpkuz6ZmhhKzI9cI0sIRu
9GBl9BZEMq43CHpw/JfDiXTesuGrVR8vjpBZxO8zq72QrL3dVm2iFy0b40+hdH48
ePpaJft8pSh99J5cFe2MW6FxMUXWXiPrtyvkut4qqdc+uMUvIKxRc0ZPlylgVePP
NqH3XRdIl83kjZV17yJUF8O9CGnre7aeus8sIiDCucE/Ufncf6/yUq+xdqkwDkoJ
7n4Rs2uDiEIK5tpIgPutsSRFLmZVrrq2TViibmV5Motlfyb8k7iZ9H5wx259igyD
COBqahR4A06UxDFC/r53AGCHlbAFVUpQJlKsHvAnFaNHciC6n6CyB3xKubHS6jLO
85oRo8UuzDXXzN6/OAqPeTojoIO4XHtdhiPILW0ARaPXdj+nxdxy61j3QMA2ZR+u
5iNXyujsNINpE34F99rSoYrpcReOmydGV/It1QxM4cnF3YzWtBNzLHfRJFreuPYh
qDyqsnXcMUttbzaqjYO4UDU5hahYyedCeglMqwhTOrpranJ/7CZzL8a05I+DCELP
aWAi8VapqKB/1qw7p7ZuaBR6QAjlCQvEww6xOdAjBT3EIgI1QqYm8QLXIEKR4+FX
YoizVd+oeYbRY8iB2w7KDy6DWiP7QdXClevXha4yFWZ8HlDtoMEMAqb6IPuRXSOT
Js7nSDQ145Cxxp2pdnMlS2kMMuWZPKzHI/T6boSOjMAEDySdsAzlVnP+7ccqUrld
6S6JQ70YfRKlaymi5uwpPa+Mi3YX2G0x4VYEJLfvDR+AKaj/Z5KJWaCUU53yi6+9
CME7+utGVyguCdboZb4X3QCe6FGH9sdRsiHldUstpgAzzW9U4fYD/6ojQbwqiC/G
k+dHxbyrrKHieW+1OFsl21qUK8S3YeRDSivabSXUghs2E1DEmNNcKwBDAVwXEW40
q2B1/H7SCQvDg5XfWoAsrHcpU/fKZV3RNJ4zk+GHOWyNf5j3ULKzjq4npFMCEJSt
v5vThV1YAL8qNasZj4gF3zBMTIxz9kp6xFx0z+YjCthnhjmNJV/SJVoNJcq3WKLM
9/yp+7pxcsGwrlqWEIhX+rZDEJlYuUp8DyPQ+DWTZKb2qrWkiD0ieSeM//1FijwF
dUDoeog6dOZqzb1pliSsSbW+R4Hz3/q4WOo52Ju/xv7rGu04EK5uYqQMcsTl/GVB
fqS4LBR3Y1oMzTHMXzkWHX2TnCT6rcC2IfBqP0Pnl/cMI/Am4S6/0sInjwHtzYaC
jQtbM+dVMq6lTEv42QM5gVOGrhNzVXSV84EcTIyWcV+9IiJprri47d3bvkD3jSt1
mmjVjEUaToazqfQO0BTxNu2MlQ03pPYo2W7RmVLRFfNMwvcEyqQfmnE+XwxR9sVm
YSJR7VXzgaQiiSxr5Bm7fVentHjdh5HP1GftFNTkUVfzVQ4jsyuy5/OspM4aVY+v
/mv+fwqi/e+IuqFct1tRkVz6DdADpc++sXY9u5Ot8uG4JHdkFeLPzBZkOAVOl4eC
Y70/sFHWBgOOFjWqHXy5DMV8+4RAJqv2zFWbmd4ZOltQ0VgMpv5iRRh01ElrWjYv
WxYGftglX3yEsgIgCtu/zC2cFHHjHnvQDKpZwby++odz7jkxTa0Mopjb/ynU5jM6
jpzmJ0hhII//KG49gO593krp6+V7Bb2/Z75aFcS+2PK9qD4vAxpT2ZO6b1Dbk09E
y7KD6gCWXTP8TnJh8PZGuYJA0LiicNqkJDXDgVNsOLh9hYNAzv830fDYOJb0AIIs
JNxU7n/mUcCKUhPOGmHQKrY78fM8ZWXaSxj+3lfrH21Dko+tvQ7XlxG5nJRGreo1
l3ve3ImRd/HEv14K3/qzMSYF+md3xlnvVWemQcrXfdCjXGKBhVUCWtOT25uR6a2C
KpGAzxuNa7wa13dvfcBMEUWYoJgtaYKDftJIzMJ8flCMPPUIIxhijej4i95m+u++
L4nQCT8zDIhfuHlD3KMYITVVMhI8f8aqyorPx6qoUDEjjUc4vWwZOV2JJaxVp1wk
Nh22L362AOsu4cI31ktE0pIIXyJlM4BZIWt8+QOZBuunk8gIcMYZ/h3QDLP9rHYC
yVnwsUw2Y/OxF357yoMcOTBi43M6z5bMrGHHYAYR2QYFKiVFXYJJYXrrV+9phl/i
OE7AZhdLa0CswTS7Zu7M0a6OFC7LORTTAt8RKWOPyL2FV/1C+TGT96dM39IMe+rg
3Bg541ICEBbM2YXE47rBp2hd6+y79bZ+KsUGXGJpsJWG/bChJ0EULYgtwY4/JHXO
lNe2jIqn6h60cGJuSaG3PwdoVGLrmCQdJoX0juakVlhWXC1eQ1ZjNLg3u+yTfVdL
c2ovrCVU754yiUhqltw12s/Yo3Qt/uhjUlsc30OVLiJ5qt074Q5XAUYV90X0OGJg
1sP2cPy3G1yLNs0rePa/kAdCQ5Yc6gnnqAL5j1Mhp0AZAoP+QXz1nOQp/4ZffVqe
h3PTzghLmxoZuYieQAso7k4SvQYD8jHVxd32hme6ZCjcwaMOuzKvYovjiGAKUGya
bz35oTvreAILC3PiKkX4j4II1KFMCx+Z5mlnT/BB380BCG/c24QDD4csVPzNG4M0
LlzO72+tGlVHlRgUcWcvFpK6Ex4jet5hQO3/Ny52pCbjWD5FoHuEuh9rFQtmbKEA
R4Gj6y8RckmuhVIiw579cLU4/SNPbvUgaO2EiWdLKX60FSHg/vY/l4mP9cFMTm25
W/uw/TP5sKBK0qeeZrK87p53tFkk4sgYQQmlhH16+vZg41mw0gGh8hnMKe9LvlHz
Hg6gw2+n9JWXFxxvQO5n48iOhEcLQkv83YIF++7XWGICxF2UisNVFvhr+R+EHUJG
REjLRTmSoT4sd1npmMJpw2vQN8+kEmDdx3YLWOB9gJvFQ0K61s/fOkktXrsjUx83
dUWVjwCNRs0+so1jWYkxF1geFr8ANSUexfWULCsIzwx27Gsuac9aePlCQ7p1ZJ6j
O726jzuwWnBX+6ei74vx+zpfNpwoVKffyy6uQBjDysr7pay1M5mJTrgTAhC5S7Qb
3EcciqYy233IUQI94e9VLRSmaUMkxXGHrizrLURK+qD8e540A9X5dV4p8HFwaJy/
QPB4tumxAPh9pSabvK+PokPvu70T75YgPb1eri6HxqY1+z1+chLh7hHJwOUyMRb9
XZQ8xlrd+T4rCvQpp8EjiKhKEs0lCiTgo0XaWdbV37OPefpBhm/8RLMznHAz/mjg
NpZ0yVAjyBfug7EPndcVJHqvqJ4C5Rk5Pi5vNhbf3JT6bk7SuWwJtO8E6E65b3JY
0CbrwhWluxdtxdwEyCgSdNW9Fe6GceGGGue/edCHZrWR4ZkS7M68F7N7MTQ33tx5
zuW/YLdPxSJIwDkxrYCPcWEwjJVXXgugnHU3L0Ff1P/IUIDxDXkJYepiddpMzHzZ
jS++XY2L7D1zJYcT5//6KnzGkDwnS4sr0vFrKCtY7jayTcEKMbZBqhanjf+BnJLA
fLdkVpsdQ4uuoFu9kTm7oFXM1BfMSqQ7ooWdsj75O99IhN0Rbgp4jULqFzH1uotT
3v6XDYvf3cc5KfeTUsbQD5xGRm+T4TiW+Ke527BVIvN/o86YVk1WsMpsQKUyCcGK
YcVqbrq0yKJMaG2rBpny40QIewT3dvtYPgzioPzXewKhlmg7XWntiIdYg/VnBmk/
0BwsxLOppsG3GI7LcbnXv1C4TF97QW3YkfB/jWj4Xr/I3+hPyVFsQ940UL+jqjKs
d83LzmrbK0dBksRiXAvHxLnyzWYsX4JT+Rf+lhP/AFurSuBlwsWAlflG1HIgv5YT
N79JZlpdxFdb38yZ/6yfCRUZaju1iQ37UT7fexugt9bH71TkERo5XTU0zyHhF6nq
ymGm8ewfg2I97x+QshpZn8Kyy/ZazCVREGv9Zc14R/RdCmmzje8YNC3AEY/5z24U
crYQtABf8EjYXdOZtpU2xcd0LgJEHYkUTK/C7cp3N2m/rQTPG2/LP9sOJPK+6A/c
qYXNG+5lmUQ+uea+0v9+9PF06AEbMMLcVTIMVqjdiOXINYaqrsiOGVKd7w0UQqNF
J36ZBd2Mjp5T3yEZKKWlWNVTkQQ4RoFx/xry79gVaIeJcNQH1tqmpjACaJwPr0uZ
sqR5f/ZVd3esoK08SUPRMGm4ly4kx5GsDn7lfl/nPPQ5XwGyFVVgX/WzZfWOaKRR
bTiaMmlQZEp0NjPtOUzW3GdWJXAn1pV2y5n6Jcjn4XSYWBCjZKZTwM5UuFI9ETBF
RGy7ts0ezrKV86DaNRD9AG8yg16m5JjD39sO/v2UXO0NEKicv/rISu2DcPDYyRiA
D+qqDAI+piYrbYuNfBFNbb+l+0cH7HXZSA+BptTDAeIqnwywxmKhRKFpzWR0dk7O
4VqxGFWXjn1H0P5ZSliODKWyNuwZBUpzwjbSH8fjg5M+XptpdJwqdtQJK6KVrW/i
/bjjKzNsn9y0UN77AGTGyk4IVsPQUSE9y+KhcXgL69QSoGEybeWNUDKgOZ0wImM4
4NMaiK3IWx8us2VO/bKUpUKMBXruTlCXLfdP1xvvQemxEHOiSHIO7BETSM3ZOJDH
o7i3p9LBaoNtbFXPEOFKS7sV07MTKn6fVSh6YUsI3Ja1xu+tNJ+h8lsBaxKv3nJo
wtwKwP3dQk5oJTAmvezJKz2RjQ8jnMUM8uR9W3knNG3RoE+YG9aEN0lP/lrMQ7nL
Wy7GBySYq1R8950OTBi3LDyHEfkmBeL+GKeeU9hxCkqsQ5UiExUn7abukx20sqWk
6tsyOCJ6lPhotFenuNcq/l/1rRw/B1P/eTJiftpUhV1dQVS7xzB6j6zzP7NvALxR
gwYVfaOaiKRtYVntoxvHYBuKlpHeGUmd7t61S1oMKTb+sKdfDO+l4XhgggPb8zMM
ZEk4kT8RKZixauLborp2xydXl2gz4Pltm+/CC5WyOCrCpTyZ6xgEt7ff2UWr3/G2
O03LlcZr26lOLZ412ah/bcH8WvP/QfU1pagBoGbhn8RINxEPUumy3LfwVkG226rJ
EWAsgCzKXJtj9fvQRhI0EQ/sjnZv/Zfk+W3Agq3ERmhOrHNfl/phnoeVILtVgoW4
6jUJP0oxts3o3MU8alLwHKz4gi4ETw/NcmcqQsLSb7uOkZjt+AFgpT23RiUs4yu2
1QmAFzKVB8y7r8IiZzYKGigEKBySo52gG9EC7B9zq+gOpqhRJzzfttw3ylAaxdvO
Zj7eCW2U1PFhREfcV+w9FOFVN63XpbR+MQjTzy0VjeEIG8+6j+mDAlhzxuY2E/pT
ItN1YUZirMxS2OmNYST7GLLmQLAiEZVtoRFi3+541XOiBU9RsiM+YBbEmdCFlOG4
wUd7tOdViapDwuGhfeyX7UnsPJSw4XyAmY92bS8JULWeHBWQwWA+C/yb6plcVi8E
CWz2E629+t6NsAGzRkyr6ORI4sqMO7xEHESgWvx/8FccDYo76ycyh4WE2JgQcQ8I
862HaYLPn2dq1xlbsZjeFxNgMNVgbB/oICuxjB6PP00gdAIKOyCKljkFGjlP9R9W
K6WYYcpU2ZU61J8bSY7TC2xDcxVzkH1aAxK+DjMncRLkSDQxoNkF1I4MOaz+qL+K
u3DBg8IGu6AtaqwBKGJYYizderjg2DjfU5N8hq5mvVT5/POYf4OQXzqZqH9rvmtf
jhVwdyeKEXd2IuK3k1DBtBvhxsW6WhGjc0ljsSVW2KK/8dne1ij/2zLAlLSzbU0H
eUDhPAHOHz+H98CNsXDLNlugpGzOIXIM2cUlP73L2+Xfr2+Nqkyd4Pb5eQV2bUGj
funRDINm+MnbnkV6jPYp3USaqOtVLSe+7cSuZJ/cshMqynCXuU6GVrDZxAv3IkuX
fxNyOlijUYyJwa2XUT3SNJFVsBwpHOvtYI+6J9GdFYFFuwpBxhGrRqVC23Gb1MR1
nkqvC46frfduurRGlK2H1DofBZvi9S+RuFor6maEQg4nq63YXzsajq4yimRjln1x
gBdTjNiLse5b4HGVo7cR6vZwsJvTHQMf6zidu+rkCozdtgcj0IkivKoE6ZAf8kfj
RlRgcaHUGS4sUVQ2u/7akO9hs9MqrfUACP8aVbetoUg59tj6ltGhA4laDgSM/kxm
nDN/P7xnVHBPTmTSiBmD9geNzncoU+1hpewLYa02UjO6fRfiKa13GubZCeW4g9Bb
Xi+lra7tkiZ+s3oN04juOsR9Kg5/kjZd0e6JVtrVkpqLRCJKVX5Nh3UzdHvOuV8d
ZWi2Gis+c80Pm+SzUyZHU+5iv0/N4CZrjV7zMnZr/H1taorbB7lTizlqXAcBHGrf
ov6+wo8H1PXTHdzgTTnM7ThNxir3znVeRXane3pYWZDW7DWLPR8Mr1CEt8E9tUDs
uwJcLdHmJ1CTQDSRcnQ7ojZXP7L9L8A59hfSESZIrtlD1ZWlt/LHCYeBiOHU2q83
GDZJ5dpOwp4arvfrnV5M44wBYYMoiWKiFitGd50LkAVwlsYb/qnfOIy1VH5OxJXM
GsQsXZtEch3YuTK3PYFLZhCBZCOFtKO1BAfK0rXkgfa3o/awzCJZpVuRgES0cHFR
W52gwb212jcUXZ2iyMgxHS+NekQt4rgVK2CCDioUVlLEY1yyL+lFE8ZCrV4XkkHm
Un9qQMCkWkFd9u66ZqeogrVS4qnl1t2vD2reAtQZ0CysGKp1DO7TNt6DTFaMHMSn
8DK0Q5ApbMBQ5qU2SP/Ioxk5vSX0t762/A/hyjfsKa+hfIymRxY65lH3D3/B3G8g
fVGXHT6SCBQ22p4WTT6O4AX3mg+WR9onyJfIi59ATVY3eEKAe+MZKUGDfPidlewk
KhAlIhV6s40p7SYBsRXYDKiQeANWeLf+uL9xqioUdWNqEWbYLo/4UzHbt73FMmEm
X57PTet1VMWMy4EFrREwPnzJG4DsyR/+kMKD53zwVy4kcMmsS1xZpjlsSWuimTsf
W2bgp5riD2LccK5bbudujXWsIea7XOoGaHDxEh+aWaEKtH9QJExd+bUX27aZV3q+
edv2hYaaRm/H7rR/nmN9hv590b+owyVaIs2E7GLmgUFmjoIWtAQkW9CDJM5hhHqZ
0aQ3fQlrU/t9PpyuvdRCH62BpaUBT0EvXOopPEvHjvsv5/sWMLrEnAXL4pLujEk6
8pptefHn7X3Id7tK8oG0yfe2C1CiyBUixCDGsnvvjj7fA3Hpj2FLA+HYMiEIaQGE
Yu9im0gsqLLh8Pb7CzC5USYV53LqabhWY6AQij7vlYYvnYfs1G2eOmK/hntRhE98
Aa9uSAV+1wIHbi0jX4mgwoZVCSXNYvaVWnVAEj0LoOSvWH/xMpdxEbFZvMROBjbH
DorrGYddZO285FjrEELQmdV7HpqLeXvy+agpki3gO3cjcnrzFgnfcqCm24B9yjwM
/jlil2tdMKeCfsEP5/0F/qtcVIqIGcrz0OYrjBBztbuNzWR93wzXQWItu/a5ngx7
OGXn2qKboLxzsaZbN/uUSObo0PfoGHN2b8gBrgFZ+GHgtiaJlf6yraONVelAC8JR
9f5PMLhs4ICH+eVXAW2X/wnaL3ujpsCF/8F8N6ytcaM//yMAuqNWd6pollo3qBsk
cayJMkTQl9CT420DQyqI0eyBFXabUO8EuGMcBvnpHhK29HMsBK9MOZ+NqGGTJQW/
O6NKiq6bKY+v+tYW4+CfYhDTCjlT5Spyeu/dspKTTwOHyrww9nrr5HGSPqioDNE3
kqch5qJ52DQTGLskbWnQzmmKp1aDGtuwflAY7T++MScTtG8J6ARELzHDZIeVnJ8v
tUVjL8ra5BTeVO/thhol3bqmYe7mNmnIcFMmeEQVMrMn/5z7FJiClsQVwF9353wf
Q6EIlPDJRgSRC6GPZ1fG0goIpt4fm1wE6+Aax7vrFSownE7AgIwB2zml+JuJnZzx
RxntVe5uTvWEdxPDUSIS8jl/c4AjeepQPEluM7vtlAQ5ZaIiMy0hNR7Q9An4RYuS
VEZLSO/1hFtYNkHAh3UOczlNCNRvPGAys/zMuK0ou1i+63TDTMDE63Vw8BHlxMAX
QT5wBTAJ9Fn/ZUF/c4VOHc7CMDIMEo2xFnUqG88tbnkYHSDP/Ns+ZioAXnMmJdm9
kiDkmNdqU8flI22nNqT8hfQGTAl0xrnTV+JGJc7YZrq11HZzn952CjmGvH2Hiil0
etYtYG7OCehWSZ4eOpNtYo0SMfV5aKzezVgrtCAvgaIBrCQz72qVQMO2eIpahiS3
S7UeqNUZKkyFIn1GPnINHBi63W5QUxYBSo8NnLjZANswaRQCn7KerBn/BVSExMIs
zh/zKOxlsNdE0KVTioNpKAKC0+sjdvIBrRqjEjo2u+RAXAwgjS5wBLsXHLr0c5X4
mkRg8ySrQXWtcwiyisxNYDi1TK3NGSEhGl177ye7XLzf03BHWyRLHAliVm1r27KS
mFNwtI3eP7tNZ7+3PK8/Vrkl2rBKATdWtX1MF40YR4VqJOEEsYc4z5697o8BYami
qYQZLCfOnSJqGB3qoc31VOmzPq6bS+JVrwoCTJkc0sFOvvGMONThnCQSRl3Ca0tV
IRYDnVwLjQsLaUCocfdhhXpi3QTiRl1o6VDIhX8qftfdyJFdCx1YNStF6LAx9ylb
wt9XyysaBrvGhYDc8dWRTP6FX9pwiaT2uMwFQlKcByaswislTvG/qjE1Y37PDHwF
w5x5aHV7l+JPPgQ/eC98WJh7DPzUEzPbCUa/bbB2GBcBZAroaBbcghT1UNFGT9F7
MSQNr5SEE18atWaTJnw5ktA4WHwGKd+s35zbvaI94RiPEd5KWLVZXEQJOlYYb+Pt
JGtYdGYQj09BRjQKWupRWW3HRjr2/t8ko/MNy+dVP1645ufX3q7B6G6yF+0foSfY
6AdGj4u7WUibTkYkrH44aND2GOP7/TBl7d3xLIq5BNbrqc2ueoFy6NUZEvlpHtq4
AoAIyF/HAL/EkqE5bFBK2FOLYLeEzq/a2w5Wrc+SoRm9vivblmYS+10AZ+lW60vN
O/pbvrBUAz2Euu7XqoCygIO1/UPcjIudWoK3NLpa4P/pJDf/rr0A0RzIvRIyIaYP
mEMiSOOw2EhQ1oK3r2xRwV5qeJ9QcJ4ZZMlkfdFq21b4bVLyayzIQu4JcM+pp2+b
nACbXaXLo3D1EuySWRrLcBilBc7XoWzIw8FUXLRka/16/JEvIxbDByPWSO2BTMAf
gPopzEOKhsu5uuLop703zNH5CEaOtGDRG0ril88gFBApoxIABCA9LeuHZSt8d2LV
bARqyPkSgpI3tKh2wKY/IpysTPXcPWrFmEchrRV3hPkH/vR+k/64TdTiIaZLdb4w
Nyugh1hr2IW58p7Wgbr0ijobcbLWt5dEuous9f+Qlo4WvvFs1t8REHkUV0isMSff
28Yeghh1/EbBsg/+jHAQZ2ByjRQWVPIgJwgFmSJYIqidcir5hQE7diunGTcSOstw
Bvkc5Mc9HoI7GStgegB6pF7DvSbrEeszjp2vZO9ngXiJagUjW6rpzUdB+IXWolQx
HYcxmyTdLBlloZm3P1QHh6okm2CpL2v6cWDPZAl9VB7FrDbScFrPexR4cbYuKI8u
TSdjh8Z9UvidlrGXzBp6iSYZytrDSEnHlCJje0jWRFX4zr+lZANWm+92A/SLqfT0
PJk6XWRXAd/NrWdMqmFpqH/ZEBRajv0/mhi+TBOKhez9k5HiHyUnTgYLQuUJGmaO
3UmD/6S5jBiTUKb/YVuJMZ4FiHGRIhfKprD2Xor9Qt3S+g1gOG7NCXBC4Y3cKMPo
/s6XQ5cbGbyng71qeQRQV38A0MjFy8fHXOC730CI/4Rbfsit/I5BvkmuguXM0JMB
ENJresmqPqcft0yeYblZMUvQXs766JD0Bvoomq4jANJxkxGKujNelGEgbzLZTV7l
WFIQ+PmPg64oPk4Q1kzOl6ItZgbTLhUgKPcxMZ81ceh40ugiac+lsE+fsETekFIL
cTXWRxBe6H89sRGrTpTQy7vS+Pp9lxOR57uj9i2zXOj89yN95mS5duOoGxdkNaJS
K42Asoj/VULLn5em8mStTSlwHvciPPBlUxUsZbKh0C0n2WyaUY77HTePLTowra22
XNSapwoI+3eVuaKiZq+cSh/sgzxyzV0QaDY2vDnkPWu85IxDt2fqQyEMnStTgkx0
jA67qp+PhjoO9+HYzH8ATByRSm3ufi5rJhqNc9Gg8poCsScudFLLKcIcrkf3CGKj
+TxpW+S+4yJ0QTTYos4X7O3+ng/r0yqiZ55L/JULN2cbQorBeRUdiH2KZRf3x267
jqvuwSl2cLdhv6MKcYtpZ89zLONKxIbZcEaUdoOgDuRs9q+3knTFdcV0S47RUl4h
jvu1QDbQmN3sY+qtOfrJLizOY02Xp+TGJO7cGxIQhdfMJADjmesnSjN4kSQYv+3Q
MPmWf7yWSNf0mrxGkdY5cn6ZdnLMY2BqfmT0wFnvaNffL4Tg7a74hAYtRzHJPFix
3HegJvAY3vK3vb5fFsvABsbDTT89H1/wa6Q3Zbgxh3fz9vGAK4EVCcxDGqvAOAbH
RTbtKPWrI+52/3q1IH1HWFA2f9hpSNSdqoqW2I9tq99PHwt+OaRsMIqoOLAAwUtB
v7lNFwN6zoHv1TWRvpSjDLVPMzGfi2cB43A/lkc04Bebfcb7vkSOupkn3w1jhCPh
dPwDWEuKRyMQVTTdj06VzVxpoyA0bIdjbAuoslPa8SGhqxrVR9/MMlvfVFYuJjBT
a1pWL3XCxmkEjysw58jILcXlH83XNGIo2Ui4RP4Yk6zLJc5YK7FJNfHr8AEHrXsz
q+3BP53XQlMw3+TL50tppIWFhurBPxd4UqLrDbJF9+vhUavslCQZBET42m5kpLi0
RAFh/RBfc3hGXgDxU0WESYA7lYRvQPogeD7C3hykF2y0mok8OXTRdWT1UBh1MuyW
sGJSxcRs65oZqXAKk20AV7ji9kGSDpW7oH2kzZcvThc=
`protect END_PROTECTED
