`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bHagItjEMc+SHSGmUlBZHLh7YANYrhU0Gl/O04RLqG5KfiV9A/JqQoSI3Uwu9uYa
Xebrp+nP8JhUdeW9c8JZiKT4BzDRfwjH9lLhMHfcqb3u8vooevQGUo7nuNwf4bDz
0vlIaK3hWTa9FkmnFyQc1zMJss2jiTKWNYxcGyiMbS1MmXDrEUmb5SWZF/XxLW6G
UEtC1f5XbSnzLFs4Ewqbr6GW4zphPpfj0ivcN/8EbrxtpNUz5O2SYHZveXvOOA8q
qz4tcWInney02DecB2OcNnsZs1j9ifkp3lqs8dHVl9gvaP54B0WFGyHTf9xGzQTM
Rz9IoRGDX0noL7tmTiVsxbM2LGKawv5cuFQnnTs7HliFf0uXDysCDa9Nes+1pP9J
344GloQI8ZFtem5Wggt+kgtaSZUbB7PBzeQ2YZ8GHUWYLnNboRRGmbkgMY3xRa7+
V3poWwFUGN29mxYLKrYplJyrNI6ziDH48/4LYtbNbNkIThYSOzBegoseor8tM8gQ
50ZazWTUq88Yorv7evqXzfaAix4tpNY8Ozd//hFniseuuvh59mGU/ykF/B9kp4E/
jF8dmQIaTuHkaONQwXc2ImNSszYQMVwTdAzpibASzVf08BtTOuFuvlqmLYaSDWsp
5aHLoCsNOe+kc1XsSleq8ZvWJGK3edrePaxRej2XLHD9ohNG2c+VhFuQ+9t9vnrK
DOt98xO/zqn0n2aJWRLzJcjFlSeaoXCBsPYTlygRmySv9Svu1oECDksIoWhOA4dB
jCK4Ka8DrPQfk4CodsUI/bCa/1Ig29gg93wb44J0YhuBAgD8061TblISw9pbKJ8V
FRz8esJp9lZCQ4PA4OL5TOA3X7uFezzIyq1C5dyU+OEHmUUgDTNm+dmyhhR4u9/Y
3KNioen7VRQEOfvzyvtble7YPLtTLpt90C/l1A7V2ha7ABX6pxkEB2wlN5hUawJl
OAGn1ySNfcyMx9qnqVYEsLx6T4TMfBfjzpU9vBZi+S25oUInMktrE9poq7Z/9Y6E
IEz579wGxYglZDd0NEQAyRrulLLpD3wTIScoBu/parr3wkfjTWhKXCYLp/6GTADB
i/Wy8IyXWgoNPFFhD8P9JAX98HAvfgiDRUFNmxe+TPjBDfLKvhv3FlE1O9Ow/sqA
38e/xzsFIdkxVrUfEhF97A1Vp4P+SATbj6yDHowfgUi1Nx3pEuSWVjc6XhAmHUb9
lCNf07up2ozmaH3kZgIaIZOCzJdqQsWmj2ScuGUIm074zbHmNLchEZSCD6dfKbnb
Ks0CVyM4xmPTr1Gdx/M/1X4dSKRsJCNdUMDbStcG/I7uQExhz13sYBxxX/54g5DO
OCSmCaDpbCsFBALfEpXle4krM2QwTRGBBXYZswg0NmbQJ/ogFrQ/FJY+UeEzur6y
WICItXGYK7Q9wmrn6VpUU3HJqNj69LmyeNbqofREFlLFdtug2DCI3mf5BTC7z/vv
T5P5c5yRnZ2CFwNaWKEPq9mAJ1Gt3PSNvtFDMqOQa5SRV+E6z1YQs2hSZXog4T4H
yWc8z4VuugLffMQh2bip34w6dtLg3stJt3iwomnY5tYBJ0Ol1XbOX/wTQOBrIiTC
k1TZRrrjIc2mwghjT9Dkcg23wHMoYmzSOibaVgsKJ0AnmfQFaW8yV1Bd9IxkGSBc
tSLkRY5iQ9gZZKwT4Ic1Kd8XhON5bUqoiUADxRgdp7LbuZQnAtRmcQkRvGxK3CGM
vjLMxitmzIzYdpyRLMEfOhUOztu6KYbtECAT+HNisK8AHYJHVAolic3UMtkOph0z
j76893x4b1GRp9eNRPdIolAcZmSPU47jx5eDjbSBVU4/Vnrtq7aPFt5q68xIEdDT
WMwcAYStDOyWif+zLT2wedqAuncpNk8SO9mbK0FsKNRfDeGL+1QYRDcLa/IXjgka
kEUJqQNIZwq4gmIaB/dPJmJzHG5Q8vqo8a0OSh7zUXwdp3f9PDXlwDDvpl3JB0mh
XfpYR/ELGuqqnmTXlAOD6ml6zs0tqpM9GgDyTTbm0sre0qaOho/5EwrU371tecpA
k7s4TGePZS7UG1h67WAkLndv7QbLqeLb1cGv/Bz3sAfyqSykWbFMq1y5P27rfTdJ
9nkEmOsONmSgiM/RKi7qmD97xiPmnDdnhru/XEYSAogMzLgdG9hq0BnZ89nOIXaN
wR3g3VpMvA/D0bqjCLHrBvBbSqYAvcfkH7ZhYE6/aAQYl6xThX4lQy3VyIsQhgfx
r3GYOgqezl8zyNl67qxjcLVgNx3G3xvoqi3G3573xZysZmkO/UnsnlufXQrj7hDX
ABb6jqriUgHY6KZOaErnXhcpLQc8JkAmEDR4hhyYF4huGwDCMSHmEj+MS4v3Kqy0
ZRCqqLcYVjiC/OGoavHT97nYNTPtTCMe56jZwt1JpHsOzS22aYRkgiMYs0VmR1Ym
KC43PO2CyQk7Vfkpq78hvf/adZuYqqRzXNEE3O67Q2fDCkxGPqHcKAsR5tHyltZI
+Sr/UQKtcoYTzrNvf3xCAhWJqr5tPcQgORaogZKlFfheZre2CSW0cGnKettsZ/X6
EIGCy2JilRNWnwwB8qStTLrMKI40xR7vg/wgzjGvQHhKviGl87XoHwoUmLV0vlmX
EXreG5UXys3mSzQyCdpIVex+6SSZA2k84M8KH3HUgkLSVLv1sD058TllL25r6Lpn
nQVMVIHs8wifEFWA/cKV58cJPmui2opSdIzYLy3jttJbl7VPiwF8wuk7nvZe8Bwh
U1BAoS0Jy95Aja6prcxDCa2Y1jSvR8BAIskj/Fxz1tusEmTNbWH9iyjg+CXhqBQ3
oFy7b38Yc/iIuM/GAVyNs9BSaGjB+JjkDwr/OLopxqnU09fQXKzZTvyScd9pFkif
GKGU38t0HYuOx4NC9qSvNIuySGLNz2y3T5WgYgJQu1Ydp65OfZ6D+hb7vUZ2nECS
Icxm/2lNIQIsfOAchxbms2VUimVMfLFoxSyYQSlrNkDwTt+rFFmEoZimjZpPmt5Y
lFYj4xbsW7WIc73+AwQ6t4NOQbHKWQJjNPyKATDXwZVDDBFZbAntrPGIkI4vC3MC
pbt2pWX/Oq7pyLimlGF7wigbOxnc1c7AZSLDTu3OA2n6UK4WlL5tFl/KLXl+2kXv
cMu+BQTZgQhNz6Xa2OJIOo43+U4RcKdGIDpJ00sIpyinaVxfDpzjzIG5Mh3dsXH8
Iku7OKbKl04VTeqdRPva4pGMAZ/OsKR4BbAdj8U1a6F9EBx/NFOPqEFSAY0+sdeK
ueLDjY8wR2XUwnQWeexUak5Tp69i4VSAhwg19QaAU1+XOptEeMhhxmlC8HxtDfoS
NaQpPNrYCsIzU+SXitwvW4z0PPpv7O+oxRYZJy77YVdNbu/iq8ux+YIst7Qou3Cs
4Ib+jBfN01lnbJfjwpiPvpu6MNwg/FCCXVdJHk8H9CXaTE5f+UsSYA1dx/80rXZH
qq63080U9KfFB/TitIEc2bX7F6+uHCWx3kED5CAsURmaVPl3Eu8XmyXXcmtMYrR0
qqM1v+YBpefOkj7pofOXwqoROhWeMXmNIZlgF4RMuI28LYANy9n3u3AjEazAc+yx
k+Hy9sOzoFOZpXk149QySrZhiJR+3hga7TBihulGujmTUI2QZmzz/1kCkEoy0Y3l
FWv0t23DXSr4LnpUYnQ0PGDq/Z3ZcDZthdEFbX4YCRR0IK6ciMOOxICIXqBJawgE
BnCb66NjScFOeZGR037w+mTyp5Sw+K0a9h6dvRy6XUS3mwIAIy+qR/L/O/LPcM4b
j6+pSiA3arc/hr4E58v/I+OIzbiL64jLNgq5BN6rDGinfyr8AbxAxbONytgnucHz
0qJARpsYniifwtr07dVXXlY+6b57SVGZrLKYcimSyfZCgUFAr+133TD/lnZV1JDx
/NkT6e2y9A7Es/iwlIWbJlV/Mgt8Y3+vK8qQCeq3FcuumPmyYwU9+skKJPkVQTEn
AhcHnt2eF+xYIhmJ0BYUhbJqL2W/i3ACq6GEd6zzMiUZ0HqeTqsjm9aJy0GNJf5O
MOqZkB5fDlBQuXtmPM2eNhTW1L8OzhseTtIDSgk7UhE+yFNpGuLNenAEZTgnAIL/
Rhjs/BHI3SF36qa1P7hxOJgZ7r0+TMi0/bYTk1degl7ccZLHbnrrZ4YkgLKmWlF0
X8KzPK6hz2kvzJcOjxIiq3vVy8XvwS0JyEzZ7QKKMXrqsJ5Sb6l0aOdBNfL0fh28
7YkOhwuZZ/rOaGC/SZMRJe8QkPK85Aj8vDvm5Uj9hgJCVRybgj+0JEOoN+IuuMr2
rNa/QTrBxwGaXJEXEVPo28gqLm76oxMmnAGArpLfvgJ+d0X0fNqvbokn3taEA0fY
5MiyU67oymYK//jL9AgFKn+zaqSuuRf62izHY7nPMrVAqJXlaRFWffNsvu8YKFMc
ffFI6HLpec5XDM4tJXnfHtkDBtyFRNUkhVDj9xObvS07QcLov9OOT+0ovg7JPlZM
hzNPO2unRJUEEQyLaMpWL1tkAYArav9dhzK7EgKxC8rM9zDv0uPcK+gfrxFrjvDL
5wCRVDQGD71b/d1hpKksIQNMmHUEbZQn//sb06bl37QtP5hAcpK2IgR2bsuCjcon
IGsYJwCj5H978W0KJjjfq3ivRh83NFCrvjUVyxegyxKSjOHlP869r9uCabVa20JA
JaCp+omxE+/D7TDA16I/W+RLBaefOWOBP4Pnr7iBsHxdRsbqfiTeIxo1xbU8xPbA
elLst7E7v/ryaoJeqkcwapkSrXVvNDM/2sIr7ThCDDGfsSUczOv+mBVEG93jmK34
YrwRRmrQqsgG+mkz6zLCci0u47Qhb/JSNtjdqIy+Cq9SdhTeeqrmIm04j5svRabY
ZPfUlNKQVqdh6Edi9JOJtSv5PYHz4+VuCrjmTsg2qFiJSNt6WYXD8jIUWmQxef6T
BG52JUs9pYgxKTdG08T2agskauE9pXeVw0x5VKtfRFufNfQ/3a4X93rlKhzEZL+k
VWk5Xm1f2Bnh562F2UZUuBExJrFeI4+0BiWYbhnao0REwejg/3eo8hFAK2mOSpUM
c53243wy6lCvzTrGBLbPPBN6ROm4URjyOBLtxaU1tT3VHfxhOOEruioqlPuMTpyy
meIrh7DdgeazIv34dXABDWibf8XhkgLlNF8kElHNc21KU+Jb8SzKE49dvDkGFhbn
3ZoB7/r8RJYUGVOzltJX+6DM1DYGrwxxBnRaoOw9k1fdayqF44hTN6Ic85nLnzi9
x78F8Z/vx4VCW3me9IASWXIvC+CPL4uBv5Co2aGf9vNV9MSpMHardQUsketoTOl1
L376mQsbalwpraPhcVIXq95VgAfic9henYs0AbLpGSnl8AFYVHf8VB6+6JxTOOwK
73aCqJriQE8MKCxDdTQflyQ0JgDmK+vW0k+oH9LfBvTg4RUFLsyJ5AqOmVLeWuEJ
jNIlr7yva7spiHD/85JpDZKSeKIm3XZ+poJX4zi1MJBJB30IsglCGs/gT1Ppqhmc
ZRm0llQzfjNC8m3jM8P67vX3kg6evrFrCgoXQmfHjRDF9DiDxpMtqf8xXYIJdlUh
5xOPX4aodbsuKS4IYQDqNuoweaexxwpE/1A7j6QSxrthCYnf6cypsU5U7hwL7agz
DiRQ80yMOSJkhqllEyf0D4aLe9PV3C8bhWcnngJ+XHLzIqCtKYHptwZdpGQ3OfND
fSqgs3CMFEMNwUUC2pPPMK5ZlfinWKSDGtQK0RlcnOou7l0CmXpsTToY4XVecaL5
+mJ31H7+2g7P5rXmzbLwmyiLqebTykj/mmH3bLYJFm+nJyBDqv4vw1VqSZf1s4XQ
j16HRc4uU6YQmSgjq1pXaxdQBtAuTfsWwhMHk7rK80VXZbSSmvVeIGuhwa11w5Wq
1L794J/Upb/Adqxgjb+j0mGC2H9rfisPXah3Q2WFXHspI/FvQFXUJfN7f9v0EPbi
H8rV0ozQ9ImqXdMgarkbObM9QHQZ64Qht/Xw6tqbkKxjl4S3v2BCwfQAa47Nkxlv
EBqW0HKlNXVedTdNTzyXBMguGMf7JDjxsljbmPUyY6s9fQL/p+nMM2rBZ1JAQk7L
3cnSwAR0TMXWoAWTOrFjsnhO7queA3kw69VVkncCx809hppYHDZwLyCSWdbp/PEm
B/bZemmtwqaGvk6fRwWMdGvg4LVh4XBBUNwzK0BIDSqeTwvhltYfkO6nuaS1sZP3
+a73RhATZnVWR3qif/avf7h75ORE4PBaWv2VuAoWWaTzfZdPh0vvX0vM3nOFad1m
oyd7mNzxhhbNQIyisJIowtWfAQW0K+s18OmeTGMIK05hFKG4tbMT4ov6H42ky96T
mpX+HM0zmi+iaq0rx+wbEhzhgEKpNL/h7HzP1F7Biq9VHb25KS7w8AqvQsBfUbMu
YC2iF8eZxQVb+PnqwD8tw14blz7QErlgCyM5zoNaS3rN9Y/nxc2Z8DW1q2eESLAf
yjEe4jxJM8C3IJQnes8at8vHGm6k5e+DIy7whMnYwtcPVm4Ilxn835etZwssMDWB
LQlf7urd95B8USJ/3pgLIVQIes7HodA7lOS/MNojoUrXlA+8PMws6ASZbxZAIo+x
GMbg7caSCno8opcFK7QyhsTFRbECv2MSpXGLaA4EowsoKjDNDfT35QaoBlpXYCe0
nTTu4ggbb8Ei9TEI8w8D9FGmwXZL9glO2kYWbeYXo+ZaeQWMBPSjepLgGGQnMVy/
z8Dv3bRteUmK4z90qA0htwKpcKv1XqFB7Bmg6OuEqbqm0KM23It7vkaveas7oCJX
wn5D3JaFqSYy0yYvhpzZtJ6ECtyXHFLyN7KITdcuSuYIlfzChgoahcxeT2X32m4N
4PMxAhuvzcDRZ5XOYY+QMDn8lYYxW2LEC0L6Yc6IQPaE3oymCxB0NVIFWUynY4xL
uEq1Fv2GI+AgLv4X1EU701YbHa623M4pnYm9KStkPmNtca3eyHJqm+RETZV4pKd5
Hr5rHHqk/GEU3Ta5/Q7f1/o9zR/oLGwaY7GdGvkTRFUblequ/9FFdEE58gCu66aX
/zpXMtD2rGt/uf5TcJYvhpz5uT6Gt78etaWJ2t74DhIryyF4CQ5nu5cO/IMSivju
ambsY8KAI8MQEfrbDLir5Xo6xPE2rbcPjn1cFElFVCenyQ64eKZ/vKZuPXRBZqAt
f2ze8oo+g3nkttqwiQjhGEugAX/KPi1AM6D9RSwTMXXqX/fWhrNskvQEG+K2jwq8
TsJhLcHwr7NPwt6KoaF2QIz1CUpvS16g2oQ/4l8h5AYLpps9c1wio+fq983z6dYU
rh0WdrCD02+S1NxC0LbNuqUxYmTyIN6DK0pwIwzy+vtQTEi+bgNjQw8uQeBL5LJ/
FOcHsvZ31rZOG8ZGgjaljzU4/ysnRj4PKzEzwU0rEowFNgVH/agLDgGSolPSRlYW
toHGrijBwbY8r33yDrwDAgBB+mtHD8yd87/ObnrxtUy5VSlaTV8V9VcCsuhupqUW
/U+Vrc+bYD/u849KEiIMSNlafPspcKlWEasU4G9/oBCTiMZi5HAC2LQ1WAwdyUzi
9Dx9RAZ7esX9NGEdvnYg05InQmbra5gVvUKBzNdCWB9lQz8/chxrLBko00BnMxtt
cFlPweBBLBfRwxiGqI1+c65CTAmObNySgnTSzC8eFPgb01sXKCmzZXp5zhrSSnI9
pF7swCKVx61/t1dNcrMlNJ+obt9kEoiQeydVugdjxJxU8tXZPJJCTTaEamRuJNbQ
Im3QcbMQHSkt7+uoyA1/ob9Pbh0ETVU7KbH+HS+raegvwf8lOuosp8TKhnKQEKLp
aOwpVeeDIXuzo0Otetk8nMAjIfx5YL2biflSn5ooRLHMIg8DDeFq3o9NYZHnldhV
dyAAlbn8UgNa1YwSZSOl4dXUzuUaYSgxGjt7KRpAns/0ZlnUFGC1Dg+uC2yJmiT2
hahpWxbAvh0LcSBHwtr1PkyQwneAKhCZYXo1BGLjbzvJBTE6AJ7a3OHNNTD8v0hs
ZJS2u/B/cP1qZc1XWVU1IrVc4gjRLkz1uhnB3v6O6saNure2cQ7zdJHO+y2Z+7e9
pgLHSCn1Ui+0rQh7l6f+nM0HgZNdb3IMzXYAqLMAnGfzzwYc4h1wWYg5luwyqWNz
5BkPtTGokVzNLD54wjlovBFZYTNVAxvvVchqE/7S5jM3vjHD0HdoTTaSF/wio5Dn
Ac+hcAjxddl2vdeY4t2KNbrijv9HuHd7AtsoCEeYCRJnsx72d2v6P7grYVXmu6h2
FixQ3xTZm1BwITeaOs+2rWIDIWarpO+dUZeHb6/N6m8AjXFRt5KBZb8VSH1Y6MKl
035+wU5IxgHW3qPqiqYjhBimh/uYJH8D0+aMODVzqlB92UIPUfD0otkaz+qWay6T
VHIgCx/aYUkPjmqaLk0sKEtPf+NDMcAZe1oKCkL2wragaj/pCimcJb5Qx8ywincE
MLE//QyErc/R8jCf4rL7SoaoKEqj36cRuze2Jvtnwl+q8qg54S/V9hj9rEnaOKND
GrxjzwQ9ruj3Z/TKux3lY19dXXx7TDNYEgt/SHdPipyCSmkE7bs8aNYcM1PaaaPC
t/qaZs362g/xg6+vpcxhIAH05hs2xeZvPryJ+CmOAsa4yl1g5Oefe6860cfbzdkY
5JujLvPbbCPifrQiIVRFylJo7xoFqXm0Q6wBwVg36hDEES7+RmP8iW2zxn30VldR
FBWKPfz2x2LWxZcWH/X22ILqG4CnSk5jRPoTLL5y/nfxSxoKtYJVi9BWvGD8L/ah
+VnCxBVZdeWuk7D1nPQyCTorGrKw3igyC4Ns0WaapZj14jQVysnk6gVMZRyUxx/W
ms9qiqgnZ+/bFlbjfeanFNQo2dtnI/grbbtbb/E6RHsoXBJl9m3pHW4JmJ4/Ol2m
CL7J4wOw+ulWzyvjCFnCjVSLpM10gpiQKQhjRn0AhagsiGb3CQ2khrm4Zuogj8sn
2LmYNsbq2KBiZBAWITTTsHc+BMUQ+JZ+OtgZNxFSIz1Q9sPzuThlKyXLVaf3gWQe
pYBY6W2cyN8Sn03vd7d5fsJbatqkn/NgGjvCN6XDZT22KH2iBRcw9T3aLmeXI/bK
xgDp7Qx33HL7J90+jobrv5nDPKm5mqzPLB7sMYZbN5YXYIfx5fHTk2FzSON3JA/C
miQfcAmIjdpoi4ylEc0XX9AKOJg254wpjwyXeuc+m+A19yVpSzO3+a2qwUwlSdIE
JwAmA7/u+HcuOCg6csaywv5sfZm1vwiZrFDs3QGe0haSA8daGczSI7MF/f6DHqyi
Xjwvp23BF/aNNGtO/QuOTnSUPusbi9hSDMtfCTo+JOx1rZrBur2Pzi0K4tPxuwBu
HVNhDfjzBgFLNbgXYzUdPoaao/ThVQTcSbdQGkeU66AV3W13LwNlHAKO682wrMoF
Otmns/LwFleGp8Rt3Ntzv+4H/3fux3nHZDOMPfIDLfanHOl61RVe2XznD+TseJ9b
575iScJPJvhmaGPEUIjsabTOzU/frOFeamKLx2n4prmnQGT07XxfwZYFY0aSywoG
nnJlnI45MMFU+s1FZz/+R0bt9qH6631RJkv6DMHjXwKPBBFmxTawjOq3Bctzlstp
FgPeouNcC5XVoEGpNqYq6bvftPqRPUxIsdgtpAdakC9nps4ra4VgGjBvabT4uNQW
Apzu4KHBszAZoH1JIs0I8dfUL0G2D9YIYmMZKzj0CtbR2MnZGbuVfeBff80VMZtD
u47KeThG/wuivzfX6N4LHvFLFxbEDU8OdFbtg/XcalykwqzKaO0j1mPuP8XVI1DC
gEwq11T4du+IiD2jqhBh8Dtpw6tAp8q1pUxlYv5Zff+9gVP6z2DqcX7UPLmkrFBW
QVKrJRMVPSvSVzB2Bhd/rO6UOKoLtM4Bg1Vpd0OCEGSZj+qf6xDMSrKpc31Zsd68
W+ktJzfyh4HAj9bvUTOd/i5ANhZDiQZ3+d1HTLDvPLK6HyaJP+Qw0T64wIBEKBFN
NQ+UqcCpIUh8uSVx5fpzDuNILTsuKaIo3zpdp83H+xiAUqj+Ycktoct6rTTrrhr8
uAviQ63hADcihBnJoXf5RNiLSjALA7igUN7MC231cu5+pto3DT+gWXq3IlcKAWOU
sP3T5KbsI0lMnO5r/SXdn2d0cF36IO726jwZoZqfE2PtwgN83uaRDu0B4LMa7OCq
MRPt37EEki5ChC+8mqKew1vWk8iiBnqHfohZjeBPhuaNYIMtH3Ajqkhkwr2xyFL2
7QNs4pFissWNBRHdYOT50KA9Pfio8ANLmjSKCB9XZIkFCG0K8d/58ffTxPK6tTTt
IVlMauZ4BOpTdu1q38iiEbRs9oWbhcFp0X0yF16vbB2JnnRgMAnTsngennxcgTVd
qvz2Yoaw/F3sbO3/4TvXLZXKJUeVK57/L/kQnKobcPONnBev2vZFvOcxqmkRwb3I
Trd30Zc4JYJWF8DucNDQpQo9UeBnOPANcz1aLRyDE9f0YDNKoxvQ78LsQqti/JkZ
iW8ed49QGj6HKxnOPsr13AxV9d4COtTbXCxX1WYU8PFFZX72dUQeyxfV8+IwYAXq
7/iYHy2TtlqGfqrLsC3OBdmbs3ehbHUUQKFdENxQzNtZ8xG8A3tE2/KFF0yiikcG
YAo8TfvshgMyMx0n92IDCDdyuEOqCf9eSxqDfOqNvoVQS2txSJUiftTh0TRnLV9T
usXF97f7BtbQnvmRIKJgb6eHcEX2A/6nhhvs16dCt5PRdSNlb8RfIiHyTzayid7z
FLD+AJlzoiVTQEacWEQ6lLTjKTRwe8xSi9dfTt2roGH9BJqCS/y9K/TWOdx63gmr
9YHZvNxNBn0ok87Y3Fp6hX3zIgMY5NZfTqyE6IMPQQYmNlQBWXMyAwcThUcFtuz4
RSMwiU4GXVwaMsDmesRarjWgDmlqf8HrvqqNAfyz9mkMwtfMvjYP+asAtPxgSyt+
6u/Jj9QqIy1XbQWzDVg9M0qygItd21ijyJw3y9VBJYG4e8qbE5tFPuqbbrp99FcA
ai1TcOUTZK7A7vW6VNhDsiz9LvUs/hnk368T14wuRPghn6M/XWDXLgKDC+oIgRkj
7t85a1XbWnU0dj1kg8EtE+J9o9aon8fbwXLExZOKqcFxYIhdb96amN4wcLT3nVla
XuGdOsLhz0oBLTs0CQJuILc9KUE0hn2vJf6r+YmS8CsuMdSz6N8KtVR5EiIcw0yW
Etji9wfXlOfzWuDd8x1C90FGP0uTLbegZFxqfSTV3Gs6Dekn6r3kTQWFdPeLfvR1
d2mt8KbavwBXHo1iIaCXCT3kL8R9lVlWVLF1V9dg3KOJKLXPqTUhusN0z/e8/SOF
cXivOiLiDGhH0j1g/LqayrSBDjU1a+PtHeGC6kTTkdH4r67YWrmof0KXcpxcl6t+
LwEamL1YMM5C0L5LpV57OcTEwa3kiJu6wUIpuxo4LWqlaF7v4knKjK58o+NHNYsR
8Ml0m3fYKqTvuxFeQZ+C4CwMivpa8YeETXm82Sv7gY8rXVyLOFoLw78XjLd8C5Bq
kC6bKIzvvXa0bIp3p6GP2kMhgThMHcluP3Hu67De7gd9lYbDoDORglGXJU2f5GXD
eyF5YqUjxJu+fZ3mdYmbPKOeOpfsJIK/mze0s20B3fYDn6muDGvma8hTcVhAx4Bu
Gzeo77p4ThnJs/4EU/JTIjBncG+xSeqRXo1nrj4usF4z85DCSq8pdIraonU0bm4U
GQhBvCHtVrllM29deh7/18Ad+6UaABzBue0OscKxafnCAbM/CdfinRvM4WDSfHhY
bN7y84ik4N1nrpM+WKu3afUlliSdypxO6u/ZuAMLqQtmaZHfTjH0hxsC6ohlTs6n
RBa5W0c2lGXQX8x6QaSiwq2FtOQOEmR1Yw7HpTHjOXHToetp/VWZIbwOeM0C4fwm
JFN41cLg7msYAcZdgrYvHXPyv3Ij1S44PAj9bJAjNDJ/qMskL9FAjJLZQ3UBQLS3
32qQOTqcGxbPRCUe6lnurix5fM38GeIz7oW98Fa53DKpiUhbDc+ccHYeP/GAuhV1
GXECzC4g4ER1P+QpAG+nEf9zHF8Pr27irZxP6YfQEw+uHBd63A9tjSYpRqo4/bL0
FDuep6KbaJSVMWLy9SRtdr+Ikh9zD4gGf1o3DJxT8MEs0uQVW2KN4xcuzvKV12A0
VGPLl0Vw0oxeEZtBAD8sjJe7i8o0KNIIy72M+p5AivlQui1yt3ezPcxVOSfa4MNS
a2XDBjACfKeqQzBRjk6kmK9gfl6cZf8pq/2yFNV4v9AdaqdUM1y/SXswsxQI0QoV
XIhQ1hrbvfDXd4Ew6dGSJ9l0MPiLeebPBg+UWkLfWHev7yRXThw1N5454Es0On8f
ab0Lrib6WIpkevOHSwMbW9H9UoPsmAKSWs69LclfAMs8l7hEc97yPKFHz1wiqXfQ
ki7tfOIjhvzKZRFt/b1qpVrmJ120HdEYsikh+mvUSA36JzpHKi7OaSNJIXfRXfja
/aM8VEavrz2u9hm1HZvVcyIrUnhCdvXPT/k9EWtfAMTB/WVEa28k+072D4EBXQdW
jvkO7YG3yt+JMB9Qu19yGlpejydj2QSyxn2D7rWC6L4y9e5L+BMcYRHZVBMiXug2
CJYyzXflkRaMlT5jHjPkf229Pr8/crCCMHGNgx1jKkr9Jwe9AKG4ItX7MsR2oqRp
aYP/6UY2t1SVdiQGpDzTDE2aVquX0Paaxd/74qgKjkimmXxhO2FH+NPeAO7vgRXv
LYOibpuK5eJW2t3BOtpT1RYkZDtGD8bvpsPXzGFCtUfjHqe6DlXniUD/nMr2p9Px
+ugsxgr9ZPtSHQOWY1ZO74H6SnPjGWFmyIvwW77AFKjWH6OiXqaMe86ZLjMdNYiA
WLFVlDwt7VWy4Fp3A5CEOjWiC4kN5yrNmdX1zmdHC86HHQ7Tq9EB0PvpVc+44odv
4VXlYoOLkiRvkyfSIQVJVY8GaXAR/9Un7OuWtZYSo749Kul6yhDYhpWLPLNrJhXt
Sj7cuJ8igrHS1L1mx4IRrGYqHaegHTQmxjC/zPb0xSQVnXpSCt493HjWCC3Rvx2P
I4w91sZy6nmZZQbTKHx6FTRU5wQOMI4vxw/+K+IxRsuJBse3xgAZ2X7rd+pNu6/l
ZK6JZLUI5bHSRQyNlHu1e0/NUFS2F4jkGOyTEV1fchyl69DXoJw/wxNRd/hmucxS
XuxUV9AmYnCYQHa+x6CMwX2vi+X7hf1CAvLRPq5QjnTX5DVc+FCOfmIcZLzCiR4l
x2E9Q7LOxOFdC924UJ6pATdyvXoUMSXCz2ZuALpulSVFUBDMLMhmci0mjXUOB+5o
vZrE7chAiEaaUp8cmFnEzDoC5dcAgY3JkPhAXGPpkwPAob2Goxcep+FwY6Y+eYPl
gllOCB+bSQO8fYdQgGxMHgRu8X5NmQyRT0J2YhOd5Kz0gPJ7RnWQziUXSE0xRCeP
sbqF5vap3UqPo1hNgRwTac0Ms+0iZvNCV0jN+/W5FLv9j2DXsv86oRSkBdiuMaaK
tRIzLxFVylIGQafkyUSNtr219TntnpamzGW4jon3NSGO3eae16aDb+Tk8Pe2IJar
M4KOpc0WcMWkYthasJe2bLQ7o4h2sKIDvpDfe/p7uF4GWwicNhcFLGlqXrF3xg5x
QR/3Ti2YIjnyGLo/Ye1/QvFWn18WiN2mo4E7+XoyhINON59Wkq82KuakFji/Vahq
EjKqZqdXIboad9m09F/gYKpSZ043tUX3yzi5kVFSeVBXyWN6Jd0DozVHcU3+wl33
7J2/6pnRckDlFMY/xVBzvo0ECO6uNbiW+LvWnugds8NaTFK0kwvuVtFlcyZ3J+3+
SMtg27MG0Amw/zC8fjWXot7NfHE1V87SwSBv34mv0IeE78gWdYzkaalpqtIqOrQe
x3IS3X0oCMoQVYQ3Yx9Om+ULhn1EV+S40lATDLX81MsfIdQt9KlU875/+hVWqa9z
zilKmtrO9EKNvVY/Aq/KHl39Lx4YRvFHvwKAeLv5N6DOS+KYksQ/M2YkZpGs7UeG
9CbT7vdFaA0Uc0+oQ5VuqmY/Oox3Hl3LS05bIvDVHeZ9xPCyM/s5kI8roh93uKoB
eRUGOBLzMKBJppSJAilg9LGBvENU9yGpju1cF6WfYh7wSzVGuahSTgSuQIX4W15/
IXXBi0tsSNB6E6ZupGJjrDUbEhOgB35C3Ba1sw8RmGOsRntGb3wXRfp9Wp53AyXt
APs10/fqBqABE+z0qD/XWsI84pGV6EuivTRNh9KchP7zLrSvaleBnT4Xdc30+UnK
heq8VTVRdNO0faKevsKrqrFPbigPXBkr2ttB+GQEJ3vWnjllxDAxxYBu8X9R6uy5
MzjwXXdbu/CWfejAdgCns67Ix1tFBEyBuaVcbKJgphfCWbJ8T2Xcf5v5MlVZOnzW
i5mu3jjpOfNCMV9v4uA2I31n9GzDNLnzTVHyF0e/AlHVFsLwA6/4NkIjumpBI5p/
mUyVABAgS97xcUyv8ix19n/fzONYHdblJlmNYAX6Jkq1PkS/gMTFu9pslhkaiy30
KjvVlzJNk0wLg8G/mI0O6dQGUQX4VbjG3woHzH2rHLfxyUw2adkXUkLqVeYkAwc8
GltpOUSOA/6j+UAHUNs7Q3upTb16KYF41CChdcY2Wxo5yL5G0sXDUKujy6BGMI8l
WNbGpmyvL3bo1CvFt66cqfnV6zC/1ToUege9UnhCzuHhNsbxMW0aRKmFugVBl6va
T/Az6FB0WTW3CY8BmekECy/P1YbDFROCj4FBdSgo/beGeRABPFLYDSr49w9iHRAR
vIQUtjZa6sme1axuN1sBjA==
`protect END_PROTECTED
