`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XEDvqJNNsJnVYd4f4v97AVQevbvpAEm9ngR97IWECqkxdbT2Q+j3nOe8fvSSyKCU
gORsbXl0JWSGRhMtI8Sb7Vwu5dS/F/rREuUQ7p4jBUrihRN5uOWol01b7RJ97G8y
O6Q1NTqFfAWiFihJGOli6t+5kIlxbBu26hg/qT8FhhS5v/BvhuF9wCKQxi+a5cYe
AhxgLKuY5RPYRywfnYHPVxbMrvhtBKTKGmawSOo3LCycFGEFWDZeSlAr0q+Bi9q6
vIx0usjhA7fgvm2RpiFKNJbOwB/WzIAKj5kBkP7iBqTUKUKlkBEYA/fmbduh4GDj
UtATo5BClZm4IPhVlIs5FjmoxsaF+1Jkap9SDRvDWuTBgqb05ORBm7RMRoxjlDg1
PNJRbUDPQ9jo5/q/gV+3I5TeRhKlKRTi/5wXzjli1PueinRgsyzP1ycitmZN7B1U
crmxZia9289ipnQWpKKuL/jMm2/La7rOCFxSRnpJFvSidVrgoxn/i3xUMoTp9I/I
bWq/y2jedavjM1IqVlzdaGufwawk1o6zUBypg9Z1Hwj7U3lAFwz6kXJBG4Lpjoea
PcUg4y2aZuV6pMJqdk89yJrfC0NEDOBBq9M2ufPSa8MU5BZh6HO1e7seVth7caXi
OttF4fJSdkgbLis7XFYbVngwzNNpBkAydWIPY4snD68zWkdjgqVXbBfCtDSMiBFt
WzbxDK9dVopI7PsI6kgwaY4ZOss2BxXOX8GTRpnO/iXv/SK/rAE63MsmIzyfYeun
qpIjGaxHq70fH5/UvadlwQWD5byUhbex5clC8ucRz/9wCJ7xq+AtohyIWmvLi4u4
IKKn9pPXJiP4M/xJ7hRIJ5aGVjv4rUzY9YzIkCLyPpTjbFb6FsybKZs+iW615gX/
L+8fUQtw3idztpFPgoJPvTgSjRViCnbnG4PWRbh5WHG5FEriIbimhNf7CDcw7Yb2
rLY2afB+DWOi0/To7LMwZG5WMspOSkawhbP/cP9UajMQ4Ao8lDNzYL6psROZfqO0
EK8f1XosjbVuGbttTO5VcDlPvLveAObN653T3ieOxIexatw5etbDuPhMlRpb0r1B
9BxTb9bkKcZ/6b9wqH1Cfi69MYhdLmU9bW5L0YyTr9lz0sMFgBVtXFLh+YpipFYd
DL2KX0iMP88+DKBOigzzrOryk8T5G9GolRAb8qvs/jGY4gfqFzzG4mt+RrbTDDv+
7aQjsliTdj5TS/J1ikIc/VviuApv7TXp/g55uvZqcNFE2QfP6h+2U5/KoA5+WIR/
HeB8ZGvuGR8FnAUeS6xgDfeMqXE+Z2apnoiM6h8+dZsaZ4IOsv3e0s/vSg2MsZOo
mo4Ag/+448CB7hS/k/cAyUEYVSC9bDFlUW95AJmZgUE0R5Qnr3ZIg3rAJalzRwHk
uNukAsWYTTjIGaj0G9zmIfa2wn0xbUy7ZG1YxAnLXdfYC0HIJ864kmII9V+JfZmW
Hbd/s2q107YxjouroMDPA4CRKsirKyBKIEGa3YcMGp8zAGlN0rDMYUbwxZxiofjm
XPKCYomg3YEO+kn7W30Mc8/ozqkTaxrQDvSoQnp19i06pJ2Z8H0xfkPSE9Lx5TPv
HvLQNmIXVdWEDTPHnCdUmNjatTRHvqL2P0ll9OD0ges1o45WS6W2OrRULAhIlBO9
zG5NV3jSSff2H6i6q9dmdEuCcv25jKp/93Aqr0EEb929ZhocUy5+oXVF3trgLrIj
f9FCSHu/CB2MRltgHXCRf7SOm8AA+anBWQPQPIvBW1dP8WtNEjwqatm76lJKs2ec
TwXtmjR1NLwJZbEEhnpUh+p3Z7GqJU3gGg1CpnjKB5QGMIamXJHLI/8VaDGrB40O
FjOwJw7koUKLqR73AY1wSgKev3qjZFGDmo5zaiFjtuJvcXSjmRvPJqGxrkk6hs+z
7x3TrIV/cNNzhXOtzQQ8Ut7RazWbZCMpq8uM8Ne6Z6r5Hixi5fchaLYnqIVseY7Q
y7u1sTX0j65X/OBplhWVGw6XoBEv/ycqXeWsTRfMRecu+w0Lg+v88L2bpgYpBF7Y
CIDRHNpN7uVbq6fPZsMyluykI3vG3ByV47eEr7IJzbcbxcEL7kX89A/wotIHSCJn
b7NCRljpXtmEkRhhPplTqUEtwh/qyUi2DNPJfgK+bTzS87Eszfq4u8C+WP7KPiQB
29pEAViCxO4eT3/0bfaAw5hp6568aNWyFkSXPjRDgu8sLV3AbTSTGQy6Tzh/SgDS
xYMdoIRu/nxH5Vd0euTPODp9e6lIY777AaWmrSsRxrLpvJeE5gFHCgOhSLWDUaa8
v1QAkPbgzQYBAi0Roy9Oay0UnVCZhlCf89i0TrMmSwVdUF7slMZ3K6ssa9/YYgdd
vUXUixGZQa75MBaYsT7zNt45IIbLIrL3KAxqsYq4R8N8KcMbD9TjtaU8XBMRt0t+
pUnQILuVnUD4Q7oxIitIZ3ZBjlnqH+Zdg+ESVyhsxiTVi0S2uinqRZCbYFSdcTwL
ZoRt515qjbHHTNz3/BPQwFUmREdnWP0sbUsyiI7XMYETkfay9nlx2UDwk5LAezZx
DMNxntHBUZN04qJs8SEJ75SZw/EoeVw9AHBBa5j1m3wXpytzbrGQhy9GLXPaU7w8
lYl+60kw5plRYHmsCT4UsBtZfIMv38cF71DvFCjDMn+n9aYIVcxW8W89JGkABV0g
qdqZ6dyRDRJ/aHRPtG7qDrTwYoFW13yLXYOmJiqVcf/zXHLc1bJM4+GGLi9R60uv
cGbyA4sCGLsWetJVrln9mQAX3FYLkGvbICyyGnvLYmpkNzMEHQcjY+mlbbIUdT4c
IJJy0Al0a8mkpzpzUQglMCx1naQocMe1qgZNG7MNjhhzJBLaFqYtmOonlGLta/4/
HoYNDTUYK2WzvvZ9BmdzNLOks2W/L8kdTOF5NMbAd+U48y45H90s4ecRA0HaGBqo
9YTN9IY4vvZpIvfCydVxwnoJMz1+x4XZp2P6Rqk6krEMv3leLu4J2vYBGIloMobg
8MlT6J+TuZnTJwIP6vIrQrUpbQxosniB6flFe6OfCshvrOdp0fwVOPVI1RfCGmTr
bMf9ieleuEYa6G1rCZRa9aIubw0obSLGRYBFSPath5JJ6pnXqYE/k6GKyvh8AOuB
XnWPnhQC2mTyj+uLPH7MSRNDUEtoDNGYv7lB4FUU0so7QOuF+gEFGXHURKaKcWMz
Zy/0D7AGwnLKnli9qA0Y12LOSL7aBJwjXP0teiJQhKDd5KhCLb+gAAVcqDCaIt7T
t/QNiXq8QIwZ4NkOeAeM1BlowKhDY9xMKkTtEFnJ/FHlL61Di/DDalBopQv6OKAF
FncFZ7q3D3Mq2EeZ4hJY75TqYbCVr10Ezvfkj14M76rkTUJpGIUAX+vy/9OxodGi
2r3e6KbV6dl8G1igMr8bdL5mTqYNDxsM4gHfE9am9x8a6gvvxMXdGeEIJSsRLzdQ
FSK5nTuDIj1mvvX1PhBky2AOZ4M/dC5ndvys0NdgDJ9EXyaNWO4kT63KuVHWGQqz
ftW2hsslr2dzA524iUSl+QJDqUaFoxBEijkW2M5b+5XT2EMVdGIplANNmh9HTOE7
7USF+aWKq+00B6lujErPeIxJoTTAhKp5uRw/NQrpdv/CGNDhdPcuzuuFBZjHHReQ
NeuKI6/5hH3kiO6aBqANrHGMlEosi8WlF9DP4fYWsKJH5xHKwmm/kjHNeOlSV9Z3
IrTYS3ATksQy565jUE8D7cfe72LEIQkdCJcI+10Vn1rmugibcspzr3uaN9xrUjJq
+seTiPu9GdkN1d7yVIlOTm3qnyQAaaIpWZHFL395yDgtKrE2rCKnmYxyyTcHxDbT
HxrSfTIAAc9pd5hQ74bcCC54g8m84c7+76WRc/fc2Y3jtqKOhGaH2JJNisa4EQ9v
VPrrLe7QwlNrsNOwaycuO/Lz/V41THjtiYRksNZI8VCeKbj2Sky5o6ZYGN6aUz/f
dIOfzuwDmGzRMT2r3QFAxR4zXWvNWwJJXtNCKXUf6lyKuYsd0dc/zaGuyRyg08kl
sZVDBqj0MV/VLJ7AIiy8w8VPsOpn23SngQpmIVb7rvQoSyGqquoSchshWsRI7tHz
+QG2LZsc2h2LfDPmbyip4M49GdPsHdXYqZXFRiGEVsRvrqwVQ1PVwM9DoMXpJ7wi
ROoNKIuS+SPkAY2rot6nt4uNdeofs9qki5XH2zE44DOIObJShFKQwvM4rXY77yND
0p13CTOAW44IkvEjSs5m3GrP1St6tTiFIK2b8qKhkiSWqsuTa0zlVmBMleawXHwa
/Wrp3ll5UtYK7M2vBFrC7s3QPUF1ikLMRSIZQscVWk/RWeBSPQx0ZiqO3U01YrtV
fywjBWSQ4kyEgwDxRh7L8JW19Ul7Z+IVGosu0tJ1/TWlxkoXLjq6W5Fcee5qbFJn
frdZS9sDDvl3cjjmIYN7a7pzJlnvCCJ5RiVi/oXYUXqCUXaY+hMjxEg16op1OBTq
uSqyNSj2ahF/eHZhA8NGeq1tJSw6k9LWPo/aHmx5iKmevoIj0nYyTSnthwg21saw
XvmkkFODHc0LPhn2SLVSBqXygmCx34VwafeNIzlp8rxzc9xtse60UCCs5eU3kq82
3eHTaCXvxN6wW5ebJNth1JDwv48095O37dR45/mXblQr+2kxmoXTwo9wSsHYqh6W
5fiB418kuxNlh2XTNpJDfOqYk42JULAz7kKrZyorLGO0bMGj4GjahCXTLbh7pFUi
WlgtK0vWdrZMqUid5oQZspVjHaD3Rm6FMEsrjDj6q9TI+EkNjVly1SDw/PR8OoRM
XVLTLhIitLmVS9Dk6jqP2MyO+f7oi7EgneWL2i+uWh/Rny7ZQM4WohXQcpxyFkiB
nKYlpz+C1Lp7PR9To5fdKhf8F+lNJoyGeBn0K+VXNz2UdRQ1AX8zWIKVzylc/ww8
IAotG/xiNZDR7K2baUIvmXRII2CPMGJVsuEb3LCIKr20TIyVWWssF1XdwLXWt4DR
jXh8ubPvC3VU3ZlfGb1Fo59b3v+tCIySPK3tSavTKWZliUrcO16U+Uty2BMRUI6v
6wIeCQFn8gpOs1jJSQKXdsHLMAxzBsQMDo1h7KQLz3ngCvQNFU5nMOaSw9qXAB4R
Q3PR2g/aR+QR0eedP4Ly4ucR1n/B8HRf1q9DhC1B0AKX9qZCaDofKaWo0zkQWzf6
20qcF8ftjvS6JhXVyvChGLh4jsqAIoqerTGespeRY/91YMHq7VMc2QsDFkvvU0sO
pA7Ywt7Q42X1y1NM8CFZtDNEsrcOjgLQPi8nZMTRh0+4zBAwJI5pO8vABor1qnVP
LIBJRR9q6euMdimnMBsRIhepBnbDsxZmpRA//I67EfQxSsUPdK0bqSNE4vAyDzwL
avRreyK1yt97kvfryL+IVkW9oEa71LSip1ISR9t240lO/5ayUMy2LBhEJuSUug1N
Fo+PGA5ZUmpMWGvf7IPMlnL83Hkw2fJpiy43pD8UVOif0/299DKneTEIcMWzJNE/
4dsbPGt5/Kuf2RunetsWJpjh/G/tnDRGHcOvskfBm4fc1H+7nhBa2WBFWNKYJz7p
0KO7r1ORhYLHK3CdvVx8aeQ+4YbfgTzq4mDZGapUxDo79E+alTSkKWyWUwy9v2/M
EtPqm8EK+nNuNp1DymTM9L2EWKMN8iuxuH0QdCQGPtC5N3hRvJCL36BLPKctESPi
YOtka3cGXJbYSynHOht+OSYTnlRH7FxXG4xJj5V+5U2XORlPynsKbo1QwL4a9zg3
jSCAbNvrNoC5M0hPSb+wLCDJtML6ajZo9xrtKbzpVTLz3xRWdTe87S41ecjhWZx9
mtyrifzgmXsqDJ2ITEKZtVcYh9ZuaLs3vzQt5qL9effkYUadk9FvDpQcCU62VhxC
bCjFNsMT3WPUw0eIZpEKbEphjUIpDYPgqVko62hsOgYdaHLHOBeDLuqomZnvAPmV
0x5KfBQ7U6SBq/cD/j15dRpu9grA/ikUfcp3ziPvlCGjMshW1eSFJrZrg3W4mpxp
8giPagJpsiPIpPLnWcXlt4bXMN+P2eQtpFqicncp6R4okZy9WL/A2lbjOwOhNZDx
/ZbSMOw+yv2s+O+jJsJaxs9qIJaO7Rl3FJxkcIyfqwK7t1ZxbFNUIlB4LTLEmlBu
C3+MG56+LnDSFZLLWM4rrOs/HVK2H2rnwZ3BxK9OKf+5Kg1ahW7HWItQT1jS+ZxR
WlTe08Oaqupka6DBTma/aQjhf9kmTn/Zcm4D+eAO+rDqYbVHLi7M2IWmnUz5Nzhr
V/NLDUX/JELghdAB/2d9lRzn8n9tQwOC9ykh5Sn2f5LJ/NDZvGihl3McMckgUzdW
6VwKma8s9rBPvhO75n2tlv/UGovctb+StJRuRNAPvhauindQSLeCk/EVaZSXlfls
4EMb88orHAPc72GXdyPbpiev+JAPD5xx9hjorVvvgdq4eWR5GNSMgeybrfCk2yHA
Ild5gCDlQusS/BdYYQ+ACm/gg6FI9lVA18F725XruDHs0pbICz05dQQfw8L0MgpS
iB3U3pF5yFqPQPuejR5dxNYGEAYfg6tm5vEq6vzQvzRP0xseZGytkH9CW4On6JC4
IcEe5QwfjgZv4ok8nVgNY5IrhRDfMCzll7RjPFDhBl8mZEVga2NoW9fNhDmUNmIf
TC9z/mF0xiACAc4GDt8rnsB/22IIQVE3xErC97LeflAX87SdRu8BoqXBjgdzBa+F
AO6aBam6/GB/9uoYF/mbzqLc9ESKP50laPPY/qwWo8LAunhlL43SfiXJvyMO/eaL
jbbo/xD+9DsRW+8TZmAZoNoN5GRaZ3grafHi/w0f3resKiS9FVmzl5/sakvbgbVn
Soocpgp2u29SyMeuSF8+eMH8k8zPOMdaPCgUI3fAs2jdHyhVtJXDM0yDwxsGW+Ne
2GrqAGQIJqJfkT8MxlDTw3yWni3ee/crOy3AB0OXzMtRp5RVzaFIgJ/7hgRsme/u
IbqIB9hyJXvfY8O2pSmOw3Ay7SY+RIdc1d1rHq4b/l4KHNZoaUwfhGwHBoNqdr1q
AfgeXM7y3GUcjcYGja9AEv8e/mhqF8H/gd5ID2qwBHRhn3OhW0hbhUQbVqfEHpL4
R/+OZXKDXs9DsxYqUptC4cdn/js2TpiFH5Uta2qq3Qyjb0LCoOWl5FRzqD2YzUlW
+fN0Gdcw6wQszf6koabD88dEGos6vUtsuXnRYCwbVmUAfpnUtcd/MbuIkJHtK19/
wfd6kJn5LnqNDLvWwj8eh8WM7QD6wLOco5i5QgjPNSWPB525xMS4GJDnJkA5Gc7x
yVuwJkKpok5o6Dg9ifa6K7QcHRiq7SyTxhgimPCmZ7/VsfgIC94vouQnv67Q0Wka
cExfcaqPPvV8/ktnSWdyIqY6VXSh48Ana80Xi17WTfi1w8Su1FIKnin+0OjxBuQL
OD2fjnMG4dRJXDwWKR7mHPEuz6oCkCTbZ/ua5oI4h8olCCz1valEFRP9w85pfvBx
0pHqhRvw0UCDGuQEOGR0pzwVApLbOr46Op1thCBFkW9um6noUXN/DYSZVG/29537
5oVe4dScMzagRDBzr7/K3eV8ZmdLTUnKUzTaWh35s+YUyeVd/QcJ3Gib1LIiU6mZ
fwHBbibi7u5A+JuqxC+N4bZ6PVKEteNwVDFgFOak/RTi4MHs6yWLLFAGSc1A/A40
KP998OON7MTvYbyX+tqTszU20c5eFYJEvs+8exmZV4RYgUd4EA7tGRjhsrqKRpx9
tOS6W2iw1vGzy0zex9ahmF5A8UhKYU8NS7722p1Ozy5xGjITOyA7L7PA/u0j4XXK
wOhqZK0M6sa0oH6gCy0A63Md0Ab7o3mFDre0WciPcG3M6oxtccMd9p8unUZKw7P7
kMQ0ai2Rs2+A/30m/0Tf4C3WmlOSZgqaSt4JGVMY+c/Ib8EaCyT0UVwM1XRS4pSQ
a/rtK+4hCRsoW9CiMpqi419o3LF21OXn9atvaKeQywyECUVo0/bqTMubTmTg99a/
deHA6OCUCrxkmZObtSbh65jqImgvGB2pkCMj3wQzNtTsg3hYTN+nv0r2ca/ZwXeV
e2halzJ5oKdkFuOnSBkfNQa7Qa+oRjExcvr8qXLL1SPjm63I8r1FKM2cvzGmjF3S
pW4KscTF3yv0eZFonv0rSPET9rYqakayefY/eEolg4aDbaPsP1B38dUBGk13KwKu
EyTBr8K31XHOX1u/FX+Qqj40RcxFutY6pNyHjDBv13jDvfRNIHLFgrOa3C4rPfmy
zGThNi5rUY6I7p+Zeoj6EMeMsyFnJ3jelPbr45nfrebY0I8JjAAHweI1mvc3Eggo
EuNlBqzgEn/O8YoqhVnR+421XDgPDp3+4AzM51cBbAFA11KZMPOOvH44j/5Trh1u
skEAsGmtylGYRWrzrMz2kIDxmKQA5EaOhAFJFtpxQDC14r5KGDbX2gPpHTkgxR4W
lG49Yt8qfV4BrMZ4UgdqqWPeW7Vpsl08FAFziXFZzJrQ7hHtZwhRYann/lctNm6Z
y5v6Z2HDLyxry8YREIVSSIYFFe8FOBmTzMm5Qp39Oc6Uj4tTDgxZXkEWgJUj/rpT
itjxTUvlEn923Pe/eDVBOs5R+rOOW9Wl0i63UjtukMn5elGkcFL7L/V2zHi5YHLC
W+4lmkstLeh1fkgRnmW4Vb03dC7ipkcHnnhwCGu/4Sb8rDSglFDI65jBytKST+k0
Rp5CSr1jIrR+SQ+AYkXkczgRv29x7PeE9onaCXTIKLSaRDJj1M/h/wb2c7r0uN6J
kvmo+kUYnZeADCB0hji/bAUne/+vzD67kqVRMhz30xxcDCegxdXok6fSafX7nfhO
Ere3lw/hnwNrZQqICt74lPSGgEHZrDa+fFoMJnOW4JT8IzBbiAochp1QyHOOPjbf
ECQOh5g8qQIzHHLQuNhBARKtP4GS1sa2xkdK5/QgiEFjF878zI12xi7LkVHZQxGj
juw85j5w9DGlAtvFEo3/DjlN/zCSfpMLaZJBtA7z5c8kWaTlNK0v9v23hhG7l6z4
6RWmcyFNAOJDYlJ3mFV8c9eqI5hftfHBuQ8mAZegNK0HUg6BnzsKunmyXMKkWbqp
iprfI25RD87xNFD9FolmW7BiuZylfW4bD/RyBnMZgCifwGabWWB2qSVO+8Pyno+d
kwhkgMCj7KYSokV+a7oL6xDUKhyOavrulKwTC9m7a3fdtserd5KjYaIZQpSY4fUX
j1RFokWghJGzDkk1JC0UsV6w2aj+5zBKPpqywPYq/bKyU1CCudwJnqWi+e4vOs4Z
77/84hoIiZW+aRz8XbDAxjFrmL3YEWjMKpV7PUVTTfcFTqy2x8itJe8VP7h4RqPk
nV6KxxROaBZ7L5nAShltAEvETdl00PyQObLBbbCtDDGXLaudWnTPZm9rlGDOzc+i
M2T8WB1MOpBVKBuObvLqpDPemOjEdTnfVTjLH2LnxZDN5/UHcTUCnA7vwnE+DISc
a5tuupCeBypdy/HaHFuwakVCDZ8eIibVWlFtAk0seUc3rQYfMxVIU8Dmm3D7tkdj
dWxUVeU5SE6smBWHxfJFhEpGXteS6/9QuX1Y8XUHW3m1veVKeEaOxcSlkw8hwdYF
OSC0Ey7goo+7DttDPHytvFVxzo4vuAaFFDuxFKb/sUpEzdvMfH1tV9EvTlFf0jEh
lrI+llnFPw1WwNkprcN0502Ey9F9x415H3bi2tqOgzzCQBAN6m/RtEZGVh2Y1aw9
0a98bxIc25kULaZeXR5XJtBT39RSp4f55A49wh4kYaD1vm8WAI1RTx2M7nYjBcJ/
9130VcTmrB3Wopm1CQCKbMOpsDidOOtDzJNdmDVeO11DvO2h+Ms38mWMYwn511qD
Jaa+1/3/67Sd2fEPl+FlDSR1eeW3QUfgAFnI6Wwbs2TuXsl6mM/jbdRTGdsTbCP3
9ujSiwdKt1cN1LBUDazpAMOJEgvqWhuH/k0+nXp4nw4Cm3X67EzNFN1j7BRXU2AM
s6CTEFq32CT/sI4T/R3JhYsKUwiPlyeMam52fn3vgn0/1aOE8XY2TwQ5uTuyfCQA
HSaZDM018o9AP0hvOW1LL9lptJX58EVREP/y5rORNgh0Ccvt2KRDWAoXBCv3XagA
NXiv5pddEf3wydWkk7Vl+j/S7+yVVsDITK5CCz1qls3d2mnCnhW1dmogfjo/6blT
M1676OLILBENP2ij/KBf7f9qLA+x1wGY8Sbrs28YqJI88rhCShflAwfH7huZm4Fb
+FuwcxnG9YsqFXUoNnPUzjWKeT8mSUgoXjZHXyzVCuChZMW4gHqMG1naH2FjWnKY
qqj3h7lg1dDp62xwDJg02lKC07WSCNC6k40HggFUVnKOZtxSgZq6gkodRDREAUWk
uh+mDMlIkdKLiP/AFG/yMSLkFjETDJblTT8syajINhmNRfmCQ0iUfDyovfKv1DPX
2y0u/wMWHo0iWluLZ9czgCIaeYM/h2pNzda73JbZZnXGJZhgSIrOVrCXOo2SFU9b
oPJtLtg/w/QJe2sAhcUcS8fTpozl+YC2mjfkq+irDwvxoVlfQyYe7KUeJ+QGJ6CQ
XkDIXB/RAmPk6dsgO9OZEdJG1oM5l7cNOzsPRkKnnNlCedQcbv+xYQzWSqpTiixD
P63PEGAMKdpxNPRcvhz7WNRGOnhEKl8jJ2Lm6uc7f4jbr1r/Jy91Utw/awRfoCA9
QsGhprgR1arJREGMVTQurAEIX47Pqx42Ov48MELywvA47RJshDRJlVzB0VayClag
uL0hrdXUwL9Qi1Q9hJ8czRBr+HMgyUSx5s9g9wrhNZGN8PSPO2FYCT1BSXKUXaW5
lcAEeZpVmaUN9TTWLGFrZKMMciu6MUegfFbxZobhCZgg/DSo6Z6hwUQC9xODiDjs
GMJkd/etsog4HFbsk82Bj4xTyanCG5FNV88T4tSi3Z6O7pWpmmSxr8Khlk4ju4N0
QQIxmnc9C1O9mzlxjiSq/pcUj5CCK4JnS/CkM+Wi+iOJ6K80tMRbo3HZXV/E3m4K
kQ3fP1a1ed+gDEaZoF7YZkG7Scd4yL9B/cSDKVb1JdQReERHU7hpYk/i4732eFUR
A8thvSAlQUHovFyXK8H96gxjXGYqfYV8sMpfYjEUyf2NurKxjeI0EOyC+az+fokC
OA4yBDr1Kdm74IodcQgsokeNycdRa6RN07797HD9KHJNp6hitYDgRsNlLTnfJGTU
PHQamkhCFfhx05ajOUshKTE2bOQJygHgoLYnSxan72FvYZZWcjawNw6IyTAlxmDJ
4UuWHjdZhX9VSYfplBW1eYM8h5wMOHFN1md6GmzCmZj64UOByztTU44Br2ABNNuS
/PnqORwVU7W4guf1HXGNPqeDe17A27GtFoBy50u8/ZJAAw6hO3EocWwDtoRonXhi
WKHMcqUZwq7x31dY0tFNu5lLk3OGdZ0MOd6NCrFGQJQce5ccExhSS+oxL/Fipr9d
lchANzroKs97N1Q9tUatY27oaafrHmaM4Y1XDC7HiNwA+oGCUrxdFTQrAFU65T4n
lwpQmp7LthuSNtUNkDrUj3wP38o7avYlnT4HnbAq8yu8eCz3nxUMIaTTXsP9JljI
d/ARz/sTxKAbVP/cnOM5U8JouKA8+sO5CeN8uKgpzn2IDMg6VPnsLqFIYJi0wc0n
IBX6A2EGLBXt5U1lUUCl5L4eqRtP7WHlhlBwAEw+0HAdRDVyKKUH4+Q9GMoj/LhZ
ThKhxLQQKp76zODlN6SDXFxh//gn3GtbQ+U1bO0LB2+T6qrrp1gmjGDzmcKzlBeu
SVk239R8tBsrWUyuaeH3TtWp6UpYzz8N31OgzBlpIwE5pMozcV+CF3VFMtk3m8iy
Lz4G4oPe/FNCEipuvs91hUzGJkn2TxKk5sFKQP3of7lVfEUPAx/7kQtOvCFUnIjb
iWtVT1nG05SOnhq095I214ShBW9SfA39rd8bD4SMoxDCnHxPaNC+Eu6Hx/neHsB7
RCA1W8WkxDIalNOyC2uhJiv1JBwuvzQ4JTt3K9l+wRyUZtZJcLiWod0gMpruwtNy
ndMLpiERTV4m6g6zqbMb27H7QH8ookw6BY45KcXLNbo3jA5lROVpfOARssolvICU
CmS7b/IMSdYnSjjl9DlcNm1k07PACkKdwnsDrlQpp3za4gli0tT6zH3tD/ov7dcC
KLxJJnFqe9PxTyFsknjhI6KYF7a8FFKqzWtalMyhUyVd3hk7Gh+t3he5TboWaHZY
enzPvH4R+Mcpg+2pkyBj22qGSqLEzwWcFgWFog+YCYyqg3WFpompLorXs9i+TEgM
xDDhOU4QwwDa+iJKCuO6U4qZIBh0Ar5LxWJ/Ycjyoiw6pQA4q8TaJnwlb5bEwSDE
7Scxo5TPOmLd03MxDXULgikLhapzfxrpeWmbMUX4BYg/u8M2quFouNUfyhA6+/DL
KZRz+ovf+R/Snur9jTqhma0u/dJ7AEgWl9uhb+oVHL0aGbDbN2NNoG8Wghq5qW9+
3VscmrZgyubtfB9stLHJl17mhTl6Fv9fnJh4HNPyv99U6lZHJmkON0LFEmcYMs7Q
mIiHU+zXS5kdqH9MY2xGZU8zPeiw6++hLxAe98Nxj8woeqQUno7JoZ7kBOnWwziO
s3iMCgdQ/uulWHuL06rvXr8oXqOOqS+Yyo+pHdls82c4CMINMNTzKE355fk+Rj69
xKa+rsyMr11rGKqYy2yidj3nXfhMjIbwU9mbqpcLt4DyQY5uCRTEy00jDQJdVG0r
p8Kk3WGstLmYuKPmVuEvKzgwBKGyvlwmzHEgytPyqwD/IMfZcE0KJHIr8THA8+kp
Rmyjy/FORDmj4VtdEFfP+9ZL3bquM42SKIoEyhxRyV0PbnK6vWHW2UPzLehaK5/e
q6+kZ1w6tlRt7j39tYQWT6HG34ryEXzTwHfv9RyQyWbxTcs560i/q+mJJDeV22pd
qZWBPz3voX02SuFxX8h3/vWHk8KY6Djn0CoCCN4j9I2NukyPT/aT9q8PT97cP0NW
TStAdbiKQkjgF2z1ATSatB8qyJx1nqTZ7Fk702zX1KF+Kq3CeUJ4XRI3Wr6ZTYT4
Tkd0aqd03BOuvtu5CJSS2oa0PZMEvc9oBy3I/NJ0iyepIpEpwJQYDJWeHEouafKK
9gZzlR+i+He9DuiiQfug1akkfbniOh0+8zNn2szZ1N5WdbSYPcMAodF4d8QJjUO6
aLWQ3FY6sS2lh7cPpSk0tdnKTcp4Agl/cYb6e9eKaGX+f80yRRJiAmsrT4w0Fjm3
wc6VcO9+dQqBFuMm7r5y3L0XItCTgQk+XoMmR2gjNQF/hHKTkuQoQao7kTYeKlBt
tMIwOKSzSUMv4NlE6sj7lQOq4LVWx6+pjm367PJjgkNqUQdm1Pd4iCENxFmtctEh
Wv2p0DHVpbnjiP7prIk44h8XCCqyGOKb5j73UP01c6VdB0QBNLzu0PQXRox8MKqt
x6q3VC20hPi3KWqyoUvRw7S7TfJ/aVFADOlj1k7msJ5JBQ12lYnY8lEL18tjyCr5
rRXKfUSmqdpcdEal0XLfTL5rIgvTjAsba+SIDcnXpxGw8LFI/44+OPhOuMrVxbpO
hyTlLi6RjNbv10RYE/SHbKZkOOjmkOn6O4UOS7BvBKC+rukBnzCxDoiZpFDKVsxO
igj2nYX7a98zyLhlo1QuCkTenE6BvhbG+5qvB9Np759jJRMRGdahiW6HhHAE/kl4
Ble+P9FwCEMXx2gGcliagGu/WokwcxiVGcmvfEc3lavG/qHA6SczG8e5jCsBmh8s
POFgPPuIi9iPQkPKVNJaJVvon+YbulixWDJEWeqDWMjYZsmHYJ2I9uU2E+gDewb6
ASZY10vmyM7l2GCdR2fmuEWi3O0TU29UDzqX8R5ayZRrHeUUc1xwjMLamweDeRJO
sJd3mhQU4EIpbky1D1QtBmLBo5LHEvFa66dbR9e2ISjf2bXoCL71nS9CsuBC5jr9
D3nxwa8Pi0P+8TSFoa2vBbDUOTmXYX5NsbHhIG5SiUMecxD7VP9R1+nFdOHsFbkk
jpwyCHUPXbyiHj3tV7C8Wir/ei0MwmmxNr+dsRPCjbXHen6Miitl0DgsuunKcmMg
SMMUMNOgFEXkGxdgJ2K9D7/3ShPHaglI3CGS9CvtQ8fEdT5EQFUETahBL4OjdPs2
IPY0tiTnAH2GmqnsaHqVrFGtNJP3Oq7iSuxQ2bqhjSIy/8CXVSjm/GXBRvjmjlSM
fhtuWjb6Ai8PGTD9u7MM5ACzKzrD88FEZfJKnmD3/DACJjyMJ32DYvbikx76iNpz
5SnfQbXDAmwRZTKCgZT9roo/rMxjjt9vDYXPwQMSMtkuqcPgco+kSrKfYK5/HivH
9rAWX6KHCvO39XlxSbfZfYirEqU/l3xVTGmKdflf8PG9TtQUeH2j730cowGWuLLE
w5YFtOKEj1NcTejdw7PRRZW5baZF3qoAmkFnkcj7Gc9oNd8WXO8kiyZFciPCnePY
9jQHNh0XqKeEhSKWY523nRzLTWoZzkaPit0iQkjMmPITTr+QSI3ZN+GataB55WF5
tJ8tfghe7cH5Zd09SXZX6D6xbOlx+qYC0nSTYXr/2c/TLq+9gw48p8cEwJRGEZI7
kIbGspjQzgCktMO+7LiNJhJCnzObhxp8ZEFp42w1aqzjV6rh+6dk6KChAtc/tZbn
BUkq2M5KK7yaXe5HBMhsAtnKJnvN2e209qyO6QaqU940QzIytSyh38j/u3KMrYWZ
honr1dmQVPjOGPcoAjAIWWoJD4JIhfJYkIQjXHhh15WwxIBSGgMx7UmSoIlgp5xl
hzW7sZigNtnUqMQies3zTuCKk/k+O6/Ky1FzXG23aLmt3J0twZac7+xqhoxEnNBD
GQ5vv7C+ACOWDQ+4jkyEqB1JiDW70MBZA4Zt3OPQXiaS6Zd3sMPX0BlHRdlE79j7
abDzNDhNoIOjXfzlRQHg+uVF37HXSwZTuSRIL9OjHVmiwiunDfw53ui7lOCIJUYK
WesDEerUcbd/YtvG3vcDo+RqzXWFH6GqCwuxIy6FhnZZgCyLRIpO2dmkLFEtlXJg
T5i7ivzj1EenmCrZl2LeE2fkiStUVOMr8BYXbfcx/KYoDWemxvww4M1d9HerK5MB
v0hHPUrJS9924SK7qE8wR1s1tmKkdsueLXv2d/kCBulIMQKqC2DRNrZnnq/8WNhR
mFDlSw4XzMkkr60ZcutvuFWb7SzD7Za+oiIQvbZEMzHSWOW85W1LTOgcGt0caWc4
5vsMrq9d+/cSJaqB3qEYjqJlp6FopKu2LDDgWdmQpuhjFeIEl5WUkHwGdxm42KI/
1eNmwKF7GqMYlQbydjpsRwKZaOEh3FGa8SEVIRz1JmwYoUPhaxX8PN6u5VC3qddT
rF43Ak6bg/jIPDmnl3Hv8FB1iLElgi/dMpKjBhkm3WG3gIzXQIla2iC2pbN6p9qC
QfXAFr5SDmMZ49V483ibPtjkL+rUsWaY7e0ayzH8iajbOymXPHHmESWKSNuPCF8I
py1pgfVd0W0QMYO/cn7/DELv7I1JCkVYdcSswRsW8UuGNaXBrPgM4n++5OUeKh5u
q5ootf6fZtEDA+rRNq6oQor2W//74BDxVdoCkbnanXbAkN1huyYpnrjO91HQ1xLI
dD6GjryglFBw5eKg2X/hqFfwmYcmIh6AMOOgiCjYzzlCk6tHvoBLV75qFZMkEww1
qGfmxldBccqACI3wq0ks5gYjU6AhhFS2ng5RUL0KC/4y3lDds53PjDYOZujYghhN
BDoZoBoc/AR8uwopKrCMdz8P37ZxvbauBMn8fyRHWK6VKMBJTlxMmdZDIUyDkn+G
Bh3eeTKYncf007hcDxVvH0xLtZB3rPmtimS76ltcs3+ezlt5XY2MxRQ4Y4GKI+ZF
GNdZCWw5y4Y6Hw1Ipr7nzrPS9wEiMdK+Klz2tXeC5Nxq7tn5X81sLhSCjWtAGCJC
q7A/4LkQZJYqquOWDsUkoBuXjiFFS+xCAX15DIvq6MpdsHw9Xe104FGr65NjxJqE
ea8b+t2WKOArAHE33gWOG/hTWK2Gp7bEFPNAtN3HIyOlO/AwEp/k6LihHCopXeuA
VbGjBUt3Cme7gkfT6EPbmSlrMtzd7ua4ZnthnjS1ET1aM0R7zPnRNiW6zPkYWg/v
R1ao8+rY8kyMLqwFrz90oYHmDorv8wpQUFT0L2qxpmz0CjqC2/S9i4/e4oe1emr8
XYxud+yF/sUcfTnnapOPDs3wm/02QD5aLWSkYlb8rK48Ndp6M3vbjluzXtflV57G
T0I/YgNTMvoLI7pdvJfDPmLleEQqgigz91qdiS4eq0gZTD6vooERkHpz9/yi+1To
dtVVJN5l6n+4DM1t6r208JessTehM3b+wmC8eY+mRoNZtr2qfPwPkY2Q+ug1LCUa
jnKA0GjZmjtjIAKKzvdDolC4bwwzRL6OWynzWj6Ge/CCnqwZ/fEQzIWcZksIn1Ab
byCWJAe+v75J9vUk2bBKtYZNPOKEmo8qzVqHqO/EidFA5xlvHdnfSa8ZRxdgi25Y
rOIRo35jbCGQ1Nd9S0ItGWZSzendmpqqF11EWliKN2TnjkbYbsd2l94X5e/krRzn
fmkLEB3BytztOu/KHqF1jWfcGBxRSRuTVQKmOIrhmeno6rxE6yzW3j2UY1BtdqKC
W2qEVhnYzeAdDK8udrN4DU1Kw4mRjw7mNpUo+fiQFraqGJUia3BQOEK5NLRoPV8R
xrN5Gn4P6d9fco0M1X7BTVZOp83l9KaLuq26GlWhnlPOcl+nmJUDCOxD+CUL3sga
2uqnIITkEuxSCg10t6jY0MPEuaAYgfmEJplNxM69rTI5TDANlw1ByicZp33e/9cb
Bgi4lllF+qhlt8wSpgkKR6Jod8ZdwIiVb/xb97cOjuXk9G91iXt6qifEBcDOsX+s
035Ommy/ZuMiNQ0nbd3H3Rj6BXIXgeeVSbWt5kZZ0anANNvAv/mmrPLlz9kpdwYs
HpjXsert1StELuOehxOFGvwJx1nh2OSfhB1fzTEH7BEpsFueO66FTO8F3H7NFi3m
eehMpHOnoZwmPugF5qCxSHHVpS4JCCeoA5k+Y6KgX3u9CnLcgMcgGkXZ64wh0qiF
uIZ1MIswm4tWxEu8kzPdDjrYU/iN3qazKDxmVbzr3I2aXhxO+YoifGkXrUb2Tcfe
ZcG8AyWfwh79KhIh0UAzvCuUph+osCKzUFVuhtDayNIXMWOI/U2ZE4NIW7el6Nd+
wj3HP1SNL6LV6s4Irh/NatJWWY1kaytZSvbmYfntnmidhyRBIyQEwDkjw8v5FlIm
xmFTExXJJk9SCK7gp7BwJ0AeTjl0n7C6GwLYzOK2gBvP3F7UMrdMp5S/xSWL9fpY
+8PCDKbJF/NkJxmQ8svehO93WxXKSClJFIJaykUhlaK9W0+2ChkVJg/0U+2pBJ3/
dNkMl5LpJ07u08j9QVZK3RNRuanN6icJJkr7sgR3JKnVICjvu9PZ0CM7VTvYBJDL
m8bll2Rszkz/BISYvtPEp1KSxX53jmcnwDI5UtL3F+ClxTdMp/VPmTZ4KoM4eCaz
5H35vlzNUFLUAoaua/4NXTQ04/iRYMIchs0d4UcFHOu34anSm4RAZx/UpehnqXO+
D4gEvNpOC9Sss20lX3M3EnLrtgrEJRj/lBcSAYVYLXweYPyaCz7tV+XPFXjMyQpO
gWL/sSoWDCOZwUtIcZ1TFkALJIaX/aa6mDh2FUmoA5FD8TGYgrtHMhq3E2lb50ET
PwOPT+FcsB8hEFnxKb7HSeJTGF28ICPQ70JVRp52tbp/24bM85zva4nw1w3Bss/A
G38Ans0dw8ovSf1OKSgz09oV+itCGiZf2VirILNCDKRji/aYtZTvoV01LmSU5bIa
vytTAWj+q3mFTjg89Zo1NknP3Fb3cvqKkIHAxyBedKCTFKYPDYGY14LEVLmwE+ce
6ad3o681p7yNIbeyzDIxgv4Gnj7WBAsI5Nl7uv6Uaf2s7JclNDMkUxnhWuL7jznJ
aKQzT0Jg0NwKu7DuL+UbQDZvlnS/505dB2AQBQvcIibvPWDq37JlGiqkXkZfpOv/
QXUGXjXaEIxIFxyd2yi+tzJyO/TAotfnZXqIkn7zrg/KgwKo8Igb7lF9zg1ouPjC
8ow7OPWMD2CXhROB2BwkKnfJHydLH1erHaAEUed0VAmNzc/ue5ZJvdwb4uP7n9d/
cZ4S27tL1EqoJNF3YDqrPxFoy2AbASRtOk3KsA838Ju8xVvsPhOVN5zfswmXXDjy
vhaKVDknEi2D44pc9hTM0SS6aRbAU9uht2KTjKyRZJ1S40ntdu35TIyC/McXBGBy
eW5L3HC5aF+O6E5jDTEV+hrQ/AM7mmIE2YTxcpLDiyimaosXFXxkuApChGJdPbJP
qvmKvlKeW+/0VrYut1U2aenlCOGQreQlRkDJZnea3tn5LqZOo6bcAIA0cmC6LPS+
vN8RDlmuq9QyI6/L9yFn3I6gEcC/anO6E4LS05pN6n+Uh3eszELJ9NgRL4kjHI4G
EV3cPpxwISflOIzTC45NN1Tpgk8q8Nfqh7MQZyyB5VoZZQuCA+O9PJzqjsHi9M9P
uQXXSy7p92b0Fl9hIblaeYQlxWRPHzrv7gZxNypf4gqYx2c0YzkBvdalVlaOMONp
P2R4/cWe/c8POrQl5qWQuWIVgr61OZjmBxW1xoFyulS6IWYTLmsxwAO0jDkIdu1R
bnfJC8+B5z1g5fJVy2hwI698oH5jPTaC79POlc0hioXbCtYjyNvMAXqsmGYAKdz2
+ZCHZwFqY/aqMChkK85OZlVPLgYSzCovP95egyOYxnzU3SAHoT6nsA4youSoMenm
tROdelk3zWgDzSvaswbZuVh5DetRlPrLgfXdXefrRaWBJu1Pu5ZUIOAnOxv3KicA
vE5Hw3DgwHoVJ4yiq8oWJ/E34DHV6P8FbTp6xpJMz6hj//VALcdTCq/CsJDbNg+n
10Ov2DXKYAslG7eKf8yqVT6EjYM9n1/z9mGJAczh4GgTpxoq7mZo0VqYIboBnMDK
TIYzuU9Jx5kjZnroEv14ieB8TOxk5pqQQhogvA80pnGof7gUgAq2N9oy8rzHfmar
zI/V/MnY+SH3A6uKOcXUicWiMbyGZ4IYhDeK/59VSsMXxjiwuTcfkzuq7waPxI46
1S+YQm4S3m41hRbC9oo6dtmhMBpileqQiyXwRZa0dejYti07lvgA/VInSxQ6KDqB
N45TpHWqE6uLohO7CM0LVxW5S8WkCH9PWreyzl50WKQ+22yU9o0VRL7l7DYzDCZk
mVumghT1rkvWyAZ0+bTsNJ/jfk7ocx8kT1qejw+J1057cFf5OBmbEDXB/z7p7vc3
DNgnnx0TYllJFuNzMpAWfHWR6+LAHJb/Sjy5kkOuyb8h8vGOkJCWh6nnmrkDriDR
HPgNMTgZmJRRDH++kP+S3dpq+fInkLmX4R89LV2NqcRgMBQd3SXdSHZYKa4N4m+A
jRCs3q0GKo6Zha2Dpz4hw9Vih7UvXkY6Df8i+3DomaTDED9drBIwV/Mn3x9N9qvL
z8Tj/nqVNj/3z01vCMBECbkd2L/ETLQiUK1XxUGrHWIoAe/s6SmEYgmlZVIJpEG5
N9gifhqR5GO+V30l61gmS0KNZWYOItgUFEiK/gV8QMtQZdWqbnuMBUxudszE6f9T
nvDYsgSvWJf7Fh14MTeq/YZ4qbZ0wkMCPLDOM63UL4ksMJJ2ZBMIe84ogWMKMNBm
bIg0cn05s6akawPSyMrvXmOxku5g4HosRvAxzM5OgWJsmEppgo1B3s383+S4Fkub
hVBxiwGZ96bGyLaZwhRAIouS43TGgfVMfuNWYSf7HJsTCGNlR8tXBrXcoByc7Qjt
SvVRdAAQOw3X0IODq5CX8/7tx+fLOKzPv/xKhsGH5RSEq27BZ/YuKOPjZNYhig9B
h9hZPmbVuJ6aHeIv4flZ/u90vuC508/eZuRYOuKugokNEogtVWxjVnPJyCR/7aAC
LQJBnWb/wj7WNqcmFXEvy00eALR4CyOTETOtRwK4qC9lX74/ES1xHCsrNaVSp8C7
U/0S6yiITRdWQrb0+LDiXICkzBrhk3VXHjJg+qmYxk2uLYE6w2FsivU/pAF2jkNG
JhyMyta8ivzurokRzpRM+2YcSwHNAUAQKb8HlInguGuaBRCTBm9BmEHTodfpzpgg
j+0G7SqOrYYBCljC3dHmmVk4UPuhUTOTotQyEoT/Fk4hif/EQ44KsIFewqwlp9kZ
ddzpeYP6fgbste5lKk33wY7UjReviWQYIM4sIUdFyUBrEEoX3OtZ1/3ywoePyorQ
rbkDiDQsN7S7+FUcXIMlvLHzfppCbJDHmNT65C7fqzWP/S/SW5hmqch9NJk145JF
gT9I6IjBf8dT4G4g/bCoSzTPrxenYY6MjImNjsQ1N5t2XKHxMH0h9+rnpbD8SQ+T
rwMcc8aSRCWnGyArj6/m5iltLO50m+pcUgzNJ3rCtLzf6oknC1OevZY5yk74E4aG
zD/sVPaacF6I8aZPTRLqxGk4xTqi3MiPBpj2+P0Ws7kDe0bgIIrlI+JPw2TmgmM/
07LyKlcyaaCFxZCzyS6peR0mmCyF3qon0kV9xdBfLjFdhGlINPESPYmwjT4o3cvo
CkLyNON0RU8md49mpuQBLbUYK3xO3Wr7lPI59k2QrPDky1KaqfP2Dn89gFpoQ2lk
DVb68BkAUXT2X+x2NQHucg/Ocio18vdBnWXu0iFMOaYHH7BI3V706GKESenatFjZ
+2oHbe7aE1cAYnsS1uC7NtXME7U9ASpKsmkLykhOTS7Yg5WihAaeNt8jx6ictO90
HD4/jABuYE2Ps4dHu2Q+vUR5UD7o49Zg6wkONQLddm+MiLMW/o9cwrnedi6TKrKx
dK+8SWhWi/nMvJLx6wgtT8H4G/vsZyfmqnyTspEQmX+Vsxa2b9MOHhz5FDJkfC30
4HDoo/5yNbVMEdrwHoTHJoyyW2KNcahprNJO4PZyPBkkSqKcC7ft6Uemiv/ribJf
8DBxoHZ/m9o+5aWr9efEX9hEDfZGuKRWB9MqN6hSVE6lPGWZaQ+3vgfyqq5fMcZA
LeG0dNKellPrBsFsCDDlbuvSNZmX3yzAbM5Se+1s38zu0SA6uls8y7zU6W56Yp+D
5gdQIF67Ewu0jwHJXSBQiQFVU2z5K+ictFeCLL5TAClS5o8ZS+tYcD5XD2SUXStX
WldxD6PsYnXhVW+FXv1lVK6bX/+DDbBn3p/oLwAkxPABe90QJqKv6GyGZ7jR3t9b
oO2VkQ3i35Io1RoVgPY4NU8FrbLsxhOlxZ0Ixwl1Gx2RGhr8E3miPDUD1xUkCxWK
ZqgKi5W7YeaXMXb7dXgG5eqEFOT3a01vHupmWFa0A999R5lazcQInHP/PfTwihBG
RqIMnj1u4sBEB91LW/aQThqYNOVLgnEj2a2MCnevJyrcH5jdFjHwGkm5lVTssvr+
bMwZulMHojYklDMugnViGosYo0g7Ol6CZBvzbhxKI59WN4oAWMcpNXMj4tbPeGHr
ml1aXFcdqHL9CTCnPWgOO1t8sy4vM0mqqY5VlbRcUZyMLc3DzmOH+M3vHS6eXO4/
ZNdsuaHyIqLYPS51e9N4KOYj1dn2Y3MxUJZOXDFSnJ0m0+SrtRe83tfwB2YQl6e1
x9WLn1OEJ6RD+9OygvQk3lCN6N2RYjXd30/niFGoNhzMo6R/6/2TwGIdaX9nnNxu
bcUVHQQyscFpQRnMmSBQuF9w5vUccLTqm0ksHWCU8RpkptfUYgfbHfFxgNJZeW9F
kzJrDiI3pEiIBTNg83dZM9gqUp8pAGTbLKAixZedg/butRsoRcLnEUWjWhfwFMrA
7ZP8pi6hwLAbbjwvupYkCLs8CB1Lk3swQ/6/MsBwOpCH4qqpR/04PqQwCj1qtpga
/pu04jWkJcx5PYv0rNFoU4YZnMPgvvLiJdpxDQUQyp/IbJSnBx9LESud17cGs4iw
EJN4J8e4ZPv3cD0xrShBZkBDLO0FbSEIYsVJi4kPNaZD6OKEw0kz6X6X0RGGb9yV
qZ7scjPZX29z4Mvv7rMOOQAYNXhaF/n4XQhH3SAFJfHU9BnSU5fFvNwUON9lb7cZ
Kz3xanZHf3GpKZxmxMDTdx2H72p9TjPdhxCW9w+Z7JiwvEeR8iPn0Lnu0RXdP/r7
F+ZEZbU2AdP5thcaoarc8UUCNns9IQiJbngZyaWYov7UU1FaAbRxaKJQaXnlBDmw
vCWzOVe76r4F2ZPRvYLOgbjIEitxjVC1kiA9HT4HoWlBQf1y4X7ZHsrq3kVVW4RI
lSciLvKoRZtkB97cpe3enGYcIvFnat3mG7it1AQ6MOcwEhpPT+TujbOdUWYY6SMn
ipq7bexxq39zkzPD8nNH47hVGq6eCOc44zxp8OAkbTKGgqKLwuco2ECSrQujgsSa
2XNbsC5IxtQwZFxY86rIzSc1TmRawNO3L3nMiA+RsSnxlgBeTEXajIgmcmAE7TyL
BSAvTHJjB4G69bDkDgw9QFNf8GIyay33tnHwx8JA2si9+WP6su35+ccfEoi00dCS
NCRv7Ooy8AT/tUbhkb9imRuCqQzDYguLMtRLeEgzSZ7gW1hsotOiLkJL5WTctfpQ
B6ucMogw1ZaZGX7Sg9XaJwfsVwupTnNZKV5CDuMvDAgUvijTsU97+8zZJFVFuh7N
Bx8yAOy+ux7Bob2A+sulARis79wyYg/V9JCKmkkpVkEseaOQL5i4NKor8ZoZNUrn
jACIfql2rCTOMSozOWgsrDfdMkW1l8bAFp2W3Dn+sGqM4Ox+aOSbB5rpj3Lwx962
t/Vndzs01LHi122IYAfYwovJY8/agGjJHbFF0VT0JArtZ0Q3q1OLT6txnFZtVnzQ
74vfHMWFiMN5tEYFg3N7Wd4d3x/XA+sJo8pdTTP3EYVQp229jxNkBqwk18X7JumF
5KiQbU7St+V4KpvwbOFJaQA8QwNvtUQis8B1WVN+Dc6CQHaLHxnTs0EZhcP2A3zY
OGWUFcnCRckc1E6fVbWF/7COIysia+fPlOpkEXwZiCji5giezThyhYLHbhm7Jd1z
6/AuEp2CQtbeqMePhv77iKdDwFEte6Dic8U2Nu205UsTJqOLrIwyRWmYpc6zSVN/
/DGeDKr+VCoAAle8W/xexvcp74byqRsKNN2BfkwiQ5Px7wET7OuKDxIclqYbDAsa
fiWh5yxQZzsLcY+6slN8C4PtAsB8NIPlLENV8H1BxgWmWie7u5ZKtAYovOMcI7eK
qZMrpAlP3CK5bU0ISiJVq4WlRgUm533sJSeRsKSchbNdWGOQKfdPq1bEoFlnmdH3
FQQb1qZpF3GYPdc0m6qYWQ9LjthkWMDml/MOq/fMgKrHtF1bq0y3NJgJhByuhjjN
9cm0Q2XYa0c7UkU0X8BCw2GCJzY3+bCe8jJs+1foRGe6XbqWPeNvJ3qdk2/k3F9m
7Ow4GKUtOX92NA2EzOgOWw00RZzhJ1U6SfN6GsvGHZTWVqzrQv36/C/TRQc9nH61
M9dwoMAYc5t2o2xdpESUb/hvt0L7TfwytXCpCsdrt9/SpNR39kicYVeKilBw+yJ3
GPGCaBfo3X7ZcXXby/AKeLKqrdrJHpGju8IxQ9UrfAr5jTz2j8yPWa4hyxSdz5KT
Tz4OkckYqUPMQQrdX2NOhWpVG1w+37VLk6Aignu0PvDqq4EdeV/o1/stoxFlhwIr
LXwsMK+3Kek8phpJyXSOWaf+n7KWoX4qxw9n4cSNN+8IzT0k1Ut4kebNOShC3Ghg
W6CR/I7XpF0mZaCpauslBg+lnGI1pH9SuW/f4DKWT8HMUZ/HnPnnXPDHIPiANfpR
Lk1XdKBdz93kHFR9EnrkprsMXQR/4Jao8aE/vNR6Rr8WtA2v8rqGZA6+2Tqj7qvr
4RICcj1E0DFHDNRH1zu1H3KszOzKsHXK4fJ7bDm6T+OSHOESXI/Meq7jVEi2VI1p
rhYmnMZOnMpdJUXK7h8jdlZI2sBAHh35WagIBq6aeS5JCyqCXRmIlnq+hp196XPq
BzV5vHFPDXGshvvjJxIgtPGCdVNy9DliTz+C40DOalBV5hTBQgaXN812CYwA3oRF
5JMjWekkIsTshC5DvtcnsHAkjSTR3LOxq+75umy1q9lU/i6v8DxE1DCTvQCXySxf
mDS2Tov6o4b5b1fSRHH/BonHe3EJt4KDQL1sVNl/eSrci4lVGeVaMMCIYf97uIzp
aDSpw+iHAvmhcYnSJuvBqA2mRIBSmsBc98Cb4bQ0qka5ky73NXiJZvGxW42Cacau
v+lfyoeBOHXUhO8WB3OFS90ozxzo/KIIQAtGDjZOKqQpJgI/NtF75sSPlTwYzcJc
WbzR8AIujwMDfI8chCZCS6mEpvs3tL7tm13xHsqGGXRsk+J8Tjs9EgvhoLg3zRyA
ip4lXp3v9fqnJaj1qWYOWyKpk8pXO9kpvcGTUIwQDO5oDVyOq+QvqYRK/SBS8Wjv
FprbCNpkp//lO/25PFAxiXVmS9OcK5Ty5tibICPcC/2C6SsJGAwEoyCqnblrXHVw
gmZjbXefcesgQHAAbDUa/sTUmYR1vGhG76TwQmwuH6DbakVZi+6E1FHMYzq9f7pn
p8rl64B8Gls5fFLHS/wglGx9PQMap07v5nMAag0hOdPJHK+wfx/vhu9Ly9wt+rlT
xPQAngvi1RTBeTG1G8YL4MoHYiMkcFoWllSD/8csxVMVke0xOWPGjHjAEqpcg9/1
rQ7Kc1+OEREcpQFXihHrWYD98pUixF0UPz7kqH7yHvgqGUNAW6/tCqeMkrLLuAtB
VzfnaMjA+UhgGg2R2mWalXBfrVyyT3c/Q5qKhlK8mpCTXqveA+y46uB4SQm7BPuX
VNF/RomfLV4daA+Z9Z7vcW8AkFRCHMgBv459RuLWHlU2oLsV6NtK9R1QlrJVNKjF
Dc5qPRRNiK9E0QZ2N8awe/5WE1k+ZzxhND2cdnWXd8MJUUshPWfjBH+xN+5lZ3+d
bb88A9kejdGFVONRYpuKe8nGO8IznobgHdNzu0LTEsxGQHvm5g1zNSGs09huuZHE
uYUEHqBK19AxeMzjndBb/MkTw34PU0Ev7uA9vnIOnLsZ6+9vEbJkpO5M/Dzd4gKL
v2uMeLyZRjmaN7RqG0lHDyGysf4e9KqBnnqIel2MODNzLlv+8CWQhlFpyAepYYYn
dpubOBg2qV/uk7PgvBvJHhpAtCAtHuULCpcJNIpQc7vM5lF9jkD9ObQY+szLlJh1
LzFsiRzTzmhV4B7zUICAAiaoXXdTD0Pn46sf++K6c9Wh0TEgD6mvvQaOZDOHQBYL
1XgkitTX3lRRnfRU7yIBwZtRZe+VHa1YGlxbyGWC4/aHVJ1w7RCBy4q407jxUA+U
wQrD3GmZI01p+Fwj9yULHYBjSO+rvY93LPiWzBRb/watmpCuVOiMWaDUgdJQ1e2r
rwuTHepscUCxAHtr05mwfbxcKMHfOmO74h7zq21TgLEbxR61FDnSUCfQLUKouLKu
tWI3IWOo0v+VbBof7WPdQMjXr65AMLfXZcSAMZOy/mUY+eCLusG6Bu9EK+uDAkSp
EwWaePA6RBY5HreVVT7p1JYppojngWISo1JjsLDKDCOilRiEkLrmnH5Y6xu7vplX
0pInT5+HShG7+DybcgobbGsCIebIlwEV5v0ekGIFGCRRBywbtVpjijFOyzNOJX55
E7aKpgeoTpzs1C8+oAWS3hGHa2HasPee8F4gn0SCOda3NVOJbtujPO4U91OrNozx
04cw/Md1BmV93hZJ6HrGPwYoG6OIw4RTso1YAmhiNk6hvjCz2cBtwNH15osOQvNV
YMEj3lm52jhlt4oH4nZvhVS3XV19zfKoXxf4u18UxzvKdMA/bwnpfdhz3Nw1s1jN
cfRpcUvGQtCueQyFuqhu31BWhpyUT20NFbNsnBuaLtpFRRW9Pqk+AslFFwXmxNhO
+rSw5rAd+Yv8gRFmhziWHnUhJfrmOFzABlViM6cmBZ2+FhkeJQW/kz+pCtpf+Rx8
n+j1wlVpJjuzibBo+BtAciWQ2Z8Wx+ISvJLuw4iIpCEGZ5cbU2P/RLXBmIaftQ4v
hHikOnxAw1qQPq9xb604KoW5uuSZzK9PX8bRC42dboR8Hrp5X/mBI7c3e7k+9wuV
RCB5xWk0csO6TebRrG5zkXkqknErdkkcVLMXoTZIwCKQ/vjsvZhD82v4smAl7SR1
bRSIeliH6Y/lbFvOAtx3v9SJNZ8CmWqcTtsNaw4KpIwABbsVuuX6Am/pgoN4v6xN
GcQAomVhjMYe0Ae7qrGi3Tn3qDp7Sv4vgMiQqH9qIYT+933QxALPzDplZ+5GF4wm
EVRpyM0cwVJKhvrsoy8kAUxPmnqxRXfiHPD1D6gyHo73AteOjIAYtNHLvgnsBSfz
Z6oQ+amUFoksVHbwKER72yjoVePVJSFoyLBvYP30mGCntmr1c+e5VLbwiLybSu3G
wbV5wRF/6XbmVnmB8lBYkMgM3CuiN6KFh5d53c8eXYw7z+VMRtIxD6XzSgNgRU6V
IeL/ivTt6L8pdDodZmvUFw/6J72uGMcwT8gG5tvDu9g4UK8x+Qqz8IaSX0nugJU3
DT3ZGEPq4U9FE1HsP15VRZvhj4RCu76vwF0o85UB4t/3r5j6zLpXkgiYSIkyPa4g
/fBDA8Q+YflDelIHX2Szs85jq8K0xmvmC/Hx08g0U6M0keLeEO6+mSDhJ9E/bZbk
AS7ErJcmYHcVjhIWm3TJBLNaJLnymLLAgaqW6mBauNdYQbwHR8fzsxTEXcySxgzX
t/1cZE59hQhWPqVI4mS5fegL8I6xAJQuFm6EYUjceeCV8H39dEbqnYeuSeACb5Cw
mTJLyEmBkGA19htk1PCd+v5QuoWGWqATfpFOPiPDea17RvhZhWwjmaLzla9YLOcq
vm5oFxTViLADDSdGJGa3teJmFQf2f0TrK4cRBnxP7hZrs0dys8v1l24hMT2KvDzI
bM8SENE+B61Wfl+njFtC0K6s2AKmUZQXKm/1aVLS9zKWQK4uCV62kjjgZUX9+CHL
AqdRF4jL3jUIwFhbjKQdSugNZ9/qIURD8qEN18rOmPsDYO6ys72KtenlKk3Ei0Mt
jymvg2m/8Pgsg3JGBowyi+3hFMJxWFAbiOoDdJuQI2opEv6wHVt6sqNBQZROWm1r
AeN1eK2TNZVZlbWuRBhG1crZMEgPzXCc5arJpxXYRez7nEK/eHzADZlkP19Aeb6/
9r+E+BIbetFBHk8AtQWNFGymeU46d0QXcJy3CmbbFGL2rM+gniAQe6LRYp3V8ltW
i7X8DeoRli9vzKyDayaZyfwH1slXAbzyG4shoKHJdn99lzh/3z43GUqW7x7u4atD
uCLju+eAw5OtufWoXr9VDUrTsnZhUr4rejBpdl8fqlJTG+UzGX67oUy0IFlIUQlD
YCQzuHK+dyK6YjeNO2QK4eyxUj3rbZWge9YMqiYeVOOwnM2uWzP9zLsdLmokt1K6
QR1z2fMCjMCpnORcMYf3a/LuiUvSQ0tbtXxawZpALObMdtTkB1QvatqNnD9edmeE
8euy7QySHameCjp2J543+ID9k8WHhrdbvgytFYUGV/BWFOnpBMXzccVMVNOlVgZv
57DJ1icP9c5JtqSpMgfAWctBhGUVnJLVGlSi/fESo0trRaqPC52shM0feKeKbw80
i3EiLiQ/W6A/EVa3lXr+ADNPeC3dmVMyRNlQUd7ocFhBKhoPq4klg8sTuum2KV+8
SlVgl7eDn6ZUw6fqVNyb8/FBxj/I1SlP+MvECM5CBL//VKDIYxsiU4uOiyZbBic2
AxaS8yegg0/sFXqyN43YHgA7NftbMm91ntJyOB9KCFAc+4cZAGTkPivZ1phuooyy
T6u/7WlEUibK1LmgOudDw2AYslVyESOCGIQPO7dFWqTZDoUFV1p6AsxRn7dTdOFY
lWfvRk4jw7p8HRs0rQIZzTWAZ75OhRyPXvjvt7BPLthqbyzbNHhoHost45D0leoa
KkdXaUVUYr5M3kvB9Q0GmOl0p2gdotG0vTg2H/kXcdBKLUrsnMGWYuDntrzNgg2x
aC84E0xbQ/I8HGEuLMh4LQnTATkx0XWDeWovncKj+B2a/2nJt4flfsLWE9kFVYzE
yARnPsmq/vn8ePEFogAxFu7bYP9libdGrx+aL3ZjIgJ6WZ9wgC2XkwzQSud/7xAG
Aek+Sl5bSrgvIjI7ynD3rOrXOP9bZ7W94zms7T41qW9RTG8jiPgEisMqauXNoHJe
/zMSp24/q0v7HVWIupkHZZ5IjVBgDVQvnAvQACr9vTsWD5fBKS15gsuIG5qHLJkJ
IkhRelI080tqDsl8XJGHLb4a+xBnj3LH6FmGz3x5kVcLw7duwxcfyohkBXBjouCK
tS7RhHfvNZLdcpw9MwvPnE5nPwRt52v1JwOdHnMxyfK7BVQb7AWR+33+4Y+n+Uhz
ryiUO6Zy4AGzrEu+aLbudvjpxcR/6DFQVTToCAp+TC+Jo1dRvR/Y2pW/ZTj1dJoh
bMiHCdI753eyFWFY70n9FsnbmbmHbKdf4JLNPNQ9fSrluFp0TcT4hgMBeKO/RT9c
v2N3X7q4xX5jn99qzaqyzJrOcgWGrZJjJfisjzXwCQXtZDkqUEGeWsdYsIloOp5L
AvrucV/w2FFQXVEDUGT76pZ7rbJfKziDBeqEwH7wS19M1/LCYL6c6z5IwCi1wr60
ohIUUOMpHq/o+XsnKC+5nqrN4JONE9JhvXTGNBFladAExN/jjzaXGkdyakPvWvO5
PTASowfBTmA/SVq4RUN3UH9dHisZP1g4rZdjd4nEE2t2lNfj+CdLdtqcBYQpznVi
UE33c0pfHsUDG40grRn73VBqIW8nWWNOttU47Vl6qWYZuYJ1gmOeA7sw+SZZv0X5
sHD5wQZMtUlrSqWcS9m+pTle1i/3H7BmFD70emQW7DIA+dI8+3lR6UGhkzXctXDw
pYETLJWDRZwUN/91fMmbTgPJ4OMO0Lwapr9NvDVm/RkRtuc2YPsk9NEB5UamuUbr
T4Bm70RmNMYgYpGWB6a6NTvvHTln7SX4ijVJfqttEfxpa5N4vwX4v/B8tYAl7eFU
tuezWZpeDkgNlOzQkX/+1p/FstygX/QmFLzHTiJWZQSr5IJsNRmTnA3yR9DaE87q
mwN1VP09+KCRexqzIG4WvPZgcY2YsuZFUN/0J1ez7A/OGx1j/1lXFTu0PKg7Q2mT
cFEJag01BJL2ShPH0SB0m0W4GT+JoFxuPWpwxnrpEs6t3w2tVyDWlCPX+WabnH1u
rnfSHsN8mIdQdqgt+N/k5dDf/FKQQ3Au8oEMlR4myLbZLHe+X0QbreGhL7qMzBbl
jAI57Us96N2OnJP38V+zZ+qiwP6SXQl2CLFEkv5adjNWetv6E/uM1/rIkWQ1LQ7L
cmdTetfOlGjEvijEOTg9ah58A5jVevblJDA391pLpsFZTzM4v8hB5CULenVQvBES
xwqCOYH5KMPqX96u26eC+PbqJz8TIYV9X33SVFm1HQvImqWyhJXzesDkhqLAjr1i
uElYp44xQl4+FbnuNZlZN5IxDgW6qnRtGKDqipAtyHIyPce55FDBilx5bJRzy8Oa
xJ6YDqpqnB1ZCOdfAPtK9ZPThUbwQbpPUjVWEVvtHKgoEDiZmbq4h8SnSOv6XtIZ
/uFHOGLLkhnbhZpNRJ4L7opP3LfOFCGZS8KBKdPRbZElhb2joplED76nLCl5xCuf
OR+juCX0qiIE2W3W0urWeBYKvcDuFyyoeB1ykLBD1cgl3ba4Pj3/GTUcXRbFK+dF
qmLvU1s3E6heoFAPkBdoJRufJk071vZZxHytDNFyvND76tXSCqNRKplXu2+DtUZK
yb7Sng6KZocN8BFmk2DNXGCOFcFbuMs3e8CbNxssnem8GxskJWbbuGZDgeH6ARYd
jb1xx7h6AyJ6ohxRZkleG5MElA6w8WwV9yOlm9O/ofKmeFv7gFfUKLLziUCHkgOz
ZkpQLv5lERr4riMoHNrVAlXU0p0xpPcznlynb2B/9zSB6iT4V+6Km/7laVMMgXqe
qRWY+0w2S/Y+6OeCZPm2tidZ7TrkVowfp/WxXi9GPshb8y6LCjWtjf7d5u8thLiS
/a7zRuPySww1mK/4ZctbIHdZE/TuJi0l5ycyUSKkF8HRZ7Jfuq9TSmRowxGpr+dz
51XGX8hrMn0idzuCoiQlynqIBHYZkQRF135DXVg7Weizg8Q+IfrcM8UN2w/OPeeR
djBi8sBVbIHFiQYf9JDXNuZKEAS5MyL3yd6Gg6wMlK64ZSvs6l+eJL+yw4neBPS3
5JuP7slfMCCjGlD6a8q0q57scQshXSBRM7+kg+2MYWi3jFnaX7POXcty6GmV0pFY
rhz9HdF2yqUfGtzPsexjADaljdLOxetJmTippVc9LrOSI2abCcucaR3waoCG8cT4
qHfF1GZhQmnnH4fUEnYBpSc3s8Lsn/jf2m4nqFk5XOm2UW3jMI/ty9Wcw8PTD0Eq
9uFgc7GLkbJW5DKlUQupskHIJC1uU56/aoYXsfESA71Bqey2TsgIxk57KckhchRP
2Mmrvx0MeO7iiswgkQ++lhxFkoaGjvBbq5opLmX6nz1f5vCzfSiW88sH1aX+2qyZ
TQqqHb4i8Rajn4Dbsosh5rdKaMB0oH1vr7M9PrrjD1neQKU2fyWEa49J4arDUhjU
EFZaPpKlOvT33NQ/K4ktlE7qTAwlvOklpoB18v7UqKXBlpd2TIYdbaDDZqfBdipz
xlA356QAZfBKKoi6yapaZQp1eB1zCLhguHpUNPSv9l0/WWyXMn59G9czi6VM7/Oh
yjbfQlzF/97TTAmS8HJRoeP2ItQp82x44IU7ssC5/ymXH5iXvd/Diy2oy49EgCBd
1jow0F7XXVHf+B8cBkrEhWu6ZB+Yr5p5CdT+eZUJBqCfTruFiQhMG/arKuo8BjYW
8bnuKfevvKwmGvLwkmNlHMj9aKuZIWB6bMTDdo53FmyqwoxcdUVaQDkYxtmi0I2R
vzTQPR4rS6jxoUdfUEXXtx6g9WNzXTHL9f+66lHStB8WUrM+xQxwiLjvUDk7/kwI
Aw8lP304neZispqJtCiIL19LrItZs+h9jJWI/Z6duhJts8dQMUbXNBa7GbVVrGwH
WKidji084oRZ9oQq45889tpJ+Bcv4h//TFMN/IZm/jfGvKG4of4/H5YE+HlbbvWW
SP/mK/g4bDL9XRH3ts7dxGAf/aGaIGxCJ5XyQd3aliGEAWNvS8xMNRFpQ+OvM2iY
/rfA3kq2RtZBHkQnHLMh15HDXN6AJxbjZjHYZcrRA7hb0oR7kcnhnd2mrjw2d3Gr
Ocx7hMGCy+Mqi3eKKMN+u6wmZLa116JuIaj8fhylV3qIrduyhkuGHMzSTYZnVPMq
X+YpdIg14s4zIwJiA66V63MUSypmubWxS/5T6Ac1KubQ9P9l/O2S1ihxjETXO7XT
NRtO1VCYBKJofcLipcU/goSZc/Txzewq4tlViMXslzQnLQ+f8snVIsyGqER4J4Rm
fGLOq0K8VEip+k4MuA6SRNLiKXvu2yPDOmAYAwYNQbsNqrcLxjhq3XLmEnvQrmsu
8UPVeDxWRMkQAuU25fMB6dCE1svLHhJ7lEX9XyFCAgv+X7w0YhpzVhMIsHrNYXLo
cb7RA57IftJ/mjFqQIte5+x4e4/Z0WAkhTYGuV5W+64OIAfWEBG6FzqWrxhD0q1O
1ZrmQSNxp50dQGJNknbSHzkgzNai5U3LlvoHrLF6B9OCAmHj6dFEXzwyR+/lgpQl
ZUE5ciD1gqDiXx3FwKgJ2wo8BgBKwVRKyBtu6OMQmAwSs7YXMBXV5QZ4COzUvq2x
VMU8hbvvEbGTLdpQBhYJVrz2sees8V/xZVzfFWFPYd+E0UotEwGfNgm7iEKJvfme
3B/09sh9eFuYsGN/fiDUiqIwwRUUCZ1zwLvfONppJuw5+OZAc1Ofx6n3IyT6YAUt
lRswKC3KDqrUmWIV55Muaje/bBesuZYmoKBhR86rcvi0Fp+8FrXuWcpR7SrnNvDS
EKtErmeafxSHNN0j/dDRVxpvGgaSU/NkXm22/cCXwQ0bXT/9Ts//kDGXObRb6hWG
hQdVEXAsKe94xk6o5etY9/PXRK/awJgR+d/osBBLL6K/5m4FncainR0XBj7LvBNu
65oTpws+zPypbXXNVAE4SeNOAHGU3h4HS5xMBssePRca0jkGRMoaxq1VR/uVB1Sz
mTw3xDeN4fZsek7rooFEPsRGX1FBOqYW44Z03xq4MkA7bYSn3BOiy90eJSgIDNW0
Cu/cXg6w/4RPXJxJdJdUdmTQOw8a2FIsJ+Dssjf1/6cGIIC7iFGSw3hQOheBUWlE
W7tnhs+iRL3Yo3UdKKVSn25Jfh2RkAojFbos4IppJmzwlYPxnVQwrmcPmuSHaSdW
W+UGz11aeNS6Nm7XWzz4wXoxHzeplKhw/Tgy/tnDud306TTCPxJzppNJM6ugOpeX
kzbm6XP2aQZ39lkMm0Qo+A1ydYaozSn6u5LVlV+ILi/V0czLo7j2nakhcEdvkZE6
bP5BC1MXmRr7AKIxBsvz7L1pJyGf8seyInoZWdB7XWzQqhuXJU811205VhRmU3R1
GqgLx10tfnmuItLHp3vxeFijXpbYHeoBCVIHgLLf6KAQlWD2fNAG08oUr/rzdylg
l37L793Q7WOn4BX6luclluZk8mPnVxFyOftxwu3VUemsjkZTPQtOfSHZT5g2Q0aC
OasRuRCDd5khjJaHPLTnnRBqSUBgmohWR2H1QMbAQZiNn/9gzTMCXHggLC2s7JeL
EA5DgsklF1G5KXw1iUnxp9ajH/wzwaQUmuBNTNcR2QPpQxAZnpUKNrYrT39u/ro5
i7yJhKvhXsmE9JjIljT/q3s27Q8wlxUjr15rODRyBhbXlImk+kSbumb01x+qCs65
QgYYdqgIRWU+5Q9YgwEdGgs0Z0OPQFmXy+h7A7VuTmuSsoBIpTPtVQOxYfdJaRZz
/azTqcAI3hzeTNAxTb5/o4jJp4gqlqcfOCBYr/Av+Csk6E2zDJy7pe77PCb3SRHD
CSTHHk+ZAM3511fRGtZUu5lD42tCr8ro3BurbFTgvSw4Ne8MBchE0EBZ2RzbNmwU
11q76Vgp1oFPemkoeeRMI8+G89rFcW2S6/RtoByqAiF6gV/rW+8UGPb5SMoXXiC2
6Uy0UNVGhGqyp3aX0gudMpoZOKKctksy0n2BEXyZvhrR8z7WXGK8diFr6TPDYoZ5
gRHPOhoQSDVj7+sTdfTy7eVqyLuW4cvXLggV6f4F2sAO6DO7JdaamP5wORNGTspw
IZsKPXNIg29/OvOxRHUVQCGsR9MSimCCLDJfylDi2CDkdWcG21tvrC3bBrgLRXa/
LzD7EPELZB5tSTJiqbdyXVS9d0tTWVsWeFixLzjuM5wskNzfxm0G37dbGB7ixRFD
0jUVl9WuHsH7m8o3wqPnV+dGi/Jl4MucX824oHMPXZpyMiJHeeVejrDp03CVMvSy
brVsZtQolGxSfSE2YfX4liKzCi8Xr90jESp0NMMAgWFgJzpClSSXMvR8fVjuyylv
+A7+iBf5GdgOHBhXOd2OPid7NO1xf9yZ2YEM68ttXJE9WYaWLZdHpi7iffHwaIlg
FFtGNYR5zI7ISbYbhbPmoywi71v+J6ITqilei+xCaxaeflC8gF8wIVh0EdL7JM1j
mHA7i43XniSVgjXYXZeVEy1BILhvv+TyrPwiqi+gPznxEdUMxGe2gFriYAsLXucS
18VACqzxf0pZZJUuFMs2islsUn5M1Q1KFNL9D6Ogyg2+ybiXxQxhR8qXBxcL/7/O
FDcJdZCQNzx0VJamQDUmdMy5T3p/Tm2XnMf0RMAR+42FFJyD2/oeKlbhuI1CDxvw
sLAktXS51yrpUgBlZHuBuDcQb/vxyrp5i6VwHBxLppg0x1gj5DYcJW8RtMopPZfg
kYOWzvcw6kq21SvoopDTQdr+f5jeufuGFDRN3PlOEKt2L8AhQKeO97WCxCmYsjyr
h5Fu19Vl2/igmdpPh3Z7vzKUicTa5gqRgQrfBxAZN5noFj+mcUrY74AzbXDRaV4L
lWJRHaYlz8Kn9mo6qJoZKL9w2PpawQeGiDU2TDbRYEa/p1TqJsN64VqTA9dCTRJJ
/3BBkquY4i9mpa3XCJrsFUzGdG2VU7KJfkV4Ey46CCHOQTyvglFx/a44iplK8q0C
aq6CHdiErlx66V2V+MyaqRniWw5kd369AyOC1buWqdjLokhVrHx+EDqHM4ZjEazq
8ZXqGaIIbPwsN9ETTxWeRnimurCswbBiWFZOxcQHEdWx4ItdQ3jcGWNnXC5a61SC
iYOQQ/vo0KWvGVAGhHvNeaFicidh9Bwb0kZ8A9/RB2Rg9Nj1g/OiVglUNCFt0C6+
ER47J5ZjyRF87cmpQZLVvwXmOLK5rmFfOAPvnM7GFkDfWn/lS37X4SyZmTj1t7vD
+2HLrXTTcKBufioXerCgdGLDxM6jR00SJVNIffXqMYEC22X+kHPk+wdGhRt3SKpQ
vVmgfxiY58/SyFt8ih3FTPQIzZTS7IIIny8LQOstBVBDtNMCsASodtLsveFi21T0
kE6EhBWS+qgH40DQXoncFSFm/avGrPFkhN0Sx7wj/CUo+1yyqzMfj4rDvRvI7M4H
/jjyxfV1F6cdKD/1H123jDl6+1yKlu0tQuI1Sw+6Nd6uMdRlD2GGaYb52MvRVRmW
zxQhYlQGW+XXeeauqTDko6QMylASBHc17p03WtA7HasmMEwjCtrXiQNgKcBWWtoV
TziJ2YLKJ/VHK7EE5A5GAGZu6wj13DAUEvVjFlpVMczWtmHsW1pk9hxxkONEmZuE
TT+9p7cucaWz8BiWgJYhICpAHf3RLAirdm1t0n8vkmB6ikOliUjYNM85JKhYfZjU
hfvlPsKBzp9zqDC+72jc+cn2edH680/fRJOAlRq7L18DBca8ViY70HcVRs4QhFLX
cW6LuWICt4hIZb/5tuJhv2wZW8JZ+7XrMGmonewIKGi4TuqPUPvp9CnNPmo65Jlj
Xm0tJgyVIcjPaIwF30h366fz6unrO3vtPyczZM7QwtXVQH2jQdaegxHDtOe0eXZH
v7O/9ZUzwaKDjJ2r2o4JHJs0ow8OLgcxzZq/TH+PdtUl89bTvLWZM845VyFeKoSl
hBwlN3WEZaVD1M1j5htEES48DE9Ku23i530Wu/l15mc/pipAHtfyjXPwFVUz/AcU
pzYtW0HGBFbmuLZ4qNNPgk1FFsPcKkXh7j8U2bnb/+b1Iafrkpvyaa7p/ORraUze
vJsvBH+7Ch+HOpizMv7yP9AM94ODsFREiK+T1kX3raI9tM1njrMrZOZeQkhRBiWV
jldTa+hB8jRTvBEkjEuXMb7gVhLZPT/GQF5S3FwG5gQ1jpjvi8BKripRkKWuAQ7P
kYb53+ujW7w/tWH5MrFqDEd+nMct9PUEZLChdUqqotGJ8piVLBf/jETFN7Dxb8xp
eVAqiM1ZX0DvRGe/hArjom02Nju1bX9SuMcLpbqp3jOvKskj9g7z4xIizt3t6Ku4
8weRDiHYRpKg87O+eU4TZlETNCekOoNCh9dA1ywI27MiT0QTTUwUCERLc/T3Q5s4
emlKTOpMrh5l/cbeE4eTUi/B+CynMEqWN1905X6vPVlbhJyO/XxMYSXasqOEXbt1
WIW3sXfayWRRshrRaZaiAld2UGRiHWsqZFfIB9pLgfr5Lp8Xqs1c+DoOOvwAdwYr
rmfW7neTSz/kUTU04QNcIS8QziGfQfhOnLWvo+y8KnA/iB5h+GhcM41VQ9YkODUF
qQ9qaBHNCwzWLE9Qb/WGAyuFXZ5vwaTvPwhWk3g2dHAvBMeogDE8arsdsNphwxig
7HrA/v9IMaRUe8mATiRkj4cLMoeaYvD7jP1Nk/gve+5zegsXkJ8u1jp73NM+8rB+
lFCQcQakbOwp8OMAKV92ADKC40Ef2td+ztT+SVxLW2HMrSGK8x8OdzJPg2QZNo+H
XKZCPDNucsburbIjFdYwG6uLrKVepx0piVccPSwrG2FnSzR3lIQvi4lTL0tfkhWt
GaD7cAE21S6U087t0umchxoIS1vjjbSM8bPdlqDl+HRYTw9Xx3hDVJblo1xDlWg6
0h3k0xCP2KaH189beqPH6hIv1Qs+dbXurWS/RmWaHPpXbqKcF2dDoUInAESBD2yB
ZT4OzTKQp5Cz072HbwhCYbi71qkI7hWi5i10z6Vie09gjxef23t66eLJa/5nSvsj
V7Xr3TFJNKGGB0sAk0IkLeLwpf4MqdJOUJQD7bdcXKfWvXATtb1AK0eZEvdednYG
OJmXkQwqIKcJOlTt+yFKyuM2rOedz6ItNm+v2OTIHrIdtkBrg7jVMkmy/1s9uRJO
ezn6U3q+t2eBszM1BCfh83y61QAh3tiJm5p0JIaIleGI7cAjyoGnN2jyg6fE8oJC
HD2cw1JFnAz1YxKdBYQQnf1JXetHStXB1Gt1E3B4Wfi0p0SKyxMegwKysIeaAsv9
L3JEEvy1WXbl/9VnQCkNZg0YeKEBV9w87Yk30dTAyLCFhXfToFiJNB+ZP1O+UYIC
I/HZrrXifBOO6mj35aKWQ7wdvSqZgtmelR2y1VnjJ4nDUEs8BpAFZ/OhISLVDV7h
w2f53LakLm3OkcNtldCdGdpySmx7apTkqSeqpWs2q9IkobbiaKEFYMEdgoJsviY7
326kCjVqTINXYfSel9NSAsR0rV5xe2XdUHTI+dXhiJMFnMvj4/oT+cpSvydZZhwS
gwbBvScYczrXBLDV+T8pMNX54fy9wUTEVqtjRBL43sxiDFqqD10oNJht/UDcbatk
fzQU3FEmyuXoWYlOe2PI9y6Znf4CC/PRh8tO4xn1NZSaXB6XHRitG0a/2JCERjqV
8MauU4NfPM9S968NAn36rSBqfOxUZD+h+8v88Dk6thfNdqkR8JjDn1ktv8var84p
x5rNmUx16P991vfLxnlSUb+k/WsJCSRKHSvaf1ZP4nvyW1MnbP85uBrkd4IMa3Uj
ysvDqmC6ikLZtdc32pul7xUMn+3e5jCweAQFvCcbji6ChCzRpO161rPibN73iiOu
XF7NyHGRMNVH6uZSmqGiaL81G/DBBB0p2qr1z8Aq6G72F4G4jY4Zy9dn2RfwCS38
Be7GtvrKc0Ezty/f4GKqUnLVFG4CgEjLWqtiA5I8/eZ94DdiOrjhQ4HALllvjBFY
WsqqlqYeB8QG0qit709f0W4P+kq4hovgqm7Bv3P2sX9STOz15gytzdnYZd16YLdE
H0bEIjznZ9j5AE4opDjD5angSoXK0BW7LRLeZRB3N5EUXfjvKUbINYpPYL1LmYYV
347HHzRryj8zsvaw60Cg/2EctJ16CfT6Z9Sl3TrDxWbYod9jxO6W+9Jk/soDYCuG
UAhXFou+yv8N5OKFLZ476UEa7ukxr9hfm+R4JwarlOvZTdYkQicb5ymlP0/7hJzi
dBDRe3ICvWKMSH4n1evvnJWHImtteiU6NaLkyrJS2nE+8aFcXaxxsjv9MVeMGKbP
1jdikVH1HZ8l+G+YvZrKOxUaXwA9Msqgxhzg6oCadkD1tASxdm7Tsri6MZ8xiShd
uylaPjs6+wW1FaJcd7aWL3QeK8v2d+LwqhQl6LDYWJfxmIjGIJfQ5tWzgl/hDqqK
Lvt2ZkT4o5oXbjzIu41Ll87Jb+WrgcVBXwHJ3VV9eP4ol6BPFd9BdMLzbzyzuaHA
`protect END_PROTECTED
