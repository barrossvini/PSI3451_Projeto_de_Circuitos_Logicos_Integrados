`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N1HOD2P7RkKwYYow1XHVNfZhrLpbZULULW97c3qkXTfujHQW6fpdTKwZodcgGKpV
OzI/VnyVn50lx2S/t6VB58Uu2t2PAHaRoj1O9B81YdubZp70RSqflgoCfstmGmIH
WAuasP5PAC4yhyOcE7cr6D8nmgAagmtrFYoh88xbfQLDf0hSJTlYZz7K4gnQcGn0
bPOLv24pA/Fk+lbGI3ptdYHVzzKxgrnwMRO6h+01gU64TmyzP9hda8KBauxpr+q5
zQiKvPsqvxE+I7bDHyuSJkT5qxUm/8FSHt/aQCpTRix5ZqbcdK3hBMKpxqjwc0lV
R64cqIRTg+7BJv/tukEQD20YH+2/kxNJNe1U0UWTkjFnE4DpwZuqxq8k9d5JRgrc
EgT/kd9o5T3fBq0gUIMinEXG3E2kG7upLLA+li+Co4ZdwdPaK7smK37NJ932pWqT
t8omFO5HDQOwnTcwOyhLLfcGaQL/MhadBANJLvO78OXRvV7fZMGUkGC396MT5Vaj
jDZpKILtmENk+59a+lEm3sHmE1u0OkyhfOrHkWXe1nBwZKZSYYLXnt0fYvb34qTV
OsTHqHbni/jNRJfBi4aXCzutFKa64eFk6NiC+Swd1rRIT4W1lsTSk8MJPMriDI8G
6G/k8F2uRHgG3xjAOk+Z0cb00MK1tFVPFCLZGKQD7YxjYZZWviDgvZxFnd4ga3sC
TQlSk3R02d2IQ963gPsW4f1Rcmo2Am8hdOUijXyagsgbEHV3Cs6xGBbBNQ4qDk/8
Sl0XXsJFJvCjtDR6kevWirdoB9i/THebtPB5DDwPaq3/VyYZnqsH7B0jBbxAoOcO
iR+fi5b3MG+zLhOERa1LurzrZKcWMHcualTYbRAwYAYDJtfbC1vS6FxMGQr6xcvo
mD1MGDh8AbNJdwfTn8Utx2MDQwgYrHC0peRQtuG/e5vYFw2PUHh/IGwfna9fSjms
pwdvVAGuvn+yuIfO56ZDFF19Q+SRW8jMNFvijKdCB6XM0yXtr/U2YVQwNPq7kdzD
jo66mIWLRZb3JJqxFbuQc4aq4F8xgOR94jCYaVm8mMNWeWXkerVFyQrbT4tvitlv
`protect END_PROTECTED
