`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DhlIbq8lgmUCupV7ywRiU5gHOYVsceWCZ8c4bjdPZyZBSzknm6L5Jpikoo5R/7Df
roj90v4VPpN+XN5UKpEaJiHS9bD8qCBpP3UpJyd8G/K9lJjI88r05/G9XdqnN2eb
pZ7kRK4tUo8nGYRplL/CSnEl/TxlP9P1zZlbeIzj4VFeTxOnzjzP0uBIb35ZFWSL
RuaKTAEM5JOcwHZON6NuV7ddu0Qz1cRKJIiAgWP3EsiRf/7Iw8ytARYUnXWwul1j
CThCbBCROBDr3U+rYb1LtPe+YSjv3zure9U/kWzyo83NL1OvXzupFtpIDmjhBcMK
OQwdVPq5EM0Xs37MfytOer68XGfNETDhagh0lQkxhz3StYB0HY9E+m+KjpSqQJOC
OB/Gmn+XhkANFDPluCe7e7Pkw+VaqxB40Dd4yWcfMP/h0wfDDLbyE51LV59Yyide
suZZyhkaqUFuji45JKTlD/CNzPysMY9HirJTjlTK+u2afvWvmXkaBAumKLAbtjfr
4Yh7/JjGhqH6aMU1rxkDzw==
`protect END_PROTECTED
