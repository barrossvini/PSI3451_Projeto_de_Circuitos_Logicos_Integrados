`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V9IA6noNKiUUDZrKrR5lafKuU5IR13u/9zrjAhrKS7AOFKd3jtDqPglkj8tRpz4V
5XbZvhWz5rRErfUIt/+6UJRA1RB3Blw82u4ZtoEMc0ncp5gDY3ur+qOuyf7zqrR2
yblo5BlEO8P4N4R3BhBipkNEFW/MPVOmlBUmLTaCTk5Xzl5cipnHhtG5cEp3CUmp
KFLHnaNXZLPeajQ01yWCzl6zQLeTxX8mRW6tX+CmJShitANe4s2oM8VblK2SnkSN
B7ck8JHqcCFwnroyhuCOi2zSWzU2NNAB7zimS806a4jGLxULGqhf2MDs232IebKV
GAun1Lj6KIYqwrItcfnMjZLLjG0hkXvjxWL4a2G2QntnTLBOE5GmvbpEAEMwcnnw
3+XissP8uW5wm053tOIDzPBsHc1/0y1+K4Iy5CdWqLFRMLi9vMCmvwKzpDMPEmx0
mf+7DMQYwWCVpS+qDrEVdV/jogFF9RFpIbuI4pHEmknhNVSBwmbgHhehAHd2/4iH
JJiDoeSmc9sDC76kcgxWuNP/dEh+fuVkzIVVLB7ETXZMiV6kiQgp6aKzHeWBIVJt
qe+ZKTmmFvc5kxC64ntdhfsFv/QYUtLttAYSz7JGJvNU01VEhn/wFHBx4n5Yisi2
RUMV1xINF4u6eRIMZ246UizXutRLNU/u7YB5TdPlbpPHfLlC7H0kPbKylI6kuDZn
I7xVyU90SEM1j7k+IjZZJPbPJwkUSUKWaxBTK5TnwvFokFKMS7mMn95JEYD1GUaT
cCnhs6MJSa1Yrzsx6uVcDwoImRacpZc4A5Q5HEaaN3UGouNXV8PBEhePNPqaA4VW
gTPUAnK6w56MJYZlOpxJEgo1knKtxwp+ivYDza7igZe7PdMDxdOjf82+iIJeousK
AlpEceojl+Gx1JgH5FHBMYxIRvAwvnaNk49tDKcfz8Hm9XsAgfbxxJv246meNPSz
fIf2DnZfDesO+9W7TOnnZAHwVRUioZGY2nVQr1ZhGxkfmWJOPbIif3OebJ/vJaxX
pTihfxgfkCXApBecvQO8HxlKDvcufFpb6aG/GMZs39W1tyQKshhUSK18oeoG7dSe
8ZWSWJKuTt67hMaYF25TfzmMR7UQZ9c4j5Gw5tw+xWkrmhqWsJAtI+q8PoMJYUWr
CZL4T+zlw6GnVCz1Yuylsxh/pjfaKxS54va9BPeuPECLLjb4bQop4ZSvpBzRQMHA
WLaUscXlYZhs9NSjqJE/tdyM/AC2B4gNy9BJ/zBvaYnAN/kBpKBWNhGFk9TBTTWq
zZzrKzWKWBl9p0mQ+JAmPY5ul2WVskl8jzotkqBnj5FQXg0M/KFpT/8JGQsD+Rwh
cUstXb6WObwkOelk6OHwTwo+Wl2wov0sb8qkyiKw0Ca84zFMTn8gvbWQFoaqagTi
TEMqsYKBVqL/djA/PRqdRoU/o2PSPzvtEKLgLUHTxDcs0KAJvtmkh71D+FPr6OdZ
gwLCAgDkSH4ENnsxuS6hVLOTgooCMpPIkw01GJCfU3OJL8yutXXJ5qX6Cvoo1Px8
mf0cITUdZ2ZjgoLcF7vtA04uCQ+HHlC/oXDYrEI2M1Q39Eg+OSoh1tU4xaDyXYNB
JzlMaOY9H4XoBEVFKj8pg7k3Bq6vrffSRzdL/lkb6fg5PxaxSmPsMshf9RQEguEL
hHTuPV8g+aFd+Sc/l09nX/aLeJ6niA0HTDNDKdIrsMbYcqCPVpRfiplKxYtd/xIu
37B0UXDJ5xtqS0utboVb8mdvauGlafLLrjDgb298Jw6JCV8OHu2a+lvf0vaCgQkG
D9LcS7uO1KqG5/1fFDeFFKukiVT4WDznqqsyvGMPYHTJirexbDxKoSVAvJiEjdcy
CFhOMyHpznnH7Nl4/gX+1qUgWpvVWNqZomWA5LC70DSuMDDTzCFrjN7PVhFseh8C
czQE0YdXF7IkBJx44zri55olGo3gFOc++NulVtYxrZgrv4QUvGxGzkiptUd41pl1
0eLwrBvj/EQl1VLE0Q964lQ3uFYSInAqJn/QM7GmHH3gQ2SvlC1q7W4rLPv2gPP0
ZahHJ6wSnQfUtPBQ09uDBMuikXQ/OkpmuyCb/J/a7OW48qQ/zNrtKJYltHMeuHvk
sdCqm2XHVMaDLye7uw6zgHSVoLKqMQM90+uBLOnZW8A96a3f6EOQBxmTy3c4mSeM
QzLlqdBp9QBzzbizMU3m8caA5C/ZF8khV/NuNY7DBOahlDf/Yg9Nk16QUXv5Cdpd
wNxWih+WW7OFCKL88OaytLLJdNOJR+T/PaR4VlZlLKpg+e5mqi8GL93Gfct2Iy1f
Of++i2NBEwBoJN6cb4KuE85sIP3mCZ3g50z9WNPM7+CmQjar2NsG5yON7TghSmH3
ahsiiR4ouZnzHu0sF+rJdv5Tld5yVOlLlyOehQWTNcQAvMXUVNIN3sx5P/Y5/8Wb
PVSaxlHxmye9ARFdAR3WX8YcOA/HQ2aswpufTi94uoFMWmPvqQXkEUIM/tF7sQI/
7nWxJW0FWvcTYd6tYx/Q7fM0keFGF68PjlLMY9DuVrO1ahdmBwmhTYSGHRBVScXV
E/0G3hSjaxWGlYngCeG0oOa92Un0Uzg4lO4/N1ZgAfbSi2p3xEzFybvsokbKeofg
HriSmJOBkhS5Ka9IbehX5IBFkSxtWCvtXvfRHdAVawvHOadyKh5wpOuKHkFWzttm
/buoFGvfV/VQn0Ez4asPQWJ7NWEG6yUnDmpPpLYzkPZ66VEnGE2jLzhhmOLPtvqn
7Eb2tayU62EEMVXshReMVnU325JTiVJS9IQ+qY88qkKyaVtIaVvx8YQwFdHOc18j
zmrLA7AY3gVGGw9YS/6G/Kbbla6viOPyB/ewoQMeKAvLhPW1qM4FnjvLyYH34BN1
w5kiuWJwdCFYsbmROYk7qDXYyYMuCekiZb4c0ifUwYIIsxiTYWdf60DIKtltJoqX
S4MiEJ1zddRlB0nENdlW8pHiMpy6UA2VZlXJjxSquhSJsfKLj2QB0mUTPcS0D3Xy
4QOzWiA18HR+kfgQsEOQqZAHJlZ+/yFYB3dNKik8lg8TxJpmveFpLOpvDDKlsn9a
YSW6vMWFVSB7+CeO6/ungfvKW/c0MTnoM8TwQn+CRUjlUvLUIMv4j82w6OFQBesG
bSst1mfsQ6vRjGCqMloLMXMZ/n2i5wJjeHgl7Ot6+J0PTrhdtzjxD3qb10Unff1y
tomt33oEvBFL1IRuk+f/oZLvI7WV2Gb6WsuIjqLMLADHSOAyTGkWKuXYpWxzo68+
Vru3cPAscxXaFQXDXQEGTERg59Envvb7L4C0VmwDx2dg4Cz8Src83gkumlD8TwoK
lQO10XS9TjbdZBcw9oBw9OPY/qYdjwCM8HN6tuF4hmGqbGt3gwKO+Xilalv8mpnV
Nx2i2d27ap4TDiyJ3fODFIT8QsX8XcEwAg3UfWPY6HKKn1tLP4BLrf/ebhzN+df1
Zc2jpXx54Kw5qJL7xsBkgKO9xUFQ39bIgVFHtMRpI/tNqF0KpFQIsrPeI5tVM/mH
Ognedz1MfYejqOgxm8hdgn09gsMMKMTphXEedXjKxH9sqU+a55wxMQ2G+DjxiqhC
RmJfXmGPn7okMuhrQGdxrlmpd0aY43OXIuY7KFnuRhn7Oo3m9dEd2iC+86K6Cejk
VtTmIJXR0ipkdgDx0bni9L5dq8cvM5leIk+hD7hlXv7zsg3irLWeeG8N++JHF5m5
1cMFh9Jgm073J1bsf4zSXmxRnuTFu8zIvB9hF5L4VSPIbAEhVSq0BX7/uNWbnBwH
D/lK0BrTMzKYcX6WXg1u+DAvFSCBTae1htgacbNLfbC/nM/C5LwzMf1mKEtvVqKy
Tj55sUyK0gq7e9q1YwCVxITzl9LSjXu0bBQeDL/v20W5aCN3j+XKKV8n+9f+LHIB
HEmL7KaJvgz2rEaZplegrG6C3TGS1oeYyzJ32LC1PipIXh6MAuxbg0I5D0lycpuI
/g+LFGJOey6wmqzN/IheFoiyUWRkjJyT3rjtHGaCR+8=
`protect END_PROTECTED
