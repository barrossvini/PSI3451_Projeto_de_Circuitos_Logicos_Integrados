`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iw+F8CmW532qJuHIiKx9mXhnSx89KVuKMW1DEdg+7CoBwKSwdvzo0psjxfTEabqm
i9OwnoaoOvpGh4YMK76X938YJgU60MAm5X1sRJ1+9atFFTwmI6YyX//RfsLVM9wT
/VJyMsq/bw8t5cPb8nu9PJbdUXqjS7s27O9TawY9uXLbmJ50CLgRbxIaKW2cWFNv
gouAJSHLNy+iAHl9N40PsVpuDLXBYqx+b7e/8ddIXWKhdZ9Gd6wPInKn9CWaqFPQ
h83Bw/Eerrs4dB5yZsRbO41mcfQ4psSgjv+AZnMB15huDsv/UvC+Ks6RKQ3h4v9d
oIeJNAeFkl6omK3vxxGdtqJaIiWTVTeGLVPLmZXcY3e+ul1z/mD7dDsNwnFuCbBR
Gzg3Qhvk1TQFBPekQHSwPkc1cPPQTaspQlgHBgr2od383n06ZAj+RlPPNUCdmaDi
kFGkk5v3d2vFSDKiKu6LWR2GulItSic+U9icIAqD7jXxSsKEgD5Hn/fSz/ZBADhy
5GfJwwNigfPqFUXI3tVSXBbGJZ6WV5zpc553WVN6ILlbTGlPYs8LjVz0G6Ep3EPe
6dk2JT92GLdmHNp5WzCakZT7qYPgA2S6pWaeHzJm5pWedtSRN7rd41+MYa5cB1ig
+rD8i4elgIw1W9+Onsfk9E8jO7W157MMG9NvY0+bFut0yaYoyIV+vwsWvWSKQz67
EstRWNJh/UAxL82K7DeSSmL57X+Ji3hsHwfR82ehEAk=
`protect END_PROTECTED
