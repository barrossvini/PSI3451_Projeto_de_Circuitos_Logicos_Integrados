`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xWb7Drnir7qkbkZICtrVlVT3WWrokLWXUGVG+VVBfiT6QYFb48v2MmLB6K07efTl
KOkF+c4AZ7O88muBb1E6AM7vq3ZLPhWQ6FAfSK3DT1h6zukqYtlpBIKlGxw0KH4l
wxZ9mbIHuklbOsxWTHZuT4dvysTKOACRKp7FzXCwMD1SpRnFIaj1FgGucswDMe3k
DYXYrdclRBLW4E2Dz3iMqJr2DmarMp8LrQ5feJQNO0bgcIemLRhynqHsmFlB/Sch
dBYG+mbtyZ+IKwI6JJmovBpsCzBAUhI35AWtK0VIRO0huJ0+x6FXFpOc/1p8DQYu
VaLofbaV4zE5pkGJDP+asiocqj5Vk5NrKLMtOL451nq4uTSL9yCbC0PXPU2/Q5qc
tH3vegrUyKGoroxRMiYzrdEop2fegJi6IVjk+RHk4U/9BdRk4v+lFErWcJv9BVF6
+BoP5DHHbO66BayytnSyd4hTzrJz81CM8wfKiNx0lUHQWBiz0w0pO7ghWwstSCLD
63f7KcNshDqXg2b7GF03BVgvafzrK56IxkjT+pDRqCjloK9sw+Lknq69mdbBMo7i
eYRZsj9V866+KYRw/fRYJEzdDsGaAsUjh5h3k81bwMJU53Rm1vVekFeAZxFGG3qH
n9if0Hgh67tWLnO+AAyK4O6PxY2qugO+R0r5EaEnvftn35E/PlW7GcOgLXXLweXi
qkl6kb8ksIn48+CtgMQ++g==
`protect END_PROTECTED
