`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FrasLNrDnh5XWWQ+gpoB0WKURUjYQz8pKnl1gCgNHx2o30oDQt98C4jsu0PaL9Ul
bOFdhgji0HqM/FE8BBKMkYEzxCT7WhgsnZb5q9HaATG6qDflPtj80jll3MkZNbhD
HhGnPRicpR4QEmK3ZdaW9Ms41H/ijEYV4WxSgRxgCadQm+gq7JyP+jPn6fQQcact
p5PmUn9y2nzQiKtNvQ55gc6sENaZ60Xu+F0mGEBSp4RPVIDQGMWBW6Oor2rwIVmR
4q61jFgVQ5RLjNNUNZxwyKzArNkROgp6nB9LUTBqogT3x1VdjWtm0glUhHgYQla2
nzEhbXN8QUHRRVmvNwA6of6dXL8U9hP2NCOUbC37xETIW+n8CNkn5NNZxMTjDo69
FYP1GK8AQUMhc9J5Bs3D+aqm5X5EG1BfeKHerP1xpzHhuSUgXRpBnwoBXaqLb99b
ExKjniHQRZl8Mvw9Q46qeR17cVHL+eAnrMFGXS/HuZ6m4jBgK1YswUyt7Fm2RURn
OgjYUx+oxK3/IL3w9BQopyC+2TzDHC/Bil8OrChego8d5NwOzlTEyq6Y5ndmYyZt
P21bgMLPqWGs+lMcALKPyr4P0UasByriwwGMaWqEBkPrJTsGydjds2NVFbjDXqbk
LoLQjyBpSy9DseQTxo1Ka+GlSnxDbMoFEw84P2HMXAJOYJySjCxgI8FhiK7mYdEf
YuKVx4HZJIKORBVY69cYm4x6RjhSNBbq84XidOexDKm2PfmEPcDz0uSLwb+b11K3
Utnaoz+shQ1rjd7FwY1AK2cF+CFDoHcx8D3tq7ep960JuDM56Gtm9Tkr/daizngL
Inpuv/z/1WGdKHo2xk6FiIYqNcGHUmeIMKGZDXiuUGmQsumqRwDLWKFwfuH2sH6x
9nrkX/u1jrBV9LY8vKEwgZVWHTbwGepvOuCe2r6k0IQTrHphKVD8RixoKta7YTJE
BQgOqBwY6wlVMyKToM5oglRPGPc/5sM0UE0hEKM1k5NL1OTv1TLL7e/PLDi3DXUy
AOqcAdWwC7K+B4T2XvZmupGB87SofQtc7zq1C7FnvTpDKzY12a9SYWQpuIHg09t6
gYypYV0G8cuAQGwr1/97xWewsBECGC6uranUFut1fgRwRJ58N/3ku6fq6KGjOi/x
VuXFkpchHslzsj1TbYJ0kpuKD707xJtVpX501JfoOSuBNcosZ6m+1E/+eGlWlMj0
nHVeUT61Nrxd0vl3XIj3G6kd+DAY+juwlpbVGNjPfSKvdq4Vcfz7YZE6+5HMkYHg
ogGxPveWbVvl2p1faL6o7WqaWN1o0YEZTJMJIPURCLMQGAxsW6oQkpdLDHxzXNAC
pjUMPkcZQcrb2Sb/UPg4KiPPNLaswkSrejkbLEw5Eq0WFOhW7sNKub5WKZHFzUtM
o64whlWeyuihidYemaK+eA==
`protect END_PROTECTED
