`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MKgqz1vXhB+5zPHN/W7y2OAd/pxauUx/Lm8iJR6CJvzY6ionZ2VNeDBZ73YoKH50
KgNp0Ql6IBQHmXnwkXhYrPHWK0c0+ZvLEAe1e/Mpu3ixn8HykKkfD6dsWWRaO03I
PbbuyJUzjXv7fnxdvYFWU7GBxXtkF/V+H+Er4eoHp+1z/++MqpOtcuvwHqx84zhw
gcyxToRhImUPgxnIR6+qq7tZVUYthYiOhVfo+ftfVlq+/SAzIUT/WWNGFgVuK8mo
aHJhafVfxipVWt2QAkNzKFwx4ljziUuenfMiq6r+ztDv6pzqKuPdrlOumCBERQV+
GFbjNaK3uyG61Ncav8ZZyTFtfdAVEKXhANtWraelUzZSHIjGS9E8osKrtzNZC1Bt
thd/1dS1KLNq7OxgHpB6GxTd2c/Fv4SMVq/2Um6Zv3rklfD0dO2KO88B9nURsJKz
J7ZrfleqZEO9avSk2gXd5suTWs3ILVNtBiEOI0OydGr4p8c7TF3y3a91sfB2A75h
tD5xseyt8EklXfNYJCF0qbY1z4aDslWuKph7eavUB47Wb5hABBKdL1D4gSFFbNkU
nBGhUZznENWm4xrphWTK7gy5vO8onZpQNQO/smCXxQXxHwhsQ1HiuiQlhgeXP7KH
bmfVw5jvJy8LgcplstCwgD14pqRl4f2YpNjDgH0ifLOCKlIVvdtuFN7ZqsmmWpUs
b7+gU8SUitk4MshiKMjRIS92K8D91K/ULFY2lXCikJvYDERzQoveZuU5NRI9K1lm
9I8/53J8Ngfl4X4vYBdwWy5Ap/wxeFU1Px2IA6vProJxRNdBUpwM6jtoVfMPZW+k
FUFEtCy4PeyxCBzCQLQ+PL2MmNb4UucRopicGIoOlifIewQTrDlAZDrXWEdqoZQq
TEJcIFaLJV0/HJiANiMwqIaG4VEZanrDlrzCKsPrM9Ihp4EWr4d0FcNDSxJqY5Kr
h4jbF3sw37k80R01vxpVa8usTAp98ViP7CydVM15GiUuagU3KPYe2yVwlAigcH+G
qDW5YiPHuh7CKTqGn0LmJ7yEGczO0z+2/pSY3y1pULQz/RY7zf2VvdiFGTSaW9e3
VbAeaHx/cEeNfWk9ohh2cRKIp1UnzQP2BTPiQYaAK0mCE6CjFXEg7ATXnnPckgrE
61/7tgiNQByJ78In3vVHpGekSNkxK8VOnkmbHv6yFhDqAp07G/XQg/Nc/znf7MY3
AFmO9qKwfR+wP3LOnZj4LukCopPaN0Sm1IxXbftm801jKNtu8QaPa/wCzaW+iDsb
0rPKtIjoOKuSBo5SF3WmV7tMgEJw9Qk9JQVHhB6vq+6XNdA33ykg5bHz8rAld5hZ
6NMB98LD2UfjgZ0QnfT/BCgMMmj0SCuhxyiDMDREfi+Du1scyT+AP5SR+dgAsnfb
/JB+C9hT/shUkbPgoRBjhjkKcHJgC855fT7tTQBUTkI+yNVjH9UYHof7XCVsTssT
lx9i39rLgpo5XpCZJRE9Cpa6vAtAMCLGDWMd8bvloF6zGzItdIDf6ZA+fhPDNG1f
3JcqjmCh6OCZypswbsuJgQMAkKv6h39e+9YpYIGyYeMxsORBB6nl4MXgtR2XHlCs
kz36Mo7+2YsMF3/KvaTRp1Rvmw1NEolPiXmAGRn26QSvbjqaaoLjviWDoaDrO1AU
wsGZvX1TN5f391QLGLF8Tg==
`protect END_PROTECTED
