`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
057f+/BDEEP4ebhVsbOw3d43tR72dGCmEeL77174309whg1FfCtzZl4EAWyKQrdT
arEix0I5pTHGDIEiYBkiKa1TxV+6lV9QFcdFHBMRA3/Xrd5HpH2P9hLIcREv02vG
hVn5s56OOLlFy+BCz2cMKxpL7sknDUgClx8/nWxY1x+bkDPxDPyMFJryYkqtIRCB
tQFI/wj3ehKmxgqMaitzda17Xtu4DrW2VYrafWuFrrHLdyxHuMPjlGqm9uEiumkl
2Gcu8o/tE9YkTTKhHbpQ2wCZCQzoVUrIWbnKENJGY5tl9gzRh4PNUf6zBtvbsH0Y
uevN6L+wXBVb+NCYfCv0wiWQ3v5f+DE1rd9WfcimAEO3tZ2kvhNIZNf5z7ljfvPd
8TSd69gm9zzNeU/Nm1kYouIMrQemd6Vy0Lknp8pqmh3wkYgx/XEj+HOucjpOTZfZ
8QGosXfxV9I/nuYDZbMhX+TTXagTGRcz3F1DbXVvOfEkdZNaVKkxIWd/9RhWmO0g
HaY9ZTxrfSLDWcb7ddGpoYvpSTFg9dpr3XQmJQpWoGzq7KvD2pBOwoyIF35217pM
kuwF0xdTmkXM1sww6uG2Pg9NfKPsnOfUL6V6Vbe//bzvVJdJeAgW+RFaowBQmpIu
9HPXsGlS6HPDVcBYM6uTHdDTyBcWmCln3Qj/NDOIG59UMEQ9589kvCDo6ZynkFnc
zUMFvD8r3afF1SV1ScaRO0yg71+AYErGU0HLWku9nu0PH8IOb7k7gD+OCG90ub7L
rhGy5Dt8RnBKlFat5eVyEnJue5dfLrFyveKvJwMYB40vlOrUhZNsHh0Lj39P2jk9
zOym80el7gaSD3YnvH6/8g3TMELfTz6oqVtABexBjLWMqKtzN8ov87f/Ik7OwQlH
Cy1B+GfC9B9n04eNqIPG4SXuyljH3eHqDdFJuy7RM+vIbeFNF6tuC9TeRzX1SCYd
0Wd7fgnzew9XDsO4CyJ/t4Eo0yoUslPvS9v9YnKf7f2JErGMja/VKff+tyhIxbVH
jYXpt6pYCDoxjAP1hdTIywigN2gU+yYmU3CiXBekrWIcF+oJ7OOMaMqhA3YO4WrC
41/wZgrwbReUnQBjTSa6owc41yTNeq9pDZpVbyQD2iPJdUPhMEGQ6MMTOkuoMEbX
mM/NO5iOOMEnOHyeo3imjBHfrFxLOiER7N6IUMHRlqCyBDbwvbbDjypSih3MGIHz
UxgcbY5E9UvlUWhrWe/XEhOjdIpPXpmWefxl/L/PNvGUpxqiRg6+B/5nLHRmXQWK
nZ5D9KtfPC9p/4VQWeMjUVZT97K+37P6N0c9L9D9BF0ewFoHC02/xy+kVeQRugZP
vrGiz/6Km62LqA3ObSkSbiVRIMlf//h2b404eItJ5rFRbkok3cY2XQrEI7a8CdJ6
h1ONmOOZQ87P8594Xx6nEFg10m7tFP/s10hWZ5Nir2t5R3q10t+5wN/WgmmUn/SZ
1g4mwg/DcqrshCekM8eiz7QfInUBjaZb4bfUiv5RJPwvVfBXvsv5R3QR5lZ4ZiQZ
JNDSOg4o0jORn5muxvvve5APjm0Pbuz1cADtyIYYpmKLWt5W16JVfp/GXeXqnaS2
8QFOEW3jj3qozCgG3nAwgnjtDKhiuVxk9Hvnjx3VenQ8jRzMj67HRG+V8EPQd1rt
kd+uBjUpWKQSIJRfW4Z5wTYonDB83AmwREYiNzrNGYkXAjpbMBHOXi71tFH/DFON
HU48f4ygUvold7KeIEF68FkHCczXW/gGRoRIYd13tY6qsUWPR1PgbRPXGVO5stA8
dcK8z3BmeXcrt0NqDJKwGu00VUJVWc8ri6pA/kRi8uuSJeQda5BA3labriSUPVpR
0mJhE2M0Kznzk/5u5lHKEVbZqyMDaV1DRvcF27BvhzB0JBKHaLcJmWajqN192weg
BqpZHeUubC0wn+NT4COqlEv5u8afJd5vzdJZrFENPpnp+SGW7Da+V/vqq1pQpUvt
/R5gIfbr0H3kVI8Nc/LjnZwbUERGpz/1rXiMeXBHK3LEHhhQRmK73Ggj1s0euENc
7Emx5xOYcyOvUO1Q4+D/T0oCa5gxdoRmvyJ5RgPw5S1y24rgNYRQq5EwajCOF0jN
XxMH9iAmVAP4K/+mvmFjgghH68LnbnMmnvKtyQpbMRdaoep1xl0rdKCAp/gHkx8g
TlVxuyvhgvioeNh6DX+oQRMlCoFNtaLbcXX8eUljXPlmflAy+0atb2iqjaTkxJaO
3cu/I9o8MTr1BMqCuW+LD1b67w/QjQf/75t2mnzJ+/ZG87d+0R1A/f36SfDNQcRS
LW6cCOap/JiZwONQKbya9ZTJH5JgSbOey65uqbVL0X2uXSYw4xq9LRZQLm5tJlKl
jQTfO2SzWz9lbG+5og8qFig8P70UtG4XxrEgutQYzJthepTVdHmijworCJnD/1J4
wwxKJnqqudMgTHnm16Xd7hv6MPNP/NSnmCpUNhbbe1yHDHrAk3nhZfufyYE5tm/j
1HMPBuhn89SzV3rKgTM9Q+YfFVY0sr6vWh0948dbTgdR7z2W35IY7CGJgfJ8f3FP
rg2tgO1dV0ob/1ua6PmxVbz/Igw0w8sM5ZtXA1JW2eZFQtqjYfDktAKIRWDlAo6q
wmZY5n7Fk4oyLAPjEN/+6y5pUOC9+sONWFUT2ba7b7Zlgtq+ubx5EsmiKVfux5nT
jzijReOcFvln0MInz7fzcdz4/JwV9qbDWxkTuerq8X1gFgG8hcY1csrgswVO9uyM
Y1eX+NOqZWITbeHl7X2AkD4Vf97Y57S6qh+A5iktR72qdkVM4icY1otwjDT+LQ9M
ZaIemY1l/qQXByZQjZitz/CnjP/YpIVK3RF/eA38MOy3nobCufFupRANKEfo7Tdf
dZnzVqrb8QGD2M9KP/sYGpo81ZG6U+q9ubbTTIYao3O670VF1lhl7HFyu4NTilSm
xE4zxTjdpuEbJdBnqw2nFvVUusKJiFtkESV+d5sHzT5zkE8GY2L/xjtmOCUVr53L
UYGRsE5d0JBspUB45sSN95+/xPPAKugLxn8pnLtGI3E17DMbUfGOK8DbYDWLzFhP
RAuVCPKaelxwN++Q0a6tpYv79O0ngqd0Uc1TgMe5nwgUbAoFSGLM9TDuz2+WbQLr
3Kxmm6WKy+xzFcD4WDbMJ9iBiFEQxnUFCJiTUmpLDgWJkIfKX4HhSIalVH50e2+K
sIzIxNSiBTqLBE/2anQpJMOCzWg61JThGUnZnTc8NDb1k2zVREfxbqX3elg7Amsn
DvOTEiDwmZzw68LkDJZipn+o2OozfDtJ6advtCXOpkzJKvspNN3DfcOMC0P2z8ca
/d2mCZ5PX7uF6HWbHDKsI4+Fqc/QLNG0/s+HkHlHmDIQytbWRJnVHnArLRSVAFPp
9Ki1VUDm5hWstRMaQJqHhTy+yFjdPal3GAGPFwbyXU8HQI8wDkpATfxWneJE3NNv
rVTrFGkeZd1HsbZ53aqNovTc6cPO2cWrv3ghKb6sRGvjP8jWl+nPGcy7nRZffWuE
YdWdR794TpC84s8oXsr6JeuzhAMC8YrKZK0Bs+uLVfNVZxp4TTXtfVI0r9vyeebW
hrYOPeCmFZWUWdBPa9ycFYCdyvu57EEDh8NFeU5IgFn5DVhpb2l1ogqf9gc/i3B0
Ev87yJhJYOa7Bw4+LJ83v33/Za6BCgUs7gxtCiCamiqIG+aSNp35SYWbt6QdMxiQ
6uwDJJ3mLqhrGBjBsxnp6UlwPiaD7gcRJytX2nGGQyfxcdpFMc8Ul36OBMDgTt4X
SlJ8oeMWOSBD6wge93lEYnriTPX1i2riMiVeikmwTwePgnFV0W5hiBUgWL7BPCBP
Oy4tXMXyoo9lV+w4WEDkT3XNQeqViFDW6ocF6w9VxsafBj1jx6gdmNaN6SuMs8Uu
zsAmzR6NQTfHlf9MJ1J0iWSpCiBcba+9nDkMzdCvcW+BHVAAinxxMFrlbaN0r0z2
eQB367SmeNH9DS+KCtrbKH3EPgDpOfDolOyQqJKRLFv2B6F0nZ3u4Dj96ocbfMCH
06O1V6QcMlUdHCWwhI5PbT5gVy852P4yHe2QOGnP42sIKYBy1sqUdlrfNdQ6zd8B
G3rwDkMnauV+PHd/Wnf2rg+hsmlcRrDcPDWhA9/sAt1kqz8aFDAitH6IOqBJQOXt
v0v6hUyW+2lcnP9CtCuRzxw6X078RopLLkCX63ryxUMdwrR7vaq26u12UWsA6sRl
f9/f/Eh5SnYYU1eWEoTPiHYT+6LkaLOCRz8E3W2RF5eJo/uiZDGUc42uRT0v8JBg
wC4grgBHh0aKxK6/2AsUw1bxOZAtwOh+Bjh0K1dIg/Uw378eTAkekcV6bn/Vxno8
EnYa0nnJRnaZG/ZtwVSypdSMipzvkzFHGrWIRvoesohktc2qI64jpous6JyPAU2J
vMoZB8ktFJb6hk7Qqt/flxNWyo+Up2/CFkkZJN2jcq2OOjrnQg0U3/YAObrzzplm
/Jz/LbkOgMorHwV1rScQIVWfs2pZtJYK/3H2AELP/kpFkeK5tYiAd8KdgM+IhTVp
qnvt12T9kK6Dw/TwJbqn7A==
`protect END_PROTECTED
