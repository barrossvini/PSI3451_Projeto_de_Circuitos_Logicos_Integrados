`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YgQiLpjq0eq0EZUU4ebeJYSvcOom49atpMOphNtGYD8MBn9X6r1OQuyBw80AklCx
wyxNoWJKzLHkBBbAmaXRFZE9JyLiv5t0FMtpxW1P44aXgFLmKC453NhS4iXIxm0D
PQiJxnTTmS9hbX1FRcsov57m7Kt9zrSxW4xEVJWOB2D89YBY/CzZCdOLTGCedlRK
4rtgQekbvuUXJc1vtafYtqj1mOgJRwLkVKyShdX4KNmKR9hijoQiO0HWcLPAqjAk
fFJy0vVR3NsgA3yrTA/o1Fy+bVyG0GQjxWIL55sCic8GSI2aq2BbOhca5Z1ynNtE
hEaI0JMFKXCEURTN97cj98ISszNMer26X203qHnFw+jc/KvtS6/rqOaxXiRDJ9vK
zfiDgIJgk+7zcWRQVR3sOiBDxRBYTcEkI6PCymTbtOuJXK+DmgfRXfJlqyWh1+AX
vXCzQDuqPoWMIU14L2tZpyAusu/0aXjJj0/HnEvAXiWKtWYf2qLIoaDT2qUX+w5C
RzVvWVIOSh3tn1zPbnYUNzTsGKhHBTO2hCFTRiRTVVoBKJEO/mf8AXH+UcS31ulL
koSTb2SXRZIb9e2DNq86zQb2kksR/6pHN9hZblLGiO8TPegN1Yfi9/Ue10M0zd+F
heKIhInPKY2JZqhgrYyBriMS0l9KXhIQUbVpf2ICWg9LbdSCrUQ/DDsCT6iiz3mU
109UEVH2M4zOswGQQK+L42yzQCHF/bHJ7ENO9AH82ni2u3xJJU9HAyZXrIQDBCM0
4uEKus72h3KUNiNe9K9ruZWrTDcjiHyESdmThfse4Zh1hcb+yysCJCOCTQGRzEYh
Q5Dx76p+mJM3tT3PdgbLkCmq50RhXh9GLVLdQWj/lHAvCRx0ZCI7gj+krY0IhNLL
SXhTK3qge1kdcykbtSgDuGH15qCANx2L5iRq8iO/gtyQi54WsGCR6GjhcKnfTE8z
jYJTBP/i2AFqzPJsPOgx1KcxPqZiO35ggg8qZjTGk79kFiG4N5x513UmzxEt7iwo
3VrQf7W9eHY4Kytn6p6ypYlxu24Se6ezYlq7CHhK/IIzws7qJB26RTvA7BIkYjAL
SaQdrAImYZR+Y+vH+GAmil+3TMoSM6tAzxQRbJPXQWTrp8x/4Gh4jeCGfcaiQSQ+
YbBTyrlmz04l1jRhM1W/qh7rIo7tlCVf4YN6H0nUZq12RN0/lJ0vXvmf8507lCGh
yngNoNfvRKaSrecahekUKzwASzGUhP6YvxkfPNeuNBDtMcWRdH491RpTZvie0Kit
sSfRO+k6rIvfp3zGk31qLUoHxEJh2OmHelFaLXpRKChkXhcs8oqn56wMdQ5IpvkV
xc57hyZcDflSOKV4s+fwdsEY8vwhBVr3AMBKIp1giyRdCMDOAwIWzABfIOSo1qC8
aXtnquHlMZqBGviYXotR8SgLHqcC4I32hQ0fhUyZ+XfKan/hxPUQ2ImnBlPItlc1
gr14lyoQTjDqj8RfH0myNGAjVAK/wSExymHHZkvj7cq/fujcaXg3JjKeVxeikRgJ
3M0lD3IH3r9AWxFI28rEaO+uprV+NjhW0jaGPVCfTkpbvCsvJthPppH8GJghCgt6
yUGZI5X0muwNNhq1exUYHojbGyxrFnui+4v3ca9O7Kb2QtpJ6NnqZKRGwtpIuids
XpDOX0YIyaId4ZN1ROlXg0q4xO8IGOML5y3DTviQLRN6S2MN9E+iZaJf4EsSdTRa
0cnZ1IW0nofKxSFVMQBKaGQNzxO1dwCp359RrERYgdyvZgaZ7ORQn5a1N5kja9aE
s18jwUVbpsi8k4AqMG+uEYzPotRYoXfjNDaFcxvDKGe21dn1Ix0uL6ndSYzOljt+
vf9UGKwsL4BBuE8VNLXmwFDGj3n2bkelsS1Ws/wJulyiq2Q4LGPPEKta+oB0DjMK
/OxEDx9s0KPOWuwAwuPtt6mKMfkACHo3M13RI5SDYzU8sW2wOrO3dxrGhflQMx7m
5vUvHBvD9uRiXKb7XHn//SB83jZKFvOKv4NoO376WFiDPhVW7KJ+Wy6JdRnEwJBn
JQr/lLaX1SPGNX0fwTrxPQTh4dBPXPEsqenYML/sIzDZ8vvQ8l7q0VBJ2PWEmQSs
D8C+6RVlWa04QP0tWuY9dUqPnudHb7szeB8aTMMBI/ZYojRNGOmTwfNtgseKlvaf
kP+D/WpAUau61hs7prom+gamrCT1c+o+b1Y1q/NjfCg0v0St/HT59uxsgYSeP+aZ
usVh5FSOCuQO+jlwpy/OkoIMYEo8iX7W5z2gm+i/AHP09Gs+fwAhIPwI3JtAHh/v
wzbhcyVbDqHTrQyS8XsVxqXS/y0s/5gSrmUtfZ0casp0HWLpmvCSi6FRUMZtpGvv
2apmp9XYUaajhUsFM6HnL8ju/MK8SDhr4VGOi807HaFQ21smEGNGu/76/oDPmerS
jdGsc8//3wJdy+f2AxRoRV6HiABtjGnA3Ax5icLd6BshbN5sAhHqYv5XFElb7QCs
r9+V9dRAmhuWk9VeiUWa6t3E6mLPElZ/hnBJw7xBa1nqP7OG0gNg05j/vR3sej/A
o9+ZroEl1jUB7To8xPLBee5syA5uMzkwmi2M4nnfq3uI6KNr71qcIhbeS6EJsKpM
qIGRpuY8adZSgG+fBzqpydrORrO+Qkd+m+DahbhHQiKwDJSJWyRG1EFPM1jja4q1
AXhfel1VDxyweBsBYZ/rqkl5Iu1HWg9qUA6lU98fVmFe3A2LTsl+oEj0KzqxP4Hy
rGbahM8PrtBIGcDgSJPVKoMHUFrfLEgBu+tiNIHuxM0yKqd9IpGK2OXBP16+K4sL
lKI5WH7yz1MIMi9C/tzvbMOUpNBc6scJmXGEEMGonv5b9idvRCstPgRz4h/3QJ5m
eQ4EnPDtDxadcNdqFJkbCZ//31bkItNNq9TYs3GdAGM2iBN829vlM9F+ueVzamSm
/zxeU3xKiUaqOxfIfSCto2lC9kdcQGbe2Y06NkTnLHIDMwcFJFhdP7lYGpNgjMI7
/+e4wUT1n5kNz6xU1tMSKV2lbyCt41VmLtcxrPzsB4/R0XIX5nCyq8H8gE7bBOUM
7hy/P2DtkkCPkEoU0Fxwr0RlCJnZHemcI7TQD94Ieu3wKr1BBWkGHBqk4+//Rn1g
XQT5HIUidbz68heQX10eYXe0rQaFZOr0NFxPd+/QcIIgAPAoBanZ4RxfkdBQPBED
RiLB+BEJ8Je/RHYIG4CPgFCwz/kviAxNXuMOIJ80OQkcmt4JGSMb+EacC0CpMOmY
fF+Jox812NdjoP9KtnsJvgzk7rO/RUMtkEyl5Qsn54nEtCxkd5YOEaAi/vTwWo8S
/Hf4BR+cYbD2LiTHnDADxzUE4BqovjuGU9Snn8nZIf4Ed0O64tFZFinQzXkDsUz7
Kiv0da6r1Qy9kpkEJpE1at+66JTydKkCKlUgB+y7HjsmOAqiIy/eZcv5Ig7ZnxgZ
KDM8+Q1AfRYPRXPQZKUa127Epa9ooTfPFYxZ2943cFFHxAlFlmdcHMB+2RQkuOHD
VkLLnly7i6JY+6V4IFR9l6VaK3DxffEVSez417RC+yJ69AlNY4Zm386aeWCm4dRE
IdYfIV+LJ0gtdInZ2LnQ8gRO3/pSHAT1tmN6ktpAVCG+SIZkFydYNkI8Hj5KmXoN
WFFaPnAhSDXxBlf++4CujuCaG1dtz4W/NtMXAy08e0MUsTTjbWbNNK/ORwqoiPJy
OogVRjBSMbYKppZXQ9sbCQ0+23fjiKMnrqePg+BZ9hwENtHJl8P5w+I5oWB46a2V
vt4DPjwwG+q5pODlNdM+XnVRc93gJwWi1cPPo0fxi8ygPzRaFP369upw0ZoOmenw
ZOohP3nKJuqMOFGzO+CZOHZe/0L3tBT2/36RAV7/IJytdag/wPV/WN4Rb1FphhHa
zY7d45MxOX16K83Pk0wJWsLH5Irq9pwch0JTbLZDPBcFp82sNeKw8CzauKsEQY2M
YYcLSp058sjRlwdSxO8XgESDzTCqrzP+J1c/Ev+Is65kCDegHeKfQgUU1Qgi4kfA
kGoKPumT9Uj1Q3E880zmFytirzE4tMrhKirisGze38GRck6kQlzsS1Gy5tDmqHGS
szG9HtSOPYVINw3jKIxlw5Y071sz7DKUE8tR1RSFHRUbQHKiFAEp3IvkEiqXrftO
TZOmJehZoxjctn0TJtr14YgFukzVdHDRWKvCCA6khE2HGOmto6WmTe0GoH00Fe+P
8XN5xr72jNE/YWCuqgjzg1TbXrRXLP4F6ld5Q8ZcNHuRXXtxIxtn7tm4jPeXVOC2
ecFusNeOF6AXEyiizzX0kaK9j7Tw20nF3aYJwVbVrRIJWQwg7p5xmAvldlYQhsm4
ZSi7DiZ/t9P9LymsegCszhQXZUouIsdZEkC/ivPB4Pom41C9K0lAFzd6gEwzntmr
FfIP6UEcb36jpSR0p7OiTm/OgLwbgbpZPJDk0dGzeuKf2dR0fxCosDy5TwqJw4l7
iRqV0sw4W60+hIHGO5/ymgp6eATYTQ6Vex+x/UgnS76umz8y7DnAXk3qGCQoGrwZ
Fl+VTpMjX8yCzwpGB8yQsbsL8e2BO11Yg7GBvJxmsZ59jstvJgDYUBu8iwvIdAea
5ptMFDYg23cn3RmJdZ6zFoKIUEQn4u1AoSB6hYt8A5PNII4B83MQAU+KCGrI3REN
+HHipqmrF2J9DWRv6vT5imJi9Z4kK5+muSb+/qwYfUWMtppoW/LnAItCaxipI5k6
gK88WH2zXk+ay55SB/oSIagqPJSxV6ahF7ueXb2CKMYJ2MyXutX+OwpXi3NFDfQC
cmMsF0DCcmBlVPXJKV3L+TjA7EU6Ukpn3ybcz59uUIDqP4qiVZMZ4gmDmMRnyELA
nK+0nfYpY4m4KLojlL+UXC9IQ85qWN/hf6rolOwskK0HfOuylVYnVDY6BvvxxKQ9
jQYrAjDjr/99/I1KfcaQ8Hp/B38Tl9N0mBv6FWE5iUTaHibopCMe8OE+r7cTQTN1
4sEwq5mOg49xkcKuDuWTNeSJHnpD0oT+0bb2oAydxyRcR6m117V5rv/ujoX7EZAW
II3SQ3UGXuDi0gNL2SxdGvEHKC6yDqu3M4Pa9LY1bhwCs4DTToSapofbppJnD9p2
eLOzDr+sH0dBkFPIE79Azt/sN4fWckOwSVVF2R+8aZi7A8P4VJfO1X1hqACNi5lw
QfqvTWZwXETDKunV8WSadpFUaZOTPs0drWfTcrPlO3conQz5YZaDSkusfJIHtJNQ
sio8U8balc+ne4OnHbVnW3wSGverrtswuUIhjOxmpwvAVhoVoo97PI6/jiNf+8+H
a1rgwHDXyuEc13mDmSF/8MjjLgIwMgkR8IvU4bJLH/XzJyhjYDnVAkcp3TKeQIfA
QQjq+wkTrS7W1OVK/AimI959gSfpGOeRFyPz+Sw8ylwwCdygxZ25Xw8l9x6gQFdN
3sEUwouckQnaWupV8lSSiTm1TqnUHH8uq4ga7Tcivdo3oDf/FEeUr5lGM2VVeAYD
I0tcmg7xRnC90GQZsHicSuMbUg2PCIJ1o/iYPdwa5uXSEwk33ByQUO524I1FM0qN
OcnfCvNIbPNu81p4icc79hRzkmcxNhp/vlxs0kqFHAz0V+j1lEvKGMu6nqrvz3+K
4h0OLrnqASd/oIj3MPUdWTPbFFItQwoI0pYYztNviMM/P/suEo8YhBcki2Ltk9PS
LQ19l2PsJcapIu41Gg8GGwyeioJrmFaRwJV3mwPjwpAKRAXsk8FrJVI1ZKHjxZ2a
yGdKDi873m7USnbXDLdypbElItgA+i60IruAxgNwhAqBjSGeKn/lDYxOSDPHT8UZ
TyzzURIwaDp7CFuK3YRld+FqKHfV9Z27BnGS8sN5eosEDsjZaZgx+TeNXMQOgIzM
skg15MFOYPZmhVVh4dMAsEXWID7NHAuyxItrwchh24+IPLjKZL6TMrxlZ5tCWdhy
HelnE7E0nz+DX4e2P/RHc3WUTub48Hy/54lfC8at//y+dqSSZov45Qob3jlhEbAF
WEIw2ktiC9e9p0cZm906LiTl3fh2Bp2aBRioAB0d/KQVgHCqX5ICbsDr1mL/ffji
JmEO9AcX2LVMIpAvaYWhRPD5hf4P8atVXH9b+TnZ5RnDLV/478VLl2qvQfx0MFmf
GdRrJhXdUbABIovQVb6QFR42DCeHTY2TQmEhf0qyrstTtlV0I7wrQPlJjp9qL43H
JfumYRtqXsk8yON/LtQLefMHYLp8wbGGPYzkiWmZ2FXiE2aQ1GmLZe9Gn9i23HjZ
qEgvls0KKLTIwB0zUw5Qzky/l3v0JkIoQhDQLkl7N4YQvD2b9UBsBfFer6MPkMzy
zAqfePf7yr97ZphE1JwOYwpti5oA3fSFMgdqrGKOL+Wx3tWvvquiDu0lJNLvSKDN
iIOlmIJBipom8+zIWMi3b11dcpT1//Q7Ja7GDhBLHbDrRj9Nmv028M0qo6T8bKEu
0dE76SvO2NkhscyjElp8fw6cMpFSLyaNQ0bGmKrsFnFyphrXlO6qVZMOGl2SF1bS
+smBU8XD7pirEuVpXw51qEIHl4MHSrfIRXulvlFBeHUbijT+7q6VGRA1eW8sW5wE
23kdHcapjCFuE4a5vTfsh/tFr16ECRFBRjmDhG5fx7sv7uHK1PNY/gjtZYbLh4b5
PstuPBFDhYybl2zgSwL9olzXa0ZFfgx7OzzD0oQqxjG9W879R9TTjY7Xd0jFN4SQ
igR4L7dAcbYsFi6NrIEGGWckgkitcA2cjcpTgMuUeH1yc6OUta4ItORBH5B+LCN7
d4wWo2YWFRyvFeayLjTsJqR+JPxkfzFXen97B0voqwUaL7wgyHYOBTHeDiMzElnq
aAN5kL0rFB6FtXFsjsExUjDDssVT+LdvvVOvWcuP1SqLul0wU5+4Q6m4ePhiSFNw
uokpQwcNF5JSS2g09Vl8y8b1791lfWe4j9a9jwVOlO1spsJOvomtPUOB8EnONiJ/
1txDT8SFyz+tp2cN9JasYyIDnMjK1LeNO5zYSUThAc+mmgGXkEh7gdCillkGCUez
Vg10iiDyOty5SZ4EBOiVOMu1cNygtnGK6NKQjej/lDjbt9aSgvjN5Fc8/EwMOgh0
tRiXwgiE/ZIJtUeJFkZmqCeqXKxLordMFo5T9VWE6y0pQJrbE1DxNq4z4HAkRR2b
QRmcTnzqf+Kq/KKBECJhS+1KY7ZxaoFJjUv1S2gV9FiAJxKdkkrKri/GuzWxSk9A
uYQJIMnXkn9gKwNJrounmFx3n7KGUOQgqLTCrxiwSp4m9hl1VAF/qom586FuCWI3
GPXqSC4Q4MIqy5Zsz8YDTTyqvxRp4YvmTCScDAwRgvf8+/8F+qdwpPtmAAxc7vmz
hE8d7pMj00Wisq/J+ejQY4pUfJJrejlwdPjilgizabyA/XhYrCGXwWRCoK1lqt2J
Tz7KCCVmhQPqBE7oNRkb1PP6xGfeeUO+uOghh3ucgRoS5gsRaw598EbFImEwIGtp
XjezXdfbtOaR/jlmuoexN9cqCqlZcDKVqoQkqxuE1cwIOgpFIHR9NKK5zVsIaCSz
q1+yo+KG0PWeplKzQtQGdQteYmDE9c+mLUDsu0IVFU7nYdQ2FHvDJIZcgGBoDcRk
O2dGvwDZrEpYgILto6moEtT6fqMPO96eDeCH6NSi83u+c9NvwDBcLnZHmKJYTCn1
Fd78FNdpDeWteo1lZhuqGM2BmW7S/iZGQNc+koO7cTnyDzEd69odD2pleabL9UFe
r+xiGOzU9SUcy/pqIenct5mKVQcRRlfVYHrk+iuDOJHFrwF1iEPICA8CtLknkmi0
zGejuYvvfCrmdxoXwB2GnAO06Tr1P7No2noaDoiyBqcL+U825+Pm1AHD82I6eyJu
F2bk9ZH2Q2UQGXk1gIXNrTEmFP/Gxp5zxfWZOyIAHYsFkHghb89cYFLwGXKBDOeS
qESaz9S2VH7jA72COt2kqavBTweJtjCm1EO40KVCd940dRVYCrviJ6zYnUuW8UBE
/o7DuIRFMS7X33ozmC6jIv4Zh8uzO3KHSYMRv5FqIEO0naVr+2PYUkdPkv5Mi53K
si1Iic73RCRQapEIfUncwoJc0nBvEUzN4BqKp54Glbb8xPV0gZAfA6+DM14+EHuu
lIPdhD4ZEKjOFdxsoxrxDL1CBsRFZbOBeEi1MjkTUS6ucZLNK2zbe6iMg2bZyGwj
kHzEtmYPMo0bTgtK5fWS3ZLLnh6WJztGquizHxanp7HqqKPtdJJ0hbCzHzFcX+ma
wlV687cxnE+9ogqhQfSgTTVaas0Y86FOlXfoxInbbuiVAv/l4ZG/24KdOoCjLyoF
grGbNaIlYOP+W8XDAIZT0wKutVBUHR4uCE320Ji8vT2FyL9piVvRRh5xCgue4stO
2L/xPFNySxEsaCN5aXVb8ISygAnlNh3GdVukaJpdAONMI6j5WC4QpVjhGcXUUrLg
Fj2NzgeDCx7hPvZW24R7l0pwiVjCK/mThpN+iPS/WZHS+hXyzaRN4TchlXADOhJA
m7Xqw1F+WXpxzF9X/kUewNyui2uqoBAWahIfQ/XM+RtrO9V7PfwgE/IfWr4WU0q9
TRFxsflJk6qJ5jfh6gb5rOIg1x2UrhmJTmpwVa83XOFoKiuTsxozScLBrmp1Z6ee
+rgaRSYAOUj2DPQhbQepbj1zRaIKsbTDYWatH6yIymZzeZjaBVibCDtKOLDNM5t0
FfkDMsZyqS7g+lkqGnBSkegnD8sO3XjHXsEKbI5eUPPn4EmnOGV+i39VlBqWb+pL
2jyZLYdNXvu0EoDniqI6AKlSKogWQTtd/msNqd57rH/R4E7JxDUk+cSA6EXXfcZW
X+L4Y7xrhxBgjtuwk1fODJd49skl56nQ7DJEmxTh+1aHwt/g04gXdSTs7ABd4eNx
z5QZN/fCtBUqnqOXsQJFc5FE4Sp8G5TUpKRfk0CgSA67YwFvfXsOvy8oZ8lJ/Zdk
hRA3c3fPmcJsB6Vc08qQ5yABzL5ntpLmpi4CCvfB1Evzy3BxZzUmgKcvv28tKKwX
eCBzBL6ZMNM8SpAX+rq0LLf5errRSf7eIZKGJd1tPFfPPiQ8PcX849Z75VHT+gGH
WOJPCSsiC8Z6nmOnPklOcCMy9Vq6kowJFxDUcaZ/WOo0NxfdZJe+TncsyZHXCavb
4zpIihnxooRk4auUFhIRDEDzcV6P7w9vExwqJvbyk1sSSufRHw3yyXoX6zgRS0IV
ONV6Qe20+U9kh42iINUtPvqvFwachC6F/y7PQli2BSVjldKlYwrSqr/uXsHfrela
EZclsfXROJzr56JsdIhfAgGpnSopUt95kkoOcGMb3hBxNR7+xcC1B06yyFNGJwdz
t5MkNfsjLMTzmhlvB5vW4b4Q+qouJxRQC2j5E3pamUFdVpO/pVgGTdqFLEUZe8Vj
Z3G8tVcfPjYaEvg+D2r024e183rEVAy/rIoQIrao4xOeqxl5z9hNiW8UBrelTqgA
ooiMrk5DNP5i0/T80Wb6amNWvl+L6x7vN9qQ9M0aK7CtSvTABI24hTh61uhA1IIH
A0j6dYYhrZ5RWzIisFAkNm0IaeJIvln/JT9bzfXY6ZnSFOq974B6TS/hbOj6DDhs
rXuymg1jRwltZhkPdJLtweBY/MR3i9lBZNG8wytXusrFq6CFOUVtKxdrholjJGBm
cpH4Xs+L3R/yLPQjKvn8Ol54e3qWvzu8aJrFB7ZRUAcwX50TLyS0TSTlPDKwVbLI
9H1PUUXs/4RBSbS7HBnu3c9YvuWXIhlLlnBQi/3t1ldpWGK15laNMCM32b1rt4v2
1K9E6127p5ppTEfKCSom1Rsg/R8poNrMOtZ4p8zdKYaddI69rhWPydzgrOj+YS3g
YEd1RtakNjgIH8KIuIOTcprBHAg3VA/eNmZD/0UbiRzUh6TnWCd80AgOTy/xEqiw
rpyFTc7DJCjqwwiJD4MV3ExfZ/YI6DFUwIMX/cO1PXgwPwO6yg2RSu7uYkLpYj/w
vY2HdHDO+ZygSHFKIL9bAe5FpOUR9eij8TPJLNldSpSAEhMJuvj9v3hvXtrcf206
YiFzqm1fs+G5JKAQnE3T4yD2xhRnoFyiSeqApnL2ISwV5CVdYL1ra1/UWWkX0B0h
2wz2ZJGefZQQfIh9U88llkFw061Sc9tNJFRopx72hynr/tyVFKi8ATAlpH+qW9vW
oMOXOElcD/BQC7P85ds1TZL0oLVBMK72HdYTPxhcotX0ltrQQ1lgmA0g2nQQiLQ1
4Yf7dQqkGnaYD4353j752rOXpF1TAU4ERtXo8brgJQxdxxdLAnOgQLV1yiNrW0b0
K9mvLtfJjUAczMsFIx912TbFku68zZbpO0JXOAQwGCUhfxUEH8UwP7KXS7HNkWmx
yy31PPbvAwIGwrpsKeqC0OTsCOTQ6H7iSvAePUumvjfnwfDsIjEJTP2KggjiLjpU
zntGfunDP8GDF1s7648AJhcU/Hhrc2HgodlsnJLyCOhFChAspkwHXuwK+PfOntkF
XWUV6Uqxc3k+/2Vy+dmJN8KpatJ0vjga/kd7/XprZOxYb6+MVWEmi9BhU3oP5hFD
7t3P3BX1BHic0nIpyI/jxtLT9bguKK2S58+QVQmLxmd4Vck/ojkdbapGF9OjR2lk
XzU/fe9jJ/dFg1dg6maB4HKntuhHUPOeiRmIubCH/2mr3MU5hsWT/YHgx/SBfxK8
WR5kk+GBOrPmqS/llrudC8SRoWD5tIkop0ZhEYKH8efcq3J8A5sCNnyQBPD8dc04
erV2FSiRpxRj7cuhNKfgNGgFAk+gazFZ0UohdKOe88hc5mk3J6MQD3k5NwjiznqM
j9ZmUCU/IvpIKIQfEp+hHtRv5o/UiblU2gsootIfAXWrRZS0oeTfpov9MhpOqyyQ
SIxBUvDLZLc5pXNDgi6VmVMYDSMQfR42Qf7XY/RhE7NO3HxY4x7zHznP/YieZvY5
ClH8YmXvtiB3Zc8D3OvJXyyCuKydIhbALvMNF3QSylqI5o77FbfeNuVP7dDfFXzt
w9yatiRygDjcKrekXDma4rCqAJYqULRVBdF8zhAxSexFryf0wEd3FEbvwmC2UsK6
Iugxo5Av/Fjt4CWc0fQo1zOa63FnORG1UV/4fGebrnRFQc3IuER/ioxFHP1S+Z6Q
3kWS03/cpZL9hqzL5kb98Kgcanz757TSdxFSzuuH6tB7uYwceDP+06ve+NFzSbTR
dRlXiLGkZw60+JchTAiURNZVDRAlhgaM1XOwKsnrCmu7FAHn24GULrYg/ZuXzt78
JxoR0/pWKLzGECtis4aIdNmny1DGbSA9p2uyJQanBL1aqx9TbNfHPfaTVaCSW8/I
ne87Y5UsRoqwZ29x4fCmZmjOUNiK2RncmEdCXwamKxiiqqWH81KZITI2A80zZ2zY
1qz5QP/J3YUUNiQrCFs91cHQk1xEmjLKqERE7YL2Lcn6roT4NNVxkbz2v91TDRCO
qgL4UEbM2WNL3kHXo5K45owT2CtqedTeYIfEWjpVnEb8MWqArSpkB64mGh4gEq4P
MhA17Cym08BgUIw93tPP4BjBtxERSnqBVLCNP+GHGQUtZYBv4QpWVaN/gQjCSw3f
LTc4aIkLhK58nK7nDgDdMmTi+gbvivMJaGYgrO/gIPf4ZyPVIb5726nP7aWmIelk
yZUAOoW5RP3PraRd/Sn5nhN1/LGmy1alH7QTp5qV4l9edtofo1EQrFwHNPWismnC
zjQwp+89KUAU+CfBlQR0N+XPjPQ/CUUiPcaVMzYxeJ1vn+6jh4iaDLXPFp+fDmZV
oCcTaTsePw1h4aONQY0m4QHaviMPbeSWXZAD/JyGDA1A5UN4MJnaJREtqdniwRDd
yL9wZlK/fxDlGw+IIdHoG1+5Fa1E02C7yVMmeCVmF2Bxz0hsmpDFnoBltHUbNWU9
V1oPMZ4HIa51hbqaqu+HX7o35F8NeehP0beGUUNf9ADfgUVwkl66Itj4dQY0jUO2
p0TTMLrxfsJ6O1ObTofMNLY3w4w/v9Y6PFephUBncGxmt8enY5TQXNeTPRrHpU5g
D5XE8l5c9IDBscVVqkhIOuyH2kltc1GMVU/j46pWnS3W76WiC5eFjkNZsjtM1jIN
YBelYvJi31lbuLhURRJwDUy3PbrH9YNZ18LAE8ZDYOxtHzaK1pwy5Uy3C6/zmVWP
LMR8zGItZihkR1Wv39DZev0THFrgB+U/LXc4y1cTAEi7maoIPqlj0aGWkbl3jloR
0F25aXRXprBs/e4/c72zvx253fj3VVFc8gbg6VxD5UC17c4CvLc+jhSx2O9nQDT/
ExOxpKtxcBTGX+5VtyvZcX549fgHU6pheDvT0UPlrkDLvdYjE16mONOMgMh8e9pF
AmyW+UL44fkQCClnG2LADX6l8iwZnkUG3LL5UH6dYpwvSg1A6aJlcmDQ4zSkmQtC
UyAR1tJLytYmb4WKxPw8hEBWGjv9PHM22Tun0KUtAtjTiVqjbls66cKgvG3mAQ8I
IA06Qltqf27Xe4brKV8wIeoBwEJwZLoWnvZcIkBR/TUTIc0Har70UKsiqVjX2kyL
qCuKRPFuxUzNm3PCuRFHygaEy3INgsPDkFzCAmrSpOMcgtG5KlPATiG3l3qXWfiM
QbdNcQZ2ksamh/fmkbemouotwDc1Wy/b3aJAFfgFaFMKs2qVag2UDsCdWYf9oOGk
YfeO4ndS0hmWjYbXf7R5+YdvNPfzqnWTvqRoYtzXcZe3Qf4ZnPpiUOyW7IgCxNZk
xVw0MxjcHbZNN1dO9rYykAQkItQsez6T0Zy2FstJyef32IYNWFURHyQaY1LC/oGJ
F+o4RACx0YIM7+y6M4Z7DjL4XfBtIqkpqHCsahjmSS/FHwyZg2rKif8b5k9BH3RM
dH7Xa/FtDWdbNC/5SVICiiHefHs/C0jOn1Q4RzyLueoonFbzXajqq4IxMDVSem3T
3CGeF6g/bEXAX0yxjRhGEwKTFTsDirNOk7v4bX1yn5Ut5IpOOOY0ZPPZrv5ugyFb
Ujtr+bUvK/0mOiA1UPBq05KnJql3rFPWhY/NOqC9LEy64Y08y+HiXUjtz97ZxmuG
D/kAyQhuH97L1fcBMiPD06WRJdiBUYvL0b2UYnZB2e36CewmBizr6sQkogcvkBn2
IOTj0904qIpT6waY2XAbVE93PIWt7d4fm5clT4L1JBl4egNh79Kj1OYkRFS3AFxn
g1jcDmvZYnROMxQ8I9gvu6+pGMXDZFjqGz/s6UNjBRlQPwvmvCvyAdjfqLuuesK3
nu/W2bayGMj9tSakrD95BrA5zyeGMUUAt4zEqVkFGTp3MIDjgnXsbI1kttImq/pb
/7cfAA1LS3UCniVv9Y6/YvPreKjlmVzPOU7KEEX9fOodgplvEeWpbVZ7jAaxs2h5
sjuz9mlqsi+B+GPn648CunsMLATjKuZ4O2f5S87klRad+jy+6iSp+a6jkRn+Gbs2
ma7BcdXXCl4Ga8nenaRhc8O6GXC8Wu1sW2gxY99EhTkqFDVw5uXAwZFGZ5RtYUe3
u8bAivClXWMWDsYzWnLbRVB7QdFg1xFyYmBT9+ltuzyJd6BvvQhX3ILqEtSb5Shw
9REe22v9ZbawwVC9GnJqBk9oMEJwrNxe5szRIi9u4fAnLdVemGql6T5Kf0HbbCv5
lpZzOYJy8DvNgoNr8s4hQqjX0UQywv4oaau/v2VS6QJUtilo0+abRE05QIEyHfgB
ERFLwrspho/e7eXMIUhhZTq/MVC+LgRW5lktkAiDGz7EG/LwSPLu6+6cbhxWf9gI
xCJkztpL1G2DFLkzUG5GNY/PfZattU1Znw9C7FD61Xt30CL5H0jagfHNnnu09ggE
lg2mP9BW26m8qoQjMm1MzpBmGTh82Slc4gG/nRYtl+A54yIY49BYKQXH4fh1ACWE
n/gLaBncykCfUbzQaXd8QqC9wYOpfGuh0RG2aFvQ3EOmvNrYcufPRdCotUwYWiDx
1L4rUpG+xMLdji9pJTqg+30Jye/OalJwnEInk0jaRf8QqFFq/4y58jkYBm2CXD0n
68wSUkniDDBfF0Ehvjw4MeukH8SMeycUpqmZ4AQU9f71nnmINhzxD/834dmrtfaA
3n3ez0KvOCn/UY2lPOzBXh2ciC7YaV4qf1r9xt3vKn6ogKJzR3aPG2KUcdQbRUBj
+I1W4+VfWewDfdbSdB0AFyLpPZXel9R/EAiN9Z3q2Pg494BTkvMlVCQSZkg6g7kY
9K0ILWhLKWUx3B/aeOB3PjoGibjYGRWXfPZ77aEJAxPt1CT9BFI4lymeUpb9yjgm
BufJMzCZvcK/mCIqhpXSpindAfTQwEfEAfyh34LUUEfa4DwCuVNNdvdKuAVoZ+4x
53l6sq09b0CIPUaj2/nZK7ELwKApfj01ysZTj0UVtxVyZI1m/NAzkfEgRart9eD1
6T2tl5c7KtDDN3cPQ3NVNNdvjHpxr+YZu0XLRvuVP3HZF8lzGFtVUUqZCnycGHvP
jhi2lckuCQUquS1FF+Da5Vyv7PSbJ0lBwEk1i9QP7qregz4kplC0NSz9bTmpnfjA
ZY4mndJfnod0qXsgiGfpaVAnDYd1ChSPTGsPw2sUCZxn5l2j0EJ+XuVTNJggAoqL
JoqgYMYZKTJfdhVKV5cr42olqSbNi3lGAa4o4tlOdzlo9n+JBgwri7Ghw9N7E45e
Y4vPdHSlpK9msPx5nybVNcy5QJY5oMAMacRzuxvJhk8bnllQU1mueQzG/0fFeUef
B8pcco+JBffhxvloW0kj38MMDLN1S6IhasBgj7pGu0uVgtQaT+K9uoZr2jjdgE06
E/HSpwp2iy9BLwen/KU4L8P4cI4z7HezkIEjm3gTFkz3vhIMuqJOBf0YT3QjstR8
e2dasimJeVTOdz7i+ravxrqPHtkR0o5101PLkg8wtCrHy8SvvXhjoF6TFJJHPzKx
NnixDEfdRMOx567phfWqjCIg3hstNewdwsh9j3rpnuGB6jv4IyYyRLw5EtNWlNoR
xsNLBoZIC99eEtZM1efyTdKQjJXJGL8CdzWvcSurZFiVpPIFmYsooy4dfBVWjnO4
LBCe3zZYwRtcpQCXbxrZxxZkFPPsi22YEly9pSjJKUDUorlqcVYnYhyfJWkz//3b
fVKYW7zXOm5YTWlIaON3fgnCeerANwMye6VYd6+9Gs+yGOMyYsmBDEWrfkyVYXkV
NVLMJnSoX1N/qQXlCOmmWkUnkOUIf6bddkF6n1fWR+ADxqXXBPT1mwy6/nqHnhvm
fkMFk7IhDERqSOb3+XvXqwnyw/xsLGOeq/ZwZ0Y47Dx5+CAgSqN9Zf/qxrX1OsIL
s7PZgpSPofa9p+BeFR4/xlkXiZty1iPpXjosdDJ26AFZPgV5gRNwAnYYSzujNF8e
CFdqCtn0fJY+v3Zj8AlYsNttDyqwM+luYSOUO5hchRI2LyRq6f861ml/y6D/p6cP
RLIBbJ/2yQJx02yGn1h3/Y3am9soRsqgCM1xC7tlTfro8LKkIIR6kOGoYPywC85E
nxxQM0tQ7YDphuoAwE6RWWwi+aNi0kb73DP4sMTFs6dktUAcsWX9HYEQbYMll4pN
GiZLpZW8NSv5DFvox537cmFh8ZzLlyHv+N8mbHNJfkj3ki8rcyZ/ta91OfmpgG1T
U++Ama8QA/P2tFKoAhRDRhRKTkJ6aXEqlAesS9QfYCLhFCUqNjZywUDpGzWoV87U
zZPvzY5aNCABnS/rKxWgPxPB/GAPhxiKAOfwrNRewejSDgTZsYGZEkpb5vTxmfbj
6k9R1u6y/YW5iBa44TM45yJgDA3D22uXfaohyGlrnIMju8jiM3Cxr95yR8LI3Pei
CCe/Jq6xNFLyhauxJcv4547Mw2sdUsUQiPFyuKmzcf9zay6B427qvet+Y68hwuDX
MJZ30b8bJHJ6DuG50mYmkyXmXNBtiXkxaw7fXZQMCca4jnid/l8gQSkQvMYKvwjK
W0uoVDkJoHdqYLaplx0EYyYowzqVDnfqMq1aDC+clueFSKEwm2y929Nrycyau9Mg
yLizEW35ZU8ilrL/PzJ2DOP0CMHp3TnmfSJc4B5V8++lab355hjOPY7J7j3blzcM
vlERE1lBNCYI5i+JaT2PsGnLDrTz/dFoC1CAhhS/iTQiC7xfj33gEYhB7zr1Bvyh
Ezfir0gB2Nl971QWgR4XZLHtRCgSm37Y1y+7mzznYE3xevx2zTffi6S71x5664xR
1yRleoydxnGjWvGpQFKeBXaUgEmU2BcErKyo2KoecyT/eOagWYnsj1YRw8azoHE9
6GiCfh50CCKRrwX7KFbMrSR8itckOTDMwEnEerHHaAco4fFVVP6iKKBGRY5qbgqh
vPhbwcVq1jynPKLWLd4WVBqkHGNHw8Q8vGyN3uD9Tlmh60TNVtbHeoBPkynO2gUA
KFvQdrizVwX8EliGcXPtr1Durc8fDDPqRc87u++1Z4+hABx7rwnuu3/D3Nk6GG+o
XfCTr8RbFszimYMYw+cjcrA5Bl/a/2ERx/jCIml0hK/GwHosvbC7vM53FQOiGb2t
qedHGfouvFRB0jd+2j9oi9WrzskSi9PWLPPJd9QgE6XPkB5+lN2MbpgacBfRVq9p
jbEbnqMjo/hDP7JEMCl48YViKb3x+l+z1AhtbuE+yO0uFPeee+oprLFo2nNW9m/4
GZf/BZ4T7VF9DTVE3r8thMeKrX100bZJHoV2pPNBcY/2JO8AIgxQYUhGj4kvgLqu
OfXI6yZn25daijVuHgSTimvP1xI3ZRcldGCumc7N2eQgCv3JNpZF+QAz65xtIgVL
U2kYSsA4zrJM2FxddsBW0WIvLe8R99AKbEYLp3MZf6CMWRR7C06Euy44ywawfUik
1/O/5jOQkdopPj1HF8zXXYWoFJ3Hc+VcjdzE5xJKTmwVICzPvDo4tyZK/txsAtxP
dKy+mbk5SI+DpXkcAeGV4/3W7XSxzEz6Y0Z+1J7aog8lXB3UmnfepbwSdflVI7XK
xENX7Q+Xfmz2s4vVi+WtWXwOUHW20OPK6D3lMvpyJTl75r+PwpfpucHOqDZpBZ8V
maSJUw1ZaEc/38QdaHEr29qjM1zOPYVrbZDHRa/GQ/jsoKc7i/Kgu42C0142VDYh
TAyQTUzk3BXMmduuqSY/VmqwV3yyth0irMMgTRCKT23B/dqDZf+k5xETFVD0y8HG
YyQ8waAlwfwnjOxMXVYktttZ6r1MeIqhVvzqRs8EyqSOiqVWBm+w52WVsAPBp/c2
4aYpUqYRz67FzPqFuvWwFeEqhFZMGWeShxLFObIcwhUiSFWHas003afE335/NNeC
G3Qznp/olg22BXbszaP9/GLWIAnj/0rgURQsNvN6AqQmV932nM99Z8nXo0dQKBS3
KcwFdenky3VQMEK6LdKaI17fLUWOvGc0eWTFQu5zYeNEWrVEMJr8BHWGLJ+4+t8x
yhUtJ9lFmm0MfP81WaIxkufo907oikpw/7EFA8szc8eHEyPD/CqKVlhIqppYmeVT
OQxKUwEZjLQhK3ArzlfQtlRgbKFLxm0CScEi7mC1cX4Iwq22Jrx6bAvDCugcV+gJ
5XSX02r/mVZR/UCJYRZC6CjYh3Z6Kcuz8HU74jV3u/6W7fClUlFCLV8QuzUuAk50
7JizUg0yS21qrJETjPtU4Q/pjoMbfObqDb00iYKo5HKm4ILgYwConCeC0mujkQU+
qKsYkRU8k0RiOBdntjPE3+k8OFAF1tqve1ePho3bc+Ka6CJ0Q7hK6iPbnrygvQnE
1LHReJ3a055otHT+bmD1AYb2UT4F7LzTXzo27QmlwLPSDwEcTymHr7Tkt31Zs+DN
9NzHgTvr31lfQRPx63eoImnsCIBvpc9k5Qw60oQoVf6MgdbssdeyW8N7v6GeC/BT
sc6Wlp6jmawL5UVGf7JsXj1Kv4bERTKqOynmWtbXUYSU9x6jcaUHAXHxqeAmSZx9
KTmeWJ5prfYV5pDSu5+nGXm3e8bRgkoWx65pH66P/85nPV3SBDShKZ8gY9XADnp4
+S5rcpwrtUv5aKacc58VaKO7KbOR2Pk0F7n6/vNRylKEF4AVTLnNJsoVpEka24L8
Dw6peuGgH3POsTsa1mzWhCqzhM9KuJbwbvVhJhEGQeJ0PN2+Tj8E5xennM63ey5S
QRAa91+V9loOJ1KPwS+Zh5A2SLJk+/IgU1O6UBZS/R0RhFvc7k1BjYy8WbGRhRKU
rQ2JAQcEu1oUer/p4unw7M/RDJYncbieVSV11iOvr7jNEYiN6FtdyIjFg9Aakn7/
B9Qc6BSzjLzGE1CXI6c7RJtUo/8e9AdXlua491cMoYNmhL/WA1DAQgCeiVsBbUs0
+STgxihLsz22PrbqXytWPnEZddXvsw87Kq8We/ZbHV1y35aSP9Xo/5ZLeidLUKyR
bQBXF5FZDKPrSojN7COdMO71dtmT3aGtZ2oYHcRq4CPEJLCO12+0v89vBo52KKvj
TDf3jWBJWgpu+dn0iUhnkiSOVo4hbmtC+GtC8Snis0TFXZWrJkBLFeJG3753+vR9
Rn9jC42iC4Es+TyJhw2/6Ta28t9fYRf5BkwAST47RbgpPssKvG51WxPMYOoVayLh
2KQy/goOA5PkZQ6JfaqCR3W0/peoT5yNseqohdHF2OZlqZ61hGhxeMMG8+S1L4XH
RssSQRc3lQgwMx9hUV1I/6iWW7ycLM2bhyJxF6L3ry2kiV8GIH5GB0DnZsInhgBC
HaMMdYBdTCm9WajRXHMrSbcMtLPxlMPKrhU/yVRJFbcPWfu4TqheKwhhvy3bFW1H
LPgGHGPhyMubxOHsHf6R6IcxM3Pzf5SG8zWdXunD7QwRDPLGTggYPXTcVpYjS8fr
OW8AsPz+M4wSyvlmYjZl/rxnSglQry6KWbqJ+JT+Z6InIK/QeGzmaiIm3FxzEBwz
PWiqADCTHOOG8/WT7LMRBcq+/uSn7GQt93Mtna6pGFMW2zEfW/+//BZv5PKsuHb7
sp7vRWiTrwZkce9l1woCuZOtSIuzvow4exHalNKGkJStegcZVvjuNVJq1Xwg44g5
6JkheO2e/fqjWHYojGuqv9yJBGsirHUr7m7wwivFjGmI3V04c3O+mv7ZePyttFuK
ias/sR57UWMXuFy5dDkavFNYSNxwuKzlnPfXD/SJmfJq2hDFBof0JBLsnkYV11h5
SeCfVC8nqgq+jaFVa97QnwkdlcIRb2j/+B3ydQ9TqMQ/GhIBHhMP4XoVRJcvCIOw
quO0lJIWYgutzcysawQEIy3B3C419pD7ML0FRHHMSoVG248pJ8s6xPbDO0J3+rTy
jJLnXfunTlr4bCdX26BaLblzg9VdQdhA+X1LHwkjjJrVTGWr34uaYq9GBpJDAb9G
lFykr7FKviVuEf5kPYIUJYU58Ti5XI7F+7X3noo/i026ZxlmrNtS8ZX1c//2Ppfx
218K2btieqBVl9Mxh/aGn8quf8PukZ2ig6Wh65+ahz8VIrGSILD26hgTluDh2ccB
XL45S6Z4zhf/MJ0zUFXPH48lzcB5raSSLw8QSQQkthfva4F6D3aR2DD6JfkjWVfI
CqQ+75SKXAerR3FaB6aACarJOQ5KFaLiuaoA1YDKoS7GSRVHlkwftQrptSKQYb1c
aoNPcvWoZULsyTH7wUl6z1pBsQvKKc6KENKHSPZuc45v7B6EMX4xv1Iqy7qzDK8a
DxspL70c4UOoW1b8RySeitOEaUjs0P4C+1Bfi5g0FE8greCVnQK2xEzX1X2OOl3K
GrUpV46bO7dq6+w80V8g9pJe5ar7qrlN4dEU4ll0jVHZHrSFpaCSzuHPP17LxlVf
67W7Wi8kUwlmPy7duh6QZWk2AndRU5Y1xzdTVrEd2KL1ExrFMQ9uauqb1c8Mb1Iy
fb9jQQyb90EzgC4hbHcON4j+bZsSJHYtpj+img7J5AcZMpRT7MU28zF9qi6Ks5/f
3HWQWckgTr4QoVWoHIEOjf2jgW9aZa7NRVvy7Oxt5shZoaD8jzu22YRJ6Qyl057N
5V6A5jnNHIy+xm2HD8HiwmrFC0/KKbAcWLJbbi+MKMMUs0xVkDdaKCLRAvOXxTRh
pfDkXBEQkmWq/IBrOxvC2QvStg3QvqS3BOjr8hl8k6BAmdaMne6q9TUxBXr4FrAI
qa7lh7sKcJ9WS/MpqA6xrzibvTsLuJYcKqYGk4MWvdClDMf+ZSMoj4o/8QEwaPU8
l9Y5/kmW/HkDTwGLwCYKAZWfrry/ZB7PZGkYEYkKOLboPRDhqwpfuj4tpHuHRMf7
jd9dTFFO+fXtjwhrvqy9iqril/vsicwk/lWSPlS0Lao07YsTUapKbVeY2TdP7YkF
Fw0zdXOP0PTEZsUu3Ck9EwpdlBmhy9KS5OElNZa9M/L/G/QGyGSUH2NmsuKHMVNS
5InnRY1aLVf0X7rOfTnAQ+0aibRdbBsTAcQRpWobs22WWguzKDJC4SCk80IB9nMH
b4btTVS6slxfpOGNe6ZPrANemKNWxpqCG6+2db4xYd7S/ht5x4UgZ3i53MahyXS3
Vk/fPd+0DoyRvjVCbInpHTh3w1lNg4tUvV6S8tYvklQHF++zG+8wq4nbBCjKjdaq
zCrAh5NWecGWBsSpq9klBdMRCPAYzJN652Y+wSnMil99HpKth2TUtFPFvw7i/TRb
qquibamT8r5opXYgrkgi2aPtyV55FiSUGFbESUVd9xgeQPgW6OvC3n47kT8Slwo9
zvrBjb1jXbXGpR2y9U+g3oLdcgz4z1mx/SgtDeP+IfgvZQe6MBycX1T4ALKpla14
1q3yk0C/8aXNblvsCiuITTKniYhfA2PAXJxetsN+xkOUlvuguJCI4B/9MqhV1591
g+W1pvUalH9gYUugmazjEbkq9TmpZ58cLOGMiCEC0tFALeGNUUbbnsKYPWhZ6iZt
Rs2XaF7g4L8A1RIKNjHoEnzhMkqjEJpAr85QCxl8Ysq/MIMAEO14Dqn1M0OxIL4L
4nNccPDs3jepCTqv54IUkPlcO73PrapIiU2WPlRunqSNq9DaHtwhTdAX6bPPV5Qy
8UoeAmg1sH8b5lYRb8hjpEBHjemK4dYchnG8CY9gBtUK5YvptTc03AdxUe5beHbK
VW0iASJHZktnbjHwa5gqB5GMEbdI+95+etJQEQQXI1zhxwN2yuHG/cbuePQAfRpP
vn45ggdoQ3BQ5+2FsNoZnpr+neIwkGfdVrKtibpSIFCC+oZixT+bpZ7GkmosKc87
Nrf02spotCRnowYALcwo7dLaT9ktM6k6rG1TuSeC79dLMibJ6+aQJOwphXyDfcOy
/7yZaPIiyHRiC+8uiXmBwXjQj5UkKUV64Sau8pOhi/n6etst8FIwZ0mqz6FT+KWu
5affgMXQpEYMPOrEWRqNIEb39O5q0PcpT/YffkWt1WmZbRhr1wyNmz6Il4GkzhFb
9TcmOXh4UG66FqwKuW780wKPTzDeFDMvL6uAP+pt+ZLqKJHeZQoL19d+AXPKQZdZ
5ogQ/bZqB10CwHUsyfKlzX7jUirNPExBuAFXlnMZyyOQytteSQfAetDUUOHh2HGr
zCRag4ogzniCW2uP3anxPTMVXE/uEQDg1s346Dk/3T3yEyGI+0+k6i4HfbWn0EEu
rTMSxWChoYLrBPjCq05furq0dBOfiCH058s+2NLNjwQGCT1IQO9rt3yeGm6hGjtK
0ighh4fbO6sKAokPYoAsiZTIIofG5QaSiNuIhde7bCUOJ1WgGWfh66rbNTVSscaj
7g/oY3pHNS/peGZY1669keTZ4Ea/1kJABMUi9tO5bPyJ4WjtKUe9rwqmPEOlfkCk
4INIGT8Wq+LqMWIIxDmGxjoQDWsuKAu+nSy1kBeckO/+4ctiuRJ8Gkx7ONQdeC+f
piDZ8qdXpGY5XTgW7d8QZnnQR7hOokQo0ENFsKBuflZxQ+YBzDn9b1eXuPHLb03i
I7+kSWUuVGAk7G2VUnxmi2iMhaiR4i0dTYCgXwSi+TzqQPDHOBnrtbReshAeYw8q
5QVnIzPEW760Quw1JH2WR5/N2hcy4U3Ro/cRyskVD0kqbSsjKJYpgXRG96RA/QQg
eLiB+j2j+5/EUiziA90/wpmufUuCTbvdPTsWS26CE593yApjfVyNjALx0E2wV3To
PXM7jNLt6uqRgCh4L/737k0Q+JOWPJvqD6wJoZP0v/0QEQAgzYQCNnI+t/rj++is
tlcHtY4vn0urW1icYB18Ac0yWMzjPO+XA2L+j1HhP1Fhh/XctPZeZTBibAmQs9sS
cswCP8ZUUAm8u4KD2J+jBsJgETEqpRlweI9E3k8lsJFiKP4VwcWjjz3UNqlDIxPr
khP7cY0r8Qnf0pdTdMMnwSQf5oIulWnf9h5yzkYK91o5/UoDDlGo9JO0xwmh2AyW
znp2O5eyLK2TBz5eHL6MlPfTfztL7x39czmlKKq4ZEFvK/cLtLmvmBNBtnhs1hlY
a9cGBZ5jvv4aXraARcSEBVH41Uw2EVChQsXjKWKcoghqPluuUwHxMgtU2J14S7rp
HcVp3jPbW4g3x2MS1KXFzu5KOB7WbJwucgm2dWjS1y5BX7AzDT1VAMRqP21IgR0l
K2sJMQOlcvu1B0AgxeY/LFCnKw3OlybHF2qwXhon8WhsGtq1Bb4NIv5JWx3xKwHf
7ClhmkLLv9/Cmf8pcIu3quYyDtG5UnTG9NPeru6q6wdH10IKZszmMWDBWypsz5lU
p5GOtefffZtPPnL+Y1kN7ffVs4uZWYxs5oxr5lgZjTj6paqdR826KD01HmsL2IGZ
hMqeMwCzl5+5iBIjvKflQu9QLNZyi3Zbld7vtEYct1sWI13dIhFWE7xytX2Pk+8+
IwQE60aSoc7wFiUZGDRICyNDuIr+1ixsVkJGz+CIcggnOOGwgQHnnM/ENVVBKf8x
y99LtKkvjV/kmih9FtcRjtOAxP1+oA0Ombim4NutuaUin8Y38RDj1sAQCTq5A10c
NTJkBis1sVC2dPsq62Mz1fEY0zGs1WoKMWcP0nAoa3UK99hv2+Zqk8tJ87G2vRS3
Ixi9DygBRoLDy1sjdNYvBPDuR944PUY8JDnAJ17KFM7v4Cnxps61+hGsucGwweei
cgoRTkhHI7J07l4YBEdj1KgrPeei2llm1tAft4QxaluW5DMcIdJ8q4+2CyA2Mixq
ir5HmfvALvhnrkBBKfh2LNtQu4hyUWSrhVX3WRr+hXmvKZT2xreMRPPduvqo5P4t
Ke8u1KBBN/wrcMjdDzXLoyVJdIn9TB2leR/pmFPQuyzFkn1RqoiWVcaJfbHzuSQB
+gmmlaWqjfC2MP843iwecphqin7M9KBLZl0Jfr6Yam54ZPLeBW5Z21ZQJeLLIkPH
2Brc+Gny067dNc9/QmvWaJzHw1PclzbeU/+tOHBTnrohPh9k+s5BydFROIoMF4LU
h17L4/GDS51M4PXVhaaYjjaH+CxFLIFW9MWqWxDpA+Szi+Th2ptW2HyB7oh7G37l
31EzwEN0BbLht91cfdGMA5xFzpQUjLLOggHb7o+ke8L+3uwK7vueTUvUCihgypOO
ee104P8/+48iI/MlVFyD4mzE1kjyVuIdGyO70ksl4opnUEsnSA6TOmFkziFuTOjK
6PcyXK7twFlNE5eX61AgW1qatbZT10KLjGNSHYmLFEn2AhhqTIf06h1+lJbji6l0
hHDktqJj7KZWcIQyslfmaEMBpnCNpWsVURBAHZbGyEeAu/9B8ZYbGelHEfe9Z2ip
iu5pHb0pd5jVGNiWdSmKSeHlxlVsjIrmVh0EAbulNeKgjNmWH6tuxWEDGbdl62z3
IpJY5mcidyrBnsordXoP0uH1Ue8CWoaxwBaoMPdPBSznwxB0Ebhu3kDcpgVFvQvP
3mw+2oXKgAjpRi2urEml8ZlkuopNA8panVcaEI/d4uFZaB7/fa3Dk2R2LwrdzPhw
zEKkWTiBx6yMN1bolG4Hnf1IDJIYamqd3r5XzfivHnVFLiN9Mzr1Qlnft7NHfBPi
5b21hRXi+363jNyoMV+LRIDSkBmxk1uq8xsozR+TJlFuqMWtfNAw0hgplAt5VrBA
F3MBJoF4wsmP8kM8sVvW0s5EV+YXXJjzBld21U1JiekonO2hSXyZB/EU0DUF32I9
fCFgd8mQj0pCfd1i45ZoVFnFGDhRH4p/Lrwv+qQt/GEiAbEYoKrlDIgqdGYcDncT
D5zCq6MNOzB+mrlCXrwiYy5A6XGwal1X3eXb29yeC/B3zgqKK5x8Ki76qhZyKo3v
8BkmSDycUqU/BY/5OuPFa+eydQ7+SShAQxOpJwBt5OknJiKxj5ZQU7GpNAMY9v4Y
R3p34a+ACz9MeyjU0xHB+7buAL75Leelzo3lt/MdXhYcHUN3YeiCFaAV2puJLFSc
zc8Z9fMMlSx7BONOuzmblGR5b3eKmPOYFZHctlcNgCnvXWYaSrF3uyKzZKLq7Esw
pcrSJV47L8RFhwstJJA0PoAa97Wkcu9FlF2og3GxTJI/9s4BAaTZ2f0hEspIz1Z8
jlQ9nAuLWKUMTdP+vfKucWlPyKPqdIgLyBY4qv7TTOCgLTcqGhNDtw6P0hBFA/2x
rBQZ5uWoyk39jkd6XqA5TkyWoQc1F+NZCva1p8ZkM+4=
`protect END_PROTECTED
