`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eMdOpjGpA2fpU6BZg+tJG1fYTcEHUOUq3A3N9unt3c2lIjTOtwsI5n6z8HMP5k7O
ERq1w9gZRqDIO+8mqAuTgnb7SWIX0owpDbomZCYUW46O4GBZ9Gu0/FXuBqAulEq0
IV4ypcW856JS041SIOElxI2ym3kZ7KptqhrlU302RNXgeb7gQLzZjMhImr8kN4/5
ntg9oVoKHWD6pW9DFvA8JHldN4SMZPZPBrBRWNetfNz2kR9doG3f2vLlD282PUKc
s4T4WN4/k5LS7lbxH95kapQX1XXyIlw6aUzqmHM8QeidtJ14HGwDVR1Ss/lT8mbB
/ljA7CknoN+GXfMYEHkYRIBDdvTSyJIc0J/R3wL5sR4MXFdT0kYerTnHH8L/iSyK
aZkAT4Tga/jkQTU0Uuux5z5TjGxNnW+DTMTXCA343cEMU3qzsCZlqUGZg23j96Nw
XvNteLUsnHIIQDzD+TbCZSoZs5DZQgIMX/pUkun510s=
`protect END_PROTECTED
