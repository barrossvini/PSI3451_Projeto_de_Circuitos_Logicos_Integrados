`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pb/lU1TjvTUdYZcY88GPjasHJOX5Y3QuteEEX/MINQEmxM6Olj4zTbY6dTuZrQEe
ZoBanw1wOHlKcQshWKeb468ZWc+a4hAe0eMdDH90iuMZQDBUxNyf8ml6QUiU4dis
X5KJRQNk1sxd6j41jQthKksppRg8fBsf0EVJLy74DKufRvP0DeLnprKqDHjhlwg0
zPadpvtTIiVfqS9oPvLadWQQOJDgsHfPA63TM5pwJBLPYUtUK8chTqf4GFj2svwh
M8b5iumkQK5WxWnJBxORqLGqC8k8JpyDYtxC+7UgIkaBNNQhohgOuIbs20DebFX9
1vbtZPOuckd/5m6L0GyGZoqbeAngARZJU7yqlcf6F1lLlusm8QFKumfBusgb2n4Z
Eh8eApVALBwT+r8MXCVDrhGgEi89rErvHk89FqxGcK4UaGfQGFOuLqP6d4btAhVs
ksVcO3sge5qqFY933vBRoQhQGNnVx9eSanQjvjqgBdUsZN6+Kk4Qyy9qmw5+s5WE
6LHKkyc4Ufhfm9pQxlYf1xqTj9i6RwBJ8YKIP0OupkNVngJxssLTM93OfeUJUfSa
P+STp1K0TNNnShVvIrKdDgotcbenudiTsYCrVpal5T/fUTHh3r/casI3OeH0Zz07
8QnAcV2Or0kIXknF/M1uzNg37s/McYKqJn5NnOtIEcPRAddtvcSJWsnFPoe/N2fh
KSf7LaCiNwcMWBxlUgc1BhMWOtQkda6v9L077aaoe9HxidYwOwdK5Dy8HsO4uP1h
`protect END_PROTECTED
