`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S4sAUWzgEDdFe0rT5LF02QFNq0k9yFpLJXHu+inPcizyjFNnGpw+SQai3GesMEXJ
GMoErSn8FU89lDGAdQB7TCOubhDUHn06ERD1pTp6ziazoORUdG/miwhcXENqbpbb
xMec23yhDqa5f+lg2MuaY2XXqLCT2emjZ72ep1ywv3ZF8PPlXaHMIPgCR2OFrGFX
RzKkm8MKogzTvPRX4Bn/v3u76uHgZP9pGmq3Vtfy7q3hwRPmGE2Fe7sLLmygCzQx
43nERxRkhSjqzy3R3zOf9h6MvTHgNUw6JWTf12OjIfYgmpie3tbXq7Au67Gl3OD6
zB4pZgAJ0EKAcLTtHRxFYlW0582z2mfgptERgBM1nOQnRbgwd2fuJqysABCE6uvJ
KFU3s4SfH4KbIorRBbyGrLz/kjMTHQ3bdIP4K02UeH/6v9O6PO46kPwPHnOQSRon
CMPJOEQ4VXZsc67H3hB4A36okcXvNe6f7n988VcnFGWUZKF91QWTdCgjC/Q3RUxd
QCOjJsLGI13aMUDC6hJe0ZFeJNv3NjpPg2L+2p0Bu5DOAVsR/TB0TBQAWvNzS/Yh
Dq+r9xyYXaAwtphte+nOgWPor7sUpRoDo89XJqdAUiW3AegD4XZRmzi3aoAoa4CC
0Zjw8y8jjGIap1OxwJ87rWOSet1cwfvknAivQYvlQ1jLy93BqllX57lzl7+5lLDF
i1+IL/eWfC1oIH3a+KL/FNPoVdSfHrBBpwGkGcyeuvb8cJd5vleEithWto2c2k+O
0ccL0ld0+EaN54tqNYjOugsQLfoV+ZQ9OPgvC4H6izgQudI8f0PdqTBjo7iPflwz
ii0lHNZni2fKSo439TXn6jBYq74BQtIfcH3ZUBhSzUQP4jqJwqDNAUzbYDE8KolI
OTa5A2GYpzeFCL/sR9zmYk6c58VkSISs6KNoKbnvFu3Edw06/pg8pdhi4iLeUJW7
1WD+NxevnJIExHKFaCASK4FWYZpQjTA/gxiPVXOtDyKE7BkEoQkz6vZdrv8fFPor
ZUlXDLPzFNoFIVaxdiaeSlBQfXECBt0cobiybknaueuSd6QlgN+fKwp/PHg+u/uo
n/bWWFnwASu3NfRGR4ie11IK/iGkq2suHrEYNnhRKiQIPPsW5aDCmJdpUo9HBFIH
k0kZUsUGGm6twiNmg/HhsBNb9eUnHEN73Wm3p6MuhBwQsfY02SpqKUezP5EDnyEJ
8ciE9q5WWEtsAOe867X1pmFd2CIk0GIZFkm99g5bi9St/oPXzaAIKYFzZKGdSyKe
WbVz+zeFuJjr21Ei7hEaEPJBS/c4IuN6yJU04kCgz99Rp06jITugOhUTWqapoqNY
t+5sAIHg8wWTUsI1P4rKgQpDOnEsIY7u1ka8d/bmhl6zV4JirrBkZMFM+CG7gwJK
+1l+GSAuEHu9Vz4Hi2A7p/PIKvOu/c0OZBabL1Q45YohxZjnBwPl5M5ZCPaJC3fZ
WlrPzciXf9h6eG+mx5W5j8Nq4bjVYvzLADUajl6w+mFxVrOj6yBZiGmThKZEP7dk
BtFnjv1ZH2u8OWPkJHe6tMReTQyF5BxEaKiqGCHj/ztujnjGyQDkP5QeeFXROpVR
uAerFaEonkWANmQBKYJi5bBDnFiOgWLuYnTrqsxqKPmpJUmYSwK+wMtTi8Rfknjp
wMB8N3wnAGywqzb4QEZeJBTuF0pmekZdoB7dHVJRCTK23RDPsoS+wovxwlJEPjkR
NKbNQQ0peUCJk7j5H6+0JNsC8oB65ySETmVg6vbMaWEr6KkrxjxmZL7ahQ49+2bi
EkpjUI3uWUtXT2ulg1YuHdOKFJGp8hozhi8NEr/Q4qmNrQxYxt+/QfEhlJweESKU
xpL0S8WLf1R9xuRHnKFXQuvk65aZ6tZdN//2fc98BOZwPhziAnf5f76I2BNyH9QZ
p8JAjBy7BRgNu6/CIDQVx7FRktIBJ9L0karro56wtdeXnco1qP9hRJuxPmAL80er
U6OIg4oFZ1DmOZ8Mgvj5jjgDAwKuzXo6m1IwgObH/V/6tCjBwBS22xbmy3DfI0qo
hHSWdD6kfPtnFbziGN0k7Q4JGtlqPDKI0BaSpUPI/iOxocPuYdSnsRnNm4sMtilq
I3UMUWKyIHrIbo38z47Qa7Y58fygqkq9RNVL4E+L2O0/fN+jkYhm0uW4TmUG5mqS
N3nZk2yj4Je3AGIRWvPEo79vzLcO5PqtepKJ4B7RoPWul8eR6Bi8SxpTXWnKIsoa
u11NymsxYqZj3I59TQEF8un1HcQktQMy+y8ZDTMAwYHHkbMVv6plGs49GgH7BNTo
GDzT65uCv9mQwvn5vUMxrKP4jvaAKfvC9XG8hb3BsvHd6Zjhnn6MCn/88eojulT4
1GmH88p6B7Hls/PmhaDyhK/IkgkGVKE8XZlAlDJDfCBe/CCMvl9E56zXOkcnWI3G
hX+x+PeQ/CHjPWCzCaMbsS1hFNsw2JgX9WvfihTYSbxLjCkR0+ylKDzwBNF8EjyT
Ki1WCZM5nXmgamLhHU30QcTB25P0woClNqdVhEtw6tD5FRn+mKxM7LKKNAgg3ZGk
glcTDVMILNNyv4R0ASeQbmdBH+3Jcl71mEwRcvK5LARtorz7rYsJs0x99HCq7Nw7
G16QfhjKSzLOb8eXnuQccs/FdxhHAfknYYXbeMiW5wsbjbvknZ2URE/kBVmMJk4y
aZDBoTDalAgEAW/B+G/n58RlL4l0WxS3uCSAqacfsR1NYse/B1yDDrs2LE5G1OLp
UCJEQXUE7HNFUMDiCfaxzJdzUdViTGuAmqAJW4zuQoWiHsSpfSQabRedXDz/lSia
VAAx4rBZKF3pv6qIyDRF0O+zG45QrD7Pb4UBtbVJxMcqQy34tstPBsbPoI2hkAI9
tvf+XNt1h9Mc715XvoTS2yGnZYT8IyrNaTQ2QLU/J3KzVXx4UiG4Yyih0dOiIvBb
xO8GulA1Ur1lQA3K1eXmwDVnlV/LCTrKLOXoqq7BILIkiq2NrXZFZFzyctGuiIyc
N3tAS++9mxxHF9/qgho63jsWcFP+9PtMr1LBlDRg1W9PdNdlTtxT7eC7tLofkhGt
Yd4ZdfEhs3Sap8QhyiuSm65A3VhllpeO3d4cihfaTiDkD6SKoAgfLI6dCpweR3KG
TcLUiJRzeMqimvjE6OkkVhuHbb6YAubP2Njas6RD3ARuEHyOuLD7aD9O8DhJcS0p
uHgtSIyFRG1NSz+MzbSyQVygmgnMmOwyv11YS3SZBNgVUAPYVzTTvT97U9zcALuZ
AvCQ6BhdHXKwykafLjKzXXMt9o2mwmqtJJDGeAg7oCoQTha6uBKHN5BunTEhRx9z
rD1NknVqy5G28ZgkdIhTOf12tFRbUC8Sc56XFWzZRty8keJXtKdH6LygRb9qHgu3
szVOO6jr2fMxH/kn8OKzhnYQQ40/ueQMBevKyihpkPcr7RMUto8Dg2EAmKSN9jz3
MEBhdp8Z0KCOBoV2Bxu7OO6k1Gk8g+Uq9vGouc6OCEYmxmUu3KxELjoK68AmCdUT
pEdI+ECxe6hQQyo/rUCQIGl4BoOzoUpAwqbjlpDgEVyrYioiRmBeX8a7GD2NMxp9
07iJ1u6AtzCkiHVdByqeMoQN2VsvRVVQzYO2UYOUdzmxbQQjvily2cicAM5kwhvI
6uThe1a5fZVAwDMfCRskeTo2WAoQt8jG2C00YAwhkseBTiv7pSO4CcV8Xj3WXrr4
BWA+oLMq/hM7gPuhGsaJm4kuSS15PFVCepunlWAkfHw0WbEMNQsSFHwpmNJ/7phN
BdMm5bothwpCLQeA6T/NLz/nxuzv53nNTPQz5+vSs8dK91ttvkI/9KEYi7WbxBeU
LVTSE84YRF9kMkR4239LqNuYJaYv7jCaNwSmO9vHykOpPtgU6SgfrWGZrovUBSEr
Nr93nL9lN7vtiNO6Qx4wPGJnhDEcSBd3xPDiTo7LzTzrL8kHMcMePGW6+lOyoRKD
TaoaxAF3wgHECZ4nEHETKBMVdOkaomvu8zzSZ2HGhzVu4c2WONaUEyOUuttQMyJO
f+j2kOQ0xjD9hNjyrVromF+wvOHkO78UnJG/iJOEVhYgTvyywsYn6GlO9p0bUH+L
jjPyw8UMWkKTzgZFQEFatg7s5XGav1GJFpYiQc1Wk/0Dl7/jQmZd/gFHk8AosXlc
qAuglwl9j7kP7wMDDEiStD7vIY4RXUpQUel3qwCRa68PfABZMVxfjVIZTCxVp2Oo
E48x+sbKoYIq8a+IUJPsee1WwlGMkBFJrcbpOELk4RqXfe3H7JdCeBCuTkFa7QzJ
BL2ns7ZPBnsbkSqjKFRB+aeDv88KKrbTApsd2q1eYoipGVtbSdGpaTGEGe6+RxUj
pKTIlL+tBkGNh60F7L8yS6uTKuOl5ODs6GjZEJu51AW3gsSyVzsAk9vYkQ9Vru2L
SfETHbK8fGZ7umLS/PIYLBG3no/gAOYAtPiVgHMwkqUzfM46UzTpgQmPigF/ooN4
slipELxsrFSDUzE2Ip3Vjm1xBhLHKTQu7y5zAupqop5mvrpcCclEAThWKUPZLGyG
fR6ZC++as08FeQi43X31BEGVp8Zza/+k2tx6KzPtCMza7lhVhwH9cKt3rzCprs+4
Dnny0LlkFsE5xfkRuqkxH8Ft9FxuPSxp1k+gTpT8XP+fAqld5N4i4NmGaCT3N9Nu
PnScTL70dFyieu+l8bkeIL6lXENYcTbNA7xrvB3lvY1AM5bvNY7v4kNYyxuqVRaX
pV7yuCdxrNw36k+1mxhyd0ZCxkAgnp8MIX70ZwirHlxNekE1Hzo2EDIYZ6LkKp6w
dB+eBMiyR4tffMw6Wxk7dlZ1C1Cr0IfS4fjIPVa9CHg6uOuM/D/J1tfsFIyroEAV
B4OkuRI//2inIOdX3W/0c1g8vxh2w5hLnVqSqxza6M7aPcbO01PrIMTETgTpI7O6
7hyNoTITKv6Gj1WP2ljXcy8IDPqQYrCmg041qwFoUq+m+dQy2+7WDLY23QPrKLd+
yP8aInyhZ7whsEDLKB0srd6LFToRVDdkLKKUMRMbpvjukWuepitmvJ7sCWKUyOIq
Dui/S2skdEvEM2UZrOEB6U8p0tr/5Tm0UoFqT+VAjYBOL+v6n/7NcOo8sOSiwlvY
Fo1IOZFSzudFjCGF/f1rt2O6YVa4o2h13Z/TY889nr6Av3jEQBofeWEZT/2PJKQt
2R5mx/fGtrWARYh194VYBnsvOvxNDlqvr6hl5AnUQ2AFLaJwlJCl20IJ/3ROsNaN
5UCygyEwbbksKSmo7cq8fWJh2dSvapP4/JiVMcSSM72fOXYNfaypIJXM4YmALbEo
Ii9VZ7qWBys8cdXmT+CIDEg/+6h1Yg4g2z7LSR14pAf4C7zEuGsx55O9Fi822F0k
H4L0JmP3WXQRrZfMmwTD8EG5QtKquP1SGHRDnpc1p77EYs1ShuIgi7MnPugUlK6t
I6aBDjR8jS9QuDJa6ZVhd1TviUhd6yirTKtjWATB5iHG72kizRIMsJb+IOE/TLLp
PLj1zi0efhYleHNWF/P47VcVYIIrq0s2JtZpn+mIn4dpDtRTuFyqeY+XjIGGr5Fc
23QnUxbWlQ85qsAY8DrqmfZV2vEQjaw1roscZ2S3ldkf/irfqMiQmRbQ5qUf5MHh
DsklLo+B//8C3Ar6RKY2QEmrcJnHldJ4peKd2raoWCh3chxdpjek/7xfIcmC3Pqr
5dfjovYlcxVi9/i8VbvUeeaaQkHAOsayH4nNkThMhE1IJqqQP0vdHmfrjQv+i53W
X2bPuMGLBDDKpySXpZiaycDYHVPCf1TGTBDnliXCnhDa2YshbYacecZaA8/odvEW
x+uPY4Hk7d8XdLx4tBJBP2DC78HIopNDEcj//2ylW4jqn+g71yP2D8IuXvB4riH5
9EwIgT3awjihxWHByCJTmMxBriF64ghrk34cz+mDkha2p/TCEGf4EvoNp4pTYeXW
7Zy+T99+Mo8P2/NN4XkHxcRU2vgJZpy9XPWD5CTOsYCCqQitSsXLXwElWj6DUs5d
ozKyWnUGpJpelknvxUsPwHgddUJredXkqkFDM8o0NabQLr2BO9IcnObS3Hy2W4LK
WPM85pu2vW7fqONK5EkJjJNeR873MfoQz+jI1MtpqiOX7848EIMUvPmw/zG9n7DX
KKA0G7E4R+U/Omna2nWJsAM/cIC79hS2Py7xSuY0e3Z/7XIyv2PwsPaAZUweCB1o
2QO67ygQEJSV3BUVPSp9fhRtxgaqYIiL0jANYFQFMsv4b2x+XEy6YOzHhaaT2iPw
Ouwk8hfrNfrscF3m1t1CzlV4ZjFEvvWhnIIz7mLSgvbd+5eerblodLraeG9vzJsK
EOPVMJQkk6QOT9pcWGa26x1mYufHBJqh/BCWPck91d1sLyWAJpLA09P4LX/K+P+G
7h4j9SvtuJ1E46zSgJWVGtwSbklq10kWZ7EjZv2zu+C6WxQaj7vk5gERd1MBdUKV
1AOhjpAN9mr2ZSseLJOP88AcTaHTzNAbox1ghBYvyXnTbdFZKVvs7LgNNhwdPcsl
om5uPumbna80v54ANrclgVQ0EolKqPS8y4Yqzt/rba06HVznhisiVThSLUYgBqRS
hoZfGx6PoqqguXVean3Br2oy42Xv3movUKqoQom8fs+C+hZnSKWm7URRx0qLDw7R
cV4HbSTow3cePaPbfrM6b8KjuAVqCCgviD7nffyCkXp+C2DwHisanl8yaB+GPkig
7GoruPTOAv4i7P/H+G4l9HUY2yF+UI4mTL7tToKXsn87beQgHJsG/Jma2y5pXO0q
6fCbL/pJXcMUX2i+LkOtWGHdHFtW+DPcMKDnDADXUflEmKBA3TdN3cM78zPUyHC0
zllXRF44KcBHoZMcGFAOBPjPrINg1oumfh/q6AMAYL4/1QcRpxmUJAe+cYcbNhAH
cbkliJk1pDOOklDSSK1LaPBneswNQoUUEiPnH869brgaExXP0k/aJm1OMnfbqGJl
SFRWSLN405N9cVcGirFOQoCqqug63RtseIVTmTGY8C64l1VKuaQqAU2sB8cAw5C5
ZuKgzSFNhb44u/Y9BhzUCpxFIisL+AtHWMK5ziuoNVnshIwyE/wGbovEDOrmC7F2
QMXoDB7zGSr/Ewt2m9cnWFcD6yuF9KyDDf5G+SKU1AP3WaCT81Afx8ug65XlA3mi
i5Hzi3/ctzCJe43WvdNFlRISeLGIHre0wikl+OduBCwjI355wxSurEvIjSfuZRJE
6tvd+PHK99qNYYjihYKc/vibRhIgiZPMow7yolwA6nRerr/v6ILp3XiFCfPvqCi0
HABvPaLR4i7swXeso0Qz/ZHzzOD/rpM9aQk5BU6YcDzSgKgFjp0BPjal0CRt1ubj
DDLt5Qbii2wuUjVowD1idi1BTWxhkpr9ZPtDLJA1S7G1N0rABW2BmVmfCiYYYxvp
qo+qFW0dVeaZLH/a6P+RX31JukDVC7TGfdNfU1eODrLF1Bn9uoC6vTYHfDMMJ9Sq
X+AvCdE2zwbZfNpfM1NXPSqk8hTq82Ek0Yl1378r3pKQiqMByMQJXps5H1BF3fP9
PII2/jeFQQMPu8ErXa70lwVFPVs3JEWr8YOLL+bALjAj602/g/yiUjRp0mYYPK+2
IBTObypk2EGh7nURprIQ+qyphwqAyclO2rnQ9CEKLDG8uvKf6RWNY3KgkJK0LjyK
mpzoKtBfC7z8DBg/ygoHr/KvZy0Xds18LTRD1VHowf3bGyuqLspYVuj8sBDI4kCC
o/k2k2ahw8C2DtUtxuNhxts1aSEXI13j926fV4r0urQE5atMOcmaJB1qOiPHZFmS
6QHV2Cf8igzZmX/WatADN8AT75xzWN6tmnN7A7lBZrXjx9+zmdwBiabvyWY7/Z0X
b1MMu3Z6ejRQaJrm+qMhheoK+E42uaPFsFeDDAng8HVlV74RIZg9ywCUItvvKBJz
S1dUUf2IZ1r5njAdjH4GG8qwOX5xwwNp1C1aeKcvi0tN+6tMl2E4lB8ONzdxj9IV
n3uRuyI2DAOXVQCepFi9NC7SKseHzomDfXbiXVMswgddfWiynjSF9vXEnxNOWiBr
hO/OVlqwZiwivLVhBoFCxnOafAueWfA2MY3fwSixEPwUSDb2ldiyq8IGLkPdITxw
TNyyUIxpaYYT+XIYX3zqKm2XbwU2Z5H/doqPUDT/+9Pf3VPc9Ya7/eS0xaKxkDpV
x0gLj4RAB4T8GQ78/GCxRHmU9ttBa/Q7EcHtIUBk4e42Hd3y5JMjJ0yJ04+3QVU+
fJTqulofAXGh71qCLmrK//cybV7e1xgeGLmdJkua2BN6hvp71zoL8c4FHOshEcso
i20TydHRi0KdDW4nar3p7LHdO1hzXx0Zu5Y5FJjWmJuHct2X2bW9GdZ2XIgjKKZw
gZ3StorUL37JKwsfdkv6VcQqqZE7td3+eAZAx1psl7XMRnxngrBuTjGd/8MrCfM4
DoaQrAHchKErHdX6OVC39kXEXoLXdm2pBV/aLJzAtfUSQyFnaT+gxGjn8uj93lnG
O054Mf+14+P+EZZvHaktZeV9EbfTDhJRDc+t0PPmE0m/rbBsdpZQ8B8HG254mAZ/
3n6cl3JEy8WcvOqYIS/nbwddjFyvgJJsryZ4Z/LaUl8LSjKZ7h+I03Z9sZA93BJo
33dThwh3oZxERZd/TcQve1i9Q2hkHjPPeRMsUgIjN9v0a07z8XW+WfDiBWvo6pcv
YPC/t/nmNkJGhkxhePsGON01ceryC6UqkJDjCFWMEH5dV+mHL5r2doqIwvWX/AZd
/wDcK194RM0C4VFoQmFfeTIaTkimm+BniA9PpRTZI6Odq9z52AAMlbyVazHPutpk
Ce0KERCMQiithEVA5IuHMj7pPDd3QRFwiRq1LyYT5775IDObGkj3NZRXjENDXscf
gd9z+wNMS3TfvrOOmIzv8iqdiALECAq3IPRRUqY60K6Y7++bnEmMzASP1xEqQqD6
wW3lJNJexr1px54GU+3dQSMlp/i/MHvhjsPXdPshUNEziZ/W5XKkfA6D0LY/Qh7t
GT4v3TCJk4DfZ7DsXOOML/XAMYm8oJiJVmuKK7P5iLLwQ7OVXgDB4TBUx7IDh2wo
l4ShW4Py2sDAKms+G0z8x/FMmyEcTchaMs/9Z1pTYjQLa3NibZt3CXVaYJhVWxLC
v0zv1fTtcg7IT6t/KVbreQl1xUsQnVvOsFeiWsdSpiXwGxsarwcvVfWn3FZuDjmI
R0FMCzMIX1dZnAVzlm7Gi2kIQWMEAfIMgwx+iwJUZmJF7yF4JryXqIsVNm7pfOpa
2D5za1+U86eBBjBiWs0Lg9jZKN+1tkKonD0UsCVFHe2xYIgq/3CYAyxm1Vh7qlyh
3neu1y4JZROBPEqxEvDeW0VSCpsLts5li+bcpvvCSY3SwdxDSSD6OR9UI54Hl62l
nzPQMq2tqk/SbXDw+VOisJLgCaiG22LGh74Dn5oUqHqEg4CyQaYyMfeQylDXbZr5
C5BMn998I8PaM1f6aqrQFs5GwHUOnIJzuQIEJZMjLarEkfroUsRxAX3wsRNUuLlV
fITqk8a/7jz7g0kT8rjDa1eD4FhU+ULjbsXYbj6+LNpkYDZlDQ+olnH4Bp/GNcNa
SrSsriXUdcoeRm4i1IerwTFwIzpRsLIDLC7WgYmPglFJxPKtHMOu8AEOLfCwft73
HiDS/3g+CX5khWS5TOly60wR93mzJomQbopzUhpe9xm/muwf54J23QUDsJmkF0Yo
/qXmlwqRh6y+XaWQuR6bLTb34QyNsaSKBk8nkHkT12hQWTjrLwcXZrerqEj9Ki47
l+2iImmuL+h1h4uxvZZ4K6VSs+OoQ8WryxHMWfLezooJHnhe8vEGRJHjUOqWXnXj
8o1n/k9yVADaEBVmLAYFkt3lTQHmPFboFioa2XKIIRkldqV4qrZxoX0C0w2pZzM4
J/SHT5uB3fnAd8/s8AT4Vd0PMcbttVGiFnHeozZE0QU+Hp779T+6rt17q/uKKXMz
AD342gVShvD7egk3Jew8Hbz/WSGtGptka6MVieeSdEdSIOkJXGLzj1AKbT5H20ln
bN81/RCImB+rgHcT61ZKDqstEtXTxD2ZNediRF5qKAisXYT2cPAwY7vD5lY2FZCH
fTnnjcZjd5GoVCbP5EfDIDu5/J8W/WWaIRkIHAC0hIzAjW9JemcRTkfUN8pkVOX6
DTSjhSSpskFJYl58RpoN8UTlooQnGz9wBDUooqrfw9WWUO/kbhmC3oMJV1KIYW8r
85SUsdAK/oCttYkBUBjq95gOa8TgJaaOZ79vF72PwapTuVf+JiMnq+2ww3KRmHBa
3zzRgJkWeqU4k9MwjmxdD72W1qfGNNx23g5KYWaN+OGxImrmri63vNPd+Z+394E2
s6OUjF/lTI1Me403MwfBz5JfOvUswwoY21p0BSvBA2pp4aUzhRXixjS7+Rw+hKtV
MbO2RCbKO85D1zFER32dLfO0pZyByJ4WivY3FWiwLhtK8WZEURx5vAvto1qdR934
2B3CBFwjme/dyDL1ICCDCngBtObePJRyTEiVLJvj05YSPuEOwOf2Nye0CzGfQFVN
Ot6ixdGMsqGIhurFmxKoDyo/d6pLQ9Vixsa8Ra5epvaoruHkGKGRPiV17b76t+Sj
KjaCHjc1tfbo9u0i8KYM8BKSFmfF0d36PZ/hgbLaB/738rWeaG11fpsaW/12kKou
Am9p+EfVe+zFNejhtgVzTPZMg2GdlL8UVknVjC/UBgcwFZXznstod9830yS1bLif
SjaVD5sH1JayOxD8wm7NpbA6Dp5doINtC8g+RlUnjFriomp0MntNpj7BWqWfceWF
pJODF4OuTp03k7IIsAg/F+eQ95Ggioc2JgaTaNIovSdC7DJlcwDSY3m9Ea7m0/AP
Q3ySulXSS1P7VIpb1X4tNnId0bRBYzky3ulY2iRphPhRfrz9N0FREcjnemqJT2rw
1+p+mLncJllgYmQ/2H8/jEa3lJBFnEJesM1Nvy15anm4OQcTAFDuUAVdOXTHPbJw
uEWg4w/JT79AQ2u/TEu94N6tC3WTZjidmK0BNo0LWLN7+YNGexqV6kZjAZyapEMU
dWXFaY2ERX0Zzpxe1QGhUhvulZqiZNQi+XocYqKpjrRqkHp5xSNpEL2JLZqnKD8d
qzd1zoPbs4GV852FbmqSOSaaa52cF6/pezZEMhvO6ohXIBX2L+n4i0jmvocPqHq4
2Z8exaO6TC4wrQeEzVCgptMOokWgY7erm1EBXvrMEG0OxH0lXrXHXH+Vho72jUxt
enm59AZwMO7YRrL6naD7gVHRcKGRhOjUl0VJbhKCvGuFWgAl8GXYIOxF3D9qQOfJ
Mp8UT8XVlI37Vt4mVtda0ZYc7YdMdIjJhwYGN1sNVU0yzZharrZWIZJtyseGSgHV
U9VtageMyVRIUO1zx3H4A/Mw/WHnsz2u3wJxioq3Kp9sTczHgWb9EBo/fN1zNGv3
YsCmYskwOMHb/s35ZuJGQ0V6kLLL23say2ysQdT4gQ8+0JlwdiZ1WdZdt4IjCXDU
DIwd+TrbDNybVv6vje5QVeJQC7a+LQ4gTI6+9Gx3FA20WeVXotJyZllorF7OawWg
+4TsWXUrkqs53pVEP7BN55xY75dyafMMpiLSn3EvL05RKRRr5GawQbA/5AuLbPmd
ZGgbf+nLleL8vipNGbFFbzFmGKRwkwoJ0wJiQ0IcwixB6fhY28+ug3zH5oJy+cab
A3miLo4B9BWmowy4cZX1V1pqBKhgDVs1Dc3dnrJqI5vnSPnbGCy74yJ9Wh23LSAZ
fPmMsHfoRf5KUX4nhABC5XINBVknEe/3kpZK8/dGD0eYKqw00hz7AtMtFNTHUS0v
qX/qrYEqEnPUlljPckZ5jaFY0wrFMd9ZWtcWOHrGMPUxkdS9nuECKQQt+nAClcyr
WFewR0ybxYTkGvrmEceDdNgo5i4J/oJOkghwMaaVb2QD9+Bze/jGI52Egjq+Y7+6
rxVtuC1ygPcmMdcLCPwjTRtr0D63xX0mn50sYt0H+WqLwNF3kjADab9EtWqgGkPZ
LYzLmTRzycObItZd5gVZU/WfUkgKJiqm/CbVH/plskVZwGm9VsYZ7NaAoCOuTg3O
zDNNYQP5LLShqo53oaU58njiDIrXtucadRCaVwr9COq1g4TEHav6DJnv94FiPv4L
4yolnSNyd5V6zGvzuUFTJ1F2gP3Veu4OWNmSm4OB5ZvuoLE2KHpf3iBuEY5EveAi
Os7ZNiNFk0borFIOWJG/snYxA0/MbtQlKRNYlyV4A/MyZUR+93raEirFA6l2cjVA
4bdK6ZJWbFbshXqnVnOLWQ37TRdhxSFTaIPiEftdVm8ru4dtsqRzGJri2oEuxZLP
gdYWtRKUN7/3lbR4oVG23Wd7gqg3blztUBVXdEs1TSJdzoHGxw8zG343xYMVL6Rb
p8gdTMgG238SgztfzV5q9gZePZoJIiEvGFl4UdZODY65M134/IZGeJwMo4szDGEq
Bb/KCLCTQM5CdrZS2TrdwloNGQVhe0DGWIqUi/12GI041F1rSbvbrsXdkdklJsCk
LqCtsrvG7pHnyiBD+0YamiOsxgLVYqbl33Fkqi6Dy7FHsRjKkiC2sYaVfKymBPEr
giDsGChs94ohQfX1LSwQhl8xSgYOWADwLISotW5VQpFB/Azo5uWvi/RvWzIHeuFF
87DtdEG35LZug2OB9kZsaSQp3t9n1EBS76HW4/FsjbJcHoHMKhEqi9VD6HcNZc2M
OJgFm5IdAq3UT+O3MvcjHb0ko7jyXkhUoNTWUUqHPfuIB3V/CRaWSDsVfuLoWf1K
K842GQmHjINfWn195ThAD0UNuTzIxEehEU0AX4bwdT6L6dYC1CbGZG0Jdjgq14cb
O0WwHtRPh7sSsN77nyc2jkgCUKQA892onmo6HLEJ+NnpJ/b8i5J7/hEna7hnoY/K
fQIqo3xYmTEXwCDiLP1B1peKLLsRE1KSQKKIvJvfWyxKmLmhhg9bZLwDTfdPSqEo
fGjGjPXxMxW/jEz5dHlD+UhoGgx7WKkHLcIL5GgJHgh2uYh2u3dYUNC7kfCdEh0m
Qi1QdWRuLwKZrh4JU6xc/g9rg9M5Lf0aBvap4qVmKwIIFz/KIC++K1FMRtb9mu8H
gINm0/nCeXw8R5JmYCfsef31RHEeq7+lcv2MYL5mY/AVCjbrjP9zmYXOAps5IySP
8Et441KAhyaKLiNZLCUs1wXOEn3WISTCHpuCNT25BwUTAaKIOY4Cj2KN8JDPVkhi
BpDWjJfW1i/LZSnQc6StVTRS7OomTTVop1a5ar9v+gs2hqgFoH4KEjdc241HESy/
RW82vZjM56Xou/3DjdKvRkTLTNdusrCy1ep6XM/oaYJRWvq5Kp4/uzcXyms2nlJU
V/gzYP76Yvoe/q7pvquJG1YiZZiSBiE172PqrWVi/G6470/55nqOAD88u9WrVuCF
hBcBv3pUqbrGbX0r3DswXyp9RYi0lggYo2b3xtkEHoVA1sGumNwu6ro9A7E9oJZ5
wRF6CimxH0+aTtwSDF6SZiTnJRDqjtdkXjYXx86owXoTpB4jtAycv7e+29LvW4L9
DGs/EXR825k910oTa8SCmPT1vFC4mqJLQA7xzdp3KP+L6JLDynJSMrCXIlNIlUzG
ptRiqB8e5UQXFVbfNeHQlT/CayUgvrQe9j3u18BnWzOf31qFybmu0UHbMPzkeFKh
49bFsl+fNM/rcZeYUQNPxV12vPFYR94e7/VdsQh5sh1AcOluDgcQsLTQOwWCyJgu
9EozVqWUO9COdJWil3TKhdB4zeHIPoh1uEwgVFNWmXqFuDFdQDxXPGfzD6xQkLBS
+Jhm46w/nni0vAwrZyi83TDr3Fqr/qbmn/EffbDuO0udYouiWiGth4CWjUeCl4J6
K4wvIiWSXTALh8pamBLiSDcthGigc360jYSwpn61Pg0VZAJhdL7q7cgmUXkaALyj
7DOJPLfW6N4V9CHhV+PS7eUHxkVhzQxEJ1wUDW6BXxfEX6oCC8DqtArVLGgHRi8v
53agNcnRHShXwBvNQVO0nJYuKJ/jB+8AiQ/WsZBBs6rmGHTwhKy9HddokFWR+ttA
/Gfv7GfwvrwLeiyr7Mhh28GFUyxQd5l9ijX7CUyGp02MnJ3fq7EqRM3fqrQLrWaj
zxnNCb9RMP/eUKz3xV+IGz5hjM84cSYiIEQrUGAwIJKD7KPsBd1eiAeazcam+Ylh
iGBgeNCl42rEQEmXTlIIwoZYLniKzy2URF5cun8u3E9x7kd4MOQdNuy+bpelMnFQ
Cu3PrRb/gaJwrkxd8HYHPnuUyX7HxxOLDEEpCxBsCrvMFkcJz/qGqavY8ThLTHeW
xNTxp8lb0pRXqL+eKXL9nKH9VgUHEA+yAjMxxlNCHcRZKM4VTcAp+gTeTmF3Bb8c
k+FDLsKhwxgR90FaGwksPpMaNsfGa9yUzHnsHuwgrzC6Um4wGz9gwnDDR2sy2bTg
QAbkcBPozlWgPl2e+tJkug0juVXMEHSKI5BLsW3oOK/5qcIrOXs+Yd2zrwxrJ2Eb
GRqGUL+ldhIDumLkp0hwP9OJYS8PS60IdPmCAdDnn9tpjpSlVSO4UXcCk4j1ZXnw
KejPsa5GJ6M+cENtJHXDunVEAyoFcAx7phBkLhLTfLGgCvpSnKzb8Zw2xgQ+m8CQ
anPIOsxnxSK8q9AIQhCd7PgtmhRplNuaSzW+B2InSJPvmq79ixCXeA/AHluP9ABW
dK08cVdHBdQ33T3rIs6HyPK7LZd/o87XPY/bFqzztLi10wN28bw3iFeflRnfO2FY
GEE2633LlKKO9DR/oSBJaovY3W0Qj8RyJg13s8YsgkDlEbww0e2VXwSCIMMEW1ZB
fCIg66djmfuyIxwnE08VrrZHxUWUGtaRfyOOGAUiKWrhrkHus7cqWOk9FlpDsmGe
IdMtY9YLuwna2G+pYhbLC3sQyYaWryUDEm0K963EUQaiMVBPIEvWfflb3eB/oXBS
QIVPW4XKGBPiaKfgEPlFQgnZHfo017jKmRwRJ3EyCu56Wka6lkbBHw8fmeur5IQP
MmWS+FsJ659ak/Vt5D6PyEmElCPsidHdeMVNctS9YZlEsuVIvRwSeVcVQus5LnUQ
ggZ3FTqD9789U7hmBcDaWDB6dyE5hXAltCldOywZAEtt9wXCuPnD6xFcSg2Gif56
l/6294WDyu8tiKO716dEPnPu8+2ZfRtdRo9YvLig1CLs5l8ecQivZieWb8Mom3jn
JKLCW0kDT4r4qAZu6DR+6o6F0SgW/w/I9HCPIGn3Ozf2VpjI7anvkvtbV+nlw5mZ
GeiOj9uSzs1lLpWF5kStilrKPQJHe1t1xrh57B+HrlpIsaVLl16D1x0fCx4ZH624
xpnvg5YoZNyCMyDH3x4t6LKhA1iGw0pAqbBUQuijpQiisiX4+LCWfkPH4X1i3rhP
W1EWbhm8QQxPIRA+nL3IGJ5dci4LS9SqFtuxLzK0qZOPHhGKe126VqekV9Wj8bJ+
1urat86EOAPW9ARm9OdN5T1K3w5K1yHljKfKBKtN46CiOfI093/+8XkpIT9YAlO4
K2P8gpDEDzw5yrBf4soKGTAScu4rY8aC0a1TGWkJbWYPhqUlAtFpNgjOD37Lqsbf
IdIjiLk3XEQ9MCWFxqgvfTJxA4upbfvpFuMxlwIaYlninbH9o6WL9kUmZ5+xVg5Z
x+YRJhu72+wUJk97FaBkOM8Lg3+pJ0NTScRW8aMKF5W8qWllOKx6JR9vhxMSYcF1
XYisxs1xVVtIAXdYy3Tovo+b6KfO+8ikvY5zVBTuGwaKDpb85BKORblZMQldLFyb
fnABPkGvxzj73b9oZTHAEVytCjRBkJR+c6VF1IJjouOO82+Ks31EM/pt82xLCHsJ
itsWKatBG+ujoGAmSGH/acOVHGnXW56b/40H4fHHnPXzjqJHSlm4BMMcA9A/Bnkl
YXMGZVJmUxaoQK42TdZN73SCnm4f9cfHaaAjGblGE9MRL1JYsxZCzszgZZJZQnWU
vbn77bv0Z9M3eQiXtdhE1gfOmM0UyFb4/enXpnfHoXhd+73PZNwcjv4Ct2MReMo3
srsPVv+TcDKx+w9wjocaBKBdZTxT7eS2R+2WKjPTWfEZh01b8EFYVybMcbOAAydv
XknoFriF7dFFtGQ/pURpmyyX+nyUrj/ExN07OjRpnByfAr4k5mA1tF1+A6H6dH9t
T6sL1vE4VYPRWJjB9jDIw/Kg8JKOAnGLTEN+ATLZLrNdK4ZYh+IjEb5XREaCmP7L
6G+6B9bMhYL3slpDlXklQA8FR0XfJZO7s584YV9Oh64vn/G5KCIHGmXeHO10ZKkB
mqBzXpwaJAC4l6fUcu5sNuZXYHQ2pnr+KVrR6+TKILGzcPl6wN5U3vcA7jU8M9Fc
KoplPBfxkRgHmYU5MshlbnxMNS2nC6zypIW8QSKE6gVwHXsiS486Z9JqHkh6hw95
nJstEy9aGbpNXfgojgdz0KGazJaEWsS7JJF5wPKJloXRMdfYlWov97jheVGSEBmD
XCzhTpMfrRGDx6vy3/60xHTLpnAYhYet2/ihz/IvZaHN6ll7D8JcslEeOTLnOjBa
sQ7XsivDSCIaSyxSc6IXzakQFaxgLnbhn8FmUJkUY5ItUhijcv4Yn5D8dKd5EKHa
9xwhZO7LDoMJdcQVqKxxNfoXrwZPqTk7QELhb/vfUMAh+WpCUQECbigh112JaHQm
QPTPMVobCX0eGy+J9+jnIZfqWxgttDOuXZyALUnbNCtMSh58Uc5ffhVqlBvbsRmU
03uf8yX9YYQepEJ9NpcDeUyr41v3KUwo3BgRK76DIYLxsheonKKfAh3dr7iyMX/m
hsAgiB6wB5ZCBhlyF+1ZvSHlLTk0WVVHzN+WcHQvf6c3wp2tizoX7KcttnWNXBFJ
2SvigTltMRByqDYyUpv6Hnnur+IQ6ps2TQ1DL+4YGfqFgJQ2oI7H6CZlkRvZX3gt
CgRMasGEHBHimCdev7MnTRBP8hrJlvvXp9j9v+Ad+wIX4xVGxqTthNSVF2v253m1
JcemTZEYUD/fDEuyTDhglTaHhRp0EcNCGK+jEcusCI4gUHQOUki3VKCUpK5Wc4LG
DM1/ZQszU3VXlv9NJXtqFqR3zwqUrGseaCSyBDK/KcOUKcad4aZtx9oTmtDDY/ms
Qfh3ywRphAvLeR56SO/bW+f6eQxcwyjgE2aktzx5L6WrhF7naXiKLGQAbZlUZimz
sI5UKCUnchadKbGVjr0YXisJxqAdjf5A5TeHDsM/zSQL1x0wZZrw71DGkhra/Z0z
iMADrz7PVVnN2mzRQawXuUsuY+1dDhomLJvifwO4olustu8X/n0ymiMNg9sTSxbe
gfSI8mZw/rp2NvdXLqJMB7J1udZQDSg8+YAwwfBMQEeEIOmOUG+DpqpInjhv9l4j
xgsOxJ1dAI0PKl89rxpW2UNgvG6Gu2STgMOiZIgpaiinUerjcJjC6cChadoswwPh
a/+u4mejOYeE3fV8bFCrm170mTtEJ4POeD6sl69N+uwMFBnj5qtGK+qCBaPZflsB
eFoTA4cgcHKfv2CfI4gzjRh95dmrX/XvRgopZSsTDMZtPTZF7bb11hKPcoN5xHgL
6+KbMGUwcywyiY1ZVYoyTsCehEiOuVmZ4YicfZ0uN7dgq6o+0MqASogJGEXXKEXo
reizLBa8gPaxUDCmzTWA+zEFQJtKtQPZqkAtdpiz+v6KGhD8TW3I7ZCLnteqGWH4
GZC3FgLxbBAlPENgqdeEsEwVED8eX9v/jMKqr97zSS957LOuetmFz/KZIrXmf6Xr
otkaMeBuiAmzrQM9CwxBeJS1H2iQ3VNgjuF43uyrAXiX2JBny8yG8b1Tdf6JnwQ9
al8KyujkYmjAi7dKpXKr6XNpCj1nLgJyaNt8bM2c6hqTpxoKvdp2vLQwHB8Tcrmb
mLLLgsEVzajBV/zKC/tSsnKJtF3PTcppJ0yK1GaeBm4r+cUB9ex5q96xDLN6AHzq
DaTHFmTMGgzuLF25NBaq6643z/gnJ49S5yz3OgeXRkgqKW0fihvlBpBSl0l7QLoI
Ck2foCNEU26rxH9MWGk4pLCoP1pEF8u41Y1YI7fhFb48fShg6CoSn+J3c4FHJ3xO
BGbL8I3upcMbnUArIR8c9LHUNWu1zeazAcn5Jc2cQQDcaooSt7YR3KzWiZzRVrgv
ADeqgWgBKLsLqYXhu/R38nK48492Tosg2HuxSDVQfnlztyTmZ7v6t6hveHBdg7SI
alUyo0H6h3j0AvDmBH0wTwW+ComPHUkvl5j7zX20cEZo+568i6REPrF9gpItY5jk
Ub9ujlSWnwJ3OcG+3Q1YMDRpmD/fPybOieVJWdRkM/ZAOxzGd8V8H9pXnJvjZRMo
LZd6iVxSN40l3zOgdvYapoTjO9BA5ZN8TDhhOIXSyKKD0/OCfjZyzhCwMYo/iOn7
pmXB7RyWHN6NZmpdjved3w7Cg6LZ+fZh9XLSn60Euy1a9qNVYXlpzizceTQyki0X
hfWQxeS1c37aRrDNhuT+ETVsoXsULOStqjlIIHlIwNFwOqvX+V/vTwwbjmP5x1cr
BPyRXTw2Fu+noCi0qJz4PVTukM5XVy9Gz0neQ0mhHMMb+Xyb2eks/hnWuhhzCUJp
hjcJKSNr6fsJMSPMlmU/mZP8s3vXnhHwhrQ3kxpaZTb8uYAfTjSseqIz2KlhNHuG
iFg6XhnImdVENCW7oglCIZBgtS3co7IeSCvWx9VVL8xi89mVsk2WaABdsaECbvzD
OebQD5DcrU6wU8h+OnFy1aarPNYwDARaz3sooSc4/F2VLtA3Jw9c0xUE4GRSavNp
Btk83neMmf6j1NLFGfy9FYxHl4O66pzvqjEQR11ugJRPEmEz2Af7NcN61IX0ZA8Z
JZK6hE1PJbCNMMuQSN5VNrzhz7Gh7oVYojVa/Y0MGI2dZjNwGoRI/4irYBo7kw4R
lrtw55g++5d6868JmWvbekTwNvuES5TA9WyNPF/ujLNsdKiHTFYqt/04/iI8i9Xn
EtayRp2jPQiJnClsjGPcys3mOG4MoQ6Vz395NjT7HRL3jvKZtpwyEmW8q04T1ISm
esLp4mHIZ8jP4wr2cP4qBdQpQPsO03/uulTdE/Kiefy+jDsnYQJLDmkhopv6b0Dq
lq6R7Pf/IP00M3PupPkAlVo2rLAze/x2apO7k9EcrfZjRDyLACZOkoy4RHVKZiP/
uKd41srLlYuEW7jiMBIHOmzIQmfn/lH3LT+CX/qYs0uS8Jc3mAlpS0uLAf03nga/
n1OSdf3KaU4uL1BXsEADAuFyvweQCHOsgJM17y4THap1TOQtlTIgHdGtUtwbqa/n
PfnqqlVIjRuvA0TGVaDejDoZ5gYCMtq3Fm0zL0UkprC9xx+R+5EOV9qNE7G2bx5o
JTUdhxrSKf+7LqSmj7zb324VLuYzisQ2BqXPz4P5lFkqmBGHTUXQyFYBM2UZkMLL
u9NlkjYWiBNbV/v8ETanFXRnwi5ttGTFTrrea/RCNLkIKL3NlvFPUpFTVaAtreWY
xflXLlDiX1kp3eZgrfKqIGMVUdNUd+FsMAShsyRNcT20KbeTp2aAu6N8h8kBtNke
wanq4QmLj4zczjphTMK9him+/03HRMuRL/AvhHVW2DddyxqCLdT4VO6H8qSGfx2F
em/ZAGi8Lpn538II7R4H8ss3Ur7cu05AdUEeWmih5A4my9MHP83IZtwW5FqVnyWe
UcwP+rjpqgki5P0SiT25wwN7Tef1P9t3rRwA7KjdxmNMUn7gkHjpcLj6ak/anQaF
sVldgOeL9u92mdx4HkCfHWTyy14L90UIcgVvwL0VNvCk0s9O0aJmUb4aVfQUQm6n
sgrL5dGwm6kDiL4vhEsSPEnD0Lj+l8MSRYz4jYM99HyYV/Y+axoBaji5mgf5gSS6
R3ed9B/cfZmBBkE6usPAjpxDoPsfb010Xe852NgVi4g9c6e1VAVNndm+bULphI8W
gAM1NKJMGjlzqOrEz/KLbnql/Dqzn2RY1MsJsvQZuXTrg7hCaTVvt/n/b456viKH
YnsKFJ5X6lpmPtbRck0sav0MgHG98qzQ1VWxNfJwsket9gwF4S8zp8MilIh6l+u5
qyY96XvRvvpKXbrwBYgfr7FH1pzuMHsI+RQXlSUNKOTOADbwisvwWeobMZCPwGkW
XHBakaDSKI5e/jWf7YqzB7AMfxT9ZkaZUpKteEyHrAWsmh6PP/ImRv01Jal8il5V
17ML5trVzRJCp+N7edBXsZWc2ds8Br8M1bC6nZBrIClNbFx1Ip++tSg7STLL6Wzm
+x8sJ7gwWmIK7r3bsxCAx/nRAo190LIDSSwYjvDRb4RQGrGlKFT6d3yGj0TX2y9m
TfuaPZLkFaPofwd3gH0+ugCeLFs8I0z1N7vZfiRzc47toA49VWMRLwWOcKvx8+Jv
GhR8e1tcUWM0OA9SEA4oLENX1IJCDuQFXDlhHBODkqarSoUG0fnQJ5NGMaocQFWE
L641VQRbI+WfwXTb8lUrZ+Jon/ZoqHQWYdVWKt9+l3li1NxAgD+yKCFpD7A+yi3o
rvsg7IPN2vam+NyMlxLg7gUKAxgML/m5AwGa2inHsQHiV1089tXcrIW6QntpRL70
S4rwa+oUhQVWgavvh1zWIYvx7a/TnyId625IF8kVM3tKMzZKftYXSiXS++THDyWJ
bhl/P2GXe3LfEbPHZ1B8/e2JV76oViFe9xb/t34Yzi2dieqxYOVC+u1FP3rvAaaw
4QWGCWeBu+SWRwvOovFPpW+BudDJevvLPiHeQYsoSvAsJFTTA8fj4QdQ/R+i5ySg
e4JCQFxKfecqzD6ZgglsP+0Am7SmIoPjUhojn+vafZwIbXOm8M16XbvZmILdzC0n
Jm1zduNFvySjNQNWiPvTAXMa4Lrbn5rjsuAgaBCupAAAiPNkAm9N010UXHByeMYG
BloC/cb027dhM5TijfTvNVNYyvbeen52/CeaEwT/GiL+ZFVxhXMAW79tQs2hWOrZ
86359r+oOSdNwsjXMSiRtxHh9mlRElmIla/ixewFw9KflCZFpWQiPPmFjW2AbWc0
BxNaNVCsIFSVGlReKEgM5brOnf2hU2I8vP2nkYbZrXtEy0OguGvMmzAhhpXsEfK6
hEZIsBO/3goK9SUzVxFx64k0tEkUBxqXfklJRr0h8J2mWBPcAeJkKVVYGbo7Z0SO
5ffvOh1/30e8XT+k4DXsStbpqja9pCIXbnnQGXNoXPfpip9qt0ek3K8RhQf9YAZu
+WXiVwNsrAV4FyjHUd1q5Hp+mwmmULp8JuZHBU03vGUac+3Ns/XadHu6/r47ZOgo
QFideSvDc0zpbKzAOyuabwbXRL8s5EuCwW8AELT5XplCBN3seGlMsCD1uj/k1dSB
PeRf6QJ5tQakRbHUUuxglC3VHZLmL8s/TqnjIXDKXpKgOC1lsRSDu7H1MwF/TolF
C28XXUiE6ijxbotju68AUK/2bj1HurpMT2fbwR1Bs5IklAj/YMUkC3y+SHRFQz/u
+hnkYQ6rDRjMAox9T0egQvghJGeWTe4t53oGuEMHmL9IizSDTT1ZcV0JLEYH7HJX
8hKDqo17pWjl6lzJlCLQ/2udc75wHiw8HVXkIcr3j3lpCK7DJLqgy0ImgwJoXsBk
1VLVL1qRzOZhun4VDJFl2+xRA1IsqY3lou+vDZ7N7IE4D8vKAz42i/y5YJhvq3p+
psSM06L6sZ0TSI3E2f8K8EffXP5aCKyaL3sr3jgupInS+34wqFEwGAvFyhTH/7pU
Sp8m/TF06Pfa8a/vab1yL4NLxymvfqe7JQYWT1vTKGe2f1wUlLhu2qIhJJTSQEcB
c1rk/qtDg3/cddYExBIIc2/EUvO1DqnZVIh26wlfhzpC/QObcebGpfmmDCyYpHBu
QF72uzaIXa4t0kHVDtVL29ohxTj74zUuYeMyJ3N0ThZmNiWLSnyjK9tBvZiVxWRb
R6GItNoCcB76J3a8fd4pL906EnqsCyWQjxmZyUI2PGkSiYFh1nNcPxDMMMI8nPUq
TmXarjXi3d3EBvVSK3o+dQ9euAvL459lhPobvD+Xz+UNYx2qn8RIOUKvMruVMjJT
Fz9ZTD3a66YMakDzJztIKRIOzgadoaORh5cjtdHvEbVNTpQbPpGXqFfAGZjC/UY2
oljN0Ylr3uW9kX9UpAYgeOMoRIQktBqH4jE5dMb30/xc+0VD8XTjASY4utNbffrb
5DCAhECJhID4u+RuwnQPnjkWjgnqo8rO+UzoQDHKNJurJU1ZwfAejkvVuZdrxopS
LaCrNciL/35Es2l7pqbbBdJ2Oklr8dDl9T0pz70o60zlqni7OIaOYVbxr/8goJ6S
qn10n68hYDEPAXf4NMSEA6T6GPNjXM42iHcsfllYfhXZxhYL9WDPYnb9x+SIGIDf
c+yNkzgsqoXgWxnXNlM1EQ4EyHozgAKpMSo2+/x8xa2y0UaNcTZJTjcznS5zXQUY
BSlaKxGm86Ae32RUwWZpzqExyZT6KouaJYROWxzRMOGeOj5net/4vbE9ihwHHli2
L13ID7vDnOj3IPkgHDz7GZRBgxiEJwx/XnKbJBvqRgc9zfYL6wGgDkv8xNlXaYDv
nhSXiTyZha1zYFtzcEBUsYARyXZm6xAY8Pm3WWRZ/mwoDfex66XzpugbpVAtVtFN
9ozejCH/JRoO84+4n+LXjjo9bZer2qN8FIc97LQKWXi1XkPqPmn6JDfZUbBKECWK
i5GaVsQ4XJWb55kz/ZUfGzbNZVF7bhSzsoH41OT5+xUyngCPEyPhJRA/ovDQKbvn
YRI949L0vIQsFQ55DX/NF33I6Euv7/7DnfkGm+mVfWuqBcrDtLpGtMUYp56keyiv
6wNYrEuY5i8H8QM3lNjozDqnYWTOvBce5nmedAL5SrgdWZ0j4sT4OzSjfHtCaqGi
NFCJkGvocGhDCuplxLIBC+m/v46UsIhTh0ePw7A7CHj2uTFucvYdLsboQA/ig3p7
5NpCx/RR5k1Tiv85dkHRl6CFLKL7q0TMDrBwc77K0j6KCQWqOqVHsLOLyLsLXU9B
gwXd9wjKwnsDnYJaEqxi9JSgtj0xwuLPQE5/tRhUswnFzxiy66U1KUKirVyFJilX
GSk8CZRMwFl/4fT6+xNpxQeembpYglo5GLVk5Re4/QkaBFq7U2U++nRiu1WWDP/C
jQP0U4K1EBocbAaN+Ap6mWuWX219rgVgT+0XmFSy7ffZwBUwDA3UOfVdWcdensWy
nhdwzBsaLHAB7cWDfS6ULS/Qx7suargiD+F5nRquRL16o/CH0IGRkcIy6T7VoxIj
0xks8zuRBZzPlLBYEUb44eps8bKiRuhfE0Zdc6znM2Ug+lIwEOnv/+Wmt6YfX3HS
OY022UEbFwonPa61PER6Li+fEcsb7M17dw5DTohLKBme3frfcExQ0SasWc9vKsig
k81ZySocXahJjwOUVORQOeifFEDfS8oc1k41qS+ENBNoy4Hr/vppGGkU+YXv+rBz
wn5jzutAlTyRg5c5DmY+YWokkjGQUVAQGRBJzOt0i9+uZnYGqCJQ5Mf6npzRavr1
5kPVEB0XlxXh+MEW6AAZ4tAzbGbADa1Dt8ffZ5MeD49DxLHHjhWSVmUyQc8Ny4ry
SWaxN0r6fhC8EqAcg1Bw2WFS/viZ0zTc/ckGIcfrJiDP2e6D8S89bq5FYfSEfLtq
CAslChPtIYOZfgtvXC218PbNGRNZo7R1uFFKK6Dcc/fx9p74Tb9Q55owIY7cnH+v
ffhHwHeLaM2QS9rggvSJpfbo8pw9yRffTYCV070j1JlD9Jlm8QWFtHSEuoFJuBhM
ja8j7pvql6E2pxMfB216HTBAfdO2vpN2M9z/0jHzu7PBobOTmOBsHdHkfuPA2bSu
NupHxVEn3w1wLPVDcMltDEiXVEjD8fzg5JW1nQKyMY4tEVnd8prPE7/NKaMnIuCq
ZwqLzt5MuOMEU5u9L82dXgDiRlk7Sc+WVEUoNJv69eQVVDc0zMiBdLHJCuy7++ZJ
EFPe8Z5C4UaJzWU4mZsF/r0zvi8gYQIItT8D5Xp6RBwVFN1t9H/ujwl10vA63iLE
3SRmMv/DoB0Rv9Reuf3ummDmcvPYz50o0jFKAF6sKDVTxzcNayEgzpFoTE+iHtZM
AdQk9+wLWYZsI66fCEMYaB7D0PeZvwp4GaSiiVlkQv6nzynDKOO+53X51RlWszJC
PnNkL68a8c4GiAzUqSyMGqQsRQykjaOkfFVCN1eXJiZST0DJuvTSTE78z3w4cadp
+eS6AR6nYz2EpQyo9kxXXUKaMGuRhD5Oc0tf5OmtPqEbbhqdWNA17C1Yl657dsT8
6HvsTvxP0ahcKt7icbUaJsi+lQGZ3ZSm8EGbn/EEFZ8K/AFQav8iMNJGqMtd9jUR
2IUvN88UHFmrJYZSU2Q/Tp2+jqSCt99mlv7KjWvPaCKTSNrCWuOGV1PEfKKmqlZN
/56m9GngAxKVxb7HM0PjcftV3hAXew/EP9jXMcGsvGotmDOHl85cRJvXaGXY2HHn
t73ExIBd8JPpczsGLcXdZe1VMYSndXnmXXL3jj6L+4rq3XhKkJGu/8AK70K2/ES5
7Il9gyH5hbxOsQv0wZdh2bGGRGx4tWLD+7XUgyOugfFqcNlf8uB9nbJLaT4edHdm
dcdLxjEjXDoExQB6QBqPCmW8Yiw04LPCd+DBD2ySJVpBzI9CV6OAdkjy0l3+Zom6
lrVhu16Sg35vh6ckFI3DyXNBQQa1X4uDt822p8l35ssRuCr8m6rywQwohCPMODGO
iP15XGsKa2PLb17vJzMLQya/yT5TVBfi8nHHLdTTCxh/a7K+I/M0tOuwmnHZZYfM
CRWUj5rHuOBWf2C/zJeHM2m1tfpS/UXsSLJmjKe42bp2Z2x34Ulc9H/gGDbqPhpz
hmekRlO7XAvOvv2PXD4GfuqomRCmRJqJf9zZnTe/raN3P+/nH2wt5luGBXiDQfQe
sz2fH+oWZ/s+QovcNnGwoeEPXiTfBoJYgn++8YfiAxebGjdEkTn8CfMk8chTfqIs
6Vi9Hp45VBRA5jg45FrR7HE0WWdY/RM7+of4blZLOFpGMiyqVK1Qv/bA1pOGXSa2
DDgHonr3CV2CHQA8GGjBo+mVuNxN52EB3j9qq1toGlQwWVRAYkRUpafgPGwoeyF8
ti1VS/AhpZGQfwc99X4LHTbN8S8SP9iL+HRUkrOZkpZ8JaBmdjyApPRiQXlqAQB5
1FzDXQjo/RFRVBNKvFvqiwvCxgRUmB1PqfhVKiLDVkjGXLJa6TloMjol16QOCwHM
ZyjtL8Pg9Vy/y1FRjfF7LIMtSzrUHUzPH2Og3n6FBJzAa3qnp8bt9Gp9jv+L2rQA
wfSJaG3Ffgl9qUdwbeWCGzZnFawoPJasZikFWR3Im+RVtYlYDxP8cBFtI4WpyVPH
Aj93CUlJcJ8xh580CKTjS/3FVqHzNYGlX+BTYqg3rwaap4K3FI9sHl9lWH0iuyqb
zl3+RTR+RhycIGfmf4xwBjE7JGMz9O7BncRVgNNFh6fBOAmAxWd/RSRnR22D8id7
iyBuKVuBlTEjGTbmFQseRelSUeshKRpeH3t/W/BRetruHjnWtjG86OHsl8z/N5HN
nnASdEz8InQ9ZfR1LfaNeozTh6Wf0i/zXW0Apyqk7mNd2W0CopLlia3l+Ide+b3B
9r1aaBRZLKB3DkAN4nGiuRSYARAo4MilRLSrXZnztMZs3KCpw45uRbTXQI9RqRJB
ylmaLmRNSHPPo+1jR3DNIW1PsQYPWJoJ4yr0oFy1fDVo7noI4DNuoz0ZioX51cF7
Mymq5z63/yhfQdRcWkbQSgnH+en6h3fi6ZdkgIDcc33nt52hfqp5qc23GK86803V
kLvXZ0MQn0lgyy4Riztxz5lBXtP6JR7HEVbs2fKLOrS4t92FGuywJghCNKfa+4m2
iGKAjPJe7A45ZYkftl83QmDeZo+bKcFiP6usp2LvA1/GNqwhWEkJ3KtkvpJXIzep
sFN5wwLZZcGS7ZkIsIwvCVBP04GfVsAfm+17IohYa3cPIQQHg4evXcYh7IwZB+zk
1GE3IAMVhBtn3mdcutvoXUBV0vKdw45mDnHnq844Fg4tYHqmuxomOsFuoPfpnsJT
iVkS63l8PKLvDsjejp6bKBgGLjOFoXJN4g3R22XstDgZOinXDHn2UUZm8kO/oqjr
wH7XLxbB/o44vUXstMSnaQpxAn5KcIaOQWJvzfxecNywwhgheO8Io//j1jQA8dpT
GFol01F7lkiTmKAQvqeeGTUQmgYFyYIzc1nPfPrAAkuRSp7hvS8i6I0mJAqjwhkB
rQnDU0AgCzQGJPHFh8WuMEV6OzxcYjk4MunRUVUW2hcQOIsh/shwOpkZ1M2ejCow
Ykyu6HfwFd0U4/Fmjy9d9/D4X+i6Zn15IfQjd3/QLzUiQP5CjgLyWw8uup8r4w6L
Ckp4n2i1fgu+wYvgcp8gO8lBxEKfQqmmIZcm7TgBxtO1lMB1/7bZqInBL3vSmLNn
xZjvrKQW6knp3YF0pGf7eUOEW8iFXLDChEm0DFeRgWThWOapF+DqWWlf5TnX5xrh
aoZhyPPOfTlpkfFXT4V9cWuUkGV6BJo2nvHl48bjUe3v1R7Cs9vpocJ+HGALcw69
3hJ87FUAszwx6CfM3nMWAvVLB7GtorZYbCn/Msox4V7MMgohSq/aAe13oBSGIZ+X
IPtF27kLdsbY+fIZV/wR20ZJNOY7ujRAam66b/CyPFJBJ5OqJc1e2r6Cwq/zck9a
KVktjkGXWeQrfNAEUtjT81Yk/bdGXZYpt4lyko7WzAlikfva5pWT/dvkofh/bcP9
YOGXpXTJG0aop2r+FfP6sDUYlg7cm1ptRvF3ajl1sVEqZj3Grx61qLzSLPg3SVTq
5AwOJJih9tngw9wdT+xy0yHCLmwWYowBiPTu7fYE8YwSfcfrRQD2d6bm2vDyQvEj
QIJ7GYFLrgvw5bSxM0rPI6PrLxqRBQttl52OHCe20Qg3PwEV879ETDcIvaBKJRbe
ELQv6WaZKhRzbDwDc+JBCzT7FcmsmP1OCDwqjcHwPurbzeAfbRVrN9GnXq0pA4Mh
b5sJ/axnM04S0BQx/if3W61suv1afXoXjqZzK4vteJ6D4Zx28OaF1BaQGft9uCCG
Kpu2OcckeMXTzWl4WsK5bLcpOZKq7WEwVdTHFDzppEd3SqqVzbEjhiS9Tl71b0in
YjMAkCDJAjJwpV9EDEzLUZgmM/pOp61XfIedRJSaj5w40tjQJYGLTqpvCs3tagzS
y1jvZV5UfarMknAeDOyViaU1UXvJDmCdcIso8fuGFAlP6YSyNRSNjcW+8J1/JNof
9HRrvrLk74xQxjzFjqKsGSDYi4Y7j4q0mKovhOiKWjYLE9/BdUgZ1UoIFT9iNv8l
Zx6jED7O4gU4IXNWMlLahybA7i3vQaZ46h5p4D0fdxADDSiRCJTtDq1/06L3B2iL
Qc/A14Ft2dzJnnXT3VI5AX2XIuypYGxW7iSmKg8999OFE/qUcPDvuNJrrwBR5tjo
pvOVEqKtmaAITZtmvfQJFLH6WiX8cjIoqTS5fcH3QRys0S+B1p10k/q5Ffj7a92D
uoAb97qeTJl6U2NEOzCNf/TbgjK6i46VxtDSrM5Z5IQ4rikVji6moWyzi1EAS5I9
p+SEtcd2KpFJE9BdkEDrF5VRsbrnaKpf939r93yZbxbWGFsAPZu8vzNXw88pjqM1
Dl/TQbOSld+TIV6exf0HJN06p2eQ3LLmXWe/KZS5ZLGFpKvI9H/r2Kr/LXXmWgaw
seP7mpk+j5U8QlD7c50sGBR3uq0RltnjWMGR8jn2IBiTW4VCYHOVhqv85EMMIV5K
jbuDAX2f5e9i1a4Hwb7QCII+wEy+CF5Rpe3IFYdZ8kXht3P1wDaVd036ijFZA1EL
+wZ2UVTOV+09+HlMuUKaz/o5JSZR3VPihDMndVSzVXgzEYF3kkaVvZtHcS7R5Ikj
M5eaGAFfA7foHdNp/ZX0GuI0/d2y6xzwbsGdzmzxpzkWkenfitNFDNa7hCFWmVzm
qIAgqjXmAr6s7uHHitsTvYFOV4rg5WHpEs2MGmGKYLk3FxppYuvpGeb4gaVyXkK+
/XcYAZ2JJbnwk26Q/6KK0oMZxZb7Khw+5I84DLbTeg/0Q7UED9vLTBHwXrK7+buZ
38Jp8/OdO3TXxFE1/Sq9uOE67bAHsB+KJUCiOicrmmyond9uIWuUy//XSmsTs+6C
impmfxaKk7pqHCSTtnzOeNn9zCvRYB5Qgv5ULaHuVE/XvxpPzjyixxuW8U8TYA9O
w37DauJdZ/8gfq9LaawuoZPJlUKrs4PYVyeA92XjMH032ycRUnglrtpCqBmLB1s0
LMGu2+wYSHdkUTtC97jLL96dmVa5Qga6S1H3SN5vUCsltIjxUvKOfDqXEw3GVDxO
kTUq0wBRQOQrNv59WJm80HpVQc7CEu5t+4mYzJHpLzC2/bqmMQUbRFB6t1/Z1lbu
fYI2ebJFIhJiQCL7fBx8RXzO4Sj0ZwlxHcosrB1GwSI3gFUn6/bOblRqvKdBy6x3
yNIMNonK0NHrNMD6SaegNi6TjOf1pjXYju+k2I+2/Rg/j4b7bTBhB4Lovi4gP7IK
05w84MKH//m9KSZcCry7+nJ8RTUrFxmF1vgWCF0oc0fKkgL1i3vF98YJT+CH7aBR
3JLmgbQ+Z2yRwj6QEJVTckSn+oIj7iX9m173CqKQk3Gt+11LMtps3zomSc1mnY80
AL3KCVxhWIPyQIvJmluFX5NzkmTFrbgo2TfcEwAxlZ6O+Ih1pxk0gAPuIsjcG5u2
DMpS37JvaQuv6GwJul3KMwK1EuL0LBDlwWpyzDXSnAnq4kRksKbvXQySmcN29xlW
vUtLtsUdBnAk1UzhU+NOewPK5uhUk0M3Tq3b4jFqeL9Y/8a3gE8D2QsdaUIYBUNk
disjzWFJvYq/Qs11GQL3pke2VItD4if/3KDAeQD7sv9DdQgcv20RpaBAcYESBQ/B
xF2+yrd4t5a0dd0bhuZwquc5b0Q5V8xBvOSfdBF8oZ/SVQkfVh4bvVKSw95uzZf9
aKi4awTN8EKz1jJE6X0xsHBkDxy9aKmCenvF7ISpZcGxq3G/5jQ5b/VpaNkGjtN+
R5up3YiIfpLiipO6LDZu9ugDfuV6L1BAAUPRMmJDH9aVMfvCETOgCVs0orC/fMxF
ZFFxD3KEKinY9Nj7gQuKNTuNeX+1rZXcIUZCcN1C7Lv/w/OawmElrzpsvDBJWjnQ
nQ/5sywY/L8C2fSte/iNEbu0y0edCe+lI2vcN9GSx5jRQjf9vgS+tQ0/mOwHQmMt
RAB82xVrgu5ezabL31ZWoQb3Gbpe8WxZT7gxNiWKPfbPcwlqMKkuSjR4NSOhh+pN
ll3MH4qWaDeW5e57Pe7UeJ5ZSDbsvxhRm3HDSrVbzXyn8QcJjVOmhJ8FUiVNiAJg
fSfo2GcD/BUMPsAP9pZ+b4nnzigUfbRT2JN3157NfSM5dlSBBbq7Lq0DzSgN0Mgv
lvdauf6HcaHoH7n/A6GQ06D6PaDCP1QaUeOTg5OzuUBo0mIthKIv4Wkfyih0KpI4
ODQPcxWo9ZKxXXEjSTUTQ/+m0Qxevy9ZQGM1IGYAJvGrcOIUbeMqenlfUmgZWNaO
U/hcBnBPJKJZ/7cHbnNr6GRSDPLMT7FA2MJNKbL2iirt5iFAGcQAKIX6+nyJzHKt
YlhpdwnxMIbN5ZbAq0FyPcq+FuJSHYybS1zsKzExEvBWdTkD1K1mFx7Yepl63dbR
XGy0xI/Z/XLdyDz+Pxm41aZleCCZz3QLNfJFLNo0+f1Mp7pmW4VhAjb3hL+3awFR
2ly0oM/q4v8NCN+nVEBLgxigluuEvpjlovzlV+VuOqeBjCrgqN9fEdaxqhgL53T3
SsWvrqcttsb2qL7XuglV3BI5FSQzutksGO7S4lfecUapQhMoNLjOUDKULYSurVoq
01STIV42qvLCUVznLDR7sRb04VE0JiKIw+vM+TFGIkUNiFHp2oT6YLcxR5bWODG2
hc2lGQgr4RDrNPBOMvVQgMLCadPz/CWdgXpQRJU77uigg4LlzH3pOpdeHPn9ZD18
gL9uGbJMCsJEkz/JF5TJCjO7UHl3itYEDis6+j4YUGpkPafjegA1JqRpLkZ2UOEE
l3WoXr/sSQJjg1YREFp0qa94XNbbTk79b86VtYrPxpMuDy3Stxw+84eAAWO/X8j9
D9ZnnFPN1TYHS0fAnO+FXCTQs2n3oRZLxowqBK/kOTyidRcZpgxbiC3NSmOFsz19
8UoZBbAyILwgWfxJJexI0VaSEloG/VB9cy+2yn1CDAof/tRN8ijmXP5lgn1TPOno
M24zVQHOhGwLC00oGjdrjHjQLw0lrRCfm9W5uBm4UzqfxBUG/mDS4aZ0BpEQ4sL+
fNWj68ECs9WedVc8E9IZZfW6a4ALkRXkk6I97xbJVFUk26E9tmNLYqKOASmv8369
F8QeNiGwQ33xSSdpkb0Q2pbs4JHpxoF+/SfcqPuB9GyCat1MqqrW4rG2YlQyYRjq
KvKT2fYqK0GNbvfBmAkuVrMjanlxeFOgeYaJVzigxEAnj0xVDj2PBs+j58df5naK
Z69VOtkScWuXUeQTzAra70vFW63J2JD/WPzDF6YxoSwNpfTi3PcUwZYLNCcqWqS+
AJTteBejowb9elK1MJ1ImpZlvUXJxesHFRfWqiMAXBzh6XM2+GXdzAS35HPojYQk
y+t6HuFFPdECGQbz19qY6zbO2ZNT9cO9ldRRYwpocDfkeZajSZm4b6Y3wYrWKU+h
H4cBM1uFXgjutS8HbYY+sdABQI9aK2WASsenJxXF762n2ocYv3FrbaaPZYehdXZ4
Slv1APDY5DxwRMt+Hky9PHQSIChgtnEikB+A99WUOE5jbKX7iGgl+j7ty/Wq8/5+
P/Emwq60MNgvS1U+TKwgweqeVlhZbo587v+gWwQOyzR/cEtztITGtF7gS23+Ujw+
PdKg6EyFL7VAJT0+B58Yi7Qk+4q82M1FWgm9lJelYDMVRkambi6ERKAQP1b5tn2m
XQ2PT7MfZQMs/1kfLMt6pZ4Yx7ZEq83O24eTgavfGZUIRXMjkvyNJb6N+AHiitlp
RKmlYPJ5K9mSkUSA8giR68J+8lgHBLpAitOYKQf3mXV5HKLIp8/DLboHNiokGTLJ
SpcGNzFuogmQWaC4o9PgXeivtBeEVNxuCQEkKuh7ZB2vLjvu4/9ixZGewGG6kMQH
RqX73cHPM38ojNvFL0JgjmQA0NHCymtSDOe9NDlbVJPesxZCkoHc9+WG/ACZiqYn
OCvvIAI7e2YQttsmNeBG8FUrhjQLD5wCHI38h9DfggoMzPSm9PzeKEcnkdumQwP6
1h9lqY5J34waZP/VNKxl8kfSz/J0m47ivtpbzuF76/DJhMuvKPq9lQqXu9atv9Aq
+/rS0uoZar63Zy62SY0mtXJ9K6tcKxavLjn0BJFhmW+gG0uRgZfzzNSLuGVXUGHC
5oaRah4LsiMRnCXz1zIWryxNkM4lFrhLW4TqG1Tt2MybeMeHK0pUCpqIe6j0xhGk
ZEaWJ0Fkf20qEBj0ZFh2TVZKnOvqLqQToKRJ9LlZs2Dm+Ljdr+rymet5m9w/R0HK
Jz6HfSDGKWltLjSLwIrqHrAUHpW2U+p49xyikedQDuOUAs85aeRsPi7Gf40xuDbM
zS8b9TeATy1vlI/PaZpIAYZsIOZi7WWHil1vUzKAY8DfNoc2nUbsUQtUfejbt4XB
mLmsxjgV1PBsaT0099r3nQ2uH2R0sjsIAsTy9Duui353HlVDdJEAEL0qvQcpIHTu
mGJIVvDpwui/RPhYZ1eXHHK7/rZYQPhFHr8G0xQ5pyuipwpNR84QFsdxt/NcUAp4
ZTWnKKyc/xxzeFU7RHjJ1ML+RdNpcRdwN778ST75PnNvyZmRVyjmj2h4jpgqklbF
qzEpObkxrzzJc91mOO27u7XJ+Ur//nW+JotmJJLJAWqGUv77QsVv5wDdoByw/8PC
oPO8ccnkKpSIq7JNwsnY7mPzclhHNuH5IqqOVKDEMM0CL31j+mN66qedFUYGNUbL
PlPDJUB0iLCzeYX46FAmzDKOrX42F6z/ZtcSlBahWlOnf8hCj4l41uQGz1oRM4Lu
Iqs//id2wBMvPJNVrzmqP6jIHgBgPxa+f+IRRceiy/v7KGigdtlXo8HDYDCIV7oZ
1n6SY29peYuaRM0/eBuBnZnIJWk1nMdOYq8sEvcnDn8HgpYq1PDaXC/zuJM1QWy5
PLsVGGBK/D6fLRs3MFh9dKmPD+xKoY+GGJ//TjFZzo+Ulqrp02DhDJjxvucXJjkd
ylGm82ny7SJNt+YJGg4Zoc7+Mg81YRc+2PRzihy4MNj5YQvXNrMFhjXGAkZmOuWW
AZFCRxFpF3qo7U+kzl8plNz9yn12Jxs/b60bl6YblAlBkY8skDuv8rYTLATAnz7O
iYYzIsSqF9AuPRzjC2akU36zpaWUvyLYpgwv/QtwP/qMykr7IlwnxxqohH0SFAEi
kxnrpu1GWBW8LXYBv/AyTiBY4TMijl9rLM6mYyRqBzmKb2bpRneWQoXXVROgFy5A
j2TPXQM4lBV+KDQWzXQXQKZKBbzm6yYEdXwXYXz8n3nMuRc8jpI+vvED8HSzB0s7
JQAe9QY4COd9VHGDDU0zB+NC+dFZ/5TbP2cgINxxF2NYXVjHX0OTz4fhMVAOv3DT
mwq0Xw5R+N7923F7ibemXM2TkL+dcO36J963tIYwrroE6E4gx2xzkhxutiOtuui7
vKjn+0R8DG6GN5oUN95gfCOaP2Qf9IPNx6QcDJY7Y5VvytUgpHN7fzs5UFoR5jzN
xhOR7Lo+0bqA3jeAgNsOiCmB3bfDqJy16WGPJSMAuKdqilWW5Hqzwarvd4FgTaoD
lmpby1rMjiDzrzj1HN6eAdYKfQPfVwhbQvhOAqHHAvzfV9qj9IlEKDL4wEB8CGl2
A/AkCFEZ1US2ConjH04kbJOYIyE3TvO2kptxzgnkT72Ex4OHTTTyHKwB51Ae8arZ
d3SMQOHg6p0SqjDoGAbWtzaQ/Z8LFK4u8nK6A2JOOepGfQ04z3GqLoABdmbSizdi
BtldcweKcs7YE26EiDBfV8qGZgSGra8OS177qiCC1UJsKv6qAiGVxUM90rXwAcIx
m2DLl0nDnINpvTOgIiUdOfaeUm5fAX1SDUCwE9H3SU7mjkUFIJBL+WSSYNcEvMMi
eBZA/c5whw6r61E5rSjdjtKiYOwrf8twfPoG49dqPVodV//wHDXHdd4j8cW0YDrj
+GW7cbF0d4xqI4tX7DQsChqm0pWnDFNZ0f2x03sPrD92ZXT7MLGLHLvyAsYodnpX
mJ0Ruj5DQGNBWhqCoM0kfimUMr2tQL/YIVy5XVUHMGO44KwbcgXX2cSwnCPsuR9Z
OnjcrZUDmzxc+QoQ20PlgqH1VPv0z7HWo+Fmtqlpa1weK3uR+W3KDxim+P3mj4WX
AhnULsJ4hsnDau+wOxS5rYCyhsCXmcDBZbbpogKBOf15/gCQ8gE2MTrBBqar6ljh
tcnW8MCARL1ME8O43enIUsg0jUSR51VCcYY7yWpCo51/+P8Fxa0zrif4uGB2Y6Ua
r8TkdZYa8BNUX1LhDd9QtUaINFNmZNuwOq6ZSiBQHYPXJ/91CkJ5CSa5TBIp6BK2
Raas2Vwr3i3JNV5SggzYdxfap5WSEI/F5A10rvd5DBFZ/EAGG2zNiMpwiEocf1hi
GLE3lINma2fhez2Lonzi9Yb6jdcDay0vTEgtt7Z667F67LTIzlMaESYIlGHwY957
UvfPHLzkefD2N1IJC11/+EgfMwZPM6ZU0SZwtl8lFb8z6GgIVXdPdlYb3ccAnuZl
KZ7ImqX7t4u1Yh8s1YOmWRfmXjCR8MNlzUKapqtmHr+CB/K8Hic5aXQHfXcgMUBn
J9Pqrb6AGJpL9clUJVONFDYpS0X6q1JpWN0PORsQb+6X1URFFy0quh7KsXplUGCb
qNLeYv8rhxcaLD2cIs1Gu+1j2foGOwHXPT7pZv20tPZzGvGX3EN7+1IcfciysFhW
HzNM/WB0FYH47jWHrQSwvENmQvhKF7EIQ1OVvx8moniFKSIARhOSqwkIG5l2ZcEK
9nVqqrwVDrARaXja9Li/b5xwzLXrQQfFN5m6eR/bFGW+qWN/FSVCeTMhQ6ZIm0Ao
j35+gBKno3hHwV5V6S2hcvOi8epjByXf1M6ZXBkZ5/T+oZyO1YuNXgfo0YdgNB35
KyZyW/+e16v0lwt/QVFq7dVxxdns0E3XGyMDANqWT6sAYxR5JVtIRp8Ib38Y6DhO
jmyXRfD+MJF98VsNfphf83zU1e2e0yDRAfq1Ih1IeKSNpLaiBlzq3Q4nvTFcxf3b
e4sK1EOOxPkpD8GItUqpoUbSNVx4EPhxD4ItCO4+Fsc0JgXIUsFRhbzi9kEMA/Yy
IChS821oZvofof5DAbxmGiPbpv/DtSR4+10Q/x/FJPgqINwfVHSMSFqApZe9Tewh
vL1Dt+dNLmzkWZoOnKIGGgn8Ifd7OUzAgCaYVgTqUNFRlTK5QiaXSDA4p+ebyayq
WQwEQZowap8b9nH4PzC3UbbuHdfUAcCg5UitNhv1IEbWoTRh6mYl0vNtvjCynnze
vxK9qEyHvYzcxMcwjM2uViJBUTRd/vgxqpWFOceW5EtjaC7yvnTMTdPkyf2W0MuZ
kNx1v5VNtwD30jOWk0Q8YPDILir8xi4t04Yoibuzt1tvacIfXcmRc3PsWBISOC3o
eC28aODfRZp1sspT0oR9M6KxGqECusAACB80Yz8GfQPMZFRv8xcihkvWosCj3cpK
I33lgQ3yE1NIvNjN49W9eRjj/mSEh9zSeTc7WKZfOA4HWZ9f9wNEuMV7qFTshZ+O
GQqknasSYGcqhrMSExMW4vVNZyWObhy+k87yp4YA+RixfDrT9E1hlAv/HTuCdGva
tz5utWERrw/ueC7+IXESMpHcNz2Qj6CRXEJ4mL62HM/pT8CTKFX/CkOV5NeiSH9y
DLNEqEpuNpDu19fPCqHca0z1H27u7Jmsmr+qrcgbAWsIgUNiwmhdS2vejABHrjdz
yhVso2SAXD7yCcxK2o77bjcbRSbo8b5ejj6AegYuxN1fEm8XSnW2Hc77Fi+bb8Iw
Qi50GqLvRsO372LPQmDzw8eEibikvghUX5Q9sy2BcPeswGRfIvDDRd7sthjdVdIt
Qy6/FOiIO947lEJW8f25i8fCNtlrPHcTZriKIvP+Zq15+B1FzSuTdKoOpF+8eger
BZEw5r6S343/b4LkvzIQQeX9YbxZn/GkdKa5pq+eYgOWaeos64FeWmschYE78fpc
sWkrpem3vgK1Vo1pVwm59YxflYKayp73tfBNJYbVHltv9Mqb30plVj/aNzj4PB+d
jhxUWEy1X2zt7PdN/yALFeLb5xLrfi0Eym5Np7Q9DhvWgit2zGz+rrq5wdz8Wfbx
cJXVWRUzYVcD3pkID7Q2S6jMmbpoVfSEEaNbJLCqLpdL4jQ2roqyAW8QMbBsvDJC
rD0epW0u80kIs1e1HDSMMIMooFflVA7dKTHpGUyKxN/wb2RCLaLQZXjiAtXGkJCA
of8/mMfG0GVA/eJWgIMwIU8HONYngXc+qWhZyzdQZGZ76WMcj5KOMWZFs8JUntpx
xdtKlQ7EqyK/aF9Tr7xWN6thKK6bdPL39z4YbqsUPJe3ECUjKnlhKdJVc1pOTWdt
IXP8IYwvFJ54quSLUit+cAyEEVxTQvWaoio273IgRiRHxqrnYb44pwswtilupUE8
XfNRMHcLYNRjM1L4cTi0qOGKDRBmXT61nv4yHycDvOTKtw1IWZHOA0oEMTFGFD7c
Mgj31z8AlnpII72AWbOeFsKHNYU7nbaivL5uS9iMrM0DO95HliiMJpn1VwfGumMG
nOvB5XBrky8gvQVqQFY5ThtP6YnwQVZppeKFL3rngRswZxxWhXLY0FHCUOkyMOJf
NHvaq8ytL7C6kD+POhsSpww7GxRnKeDo/jvJWzM6iTm08LiFUJ0fJIPApzFOho7p
1BjW2BLKWzAp0WGlJPYQPPw4mxRLeCd7ybQu7MNblqZ/0EodclcAGL7B8JmoT3XP
8zouMKDLZ4Q35sVsHUPtUexLbHel0lS8egM26MKGH3tUwXj0zvpJ0mDg8/5WUIha
LArIy9A7txlpOH5XtA7zbv+pICV9FX6xe7yWQEsVXK45fNIglKNkfkaCRNu0UNEF
OOdL2481nTTXzzILjxHn2ArZbj7khVtjTM+bDYCvNzWNXz+jncIFBUvpYkzmNMKF
Lf9+wu45+A5Ad8BXv64cRWKU/ilvLDBGmXX7KZYt0tfe7f1bhEdfb/0IegefqnXa
MHzMUZYZ6Cwhx/XlXJ5zoWs7ZqJ8Cb8tFGwXcN2tOF276t/2IWO27/inlBgS8fbG
s8EmSx+HFUrJhtlQyYg2IN5EpZXlo9nKdtzeanaJcxsSw+AZm7cZH3obUUNySRVe
WGxu2oFONiYg3zDFFUoVEr8pz81fOn0HZGBaQhH0JA8UNUcS0KZcCU9NONSMOaCJ
FNZAK3XfIHSHFgAwiW/vciHh5mWHaopB4Ei6wEivouy6D2JdEQRAnRPjb0lpcE5n
vAXQJm3RNXTUZoTbtpgtxDgTNmq0tkbGaWBihHD9DDz1gdjlbC5gidTKm6sJUOOe
DNAOHbIp6cu3mjTlgSqkOryJpRsNvj2omIDSQeEfVYLPkkxWksM8jYRM/xzgUz2T
XUUsIIpUECqCn2BEHFrBfu5s48fC1DhDG9PBwK9ey7pKOUMhfznk2ldWxzKxVc7H
wokvfjV81NdLh32pdOfeHzZ77kKUo/cVEUSmT4MU11RmIIDwZhL4RpJfjSNt+VwF
/Jldu+R903DYYmXp3ZOJQg8fPhlyOBwT27rFgqahCJF/pQPHvqq8Ipx735s12pXR
Ka/Dvg2U+iCPVmdGu9LVN2MFFGkHUKJ66QIdzICkbkZILNNZmxRhlrKq0dprV+nb
PSyfKfB3IgIk2zrmS5PTJTF/5JRR3JLYx9h2+WYYMCsV0x3tpJJFqq32sQjt64BQ
0GDs5nDYoUNACZhPPAPcapbzMTdUfO31vZlbEsqs2aQtDqBgThQDTt9n6g6AE+tE
SbMFabAmDygX4kT9+UZ5lzvU1daAbMQjbBl/jC3IUZEoJB9k0XSyrPCeuRbcPrpH
Vr80l8wnFdMEX8thBpGjVZ3Tp8QgMVYWvvxCH+Qn06uVa48WxYBd+xz5/d0rG5+9
JN51YnGORf88cj7ytNf/AGKzkkceGNbX9GApmAO8YgfokJ3yX5EBjByjBWcBEpVl
ineH/d486ynGTRGxyNPyKEf2mng+Y2CVXh3SN9HqqL+5gGk/2RG/fW7ZpTevJfvO
i/3FD9gtllHsjye8sFqgxf+BTE3Ir0NefM4ydiSxd8lhZk89Wz1BLBvojgatM2le
pnZKbueCT4C7ajcAbOSCYBdON07khIdjnNWkmJWTON6iirlt2d5Fb5J44JY5jbnK
E2t5KtpQ9Iqp9NWIp2bMQB/XrAJAYHjDkayB/rPEAShJP29/RGL/XaX4rfgQ7e/N
bLi5ylpWRRay2XlbBVOD3MPFjLVKT4XT0XdHd8cEBEhgfrvUBDXGo0v4jrIx+dvS
GxjHm1mbzyilIcbTIci9MhxUo2fJ4OXi4vfgJYIZf4Fxj4AJO9jQ8eCTpmzzmY/Q
Jv1HrrOh+odYdK3yLBTB9bJpw8kRaLD+4LCBNEkJtc+0hHhVt+PIHVVetaGUA8k8
0Oi7GI0sjCxAp4mNH9kiHgR2tnmaambMw6o0h7cbT5tdfwrDyMFXg6XcrUeTBSjC
9EVAeYNrUItjqdww9yklRHC6/XzT5OOtbOnQM+bBmp3zPbvaJ4tkAQ4ssPP03q6r
NhBOU3D5LYQBNhvtQ215hLnEQDcucIEEWRBw+cBLdTq4e5OcaOZ5B3DgtEKqsG7x
DlNgLRc5ruy0M6gTjPwMpUQXf8pCbZ8pZaO+cf3oTPDC4SF9DV1SP/mizPBgOhm0
9Z2wM/1bfmu1x0SJ2vxR46W6C1nRvelTU4WVWxDO9AcRq/voKAhT+W2YMU+lCxUC
RW3yD00uLfluo4614IZWxd4KM4sb7usLWA6kdug7G7XWRaZoafVffXnS60cfmrlf
FHZmFTFsjmbpTm4Mr107/9gpqtmpRkW14VGiWzk5omn9yUDRqvUFaoHkEw0wnT61
/XzX8pljWBVfoPXqWfezVHpMWaYEVWxbhi7kYPm70wr9wxWlws7oL2SPaEY/bihZ
46qe+iblK9IMirUgD+gHPOiMZNj+XDNzcQiLmws8tu2WEWYPeRN6jucTG33D/L1J
vHaKdrtFNKZG8cDK6zcEqjJWbfiameY4Bm8Bbun7r1U48rhaS3l7V7lXZddQmhN4
OZHmAAjm5cBXq1DJ9U/8IKQ5n54X2atbYdxg0QcRq0VS+9jCKkgZTZ+UsW3ALBma
k39DsN+DK5UXGHNeDrdxmVEg+qxGiuA2nCqhkGm3z4YWHfJDNIjsyA+mCX4lZD8b
CzBvjM61DRDeeIsQkVwAu4l5P0rO6VjItfFmsIrcY/kapUfodmYn00x05hT1VmTV
Zeft9rO8lHJ2bWG1PLPb58Nbd4mu2tsoTmLrelyfZxl+CVx5P25rhqEHikFlWqMl
NtdpNyKixau/iTi5dpS8KOpSQLLA3KEsj35+YcA+wKbTSJ0Ec3tcXnrzFIDpYWml
Jez+f+3DnIZuctAkvzxkf+AcwbFyKLg/53tbWt8qQRll8/r2dP04ddMBeq6yOGrv
McNFP7Hv2Bwc3PEnWvS1RsMkk/skZ8sY22YNqwj47HHHh8OOK6G8OW0oyMlrSWSb
Y1CjhIr7w5c0N+PRMLXbBco23Tdsf0lwfuygHfc2w8wZW7c5zEh+nmCmHb/vMENl
rK2ZAYxeEOqR9w9enbEG7aMNJixF9Chwnp/7B9c3nzZMaq52PB7Omz/J7kqivFwf
BjM3YpRkdwGgcCEc1prwHPzlT6gD2fWugMTFFgXXZHCUxD8KfTkOM9UlPg5jZ7+e
bH1x/W/Dg2dAFKgrGpdBWiYgV4h8bQND81+AZbHMo5uV+dsjgPSu6Ecq96TO962w
ZjYJP+Ty3p8HPDBBXEcUPyyjcurCsIuZ10sO+XwzeTtPuYvPRX/cbduJwFYAGE3O
pnw25DnTpXK7eKiT7SpjEQXiEO5y4ZBKS/VnwseTu6g+osTIQsBWds2BBg8p0kQs
5goWTIF13CCx9EUShuWPtEIvqFPHWhq959KHovLx5az/7OHl0H+/+M2PkPCX9R7n
i4lHywTlnohVvv5PhHcR0rf3nFUD2og487vibjDkZw8Ymbo0LW7ox/eb2u7AQbEx
QupOwmHKvwfz9NR1lary0zSCRbfdIdZEr4lVl2+tWVU33tdmyuyEhJnvpAZ2Aqtu
5cGFzbRHL6k95i+qWs70xhzVN8Zk4sYp9LaWJDNfml1nAxMCZNJZNx72g6rs5GX+
PSJdK2Wj6dDiiIiNHTt1r3yMYtG+JRK5pNJV/bOvSk2KWQSv+vkkzOty3kvSKorL
RTQ4xAsA0cA4GqEv56V2pDi6rs5reJy96ZdmZGZ+2P1DDUPTlCX0gLJ0mSn+Liid
salyWNkqhk3c5Gac/6OUJxliI+ARLCaHA3gCl8T1PekiEWL9D0bs8uwNP5aYbwQH
dAsJd7QpOk4j1bVFogTOmpKuqd8ZlIo6ZA3hGCKI5HwwhytVdUPMSej+Jvu8COAF
Fdis5/qh35EDJWaIK45WcFJWDdyTh9HkR/P9LRLjLNRPlj4mjyi5yyqvOD05tzJc
DlIas6ghzyXODL/M6fv0/Z/zmHtviVQl5g3e/16RwgkdSyrbwztiv1qNDETSn3cy
5gPf3KImGx3n8OIuRnH7P7fWiXSdxa7lZNB+D3acparSGj7YLp8DHu2g3Ix9h9mV
BQn/D4pwVOc90sO9vyCHgwL5qalv5rDzU4Y99MCFHHWM11YvZq9xvKB92g0tZJb5
5lOn1JD4+uUI9jGDeY8agGFtvl+ROsHKf2GcbiESCo5MlM5EAHpaFG0fNbbAH8pb
S/f10I5xjR5FaonXQrsdec+HWAM5neKR/IgOankWT/3NfDmuTFcO0OjMgXPd6v4f
K+hJtJN+elILIlCylkhuq1+0h2msvUZZZ42rQ+4ZqjOP3Nm+djWp9ehk1u7VfE9J
aD+dHvjO2rDNtmbskv4CX+vDsTlbLdeZKyyrbL1zOXre+AT0E6JJRmHCEOfFDvK0
kdE3R3V+W8iprAYWgK4c6637ugsVIauPFs6OZbTKfyMWVWbRe4KRVmqUvnzsRcPg
WXNNnQyPO1imTjxrEUWmKrYpRbFYh4FTvevKYesLe204S47mm+Nzwo9zhN7oTgKi
jptMu5s7PDcJxKHc7zYPcklLRMQ4YzM7JNe3PbAAi7acyvW5jjX6zXt1AY6SJ4HA
x8AcvfBRcvmzkdnzb6F4qOsJRWTEJELZS37z6acSjZFYem4/FQnkFtI//1AP3jwl
tpDGDzeAFmis9RmyyrgczU+kaQivzWOMxp3qxabM+JfR96zxQTEQfO1RDHuLwZ7t
UIHVCcZiShSbg6wGMf6TxitYtz3ipCyO+NFrCWs244GMXBSX2170Ds+vMSxCLB+v
/lDmuOL9FbxzExWmLrIlHn02P0xhuoimmpE09Vyk1Tu/7pgVf5P+UA1lK43YijfU
8cTtTV/r0iXdN0KNomO8iF5Ok2JdUeBpWgi4xOlNQG73Ntf9bxi/LIjKMkgT9OKY
1NOqJoEw2hqJCB9oJzFZofDdFEes3mF7wzES9B8qAFqYrBMotHyj00JOgeBDEbzS
qDOOz6WETpRjpbl60i8fr8bI85kw168o5Vsg1UqODRyA/jbIGfmFZxRVTqybO1JO
n0GY2o5c5zSeRPv54H8qe+fER28Qdlzp+alPUmH9UEINKcJa6LnfA2qfEFuHe8gP
fquvjqCbtLCNMJRPD6IgUmgU3M14HqClERjEROYqHUFqZ27U8Wcz3rMLxGuMy7jN
bFCkyLxlGKQVJqQnrGTDb9ko9EwieYJdb/Bv9/71ZRbHFn32xMDFhjSc3Wn1TuoZ
PtUTj8yPXoqvpq34oyOOqBC76UEv1uLBYzPfgDWx8AqyvncDiG+klNCwF0eAwwAt
SPDOsCkzKfb6VKG1Dv2Wur7lPSVkjy75qgR6xh62Qe7iPa7NgoOWK75NTBP4L2PO
DHgJfonKywEUwF45i6+ZizsjIELT82j4ymjaIjAEttbkNtyGwNjOUouwesSHXra/
0bPu49u2/UAypbd/xARSpoZ29X1M/Tf2QZSQkCD8dVBdcNfKc4KX7hhsAnra3o67
hlzX5bH+GJnNg0fFAC+LhU5VWsBZo025RGtzURJLZ9dzPrwsaN1wJ/puG9emju/r
oaRV+Ryf6Qg8qlIhY56kIqBdrll16xgp+N/8rESw9cjpStXQ/uPU4cHc8FWP6x5X
Bw1bJQ+f7ACRfz0Wryy8tT6Y6ybvW9pCLy00EAX0K4w0z/ooyOe4TV5xwrkVocyh
0kw2ud9arz+29zmlIaNq1/ZGbPctvTdHNbUVrfyiVENdWUQw/+3Tr+baMVBMflCD
LPBpAbL+UGFVeLYFGh0xJcaQnrLYJyMrWVaRXlsukn4q0lN5sCVP6f2QsK7hNXoA
0UCvZnaNS81WBTe1QJ1ZJ3BYoEW2uEoJoRcqK+/vQpYJd4rZZ53iYcqFid654eU4
bAK8o4zJNrvLOCVPu/f+L8H0uqMGWIiOsYDwCnnQIW0pFk8Qhsf5TZQ9XqHPRdlv
7TGgU2krF7HOn6WReSDrHLNad7EnC4HK9VSpqEEuwpykS9Jk77Kq0FyTeYLlKFVC
Neql+JzIFpap37es9nDhFdQydbwiSJTb0lA6e465g+/q4SDZduGZkkGl9mL6g2+T
+dw2PaLbMISDg7OdUCMUXJG8c20MfUxZkYnv4AaFth53UvHdN6YYESzrn+GRPPlI
CLqFnTU8327Dz0qIO2C2Y8qeuv/QepW1F3TRdB0nSnC93XrIBACqhhPdQDfLI0Rc
Loku3xTN495mn+zbgHeR4dzuXQZm/VJRBlccs5go8Y6Ubz2I3uHN01zMqeSf5IoR
fV7/r/yG7bHZhfTEhN6f0DF3sX6Pb2qRICvgaVakUzACawZ68l0UQafNSICtdimF
SIPkd4/XH7OKHyWe+86cBEzgO3dEnt4yiLx1ih1pHxsRPgMp/3VFsHDrknUSGaRh
wwObOuA4uO/TmPlSkAcR47VngWLwYkm7YFQ6bnu0POdUtvE1wxNB63GV5/OTt33U
5n7A/qL2d+HaPV+5ppBVo1lDnttBzrP7P6G7c+3Q6wQfgGT1NC1jKiUldhrVPKWI
hAql/MTkrS+Cl44yeknJEvu6v6SkoNs2yRWfMYKFZSFMqFViZw4whhA8N1qHeGe8
qQFk81MPw8EIqvOi+tyR7loFeyCeNaNFilOk1QARvGo00YmwcwldKbpkE26GhmhQ
VHbaj6pWk5uJThmpu1cotqeBtNYb95/VGkFiyAcghISWe9HqeOLBQGSaSfEd9dwM
pp2maoQXYbh5skPM6Xq84hJejpym3bIlko32aSRp+PByMAAMKkMT1AXRaXImsf3O
CsFaGT6gpFzVa27aQyEU8qRtDD6dI9g28hW8s17W3zvMRrgeSXfvSmlTyrWhNPGQ
1jnLjowtFirrSxG3d4AiBC9fSS61KdbRDDmLBfLejnohBocE8AxdKRSuxcbkv3zU
K1RXbvX+5ifbIsBczC6x1F1nZz9KEpu5iw/JOLfyh8KCUjVDFDgbzMCtrZManzjO
WbF4IOd5JsB31vrDnIdRFlOU2JgNXqczOsuxYajhP3DJ+ZwEUJh9GadoP7EY9fU0
ZjHDAgelba6Y74++6BpjA6aQCNye9fdvffyeM7Pwiv1ltANOH3gEfqXNsIKNN+YS
Fa9lKFKXHE41i5dBADMZTGWRVw2JIkl8V/OuVKGzp8c3MK8MA4v0LYpwrWAuFEUd
GFHMy0xjDikGwaqoaVngiYVbR6SiYVmTJDQeB3OSIjeyKRqzlfMXKNiUAVPVOL5v
xNQLducj6ODXOOhYcToYXFF0OCoA+Mt4eqgR+chSPlaOL0LvbkXHfjJVCVkTcAR7
zAKygONwhWHSyPoH6NGrxxW2aMaAJlNtiLBx/pE48nKtgqAbFPnK/m8iBAkKHcJz
a22S8VP5y3HQEOWQkYxAxs0PRyCWpzliIfqdDZa9eHH6HRBRjn2NwuXzypipanOo
HWbroKlxt4QfbeaIs0/Op7gao+PES92uVGV9hhac+7bDzNH0Xfv4iGjAN5WECzkQ
i8T1ubBWWuoEvacZw8si1VU0oR2bWjnFo99+JjC92GNcKoH6Tc2R6Bl4XTXQBtwb
FbeEvTojAJNUHd8U9N4XgJnA/ZFBfg+Y3RPLhlwCl71UkNzFxNu84fpp5QlKoVxe
wdrM4bZKIWfgEIPx++ROsWe/6QceuXsqXkPKkhHJAMMZsPjk3MJ15vEKtWq8WAEW
AiPzIwSmMZYfqhaceLBRL3mTXayfzdDrZZNjZTbJ5F5nVe3OKISiE4hrU3Buy/nn
bpg0DagO0MH08DiaHNbyBmU33HAzbzmq4o9u9NA2AorN67as8wBQOZAGW8xId3Gn
onOyylN2FhN8Sp779inXfcCvJ7tyDN9rHBr9z4FqWVn6c5Ry88J3jZhD2E/CAj+9
qMGaJcOVJ1el4zOFx45dqSeRzILLTIzE9+E8BSpAk+9V3q1a1Qy1yYhIQ0lnaIrB
gE3felXYdZpkrJK6+9k1maoFI8ezOg/6NpRbdJp6l73mhapAWRsKaq1bAjl7Ze88
pK+5g3QPTidAaJ9vePl+NzV+GxLUb3TK7I68yZlPDwygZuXYMI9VrhsGIjtFDe/3
nJ5BBA7EuAMrX8LUi4BhROdKHUi1BcgSpZ+zXkvbwHKLKe8vDRZe5BXFmduxmnDz
2LD890EQiBZ7Lc8YWLTWyaQnMyvBSiO0r7gerN9XHkDM43b1iksV4jvEgbyzCAn5
vupD2MSmZKh6khQhneWkWEdEidrORZQgBffSNpUsDtJ2kRyHSIb2CUnkeStFJ1N8
faQFQhQ5ek9imsl/vbxv5G/priZBdRvc+dFgIDXbgJh2dRaU2leW3MFyHlg2fSJq
zE3o3U7IegHLdtCVJClKaVbMgVQsMJloAcol/8NJ7nfzvV7EX5eqIN+XvzkBL8Zz
8aE8p8XNE/f44qooyEhtQc60BclCmQxpVSHGPKvaPT94p/gT/y5akCjh0ORf0b1A
d53EfLZkpX68+z6nSqX4iuPh8zUJa9QRa5gCSiriqJW7y1sYR2uAIpvbWgrs628S
oQr7lqbBDJEHm5DpkzwryNZH73WM+pVV+mRs5UxuVMgSUfJlM5/QqMu4GReVjKcU
SKVr8ITwEOWlXX8H9nZLoa+b0zDBUHDdbStNkFHBVS8v9OmBqP0w3BKdr0i3Pwwv
/fAnhz7depbOzWlqAVhUrvYkBVXt9E15hMlBEkb9NdonFLwk3yZwCGLzWk+Sz6fk
yAqP/7i5GaKoRdvXtvWGv6fm8vPwD6d6XzqNaoWpA6KnGdNkfqR7jEuVmGMUQFFw
ubPuocp3hpOEVrv3ZQJxHQnlqCUb891rLCqg3UeSEEJzH0OL7IUmN7RLy9uWEBhq
0KZtAOkR0QYKdv0XNnH1VEgbuT6v9uKNX91AT/oCznW81xSq8UcY0bZJllEXos8U
z03DKp/oUQXwAoW8Zy6KvjuFRnRY2D/ZVJhTWZd27RaTR2zHkYL7MNNPo6sabfdh
xQflO2YlFjSAkteVIuCIxB7qJowpG6C6bjodu3Iwoj9fhGelpUJ7dk5WlRsS9R0i
HkqqtnPGx5gvEYAD+0fZQ/dtCxhAjdV6JWLKc6uyiSKEGk2iDtoIsv+6rKx/pLKl
h0rB19Pw5E/hbr8YQK8FcmmjJEDe3FomCeXtVxuXnWbnnDjK2qq0oXXKHUcxM7EH
yF7rdgMLb3XyrfQLCycorS/bm6udfXH4aRHeJCE0XOQ5PN1Jwy6f8ICgaN7cOnXF
Wey4KWtEoVgUWITvVirGNnE20XxlL4hQnEYiB2vg/jQTpuxJPhWvjxsna27rtXlb
X27ZCub4vytDa7/r52Gzyj9rFDEQozP/hFNsC0QGx5i8XPpkpBQn8a8Qragj1Ibz
mQ/LRRnobgmpekh/YZG3CzDLDcq6eWWQDz/GjC9RDTBlZqKz08UXyRqfuuO7IbRo
G+CZPxkZ/Gs3PSpyv4C6A+chr0WjLMTBtqOtQEjSst5eX/mAOp9oPmqBxmMmq8CG
vqX/1FrHc6IlSnHEEFbdZGH4oCBx8cmu940aCz6HqLi5sPwxkxGYr9DRpIzxaOgF
iM2CXayGBUQJfbF2yAeassHqPaqk2Vx5RJFyaCpRF7QMlerpTunj2+PM90IEWXr4
njKdocUTwcmZI6IMK0Jsjiri3eHzasNpu7pljZT0X4ixRh2nzQxavgC20PP7jab+
dxj171WMlJVIqrOAd6kCXpCia+U4O2A48gC2lwq7OUpvbGQBtxxXAwxzp3EenTHQ
GsFbDUcKw3aYmvrc5Jg2H6+iL7CFkPAkexutP51LwU7ZzpfVpLIeVDGmNJReVi0x
axmkhK6xTCC7Io3EetpWKMKK0JuOmJ+fGUUn6t+HttDKUbKClnnLKzkWFF7YXMS5
BOpZpDkMmiDpWlU2nsab33Ye5FpuHQRwETnC3jNyEcD37ncMGaXQHKlC2i31kRnH
ctYHuhe8aCxlKYRH5AJpAUwwCiHqhBlqPVbm3KgUKURl7gyzu+yN/QppkhkYX7Z3
kw5K8c1TThFPDnOl/+80xNvtl3oSUgIlGlTV0B2TXur4hXH9US3CZ8vVBklPtyfn
D+03piIz0ON9I9yRuLiYqZhO0rSDyMzFlkAByffDchiLsgiV0JKlXig3LYcWJPNi
hTWsQHkY99YrdfOMe3XiGIompj63Pg7xoJwSGrEGrvotmbO8IR4Ly8x88alRL9u4
dxZnc/oPd8XFbhLcuurUZyIxUJNkzU0vTfMx2fAyTGDu2ilObNcy5B1cgs8ioEaI
N/uYfzWInUL+oK4ikwZU5lWD9K+6USQvrg8mQnf3d1z/yMz6JByjBM4MlR3NAuzz
UiYLDHri040fDSinLSOZtkZC0WIBpbz9S1nlEWZHoUabsp8ziBgEdeGZfmpdhw5E
Kn2vo+zpEefypKwDcFKs4ehgU2S381Nwb3/5Cil95IK6HIfoFDHLxiEF9QeHylFC
yXpxSEU5Hc++BJ25MRVj2TLpcmfuXcZ3STlZoPmDT+HS/+o2pmsNqBNl9A0t65BX
1C37QJwCKu/DrInJgMq398Qj3f/drwmW588+uyb2klc=
`protect END_PROTECTED
