`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
04KqNYg8JmJfRVwpVtGgcWmk8riu0eMPW+hzOwdoKAdLvRXX0OOxvFZN6Qq26EeZ
FkhjOStcgfmUhErgwXSVik6k8yksI34idmX2du4HlcQ2y49ejvd8hWxuq8CodhKM
Q9vU1l8GT58IoFjJDlG0abjxswUZmSXYsvm+TRMVQ9Nuom64oth5c7edG5Soy75I
Nn0NJ5xqtuVmXaSBAnC+2hhdnHR+VbwPRRb5NywEe+90KLBnU09kPkmVgwhup0lV
1ZyuCiI8cf+x+jTVouBOg8lyovq+DGqvdWEOWwjhvJO1Gr3v3o6YgM931U7sSYTj
D6uQs6KY50L+XrwltYbFnw/H/KNEISaWiE+K5Wf4JeXmkYzbvByloY1uxOEnjGoI
xi/yTRwDtrT627SxD2cIawOzBNRm/ANm6Cq3EoPaoRfM+1aqBAyN74nYu01DITXI
h5va+if+1n7VnLgAOu8Z1/t9oFMIZUsxZIafdZMi1XDe7dHUW2zKH7I2A6cmw9eR
JXpe3Yasg4uOTOoqK0I4+6055V+Hl7wzqMdd390XoKaxKfHkX+cT12GFuXO9piwT
udr+KJYURR4tdCjwcyoBqBD8s56QwvYh9tY/kpMZI5EUDCofdbzDiEm3NjG4Sv4A
l0vtcvOZ5DzZpyjXjww8eU3EIbwIW3jVvnzzC1e72rD2vuubQhZjm1A1ZTbV+AyB
CbT0MM+wjfHB9yg+YDunew==
`protect END_PROTECTED
