`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ahJUpug2R3Z8Ir5gSNFXxadiMzqPYxMPkWK1XkTNZNS61jAPOmYu3ImN5pe+O3Ns
pV2wJJInw8OHb22FJ0MlpYbADgVn1D/n028pYRTT64tPtOuWvslY6NMEgow/TVqN
x70S2EkPsqCbIBBnsjeGh0W9536bzjLDcylxgRdxHu4qO0okMzdSwpqZit79seGH
dFgwD//LUx0fnXkC0FZETUPPHdklqeIjwVRMqwZQNl5WfpfUf6dChyS5hYsHg7x7
gA76fb/LJDZjV5sEogXLEmXTv13vUiyz3VCd7iRvsFE3HgoDeSnkrX6xk+5ZcmkV
9m8+13kJwJQa6b0/lS7PuYN9+GWYHMunA4xkcJZGN/trTWRG7TVz1lmsWAIkK6wW
EwulhhUg24XTo/8gYqBmvar2cL723HAw04cMI4AculHrnKQzGa8hSD5wdylU+d78
GjF48hfL405n0NdqVl4Hq7LfDqY6KH5LWlx2X7ypj2IkSVvHK1aT9cZPtiAr7Z9p
`protect END_PROTECTED
