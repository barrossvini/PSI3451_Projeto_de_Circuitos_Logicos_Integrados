`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XMT8353xzAR2OCNgUZlCm3uLOlClAH3QBvDdEMmx8v8Cb2fmbr8Xh0ihe4glXA69
ISnXncLEDQUvWf8kNGVlJ+Se340M/Q20KiMGHBQBFFtPp39LNdt4EKn9AWa5aO2r
eNH4yDeSlPcTSDBmkF1+PHGlFwdICR33VZfKeOXR/0V5WZ/94lrL/o9feTZvv7d7
dBehGhyXYVTe0mRbXvtogXbzTv1XMoCpa8eoWeVwFWHOiFlMNp2ZWUI2rN/4ghUR
A6s9O32oXvlqnKeD+7BzPTHH5TA7ZmmaXDAi4sN431ByuU+YmNCWT7ySpJZdhG0M
D6pwjvYWiw9n3I19T/Sca0npl9cFaPOE6UVwIMpmWlQnc0mYNbSNoH44WVci5Ahy
x4XOxyFpotaGICgONplfMqDAfhcffUpiLWTKNq7zRWQ2pVAJEjRyaxNQkZk1xVJR
OBL1vHALi5HPHmcatd7XNiLHIhsx6JIpnHT93esjMDNgX+DVvSc88eZLHWn3IqHz
cEqDYELIZh3layi/80JzYNgJ8dEmMyDZzV1X0qO0+b+otKJh7/kSMpuF+jHen4AP
m5RpMdrW0AMrkCN5qgwNGaWfpNM1loI0AtPSsCEd90ib/noKouvIfJUnmaJ0hQMy
GOK+dQds8BtMrSMWDdC5MWH+LoKgpxyWKa2QLQmGI4f9nWWOkLnUFM1QqL5/YnBm
QrAZpwxPyD8xzx8NNcp5RqboIisxi1PuhVlIkHCt+qd4v5QfsTSaEgPHWtW1q/vi
y2EwhTAu8FkqUkLqhvFKAIegDe7SZO9T2PviQ3HtF+AVOS0b6SVUurCmxKLgINEa
gz8WyRfyadJ5jvqLEj/VQukx//qjZQRp5MkfJGcTET2i8S8/cHLAPJ8HTVvumGgq
3+VnctUkp0zYMrf9d81ohsWvlzjPp3EumjzEyPgL+CU=
`protect END_PROTECTED
