`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7RCo0iSyMe/N6vzVYSl3zsmbeTH5ngmCPvxTlmwB00I2mbNVDLMv48JThTq6Mo/S
kH9zkpJpngfwbD2IF9GeBG+CJk05c/X04TAHlzb4XVzkZidWCnszwXBNJW9WAtEs
vQivxxZ8aONHYgSXAX9KFfnfo7ufP0vkpDDNiptGgQHD1szcXBZPsUUmsXvilmAl
YJGU12iTiFAH11qrAOaHQ0XM64c4dz2sHxxc7SRmVXr303nqPNFoVeXE8BeYUzAP
f4q/syN8yzpOB+gAfDUC4FYeRqAuCR4pzs/J0bD6iHZbGk7/g0qI1jdMe4cjga0m
dcm3eDlPm4uSWBJf3XK6BXwYPsq6tDB2OOma3IdxTv4GlAGdkJtuvEILeZLljD1Q
r/V5pkUZu3ysxqJZF7Pzs8CD2Pw5AiaKxGT2Zcrj6lN5Xg/H8BA3zuYLpMEBteLv
8gOfRzUErbSeMLKT7xh13WNwmcHEybkmsPEMixs1LlHW1bEpnBErTnJJrIN1kt+K
UjXiiUDM+f/qmaaJnsdEWuXsSUzGJIwJloxyXGGKRvdrE5q2LNUe2gI8KHZoH+b3
pVrTQSNugtfxVCMdkmYdDqVGXGc5JF9SMXDHVbB3ZBEVXFp5OnUMKgELi4P1XEiT
Qgznl7DwhEMW18Gyd9+7qA9a3aLlX6PnAIVDcTsqlYsboGDpN/4P7l0w9z4sRcvB
pxfImPO3+VLFLVdjf8tPwTudToQpL2OeebXkB4w3OgU5QECZ7qDD8E55vILwkL6Z
NJf4cOSr65Bd7VLwtxvekYDOS8fVgTnoDllXSqcQI/iukhqcIwAJIwRpv4aEFANv
bqqdkaPYtai7n5zxqFrUO9/02RMHiNfSFeLXuQ2ombb8vk2SBavjgzmwCEQzrB+G
FYL3Jsh2AsPFFhS5a6jQ/fDvwVC4ocwiEmtf/PPkGku3tKINwq196DCm4WMcL1Bl
Mdhvjay+IHLHO5UxNsC97LVQ1iYwGF2cLWKIrWb2iRWOhQtzf98bGiaac+ClzVHE
wH0gyemkVbPze6DKs5YwescW4i+UI7RA9kv+p6Ud4wpm+jctm98Ahu502CJBSBqv
NFyl6ONFCvL53X0T/iv2hjKlpFyhKubX12Udfb1vPvTUvaClUFFqQA9Jhe4newv5
m3zfwgTXza8sZbFDixT5U71DUA9mwgszCMVsEACDPSPXMY4K7vRZHJwekMIBiVXP
wwmhybsnSeUhHPc04wBcu029HeR+NyshAWOif9vv8zmE+P+nNLjXW54PbfbroMXt
QKWn4sd3BCRvsDMy9gkfKf73Ddmf1CWv/kG5QM3TstUigtgrC6bZF9eXn86EQ9DB
zp4hmkT0V76WxbGqn6U2cqghVrfbCfPzYY9JxNnFn09XeUMX6ylFqqaBrniqpsA5
id0vp77syNqRF/LCXl3qLtg2B2iy99I2s95J4bhFlcBArBgaBLw0Op5BWaAmQe0b
qZwWAIM3n8aH/oka5sSb7T3wZgqYPx6zdYz+jaJaCyMUhp0NAni1SgL9V29dtfAp
3XTlem8xh8ffCRbzRe9oEPDbnB5JPGxxQZWJMGUoZkVfRenXmnqzFS73rbZmIvvT
eurURsnN1HLoTU+VW2pcSUWlfWptCZ7P3palPA3ethPNjrzQeC14P/ptbH3fkQCX
MwDD9RrrAPnWYPZwirffQa0xcQO/sSZoZcp7JLJS1wGEaPEpS2N4HrqafHPkrx3e
d5BfqfsMrBOqmBL8uKYYMJYUAOuzhQoV5Qv+Jo/NFe1MgKAuMsyDrRHuS1Ssq1Md
OgztmpkZqkRErGT/VsEnbA==
`protect END_PROTECTED
