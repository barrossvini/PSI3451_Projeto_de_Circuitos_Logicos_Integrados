`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iZWdJ+igUjyAHN1lKWTqSwAbAtVILKk6D99hmGUHtskR8vAOmBE2Ah7leAPtSbK8
yf3BQNsbIJs9KhvYihJ8Rnj0cGqq/6dBP1oLc3XxnX0I3eKX6OUjUY+wB3u5sm3t
ktJAP4zMy2Vn9Y0YogiZd+rhzkMpZW818iCVxY8wHaedHljcResjWd74yLWuOg06
z9vO6wjnZWA63WEtJf5zftBj7vbgi9GdYgv+R3Qa/1ubUxVkMXf6gObzFyc69t72
q50I30lsvidtfgS9WxsAE39tHA3apBtY6cDHvgR/2xNdiiTP07dInh4+vIeoQwkK
XIP0a5ELWi8mg2w7p4p/xTLruaZN8R87GCCdTcZpEhe/jxRvB9CL96ZGVD5u4Rra
uYvEJptDdWNgyoVZ1ujG+fhqk7X3ODyx8vr6/IHtxABFDUSkDGJNtCRAXbp/+XFA
MwKycOwePmfcvKTtEa8IAl62ZmFUdBzcrlmtiFaw/bYTJLdaK/+i2/FJAIMShd8Q
82gXXwZyW+iBTHH2v1ZbMJ8TmKI/kxgQa06F46byAj4TbyYoCs5JaEJwdJV/4iJk
ZwwxzZcRnZFEWHxtAJriaFPRFvmnvIWsVeLSX4lNN2DMe78im9F85eLupq23uMvJ
X4HWkS4TZLtl0vP50Dv65Id6ZSXo0kWJ39cq9OJuETGAzEWJLC3kM6Kg/UDo5zr1
//Th77bPcrIHc2RaLpfYy+eZYGCkxP5WkfLkbwyq0mRKmsuGm6R4POty1+js6MkB
kf9Ok6Hskbd1J6VL00C5ckIJNjbLnCIm5kpj42vNFXoSXN8d4/ZLEB0WZ+O5LOV+
MVoeCoOoEFnRe8/arNsqCeP6+qpwRxbnCjYaaHw0OMhEVVmwnidh94ja3RJBjnKA
jVmOiaNcIk/1wshegrpKOV5H4EIkfPgcXBxcMb790QW4dsUSrqW46VEf9E8xRGpV
ttBbKevGNDKCUi3qrp96bni0tO+5owsB2rtvPrbBsfulHefKihNv/jWKWcKBka6Z
ijwAB/kPfcqXv2wTBoIslHvYh0zctrVv0bOUJbNkqE6mYCvxlu3m7diQvTFDd/fL
By0BUOVjrvWjKkkHx2HixsUGQ5+vL3IU7yJ3TMF37eoGPZhIhAHrBj4+Zzj5N/FR
mmCpjXgJqWISIgsUUBO3l8hhPT3t5U1kO3dGNLHtoK/7naTWRgAUtdPkka1SBDdv
SileRZdv7OPREUHtsiyUFEIOuYgLkLDrICcWWguZ1Bm99z6DTqxdYpB2xbZPPk7l
y5XEe1JLv+WcvRHFHPAtubqWuBInXATZt6UQObtR3ZkJEADuhWiJhNd6fQEDny7E
s+CBhGeiVWRH7mlkX0x77sGFxm/i8NeF8tZ8XFKCwiWLsqNevSJzHXRQAUcOSx1m
wVKgem5DAYA1Erhca2sej4KRmrFRoK6e+fwCYYgSfRy0WeMR1Bbcrm5nO/iCOC6r
LWbdNlejU98UaqUBuRwtrwZR80xRwN9PRvQXYQ1/Qv16RNpmne4I/sWuztzsYt3w
ZBc4nD/lwZi/CusKYBZWpWxtbTdn/lkfjUAJ4wBZksqapelXlpV2qTj9IgqTH+NS
Cu8zMeIMoMg9SiRfkg5nCoDH6LrDdLHrb7RCgOK1RIdgOJh0gF5qFc1cI7I8eYVU
lluz9aqXsoJdEtQNSaSKgQJF7eUpRXPCnKp7JCJ+4u+wb2W8STooWGKoAOkKBEhg
sb4sBldTFjYBqs7l5MToPXxgS2wg+ZuMSFVT8EJeSFXEQ1Hg5lVZ8kq7GwLy3dH6
dKVSytyOUcaORH6wTFjtl4nw6nldAtzF98tnI1v40utQkFIk6vymdfgCL5Tfnl23
C/rmwa7Efo9LXAn6uw6EgE40r23TdJljPkOc2/PbUvJI5Jiv3UKTrS1QBryCNNL6
0nKPGCFAMur5MiKWEK/N+/Fp/A2CSTzj2mb8demr4fVK49FF/9GNoLTCke5dIXjH
CfpQGWVViHg0ilwKKauUf9eJllxQ/t8c8DjbO2DrkPVzTMcdzsNlNIdDybJusdyG
uLFyyBjtTiyPgWV3DXL7A21gL3rboG0g/w4uFo4OKwwpmqnZL5dOAxNwGaOAzl49
un+u4rg/nYriTh086GY5YoNV3VuNcWDh/yCdVdAYq1zPfG51DKNQc73GZfwLSwBn
Y6rrtBkk8uFb4hAFvwI2EKcW+ST5xQ0Ma45Trq7KZwjulA9uv3a3SLLrJcsALliX
xiunsva+gsUsV8/IPktGlDqFzXNM8yvtzkKOUnNGI7GH+CsQNnHFMv8p3FX1y+HS
m9h44eX0jFS3aaOcMqHUOyjvWBI1CyeV4M16YojQI5lh0GbEwFrE5e+2kuT9LO3j
bBdHDPJY4TPZgsXMtSaxgkFpGSac2FhjKW6UY87ClHpuZGx8reE8GOKQTfsRUxRo
VzZCnaXG7rXPBJqjzoi/Wvu9HdriIF3koXhL2iQgpFp/hDjLG3XBPphZdJmHjqXv
gwChwR7Jszca7XDUNQpLKNq6mNK4n8Q9eTlRSGvKxlRnTtZW402hHow0vQQdq0nT
c/i8EGRVGoiuZiK/ddXOPh09sGQ2AAOHenZXkO8jny+5BNYT/6znw/LUUbjKeqOR
rHEK88ofbZN7HGYn9AOaX+YS5UaHkQG3wyVrcIoQ/Y+Bou5fTfKE3lDUUE5hJPhm
YxPp1dZcy+d0a58Kb9CXDJUbIi+P6nGnX/+GtHuKCtK37ptpz79rziJc9jGjGBXu
XUqEUZ1dKwLzqaff9ixxcAh645x3tJqOm9j02ZwvqdhxuhoPy3GixUdR1O4ytxzv
J5lra9Qa8GcDbOS/41ZZI64WD4xCvgdUwa4VjleCnyIK4R/TkWIg/QZ/Kdvo5ZQP
3ubKm34ZL/EJ1Yub/pQTrPerl01pcL+wLE2fXxpwQbi/8BnYqBuN0CxKyXDrnwj7
OM0USWNqD3T6XNA4fLv7p9sggReKkeuULtRQ4EWZZApQOUQ1HGGawHT+a29l82/I
IoNYk/aOVrHl0rN+neJQwPwwfHpkBMAhQFOvV3dtenxqWhbYPdl0+/yuqSiLldqZ
JrQ5UHrC9F/aBiVCO+IVRls+49dZATovmtzjcghc1cNWG1Bq2y1kPcKGk1J5nP5c
NG4GU/k/I/BL3Aw0EVeS94tswgSEuSaPUJEwupKmJkKhxVd5w+BhAzzVWLbnPKAH
p2SD4bQm2I2nS62AxCQM58eq8y4H4ZuEOb2cPmqYhlupqcdC31ttSnmu+OY1hC7N
NTTW3HvuOEusKdRIBInX/4sg+ZalguEOoOIra+iAt5XK0CgEDR51m2Z1wembBTUU
02KyZ2qKBbnHl9C2b5Ly6bN08cgfAj+GCFzL4KtQSANaDMpnQ+9q4T6McKPNpGTu
6RqzS16Ushoi6yQEjihm7lJrDaqsHwzLx6nGRPAKIPmmse9m4Auz+ykX4i6RuGPQ
4E1h2JycXXzel7BQjJQdcJyPEOPbz8zgXbPxat6Dr0JCMxSAH2ODs9ymGtWslL7v
EtOVfbZG8g+15rPdi9X2bnhy7zbXLO8LsjlTFRrlB9eTrrBmoUvZ+xCXBpv4lIIn
XGZ0n9T0W9yy8gmWZm9zb2THtbSALl0Jjc5vDxnlGDTJmQwbJYObM6CUaMOBt/mZ
wQX1VIJ+M9dZGQjYAAcp8BJCW+O8my/Zww9UX7ERahvHtRUiwEDKkIHTwiW8DNVC
E2DqL373aldRNDNJZNSOZX5iVCYYYA409SA3j9e/4BiD48svFrd+RxHLmhVRJE6U
e6/yajU2Bk7pP2Ba7Xs3eSiryMHzs47pJYp+ukCN44gmW04O57L5gGVyJWPGhrIF
eHViUDgVC6ixsFIpieLwd480RPAf0IW4FV1VWadvL8rhi1Iw1an5ItFpbLHumEyO
O3Bk7QBjT0KXfswrn/zVNmpHs5U6yBw6PlfpSOt9pxZWmOctbyZ8lz5HH793WjA+
PNIghaHH6VQdf4Wku59pTHx8kD8E0JBEaxmWjut9wezXOuohybtez+l8xtA64Vs/
4JEMkZr1RM8jR4A8pwuidmUd8h5VUrT1H+7S00o7O4qTFkedVC8sQ/lySAlld3IO
YE7n6jXaTwwW6hGuyQQB/uhqmQN8COe3/UNXYNJ13iIWcQU+PrrlY/RaVkj9PaFn
e6t6DnEpmsnFQkONyNDcefh+OmtfdU1Qb0dlC+D/Ea1tlSRoeTwUqtFa7wKpezOE
pc3SF9/D8cQBxojWP26P+TJnmw9hhcQgVp38WNFYbhMY+FO/262bZ7xr/9LhReQ9
PPyNONxOLZU56lZTfvyi7iZLtTxJOsAZuVIJLXB5HZ+BPfu+01vQjgfNEaUZJ7YD
gCJxZ3miGkAF3Fxempbc4VF4hy4ckGDnxdr4tbO11sTO8+lwb6aHxjBQIoqyd8m3
nqzENFzlu2TVzQijNbVkEWJ3mw/QkFmuzN/u4TGN0eDWNhPqPP2Lm4PQrDkjplVV
4is71OUkWbAS7eWDlqrM0KDbyZVpqZgPxhgdnbkj3GH7fClKYWfLPmtNr/IX13AQ
otshSCYs19GNfTjdW1qAfQ9Xpbo5Jmozxdzt7dY9tbtG6SWzevhRyBtmdh7JRduQ
CdQhNQqnAepwiWdBAoiJBPYx6fK06Ya26FtFdXUAlDMsdTKpuynDHOlR+93xrYg/
7m3c/xGi9Po3paZBzyAWj/4Og2cqcZYj6KfBOTfUWUldw7KhJYk5SccLxnjfkoc/
GaRDl8IvDNDkLfFEGXQ1fahy7+8tb5E+xKq1I/wvSMnLWwIpWxiFe9GAO8+bMe5S
qtTQRIOdRLnS/J5lUWyAM++l+QuGzYIgrd32KxJh1RVo+ysKCS8reY604WMqIhQD
JzyABCKgksPXpeaoU/WyCdnFSqVIAm+aCKUJgaOgItCmwWMv56UgOTiuiP4Sxrjh
bDSHGxDfWo6tAO1FviiUHZElQWCGt+uWtdDw9befY4Xa4TJnn1X4O7szK4IXDxJO
MSYBx8Tr7Py6XGWA/6xu+298EHdQbnFmKW7d/ZcVgUA+siUmBUTMhaMz1EqnMYiI
prLigU2mpkwfiVJx2Dn3ZDycB5qcHxhrzbLv7p3yb35xQS9K1ioabJwf2mBIUt6m
XWaNDdBduEH8HebUBiQbyUoeCrPZClzLsiXQiQGmcmlxhDuhYYYQOeyakk3BPRF+
OjkC1quHcqNrrTuhjmjxtF9fBA/pmru9KLRCw4cBQcayv+TlrC3xLZPpWYAPMFBU
rpXMl88uwMe16nk50/vwoCx4Pfzatl2BGqLwuSfQ4UP8iLeW+N55qpu5ocyZjFkC
XXp/3o7avCpv/FcCm344PhfKYPZUZ9eo+Kj8/U2J+qucMXEVHJcf2KUQyQYRo2cL
0LHWQgg1z0L6Kh5RpFTVPEDTaErUF/0HYHWswp49CiOvah+iv4v0YEjRau4JKn0y
uTN1AA0FZaKn57ibDGPNZ6ApF8RqhdxpCklpyNIIChYVzRYuhgVtjfYgzaszB0ON
VLS6t10Uf4CXo1JfL99c2RH4tHxkGb6D2mPdq9J1iLRFXZ1twIZZ/ocRjwdNpxAb
exXtu+V0fI1m+jWqMamedkgCGlxT5rIZgZv6kodPekwHGv4ayruZDA8qQbYSu5fd
Q6yItX43L0vVAdDBb3uAzcMc+7+HSoQxqkCQ7Xv9oJP22vxrTTgHmSHfk+oL5pqF
mLq+pMBrOhQVZMpDhhjbych4YsUr5m2uAGoYikOJynzTiTZ/hgyNVEgeMeOGQqQu
nwhPZHNnTE+g3QF517pWmUchIIOVcqcu+Jt9aex8zMZpjtCXphaXLqxIUFQoA51n
SJEMbkWo67+DEdffgywlkt4RatMbBmJyYNrAYaCSP9LVAxO/Ugkb62cvyDTwL79A
l3M3NFJ45Bww89jNFcQGJ+Z1O5Ns981BXm+J7t88GC6TBik70hPRiu7/K5kyGHbO
9iZMXt/FM8Eehd9Y07GN2KHplaymzr1JyJlwL02wgAlS+zKN82AU++9GvwH+i2JA
x231CNJuRShlH6SDRK+F4knvlvnyUCBgC1H5qYlDAdZSHY43zBEFNT87EvEvlkpt
h/LYlIBtcUtyULsDEtOVflyrPHA5UAiGORSAfSolnK6QVMoeIj05062i4E8DWgD4
XEF1rYRCOPYPBxS54na9jAjM3o+5fmT3KIyjSUely0IpIM3X0aMOmzmdh2r6FNTc
H24ME9wVfxAC4jeQnuzKT0HHC0ZNhvTp07WRBPbsWOpcph5dYlXLZOBeR4itrfBf
DtUL9QxPcdjhyALu8UYMCbuB4lmg8hmpqLUuMkyZGrN/OU5N61K9QmWBit3MHmtC
T/B5zkU4uVcowI0tm2yG4I01Pw5cNYV4++BUZwimRDdjdN7sBNvmWBRIzIyWdwb3
8CIarVXdU/R8eQmeHIt67ISHQdWio/QryPDtNvIKzB41o0ttbXhs/98pe46BoW7M
Yhu1xnxWygjEycqCpQCZJZ//08phg31W4C8dh1hxCYyKqntOBLsYLAo55zrMMaqS
udu3V4a+mxzGL9BiUYQX5s68XLJtJpfT62w07x1rsGPu9qFOqxxH7W7tmr54IHon
DR8EhpTEIkEhPm03XQYTqpI1rv8VwgPzhljV0EnuWThajduEQhO+esBk/ivSBHYG
ql9fojm0mWZ3Sqj26CPPael6l2joUPNAMDSBdO87TRis5Bp9djgglPMzEXLjgbhe
/Vqi7liGo0YGCtVf24ix5JUjU2f6mwXgUc7u4FzfrIum/mayuHJwT81zjcjFyFxl
EXYDvWQA0FKjw+zhGRFDtNzwtqBPtmeR0E6IYDAV8f24aUf7x1OEjhrhavu8QoEW
3hZ8bmM5IB0nMc0k13sX9TD0XeGsUKnsda0LdXPV1VQc2St5WbFk46ZNSLs7U7jL
VhwsTbT+gem+3JypkWTE+8DIeEQuPfM2qWdZFVJiNq9Ig7SwE641KFm+SO+fJ762
CQKqpM7aiggkEDyZ4To+9szVb67Wi4JtOd2+guKPSJ/CCTr4JTn9bWeAiRNiq1Qp
IyC8yLJdH6prnX9xNUdNKLZnDBWWIG9veF1eielxy9hlmS+Ga2guspTwO9RDLgUE
GNW7AIvRJvSh/gBc4mLaBHVXp0VPkXs1YdRYGO3yZCQjDTnWGkQTB2WVeqVM9ban
QMPNW9OF0u0s8sjrpLVFZ8Tod45cKx+i2bAuw1L+a4Qp7BivPNa5MCiUeWqHI+Ep
DmTTxcdglPzSOQjK9MS//Ugd7NDwNa4UdxF3P6DGU4EI6rbVQcLBbx3gi6FGhVjL
R6ffDM6D91A9qkaOxsAZHixkKZEmS8dEo49yRIWKsglHdQAhIwO3loUQbvTSG7Xe
4v516qjA5IoWpSFXeiQVSIOqXkN3FyMpuW+G4iWRa8Y1PCvDvttZ9qsb/CaurQVN
jsqs3Qip4vpGRrGlC9BakCLkkF+q9rg2HdX6jgB5VceNEM7gvzo/0/P+gZJyKXmO
RKdzHk7cXatTqedZsdD6OFk57BEFU/n7OOGQ4zuHhJQDEFUZwC88EHs7+vSMpubK
F5MMWuwXb7P5F4Xnx4y9QbuuPZ5IQ/CWwdG3ExozcUDTosqw1OdRgCK0UWRloR1s
Y48jmXsez+Qe5iAHVfeJn3yzSzFVIyJu03MwG7dbgWPLvfMPWyyKO749EeN/voJ1
fBsxqVtrnDaloDTonGcg7T7UGXd9MFeSRrck/hSWNZSvTIXO8g1djnek9fz+eOBB
ZkTXMVyFyGeLO+7wgPMjNdq/1V/4JxsZRC+8Ho2MpZBXMk9gL9QvyzNSc3vg8afw
S55dR7GE4279lNIIWGqAy6yKbhFASJZAZhHd+9N7gR4zMdiYW7sKO3Cw+kx9wQle
ChLEthrUkuQ9cpAtx8Qqnt8D1uD2AAil7G86Ni32Zw9fwu75oW2xkxQ4V/kQzDtq
xDeCD6o+uMsnWFFOkHvGeyrY5ZyDmUDMKmfJwdi3MDnqez4cnKX+Dv6CiU3gVxSG
`protect END_PROTECTED
