`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zg6HXUloyaTVo/TKxBiiRXb5EbTWwJHLggRxoBPap3ug2LuDL/dhce9dj8tB7qoo
SoA6rA/EhR7h+1wbqPk2l9trNhZX09AvBcULvunP9/kHqzVoytyAFFfi/+7x5CAW
5D2diX8I6POKBja48l4Py3zS3otM1ylGVLsWYNhsOqnpKRvdvzMyxGCEBfQLk7C4
nOPukBqm/LIgs3KpMai2vQUN2FYPISnK50KZH1x6aTEeHCUkankTE4I0G1R0YLZV
VoheqUPrErejcR84b3RyHZ4gQo71yauZIWrNAfcFCehpJXu+OCsyJZULE7EuU7PA
jQ7yT4gBRpb0ejozHi//BtlWKVgq7FjFAw4FNYv+EGar61AhV0ioWGHsW7K5qMmj
OpYy8gOpzuFIcLj5Lt7T0jNaQCOscYhEqoHZBfoLDMXdjT+gas2fqxtB5aCmP7Em
8Vyx7CbyT2Dv39nMBBQBdn9T7jvX7ip2YCqwsmqVB6c4TJdtYa1ae3uoPkKBpArm
vR+BWw6DM+iJi519/SARyRlgfYhuAqF1Qef8xO3trDcJKI4md2b5M0PhY/KNVAId
plIeXGNhJ8RGKTDBLL0IJBq1Q1KG8ygi82TEdWCN4vCudODFBzIfDTXVjXZLEHpD
ntiy4zLnOa2RgzKf6LAuqexJFbvH9fynHR4219AIEywSExgo5BWEUrCoiopWZ4Ft
MzF+58e8+OWGcTiLDR7QjydoU97eOSCvCyD+zbdkuDiqv0H6gE0xHEZn/BP30QxF
+3cppSLHQLHT7LE2C0O/fI3y+YrNtqJEEGtI3BEvppBJSiGFayi3IIBgjEBDfB05
v+Rk92Wjm0uXUHpqnaac3acNVKycI3Y48oeweuBxILFiD42piIhS8tlxL6XTJslW
kSM+7SWCv7PrqBxELdrt8R6C2I3n3Ezs/XtQ8mpnxt9NFS+zZaGNUCnzs+b6sxGX
MBYQAOgBYk0sK/DFt2APCB5etL8beIC9XUEHkAK1/55Ui3N+N3w10o51GP5Z8/99
Opf8fAGZaulvpdpatBNMyhyqX8Uq+wC24Ppg2ZaSpdQfiHY7mgE7i7YC4OqdCDLY
clchvs6rEIeXgVbQgGl9sGE2XOAs1U7ld/IL3tigHZ0woiibVpGOW//5xQZEGl+L
PYRbN70f07MW1egtRALTqEYwJ3WU5gcSJVkdHGD1lhrH2tZqX9J+cr4wywdA64rJ
+WhkaSPgVPoth1gEANJHA0cg2CA9bEpe/2D9AaLEJP8IPKLVV6NZ8uD5cx8laTNv
06iatvm0rdwHgipSMiqQze/39V9gs02vZ0k+WBWzEMr0fr00l/KrYhXdODP6/3Te
zR4Y2k3vkgJckwq1RLoWlm83iAhXvpvjfk6+iOemHd/pPQATy2YbiJYKtovDXFuM
9YtLMkuY8WTcma/dvZuazLplyJy9Y8PDjFIVh0tWK4MsHuDTFFAv90uWeGTkWlM/
SuPyjIaCAkKxEGVhr1a8EWNiZ1C7F2KUXeVbk4gueZzfNhHNA/TKYh8p1p1NNnIE
gBe1ifJ6lqfJU7/t6DhN+KQL1QbgMfDMesGNEHnoMV9tzAjf552hs5dgFHwDNO8a
pmjP1Xt51bCAM0bJ+ze6YSIwTEBmy9HGoLQHUiPI5zfXS2GeVEWOVP10EDfVEVhD
YcZGVzSOgMg0myweOzYr65ysPU5IVhdUH0W1huR/WRrrJNIHFfgz3Frcjh2dKwNv
iTGI5vMydoJicQX+JwlYBTTxfr80Pvr0hCUumTKCs7tf0Y/rpGsHPl1owgERXKCC
9FzbRH0S5YUDxJHJ8/m3cRVgq1cU4ub4oCMqD9Pk3CTzRudlk1/iN1+2Cu1QVyo8
fkOYVwDb5oZYHGajs8QCjtDgNbVSTCqnOqtvLOPrq43BEKfOsvjUaPCsr92MFDPS
jjSG9i0jcvqNUxrdDD0mkE7hvZdV1qTaccYcl6z6FUk0+WRJPhtfsCxoONv+ZJwE
1YqPwHaDPEMVpw40WZL7c/IBX2NKMzZM7mNSsHi1KwnZ1BM/qisY8EjCKzd7Y5Af
TT7gx84jNJJ5XjrYE+jnRb7uir0MumtIAkFhTz2zeGWrLdoSNw4iUYsjZe5Fp0FH
IlrmuFWXSZAFs4ODWZWSoDjPbql7STDYdiTihH7hydNmbZHuw/HUO68hNf1Vsg8e
uchH4fpUwm1qyhXexmovgjoLp3nbW0pOgOGq9Jmj3/56sQjPE+lwTQLYujCNqhWg
LXdsyoi2ntv0YgZWZStZ4F9SOwF3bfHfbvPblHt6hvNA85jJOBeYCVXk3QGckJgm
W9S1y+sIX+7WIsomfS2ak7JizeBSc7MyIBuox+LK1vg+VUyRBTc8NrBj+ucDy2YF
XZ4bR/JI6OJLOBuIgZ7Aq5i8qI6iwqM1xUyoBvOfVa9yCO9ah5BDCS0cM2WrnckO
xg395BEySRMj706m5Y9Bw41XkzZh/LN5gQzfZoNujZ1Q0gei5i2HSi+WJgQnAgRy
/8mGc4x1xzqPc/6RUPyhvruPBoc/T6uVs7f/JNN8liixiWu58NUjfvlLTy9+DH1t
f/LsNtZsfHmwmhpt5wFR1kwHEShLjWMz7uipxQ/E2Z7rRht8aBKMsoq4oiN0/RF4
eR288diSHJUy2PqXNRjZQRChv4Nf5sD8iMQLI7q6PqqKssIe7AGt2/LM6Vfic2/v
Ko4sDVdJas5uZz5Ok/LgdfaI78IvXDvFwxgo7oNHlc0jE9Np9bzpyU7bU3d9nUnt
bDdBE07C+IQGITmLg5wmU7hulodn/EMMlIUeLyZvzyGvIOKCDNJ9c7mzu1Iwfv7U
rh56PZo61ta8tWhEieQZuI01WJcvT+XmUoLBK8q1p0gQJ7NTsYg/Hhl3TbqmmTzd
6p1H46Nc6IejQUS5C/0XlGFgavQXpDcPaPKX2NrNgDgSdSGYOYo+HPN+ZDGq4Pw7
nKrGgqrnSJlIG+O6pDMsm19AhdmWP8RtMHZIfOh2Bj04MPuSa6jN4TsYM3kkZ1EA
yVnRYSGZOkb3kWBokDWJI2nIq7l9WI7h2gbTNet9ZwTzz0sDE5WovcEYstqwjphL
UsBk+u1z42Edgpyjfbms6jMhNK7BYqv7i19fpaCf5Wekq442RL/IltEzAogCg8ZV
RuQHBNJ6ZLuHUcr6z7/elWfxxIaYj1xKc7a1ZkNAURp1LvFMbIR4jKVrsd7VRv4w
os7fJsQWIWiUO1QEb9qi97dMiAAh1hX6Mud7R49g4TghmalZL6YpxY+2DivvirHn
OZI6adECmq/v+wuo95yggqrPEAMRlLNzrADDObg4h/bGMd0GBIx/jDky9dK+ezbu
hgPFXnoROn5qqXp+s+kGmWHOD5ShR39fUfiEwUxDUVwySxiWlgDtoQG3j8lVqAA4
9SyqX5CA1cgSdnUb+dK6aSk6Ga9dfQeKY5rdgH7/C+hSBpnJSTFxcxPCU1vF5aOH
9tXb5CwRXE8lAyr78GguoDvdYLvcdzXzd+yhWxKVdX9LhT3n9Q8mKxx7jcLFfsvm
cU1BKDO5+zdDJbzlGMbXHVRln3Q30y77Wjom5M4Pcx1wuG1fUOaEJuxBax2QJkxF
08Dw8BTwpLkHBx9iNscQ5LpuHBpWi6CAdGRr7NvUOtcOyXAo9zkmad+dp5RIlcmH
fTuqqorHr+xOlZ9ysz6I964iHl/HPjfJwE46b/VfNLOT3z15yAK6tv2E9CcuqMN/
QHb9RhlOv6uuPs81G9WRCkbjt0U6KF8XaK3OE3KRymPCJLHxVmUPrvQBdLiKrWyt
W7QXHbS6q6JYGazGEzI6+S/xCKxf7Ckye8i2AW7stoH49+9s2MQ+hyKlDpskQDcV
vpKJYI7an7q4lBXqmXkYfiyqfxnUghWjQHelw71yqr8NqxkCpRMxjp+lD4FIUNR4
NLYRSdUVwEaa66CI3qdg6pGu02aotO4S2xzkuLEuD8WiyTYaGQH2T5uKP/MMBaCh
ifqjGWAW4BdWCzy520y7vQ1NVs52cdAc26vdF4qRvOPhptxSTzGN8MJGiIO/c2jt
khSK5Daf3GHNY4H42Dbkir1q27QSfS+WlYYRDXVK/mwThy6RqDN4d4+kxa9XBBB6
ZuoBenECXIFWUC/2bzCCbfTHZOMe5mqIqgJ46E0cxHYKnv5/SS8UdqVpIXFLKqhf
jbjqx1yfnynJWuzRWhe8bzdmkxZ4anxhRXnKj2V8vy7Gyuh7TOCSiQ3QN7bXPhgv
F0O/F+AZWiIhrQFZOiAYQ1Ld6dyr9QqogHGwZZWe/AZP7uFwfo4zmUfYt7tErgs7
P5uiic0Fx8UFzN/XvwsDlVU3MPsAxtYLkfaTjvrpiqeV5RxlBw5dO8Hna1MwElBR
nK5kgfGfBWV5+A/UpiUB3s2KQK5uLcxsBAtTRlblWvSfhe3mAAN6Yq+x0GpX1x//
l3MaqdSZy4422+na6SRMraEZSItXFaoR/cPgtlXABANPndxkDagxKz9Y9zRaonuk
D2pzmb82ZXtaCA3eMB8HwDr6tb2hRnGIAZNJdpGcDBnGHhIqbHAIIA+6gDcm3Qf3
ZcvDZ5uV2VvSeVL6QqlEXnj7EdBYz5v7iwaNkggppq0n6lRR5sPYO4K6BxM6sHIP
`protect END_PROTECTED
