`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jmS7SmKU+peRfvaR0KpSmmqNP89o6PA4F5P6BM8mw9FfBAWQlMw/p2BW7NXAZNTV
J8uu0TMAmp9WPdWLJ5Bi+rf3AXWnuIMqLWOCdTMDb8p+NRsglFlBIy56rKkFntu+
cob+oouLGDPYYqlWFmkQUEEbn5PQhBxhcR0jiWR2rmN7EkWbPZRC89eRQPBHseRL
K8GZPyzSp/wbXQ0OnY/ZYfH6AZh3Ff7Ej3TXD+6/mYwB/Orwy+M0xQxETx3i13r+
eB7FkJLw55T3e7v444iE5gb7T3kdSk4/dwZQt3hgx39AnKYgAD0Mhe4Q4HP5DlFn
Ir9BMPsQm8aynj39pejvCP0ToThqCZ5gHYfu+jYrzp++jxGgcoCeDZzaYEe//iqN
xS4JvaIUCeYfCS5J+RfphCAYdp6+NqetRUHUjqkgjkXn2L/OgWuDlkPkxe3nngL3
k1F6R0ZLzdCuTFkdrx+qGmDaLVpLz9+KKtlar8niODmHDkij3vnr2QzIGegcTJYx
XH53Mf+MTxyWlujLLJgXFGJPGYWlPa0MFw5qecolMROksFJljvg5Lxzhlzp8SrMt
NyXpfbO6SR31lfyHn96xeEJfbolfQjj/9QMWDzOo3KlaL+v7eALwT+GqumZsGrEr
7/tpV/lid7Kbvf5qt3lCkIDYs30ciKyS6p/7V2p052ZRzY+2fK0P5OM1MXSbPrw1
/gw/TPFGJAAPbYfFhOqSqL6GVK5wgpco8MYOGbBlk5OVFJuhkig1b4VEo6VbUCVD
c7tTOdLObGfhCpSfltKh0AKebwlmdJW5GvzUMDfgYN3G2gguRiYSbmgInAnxZcLV
RPghvgs082Rrc5owQNPuzX2zpfuElGTtZoY74AYff9dbuYVcRBu3XkXms+nr1DMt
rzLx+g+oW+/vML+u7IUs6amX+iVSU5GIc9OI3Jp978/CPxmNKkpsDTTrwFeZnjU5
yu+JaU5mX3Mig1k5VOLU08aS1Qdt0HCzs0n/pNQciS3LuNX3PnVGyruseJ1ZQ+mt
jLv04Vz4ZqWnAgiXzFZwM67Ez8/N4HUR2XZrodGUCf/cgXCJ1s9/eH5iGsfL5yJs
JRrstI4S3fkBVWW1lCaE7YS4cuvzJ2KHT8nb4cY0vdhusWu741KO3wFqcIv+lmVv
eKDjiiwEv81sZ5fH6egezWhdAIfz2KIakxyG1YaMrz2i8Pz+jEdQrtQhpcrPM3zN
Tcihhp0lHwSyXB5UJ8u60dxfSMVAlpMEW2+Wh6EFPxSlUI7E9tZS2rAN+NVDRrti
bHyKBDkUzGgwhdgdAffuFvZFPTNekZ2liPx8Mved86ocX8dmUL9d48yocKERHndS
0eEROBkTQ7ll3apu/LKelhme/CpCWQCY8NU0rW6ghBd0stcvPXh0zxmak0+xKwiC
OsSZRhbjE5RJwkC368CZPG4xJ3eLJbvdRQA4xRjdcv6CK/HxgirFdGlaR3yjxwTr
yoi3Tw612Cs6ay3n0gb0OHyztF8S6+6DXDpPr/YQLkOIJeddU/imou/3XdHy7HRG
x1KIC4GtpyVLINkqL7dP+HloI7aQLQjZdx2wtEf0czA85YpgN/P2T47JiCm9qpnP
4xlYeCMe33UJnOAYYRXCFpYpU3RyQHr/65CPT/mOkmlU5i6aaEWpT+OCeCYthijE
ERUzubQ2nX4erU+99aVatRBU8ZbhNSNu7yjFY5aCB22VuHUImVfEwD5rKKHo0ydd
5EhqYe1JSuUNbSQk3SX/tYVWEoLWNns1BhXdKbGuUmHTYb8zSVyO3YEWM+qwBZu8
AtpPDg9UpZzbbR1eQR0lAj7S+r42HmazWu4ON7U++ZlTjI9bLd6AouPCrHQifuN3
oeskSsBLPoyuPlcCHPa0N+L94zkiKR5Y2HsNamFAyMIrCwxnfAjwhUbm90n5lpL7
vToJpJOJLXHdmy5bkoMPSKtOLa+KXrk9v30I+UqTOhQLwb8Uwo8N4hzBgrU8XGTd
keGOscm+j6ZgnHCridlb86a27Co+7uhAVzil8AS3telyGApht58xoVd7pwMTZ8QC
o+Y9GWAH3sJUcIr5hA+EGkUi5YtarWIVrTVVy91ngqeCuxbZESj2ldNgayxJ/NjK
CGmhPEIkIsnchLPGKsLYVZrDxcEit4vAjI4c8OncsNKOUMBS725iKM/aBmItzH6W
nHbyBhb/xp4T9JjAe4YNjHTGCKUvHDEX6LqenUPAyss=
`protect END_PROTECTED
