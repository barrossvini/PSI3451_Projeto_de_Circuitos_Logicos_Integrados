`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4UFMZ3udUcZlrh3+gHDCef5vIZSHgwcd9fCoH3paOZt/CeMyn6flwFDS1uBE62Xw
fMw5WO0ZP8zlWIbWLICIz5L/6yy30Kfd3EQkQW0AyCq/XD6oXRILnqH3nAZhF2pC
P1joidVwyrfMR1Y1Dma+W+L8Jh+UDUbK6nMf5+7YcAa7p4aWVXHmCtqAdjCTDiRf
KlkGrReMJaV3iFjbuJ2er5WUolT7WwwOi4og4WHSiOVf140iyex8oPmyZYCCjPE/
iXMdR/irdzkww0hd3NJZY1OvQ5i+qf5c68VUKpdajp2BE1yVHsYMrWg6HISVt+qP
lqgRbn1neI3r2XLPKKJeWWUjOgUbriONpxsS47AsB78eGh96Acl6L5Z4TVyDtXK2
d3kmbsjUg7LraEoK2RUZ6Nlcfk+cK2oxG2h1Gc5WCh8MZn7om1dS2MSeNcyS7j8A
YSeq+LQwaJqHKpTYJUJr0I0OhoxpFmT9MA8sOog+NgubbZ+EIXYKgcysZJyz2877
UGENdsuapyQRGzIejjSChrQmQ8X2Kd+Cwmz/MUJY+RJSgUa9dwkMbpWxwNS/lvca
AbkmkHzjfnL457KdnkFJ9qk0I0TtutkotnATEVP08K1S5DfN3iQteJn1D+JVzXsL
ZUYp9XdtnCFOkoI8jHlXBFxwEC3ArGc7FobvzCnfjMAUQkh/Z9k0y+RF+LMAlU9c
+sqLUSriRXB9J5qe6j8Otdco+jS4YrzNaIJ0zWyL0yDutW1M3IPYQCcpYu/TG9w8
0H8EV4rfEnU5hc0RZhdff+305x0Jstde7uL0gpPkeHjeAFB9MIwQAvkGjL4beR1R
S9voPmxdY4BAbM6ZwaYxJhlN9GYiKtyxloRxDxwengwMgzitafh7w4Y+b0qZm4CE
/rGYkrJ/cnG2gDXOI5W7lPu2YaCPVtuF6jeeY0jhhR161rsNWitdEugwXQnaKXJQ
52uOutcbeb67oG5Xt4Qgv4zJ6WlmsHD6yUaBzKzV/jyPAryic2bxwMtP0c+Yc+7Z
E8RyB8YAUbaPApkLsz4AEqOtuK+FkKNSgNnJyF6/lzK5teYbDrP7cDNL+F09sICN
hNPcmpSBEnbym2fyOA9ZdRebkVjz1zEcBtOer1zFJrsS1E4MjFXctJfF+df0MuXL
hrUNMuce6q+f80Uu74ixBjTYSn0fvy2Sv9NFOgjMmP5oNS+G6DLCw2yHc16Rcr9L
MaKiEd4zz2tsFdFKSFfB6XrRA3hliymwfWOqMUCBltN+kLJVkp8rF6Tc6FycmL7g
Mj1oYpVQ07mPicBEB+bseNguQ4e3aRd+Lfk1Evu6mLlZWb2yyjUw4lqnOxdvSi5F
5KFNGtp6lcIFi1Zb1A5lhIW7CmvRvanuy8Z7BQJ/N9VcaWd1yUxlK4B+UnIdDzWF
tSR5+RsSdcoMlditU2FvatnrTXAnjKMW3cwctw33rqCEVpwNTpDy9EXPCTrIYigD
Dh2qGU6lPG9vfFf4Qkfpi3eTH8f4Whvs9u070/qcAHCZyFh/WfzM2WiSXI+KOf+/
TBk7XSMrId37669csH9aV8zx/wtJH5qxU5poFrAojvAri3l7wl/B38SfmsVp2NOp
9POv4onaMx403ztgpu9FaC/mElqOe3pTYR0Q9A5Fel87b5lxgjb30S8fYQC9qmWT
megtHO0p/0gxEw0VYgRrqW8CPJBttGNqjh23i4ij3rmMpgsM2pfySFbtOeENYrhS
MnOHZ9rcedI9/5nIjejv9ox0kZjUwdbFUKpIG5VV8ZjkHHXzPo2SDSuALXmjJd6Q
R8lcz/KsEgU/zahVHO8s7OaautyNBaiq4UGKmASgIxx40caT1dylZlLExFriWy72
87dRvImijyf9epd5ZOGGCs4KJyW7uXJOd6Q9XftobR4CJlWmHjBiOhXN3lgeolil
obJR/Tj9HK8iMq/v+HY4+47j0+MuUwNvkAOSW2yZ29wZABDQnV5Ke1PCKzXRMhH1
ZzKVd9r5LiaGCL9/c3x0GRMkFyr0lDdLRjQKzHy4N91WTeYESZuzBZLCzgc9pEXx
2Az/ztHuIQwJHfUxKH8xs3IPsrB8+Mg6R8fDOB/T9HWj7xir0yYi18soMHwEYmgR
AjZoQgv17wTWzwqN3nhGFKUSXOHs0/BJNai9BVyVcFxnZk6LtYttoDmL0m/VGSfu
/2D+HVN4pO/H3/A3ipjn7KP8P3HWMUbw7xOa0W9vQxQVFlnwatpXEvJ2JSM2FkQC
pyV+h5CDn9Z/R6BX+o9OqFMe5VeIB4bZG0DdyksW3olpCiqdqyM/H5xTqQ275cfo
SRfZqOiDGl1KJv2K72Mn+L/UyFT5bnIDBuSan1lmNtlqviPBnsMXDTzzEc3Uq2cF
hZ14heGsCpwKcY+OEiu48Lq9FGoHxVbBTWlZ3BeX6uo8blmH3gPavKhxipmDbByT
PcJDXjthWbfpsu+4/IQjRoPRyD3Sz93MuW/oXkSZBPnZsYwNQtGneH4kw9c186Ig
HTgm+DLqSm6WDQi/QXmjOe2A0sXeJSQlB70o1GkZLA0=
`protect END_PROTECTED
