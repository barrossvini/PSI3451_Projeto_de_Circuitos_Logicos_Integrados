`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IQUOi5Jl7E+JRJjKPyxBp14SKaYIePJLPqdaueM1AgXZ4VAbX4uWj4faABKpSHaz
c8JVrdaWrUjl7D/rkMRVGkkCacJiPbD+gsXTWO9td9Z+xHy8U0Snns5jCQoy7jza
O3DFuYQgeRFyJFZ+iHpwFNJnaTKb4813Lm+8AfZxPFssmHpOnYbhpBRlfKnEsonk
S+G0PqLt4vdwJUlLoPeEHmMaqEZAq0AHG+KEjnRgXSu2OSn3yoo7PQ1BBAkq8CFt
Cx8YkCC4179y+Or2e0Z6XSVCxZ7fa2x1mw/2KI4QFQTr6RzS1wLV/dgchQGPDzNk
hSJe02QcRlw/tbrAOfizmV8Y3nLJQRaEVoFi7qQsSMwoDkUwIT4ZNWwRx8F/Wnww
IPaVIxY+4BHgKdLRnQkOD91wGCvZOpGpunciL2o9dP4iLlAOYCEjTSekq/hzNa79
NaXybhiN49tYgJ7wL5DqLR7Vix/nOmU6eux4vhtT12Pshcy5NQHOp4raz1TqsYj+
DHQzsg2Wi6BuT+AA7/WKUIguqf1c1ViLO22HEeVea9jpfs8rzZvbfTJDrjqsPIOh
6/p6VwV9wJLPCzXLS1vwuhNiiObiT3DOlZ9zOcpypYuChSTYT48HYD5hJaXF8P6B
i2yexSJhNF2cnfJEZmtTRc/Z+nagNzB9RKu9LheKepgRX9FYRu3ajAGqYcKtbxUB
bhv9OrcVxrT7kyr2qS7AjRtmGvAM4hyKiK8zrPKa6tQphizFmHP4Qso3VTkq/UiC
93BSlaWRWEkX55sFvNRsHqTKPg4q6+vt6Y1l5ZYnUFmBrizUbm877LpLYGu5fnBE
K5WefPbI3MzPxLRK3B6w5eDit/q6c/WpN8FB93twqJW8jMZCqagaqdd7n7mRvhQu
tnv0jwBzYyQTVCXUt8p3SMkJVMsfzNrBEUeKf/iAtdUtZbwYiZKdAkYyKuUlz9EK
SYVKxRsZ6+v7HzflBrIVyMluamci2uxG552aOd9S6evz+PU7gsZgOjYzF4NEFWKx
VlcykrSKlP6eak7ikJcbhXya6kfghXFb/LOnMSNyC3cyQs66E/fxBXJudA8fGurp
FsSbpLIqTZUda0JeLURbMkOQs8mF4Bq3WwtbryVoAjPs6R5w/bF7qAGKrwXTXzJP
PnRa3f0KvpTbAolZT0ygmpMdDPvfgWZ73lKvsiWXThEfULy/4KaPREoiZSgzLjzX
ByRHgYR4VioEzlet1w+DbmDipCoXpxq0/yq0OL3w/iY84ZSvtD4wCP/I+vXCvS9I
m+OGXfgubI5jiOF1XpsEe2i/6yQHeaKA3KNSdx9ktluuAZItJQ/nx+aXVQPmRPt4
YaeOYLsHCts5TPo7tjeVnMgKbdbOn389jy0PgO5ltHid+/PQszjJPdCAbcekx5zs
iNljnCzGXRV3gG4+1ALBMeRO8pPUrWHmsWG9dHFc2cLXVSImyLy0WN1qej46/KDX
U/0CjU2uoF8gFe/OJJi/xN+G8VHcP0Wj/16Ms2QStw+NW/CKVC8et9Oq9tDDf3Gr
M6Wf3aRc+AvrvtQDWtsuH9w+T7XGnU0gWch+ScIzqXFXlk+RKo4URVxkRi0Ona+Z
Xxv3tZC5CoPUh/vW/mhjCh0WsQx3GaRNt78ihC3wZVPHR8uZDl/6L42ImG85V97I
47MXBVQxEcLcmeAq8P9LPbNSI91EYsghv53kq8ycSZQwC71yuH6ZASUm7qe0FOnO
aEqOpumdzjE0dBl/cSmKwTgwYrhFmX6EuErwWmjUrOi08LapKP29bwWEg2Xn+96K
7h+Bfi0NCAWgVF3ej24B5QH6R+PId/+QITASwBHM3xKJglEn9B2/Peaa0UW4K6CF
6ETaZQ/6dISsD/V8AwLQxbUmy/DCTCKT3vGPFwBGwL3p+VN5TfaDrtRCvqyBa2xa
fYUPzBOnabUnOwgONFZt79Ck0Cs2d3h8mZZOy7CeR+pxL2g/OBFLMqIyI4LvRX2P
GrXLzOWW/3VgAS4rX3PYlkNCWmda+ePSHcpF2PMn8pBOSy+H4F6/gnheflZmE46R
lEJm5j2YHjYtODUdSD6A+E6fHeNjS81dV4IX5PucrLbj/lYX97VD51AICZLfE4lX
4Xw9Xrx2RVeTj6f4OQSFafDI/x2rZt6dWvEcL1ZYrEB/tXrdoqNhh0Zp4yBfk5FY
Mb93lUF+NteI+MIDHHfbPvEcYqQ/lSm6gYP6QY4OpK1cDiSUcvV5o5mJZ/hCPevm
5Yg5sUOs4c1S07tbC/6Z4gzJCLnHbz4/11ty5od69PxS7xSmn19F3uIfTU3tRGnR
7NJO8+JciAgdY0YZjJTZ3HufdxIXB6pT9Y1CvCuXWpMjCMbnBvam4PywFVvBYVaB
FNu/ji4p5PSNfbCu3i4srQ==
`protect END_PROTECTED
