`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eGFJ/LH7PkTblEY+hhpSzJceJ3sfzyDoKseEZ0gNElb/j6No5Fa5Cn3KLPDtqxj8
TwViNIQwEPNd/GvE4oq0d5kQnqhx5MMlj0mRO7KLdCpEBYw4R9baXrtIssrR1SLN
UY7mgfpK+cQkFzxvSoWFcrgh39IPPmNtRlNIdgQ2CrIrqNvKPl8t4Cqjfk2UbCQI
t7p+Dy0l2uKjVZBM0zdM91cjMsyXLil5LTttvWCpbxeZdpURvqVgXZp1hl8LDZF0
hFgO3/TiA8szkJVw87nIpDzZGB7zOv6uMq/nxVUjzgky/qHVr+WJJOjBjc3K1gZ9
DUlxsTaIgdzqpB6ufF1NTm/Csz9sKctRznXLl08XbiwCJ5btDoWhkau/XZJ4FEwR
+usoF1NL4mp0LQ/2kVzFBaqTrUe9Uo4yeM1/bvKiykcAhIELfl5vpnutMLX2U04h
cRTqzHSjF2nFO9yJyeCg5QMfYnYXc95WiNw6ejcgTGhGcWptnshphF/aEk33y6Df
U+BVEzwr24GC5jFZIsKXVd2hXJFqAjRp1DTGJWlnhBjGjtMYN5UeamcspNr58Uq6
pbUdvKbf/l1y7ctgu2rI1nxBg7M5r76NtVyDye3RuXdfpFY34p9Q/wAR+31UICj8
VILEVhSwgr8SFLjMhzPtCYmx7UE4VWQqMARZukENTlqnsHV1TC4LhGa7jtLQ4vyH
NMinWn5LyA3D3RnB2OE53i5hjGkFsD0eRrF1n2BS3+2dL2VfMw+iDolO+s5Krceb
qAQdlvikolC5f/u7fCsqghLwd0ZOUpP92tqJTRB4IDXnE3QAW5Z0wqvMiaWdQhhi
sz9kzG6RpmOJFaqOF86CgEqsTFTrRGEIYdZ5xULPU/OBmkjKWhIvwHn20p/s/h2L
lf3oQhzpiKLbPImSyoTITojmC2PH8vCTM+u1eiQu33kfxhphdO4f92Phe53LlvQx
IeH4zZwhvhf0XSQwF83a93vbfIWKNQIlQMxGq19+ALfnKH7HAOj513RGAORXqlux
njPPwtkpX4DJmr1+sK+Go8/aJWZbDbAXWICIJWcY+ChAKE/UN255u91+RqTf0jSH
b0/6qAZ/RRONIqjo6/w+luWnYWK1GNOuwABA3JBU1G4SVyx2cBQHGNliFjJ/To6O
wbWuoO/QYdNYmmNU3D+P92uNAdEvmkep34mKtP6vhTpdSd5LFeGEGIWaAwRA327G
YGN0Ne2m+soPKKShmajooX0OvUsK978rfczj/TQbq7LGN2tBkFmRgJvzWiuuUUUu
Ik8JcyZBzMVDyXN3FxiiDzp+vM/4ACTewwuM6u1LB1hTgMgEuIzvnh4H9pii1F2V
5Oxh7ndfChZdfrjN1d3dCI/kryCt/6fWxZTBOF/2NZSAd4TbJy/Vvv5i+fLgKbSC
lqL1Uip9Yvlumf+0C0sGWUat0EN9+DswMMnOQzJsi2IwZNkZREWB/Cwtxzgf8hjX
26RhlhVKUfz/tfRh3N4t37X90qrQvj1UXczy9iLHQYGuIK09SxcuBArZViKiLY8+
cHyq4O3jMZ6D5fICKaczqdA51gpn0Yj8t3Qxj6wVAvSYfLgheVLayy+ug6xLS6cG
fDTnqUMjoZQKugK6QqgUZmlle4iPFpGUsloVpT2siu5Sgzh2wH1ZqGnBGMKNOoxl
y5bQgt36Ef77ChJDPIgCUiP5xr2y2+b8Nmhg0bGU1oAK94StaLwu3o/mptLw6va/
wdMxKaVwHyqHCl7xvS+w43S6V7DkJ5avuiCgF+ZLqMREkB1XGB23QAqwSV7Ape77
hFx0FD4U4995uXr+vpEigfL0rPsvPRMGYYzc7oQK+FAwj0UHdSUWoH2rRd5TTcwB
T31FWPdlPi4+KSGe6RyzimbSieHiZ03FWwfY7buSL4MyDVUEmIX+pul5C/BxG6q5
631f/NK9ALSLsmGsxWIcNnV0DaijZODrHFmPPbgN0+2eaez6kYPsME4cmJcXdHlF
GC7s0WUBx9MS3ZUcpcErZvDdItIw8MWh7rcWc8YNQI+iMklXKmYBxfPZm8434rXY
iiKLxAqeNv1y2Lti+NzjcFxB7njiBr75S75EJsnCgy3InRwxQu7K6S8c09XCGfmZ
0NoPeYW8FYXe4OQfQQIhOP8pnMOIGPEDjk2EXa5p+LFAz0bQW1l7jIQz+emD2nAF
q3wSTo1HVh163BtxLspjE2SjjcjSmRgMzzwxE54udVcUr/Oo9avkhahu5T4hQUHe
BOUl/oz/TXZ9CoFyvgfc458LkbQsntnCA2JsnT7nBXVuPj5IS3q2oZaV7pikqSgR
RaWHJeQZKbLiH2hHfHW8vwKhImygwgtAHOgLkbNR2tOsk7lw4uWTMug8Jue+eSwx
mUKDTPLbjwt0CU04BC+hJH9qdKtxwPA0NVk2HOfaWx/qE5IQW4PTHEoa23dtSvco
Id4kyltm4hkeqb+3Q1MEnoNm/zydHHVPOATlmXC6Ww0WqtO1tFkJidIQXQgq8ifY
lplNzVsiQfJALUfzebsN96D31jYfymNVhwKkxXy7J+PLOpFdtL38dzttws/tJEOl
ratG+Dd95F4HzI2tfshuXUhwA6xHDLTBOX624KQH2ow66LKqhGaRg0FgDb9eUA4p
/e34Fn1F/3Q2H4bvfiaGn5SxOVwp94XONvRtANxgxgc/fmbGiNFhZ4OZwZsZRd9W
0x0WzfnPoUJzNyc2OnGUqH4s3Fak31hxE1yEKZ3Q/Y8bbMriiqUAsjflElzx/HK5
Dv5MfAkulR+toXVubDeFImgUacgVD6b5cAHt6NYpRZWj9bQGnRa/g93wPFsHhsH8
S2vHKGfVJF+7eFkDO9y6PQdwDEJasL44jxahCl4skIBj8DYjPb3gQXbW8ZGlnnEx
BuDshcJ9G1t9LlgevGwuYxVYCD68bWcANs5xICi4vsx7Wod82pyDQH4d86qLF71Z
WJV7nR4Y8sSTX5O+w6u9frXMWAcVRUUDRO8bUtjMWjSMUp/LchBGbG+yAY5LhPc2
pGRCDqIqje4jQmhosJ1pD2hsPT3sOIkRXyEid3FiNiIZLJANr3rKVgNXlQbxXwMS
DOdx+D7B6I+7+Va7hVGy27VBaQMWGBqATdMyvxtujz2GGNlBCY08S+Ae/pKentMY
cgPWxRFeoDj1wzk/p35Lykvux1ge5HyZbrFZ3GnFLmsrXyECNWzXz3WUAAjNnXX8
EoLea08QYY0MzRTougsTi4itG06JJ1CZONEd1+Cg7zsOwdVDntzXwu7z4htfvfgg
JTPtrDybiUIVIZDj9P6AjF4PWNREK0yYRJslykAm1BT4NSfbsSyIAQMLK/tFILJ+
2Xpq5qaCZwYagXHI0VIUZdeafCwVjeTsd2T4hKt0JdQxofUMQGXj1Q/kHROio75y
MNZ5R24lge8ZVzZyj6R7b54Bwhuk696nJZbtBbM4AH43oDbfGZDmKT8H2ZEsLKxL
jNw28liBumyjVfvOnCSG7nuJxalJxAPbhU3IQhUT3q4gCt7bK2NgSbYpvgVCRD7C
qXGOlpuaDSkddUNBi6xuNdrcPRvzseHRNFmi1bFrRxLQs6vYHk5cZilM857esCPh
0pACCkkKZueoBzFVduJEvqMW++vXMh41j/c46SXQ4jcxvovNGcNrbLXxhZJEPh/J
z+V4LRdzhwgEO2cas7YtqTRwc2vgxLbeQvlREcq44lHWREox4wjYoioDY819BHPO
6307dhQMoW1J1spkDE/lu9B42WRja59E9ftItJJrYMDohgdnfFTMIOkeHgw/OrvK
OG0F1OulvDneyapG4G8pYnjQkMbvZ2ejKAJ5KZ6ZGkEQDwbOPe0y/LR9s8CaxRKL
aOxdH2bEidPlQhpIxkEBGQxURC82njby+qUiJe+/u0MWAHs8Fj38tvccTVQX3uMA
kUDxVPgfr5hj1Ag7kHGp1seSXWUikeKh1QPSje/yQ5Vhy+XwSFSM+xGHNJYLzjLp
xEHkWwZOjFNSe6gpm5xyKBO0c4O5K9HkOlruE+55hCoUiskqxzuyyycAIZEsR+AV
9QmsEzIPK7cDPBIEsEz0GgrEuu+pd11/a1/4YZkqfSTDyBOuEc0CIy80ruPqPKLx
nCAqhNX7j/5tIG8BPzyYC1CvqbDWEFZt/5Z3vGqPJdiekEl7PoTxDzCpXw96izE7
Ci62iA6v4EAMdPG7tqnQfiblxtEJ9No32BQMo7rgbLVuN8hvW7gGCRszmFDGstgg
4vSaOtoXDL5qFtXDlb8ccQMYAshH+6B5a404XqH9OG2l1+LKtWRhzS0SFKRjv2Up
VvEANqU8f6rd7fisDuPW53+sFbpsQYIWrqwsAN7dGX+yQa1BB5NvMTX8DkYsoh8H
qzyutaRzvKHNthJxi2SHYJb3TbHlZhR5pRRbOg2Quc5ZOcm1kzvwFVTX1OLCYex0
K4o+sVjo8+GomaMURGWVx+oqtQ58Xw6VaYZuTQNevwv2ZHeBp1hQLXmN2jA+j04y
Gm10ZcxO5drvZklHgJCm55DrPRR4zlTZq9ITwt3nHxjYGUZGfd7BlHhfYd3fFLqd
8trGyuvuqs2yq/l5ioZMABw4nvg3yeeYlL7hZeoFrVTQVf3OFGrWSPv+cwHyJT8x
pFIrpcEJenYwj8tT+sh7WCwizZrQiB4yyuhNcfc2JbOGYQfiguQ51Z7y94JfTZGQ
rIJurPfI4G76LZseZnORHC6a0mQlFFY28dlwauY5GRWP5cIVd1AI26RcfpTcgQIX
51BBijw/5OAcKeFD+h8lw2j/QZ2t6HBFjZmt+UQgIKpWPu6Jsh3jn1d4IU/RB2lu
eavCqmaClQGs+CpPSLNuGp10OFCQtXZvMpw71Ff/thi3drRYzVkL4WZgutbzN8HJ
SmIgQDmgC9Wc5QGSGa7FpMtbopUWUrMmq8FoFI38u5t6NFyPtRVqarxh3a6GaKv1
I0DQMAI2NMSyR/Xu9ihsV2cpupB1cQgsLbPPEmtNA2CPG7aq+O8HfVOu568KfzBR
u3pkFFokbCygdURSyG/f9z+fccAcERtFpcL2qB/u70G8NNEZQh6p/k3KPdt1oJf/
LV1enmDKhONqB0TesFTV7E10Kc3u2yrzvwUH3ehAd/bAjsM6eadecXPG23DJnajh
kNkWYz0L0p803AdwJmGGc2HTb+VZ1dSzL14xWS89U3PjgVyeIUsjn+qfZZv8mKwU
WOrwA31sdwf94sd7QsOxPztq+vKkuEH+zex61MHtMRAVvNRorRpnZT8B6IB8wTIA
aLfNbleVU0u5mLAzyA37nlKkiQ4GMnlrahbkdcBBFPUHquV/r3PksxtYUGS7vRNz
dmr/dcu/9U7c8fG6vVwcMm0ennC/hu8rospLb/KQACb0VUO4L5nA6W7UyNxVNrlg
Lc6gbDzKCw3XH3Ek7yjbFSjcrDQieFP5nD2ZYDRQR+/FZuKP9Kxe3bPafavu/1DE
LD+0Kowl9Pcg/FPgkDJyTUo7kZyRGPfP1p/dWxa3meBXh+3YigCHDQA596hS13co
sltht8HlH3zHhhbfXCmrze14jhMdXS+BYlcv7XhDFIGdYZUPJX5De0j/ugySyIFR
yfSMN2pisZbaT+azSNEPDUGmArs5/u7upy2N5opZRUGgpBFpiEPJukbYO8e/8PyN
Pn2j+4ohsOjziEFVTxnkvcFGYh4SnJGU6bhutwu1O2hPd2mJCncwP5tuWDmJBjU5
zsuTJjEDIcAc7Qy20G241QAxCVBIOBso0Pp+ifgYRldQ8bquJC5afSb24YRKdnwT
fpreHn8WyO3FZJzOt8VmlnOMBVmdykeho6fQMZpxadObnZJg0NomCYLqryqa9ixy
PZhU1MFmCfu/A/2PlHVLHBNeRqAdA4che64YrvMXZHLOAq+4Gj7ihuI9kItRJl+8
DecpeoH8JMhD5WyHe3KEaYyMK17DtC6KGkQljYV1D4oLihhauKip8ZvNCbsYpVTX
fvmtQotuWb4dJ8HSIiLaTRwW0g8DPh4nmvZcwcboJmaXDoFFr9m+ypS0LnkvA68D
knv7xa+wYDVyE9573TbHkYDA8oF9OXpFOxzmg2pOZ0rhcV6KgXn7Y/suDjr3pKKP
kYkTLU0oOtBcO3kzxmFk3T/pNwoGuckdO7xEa8lxh+Hdr1FjRa6nERbWE3AzbChz
GSRsDCpDAr305Hh1VyrpgFKubahUDXP1UYyXgBnYp52x7qZpUoKDh0YV7gVMAD0R
G1Kso3TehTh7CEGDtdDikESrzkw1EP0R58imGIbe2bPgSUs9V8yJIaH10z7zx4ka
yO5wVSz8o5OLx8RD4ZJQDdP8WXrWf815tdT8BztoGFwOVAVc1cMdmkGRCyMxkyA1
pzuRULLngwk50FXkQOX8HppnihOC6orj47j7jYUbj768Aad3EGS1y2+Vci/3BJyw
SID0w3DFF9+B0pK8vyrIneCs9bHl1gAzRtdCO+Ony8x/rNPEBLVds/0ZPx6StcyP
uaoLXf83WJjyyH9Vk+yLx/LpnLWkeXBA5JZ8TCOJeKcH6eN6SdwZbIJCZvAdM3ff
a4S76c1mQ8yrrCdzZ6rE8IrimrZNthIkl+z9RSoK5JX/j56Uy7DqJBd/HXsoBXs2
NlzKqwEzETQdTQM6uWAexpF2U/wWJBW9yI1jEXGwfbsvpi1jRSWNJiXKi85qKm5U
T9TSlYsxpyjMopMHXCCBdAuAHbS1zF8XKhJtJ8/1GdnlZcid3y3uUaQ6gM5v1MV1
touwlyDtnPAt0+E99WesAEEnaIJ5EGfZQe73rjxWK1g4jV/M3KmIqDoCrUkSxJkM
31xHOV4dhR+G/hJux7MS704st8yl8FOalYu8pZBTngaW9xEGshpGvYS2xCcFUuVJ
rff0hLfD4GiMTCSaiOytMLUX2woLww3w/sG8kVdO7/9c2XNcbOghlKPrIh8dDn25
lEn28A4PVjuaOSqKelOB/G5DX1GVV+0lXff/+nr2dcNVtrL34R8Jw9VvgM41+g6l
wQI1pIkhxfhlutsiLAGvKLFpTLnmfUHIUUgFSHxlYCmRxnr+8rIcYMBwl2z6c4TY
4Aj8n/DMXS0k+SrkDOOxO8HkjhHpk+Y6bcJ5xgj9sx6UB6KM+zuCdL1FywGZv7UU
nQdpb72drF2msnAjKMMePLrPdiWRs/q1xdbfVPUTqa3F+dbbrEp1brPjxCybL/03
g/5HrAi7Xl/LXr5XEBWP53CZfNZajNDGpQKfG21Ir0LAnO4cSmD/fEGj4KfkWfon
hdNM5qh5CMSXCHO9GV7qg9f/7aQ1S6mRDV53YYWTNUkYyMFYyHKvQMYaogQhrG71
9FnrVF4YQrc2IUzet8/rRzKcGrXblc9WK1IYBXkW5HZj7qRxjYOFeZ630VNdV+k5
pD4vcbFCT5/DA4k9J7pw8SAXFm0XceMuZ9+iMhoMvRPbKWhxFfK4rekYS/30pqgO
XvNkoGnmAlUrkghH0ygkRyTq/78VcxpqNsw8rNY9nmQZR2ncbQPrzYlD5pGi5/x+
1GXT8BpmDcQAgv2U297XGTJj3qpO/UCOlslHzUm3RJKOl4vTDvBQ02FWYl7u1VIl
eNMclvut9OtpnyG6mF7meVY2agO5ncGuhtH/QpveX+205/bxuCsIkUE9CeUNtbeV
xNwawtDJfEygQ7NerQYo1FInx0SRNVQ0CwWAAbl0A168h23NMvfWsN21egX6mTll
xcTilhgyx1xMo0vsM+DCKviWrjPTA3+pYOAUD3LfwtLa1bYfTniVR6N2aXrevYFF
BfQiag+htiY8Q/xdV/WjJjDq4yV9Zmdh/+qqYwouaXfZAXe0MxWfzu447KuFgbD4
ImbSWibU/6yG+ctn/HZMc1EG3WIZPY8zTpaoZs15AYmTkWXrzZq9v6mLkta6Q37M
hK8yFS/WMWhBQCvTnMF2Vf0MAOn3OtLEv8yBndrTUiR+RLiunKZT2Tmd0vBABpxe
8Y7k7yMI9FZzbKlTdnVHUGqEqjMmJyVPg41bBHxoMoM1u9nKv4M74MiC6zHsJtfB
BBpWknNro/oauJ3wVcHMjYYbrHM3Xz0C9K3rW3OaLUnDwAKUOL18u8aIV/wOBX5i
6vRbLiB2cjZgcmygns0onxEYfQRIXyb3K2JA4PTP8eO5SJaVtTKMwYpvJBYgz48w
1ByAjtFsOgaqBH0SE79CI3h/Pc2WzmPl/2ORbr8HbgmjmYoRDN2bRUOhJxdAGVuS
5bjfaRVxTA3nVqJ1WdjMuzAb5A6VKR/JXkDKehyfpJXylG8vCse5dZN+POZykVi7
ZdO9BZMllmZmW0Xld4YKCnUaHHa8vUMyHNyqw4IgVM986AQVrnnhECB5foiEn2pP
uyH0isGeu37E3KIfv5p3dpXrrID8+gH9qntLOxluopO76oSYLETMPyG/HPY1p/GN
4PKmHXuJME1pRQMKp0s2c4BR4Hb8/0NBSHuNduL1O/fRWn0i+Ku+sMKfycaPwCTF
N6Jnu4aMK08gDIc2LwrBI2j9wHG0ZrPWY9EIqFnI+Gpy8IxLzDKlDC2oyKmbW7Jd
uZ7Sj+EmE4wydwalbsWv3mUculO8qwEMGgdpgcp0ssK/sTyIlA/Z/l7q6/1gj2bj
fjI3YtPGYMuOl2B6GfB+BiIlzYXi5P8jwgohukrzhcAlIC/bsF1Ix9FpQ5kdTRAs
q5ywt1wG57NMP0zjmSoaeFCIPy+hwdzcSXs43wppwez+YzRnejxqzByIfGjgTTM/
zSGUXfZ/2i79mBIJKuuD/U+rzmc9Vf/HkRQB2kVmFm7fSE5jIYtPEtJA1kBHJexi
ues+NaVZpKMyOGFXmLHJXMgIi1hS7579R7oZtDB7887dekhAU2ATmkqN9LdtFnLU
q9ABrSc31FyT/1/FsM1K9VILN/UJrYO2OSZGulGAAB4ZGdtQeb7ZWQqf/kjG2plB
mOekrS8JwIHpnvTeuooYFMkkuUcN2dRB1jZrPlVSTLROIV0fr5DcvM3NtZAOdCoC
yR4lOM/fiKmwleB0EMvFQtXGdy4hvF4KBVMIDm+pWwHTsVDzx5+7442V82Ct8kDj
UmOsPva7eylOYmCK26b0gjoYJg8dotBryx0znsMtGSkHcjPEFgWOV1/HrHqQI6qs
POMOSq8mICVIWu5W0D2+4FdRsGrN/uQHvS0QdCiw+3n9erJBgYyT+AlOUAwR5l81
3WtGlP8dbhNxwNu6C6GIugRRHLnLR/ASUbUuA+tqPdUr2mGZfQVspH8OVBl/8VdP
YscvWNtsbGMn/bbVEvutaYQ9SCT84TLVNAddsgHmQnboTna/wRlr1rePMp5qGxyi
GZA/W6jfM/xfKku2Qm0ent5wykx7YI3MN9Xq1Zb3vChqSUYYtbrs1adi1ovu5hZC
KG3Jb/1Ir/zONIa3iDwGRTX5vXxcDE/9DBcXgg0a57e+y3HYKYIG6M1trhx3kqJr
BvLOY0s3JipyCX7rnr6i+CjebozzzpIv2VYRa7eayCzBv4zxbEGpytYYTZv741tK
0JXyA6837GyvlP2BBrpZO8BP+QDvBVb1oTNupIdx9fMJoagx/zR3pOqqfAsrPiGQ
xUO10NvqQWzQNwgINVbg58/8nBzD8A3ROEB70cW6VZT8q35tLJ00uxmUleLr9Jmr
M+MzXELXgxLSSvVnfPY8K1otG/8EJ5n4kQZ2mxRK4rL5I+/EwUngRgVeSFw2aAVC
IlbUANFNur9L8ANHdJ2ekXAWdvlsE2gVKwbCAO41IhFTLDEVH6CIEGZ7TFttYbNm
JkAAsuTaFeT/OjvAVJVI0CasLdZLRDgpz1idjIIeoiYNsZcPkXRx/zL+R6wtGI/A
F7ib5inmNI4RoUTSUsnxtkJffhKbQOEevV2ErdMBmmKRAWBaRpGmZ2MTr2RoMIpd
wPetXV3NKkwyj4ETkWyN2V8M7CZQ0gSSq+YU9oUOS/mGvP5KoL8HRsMVi89ZpJ6U
1yRx1lec8j8KGzxQ9lJ03KLhv1axHZ5cCQPW1iYhfks+yU3nQrC2d7n00QiEEYYI
zni1CtaLyi5iyZebYQvGq+ivvBvp31ZZFAa4D6FSlsfkHNas3UFQ7YNOXKYSIPEY
uFxeYwbhvKjBwAzABI7TUPMRc1l4psfwNDP5MlrA8KvlYClJzjWxelSDdhF5izi8
4oZKqZ5IaLKKC0ckGBZRp7Pd5SfjY2GoQIBZyGaI68zL1wRH5DXMOsoqASbwT8Fr
3zPFM2Fc+QkXDBQwjkMEia8dcvXPA3QjgpVT33AWpPpY40V1poC0wPQQ+YMPP3MB
HJqejlktDmyK5R9AVzijr8BoQctuMComikFmaT9Ul9yUCRXsmGO+66Sj/TjmQbEh
jsfhmI7QpAQDqRG2OwZWq2XEf1+Z3C8Ka4F0RFXhV+bT60yy7vVZDQMxTuH4rYOv
bGrkb2rY1HvCKfwKWWvGUcAZpwhuLNGnck/ZNCCEphHCjR9uvxccBLKCvAtL+HYq
2S/9KdVh5/4c5s83Y3s+pOH7SSvcL4eJu0rueDTBP8nlg13ZU2CKBB6Eb6aeDg0s
PcvOb/XuEBCMShuljXA/NA==
`protect END_PROTECTED
