`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gsyF0OaubQoJPGWqxOAnOf/wxD+cedWr9TXLZJvW8uEQ7fgQa8BZkiUIJRrVBLee
cE5Qd0ahOHUsLHBX+wXCdrw2FnJj3UJn7gvQz1ri0hVwM2D3BCB5bBh94gGWPUpT
Me7JRyVEX0i+WKEUo3cPWklDZobG3nB0LO1QUFFcv5nmz/6/QmW4POqCiKwgqY+u
CKb63qliHF6c4bHbyqeNQMcSfWxZHgqTjV63AV6plGbnmvKY2oSYRXlVUaVc33AW
oig/0x4fPBoyxs48GQHKvJ0XNbY7GbqODgM69Te/TrJHvgd9rNsD9olv5sjfcca1
G3JpCx6iqTSlLFC+NTybjHd3wZZkcHTrxm1C7Yy3P1cF6s1V4Fnr1mT2MvfAA1B6
yP/jZ+6j7kyX1aeUIVYF3u2kjGkfVx01+zqh7+CQAeoAL0Th6h88yLv33ngFWNQ4
PZwdR/ke/PcBg2iw1Jr3VA==
`protect END_PROTECTED
