`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H3RPqESTxpco+fQYr4SOuIf0Rrio7dsdKb8uGVpvtQ3k5FDs2GfmJsBRH5jy3GRd
mGgl8dKje6x5adg9/lV+w4o+Ge1qhVsNO3VbIBLZvTXv6rGNVMh0RQnOaaEshzhG
Xsr9nD4j9wgIkk45piM6G++FlOSyZTv5/RGJqKvExphglc2sPNOeShVNK1lO2br9
lads2vaCPVwqG+u12H5km15LU5kwUhyW6+NMbTjy6cCd6w9cVpk6CKFSpYVnMQE4
IYTZemSTQjAQvS4H4vj2QOzIG1QkNsvH6QxYKBYDWPlQzdcNhRrx/M4F/k0KKIqK
dei4ldiabPrv512nsyT4/78bx68GoHViSQpGkShEP8zjxoXjgPEQJQ0ISVuvhwvj
ovspuHG5OmDXuAILbn8O1cZjO4G0H3EGsPAxNDd4uPq6tjBYi++WO7mOzmib1Rw4
q714hKaFDM94IH6eA9E5QrSO5PBziALxyX4i2QKiJvFPnnSTlq4mP8l3kqzmUgjO
gBP5ig1DkzeqTz395786y5trjVKvip/frKTN1VAUDEGMm37wYHfWItgxaGMs/kGY
ZuSxcNhX1g9f8yUQBVbMOjYkOVivRndk9rhYXQqrd8GpYDMEna/5kjl9hy238kcR
x1XFtp+jvWnJrHQiNWhaMJo0wQ5nZiBCTREe7qcbPnhsZi/FeqtAyWXmJByyOfHT
+/AxNPuZwjJJL8yJj9zlPaFHN8F+CCKnOha4h+csQLG23r958FhEwVMiyG9YaKob
LbNqYpjGcPvyRLNlQRUtjAc1s3OgQUiSZMmb3XGMtjM5ltYgTE4WZ92u7Uba8BlM
zyZqZVRqYeH50g/A6s0vDENsq5HlODm9Bidf3B8s+txQXP1sNPcC+LZFtpvicljm
AYa3b+/nXiCPyut8HSbjVh7CDSrbLQ79bDBjfKTUMZ/uCthi5M9Vc//pBA1Yuql1
6yeWSaLQ3rxKdnWx5YLEbhwQ57pSNu9WUIjlJRPDHj06fYzI1TLedfEF4FpecVkv
Fy2rbaajb9OUF1y2Yr+ULxFlDQ074c8CcTlE/W9xED/c7T7D7z3WNYZBRDLe4Yro
UKaXsrDxwlysjhLXM2OevTSHPfS/o8F965+v0b9IWLbqavI4xTbjp2M3lBoj5Ns4
vk7SKMgVG2Mol68mWiaTUc6UC4nbsFjuFriLjbVvnNMXXVQyEsCBBMcoedq+4iMC
DvJLlheHYiOpgEki1xWdSItotVIv+tlv83b+JdCh8wecfP87teuw1EsRUgXwMA+H
wjDsyzvK42La6PPIaqS1AxesNPvC/4E9RRG4CwylTLX/CDNfva1GxSHIqkJ1Ht83
r6N+5nieIsmfgY0GutxkAJUb7zCe7+uFg2iamZ0nPQQYjZHi2g+Qte+045WQBxfO
naIpUy8OWZPe0UzopJiSXE6ICNW8kLiwHkkPYHMyv1+8kJe50MrWKazcTdZrA1Vk
lPQ+ySPDR+IjQEmvZrw/mXakx0L0EudZJQVFyhTFNM/F+FZAz+3keb66K8wZKD+F
CwIdVMNdjA8sTQo9yby7h8IZh1VwfB2FYlJOZ3SIIzSYd6DWM2bXmojFSpFRGBNC
lm2Z04wIsnuoz5j7IDZuXDKj7k1+QFlr4GJcaSzRoUg=
`protect END_PROTECTED
