`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WmDU4l2K5y2crSbBpI4jGFdhK22KeTwuC9gIzvGGHTvTSiNM5divqGdRJcLWDKUa
3iAyzq6NTARDKJCW+oTfTNlgxNGAIH3yExUdmy/myqQaryRhTWt7edLlUKwLqVay
ZkEle+4oCvIsJzqHMPMZX8XAr76RLbxzjyD/7f0BzOOSXPmXewA+cOA3IBQRPQpn
5u2V4i2GHZGswgK2FmS3EQSS6674WSs/i0EFKacn+ArQsM7v4wndXm5J8lYZvS/9
ir6u2ZUbd+mbMPjQYBDkjBvpHoCW6bTx+a0tDIFvwRqPriIHlKyZR1q3E2C52bwf
o67D0sumNM+xz24wSkJ0PN3nj2mrb2sifiPjqwoqvK3kcRVvWqPWd0DudPLe8GUj
maE0/phtlX3sohnILKN9aC3deCW8Puh0J6HY8J1FKDuQMxaMguSWl9buPFhTBz/g
tdnWkeHJgI76RmVw3Z/NgiYdFDA9yQi8e1IaPS96PGttB7XfkopamFVXIIq/2HcW
wmk0OSkflVeLYFtNqlEkHE2fY+6rC86aJPlDAWLrQEt1nxXVdwwAgIoYTRbuZlfl
69R4jPWTQ2L9VsIS1Qw0BKBPcpKpMSYXvpWUkaW86ZBznfUj2hoOHVf+m6i7QTya
PvvxDiOlxioBHrm2fI9EnGvKu6uH/yEspBD17CnYtKQm91RB7k5a2ZYxKrN0+HC6
V72BEKze7/CeIjs33FLI2wehKdaDsl5nfBw1J+JcmvS7/L0orvX7lDjiwq4qPbdO
244hfmf5SapIxUt1kDfme2T+8+eQ4259uiPBdDXb/VdTU/rP82Pj3q0F6pSO7Wmg
+YMfUwftdlAeQrLLO7kGfAsXWR7anXHoq8DML4RUhvo=
`protect END_PROTECTED
