`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y+o3CKx78RocKOpX+vtIqqm29zOO2s40jfsivcuPhz0RcVWWa43W5ZMjaRYnTgSG
ipczTfbLhWFIi02IxmH9OFX1c68T2uSb/UQRAxDSBZVHS3+/l10ASl+oCs6fwC2J
XDkML2DZ7co1i6CsDW9CCXlFVNVPuyoJgDcBKBlB+8P0CvGn5fx/TULkgG+sRKBm
wPWo9CbBK3HhRSXQuDa4XeD8OQYGUwrLwG6cdlEXaZsD7CAp0qmiUb/EQ9uwNv7/
/7v7jj2b3BROhAHX6dfvwS9mEONn6cMhyiCQ4napJcdSkpWfXq3/DuytP9MVIgaV
TUXl1IPYrRrhYmMTyYKkOsop6vezgdmN1ywB+PoqyBrD3l32Mx4xtEdc+7G1qSRP
9wO83dttNTV/U0en6GwOy6CqNlD3W+onKnj3LQS/C81aQM4jBGIVP09d5nAL9u9P
XdUJLS5Nl9tXkcSEsIcD7EabVsQBAJtsA5w6598ceuRKofoXxjsPD1FbxBi7ie49
o4/rT20uVjNgpR08Mmx/iYLeyynPrwsvhgDUiiN/mnrLVaXhQF/7GPF1Fdx0SDDn
+W2597BLQE/6h+0wu1WC706N3xX1jmt1Y8rFxG2BlZH82RbNVtS4a9d2HZ9NZwsG
AkjwPrRuCkyW8jtXM1eZBMwsqj4lPRSVYnXE29z5KX0pfga8G9M/J3ynha/aU/nX
ddm7DNheD+k/f2MiAUHYJMg56newVZJ2edWXknNShQF8NJBsVcB3xJn4R6jiWwbC
p8ecW7yP7N7vPt2GQ2RWilSQsIOuG/apUAJ8Ee2CyKtlrVjDU9KANBPm3rKtdCEb
S68cKZzTndQFvN2XeOkF1lMlwa5y0x00GYKqwGrojjFG0+9Fm3s2pYWW6bl6nNyP
GomaBkcebgodezgup3UzGQjpS11AFBdsTWL9SX5hZlmYbx6XCUebW+TDBiL1qs7I
3QMF6m+9hECtLaJH8+lER1KBa4fKxd65FC+siDNw0AFTZzAplkWUsPk2nadyWISa
/bP38LL8J/7MWa5t8WDm+f4c4zoUc2rAkYyQp1h9LFkHsywYUAopx6JX39rW7ero
ZJN8oDca4S4Rvvh+fntWWv1Dnj0wqDOr+45X0neco1xDVqgNp4etYtD1ZL+5/FYv
ebPHAycne120SFjfnVSC8vubMkEkmfK3N7jza0kz5UX8rzPHHWdZPiatC7HdkqHT
uY1yh9Yl0z1ylX8KOKyq+Q==
`protect END_PROTECTED
