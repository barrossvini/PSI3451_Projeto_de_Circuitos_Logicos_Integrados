`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7PODQPb4IS295hZakXgFVp3/77tM6U+ODhtoKB0FykSxI1Sfl4n7sJB959yju74l
JvQhdmGufPbFai+9u53ntaNan6XO73TCRn71XYgb1SuNaBj03xqjc2Kk7opP61w8
ihk1N/vSAPpBK8+AAt+LeY8GjNZcead35y/kkc5Lm5Ztp3zJraA2cWV98ZLpEozO
bCeX2YKinCnXs/MLAJSLWm2LJIQwRooypouSuWlP24Z8cigYZs7pL7JAGSOEZvq9
f/DEwQvfW1qOJDS4vp4BYn1fS+fc2sDW74DK2Mzswgbq21OYLHBrsZTmKiDRYFrT
qGJkFH7DNp1Bu9n2aEwLAEdviVlwl2A9m4GrPKMpAjEbOhIYVt5oVOj0qF2gIqKg
/WnIoN8cvE1fDAhEdvSfSu0zjfJfUDeTeODGi73W3QcCYEgCFvAFo4A8z08OnXwP
Je7F4Wi97Fim95s1MAaA2XgdqBZZQDGO6YqZaLtaaX7K9lOEZznczz65bqm7DaGt
+OBvXAbT6Vg/P9L4qUxTTGo8z8h0KpzwzVp4i1fLzqxALU33CkHk0aRLXz75P8P3
clBagRgtFIVqqFWvI4K3e4IjZfUhCRAYz1KFJeTYWjlpEWZo+cSrH7iNOYkfNqkE
`protect END_PROTECTED
