`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
36FfbdoTGAZVS52JIrtIBcLO8AErJHH/3fAAMjHrQcBX2D4+7h2dbqk1T0RMAupm
LuyfVfQT1iwwIGGmxaS5xnmn00mTAW2YbJyYd3H0klaeH9wvUbjry9RDwqfybHZ2
1f107vq/WoVaoVjHpZAv4M9pLhNTcXbW/mk75yHPErBGI/r3qZ+Utq6VnOE23W8v
UcSvHnrzXRyIicQAe6er50IA9gNSvERi8SLlRtr+/22YStyBBUj5z/LahJIkzI14
EZvsdlDWVANJ/4RHKkeLoJg7xxVuVVcs8agVeFeH5ZGnXDhHKHi2uWSM67Q9sOtG
KdR4D0aNLW1WU0/GweG7eTyXbB05MTubxUUEk5qfZ9qGqjsvnbyIsw0IMwRAhNvq
/zYBx6Aj0yyOOMTqFV59pk8iKFG55KlWlhdTOlIa1/5fFkh3oAgCJfc2ABaYb4C0
4icsEaPFOOVhXZTXIt67wWHqkmR9lSyzyBJp0MegZELPH0rDGAwPgsisdJzpuCRn
QGYzi8YXav+F9LtZ8TgbA38cE8/+a0UaLPtxAg3SVdKEZ5lLcJO/72iFBNcgigkg
sGwtML86tuDDda9zccDl6v/Vp+ZW5KPEOIjVGhGaESrJW6NuOfvxDNHjXYFr1cjD
Ch4zjg9Y92YIpmx8wRUGxu1SsZDDk57cK7WV4gC/Ofrw2aGp7VsZeeq9xDUmhGCN
QVWg3AZj53gIHrMRfrGFDEq4EuB3Miw5MHDfKdvztSKV91TGg43QYJW7mbmpk20r
81j4p0SZBvMruIE2h2Vx4F7nqBzRMoqEl2ilkscNLK0X1ry5eHs6I6DblaWClXmG
2vWxlqvSxDMpFEEm22/8w6mS4k/okoQxCC/57ZA76sSXwiclqtc2T1t8JC3sJ6oR
2xkUWy4M7nYf5HKhkmUayKfENWjNZ88NcxWE1rmeORZEOz+mg7fPSCniwkOM3MFi
ybLciGYnBJ6PWIriM1GalKdnP2jvwsnpACHM7EZh4KjuB+o19n4MwH5ro6O95tzJ
vPG+cHCBNrFz2GEC1OfPYrbCYGKL2VPm50ewS1i7eMU=
`protect END_PROTECTED
