`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z1n+0JGPKOstZ/SiwoE6RxWmLOkomcHMYMKYRHyaCj6E0o1ebypWcUE8rq7ATS6l
2x4fDJ2jExQRRR7Azo5uhyXuvW2K9qbNtRK5T9VV6VtM6WOI4O4e+uq4cWwMNu2c
g2ocYWGiwxMtRYnzTKYIBAcAKPn5QL2d5Ulfny+/wjpLuj4RuHcUTv/4KtDhCGg4
emEQTJhH1Dx1SK6FsmmOv6U4MzjIZXF/l3he6KAcgJnjlp2ankaWwHM0CoIcw1h0
tP0+tbssY39AX/1Xh146xfYTaAGrFMZFyxQJzioIN1pvyqyC7etch/mNKWcW7v06
iuVUgyTAjW+oYVwH8P7CCldDZ/c6QlMTvc/6NrgWsvy/fZdL2+r0iQ3kG9x3mrTY
Q6adT9Z0oEB4YMmfvtSOQBHwgh7qOmvVltZ+6YfbUc+Suex6BbU0eluNJyNZA5v+
QOdE2mHQJB6d5tR+Wt0L0bRMWsNWtMxQnc3s5sT9I8m050TntpBtVVzg1UKzM1lS
srIv326uOHO3gNfknXfldN4oXTM93m4kAOrTsNwtMgFFlaxCvQBRQrcswGB6OjBx
5Vr2IGmtImSsQI6OUBPJfylBlJcheJyWdkzS62YnLt/GUmVpOOuBI9Y0i1p1Y8EU
w9XSH95ro/q1e7EvVNaaKudyRaqjXSjzcqDpnAgrg0fnIUikYU8lhQn2PiVu9je9
TbTY3J6JfNV+Ly8ZL+rnIjSH3iD3lKEZALiOzR7iTb2E44EZ8O8t49oR6gpch40a
exDiuFWHRyNKbHVkZrGrGGiynthw0dx7gEA8dHfIFPyH29JV3yk9TszmBo5o9Mjd
ymbT+Btug5rvcEdmLq+76u4jO110g6TvS6++GyP86T5z03Lj1AAvix3KB67zUqwL
Z4shmdJz/64L6+M43HJO5LWgFaRR/nhK/gH+RYmW3HzIsJzbix/4oxMOyhZvt4kG
`protect END_PROTECTED
