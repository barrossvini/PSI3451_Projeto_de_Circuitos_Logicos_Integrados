`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vU31rMaytRJqeuAxZ473e4QeBZ21twbhsqJ+3gIxQBvX+KdFNzSjTqOTm5PZKE5J
dB8X0gWalYKVOPp//5Su/ZoCjTkeZn3LYHExTitSNNLv4w2IY774U2OdHOokro3w
pr+A2/eC4PxMzDsFWsWvWLxaibhA0Y2oGrJMffhhHmbotbdgPWlwRBLjMmR7mJW9
N0jp3Q4NQ5sunbWEmXHfC65i7+4ejI+X1kH+bKDX2ZAAtJtu05IjJw6sQUYsTcPi
rF7+QscWFle7b9vsfLDYV5rudNn7ztWvUuRFDj28Yk96eVyup6TafyRPvP/rMtHv
XNpJZJ5y3DGxouujlwLKWEWoXv63oQGNsJfgVcqxQm3UqvwDFt1fHP9yhWf2EIAU
cQcRtGl9vmnxnMGeZhjaJn6H737j0lZRurEu43TGwQ5r3+j9Ztsw9R22kN9RAQ2Q
r924hMKiAy0cZQjBOnbZP2nBUBvpzm5HNxK6bmJoLe/EKfsYSisNOwXds7q0Gps6
vJhr2SrfpZSwxvUb9yLEAR4qSmejnfMFZCcUoDTdEGC2zpjui7FoJCAwiBqnou95
fKTZ250KF9zOgmleeWGSBbamxU+DuwmMlLRVbe6B1qNeruukXfmrgWGVAw6FwxNc
/SjiPWZd5JgxYUbHE49HI7g0a5R+m+7N1VM0ynJChew5HsxKmc578lUC5iaqlLBH
GarmiAMRRpi+W9OcBSWSTJtITVGApu86ff4BYT/vTeFM9j17Dh60JSN/goUCvdmB
jc/VEw2CDCGVv+6cg4CBdih0ARPiJFATy4wIblgXvm9HPLuGWSHt71FSmv0Ru1Mg
iHc2bPVe1BwUKRtLMqOouX6h+27dbVle+0MwyRCn1NfOzrmfVEEzol/ZrDQkPO4u
nZrEksY6rlKUQRYXSO5A2AmZqSA1an9MOfUwbtIO53Vu0gss+GXo0FQYZZZEhGYf
uk4jetkYd+urkX35kvv/H4UZfhyWKCJ3mp2TBbfYlFsP3V38EfxH6MwxpxdLFNLc
cMbpNmDpWjeGNlNx/1NNbc934KfO5ZdDfHJViPyb8KIRQvZtV+TcUHer8zjbzfku
zpUS8NdbnZTP4R3wR7ljydYPvy2beVQhZrh3yvzn9xRHzPcpivJFD8Q56sc07csN
2voC4bk06Zm2pAmsdkrNLbIoAbemD3uehImaAs0greiylJSXOo7SSkXTI9Zi7PnD
xAMz7afH+ZbYCL1I0V5s+/6gFuAXlLz/ZncHrspNNjCStn7yvba5NeKT/nz75rRq
RLHaj9WqlnaFwcCAGCQ05/UKs2cyeWwQ07L/SIFDc4Fy+vFASHhUKWSG0DKRCZMN
ehvlOuvRXtFi792Hb4gok+DFFFXXQKhCpc+LrrQJu3LGkVulln8+huTGbFohO4sJ
iHFmBCTZGVjLjXWuLU/7jrygn/vgl7NK7fYrRNnnXSMjZEqIHFGcRR2KwEErqCXx
+6VeeTpYiE345gIpGg58PffujlhgKwjdxGXY+lx9ZYFPMkeoc79d71UA5HAUmQAB
5kFoYyZxjqF1X89GhuQlPcQ+9indK5jf0fexV4qV6gmc/1xvN8goUkt04knvwpr2
xDqvp7WFklLwPKWKraq3bMGCROBh1Qu77w/oTwMow5sjAT2ke98cdzAcwIvgSRXx
shvPobHnPbflxJg0pfEdxm2wR3PADKFXdO46VzcFIqe5Qj1rSNBQ4bp9NRcEYVZK
OrVfS6qlsr1JItb7TGt7OnEAlyvJOQN336vlOBRZYa5h+COAomD9QS8AlWaNyMUc
Kg/fRoy7ZY13dTRc34RnUGpPuXiO/3R/Ba0zN1xqvg3Ncg+QrXEXcbp20oJ3cYye
67fmbd2vKq+3m6G3C9VPtLctU8N87jKaEgsZTxu90SbAKpneIwuomIST3Q4Py69C
BmjFtI8/CaZCn+UV2rCYFoUauFEL95h42DIdb5tEU3RwaXHJN63FhzvM4AulT5wt
Z5S1a2XaB6BXF9d6df6RBYW1AUfYcUOPS3cFFIevyB2h1MAJ4K8imlqqBdDQOGNk
yNc1WHERonGdkCoU5KsXkf334htcuSkZymatz/ZTHU3obzOzB2EL+3tQOnvR3cXh
p3xgkLRKn2Ggn58bx8bjRsnwAdE7haNbjpuCBCS+ZVWoAbfoRWitawYK6l2tMw5c
yHkrg1iydHjiLDM/TEaJf1HPRXHLl5bLm5PSuzL5y9pN35/2ZRguEaUpaA+DPyGj
ozvxW6lxED6tVV+HFlI6nw==
`protect END_PROTECTED
