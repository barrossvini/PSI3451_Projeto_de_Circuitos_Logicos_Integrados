`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LKS+LMq8v6/9Tob7GX/3e5c05LVC8GrSn13iCGxOR7Pw6rJCj2mTNvXzVrHbHByW
IP7Y1bFVNU0vPg2WVewStRe8BheeKcYohfzshXtOzzrdNmazfq7GRYC6ecYXtr8A
PAMJ31SnolXkegk6DjVF7PfI9Tuwc62u+9sZ2HQLGdQpYUmo0TN497MR5YYV8rvX
8IwnPN1E6oEV5bQPWSVvXdQhWxmu6dExsA6Phq9cxxBE7HPRIyd6pD1Oj/P1yzHW
LPJiIV+Sh9GRVKUjB5bttFqBcsSWAP9mVvAkr6zDQgNs86ggXbt/n57A1VPeF/xO
yyo7Ue19PrqmHTaN1Vr9T+PJtp69vmi64d1Fr6E0EgBr/p0WiCIo5bkqfvehinsB
VQrBJbkeucstI2j/GDHY79sKGYRFmudLI2wQ72Hvh64NEOY+X/xniyKHsKKYPdWX
4XYXKMNdtkRjBbf3uke9zgMfwRK561+XlnteXi0yFoMmIsLZkOr9sEjWcuHbzs9r
bRY48llx4134hPHYq5RNQ6I/6ttG24W8CctNMtmMvJWd2zesQy9RIrCkS3MSMJ+A
qWBn3vB7GJZwMouTxrDk/U9+JmxECW8ii/W6F5GxxbDHql6yj/zybfU8C03VsSYb
YF9aOsrJTNqUUixhGjK+TO8G+NKWeLnSzHNi3w+trmcARQMZWvhFZwpHKpOLrLl1
4tQqGejvvPSF//4E0g78cIzTLYQ8kcJId/tOhS41PDkBlvhK5VVsThgIoHRpildB
dGMkuDy4Ym/YpP8CBnFIkwok1N6gXI/D4iBhWEFdf+Bsz3hSMW4zM47RpT1HlbMu
FZl7O7k+Uptyt0D6V4uX3DD9kCejEzQl4YlF7JipSN0=
`protect END_PROTECTED
