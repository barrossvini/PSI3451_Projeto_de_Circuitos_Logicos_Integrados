`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CLBCejn0mxfdvMfRoW4UGZYtc1Pbpnaakr1WgG1OERf4doOcGIBPw0v1m0pfYqU8
XsE5doYtftqL7vKV9aifnWPh5Zc885tJuh2F5jZw7ZpTPemR4SxD0x0b07TTRshc
+HW7+qV4s9svi+dPJtcyDJ/gt+NiE9CIoLyweY/z4i1UWe3x+u91h/QF6HkBoQ7u
QFqm7gmJM8S8wDtuhRTQmVJntCcHFJOv/qnVBS9Lp93LYlqubcmvRJ8XJbvvIq4i
4eyQ65dwALHQZhulsNyIC9MHFZh3t6D/o+BbwSDyuhDd0iwJ8jvKAZc1Mc20o53T
RD5c6AreWpmcq+xHUSR10qmerIUV9HBUUd1UhG7ORd57QsI6kRMKrfjbTBWCjECZ
pGeIjyYufyRfCKUGhZrkddXanwwWfDXydbOPK9jG/jEmrt+NC47fdNHhRK1iqQJi
ggIjgAsTdPuTtZtO4NmV1AfrjJ07euoWtXdNe4k3nS9UEBb3ebZRw0x6BgGfA0z3
/QKU3Rw8vQDxPmXNSS41/Pwz4yuF9KtC1StJfYLhcSiVY9D6UKAGL4eT7gEgUOuQ
N9PhAuFfPzTiPFbic/NmK6NX3Np3wSowiMlIcKa8DVNBRZ6NNnWYNDw565I7M3cp
wBmUtf5iI8V473PLlM9NSUsIW5XBSWeR65GviC1GtkRnTGbYjZE7vifc/ghQbJFb
QqvXCjB+9rst4zBLkHNzO5IglVodgbh74xzAlhGm2iPk6n+rOLGWE3rCPRarTuHh
hwhf8KlOis1opBpGzyWbwIDVjqS4NKd3rBVeqot162kCtxsY9yQoBZJ3n+78S7K3
ajlb7hs9RAl3HAdPJbcjNQ==
`protect END_PROTECTED
