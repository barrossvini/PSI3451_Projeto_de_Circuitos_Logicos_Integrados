`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jqllOtQRcwKeBRTObC1nrZbc/jwgTkKJl8t392ovtPm45t6Sba88hxe7A7vVLT3T
S0pNb8wAkHX8ZPlQygdhyt4ZdKmM1bEicGcsQFYwWhmqPJsBmyNJakuvJbooWk6m
Zua+wIi/TPFtNEuD5l7lBNl18YXC9dy2cIxzTf4YDJQxWMs0jk4TCxVDjfIIMaxR
nU7Kl7TcmbmVVyXLo45f2dTHbcg1EO5NyZ1E/nGfO16GiNPJliEbvaQJXIj43obt
Zkx4t+rmGdUdxM8BWeyCz3UizJhTbvI4bbTxk+xTVRS7gZEvbYGmI1eFLSUqWoXo
JQHiJLLEpZKtxc3gFGODKiBptYONuG7EFbjh9AlV4CuHnJfwgurUt9ksAXPL/+qJ
Y0ovPEKUwkczb3BgrEGa9nWi1q4XAqtGh6g7poLRbLGTkMQE+/bSuY8goIW87bfp
3JxSl5XiifJsuu9507zXukTBQ+OzkVdAABaqDmlsrebSXU2OAbhnENTE5Ezl6Dfa
1SqV67ZP/dO5MhSQehSVT6Ke4ZFG7flmZEHU+k3qGcLdTqItFnyQ6T8lmZ0hvYM/
AQT7GPAcdyZU1KDeOJCFiu95DV8X//YtNTO6HohIH1W0gsntAoTqct6qCuBoGtZD
pEdw08UgvqL3rQeRwR/pKx9v8GDoqQxRdlbE4csq4qgajPXYReABmB2rRuua76Rt
qHmcoDbxUqJ7dI+DWDE8vjtYYjKPyXdvM/MkmgCsAiDlBkO14me0ebjYrNLiydu/
KHG0qLakTuJvRMEvYFZ8L0ck2bM+Yb9TI7wdTMBERlx8XkHF8u4n9LEBDngwKJX+
k2kb6zAJ33OIMwN2mgE+8E/UOehDY+dtmUI0fbqDnMAt/IvLIdWwqQkPrwogeG/t
pAbPDIu6/QBJY0aLopaEOSqaiE5Cjg1Qov+jSk77ql0hqechIUd3UKKY351/7VYo
Vh9Csk8+rlIq6b65iKb6m1tj39b4O+Sqr1LvzqHKgLVMRcmW/qucWoCOvmOipK4V
9SAKTyLCmd7/dNBkJQWDBDBIozUXkXY/WghmwrUW8tkk38xl/VYNd6ZwdTuq2UlL
wRtxMRQjYP5UXRWYAAnccXrfSOVlpKPDiJ1K0bzXYyFcZGukd9KjvVc36yr//CH2
VJ4HAd8tQPn8GRyyXlK6MVLncNWsGUkrL50kEbRYmFUV7Zp5Mk4ptvRmm9+Q37Pk
DaYQ8Y78SOaFEUVHCKMRRRbCPuT+E3s9I/QlQynbHdtA6ek1nPiGEqZaG6KIt1JB
9HiCcarwxNzpQwqpbt/tZyr61BcmJIbtAst0WRNEdswx6zG/pDTBWD3hvTZ73rm+
jeSkn757OPEqHW78TpHHQ61/6cj3fNcskwALmxB1dGO/0znPc1a6aA7gE0pGiV2P
KCmtnmt2XBo6ckPo3O23fSnyQH1xZZE8uaj4jmrqapVN1La2LdmdVQ6l0G7mQut/
x3ncfV5B5zfmlNBRcGRZgrrTjKLIKU4Mrvcr/gCTo3g=
`protect END_PROTECTED
