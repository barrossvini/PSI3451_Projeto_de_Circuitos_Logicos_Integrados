`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rstAhX/sW7cUFPm9BKRZF02jJN5a0aDbpqmsUmQyqkYpKOuOSy7Mt4+ImNLOWvqK
NcHGQ8nnzoXM+0hTgceZd3fH4X8iRw/x9PB1s0GOtJyWe6ecTQqP5Y3vmPKC69Ul
WPc9YGAYDASCwsEhnnKYAqiupuavd0h0dWrqQrB3A3Hb1vBFayEQe3gxXLGbasjn
iBNyus70oQQvtP5zyVJtoSUOGQHW2Pq1y8w4GqlQ+7vRsPuG39Q3iBuvvjDf4UWC
aM42vePzy9deLS699Ic3qlgJNqArB/Qq0242iJen8NQlth7ZtThZr+kYmFZJu49B
/+fkeCIskwZcX/WrRsmgrjtsVGJghhw4posVowlnqWGOFxHYAIIHY+4JO40G4Pv9
GDWtSkdwHateMyRgQVgjYl6rYeeGioxqw6lKsyPe9JsQfp9IHTUKC/U29MYf71ZS
4PUTXFM6Ea0AewDuJ4k3z2OyJzDakEaOA2SqEvVcSSVvOv1qEuXoXtpIqqPitn7P
EUuWsf5mkPu95YPY9GBBi24rdVYqAmsjdruV7gr+voWNjvZx8ln7keslh929fNBh
PgMI0LHfRTRuBXaHOviSL+LwmfBV6gaUcMLE0asHsVLncK14YI2w4E427EmUu7ik
6+Jw7PyrrfbWioKXnIcQnvo9fTN9PyLNE5O/RY2lZ0e8j6i9GyT3CPArzwt7LKwG
ySlnTwRgo/+QMEPX3UjV3/4oTSDQuV5nr/03bEWRyRcapHbUx2NThSGNTEKkeimr
9UNSZFtb7/T7TmPaM2RDtAKiwdjTh9H57lhFI5gam+5EDtGNYI5qNbW8yHWyqcxB
vawT7rdMbru5IeaU8c348CBmqgzwtamyGNMTY6twqIY=
`protect END_PROTECTED
