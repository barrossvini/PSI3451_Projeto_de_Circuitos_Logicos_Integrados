`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i7DLIP6JT0Oz771F1tEZtoUhTcet9wvGGFj1JNFVgOjmKnfXYjZHlexBA9EefJtF
yQWwfc50aP6MFLeSoypLzskFxR5jiXPnJ0Ra8o4YaWGv6wS7t6RwPs6wKY9L2Pnk
ouww2nRyyVappX38rqf0Z681eLwD+ROEh6F+3Nb0bixDeCl2USqs9GVFV+AVOB3X
IzkE1AhVfrP8Uy58VAiO52oKBV+3Gw2K5zGDUYGwfH9ecQPUHOgXsiFG9+h1ffTr
SsHGiT8S4H9u5ymqzlET7dxJjfL83FZiX0mvXFycxZqNiz+eeLLACq6dRt+R/eo5
VS2geo7LP5fiY8IoEvaWowrQEIL4Hlvu1AW1AurCDKEodlgRPFxnJJiBaZOe3jd4
Eh8KAoDIF0CmuUAwILkwsLXOM3X+ai87h3GsdTmxdKNKdMHdWJJrE2h5VK+HxWLO
GnukmgdT8zwzKvmgXALrJCAsqXLInlHGnfprEatDi2BFXjHsGOkoaO1Aa2UdJv/Y
DOp5UGBQtK0QrAbgjzhqnCHVvrMUZMLoPZo5HcG04c/tLeyDGXBWCWVcyarqLOac
utZ7MeyHuNgQzvxDzf2+qRNSjd/3jzv17yCxNu1XgXdN1Ej/f+gzTmYJirUwyKEe
k6+iDk1GipnGaY4fcwCYegukJ4Ex9kVNQl9F6JgGz4xbG+d1Y/KF8IUNx9FgTUCT
c0OGQ+Z3koTYv1GRBu9Wy7mKKIRpss0Hz14mK5Jpm6SIybkB1v5I1ja/9MnOmy4F
wwYxNg0sRZzNnpSkzxt8HFdXVOSumM4p1F2APKykUdauYa6bBpVTB7gpJA51R4XE
sDKesmM6rEUfU/pqEQ8LLXi0bLe7A84i4dxgb87aCDapnJq3ELA2+CIXQvk9Nw4F
ZDpcBYC9YchqlYEKbt2ZP2U39WGRDbPxWXJp290j1YVpy9PjoqYOrqsrrkOKMSWr
CA6v4EwAXHglsSJJH+UnqrorRYhANwsV1TbGtCrJdG0odQQcjLShF0TyMXLeAn5G
EIvv0iRsBtsXQtGNLTHRv6kSuCch0AkeU0zuKRlx8vD0LkzpDSop6rkxZii4EQ/L
Bd4N8bxm4FO6HJjCa3gfzysoC0M6m094hcsbqcBdoHCp09YjyyYg1rwqlHgDRHc2
wnSnVDv6umbD1rhGXTbvyU22QWKmOGpx7a8XZJhbsWc7Pcbj9ptO7bXbiMbmaFtv
LAPn1aEvjjt2gBpHZa/NB/xI2rol/aVzEqySu+7tjrM13a9P0vga0RTNjFH7jdGV
uXle/wI9hkV/E8bTTAS62+kc0faQ/AuEwovQSQ55MhUx8syqFRYkP95HM+iXz9T6
HRc8IhJKBkEbzN1OvWTMrC+LI6EDTTbQ4it7n7Xj2u2uebq1qRZ4wSqm1uit7nNW
OE1p5IawfvkFgTRU0REL/ybNdgwy1i9UrK+59mcobJdYzOCAXXzng/kdGIGc04pA
eD0hLIbw76XsbeEw/AcToeNNW5li6illnRNgbDxbtfwj+zljGhMk88tDq3wy6VEl
7Ek1dERQtMdKbL+hABAXNjY3XFR+YsuZxe+QodriZLhzdvruCLcbFqyNRdMqOSG5
Q9zqWu6jSBS7YupANX0AZ6nHxroxU1pFoX71cdAXVXsU6wcgmMa5YwwGoPnfWcT0
yiyY5MSkCl3GJRWmjwAOmnEc6aDjhQwn8AQ7BTplN3djUsy06qk1eQT1vdyzSxsg
fUekdA2uw9P68aHdcbkLbAa5VqO/CY71pmYJqZsTVFvqGkCCTWhNK0toeHbPFWbO
Fiy4opT1cm29WpgHoPCbwQcTYvUf30DbrBbDuscP0PH4CE1+XrhsJpSekspZXKkO
nLzpU0a1FhgGMtxaeV6y58qg43c9WJKRFW118Mj4ZLZChRYI3eFjSbIbvpMRk/Ex
24w1zS/QphcocAU2bOd7BNSjQ9CjxHfubvMb2ik3zzsY3QiMV97k7IbkVSJucYpa
ZjC4GFOU3vaTnqSVcQxAfrmfq7rbyr6RnTEaoVsWigIJsCguDh2+8AAtCl+0PTsh
gfjXvGVmVe8JhKv/1bhGJil7Y9NQPd6mqpTYkuvGs4zC67O0j5OztnI/WFj8D6PU
/2MXm47uVV6Mxe/vfcuNePzGdZd+/J1dsHnuPmTFCtAPeEgSWIvDj10mbfuNYIlI
TpmyZ1q5u1rcdoNqIk0nazyNFXkG9lLxWUzXmWoVR2Fi3IGkL0qQMQ8W6jPHbPgj
uCMlSKXXssi+vNV/Iv96Ri4CnsVjqRSO0I/tRTc1RShzPRcmOw5acNmVcrE0Dkvv
9XT2HveIA5yznNC8Y/eewFs54rxQYcuQndcTD2dyBYblkknJh6+uI8syGli9H4Uu
jytsCjgLfIYUPKH3CMhNzJZcmb1ndyw1rihCZQfQhdQAca3lk+HVsx2eUpqp67aL
u0hlux8JWOhzNeRsv27hbAUOMOEY3Iys9PgBbHKkCKpucNFal8PrwM2utrEIio1Q
xUOaZjTfEIKgcCMlQImLxV91Pp8R9uKWpXgAFqDOLWEksZSu6H9KGwY3RQkKEzkd
xjItThQYmZqspUMXQsGg1aVaRzQDmfSqIMpwcYijcUZoKoWEiymXjCX1xuI5hxNU
SXCNEiWqsdB4r0MX915MJqPwZ5dDIXPByYTm0Af5nznwwF0WEKyxoGO5I7PYaTFy
B58/0nrgqxtgID+dzN/ay/922eDrfQ9Gdcgwy7kvT7uvVZ/xDerkVgYSdI1UXdmH
zwUpufBFUZbepG/g5HVdWZSrtiR9ijLgs7l02ss9rR/FReW2mmok4L7jKnnFESQf
SGGBcpsfKd7mFkrok5ZbUpbiAlRQk5W0i+F7cwLMGMd8FPARdAVshjEyERaE3x6/
GQx9i6cKZoAV7w3mx14FZYVmdFceLLeQJT/nIDwsn9Qw5/g1tRG5A7dOu8jcgerU
1P8QYPPb9cUvA6B6Iin5HyG2vDe15zlNapteiIlPdfM6su76374vlxk4pXLgeFF7
6UhfR+2PurOlzjO06rjtwvqcHEX5I4s5E6/Kko59kQkkeUs8rtYJARSO9//8TFud
lKS8riLpVNa9djSGIOaicDtBsxvANziaPnGQfJS6MGO4gbdDzFg+MZrGA/1Y1Nm0
NAKjy5OFULD7O2E971n3+KC+hsMRzd3BjWjHPMaxbz/bQGTLuZDa/dLDwSMNToNV
WdDq7jUeNaWGmTdLbd035F5HIAN064H20+Amx6hpQgDmL9/xWui5GV++ZqMwUYD1
AfPax3PUV+NYlS9W46PhpEM9+gPF8DsTuOT2Qi6HHpQ+MTThSYz9NOhNZxCVUgEP
pTzEBeh0Mx8mUnEwKXj25Lg218QygNeFLVy1oQPNi5k3+JopxE+6c6ZCGARb2bPZ
i3QmCC3XNj/0VBniZEyctYGLeURvpKC9nuxCd+3rko7abXiLbgSAXU4Ev1Hr07KW
VC4tGLxoduemwQacaXyzgp/h/HxV8LU/pSuUFGzuMTn37LDpn4eMaN86rhLWBX6d
u1rwn0wisA635kbBaahDBd7U/lvAnni0i7AT1pdlSH7Hhs2GAKWhJGhzqHPOCx6B
cFS+2/TIMotZI1RvTYguifL1A2j0kreZZL2RgORUPYffglyOv2aR/G6yVDCmeKby
AL58S0tv4XC18cXx6bpu7icbCOG0BGcYPuXbpp/8kxT7UZBbkzLFWN2422CgXaZ3
kbOFVa1yiJPuvlZyUJdz9UvwVDdRxLpnA4WgqtsmhWIaDlL5oIQ8APybc/Y+lsEn
jGMtGgOdJB980Ikx+KY37H6j/6Qeh6XHe/hX4l1NwusKJ7YXMnrS3YvwbS6TCL7d
CMpaZfJUC1O6BFtbqs1q9wYBAapi1gSZY8NjhGzSqSVFnWcC77t3iN3Cel7XUSUz
iXlke6MFWWbLCCGhsHvjE8GzCHgXrVsKe1xO8UzKIBFVhOXPwffVQQrfRmFOWdSP
jC1PNryWg3ZEfMGdzF14/q9gZNdipAai1ptB5TvkTlwuctZc1J+Fz9dFQ4/+k9aO
0qYWYHm2OUcdDhfCStWXL7S7shy4rvvxt88pB/xI4JujTCAEZoUqNFb5MEfBhvVv
eRnQyWQk3vR6tAUs7ahqJr9Q4shVOK0eWtouEk4FcijxcpAt5t2x0BXF/V0P+9Of
qS/LvaP3zz28y27mSSPMPToFJOqchDqRVWmiGAjfYLIq1pDM59t7g17xxay02XEY
0fnqSi10zIoa/k4Iz1r2pSfYqxfvdc6zpva081f4STwljxOsLwaONnhd+he1PUX7
QxRqsTSlD1/v74k5ODQj1kUCdt74URw4+P65w2I6ADoY9u3TUNG+HbDMF4L9KpCc
06pYm7dl6jQkYDfKwjQTj+nz4SQlwOOqaBPNEBkpoOL5qfvawkTwA8und18R8nVy
gNLGMBT/xiTCb3P+EB1K6wTdGuigkuKrbhl+utqQWF7vEO7c4OAZ2b/JgtfNsSEy
EhO/8Uc6NDaES98Eutt4YJP4ivvbvWLo56l8wnWWR2kD1sZKLQGBuH8z5xvrfNit
42rypqPupJg9xD1Tg5N0giS+PCS4qHS/OJNymu2ER5dWabjnWZq7BIYsHkiV48IJ
q4GJGaUcMXezQTX8j8g37VD4eaFGlImcl13qkayj8aTaKEE1fXTV4MMiRqHSmauo
ih0Dfn+IMap+F+gsaNKXpIZ1Ke3y3ESO13X29vgoG8BO21XFHaL+hPEyYR4/Bm4F
wFmC0xj2nMsUoOT0IT83gdQS4pdSjZ6LCvklXi4ndW4fai4g0diteLh8E8ECqa5U
oiZFnbmNdryTxQ9FwvFlsKwao4ratgElokaIMtC5RYYwO4O2WsYXbykOwg9HRT58
YnVrU7noIKltr0Ss+i84zvaaJr9lHAZ1OTjM4W1VUUlgME9J96ku1anJANddwlsH
ShKgtaVu3NNXnqOGUBpgtPObWkuer5D5c/XAaL1AErspBNSfB7DQlruXQQDSfmHM
sAawPD9bMtvZabzN/0yTtaUVqnn8rscKPqJvi/L240OStgJzm+AVXz6SypHan549
uL9+TzY8TCcL7TmywK8ymAab2xJ1CUN+qj1/dUOsbfXgIZP65Oa7xfAh0dLyvMxh
is/68qjvn0eJOGYBKAiLnjqNOWS2oIY9poQWBJB4Zg1G3Wbd7hh8MVyt40hK0GPK
RccRUbXBrGMBAQfj5Nj4bHpFiDvfEZG+mV0mfT/gVLnDl83JAvBxk8zdWf+XuJ2Y
FW0E4ROqJESM/NSSNjYYo2sWREfTd4tnUbx/U5d007r0MqNWZTDWiowgF3Zg9iHn
N0VYvJBc9LRCeb27e85zWTOb1tUhp99gdSlFaIZQ9nGOAfBw4LWz0CZv2dvqUr1t
1tnLpXPvW2oa4hGmcuvG22Qj3doLWep0z1Uj2fsaaUqluiFhoVfLEoeOvSMmcmTu
FNfs6nOgeUK7MsQxiuTPwaUl+2XYbvevcHbumJF9I76xeQ/+8siCbdydcX3NexfF
1NapUXhzvDhUcG+t9bmXzCaAX3/WRR+NZcvV3b849ZIncliSgMVR9/9w9oC9JV7H
Qv0gV33HdjTHqAOvZ2pxswD5KNPSuWFZxMJoS4TjEfPqcXHSnbPDF2XLpaOeC2Sc
Ge0n1O/GS/AYdYJx5Af+Uo9VRj9+RhnjLRMijBGBFlkP3helmLSxys3BE6ceTPIq
ODaNZA6uLv9a/LOTYh8F9TzB4TTfkzp+MshCsMo+nJ/hvFeB27ojdLxK8wLFaiqK
OMD5uUdlsKr7NJ/MTh+R4NCZHT2ZWrdu3EGpmO0qKHp9LByVTArCNjwpWWfq3pvb
rmzIRG3tXIoosQcCNk4aUvbGxiXu6o9feIMsnswTU3QBhUNlqaW9JlJWosS+0T85
yZC2MnWZH9JaqeaHrn17q8KkuUGh/7Mrz8ugWPzMM/jv+goUzBx0CIOD5BKaayMN
fr8WR2beBXxxbluujNxcoM1T8r6CpA5V6v9cJVGlkpAtWawTzK06iB0yFziGzS+v
9e6Uky7OpFgFzxETSfktaVna9Hmbwu+hVsjtU3agS0phN7YFWQ1Tnrb4dB3BqiUT
wN8qa3dexe5m6gd1EX0KOS3fu/yQ3RvcYLMuUHyPb+XDHW7jkczs6B6MfcwxBX4g
3VmKoaC/M+L6z6I0exl7GoISmqplsJGYrFPv6Wb8wTUe2qOtBW03o4D2JJ9IbLp8
OakaL9xWB02ZvHhih9jn0uN6aeBs03B7KjvbTwvkocB0F7nBQOe76v1awWfuWobL
+b+k6UTUxoLFmyulrxJMO5JLB7FBACEI6ufhwnNVbz5D32y4FnbpMF2zAC9bRRAk
4Le9iP9esCo//cCss3BrpbxuQ7stdv2PGw0zWDrfT2jahLUAk2Hf+O9Nm/LkEuJd
F5OmCfUwUFJsIQscGOTePjc0vMcA8B1sNWYXGWrmnvO93KftM000IXK5mI9yEVNp
7KVNcxQNjkuUjMCcQAisjxT13UJrTGp8b/Mj6akA3QtFz1Kq/OHDWUapA9kI3qPU
hA81h2Kyoz7wxZRzel+xHmQwjU8NdxXj3vbj3sqoRHzucl51TQp9LYAI94hCImzv
ucmAOd9v5/OLDU7nxBT9jwdsoSCyGr2OvQ1Dn+YNzuH9Zhlv25tnfJcxsEGBy+j9
2DPP8+Oaut0lie48jFSkQ8A9bolnSvMaH6w5FhdLKqYGJOz6Q3PnBqsW1FKcHOEs
fMEKv5YnTNg+By3zONaO+ttRKFEn8kourxytpxHJ+DC5eveCNSalNpmxSq4MrzkM
RnYpbLZ+zj4ovGr04NndaYDQJY09FqDXkZNH2f4XVpV6Qk9Vd+LjOmQ4XRTA4orS
whjtpGP2y5KqFCypI1BvEgeh8vv7xID2OIwyjDGcrWawAYREi7Pu1KXbf0DGVLDz
bIGdXDR4jH5UlrDyld+5+V07Sy0sFwVT9AEpH+W4Cxqfd/RruQF7MQkHUdWjcy85
rdoExEqQtVszl5t+5KLEQBcWXKaxcOkcVq+GAAqcHMlM5+ImOa1ulaxzIDBC28Vi
uH48/S+qZ9y1b2aFKxWBbavaMpHFByHHaPhDQ8dAPJwP8wSr75UuYbaQj8zkiinw
zhniMMOuOtzHweftenj53bTu2FI9NLNgCqEJGW5po9mMGl+K0R5L9SozMAQyYDWk
tNsAT1KwTSasiLhKpu5QzNeANxJ/uxtw6G0UojMA+ABZRFU2c4qIAe5sGq2PJrF0
Gkxsm8eMZwq++geh0EE+p9ZgqgTCy0f1N0tZN9aDnPFdLyplt7Zy209F9gJNlYtI
Nqr7XnYOKlAtjUny3wOoyw==
`protect END_PROTECTED
