`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vh4sKn8odFs+BKWWcfPuKQylpoz83D5P6HQT2lDYWLVEgXk5LLri4ZyWs5prw8n/
2GPffeZRx7Eck/tTdmGbM4hZZKnxEknRmRQZnGN58DZiybPu1v3O5lkfhERDuIf8
S6vFK7mFG0SUJoUaIWi9/Jt8y22AocPdHGM+l61VQcr3c+tE+qonCbJ3ooEDo1K6
Wdg3ZpyvpgBptSbOn+r4+sKUA5iXdyk3vr4XJpHvJl6z7P7Z5K/ZYwAXOjzpYnR7
fMyE4IZTlqgZskOMBBU0SgrK5xhf4p5+ss5Xg8FcmriwFepM0Qz73t/tvTZ1sddP
AduO3t+6+wL2pQ87YuJ6yZIxWEbimEe9MFrR5aD7gd8SPFRoCWP0kGvrnXkmZ801
hLdgS8+GuJQbUa7vCwibRI4UoSqry5TnkX7iRFw5fobsFpZS9/A5/ET2aaoFbuEL
ST6m/ooKiBtmdTJxL9+uuzchkC6cSthTxF+7hh/k8gT9oyZT4uoBY/RscLFl7k8O
CGTL5vK2I8f6Q39p0BoREaswCj/eJLMq60Z1M+jHBF/pfuDfaqqiw3S9Ax2DT/jT
MW0Fai5pX2Y9G7tL6nz/R2HAR++/zZ3PEF8wBJeCy3J2JCvL/tS99p3hO96F7QTp
RvmiRbPDa+l1flbsZ7NdylNQ2i1TUgZwO8Bg9xLnwGZ8xK+Qo+LHlvhou3mxdAR9
HhitrXWKc8yV59EJcRY0GYE7666Jg1fgn5iD9G+ZVavKn235fI+0e9I0/LKyHYvX
UYaWC1YWyLbelE1zlOixZNuz7tHYV1o6xvcONSrllI+/qgjNspALZTD40OZLE+sf
uY8wQMGvlkD8hp4K5eowdZc4Xf3nH69HykTs8h7y1fYyfbs4n5dU2ynVBsJbrmIR
FF/p4fA8fvtSj5foUM/XuGXlXjrwb6l+x8wXO4Dzdb3auTorVL65hCsRpQrbBnzw
`protect END_PROTECTED
