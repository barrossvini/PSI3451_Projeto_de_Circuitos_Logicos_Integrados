`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7f7Zk6RJhcJOBhhhzDP3JEAWLV9XNfFAAtxhBT6gQXfsn7oVsJSoNOhv28/KiClr
2cp3p/vUWeTk3DOcpUWdK1sv0SLosbB5ldgYvREeHgGqYuMf10ORGS49qLC/4a61
q2S2SB9TpW8MWiZaYI3Ygw/gFu+8FYQJo8Srd9WwBK1mkYnloGo2FHhP9Vn73CwY
dr5tC2xgq6yLKtzbLLJvoQ8KeIIbmctL/Pbdl4gZbkPpx0IfAeX91dfrHKylFrrx
O0cMIiEAH4pyHhq9BxyLsWL4SYOSI7xQ0J4K/dBOKSpfMhl2ExmjaFgpM/lOD6Mo
JkhXYleuiIogzjHmLS1nnplZ5HgT3V60POgCJ9ernxh0vHVIEuc+4EqRJQWSaadl
NcIRBYilysWQvvOWBVQCRdYhJ/d4AQ6OVWUI6PDXsk5XowSZs4VgtktNfxgIUlOs
2pvzWaU047Frt0/XEc9WHzNUNtYuB8YX8m5TFOYdhMSKXBfSGoo7B2hPK6ZSV3bg
O9Nff6UrqudR9XNwOZTVmiq6XGtPDy2A5ZSmu7BQbYQ6TS5N1kna7dZ6UOPz4XxJ
/WvPSwQx2zuLahou/vzQzvrA6kOfKsRnY5TJ3tTSrgpZAPTChkpeYo2cK9sVVs/t
DnR+iXhzvImyvi49f8z1wJNWEz9mIsJq2yytLhTDEY727TfvNxfV+U2Z1eeTkv+i
jvyAYbRxJoBJSdcMlDyqRosYz8GJB/rSkPM9d4BXl20EJxgIp6fBAl6r9Esk97+q
/nPn0A0fwyHUE2EbqZMlMu9Z89uXkbLwLjPLFwMNEzuG7lgWnV1thEVDULXX5stf
LNHEnT4InILqDT8hgF7O0Ro5SZMkTwVIddamX/RuVRK5DxMgaf6b8rgjxU/zK2Ax
5iMHBpDnmm0PkBhBmtUzhTXWYy8KLrRGPwUzHdyHHhtiDd7Oue34y4CkINRoZrp3
JRDAgx+7w1QRuLf9NZEiPN85n0VaQhgNNXt+PsSs56umbkrh7vHyiyrkVvm6n8ap
we24yeLKK8lpcfjHGigkA9kUcjVzqkTLlqQmzvkiU1sD814Y8Pjz9ZYLtbTmnKKg
zvyUm1rpd/hEFBqLq/cVlExqK6EBwpL9D+peLnnqRAmgUg2SRvddr8u61bTvlni6
xUhrZlekefeTxwT0yvrHDciHHk4+Ptcn/dEBHqV51RFWYp08Ej+tlmV50gk/oC2p
Xt4TxmYZJOU1C9PniMp5N5xSMavlWGKMOLt/tCa45TGplvvTpjLiOudkDxnhi3Cm
SyJijnbxskzBEr5tJbqH0lWN8Zve59KjNLeBGNn6n4yeYQcJw4IoVh73QvpSMrOP
ZqC1GXUMQEELci3m7bWtvHWLjotam6XKMUCgTmMaItto48W8z7vLXsgslYTpmIw4
omQMjjQsYQD/UL9vqGQblVvVAC3JKKR1Lh3lCh123UrjOghFcOUGtqkJBYLpXP+Z
ElM+8e5MQKiRdxfGRqPqqT7yrXF1UDmSvTjisLUemAvQGtvCjtZ88YFme2Wy7ERa
VmlQJqoZ3ZkpUOlvyfTvZcgMLCj5I8iY2+tyuPMlur9i9yNe2IHYanku/gozF9z7
Bcr42aKNPaOZfTFlziRsHNb7AfO+DyXCINkTv4C/uZTPZnOOEWS2k1M/e024IL53
UoLO9K6+9ExxjL5stLSYVU28yuir84ZqX5JrlBlQ/wFGt8ujqa5RaQ93m8ARPKAi
YvRH8oFR/cOE9FwF4HXwgDOlO59nMNOVoONIsQwDhnF+U7HcrNh+mxj5CRfyQ7Fo
qlUmyeVbBZRMsyrgmTrq53KtuFnpxG5TBqDakEja+jP+15lDb7/Tq0aW3/U7Mfiy
GzCXhOhU7uMtQJ0q8z9IRRRzHmYC6GgWGRE1DDXD5MLeiiJ18wJQe+zpuD94a+Sj
EgNpKk1CipnwFkwSc6DLT8IMsUWCRmAGyLSi+QSJEvKPMbVtFN84K6prWuNC1O5C
WJQ9ONAG+2oewvkPo6imqBkEdWkb5RKPI6Ly5iO2JhXw4/j5M6zbybzVHySQXo2b
6huyv5NIQkrQBq5drj7ePpxtKa1Qnc3qQTQmHZSBxNQy8izvDDvYENI+oJLxNZtK
iy/AAVZaTthw3J2Ydh42o8wyarI86v8yS3kS3Tg5OXqAcylFuTOSt2XCozACKfRQ
33FQtMxJhO1DCF2jEmc/OGsnQfoBIvoUgKrU9SiwnxRDWVMOX6QVXzfXnWWVx088
n1+wmM6sVYp/ASjPPDtJDRbXKRBFif2daJamcFrHmuzxGkU2viXs8hEQBoTumzx/
q/d7ekeRrfPq8YkguRnkaHrpK7qT1pUgqp5muLtoJsWS0jLym3KRCvtNfjmC8hBt
3VsYC87RZn9DxLV+B57hxWPIzOmvaICwJyTMg6BbHWZgx5pCvo5nrdF4j61BX+bB
58ddQnAbtM+mF2yyt0oeRpkUv8tVyDvF1Q6Vx81LG9di/ckhMtuVKbOLkdpnWZ5J
8fSQdmUJYE9Ms+STChb3ymi8dxONd/scIg5Gp12rLhfLQ1F97MT53LNuGOOTbPHv
8jsO+AW6UGz2PuS7L2K9CogENuWFSCqXKiYlBirL8INfKPpswtbrH0XBoFV+9JwB
qGoKCQJzm6ajpIy55jn0LvzAZ2uAaXwzw7WjnXyPPES+JkhpPbhcIHU8ulpAl/Xo
oPIsZQujI4BNM+Suu+lFyB9LpYtQyKrBSoccijmXotjI0/lz9XPRMi4i7Wsxq7Fk
Z8/S2b0Jt30SHfZTJCaZHJRO/L/rbuZQPeQlHiRZAHt8OgrrtEJs/2TkCyQ6KskR
dOy7CNhBYs1sgl/YTOU+P6QHKu0FXH9gTDmjD1zACZsJq6S3aA1Y1fabnohHX+Dv
C59l6jnarQ2NkpCObjB6rzN2ubvUXryQwABAKNHiQY8GVgv145JsH43/8jTZCe8j
4VqWL97IrhWKMQPsWtgR9fR+KouHkrgFR26uQVfM77Gs5PlUkCFBJaufpvB7hcQ5
+yckjpoqqt8YdnhrdeaUDIV7ki9H5QVTOd52XG4EUr8DUH/9FBPSokDFCcL5KUT1
2PZT/hi8ALf5/egKH4EqEtcDa6+VMpyyv5M3fV0BORPYxoJxYGH0r4xCiRoOGeHn
yFSL/FixEbJpcTNwJS+p7wLb5s8QVag+vZQei+FG44LLRpIT8lapvmskhEY8gK2M
t4puDuTLXctBtw8NdgVdmbq0YtVp6tC3gXQXES+69/GOmZEfvAGFH2zi82TzqSu3
uucFjp4HWh2DkGnHlrkgMHbMt7wn2EnK4B9vL3RJe1FfwxmsRNAsSSBHODIOYc44
AMs7p6i/SgqMUPpjQP9RdWqvzl/I0p96+EiXYj1i+tYCGnybd1rcEIVAUFUj8YMY
WaER9B/2Y7E6P/3VqsHUsX2Pb+Lio/ErhzCfAKib6iZ30VMGCdpEMB0oTEOLzQ2o
LjIRp2tbtYH6IHqReAsog8yDqQ9ecQ7F4UD6KOC2p9zdITS8moJtECowJSS/fNFH
br7ZdTlDCCKsPQfjyneUIw0czeHGGDIPC9wAcYnbXNcwtWKS6pqP5MT4qfodLXEr
limK3seqkUnYHUsJ4wk7xdqEPyicb4i8uvt77KFJIdM=
`protect END_PROTECTED
