`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rqxz9DjZgK0/txaB4Dc+RSn8maY4+BzrHiZXXNeJSyJjieJ7vxtFVCL087GAk8ds
uYnvv9jdGv6fS91vaFQrOLI9CGDwtbVnssI8XoJcNTFoD6z6S2xKRKktm73KqJEv
dYasH4uBaSRz3Cxsa0PS5s5eGhTAqlUM38WfFp4oLrDzAN8r32yRid5z9HVGjqmZ
OWGydHjU1TCinByAaHCw71uAcuVzlVmKph6NnUIz0u99sBSpCfBa9U8GUcLfphg6
dTcP+IPA0e+W5VH86Knitx5OB3C5vsOHshHSYDiz1TxQCBNGrJgzoCIktCo4uD/9
NziaHCNtSn+CyO55rmI13fY6PesgbEwCzI8FXz4i1mnxdKB+2+nXzOFQ+YwEWhmY
GhkOBKOLPvJlf559WaQ9wbwID6oNWQIGCFoDNO5DytQ5gtHaConBOz7HiCEFiKv5
BgenjDGg8IVvfK6NWdRuNzcU/D57f38u+0MO5WaZJCUQ5YVtdlBU5BeQsJiudv8G
WA8zbccn2TszG48jyIq6jPy4jOau7gaLN0Q1lLOgkuUzTZZQCzHsWf6i6iam/6ED
WK0lhB1ywjFyJi/2Jk2axvbnCxh/XY+a6pw14VOmjuBVu4sJbP22o0pouQdumLxg
ikY64pkH8l0ydVa895tK8hzDmwecX4Tah9GHnE9o7CCLClTqNef4YfVA75APQQ5X
Y2+FeErnUlfYaDh0L6ewVZSduMycryejgY3Nx1Z+nmyRXuuVER9dwDbZV1iQUldq
TEDGNSbnXJJ3JGkimaql7Z05NGnktRLd1ncvDHLZ6yKAHJmjqipoPmfjJhTv9sYL
K7EW/WIg+DDst2BmiMjOqbgNd6F9eYHFK/6zIpvLT6AAw7QYxs+KzpRFWk1EP9WV
dhhl3FHPfEPOcrGQdnHTYClmKdTHsDmyP+16N0BFCw4KVPjZLpUw5jmaZ4L2DX0m
XQAr2vuZYI9W4uLeOoAl4bmYHEJ7yDsq0rYEn6UYFCZqDaLFjcZ9nICewEJrSr4a
4SIjLk8+HY20+B39bduTLVifqbiBGqsHppOEPSFWF9R4MjYr5n4UM1vQ/+GjeueQ
K5Bp31tvZu/JjftN533eGNUPsQYRV7z5mFCOoMcLoIeSLj3jwVBs0uP6mAbtDUaM
psmBPqtM9TjZ6mOAzY9989Qqa4tGoFaEgPeIRmSqbhOlucACXtB/e96SKdkOBnBK
bHvyjFQ36tIkcEJoE/lhOi7mwpbuFeBGQC00ZcrYMecDmyAzzAQW4tUIycwWeMcu
Qvm/VUYJ2uD6AXeAl0Qxd8QDC+jJElunfy+XvbXfme/vAJdHFOxnXDOw+xYdCPlx
ntB/VvljXWfLLS1LlAQLau65CQMwUxhQrWyuliJiWJgreR0PnKDRIorekc6DBGDY
`protect END_PROTECTED
