`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tc4byOqVksWjXEUavO49jE51rGFbvbnZPnHDitxIEa+QImuoELz7rlgIbkZqiq3w
Ni8mrTQOnwUojYAnAUGQN5kQX/v7QExU45KFSJZe96HViDbH48lBdVsLZTwif9cz
QkruoqQhzak806a4OD2qytJFGCpKa11cXr4tzwSL+Zv9zeyVm6zYzEEJlD14xHAV
FZSInYWrowfiFyOcXoHFO7wpzIADGEdBdFAyqWOlB3/a1RYe9d6YFel34jU2uGv5
rnCAWTyiq+yayMRaH4CfLHadWCxZbB8d0IAH0pfnhA0DCUNndNCAtyTy24OIgS7T
Z01M0U75q8zi6H5g7aWwOHr0+ohbJnkawGUkbNsDdQ3p+EeQ3TCHBtfKrb5nW9Qn
1l41qPEic22BHdn5a9YlIdOKL6On/lmmbPdkGK9bWp2fWaIdzX6pIA//sUnbvbF5
DC9r0AxFkCr9IHJteP1i8CakBoQvgOo3ocpLpFON1yHa5lzydjQnSYsUB7u2PjOe
kcz4P9gfiBzVUQ0fDbfaHEU848L31Mm55OsMrjrQzFiQ3isCZZd/kGJ9iOj7safm
aDRh3k6rpg568W9GqKzjPePVHwMRwt8dBgoC8EkiVLIPnVEHV50Aq4p1SYn3nKSV
H/c8N1wol+dYz3iQfXMoC+6pMjBSMXu7GVG7uygDrnaVzbisSpvKaqV3iCnxJUub
yYGxfu7AD1fxSEeuMn2WHwQaDjubQx1IHRkbgAxyoBReP5AC/0JQXkKimY3AMXCV
sVvYFOqN7Qm6ZGmTOXR+07gNmqx+qlGz0RUBmZMafGlVVx1wuYHh/SeOsRfFE1Hg
RX4XKX9NXn5s0flr/LXc95IwIhLXwEgvilHNBNimBaZKWfD53G1FL+VqyFSfljKX
Cdq5FUUz/svrhZSeU2lCyxSnr2wXKHfDjUIpmbGWu028OEw6bRda3gK2rKpWnxiY
XH1Y+qxtcTVlKm5g6sYzKo2Rc/g2d6MIH7bFALEBSvUky7qfrvg4fyUDg4L3wsgu
008B3ixBtRcn4Q0l13ivK2C85cVIS0kU98yiE5CCqiT4wSh850SyvOwRlL2hHtVC
AmHnv8dU01sjgAWWM82bizS5ob9AojzRZbCVKQMAHNvtg85JTI6RxvOVXmQMY7r2
vu2GRouvlbYzWJaEqmL5A+BduzFPgkAdaCz2t1b3moHs2u3Kto4hfne7oR6NY/0L
rObeuEwXQsd5Uo6KKMEcDP1T1YGESdh02RHQWafmUSiH6j5taw3Y4wySVUqJ1LDp
nRkVqZLyBP5URbGFoXH3bgL5mC4/z7grcDL3z+759WHvykXly47c2HC7TrUt/Sz0
iEwGM/d2M76EVwnW1tzlJ6sfu6PZIhLUzB8EIck06Fr/MeOkz7OoSU94hiaZvKHY
U4VfHp5dJILwizztwb4huIL2yV/84qPBQO0YWewmOmne4xexd+Fcm1pZv/qFw+N5
5yXm87aQ7A/u+5Ri9E4HfMvQLITy1VeEA0xPRVjJIRsYMrl1Agq525VT9Kf2AMzT
chf4rGqUYFHzvLEmFhKuQ71mPSM9yxwY7vhHF2P1QhHA7G/lAy3rZFjEKxm0H0qw
s3sSU3cC45m1HxcaZi6kzumrJ2936Ew+cdPlSENyDdcbIRZKcIvBwIRbZ7AXSQmS
rLFL8fEOj5QeyEVIp6mc1uEOvH8MnOr0yuaEj8sIX5404pX4MKkKkJQMLtZhXXbk
jeBD7811GBxBiq19ac8vvsO2EEKe8ldm/1i+cT1JxTT0JQ/P8jTk3NK2xAxffI6r
ZI8TovgFjkNtzBgXq5e0m4ssY10aRmX9lEWvwj9kNxuOuxK5rcyiMxaXGMy5GHi3
U51GjiSF/qoEMuT5HRZTKuQpPIEUtpWHVwBcxbK7vq7DfouPVuK9rBiLN7uc5Fiy
R9pqIKf91c7Zpphf00JrEMZ8k1qwZFyLWmhK7V90gzFIsVWDoWhkXZ20wv9PLheP
Zg9yEQi7jldCXnlWMj4CJnh86UMDzEi3IAxvXlAM/ToWOQ24im1/pBYzzG7JpEVH
VPxlDx4Q8MZ38APZ4fevDLhdOSXHv9cV3Yw50I+65iEZeQmSm6ZRhB4Sa9gY3gbd
GZfiVtowyPZWWRwr7Y5unGUQ4T1vAxvzH2M/n5ouYBrJolcqi1IurcOLgmy/Z7zB
AhzXKjJ119/+jLA2MW8zbbxNuunnJE7yui7tsmWUwwMyGss5aTlh7hKhkbyfVkA/
9deaOAld2sIOFP5s6ZuGYHzXJwBk6DmKmkVpZYOhJgiJfX6os1MJG8O+NKYKM7La
fXK75DZY9nTLLSJT2ZlBRq7Byo3njGpIDsRrYNFJzj+kj8IOGNd8iucqnP2QKJIL
0T3QQg8TjOkYZG3V3VQnho8b3GRrlYLEZ0IGibBUc3rtu/RSeuhRDa9j5Bgm/LJ2
DrX3VJmLFo3zdOwElzrxMbQ47bwcUPxCJzAYTMz41ywzWcWbUWMHUq+aaNtfx/Qk
wY3LoK+2h6XDx9B3wlM6Shx2tyT4ON34lt6n8nhdP9hS7WseA1hRZW/sRyN/Do5z
OfbHWX1IgMJpatvRwKXsZHC1DJVvffrsLtU9a10aScOMP3ml65vVJoiXKFWiC+hf
eFuJ6zhxfpOlqQeKck4jPuAS6jqjOilA1SaqeKTuhwIlJy9s3tr8Fqk7mQH1WnlP
UsFtZSXTPoq6UNI/dAkdPkgWIveyBedHRH3lALeQL+AtCjEdetUyuWsZ2mO6S7A4
FhXKlqChtHY7lzf4zVXY6bXx2rqouACsRGbVheNdvNhSAfo//9eyASuuwSOwwBEQ
TKoIApkJk5HIf8oqZ4cIiLUNhebFYV0OWVK/qzfQ0r5YRQby5QXi3RUdeBLLg0K2
v8SQMZjr8A2OL7J1rDStxddIrCYeeNBLGhNCLjSQ5reJKv7fvf2x2lULt8I5I1pa
WJCcNTxdawBLAsn9u6uZfDWihcTdIFanw+Xt+U7clfocCY28jp2vfbfsq7skW6Fm
bbdH/5dvmJU0UhxPO+rEq4qDgSQeHAoHOq+q4U/QD+Pmka0DMBAuw7IZ/GYgmKZk
JNOtSbPQvpJg1Iyfqi7EgFMdPxmY17t9nml9NPBIiY8JNPLqMPvclVsOIhF7e7AK
9NfhZZWxcvbFCiRUw3FORRCgWJebYT8b2fDquJNQdxePsGE275SURI2lBKMWjtix
tj/KS/Oxd4YV1+YKA2S00pmikbhHtg1ZwEUnhe1HFLJYC9TwPYL7bGb1DMo3iGiW
8DNTqCba04Hbc1/H0NvvPjGKY4IkhbqnZp5/MFyvVlDyim+KTi2yOV76bgmMW+is
WwnVVyKTCtIL8mYWfCMf9cEolUyDm/g8tvfjwCELdFokbz8cuGpIaBGqiQKB8faU
oMtCv/Kh7K2qw6lSTQgcRfheOoo8vmePf5kRJQBp7rPayTuLv4hv/5jkRcEvvwGW
nBfO6oLL4+QzUPVmkeZnJyb8XW7FK2gWMqBaRQIzuS2943xXyiEqqssunkgB4A3w
RTj1+HHXxF4e0eoaogbmus72hxTMl6RV/62K8Mi7KrFPZHd1wMmTss66kS+0Zavv
EWMu5XS0j8Sq/qTY9WuowCSZXPBB/JGZRp3HnctlyHr1gQRJcLujG8nPtdCCEhBB
ipxwg9AjDMsCx7sL+EwGicBWKGcog2Am/1zcPk0Lr+vyZ2U4W2RfWxRpQEOKk3MC
3h8j9GuK2aPSpwkiwizfqRr17/PQeQ2jBZwuXdUzhbxo57j/34aBnIqdfa+6K/Cc
iuOvEg+xNAZNNobdAq+jZYvmYUedr6ps0l0bUDcrUU/sD3/ZX0mfiJiW421gwChZ
etjVYdaEVSAalR+8oOlovRHD6JQD2DaiENlJ/HWbMG2wKNapc2DV7mJ7aJ9wB720
TmQ4wpqNjSJdL63i9ze7NmXQd1PfnQg33HIeHIA/sb0tLbvhO4BaS3i6YqgZQ22t
UHPokiU7agR24ktby5wx1p5NvmXkCCTSFI8pAWnpz8iu1n0IS+J4seNtJ1pqxyAA
bUJ2EviVmLoyHNZTXEk0fGz9xtw0i/pOBp4Zw+sKADUvH6HEwFQlUgWTVtPmP6U7
AE5etP+faJj/FH7QxIjGUsQszq1Aux3NGAEC4+JwsTML+pDRvxnoeCBB20w7WmzH
Ny+SMDPnkLs4YhxnlXgfeol13CWCrEuQA7uZ4BvG0ot+1uHVs6cq6uTdoqdRo7lM
zxvDTH6DN0QbXv5TqugK7lV4tbMyXdjfGAsph+HOvwIv/JGRI0FVm2RP/HjEL55j
9/bEHoi8enYVvnUaHQ0KofzGzDqDsqgDXE8SmqLFiKarCrYOFAKQ7Fv8eUJRIQoN
yKujqGPQiwVE372+BExwI97tKEOrTynZrNS5Ug01HQWM7n7duW3C4qwYpynSxE3r
fxxN3gAMS71dyIGTZ/6ZQjOafgPL/zlR8BmH9mQr0MMmHJP7JS+mKWCIkxkCB6OM
UTaTYHptIyDKbWxisCkvBd91uaPZIR5SekBekrWKB2Uywjs5cZzsNN5SHBptf2Nq
98om3wAmwS7KS/e2+sLNq+bHTbhJSr+OLww89oQYtXbQ/8/KMAfQ9KbFc1fwGgMR
q+CVaUvVHcPjvVLMzLRptl8YeBdmhhcK7+B+QFIqTpOZudcwiSR/bqbDUBvg8m0M
p0S5mVQQRXIS0jKwAWdX/XN0EqfStPoHtzkun4l7PnFJuNPtDVzHglQ4JFPV9YwY
oiOBkLTet25acqlmzlkh8LTzMG9ODIMYZOA//MSgSE8Zyj092Ej+clD53FyAxa1p
EmC2hJqFlk0YP/1hUY2oyTUiBMT6cDwCVzA44wvGk9YTwKFt5ANWGtItxuBkjxeG
hxvRbqlZwgJyN07vldWUtBjeYYqDz1S9S5AlYbMyonp6AeWNXpHVo+S6ozDiCBI+
Si5enURSQv4+N3N9ZWPiQuhNaR9C+I2BaManJbu2D2Sza7/7HvNSU7vrwPBubV3B
z1yFyVnKWY3iDp0RytIBDTJUPqFbxuUlEFcMQJvG/05MfgM0Wck0HdbFcHx2G4SY
0V0g/fIvQ6WHwUF5BVjLI5kWSvpAZZCq7PQlH84xxut4R4zlDGeBV+jUEzre+lKN
Q1BZs1zjBgDaeW9eI1/c1RYe5+gNLjUAIzTDz4kz6z2/jqEbIAd6z3rImS/TMI2s
GbJBm5HB3p5By79g7I0hwhHNmZRgn4Rm4uHCDgQToFFhvURh9O8tMqnSa0J3+DtL
e2UTCjSBihhPIsRqnUSD5+ob70J/W+eNmGFJio0yHckauSZI80ZAynKDQvyEsbka
9rZz3KIrpZq+oMx28rX4ETb+keIKELZRnmk8gB4Ah9jK+/fGTgzUC29joWqwukHz
HDpxD2MZ1PMV9VYpBhepmsr0ME5PVwCZcbTFqjPf0owyUUB3rd+DfKb+E77DKGU+
5HVKfxSrrCxIOh4yMct5muIEoQIVsZwRcv+/jk4kVu8EHIXCBB43L6XKMYw6/tTV
qov7YmN9Y35Y4K84DICcDKwG8ODkfdkZQ2JpIXCuOp2gIUrxzPP6Foy+thyj6l0J
9FBh+p7Slee4yRjqGgkRk5yaXX9A2TG7BCtV69vY8Nft4t7gDfUP/NUTqrANKbzc
DV6aJjfw8YywoMHEvbSZdVEVOBwtd5+dc92sLik4osHxAX0xKCa7V86N4wEavlk/
bi+GUU8hBOxSsInqajERBHlI7+4m6cQIc7YifvrCM3ENwQdMDY7v4Gh0m0MDAOPC
epE1W9ouhTmolWGZmhByAwNN3zz0/kOod941XZyoGl6KuPt2DCw7EEtfbHEWQSw4
xKOEDwAUvzP400hPMJAMy5R+vg7hP338HTgVvO1TMAXbhsJwjlnQiX0T9M5N0b2B
WR9mSBNGh2jcEmaoaCa0lEZGSaaMeHc/2emFLwbvOFNMt0v6SPhuU3m55ioRYnWq
pm7V20PKW/pPi9dzCyvzYUXufwWSFYKlJMjHvxLbwJKCz7RxrnEhrJOmkS0pgMUC
4uQg0BoftW27VUVLci370NbqoENFGDE/P0MOPuNq6pZM+S6zvV4ako+IgHZNcyIf
eJ6f9FOWseOSaPPQ7EBLTdyRY+Duw/yXTdJD07vw4nxP10ktcnnde3OTxYZ1xBm8
DpCVQ/jyrM+33VYJZB8FhgzSwedZDu/z5QpnU9x6wTvQo8UzclprmEaQk5AeoaxN
s0U3QSZQbRTy7+ER6Gw8OF5Md6wTSFhOPOowWw9UjqEAPwVcA5kOFvKawLFsYkrD
DjZ6QqEJRgzGk1h6K8H+4G1LwioRA5ImyWERnZKEauimSuoqkSBjRFpR9jnxyWGs
ZwPZwxDCiO6dy+VvwCnjKCrPTKVBeGjt2WuxpIL/b1mQvfzsX/r1TuIDRkTyXMrd
g6Y0y0x+W+t3MeMUmC9xIdLpt98O4VyPRyMTr3GpSew6nC3CwnCpODQu6GBo94N1
HEYdR29mHtAM5UBM1kMWPBuFRhD00837e2quZjf/S1upFcS8ntbbyxlii+d/vsy1
zhNX1zXe/iv7LvLvN9kjmHgBY2YZFwcldTvSQnD96Xi13kZWDQnZIP772/uPvy1J
5tgV7nGxlttl6DLgWLG0u9gyAybjNn01I4DuiMGmPQWKY41AWFhTDWup12ojgLs0
YTu1X+ofJtL9YjRJlSNvn1oeb9QslsGhVc8Cp8EbjaEhRL2DEujmk4zqxoHWqLUa
9YcuqHil+6Y00dEGwYUvwahNdjE9EndgfSVyqPW88ARtRkH+Ttw706+gW2UTwzPZ
hj28/HRH1o524mmAsPa6V7ctCeUnye07QTsOzypenw/selK3dxbhlT4VSWXSdwjQ
FAFd/A4Saxp2qYuE2E0cexZgavbY4qR/jxrhfu8dVArSyWdIGIyidjtZEOLTXEoK
A0Mr+ZjuuVwbPjnj173n2nlvSsCOvKxdMkMcCmhmVJ8d8MyeCUmun7KaS20N2BdI
qR+i0KBsmdKP1aoUCbN+GCdYEuLbgvu4nbB4Ft/8b12UArKhUZXPvoOdjnmDo1SN
IjoE4+m6ZK0hs4WvWM4kcjFqHEYyldhXCiSMw5stfcf5YsRErNXikPyhGB4nC8t8
fIguwbVdZQgOAEFRbKVBIGqBR7d6h2O6w1QgSvgzoGfToHTIe4BA3e7mdTGMZpnk
9DVScnILN58wYylJ/EC0bTEIpkHaIcOZ5uwsR848bA+3nOO6aK0XR9IZ4QX3KLpG
piT4eONmNBZDoa8nsf8MoxBrIWvS2NaY226dn67kgruDJoLmnslVgcJ5OMIN+ljb
NBlCAbYxrPz8ozZ6b5AQQ36pYtNDu1VmGm9KzAyzxVwWZLjMfW7OEVf54NwmoCvf
g7jN2INKdp7y70akJxsjz/7V+Iv9oghhzz9+JmQqpOqXj/NLSvgTNMwr7SXvn/bF
yLzIFQ9pBnl9hTgkGTrV5bXvco0ug0qLO3UmDBLyoibmhg8+LqQWfw5vkH4h/Vv4
V+zWwJ5Zvk6jyxnF620jz37IKPhZlvdEi+6M1jzFQgPv04i0+1KjcIoBGFiimj26
OafET7CP4mX/duoTmwg6b5k1hPlScaQwI20ki3EacC+0OzwPkViCywvN6PRk07Lx
4eTLDXiMOSuzhgbs0eP8i7Bu3b1epr3Ycl2lf1vJMGRdrd4pabMbOemeBXgUxqbM
I9jdzYlyLsg9PLz95Llto+4g8Nx3YyhahW8OmEczzpsgqLRsn3FIx2sb+iKea0dC
rBAwYYiSd18woWzwvHJ0YCVziq96X6WVbpIfKQESFeeHAHgJWG6rdnaG/lCrRRQR
4uv8omZMDaLe13bnnuJREuPUqTvenuqr7oimvqa9XPLFa9PBR4vzDNEc5hSrYpop
xWOTYpYB/dR00Fqn4lYexhk4WOzi4wgtFrAsrFa4DuHaCaC/97Sv28yAB/jrIqBb
Gdpmta7/JvUzYLaEgvdtSe55Lm5D9F+MHWNOAOyE1Qho072gGU8ERBygM+YuePT+
a+5lltQLzqTvZd3dlgxEExAlZWiap2etuaYgNvQf3kiZcP4JMlCXQoZAWakYzfMQ
1lFyfXLkLy4rEXoI2Zey+grR9SDiNVhQ80G46vUwHVfF7f7Widrw0kIpIt89qlDT
V20IVS9yD0KugKUriwSOjL5UzTkkmv03ab9d/14DagaMJEd3eTWHcDoULoWl0yLB
2xfZh2TsGkkKMcPe/CV3Tm2UuwdyGCFRelKdaIm4caie5qVyesvCKfsgzSKoXOOT
xyH4oACwgEnKFgZpNoHz/CKMQjU2HOG/s2Y9XcFwPVxgHGfKk7jOvMm8DW7UQsfx
bXaEa7QzWycvjdCxVKWbOYdtX1nefvrDVx4VOXPYuJ6bYSrhEgO/R8FhK8utdf1+
rgfm1/+8lKHXzOtORRwTipjna5rl18ei9eQkjL5zrpRSV5OWDlYO3xCW38+mVwLD
mewBVk1qV4qfbjBQn2J096qCXlwcCvjxYqketh8s0u4CSy2JRBH0lSCndZz46zD3
atSg7oIn7qEafLkmOulNFXUeekpuCASe1tU11SyMvUBTkvfSGkthCCcJ7sPpKvSV
TDq1RxQUlOinyF9+7zSRycYihzu3uiIleHL5fqXEtKHRMuQWkV5X1M+5MQcOMnao
oZ0ZPz9xTa1nNmqkNALMQTSvuZdrwIVXInn4qa8E5fQyt6p8aV+5TvwPc2k+pZjl
8YFaaFFwAogo7TdMPNyCp/sVah7jpIuO+3i2E/zq2tZwqi374kM7KQQLBlblEFyE
nYHxi8v2O9wrRWiXY7m2PavTeu4/eNAVCoNT6Y1dAS+ebfVgKfbolD5x+kM0Zffj
r/Mto8HnKGPDndtGQ39WMlv+/D37f8J6HrjIM5TursDYFsEMAndZO14RdLwDQXM8
P3W3vjsh7ZjVSwKZoBZ4Fi8zGGB7g4c+eQJ5/rS00R7cPx6wYSI7niC/L0+Zp6fi
bJpaU1iem9iwwHs7/GufUyeGOPj54m4R1iryqxLtEDkr6sTfeVXgYxoarWMVBwd+
63AXSgGz2m9sV/Rc0qssxH0CIhOxn82mBFDzIaEsYGfzhuiv42tHxMAUFSs1azTh
BLfWcGkqWrEZU2IoZvmiie/ecxb2vFF6I1G5cNb1Y2A4PNHK1L1kpywn4oFLyNpY
mSk/Po6TVHOdGqZ+tNoqdm9sK4kxmrwyl+z3Xfq8DnINh09EQ7Fm4PuZDU4DWaAp
iwFIjfzgv9XwyEnIef7rk0KNpdkmqKBWsCdSdvD204Y1q4TULPU3Mg/d4qrG2jy+
rG4KZ3UDVWaWERZ+iEFkltgfWR+B9lDPthlRIc0VACC5E/PhlHKmKDw20gPTsfhs
ph4IvDL8A+yAxemiikR3M24AOCEKo3CgDHB18JoZxsszOTNdRG6P7mdEaRVMIoH7
h/TAZZM4ehjF9tXLOgsDvwfhTavvx7/dzkqoKxSvsd3F0UkOKkwCQ6VoXqwhCJnT
xNyMXWzuxhaMVHsNDpZoqcaYFfKCcZ1CpSOS73Jwzm07zlzhG4clEZUX3gSSR777
LTF0kyjCJXfkuILE4RV5xi4UUpr2P/eVERNBdhfQzE441qPDG4FMfdsEgEVzavlm
Y5QcN0t/iQP+tBeDqbADrrus8L+utssFkgBtcyYPNgSSMsiXzkGIQRG5vmiJVaUt
yaQbdeJeO/11yZF3KY14qv7x/8u59gX/tC14CgxJovHfM8ScOmPyWWyGQ5M9Poq5
UP9uTYv793UD9HyXjd9eO710V4fDNV6zmUUmi7rIQvK0GlJN5sRSq4+UQAjk9uHr
awYvbhDbHrd9KtR4UtjId333R/sask2fo7owxDQcJr1V50DeJrE4Fdi34w/d8ovx
LgyVoAQBl13Kl0X1RdNsRLNFyHDl8zQDidUwAgEcnYSBwwYsfug1+xoXgaZDRCb2
nZui1gXpkrNhfdlypZwBYP6awb/XU360FZiUQ8HlCrJ/S+RTkJ/dOInmltJcw2CH
VjfATsqXXshyV0v/rTF24pejI91i8B91L+JguzvI7pmRNX9DIoGvrNYrlrlcqlYr
XJTJjo+FfrnP1V+h0gSz4fSiQ1YWkwbxhebm1EUtL6CIpPdW3TOEFHfTJBnz1w1+
uOqBgIvXXNFJZDC2UsDBPe4iml36E+mkDaGTDRKqpcmUA7Zdbwzss2WR4t9tOxab
mMtthXkGUA0F6yEIfQoi+CnU5azrgxcyjWAbMGSnZOziVTyhrHj7SblqUVl3tKPq
hHFCy7d0Iqyf77Fj3tSfxixqYsoV7grGvbGH9L7R9KI4mTb022HpqQ8OluWcmrip
pGfYt+1h9LKYBxLA+XhH+uqwTR4nijX/Bkn4g1s4QDCBD8AVm6Ip0N4cuHXbQTci
6CB0truTfI1inO2HXED+bDGNejJMBFTv4u112Q+uNJpnXe1yfIQ6Z2at6hohP+LM
jLeZFgsI2c++zXFVtSXZ4jILpTkTAcPzaxP+tFCFnp/feX5dLlDNdM3FhIK2uH4D
j+lIgkRz9pN3WAZirpnznS9Gj38zKaC5nQz/LKbSELZ9KmtWPiZBMo7p35UlPfhn
/9amMr23JcLofq6dLYdpZEiN7/uPEyXm1osND7Rg4n0sWocCgYKvzZ+JJNE/4fMC
QnMigp+ivofLpgYhDil3phy7prnE4tsGcpSoMkstYifNyOAhHygVYpkxFgGoH2XB
JjQIztyFFY/ctoeDoraRO8Zek56vE381dGcFuiOdy5utoVI9BurZlb5GvL3MAegi
k3NHrvDIWlkIS2ykGiczCmrFq7bKpILP7zfrayK53HeIpC9HahVu1tQJ4yf+qWs3
ck2mn233+PVBkry+9ifHk5ZxING/Rja7wSAp69ZEXLPOo9UeTzILPFzndu+QHC1t
h2HlOrisfZ1GG3U0MGVUtcqm8XkDQkvbrqnVM0STdjlVOQXK7UnH/Pz+nxywyAnh
LBrW3Wxf1gxcYp4P+xeDoIPn9gTHgT5puhIgAKOUksT482DJiJR6OprpqQBB+i1y
atMlVo2nWm1UZToSf+a088KYGBNSO7kHVrjrL9pnb0SrDbP2OL2TO+9xS6isUAXQ
eONkPmNCZBD8Ta9qsfrbZ853fYRPYKZb5Mgfa1P8HQbI6DHNIAPEiEplBIxnIiYy
G+WDUTez0WVQ5KLzQLfqJ/j9dyesdU0t1krIL/4sziRmQ6sWsLkuYL4iLaLqepm3
yciBDLi2xtMwrPPGMQ1xdFn+6qs7atWVL+UCiXrvNGXiCtua9lcPmNuf0lyHEnak
8okrmz1Qp4V3ZJeeUVv/MXP+viv2mn0OTxnhU1Fsd/hYNJPcWVKVGKM25+JvJJkV
/ppc6ah0mMuj4Ug3kNPjP85TmZvrh8VpL4mIDaSb8EzehVXP6nU7cOO1a05tx8Pi
xn8PtjKwWsxCOG7AbMV2Ir4xSLRI/uMTvpUWkG0N6I4Rx9+NoeZBsXlO2kTp0glu
iPCEomQOWn86oJWmUDbUMqo7zjynydXh2O+hIfMclJpO4Z80/yYRBBV5e8oAeL7Z
/KrUP4pl92V4W2+itNWrJCo6TeTwcy+Gnm9tF0r4CeqehQIn2Vny0vyj0+Z4G3l2
y7873sUKXV3jzr4GuWaczJp7rvG+JDoeEw+iHOMnDoYsmN5TErK9OR2BSxpnpKxK
26cwcP+LYFH1nGB7su8i47jcYtkHpC1mEM7DP6oN/z/wemg2e2SF/gdwcvuMz32F
j26RqUQXpSZ6HwaRTpY1L0MFcYXivJ0Ec22nlVnm4oqonfFjeVH+WVqcrTFK5asX
x/T3OXHk38yKO29pdXBX6bPOPlq98JeLtgF8M1dNxMmlKqcjjE7nwsVIlib1Cwof
vUqsuxsuWdYQDkmSHSv/4jlXsgrCyxmUbchV9qBLU44bfCX1Tq1+og5yzypRR92P
VLfKem0FoStiYW93bvh1qcDMqg6RQiuwdP+2WnRUXFuCk0wVmaPdLjllbDFyuB6f
Gsp/TKUmOW/KKb6mCKR3MFGQ8i1eK7ZM/PIkNSdxXJrAhcGBXitsUTF2HHbyUzzF
SnA4yQkcbz07fcEnUP8oW6drR2ibmpZVxSG5slLb1XCrbz11LcrIV7jLMvplLRlY
NuwFJD86Ho4kkXDKDOTz3aUATrx+HjNkbVdKffYmuMTcsblkzxGM2YesIyrVbsb6
i6rPIUfWjAD0ysv3McXRbCEbnt+I1bRMnTPCATC19HgB3vpNNlaU8nZ1tFowQqQz
k5iWkOR/DTJDV14LmeZlHkSuNgyKYJuIGVDDFMdTbW/4oAp1sUSmFvtQwYQA9GuT
NW4tFZEakbWy3XfQpiQc+K6Vm50olsnjoPy0+QoLBbZnwJCrNnXFmhXAMtn5XmV9
lzshNvxJEk6RLZYWsTdy1pF3/YGhqX84bE2GBCcT5u6OaKtV/rXnhHRglxLvI6pU
OilfazCsXOAnD1DlKBeIS5Yn/IssnS5O62LOfBe7FIailtIj25TUSvV3YjUmzavs
sM7ybPx6w8EVjPzNCJi7dzvDkV/pF+mf8cnUvEuZkP1FyAI9tt44tObP/nBDZrOT
iXjeuZb1ApnP8ic8igi9FMuLPTp0txWrFmDyNUFGJG4H59iAauDgMr+2lC5sOZLh
7dkAvrIY+XzETY4UbCz4nwhEEFzTCdWZxUdo2bgkByabtEtTrKL8jz3s4UzPWN1z
EnzB+EiZfmPyAEkYnPTB1/KxuZr3DcdoQP4YztLrZqnsgVjw/Io6khHWVdqJEXJx
szNslMF7xuZ1peK39XPY45GfIkhfWFpgAjAL+iee1PCY4rqeM9cN3ula/nKPIa5z
dRDR9s3/2zRjlIK/h58pP/vBqn0/w0nN+q1kU2SvyHIRdFa0IN6ExjRgSXR1si/t
zRCHmU7OwxTncYuDCNiYtvjZFDf7PGIQQ96/4L40CQ7sTNvYPQhFj+ZgUvn48WOs
ZYHu1KAR5vLlPhfJI7poxjVYul7kqyob0ZVD1S71V4I776JZGKx+DWebbld2nTFv
ZPe2DNDUrxR6xXLjCRHNJ8EQ2K3D36pMMeQKWanjcfVvOeQ4hY/kRvW8o6L7mPzE
fs8su4Gfjf/icInIZPBYtvG0YgE/7NEsunGZSv3H4mNDVlnYUGU3vcEPOKV+dbiu
yAeRG8lgWwqGpmS4i68EJx1n8c/esB7aqKer1LqnXgTYXvZgPfQrTdFWVlL5VR06
SbYZJkZ5z9ZX0Buklr/k4rYLj57UX3YEj59H8fEYt9Q8ZStEsM8VCH5AsSNNOblt
1vxE1SFFXSGibKYY0SsYQxFy386EGwpXOWZIziJO0wodMvfQdhO2irZUj1v9DxG1
dvRidRvw3KqAQiuz6EsRg4BhMf/eTCjDHYE9FT2DD+tYOhtKlnkzUN1KRbWDFGwR
lP3q5ZYje1OXgqq9uOfRfz4IR32c21Y1Z48wKnYyNQMmeKylwxm41wcyw/yjX47I
ZaeV3nM0aKZoKB3d1StAMxjObuD+GtJCiCTXTM6y3gIuAmCAQ9wAOe8rFcvtZXPy
GZD6BfmlSJykgJnA5eFgcaAueDZgci47JyBitzrQR2pEXk4DYYvlKAkHGA9YCB9Q
Hs5pIQtnSrJeaXYpQv8ddRiFV2PpzwMkIVaaJch8dK7MxpgBe1ojwoVC5DbyVNA5
BjQeD/52855+fJ3lcMkIJXZGNQIlYdPPreoiis63URkc/+Ubh0Hr4hG28oJ5BQ6W
m7AVHOQKXd6Y4ezEMZNjYK0lGno/CItWtse69Gl3EbkykP2tfHLhY8GrdT/mXdTe
Mv3P1j4XlD73Gi07pYNFpY6UxYwW9KvINQXDoyoxTrSmS5qmy2heJoVqRAbddSXs
zFd15UCUbROtBhYSK8UxHub1NpFvTnBQFjVVBASoc0eOfus6ducwLwBe0+YET712
CfMjjCEwnlP7B0PPakenmCd/+LruhHmwZ9FlQrqzFEf95AJaFxZrVrTSbwllJKUJ
XrcLYnQ9gmV9sCfKZ8yscQtKzlTMwNKazjMHNF6yelD1Rs8ynt+yde5xg/B/kp2M
isS8Mk9msqPRtBSJswkENpy2HNn25w5ACmiPgr1CbT7Z5uW225Do4eIqmjNOXe9g
lFVx9ziYxilNH9J2VFEuzso++GYrWeQuIOuB1VuJaexZ64Kiq96NqlX2iWMAIyex
eUnKxHYF60L3u2GWp7o7vFboXGJDNz0Qwnderf5FrFm+LdIclPVEmtpqkggb4wNE
FiA6p5bhIYPtcbtCXKpInFO4yXET872aXx6g10qJBLkxySV2GJZQR/r4j5MJqB7/
lAt/2usGVT8rc0AK1LrE7Ut/dDqkGPwqVIho2/4a3QRkb7DtH0cEkrccX7uerZiY
nM6EkciI6XvCteX3Awb1mJbwWpUN7N4rFYlJhueSiygC/GDkEREHq7hqJQrZu1Cw
kK67msCLs6l6LxIeI9ONofe5l0CIE65LZYG2bIx2h8T/iPMTk+1NqreZNKPbsg+o
xmzR6znBGm1U+sD2YEQlqbctwz/PfpgSBhxZ+s3zTqy8P8D6wOWHJs8O+Kez4HPs
YntQIi357hCNhUquNpV8pFlyq6+bTUPKR0bY8j5T+MyVH12794ozC76LJl/UunjU
Uf6L+ud95H3FtpQJxOvt6vHSiacZIOfYO9qcDkpRNeldwWnmOuJPooc9b+4tj4T4
AMUg31dBV4/Y3MAz8TSO0aJ8r2ulkNSQ7ZZTTE26C1DlXqyT9v/lWWl72Pv52K2I
uqX59t54csmU71oOfrK9Gnnq9YpQ9Jd/RkH8NQ4dFK4mtD/gqAJsmahHA+iPcgiM
vY4U3jZFFuNquL3RECyaHJLN8j18pcs+Y9iZ9b6x7IyERH46C170uCM8WKKkBzT7
ESdXDXN3nqVtQKiXCCRlVnuMyZWt2/qedBGbrik9joLFajOpzv2aGI69ucJd0j9Q
vU7fsj3ckVDx4zqrNh9SAXCLD6OlfjzxZkACFnf8kax9v7ID9QLZkhtNeO5a6BzK
SyGOSZ4GqDWvQx8Kto3WxDZS3yilzZR74EWdx7TMLreflugo+YifvmL/IeS4FBUu
0RtDULNZcLiSW2KGb2hEyxJ0PUQ1JPEc4vdkiU+3WY55SlAn0bgTkkiRtdq80hrI
VXd/eOz6HtC+t8BImaMbYkYT4xOEQVZ23erLWZdKaeKSYkdS4pqEW/32ivBdrHJ4
qSwmQPTd0U+BpAVdwZ2L+cDP8C6Z4Obg+/T8PR1WE7YZKSHCTbZ4+Y7+la76qm0I
katZEViNNlRWUAi3vkNXtEdwLxcxC07CAhPzOT8Dgoq1D89to2elPTnWoz5WlxxY
Xmj4ygfOR/QSvGnxMYlazVqyfXtBflFWFeZYZexK/xrrBh4iw/gpdQKfBZgg1j13
/PEOiKmgZwWnt7Pr1LKc/EIAeTcVdNg7taFP8S0ZKYLJ58K7fq/AR6nAd7ZaaDbU
dFzMNWf2nEdjooJlYWpCOfnonQd1xNLQAxpA/DLj0iNrU1zTLIb1VTiiNnmBRaIw
2KfacpInh0v2eZ0wTbU6PNoUBwR2rLNFwDTy0wv1J5H4tL5Px8MxS+V4MPEI4C2l
XyO5y64sAV+nRg11ECBgsZL4mF/uZKEFZnochPPB+aU2OBj4QfUPjKFZrbOWfDOT
0P43KwCgYgCGaIF1A64R8M3fo7+Qg1iiAO+Asi5ZSm9jkOYDX5+e4gbjhuClqXDi
gxsZkfcRrEU7r0yMnak0IsaTj5iIbuDHc+Rv67TrhXvGoqUKslyLhWq+T5tpzhPc
7LAQOeyxu0ZbTlOK0sihekvYbYQv/mdUj9GAo6TH5Ix8w0f1l+GwmYOGSUkvslLg
xux00Yhf4O8YLGPN/Sa/9vhDd+HRKYQcDpNCWSXbkA0uoLiodtaaT0mhJuEnVxYi
pdC09Jlq5p3vOpygi917MifpOh49XDvEkOjvSZ/rESZpdoru1FobQsvXcz5T5eUQ
06k4VCwNfTSfFrIs8BLKKXPyZS0Cd0kF5MSO85RtwlOxvzt1tPxkEElmI1YasxKo
LQmshSGUnkcFudyuNZxpYvyFsVvM9HVkodXvu5XWd3QBBvW8XtbbALeZ3dUx8gsE
WsRikrmFIaNBfLR1XNKL+B2i0K76tNMssKJRdPwHoTsJ7VbVllvxZ9r52smMUQsF
HfIp1B/Qa7X/B+maeJ7pjndygmvh18KnmyKIcUf2PN2zgJJ077WbAf5GHcW7HDLL
GQQzcM29Sxm6e2yupPrzLa85Mh6c9sFtaYs0kah7wbwzPL2q45JFQxNTlzeDLitw
YqQ1rRPT6S6+RKfwZYOA4ELzMHuojoyG735QIn+dIEBsyPkkaPXLuqZ+wikp8D1l
Q9zH8gaBSXvcavAew+cpyqTf+kM4vgRUmBiYomv9rr6r0S+sFALLxgTtjakU0S+V
9ju7OAaeIi0luvggrTINBPY9UwWmyifYItmfdiXy3LuOcw757tG7U6KfT/1k2cJ+
h1bNCkr4r//Z77C4M5M/4ERmlljPoej//4A4eOB9pPP2M9rvZ4Gd7cGpM0ro+vh5
PRw2EYS2xuNDaNOjj6Cfxb/l12DLTz4EuQlncB67TzXtupSclMwchJtKNPpuYV/1
w4nwlFepMCFod8CtIO4sFB74jpi0mhPg1EXYqxLfjbs6gK1giXli5nQSQUBefaUy
8PsGxNlT1GtY/E6R5MuBHAh1C+4QgAMvCW07WFOwheUCuxIYn5J0Wk+pHzYMaVEY
5DaQpYDiHaeOBfX2l9e5Og2l6G4ByitQNe+uqOUjy2w6ig8RN67zotEo9HRvmNBi
sV0gXptKGUPv8Tmntxfu7j21RDje9seVJRsibcN3QHubXbOcIT6EFdBv4nHGLGEF
OPqkHuKfgrNZ0dhvh0eccgeO8D/P1Cfcsf1QYcVS4+I4cVSCDqUGaClfo2zI40CA
0fqGwn9YKj0xGy4y07l8Ppf/AxVDpYZmT8RjhkgXoSsi1nY3ax1DM7Z46LP+PL9S
7bBlsg9XmfTal+GoTbdKZmJ5qfenn1xEl5rjJijD4E5EQciKMDGGudCFNJaght2Z
4Fb5kO2S4rFcSxZS5P3acJIwpIVE1UcMFP80MUpgUdU6q3zR4R7ZaU6PjFKd+vJp
60eXEo8SEop7GINnefMMdNHcxBcViwFo4mO54HSTyukMAVWI0HESRwpR8xKASfDw
5whCsKju2dQBZ39tzKebN8rGhwDWlWcPUeQtJWXEAkZFKxvJz0+ih3RgFakrJAFZ
PVf3QEaVfmMepTGMh4jy4yhF93NU0QVXcm7TxKIpSVPkRnpZ5418p+ZVyZRvC8H9
89DEuT6zpaJAydBuWbiRl4w80W5ofA+H/2LnBzoOdwapmEGd7jiVUDlodpEpbaAc
NHG//dACaG5Yoy5yMtfHn9c6pWSqfGgoiM28WfNdF6ooRLFGS3NdmM+2XGYMu0IZ
MXlCKLLDHtTxor0Uc6e3000KQs9Nx4raKynvKka8pzn3zZpigyAg/Zb9iJaZoZQ4
ZSN85KTAvlZRLp1qLc1Sscasa8RdjlTBwEGqY4X4IbRM3qQ5qAJhfLdy6vN9uvk4
1Is3UJHZsIOy0E1JpHGc6ou1GweLv/SIlXf1kOiIeX7G+TFnvI4WZKCfpWqss5Uu
XXVSezqmsuo29meaM2dSbad18b9XwSWqL3gP0W2qNNLK1rH7ZenyVi4h9OiJmi9O
IjpGEXmxCwWtajnfO54OvsDkxarGIewv3B0V7EqdPe/qu9OU+P7Xgwk/1pga47hC
r7cGY8f7Mg+/AmvK2qh+u047tPFUeSQ57De7gcXK9AAvRLBpQo3Yr+U072yiIoyw
bNWfu+vV9tcsxQ7oRVGMgRQ2IQzb2yMhf51O/qoMnLK+L0MPOESI0a5BNmkIXX8e
LNTdmxgwqqMAOXQCqpZO3AOe3kMLjeXNsfhKlwwlexEVcq2mQX/+w2vn+DuAgjkq
6lrc+DZV2iUWbBuZTiburlENK4wsu4aCp3TnaFYvwwNtVcZkcdrHBuSqaz2f3dDm
W5rxq2h1lKcnQ8Ghn1Jeb2PiX7oyPe0ma1Kzz3b5mgUgI1oIzZHXNQk+RTGjuaWs
yJCT4SfgtxejeCpdA4JQX0rXI+6xeys54DWrQWsgNGTlvcmiGJHa44QlDHSYqw9u
kF4EtEyhpIhDotPdLWKS0Jr8w7ClgCpFV1RUrTStOkZnGOuZlsWb7UoQ2opJn2i/
LZlB2Q2DagvNcfS+hfi5qeCTa4wNh34toyeReqh79I//USH3q2E7KTN23ancBP4h
IHxl2TF1SRNmpPqPQ7/EJIre+8S6JbiFgvnv52uZgc2ocpOxjYDOkTJodo3/bCRD
DhilJ7DYvc6PCle3QQEzf95lQfpjjXGZtKY6YgrRh+H4JUsIoEHtHbNvdqBTpW1n
WeVuTeiSGCG4WH9+BYRLLcSqy+LgIZbsDKjB1A6XPLHNe217ojTdWobCFYc2JK5l
Wt8xveY/Z+DrKtxotUBYL8AFBAtrjZ/A0HkTX9gjsuMLfv+Bf0rqhycl7Fdkf4wI
ry0ztiX63Kb12SvQkuDf1WXH5ox3BDo5x7V6FFTG4+o8uP2tVRdu7zhs63DC145L
BEH/zRxKXEOJ3LrJD1bExnXqQSLe/BqPzvHES1/cshWsdCW+vXOAEFIFTdhqV54u
+XcdGDKbXXyTwYzDOVuGmK9CQjUzLPBk3mrtUFFcDOrgL0FKHuKka0Wdf9QPYIlt
xFwImzm1ieyPhih5IwQverlhS0/Ry7tdUxJvz+wyCGzeus22w2V5TnDBLNQSeNTy
ABT087g9YKHUc62I3OknIm1pyVBJN/DGAE1oWPXXa0sNcwGMyjwbl72GRIRjsoHs
uYIodo219FOA9pyBxKtxqt8RfFbMrNUqlR9iGxpfqBU9iefs6GgO78f+yTo8xlSu
fKqIQF/rUC5/+KgHd62SrexmXbiAfoqMJWkrc6xL/1JVy9/oX6+dUhV764N8uPLp
16yhN1VbGxR4yBXE3AtyS/co7QkuWe/3ywGnid8rlMhMOvTTe2E3gLB/h7NcVqiN
SBFCA4kwNySZdsgUN+QUQA+7943w6pVpgiNYr9VFIdXJnxyptyw87Ehrcb+U2/Pi
YJXb0nitCAUq8TNmJukeDw8csT3asXqjRo81KXRs3za/8NYwODBoHXz4IxorlRSA
ki7H1dZ2ecq/Ob/UqYFsfGLaB9E4eUT9LAciqojxZHHrLBQWRNNq5ZTJI+jy3ZlB
HFYA/K8CM/Ax4yWynSFbCQq5r3xtPpKgY4kANpHidHr1oB4LukyUm+2Lt93x1Ckx
84QdhuOyBj5kIJd+AhxOinUPtSGp0lJg/SU7ywrNIO1c01skeAQQYj+UuyxBpQTz
sC3TOcDGEA8/LSB6zCom79xbaobU5QCY7UXXxYAGoF5uyew0v1KZ8hymfhBZNo39
i5FeDQdPyGS1JJ/lJ/WctPEFWl4zMVHwVM/nCFtOUXiCL/7ezZy/XOZLKL6Mf9Y0
R84JIUzxveS2+NG0JN17KN4pZs13ZngoyFBZsS2yWzUYwvojnJRZQLe61WMwhwIh
Cumd7Xvp50B2oy6B2brisYHJYGq6YDhZo2XD/VA2DOzCOGJzDkduFWx54HRK1AiZ
354x186xj1VkpQMyjUdnt/Xshxvh8UKxEg9nV207waOzDiXw6qQUaNK/HUwaHMX2
kqsYE4l9PjS/9tvdMhjzk5OG/+XRR1ZB2y+OmZmbUp2Q63PWDG3Zyr9OUFtxyMPT
u+dOIpgVRxbVwKOIdbeJi4QfPz9WNTxFttXp8sWrPiXov+HqxJIgz8rmZAzEeY8r
W9xmp4+hvZ3Xd2xLXq6oFfNCsMtAxWNJOTfMyrMnTRmB40mHGttGhIO3FKYNNgnR
skcWgDETIvdnO9i+BZ47d4IrlW/Linam4ztS9XvepN3qSgJZBblfMFU9m3HweQY+
7494IZ/FtcLF0giSRZHOB9svIu4I/twchJrx+tjw7F7Ee41HMreyhJeaXSGznrWL
VImL43mT1QbSYoshZwspfttqpeDKbHHXYR1T7ArP9OQATysvEUd0V4G5hpW+47H8
JqDYfXC/wBihWGQZ3ACc8ltdtuxmL99ehVJGgiozSgZTa5ci5Vv/4ruXP6E7Fmbh
QpI231Ct4AeKvIy7rRPzYRT8PUq8nR+HFPfOEwYl8E6DI7OBvgKDDyBWMI+T0Q7s
xiflTcivcuqXfv5G3xpc3woq/gO5TB1G23rnIJkVmq0cQjv0K+Uj50jaZog7kSoC
ViWtTqEEJOimA6GoCqraeERPpfoHzktgjsEIAWS6dR1ciooQD5EEjfyou8RAbsPT
CVpQ9uhXaNJ7jOSzF+1CiZMb3rJFnlrJIeMekEpIxZQiK7yt5ui4Zzx00LALFrw7
gxMpmvfrEM5+NKYuTpcWrvWffQeXelHUt9XS/tWgpPzj2tg2fgCJaisY2qGfSmzi
yzHXVwmgExF7JV/LxzEq7Ja1ALq6sMqWEKTr5fjPw746N1G/B3kmk+Lk+0sp97XV
9aZX2W+6MIWrHjvuRzHn57ac/JL+G7c9pvrzRm31bR3nC7HTtgz8ChravsqbT8nT
ls5A7BjJKuYlEwQhhexDyfRLyduy/h3Uk9+AS7cySavRXxiXjKDdBUWnfL23BOsM
clWrOrLzxv+KpQvLcMj+4amlZ5k64mKW/T8XomVyCaX2YgmCfgWt5+X92HfZT1Ye
+13fT5oCWmwL4QNDjADtY/rptfSNzV0eFuYueCTfe5xqWaOKGmWR6eA9qNjwa+Hi
vjPHdpoBpl+vQ6UBsXok+GBlNIefQjNZvzdUSFOv4D0J7dZH02pwOGlT4AEUZWef
wSTnjafPGwkgcfTHw3ZV/9vr2v2g7VyyOy3l73lzhNlmEg0fnZnAAoi86c460hf7
Z741wdszaWLGycJOgeTnMXAUjYeqsXCoOOOSaxhmBwaMTQFuP6eYpPKkY2dixe/L
SytEYFM/O0mlfcMIPchg7lop4sLgoKHXFk4A2zgNktIAKdJNGZaCkvHjBjqCWL41
Mbt8vEH24Kc7FH6IwhLlaY5jto9cvDXIkrOp9uX+iVTV6lBpstL+TTAGewFkswRN
tbjtTPMc67xbxp9vd/9q8EH26f9vzgJ6XY3oaKaW5Yur0pUWNCl81JXUZttD5LNP
TYgZvdVqdwmX42kpSarBaEwrij7gBsw0qE8rKLCsHsUovVLEtT4O3ozUT3ynCCCY
PldOrkiVFmtRiGnkqmh5OO4Q0qmIxyX4DhxLAGX+dJ3QUFV7Z0EMdSwHM4MtH9B6
BiZFmqulrhN3knu4waXJNQkAVwmqbsqhhtbyuDF/uVWQUWIlRTmlHbJ2XfDY+1LK
wrmAux9NRxpRRgQH54hX5Kb1cG16z8Ws3NGDnpvVg4SJQW0Y84aUzHsUFkS/9R3G
ZhVr7I8baRB7FCsLu90Y9Y5uFFhlBGdak36+efvO+juJjs+D6QhFSaDFaVdKmfCI
RjmcxaPiUV+XJuRnNlP1ZG7EjJkLVeVVQwc7UJLuOnktwbRcm3FbFMf3qJOqgB6H
h8yIamZvgIO0+sEaDACyjkC2iplBRJ5XD45maGqD6t8tuT1l17yv6eMcqzCyyj8T
4ILTawXpg2vQ3zCtazEmmfUgTBchqgGUGkdBJ3dXxGPL08ewfkzWT60AU7qdNWht
ZPp01DB4YQrJS7fIHRPPBypTJ7RUhoNQPogzFqSUIgnCA72uhTnU3J1JP+/QenxD
H/FvfdQd/9qPQFvIxH7LS+3iuif+sIXwQL31eWqTlhjye6vSrxFT8ks+JAxL7Tkc
qOX+KAnmt6Q5RfyuIB32uTEq+ERosff8bIkyrUw5buWBr4Dry781ceZ0beBA1+e6
MxF7oX3WBzwzcPGR5BfmSBoNOaY4YEaousUCFLrZJMfopdvcOIMCMxpEuAiEr0e9
XR8ViBzFM7pWGS6vB432IPMDKnwsozAcUfSsRhppREj2yktrquD+xsSkICcfnCyB
aOKmxQg9C1TM4SfPSEDz7feHqyla2oUdbp5t3ebFjh3Sx/iChaHnyopH9JQA74k+
nD4ezmJCXIuKS2pPGtPfC1r4t9AebFjGxWEZxT1QFwjX/+eFJY8QS1zArVu3fkA9
cPhFENOEDQMqsoofjHvBZLMaYgsIkrGCcpBku1NOBuCoK91Bny8mRrcLIrNS1A8e
D2ym2O+0yv8r5/7Zu0YuBkOV8UB5lTosHtcFwmWCTUKzj+mKiNWfWOJB7lAPLDz3
0Lm4KpmoE16mITYJtEUtIv4UcjACpeyd5cvWgNgl0QQ9i5mbX3EhG0YVNpXBBZGT
8e/yol1BVKo3XeGfjcVXyT/33hGZBaCYr1/Sov6N/8nWJgzypRS8+sCrdmGkWZBq
dPW7Nj6MZCtlPisPfCUAVx0kgMHHpG9086tQEk/ZVyEKU0YXrq4rf3j2J0woqX11
p3AGtDhZWBoedjGwYbv4NEJaDuaTn/o1R/8dr5pfza3eXmiTNT1v22MEyqEXeqZF
H2z9Ui/qaarvUNKwkBtAuelEDMKSS+W/tH3SOZZpIgw50eduqPBLznRGL62QPhI/
0rsillKm6BK/cnISrhA6St56M/u+6qNHdR4gbHsYj3HR3+fod5PUVT4KLAjwejLU
AqfCDEbH23i5Uz2WznatVp0qc4MyZmRr2XOqdM2Yo3I1JOZroEsf9P43kpKiOzbL
fDpCWA9lNpmzOviOohTjS9PGqAVhYrlUTy/LhM6AQ6RLZnNxUWw1rfNj9n87oVvF
W44PngmdT7FWKPfcWLyAN0Ib5POTn9h3TD9srpHX0q803/etSrdoy9ccCVnhVm8M
5Qc+YXo2ur/VOUk/LXh6SfKIfg1XtYchssx4TRVDNE1YQQ+ngeL6SkBDG7ae51Os
StlAKm4X6mVWNfU69CU+xme8dqL953CEzQ6FhH6i7WtWBGkWdI5gHqH3O4LQ1JWm
G3nIdXGJHEH5TW053WvL0kGcpKLcUwd5icCSJlMkNAmHtrN7ZQwC6bG2lrmH+zA3
V5f24hgDX8WR81aKIyG5j8ayW4VvokSW6KnQIxvPhq6WEumYlrFuvSz3yAxeq8V5
tONrkfeLuS+nzBcMsxikgSzqZ3TAWJDQLcrR2acQGOz7+ec7YRlvYaw+jjRo6Tpc
OT8dUz+hpZUr+N34bzayYGI89Nlc5JYEZ3s3bSV3LG9A8hP+CWiu9b8lsnNLJ58C
Jy/DJRJGYqd34T9VfkvWTv2ggAuHpJVk+K/DOBSoBH9Fvcmi3SIulet+swpHE0YD
UFCky/gcnRhcIKEax67JZ+RT94s0/1tSnazjoOq5hRJdJn7xNrVWzFFC14UWYx4h
K3MhITkS+QjDzDOwNoC3jTrhfGkQ46vozzoG9UzFuRYbmqTrxZV5X1jYh9ObjXbD
8TJinfPYkQmDTnEF977iDS/5aNZSb8pnNwgjZNVeN+/VEqEx39GWE9n8Fm1yii4b
+YH9LdUmB7oM9fSENAVqA0PxaQMw6OzR56MYED9LprDP1Fv/QzXmNa/GYe7xfuEk
qW+MZ2k4OlJ+mLnuUIpvK33+4Mp/7K96i6SYhS9O0V2cAxfPvDVAdZ7kcxKGhEJG
sESCrCTsVlGMP6Vwx0SU9X/VbTqhzyfnbVn3nm7NgGt1xUZDkOC7Jua17+uceWZk
T2Rxn+UtwMdET5cVr8nWJXLZC5YbWV9EYpZMF13qX/bFbOgkpTHhz0xPcXrRV6Un
AF7SVnACWkulyysQEloOXsHe2smUuceOQbEChXNiyoBBFMrDwMoewIOpHbTFhdBW
F9bEvSRRHbUrDkQ+p2zEhiVwick9JnkkWzFpNO6PYr5o1rqMVdUXmUbxY+qWYKno
hsdQWfzzYmd5/nYBI9VNbJPxHXSM7rB7VR68+FsEakbkX9HfmglKZH/7jY9F3y8y
00OIu/4zlnT+P7sdVWkt2xciT6EUKKCxE/7NVdE85iT54LqkWuLL2ECfq6FSVk5B
2nCM1jnD9YIfjlTVs9HYtkOsa0UgqMYZuIo7/c32c8e0KNdMDBjEUOrz75O4ULlO
VixKgRCfhB0aMlkwvUQmUOh3QCccTDzTzEr5jpXKO2fviCl+m4CZ0zmel+CuzjAQ
Z+B2X1CBZkJqYzRTIlvo6W0Tz5RN6h15UwqupetctuIxQjPvPQhCULe8W2ix3HIf
aAN44ONLNLCYO4IP1riW9yio+yLS3JoyjoxFYAar8O9m9+EcKdRcILvxIry2xdu0
id6hb5Ydb81qtDq4C0Pl68P9yoqxEjbl1Q52v5yDyUs+iGy8dY9/UhUgDRFj+PzC
bdYTQt1OtEgrjbAiIWTcAPY5UAOXstnTy5wYXIR2XB0kaJWe8XPzes5r3/ql94SV
CRLnLXtr2q0GxLv55rVfN7ZiyRx6U/pKaw9Pd5R6UWAAqd9jqaXpO/x5J5pWsG5Y
qaV/R5pcNHcw+2v3PbKI9bNKINJvYf3UdFKfh1eat/FlZCKmqMimvX9Ibz4yVDSu
2AaQ65gmpzYbT975L8UzCrYG46SH6LD8eAB8i9esehMg5dVb2/UdT0ZUQ3BHoA3w
XNL3L/US0xQbdAxCv9fk1C0xpSMDWxotRwiWnyo9U2+636CqlkMywxcedEDG5Q6H
injjvKbaeKMG3Fs6O8BVgLDqRT2xZw70lsUoYwlmfqibvrK30NpIU3kCGb8pO2mu
Kwzdep6KovoRCqPzzOpBWD3ssvos14/AE/6NIQUngCcGsekth5E62duP/DDp88sl
Top9Y2jPhHnacJtF6nwg5eC/2E7B/usm5JYT4JNq6K0ZzOWwLomGhtQdAz560/I0
VSZySoPrNdoKN0qa/Oj77wKlF2luruJcllX0NeRabFtpqAYIzwAp/jzRjbhltzSG
uEjVX0LR8TynESvW6Ln46afTjRew5Q3o9y/kSDiMWYZYI6ayRfPBp9djtxt/5uDs
kmo/D9Sn7s2vqdtjSJAiIJuGC8I5TFF23yT4I1f7fsJqRX9KI6O1LLLNICo+y0Xu
nTIWbqAAxqTy9yFdHbODI5W2R1vGCqfTh3c04VTWgdHKz4ro2Tr1TdpHy7eh34iM
tYXuRzSC+5xbhvUdmykaMgQ34V3xQZu3eFGho6m9qU1MMZHDL6knjXBwUZqXc4W7
vt/+mBEId2MkukwwaZdhn1t6yMXao7f1GP2zKeIJzgrvj49A+2JwoNpZ2Fc+KZun
cBfpGBySjJe/C37sy8F2NCGHOE/fbzO4dMUQt4GByAvbfrXbHZ9AnbQfxlz18+/Z
a3ziy8g8OyYT8C7gNnfgqQOKVMptriSjhUVFvHB68we5vMHmok/u0mux6AZ6lM2b
+L6EV+nOauMb7GkPXWHkmvf7+J2VgN1b+Oz4n5lZ+2XIncq+L2MsKN1tIjlAA3a9
YncfLmr+u5yHoUJa/0r1WQid3qhbmtSkRpx+2YI2Ep7phSEx73b6cfOJi4UzkhVV
Dd/CqdmSs7yFvS4V2JC8s1NK23EVbF2a84kbz36Ab/X7U6zI3NQTNTw3BKnGLAUH
y7xKau4vYfLOwGhNHZS6GxJzX/jAZ0qMgJHoRRqN/BdEdlThY9PpM6icUj9DiARH
rZYwh64xkacKvFN86THQ+LPIjDraQoIKBq1Osly35pwzR8f/TmLJEINQSg/32kak
x8gDM343gosQ/NK8cFQ3Zw5HyMmbgrzdyOM7hyeiD5OsqvxIAZFK0esuR0ZxrjOY
hRWSrghdhlAiHW0N6NBfuKIkmCiMGdduPo4IdBpQZeXBo944SCi66UDGFDqPlmeW
b8zRIMCayVtY8G/h5axbPKmJuZXyuw/k1aCQJLq8XrKqWSi/ywcd8jDFwxHs5Mt+
cDACj7FJJhP1sFXMVBxwQH4gG2b5cV6RhPCNJ/cWHUAm4eIRDwh/Z6ARYfQeqGtx
80epXNe/BWM98SHKXgBKlygFMfbTK5uj2Cf0OMinZ47FTxPLZsnovXEIgiuh2X+z
O8tO+TbRN6Um20fRTvrlCeiQrXjopYVpXV1xlODvY3dqSWZ8GIe7VY56w+c3gDfD
TP+XpFN1fDzH/UjGpbYyR1UY/A0hASiWaXY431FoM/D1ePxGLkpjEUwj2wXgrOOo
/qSO8Xkilg+526NQvy69AjFgrFi3MGMvehZtTw0zNQpJJfmdBT5TlT6CGh9gzdf4
92gIcdKR5qdStacw5U98ambq++FKfGjN0dPxdMfkqi6Oxk0hgG3bRDFkvABOIfLC
vHPfvCAZA6LJCpiorZhfBNEBNmzGv3Y/8bxSkpVsYX2HtAtO4RLcH/Cnm0E1p95C
1KCxtPj4gh52g3vumtmBmUXnwdKL16wePC80TiF4buawpUX+z2NB2OFOmHUvfzq+
rWBDh44Tzt24pY7cLXqcNKhfniK4VUwoW01cHJ1trj71+EMBbWetEDGdzMmfb6jA
wbvyjDhj+4PbkrSo+lFI4FT97L3UtzgHJniQ8juohtcAf5lUtc56TS9WYEPowGG4
8gMx5dOGfGS2pY/+c7kq22QAZ/NkcHNtXm+01VB3TxGZO5HADbwBpT+Rlf7dnJAL
MW/+JTR31n0D3qYKmYVoEH4R8nWaCFh4eWiLsZPKomNYfmvhvZcPlXhXR9EjLbsf
bFNtc7IudQXIAI62EhhZEr9dcXc1jTeQ9qOcXJF9ITkA9ViDKG1GuBTnpOr9Fst/
KjWvjjyzy01seo7U0t25Cw==
`protect END_PROTECTED
