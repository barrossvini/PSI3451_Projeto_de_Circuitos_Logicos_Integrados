`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yihrs9GjDsjPNeqJ75Jdx9Y9U/QWjifSDOEBe2UM2lzoyYfWJhxpZ7OQtMZPQj12
wqNvwVt2/wLxdPTpu5SBimmrkH+60fer2PZgvfBWD+y3qgsMWpEyakz8m8iAOIWT
DUsYJvGmgTi5xo8TAvxdkMP/JbJ7tlkmWusauoRNx4lgtcXI1xlTE86LTs+FrYxm
U6iQKGuHA/9WI4GkhP+yFrdJEDuNFHDu8m/XvMqGE86FNYdzj2aYrEEytM/KP4ss
XQzgyIfCnAOE1mT5GVwt5d8b33kmCfvrcbGWVXpTyP+exfpaxEVRw0zrmeiV3zUD
lVsWwSKhRZE51b4D6oKU4YqyPUJNGhFXG1nHrpXtpw5URpvRMzXwzSidK9FakPCV
hjh+yz7FB1rfwaypRZUbYwOtmSvYXudl4z6cbXFt0vB+WQS2MFv2/DjwgTQyaHsS
LQ4X7IOv7dJrC3ufPNe21ryCyxDJSVOvWLj2nD+vOmeXWZcaDuHsJlAXvC8xJ/yM
aJoCuhyg8Q3d+6vkWxSMXtjnXfnZDTKsqKWqzzGtjh1Y945RAKsgES2zc5VJsu82
iEcOMwLQWGUczAZi9wrvggbTgT/sV/NR9LwriUn3sauOk+Gn+5rGW4VvZ9wN1LvW
uPMNyH1hX8Bf8015KSPmS07J+0WcGEBhaI16krii8ogTCSlXRUKaCN7Q2pDMAvHC
QSgKN3TTJLzrQAYFeZBkwX8GBXQQN+55z78+1z8dK/6hSEMgDKLTnhBIP3IVKmyA
cEGMVJ5cGrXDGfezGf1Wi2giJjsr/bubp6EK/1cEDTN7RV9v7VknfItaNrbNzZIi
i6PAlI1NSHVv5rU8kzTp9zc/JAGGNHaaxdRnul/EL1R/B48WKi+B4GHNxMakC5cr
WWWJP3VSdJvaCIRS4DgVFWs/88O4+bQnyD9aUmwI29SeBOKFg2Dx4umJcPxPnYBK
YVXDO3m29Ykr+8EjUeRn/Rlnn43cbvDh8wGihQQUbGjAvrEzgXPpo5WFf3A2XOPG
CDLiIHXGqNNzwXIiKWxfyL8C5QZCZHM6OQZzhplDKNOsm/2Q+B3mXGhxEV+M4fUF
h/nhFntuuLwYvCXHVKEX8A==
`protect END_PROTECTED
