`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+MTLLF6clB2pmG7VmR/GO8lCuvErEl3jiMgpspArTTZ7OWIEHlBDd40FyiP/zEY
kiWKfAX/ezrUMF5H8l0uW0HtwAhQNemNPQpi63SlnhYeCvYbgx08bQqWI11wL7PM
gp6N2COXLZONORRUr/VQm9ySFZqfdd3HeDlVDDof+y5iDfKHMsMFJYs6jJ5l0w2Z
n4TOPD6+jrxU+mTPH50aueKykTpNUeYbVdDPmktMnQFT3/mtFw72IZOL/IGHoHLG
ocscN2diOzGtOkNwjjw3HmYTqgRCE7sIEoZQijFPJlAXlLfsv8aGmVyGT3WND7xt
PFr5wPq6wBgdQZwH4qg4AeDlRZkhieRtpvdyFD1i8RZ8wv5+rzaBVszGtGF8xjLJ
QRT7vIb2XfcfGJJ2Cf6GV9e0nAM9sheaq7BgVsyZOQ8rlWUjD60Lrh7ax9rMQcgt
VzoZtPPNcncZnvrc5wcERt0yHIUb3eyknf2Fzxc6Dc1d36IoQFcvfVG6I2BA8U/y
ZH+zdpA8FLdZPKpru7JQe8vocY2Gf6mqcgwotQhBIZ3WSCy5jrULCEu98LYLLQqV
eb3ahrUR3huvF8r5QxXSMUdiAJHyni9aZwQ77zzhDkTzwV7VO7Q8/uuGIpVH99Xz
Cpl/t49COo7/RIvqeG1mYKtFl7qpeanKOcqhnl4tiay5Qd3PQCyrxV0FERA9mhVM
`protect END_PROTECTED
