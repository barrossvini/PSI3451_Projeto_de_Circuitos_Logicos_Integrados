`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WU8DR/mI2+Jiz3j/H8x9dtBwWS1ju7tObDIZifH4AwAHZ/WDO8Foh4AknPRyKPiW
0BnbgH8U5CHRH5zYqTM5AQUTmiBZaY5sEtAvB3XQ+ipibgq87/PIf0El5es2xLnZ
ATcM5SZwsmraht2izA5761ML3xrIfLAyZwKVAfEedFNVNPq0YmU+AZM0KuFx73u8
qs+PLk0bbqgMKhBcS8Va+EymNGKluXiYCsYQvnt2vqkqnbLJphfA0iGEK2XFC3ae
Q1xp2aKX/QdAdmrK44lY8wp1ZWaVmvRLXZEBk5ObFBgbiRcrszXv2HOFg+liyiPD
K+KdsCX6sf1E34L3De45zhtv//vISoFnFoOlYOAVGrowUsEfUk+2O3KjIE81Vf6W
b3+9xgDw8jz0InInu/qX74ymMdrJUtpimiESAEhUCK5Ds+t8b3dnWXhKJ/RGFehT
dDnKfRd60KtHBiQAPOiG1gZVWKMuhiPqalNCne56Q69Kd3+GRMal0ysJjT7QDNPa
m76YYTJnNMwDllOWX42P0X1DW4iJrxnQ24eTB86Ak1fxxaatzy6JmPUZ/sxETh/r
KEsV3b8cIysP3FRWxB+WsyYUyW9Lo1NpUWkK4o0OsVbsj+Yyh0mxjUQOpsBPKOMt
1SRF/naySwCSv43nc9C0hccz9r+ewHnCPkACfd9cjmSWZoyQyT4ClWJXTkKyGLED
Rh7cTCZwGlVSYVrbiTsYoUs9n4sIJpgDGcx81lo8Wtlf1wzUf20/z5psOK+BJRoT
fbuCmoBkzslXVn2QkrFworB9GR869u2mevbpPIpGNh6T8dq/LIh7rhWn1TmvhixR
sneOD69eNaXcPsyYpurCbWmoAlEUfMkzBUTy4hg8z58i0iEtPUKzLyAb7lZ4Y3/Z
SsDK94FMOmsbyNv9ho+IhS/kPTtYyD1+viueQfOzE9E7lFnP7aa/Ymo7yc4GptTd
waRhA3JDp5LrWeW2HRJIf0MBMhZQNI+YG4ecP4BnkjVKiJInCyOS4Ren2zQPLCry
UqqvmiLgpF6/PsGZ9spgXPKMe0rHnaWlgKZnBMcfs2ur2UFatWVOFsOBLbnBQiRx
CHLsNTBI2NY/5LTSSlOrbYFTQY3Vg+nfFotQ9SMwVKNLeDI/q1FzHw9uwGeweTpW
HDTSfSMcBvHVM+b70WzXZGC0ZxSnknymsFN1hFSR3kfcSBrC+cop9BVV8/XLfYnN
i/yQ48I/PgfyuVbmL+IQ7J36D7g7h00D2u+HNAzzXML+ERUWo8UaNh1SolNoo8mT
yoRJuziP3dp3mDcIEhrG27ex2naIrLWI0XNpAqH/5WSw6hMA8LiyznuQRusQddXg
uUOOt5a9B6q5NnypseTHmgzjuj9Q723M89Us28nOctcsGTOttWfzf0wdrnSb5p1M
3PRAjOoOMKvmz29TqxIBLGDF+ARi/JJnOuXLrkEGESFUiXb1mHrZMMUOFedQuVZT
8Bb+vWoZu+B7bmBRpg3Ea/gvbqxBuydXiYm/PaojFhtQzjBG+1+a4DNfsK2k86RW
A8gYTukmatPeNsLG4LaTPgcG7+pv+sIy4RB+K2SXORFh/hCYayA/vgt3x/4aQ9sM
GWsN90lRs4vaBGGrS1n5Bt8Usvq1s5KrseULKMF6wNdpdRvteAxjMVHbx6sNtUs2
aYvOua581kvgDAXSt7d6YA5zb5Mg5eyin+bnEXdn0HvwWtyG9hUv5TPCkwWKg+4h
DZzSUJh3pvKVuYg7FwKrpFAfaTTTQWJ31/vXgYrI/g4dk+jl1kOeG4HybD9jOyYz
hD4JOPYhYzNWeEtIDKQIvSa7scWQGMDlD/sYS0SvWVGX3KT9KpQDIOCV7N1/V9ZL
II8jDhp2OOyd0416QJ3xtlBMfHp2zUluNxSNPME1XPFonZhrx8X7tD4RDJRXTPiT
43OeoZxknw0LgdxqIiVsC48bYBtAuJiLYtiiPypeekZPqrGdN2uoWwo5wMtbz8HZ
2S8FTxj2WYiJdHujR6hJXwRKgV586utt6t3RE14mP9LcoPtWNMFKJNb5QdQ7nO77
yNA3qnzZ66mutgi1712b+1/3dcECYNq+1rc4glmjMw40LlPx1+mRpkMjla/9Rg9M
Sl7Zs0x/v1Th5uLFESuT7mQG7zQqUgn3gwerhpzOQm9f09uO9EzKe/7TnOsn/Y6q
fnpXb3kv/Rggy8fjrrWnaqomZXkNbmPI6O0Q0evcexHiDy78sMnOdodl6fQSGk44
1HiaMlxOnEGGOGDsrZKEVnkqwc2QoCpREAVZSmEg6hNpw3kYSe/Flc73bPoYNHP9
ZB/08m6Hj0x3T2NgNN1CBhJPzy2DXT/sHTKPC/q7yshl2fFFY30gNP6YWBwoB6TS
pvVNJ/kKQHCF+bAtL077eWcFXl7PeGMzatgWIXs79V6INjsSI+GZ72nNCJo2FnyG
d1QcdmBwbSL0c30BPJX6b/K5clznheQYUtzZVCo8ZQMFE2E1Mc9JJ9vXoO/GGp8L
ffcAg4vSm3ZeyFSYIpKtOq/EEQuc8lBQoPmbj2HaUqfec3h4F/dIw1qb3vU5ajxn
hr49B9B9X5AzuoAi75rcJvUPMnMs1lGbSCt0dxhlRuVqc/6bXzuCgtY8xlISQ8Aw
7OH6zUHKD/pfZfo/tySb7HqwysRp+3/9RbH4xXnsC+FsF47XVGR0ZDS9BYEJ1Q7r
CcRVJ0SUdN3+eOyyInzZAUqfl4WxV7o2XmHJBoJFM8ewcmPsX3EI/2xAH7YQUn9h
5E+fTvMpq7epYpZpyAJK7P99AiMaCfaNWI6bx3jxj/N3y6yuHuLZJ46DjO4Oc/62
tlVb7RhK5zP+yNa+HbXn9swSozM0tUIYpE0ZYfDM8QsNZS3XApuBFCM3x4WG76dr
fqIIJ6R0ndLFmK4uhqkbDwraB3Zc2PYPW3j7gxoVLL0Y+wu0RX1yIFLPkzjbFHUb
h+ftcQpcc0Hfeg8BFunb57a2U94AisRifm+iQB/GGYe+sqDlwe9ur0NLVc4gEoUm
jDOCYX4uPOpJh5JO2JUO4OfKMlTGnq8dDYD8v9k5+J/aY5DoUdWWX6TzxbtcAR2j
Xf5ysB0KB6pBwC6L1yDLXCIeJl8mUgUcYepXohRCTcEBbu1Xymce7KsEGzwaFc5y
FlSi2BoMYoPy9qv9jbPR0LUK657sbWkVBtRwrUFgWkm/A5Wz/YngzNIKy9ogYELb
0vfR6GkUJdj7RixPIhvaypPh+RZydpxMQu9dsOA9L5rbphdaL3tCSw8cXe7c7MB1
nPHlmzLlnnaWIbvsscS52XBcV19ah05Wfpo8pMdZaz5fprYi9+teVhOpbjllmGsR
EkQOhCthTmYP0LuqYHH0yqezLyca2LYHITf1K6jOyKacjfyMQsxiyGdQbk4hgQrh
oYE+LHHUBrxKCShN6B4tX8cZbwMTW7B82fAMhibMHSLiqrDjVEce1Xhhd9SybUbl
XtY6L2J00Qvc9pwOoLU+qbArkZRIbo4xbkMIZwMo2Zszq3/UPbOftc/GMSxywgiO
lcsjWZM55lrHt1mDIh6BtzwnMUvo6e33i7fHcZKSjdnTZYNbDiTDqAn/FGcvqABq
yEE4sGlR2g+6mqzP7AkJWrRMiLOryWtN5wvBj5Xm1cwxPFa7/7Is8kTWxqacewuZ
2zOxUCG2SM4NwQfyuOrcEUJWU4c3Hyk3gR1m6Sey3imXSHKVmmQ1D4yaagmKptA5
HxnAF8uaiJHyLmpBq5udNYk7PzsjbIlO4MN9Co2r9u1wu5LegnOCTuZNCT5fmTgZ
w8yh/dO83hXutT4ZYsqD+DTa8QmiwBYN+2YwJi3ObNBBBH78xk2OVVJ03B2x2gen
u35pqlLFtlmfodugnnbeVEsP2Uv4Rtwe2tRqBwzOl9+2KdSEX5d7WTIhdGyfBjm2
kkLHF6yo7FFugbErCBHmgKVBTaEaZhIs4Xy0DJ8OzDbfdT9xvqT3BNHLO4BSkHON
YW1VFiUJVSSLM6X1LqeS6S5q/8SQCbMFO4PHUuydXcbmBVYLH9Hnh+AkrLw0AMJs
PBG3N/BfF1C0lXgotD7PAkWYdoyT1BnbW5WfhLH22TVWMudaZd/i0JSzoWiWj+Bo
Wk7ZJxf2rpUdx1SNcYtFey0XvIH0WwVBTQRTOqFU4hOC/COuCC5YFQuVI7SecDpW
WjrfrYYD++NptVhUD471Sjv2E2wm1l7wljITq9flt2+d2D7KwG+8z/hlM6D+9bR0
ufGIQKThAEiey+5l8+MSGeV6+xj4t6L53ktPbBkClGwe6oGiM4uZ12MSYGKhDWhA
r987XM/SO46fPUB9hmj8ICyl7fAnM6hG94XpXQNAv6npxCbMbWfV79Xpnv1vYhkw
xVDAxgk5v6NG/Sgzr9G2ElT9kHMS21wnrdwUyFfjL8RWVLVRN6YKOPiemqcujMFa
E6cmwswz4EsBsrht22mlRJ8aMRl2THmMa9IQHMB0BF4XERCdVa3sHzaSlLXKMOOQ
fT70Umo9jZUSsTUtJll5E3eYwpoPlXy+CektjdQm/nA4n17sgtmQbA5zYQVKFvA8
g1HH/vpQaju4pNQTCoB3LgMOR/bqacq7+gHD1T7+nJ+gAZliLbM4ztpka4wmcvQ1
825d1URuTufeQ+3azrGY6HOl4jbGPuvByNnMBJa6q3k+0w5XlOFhighh96wJSLvc
OX2LNNsa/Vu62+PocpnIw5TMvYmE6fExZW52bWdmKrTznNUYR3n3WoTnplVjGfyJ
2xhRyb/MluHWd6T0744LqeSHMwFk5YBZhBgedaU22aeH5mHBYAb4GZ0M8dWoufNW
0YicTPYUw8mbewWGK2A8hb3dubNXVUU5sin5CdQ+3WfDPToOCOVf0YVrcDzmaVqK
BhBG37DdYRjmiEcOP9XiHO0DzVFXqKjDtMWUy6+bxzHRLEPcjmIsSN+lrbzmltJB
sHjoTu41PXhfOe2tNu606RWBAjJMcKbahZI72KjQ8WPix5PYLj9G4Pun3K/qnYjF
Yejg4qlgLDW5QSzJuRzkt2awFJzZFemlFdoVtFO91PhhhZD3ESnhU4UFt55fSosi
Z3pVIVFZNSRuJPiB/iscuHHLqq2D2AjVD/BHzsIngOkLLc5kGWgdH1VI8QoYhGCM
BeAyuGd2yjxSxU/npX/nN1x8+sgevJ3BCQP0XQ/SkkBxiu8Qz2WVHZarsT73gXqS
+Ij42wbv+H6fZAUBkaBpPLyKVu5xfrR3rRCLU6/tvK6RS9V2zqiJRnNK6+UwdTLz
5eameIL8UVQYpk538+02jrSEHcoZefQjvaeramFSbQ5sVE9rAlmBYTzr+JeQkQOL
VC0aiWWVZeWgM5Qj4IVETsBs9yvATzPrKTiBExuVFjNer4EWovWvHff8AkCxQcCF
8mYw9n1FD02qMDMjwlTuN8efAA8xAJGPeYwRpUmJnRpmvoybiA/pofq+K9Ow7W1+
o/0UhhDx3Gnm5BSTmRrsDBqmS1XHwPOvKyp3fq12dZ2/ZQdDo1TVHrB52bOdNPxB
CIeYMx1tGV29ZGgRqsBYi5MYg9wwp3yQRG9JRYdyttKWCebhtJXbeBmI2Nl0fjty
WabZcidoTbfR4Ida54E1UsZKzx6F6udXY0q6/scR7uYw8ql/uvLbfGsBNQbs7iW5
sbHp7dM3tvZbkAXkAYCH9meSApers7+MzK5849cZ9UDJprMAuGfPXvn9d9gtoEJI
2ZABL7sYwbF/8Hq5fraM0Q7jx71j752IEcWBuiU3B4XT94aMivIvT9wmHWbJszRW
GXOG/hPsuTUiU1PUy7tlAUW5RfJtxlTXifozNjV+QxAFgDwqaYxzOYx6Jp9ideQB
MjjdvtBzd3lf5kA8FCYu8gPujvquEjjWSYyhuh6t7RNv6oml3emdx4WIGJ5Sbszu
fBDG8chk2tw8H5PNIZvD/9JCPX7O843Qob7rBWyuBADiyBoaRE6XM6dv/nRMWyhh
Ay2hPoqLRso2ZS3kIPL/5HsAs0pIUNXp2EAGXnSWiCU5WlOyuhpvCq7YUG99VxFF
2Rp0qkzURgsVGbtmNqEsGSrXkqR+2BV1bXeY0rzl9DQitXkC7WHCvXjtMik7UNA+
NFaPGAEjfpXYB0XAsyL+YNBkMm9fnLxMu6nX3MB/RLBd7jRXD9XglR5+Wl4ijmnu
gl0dTno/XvkC5W7dfpR5zY7zbx8BSuiVl1Yxa1BHK89uCb1NCSXeHitOzZ4yTNPk
hycgFAhvpP0AUyIRaLdNiOun0lxfaOzenFyvgsmRsO4HgMzd2dfnWhq0vnNngL9p
isSav7pRvmM+FiTNCbjgF3iwstgnERFQII+qdl0B+1uKCc6+IWmUYOvDpF58doyw
oX8V7vC2jrZhNaxs80qme9Na9LExdt9LN+0WiN4MQTtmfiwihOSRvk+FTzHB708T
bEMNY64IkGLimKy13NwzlI52kfAOUfM9ZpVeYvPYHl1e3xXOBN8IzgdCfOKwfZmq
A/1D/c9i928DXqoWjvePNOAd/Wfo3wnfABqQJLJWQoPst8yZot0Lz21Ld9riV2Mn
eAHRxbqMnGMgwK20VKlgwoqkqKCw19nSpui4/+u8a19xqfrUPL7slboFn1Jz1Vc9
OFvZk4A8+yU/JaXVvs8qGKzXYxDnDxOVbausn6+axSsDSY9uxQLMFXoSeZlQvTZb
LgRF4nSGiGutlM2G3B48/FqQDqwC8gKB0cERnnA+DvxR+0nlXttDy6q11PMRg/LS
vyWYuDH+J2gOrG8a1JMDcAFBZHu1LCMXJBY5U8zTbtv6tSV/EESqeSsXLlXev2p8
nsInUnydOxrRbg1fQiDy80wrR4HnlJ3WF/pUFnAIm5vLLkb+6CAgsICeVJnZuiMW
sbZvuRnuPC+i6T87M6Xo29msGojUY4iNu1S6nczOBVF79a/o+hx+cEGVW36Wpqat
1iBGMGeYsur5sCqgwS8abwHrHNdh+oA8UlJ5BP7um/6zsOYbNN60QxxuVRP7MXa+
5SnMv6yAcOZpXV7uAsL2gTffnxHn2IjGbDQ/xegUpAvHQJfbHkuDGwAWdalm438C
TotSKrdA3BJiX8HrzWY0qXJanTLayrKHZVFQZ7JouOTwQfYI/m+CJRNgiChdsS+5
PTnXcU/go9tTkitTZS4WoAtguM16hk1EOWOXtLz2Rc7cVtZzlDW+vATsoDDMdfXd
6ZwS9zpN4r60jqq5Q5duHx4BIMLFtUr60eeBC5uGHBEleOii88A6/kfUZXxtAsta
9ltdbGDOIzgSGku9CE3iCmmalf9RbgihTsLEgE64a7TCH1N9UfRcIal5B0a1chHh
GoLYIaYop9h0AYX3dLTFpdDs4W6hNlbtd+c1zFnAPVOONXgLELPdv5XoNznzldq6
klW8CkxftulMLcUHJH4INO6A5PWYhRrYusnv+FXOh5C4bfFIHuRe859L9IZyiAG6
HLCFJmtJewl+pgAN/zfIzOPFWKEFmHwDsuB9QmlrGLXJOqWcVL35gOlHbWUoiUQW
APno3YCwHmmBU546DVFUfH2zvvCqJZ8bDrR/akw3utxei9UDaA4NmOsI5EHvDaMX
NiBI4t61QfD3A7VAp67RkbE9SJl56H+Agh+XAzNWDZHst3K7dsMZQ1pJ8Nh4N6JP
AlD235EqWtcBvAu0UFIMm42aP6ycayhNDWAG0ttau0Hd8TNtCXdMPYLkXIXluqgp
JgrVawy2OlK098+ZZE/5EacgOxxTImjaAJYj+V2ugoAY442QaI0tFCjHBc+ea3Mx
taF0qJeBa1cE+ztWrwZJmJMQOmGocEGLYYW6BCOeFug6IpRmYrPdl2+wMaarOlCX
AzEy3R1e14GcBiL34Ru1ovT011Slm+2EVbxCMWCHMWcNtlKBabJ4ANsnc2CE8Lgy
j9AMXv4WGdvlWDva7YLec4hYqMkuKkzwn6pQaiQeeYmAtk2eC4sxHrayG7/P4s0F
TGnCdkMw00Fenyb6dH+ZcJJniF9Mz4CuF018SIjAe1UuZIBoN8DDnf3EMj8QCbKg
YZdyjfbjo3dmfoMnyROdocXPK/PodmV6JBClTEAvIWd/7gAhHQlIGdJeG35+zc46
wp/aH/KBr3cks+rETTa1gOhg2pmyxZMQlqFdT9M19v1N6A5jR5WMpLemyvfKYsJH
KNmhld5i9BT4EUDOMcW7MGa143TAnbOnuUznBcbn6ArYnKNCa5Xo3DtaBX2WQ2RM
Q8WBBtsdcRH9pVGuwSzpweT0d7jorU9H+lmS23YAmWsh6t4/4Y2kQ0IMr7wMdhT9
5TfpJrvHY/zyL4L7IfFkq0kOSyH/IPizz1KwwnRmM4ni+AvYdjPUgXwHBFcbBdtx
nt9bD9RqoVpNzK6/RJVcvUragX1gGpULuBoX4wdTf1Nbte963n6f8eAXRJwYyktu
CyWcbRi6ty4VgtKYwsErJEGZM5kwoVb5pMVNMXhBcOCap64ylPo4YiGr/sWqN8o4
WSbyEHlb69TerwOU93jpudQiQ0rmRIlvgEghc7000/T4+1ZdmyDecl54sVxJSetD
3tVootoXn2vVH1npVAP5gHC8Jl+lRWVd0wd4x+fEczYLnGK7KDxnqmZ1tqOT1m0h
x1Uae00CdURQk9B447f1uWfbzO3t22G+ckP7GQL2ZHU8eyNSujnGytwRk/MbdGhv
OxRAo88mhCFHLyu7fIRBUBInOsN7lspXhLLZvwvSlTc8qArVbH7tA+6mDSKvzOqg
DabNqcJG0PfPLCfTknElKjOIZX8i1FK45TvGqkAiIZWGkPYoJuUEudFMi2exyNnp
2kEV52mQ6AWKwOW/oHYYWU1Pi8QCFqzPwBR5STeGO4VH9jawGKvZ/60JPQmqsOJN
QNhoOCYskAxDi0SjheMCltJoejN26VbKRPXfDUAAT+M/Th6mapKszlVedKDahgnT
jlNrQqQR5RSBqlO7/d6cCb3PksDpuh2W9/5ag1EtbYNaN9Rn1qGn6AwYvIzpdRcV
ghdxRD8RuVhBoIpO2s56Bu2fZsusYxhEycccq8qbabXI8mPMsJX2l4dJua1u+PW9
ag2H8dC5bNZMXqQLU6wXBo0q+zbnm5CenbDaCKwvn/SFaTCAmKm50h6UIl4HwOHh
JTRk6gjyeQP3UMKJBfKoCB1DNtzAnCZTRYMkotg33edYGBUhOIuF3nYtCv0wtIL3
kHAElCYkTXhENVmTIjgr+w/FbQC8fP4DrTFXbDjC1kGmPnCKXcsVVT3S4VMtTfVL
/d06kkbMEGn0oF6mUibY5HEbEtU3xtf/bMF0MEgTNtwgxHRNORMA+l+ry3SA7cJB
/UWonc4Z8Lyrd//mypFGJtwRyQKj3Z0yRA58ZMAD+qosyDZUp8DAcnkhiAUxtNri
NErcfnP+eYcpGts6iY2OJ6qZFfUrp09FZDx8k7PVJIPnhslYewUAuuSv+2Bcm3tx
YLD3EOP5rshRoKam+nAVmzRBTRzdEUbDuohaXKkpbW5qHw0TcsOmUNQ14agNPw3r
diQeGpef3+0aCllN/Gvaw+/ph/XMBzJvRfqCLC4WOHKp8Y1ChfvvBWYIU5ft8UIc
+jCsDrt8clTaQBx159NkANSO0gl9IZu1yUlcEL+NCsrtHC5G80PIiMYGIfLpbsa6
J375QSN/9cH1hkqU6pHYgVqdNe143PjAAWU8d2DEwaUKtLWbNnTCEMSgWLr9DBUW
VUPgMDysG6pDD6huQXklkZPGnVn2fudeLlbkMwDyaPg3zwv6BrpMtYsF457CK3bT
bs+7mlh+ZJoS9ra7AJEnhRrxXKGKzfHE52IxTwkXzylXW42+/APGoP8JRR8KwLN3
BCvyTvyQaXX9aEODHwTwF6xPF8i8RwSQgaYPJpQF/8QHQeHXz9b7PP+GGWBdcnTo
Pt0dNMTkX3+bg1MSD2IXycp/V3GXBNn3ohzCg4tB4QiyEAq/38BJpp7tsLlDlL6t
Ye+Du/oLUNf9vfHbfURN7UykJ4/AClH6oMp8AvTV9hwwpNL55haJcfhnV4GBq3LL
phmmoADBWUBcE6Wh5EKbZbiTVv8e/Q8ucUNlFyBfrnE6LxQSMl1hEprvi12XzGnN
KVaeVVtJMh9qAuakvymLpss9DwQ6eGQkohQclK+6osv7Ox1LJEmW9Ltko++x4fK2
49YbxMHCDomQ1Otq8OVmGe4DnQMggBJ9A/bAWqS2negr9K9nxAvH3NAZp6XoPTCU
9cJs4OzaWzdjdgAjEUNN3TpOCAP0hlzoi0w4Zlq15xzuQsebKxSnvnH5s5jWzmTa
PNpKMT4VjB6gOPyzTA7zew+lB6hM0NGnLzFICA+MA5zMksvXhBTKwjRLuLbYUBU4
bvnrSfSm7don2MvToy/w1IuLEqw3L4FcM0ylDOtGO9fisHSrTLIaXw+veL2Q10WC
hqHek+C6RvhiHzRFSbOCKXo3Al4MUG/Zj/7iZ3EW6JWWrRDKEk3UcJuDnbmGQZuF
7ch9bTdKxm9WCnF/Zc1zYW8Jlk5umNs0RRnLehLdk+Bnlo8m+ggkAXxpovI5lTx3
bFIToCYBwg0fluEFPNU6UySYXQJxwGvKfl70cEHsYxJd3NZ2miiAk8hmqPqQP9Ak
y3CPoqxZaDWMo7rqsuFo/gq5tPfjZsvVBgf9trVAqEXNSBFdUJSKGVwMdVvqLbSu
x91zpFDBYTsOSuUiS5f61jl7oymtk9LPk6OP3ZsRhR2LARKUE2IoWJPiA81d13FD
ceE8zGuGyOu76Oorh1ZleAhpKaYQwuozpDIvjMyo6xYrnhc0YqgVgHzB18NvrwfY
W2YeG4KspjWsDWNhaXeDye1s/hIBRoJFKzhHFatsoe3u1OLRsoLyRG8Ydfp3pwLn
d3i60f7eHAkW8tcWf8VcnFvHv0OZ6CLBsGuDe2IS1qCZ5ksaQtavXAMfpkSW+52Z
prc1JKzw+XhSHd2HmYB3OOR/T1GVOUTT1BMO7PQJlc8=
`protect END_PROTECTED
