`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BQVs7bwv+qEPWrUDLixka3RnU+T0aPHxZ5lGQgCfVJ1D1QgZImDZDaNDoTagR8wM
qgufVD1bQ8x2j9h4eR1QCMXRwWJsGm2Q99Sy4cUqac9oLiApymdHikRqcRtxfSyM
bIaxq1bSS+IsZM1EeJj2gHeFcb2e0W9HunMnAmjk7mTGJajAKobBkg+E+V4WDuBx
bSfOvWsBVbxsExhibp9OI3nNHGkccPQmNscnWjl6FhUD1nWxhcFxzCpwPkLR+5wJ
rPbl8IJX6CBCf9jo91gzIyJRbamny6yAbZ8/yc1P60VL8QpDksT+RiKHvWTWpZkY
tToChvLanvWQu4syS4mOqD+vx9VhJ7oxJEhCisK1fmsI+QFisScXC0Px7GCA0IjW
EcNlEXLFogFPB82IU7FFfzmny7jjaI9vf8aQk2iUo4d/ug95m6qgPzGuaDTA6Rmz
gMwvzoXXzK9qxIQmOj6B8b/kunRveUHeb+A671djoA0zVYIDTwpaVZsBeypy0emA
2pXG9VBzIQwVVVnfsnumIA3epyU9l+41c0Y7ulukeRn0nZ16lT+JwvQ8QyamLP/J
tpNmXhh/ePv/vkvfA6iGSLHMgma0+ACxnB2g6ckGu8UkTIdaUrcD4J7AJGQLr0LW
TlNyKzLF76u6GSgjyddtXTh2HcQQTBQ0w0PcDVamCryiZrrxSdlg2drRbpERV11E
JnbxS5zY9kf/YW/KhB/JLfrGvBilIvYRzmKk4l8/wXQKQbkB1NVZ9aLLw6Vp0Cmv
BRrk3OHBU3/y1sEhquYAnmDzkrjaDaLEbfIbgzK4jjcm0sqxetQ+z3CYHdynZQ0D
dHqbleN2wjdjgnrVrgXBs+xNp1J3qRTXY1aBVTWWlgwrIKGLU8SgoR+1e3HMJWw2
wTPBNXd8tmQeSuiv0qz7lwI6Oad6lwfTzAQ0ash38kSwBrEukwn7iorV7nuCmzM0
7Qj3UFOTfBYRSROpG1bb6c6NksP2ZVIrexR+0rIvSbljdh6qjS6lQunl7jylubEy
Qv7Bzauf79tkbbgMh+4kB+KmMZNdyyr1egifIqRZ7T3dLgpdeikx08WoMIONknB6
tezIoRNn+VaksLkHXiQ23g==
`protect END_PROTECTED
