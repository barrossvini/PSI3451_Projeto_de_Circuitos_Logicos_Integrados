`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FIbn78zRw2XzsdJwrW1SZtoA43FcO6g090wFi6FrnaIbiZ6im1av98nlpkAWGJ0a
27/qrnKc9FKpzM+QcA1UCDTP0TwWOkoGl40WtN6p5Z5aus4BI+AWeaKppv2yyTlm
CbL7oIEMyzMbvmtwRuqrd0tIluM2ZzUHRAseaAxmsr0jQb++Cm7bEn5WAH6XQLpN
OD/N3AP1DeDM4dHjnSKivfwigQrm4/kEfJhBBZ7i9kHPgZmuIV5wFolpTu60DDAt
fD9N2MUnshGrgduC2HJBdZ9F+7IPN/bSxigDan+bXGK+Rj5Pm4HwxWpcG97VH8C8
2SAhsjYi2b0QU/WRWc97YWGCwgIYTDChXiaJgRZuQMRgLPzcwrXZcO6Niz7+uB9f
ZEZ3aVqbUS2bhu5czLCpomta55sghP4KoEio5aGseiNJyIdaNTUB1JJ1NVgZo+rl
oWEouPCAc47g7Vg+Lu4MmMREzo7qH4KJheqg5gXivKkxy98gdh0TgdK2KIkMjNbD
GdCuBfBNxbP9EL5BSPBQaX0+D0fWwOY2U1EBnZwr6L0+bCyaRwhG8DqC9sKfkRBX
Lu+rvfxsAZQl0N0++2LHP5/ijuSOO7wSxYb4wXLXrdwsGlv25ypXZy19ojJG40LO
3AP+HTYD+BqQpzTweQKwj0NkAFKHB1xpbGKngwvNpLlbSqUHzGfb4IFU5klCrluj
elbDtkcIuHVf2NjMHUrQWaPKlgVVsBVBx381UaIYzyh8U7xd198LjWMN3NE7PN8f
ibW7wTErMjTtLc+svSe3+WTKyKhh/0MKHOhdWI6NmqLr41XU1CXhszUhJYQf+McO
L5berWSDW6f0nNSxtfVzj8/LakQLjz/gIItMvwM0vcwieIybVeLtXdF8d7MEFgWP
kfzfOuJWVxei0Q5N9+YoZdGH0GqT0dnhC/uBUqsJNIm0eFuj12NavylScUkHvCLC
QyD427TX+zfiojlP2mz8nywQoCme8TQkDWu5VjOY71DLWpZPidT74eGmvXp+X5eu
raLE4j6NvbrALJPxiIUxZ02TtPY3ZphZImsEwi1//nEDbSwB/PpIUlC6k+RBkZbb
pwThPoFWfPVpRpMIuqnbNKWqs73idqgVTNjnn772V0Z3UH1afWj26UkuaM2PjNdg
MNbm9VSVb7YjtAHeWIG4ng==
`protect END_PROTECTED
