`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HraB+G3AoAhAPDPeF3mHjqgir6SXi9Vn34Yq+YIBt8suAxwCSlExEbYcrVtVLAIi
MJD8TEkQhDW13fitViXLANhVBFgGuHJ6lUqGkdNpnNO0S1Kpa2Udw8YQCBCAACZ8
ko7KDvl4OTX46E1HA5LmrACEx4i6BnldcjCKaoVIVZASK8vbD/dcwGzLOuyyLyFN
XRmdr9xvvY7EARDtm7O72O3pTVpa9j8Lg1x+I4RQaFs57qYy4e5xXJ3gfCtEXnCE
hbty8/bpPC1yd9O+godmS4sml7eleMzSV2QLrOp9uHPMWWCWOg2o8a8QG5kc3zli
R8WpTZH/cG16oJaaPeNMeuQ0IdVzC+EgTCo+JpMAIEVE3KpN3xsG7RBSG8/itzI2
RHNYjBZnL5+8mw7n+hZqK8oT8c1+PE5lvG0BEt/ypt9e6v+Xpq70LvIv5/vLp5eN
DQEEcDGWWumKaTQPWqri+5WmUTj4ZXanxFtjpvfnTVbYZRp0Bw426VCdfwsO+fxX
5eG7UKKPDR4WkdxICZ+y93rNfIphaSQ7/d9oVxs/K0Q8zLsD4TQuEU9fIX2Xg9T/
XnyUdFxapnYnCsrBlQCUK42edtMwcaKIsnT8RyGULSRggOaverFiSmaSiEJ/ivAF
tYMiHAxAgEsUY4BM1jfjhN0htsyQTOmFAVV+XGP7aHrLwkZR/+ILFkiPRNfrZhRX
+zkQvqWqe9gnHjKnc7L1GJiGanKFM8MjTk8Jfm57E07D3aZ4LUIjNiJ/cEZ9Etvb
XTDwnkrNIAcc+rMum/JQYeHKnjztKd0MMJYYmwXEwDNaL57ZZlu2RilDx8OltLFG
S7sul6Z6WBl/0iUQ8B1Fbvl/C4nXEkReXiltQya1yxdYWsQgIX75KFjaIEFinZnh
fMljLjaJdz74CmV/ToMSoOwEUsRAE+sAzkoWKTiJ0/ah7xWtBxJC0h4OM/4dmxaF
ksVeU8ldI0vg0l3jmtrJ7ADwJ5kh1duSKyeYbbURbyMJfRh/luO8dg4MSjmbLsLN
1a0ryFy5fCyFqJ/TVpm1knpWvu6NqIpmLf9Wu06aTnXk5aY1qDASknsDEOVlbQO3
6oQoK/C4kUBnhZSpgkD4Fz3lwCHSgQADoNam3f03Ouuwumkqk3eemq/PWi2nlY3a
lOOPnPG7IQtaFi4VSog7JVHJoS8ruMo1xwp7PV5AX/tiBLfiOBWRaIlWdNJGNNwh
RrvkPNCcJcRKlA3Fm/3JWLQSeC2B3ViPZJd4YaCyH9sNUPyXMpHOkiPHwC+XYiWM
HMToggE5us53JvGOBVFJ9lN+8an1O+HXu5K1XfdPRINrxa87nKwBoV2ZFRRuTSWp
oMTUO4BRKF0ej4jCxnBcpzAl+z7UmYZgX7laCxRYoetx4qssnkB70BD7gDicTSQr
EvMmIyfkc9gm10cr3YFu6DwXqs+pRx3L+9Zpm51vS0wqZbzn6GCHr5oe3/wndvJf
tJebS1/MRhEPaE3TY5zPMuhTjYcZlXBRJSwwE0Gcd9bKRlSTbOk0qEH1vu9+6dpc
MfJb2ImKDTC2ipHlb52CgjyIr2NxPSqoc3Khdo39WQZnVTFkYwzNr2z0lNWOrPOU
lKNJBap26gYb6NncO+bPnRWr0Id/NeWhVZOL07Sy2w9cDK57RGo6ER2NIfc++Dn4
VMniPxmmm86Ux5HR1zcrLLP1Jl5iNpQEDJRF1aafmsLo8svpfezNHJQ0SDNHLq7M
OzKU7LOzcYbePGVriYqhC4/SptnyrbuLVQNbCgLP0RKuC0tc/fBalKYVilNhF3Z7
qvGmkevjkh2gFI1LvZS5tHXLM1TCItLmNxoIdufO5NsUAiJHS9DwR2e9bJH1TLFD
fdArFMCq1GGYN16RPoRfLIzRP8jYznGdRiYXQsF9FGaHA/xfWKlfeVvF44FxVVai
dgn05fEE4YFfRlAi5WjQPfnInYqHnb4WEzPngaq6Y/zoOiPWL0jJr063EGAwmb2J
9Lla17xebR/MxsEENXf+iYx+JlTK3S8BDQmR0hBVGSnVku3X3a0kgF+4iuV45eZK
86N3NiCUmqlYOTWNSlac3iVnoE9OpFXZNYPQHir7Ituy8ywILH33XH2Lb04Y4Pxb
YfIoeZ0kHcEfOvZUnrgfVtRRyfD9Ec0W4YRsNI3h+nT73cQo+uAFehLVvvVMgPI4
1WrsZlhW8ogu8mz0G/qJtYqs5XsUMKpd+Fap79T8yLenkSGoG8mgHqgjnEp+Dq9F
ZtEcN+5BpmYVFrWI6AQ0qpB9FpFOugE/B134NLMwdF/Z8cPhOpZ06K7HMO5PVA+K
w+ix8SQIC6PeSSnTL/aH3wKkfjuvhZ/pCM1dHXvVoWi7uxpv23kiEbLNyn+eSHys
jJdO2vsRvjERHB9DdLAAczfI44HSeu35N3d90K1KsqLMxf7LFm7xcdvGTwVrN4MD
HAYEB9gDjclqUfKTkwuONzEgQQTA4Mwuhje6/7qQ+Ae5TUsYAA/9ulMHqOu0B1cp
PD6mWSVOKiJ5ZaZEJHW/32BmFHmxxn/lL3HhQaJEwqc10ZToX3VoOKH9+fArRLgY
GANKzeTt1kmkjMN/Nejvq78NM+kOrhq+yjECtCD6BTsKs52h1K2nLr2jyfDwk497
glUPdIV3TrGXOQQvP9CcdsMGu4PjOuDH33fgH8mh009d5cAgXOZdPKkECroCz3a4
6sN3Ln+DN+xZyNy6yQwpg/4mGpOCNQKKf46ycBZq2oMoC14u5+vJMM6wym/wZ1Pz
n4olIoWC409Jym7pellRxCqRM0CRTbWygCoTyArTpjTCIftd9RkqFWDgxaM5FoJB
Nf/E4GjiQve6jaBy8SRgJ0gV34BFx9Ovf+rfPmwpoM+6+AMY6uLjgLe5OLjXNs2z
WpfmSJsBmzv3qWkLQSZ9ShnNPGbd2byz9cfUAyg2fxZt0DLacvPWfkwDYSLbM3GW
DDtAI2Beu+F0ZfvHDBuHE04lQprFlEieok70ZA+UA1RAUjCMHL30aEFMlzEWJ6VV
egdOJ2qg98oK0hZ9m/T7XTgN1zvtONU7v/lsLhs5IIs5Koo/Cl3gcbnFaylHijkG
qSSJTBclmDwdqjgqb7ivwLdy687Nc5ZvhLAmVwpJng8/UwLNwL5NqjDYFYT9DOvS
gt8QWakgkbqjDGuChSnEizlBcWmIwoCt/k5n+7GeWILxajiahNbJzxCBtJ3O4zGt
G1ngFOAvI4P+YB/aKxonVca67J3t59idZ4EDagYA6yBASQOUeDQ1olL3vqmjcwHX
pTvJuTaflDjdV5jE8DTagNdjWBbZzPoNEJHNXFO6RJ+5oFZCuZ4W9tg0kA2Ys2mp
WwtVInRbiP68Odr2NcthX0qlH7gthxw5mMt0LNlYz0U2hsgIwyFgmAH+NoGfOBOs
9Ub3tZbOP2e33X8jHzJQHjC/gva/d1Mxsp983a2yhEGLA8RYwAoxTVBQuCIxH3M5
DD1moY7ii1Esqb2jjux++trBEGvcJO5bXbAZ99q7VXegVvVCVO4KSfuKW3qTNgsU
7k2sskhHBhFyf8KRbRil8SJXKFAtr6NGqIWszMGX6USH/tUM1YkYQ3REKo0Dawco
6q3T+AEvl7K/y/LNNuTKKECn5Lpf1xm1hkH+xDxjOafBfazEuKzU8EuWqIjMGr98
VWKANctMDOAzUaoaTWdhR0Cb52M7jXWCTZL64Efbs0rFGSmRI3iMefzrsx73ZdPt
i0oyF+FHtuguEVLKmLz6ANkIfzFtJYWOCb4JwrdOD0kEgyrCr+wzlr50a6RQREvc
JGqLqp1CMAgIB5lfGk5upMsEBpIni+Vc9EmjK9HdX0ngPucv4osKgisIPNI5QKTc
4eiAtS/DOxe5GBfkt1WtNS2g5tBk7cBRts+aAB7rH0Ak0g5NTU4DbJPTNTueLhTG
f97wtd2L4S0Wo0DcP5RrDhgknxhQl54Fe6y/8gHjON5k0rI/yJB07i1p9af3QKYU
7D7IAwNy+Zzw1L9QuEGBdSNInxZLB9oZfQB3Hx1ga2+jhW9ncii8AyNphG6mu3P9
M6xoq9aHJIEf5Gqv0Rp+C6ThdEFpyqbNY368D/QD1L+QkJvd4uxuKu2Qj7uGbOyW
us+iHaKHgS4buSJymo+gDSfirG/MbA/Jzfm4qf1Bhsb13B/bxnkJe57JhmUUa61v
4lspRPXw6btGPGldH/gn21luzGa6ZGNrvltgXw/sj5RcyCi4xtIdpjvP2SWPgkKE
POOaDKq48heEvCEMVIEE1U1dBveqdWLmxtF820Rq7+Q00kzgKml/bmFo7EcqblmJ
oZmtb2Su5d9k8uQIO6ioZ1jN0yH92T9OSvxJsv8vNsFbNuXq1WPQbeyjcIZuBCo6
PZEsWvxoMqmcY9Gv7LWjw+1sSnDdVp0y370Zl0qiwuJkT7qF82Hz6w8IN4AME3Yb
3YAGFrTTLVRq5j+Fy5UH8JZTtss9lBOTs2SQu4UEjKaEwpaMSbSNVDzMS7BfCiTL
WuGAZn4hrzxrxQKJl6gg7E00SDpo6On8xS2IBXyW1JsDTc7kyGBxIjN9lkdL2Y/C
Zhc3KhIXFhsqyP3Ct4adDRkiE476m6yLEzJc8qiqEyNe5xICqGH1DroxwzKckqqi
SJVlACvacrpAmyl7/VN8xMKuCw3ZYueblyP4nsaeglXrPmD9794wp++G7AaKpwZ4
KeyBJfUUj7DYoQtguBOu5VyVmC94RhYUSXWbaim7+vhK0yLLVpfXa7ACPUutb+21
o9+OJG/t5uQlYujphfev7dNVvTMsDxIJFRhWvmSKlqIIAe4wHUKF2wofw/ji+rfY
G+zIn5Cs9edeSrgVE1W/Gz/sPemjxDa7Plz162MKvy02fMoK2LdcfQSWezwLDzfu
CB7iP5YEBIo/nw5hjc6kE97PrOJfsBXuXiVNN8lvojibeHi0MPGA3suCTY8wNXfX
P9+LdAHbAPeazFpZVc3wvK6q4fZwZYQLNKeAY7Vbc1T/zv3gZflxrYFFGAJjkFMJ
NK1gdhgHLPd0ICS0zgl8B2CGmjg5IzgKwMP1C7IzqNNK0hSu9PfOmKARPMfN75qZ
XftVNrjFMbtOSJX8dtgotS4pUCTeM8qQH6q23Y6j/BkfOnXLYdwnbwymnQxDVkF+
NRSOTip3xnm+8femwqVHRtJJYpEO06CZVzor36xK2rHfI93wG0rwuYdrGSDm9WI4
IpYaX4G5TUD2rySjbdEbch0onrbkhlS7VU7DEjKsTH0I6E6gY++V+jOt+kjKXl0n
z8IA6FmUKXCqmGcKD9qSXU6wZ0hE/twGdx4v/EB18jNPMdwNubOtak+2nevZayd5
Zn5fWls7sSblmy1pHhPydxRTUSvTk1jqBSUtgICObiT5qxmVq9WHsBAMdY+Huixp
xqyQ7NLNbmhNPTmvQ9DD+ooKSdWeI1/fMHmSqU6F5KwlktcntpgaHB/KYS6ML57J
6LOzeMLKLe9P1gvQg5dcjyP3eQUDGu8hoTM2p29UxtlFAPFuVW6pqggssi5mE+RN
WOptjAC2fgMXusH1Rd8U+CRu73QpWEUBRt8RM42tEKvw6UFtZB6gA8B7oLzhFZhu
daQuxsXaxKjaRoCuyWg4PFIwpJFa7o6/vicAR9EeDgnV2abv1Y1evTFH95eZsxmg
16e2SMfYTGZwd+IrVyRsMSbcZk8SNqAo7sISiRmZJ7uFUiZcGugKn6Pm2En1xI5x
QyoGmQjLBIkVrn+AY/ZyoFI7dUnXBh1dzNuPb3P6tha97qgU+t0AJgo0yPb54R5T
Vuo+MYc3cwL+3uPXFT/AsXrrFSVtsBOX0LP6bLKomCEWYuKd+ayNEf1nzTiXpVTs
D4bsJbJUbqS5atQ6kZPpQ5RWMJ1A/19mj69vDvjJUF12pzqUZRlLS7qzyjQE7v6N
ivFrGVpkeIyDBHdaR7PHVr3Cg8g/JVfjVFk4m+fz2aqh7kTQGq/DQntaUCh02T9u
O08l2f/H/ncmXDyBaFq3Ptwxod57tBpJ0QEw6nfA4vD47sLIGA7/2rjjH8+bNq2U
TEWLv1lAXH14D2e+q8suq2OIj7MZR0Lu8027D8ZFRb2CkIjCqqwMJj4zJ63zDMdu
tooKvtPKSADmbVG21KzcJwAs6JL60vy36MCcaQxZsby0W6C5rqGLGe1FekpC1m1D
VCjFVx6D+jBJJ7H7j6KOfrxlKxfDkj/dPikzWxQaMoQo9/hAb60+C/OVC9WBIUGb
j8Td079frg+RlzVKXGeMyfJqvcoeh0NZWpkHoVt7B/dV+lawSoJzfptcHhlwvWyO
Vau9ByKl1dUcefGPv5yxMCQOd434oQqpw11KhSuz5EcrGbsjT4WOkeql6/CnfmAD
eCZEg8cXRwci3zjBp6Uh8aAWdTC2P3sUNNI1uL7j/DQdl6wVRoEqSqJgQpc1f+Mu
d31mJVbSRKBYLJtg4iyT1k69PgS87SpkbckJ2m3VHnvCspXaJP7qTXR2JIrBxGmR
VrkmpLzA+xn2Fj8whOViKKQUG9dIWIBOvHhqeLO43D7knwwW4flc4tMOgc6QYZXw
Z7iXQZGAnpecC/svgEF/ThMGCOyjXlOvSssJmiVfj50mtwFYDZ5EX9giKLdRP8+x
Qq8YRT3jfRlQXpcrIzFGz/bViUm06SIYM6TlOJZmTKogO0KhGwtolduW5fRQSj1n
xut2Vv4FLJ5t1/NrLI/7daixEzgOQPAhbtZoyWWPe0hwMB36iB+ULvUeNkKgbtE2
amziQNgYHRNVK9Nk3FCJh5V4SbHVCY+tL1b3OI8I2pRkydGUJIvt7DVJyhlaHimq
p+UeCfeOedtQlOUFEuiljvxHkpzpOcqsgobX4dkCX0AkvOBSgAmgzq6JHVAMVi3f
KEShaHYBrR55GBwEzeS+yoNm5wBO4eXbU6ISJ6BCcQ1MSiRzBysP3OB3aMn40VkV
qmovGGLYVHLhbsb56ipaz1BVDNyJyuxZK2oOmCT7UZffiPd5oBoY9/7MbU51QRG3
UNExJ/iGlVq4efEVi6asyeT+QdEFWV/w/7tP4GqLbz/WDSB2tlvGpGQQqP8O4Xgb
T/yjXt4QJU+zuF+15sITB1KPBCCPO++CpABiAFy7HXkB4lhEdWPMVg9oUZMl/39l
MmHd9S9JzoPxYccWnktHl9InvAnlj0pFHNaZ8B2wAl+UR8lcaKcw3cBLJl5BeeGd
hUf64UAWE25eSssz+9B+QmV/cNbkSq0eYJMfqTv6tSe68a74ZKHJPQzYN3kx+viJ
JY9g5OJk9aZMJxTTnU97nFTiBhR0skYQyXkPVMBGGDP7EsD5o53VMdwgdE1VBxxk
6mkhqIZh7TofKivvygTl9KGqoOUYUREP/gN767IfAzIdT9exEkCpOkpIw3OlNR3N
kwzr3kas/ix5nTMuSlWuNmu9SHWt/CibuJxlOGLSnuWSnPqsxEl6ez4NoHSiZbik
vlpO+ptbV4RnEEBrH0bxQOb4/47+LQrWN2QiDG80XMOduASwCEm3cz30rngYeFoC
hMAxIOX0J3NBdxVvk1nVPsKDbwLz24Ld74Novr3NnOIBZM4DQnziAipqCgZbsmrc
TRQ6ua+Obxu+rQrL2p5uF4qCAfvDwv9U+qecadgF740OLnjaUDgvtRojRSTcvcQ1
G8/1G1dDBMGPEbuuc7eVWVs6VaK8zm6vNfjk6Dc7cU/M6/pakQXvVUCxwTNNvAOu
JP+rJJELAxewL82yzQKETDu/ina329Y+2g7gpz6i4FJjzgLDwm/39MDxGHT/NvWc
QOyh7VH4RtEaBw4n31YnjnU9W/6YXQK9bG/JUZfEEdpxKixMiS0I9en+pA3p861J
wYpCFZ9AuvTZTRUdekozKy8HUFYbsqWu4tGZFaFMJ9NPU0xjNjsMip1bK9W9pAGX
X9aX2GmbTZoJ8X83JCn4ZN3m0FLT/xstLPbHr4vhGrhQIAQDEdAA+fMnJX423jG5
73zRQmEkww9IgGpigrX29qovs//YMKQS3lN+t0SQj4FXo9h1t5mn1ArsafDCBshV
j9UtUfAtkBz1LWsRKdZTfVplGyZMn261lZx6XdKRBaECkpuTPIU3CQl7wsWczMXQ
fq1u1U8avkjsrT0XNIECsfygUNQUZ/ccdOQHDjiGBXvGzzMiTOm3iHQGK0zN/ntr
c//pa7H9sOXCayUqTDEU+8Wek7O6vG9NSSrKXe7viCmaEidYM7Axf5X2tGojYdDY
AYVtLlh6/5937GtyUa3QccQN++xw8gitJiDBAtlTxUEgdE8XQWbITqTbEoWH2VD2
Dme9xzQEt/JSJqE7KHL/ay9FES8qoFiciDXdQ0IpTx1iaQHPUAbp9BB18o8mZ+uf
oLPLn/XXBh++StNae9DZ8ea/1i6ARyPDFRCMTmV+9pP3LVkK/QxAVS+Qu4p/v1hJ
7dTHNhhKcYb1Uz15mMFYyrjKqgAAYmDhgSbh+iBz1NGN+AR6eAArDAcTupg297fO
4gOb+WlZrAids8stSBLePD1EDce7z6FQ32tLRV9tV7Ibg/4M9ybpsTpi6JUkNfjm
axb/RTEBzAo4PpdyD33sDNlr1LY8j7EJfmOkJEajQ9CK/Sjowe4BQMFtgCL9w8e0
ZVghMU2K/lsnSR16WEDc8Qx7+SBuj3RtUUC2GnH3byM4mLLC2dvlK1fbIZn616SN
QLduSBdbyOlkpetgzyuY9MaJX+sA+auoLIqBXR8JI+sk959hk1Oius+iyeVRva34
ZKOeSe10xPl/3NFxcnt0lCWjIbSoC711uBzsoG6ks8Rlw3j7Ocy8JzZFfABRroRE
Sf3LEt5U9DEWMEr+ecHI/z4B6zdy/eorhsFFlegug4tMe9O0xMILvkdnEoBZTqLt
UqKoiemub7foMRP6THwoKeWiRtemUobBB923krFIi2kz6eOR20bbg2/sGuW/oJF4
TObwoe/QOJahFPRui27zrwvIIE1OXro5dDzNFR5hTkgaZNNNl0qsMDH9nO/pNm7f
rwBtrBfX6lu1VdYEkgupLv21YAYU/Fhsn9u8e8KFfyVoVIj2C8Rqck2quftxcuOe
gX77b20FWRZSpC1zCAQWrJMknzlxdhp8v2iPFgZ1r5YUq5ngy1uBSjri16JrW3rh
gBcPLT36MPtBQ0lYCTkc4tzM/T1sO2wAQW799ns1rjEC1b16aEm/orFZi0wdC8JK
RlAX6CmfOiP0Rs/WTOMAScIFC94skOu7cBRQ/EpCLnhvge4HsMDtUOrD7E9mnC4g
BVNDj1wgkAn5P+hN6aj5eSG/q6YqZ5x5IhkLBm+8DKjNlqS+2g4ODnWUdcD+3MgN
n9LdifCvmeuCvB4S4przMiT/x6DbOms0xpH5W8HSIa5ggcxzb0Fjji9zv8E4NF+C
gEuftAaUWSbBzSG5CrtkpOjrOIGqGbNHruRFZkhOKrWWIjbbV+WHM/sWzhM9MBJm
WykGj3xkR2ZSlLKp4gZZjJO9Fh2P/QLe4HHHrUcoRXmf7aGVAaJZJh4U0tjH9FD2
cOJ7Y5WlMGS6Vp+cUv0DARH8B08WzNy9nXtzLdBwgGu1uI5lXncI9bMRnX/eeaDu
MVFw2X47910yxIT3eGHA9cSAJI2K1aCF2B71GOJ5Af38T6TG285pvdemyEe07H+8
lLWqI0jebnCkT70mn8/onGTyp5OMQxZq+byvCfWwGbAM+NZ07Na45Fe9vwCiVnj/
F8KMuxs7IRzkGZrKgWs+yTfgNUhB/4poPqwI8IBRh9PdBqTzFoBVnJRuFKZtoiI9
DLIejatOLFwim05WiSIVCb17gOeBzmMdXZPiBetSPQ4FItTNyap/YQhEebSK3SiK
L2aLeFKxVSelj+ruUZyD6FloEWvC1rjzFrPX4nWY8Vl7zWRT2oGpxca0lJV4KTc9
J7e3Y5p8ZwHdxJ3vr2mo8SGQPLJZUBJRMT7Giwr9b4GUj840tKfX0UP/axn2lOe+
ybqq4LjbJbMhZ+BbA+d/oysfqNDa1CD4ZYrwzRKoifgqxjN8WUjXrO9WOqSyG53W
knYxa1P6YQL0GbBPzf6LfVihuEPBvs4BlbvoMK8wUdHCnAUbWriV0KMCIW25yFaW
rHtnQ44g/8TkzsgSoXtU621B3o/c6UoNAMSf9eGidy6GsQyVO5Z7UVbIfuiBNT1r
d8A3PoEE9gDtbFpb8B86yjuBiPqCxF+vC31U7YWXS+I1jHhSsS21ihcBtBP4S3EA
EkfZxOd+r/cWZLH7vO54hlFBbdew9ryMYDv7VlbSxcdzOh38pGfW6m4GsBG80DhI
g6NvmJb7m4SXT3FG9iyt/BYk5rlic1ERPRyYvULLSlcQSoXlYPntsqByQALiiups
faoBe4jYUij9IW/yr7SoBsY3x8VrNnW6csli6cqQjRorIqGzqx/orwlr91KH1s+k
iWVUmLDSFVnyXn41T1rCel8/vo5mBokjIbmgQwWEMUcSaVLnt/tvTIbFi1ve11Nb
hYFmEIuS/G99W/XFK+0nEhKLQRpH4XaigbxC/iSEeud55a/fJU7k7+Pfpz/yOijX
zXtXYMaf1MIdhR2hwQKYt0DH7Zu7xEsHsvv5OPb/VHWVLinS0j7g7zCNoyhexA77
dVBw5zLJqVFeMXlqhdbMzp7w6kPtgWEWxwTpCRxSsDK7pyECcdNKEzNplLSL8yOs
VY72niBkqVRd6oYVukRkDayYywoHVqZSpcEteD7MxRYWP2exTvnpi8V1VVoBqJk0
sTYhMATJSAy0rNKpYmg9W4PR/LpmQQdC5CYTZkqDlU8WjOVJNky1X1O+zFnc7rXn
/+E0m5yFMlD1HrcHYLZZGDvLYqwGxiBcod1nTU6pQLjiS3X7mxCmN0GLZRENjBf2
UptZ2JwroGblVmWS4i3Gt2eRkP+jESrc/Cg3ZSiuWXBHghxPjfAL61WYpoSN5mGy
Ux3QRoBcpJFbLFDtI4aqBtU/SKe/DZttLZkq0W1LY0sq94WIh4qFwu45VsY0R+bj
4JQHxYqQHz5CCMFXHxJzFWmuAQbXsNum3icgaHzR8XD3iY+RtVC2fqUmz4o6EZOw
fBkYZa5WXBqdv8aH4bOcRxZGIALTOLCJDW08AsNePZdsmescSRO72hnwM7Bn146v
ycerpTX95yeGWvO6gcmmddQIZR2aGFLwWTcRTQ8dHTBd3Z9QXCguIA7gD6VHMhe2
d9hv26YRhlx5xd0GxSHpAu2nKXH/lJEHWd8NSQwpDEXcGgTolBX8y4HPRujuif2J
2kR3vROqWo9ULyz9eJ2qX3lTt28SXGdOYiO9rkHIp9CPz1URq49DdLlMStLRrrr3
Es9PYI5ZC5cv2YPPBUHb24IYxywj4HtUw1Z/s992xZlnsFWF2RgTSMpqT5w5YJix
IapEwGWAVaRzFCCwJCy7j/DS3lGRedXzlaP+E+IEKnKGg37T8i5MrSStqCVgOzOV
RTJQgQyA6dDvVqkVoxu6bre2EDoYdcVKf0h1Iewk0+NsBmqkkprA6QEVrxGDbZAt
3bq86gBM8u8NqtR8gkKhJ4DzMrPu/4O8fEBVPk+BZgrSEfavk3sLocdnWW2W2coC
hFnCoZ3RtUIaYwmJQWJNoyfUdAWsxsvHtQm5se0LizhwvmBO8qz/KUPC2Sbgnln2
LVo0JoFrvGqkkUr8Cqod8yfTsipwog6CyxIaEzzeTdabaeL8ZrM2ya2U5eGqY2ji
eOZolMj6qgIPjsyvwXi1flbrUMY6TBTk5IuQINpI5S1fOx2TvSL9VbUu02sol2Wi
G3EhXUMVuidRpHw+vDigz8cSPq/gf6jFy2JZYz+7JgWnSgVgK/7qjOA6xIay/ZrK
835hfyaInVb/WNKd11N0yLYnaVy/ttPF3fMQ1+rD5GEtxg2pyYGVKCFG7gmBWNfR
8qEsrZo6p72mRskdi0lcLxNwvCYQb8cqZm2bHt/sGR9QAA8Ki7G4VB0/iOD+aXN/
xTYZoBbK00wSeNQ61H9fP/ho3gLKrWOrpQQRNTXdjaEdtipyx0SKQ69yXBuLVNZ8
zcJgfv4uKwXwvNzmh8RvTAzreTB+h4zidm+gSdfgGenjee1LiEMd6qKwNc7Z8wXX
JrDqAnR46BmFQ6lsaPHxPfZSQxc6QEtxjhBGDN/DEQAR/Ggzmof7cNitOlwT8VJp
dIHA4jV3zcCRgQw9kY7n4TSEjB5bDxyNzv6h12KBb76w9hdrEXq8JMlZypSg5MS/
KSmfWsKvdpKctDevQEBIbt0FlnxrZFjZp2W0ThcwvJvhKEGHULBxX/UW8NjylvIX
IRQTft+s/9J8+O4MWkOfsCK+7iQNLxxp+y3v0opNE5N8VTxpUXY3WTDkKvu3LYHW
z5MB84u1VYXRFFpC9aVnLI8xgX5PtchgzrT5eQshDUpsHt3V0YIJMB0IcKtdWqh9
B9zBBK2FTVyxZ6wtzL+JInBYoeScHle/QakUIF6YqGPplr1+CYF6gtLxvFIhh29T
GzRnW1K+m1m4p/3m/HmCjFVIjLcpeoIy0Jyx1jL8w/MZG33FWGEWfQxe928HpKL5
N9/q+ppAwZ5++JNi/wGidxvLF9TTQxSvriIg8TOsKaCXbyS3ntJtLLzpIvRid1yl
ElZ4KkH+gIJGe2UQuPS0fMsUY+vR80etD2FLnu7WbWVsOTrvL2JNGFn0KThCd5Y6
iBHfAZ/W1gCl4EOBoWGT3HpzJv+xATksKhszIpka3EvRtKjNoTQ4iQFjlgDIXYpx
83uxFEZjeoR7p/p0Tj8UZIkhyKrMD6eYCpd3IMUBqz+1Pu7GhBYphbQYjPMEjo3g
kw8gvPa/NJ8sKerihjyO9jAiZXVyjeCkzN++uuTl7KH7C1r8xNI7EhchS52zhCqh
EH0nC3IEve9Rkia78E9Z+pJANumTPrcVUJSbevj8fxepDheV9JPM1McyEGJ2AFU+
KTwxV8SZFiR5++fBdNTTjs8mbZ7FVZVh2/eTJx+GVwgrTtfiUp1m+q92Ed7MTkpI
bwpMuOrEtaGQfv+T4ZWSQ2mzsU/wXhyuLiq921tsfPHDKhMDdFYWtbZVpnJxY5oM
XUWaxuBcywZY7uaxLpcqCjBP0NAxk7HwhNQPlZrGCB8oe+eAWLgD7J9SN6yJ5Nrh
OGpwKTgMwx3saQvNGse2nB2/8LiXiuljwv7ALrrVRlOxg1HbBtcNeW5qyF+cUa09
yzR7Hna1ZbstmJ1AsjKSUiE8YVONXur2KPsPVn0wkyvEwD86UZHWq+B+OcbPcYIw
3ZCOfhCICsWmR6b4IaJ1CSywAqtvLDlOro9HQdL2w29w8dO6f/npKBhPVhKsY6HA
amA0ltXic2upo4ArQUUpH9nSLsSoJoWneRL2vlmIEcwFO/SsdIl7RpoNWwH4P2kM
yxf70aGq5ZKbJ/biWoq05FTjCT9Mx5jIZvQtNdrlaBTxVXCRrZ2otaSgkCkCtOe1
As4NjTfq/+5aJ6EjMYbwI1okqqSkYkZ/6YcZYYz1Ksmiw9X5dvba1KwhaJFVw5Oo
b+jEam3gTOGUuyK5TgFzAhv140YeMdVlSUeYX8N25skao3SJ+Ps256moQT86KyKy
9VyHBcIWZlueBAwN7u0gfYgJJYs7fhoZmJWpfhApcsmxy46HiKsJU/LxUGivBJNB
35ZPt1zXzO92AMWXsTl8aX0og9MfXstM81drisgVHzBr0ENcj1uW9lWU8/dc97ry
sj6zB+e/2+vqTfs4umT81hcuDsDd1bfiZeJPIyB1QMtuLlwokKWiB5rRmml8GbuZ
YrX8+dlUbmj3XsGVo6hrVC3ofIifndKW5plfxXbRjZtDDsElvxaFKdlgnS4S9PLH
3e0ZC5wWPW4fzcgxxaAZ94v75rgZoFmSIANpS1vt4zqgiYp27b64jhnYVQ3nWmL1
Xm5IxPCTyRkLyD1YQALiI8ZNmcrJMVvF9BTZ/WFifcctoMOdw7BOwlGqlWcD4h2h
LKjKHs22V704vHNh/vGgVhFl8QQUwOVtOhGi926t8I2MyjnOkFdbzRaio5tBsMul
r7isLH/R79cqH7INXSl2+pLbFIDtTafzEjUGz79FB2yA2cLnVIAPasM54DiudXWr
G84ImmLFlaGnWLVUHKg7i1ssemWSaNNPUrrOc1DunhdL8bp45l6STp5UYYxD+5W+
BfGTkbjFLk0sWwC2xKyentqL2A8aqQPhT9L7ahwV9ft/pmIRlDPNQPCj65avUHCP
5LBfj9YrN53Un1dvryClIBFkXWSmGXTvNVW7EYLwEye3+wYpusgIdXoM3MgKXgCH
Pibh1+ExQ0MX2V00X7onQF12vDJogoJyp2hs0mU0CfmXTOHPKBczAgwkdifQV8Xt
OmPT9NnX5q92dXFM7deckYbKCv4kJbKl+8iZlrD+90ZcO4dIoZkWjXrXhK0q1Eht
TzMNbvX5hYJ9tuXucpBP7zCQWBYJrI/41e7IuA8vDo5mhwKJMd4p/Waaz/eS3c5j
zPeIasPWvOEkx1607B4kvYZl8pTj2eyh1cF3Bec6KWubeYn6+JhEh4MWj5Oe0dIk
rOZaCNfYfmuYlx292q9d0yCxaqturQxCTsoxdWf4/15KmHK0pxJoK7OIpjtwau/V
Ru930PbpWN4KIHyEMnBQ2j3mZobgSyTW19dYysf6Ei2vdnIEYFynMi8v+wnQcifk
nngm5+LvQrOs8NUkcMHAbydFUV+SwGHbIviHqglNWieZekh5tdPxGQc376ihIOLz
cKwv2JHoIlOUoFIwE/+iyh57JLIlrRGvivVPpbAPctiytGT34wV259Aa9N8r66SQ
9SNMkY9wo5PY8LdkGwkSm/UIXpHdceSqRDSAtbkyKWi+lj6OjbzYcz7kpAEz/C0Y
LCBxKxKvntdX9ebC6epX++lpho3EAYgcL8mqMAIBwCAVOkvl1dWqwocpLej1EGDK
qz/1k5b2jSLlfOiELvuhGZpbCNvA/p8Mmwc6PNtw5k9WP9LUsv2zJGYvIimoy7Cm
quaVp6X39XaofiiE8qIjEaUlbuFW1D8di9lDJ9tj+9qDsSbDl3GMONaM7NU3kKk8
m/Pp+6cLU7dAQe/dH8P3yZ3W97SeoztufXhCct1xUzIUkQIbfnBB1VWOKfGAgG3S
iazA7ilXaOQQmjB4frMszj+wC+2hGQVZdqT06QqsbOq5iXunqZWD27RQq7Q4kK2h
NYfsakVjaeR7vicOuwJtD24f9C7T4htvGsGrBF3IhAQARbx8zboyx8vdCF0RTBUP
R36HI3R28VxHgLr77/cAxULGPnCJ/E4LFR38ItYadgFHuTYp3s31JSsYk0XubkmS
PvtTBNE6PjRj0ZTOXjJODjotK7O0pd1fNCkHszGhqKhKJoTIkxFuYSqej1e8Exoy
TeRi314v3nKXjRWliUoUbOIuyC27ml9Gtg1QuJ3effca395+MLIhgrkDgH3Skdft
M802HtU0Js8JtgfmZ1/GqzfWl5fTbDaGtwP6OlYx5s1Rx7jq9Qpyow1mUbNMU8ei
q5l6FukbKHcq5rJYEKKt4+a5bXpTNkm3XhjcSPSCruS1IDC0cOJTcAXKlu4MFliJ
3k8ZUjjKeJL+I5Yc303KngsQcUYaTvBNnNDi4NIpiKY=
`protect END_PROTECTED
