`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZ07ZYEhrKVB01M+8OY3LStNA4ClxTtEIR5OXzFcmAYYRAtsedj9OESDNKmzESOP
fb3yMyUKtJVxsAgamFccZDELvve91fPCZNYiuRuRDveQg2Og0CUde2yJbMcYlcvC
8M3XqLJCREf+boAS93aFoaB6+Lcbyo7fR6yrJ3HRrzE3C4BRTDkoAz9SAkEvcGah
bfVPuAWxyxRYH1WaQ4jpM3ieXTvyolYJYiSkI/rzEDEUZxOD4odOe1TOvH7etW4o
njKuyosGXHa2hPXHoT0YmgDgJSD8uW2d638oNJxxWWNl4CghwhL+7IGy0Nhmnodk
gs8afn84nHRsV1hJwFh7raGp/cS5011CntBYvcIWPGtTMgJ8iIDdo72AHz7ahQl5
lEcllTlk3i38j2Dn5gUpuO0xXn16rO8dMIUAtTkltJpcr+xq33rneySdXuXaYN43
oR6dSPo4r8Cux74yap258wcVLwiwLtTLJnk98Q4KFfxV1dbd5Gd2/lchPOhwotZS
x7Md/C0mUDQbyljA36xSG0gj94rnL9dEW0+no6X/nnts3WqHXIGwRcbf4PWPc8qx
n4YLXXlfwUX2UrXx9bvHVsxlrj5Wk4jYza8C2zi1OgzyXO9Zd6ZyCP4MKhzZtVtu
prYkXPZNsYM2KB/QUmnRqlDFFEqxlWO0o4CZQmRBS4m70hYWSaTYSOy86gfdsq8V
t08grBQL0OhL2H3hi+U/tU8rjKDcKT5GTeHEvmXxmIPKONtRo2c7XyyIb0vdIva6
c7n4wvYq0zGJ6+qi2zU8fZsK443ZBDg36/DqB1x9NXgK0fc+3NmpNoGrrUz8G453
2QEJyY6OLiQNirqXL3q54By+RpgNJoR34WJzOYopgaIq1sZ+YgH7gLKSChepvhXB
AJhVzW6Q5txQfDjiXTng2SUiTj0T/fbKkrz7QL9robSexKtXlUyGPxIvIIyykUVH
F1TZmRRsgLB3sZRWdoKp2/IpdorVdABPHZIFL1K8ZiO/pfYBQBSLEczWRYJghfH0
0m38ufTTkkXOAte94efSaIcz1Hjpb4b/7CYt8Fxww9MxaQuqD1Thi1fotbEiEknh
O4p2vmiQ3Fjoeqy6TIYYHr2sYZ3hrX4KYCXVD0oz9F38sfTUZXJozQtcC9xGAWl9
fFkwGrnA2i/4JzDf9N+DcnC8VYpC/M7kK0D2+RHOVEDQ4hylJfJZMkgxVrEVGTet
wXiCAZZtCFLQHaK8xnhyBzmjzV8lZP84CDkU7L2Xotu2oLBGi/9covlMYp36wOLJ
v9WAtHR3bJpJH5NbBWEJHATiFDwC11WN5+9gf2D7zOzdaD/rWNZRrhsF5+w1UI87
UEIvH1A1ntMm6tLgiJp75HhjqtDWhwYosG6BzIbNGPa1v4/Ks0514Neoenp8vLRo
sIT4mksgF4vJYXvbylJWBu3P9sUYFLbD7IA3zAerUBZKKe73MlMCM+cK3yhzA4Ll
Lca8lLMZOiSa8SfrGSammiJA6wlYU7YhJYyech/pbJ/RzFYPD3qKdMn2gSY5O+av
G+yUXO7jjbB2fdlSU0Sx+zL/9rEdNLzwMtk99u2T+IgTWXFWMyvMul6GbuYYAOin
rqySUabRogTxgyJwP/63GqfQPH1sdtd7Qxe5EVK/Ra54HUXN6CB3hIdQEabigerX
8mDoemWzu8fAiBBCvE6ZiI9fzq06xeYFsXXhKujO2bSg2QxArb3Pc7sfNxulbch9
/C3w2XEW1cSogiSMSUoQ/OCoZFJQzChI5rdCDCWGtSoWvAy7WBBOrkPRXhqICv01
v8dncEpXAELjZEH2T1RlKEr+Zyj7fZLpUwb6JjW1EOgvgnEuQBC9gqWyIIK7JYiR
SndiRp6jnzaDPcgLb+EFVLUmzr4jOC6tL5jzDhE/WXzOKChjpQ5m4PQN9Am9PZPQ
dz1lRhGr45kFJeJZwr7a0c8hB1NZRVx+ehXi/pXLZSw6vuxpPmMkLmrTfGW+bHTT
bpab3a50yYr/UskvJW0Lw22DVh4iOb1etZghDIQkAUNhNldcAS+QdgZ01iPYrQEU
5dW0uxR2Tz/C6WVQddhoplm0BYnv2ogvYLb9mOCMCBOOdnTJ95/wL/tNG4UplAro
89ptk6Eavwo0MFKIrbKjV+zM3KS5zsK6yuH6hE9USLMLNo/QZjKwHaYtw8UZWv89
HmIPlZREm9/kLj18B4RU8WN5J05g9VeHpNDTuHhNmRcpjJ6TVGKwQgha5GzJq4Oz
K5fFEtNbOR4dxh2XxteqejEn55Q6o160CfWosFBbfZwQpzASanr/FsoTJM9AzpCt
ChKCeNE1YGqxVp+q6wVClGiVUd4axVD0hyD32nObauOPLD9mUOp68qkfpLlq65Nz
SndUFHB0f1XjyO/R5j6rs5edB9cj2UWWzz2Wkk9aTyMGSyYVjp7omQZdm3WASlWd
2UD1FS2J5wE2F23kyeGoVckxslnBIYwcm4R1gDbzh0AVVcpN01J5RhYPfWNygnGa
LPSlwIkjvNeRwoodzdBNQs7ZN9pZ680Epyh1QKfD1nG8WKQIx7IlhO6pLomX0EvH
dz2OcYQe/NoqA5EWhfV/Wzb/1zymxQXlDqIjMeO+w/fQ63VgHnWeDyEenTwZcH4a
JOF0C8Yeb1OBedwUe2WPxf2cy3Y8fukqytROjgFOff0GMylaOWbQHieu+zc9K3BH
YpiAVn+rQhiG35ZKaA2DTgDYNSJ2eJIAb7dlAfZA+JFCcufeRZffZZKj7BPijLuK
edZ26FxZuX3eIVxc2scMzVPWpz3HZoubqrVDmka4X5yvuyUCNIjVxdE2eSac5nEQ
OKe2M/e0yB911iYK5cjGfivcA6U2HfskLqLL/qPLTcJ89kdiMhKdWLVn2H3w8Ilw
sNXH0upRyS4zGdzlMZVncOXWuetaCA+PO2V5RKA4UGQqTO0ulUPDDY8o3JOHu4jD
jtd4d8sdd5InVnVvnfVdfC49M5yBs+yL++6sq9dRiesIKQt4D8ngmCz5qIlucbm8
ub10w6jdPtBd7bmBCWgWzdgUWsRX/WKt03eiI7tJTukYvlNB1wxkrB6VNSrTKgc8
f5ER2QmztSzgw3dLVcZF7YBi/lRz7C7iwfMk7EsiG12b6vXXWutWC8g5CdKvJJIL
GHSjU4Cc8JKNiqPAKwM/51ayYnEB7VxTUFz83qRsWu4cz8zBypvPPJykPseSrAie
dtit5hX/9xIqQZndPQkmRxbpnBBM8lEGZtVIcNSblKuN2TBj5I9yAbfjpquZiMFE
zowPg9P0kMMqvj8T1bqh10DHzLvNuawIGyoyHBCIB6CBxVx2kLUJ9dj59pH7iGz3
k8tI/Ni0Lvylm3LFrudP113DmLsO4oxXB0GH5z322GWWwYyD8upShsAd9TWPlowy
KVbJlznjgwN3x3F/+9hOmVhj/DmZ0Mc1AZ6Dmn175J5NygiQpYJZzRXYyEdaIHxi
VBp7olmfbFlzEI8hs5aHTVBjKKQwhRELWhPfBckpgOa49FCbj/SvsP2rbAI3U98c
JDzIZ22yuYI6opX9yW/FoxTBBcubttqZtbO+b4QSUZoH+noDk7PLRMXuXmyWlZaG
/hOpA9pfhhEnK5b5T/lTYCR0hfln7M4u0FT7rsMgz0t47PV7NrdlQ9MzmQRprXkx
XghkN1wNVeG0QmOwQsHBs/iQwkih/c6LEvh2Bcsew/Lw+4Mq55USorjHbWWY1/4P
ESb+r6h9D9gnNlq6jsyUcwb4MQf+XvKT/gmQMBFxQNOCmpx9OiMCb6NqfkwAQtHi
nG2NEq55WmHSuOxILI796qXX3rRXwuHVs2lYdKsxqRZOX8V1XJqsvPzW6Nl2HPV0
Gp96kigw3LyfUcRfAQMHq4IQW+Wn4bBlhF23AB3H+NyCEg190ev+FFWUD2ztBA0o
5Tag75D51pBT9FwcL6w5ootKmhRzt6UH8TC2OYZno3sirintUbX5KvAKdICQK6Oe
p5KF7IgWJo1KYCLT3aw5MdLcb9Qkfl/z6Iu1oogK0bE=
`protect END_PROTECTED
