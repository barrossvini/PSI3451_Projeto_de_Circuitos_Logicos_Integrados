`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDl45Y6mkgW+YHqqUjGH62jiVVlwZGqL1J2Rme/PMCRJFqDBgFztFCxnrs4KoaU3
EM/0+CD1jykvi14/JIYFbHNXCp7vWPaGCjGE5WdHhLh2VPxNGNow2DXN4wj8QPX9
Zw7lU/KKU/R/8vGKSDIo8bSvga2q2RzGGgbHZkj4UHuphNup73ENKOPZ7yzDOUBM
mT6c3E5dG3DUNP2/szlquk8EeBCfCM6w7Ig/4sv38GW8WepjZy1a4wF0uZ7cNH2p
0H5E3QqlqwHNxnhVfW7FKy4whf6yPepW3Ks8XCNpxah9wl0sU/ziPB+o3HPutO9Z
Fmd7wR9GqP7jTEgZltTXF61+kQ2c/fvj9FwAsoiKUpNUb5Fa9YvsavADrCG/+4e6
keB6KW+Y8XFHEZMJEGNnRjJANh2ItJVUTLFM7fF/rMYC4w93Dpq1LUFPGNk+z1O7
zVpEOuT4nGUrKh3GaYh4sMLIYxbVo+MmTyyvdYg1zRLnwwhZY8fhneZJQzGK6bqS
qDj739qS9AHoYub+VgpDgThbki7lO8m9EB84qgs+Qc0LrnqFBYNJvZO8hSiTOFKU
H3HwUpcRPZ9SxPzIYJ8uHsCKkniNTL2ANvS2e/iOe8AAM1paAArluxmgETssmpze
ZLd3MBIjMJ2s/XT1wsAEQm33y/aLP+PE1PX52PRBGUVZru6hjMoYQSZGUngY+alo
DVU2IJeIv4NeF+UphqOq6NcBmRRFjYj1Y2QLO2bB1QzVQ8RsEmj50c860f4c+ZAr
PxCf9LkTUW5aab9j/sIE7utn+Gx35sRXJVxtDB4vruvvxhCjm3+faht6Ib4QTxAB
qf/nwUa/q+L0rSiLfVEz+lYsH8CeXL5REudte89iwv2Uby2TWK2CBmV5Lmw09rWO
HaVUH3aTK7eUe7RZeeXekWw1Abarve0LTihVY+CCcNpyBJCYtkpuybFfWK6qDhJN
umgqblCJRVGCLwqDM1nZ9rzuv/NF/yd/d2myJ5ZO4DZMgOwL6MGRYuYMfwaHtE9O
5Eq26FtFcGc4owB5rCuWSaeAMNuewEGq1IufbPzLdIY89ceUWxpiiApmnYhpPREY
`protect END_PROTECTED
