`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VrCTdgOA1Ia1AHxMYThzBP34j3vTdPaFHZhMKz0nd6ukHB31/nCII/EaeMTLYE5M
MDJqx7s1LMChtxR9yPMsquEqJcVjTFJvT3vUP+TG80bxuOJ89USuOhUbMxH6d9DC
QPvOFXmrkUyNWmYOB3NaKzO7tRDC+FeL5C3WSiQfCh8BPUknRK3ZQQQkzVNKjom1
80rRecmDV63C85Aozwv/vIGV11eOhVp+6R29BknXfFgNqpwXqzcWuGdu64CcYLw7
1uYmr/Qad21oTH1DE+6okyoYGFqZixCZ08jCkoTjUY1lXMnJyr1NpGcu7G6h0Ovn
xQohvQhGUPsgyJZdjkcmBvlHkUCwH+fQz7B0kplOzkL60a7tjvYNXmvZbTW2Pyse
2iHuxbfYqm8hEG3zAf13jzhcyiWTe6dUz3wiv9MCLKXd4QwlK0Ytp74WCelZAnhc
OpIJU+zOi2/ig9lQMw1CzKH622YhWYQAeYMVj3cR8mloMGcFq0iTKXOSewnvsBZw
sJtsUVvg5j+B3meAWHt7kCQZtbI8IKU9OWOT3cJ//relOe+ucwptryzWbkYva37W
rvRsrF4hp4cF1uX/G9Vl/w2uGouJ22Gxads2gE3PfS6VMUD4SxXqzQCHAmpQDUJc
IFSieEr8WorDPHCfclXLfWEdbvq51BRVsEXLo2Rk/DnGAya6CeYNOIHsRuTUnvp7
g1e6akNsh4gmWr/HUh+yq1wHG9qU623Nvjj3jS9GAYZnPaT/LQVHqY091OfZSg+9
y0IVcWvHhdMPgkXU74Lf9R2vb8UzXr/DNcwGmpUoV9nR4r8eRETI9/tOdBH4Uc5b
DuHfgXmF9sX+djN6xg4rhV7qImU+PVutrGkFDFDo+YjlxBC7vxZhsagNHTGRaBZ5
M1ShvDkCxQuJqnrcf5sPukaNbhFza4Pyfn1I2ZtidR36DgpYThgCldGaEGzuWCsj
1iFvJer9IXd/RsrAi1cfMo1YbvP6hu+4k8iid1EZeTPhkKVNoShd4DLOt8RtjYAm
+8UkoSSXTTwJEIFveEkvqg==
`protect END_PROTECTED
