`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VhBNYHIu0BIXl9eIcSOk9YYH2N8yEW1krryk3IpIcv9InNbWKzT+fr9WkAvyue5W
nMRY4N9Fj3pYuxtqvYPMeKsO9gIxLTOznIb5fWkUjYYidRipuhW6P1jgBhM6Y3Ny
9i0414wVJF47rvEEOpArrlN1/qVeNH65IRozFaXQUWdZya8ob1LbovMiocjLUqRx
N6LAIpTjUbtR4dFAzVr5NqzY2GL9sOVS07JZpij0I4J5F/cmJWiuSEzUstqpgK4r
gId8/pDCQP5yXUDfBn4I2+QVSFvoYpMbnuQLWdwCYTLkb8TOIis96DI5xSAkJhyz
jdDcyTWdCMt4/9+2Y6jeJQVHlTYTpHFEA03TQa83wq6U6nwIjeXDC0mjV6I3MdOT
i7GRSq5TKs2NPU6miZ9KWIxUhOJXOtXdI3xFyAegmu+Z/UG9+sHFNDblpbmm40UJ
kLBMQeJ8/HlQrdoGJX9ZXtTtBaExg8u/y8HvewejhzgwIusdQHczO8KBOLn+nQci
xnZ7BOeYx5XIhfpsIEX639HKxfMKrX6lZ4W5wPgy4+tAZtXTM8ZMtnAn0cibymcg
6hLyRtS+iOo0ygTpZwNrufoddno1B5xQQl7qR6dtjMFV9t2Cx6JC5ulOguY0ocjO
jRyYxkhF+v0L/9dwgrVpsVXQyc6I5feY62ZlVkVdffdGA1lITQRrw6NZ6gZBj0PQ
Gx95beOQnp34ECjGmeQq58oLdmYmOjCrvm7MPjrx7QihTSVl+aNog5H3sWjNcTet
47Uqy7U9xmcCgsTWmRyBn94GivVelEPcczS3HY7dilphk/WipKLeRB3Pd35OudL/
jPA57PhQjswnPK1wX5Jy8g==
`protect END_PROTECTED
