`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
njaWuMq1Lrrj4Hun6Yh23VPLQWP1pr5K14QUBIW4Tm59kBJTlPiWoDbicBdhB4ET
c0DOkA30wHcCDJGfIw8ciMZtrDdlInVqDrffno/F3Spyu8GLi7rjmj05OJ1qNAX+
UIXLHz/TH37MnayaAKK6L37ZKB2LdiqQd8AZVKR8npWRcMTzFFw+3qssVl+wGknL
wxKxwU9Emb8ASVSmSiJ11l3Gkmi+0Xy2YfaMnpE/zywwXqwdK4cciWztR3p/APby
migGlQveg7lL1mVdbzaqDy0GDRwgCJ0BhFAva3xeDTye1bb8+2P/EMVLr+7Uok53
aYU2kXiU6Kh64KA4hfiUQ3qhk36PyFfKW6qp7MAonF/Gh2ItqATzyKIqGVypayPC
+yWsppyzBsrshEhMtubWZqXQYkKrxIYCrifQehZ3eZNVgclQ/U8yeQGssTgOSfOd
0hTSJMXVN5jO0zABRrmG6eJFJH1uMfKADhrvoH0LWtGRSTf5mqrLTOcPp6DcY3aP
bbiBDq/Xe+LnVlWTC04CUARpTqko2tGK/R8L6N421tpmyevDEh5+seC6nM6RoKaG
lHI8L1OUAEOvuEO7m+Q1b/pNRtzSLCwJWtiJ5mgN0Gy0H6XA0+JlqwaE55w8+iCX
4LOkxXOJoYl6Hsauu8oSh88AVqjcUvho1+RCpxoMA54KrtKFT/R+7G1J/vtEZ6nC
tJflxMKM7+ATmcDyN6rSqnD3YbduDNSbHlFx5RdtHYdzXGcaSPAuGuZG4594nF4h
lJoviYEZyh2b5FMyLOXxYXpPU4rUhD5RLbsD325XXRWTGuNFJn3dvIgPDPDVXpuO
qUQPNXQTEH1aTVq6SIiB8Q82jdIS67xrsgqclePmSa2XBEPOA7TCbjw4f1J7fHNK
w7cpLjWStG1zqlySk3S6luob2dILDwni7h6PLByxHfP7VQaz+69FLeQ5PoRycQCk
WYJDt59TvaCovLhhIU1B7xYSeY0ZRroQP/EW2VW3J9up9yjAJKvubkIaxnTaKyOo
ulVOQVsMKVxeGqWIt+OofzeJtOft7KZMDZYv1bGl/YmMSXIlBBjO5CwFo9AJYhWz
QvGnxSwTGI8hbevic9W/zbeWKMpd9Xv/bHXYRkeztVJGqq9V2tm/NYtZiNrGpi7t
dIQDlDIAfKTimu/FxM6+9o851gcl/zqYcNs32TOghnjzjjk1F2PvV6XaEz72QVD9
X853A/RwgMUZ/q5uolNwpdJ5kB2i6qEYoPcJRxDwcm0GhadS3nkywnLD/m28B2M+
sOGz64TnVMcCQ3nbv5hWzO2zQiA3FmI9PaXloel+d4YbnRZo/E0flf43GIu4Xd4c
lj31CtnrWbqlx5jEbkj1aAFJtU2lQdqtyO+Ur8pCarL/ixF1TJG/a5K/RVG+tlYH
0Nx2g6gRVcAHBQgrYqrYR5vBMTq//VR4KoJVHJauG5rR7179UH73uDTbnRcKRg8u
zAKn7EqRDVIWFdgtaFc4dvISqW3T1IFUTSF57InZHlZjmSPlfTdVoljglD/HkT6B
4FXsculFa+ONGskei08F8WnK4jvjsWcWMguM/MCOJ04OM5/n7vtm+7OgCfbP244Y
7DxWrccX+oC2m8YLHIKztVlpio6FA65pNxEafkCUjv5c1gn7sqJUuUGPc8OaQ9VB
r8YY5zKsmqmdISHCUevUsbe/fgNwA1dDuVPtpXA6kboGYMANvD1hlBD9MVsFNUzV
Qw18KoXQtFNmIagPtt90FPPXfCwbR5WdUEs+W4I8BzFVFWwCmEjs9CAriHo822jK
65kuAIE2he68fiyuA+FN5EpnAGSMQXvNYBh++LKc2w5o+0GYmCzQpZZ9j3vV/+ih
6Dvnfu5lNygIKYQm1wHaCi4FCo3nr1ohwfTGKk+KnlAzoF0U5cGt5EUyUPDhecv/
yAteK7cECUPR6WPASbSVb40umZS2Hi8infb7S32LQhvFZw2fnbQL3MEnOpJUq7j3
e+IpYAn3hfdpcnxo9Sb4fI/cmmwDKvTPvAfRZx64eSGTd1vJ5cvGlSVRgcD/PUnq
eVKDMrzRLkPt7GyOc6Jfa6Y4KJZlFAmnjDVLTAIqH88w6PM4cavdW0r6MTJ0mNSj
CX8Dq0JbbRpLX83u5CE745kUz1A4sY/goabBJp6dy/6oz9RpY3fYgoK9A9DFyufE
OSJ6SHyLx6/WOTZJ9gHtMp80h3HTIIRe/4IQcdnHXCTX+e9USg79gboBhTgLFI2G
VkMiR1xe4vrgIuxkeXjvxFmkfhpJH8LCIDC2kq9cXkiK7Ku/hM5LdL8LC4i+59PZ
MY7Q4iXq/Es2RKUfgPLkyG2rDMX3N1A+WiVZt3K0CWJhnf3rgH4b+hCvQe+oPaMO
jYkrccYzwFEnU71vlk9ftJSwcAL3TOeKy4flDjz+SWvnF6aHFR//ujLgeMeKWJKT
9S8crEk9DMtB2TTTGxiq81S1G45BIIyRazYHNaVTD2e0jCmT+sYiz1BMgk3eE46M
ZZco3s5LY0rWxMOI2ZYze01eo8Mj9DBp3xkuYhroUuMUp7tndZqOgSP9WTJfeqez
IuzPXH6yf5ElUsPvrN01ZroXCuu0IKcBqte1yrQMpmY7lO8lYnPYHmzRnbdA3q9U
Iy6f6dg2aXUC8MOs06Pc0XdUDfAjHbY1Pu5fvTh6DIqVaQiriL7H130H14kcbu17
Ath6Uy0CcUEKU/Eyifuz++7ZDfRMsfgRdh3S+AfzA75PxKOQg7rNToGLP/0c4jpR
RmxG7cUX1nFbo3lEanFfGC+Nndgrx5Jx/mn5TpIwenBj53Mcib67bhcwW1Rb8Etu
ZHAWYsRUoj/YAhp4Rsd6piWqe1SS5of57GBvpcRne49iAD8AR/mPG+6TKhCaUMas
uekl4EUUoxEN1uGmjdhnaSdCPPsYzRTi/Q/JLczfHPSnxmbOxPd6qQYK9pXVH9SG
IK48mti1+SZNuDJtQ1SR/wqTw7tY19On/M43grD/vWEh/ncVw2nI2+E+5Yoo/1EU
f9AaiIOzIHWqyfcweZPow+Qk8mmwtPo6v9tjL0PUmtfQd+EnxjYb+WYBWbRvOAc5
fCRv1MqMxy+C2cXTxauYpjnVxGpU9zzcv+8gMCxbiSXe55WKTusE6RluvRQjtcLa
KW0+eXuCwgA9uN+z/mu5fSCO/NzgHz1ZH/7jTDBM0utbJnjoEl/Vt5+PvXFdM8g+
ZIWjKEzNny8f5IDNRtve4SixeV7itDM4BelcBoHLV73cB/4NPfy1/5D5F5mxX9mp
L1gPCjHlcYOH5g8HPnU845j2JSsezL87VZ3uZea0QcNopJ+8609bfST9YqM1oGlP
6rTmzDSV8kwCKqWyvkKxZG7wlPVn5zQz2SqYup/sHHVmmNcIp2Is/eIAC2SCI8Jv
uq6xA0ZhIjhZZ+2/SsiYh9xZvB/hMOd3HSiXpfayKkDxHs0zjylCEk66eenKSnG+
Et5lvpf5C5/RphvLaiHKbATrUlFgyyXGLQ+Y2DDxY6X8qyOH6CkGIK2Q8Fj5AJlZ
gpC2UskMILlZc6GmxEjGmqp6wodAYngcCMmKGNmkcgzZ7XFdqjP2TcLpdwVz1jIX
7uXCDduAmgLJdMlp6efJ31f5lnK1afQ6uSPJ0sGMDAx7iNt/Y4GahymwM01BEJBQ
ipWiM9+TOLT83z9yRkzfUVmmOqdwANIcP+6ERNsAC59nF4rAEyEsJ+alpDdgNCWi
CW8f5ZP8uCpSQMoxyiE9jRAvCkQWgcBNsxMwrsVM23HYyN6z46ajug5FZGmnntDA
+ID3E37Ui9y2d0nYIV2SPlS3YEVo2mC8z6flnLvqquZfMF3l5DejlXj/0O/lCEU7
yeC6sqJ6e+u5l/UXERhR5UeH+8w9m6BlWqhcEvnt5imst8YgG7XnZfroOyQS64Oo
zQYSf0lVNeftk1mmfojYAFMJ9YFmlfzzfMWvNnAh7QYmEQi5Gc7HQc3woK/llTKi
2UHG3ClWtTaCc64JMso5PWgbiMZyqLbAMXfXA6FzAUEstvqIdQK7u4D7uWWc7zyJ
GJQhpjMaLJ/+SL3lcuNVkziAKw5t4sCu6ZOF4r13DSL4P2rh14ZYKHjC9nDRl86p
yC3GCqPUqbCj8h6TCZ5Gmnqo4CLWEE9Yih9XMNFEvGCJo+evB7pkIO9fSy57GLzS
CEDh0rb/bKGf++06Ow5M+936aQEkSoTPfbSnnQkoY9BVkN4D64srpZM2+Oc0saeE
XUA4JPconqCKSs7fLziEOoa8YyRGRc1xbHVCn0uoQ+5So63iqDrAr2mJGtKkxUlF
w+s8J//KRPLDRnKkTcTXrul3w+e/MB7YMXdAFEb0cYjIPGuiG1048Ehq+WpEG1lG
y5+LMsTKWUikdW6zWGBwzBe6C2A1c7XtfQKLJwzphCf29aBm7Jur6tzdzODNXlUJ
wKKP5U8PXyVVap7aqhMKrCpWccPh9d/88Y5k3IEil11Ujq/F3uL9M99opBpvZJaY
SsJlzuEonf6/Xm5JWgsmAegHw6DSiWiNhOpzbQqY9iTCFcDcvRfWB+3BaaBgtGkR
+i7KZTNQPEItmipMiB4XX9/b/sw5pHbOnZ2KlcbpisCiN81A9T4TRnC0seFZPE2o
p6zjq1hJWAAZw0gK9aEUPSKr8wIIO51DeOKvxv8oLMpKOSD/iB592ObyQA9RYNQn
PYJV14x6TytSYIhRbzfHYJOcd3ptPBtjyCnucmVTnBuSNkBNg0tYflHh5GFoPk7/
hou7Z3S8vH+hBcymBtkdMiw8ISJy61SfA72tAgqIwbu0eXlTmj0V9lOiznSiBpIp
RWGICFpxJ4vHh5I1gdtsiSdXOqjASXKrYGCO1y6VNQ5Rzv2pTgMze8SdKekHE8uT
/zewyAIQvZI6cDYrwbkEdj3nydbQUMfkYMmxP7LV2QKUoFWPDPb1r2IQF3G0gdId
NosnAkYR0DhzAnL8djHrDLvgNMB+COCqYb+0zi/skDK6ndah1W/e2Id/Td7r7w5u
y3aJZSaedkQArsgQVo+lQUzbm997xuK6RN7IDuQGhg87OIgGFTirjxPcg05d+rOB
rPepUOS1IzHdnRR+L3uGYE+2n13KpYgbFqln1Z6aASkeiHwIDJflkUyo7o6RfFee
ncTjXcM+EbU+cmMw8VRadiF7znkf+TpscBKKEnP1vJ6AFS/j9dTERQUL2O1qas4Y
kC4RJrBV7I0mSBlV3VOugXW4xqMHBJ5Hii5vxuBz4Yzvswvaz3puw5H2elt9Gf7f
IlA/Dw8yQsXWx2cYzi+zJv2UonVyc8p3wPskojbstAjq/oAGcWwDadX4vktM7L65
J+osk/4deZ2aTFInFacDVDRiWFBq8+JkCNebsM2w7hjpmL0XB5gQnsQgZK1soF0v
vHxYOvEpS8Yrgt8vJfT36ybOtJWwtW98O39sjzSeqHVX3dG8muR0bUu+ohT8bv93
4AkAxSDC9g7hWe86kG+zdpDS9a4vgjMBkLqlr0meU55CGYZSezqFMG1G0uNlRoZv
jDFVihggjV45F9fLNM6vTxWt9ACfSjx4NlXY6MBBuwh/5rD6sENzE/xWBQmGtnYz
/3IIdZE+eYm3CQbVBacX3TZchx3HSxwsjEhSycJzUyWZUSSZYTVZGUAql9Yp8eBU
KRPm6EM16cy/+x//3nDMwKvaCfgnLY93RRU8C0HZKnkMX6YmEzFgrMlbX9ys9dtL
SJq8ePKgtzSwMO+r8QeQP3mHqXoMDsxXp8D4FAxgDyM5EZNM98HDaOpUeO5hHvXa
OyN2fljlIh1RrcezrrtIU9KcR6g76tn2mZT/QstDskfIGDk/tlPK8wdDzUNqtL2Q
KSs7/pYXf1FQr5IpV3fEJ6s3n9TKFbKc5w4BMvBjdICDEiyhG3ftNvNNjZ25Qwgx
ugr+UUp6ePxkL/aYZsU6QneEv2J4wZGd86ghl+Sm/qmT6hbWlaRFdrOGspCBE7/0
WzjREdwry3F071atFMoLTa0JAMv0DiP0yTG4onli415QqI+e9mkSyYWkfgRirQw/
vpa4Yxm4xw4FObvgM8MBLjBg0B7I8D/GU7RP8vJ/toEgN4ZT9TOHG1en29ju6+kb
ubQwN27ckNxzXXZat7cW88zjNLUIleMUZ7PHjhLQB0tOaorvXF9BmBfHPt2mMcwd
z6NU8q9STnZ2+OaWsXDYgcSbl/ETS0aoRkk/WZtB7v4SAncZg5aENQFVKZgI1hhH
bQUYHZEf6ucZlJviZn/sUdFD3LEH73vtI+plYlPQMuNmgYpWgBKhBQCjTePxa31q
VjNs9UklkuiEJdeH5K432Tn28LgK3TPbBnvKzCGKDDkkJujyO6zDZopE2AjBzLcc
MSx7RlI0emM8lwsjniQQEMMKVQjwXljfYDMtuLKiZpAZW03NsELL0KX963rxVERG
0r4bFNlM/3o65i8Wwo600PGBtmW8o7xHJgi1lR78vU3Nmt5usjCUGAV49jOR4jQB
aZc5b22q4761AmlUKsu6sVWfxhoJfCalv7mTJyq7z6dQRpHObyVCQDhBW6/N05KT
VSKR5j7B7n/DEfQQrRDPMOGKKnL4E/eQWvqdwZEGyV5NmjNbR03sJXbSeeVL5Tjj
7vbA8IbzccPolSuMeWsIXo4WssKzM+i35aonYLcF3RqdjtCHiFNiG55T2wkJ/WoA
IWDpIiNGk+Wup80PNGr6qupJJUF4evDX7Z7cMCbsuvmNizynqaquHnBRNOWNPxHY
l1s7dMT3ho6nT3y9HuPh4Z7YxIdV1VP1Q8RXzRu9E0w=
`protect END_PROTECTED
