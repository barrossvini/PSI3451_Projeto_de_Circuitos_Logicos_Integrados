`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7dw+FrqASjiL1Ww4LnxoENyCKpPCYEENW562by4dxDMS53+Cvc9KzNFRUlCes2UD
pWPLnV0xJoY6lbVDwemnr+rZFi+rQz6XmOXRhq19O/0hr9usxx144iaDMN86fzQ2
KsV8A/iM8P07t6M/PO1j+Bi+TgJ+yhcrXeUhtkk/frRdl+L9pBYPAKyVOXHgpz3v
tphALcpz4UjJunhO3InGN58AktJPzN2S0XYS9gBZGdAMGonbV7WNdJKH1VlJNcAz
bXMG1ynr94XnOkd4kZ8y+YXyKYSxC80xCcAAlS+gk7/nkif7FlN8KUtekNmNqbv5
vQ0GeQrRITFwi3jOm0AFl+uWcZgw2WyNirn935coa/XQwrRqKjTguP2vbGFMtl6x
EetaG7j8XW7Mvefze0nKQ/KQKi1+DdBZRNH8dzOqSkUV0HpbiKj9omGu0dOgblnc
8pog3ivG3kAVbsrHfIQq0vdeArl+PGmLvg6Ofx7Q6G+/jYdYqjwUnShqMvm4jcRv
2VzroCeiqVZzQbEZh0W/Tu9qyzH5sFOwMh0sD6v9WLgfhEvOa4HY6qsMvfbJfBXN
bDZrxfk1siNvr2d+zXj+4xnZPhHPfzAEX4FZbTVnDIJXTuC0FevAsUCCcJbXQzWu
f0lpRqJgtMewMHfmU2xELtVSJTfztGA1RrU4jMT1n//iCdZiWx+6NYfhNNEcfx3+
pq04pXIXWq47t0Y6t8XC0IyqKXAF/XfuU1uGVUMazDV3VUJGQPoWI79Sx2iTqBYL
fStvS2CB/4zL6FG41GiUz+i6aL/s5cWTNMn7mqBb9pD4rFL/amlSA01Bsz/N6MI4
6Qyx2sMTGw16vyq/lyM6t4IGED64hvaRyXsHaRAbZldVwJNflHMkvzIlAGG6mC5E
0EOO12hifjkO/XznZZnojsdHMcIR81KKo3O/mMIykmYlkB2vvLkLGzzHO7ApHOP0
`protect END_PROTECTED
