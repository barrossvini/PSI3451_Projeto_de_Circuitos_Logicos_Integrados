`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wuRagJfiJarueq8Gexn2eOtz6rJjeoPk1iPamCLeApWsbCXtNLibcXG8v7VN94Yj
FUImJ1VlFN6vQ5aW0AzUd2/i5g2OfmRzPRKoAOteOCLOukps7zJFqZfN7gy1LfLl
MlDQEoqb3bkDUtUCdSBwAsm0GQcD4XjGZFZE+jpEG0mlP0fXnG/o5l6O6owoikAc
viI/ShhWC0mU3CRq7SYiC7CaqGKU3CZ3hLroG36+gF66b0ESa9FVFtF8qmq81pI7
f4JSApSvIj5XuajtJ0c6KNTUsvP1elBM2sEDumWW8P02LFGz/PTp65N7hiSux/+C
1NJgp4ebd4rwA9uZHUhn3WXKRGEL8EPkDzLsHrw5Cl3Mfa08JnBZsIYMmTyL1/rp
l2f4gP57U2m10VXsmYCdC1u35Zv6wwk3JfIgDRJfLWBdHgqO1wMDrRZblBFiHN32
yAbRni7urEwLyUDzO/esuI2m19cytmb/vclXxQYQynyu6j9WK+tsjEmE2Z12G9km
zZrB2cSwMtwEim5de9s5a9rzep/47mNxp/nY0WyYcXFY2r57F21r8u7V6kaBgQKA
YbZRsgPLIXsUjCNXhWw4jh8uaL+YOzRgFNfmeEPgZkTuFa/lTw6tg+hrPiPm5neL
Yy/LoqtuAyLXR/TWFSeCOdhmOsEZtEeMxrQS/2JgQTf9Vgo6M/wMUq/ybtzrWeRl
BViNa8ALKuLP/ODVpmAttgwUNVU9LzHBDrZZXj6eVDVJ/eWvVmJA9wzNIkwe+VOi
XKMiQkJnp9pIs9c6y2pulN7thflnmxOcw+3CHeNo8g0JMF8OYcur+VJp/ZL8lkIj
pV/Vd632rYkjc8emxA8qLYgM564j7XjLfLAB4EGQrxoiXmMWu9VjQAKi2k0JtBje
xheSx2zTloSz7Be9dAMeiCUWRSsTJaYhFSAlyZiDlG4Ff0xBPUP/KRdQNU051pZQ
dyHxcLIveJp/xG1VsYPb9r7tJ6PSLhqV4ENzRkvLGC+rG3jxclApfzDG8FwFy1/x
zvDc4HrG9CXovRaJ6/4DTY4B9iA/R6IpHzXzX7yQFD8IYjU/8C89/N0o8zAi0WpS
cx86O+5L1my4k4LFifzSU851Ps49qp/uiGFSqWIPXzh158kKxKFsPmwlAPiL5kut
ORHCLXuy3R/KRnhjEvcR0on4gPlsMKeWTXkY2IdF1h3tNaGHik0qWqdNWcti4V8J
fl3rb9ZRhEBQuO5VCY7lqQ==
`protect END_PROTECTED
