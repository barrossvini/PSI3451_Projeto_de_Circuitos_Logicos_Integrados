`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VuUouz7QOcZo8llDKwI0jIn+nXQ539oHorACx86OhVeU17Seq2MXlPrnnML2WhRF
8U/kZR25rJTmvaPXnt5MPvqnzXQvMEEehqp+/VbyI2l53bhgqVGrLzwEjVL0G7IQ
Ecpma8Wwl+7ZRz6TTFih4pU18JBvaMs31vP9AaMvOGwZw8PL4zx09X9jWQNTqnDt
pwLtyk12516NO6NruVd5SFjcA8e9X+w6Rc4MU/Fi2qgG2HzLKye9bqqPkali3VFC
bi6UBrkBqHc0zb4OAApYBVknDATZgnsJNdPAcHq7tZjV87oCwIZvo4uRl+zDOnbM
nUZXw7NQmQd8C3QjjgofnIAThGTEoKo64tABLXnHAzaALIHR9vOd3YQPWTTh6vMQ
UMHgEHxXapvH7qGpxjSxPylrDjUO8s8gb3+I4Ml/qPoSp4LKEOY1VG0EpoqJZpH6
AbklkESR+Yf+RQb7+5svnQdaPihzGZaOUP5s5JbCdVUKJlluqODrVsDTuAnXm0gh
rKlZ2q6NV6f/KLpTyhaNikiEP3QJfWacetpJwX4ZPvfJNQn1J3BfRj0Yk6kdL+kF
B5KRCvVcT884oJdZwFhBmfy7KC85nuODE8Rs3Rg5EXUx1w0SaTDepfSf6n+KRF4w
apc0sQsysD54gwfYeQkifoiL2b2yVE/EVQZYaBXH7/ho169nEgyAliI0B5U2RMuB
7AIkM4103Y2NDIW7rT4s7nzimuoII1h9/gqALE1SM/vgKgDQFflsAd72ZDPCjV/H
QbFDkz8ksO08g1tgiWKvtxq26WAnuv8kmeK9kYMhPgjOf88FuQboUVgZez2F2wFs
mCSt132lxHrA0TdfFa8wwHkFlDlOMD/7lIs0bnBG4+lvDh7+b+ypOseoNl5uTe1L
jk4Gw6z19KAjy3CIVCw8UXx+8ShGDsD1vsNfkKQxpHxNKFI3wNSVjN3Z8Pf7ra/q
54C1Af5hkq/YSQ9znrIb/QJJKxH6zMXvvgck9veQtdCX47KXgf7Z9pK6UUQOtRhl
d9uP/sXzFLQXC97p4tUyV24NYzVH6n0NCt8aP2sjsQ1zAKrEGELVluvdovgvrW+v
kDYydyGyvtuv36FNeNY9akzCRcsFQFsOoeUQQmxJGTpSctjCh1ttXSsDlYe2PF2A
m5B3uVuGtYrnfpiLU+QCy2J+IiAflqOFFSgaof0rZ97Qny5lmHrcczzz4mTmtWKP
5NBo40ewpS8mUREkK0hfk9QB5GZZZROFqfZaPInl/zlLwd/GH5iSe6LzIg7E5iJ7
JTVy2Ylvp8tb7HQCLvQDmH3XzB6x53Nws9Tv82bN7KxtixVoESOicBlGioc6sH87
3PHLpuXjJiyTR2vWIvdmJRgeoEY2/z6fEt96kTX7e5iAyKcYz5BbAwK9WQKj3SjX
1Qc50UEidjakVrHvYiETTqA6McUsBBS0vsNvudrWz+MWBKeqNOg20/Bs9hJ+m5cB
Kwtc/xkENZq+Y9Oa+tkTGhuXWRoS4BaPg86x1oUVyesTSUvxBQjA4P/JfmLWtGn7
0oqlO2n/XsQf+lTtRDdUInjCJx6mN4vxFMbNgY71bMpAwwCOXZHtwY+/KvHdZHh1
0ktBm+gUHVdfdGRojutFIf/IXEPzq0vlejTR51tc1jKWwJt7/b3KmV3o0H2lJ0xX
t+8FPQQeemLGF2VG+mMJJ6pVo2iR6rQgV4EkF7cNKFy07K7TosMVdMRAcvuMdESS
fZz2dsX/2hIdtNiqY+QScw==
`protect END_PROTECTED
