`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KCF3srI1uYWLQdaPg8rFKbC2Eq9ClI0Uk7+p3MQHf7m6UOro2lFTwKzeder4qpQk
T/ZG+lBUdO1dKo0DQvl3OYThka0Wil0i3Ay/A8SPwAkaZ2QCGkYzUREb7KNsoISQ
9btev4yetoC5HfDcaV9gmoi/w0kQhXF/NhmFRf27uQ8IJmKq8/pjge+LOlGo1HW5
8klq/qOcRnOuW+x85YDUPBZ+M703zbvOrGAS1KUTh7uMVY/Cis9eIvsATqaJHKBG
4EMz1HPEm9d9mf4G2mluNJR1vMtIm0NgyIKRaPhitje+pV3LWBpkihqxJT6O1E2R
bEyi4IPaJxVJ5rR93J3uuN5VmwahQGYRFJHP9rK2H18HpjlKIOK1ibV5yxUxE9aF
FA4SnVWYuw9NTAcN4hjYsylQDiEPEyO+9eEj+dJnMP6S6H8IVLNL5sSLmwKCiTwI
iTq3zptleIwvyC660xj+bVAXJ0XQId9GhqfX4eWSjMR1yYWgHJbjxX7m+cLqPbSI
TWHy/NLLkyINw18zHNUOyARyNZWGK2lAM6A59B3bfd2jCYw1DwuOmB/EtOKDQb0P
WcMLTvJHrsED/KhGfkVxjPDoRxGtNLSlaWcKWYn5pLOs/CuT1lXaSzRs3kj+E791
UFVYh1UFZ0uMkfovR1tKbhz7evzmwkhkKseuZHMvoO8TxzBskO97HAuVAJRHCmgq
hzw0co97A0/3YGd+H+IqvoFRroyREvYmq7ilT0TkYxitgzzf4M816aopiSWnURUm
SviTLnprvto4zXF8rsQp1sRKlzBuyxR/tkeyYMv7AWGx8whT988pBRiEHNLXJBq5
NGA9DyJutmgu5wepS9vrdqjP6Qkw5T33WrnWepY7uy9Swz5Jp7zjoH9Z4orydhJ+
LSo2VWkApSyLlWgIAlDrAaLlLKwJe0oOuWHKRAxaMEYjyYmaH6eanuNXjKmouPnn
2fteq9kbItsOijvPyCEvTNLPfG/bstBIovwX6uraPkf2Dsr3cMEzaEko1QwfrJJa
F9aCaRuSCaTaJqv6hS2iT8ODty/jtR/kF4ZV/Z8xl8z/5rKO7THBGF+XPfJOheer
vRj9W0/5wC7eeF0H6z/b7jZNnp+4NR2lJSfjgKldbGvETdBxG0/kmzvTdkIr39p1
aPE3W93UHfw27Tnt8wih45eIuUgZP4iGRRgeTxgo+vZkD34rGANqsYWKxawvFS6y
GOFU5H1MGcIqebI9bwQdpfZh1bc6bFnUxlWoAigGtSsvu3+A1scjVPwX5vM4WqMK
OwCf4Zr2Jw48awzLZYnmzJ39JmZ0UYT8cKU98dMrdApLjk/EfcUgGO4PlPA2gJCY
Q1AJnpiLnSItCvEXwLKUaFo24EQKm1csPrr0AQUnXhFEql6jvvXlmUz9vVKn1Gta
CKJ4oYLAo2V/NFunJRhdyIqRf/5l9kqJ9ankPvZk/Iku02bsS+BPl7dve2INRUou
h9Pp5MJYGPMLwVH7YlawCqiPMe6kXHDCSWLty003c4FVZX/vhwS6BcV6xF+UysZJ
K1Hbm/Vpq82Yq2Um1Do4yQKRaKQLf2PNdJ6G2nnTwOOIRuInmfF0nPJtdRVNM38m
NUlPxNtYxiKxz812EKbwIvYwlv4fx/ygERKa3sDlAxLb3ualk91AugOj2yBL3iiD
8wsA4PdMg0G1/xBkbH1/tfQ+t4C+4Pk7FvkkpVcaGKcc4ls9pKp4dh0k9M6q9XBP
gjL+6q2ngA83WuXD83KpJY2CfF4Y6kp/+ZoEsBTWYMvD3/B8u4jm83tXvMS07GhX
YRKJTWuZUcSOK/stErXbNk1iH7cI9R18g0KENkKV3u6jnyrBP0kAdxsJrWiDFHQB
zOPs6u6Emf1viMVjlevtGLF65eYu6bA1r8aSp/RLe4k8QY9KVhcI1eqbp9St7Kqs
qwBQLFOBhh6K1jFiwq/PPjIYRYFJR6CrEUQxIcwAwaY8s0y5XhnlztofJmcTSYcg
EJMChTVWNJ3B4peFNWbWEVCbysq1Xg39eyiTiMUDxQCE9nc7cRGjasgdHOrMXXLz
TIe4O7fMAZWhRWmUsA4oRumyD3sDYDmG922LbBcsX1MRNOBLxqT87rj5IgPWb9CI
TS2KDgXn1niSEOnaZW3je9q1G0LOOULeHrHOZFvmJbmY1dRO0Uy/VBWJwObr+ESX
QMpk6mG2MmptgB13U4WnGf0AlKxuwq91ro5ZYClMrX43WiggR4hK1qObiZ1J+FdZ
i7ow/xYNSLNmV8IMigabc/EvNYO4IOXkggYd7a93xeLomMHKdPvUs9kz/5Yq0y5A
jYPY4onXmsjUHjT8HZ+x2jEqv2aRFv0/66R2WyLugyZsZK56Y/fQTkYV4JV/n+/Y
s7oBSX+ztj4EFtWZhrzJVgDIgVnSzEr9kUOY3WtAEf5C4zzLxlewFJDUCtxy+PqN
HC8TK+Xkxs95v5Pi/W0R81+ZkGtTtEQESY2DLhHgYdYlV39JzfAi1jvucTUJy/LH
rnQUwUukdL0Gdj1jGWMScBFmsqNGOpJzbB8q6LxMoySb5phBlv7FRvzS3kUrD+c/
aw6JQrBUb6A+EhBtdWpbj9412SlQR8KA2iHEDTkLGO1smu+WNu2En/wN3y1B6J2q
r6U2al81uXjSxRmGu6wC9ei0SRrrueXdkKdEbqNvqQUEIMU9zXmwRIjbzqSMc8tt
xXWnsmT45PoAbAf/rnOsafhqUcM35lRLFNmsSTIMJZrI/rVuGKp3aAh8slnyDQUU
LOLGynJasPwlSErkRNum210+izq2JSrCBzdX8f1UzjRV9E2UB/IC86i+wzwbTyWR
9mNb48bYIBNuxXK+oePC27irrJuKuGw/IeuNY2fSVb38rbFBLf83oxSfqrFtW0Ik
9E12T/X9eDqdw32gA13KYPCSt6pc+1au7tb+sfK0vecyx2QMSSALoHPd5cygI8mZ
OFitMe/Qx6KE4kvDWfb9LtL0y/Un+9TxhNKo1+qIdLVWHdLHb4qT1ZYCioBCOTE9
p+fgWnNhRDt+9idvvnUAgB8HGkzodGunSeQml1XOBvKzxFgKdgFsbGGrggvpR0GD
WnVGc5lFsKvKq6Y9mYB8VOPY6MxOd4uYeIllX6kVoApL8NADO94yoJVhEJwdvMFv
oTkr+dnidiWeIwP0PLVqamgXE6oxPvmjamuuGQQkbTM7uVXkrZWYhUhM0Wpc+DM5
yzrVlzZ/aLl47sxGcTSFMMb6x+uekt1xxQri0Z6ePcexi5l2IzawtVNynJQd+ybP
PWB7DpO2usScps3uNDGRlPSKyq4xZa5hVtyctdXns8Q/uX4STYmf9P1u5Mw8SX46
1fP6EgqvzuP9YBMD1C0n2g==
`protect END_PROTECTED
