`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33xqx5mZdML+OmmY76Ylwz5SYjXqPG/n8+VBpSuFkblEy/NOpMA/uFgc4ncrqhAG
lFp2uevsFk4DtGsFOGGgVGMQEu4TVxzYaAQZDgs6w1+1gMWT6/OGyvQqkxZnf/MO
XEnEA4JK/WxGDt2lIRBbcySH5w2tV9XTgSDMgbZTy367qnwlmaM80bL+LIac420B
HozxuSBwhDKKI7JDvt/bpGIn5uL10Ij1W9EgLOZCzWVIAmmQaAxFRR4M6IC/P5uf
EhYrWBk6j/OMLKWzu7TXeR9H4NlK9tDtmmwIp/V9x6nkNeFNh7RBwSWWyjKT4MwW
oOY0tepfVfA7h/atyb2E/4UDgiFWNj5nbQbCY1JiaQZZkMORs/MHaO6iob+JX0hq
ah5F07VWOSrPXck03Csp9EmWnGLbp/iNAwNQHNxthzZITs6qk9YK9vuCGW5k3q9V
y5UXh7ie1Nf76gUQl7YgmlGAyzj2O7r1PZiLqb2HiaiB1O+jbLOgQhQYoJhWooKW
SZ7N8rVrVKXuCYy1Pay4qQKBo7O0/tpUiRTbofcji+CxXagrVPNR8ev9Ffert26D
emsuKKUDab9vlELaGP7CjiLWQI3+W69mF/72xixfx442eSVdzuRcbLxaJPc7zUkP
DiLzgEM5biK0HDCVy5mIC/YLtnMBb8qsaGTZ8XCEGhjSCYwQeJOuDBP0Z07qJFAZ
aYgQgJGlKdy/BDwbSleceoss5znKJwrc8Qp+kRuCALvCxotNy7j1BD0B+fk7A6rF
lQD5gjCbgd5paJdHqEG2qcNGF3t0DoGYXdYJuJ+PzPnpys4EZbPwO4Hm06YlI7Mp
CkJ/t9YFA9C0yEttoKz4gcygsFAUqPNzTTahIPBN4NixZZfcEP86GJH3Jfs5xCxX
fooX2Dv8/XrVwBJmrb4BpUpzh1qqvAfDeiPlLJlgnVyhCC8vIeJt9VAlU6vihKJG
cTYRgr/WDHpGq8DD4MBjrg/QF71iZy9MTqQfZ5u9cEV/MvPd1F06/a/eeLPkFl8j
YqHYNBWa19i6rLxO1A1dpNXUxT5nl93g8CZJFxOoFZDv5IpDpUt5MvpZ43gutkfn
P62sNt2rR2Dk6sXxD8MdL6QO9VtsQWd9NFbbEwC4viY=
`protect END_PROTECTED
