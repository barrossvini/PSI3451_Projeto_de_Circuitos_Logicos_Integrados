`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZDTzDvg/PYrc2Ls1a0AF36psnyuEcT/pCxkPhZqHz6TmDKCgVUjRVgfjz4ebcwJu
a/VOC+DsMH2T30g2uXaGOqF0UMxc4zvvymYaIhfWIHqpDtEh2eMChcGCdzSOckp2
fDCcG2SPWdNHWuQP+g8AKoObQUZ8Wrk//V1Y431YQQFRN2xikoFPbnZTAY83JNEr
ayNTbYyhgXfyU9CSrWnXFAtKVmhUqVOPvo3EXCoBI4ZxXwctvO6GJDQFKejsnNvd
VVlY0n2Ah+EA9v0XzrSO07urpFBAillVxv30Mg4WB20qsMsDHQqZ/w2EYdozG6eT
UR9tvdCGYTPxz0yNTFGB0Frvzv/4pjoTWXw06mYwJqmAqlo+VTjRSHG4AX6w6sle
B85gOUHnN6gJcp2/Q8FCjBiVfq3n078a1tuiKh7wY86X/FPgHRll3SjKs4cNOf59
SpElEic41BkxI/SwqDg7TclkAxrmKh/YwRRZQsNAUdwvUK/MqWrTsVvToKeznVld
FtapVm7Ihn7u7HegYzXywj/Lhmy7OvP4mWzDtq56ZyVfxVBdwsGM8KObdHquBKYW
497wGIOw/BwW8qXZ9yV6ITtj2sxiDeMb/zq0UI2Hi/Drfl3YR3zmsG6HF9yvj8G5
n8NPJ7pBWI4u73C8hrE+X3fj2Plplaeb9bNiDBqTHTBvG2zt96qPyZKwQP7l3tLf
`protect END_PROTECTED
