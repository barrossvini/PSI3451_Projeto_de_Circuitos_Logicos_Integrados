`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UXNzNw+fwTwLkPF0lxl856HbY4fbc91tQ2+MdRtAO+vgd6uQD3OORqW/jZk84lqb
lTXSsJtoLDkSR+pcfv7eVFnG0ouWokmzReNre27jt0TbfH5zwMSCtKwovpcD/sGH
eSng20Bpm/H98oC6vTgUr/sxiDQOeoVVzLosQzuvnd13nYU+ZXxX+nrywMcqnSHs
tE/pYUP8znlihApw2uD90wyZVInoZWy6w55DjyiHEGfYOyrQThFg9MdXd0W5N+K3
/AHmmNHqRnJh/Um2mAKB3B65au0gCJzYAFGEweGAfjdjhzV5jY1rRpri16io3tDM
b8S71RoTtqSQa2JujZkazCULr6DG5OTwA/np4LuNLBwBPpgncnsHeSTOs8vnKeOp
SOocw6E2EaE+CSODc0KYNoAcIdqm8+OM1ekkbF9G/5u04xhWXKHFekrnmNW0fSy2
6HthcW8fIsfjdPX/3S6sdFGL0itIkUzbC40ekjJAmqOmjzDMv/pcHIJcIKDvHoe+
scrSAetOXM4A7JoDxsyIhtxegezYR3XsHoKHgFV2yJ4BPMFNqyGnx/aJrXZqMce7
SlniK3cRIDQMBwPYWpc0w+f4bzTW3oTlwWOdKwijpk87XFk04Eyzra09GzJvtEwN
8hgpiTheCF+J4HGTrxUxPXdwpul54OhPN0F+1oflW1KVWrJJnDngxo33PCl/bA+s
4gry3OC8SIWJjcdTnv6mTy9qQ29oFSa8hvj2Mx/XuVxFtSBKZZOc9bMKtixtrt6O
x91O7VwsBm6ffaJB2j4HY7KJzBSdg3OvRR1ezCrGAH+moqwJkNtcFgJDU2vR6S7L
4SG19ZbF+1gOxGuvroRX/FwZC5zvHsOZTnJDU5w2LGzPrmvb+/qjaS1qXOSbyWoU
+YNKZ17bGcyMqHEgYwdfe/GKHKvaoVSCdR9YQyI1Ox8Zvw+xZEVdKV3kP7aoCqvx
O6wnLUdYcc5IrCxdwUz/4GGKHYCG83TIH30HZ41I27thYs8/a0sageOCkRnuRxYg
SK8qGaRzbDNMSAvd7EuED4/1reP6tiIcMFJvoYtEycJgXye70jai4sOih00SHYKa
UVpC6t5+skW6SQj/gvRc8h2fX0D/fNZe4RZvu2q62o1hQsbaDb+Bg93ATB3zfNKd
9By442R0Kcd4ZxU5MWc02buDJU1TwOX/NT8FvydKClF+XNK/mHF75xEZBrvnwozb
egYTkRrKceA4BRAcxaidSKMyGGYBNSDrfPfiTjzQTDSv0KcwCxhYWhy1v8kGYKpw
fIn8VcybtZ+WBAMgU5xJWBVHLmNhWyCBwKc2r49cvJkHYe3cBpfBgTc2MS8XSI40
JtOIpOCyWDfSBzGuc8B+UKv7OQakyEwdmO9+hr+1wJuTWRv0xid8WyZ3mICZcBGQ
MH3MgC15xZz7y1wVX5WyjZcyC6y+kYOZ+vz8QRWlnVmnRfYu3zPLaezPbh4WQIGH
bePTjdbkKW+me3dWBAe1f5fhBwwVzH5wzNW8N9fiFAYoXuvuuh93u1CJ8QSB4XaT
JP82TmMQ278JZVMhVpD0rAA5sVVljqB8FwmQk4Q/54RX5sgx4k01pDd1jvjkmD9Q
V/ndDklYLjukjQ+0RCl38ztaqNmP3/kzUBRpGYK+B1OUx3bJa1URPUj+RJ7FC/yF
qj+J+STXOzP+XIX5gfeOHIb0ryWZFOkI/UWeeOKYl5OPP1jJ5q84JEenhfDWmPMe
uZVUThvpPKO7+SEdEwcaJvQIWSUt6yuqdOlP5jsqJGpXJoFWAy0r2ePJsELGOZTQ
ZlgmUegBllGCg241Q0ZRv0ReSiC84xc8cIjHhzWlcpSGFD8FOsABsGY4Ty473a9V
87LdrcUq8O4er0chzjDOZ8R8OexRV2gB1vQ8h6fOn1d8Ie4I/5sIeHbOFvfXUoPU
vAKisdCCrykDv/JxiIDUw4u6OfXWFXuW+ssNXc7Rj8O0ygLol3yGHuB+6hOHI5Gp
5OLqWJ9u08stgpiAWwbfan9BTfFPfh3/iKF2zmXTb572pGXLBLmFDyTQYEp7UbAT
WhQ7xPg99SLGEKeTD8Mhni2U4CDF7Wv2pLp9wXiMQGtDseF6J3qlFAGlKEAka27v
tWpNNFtcYdDYZRS2ZS+7N7+KAuZSMu697menxe5r9QPzYK0sMC3U3EEY7jo/zF4j
/Gk4GI9feohb9obn0vOkEInMNqYNDwU2kzQXuFuCywyAe2nbYKwKaZR6Zu/hmto1
4W8jnco/f8XKLJEasV69Y4YQa5Yn660mb2f5YlIVO1CtYlOEkkr6vwTdj3wqKZTT
ZPS56lfX6Nhw3gEOSTCCErXwLllkEllngh+V8ITKldUuF/4U+TgQ0skTadrXatyb
G8T8TrWeAV/rSdspJWnFGvLe7aOQI6CQC+Rlwcf43qB4BI2llScMQs2qQ0syCMvD
cPhhnSlaARwiXFlzuz/l84vsrgwAVozFJMb+7ue7kAQzWRdblh4oYxiRcl2fcraI
0O+twn1RWFe+KpLiEoquXdWAPipajEdCRl1xXFMzCzL7XXLOvofUWI9tLxy7JCi4
xU70McY55pFj0z+FUJBcvGvcJImn16c68MvwsjbEi6+rMnj1/M9dwTE7N1Ofsrg9
PD6CQ8SHUmabW57he0ItuRjsSvruvnQlbz8qu37Ig3FwOVKGuFhoomae6rZlcaml
XjcN2wP0nnDonYXEycB8a58y1DVvpFmHKcfBLTaQXGxmhnNlSElSWPhb0g2DO2DM
W7O2En6YaVBYspas2+WWzjq3TBip7SHn62hTAEkETgBOXpL0SPpBpO7ErNfzfcdP
t7rldz4AzePPjl9lwwnDM5UVYzp2EVwy4DKGGcuGICquR6O+9hzDyicydgy8Z6Pu
3vIGV0dhrTNVan5wzoA2T3axPO7MHqMY7q8sFJJjLT0ZucYQtH8jMD4KnoFVJ5cy
xT3ETOdHYV2aKo5RF8rhoxRg2BuBYwVMVdvEftJAjHBd3z3tMTVVr1h9JdRYHtfI
FABMr/Uzf+aTeYKUpI4ZpFUjMFj4Lk33qwWD22o0b9ueYWQnLwoseF6tPMJtTucL
8QctaktfuuySXC+78O2N5Soy5HYjOFBQcC+hTFEDX5YANZ08/O35Cpo34EybX+gW
kszDyDzbhGYoFvb5xENSPDqp7nfDwvvcqWyexV76QYpbu20c5jIgg2ZrGEbCt05+
TFKkEvqgdvGwM3xXkMdhM8ZkizDZEnBzjnPBuZqanz09NguESqG9rW1jkxCe/ACG
zWtXOwp9Q1c3lFETOe+54qq9eIm7hcywcOxjSRrdJ34oJZ7ioGv+6Yw0+/BHJs7N
lk3HdjkE+GKD1106Ivr3g2qvrOLPBDco3U4lvabiIwBZd+hmpmreZkM/gB1Iym4V
HeODu8nVdkEyz0rCj2jgGi9UprGnVGV9zQhnsIdVb1tjN+9CxKkBr52sL7PRy/UJ
lY8OPeWB+S1pL2umEsWZ53/2HvbmIuNvZXUM55+bbU/KTzacnJ/XQqH469aQJCYD
8buoiOrrHsKYm8g4+//Ubo9OVWD6BG5fSGLBuB1Avsg+l7530Td2SNBjAFWoeQzs
NqjuZ3h8Yjb/WplKs76jcpPiN4Tiq8m/adZGeHfnUnKjPcTQw0qOEkcbeOW6M4K3
7cqCWygnh+/tBsw86q0ytCMbY8DEpSn3wR41YzUIIRCc17WYlktitvoxnnBPYuK0
XVi4Z8Amb279lXGSkS3SACtVVtYoU046i/U50EjaNTD/t0+QuzBF+p9b3VQZgfTj
yjDMc6cC0Ebzuh9L9zwUtPT9U7X+fogjGNuGUS7DZWBtp2LAutDt0GFU1x/nXUB9
ICgcYMnNJYyB5Ls074KrQJhoekC29e6vDHcbGP7+I0XrxVuPRXFCzOVTyUzEQE6P
TKHbB9XhnzKyFg6ZpQwmNYQgCl+qkXitf5roAoABKkIAd8sYSMyLfnp+B5MpGfSE
MjxaVdkePCiDE2PVW5+5K8WHVV/4zEvFy8RqAsqkGrMV3GEe8HyxXs3g+xz1YsU2
4aHtqsxrD0weZxKjpRw5NkBZ5ETfQ0rEfNlcBmT9QgRTwT4HxdO1aaMVs8rJT7Za
4FAD7dSBewMbZ16dJ/TqQ+Byl36xdqvzxv5I+9vSFMWlcBNCbY8DYGnILoUMKt+5
wxTG4YBrl7TxuqnUJoCiDPJIELmluCG6pR/eNAW/pukRJppVn0H+t3bQepmXuPlw
U7keIMzYZE95Yv51VspxNOJe7awODW1EwlDPEaDjIWovQaOkvZJ82thfBkyP1Wtg
RxLCzHM+Sw/KTXKzHgdik7Y9n033bshnLRdYKZGFxG+Nwo9uOoO3q4XBAM7mkTG5
tu1zTdrLP8wso+CVG25Jth8rzL5QTa2MBXDgMOTkJMoc8q6vQVdPMPkS0hxxQuXE
oGZuHcdpaYitTxr7VX08BVO5fC7gLvk4a/C5xEEzSUNE+izL/I/K8j/EJbL7dMSb
DgrtPK5aJN+etaiypw5Gx9wzRfiOhVpquizxtLGnpUPT2s4Jz8QvQc2w+Urvh4V3
ow9avEk0EQkbGBr3n1EhQdX77vSPcohafhJGqmNxDSvBtDixo8+iOD24zMvrTg9K
`protect END_PROTECTED
