`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cRM+sZmkwfDAdrCPqlzTXuKLcFvgxawVfxfNeDn0oTTZIJcfMJ813WOiFC6gQwFb
8XH/Z5KaRzRyLwOgbBxXQaTIHoi6g3fiWlboU//hslKXtbqpYy4RKk4OGbRTnH4c
t0KT7ajTzDZcye0XSCJH3O62c1HbppJMA5ynBKqqAEbHT9rI9gm6/8dth9R4SBsm
oE37V7W9qA0TUlNqJ61FWdIRdUFBZV0PI9j9a8tEAOFTDAH1i8Kta3fTQdqCeCQ6
HDd1xQ2JVmtoromn+VSk0FG9LIoO1CZSUcBV2qoIb2XNw+XAU81ueSRlz3wnxRmY
CQlhXv7KFnPWWpFj5GYu91hjzIqIRz+kHfnDqoM1Zr84eHA+fD/pKWzL5AVPMLNv
ry3e6LmJXS9/cK/QhiyXw2YlYxP1BjSJjzcvqV6pmoOYImAP3IVuQqRnh1tXVGHd
4XwRkoab3GI4wphsMkeqVT6MMD3Jy/ETvhtft4dGfbl6mSMoarkFSlwfXvMpoe5w
CCcZnv+0eGKAEjaaDk0aqXhqHBtJP5KCZmA0WlyMw5VvffliqhUaTsMcHez21AoW
CPrwx2VGdc7jYrtQI242G6qlkQh0ILlhvzRyIaFuo+HybwgHKgelee/tgDiYCCEw
FcFsCTFmZt+IBzzSsJa61L/GJiQeFyQgTKj64QATyWbWgoGvROlBWkp/FpYXsuK1
vNEx38wa2i0ZTv1Jf47UxmF55GJciloSxCjdWs1iPpVOPgDnGupp1EU3/KzAXo4n
MXW+bBQKVU1EoOrL7TZTBou/Ar/jERKpY4tEBxUPgjwERQmz9w/dx/wd5tEDNS8I
Ksy4Xg/pxkHDoy9ZYBCn1A==
`protect END_PROTECTED
