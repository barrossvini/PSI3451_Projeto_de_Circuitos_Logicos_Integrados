`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VcPg7/aDPjE+0Yn6c9SfTvvJmcknDrUj15G1ID9XQevLOvC8K2lEXmYFBU09AeYf
FL7jxqn77UcQYcR4bZJbIIts64DqAs6zmNJXVLMZbT7FjBDm3f7AON1MFa57RtZ+
sRQnoLB72frAiPriQY1nDsdDKaJeRq/ZlBbZCljxcKbEJFqQeOT0vdYl7CeHH0hO
XR9GAX2ovFHsgZ+FZLfQxjg2Sf48VK0TBOfNOgHjWmDJXb0xzAuPsb/bs1k0byTs
SYq0Zn71DxHpind1gmMRvA==
`protect END_PROTECTED
