`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NJPrH7qpEqZhXj7Z4n0K+OKAF0oQ3aDfxExeYBVDL09wTXHFOSGirP37u2CRfs3G
Y21UmlOKSHmTjb2Nn3DF2lthn8yeE1Cc9oKYO/7t1J7BoHstfT4lHjS3SYAVND/A
SZshvKY8I/vmGGwEskNs7JWhfrPZrWth31ZNYT2+jssErKs1xZ4XHxs1TgsP+ZVg
1l82uh5fdwuAhNSyOYdFTgSUaPsDIx1AQNwmGosZ6jX8AfmGeDjSlLCQHWZcGB0O
oi67nwARXXuBczYEJWtgHc7MROGxheSzRqM93sUia5Dq5r4IzFB2MEevyxeV7EYV
D3nUPdA5H68nIJhFF2npxEOHAvVrUdZUFNuCHRDQLQpywsLzm3HPdKmjMYhpNGFw
Wmdd55AfhdlsN+wQokxapU8tGMZP97zIXt6SRqP/3XEvNnanJywPY/yGDdUx9MiJ
PQ7d8PasHKE5p1MhR8vBJzrraa6He4Inrp5+L8tHpyoA0D3QBVOTL0FRmCQhf08b
mMcePbUsGvZT9AfAcowOwRazqoA3TXvsgf7A2WuNRZmWdjiMqOBd1qFMm/vtthA0
AeoqaONT9aXD/MFxJswAP8q95rsocvOnX60md5AwmFBBR3ChUsZYSAXd70olyaB+
IBwsLvN0iAILeSE9c4AWGu/28tAGnZ3YNBuMWje7VaUd1DhFOrS3HzJdAReyNSpR
NW65Lhe5eBRVwtyPYY/FhzGgK/Di6Q/u5QzAmbc0oE4uHClbRjDFCVmIS9VWt3ic
5lqXh9Uv10i1M7XtGLasuXXBTBBZ7h7uqwkDY4La7X7x2prwdhyycl0x8LWk4+vr
SmlOwZGhWfpy2VpbE8b7Hg64BzXscifCQrRQjyzkEMyzPyXeG1vqZWg14yosiOUT
Qy+1o5QX5yagOrXu3Cy67rhX65E00gANZbWqEjxlP0aOs8hBTiBetdeGWR3hO5US
Pb9hbrZLPje1+bR5IeXJfDI/vLfDp+Qt1BMLZD212GfROoEka8bf9ZNBsKuA/u0v
p4HqJC5AoTaGlHw6K70rQsXCCgUQFdakKtrs8aEi/dM=
`protect END_PROTECTED
