`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ghzsgdIlcg6qVN7J+6GuMAc6j8IPo9yYYulyzlyaijAgq9vKrQAvwRjTDjgsvVUi
asbeGFSn8VBvVvEUoYCCsya+Ct3xhP1tK2LWb4URV+0AjauVHm8TDz3Gyv5Ah5Gy
ebq4lXkjMG+hwNpmSc6STMLWNSls4U5MEZqMPV1ldAM/ThYBeim7SPvNnOxFsvlC
Y7+fTEOuLZ3s++TV7QrhKg2WyAOqA9kcW3BQVrTUFFS2qDetpWy61mErqTheZ36C
F+XxV/qBoG4UMMvayshgofhSjyYCh4EATb9tafDXedO1XmoaFpDP+4xD2BmmP6tD
gBRSlBmBowgncrV5ZXz5SSyxPQnEF7kVT3rkD4RSXDAhkGcLGCcU1JbaD8wUIY8Y
iNyGanAtM/wrj47NsY1R0AT/Ps93SRI8gO3ur0BwAQXf0P9Ss9sEFhNaBXAZu8Dh
L7NDWd71qFIqY6Wu5ID5Jt0sXTm5WwB0Y0xlc5mDagxEzPKw5q/SvUKMNEkxrKE0
FYViRKlGmJ65iZLjbNVvl5n356s5InAMmrFUToLxi59B2W7zrYHobeyKBD2hIUwJ
CVBnhXqLlyEFyVv8BK7DWypBonZp1gA0UNgp/YO0t/W0/pa6buEoi8FgHhog5dAT
p+UXSVwHAFRPLW6Ue4Ve+JAFsIriyXKqf/Vd/r+r5KIn4I39VBTGPv8pr99Hcl72
B4+qkebnJq2i+INTeESm654NvaBVlqimGw2ENmb2h3eV/XhgHQpLhtxNxQyzd3oq
UbV+1lZqskyTa8SDSnQa1pLXrhJ26fjJobUHTBR91dtmlTin97+wBxQ8nJkJDGBv
qrZ6/+B/k21gxQrWarbplSNd7E0wpdL7ZAu2+x7YKh6a7ut4+G4JGmFG3Tkkb4ti
MnsCncHiSqb/OXGnBqJdKZIR0flV/T9hCzQnavh1DzfMjYHFAzneAdbQOgI+vKi/
DA8aic8CFdprHkolfiNYHMip+pjKLeJpr2HOkOybbk86+76H1+fBcEIVFU9Q++v5
6qsN/6twVdRq4GR0MxivHzcjaszuMvFy0MoxtVmP9EkGEq/ZFBpVXK1rShJNAUUe
I1Hm9WuPbcLHpsd5xzzfps9aGHsVY6bx5RWNwo7THJLQettY9GEiDF534Q7CpTSx
ORhiNnzkoZ+Fuv2lhcyNRXpUszSG1WsrDaqbfA46YpIE78FJBHoH4jvjZNycomsd
zrKPqeuRn5DHxoyYpLFPBWmQT3QIz8Zs5gb9LSV4olo8kRjmvVBjQuztOmU0wa42
xlDnSVRzJ7H5GKdDT9/rOfrL6o3a2pbXAOFX7QrBchC/1lYRuu1O3hTrtDUhvCAX
+2Z2p6SpYLSvNYeHPHuvbFEtwuT9K8rZUT7HMx9kXj8ZG6EK324IDqZukaEklcJx
D5FAjX5tLtYtK2YXb6M1Gnnl7qznhHMfxePk93HC9XEpSaX25OTTzVIMS9k2F26b
zmtjCDePK7ZhjBEGIHo/cCAR7zTPcCgqusA6WAC1hCltaFOxzRfsZy+kV9A1z6Ba
pdSONEMeV41YwyFRx1aj9/BdZcXn9tg06RQ6WRY2BGQ/Lt+wdLBiEm9JYA2+/yOS
ZxperjbBBhND+E0Ne+t2dNoIv6gO+PNuyJQJAuzN4gq1xbe1qwU8Dp5jtlUT/CLY
p7maq0Nd4HSYPj1qK62IBnrWT1RAwBhwFV3xMR1VN2OKBV/AXaIUlfM885APHr4Y
HnwMfxwUntbtFJnDnTPbdjgopdAhWPzdbt9o5Ogu19NHe/Urq+KfmEdorXlTeE6o
UZH4hgtdJT4b9DtFa/Ao1HiPyFmGQ+DNUEj5l5Z3MjqIXZYf3YQSGIsmJB5D942l
CyZ7NyBgzVqjmIZ4kdTL4wwQa1E9sUndc2i4QlQ5kzJlZcKW+QN3TVu+7wsjDV62
MNwHqP1oRMKtaf1N+lflTjB4aipgfJOUfEnqJdGoS+TF2pCn5LjiYUn+m2PPeBoB
zgeGRNwg+2gHmTwL4NCr8NKn8WApD4OFPDZHw0SlM00YxQvg/DQVc01w9txQB417
iefGBQjQbjTA6Xqr4HRQoPFnZEsZ9ZYJXpzR6pira6c8QU3Y9A0o5tLdoHsHQloy
Ch5/dcGpntHKoYsfO0VVh29fUYRMsDFwOG9g0iholRqD4pVmEbEz/hPKdsQsi5AG
YZ5X3FMZjALbX9vz8hAwsM2AzxuuD075pR1xeu/xCJAY1sKYqpujEgadhqz29C2O
Xk/tO2uBfw0GOus3a31rTLGYgnL+ljB5+ZiW5vNVUVR9765UQm1TGotywbPV+HSJ
qgDn0hY5Lp0TroBlIdB0s7VLNVD8XLAf5gEGNe3ld7h5VcdBKvDin8pvVSDWXN+3
jrpKR/T5nLyi0WfK9EBiPDbCj3hTn17LzDw9Re5C1fQIWdRNSDJYebDLIjX7MnIF
rWLmwMG8EiEDAF+DopOLATMuEHsFFyUOPkNmHOxAXePVlYV3InMh1BlvDBFucc93
t2jNTqDrTjkVjfn3NCOvyb3jalvfxAdwTEWwK6WYjovnPRTHusR9sssp6/erRK3f
WfYOliyuQKB5X2I9fyx0UFriE13BJZ/IwyIXt4IMg/xi5NNEa+L9U4S9hZWXZ25X
sDYG5q7fEz+ol0tIdLbhewflHA7rUzfeMqYwtS2dVrj24TJukMNQCKqG+nWJcEyr
oxGWdALzrIPQOxO8yrZg2KhxHNsojB6p7DRCAomlrMBl2a+tkL5w84YxTitlOM64
ObBS9sN3X+jejT6AyEwJ+EC9Qe/WOVLXkbsU7S7wI12HxvSf/P/FrnhYu9d7D+kb
wxj/D5Ye0ntFbhX/2s9U1SBAOALrRmSai+BAXcQyukHhnC1OrOe+FDbZCALbOkuU
rXBszZFs2MssSQlQfGdRhF7i6W+enscYtYhfeT4d3R4xqnzMqFc1MzolYuthFRHk
/6tXYuZCPIL7bL2Pym6tGMJ2C6dg3EVpfbX3de10y+vPrUtXmiz4FiUGSKwSQxcK
i+l8v3uu7sLvgxcLAho1ebFz/gEOz+SG+aSjfE1jMXVzvnD7hn7nBae7h7cTpoyq
9uuFN6PP0F09GZJ/Ce3kwD1QCY/4wc/E/HWOn9q3sKy/4CzWffLY95T90kkasGh5
pTPw+Y9UTp4w+jnuUYcMBXSzhz9V6yvoJuM+yWMhHlEnwVxMYO0UEHtI6GaeJIUU
Yo0oYcUid+wTwgR5m/v+NA/diF2JDdXp+jRXVplNUMUuVNjC4AJvVtStPLDjdZQe
BuzVY8hTR97fxYWSSWxmvhr4WxtU4v7jh+j0QfV6d4LhnqagQfr+LFcoBjOuSBUr
cF5pTzjE5wZDLOpSxw9/yNFhJLRt7CW5mwT4+2OkWWWdReMvhMKc32Ri2DZu677k
m1mQIWlcNhSDpXUKuLbGEf92TGSBFJXnTFOHlaev+931w+M1++7vEbNPAPWjh4zV
fV5Wy5H9G5f4R/I6ZVQWfg==
`protect END_PROTECTED
