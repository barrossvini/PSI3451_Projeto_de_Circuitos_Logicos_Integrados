`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AB4BGHK2kbEgMg5gti/frG6zr0ESAomklJ833tbJ+r8OwHD2/c/Xy54rUb6tKJxC
ja+YWpX8w0Q3nHIO+JLUE77jpyptjCUHh7ywOXXxzlJdjjOLZs1ZXsmvUwSijmDn
nh9APmGNwvo69ONKG6gnC6S1bIkE+SY2AL61UCW1mno7oKyRmqMmy4xu9pxE62t2
+JgKM/uRMk7rd0BBdu0/81Fi9hbSpTkavZrJqT+IvHPsbpOjW8rytN1tEgnUfm2L
jP1eSJ95AQrTVNp3KNvq9bz/CI6AKSgLph4iyM8ThHZOO2sTAuDDnjGQft90BsMc
nd927PXqpWHpHL+MJyCcXXVWmw3cKP32ut2aejCw5Vl643jj0LCYh4qQqxehOTTV
Da+QBr7FXxImAz1QXe0s5uWyr4uge28IkmGXRicw/nQOwlYQFlxXC4buOJtc1pm6
rgCeX3rgGJI2isFYaeXhzaQU48YRTU56EIrXN9AAafVATHux1ZH/j+s6AVMLFhLn
B4DvI/O3rVutjMhidkdA6qqbszShXcM/W3FOx93dnx68PgXOltX0B2cH0ridsG3R
LQR7nHe3GJPSy/V5F0fUGm09NEmT6Lbe0IYAnpfnlBm+q0bAVief9SrpuqJPaMX8
MExW7YWwFobFVEXFkpv4DTI3YwXYMfgy3EWBzcd1q1s5SszIccYjiedWoHkQ7L97
p9Kgcqh4xlbq9OAOznXtHwvE+ridQWHYlcQW7sYaU1oIeOhfgLDd35zmLF1JPYIj
9mEUgp09CCTYxumUGgRhAzXUmVYc1owCrnhKSsUt23YBpJ6zOPhSZAG+CQogi585
E9PpuHwnnsWexPWPQMNo0Gcq5EikYJxZJckJGd0dT1ftIYOfB3iyou7hHDkwI4wD
YKf2TWC3CXUg11q7yZCcH5uKy1cuSlUAm/MLqBHGQ1KL2nmaIh0tt2Ny9gIDD0HU
bbVFSQk9nZ4TmbReIB/iqqTQuz4VTlygRItzRP+5PRZi6Sio+nsZBJAkA8v6Wtcj
jMs5IWiJ5f+P5ciqjFXMFmTrEtXutjgU4DInEr9u73fSA/OO8bR6NgPQKzuvTNkH
vIpdXzssk/LvN/HxB5hrEq+0r0fKo3Z3rudZnBxF44aquTGS80t8gDBlsEbtpJGu
WgIiK5nwOXvwVwQByYj5WSNGEzS9OxvRnuu4lraldlLGCwLfqbmQUD3DmFYlQiA3
EIKh4mxgyzzLWYVG4nRB4KagMWXdgfcGS4Ias6W4N5yS7xfK6JUH3ZHOP5nq3x2f
c6iVcqWadIlLyTsK1N2YknG7U1qUHhvAMjZHIOcM6MkJik2uln+2uAq3Puazv3qW
U1eaxEoT8hAve88yA1V4n9/43y+fCKVH/btZYP7kU5brRjPoh4ClG/myLiXAetOf
BVh07RwmrSVj6ECNNIA8Cj0L9A36/SplaDNr+Cu2oHlcCkjCCHS8HSWy/vEG2uiY
`protect END_PROTECTED
