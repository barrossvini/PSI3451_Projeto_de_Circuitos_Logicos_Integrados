`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UjomtHv3+uh7JZSSMB1FvtEJg2Rbjw8RYMkFI0/aPGJ65jYDQ9p58HEScFGTv6/o
0XD8vbu0dYf4VTiNxcc3Dud+B0AXDXEckhsuymUzU1Q3Xn4xN45O/3i/P+rB1BTv
WGLgiCwdhaDLCemnFRSppFelG8MLnDv9gOXjqqDFDIF4Suc6fCUhz2eyzOzcLkdE
k2r3RqCzYadV/eb9zTdfJNMom6KGigmCEm36UqBJYTWgUJLU/oPmkm6TYVQnJM7a
lbpCG2dFCMLWdvxtyrpeNCSH6M7gCWV1MP9WutBnmUxWp8tqcGUxufHZA+8Dt97o
iSOxw6aOVHv3MN8aAkoUDET5oKUDDF7Z03utNWHFLy3iw9nXvaEd18BqHpsWgKAw
Vl6ntxwvk81Wjbi4TPfjT7O/5VYYuaylCK4jc85KsmMBQD9vCsFvZYSw+VfuNtE5
bRxPsHAYSEVcR3hd4dtsE9C4chN0A5Dt55K/37i+30KWdFARY6KJa5fJk2MGOSnl
TMygj9p8Zcwxzej5w01oO/a7+81K+yuL8xAcBlf7rs+Dhw0Tk2XzQNLGhBtkxWmr
I/e5adc2NZEk5E5xyJLpEajHruOr3fvBkZRZI1YvOKPRA0h12zBlKSB3LJL3W89P
qfqt2XdMk4PE0m9h1/JR7Vb3fHEYnaDfnLLFHiX6GOXoNixZnRPH6li2XbakGeEZ
0GyK6GDDg5QDwzZ/7mN2U6phfobB6y1oQ3L7ipqJ8OWtrzPvsSUL4dBjgEACvHNW
piiBDG6QVClyaX5/pVeWiIvZf1xhkRrL6r8sCUqBNrIsx9EbbFFg1EHk0Nw9R3Uq
ZkVwXyIX1ES/Tei59UCeXDcLAw6kEFpT6l9H2jMt5eGK8Sp6m36x46gHLaVDTxJE
4yFQD9Lcz0553mjbZHVR8phvQITaOOF+TQx1/9otC6UDXaqtRm+DBORbR74uzw7Z
McvLdMAO/EZmkbggr6/GynTe4dfpmBH8dgNg6uMr+jobXTVeI3g09WPPsvS2gUBp
QkRdLx7/sNyDRMTZ0YlXJXxFgKin54dMyMxqzAaOslhnoDYsX46ecjNtegy+DBGx
+/8tRglKH57Pswn5dyQ6CYCd6uJqqifbb1toVZvHTwtpj1Vb4X88uA3JmCOjEpK1
tjOg0gk1EHLjS4pQzO7jKisXt46TQ/4DMPnkTtchQrSWUsVFxScaR9RxNvKUh3oS
n/g5u2v2MZaoI00pl+uTdRbmkkRSwT3K3+WyLuSBF6VpDGQD8+DLss4VCdXs1+Ui
sfaGwCbByrp+g50aDag9djocXAHM82WZpdEQsN1b8NCY0XbpV90OSRDzgcE+PQTD
ku5JdialLeqQu00J3AvYJqpNG9SyMlIUSgLaZWdgOXObk6k7w6lMsRJL/5gK3jfM
Tiy1GN6/+uoD6hOk0zWyVjgBiHKT3fshYJNVJuwKtQlLjfUNPWVkL1GyOYH5Ht/R
LpI676gIcKJqGHAsy0W+L5fIDp+4aiolkk9Sf1dZtgeOYlpSYy6tmAcDLoi5Eytp
WDA3onUx4ploz4Gjw2vGKW9X5h4C/mcIBn9dJlSL48gs8LbcBGkLQoQX0DVxrWc/
wyuPP1zGgCzV38pSB/yw59aZa67HvXHaL27Z7iqymztEpBNjMXgndquvFq04yYOM
qBJj1xZupz0PcHo7TXueZ8v107c4oYEydOsTTu2thSE+NjoTb1RtopIGd/TdaXGg
J1ytmnmAZS8cHC08FNuDYTu4O597aGKgM2InMALOoqOh9NVilTCx+VBxPsRZ8GgJ
hzBP2wKaWd8rJ15bflB66LrqaEdSaL28tx5mhvdaavpEyiQZf9TIV0MCVE/M71V9
kYEs0hTeiaB/oDC2UySq/qVyBODURhNTO7SwoG368G1f/r9rlHt7sMFJ60I4gKbb
5wexTyWqcMd9DvgpRbnzd+xBOIt5/hTN6Ka/HoH9WLw=
`protect END_PROTECTED
