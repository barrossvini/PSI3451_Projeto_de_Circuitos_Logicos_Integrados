`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zroRKFsfDfUgcTnW81m5kxLXymSR60rr5wITV5hAgkepXVAUuTuF3wdtX+qeGo5j
AjP6I+c7SZJ2GPeHT3oQdRsjfF9JuqRrCFtyHC32FQK9eW9W/EDhTbcPrbWtuYCf
qGkQE4awO8Tj7VPtQGXP+ysLAmR5VGGqqIbuEh0sRt7ZCaiHUffdNDpWsNYERXiW
0Yx4njpxwV/EDg69tvL1jOUUfmUNcgjRFg7IBVCoPbgATHLT0y5CdYkoXmhqLjXL
80VGIDX+JP24DUwCSSY99fgKGHQvFY2exKh3XsnYeykdCrMLGZp+nnVc7+0gfdpH
zIWLqlzcRLuugFPuK40B2mymQJgNmxvLq4wCSdZIsHSI0RiyQyj+6iim1k0bvm3q
Gm0v27NbhYBQWDZC6STjL3fJ5s+drQ0YRtobj0sbdORe6/rlhRUOfzQqrKnAkNM1
+/nEFcQMWOzXDTneQROW5kebXeoft/Ly9OuutFBfFdLPx4rRUuHuFDAuwDV2kp4p
GXBZEcbSX0mbdgSBSfVw3aQGuWZt6nwGrr4SWeHOQnmeEsYtuG1qiYhnNlPzNY24
Zfx783F+Hj9RpG/bVnD8Fok1Z81352AgoOk5k/tXhAyrGp6x0duZoGMO5GHoYJqi
tViGoGxXF9zuybxpW5qt14cO/lvYZG36aEDuWkhmZrOtqklfiXlWXfZDb67UbJRk
iT4L3eapUN92Ru/6cHnqdV5cFhay9iL8c4O0q6BBu93jcpesHZb/IcAMqEjaQVdv
UcK2iY1gk04ttgM3GTRRt0tMzXy3RNOXGQEk5CBw1fu+vPWOrnLuDRaiTMSAZ+H6
cZVXrjB3GpeN66dUW5w96wRecQhQHFxaYvFo1l//x8NEuh0g56/RuVLw80bqMM7m
dJs+AakZiHlvKuMW9vGmZdLST8MfjdR5SRzj4P1P8SR0LT5cTDSTer5WHgFnQ1fw
M42tacIk4276kgiIyqjZrmda9rox4jXTc18D4ZyysnFNrReWw0thPU3tGGQZg4sG
LJRre1CoNCPoCp4zE3ihlBiU9DKx/xVSTBQ9v396TZ8+u1cR7G/EhrYMrI7ga6jf
n9Q1mIAsRp7QYRiGUD2s1l2MFeCShZqcimFasbDodUiotYr5dTkqVUcZjhx4ScPc
6NUIn+YSaS9YdfrBOPRf/kpRihstMBxmwM7BqwsWXetHCzAw0RxGEw2XJV3jnuhg
HH1xPp9o+NAm1FSGO05/jHKvSG6Ztnw5DjIGZbdBBNh2gkEBi9SG4Dq9tm+A57+D
B+nPXZtHgZu7p69Mo+GqVluZa5AhFrU68jR0BvFekHmX2jPFq1UnrQMNy4C4DPAD
EL2/HMiGvYADwCJr9Wh+Wu5Y3x0n1s4Hd078F5GPzzpiJUZXoNw1a7hMdrX0IuFH
THHRnGpy3VywxIde5Wiqxg9/PeUXaU5OJ622/wSlBpIwI+2b17nZNUrgjnzl62rj
/RIokUvVRvntorGrPatiJpGqUWLWjGVE4WjOLyxGQr5tK96sh2HnJsQGTAED3fHg
7R4Vvu/eyhm7AFtO+lJZFXrfdVCGb046CpmUp/lvsnAbcjUa2r+0TwHBEahGX40W
1bfA1Pcb7jJLZmXVXR8jmdGwOvtqi/rU8My5yAgzgi2uovhNYjxzD6ukntNDtHnl
/EmXzBCgC2V0G46oRIMnhH5bkAqxOIY1CJSS7JaY37wPp9CRAkj4adMzHGNcclvb
inV9WgagShch5yX/7rMWOi3zwdLyXgM2shpcQPRzHPmgXe79NMDb1pCuaImXsz0B
4ENPTxNIiDSVB6J3oz8SJXHEMtm4JW30UtwuC6fncD0iZHPR1I/GL9RqiL70P/fl
zqzZ5UJ9TQnjplBgHDiEG+xQHzhIIYWUPgVfcyJmkQlLaBH5WSDJypOPqdaf4NhY
1UrIrgKBzJjUg6lcQFwViBWsTGp0aZRdj4jFhbgzBBVm4oIhqQ23vGlr8wb6LkRO
K59PEosK1QJsWMKMDHCGrR2PdHkzlMRjTyTSMkSg/Icb1qhKHOISv3F+YFPWXj5y
nqQRBAOrCplhCH0lhgqLbyiv828BGM+C6LxEADh3WtYgWyezxKhG+E1/GgiAaeOx
crUmIfKOHfDb0S/qlMhjmIfgV89kOi+SUhIDVWeEIkfO3s+0EvPkTz9rpCHHSTzm
GaNyMpY4VneB6924+bVbXnFZPRz7YoxZy1T4rxlbu1zVjSSuHy0LzXNsZBwGto5m
eKBfVviEF3xI+QhRUntBFE469gE9h+eyXncj4trgUyFgS4yZ4+Y5Qe/3ysFvBzrk
LQkYuqtQDr6JafIM1QrX8cY2pakIUY0F0cNLpMip5gWejQdFcmkrZQjudKJBsXiw
BzSMH0pGyzZH5EuosI06aSYuTRMynEN3y6hv5340OneJoIor19tw+8pPpo0T04y4
WqgeKKyyC3O1wwAenF4G5mMIUAnDVgr1cXouxx2De1ALXOwQyBUPoZITY75dq381
t+p26d+L+rgFHeNED74dMKsqhLMkKSjq/w1HpRLF6s4nK09WgmmJUIq9P7Jwt/6d
s4JcmOvpdZ8cd/zWLMtcPRycJvulCbk31k4B4F2bzbAjwYQn3xUXJTF5ssBw4b3d
Lefc/Eq0F/ushnJOf4VNRo7n2TmCYG4JIqE7I9gmGIs5Ry0k8jZvdy3PzOA2+A4L
sKzsKcuoZVHdKHDglibzyw21EUSBSaCHcof5g/IIyiAzjYAGD+UE1UJXbUaH+mPD
yvo1yPtAfFwjQxFGLedY/bJPXUSUe+J0lnxWr/aqnghRENvqoEjT1Jip0gFhD0Vh
wzNFHyVJZR2jU7gZlMUlZOuUn7YHEs9BwnL1CO62M3RgcgZ7zpob7fZF8KKgFjOZ
lRsMqqo6v0WuZYl0cHQqtXFN/I/G3Qvr3RQNh4VbPOnB2rnVx3iCVhqT/3PGK4xj
O1U5HRAp20ci/xyyvEP2gGTL7tK3mioN8vxjFuf/vBNjbFQm7ElB2jstNe1zngSa
XTV7RrofuZiT/vC/ZIoe83orsaX4PpfDiUKTk/6gffjL866DiP++54PnQt/2RcR/
W5osqYNBU3u2I95lEbnY457mfpC5UiFUSK22OcrJ7nUGA2PRGp+zsoXGbOL9dg2I
5K+ZkzR+E9K+nAmGPvKd16EnejfIHsf4J/jYOKQpwrMt+cK3Cf9JOFbLI89cw4T3
0FZuxM+p2Kevv1NK/eAKmkR+SEOClk+LwY8/TFe4gZ/umPpgF4hP1qCDzp/Ve5QG
x7mK5BIedzmknCxhy6YgOY/voxVREy7wytd2bZO83iLK/817+mWDZ8zKuRFxawjt
MS6WpkS5u6Jwi9HlgDy1HddAZvUZzOZHJTSgfNAoWZXJ5ILygbYVifOhecWsnHki
e55yc/wfNW515nvefkoNhfEw/Aw+6ZQQbU1V7hiEn6rBtevatKL7vPkt+nmiaxj6
MI75QkjaPqJjZmYTuVFnSibkQTwh6o9sdfIn++B+iyjwVrNNczdsiR6JNWiIyIQY
4knHjvIbZjtq3ewLHuxMKD9Jd35elJ16VGDIjKlTZkHF6B3bFMZCKJzhHpr9joOc
0oyIFdL9ZCfPzg7HTtGPSW+/IDesWKiDu2MCdRgm/yGmoVit5gHr+S3wRqmC13ol
zdJDGpyg/iTkem53ZHR15u1jIs8xTsBgOh+BQtQXOXIBKZpfbeb5ilHUWp6Asz+O
oDFPDnUHH7kq6oMakbvdtB2nFiCqEYu84enHbmtWwZBFNwD+xf0Rxw04gpNeUqNu
5wsNZllNbgo7ZKGGEYYdmsMXGsoyYatRQQvPfM+LyYA4tdD37+M7hn9/SngYXfaq
1vs33zZMo2Dxqjo4JpXWyzUpe7laucacQJ6FLouvw36siOhRZyFhyQQeUr1mHRqm
dWGcYhS6hOKbCXSNs+T/zBShrDoZhwbSB1CebgCkEEuFInF4mRKBbVHtepBurGyM
A/yKLsCbpi4f2a6VzGTf5qXPvbgDvOJvcLcMOC9dfD807KBDARQFu1QSy1WthtYo
x0dOW1tTD4f8rVPpA8K8+BBQRXJixzWTFexRQt3jbjOPByd9EBsngdDKdZg8W5x4
r8rTG2e2rur5lOzuUqaWZR8E3ZrpaTJOBygx/ZDGfGQH2dxz2o6VAGvB0MGExa+m
+xkLRxVSsNyEtlpLGR5o2HBjOTmohgHo1ZohCnCOr55383glXoqU8ucI0wS9EKQq
c7EUp+0XdRQUUaFXPqy1pwO0S5Q9rWYVaAwGeEuVPnhE9Mtc4LKnGByMjSrVucTo
ccpaevBiKpz/1w/uMS5pRgGtRS5pmTX6KBdxm496FiOQeI5P1L41vIfSHazNxI4z
boyZAXQUXlsCKfxJgygQLJ5OfEylcLGSjq2wYveoR51OZDT7xIZRqaLeun34oiWQ
13YFMrt7/RRiSuZrmtC2KTrPL8pkJ5h+C5NK0pguyMpO/ny8qZQJme8rsDYWeR4A
1B7bGO7EW0D7sSG496g/HOkKCVcOtnkdc2hauu/5Mpk7DhWqmJkXUdB1aSI5nnbH
DyVTyDPkB2F9rCIF7czaXiT6c4BC9be09mQtYi3NgHSMjr9CVZ/t+5A0jDCWc9Am
klh70VRi8yS0HnvGG38e3h/O3I9SHnmKp1TawNERzCUVmyNXCV78Iq0U2Z0mqjGY
pJNHJdcNQziBq2AFHLVQornzq0b/cVJ95fU+NS+htiJ4LeaTashIqQvjvlAjm0OW
jNPwPl760qGyT7VPvoopRTa5mmdrz3wKEkOuCCcaPrV7yxTgVDFJQ3SMXjDoVMtR
v6rezxjnAWal6H+/NAKJjcM9aV+ft8BsUVxmSbhOb80Cf/0casUyy1oQVQ5PD9qq
apSjE0vZu65Vq2w9AxYpupVlaLQWtgS6FEiab1Nrbc5kvifjjXpvaW+3qXgNi2hc
7nsyOik/IMJJqwj16Q2XKv4lfJQ4KMEZpXLMasQzv9kQx6crYphmE6Im++fveeW+
WzaTnUGXkEsEtuALoTuVkoiW7pqD7Q31v8F84+p06E8AVtiOz4R/ThgCSGOwxlUM
O4ApNC8Mc/0EpflntS76/oD2uQYFRHmHVhgfm/jLNcE9OR9uOhWFHVy/mesAZNsF
tD1f3WE9u+4ludHJEPAt9h1KMulXESgM+vGBW71H2pKcsyq86Qzwxg9Zh5XxyzX4
xFvSJDykI28oFuvilz6SLDa9nXnN4nHx7OyNzsdtQofpWze3b6japMRr/YM+bMUK
VuJd/uN7JvSuxXotJNbbjsPVBM+o+heLb93irpGQMtQGdSVvZeEhukwMyOE4AOVE
B4JYr4hWfV7oLDv/vCSKWnCZu1h+UWTPRjS+0ajBMdalBGZcdCZRFKHjAgOXAie8
GOykVduOXE2/dKWrELiCNoNw2mBA8f13D91hj74+ai6Feq1e1KaxiGhvKB3FSPcz
MsZHkmLB053irIRq3lPYbjBlZRZ6t5hsYjGySrX9PLirfMt3xSBvUKyC5YprVuxz
GT2pPD8fob2+CCq8uPRKRI6Mwgi7tu80xPyObPTniCjJpJ/4KJpLQ6H1xPEyAYGc
2bUUz8NSjegA+vFLWLpirNIJqxVuvm+FX6sgqXOUkxh+LYRdbE4HGPfCTaAqS54n
ZICuZUhetCpIYtJlFV4ieqX2+WhU2LU3fY6S3zJf+3PxxgEDcb9zfmfZjmRY8gZE
t2UnFZhN5aOECN5lS4oDgcst1OLxBSN7kqxtyaMCEz8EEKSQ9mgc3n9vY1Kclsgd
ByfA5o5i805r/e1GLmPuo6EsNPip2aOA4JXOX1RPap4ArftRsvxi996X2mxxh4aV
5NibTeKR1yZV+AClzEgu9W1yZjGxgfiYza4H3XgzkVhJqBw4qvVWO+6uXTFc2nBN
oiY0++Y2UhX97Dw1Zm4MqmuAVe8cKIFFtSZ/ZzmOf8/eOV65I7beu9LAhhgTgKeP
08hP5+jyD3ERH8eT32GpUAxk0cCuaRzOxynyAGwhcyf3tKQbJ+vtaL/jBJmGpLJf
T2VjNS15PwR07yiobVnCI1hBV/KQqdWHydFEusO1EWAseDZ1TtlhNvpbGeyWQzHk
8u7t7IT6W/vXiOvKB1AVingX24KIl1pLkCAy3MZB7SpIfaXOFtOqx5XmYKGRZekb
/erZI1qCK7RMzRXFCzN/q8FaCEO1K5XMcvpd8ioc/Tb5PCgBqBRXn2WIc6T/V3/6
Jw3K3XM77Z1ayQ9xwkAdSE1qua/Kh2u1Fxj3rTI86s61VHrulc6HQ0cNH5mGVvIU
flfRGXmF/EStRmhFCx7qtaSgNFVeC6THiV1ujdn9MsohkNGyrovpDnpZK1Kqsfjm
Xa989gG18EEfXgAh2n4PueRs8CsEwudmg2QLotR739RX4lI8jw6bSnDn5GSIyQ1T
srK3Hw16OgdI640wwskh2VgxEL5+orjTgO/Tv1MfWxruJEE1XMf5HrrGHAejdQ6Y
Uz0/Y38fnlU6oLgsJjlD3buXZJz/hHldZp9AhVyHR/zdeiIZMUrQQAWFKlgbefFa
xDnclFsA1lroF1L8uqFWvlBNLy5O7F6NF4F0seYNl3HGURtmPCik4bBJBkL1QXkQ
V0EXwZFIFbx3t48mr4fSKt5J2s7gwzOXcogmSCfLHpaoIIkHL4yW5qCJvLlB9hSa
gHlV67GJ0/10xVDLkpenPzrAYPF9y/Qbtuv+6VL1w4PzjOdlAuRbao2ph/rb1z/W
m9QWvz8P2Z1wrOO+CBPcVgB7aIp3ilVaCaS3bKYOcd2+Szoq3QoDI6QeHSwaQ5E/
Mjz0Z2c3giliZ5fuQuBApkEEIxcSKfUqHZ3syV86HE5elvtO+qQoPsWKEHDxVuCd
p1YvcL58fBi7YE2JSotdca76rpSgEof1vXKhPJgZG9GJGq0vqIkOafXkLKFBCF3f
NoJXN/YEUPbKtUVleiEhW52RewOtRC+Z/PH/iNE/wYoSuHBdO6vaJJghgvnK79PX
nMy2UnMbmK8I4crUSekrpiDHoanpBht7ouHmruC200o7njgkK75+waoWUPjqZ5YK
MZq98nFtvPFG6nKUjQ22PULcUD/bKRn70Dc2mq8KgYXDi2D9VIsGaKw6a30w9qFn
ClGqWlp78CyoMCei7tcK5dP96J0Z+RcIGuOaqhIVuhFv7N4V2KnlouKkUUkETvVX
217jVlSY3VawRsSVxBDGpFCj4mzwUFquY1X8p70Y+N+lKQYcq6yLd14UO1XeRtlp
0RvVf1fQyE89dVIm9i1HGXyLEfmtxiJfgv1I1TpoVpigXPZ/84azAxUCCheReIbA
tJ4FWVD/TsqIlDw/DJ87MGFtYnnjRsWLz6LL8lBhNbllcmodMRRd6ibMkaDGEllS
9WtESJ2hRVx3pFAsKRetpLP0FjpEUpZ+lnD2Sr2e1twcTHgejI9bqBvse2lLan1u
UajMWfFnBNbHLBwQq439aJmbDmXGt8IH/nsGvj94GetsiXvxh8QNiJZJGbcSwL/0
ILa6Tn7pTnLqw1uuf9HQZswc6PJZRVjXkgkLosZF3BhMNi6xwb9yR8IKMb2yS4Zs
4CNaQFM4XLJv5otjxii+tbZf7nvCSvbAs3eeZi1wxdFX98uhxN5RM+iZgAcpUfNl
ir3GW+QX1oR/qgYymeMkfkYpyQa6w5pGDoSfrm/DwnAdSTH39MEANMvkIYVBmMDK
Jg17CvE1JkqeKG5RgcgoMAl+2TiWjdYmXWsmrJBUDMmbhl9+qR1hBGiwvI0S6Jlq
Zg10HYb/KmoOzmpY9xxUAkwOBfN1t38AgkJ0DTCUIkkRei5RX0M9UBDyu6hmoC7a
8xtgQ/akIfg1BBwKlM1TE9vHQJFEaM6RSjNcF3lNy0sAgA7VpySGqIjqvhUttKdK
hcWFXeKu7m5gd96KVP3BnV1NQn/RB4X/U6buuwA1irwmapqZj7t2D6RwH5PQ1rNI
sIcxGbImqQsKGOUsfPGvUJ+uSC057wsvw946/AEndzsg7NlwaBMVKG+qLftkAfi6
oTO6MLFqUgD9hWfmXF0YAST2pQ2NCu6XInhOiUWIElsbQl+Gim+fZDera6yrVTjM
v6x3H5xmx9npEpqlg+GEZJqEZKBuYHMWLfzi3gb04zWDf98K5QPjaqqtQKRM8CGr
VyjTR0KgcII0OggMbOzgdLACGmr8dsGCdW0xkwsxoyY6+5TLZYZO1AhVw/WFIfkF
Qo22Btj5v3zQEeyCEOg8ODTfCFkI39C9KYWd8yi0VeUCYGgFyfQdscIJNmrAxLeI
ZR/EvYDLbnzIO2ZQEnEV0p11Ei0K/Sz2SdNeixmVFL2mJ8b2lrDnMcz1wsBxG6B2
sGGCou1gQCLMQtc4Kyud5oZp5gxLzwOimibCEhX7y8OQXMp7mMf0P6u3cfpfEApL
9tTgWi6pZdl0f53eGmV2aO08OPHw6PwQ8GUc8CWoJiVHWUkk9h1q2vMc0pedITP4
hZMIfDY0F/TX3LzfXaIjRn64s1oUfAHAu8+OJsb3VFzvzBxfOzoTHy90VIsX9S4/
W1fqUZlbiXADBKsGRajvBMtKM80m0ElTFYZcs1DU8PAA02E8NtVoB7vdwD+wtucR
j8XSs4CaiMZyY+nqjegnkyyqoiAZyP5uEG8zsu/7e5hhH+uu3UWyZm9IywvQU2kh
+StyiAWBR0I4YiFjvrGKe6YJ/l7ODgIfZrhJQcab4jevawLSY9ZvnztMT1qZsrrt
2gW/yET4NGEXQFAdAdf42M/8elBZV+h6EHziR/GgGOoPazDul4NJjbjyT7Adr5/e
CxSQIWAFAJ7mjhCJHjHvujjpL44b/hgvH2M27Yc/7UJict8FM929VYfXrJ9qEB/b
Il61idv/fIoqRnK0EKirThZwXCj/+CXQmhgPrqSSotWtUNufgWD9bvv7MAc5BVbT
g540fdRb4ZV+CvWwNrBiNDTwygKm4iFcBD11p90RIUxBRXvFXwFdxafWFSbGexPC
VoZCZxkmvjIh7N1pQoI5dRBpYE2XORy/IsbLqeSnAqpx6TecdChkSpPb8x22RKYa
zoTSXzVp7sz2C+fOkTGdy6gyus7GkmajXBQzFIBhrurpNgsJeAqD34Uv2nkpArDs
V065Hx28BYG9thOmKgz4fX+y2VjxrguSjIxC5VkZSy18Gco5Ya7NBKLIXYMDeIDe
3/3gJcdpFFI0eTzviLtk1cRYEXGcWFGW2Y2g1eq44RisKdH4wBtXe2FX9mbfMJIP
NCPoCF0UeqrnhQRHSv1+wW37vnov8FxuzNgeLqbl+8BiCxBZzFJJM6+SOh5tQqnK
50NQmLz94VbfrSp/UrWQe947oV5MLTr1a9PY5xEWVtJhS24LfEgojGIBHjb5ckAA
f2Rhegp4L8E5tBpB5vSHNgKFN7XVswI/fkQ6NrpFgVtWCtSyEIkcJhkQMIE7RREe
ORvThy9QBU2Ekf0K0C8y81HYQkTt/xnQwHRbW9q3ie4mmuJE/plcdFXdxa9O1HOP
Fz+0VnrN0HQnt28ncQyhK7xCau7Tj5T9ZVicWNhAimPp7UJR5iaitEJBLg8Xhuch
O1ptYSHVkOFMoHS3NUvIU+zz2HwEVwGILLfvFVEgnMv8jeXF9k4TVG6fZHR1hYjz
M8tVX25DQ+kXEQfhWqQ966LhsahdZ5eQq9syHm6Mywgl4bhhVOZSXsTEqrGrB2IB
Gv7ggI2chc4IKAflj7v+orx9Ii0uG8m3aZs7MM35udxRXijxhnhV/XWrvkGHmIk6
TVEcy8DB2++/QfaFUZ+l+27BRg4kuuiLtYY+r7Fv/ifkq4bVKo+kg8Tg5QzF+O97
VebMU80jphQ5hyb6vI7prUod5UHLawD7RTOBY21GzjE8oxw5N1mfNQQPiZ10SEi/
c3Mpi0bcYAePhkjAWY2yp+qnVtgtYoUM4vFDdf31bLVSeCAICHNXdjXbkG9LyMQW
pKZWBZh0/dERhjiKzWvSri8NCzQacOTfuJjFyHH7iIeL91iC93AvmoTvZCpay+iQ
ZlElMqpMpOwrhZQ7p+vo/kYQ8tiw0bAkm1u7i+afvykQL2hOYTKN/C9sI5dpXtOw
gqxErw37O6uCtNkjeRwIOY8NrumVYDfClqvXh3xB5aYDopVFHKgLlZW5smv/f+el
Qu7XCxxnEcKVaIKBJ70VrzMSpDOwdPlPXsEnkokc/aAADt8jdayy5EZXL8qSpLlm
/cWTX//CIEUTF/NGpbJphIRCm7CLxIAKp2sAp833/eOWrBDE88iIbUtjALyYIO5e
2RhcQR2EfdEYVEpQtbR1sTcBDHhTmU3ANKtJ+ZaBFnKlGLB0LzCquM7hjxhUtAWV
j1buIZELIcJ8/QXYalIHXqxAgOXR3oot9oC9EbqHd1ytT50nrhh8i0gpCHk5/qEq
+PDLAjO/omB+pEd8wdF34a0XYW5lLMnY0BMPmIBYqWXakjztC8Oxuk2DVK9OJTfT
/ooVqEs+o9j8F8ATL0CQdYQzIdjVii4VdU/XYfVpQV1vOz2kgfGP4zYDsXsKmYTd
lkhJHbmLHSm3wgymjCT9oHleEnvE5TOFRNpXYH7sjCGqQ879hjJDKyRKPLt+tmUT
UmnLt9CbtWWTkVUK/UM1Xz7pTE2sLWQ+rUi3az8pTBm4tli//Dz748+2rXG11WXy
wH3s4wdpi3MpnAmJpW5h3xqyojR78SVeWPkBN4304A1czTn3kRt6QBYxcPCvVKFp
q0rpfZgO/DJkEO/VUP/8ipLAcMhEyLOClvnKq3YbFNUV6jFVPrtEQT8w9Znd16hZ
t5Tuqkb2cLOFlWkyn6f8GEu/Y61MnmPagTo4MKPnyE1pac9Cldmv0bGBtbLuBZfT
tWmVBQq9qUDA/gixb6TAxFRsk/jEY4fLs21F32a7sMWojpEoyh0Cc52HyeVa6DpN
qKjiNfCIaj78Tl4alLQLaY3qGZhDWIgFvqsoC2ls/nmyC1tq31+JR2oj7kKeIybm
8teu20lAZJgh7DrenbCwxml5B2rybBOkX/W5aCRrRqJLAHJ10h44bsI00d9nfuvl
bapeFlnUUdieEiVklPtODeq7F1yhfUM2Qs4Lt8xsPdPKzC5JiEmp1keglnQRVkgs
bF/USN0UjKjZyRJbSDBO6jGnt0pEpwPUV7ueeIpWkG+1K3Vsm+7D9GLKNHZSFHaQ
pfGFHm0DWK9lf2yYR/FQTSbmNzRnu3VOoj7QNz86GQhXA5ioyeUimonlbdlsN5Or
83o5Cq/EnyanVknbUgZVquGPbVVaFqnhLFxhYzS8tWgaqISV0t4ILh3JImwnaCQP
U/Dx+MlGuWe5xv+xX1OnbJrhmIdPR62zsS0cOmuQn/FFwKdMUOFQb8D6FVwAoXGF
bauX48a156oCYCliOaX/FVCPSjP6THX5/EwF1nFXNnGPNDxWGw2LzYL4xXTm2yrK
JjWxrnxG5lEYuJf6RDECZ+j9jT52CPJW7JswauGZdxknhmnvaJDCLrm5VwVbTR/f
N32RkHV2HpoZyvhGjGBlE/xMHRLQJwlXF4Wxvkpb4th8Y+8r8Jad9RGs6LgTvU3r
NLYF0zb26KAh2ceimO9ie6kmNRlUmFkEx8eiinyKKl/1jA9Vo936qgD6G3HY8Xmh
EkP+9DVvQCiWSw7gR03BDXIaTMkRyQlj1yB0U3++3MTEapjFxgBhAjKuaSnHzaxD
esCSGrPCNskCw7pq6GFJHHoDEeHHYzXhCp8B+pHkDqcCwCaT/UXLGfzqo3lJtXp1
NLX8gSfvR/ldkp3uFcofrFy9yvCkXMZTJpHjQrYx7ySim/exuC9WGU0Co4qj0jdH
aA3PcEiF0YREFh96bXHU+sguZ9vq10u9DTglqAOfSah1k3IVXkvBDGbaYCYlNXhT
u5+KS5Bz5zoUPKFTmfHHowEbDMNKZ4YNj+3IiVzxHNijGfnMBvs5rOM3GbKKmsXm
kKddL8Bf/a1ZbTYIVL96KnLxOOUvsFCxuNCGfUqyTvM2z9liYlEwo6BOMxsZEzKl
CSsJxyeJ9EcOACWTj4Yl8FOxW5Wq6xHSRFRoHwlg+W6+4qseR4RywGyW+7xEG75f
7mvVtnWsMPi0HIw851ofWqGfywgFZIL0lCNp9DEdQV3DpkmkbRG6f8zo9X9mXARi
tutO+iZETGEHqhKS24CqeDqd0zw9dS12oIkU1fhFfR4GHFmDz9ABaXTLwZU34ols
c+a3A7Fs0jUfpFZ20M/3kbqodQH0/IEWCd5qDblQNZMVymEfTdobgO3i4fTfIWk7
JXm/VQMXFO23WhEg8J7WOHDbXvf/755Qa/ImGRROKIUV8iUdkMmd8PDR6/CHOYP0
bV3inI5HEKwkKsDG1MeZUU4eTkAvSbNM9oiJpIDkjQsKdTvUhPqC3KIBj9gtoP2E
I5qUKjMJdaj9gQg/+pKQmAt6o6OoySWluGfmzd9zGEXxXMuZ5TFGIiqNLRXHJQ3t
EvrsAZZjH7+Xqj84MP11TtwdDvlu8WUXOau27Xm95qoMWmlfhsF4Yy2NBCSxq7iO
GuaB4tRJQDh2OQtiOTeLEDVHAxUqTkuLzIyFEtUPlXSPLy8rut6Zs53pku12YNF0
11WJGNYH4jxAz+ByS4n4lqU4dMYdh/8UIBY3ZR3WpYJXmPZNTfoExhutKdcebW2f
mKGFzWv8VxJ8LupGhS6Kf/8MDbPVzYVMVNFIJYVewPKh0USeFX5zU+GSxWJXcSPP
dtWo9vgb7ERjP6ixilmDiIfq8+ZCs+JisIdDdWFhfbub/9FKDT8sz8oYqtPW7p28
+nf9sqIWakbzAH+Nol+ukXwUGSZsq8npKjmVeeSzrNj+JhU3AXrFPN8A5UQLMggc
xFHvNILZuNqBqi6IcKoytTE1IwnSmAguzuE6Xysso7iFQXQ593vk3pvQBcgyBbnV
5eT1pl04cX54CAf4PDe2qj477sQifadqL5sgZuNqe2jRif3WwGVnmNKviQZMoGTs
LZOnvU0XJnFyn4qGSv73PgMgikoyVpe4LdM6iRaMac5bDq8jPBpLenb6tcbFcuV3
LdEgiPoaGNLC51TwRYEUO+wmDK/TQTbe9xQxVwv840ixM/ExJv2CKXIyKurYxKJi
Kf4Jcdw277ZyCi/UWelZ2/tINvUktoCrRuNSQ4Cgr+wK1v8fvNYxAWTlUUU/Ioqx
e99LSz6Fo42rK66zhF3WmVi7v9lAE5DxibA0IgSKLS86lg4ctproY2A8qeuFQwqG
PQ8RcPb4TnZslfk9qlYnx3RuxuuqSp/zOxFEvT4DxaMB2Hr3DPs/4MbILfRTSqXV
n6UeYk9lO0fU+PmduvbxyY/WxcKKGYZ3mD99Q7HCtJ07y5Hrr5LA+ZF1YvmW/mGc
RBttEQgWGYYSzSeYjTuHW4SRiiJdVJ9G+4uH9M3djahAWlHgyylg2lo6RA7Qod1N
oEe6/U+e61ErVruXG+wue0MPT1PD1MdMO3qMWS3VkCB6tSIn2g18yvik3MHkdCtG
3fu9IS/N/JEr8jgx1wxISNV02b0UsThnr8ZrbQDb9EZGxdeFlBi/KDMfkYaDQsl5
4AezCWKIwn38fNDPTC1kcJqAzN0XX1PsFCJhxxj7/lSp1aigcoOBAq6CN0QxTMx+
hXjnnIbGuuKJ8KHdWy6W7voB7kZk8pQMcW4VvTCKyNps7VMp2P6o3NvLpu2AOZXb
vW0EBUFjaV8sWoBS8rcNlpzJShaoCGyk6vEF9j5UlLKBlQgh7WmWhks/Ih4dd2Sb
+Ld1DYi1jEk7S1Lz/V0Xm1gdeB45OQcc3fl8NZdbOCmCkDNCGGNCeEi4qnUDjoVn
fGj4JZvv6QzHtg6iCrqJjhetINWfYJQ9CQHtmh8Q9o52QQBHTE8v4gn3fqh/0S1C
448+JzDGFRxKPYsXKuRHFHhu/q7RHdVZTMl+mi4Ync4HGwWuS1ilGJ3AU1vie7B0
C5JAXzKZtO3xLkdSmAlqeQEFXq4610fCwjnWXqwqIgwDS65zGU3M80nhRf1AHJ6L
raas3yqJgcXC1rwsPcy33Zujk1qhL9iqKtUMMiPwn9AO/cM4UX8vc7B3MlM0nJKi
3iPa0mX2wMTCaDlajpOOClu3v3tUmP9A44jOdCgF4kckychut03CBg3m/tdZUBJX
OVZnUnrXSRz4tB4lT0VcbXLGUGQFfBdzXSnKnHY9ZbxpmrGUC3JmdFbwmoq8J5c9
gbmugaLtu/CdzCiyDQWCkAIJ185U44TX5DrvSTixMf4FHOXauzpZJUwIbHzb8noS
0Rpy+CpRadMgSSmVNd1EdeEwf0ikMF+jlGukpPFNRtiOcyu/tGZZIsCFVewQZA7j
oULecbKfT9fF2b4E3kxC+iu8xGAd/4TRFBazWlgowSJf7TIZWIhAB8uyxfckc2Cn
1nUr+HjA3hhCcb9oCAlrPjnY2IEYLoIjdi6oTy0g1DItSnB8hAGmlalpUo1v+iKM
5Mx6lFLWNmRZr3Zky9JpfDFqRbYDIlJSDqyCgHBT2r80AF677UnRJYb1WhbTYP5U
TJzRYrrVkW4xOYnyc4mziwEOZ/eCP+SZJwnOYAlX6xjf77MkHBmHxpUlAXsAdecZ
NFKMN/lHCzDeMDDRaQPdsuHdjDjykDa63vHgeurFHLTV1aHSeGMNmMwsv7chcylN
2yKK6rYz/rDWfEz7N/PCTkMR225xy9QtnxXL3C3rp/JWRfHTx91r1M6DDAtGCPqJ
/PGuzfQzLdnxVImcKVgcBa0X9Zy9nKZZXz9D9KBU5Rp1MwvZ4m2pSU9I48fGuGp4
wLM7BISZbTuKmNSltBY+Pp7AkU4mucr++JM1hFhl/VD/ibMuhn2eHR2++ruWbpTd
9X7K8u3NbJ5z87e0LoyQWQ==
`protect END_PROTECTED
