`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wUfRcnbfmx+5UHprOAdITnw+RaRc05NJs1DuWAUaiX/fVU3vhlDoxnEoiMqPQnuw
rvWViARucUDiD/lNa1ICd+HdrfkmGo4zDOa2D5ernLjjbGRKZaXNqnxwZvRQL18Y
7juMb1WpFEDcUVodTv/QxN9YIChNS0M8ZS+Who/1W+wipapRlNljf2qleNh3pfdR
icnwFirwWgzaIOSS6Zk9KEADd806n7RHJmB+CGH5JGaxfiRIZiG3P3OGdzbQjZ8N
2a10AKFEIzxHGAi0Kr2rhGkE3bP6JfHoxlnPwFfskWhyy++YhCEASEZMfTBn5vwh
pytEkbtCv8MK86SbiE8xxNB+0qgIICZUQyaMetrP10JhFjRXQcj0W1oxErG21dZ4
QGqfwQR0wwfI4J3qMHa43Fd8yjRJaZKiC8C6+4V6asm+M152+KubZkL4DTNDb7g/
d7a/4yKDgDCESc4lbvieYY4UAfn89l8zYCAyfl3lGI2bCSi/uWeamgPs0Mk8TeDJ
zVlLg3NU0oCY9ex2aDxmlA==
`protect END_PROTECTED
