`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r/UZ3fGheSEmefpf+teUqRg65KoinXw9i9AA51OtJRwGPGz6plANSUcgD+GdKDCt
vNs7B2SK9lO9mitGD51Mc/Sp7/wLH1rqXc5nPwwA9x0tKagPH/SNNeXOEF16Kd5u
Q72eN0TpflqmQhv+HfH+90w3C6uxJh2HvWMwt3ethNqI5kp6kFxP/C44aHv/zgEw
/IoVnV8u4V1VIjOEGxz+Zuki4/4ZpQZ9m1k5+3odrRp0K0+cam4JNuFFvtzmApjg
CW+KS0I6+FwEtHts2lLj3WtrZMv03yVyGpiLuNzW4LH2xCuw3e1tlbyO0+botcKN
xfrjTSK7jPEA+CQ+yp+07uf+DrsGl9VP5a9Do1JpWfFUZq+fYg03rftxxSVEvF2G
q8lseYF5peIXUFTjk0Fclg7p7KGX5rAL7M7tj9r1q6KBWWrxDAVG7tLiKs+PsVBd
3rMEz25d9A9KKK913CWHYcJHUgNsbOCfR5QewjOQKCpLqvO3B2NhP5fslIJ+epv1
R1FQ8jQ70878DMl/qTLXnQpMslKfxSW2t3gyJV4SsDEvaeqK95FXVlY7RtBxlIPy
SCQAxZhvZRfi+VOXAg4wFCvKyqFaRH+sCcDTFKX6g9zNf2Sket8R5NumYGBXHFp2
W2bYKNDwxpH+U7V9nx5Zf/lU+kWwexOduthj5sMldY7GfsJe+C1ymSi3kSs6b61j
xtuBQNMW7M5sMX6eBTEgM1QBAjWYd/uZK3MtJqVcYKb8HtvgG3K35wrp4XKsDea6
2sMXuC7CAzThOk8Vxrj+KyuaPW7D6jdmhibqEByGDLLtsBFXZaRrndZJ1VhFmIny
CzoxsBRu3VzF3UpaZx4SNxl3FQt173NxVjh7BYqMIeJLl59iBLUbJCFI8WOl1Q+D
ZBE7Bmghx5ECo6IJLBPdVu+FyPjsHcY6SfIuj63nvqMEU2+b8XPEZcl2VyVir1mi
xJ6xixpYC8J9joU5O2BPliWWtWndBF2hHYdASsXHdhsGuFcHeBEWxHdGCC+l7PDV
DU41J6LWE3GamVC//LUyFooKpeYxGB4/ujjXDH+rfHb5q+AwHnYE5d34GQNslj8A
cJHX6ng9dgcjAYy+4y6dlINRK0sqGGXl7e+Xscb2ezbOca1ALjV/MRPB7Qo1rt0M
Q0PzMylaCHvMICmVUfFnCKSaYLCqZZ6naJNVygzH1+U72voBo2JxTGF7+doQWhvV
ULpGmJomrMxvkTn+mAqAH3IFaeyaqR8bPBW8aFSX5Ml5Fs/n5fozWEEqXObXVh6o
jrNGkBfI9WBD+oIvsoD31WUQuiRWl6HHvWY3M54bOQiofjZaskFnQx8q5KhCdFw2
vtTPdqtadZ9A5t0zoiQeA7+7BAFyOLXiUlaOHzmjh2CVZqgbOhuYONShM7ZATcyI
wVFR8sHffQtXhxaxHo8ZLHNB7PvYcsyrMN+f0LjjjwNnGKujoCLOQBMhNg7LseYu
BM3sUBvIkv9c686KRVKZf0WkIkFfJwvmt83PwONnPCA261dpsV/gD1nCjfCwY9O6
7hhHMqpiBMn4as6AnU+tma2wxn/rHAnKLA1hbUuZELI0ZheZ7qDAvZQjCakYFXyq
xmnuRb7DxkWPiRt8L8FNSUsY2Bj1XNJHCcc1MV9VsROAZJHudpo/Ss7NWGBAyuLl
xc757rw8JK6WnW1LLVDwKj5ekBzTJm/Vzv78ABythxNAWQWx8krpMOcD7TMD/Ly5
HvOOgB5EmfmVTr71FNJnOvSJrG1wOufs88L9QQH/uwWxUk+ljUxv434x8gQU8Nl9
UY8PobJ9MPggi4WKmn+uIDFzb+qIXUGXg7B9wZDnEEIB692gaKBBgNZTWb59l2mk
8DkHrehO0q8QVfBcF6kNinje2k5vUP7nQA9wURIo077cZ75hYI7XKDKEKjnwgBVa
Z48zit3jyRWHUA3dirmc22X51BmGrpt5xJ9oB3avRR49X58ZunowQ9bdYxJqvamZ
YF2Ay97rpNcWIVtrE4BntRDFIqTR1e9RdmaK4QS3Xx5tCrfBaar+hdDKftOTQdXZ
f9urOEY4mjMGCNrqFprZakTEhYaVO00xaP7svrOIM3qPjSXx8uerFYmAS4KG1DVo
XsK2MM9bjTqNJ2M2jRuTBYKlJ91l+1IW8IRdPTRjpbFkDMs/DV0s5bpCc6dAnGQw
dQynHDzUvZkBlUSxffOUFjfxRhhKbB/eNCSOF7YfHEkgQ3xyUgN16jKV8Yy2qxxJ
x4dLcv4lgHp+X+t8F9XPpAafidVG9MoSgfGxvPf5cJgXnzRZ0WkFmJbCB6aGExcx
56eKFOW+lGZDctto6YJ/lQqgUqkPWZOeHUEj/jFCA0jrgjOcYYfIJ2ZTq6SH0zgC
Nk4KyceOGJdYKr7xuN2nfTLODWonCcJf327IVfkLdHZFEHhbf3Q7W8k23r8GmY4Z
fxRhSw73HZbAOlfZwWoZR1wa/jAjzRl/RWUZuP5NShwWYgZWKQYIIhXpJV3BpLVT
ufQKYPuTNbA5ZdWVF4a9y7GE43G1vzVakFggZq3x9q8poGIQPKfMN2ha3VKdqRAO
NPJ13lqENjOMMMsAcTmN6hp35PczOo0KnYk8yS+TUEUGEQ6JiGOhzfrxjm6pL9Lp
K6zJCWO++9ytbVI6NIrRYAVQKF9MrhwBhgiu+ZIi9FIEbVp90xO+UFSo5Ax2bm/7
g+WfW5mcvFJpOlFWlQQ3ZmBpTRSQFS4fyfY2YWr+/uMpvUw8xLOOdaNBdte4iF0w
gDwQOSDOMfYA4Ur64YlrC7oHKlXfAklcp3gNleZy9inmLQm11/yk+ZukJZeWRnfH
k/x+4k1qFirE2CnvC6GzWFFleX4Lu4Te3W5V/g24jX2LGScsEzV3gCnTT6E8aK2a
5WY2MruYczNjYYDtAQ8RraYxF23/EPUkcanmr2xNfgl4PYhpK2i0goyYo1aG/SzU
aKpeaKWNyqkDmIP/75cnZpGOQAKsrw4gJ0CrvwBL+RmSQlgy9CH7AelkMBw4joDK
B7p/3u4764N9GWC80f1fr5jAMrSVXGDL0STM7TfHzSKMqlT6Sbi/HoeKiCWmohiu
CzjcsHNuyC2CsljI+UQTIF5YGqKSQ+hF1ZhVvg0CqwHkUU0bAYT0NjRr7SRwUoCV
nDeDg5BRe0yT/0zczy0mu6gtbrvX9d2/AB9jjgIpPtzoKeCicJ7LzR6tdWXraoVX
SFmYPddQoB7I+YCopXdwslhsOp5tpKGWp7UWAYp8rrNTatrznLXnMbQ46ApYHUEn
ATwVKTQgsLjfjlzIJmOgAH6WxM2soSkpMEQtgHVSSyXak+QREXmqsSSAtQV/CLrJ
lw9O7HwG+vqwhyDHTo2HVmf9rv7GKLROM5ldepBqDqujgm5ogN39x0khridmecg/
T/oCzPgvecYt0/6G8WMToKlIz5MU06/4iVbz4oLl0G+YPrD613gg0BefErR4TYgc
dimfOmWYWkF0yBJbPgQ1cQIt9fo6jcqDGVT1NuWBBz1poTiKZRKx2iNFzDVhoIIr
9Ndoya4vF2upeXsz/ghE6Qp2IrSLrg8fvdGwRAVYP2vVqNoMagVf+HB3ztFwaifk
PPdkBdTgQ7EBV7xO4SV2vRnape3B3Dol3MCcef6dTODBEDOrYomRh0XxbNKoHLwv
8dOR0tghIGbdsXOCkg5KtrnPx0iBAQ61jd44dXN1ZxDpVK6w4JFuLbrAlk8JbElr
N6w7TQZt7D3FF16NfdV8oIuVpr7+nXJP33BFcvBuxeZqgh9lXHk4V1aS+nkfUG6W
YAUoIWiLU/dACkT5t1TtuAMdq4W7K4VDbYTQublBln5z+iZfszrdCr0q1hkSaZC3
BzT6qzKLp9L4C5BC7JPSZqxZ28Br+WqzDPBKRPngcIXXhTwiTg8YO/rFY2js/7wA
gbJgsOBXeKhk+SrxEQWmGi9ma8LiO1HQLXOKWulM4G7xypHrHzQJLGlcklS4aE/R
Qhn/LyaztctqZ8ipKGxWssidL5fcZoPQeXwUUfveaFJpeXYJxozBH1Seu7DCD8R4
L/r+7+OsuTRGO01+jPaUPEChNJ1TdJCYH4pL9hVPeRXVlWmoU/R5v22IyG4dmgc+
2jpk42Z1StEUW9MJOXq+NiGvJ6DwcaOkKz3wcKEmw3+1UPVKZqzseRHPp6dNlJr9
SYRPqL26OGO9a4NILq+I1Vo7SbIGggc2GLi4hQeimjbKWT35XZ1qU/pue89EOOan
XaPV8UPFAy4H7h8OgvsXuRdHEVfPp8AsdMlUeJPCku8Ch3SeZ/YuNkdX/t68d+Eu
GFOexleNs3u+EJJcqYEo5dlgXsdFd/V2WNdOa03R4RlSVTwfqOdcB1hZ/n4DxhaF
nf5TWVy6KR89Jcr1743On91Rb0mhLvTegnQtVkGS++jvNFvyIx/eD3DRloSGWu6t
2D/SxPCfSca1/gl9rBKwQpdxR2LUKjbZXxBYicd8+INolsDuerMv+//rez5ROa9d
xj3ba3WoyFbn66P+zxWOGv+dewAuptirgLEk2Yn30N6WIO9R5PtWRAMR0lV73s39
Y7WGDg3y+npGOESzfbJfMhYfeELHFK5+frOog4zk7cGjCIY2sOUwQvEeUCa0bGqj
8Aj3BT9loRozx7g1pumA7jytntDyV/qQGKx5RR+SsD4SHX2vaiLYAxYJRgaJIBZb
wSXIcoTinLKtL8s3D2vMC2Ewzm/RSc/fz9i806gN+lA9xciqB19LXolsr2Su7+Hm
6W5JW9S9fKZ/POsFXd28TEFJNNSmE1ZatRqMdwiBux0ac/jMSKW1j0otk06c4RYT
LYENc8ZJqsMDdCvlQO8L77UpEMuFjP3qZ1wiHm12YJM1w8jJG1jnzdMGORYezDya
wP3Xm9p5Tz6ZTzd8PiZQqe3by1r7War2iPuoLqWcYWEmHeGE5KXBJajV2yT59ZYA
Y3ZpytwjEeaoMx/LGquMCd7cT3i5MxrDUYu28tfVrGtzjZwh2XI70HRcXloQ8k7q
jlZjzEJSsk1ThVrC4lPUWe4X/vcDmkh4VYWQrMi24RxmPLT3/G+I1o8AqUVofUfM
R1Qp3ZWWmUl/JJ6IqSZeGy8oSDGuEa61Nf5tOzerPrDoZgxQzomw9JkfOpi1y8aG
P3zCXtZTNmMJFdgkxZGYvXF31/+nJQDuGd0T8uZdDolT0DMuMMcC/2fwWhxwR/r6
+Xp2PRYE3jQ8G0WwnHe89V08ymsABYHRs4C3ekTlXQSP4w2JUaCnsi5I6jXiuRv1
g72m61vh1xvMb9bY8QxgLPL7hV22KgLMtZ/v6x8/k6fyRAXGGLwMwhQCqMSZitOw
4yxh69ZpkOGndE9a/bMs8efJlzlv7pbSyY0jgsknNWOtpx+5pD1avCIOOHoJ3GhN
sr1uIO3sG2UeCAuO5EknMNB/Nkql/4nTdkeLdO6NWG46BisTH5vIb6JY9xvwqsZp
sBLuy62BMnVxC5lgM+RBzwHQMYpC3/nRz2t6MWQStHcZMAevwQu9vxBkDelmfOE7
0XXvAOv5UpBeNtmwfpw2D7uPTC1R8O/3SZBTQmee4qRER0zTopo6TJ9LRL+8ukht
o6E9uQc40HCQKnFLAjDdLR6W/0Fal3R+iUa39IgGTxXQsBbrBvGrVOTogC/WxFnK
BueWzpCwMM1a/AAy43ML6pE8bML1u9IDV0z0GjYxPsa0qJYsRE4YfJcuemClMlvs
ig48eo75dcJsE5fBIOMgm7/4auVB15kH+Ao5XPfWH6ruY8HFVX9S/dkJyzLdz/aN
B0PR5WXWJFgSdrXp7XLxlg/lvfwqqPVUxkctispr32F/GUtn8JzWX5zWwFN76KdV
7QCMQs62gc6HfnKIXK/bbSHYp32CJwC+t7ZMz8SD4KzjzerBagN47FkWPORmM1r6
cVvjvIPYbQv4ttcx7ZQ2P0yzcBjTexC9guzGV8DMg5BF1aE/DlvdtkYJtgp8h0ys
CT/BjQKQwnxcjBNRyYvKSFu18gYrtLG74arNc107xPmEycBSPAj2uHwv/VqdhreD
ITrU4PfrEX91+I6P/QKLSV2GvDTQIQ//M+Fd7cUPb4dtS4M+94/0DW6/hwSgGZN6
SeaofBlN7+JJHJK+rG00dfq6MxUspBITUMIgQT6Xq93eQSw3m+BhRe1GbDCN58u2
6ZMqXmeQJJYLEcMz9qleJvh++S3F3t+9iVjKsFgWHG4LKjnQ6QG5mHHFhBIAjhcW
M3fHx7v3/rC4h/5bEVJYxitW1PDJXHSTqwDHLrk0edl+dACrnuPBLdRxfxHFzORK
zXlF25wVBngpPBRFTQ5DkrNg7MLLp4dRO4PGyVsawtM1O+oQlGpy9oFMdBy4ojL2
d1tbWIhUv7raF1SyWyU3bJxm7dkSairrj/xoFMKQk//qLipAeuHU0zlRD1OxJ/1w
czRQJ+H9CeehkxptR95N4ffwOsElY2YDKXpg8lQ7Q14kdn8vciHt7xUlocjG3MBo
+zq2rHi0evkY2V1k1nFDxiV0mZ4KTibKEeplj3LeBl4bIkG8cdHlYdxx4npn2L8L
WkPeyUhO8EBH6mPv4r+74R3u9r71LrLQn+3eH7GQpzlXE747WpOkGM4Tu+kYg3Ta
hgFkNV8OwYfkF5Cz2eqr2IRq0QlO3OwrjnnEfMM7MUBNUokrq2HQ1OFKSZlkZ/B/
McQTPgBlcBQU1pqMcEE9cFi9X5y/SzqF46Sp4WpovFjeRU6LvOc6k37/ET17cglU
0r2/EkiBJAB24WeFdKVgy9AbjNJboL1Hgt6i000ORxXIjR1mYSRuxhE2QaqJIKEA
R2dedxmw87is0pY4peAZT6pAJTIzr+Z9Cj0Tu2q5uyuBeUxJNX8wDMouA356eF7Q
MjT4Y6bsoWKqR/c8XXwU23pJeLTA59v63PlW3eDyapQwLhYuscp7LdZp/TRWK+mE
Sq/ofCQ1PlLQUjeOaQlxwSGR3NIMDRWnuMZzPLMjDrIotj6am8EOlbvpxGpWWTHv
jfyUBy+evsyxfSBuESLjz2RwtX8Jhz4BvpzZuy/y4Pz6aAyVc+TNk/FbTw2OdrF3
WAvRimZTf/xFZMd3jCBq5ZhGpj21jKhrA3mNriaYUX2dwS3Taf7pyYXCNx/EQrPQ
HDwJDu6LaAAxKqqZ7v+uE8otFaFL+orI7FKiGO+E5evfHnNvDCHZWnBPYBdT1roh
EJlZPAjuqU5pZlbJFmPpew/PtnI5/hSdc9Z7o2zqxpgiZlFiiECJlG8p1b9ts1+E
FQoDQkYqroVNK38364xJb/rXOpOMlDk4KLoi08oOXlsCgSlTNuXxQah3LDge6pwd
h1I18A6rEv86w6wNqLEOnIv6pSgDmMD/DteBnUQsRUy2ZEVcifbLITykHdumUpav
26MY7edlpytkWYqIVWrqYmvhs5UAAv1NqciEprW5PWhw5sQJPCqWTL+a/CiWznp5
b9YLcorDg8Ui/lqfpQ+L3MIoEf077/lubggzHNBJi3x/OvgbsjhZ60Xb+yEKk6iY
9QFAkAa/Y1YC1NPPBuW1XbSuv2sgSFQhledC2HVmX+wRlEe56GmaFe+zdgW2yMHk
bfKswS5igNmkjbSYIykNtE2VPgPZoaG0T7sH9k4fqxlQLop4Gtq4d4mp2ib30T70
WJVUYvVHhUts8hOBMEIGIAjIxODjLEjIbekD9/URd63Pp3sHK/l2EoUExuBy8vam
R/opqYXufoJ9CrarBmArH/B2g7IcldzApf3RsWgphqK28lU5go6I950xisQataVN
wWQCXQ7bR66mILaZ5TftNvKKoNHr9B3Zms727W2IufKV9xJ9myPS8Rk8VxzJ0N4a
IUj7LQd4ROfR6ntYvk24KUpQqODS/Yu6Xz3iF/A8nf0j0p15yMkw1NubWFu2BhTD
bEXnyMxQut1XwDT9/uopxGVQ25f16xBsriYCT5fLvQ0RLBzHSJTD+7kcVr+6Dlln
OaqfJJ1HDCblXYSBWa9htNmMGHWtn84wUtV0Qit7JY61Ish692gsdkwpDbOCSl0U
SQpxj6C9QgKVkp9x7rBvv3h6EHAxEOPL1dRTAWcmW76M18v9jLbqAlTOXyuhHxZj
8TWE0sAOUTWss8XCtpzx/6z4LmTBMqKV65m7Y7y/aRB8YvBRDZLO54/MWdvlFlOz
PBPhESq3IsqropU3IpT4YWZQsVTIFWddQ+d3auTkK7t44WMZrazhU0UBok+Y3mCa
N6OjCKEsSuq+kV2myGED5gh3uqll3tSzgv89D8TbohCe4z7cA07fZcYqIOJ9aWtl
7RrOLO3IkZ/2LzIxB0Y4QVND82A3qKeNG8ExcnnxVxvbj1EW5TSO3ehXi/AXAPxG
ne8J7CeMmlPBzIbMzjP42qpXdkzVOiA30wzLOVndDwwIeR5of9uFaoWGt7ca6xsp
nLiovxwaPlJAzObnS8Q7IcBsaKwS6Pad4i1npv9iYPjyrImqdlJoVaYnspSGlPkK
Eg8DbB09eCjKav1/QUfA86FmZP/zT3fdpdZQvPHvLIYyImZEVHvy0gsdEeXxqIei
guHiQVs2Bz1ls1T/fAVnNbpSunvWvCbdFfUX/bTWH6nbOyna7AvQnoO8PUkaGSI+
/7Ex7KNNWtZzH6qnpDfytcCAH7yTG+Tyu/PrzPyyo2suXU1I4DnNUmqtM5XOUxCo
7hrmUEiyx0T0/k63xf133+YYaD283xH3V3gWWqzN3UCWkPvj03CBWGxb3h7hvMow
IdeElwdVIkB6/l8OBvXWJsd5g7Hqy+1hxWBZfGUHM3cdWPzTDiapUTh3ivwK0uSy
8bCDUfQAn8jsifcD+zVS8SDrWI5icR6yd/3eUqmsBmfKEkayV8E6gbX31sWHNTyz
J+aqZYvY0ZdYVi2rNdDb4O3NXrOs38pJulktjxJVa+P9My7eP3CAoyCuAW4aVzPz
lkLpj0xy3QvRIjG++C8QtKPD2Vwv0jLle4e7r7djUPueUgzkvxvRIzCAiDmdPX+l
1+2Z4Pm0QZyi/0qBmfaG4v4F9H3aVuE6DZeORNSlSrNz+cO3Bmf5Hkj384zc3laX
MeMPsKXjhBnudybMA6KCCwuVahyDF6WSiZUktlhM8ZO7edUozd115MGN54eHE5SB
dkCjhR5Lp8LvVZL+xj8FsJKJN1Pi6BgEFyJw8p6kp1vKAUvwQQa/5R4sWMzIyxo0
KcY/SA3YBCgrAwMLA1WO3HhBwOEVXVpTojn1t8xhK6x5Zl0PS1B/jRyLBHE+T8hG
kFAh7+ZK75KRkLtP7/JeBTGD3FxTgCY3P17t3qIX659+HtEvzFHXzeTTZHlwMObr
8NsmVG4dCPCuB0YutNusPtA5x0m0G54r0OSe6k3CcOhuWhZWdnlw28qZd6hJLQ+P
ylhx5lwxmo5xCSsQiqPh0sTWA9SL3KPlmFJi6+duCw5DEW5HvWqPdzj6zj8RHieF
J6QOv5EZdGPh5+dEWWeNHOs5IX8dbeVNMogPQRfPfFOlyDCIn1zOGe4tEzFFFk3E
dLLZJ361mB7WEOLUeOcUw2bLqoEI7gucR06tdthlTYVDYzAAFuUTT1oWzZA3BXn1
C+zMKciz93tllY/1oProZBkpCeYCdYEO1Jlozp+nPnCasiFVltsFJQDjFjgfc3p1
sqmGFps+ZjemgI2vFTzvW0EcN3dv4haPQhXAFA5sgolNKv6w4RPUFt/xdEMyOsge
XpyUKxmjLgTvFNREREAAtOePvVrwpkQX1lIJb0tnK+ceCs3k7ydMXo3YOh7JyBYR
o/rHJL13a51dInoZrOB4CXqDET9jsm3S68RpoSdeLDYxdvyjt/PPwdYlH9gAE7V1
66P9Q3Y0c3BaxRHzB1DW1nVcmuUv/7D46MtgMk1ohK8ZnDnCZjGlKVsYmLBwY2B4
F7b7QA+GP/EQwPeGilmE8UqKt2L+iF/gj2fgPGpWufUyNJGSiQVWDwIk68/ky+2/
chsPCkMSpD4rCwxnV7v5jRpdsV1gkw8N78wm4L3Ge2iEwqgcAVyN8dnoFrnIW36A
UMZ4Axx26sXSiV224rpjJNXmMA9ymy8j3NYC01+my88vkHhXFk6c950vpY1F/Hd6
Z5Ai4icWNd4dqOsL6dMRS5ll9c7uFsmJ6wz+PcTtWf4RShCHZvIWEt4NNnewGUmi
Wm2iA6yyP1LgryStZGimEU6wSJk9y2j+f+igVWlrQGJgTaTzLDZObL4F4vYb7FI6
v0khWhqloxFAX3uzGA1LgYckK5KfOFubyuJi95G55xC6RXvjr8kJ4pSNHtm4cAPi
QE+im35C+kDmdBZT4ffNAi++DByi4sQq//DD7JBtxQpp4QH9npS8RHgRy3NGQVvN
y/eLwd1YepD037LHIY2bi1GVohmcVz4QK6N0vNzzFSiaDBqeyB1HkQF64LIA2lYB
hik3AL2dBzaJ+JFyV7HcpXP5qq4hXp0L5Be/LkchCoRiF2SvFZsSEZBL8JOTGKpt
C9tU+6qwS6sEZY4nrlehWl/E+eHA4MpfB0YOE7+Y4IZUKwEeS3NTlRWXX72n/ZyI
hpZWcWMDmx3RICWe5yLfcpRuyepxIAV4QntnSrbs0fNVV2ylbr7bifEMkxhb3gf2
HozsI/XhtX56eof/IVrpj7sPFzBC0YoHFZxiUOplsST+7AI92c4NvC7uMymYabcH
ngauOCZOZM+MmheSkk3jEVnhiIUTrMFEoscwx3SCRX3o/JTDIMmODbcttR76ltnc
RiJJj2dAJCS1To1Mbfmz83tbXGcEXPmPbSTAk4Rbzvw/tumUZzH8wq5UsN2Uz3Q2
Ou/nNgoeEQjSeWGzukrVfIClByts1p5O28xcdIOdxy62u2bLQE+So3xvT0LIYxIj
nBFWE1dDYPacWzh0zQjbuESLtCOzuEQ6qx19WtYJzmrH4Pvgyk3fn1Qe/OKJe7n8
8Mw0Jg6K1GclFDYZcwCjy1n3OiXNkVcuv6BfJywxDK+S899lyO2Z/Qb9F77oe9w2
95eRX5stKoj+cGi2pK3umd8skHZoYag6Kxqy0iP+re1i22gcJTCaugvkHb38necz
nMibq6dtQAOHRnZ9yBYcqbxgbpQIGAkSvSXty4dqyZbN6Q9GrPdFXvCqgKMAOP5S
5I9uk+rplrhK34zlHLZvrUr1HGVhAHF7/LNwEFy2PiL9DSstyQ3K7cl5WM0hLMaw
FmkhzP4N5Bjo8O/92IhnptbyVag3JZFpD4AvekdwSVcLHPBX3jo6HehAFSb456KL
xUU9Sf4Ii1x+7sB2U797Z83dufeMoRPQ6Kz667xb0DeBkx4uSPq7GhUmNkH945kC
o4bVsi3FMMO9Zd1gYsRCKFk2KgnkzgoEnAQyCy+V+VbyiNOhPMLZlphbVqS4/tnf
5wWakkjMBuY5lJc0QVKEDtJtQPCKYAwVvdwU5zSnFhaXlQ+fnNE9DBo3px3CjLND
jX+ylOI/6KnM5601MPUsoNupPVzUDDJ1qLg0VadszXuoMEccKDWJsqQ15kG8ulZG
ia1hbJ52Wo/SjyIeEmNiaWvQ5IivpgYa0YA70E92Jz9Li47G4nlhO0409JwgucI+
Ez074ovb2Uzcy/Z0qz+5LvHxDf9LWevnLEhrUIFxbk8Zk9sNamHX4CDQjpQ7Go7f
w+0QAVhxGqG/ULO+zGjSNnujC2QxOpnE0yL+bneb46K4cbtO+m5Pb5bHsgykPZCw
rVfnc6tViZlt70vJ3SocmblSQzE1ovsa6Ca7lWXT+/Thw5jvbYHti+Jf9dO3y9+Q
6O/F6Kx8XhJ4QH3xU/axkN1SXlvLRAM6S/Q694+aIKFEyhx7GHZrs3eLgCSFW/Q4
G4OCfTXUVp4l9jSaMn9G6ijWzb6MA7COO7wuwJvbGDST+USh7KKPIunDZ2ApY0bq
uYfDYAaQA0XbPwTgxSnknL8xTChf0Gp4Yg6fnYgq8aSjWnbQbC/Jc7SlYs9BjOkm
OtdP37RPbpRMEdhrNPCMNHsVG/6ekukidN869FhCdViidP5dbhOzlAyZO/E8lMhM
LfI44Lb+s1VriS09rewUhVV/Su4bAnW4L1twDmp1zHnsobYWDcHdzLgieBkoNHnP
/vWbT3Id4laSx89gtzmIA5G0Nnb1Msqpdi0jyRqTbEUpuPuI8hqZYYHx/hFmIQu8
wEFkpEXfoPnxXtmDns0jMmNdn1zEVj5k/ufA+gfJvTnb4SOXlmXj76ac9D//44Nf
BJxoIVyNd48c6d6ZcaODHo8P+TUx1FtmicKFaRIuibjvuQYvIqY929iR8kUiphFP
2vGd9htZW9oMSgOn+FR6r0fWdUQiWAlmuV10KJ4MIRWBp30BKTq8jz5ZjXh4BHz0
+B5zqPdaCWxwCUnKmMYXsNPKOoqXkKUZFfn1iJXP7vv+T1LOZZVGXOJW4hJOlc+j
JS5rQTVOhff/3kUj09UsYpiqmNFJDqI5hG/0mnpif4KVPxk4Z61Yh3zw44XW2JXG
w/2EXGKNJRQyQzPSmT1JsXdDhyrJ9vzq8jTuIcCPDUsMfq0cR0GMYlazNoi7igMG
3X88LTJFXXZRHfXVCJWLHgy5mJxDH4kUpWpREbrs26dZikBfQXfvb2A6OplT+9JR
06c37VkQSZ8ZRtqhJPdbMhaE/B5EiM1UqPpJ50S62OoYKAi5Af2aICaj3E+CENIg
ay4W3qLUQeLZN4u5T2jxqcYyMgQCH/SIHC0YCxMSjbtysRWcv0Jjae57259IwLPW
muNoKhsnLfhOWBhgnUUdimq76zDcFY2Vh9YShdpYfgFF4zfBkb9aS8Jl4TMj0z4T
hSRirB6cBuUFeOEvo3IoiBl4reZ2MwxpbD0Q3rufxjhu+zvyMc3Aa6kamuFuno6v
7LKyDhQn2S9VWyAjwG95e5Gyq/dr84mwB8aQOqFWRWDLqkeuDrZJYyDNsiViHXe+
SRBP9scxZkBYSGC60WozV7f0yZiZ/wGQNR3xz4ySzIYxXMAPTPUR9bHak1iLl9EQ
pwajXqjSXxEtW+3ihiw1fRYDrw++2bfr2UFhRFvUTsW3xWQ7yaAtDoSBtxk5Kedf
rNCXxvyN3er8oeetBi1z7Vf/xzGvzszqxBKHwp2qPlE39g0Bk9HkIQwEYv9AIA5R
mWHrY8A8Xf0AzBbcPxnx0SZfzRrgOxV+ZYbXNsOVbzpyRC86ls2ygmJNO+XzOdrD
LKslS4Dpi0d234AhDMUEquf/B+OycRzqan3iRa3DxChtXJhsZEFt9Bo5q2K6vF6A
ZhelZWIjz3HO1peD5gPhb2aK+3/2Etv1FdhaVuvPMO1IMXG3411h4hxJWzJ/OhgO
hdhSl/IziE9FJCGawBC9YYfvhyTaqjqqg3/YPWw8gWwOwpC6iCI5tLIyy1pLdg4V
+ComB89SpGdoXsuwGO6lNzcwQ6YGFtpszGb9nIKaQVHczjoxTOeFQ3sWiIJSOvvU
ru/z1RBFiBGWErcAEOGw4uQkcnK7of8TNBDBqegtxNt7K0T5saGo1qazMRJ1kUe2
qHh/kvW7eApNLZCZM5m4u6eKHKoogFFEGSEVGqL7TqEocsDhEuQRFMCX5pJHcESe
4gsMWSTULPAKZ3IvUfJefc3ZSlFwdh785X7w5S+HY+12LGYb2kD6dCyKYJpLy6+e
2xHcC1AjFysKBXCGbULkEnos5tu8e+aIdt1pYQO20RSGTZw1tLAum5IChuYjyD2l
IS8BvOPjdeVxreSUNOrld9W4D94K3t4DtRrD2VZEitnNDCT4BXhn2ZkSFRbpc3x7
vXRuodhrJMsO3vJZLnLCOq4jlgfW2U2EGkVoQ8D5fV+2VXg1jlwJYomUOK4YyMZ+
Gclhmp8EpO4Ad1Nw/ABZN3lR6mRBKOrKH2a5seLjXD3HDZHy//YVQr5EEIwiXhHR
Y0PA6WnhEkeo5qUz+Z2hcZkR/mGA7linsYn00YtDlf6/KIOIRej/umlXi23xA3Ze
MzVEiWvM1i8s99Fgg4GMCC+nPegwrSxCQSCJsyCw8prvJGe213b4YGmQz/z60dMd
Hw1zjb30voILdg7CTqclQOxRmJfqI6PfpVEOdwVPl0Tg0kKeRt3h7o0g/92rv90M
BiLe4ldyQZ7vA9SNzfzpXCKDycWeXnHYdJamGXfkPO8VZv6V8Fpz0a+ALyLxHW67
6RbHWLgH75UpjRcq0YQmsfofB9QMZ1093SsdN0OfiBVXqFPuqDwkzTM8attzqaAR
v+NyEJ1hhTd9C0pCmqspTguF1nFjCbGWTs1aMEiVGU/+/vSAQ96gSg+L4e3FNbpO
hjZigJ5ttQWjzaFm+Y+ucbxfGOsMNighTQBt+WJ1bciVtzEWfzPvgPSz/CwsqF5Z
ToOq1QIjPaDGTy6FbOjttVdAhf2AoThymUsDcf1Sw6lk3orDtZ185u4btfMr6Oci
Q+zS4Da8OZK5J16N607i1pwNsH6+HMXU4bQV4fI0cQhRSezBOmBpsPSvDDiRRb9l
YV1VHQkZsqUoqFb1i70+cKajAfeveIiuC339Fy2tlqz/ho86FFHuTRaLQlVf8Gf9
3nEaLk66lucq5CNJhgT8Mp8L9++JdXT0KQQei5jd6dNaCRVRCD/hhehskQWGAH7r
yTnClxqyDBH64FJqfpUmEdTEOlXeRCQV2GoHbRh322c6YK6xdaxcZCl7oMqgPZ2G
2ocTtXfCdPe8T9cNCf+sej6IRZkV6s+yDnrtVoard0kdwDU/ZjXiaElFgczNW+97
6MgkluD2Z2tuXxeeaQVUtIxJ0Ste15WiQ7EEmwle7pUaqdQU/aAZ5OEsc18kWn5L
ZsJ8/nQLjfF9dxPVchJSRQizdc8Gr3padg0l7YMrDP4B06ZIofVa9HwRrz7bNEdK
AIZzFvHRtILRSbJfEi2OnXB//i0gM59QQHYNJcIahkq5FC54AEQbXtVO1glMlDJK
22G5qdihikxNX72hep4fJrIkL6omV3+ksKMfdjcAMa+jz4NQ4WWou0BECP2fpqtx
gm5aCrB1qi3axG1hYrKWPLxDdQyjsRdRwSI4BjhM/xMfzFBXMW4SBsSaaUw5dDxf
HZSTpi+6PA+fNsKYqDcJAfSg2z1L+tGGEqI+o91YF1G4Hgajv/qIu4R9tYMDIkpB
c2pkYL830Ju+2IjRaWtxK8IYqtNnq0fFxeLhP4atsQK/iHHM3lJD73v5EMqvZo3N
rQMXKumKAYNY5O+Zu1jBwYaN+bOSpWgBLPMrUQOjVpYBAyGddUu+MTm6XSeXnfwp
xUzIJrzuewQegWNdCaSO5+7+51hPxphAI1bASTXlFQ6bIponOTmU+ycZOokcaFvu
jhx3NjM7tTPNOXCJDEAt1JFbgkr9M3nmksRI+tMFsQLWoy0+LNTrCM2GoiDNYLVV
7Qn2MrEaV2IXgftnJLDgHWkpruCRCSfg0G3qNoXqYkfpxnK6aVvjli2teGoXEUuf
CUb3x7ENXG+T7yADH7iX1qA9Q4cjVY4v+mQkGpRzI+f3MFQx8GP0xkYwMz228r5A
WNTIPpNAkstY+0PGL7JYHJke7Uff17Cr0YARukt2zrhCQ4Na+DK9QMA2dkVggGKC
jzIdBG6n7WJjG+X7G9l10tZeZIF5BVQwrAkwNHnE1AVTkgnh0eqbel/fcJMFPM+2
GJpkagR874IY6c9ySQMK5D5leD/EaoRPqNfgF7Rfz4oyW5FIZTIiqPZIcuafC/lK
Bs59iK31O2pwIhgz4YUcmXfW8pqXXcadNAoVFk/FXByHpv7oRlHbm8aRgrcJTpa5
lIHEOJ4aOpr7C25iWdx8jOGSV5DF7v8ZZ17MrfJ/yDq56MmEBuZJr5SKlwebjhDb
3HpOB+W0UJ39QLJ0ksKyj01hzxTFm+2tseWeSFMmTDCBx+xoNpNy5rrnKzW4NfaZ
ReUi2tOlDCz+ybao5W8Vb1RztrzWtifiuVwuM0ec4NzTj43nyJ4DiLVYFtx6oVAH
FTIEvWWkIzi41D0r7V7Vv8Kf5plaE9h8sT43X+zPWmeHtWaBDKlvB9pnmIVktMsC
rC2/Hgc1Itk28JS0TkBmcpVV+pv7S1/sASzx8z/eAlrq8LzhTyMY8ecmp5oBGx13
AOJXgSPpHNe/rxf6vPrpOkiZjwUxrYdZrgwPvXKVYL9TMO1YDNR5KwJ7nBCrkfqF
mygL2zBpcGg/OysvWRMrEVEJv+q4MgsiwhHhFT/DsxDC8gBXONJCa4sikavWfYTl
UzaU7EHZcH+PWlhW7rIZtb3HVZs3UEcFBx2YyENfpkKWnAJb/uD4926l6IYRUirX
uM/Cku5y3Jl+kZbOlbDkGI8CZh+07pIby6JNSmrIlWQ0ZNZLinJGlRFZkDU4z4DL
7SV9jaMHpTr7QHhD6nOquB6GWz1a/XHfoiO6n7Vl9VIPu0hMG6IwIfTZrWAcAE9c
ZfM15NrypIH64xIzY3m8CEVP5GGdd81ABj5b0lQgfcUyflqCyzvkVvgVaJGYfbGB
YG0cZSSwtshYXmE4FQqQSvPgZjE+tDvChg4KnNDSXbxXnMujVW/AuxS9Skzjt7ba
cV3IQOk/Lxd+phGCF1EQ/mnpUiEFZf0JdpwQLSycCwbA4MYUxCa/cn6MvNRQSUg5
Z2v18DfjvjBKVRjBOz7DRgCUIkbljH6D5Mz1CJ2Ka4qBSNA/zS/BUgUCiHNCupPP
6diKJbLB2FNsxzVtDW4HgvnulCbDjPwPb0UK6+EDuMEgLUssWfGKL+fQ0UecV1X7
2To2lV+t1ue1V0IYOLH0QX3xJ9qGbRtMTcbnmauxmXy9cVpRZWFWxo7HSGNLRsK2
A20HickfpbksweqMFkMpCIqZh1tgJSvHzkq1uldZ5Eu2gAPyZ1KeqH5ZbNBJkN1N
4BcoZPjkEBIzIIgfsqJ31bCFVkVhyAy4Nem7iy6wBBcYsumErPtpqImzANIck2rU
CiWDe8KQ6ID34t4Y7Du3tT4YuSXpct5wig28NfN3bdyiP5g/wULIXhxRrjbVpLmE
yQEwyZX9br4TQTY3gJ7JIBkEwE5mciTyPqCCztrIxeDRaFnHBuySdiccPKECuGc/
d993RceCL5V5E+d309KGp3dM5i3BZXlyMFoGbuQdpdt+7kbHCLnS5vr8QZnkq8qS
K4Hw1L/9qPpur6yHXCDS66IvZcf4fnjJla+xp5bmA2JK+En64RtSa5MVaKdhdPwT
tuCjfrEv+R9RhdWjHQK23N0ucCPW5wRSt9w05VhKRwaEKhpZLaXu+jmZGGB/L8o4
ePuvy9HaXEmCrx2nPvg014K7nYI0PsnqoaY1ecZj2PXA2t9ix5V/gy3WYA2z4UCC
Yi4zkYLAkFXoZU1N9xELCjbkfcrJzPtwYhqysfZjb+xZEStq0s5cFzLtfMerdVbR
5/H1WI+k13gFWwqGrHez79Ro0BwWcIHiBQOMtCGTKxjUaEGs9ZAWXRCUlrlFelb7
HQZlMuBW1W1lZnzRIGt7V/3+Ac+doAyX2dCiQRs9W2FILwGPkkXi6EtqDyMWYxV/
Of4DKmzi2EgWHbEOchObm5g234EYSUOzvO47e5Ketr22q4V+2eSRNn1/sArrHsIo
JKQKdpUHouEfBXln4B8njRDIbMoZPAsegzf8w48xcFgnxCpRcA+rBnM68HBuINLE
NsCxMkJDAsPYmgSP3v5kYQyeX5+wuwGJmTBgUUjIdEJS2SlN4JbnOOkF/9KJgJ2A
+FCetdKWoMPA1UppIvRQyvphR7h6ABMPBLPE/gfwPDboNZIIoJfw0IzOLyF7sKhC
Pz5Zi//Nnh0l6mUfYqtTl/kz3sTFJc/me40FEHGitrpfcbEbvcho8ko75RGumcma
NIl1HZRau6gG0cbUPoyVL1e291COLrbQd3r/eqkTY2RI9CArBT7CAjyWhUiR0D9X
KkU4TL7Zp3SpmhepKds7Z/aipGQvGlXxSL5yaSKF5vgtV32tXKAYCFIkHb+S4RIN
lMUsnRv/wHbjCpX82HuUjckJ7JBiFv8eE1YUhIhR7s0gTijqGmbV6S6NgBLaZt3j
dEuRd3oyymzkpss2+KJcOSryi7UTXk8LRKQQQMrRQ2ceT2bL2r3YbzPT6aYsWSE3
mCDcyxOJDtRKSjJCJwCOsuFvdEgm9uKt3KqG36vxNB8fEf8yCWhWNIrWAuloSKKk
TlJlbj7HFGX+9GV/AV3YfnV1Mbatpdga6XsTllQKwT+wmUeMd3EgRu6L4a6MAvEq
ys/DirorhyOwfwkXbjFoGXAEefGAQ3txNoSm5a3IJyTmiusc6AFsBuVx6UDmyuiw
NrcqhfduaCABI/UCXuxZ+g00uZY8BA+OJAU86WIbC9eMtU5QUug2YLWv3+bUJGNF
abHx4aVhsSm2NYdkB4v9uVDBcjVvapsH16NGCTVvoirwZXh1leGKTLzomYCdU08x
tGg0wSZ/lUVwOBJJYJlD9I7yxvHmaR3DXhrQ57EEWVFK7VVlHhBJSOm00LvQ1bo6
csmjU8rCVdPrsMgL0H3WZqINcVTJ6+hXYP7AVLt85oHfpt7safjdFH+YB55bP0vc
2ZjkA7i0WBq+uDeUZmQ/Ni8rr2Upf5K7XQ9YqgJTB9eUkXXOCVumWo4ktRU9OxRo
Llcle4fGtli7htuLRHtYeOouEoM0iPDppzFzciS+rLmfkbsAPO3GXKvHx1oyRnMd
SHJHnMhlYwrsr6gjxQv4bONHA6kWSjai/rWhsiLmaBqpLaRqWzm8b3y/E4Nfqv42
FlW29noBiXmnhME2MQn1Qi9yCKuvAzr6HR1R5b4SifUPuhsGxXtFB9XJ1PezeaMV
UADWnnYpPumx4bfcXWrhfmT5hkm/kfZnbCy9SCeDITO41AjvuaAVhZefYpQ1MM+Q
RpsU5pnHVqVFACn72dO98DfdQ9AaC7eoTn5hZrVBDaYtKxz/obIorYdN93jM1bVM
MCCtT93W9hTTXsMneeT386a3VWPOux7eNsmRlXuo2TZ3z78gyPD9E5crRsCP8+Px
/Fp6ziDQr0+5GCY313MBiCrzcejgQulW7jzlQwMcQyzydH+YBPSEE6SoJrJJGcLz
PtTDYeiplXIQzFQGWia+YHoHcilD3RRbxTIPX0BsX8OdBU2t6T1nbvwKFI0fwLk1
VHYgVi12yMcSaxJ79JiqUD4LViEYUCLvZzkAw0JiRWtNiNujHWFtkGMJNGX228ZE
+AFraaqcO5M82re7URXBGhs5ibe7b6ISiPX881mmJXKThpDOrKpyUOt574n3QbNH
lhkH6XrL5yqFJ5NmgnfA0yErs/+qzxATENSDE1ki4ewQZu3+524zJgvm9qZKexQ4
mnuF+gEvTumP0FbzbhDlR6YI63onMWplaCENn4ahpfo3qY37W5L2ZwcVW6SJ84tM
Pv6r04jLZcisaPo7snz5hEfYDBWqFjbdGybCWMyXY7622QjsxSFEvzQ9Yv5R0nvh
iK9KleGp2sEyx+a0j2furP+Okn/M1fBxDoUe/WNbWFXfVj6i2oaroRPi+gX8n6je
d1AH0+3u2xZr8Ry2gCecVlRJa9fhTZnLMR+FEaK3hjPME1dyouc0k/2rHcxWcckF
a+h6jIptRKe5ms8ISYIOUqdM05kdjZD7q2JjJRtTPO+iHPWqFjw25dnMCpQxMLit
zgzL0OCSlnz0n8/uO0CFjijl7bN4GlWMTqQ+PLioURZTYGL2i/6kEeBnYp5Laule
JTCzCLO+gD/DNw2P2y5JnSxjTDNnM1oBVCI4QsTUkcbcwXUt9E0bWZUP1f2kn1Ar
SrDbETB830vvyoeSKCmt/oZOyyIYlitsWOpWPZjF/craGS/0gFiEvqGpl691Lmak
kmBaCnbKE5o/ZRsd+e+BCXUGMq6rvZ0pW8RQVjp38y5DcOHZHi2Pr8alDdmme2qL
JofZCwG1qsMC9uJEiQ+1q71r5xvc1wW6v8WvF0URrrx2M1mRmSCaxokiInqknTBR
Z6jfvAhR7E4XrTRVyc+C5jodARut0gtx6pPm9siXwZ4sQnMoVby8QAF479AYMfRC
n5l682dn6Uu9oDpXbGmyECnthOvD/Cl6sRibYChVMQb6Hh2CDTO/Dcxt7nfnF95V
9Wbvi8UAUffUtu8891HomanGcYK0xwyuZJH9uX/++jADdvK1MdcXFhOq1GuLH1UP
mLLyA7MAIMYdd2a1PrgRtFCq4MF4Bfy0zyrk0O3cvBkIKhOzvXQudXe1qUd+NHYT
3sDjZhDh8UN98XHtsYEAfUgba/LhsIpECWB73WXmRTu6wqAQhWV2w6OnXKN9YxvC
Sk8WcfU+zxs8fUCt6tZyp2OukY3ktNRoNvHzE+8jyUdWt5udM3+pj4rlWqZAcCbL
+2Yebe+cZEmxHzDozi8MRO5yDsYvQDCNrns+uEoo6l4Mkc+yIpxtBr72Y0xDyidG
A9ifhqLZZGKtsCEpkstg5p1EpzoHsjgnVDk0n+oVauSWo4q2j2Cu6X7xznnQDfiU
UxcFTCH37rFFBmMQd5xw3DMMlOVyXQ7qNVCzfLy1NX3bGYlIeuSPqSwg89SPe6Sp
7Ed8OpJMQuhn/SCKkQVVksm7dr4us+kVWACcUetV2CfLssh9tnH9fJKwASNtGqqD
YNzfLyCmARwZcU59khJmbydMmzVcPCpdvI0lavqRqp7h6tvbyxz80JxORo2oGna0
LQ/l/65LJCJxzH5ZZH4QhA984PazIYa3FuMijNR8VgB0irhEAeqJoaUvJygJhLR3
Y2pmdHrXlNn48IIx+XGXKA7K0DYU9Ubejxb5aQHyCLGM/gR2NxFKCcLI2kB1kcGq
UnmASAllaP/t2vJH/2y2O5bFFJX1u8lOhyz3zArt36JmFMxpJbyU/Bm8eAVqiAnI
O6X3nJPT4rKHOaeLXCcZZRsYQG10oFXpIR6pkNO6ea8u/wZSLihZq1EgbUpNFR1k
G9IBDB95F7WdRFy1eJy5KOqkzf92h9UkNfd8eW2eJAssAOM14dQns0B6Du1M+gDO
pfgbRaq3Es8ZhBBjI+2EjPwrJpRVpvGVwV9J52M/Tyk5d8JmkBh7gnOSih3VXtxG
/j4+y77b8S3hzfUDysQphiWgMY3y3sQoJUvUeQMRz/SOAHRGQid3rzh+8/+An6zl
q/vfU2/JmiqJ8cExq51LaxaewQU+3g7ZO3SeCuoecrv/6hRhFXuh4um7xWZhZGcg
dBIFYPwwT/EDcKXgnybi79N2rKAQ7IH6x8ymbCFBXpEqAQ1kPh0pgbKf1q4O5zTb
IZmYDinqA8gL2U3on1oiBARwfFsM56015BJwNb3X8yL0yECdGMJbjr8gxkvmHEu0
Wu6kgxiPkUsqvC/m1ASOW+djMJo2MqGeJbohvnTcGHRTYdM3gLKnMoVii4++I81W
PhgLUH6Nj+Ktp3oxYZdcOKgUy1gQ4Rgf5Vx4p8AlbVEF1Zx89iOet0fwWzrMvHsm
UJRnRG9nWstJ2nyjLjFF4lJXXnkRzjTTFEu4c1kRtAcX5hmnLiLvm6kkmlP2ZwGs
DvrDEHbVlidi0xAYekg0/FCL5u11Q+F6W+7HBhWejHGzS8ut6VG7p0eLkOTSSgGV
EwuTKlUS9Cmx3o6aElIErInsVkewaJgtIfyoWcOf6lLKzvoOf38k36qy/yLMxU37
W3x26A1NTj0ApK4Q9fXJDov588zBoomvWFE2fGHPW3B/Uau8DDvVIyN02fBPRlE/
OalR3NgldC0k6JDjLRQFse9GQO2jnbkB8Cdx8hvVPCdoagAhuSyu/jfP03Rl8BI+
fg1+G0tFh+enk6MOF7kYwlrLeC+SV6DF99UPE4C8NHvaRtOGsGk6NvvSzt4aN0Pd
JBNhxi7AyTop3hUTvVlTqF1umqOKO3Kids27KtFnPgse0SZaxKzmOS/I1eLPAqlm
UjC/YY8PvhKErckFP7ZUyYlc9H5vDlAwbp5Zm8QMBdNnfXQjEIo3OCzVndqmvyyH
eqL8VabLFaOU4JRVoe+5uzYWb2Kqyf5A2iqRDvShDNJwf1MPTzKOsYQmBgUBTaAw
NZYvLYphrWbmDfBqjy2Xn0wyd0bhNjPbNxkyWHzbEncogZOShHmTsnlcR1Fozq7X
3LTJJRx3NZ9pbqPEMglzyZ9rZggqnpkwP5bT8ptXYPTkxwRcupTjJvZS9MEzwO8a
YWxvElPBATV6EBFut39BU4QL0bTwDAX1GVn/SDjMCtZmrWf+itrRh7VQ06ufAsXB
h3piTu6ntgeKYpzW7NKBUlqndwIYiW+Uff8TstCVuoz92Rkzd7qBErCX0Wfwabwf
d/R4zpJ6bpZEHDqllZyqokRuKT4+X+M4acVCjbiKLxfUa7lQsrTlWV7dbmLvWvpU
hqPrQ9cCJBBgS+OHZSNaZ/OKqrFt3aB3RrA0sGbLZ80GcQwakmbSY5cFw/x301DY
eo5tUsIkhC5HvkNoZjglCnFLBlT7k2uPr9qvu46grIt9cvxA+11Ckkzc9a3DbGcU
xbm6fsBp7VTZgvT94oee6u+wscOSdGIfxU12l3j2+JF0auFr7IPtd2mk255vqNz9
wY1hiWtlPHrwl/cDOjKvgX8403Ag58NWmkrl0NLWBOkPGXH7lSpBV6CyQXPJXK81
PuYQAjrLFzlOz1unQ20/XXhQkPf01Kqnqpas4GDeEd1Ikprt4fpw3bvOSeO0+CFb
ie+kpRQXlPG9nC57NffbyWm0rE9ptOaGnSfrTVT1XK6WG7SZWdqDsq41lASZBHGG
SHnd8zt8I5V4ScKa+Q24bC2iFUFKo7u378T1/C0y34r1tSOox+POjfadAd15ayb6
BTrkI2RpnfuIqMwynK8SsP/AAHTtCw5MJrZbTteWcTE84vYK32uYGzFggk4HZ7TY
IkjFj+Vg6xiC2ahLGEghUM3Yg6a/JMX21iaaNn86yOUD5/wA+HM7qZtcu+yKzhGW
VBkWzzNOS3uCm1M5/UarJmLl/llajgc6K1wG+7T7UvednVIDKbECu5ZLMyHtJv8Q
tsds+JmFwx8maUIRBdm1cIzXq0ho/QYm3e7LnNcx+Y4mkodD9rwgveqn677WumAZ
dLMeWO3GCnrdew3Mj5oBnz8i0VEFUsLdDHMybWJrJIWaB+rMZJPm3z7sg2fGdlgQ
9GvCdwUIBDKZXX+kJrz8MKz3SL+YHtPC8RTh5JY7SfA4yYHbk/3BlX1tBYViaiKQ
+RFyw5o+ehXNG+QoX0Ig1NdabDbmtkZTulIGZLgmp0pkmHA7jatlnDk2UwmXGv3v
+ey9KmjGL6G8CC+CjFkt2rjrzbcVcr0RBJKqq0xjGqlaZUDyVvkf8V2gpGSBHyMU
HcZv/Orpcos9RkVpQnoXygeBryGboPfL2NYXhLCk8UK7fJFMJZLGRCSzFD7WyVa8
yH71/6Gbqm0AfdIwzrT6e9lKGMDUX8yeUYfZyKJQQqyLdcoE6S7Z6OR4x1JHKZkC
UCiiqvhh5z30vP7t5U+2QhtO7UGAmz8JFLyvbrmo4Nt/947xjdHFGojfnBAezmzp
9yfuOZLlS0su0lI2c6sDwpRm1i91PAp5RZhhcny5hQOxnriwICSOsJNY14SpgaRs
Ux6V7QcLmMLQHPmN6G9lJ6kh8Hc4SLqt58pzrl38iwv9xiovxDubcK6q3rLrHnGP
G4rYYGcImfuEnbWnMIo8aOqdrYP7UfweDixMXGQN/SdzPGjhaaDOuVA1DpP1Mg4V
SMLlWifG6vLXzoZydpiTft6bjaAZlI0p0BLXtS9rRevTk/Tf1b/QaSexWX7yldlU
5OxpBvR1njB/wIkx72kSX9EqWhNurvIQXW4vbPyUkgY+HhaSoluK7p7lmiW6ZStX
ZnMZdiHF4+WKzIKgj3bxY3GOp23tRSeN5g8j6s9YSqVqiAq3M2Ij9aD1iWDBfo/b
raQ8KApZZ1CMj+qsPXwQfctJkFYuzdFWJk8+JygxNgnngD0/pTEHZ6z1rSKmLjo5
BdwUIKwHRjm92U3Mvimxxsp8mcG5SMKOA0WauAfei7eu6L6wcm13bXkoKABQ0+Cl
xeXMb8a2ZCp0eMcXEaZXdmg5l5CNJWhuTpIE48c0k24PevKwQCOhc2wLBASF6IZk
8IFhv8hWXDB40AzwICWrlH+yUTZD5ojZ0l1011PWUR7Z3k85hHJufZeLBmicd+xd
FKOYA/NmPGZdY213HEnlyR85ShwjImryh+lzeKj/eTkmaPQQcfTrs3oAjYNqoY3u
c++CJ5q+LUSxoBLNvAqV3obe6VLNBT6vzpFVwQOG+1cGiLB6JyuwMDSSdV8kPV0p
CCdAzS/zDXPddh9epj6X5PQfdzMeRKmGF3QFve7kjmjBwksKs3HGGoOY1jBRRz27
EPMW/PA3yjDwuLlW4ruAZUSQKuUXG6lVPu6NHPIAnnhSWAEQOwJ4o3xE6ENJmQ5I
+clbyoYM24yK7QCte544KzZqWxP0VNRMEZyeBmdeypJNv9Jhg5M57GA6v0oQaaeZ
xonaqL8rinQa5PWFFBj+ZeDokaneFwtaM/fjcGxUWi7QeZ0YhRdPVhiPVzfMI0ub
fpSz8GihI8pOwGc5CnpP4SzuSUpHVFf/Pj5TMqPaQniIdTXMYvmV0rq75UbFIEjE
ykGYlN+HlUQOYE0rEc4tquvwNs110eMURacQNGaJqLzArwFFGPUIBydU6CXSnsNy
toy+QIZEVcmgVfoWukFE9Zcs0jNtiEu+5Y5KKSxZRV4uEAqsNsu7Zx1VcgTQb66H
C7VGILwMWdi+jFcuKoMGKUMX40DTdpZ44J2PO1o18C2QCs9QKAfdw3ubG5jOWlay
UBJWqpx36wwAOcDFbSHPjgV/uGV8eKR4KQTp5l4sMpotpdlfG6xmffPdPRvJp8MR
W6VSB0b3GvNGiuxz4DeWJ16GyILoMmsVSpCTnErBiQPbWgJKquA7HAnIsbJjP0fz
CSDg9cw7XxUhbAJXSM2LV4UsWXOJFKUb1E2RfoCGp8S4EK4R8VV7ZMyiQ449cfIv
W/k3JupiIWF2+htwdmvAjuxId+9bp7fTxXLZ43phQP4AeAmrWvr/Fxee0jW+4FQa
DNQbP7qqsiwH3qB52ta9iZUGEmOFIGBpfNu0MVkS/kiUmdLRGQ85kT3wDpBGocuP
HAKPRAn8d3mX2XIcZwIhJyIMKYAJs8JWF/Fm3S6n7RVCpFi3BEKHiz0hJNGaLgx1
afR1zSASO9qDGDPzUFId0Rwe5bell7Q9SzKYMHP2m1cCvHoyYO6l4ETwacHqxpxY
E2MY11slQ+KFZAzDtkKLa3J4YlgjY+umg+QkvpFBeKCBZFVQJd5InpdJL42tnFT0
Ci8/mOSe0f6oque5oryIRH/OBzghLtCvKgA2qfBEXaZAg225OiDrIv62s9m0fq9b
o3YaxiX5y1JH8K/GopSLI8ZAIFkbsrks0NMycOnFyupnc5tRue/aJpXGq6Zjv024
9CQodNSVEPPzju+oqeIJmZuKzLnOoK9f+MG419fGVTNbADqnnRcdr18nglSwgBhr
AphxScXa+oJZzXKz3blEI3SG3eRZlNSN3CHUrSY2AlU/Jbskiv/KJK7cm/b0/Zwg
ZlFvZ8AVl1DhEWOdLOr07prEEE8C5ciMcgx/82CEx+qjhUrXS6mD/bQ9qcChsXRb
RYO18bE2EmmMFZRDW7qNbSHLZ98WDNRsi/yQA+BW8dB9qHeWAbq6H+2GQlspQ7dn
gZ5JyqH4xEmMt/CdBDKVjNqhi+rkewjwCnvMfk/8/rFhcqu4yT6d4mCh7oPNjWPp
738t6brN7tBTgHUTVlHyqlFz+APeViIF/kC8jeAMJU7le7sWgyW5rWeN4mzuHIuK
lyQNlObZWrTN1YbM7lAQh95Ka19M5iN6q1j9tpqL7iIHk+GXyNtGgTjt1rlNKIX6
uHvPV3zRhyuVGcYo0dwiXCr/0PvYzOm3UNj5s1eQsQmG0T0C3rb1cdQc6ItbSoQT
z9Qi1JqOrM71hG3dWAmBONGJpzSuF/EtwgEEyuBLaKr0M6MCrSprUos4HSQ/C1Sq
0tSm9/F95lYwF3Qw5Zw3uCu47dTqaPx0Tadp2vY8NT4eRnefEzR1NhSOZDtc5VLt
31Qhr8mHB4RfD0dwXTNtklcHgogrBtOAsnJLL5UJFrRDywp5mvFOhOJLi7KrrKiB
wDBu/QJjVddxCnFi9HSr76RVJojkpqxOPlXO3unQee42pao9F7A4omTn3IRCOV/A
7tnIM2/F16CpLojxraQAImZTBS45CaBdio0pL35Y/CG2m48fsfeh7re1QVoqgMWG
wM0H6YeGFeq+vOk5faMQKqHIX+qQDKQA1g1hCtD7Db395SCQgnoSmA2ZL9F5s4Qg
JptcdPlb1GwaKgabBl9bn+HTsadUlw5YLvseFWpnmymXlYBdAVhBTncVDdsxS0OL
P++KSVP9wNReRv3srRql/t/Kh/s/xYynBUxGt5HG2qE+4pan0UOihPSUi+Um/IEM
LlXiRSWtrFKwihHyHJqJaXK2IP/BMMmoPgL6nqWW9HzIfFA8+CJanH5/KCjrhbP7
1g7X18+gTumxrlbd+0RadrxVMdYd4KWj5LDQS0qczdXWEgpCBe0R1GjavtewILw3
SIWqIRZUsoE8PP9ITrF2g3S4cgxyEazkGeazOxgmYCWI+PCMcU1kK3Ph0+2qvm5r
qpjitE/dbyWbzkfepqcHbXxQ5nENqs+T5kG5cMaGSsSfPLOSEHniLNWJMbGbESyL
+jyDAZ43IHthSV9e/6/M/OCgkR1rJzQZct5TI+AKaHGTuh9YHi15aCIszxWaL4P4
4VgfsQIGrht/kpx79DAodiJdK230inYx3eHUDg78EoQ2MMwXOkWp+1LEi6qAf/Ps
tSqEYg+Ui4YraiaymN4yzdzNYdZumtYLuLE3L/VMo+VYSLyeWY73tsPGkX/fdGQ/
271Vge4Ze0tz/2r1+PWcAGdeKl7eQb82cwtCPJbGmG8drYqAPTJncyr24uU4Ja2R
z24OJxO3ZPxlwUn3FwEWULTzl6wkhP8ebiyFOvlh+cQB1FmQAKyXN2gs+36v3d5T
4Z0IfDuU96qZfbwVLUmfHRJV7xW4CfPD3kn/Kg/D5GTytV76YlkHBlL/ypZoP59L
k1aClVtes7CusGA5BEYq3BGqVNyjTH0jL1Usl2aY7DygjWmcR6QeoiOFB/2ZQ1pE
cFSmM7qgbUvm+ppmHtY60HHISv4h/esgvUAPXmYg63fvkqqi9XyI9dgh3cGC3dYj
Bc4xQNIJoeB3wKc7R1UVhGfDUpNZvFPhXRxjiKGkiKfHlf5lXNznQwcYRu7MhGDG
5KcFc6oSxp4nEmJrwkFk6gT+UkSse3jVXJ5Uhr2g3nfCcsbtyplKuhcR6MJYlFeB
Lun9b4HDf5GzwIRNcygz+n1Tyvhfx09RHgmSVwSHVeSiPBOrN9KqYIjG5qURfQzm
+RAzX2HYMpqWMwQZgnfAtqDIex9Q3lyfIDpnG4Drm3xdj2Ur9cNBYghKQGjXpdpA
w6u+1RjrPWUy/PMozA0B6YZ8xwSXa6/Xapb8cp4zZFRb8orZkYr5sUyX72/NAaXs
xWoy8IxB43uZfi9FiTwtldv1+bP5PS7is+02sR7fRdoT185XFLU4yMJS2FjXX4P/
vXB7ypevp85Rd5Q+bNVCdJuqC330i5eQOMjRNGyQ8t4kVfZ7XB+nHOaP+FhY+F1H
AE/5FYTUMPn/nMgPQf9UMO0c2J8/bGb3d9hdXBvC3EYe4A1mnZ1qqrwgOaBQD8/f
xhIKKLC2haEjlrvD+7WLHiGegoKpDG0NIkBiAfbdJeEZ5Kjkw5UZvy3TH05biuJP
1YZCxRBiXMfFVabHpx5+tokvAYIo0+YTv47K5uST+Xn10i6KmiidS2guVbmGNObC
4bXJ33MAGA16YiLhroIXKRe8TF8+Mgg1DzcSHxV8yVz2F84Api1oPecNxu96aJeg
DcyXJHXq1XcHq/KKxdjteaAOo1zAYWQrTBIhiU7okeDLn98/1OMNF7nMhr1XmqhD
D9QgGs3IVLIxNPn62IVL4LDfTzfnIVPGpFWYZ/meBIxrrccGe6cDRhSYFnpkcSXe
dh4rTPi+UYgb7MV0qpBf0CoE/eLnueb2CWnUaAXbMKlIc58u6YmxXe64MQVgssop
2N1FaChipPO3XRIy7gPJ76FijbTX8Y5N4T3Bbk9mlvAHa++mT8QNS26l6vwjqU4j
kEFhqu8bAomtAcKa0OfK3Ws9E7KhZvZjZ7SY+4qeJHadNGsF8CuyG5kNQ/HFRkym
64+F1gukCwX7gZ1W0561DiGEX2RXwRzBIzwoHp0h5/47JISE0VONA+Q956ou0n+J
AXQEHpzJXGtF/bAC614MIfmljhCioDkh4dvfoMUNjZ5oFep9oRDdsYDl1EQhiKLv
+IsdJLhvqF1djVzNtmNiJNmz4Fsna7jtmRsaM086p6ZPP9SZK/FF+F1ysMbRTZ30
BlD3TPcqyAE/XGEOoTMykEohAwBU5bs8qwzTXGugAlfuBVJ/hL/wgQnLGcL+eg2x
GDiJ5XfunGPKJFi1z9AUbtv/FyUahizQvZW0vOo3qAId9eqr2PEq5tRR/8ZKaMdC
aoE6084bRTl9nsbn1uMNwHJU9ZQESWA3+so4pRv5UVlRRTOpHs5XfHhwJ+JCMBkj
yTRd0krfg2eIjAlmbZBtriB4sS1rjZ/PYsd+bKvYNKKs0qXS/IDo2MoSaahvVrnv
JIXqn5b1Sx0ipvEYNR81aghcIFgFwfNznrfGyTQTpqnU6GEJkWRV3We8A8aryryG
kzSNg9ssMSDI0J5nQA6+BGIb1x5fuGRlnwohORYfkmmpYjP3okSACqPU/Exyg6/e
dZ4mCv1oInNWDUWuxdZi7uQmkJnp9Hdbku/KBBSKrnxa5x47l4SvR0TUBi7/Hnnx
dCVwUieIrLDzzqM495InErqRb/oE8cma67i6ETSs9HsBQTFUh5P6jk3g+zcLRFUG
njUf7SmoGvfQIhc6ZTKU7y6kDyyDUxfrpa1hW6G/3FLc58Zdt4quF74E+w/LYMn7
NpdYVpAnwcbsvp3MtZJ3yw9vOUBiYemdsuZRFIEJyMI2m7WQ2SdaKSMc11KypuSD
v4Eh/enNjs6pNVG8DnUtdqK1tKBsbn/omYeCWwUuF/pMgNOLzOCjydRXZUl+LNU9
AKm+tSPpuXtF/ZvTqN19Ns80u5giv+b+J5B2cZuiMSK3z8zdtjz028y7Jf9jPQ6p
+B+CFD5eVUyVOHdTaXDWa/FPz448Fygmv/twLyZ4hp8VyVA6oSpDdY27pcIo58fN
DY+/WYMg50LxNg8PUlFWpSpbEysIqMIj66adXSaDhWzL6T1txYPWqPJ+DzeWLzQG
YqN8C7T2l1Sb4jAXga690rD/Tc3GPZdxZt2djU3awEoswJn0U810AEWL2Whc053j
Luff1Wq/hnywcNsORtUXLKXTirBjYaNKV+wB6xQIrkekg3G+gERtpMRKP7ox2iYE
lszdJmbJdYsMw5AfbpVJcXYIYvMa8UpeUDPyyfel7szGNwfC0nBXxHGCplM9giws
z6qvnvp3Taj9CXORB9BlVtwDyjkCKv3YkoZS5k2rPJ7DoCVlHcXBLXHGQPQ3aEUq
ht9ZQrzsKKgLcdT+QrQRAWWGc0mWxFliKii9nClvv9h/GGfXox+qK4jvq2vThij6
Fmn9tO+Qeh7/aXu41mkiav3LlO79neR7jZadaiNSRlOETRb71z/V9R9PWmQTNf85
O7dy/l7aBPCu1X7rwqgvWqI2SXIL/z8bhztSDeUdi7kwvI4oMp+E2pnus3QYJwr3
eG9N3PZW5bL2gClyedLrwFUM6O6kdkxpFNXMw1+q4sSm9MlyXIh+pom91EDZlcAR
Sv0rX8nkrtXmqfLSaXbNrwM8og3FtBH25oJfyPFbXCCvnrM2FAu/SQE+5jh7CMP5
Q4NjWgUdWZZOyC1Izf5QhWSNUm8NKKhEpaegdN5S98eIuv0sYtn940dXMHkAkijF
gOf96aEl1pGNO5c0tMGNRq2bSWOA7/OICXcpBACYrYhSBuFt0Y45nbbhn+y8A8av
nxwN5snSMNEoG/22c+wLUwMpuIew/b5mL/1vcidFvENuNWHB52dgxIfo4AOFiDaQ
HzW4PYpKjrwsj97UXr1htyJxI0yMcEYhB35EBbUL7vru5pCr08w2+PWZ214JMl4o
H0RBWXfFJXy2mgautdhShbYMtx7r/gUsUwVW/JY0PDWmQJovMLlI6QMPk9HPYbvJ
WykA6iCz1UOWCHeJHurME+gYoJmkYCwj8Sr02ws82n6+y/VkmtPfiydbnzQY3thL
3l4a0ojeg1IFdkwMpzJV5z98aUJdsUMjy9LnJk+HIzyl4MkhYdW8meowM1wE7JJ1
BVmIXr8FBBBQzptC15RLlOORPQm1iqC3cA5w87QuCikhExM/9kAz/GBcnF+NEloS
SXYbJsq54/53N4tR+/dLkdAXGaaqHVjf/r6xjUm/0xlCoKDdpfsJJUCToUl2AyG+
j45OaCHbzL0OAVHnzAh0AsOFpwFnxA0mbdh9YiQqw+WHnKiGKcLKkeEDnvFrfqzs
hl8XQx87sRqaRRnE2PTjZRXyuD2eruNxdUiA/WIFHWx80nRt09nWsMEEEKav5FuW
vK8U4XsAcHC0IMXEgApMNuH7d5/rsPub8XNfz67hRlHaC/UGwNOPlAmVFSqDHir3
xRMzrNdKv2Yy+CzpiYBJ3QVVIbJzkmaE5rCqeFDyz1OQ9cJ05K979Y+eUAzWAmpY
ZxJyJx01p3ib/Ch/elDaz7cezQXnImo4dX6LqrZB4o+goXF1E98UKdFfTV1QwFl5
c57lUY5EZS971aCOX2lrIaG1OQfTLGX54Kx2atU1bE/0qs8he+IefIyyYNP3bKmq
FokOUrtI7feNqzdBqpt5/4McoPOLExr2LAN8QKza1+GIzYHL1bhJIhOsJxe3803P
7vfA/jrrQ+RCseDgsvpq/nUAozVKQ4RGZwGMVZ9gviP6zeNcpCwxKw8v1Z40EyVY
NdDOHcGi0qZNMS4q4D/QA0O9YiFM4J+RDUBzeOVuKVQGQ6OELbdZZNP8hvzBQYMo
RVsKq1dSPE5eAWfRBfdTeCThlxDq6JLwo1P9dq+iAMeg4fXyeYNDw8aMbLPb45i7
q2LE5nKgct0Qd0SQfTG5wnqbMWI9D92St50cZvosQCtAH1xK8v8WFV15jwT9WpQ1
tB6QmaQYeiDKWcuLWYGQ68mwk02JSnh7Q3B5gm8+RAHfq5Yp2IykCVlZ9xo35QtP
ypVAbdz24iycOhcbvPDW1dV9Bv2SeENu7OovfZY1UE0/Vk97xF2/fl6U4EDsK9C6
ew7IgMSpi2c9X78rmSp6EfQrCiCW7v22HaOsN15gbqnknCBaf3LhGlvzS57n1KdL
IJmmxhqtZWi85B0l1cS5HGbAEhL0Npc6rRDlck4ojAxa9GYI0+2E2tFOWv1Zj3XO
fwwhM3av3VYUdaQlNQASDY7jRE1TACUlG3ms+gZ93are2F0AAlRomVfMS1tJ07l0
zJxOOxAtN1JUxrNhohOXqhN+nPx4QOTosvvtE2oGXrxjlSKGvMF4j7xvVp+YISfQ
2mBz13UUWm3yQ4n7Go+wd5I1aZNgxNp1qOfb81isGxv7f/yZb2UKQQAfXgQfFN9y
7+FddkNRWxgK2R9VRXdGr/7xenC7WSmGxqdjPz3eZwwGh51UVF5TDtq/N0fODR62
aDK/b4j+r8m4ZQ+X4h+JtrR8v8y4CGko0R8F8ne4OzPgRgak3Tqn0l2hgv+xEZOS
vfCb6K6T1fLgIvxgsdZt1LrhqJFoB5yesp/M+HWhdTgOZ1SKApxP+Dm8nClF6eWR
zVRLMZ0JuC0fzY4HIzajSpcCMp+IC8wiaQWZhcflOyf8tC78Gm5w6nGflRuLT76W
NkvI84K7NjKix19KAhzywqG8h+1ntK1mpuURjbnZxPwDGXtZJWRE16ZCOUXbLK8M
SKfWKuF2iwEvdL9cTGqkS6eU7i4lNfQt9TIgw21klvNxy3lUZUSDCwWsLDxTsSQM
9tJZv5x6FSzwLV3/j3KcCkAgI/Zi+DGA2JqlGQMIPcCbJ+5jjKSrwjT5ieoi/z/3
hsouxmUVWhYd43sLjVUBLk6uzJmw82MeN4+KiNMVFIlkSxBwPSwV+iLW6jWOXnP0
hcLlxa44s5Usn9L+vqLa5WEXEjcgo2In8SSsV6W0wB/1F/gZ2Uet/S/+ykcVdPhO
/5gIN7Sl2IsETD0wceU7+w/FduAtyptxWYKkTm4r6JMrfcsWsCy/3/z/5yD+aBN3
UAVMYXzbHvEv9q4347ohcZ0/cRAb8/vORp7J33cARBXfN/oPPyrmXk9f/SLibgPv
VOMstf9yzmejxeOj1uEDrdF6Gd0dzhNCRIm1CiIn1krbGrTEcMmUfM5TfGH4vqPl
G14a3j+PBFpwUV/Vj2klMYiIDXqWQaGmcdL3UmNuyOQp1Opu6PQFGgCWc84Hu/0T
oCX7eO2a/SSlappgyQk1at1fF2fXEKzQ0k/9GiM2IYt3+fL1D6ue+6qXVzympz4X
FhxmvEtJH+JgIWU7HSpQUSqD4oAP1AIPvoh/4eEa3KFREUlUCl1UiIo9MN1sp7Jk
5bXnRE80GqH5IsC4i4By4tEW/BpY+TgE2evbKmpwYxzG+FTUjHq5YY2ZXkxqd/VN
X82IM3e1+VyWdEXOB9PJmVN9ecKCHJIKIAcNv1Z3dxylSEWwgf0ledABLN+034VA
cE8cAmxptwydzl7pQdtoo2kSp9L4rykx5Bi5S0W0g8EPLYMyrv55rJtc0UOukGhL
FJtrpexpy85pLHacfaksa39I4buYT+PQo0MgXSn2fHLtPrwDAk7Mu9RfOdWgPIgq
GYzv/XyNeNcdbMZ7rCmnweC8uBStkObC4Iq5i69YW0wXEK2CyDS0diTOrbqGlxwm
UrUv4Gv2/bAgnlcURzawJ5mraf/OO6LCzFnACH7mQUAl/uaRPPuazd8GBSlWfWFr
DrpvPxvecyGLB27V63L+SWvrK+NBLDIvZPyGIinA4rOSNrzRLq4EwRo1+yQyEmQG
tsePPE2AaTox8imYhCapGXy6zXLB0/3RaJmt6lijuiCEljtD7cY6KC5mnui8F8jD
YGJg43DECmPJZZ9chDU1ZACyEwM/RW0a4X3KD3bIha9BlmDB2QoYjRx1PxhHAcvp
MIAUKXyDC5GDnbilNJqNgdjOJKpll1qChA6I9EAdTF93dfsOYDhgUOd5nhHmz44h
YGxt2LEDuSL/QpsgRG9gWZ//m+NJlUDxI3pKVOS0WeDMOUQU0eZpsZMJHjjYsxHL
+4sn6cxszvg2GtBKpGiULjBj5QuImYJzE8WLSuxIx6cYgbFQF8EKoWGALlgN4zKQ
tl1strGic5lfGhskb+9Ib2o4WcWz+6Hq+6QzmpVkpaxQ9+sJOk4boJtQ7Ft9u0hd
dTimNa2ileG8yZMjaQdkoStRG6wnSZRte3B+DGHRxqSM5T9HrLbLqmAbU+opz/AB
c/nnlGzXQpFViHyM8ThksiIb2HZJpyfKZEVhaxI9268/56gDz3l6SmQ3ZZPLll7t
6QRNVd4a5NzGWokNlfrbxsu9glYoa+bcOy7yu1ueexsr/C4yloSH/EblwdzYxQBx
7oo7UxVHv0KhWCFDWBJoA9//qVZBYrYYsRShl0x2tv3zhZSNugSRdv4fpQLlrppg
t3vKzQROlzkCO0/vBFtUwFEGLatMnc4NwAXqpf59yy3LpyqrmPKr+WY4DtfFTaDl
J8emqFb+ErjGH2nmdemnoI3f9SmrxsaCEmWVmTYlfnpylQDyM5Xq3RH9MEOVNumG
uh4YbwDCwAKAQnPwNSNd4GCdT9UonDNu+mIEeZCY24oTpGnYunZ1mijoGizEX/Jt
tsv1DAFckb0sO7rR9v3k7PINxmh0Imy0//L/x3YfUvdcXjK1gF9+BxQCuKg7m+Hb
sgeVRCRP/ZqcqCXqAU+xxfJGdLkcqdf/c5uzTNyzschMAxP+VC3Prfz8kxZcOoJ9
5sSlQG4mj/Gr+CRcWLXJe+AQM+Ta0VBOZiQRgWjwXo/s7vm7bOMUz9yQStoe3jtl
hBrfBYURGTZ31cIW35CGupvrknV2jDqqp3tkCEKWjXaI9yKENdob9aFYuGG0rvia
IH3byJ6usWZXHoUdKlfqFgG4Fg2Bm3bj0OqRmBHbmc3M0FJmmQTXprrh4MscOL01
KLChkjt20adA49V//KWrOeUunuEmBpmM7OApPNG23oDRzwxfQRx2GCWk5yxS0Qr/
dJekacmUydJY9o9HUpN7M2NmNOHizhmZ2tBT1VahUhEcVMuLc+KEfDSrdPWClcT6
+DNJGWugS9ng0tpFudON31hD7+eSFzJ5bKuGTjivko5fcwZ/fImNQ3v/mrnLED0h
VXdTvkTY2cTpY0beKaD8AxZhIBOHRDZKmNWEQT2tOvadr7C7qtKkfernvNSO251h
ZQmXg1ohzquSqpdfO5XtFRyke2eJ0ZPoycfq4AHyohJVQ/AfXMIJva8G+dhxTF8g
azJbassxZ/KsFcfnpilnZmhuwWqlZeBJSmdy/VU0N0HD7rCRUyw6NGmhaLzZYCdw
N5kGYGHVPC/AUIHd4uCt/HAgxxWQpU+MIPzndsP/Dnek2ao0YpDiGVBhsib7ewgl
jGh1fh5Hxn0rd5VEBsvCdxs/kmctESPySsiuK5ZWMd4FaIFUxQF1vufbO4xSt1OU
MT5DLAlJsuxLnzT9yUAVM76znIE2YUWfEPsE1IBCxi77mH+kZ07hB5VNV4yWPqIx
CyVqVErI9/u1oXqy3PwmomTTJYUQzo3nTYM172iqd8d601x0C6/n3yLJrW2EjmrH
MHAOBQ5eJ7qHEPhlmSIP5xYQg0I8rjuFiDGnCmrIpGK+P2CDDXwoxHiFuAWf8+bp
5nbqc8MWWjfx6PHihfGNZJGmvnqPzSEGc3bKVgYEHswLyeC2/bbD18i8jP3YeMo9
52k/cKHUsaH946Dn6Kaibj5yyx4fSw/fje/AtZmdPq/1D+G/oNtamiMHcra3sXZ9
xTRJZFU8RuRXWm5MWSswZqCGDJSnQSHDqmuuVuRXANeNMzkvOOOgzFBJjRGx0UJi
xFLSXopyYtPF21ZT53tXPNJyN9Ehf9cuMqVs7mSqqv6Dlxls0bwtkZ75veBF9izu
q5j+x2SEFACYQDr7ic6cUASrEMn6AsCvcvtvxJ37+qlQPXREhD0hF37gjulhhR2e
HzrcTr4giPk8TSh+otYivDNP8N7JWFvabnhWfa17/qsBspUdm8u/gG1ODWjJXyAg
ZXnYPYkf9DSw/jC8bZeTRA90SfUDAwLQVgcPBmMEXPJ+Q63SwKCk8DCyH2t+0uNM
/uPSl86/SaggRiGQDBjoS+kKc14ZRiQYV0wFu4Ds66YfLvXvejq96WbdicGhXyb7
XdiYMMlTTwQm6+AK7Q53ceOZCSoeEwiw/zx27YSAUokTtEku2JSvB5iH3A+f4RUy
DIx3dhOjqz6yLaExob5yK+vkEwFi7Dt1zLjVH/6ks7PVITy6QnRLYI0ShzPlIPnQ
asHNXk7Ddr2hidNuSB+XzlBwq95dCLamIF12IBv9+vueZO4bEQ7IM9FG8BMfe9Ej
mY93MsL8zZGep32vr9AcpuvF0g+RjHM3k+586JVICEJDj7iW2fW84cmXgX9i9SVh
Z8pCC3u3+3l2AYtNzv39jvqzAw2xeFr91fOaaMeKoKhxUcgEtBcgWECDT6SSn097
hg8tKvFtjMpbjQZqQ0jvImiPLBfhuSRt8U/C6BqiLr8nw+WG2iZ9yicpEnCvYNty
ZhCK+luyh//tis70O21HFFHP5wVDXov6Idsbw6Y+AeG3JviSZc/+zCM5F3lKCULu
yLnu+IKgGoknwauaOutAnNTVGddR2UCfiExEh8tMsJdonA8yqgAQYr3VnzyHvi5O
LZ9zuBq7zyVruzKlV2Yn8wYLWQldAAvvayHIiUK0D4kfy22tNhBpqkrbmcyvVbRr
yXmef9+NxAzYvio39SnK91AfKZ7VKQLQOx2ZqRqi8E64QLDoHISIDPl0jNV+7ilp
3M1ozzGBtS6fgUEN4TTkhV61xe/NVV2iME1jAV68xhsQiH48GqxLxENfyxyRi8Js
NftL1zP8j8t/QeNsFEd/T1IzIBS3OFnIAqjUk0vl+Z7yge0YG6Y2Foh63BBtFK5H
6yrfNLg+SLsxMDwXcCNJWB5/oKdwvYxmHMW3B2tBVj6enzyIdQ1INe2AjAlRXY/u
YeABT3lMPsUJY7Wx/zcEgNxmUic/Ue9mmhQuHWLcc32+IvklVuDtZPiBK8nb28N9
8shZPFQSovRFDv6J3oQpVlZIY38/ozQZQUSDHDzskO+nkHhIGsHommRVI5EmSzuh
2vHOyy5mRuQ3BvatKVkC1ufmlQxm3Hs1IbQwQGZhO+Itp2bMJU2FQIVdVzZXkNnr
Xd4L5U2WRp14Tih/qMooKnp+uVEs+2qLmip5tJNJwNwBniavZsNankl/fmsWfFyn
rIu+iGEu5k+9y4wO0cT6QZ14IUkiTxjQLTDBEhnEDFe7N7C1UEErVD4+WUpHqIXW
8AYSVnU2nn5r5uACddgVzeeoypwIdQ91rMl/J/GTAfmT8g+wzym0+kiJTjvtp3tO
utMWmbXYfF8gE2qoraw3ACA04JqZ4ycd6HlcB1eSqKfhRRVDcJTQMyY1BTo53yEg
pM3E3r+0yxJO53OafCDre2F3em4hEYVMaKjRRbN9fjxHRwAQGKPNb7Y4OLP3Z07L
U388bIOy6xTLcm5QlocYCYPb2ZiqniZGMHpY3/pkulvvcrBXd7kSUcqCfaxoX7cP
0JtrKuLowuacApVn0PjW8K9mAUj1yKtxzbyhDJkKUOrMcaqCAp6KQSj1UjmTOGZu
ORcZ2tuW1phkTt3L+RtpChNMXhwFGnXUufyHYOs5SJMrE4j+ci2f8YJhZDQ63cFN
/yU4FlobZspjnqZ5XoOKkJPwiVQukuv4F4ENiug8PJDUkhO0BeMqwHKujmaEFJYL
2npIKcdFcUUolqyFhBJBcYBlxfs5fR/OSaj2wS35dQ8JkIM7GRzVl/UBQYuYbH3L
t8nDHO3xMFz4CYpKq8c7YvfkUccMXwqymh+aq84867rxW8yyKW10bK8k3eeU0jnx
zMNt9SYq32weEv+HgIF16D9GHyxfE62AVSeFG87VU1GIlabEXjpWq4hAdmpEJCs9
nAhmytv3J/wSZ+9sw9ml8ym90T+2Q9lerfrz2NnEUmHJHHSN2jlrlSaUw7rm9E75
zguN421Rooa+7GydNOQe0od7GNqkDQINIZXYlShsuquPvVvHS2Ta4U62YJOeBU4C
L0YIwAnwdvKcwY1GTWJ9g67JjzfwRaFUELZbMTi6ZXZX3/6IqUHUH0PqvzIQYXz7
kysnkQtuG9U1LubQKgzKcYzNEgWtVjw3JOB/BcZst29odERWp18l0xLmA0kFjEYo
hC04s2yrjJwhIPEPQ8KzlbjGw+vZlmSPTBtqQQYw6k4p+mAwCejErRoVUpy8wbJM
7INL5msK+RtcVjtNOGOLh7aYNV4iK4VGV/dMFXgz5qHDpNw7os4LoGL/MesMTPZY
Tj8LBfY2DLQXJfnJbrypz+1qE6blHGziWWeaDUq7fmRmuBlnek/miIeCZGzdJTwE
m8yoR460PdWtGlUfFcH3dnZJ6lARSJPu2SSmbWalNywrbpZQMrei2Ykcce9dj5Cv
mtCdjdUF70I+HdTuZcITdHHqfQUG6Gl1qFRzIAnaXjbMa1BCrKvl7XR3wMxWT9wi
P1e50vl0ACeUx7tP/WNDd2x/uWd59dqeQ6SWqPsouDk+W6+suaQsyd/0e+fIqkRk
PdbeWmZXo1n2/pIQDki1XyKa3G1dBZIoj2+E/DCxpcEStztTvubvgm19ISnHys2D
+I9SPqbPetxeIPJWYYPW5kseu1JWTqcK3ECPuXHXl4SL8CUxlrIx6PeFCfpJ55Fb
UEoA8MqIKkg+qZOzL08qPa2DHOdznEP3vXGaodNLudkycOxN1IPKmqvKv/zDwQrv
uKvICz4iqLS4CEZ7y4B3amnF3WOIjPdHvawMTB8Sb3vtDWkk22dhxWiEpfXE7ine
bB4f0fgjgM84O+tMtYUf8du56+Mr80dBUeZjyGdxei0RTzMuypdOAjVm8Rl3ShS3
V2GnvKyWnEKCwXmZR4SJbx9mmWt1rafKTOBPswPMbcXdTAQM1SQeIbxT5c20sta5
Jc6xrTVIgArtrHldi9o+YlFOfDnUJSLVJEAQnKKpXhHb1Y+AHDg5a267dghtsJ89
BJF9MUschk7fbJmR7QSew0SgmMYVwQgXaJh1sgNcBEpo66t/55R1Mcljp0vs+CnD
AgwD7BAPAkOVmdfMZ8IDGRKf8XJNVg5A6J41O8ciWe+G27nFNi6azy/mtSIoZkbj
qNbNx3PNuVU6AjSS6NiHR6auzRggUIONANKEVcLNOUQqN/lDVk+w0tLAYzi1EtXr
2EdAZbxZCWeXVIFsNZgPivXsRBKS5mhntRK31zSSoVIq4HW9XjCpVCH3KodROQCI
ZMCBFhsPPYXlNekK0QzF2lhU/qVQjRxgAfg+v4XzBQU6LDBteMsAZSH1NlyeGhT7
zYPApVCo4sJtWDbmrLnVtifNy7qhoyX0SRFp7htGzhchwaBMdDlZuE2UedeiLVgf
uy4vSwjcSMh7D7BvJy+jHlHkp4i0Tz6DRdQ8ws7f2SZDaT0YjdxtCW5/e2tq8YfZ
mFdrzM5ZXoybmMmPvCc82iMNhvOueODdniBjTmRVTs8I/itY2F8wcp/nBlqzRaw4
aokgTLw8U44Pv/Bk2TWTzL55sEkVbTY5igrqYrYqXmwnoKqudZbpq1B9qCCB6iCZ
XLcReuhiXQOn1pzPb4+KaQepLI3EhK682YBN2fgQMx3hpxDeZjXIlaqRxG7LQySN
6P5QWlEvBoxndUFbrC+2meczlcbv/SZ+saET4iuH+j83lae4onAsYYRBcul+nCjW
OQ/fzNpEB69tEnTXm+JhQrLj5V1USQkAdzPoZHs1thyWXQJy7JeBYRnLbA23N3jq
/mHrkkpGaOGfi3py9coFM/E2LuRqwAuaOFLgCn5HZVmbLX28fCtHxQrBkJG7pfDx
XScAc7Iwmps5yIGXZTlOr1rWFMq0r+pzkOll8MVPW6IQDDzSBgchjfSavITwCRkU
W3ePcVW12f4mMsbJ0RhTT1OAV0DdbGI7Etg527nacLNkBtzTMb/bCjfr1fbo59Pq
f+nriK+0BVBmNALWnujYxzhT5dbyF0iaTBEr2GVDk98kaGnhU7xwzwDcigY863F9
Qs2cI7QA7tOmh7bPLNlkulvp4Du+sjzv8G+RBOumfHLhyZuAo29l6JR5k16oO2Zx
RTBkWnNg8yIyhlAmvVpqJfasbFaYqmTvkQBU4czXdYGNaYuSUOlmd2vpUaqNMg42
wOdoPJi06X/y4JJJN1N6NaKYsPMN9kQd5GqXeaIBwRl7L9qG6r9XYqQzM538CyXG
AAxLsqg/0Cvx0dDh+oE/H2BleaUesjq6wLVIsMPdhpBhOT32YWsIQZXO0p1rRSru
WlAzZ2w/BQOp+fwvOj/kLaHOhZCALbCy3+PQHbQetru4EFqOFIHgXsQ0tOMfcJty
VR5T2ezLEP/9JFTPOk7Msj5DsoJ7bFnSrPjpO/F5YIunzr3aRM92laEz6H9QW7Qy
+rP67JwwYjEiR+zys56hftjd1aDzkpB6XNb6Urrgw+R1rFA6rcurHf1hm7PxtJ65
hPFhEjgPsOM1JZ9D2VuVkBu6l7igp5gj+03Euhu0YCSqMXLAET4x+VR6MpigEs8s
6wP3yvLIYjg3BJO71RP7fiKZlG2CvcT9VRL8VncT6edbagueqPU05v6SlSPYdzR+
XjkSnXGkir4nT2FaCOdTSlndT3AAVFymMUKy3Unylzo9eEJVCN4sK+l554DKiJJ8
xNo/+eUqoES/n67MLMXjN806Y7vD8PM87PoTvC5offTxm6nn3GOfpBsnqvbuWBhd
jxcNTG1sIaGU9sZE7HRQozX3kTNhLxUGd8r43KGaKiyIKLu94b3Gh1NHjdkO6md8
MdJtX0YPxFPTjkmkLaw6Pfk781IpVcClfHtJfNUh8/fG+i6Z4UJkXk0yyQjG4YSb
mQXgGr6T22DJ0Mt/msN/szAoq66LeUftnnDRUsXyrpujn5+GJOFyUw4i2yY1pWCy
MxC3d6INIdYIHUx+Tvu2wdNfG3gUkwo9ZyC3ktYbmndAtGW0XfYGHMxYjEYZGdHt
HesdPCORm9Q7zR23SQxDYbLZPQ8adGA8GPXCKudNjKpR/o5n+QsszhwqZfWQT7x5
jwyn5pxyXrh2vIR+QU7ikvfGysTvSlBeyaCAVORUqHZ7vaQcs/pWwajZyT+z2I3d
gatoUUfX+KrWxUFU/16q0XKjHDYSIoaQNL3Jt/tddrZafLzXKlX6F1ruxzXyQ/Oq
asecHvM9Cwb/x/C7VOV3hUjAPA6OgtZeqJHm9y+tVQuDyqsC2wX0DuYlUl0ynu+r
RTWglQke/DSK/cTjRLxANjmNhSdS4qCnKCW8rzhZiN6B9+fFcwL3VGSbQt324uGv
M0CpBiDHBN9gzWD3F2eOnqcTz3LOt+LmlNwOC6KOdG724oMkSSt5mTJfbRM2KcWC
72N+j74Q3h6rwB0Wbti/ANv5K9eFvzGjPGjk+4B1G5c9z12T6kSHLdnJjVJmO5lQ
pLr40jEe3/uRzMqAfOORKOxv7ClTOqt6poOfjKWMY9R+/fbv6WMANNV6Gjllvos+
z3Rt2oeJYeuwRukVCWLL/qAYy0An/Ig84rZpmrC77Mvre1lVhXT3NiBnH1KyC/d5
2FZb4KMish1wToO+CBp3TifLHCxI40HZ5SPFNZpjQvHXMokG6wHt+k2VlRyRUGky
ZM4t9mh/WIj8ZFGHxQB9IhZTcpFh2nU/Zqma8D3cyFIkZMkCvvfIkCw6aNlvuRZS
9I7jj/pFy63BBzB3kVMDEP/wUtub3tEHiQqk72SvBnHa6UD2Y55Tqkl9p98Zh+GF
bbA9hZIGH9jeuRcHcR2Zc8cjDGHU+jwMVgNuepDHZYyQFVhwXKl/OAFE0NDLYz0j
1QT4kWoU2gflo3L/y5BMxZINr1n3Z7o+gThBryaanLuQcGQhvJxcThlWi0321DvD
7UtbJC9G/1Xx137mGSDDfax+RnIhJcc4oEa27DHoetRhFLLjPA62nHw8HvGGqDbG
1lS2aUmC4j+0+0cULh7MgRL9jkM8JoNTgiPTsHrAp08WhW6JMSHSX9lLma7Ir84a
SOWpP9StZ3R/Of70CBmxEoBji0dD5qp1p448wN5pkdp9BJbIj/c9x3aAzg+vL/Gm
UJPMXG9vBeTw16zqNGyzs4ENHSo8DvvXxJRcjRRwMo7WkPDm0K0z88FhGTBzg0uK
HvmWDi0NnUXZL4un4hWqq6JpexIvNPyJLbFiwQ93zS+2SDmcUhADjfzJpOXAPKqy
bwayN3F0OZ64s5L4MOo6t1+rwl+SGjHkxkgaLIjzLQqQj3PzqOrzwvSNHMrvY2lm
jMbzKZ2oc6yI31XoYGCYOKN73UR2k6JLPYZxTwrFPDSF2zsa/BkeOM8Ue9/Ten2b
uA1QsTPrY4S5HaL8/wgEq7r9C82qFH6WBSZfKyw/M7WhQs80KiMVhyUc50rahTBK
v4vAvUZefxJOrRTvMiRgLfAuXm+rhOc9iWX3Nt/BnDVyLrBRTxstygHSVMNB+dWH
MQ/n6koi1g9LvQGLNy8x/0M3SL2s8EYZQ64j927OT0xrC0q71caO8fM8HLCsC0fh
IFfN0bDRUCOtoRblZsPiFWGhgXjBzp6qNHSap+0wD4ndDrEkDuRKAhLqfadY5TAo
XfGOFrj4wenNgKv5mLjY5R1yvoGAiFKKUT3JdjPVySOTMwzIJX1KGRwuHr97lbmZ
Znzi56SYgQAlACtykQQvypOnBW4+EvCBPrjhV39RedM2HOZQ06/qurctstLLX83K
JR+WaQbb5cO7rb7tdqfVPjxo2ntr7c5r5dU11VWrByUsJCbpVn6Egr0i4UP2nldt
pMkS42qlZ7fQ1oVOtcQXwOOdHrpXTUCccb59QQuymFtOlOBi4plXI2TIjF5rn7Q7
GdTyyMj81YfRHT+XYPkYfhYCX7h+BdKYay1gziGSWhmzXLHwmTdbHn4N9kLkVgz+
Nv7Ii/pIMZ6VWxX+FzFxahbINorVU4aNDx9dBBVTeICnsV706XzCcWq6gdOkgPio
dmpE6tjnFUEKMuTTAjFyOg2Krcfszen3HtUupeZPfY/9Y04km/AUjvQG0TWlJjta
rC+k2ZdI36ng4j3ABpaHOdvPUowixA9XvuPjBcvWay6IoyTtsxt8qzmG+zZMlcUP
z4iJ37OMGhmtua2otOU5Ic7o0joy1CzNhTOl1tJUgY7O3CqY66okNjmjDMjZ5Fv4
IefFDMGYbRzPL9JMmIitPykHDjWxXN26A/FlQ4mERINwsw7fTwRN7gdbdiLMY+0p
zRJd/bVEu5UI/zfhF9z/47duWNIe6OSjuzzHaFWVIqwtazOWw4yC1kpFS6YvkW2i
zviHSvJiaDWJYjRTYzsbi9Ta2J5O/XwpRgVJ8dAS0aVO1JCXkTcFRw6Ik989/ZRy
DvBoY9X4fqZkGBwZAwCBgzwAQRMe+4eeS2XUNzMeBqhyEWtE2LvLrchf5x8ZkTmD
wFbBVdjYg1laogzKV+ulzD7NXpZXTQwyYh6H2RrPV3Nb3kTeT2al6eWhf2gNQou+
TJ4V10+f1TW5O7y0qQEdaIJdGmCRiQ3M5YLd1tdOhUwH6IJxxCAGzjYTGZXoYD5y
QeUkHjTOILwI1yePFOJbz8bqawi790SMLD2aiXqheeALihmVhWamaqCRY8Px34X9
2ECqCfVd/MtPe/FUFfXwE1srZZOPPXpgTb7TacTXoSQBPCmPgzaX6XY3ywQ5q7SS
e/5Iq1ap19KHhI5guTlOUNehKTnk9Bb1HTkP/N4sih8BcoiXXLHPVMGvgGfKzZ22
BJPllqmCcjgOJezoqPQHFCi1j7LR2yJVDTvrk/nz7O95QNugOi3JYVJPSeQ3NY0d
rgO7SJ1Iwkn+Z6ToKA/rSz+D/j1ElIaNNelx6NyDqahL5k5dTjdVZISliRd8P27q
iQ9kH5Ptij9OeuWY7TvvbdIA16J4hFPOYyyqQ6M1n2+Phgcou1T9vcTuthUMl118
CooWLsujoOFEvsMQ5/tVhHbueu8RU9Jl5S39ERErRouXDr4XMJPFBGkrvJqy1xSN
Gopv4cDujjzyS/DLlrgdpoHEimaoKDX6jF3hQvLKrR1pRp0WltlfjGFolmuXnh4v
jWWdOMFq4d/OPFShnwisU6pyXrVuBExEolPbHvFvl9/mvwokERYN6qignPGiUJm4
3OyDsggNw38jgmttHgz9oZORJ3EBixGHlpPAeh+1vRDiObTxMS29poOyrqY6UI+M
WuSQaivkvk6sdflGfP1lEwZ6y7gDzfAWsiVnCpC6K3xmF1bq2lZoHLpPHEuOny0t
lzOH3GxqQdUNrEkcFUUv2U3pbRZEN0E5YcPjUerBGTOzcOOaSrUjXanGZk750qbJ
MwKnp3l3q39KGt0IexaO8iNMipSg2QCmTA6zTnD6QrnbESN5WydjQnHiEFAJAJMo
ILDS+G5AfJ6ols9bZclx3cJusC6KmHctCVhVqdMvXcV9xaw4hrTATARLuzAYq4lr
3du9UabJNapRBYI4T9Pw7SnZgxuyWOjZipYmlm8rw6tgKr1WHYwACv4UnefRTxDI
MhruxsYNiw83qMeW7wBce8/AwRRoX8lP1h5gLMmokMrSda/cykjxwQUxS2GZITap
SGNc1+OBpiVXTX7gq0HhRwWNHcwEVdpQlwsSmfYMPTDNLiw2IRrw9+aO0sbpxVU2
YYHsu8qjYFuqnCS5/wHADVByByE9xsOSoaKZP6u/PUUhq/bpZFYwgTpVlFA5mhce
s2mPRW5ueLbqGETawz5ABOJdhMLa70u7l2KexvlUk/tgiJG5RgVMtEhkdjFlwsL9
xaQN/K5BgMsbxzoGU/muoZK1g8O7OV6zZKNFtHkAZl4uqYURQz/t88U6oitn/itA
PzzHVWyOux97QvE8nNx4gTKTKYXEjR54gVkbZfQxVRvjlm74nDM6l6yLMYvHYFk7
ZCO0K0AX2u6ephwNgxNkGI5V5irSXeROGk7hdA8Th1iQvi/MphMFZDBlf6ObUwWU
rsCr9C47SlYbLRDsSKnEL/lTK3MZKL8Vb76mtBL3Y8hVPERkQ7q1vTDj35CC812D
Gpz67BzmKsm5Z+WF1icH1w==
`protect END_PROTECTED
