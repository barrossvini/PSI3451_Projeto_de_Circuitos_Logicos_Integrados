`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
raUPPyMZrkT5Zzb2UgbNITGJaR4TOOVZ5n4n+Ur1BdHzTtWyEqlSPOqbarMq34As
gDBkOd513b6Pvs0u1gzXXcyYzm+io+wrSbLQWxeZ53jK7mzr8C3I1u4f0nZ9ueki
a30N22BJqP1GsI8T//s9WEOTNmKKoP1GzhqbgJauB+pLAGy6koK/xe9bhi/5uEaQ
AypimJZsgvrkNma4x4FDM0vWa2Yo0QBnSOqKlLS1ZolSl9O9Hp2DWZeAtpcEVAAr
FaKW15oi0YSiepkRPEWTFSsj/jR0IPepbUMgX8/glBH9tqyC//wDgMvzFldRNgKz
c/Vx37Dz7k/RO6Yio1gR95erQSf//TuXoshL5HOnL+oWMdNscSUFpwWEXLUezgMy
0TCSk6gJxxrMiD6KuVRmKy7TB3bZujEkX6pwe4DHAXnNSrKZwN1o9fEEDjAC8s1z
Bo9Qtc1bXlqmurncI4tscDwCYnc3pc8MTqbvbq24b6V2Ew+rwBQ+G2jbxQHFcXfh
vs/8hrPjIVtgx8kGSaLQbVpZFa1hHff+nmJP4/IVTvwIw09qCVH2ABM3EVUjM6H/
tDzzNybcId47JnhA/vjL+zUzjEV18xFQoUH9pd++sQ+ncHz+M/SgQETLSCEiqiu0
nJchRtHiXZY8Ybxu/GOV0R9xXXrrOOR2r+BwW+JqFo5Ny6/JKw2G+CqT7xlsRIt0
tUKK0UqbHwrKUMZAWIq3gW2oPDFQyxbtbGflBlfc9nnJzTT6P9dUO3dKnFBKkE3b
O7YW3Eva2PU7N/qfhqkeefoUR5Yum41DX325XWQbR7+x5D/KOmHydtq6ZonmtA4v
jBl0dlyiQ5RFl4nC8+le297KQdTdXJi1sYxmyZ1YD1hw5cdTWXmENtDMUwgGzCrm
fsBKU5EKdQ55VlGZkv5t8P8pdPgE/4Vy3043XZ0hYLxHrpBcFT5vsZRAe7UUNMwm
IsP0islKb3gO6X0O1hMC/4Yd9DftLDDLKGfiYP8sH78DEWHJIcdMUK+T87nzvpqy
FaJNcEc56q5I1xNQ0hJoM4aldXiBqMMRUAWLfJpRurx6hxt80o+4UGl797ATbq5N
RqkQ6WUCs7ZrmRenb4SzF1Nwq6EnC+9Hqul1Vv83siK8r4nk1VRdkJZpA/WVEFvb
b3tTVz9A7RmiUNR5ANqtRTYme9bywAuimttqkFIWembX2ZDD+E6DcrABbksDK7p3
g8heZu42Y/hmC2znXL8sv9bpEwkAw2RPG78MvCLbSS2PQPMsp+yoV257XecaZmal
nURco6bjfXE2yhqfUaJIbzDrGFuBFNV136kOPfYIEgf0wn+BRjM8WXB+R2RMxrf+
T5Roo0aMjjA7iQ9VzdbkqI++Q5wg0DKGJoewtxao+bknyS/LDfk8vgXO/u1SLCXU
`protect END_PROTECTED
