`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZwO6/Yn+9iqxActeBnV5xrJUUU6lCkvBmagsGclKo4JweqTcD5KqDmrxncZq3JS9
29Z73wcASHy9CEp/sPR0Kq62YFC7BXuNbC8/tPJaQKrQd6wmnn4NnQe+jqJK8sNM
85WAVp7EcMFlXnwZDvwcwfJNQq1Y1z6cD5KSHgg7Ea7doKUtZ9cK6gBrr/nIx2c5
X6mZ1hTe2kI7ndEekt56DrLFDkK7b7tio5ryL86RipbpgIOI1+Dxb0PnPCWs+frs
WI0A8lN+teDuAwZ9jLYwICAh53uK3xA3vVJktbKCmAZlrimv8i8oWCeSdM+Fo5Zm
qh1camAjqQ349flmnk2XVgz1oHsWF06HappApKJUxDpJny7T9NAPo+f1m9hGMRmH
05z3bxNfMetk6pvwIXVjLYg3LXp4YWmpyxMRJatBM3OwEHPfv9QGADYtRIYTY8BB
slrfiJvn3c9vCj9tVnIYQTM/ispwHPKh8wGc0ucCelTVsFouqOyOComWr7MBnBtb
lSD2aTfuhTUiBulPptx16A==
`protect END_PROTECTED
