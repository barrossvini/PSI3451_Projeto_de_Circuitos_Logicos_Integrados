`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7+NwbBxEqwaopZ8/5Fl1DlQLuTINHguGwAxh+qFDM8MXZyK1k95xoMYuh9u15zXh
sl5qe7/ifINDbom5GdYHAdG7IUwcWAJ9l0h6COStcwd9ESW7XsXsIMq+CuARvFZU
XLmJLKwPwq1VWGXIrctIAboKAlvynwVWZczkZU0zm++GW944EXMjUUbXd7+j3l6o
g9lq1zBgbJR3+1h9E/wfY/9PztCjghj3Wg58A8i4GF1zAH1+LmGijG0g9M9bSZBL
dI9Mw+EGuBBOaIEzV/caR3ZOrnajotWf6e81d/W2qXGTt414QBSCiBbGDBZK1QZC
+AHdYVTXG3ir2Giad79siaMgzuQe4hFk+/IEy2Ygrjq4CLA2lSRlBY1YNn7SHhO/
F+KQzjBzkM/Bf3+M83IrR+OFzfvNj5fuqquibn7sx6mOkkoWIRzjumw75lSrlLhL
8F+ryFH7rTxCjQs9NmCS9JbekuykogMMb//RN1kCbe4IUhDnmjOT3bC+gdiC0W7G
ADP6saxH6kpWK4KRvPK73ngV24Vin4QENMvD8G3FDd8kCZMsn7E0mE+sivXhThO+
mhHhS7lUQv0yEDNHXPD1VAzO0dwQkqSAFPckiVfrxtZHfWzIQOvW3LkVCaoA3hKj
xhXLizABdihpOUtBcOrbWlf/27GgKeF1+jxqYzvLuaftXCsTfemM5REb4ptoFsA8
tkcrywnHIk3gsQ+FyAyIEf9txwcra1BpYzgScAITk5h7w6k5p2WH27YUWaK+Qqh/
fBMpPyQxvcZ2CSWMqWACT58QAtSDWeT04BKWal1yTJc5HRbljaMKlb1zDoZG8L2D
syumrYCkhtxLlLX2FcmnuJdAA3k34vZ1Ey910aguUm3KvyidsDcfb98Say1TLOfc
C7j6JzOPz7u7S/cS70zY1J6ZjEIZI3oFJFPnlL5fSJ4XN3tRcC7AqoWvN93n0dLE
/7ElnMwEoZ2L4h3frbGTBdluzlfY6jf2Qi0y4YgN987wO5Z5iJqX4F6QYqK//KqW
YKZkRGlEEMYyq8eUBmlD5YdL+hsyClnZS9aAaQt54cvUoWyzEuj8Eo0qnCSFtWbN
nSFvZ4n/LtLhpKc9fhlPfCOvCnl26aDy8bG35fYoxfqnI/UPM8IXKNz8fe3ElVFH
qGoYaF4Dret1iiuBiZjikgq4tRJLSTpZVWekWRZtHCZepXeMPJqYooW1whHFp0Pv
MBrhykO2qzdhUm1ILwwEyWubGsAxL6LK5kt1zj39JzYcVrC557KeHbKG6wAWjHD9
IPq6ntNA3ktXjB1tgGWqOTArP9zVFcdSg763YDGBnvwAb/bo5HkkYB2kqZkjrpRE
SRhEkqfBgwTFqnNE5EeYgy6rDJi+EzP3EF77u1TOJPdq3LQKmq8E1ZVFxS3i8ZKD
0VQ8moiA0DlpS8DpIUxiPdP2AlIc7zOFrEh5fWtClJQgKGKi7M9PcdwbSz0vZKgx
cgYTKkK4Gvjr1qYWnEvgtsWP/E5pZBTE/2B+KkQ3HAc9So5tyg1baCDFEwoWDGnA
5AgGWjAPEauAgLFiUNoasRYR+Q+VMlCBaX7G1XiLXD9yX0gO2mL/O7i49VXwxnzz
kraJFh/WUFHFnjzscHgSmPzGCv3GJj80Rl1Bp0hkd/+sRRq/ftSS3f4LyDf5iXH1
iKJaciG1T5ASDZN9iixUvdJJq3JRpwzBXVpx2R7hOq8tGeAui+bb7pbYzycbcQbR
hMlekmB22s2G2v+C1s5c8UWQnazZmtOoNyDfironQZm7haDNwmX52x4Lb6tNoP8/
flr0ruvAMN7agq/o6grOCKx7Le0jV1HRRqFjk/6xCWRPPzXbNN4xu4hO9EHJ4mqQ
dq6KP+q6e61hzg7v9wKXXNNgPGdMtX+mcmb6ANzrCM0bq3WPjPzUKdYVOBaUNVnp
oYR8zoiAT0bnGUrkLVxDGqFJmqD5sUduvP6OEVyE4pMiJV+N1UqeL+gPHNTd/bMX
6s8Km6iXKcOSwIsEWetFHC+mTUD/Xht9YiJHhsSWn+9opZWKsKmNovZh24UNLd0O
QBx2IMa4ggnXOh8hJg5ScsP5xHPHlFLFnJ23fCR+JTU9DKWzSqNB+YHm0rJ540qJ
McneSPe8PyCC4Un1uCgG+8PsMwwl1Pv/ZClN5X0/ysJB1b9X37UiiE4DEn/7JsR0
EXhZavsxSROcAPfdloHHShtkPNNhS+4NpnYLELzQlTpyifWNgVpkt8IICuwTHYZG
RRAbOO5hpXeGzx+Ivs1G/fY+/G1lE//jdYPcV8PIqgPsmP8yPCyw2ztp9HxXbraZ
yJ41xYF/sXTSOfYVyZo5RE7kXf7kadzvI75xzw/HjEEIuxSJqZq9u5XPPAFBxmQZ
EaSYKKzzVny2Qk+76I0Qa1789bM/29dqE1AR7nq7+STWSJJVEPtEOrLXNGtVonRg
skcSS4MWXMeAk0fltD9Z/rJQ6cfRbgvM8+nowawX5qnl/J9fpKMOpTgGY+Pk/v7/
VOFH228zhxb0JgjW/JhG9J7oNoItnTg7verMOCDjxrsd4n9AKoisRpk095ViBtPr
rRxbB+Zx4Af0eRihUUjzhQFDAgF73WiF9Rl3zT0bt6FWXKLLCAcNvtZ4qStDXFqC
ZA8f5Re+NoP8XMRHXm8tUlVp2RVzrBJVqzzw8Q3LT0dCFIUnTzKc8gbhndZQ6Kqy
+2hRL+Q8yr16gS3qi6aV3pA0qYBsRoIeH2kHme9M8g+xRLghDQszA7gxuXEBD/Tq
5+3Ta5l39u1at8peHCyX9QFjYZNNZ/GQc1F25tWZxTxXADEODkA5aogAMov6AW+U
woemGNtYcDCcreVFc6W7V1oicLMmi52SehpCt5tSUoX79nDvezQKRI3To6PnvAkH
lDV3nyGF5valG+YhQrch9L5z4JL1VdwqQ90PMvTEywA/8H+ZyYGkjPh1+tXmQCgo
zNN4jgvXpcbQpJ9F75SRLNHe2ZDYMw7pap/jtc0RitAFzQlYY7TsXf6rFHmlgre4
HDvKiZHFbg3YvfvUoIhQQPm5NGwg3zNcJLC0X+tq5VEm1tqxxan6/id6VSgz7QZq
M4dqz5lGg7mXR4RusNQmakekamqyr0cE6J9vq7W3Vx18mhS2dUrmu9NWBp5xO2N/
j2hH8rQsduPScOu114VhKW1BglzKmWTsd5L7UCO+e/AKidkU39ja7Bx83cXVkkVD
xTgZ/rVOT7UR6zUPNkdEAnv7fxHJt5GebiaeAT1XaFa7qqBekVjoDKHCuYiFwNVx
JVosgy57F9vv5S62w696k4xCk+k69mVM0ahm39XjFET4S3wio2y+aXPVvTERfmkw
vMlNRXBUSb79EigY9mptk/ntNSLJeMLXPeLXLvgEse5Sq+ecm8hUOA+QWyeuQA9h
QUcxi088y+uEncsi+oocQRGQ6nUP1nHU5BQOGdE5MjuBXmg0XC+jt68G5Lfx5/Fd
p1q/VyBaHLzkFKOENpXVtFu6hi7Lzqkj5GzPZbrtO5N20jo6vk0Ta40Aq2e7JXKf
nwdtT6JnHdfrzM/3HEAw9Uvp216RIXDW9xxBs/UleeHwu41ftye0uIEF/LGGySNa
Fk83t2mVucieLC60g7SgCVpl/eIrnzQUv8OsW8Y5dcNvd0L/Sz/g6tuJNiLpUjJS
zHHaXu+x3c2h7JtlOTsuz6T0731B+ghLNfnVTjsAKVhW02JsdOoziEwW3+Z7jTyF
xKLaJ0Zb9eG8l9M8eHxMMgQkdgMwEhDFKsPd/cHMoHcH8cfSx0UbWZJsAdSAbmKu
Zct9xiF+1uO4FR1Z630zEmuoBqt9H7nMyR/KQ78hgHP2IsQPz5COzGusdDpvda9M
VV729aLN8vtphde9f79nyY04SSSVIKNl5E1DmNr6syY6eOjCVpq96P79Hx+vyqpI
D5MaoWj9Jt0JBz7MkcPAh43jH8JmkBq55jZL/YCOkBGeUFwYVxHUysSvHP+5QCzd
eQ+VxRfhc6NFkvdYZeMMA9ErPS4pCiFoUKam/9dJVbtNOVUZ9hBnIA0a7D9lHX2F
4m3tdnwj5309aWW0/zzPXCu3bfp40I6oqSjrWuNi+nUrzi6yv1TwF0ZXyBh7CN1V
Qzt5/poq5YgnyWOma98iTCKmKgTZV6B1eGgggzMQCu0Xw22PoTcvL/mcLmKXHLUZ
sSA6nUozIppWGxcd7gwHkv6cBlsTzoWaBlKK0gbXNgZChAHN40SeG1m8hT41mw0v
RlVyxQAdzZB/bCH5RJQzKk98lV8oA3ZZAt/RinwmsQM8n1Pr23pHetJz9AIvKT3J
ds96OxvsukrvNSTde0n3nkFJHND+EqEfnzj76CGi/AlaKjBbU+l6jh7p8NzlbxAj
VgQzk3958IHG13GQavehpFAOcO98e619q6TYNnFKgHvXVP2sI55bmhqZPzkwzBov
7QNFOoT5ggK9i+gOC0u1WWpJFHDQ94mm5/kL4dxL4c3WWYdbUXGWRdx23yg/aOt+
v8VgQyOu1SbxsjSP/Ad0iwX+qpQmtmle/WYAX6ddR8QNecGSCDZ9jTR/PA4cf/n8
8rBsu6sQCmpChhu2F7qT+3p9KA+wpumpkd+J0tIee4E9+B1guvCUjBJUZilWtbCB
WeBZPOrVeJqhS5HjDNnu7w+00Hs0oELEz05FtHHgCk3NO3r4sTIr6tf4fdpf3oKf
bKl90cckyCgvJTEtL/5xRvC1cfb8LC7casgdQmGGwG+uOnsQGbDrzGUuIWN87V/f
eFxlgP1/cyuxkJ0m+h67aBoX9EJOdRaGTDkXIhCn1TQ898Ck9aa3zLc/SI685QaY
lqPlfMkDJNgObXeMNLZmSz+gp+FMiwHEpOvaJNIw48dMVf8Dx+Hyl8UJS4avVCpc
muIwQht+FzPyuLEKy25Q2Za5ICdR/X3JqH301eZygflB3hnQnjEEZFPIqrK9nnt2
SXMWW86D2c3UcYo2Gl108hJbhdaQ7tpuQOdBnnhWnrgF51nTVtJ75IKK81WSxsbQ
t6zpaXL3DVnflDl3lrnA4fokIYNGrbf6Ox8Y8nFsK3H1wDFh8lMpZY+YWVsA73Ga
S/8Hk36hQrK02W/ilEGPlemHiMRUR+n4SS9q+Q5Lg3XD74TYaxgnipvU5/80Q7tm
ewb4JE+TjrOdzRuZKlFJZswFmyjBJ454cAM15j3pexM+clBXI5sFz3VuQbqTMDAm
mAN/CgO7lz/laobIa/AVxMCjZQypbriVoIwXh+Lu6/v+DxhRszrv2VP5XZQkQfmj
yQ5hOQkhEQanBXWa/Ja9U2xblkKoXJfKWwayk9K+HWR3Q1rIKNazYDD+7/rrSe4r
EWuY6lvoeK54h5Wx+moOqBaY5B35k4zKrybW9FRFTJpDAHQtQzIrQ9y+QI144yUa
ezsKDlt5Pa/BQfz2tuRi6t0bQPM4WxiRuR1FP6PrJBFZDroiRXjxUzTaYi5uuDrg
frbZQFnyct/VuH+Zs7HSOGUmz6XNaIfn0pr+8JmvFioshfBeWwDUo9OhpvMdPmcW
xfpU7AJIrBQOc8CYATIq6Z6Y2zcqI8IIm6bRz4jJ7VVie02g0LcqALZ8H8e9DSpe
JxvzpEgYAfRPuY7f2z+/56xOldwrdXR/Z+SY0btQJerYkzmakSwZQig5C244M4+G
I8xlE7BxMBkjGb/RQKVN0R2WKHo+72Cm3jWxh8G2l6AhPE+skPgdL26BasHWKpot
WVMx81uh6cQ4ORLY5qHZGxDY8hgU5KDM+6xaxNwBpR1vjB24IYDYIz1xfyaW+wgl
OGUKgOXyCXlIK9hnXCpcaAT2Jy0+MHN43kbC9vHEBEyHskOrWVSZBmx6b3G21Opr
GWIpPnDguY9rbezHmoM/z+ATIR7q6Fo7NIgGLS10HOqhp+EUiHPj5b7OhKKFPC+5
hLQ4i6pv9b5PLZOD+PGyszzNfa9zD8Uun7RUJquyLjxA6o/1zhIjUz1x/Xpsb/rD
+X+R9h6AvKpBjME+XbDgTBoGg8TaS1gLQGSbc01QCxbxQglansnXKhi3IkZdXAfm
PpDLvnhDyPuJYnxDFfPyBn+dpVvRdwA98bCILHsSKjFzlJD/AKzU8suvrpKWqDsB
ziVQWKNvNK6uufabzuN5WMBIkrh1M83cQdsOcJtbg1bEAVWdT29BR15YMZFZfxBz
w4wYx7CIvdYjmpVzDq6pdgMWqWyY2qMShuR7Sf0jvxaHY5mQSeoJbWz9afPkBN0o
QBE0/UWsWWZ0zB8iZuoFnN08rniW/h/alWpJDBP57GqKlYXqxMziOvKC93TuP+0d
focFdqldCcRb11xGF/FdxHY0ESKvb/SWNP5BJ79di21weiaOVZfQzCmxmIvZm2+A
7affrOjSnDpEHMXZYQKsHKlDR0vcWHQZ2kUiEfER93M5MXhKwn1Rxc4U87v84Ibx
spfIcmYLZIIQqh6hAJ8+XPVP0utXIvphMLcz1cKPzoVt2tUMAlDXxodNuH4bNGuY
RxebJhtVm9tGTPEJ3lqkhdBcKN6rZ21pYTSy/AYgpe6K0eLGEj05L8kZkZ3SBR/T
s2+m/9/TDNFA5CI7WEotQrd8ZlHuCQt1uJaC1i+GuaBpCitMsXwGs0V8OiOkMzne
XIP16SDOJF3oopVHZIgyaRbXfpYwwqowGO86UpZA4+ZHp6doBGmBS+P5/o0KBv2e
apo3x/YajcqgsM5QX1Xpt6QT5/Uhs4htMVl96c7zTTV33FOqY653fGMofUzHEk7z
Kf7sCDAutzgPzzM3wlV3VWlXqngvz5+HBkBIRv22oXrc0ZOXjVr0TEYII/8sNQGp
2XeU86+sq5BcCqbV+yGZODCjmOcqfvLvP7qg+OpRJp4KGR+8s55NFeTwPwZi9Bo0
6qYuU1J5fWu1cJGIqs8MbgB+IXK2ypr6NQtXpIIQMdrrZ92G4i9pMtsz9BdgtLqu
m9J+7d15HDpH8qd3yUfcLwavtDfuFO43n6RSxQpmFdoceYooocAnX59HpemmgpKq
hKzC3FViRDBbZsXq0luOnZvGo6yyJNhbOpwjnapqiKthNcvtKTEA49F9MqIxzOjg
YTjClkVzKNH8sD87yARrMqgQD6qOcFblj19Ha3tBXPfFKMewmkLKZNxJ44WoQkeG
3mpkrz6t/4nGLajcGhb+U8YZDDjrrVzfSHv1yAmHdwLoyT3dEBBE/yMWgN0rAgNN
k8UKPnn/PStxt83ZKThJiwOruy5ikiSKTFhEB4RySseqQg8tM21dgewEv3KLDqRU
x6iSIB1LNqjlaq1Rbr6hZtcNnfkI6f9LO0/vKEkwx/K5yys9xJAxvv05BbqaVncb
kcIxvO5kiBqc+4uqKzKpWt3jIn2ZAi24YaFgRTSTvziBji30w2DTHfeB1wgs8K0h
dWXQSM96wQw5zbyFRGdcJ/20/NbnFIm0dIQqVRLdcbn+jogC3dsbx1T6wHUFWfsD
Dk6qzEOFBs2iUniN8lcFlA0hhCpE7HUP2UzC6H8HNjQXzdfwZY+g5P0/vLRJE5IK
bWAl+fxaQOKQf5DIpxrQ78jW1KYmN8iby46QeKvD6kcPAapFJ3gXkAEcYL9sEZSA
fVecZHkkh4aFMr4/umBZYl0DqjIkb+B3zBxPc46IermO8R2Psui9G6HyIYyBbNlu
EtHZPBGFrQOIUXovsJD/hW63d3aMsKYhGFPPD3FipdZpnRhEtTCvSTaXvW1UYVv8
4HBVeUKoqGLMe3xoORWtvEjPG4viMw5Z2JJ152rwbvS9i6XBy+Cwy0QZZTWS0QVe
gHfOJ9XEbldVxu4MqSNX5A2OXOk3bbF6BA3ttwuHxf6TNjZa09C5ZKaOcxXJpLim
YjXKpgzmZzjmpbQHjhiGCeQ/kuQbWU6X7AOlBhuv5JQlOHzFPt/uSzRbgz/axOm6
juk/qt0rkcAPq6m+lLytY1aoXu5f0TPtS6T1Bas56xNKNiwylFE1prDxyKFnEFEM
TLFsLtvo54YN9XAi8zATojrC+fdUOxXx3mRXE2gVoBZpv+Iuj0QYyvcgAAcPL4ln
ggpsEp0ZU7CXf2Wj5LgE7iqQ4vvuPB4Kow4iD5EKO802TMcgeN5wEl7FaH5I78c1
rianV+7aAn2gbXrElxzlDlDU8ocjNw3koSB0p08tmlqQrbpMIt/4MT02IhPsKfoH
7s0wG1t/sXhRZ+Tw0ypRyQ7LOCW51M3OQCTinxzy2ZaeyPLtPtUl4olNRBZP7rom
47r7TTJlxVfXK/9k/+fosUzmKdFh0u6tL8j099nX7WP4TH3MO2hBm3qmnYm9s5LR
7I790Xl/TGOO6kVB2u+x62aHQUupjvIStjuDn/3TKb8z4HBpBXMe6h5ZpuqZfRmz
N0qCbKpbTt3CdahViNUG8VxJqYI1kxzNVrMxpVD1EFLZJ1C2YeorjjhN7+krss51
pOlsgsar7XF0ylHh4m2Y3Det6+nU2+mcigD9QiFOgzhN7smRg51Ckgkar/RBqVQl
WvxUV9FzUYabhlt2FJyEIz3smS8BSvMKpOpaWtPKRNw7bh9I1kHYN737Op7FtVzY
81AOhMSgFEGe7K6WCZYyXV5s3LMDMOJwciisHj8gcnlvn/pnA9pz5NRCXrTLgz+N
W4RX6PqtcAIeaA/Qtb31dm+DXoO0Zl2lhSVapk7L+bTtP4dY/NGywVV3XoG+f0nI
tdjvOu6S7uT/PlMRdVo8va9bCFJZwRb7iQob9LUeGNCqJLwBS4Fodt03BMn0LNjP
Teyekal/BC5B7/P2yCk1Iq0Pc3OsssgDAakMMhNtgKyDFN/lDk3oDDzFu3pMhYkE
gFfgSkg27evsAp9+QXGVPPQw999d8rRjzxyCuMlv49goihTAZkmN1RtW1o9iwpJn
ZzTch4+3CtCAbR8bZ6QozPjsf/Sc1T74aT+zy/XojIan0+AUjeSCp6IswOfBPDtI
LvB0bORL+vopcPV03UD9Zb9QrPaEwut/vio9gtccVeUG8yk4D7+gHTvmspPbA5rX
0u8BBpaKKHY6OziLmtAkkwiuEF29jK/DLIA1Z06BNvTGTf/zTkyxYvWMRdtWSVA8
FvbxT3t11o3UYVAHQc7OC9nhsShFUJ4PsojRMTFqg2eqINq3b4XaDejUdFvoPfhH
ImBdbmtCwxl1Sg1moVdR17xvIRArnqMnQ4LG+U4E+PncTJ+4Xr+U4j9Br9NUOtZY
kK7rFYYyuyXE01lI9uR7uTFqdDjs5RkeZmnfXwGyA3ZGUjxCxcGcwzG7kJgFz/Vi
INgXc7XGgmyuIyD+ZPZJhthJNxKCK7l/CuK/voVTDTagRSLlBJxDcKTWJDgwW+EL
6OtE4DffRy7jdaXySXTZJCzXVhzwdaoHm1T3kbAizue27FnsVFpuap/ZyVYvfDZW
HV7Vm0XP2JOdb1xMfBiWAxDj+Hr0drtpJe5QeivH5GaEUd9L4pQEI9h9+Z/G1hzk
Y636mfusXlaifR+YrlKaAdHb3w0rfG1nYCI6YeWLlLGShn6+1508lO5uHosnEWxx
dMCuMvxdFBOjO9e+5onPa5+uVqSeFNpbOZEB8GeTPASallVCswc+uC87wdjD9++o
ZYrwHMub6FkltwMuXxbk0OyUytGVfLbBfwQUBIYcxMVwLBDZGbaK1R8YaDchjU9z
q0tF9fqai8pOENWqnFJsldwiSCRhqr99aFBLa48Sj0Sk3JZQ6/lu1bqfbPRiYIEL
7Rqs9PCoVmf5tNaeDgl9p8eXvxM5+rERo/HPwkWBAAC+WayXtSdgZY2Z8s4X04UI
xWeu8dbX8j6FOizNG9ojLN/0FggSVSVm5FjTVmAQtubIO40q4aIlK4aNI/uT1tbP
MXOtcmf14YFXr2PSG2aYBdSOrOKWhLgGs6bU7aFk2WW1vYkBHLUKhLFUOaRQ2+/W
wVwuNXqMXF3Bi/4/fdJ2KnFsE/FUktaYPr2Dw71nXrInnzKGANZMJYZzeN6hVvL3
Z83GTadB7zegrM4eEM43x9rSSUsxsEMCabVltObmX94AZL5++OogsR/yfP+GaYtQ
Gj72ow8EIQCoy8BhVrRCK9OgKKZfXZKvfNVbGjLDSefDJvEz/czBKBsO7vcpbCsE
M2VseBl732BuRzdMHcVAC3DWdKottvHv0SYvfGfGqx0IGmOCSewhhicVgbRVwgiY
T5C0+pmqtMi41+Syyk2GjbGcejDPo2uVx6lnRotOjaIiVKA7NzeOM3WjjVoMA9dm
PEODZoKQi50BpowQXIdK9Yl+7Q4ioLddOWlj8AhpIH4+z1MXDqWZruwKdYIH58XA
iu70duVg111uaLFaSXL7P8M/xbz5GOSnlld5l5sfDmU4gEG+ERC63o8B1za8inKd
JGD8PANVFDZ1an/UP6mSh5ZgCHOoVA8By3opuOVNxlYXKgObtYl8a8ir32kLBHJD
45xQ9G5ce+t1rA1eO5nnfC4/SXUFjRULNlG3yxhWMl8A+99oOiC6TuH2xW55oUny
FT+JpCvroiqjWDGEYsAU7Mp3LMC+8I6VrxtoqG64nyUnFi2kIhmWnRliP7RX+3Yz
TIi61CF1FKKc4P6igjJ28KEWBUhRGK3qwSrVHk5TYCZ1lT2d74PgH6GIHjrTCSx9
8mr6k4nDj6x1FONTwEXusRtyr2Q7gM/TkQI2bGX4B/2sghZncO++LysINCG95r8U
+ic03regHayZ4Hopjf9oLoPoDCjmV7D8glgZEhdeb+6iBvaJumxBj7lz4jNv7jsS
XLetM4QejK0zmV4NpUVu8TM4zF54Z/0DSfe0nhMOaVcaBjuzK1ws9KfV33a/M6Ju
dBKHJ2+VAEUdXsIgBzoFV7IkYs8yR4EYgiblNhIRw1X2ajRTNQ+sLdGV7rzEuX8z
pC+ZCkEeLl/HE+PMN+FGMnxfBEYEiuk012rpuZ4AlgbCO4uepYpMnz6ZjCtoeCNY
PW3hmIuispqmnzVzdy2KZ2/vJgm6dEAKR5vf/YFuTI1EK0CHRbxs1ycy9CTED0gw
0R4uhGJ8BoP57551Aht8N4Iu64Wr1yKRHyToNiAALJEjW4jVuRbrAWYrBssVTAfe
8GtcuIoGWtwH1FAvtksU13/ZDW4Vo904LrsXX6DOLz/twM3SJVk+xizI4oaqFImC
4/cKQ0XTgpHv5EbaCXhmfhMn17BTh1OzJHNdnf54HyicZ8f8G6gvH2fZOA5Goilc
9LrMwe++R9jygf+bhbQT9xRdmJqde2nkv7/glACpzooixAivBwkOxvB+MkjWYvs0
M5qsIbOYVYHbrlOabqg2onm0yjdZ7/k9KmyyfyhFAlVcrYE2juFE0yFFDnpudt4w
+xL4kKYuIIeG34Wg8wr+1cDycraXEdLYurv61fw+u/mAevGE6viwZnvJpNv38gCJ
RZKofN7zAyJRhX5SgqCgKL/VhFSXg39KCObD0SPskho9YXmx2TIxZY98Ag8UEU4K
UvsX968bs0j+zwtwISOAIKxeL+G1kFwqncJx1jOiALDWp82MbUZBpA5lYFqwNYy8
qByUjOYrBDFKnFMFHPqzRgLJNWyDGq3/BNlC7mttjdQhvGco8fihXYX3/1J5oWmr
I1PsAImU0U75zDEgpz/Sg49n96rK02A9Tv1Y1Wbx9obNPfdOOJyhA9RbhrI4P9xV
2muOQT39SY82ubyrarCtMXR7Bg7VftrmIeGRSfGaCTTlbxn4fd/pUlxGAljcGuVt
LXICng5I2IEpD17mHwD0h/xMODhOqulkWRt1cb8jKlIFAr1Ciq1u6drhBKA7KeIt
gRJERl2aW9m3V08yCgRNA+LSDmfbUlC09bkaII9E4l4M8fCdXANcibcsqK3Q/xD+
0qUpTE5mDj10mDLJ7D9WxT3Ne/b9QmJcRNXh7d4hGVW+hMUe2DpYQX0peE1aPkJb
WwQGyBqnP7HME8FIPhiPx6hfymV2/2zsHYu9ersdiQ3rIZRUmpuKeiTc5y+dmnqd
ONCjoThkO4zxJmBjBSIUOSS62v9Z1wuQSfAw1Nj5b4qnUu86RZUFLIcuqKoAi+hw
hGRpcfU67LtVcuwrrgoW6XIKkmLOZ9pfeBPOC1a2sIDhaJ9recOEPOmOtcwv9Q20
jR7VITWVeVMyXzepMM01V3syNDOI5rMjggpUMpSr1GmQxY970FMxXJCBy0ibnm/f
CaROZjGoJg6C7AN61Eb6JRpk258foSbWUPpbYbYM5dAZydFElEVg7wfAXPkdi7D+
M0sVPtOrBtpOEJ0V0VqWEKyvvLNWB5UzLbO+SeopfPX/H45DXhjpzBAU6+BWcJsM
xjYTHTsaJ5fa4oSWTCluxotRSyvy23FLaeEdKRI41x4626PF+v4F7gWOJn8Vj5Lx
OARjmbsMUrFPExe4c+3oAk9lGhpMJTnbeLzBhj9m+wHElr21OCoAHxc3bJ1aT+Gq
0v2uR733zcDiRmf8l6oy2z264YoasSLCL4IfwbuEniLEgjyoJK8YPNwfhsmVmpKc
5mUuNNKCN2mAUvcrKL3b+f4XXd6910j9SbBG2qdb4UgHslGnpaiB1bex4GCAWqq2
P+07UplZsQPRrFYTTSBzNG7Be6rNMj3Jh9qddiWFnEWbv7/5O42wTt77ejHxlEvk
5Km+myxOnqGMppyAnnQ7cPZy/fRTpmToGRmSGdsLK6jOxStctjwj7yCtopC9wtzC
xftIFo9ey7SdX6RdMt5QZgGISueiaP8UjZd3scEN4C3PJAgUaWkKqrzHtw2xzJ3M
ZgDTtXWOm9hinbjtdNlsrr49WB8SHWdc96ohU1KX3uO6bvbedaijt6AtyWJTlgsq
AYCbgsJgrzzo12D+w27VrCPNKpHMFN4txJdxWjV+f1YfC9koZpg5opeuVSqruqj6
s/c7k1opzN/VioQG2sIIZBnMcZejFMrWc7EK4I1yKKcPDC5IdT/OY64+yP/lOBk/
C+y3mZuAt9+n3ZEY9wDNT9PPFQsxUiTVxFSFvKxYZR1Y7efw372xB7JoC8GbObIg
UF8WmFHaOYSS0dHlwVhKAkt6PCUMM5ZTjRjsJM2Y2lnNvYgKLHewwdLefHB2JARH
4SqTvrW40egUAmF0Q/kqs9z0/SZ9tYfZN9ep34PTqzfnk1nyGhJAirYPMskuLkBw
omaHO2B9C1fgp6Jb2a5p09KrOuzqmEayKgaYE/uZBYEq1IwR0jVZTUbhmOTH/2CQ
DuDQIVPrc0Q+8e4unFIpVmfpcK59MU7DGB9CuZj2VxQIQYYPwUK/g43ktO90pDHC
NpelEbpw+R5DfDHyIdcrUVuFb/XeMu9up4wlqD7k0SILgd2duEmDmtnPO50Fm0f0
cuUFOJCWh4tVkVprwWkAjKAMqHy3lKpkt+zwLZkApa9EeLWbapOBGYMVpg78h5Kb
+3xvXHzIPKLeS2COaYLIzGcSSVVbUlQNn/GT+s4tvfd6G8CQzQRUMLJ49wV99FB5
6A5jcxsQ6+qPCt0hr6wkNfQH2WsgV7x57phC2ec6vpdKB1g2BNAByXsbVE/8Vm55
3ZUoai8QHut5GceoikCHIT127bBfVfPQxpPLdecUuDKCASRlzs/iXcMh9ON2mhpE
UiM0eFBXjcyMzqkqkdJKbGZ8Oqiq/FBd++fsP6GpDg6dbjvaZU3yLopdwE9AsLKO
3mP6z5GMME+hHECLxreGvA+KqQ062bxF1j5hIfVhRTF3NT/NQlOkFXSaO/4Ueoo0
YsRy/KttNUeEeXGz8H+0MhejSsBGBgeKFHZOIALkBatobCouYrE2vX3vy6lpINHc
ApHy3yyURlq+l6+OtgNU8sCP2ag2ayB0u2YXoQsacMFsWgTvjzm/p/DFaqxH/0wA
Zi+Sp1bRTvwg0UOOQ+UCCBFABsD/KRuMGcGOufjGOGYwVljnquFPbIgEYiY52SlF
KQnW4FLjozWx220hsz5h57FQqspgZQMAauXGH/meDd6/KxcxVPKj+Ondy1OmqpWR
rPlszuq7vHiOv/hzsIGDwRSFcHNotC7Zk1aFZduDP8hgGxgXNhScAZv/FOpUxxV8
cUMcRP/xRMr44xMqwIP1cq87szJCqP46bZZVPJou2bhd+K7GsrQfUiwDgQGKgBBB
2ci3nmgYxhqE0o5iysWcoyR9BniJo0e+pHGcDbDKbqtj/8sHax1ZcZFgJAVnlRff
lSwzpM22w3DHskAIFy03zdNSS063MatXlpFJPXsE4N0CYZfcoEZdnJVhvs7p66ap
rr+t5Yeir1f8d6cgkLmEOlFXG9ub2/CAP17ghJ4DTxOP920BkvvZD3xupVsiQCj8
PIf9ErafTPtuxHBH0a2C5kk4b7v9gwu1rM2ql7B82ESSGQxQVc85Rxs86xWdwpuh
PZh4MlPm70Zwj40VIC8tc+7wnGIjUheqCmTdJvrs2eanonzhEosWdibfmtyhPvLJ
DN4uPmakAw+n1yCiP4S4LCoA2azhb6c1MyRMLkRx3pzgg1BbGGLXndBH4YgGgVHa
QeqE3VCHkRIwz5hHrWxflnSsFNjiJZzBrXQdNR4/dyUlEbTVzUx/q0TrCV9a5a3r
rXaArt+EZ+cP5iMsokAxl+yjIeYV2IomJcFHuRrGlQQjSqC0QlG8ydlKQOcJjuuE
ejya6z/pIA4I6sDEmVy3AVW2vR3/DvnHp9H3tcuZ71hMjaGsBPcteQ1pHK9sCdce
75141S46iiEgNQb3BltaPEAedyb8c2eOWY/skuv6U8sHCz1nhChqoLizamRoaTxW
0L+ynuzR2B6ElDlYpFJIQfusAdTV1E4B2eIxNtVTEgVoMdQ8YweZE+2p8uCxBEQs
wThybTLDF3eGercTLD4Ab8+HewmuML275DnWeguC/sfzYuSFByRMLyQ3xgGhViFL
ajzlerksGzxB6kA2yQyK+52v2deOQFkztDeNae4Th13a6GwgvR6zLs6anclrMRz9
NQ2WoWNna20g5IahggM617N2xgPf4LNa66+4dCvX5vPmwECCL8pEtqrUcFGpMLWS
5DYwMAs/6F16WUgiMhY4AdfeajFJ+XQxs3x3c4ZkmXyScHEnNImQjJRPAFi/4vFb
h0zshIQc1HcDp6J4W7gBoABh49ZIKmMg/LbuO3B3AV2B7+gDJDKQezSxLFWu5wGr
06mE5NdvHi9KbYmX8CzJ8Ry02EZCv65W8thG+x3kEW9abIescq8FfUNzAJQgq7gK
OEd4HtjdzZZ7OWxRD+4yWzEU/4b67hbAfI3kW7/bsAqF4AAGcL0BsOqCSUwse2Y1
GFmcv1w01aVGYNyKF+ki3gX7tOsbOg6gSZgAPOE5DZwBzB1usAc0ogBfbDpwluaT
FJN1xbjtOKqibW9kPT9AXetXXuV7OLy+sGpris3iTFavVAuwR7FLZHYuY1wYXN7T
T4qdomBgBHT5CS+ZGUsf2REzsUNuOEqUDnoY5G7LDrhHmqqsDp9BDRXwbrEO6dED
ssKXch0BxyFx2KRGUpOI1lX9jzx4TQ/1Ppko1f1xMg8GpC2/pdeibl45VoFquO90
fkh4v3DZnWK82/DU7HlHveEPDVsMpNiLe1zS5Tnop9WjJ0+LD/RUdDSSNkKwIcTk
B0gLKKKnT7d0or6VzVMG95P3/kJ52BCqh3PnwmJVUitH2bFzvomk2HV9IE3wC6R8
5cC/xTOt7XqEo6ckoUWiGstfGDRbxuWIZznjY8RCdMdaJtb/Fb0HDXyUCebvMHu9
Wha+KUJC1Q6S/oxSOiYJAlbycdr78LDW7Q48iDLJXPO7CXTBd9WOEXmkNi5fzt24
vGupEAqaijxXRcj+gdUoBUE9uGDLOcjEfvdKPg/RoElcjKcaaJlrIXosP4WEJuLO
ZYEz582plz0JPvPlIDSGIxnsSzTNXj3T5kIitW3VngaiKbbd+1/WRjBj0OfaRWLc
EFQ4NXAtwaopObEeo+3phYqtIcPeVIN5KT7YBMe0hV6kvBShoXR3xbfv9CYc6YDx
B1v14kwKmMpUHj2EfQlXltA3BYnomMxHk0v5AcDtwe6+qseao/nF3r7oWYGGREFv
nRHrPtzHdT4U7HHrm1FeF/wgbdNUijBdcOfegcOwf/U2sWNFDz205Mhhvh/iWQgK
FgsyhDB7Wq0J/xV92veNi+HYfUyXd6GCUdwGV+vTKtMDy/akQkmd0pYEro0NyBA9
zJ+zmmyoxFCJKdVrD2Y9TG3GnioWTnF5mP1mrSW7M5l3haFbHwo6oejq8QTbLSb7
uHgE4oAh4BE/BwjHJqxuTlahfLvFTUng6hDy0x1oLSmgsCzyrw+M6I1qqPuI3sww
ScLwf9AuIYZt8qhDBgqPndz9a76ZxcrT/rxm4zYdFtfdKLOR3gd9oGw/35BzcndW
9C9z0opy7voLeTM0YDIg3iPmH7PB+v6nRmuDjv9DoyJ5fMNBhUVCzda89qsstxwn
HNyGfxNfaVBq2yvbkj8tlEufPWWCd47i5paWvDDTxZqGcK/QWIQsY7u9lc5Z68ve
k5048YcSXftcgx/cRIeTMIaaSqQkfK79xRn9hA6HRX5TCZlPEriAwNPknShpD3OS
uCqbrl9YglGfrrC3C07Wcq1gIX6315kMXnUFdpqJBP/BDdgbmtoei5q3HzXLkmZ0
np0wYKAIPHgJarhU2/su68wIOnWOVIp550cUkI8zCxhuvDi7d9D1CG535X9x1px/
PzjzGKaWDjGN2G0k8BJ0SAMWnJ9zFagyz3mLvAoezHBxHuX0wP0Kd6csdHciqdPp
/Wpjxcwc3zaM6BkFyIXTPgcyC3JBkaK2RRvyh4GLwgMG1kZid4pNqOkRJuO1fMYh
4381cPOXaS1Zx5Flxh8BrKLJ6wyHkWOoWoFai3sBcAEZBWoum4MqTrpy4hhP53pN
ee2gV3Q3eIZ2HxhfiVq7/SsrH6n3b8JkzWBtdKWRKphRww35v4vR63OVSknas+dj
4sxegFW+LnjE1/6BuYwHWRbi1VN/q3GNf9gDJGbNjaG1u2ptfc2OgyfdChCeDgT/
26IT+R75bqgXnPjKXcj5jCcFDbjpqY0/w6mBcszSWPKe/NWIxkpJjBJp3w2Nd4Dw
5x4hio4ilRia7MN8X+d3MdhCrjM6aU1MOQkMOpahCnyPyuKqM5txPosP+w/or77c
g/YDHiTd/kPnEBAk4rav8YanIGipXKHVbSlXPm+UIhHEsqYnRMyQCZxQp/bg7xXt
ciIKILe6XbOOGuhxEj/kkvZsHVmFKJQsk21rmAXgWFAUM4i0VS1V9kEvXPNlsRo4
0LVmXJv9JYb2GSdyK/OuZLao1oTKgMnhQow1h0nY8vPme+NeBPeh4h/ETRucWlVW
upan0KIL94WecPon0XSciGH412slEso7LWCipLl3BmnLvwn+9Ef48rXJycqCj5e1
bFMypPVulZGpJ3ZrQyJxeYhvsde8VT3xpMgYNr5cYHi01jl2RJhuRFnFi1VoYLKl
qoLyoKNIGOrntSmNta9lCt3fHWtGQEp7ZcAVWRrAJ+0e4SifxjgAV7sW33QdQ/78
Xvy6qYVGoB6ttlbP4rj0ctaqSvatcqApxJ5fVLrRUn1QgFVBVeO+jUTafQkfXZj/
99DX/Qb0U4FvMQKB3y3Gm2+pPeEzd0z446s3mPCBfwmIRp1fsQSB2Z/q05sAC50A
IytEI70I8Jy3nAsvrURkXiQQq5TFyF+2Hm9nct+j8M+3kU+3mtlf439BY7BqaTFF
gwrYSHVI3vInDL3fHCzbapx+6LAQBUuUYsfpC8MZNxOvAjiDnlrI4Zki88ODBdWC
L7+EBN3fZitC2rUjQC+OlGKu2L6DcniCU3NIPrEo0hqCujRdbEdTi9fuwnHb3iqw
WsPX+i2r/n8RjjPmOACM7da1AhOj827zMOmOmSSsi34CDI0ep3m7u0QC1izuhugK
2wLqA3Bz3fR4t8S3jBq/AarCngDqEs1pLX8FthDVlnVVIXKTWIHTv0gdK+kqQUZ2
RgF/wW9xPoqtVK0nQEF+XjAZTLfJh3mkBnuyxBL1P7ky9m9ghV6hD50Z96RtXCP7
pkNWYOH+gLFtzWAzOMS5CvHybxgu+5HQE9T4KLCuH05aXSC0jFKri+BBQ/TsXsLx
aQWJL2hq/0YyHXgtz67CLgT06eJ+Alb7exiP60vKXJvhN1ZXTjNtkg1d8T6Aaerl
UbRzw1QuMnvaiFT3oB6ZJaUDjRC4YwpKaeiC9lGYMelP4uCZRUQNHfng2GK7E/bN
eDNYk0bZ3elnwYIO4zX4F9E/Fw+ZWIYjRPEyaup/HrvTwW/bgI1WxLD7FAe6MmE+
8iKqCQxQSU3LlIxeKVxyzHEmk6fbBDcHMVPOgqaFxlsbDZ8CJh5FQD0U7g3EbE+o
JlEQprw9t8cNJTxkmLanmcSUpevQ9iaMc7Xi85xg+vdQ0ZNYFvQpNIFr7jXAYgMj
Paz+GjjH5dQ7E85F6OzUexpwUrAxX8+O0pRvI/bdoXR3dm856wwGb3u7dqRPrZBr
MYaMHXAF83UE3PM7dUCKTO3oW8lcurDyQVzcaKVtbgRMuUJXRTssP78+TSAk7xFE
VE55c87EvtZ1k3tcWnJPhQjITgmcRNZ31jDBbHq4G5YK/YZuYZo/klGHuWbQUXF7
CXqLswZG3mOvLIVw7vR8Vepe+hAWh+efA+DeZgmGkpgRN32h6rhIM0Q5UUm9Zf6E
WhOruu252Uk4iiBpAiz4ybHAC/CzXp2k/QSosmqoUgwjWrIRLtJNlhfyibZp9SDu
ujZEiBLAyHGeW+pGniM2Ya+h0iDLiMPF7RehTg4nhKpvEJipQ1wdVuqw8iJMW9sO
APmt8/hqksOu/lARUZbGayeok/AQZhDWF+EwZ624vCUm9SE3nzZaEsYo7Smnuw67
xzaT0sjgv26Np9Lii6XFz5TzS5JYRnIH/zqlD5qvQTSjozhrBdP8Bh3QcVxjZvXT
lPoAnbWGMwMhHKocbQYT492m3Wi1O9M8Rq+KwGVObdZUMCQlDqAIg/Af9ZQHAvMz
myhLXHQmihQAl1ZRF//P3aL/pXLmrn3CLQ6JRUda9Mr1oFncyGHCwx092qNw8uA0
eTWrqa3+QfMzQ0LTbpYAIHPko4lyEsVmjrgpYlD3zJLUicuP/dUL3DXfS2lNz7Fi
zgoU4r1cRhyBDJ2Nm9yiBXv+vvVpzGxtF6uD+NetHETCe3FbX8F4qFCLFDJA39Fv
c0/Br+XlUeJBNTLH+enhMYjzeXYt7naRDfblK9r07uLZdEwiUdU245Cw3cBJ+Ghh
jzG4D5UdJtaZMBJjUGU8LHRw4aQEJUAbvk9K2Zod3TIkrRcTlTtk5g+r5WYDYPQg
rJHE98eNU3B/IEk0Iuu17eat8aDdksa6FM269JqZ+rRkrnOXTeVgj138Tjhd9poz
THbTxpundbshwoe3xw+mACb29/GAS5eMLFunUWKvQpBAmox6CM/CsKXGvAy50KVR
8CQWlAHreFNNJlay3uBMsi1Vj4K5MOWOT5+BtzV4Ye/LHsxbUDKlnKWi7fhAbP39
233FOiw5ZC5ofLHWT4z4pQujudU1eeTpu9QcxBDBGVHEN7FkOhLpI3MdIDtqiz5c
FlW/ltnfpwlHs/Rw8qvi8Y0q4mo2zxI9ziJiy7VutGR6KRLTc5MQC8bBUgqw64GH
k/9Ql/wtzz/gq/uqT87hETQFaIIJxeAuyzNz6+OLs94eLAv6IJdrcizWkGQgq6j6
HgxEkaQQmww5NadkYrJ/PYjCZtX++OqETC9m1y9wS6MzZ6JE4NhojBqdlwgpiJNf
0N9INXpY3EdAItwbCE4YWLS/nlffZVH86MJfEtsn0bDJ2woRG/Yo5gEeSL9T2e/q
jBv64C0RTo8YkQUJRNWQZY8s0Iz0JSH7GXrB8K5X3rF6RwSFrV0kPjdWuGCRV04J
woKUhS3oAbihsz1NDkMrZrM/AHM7dAtFI1WO1pG2qOX6Iw/acXiSMxaxHOszUNe9
Y3hczcZgD3OfEAjlII1A36tq7zJ9d/vTX6aasTdBtld+hI48FCe3Iexu0qkXVl01
T+tsjmZpTm32Y3pdlKaZER3Swhe0gEDuj57QBm8SJef0vicQv4yx2sraNhaexhhI
rO9idE2L2k/hrViBslOCyEemQZo2V/2fYYApH/0P4U1beJQNU2nbSA9kAyD4z2FK
4CCXVlQ1O1qfJWudRlefcbwTMKP7AIAawUeQX1Ws1wKPR3H3Sd1mrjI1zMR5MR9E
hGztqraLSKIMH+aZcw4S+mXi1m/X/J8XsTMywZfYmuy1d0NyNiJWCma/jgEnOrWO
1HLSpEQuEra3ZeuE6iN+Fu2EJTWdC81RIGPgniZmX19XUkITCP93jTIcLz21yooC
+e8AJKI3Q7joV93lR1QM8AsW+3UeexFBKgebc5HdCkDKb6k2obd63qgDA23W8RiH
vtiiATJ7LOaBTtaOTdUGVPONKtLzOGHT83vU/u79KKEZx9CyjJ3oUo/vYU3645iF
icNl1S7SOhRHM/xDtZkIbZyhCFDq95f4s92sQDlrqZT6mnxbvbrbxOrhNsRni0Mq
1uxON2j1SRTYyGJpxNbLfi4878XRggdvAik3tdNxHcLdCsdJ3jrX05JsyiHvYqfk
mltKYP+xb3Ox3vvrE7oFcYqczyLYDuIxC9wRSQovUYBRKcToL5fM6qmnCsEWdxcQ
7wjbJNAKqudBHB4uW7GgGQwIi+R3CwxPu6ipRF0nmzIB0484N6Ex9kJZL2247ESj
RqmudaXNt23xo8yX0KOskjOIjpsKwgbvFUk0bvj94W4Gka/9jocXNRoq2SOy/CTi
IuenZSvFRpjDJ9bXpWXPEIp8817Fq7tPvmyWIh61FV9MoZUVBw224CULfF563CSZ
0iR9/HChuw+qqFK/bD3wKz9IcGEn9SHGnNc9wKSERSey0iMs7F0BE74dSOzs5Kgp
5J/yweIQvV91tToEfkT8KyQZFUJdFjuoCPcj4k3eDB6Ry9UM0VNtHV86/eYjjUrW
F5d0Y/8luzu49BFn95k9b/DP0GXwMgE07jI61ooodQiAuEWrEbANHtOsEE9/FyPX
BPBIP3ugbq1ypFYZ9YRF5PxJG6BQga8lZzeygvtDk4lJ58rEQ7dHGyIL9qoiDgqw
7jvxx6bkcfwgzi7Ko/2U5tD6qpdBHuswHULcUDebdIP+U1MWtszBIZP2e18iYVlD
OlNANMxnihZ3eolYmRvvSu1RwUTPWu/IB8q4YGhUy30ofa7T3mXLwddrP3sY6vyq
MeScOKXHH1HfgMoJRPs+owhjfLewqgTrx7h8j58l+qy76075juzpyPqGNxn7fMxR
bDvQ3G56U/2YT3Q0+k/2X61hbYguxq+y7wV9dtSwQXzEHjdbaG4mjvrMIG/0cVC+
qOg6iYjDzXFnuTxInRmcxOpJpFQXnQ7IBQ7p9dIrqaB2Ut/exiOjoCV41XNy7327
B7Grix4jvxgknGwqcmDX2cIeXHV7zfnmAqwGOkuAoFTpBIHQOhJxyulcv8y+YkC3
5R/g2IK7/Fn7QF5hD2auqaJxZ6GEvESbZxC3MGo75SLxtTTRb5s2xYKQSqS442qx
WDrGep9JCA9+bsVeXWpT7Vmmk5dlpV+WcVeFhY2j3GodpDtrevf5RWmTFqFWWyOo
5x5dV6IxrlonugbkRsGiSsu5nitFYqMNxUfvkdy+my+/k8EPzB8G8KdtFZgWuun7
E9w/gPFh9kqMvwimY0h1276aunBc9uO96KMfKQJGXBQ7C+0xBZnC+IiypU5T2IGo
sLgVO4hJld8jRY8QrjMQXsbRugYk4vCq4AkQFCCxaPfa6VuA8MfQ0gt+DppZAVhO
/DOVdpY3IEpD4m4r7v56NOu2Xg1asXqr3/1BA+XMAuCI5DFUzzpSobzD4IItVSZP
QGI0UPfP8tCxlXpqgc06VjgZrtDdG7O8KE3iZRMH7AjB26pzjd1thLrjseIrqN5R
FrrQRgb99qKF0n8kKU8qpJP1DJNjpiJqSggnI+SXkWBMmB1tpXzHKpQBT61hcG+f
gIGcGx3U9Qv3+zWcic/Q9lD3psxCjuGycrzl9EHkc+nJvX8n/NWH1rc8G0Qnmp92
0LmWxcIgAlUxmn5T6KLibwl4M5kKfazChnH9MaRuBHN0/tVaRyX6etW8hkVrLETL
wogVDEX/UbYO42XS+r33iK8+ufbdzSRKpf48jorfEnejTtIMgpKIzJa9a5xQSHl7
GoT2hzFxKZqgpEDsgtAFtxjP5YiF8K9BZh0veUxT3S4mJfbTfm9KHHKhHlElFgKE
0ZfstHYd9asEPHIiUReFU/1xCWbpdjdGJn21BgId7SBSfPKwnptHj5Pv8HidxSkB
bnJ/CWY75oHnbigZQ9QDoDLB+phedEwW+9I2W3PdnfC0nmheAa09Q/lLMuqR738Y
UBAYfHNgInE/CO7w/OVY/KA/qqPEQYk+zbJW7Fkn5pMZOBXHTXdGDSjhHwdG2j7w
symbKNhAD1Z+u5oqGPCuHPuENn28/Wnlik9CyMWXxlgiHVE0UYB4jv5j8U7rCAl5
uxszRQwAS9qIL0FoiLTU+rRRZLCTycU26FLfup81a++/SLsu8W2wH+wtGekJK/jq
xyJurdvvjv2rC+NC8Ztpd++G7MN8isPY8nKAOJjxHBKAtWiK4gs1XuFA73c+qucW
qN1gMMIJsKufMddkH/sWWTrJVRnQONDa6595VLffAB6OkUTVgzmVH2D576dtq1C7
jr7SQ5fzk4C00TpsUjFy3GhJaOK0ubSKhW5vUrTYMktdzKkKTdLyY17wKI0XNdRp
izax71MrIDx0Bgdi0ig3LWjd+TsXH5dJReDyNa1M5keLdYksQQEA8NiOt7jgdEPU
ZirCYpWquInsR999bAJInlrUB45keYh3sG43i/AQs+gpOoeX+dPKqaaSLc9rzNtQ
A+zhHsmfNsq/4tD+YpdEquUHGyNIZ5aatkdZoLRA8ejt13tTiZ3hFzVzDaxgLlgL
gcGT7DADJaiHY/bGqFZ/gHIkNfCzLqUrFvUD7rqG/gXWCCK6wXyj+CIidHtiqAc3
IDIzl2vg0M0v+law4nkS8yQ542B44mbsOg+FofQRN51p10nntM/o26QxfgdSIv5S
glD97W6uXjpa1C6fI1cC5Mp+qD7/gjaXkzfjiRnEl5Tbr2OgrHu/xixJe810J5Qa
lbOb8C/3o9v0nGVoKcans0EE7Nry3CFrDiZHr7wDWwF7GcOyd3Y/C6J36MoYeltL
xgp116C/V8KnQ9bemeGhKU3vwGa3b/4o4QsvOnnLgsIKuZDE2EToJJhuod5SRec5
H/DTIbnkPl64A+1BY23qS3u1yScvTmGPFhgf4Bl7/V6LdJM9EEu8wBJjbfLgk266
wzMLrvt1gNiZ7GRnRI+EJOXw7Tfcx6i2MEEGLeEzNj+J4kOi0NUin1GGCiUjOHSi
XoWrRIupFE3qsVz3BkGkBogBSPP9VnKk+xWwwCYem3d7fBonpnblDDzCoH66jQfc
behcMHuokDj55sFBk2NyYjhXBjfgCQi0r3ltnkiMpvUYmPLLwOMYD7DCr38k12T7
Nuuj+7U16akb6Tk4MX4aJGO0JGtZzeGCte15Qi+1e6NDpgoeZjD8w65SmOFq/aRV
LSRm8+FeZ/029HMkZMv+dcE0Bz656vqJowy8JNoCYd5Otng5qGQ5qFSnTV6k+Y/j
EdKVuWNP1y4XBUXhAQNMyqumYdy7Sb9Un7oMuX9oiHfTjcFJs/bspfgeOHjzP7z0
byltyq/HQSw1Voe7XyIKze/+EXxqdGaU6zAqrMGznoW809p+EE8qB+ymR1iP6xIy
p8r0Bm9ehrMD+DQ9OK3jOVb3ck+h7x7I5K3vG7oxHo7Yw44G2c+NFwLvIzj1Vfo/
YZDwG6KA7cJj01KILBQevBWOZYdMi/E469EyraDcxTsh45JMyIJ+mwF6i4zaybA8
bUcsRim9/sdcGlNXKssqJaXyEVazhnkS+1OuSevOVqsWZ+1q9x8DY75sP7IlAIgZ
7hkgIaBP2F6yCPn0A+BW1WWZLvnFIPIjSyXN4MN+HtwNUBhwkoKcKG/1MEMS4fNc
BsfjDvu9DxIZnWdhYIKQaXK9R9Bp6QPH7r+gpP8f4tdcGpmgGf2eKrWLoU/QYva3
Fm9Wwel8iCcYPUjTARZOt9nymg3R0cfHlqT1fSc8Qok9XYmOlPvzCTq4s98yNWnx
NtA8ynJxis55faE1XZ26fUYu6tFc26oQsYGEiCWbVMq1sN9TR01IClIuVHgBIOI1
0BYj4c0oTsV/2hk5qkOkrrZTfBJzF45KEEBSoRH6xSqt+iVBJEKdwic7sloAiaPL
2QIt5lG6UXpax9fIr/aG1xYkYD+A/h/JzFLWzSX46Pmj79KMEjV5TT/QQHlb1CxO
UvRmOtvGy6g+zCk2z7QlWeZ0IgLX1lD0upbKIy4k1JTT46C2Af23qSwtbiAGoPT8
eAHW5TWQuwgeKGf4qOJNYmHFSQHZAisDf/UoZGzLX5TZEnze780Xf1b75Vmzl3GW
Cj+SSSaF+Qwf0R3aIAKsx375rWHls3CeT5QOE/d80Y0GMJsaVAhKCxoXiHGZDJSD
rDIlqgTFuVXC6hGmgvlcR0pVUGqvnArAQBNMTug6bD1qMxXQliFvS4HQhSnmDTFr
osvaux0UZV0VpniIt2c8H5WcThkQmeBH2d5tHIjuniSqnOUpNoQUfiBrj/HYNqnE
vu8tEMHYlPY1tUxv1jGSbMyNNS0cMlOR+1gRqR0tCAfDG4uvrDPXVSWuqk9RGz57
/GSfVdM7JwiFYFiiq2TQBEm/0XUSwsbz4CxmF3uChOi7eq5o14UT9bjy7ixtIR3/
JrvJ7Z0hQznAszkBG0V60wdUOHw7LhmdDVCwKM1Vk/lP/XA1iIHLiIQVvPuNiLXb
S6McGlSwuh345tZ9zm6ER//qRCpnkrt6F315KrHMV5LrSEwAUAsZcwDIn9mH9ZKU
Hjjme79m8xSB7rBtAP33R1D/lOohBC66ZYHVYjYBDxxvIfvKCKcaN9aG+gb7CVCf
YX/CTAh6FXzG1+6nwp0YJPH8YQd0cuRE5H6XJYfnWa1Kik10K4eCjNdRP9xEgswA
kaw8NgsetArzqw2Grk/RDBGzIJiic/AGl4cQvd9PFH5Q58RYPCrTT9oWQ5+9SdNr
Le4YYU30tLc/j154o+Q3K9buSJdgMyM8G5nKfore5cLQ+mI415dW0pQ9GYwG8bux
wjBJLTICyAxyFWElAjVX+4d0k/GdUYS0KpRV6tRi1nCZv1H5PbTyqHe9NgeYse7S
aFgTvBnmYTJe2IrLuPC2z6t9Ip3FFtBLCrOcXesYLZog1HPSZbr0Yyq9hzEAkdMB
NTcKd9cgfilC/qeG/dCyl14pxtzUXKpA5Bi2E8GxkiwqvKUXoHpYsfhRd/x05ufe
Ay0FFuurbGBWKmlEUfe31uvROkIOWta/iA95B5ApnwhG/WLFnOoHVyutjKYIxxG6
gllJDhL1GLb5321V2ZerPVks8yWWwIP4Who6fz4bSxaZrVfNkDhsV4MVxxH8S/OV
mNzzanjwyiNAvoeqZmbKTvw8GcjqSb339d6uW0wp8p8YuFck7bTWwrFv8Tb/jbv1
D7qJR5fL+l7bQ9qo7lfadE8TalZ97APCR1ewpZ3b5JT5kppoWu8KSRQodw/mJFOG
R4B/aQ/j7bbdJ7xPT0SnJWjb7SVb47r14OWw2YkGkSyp0K9NfgNgJVF7ZlfBAwva
NNHAvzFKD8us9/FGHx4i5E+rHljC4wTiM1HTs5YvbPFY1AiYb82mkVGKdNIIVpOu
wHsPB73hyToJTFG9a4MjInzB8DpVEyGjsRXEABJHDYVsRSTYn/g3N3VO6j8MBmx5
xOy/LIV0jiWqWbdIu+EjHi/ksMHWiAkOUd+DgvONK0xF+p92Q7Z2loBLjNqp8ciA
FieoV2sJeSYZomYwWl64QXpdtXTJupAFtlTepXQuPgACoY4AgI0gSrQu6u4Ay56H
ugwIGJLQRn6Zsbm5MAcLd3GprAmEPr9GxAwWANAuyOnqQX99Kz17wfdHZG9F3LkQ
tP21UNDy6TTq99x2QLB8BT/g8BSFqHhGvFc+zUMb3AM2m/R7miCYJR9INu/6R3vh
NbeXX21apZ67LuzgVaMO2/PMTOk9d1UeJiwEep37TEp7yajOB/EHJx97CmfG1jeL
29zt1441/wcLam09kbRnF2Cwrpx6uJgfop/yuQa8MdmwL4ar6P9Vm7e3Z8aG0dE/
wtdGqGJ+wxlauLJO3XCDbnT8sOBQB5UnXQfA8I5G5njCJ/egSMuF5v0bGAm7/haL
62cJFI2oWDfQwPkxCHabXv5ePizt63rQgR/JZlS/n+/rWRDm+X9gmq3h7zo+R9xM
JDA3tOhz+tR+fNQUylnALlVtt9utJhiVWvGlO591bjTqFeVsobGTPokFMpjC9hQ7
pD5CRu7Gv7X3JjRFIrLILDdXqBAJaqtTxJFzrN/05Y4wTkViXdhqGzC5xuroTp/Q
kkvd9OTUKwVQ/nJfoVYpPuYsytPjWLjc7YXon3n8YfIfF/96+Ys5benMK+aQ3XQW
M+XnpdfJM3OwW0Km9Qp1nr2YoQ5ip9v00OwG2J9FcXtmgB9Eoozwp0uawMW1RkTD
LF7i+BxFK3bfX+fglTPhfEV6R1a45ka+aHg49289MZEIJ0iH/B5IvHszpJnutbtv
UR9hOksC41k3wmYLFcPAb8rf4XJ2+DZQudCGL8pOg3IhRMlL/Feu4yIr14rp6qy3
rmnqozY9nabDxW9vGr/CWB6hsjIVhLQsG/Ot6vN36vI+lBqy+gDoCKgUCu2tqh3I
9PPBW8NcMBkmvAxaZnIvZN06UVrMeFPKAY+ni/+7cfH+IQacpYJHvX06xWt+zAEW
F2qoLGq4TOA9Upwx5mAbOt8VGypzBb4YjNuywOw0li/UtVH5gjnK00XMKPu4r72c
g0qRhFz4M7JeKr9QfYp10k3jjf/bNzUznCf0rxJaOAhL3VmOstak7yzsa9WKbkQ8
65jTBlmQeGhxTWuMLpiXTwR5TBoW8psD9ufI7R0cvHFCM66ceN/7d/nao7zOdQA4
p/4mIFvacoB9Ecs+5Jau7k4UuoX60E494RVZgyNSs4HzNBDw4Tdtkh3vCB6NLQ5l
D28NnefCmcNVwUc9gla/0bQWhxW6YFe3s4evP7TaxzKQBitKFG4ifdYmL3wmWafN
QCQxRzCKF99sxY5iKtDRi1Lp7Djdg8NvScysfblYkL/NkCLv5EMPa2y8MvuLM1BZ
Cua2YguPOT2DgTZeUQTn7Ek9tva4chTysLnUDL7TWrw2kZ74LaHG75fEpvTJUMy/
89DY64QQOU4NENBwlPnhWrKgiAqmlsO9DIfFCEOXU4CHN9TApNEU+FiAYP3UnPZ2
v7SXGf1qvN2uz4VFPKj1bMvJ7UNwOmu0/CoA+WftmltJFXPb1J95UR9PQOaqOlQ9
K1K1GfQ7PsRZZb21vp66Bw9DHVQ9rNVkxSuImUFy75FW5fHKG9mkzkfR7EIP0jbb
5HKddAtEcv7NHW045m3I3V5IKkklbqwW+n6HnjtxdJ/SCuZ2HmqKa/EY2hym7CIK
cV5eBN23vlyrVL70hcSNV5XJ056xViCvwge1Pw8gCu9LHEQqBFz0qcW9P6zELrVC
NyM9YTJsAlMuHy3iJwVah10Yg8bq3yMH4APZrIcCnod/XbC4Lcaovu1BhazSavF3
ExpEegYUFwwFbjcRxHLUmjswX8JGSF2kn2xLoYZSrRZdwfXyalLjD6K+JwzTN1mb
wQeh2lFrIgxlVVsM2EMtwz2EwFGF3xYRpXMvz2vdpz17uE1yZ5QlCGjlZSDLZIyV
WDHOI4dN/lMjQGESB2csQy7FS1hwL4E9wPVME30srVqiHecgYNKdA6RfPg+KSxuK
b1ZxgP+kToNZoP/HxW/ofHYRP0zGpr/0Z5NyCT7o9/vX81yM9Rftqhlb7oGbAQs/
zK05YTANXvNUhWL1k0pLUv5ILGpg4g+zH0trRoZwpe3/4/zf4eVQ/CwLNDrROOuv
5t42z7WOj8MN3vXXEAdGi2BBpBtQG7/9utUmnMH84c+DumjtwWd3pAVkEn6Hujnc
sdy47JV2Q3R66hZtbNE9715PpkN7slIHNHvAaLDO6K8gnLuxYcnfj7LPCVyrXOx/
/+HgNFdSf3yXt5Wb1ie+FPvTSFBOWqqqOzCUjtaGjv4E0dV9taTEFk6V4G5PMvMS
NLnCEUPu+QzvVYivUMnb6LPh4ev9SYznyP6oQK0DaLxxbH2uvLaqO7P3pvh4QOfV
E6pTqw7tvjZUe1PqdQ0YgWhf4PGmsQ5CslD2UPxTfHiJSsc67+aJCWb/08kNY1Pg
egPnJIIwuQ4yuDxJKkzXiDXsi9IAYg9Gqv9UncNnJTFNUhWcRED+v4wzw3/gx+Y6
f3BTCZP9xjlEZcopOZLjh5CR9JqtHEU4N+4/P/kLdecmdW6OUaQYVDv6FWz3Urtc
1Bx9VZxB9i9YU3hSajo/dXyZn0YyU4a3/gkqJ2MpMmrkendXq8S80F7f8wSr3vzI
Amdgz3mW78kyr3ZFhpXI3b8TP8xa+gUkBVaz/o1ArG/A32RcsONNj9L/Rtu1n2vE
2YI9fDQN7LvgtOA26gg/8ab6hEqR3Mcc0BMxvEMM1cpagsQz+YFYgzy8Gfr1USIB
VCs78zU1DZXboz1XvuTlv7lNWkHBxBeILQjayeC2JSuHfdS9le+a+Lmafy190wfN
Gofi1p/JOP3SdLOcdUfCxO1wUhQmzr0cuwIHjuCvCuJEm2KhkiFQf6ZIC1QUGcwh
6lohpGzbPK/DDOyjo+ZFMA5qHoGMOlO6rL0MqtB0sH+K1IjmDjHLvJ2p4XPajmXt
iptuEMWsfl0gwhAAsoVQ9Wi7rwxKztXwQnb6avxfR3RNSZtmjhV6RDWsoSQh2fKd
4jIRkmN7uuK1mH8Tmr2wxe+5sQS8aTNgBV6gZ9c03E5oo5E52LiBDcI54gx5+Q3H
rOk4eIovk59vdBFqBuNLsDQWcIk5IjDF9kVZMG4N4XHIfS499pJ4WLTTclSIoH+E
uUFY1NKDCu+0hUTXa1Q7cdhp+3D0Sx/Yjv3pfZk048sEinAPkM352v+3rn9akQp5
s5gRUoR5n5sZlJVfYm/8LLioIp2xvhvBMLn6FMEOEe+86shvnx5neQG3onMo4v4q
2ngIptMtf1JTHrVXlTF+Cfo/gvA5PdH2qyL4a+EMY4Q/DjS5TIBoiTABYnsCCHGY
llywh1D9rIjUvL0OKFnEinAbh+9+btZndFHZyNuf6bDhR9HDv5cheQCuslt12Vzd
toTeYNfDPz4sVYGYjOIL6OIl+Fs98qEXirxUdGAjf2ueYQsTqEjVo5AB3rp4gEKZ
Mb4MS7Yb0hOKFBqYOXnbLbTF0Q6+JbkLDjmYxgxqFAfmA8T2NcRhpYdGSviRjxUV
KdeEOP5RDyXiDC6zNmR8bPwWie+hQ+z9tyjWiWj+4SKerD1Iwbw7yJ68vCJXuKWk
+8ig5B1I330tUWrDwnK+23dqH5gKJPKiQH8u6UGiSn6DbH41Gj4cc4fG1pir+Y+6
XeOTGeYqUAasxT+LZvF6I9ZYM9q4SiUhR/Cim8TX/xs49PmHs1Zf1VyBCF0Ungy8
1khpF7e7z3yRwVS10IXVkKGSicFClwnfrQuYzFZpxtZ/hL4/16qF9hrZ4rjkJXs8
UaSoLgvjIQ5LGjs5/XqiV2EvkGavoW++8msVMjcwgZNQu89YtHrI0uOG3U3NF8Uw
PRpuJWO/GIsT0VodH0ktSDfUC9g5kWeYMb0SKxMiCtinvoLOtSazxEUPkDgk9W9+
MhVmzYzTXpN0YP8AQiT6gnppPb53vAt9E+g6q/XNIEIoMCYv2521KVjBpaPVZeI/
KFQR4lr4kcFk5Yw0p+cBZ3J3RODwpw2S/T/4b8wk2S6lc70CiwjijByVAZG5DBCK
+kO2UXnmUo1iWXmOaEO/8+n9Yo1vMQMXoJUz95Be4RDXC/dhSwl/7BrSu8UoHxDA
gtrRq5QpGBQq3QQTKW7sOolgEbV29x9dhEhs5UgtABzw2MaN52W0Rm36jiq0L87y
NFkb0xx1N59Ndz7l2eNmfbo0JPgsdlhB18GqtVfSdWC6lMfpqdnCUmE9hwjc2QLY
laTv55KjeiWTiMwsvf6R3u3JXh0Ds1ehsggQrxpGiE0R+5ReA9ihrqiOSDuQda84
8BhiJrwQRUslW75KjPJ4cYTMAoQMFtiso1Aa9hEjXwWrUKLGPk/StjhcWXnS8EYF
4H65cZGYw4Mjg+L7HaDdQtztVMVB/lRfsZSxmG7p9y1oM0Q3s2maY7pie+rdFnC6
NtAX5dDB/GLKqXMSep5ku14vIiuSGogvMAcROtHzhaLW+udScb9o+PQeJjBnKsbb
dsQpw6QdqunXAsEn/TlR6nYIa3HGEK2wyoes2QUPkh9Li3Sjb4adbsx6+WzLYe5c
nZZvHlvhgl/Q9r6hw3YiaXNWg+2wKV2vlcfdMCrjEYUbX4JzVb7QSyu7KSm7aE9Q
Dp4KDDyq4n/DsgKScHgKrE8LAzKCO2zsCDL3MJEQ+SRqNvRhTUaGP6BSRUl+ehvU
F4K10K9AXbm6ttiaD6vKl7hUyjEFz6mR3xw6HO99YK0ckD7/j5vdiRx9856Dm4CZ
+Moav1RvDmBVV4ff8zEABvDMFWioSS5bjWXceOxPgMeSjKPVoZcKe7Q3ztFG1uKb
5qwl5Lxs7QiNCIlFdaXTf2g7mqWQKfsM4zoy/u5eaBDmuIOSVLgsjplS/YqndWKq
uy15nFdNuJ+cnux90bp4l0SYotesRBdG8bhJZxhMNn5xKP+ea2rXQxkAW2axNPVV
Wl4WjRIDLUX9eVTK1N8toMT/AZ8USVZBhDWvyJdZKS1ayavnl80KTrtY7RQgeZVv
2kpMKfWxn814YjTCdUtHurLB5RwRICUNC9c6GU6SRpupXbpTdOus5ChyaiRkcS+7
jC1u9jjYFXJ28buY5/SthpfcwC2w3XebPr2inKbjDSwSWqOFRvJTbzOUBgSRAPlD
igFakByeFXj9DH7b8i1WYNajYI1MRpx00KjBuQY2/aFiGfv4zEaXpZMQXiw0D4S3
QO0rnscO0ID0NPCeMmrgdHd1WOxSja3OwLE3we/4JUQ28wj8DwpDd8hm8rP/mEJc
Qiy1lmthHLWq2X/IK/jB7cOIN6UP3vDOAi1XP0/J5UFGowTeRV0CNfNFvt+mlAO2
K3WK2AusUOweTnVgV+aNDZDG3g2ZhfgxtVvwKUF9zqd++gaXt0XGiTnXQrURHwft
IffSgjxOPptU6aIw3dc05Fl6q2UfbBtBufIgaWmY17QPQiG6OEODubNy/lUR2hGD
Mqn/hqgCnljRvJltWZDCz9GEqbjjEp5VXKagx9OJU+5bdd6rq6UD2/b+rSMU/Xdx
d2dTal4pXvCHaFQyFvZtQc4quyhb49bSNAFG6zBPJ/6bal5Vy0GbTkLXkdZIMJkR
NNfsCG0VurliiKYrKyz53r21oKXJXSSQOJSWeEsxQC6JE8cUAOfzCSkxBDhyP9Ze
+cClVkfgSosveLn+kkykd0MSQi9yc9ji65j/+GOfyaNoRb7mufBb8/FQ/3k7KKPZ
B4644VoPNiFf3QduBV1+/DXwgqwAxnT51GnWxBsRVliXgYk5YCtMicAP3skHZZTd
PQ9TVNZjNHrrb9Zn57b8X8KvYSEE9Qz+5/eim63DlUEuB9KF6sS4zIaIxmKSyJGP
ChLuhSCB2PzX9QupTZP3XJGn2eE8WwYIasnt08Lhg67cSdegZKCtEt0bj4rZhkC+
jcQL2XATHq370ftk4NE9ru47XdW/LbbYyyz07/6r5eBe76WCGO76pnu660Ds6R77
yqimoGr4NKbI9YiVik/AK97RGhE+LOTEfTc1E1MI6JTQmsuiWLPbaDwlpfQBDgM/
UYgMQHZcXlPURsnobUApBrEHi+Lw7FuEVTGeFQlgFHjDbmU9ALMlju6/+cq/ErYS
sOkzlzgieoP7Usz62TEttNkmMt6YDGgdoAlpENJoT5bvWcR8VOT6qoozfsMA+Gie
7a/vr+51DT1xopDJ2pu7FpbMGqLt+2WLJyn8yigV8PHVqx8O7tERg2/jr1XXNVnk
C3DJLd4lcKVH6HWKVkKm53AmdHgw8fajO73lkYHAJF77UhIxfaCndgw2/Nj/xJ0s
ELfciYDa9x5pXYFJ5PzvaqhQBHc3F9n3KD2zcglvNtiss9sBosK6EAAYVQX3mLxI
O/mEE0NANSI8XYcEZuHOGbLKakFinykTdgK02gJqf9qaZNG5x+d30jzjQ/AnGR9U
ECc3Ih7ErZZgFEvv9spnLaNMj5PSqM0gwswFsQSZ2Ctz9Ss1PF37NX9B7hax7hTi
9CTzJbvLXo8DaSbDP0/EtHVkJgGvp8lOe6O0RfjDTVMfdiNlhATa57F6sl3K7vPI
iAw71tDaHhZyTFmjnL3duQe+hQqud9bn3atOLBupK9lHLbYDKTzoQy3VBLmZSaMS
jTUUrYB/oBSB8ch/8XsnOmntBO4g5B1qdH2+Rxjj+LyMQUOrUWrVNvgHMF5BQ+o7
IWyHWhRFYApsBY7F+/cxNAmRRs0OnLT8JYcxqjQFOutMDxAu/myIimmD4AcMRuzd
0CEwMyxO8gyCPbcGCBuPQf6z4ZvrB/kKm4vHXqto1k6bGWlFcOdPLxhowuNJwnUD
kaDYPZJkaeCE98LIYGsQ7A5AWjv8hwKPTOB5QEv5+BNwW08MQTql1cWIBbBsHaYH
EqaNgzBQU804xW9Trs+VljHtXNwsFKvPH6/hJJPqzbA/FfSD3aafgjwbcuEPhOIf
hpz9ozdl4Y6Vk8hGnwXE0/cXNQyOPQ969OBe12JqvaW0ps7liWbLVRNoXLEgvf1b
y3NwBH3ADL2xACP7O7U7TSmCVaKdCfuVP6hvj+AKjBUNNRLzSUVdyUDnmpF1P9ta
0y1W6Pm+zj+toRUNv1S+ARcR3pUwIzX2nja7yZcljx3HMUL0nGriu+G/xhIDyjHJ
BqXvB2ySU9nlbIV2gcTciwf896Tma7vmpATlJ0MSnhHterWncf+1CrAr2EipUvRB
KiVEbboPFbGvvLp5BerW0zj1w5TUBNVIxDVsWfGsHloifQMwfJ6AGZ3sYIb4WFgH
WMmwbrb/J+CWYRtOCk9Pn52wXghVWkqBxOEDSY+X1tiiRHyeywCDRKY+W9R1SP1j
za+oYZRGU815LQB6/eMomnaHxERJCvJJV7YAAF6qr8PGzxgoSLSoKceyZZxpgagz
xzJ2rB1o7bUslvhT26Oo7IuQ3m8Qmvjw3TKHZjc6J/N2+tWA8aYcBGP6tcyGaAHR
J2IzgE1wwyHg2ZS/sYtQW0P7GxjVD4TxYKv3JR8vZTY2TnOk96ltYC5KukG54MI1
0ZRX2Uvj6U4RQ8Gj3HLGYWtgq66+s8cN+ROrjT9QMbWHIksnNrke2k5T8shbrx1B
ySGJemKavp6iOARUvipAMLH4Vy0MGHMxxc1rmfVT3zIJwAjrz9znqvu2DkrObAAu
Pi0Z5AiKV5I0E9qcx2yvxMeBeD+oeLXWTVVl3nAqLZ6jXzhxNiXN8RBRoM3YOvHy
g1win42tiL8rRhF4WeA/0UH1gMOCfQZBns8D9ZwfEV6QrHU87HXD7bL0N4XT7EuZ
zeb0WbXHqrM02ZIEbsozvehnO94MfqAAOWfaj2aFToAkl9XG767GjF4Ehn0yZgRr
RZzrHVRIjs9PwsGjvMKGov5TVkkZFAK0CJBKrEz5k5Uek+vTU8Gu5h17Cwaq/KtN
1gCmT+I5G0K9SVWdTete59zHle6vizgWwlc2ClWrA+Pb/hw6jdhJ6zMooxHjtguN
6Xn7hKw+ss1vyJiVlV8V6CBHz/zdXW2HwuDv6ux43zs6Nz3+69jAZDS07yZZPEZE
poC7CvLVg96I7fZpV+iv2tu0n4sMMdjsIOM0OXsh/hSfs7ScVemCOSPkbifNsyEW
av73qYaKkxzBj7o7g3PZ1pgLzPFp7o5/mwDwgkSZgS/NN2NcQVfoi7gxUaSfgobb
wVv5t3I1AG2w4QSf/cMWKq43GmbE/ugzclFdBMMtQrDocSLqgr1KM6B3LvUi/ntH
hQC/hwEaD1AWrem2Bu0o2q1XL8n5aHB54dVpMUAGCwCM5HZBnZkgWVIa/Q7pMg2O
7gRaYXnT/hE5qz/29efREKsoDzgwQI79WgvVB0a3ei3Hp6m6slOESa1HLMzm8nxa
BscqvWTiNe5D2dCDTwELQ2/m75rW51bwX0glfDdufXlXPGGBio133p8QqS/oYQzv
KZaFlHFWvLu1P4VvxSD9fxw0F9mr9KeTiqqqVBMI9Ctl0nG2SXpCtDRCVj9pRzHZ
2Gi5bgWEZZoKmFxkp59yq5atSZOX/35glawVxd8lqQcTdihVO9hqv9uf8au0Dv6H
8P6Jr/mUpmkmNnxsjL1Xee7HlXEfCkN0eGW+Q1H8arU6Fcb0+r9RVMcsPv5DJ5+M
gOxuQ3okN4RhRKPwnMftk4IROh8d0dTs/LAejtucw/g9wsRxfW7g/GQ7pomJzTPN
wWrKEOltutxbS57vF5Clig/HqGtxAZaGUDuEgof1xemu2LixzdvP2TrM21B0Pkas
Vbh/EUkK+CRbImQkWYx1kh+DywcojFi/zyMLy1TuVCif5Waf93mQ5RnypJYTSu3/
nQc5NkCpM/lNGKGe1FoitIq1Fq8ml0nMDNKNOiKhw9poQmreG2ndxnEJZVgn18zl
A/5mAqt90ZzyfSqy4NyVRDgGXap0xeJ4azHfjTAoi4wDwRMSV6r+QoMHPJYXxK+Z
QnmZ1KaC8LIcylDWv8523niqam+sTj3KBfBrLjJJoQ26PqR17Rm/t5NNCt/lP0xO
u5tNrtNBswkZot3hyNFZsuKd9mJA+t/U2loG9941yNupiWZ+6X6KAv++9oMVCOdd
S50jlzHIufQDO0OLoyq0+CVnC4K5a1zT/Zp8tHRrOztkTDCrbbMQXrkPYrGxXPXT
Cas0Dn8yZIPRhXOHNaLM/78uUwh8hFbOJ+lk32+Dwj87lSStW0N/0gzwjwqqOG02
K4iWnb+0v5vYn+pXL7dSdIHSp7CPIxdxQlYXkBmjfWPhMUXq6pLIq/x/asXmoKKX
5ieRCBeTCtjA4wLS7nmJ9xbMEGBq07kvApdtv93IxryXzkIXe322wkIrGiL8/TPP
053qC396AAywmsPefJ3FnO4XAC4tbSMEY4QX01yacVWCE8p2eTpIkb7vhd6kehRH
upmUn5AG3u9Wx+kCAdlLFkK2zaBQGmfHxiAA+hvsEMhtUEX5fA9vlsMWOfUrP65V
EB7DSmP1iYaZ+qBjZ26Qbufiwi4QdMxr1BbgOyaDhGYqF09nxsPgtNWntTQbgqPA
Zneq0KQwjuzNsloF+CfzlUV7hKmypfM+/QVcx8F7ck2YMJ96WGHVPs8CWLFjA1ZC
TN1S2Cg7jB8NdcMaggQ6JvYBP0TXvvmG2DBbAjOvJL3O0cwvwq04bEjXjaxdlX3s
dkexgyY6Mj6znGVv+nDYnOwOqKQ2eY1KksoKzaLS6drOARkRxT7GBJpq/GS9lUif
nqj2+erz4SN4OT3402gn8pbQ+/wyhcR5DajiN1Nhi5qMqdhnNq5AhA/MTvb6WhKk
JeupQnrnjM1eIgcvrwWYwiUEzojLFolTf+VnEjQdp8fiV+J/ZMDk/RvRDxrrteUi
YzjjDhaV6XjaqUx9AEDlCo9Xg6Q1EexUDUIabL6DNYgguteVeyMvC71ohg6I7+Ma
jGCzoPbZIiie24SuUfV/j02gl5VMmNXzejE3VxqDBCxS80Hk7Uh1evqoXLYAmlqX
0g+PSe3Z+jyYtmmaWxmf9XZHu0xpdLIpT0/ADVLOZQBi0nAwmLVZITuRCtvO9MoA
XTWMrMPqSrONW0AebNkobwwzp9E1/kLSzpTIaVH1KRuhYtvepM5yUJ0y0InSte46
oKYcqchdf6gL7PQWSPf8T0lsORzY3okRF0PtQoRb3EdaWRegOyLKBFdEMg2dhK87
2h7T7uGibOqFYrSAuIiFPri/G1QrsFcHlVdGJJOq2h2JqOQ9sO+OSgKck96w5t0H
H3kU8zMBe409srY+YRcjzuEYyC/1cE+43i2qvGQG3r5qCkKdDvJ61kZevBruJ4Su
tj6fHKCb+Zjxb3X7AkuXIMS9UN8l42ox1yuEW7LmNC7ISHfMdI61AOX087V+OZG0
efe86TY8bAbX1Lvc8Bam5JXeMW0Ml3gMYnlEiahFCfHn8q8ZT/MzF9QcyhAtLY+m
nrPCthkjw2/37GVHG6VzynNDwDQfXfvQRoEh49oxXQNGnoCzzcUDQCPM5fRqv/Tn
cux5nzs89Iz3ISTgAG9sxYH5oPfI3OL8MAgI6myqEHCXWrKEBKhuim6s7+SyLz2L
ODVOtIAn6LcE9ELyYhoa8PotnpAMyjC3AjTG78lKOyAsmuyzNxsmq2nF/45d0dtZ
O2Qe/NVwprDv01/UdKjC8t9ebkH+6+d8jRZJb9ynXo6qm4IIO2cJNdHjEQcA7gup
78jCUuk4n89vi02CfBcOSeKFbWtzm1FWsHTLyfBHiH5KVpTPdgqSGhS95DxTwnAE
hHG+3D12p8qtv1Jyc95SYMS+awu1zEUpwDQcm4lAMukwnp1g8fYreYfPuO79ihid
PWQqY61ftcBPefR2ZGNY6TgeGJhDLg5ZPpKaBzkJFrKqb5APqFeX4c5ZG6ZtgK7s
sYAMlrjc03W8Zg9f5FF7KCpIL7cw05kutjuP1glNVnHN/Q5VUq0WKKTyAuKXpxHU
C3vupyT5kFtQO3uEujCxQAJpMGNBBP2m9l1U+cw16n1lV3TX8xQB52V40T9yXHQl
Q5/Hbl6ufdUVJCG0rSW/wxU3s3LYHqDCxCC4IuYrMU8FeJazXXMD4GkCy+xl8v1J
mCEnsnqknX/zysZq8RMO5Ru9dJ0BjyBMOzJBhKeODnPJptIRM8uf44HvMXlKHMTY
Y2ZHqAmQJWawAANohiMgpT9Nj4ldTW8aFEH9b7T/+G1eKY+iIMpeo254uv1kl7Dj
W70UKgJoAm0b/d5RmeCd9fWhkyhvrq8mu+0Fvk4UbpdibKSICBM4cQINQhWgGJde
N0A09B8xFLBrOkBMfbyCStuN9r5GIEf0OEAWB7TLzTeDpEIi6Y4I1GfGhzlFkKt6
Is+JNVHzIU+5VfMOya4ohlvV04oHt0EETpF5r3a2aBdd/SBzZfCWpuwI35hv+aIM
34vkA/PSsg8IBWgzluF85H5WYG5Ahg+kChEHx65fnBXp1nGNIo9ZuQQn2FiDRf26
0JWKZivwZRMX+UTUHTHtuDhbhajrPYquSATPuc0S16UUgcfreWVuPG6vNqb6PLAM
mVdhQuz6lZSD9Vz5gg8xFny85R9SUpDhdZHL17fyaYgN+GGxN6iFY5010TRB+VXR
p/FW71ZAeJO3Cq/R8gnmRdYlzYrlHM+2OgzyzGauWhRUn4S5QEnWli5wB2P6tzJb
Z2QCa722hCWaR548nz54DsTV7lcn8S9ejc2RgnAQN8BImMr4HrCLdZ4E8MNJLCT9
jDv7+Tw3dzmtNd2ZInBOlMtHHk/TWNHA4ls91CR/qWAwiq4kcLmFWOqKVWICiDEA
60cteDA+zmwB7BfAOMQ+jjB4tYDu0fIex/ES2S9Rc+/8Hb+e2z3mEq1fTP4UhTJl
byWCg49xtOmj5Xm+n3GGioGct6vAy6eC29gRJFS8E70Rbj+2QbUt1scisSzdkgcK
NDWrb0L9r5V5Thm8xo5sNaRiegOXQmt+kFrcFbrzZ3s+fSxBKOD/6EuKn2ir664S
Gxt+XAN2dno91QyTT4w692Ks+KC2dpPEp9wxI8iexizuVwA6yodmlbEyO1WqWzRI
PFwaEpRgXl5p0SCVAk+NTYgMlOQpFKCQ8JYDGIX/ueRLKcISHSir610KCi9htyn2
ACSNLKi4y1dzAH37ZryOYi/8FLxbYte1HlkaF0CbWGaUGdQ0lKJYIbB8CXGWNdZ8
YXY60ZgC3BOpET5yqBDT5oGj+fVjpFMqtv/HC8Mq1F9UljbXk7M3VVHQ9+0iBiH1
x1d918hsHY72KdRi8AF9XKmzSNXejQnBCU6R8ekLzXOPpFOVVgDrIUF9uLtojrz+
vT292oVmR4erpDdXnpS+XKlO9vnbpATmOwP1dh67CnbLHkqfXP/Lth6ZjgBS0GGk
bI4Ds9vfENlix8LkwU2EUz/+LqR68pAerrkvLBpWkv1hk5mP6oK/2aL6a2L8l1RW
RLCK+EZI3q0sOqLwJPtyWFKewueOHLEl/tR50GmSFg6XUhGiVirRTh+mSmTOHk+d
2pRZWFkLAcuWzUx/l+qukJY/A5v26HXB0ibQjJuFXcsj2AMhYuj0cWZPKIRHYKA6
D3udW6WPlHXtBKW46jm/f37OKs49Matb7At4iD611sCprvpyMEgSUbs9sUgvZ2/4
h9FecLQ8wBfbZ/3GBrIrYPlDZjELxYKQKh9XgKf6F8PClm6PoFIENx13hhy5loRw
BMScO255A/t2F2rr4F2j0/N2bciZ3Od2GpJjPHRgM9SrQ5Yxwe23NxOCiYMKdOfe
FmLWLPHYuDe1KDC7mpM0BcycTTyu1QQr+TAgqsqe2e/1iHtybMiH1jh3O3m2lxCo
ZBayPYe9I5xJjGcfM79QT7L57H4jfn1MkBOAwo2NnQzhvGjijEHIj2SFmn6saG2g
Mv2ERA4GYcoDNwoMWSSPYEnISpEjU66DbTdAvvGtzVTCJWyXvTGOQfsaB+AklpGX
HiLePXrw8iilOD0GGLjS94HB03KfslaqPETSf/i5hErrwKHoN3+tfQFNHemvwHrp
+UoFwRsqgyb9oWBYoRxclqfRWLMbfS7Co66rb+2tsquEyy4zBwgQ++SHrcnueDgP
bc7qMSIJ/Sp+QIqdguw11bXbR1WcoBJd06C9PhLVBJXrJ+jx0XSbfVTB5hDjPORR
zUUlF644dOMTsEBnOTxkOCgJCx1XOeLisLZJSaRvW/AYiTkBPXxVVUXThRt5bWGP
EPAdHcdvFmr7/1ZbhaVhV3ZwZwLXqQ2NmXXyjg3AQY/PYBULD2j5HR4j0Azz6t+x
UNV/rpaquNKisgty+yQVkaURFcPRNM/e96NyKMyHa+O3flev/KxChud8f6kCCeEn
9irw1ZfQIMgrO9eUfKfIbPiFGvzDekx+AlXkW6EQ8oS3HDfbir4crakNloL8IlWc
L5DjcHjR0lea7151C6rtLpMNEC3TvmR9KyMbBP9oEDsWHd1reoN17cMHckFT2g9E
P6YqwLZ7UkPsnQH8DBL+tUFj4wgT6LUr8HWfvjzXpogq3BL1q+0imYwZOsfpfXlt
G/vGUXYRwUo6hk09NNLf0gx48g9KSPEvBYdTCGrENOI/DySSQKIVpbfzCjeHKLA5
EbZqVgw1rAJAXEr2NWtzhQEpkxREWMtxNVEIuJ7O/0WPFw1I6i3C+COB5URoAlG1
ja+QrtBt7Bj4WxEjyzeaE3uI4z3LPt3WOjloBUyQH3+QOZkA4UhFeNHtIrx6TjkH
OQsdqiO05sWBHvyvT0CcYYBlU0zOvdGrZmjxVJSjKP3HTlJmRjtzAqv8KMpMowEH
XQM29rIVoqPHeuCWqJbsya4hORQCYspNZXlmcFpLRkJnqDNmpBN/mGb18j4s20Ds
4UAR1w29zmd6g4mkT9XEDh7wj4gle0IbIC7HNoHtjqLhbdqV2I0h/Q4UgxhI67ck
chRQibg3S744fzcB2yVai594D+Ij+JQeGcGvxK+/IWCXfxMl2L9UaL/DiYkjCHGJ
0ElkZkJCPGWhY2YzbAYRDxYUT9FpRAAfG30DTE+yIzfKLPmlet1Yjl2nNrbkPMvp
ukhFT1tCxfi9JDvpR6EiukRprCj6CTA7kPzy2SakjZPcj/1WdI9uX+rrduvz+b3x
Ce6DBdk1cCQZGEx0QmDlWxVdyo2HzsllCuqFwzmE1k1VmR3pTrTU280nfGxTVJMe
ly99wLj//m6qZLP6sRS4RCbQfnpmixWsp6eE6+48jSbOuw1GWoo6J1QTRgowjH01
bCEY0pYMRZSuAPpdDJ6aSzJK7XKHeR2cFi0IRB0899PMtoGa4pK+R3Gp0rs9bLyl
SYPpaFy4/BnfARu3Ui68nKEnVW2OnoqncVp9faQWSS2xCUD7OrXAjnFcSxaYTqmW
hqj2cmhVUM8sxNMYA+gbfiw25aXcVQY987Zm4jx+fLGh4NaSztKH6M+AJmrSBxiB
bCHgy94Ee+4OxGGSqikSVT9QzvdC2IdX41IRw5h9e81JM6Gekjr/CfLsLExOfx8z
OtNKSZH+B83OdnFcAfJMtkmJ9RFKzSnjz94Sg9KFVBY3yAAl/ciZbc9/PXkFyNF1
IiP5ubiLa0mDIJdpx8S6Cb9WwuWsHKFPHnppGdTMffi7EijzZBHKxPKC+J5O0YKf
/Hipwtb9F1IwPb5Qf0cd74erMkwywzzt99EDZRX4aReYx4Yhww0Ar9H4OQd2cL4J
+f40q/FjtGpEoX0YKKFdjNAiv3s+nVDNoQCXfIk/bR3CnO8jc7TBxJycOiPWYwn+
wa9W4JaTeQi66OE731ckDPdGiPRdaQi8qi/tgUWhv5G3dYLazJfUB+42lfAeKiGi
ukyYa8iWADLAP4a66rZ6X1rtXZ1pLBJzrS1HQ6u86jc7vKNK0JawjrbIhLCD8G6I
fNYdF6LYPJI7ktTKUil1zCLQK5Hg8mSJ0uPQ+kKesB7XeP3kcdLqJprfHsF/h5yT
5DadeRafx39cfrpgi+AuQWwvMr/wr7CoBh7V+NlfmNHU+Hq+f1UnDFTsH71T1lxK
D1W0TqDsrnJ5XRmuijJO0Jlay7Opk3rI9pWX79kw5aYuB2H2tzTKwXcNOCOuTZJ4
tGt5K0HupsCdMuP5NuNHSjmfgAQ+LBwg4sMil01y/5v4Uw2JW2v0dvVeMvB6Nj0y
fzOYYU4dFhEWL+5QMVNSWgFUKh/ZzW0uMXxKc+9muiR3lK36GzxH+Q5Ud88Z1EKS
26kPgQJ/w3zzyQeA+Trataq8d6HsNhGmSJYjiMpsKNNK+QW2uSAZFC5Xk2AqAvRi
W4OAQyi35UfeCbnm4xDQSvdYpcS+jRPnooxGr1Quy4eih/PRrYfellZPU9QjOrfr
nfAZwKJIzPa4M0Qjc04ILrIBOM8FYoItW1w+EjCYSPgLqUqoLxC640dxA+ph1m9R
0iQ5WYzv6sI2wj/xxKnk5wt3Q0qxA9JajMl7hz8PdKd1LlzhtZCH84ou29BJEL/i
FNokmmDx9mmTuy6UzzXTPa2/6Nuz9QzA6v6v6Kikvm77AUXqlhRmD0xu1KyWg14i
x+SAx77WRPvriBnWdR4YjsFC6CjZV55lSG3jbYASmbXb5AmJbNpsni9PSkWC4GhU
QVzpTQrf32ZJXSM5MaAkw72mAoMJF40uZg9+V+/Q7+Q3d/B2Sl/iYgnCEskS3QOQ
CDGXMEkR1UfrdTYiY+QixHapbH0TdNuGcOuuvYsKIee6BJjfxPgC67bjw9Nx1hW0
Vy3ITDoZs7G9t38XeE8imiQrlUdq6Rf/6KvwyYinKaSbiV3S2GKzdIGEscWsX+IF
i2gSGvO21o2dZE20t4Wj2bsImTOt3KT+yczuWvqanx38PQna/GHvbyRc8tbbVlOd
k3CulnjHA1j0bdJ9FqLSrtw//apimwlaYXEvzWpvvyvsVqnaopr7SQNgEQooh/IP
kZDh+Yx4dcZEbn9M01ZUcSf2jweDUl/UGatXL82Gop8oHF+FUF5Dp9POabHqEdX9
+BuDeSP871irKWYa24mxP6hc4CUOL/dseR3AfGGle6egSjKSyocr1FM0ccZTRSi2
mAId0cfNv1DIFIPoanA2LWtBengFAZklOCbF+dae0NlPB3nGheGOp9w20ux9n3vD
72QeuurqVC3riplXFF8sg5rDE/1HZRkmXYDtxLjeP3pT3PZs8BIqnMI7KX6lvxEe
BOsVbUIh4mCWzrr4g41HxemaOQrjdpHjTJvsChRVGJTIwXmnXG08x+/7rgEXAfVM
2Fc1Rwv4xHjAD1kI8IcOAN9GQHsEwuvTTqIX3k20gVPanoIqU4aTI4gTQxwmrm+p
HGvVvrYjLkwagTH4YkDXjEEw/aIGyJotfHrK6Rj9CM+gXB2jvEbfI++qyGQgzaX2
G+aE74ZBtjqsqJH/zNnzxidkpesa/ohHhQSpKrnU79feqbDJ1twiAWrDaH/NeiEn
nElilxtsl29njm6eByvOgPihtJzyvwmqZX93giKWN7BRW4bnnFj6xGxMnWu/ORWF
P6/fUaYOMSV1kIWcoGRx4rtQoOa9FyVPUzhU+efAckoUV+4acLH9AAgI2eAiyPWo
tdJkJIN4aoQLna0E9KU5e22V3JiyM6OhEPxAzP/Ou7ltc4TeOrk86ztGpIQWb1T+
uAcaYzPMBiKM4R6CFtIPaKI0E6XmSCbDot98KANOUeBKVzbRqFnGPGoRtTJO9CJA
ICOc2f8O14hw2dpSmUQSGAcdPDz2zrgQdkLIvK+r94kwvvrncyIrWXA+HKU6NYQ/
UDCZ+1lQnRj2TZ+veglJmRZZQ0vuCSfuCfJRa9L6mZ1oHowokpmrv3u8erm+//mx
IIxjnuRRqK9wzjRWrOk2wAyva+SKvZUTY0T1zBZEKs/8ghUb5GfvF9aT4RGUg/Ni
I8kCksSdeYbu8G2VB3HvhesZhNdOv7nDokYPSt6qU+MIGfrL0x/tLPasurQxZFko
4/0dihGNCdk2h3e9WNuBlQRquYA8x+pJgU5CZGesTxK2i+SAQm7BeKZbln9NIQse
cokNnA6Q9NOxHrXDn0DI6XuNdoznkBocBtyudNZCNPFSm4XUvl57wmezJTkETISt
zeS874tiakpWohy1bBDCxzgwpWoRoVeGqn35RtS23zUulBIx7xm4IByh6EMAM1lO
OtrBZgzL+763k3Qj9RRgLVq4c6C2cENmnW6+WY34dhNWEOhTjxB1c5ooTxDg+m+4
VxrloRZ/GEOsntVOoS2bVD1ogUGTorRTIYhA6PWxRxDgbsg9OfvJP9HaPbGV3yhL
NEtXHTyWvl7ozfwLH+rkJGwcvqA6CXAJ4i+yeeC+1og8M97rzWVs1PMh7j88/PKc
BajiwSbpPAeaMxVvzsLdpKiXT7GPyF95PMJMuwh3bE+o6P4jQfu/OKv3hTg6+Fhc
fB8KDKlVi6mevetUTzjTz59mUNJzm5MaJjpMp24WWNXE2dW1Fzx/zRk/+EvOB30v
0qCi7oJqqNWm4E0v4m5eSAoyTFGnbJU079Udzmxei9LRwPIaPNHCeOY+RpseWz7Y
qwGL5LCR07JOtjsBa6XZuoQxarGL6FNdkUz0KbnemUImVgggJfYg65rVY8MMJFpX
xsXrE3iWodeNoDAlwmPB5pG+7YGSzNRMZJ7HHqidwuOdGLcSAZFdYZ13bzM3u1HI
+R8bCRoBrfiZ2jYzAiBshYwQiKfshziOvEZZjftj2UIAbfs1Za3IzmrCVlTiJL89
HYk3vsDnRXcyVl2iMJ+Xpg8SawtnqK4uRIpby3guSB6fCIli80b4KojQ500HxrbC
Kk/4UajQIPGWleyIXo9q3ksq6HJTAZfyGagI/nAy9peD7/5iiXxsf+2XC80DS90d
FlzGFWCZugV6cZwgsJwMfsKPVbBQNc1rYC07amMEdHl9sQRiqbsUCyyZbtxMW4Hv
XFbyprC4UnJDm0bfNzzIH814eVGOuSBeCE8iYbKVtGifZrpXfQUICbaIMwMEfVXa
dMAfSQg5epozTX+yi7o370jl4y+UlNP0barHMQ1Ig0CIze2NcRxFPRJTXDHhb5vt
gOPhoWupp2z+Q8ftVy+wK1HZ9tzKqMdYhvu0U/zDS2dleFOk/ooNvByd+F3xWUa+
66WnxkafScv3DZhXbdrDiooRTfGcwC1QKJxcN4ZTktGtpgoj2K+j6y9KWjJ6cFqC
nrDb+P4QoHJ5kx1ohMI1uSKwrlBGExJYEqI24AcGYGatRs+tWTPeQ7lajIUoWVg3
rT4UVeN6OKkF78OmDiqdJAjxySkb/SABlP3VhNLHX9qscnuQY39hvd3YIW4QUTPe
DwG/qAfDUXUd55h/IQfGY2j1uD3W9JhkU0BpPYOpD6Da7uJw0XinjHHeK26VADwB
N6+O1cIHsusFq2No9fA8y0s4gksqDFp6RnNmHtopjE1w0a/eRSdS2PYnqXvWxWsq
cvdnkDFhEwKUcO01RizaEbrJ2tkmPoJdB17+mimdtqG3c59eBlU862wGdNX41wki
c5whd2gm3H05In2JALyvCN/Hxwv5cIT92iwJsfsIcrZaz8SHXngbxaTetDcOBaVK
Z9IJ9aPJKrmIS6YY8LqTjZ1T4sYOtzd12KW+GMWytSD2/tbccC1wOe5xmryACaGz
y0iltcfxwoDTMU3VcBOu5UDEqKY+pWbA3s4s4QDK4nRMCutcJXOZdJEXYCrLEiYg
wXjtXRebDhbC8pNokpHHuuaxOxFBRYMOsk/FFFj0P/oRiChH3LIki5c1YK/jkRAC
ATyUHOjUlwBA2RwfM/fYnxyL0Db+MYvKoxiekAYM1f7MCm7+FcfDmdkHy+6KF8jP
LGpgU/dozHtl2QWg+lzqPI46Uk1WbH9e82HoEocN5JWwjm015nYc8RYRjg/EdKiQ
wEDIZf4YSn9W19yYGY7qSR3NopLe0r/yynQnB0OvHP3/Peb/sGuhyFrqfFZc30Wj
lpl9wkTcjt6Ed9Myo24xtgxz7SQK9qiThJGkVr8l+cXOzAiazgmshYRxbbTkPH2Q
Q/HEXD5YtBfoaWNwKs66LdaAZkTLS+Hp2aRDo6DVQYJWno4H9t3e38TFYnntX+9S
lMTkQhNSg4kYYAleqUkWnlmDf73MFHaRjTTP9+caQMNftUbU7K382WnE6+e+XGhK
VyN/1nBGsmn3MoGZiIiTjRwJ0SHOZkOZrRAHFV9ybCSR16l+3smr0rNh7HghXtIm
rXl5CFQm0ChqOK8gzBcz82JSSS1OIPXkAKlGmiotIdHXel6/hGn4w051kaDKG/gJ
hy6TR9haWTu7t7udRPkHhJujZe6xe1x2ZBuvnvBLBPc05trE5Q0oOULXURm6eWQD
rzHyKczzRHWjwCpOxCjoZCWkBCOPIO2AWGJXD1UZ13cN0toN+QslGwwhSqspUM/b
XjMVn8vsrEp7mwcwmvWNzR6s2u2Qvtc8W7SsnSakUH3rypaz+hSbBSwvmn24Vz0I
JmXYLP6LTPB/ZqXEEHs9P+6atkdaZVybeWZp6369kJvhGAEM48yrlsoA7Glae2/I
nF1J1nCVL8yfci8mYpuGqm9xhV/qidHEtBL2VbioDvL4dkzdQOfYk7e2+2NDZwLn
u9WdPpyFgIOIzUYpvSMIFMDMFR/bnu3bUQlHckbvc0uD56Me3Blgas2qIDLQuiat
dij6IuYRAHbuelE5Yh4ZEfuC0m1mmH/YJWztGH4I+ACtqZ6QcT896dRV8QDkXbnh
CfEloOlKojvUHYxsIeUCANwk0dK8O1i453MHNoHnB+QEx73QUAIyhJMRA3/b/2RR
5tFJaXUow/l/U8wmBycUPl2FU8gkBxym9O0JQdiDYiMQJsVEKZ1cy0s9aGmGxDN7
wYdWSwNvJDtYLSGk1VsKWDZ8nMqOj9OSbIvFN0Ke2u1ymtxwFN1Nwx7SoTWZ3NzN
1f3+LepXT7EN/aVISWDn1p0WWIFj0DqUEU0A5EOV1Q9BeMdpoD5C4Z9ltzjN2hBW
+LzyASvzY+1Q+43b7/Emupcq+F7pONLBi9ReXUbio8Q0AsnxVp4XBG7Unp7ZWomd
f+x2K25JkhxN6NeyXq3bpv2Ni2teW1lM3bIiUxiAWPkcCMOVVuw6OFqbEH8inlGB
xeq0M6c4qPq521n6SC41xC0OXsJ0hzDavMpVtwwtgB4VPSotJFKb/zeiPagVC6kV
PtlQezteOVGZcXOBNqaTMlCXA7+uRQol3lI7HNw2gTTs5ECHuaN2zC2jykWcDTle
0GdPvzbUBZKCFhmRgL9SGn6Vd4dFgkrVdHX3/xodBBFn8twNh6gOXOTdiBDEcZvm
AvR6CWu2eICtuucBW0A9UN+4Tnhryq+lb67uPQ2juBKiJbdMiYRa6kwZkB2zZBxf
9k26uOI0IbVIcdNfdpp03AWi11LxqdMak6kL2op8GDdQg+XNyuSqg6hS7V619k8Z
2M0rR3lMOvzEEcXa78uGlWK3dp+ul4YEJt62aPGzoQBRiwH/MVbfOf8EOSzDdZMy
m6krryKQec1NPUIgSw6ymmKkwE0LytKt+GyWEqnM3M1UTLBJBQHaCpcdH4odqtpa
MBNG/ZEF21lVm6QE7YE6IN25om7dNTqok1PpjwTKdz4034/YloNXlEvFCW0PUutQ
lOcLWajHJX947pRN9Z5SoY0/7Uj8SJY70E+kW9rA/MogNTNjus0uIVmp9Mm2udTn
rCO2hL8C1rvgvrnOPjx8YtbDnyE7nzqKtjyvrD1zKeGj+Jl+YYnMYH3xdsk6p2lF
7F875+AovkhuC+rAaLeelbwHIYFmDqmuXNCKRYLfloiQD7VGiqFMilBbi6/vcczO
ETx5GCcqbFerYRs7m6dY7OM8hzk6hKFV1taT7Gp4O8mC9Lv4hNb1YLejmQvBVYDN
wOD42QyNMFzAOB4zIB/dU0rmXWTVzV0DiMfiQEyjvtkSSj5UyHm6vPSNiJ+hElFq
rpKp+1olxXYbiiii6SNhHcufu/4XzcL2zCa28z+GIvjHqKNGA+QisHNP7Rdvez6I
6yTAPFibK7YXVhBrNMsy+jjY3FiPWKaWpbFO4BKnHVQFGQtOY28+gTEo76TIGw8o
MJPqN0uMwQPRtNKDyM2E4htpJ2flJuH1eBPLycq78AOwW5ibiNcOLz/kO+nZNwKW
62sbgMF3nzPj9ylZ8bE9++jotn/L3qIMw2Jad5ZCPUs0o6M3klQuGz6O+66unjtK
IHnkBfBFz4r5F6PAX97hGXGJcJQ4kI1DX0+3ccgSaKnvNa1WtLGUuJwQbPAyKLyZ
I+0oAl4GNfXwe/EOFP9RBqpbj/ez94lWBFyY6oQhxcB2XaNDfpJYU28PulUU/e+6
NgP7nmlxKTkwSU6Su3CU4QkTlVJm4qtcfiYcK3Zzh8MBd2XiTMXnzG5AWQiDp0nD
WVkQVq5NO8aVZHVfBAC9OJL4H6BUxPeoYwF5mfFJdy/y/vNE8ACSfOUhD3zOX3Or
i5ApwtWmp9s4rzsnPnNYbCpRx/N/u00j/EvtAk5ZIMdNybTDty+2ToD2dQ3MIlR3
AGOx1tWVB7K8ORVJENXS8Tjih6JkbGW3X16Cz1NK9JlNLr8g5L97yrY+7w8ZfMMp
kh0A698L43WGASzSDFlf5Ac/IyBDgib4+qtBawisHbB1qLJRVyuavVwDcXGjB5vs
9bU3LnvFghII7accNxr52t1/yN34VZEWe2smWVOepcyzyFAXb3P6ryMCYDVPWjMG
qNlrgHkkhCiHXNIiu6jrSnQjtq5Y6Q9fH4jIv/6Uj9zFckXMX7cuG2z8u6hW8mRv
8W7kiXU5eStYCUPuPzkz61YecpKXC4wBzYwchAcgP3nliZILXn57gVmB/DCZZ6pM
D5OnfkFSCsCxsTsEcqyYLmNYLGbAaPwzyg5s1ELX6gxEr1sqWyd0isqjaH6686I5
Fqahet8sHSvtg/afLNuhigGOTGvWlf8CFRKghMtGks463+z4D4DYVKPOxMKiYocO
S0VIhkG6H7KZABdPTpm+DlGnPBhGrBH/nIPF+9DwL8zRgqbQuEbKzucQhYBLM8aC
Ytq37ned7kdykr9VC5wlOCgat0hmwGGLkMcxJd6yeslPazS12jtHDQZkEJfjqRrv
suuMUrKi7NNQWt8f2VA1Q8TXcyuNSspFxH0yihpqixfz5jXWsJZipmZeldcoqvgz
5iiVOgn86x8t3FuHzMMxE9d9PVFlNsc1wviPYw+2r6uMEmJEN04kFnWH8BgVVPq2
Ec54jfxYItnYf5cgLAJCyj52p4FrwL8N6Xe360ond0eDO6wk3634L2n+BbPsey36
az4kTeeMCd96GQF4KGGTnwjb/t8BhesToPrFQSOiIIQ0L6qlpgZAGKhu7FfaSmpM
amL8ZvSXgIsj8INFbhl7+VtbKfuijI/Ovx0Go5W7MrP2xOSmqTc4YdlKBEFBczM1
w49M6Guly0lXQ/3X8mK4M7UqX1mvX8zu1+eWgFdcrxmWISbiOAvqk8ddxSluwJIl
t+lFU0h2CxuzbCFHLFX5cFrFEeI5e4J8dSQq749A7Xs6cul7ShVZMqNsbHu0wCQO
rmDJvlRJB/qsRZseFR/f8lXVmdNS9E/FhBdL4WG4sEMsdyLiDGsOd5lb/pLHSACQ
6UFmEXqyBGjEf3kLdSllNL1OFvqRjeDeudsF/J2i1aPoYvhbK4twUz29mnt0anr4
wDyKLzjH6aoD5Lj6jA3PzIJMJBaGWLEhcJgmopfb1pCDVDH1whqQNY2LqVlqHk92
COHVBCBUc8rSjk8wNaNmz/VpFcPvJjZ8odtmxaoaAxq+Jtb0NUeV8AePXcpnZ2SK
aCCUCamalq7tZJDK9TLvodOW2cVQxa4l5RJcx5QToP7YCIQzMST9D95jM+gQqLJ9
7b+o2l2a1eQ5/7Lzacysp72xDNndFpmS2XCl8D8+hZXxuTkD3QyIvvF+HBk4F2gB
aoYgy0BIc0Zy0p2KZewrUd9gv8rRYG0KaZPQTLqI0uhiOg+YgqdzIQrbiFwEXrON
WMDC/FtaiCsxE6+wPZwlPbAZK23S/BgJMHEMCwnjP0arKzL1AhAfkfh8kowoRWdA
t182IIXxtNmcO928wrDIaMgApptmB0nDNj1q07O3xJTXDAhTDzfxEjb5sPvWqQfo
Q/6qbfa0Pk1AY/oDMdyIuoEivD4wRZdV7+VIL57OCUAQaVhciBOC+8IRUB9c5nwO
rZw1JkIwjnlcMv7F1OFo9ngePF5arGKwH6y88d6qOtfJTLT2yIQXmi+CIOyZuNcK
K+PGiYsm6Z6qipLxTN4t5XQ3DiD/9Fw0LWrnrQcM+StlCltWwIsfLwz5kXWwJIBI
W55Uc0WNq+SI+mcunVqIzXXMuMYQcxvKMhDt5ohrsBRWrCdRYDWNxt2A8u+Yv8KH
HpUFqykbWl5tkz2RT/d/nzNqDG7YyVmYJgM+6BpA7qkQcb75jBeWxOpCk2GKGrq0
S3Xp+GTM9Y6PfMgjW6C3+KJ7lHG6pg13MQUQKP5eCHexzDqmBetAlRc88Ji4Avs7
LaxB2FYFT898+3Z33XfMutAKa7mfDGRcHkG7r9bAQOsTVGs3cJYR6siNgvwkRd7m
7KWWnAXCy7JBlI3hGXJw96Sl9gxrbU+gQULTbyxYHDihtjdnT8isRsEOHjrqCufi
J+SyDBd2FmmnUJyp7l9AtbeLcWH//K15ezcZUcOgbau/N8H4nvmq4NFoSrnlmdaq
yc/aJECpQDugqJjXufg+CixOy8/DfZZVNR/rXY4021mBEg54nLupbVCi9gLiCqTk
nZ7EYHrHrPaANi8xgMUICDatAFxcZweu5CXQeTft70GAvmQs4frZf74LBUWcdtoR
qPn/0BQoAR7MKQoWhb+Rl8GKL4JHNfVyr1ZGSJqj8fvjlrlZGJSEGUyGMGHvCXTl
1b20rnsZAPBwdDUAPI9PfKRTKe8CPUlZMtcNU0npdEbG0cW5ljBNGbyYW8zUksTD
MFymRiksoKdHAtHTpnJ9pjKU9D60NRGdcWmEcgGDOLWvXq7jWw+wcSZhsM93Do5T
Bz9VTr2IIDXMfNLXrwdw9zTnenVZiBZIiEtLX4o8FE7BCCNDxFn2h/YkJJ71B5Cr
gP0UseJZaf/KxnAfolOZQj3IboMLM/0SNj6wHOmb8VrvyVu0tyR7VNVABBInLjzd
CW6Xo6569Sws6XaDHjG3v5DDdIN1asQJkM9q7CZVwGeaUQLpHVfheRBAKZ/stu9g
lzAN3XG4dB3A2R17/SiqzfDWtgWo43rcAIxxHEgesDJfgutphYJA/BjEAyRMRL1M
Vbq6JbUAYIOP3/sIoir46TEi3AK3Wd88GjLSbu8cw3Lp8w+bUgtcd4DJOvIHDRB5
IWiW5NpktrmfliSgTEi4n8CD4wV4wFl47lzV9ROTJMv63osfRHa1PvveUN3okXn4
sGWXNGSUk6qZFnrBWEfcCX9fvXj6ykWFUj2sbYO1QOjGSsAt9ckHCoCP4joflef8
2uHj/aa3ZbWKLFrN+oLHl6BroMGdzZhjViQphHrc31BSgyT4zJ9GlPNE93obLbG5
7oUnpQSK4iuk8g0OFFcfgZ7J/0YlxcKcWT24YaSmzI5U8UjOmwJImaRA7VvacwU5
WELSY3fWd7Fv4QpnufoKLJdh1Q73MMs/VgSc4jBPe4YHi8ECkV8gnMnl1fhb3WMK
I6xsgGL+hKoDmSOmiKdWIy4V3nPZfRAsIGmHt0T8u2mlwXMBJIB0d2BGhcvgXsY1
eyZo7itHLMygmmIRcC8Af1WTnnUJSFIo1mL/DdBRPeBZhYYCzd/sZHo/HvxeS4To
y87olHTRirrcbRL9JoJV+MTd1xN+0XJDzrY8Ky5hjAyL2KyskQ+zfJCAQzPayPR3
lKOdS1tgxzq9NE0gemsybShUuY2lQtAHO5+K2CnDR38S0EBYcUZ9qy9K0DSStm5z
gRxChgBQqaylXRRxFP9pcNYVCfc8e6z2N0y25cWurmN9x1144Vv3NUib5k88vQ4Q
2uZqNMVcxlUJ+FQmkghIv4aFPsEx6Hpor4Q8s0hbCIWAxcJrLw4p7vFpFLm8lMo1
0R1x+Bk1+l0e8m6cg5mZAQ/PnQCwgakyVFmNyhYnsRXF/ndzwf2/zJKlmizQn5Mw
tSU0dwygOZajcCg10xF/c2Ajf4QE/8pHqq0wx4qfmT/sRlWB0TAh2E2a6P1GwjRk
ZqMo68ZqRI3pJisGQIlpHYXR45LC3zYYabhA8hNre0KJuTdBByeerYpIh6Qmu3Tz
uhc/TGOIPmsnAushYB+c8c+c5TqVTL0hcLz+7IOWQqVqTCoa0cJIa/E7BtmkfcG2
SNAcbPuBrG+BWleqdm9G81v//cHbgEidtT6WCPFNmDi+y/ZLRFvFACp/dfNwyQjq
5feJ9RTQWEjxv2vT/gz0TaXTXaREaAg4qDGundFo7eNauZ1G0ArZwGT2e4MHL4ED
W46CiYcy/7lTHjOJriKtXpDfvZ0tKIY7o/CokxGnJ7C8xeLyLDLli5a97cygva3j
tshPjnxOSbZyCwxKCjE257Vs0SGO+5g4ozsbxRQ+U29rSzCtOrsFL24Jm14qYC/E
lBWxbcPSF+FrsoZWMSaHTlXtBS61ivrPwKgwWFF7rT74OP3iJS3b/3KrJQHtawZW
JsT6jKFDw90bU5JvOVqOnhsFSyjvGFVBtEvnuYX6uN4QF7uhlzkC89vQ70VuQPW5
xkf62lTHyyYOqHStaVenXEubP/R0zIForKU4JP5aMh77JVfx1Cx1g4SMOfan46tp
OMfwNOs8N90XnXrWelQsqtbJkRgS29L9iC/j7s9hOLFYwdhGlqZaFux+cwiUPHyg
VK2YDUfz7pLJMS5txDPmK6uII3/hzt9djdMVspYW3EjGXozByjsPTXd8LZAldszb
t/ZVKO8bkfG8UALdykbeLjbXSEN2tcnepn/xP09ZpHecwMYJlT+WraRi7Dlrl8Cn
L19R5peWIuaOF0Jz0fULPLFk33cuFCoHUkXL2iwrtW4FA4eJr919v9Zf4w5ZQqow
PSxxW4dQrfvrVDpE4NWayt+EDL+LpNnACL/JlPTdEl4qxac4iYvr70d+4QAron3u
KgNeqMBragpYng8YRpTmBIYgc5GpT6ouhdNT3ZLXSpvffBpHPiUuMWK6N/i6mYCf
3tV+z8rfC3Qf5GFbzjGygWWJvPcdFhfyky1Hu9fcaE9BCtllawgkZd6T1tXpYqxz
xG9PtP5+zS5u3rOgGeyK/MEOrN2pMWGW4mIvAI02E967P/r5MDNBdbUToNcEX824
gzw9f+pYfL9aLfHj7C3e8s8l/ZQx6w60nIglLqGrFnzr5lRlmDG79wA8EgB0SMaC
Yw7SpPkBiLduVzUC/waIRtpqGWHwKNFzxqs+vkR02d6RFsiaV9zt7t8UOu//nqFB
OZcv85D49v2P0NdWOhcy9lepk2N8Cyk9ewJzkahPFxa3LmkX6CYuZtjehwwpgqke
0/FQ5PzqQa5N0TNn2+uBXwAl0971JblV6iPLcbSQ1FMOYJ9Zsnm9BA8kCCawINCx
ImA/qfpZdiBqxbyzH5BX9VB2/t19kdUAf2qM3xS6IK0UmTt51JqJorLvTlXejt35
67x32OIoJs8Lk+PcI4gdmXNEOccKAKhgocarVIZi9NdOLnLqolhwkOwUreMzrLdR
E7p2x2Tu0AnmD4d9TRS51r0Mb+tsGlaKkrg16OmOmKZWrCVWf5W75J7pFuyEALPi
qxHeOWGb/Hd3dMqg8ABD8QrSihgO3VJhLr+kTmm5BBidiej7g1jEZmpV+40EG72g
1XM2VfDnfJRJdcWI2HCbvT9hAESyBTMB9UcW4ILJQJmPueEr7Fpay/SmDgXE4mms
PZ24npcvJrl+fQMH7pJnqkUzJDXJPYN4hMaCf7IhrgqORWVhf0czjlt22zS6Vjmb
1gznnB8eZ3Xe5jNg/8/V9gv5aGg7lbkXQBDhx/oV8qFljJJThbli649MlmsQ7iUJ
Z2CDKljLTLq1uyPyB9JLEBrXugCFKJ768WUWwwm0V8VUtKXfHx71o+P6y47k4yxm
MPPpB6PQuLJFJcEYmMLriicW48nLMfpDiL9nNIdV2iF6qgVKNB5qK6xPy3iDHnNQ
mULTYTqM1CwZctIOT8AEhDu0xXYr6f2en2HOTOYVIS5EhHuPVv/8d9sH62QKVQNM
6LV+W8TP3ugOtagSGIGVUybkv7UJ5v+No3GNqS1ESwms0sFJYs5o5gv2hKmmI8MN
jWTs+5f8HnjUeKln1Q+ZpO3sr2yXGO2XK8Ke2sxjP/MD3g/g04TCVPV3UwZ0ggC3
Yphl52r7vgqs0DxuonhR6T6/FeZnWPLbCoUx8KiGSA9KXf+UvRxwZoKM3Gb9IJuH
gxOU4oU5bJR+e/FANTEN/HJob1KfHVJ/5PzzJEegIfuMdwq02EJjsCky3UojL8uK
h+jr6C3LNtyXAk4nvGwSpUkuM6AdnRLJSlwhRCaS+e7TTguyb1zYrKuFDyvdS+W2
tTzaYUYxRi0rLPbogQrz4rSCCiSNNSYK3K7YZ7awYe+pDZCwRqJYmNHwHqqGY5Us
Gta00AdxKKg6OvrruUnOcldEF2PhOvsN0a3UT6EZX8aHiY+JWq09d7XU9WgWwmGh
mxo3i+fzAmjDcIEdyiomGfqD9nWcc8r2e7O88dVxQJmRVHTEWOOPfnqMfvx7K8LN
kYIEQCFRve9wqxEIEKK+vXysTm6wSW1BU0b8lZliXjrs7skBDsWyVuB/BmaazCvR
vC9KWWDOVl9aleqeKYr1yoeET2afzYTehBOAJDLxDwgG62kA21olkMkimqIcZhS5
nwwbTCpmYFKdif7aDiBDLyGECtxlAjgcxYLVPLPUc9HfXhLf4J5FAsiCO3UtMQUB
k/z0uSzVbLyWvBTAonWGK9laytmECXCfa8X5r+gKjmOISF7sAidf2Uf3bf7+vREy
Qu3dg2R6PcFjrsr1qX5G+sKteDDgT/OAmtwz2/PEeGAT+YDOR+4KrLtL9nSwfTwO
zlt9Z2tQSgQfA/bbs34Y3UyW/DlkfO0+3Gp8LM7r88J9SsdlbyZGRISYcc609zYI
4hqoaZYTnrIZRnna+PijjY1LgEkj9XytDrlEX64p7y+f2xlwM9zcvNhbOkfc+kdq
6yZA3aiVg7+Dh/d8ee6vkJXqwY4gpHeEfw9AwcnBUcHJIDlOLjeYVWXNl9AArJue
Ot/F3jB9QFEA53mJRRfosBYRPYapYOL4Dg7t1uJQrznc8lotivGlVfuTy/KgRYft
xErhIsBxfVxUkF+RdkBTwN0UcsypzttsACeQxVXgUdS0chg2YKjwlb5kmsIHLy9J
NoC/bKkR7Xjr3ZfVH92qlSX/hbL6yJCWotUwbF4gR2F1QIftvmjZA49LV2CtlR54
qvlHlF207grmidqaVF+6lV0JW+QZbxuw1rnhy8nGCmgbTJD3LaYbY3q13m/uPXDM
nIqrMGzzXSC6wzuifO4Ay7Pd1QXPbIezw9AjLXbA9Y1uqzoqkYxZfOrcxV/DyE3I
SKnxIsW0VJ2Tb0wsjNhsF/uN5Rf2riyIjMw3FaQwdqQ04gZNsvBf519ympzwRURi
C7ihXiiuhpcHxNj9TsFaUkbSJ4R4JgcGsumuyRMWncwD4zZ1NFC3yZOdbJiRFdec
YV96eXhjQfD4+Om1PotDjSfjXsfqUv9NCLcJeAQmgvULuzZx9ecJtI6KEE6MfPQZ
u12oZITWqwaiM3cjvx1J6x+HpgV4P+5hAMVEEO1Hq5Qr06g5bSdxvWIF8reK0SXi
ICo3xn7eN0KDyEFsPolm2JO67I91VX1mdxiz1iAvMQ2nUoWXhCC8iqJdSG8AKrt0
capxVPiyP9UL4vHdbQyOltHIDMxzqaLu3V6lpb0gYi5jYVwysb5UksYocn00uwU+
aAZfMTKFni0ua6TjVj/0Mj+BBTQZzpX4OOCT5I4EvXkg7Q64i0qr8X5kSRLqg6l0
ce9uLDUoIHhOYd0psmKwsuslszAm+UF0nKrCtPbR/hP12MLjGu0RAWg5FUhd6jlh
6HieLQvucppRyV/K4+Desx02qOHCpQGleq/o/66ELv6DOpFaxKYN2r8Qy6l+yUpj
3UPgVJmt6YKMV1kD1IppKdKWmvIN42OAInqx0c+phrBe6RFMK1zjaYoYmqOWFVdg
rTvAQs60YTa1unwTaplihmgBU8y8sSO8YtbXLix2nKqRyAXoHdHUY/i5L6KSDgiW
B+htm1RYDd254bwHsOrs786dx+6yVFLSn8lN89OXEcsvVDcJPGUzqWGEqGCstEdJ
U955Oa9JP/ecIzjaBXCjQA0mp7Gp1uXbe9RzkWB3QRxu/5f7u7KgCUM26CCxvD/P
sw3wS8rWqwh7y6dGpEHFP3j6cRcgj0q0u86hSmPk01JV15dUewh9tm+J5rfARUeH
pjDh4PzQsz+2bKxp7KMY5x9fWIsay8+Cw5rNKFUzbrfPyh5WJ9gAhRCXknj0FDjW
7rKSxUdbUcGLuVBexrYmsgY04E+QudrN/T6+ftMtF3V9pyvbcow0cjpUnK8fqdW0
mo07i0+6+OElswtlVjKvJFQ0GwQ38LnEjIhOihjD7yt5l+vZzCRHOed9MUgl/IWz
BSAVeGd6InkqNiRkKYrbrTgaAJ56H1jBH6pgPoSRc+hs/M1arrFS8r55kXYy7HIP
+40ZFqq9Ceup1dVga/prOwrRrc35ADw7QbL5jsVNRV/yuVXANB61hVYyAX4kCpy8
ajYEp927gUFbjTXzE+ptwiNARYHU8jxzn0+onTEh5cJ88N6bXOepYltCu0p5ZAjl
QsqPY9eJZiT47BIIP0WckipMfkZiwjYY1MNaT6PHkqCxXU9VhQvTjNiS1Dq9b1Us
YHtW9gKaw4Kox9n4J2C/O0TtCZO2SnGgQbsTDIQ95HDByIENxZWLuvNCvylWhKMr
nLQ9p17bBDBKm7+kQJCK6yylBPTcwbLjUNMcVFLevb3ut/pQx52sjLkAV1PJumX6
l9MgqkNp0fCCoBYIgnLt8JhVeB9ZfNeSuKINr4UbcoHGq9MP54V4meGTt6VsHtVm
VphDFNlb2yLiovLKOCrvSthRPVIkQT8gzGW9AMhiSJX9J0is7Vi87KqQQHTPkQwr
clxLlSgh4LzAFQQIMkvnALE1Yi17s6iwqr/QCMKkq71YU0InhxuTXag8cFLg8C4G
lshYkQhnL1Xx92FXEEjKERZnDleSoMeVXkpmSkENgMCyFk+zesYfGiRGYJr7aFq0
NCxMLhMdBol6avwLNd05jab1Mzg/9T/tj4vXjVLtTmjEXEDpnn46oby+iMuFedq7
EbmvMPJgzbjxxkQGBxqUxgAfes8MyGO09NMlSvbl7oSHdB8KGY8ViZ2EhapQoSx4
xz2A9BvAVRmb/fhKnN6ORDFl9bpiKsadLNX8enrTBbnBKsglSU1nq0iXjEcqRhhJ
1I8bfnsDGwTFJh37e9ayDNl3Nwmf5R1zF4dVwarkr8uqsP8xVIWfnpLpIpSQZnW/
fR/JlDoPBF5bzQooo/2yNu9yxzy0fYTRlV5SOFFs8yGiyr5AP2GsdjMp4Pfi5DW5
fEBe34IxPEpjUFLIcj9uFmosgF5IyT0mX8K4CEI/fNTvqUoh9sewCe5pDA20P1Pc
VOxJelY9lfp3/KHiIuyBteUO2nGFq+Q19V0uMi4QEQTLqjYR4M3G0Cx85yx5vHNj
tM9LRmdiowDwpLHCgRZ+ZEPCHhviLmJUH3CAexL6axHNBaXVc2eUihGg5HR0EH1f
fdnFIkLYUrdvVCYEkyYB1cspFFuMZVFE1f2mrcBtJPDcD8nnUb/XYLKVyM1IgDPq
s/lVHspNpIFbe7Azak4Wae7AHs+bonZZsnfRDHmRa/XgDZmgjGBP8fidALm7xxOv
qIb6uRXtQRyJOTtxZ5UufpNE62JiRL1pB8xUSYl+46vtgwbFyquU6liyp8fjjAUM
D4dUUIl0ba8Kjpe6wEjTsqzy9JTF7ULgrSaebM7WxoEYyJCRC+R4koNwWPBnDbqe
qVQ0I4D3TckaK8MncgBB78j2yOWIoOAUItw2TAsBonDKaHMqvr57dj4ovtkhjK5+
P+qk+e74B1qkf85DCAQbZZueYO814lhthKHYKgK59ZAJ//Dcl4eaH2X8IqYrVivF
+Lr8iRmZ5UX6Xap6RJivHQzFD0raeMJHuuU/pO7GZmuvcVbqCZIid5ZAY+eJSMzB
TQaKtRGpah4uJqK3hQm9vg73yhw6apXga8bOWufTDPYXWRdBiZrgbcmHCeh6z2Hp
8bHGgaVqh9j0KCLTo/U+moPyLNkSeGMarCOk+e6hXl4crChccGSKeIHkVoPKWk/c
M7l4TIlEW/AM5nCwwbq+dXVmRbcw9SQtq4cVJo3F6C2tBYk/XfhU7+PfywKIOFlK
iToeO31MypLVffa67npP5pBVZRD9nHARClF/NIuTKNzE3TGT87odx3n8mFeuXaQ5
3w0wIGOdR9XZD1M1OnKsi5rRIu5ok3MfAsj9nqjIxgRjSpPwZG72sMpwEDIfd4gC
EynWDGSjyCOoBmNg3WDqmsFLiUU4tKIVYLZqAW4nYgqI/JVO0ADL0182Dw/Uz/k3
c6BE1br/oSbLJupIWSg58G1llMgLyHY9wkCxdXkYDBY1nkLLDpcMhcZEDqhfdyNL
1bsabiAH/L71XesHyFiUqT9aVg511nBVyG+AV2m8XxXZIpw7HkWie/Lf0yaT9IV1
vTHXyFZy9DyGQZ1Xculo3Ru6Jhq4xo0vyeYw88okrrAYlJzy/njHdtsmFtYAKCfs
0y25lO60gQgV2N+inNvFkpnuwaoDY6dNUIHkQMbFiSqY6tIE2f81WEJcLdZ0hUc8
AsD7m2xz+KPSTzvuwvPOXo6MebRQAKdMn3FErirCixT3UjQ2W/zTrEPVPMXm0szo
DWJoJmlNxq9frXEbeCtDbyJ+Lv1L21PJzygck9fSVTmaVmpSRL0ubB4asuOpeXgc
S3XlnLCF6vAmSTW9fIGVsq9AENUW4qppAr8gA9ZIZqaR2iPV6OUP3Y8/YuBgrXX+
rL8t1tEsZ0gCPykXCyNuC/ODBW9RVKzv8+tx9Y8DXT1hbrwOICq1ulxYxAfT1oqA
w11cj1m/eEfQQ1unIWBf/FKojSxhVW6bXGOAR5X5vH9JaPS92mq8oco6Gw4j4PNM
rB2tjWhSp4Jn/nU3Dgl5zCjTY39i7FyYJKnNspjeg8yrIL18KFd01uFT2+nsKExJ
FPwMNk3o4kw1qufEV9n8ifOJHXJqrquAbYCt/n0no9EOHxic7lAgv9tt0sGf24A8
3fYNo5JUAVmGgzcH0dgCTpxvExksnthU4ROASoW5gzWS0s1CagRw4z+PzuLcuh5w
TDzQZaFx/QmTS4O9aINpQNiBSI6snWckl7ciM91AuioIn6kiZuqj/aXgj8Wg9O53
uS/lXkuQbJlNnAIALyeMpk8x0Kd2uv4nVZSzkHPw/e7PxeQMu5pBek96Yk0QG7Np
ZzjQ8mfn77SOL4zt8NNjX8HyVWTO+q/mPJtkjVP3Kvfv/xoaJb2Jk32KZYi5ATkO
n5dMvjQK/mvZN1n4A78QMjVehsoOmIjO8hCSfg/IX7NSwJs+LTHL/uaC6GQ5eOTt
OcBQnNkr8CFRvRjQIPG0XVXiKJNiyMDMIxIS697X1h9MPzWdZZaisZAWyLV9I5/G
y7tH2AZVbsHuUMvd8CAZI4sRHHLcCAIBqWW6yOjGgRntYkpWqcwqPQhIjJhAQjkh
5scSjWzx7OvuQFr3c4ABbSrkQS+hkVdsE88Anb5rTTYrE7SCFfInBlJ18IyXEs8D
sriO6ZB0NMdMjM9BAnuXp+UISMnjjRyrykE0qcU7qcbuymflvtak6RRMWfvIVwbx
zCYbZDSyJIwJUmUoIHJ+qKnfO9KvooRY2jplcp52LXJaRLycZW31NPyxiCLakcM/
CJaUkAULUPZDSBbZ9sA/dlzXVFoRDXdx5u3xTg7C7mYGnBtKb5zPiw4KSBlN+oqK
th+UttC9PDf59lx7pi8HpTJGiYXc8UcsHWQbAjdibXgDaBCTbs5hn4VT8VRIveZ8
N9p8T6rqttpawxsHLrWpDEOCVVFNW+A8NGVoZg0xdylBjjlkOY+RC4ZU8Ln+RkxB
PRvm+LY1qX0+BtI2nxU2YCmWAShBu63Mon74jw8mbQYlxHMqL0XGjqp8lx5Uy/wD
Z6+SahI7Z89wmrBZnWojcquv8gJz9WTd/vZfBwRtn7UiviQhc1bLJEhT9He3ZMkc
K8fYJjjX2CSa969+XC1phcsxfHRTDnstQ2k+NgXxL5zrB/pnBzjKd4Vn1xRX5kuW
UTS8AiRB+Y7hmxnUxAMC+NWp9+PsAhelG3JFBVNdXMJvHfaLUEAPWd5umShiQM6a
sEU/LgbNvCg4snbUwVM0B2xpGm/wuYwiWoQaFuTPCFr+0n+0oTajJDLLL5qwEBXE
PM5mSf/Y6vHUKAI8j6Ydx9czL/MYnqlbVv3CKbe+RtiPeMAH/R0cxOkxOoiw42Tf
vlbVqR9eT2Q8CYIp3Drg90BYOViSIA5SgICl01v25fnlTP39Pt1oONQ+BerpAvtP
/XsfRW0wlEPoGNDK3oslCrmZ4FE3n84tuLJzm2d4v7FyEG1/Fh+fW7RpALumlvEm
AcD38LROhh02/BZg1TSAmcJYsKDwpM8PNkmd/RBg6jtbxDYG+aMohTLQ4lD6U/Yb
VIVR9bTDGuBOoGahrkeIVCz0b0HNFd7Jon1KyIDYOd4Y05wg8Pcr1WN65E8UWQVj
A7rFJKyrIl4+NAWcQbXNB9BwSGm8jLV2tyaHuHFx5idABOzdGBnETwDh2p122l4j
tLhfiQ3KiLGgHaKGGKkvG5nx4/nWPZ1ZPrjVMRRdXvE5Uud1COO+TRKYbhnDzE3/
ZAsHoYATu5arxPgjt0C/v+GK1WgvNQVPWqoUl892+O/yySxpXmPDVU0HPQdNoq2F
hJvDdRao78VRqbz5iA7vYU0qZTE37mSlyVApWSyjzl1gWPSeTl/TBIfUxFriwBN/
TOvFrCtTOoThq5/b0D2XVLZWHeVb6aHo7TH4N+mQPPKKh+qyFfTj4CMNMHrdVvA9
pAWj7gRbjKi1elQed0QxPkXO3p0XdYD+XVlGhFlDNYjZ6z2Fb182Hapq659+yCEl
MPGTQ5qiYKCcl/e2JmDTwycxeGix/3qyYgKzjjLf/U+R8Dac9PffikiytNTo+hxY
haB3Gz5671TfLvq5VlbHIZ58QL6yf9UlxMsn1lfOtCaQmLjzH6iRBaeUbBOrONoy
kUWJbIKdwl4PpdY+tTEmucIivyob27mGXdPICU5VoqF5vuKXwmwsvWm80FmgCnsZ
dEz0g73mgFr2YVv636USMW4OhIYz1lIlHdKdx52nvS8Y8DwON+n18qit88XKe11d
ZlQXnXHdKhysk2DHbvKYIM4Cjc456p8nR3kaKm5b0gMr32hJ9L3lHB/v3VElMmbr
B1uOllmekN/SHCxZyccVL4AHpRnnbkP+fkHqPNpj2h6W/vLFJ0T9YpBchpt7RYe/
UWTJh+ea2ynsSJMvOjTTFnNbotw1FBWfSyRkIQMJGmL6M5hf4xn6fq2kKcYIixjE
iX4a41A1o27wHhI6BDryi2ZJSUCMmSuxX0YS6Rww8hEg/2nIIXwMq/rhU121tbph
N4T2kgmC9ElAVVGH7GDMeqxcLDhFLZq0wRH1UKUmj+dGRsuXfVtIP/M7tyri0pBo
TltuF1dH/oWaGVZ/O/i2X5AHSTjvKKHkZN2b/w/fxsSvTRFgVys06iOPudIcliDN
4cchLL7tP6+n+Iml70UqGy5qRnRwPrpcDAWzX1P/FaIp7r9DQdNDztMHjPi+dlbH
65Ils2x2EkoJrIQ2F0qJ2EkSLwAl+/w+Bg2FzB3V381qexetJFUc188Q+nTDskVZ
sxXmemO0vNQtfP6oDlLbLC5V93beQic9qBTFVvpPAiMvZ/JLMds5yzEnKI3Udqm1
VxTFOszTelysfAXtWPxSjdaSknSNdAHlzs+itAUH75YA7rTeYJ7GMmEzHPySZOkA
lfr+2QTZ2pTL5ugHANhQvqvuPLOtzO5SDDVux7n9FL8FAMfRqhyelPhnhG02N8Ts
BqCJ21ytPnGvcc6nbAs5c/MVaOsJM9w4jkOAIcTjHzPAEzq55qE7zg2+jthebJ/R
zTSsco6Nh1Sk+DfGL63aH9PpZ04EBhYSRaU12/42VrtfXkpNq2wc3tXQqEhXnKnd
LxIbbtk2HVPdVYIjmbA8VZIsXgmnNi9Q7nv5kRdlsC446XCaS2bUztW2PB56FQRc
FKvHxL+6ul9icLx74Ajq2Hxz7uAPwAkVwVupR/40iBNOCkE2kQKRM5d8wYf23F3Q
NtH+/Z1JGXZXHgeESu5uh8HORBxZxRpmZMcVyKamx444kQGefeUt6CKuCpa7bx4n
h6Cj+YmLj3xfyRfyL0548Q0rEWyXAkIicaMa9DTxAFi4Y7MmBE3cySZFCLoOeypQ
GAJRX0z8oUnm/RfUoTWJEYp+votIwxoLXn3TSGa6452mTGkvgte1YlDoMsc2XslC
tliuqiFj448a5i1x+hG6em/BA3g2nP2ySfKL37awUl4pYyUUkcEbygHAb9pGjBRX
+PJ+0xgJ2kEv4eFWO+9uwsMZPfCcrq/flFO7r5eEZHnKVYxAiW5OgQ8TAuYPG818
JWW7FGW1fRCS7tRaa1YwSkt67u7RNaznPct3beY5tyTsS6Vm4njNRB7DNFIcB77G
BipmpvOzbhXpPVY39TdxJPWuiAtSNrKbAvACU8h2VIKrS63MfXsbFZvsmchaxFa4
s5UPch1jdr+V6MtY+p2SIm7quDzX3JMQWyhkBXZAp9cPPwU2mXW5umIdDBUvtJNl
CLzjE7ZeNm5fFCnjjLGk0Wo1yXRSGNzTCeO7Dt+eGaha1YK+O5lDNvbSCznhzuIW
W45wbAhouXhMmbqEjlT4A3si9kvBo2Tb5Qaq4+SNRPXovHvXeya8dx3+6gke8ahl
FYg9gXmGlD2EEP64Cat2MQ8UBQ5e82AhV/3YVjar7j2aaJmk3WMYbcsmmDeqmpmN
oNdk49StJaWher2Z85v9IF/YwLHnybhSfdPXrI0O+Udm0DzyFD6O3pdD3FiN9qjX
y7c624mRl8heMm9fBXfYdYBwUX6O/pdteF+RlMIWYzIszBBNKfZh5R4wBfCI1MH5
guoP5wrcYxyiZuG7TFCBXLOXW1nWRtDuPUFZtoZz3Z0mheU8s/L4SToDSpQqrfZZ
SKba/xN7yy31HtlGPku1sBW9rHiwBezs88D+WuJ/BBJ0igUJ9hHIJReDrl1GlO9k
I1SUMdVok2wNDmA+vn+t/ghbVLdc1r5/3VZWk5cF41y0urNfIz3HDgNGmMUUX0KA
GglBkPRGv4fAc7utQTEmhi8Z9/o08JhSxPIxqrdqhR5OwbpmCk8cz2ih8+JV7K47
xI764mwL/ahHDLAqMnLIHp4O6aHUfhX62siZ28xFhdjFbquQRPvGg1Q9wn9HgmvS
UoJXIRjm1Ss9raW9w5wj60mNQppxzmTRdkqP1Lq7tTIrgLnIUjGCo0VQvqRn9oR6
HJb5oweMa8bUaXmUKxKGUOYdY0uwHU+I9Tkc13oAXGwe+krbAVfqLCPFzzaoIlhz
cpg4z2D5ickNpgDz0oH8YwQD0DM9qkUhnPD8Oeruq50tLrL/6IDJJO0Gzr+nXIYx
4YhiVQSnyXXWe7ye/Fflt1T0MtrWBPsK9JfzoJaI/1UUqgk8cLeaMiiY2EYFmlmg
XgnyJDdcmL6PmHqOsTcoBes2BP/LH0/JTGtUYJkY4bxHbiNe+z/fqHb/lRXpNTEz
f90Aejr2ArXnFnxYri/yuqbdUIY/f6q6zvAwXLwH6ej0VYyxtvOmJ84O2OdoIXh2
RdHWgMHIbURImKKEhXchl3swXM54QV/sm+j1zdK+Z4nfPXUn6i+ppILZF4Br6kaU
dDQG6LL4TbcWy6KXiPRQx1oRu23zrr+rdRznfkSVrdxunWa2wvEOIARoxlt+u1t0
TMFe3pzQil9yUTQM3ZI+Ut51b1hE6+hT0Z9sJ/ElwT/DBT72CgEKPdKi0jvQgxF9
qNUeOcWnZGu4ykkBOpXZ4paz7SByu+WnmIMHNsXxTvkMirdeucWs17NQWc7e5wp3
/OXA4rpNO3eyFJ/pbj1hn6No6s2p55C+OssFbDNXboiUcUHla6hpyl46vdBdD/iS
UHSXbtMQ2TsWARcoJUbcxoGFMIwCm+BObVi2crHbFTl8tPFh9FHOtvoeAtrBHuyx
cfFCxzPMZZmfvYy+jVSf9cUvHHPzUGE6JE4acra0aH3rtRAejqXdt69J9oUlufRP
dLA39/70a5WhL7ndJmvcv1xWSKbWF2thBK5nFtfddlCd2aETEtTgB+57FKxJ+auF
dr4JyWgTfJMjuP4/YZu/S/RT49mkzJNsnz3XxFfvSfPYg7HBOq5GX7RXGSTn/IoD
VpPDscFWaipM06A+npMCPnv4rhokMng8W775zCuuua8otTLALo4h9eBvCqL2kuO3
M9kbZNseHTEKnBN8oro4k80eHzl9fMXI5wLzY1g7ScCNZs02IG9wPHyXXM8Y5H4j
9U66+ncCJui0Vdt7SDxGfrusNoIdbEgQds0gLlRSYFcGUzSoGNlbhcp0Jb5tlUV6
yh7IqrL9g4Ldc7S2dyNOrrh3pHUanyUs3UkkQcpNAujtJ2In5vBR6Vv2eJcFiARc
myH3AiEb1T7Mj0WQxgi8HzVYVdPZxbLFSVkRsxBNogHqC7W4mfPHBejZlhQ6ZSzq
N1M38HBY5bU8LqEcgeU75YD+//TO0rSqRyo4yyLRUYW36BXnTjfngKCP0efaJxBK
dZlVAMwA2MN+FvNhKgqboNrIZF1dq9f+O5rXwqKPSWWGjb0mcCS9QiYQnlJ72aGz
FapRGV+4hhjNTEuEgB4LtUoILWX/3DHkgRJmLl0qyUh791SuVTGIwy4KYLT+mLpK
D+BT+9ffE44Syb7Mh5KYlsIEOhkaamk3TypzXsLf7oxCM1BV2egmtYMCihOxgaOQ
Ckn2WWTxDddyyhkFjlo/c+rZZkWkIhP6WNDMSt3b5eohGq4oO1nfCztAx2C7OGs7
yi1ZuN3JnCp7XuaANJQkYc3EGXLojD7CfmwR8X67NLYxNlGc7PFJQlwF9W60iwR1
wDGgkkJTBfQqJ5QrPgIwWSFyIp6AKIeL9YsCIsH+NlDWQNRQQzCk+y6nB+u98P5V
pgBbnIHGgRw9FzTE/vXuux+Q6/rsfPmI5yOyWl0AMmVjISCliiiMhn1ZVyi1JsJP
w5ivWDUX5XtsHkjq7vWTA/+v8bnKi1NYAbDI4W72At2iT1JwxLakWGDMG2N2710D
66tQndXdMDoAqEv7R1Xb6t1lfKPp18wrUsoPpuxlTgfmQNgixdSM6gEitAlv73yA
o6bZGVMEVDsFJYMGnWRlWop5aCs1FGVLZAfdzzhT8nG9buZBLEArJebZrfDReGUZ
CQGIXDAnekUGDltXM0Yl5CioCHvQH5GXECTX4wyZAbtSrbEODpP4LlCaJI7GAL4p
nyXf0iLW+VIdYjN3iNPwRycw4l8F5JP/kmgylu+PqVGXbLBHVDwGpkA7trJVzc7E
lMeriqpWdTDX6aoRw/1jcVtZ9NwSC3bv0LjiP6BFd4LPAbJC4WB1uiMBwgNybLe1
OHhMrsfHiETGbLByjVTj5aNp/vZi0GPhvpg4qPJfZ+54B+YBaMgYV2k1IbS2IKEw
l9Xtlcbe1mJbbrQuQAU2VsPGgVGFW86sabmGYJ9HkJXh/n++NdvIzpHI19u/hsL6
vfhb0+kHqOTzx9HytipfluviOItGnFPe9espm7ZKUzr0JhQC2Y9HVKgb1RckptLG
xW03kSAKOmU488FKWAtliPFiZLgzSqH1iMbUgWcQ2Km7hhSCYnaTI5juzLtJztaM
9SmY3+erDUjYQXYwnEzAGr8T2xXaEW0jdSd725RmHdm7BedB8kH44SDJRgyobst9
KbBer2UtNAQiUlPO+KFMQrwE5MFNQXWHuLMGRb0WvJhvtKfXI98nqtiexaL6nQTA
+vSYzShrM8P/uJxyJchadfPOBnXQUgQTFJkz/zM+zZi6JJKfWjsvvNa3dCys7nAM
RTi78ElmKg6XXK1Bn3nsDy8S1IXiF45kPOYtDG+EZVoMYbbGJnRGTjXWOjIdxRt0
UFMfwfxx1jReCkLMxMzC7H8Po3Wq2jYBu5MFaTFlHF5oPWD/ZZG8O3S1HmUe39S2
t41eMbNj/SpXuMgT6t4C7XQPHpaXAtNVXss+RFgwxihmldjLHzAZTuCuOWGy/VaI
litcOhdLwBxG8SRQmHteFvk1cAZiKY+LvSlbKvF7ty+u1HAuaAWCd1ALtAO1ufrS
q4oz9v35IBYEqYMv1nqdThmLjOysrX9XRX07VWOCXAZYyLFny1bY1B89Z4uTotY5
a48O2YrQ/AXTc/3Gx3VQNYZCs072Sj+NCIA6UVTPKzAMubf3z6SU01kTsv78S/Uv
9/YY6l3TxIF3Wam4nBpBu+nSXHJ5OlHKL8bCKKyVPYKLFa6zjV89hLr2tY0lfCzm
+ni2bUQaFXGOSNh8Sy0BvJrwsz6Og96NW4MFwAJ8x1PI1HRMaCFQM0+mmIwPgbY6
ClFs4udYgxDdzMvYGDaTEAysKX8zXiwX95q2yRpdc9hvZY1gw3gj9XRX63/IUSyn
EwYk+9g7tL6EwhLW/n8+b3LOmCM0TEcNM8qMBmdpdkPdm3t5Im+JFwyanbibbsXx
BnJE0sG5bgvZjACr7tXm4E7QAuJcwchhwadTv9UeenPr+OONEgWEFynYA5y2Zue2
uvYzhthFLAc2T2m/iyHq/71XOyZi4G9YPlWcN8sXDZAGRVumTvt8z1hQj82KyCjm
f16AgJNRGhknvPlmtHx4YFW9AvWVs5lAUgzBd8sglHPaa7Rugx7P67cE4C7yRbrH
3UKMZUMgqltw836R2Wbz0IAmjR1AXoKUfD4yFP/vG3UmQtAqzXUFB7FTjj2qnKuI
6mVn7q60YRX5qk5cW/OR0ouhJFrZogRCWv3VsfRnOirqoNTuX9A3pR0SxaUhNApy
VuuI9DLUhKKWQCFjp91JmSPm3iOvdEadpiEamcmnpgixrLpteJS7O9svJ71CDQVK
NG1Hb2NtzepEO7g6rENktwpK1BmDpdzSi9UI5RAZ2kDR7FCsIKp7Xr+Kgt/kXMBk
19/QaQ7ab/GytNHiZiL926FQFmHR99xsmzinxq1N9vzNQJriL452T2HqPXi5GdO6
wNqdwDf3mtMYX0NMgbZuQG7mDoz8vcEPlCaF9UfJ99q399PQWkLN6fpc/Lz0nftR
s6OxluJMAmUq8xVt/rV7Wa1sxLT2A4JPB4dCYdla8So6IV05NqsYUez/oMMzjbEJ
CGgU8a1yfsipwLMzxWKm/SMRyW7vvr+QLcGJGaHmr8AI6w9uLP42vNKhVfUfGZdg
uUnWjrOfPo2TiGfEg4Ddm7bXPK2/b+6aQqGkyE65OPCqGM8K9+ux8dsLq7Et1J5k
v98tIDC1NyA223Cf+v4rbv3A2nlFAQBoiTB/jZUA/CEPFNNjLDgIUw/fsNz4y4Oa
YlfJDXqUCQz9Ehl/TlFuOOVnSy2hm/PyiYEaKFi98+8GQPoA9DNZRqJmI5BSGl7w
6Lj8zb7HQS4DmXJQnOOzYfPoIto3CFOPAyShI8tpd3LAJaWFfw1nrZPdGykR69xi
KYb5mRcvVyjzI+cc1+RtGYPgGN3Zi8JDje2xuDrWurX/yfKttH8t/0f+1p/sr6UH
rPk1msKWqgsmio0KWimZgn4i7cBDYMOxLdCUhlGWIfblOjb0ve7pfDSeLKp5/Ped
1XId/8Kw1s2hSr8k7Vo0KNTkjFecVNAO6wPrpH1/qYPyoxZzKPoEKygb3C7r4ZCK
KbRa0L+gSf1v168Iwkf4ML0Wt0f7fMRVYX0a33zCKVJlp8Re1ea2d0W3q8RtjL/c
izDtunbj3jqzAxda19aq2gHeuupVldD8DiGtSIQ9FmxtcsUvmAbT3A3cwxQWqj9f
IQO4UcZabQoEWHIh3FM7bDldF02ReUlYkP+/r5mQ0Jm2gACumuv0qW2jctwKomxt
jcsa5WMMhEHS0NfVCqmDCQoHf9MsAYwFKFlkntTv/lec4F8Cu+EeYjsnW5N2ZTu5
H4F291aQqSPfTEcXbZA1u6fPM/HxhOKDdhr3NeAg35N5P7kaRkmzzqD0TtMVwc+E
ZKLJ3+VdbdXv4eh3iHxpjmqi7xZvhFHgNYr88HhwaCrICVPIEkOsSvOmZxgOigQp
EP57Mk0TSUWX/aJHjTiBjDk9qWw6fU0a02EeJdqyEygPDGa6xH1chBuCOGX9x4e/
rDRX4p4o6mQv3cdV2oIfFLMQCr4zRQX0mLNJgVqjF1wuZrS1llnXmt2pGCRmmKva
/Z/Mfd3CtMwg8eH9Ixs8qzmcu6e28OPTR0G+uIJxS9Oukn/0XmEmvuDtnBTArswP
YsMvY+2w3fa6mW1lL2lOnXJWOcOtxK/ege5qnQMMqZJuk2sB7fm6GhWDGi5dUtAB
qL41s56P6kBPIcxQurs0D7SBTyKN3lp4ixvgbBYyAxSGWD54JlBoiQftTI375j1q
R2jA5LgUKw7WMllgIvL+ChRIIRH+K7YZMofpXQG5AimZAk/aKv1SjGXpwXIzSNh1
r8mS2bKl+wTKAnmM6L/1NeEnb5JVInZDl9G4D/jOUWCmjBKuvjQz8OrubmHmG0MU
Il0PPwfr16c0jbGQHw4motUQ9A1YYnflqO9FMGoK0Qm47gx1+soJNKUaT6llL4P4
eqzG7AOetPCCW78JN4GzpMLz3JhYpoHW2jLobnmw90F/AyAVtfntYqMsxrlweKiM
qC32YrdfI726ulcwkWmaYQFEUlpt/FRpBxm252C+aQdIF2ygB10Wyns0Zc91ctAK
eBPp0sHTWUsLbOCLUvHa/oJKxOIQLFQqTD4xPPF1ieF3Ixv/4W9u7/PPZCTK0vZX
8mhRx80v7WTAqm4mx9FoHSdDPP4cpFJxbLmgap33MwTLNeUb8YWcRrcU8T4oLwMr
VsjFo8KH+MBULnQiw8br+9UwkJjtkaMn9mQAMkrVQnfsP9CZwcpH+M1RnvXpfO8m
adeAXdpRT6LaROl+VSNWUnzsrRUVJG0lDfOF86QuirNLAjbWAzbYKZYGUwXLt2tb
DPcWTmUntN9KGL0UXYzBivWvAKy1HZCcW+HLTndbqm6nzPLd4fqNclkE/PZBIrWL
UinmNuhnJyOfhtW5sJtV/JjMNkDzxtAgigcq+XXPBLzalo4wpls1x/IP7o4XFMsp
uU3snccmr0L+MZYIoamJMt903x36Laj+qc9Kz8caYnOPocvSv1TQi7ZD/3fdoKqJ
SW0Mv3E5I5uNFv0ylaK5Z5ycVuajgwEKARpBWpYh7dwOr4Hp/E0gYsCvX9rUj4Ku
VTyizgH7dnE/vWyE8jwG/cQ3T4x2DQEcZKF9Lbxd/Sk/UcJAb8wuwAqJBNQPBCBk
y/mn6q4+vyfsWchx6z9gSCvtY7ZK2GORdlkqPLeYtH3L7AwDnE5CefS/LWBBKhw6
HWPYFC1EhVMO85idIxcC82ULcm2ggTvpYFi7E2EbfZfpHzhnew8VIboEtdZKEeBC
hRqZmbEsF4Pj6bVx1Jk4HvpuXk6cmK4MNcnJpP1bdGiq920GnwhSHUykv1Rkvx7p
70XLc/CF17zN9dlgY+iVgD0OHykp8FnHAY0wZZ2A8XY4w9eB5Vb21rWYxfMj8Onh
SMZfcT/F3TVJDldssHOOhwmj6yxtq5//MVccEi3PdSjfU+sjuqbf8t0XQrMllGBw
2tvHBxIFH1fRRhuBb7UKLJ72ygJSlm9fCAdyeZ6knhwnfrOZ9Dksn3L2cG25fVjm
BEohOeRusxbH27Jvqi851Y7czi9dLAGFWci2tlfaxvGNhDc7whcENFoO1MgDxweT
0+l1vYXYUVL/v3sCCbwF0QZynRDX3hYm/oVaOZJCFn+d6EeaJwQpcc38buBthj2p
k650adUPdSg6uzyPthMkZBdCWHDs7VawpqCwET2ZaHScSAzXUu9VrNRERmvf48rb
u1iT8b58KsNOdVyrRGq+DoaTm+AcQgquV6Hocdi8LFbvx3/FVI26LM/wuQEvqO5w
2FydlKvG0xw/6Py7RSoSqj2KQWDCpT3RZP1sc7VtRtWGY8VNWMj8+h0gd2i6W1H0
FyWHhGhOZCvB8Ghvh0FHwENiNlFXIJaeZb7H2by03Ar/lSB8nRN66HbHAn2B1lbN
pCxBR2R0MNU8vbtYTV+HX5BG8DiXhY9fE3O0Ktg7fyxgikY+JFMoiENDf9rvJ7lu
bn5tlUzN8q0vApgW2regimcXeUlVetbs8Yfz6eBiTqsZTlyNxYJrTsavFa+3uRpH
W+ELy2pkrsRxRMxvqZH46h0tzG0mPoRp8+pbb3W2TDnu5eUPDrNkF78A1PVflhdn
eH8VVO/8mRTLCErDzWz86n6+5ymyr48RJA4Bo5xCDEdNkMWweNMcO+zA87el3F6V
AJ56FQrV7IeUIzgz6+aDcMp4IVxopL/WKSrgg4rJ9gzHK9APD19EsqphHoxljYBu
eItwrYh/qOwsDCCP2kQxFWPYr74+ZdHH35WJ+so7WU4VkTEjYTiraNCcf/YSGDv6
uK3XQCFbver3cVtRtzfqb8cMwJZGt1FEU/uSOyJECodf3lo9sHTWSv7WVyNJkH8q
sSSyMRFIq2mrWU8aRnW8Xb5EcQKYkufTiWooVE3mMAM/b/KKc6nSoOZ2z9vaCcP6
9GdFWDoUNBXg1orGt9g0Vkck/a7pDvu87WIpvL9IJVkenYINc2Ef7Me5ld9Dqvj+
4p+WU/quiIqoj9C1YJepvDrdj+6Liu/eHGhaO13SGYcjkZ77v9zre7ggqBQ/5FSh
pH4moHYTVrUczPJ+vPZOxbOiFBSmCbMKQlvhreRIPZu0z+tLdgFIBRWKok0wF10D
88wdPM6TKcjHC4qO1MfCA/dYZWDApM/sfES1aBMaekSi+RU6fgnyY4mrimJPbXUp
Y0dA2ZFeBxX3UCmFq8a0t7QeQW9TtVHoDiZmWWUcbtrEk+F6mkk1Q9WP+hacf5Il
aQZX1WmGIUlb019d+TfzWrd8IqPv6I0hejPvh62Sui803ztBreR/hlir8auczRUa
AFETQ+fgd2xBcgxYdvcg66PtTmgjT4URYRUcwJrVCuZnwlF0nBi27Cn2jQ+l6hU6
L9PvmggIyUQqKOW7ceuHAsdzSDwo4JFd9DHxxu4H45wIBVJwqO9UD9bdlEGEQzTs
sdEJm5h1iVd5jVaH0VuluXdV+YgLZ4ZxSzU69j8DDmGVxu/D8smWYDMMvsi1t04L
GsozgHG+p5g/YYcJqNd0ump5FfylJUrHlVBgHDc1OnzlYYy0eEPRcFPvmQFigtiY
S6QiGFo2IO4c4qNvEnY+cZxl1gccHIftvDnRnbjesrbwO+cdpK+dCSVcJtcL+98k
JmzijSjmMw4/vJ8iYf/M03cOoERAhVZdwmEB/0PzNb/A9D3yXcgz9tGsqeaAgGUo
H2xPPTwvWZkVZshxuTIVBLCdYXXib8QaUsaveV73phurdJMXj+XeN2AYrYbBjZXA
S2JofbEthDiV9nzNHuQXRoANjSzj44mvplvFpY2SM2pdVHSK5tYvggVOfI02U9r4
9s0wlfVo6alLrIIyLh2nfIVydj69qysgzzSPWtkiPZWsgYPqI0kPq4IQ3MEbdBq3
Rkka6VOlxNUxc76DKo/nJOIdERgMUGegFxyvYiq6y4tjxO96csDpAxqX5UkNSjKD
5Af2Va6c4DpBHS+3HC6GY7BH9065QZqeXQzpX8Ah+aWVnlDB6hY1M1wotu2Vs7Qu
/439XXHYH34ET3nmtbCmTSqhmJVHNRdgV69eA+fOkUBET9uI6wgPxdaw9/nO/83O
HNLH3SUBCD9a0MThvuA2bbiZtqdRYTmHCRvfqsF5QadnE1O4mKh4ruslepl3ZaBc
LjYZJntEO0BfNTuPq8sSCqOR40Pu4jS2T5ptMhXuouCGvrcCPno2q22Zw+M+QfzZ
ABiTgUMr9mebmBr+2d1orTh0ZSmb4OsSuUVrZa1tBkBlBx6h4Cs6xU9fhhJTRCav
w3G69aqkiF4rqZjeMojW9XFvveps5N+FPwAbWNGvyucT3ue3RZQOfwlUep9kM9Ij
SrYXsIaBOoxcHfeyGYOlyF6FLASCkalKYctJGgccraxJJigKDG8QQAlbZm5wdfZL
1zxvSlcRnnuV7YcibTBohoaiLXGUDjLWEqF4s/4yB9bdnK0lVeHgaaegyLRKaZc6
PoHW2bl068jJ2pRmB31KL5+yoGHcJZl0KW7EqTunQarih2h4mjy8/ez3suz6uMWs
9wr1WstoG1Ii2Z3JoC1YPXRz2UqCmwX2eGLy2y/00EggoVU4zrsH8xUyyQcKtsdp
7DWuOf0++x1wBw+XOWBLHYkQ0G0XrBZDMzGSMtTaFk4ILMOCrmDJ4J2ux7zd3Jwe
zJOJCfHma9PpwvZsynBPZpaEAuM5v37+IV14ehYwT2qqmCUDXaK6PJB4dm7yH/Lt
MiG+D5BNkn3clOROPdI4R/UDMHDsVP98F8nptggO1x7ZDHnSSjm0yomGhAD57n0z
/Hc58hFR7NJ8enhPI1976IyijsyV1rJil1Mg4kgbzRnyae2hTfWuZUugt3Em/7wx
M4097QMM2lOS0V7FM9NzmYaOwzqqXrhLPKcZxOnR7FJbt4xWxVGkyQvMpKYwEFWl
15UR7yqxewwtmAk2hvZRRvfeD7G6GFmsZUzwqI53+kLRZwZaA4OukBE9hvnfi0Ta
6WSKa6aa8q+ORdw5QnkcROIjEkZySz1bwrm+js2X7ZvtRaToNZwNzAfIRaMfI8lh
ufpRajuvBxos3Cn7ZimdjlxOTywxq/RY2i01UJCubkZf+x+FmPmh6sCGj5P7M+o7
34mfKCbSS6PQ6fmn7Qw68BAX52G2llfjNbF0L2zWvgRs5MvZ3N+cmfcdhHgIKU8j
jN3SqmH6Y/5CrfMk3FYYk/K2EPT+qmAYXC0L1wL8cNUtfG/OVDTmD0Rosj8XRZMV
cf3MFJeB9+MW8lkcN4LO2TUmAWx6ZXMr5x+g9e1b2WCHJFaUUQA91C69QdKCf8fw
MiGMifYs3MfPi5912g4buZjGND8tix+Ol8Yfqslz1JB+yp3d5x2qhY+k3rHfo6jC
2VUxDA7HDo24G5tmbOCMrUXpiTnJg9lLjjplgAV+IKW8AAMYZ1W2I4+WifinDkDD
NSJrzzzaU+cuvtRV6XO8vf3E5FkEX+Tx2l+5hsX2V2PDlxDIhLCHf9Q9XU1g5hVs
rzxOS0RMQMGb3rj+8Rhp2Qf4btWU4KmiHEznCJBMeTBENYUu8npOsYUYZ7LcchLX
t7xvryHaN6DgurOHPULfrZuvtlRkm0t0ojioWdYydrfz4sjBSaGxqoqUl3eh7mzr
gYqp0znIBwFpDD6b0Jsnndl5YIU8GlZuo3/DttVwiF2aHxEHkVpqB/BdPiRzj1Cq
2TE/lVS1VBLVBYpXMOhhcSmKJqA9zgpSWZxIQL/9lUcxvqrQ5tzA72kkCyLcfzI2
xsxYTXTWJrCRq1VWiZ68NBfKmgHRp9ijkB3o/ZwEZfBUqCjzb26i359o4fkmLurj
QoqMziq1StF54QQEWg39ROZYO7+GVrHRMX31GoFe3OadR5+vGPaMDIJWcP8MQ5Ni
SyIPhZOhWXa5Rf1s+kilNyeWIxCYL9UsEtF+s0Jf5vaRNdwBY7FXgJk/r/+n01rg
cubg5Isb3mjzP0gyBUgikhLeKdNCOgohu7MzuaC7O2yTt395/FnxH4G3tDGFBcHZ
jGllohkkvVOWVfMu8yrq+eKtFRV26y7Vyw91V7d4egvsmHMkxu1m/q4C5o9TKx6g
wrnU2SJdtOpDRIFljew04TGpMGfwga7qZXjUNnP0TbCxwZFfmul+3EF3kmjz+JIl
ed2p5Eoqi4nHkMObqaSsv/6Eq9VscHi9NplpfLInOKbN460o2GB6XWgA4IBkuWNo
Bx0VdoYQ9IhlvAAKBtFYB/LMQo2F1wF9BIk1m3j96n6DvyMD3qaed80hjtikCLmw
7PvtfVU9571l2RGXLudUFXw2gYYaqzQXfofgx0s2t8MotxQFqQnsko0P9Swyze7L
u/X62F2skyo4oYlhkeEB3tHJxeYwRqgNNTJZR1S1Ckyh4qwMRFcqPY2ZUcxy0Bl9
MT/LklSwFP8Ih2HkyOU/iInPnBXxrfuAEq0/3dVzJGbXeTthVXHy1OQhTGQaXiq+
uFm+33vjKQvqSZarf5xlVj034T6bTOQYkoEXlwRwLegIQcK8qcapjUC4GPptkUdE
AhDp1jmS0FisBXM+xUPzB2nFErGgYDOCfy51bo6a7FwxGt65A3B+Q4h7du/cZ2tY
LMFaWKX8BYcvRDg06PHe62IVY744zfGpFmCb4NCiGGFz7cT8/+EqHT5LeQ4uO7os
s+rD8R0sNutcAE+e4I/qwxvwh7JFdmNnZmWI+Q9x1p6nJ28UrsPklNcFZLrTRWcB
fiBiy0JOaqfdqzYP21qabwjOjVZ0v+zOYO2TCoSaq5U7kSuHiHXbEoI5L78QWSWQ
bU38v6RbZmB+QVSByY0rhBQY3v1rf0b3G6pOGD72IOhZtyolmqI2JJxgx7RFQpXP
aCFwGfMXW3v99ARfokM7i3lZd5EVBQVzAuU8huWFRNh7g/cqXe/ibiyKWQl0yKSC
1fR4IR0wmZBL/6JrRbEvCqgQIQzSDpdzhrlQukvn1FaCfP4Akrxh/zQhrboSOHjt
pouAJSUhnHaxT0UVf7jhpCbHPt2nl6A8zk6iQAlt4ySdeNb60waEVRUA8JonHBsv
WFt+I74zaiPEbEGrIsmcdfVyp3wf24XAfqEY4NmDdbSO071KRBmJaH5IGghTwF0+
78XMhaCA3ISYaPvorM/h+jx498ZU7oOpn3SFRt2mmsNr77xXh2EmkvYegcV6Or7+
uVU9kobqPBrSDcxNM4+IvZFqSlyJJKKX47W77a2KfxRbWsx5hqFH9vUxr4jaoiUf
PSOUcqWcuebP+VQMXHFn5Ro8hh4gc3OXmFwMG9RUvBW05UrXXwhnUO/I32gisx2H
8wNcA234JfItg72qs3sOUyQ81z+hvPr/YT6o88ERxKM9DKzoRF+3lTzH5PAj13L0
2DJu4OSXKcly1U80qRRYLyXsWtu6HOG5KD6Tgu7stvC4dOKY0IxKwfARHL0tsopB
MUDM5nK6wM+W1QJ9fZX4VoZwMC9QRQ0yhfAp8lfNWkGay4E7tPio/ufDW7p0PMx6
RjS0+ejsIWXZlK0uMde17m7+fqY1Zyo8Pf8IsknE3EdhAPaOeZeSCPgV3IWw1dHP
QrVMub+BxfsuX8sNU6XRmOBjNPR+lfn+rjpkRr6BGlQH8EWwq6Qcxynm62qivyJM
hQGkEXh7FHXzcAeWCK/k+K+tVlGT0kvBW0SWjHkRiVq61LAcLkFtKl5sfp0RcFkz
YrZ70ImJb3UI+gxLMwRguEjhs5yL0DFq9BMFCfa1BhN4zCdydathjN9sLgfXY0kk
O3UI7MpckX69TidJS4sE1gZ5W22UMu8/FurXQ1GZ9CkGOxSp+bpnCtyP9y6YzE1G
fGYgotooMTP2dvHdvGlRxE+Vktxe8SP7eTwLPM5Tdqz2mGRZRaJezDDBwsr3v/Yj
q0RsUERUlILop+B8c8Se9aa2PQzKncCB/V/O090AoOJrYP6/0WZ7slnsCpK0ccLW
+WBXlRoT5j8slWxSR+hqGlSeVfE5pCf+pXHwkR/ieKBepimtdbxGM2zHGNJNAcxW
vZydYz8CU/xut+TfWWc+r0+7LdNN/TBJqvTVseGoa1aruWEnPz6cFnP5MmD/iXpt
iweNxD5D5Jly7BjG3OM/3UfIOXBRPd9l6CWdA7RrHJWm12+fANq0yj6xy5C1rZcQ
Lbh61p/8IyiDU3kJBQpvbhAjw1w1skrezj/R9lZd7BSRj5UHaqmagRJK82tQpgEp
Xf6jPyAFyDF5D5PSYBIJlOPSSRcO6jkPfIMHl3J6VJI8bXvWbfbaHAjLhsXiYPDd
Wo8Y9SFnA6nfSf6nlJpY4NKfxHRXXLjBGeXQXVC6nJkid2QjG5LNfyuMNV2cx+1O
UlT6HnaPMuOlXv9UIci05McSLts8DylIXmfoAI0y7tprlgAYaYLsubUrgUQIRwnP
lPYayZlBd1xLprSdNiw2Z8u9+0xjqtnY7lx7HQ+gBaor5VkKr7RQShKtYphQJC86
LxOiJdATpgSfJpbNn7JhQrkx/UVjOw7GY7wGf6UN/SU7R4Xuf7XmAOBlDKdIsHLA
R23MH/naR9VgBurB+dMn+pQrcd/BZSLS4EE4OUL5a0hVIYK0tghUj6CxABpOFOsj
rIltDkPwVK8R1MSq+/UizM1Zb7wK8rKaqcqE4aKkGLrfCrIL7FwHfIaBm7p4tDRO
jVNEAPHDzZUeWySap8HR5kCJWGoonyWMsnuQULEKCB7/Jtrb40JBYZCQSsJEA6Xl
nQx/knAJ7Q67YXRDB//qP6nNfVryCt5tXb+vH5R6kiyNnGOwqRffxFWO6vHAXMiv
pRkvS6KyQ0735o6bpjFcbLA7Qm7n+zdpNoSFlyMzSsUKprqOAFDeUXfqce/3y5O0
mTsDZ41lRndBX7Vpqwn+Qm6sETDzGQSyoAj+y0rR6xxdt2L3QmJhnN+mEQGOp3F/
Zei37Gl/tr1vVVK48+J1XLe9d/S8D3pl0VG4jPjfJBCttNoO2K2ILSUAlManFMra
+bln4SplG+x2bnQoUZQVEyP8XY5k5Mdr0bpa2Rw0xa2R/8Op8+R0LlaZWlOkDI85
5KWcdocTfTtOcqYUjYoCDMczo6OCvqJtbUTC9j6nRZK6w94qtZXjE+a8UBI1iGXH
QQmfStcz+Wg/YDYjHNXylIk8ybc1S+844gNQM3Agv4zTVO/iBEnyyT5OdwiesiGH
F9lL2HLq/R6eaqm+gFjMRTBuTIqFcOaKNPlQn3fTCYqMCT+1sOYayPbjwgyZJaTz
LvQ2lRZJGoCmDGWMtiJfYwLePxOpofbc7luSIlnGuJLzOP6aJbzw6mfJFg+l2dF9
zKTBgfoKbENBUw1JF1US6NLejnux6rUoBfyAKKqlVtG734qbKhCzudnBMsbKJuEC
nUiAQGdNfsJWWJR3VZpHMjn9eKFW+lTNuUdR6zdluxQzRIrhfUHU7tqy0qzXPI7E
PbVIDFIBSRgE/L9XQKg7aUBlZL8u7dqEb/d5vb8KbMfzLZS2WEFmM20zM08W/g1/
SM62Kp8pASjE8GW8Av4rCwxtWtcVpbm84Danzye0GyqvMkNDOnYRkXJRM2KLoT8V
30d088SGwNxoVj7AubmioG4p5LR6HHUiWSgEkhmhk8igjjBB+rtYaOZpduhm01aF
8jGBoVxA3hszoFxd2ZzcjovujMCXvTFIh/gspdSPJPb365mkMhpiOOgfI0mykJ82
MubNXOjAEDX1isgKJQla2SUjqy0UtoFkD/F+QVs/O+n0u/RRnwEnz7mRtqPNSoCa
+tH8A6Tpw+SPd4xr6lmdrdXJkOEAf3rlQvnxQdoqJ2cAMrvCal3MxwAl8MG3b8wv
PWTGRxxkb20/md8UcgvxV95cAKavbRYOkXYS3Hm+rmLnaXrPvixnNX/u+u1gl9Wh
XkTTDlZ3J2nQ8C5waGLb5wJyQcJkF/PDtCfdCRhbRpFDAJusSInm1o9625osp/ha
Af1Tl5NxG/wYsoDZ3yNbqI94NO/l33AsUTRU/r03++AIxZabsEeYY/2UJXMFu7jx
8GXFuSSrhzUfLNrnw7Nh8GIYjs9/TxJWR+62AZKPIo3hQK/xCrE6TYSBk09er5dd
yUbRfZIElbYDisQU/6EDG40u+aUJ7fuHZfed2snOjTgSiTvUBU9SSIFfWrQurT5q
AeTLrUPCojReQydiemITwXZfGfGV3Oe0dggXlwn+BYytDGR5xgDXdzsS3cRcPps8
l3MN+Vb+VuRmf+v+W5qKy4Qb60/GGiV462yOqRHA21tTMD3ULNf3DEAXGQx0VbTE
B9ydVv/WDm3S/0jUvRkuY4VGuJ331O0lz3CefYpOobOIk7dI9nKcWboqmN4eWYQ5
JlQlnjX1iuZwNDSqojnD7mMrku1s7QH7ghlob71JFRQBZXy4rcBTgiWA/BmD1WhH
GlU4OCoxJmQXaD2ipaIIxwWXV3Z4ynPcMN0NiKZ3IBg0sf5EtY7gauZvw3l9POe9
/xKtLT4MOPb9fUCLkrAJ9OwkK4CS/RlCkOdQSVGkgB4OXu0d4ehPNMxGfqrf6R0Q
I55vf/wwEy8NLanXnVmKFuRjsDkfEooXUub8CFGiuSGvXgMcOo0GqYR1res3j9nd
MQ4G2gsd7VLybTVVboyszchu0p5SxVZHUDJ9l1nL8dxep74PkYYyeck3XNE9N5jT
5K33cDwzNNcycH6O5HJbyMH11lzwYlwY4a7V56+5Wdv2rY6ojQX70A+iwSXtQGpK
6jFScNXyu+BTXs4yn7zOYt0Eqg19Xz4n8QdmT35Nv+CHCAOP3w5qBQAqtOUN/th0
+CX9EmjmkBE+ZDuWEOvsA3gp8VXaCfp8t2TYxEEO52NvlifdQt2PRcA4R8Mq946C
v+jhX+NXR2zvC/NTZz4plaeLfH9kOSwdL3Kc+yzSA14Jd+gNHU46aZYyTHRJSXUh
R5gZPExcq26/K0zqUrf4/CfL8oXa9/LvDZmaUV75hQETUTF05L7KPjVVtKyDa9AU
EqKAFRjDbDKBug9MBuc2pFYqhLquk27kB0XZfhsG0Ursj+JeVbCZhqhrBaceHFDu
u8WpHg48XPMlO+ZsD8TGYxOvb8+zEGHwA4RsMBFfl3292BXT1ub2yDuJF9QFGLea
y+2c+esgpvVjTaRyb135LSWSqWLIHEc1QHMHcws19uiUtneQXRCfC1e0mTYqReY/
XdQsyxZrRZpDbs7CkSSWxojht4rECl4tyHuVDV6kpRRsh1n/kXeBgEIxYuzstT5w
rJMxjnMXpMfKCzqXI7deZrNGMbOR9uUKkP78V1c3ib+H6cTJZUqyZMUm/uKevJap
5w5pl0HEUauEVxBqvWh3YM6Thp7TQTVvpjrG9a3fBFaFbaA3AplhC7dC1JNtcuIb
MT0ZUuoOxl1UT62ULgIu2foq7/aaGiyQMi3EKsMXGqRecEX1BkDRYOoQ74rBk2Nk
UIoGF7WjRaaAVUlqTXQK6csKTvhuTF+sgRTi284OjIBBJIrH94urpl/ySEvwOlzE
IDIfX88Ij0+GRil54wvlUpHToKWqn68uJaIXxs/yjEUijkAXgNHGbfXPHC5x51oT
E1tJkJzV0/yOdHeit0r/wSzegnZyoKXYly/4WUUmLLp81oOlGUe/d2NHMdnGHwuJ
8fbBsy3YpC4vgS5kxQgYqt3TERA547EKzYTTjhXiqDBJ0YeeQGicIvY0scf5yg44
g1WvYydEHBZbSD1kQJh2XoT0qbTmpneM/Wqd/SaAZ68niHCqS+mAGkDAbXUk1k+z
L/Vl0/L7HS7q4nCY5GAt26pcRuaAEDlfuXPQm8NlxOstUtFQIFGDU99VosDszw3D
rKlmydje2LMRMdG9+R2NoaQjOXExhWYroUyUuj2gQw1qtWa9Ok5x4zYbTl/vf4rU
iFJK+7xixUbiTLujXlQZHLnNUoOHhtna1dd548pBHSq0qjKGCFRGZc4/lnUu8nRS
6p6f/cuLxhelPVKa2IxtBlMYqAdaIM3dd+tBzhWelIx350ZyQ0GGHxscko2qKAsv
WxZfIvRYffguw4wB5pO2AgKVUeU90pOkfxvdEyaDdbsL+G4HFtG1/5A3r4HgfXRX
Ihpsl69PNxWfCck3E16IS5C2L2I84QzIPHkXMwt1ouqigrXFks5tp8pl6lL+LLLw
8FIbvENPC7SutaefQRqH+AKH98sEWxbO39sqdjTXFIBzyOgzFTW52s313f6fLRrr
uy8cPxS7XryE04q/IcsM6ZIamMaXvC0Vx0AIgKEIyoslgC63ESxKIIlCKS3mfCKm
MGPRmGsZ3X3k0DKEycK2V5Wpa/hC0wBwjRpMkgn+S1s+wrHr6Ke9PIl2EXykpVpk
nrJa+amrsVwF8tqRbowAm0V7mVAuLeiA6KJa2/X+X0nymJsNz1BaPJoUYEyruxGW
odvj1mvl+Vvj3RYKipAL8Dc/FXg/02akceFY51TbAAywNKrvEJBY7cadLcNO698g
GBQUs3mIhxl2I9oIjCMPNK4N8d3SzNg2fKdSpO9WhvGyhGO0lCmmQBl2tKsNC530
lBk1rPSPaklQv2mwn9wk+HqhuiKyUnZmoqK+ZJmfpkC+zdjX6W/kFHKLP/MFi7Pt
0MGt8byHTjOb9dHXBXRTGOPm+ERynW++1a7xGvgq1R2M3g55v7ZuJSeSYnonfDoL
sPeSDKD//Miy+3pCuKOoBCnlcuClpVwzAwWoPNVvitdERjTLmxXUcN/0hUYKTSrI
w8Jkerqk4d1tDVRo7owPTRG3l2DRrUDGBfD4nJUDwUGHznnNfidCJOvuIYpk5cCE
+vcRKDn7++zhtImHzwNdbo88kbPWxYw1cl0OcuG0AWsDCJTfrtFG4000iITQ1hr9
WRV7dw1xYl3CklWyq6vn83I9x1T6nRpjwXDAZJ6XlNvW+mMSTLxK+8XvN5r1O2j6
l/OgkB5Xk3n6ClGfqlur4oa7onu0RmvMnAAN3tZ5/KEdyrx8bHHA0RsHd+KsE/PB
kr27s6MIBAHDkA6jZQzWzWFgegioxsq9EBg2Cl2b0+zFRAxYEKlHqAA7xpSZ/t+s
Gwws4wcWlFqsTz90pHz4KOBpcV1+ecFZOPw3rjRi/LbxbPxbAyBIlFHoYVjRJRac
A1T0S3jVupok6SvEn20HyE0LwW3HADZMFU638UtS5S9EALserdm/36JXZfM/ncyo
CYMQBVKewJj8+9+ZCdGS8aBl0DHqURf7eMNz1nGwdcLFWBFKpPi2LZ7aBaRHre7j
0xE+9PPCm3Gz0NkhJc1foKwHJy7GR3wju03CjAKgX7DOheGdg7sbtJlg9X4CpbEw
ccNEj5Hz455nQ8FFuTNBiHo+8BgJ5wt8FgtjU+ueip++OH42Szd4T5czklpjyx0g
BUulgRHuzLqsuLeYAII8ofxtIMdzlKghA7uj1+pXKK1cnnBBaOLghB3S8HmIpd8e
+FoXY+WX/vjeJipegw24HL3Txg8akB0mSlFk8XyOYa3jZSLwk8RYRq2VB0TG0LOX
OO9TPP82ZdAHLZ0O49QOObJp+vmPyjitISnaUt9Mm102rlo7WpDX2n1Uuk4TL6kW
J08QmBxkK7QdNvrnamtSwk0jMdgOUbrUePQHosVsJ/z4XL9Y6WjIVqn8IzsoYITG
UdMls09gtBQnJPdV7UalyCmOnsgpL6x5ITiG5YQY7JGK7FSmNDZ6COGjLwOI6q15
hPlYVO7K9tWIK03tNEWMrTsZ7jhhlrn3l3AT+hcO0lPYG3k8TQm9i5Aha8WLLWVc
0aZiHcgAh9ylD8jqQyCeoSKv8v4kvqCdVdWtBOgLPsaIeJJLkoP+ScmXRk6Hoak2
a6Nyt5JJ8k2lu5vnm7vDW/gCnHmDxTuI+fuoxC6qiEQVoT+GQFC8OpUHX0T0H0X7
8BAzGSoItjWz8YMcvkac6uI7fAbLBYOjZINua5n9i/Ls0yiS4wEvAw1uJ0n28B69
VVzEC2y8oSzFLxzARZ+NiO3sCDzByqBsifRFqbMYO14gDlH7bs/hmFilEvztdXOY
oMqrkmp7LqTYCrnspq+SHvM/NITpCO4YvvBBEoryzylITWw8uvkkDVXh6ZwWHWUh
g6iJoQqijNcYXn809f6uMIMpV76ylUKqvlFinw8RLj06FA9ZXwbrkmE+E3Wzci+G
O3xF+GW1rBGR3vwXdjz0AQ7N8PlXOQG93t9pcldhsKrvH7Tj7i6755mgNn3G1K6Y
ms1fovG2WwCgmsGaffMd2KXKmzfNhreCyrVPJ7wA2Qhtngbozh7QoPCnnzCI0Mgt
BWanXVhSNjHauioIenPlwY7NnXUQzaMEre5gkQdU7SnIoqwZfeLMVGi524bdldSZ
n9iwDTtHhCcF94OBzgibCFTNFOT+gHSjbj7FIWS7/yK1R/uwpOX4JCaTYzHderwo
nuB5228WijHlELGJuAMWsqBOpc1h8whf/XOmUiaMBZ1EZKCEHtByG7RzsmMGA1l9
yj1wmQdC/hsMJz+r+F4tjrR58+uxaQlyaYyJCcut/+59DrI9xueaEjgvprw6rw3w
v/AD6XTt76eo2TXwt41bdwu1C/fJD0NZl/N2CO/X0/qy6vQuD8SFrfDIjVf/7fWp
xQBYtia1+p8eH6+g1XPWLTLbM5t8cPl6yu36/T/6pa/1sn/eLYG2fe+qQ/8ySR46
EnYaX3kqxyV/FkoRYY0oQuRA6Mg7u3qDMCb1EpYWfvI3Kn+whLPfA8h9KxF4Uopu
VRwCrUUR5LKC7TC4yjOFJaPxzvQp62l+/E6aW/AjS0p8N4TzyIDTkFK2pR2+ghVM
EiKv184iA9oq1OzgtAWnfdLZdGYvmbmanDgrXDYaTbI1+OToaztSYYyBL+Hv8KkZ
4bUvgvNXmWjB2HBINFkNVORlQnzbNet80LmpHZMtTMSUS/ArEHB38ygrHyBdRfdC
8p0T4tAFoPYKCn9TAXlHOC12UbfHVBa4LNQIJgWix1nmLLXtJuCN3ZPxrJNqTL7j
j5HkT+YHlMIMIYXQZy3jquoqqP4vzKCdfAmahXhiomMYZctUig+Z93wPeMZYH2S2
bbw5pXnCIVllB+M/ODt0StoCXX/CVt/lp+SnERU19P6lwGFM+nooVWv//uQrkEPH
l0Eeia64pFkJc42WLwASbJz9vijrFdp9JGuWA8qbpaUcWN5583BQPQP8ACkziEZ7
tJtnC5Wzow3UjF55KePYvJuGX6ECUYg0+6Qv6TjC+Zdl+aGRT/tpHiVsKAXJbUYC
dYko1an7j59zrgCJsUTrV4NLtnvohwEFL4pFWTftroa37BZWkqH9ekBF0CVsQOLa
f0OI84cbPkjIyDJ76o4aDAjG1X1RE1RA1Etm9ZONgzS9SKgG9KUK4h0lk8xWlCm2
4rlMgIP5Ed5SOGsIlH1Qe4FuxkRSsh/XSb6PNfhDD2wdTdpZeTfgyf5jkCYzCzs5
1iWFyy+RyPvFeelZf25lianv4MyDXFmPIu0YVZz1YK8+kRqOR+wgERcMOlPDdJuU
RLXBKGo+b4G5b6SHa2QQ8+37nmyvKXIYJPFi2cwqtsyBdyTT0saCstQqFORjoSZv
YbMEdudnoldFel2QYuyyarTxhIIFarStLs1eDdX5e3pSzIP4sGGOU+oVUjsNNGft
qcfFzsT2DzXQXLniSMVyzFwnFcIl+9KhaL/aj8g+86Jogm3ojP33xxl8xOSiWwnO
ymdKskoxbOZwKEFqzD1i+1f3LNOa1Y4ocjh6CgvrMBzJ95QLZdVHrMHbFF9J97Hh
HCJyGhmkOzHI23fhPUdR6Ez88Mh8NTqP3iFtc9euN7xP2Il+oC6EvLpUJNmKqaEY
9SFFCL7oWi2LrJsdPedFGLICpOO7rqekig+HUaDdASQTbguLS+NfFr2Vw3ghfpkg
5DnkH7jnNC4FW9I2cxgOXRzIHz2fqy4Q7egGACdIeCAWvq/jYFRoxaA+SvQ+13Pu
n5evx+0YCPSTlwLbyFNmWv9eBITTCjUwkYZjEhSEjmQre0JUBn6qav8z/JIEYBWN
e6RZ+zErLyqD+UM5Qt+WEkW8FGxc1jdyRZhVJynluIh7aQLXth1AL5H2t8gY2Drf
PSPa02uL5mO0Vjg/qizFSDF1hZyB5iHY+RstJGHRCsPbcQi2rlhw7PfhuRaSqlx2
0g+V3QkaRo11QGb48NZzPvwrj5ffzxkbwa+peZDpppDLjCmhyaBSfllobMbpVcBZ
opQ5HO1aXZNf5iLuJF2l/vVzNobj6gpHtR3ONC+O/hLYaWMTYMxgvfBdOM6zhogJ
DjrYuBMts4Fy83gk7vY8nrYVuulmA3NIbJWXqW/sN7gvWwt7HjylxeF/FG9chba9
Xeh9gOaeZ2UeHJNq2+y/NvTN4D7nLZPFODfv/0RQs/6vgObQnPA66jvh5lnxjv/7
6ywZJts4N+wxjYiaRmbp8CQ110k++bib7JXO9xoFQvaxhvkUCAy1HQ+Fi7Jl6HpO
1n2K3jXhCuuEqNV4AJ4C9yBsrFWqdkKoxCt4alaRtbzgiRvH30QdRQLlKkFO4Za2
qWWTRGUKpA/YcnfrdmOCQ/VBhA54yyKYOIzotOoSio5Mgfx/QoO9g9MqxMvVgGFs
bzXGkIz8+4WltpEopBF7A5daGx64hRa3U9viu/RNdbTzxFA63JpV0tHtKwgu2UGr
UREye8KfazzEcoxai18oCXCWDlNRm7k87gq4c0G0tAXgSYIpNI133OgYCN+B5opQ
YXIqNcvz4S2jfG+pba9FJUpk+KAv8MR7xOtd8vfWY50UIo+5nYiiDq7VBYtO6UqV
JKpyaag5YnJf7isWaYKMjcGYnEPjPpvTflaaqk/ri+r0/hjg+Vmd46Qhj/tCIMnF
Mo7nDRHMQCzx7EtmUTpcU00kjvx3hi6uOY71/aboLerVcetrkYfJV+dB0v5Ovk5y
b0xRCU45aJlvb6D18n6L9gI/mnkTd0Z+sLSde/1J6xMRJrQztR4Uxi97t/iKLMo1
zLTwXT23wcQvDI46Ng1y2Adxp3HBUYJ+3SfjO7cBwj82q7cQR8XL/eo+lnmUH5lT
fNl6GMAbtGl/huY26/PsSqJAVYLF3K3Xx6a29FpbbboHms+S2e8CcHK3aeyqThWg
TKp494HJnPqYVHQu5SV6a0TSth2jHRpS5uCizd0afaJ3D7iwWI0m3SyFgv8IykZ6
W3/ht7yrg73dRrZej3pOihZndScsmVn+a18scY3lqomvwcJKngpg14ERV72thyDD
ItEGizQag/HbmU+SSSwI8IFq1kQd/L5Vbh0SaiAvaCLAzUUQYL0upR33Zh4GG+XE
mbriSrvjMXeZ0g7Ec3OqO8AH9jDZlqW+lpF4d6pCboC7fSTCESd60G6Y04CG30kF
/5crddu40/3civ0NLTMp8pwINflLgIkd0oTZg++FV6Ib5MtePATmYAsDYfhAsPAv
Bt1NSpopQMmIZ+OSW2cZ1Uh5ZQ3tP97xvc1A5r9aCJDnu94ZSr1yFIItzEqvHLAs
WZUlrE63+p00rQYMAeyd4Z42LFO8ZZeMDQ//YksyE/XjpT43GtZEcNdTR1bPiZaR
u29NH8QiNfMc99CkLu7CyZGNQcSGZlkr+j4yN06E6zU0/qogjl2s8/7ByvQWlL3F
NN0zXCgFhYNi3Hclk6R9vBBYmLOeE1kqYeQU8NMWRjNwMDp0IjUo+gzKF8x2Svg1
4GhyeBUHBEPC6i19CLJ2dI5k5w/6EhpLM4wfxEQtMSQeheU4NocIrj46WS2Q1oOK
1ofMKcAF83cFgOCChlujgpeVWlOXo+lhU9Oj/OIIsI82msj/OHHot3rikTSeRYNr
bOfqbOxvonXYeMWlem+BWogWlT+qotCgrOhvO0H9sRqNjGUgrOdWZZDolO0zS7/8
MA9g7DC+Bor/YCtFSLSavDhAzNmQmWSPm0SAfijM8RY9fLXDYObp6uC/3kHUbPzz
BFza/Dh/pywsZeyJRX3cga2961emrq1yffyZKeyUdc4riFnu/svuvzaNU1wzMHgT
Ka5Dn94jb454PLwExsBFFNVa6NOeHlJvoW/ocrPlDct7TGLXdhWDGstqOX7elCaA
nu5wBinQE7VJDo6L7IXumfx6lbHeFBf2MQrHaPZUp0DbXePQ5bUuATZMIj6zar5X
Y6CFOvClWV21dfscvaE4S8pvImIySyb4Ccx6foYKLAxLwcG92ti2CigM5foI8tuA
tlFAqZYOMHfJkZf3VjngVcmLaGej08R7NuHbYPsdzC7D4wX5hvtqK3tyApP+Klln
JaW+/ffm4b/y8oJ0pdfC5gKq7qilq/PXd/843Giw+s+oynNdPl/z+eCwPvr3gOf1
0hr5DK0x+QlsKWnm4NYvpQBuYNVB1hR3FAW3mSUHnOV7to9H3l05jLeJpyiEKMr2
kPzzUgq9OgCkRMaGpm252dmGX7xouzpH9nInoaSbx72ZvA1DqxsuC9724mZFa72z
Qxt18URAuSasVz8sDVglKMUef9rht7bUbJ1Pb0jqISbRqMP4oUsKSnby3IPYCkxb
d680oC+qd/vDYQAToN8FgBnboGfotcyM0F5hGDvQ/ZXulL0eZuzlG7rc0qGCHo5s
DTLLSFOvY2mYwdSgv778t7+SwuxMlZLETTc5cKCxklXBAKDw7pVLDuCifFS5WYTS
WBvk58cpr8NGHiuWLiDS3apyN1XzRTOKzS3+rrBo0RRLow+HDAxfpcFmaFLJ8+9u
2lY+XOMdPwLlWTFB8pq6uwv+2Pf5VcLZURdkVX/7TvqPvTrq+eC/Neiv5QxF0EM1
pGmJBbdA8GfF8KWKbzmTuSiPuujARZ6QDydGw5Aj5jMy8ZRJyIoJrrakm4lWI23r
QHIFp0mMUCc9XO5oh60hqwHljSBIaaZyUByjv577Bhc4PzdXjSErKE9Nm2tKuLDr
FinLWY1bdrlqVViQBfJhy+UoJkqfRe3H5BEq1IuYO4Ehw710qSCkT6RHARRZAsIg
UBRwH1Suxk0+GzpXlsHY51Zk076lfxlv+F6urCVhe8MzrroSj7nuysdm+YRSLiYQ
XM3jQLVoRuIs4nHwOOXpdS5pOxg1IAGRfQAjorqCM2bfl6wta9j90FZbkwXkN70s
oCYQOt7Loy/i0N3LWqw7T6u2TErtH0k082Kwxt/U4J5ExAvgZnAQxeFDqlo38Rqw
/La0rOK2II90yfPG7SWvIrLMKGPhWEY6ENIJLnizCxAhj8gky3mSM+J8pDWIfI9l
EydKMAfbTzOIUMGyYV6nA4rvG5PtiPLNUvZVFprVRbkKYmajh7ww4+veNOBlmDAa
WtYlnGZmJA0fTVRPlkzsbQyKP0DcBAG4W+/uKyQUWwI+HGCxqf+iD4/UMjFttTAy
8FiviEK5SuMqIoonx9PIL1htjnciZDxGlxzHvig7WecXAxn06YSd61urjpk8179h
dTlM2zk38cQQoYi8z0HnU47JGnnHoZ/h/ZJWHXstvbP5th+CqHrN6PK6teK4KHDb
Nj9OsxW/Q6rqVl3XMAmihoyrcJTYTE3HFlaitOSknCUhqhESJ5GWqUzHhAolddYJ
Sj83PZ7AyswGrbxzP6UCX8Aex95rUtGWmPaTwxFZACtYqJuWfiY6R8r0HaVyXWKV
4vY7Afw4edRCoz6qQ+3k2EUfcerOcpZ6c9FnU3OKaJg7dE5zE2jMaw5yU2TzkZcm
U4hIU1wCWPIy6OkReP0KLVg7A1F1j5eQlYV7ZHXckvzYg5WXiTcxajtcy+Yn7WCo
Ae4gi7iC2GSjnS7fFZbmuK08Zwvq7Sx1wRjv+zU2UVNTLZt7IAQZU1E6POrLfwd1
F91dwk9eDH/FALh0KYNOG/jAinqEzvVe132jO9QKuRC4BQQh4BxRtbWB79XgjcbK
xQkDnCthWX0MiyEbLVe2Fx9zGtgM0VyHquaBEaOSKzE/Niq4oe1pyqnQv70kF6s3
HXs7LExaJKdEk3NHnIOOsDPg5tbybT8zV0nraeL5YbxMiov6GSS67ZRwou/5lPwE
ZjRrPXWjQgeKKFGYIMCMdM5JhloahYi96Ag64ZG7AqJnxBMN7YTlaIjmvLipfD3K
tIeLWagowCcNv+5x+1YM/MoYweed/F/bqcJog8ZAAw6H4XlZO5x/ULyzeF71XW3D
MLYpyfm+K7dGtrqm8xcIjqc7UHG6ukCGtqUsGwEJyx/IFvUFp2QTKpGQSDxHr1eU
mddlUXpYerIx5jgFetZvYIfvxiDAFL/uX1/wuO4xK9NBJFr83XorfjaX+ubZ10oU
HstNp3/sZdB9tbaCDvHOrQa+WQPAwA3lSirFAl3MQrZNtcckedgi0OrNyL4ueIb9
ByCcvECdHfhGyrC6L7L8C8WYaoJHRKxqOPbBaI7BmDmV1NKzml9eMqzh/KZx3Mmp
CPZZv5IpYYXsJNl6pOAo1FTvcD0LhLJPWRWLmNOunANM72YuAviOOFb7wtuKopWu
CIkhuimz8gLapPcK0ltdocEqjXkGcNr3Y3X1ug9GZHZ+0+VNaZNJOWsQuF89Dyoy
evXZLDVdrCsKB7eW4Uo5tZ7GAPAegIYBh08AE1HbIfAWr0zvPVN87AyFNvZiEpLS
hDbDnhu2pOhH3xKAih4ZqbcHt4ESVkY5cGswVF0TlRlJz0Dd5lYMYuWId497prTu
rP+Qw2voee7blxjpUUzn6gUhN3cTQoaq6FDIPPUarbg+cm6GclTan7rabSIaQ/we
0OGECF+QrzSFTbijeFMixfnO53wkduJuv2nBdJtQ3UOEVxp2hahgzk0ziOjRehv2
IzF5YZD91DVGRQ28hkW0VyQKIPgm70cXqKnVPuhdXqNRRbE4RzDP9vbgqNyRZcHi
aurBl+Yp6g6BxPA6RdQ8ytaazN+JxApRodlHhuzI+AaGxACnFATk5aQ/Wk/JnlVs
giNmjSTnP36OTSSZBFBXffIk1/45w9K/q7VduUX4PDH4TqiXJoKtEJrsUhwS8Tbx
+eKSZ9DskwyfRu7Nef8ln3gNBIQi4thFsRwrNEAhkTt+DSlELR8+pEdbMbb1+0ri
A1LHC3H/LpzKHnevuaOi8BznN/lrPqjIdM5v3lJdCg0t2FLqgiVuPI+7w1aB74rN
Nnwz0fI6YkQmzCarPKDWLXY4NsYUQgZVLsPsyckeqWzCAklTm83Z1FAd8R49qLC3
KMvRnhbw3h/d6p3RxuSlvtx19ATnh9hJqvC/T1j7ZVNF2WLMVPtgsA3nu5jnGkzk
+SLTReqdDL3hI8bPc0rF8Nb1WT05sXCARO1BHjYvnX5pnR6DXQ95JOhs90wj+EFi
6rSJQzvFjYaGGpXeYZdcjVit8Fp69pKUi7RpsjnQMiKq1La8GTPVj9JpkziZ+ind
jcIKnk2udXcQvIuvKRsA4xWvwZEBCzCgkOwcSvAYsr6urb/ai2CGm2pP36VZjsZt
NHSrn0LkmGZJC7HU7mDkhhlA9uIlPDy/Y34933Hu3pAZ4vztTEIyolACtoPnPKhz
v14m8bYh+C/kNEgSH1592GbgaQJUowf9jJTspdlzqERP2FxoLyC4O6bZmkqH8o43
N7uzNokB4ZyvTzTm0lnZiDJEXYSb1VJ4QCSNav/PQNrSFNombEpOhw95vsk2Jrk3
o/qGh7rto6WpFk3yjgt9pGD47v60HpcallIUTZFOPtXROx8S9Jaz3IiEQjsG3SC9
My/Unq0whKwfJDRmzQNnqSiTCMQPUFA37uJXFPiPmgV3pMeVDjnPEt2MYads5dHc
BRk4Epfgtfrq4BRe5nJpiLdHPacYf6BQObxLbrOmfUmKnReXKPrOydiux92fnWyP
6X+D/X1alVs8H3eoc9iJws59CSGnlmc/A54YDPwnSJLO2KftxTHBH37gtxhtNx4R
hk3zaacs3CghB4bqH/ZOcQfbPQzP32VdlmytJD4x/iGox55WF+QIhyYkano/sFKG
iQCVCBKD0M+Md1p5+qVA+nwd5sPVGXlAI7T3injz0uWR8QCHTl1PgLFwXDT7H+wu
VmNC020vp1ChASVcnLJjfGuaUb55kjsnD0P1/J1jnm4DHZEapTKB6YA8nG0kGz/e
2jb7SRxhfNqVyrhBlGZ9aI9PxnWMrIvAr6cdvYIxkcd9FOpLEUW+5VQV+gfAFQkr
zeaF5pB+O6iaxR2NtJsaZsecKvu+rNjMoT4OPf060+BCrNvAh990k004mBdnactG
t7P2e0OurSI7cuproYhien1RKwLbaqx+ONmmCHi2eUxA0Jlra/31jqJBjYQFJ6L7
H/XalH0H6qQMi0MQ46BFxHURRGsXy03mXhbl9/2necDoz0h8VF6jVjUdMlPU3DuA
+IKMpfhnCBOXUxVGRMdrS/4j+OtuwDuJU8AjZ16UlEsl1iqJqK8IbznA+bsa+vBL
EBkFniwEaMYtEqB8o6TzBGT/06mAY0UyYso7vKFjhfaA/ToUY1bU/i0m9onq/7rb
m7WCiPDJuyVFLu5bI+6c0NyV2yxItTbVyS8MVahw2B/mEfBtEule7io6cV8sDS2R
zpGQxxPjbA6NxBynh8q16fRkd6+b5OE+ua0uceoI3aIudIoUjN1H4hPolM9UX5xu
XTpR3AUupXB+3rWO0KJhKnOpD11nUjR7gEdWIEb6lMdGCnfvDlM8b7Sepq2ZynnV
K2v3+Ja0XRXC1Dq7UnLQW3Sq1YUXZRFy/Kv+azCu52FMHHzLPEESOv0ommHFrGxF
QI5l8bCpmX9YfjOi2NsfsAEkvW7Vj9RgqF9h+gcZSkrAifxrI0RyhipuArX82JvF
mZgo7FG4tiH22Km5QTnmIGoo32LH1VjKzGtZQ+75Kl1/XXnXkqpEVNJIKoYT+vfL
LCXVehyBUa+2qO4jKwL0TQf8F0we7itFriZJ6twgUyTn0zXeiKUE/w5mwvWQ02jK
OAbmdzIG7Gdo/p85g0LSBcHewgwNUc99ew3l7YPIBXoZMa97rmMMzyPnradJc5I1
AmwkpNWoMg3FUqoUyT7CjLLwEeXYDTj3N8YzWz9EMvEsGHlDwa9XHrfP9gl0mnJJ
BhtYMyvA1n4I4wz/oyEPiEB0Pygi2taD6zjpWt5GXgSlLok6PbMZK/YpyKWpli17
1mpk8cTX3CXmVO6XRaWUqAIrZPU4Ac22tQ7JRb5Vgbuq5vhb0tK0CDhrqtrkT1Zz
tY9DdL5/YnAVOVKCApY3NiWCeBqT0iHoCTizX7kkCkoJCHQXeoOfR0DYFcPSb3P5
8Wg/1xdBuHnMvkFG21M2h5qZ3v00Y7WaT33V59P6Q0cuHrTsYgl3Jtjp4+WM/nUG
MeLRsED0hoEPUegDpQvjcw63nAL5S0LUV1hsY9ONj/K0OVWKSIt5MX6ynH/tn/iI
jV5FSj+KiO0y8ZxDlbOrlHq2SRRef4XwX5a6zgftFRZLRyYWZOItsb2Q299JD/Yx
gdVDXxxlih4x421HllC7wGHSQA2j+xodcN6kYz+RvnRi2frnDRhmXRKE1PrcJoBD
tVdqqfpGnBecoNALXdKJuX3dMgBqTJ4NPtnunJI032cd59hEn27Yeja5C+XEnjHg
4v1XAtpy1y/bHn7K02dvWxYG+83nLcEadHoIj9hoy0qePtpq31Fr12Lnd6rS1gbD
AOhYePKEhTU0xdH6IJ4GwAAyNAgprK1qWRVRr/AdNGDbVpCKsnyIq2JKk6oIoGnZ
Bz3vFf1NZL3caWd9aa4+UINM3b7uUeq0bxAz0jqRnkB5/9XcpUOsVnqfGitPXDI+
B2yy3f5kgwq9lyNozhJ27hDm/nGneuo5+VA5w24L86r9n8sTmX9SlkauAgCfDPtI
2EQLJkb6xhP4iBwYkoWXxtGxSxD4tt1/S2dlBW5qfQXMd3cZO8A+BuCcKE4lBXkq
VbP64N+yyqX9B8CXgnQnbqI7RdtEU4RStpSwwTwhxY/drwEPTQfVXoxY62QobCTt
4/sunLQ3h4EYehf9PlXYcpEmbLcRQL0PjfHqHo9uwt95pLefR5pzQyBkmZDK+mYX
9P93pa+XGOsDr7p1e6lc3efdN54/5URHZpop5fWk9ySXHEeXIK/qkudrlD4lmX6e
YXqL0ZpXnP6+YTCYshLw3y9Pf2M7yfmInp1+lJ3YIxpRKI5ha0ClhaOhz3spgF1w
WQD2uARQKlYuyWwR6Qqyc7ueoIDt95ev5nZqBpGjZTmmmE+ZRNqn5K/BB+L61ZqX
6U7FiWhhaPlI06PBQ4P4P6SGEynMtudNdxm9/j9s30MaWU/VCOdQk5tPVLeuXIhu
GhUztTE1pQSGGQAOZEVKbDFCbP8MQzTZMWtA/3B7sGJkr90Y7Anoa5XI2F4Legc2
MBL2uUUygJlOXmS+5KaotYrKNRneRxpc79eGX2NS7zVHOhfRZ7AriJIUZElz3ABk
yqtjOcfKjBMMcxRSAua6O5yPnfAVQR3KM6b1FwkBJ9PEij5hZASu2tOwXQsKNsxu
eac218bTuRAuF/SzyK/U5KW8ddHHbWMNIiGQW/5OJg2fIVQ4BogQn48hPT+swOWj
aaRqRl9V74jgnsmGHxKR6bQdRrkgZVfJ+d3J6TaMenBQ75paOBFeIK8cT6VIVjEY
jpXkOu+LJKNsGR3BNcxh7dSGCRKa7xbXJw7ducxoG9zwCubzRWx0HOXTAPeiCyKx
QjMzXwkqf9Qlwz7RYK+gn3+DxT0XYrwefyqlGdFTL/T1rDc0H3uLpSow1KNaCAKT
X+rHFnswHeRgrnWB+p4/KbNwT07AbpBvKQM7cgZd+XjZvegX2Z5tDBfR3mUDpv7n
1OEz4btEEA7lmx3eFvnYb4lD3VkgLftMfEFZJx7VjDcDRjXbtd5FBos0WoQhp4ge
0bnTLfQCo8nJosBIxAUHkdgzfT5tf0XKxVG1tbErW1h3W01JqeTHK1ljz9gu4uxg
KDa+vM1GTLiv9QO+dn0RnGJrdUVTU8Mnhwz/UOu1Mh0Deg7cIJtcFcGGjRwZTu7M
Rhe8LSwUhLP6Rsd0ZAuBnUxe7b9MAKputHPcbvWhWyn7h7K1oTa6nAOrDOemE58Z
eNfLUAapZsabIkL4pPtUHeU2M4AVv5XLrstl1SaRBmaH6uCuI57QdEHYkqaNASRz
qZHSyjt+mcoLGsjlNiuLHFjkAVROd50YtjIwKEAMNDFjwYQRYpEyMNswNWb0Zjf9
PiEjyCcjlOF31L0Ah09uhgV5peIYwFrpfxd7biM+j5XjTe+Yrlcxrgd8yLWmk5Nc
VVVWYI5Z24/BDOtA6GY6NygxDbNFSjSEqL/DCc0U3fLTeQ4UjbSnB0WWwfY49tbe
0h90AOEL76OJz3jCt0/t54eBvA/m95WiAfyiE/NB5qHH5o3vfNWCd/E6/8ERu4MS
Ytvd8WKD16ADwJfC5m1z7H/jYAtYNVWbG7SYmKRUX8HoSkpTtk2oHDKoQrKiva0I
zdNrwcVRbgzqxtal2hLJPgtS297Gv8tgfDFLP0csGBjYeMDrOQw54lJ85nRyI4H9
4hhj1e4CSdhYxg20zDV7FUs1B/JfdBlKEoOcxyBd1+gyYf0EX9ezMZYfvFHmILoU
H9XQg10zG/5IPTYErMlln0tTBfhjAl615Qnj0g4hoSN1pBC3fuLcUTNUFEOHkk4o
5+WVDTffkmUDtignHJk0edwIrAgE65tTklR0qLwK2YzPMI/sLqfup6/ZYr8+XqwT
rrLEhJdiZ8FUEe5ts0j79chYc3TQZh+f59AZ4VtvomDAWhJz0ceEScLY9oUWOxhi
x9IwnFB+uk+flqpfwEpqXfvdhimzdt31rOObfFJo5ymKEq6BwiY2s5jwSUzetZ9c
sA7olZ68CexOWUAYQu9zyLCbZlK+RxWF47rbLCOkZqhP4lBfzv+5zYF55NXEaIjE
ZuWaIBVSy08qRaeuIsFvnjvB3FQYEbMibVSnIIhBN6B60k65SvHrshvOTh0mfiBx
ABVGtzCXgWEu7qrk0ef6Nx8lES9jWHpcH6h7z3mXeayFb5Qed+2nJvjCQdXi4qEx
h3JKC17zFhEJF9O9yrCmDQyl0G7r40u3lt2Vz+rfeRBGG2g6F4HeZ3o/rn7qZ9Oa
s+Ektlh499qJcjBLJKOHZ41oHFrlc7/k7ezvQ4fodcOgfgqA4g3jfmL+mqnww063
oLGhJZToV1FOTxgAXVvmWOj5sqGw6ZY/ZZ225UZTp5/R/78935E9mFXMP/FUoanI
h8ket65Iv0V07M8h4mEDuXaL6Kh4QdfGnLEYe4KxuK1gN3UGynqyqNAqkOoOV7J1
0ped4Tgb/nKCoPaliHGx+6DZLsIsyxtsY1apx1LHCK+f/dT6hc/UW4+xkiimwLhD
L+ngkfdFxlXzOqAQN4cXl2v/ESBgPXegblbuzlCIOqS9leREM/Yp4HedRjmO7YIK
qg7cUBNMRRmkd/SpFABs6uczt8pjHOFcZgw4ZpfCfc9a//+6mZlzp6qZJSY59lUU
Czphbc0WDMeVLfb40ePwEU7u3PGky8IiQ1IAPzxyqWv7NNfn9Cg1ogDXFZslaUyg
YyoEyuVMiumUmDhk8hmtaWCmSpcR3gdxesQFk67mFCiuUA7RjFPCcj/BPak3fjs4
TEGMzh0vVPIaLPH7CJZQr/JdM2hMts9WY1I0hsmchrQ/nRYtt0ClF/azt5FkVXn2
hZaTx8pAhmhTA1Grh5ykGpiCSCdY03a0NoPnzFm2uhoP5jvebNKzUUltrOgez3Ju
IGxsOkFKuCHw5jtVkSHS3VrS9MITRq+hw77CwtBxUftGBfU8bgO6KMHesFIWmH2l
qz682IvUkKPhqTQjwjFU8SlWaUUcOpGv0r7+R72taBgN3pPKKbYAk/XVFZImU798
LPKc5dHvj1jnvXDCdXIylParGWbUC1r46hWQi3flhoP363uQQLDebjUFtNivzCs9
BObpMlNgf1JfC0hdOHPfElYq3JXV8tPrGCNg9adnjxdsSRB/D3rpVVomf2pcNp7C
dDZZzeEGjh7UlGiNcegEoRf0MuBtN+qy+eGweSjyRWBw1X9LDODYyJKwtT3/UisB
eCZLKmO3oLrmQqDQRpbd6qDUdDb6pK+VLNCfwue5ixuBvSUtkt/smNu0BVxhITdc
ae+rVfPdH9BQryynn4+g1SOz53SJseeOLqVxH6qbSZihhn8XJ4DMRjC+ABaEqRVw
osj0LGhPze1WY+Vi3bsvRP9RZNv4+FhpBU/Y7iveddloYWJcDFZwynI07VIu35gf
C7c3t54f2G7zyL98mtwKQRpR4Tr23LiBg8H/8O436Ob/9icQfuHNVI7X34dFyGYQ
d5cm1Hr0TTI3sac9fZlrOk6CEN+Urjaq9Ra+FwlVCC4a+djVbavdsebIYtZmw1Ia
+lE/d77ku87I15scQBBMDtxt+W6DEiEsz4OU7R8AIGKjhOmfXGpTbLfpJccp1sZj
8kRvLsVswvn+FColHPMxgnqGpghbvQW4lzHfhCGaH18+FvpxJC0JLEVBdpWE5U4F
wY1R5dAgYH0wN75alkdXvG1OoRsG++Tm3GBOSeDVFUyeAopMibaULROorGnrZmQB
IRyAWoEaEmLPWAugowenfIYBG6dRK3dBSMcIsjbnAkrVfMTiM1OsZNpI+l4YMogS
iLS/mDu96ELugFpzyBCdbl+XKHKwogVvrfESYlC2ivVSgqHqGuW+dGqJUkJNtKD7
cGC4T6PsGkH+BkwgHEbTjtqqG37zs8/nUPUIzO3G3Zikn+baYEyolme3nKCNehzd
/4/7LKAyCJzmEIxGhecnYmd/3gnvUpOo0WqD71A8u23FIykT669vlV0R2kva14EI
oBrniUD5kQGr2syiFuvbsvL21eFmhC8L35TNNiaV1txVPzdHtWVtLpbnLhQTSsjC
4vq/klIG41MxMWuQnm9X0xq52hLaIexmCG0hgnSUb3pn/LT9yNN8wsuJuAsAQG08
GZS0pur2nvmh9vncOFRsf8jPT4DLUxlhjKJ0Ot+WVt9NFKaDhEf+0K68rW+JJ7lo
vOv5XB0tHyCD5Aw5hTHJ+TIEvpg8WCcNGQh9qrEOlDOd4y6T9N7MN9xxng3Nym+l
7+rf5SZWmo83gHTCRBf2ToJi+6VzhQSJNLdX2N4jOTpEjvt5+W3c5nF+W2ZFd9xd
CbagF/gDcAYP1ekW/aAujSDHwP7gEdpEroRxz/uBq6Po9/1ns4IjD9L0WwMjnOAH
uxC/IRmUkUiSZH7/n6VY9Ddbs7xhCyspJZG4FSrYyUPIr8a/Hk/SrP2dls72zvB5
VSFiSIGbu4eS2wuBZtn9gQ6ZMvjbmT/XVLGMh7KaPFYZb8TGVorMzPXstVymZGB6
UgvQySE8wo+rtrd3CiO0rL7BqadGJ7PnSdxGInvksv7L8TKuv41eEbO73iEZXH4b
/T6+LgpAN4yX4xz8VCe6t6I4zhTL0k9HCA+99yQpBg/A2CnzbadyYUYyRGUH3qu3
znpuOr7jmVdcxR0eqJlTeRdmZFAuUd5vs+ASlL1cuiJLSA5dU072qZplUoY5JOSY
7062SF5QX4ysMGmbFRvjtYEDVzjbfS+nhNil2qYjAZcNJQgoS0vLXWngbVXfXdRT
KqBU1+fCLeoW3zA2hi8+ja2ID8YeEzPr6QDztvpmfcezTXHM3WTVov+w906VExCn
7gj0bCk3eXp5vUMqGIlKy5X2pZ1BnKcp00fOT0eaXZNhLJM/qpUS77eZhRv0iD6M
AiLE/4Z3b5TOm5pnQakx1pxlQna56VXUYStuURRBR4R9Jz6RcP0S3aKFVA0r5Irh
2wA3W0fumnm3+dPnZ95JDnYNsKZFwsvvJsuaUKfC69APYM1skngg1xFqG9DeLJ6p
QP5B5qYHUM7bwpVQbB2rBvH6RFgEIvIQeF0WCeoGvD7KX6oFUz4tbwyn6kKZbbp0
kc1potE8c10QHLmnnN9JVY87lIIQzJ1M1mJ9Cko6NdLhiIJRVuELy2UBRvMEaQW9
zfVXtVXUcMydszM90kzJNBILwQP+KaZlP04i1iKKeaFNI6hmkJ6CxpecVlXNrhZ0
0tBf5a/TSdaew6JbyfALcqt2sa+QwRaqvs7oFmdEVx5Z1gCoQYzDIMamtRHlB9K3
u9H+KddJOtYZIIcl2eyALI1+9oaQ0CEuuPwCAziTeP1BX/D+ZnmuIuFpw58xZ8Bn
nZPwxlNQHs4O0p+ppvletNFFV6vFXPCJ2cjKvYVDelk+CT+5YU9aQrqa+X/zwrgH
7luyLXl4oRwYK07RSl6iy9mhwInahxUMlUlTOov+IzEciZR55xYgMSwlyabWyVw4
DqorFnd0s3zRaEvce0dTulsPtbQEwFDkDiG+H1sl3pMufBBQYPqeq+/NJRFQ91/u
B8Y4OePBXdyzqBYuNn0O2zjYx8taVut+ioJEYp++H1T28fhWchQXC0e6zuWAFgxc
0TSYCkjDRNw0EfcScdYMX28Ka0sWnhqp1mKjKPheS/lkDdogoqT3Ef9tMlxZ6k9k
QttfGXcrAiSrA5YiojDCB86187Bc9O9ZHG5cwAf+wwIyGnXhnZaUUIGA+Wmv88dq
4OSYolVT09z1qGoneLLyoRlZXbdGlYTQ/49UjFjZUyHtdFIDPOcQYE1mdCP2oxwK
Ojl2xa0KKSSAxzqeKU7xHJ2ZEgfzIealtAlr2Y8JWdIVO5b2hJ99GZt0w2sTiaVs
4rB1L8Gx3FTJeBVihv/mqf4p/IMzF+OyS1Djh3dI2yj6/deLWdwX/B1r3h+6hOwm
y//HdHjNC74UWGRlbn8jKgSV9fPICpjrlndSuRYyI8YOr4Hex40PHMryHGb3oFPm
1EjNjeQcuO8zeKyXbGTPeH/+l55PPGYHdzhScvES5Fq6DJH4J4u6+LDDUnkRnQwx
nuljW4n99rrcJq3/bdTJHURjdApGh62BUR9w1I+Czkpt4M21JyWL3etXOO7MqPgE
9bSkZA/4TxcV3kVGk61hdQDvyHHJE9n6l9tHeWdc5z05CYynw6xrnnA/MxgZaL1Y
7mzUA2ZnnJZb/cXGbYr864ToPfXYt2TjAsa22vf7sgsWSNBc5FsV00Ll81If54z3
sLYAq/i0+aLgrf0ghbzI1rPvN5vGL8DRr/r5xDJaqVU3qyUZO1flf4m2/AjMw7KX
aifnUz2+hdYyT+X+LsFQmavvgInmkmazEASduACRcoHbjSf5Ix0vw5Xz6jfOEVg1
WWrOPUjDPH5ZsbtMee2jeayNAw7H1dQ9r6FCMSArp4W3C8uctpOD3SEXuhRpIkH8
bSdR+Fik2cjuMwwz3JE4H1PtGmdLTCoy/Z4ZnpHb/UocS01i7G2JJeJv6NtBtwy3
r9AAIthSalqX0tOgJ8uv6H4NClyAp7gVENTaDSmulrOln080Wm4MPDDSW75ZT5eL
dWMqKwMq8nHRrl7ph+5TBoMx1NKgvyRDOFKgk7jOT92uYiPm+lPPeBLDqrYOd81x
BLqlMqfyPn/PJ0hWYJ80mt2mjUY0R6FpiESwpdh/WttSzXtjirSjbgEbsdZj3Ewf
U2FscM7Ix95TgyI4jlIU4dM60SRGgYIQ/DXmw15SqGvWB7JVX7s6HNhJYLzxGvEV
1AD9tdRg+sr/cHeU9ZmsbHeVMExDxZ22vqpy0GgNi7g5paWqlQIP4etmKCnl1uwW
q4EF1TLhsBgKzxTi76v+lGhkvj1uO2ylQ0mFu/kNTTWkR6zBoDRgWzQTGbIW74Ch
YFkZnz1TKLvgtM5K3t2OCfPCpclsBoNz6I+z4j/VqExxkZZ/4rp8uC//GBZOUpST
WV2Hoqx/glkKRtVwWiem1FxnoVbVe/Kqua9aWTJY/CKyL/3tkIlEIJYAnG6LRQS8
GSkZVeuXOqjO2Bg50TMnisV3FWY2KYuptMgOONB82qY0s4JY/XT0INJZxIvybHum
Xo3vh3kRDnT7X1DZyLEIgLWhF5wrpOxYQm89XrDcur+fkd2pOYT/7iTZfmFeFjKA
LOtxAQIzxNdvFQwAIUveDkb4ZA6LXpxwkyNez6+Uywls90MqlIvZVe7IytLt5nno
p+M3W+GABTLD1lClrAwaNJml0ubBJNNBDJng4uXNluiNW6dt9UfyeeTn9WtTnpaY
NtQWesNuiB0MoSkYJILgtOMuD+c/fvqqrr/CswyDdnWuMncDLM1ZutIg+vyDDLwr
k9g25gfHs/6LXNial8DZHBgiqB3BkfAVUB7nJSfPXS62uFu2qk9oz470d05mka9d
Uem+QwTgqGmCsLWNyqnod/ndU5e826w65uJnJVQ2PtpMs2HBGyHPoYxlFoQy3cdC
W26frTV4AxS+w5fLB3Yb5a1hkKAOpi+6gQ1CWQUgy5QLdoTWIZs7aNcc3x6J7ZQJ
JAlfyJnpn1I666rPrTwX1nrJ1pQkReU+P2NrYHRg4RgCKwduoFZAMSP092DveH0y
heDjssWgJAUK6tLCcGPYL6AFbuLW6jasLRDzDSS+C5vayce5liXA1O+UNEO7F3Ia
ZR8sOhMWS39fhvZsgjwLXY8najW+9kC0ItGbPIDPijKCdCo16USZhNs6wc0DcwOh
q8TwAIlFZVAyzJt39Xr5YIui866lI19YE6X2rBVnfY1EZX5654S7Pd6tQMvu5n6O
apXWniVeQwVGKLmp6ZMduIDq+M1P4lXoDeRRz407HerEb9rcipCAxqcNA/ozgBy2
6ZBmbTVa++i8uV6OhqA+eKWiWKtGpvhVnIlWdTj1Qcv3W6XqMnAtuJum5vWHcZjT
yeF2YY2aYfmA8bCdqBUjvjvVifUIr+tkGlg6qKAfOLyvFbyyouvn4k0yMX3GSZ9P
bR/s8T8NO21sIsfJY9Hho10uW/QcYnHXPhSaZc6XReqIskk8Gmv+xawVC+PM03S2
Jkzy+R5lxkjN/ZAqDVXzSdpchHmohpWzH100FJ8Uk4sFFWGehKu7qpG3rjPvRqKM
hQiikFdrO7T4tn67CKW17fxoaYS7TLAvWf4QOSivsXvz8cqDqhvmWJI53Phnliix
00gpLs35CAu7Atbk2QTQLR09/+H+KZAY2Do2ZBueGAKygsbRS2Y7pOmf2IUYSedj
AWGuIDJ63h451MEp5oTFkum+r/SZkXNaveblkKev4UDQPt/RgYamUro5FBrmmoNl
vQ/7W09kXPFpdxgijca3XSOLzxaz48MS64lgEVjVsnC7wt6qUTls1p8zgn2NCPul
DrztO6ju5gvATiZ2BPrTVpuuaFzOftzzMgHtudij8YCDsPy3fCVj+msApSEAPSRh
CBWJm7JAR72vH2DQbZgjssk59XIuoLDtJkegNcT+J7Dwab8v/pzvn3q/v4fUKIpy
M1iu3h99YSnSZSSJUiHlEtsMB9Ri1tDeGxcE5iOlHouZ6BVsnEnwuVyiTy03zuZa
EKeltvjmJOnVoI6fB/CDk4jYVjBinQrQc1SZHVV7SjJrPFDLNKChjhuprKKvdbbt
RP/K/FktfEyHxs+9dMvQByoCa8VDBFlDB8Ncib1IVtE4JozHepHh79mKsk2MUWul
G9Wcub0nKDEqfmYKQfkuVjNyqdzIzSxOGiK2V3dbGzejSyQlDVgXrE6xO7HZhxIu
iO7905qoSXnFiZpimWDZwOX+guZNNgfrLDxVCX5FClYdNnGE3JSz4NCDUhiB1ORu
t5ayyhqV440H4JXYNv+25E04666UB4sZIfne7JYZGxMvRiGy06wZ64+EdJvT1+Qz
O2fu1MVmzc6livcPTJ8+trxch7wVELHDnT3xPSW0GmT/j4tKRjSr8wiMmeOh2Qd0
5QLHYRtQguxyrOPak3w7U/Z2Vhj8Jwo1CkylvTOm436D0vtWfdisqlVDOorAaU0V
Nll7HVTyVnJVotwWVg2qiy6hksM7HzrFTz+Dilr4nmBlYfmcWPpM/9fEoVhxRNds
V80R6dn17pooWWY4zQzHJTR7/yeSiklePRk2Ozx3g3sexKPFn5m8qAN9qV6Xij+w
rWMYwYeph8eXgXgEbSAFCT0JVJa9KSaKePa2OV4UAS45BDIcNroqJR50wWBsA2Uv
xtDKqQh4k1WF/IGmAUB0PTGOL2ZPWBHi0i+wZdl7mmLO2lmvhf9VzpAF6MI6ZQVY
5V9kiW/y4vOZVw0mDWMsHOI+aTww0HSQMJfgrUGgRsAPa8Lyw2jGG4GurSZWDsrT
djLFVLzb/aLGRUqkrcnB5Ts3EkqUrC+6BKbkqOx01uIS7wtGtQmrWU7Pt+ImfLkr
sbijYXZueBdSe5EDgwo7uuAypAEIq+s+uAzGVOlSwXa2VoYdSzJcOjYzh+YPsPuY
jJ3/qJo5a+Yk9k7BeWub5rWpaJBEnTsbYmvmVIsE6VUx1TAuVVYh3wwzSbdx2cJp
UAtnQAomZyIhN7jemMJ97PUOroRaPLFESGAV3HnyNOBy3mqgOABnozsRdbLY/FD7
m1X8Y2ayT/9MrM85ur7EeNBjyIRFDigpUHd8ShSzlV7mQ7gtLavk7OWgHxNxkEnj
//sVhDGRugHkmyRtPlnlVbB48RkOl6ciFPZeEtrDx7TL4EPGTpfIZEDhN9c+SnLO
HE7oUIqFxS+RI2dIx4fCFpxzVnapAt3r8vAa3Pgrsc8NKPsYq69YNtVurSh5qCV6
hnzpu4+QD0YbKtmKO/vGnvNXJAnltgf3QHRsQzuyFTkfu5IKXA0wMV7Ydzh9ltFy
o4NczbNTAvfdC/TSXh7xmeQGtfFZKqlIJkpSBnVIzZJI2vcKgWmZguqqkCpE4CNi
a5yBwv7xvAW+RCFxo3uqCqEMiPE9R7oCCcMS/pzF9rtOx1n8pOaJSEU6XfiR94YO
ieK35zvuel9FLjyfEekS41QMxU2jRIsBLo1/6zvjTRg++pqnUHJE7DPQHZA29NZx
Mird7G+qJ4SSRX8lcGgcHbcFIKmaYEO1887AP3IR4ZDoLlFW8RVsk00P0nKzlOsr
PbwbY9NZreuRhcIJlrbXwyVoyqXiT5qnIP2ijbMGl2qCCZtksFqKKlJUGHCU5iNe
mj1uURVKXsDoFoApb5Bp9jBvzVdlwn61fjGVERquxhvehz0Q5/46mAZeZvmN+XDN
y40uMychWokZ2sJ3pngjptfXzs+rSAkhhem/kUDWIfBpmz8X5BGe7GVdTcxYyUnc
p26ccZN65ZuNSWIAAe5pvi9JQCmicud088egDAzXnboj6SqlcQlQUuZRRWscFom2
EhS5LwPghddTkV+UJbGHxH8byttja/FS9VD/Sb/6DzSUxdJ6ncy7AC3K6pzW94sG
bIMaJdVhvJH7FGXnLjXJUAwyYUxH0GYSBEvb+QBGWQYss5GX2heGnSMPuK65nUsj
sZF4y+QkMQdT3pM0XGADHrI3W105cHUoc4jdH0nK5lNPh614E1tO71RBkQnf+4h+
YY//LpU/nHCVR7fgK6Ft32dk4Tq002vn7gW26d59Dxgeq2ntY/RO1iiBFQxistek
WRB1pH0BFuoPhZI5OzujFiVTE3p/AvUfZB8xxtUnMfp6XZsET7T0smnocznDqmh5
pvmI18yJQDh9C4KavR1v7CjeXW6wUkcPNIsAiliTJOnLEXuXHOfQlyrQjfSbYD8M
nSpQmxjlQrKHJwff2CKHZhm/B4XvaF/UZW0WdJbF8E534noqvtgLhg0zbcx2IBP+
bsZIPbkS+QJJYp6kX/1y4gUhHZy5DWmC4nXnc10y8kwyhnR3Y0CgmCp18xOhCOik
qUVqOeCnQtWFZx26U41YgqbrI94fktKg0elJ3ewneQzkO4ALK1XTnf5LCaCgTLA3
UdAzg+okGapFw9o2RnCUmW9s3pW2f7/ixpB+zRZ7dB7CEmhUxzxTGb/nxKBtiM4x
nrZ2S0cz8EFSzcY+RxhwjqB7nFjfdLllrTpNxQ/Xwr+GwDFtI0AHYUBD+fWF03AA
OLkVqh0YZlIPJTTPY0mkAXcK/1+tU2R/GJUZNEzvHHXtsqaW+cIKzKfuHQO4y3AU
Kmg1WGDWSLgCqk+ZPHeJ7SsSMvn9qvC5nyDusnA3IU8xuUGDBpEf6dzxkgA6Ohuj
+qHGg0GhVtz+6Y6M4SRwgPBfy4DrcA4/w1pcDk3W2HCjAXY0mYbdrAUoHFTs2TgO
xDb/IXHqCuxuNIGX+Ojd/36UShMESYPCb9WoHe+X6P5FXJZyJPgBH/9LK8wo35+w
eyoYuIWDykZIH09aYMOVfInZT63s2MW3TGbOTpnEd013295FI+mqA+ZXX1xEkaai
T7uPN4BLa3Xy5ezVJLBRNw/UbxUblEnQNQm4ZfThJ/h+cQSjkTINR7ACs7dfloX7
BuWgGGxOtjDRhLvp0qgwmHb6oKBE7Hc3LlBZDvE274uetIcmwYkrqclIkuVbvZge
DEgz4uhXTFr212KEIJ4ehRC9uAriPoxBprNqPlPBKxFWY3w9dQE8ldTO8wfZXZMa
6z3BpY7doATIEbx5F0aJdklgd8EwcLShT7/aThagwv/+UzF3PbKVpcGpab5F1m8c
odXsmJnBuhoFrzJw1rOzG959JMOpd745rtryAFS637ubiWTTKdJfTa790cdyM/Q4
sSq+77HCGOET+hDemD0YvzdVKYc05QhDK8DrsqjBOFi1Bn9AugaDcL/VZLVkJXsz
eFGQoHqjGYWqzl61hLHwaDu4Uh5Nx7EWLF7deaqiHZfFXq7We5qrend6F0SJCu8f
kF1JBm/245qqoPIEAFrJR20nLB4IP/ZxKURIIa8irg9FypvvR4Rc4Jzpp6j2VnVG
6a55pvBgK4CYNjZ6dKEVVsogMManKDKRS1t7gbdHp0BQUpeh3dZcinl3CXFXcEQs
WPJnwe7cB5yOvDsN/L9syWu9e+eg5d43asUQzcGV1YCCDtaPJVHfeF78jqR9w5lp
aGhUe6ERs1zNbyDta34tr1kp0UHR77Oa68rxeaUUsnZgJv+qmg66rRs6iwSp+k33
ebekNTOGsZRNCWMMJSrw7FAYdk6kde+Y5ZWAmHpMXW9etyQ0EUC+cMVZMH6RGYL9
NPaiO+iKd7ZqUG/4rknvHqcY0gZOsmpYPZ5ytKePzK59yOxYeWR+vyePkEDfMRPi
QGRdyP0o/8mtXhAkZwc5QoCt2IZWSqYfvW+NNY+SEeLKJUNv6+kU1mEcH4dt4XfL
1OmwB+R/Ckihj2BVvN/N4xuhDPnfVjHBb/kKfAncJUR6UEclKVY5zFAvSdkESEwv
EL7FOtJZLtDGjzxfXAkamilVmCKqHBjGKKbsVeAnh5fsqGdXxRYfvsZ5ls1i1ipw
nTHw4qwXnvBJjEmhZJnQ1aWpMAmKpM+o3Jq12mLHVK/zgm23NdIX9l7tuyoqNsze
DUxrk3f7bBJI4IfHHku4pqcKRfLjkZS42pTD3wQ2A40HWImQUc1qwK6aIkxOpJAk
yqBQCob52V4H2OWFOiZNR3vgcC3TiNd/+QP+fEjeRpy0z9UXYhHnzdjpRm5tB0Hz
1XQcpFqubafYkSpCkm1k4wNMopEiGjDSkK6dqcPL20kWpaEOMOL93e+u9sp2L7Dn
I0/c5XwEn98yndA55MxNTLYL7XJ3xPOGJsS9fKn1h3/NU8a3rvtip9ucWm++jD7p
Se39NezhAJgqFOih3NeMRrVxoYRtOifZFV0YmZaF0Mqr7FUi9W7fWcyIwTolrDfC
xsc7YGm/RvtSf2j18cl6nosBq1pFAZCqFdrpq3+5FRKfzYtMZRgnHgsAHNZddsha
mijfjdzlQxPnAGPpV1ADL0/i5z3NG0NX9G7TJjIiNW5lOsJa1FsSYJ+gGPze+qLw
g19b6ZYK8g0yETATiSQSmx6Ivtkkl3mzo7kjlsT2rcKrqZTQHLLqfilwWJ7oNV45
YLUqmhfWAtIWZ+Y2/qI2Vzr+5b8UGcU/ImC3YLGAUcrILFv7spzlYQxm1bMRlT+V
SpIgeVhGmp+ZWLMxklMRwMOtNZQ7AzaSZWQi6ppSTFXLO6MNTxbA7OXPaJQRkXve
tv8gmvQSukm71YjGmvaw1tHUpETaPihB1Ka3gHU8QP0qRs4k0+HC7fGsKASjiXht
aKrU+ghZ5nezGRy7VM9JEIBzVZbVuc9Ib1W+jzvHk6YTbVcVVZoLZ8hWCczkO4Bz
DBZ6N+8fTeZozVMseaVuyh/jawxrM/kYtLDEMvTy9Beg0beqcAMjtpzk92WRIPVt
JpSl8rcA/t4taeA6Ixuf5FSufFbGwedA7wuyq++HXsB71hTGroSte+GHHvLrjabX
9x/H8h/f8lHrUx7n0GCvjAjf0Tqh4DrlhxFR5COutpELMNLk2REV6aEWUjFEmtS0
VCtHSlyFS885583Q8d2HQsSt5hMgecRpW380Pwz24L1F2HTOVt7EuI2QXut6enKN
isAUBKKTY7QvKr+CiVN22wPoUxHRPjxDhoMgP2Bkws5EJiYqXyrIqmxzyypQlbq6
btFx970oeBoRQRmGowWwSHi110G5vJqZsoq9dwjFYCH8+6fIT52CwnSzjjh9w4Mu
K1xbv3FJUCXc9cgLSagCZY8H+o8RKqRp7AxiU076djH6koQuedY0FzrRvvzq/epm
UEViHY2Wvl8Ucxa5YfvSB3ACxd8VT0QCBxWj/GJ1wq9zwRzpX7oXjlkqhHKd4ODx
y5RT8saFDPAhNByFRW+MGT2Umg8kSI9ruAbaYGPH8rYqfF0BWD4eO6SP5u4EMTwx
ERFuhv7tVRfW8HIC38dnvVC3tbP0iuIPf/y04++H9Wo2r3cvh1Fzph+TIusgRt+y
rc3OQdrrimLehA+7WLf0hkkthTpJBe/slQuHZyzsmx3elYk45G8xce92hzX4817V
yUxLYQEkBnvjoERckATTD5H9zlAFmCSX9MdBAKasd1zn6RviTnxA75o8rXTHDYG3
YlvGnBszpGcqvs+fqBg2YEPj8Cjfz4lNMGX8CBjw0CAiYYPqRzN/WgWN6SYjuwvu
QOiFzvY/WuS5TcLlWyAIP8YB4uimGkjKMP4D95TVyj4sWYAmknur2jgQKAjIzhzR
hjKIs0xqZoJk1A8tmHv7rm1Bf7f1zAVXzhnp3eSC3vKK9MpNKnxj3XCXvjevswaQ
PXaoSobp55MiH7geiNb7XSNklRNt4tgFGWOlOLqrLO0jcw0E3ryJo/XliuYhdznD
N3Q0c8GshYL/Iz0t6ZvVGmf0cnA53jinCF8Y1emo05biPFCttYpAtd4Le25kebEI
shOumGMg18Mr2RaxMa9UkXHeYdWMBT7YCG8KTwBoQZmGVervJiCB7ZIVXfHrO0DJ
Cr6aq5RkN/lRtbUzbkhqxQvIrQ/5IDv2FbjGbKvM2giswInTgysVukgQOKjz+5La
PNOcNwnRDx3tq58AI2CoTwYYPueZXvDwLNOY8TwxVAw5hUcidTZg7xOO2khkzVyC
ctwe0YNEphDBOcCOjrLqNx7MmhWjLyU0Au+nT0iPa8Yu3rMaN64sVskZmgvsFmZf
afY7zw8ZaLkFzkzH2OUqWtmk+U5YVHevJRwOyWYZKTXSOYw8zxSyHRAUohsvEK7K
3827B3fOrBKk2V2XAfvWa6Z+sx3iTVBanP9dSGVcXxvVtO/7qRRlwmLekXeUwHYf
cjR4gq6UvPI6AeKUcBn2Qox/4KJGGVOlUGYTs5eDw7NnCXyAq8itcPZA8i2/x2vK
MG1tUi4+xgAd7ms2LRmtqjpB6OgUnPc5N+k6yCVlFqSp0LGIwO9AITKy6cpoYjr7
jYYBuoTttWFPLaAGXzDVK9Xf/dWPurDIFO875GJcQkyGcdFBCvWJOI27inmInvcl
V8AwhULqfTxwkBijP7EI4a+XF0bIAJWDQKck/46iBwwfBjNnHsiaRw2hqp8kKs2w
eX8Us/wwonN5ihpFfHXtDamREdFBavpXfFVR+p2BNruAP64/swNa//IhijFBt+m0
2e0CFeTUw0tduLrEQsmzYP+riHi+gFHNVc1Iuhwn/72FdBf2rtOHmJlJ7iYkefuV
gB3XGOUE+A/Ot1Oqr3CX0WfKAF97bVCEwoqkNFlWUxxuUfIOXAPKiEYxL+Kyd0a6
wiVD6OOZcHaHw5kJMfBWrnBm83zLxufO9DdHA8TYmCU3V2wIl3REqCdeWA+w8KAJ
X+8hJ9O241XX26ojhoC6wpbTd6ULlPSIOLnaNU0Bcnes8HDikL7MCWyLZIp+5MKU
SdXzdbSSxkPrPAAhw5gjwsc9OCS5DGy/2QOivKq6JJ7VnB1nPrlWYJIQ8VLw0mRz
S/mGsCrFXjqDLKSd2FS6l8wqL5SL+l/WMh8NXLC3wQSbMD+54HyA98hO9yXMjKf8
LUUiPlHOVyIVwP46APvnujaEQmwdk/1MDYzhxRI4sW0KO1NV3eAwnfgxVgreJPJ0
ux1ughw1CVCCGi/Jnx7iIDyQ+cZFCeyzNDVQmcGoHQOR35qRx1wv5hptF7eY3kpC
J28j3n376V9aHC+ZGSJhafjklhG6+o7tYXukWMVLJsj30c7NAZVYAqWHAcTeymLm
mtyCpmClMjZtdmkPQT6Q8saMK3nFu//WxfwD1olKuaV8AkKz4PB/VPqm+QhiJil8
D/W63u6ZtseGjqHttxn5hoVWDAZQgEfDn91wgyX3uJalLKCDZm2GguWP+mLL9wTl
ELnWBdwo0ysiSznZtbsmBO3O2k/ma73diZdpfqrKIlHx7PyimkgKkYIOfwNKdb+n
VBQWlzuLxGoRprnIh9AeAicLL9IjeAc0YXJ1rDeqfr4EiceB0xsqz9k0+H2aIUEh
dlCMXZS83Q2s3Rw3cHfUrCXQCoZM9MTprlD7CfEzKFg30oLYMx0ZBg3j+3xjKrYo
5SwssHk+DE/0uD+fD8UFG188Wukki1s0zoxQCmGoPW8PIWfyU3qDJdgudc4kFiDk
5ayc7U2C64wn7xoQj/VHSaluW+Kj35EqHGcONWCpcOHnJs1ShEjq6s8V/hrzbVBZ
V+VECFR/E8cxfKT/JC1flPPDJ3fuRMX/WrWmteEu14jW7NqYrGcjPiFnHG6XW+Xd
HZT3luQ9hGOLBAmIAVY1byHX2KDA3usAncARS4j95TeuxbtTUyfPwqXS7Gyq4m/x
z9mImm/7x8jUZOn3RhPFn7hsE896e83eOnU2gwU+10y9c2bh2PdLyJb4/EnTz/u4
+YilzjxId0wCMFWFZbbhubdUoFZaDEeBt3rBSYrqej+z8RJmO13TnOj2uSmJdCLt
ja0LjXsgTU51oXq0DA+E8h/Lr9FDL5eNxIyhNMlvTfN2c/gbqb4LYE8t3wT0jai+
CzIIj4nDDXQZzJWlQufxHj81OeiJsyh/nE46cphbaa/VN3J25G2AbCK9jNttpOa8
UzlkbDKGxj6l0aGVegkW28T/HB4IyTI+2wNvnBVw7hPMpxLBH4uf9wc16Q15zUW0
V0TYspFEEH+PaOeuEmXZqrIfixeUkaOxKRsN8fXhe3OREFvUkCoLiGMsSsKYOz2p
N8tLincczVeAoojV4Sq4rl1p3vHWhRt+/UgEZBZiDeoAwqubIeTx9atHNZu6TOVD
xz/Wtx6WXHc6Hw7MXURdBAB3bHodiyWJaZY9/O/AHM+HoOcQNEKBbt3T6zTdV2wz
oMqix5moLVzGc4uyZ7IoQmo+IDEbePhS5hWsREqBHKUkvUlhUpcc2AAYTZ38UbtZ
p5BkuRUdUaNdmGv1T4uLs47eYfAXH8d7+Os5ZSJwdEpkUeGj7j9k5JTKWaooibtR
e01xXVD0H3gf4AtYGUnmUxphi0zwdub8t3rtxyVBKVLhomsBiNzmHJ8JxDdH/wHE
ogIcZjtCUQTDP7CHblq+5GE2cqwBjSKLTwas08RbHWtcEBwhij16n1FMxynuF3RH
tmR4fWQ4dncTUuPo0pIj9OYMxRH0vmlxHFOl3aZRZn6DUV/veLZVoTJ9su3eLH0r
FT2e9RGNFqFqCsK04ih+Mqw+ZpGakfa8oAw9rM22LR+dc5FovTqgriWAqm3boDuc
CLhPn/Oq9v4n0hFt6wYRarzdi/39hRhSUPxlx9ANtU6kNBTyrj82vmUoCPlj3ivp
QVsWHdZ6RHaKFjtArqcLIndOGVm72+Jn0O6Hl31Q/1/eERStwjACg2tN2Pf7VYbK
VBlHNQh/yQYbbTWxXL3dRRLfwKOOej2wE8e4R+o/c5VyCth/WOxodBSjyKWz9ZHj
r2k44+D3oJI28T0v82GzRqup3lnvcN6iyfLrJ6JkRvwp+mPOdMZFyEPz5nfNn3fE
YbMsX5GDMQFMxWs3MkAvGx9W7GathKqPbgOpUbbtr9Iz1kuV/K6N0hZNidw3hss9
yT5uqqJrSPOjvIfp1QSMNTkZ5d15I/HIT8P7mXE2g0Mar6kMTHB8v6WzwQtJ/93k
YGS1bH+R1WmPJcOQKBo2StPiNyASjOf73K+zDM2WIKzGkjL14QwrM0A3G1qZIjGe
nQg3N4NdOFw3+Mm1aA31cQSFk4ppcuDcgOzJLmq6I6wTOroxbz+kkga/NaoVNtNy
AoLAHgK5UzQviJ9R0FE4ByU6nna2j3Uw8M2SceKaWaySsdnecEi2cwGSz057C1NB
hVPYCYE6guhbK8hi8Kv1jABGPdQXlOLpD2XoRkgpoTe24LxiV9PirWpRZAdKLAAr
rsj/477vV9w4cmkusd5swI+oXHKvESjappMtxoouPUq2NRZg8kjT6OHOPwPH7hg0
z9LU+LwA96m1X6Bc91E+XSepXY4ufZm7OivoDs+dmBdvEVjEyQ0Xi8+dJjLLAc26
b5uQPVfEmwInHV+4JNW8Xe0hO2qj7ynrjjJuhquxBU8sBhwFPvoEOISqhBo6I3a1
XenFFfQ71inWfPEoRp5MT2bSd8Vd6ZNPJ7rRD6o307LmAz+WwdVocmRYvp/DWOLA
RbEQ1BuoL7RpmhXJBNI8SxtJViP+glzITRHAMARzlflbamTBXlzidIddAVEn/FGY
Vbo3yU6GeCtVzm6bk6XQ2tu+fGAPrhYu5UwiyfZskaddVRS+3YYVm9MnvhnWXHPM
QfyyIojnoZnIooogXgMUag29hT+1v9xEl9BhHW68bDgj04hPsf9GizfdbHcHi3IL
V1QbGVk9cX9FIPW5z3Ss3bQR5G17vUdQ67pIqQCEiDdHPtAiG2asUMPZCu3LHIEF
EG5XQZ/H35hJ6pAr0gcMbQZixp3XHxA8MM7M2GeTb9Z7Su3SATFYQW27pgFwNrYa
zrgof1F32Negkgrv2tcG0ohUSCdAI9JVdxoE0KxrpQ5rkLqWY1dNibALIuLZYo/b
jqWqH48CuGUXOGJJix3Bf+/j893aHE6p9Mtk6GRwA+TMNb5vZh86+6dYJL8HQi5+
2y9tG6mz3kIu7a6ioagi9Y/m29jfNgimA1BdygXxeuIyUmSjuBRFbQBlwKsYLpfr
xTMPsFrDpEq76u3AEyt3NATXlZX1AMwrW9G4H/8GKs6gmjgZjHBWcPAmFYTm9E1O
A23J5v14oXEcB10/PPy9GKzVM+MJeCfmHS9h3KAr5I/QHexD/hdrpch3Tk8u36t4
k2m5bdpPVmZjwBoIu7iozEmqwDP9EXZtI2H7oMukHsOy2YUdg0dzgDLs+wXp7tVq
LQ/LeEoxY2FNdW92ANaMb2n1vxUkgoYwGp3J1wKQmg/CT1Q0ib3MwAp+JN5krHPI
W0/D1+e55BrkhsDoKEHB36NAoUSfHALdu4DGEJKWqLqRqLH/Rf8PMtPeYImBhiAn
QvNteHB7OTzla1ApBppyUpVeAau2b+hSOztdJAYQBY5Pe9QpMpXSQ91svLCrhrih
SXkC7HCC5HbGlGUOzJOItojf0ez/arnzlL7uWMyg/DkJwGGZJaeViO58C45JrX2R
3dNULGdnpBLGHUPwcfnuBfdatT/J9gXCsYLmDGd+fFTDFpNARayimotWDM+vPYTr
g6iSFFafuv9VuXx4qYh1t2iCBI5e2e0gap25UyVOajk3cOQYMhm9XSLiKf/399Bo
Z+pO9ZDL6UfEYlm3kDwffctzkMrniz+KGHiTlLuqp+pE+4QpQbY2PJj7MfZ+x3K4
fM4pyU3o6/TbS9np3vBGN9SSr/sYubxATtLMtSMpqbtfyElW+L8eoaz+NHgtA/o0
cdOfo4hLGZNnDyNvUKNa4tC8hdyOGqo/KmCAEw8NeD8g4PzDAIi0yssHXY4P9hVQ
0G30I52UmQr1sYtkm0PX2/suo6RRdkLc/wiyL0b4GcYBiSLje12o3DVRxlpOpfIj
OXYu6MfRGUng0JYB533wBD1AA4r03rNdnXB4HeGuKqw=
`protect END_PROTECTED
