`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zycQ84gNYF3CMXn+cUpMMlGwlcwq6+1L41ewF9Tb1LqIdBsAuqQ5nA52htO9cFF4
R1vRDOgX28iooEuSWns0zW8VVAImndJV/FjvqubozkhNAhOPzQHLkTfW53sIGDQ2
BdS2EOTpvs+I2YW8Rf8A9p1A+Q9aIACM/0gDsuGHuiQo3KhqO+tb555vZ67YAnmY
vzRRQBNao/b7JP3Xh9hBfMeRYtj0zdXHe5/JE9V9hKnf7U66LH/D9B0ZtUPIGVog
N/oVIZZJQSQwK1B3LY+6lIbxzOGuYMGaS/ay6Wce//Erndl+fw2+GrXeLP9NIy5j
cMo6tOwsf7Gqf3q5BTax4tqX7YvZpKWdV9Kpj3/n2IsnOPq9qRJCOn3m3vEMOHN8
9k75XiFQwMbkmHRyV/2hhbebdaokz1H6MkQzs80YAsLbt2au//+G9jFnSlpueJCh
baLqssduHl5c4Ltk12630WRAPEuUpUsy7HzIVp54mNzcA/dvTpfZkp0ETHMdYTaI
l4pL/ggXakQe+t2XBOLgdZsPJkXRjJIvnq8shmwvEjEKeb3AlrL3cb1aTpNyIQPP
HblZWVXs8FNK+a+cbCSkx5JJBOMHdqre84NqN2qBjEIdaY8Tz6UiuR/9BIgWdKpM
QVGVpLXL+cJuz7atbWCKY5TQ6oqFvXjGNgqKshGBZUxtZa4q7WeXBJD/Rdkawa+1
N0TJ4+kedislhPBnlklIJTj/dDCny7GH7Hygu00ViDG+0eCrasA1T3a25XEKsQI6
SJofosn8ifO+qeRQlnuJeS5vYAn9gGwCjkit/Cmyk08GyWuDnEqmyXaDER1ZxE3b
GsYqmBjIQsYfeACOZj5BNQ==
`protect END_PROTECTED
