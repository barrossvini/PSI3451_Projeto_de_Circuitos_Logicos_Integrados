`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zRD4bazFxR63NyY8cKdvwNT89KTK6W1wUaI4Eto/a66IIGAgaDp4H7QdUDb/EhDd
9MvxvwnKBGoQo2rLfzFhmbTJQ2RZWNngIIyLF6ntfBvvJ4T0yws7n9hXfLrueYp8
TTbYMd1BjgfILYUtNMhP0VFdp59PAI4HzAkiE9opMH9kQh54KyVt5HjH2Sj+ykkU
Nh6DeIEbn2PwJb7R42nPCsJbNusGrEmrPO2IsInF01mea1EUVPItk80fQyBhKFL5
Vr0zFUZ9nAd+CTLbNDo7BkXYBsCfhqFul71yoKrMGQ2/Ahq95+flQxMARgDJ/O9B
LGJTAKeTiSkJfyRSLSjONHHXI6fQgFRW7J84FNQKQ+LaPyl9JcheE34DUSc1cvie
hDD2H+xTpg624xVKT6xpw/SegPcoxViDxMiKSdLpnH6C34a2KQ/xsoLwX+eIJQ1a
g1EKi9Yl4zNqmyWaP6yZH6MCnczONUV+bOFKklEAws1DtUsSkxx9MUzaCDaJe4f7
IRR0OQ+5Y0OcxJ0REaRqWweNBumlbwptmyBG3DYE5mH1NF3Vnl+0q3i0YpORpiR/
venkv05ZBCHJH0e36q3k6HEkfJrokVMFQ0Tfc+Om/oVzlCaBjxNYibzB/AyHqLnl
ZuZF9MSnrUsQjwz/9obHbBqOMeEHsFG/KNAqUS9avukNeEESIczEhGu/ENrJ4iEN
WiiXRweLgG8GAX5atWy9+jvWlaKT3vFNNyI2oGL7Ay3Oe4WzTcWhMSPkUtv9/p+Y
7R7L9B07WxSOsEeIbRW39zOaPK+AEUf6e+tyPqyIaIthznTmZB1SpOjcyER5eNwY
RzH7W9PL093GQuXP+pqq6c0De7+vn5+5/Pmsux4M75RpE+d3dEd8D1gM5bhVd+IQ
9mUifhTyeZKDvIrGDyls3b4KCtvOOog3Z6FNU/KX/HTHoBUac5DGulsLO28eY/YE
So5lOZIaEs6MOcBQgbvVCSNaWOXtUA2HELZys+uBASeZCpm/rbhVC/eN6GQGQyRc
+v7YnPn2cKPK5WPBDXJwlY87fSq3alLgmd4/5eMIp1iaNMInXW6uTY1rPXbZR4ai
hRJXwaAOxAxnjP6BfO7aPcXtsfrCoSxvwNHKIM4lSkTjsEMRSdquNAQTgLb4mutC
l1npFPFP1W0cOSHTOBN9bp44BlFm1cAqyH2Erw0tsO9d6F+Kjba2hQYcnjSiViwS
Tn4kdMjFhQoT/az0FsTwzrYblBFBtQb0pcLm7/uQ+8X1KnGDfh0cklmeM/NJAWVG
QDtSaE3vyCLDxG1Cm5gBrt5TEhZ88wcMDN8lo2auRvKGjHDaKKUaNazoZ6VGAQ/5
DFztqhAGo6+PW5JKIF5/xRQno+ojbjlMLKh0mSSOKWMkmm0h+bSGq7tXLYM+Ean5
gb8dVSRwRvsEe5zBL3ywufYQtIkVs0Q9vQPJdayaTq22c/gTPJB9wud93vjWOuPB
HKKQcRsCLSc+KUf1K4fesgUHNdEPw+U7EDAjWMvYlLrbgdp9OjPyGr9az7/IV3Mp
uWj9uwJg7smUX2ej7/7oC2CMpVfG7v/AYHKEyaJXzZdXQRQt8vgps0FaFasbSVHW
p1sP8M5xVY31zegdT0BmCkn3aQy8LRZhbCSp767fxoTj5TFuipwgCqd16hipCXFw
`protect END_PROTECTED
