`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RRgtD/rr77e37AOxYWhmDPKM4ukMmf11tyK2Alv/VjTT3H68uWZAB866r0Y9NhuX
wGJFWgUeHZkZjaj7wX7U3r6OA8JhdKRHnpTMYQZBiLcxA6X4iZzxwYpDWZh/XEim
F8PrxTpazhPb1TGV+FqaEgSn9RP3KIgk3jNVfrVP1xpyU6QkxQrJQ4o24DQf0u95
kGv4cKwkkFkSBF8a6fkjC+KNucr+zsCBewSc+gwqcI3DG6XASQRdr6mmtWvkjpBn
CFYBu+vEqCMaRnCF/DkhDsgtpCFnL/f069VeunUqkqVgcz6sg1RrljtnuOTj73JH
Phm6wwC+Xosu7QRrRwTDNJLlB+hp3SnCzrYRp6w2s5LQmItepAKl7W4S+Fx56oGl
BBUXqT+ICPo8/IQDEkBKrBkU38qWU6bfTnfi83ocbNtmP51J6t6GICIDO9qo5q4d
6/K+/F8HuvviDhMlRvodCa5PYv/CzcSM3wyZ4c2GK67QAYNKfExDeS7FdN9b4WE2
gxYLc8pEG8l0of6Nsu4KTw==
`protect END_PROTECTED
