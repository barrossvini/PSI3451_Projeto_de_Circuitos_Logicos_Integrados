`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GXcs9NRpUymwKqxAXo+aDlawGH9fymsNzqOod0cRcxGZTlITHmj/P8y9d2Z/iDXZ
Y7SacXlQwTsAP4iuj+RdtEvvK3x0PvVeFhByOHqFXizIDCYIAQtONE5BuS52uwu4
IirCweV796Dtr6/kkAXW2k5yBdXQqrANkGajVbRNa4HmSuY0J2YrKZTKd/5rPLsg
/7I+lkgl0HsOkuDnLZk1wTSdj9/1gau37dxXKQAD2BZbXDsleRfCcQI+geGDUMUK
EU5+FpeHcmOwjXDiI32phSIzaVyoFNtlWga6CLc4X0a+IsY1cYQm1wY41+DFxcGr
yTxOhZTEVIk7bl5fjALgxo723YSEUYc1QDM2UQpP7dsvHcrBrY79Yz83aX4Hcr9w
eNOSul6pPgil5tN7hsbG0eamZLyQBOX8obREGasPZiF1cu2IIYZE8RJ1axYP01NN
mojmWFsao+6/LnN6RKKLb8ncjHu2MDuCO+mk69S+cGHC5vmQlGnr2/f204X0AjF4
veXxBjNBeXnrtyf665BM2ugCdSHkqJrWz2iDIaK5LbGTE723UGpnbVaU1MIBsdVf
ensi1EjokZK/ewzaKJnTi88i9xYDHnbUPkKODLq8TSksTsPjc36M4H3aEnGcuzdT
b7i7a5sQzDeJhp1ViBVZc+KtLl2X5+PIJcdG1t5MGUHY2AzU7o8uzdEzznBdbVT6
SdPXSaipw79T+gNr8LRW2RlrTlRjvd2pkNhkfIhV8lI=
`protect END_PROTECTED
