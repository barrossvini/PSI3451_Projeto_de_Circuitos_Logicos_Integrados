`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NarmRf11k4vceztWG0W7da0hYvpJS5X7k1qOzTVj9L/eC6CdQdJfKu8U7zmdiTtH
XDlLc+gkjk8MmxyebZ2cnmc3C0pff6ZhJYd0V5Uy1EKbSaGol7Zemlwm1WKcHXbT
yobLFlzPUyrBlMrJuuk1kOwE0RTZ1oRavvt5n2Kenhhm+R/EWdC1nrQ9+CVCx0ae
w3fNAWOQfRBNVcJdiog+qpMMyXNznYaPovVjaXMhNK9zgnRuMw47OCXmvou7yh1O
/B/dHvM6y8cidwOyQRGEH7F8N/UtIUTyAcBjfTEMUpRjfb9YWDGxZP8qu/ZdCJw7
sr4x0I5Xp/lHAwi0nJLRUvuzFACbuV8wGMhczagtGorkT4DYFjG7oRVk7Q1uRSEg
rHXi+ivQsOGXBZwzJvV82AA3iake1kY0GxJVIEYwPRfmKI48MQzPc2g8i6FLiuqC
jgR1QDB/deBMT8+51XU6oCg0UTQhGAEddq9bYh2i6XHbwXoTRuE+TyRK5FhvcbgF
8RvT+fM/+NC09PtZqNJdruuIyj1ZBNhpwnRGZivF1bbB64SFCFW9JrSfn9ggnjBS
1KjGmUF7MOEfewKv94GGOAixjDKhH1NQh76oskU9J5OB5ASy/sTrJL4TOwcZFdZR
Jwwu4ymZhpKfJgccLCOdcnLdsdRsVsc/GZ14CuEZBnkQX4Tqcp5TYuSsysACvEUf
ugpd+3qjZkRIiQ6EqFITvTdqAxzJO+rFarhI+F4ZNVfHz04aDjht2WQQ7Jv2Ak4e
/D+6sTTChyMHXOGxbw7cSHFANbht/ct9UGYf/STOA+vjstjuweHmFDx7hRPaBgZB
glTqr5w5ZXkZmtFuvrWEqgVwo6cXHoOewiWDweI83fHEWbUCl6qqBlDrTbVnqQkU
nCpvFJxfs0C4dB+E+j6RoKZbpdB/1tG1xC+YoiuU2ATRh99+gWV+xJHwl21+wUwm
lfO/oLkTkmPTL3PybyCuFAkpQd7UqYjANFtYTAhvgViWeqzfv1eWYsaJ0eSsmO3q
SQFlgwXdv0135PQmhA4Qbr95xIhUfDh4aTSRvzy8x3P2yddGphnA6+Q6lytJ+BjC
c0Za3uMEtvZZU+aonNDu3qJRBctWOVZmLyz1H+7HrwXlJOlmN0wumVNxwPTbZiCd
QRftyPI0mDReMmHF2jgnR7SuqofUoEX8H+mQzlZGvuEHLv73Y0Kj+WCUPLYSBaQn
zgVZMF5BVJeXy3MxpPfimVGhfRn+sTDPDmrUjHpRo6N8cJzgKNzEVcxnLYtWPWN/
QaLiZkOTJnhxb85oX0+nAHgIq4muHBlJY0e81xLVmVGZP1xYRAhVqxubbpSpcGgI
FxV2UU99ypBrexEwJ/YL9QUr1sFjzvnMgW9ni0Z587jEFx0Bszl4wJ+rMweANmS+
aZDsGjuc4RIYwFk83foc81fOq97bG/RVfnjlFWMWlnlue5i6i0mAPlYiS9STZQeS
glNuRc7ggNej18btJp20JbBVyNxIH/fBzQUy+R1KM8DCOgMQJwjPc4ehKWZ6uOjH
dF81K93fJfU3aNylaznUFkkcuvhd1TqvHxbWNFDYN4YnVHrG7YRWG5regz8uqmEv
ajzBgBu6RBgkQdq/CzXw7amblgF8zKuL7/FxiCA9Gev9Xeic/J9mAv5kPLF3z7jQ
Aw4SVars+6Fbe/2nUlJjBPqd6pjRQiUde6kVqB7n00r46Mt362x7J1S2FYhinbNa
zWdQ/vIVByp/K+B37xdQcjqDxdD+GNRtpdmplgOY3WPkiwS3GbwJR8Uo3H4M+zxf
c1/lS1FC4qmirpXu9vmswM76hRF7pxNKhP6AplnY/B68BbZbZZW1ygGEYXJUdMa8
JVJSoUNB4iammIjkW1XA9zplAtcuj3wXfx3h4010AC/bweCvOj6AahZGFOWTjgjP
FEE2rzWsOLD18zWcDfl1wSyw0/z8myDZyP4H/fzrSK4tFD2cJLiAm7a2DAVhfsLY
OF9nLuAwwsvceLkb9A6VCgFwaizZfJyVIilPCD0y9mKRUalMa48UL10Fq8uDC8IP
PWMjkZZ31IvwjxqPBPtZN/5mdPy55csfKljg/PLcSCDVnsaEY/Ur/c4q0CrCNPH/
bf72I/QkSOXdFrRA3JsSXqku9HXOMrfZACMiiD+gyKQJMad5jLAemlaTjPHVusXM
ilM7mo4yFqJjZgpL1KPUFX3gRY4UtGYrwvpDKy904Y1OneaEPqxn9KUgMX6TuG5T
eW0+pVxfkWiEwUCKM0s6MqlmyYT+c9ja0f98VMXhWmeGPeIZGFrOeQE+gvnnKk4u
LIDg+33nZxEVBi1cogIWxdJvrczbYUA3mudVXPX2Dhhag8R/9icW0FXHJVwpjjHB
7uoHiTeuyEYdbj9sGGz1Y3uwzxyIVXhZfD6nznWpCsx/wfx4xb5VKVbKcIE/DrRX
rkgnQpaHLQv/tQH9G2TEsxd4cPGPG75eOyDimW0IAs3hoM1NtTrznL1nC8n0/RSR
sw30ZQrB39jqTzy3g38nHWXMXMStBK5mN6f5WFnWBGwy/qS2n8d5fWQi49H1mOz8
L1+xET9b1BCpCD0NObeNxXADbztZHwR+al3xFo1U1SRkJIVybjRhychGURj/wYFN
ihokmD18jedRkXeLvjfoK3yHyDW9+VzdHkmYiMOPVCPBERtt+4zDBfsJ+XygMsj4
UXPrx6z+EVDWCmrN/+j1zOMth0j3mwNIuKc+v/mmuOK78D9WJEefPJnMHcyJ6AcY
y+C0VZFajUOHf6twNDzC2HeCXSuDou11DMB+uVON2VV4fZHNyRmB07k9avWeCbG4
MOzIJp9bwU+2qKacRMyJ2ZYE7RO+E8fLxmcxKaXuZcE=
`protect END_PROTECTED
