`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RqO5NbbeyGr7bLLptmDq3SgCzKT5T95P60f6wwwmc1N8Sgaxol2FsfV8UBRDW5qB
sEENiIs+jGasIUrBebbAKeWPAmLgxUvisSdAGKe9kx4SDwsZPNsW78q4iQHgoOma
FLdp8joSh5Es13/ZMJ2q7Mif+Jg6vdbuIgsqYWKostT0Zkw9aBUD8i/KwGx4AXlZ
qCovdFjC1QtyMh8lBYxMDcMfpDr2UnrOVWaIQGK3Xar+n5JsIYBjjyuqzbB5lZ3U
8jiIpJbMB8f9azpuP/vcwg==
`protect END_PROTECTED
