`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uNuAq0kzqOurNCCbIu2mLmQjk70irXgWo/28frj6TB/DjSV/5oV+e7s6kVoGzS2I
3TKCIOaQSkMTk6MltpX/6onSaV7Dlshbicfsdrq5lU6b+61L7g7m2VGrELx4BTGZ
IqJ58KIbC+RPESQy21zpkWSF6AN3gZYzZBtvp3HVUBf2vRPyOH+absarqsLvxsBB
msptrPLJlYlhtR5ntcQbFAoKmEH9KDOUUas134L3m9OVbIEDUgAtuV9MS8A384ZN
SZKeQukYliaVGh2O24wuQPYF9bpaiGJyxrSMDyBcL8t+WiRvqlcLVH/lkN7Xl0k6
4H2qBEVq2VH6puywSL7gIkH0BR+ExWmKrhhvyKXaVrTaMembDbQ4E5HOIEiQDxpm
MDYjrvnm2332sAemnHy5gbklojfwnkfU6mSBMkALG7Yog18GPHS1p7xM8Lk1/uMX
cQ0d5sjSYbm7iUnhIYk1ZUUBDK8bCZKQOoBG02jmjbnz15xTz0kUr5+Q5sWij/Me
pdsRFqqDGrakWOWaWf690XqfsUjVsUF6sMfIfjBFW7sHK/HBzhu2yJ3Cet4sKAgA
cuI7Jod6LmQKTTNrZ6hIF1vtNQSpxq0fSxgZif/3hqyvNN8dUoqcuyKuIFlfO9h2
iMSreFZTdy42Xy+J+BiN0zQe4r7/ATt14SM2Ne0HL0q3z6kunE6OPzt5ige6l9xM
B2AIYFRCPlrQhKED14xL6RaUsASyx/9HMeLpzH2gN7yeSCo71YsBjJdyI8jLfeOe
5FEGchKLbGJRVdfpqz9O6nqBu3bDxyUkhlcToINo71qt6jWQpXqKZlfOyuyl2DpP
wH/UDqdMr/QdjRGKALJlUB+SMZDuDlerxgxgT/zQG2yPWAqW0YZLYPKWOC5i8an7
bqpVj6aTj3I8SU9SGB6nhBvHnPSAIY0hENnG7xS/EvVt883EBh8VtcPjlf6UuJGl
+1FER5sxq709uhCJXaO0odZaPVVp/W+SLxpLNewj4bbjDz9au2WbvBgqlSL7K0TX
fF09hfImUUSGEZZib9P0CLUWO3gSgg93M1/q51MtMAhi+8UkhVesGs6Gyj4ST5P/
BSkf7gDtyxxtFurD3rvK8ZzzU+tBZ6R80QZVPmPHYVQztyIe7+5SjWbxwU1Izabw
MyKMrfhzvePVNg3khBkIBrDVxcFbSVCYSSbuonfrnTc1zXWk30i9QDiFG7Mw7HYC
AFv91VkkJYhB2rM19atkba4SM88jl4HLLTPLTAu5bTQrgJKFdvNdJD3FmFoOeGgZ
ya4Gysq/j4Gt4EH2z+UO1dMoVgeTuL1rfCAFCg/EPSVIxjvcruN8gwPlVURBh4wx
sQ4/HQlSgNAEIOrfpL7fiR/YzE0BdBddqonyyVpbGjbc+CV0d2h6S0ShatCoIogl
EgK/QuPc9HF9ca2UPKTGl7TsdqDs+rGChbb4WZft/YcL780TcI32L4wjFcOAlvoD
BjEeslnWEaWN8v3ZJj0nZk5mRS9t2fPOr/g2tEx6m0CaOZ1myq4ZHBVeARA/P2Gy
4t/buBWyWLb/4Ve9LyJpVaMhM/ibjH5thjkV746X7ea+Qv4K1RopCPXw1be05Lr6
4/Kzu303coBw9exbJT03L+K1aBPy2kiCCWKfemsFuCim0en+4hDm18E8cQf0AYHL
GwG1Q1vZ+4/fztmH3Gh6YoWy0joc+rCpVgEUrk77I2QGcMsvG/i5UwFTNuMxF7Pe
lvAA/YyUQqDjSAssT2QzVlvqYDhJZ4txDcwoTfZuiHLQqUa79bhFQmWJn7IqRFy9
rUMRfpb3EeUU8qQBMnYWfJcRUgyAib7/iQkbJV46aR8c8JDnY1pI6RBubmIfXDdL
Ed3HREVMBXuVRItmJESf+w==
`protect END_PROTECTED
