`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
igJE6uzCd9r3kOPI+HV+mSUb0qh03do+Gs/csOG9rzQVRsurVcqqT1pIbJNWJQCt
Q/rYFvaGKk3TU8VlOG2l+4oJOCpED1wWI8QbrX/m2o1kyFOWneEiwgghLZDrwWPA
mCVvzhvILiaYGv5k+Ynu7HjD1B+Hbr1vs/f6YXm+uVCuJNxcUYUXnjPRu1Ncqkst
RiNb7ps2T/zumBborOduBIqiNmBgykisTWNv9roDD6R5OcX7sNOuPaSCIa2E82Fc
kVSnc3R6V+Gl+tLTVBGTN2XAUo+8rkUzbVUQK8PGh19KAp5ry8PJ33jluqvRbDGQ
ja41RLyxwXSCmJsRMXgW5FF96Q3jH3SZDMopUsHBDSvX3VXCXyQivruOkzc3fdFt
s93FvZGL2egcKFFETF86oVRK3W/+1P+uUc8AjyTj/+SQDzyUZuVc55ZWOpqh0hV0
6Qko1a/rUmx7kEKttczAYII73MLK/4tJpL0Lrz+/mBkXJcvOmxibwMEJYhSB2gp1
Z1N13HBPbctGAs86C5z5GF/VSbIbtrLZPLaXKJ3LSidPcQqumOrkzj0Hb4enpEjU
nkwrLdOoopHYkRRVVWRWTbO7dZen39OVxxaw01bwN5/F8iFE9ZoBdaa+yiA3fBxD
HjpqTKwkSIK5WHGEWUPxSR8bbopt9PK0rHZLETtcGp0AtVRj+q9Tipwb2O/Yyiqb
SDoDLZDDHpRoIOT50ilnoAB0ZyUD1g7uqRloVa2DuJ+TYBM9MxdJZTFAjOH/Sdb/
hvpoT74Q5nCUrT2LqykBqUenFNfsIA92KspyoryBh3jBEQJwKoUF6qLjMYg4CJ1b
EAhc20u3HK/D+Dz0t2M4sn3J9gUzomqwZZ5lLBuqYRle1HcDFlWzg8vPI2yptPcx
RUrQ/MIXTtvIjd3myRSre9LDd+vJnL1wU2OtjEL04I0LoiJ6pPJyKWbbFcyVMYOx
buA07oOlMpBsQ224carNRRiLBL5Bz+QnAlDvZ2qyPlp15/0ykANauVCFoZ2DZwv+
J719SnNV6C5hbk4J3syeE/OzYWYXOSIFZQzZDPq7qVnEsLZ6Uc2y452perldgAWj
jnpl8u07O9A30Eq76GaBgS1AbVDFC/LabnGyYevNPkrNgbCsM9qEmU1LJ8KH68vF
QJJQWrnSBVoKW0+8M3l8vEkPmR2UiY3fHSjwKJrjbgUHL4M04sdOilxV6wfhb6ff
Fw3ZIbWuBz+PurMjNe5WEaNKromv5Kn6ny4qP41pSc8Ts40DKs0mDp5ojqHaOywp
xK5FOvk4QQ1UX5Ry2/Hj6rhEY0+ZXT91bnhl82I8CgmRA92KsloG9q0+kGE8GCHj
+9VtAxB5KxnLxmpbJgOqKMSEviABIQpNGe3KAX8ivH3DU5oXwt0KOS8ENAd4DcDU
BW4gCzGuVmfnKeQMqHJs5Y4ZMM8uHbKt2pkB8+FhGIk/rMSIZRRxUAWEo67We1Q2
O1Qx/7wCsvxhiglbSHKW8LoRK22hJMSkL5zChrXKrR6XZ4IuN8yA+ht9Fd8TGXo8
nQk8VPLjnICKJ0FZ2cT2GoZtgQlgWVcSUUFHpl7lXx204it7iZyBAQhq382Z2zTw
LsuSjLyaNW6F54/7FsMhHBK4bVHvVNqqfMnxTcBIxJ8rV8Z5Vo+zhey/mMHgpTWp
KFfLAz7a48kKjZpu7FkR3SzLEfGwT+fsnFWy3CLm4WqECcI1r+c1FPpbHUStL7yT
9dBFU2XC6AY9cw8iBlMvsO+MwVbSn+meCP6o3s1Px1pRb3LYI41Men5IjaQEhZqK
Z1b3YUrYaeMelKm9PLc2eiUcA3LnybSyALkdg1ukbfU9WxB4SAFAmF2sQCIH7/hL
4szGvNHSK6+bH8pReYOYYKW3YFwGKIBlsY4vsBpXPeQtz8ycew5eSdOVWC6/bYMC
XzNvEtUyt8N+XhtS/lvAyrgxAr4lQ9kyelqhRB238ELVDUH6Q4y4rn3v9kCNb01G
iuKvUgt00g8RsA+5hmrcBBhmxz21XRnAKeiNtRjk3fRT8YzsRd0atYVSTr4U+SQ1
pBLFc/sdlLP8x5RjHXznRRD3nqL0QFmetFjnWOfU1v8bUYEC7rSTAV8pw8HTq+zm
cUri6UnS2KkidQ0IAy+uokBYe9Rcce00Q0qnimFawYfnTjMJt7L6dEj+nKGFyPuG
XZHExiaUxMrbgbVz5JZIZVrdMWRH2kIlJN1amSzxsK30JlsFyeIsHiMR9ji4K+3D
FiOphMcVWNMSnvyhC0DEjgB9zcy+3gzD/Tak0cbWN/PLok2KHlOarM1QsmL6k+cr
E5sdl26yWrqIyG18kWsLeUnxYyPrY8L+WOWv88ltSudwFrhlXsp51rsIFQz5GoAN
41+GFbAuEaRFv5osbhrcdyl82N0xTXv7TGR37sGmEwxRU1+3rLVbTS8ApMpqMM9I
qywQrrTKqSiN1XO2DIQvcq9g5BgFzJw3T6bDLDi6hDyLcYjDaUEVAVuWMmlBIZE3
15HOZhv4PWu1a6pEyGxz649YuUnxADOu42cUmv1edHk/cxh9ZQ1LuTW0Of0nlx9I
NGkGuh9Jl6coNeNNWZEM87j/uwplC29tCfRyAdp/wQV/mdgdBjK7Tj2wyldvDxDK
PBeR6OtHa0rEnxq+nKeShsP+lGoz2+AHpgDYFQh1bJzLh+O5nVXspH99LKf9trqY
J3LlKe0t8IlJXRc4Ntob6xiDx7C4/YS1jS+O54IU9+UcYFjAkibV6NKJysd11u0b
6jii9LrnVIcbjUXxdrGCl4tKMwaPEypxCORworvU3Mc8XeFtxiJe74Lf161g2qh/
W+z/GKUq4jzY5Eqv3Bte9UsreLe9iTtqILcv9vjxA9k=
`protect END_PROTECTED
