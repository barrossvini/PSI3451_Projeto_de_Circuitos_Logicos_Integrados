`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XS11ekMKNeNmM2BUw/niZCFK8HO5Opc8gDoyqpAzVvU8SAnPzV5zw3q43Tq74HYy
HuTNkMPERytvRUcXo8AJLVrzGzs+69IeXO4KzZ7VV7Ql//x2DfeN/coT0KNQfwP3
otvto8I9BWQWAgJVJc38i+20YPrAsALVj78HfLBCYm3lSbIqdxnQLTKvkA8bF1J8
eoZkih4YA2KnfiQVf4vUS5XJ6IHULigQvzHLKabfqvF3R+bbb1+iORSfNyZdTSWZ
VecFcLXlzvqq0ZALnlxLGDStDQHW48pnS7tVyg55897IFlN8TdmSdKfvC9vnp1DJ
tqdhi0yjNuJT4UWBav4ayWI7E8I9VwR+xd3GbN1A+2NNd28bNhrlP2cWo0Y7BNGk
OSqAESAp0KO85aDPR3p1SvZNb2wDZ39l8heDM3FnOSuysdhXDBsgKYAESmKay4oR
w6LoLZ7rj6S8mIg98Wym3AIMCThS7SuX4bVNyY2I4SEP5imLFOca+Fn3A518rOzy
uU2HrR/hkHB4wajdminJGZuLZb/yi6Qex3K0hkiA7mF0h1Q9Q4mIJ2fz5aJSiWMM
ZTGWjivhBaqm2S6AVJBtjBV25OHvIiv0pHNJcDINQ46iomMc6IOx8DQ7TPsvVd5x
64Mq3Dt9LAxGdYKsOw+jsn3Be76OblL+1my1kd8O5Tyh+RCqGS1vdy/y/vM+AYTX
G8jvQoztaCUK7a39zRa0sPQ87uVuqkDUUJusvhoQmF2OFK0ArF674qDZ+ySswErp
FsyYvQE6itv4IT4qFwauFIa7pwWDJXJ342kVAv7Ihu14U2LulP23hMxjFnFnjHvt
8asl56B1hXcHwFjsGk0Xy1TFJCGX4YGWDvMrLguJe1anuli+iLOwAqQo2CWJ/WKm
VXqY4CXgv/D5SLLOqsX+hM48mrwvZNkC4NRrdG5U3IGkujJlt/m2ySzk60nHkIpq
VmcbSqTi4os+U19CmegI/Am0DtGZERvcUAV4Gb0iwd2JYePafaSjPhcka0fDEd4j
DmzY8v6J2SJz4qhtAcn+IDuy8FoV+hB+oF6uvKyK/rJXpA01/oNHfuiXRrc2uRrE
vUmvowgXAOvxKlzA+dGYXA==
`protect END_PROTECTED
