`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YB57PgRSQ5dlaywZrDb2TWKMtEjvygs2bl0oKU0gxKCgDiRF4iceE+0RW1JQTKyr
H5DxjIiJjECe/lH4cLFcUFwn5jP1pp2WjM/FhAEnWyn3ampdD6vy+QQgVHLweWAz
QDzOpI/npWoZer43m7+/vPq84bAQ9chYQYplvcGxyUz5m9bCwew0Xx+whOgKDEGK
whXO0ymsk6ThXyuWZWxb0bn0x51KBZyz82LXH8Qm5IaHYM36IMooHoUaWSfji6Jv
21eYukKRfYnD3ifZkK9rNTcbjxw+qjwx/bZD9Wy85H9haP0c0230HVeTdAlIS6y0
4DoXQac12ZUw1Z/a46A3RPj2HkFviKa0zi74XE0NeVJoDnHkCQkcwE7bKma8NxlC
PsJkk7ySZv/6hCfF0tGY6PXX1qg/AL4k2ECnOpPYBiiE0eqBOO+8cJ5+c3YaK0yh
n1J3IlxevuNohlsgd+t1GVwlpd7Z1+nFiNhDKArzexFM5Z/DgJnGk2YNb81nMClq
GuxzcYTn0aEg0CPm1Mng7Iiz0zX1InowaSY5KyHz8ScVTlntlcx55ZalSfsSZwlM
neLdOta3YMcXBHLH1ueNAsvT2y53pnFtYvVW3fa5FlC7WAKMEoyteKEpgCSHeCPg
`protect END_PROTECTED
