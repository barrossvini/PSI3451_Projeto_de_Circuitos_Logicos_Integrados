`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rmT615w10BMCgpPp0F4aNb7gJI6Qi3oeoI9sg/05dwHXQ5C6knToHiImn7yFZMAR
6t5/PLufcdSAPYbcyLr8kvBrrPZuh3apo0Xqo6WjOEMj0nc7MyPBkr6/yKcOp8JN
3p/CpfIKG5teshfjF3eZ7Vb/iUh3xDepUbirNU7NJXyy2p6NXECARz/XYbmFjMiy
30x7JU8WiP0TDLNBhIctRHZGx/KBa7isH8b7ZewI06cL5lBZb/mioi77nUifok3m
ZKc6eAtPko3kJvgt+VOzD42rbMlsl3fmFyPd2ydZdwhDYnRzmS04moKhikohlhdH
xoq+D+yRKRBFkizs91QCH360iGLC1BQy/4kHk0zdXQKenDb0A1ESJsfQxUSsAOdX
jdbW8ptFQ6fE1+KUki8ZihaofMMww7aYZojguFruyUDLPw3sXgcmqvmNEPj/rCmr
hFc1IkFUyj+RjiVdvMzuphMOmpP7V+u2GkiduhBoT+DB9e6/BkGhQ0m+l6eXomTq
CLA9EvYqJtX4u1kFQUY9OtrDudyCl7P8EHIcgntgG4olv43SZuPIqPM+7oxi2E9M
Z/SkxZr84bzK1OkHYXVkl3qpyIJefCEXvdNp+krGOXs=
`protect END_PROTECTED
