`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vlv3M7mF1HyMjJ5c/vahNZYVat5VWWgoPLBLCVqSufTkR2NjkVkLRofaYKIo5r/S
VOhalpO42+75FuH7anog0EWxLybz9V2ElTJNfb09KCqVhTB+9WV76Yg2PQefcyrX
dSin4VD7/BRlkJOGWvcdvepohubitnjhU0corPJF37Dle88xX7NXjhJin0zuoP1J
yC505il1uwi+BPAy70wqlJu8Nrz3vpj/XNJAkJrXhx21y1HPUKBK6binIVC+a8V/
uJI8GcDpy4iprYD8Th3ApN7yF0rUWSJlazgAaz2F7DV3Z0WUy9Mskq0jUrTAaNFe
VzSb6Ki3RlCZI5Bx3Hq8e3CdX0duEb9n7GpRYv8voFHFnxBkjFBMWYHcW7K9Og1I
RanrOS1Rqyy6iXTohiT3F2hSGzNkJCKpTnqOXlVx+1MsdUjFLpg41xAP5V8tbDkw
8M8aYNXHGLNHDljZRU4wV6PxjouyadO8ezvTkPF0UvIlbTduAzMTbAIiWb5fVSRY
WwPiSQFfjuvQ5RwFquXz7jYseqcMzRiH1NbcnDYfazznea9dFzqRiYk0ONv0wywt
KfGdB1agVevzTH0aEqe5JJDyCK3HPAvs5Z2LpJy1KnpmxHQSlnnxu3SNwmjRYD2V
gcpEj2/uj+vVsk+E9mmLA3QADTKM2riWU/00xPLf7qgYsjLBrJVM1RqrBJtHbVbd
UsAZN4PFb4zh1ahEK0m9lIgimj9h+NmAgbxlXFoXueaHjh7okUkYRwm5Sh2gOTSy
kmfz+9D2h3JTw4Qtkpt7ePYB9vYzPBEumnKC2U5mPreZhPVsYukIYwa5ODJ0SVER
48HHNlHlrQJEx50LaEU0MXt0++02EVmiDxYP7adbBdMzIHHWzbviOJrm2FFgUidl
xkmJkJUSId9KB6BDMCBXj26g/e2Mcu4W7HweWeYbWcwrZQ0Y/7WUUkcLjbB7qZgN
MGWoLPtcik3DPz/ELP6QS0+mtd17kr0jLsVJrXc7q/BhKtY0DWjTk6PskOt856HG
3XGwsPkrJts8zYUg67DBJYr5rUdcSRw4y/8jLOow/NCDVU5dSHZWGdOfnpFRr1gN
mz0y4nV5Z9Fh3Km1xc0dE6VGrvuUDM0fapYcIAftdQSEQHzdv7Uyj6iOjCbSy6nt
kez6sDwgH0YAzsuR/PFYkdQq5bi5CEhHNdkf2CQ15HXFr+cl3wXoo3Oq+U7hIus1
gUOB3nXELxIz+1ujH2NLTuIL48Z+sUw8d5I2HvX2suV7pQx3l/TRRNV+aoHg2aV6
Im+jOw8lFgwnNchY33u13yW9lfDv7P2XU35qk0oibyOCHvk4oSQUW8CFPrgauOmV
xaptrTH6d/jA0HG2F2nnXfgU7tIun34a/qktqBhLGYsaNfCuTtG9U6LxAREeFtfk
N5rptpCzulp6IQ4kEERXhcDjR1IbWo+8245NkYACwwBFighDOptlQaliC8C2SXFL
mSUZuRd7zMFMJagyromGGlN2QxpCj5/A7TO1f32vNQtSmfMsmIIpTSnHEOYwUL/e
XxjWryiI0cwpAVnziSjOm4k+C5LsTBK48FyoF3HhKX4TEV6GZpyxIHRDGj2XnFM+
ibiwl+iXP52WWPcJwNtX3Md5fjXcCRB7wlqaxmzUekii0zRsu8pUkGlwCMbpMfYg
l0C6TMjLEzn5mTIOPOBRETDpfkWmryRrxJPTkeImsTCZCoSgeGjXlF99fsv9oYZs
FK+gYORjroX7NdEoZekuKceZhmOOO3Zram1wx3I38Jgaev+AwzVEdYMdkXrat9zW
tleh0+6zwSsLlXOKczX2B9w2JXa3vhpSa3ehiwtyBFtr9UK4OrCym861OT0TSDBe
+/DI+inWxAftCurb2nZ4+sMh+4hvql3Ezb9wVg4mue/DCulN//JzLY0XMN7oA54t
x6CetfpwhiNf958nPAdsBHCno9Vbokk3J1TPRwwQ2j8fpFPC8lWUghUJT718Wotv
2/H4pRr/xWLJ6M70qYjaKgppmtQlbYCqM1cnZxNKAD157y6fWXGri+H+IufhK2Fx
5ljNBJ61XEmr/R62kPluKm++6BNpaUBciPazBJ9EqWCRg5BesYzXfB9aLgKuhxho
ZtnyadI9vDCagufgNuoqwibgdyzJ0kHG3rdPYG+2lRMR7HOhLlLdt2aK0I7CiSIA
sKEx5/aVjKJcSa/dgDNCXaDUIi/UGRbyMLLLleOFXq5loGDsrv70p7PpByAx2G6m
+nfjx4ZsmeWhmehnebO4CDRSSARvEC7i8PuXa1At8S56ffqIRY9zAAWDxiNZJYYv
Tk3bLVx/wuhg1b+Dkne7uPASFc83azXgeTVHqmbpAk/zD8K+piB2ojFDxOLcclKt
dvNWFJdciLeGpmoT/9YyJHJGZVtkcWMHAP4PAL0LFfljUFQ3KZREopui9gO9f7Q8
kuwzOAFPipt4Qt/KI4n0ylCJFektUqZBR2nNhfF2RAkZOCrYPOnehvjh4PexspA8
ZyaWjCe8Xw9CDGxvbDp3Mu6CwJVMGJ3o6pjM+Ol8y9D/4o6GZc7SKiz+/K1Ah7tR
J8mZUI0JML8vtacOWJDaKXkO6h6TXXzAdCKbpgRKMu43gb/m827My05E8TsvkVGT
23/Lx0pfF7CXacswZd8MsQBTYIIBilnQBtV+gZ/WtV30WGuxlpV/oSIXp7F2Egac
7/EqOUp4I6yh8XDJqTlsyRlby1EnhEL699No18Mx7aXnRP7egqZj9qN9M3KOyDT9
xt5sQvFONicTYJj+UQjMOHezq10JJlIixSCgebFBM6ER2m4PEyEaBFUnm9nvtCfv
Rd34/JNcGwd9BNx3auNHsQ/h+hJh4C/TwAShx1NXQ1/rJZ5wdS7Kfg1AY7OEsiMm
ncQ9ZC/z5LaH+c6cvIJMpcOrzZh0UcGdqmI0hd0/TYZtm2xdAT9Ainm9MZUDYQs2
Be+JpLg6oXm4UfNJK2T1mCbtvTDDESJEjTX25IUCdjzhixm2nOWUJ2OSE5C91EXS
yqqnpBZ3rGagIqnH3YdWcOJJitGS3U3TpUR7bd94bxBLj6KB8SC2BaRSInZhnE9b
hvCNkm5KvyZcQmzcgPt4Ozlr1hJeNY9VeTO+fQAUax3fQDC0NZqj1DTB8/yGH1TK
vyjiAZ+hhJ8mfhkVoQurV7IeydYwH2nOAICyQ5UlaUCGBrjNqW1QMYtcaSKT6v5n
bi/27D5JDljoF+yXcD2w6Nm8cBT6vJ+ERq0IaOru7f1Dc9NxP+8o4VduSGQc0Z3S
DKjE4us7aHqCzAyquJM+fAOTLxwt71QEvZ/7QM5UncKDAPiQjipM1ncNIAH8XStK
hKmxRvqO2bGneMyB+TYoB0g/jwJ+oQUrB5VH5UWp0Gzk0TYf/tpqGWQtYH2nDb4a
4tJlLO/Mbt7qRLebN9+5/uJLDVWF4xcajPIjKq6tUF7m665tbL7f4u1ZGKlyXW3T
O3hHru8cbGkPrKVtPPtulA==
`protect END_PROTECTED
