`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0qzOH7eCayLDFiDsBX4MlJADMVUZuunElRbRGesN5hDCjnxiquUvVndumd4TORvC
ZTZnkP0geLZ/+8kcvZxZoOCQEtayaA19/lFCGaJCIm32D3Negfz1v8YvWg5fkgJ0
aK4Rvo3pX/0WHPEep5iAS7om4qZgOAsvuV5a6N2sjikwW3JQ5s+A0JNWsx4lATQg
QOxBtxF+CPt73M1/S43UUKVWW4ygAo24AGKDe6RAYzOxXeof6m5cvpCJ26A64R05
L8Yt5WkSPaASXqLsU3Fl2SWSX7RwDihnnF+ZRiukOCgGqSw3jegTav4W5A2bvkEh
khOKuXwswAYA8qA+5QIr+NBWqA3b4KjQiNCU5MyEuYjU8dGyIknQ0eEUtGJihD/v
1BXLsmICqvL1nfOkQZm+TKHcJwRO/TGpY/koaPk/Ign719onmDPMqHLEHw+pFr77
OG9lnJSeePn2+vV+NjJC1y0Fpk0wArDrPfoH1x8DCuk1MoJ8xexSt2+ET7yCy7eP
Tw4z42paW+r0JqCocuLl7bUFuVCI+bvlxC2ieNh3tu9JumOGUA+ogQc37WZ5IeB0
ofm6KAFrzOUJJEh3VfyW+Dl2/RIIz8ZoB8XswZWqJy/elWyY9T6wmoQwM6d3eSiQ
9tZrveKedzFVDK/enMAtL3SGnfNhCJpkWca3gK64MW2kzdEllFbL3Z24wZthhXxj
lriCoB0hrmgcsFUJvtWmLxErW3s32yK9s5EyhsQmwH7n3ieVXTxJX2zV+ao/gW/2
+Vck2HvwATfeYCL4uod43U1xq7zErtMESeBPmvOn6WNY70jKaGLMax+xDVqLRHOB
xw+72Rj81Qyfg+uh0zQlUvLA7gNTPCOG62hdKkc9hT+uvUD2JOMrKrjjG4Lv6/w4
k5fbRM0i+k8yRR/8+x0VorRezVWW7ezD4iLtW2nDjjV5hT2q1HKqVW0kozxmkMFY
b6ffaTR1gg/fguhF0tukzVDEYCSvUthXdA/wR3BEGPsRt+01B4V5Arzh/FwLg4Pb
mA48MhEVfYdpPafWlqDCrtBSWRn+T9q3Ve0Bpu4ldH3/MaTGNLCEfTD+d+yq64lD
lUSqXflRY8wcC2IVcL8jiOnUVZ0DFKRy+zWJAjJqoKqb9ZAeXpNzbHGHyl+en6Pl
dKq9E62FdjZkIyuOdA7WWhnsFuACaCjxQ1pFmYN5SjAh8pGvi5JV3YB1iKdTQp9z
2ZxhKHSFNjsGCgLsFvuBMBnyJl36pVkdZXqri3fEm6w=
`protect END_PROTECTED
