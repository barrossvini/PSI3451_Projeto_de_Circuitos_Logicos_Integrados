`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CchjYGnCdoeb2VtM5eW53FDiSzn+J253SiYWBULHf3+xM2iInEnpl/pj7g9XMqqg
UZINGnZz96o5kvDTyJF0RkytoHHEO9eeWrsPvOia7m2h77ic/AqEsLunrK9jbXDK
e+CzXjf5tzhjE9Qu2NrSLXrmjdcg50Bo9u6cmMD4uG89V2DPH88E5SJ6+M2vB8yj
BpqIN+GBqYeZDDb97Fd6j4/meLuNjg3Ss4YN+nUCTCOPn0tYtUYuAzOAEetYvind
Qb/yYmIQsiKoK9SE3/93B6rdk997yylIi1rsk9qKJMk2qZubfjqHXsQW47Dka852
ewd6R00fLVeiT3ttK1JzldQIIHjK0pRuUyW7oaYNp4NUGhUdd77mCPBVSfK2l6T/
skeeAxcjp/9tkpNhQMH0nBTcHqElpgINZXIkrmZCmTWwr5GR1/5pj6ClV2SO7K99
7YF6k5CUf6PJ8ySRckf82YxC7D3chhRtVAvFoKUyl5bQZeQX3Y0/Nhah+beOrVKG
Edafbi3wWOg2hSG7O6MVQaYLQDBQsPVXVT2MNc8z9GUZAEKxm8zsnvavMYWDFpQz
R7j/xHN6DmIlYj9V+Au1lsW8UoNOM5YWTnRcYxa8S7W7/yTdID0WYw6xssIkYz8h
7d4S1S8RTqvahow9h+WXe1WJPKU9mAQvjyfXl0VlAMR3Obj/2iLmU+p5savOxWcR
JMFPEerypJZwUhsxacPRn+k7JRoIjOPD/NX8MADtWtEw8bpafTKrRYApt+1+CQY7
+T2sBn3qDYXENYEIex4BhEGqtSmW7C9vEPLx6Ycw7Iy1fXdqvBPQu9U+nnhXRl7n
AkxJyfZ5BtPygLID1TFB/X5m1D0f7pxBvrZosjxsXCdzKLVvwPZ1Gxy9dCm+oltT
qYG2OkHAGaQ/1mC/YPx3IfN+0/8RqO0PdJbW/l0D/8xkKGSh1q4MwRBoymlabV0E
N032f+O/vnBJGkK33wAMWkA2DKspvY5WJwZ+lb22vm7xAdas8fmhd9DwN17BYMLr
wJWu81wbn5pxrKTC+NaC4b03Cte/PEJmEBQpkn5bDdOB+oEoYeetMm/6WUXYRv6A
BGCKyb4VaDhiyDsn4spN2/Rch040XWVN5BsVZZSq5IvcjkbMhHmboPtsfK0wFylt
qm02A+D9FTW9MKXz1T7Ov/2sz5mLi33WDYhz3E66mwfpKCF7VLSHxeengKYxukEC
jqkKpIe99AgREC79DQuovRjbz7FsrBImWZDQlwWta9oIbiyfDq8W3zcLaboqrAk9
`protect END_PROTECTED
