`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0L/i+cX/cWb6I4RC2A8tIbVxu8Kim8eSIWFQ6gX32VfEjMDxs30tdk5r3iYq1wPt
pYzmqLOAa/65GZzzK8kwxobex73vr2qAqMh9o8kWKnDe7IHsoF24fFbFN/R8SeH7
4j2DUCfPDlSTYvPULSckhmnn7FVzhB+s4QpjiDllMwv0H7dGgYezSdWXTDSk5UBQ
JeD8P758Hq1KlIV34KpeCJ+4oBnUZ5JlQN7LAxA4uAVzj9Yu3HkbxLRnCqdZRFlS
VRswBUpV9m0ETAVZHmuTSZOCzqon5MxeI+nIZQ1cru93rkVJxlt3pYdp02CfJ53P
2Op4O7cyp9pMhtAoU4myTygagsvhpw7NvbXqhjbMcCmeKDPFrR9c/hIXTFm3RuDn
W+k7wF22VC1DWqWZbmPsnWLEuuZ1eWkCxQ61HnYzcdA8+piKD8izREPzVEXJB3DD
17+WjfODpLNOxt5jJHcZ5Zl6bEBJdui7pEgjNPo/0sRQQZeMKOE4mP00zOYPnY9F
en3yg82YG32lWlcoc7z9soKU3nYiI8p7DRowYLeKWc5ZpEKHwvLhxPbJn3leTY+g
L0Y6JqKWaw9KyEM2mCTt++U6RuSFhSUE/kFNtpGosVOjcZmgOZT/L8gdVLBL7Fjq
/BNblZrq/nbEkEv4KlQFid9+S8RhnXBk5Kma4A5NTv7d4Nhhcd9UMbxLUnASX5Rc
/c5tKcWOMvSi4tQZ8DCpe2mFf69k+65SxvXY8IGg0EI=
`protect END_PROTECTED
