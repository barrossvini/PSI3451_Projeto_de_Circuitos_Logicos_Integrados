`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UxTgYeryTaxwuKLDDJ9dk/Qbua+TDuCWx+O8dZ3qoVrhinTB+EoMgQO80X6vIoyf
ZQ0k5i9012Y3ng94u/hLrDTCX5IyMQ92SOxkq0v8PJeiXZcEk5+O4fIFWfR6tZZD
v3HduZA3ekBrSDzgBcRskqBNseNLg8S8etwBwy3lMo9m2pS4za0wjK626FHiCg6u
5ApIbfYyNtTAiBvViJzUyQ==
`protect END_PROTECTED
