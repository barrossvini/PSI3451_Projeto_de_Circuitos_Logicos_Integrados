`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9b2/M0fEEpwuP7bdR+N5C5Z2g9vPxu0Z3QPBZE/d2ooitq0oMC7V/BwYHf4Tp3KB
/hbVPpsjxN3+/pFtjLZyYT3L04bVvxc7+mIFw3DJAtra2LLK+OrSJSxC8DgO7YVS
YSogMGZoSrMR0ucgiUXVYzNmUP9UFd+5sRRiPdoDb2g=
`protect END_PROTECTED
