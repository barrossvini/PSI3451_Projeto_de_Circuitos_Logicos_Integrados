`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2AesYTNyn2cnimdnOcL4T6JqtMNkIS1mJfuZLLA1mNDm0QlBf0KMTuc99pNBVxOE
heCeQmeIbWLnYwGiFVIqMaaEo3XhODyVzSNDcDfowyqFiEzrNlT6+Xo2ghKKhY4/
AyME5iH3q66kOeRF7KHU6cvlcZVnH+yWcbAuVnT/Wi2RQK8LomeBb+Ym0WAQUqLb
jdfKxftJUB1TBZ45FOOqPKxN6/NUWoRkm3HMXwohcXK55J695oXsOExhBTsNVUbM
9hFlNjbtoc+5EZL0NRrR3x5xR9XJDURJUieq56AQPgpd97e9u4sh9m/GT99mLi+6
wmdDj16P5+lRjHvrialpXdZxqeFcQlSiUrDCgy8pG0FBiQCs52qVgrNNiKe9kc5s
PsvWchS6w/Kn0lBl+KkHRKz5Sm8jp5MRvzPjfvljZ/m3EMiZChqsE68FiSdVj1Pd
zzT9MLxRD4m6MO/BUM/wx1tp8n/34JdqurFatzjC9cLYLePiM2wYaXtajCCEL85x
XduxCAdanW4607vinV280thtFbfCGXKRNuJ7aAfw9badqqwPbsPUxXfQCJ7pwbpa
sRv1afVXCUyeXjI+H/QpWU4PuVDb5fAcWyDaPX+UJdNqCYzWBNbX3d71qQMyxK6C
mEWJ+o21aVbDL8Wlhia0rKq+CRf1cV5m/rPc/q3p3txTdtouJaUjBQQJ1VhCouau
8Xq7ptOPiFENhjlk4duwiO1T6ch/WkKEFfrGnV573qT9UxJGkuLopJIcaaXy4Ria
tsP/TUchzZu+euEt5WsZJ15qmh2hGhevLeKtrO+oAJI34M41SNnw3uaZSWHwQ+ZU
cGMLaj22OiDIrnqFC6erBaocOFENFrAeECRFLASxlAe1waIob47bMf/3s/EZeBW8
CpxYKNaaH8SG8SqalBa3EZodbKcscSup0zHWniKEjoODsga0GPTRtb0CZ4q8XO86
zpozYsjcBWD5WMtHLDI7ceD7FgLSsF0MrD1H/WSZKzyDhcwdFm52wnjOTfgPr8rc
VPoVITJ5AMFv98TMfBpokLPaQFOTftdSxOKeiuSK5fTUOqwsGh/UDraTEz/WIJIV
sohF+CErZ1TlHn+uu3oObAI2+iFZPj01ZBqZFUPyp+x5voR6pWfJbtWPd4VGBeNc
ERCViIQ4O+ZKT8ap1L5j1szOEbpQmv8Afcvdmyjl8+QKwlaMGG8eyZ/tIvor0AbG
yAQcy+mtNQ4brvhiOWIXX6isKRFU+jQZBCqbwBbkrq+KyDAjvBcJsdlseNc41Cuu
X93/TFOjKm9psquldGRY7b5CfdzjRlkFQPYebBC8Xnzim5kOdSuHxCJGGpoIF8y9
8xB3tepa9GerJ8x8SZMlJZhvVqQRORc/0isKhKMGy6jXm7WcPDQJtf99LpHDraI7
0XqT8swI1QPJfhnY42fUc/v0J4/ECGLzJECdL+fJtc8jgefOtbtsyofL6K1Wcu+j
9vm7ulF1z2Z8zL+Yk263IAGnqibYHk47zRDktLPLgklRzJ3cCHp6SZvObIKSXvMS
+sKDDOuWuMUEa6fbFoVrqX7MctcL15STIO0ONIPE9yqOjfRwtlb9RrqP+eHvCuZV
NUWOFY270WP7AJGdOQ+N8MEZPpiSkuTSiFsXV5o2v1SkOlhm7RYUECXjRLIXcsej
BMTAWXT5+x0vSbN3arTkrMJUmaRaTEgeE64qbuYEEudFw37OaBRFwVifYcW5fh/j
xMmW8sQxmY8LwNVZBUEa7TbcGwzZ4DA6pfxcx9JGJ1w=
`protect END_PROTECTED
