`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OsjZG5FCTWbJx/S4MyaeWHEjyPmZze6OeV9BTGgFwFGCJUMgoOjVxOxQfke/VLsC
drf8amMVRKC2GDBZqdzw+r5/FopzBtGalFY1cMh8R/4FqQBFwjE5AZAZwtUz7WoY
wbNXdyUKF+tczzRtHwu62D3MUtJkfaF/3nB432cwGao+VCarDv6BYyI6L9I1TFnq
tDoWx7GjpPOheREKuv3RUs6bXLUHsbtVxYwbe0YeOHyEvO4wCx4C6YlBTDNXH8+3
kDBZ1Yr/j5xec9wf3ySxhOTf7wcvCnNlyKhwkpp7o/WERxkpQM7MlH2hakzmVF2o
Aw/E6WIBEe85Q2MjnKbR/6id1d9xllc6uh5JMqLiRHpLprYnB5Sttf0oV2hiQ4cG
o2seO4rvf8ju05D38AjuJnj5mo6mgnIaFGXZh5MdnS1hWC2kypNqkEVpHb1iNevy
JDLFfBoy8cy0CbRQj+0XM71UlqKQ18YhMtFtK1iiFeQU4dRq4EoFU/e+xo0p/wAk
731+1bcVNRoV0s4//1aIeV4NDK8Iz/XvYiQrCfdhmZSPO3Ef2IQRgb695azptGCP
/OwhySiDRV3XA0BRdJ5kQMYGjyGmIIuxEcbwVC8lOz9gbIbs8Dppk/5muDdg2wu5
P9iCf8rf6Nq/plveG05stT6Wl0wciknIDcbQHdSrPAj4PNvvVZmNRluT0Ydqig6P
nSAPk0VPso4iYjVsxwOa7yc2vsnJu44Fc1lG/2U27dAWdhbmR8VP6Zlb8E589cyj
SLDnxskMzkEYSwlwiW49Dq6wU6kl3fvGrQNjwfns4gizjG8Kl3dhnOR/YN3VS/QV
qAkeuvKK4a5Fn7LiSuOuAVWcuP9+A5fd6KDeNExWDxJ2SPUe8emiuivXkp2jiMhj
Ir8pvJ1fx/gPVbHon0KiL7CovVhDorsqm3XjIauzHW2xMjc0gXy9ITHOeuUQPmnt
fwpQ7nr/KBsi2YdwWyE3Z5ikes9H4tWw6WhAa7T1R88/D/3nNwGKJtBM2XMZa6p2
8iUHPYJdmvgrVoGnvh+qecUYVv09mha+CDrGt4wX0x/0E9UeeBTqTTavZmUAoOV6
0AVPF3zK0XInJtxoRoAYEL2E/M7+qYQZKXlSkfCN343iYB7Iu1hZoB2phzIRvfUA
kzV5Y/E1VOptU6CPn3rCiTV1KSe7ABZnqj8yXjWfpGOZI3jZY5QK+5/0XriBfFLk
olBnlehXpmwTcgNUOEekfezkk3qWZyIq7NqnxQvGdkkQNpc39cHWUMUhaNMNerxg
nFxDso/RxbkYnGZ36OWUyt+LSJ3rHXO/nkchK3u8eNfzSgXZqfhUgFjr1wA7QNKT
SqCc7JFaukdDJ/T1qLx3UFvwqj1JeGcUhib8qjBK07PpG+ufu62bZEhTpZ7MwfSW
/MvujIAITbwaMIL0hnV7JezViYL5dvUvwOJWOrTwIPJsstPHYXTqupOZRvMh7BxC
fDEH0BguF4aWxlluVzejQoVQEc4ZIczxdG5rWMdcf8OrnJaOXZBFSLF+QbPmAohn
nCeJlFMO4/Rr68fBaM0++yEEAyKvTHjl7tjNip3PlLs1ar62SsEGDLttuNnTK9bB
tj5XJvQXsH/Q9aRapFMwRoLnRr/+VjDD88JSICGDhCEBWlzA+AK1RDFF17K/H8fl
FBUBLlFyplfgz8VHUhrHCU1+TnzbGD69UvCcJ9vhmubT7PTYLmzaM4yo9ZFvBKs5
4G9m4z1seAhljNg9PZ2yMx0FHtGR8faTH8OkjaupxFujGX9EK9BKgri25epvZ9Gz
6vQ5XjRGED/+fmQnH7gW0Zffxr86DYdL6z9qecPPekaaQq1joLbSmlKKal1ibFdl
BFub7A8j7UISkJ+EcN85mkTSvCBSyqOLF14FYHyO+2VKANRU4bzWgCFAIsk4MoMV
YrRJNHs9SNTOxQF0MwX1tEF7ZjlHWTq8DJ5KKr7j2RJxopRlTn5nJCs7v7icVZLB
hPJkJXMH1x14jtQmInyJkiHqDOFtIe2gaOPCkz4R3XFMUQ7z3lFQqQyTD7+vODV3
Sq8StwccxN01N8U8zcuZjrD8S4oal5iYP2lwfB1Ol6CJ/5lOt0XGMjqlyrBT1Fig
Qi6aGsWfWxolx/VN+A59Qa1TZginEzYDu0hAvPyfHF6uC/q7Jtw5lc0cgrQ9CEPK
RWuE+uKy7IvJ4Rw4jktL5Pa7L+nW/QMCtRGJjZ6gnRGEhK4gIbJBDEVhSzbIcW2G
KVzzZD0a/w0oAsp5K+2MGj89SuWiLbQXTmYKPSJOTDCWiBEV4NrB29LoLK7XS2lA
+gFUm2ZSLtYOSjEbwrpItYjonBLHkBhOlXl5a+SW96Dak7gOwj+sVeFRu4bQfx26
`protect END_PROTECTED
