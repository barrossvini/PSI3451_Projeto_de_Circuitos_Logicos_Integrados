`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIYqanFrzjyFotrS2VutfcNejthVXITcqrQI6RRz6qCejeD6qnCfVUca57Fu4Uw/
12vCirkzvCYO8Y1tDxMilPlw82Vw1KXjZP/mxPtfVu9PGNLpy6t+cnlL9ZxM94XH
s3crHOr7ErzsqssAoTkb7TT9AFS6fjAk1jxaEqtRD0/2Z+rkk+oG68Jv2x6CU8NS
lJpAzQzycInh90p4+5htk6ty22NbtjvFfYwhZFLeyViyqeeeCUb5yWDLTIDfT11r
T58FBYHhm40yJGNg/7XnWTxk3ECydgPAYjipOrofRUivgJj80sfSc7JV+2TLakZk
h6DEq795oNV2eyDdco/GHhd2KPo2c9he+HC9uwdJQpYVs6E7OQ/n/egrvNZBnO13
qqTLi1URKhyoRBu4qShzRcAR3moLC6DdZzSbkd/ftLFUzeCtku7z9kExAJuj+7yw
1GTPThwOnFCiK1/ypNiQKLomO/v/iDFXA4mQB6lnWw0oI4Caq/gkbXRxzfUUOGYk
Ed+TBUkfrh7p1nHOPYb2iEm/8zD/71AZcf6hJBlNgNLwJagyrYXCm3a+WnaRFIF0
4HKA+hYxC/HimwkxN9PI826WUqcWUjgAnic9AEPSzaBOMyJHL7FRjIk7pDs0aVAK
nR5ZIyt9kPyja+NS2g8kSAZ4x1pngCM9QOv11yEDOqDRLPiTv9Ra7cTRMh5ujHgt
CvzTJcIlv9wEBeBfylfyV2tQgeJum1srMwkKL7ZXxLYbkURSaHcGp7lvMmghmYrD
l2x9WIEotmzmqESlaOM+AVR4N67EvCqVveuPryAlZux0HD2s7oSN1ii45bJDHrtA
GM2hNFyCCu0J2Q+GIxzctDWr4swDUVYM/OEXG3UxzByAyPT0X6KSV9mw8lAeCPy0
4hAsy49jqrUI0UdRjX1P97mQyS0DH83O1RfEpNzGGaPjFYaBfqhM/PYqNpAg7FHD
veenYDY4B5gpTqtx4Mrxjyl7dAN/LFf8XjY/w2quyucjlWIVOMUuD052x60S/wo3
6jAgBVW6TkEMd+Yywm+dmTlmK6DQboFuAkhR7tZ967sMgHbPWwU2MTDr89a9X/4P
BFMxgATTEz3cAfijArwh8vDlTRoAgWlP+apa9fxcK9PTXkSPgXnVX0YLpUSQVTsS
ojrO3Nd+hSwVsVVS2UDUnapJ2hG2J3nSjZTzkkSMBzQwAgklxTfZ2sRE+DY2iE54
DOphNnT+941oA0QFGWsTFG+i8RFdFI86ZtITg4lyzKdVQRIHmgzG0dPdJ1w6BSsb
tM2POPU7R58ShT0vxMoKAaZlm5YvXWcgwLkhaXC61Tzt2BRRotQVPLUuHSbDUWs8
GHsSSL5sDWgBAGvdXhZotOM8gOBfq0JbdYoMnbNN+Tq0B5Hrwi+Qym4Pgcgqkmuc
95bJYC9lEkUex2CxvujGmoFXD/QmPMJExwIod0BQe9U+XVNne5ZcI1+ORkXVe25V
ECvEzUGY4nzlYP63Gbjk9/aCFVUej6m6tThaKgsYN8d/EHgI3dMtgSm5v6KSu/0B
IVBH9/v7w9eB0dHyzb3nAxJdW4D6xv5KO99fSxXqP/flps0Rtb4L9fd6yGZ9fafX
N9r+YxyeY/PikEbfaEyLtdqRw9iLYfOpWTvdoco63BidCBsU7pqLx7F/0uI/vsSF
j6sqKCyHYCgDHqJN9FnCLzzNhhe1X+yxTAmscz/o+S2y0Ulhfl70Ucn3JUU/6E1O
r/x/I8nkVqnJYXGr+bT86WRLDbe8ybXst5WUIombYLK3Z1d0zoDRNZNVRxvHJQHj
1qLthZFYXUdWlVkXBgMKi6p7DHqs/61V2b6lBtQ8xXEn2xSqJPg2VsIN8KHS6q/i
6yOCDpKHk79ptMOKlJW6YZ39adl+5md90ZYEKnUErDxWIWynETr4HCHRHYiuWZiP
rXos35CXEMuDztn7Ur6PMCOe8o4B1Ut89q3Un5D3zv8LtlYp6rt/w5XlJI/xejLp
RASIYREeuSFwlwXLg4tPEko2f5L4DfJaV1Tg58WK5A5IVoMLsi05aeotw1CX1/yX
miaS7K5quAQvXQf6joysEf7hikT35sB8zo8hWyRplowv4ReEvHUn1F2BPaQv/eHy
EaZTmbb4/UzoNDCHw7H0wULGV143QCpfoWXEiRTu3I25bZc/M4mwPhYuKs8Tvcc7
pr8KxpWQitTAqbO38BhvH2VnAgGhxzzlIb3pcsDVrT01TmQFKz6b8KdpvAFKmQ86
+bTO/YYwSB4FUR4QjbZHdU3v3rkQehqjz4YlmwtnJd1tnFH2KIwkcCeEUAjtNtvB
Ud1IxvCnVMR1yOpQGTlK2cOuR8RWoOyyLvYF9Pwbn/oulqh/q8bsYVZMeHHgE2NP
xwjmXJ7VpJN+zKw7eIFQqbIvuOh3Ve6GS8UOYrvCzU4Zk29wOzs73PRTccYJPrIN
zZfMflIHEnAOoQ9xwo97Q8+4K/PGgHZ1SxX2u1hRlzeap/fM181xvfD/OiTHgBjk
+8fScD4N6WCjnwE1qhVu1QmwJD9zimYZj0lDmmizgpgdrtZCGgPNnmZjqmgnDL2F
jqlXKmuORhumh5n+o2QmjCAkt6MNH3FwSmBDBryh621HeW5JUj7X+fh7s28mVc/d
Ehc6dmqApOjF7fb8HHurG3w/DX1Rt7y5iDx8YoGzdldLGBzuXzt78p7aQARer2jQ
g7ALc6LR51S9LfSGBODidCTOhbgNKp40VcStYDCHxMGg/jOoGrCmnwVlx9b1FYJr
z/wAdUFCK5DSakh3ML6pGpG84xogxKk7U7Fj+zgEUMu17a+GbSsXrL5nY9wcMYc4
OwS0drhcQDOFcJugoLoWy8RVRG/vBuNMakyqnnBJQ3x1I2uAUVI3DDgLm7GJNCDa
sEidlwK3hjJjpcx5PuhF6Dc42/twxQicND9u2nAwmqKfvuGnyB7uZhSEaecnvOL1
RpCQzythvuIzZlTbK4rePoDKlneQjSmJVe3JfVgjRNFYNqSrW990NdYLd+4z2y1e
QD99yLyIhH4LHJROV34lRMfWJEPUSuuj24RWzpcTP/9dmBbkg0x3B2p3D2fvO7sL
sbWv7m5D+3D4MdgmM3tJNJmtObaeOT8tcpwNnIf3s0WEwtmsLzpizZlGWStWoIyz
tUoC56JfwXLqoO5eGpXVrt84qdZVWFo+yOtTVCbRK8bArkaWq155k0yWXPXg9vod
p8rDQv+g72r0oPZt4ecDG8x+mSSwHL6qcCQpN1M9KecxUaxzgKggJ6Tx2bExHFhP
NgF9fc1mXNgInIyeFZNsbIhj1OnaKgnvgwloFvAhl3MwbaIquIlgpnswRXRZU57x
ePEVztICxitLONN3cvLKF9OKEGevWMexzd+L1BZxnIqscWLKc+RYpH2Wuo0o0f/o
e1ROzDjE2ZN5fJq6zNasi3z+/8E945/4CoBuR6xiwf28Bfsmxz2csD65rZgkNTqv
DP0UwQ1p+CKXAkLYuq9NePF1JBLAmcCX0dTGmOU1w9MzK08hcBU658TOihU7+d7/
oIPRCH1GhFJmxUbIVWYMNh9f9AhOLAykCSn8xw29UF2v2zbdxD708q4vmjuLB/a6
Qn7GXimh+DNsed1HHB1pyZtUXw04Hej6Z4ya1046pue44lfYQWhBu1Ep96jzPcWF
W7krWiVOCmIU7aoYw64xzwNFw7VJp69TNeNcs/YTxCwdtimLYHPGGmTXdgBn+NEd
Hhs+LpeRBgjQBUHG0U8grK2HAGO+LiQn/BNDIKOLXSDvd+6/PLZuy6fHeUv5Paao
EmfbcrKnOZAlq578UhxGIfhRmxesMYTDC2BKMq6jTN6DNxURNklnEkED5NENPWmi
UCbUEn7sgMxDr4nWMxtBNrH6N+v5De4F6YBQaiv/moITLah0y6sWE33jGaKKjm9Z
56gY7/xO7sCEa0c5c9hJkT94RqDZNrvmcRfn72ohFQLVVS2KEMhTxYf0SSodnwsA
QSzAidkcL93CzlLKXfUgHKxvVbD117/JJgQpy84t2pPKJRE43XebHaxNTw0skf2T
Z0M5m8cD1V1AvchrcMoNaE1pkrkKym4+/lzWYbIe69SUNCNPdqJqd47nlxkA/Owz
/+PTA1fN4Tsfw8OU6E0SuwfZg/6cW0ovyICqDzLBK87TbPCSdY7dYpGJqAxK8tzE
Z+UqaHTZ8KQfgirCqTQJUjy2Z2mN0nr1FCvVB78fyV7Hy4MahVFjbddhBhDcl993
OULdQAimmTvaZAx6HiW/xasCzL5Go8j9pxzd2PVXEaC6oAUXmUK5wCKKqe22LOAx
TeuC2EYuW1rls0fKp4my/Cr8bOzoVXFrvok4yPKV1qSLjznFzJyGIC5zfoOZVkzT
Jsz1IAgh0ivmbEHd1NRsbXF32dJTmxZDmRFUIZVtj/F4fFTxMWMxouQM4ImhGRwX
4HYV0tLv/9lEGr3gaWpI4jGdzVp6kqkUWeXmrIxiauMrLdDOhc/4t+CZDbHcYSk5
KvJZpPu+KRfQ8D8jg+uZhezxJ2u4eo/tKq3PhTO5Ax89Ml0UdWnJSsF60RerQ3D+
j0SsjXCuEiSggoaCtInCzOBaGvkvyaxh4HnJT4OGgt8zutztFHEhIZvYwuJLKJYr
tm487VcnulJcZnKc5D7rUDS9UG0nzsjSRn3OPhvyR+Kvwd6hAZ67uW9s9ozmc4kC
2WrdedsZChREl8j2YVw5atEaux2zzOJvWF00CHeZvSdMz/gBjkiIyv9EVVpD2K0U
HBTMp2TKKF84xlPgrdlrqNlKUD8deiHk5WAOS20MvoHndnaiJEy5YpJ011nWwQlF
+VYXE7c9t4AZ+FNeAeuaepGnJEuLjkyf29HyPI16ie3kMhkPot6EXqXhaIEYmEIA
EKHPCL2DDF49BAUQWD137vcL8EKqUKkQHvqrqV+WKwrmYdo/C5UPPaq1rvJssN6v
UFFkOJnK7gsx7molpLr/IaoIH27PxGUbYAyG9Ujwk9pG/LdVWormarvAMJt98lY6
E4dLzEGcwmn7+IyaYIN5MNczcNQTEHM8r3PB5hYUrr85989pmL5ovKfC53cj+EUz
YnDraCd7UeYR/WtZika+6YTsW659v8Pp/gd9SwOjKRYkR8ymg3yhiTgOFlTRtPCA
eXlQSDMp0rCnqCJ9ourl2EpA8u6ZMhbu1lzLBZcJ9hCViAI964h8a58QibytJVFt
G4G6w9/EY69HOApXEpbCm+kBxTR4ofO4y6Pu7WSK3vKBMZOUcTi4lqmqMzsM+m30
M5kol8JJmBdXvp/jNDHR5CZQAie7jyQ3qk48foRT0QtJU+kYSbLNB5RmaYDEXfBD
GMDLL/tA2QRKGmDn7mdVsxYDyllBHfIMtmomW5yGHMTSL9L6r/odXLIfsMUa+eiA
WuD6gjZBgT2/+xJsOfBonow9FTqRA9j5FovF7O03xSfKekQ+g+Pvnok1Nvrz404P
N8Ao5l1evfwc71iOM01DAyyDCGkJeSg2T3dcAw7PeTCB60fNicF6E1phoFffHZ6T
6k5ufhAgEyAffxRg3BAtrnT3Zw0Gy65WfPBnlT0Feyy48o+/p6j84s7vdN12itzK
sKmMOfooczwLWKCfbF7ISdlvcFqvk9JbZwbUi4cL9U3fhsve1Egb/fLWuyZXqN/E
DBO3xO/5JpJsPalfIsUzJlaT9jbvGJ42SBHntBDc1DIMkqnyn6PpABDxKuBPTDBr
eurKLX+3jQfUsc5Dd/HFWY0E5udqU3pW+CvzLRlLAHpKbyy2ok0cgXfVryUPb/IN
ZRsAYxDrDoBE1fqQSqtqEkQtskPcuntnU89PB42aIVaaBj9pl6/IK5zaWCQ3cM19
S3pVPgRgKoMBrjw1WZgZdmN84bj5dYSUgprsNB2Nx22jMTqrgkUPgmZp707B3x5j
8FfkUuastVl2cZVB/r+zQ3+tmOOgkaxNTcz/3CJyrAR6O1lmcwNUizQuv1EMmDWD
Cblj2LY668s2XahTWuD8EiDp8p4gp+QvQ9Ti1tArfQcKN4CoC9M0ktpj1uw9xckE
AQ3TB1O7BhHhSdrSI1SW2FQFhN0GOxK2WKJd5QKe7ky4LxPJcawUw51jC/0EIRQb
HuSEyYUkK8vV3hx1B5qpPCsjqtGWdt8caOQrNqLERGjFbMTgKFnvCXLQuJXbUWoN
NJwnbQcQeFW+GOmfHQo/oM2pw08h8pbfRWV8yscisw8zEd7Mi2hdv/7q0dqG4ua3
JCN/LWgUTmI5JJJy7orxajzKVZhJ3gTswp5H6c1JxjGQJmsg1s+qC1sNioUxUpIH
6hnh4Y53QrcUUiO12p+UGIK5093D0WpUfj+o2uOSPU5HQ6I1guliqrL6P0KL6uPq
kH532LU6wq1cDc4f2bxZ8KnFU1mIboAKXbGNcqyfoqJsK6jVXKOtviuWRyfkl/mo
AtMPFw5UrLmAVdPSRigqii75Dazcxioc4fZj57ffAC4sdO4ES5FzbuLy+EkSwUBz
9xO1hbyOuSW8qxhrXTWfeLTtBEWUl8nWXHSFyyeAgp1edLCqdeIdDSA71VrNBLoT
HRdf1sbkrsSSTmC5uKzrVqo6EuxslMHyyiq1Ww8nnvIKuo2rfq6MgnMrpu6+NNQe
GQxpttaZGOcQTt1VcNAXXWP49MOCk1awmdmy0cRbdE5Re4wXtc6LzRlW5qwu2pjM
297WNotFAr9OR4ZOVV11Yf29mxZKg1s0bmE48fms7z+ne21rvVoBiQ9dtBoQcXCU
zjJE254Hz+txCTn6CC4MOaISDgeV8fNb/oEo+uVxiGPXxfZmkFI2VuenBL630VpE
4XrcxcUweWaFwDX26P5jJYv/6BNxQHKZx7McXlQjx0TDn9+jKmPp4jKya3SkKVjr
n8x9SoGGS52cNUT3hYSUW84sgUtAz4zW6DJa+ZKvOeQH9j83YQFKBhTFJbZ6UqJE
aNI91TeHE45jQp2KQhboabKPDJDGZitzROAUVJwH24bwHVJyKkuf6SrfilvYefJf
qbPrKRqa3KQ7H8mQxVC0vHpZvVVtO6NH7SckclWgsFqERF6rQFYkshLXg7162KND
hnmouVtu8TWU5rEQD3SOK8eGz2jLAU4vXGVUmLgMmwQFnj+evMD81kISPgjw9r+4
tj5f4GFzoJbzzc6Puyb57yiV/xOd0hhgSV31czWQa7lZWx0rQ5i6wBvoDjnOmPvM
ZSkcFH+3TSVZnufa/FrjXSO+S3fMWiZpqXtw+w4VUcddpEMGfAGVqpwkRZkaAaOV
LxNdgKEoawVcJDVZz3AIf41kpOT/EWjnki4hIvKI6/B85C0oDZAyV/lloroCWC5X
M53ELcGagfZ0fczRMxHg3Sita/3GwKr8FXryNiD52YTWxBxrJEBYJsAlzL5cAuop
RrM2aoDZCAKJHsfOL/6bt9XTe3OeeXZL6b1O2pPOTGUB8jEG+tO59N168pRYzS+T
d5hiEye1tJO+1Stox+rVmsfeIqcytFy9b7GTXqpxQ2ekvuIJ504bH+avFvRkdXfh
7rAo+H3f4ozPJ1sCdfgLsnV95pUW6RWSatF9S/dZQrZMcDAJRsKLnSXw1yUYRqNW
A6FMgQNGJkI9kotnh4UKffIkJb9KKA+u+FU+DMJTEKa7o0bcpyPDsdG5rIUK/tre
zjqBdNm0nfje9/DUdOFi/aUkZjdHLV8FxDju6R5+Hhy6R2tRq8Ev13OPzZ3rp/Xr
HIfTG8TXHu8BZ525CBJYxpXPZ7/gLqWs6QkVva1IOflSp/unuclMCyl2Y3RUTPL7
bonr2YLHwigGD+8ffLSxxOj5Io1b/3SioNmm7mG4O31W+yGW8mSdRzZUE6ptRS01
+x1uHAvj3NTTYa6ve07nj6T/MMN1U5Rahaiw7EhuDU6+RkfkHacaJMCldGo+o7W5
/DII1YAyb4oFf7el/oqRPeiJszZVFs0roCCTeowe7k5Vq1sxq84igxihtJV6KryG
g2xj7f9QV5wIPO/ohrsL4xN44KzHapX1XguQJB/3LlFk6z7pNYUAcp7ySmzegczP
oMHtkySDGM6JEtvk3ou1wWvo/Wm14JkTiszoU7QYrWDqEl97IxzqzHOFFJArPwod
PlR4AiBQ3Mlf1MacAN+S+U47b1tfFnPGpwGss+RxZNwtwIt4aS0JPq/4B2yh0r6j
hi6kQUMOmwqC3AOUdPq6k39TEbg25i7oQ16c50NGZcApTcxtT3dE0ewsxAuZUGuo
mEL+La9jAMYaWM8bfjoGxF3GyOIsHbhKgVblozWf22dLJmBk7Ozwu2YGKH+kr4Tz
i6RpcKo5U9yEKAw8UQfXOUySne9ezqzrAmWW+IxerSMbPvDC8fg1ExTxhyG2ZsVc
OX4MAX1DOURELJznrZowZwu+ccMSIc5/wwedzLUmdoH6YKhWmvoU/78+cJeS1hN+
t/w7vtfDrta7aorkn1YIMKZZJxdOJi4rlbMkYm+PAzqKL0K8rDBsMAtfpbbwzKtp
l2zCskm/sKAMR8aE9Rr2Y8X5MYfnRm1P2PIdW25r9pG1/f0JLOq9kiepiQ8cFtGC
wPCt46DH3tP2/yvWn5aBBbh+ivH2uOWPLEyCspyn1G3k6PJKW7GPlTWzhcu3pdtf
q2w4UjMqC5x9pzew5uGsJMYrbJnYNRjssP58dyV5zKRNZPdrcPHaTN9UnOnfx3AE
/v3JQgmenughHfkWCI6LkwGFJH6A18PbknJaw4AoVyLGLtLbY1U9Hv8x0EmW/wPB
4VFXqoPojXeO7W5F3Va3Ys3sD7M4gWV0vZRIxjTXx9GfQrXmGnSUsYlFtxaZGdIV
YgoFrJVbiIosyCh6xLZwbKTMzrAdVpLw02qTuNfF/Z0l36aY00aIAXNirRYhFinB
tOagJISWejO0WouIKQAeFJQw9gdNXKr9IC9XC6ch8d/xEY1QMGHdg4IU6LfU5dUl
tzvjMAKehho14OxuRkhb/4U1veXaxN8csnv6Sq3O1/vzvPsPjEk0Ym0mcURj5rmA
hkg+ptens6WUgs5BoeLvv1oTE/uDzM9nk+VSYOHQDO6p0qq7grF8oSSv2RQ9Uhtb
gVQz1EL2tXx13E9cZrRTD9wJbET4VYa0/1AlPWi5HaqSyQQ8t90Kl3l256nCzvvc
R3Dna6sbyVh5B90HwSYyKhtfNrh5Sy6wXxsm5VMXoTdhb0T1akOsBsKkWPr50YnE
vVaN9OxtYbeZ8lViw0nTf6jjtyWQBEbfKcIrlqm/00zQvI2ZCM2X0FBehrgP2y3G
SfDUGJrGD/SUSQozsqtJgccIBGVCsQqIjVG9MnAJ5Fr97i7xW7GTrfJoefR19aDp
9zpXBxrK2yxcP6VcCfUIkwqK6FbXFR06D8Kx06Eg7fP4NhlTOn8d7UC/E2FKlDic
XUk+TjSJPgxaIJJLIA7ZWnxVy5aZ5jfnpi7rZEH1uY7Sk8vZ8dLwzwy2KKzJPEYD
DlYE/VOZ1gdEGVUX9qbvUrIXpmQ/ru8V3d7Z46sKeFUTNLopioxtd86P0NwJm9iv
xt7sjQZMD1vBgsSLdaR6qJg70dVyX+t90xb43tAghdwK4p3MpizNxD1bxxJLggUQ
IMDMF8cNPuiKEs4yHFz7kNDZwhhoglVcszjZHq1zVEzZxGPsKs44ZepEV28fW7Ol
/7ohbf+ndLhoICFyR+/1UamAMIqx6BFgAgDv3V8jy12ZZYHTzniOThR7aMsyCzuc
7UJrKlyjGekfPNas8MPp8lATqqCN/5ieZAjDfoZbZiw0fSqRHJhi+OawVHuneZpX
usEam451UyQ+OfkCoEUlejoJwPSxPHcrB32QVImcb86MLx/NPUxcmablnBs/dttC
Gse2pCs9u/orRgiZlShbfz3kDUhAO1jD3ZZEobfVFvCW0pn6xynuEEUy8Ad9+750
ARYBCzdvMBg1B47NZNG46ADuFN+ccLpQJgbJ9cC+yTBoRCVMJ/99U1fESvMzp92H
PSWuNYHNI1uP9A/hsrc1UtjCJo20y+N6jQCBBkWAl921MOJbgkXXcQnqchglWdzL
zrwbBqeyzSCRlIUB64ZhYyKP4ott+P05ICwJiO7VWJI0l7z37lfR0189UERyt8MN
FUW8k6KppIynXIcxZBmYUGmQSuvKHhdgeX0B1VQrHaGp+pH444h/DJcB3q7pIK72
CC387ngt4Io3Ew+1en9Y4WWDnjcpcs4rYgTqJn8EO4B13RhADfARkFXqdPdv73lS
KH0EUhyT7hkR+lBVAvHbxfD2pTcIdOHshLtqqXs/x/no/FIS6ZOOPpRqspc9ZOXZ
79u9A4VCW14X3P2O9rAJ1o8PSKmCMo3ZHzsUS8wwvLtQ/QnrzWih9czMqrRrG9GF
OjrNBp72qWCy9l0no83OXoh1dYOCSCoU2xE2eT+/SvxOtmPs9g6kmOsQEWLxd4Zk
ZiKC85b+Pf31DiR4iSxwtK4h7PA3xpYPsw2LCrTIeoXUtvi+okMqflDnoliU393Q
wkkqRm73ilPCKQuNlYlwsTZJRSZWm15KJ24xayGeDHrd0ni0xNHfOZEhoLlXFKhv
36ndO3a8rOXzqrqPC4y+jEnDeTo6JiE9b4SCnGMTEB6URm0rxm3u6ogzx1anRxFe
hoAPBLsUCdMzHICtQ8uV0Avy6w/bItZFXztG83F3CJyy6YZa0Nhg0NZQDHGSSM/p
73euFaZAIkRr1h2iL2sH7LuX2RTAYjNJv8e3Dr9zi1QdDoD/8FvxNXGCXrL6I0LW
6BNIMddMT3at6KqbSongiIjOYdilcOjP8oyw2ntZuZXuR4O993rPrtcLOuY9zKmK
gre/ZiQt93KciRmgNjR3RQeRjd0l1MBMNPUgdde26DxbqxT3dPmRPUn4MrOH5n2c
l5e5Ul52hY2Ax3XlqD1FWgORjSGjCd8AGlqsNGfYhg2DcEKTPYyVJ3adFtyZHb52
E/HpcEbqww7snfOdxOSh+pJ9zj/25s4tlMXDFUuVJH8AtQdG6Ehy9AF+6Ews/nhJ
oOctMEFiWXzeRTKh8vUMiYJDwzu9z3m/L/FTCg1HQWSODWGEwwtKjJwXA+21vnRs
wIWL0jYoKIFx0DMe4woM1Q51wWG22QoPje8Jci+wGrVOwsVlnqcyyzjIg2AcX2dF
cnY4fU6oyCDthwliGWOjMIi6G0oMNF59J7UgUQ4AI8CDy33eBNSOz6GBhiKph507
+st6Q42m/tnDMkiEoUGI+t11ubQMnykO+UgpniJo8llvRSMDLSyPOr24GTPMwlDs
9quJhg5HGlIEtjMOeqGP25TJMn7hJGncsH0/SYVRMzticMEQYwNj096UZChUjoLW
phVt1SIjlelEWj6eU2vJL7GfHOEWx3cIqopo+skRVT2/Hv/H5Yjf5CKgLi4CVyra
cbmCd7tJR2uaqTPOvKDfmWtFr1GGh9MMGJ9vXyyDf9JnPKQVKhYnln9532YFhm1/
0R7g67ZzluBHt7ggCuBxj2E7QZT6JhQs3s4ahaIPTDJPQrOdLThdld6tjktaKmRc
y4KaDHO7vbE+MesXUHR5R7bgr7sYsvX43XEbItMsCytUUxlCm+IKl4aQ7qT6BEea
4iT0tpDR/f1MEoaZRCqPyU3RNvFRb/1pFGfjTxgVI8rc4d9lHnv8Caj1ShbiFcPv
eW0jr7gZb0x/Ay7LLfXzF5JrMnfhx9+unpC9h/poudr98DEwjAXk9xOQ5geem93Q
FFAlbS/sj1s3E0aVvJl0VUmuEpIKhDL12vopOftMlIgqR2fjXqDhVgFvqnqXe1Hs
8K2YeOssbWmOB96KJD3tHpybhwVz1U+gpaFVpY+PcwzTKnr4qcN/yhPyh6obh7y8
6j6ZC0lqJfheVzom+CIZjd1DTSG55AKbMdy/YtNCgj4qbTPLUHspTsMKAhQxC6F0
WgNTNT0Oeu1GdONhROKmbXEAdvmtiIPH1zJIU26H/SlLMg96Z5NQ2AIJj9PfITM+
cnw7fhy8wvcVw0oJWuULmMGBHZ9j5Vu0ehWXbZ7x72JzJ3X1Isy2O37SLWxCwcOt
qg9A6t22ZMLFIEY0thJHlL414Dw3lcaywWmlwkx4q1qiNOYiE3RSVVtGAUJcQkDj
VDqCR/EMCroZMQKrRGq3PhR23o2OOJ3Tpi8pumKtUfz4NJGTPNBHipFSidZhORnR
Io+9X3LzDzCTPkQCzGzs/Co2VUlWJY94Zzzn9xIJNIt8yHcka5U+cfME1xWESy59
ynm3P7dBXy+a56exTSAvcbgpBcbINm5M9/Ho7DlbBxuSlWNnijLxHWkQtF+/KgfW
Jfw53o3ZepoNMxOF7f285jlEtS38vw8RdumNU++J3ZkUgsy2FyVPmt9K+i7X4C0z
TVLapWYRdJrcwFk43Huyqmc55T47veQiVrQwxkqoQ2PDmojXvQiJAxSnAyv6YxXj
Po6JY8/v1wUftRjz19WdpLlZuXZP0fIbmSTTGTJA+l7C4a3XaUga82hlF6wvYaWu
2Xe5xJjUZ4D1xLqGjwwRc2rQum7LS+fL4z9iaoKdeAw1bIrQgYHow32SdzMJdGdh
VDuwDVyPT5/thw21BJFa0CSgcI/U8iubB7WfX3J26Sz+E9QHlzKceVzUeQbKQ7gw
5KP4i3lMve4mBsB/EavVcJ7RePaBLN95sa3QVieDfT2OdCzIM4+CCNuagV9w5wSU
UIOwf4AeUtFnFcY0UQ/lgd2vtAXUmeTnELS3hvvAal0AI7Zx1xz4wslPiWvG1vjm
aUl/vjShRMao/CNqa/oSWScAtL4WVuCQOIkRzvLxrWFjiNNeZTIrydaajlrT6j5k
wRfUZhg+W8zrpDlCtMiGufGj62UCV7nBflbwGCG91Y+F2mWGhr+JiqwjemtsZuXv
YGRtehpX9VDaIGYXVsjJFHQDSMc1wBZ3hrDLGqF4t/f+tya2Fzx8qUS3K5ZLGIll
ZZSX+aN7ObmuBRwJ6oa8/uoDSOBIMVamxf9bcUmhwVY7jeGZMJ9WRndHwWLhhP4k
FtFy9ncJ8bDme8apKzvwzXNih1nIEb3X+Vvj49UYFvEUhg+MAFLDB28ZTJDN/NXn
2z5tdbvMblUtIIH0blP1a9UC6d1Q6QBOFB35N61+af3G8n6uPpPhgNSl3uswTfZY
dRBb3pnAIG4BYnWWN+L0DGed4TOCVF2Y4THMr8WHXTUVICSCdGYO9l8vB5Hii/Rh
FBmXSMVH443hZjuxBalPCE44drLiOyKnjUBhI8dErA+G1jUtxcpiceKuP+/gJaCE
FkSW6ZnUQf/arX4DbOVoDgkB+ELbhZq3iTNFHhZZocoggNlAKoxRNNRVV3y9+9Rn
iXoAoIgMbl403bkldt0v9Y8LpSf4DWoJmhH7dx3trgwDE56RNz3hywz7YKFsX7sO
EmdFaKasvGl8Gr4UfymrrOuD4BjTC6u2CdtmBf/orLDitcZv1OEUGsh5PjX2dm1e
yvKIsLiWDzPB5KZMX8nlWMAHqkH01Z8nzaGsVydeRMasgJJK3hNJ4UjCPVsQcWcR
unnWZBVx4e7UE786h5wbw1IRazbDqheelQtZlz+E9ZnDtd2sJO24TISMDbCuhBC4
dwJMs+YL+jqQDV0Z4aQiabOMA5FyvklYOZetWGLgclH9Xqy/i25xISG0WPuaZCj6
LC2xHoUDhtdjopfrboKr5T46TXGcfQvjio0JtfcRaEficdXMZ7idsAQgPqq99tag
BwypcPWBUYBEJYmfNgWkrxGppwwWIq9gx0MxYH9DT7pQ7+7+pP0tRTRtc9bWgeG7
HPPYUePMKp7sFS33rzm3vYKSEX2cwa3mzbSHV1I9z7iUgxaJ41tsLsnUE/G7fS9N
HDX/ViI/KEiB9HPPQKXOsVpC1xNf6n3iT9PCS+eoKyiroNEY+9Kx09OdLJwloM0Z
dlNICvJbH29pyYJ0Vv3zGXM5SRi9mkbnWP16sU78QsH2p9JYhFSfiZwzJ4SEiNBL
+/RxUPWgc5aTYVU3nawn4zT5nj63qcHfHre027ppIDRggSA5reXitGdT/VHKaSQR
NwooMSFjO3BbfK6MIfx9XXE4FP++1P1DvmxysS1UfRcSS8WuDIGdpS2hdcwk+6sH
VBwUmh88zBVWuQwSej+INfTp9crFe6kXT3AbSUmDPpNWlFTNDQdi4igLfTRBMFVV
rREbPTvM3PBfmP8FSgtabtAUQwiEutB+ax7MRjoe8Qz1qh27RocpBocjGizfqFg7
WrVyV53EY+5UOzPJ8s+mhU6MIAJepKBLN7DszJmPMM/qXP7YawIXgO5gNkvyjq5U
fIW+drWRtkT4zVmjtYzB19pUxWVBoBOLVOVI5XaNApz7I3OcvrjImaJvJ1/kn2Pi
nwsjKXSJ2q8tWfYEl9ZcMiO1Sp3kTrhz5skETvKTgbGI9GV0C3FhDzKvBZWUVV0q
uyObOeKj44Mu8vLkRZbXzktf9i6JFhhEn/veHLPTafwJEQXlvWyHJKYzOZBo6uWx
ufJz/VQzvhyOrOzBfpXJXScbSJDGU6ND+mGZWYDnWnRRDKh1Y3anIrR/hxHGX5A/
5zHqbA4mrOU6E/uAOBtA+cMcPXGS1j8OXOlsD3PBCWb65N9Kdg5hJby8ddAtVGea
sDJaQf4UuSCqPLssSZPKyZhPnxJ7noyewAwhWTmP0ny/bb9rI8aG7Nu73RmIbL4R
wnT6IR12hK9wEmeSoWpg6QRGAVlgkKJy1apBsL3Hm010w9GVCf/rwpqGlfpdH8g0
y1+Q+uPcdVbQxvAgT65xg5UGh4Ny5Xm3KgfHsY2wERe/IXX3RBshjMZXXw6X1yRJ
SRX+xWEE7whHJAWaNfAXqrgsa3ppmpCzDZPV2aCYYqB1YtQiVBw5gfuhhqczchXs
uIEndj2wF8KRuErZyxSpqrdQ6I4MMiN20zfqaeT3V45V1ipxc0JeRlCvo3rP8yPy
DJLU01aH8PsNg69+HMb9DNXbFb/9OaGZp3hbhuuAEfDhsTYTNQTy3MXqHBVXaEa4
OWhkHF/Jre+SPR7J+Sm50SJOj8fPHyBNOUvDqZGPvVTsgXyZAjOV7Oi8SUxO5k75
2QXFWBITT2Ze1a1Xjabz4XJd5mreSyCGRDxM+T38jOW8Zj6Z1eEdSEVdg4krg69N
r83ftQKXCg4EwCs8UuqZUxEX/1l38BpmSt49GngPsgN+aYJoZqAJ2BEdVaGVgNXH
9bnQOVpjPTTL2Ph/14r/Io5trWJ72Oc/R7A6EE8bm1qF7EDwXky+zfqJEm8DVi6b
7BkaiZ6HhEOng4NHXbY/Wz8rjYNleaYikkI4BXCOUltY9Ax+jsv+z9RAkWDCvVpX
jGSGo1SJCd1e7mQ1HEpICU0sgXUzPUzzHDi0LcJF8+8VdnAn0Y4L/ZH8aRbGjckN
SCZsG5y2bmSkMengxnzk2QhSvbRnF1TskK005EpOkXcHeGwYysZG4L7R+7k+kZuH
7n6XPrX7/+VL4LJs0ehmdVUSVHBzGrZEeU8psoSXPsa+BF9RjLddG9HOtehO8Uas
z06psv0N0QMo6EDiCbjN91UlVgTos0ElgcQo6dKonoswh0InBb1y26VfUOlnzrrM
X6QtBfED+UaQb2w0JBZfReFl9Y+GKvghkWURuEEofK5xKBMMkgsFFzUpvQy8aQ/y
b0pHklJHVaFhXyZdpmoDYnad0FMOS1noZV+yjJks9jTpXdF5HFQ0ozkuq4edaCeM
GAST3R/5uFzrAkUa6VgPkhxJkaFbLmvs1r4VqQ+8uIiaP2xFdy0MYNUD4SJ6G+Xb
qRyWXY1zhSVamhrhKoSsW1BMrCQ6O1nqdBqPl6eCeDc=
`protect END_PROTECTED
