`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NEgXaOlKc/Htr/+MyBEgZaq6X9cI+fNsfLT70xOFDYosh9/sMq3fSKEPZynLCYoz
s7+CFl10DiKpPNEtrNUbpfSDBb9XBWRcIzGm6RF7QItbRq2Y0WL6I7ZUHGeJdJOx
epHGYJhRWWUIyJaN+qWSqMZdIkfjuVu8Goz0lllvL1LKuYH/l7TW2yYlNX3/U2yu
Jt8L+5wWlhquCjr10Rba+79rK4FxObV5S1gGk/5Vj0gmMl7ExMF9K0IO0pnwOfsl
e1nrcQXfXDQdgg1/Ay+0Afsk1YJY2bvpHRQ/nvwzMVt6y7Zthr2dZ8FacDADDdin
GNJKVA711clXchhvrG5uu7YCxJYMkyM6VSskGtdPNSjXGPC6mzQYAtYI4QZXn6GE
JuJojTVZvDarMwY0n6JvFQ2B/2ePAz9uo/0gnnTS278hZRDSlWggYYWow2CoTsOO
q5RlvlX+hh4qQ1t2TFnVSgBy4juq6EHOVVyzKdmPXUEnVz6YtT521WsoEqQdfLv+
eRCINP7YIiNt1zQR3UEnFQSz0UcCkbuMurr8s3YQsX87eCq+GzgFOw/Ts9io5Xn0
gKyjyM5PomCamz7Ig/HqdkNFvnP9sgbJoiEC6qjkKZLNNHqElFY+dplyOI5MvLTV
2NzF7i4gk9GTiMucoEXcI1h59eUvsqnwoc+h7kwptgZaHDiIAhgCqqVj2CA4cU7P
ZsSbbqn5FXgjl2pRkuGr1a37+VVh2VwEzzEWufnV9F9F48aH9V7NrkL971IFPUbU
fuCDO3JpjfC4YU7GGklyGdqQ84Ogotucma81wtCcdBplfGlkEab5SGB1tyHdDhgq
`protect END_PROTECTED
