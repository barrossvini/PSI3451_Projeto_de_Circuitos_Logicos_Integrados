`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FFfvmRAxJSGF+Ezi0h0yAANdTfqWFruIC9PnNsQSDeMaWYDXvAoYJkJwUKHy6p3s
U8KnsJ7qYtkFFKzjnvfUml4tg/cY7Xt7QytnzKX2+cWuAU+zCEqtqcR2/vuhQToS
G0pLS9tdUaN+zMJ1jgpMySC2rKgM9WfQnhu1vyhw/70KiwviZ68v87Az5roWivB7
bp+x46uKGAna/al5VnEwfha4qDNldQS/2lqKi+GK3bJPe5Do9RaYZ3REVr8ZhhL1
zVwCYqg5FZO2Lg226xUXzFXa8DCVkEmcDvPie1tpV7LoOxyFLGFB+gCGKsfLjvOx
atesNRS0ULsbsrRSeemgpSi1A92SqdZBWhPzpNGIJfgEXl9UzF9yShPnqvEJXXS2
uqlqSJiI8nfnXgabrpBL1Ask7JLPjQDTuai0YlFaF2P/D+AXgySA0Ztc1E4HmbtI
peZKHF1tmjgQ7mQMXTukliupBp96fVSDwT2vd+5xrvuNgTxDENU7iVW6asIHhLf1
Ny21iwHoC0dIhe43A85zl3+OUNsjWeF5nUoPr81pTsDD34V8TThf5qvRVwRj/Zo3
hzSZUIsBUheRG6llpsimQKdfqOWXI6BbvlEKvt9kmcifz4iop2/YmplD2uzeMSdV
w5m1q5JgihujljsZwIUbPpsYmeilMD3UpuuvfkTy05tTJgSh7at2Paaf+/4TElFP
GPU5OGbvoZ/SvwSVQlXClZL9/erAfe22id8KwrhXJBTIi45RhwP6sz0ldVk6vHu0
6IoAlv5ufR8QSEZhcWfYqXWN6tKYSlpeZ5eEUfgax2twLyaxJjOuiaev1ga02shN
DJgu5was7nEDj66C1hQhk+iKFdsTF6DnW5TTTq5cECVig/9Rx7OpdoAmr4z+6K+v
FrS0urjJBQNvwWrAtX9KPlavO+0kmf9UnloDHb4I7bOcvHmZGIgUS5Aro3sZ9a33
nhyIEtH1wdRvvacwSjLQUldZsP711pZAWqX4Nw936O2kbRsbz+fS4OOMLYYHO7LX
sGJ7GeeP1zOQh6jB0gB7EgvG2rTnMFyIVNaaYWB7PeG5EKppCUCuKz0WYX1LADyn
TQtVc8mW/TQnEYoHR3CQVw==
`protect END_PROTECTED
