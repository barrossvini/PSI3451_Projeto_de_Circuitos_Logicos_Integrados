`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+sBFwzr9QFE+iS2Dt6oyGgK+AR9cQTktibtvmVdf1TcG5IpVjzsKoekju6L8tfQ+
w+5bzgX6oRKN/mcbSI9KTIBFBrVHbn1VIn1f58tl82dvPa4xUBEuL9KAAbam8uKq
B+G9wfl8YqJxCqjOqfP6lPs4CPT9A49xS/MfwzllUx2o16DoN4Sz8eDmaywoZ1S6
acJKC6UBk0F8zfXOzkLi07lbIkYBmtgwTZw4dW/fNrvdcABbtuiUjqgzdZjBNWKf
/jR/z9lceI7HtD6xjLY9a/r8ElRH8LNWZhKweINtRhfYLpPRjAvJLwOGd8Z/grYr
aei9UuEpFQAH1Ac3gY+mMdz98lE424l+ChDgjGV8I8ZPhlieBoQjyaEZOxIUMZrY
75RF0dScFTtDlnBlrrgU7Jya6Ov24g8QDNOzGMPVcrp+D/dRNGnYJnQC8TP2uaP5
TyP/xytlreejRnjfHxjX7MdFmZVo2MkUEOvSilC+k5gdRwQHgxLuxII0MT2ezfgj
0HCRhtyiSSE6RE0bUHQA/IFhnHmsqF+/sYw13s4w0WqYLqVjf9m94QYL5+AYiPjH
15hki91++wWKjImayXcHgpCmkw5/b+sUUm2qRGuPOsOxWxNvunFYrpNtAVRPPUm1
Ri0LPtLAGVMkXnP3I6Ykyj7Vpr0Earx/OY6zOKDBWOPxlgGok4Paj0oJDaT5uuFA
tJSoDuhUMx6Zx7qmfHoma+memFPnktqHqZ1hez1aR6MSMun9dCmfIkhxRZaFcDVO
L8R0XPwHVMCfhgLsqXxswVVgGfBKZiF8nmFKlDt2B8NqACHSZF4thjmw1fGrsonX
H8utfzFTJS9XXb3Gp+cOJsRy9JaHkJH/jlYcNGeu4eBqlDHOEBzfxAWg4QXInwUs
xKQhiLin8/gnMkwbRcq4WWqr5M3TWxkRm0CyK/77UfbxlrULLqJLfBATGr9k/8qA
KaEWRyEV+H8sndMN89T9Ri4Pv2YTXVCseETujBW7igXk+Abgu2fDJ+zb6Q4L2H5s
0VThJMx6H2mdiHAr1oLF9+9N57f6/3qbNJTxcDMN4KVPgIBSS8d52sbEbolMQkRm
XQ6UtmyWCxjhclL05QPQsOAxLsMMslOREjNx8e5u62Vm/ex+t9/g6eH1JTJkH2GP
Bdl/LcsnaW62C32o6Q1YRvs9KCaPxvw4yGrHsedOjRxIBeUauyMwi/mfBTKnHdBO
qtq2uTzU7Nom6iIloRCWEepHhfKKX+p2Vb54Qq9r0Dr8DaNOmZIeT4L9hycnMUYS
fD9oCxzsjZ2erB+i4od7ylLVXEmGaqttzFDxg9L/oFFmutVlqEr211jKiC8uUaCH
VPh5e3Qz6jc2GNt+ERc4ahWZTnYYT/rjMlUNR6NZGhpYyv3115Vi6Zet8IxxCJFe
usv5mgJiqe/7F8iQYerypMqPNP1iy4qJcZKw3WEMNsXgO9Yk6861YMr2uG5eBaai
QLK/IPuS8p2RpEFcsDLYCHrpVFZDqD6E56/MBTq/BNcYMZJW/RyUrIap4FaIn/G+
IHi3KEBYSzntmBCGuM+NhfLfv7vH6+yDf0qF4DYncQ1aGty1JyoTtHSikEg1Kn0Y
Q98A0HIRPeuFBks49/sIXW0GYaxvvFityDwltiZR0XsmRmwgx1Lx0eRDTfXZJTZh
Zcwkk5+/tLuTBMbbtDnJ4TjfGMO1m0kyIg8d9U20VfDiMK4KAsgWZAV6S8f1jeSD
qSob2aiSNNfNGM56yI2qigLL4DKFr1T31xZDb9EdquhaFrXJOIAKQc3389NbaS5F
S0sHw7aAdy0dlZsn4RtDWPyJ+UfIxi/mAbeT7TR9HQ45AWb7k61khdoDjFg0IMhT
n5nq3tz2LKej3KAKjxAFPARMRk/wz1vWbyRo1wAIh9LIsLlwWzeYMBMVHP36Ta+s
00B+ngc4UKnH/auPot/rcPyh56WCw5KXVboIBlby6yye/eOlos9BpiP9ZekxO/bJ
vtU2p61DjtOGLz4kj2TKK3l1AtMF5Zk6Y63Ce5M8MCOWqAY6mJDNM0ynMUw2hkp3
Q3z8v3BMKVLPYHR2aDU7Div+YnDemc7CkWkCsbTqtKehDwW4Yq08lx4iaeQcd89x
pbRxxeFY+PdM5hZ2hmlXqwIXcNRONjby+GGuY4BwfNjn5h4AAJe4MmuApBdw6fOK
Hh8LODZNnTLWZHgIC+5iDHrRXLYODt2/1l5MzwO9wm9duZUbuFv96Ku9CEpqHp7Z
YJr0gIjpu1TDh5z/PCqqvOpZBlfzwi1f3ih7TZNyF8zEn6G9Mxr6FZJJG4fpH+d5
1e0ZOuJ9d5PxjilxqdEbOyFtvQZZ78l+bPUxd5g5ihTgB/rZFSEAXBk+4ZSg3DAo
+JCuMPO5c4VtwsM+y2YvxQpW3OrvB6FWgTJhZtlDjJCUknfJ4pV+AoOW/jKqvUaD
zNA87JWoaWhnTKJ9eY6gWNOs8XKcRlk5mOyK1ZNZt6qBX6IbBVMLWjG/1N5CoHVY
kPtT7iHPn9I7yW6ykQ8HVQvWNnCBm0ecTRW7f09jqS4loe/IRhUqhmOizHh6qnlo
DamFDXnSgg4J4b3DWNZ2pqaSBP5/dLJJ3l+FQFTCWGqyXYZaai6ml220ph7a0kiB
SDQaRkim4IljjC3d2hGe3AKeSREJuoNoVRJ1sRv39Y3PpC9pOc0PLxH7g2YZJxTp
dFX7lN4hYU73daglmVqetdEnojAXmQfGW1zm3NvdeqBKyZZCRIbn6CSgBf4uL749
ji0Kpq9P4YvASgk7r0MBxfdFgIQdWxYzd+ol/x5kLA64O1MeQ1SaRrxNi7rAHYk7
Vl51+ds0Nz+2L6u3uV5QjVa3WwgGzqJt1jeFjAawnetstICSqFfatrUDeNVphHgs
0xl7ZqwPn5tT3QvAnl4mRMM5f61iIeouBhr61D2P16WprYLVlRyXsuwh6diQh2wE
1MtzZ67vgENs+ywoNH8AkfEENiG56erFWBLzdn1+0W2VgIVOoSjw5LT1XZfe7GmP
FkONg+66nXQJTmGyc/ovVcFFPqBGzPQZP+Sp7u1edOOFrx2F/DKkgDf3taqkYrtj
bCgLcuWe4mgUjVUDhgaSJEAguEVHGcj1BHQccKK9yYgVZqA1Yi1sxbHYKtYH75l1
+3tIasAmes/fbn6UCSm7Ir7Z8YpkEl6ABQfh6M1z1FrRwhrA0IjhGo8j4RRhp3Wo
JWfC6wxKj9sdU5ERlbCz/9DmrFpB9f7+lEzOlMaXcyz7f6DN+eUQfTtpOGsgBG7i
Yp38NzLjvrA9UZ9Z5bX01SgmfRtp7syvpfVHLgGewnyXN5aazrh/oYmAobAIRHZv
Y/YSYltKn/NnuzzeWaXkTG5x44FOcF2OMDDZ2L/q4Fsh4Hl+oberUotOHJcOBVaI
ujoUkmDa5IfxbUCvGld9G8cDTdPoXvaMhj4AuG5idx7gpUNrVShcHf0MWoWwN61S
GpKiE91CfuTISyi0HtHmNoWqODhjyooDLYqQMEB63tBThHMq8ars3MapACEi9KZJ
neF4q84eFcmOKRMdy/cGF9l84A+hahlbXwoH4dxfIlxOCoIAFfMkDYy4pfGELqwj
+16up5enaf6Kou2y6RIRFUWzf12oQNLaZUwC4ZmaI3Vp4DRnyALBF7myr6uhWUEJ
OHlyeznUHOwzZb5aiJ8lj/iv9+nWZlT7Y3EIohgDMtsj2UuIiENURf1X9hQ5ILfW
7NeYpH2pduxh2bPRT3ysrzioDLEHkaVkPGe1vYcEExboxMLc1MHpedZihnqlwdKP
gsHfPFHphmuzVP3Jldc6dVIhA716qWNfWzhQTrJZPGkf6Zfm0jFVLz2SDnpjrDxt
z/cFapYI4Lk6eJQl2Zg//yDNyesTb2l0yUUk1Od39gMHaOD1cHZlthFmSHJ1nauB
2MjlNV+sXhCSptcP8tt7iyMX8DrxALWnlj4VsFD0Lujf7+cn4ULWrkBr2I6ag5Lq
v75s+1QyP37Xc7J6ckf29JSfqisyys/dy7rsDsg+zkDNHst/jV9X/VymqiqEEcrY
v9BYfjRNC0LKAI6gxZ0RJeWO4t+OQ/0aQFMGtOSkc3FU2KDdCnKr87QB0kyTWAOx
2EE7RHBybuIRkkkvv+naz0hp515JwH3qlUtfzCRwGAXxqkbcVTrVZhoA8XAy6qAq
NT1cmnrU81kPlvVjRx1CqsM/dsV0a8bHjwTq+rEZsAcQcUDkVkKioaCdjmsQcNhq
P49fwtrNeuzwumIRABJ7teU6Xgkb/PIDwAQOSwAL+5aeURsFk4jaHKO7C0wfj/22
13RXEt1JI3zeBUagqQbM2+ScoB20mms0PTbVIzHc3dVu1vwkzzIrwX0C3fU/wEJa
pa8zJqseoZiQywVRlaT5CHxAJf+PS4JxExy11F0BJOxEcTUAlbrJ/ApJOFOwSmb3
ncIPM9tFWwOMI7+eMykG6EUQJ2WtR8K4mizFcXYp14nL9vMokpqZx1zQCds3cpdI
vJcX84AD24yeIQRCK6cAShec89/qgzTCKnodNBZk0m1lkgEZXHkuXvAKbbtqU6gT
1dbiC/4/04X7JIQkNl9tqg==
`protect END_PROTECTED
