`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTKnQdfpAyBXQtrDpmZSwIZvxnJgrFCtMaGdLL9HYwv/SdA4tThazETQcm8E7J6b
ZvdoMu2/AzDUF7Vb4QiW5qyi5T4lWMUzTm4ajnBD45Z4H2RK2S3Afdm7WdUrbhBK
gWsTv6PPAhWVfemktCnSN0qdQ4bumrI5QJyiIa66XMzRsNEzjLoW+Wk7UJ+J2h0p
5y96MjueLEM3pMX4EXr1r6Z+PblB8Gfg+Tf64FMwcNe3DAP/c3K+DaI4bmbsR4i9
ZcFx6+qDvg50i0K4tJlVUEMYfMBqN1gkhSo1KImiFuLETjKSy3sppWuv6gWl9mCJ
7Ku5YkaZovQBU8julRTKqLCy6i3+csVnum3aLNIOXUugCnML/gWNw98gj5DuGJ+D
5hANSHKGmqI7H1wtkXB/z18AULclgu51/KNSsq6oKNR7g1eohY5xCVdWMIMETNqV
fpUj5XgZyULWjMbuXLsjMwPeBPQzTsJik6kVTSBCXuPDJjWh2BvvhGQDVWVudZG6
3NAZcmz88MVUahgUgHJ4S+t78nDaI1diQekYqufGVOw3CUktWkrXUhU9JowG815g
ouLLYf6ECyfL95ICJRo38/owJH0D4piSwGgiKleSZ4TBmfQKXjlr9jkh5RLXxP0+
00r6Jtd1VMLROmZ7rIBW21L8LhDMD0VQPafWGe+Uf7j8MXH2Wu77XK7NfJZgFuuM
e6LjuAyEohFSOmRR5nMGrQlVy7pwX1iB5Eea2J5y45lnBWIUQgzYmaFQGYvsmDDX
xs+jn0a4AAr/1dioAGRKa7Y3sAqz7cOIqyf74Fcj1ke2rAAX3ccK+vAshZUS52mO
2ruUuGf/7HGUPcQusNZyF3sIS8xy2FxDdRYQottvamu0ZmErEllJdGcUME2MR3mi
m3JYY/A27ylz+fyRRN6wrvOrFyq/Fl1vrq7hVz+bs/aYGgf5dRaacUVpH39Pzvqy
Csr7HuEEPb15PvDazTk+xjW21++Lasf9kri2mktS+4VINJgLXmKdQj89iSIL6A3y
RoGFE/oRG2Il4Bff4nJekZuQzb4hVfJDvrCYhBay/NIQFteRcBpjkc9rauKHQwhV
uDhfQDaoqwH1W7iDDrOCLvaK8Se0aAVAaNgtv4j1qF7aqVj7YzFYoH2TMx6GzVNO
znYbTwdwfPR9UilWgwIE4VGnUUEFFJG7N7eijcYN7DbGF0rchy0NmW5v50sWySDd
5Ehk6LTTMQctfHZ+G2D1erpdm9ZqcmfHVV+mthKLrvWdY5cmzqlOsCjDxsAGi0bB
fdDF9pWiitBlU6qEnSeNLrii5x/ay/i06eiYT3Yd+iAImfp0nKJNWuz6tJUBi/qq
7nZrG9KGo9yJOs12Y+guH/1GXeG3Nik4G0nmqNiBnUWTlsjGMl7mnhgw5CoTVWOB
VOtad2PGijs9jmvVX3gJoi8gcGGKixp+dKewHmA1u6TsuOKdFHBdfeEWFHytmnbA
48pJ4WrlhQ1TUJ1Zi3f5jM6aGyF5O759y7YjVHSmfUIN0nT0bHeqT8pkeDo0/Y8X
FpiaUhxGAz0qCxvnhHRDxTi/6wnCv8CMd/IqfrlpDN6SevBHYxQRNiju2V18AM2R
oVuG+DreLIiGzznJb7TxBgZIf5tsK4Jq02JKMRAzWR+JoLVccPhowOxkpZ485t5Q
Fv7+FZgdzF4kVaPp4+hJ5ULXdzMNkR6s3VtSbo6fVQ37yQnE7SoQMOSxHceq9z2w
KmLwYAL506BA7Jhu6rJdTbEbCxsXYkgTRAbe8imTqVurRlWcn+9p32Idj9TIDs3i
DxTWn+u2KnidPJR6RSi/u9jM5lLrJinEwHVJtRn+MFC1CDcysOj1siD/QcTaP6bd
LzfvuwKf7tQI2UWczo0V7sxsiAbr3u0pTBFK4p+mRuZNmhKF0Prq0Y+Ts3W6SVJn
v2ruXW2GSvsJF3zh1D48oUfBpNGHh+iuahCBUBYoKuAp8XY2+oul2jbaquIqeuqt
80bUJUlIBf6dfeJyTLxsOKYRKdYMaL+3idUM0ZxehHTbMf92b4ox2EekfDxjzH85
t7B9H/JempBAnxSKmDMOgcmVJc42KpE9M7V9CIYoxyN6zbmcA1unK3A1cvBqamr5
pjJuujnROnFkW/N+ZczOcCHEMdn8IbfdjyPgr1AHAbbZ5vblJa7ygbpRlOuW5NTF
MVM/DjNN2Ppp8krearRITNMnVj9aRqlMLdrkbaJUJ3kd3Fymut3fF8VszSzpkZlV
bFLzO2lJFW6xsa3ScUJl+6UTEsbJ0vhSpeRstlvenvQ46Zp/UCfNlC6JauSehWYg
200tHNgVuiXn/IVEwzrbode1jYjZnohpqj9X9IgyHKdWWABpyxYuprc47Dl2beTl
Ew9h23vIbylLVGL7zvDx5Keb81VCNSxEno3LiAHG7V9/rE5te4wxpYBwc+5Z9dAd
1mPMFHZBfJZ/stUB5ZhOHWQ+MYIynPyuzVW3vyhmD0NF0fFfkJhBBZ3fxb84hDMx
imZMS9+fGU1wBGb2v5inv8HLWcbSIW1s/uSaLC+poCLDYGNsmHW/+UQ+7Iegkj0h
09o+W+dlJTjS5SwjonDrMoetVskmc5w5Wgqnd1cmwRMevjoxKtCC4jodrAuk88dK
hiNzEDH8f7uS+sYzaQKvMgKY8BkC94WjubbKNHQhWFICbbNgTzKx23HkP7oFfSdx
th81eC5ePiGIhWZnG/Bd0hBdaY3p1EjYHeCXUKTqvuGrk21INehwaPkYC5zLhxxZ
QYhlGwJjEc9hUW5dsf9Es8pbTNJWAKjKWjyewS+KvmHGMJp9Moejqy/imrNT2cFH
Rhd1kJkr5/HbsQl51UFoOMKU3VKu/55C63+4nNRTYIMy1bX4YADGkFbn7/vj4H22
JGpqRJauxTful+SOo9EGvFOAXUVnvRT/bNz9q9ilCXLpS3W6ucR7sLjZqr2dE7i0
gm2qdncrb/mtdbVyQaf+iAXCZQjXy1tm0fuI5rCi2xMemj+JXZ+jBCHJdhTX8Bt2
gLui/u22Zb0UVAzZn/yAjxgZP/e25Yv6ri9z0yY5ZZ8n1gsCaYuuk8SslTo+q+iE
CaGmJ0NpUQbmQ7mv4qYKAoIPFRA32vc3QqRqtoEmoKOmrBD4sfnXIZN4bzhWLFFs
opOILT4k4Ts/osvFK+nUb+jGaojzHNyWwtyqdERrEQjqTjWQlhW3ioKEb/+Y2t5M
Paki131VA8G/4591enhmabIIp87Ajai/RzHzpGlHQhEC+OzLla1fbG2HSSEDZ+Gv
pd3zi1fUmEt1plfs6vXyEir8UK0gRAK+fYHp1IjgOfHoyW9LJyBgQSFkoK1TU9Bp
h2aAPtdR3ici7s0yMlJ/C5Oo+2UICplIhQOKbebuIxVIiYb4GN20eLR35sFSFOPg
JSmNm/6ABl4v2Iv4SHVTPoaHIw1Gsj4meneEcoy/qEwaQq700eqoUdbWTbWNG1l/
YUwW58woY66KsJL0QsqKgjzUBEVRCPG8OMAJ+SHF4RNLZ9e/Osnnv2EHTgrTKEmb
9f8Kb06BmrAZdPe7t/clk2ak6d7WOvKO/1ovoAa+7XtJ8zIZWCxjoqI0Iis0msX9
+tQ2sOaqtE/Cj888L3OPS8iNsjsbnT4ofm7aZVETfqkyANoO2EfQ4LSW+zxIURRO
XwIY1J4XP6a9hQmeZVrT0T0Sxe59aZzz+ygpb5GnR1UuMRzSWrGolwgtiBlK/CWH
WW1iNSQbPrJkV8Ep1HEskA==
`protect END_PROTECTED
