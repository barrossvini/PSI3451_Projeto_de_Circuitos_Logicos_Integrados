`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gpgqvev92gJMmZJW3WM0dbv2AFMTzTjVCdZ/WeOxx2gmze6MiBJRWlE69oy+lTuq
5ntYJ60aTnI+B+puqTPco8WLzP2X9SJsSpCORLO35lJsUtnCf0N3sFXj4EDhkhaM
3XpT8HweUPqA05O6vSS+yePYFQZSqfSRMXWEt5/J5qTPUnpT9vnijOeTQ83Syi3Y
YaYj4r/ToCbVOgQn/ervzjmwZeGQtjdCssiLlHdYvDe3kSgeUpOGjXnqB97JUaH/
WDQffdqc0Hn+wx6DdB6PT2x8a2c1H4I6K/WVME/FDD7IiPiJ+Hohu8dlIO4ogvk4
Y7IiCy1w6/4EyxyeF41pdKDHrIwYXo6Jdmt5zq3A/RTXCZx9/Yh8iJNY/UMSOFJA
fCLQA7huBI5do1islADD/YkTiQejl9rVM6o/CPQXiY1sR7CjvIfLz/JO7e9s+fLi
Kn5JTFiodXomRa9pwoRyc3mAw4aTLXrUVRqRx6q56K1mGD9CGjlzpKndxsnS93vh
8b+biWFKTkaqTf72vOIaoyopfvK6iQICp3Un+unIU+PG7Ew1In5Eq4cwAg6Vfmre
oQgXOVBIBAnZV/uT/tkxEuA5USKKHcpO0xJL0zUfxSakM/wYayTHpv421abDz3Es
BafsZkUNmWU3R7u1oDEojYP31tLIOQH0MzusFH65wHewoXLWNyB4H4S62OUQVyOz
L05pjWNZXrWMeEMaKJed0GCy5DM80U7DnizAWzPyDhaWjp+uuiIq+HHZL10uscNf
D1q0bh/i2JNaELuaogU8ZATLekpEmLZrLze7k6UZ+rj/2dbdd/mNHm3FVP7d1x6y
c7ZuHsVHyvyc0S0/2+AdHGJSeCN0dr0jibOnLPLeFq5UTBRADp2m5NhN26CPPpmG
+IkL9SWMl+LyrpdESvsbUGWTyTqsuzWdh0dbWMxU+PGahoW5AA5agrRSnc+D8qG+
2AWMjI3e3Fy1R5TXhTYnY8Bss1Sl8ffbxmvyUY5+xRPmFzFNiDWmSlsAw1AY8+Ab
3Tra9cIeKBk0ehcwAe6db1wtMCrfGidxukvUpB8u8k7Ta1LrNNpuJKdIupwWEEBb
9WATRi5nt865fU0T4XYYPaZWZLtSTP00kQwSg8RL5LRMNn4yEuISnt6Y8+mtZ7Vu
0IaBNa/u21ejTFKXayATm75N+sMacJT/qkJXAxwsr3eRe8OJjiGL+q6hdcGZsR7q
`protect END_PROTECTED
