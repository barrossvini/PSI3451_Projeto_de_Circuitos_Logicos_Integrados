`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3J6YB0eibl+VS+sq8DV95XyF/QPvxXzqccDmi0wlUsMohIRZSH0FP7mJlHiUQ8P9
3Mrae2YmrUSr7w2BugqvG+GVq0zgLhM4dqEDIFjf1cnd/S7i5djPfezgLLWUErTX
9hHypGV51B+cjO9ZFA92k8GBVe9z4606boVeZak3PvNHvX3LiFVNPNMSISSX4SR8
qT+F/TT1m3pbpcsWlZsphVks086AhCRns0z1pTvbZ5OLpnYViOySUlRGYCZNG3F7
lmUJqJhwNzSFo3DiZqTEeCducln0t8y86UR9zH6SGBpm3npxO4ay/8gB+8tY9gNo
f0K92dMc54rv0SIP6W25e5eL/+KI1Cw+v06ZVwWIu0RHp50LSptt5eJANSp3F0ad
A4GIxiGXfR84qRJAh1amVurRV7tmpFXx5s3EwPsZpQgwIIwBPt4FRDS+cdMzLop0
S5zEIHGxlnAI5RTPe+eyoft5oVbpC1tHvLiSbCKH2I76YuCRiAZ2+a4B32jDfCT/
koekCIgpO+YsQh0A8t/pbZSvee8XrsIwc5V0rU0m4+799oO/iO3NBixDdD7TCohX
ZqbqEMFcKF5ChaWnpHwVXElQDYqrG1g48Q8rUqDIZn627K4ZHcdrblUOsC62y5w4
NLsC3+43M4m++EUIAi/gFP9SIIr6ifRlXKNqfS0wsrOoayYGp8u4Hisgl08cxIrO
GCKjxvjGoiuhuiiz+d+iF76wdkvSZpZWR+9aD9twg7pAZ+0n7uYcQD2FsO7/TDtW
gPcJ4cZXEKUcURnVlt3/lZEqKmqdsjD4Tuq7FftViCPPS3DfrKpYv94maZYVkezu
ZeqwRofHBk9UkiJOpz8iJD5MdqMUOQ2m/MBFCznVerrRbhoVUagwYPz3eCx/utn2
`protect END_PROTECTED
