`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RCcfM19G+YqH9x3wvKa+OqEWGlWjQJpdaJDvjyC9oibQxI7pDOGk9VGWHRg9WTHy
HlBw+RQgHw4ES6T7me0V4rgtBxu4ndTIAP5sG9mVIFaRRiJ4ICawKdla38tDih5e
GeB0MXL1q0SRc/ivBev6Ffi89cpzhooqL0njT+LLkTpfjQcdo6xzBHgzgYCOC0tQ
XaS7jBeZvC13V2JdUHQFwlQ/S2d0IScrs3hPTErCkOGXIfCgrcNDfYIaMIH+CiXa
KufaY/a1jpjW3QkFaIiAed8IFbdZCfc15LcQgzFeLcsKlSvTSogVUmKfYJ6PtOIQ
ovG2XCT/Ap8u9vqHwRQgv2FTEGAuqXFzGcW4kvrTuirFS/0qGgZyJtOErhvqhWyT
1V3PAVU1d25BZs69B9GFr5dmL8a0K74Ohg/vwdnMEXaRJnAsKbKQnZVb5nCXdr5g
92U/8lvXtChLCVdgjGzNZnmTbzcgPWDHw4RyAjC9o8YQyjeOFhyp5A/KmWg6LADP
+ywOXozI6BVkaiXjq1ajPyQyJPMDYk0RWan9sSF6LkJi6areMEClzMNtStBJmpDH
dlGepgNgfmVghgcDI19orIB5aHOLTTS3R0V95qst0gTMa4YO1Qa9A+vvo8XqPFe4
zs9cdiDCLNpuFVRTWIIAtqSdz16ebZ9URkcWdzi4iRyKjbzCRS5fXpZDRCGxmE8p
HatH5NH6GR8HWw0+owG03ogZYrDoahUWOh4Hk1bW2vPkJDsWhyROnhC7qxR/TY3P
fa3z6oFq6/foU8COewn4UUbD7qsZthvdvrf8/vn4xvkPwzfgxXebnp4xd5S4R6kI
LTcYIt1siEJ6gnPe+aCBwESPt+CAQfmXDFzsQ52q0qQeVt/Zfv7IudMFESH/HL2m
846Xw6A53p41UZecQINS+92xpNFsbCRDQQumfoMgz8kJjXdoykukHJ7XJOMM0hn+
DRRAPE2+V1rKl6GuBnE/pWURGOlCP/iFpCPGelXX0qLlEEXq3LamN70KIvyLVHKv
SyIgYucq+A42hDZoqNvEpEnAy5GZnQ/hDONuze4FbQ4E2QCcOOKzuh4EWvJiU3nV
sqHK57svFdHesTMElO0MT22KddVjik/fgxCJNPuiQdAHT0hLfmzDy/t2sTrpQ3hs
J4KbBcUZZcHGQRZFBFs1jy3fFw3FLnqzfBMdABs5aIRNCj6AO+EMOcTKr2kJ/FSe
w8niqxmeKnNw+j+Dnb9nuIr+/TsmWNZTKe6qybuf64JUUNcgpZ79DosMA+AAWzIi
8olbDajAi8iJMlWMQZ9KZI2sSr4MslV5VM97g8yGUVwCDA7RvOCcHFkQEEIYh9X5
kaXvoU7I4JSwHia1P9qeNJzdCA5wwGq2njmUNV8VXnWsTR1FwO8Y7XsBXBH7hT+W
v3T6uSn2ejc6bfs3yl6EkO8t6yCmDeiEp+XzifbW/epQjQITzH2GAz5uJAIE1T3/
sBKbGdmkghlOPHAMc/GsSg2H78B4hSiibbAzAvACeEcv7OsEjMEF5dAfRdyDt7a+
OcleA+2gkjXvQ5hxeWTvCQB0GLg1049maPWTbR8BhIV8+Y38iUgkeBr7WbLYQfqc
anezsivzF/SFRwbOFMSTPpN25gacOQ2cANXoP/elqSUGCl54aVEZnNcYc9ZXsPAy
ovxoSMHsQ0g57lWMEUrGmvk9RURwhoCVMBb49LH+5k+IGPYK/R3YW/PJ6MbxPYwH
z2TdYGdZTkUMm03eiu2jBGy/1a8K01RT2m5HXS/B9AoF9/1PNhN8aVZuAKXCohC/
xukQcAm9AXWH9nvfIlZ0BSe2GEMS0wkk0y87GurcXamJVzDiRzOHlOj7GDs1Ee2b
TG4hS+q+eLTB02alqtb/zcSWrF8YcJlOLMa4v/WBzDKq/ZPrMVqDmWpWofDVlNVO
VC/1mMHB6HT8TGAKj+5O/kZjTcUFTym5edBIM1VcGUl33TAkn1QGA2BKkMhCUU9Y
uF8kute9zEjpqbLIbP5IcLZ6Jhc+TQkhMH1S13GG65mO38Vb2XZk3qMjoTbt9yLD
nu7thw///afHFjJrGyFoWYB/ANdqkpNliKc+n2kZTue3v9haMkcRuvjLPjXQU50M
S3BjNt7wqOICnSX48aKPHuUKBj4E/t+XsYIEU0xKmzp6oZQslNj4eQc1Iw8TnIPf
Ix4f9sffz5UjG/fhp1sMWWRX52XvLD+chTraL/5+tKG4kSgdFyccWF1zEFrH16KA
voMc+JSWlcvMo1TrbVSncR1zlduPcyQ+RLG6kEwd+yS37RgF62wPowWsc11ANong
gS/Xlfv4qge/PKuDmFSezsXe7WdbpDgjmKEAMwqgew2HHSoLEPPVA3/GKAPSPVzV
n0vHhS/SHk8V5oniAk+j7o0i5Nq1Z0VZ0IPVmz7HDqhrIAVsTUz6Rcp7tJRd8JSV
lsU3ph2yEdcFtseqtfPU6yNv6neLRMFKzoLQhEGRqk2kXcOs2/aP9kHUFJWy4m+f
hqir0WPwUfEAKaoNQJCylga6lxA44L9heDjLxPuY6CBguoqR9IlgXBcSVEt2GvVr
a89WK+cv6+9NLwBG8GC6UkvLXiHUQRrrMgQeVhwWmVuKe64AJrJMdZQ+AMgjN/mY
GBviikF+zIeovWRpWsZfy2qcJLSBPl2jXfAaQ080fLrjBupqVnFVWbet6oDsORwG
cZgpAUXwqfJUhCOjN4kC6934UdbvNSPsBZPImjeWODvbokSnjxfvDNYK6De2Nlpg
xwFSalkq8X/d9FIh410zPyj0TQFFdTvWli2Smo7conuKjo9eGD0HkoWa9qRqxa91
4Xc15zjdmKd4cZaZaOCbMnBdXj+TvDfzhT/8CSj32V5Z7pSU7opxfMZ+KSsJDe13
DFjJLprWjVMzx/dxhL0Xvyuyqzev3uCnVW9UvCawW63wMTnwC6rvxpwCR5W+J7Yf
OSEfvtYKtAOT/O01maq2GTSRHL1tG/WZXIAIKsGtq5YDfn7iQGGl9iEz40Td9TPl
ttATCE7PmFSYrtdwCW8LtCJLRZm8yNLArW0Ot3GVT9lHl7qhZ1f101OuKrdpEmqv
+E8CZW/6tsi05PhDwyXbdW4fGHkyGLP2/MRublMNEr0SblQrDYrYLpnEjjtlAgve
FeQoz+uDcSF0AAtUNlcz0r+mJbEs9SmBT+TFD1U/Br8Cp2RSDTRcJd3NjNLCDvqt
3bFvmCTpgrEKV1y9lFawXS4DW2wKK1XTZDwrE6DM410CyXhfX8y5aON3+OqJIOZz
6zSHBDOnN2nWoqysGuxWe5pWpfJpSKEyT8+NkzMbUmMGt0u/Std3u7JfT793kvCM
Nx5g5J/yCobfDBZHRaryvgctHOFaknVqtYbu/Q1bvuFlytVvGLau+rjzS0ycvqoZ
FbOOqAdMb4tr5HWIQzz7TE54UgBZy+kTtRj4Ikc/hTb50oTb/Y2JCruDy9tdd6uL
Eku12rGyA3l8BC7YB6P42f4Th8lKlDMnm8pDgqppKVzI465IQCmRzYbN4XvlOYg/
2qlw7PfnEG5GBC5N2jLR8ZS2mOzkrTpoLYTKtoLsWwa634R/1GXqsejyMtcHQYNA
LgbxC7+itfl/tW1ITAxyispNG0F9pX/LLD1dc5caZZV2XDHXcyNlmJl5EfVcMdXe
KLhxvStz11BPHpauMaMZQ1Ma2hyZ+W+7mP81f+ZBiZx1oOjVuVSBUIwEPX0rj054
XnglhmZUpaHWCU0oFCyVccm32nphyKajbYllxc0HBpPC7Cqxv5/u4o5+ehB41M8V
jSs6C3cga8fa5lc6MSOKgXtOw6icbZx0Qh+2t2kMFvWRed5xMjxrbnTIJ+6qtskL
S12uhzid0OFFB2ea4WWdhXZoWkkNftHVGZv94yEGa5iHFxY0bdPPuw3eKUqhw7+G
VAwqrxv8dO6f0ye2ms+BByw30v8phOLlSKN4F4KnzZz3H6FOaPls6BL+uhHIQ1Wh
IW+YrG0W1fiUdhBMsIluSFGBg3eraQNPbjC+Icv01bx/Ae7KzlQC1FNqDFBh4JjU
eOgZS+KaZaheRRavsB0LLHmJfOpH4BHf48ZCVQXfoHC/DgvHjL15dlRQVBl2v/MK
d8a1EW6K9BTuF2NepsW/2uVCKkXmPyVm62Vk1Sz3bA8cajuAEtufS8fZ/BEZtEY2
qdTGDVkieJvntLfhWcOVaTW1nux3kTgyPnVmpuKw5mXTiLhVRR6UIWWuIfs7utt9
6aec0Zm6f1Am+FTuoNVfkMUlLcQG7mNLesuNIG9I+KFmY/wnyARiBgLIIDM1l4LH
UFLruLFUwq7I5VgHArHrMaV4U9v1FKjjJKktsyOhmfPvGEFxbTLWoCsYakNJiBal
rK1uZ79IJJtPCkI1nGxTpPUNSFMkuX8+BAihhkuF/uv/UWOoEtU4WamPukLMIal7
7Vk8ErLVwjnJyiVbvktLHr+x3TLWB/4J/Tpk13q/WcYlBuUeIvOpRdz3EtFKbBpD
EWJ0RquyjX6bK8oqcvupL1IFpCIEBRlT2c8AsuNZFZNAtfOc+dAceK6Ttfg6+QfG
UwaB2AC4Mnkrotg3qs5qQVXIyWg+LqqhvI3zL4QjN5nWxV4CJ3lqspYtjBqzWZ2r
p3kSeLoO7oUZIYwtBimfBcMl5/Qec+k9o7s54boTYGBjjT6SmqFIttZGKzoWru6u
IdKw0IFwfmFAk8R+EQ2ClmU7gmd44P2obNxHCeIy7E3Dus4cVEo6+igv7qRz4OxP
wRk0kpsQJOtfYHWJ9y7JnKYD3TsKEmrgnyw47Mz8T2m2ulCFWydAFGQPC+AqnYbp
1T1yhloeESr2U6ghw2vX3fRAOQvF0OSWFrmLyLBhq4/9IZBRQkM4/akwhmlNUEpS
mU4PaH4ESpO9MSYdPf8H/Y7J1ENZcBF9GXBkzf26x6/3amHeNc4+SoI2pHFp0AJT
QZOIeFGJDaRFE7YOnSmrDKA9xM+ZX8zNBicHPmHw1lPoi1CuYB6pRDKseWLjNRyo
lPUwm3VQUbiPwResv7xAFdht3sUl6K15WX1dGCE/UmuKuHwltKv4NrbuZjYvfPmR
z1bDKHfufS2ORztTzGui9ub7iLLBn6I+qI38dGJKUprhg/w/YHE+BerbLU1ESCRd
HDbprw1nd3iiIw5d/SqoQf0QHldSZfYy2CU3yllLQ1bQ3RTAv7APctXBwYKnZkad
lMpqw42AM9YFbSEIeGnvw5T4CmDAHhhFpbVN59WWLx9dOmBsu3jYi5Z/lUJttGc8
KD5/Btw6rRD2EEwj9Nmefjz70gqUIhoXiBIL9yfrL8nQ0+D/tYqG6TW3StcrQvbx
uqvmFswwMQQ1O4snVaeApKf8ApmfPCyxgskcttrTlrIh6uD9z0nTYNO9bOKFKd0H
zDlPT1vRs8BzeU+uhohusshPRyHnfBqB8MK3iIwGRs2hDm9fdnjRb+m6ZNaUl4dj
Fnj4wM2EVCiR8xS69VJy7UK3IRedEXFYZr/HMUEFhTc4xVPGE1SU/oO42Yk6ge3Q
Fs5MV44t/5G2IG3QvtksiRy3eHh49ra21m9FEotXIrMHmSrDUkLGc0+JkcedOni/
SEITg8YJJJkaTRW0k91iK+xtXDE/kKn42682CG62kExVhonCb3KnO3+mspVesNCO
3ngAjwBpTUwDC0dHRD8/oLjv333AlRiEPkVkXqKpUZFAMzvBmT59m/MYzfaNzOVa
0GDRDjtBhaA+c6s17KlYuyfRwye+fuE2HF2yZxgXztq4+sNz2jQrHnkzSqjhR78+
Nrga6k4pOGc7aCa3TfRuAMsM1Tg5AsV876P7LHatedxEIxWzPfjy09s4WMyIwVlI
OH2li9JjOOQHUiTMIQp5YsFPHiveVD5pZXefvNnkr2/mYmINH9kwyQyqdlbquGBL
jP/sVkNDblVm3kFs4U5FVo/wupveYicQINiyHl9Li/vsEJUs5pRyotUovv099Arb
VrTxKfLBdcDq8rQ9wl5eqFyAudys2awG/qKdWfL8HWvgEcFOO6BquCUhhKXCcagl
7uV4neDWiShSJPqgCrLLqqvpZwrlPQI4bA87XIKinDxJdyc25SNdaQmN6+lWO9xO
lkEyWV4mUnTBM8QdwtooL/4PtA9DHhRakYpFgEsvTFmgs+Bmx92+8yyTLyKCw3Fu
e0QXeYTKyncLSaWX/sOxcQqjxjy4Ob2znCluX/ouvmRq/oH6+CRqK2vMfy0grUMS
7EgGSrw5S3wbpPN//WsWxutU0+kBxufDrQnOjkXsLX8/BkmS6M/XR/ZJEp4A4V+6
x+L8g53ZWckxxXBVGezzV7cPpDCePIZ1+PYmx8KyL7AqHHo2kBgnX62nHPx/g+SF
ey96gMUyewFvfJGyQO7C2afAyPgxVdpp5HGW53MK/kcULHE0glFK1AKH7a+ncEch
ih4GSAul18IoVYNlX9c8lOXgEPWncRY9COOPu9frgT39Y6PRplBZmmz0xJxAgwoZ
IbuMoWQ8Oh8N11hqgfF59MKfLd5/2CVfdWiNph0m4IeWuhLcs48Rt41xu1zmsWjs
yIysT7G3dbG8CAmSLtAZYYQykQm2gPc4jwpyTsyNXCCvRDSjVtBisEkJfNhnTAhL
BDlMFZenn61DFnyt9LF8Q4Me+W8u8SaPNCnyD8NbNXxBt3osE9AvsLP/IyRKZYil
tBs+3NJcr6haePR0dQinnOQqlNKZlPm3B1hlmeODcAJ9Al1cQZdXvM/y55U4A3NM
hTxa0kTXAPqKef2snxaIl5VxwqFLVwHE1EhNV/P6KiJdWZWPsrWNraw7jP0yqvP2
3vOB9oSL8fU5skTgwrEscYJcsnqL8rlidKYjvwdoFe6JIPhyYh0pydaiEYdV7jxl
hxPrHBxcLLLSc81pZvhqt2PrwyhoOI+SDQDszIqT0sqd3tuYYmSoIClrqqCUbS+N
qibX4V6SE7tk1Z1AxDf17FL4KquDBKkIYxOtEiHFR7tm9OvuKRCx/9hUekUWVnVg
GLJdGPhQflDiydOmppQ3Ys279uzm0Gxz0CT+N5twVq24zTSSzithjHwO8LNgaKr2
NwDS+4LGVizvmz/cZVJbqqR8CbzLIxRHipFUK6dDStkzxNb+aDUEVVy9QtA0x+tQ
bgTSVewmSfwbcbhgiQ6eW79ac4eui4EYS5r9pWhawAflKYV6OI28CIHg+eZXDTRJ
rRrRNE3IL68cR+JPHlPlG/eVAy6dJn3jOLuWLbJllnjBCtE7w1iUZJ5fB/OxtStN
FDJEguxPAMIiTNqYG9SJyZy/BUfI4D0QNufcYXAPw6+d54jTptHoxZIdsnXK/Umm
0z9bAP99/mUKpc4mASHDIXlwzwIe7jkuXuduoWMokGBQwqs+E+DXRwl3nPYIwwsp
c6CxMyD8gi7iuaVEbGZC+v3gbKaVVtKrlpAPFZka9Yl/BKQgNI+QqZi7BR2sHU1p
7T4N3Bxq4WJ8x4uBsR6pXll9nbQTDKt8jQ0uURLhpMT9cuBwO2xAY0JKnnZTxFX2
1GUulbLQv6jv2GiZEF24gAxrrgqO2thDVRKOOElT/8YvUKshJJ8cEdazrVlZQ5OA
UaMXsaf2/PaClwxEJ9AnHjBaUPL1U/Uql756qhpPuF18owjfNGphvDMLNh4mpLox
9K7A4fwX1lGtXRUPdSoC4UDAoCXC0afutDRF31mCNMPVUaoisbC+zKvMDOP0tS/k
VpT86E1lNooM7nZEpboSMNGYZL9euWrSjlkiIzimtgRzS2XI/FyUXR9HaXWC/bgy
fMv6xJYdFAfRixJroAqvlYtHwY7DDU76A2kTY0D7OmZSkTofqOgW2gqr8i+783ab
QH8DUYCHX9TJZBUPNHlLvKfPBs7dU0TZ5jtiFMCWwFHHaDoTyJJmah/SpmcP7tzD
RppDkPfjjQ8HPRI+l9BaMnTQ/XIo1/gHEMqtjOAb/8pmaiqTspGXt/YZx5hvswXz
clfbv0+1BWI68UGc2Im6kSEq2ifo+DvIbMx7qgRh5CT2eyGeybRPxfD2gu3jHTVT
Q4LJxr7suS7NZvB65ik66twAsV2ROiuTViawd5JE4EwSWhwuRDnL4uXPbGyLO+cb
/5O6k3lOC7zqV7Ws1bIdNTjNdqJZ9ngvXSKScNudetjhYaJa7QCXUbF82MTk5iIv
L07Up1aOACs+Jv6t9552lLbfVud9yD8SegwsS/IP396CpKMKKnMfKUq3qivNaXjK
sNIxckAZl8RmnaytHQ+fFwMAY+HL1QVm/exFP/gg3yYDk+uM6kx1r7BTblYXVH5U
pR3WYGgy5Ca2kTDV6Dx1PWKfRmImSwiTCLsKWqiq1zlv3uaKxnZI43VJKs2pC9v9
iOK21sz1qPthpeklumoorOlD6udbrLeF4uRsYK5gjRLreM2eox8+wLLD883+wOit
efgDNyVJjhZsHI1cZZ0vIYj15AJA3waTQMqEc2EregoZF0xoeoPIvGRLetP/Lxzh
gVt0ooSrmfKE5eY7Ahl6J+sEBjQtVGqwu68k2i9Uww+u+pKL/vs2n5yd/RENVhfy
18A6bosXUlKC2trggvlex2H6ZMciE0vAZ3W1RCxYNfPiZTupEKBUPbi5+Q4moU7/
vsN0wsJxUtpcCvzOXZRBGmGT/jEk7zmSdmCAhFsNU6VO+HvaQQB//16AKb0ZtBad
uEzDTK2Z5VJ8WN+dN7IuXTCwwfPM/pFxSsRBpK0E2Rvh9I1SEJab4lKnPerE0TBk
HYaPa1IKmnc/YUYi3J7gZzGszchPiJKocS4bGI79WdDUCnpJQ17gEv+1DwC89xWx
aB7+WJM2/EDXF/EHpOTnnJKYcPN/tkRP0wUqbE2Z/pqkrXWAchxALQMwtkTk3hJI
w41vbjPAX+oRTN7g2z8xEMgHslBYYzj/VQE+XPh9NeZ6mLgxDNF7FVvzd7Rgx+A3
yQv8iTlQJzlzL3AXeNvB0F9clxdeIO5IOtdokjb2SjB+1hpbyEVDdIZNjvTv8dCv
5J39mfOwuJnekhY4E9RTDqe2g085Z/qw+ZDOuuO44cHyHTYEVmq3lrgvUjW2BCBc
PtF5Ja8leFT/noVwHY/kLVcUygeBbb/bifVEEBJZefs5Pc815xd+QgxESHeGGxmG
WPMCCBof7ozWL37v4Xzv50kDrPtIA0tMdhXKFZrTcOUfBdMI803h3bSrGNa81urF
OAVVPr0B8w0KiAM4yocw/Uh1z7jtqYT8wDM6PrFYW+MQVgQGx2kAC4vhVGvG8kdC
ORb6j7i4hmbotzebgD8QijdSq6v+J2MdqHchcT/gIAyb3xXRz+CAo3ZwhOo/cyDi
yRI46Am3m/lSra0o9EA0zKavbSki2hbVQJ8ZoO0UHTwaRLnA91Rug3Op6w772TW3
7LH50yjtxQflWulixwp0tF6GrvCLc0cx6en9UIg50nFj16ump49QTPj8QzMUlC1T
eT0N8gpwlA/5KYAqLS64yPApcMMLVkYkZ6CJfp5/aGypslfuRvBTOjcumsEXB82L
VA3LF9FhtvDOCAEHbGjElaIzl5k6n5unSY4W8QVF6EGhLSHuSiVq4YuHExZgItfZ
0dBfmxTYEb64GalBAkfj1iEHZ56h0nuO76nTTtmMAk+eqyjHwCI5MqS1FeCdSkP3
pzPhnfyXZPTs1zAgFiU9atR69PDYsJilxrs3yI4E46R5ISVJkUdP//ceO3ZAOO/N
y1cdEkcsU7jsfdfjSv9b/fT/0UklJaxXc+CtyHdRhRjVgZzcG5c8JBhpVT1t5nDV
2Un3HnHXwtd/a8aS7yql7TkKEdlVEL7QYE4yfBsbt93T5iN9ImLUaXbBqGvSQwwu
GA32nSkjSheEBV0FlcN28W2xo7dIKFGMQa/N1ZaY0HQmTD59AptGjS9SZKmefFXH
njjiLJTYBtTFTDkshjj7W4GlsYT31T/RUr8pnUE0cVEC8vN9P6KCEiIh+fyldPwC
uqifH+HPNzEMs5RyS7EpqGdZkyIAVl4G3H+z0mQ5KIiuFpmLYhoKRzOVPwFVc59+
E/ixA3v0Lha1ya/DzbGkVQ97A5ZpdGpsr1p7SxCNDp0krEswVAtsJmdq3cXxZuaN
58RZnwOVSu+cgMh+NKZL0+i6ySKXvtEyRbI8U1sFZsP4HTgyyDjP/lXmcwo59OA3
8r4QJxmipbzN0+xxsVwKQ66dEn+IyNEO1WXPlmbUmYKx9T5ZHjKrNvrVl7jllMd1
SI6jgCsK3aJcjYkW0+qUVnJwI8l2IqlwY5YkmQK8SSe0yokQDtD4IZtrqnxqjtfu
J9qSRuATtOrDx8BeK+u4egiGOuBBHS3eGAJNKAR/TlpsZ2ZyuFuwCeW1HZMC4uh4
ON9vSDsLUibp/9KlnSG4llrEBIl+E2nRhSRxuOyFeJBeOrSiIUbcp+WkBOVbrRrY
ZMaRV/DDzbzYXRzrjIyw93FVH5kgFwjtQC7plA0bigQMOXvRlj72Iuu9n8IX22Wv
nwht9GO3/Iy4SIwWv9yPCMy+tLUd1yx14iIUX3X+7/yXFcf9+JpFXHjsibp16Vq4
8QlMUCiGBl3a8BBnO0EoLfYnZajCThVkpKQW6DoUJgM4paRxjSvdGHoRhZCCt1Ws
qMwglRrfmVqIs4Mt+q5BUfTe4/DtdPwhhnSW4rhBCoq47T/KSnpY6UzMJWIo/j0Y
jYiMJPAf+xHJ5ChNhcQOiMe1vnJXxyoTOwEYf3MbZcEMls+Dy+83kesdveIRPxHg
oWmFbSCH/HpiF7Lgwl/l7AEKGFqnNBb2YNmd8RM8oDny9iNytxEcV9y5PnwvISom
HBq2HeJyNDBFELAE4ngXFtU8mqinGHVKAO7yQmyHG5W6ktTBrqbqCAtuJJa2UlfQ
Ct0s4vh1myAVoTC+K28nQ1y4srvPa7d46/CxMKvGnof0X4/KvCwAKWMTdGB4Educ
9GGtcwKtG7W2vSk9jkJulmqV6DzLfDyamklhO/5aH97rRV/BK4qu+SxEpA/+Dwr3
IGXogso31zbQZaBVh5aYjNLFVheW+lhFEvwu7J+7OcFrBZer0YKcM428pfOWiL7k
FgBPN5D8LvwPxo844KUfAXCn4varFMZuCWbxXoxWBMrsp/6KJ/gDN8s0DLeem9C/
z8U8qXkMkmGI9QbEe3yHG1gVVXsWvWVdHpYfD0AcZMRsn0ORuyRJZAc8EiSDM8jA
PrFHr+t2NERDsDDER40dQ3g9iwJ7dLLwMTt8srljSkPKNag8qSz0SmSRvpjifKZq
1EgyBZdexJ16ptm2PP93LEhrLzp4nUkJrI/ULz6liwAbdhfx3PgsUMeEQQGtKh1d
mn6l+T0LsPmidzEBvmaWCYBufP3PJNDkJ5HzBMiSf93fqoJ8SRRerwFgOuQnawUt
qXxHP2EFKIN4/quimOem7GgFA23U5SQQ+Ctqs+HmNIcDwsPUwo4FRhr5zOPNLAzt
Z7ponh2UxfTkeAo1y0fA9qi68bsYXZKT7W1JBXiBANFabanPY99KEigiry1a/T9h
ZU4uwVRDOvmMSzRp4x76eG3vv1VZUqORhYrnSoBs4P+l94ReznQI29bx2GvcIZaE
bsaqyct+f4C/v6Rp1kC8wDMm/F5tKl92XJJPEdJobtW9jDAsR3/qzFDU7byQL5DZ
9um/eiAnttLGMszUP+7aKx4Psq5T4ObX/8TeoSWiUTI+YGRVw4CQs6mIx1UK9AMa
CFLiOWTxdFROL4KzSYpC5yYT5iIaZk4PQHGhDiO6d8hXApKFuAudq5JM5b/MlF1T
Yxd8GhISZa+E4iA48mSrZNHKatNqCouRCHfeW4yth7BiMRSs7C0j6uvrXY6syC9b
XC8WUxRI8rq0iMqDAd62jkhm/7LhvGOZr2WXj68qPIeUscSyGJumw/3rEVzfUw6f
O1zsIYf7Z7P9HjkidmeVMTMMu4901CF7aAqzjEjjXzza4RFX6dpCpo/DaQuFsNCq
ELBgAL/ZjnerahcMFMeKZzM8LMCdRNxfwfWeI8GB6NvU1A4NIPzjNcjPNgSW1oIB
+S+HonYFDAWIHhddZsPugmEAEPebMS/p8x0rszhnD8LYUiYzHeOPPxuHqjcXWXCd
0cA6rxzqemiXqMZc59Natt9dQBau+7AVHxo4AjvccMjABudd8R5pGrBMu8TtFE3I
ZQbPe5qCK0Paq6ivXHpsFHD/c4fp/zadvMnofddy9dQR0hmNJDVo7vsZmdzBVS2I
5pXinsjszwGeW5PgrDY4joHOJc908mItB/6zeoO9PDK7jpMcLdKennQMF3IzScBE
YKfKCclbN6QSAnR+E8ipdLvwzyGTST8mtJFbVvBJ8vu1ffpNeYPk+GqSrYD1B5vG
qh2hVqEWbrs8Dgj8MiANFdUlFW6Cll0JeSCMPgoj08wJw4K4PMzfqfwPYIJqQqRE
YC4PpPL1BEtVNOjy9ic5zQdpifjAUE3JhJbEZXYlCAU38Ix2dov/v1ltGn/T90Z0
wqjIeFJtg2piyC28lY/WaKZZTXVp7O7aAfhAjqKFyzYKUeTCcvipmgXZ3/G0XjL9
M6tMCX2pt/0YhBka7lk45S0IzM4qbOncrrAu6tq+3u0CbkAISX1JU8YZyhlTBEkx
55WN734Vfm/E3pQHUR0Yg0JfeYn41F8OMsA5ikB1xZ9XZOU6MZuJpOBraPCA3qPw
Cz0vrVNu9Ke889zAZdYa1pZkyS9DJ2v3mlnqu6qKzr3T8Zu1yNwOrR0Ygl0z5Y80
OvvIAoeEyYBv7APqoDCra3Ve35qBDbYA5gErthzfUTL9/c3QGNQuXM4EEJkybl5B
LvfZvYhYFSgC6dMcss3xgVO/vUZpEYEJuyawAr5RZuBLGvA4X4Zkx+WL7biz0I59
DwMjFMjKssPsOSaz7xn9/Ol7yTXUGJcNRU5J5xodYfVt69uM5wBsFgIUc/iwmQdx
FCkMEdu3rqjQovVoe40HHR+WdrAfulwb7QJqvA3SHDPyDZR0fq+8DrdpWUDGIU9F
X5MpOL+0BaNgQyMbIEIjkRtCOlvLhLib2ZehyBZMBRUoHyzl8O+AiOGNF7Ryc2Kz
OWpjf208JT632S4MiHcFYFm3bFOSJqf+e3H1FUHUZhxi/g2r7iNlgjcf8Vne42mq
0QLsjWzEH98nVMThtEeHUZ9ePUhb2kzOevP2u+tmWxG2K017UxGR4DcAEoBz5/Ui
jHx9g/9BS7jVp2Q3vE+EtzziIklSWdRGg5YU1zb5/P1Up8tTCfnCDxcG67yVfPh8
5DcgUrnffKGNB+/62WGmu9EEndLImgmrQReiiOplXA/fVBNYXWkEShF6mDYjJEv+
CbHSMT9tHhQoyCP9M5FZZb8E7DMgzlo4wJw7ULyFxOvKxn7tiz238I2Xz3QTiAK8
O7PhWV3FcBff0bqQj1HeWw==
`protect END_PROTECTED
