`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zXiksrUILlrFGw1HiTVUUAIVhLP5i+V6CKsC5c9rlowMW2EpUKlmV+5KBtRzCtYP
5Wrjl/o900/MwvLMiY88zsNvBMfliBtEuQr33zELTe3iAVtczX405GWYuycCWzic
wlpZeQFOYWbLBZE4G6awbhpSTZIevSwCwY9G7EdNd2k3n6cJkl+xSre0I+3X/qse
LrrT4GrJOaZM5ttM5d6Ip/qjh67IlXn/284FXrvMJYbLS4R4NAOFhhRs0NhF8koy
5Y5BSOPIg5MEAjFMpWp6PLzG9F+zCJxo8ybIxvE56QkrdEVyjh5LeT8shXcjuWsn
D/fYKsFYZWrV0KDc2siv6JI1eKwy4zKXnPMrQIW0BNgHm0XM1ig+MT6VMYN7V3gw
XfBPeaAEHiM7cCojiMqwXGxBzViu6LWfHgGFMcK/LG6cdRsJOE5GAnZ5lohGQWif
6sXvqKMeeoJQIiYJKOUdFA//9CLR70kYKYUwLjSIe0px7OYr8kkTK6TdxyZjRNPI
ieiKylr4XUUp1D7qyB/fIi4gfR0gpLFis2omA3tp/wLsm6iOBjRsNQcBY726Mymq
iktTxqk1PZOd6wUESg5w7hE5JCAtJidkMzgaAz/4teQuMCaIdnc/0RkAnAevUIgb
L7Z/0WdGLOFAATkPMKXJ2CXSu4vp22JNIXYmouzp3Zfm5tkAs9wkYEUNXv7inx03
rWubr+oHQ7hzW5PPIrp2HS6z9orLZVLILNf7nvaw3d7Y8FsDMCLVfWbQVxmIvcIr
3SFPgOg7oxZowb1ciNdZIMS9GVUHV4sXK4geJaAsmsd8PNv0QdEcvxM9otEAWZB4
TExPzhtC2WGvg74ZyTR+nK2Y2hoE3rQWYegy7WKMO0+/h/aQrv0OngGvXlRKs/Up
zZfhZ/u7KktBFcbASS3OHwNBxHTqBSOm2mwytg8KfNpvifHaIrEIVeuuzMmifdRO
1o9McVIa3Snlf8HPqOaKJPzJbuHdwI9+NtvUuWDPxQL0QKkE5A9x1CZQ0gvbjYQF
jzpqdy5PlpX86hxv0y2mO3uvnMKQhJT0AUpHWbb/Fk5rovXls99IAn5URma2kDEp
Ly46SMPatTKvfr2ckFjUzRvjbPh9DrzQT7urZk3Xc/1110d13APxfItErFUR6dsP
xZbQZU8Qjc/9TaWGvofNONprCfJwxm/bLp9WwlOrGM5TYgKn8OqunZdYLhmQQ0LV
JAZ+NksDo6s1+WRQ7oNyQlYMzi61cdHh8nG/q6kwiFv/aI8BThWHsIp42dhwVNoY
vbOWeJg6SxBQrLwNzhwPTgS5xsMbWkv6kycmRWjD3NU/Gdwch5bx+LtGYay5i2hp
L/AgQIhjnMvMYwHJ0L+YzKPEaYxSqa9nru6hgm/5RbG7Kv27tfHXWa75depMDheK
LUhEz3cmchFLzQakwjejkM+EYhUFNVM7bx2M1bkFg5sduuvyRNyt8t0DZmlHrBal
QCkjVYUIUjvGWyzya5XYS1jZtdsKySj88H4nvI+OKVIIWfhtMYYoE6WLItL7EfSR
FEC8Fduo1LoN1lYsDwa4tZKZvpeN2MT8l6EgJ/kG24Ne/HyjUvxaHQYy3A/OHWaV
2aU2GDxXgXQBoxF/w8duyZWeyMIcyGQ9gyQMFIfVYEoeTyW3BLKkRrBEr+4xlNGs
BpT+73VVhCGJQxWLNosFrpEu/icFZBfBbIgTvzhS+JvxUElG3XeK5CCCKyeg3G8l
7VJeXvlBUpAKqf8NWvfjPhSjUROaLS0uVvCR4zVaiPLRCeJkZlHCJxh5KEy7+f6r
K+Y24hwHAvZabF9KnEwTPDCXtth4i/lTfo0qUwpVDn5DoCp2+OeayDtKU5Llkfhr
3rHfVjijs5rF/rdNc+Q1Z+ixBm+z8P7dA+uichwx5RPcKfw0DEi0wuSeBDYaInPA
8uqXrIFXPXblyqPcf5Nwev4MTOuBGAsabkOQ57Ke4l8Etv3k0QENlpMVgHcz3g6D
z65gfTsQ851YhjFy3oCQpAp38iWAhc00MSw9WhEaXRztJXDjKxwRxGmOkbp/uQNN
Dg1GTZB+OjSX4oa9u4CmWUiw/ZQUXsVHHs/GS0IducBEabhu+xokJs7eHf1aZlJj
qzhyM1bytinA4R9uqDPQGsD/6IJ7N8agsg3jEUZWqbu/L2xyczIQQsR96DZOecLq
MEEd6QeNNzONNyp9M8UXGTNzoeX1eZGu6AEMJIQhZfLAsQXNg4JZfs4UuAF04+qK
nocoqwmBO0XjUN72Uswf5upCxb8iL6FfbuumlChqf9xPRaBJL00Ptaq30AU2LwHI
GVq8x+k9esrfD7wE55e+Gu0BdC3l2V+TrdxpnrfR5JZ9KuECgawhgXitLdI5X5SV
1rP+2+bfgzSe+mLEpOcMr29tvdl/NUEQAc4bMROTn0sqv75Zmv5zpSjyUAYbKyaD
Rxx3VQCjTEruM9JXRtL8MpyRAV8Mjsz7YxkLGmWjlhWyRssuj04fOLnu24nJKIBR
eDsZTRw/Yh+m5wM6AozwW5Xb6+qjNIDV+N/ttjgNmTa6oS4WbDVju9AVhVY/HbvZ
lwVV9VS2BQlJj5S7lasg0JR7fvXLvrM04T0n0PnsJLcogfZuFtJU1V7BySon67/Q
vLZNwl2GXOaaib4+U3y9Y8Qv/txl43yAreU0WXkll88zPRyjWZ7iqrxNJaTnAQhd
8nzvGET7TAUBsKmPco7TYAP3F02x2wFDoB9RhqwSOCHNszWbha7WPstBfAgKqD3c
mSzTOUGUdhDQpB+HEwRCVaC54r0JlHAWuB+6IP5l9T+oiPiZaSPvf+vlw58TD6a5
GS6NQhsiMqqm37x8leRwPhMbCvh9K8PNS5KLKmEMM5kecN8V+WnjhLds0ha0G52D
94vb89rRAckt8H7inwvCG5NlUCAFoYBS38ds0hXhZJqUzo80vIivMLn0bK3DmTCJ
R38fQMwpzM0ciNQHoGfCBlbPVwJ5p8opr0gsXVJn+mWFcFwrb1YwK9lbsxVfgeaK
d6+cW4cMk+Se6iezlL3dY4zvq+qBSKiB6/nBYDWHoJYhGy4ffKRYu3Fn1yVjSokw
jJ3frMGocv58CcmBGt9YpQGNv3rGcVdGw9IvKVhSpvWFeC5lZuEwjTZnlPXfjVnn
RWb1G578VF6TAPShhRJliYK8yyHKf5J7sE3dT5IkZW7jRO04XZl5VPAG1iuvIz8e
QIT051N+1WnialW+immJunjmR20u2oAVY1B5fZSy+f5naBJ9gQhCTgrKJhVv60eK
3W5qLKZkyTIBoBcKGU80v6fhfdJ3CXk+l+fCccGT6LE4N0Bfb/UbLSY/nML0+Xpk
UEZco3siLw9VvyG7AxrcA095SIsa1mHXJqfJC9B5KzCVWG6ZkQ/Quehc0AKSZGdj
gbVyGHS0CCPqp5Hgu0WBGP5urnxKvxyJntAEFZpi/P5EZV0swnr18BdjUwEwoC9K
OnSOOcW28n9o5cH2yTdvTxzSY6UofrVxJux516Mvu3Ifvzc3Qd9BfW07X0sOVFpb
5hikRocncfbkVoEUAM46/0W+QU5DJG55VXbJxoW4HyMWJ5Ms0H1tJDlyA7+EA9L2
aKJq+U45UshT7rsvU/iAD/VANl8D4lAZAslNUOVjkZ6rw0OgJnbtH9NGJTj48tyc
CUaK5oCNWUJoIXLIn84+C8YPXJHJpt/ga6D2aFvMbu1iJ8PS2GXEDtSUBhs6l5Ee
C7OKQfzw2Opg37Hn5zj1tR5W3uxTuDtDwqbCYD1hPzrlnjAkrw8fSgG4Wx3FrRIo
oBe5XDuFdlqs/MlDPQWSv8omnkvf09mqWivg2DIRqqhZg4wH7i2Q4HmJ39OaXXSi
CfPxlzHJj2btlyY17AU0GDGjL+hsndfZ/CwQ+mr8zM3rj4w6+v0Zug8tlLCM6Huy
xl1bT1fQbaRIQJgyI0XeX70cT85Jr+8JDH/oS0E1LZZjjODkLF4tJK7P8M/2r4WT
6CqRqaX3fMmt+49MP4eTUkCqjcSouDHvAaTjinpf9G+abnLQ56GcMXc24JL6HUud
X5n+pHUgaBwm1LzR9WSvwMd8yzR7zgvVwB3ib3fWckBOLRhenlvpb/OviyBpblkY
q6eokf4xA09UZ2JB8j3ORlYL2Yxe8BGJ0Uu1vkaIeq44byYxSRvLzpMpGHE+/OVO
78C5VR0zVjTKCyHN/BplsjSLpv2kK9BkU1bSS8mI2o+Q9p3ucHXQR45M3UOTMHhv
VCe2covrt0a0yy3Af5cJPpuj/ZSIYpEsqJtI8HFujz5EAFvraVcY1FjVDXslIJdL
E90w3/q2L+tIEXWWxap1RPh8Chy0tUgOY38obwKdKg2jNzrlRORHvJ9af/cuLbl4
/uyZJ4oeJBQhWkS94GuCv576vVGg+Z5bsLT4Uy+YMDvpcpiy7aNVgKYcb1AqsGt2
wo+nGcsbtux7D8Ay2TJvL9/v7VkY+R1owkM7GpAYnGCEIHtr6aSVYX3M7rSXG5pC
panHRkxE66Js877ufFM5m0gQ9O1bhKnM2VqFnNgTRm73AopWlmkTgF+m+kO7XZW5
s8EeQ4pObOQkbCn5dRtuBZ7SlGP6b6BhdOkz3EC5Fnk4bqLwSllMBg8m6kJeW+21
qqXYBn062IUjlpckHcbsx7vLY7j/KLqGiAoskjTar0CNBDXBMfA2JfVLhWtdgbnL
53iQvEgLCFjhFiu/qG3zeFjldFHwtrtXUwoEA/MBfsp16AWZizcLxDWot3qRJW5r
QwfBSGDpgkFe/xhLBKl865DxJEqB9Yx/DIPGYgX5kGSNr3Ocnqe+T8N07qGURNuy
CniCnAciPMMDq4cKrXW/6Ti9qoUgsrx/wDaAO0e2faTNm5LV34KIsiEbmy1SlNZv
287VhbplhUb9eBml/0OzAEJJtYZUl229xA8d+KA3bOo9jzGGPO30CUlbMYUi1ZJb
pCPqn1QrTrrrLIsvyI/zZeCRXqULdjfohcTOYxLynKAc147CKc1NQKzFRKSjtwek
tpWTNwk7VsVx5ER4XpIUMVMgAzMCFFlgVwdS0FTz7Ip2M7GSCEgZCQ3qkSiy5Yq9
fZ5qkt/K5JuzMghogUY2+C5ik0flle8sz8ZZ8oaeoCLG1TYdNo60h0uEaj12UyBP
7pU2kGrOwWfzBBbPVzpmhNRzCi87kXZL7g53wpC2D8l+HzW7rFDI9Npp/cyZLXu9
l9tLq7B5nSSUTIiSbHHh3tIKM5r/XP0m7W5zewlZZ13jZF+k9g4/XxShI0zC4aKI
w2O1DN+B1NaFWno+TIrL2VBbWGebOR/oivzq9ZqdLpn2yAZqgPRfijvLG8nMO6Pa
wuqU/SWSdFDB99v1wpXSqsBW4W8fqEeGD3SrDbugo5Sq30OO0kO3R8rurEsmp+ye
ZomhgJIA/bX9hJ7+FbVM2wXjBcmAjjV9oMq9/BrzFflUO2oTJla6zVmQzlATzGZg
qegzBLbHlDtH1zgbokghUT9IAZ3bp1xhZu5A/kA0L6YlKePy1f7XKx+7fjt/FJDM
NtyvFr44kIqaP9YaxyOrfbQvGVgFkHUnpfqfEEY0JpuhNAsZwYO38dTxrSClpSrx
flawORQdvNMHWuz/+Z7hLvGDYmlrZu6HBg+fe1HV5E2Utgj7GPsUrdoKs4ytOZg1
RpkDjssuiKGuy0+h3e08C3lnTV+0gwGE36R5eWQ2LkRre6yaEY5s90TyBKbKZDOr
UwueNRHcqLiOWbCDC8Po0JzxEE1RB3CAteQp3Tgz3DtRrkYWxkpKDcaswvbD7j2b
+XUJ+6KGhodc47oLTKbsUMWYNR7uFM14+Z9osdnmwiUbIsZnGrno/35uvglzTZZr
Be9+f9CHa9O/yK5YPD2qz8IDgJ/62801tfXOg51BTsMolwls+DLM8oimpy99Z+/d
bJyCvMTB9dPFBMpNaFtebibOIxHNoTQpJ5VFQ4v4aciFmS8iPA6obS4jrE7sYt+/
hb18rM7CDJqIdOYKa9eC7mbFdCZhG5WSMcM/Yefk8JJgsuVsn3a2ahM65an+3xEe
OZjjrJsmEcbYcDLoy7aRpZJFNjGbG6eNVBPuyUtPtNEzIvgKtLiWu5HQgqCRxj2A
lfM7vZrGkniyYU+6EDEUEzaUg1REnPYuzFucqg2n63ev3m4wNCYoxmGxEd85kUCv
HviyElt0LWf+5RwhO0FIradAJdwdWOoz3k9/eb2S2kh+VLqeuKQSgzyD30mbsSVe
qRP9YibpgfS4AdysjScW5RhyhD1Je3tIehZGv7NovRslH/chKUcrhNYvhZJ1rckN
5uXhr7N0v7rrk9ND0gLGZaKw0c7RIBAhrUszkLNwzWoXypki3x37K8z4UueBo5Qz
cbSSx7mGrK2vhzePRMn/ni2N5YZ+Bm84PjU2pDqFpV6H5lxs8sNomkqWU9iJP9xl
60fgePZmtTW+n5CtZ5xo54VR3AOSMAlpe8etP5msTPTK8K5oDNx9Y1GuGbE0lVhs
Pb7nMTvBxmU9vYXntd8axpvE+11j7ZV2TOuH6pJIP+3CVCVFn/VyqWUm4/OBBcri
qAB/YZuup70U0uLcJtTkV4iTcncIzmr81lZyKhf1tSWh8E0kHFu3JrRio2s6SU6y
wnfD/89uupLxXJPv4m8gY6yh2MthXuJzFUzdeqQBEv2Q/QZt4eTXTktsfWzQEacq
ArUMjDv/LdLcAI9xhJxrwxVMVM1//gbLBixQEvxTNLq9Ykqk6nauAvEVw0pcVdVa
tZlf9Mx9ntbtq3vqKMSdYIIFtXP10yQPRYtC6a/ttyuZu2GEvgeMURHPA9y+7e6p
vWPAgdCQo6dI2nyRLLb5UjO7SJFloEqQ+toSTPJLXR+VTDorojC9F6MjbZVB/qj3
je/5/hWIosEIfWC8bnRVKNWrhtYANPpRVGjckPiYc/dGcYoBR39bSuQjYOtr/kuW
Xq66P3JBHydcufsIDdxGH80g0hUrfG2rZGagCzaL/sdKY/L+vjSNuO+m4T6n6aXR
WwUTfnY1EivRUexWme2MrBHQfA+NwoObskOBbJtCFfvcROVUKVptE36MsWJrxEMt
7Bv4h/HAu/P7NeYRa9F9+l4Isy2PYxiuPzfJN/hccr3maR01A5hzhpbRm4SBifVL
rFaV/cLT7EcLFe+RLDhnv5FQaDAIoK7qGmmKGiOgfF4FAovKf5mWSpfMJ9SUWF30
bGQI3GWypQ2FwUknFaoXo8gL/zP5Emxfc+WE/jQ0hk0gbeQjGvjshwYr4l6q1jMt
zYuZN3tMYzSGzOZeJwC4m8bYlD+e6HPj3JZRi39adJiKrOnWeliQ1EeMefobktdn
xwuxJj6EBDqzPhYat47Bj+7ytYX8SWHdH4JLKxqPAJ9KJuYTlLhOsvJLR+GHY/X2
cZ/0jI+VhLKTfud1xl9QtTgFHDV9WR9zAHTj4/XRKazSC/ilZ2i4DG/LJxGbXQNS
Bh6IQEmo/tPTsAmzaAj8nTCdQkonljtRKo2v4c5zknQdTLb6FHHI6hoXLoBLY9HJ
2Rk6Qg+np/NthGvLRR1tZX6Ay1q/OGCTxQ9Z96D7r5BnRtvugqWbpBRV19j3oS2Z
OAK11F9lw8XpviiRuHkFqRhSAPZJpzI2x+Tnwj0XDeEWa+NbIMUTvgEUZeXVtfc6
LKWKYIMDFp244usKiRw+QpoRJ3Ru1zlIan8TFlC64wa5wdi3ulNFHgCEjYuypEYe
8hdDvwMbRfYM80MBqkT5ZYxe1FO8jQ5aI+n0eZF7vx1EyKNIW806SoDehTy2b+J/
epnMaeWd6N6qyZ5pmdbZjUFudG2osp8umzLWUwvtw3P6FWrFkHy8GJtSlpfU+wwZ
WMmFlSbq9yvoTam7Ft3WP2pyLzJjflCltB7CSpSR9tJY20vkEdyfgYO/rCCzw4OM
TdvYGPBKqJ0VObVBWLAIW/zC59iKH9al8ZJAfo8mPICUt8LK6VRGkLlyR1+gKI+h
UiDczXB0hkHTdxjWpDJ8sujNVfVcKOfR+NYbzOyhyQs3hWKLA7dKMJVy/DL1w4Oo
PlUPhb/Wp7X+4Db/szFf44jA/70GEApsJszr4JmR8oWclPBDa0u4aH2dktp/A6Xk
STtMPGiqK9F1hyUucUTcDhdN4FEFGIGdNze7htVu7lwW79Cxt2fVq51VtkpCfD3f
FGlvvXV0XuXGmz6lrIN7w7eEzuela5A3IwyaOGSTN7zVTyHCs2EsMFOciwOs23ME
E0faZEuLUUcEdBDicyce9ne0334FNE+ElcJCPzajLs6Es0kPptdVJPxg/4dBPSzZ
oa0w0MLwNkbq2jEzFlAcOJFyyGyn1h6oRnKQpC7vjMnh4YHaJAlw89Vu76lPZeFk
A5ZgZrICfeZupxy9x67Yw/3qy7EZCR6LYnWRyI5YVBgA9J4hPLWxSIaQCT6Rnwyq
KHH+oPY6RvKjLJdKyXZs3/97L7z205ZH8ZAqhiDjPbF413uChucED0l9G9rqOZxg
Likcqd3nxK2lHWgCS485GmGny7ERL/sBrS34BdLuUVGa61IOukBSVYOePp9YXE9A
7e1x1+ZvcaYSLUqAhI0ZOySnvpOcmrJfhwovJgqozq84ZfdP5cg9FaO5fVB4aWNB
eFGrYcmGVKScih+yDm/cZsP/KHh019kQED7WJiReGbudNGgUkoQzhyaQzIlm38BI
5pvvmIv3ZtGN6lesg1CHMexm+jtDk1W79OedTUyMC4necjoHFcQRiNHjpd/yKUyX
cfVOeA3cq8lbdfZR/AfbD4o56mkQsiFiKMYpXm3rvE2+vO4yXilGVnUTTWQNdZwZ
6JbAm+6khf/DQiD8d6iB/FBcq13eNZ7yF+CFFfgGaQxforUKjIPOwgD+VbFCCcLe
JHP4C5FWrQTgBk22PB2+9+Kp13Kd9R6seZ0sX2oic9ewtqFeIX1jWYN2Og5XtHjY
gegwFz3CedvUryXBh3Xi4miJzCNegqxaXWoHfiCC+1/VW63MbBNiWMee/d13z+p/
D5l8QhZ2a68Yaoe1mzAd76TA17sRk94fvn+Dvvu2PIom1oHVpr8/pFhI0fSpEovP
zI/ubA3ccM+EsIEyBdBDF1ww1Zhx9DEASYCujAXn8JGtiQ06JTggHykwXhIqufhM
tzTXGQ+W152xJDCRil2B0++3GVUXBszESb7HStQRcmRoGy4f05vXpvGDLR7m7gtb
vUDLefRn5jDcc4/ZozoUFrp/sqBl3GrnH7Wyxx72tVVOjgk+YhB6TN3T+ymqM2rY
eLTTvK4lIngxS3ZzgwLCl2h5rNB9hMZkgaD/26CXmcw6LyFBPBYxut8pfqgXvyCK
PQpeMSnyIbZJZvtVd5L6HwZi0yHZ+uWbqSpUOzQi9w3iTIBJUmAP+TgPAP+xop/g
pjpU3DxSPjIEd4tjImdUA6vjoIgxdEzXtUOlGdf/8ncMznXQn4oyjrIzti7RadE/
Ip71HfwnFsdsoeK+amHG7Jz52LGaVU2WPTUoNYCnglcDwx4Wxia5SgBc8AFie2VP
bO4yyRv0XL8/+mWHQuZUIsTk6QSkwqFD5fpLvuXHNWmukXcmB32Ci2TjV5HI6yXA
AWsrUpDcfb/r+tfx6BlOYrxC8d60lKG+V/I2LFv+neYgLeO4LbTHxwqYlkFqtMxN
fESy4UGwrny/H36wB6UtEOu9zh7lDHNeDWjC7eGmV4rSAOjUM285fQN+QMFLJ3a8
2TZKPhoTzrSZc0xmhy1Vnynuwt679De8S/R3Uf9PvCYQpMGqW7HcI+igUmc+xbZH
kymTwRmwhfutJWJSB4F9Ub6ZsKPfFByRVWVFg5QARpiq547qa7Ci50pQimUn2/XT
6jWN6xN2LTv3PKmRMC+sfk+WAZe3XQQxdc9K6NuYRzQ+BCeZq5vfd3fN4xtkgERv
WDkM/4QGvC6F1j/3AlYbe7YHS8Sym7gfJELesZbKljcIWyjFccL6SEA4yD/HdR4z
7wPVV9xomN4+R7efu25/p/hKtdWDrJxF3VxVv9vGtthKTlydIj8FRia+5x1xklCa
xifE8ELv+Xh2ulclqa54jdSEzEtJBu+C5naKlf50GJShWNJKkG79CNvUkueyq8wI
hEpQSvKPj6PAHh5hZS7u4hbF2BBjlXaVdHefHXZYYzKUch54QS6q/NDzZBpDSjrk
vVsfpXXn0g6uUFYWwwz6QqND85EgCuv2FxNO55kUDOEiLOZWgS19v7Glk6imozL9
NoZ7GL5yj+333NnQ9dEg0239EtnQSw4kUwnm//D7EQgvBxTVCUCTC5VKFD/1T1ZW
8ruI8uSiQYpP7uDiMY/AzFMLiz768Q81eOs6vLelbaFmrtPum9dT3aSURgCEOt6n
C/UrBsKwED7oHwTa0ZQ0Q8W+oiUqYw1ruo48xjSWLz2l6uHotiyd/emcFz0Is9ej
LM0RqEZDyA19+0GIfDDMZjhn2vHREuo+DrFRXNfSSDaeM2B+28cIxYzhnYJI1D2c
vOI9sDrgREqTfGLA+RoOQ+YTD/EKH9YseaKL675mufK+rYE3RmTYDQ2AR3pFRDtB
c9Gt4xd/5NxufBiNjSUhXg6jouwocE4O6bENJp8CP1n0nEUNQ3gjWevZ2WQnFoJx
/Kahad0nvfthb1WJoCGMoIun53msE5lq88mAyy4IWHh5uR5p509iMGkbHybwAk4m
+y/JVoP4txPpxSzKBI6JEVe7zleL/qSsWfka/fwEYvGEREBXyF3303anHacWF+OZ
RSR/+dF+klnEoWZFrOQYlyXvKOcJd2wnf5LqA1gWj/rlZQ98vyOg6p4RnRVyYkA7
czCooxJV7uHPk9cpAUEst83qN31AvwoQglJeuRbe1CGQYnbWFmMYUpmWfeeYj2Vw
u8uvyiJ2N9DVAowaJGDsL+qYF+1HtQJpzeg+06byOIHgp++LJ/gdx+9kHVy+79VD
uOK/JwKLW2CFAievPAKpNRQcVMTKxNwuUja8otNiJUUrKO1L5sfK429X2mmHemzX
JT+vAj8tlD74fqQjZHlc5fPyT7IEv0oa4vAUXcTqBhLlzW+YU9zq5xsTa6OoLyNe
qsoJnGKuae7icbyFqA+eN0ltVazyxW9lQxf68FpQ5ZTAHgOf9Arw9TrlWtTfQH8V
fIeSdXqlQ6bkFyaiuS/GfvxI2kwxTXXwmJtbQdroT3s41RbwExZ6dXp+Rcq7aVzZ
IKjWgRLZlwqF7fs6eIr1EYvt/vL3h5kr9dOEwva5aTxyBe2XqOlF/lGEgziEG9la
mouikZhneDp15AhJjJucQ9k+PQy/6ur2rwa7bq5Fi6UuMT435KSDGrpqow7jBKrB
+sh57aY0zUvFD9K0m9MgSnSmP6jv34ydtszgbiOe95lB3/XolfezyS3z8take16n
xBuJsbGIktikggWAemckdTcPYFWAfDAzlcTO+72mRucOjJVw6HAsyvCDOLDf7Z+F
ssKCmGQWu3L9xlujYoV72IYNlXRX8T9xFcgVCIBZyd2CKoGuJ8Nl/nGT81JwGTlL
uGH5fVgI3orN0PMvCnZR7ewp41f26U00rI3zwRKrv/IiwS1yYHmj/XBUT1efuxDh
lg7RGNiiaSOQUYr+He0XQCni/AAPd6gYM4O6WaMgW2tYdJ8Y6mLBr6xteyB5kBmR
Gkk3OU6Y4fD02pOOlbLduR5e99lg1kzEDmHtsdEdEBSZcCA/354OSI7lFhY+SCD9
JtGwGd6SrUXMirzqBfTTIgJHuNL+7ocjYk7A7A1AExyp4xCLNsCQMQGOXFdLGlrG
0gj2rHTmTIhvbynu4Z1inb8oXcLEh3idgoIXW1lf1uUpvhv+z/EEpg3Id24ukmtO
Ul8iL+y1CtrfPtgXA5KMhSfbddxCwRsL3mhC6laO4AkEyEDGH4haT50s6robUWFf
eHhE6z4u8GO8u6CwPHDmrJHqvDkv1Q4OD22obslWHSSRCfVo3bg4lgvSBS/ux+t5
r5d6pPMjZD8DJ0Xp7mWfidaiD+GhjHfH05QaYBIBRdYcjKSFVUQ/LqPpQn1emHly
kLtqzltfasiLfMPjCSgR9GRgqn90oo5fYakxsghGnoAMwjZyrvs0K/kbD180gaYf
MQOpTMUMixGJ7K61CVGLIoIrF0S6PPZdL/3wzeEp5fEj7B4u6nfpA3/bOYPJbhAR
spkMui6G+l2VhjCICpsadbyv5u5CeR8HPNEGQrr+ZfAXwjVgXmIbyvaSIuq8hXyw
4I2lNIdW8npxOg9RPmxr0jZhVGSup3ewUv9Pl/RQIiOzZ97pfjWpAY+AgnS6f9lp
gVUQcgZm9d1M1sFHGMaNEj/Q15En+vPrs/ErNf4LKXgNuaamS3rSv6y3sShyMkgu
dubsTd9AJCHwUujcCSQS5mNcqfGkF1wvFORQkPKL8JiE26G8maUE1UnKJKR6XcL9
6tZP3AAEzqyeQaKOJn7Lo+s+BL+PXwbWFbgOsb4gNWIbE2QPihWeYO+0SvRmN4e8
CYPAtQEpZbBZZRC172M1UfeFKZoqzh2LonXCxlKiblxcaVdDpIWlNQMUSFWxIM7K
nKC0qrT+VVaoVb3dxY3e4PINx51TwWVX8Mml1y8IzYDdWNsGJe0o8zlEaZzUWYgA
zfEfNcVcxnTlNlE8o0aXYeLP2rmO+w3puhx5CSqTTICcih/ZK11lLGI37EoU49OA
irUEwX50siiUa6UlToIM53OcvSNH3jZaVuObadnp8qjeecbta9+jgCC5s67qaLZP
BAEcVYmprOnSOmArrkU44slWkf0ukq6mTy1bPAlTe/fglUU4Lvt1PiuKrZe5+rE+
ZU1zDfq5A6hbPED8EQPw6Z5Xy34OEeqsIAXxZNCGeFjMnebeaHf0SbM1sROz6aGD
pGyGj6cXTwD/aSH2laRkyMAcTNVEgIivmSp36eWVvsjAmfSTdClJnuro8rkiW47u
rGAFR2+f7Wx2ydX6FSfvDK2lxx4oFYwT/4mvm/ktV+hicGvDSV9lKQYDQmM2zHMZ
kzHQDa/3kABdzHJ9LNQtytGvV/pJ6dOcRobBNVUNtfYi8oDjCiesIJlwJ3CzrxNW
gGs1g9yRg5m+UkY/EejQtPDknGc6HIiFJDilB/eZjtt8LV0SAv9LYRcG9QdI23JN
g2BiGUX8yMpevHeFRc41nW3W8Gc6+tv9bKpNLusdRCEcPjH4EmqFsEwdePvBRdOn
+CppvWh/rPKj8swL0rMND2zs9K+7Y8t96NIlRuh0TICuIPWQJ/nAod8oSMcT6H1m
Re73JSKelsIDFbQKcEcPIA658FvNj/AOatyMUyYKmWornHgYocLIb8KOTVy8WjZv
ZCtOvozqDGYgHNeDjR1tlsWrPLCwSDtqp7Djd6NKgI7a5Oj2VopxkLtJ48uzTNBL
BWe1uIZvH52SwqZKXT78foXxsFPz6x6YAwPmTC6MwFOhDiFoI1WC5jIqC+nuBccY
mFJf3WGCsHBCjclDw1VRBPdnx7vWYzxUvFN+Ps/CqSdbZzivNowpeX0tVK+6rghx
ZWeGEUNNDi6vphMLvdgc00KV45F5LHAJLnMQ4lNLQ33Zzy6/hefV2Fgt+j15Ri+f
IbtSTs1PtXUnWw2YgofX2T12pEYzFIV/Go3w8fyV+ozQ37hhS7gTY6BysZbnO/X6
odYuofuhjKX82CmnZSKejzO5nuqpIBsA2lFEOwA4p4UG1pw6qOidxo/CY1Ytr38y
RuotTMldlXpDpSac4RDPhRu/0Fz9qY4ueIP5oellO4EUPuVXRLTcP7BDWSFebY23
DGd3zHksgqd6tEyG2+P0bwaDOwLziiOMbDHd0mITVg61z4arLTngThAy5WxzIfUV
cy2fy7+J84on286I0RFaUNgkYMU5PwiaS1hBrWZF6FpGirnWw2Own1+JAhwfnGzG
HQTtCtsfgijY5cwHM6TPRx3S5B5z/3tlgkN/sDvprnvjTiO6cQw+GaOsunUywqTE
nCvDrSgx+SRjtrxet38N4oTa0ZOAGXdNnqXus9P+OlWTSFHpBrC31FMu9q5b0c7N
+aa3Rz/sFPP14Y0vTS9tTfjwKI4s1bhirjej87mHUbmIDy22/QqnYBvYd/cpGp9u
BN1yfRatHJIMc7ake7SXeyqPCCVIC/+BKHFd/IxpoHbrnEs7K5pTGJsGJBFADRYe
ZfpOTP9gRQz6lMS3rzP01ZgPX/W4drOKG976wMuHKAkO9kFXVB5gwfjNFKJNTlic
+vHDAcmpVoM7GhefU5khjJV+jk7IgRlOXW7FMOZvonCTDV+FBcriKTb34l8WiQHt
6iVfYxyLH4piB5BxibfJtHdcKUEiaY5tEg5ynxd6K/UoW2ZQS5+S0k42Oz+I8gPm
oZEyogcuCcUH6ynGauPN2IHslNLjJ44ynpGy0zm1Gq3c+NdzItELPjhq9R4dIWAH
LVBj/7P5r5B9Z/rVy8SEG96h9uPMkcKfFk1Y0cYc4k4SLsH2oA5238feInF+arlo
JnKz9TLO//u9AyhyfHzlS6MxSpPx27W0J5fG5nO+a0/JGtP5OCBSEdhV38Kn15/p
JGdkIAclwIuURNXh2FnUDRjibjSgGTc2J1EHLJvHfYvEkt8azqiOCw8rxX8ylRbN
E5k0OERKdvcOCH15yeKLCOLON8/i+KeIT9w9fVYQqOlLSWfJJJqpc19/ewhv/wyv
cbpjIaNxuyDAfQHFGm1NYb8ZJtQjDEwyVpLOy22gVU67KkfJ5g+NPQD9iYRDdbw8
wlKMaZuUnVJjF+BHAB/L3UnVW6bOnS/9GkVry6RwVelO9yH0z8EUS9Ac3n8hwmdv
4xkuID9iOAPyoKKeGVtxnVxJzNEnldekU1DPAOPCOmkSbkt/gu2qdBq4asMOpvMo
TNmeuc3HhJ3xJNYwJn5+OEkFMjVqp1RF/5a5IjmuMmdSkdDM4q62G9JTE6EXJmLt
5sCkoG+5blSI4j3BlIsyl01jq2h7JMgAYSb3TFVpzoasKY4docRHF3MUO8UNAnXR
gm3q4KqAkVsJLwwSKzBDnauamYAnGmMJL3gvB355l5bNgHCpKgJOHjsH+oA9Kuxy
ie0KxM0aEmmOogPT7hoR+YmwLQrM+adxH0kD5757YEzHWO9GDdH+e4p36MRLKi1o
7G6oAvcowbg5V0ecRfZHexDiaIcwvL+GyUWzRswhkqI3obW1Vk/oQwSph4+jVJoC
Q6KcyqqE8R/cUGWwopEQqkiItwaVJcKEgDX4rkGGaf6iVXTRrAjzGj3j58nGtw0w
1wlWgpneTDbyAczA06Bl0yHyZPsd9P7YRaJFOBem5VVWmOyo+qeIiET9JTI5PbeJ
b5J3C0a+P0xAvOpNr25eSEenZNiA2ztt0K9JwiKWseU10r4RtcUxnoH/bUdqbTan
norL9gcLnOStO7gvnxOtcnXJ0h8byvHJDui9kyDdWDbNf1REXnld90zWTMnxrUSz
eWgK3Wt7s8iCEQKrGVqpSXmfSWFIPWd5mMdevUOChj73zWRuelLdZhBbYr0l4Tmx
8h3Hv4j4lfmqFqDK+L2k1Gt9xWTPgnuxnKMTSm50V+SzPuwtG9Rk7xVPM6/aVuRe
w1VqobG1bmlNFavZtcKxQvkyuAVXBTS16PQaICW0SuloFlNAXMNcpS7/gpIapmdD
XFidUX/2DuQ4MB3IuJygFBcWPyfKf50ienx4GrO3LdQRvbW8nxnwoRVWSjonNwaU
z4NtsRDRmW35t+onQ+UsJBtMgH0Hk+XrYBtym55885+2pjUXFnQqX2ZiuK5l6uRb
Ki4tyuUIxpYosvQbTfp7IrObTGiC87uOjJFNtQC0z7imGnJY1MB7gsvOgkpdTpOE
n0ZfmpMhXV5zkYEdRQOf570Xg3u+nz5lsZxLFtdSEwlXtsJAleZbtsUCLWAjisLl
HEAfZKXj3j4zdaH8XaqWYIvrBgTHzldyUCdP8cPiqkIMUiZv0RNOc729E7+CEDJj
B0KUOXteb4NtSmygth7Qmv6GcaX1TKUXAssElQJhCHoZg44GIgqVWFRYxNITeN2n
Pmh8y3yyGeLCVEoWIe06KifWpdHfcUIBSeRBSTX2zEyAMjQlteo2jsLEqJGhsbGv
+1qYZTsseRAYgGq7bM69sRck22ZmPFYpnsoX2GWxMZYXtrGHCmGTbN51/ze4sV9D
iNYMC62MWW4sb/DJkLonkUInIW2Vxxc/4Z1MiO2USKoyQKDC+ZC43iPKoF1QnO3R
k7MW2Ug4csH0UtVeOPW20DsLP20THAnfYeFU+A2cZOdgfC4zGHpz8/qWZ5j235+z
oUiY+Tu12E84m8t2waVbihh0rfehwWwlJQnizJZDCx6PvhjAmHfwwIDEGYVv5wYf
s/uJb5yK5jtpxAlB1IdGxqmvrQbtWp61o2LizwR928z4w3zSui43w6cA6d10/wVk
VHrOSiLum3cfG0/H75CikUqLYdRtSMSvpVEd1u6zXd7LTDkBacFT7/b1d0jcVPNR
GMxWl9BsS0cWZ18K62pmxXTVlTVcG+AP1K2UxG5STGebS/d/ku4T5fUwNOoRexUf
uPAimdpwMb+u0c/Z90YrA/GuYf5Yy2fjNvWTccrAKJgWywNOn+rSIBZSA3sA3oeE
jBe+vFJ1BNXy5jMjoPvF4wHOaJZuQKc5NisoCSwoV3MmsGiAWHtSbDur+ouc0BMo
yX26DJSOfdHX2302QXdpUd+xPSFb6UK2g3EZmO/5Z/11Zq4wB1AZ/i5UFVt9flRq
eWdANj2mdKUQm7FeK2Rn7l0A/c7V9183cGgRQxFLgmc73K96NaSrMJtZgBY0LLOD
+L8lEYar+XnUWTqpy60NCDvLkSktB15PWL/SNTzbncsv/oPj/afE/DtkyMNsy0aV
cxo4Mmi1bDLN6xazRKC3YurHm7Tv5k/9laEvWKiPaYEOeiI5BppPLhbxf3rsUha4
BeiCin4LHskBAlpIeEYWXGuGU1/qeRl9coYf5KSk97N8PX0/esF65V+MpEjJGdOz
AAf9UCevAFMH9ToD1CFeoI+dJCz+3RxaSuRukHk1UWmdkv6VLCchk3z4OXH6sPM4
Q8DQzlqoYZ007lHnc3ABcSmBL1Zj8C5/uYqCmSCxm9zbx97EnGQEndDJHq03xvmh
Pr0COENXIxYDP/z6bf2KVMC3zrfr03SLH13mH9ohAN4e649yofnBc07b8YXdT73w
Tc5piNSwbP6SGKyZWpKu3sRhYBDqvRFM8LN2G+/NSsRy21BELpwivpHgvkkYudlf
K+y/MgJEekE1m8Ekv4uZefTtvB2nzmSCfzoCzED2HHBAGMmNGRAxzC8sK1HrorEj
GXYwAL8i7BAII5ITJ8bUjeqm+q3meNCnNi9tuvJf4tSSR+xxxjs9umKJNLfY2w2Z
i4cKWYVub23Qeq+JQNafwOAxM7bBh+kWSauizVJJFUjQDW4U71K9YZArhmcacvR+
Jbzhq0azp18+nFGnXIV1OdeK1RNBnxl4EMwPcOTA5jx/luasI/NODfHiatGbGbuh
Craqin7EHFznOEXlOkbwL7vlDsYjlvH/ehWaOHK6zAkI8A+wzEz3Xdx+xkNJpqSR
iZjqUMddxWyN8j7QCq1URDMwtAYa2S6Ed3AdaFblhLCN6w50jWQBVwhMGuEdqi9T
pxexLpY32G8QXOfHjoS47gUMUv1ZXFPlXTuD5exuvY2MBWQwMuAO8zjbzYWbgGvM
bXAI+4uesC1XjWKYTU0qfnkexPuBqrctL4HXot2pPocWiPbEwocgrxZ6/xmMzWKi
Px2s7PUoqlM1mdhxFJ1BzoN3bFm+2Ar7wfd2HtXUYpwcofdzrXtxG/RKCYKsyfrE
5QMQvrTgsjwo3kSEW1YiIQkcVm+6qLXitOY6AF9ZIKrwiMCXr6cV8XC3gGqnxqb1
bmv2Q9RaONv2c2Pbr+W8wDHAy+iQgqumpwQ/rgrQ6dibU21XmaUhEcZUNLtSXySh
guHIYQfL6bpopgPAvrAm0soLwT3R++XWU/Tn6fkpLS0xeUhxd1XfpCFT7EXRcD9l
FYy3DLG6kEpElSeiAiE+f7CtBhZiTNrX4+W7wu7AKLljAc0HrLzYe9XWbqzgBMR/
O9ITWXQjjHvh4DoE0sInUoTTgCQVubR4cr1ntnZ0MzzA7CNSBs7RHBI4eZTNSRKl
fd+N/nSjk/J8GNM8W7HLoH0GsD66sQXbGJx/SsveTAE3bji/JcYmmnY4CzRz2J2x
RUQgO2nNs4wy5vTgHLv8Njqi1teWwHjjsyVakVvkGh8w4nfoeTcFnr90cx174NX2
PN4oYle20cNF3h7ffCR3fEaT1IXRaoz/uPPtQKacUh5EKgQVyoybpvufnjP7G3E9
Ds3g+/e00CMAQ3ecndwIuhrOU4kXI61NY/hJVcntsFiW7SKYwz5EAegcRJ1b1cHb
YiTPJrux7TUYrPu2Fhf4FUHs+qD5LoWpFNq1WiSifYK567M1+QlTbbDuoievDciy
YtANFI6O8OddPeNI3jzw1NITNIeiAUDE+EVgv7J+hq8lwbj0F4OMJsY5IHAcX9zZ
wiT/vUP2k+KR+oLj+kojShUSGmrSU3tUs0VqvumgTEYG+RIu94hGvHFUXn0J97nm
H06154JxNyZSe13+14OOMrUYOBR/Tz/gzhP+ToHyZ5pkSmG4pfJpQ4JemK2owtTc
s1465omCCD3vfcOiEwymY/FYAKVwlky1az4q2gq11FojPVF9cptA36GlkoPu8lfh
K7KdC7gpusCG0q2AFZL45uIR5Z1alMmAdtK8Zwc/W6SadfA4FqfQXkLU4iEM3gJ4
/9xo3yyrp+SiUaX93Zg7SgOI021O5OIrYe4/SiCRQJjqKXTzLSFju0624y1DL1Vy
AmHp0hhY5Q4Aq38S3W55dyn/ql8vhXlLpj4sQwA5An/xKZt/EGyl0dX4XdMR/eYb
B1FizduB8xgt1VOchRLhe5VjeIZqmavHw8Prx7KvwHEXdax0ODk7MJ9jTLa1KaRC
yhebwCG6RxPiyTQIvhpjsD5MqY3CSEaXXrwgC/eTEfolnKAj05ExJ3VqKvhoZq5w
DRTbmkB7wui8kU0EzLDK57QHmL0VFUK0sMPf3iRewgqj07eiMJzO0A2ON8Pg5ZMI
6+Frj2EAmBk5k+aSeVHFmbrLIiut9Spch2bc7ykKTwbeTEBafO/jVbfjEJew3Vwv
L4FWtRA3lcGMyo60sfbZNfhGHo4fngPn34Ok8Pfnaf8SpSXT8vIAMmQt9l8npFYu
4jRjFj9lidFUkLZoVHPjvOSf5FlkY2BaJ69+MLjXEKicbi4Z7Vw7BkoGgIAbMOwL
1W+tL2aq5egf89Kt/oz3oZb2iOR8Z8xv2siJ9cCu4BKXgPuajHlaQbDn3W0f0zjp
NavkRK8fG6hF7PK2W+4HRUuuryj5pcbE+9tx1XfTZr/Woc+xa4wcyzlcJwbJNTGl
52BIB+H+YZL0/PrJzFdX+zPUD0nVujJ7JfNKY4mUYLfQACJ//YUh4VBp67RyYsPW
fGbXXt23HFZ3okqZIV1Quo7771Qbz14+z3CExosm4FLNiFltMpZrNe/9f6fvfIZX
eyRE9LewSlje/M/P41BzwR2EPHI8iL95moDrrX/CXmJuQvt/4ZEWf0g9a+cgbCt1
IAexEdbSrEHK4GLcFTjxQIqxfG6/Eki3BKngMKWtmBMxupokGo2KptTlOp5PYz0f
iuoye5VhBmJuojFGuvgtlHtXMkyWeFKa4SN8RNSbZReRCSeG5vsmUvYH1vZa5cSm
gH3DopeGcO8fQhhjjVJd1JD3rbjNKNuZi03WHxmbw7t/cQPt4/Y1z5qgR44jQPWQ
4mhluyGM60RdlXVL0TH1cPwuSMqz9WR8r1jm8mAEzmmqru8CrpLAV3rvQDBR4kJ9
sY7H5pT8Y3HD0PD3mzzn5QG97uf6wbI19+HC3WcYPN/1fmreL0w5YM51P/fKUInb
XtYENcvWWLv/I3Ztsbbk7WLrFFM2BSOv2NEeQ54c5i9xP5BmhxOiJFRcXLrFdeHy
mg/E/X6od8oosJk1s/94xvyNLlSi2LGHCDtSfgg0wBt7//k1DnDbJNjFYMvGqniN
2Z4DvCCfsZwr+JOkENnC60HIcmHO663Fec6hqW4lRvpCOKmhmSxlwpZOK6YoRWRi
T8wscHUvN40cQ6l9UVdFrlw0XDKLQi9q27knMY6MHppnmFtsOQMkpJrmWcpCAwFY
cweRPzQSVb/JBWeKTu0vS1+/Hr4PcVrAYM9JzMk1M8fvvBG8ApRiqck9kmTeOn0x
x4T105W/1IY2bfiU+ygshS4BhIhq1mgU2ecBZyrfsg3G4fosbonrelJsFDXwGbJH
T6+xVYUDOgblCGG1nTaRNIgi2EG0UTc91Pv5R2mFcIgBe0AMhNwhI27XrQent8dX
UN54oTV6csBtduulUkRSpm5c5NGjNXaHF6tevdYjaT4OGNFxMymKdgAiuapY33+G
5vf+IImyg8eF0KxdzJTHdYCvORatFW60frBche4WQFVoVuYfWnPhSiW4Nw3IuQU9
fzspZns9t5psythny8CPdp5tyEyroblcBJwBeFL0KMnROxcACLQ7IZQlaPeKvji9
Xzg4Q7ng68uLGYAJ2k9d7KELFFRb2pOoZApDu+BmfzKo94UpvBlq+g6TEqC6IGvK
ad96v4Q+WR+AhjEod+pQZYIgIyH+L30JDTaT8HWdItmKouzHzvyAWYIbp/jmCdEZ
CjtP9YPOju3XheL7fDMDhKLyrgjz4e93fvhzNyYHG040AbJZjRSzvxvW0OmEy4U1
EmpfA5GHs4YJVxPZ9BJY5/dHQPj+vxHSqT1prt307sKAcb0/dHwpu2W38rLZ9yR1
U8U/6hAfSFri5xsZRPeSORTwoFSLUWwQarGQSDu4CBDsljrMYV5dXc1ptD2rPYi3
rHEYXoz5mUSDqf34n67HWcbubQIirSz8KiMSVHw1VyIP1P8ptBc6PlTFz7Z5DUle
AzxbRzOAzuBADPCHQ0Ozibj+vqj4Zt9+wXwMul5ujAvPLsKRXIQVk2DjVcfy6eWX
N5i1QZt9aOpDo9PCISQL9Klegyo9JohoePVSylLQ+slkbJ9Bzdl6Bhr8S+lcL2mY
02fbZWyKSjYHsoNKg9BYUeF1K28Al4vILTG95dGXWVr1GTHeNl9s7P5T839tu+Xs
cISoH1dShR2Yf1pf0QEcwdB04uoMFqkq0HFKizLAmyadumtcG1sLp2F91kXu0ga1
ECUqqmZ3qzX8mR5geDAvFWIz6dLBqck0oyw4ixv5+MHZF3Ogp5bmkjH7CPBbVKQa
yzITnVUHq9q73bdzvY9IIRfdsOGcPLgvs3Qemt5f1qUNMz8YP5d/EfOts5gdal4R
Cjbh6ogzdahIRBzG8lFP+U7aKnIkrNZVA+PEdENXPX8op7i71zDRzvSLGU/GLIor
+F6rU1W9VRVPmw71zR6YhWPwg2KematVWDJGWsmqr8RKQ7LShX4dLZLOEzNaM8ia
qxy+MS+ba/AlT4KSoyvABSHASx2le3NJtjzs+qIDH6HN4jND75kxr2lYNme05NpJ
G3LgbAA4bxnbemouo/oLubNh1cZ0qAlCDlMyZVHJPfftidQE0B80e1DPSiC/eSqD
DVuSWAkwHBKtTMMLQbDsZx8VRNpWkvfxmYjOVkyepUR+IAALw1R0t/3oV77K2zst
2HR17d1Q/0YtUcx/I/vmoRt6ZQfT2hcBrZAjPSnxKTcLXGoU/y1SorCzEtFiAlhQ
yNtsCiO5BQ0lF/Y9Fcf6j4j5zcGf8epa4SmbENK9YqhH43gghRMcxFRHQrzqcqF8
5wPiS/RpMep6/5LS0uuRFamek9m2XJb0lu53dY7bQRJ8jvHF3sOLorTOT4qfHwD+
r6QDR23ZqUhhysvSx8a6pqLkdi9Dv5cM2ekV7FDLbtP48W6Oye7sYlE5fPfM287L
K/cU/JDTKki+cL3aVtdp9vmLKcRPfuB/xJQipYAU3nDE+atPuxdNJgjrbrtoqotq
u5+jX52hP+rQVGj9eQArsk33zzaemmxgf1MgUHhNnd30ALQUI4YKiSrcOIKBCSlS
vpIo16YFEoLbeFLvZ0wXkadhznSm7r0i5/BPW6tBSNTTtkAHqGxXFfzA5G0cSnw1
oepCxcEVsT+1Vk6YApiZ9x/An76aCkJr2UoMjolBq5oICKy2aQIh6NNn+iPVMEad
rCIuIJ2oovknPx3tqPuKlnCSRk60J5XkFBG1SBNbZhSF1F69pxjD4qZJG/BER1qC
HqzVOLJ23K+829uhiJzwIhQkor0CXebwRc3AU6Qi94lqpkGk9w62BWyRS7hPS08D
SSqxH7HGHSgAA1ZNvUb8YuNRhuWodn8k1hv7zcYkPsAoTYEzQdTnLX580nyAwTnh
cE/MY7mpXP2Muau3/NWSzvScYGa7E4Xpj1YKsW2XBHJ2rThgXeLJl8cCXbb9kHZ0
ztoa2nTj3kQcMtpDaKlkrXo6RoSlEwxQXRVDEpP+yYCkjf4Ya93jJvibF1QHKrUA
2++mmssu01hOnQLxOPPdYQBNGWDiZTxQnwF0/uapR2+kT6urMAEeQsngHANk1eog
ek/7CIZ4YPiQqAfLEIyBfrO6Y5DcSnNaoZnkwL7fCzfJy0ieqel/g4V0vuernyQb
fsIM8sJOYWDOo4pnLOxVmc1vmoa11wociPnKyE7W9NKSfWeXfZ7flIcq4zgqB2cB
fngObgoMpYUX93omv5oTIl4oyP42bSqkmuAm/zs+xiLAqEjGig59Ty5POoW3jYOg
hJFgdJv+P0H3fKVb0gFSuh/HLXO4Ek4wAWCyq0MTrTn1xunACahUiJUxj1NihY5c
d+IsI5L9VBJrtdtwEvguaLyl0OoH89z8l6g1Vn17qb9mBTm6C7Npw9FSgCM3R1Xk
8fn5rXp92+SViTchM9oSUVMFqDYWLvXbWLY8Y/3+oHZyF6yluESJY7Ymp9Q+2sCF
2qDzBMlzujDA2J+V6bSLwHYT3SON5RtbL1j6gFSeimrf96/oPPmHuEkbiKYnTzXK
9OuZBsZQhxzb8nNaQd1xNsrNXEpUTqajAcGZ8X6n4OTomvbZPub/eXt54GOCoHjv
K6UCGSBM+rZDYlChw8lOP8W/6aRXPYVb5Bazyg8PhubalNYr3AfJp0o5on0uHELr
nP+9X8TDL7ytildzJ9g5NC3zjcvmeGSYrtRdctANVFcHHqDpbQ2sfhY0GHp5kQCo
21AsuIZBJY6MS5w6OsdaCU19Ex1IqGBH1ONgnd2Q4o4INtIcqFI7XVnyeC5x9uDz
dbO/2w81X4nCLmPKARwt3frTeLGMAbVFtYIGRDZbgclhWBKeJNvtRyVGZgeKKl1L
GpD9+Ztx2H4+UE5P7/ipWoNw2qdFgIPXuys/0PXJEhUAg+INfwRug+MRrC+Ch8zs
Jjan9VAkM9COLpk8DN2r1BajkLEa1y4MD1JvzU994vHjgZCOsfktYz7ax4uLFdyq
NxwbXq+7RAWnbsHLw7Owzjbn0yW5++C/YXtEtbE52OhRvgd4SUgJmbh5j2CYXFdh
9fZQQbCwf68HQRvdFsfR/S18Ff2LgZOwuzpt4+GyRjchyL4tUJqARDZvCPzuV6AK
OjqR8jlx1DfeoZETzldxExzcKbk7Itm9H1ulWIyWoWK9Jx9TNKY2GSQ5NqCnaySd
T3yEQrcNrzF/14sUlvTu0WXOOC8sOIuxQSthq5neJXAnVGHNdfy+oXjZ1oHlNAEF
YDTSZEdTg20h3dhTXMxTAi+WK5o9r1a3D3PgmRUriVr4eauRbmy2xL9rq7fMLDkv
XAWPBvi12zitI0Uyhwio9wb/xNSEldQtoxb7HTo+pEvEdB4xoHWMKHsPQIBIdv5R
Q2k5haxkObvEKSDDUFpJsQ5IH0yx1SaiusCK3uopyBHM8APsCxfX8qlHso1rw3z0
hXdRZlZwIBleNMuW7NNthu2qJ5t2me1lrDaImhGE16H5aZb6J9Nqcz13Kr0c/Pew
MbHTK94XOQ0GESU1fadq2UIp2VHr+Jdtaji7tUhB8hQE2jxeGzjfSnLzVBXHle1d
L19eeDk6CZxc2WfHDZAr4WA4W6jju3RyOgtk70f0Cr47JnODu9rgQiOrDWpBPNL6
Q2R+EoWDiglhQfP9BaHZL3WlSFgXfxGm2pVgbXU94Y8LLURlIeX+S0RjyQph/f9G
cN3fTBU6zLQwNKsWHS2Nj8eui81BadB9lXLl7FL6E1CTSl2OB6GBmri+oc+WZrTt
P3c0vk7JH6j1AkfVz7NtoJA1vNP9Tw97xAyy/6Uq2bq3VcR3wIdXF5Py5ubvRSH7
XHExCUxGiXHzmVb5v97N2UiHNmkgFxeNKch7+mc9y0amVZY5U/Ol9tLmx1AxXcwF
k61mxbmhr0//uMJYg2+DHjrqSC+CHbRVcQGLoSpeCYoo7T4qH5SPdYb3gzrpcE8n
i3WJs7byX9QtrtJObSRNdPWjoSeTCe4xrxkq/bYagjmQHWrv0k2CLfCMJxLEbwGA
W+Ms5Dr+MYp4E5eKZ3oF6Aw5Cnms/vShEPe79aXX3sH9ycB5j+NOBhUrHzo5Srxb
1smj64ILBQsXjM4ICYqiMqqWHPFh+qUx0N1e2aizq62pGmM7wlAEbO9U76x7h+Eq
ybpnn7v0xM1e428attho52/P+bvb9Jo2Ai2xiyfJWSMRsNsvGejVZBpbQsnmZSBd
VxdmiVSfuCXZpASqdhpqEITLGs3mVnqCxyeb/7x1JANqslr0KostXl3BAnL9C83t
BsG/7c1rmMGf/d0twLNxfBhjwZxsiPU8nu0Ja9SqUn/U0r2BwSaurNt1oL6MGrH/
1zJabLNbeX1LxJABZBUjjUkOwO2sq587vSVWHR3XF1S2u18/tdnPWIIVIuG50phs
0p02OIM8P+iwddeEC+FmPeN+Sa1Yd6nLuZFuykMsh8BSX5NzapKtkIxRCC4t3z8i
XYNEroiAMg3piBOfTz3a/hV/fR6UHpDdfF1yJXBMFbWpHAriMHikU/p9RKA1/6CD
FXw9OZ3JgU1h+taPyH0Vo/7xJUto8tkpuIz+wwTVOt4i6qpIf8/2XNcF9HgWfFsz
bDYGASJtbJ4rT2MBWLTxkBhZIKzJPEjixnbiOdQi3DsI9O6Wu4M8LnaVmVxQntbi
fqZ6LGZ+i6BKxDM8N6/OwCAFMCB9oo3owujlJYUI70ya2QXPk5lrjh66tfAQ4RO7
r9N/C8BZf8Pw39kucKlECnRY2B5ZzfjTdFijYBdZNlqZWNtVr6chbz5FmIfvg/c2
h/+uqdH1XSoBKybcmcPxZACXvysgTYQDxQ2T2cJjXpDg3e3khBOZrvzKReGRKI3O
lMbAoIITMD+0fgm3qLXdWZ5ffGgaj9psit32A+f/8pZOBxkoG5h3/348hAC8K9Nt
ieydCTJoRMb5GENV5gb7L0HGpjUurvGVD3m86duk3u0DBVvu4b35PxhGHLnAHq1U
B9pc1J5T3m5vsQgI8+0wvo6YmoXWUlmpolHFLOw12nWcIqnVgjXvf/vAqurHSso1
o9ZAJ9/j1WZS/nXDjDrDhBQmd5dVqVXAHwgSYjIbSq4/T5TQJ/86ZoH31JEy4wE3
Uz3Np/VTahlcsCHsg9eC6EZU+b5ZrrtZom5LphOr/CudCJFlu3cXYbSgl0tXXgIW
tRcvgt0ztYpGtWtrK35o7iCiArQZOMNimiXtQwAgCqrNgkqR5KkQCwfrceK2kP0q
o8rqZx/+7e+rbc1Koi2TYOf/GFe1M9SdYHanFfPkSYs72K9kc1zONKLpSVgUs1st
WuI9PaPr+FdS0zVEcKLd522W36ot5EEF+oa1TsO7yxA5UEZz5fHQsb3ceRiz8RUU
0u89oPRM5nJ0eAqlB19lEIyOgNgNoO1jujdRGDwEaLdWMCrhnswPyyTb/4K9x5yj
eMZiYb4A20kAomVNDsOtpVL4Jycy1mgQUqXlCwMDG6elAUBKs+tQvrBehUNSP/XK
qZVur3wh/miyYhdWHku/1QcK5ov/iUTE0+LzDz4PhDcthJAufBfmkv4CNuKHseWS
GCA1x/LKhFohAHTamjGFvFXsbrdiSe8lErxfsit8SWDdCxUJ4OIZcgMlFYswvYb5
NnBZMSZY23pi8DignbrSS6AKsFVXJ7hmKdMZSApxs4VQOulbfS0VeQs+2dLShncU
HqB6cpAPusUK+fc3DWw23ZODcee2+xBFizGWQTh1nN58qHbIdm00lAJO66ZvTf26
SRCV063tkdwchCtkWGd+PQbPnPsuSaOhLQc6Wh/WHKtV4Kqa3zqE29QWCrUdhNbc
pSsoO47CQW/cAVh+EMgXRGTapUIyKLaNLcuwxkOMy6TX4UwsVlVSobTlM3IbHFys
bPc3Ewz2vdDOuNa9AsGWO5thCUwPPvq0tOT5SbHk1l43qBRUoDbi1cmO3sH1Y/wz
XwYMY/1EmRPLj88ijQTWMa7xZLCbrartEEq5fJLYgvtU+9MvWRxqoXuSHgzy5W3E
dSbS4US9jTGlNu/zR86yWCZsom7OliyWiF02sriA1GpdzCh4ft9K4a1CYDg9PaIn
44B8Wrol0KSFGmHbk/Cg4G8AC3OToHR9h0rRK5QnHsyYwJ25Ux8/RW1L6UEUWsrB
0oXSetn0Ix5FjMx6acBfp2UA3LYiMJwnXZ/H9Oov6mG8OpfSwikAhMH6c2Hjt3sg
sWxej8BUgU8e5zAV7CyK9aRA/5P0+yWmSxaKONd1VuErp7VqW+f4B6P0DJEtp1Rw
YWVaWM2CUtC0RLBLfAyQbVIQp8hdyDzpDzVs+zWzmYkymBA3FfCL/NsjMGYs2iZc
I05f9Iw/7DQ4O89iddHqFqr8pLdLuQb3g79rpDLTFLZh1lEEHURCiRXy2EfiUz4x
tNZUDqUBrepZTOhK5CDOiXr1stzfrOwrGRTE39RnRw8c5RyQXG4sKOPN26etIXLX
31hFNsvJgvYNdSHqijVDp7t3EjVNeti+ZTVU1ED3eaW6jJTJvJa16F8tw3PPof/n
QeQWCy3I5Vmh/ppD6Dp0v7JszJ7aTTTzqw8uvSRkZqwY018SBgu2z+sUwkmOFE73
oXEZ1UADRdUdFcGKL5QwDIz35nEtCbqd+rAh/rOTfFrLo1RI15UFJVbqjpJxiCZp
A2/SNgBl9V9W8Z5u3KcdHvaeam3Pd9yI5bwrCvScZCArIdwPJX/Iw25JAtp77RcJ
688MZjmRVaxb/o1OwYTsz2cGEibWLIWIFEJEobRlDGqEXFKkPCj9euzLtXSwEnFD
X7SaT7OpYYHZJSphxWPiHii70cQ927rNc4WHV9+JbFKAYsLZ0VCv3C0I23lRS+gm
rUan3nsL+1xa+q1a4LxqoMzg9N2qyGDJRwzL3rBGLU0jPMUewqx8E7Ibq91bhVij
GHKtjaURAC3Wo1rH8gitpojBm/+TiCjGE/xRqjFQoeU8jTn3nWOoY28glwo+6WCb
oKQ1AC4eaybsedwH0CTmDy6m7t2FWxd+cw0IEbtye6PoggHViuTJPH/+ZAcC2q4F
zzfhHvOhm92MCQvWFX3/Q04btw1UJCErLyUT+ETtTQIrvHACH+E0C6bwV402zxuM
Am8hULO2as6rTLIztW2VjNLfd3snp5edegKqD7pMqZGEYxrCzIrcdOlMQOti/Fom
ctNVUzYc6IWTSgxM0d/TWhrY1ZUTpm0bgks+OnGRtd7ckKbRArzL7TbbpmCeaVsw
oVk3Oz6YaIDvmQXzspSQiSQrzm5spPxEijCdH0Mdm9/T/DHfsMdl1X53e9VLMVyU
sj7pNDMd0orDy+n0mvpf4N+JsNkBwkqtyTtysgTDH7XGWao0NsqS+wmQSTwWsfyY
UNzD94v+CXT2SgQtupvmTBhPbc5bDXcbz50rY8c1pfToe6nNldXnsNVA4iUFOO1L
uFbIBcOIRJ5mbea5ljehhErEW8xeuJAdH/efRSHEdMJ+Soc6KWo40LxwL9fggIxm
AGr02lPprfAsfySgTjHW5tw2zBPgf1kACXz7AtFkAZ8fXMHWwFl2gdP6d4bRNSHh
pQqPbEe/esyjKtoVre/OhRZea9N5BJIOt+zCZa4RIulHxktG7qMCAsMh0soLjsXA
qNpnFt7fVPlb4b9BK0YCTRTvA/pU+Yjax8RCxC7KPml9l40IH4Wm84uH9pqnqV7s
Fld6uujtFwoi30DTIZ2L5wKsNytNyue6c5lQGoyguS7AzjKDbTLlyVOln/ROCFbC
oBAHphKNpJcx/YJOMlxPhThRSj7wJXlptTsxcfvo/HcACEdGRTHRfwb81XERz1cO
F53hWENzKKpTAWiwGuxCVjhLxmetyX6bpXqNoRWYANgvOoem4RWNk/nLGotYTS94
D3Exj+Sb8L6ab0OGq3hjXFlclJ/3wvwNqsziwV1wHREvkVVaZnXrohh9P6jN43hu
G87lVBqTlXzCn1uNDB2E2SM8sjKjsMd8QTp22/+7tHojbfJmZnNBm/Zh1R0x9Uql
Vbc+KAJefE+CJEjUk10q5QZfOnBzMdO+TRaVbu4xRdzGBLiU22x7C0pi4/xhNpAp
YZ4FNuKXhkDzyIcNkh20S1x965Dl2NVnc0agP9NZcFrZB+sVb/NLGUEmW53J9kTd
pIwL2PbkIiHOOrs2opceaeqCXjvpxn4wUcJkFityF89ci3BebLPJ9YD8xOUsXeQ1
qv6DBO3JlfojAfbxbGzrUsxplg0n4ryEPRaG/d/RwBCr6XmmI1xMoaIeIhS4h0EC
mGhc+tQZKVpPBfT1d2ldqTXJnfu+qbh/AiaDq7XEe90NVB7qxiz3xq8mFhNwmqwV
XKbO10Jh+p3IK/axAiceBmiKWWx7qePQl6roGiiC/rGslYI/meZKvTVn46WX2EzL
NYCMXFMhGsg9CPjkwAMGdBWYMLGZSDeR4yAFBCuEc0SwBAJfW3gjn2GuP3NcdXSU
+jiruo8v+DB5sCQjjRvptVy8fczHj7YYXn1DiKDCwTQ6W2Ioq/v5xyhxwDFwbZIs
ZfSd2Q3hbcj8VVG7mS6R669vaDf93zwigC60n9CbSA8IhdSRe+6GAIgmPn3Xsa5v
5RoFSKKd+31/S+N+zmKPMFUSHleRCbc8tKgUzN8ni6Ra0gwSNxB423v6ReewenBe
zw6s9qIiwlJbmVPML9GvGHSfTVmIwAiIQvjCyyQynd2BSDRi64ydA7uibSrK8o5g
fWSNyaFQo1oGNXlZ5xTSIROz1ytqNBin/1JP39tklwxr56jQCqkfTWQD0uu+2fsV
YEewz0lxn+6m0yCa4TD5YvKr/BWA6BkW3PbQ2+NLJxHz+eAw1OJiAKXCtRgAI17f
h0evTJFOkp+UXaxWLvVpdwF8E0BtjKhhSjSJ1ntjZwyXuHnPCi8Mkj7djsuY8/Rp
1RG+gRabZxIOq7ILoEDoC/18n1sptUsNSCNasaAiqJTc5tZ6hX14z9jplXMg8W1C
lSekalg5WexMudLGUQMme8QK7cpB6W53YdtqeB/fAwKz4OKlYCtVuP489k/HP987
hdOftXExrpbM02CpqZiFeJ7ByVteVdoj+NPkdxqOPr7Ubg1ITnv8ikVRY0KuiikJ
GkDavzByRqsg4KIVZjzL1pvAsY2ILo2LZuVC8b+gZczn8Wu+uj27YZLU1JLiK4GU
N9ModCCszH4+baBx8Anlo7E2q0woYBhmZkneZo8460jcqQXJbWARHjqWsWLua46v
4s/ivaqc4EQcr/U/JcLG4LjFDu6SINC9WyD+soDUERMQvlCrPxNePD8P/IAf2Lvz
8j4UAVFcAWg5oftJuIsMA2Vt3yUMjPGB26mWQKtuEqMknuKW69VJ4EjbetrRP7al
VtYzEDHqJbnbO6Kq/t7e1HTUnpflff/fyJfDwt2NLuUfuWW3IHKxDS80Lr03YGey
tej7HTYWWaRQFhl2NAQDBsHPXISLf9K7w8icE5LzyzQwFx8bMy8ZD8s2YGhVemcl
w59ZOw1BV/1ic2bvp7MC+r7QBi7LWAUtvw0FnJ9R9uxbm6i9PHB0v5WSj0lkBN7L
NbP311VrsXbQFDcoyu1R5xZQaHecrk51/Ddg5VE2wt5KLBcktCxOQLnHO3M6OuW2
AHQWE4Wzq7mX2fGIAObd6hB2ddQRzeFWH0ntGkW/JNT9fjPhs3x/eJa9JB1lZ6Um
/Zdz6npuqSfj1d3I7KqqkUpfr0em8rIzsFzZx9Q/wyKNz3rFzonulGG1zw7j+Csd
CHNE7N/O4/fcrjPBN7Fb/krhp2rsSeWc2/FsQ2As8tkLU0R2aLHxaxQzmh7WHHQO
cm0F86aORxQft0XyMKKw/goy5hTaR3h+T5zk3bKvUgZniYnNLCUHcWoNPeNhGOCx
NiwBwhmzXN9mkjdkn4OyyR3/hDR5jmHuDlbYYg7BzZmkoz48Lhyd2Qc+6g18730r
GzJlmJ8/Efk+bKm3tSDU2Grde//tgDoWNuLK0f03FjbJaVdQ+LLxyNPAvDMNHsMT
yvA2QddIxO5/6ikd4XUGMZ3dHrD4zoULWQqMeEfK9nAlZBRG5cnWM3MROKY0+L1C
1EYb/C1kv+PdeoSy/pPtYug5mCzzsUAQ1Z+6WeiC/Rm98JDVhSwgKuqeCa+xSn9j
ak0iTxNYbZhmqBXA6A0uygCTWFa7xSBB5TW2elqMhuoe2DY5WXwnaUpxbk+HASBv
hXVzAfz6G2S877GcqAotuBOQOWnek4fr0MIeWCmNers0bNnRnHMYBOuaqUbmVWZz
UksLBORLpvoOEzG7fT3qU+fx/aGTw4gV76xBsaP/p3CUw2OWO/8852yYNdTQtSpD
yJ9084SBwSqBvDAnpocB1fhQh2DZeGSaSiYrpmk6Yw/EO0xVB/5X0pkVgJKi35sz
lhyOgogDMlFg9rD1pRZ/BgpRYPYDKUxBcUFqct+ZFrlDTB6rI7v1KiAtEElyF8oz
5Ii7kzlySmwDWR+CzHiLYkxKhKbU5nk8gr5DsZZL5Yr5NCpo0Me3iQ7lOcBpB7nM
6PlSUdcMGVGdjp0HCCj/CmooRtTW5sp0Jggl9JBAPryrDbupRELrUvUfCSHJ21SY
AdrtxOCUWnOHUneusXTnj8XeP1smXxZg4l6zeLjHXnSNI3LcHP6nYp0DJpW5NZXM
rVCP9wuqK+REVY51ocVkUefIfHolGoDj+1Ogjwt9rFIeadBJwseJwEWQxrP5+jXw
b2FM+Qy3Ij3fnkbvITGPwWJ600gW8DP82dP7w3+fyboqValG7BN/SczTkKEnhcqW
ICb15tFH+VKGGfwn9cN5Fu/uirosRQet1It74CBAnymORtKLdGtThf9YmOnYp/KQ
yShux5j1y+nG/N0FpyiPGbM3C0t2r79CdgfyOk2x2TvaOl6nGw795UAKikRnNdJb
h7XrI/qV9sMBQihYhcMGtAXXWun5WteuLsdniSLDu5+0BOmkNxvBw9kTgpRhluM/
ut66mLT9V3xFaZky0H06TSz/IfW2VTG5a8P8xiNRft/ANTLywqihBdSGawzD+me2
xdPxtL093FHzomKJ1EYn032z9kZoovgpQCo5XPUgxO8ErRKzZZ2eoFF9tZUL4t52
N+5Z7alT7CSKQ/uKIR2rqG/kE2y1Bv/GNi7M9ttt/wv+kCER5FRriUIl5UWlUTSj
fzwVFedPuAeWxnbLK/24Rm4cmd4eDf9ZMOKtWhioXchG0UYTZ9/Nxk5Y/VIs6bla
UmvYKbgYOMJziISN0idwvXiFnLADL8hW2vCdGyGir+f3JKSfJaTP7gfE+0EhOEt/
OdujfWZ7Oie73CEF4WhA2Q6zTJ1oKUFm0rWXWLQa9WcuA8GZ0hDB64yyQK5XaNa0
FQ1i2zeuD1QKG3LCaU2CmUWxgiAm51T8VyD98Z5ENAlzj/0pJ646CVJp0+k9Wyd5
h3JJj+3K7cNvvOkicoZol59UKKX2MqkOAq7a4JCQhjQdlQvgEkbGHjOT58B0urvl
bJKZz59p/l8asPsWglEuWtuR/i+nHpPKMGhlKtkogJdbU1h3rqQn7iH6LiJBjNLJ
r9/V9ahDXOXcdpo3GG38PTRw+zlBHTscy62cCtgOS7oylMSOH3BNq6q/K9U0PtCx
52y0L7VhC3cBtOxudqOzQT1ULESZygt1bUB8P6XSaW5K8RMVlyYb9G/ujyiFKQ/B
o6zEcfJc1eRme9SRsvoMOJN05ShW9vNTSj08jabdXVJyVEbZLd2oTeCV/Mgc+RAs
G+FgYIQGb20PX4B4R/tJVyOe4Mi0iGc0tYpib8vmq/c2SxUVKPgjk5VB9WwidO9q
btWUNS4zeCqjsuYMHCB/YPaKaLPxFBqDAz6s//cy8vRlHulZ3rpkYyVsJt40NJFk
4/wX29FbUe2kGDdIp3TjgbzL8MNxqHdNPDc5aThFPS6m9MSGYTL3sEBmgbhLr58Z
pdmNZVX/Bl0I2SXtmJHwhcbxf/hNsFt9Or+pfl+LCxFvMPlIW3IRur5MEAfJR/tr
Ow1p2CqucvflPniefw8aspR6gV8d8TyHHAMKWu3YSAhcWl/oocDD0BMNFqOcnqh8
uXF/nUUXOcT19Fa5nAwNa7OAEXhV8PbaTauAosaoab2Knkqgj4d6c5Hjv/15J9UE
YYXZbuFghEo/tuFSVsBXhf83EPrmY/SvxWDgBqc1Ze3gdloP4Ow+pmAXM/nVtmfI
yZI2yVMwjte8RP0P2djZFazPzul5mFjIcGkh9SiWFqqtqvP/1nl92DbBGVo/izB7
LbZ7P8NQMX3ohyEg9IlsXB85jcCRyoTBhD597BFPKo5aBOAmZdDjXh0TDFBCPyLD
dCUDQqcKmszY3484DryWLL4dbvdC9jlImEi8sysoKAYuVJYSIOcRHLClAvbkt7Vz
LHwZHhDN2cCQyaL+V/d9N1+oivoZDCluGUW7k6JArQzPw5+twEl4EetxU2cjb8xz
14fcW1wHQw43RmNj/YgDy5XpZWhXctinMRYw0IcwvIBqAk6YYdZNv7LSKyVJ9rIf
5EKazSyErwF6MxBCumdFut0UUs8CZMkyNRwnS35BJ+nsJPlgoUjSjauwDoedXRMb
J60gLue9D7/g37rjqj8HkGobHmY/POrHsMytwyTakPf6Uxv3aSU5ac4G3cTvUOaN
AY937fHBWM+rQnV/fuLi4RCsJm92jzFugBNHbX24/Hpa5ktC71y8e18vebRQahSI
9uFIH81ajrZG2X9QMGfGWa0JpMuQ73al5m91kcaw0d+i4KuKfG2PoUxMp3cPIbkl
498N1ZVLysA984kavoXd6lsaQvJMeKdv/f+YzeM7mWBBJf3Dl6+mqeVgreh805ID
zaK8D/YcbvnlC+hFqwy6dGvudZg1iRu2eQwq0LHjFBtbDT1hXoh0olVZHcYvZR2O
L65IpPiI6aZVHi+lPQaiaAnR/dfho98HKdwjbRdhpwtIWwZCAR+wf88kz7xF1UPm
HOlrOF7BceXkN5s5MvPh5Yafu0jaKtTlAHRGemQAfsg/Y1e4IuRIa0pqIgF82IjC
FY8GfMeI6wMIiGuX0KN16/+VMgk3Ss4FLxd8Kua3qOkHFJbbANxXKxRNBEeONYE2
GrBW6mbdizbTT+FmseFbcbzPWHyhoiaRImGk9HqqbPRG6M3xt0M03mRWo2wpK0BD
MXp9VcY34DxdYRHM0OgHvrDHNHeC0MopFpRoME9mykXLUwS2U4Esk4/AYhLnmip7
EAK87unX3eSbPjufxbcK9oyWgv/y6p9QWb7ZiBMEWAjJn/qJbulpcMQL+pDgLwDb
xedBrNGUvTTvaZ2rMie9Ug13FAQ9ju6Aj9ZUKTTEhMKm65YbBmjRkcRQ9ixnCNBF
6ShgWAOgjgKvu+UIymxgdfAceovsK3e/t0pHWYN5uO0J78BKhYG2pZZ3Vgf9kFmZ
hvT1JMpUeJAbL08+QKb89YLI1el+xBMjvDLBNXefgW4FXx1fEahZutt/+6gaVWPW
C4RbXoDCLmmIIbBSXEYPC1oJ/Y2j4yOVjoEZaXpKB+KEJbdL+B7ihi5HBsAKH3Fq
+xVRYrz2Uv0ciJNpc2YcV33x26UPSU54tOqTM8BjdnW0iN+1al55bbAI9EUMJcSD
mVYwCsMrGiK4aWA3SWntg+i0avf2c0ozj1yrZ4lmSQFCRA4OozPtuH5Du3joHV7R
Gr9toe/2GiXceTp3X7ms/vR5i9CszihGMHAZ9Hps37JZ39DzgmzBsZTvNo75i41+
AK3bXyJcz/12bex8GPd9wbwkCBcMAo4BZ2XoAsmKTOP9ZvcPbkIy1d2bO5Czj8y/
WtxbYeu5eAZkBMoC9dYcW+9PQ8Ss4rnfWrbODJ8PVl7jIKkRaTtuGiBO2Kxe1ruz
io8BubSKu/qIxI1HcUNXCjMBGUS8CKvf8R0iKLI+rb4CnfLmRIw+tfXMSoJIOWvx
/gAMZff0jWxGDzW6ZoGWPvAJWuuwmBYbooGHKsbUptSsNjEKyc+mtTVboF7eM9nj
m9YmjfEwdjkdBmzeSieBYCjk1QBb6/asBIsL2mkXT1WWYOWIiy4VS6N3cLBXP+QX
MY3MkSx+nM+xkGCyl0MDcwde8vd7RG9w4k6MlhULNmRy8dk5nyph6ijxyViLgbsQ
ZjBUbPBNjkvc3LXQeC96mqHBJqkzUgZ3c9EUsTecQn6aH7fRSWA0SKcwir2do3+y
a3cPs0qOqncT709mfTkTPghcgStjrtIayXXr0qLHscpycLPU6EOYGOZlVggKrGGZ
iACnOhQtUiAdFiTjgBjNdaq0geIn8K/cJUT0nYeAB3pzstXVY0h5VyuHk/gzdsE+
3/OheWyRaUqMO2s2TBgOgLHA6mfkPZf6Ly5g3h+DbWhoZ1he1YsUkRBtqaBoe8Ij
FCWc6XLitlSs/SscBI/1VGzuqgheFCRGv/5R3HB0RhVFX9k6Of7mQwreXnI54fF0
xioUTgoBa74201Ea7odUvseNQsA3YnLj6/GddYtrIU5RDerszd+i4SLRX7EEmi6s
2u9iFl5YDCpD7s09uDTds4nczypCoPgHm2ibyB2Y9jepArVSgPAhmqU8zn2dUCGy
guVSTBlBvnvti8mcbjqX7VrLqbL6dGS5v6RvxnW43/jZhBbaTWUS5Yg7J09dTT3F
g/FKNzEhiH2WtgxZcHJ8C3p5ol3KR0ohkwctfu/oXtCYuL2Ep5t3Ol93lYp6AGVU
3/aqiDGX2YTWjUZF8QRptL3AKf4nyLrkMLT2ZC5XJ7LjqKXB+3GHagwo75n/7SO0
OaXe8P5Y/5zdRBvAQRY4Ormp/gzzOGAQ4vSOBsORIVPAA6963APJinzIIFC7Q6RR
LHlKYtI4Aexqi9/T5S2GHxqi3WBjaJtWkIspBTkosnUEL6iV6Xk7/e5UBr+stlQ6
KjNM4AEpeGWhoql1ocVagn7FZKgRmj5vhWjot8uJ9OpFU6qHqpMEMGnCC49CJw5+
AhPw5JFxfSiEiS8GTeINRm6xbYZ6D+2qdUCzD1OiAIVIU2yYHFLI8Cbm2STvPVbQ
0fc72qldKb3NRGb5CH1BD/NMRiDhjcZ28IPG0fCX6I//aXIedxujc44kSgmbp+Vu
8VjHTr5W6CmkUOhjSaRACTQDc6uEM8HrCpp5i3JKSpN+W0ZIYeS+tXPt9EOa+Jl4
a38oBCcsfzbfIi6Du5tufrCGFadBO1x9Fhm5XI+N1676YYeYt215pdmxcGdXqacy
poSkeAkGi1AO6ugyXIBO1VG7bMgIzXTckO652ZAiYWTAQ5fDnl6Jz+O5LwaFS/QZ
BUftBrWQ0BNI89lPG2fzzxS9itvvjmaOqIDNeIhGrOC2tb1N508ibqqPXn84dbnh
JOZiA5srbUUlizzD6+Y0PFEQMAyPtx+gKVVdU7gVMDxbLClJM4qTyRFZ9hOtG8nj
yYQGFYRI/i2aUDxmrYYTqLWGk5CNThIE8F5aKEKpz5YzBcyr/UIVybJ8Iy2lqcDn
LnfHGoSJISoj5i5X6VsKwJkrhVtQYzeH1yIFekjx244z+1QSwCY+1hwLP2aF3K32
aKHbOfiuFHBgq+1wKFmusZPNgmaAfpNcbYmXVw6hoC5YIQtGhbbziYAx41fgD+wF
1Ncg4MSK7JklTLp2c5GKoFTg7/LrhZ369fvqCKPj3HvbODdq5pAhkVYLWeE04+yx
5HXeLwKTOO98GmTB3a9Trmpj7Oogh/cbpkXtFUyaSJxps/e38vmC0vDaS9sHxoOU
1X+eIu96KyXDjja3XlJKgDlAd2vrQiISGubBFuV2GKu9Pq9ZTc9A9NFx+lYCfrNr
SMGMSDr/u5DNbEk1yo/JC4HNtpVsM8jbQmFHA6GTt4Yy89DO/6mDWpeNlo9bVh/s
1i0WpmX/Tjs3Le/HFPMYiChuLvYegKEyLE8o3h++/D1KrEnS+vXijsiVHkz/uWkS
GzLGxz/FyxEJm4SVUtZP0kkhKiOekOWdC+MLlAhFLoacrzNBQTfOFh2Q/XDA5HQh
gASTa0dW60SrtvKQt4TBNUAygeFMizNgaVj2tgix8HrU2MYQWnxoUjxFIE+afO9Z
ChcJkqcjhCxddOUHm8ZwtqfiRNKRE/Tax43IvnS3NhfNyx6VnJT1YwGt1bzMntkT
tFUErZtMegs8vPd9TGJslyHDb1pFC784jTvzqw0HjITWvJzGM+KqxENLBc6E3z71
WtxJUHB3450axcsujAZY+Eq8Vr/APGabsYHW8523YlUvVPs6JGOzPiiMpaiIgxk7
IwS9VY23epSLnU5fCa5kUv+xLy5SKpM1/hLHBFY+cfOxhWMn6jVRiTwxL/w5AItG
o2hDim7OAiT9sKEb+8r93yHocC15e4RYQdAI53uI5fZ1iAvK7FsYxEcXpTizhqd3
chzcLPOxF8RsEWONu4WFREFZA/sv5voSp3SDMfxBrDxupkiDNXfR/K3y7smpuqU5
qQnNqpNEIw6FCZOgjAyjD9GwXTZ/faY0LfHiL41QI+QYH91cXhnDYagdyNrjiqWB
VawFN+xHGrivz6zBaQas2iog6pWGdp8clplYmVwICvrUmQL2tpQanx/PPaUQrQRZ
3+hbaXKt8fpRVB/74pbjitw7kw4SwyCvuIT+5ly/IQRXU69Cl4in9xjPf6mvkgu7
1WR8vbC7SeoR4pCOzzIGg7hRB4U+Fb6GrVmILCknQkUMPGJl8A/pr75ILepTYPVL
NTriF52DYumeZTzW0Hn4EntvxA2JTVxkBiXDV1DfZ+YCC71/VCLdqla/wVYIRDHf
UeJuM5BMCfTIChMpXg+UR87vJectbRylbbywW8uo4GDhA1hTufvWFc8X85KFiGV/
HFqcqVc3efeUlmUbgNgXcetei5CBpu0pO8pnxk2JOcy8pCsPe8zil+5Ftx/Q2MCP
+NbPzIkWlDh334FqXVS569ePiUnT7FESsXFczukgAhUXG+zwG+34NlX/+J2y3kdK
niZev/RLLk2sGh3rUVLg2o2cLwPeaRwNqu8ZNJHypjbU/EtHHjXawFix8l6Yzx0A
dEaDd5hh1Tj1pUF33IgIoc2H5SzI3yZIYaUUmJz+/2X1HKMRYmFfJT6/9ZnsH6rj
XabjGKe3UuYRvIPS6opFIzhmnzKhhngMm6alhZHkMiJAFgSTW2xgvBN9hSN/jYwL
CES0en+6I+yXFbxqj9qTRYy2saP30YXwFzvxhJt4zfVsqlWEk3pP3Mf+shLG6Dzc
MxDn0A1ZOa5YZpPav13AI9vi3hHwKqYKWLrBDGKcCEwCw0Vale/i72heD9Ocjoe/
bgzG9VF9aZj6bM2oz9bzrfunZGkw6u/wLCuNnY/RP1OdZ8pF6THvThv5GJ0E1Yqe
o1a7/nGm4okE2DRpxd6isY+GjSS0SJ7B8/Rlvq7vgR5mg3z26NBCjmb3xWtPlFdZ
/8nahDGyh42MTsI4ChZVyfshkYiLhdrCWMNwOkZGESb3D70LLAko3/esqpX5wiNO
JqdPYzqY9GUHtOHihlQA+Clj3sOkFSAM83y746MtAb8PoaqIC5p8uNBai81UINgJ
qvquBdEIC2BERTpTtKNM7wrbXyrwQzgf8FwTxNWcyJ7h7eKzpHe+qlDfVX5SKTE0
+wbWCzBKKXxmVihLw9pjki9ylVhVdixFs46zzGjJ7EzDN/0BZAutpbVn4N7dE3pH
13wAT+H1c5CSWkv44BgUssqfZgMTVgSqmC6qnoqciNa2SdnObdu4Dp/DfpXZe8fi
nny1oRAaYRnzGTqsmm3mSInP+4a2JoHseF+AGVzrPtrvMgvqlqWQOcK8eEhfntoN
+pGBQpJOzn4jmTr2OrypKw/LJKgWJ92c9RnFIo6c1L2VCsp5xBMt4/JsDs74+c+n
UdUVYz3iQ9gDTqiTI5mRv3uHEFgDFi4XZOvLDuzPilEW2UWIQatiP2CZjqh/0BBo
GdemJnUfC4C8HlL8dPyv1olrS75MoasKmKwi/D6SR/hX6tx9D33afpPFVSM+05ok
tWA0IfZ02bhWiD6RQO+aUF6i9+NSo7jPLHKDJeOMPJ8PQu/4QZbCwqom94Zw0uDG
M3DwzHr3BFIIabX/qyT0XOLAWNC1j5SHdrjKu7nQXoNS5OFTo6Vq9qR6gea5z+Hk
uT0NZ6giZN8u5Er9BnU/gUpNgX2mnOx6L1F0pNXdv6fm3hFniBnvEGGlyvvIKE1m
jJmesi6z9jyghE6S12pcoJAzese0ghomAVQpDMbZOpovTc7BckwV+49StXGk3gmv
1F8ATF1uKq45H5PjwxC1WQGGId+Bq8xFUzEe+8lRviFRgBTmLZNX/wvYVOqKBZJJ
PsmNLZVGibs1mR07MB9SAWfF1MstnD8svskQqQkpuqAx/7d/uVaChtJsvlucIyE6
xX2TmSbFY5K+Et+p1GLzt8eFuRRWhh6OfAi6vvW7b+UWkNmpQkCVexIaiReCZzTo
N9lqtBRnHWmcax4P7awLPbMKc+mE6lgDdZ6TDKeeUFxPC4bRPxUh5f/p8Z62f6/+
Hmsxf6NIH5I7eUoCyazAmueyE11LvqpjtCXHlC26mVU5B9yfs1PfIo83MFFpMrd4
7LhI/0FSdCWLG+N1gY8Idw/EFBxp9hW5pZDdTom7cAv1t06DTZ51+1BWZRsnrTla
vfhxnEFEg0MeCB3ZFaqkOMUaq+M3i2Q+uhr/a9TPal3bBi6RacE6QhncmmDMYQqh
Y8wGkM3CZyrocvnZJtF37JWKkFNRErSwRFSLj5ApWS+gITK3zKtm7qdBaWcoYRxy
BnpEQ0Sb67uMz6m40tYfdnIUg0NyzJ9c6bwpZsZT/4mtjfnQZcEsjpKI3o+mycCf
ydqU/ifV/+qiKFXMPjvSzhD803WZWdrPy+5JovYfFwq3ayuRcCgoOVt6PADlcNik
X5sp69utP8p1VViFRXZ2ZRdVgVjNdFTTuSuwBjEyUq7zRqxndruw4dSoU3P8yE5p
NT7f082ZCN2iYLMwiCX80+VYtlWtZkkAIQlsoJ+Rn/nsjbQkBzRw5Ib5ToKmW6br
qPsMEwnRGSAhBZe6nc6u6ZfyYRmsbA22DjwMDYE3GLk2l0yayv87tvlFPwJIDB9Q
dCKUijfE4lfUVhh0mtsecj1SqIY7QHzrjyWCyqxxIe8pM8R/LrJSCNI3rnj2r9gc
F6qi4qPEVyQh56o7VncHCQ5+KmUkTCGUe1TBcrt/R1p3X4uyOaF1PqyvlSaxA+Fx
9LL48+H4O8duBVH7ZdHyRJPOfmEMEiCc3WE595KoO8fjvIFQju5Dt4jgnl79E/cl
nPpdIFqZQXDH44OW/wwQh0Hg/J0SA6g7SHPK9ELVLYRBDcdRsxlH+O0O6gzFKrDj
jDmOAu+oS+Y+sFHPCg06CFdHCLx7ZNpxvsbJtp72xWI+IYNSAJatIHUIr5SY2ng/
kc4IpApaX3zll/qbGuGs50K1Q44pvWukQlbeQn9opxgoAD9WF5Kr5p3Ugl6hdDdc
WP9q9yAsZmQ4VB//qHPURLL98gx0HOHjBneWP1ChXKQJ2w1fxkIfaXQM+S3rruqR
OqjGI/tC5XEuV/N5+QA/0AlAWs3YWcDMVHPYzSzSSrcqRW1Bb0EuYP/2+0ghoVRA
JpXgXi0b44NOVUbg3bKM9mFJp5hqnBxvr1eFFuzQoRp9SFIMS9yNvO7E8DXCwycC
ZHlS+ETo9Yw4e/IOCDgYpX65z5nkeyTGD/Oga5I+BQLNfoLc2t79t98Tatzs8hDb
xXf4jn/hcnHAu2ZaMryjRtgRHs5yS0btFdNlLpq/5ZiZqwBR4+86ZtXEu7pTJdQx
xHnvpoNi66eUlmqDFc99o30xf5y3+Mf5i4GH6e/P+bVJ+CXJg3D45oQNxWMEwQcf
6MOBrneLCfu1KWI13OcNY+VZDfr+JpfhE805Jv7RwTlMx2UH/bswSFyY870yi19p
6kikd/oMtZuEMG4vX0YeF9GGiFCNJShoSLllVSYFiuFJ2sGZrZnNjvnnM7DbSCiL
i3MncvCCOf379/dQ9um1yz7ekaacUnFL/xk+o3yNjGkzO15N6KANyddykgE7sQs7
BRDM9BADlAkacXwOEd9XfyXDRSpW9aO0KuB0/cQ51WOapQ6PZZHBRRxEvYAWV+gy
ovAD6yzb1TWQbf1UIBjZvuykj4NFhjghmQRPDKm++y1yF1AuwbfPBnYLhinsj38m
mpQGNDfNM/eOdsaXN0TugjmxBfS1wCqIfRDImCw2V7a5xwXvN3sSJqtj9TFgEJSn
42uaHjOIAxQfvDjHqF/jfSj+4cmQK26o1bySlFvamrCvpIA7Tg2DvhrF68hPmfy/
WfMkQ8GxedEFEW+UNYwTr5792vCAWqVtIvs5WDnBkEIQM9whcjqn4tlHCDDbquK7
XxUBorObIJyLWCzmHEnLLTKSRko1NVHICbwVl2b2Ca+JFE/Ckj0qY1NGb4ysgsDp
wlcqnpfXQCbDfLdOpvrYr1YB0R9oAHFxszbIIx/yG51q/ThlxOgC9K7qQgK88732
gXjXarUPj6HQwk6NNmlH/XzJ4xgMyC2tQId21u7HM2+ChKJEouOZyEpMaiQmIw4j
LevxCTMUM/uthNo1DB1ANEue0exEgbj1D7PVsb2/Wo5K+4C5S2dtukAbv6g7aIKt
HOlwalXGX93yismMh+f0rH99y1tkNN7QQuZomdhIMBa9LqyA5CrMjP7iBmE+O7gg
s2pugb0xIDZninLFVWTGEH1/kW51hZk8UP/RESMb3wGEJBspGpMCeNBQTz/ocOqX
eCNd5D09s64y9bfmmlzA9I37ahQWAuCKUnalQMqKPutSO6IimrnPNvbPxvMGnLMQ
8nRGf0kp9OFwXaRh2lXbKvTGR37iuOVXkuKtKJ6XQvdO8Ndnve3sE/E4mtJgxqVS
rfAHpOT8Si4+yPCzjsJZZpzKhTF9zdiJSkPOSo/zPUpRG/wnaE64k3HPyp/SB4Ds
6hwsY2GFZeQwZKccv8mn4DGnhyP19kAYsPBLwzDYtAebK0b55Q/Tfs/PMDMQkOmt
hvJEqwe7jo8PNnsoxjNODywyPLokIcDjm59EnpRgk7gk+d4dTgOBs3dhRp7/CN0X
UrqylsixdKvTIVBGhLtmhC2ahk+M+m8trh6in/3e/pYztSaStJO/oPbeyl+qceYO
T7H7sGIOhlZzSCNbLvdfHukLLXTEkHNNpVR0Yb7Yan3Edc2gcy+c2iSQTWFKVheO
1arhhW+1qPtVh9xB15tkeu7diB/jSsC7lzC18wuUKKQZZAW4fKut+bFBAa1A5XEV
TxUfH9LhOuBGzXTbG5NI5ZoISwYOPl8udKYSPjUc6pYyg/jBmryXH2SRaTt1LA0/
h9q3MukjFfRsQmApdp5pJQq8vZ+XUY3OaPSiXdQ9D/oQRoO1jgZlDycTekD4HbZo
nrX2dOaHfW71GSDvJ6lgKUJTQ3kMwamY6iIxWC+BcBO50PcldRxAusnoMY+THC4K
Xe5sfZktoWI8knLJOxpDjmt8ArE2La1ZCa+TjbboEhpR+rJOB2srfBFSV+h5vhzV
Tw3VEK3lYVwQ9ku3pPRCLowFSZ6UKghadeW3OOl6tacHYHDIp4gLBaLgQl0uKMlf
cwpqJdiWNUNxZ/PuUt8JZHHLwYG8QsGuB3C3vLs1GaSG9+uOVrIykjTaoM3qDjHW
y+XMuhOqvcNM47nS4iplCTtKmWqPgVb3UiG6V93O7FvuIeSVd+ry4hUdlhfdED2l
O5EA3pOQGxHUiZv69vCbki/BxLDGOoE4WG8OMLZRAm4qUH3B9ktRu82GetOBV8rH
9iuCR6stBFSYTp19draQ+p7hbihCKRKAg3mV/thU4WrmVetHFosEsFacF7CUZ1zV
izA9o4b1O2Utz4ymCRIotJy3ODswXNGObT1pSKHzPnFDQV7ig454a5hoOhmsoTn5
UVFqhiffZCxz/dbFr3kn/+61aABYJBcET9h4gJ++EqCxVXb4xR7u0tG5tLF9Lf+F
JVYuUYKlbw2wCX1Bm1UwpVKcHTg+T0RoLhVX+CIx0leP/BCTKzKe3SeXBZJoP39N
U5y72bld7A/gSCJk6hIkXtJeVTFkqNOZusk8kThkUDo2MMINU1BL8WhgXyToglrs
uVqyY3+LWWd6MqIuY/jTxtFprEN2P1wMseWP/x6m7PDlIBLy309ALEIiHRmoxJwe
OreCI4fqFVqK8cMqbzlL4p3UbuNyxXbLF1iMLm+vFqx+FH86kLf4gCWdzIkW2+kU
p4ZrFzeBI1t+kkYNPtkk4VhLWjKbdzLbcR05e9qUxQh+UCYZP5ksXf91kFvAkLPB
/2Zu5vzA5ws+ZT8Nk3eeAvBdFlppBmzwSPOLFASN02rHvbQW62W0KCvsbVi2x7RT
OoqlXWJeNKVB7CCVQH7k4cKM9KsQRd723gQwFVg+K4Gsxl99IR4y2RM6xtXpChEu
HXd4WpUeYeys6hunBGP3ViNtk/bOH6Bto9qeGmvkkuOMBGhemk7mZzFGHI5mRrd8
LjatHQrf7fI0BO6z9g/GtcDPwfE8ykXWKR9cueg5mprenY00JIdkf/MKZukYsxlt
+oVYI/nVr0qoK6gTMC83nMVPAdlLzI1WtToBswF+vVUq3KIp0AKG/RVbYFZNq9/0
iuaAhBsydkOGwL7ROGb/R/9tvBA6OPXg2RLRYuHq25/8Nm5LdAaUDs1hxYsD8Qlb
+Cpjm7MuKfZW9QF1+jY3ylhSncYKPSIrQYvhw0vzf+5VyboLw2/VgSWwriPd9YpG
J1AqRujl218CloDnBu+rvG8wc1qYAlKyTxVPpeSeCxrhnUh44rDdagfFLY1XnFEf
sWu0r9t83s+A2Lj+pLVrp6qs7Rk/fwAmipJcQI2ZAzxllX+9UliPEqU3kc9M910u
LofcigHxKwOpAqQ+XIhrBVF0JGbvZcuegrHE0VkabYO4QVVynMohI+T595x0zq2z
X1g1D16IgD8p20Hk/moZ+dsIgsZFPC007GJPL8GVtUXOWc77Akew0M6yGqH/M5Aq
TusOnfD/bg6iUX4Xm+ilXcke6+SH0uLDOibZqNT+xPFIhwF0kac5omOaJNYau3Hv
YJnKO+HAXBVh4tvCYq7x3n523MlHzQJyDwUS47RxUF/GHiw61WSJRfj7UJsZVlx/
9Q1BDtx2ry2v3wlZrpJVX21Os0H/UgEPai92zwu2LpH7Pn5iWYi/bVVQJ49xfpcx
hjNtpdcmiFDQgu3MudLA5bx3qWLmqRxVOCnhJH3hYzPo5miu3GM1Rz/taBsGaAaI
S7u8+PN63/m72ppmUKK+jK9TXe6Ttck24HHM7DpqKBQHTs9a0vlcsdfFDwGHwkzE
atztYIm/D9Z/gQQQ+55bAJewDOMAzna3aLCCyXKcdqOveCORdPQY4W3lu61XzcR0
6G7QgPVjo8nlM/fIwUSYA/cBVLOSop1Iieg9nSN1dZl6o/FHX5DzTvJGZWClTW5P
ZC7ePlLW08AE+2s3n6H4mp6MLcxSDjwvALcUHuPieQ68/vE4B14U+v8XF+emnyUz
0t/P8MFsSKsqdl1yHZKmXgHfYOZ56+eBWQt4PfEYhh8KbLYKzYX95xrI9/sW1XLQ
dUSaWrFSpV0sPtsjatA5N1MlHNWrc2gURwBwO55Rd0+yXN2wFCK7R809IOz2KH2V
GHLA9iDWXXWz3/lmIAzjK1Khh738zGX33w8ZWZmWkA1BREGHm1Igq0nzdD4WSCoZ
kLmwyYjMU8ws/SWQkRhUNi3DAkxVA3rRjMeWJ0zBXHM+3IMjuaWAXyoWxp08k5uu
dZPKy1MajT8jlAwuF6Pote4wszXcBAxcptu0mj2pBPmbB8hRq1M6bUX/4Lg5oEJ0
QL/e4jjguz9bZS2MgPiKDDZFYVnGl3I+YEii5eW7Oq7C1KYMKJT3hmgATE2q3Y0y
WqvJQ6ybcpYlLafSvW60/BvkFswmk9xws7wZrG4AckBm+M8IhQ5hmHGDojkdWrJk
EvJbf6ZT+zRQ8opzcW9G4CM5/JFH7cjkXa0UJdm3+8EPHLVot7zS9wowXeP69O1E
lIYJAsrP8j0bJedCu3caB0vHUGpushDAfkaJ4q4kfnKEazlc3diIDv3DIzcy3I/G
dDdtr2E8y2Z30fkW5xjBBElOIq0S0CS181IMtc24+CJYYlfKdWRdLWC5DVWXC1j+
YaHKk0i8cZmEMzxOOI8dA3p0SWZsTEqN9dgx2iC7Cm/q6TnwX+mfIOJS/wsdU4ry
wY8lMXpNxVkoqV5TStRS5KtelNRQmm3lVChNewhDybsM+hds/dIA0I3JdriB5CBt
ffDCVQTXYa/XDtAdf5IdoOgWkvp/WYHVpacjloB3yVFFIycW2Y3oik5rID5/RxqK
cek0biwggHNkhTdRwFCqOat35mpL39/mx5w6JjMb+x7y0EIa+IXUaq6IfOnpTfN5
j2/+oiQLEIPVZABcGuoeM16z4AM3UqduNZJGgJTBTpDd/MgqOhdCiHV0ZUxiaNAB
FNfgejKDQa88YEvJxWvzMxFI/m8OfC0RfEr3XtNgikzBwXx6dnHhqPPDbGVNX9H8
rFHBPggol52pDaqrZQNylKJMAJCS5PdO/t33b+CuqjLm/86Px4827grokTnwRXmp
bUe/89FIFU+yUecZiGilwKKa2SWRIrokw8t6fphTbyWExtkE39FYXyTC3uVxgrrU
oIY93jp1rzNzl7l7M3TBvCucA8CAsh5RfZs1C7kvhpB5SuJsFnWNj4Czo/ipW1BR
18YYcdsIEgQfN+zlAsg9qQbnzMlnB0x6x+dUtuiGhJ6LmH0eISVYaxl2euwDA0fs
tRSfp8kkJbIE1BTJPVvrnQ18l9MOTuGel1+Uq835g8+8mlinnMP+COjeV4TdpcKo
C7LLapggmyYhUr1pUa2RAuFSrEkB3wpVtatSFEeV4VUJgqEOpQYZ60yyiQllJW4J
lQhT6JOb2AwWTXY6LGCKqY2cXw3YpdO7PKy3Qrty6A9y7jhaKXL6Viqie85In0Tu
baUZWLFN8SiDiBmbhbrQOJxcdGftySnQfbJ7/oTc0qbbzu4Hv4mCtq1xvsn0rB6y
0GEmdDYIOjbYdWpqRLiDbEPHG4X+Sd7NtdHoQ/21glb7bB2LCj3WJCtOMk+KHHhF
JpjemsBu//S/fkrPUFI9J98rHSGOTecKWwdxrOskzPUYeWTT5abzlEL8jZu4NLC3
6T8K1Ft3K67IvwxAnrQOdJZHGUS0ACmRQfgFzK0YpFrIBBRqlegRkWb59o2Xojtj
DPqc2+lwNPyr2ZWoUqEUTQf3MMXrLrtUMMKEiYIZG+J683qApfZ5wbuUQaXY90Z8
0O86vyQwRty6BUi+oDuMrObMgR6bt+DTJM2O4EbxZGctlU7z8neBa2NtvMLKunsi
MTG/7jIWECuBNQ2I3M9flI6v0oXO/UDSRj2J+2OqAAValWTqGJ6eTHmNvAbCxo7y
X9UPkCSGJW/E3KCoAHAf95PV6/q9XLtAiexMaGre89VS3YNzkXgUViX/QwzpVmxF
V6Iv/ys2qfldofyklWLgRmAZSSmjqx3AZ/NEhjwiKMYEIfFJhwm9FoTBOqVsvVxl
q4EIuIHOt9uAU285aEHgJb3uoW7WAGUzvOIG8H52xoaY77wiQ1ENrq+kt/81/pZQ
CzUPLW1Fg+5rg6Q8By2lJF8UPxIWk4nLpc6Bd11AmJ4ZCQzYSehhEOVWfnHfTCC6
NNoFHZTf39sHBVYxpE8ywtuIBVpSidgBj1/hweKd9KlEWjZgwkYqfgl+oGJjbVUk
sfMoi99p46qCh6YLw604frIaChdVZiQHYpW1I/uW1pF7o8CMcfXfdt4cRDv5K727
l7dkl/X4KssqUuz60mHcva4B3vVKiJ1ocdB0+OOb3M90L46fvEpoFgC6jaCnh+XQ
HlrmqMWqD0Hh8CdQ3rpbfjIhL9f1YgZp10/XuvZeVzOah3JdwGnP9K8RBV/dnzVV
foW9ly9NJKGf9X19ta2UdV2teSM7OI9nOwoG/aruoyxBMx8gbbUlQBRU6YkVKZXK
/j3rIF47X06d4JNrUdjaLx3QNWH15BvUgkbAaiSq3jDmHj+gu+xJsq/xuApUnLHA
mZsOUrFFkHr5eCWyyyy7Y1LW427JQRxMQpuIt7O2J7X3vAEsoyXrJsqJd/FVI5Lk
PsjZxBJ51dgeWFwWSitNAjCvPUrRGUwKiXWmMX/G0/JreRo0CR5pKTxkGV6o0CO8
+z8Oni18UuJUM7Pp8le6H4gmWrworaD+FDbE/qO+Cbe1ubd/nBEjDfTns9+3wHT1
6lQO1+Kah0KsAnyxrwB1cVyLFpKAyb3VoaOstjCcf5h+pIvXMjDUFQIT5x1NcoHJ
2ONi099iKLXbRY+327oBj4KpC5DZdz9P+lIHY2Ncp5+Pe1GBEz+1V0O5HR2loJj5
fqteOo+XscVPHy6GjRZsgMIHW/PBst0Hucl6pgFW55KWKhZzIFlxxrMfl98jfTnh
SOdU9ZNm/R9qwx0pPZNtNALEiQvzl3IgTLOErqB3rMj77mYI0rDAOSA3jVamvuQc
6ZjpAyLucw6AVuLXvguCLZs4JrbH0YcxgbDAV20ekO4zJjGr52q2ts/Euh9rD2Q5
jYkwRCgSLwIZaqHa5hqB0ZNdkPtTVXko4GBcz/53ypmW3jQCnA+w//hsP0WYx0Bg
LrAK2DbTvW4j7XBM35l6s2TtFSMiAtJOIPLYMOHofWpXReSnurMTbEyfKtOWFeHG
7BIdXklVU1kiWM0jOCxCc1KRMgF/PI4JIwECN5Sbyrs2iW75X6ZSSXpLDXAlwvdD
S+9nVZZHFWc+2mTAQBXUpKzyMr45JbHoK3mDLipw5JA5dJe86gfxzMC4uee57ExA
RsOoNa6RFamc4+QYYuYzhHsv+ydlgj6evuamfYxunNZRTBkvB02qnW6Rmq4Yy/oq
+R1MXg35pR4FXL4aU1TDlkCG1WXxadU9DtWpxy2RKkH86pDPoV+HlD0FaBW+W0T6
CbMm022eyk0jnoCMNCDD9okD2RnJJXF9EiELYHg+FcHLBHOOlpsL3oaNo1/H6c+D
LZHjDyCToiyR0/RJdfFdb7EUbAdd55nMlLppDGd6+SZC0NM9q0fwxnQFswlb/IQR
lpyeOoHp/yFop5vzm71vKL5OQLavVPzO0wk2gmEqx/DF+hCnQ2JrtbH3hioKAOmy
2pCzOblPG1rRusfbFKPM9b5vdI3xvch5mFlQDVD2wMMd+nztEd6GRBh9U6h2XgHZ
Xu1MEaIb1E8H8DoNrHzro4IW7ccReTyF+dnMdQBUujjjMMXdhp4T4CyYRHb9Muo8
5paOpeLOkUeBbyB1oTm+Qk9R5H/4LHUU2KBtU6fJCMHhHN2AO8XRlzs6EHqEsY5Q
f28EBvsT2+ErsTzq6VEmN8AVfKnWaLGsUCMuekVCjiV3Dq90hbQFmwqwsGUqNiLA
RHQ84Fc2h/xAbhCZtqXSqApJbPrFpqwUgAeW4L+05IyYn4FGyYbG2yhBsAbgXBT8
qWF4ZOFZebx5g5YxPmM4edVfiz3Bf9VEosJY9etS43Pc1CQ2AymRVAXcYk/D/r7L
S6x2FMEyAFQnYFW68k9aEN5psNUO/YszIvZ3K6Y3pn1bMyfL0CTOV1Oy3hcHQ/53
hv9kp2JGDtfVW5E2OB3xpMaamvbQgTSnPipwOQ+3aQYiWGMfkVANgQyeSC2ap04J
3a6BP27eOiGE4GPZ8006ZxmDkHjLW7KRzt3kY06FJ9tripk7LtBuDBy3IyIcKeSa
muLJNboakk0gwDdIn3WfQ7jmMft1YtvB5WDIob5+qne+IqdyMwP48sTkQS3Cjvwi
Leo4PODj+LjrlwX+LKWIrd6FVyXR3YrPPGGTuwZUd6oiaVF0ff/0xGEawC89RqcT
c8V07bxSwvZvmmAxihrdN2RantE/Z9VknGjxAwARPw7qkO1PZIEhP2cDHRoFU+aP
dNjrmqp33+tBdoMzZEW6X/rlAGAYT/V0JNQ9Wj4+SXZayJBvSUfG470jK9+8RP9G
njOMX+ia2y+e3jdDMv3MNQLQ5w0ny1uiTTaPzlZbFJu+98Icr3c9u7xGY1ov99jM
6I51ujI9qVXBm73SCXGAdGyp83VRweckleBj4uf1mNKXLvqI36OmlHZBR/pyloLU
KwIiG7rt7pPo9jJ9LMBFhOxaK5Gdw9W5pABlKXKrnSFKPC4+DGxFE3NG6xMfogyK
8Te81gcHG7Mxkie7s/zoZvXiLHDXqtO0MELAzWqmrv1mi7OL5uIeAawLGoa/OybC
pcFP3X51soDqGwMXQS/GPuoYS37RWSPz2g9bzIKy65eWTWOAk6Je/UMCOIS3oCuj
rC8xWL09yP/yOc/HnPCo4lG6Da3GEMKUzQOK4cvdXvbS3uicxWOP3eFlWElq8+Oq
YVBhvkrbQDZW0Vs2z0FUOERCTLmmIEzDnG1WvwJDQcRqKiJVdPK9v3s3iBkGZyPy
knpVGa4T3PtlnvanrbnHAgpbqV4XUomQmv6PHPYpmO5vxQ9Iw1FPLXD65byFPV+H
XzozYfAg83m4OYZzgs4TuYfuSRAUsPXwdGWWm5exkm1PRwTzXEv1by7F4gZnqNcL
YLC4iiEGlXKh6MM2fabXt7F4ulFLWjq2//bv1EISylYmnhztqb+reA5I6tGxWDmQ
7Ss8TSeRpphbxUE1DwmukcnQQvJcCxfavRVExdc4Oov+HGv6n5ySUwAjPgR4mF5/
GZaF/vG565qFn27kkRwFtII91xJuLDzeDnIbgLHGwQckH20fcCcI6GSPULJsXvgX
EfJr0Y7AFzO+xyz+OvJZZRrRBAcqVyhNQZrFAP98Y5KbcxLrtDSpkH0XfN98eGGx
aH3d5EOHDjURk2ZUtRZOQPGM/E2dpaaxATe7viofqNvbzRDIo0994+e1auspkItb
GfO0vVlBKfs3sOFS6K436BcVuv3T2d8nAgwdlBomjjPzuM8DtUDgfW5hdQK9dZDW
lZKuUDauIkmY+wwOOA9FrxfSZkfda+j9U8l08gURu5OU7/lVUFPTwRRRBJo6iE7m
H2aX1SjramklIHc7hb6TXodmaHSUrUA0RZz8MQEnM2q1gcAClb3JNhd2Lu4RMUos
3HNmhuDVKYlfhgkJCa58Y4Kyh7ZnfKs7GG0YO+hjLOV5PUarRYmdUE99NXuK5Bdm
wDyYlu1otYiyEioxJV2+9xdeJGF+xtg1W/7tCSxUeMdu1mW4Vo+T40di9t2tco7J
+zEjsykFPlMRKVIAjvyONQZ04rf3EhC9+jn7hxZ1yQp2o8+7A76KmIVfi/U6LAEU
XBs7U6vmUcDo80kcEmKnK7vfjeVs5KnhJL0dvrvYCrKM4TavdE0pd7hiyBHJZKeB
ti9m7OVGqIeNo09l4Fb3FiA5Tj6KL47Q1pKEBWylTvR9wMmsyu+2UXJkt4Y8JF1v
Qljm0R5gg3R2/sywgTyxGFbA8YaEwkWgMOvCBZmR5n1VMoVJT23Zaefn17/dQNYN
JmtckqsojS5uy5HO1epvc1YMGg+wN+B/WL3EpyZ7turlqa9zHFhQq4mBzKeOyl/9
DbF8jovYi2AqIreHQr9olfOEaceE601XE2fzOHGUjx2K6CDntAwMV84Wi/yyKJ/r
fm4NDtzDCecfIMmvIVjRxc+C4SE1JLHhxDdfEg8/ZAHOVLB882mlSC6t9jF66RMR
5XbpCXlD3owbWPwdEH1/4NdkYmzY6gXRkUttuqkes0I29nvohBdfKtW7CO49jlWi
CytGHUAUu8jyM06x9UxYtXOol/Dl1cDPQmnzN9OpIiRiBiIW2wsvCKn0JIaAXNng
GItCVgRykEipndK1JNb6TQSFNMrNZttwxoXQh6DEguabbKyJwBE7YMYdkxIQ+f/X
zf/HuW9kZCIsHx9xGOfJfqirOubLXTUx1/meXwpwIyvI0ZcClxQe5co7ozbHrDKW
x5RFbpiUr1TpMIL397y5zxuIKAS235N4JMXmIdcQM9Dm4nfFN3ZQF826f8Z5I0Vc
fT1cQsyz2Kjg5doIpML6NghxLNWOkQ4ZMqdW9jfuYhX1cBDkSPldr07ZBwXmz+Jp
yh+K4XD3Zz23BkoBGkwcsBMs2Z8vnvt1NWItN5I65gV+wZ4odPl2XZSIfqrK/6IT
/kWbKpGxHECSdHWX8qnAkndgA7g/7UBS7lO9u2jDuv2/uP3b46TtErmY/D0tp5SJ
MYAipeUOfvwXh+9LN7nsLThRuSqDYcdEOl4dTfsREd1Se0iMsF+VUJyx50SMvdqV
TkxjqqCmlHakZyt9Qd0JjS+y+ln+/NK4qC4D/PkFAWTecuRUn1eV3S6vB/sSr+Gf
KlM2aVNinYQGEqm8IJSghDGBPuel4RA+GzbRiVlLWkv4iECv3eEHFoUUafA3dY5d
TH8vq4JDFxL+j0n0YEXl9CpwBCGrsXNTxi57NMsJ20Kwnx+noSjxMt+kBg0YM3da
oTECxgWhcjKn/S9GrGBPhIJMV4NpXKiONmSGru3e9CeyiZAVzGEZWoy+g1xIoIDB
pRnJ3uOKQtbsuCzJHZ64VHvucGV6S1Nc/vYlbfjuYSn7jT3B/V4/e8P04oa+2hLG
iMmpiHgvocinkpJYDTwJXjO86YRrFSDr3WM7t21Ho6wyTdNgK5UjggwMJD8v6uIV
6ZlFxQe4egzKBh24wGrJSL3Y62j4DkqHhRoSDYk8uFvbatI6L1xx1+QoYTCvorfo
T6BhqJkPYlKOVkofY5aCgHvDYBPOzSrN8/PucX2+8XG38GO832DA8qDt5EhLV/xJ
lC3hGXBcQI7YWUtQaXHJ0gNzaZL9D02+AkY/F2IbOoWiBHooEZUAkqJO9xroKtBd
QCEQpAaps/2sNIVp+0BJZfKx7ewsaTEVvUY/489YHXSZrpSUfQCbN/LxwbP07T0P
WaH0WGFlVLHVqtGSuZlZi4+YEYamWOaOV8r4oB934koNQCmWjWBEcSXV8toXXi6S
UZwiXRAaVqAEk+8QWxTo8+ZmfJmsH/CUNUpiUkg0YoKWZszd6v1tW6Qr72tQaDom
RNeLkMLMIVFVhQhunyRYzk2pjl0JIvuPZONsaWacvWBCa6KBtot5P2uHh9E4sNKt
O+DhRL5xG68PIjgFN+NHR2aW8av4w1mRlPttBb6hUTREzQi472OvNhOszfIbzOEI
9V3+SYND4z6UgK8wH7OKrBZI41QwRFKSs7E0ZcqwynuCxSCRKfGqAfRcCBv639CA
n9kRRpMorFuzGLNp3uRIV4Il8CCiuSuaCpENH+J/SOJT72tbKMh+4N2NT0gLCRgC
O5FeYS1+de48xc9vlYAJiQ156exrfakQUprTQ59HRh2i+iDY7lPeNLapjjvQgxnF
LdUclhmd3qewVDAnVqhFtwoKi/3yrmVUnuwRPyKI9sjBSIeBc9eBDFgxCwyCXLy+
npSnHvZXn4rPi8TyZr7gIAeXGmYkytaiqf5++V8ygy4LD/V+x8gpAyblsT0pmjAX
l1cek6JlUXUFkY1dc9SMrjHoe9xNU/eeQBVmM3tnSQ0luXTyzEd5OLj4gD2dNjwE
FUCciZxZf0iIapOBN25wK0VA96KV5P9NQJ1zPindznLwlai3rnLdYKbh77+5qnAE
PoVOtIf6Q54JfDBiT7Pvhtw0TRP/W9sDGp6rePTklfyis0sdp3/FAIB/n9EbK1iL
M5r1MlIm/eCWmUKRJaZ2wklNqEqsEtepBZG4u4AQj39UgfOM8OQDaitxHmLh8BQX
ySUPbARknqosrISs5tdU/B0jZ5ppX67d2vtFM8vhYxopRtnPMHwWS+L0BQLo1Bli
/8D2lzZHZcabHHJuSawN7zKinymAApx6qrLxLey2pdYgPMEe05QKTlO0E8gyoJ52
7jk+YSyCC5NZP9men/7TL3tt2ddljCuXsAmDj9CJHfp7JchE+RJsdISEzk5MzeqT
we1T+AuW+8xmYdK4XL/XW/lQXk7P+paWW2FM7ZIVS8UIiOPkye3Ix9Dcwb+fjtil
Uiz5K7NCwazsnILNRppkaQwFXuJeqzN7AZCymk5FER8OJXI1OZ3z/t9jt25jea6Z
Hi+r6UjVh42kAfU4qksYFoHfCnhdPO8e8xAKxD4pEVdjxi+YUf/3X8JYvPAEeZs0
oG/UuEsMEwsXvp3LLFyWLA9FwmZjezvd7OWbbaCjpz96kWpQPOyM+L5p0s78j8vV
8/3OEtzAvpxx1OsvMbiVlDoXLxaAWrHuIkcCMeoqo/qGtv9NOhXe1x4xquVWEnUp
dAmNxLj/CjMWZtRfWgh8cgWHT9yocJD/PGvzCyqfxMJU/mexUVJn2SWqwCQ/3Czu
agWXhUqaVOqZiupX0HgTL27U/mghrwAfuA3EN0ow55JjVxQ/y65GNW9Nd0AQl9rx
5PyVGnVDio1bBnFBW3dOEdY+/jcAX2FdrgAkdPfAyDrmUp0Cvzr26XqP+XflBU4x
eCkr0sc7ChEBOggOExgx50ujlDufhiCaSWE+VpWfvdTkkv0ASzUBJNVdmbI8Odd0
upBXMENS/SVWIb8hNpEhR57n5hguQvHdCXiV+LK/Iz5fshqBoYlcAIB4qqpbBrfS
vwPwHnuNicBg9sI6dTigLnz+4/bRtehUnSF6HD4W2i0o6LhBWlzDSSokzfKJs6VM
OqVOm6OZN/pwGnolCLTpz+P5vbag1x3VYO6kz8E39zVUUDynJ9hATi0VwZMjgnQ4
JOMtPJPHY8iAK3zykCLPh4ZJuNssED6H7VGKJVD8OFnyGIB9wL/ybHd38SBqPius
sPTc7Owk7zhW0REJyHcZuv180an+P0PbbBqdRmQ3flNaKMAsEiFDBTmgozlmPxaZ
TNhpFgJAsQQgIrYSsrwzx+gWmV26UklgU5fyyUxqIAZkmzthGaWGMEHUgHSbFN10
VrIRmU2zs1fmyYldYgLEZWRjgGSt/Sxs7Uc6JyLJDaZ8OYvhG9tpQvNQ2k702xY0
x+irset1wj2hoORuEimcMF9cg1Rne89JbJZJwY1SYjWu/YwMcp0flH1watk5U0bq
i4bxd8PPdFNYILKO7tchgnZpfaPAxzsA/jCNwlA2lLG1LfdFhaia4nZzk4wHDL4L
/E7fGFGBCBUzSi/13qcQeZxSKl1KBSvpNHrIkwUSh6LtBSVSWRopvmtRrOHgDBgl
fx5s+SOXAw4jNiEanPEbIXKpMLQn4N7vyxHfLhjeoDegwMFvsEt0ZLWgQ/cQR/z/
OWO0GeHROa0rjxtS0APUnI/GQB8MRUOwqNq+DC+5cYd9L7gclaimCdAMSCJJd2No
b/1aOpzLWOzMM28blOta5gvcwbisCtStX5sQuiAY+wV1XKp/AJmIlFvLylXfPnZX
d2flXnv/WOcVt6KatS/jpiOOoMyIRsnMnu96u8IjBxBeOBCwpzwbvgufUe/SiPP8
fafN/2iu85JeUPI8SUJ97fLITfpxwoU3JRSBHxMY85fAyCu9BaRGm0Th610B65QX
nl9SNm+kNPrW+ZXrDCBupgw7OhFtcmi7O/xOlWhqWmzrqKZYRqHno+bqo6DP8cFb
MeYGy9nY4dIW9aDR7/iSNOUgGmaOxzUVbkO/Owiqyt7uwjoAYmdnphlEK51X38q/
jX3wLOtbs9JbzQRAdKbwPmZzVsqZkOwzmG5F1V33F9IH4e3p7fc0FM90WeSKBWIE
Zht7TOCYst0dX0atSdR5E4pdMjlXHv3b6MwLNWheD2pO5xwfFZ1vpTQUe5+ippEz
U441La+CK6K0pFfK8bKPQI3IwPRPF03741smAsghqfZDoNq7H9qaWx4jFm2VAMPV
sP5NpolzKfYbzcvgdVZjekq3W0FSyK3MMiI3KhSeE0qA/gTX2ymOawcEtjP86F6C
wjZILinKGxdwdBn4/8fsU8rRJeESDvvR0EO4gu5x76cDL3H1k/AxYY1lQBFrFLXT
PpFCUGDVRMcl8jHHvMoQ0tycP4dX4X+TILdHHL7fpLvkL3F4q8TYgqaOFzsgrSEY
sFVOlv9G642XkOO4vnsvEJc69bSmIvOs4BJBNtUNMIt1jqRZBBjKY/hVGZzf/xM0
Pc7XnqUjV/LlORbvGLyjgZ3FShimPBZui0Vn+pEaQQSjMYJJuAYl0UiS8P4Q3v7s
C50ttSzwfH1KNySoHSfUI6qLkjTqFM+Ga2hi52Sb4MsBBCU3NgVXnTC6VtgzJgJD
VL1eBjnqqYYAAtDAj4Bsm0dlTg6bo5k7tMHS5JXiHVm67an9ch8KEwv0cipxg1XQ
qCPqj9ZPcgZ/NE+5WQZHOR/iBt5hpLQtCyYlfkpxd6cV+BQwrf1nvmfIKlJn+onC
aU+AT9o65skYz2WrPC2FiOyzvo8nu2dGXrhpKCW3xIOu6b5ISBcaKjifw/XrLp35
JRoFrq4JdyvF9bhVWJ52wDf/GaqKnPVqan8tD110ToBv1gFn9tU0X0Lt7f9HLo4w
HyghPmT8mLzCWnFq1ADDxFHzcTxDzeS8+pN+kbmpoFfF8W1P0ES88R4CoPaoSW9y
ziEMmEKgKMFEBHCn6zxTG8JgLRUkiuZRdX/6gttU43UTRHX6J8u/1P4yCRh3uh4V
03niGg3WjDEIWOHOG7HPiuo6l5bz9YTP6sVoSDzOo4HZxoOWifAz9VTi+E5hmb8M
FSXXCdrC/Ux2gsGxgfzav6SyiZDzy68UiZ9b6WTHN8aC4kpIU1mL+S1eT5EmUQuR
ZcRsuvC6KEMFtoyTamlY3G0c4ZuS0b7SZVe1/NozLmep0EtPrNjWmY8ysdFPrrcU
Mt6sEqS5zolk3/dRaZHEeZSsBKrxU0lg+VhAwJa89bSyhdFxwAbtVZQOsl2zNreb
fTKfsfxIi4n+xTLI/SArArAksobNq7X9N6p4lavZODL3MB6zvvMsi7hqgivkASXZ
nobRHFMFGcNCc3ng4oRZMpe31xddZNFGZrzftBP2yQwf/EzAFUzSDIRfyDgAAN1h
xIaYAVoaD5Lq5sFPF0TKFC4lerQ8S8C/YTQ39ne3mjZ2Wuad94XASTfvd7xc04dG
3zQxtlqgYCnWPAtd6CEttAiYT+2h1GjBySQ4UPf5856ZFHwFzYxbVyIXoS/icMHf
7iwvS3/6fRVH2QxbKouxGn1ZHI6BL/sgP3H/vHMsKChjeg60XMbMLs2QYVJcdjcI
S5A6razRfUfFUyzn5nPPgxVemmV+yPWPZ+Y2NyfgmJxRrKQNGGW5nhEzooTe+obI
qtdD43Iq2jGB39YN3koocEOFf50t3yfM4f0BejKIrs0vpxX6kRLonv19qAL90lGU
n91CQyVPMLJaKtiXJohVJHW6l9SE7wD8xuMCA8134M3tiHiym7NwUE/1uvX3vx4l
ybjvvqCusN1ZQSG6/PT1JCTWxNZRxmA7u6Hbw/yoQhInuASwBTJXFq68Tvfaijkc
ZLTDtGKvaC1Di2jtMmiyUTbh3EIGCPPbw7JNWQVrkzsEthCY2MvrCsrDsjijQjOZ
je+iLdAHGZEpePVj0H9MV/qGgNeQO0JwgOqhpiojokTpZ2XIQ/2eJzlDXjbG6+w5
GnmDy229P6maLRHhqPo1zGybGg7LEgDIOs3XRt02LTRcMGzpFKcn196bihwlzI/x
sf0A9PA7aozi2GtYRTHsVCJUIss2GLV2hNqMDONiLKdUUZ53C9nVOwy7/VBy5zJn
zV380/3KAg+99qkwczMNjiCMbqfjtwxegU4Uh+YNfnlDGzIlP0ejrsKOeJ5NiMqw
o1dUd8aDsTxORcVQMbCLtEk/NgBTXaDpQLYOwcLNdF1zf6LL3sIH/yAt7LgTsWds
AEeiCmVU/B45SAjOJNRQ8lTqOFQ0x9/Xa/5bobeUkrvlWuMnK/CZNB9fQ39eZR0z
8MMCGPWB1grRzAu2ZUMH3wv20r3XdtQno9osd4sIM+x+ooaIb8kvC2DPiuU3ezsp
DZpvDSr9pxEvAQcggIjRk3fqlSa0+g9OhOJ4jPjckaSUZpD9soHWMy8l+/7VQvVB
3OUw1eFAs8nUntEXhB+QBKK5MSPF0lOMc50ho7Rj66LckaXNjWw04McWanH+bewi
KXIQ1VMwILsw5LLKv7iVBmq09/HL/bw6R4GwokIeRZPRLtS7lK3vT+MgGAtGt79Z
0rvLcIaYveO9du8PpkzJNylS4pxz1Va78wuFiOsSyMJk1uYoX+h7EmNMHOtHmb/5
kFVIo/ECFuHgTlnMuQaAe6mXOjXdxi4oZhLplfh7Y2efcQkDJ7U9Np83yrDFWFio
OyaE7iRL9TO7cNBWlhfB0Wr5dHK1w90ulb+KKuy/6+UcX8JeuqRdIHk5ZF65WSk+
YXcN34dw/BRH8sYOjLYzatu0vm072E/OXs87o487LNdCDKWeCNzwMY8CpSoAiRMm
i7fJqrpogZxGN/WWLIx1SwaNJiFsupZt/eGPRYq65eyPlV8bgNGP4G1gwlVzfGQC
f/X8SclpngD+wTIQb1n9oteTSz9d13ioNvxvVDDYwnhQOClVmFAwlu/ttEKEY5Qd
lAYt2tiB1efIIJzimWel9TALIfYlJDl+Tlzo7KoCOtSgg5Ji2yq/jOde088rCXKo
KhOvq6uc6oCRSFJwfUulaKG3FTQJAen4gkIoLhYe/sCzorXj5ZMvpF31+aMp9/pg
9WMz3Sly8UzSOlBR5KCXvEIBcNer6Lij2vtI2+ieqXN1xp3Xs/DM6hKI+Xrrs+fY
OoEG1EwEVyAcJ6/GqLt4u2bRaYoCA4CBwbXnGOgb8X1epMMWlh2pFm63nJWIcNf0
tfejLl3Un0RzLu/K28veXhjEE+uppngSE7Z5zDHcqEuK2PZG7nJi5GY/ibK/eTnk
rHnPMbmLrLYoihseiYhYEfjN7GqaUaX50Q8RiXRrg5C3f+i31Q8wHCdBOS721MmS
BJj7J8Oq+ea68qPsK7F1Ba0NDEYV3jblzxRcVDGwCw/QcqJFQYo2V5KrdFYb7Vqw
O7V85Fc953GvvlBU46E6EYVFHreLHptDJVJIm3kM8HD8mj9NXhhMi2LCkERa0+i6
gMz8RzSbPsNiFD8OTGXNFCAzia56o0/fnjXNDnS3u624CxpNsQ/L8B2d7fx8DRal
4Ckue1ptnBWGMjARiuz2WaeH6KQG40vCJZ8GZVmNXVsBhuDfqtJR4Te6ady6vIU3
dm33doOVbdHB9fLf4T1ELckBnMsgod47QfjqY1pmbZR4r/q/EbVQPk9M5Tic5vWB
arRy3hrxLHhWs3R2TQqWkUkb2IgXoAbRQROwBvlCFIqr2M+hHZX/IFevVrHVZmoh
bZJoWUSsLgm1l4uIHqlyE63BLhmX/W9ed3jGRiyT6xvQbCbP8JXZsRR7kZeu44K9
uoqj+ljumajcRcE5eId89eiyhXipdfE6ToJYWIZKSf8tJW1zmeObEkYwz5A6aaCB
vDVjrJIg/xG0WiRm5HPwWeK+vVwME2o3C0hAdsLAYgis3mufRLwc0DugBk412OPR
/xbiZ/UQFtOa+/ovOoQzJnI5hrCz2p2g4IHDEUpytX+3RAbgf4OvivR3Xa3LB+R9
sA1MYoKKd4PiCHhcrpCeSgWcL8CcWzdiompS0rcSXO73SqpDP3j+amDdHj+F+vpC
h0K6TVhCksejDsbfSXIW8oVXkFok9B0SWRXRsccbQu8deDS6g3LeUxh96Vut985k
Zu0WRtcQ4xI6JIYtdoyYL+hPfbfo8ZeaWKhkQ+GjADzp7rv+0BZYWygt/ZKY4aeX
AJ/ftaBtboijnhHhKZpaK2PyEScjTkHdlt5nZZGiB+v61JD0mBrwUAIGYVIU/pvQ
XBIk/ZewHIXCmgIBCFeK1r+4KW+aQNjaZ0GBilyuS/ZmHkIHtqp9ek+Hx3nsOEkF
wpzCkGIETBdcqqG7MbTB/YL1Qfgks4T/a0M670lcuOZrUtpq3sB/DWoF9nTkw21q
WDROx+sGyNLlISeGzm/Cw8UnC9SGjf58zxuddvqkS1vvX8pgqUQaqoa+wYj6+by6
Ir74c/ltZbKSakKbTv4aPqWafC//678Q2QPL5AqMUjo2vyawfj8pMPSAnnfTD845
d2UHm1nCiwc6FmiKuj3AfTAFHerQn6eALAkfPMGTVR//t4xbGrXbwWpM8+59LOjP
kjm0FpZixcWKflSUAWL/QiLhEXITEiizmBmgycDChFL4QCq8gfoezwWZOeGtiMA5
KGU95Ggk9wDZYmkshRsR72f5NH1TeirlvIj9XG2hfkmMkJ0n9jgamEB7SId3+uKv
wGTqycg4zXWYNwV97q8rn3FLctEdbnPMtmFNIGCYh2seDvyPQzJuvexwQXENj7JD
1COH1b6n+RXdJIVUGBLu/OrWR2zOEW/6U9Na4BMqwXqTGKeYqIsylVuE15hweIaL
L8lQ74vlvtYbtoywVFg0VDwvIL3Yb13DI25I1BZMtcRvKBHJb75ioThcF5SsSu3R
GK/oR9XluOdGrLs6hD0MAZYDJl+uWQLSYcwOo9JVsMGULrUwWViERQTSyaRf3I2K
44LT7J9mJ/mzQsGeR04Lmj3GNSkuFsx9a4csyZpMZI4+lpW7cLziDcfG8I73QYWk
p4rblTyAMp2QKFS3G0Ul/dNnG42kC2nacTa7F0Ow1o5YSocwcKOHys5ZU1m0MvS0
Qhv+yBV84QChTyfNM/M7y0Y3JIieNRawSwN3RGXvQ019kY6woY+5UEeu1Z3RFMqc
KtB4V5kEJN8Cg+1IFQvblO9UAUYzDjTcPq9KAR1oml8RIRajuKtKCK29khNAUMkK
KPz19jDKNSm0ilrgQv0NZHVciHcKkNR0ezwcHASR0+UE2N7g/59gDzmsUFwXHuY0
vN+Yoc3GQz56PnvwDvw7zsUIYuYYle5+oGPp9rLOoKloJffW/fja8ylWrwP7V7Jx
2em7ymjXXaKRk7NRSH93hjSFE51XXmtaYRILZnx0dT2ETRNwGgtHxai2/u9+a4aw
LFK7zACCmLH4GCODNwWrO7Qt3FgqhTVCvgSr+iBEErsXMib0tcvHI7PMkhElPLz5
6zBfzxksImlti0qfESba/YME3sS06kavatZLQi0hjlfVtkReYFDnwlAE/3J7IeSG
kKPdW+cVlQsktqMSfHw1qMJKJRKs9ERt7D3tXNwldrUQ+gbbUx6HQyE0grNPdhtx
X8DhlCuvxAjaY31PzF2nKjTPNf02nn+XeYT4qUB+spRWPEv3lx8mXTpdLJEGNi4n
5+yJeuV0+yY09y/tlM5QYwGBAsl3dIRK8s4R8dkH2eYhiKvCtwMiI3oIv3ubx3y/
1aKDDzOzHNr5Lvwf1pgB7Gs/YBWZo3WRNjU2GvrOuaoO9SF2tU8JH5sAV0AK9M9i
iMgpHTlZiw7sg3DyEpdIk39GXORQp61YsGzX8s7Z6YRACfSJdhbb6mlcVeS1FjtX
5bWB/rMlSrvILaQNQY6IgODesmn8fmRp5Y917M9KRX/dcv45EJ5bkhavuMLyxA5v
JMjbSTl+SjpKGBX3GEWfPpxlzYyCKPb5NdpPxX3YRTY4/M1q8rcHTCFKId2AZb5D
C5FWXWBA5OcJZoZrPPmQhUAcnoIpOXo2OKg/R8deADr/oLHR/cPuamFw5Ht0UT6l
4gSMs5ccc92rsv+vl8KntyZwAVn30arEM1DeK4i8wy4LY+ri0f9xLku0X056K4/5
8WdsHhEULU/nJA2Ddz8jQlVC1KqiBmP3FRdER+BZgOqVEWqwPPbFQHLXO738b8Ob
IduP9qpYApBlN5H2e284Ph3bxBpyY8o4mL42ZzKipUkgso9kRHet0mFw5YP79eYT
5Hp0WZ0s8FSGIHgqyWAn/hLJ3vsUBH7y9u+mbwEu2QKryGcTspvHKXOHTCJhbPVL
jVV/tvX7e6DGifiARTBOtjYW0+XSWA+dDF3XRvMN6YbPVJEMPiHRzwijUiClGZVd
rcXZT4Kw3BkFTNgMu3QtgiTq6MRNh3nI+5Z8RMvmtkL2bY238gWfdzL+y2nctfqK
xC+qfLT05Q7qMusA8UDrapAGKycZacVtpe20DPdBgdD7fzGBkj2iC+s9eDmXHUGW
yMy/h8tFdz9A8XpxWP/Qh+KfWppfZfe7K0v/mRU09dA+vEk13MZGPeAvEK+2WByC
/D8iUjrqOUsUXZ4OUOixV3t3BhsiJv2qmJclNqGUzKeNwg8Ahcn2sKZwoKTOO0ok
w1LZmhs5c3Zh6v0LL+Pahb7nLDw5wACTfGtehOVxM9NsQrH8aDmWCYeY4tx0aQWY
ynqNmpaskEi6UAs7DE6m9DzxpjauiGhI+9M94cEVy9I6lmVdD0qw6IcGMFf2N5ai
z7+o0M+jCdKphEKhoXcAl+0/R5J7CYZp6pCDobRgtOFAOLHzNZbmiWbPG5UgeNKf
2EubeNHtujxvz2fRPESrSfeo6z+BhFjsQWQjVsvJDLhq1D6ekNk/LTk/DqwSYj9W
6ZyifrSar+MXDQrXQiA2rbyKIS4ab+ec3Yqd9OPeO4uZ8Zjfv/lXRIR+HUlJbV3s
do3W5rdNHvGj3vH610hd3gJ6CqZoCApO5TQKlrzeptWsK1NVYs0As/qRukGG/ITr
v7nO/lry8tOS+RXELJAa4dbM74DKo1GSyiBsNVJdSjlHhF1o52yxfQcfzQxf6kaa
2Ydpr/I1hsuEfbtcM/pqkEpJPXYNtXg0WbsyTBtRmcar573t6SgfHfqocg+lXKa1
IiRv1iaSkSTdV606WXhRrPQNlQtmtI+BkziwueVjcnq0Zc+XbuEppDn7mzJU5ZCK
SFmr4JVgFG8GdOK+ACXjzbR+wp3/RRs3n/C3nkH7XM8HlDBnmeHVpf/YYEeMi98r
zLnQVDsTWbl6Fn7bulJ39IbwhLNmdFAtOyId3EX4fTRjK060bmM+H/8I+UWUXRB4
GOTmPefKQU0EL394Xl9DEKYsvx8L2jdyVV2n7wzgpL+VuuKuS/CGrHis6LpAxO/i
DiJfWfQtmvjmOjrGX1wex/Q0tWSgpK6BG5DN4d2cX4yYBB3uaSWi3f8kPSTJfV4p
PtlsV2IxieDbCQum94TQIU4R1NOZaEUewCAYNbpdp6gAxfslG3izXVwanSW3WVWh
u8T+NWxEti0yaQpQ9xTW02Nqk57LPFqyJtiBb/ndT8DXPXvetdBLQEj+4Q3Z6Xok
7mGHZfKHpfkxn8iH2GvvsU5fsONnk1I1+Fd6zrBmfIT3duHqaFsc1VuugAA8SH4C
eNhjD9kys1sei9yj++MkOhidRH4SULL5Mf3CcyKCHmUyHKdxi/tNC+2ue9Po4+bF
rDGT8zQqCd+kUmpYVvllYoi+BfOM9Yk0AWYFVq7aOu9HC7L6w9FoC7vZlPPnrQxB
vlMNszRJkkPb2scXuXUQ2e0K+Fao1FIFFG2BP5A31pHXQ1A0NwBVvAPFd8tjtN4m
27pL875lPiUpzwzU2j/g+tVznv2EBGds5TQOW+V+fZdIApnuxUTECxbCEYISQfyl
DtnZE4qqTJ11xZ+sEHdlnojicDTKE7YRMxQCkvOKLt7SWyzjcKY+AV3Y7FpoPSvE
pqQmg+HC5PFGQ6nYqcpQKaeV87jW3dahqwnbF17bWy3fF6QYcCbGjYfapEpMx2DJ
WEN3kzJBw9i21odObOWxQylyUXXUn9zo3JDwxnb0wZqOrq4eCE9FdF3Z8uyEf4pl
OfJxhnfHrXr0YgmlRKR+p6r/jxLekbbf4Z33w3DVdQrQ9ZuwOlt1RCJKS/MHvhIe
/YHdSibST9og3L1XrKI7EGEVbDtk0apd6lpco8N9nWpSzI8nSMMqZ16VfOcOaM5S
29D1xuRc1RVrWr0Ax+sCFGOLOSpVgeUE6pKBWelo9IU7AKT/TwbJv9tdAHUt9Uh6
k261+c8e3JThnC+mtcFt35mdFfycVzTAjRnEK3eXmyCLvCq9MhPO3WhCXRRmSnD2
NeMj8OwfaU6/S+mJe8U9S45goIfLcjk2AvT2zqWliNwKWFKlP3L2H4eefGal4Wxh
olKGwFbu+ZjEHjU6LIWGE22Au+MzCQWC2AY7xhymSEvuYHA8JLm9yZbDTiRypxEh
tT7qQVSZlRQ/u/cr8MKylPf8ybjX6QgRs411iL60hfJTT7QAeFjOE18cvkwN+Vqc
+sNOgWzdrUgGETucblO+yAhglDJj7cZnQd/tuu8MbwKYQvhRDN4dCCU/jbcysGsx
O0SsTOvWd2PXMF3xbh3GC2qYlXVYupjOlw+Kx54VOgKi2WbF+yZWWR+cSWbBLrfI
UNFCHgDXYsSZfoXWN2jRN2oxwF/6utblnwSVndMlankzP9ZTUOvWUg6U9Xy60aHb
eZN4QwxgS/bm+KO6NY+EdRf0TrwdJVnYdvVEn/5KU0cod9ijKdvB1m6Bb0MPmtad
0aINE3/2qUTZxIuGzZiNrjrOq2pk72ju/xUBZK9g73Ip3BPAP9OKRvU1sreBIiB4
dbZbAcm3+tz9nY6zwyhhCVUmnysAqKMhGnciSODdGm8LjfYkTjHoS6+PwGDAyXND
oLHdN12U8Z0mz2ZZTcOQvLY9h26LQQFon94PcQ63cmCqZjevc+4FswlgGYhkujV2
5ZXA/xmkRJsl3/9lg+jdQ6qHv9K3pONvn2NmtOuZn65y+uB7q9MpVBrY3oI4Gg2E
SXPGYr+qZz3Rr+IBtbvY2WavfQ2Xd9mZBb13VbgP8aGYfykcRFAG878jxRfrRML+
H/B6Vv8K4pdgzitqIdg2sSMUY7Vp6EzEbrwgK7zq4LDptjnFITF36+KgRr3zpt7d
/lLvLWJvVnxfPcWPVQusFAhS1HjV0jBEwdvmRxGOBn+ptJBCgvsi4WKO/+ZtYcgb
VkzqyGrPhjB4gugmnjhfOj7BYJVG6PwcEYnf8JRIvT+dGFRhT0b8dMal/Gkxa1r5
d8I1lpA5XlM4PkdfNYhpVMOs3gvqJk4+Bg7cWhaw86X8xT23KQH8G6wUajB3R11p
kUbCGGRUQ94kLsT+yrSWbAeperC1Jnukt1USTqYVD/i/QxACG8CY2L8Ror+rxsZ+
quStMhylJBEYlvhcgWjlTwXJqkmj6Z0G8Lv1F/diky3C8E3zbY51xoWv/raoOzdi
JC3STIhV7UiVspEeLm1KBYIS9O3wsa5TTlxJyXblmLCIFLN2Au33xK+zVZz6nJ3a
vpKjRLJWQYYu8xxLlnEvLJYVOMeMZzrN33XHgRR0R4rFQ+jKbzkn07y+ISgbP0nI
TwqRlAhVioxptz/kZE15/XxjkqB61UtYNhUqbZOh6p0VHuFmEO8DwwhHqZKfRFkc
p7DOQX2Lo+r9UOVV3oGK3XaBTvZid6jg6el/hKaeyoVg3uZepTT2Th6QncAk623H
3hhQYg3hqPUDKk9ph1igI4h2ps5YKu7FcGCZNg1QLn461QoWGj3KvTSNCCSbhz7o
QnloC/kZ8Jd7egX3aEakJzu302s1qcMRBTqrHm2hwEVbx2xnbkbfZqallRuvOIjO
zE2E/DkQScYLwKRDfVGqQnOrbSLcqCJRdLBwfaJiI8fkhynDeRWKJQKLYUQ5c/JN
1ebzhT2xU7ZfYsWJ3ji0AE+gKBupA2zLY4QHQ9zFuiHTvjC0CPhJQeVZyMQ7ea8p
Oznk3RtbQiNceG3ey6EL9PfyazXP87tUgjY2XL6KCZC4UBq+0TR1XrU2bqujyqJ/
cdxm/n4Yc+gJpNjh0NOUItO1y+J/qBAPD0Efr5eAqNuL3Of3in2GI7DsUQwb5KJv
h8aqBAbIXZ0gKmZjcp8rn/9tDr8Wa8IWIMvCiaGbi1ru8vLbzKZmNyEr3CUSzBHt
RmZudhn3JeZCNcsXM8Wb0lLw+E/QdsHDW/ApI4NdN1V7OQZa+i1Q8Ur6P1B1DbYu
5X3+GVYsQSLS24U8nUfK7djoEHZ/Hoc0HdMhKiCYeeX6SsMpKmWmvXL3EwpRbs2E
Kkr6QzXnTbD7FQqkuD37uDRggZNnXa1SP1mObJ55/UpIicdeD8l19Aq7OHUA5ft/
EsHlzVPd5PTB7LDDBZkshXFhjPRvjxyBD9xWOJtj5/P3HpfFJp0B+60FMssRWMKs
gWnY99B19Fm6DxJxS6tyEW1vru6cE5IF7TKX5GatBne2GTM0689Jx5F34V9ptp5D
zHtAxABsFiH8BUIu7iLCvtcE1GEFrB2Txw3sPvygkWF96ARHcTl3DrnrAY8CMTAZ
j5Fd8FjNpTnGmCofIBx0wy2ylIbysDHtskqb/OA3OTczGys1OS1ue5N+JrCdlGbe
7GvgSrqPZzdx20zmf5ue033mOLYqPhDQ77yXAD9s9/urvPHL5pLU9908W0w3FvKW
0Nmx361DTSmEfxRB8u+zqKH/na6a06iUwFIpTPA34+E2f8mDWICncNOIMbGLz4oG
oaC6MW9j4lhG+4SpdaH+ltrcana3Ae5IYaPYhT/pd/xAL09LklboYkY1w+FnlhhW
rAJO2qSayUNj92zieM0AT4sGFQw3wu0u7t3HM0gdEVw6lNf0jTyJr/xpMj/s+n0m
ALDdhCh9/0SvlKCrdQsql1TS8LD41Vz02nVxSBykTfU8v3avoMuEdJfjBdF15j34
7lvdymnXb59mht7xh3/+kadR8FMzVKWAz2Qd3rwvOdYDQXW5kkSo87RpACSZS1Qu
stDIpUNTNmnafAbzysUS+8OVOCG4VC+KGy38OeiH37zD/CzXDf2mn9LEpOFahvXR
t93DbVcpczD0POACGgyC78AWPb7oAVnLWrrPDjlIfnovH/pPXOE764Jie64R/Jri
AMYyHz8SlLstn7Ch5ULcK7WpMTFKH95/vlvGuOiG6b4H+4K0Yua9PuQmUxewq+eN
fwvGG7ZjYGPtD6tmCzRUzvz2zgpya2QEtSqymjJ2A51cmrWxCSdCxTaN0X7C7Xbm
w76rMlm6o9sAm2tvXLjeMk4dlPi0aoaJ7bSLSqnbHnsU1Q2mf1VVM0XEg/etLRsR
GMucyGUX10B6Dv7jH9j7RSSHY1wE14l5D2saB5XESLIp9qkG22p965N76XsTi65b
un59OtFExsDTYpKH9Oy7o/RYjplg99JIS7j6yW6eRuDAAnui2dZNXOAE5VFinJdH
l8RWEOUXW50odZjgmsD1r7/3Bq/fiCC8yBhEZWDGPk4RnB93FJsGXftmJ7pGS9vn
rSdiCcqIydciLtrjgxjlVt2K9C4xxPwTVdFfFhDQElbtjmOsrK78Uq7/vVQocsuQ
xg2jR3pmYyQz5y23EGbkDhXH8j/aoObYScbtr8q/2uMIdCszTwGWSLwq1oufOzpS
UgAvc2FxrKxAVLKn4hlpMIPZlkaVQmIRwgJs6MbOUFdL1LVo6pFBrojTZoofkM8v
zOXkR/YZBMZBGIKStWszluYks3+lLG9KHmrl9cXRTnpE+2XMWxrAE0qyZgOiCkut
CjrmJVTqeEfX2Y+8oy5czeLuUZlRqGpgTmJC135RqY+Zjae7evmwVsv41NO7OXCU
FwMk1kK/m8DwSucHc5BUVQTwe/18n9leg9JWQ5qJlbRrHZlLwKdecSWhsBzt2bb8
8TnlRY6LxwQn3BkHyWY2/9opkyPFC7rwCDv5c2gyiElvDixHEZ48ZKChDSCyAkvX
ayF7PPRPyPnY/u4R0WV+n4ki5bkmwmgmICkKkH5NotOfQbtXDTd9q2Rm3CeRbsyO
gvDkE3Ilv/KGN/r3m4ppAHbRSsrvEfNLfBS//Z7IpnJRe6hO5K1YRFTSgFiMVTPY
E9S1g41v2YAoagggotEgzNcVWPtEaYfdkSVECGN1YnClS429K2Jjqlcbe9hB6Ft6
wkHm6Af73n9vwE//A6QXYT/0ceA5FjE+gujGD3kEXfki/1vVmQplcSaZBi06TGff
Ps4Udkq9RbAPcscBN5lR0sUoVRl/sS17CscwgHicGBI+/L8ydHPu7fAHuJS2/I2A
NKrkwaIMBE+1Y6Mk0Ra4lvJGYbGApA3lIiMBi23aUpo+/19+I0Kbs1M/pGr+uzGz
pvlZarYVolpszQARE6KioMrFZoGI7xYRryKRDg24wi7Mm0CCA+Fd4RC3PhGesqO1
bXv9po9mVvur2+c8f3LuAeBF0MEDXv4Mc4AdIHqTfL2y1/dxrHiXOihp6V1bfl8e
EUGXTzWIJDF7I8YyaIN0Shctho0mgACwGVwlU3jqLdpA8xxI/MacvFsJ39gY3olr
wX1DSIo6WcJRWYTZTcBlgqs/M58wDMeX0vZqoi1nixqX8xJFwRXK/yGlXbow2Wdd
/uikMF8Qs9nVOQ00MlNkhNOCd5nCJjJeSKqDsYPkCGW6etXOAC+gzu74cExxVK+I
/KDAPfZY8u+UaG/XacrMkdVEgAHdfeD2gOM1BawudU492aZcQBnylcpd65Ejf367
4xYNvcCA/4J8F51dKUaoXWPJKvadIhA403d2CfV7ZaUdcScofH/AxAY0Dzut0b0Q
PmL/z2MtuOzmFO9aFT+teMdilyGqoa2/9TwkyCwJxUDUsXw6eGytsFsP1KoktIrX
L96Dr6ZeAeGmS9h+KXWdWOzxzdmF8Ge+eNVuqp6ROgJK9KBgzMuw8g+PWl7Npvq/
WQW/1Wweo0omwLg84uAL13RBjHRpzJkVCrB9HRXfjClx2ZIpgXEvQpNEMPZTuPdu
VYqW2bMJXphMyJfYRtkfLEVVJHezGJcg9bs/jKkstSufHYV0P+NJFAyOV23C1b4K
3oudResIbe3KuSfdfVoetcm9Pqckkud6PU4VZRZ4E1HPx41mYDUXF24+r5RWAEcf
iV9CAJtSaY/JW2qnltsfC2f5dGmpGRDVtYNZb7Ltx77BgD6dbBj6KDtliQaqruKk
ZfTK9MzYrEiYxelqv9Hjl/xB6ZsoomN9nvJSrirRuS/CZy6GmaEsqIbmqIdXCDQC
6Jihc7yETVAl5DxjWHQHUUFtAM5/lOhBOfKTFXgAJEaUG3bw1ANvtIp1qb3cN+t+
lLPEvxlP11MVs6YR8+sbXGraiZN30LWGqt+yefXxKZHoe8+f6hS8EFGGZZg2B6i/
kkOyXwlTocyzehtKwj4Zq0D/uyimnEyBcZqKKTiFLpdMr1Zvh7sAZttFH5S0UMpn
1NdmVzhuSIRcZ341X/+wQ+uQ8X0eUz6v7eWWgdKCbYlR6947laeq3t29JeSchvk/
uRNhdu/N7TJuKmsl0/0pKt+f/HHh93v5IEQRKMBasvw2JF6Xb0iB32eeo73MnjHv
+euG+uNVPYyMxj1ZVvpjTRshBT+6/NqjFA9avZSdLJDotozuxHPE3lbtczu9ai99
KcRrmE9HAylHtzkCvVTNZZifnl+/fd/UTjgH3W1dptsLwWmBGWPa7LtZduW0mMlG
PLMAbW6mM3b4mSzWY0+zJKPOB6541SpVuf14qL0ARpf/qyKy2gKFargrjXwzqUx3
52AsOp+CBqN6wqnWtyrf8L04hdNXKzo8R6QkPwAsUtl88iRm8lBYogzAQRTgGwvk
kMKrIMLHwP2NkfQUxeoJsr1FVgVYNJdFvNfDA7pPVLYm2TlWRwAWUt0Bk1yQ+UBL
//l54U3xM858kmqN+NqIEFTdDW0YdhvRGdNIJVoWEgBL5DiI+Nj8RfWunPvvAC/8
RZHbCO7vAMWn9fInu6g/DtT17mNYtYJNj59BUIVHqNeuONiufIBoKKHLFDzIdrr/
LgNaPbJYAsFjSNK2I1uk1Nev+c5PJinp7RFxzmzuwVNLCwWZH46v/dhIWOf9QFz3
L3ivIoAxqHUwAJWevpL3YE7gB0TpDRP5zCW8IY0h+8wIii6mq9IGG/MYsa3kz/Ip
6bQWBetswUg+5DbXhifMD94HuQx10WYeiKqG8PtE6SbNqpx5JDV/7zqIi8tP6D87
0PJgGgNlgxvUwpHd1wCDAerfClcr3muaZCz/RRfb2AaWNw89GyIMgucGYupsmoPF
qsH6+PqPBkHhxXlJIYux1i06Q6+U3i5qJFCmy6R+RMZc7cSJ6t5rKA/sUAKG1ZRW
awLkhuSle58F2pgd6525hS8JmJMxQozt4zfOhl9i2qiCk1Asnq0zqMtoBMq4KsVy
7uOsuljrh5m64HyEDVSkcttKViCKTN77YAh+bsVtiE6CmX8xEeyi/x8N/7FQg9bY
UTELMx5LlvuMzA2Ec9S0LcXtFdNKf8eX7QS6A7PvvzXSqQLcPK8c+3JZPH31MtLK
FoAwplCci6/lGtYtfahy27IWdSlH3UMrX7vX6ugHe9Xs7pJ+BMQlsYGlBFjCj0Q5
/NkOJZqXDqYRA5Xi7uQileBOShWg87rIUHS/AOATSUm1Jh8RvAYSqk8pzWCuUuyK
2pFPN2AJMVAF6njx9x3HO6J99DDlEeNkdKZTrDP2hA5ZMeT+boM16RFA+d1layKy
ToXrLaIq7ccRAP2MF+zVoXWqUYBcPIXUr90ypB/QkqMeksC574cz98+t7eg8fWb+
f3E9jCj/ICrrVKrAaWpO0EVp4TRPpm+vrbkTPAGQp4eDELZk2TO7PdZwF4cZ4ESY
73+tovkkftHwFmOiDKWmgkaTDk9s23yIi8fAR4/sGuJGfx6+XWrXSmKG38tywfI5
UHnKhWjAVFiEVvpL35w5dWKVm30f81KkDzORJyySdv/RSDmV0l9w4sRBlErWQQ53
8oubjzI/j2V8R1zyo7BKoXES3xqI0dEsyB3sQSQ27LyblvwxZKhVCYiLwTvGMvEQ
QUkYmHp9om32SVeIoLunUBJCw6oNYbgWSkL3/x8HoV9hOYtyvIKhenYup2Fr0oJD
I14PINkmpIeweJSMzkFhLV1Jc5vJSI78YxnbiQND8MQjcxrEmiAninq1z8ndpvWf
s5FsjC+46vHPcpPUqAydT1XLnLIs9oArxUcsORc0rtzHIVeC6GM//2s3gJuUbA29
Zgrs9pWirg1DOP3YT3NgrB/7cLp8PEYN2WECEyfpsduzVRfB+6gO5RvSGm0Je+EP
yyoS3H8l89m8LzJE6P7FFliKkpX0onVXw36C0slbJf7fNIFtnMQ7F5C8xenWk8/C
w8n4smQBvYMXUH77e9FH4gA7Oea161C0jjvUp48MDHVdaeHahRtqRJp+LX33tktW
5TctJ1gwpHfvPQ+jsK52/5UI7v7NEDk83ord+GhqFNPV/XXAm4cfQ3B01On19mmB
H0X4j0LthJFEBnaX2JjY90rUYN43KBzbseYLNyAo07uSR2YxH3vZOt7BJYDH8cao
kJIcnT0G2kjLt4WQiO61oUPJ50U8fUNnJAnK8y9chhibfHpSFgaMC1CtsugRxvdL
1eTDGzJhGTBEY3RfGP3vQ2RAYGUI4iS+tJdwCssJk+6ov5fzuhDIT5Wwl/ftDsNg
l1mVdDu6wQzsAiAP0kFhnshSJJNIxCAMOkhKnOLD6GVB8j9bIANYspd5emRt7oMo
UET5kLZ8LCQ7oy9cONl1c1bUs4vtpYM3da5AFxm9Rm10wa+8PGPQcZKdQjQJ6tRI
SPQOam+htfKpcWiLPEM97pE5Dz3kg0+vbaYeQmJtU1jlP5tI7emQdx9m7H8Xn92E
glTZH1WdghKDA8jYGZBrTBZrvSf9hiUpP4eVBh9NftZ9lttoTGYTR0SsLi81L3YG
4EVv6DiTEH7Ek014SmFHlhE6e2vdkQ2H5otZvW+prxeD/PWuSMdsNtkevMrdtSX2
g91mDpFHm+/uU8/qYySdZx6RZqcDNTEzQbkzhjyRsVovjzSZ3zWSO2jyu1HN9Tzx
8Gyh22HdU5BE9R6RIIx4/MogriTK5ioNidEhFCQE/+qhLGkXhDl8wSMoPuM6rubu
LW5VqnBxuRHLwGvCEFFTFHFdxtqwy1QD2RFe5yAsvENDvvhubvgpytT6gV6y188L
wAaUsWKomksh70XHE2VKmn9xyCFEjSa8VYSjnTIMnesbrE41LnSf0xqJL3h3m3Jf
vyTJYwZPncN4H/kbR4yl9ezpRBOu6xL+AdlGubZnQGssRmzuMr5iEot8byHYfziC
IpUrqbUiXeo5LyBZAuOM4ksVu6kUFns8Q4FWp5I5mgparMgoic7I4CJoT1ee5okU
3Kb7zPh9drIh8Wcl+58tv+evwGyGXfl3xgvVbvZkrFOtqkY3khtPptAvbW6WuwGj
ANGOuaT2B6Kx0lGuO5AgLQutTI76KZ1w703xVs84xnJwMljdg7/dCjE6LsKo26+1
YI5O0bicq6DsxaJvmxXrEyFjipr4CMdkrKSJtXeKK28Idy+9Myln2IBTtIK7CXfW
s3h8hQHo6tTPnsu/bH+9/axwvK9PMI3mWqGaIObOGagRh6sOL3DCLIP5OLm+Lroz
A01fc91SEofI4m/Owo1QLeOgKEOsbzSYXLe2GKVw3HDrMNN2avCod/YaS8fiZ5eZ
1HNk+xXJ35hOeNOzlTUmrSlVqzEGUNYN3uU6w+JE/WHRucoq9iN9Sxi22VG/R6oR
uatifrQmI4+qHFxJ4+v/DB1nPn0Tf7dsxA/PiI33x28CrlQezHOgCdmyWSBLuUCb
JTGkXdK0y2HCMCKFtJf9Qn1Jf/n0WTc/lzrkQX0U2dCJ2wsZnDlWcBItIWDmOEPK
+Jxa4Ql+2HULwk0NytOFNo8B/3iYPbHtv6feb71if9hNStkGCZnfAcK1C8spG5GV
sFYjnruMM4qVof8aRfoh6Gf1l5QHYYVpMaFA20VZKNuEtODTRv6I72uP0C3O5reK
YAnIrYPbQjssn8cU6YocXBjevDnHgZknMmLhURkxz1TiuHe7sJm3N61J9IKgBCov
J03h4NN3aP+Zagw8ma6A51PNgQbvlItFwBoGHOi0nxGDVR7NphTerRUoEV6XEGT2
2uCWtzckOT3CK4GJhxMU3snhlk4H5IZCA4UJiPMU17jq2HPDsrX1jIBiHXdl1f5a
FzNxlaHwU+Qk6Wmtg3qSXYReC4gzr6zokBCzftQr5oCgOEok0LyPzL4y4wXgjiZz
7w5qN0O9YblBBkq8G2ePjUvRxaVXZF96NdaFh/HK/sHboyQpI2KGNS4j+Ui2RtvH
eB8+jKFx3g5eoKScFKX0DH9BCc2QaDbED/DB10md2EYBalHE7zIJW07r4F6cLsZh
PuKZNkwq9y/NYMctw1CKCdd9KJDhjv6ZESto8i8JT1dQZct7kHC7iah+0ldnmx7k
QhOtGkqJYGpu231X0lxpjlxQZqKWe/QDpKtcBYnbZKmT3DcA2Eju99n1uJTHVK3k
uhfr/Uzqo4cmzwl0aFOBUXv0iuIaBv84SEzBtTR5Ac7mnUPpXHciVKaUh2rY+m4U
6SRk5p53o8k1M/8U3tYCdM3ay6cT9EMXr1fSgvpYcmMObQhAZ3tO5Y6aeevpd94j
DAMT/R53hF0qiKYyOCYw9HrS4Ng7jz1EG1XGyKCbNGsa1eF2ARGImI30BIv+LN5Y
NOMKk3AkM3waLx8ciO9c9bDBz/omgoku3nqcRgkGQrdmREKsVwYyNQeL4yInz4+H
uPN4gr/Dh39YfLRIM9OJgCjv9R4KPbX0l3JWcEMXxeGBZqH59euTIXcSLlPO7vD3
CW9uCJfgQOgh6ycmrk+zpWZ7rciDfI5u75P0PJFd9nYN3nVUuAFljyETcSETP4R3
128wNCQMCDFr8M/2e2dEVhyhYzb4DbMPSz5Oenw+9MKG6EFlAP9ry4+38QxEOFOQ
ZLF2y1VAOknKqZvYNJKQi2rOkK9XVQk1ga1KOBdtbWQVOyfPvgac3R2cfKld5NjV
oAis8HMpktrNLDSK7ZJAKAAvBLyF0ckvP4qNzfCkmIOhGQH2Uj8j1RsGoSiCv9VZ
3pQCkZjpmmYmK7jVQA6J6Cb14QY1c3o9DmBoz6HRD1IiCT+GbaGByF9eJ8Hd9WZF
0Ky+J7GW/P5HmiY06Wap37l3XML0msLaPo6nAbzVc3ZjaUBe58m8rs3hkUIr6xCO
KM5k+syoUIdHdqzDUglJqoG3WKLqtLx7+wWyOEjJ1gqkVKLNYXJ6dRe9uOVbMs+x
+9LFl4jDnsLrynKLVE/qCryMtWRjUQYb8CxZyM/TWza1v3WXJ97s3FeAdTwpNn49
BhqI5Nd81J2VW2dZzcB8Gm8HmUUoNEBWa2z8cjwZl8O9y4aJM9Vxw/fdUelB3JnJ
2x7sn9Z9KfZQ0zVESEwA5GLxa0ST62vg0ncohB8K3UXrcVF2IN/rC1Pezs5V181S
iRrgVzi8fHRfFDKc8Djyp2uEF7mIo4AyUcx+kmF9qBgeZMUxpZeloIrsCKPRxi7f
CWFOq+xSf3kHjSzk7zjjvkrN9dVIwl1Q60D/Yto4ooqbW4TWDhrEsQ56YE0kwqSk
9gvhIydSVtFu23nil7QbKz1i2YLplY252yEUIIysjtuVIh+GT0BU5jJ7OOF7YMf4
SQyFEkvoUIl56aKWAp3XKS4ftY+KvzkWH7GjLzpcjPrEpYZL0Ij/e5h2OPOAujtp
SkHszYvSvXW7+SNilbF14Z+MpLTAgMB6OVquOGdeGNNHEWg9DoCNz+QvhlBJvqnn
CC3LhIALDvqD1kD8HM/81ntMbmeIn9cWla/XZ2Q42lt7oM0/BGxyIOvdHzqXEfUw
8aYHOYKUxjRXxLdS242NQH3q9ADI1nvLAN6hk5k0vNnk8YvMHFVEZi6YnbcPdnUr
qkU51vSXFFsd3IGMtqIOSVSlSUJzBoAzr+fevsc4roM29eMEoI1ZP2sbyW/PlUeR
N6Z2KxCCWDmpQVU5E0J8wTnvJMOLCUK0qy51ttW5hTuhq0Mj7CjR0FkuP92xP0ep
ABTfa+cT2MqKxPMHX+flH978Z/z4GtLV3j/J/2OKyuWAFytyn6EQoJAwHtRO8z06
pyEJs+rZCycMnlmD2L+hbLhm27tJqMkIfPFiWZc4IP14GlkmqbqhdSpgzfs9cxAH
O+P3Kyqtrv6iaFe/QeLOXhTtdxofO9LcgJmF4TgZQh4wSBo2jwLsWoj4YBsi77mk
iLkOCHw9UCrfEY1xrPLj029fO1iM6+7LmJTgn5thQZI22Wvuq7A1xPQmPM7+fyp6
hEDhHmOTFY/2VieRNO9iT7JHqWgkyRkuDS1lVmJAc7XgYMAsZ72iaPmdybe2wjXM
2sM6oU+Q/OuBLtWqXR2H2+Dx+sJJZ8mRerhe2tNhvSJHxwai8UaTEvwDqh7Fx5ai
W3krYaNIf9tO90WjnjW8EVpKPiunKd5J1F13gJ3k5085oy/s+o7jF8eNO44fsqmI
UcD7/gcKlqJoDAkfX9FMkBGeNDhxNtYkRM7EFF5XuwiLOlQ1I9DqfrySlS4aStNJ
SLcSOLJVeYOr+vNObhEu/ZPMc/hQF1bHbJr5DV0gbpE6ZiutdsXcObL5kWERJJNU
qNNI7yikW+86Y4syM9G+K3VARzJn21zH4WtwGHEVEKbh+lTSu+093NhWRmxXdqLn
eS9u7UPDZQ9DRJTVunH3hjI/HiwbJaeRk1j4r+iksyY=
`protect END_PROTECTED
