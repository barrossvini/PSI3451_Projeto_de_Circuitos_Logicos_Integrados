`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yFC4kLCQ/zZxuNMp7zt7WHA/xFE6FlMFkatC4e5l6fKQOU9aulfHn6DmWLMSRKBX
GdAaisas/Pgq0egTBxlhlEnNOoBy1JDFrtF4txOvmZqtAE0SQOTCB85KZ3vIIZJx
vtxRkNhzBUiQPu6VQGiHjE5Vbe0mO/WoraeKOWHBuaFEssZx+XbRo70Oz/FcK0We
8nYD3dmpLuCXqqZ3+yEe0zOsdexYOjXB4FShLNoJKbIjp86PkCyxphK0ckV9wSQD
2QpXdt52eJr1n3r1khZgrDP99REchdY9TpXi4TmEcxJYu0D8ikL95kLYiF4dLxPV
vC6A2Qty2tHF2JVQTCTzGNpNZUWJtNt+YrzkMpO8LZWLCu08qMxYdXgbjwbSe1Pf
hSPG+FuqUI17Y8864AF25xaaTbseXK7llPGSpsFt2MeTLa6TJ2/yL7ErBt2hg9tb
97P/X3MdAufBvAJTv+7It/NqAQ9BLo3vCPwz0LJeRu5+mpD/8MXC5QFwBsmIdP2P
Mql9aatjeQhnGyx85qvjIebBnIl68h9RyEARVA48bTl5zrfVRV1XVkiKCj7YrDjT
3xLSl6CvNwCwyKur1tsOeqrNJK6GATLwNziX/MEgljIglI8sJT5AEgF5p28RDds8
9A29YRpFWK57yurgR4XrlFl0iI5dwRaNINrkUfqNYW3+0ygNDL909jGmA+biVKmA
fPHeJ2hUcXgfPURoKJg8eJoNZc/UQkz4NFy/kyKATmOuoi74FrnYlQYEGY4bXP3a
CCGWcmUyZw2e+aRQHYMir9pLZFvuUuYIOhVZNH1gSxMBWg1+qN1cadDnbQMuU7Gq
8qwZ5fgzmMBwsxy9qFyWWA==
`protect END_PROTECTED
