`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q2iit0WobICA04qoXbMT0NEiDOcTAJlWuqKQcFZ7uUWuEy5scr7lNsX+Su/CDyMg
X/OcK5x7Nwn0QUSWbPfiNmzA8lSuyS7kl4kBSRp/3tIFjfykaZQKCkwa79xyFnCY
YJhgTmIznInX7wZ7DijPgw0y54qcNQM8N7qZaRsjLi8DPMa4sGBOPRv2IDnPOpy8
sSqwbbwa5b/6Sq++YTMwgCibPTBNPzd+HdtI7ogafn271IpkG1ibu1JHhvbUONzI
xnV0HbYIMOHKb0JLIhq1RNvLoeQlyIk6ZxvaJHKv2fsYu8eJIgpuy3lcHFxUKmWu
IKc5R2wIvmtZqXsECbkEIHEqN87sUCPUGwyf6EfDBa1+hSYezjjJsspwaigwWkPE
hkKbihV9xfQQOBehDuRS5wRGl4kp5ZH3K6+WlIbUACMdtSnFuXxmmjy5ZCuFC/lA
P220kgHieLYHn/TNFh4GOEoG4dRwQRadgSZXFmEN1InqGVQIHMv/s3BUc8bqU5Z8
6+799S+B1z80hCA0lZtgsKhcH4GUhBlmkbWxRQF0b4YzlPEi0N2IOIQ0alLyqoXJ
yYx8cAvKd/e07Y0EenSSJXL09cvx9IZXdu+bpxJm3KxOrAN1/9r697KqxcS70dKc
eAi9FG2h5jpFo/lLKn74T2CnVQtjCa7G40aqZU3MUMMxjhlZ6AdBdJyxT0ezP6OT
PpiY7F+Nfu5vRhgQFmdtnYtOku0JvCYk0xWPoOUYZMXJFZ6CziSl72x9ZPIvrygx
YmbMlS7jPaeR8urrPNoAQUiIqcQllOiY3RoDoCdxiwDkF6a3Erx6GE7YFj9C14C+
m12VZ5L4bV3u1DIaBbxh+42IzYBZIx4d2ARRe48lvmLVMBowbE+Ssp6i2KKOczNQ
LUgK1XtV+2zdvi144RHcOVPxQjPaE+1ajozvGip845lzaogKymYMm3Fuwq6c9zih
DJ/ZnjRpwl8lYRHRu9iR3MdnLDVpXYmIGre11UxPGpO32XGf3FLwpxy2zntEFR6V
8PcCXLayvzSN61gtVhdup2b4Zcw+z0uTpCOe87lIdbiRqk4wS7Yt9uecIkyA/u1u
3hT0vEVRoC6samPEt+czf4BTErK3xAUnCoRbELAeYTUsvDteMp2yVljlTAFC3Vzg
z8ST8IHGIsJoD5LqtJFbDucb4H6kX9hojhVnGMQeQxwi5qAJRvtpMtr/HW62j745
uto/ioiREEvfHgjY25hISQpHpJn1RlwjaKjvSf47DMWYppoZvpSWG1WNIimrkmQS
8BNUUnT1+OsaJPBF4O6ZbG7+shJiy361OeNnSkrUrSP81z6UV/VYiXvk790gutes
0cjXRHW+kt6uZJY3V/68Y/dQAIPmxen5JRKHgNHHynY3GPbVJkAL8F6FsQhWoCuO
QJQN526nHFyFBuopnSz4XdYwti7A3iJf3GrcRtbwXYonxD//yPTSkDmPGM1vnLRc
OPwf1sU6iRv5S/uG/Y59V2RjNgG+yIMNPvkzYQfCRHQmWqqbNyLdG7tV9pnstLcC
gyqijXpEX9RFgJ7zc8YggBW8BwTyD2G5CkchXAIMgIBNzqX/6Qn5LULadE1UnXi1
QG89pdU2DSM9bOEYk4WBUXqdyyECmqGwOKsyl6PgWJSeF8J/EHEzAhdJ502o8Dg/
oXqcoDcVrgDN/1/6PNsZI8ZjVBQyYYGkHGypqvMI6+NmBDNizCQUl/hMxSicNMcL
aMercvpGPkeU3Is3exzBGprLYbqoKIVYmEZLlVWYzOsYM0mIVt+B8uQGsR3b/QU6
o3QY/v18ZzzkejSuaaSnEPw2C0Ojo21rQmwowqvHWXisA6cl6qoyBCdxtWrFRkUF
JlpKphfUuS0XJ89FAtbRPZdUvdFbQmvq91hu8aHCnTG0MbLvT5/kmu7MWvHPjLx1
PGMzchnZYJVNQLZRhDZJhjO/uN4s95JBXPff7hFo4dPvnkM/tzvqepXRg3UAdsKo
9gxUMQis5SfIvWigistfA9y0AA6C7M2jOlX2CgbPN/uGqamP/mE9mg7k8ml6F1ts
wV51lyZZOL86Xgrzf5Ugt7cvldoBAAS31db5JcowehrEJ+XXDMw/JcRJlvMKGeom
F0RBZ7zTcWDm4VEACCq/z0/lWbHg8xAccUr+U+czURSNl7LbqWCqnP5ZoTuJhj9C
58RqltSUf1aip0JZ9czuQOrsjudf78z/Y/dexY7qdzPNkNlSWlYaE7v0AWIBmhqy
dHp5l8hDdCRmawHZUwvlw5CzTvYtE0OBJ89h6aE45JlvVbuBEOLW4RobWhVOJbGA
ZWNLqX8Sk8qSUA2fSHnAZuRFQJ0ADHFCBQXih00bprzam1XT5SfbL5OiDgAa2cXL
YuVgCYr/+2aw5xqL5aKpAZuMlU5VvAYhAo+2kAjN2jHGoMmZMOV5kkH1lbow83uJ
lyVl7C4C0vHbqA4smxiggIHsdKnT5dRst0+EP8gaHS6mne0i2GXwNOKIkesIW3Ox
1bhc9VLCFOaJcSYMhUoQ2M756JglVnnI08OVdxP3QkCLmeqebwmlRJnNfcDOsNJS
bJ+coFrBlu95o8f9MwD3l+/wGmKL0isM9fc2m4I6ktwmW0pROistHOjcDsZDSlQ+
CRkh/yGAUM9tOARRNsh/rHb1l4z9q2d0Vf4zy6xiiQcCQmOQ+tiKO7UeGPks9c1i
nZf9rii/EKui3Ovhj2KHv+84Mzsy9f39QcLoRVzfPoZErzuH/h+K+fQJYk8dKF9F
dhtwJ+l8nAoV0kSWjrLSmTFrpL75cfoYGbkQaEVRnCIgnpGEiWo18DEy8l6zYqr/
divaHes2JsGfjeLtuNboIsPe55vEmXIqAU7tJAaa1IBErIN+Tzdy/YP0DZ+fP5Fa
o/cuLvxW5jK/ttr/hL9yHYB/fIFVhzGEtM2zUjT/2ufbD1Vpl6wOj3U3YVPgBCP9
viN7CiKkLAoL6XdXTGi66hfrVzv2XUq+QTg1k46hioO0i++ex6r4yIzESSkY5cRP
y7i1D+dIU/Le1dSHQFXoQzaVxIJZrjucqyeLd3Ju2ynSokb+HyTXQwwlLa4OlWg4
HFHDrql3w1f755nxYPgdZ51CvpNHRvUlR23FAeeThw3IarX0eqabmP4Jq0IL3dF3
h7mGTD65U73/d01Fj68CiTmQAGmmk91xcSrgXyBWk12Vg/yD7CbWsOQqg3ye9z5g
g22s3z8g7qQwAohmS498UI+5a2VjCHKR868wHOhsECN4TgUtRLYcbVXeRjfQpa+p
nezaWwGsyAdV2u1J5+OW1Whq7D8QPrFUBhBsWL07/EX0xTDWxUliV0B3AJodxxJG
JfcvX8vHoQUPURFxC3VeFwXkbNknRl7cNMRCZWMJhuGhYEc++fPZM4L5SsHFfNxV
lz6xPXFKhnmN1riCTlcW7L6ZpcTLkrlT/NMgpIPw6ZoYx/+jxyN4nDyaGqiwtglI
kLnKgBuQQBz3rVJiip1RwTM7QUYsTs9csI3DcrCqhnu0PXWXil6ZJlsgkWpQ1QMa
GUTFQAJnqe6SHj/+mbYf9k3GFRUomgM/xbEmcNp/k7sZxOjQyOCHiCPdyJE0xGMw
2Ty4b1EzwyAZFia6P2KuKgspNHvC+r8hARXdtF5Nmbks+NkBqUs7aPUSz3OcMFD0
dmob9LoTGlep20DGn05R1+knba2dcQITB056r+AYX/Y1Wp7NXdYpcCHQVja6RXIT
QxsEOPi6845YdN45CNBJNLW3IK3Svh94HJ11ioll2rLwugkFsjjm1FlvpbkOezYZ
yHZZ2/7h1G9g125PRRh1lgFwxRWbCL6kdQrwkujPzDMqEUnJPEug9TiSp/Tuk6o7
AWxHrAzI5oNaUy5W1/q5Q1i7+OHEXC/wpnkBanPDkcM8AraypDXDn886ME3COXJU
f+E5iF3QuBSoHXy+zXUi5/6TuzYRUVoU0a/z006pNwp7TeiVNJ6PIK205m9HjhkN
QaPyXK/2i/0bRayFdYD+1cZWnnOaPsoTcCpiA9yFURqGQTy3rBuOWf1hxkGuUtDl
NCWWbFJU3FpZ46pYY75P7Cgd/OVe2QHeTajUwUqBvUcSdhBTG0X0b/V54gy4VH8R
6aL58hcRodYVnD8VD+surKi8VNF3Flld6X3oK3UmREQ/QE5lL8TndLXEKiA0dtpQ
QtjaoPI4Hx/PTaBsO6SFS/AmETxuvVkz0j5Pn1RNn4woWgM/blsX53rmksf8ci40
m9g5ZkI8HzbiWxNs/ukeCSwwavwTC7cb1Y26im1Bo00cocfCJo8e+d/iSrI7HIkm
qimnUn2Jwy53oz3h3oaHXQtzkiigB0i1RJh/+yrrl/lTyCPRGfQ+pVp1nRDCKtv1
zYHsfcXSqsReAf1w/nnt2D/hvrDWHmicWGSKbLY5ie7ufsTlIyN+XdWLRoI5WJxD
nn3VSVj276W1j5RZt+NcBYDYBs3YyhzZSTzDu0oXVp27dkfWuwNMQKjFVFspCd3n
baHejLJj6SGlgGKqw1U+BZ0DyLBkqMqFk+I7VFRfaycKA8uDteW4IhNg7VVy89RF
LK5cbuNp0eDJL5qAN0hJ3wkVTWzqp2M2e4OlVpzDuSPlkMlpUJqE0ddz4lOI9Upi
0zjd3GvFD1TXdnDwAvcKIKFGuksJo5Wo+DFzU3WS0vg2WIlJPsTlfkjVzzmlFSTs
fqC8eJTSSldXpsOy8IVcMoVRSeNdjxqY1oHigraKhwHQYgvyVqKKkUPbyOqjrfde
5zMjRYI3cknDfnXsnHiJIujxT+W/kSsNxa2p0rrCo4sXzLP7l9xlfyqpQxQSnmu7
0DqxMQq6MCsXbdVhT3XIPscRx4oDosA8Ouqc9PT5v+OfQs1VjCHi/bjifByJDsbN
tj6fpP5Lh0yWTERbHqYR9NbAcSaHQe3UDABE3SmOfl4hte2B6pwKt2DvXyIfAi2n
bQv3Ak0azojof0VIMXVW+InErAj1ExQBoejayJRuOQ4AV24SnoXzrIp+j8mYA+Qs
/ZI3e29wxAfuwPR86Cv7se6hyRgC2C+i56RBvBPIKq8LaLj6y8DeEsMZ8zrlydXD
r6iMLR/Ank4mmLl98QnBBjxwqNvuCNmUQnbD92dCX5NvG8GJm/YqIy1CvV4kT6J0
A93nZMx3lw0F49cSwieh1wALCK8LH2Mgv+xPyCBDn3hw2VV7D/yxaCEoi9I3uxIE
7u+ZD2emIEVSLffzSbblXJpJ/55PCw3D1+ZXViXjRFWNgbOxvAujkH+mSxVvbFan
XF3A/HXAVNiw1RGW4vA/ZJUay5KidVXin+bFJGTNFL0owwkQ86VanMoPrvRclout
eeWPHhI/zu0NXttqzikFaZIpowuM5Ixj2+XY50kkWt1c9LaYNKTSdQhvZaKQmtv1
KD+1ED0/FjpjsmSrXXZ+gf1EEcVmFn42JIvToRu5/nrHhTeLiQE03dJxoLMtQ8fq
WXziY7XZ16zzXWu0avl9A4RvkmU3DXdi8bcUAKkj0j+YGuGHJfoEFLSv8bRsOlK4
flUQNU0RUoiatoZ/sgeXUHG+VBRhVfhTbN9HZg7sqVjdGRHQaA2GYhFPnhf2viAh
IZ0VIHQZzMW46ZRCiHS9JhO3NwArtFtV8t5s6nesJj2QHPxdcnIw/aMfqFJsY9Bs
pTezfNuKzM09SqVcKkN6pJAVNuz69W2avqjN3IegwpOeGCkXlxHOGjimcO6Y5P7I
hy7V/CaWi0VIO+c3u+srKjJyYHXpCjdqRlIdLwxa4KvTPP2cqBF/YOzmFu0sImpq
NT7XSFOj+nR/5i6c6NkOmUEYcQkQqNeGNR2yiY4d6tKiUo9CpLS0pg0iF4iqOcdQ
gdjOgJSgDGVXhOm2UcJ4lz8plEaGkXb4CR8Y1EuPF96fRyFZYXo6Kts+19ya35xC
NHiB2t9XpULX1a8sSOCLCo7dP6zAqRMQJVNBngb1T4B12CANT8wxj9PHb6K0O1Lg
cGPru3gjuDPNWnjgqLCxnHUm0X5oKL4C9Q4SpCEwZrVh9PVQ88tcBm5tPT+LLoh4
MpSArbHR+IXGOz/8Mrm99GyPcUmgSM40PqFDPhnEz9ngFE7d+IZWTQG2ghgkK90I
Qkp76HqbC7AGh6uLt0ywaeOb9+UxOpKnljpqmYynwETEEi/++NNZ7SzMx4LExFtO
F+pyTl5in/Hroz2w4+myUZv7kzZjpCq8sJCuSJdQ/YFzcn8AYfjp0m6zTUuysrro
ClQSNj9Rty82xDgC3hM/O45mtuOBd9yK7EvXjlb/mXhiCuHi3Jun+/eTq5sRIUPn
EOxxLDuakbYO4q+/KRw8P2qHt13wOjob2DZhfsaqk7aB3sHwS8fV9mWl4rL3Rods
QgQaKgHZ58Ns8TJ+HeSiqjYH4p0xf26DJwqiaahyd4/Cp5NF991nHInGt3si2YNU
fb3Ef9NM4FhTCrFNYV09CddiuFbjJd5GkHhi22uBInMtb+EEDBfGLSnMMugGor/6
u8wDI5CkxL73lRn4DQebfpUSAsmmk59WA26H4r4SQoGbGcG6jL6EOWbbtv1pLV3M
Dq8y5Oqr3t4xEbfVBE4Ah6W13fhWiGI2FIBgp+KS32sPvcPnv4GKj4x94OhReH00
20PmWrwdsGtWL/XgjM14otOK9iuu03KajYAF8yY3X1MYyJeEb7SHfjYFXJScRuCo
JnFoaHvc50/rRPUktG5FGtdT3SftX0wJFYkmSZ1xTwHJpILjTVMgu+Y+jZaU9HXQ
t9W/F2/3ymddmNXhhSgYnfbtqRhu9uvvjqktZJiuRt9zA1tXypN93acDC+vlGMi8
C22jny0CAtvVGh+bEwkBpM01x7xbKwmmWSoXWaqgbXINmgGVlszi1UGCafr2r2FH
VJllrftlbv6I8TcycONV6+838z4a6/LPL0FkuFKpoqWa5d2RZupqkMrJudVkjd+U
3cdLf5RhHn9Nt7FXV68zbV0zUtnFcIsetfhDCpwC/aP8X1pTmVxgExmk7TvpoxIz
9CiCgxmRSGbp7BNd1e4TRYXpMVc0ndgm8VVsZBRaVEzEteC6vUz4tV6uBpMYEan7
vTKt3mlEJ0cjJIt2f8axpUQpyJ3T64+MoB2oo0mFP1tjvsnBXYUxVCWvdbOSDugu
if8+6cbS1Iq8a3aRmlTaMgCzSqglcISqXJ4DunSYqQRQDjtjEzpKtnWPT2/Lq+k+
XCUyI+mwOfx2Bmj4TsLvrMIRR9Uy1HGnvbiFuRUg7GsY7W6krs9vEiuOYBQY0KP8
E+tkRkAorNV4JW9l3nKHW9zd2r0T4QLMqbC9LyotBIYl7ihqkKgH7GiXnKFawQc0
YPnbUy0HWlFil7zyQ6ZYf1oeY2kQ4UWsVv8+roIABGtPsC2mYXEzdZovIRyImnzh
yYb0Y6AJJJWKc6yJKS5fg2uw6E+QRYmBRS8f6QsZse9StN5De+0mxiKXLfo83CAC
ZnV70VuT60ZRayR+13AB0i3YRh+rKC7arYsRMzkoI8QKhvJgiQq4hM+rKE2BFFf9
C+sTZ5slNKDew/TQ7p3fsSKj9kSaB1kKh8qJIOmKi2gXK0hiDIpGTULpzRf/p0HK
gWTwmXgl6Wt/PDuUIjUolgosSQY+4oSYyVYOMk2C7glYclITsLQCluA8hs4UvRUR
HljDhlEyn/IrsOSS29z1f8J8rrIxzPaGk8YWL+GD34E8CKiCXihVbZxHdQ1+7FSO
dOs80EZDVGZWGvy20WN31Zu3br5SvtSvXOyehrMtplWBp6eZytONAJBMnnDMV9oD
qKR7OhVNxbSbl0Lk0HVZQtm8WHdFFuGU0JmThlP+aY3XhiBWQEyQ9zBAfILJkR4n
WTM60aoCbZpBZ8ostW0Io4HmTjeHHeC6ml0zNQ58RJBUYcbcPaZZZrnfg6MnBnjE
7EfBkv3AQG+TLER65UD807x/Xq6PbBtaZPQBq37HR8bVjojomaqeY9eamJSHVuoC
1NOA/JD/fSMU/rlpbxDAqHHuf1Vx8dgGbputHBux+uPb+0BGnLiPKohfsbjkhcLA
4HmyX3JdNJXHpypR7xwFFVVigPW9yLSOimcgHz9P+FviIdK92M7Kf47Il/PJuxUd
G8EbIRLhPA82WVUVITavwZSXG7gbYfn69o3877izjQVZNnPNvNxYGCM12ZNDBHQm
fbpCZ09TlLG1R5CCk1wShZ1VcSm8KGbbkCTp+d3OuMNPR8sEoqw9M452BqFnCnSP
uHV02B+v70BjfHEAMvilOkF0jLnwCvWMNvMiv7fhSL2W8vJhTVeClmM0OyWKshZZ
eqYjinGu+pYqmf7WkWy31m9NgfF1ZXpA+eQ3Jz9pbO92LrtrsuJbsH0b88uFmvzb
oOK1qaemxh/3XX03QhmG4e2SLC9olobZOoDDIhA6R94me/k5kg3BXnDvS3c/EH1A
k5c/b70GQD66PvlaQC7Ni+ZXAKsfa7S3iQUv6K8HJ6uxWywH3QzS8OTAW10B8GQ+
enqARgQHnUc9EzgTHjEDOZ6Coce2l3iKddMe+YnhTszCr928TSqz7rQTWyUz1W5q
qeoSDLwWGPgPU19hQxNkuQp2b2WPaF9zQEbxyVsx+ZhAaOBYhS5SKdMiYF55FuIh
mNilkDOoVPkxoH6Pa849km/dBGKA4jm3p+0AN//jV1BXIfJ3z/lEuvR67e0uRiS7
UQiAr3IsyTfDYxAekkZ8DIeNuZa4OR00K90W0YH/UcSZJ2uMAuAM5g/1Z2fLEzGL
xz/yGka/Fx4S8OyZaPIQLNWexaROxycjNzIq9tVZ0vNyFeE3GS2me3Gg6Rk4VxZQ
Y12P5F4VRy8qamqNzcprMpUwFxj9u0WTINb2I1c8BBMC3cywpb0ZNmU4WKcTRnms
e//kU2iyQuk8dE5/7759+yXMZ++X/3GctZQohsxwVDUr/yDWgWPqLbhxtA8BTOh2
+RROLZmoyMPCYF6MsUSHNtCu4ReoGhzPcLzizepxmA5zBlUeciDBbgR+Kx08tpZ8
9X0qDYaBe+92aepx8UZThvSk7Qi9QDwIDHuwMdjdskSL8wV3u251R37ooHuIHgDV
iKXVTaCkKtwyhYVrS+JQJjbEsi1rNBt74WiEtSslcFhDwT65w2ly0HHeJ8+Rnx2S
Xji9gZybm+SzqF8vcK1h19IkIDVA42tsMMMpibL6RlG11Sf/9LxPakWeNSi/LoDZ
iEcUCCwYnEmcfodVuv7JW+5E+by8L90XPPkWJRJq/Dvtf6auAy3iFLzC+rdOMfEz
1c1Ju/zk1lCenhqkheKST8hFxp5zB5hyO1Y4sBJYvwHgxHO1gDQikKvfOwszhUcr
WkQbuw0pVAlsBcqjAir2mNzVHHKzIhZ+RYpUJ/wA/pEBKB/RGfAP2nN5O3ypd8iv
wxIV+EFYPRPeP84735CnqgwmcDahkq7cAlP4QFJ56blm+OmnShj6PG+zs/Q1ozIv
uquJepw8Zt1AVdpOXq995x7uKiGRxeNnEt8mvjGRMRws36uHoaUomAX5HVGkX3aW
MWhvnv5Zh3DFQAV6cwDVyfRGBfTNsaK10wBDfREw26qmQ2E829S+Wqh0i9jAdLoP
jN/mp4yumSGW432I+WL1Amlw4A2FNtyPUSXHmUwnSODq7eTKNCKWhcSTh9fRniN5
VAs4HYgcYUnOiFZ0mSB/kdv5CaWVSSp9by/6B+FNyBMFG70TooPeaVo4Byu32KoP
mqpLRn5Gv8A7oo6kedVmiEl8S5S2kL7WutnVf5Eaz5pzGHX5zI3yVhIdxhcFBOwv
wijtbqacayoDOAHCKhEv4c417LHTY28MLiYsFZucA+0k9/2IPI46teu2Yapfjc63
G5Q+FCHVZg64VQFhqc/pP2megiIH1d/6EqZoutgtLRq+U7N92PuVK6WythSH4evT
QSBZw6VNswkCajWXGStyJTsUrUz8UClgBw52P0rCHY+Pgv2/8zoHL426V1UAt+C8
9w7Or7DdpKhBPJ3x1kdDEnmcmSzebpBUR4vI2i2P2ycs4thUjLSfESTySTUhxefA
EcV1GsjVzlQ0v6U8ojv22oCa5SQYG5LZA/EAq1oyu5k3h4dNNNYqmFhjeZABji/z
aTCTV6s1eWASnBpYI8t/OfTL1dD38Ii6Qp5zDS1K/O6m3oc30mCyKIRKCEacWtsk
w5pJsuHdSeirzlo4wR2yAQxyadSC2FE6OelpO6OVRipd2nRJepazfRsPtaqvyhi2
VdfMaQazhrGva4lpG9Qqn9cQnbc0wzeQ7kYUQRl37HW1QavOd8AfrCNrwXqbeJAd
KZojomHBO0+kmPo/+7nyH36iSKbA1JnDF4fwxLXq/qoiFQZeP7uWm6qpEhyqsAdK
bTZ6QG6bKXFRaHmJ4h5u+vRTsoieWFMncIV71f+C7Ac91yhmo3vfyb5NXnUJT4h4
iz++YxnLCSlxblOzzbmx2wHA2mGOW8C3Ch1OV9fWgtHpzAqHn8xYkZeYRlweb6Yr
hUFYE9Y3bHPln8SXFtOPOXyIssgFmfuon2hlSpn1VAE9478hfUxRqJs7quMQ4Pgq
AzJaAYTictNt34PWcclm9r1YtDG/bb4IZIt+IjuGY424fhOlV43XFPkASG0tyRr+
9rZxndelHIZ1rF/twa+aw8sacpSuhC+Gsy7hkGtURWineJhUB16uBcQITIOPB8nw
C5gn8YUo852GvdYOzq0wpe45Ie6pQbOvBlRtqfzBuIovvWdHJInKO3Ut2/g4aYvj
ImYmNpzWVLbmZKCK3M/uuwf0dRpbi3UdBdtAJqOedsR0vEr+ONVB12QlxgwrmBDd
UeFksSFVWecvM8x9IVVnuNdIwZMMp0PSjQ0Du4malSEdkcmHn76y8F0NSfqcmqDM
zzQ8Vh/bGtq39nfNQJ9qQjJGx1kXXa576Bo7m9eYF6Wo0jEtNuwdo19YrjWju/C8
plT2B7fUvO2m8+keGnpjhcowkyIw8wQaESgCZ8xfbaxvShN74Gbhmtjp05d9Tei/
Tqa/IkJoSwW6JayZdTS+KdCPnWP4BiR7yIR4/bPDavpGCf6DVLzXo4R9Ibf150d5
Nxjh354p4H7fB+ggpNODMICyHB1l7EFGLijHqQaBFU6WH4D+a2bmwiavnU6SyeZb
J2OWskHuAY5wGT/fY9OW64KImwTBC4QTaDHYbOHFovhgbMM8QwgoxbdpkipaiA+R
3j+VwOJe0hgpoPQR8rz+jmkx6fzwzbaIiwnqmDbcsAQjOFGtW222iUY39UgT3iAW
zOX8ANuhwYB4YbocMN0UQ4xVI+0RrF7/p9rlYlYNJ8qDx4ycVCtytObte0/iLm41
VNZPkKVh0RfUNXYOPWVixSCOjFEO4BzVdhXTKW35UhwzdgWsx67gbgQvFmK8JhTa
aa1j1HJ9SgOQI/g/th1VikvFiUhWxPpSkygrXo+S4xEuPW88kjIus2xWMkRTJNMa
CiedZeeXyvnNmulX84gMwaNcguVVgKQzz7BVAz/YOZY7r5L7C8nKrAFI5W/3xMz5
xmAiM18TAH4o8xZ9Guz62q4cm6fuIuUI7vbYGT5nkDmxD7Omt8V1xupJC/CvjJaJ
wyAcED6MUNmuUlT8BrubSLj2KUWPDniP+L3Uf7Zp6zW8rfWIyQHwCTiEFKdcDMGH
1p0ZU3XagqhPI/YOpJtSzeVwgr5tcNT7aZ0nE0F330bmYjFIzrBfRvw1sobbLJmQ
vuSjloRRavJ0OgKdnIykG5g6BWoK8isMvGOhkFNouVeHHG6rKB5TVTvmA+4gnFUr
+k/QrCECaiORZw8Qfs58j2h9/QPtilYomGI18Wwz2pF8hGKqPFJslJMgqfUfRiaD
R+rNyyJ1jnnd6G7JQlPZhHAo+j11Hjx5gKdJ5Y68ves/d3WOQ3LUovNjmOm6YV0D
9fB3omWAKgxU26ecHTduVyjZgAjD+iLeErpaDkelqke8+IU+XIh69GNg30uTZ/0J
S05I9T1IU99yxrlbd3EWxxwvmegSiEmG5QdKEgCkqw7im4fmSg56qBPdL9MXZwG3
YM0AKYEsBBYZ3MKycMDj+Ay9NCmtNQ1q44rvryNvhDx0R0RmOYcn+ANeOrcqBhvV
547l6R1rg7ch9W25KbJvXZd0TwWfITdQcXtFxfIwqp1+ksNC6/Ja4LjjUA6BQX74
TEddcqy2x7fWw6y44UnpMkbuJoBWs7gSas/hg6xa7e4zPEWKOQ2ByQSXnSMl+Qpg
RZG8mkgUxUL2j3aoPQVvL8lKd3xJdqQRCeTmtdnhJyxDUJ70guT70jeVIS5yPF7E
FUkAD8LSuqngoOleNAsLp6tCfuURBdiqedwE3eDoFX1UsLs6Wk5aevcvyyHUb/JZ
3/CcfTicSl1hps/BWbB3wR9fWgrcqjzca+oWBPCVaIHSOCmJoLGJ7dCOQjMIJxGs
owRkbwwEq5FauYZyaPvLKVHe069GXBAqnW9qukpmm5oPqnNFyDHRkLOVCOPa8+uK
+n4EltMQyxBQpAOiugZET4hD8AU/zpC2gf3YjGIJa5hHmEAD55RlQwgQsujgQh7l
q5vWRGZEbmYIpV9bf74bUJKFsSnIB5zACjxZp6ZsoERVZT+OQpSIGvAN/QSzB1QL
LRTdxZ/jR/z5IgkA0mBhr66A5Q4GPEk6+l8fYzduIP6lcmmvmfrEahCcXDF/F5l6
1K9uWr5pKs461OVoSGcw7HXcc/EyFR5b4+36OHoD5RAbDJj6m9KPOX9Qvj4SK81T
frlg9juKcEMO+9UnzdV+3/Dswh8Hx/B5hBwY+yrO06/pTXYVl8g9QBvvoq+UZhjU
h7ru4hVLt11Gkp3M9b6zSavcY5E4/eXb3IToXGHM5WNgwrupdqsW3bt6pYVqUzts
96VLQpy0VomT0i6rSyUyp4RFOTeuXkAu9ZobSnH54+cKbm46De2DS8EISDwEpMUL
dyCfSpjEZBxTJYi3evHS9wlQUm1YHrrvNSlUqhhbTc5Si+c65fPYMpd6YsEUBp/e
h3VKH8ZesR+TyGWXc/oWmrnBK3ngABTeXYwPxv10BxLpOKbFIZnRyzBNhT00jWIj
FX4fWshGVIo5IRUQbBVJU0axJvUMEuySPGDkJRv5/R2P3fBpRLATD85cT9Efwq1D
r4rMJVBmFS2Tu5SerPcM3Rxeend3jc4i4O13EToM7nNANJqlcbJwGaMlRY4O74u/
HGiVmDRZLTdahzvKi917OiVAZDLSsAyLpfrz8PrRXnwRaUmuwbJsCTdxGAC0y77X
6e3MzanGVzCs22czfrj0y8HPWmA7Ey0HqL5TVvVSt6dnSxSiJn3nAOd0ezlnIZDW
IfBDUaaTYrgEd5qN2175nc2wRUoMoXL5NItPGzsxETEEhTFNc9MYXhgW9V48zxdq
blfFrcnC9y26JwYTwDPIrf+zGjv3QMyAM6aRrnYs3nVNFeFiDgWj1p3iMh+5IGYG
LrVu3oxzbldW/uIGf4VkGC4V3hCnCIfifL9DlEA+cGa2fG6BZWS6rszMacbNbMpo
i0yFA/5QAtcP/gJhE2IgZWLs0fvA+WlC348nVCnbzZEDMzKGVqdOVxxFgoAwOFoq
wX/tkyNdQ05q1+WKROhwMtEddjnlmkgXi91IAaSrQFzst47MXQ8PA29XA1S3t/4f
xxRRVVYt7i0W86XNlXacl/hFgIIkjmWB9jzG1sclVb8Uvlg9//YfMnmFyZ+FXRrQ
Bxl4TRkwBVRsD03qtgIWkgWFuXox/K5MVN6hVFVggPZff7yF6xh3vl3oYpQo5Y7d
3CuIePYhZ8Mv8tp86tHRCWTb8a6phLEiC5jKwfBHIZzlTYWv0FZNOrMT0uE9l1Kj
T5zh0zU0BjuRVCnrH3rf/YY1t9C11Yh4WLHk19vVI+1Vos5D3PgDMjN4/WPGGw+h
k+jXKTSceYWM528k8QQ3pfpUTokZbLBJ2YkHTJn2FysSVZtbzfAtuobSWR52dTVy
S2Hv9dJUbXE4l55/wLQvg+WnyAymT6dZ21hOndWtAthv/VdAT8/8S1JCmwZuTlL8
T5+KkcZ3V4JozHG7cE3ZI0f7qm5wZoZWfdzCJJBI7UqZMonuna1RJn4A3FNVfWkL
CSg/y5h20z1WCgwj/FCxeuCknbCdnP0Ypb8XYTAiPzi7NL1ez5L74JzMqjWmm9K0
okRvLgMXD+ksItuGjrBWYnSeAcAtv1yJcukXyv6yZV5veP4tB/ymGrqNilyAUMwD
e2S5WqcsAKSN51XCCTCfqEaoK1h4aOrwimvzcZYBlcpcIJoB7fLXc4KcXgweRITL
l2uWNxUZBHBdTWa1cTduslPtgYw8+vbCcIkBLJacGi2enP2JRxbfttlm3hjaTEyf
FzidYjiYFsZ2G58WaRFghzLoJ9TL83RklUNfClVWv7WLVWVBIyjVuV8vGuDHTxit
WBrqHycssEvdravsW4HP0DP6s+6X6mWGhx+CI7xZeuVS2h7dGXJnGjfBxM0qivze
/3J4/0nUtoSaBd396uYemRlZ2KJpVATrKgh0CRa1QWFEmkTJjeAiE3iEXrhTvCJj
/KYOJQOW6yjV4CupVUmMJU+Po/F3b51kFwvoe5rCbwVbczBqYmzhXS9/Xc6O+lMr
K924B5NI6lRdHwCzPdIirP8SxT5fXwO8OaFdyazX8LIG+nQNIpzCqrKb4QQ5fT0k
iw5BHLx7ZCGj2EFvk8fZpfKmQGx+Hqk8/WwMYhRgx/EzlMDvlAPIsIAxXQ1771rD
bDhqZyTXFD3yDSkwv7BVWZfqyN6HY/Qv7Q95v78CA4vUbTj3WNLsax7tl5oDYpoC
kq7IGpD0//zoX5H23DU8e1JMlvFILhTP++2HmET+ffeIU1nfxZa8uyhF66zATqVD
CQ6mm4XIKKUBuBfoZb3mb46RtlRxSGSLyHLssIL7s/7o8OUOi3FDGKb9pF4cmtvF
UPzzSLk6xuwFWDqAAa6+3lLg6u6W6Qr0vrBqrhztZWWVJzksT8xjZ+EkUDdNOP0d
M6f1Tmes1VBvuLsUpXX6uyxVm3euoPWj00F8JweJvzal2Y5v1kwicI+Q2j5km5yy
08Gb9JFDy2+jwxQiPQ/g0oAhP8mPO3b4V6Mp/dJZdcCiRjMnAUB3/L9frSWJILJz
ZAJUyHVCkbZQciXXVggO2UFA5A+bO7M4u9OcvFxF7tja1ZSoMfrmGNfvTQ50Km9J
+4i3cbIFGwglhWmeQ0iF6UelhlZBjD0Bxw519c4BtlJdD1/MVBwHoQ6ORU/MZcpT
XG6AdgRd11LNjmPYRIZsjkUYaXZIMTp8oElEd0XRvOOgKhuZ6kCey66NPE4gBblO
U6FzW9rweH2aiEPrz1di8Ibk5+mz/jUoSYQMqu4B4kvPmgFrPniZKiT1WDi7GpBH
cYSg6zXIcxlxeT79KMd9EiBpwdzR+qVLleZ9YrAzDRFcZolZKWAZRuLmJUORr7BV
vAKH6YCpItRRP/4gEwR0NVSiHPacx4aATEeYidpz3AzFUfxm1NTPpZU2+nYDmwzK
8knKN30RoRohwLI5sotnmtj8KaYOOHYVHs4Bew9MKR/r+/LX+IJRCLZgbXPibuBr
5hW3UJ4xjb87tMchpyOsfWSsKR3iAEGdxWYcKn7BgYjHrQjSKuGXsElVUNp0LltO
gQr0MvkrRUheS7iZ+AoNoVILbqwr1Wqqwq3skMuj9IW020RrAvL5u2YhLBMiJq8h
1jbn1Xvzs9N/keyvPvXUbLjSNpLyAOZ0ID+9K4XwyYnp9NwxZ9RTCPnKXGrXsDij
Ymt71WBstlxLlTYl7KDg22+mQR8VhySAATEaZIf8zaeBAwMAxWXcU1kuHYH8mdF5
vOaTnSZhbyezfUeeSoYZazPSQANvD58F3BW9RUdJQbedEGzSQH7PDGXwxYUQ0DKN
xDTvHDhITdaJHs15tgL3Dm2DQ+dT+ShDif27paIfVugpQ2Yg4AVM3Qzv/Achp/2D
cj1Lg/smimNGsfsD773aiJTNvXQ1AAHx9vFEnPT3KTswlNlWC8t8UuNvankWdua5
tPuWQ6OtP4Zfmqc5IrcuGNwb9vVClvli2OfEAjrsZ2uGMuI7lLB96/zMxqyGNgng
KZ7YJBVg1aJCQGTwVZwKhS+kNAO8yd0+JI6Yk7OWrUXYPD8VYiWAHXD1moA++dFZ
ZV+6aRaXTXleEEBgAhvYbTW+nMar8amC4PHGIk4rCHSTSRjsY1HXscetefmkY8Z2
eNpB96/I0a+3E2nZ8IgSoYQ5wyKH4SYJtN2C2lHscrK4ASutWmL2PgUHFxmebasx
nqC+lACca9qo0P64b4y08Pdlq6pdmovJDg/OtJTB5CCxQJmBRoHm4nxEIFy5+RKM
u4k5Gq3aKrqkHY/Q5/eb/yP8Dh4QyVzI1CgVKFEj/FC+qXv88HbRLopzPUoCoZTN
FgjjugnQiHg++guA/fypoXLCjcRaot1esNALiNTjqUmsUXk44bK7uaR6EDxaMf+t
dV7mTwr+Za16SZRm2TeP4kr0Nt1+8TqO6Euxb4dVZ+Ku8fswxpEDcOP9+bVspqOP
+GW21h3Fk/NExGh7EPj3c8g+S3ijcQppkEulCelLFaEnW/yMA/rnV1Dsx1GBMdYh
QmcZHLCoE/Ds3+eKt9Ce5+1MO3pMbeH+EbQUEgj8KwTzeirtSJREyGRGZFZgIXLD
IPAzmRt9ckngfXhrkmgmQgKpeSkTeqpFLQEK/o7Y0cZsr5RDLV9pml27HdQxOJOO
CJIquER6O0wDbRmC5WivbbXAQ2Zs/1yV8SOhCz4sHyLTdiKaZ2T9o4j3KZnFxB+x
NUv8tdYEt3cNV5+5nB6cYRYEE+ftNjGTbgmbyvBd10b5hL666E54oDXRsXi0wdlL
/rpL3tFMvW581iASyyIeHeTkoCsuJUqvm121elMcLOoQY9T7sa4NFagum+vMBPKu
Nct0xLNZZmdrwLPX64yJxL2QiKdBYfmBNAlHxm1sKrzc2s2j/71dazgM/aNUd5Qz
Wa9YbRK7a56eq+JY8JMgIc/9yJFmD8c6TbvOjSek0tVn13dmrCRL0RXocpJ5tpwy
kXkn0dQL8s/aW2A5a0G16WVP5VC0G6b0C95xCog19NgyFWYO2Pw3LJ653XGJLj5h
u6o2SAvTzjOizMltFhYWhRE9y0eEAIe0jOh5PPuSe0jMJ0l0J63N50HuGupdOWHL
c63fNu0iJlObzKXHSuZbYShcrWFgKDOoREQK7zeqFpTtpzq9u0+rjOHyVv9wdLJE
SacGr1/AQdYg6ut9EEf6m5M0N5/ypoUYBhMDzQKBPkEdcRAosmJMahjaQdT3I2/D
5P/08Mps40Fv25+YGGaBCpeL4YU+PvMOCTxzsGcFtKEUOTtyaeMy8bg9yLDDYfiK
FE7HFDQTGMgs3AL5SZVVpKQOBi38pOvrkqHKyQcUQM2lkxP4aTzoKmiU1PYbtyNT
GO6DSka/i5GV9/iCgRXFG2ooZg5Zwg622X0Hzam4bwgqymNGetAKKOB7h1R+1IiW
DQ9Bh2Bzw6eqgLUocLcmP/jhwpXWovmUmrObfxleEip9YCkRYRIqkQSzjI+o2Ndk
bN+4+Uy4c1ZQdy8q8Zcoa/Yq8xS7UeZ0EpXEiAUQ24flC1sKtRyMptIxGtemoZzM
t+xtv+zHwEXw5kh5NCO+N/4D502asVRb7aiUJ0wwr9cgS/XyBe2E9DBn+nOTSRtx
XcsYLMprgsSUfmh4f6X/AVHTPoRm0JFvdtu0WLAuCNiXJj3t2jmRf7j38y8SYr3E
nRBZecS3AxeZn/JZkGA/HFN2Gkk9mXtRaM7vBXjQXnIdCkdts+dDrsAuJp1NS1g+
2ZaJ2VD0fZIg/9oiO4XVFduQO8tv++xtmeO3VjVzwZz/j54Vzk/ZMLms+QxZj3tK
L/jycz21rMH/VUGFkTZSSaBTJcy8Ttx6ue5cXfvpSwtqNttNM+4LBiiRV7/8+kMv
xHH6P+6QjaIJz/tQF4jJoESNEr4gbyr1flq+4jrrNCNQLlwaK+9aIWV2E5ezyA8f
8mor6byGg+guHGopcuJ6os/flajkQmxFwUmXrHP1yeCFjb7jTTddRl2Qr9p5saVR
m5ho2QdwotidTrfATMzNIBmwWHiTyGHON7FJnC/xYIm0Ezu8xHl3J1YxUbuWPU/q
LH+0wsmmmvOeb1zDWpDMqzsIjhfH63oerXtM+JfQSrDrcniGFpK4kWaEGrR0Tscj
tLoxIc6wkKery6rmD3NBQE1V9i6wrPtApZqbU/tyZ/XJmhBDG2vk8bPNVKvYErPA
Y2Be6NOmiMWsSD6hsC1VNs/nwXF6CxLpcoksNGaYpaYYE7zTyQ48s8FtMQpQJDqC
jhR/oB8lZUHX1JIes+Qg/qlf/4hU6KIv2FdCCuuz2ZOKtRaaNFit96DRkRTGCqtE
/u+dYHWWsf2fRVlMdh7XiPryEoXqB6TF9pku2dfozMGxe/zAUIPkcGZUVNwOJ3JZ
66F6mMGj+tuaez7Z5B76MHeiWd9Ii5lRlRXmrULt7+BYLD7ZqsT1BwexJwOSh9nV
xw2KNIrRcKb3ACS/DclN4HGYnqKUfr+mGjiJniVfF/aLW9H0x6z8ZA+6/PGDi9Rv
WvU4SvBUIRb/6t7lmJx35+84BUdQgLgcIxq43l8Pk9JoDDuFCnjk8fO+ABfTXX30
rKOOd40ZxG+Le7x8qjWCYlPW62DemNXViChxZT2+9y6fVGrE2Q9DAScSQll9iqnE
un2qoe1T70AZlGzVUz+7IZcXTC3NPrDx2ZhEJcnK+woXMis8AilSjAnYb4TS/qa1
sm1+K8Z5EXp0rjuRgexqwtJYyMfUOIt73Re5Jf1rlOHhTl3eRg4aZnHut7uaRMYH
/SgeVhfHVqvbmD/G6WF1Gr0ISonLmTvQChRWlkqbinadaUH67BCFPcOVY1ITGHrQ
NBQ2IOPq2Vnrxift92rrAmCtEMuf5uxSGHh+PNOlQyCuBvTuHkVM3RHY/5AxzJks
nVtp1gITrLyq91OXX74/aM9/hJrP6IdXWi645FbkFxqJ+HcP8Q9vWUd4BaeUlNqY
RbHbf5REBokGJEEgPjC3csbte2xobORlHnLGQnPJRTDS+yx4xwW812HdUJlnY2gU
/zvn6XlCJZRUDWXrZQ5c1fPVGe/4ZzN9zGhPKkDlFA7XyDDT4zGRNnDe8PiJTHtT
xAoD6qTqpUSW9/Ozkc8QIM0XgIC9SF0xQWDzPWlel8YeK2HjZo4mmEcH5W2gP8RQ
CSeYgRGYsluBwKoNAbqZORdcfLtd/aOoqs0/DxzsoI7WMS9i+vGTznKmqPZVnlK3
K2Qfp7M8YuWhl8Yh7zxQDJrg79Rha16QxvjyveD9sIL5lNXHPu54QlI1cx+fFY1z
3bkd0GQ2OT2Nf6OWSrSN+xVGi4nOIjuz009PP2N9oaEmJfXFnPv4WQ7m3pCox+m3
JM8UZSwRZp7TTktBlDyL1PWyYDZwztRkPrsnjw87bGn9idG7iQXIwiACizInnCMh
6dVvtg/xXjbw/VtCzegSsnSA6bVTWGySbYeSYLU6nMhuoXvbxtW3eQYYeelKYBJ5
g6ixfiYNP1QCwsO8bAtXa8BXF4CFiUOShZG0WruqgwSclxZ2iBL85fcb8vBc3DJu
elWiRS/c0hlBxLFqWFqiUCULhZ9n2AlOwoavB+xHmYR7gjKWYC/qx/GFWYyaPqFK
x0q1vUSLWfRgit8ikYXJPfbBt4FHoG8Q9gT/3UoY06ZsC/Mlo7sC/7F5JFfXXhGn
yxOw4jwU3Knz8W3fuH7bIAFTUSluNJQBSsgLpNOKRfttwqhjY/142a18F9qBOf3s
YQWIvcq0VxKzCJrjdgn96sL7UC9gAUWU9SwG1ABFuZI71th4vrkeukbNXHV9UeeA
uL5hZiZFFH2kPIyxPeR/1WeQOdinXoiYM6ZkQCdrF996DpKLPPcz1PuJVMBtg0Rd
/Zdlytxs5VPjJDE44CWdP4XFacIyZc34rkwe1Eono0z35aLpS+c8Xg7XH/tWafJc
zKc2ItrJqI3rC8xIUUsQV8Q/3O2GEpSd9qsaXQES0mYtx7dRmNZqa4Zg1Fx+d0bc
LUoVeBl9Q5Ijc97mQONqd0PhMlcfFnkTOzaxwPcTqeoGbW/ct5IoKB2vDKt0w26/
VP2An5g0DouTpdT43u9M+DRQV41uvTY5Ngj9RH9pap23w7y9xfvvBym4RHZq8fIE
BUrAq+YtsAPTy2m12FcBadWd3VvTthdP9+PXnmt4p6v9owwgsMyZMS1m0hLdn2TG
C8nYkj0qCku3QwcSFwqg05Cu6EL1LPNzaUvSLk8IFjV5bHUYy71u3sOawrStfX7J
9WsEPvdER4+c7xFz4htL/bK01/C79B7X+pMTO3p+/WMhm9ID8gHOVA/J6KH87dpM
UPWUED6W9WlhYLZTdlG4RYLLSILJmU6ar8FUTRlxT86X9NnV5fA6ndrNQnbJSEQ1
G6FqxxuU1xcmKevxQQ0SCav9Y35TE19pfhDoobsKjYrLfx//1dXmB2H7rSGQu2a3
AOTbGJaUO8flwT9QuU5/vX3OV9wf0MHl0bkIB2ufioY1EeHZicAH8LDRXl01HiB5
LHKM+lrr0BFU0bn24/CpwMD6hcdqYa+Wo/SuZdQpjAObAgsmtoGfS5r0FDMWL96w
vKAPE1PiHHl7ugBQcYUllzupqNd/ZgmGh3caBFvjJsV9MTU0qXVAUYKLq+pl/40a
xOa5ZL3KDptw71u46JQet5xpM3p2LG8kX2X1QMTm+2Pdk3WYG7GgECedHARFz9ml
RHX/QBPcgB0/u0mpTJz3NBrdQFRTFj3LHm8jtFVBuylHV8jSCJzk4cSeFi3HjvTa
aokKSuDVJNQxC2ZPdyqKkcDw7IQfU4FebEh27JD0qJtGMo67CG/v+kkOCwG0dRuL
kagCgrqBC77GA4SiJ4SoEVxoJBnuv8hpbXK162T+HVNaNzcSDUj+IBQqC2Cchvza
sVIwQ94TrF07XRSkp0nugdPUhglqD5bmuFOeAJ0VLLS8f6zLzyqXtn1pC2xoSd9I
GW3SDpW+0wdaRH+mbKvGMjJPyR7qqvvj0LOFz65PmfS2xVcELJ8tt/XBY0oyrUQJ
p7WA9revcCCLHupxchFEVkc3EAMbiEuSVXvGfiG8WbzHEW6NwyW4f16qb+u2gB4I
SpOSyy2yc9uwth6SMmOdvJb/yPUbKNt4xAyM3XrYpc50JyqDt7K0fsVXlTsCG1/E
whwgtPK/iTuz7rNkPxIAezvUGOp0H2Y0YKCzAUddjHPYrW9sjwJ5o16GQuOj+saa
oB+T3eF/Jambsq5jok7SmSUNwWkwXyOylq6uFYHt7ajr3GHcLrc7ptNegeXQS6wC
R9nqBtBYqhqp2LduckHKvduAB+vCU+9Cv5YKAudZMGJJhJybt9dVJAKPwB1nkg7U
4WtKhWxvJxc4oPyCUDq5cps3UgWpBCUbfobj/lVNk9s1jM9wxzvtCIwQQyCIzUoY
fjAFZmvepIce37u9ij62dd4kX7Oa40qeHr/buDsDHSTxQ8Y+r9deZUAYMVNwecRE
SO9ExkbfATCjbYxpPSsJCv7ptm20Sb7I6nW9nehi54WQ99DEdiFIwhP66nimsFVt
30bGfPz0s6g412OyqrF6qr0fb4zXh0M7TadaIWivbBWCabTkXbaLtDp+T1MzMNtq
LNVSZtGko1P108gtx8BnxD+xsQMO7ODw/qS9HsDuf4yKw1AEWjxFN81291qNprHW
dPoKMUE6zN7Z+ErZW/bPrCHO0KDvBRUfvd4eEgxrLLsVKuX5mVBw0tYYVyv9jJxe
WzbidkZVt4asSwbCCMwXOiCQMf/VxgUWEcXIJCJqf/SYpof90yLg0DCVsia6nnrs
/ji3cVlolbRSO1GdG/mbmS8ofyGK68XH6Xkn5d9QdKA5naDHjh1U0t6tKYHZ8Yim
TJ6kUUdBc0mSt5MAGCg2rX5hQvXsNHcEQQw7bctk13Fm1LlMm7jrV3hekl6dU0jd
RO/oQ5UeKx9exY575ILYcdZOlXA14wTspG9SZkEVEE5ApHG0vzgw+r/AHMbCJOsd
IUnxjvPrZgOOfUyH2dOfuw0gKBAWae+Zo+09mQXcBC1Tuhsb+ekgRZbPQAIWLi83
TcutUucPLYR/G2BeT4kvUmxgrP7BKkHMWSUyz5PdU9J1oaxWiXI+piDnqXATY2F1
VLjyLpbug0lXkaU5glm8+M/p+XIPMrOy4FmzGDjoyfQJNpERoS6F1vm40l90bPjY
VECUcL9Qn7LCvzMDjhV27i5f7uQmi7RGtl/LyZBIKcDkHvsloIqJb77jzH61a+Y9
TUsxGIckX3U2x5REfNG0WeRlcyCiTngW2aqMXQ2RoqiOoGiT9/3UoPA+NbJCTmAW
nJP1wjKFjpqZyuAc0Cr1Z8sM4b7HO3NfAV4A1mME+qBq63KpIPX8oxBAmPVa2y9A
qpeDhmGQg+2rmCtPcH9KaggDezhb6W/hUVhS+vJxwgWRYDlltmN4lD2dlTW1pmV1
dQxTnzAa8rRgUZjHGe4zrUxIVHEVvAniq5gfeTIZC2gbhe6gPNLGZuBRxp/xzcVH
l1RXlphNHG38b/w36baQXxOdri00Mynh43EcYFTpyhHFATI3yxUq3tv+HguI/6Se
yeZTdCrA15VtkQLfjiYJNPUM4oAt2fLUTMCHU7h8BSL47mv1wnwTZHjyAHpyoisd
4Jai6liVXWaw/m7yhJ6dgMwK8QivFVB7DNr+2jD0RKVLwffDPAg/ZuiADyz8DO8n
KlxsfawhvLIAP+0eMuozV1f1f1Pa2jr3lRTIrD2r7x8rwEDNADr5WI426AdGfOkV
IFj/1dcfVEasKFJ6WPOrRtlR5jCP3/rd6WnDUvLUBMAMbVrE4i7mnt430+cpH0u7
bssoRHw5NylhxlqdPlQh2yoBj6uvTLyAaKFfXa4Rj6olkR2TZ1G9Dnbh/BEkT7bK
thQcJVy06MNEXNuPrFX6QFPrdn7Et4PHXUvlVXXnhQKXuW6BWf7ZtuPAP3DU8UUJ
pO1M4ICtHzpLPYAt+HwmGaXfY5BYFR6AijwiLTrU8CqI2yrjKwgeqLT1kHmwwSBI
J1IoLhJlw1bbUjcXMGy6xzCULYUL02mWti/lcSVfc/Ev6XtcxzUu+a+FhFP5SCFX
VwVXCljAHajakaauM4/hbpui9s1k/edn9SyV/SZo5Ip7iwPl8DRtB3ugp+naD5mk
JksJ6mODXdq9ctzrAEjh++RyUHCRF5fzCqZFlqeRe04t5rNX3r3/tOrycFgoTiif
pk2JfM2Xc40YevxTPc06ilKTwCQ6EuBNriT+fC0w0PPdU1jntnuL/wfCzIfzs1wh
xp+xgi3gHXb56/a9vFBeZgeXExlaxSrieKje9QA17y+XdnCH6RDooYD27Lxg/rl2
XW178otdqqs0SzE7TMwrQcpNvVL92BnO8hJ/iI8TPh4dbbipdpgHzqZAEjKq53og
P2vdwy0QnXlRwLPGOP3tq3jt3BnBUYV4bI+BvoGDPJcmEn/R834ir3RC39+31LBW
iYyN2Tqq5Jc1Dua6QaxepjPDwR4HuBLRiPS9bZvyExgO6tZTEofs5HcrhAaOsmaM
7mMD/mYymr0d3l5Tb0P+dOBco6Viu9mXWFpwCKtQX5UHPTV+6TlIrOmN/VyfzT5y
zGNeU+k3PUa2EiYnmCE0ODA0BMLsxRpMqKd5tQu6xe0i5VEmLQfjkYusIEGEKJA9
jJ7XlKRRe/SzpWli9El0ZTZFcF6axvCG1ly4Dt6IXKNhWrYMKeBbkTD4B7morBA1
w37Y4UtTqw6cXD6l6uaw4w9zwDjU3svumZwquMQSv+1RoZMKIULDP4EB+1XuYcSN
AyQZWNaAniWFREDl7Kh6/PsKgbz2bUrebzu7iluJsiwcEdMq+gIyY4fBO8dpgXuJ
HOey//Rx1tEZLO4W7qwqyByZdQ6HPPZ2Kox3yviDBby7BIrs18PfCF8bsH1WhlVm
gjpgxWHv1Gl7Q/pzIpeCLb4S2jwV1efKaHatQ7Fj/PlI8onVPXU1llIw+5dwtv/1
5NR6RiM8beRVMTXsmh99x1kd3ZfN0yxB85jdQbpH2nloS8GWFoyENsHR8G86rqS6
WW+iSpcMxLGN2ha80Mb28FZUvUeMTtzWHal5GZjCV5x10YwsFTpjcTjMfTP7VYVU
DRJtQWlekBzjCxvbRBk5Woh5tMefDbcGDXYeglFYhOGAX61NH5u6wk4ZpImwl5PJ
Exu+/aZF/2Q+D0IDhf4WcNJNoeCpE7Sw5qqDa5D/2OeQFixpC1i/QObmuevykrxU
xSkbvdeG44j3BNtWt7SpUlAhQOGGurOcnikaSaJr/vTFOSqTwuY3gURxPpNqyiIU
iJp1MaCohBjkZIWEh1kM2e+2hNGXGm30iR7+VBrkcxgKUP+2ttP+Nanir6zpGLmX
bm+ZX5NL8keWK/+n4aI+jY6ntlXDCriWjk4d7d4VLk1e4D61neNTUyjLKry9g4bl
ww02HkYB0fCj/kC/BwbmI9+p+Kny8cu7xtem0f3qEjvqNf+0yXv0U3yNggOw5vND
h6vKY/vP1QiSVnJL3S20Q7hegMRPWNWKkAO8M2eC3AB0aSBiAFD97l5AaBIGdkUs
vw8jPcm5s33eCpV4KnMlO5ZYii20awEZol4EOhTD/bpwxbNg+IZtyi1dbp7d3DVV
P2WnulQ1JhT+Wi9Wrtbfg1r2rysCWigiNr/2mbLirJKMfKpS7RcaUIjOcadGpyGl
glESVz/wtaHfD/LvxFSoxUtKSogdRzQJiqTbiLkN2iwUYZb+sj9RBmAsE0AHPwf0
QQbZ/uGN8nK3jif/SKNDzCvJukUcJ5r2Lp3euvymA2odtbCEkD1z0kd8n3K1K103
hOBaqTni3Ibehjpo0EAhtBI3waP+rRMkf5fQbTDXCKEYRBakHk+FOtZdE8CiZXY0
Y7HHhtcEJfycVhv4qjAnZ6f2WZeZQMur169m3p/32hRQPZ+UtrDmW7Fgd3qWAErB
kNtDWMpAiw2zTt/lr5Qc3t6PnFOWn5JN32QJNANfUtVeHu3Ps18Dzg9JUYWi/NMv
l3a6xrOj+Fv/vGpFAwroBF+i1CwCvNUJykBAsC5Be+FArAFINr+k4iu7GDVfgY7W
nnLs5QtRwdHyi3XaTLqadY/3QKKDt8DFVFi4TWp9HeQJYDNwYYjueQJb/Aw6D1Z8
wzpykVYQefCstOasSmO7mUixu4SkqN4fZKqn9GgfL1yhFiaa7H9yLZ1ziiDshpyo
JWjAYRijLcrj6qmDT2LWQhQHiq2OoeJagx3rJJ7OvdfBSmsNjXdiT/BWBJGP19C2
AC6IrDH7hf7TMZsl2FjCIuz8gq4npwLIURT0OA4wYU6/oQ2oiKV5T29MCkQNHXby
ZLGo/eqN2OXCdpRWsxl0NWpk1Cag+zsAjiuUYYzeybNch9pQFGhPFgayti6n5zRG
YcQ9se/caHSiDKKGi+4m1xQY6Tgvn1GR2m8aBUrKKvwfPTkVEUa32aNpy4edKTik
EdUdXUx7XJ1ZENHjVxTJi5HXHuya/pRDq9OBw8WkTCEvuBW7/k22aMx1YPAtZJQI
xrZdc/rplbdxESOx58y5DtXk2DfeEKrx4EQdda9kSE1j3w51CNmoRDLlWiJyny0x
EAAk1S+OrfzDC5ACdgFaAj8/DePbwgXSQH89tqUEnvlpfTkp67O7o+y55w0fPd+x
ZRSRQVJHzxHQAV2yPgEL8GPxT9O0MoA7VR5zPvqxeGvLjJtNHZJQUZsKsySAxLK7
ilzrFMsQ9AQuRMVdZgwGwPBYhXHLjP8/NWKBFacjuIQka13DUlLk5Q3tF6jYbo3j
24/C1297NCbjNOlHmKaJOVv0HGe5aHauUZcNS4auwF0OCbtcFVhM8I9QYK3tzVCy
owxIwc3HqkgPmRu/7hfGUt7NgMTn+OpkLDTO0X7Vo1MIt9COHmw7vlmqphOuto8h
T66gknuvAi/Lu4hCkfui3Hy9lEecQtSsOc2IKQMlA3f8D6kIpbvYOPFVNiz/F0Al
2SIqgsVrPTxikr0/MleIH4YSQFb4hvumzDFFAbWTl84I+Nw3nl7vtPIKXEy8elRA
PaLUjkJmS3YcvNKj9dq8MgXscOKQnI7H3XAbPfVhVsnRgv11xBSPmX0GN1WUTOdV
HyyZ0QtJtsGZGch0dXr7+1V6leOfc03uLXS4LrV0zhpea5dXC3bS2F3o+8QH6E2K
mFBqzAJxaGmsrCxCw85pMU08Y7BolQ8/z4Vlp8Y6Y9SONw2Pg/jA7GJw4R1CmOq1
JirRjrk/ask9RCgyPJylkEftksek1jvVXGYzt/Lans+tRnVqWb9Tgph952D2zfBE
1ZmXc7XQt7wudcIEjsDYQi3KWS8qmyBXSgD6KEpc3GTeOR6+TOpBvQUETekMAk+K
y5pfo6v6F3UD8LMyMInatHUhhzIuFGZRiG4AUtVWXMidvF7o2crCN3ADsnyGeOHd
id4kRg3lByR0F81eg28ZKvXx+Vq3pemqCj6M7KC/9+87t9P8yIX462gE0SOf+uH6
H8+rPaiqR0X70qLK+R4Sh7775iShPaiFAN8DQlo3VJxAxNhl+Y+yKC3vNb+F4vP3
EiOUc8eGu4xlCEuEv25PdhAsgz4XqqncgUpoZSst5oEpQI/d3E2Sm7JytgQ2q8B3
CdsPFm9T7+dh+GkJKIBR2hE34IXKe8hGQ7iGODbhyA91UZU/UkupwvY4r5TgEflv
8TMb8DkoT1MqchAjyRxgN6o+y3WFVaPCiO7vKQrmuAKufviEzVMh04Rc5FGRxGnL
nAYQ916ftfnP6Ao7D8iAJAI/Bh5QbIw48LZTd857JiHgZ3gH1tgC9f5VHkcyNQ4V
z1mZ2ewtWgFqQibbjTQDEVlTXiMEHThnR+bBBceaFUZnu9di98plyCCJp9231FPZ
BT0PLsHa/4jjfqy1IDzTDMIHh6+UHBPzDfaeHkTg2cpEmmi1GwEV+7SelhOyqOwK
QwbFljt9rPXF+kaXHc9/lQzAB8njtqoU2MQ+PcitIRhgmhSHIjsjYZRHuto9s6Y6
OBz+5iD4F/JiF/xmpvVWgOw6OXStwU0SDQBjmUwQQ5EVVf4X+n6xndNYhSyW32KR
Vj+frtg6LRfh4hbrDYbGgvBYs08+9ehcSvv9C1Y9qDZPCbtCnOJ6+9OIiB0r/gjn
8G5Q/JqS58sIo+k3FX5b8adRY7oP11jYa8JYCzFsT3bo0pH6HoL6vwTgMfMObERz
sl60Rpi2KbSLNCp14MQec9sYC7NsDtCw3w72NMdAzu5mZCLFP5+lhTMMQ1VExDWH
Zinylb8CqDtK9WJehV6fn9qIMsE85QCZq+mtaSdfgnYJyS3FEL9c0apvFZ6AQcV5
4mHEtMnfyaE7HIotdyFkrbIRYrvWZba3mvfFAtELt260aTvG0+6eQL5wgNvI4XEt
QkTTWhzH7VubnrwxMN1xEqW5rz/55H807tR8tMtEWGTzzZv/L9yq59NfaNDn97wl
zyEz1ujntxkwddJfV9GfPxHxc1Yfuq2lYa79062fLRtL9tC6lO9EPszTqoMtzIeF
ZYGVAjAU6bBZ7V8rwZYqRXPKvFlIgo4Mv/QXKA1BTESRkgqyi+DgIGUIFAfCC7nB
iME8oNq5Yn4YHn//F4i2G4H3hVDu5mN7aaZ8B9f6uVuM0wQ3RssTSAWkTOgIHd3d
evgkjTaWZdGHgpmM2AcC7dNLTE0gK4P7Evkn370lS8kDr0STYLWkQLLJtBPcWnm3
O4oQucLn7c7A78GrWfG/rRlb4ZVDXnHrm1L16fyPEaFAtqnpOmJwC96+dVFphwdS
KJcIhBpyUQ3ygoicGf9JLdsnxO4naizb+5B6V5g+b3y0BRFjPJCobY9BRJ1MnIr4
UBakaT2pBBQWZdMbq/sUd7xo0xJGgYhnXSRCpMIuW74ujdxOjGEwCBW+A77ePHON
S/X0wMBrOy5JMW0dQAFYzLDR49fGY77jVAQUn+HwyjT1MXNzBd8t06zE0ZR9Ob8d
iFpLjRhWqRXJQFz4+2GOnr6qM/he9tv65xkjm0guue9kLyBlt9NbXKJnT+8Ioo2B
5moJ/TToBkyFUz+eUH7p67lm5trslDftVP2cgjLtvyeLzD9zbCUle/qVrm43EyQV
AYAaBI827yv8YEmM954c7Gcsytsf/ceQALO99qJSpQWf7kONEb+5nhn6PNuQcAhd
iM6PvXwfSoyU0m7TFTgxA+y0YnNL2sRvyPFExt5q+u9dk6460dec+CWx0VXSUW/y
UnjgeJnLGg1VMCYJiFa/eSpo0OBsQqCi+jkZDVbJ24+CpAWaCZ7Nr4WaapZPq5Su
XEdlkPJa4s3NVjL0azr4aR/YGxnRDVLoV6rVwuKo5A4tsUnCtBeE+NVlGdQgl0Dx
Q/NvlbWt2sQVDJSUX//WN0lznV2MAwtrTsTQdd68mXycBzMy/gS+6576U7MwjxVx
NFIoPK4M1TOUKz+1/Cfd/ivoika7izhnobTPNbplmaAe4sIGKgfURUkQWTUtX3YK
anpJht2M2q2VNr8kWcpgmK+DQJ139dD88gtHFU4YklYSFaZvCUBLvjJQCvx5tEUr
lHODtH27WYGLpPAOTamR7hW6nJjkTkavmoGfO8YxlpExFrZBLNNcRVWNvjlgIy5g
VE9qCteh71dXKdVgbu71iQGZTAlskmPjbmTztvY0q8QJ01goAd5v41edAjnHGs4m
lvuOMDwHXM1lsTQoJ/KDFGaT3jDJw6o5fFfiNpEvWK+DY1phzI7XPHdqqf6W4T9S
HptJfqsVsy1Wo51t/LYS+JNGmyoz2NvrEapn6O9K3DjAy/39zAoXaJLAJHc8T0Bq
6pL7h4t0rsDAs7TgRbstWRLk3vV3G4gGsNBF81RXQief1r6BHhb90TvYoiSu5c57
gtyaGSg4BKItuK41t9NtohyKWa4LsYxX+SKYkS70DM8AbI7SqPSqgj1tLmMocyIM
+GIC9+cVckzJ58ZVV2tUxnKdQVN8Fr0h93AFiNX9LMH2ht2TA7EXLR2nvP0GLB8C
X2GAhbTpzf5y0N4/97QAZBoD0Fgagr5ICKaIPj5Ew7n1+XH6fm+USUu/hpnZGcze
BtRFrOcZLIPepSy6hahF7o6IutkIwncrRIcIuq7d6LkQ/Bthvb09swMv5PsY4Jty
nx2r4bMaxae/2f/8CH5Wete2mk/37EGth4TyTirILTl+X4NHBEhpYdj+j0zwLN0S
1+Y+RjqXMd6jpLNaPRdrldjjbFS5SXQgWacOWb9NMvIGMlXSeHngw65WpAafomAO
opc0DUlHKR5iU7VcwroVSlsGLfPjfRfoBkeJR5c6NglER+WAMZpvyE4VcZIMMNOE
8ubUH24puhUafa4Q5QdXk4MuAelI5l4tKsskEVn3+6G2EbdH0LIoyoIZrRJJvd2V
Iixy8HCHTp9z1Gp+vGVz5aGhVr5nRHLUtOyUlhflub2AAXkXg+Kiu2RW2oM78ksM
0jvQyXeloM3s0/QhpnjVaYF3X0h2pnYA7Cce1wrqsch2xZy/37T+MHQcFD2LSBhY
6q4Rzd4ZmRGLfjblQoTWUeljgF2x3jdCs0d/U1aTeyPLkv1xTRxADpi3R0nON7iS
sYJG50NnOCptb0LLnBR4b2an51I6eMm2A4LGFNyQIlEbRts4wKtaZ3XMFvq+7O9Z
14CdV0kyuFn+4VUNqEk0YUP1/mCEtzJrOhsYCWif9HoiLvRV4uLvcQzXtZR4XJp4
CfHcCWXLxtk6q+M7mp0cOhaCa5P0QuIYNNCx7qO/qIDsXNBfGGP5KsyYHZ2qdky1
3iCr6xP6phULC37T1s5nS7nOH1U+T1+jUCjg3rwL6b8WhIaar7puIjskSe1ZstXO
b8rP1NJ+kg0WdvfgtOLH/jNJIU2PPxUeblfstwmJCoervNhujRASOXQp79d1txPV
tayy9dXAsLkpq9r7yPBBTEqgtzdhCdX+IGUEgYQr3f610nPHmIgFtiUJ954yBRKN
gHxcFSfR1bbSga521iLUy6JtBef23YuFmfpxwWM8XXS5dCQb01zTCQWG01fk/sSX
M1W0Ht2eJNkzbA5O98D82THsy+Dy73qdM6cS7P2HbSWu0XsF1vN+0AXzW1CZhbwW
IuxGAGQ6rpm67f2NTTq5WZwGVtOLZlYbHTfwSqq7XzO69hJsyKdHeDH9Kl0zOJAm
JaF8UkszRtx/7SpD3Ae7HQjNOEoEo+ad1YWhIP1Y4lcOlC/3YUsGEoYMUhJjZOuh
XKDHCgwRAfeMHuvHK07fuMqvqray1tijOTJ+IQuTyiMl4WnZDtPf9dHaJUG4q/U4
xR1QSjTvtbg3iSolleKfI9g7xPY1v2zH8B+saz2ttZCRDf76OBLl4TVC99RZ2Sy2
ev2Hu3idrNfnTzwX3jeIzA3D7gNoXzvQ19/Uwm8a4LLDMEpeGaEHVtkh3k6A6uVJ
kGk1uQzSOSbMbsi7CvQbYk5u5p7BA3rn3m6mQeNpf5zDGevDI8EqffZ2N8fsVzDX
IR7TYGLaPj7A9yOYOSZu2uSdnu5lkOmdrpDT/FWcDiA1qIe/t2vMi5iKpy+s5Ufs
p1zMXwqbTQliMZTE9df/eh7c7JXGPX9wJLVWE6vl+PfeXNhN2+8YcqhOVddLAItV
KPRZ6gRoJU3uEpef8NXPSD0QWNEFP3D0HfXkYlnIw+b3HoTr9tcvvN2tRSaeKHJn
EdsyUz+xq2rTbO/cRvkch381SYe4WcxoHMpjpSaDT5GSqa3Gbg7wrgMdxrOcnNpq
cYoBvZx3IZ3E4ejAuvL51shuGmw+hOZx5BajYNh/tJfylww3lzj2nTVJwo7FIcuJ
jqVrBn7FonF2ngYcrnN3RTok5pOgsaanrt7eFU2msYQy17Jtna2m+AqgYhWfIhbl
w/hoHvh8z53tbX8UJBUYHzKILJnMI/e6nQoXaM1CfDn1A96s07N86/CYBmtlDter
FSqw/wStJN29Jox6PfqDVwiGcfZpf4zCMAglpCqjyAt1JIWYf7TSMT53wdXnylVX
GSpl1iaguVrgZeLL+mKUYfWfn+Hhsl4rpxsxozjW0qb421dt5fLAfhTGxLgd53x2
6ToGJh2KWoc3R2vL0eHKLWSHRqXs6FKNsYBl9gwMwyfyaOH3CS06fLPoQ02xZte1
V2wdXPhCtfcOds37/dsRVavchDEr1vnMJi6Tbhtf2PksYVZxb/MnMq9tRzRrFFiA
e0ekRVTyjSOAlVFtvDjfsEAhmQCLI5Cij6AdAbemwaiWWkN5Ws+wb+ghK+11kjEd
JiyZKEFSXACiso96Zx/fNMto6jPVbxzXvvVJ/wHbCraXs8noXDrB9td045Oxy4VU
Nx9celU7Idaqhz28uHrBvbrLvx5aFinaijuAHVltza5KlT3mvgiRJ4RNc8bKLlFv
QLID2BNHjsKB6ZnCYHc402Q4GcVRJkeLK38RlzpNqy5761Npj74pnOWQMjQfkW9x
rIJADwCFU9aQhY1C4o9EI1NNrbi5Uk+cWJj8OeUAY1lXlOYWQL6G9ZDJAQgcO5V/
FHBj4tda27lfkIzuty1WAo2tFTJmm/X7oyX3s0vbvTN2npjSuzVpcbNz1RoQe0kr
+meaqZh95vQceJn25oZ/J6tyEnCPDwGLqJ/UughaCfPCYz9xXt9e2T7r2mPGh6Wa
IsCp1AHT/hNKS8ujQIYmmQxlIegu2nLlk1pOOOjuVmlHRNLuSh1//xoUG7k4i0ng
f3CxnlBwmUcj3WESxlppE56xLl2ESsIkVPdaeYaO/L9oIAiE+IXmJrZ2uPowaJtf
fW9RQUnjBoDQ6rtjUwGExZOoX3fRqIWxTcHPwpl4MsnmYQDmEo6e5swofzpBtghl
g0SINF5Rvc8aXo9fFHqwEd+38J8E67MwccmN+3u9uSL5yfCZbmHOdBh9kdQtAYyl
ye5mPu3Q0LbDJ1cXyli5SP0pTyuzTLgtYQ2KKI2nXNs4C25rVj0ndk52JcoUQNKc
YsWlXmf+KXrevYdR/JJfO/E+s7APmT8SJ52VIELUs7vsmgoYP3ZXwYPgy4EI2FQd
qpgTuAM6slGsW1IWi9OnVqXGqOoBaKZQcqpdouhUMeXQ9wr5oyjASkooF4TqmxU8
q6ouB/B9rg35mcejgHrF7Kw//F+NZqPE0FM0KqI3+CS4IRQAXMj9cvpXp4920wnT
QghOSYat283iGWA5T1yUs01Gc47MY5G14AFMeAUR+mrojS9GnHSsDuiqQ1DEgbd4
ECGiHLhJHfleZufu+E/FjxFatSyPmcbObp8Z3bCq34IBZVu/7vE/qitDa96Zd4ip
orjYSzGaDL3KnrI6W1X/WUTkAOWBLWznN+WQUqJCd8/HqecWHE9SiwRAFPSHzrWT
WhUkpF2J6hd6Z2KPLXu56WH8/hlDdbK9tyISwOaMbJ4JZ5Yv2L0UHysEA1isYd3Z
djj2RfX/YRVHP8JtTGdE4/o1eUxcdx6NJcQ/F2rDptmr/91tZbfMDULH7IJ0HZZG
ut39QFwPveQqceyIWsD7REzWv3FFbn/st60aV/SNYWAFfIfyUeVrq7xEFbWQemC+
3mkZf+WRqnnybS6gBWKeojnB9HmrlqFAxDG4SFJIrvFfBhfrj+He2aFbmkKjg7tC
Ndf5SDiT+zbX6WkzoxhSwXzIQLaq2zuKX9y02XO5dsYL/ccpRuSqp5LGO4x78Dg5
7aj74/DLfXYhOMkZAh8zA7/0Pq0k74ZxGuXLQY8okpZjGP69eNIMaaTxiOnZs2iC
j73vg/9C55h6e/hzuC9FnqxPkA/vXQ17BRgkD83wTBK+WrFVZ4Npq01kB7Z4dLHL
hMfJ9k45vvO3qpFB6I68t0wayay+tkPdOwCslZpA92OSYLumU8RpvCAm0Ohpjbma
XIf9J4JkqwNi3SmgE5alCWNxv7gFAxgKK3aWEHCZDrv2K7bpTq45hZzKhXJ7tek/
R57GV2c+p8k685K3jA84vrJtB0Bie1urBeAO2h1HA4wk6+2qmvITqW4NfTEZan2J
MOz4xmsDiA6RBSAbHdKRPgW3y73h3DoJZeIt+cqRhLDuVhpwawk38v/wlSSnieNg
YJbFW6s2pxyBennJlGvH6pZ5i1Q0quG1F0cd6ioKJe/mQ9jRoyN8obOq2kw6RHZA
OMkuyYl7JcYQYI4gMP/ymUxT6xxG0CE2ceEjNZegJOt0h2gMw7m81DgkIH2nT0OD
IvQPm1cLWD8LqgMJpsKg5Z+EOjzUWQ7698B6nKw+uemIK2Rn1lmcy1BGKc0QlP0r
5Le4r3qEpmZF9/S9pafbmsz0L/yOzCCBy8D0CVnNp6jX2v9ldw+AKn+o93+8wzdA
MLr/Uogy/lYvOOj3K2lx1UEPinhXxhrMTza0+tw3L/1q5e23is+3rQLHp+Y/oC25
q/06edirhSL38EXM5fjaN5MokWZaP9ERrW3CJ5NqL9HXev1QpOnKzODa4tN6CW3m
7WZLYYGdsZbEFKQrdgC/BN2/Kfc9cXXvjolZ/yuGiY9/CWvMRRcoTJZx2drJz/YP
OUC9kYk4Pf4mCmTq5tSNSiM2XTyquZcHNFg2F3X3FGnTQz17cI7jNfGL9zCMm9hR
woSxQTLwaCr7kmLYAi1sp7KG9f4gOGLCIpL3PpDJ5gZko85boQKrKnYqF8lcm1EZ
5P9EiIzwkVPo6rolInxGkmHvEACxIpt+jtswfFGupMLOzw9xnudSkVoGWytgPRU2
W1bQOhWCbhS/zXfJ9YjS91ay3M87Zw52Oomr7HYTLHkDZhhI3IqJFcUo+ZApmvkn
T8VWfwMIucMqlNFMFpFS0UVYXutudoZd7E7k8CCRTKzwaxIWNiLNYfwn86h1EojX
53oeWi8HYgxaX9gEw2X7R+irc+k47ZsZSwsvfEaqZvLf6BwBd1tkR5uv75mIOfBk
TVUZcFQ0ilEM/AaVMpK+36QBjTCsKulesxwc2EKNh+f8gSZTjGhKbsPJDJSnwwO0
03Yr/ZtdChv68UG8pBC0kWd8svWdv9GBroxFxsOp3lKbPxhKUTjTa6LOCoURwYQs
jbTWbLULFog873Sv6f72VJ+P+xTdg3QQsNfIORJXUEAn1Gqwb1z1s4VC9YR6HAYX
Q8R+l6ZFPl10ltVVUfpyb+Hj+b8+rimMKZb88j5VPNdc6J2azn1Bbn+aQdBM9JZL
Vmk9mZ8rbmbBB8pr3dzdHWZSzurKoQbWOlU06+w6N+nUmiGh/twxwhcyUBCRkbHL
VrR8LS/m5ONXmgxwcdaZmPcxd32U6KzHi1RZxqSPf6nFg8R3nq5IPn5terU5e+60
BiG3kRCwFP649BUUypg5Pt25FWvPxZkTNIGwPkRKeIlYxXfjRpYHzw4GoIn4FAE7
gnIgZIGfqZdNhSBH0D/xb0Jd8fVjv6d3QPkO1CVr8OTDEvVHp5TzysMprrKHce2P
DHe5YoEROv0NEmqFoXaBtk9VoHTOq3ZrzyKbMRaG6ALjCGpHdr7tWjjDg6q870dc
Jr8K5ki52zpri7tEqa/SWzoUhIUL6dAB74gW03D2tQHre8xETh6AmwzalGwDOLrP
AiZsG4aJkOeXyCF90BAB4QS8Aq4O0ZpXN16coKmDx1/sf30DGa6bHp5kHsNaf9yU
6oyc1Y3EiAJWbUv4IPlOosRsao+N6ObEVf4TCHJYkGyI0ePoqQvyOY5pXFjyB1qC
qCQ3BdVcYbdIEd0aCDCdvOyEVtUU1Fwvhpy5MZZP6Bmy6zApECWDMW2S6B1IlBGm
rYy/N/o/7AUSiQ3ZIBCV2Ed2/Bm23j1/Y/QZKa1oaDWvLO44KdJzoOgF0biv+yVK
C5MQkWi7KMq1+7RmH4eyiWwegJjd95YQt7QL5HJth9opSDo3zpXykzgDSNex7jYX
eg8w9ngLTaWbw8S/iOuAaMHWUjBNbyr3acxULIE6CSLfFT/4U6RpoRCtnF5Etwyj
1oPVVKcEgDEMEFszenNm7MYufB0FRXEmkJeLeDrEFbkskkZOzVeWdkmIhyWOFGSt
YnCw6ZPIPG3r2Q8OOyuQRkdAxyB9l0rCWm+24d5LD5d/8nKQyozLE4BbmEGCgjbL
vsQoSbsVxtjhEqtQgRMoLd3nXFi1JF2El8MPsLOG9yor+MURBfiIx6EFqWV4yBOU
MbtDHonf8qjRSP43+jg5CjK60Q+HC3glZgFn1qR+TOPveuGV8NvwD3bJOYlvYBF2
tkpiqouk5egJh5AyQmSGzl+jacxj33irAK+fOF4tTCXhw3okzrlYILzczEHscOQf
S83rwxu+MP0t1qjJNOMh9XatmYQzlhGaugPL5s5pLZQQvbLQzrjFwH7AvpDtB3lN
B/dsTlAJNNGLNr9N6TUQ5v3p7xOazW4Pa8XSQwa3n7ldwlY2H7lnKMoFLVquJnjC
YKJ9TQaEKWHfItbIipI+d/2V9adkGSdEWmaAcdd+cdeA2QxvLQymN+iXKmg/78ux
xCX/y4tvqF0bcL0z2QSIah8p0CYXUhAfIjCrLa1sXjOleBXnC5vParx5aUhw4PMo
WwwJswFFC6QGpCDAv0MGVthX4LowIncPu83KL4mcqt/JGr73fzrPsze99UGBsaZM
c1urrCsi0bDdlkrEDzynZ9ernpS7ZpNm4Yrcf92HfAgNeipyVqmX6BEcdig9+q7D
NUxq9dpeWhTCfsDaZSXFRm6oipXVJSMqOL9R349jgLOWk7otTCyXDY7zepeXBcMo
vi6VF2Y/UoB1HBkl3kX9kdYUVY0VTY8a87YKUmbYld6ctcffUHBdJjgY6rxfnazL
m4d/2y8fBxQh/5uwXxLIfd301+EY35ShphcZHa1qApm0svHGYiHJ3DXj2yiHgZBr
g9mcAcL7mh0wFnT+h0zQaPEbK3KKIgIirCw00+FaDTcitxzud4vav+jBHBCeLQOT
b8m5WfGdEQWPH+5IHXkKa6irevvNeH84wTxqU/8z9fk2Bx02aXxfVq1UVdJwtZms
BnSpoXwtPKuF3G1IRFlg/oWK1eUKH1FRy0XSgdJUXG9IcWcfFFRlYvOaeKMmVwCX
j3tlFVFZ0qHZYQj9THZvtJ3m2hSSWHtK+JG5WgonVB4JOUpxSDa4L+vSD8CsY3Mn
oyufC1i2oCCIVHXrklMO8IPZ7uCqI+Y5TiWQwGWYcAvTSwtrDfxpZ1sqpPc6WgSm
4zhl9hY3GBrSiV2J5YL6bxB7b7yKnHiU2vcqlkZO2sy1q5N4tUA3/L+aaci/mH30
8h3G6Q2SQRXJU7h14ydFXPE/a6Qfzpmc5Q4xVT1UKnTRKCz8xdqmCQWuTD4gFZ0N
bf19jbc2mLQ9qdpQ5euKUwgM0KkgQgVloAlo+tGeUwB3ilRJZE802lIPUq0FyT5j
lg9ZTidu88ObhcHqPmukZOGgtKHnK33NQlpzoHl/oitv56AaYeJ4I7Eff2a7kjVj
IleXww2vQDRiZ4BFWUwF92YKRXukl3nob8X9WYnlkjAlg8+8NI19HsATgbmYc9K7
4G12+z8SeuGaPBSOciAUyVMSeb8iJWxDBsGIH5+Zg4smuyx6tG6tN3toFknt5hhM
GJyT+SrPbT1XAVfBDdjJ/S18H+JBm8KUXEJ7NxgptH4RjiFfVAWFWXHGu/inrnDz
QToPg6f7irVFHOeU7+bJPTyDT9NIZ/oB3b3ltlI5CdaP/aEihIjuZj5vVi9Aoh1C
sNECrn+5RFWs98n1VtWTqoUx3g3pjSWXCr7+ypIQkDmG7wzpjwqKlr7CjpLDh+9W
iHnOKzmv+bV0eUuLCUmAj2VDetDcuhc/jitzerk/o0He+c3QAwknpleOcAa5Lyl9
pz3yrnibJSauoFmClq4mwmz8DWNafWtaf3y+NlM27lWDYPOGsj6wAyXFkm6xl1DA
vEUK51SIpeAyz6aORnsOj+uvoOyO4HDj6hD9r49x4H1SJzKQp8xpkiXAln7aq5NP
KQ6w8yWVBm9IrdKUYxErd0FxIVqxEY5XcVSkwHVRbgmFP9osNILdygn3g0k9U5cm
C2zNNfXF6huVRXNk0vwISoGomCPGUVnhpqopKXuD55MRZA1ZJ/F4BiQ1m86/+Rxo
WNbzQkeC36f1W1UfxwhdFf0xigfuH30PCxNtyknDt3T9iyVAew8Lv614cLZBujmC
/JxIyQUILuGVtL/Oy3fn27yBnxFZI799Tl71NmPtwdOVn9jwPvMLU/2cffI5Wbk9
emGxI3jMMuh/RCsAw3qKDIkEsW02YaUJck3SEC9Znjk7S2B03Jit9ForKO1zg/C8
EZXezaev6X4GSZp912iAtvXFeSTDVF95xQMZv+EHzg0g0OvF++E97ohD610ujSTB
Ln7pG5t5LRE93Tf7mlXDndWrrKbTkgh2NrEu99TmfzROxnmzEI6DHYLQ+DpJgu/y
Zlw5wGzVA4CjpCS85KUXa7pDam9BFBRlMd/3QnI2qLnvVgpwLxtbp3VhEWJhv31o
w+46WbZXLocZmnsRN9bCiGMPf1cbiHQbCHPEsjaH5n962MjuI05uoa2Qg8zz/Qaz
N0pJPaBGUZJi0sMtKejOlnQt1ki6scsnE3wHArjf6SbLrKmMRKBgIL4lY1Lmlk0x
8U3he/wowHvygBRwJg0qZqODClxLaaBMJquU2EyPRbAY1JCowToygFyPvkce4Oln
496t7A1R5+14UAVW5muvE4NpdWOsuG/FAmkIuo5kAli7X4bcGHX8n45HvnUCW4kY
0wdCPTTR+HWpZ6SBrXQrntyUAiCwOY4Nc47o7xwSbbwrC9hSxzix/fON54edfD4d
J4cAB/rve8YOfjMTomyvRE+1DatGpretn/GrfD3GKnyAzN+0/BXRVPad55eW8qyV
l7emyyoB8COtrx9uJYf5UY/EbdSI0uxqu8cYuu3tgIIBSDaA0oRffG1DGsfjSNEI
3nLosoDHFjzk1ERE/S1OwW63xXYNu4Fzt0xo7kMMaCOammMwCFtBSXmqXdb2t+OZ
wT7j0oEU8zxkwKhqndmq0FysfePDXPRuYz0lM4HmJkHlaVu1W76toMR5d6TamoLZ
Rx3+Vo5IE9Dyav7XOPMb9XqQ9RoYSgMnNz937n0uceB59QHIHoF8l0T1o9H/ee+e
DmJBZcSTAFwvh7mL3beYiWg5UtfET3qbO6TsTc9AxpsD2WbkJ97SUr5alAZz3yXF
/KrLJiNF7Z+5no2Kgj9QEtEukDG5IpyybH8w52TKMN0+f/p7brNkYnUDeA2b7a9/
PxStP7p8sDvhZEHHxwc4Hq1ELYsGy7bo3wueCeSeAB9UPiw5+nVPki0m1crJxHFW
ERVWV41/fTA657Hmc+mcqEbTsCczIftfh4GhmOAfF6wvcaBEs4eTNKNwnP+UPJb4
keDeDnNBmvtRLukeBgRszkz9GSka0d8aM5w0+Nqg9jWTp+GvX9Rtk5ZCF5zV1+Zi
g3KG5PlYHYbsoQ9aD8jA9da2AeBaT0Kpp4P6OsO4dgksLN6UhapO5chBCi6qaAoo
43sLTIBHtoR0+0pM1ALx1XI/NhGsv818zSdkWwuiy/Do/TJB5WtkcHC3VahE2tOj
t+JPxovCu1Uds4SFhU1AzSXcGY9j1dSxdnFUEvNGqffobCAqUz56rG4RBU3ABHnB
/9zKC6dVEb3e94OZ8C4nGjpwHbIHb7MkXOJ6nonM6VljSsaTuSaN+2l0aM5Q9mza
5vest1oOLAGI1DbQmIE7RoURRY2QBxBwR7iD9bUlE02RgBoXoqHLY6+DjnmVmNgL
JuiO/teL1NxEngY67iQDfDOYzjncNq+0a/HLLTC2Fovd+LmeLITRIY8LY8K3KzsS
X94pA5BDod31yajFj0VfXbWZLXsYUfoc07JmUvEs/Hh4c0/tyYQFDZ1n5hBLkJ2m
j5K8R1HKydJpSkkd9EeleO3GHMZPnxOjxXyp0VoFhdRreM7C+HUQ5rYjro2AIzI3
L5zVGAYdJM3qBkYFAhUs0KGDORqOANXN9F/nkPeMdRJ3l/HdAzbwurhF+kjoap+n
iTeNlTxd01gp9007wGnxi1wOWieAlEKeyuwW12e0OltGAdxOCTqWXvMRQQLVwXCY
6U6eG2su9toEIY8DI2BMcPnx2n5QRxgCRE5cuP7egJem19np+M83gs3eNnu9AtJD
SbHkNb03mypqsjsIf0Sv+Ujacv6bMEN9lc85vhuy8LRHR3EWdff4mICHFSa+vN3+
7NsrD+FjY+lwb9n//Kx6jJChVsth3mfFm7/2DIA5noUheFDtIodRg9HVOANHMcJK
TgUZwBDv1AmczDT3lHScROgZJGE4PwlO4ePh8jNBn7sYt9ie4kgW1GT8Jpj5Zp31
gNKqg6EnEgH79BuYejrqYxkWZknEvLTCmNefwbM92cQDOuZiNuKKCJ1EgHXh0lVK
xQg4wk5xI4K6eGn9cdrcQmpkrzr8zPAczu1Ro1etmNd8Ul4WcDdZpakdb3+Uc+Eq
QT0kcQaH4sBG2wsbN+CVvg45O+LR00NSwaAYvRa12fpAMGWiBR9j7c8uxIXRIr7a
Y2MkfpVQ07dQJQHhnY8nhXoa2uKGvNEw59ExNgSg+L8F0QOggg5TEdAomI4opNht
X+XTNPHqz6ETyKFJb8/rTiO2INNZXjqWOdYP+DAGJ9uJ55SDvyWq71szLZcQWAY4
kJW/xjxr00WTnBKDJncE9Cum3FqCXDasS3wgEMDqi2cRWL2YXXtOZJMcTy9cSguq
gCHcRKF3DjFVeT9S+xJXwXw2XUTMTGpUSxhPZ84Lwpw/QoonV7HhJmNTtELugNJK
qAu/F0hgrNp8o1hKPHvT6jfXvYBoLKfZDVUybcExn6kNVIQX3kk07ZG7vu9Jjg7t
F5soiUoTnVhJnSkfHWjV7qTfzSahhbCNAe/yLvNTmHHScXvb09xvMTeQrT4GVg1R
pKd2tUPNWIq86QFfkvsy9lCXkxxHd3GEjxY3vpiNhNPhOb55hZ2brA/6OyRexU3+
g7CWx40ENnAbC9E/i3aOpm6d2U1/bAP6qgVKwdwxLHfGGh/2WBqnQIFk0jc1Cxua
oK2MYkkWhao0WxObpC7sVtgqPtNH2Y9x2nCweNDYZ4+QOuvjboX7PF7wVSKtZDeP
/yJ4hNB1QaULqOG4iGTRur1OTLKODAcW2uHiw62g5fF3nvg3WCILBJ/QkMnFQe/e
2cMiPh3LUSvQRVVvcC+yNxoqQQQ2au457Hil4OV/f1qsryrdI77Xcz5Cnzi0YLwN
8RxUL/GZCLMZl0f0p7dk7CMb9oShUPFKwFg4Iyp2dr3LT/AiZZglaMItfsO/LPn5
BawfM3GffSoCz2XANyDNvaROw749GM07aGJeXakP/gnUyydXJ13q7SHULmumGPBS
xMxeUpye5M0jeYWhJpRtC2S1aTR44xxjOcQLF0xUx1hR0hrmnM4sQZyOCfX1sCzW
+R05E3eFQQTUcjFprtpuXHrdm8xjONw4QnnTUCwpsdfmk/zLxiSXwcW7rte2+7LC
vRjLRmF8Vwb4kSvDF13uTL7slEzvKhaqjAnpIaNd1mbyR0un/3X/QJ8QIfeytVFB
QcdfEeVWqqUFKKZQmBC4R7YRbhbR6o/8FKjWYfIo/cGY1FZhRjGGXj7l8Z9mcCgL
DlyHTrC1sInLAW64CkN7NH02hic9GkUlyl1WvtCFUt/VDsecy6fPYZ6BRcgrHjjA
0c1Uq04lQlWUgdLo690d0Vi6GoteZPn9iC3a/bLlhyggRhDUmjWlJyTCw3/xMLbj
Z0rRbicRR8XzZNbIFEBunBBjl5aKI/Jt45G62a4sozDXz+SntQeJApe8iCp4S+Qd
eya0kHqWVq981IqPNMAVx3fzPjCtMKoN/hocgMGT/pG1PWZm/LfG5xhxA1VBbU6j
9BNZISJvvAdSQS81S0amsaG4dgHCH88YjO0VvLey7fQynuEIq87THcOGfECmfszA
Xocojklrz1KcFTisu/IdeYQ5CZlscIbIBNSL+W2sXIj6xf+xI46fA0zMESBmh2eN
E3IrYqmAYX/rK3WkaBsft/R8Ywt2PdxrdPPtmFCeQO9kbjMx3/m8UAQ+5ru7UnN9
Ed55JfUw81ZEoTavQWhlP7J/CGI4nPxr+ZSaZ3J6hEjMtOqFpiR9ml83QQTnABz7
HOFeS8oykUIIBniMH0dVZPUSMvdnWwE5mjDC1QLWOnDAYcKKEGBazZbqQiqumeA0
2ie4x2x/+ZrVaMzSU5a/3gSQuoQw223KOgOzSZWoa9kMdu6mTmoVa0BS4Gn/7dQ3
QJ7jThRulkaNyMiO9BjxTqmrmBW8mPBYpr3hWDF+yKtmpMIOQLBzbFiFX3MEedWO
WxleVJKpX/XdYxYVH/PyOMZ4QHXN89z7JnIlwzGW/0IhHEIM84LTXHOKvHdji0l/
R9TsMyVvJ8WJV24ipfcW0m1Kds+SuVebEoUBYoDXpOZXvNR7BAYXJ191vnpZSBMY
Jr+7fUhQiRD0VNnOxAgCszLFp8+hHwrXLsfIV5H+tIOwP4eh/M9/VcClEi+jxrH+
SabPXED35OYzMLaFli4tFqErUvU+YpSJZDIr7L4gnL/NMy7n2V1aluXlBjzR3H09
jX+ZwM007XYFa3RCt9jGWnnYvxhaf4B2yvB+FyPrAoxNyPQHFUPrkhpQiuREY/rE
tM6pGqTokj5SNxAR7ukg2pdap33KGIsj+6o296zjR06hmGDWkWiKBiUPOtnBWdO6
M3TBGtV4wfoFmGBd3vUWt5YNSsxGsxsRSnwWmXQ1/qPTz+R85FexXdVhD53aXyC6
vnMp2YDdZPmTOxYF5V+DKEZn9/xUlrVVSbZ8ze3AOlKtU43JVcGSyq4Z+DNRlxLU
pMDPm3GvOsI8Nrim6HsdQyWgmidqyLxDmad1kSxet5FXga0zLEEbXPD6y8UEMGCn
3wR7J1AFpZqtF9otzhD1kG+WR+N0rm2wvBZprBWWshixRgK1QyJrGo0YaPwC3+4Y
UZ6Ky+BW1tamg8M7RMVJhw3R6PjDkPLsWUZcqcme9+yL42a2EINCQ+ZA24BfjYV3
nQliRSIixzM/0dZU53xfxxK1KEZ9aNAp0AFUO2xzmnXpIVCLCxKndQBVDHI3hLUs
tO7zSDztN2YUl15iCojMI9yhNA2LXBc3M5UF0xKQz2tMWvfv9zYfhVHduE9G33l/
g1EWLw1XcdjetUOJYuFDwjEbUDMxqUyH/XrUIMM/19oadfSx/KaxxptdeuX7fXfn
8VYKjOmuKLJ5i4cvZBCYzkBj8oOf2GjbhRSav+LaWd29SxsvCsk7OHOQ+5JsEvRw
aPk6lc7bi2MLq6i5BTCc8fAbUR3AmqQto4JQZZ5wXrtx9UbNFcKghsS/MHTk8yE8
6MQ8DES4hxChITIpTX9Di2fzREP2l3+QK43kV/kKUqZX/7UM1m8eNe7V6d4sH3oY
jdfZMEErN8oixm52LpBLfNXUPn/G9UHplYE8MmeariKHGklqivh8KS9wtE86duHA
sr/hRYU9m07eO+UotPE+e0L+RG7YnfqIMYsfHhDXAm17g+UBfLnzhaot5YHREOeB
t6jn0RIlm0qe8rt5nwac8Va3nX/+GWN0QdIS36k64MLNysw8kKA+Uw64Vl0UeGUe
/e9H6tnLCOfN15rdLQW2x7nyzfYUn0E4O4wYOrx8nu01XBIlR0HVF1cSzCyBPaRN
DjvkJc7UfwwvR6ufwJcH75IpjvCPf0jHEIYkf6iGdPmll325PiM/dtCBQoG5OXe0
GgdLW+ewPcn8ikXJlF6GFunLk+JruBtrLagkDAkSBdeNsv+2jgnN68FPtLvzSrId
0VWCj+XpmhuHi39aV0YdN6gDuVwDnlpBOjqERFMXjGCce4YcNpiEOhjHm28jwVzI
dXJXwCB/LYesQ/DOE4oQVZN9z8jXmr66QxMJZO68AkRL90nbt9l3c/D0jguFhfYj
aFZULcdgBG6iFEj/MXMmvlmb01392L+OrWtII5nib7jJPornwkwqwNanQAyflv/b
VOcydsQ3mEMjQJfwEiJnJlZseL6CN0vz9V8nzAuhU6Fev2R2SgQr1DxpsYGtcRGd
V/cOS9lZEyfwMJdYFNFndImWdwPKvJVJAcPBFUWliA9Z+Um6p/vcN9e8id7q1P7M
fyEzG5v7L2nmPoi8p57V87/DJp4SPR3h2JVzofhnK8AOGBm25lKxmz3buDPavnkt
GFjBIFTrsmIlTROHyjARCM2PlPzAIbi1yH9VCkIWYGfectbhqJN1UiAXnoT1DXCL
TWIM6etj4uvGErQN20uA+TZ5z4rEU/HqbToyy76Z2b2phvDPji9YbqgoXbIXc0XE
KMo1w0NxltoUDvfJe8yOxAPrazDQ9F2zkcOuzSobATZCVIfNpJxwNStoxdruAHEq
98zjrpd9Cu7cenAsEuvOsVDR0V3FW2djsnvq+7Yn8Ugzx3Y42U0jxRHLm8SMO+64
FxbMC9E3qT2NO0H70mqBHBXJjV7Mvhh2J7yzY0Z6y0a1ICgaowtvEpvWGY8DA/aP
IxI9oGBKX+3msnYPfvcmqZiwpILiBYyq/BAB3S5rp/LNcNj3RYqVZ15OwujJM8xk
GYtgrBHcAITrlGmjf9T6TSbe+VeciZ9VQ6IkXDlshPdCbymYQGJKVc0oU1DtgL3M
rdh/ZUH6LfPFgduSbqXorCIAR6H94Ojcj6RRVul7Z8Bj+zR5804RYtQMDYT0fVOT
wJIrYH3l73HuUQQ7wuKR78LuAtgtYEpuL/xCvjkCazMFN1k0ES+lbAcn+I7NsgpX
aOOdGp9LtVB0Gh7GU+h4I5ZTzRBBuGznmTAFCJ5CYE44twDbyLQ1NnYDA4wy0yqr
KWEukW7IICBOfaSh4AxhBwFqF1x30TyfZfCU43b+WHa48BrjXR9eOYnR4hyEVkeW
LJ3XLqPc4fxgF70YarN+OBxOJ+YnbhQxaniK3jF6g6YTM9f+2IRHWFGJ+8n9CygA
XYCLq8bUJPYhAj5Im+Uyu+8GeU+ZTy4wEvPMAgZn8uspwqirLY9oaYK8R2MrBRgb
cnK3vezcC1St+4Ev9cRWSdVQV4DAMOtmjcT+O07ogA6kS8hJjlU5Qy3ttMsQqtXl
53AhlwMju45qoWTbtaptJNvNI5hSHy40jRERyEoR6wabVfbwOlvCR48L0FLm0Rcs
+bHWlNquYY9v0q2FUrbf7bWuYPPwBkyO9riFeYAvt/kydnwnIJVGhzYjHtq95ScQ
W2lA6QIA52cDZzU4QHDPerWCMxU2WAplYukyZsZrWX9nRvYAD9tGSCSQIzwG86ap
EWEwuaKX5CKVgoNJd4/McY6T2SYNAnB0RzqQJ90/8BEoWeedvY59rugEAD4FMMX0
Knyj2HPY7aIFXUk6s8QMIB/BCUSTqHV2u9xmjPYps93idinQ6a6yWJZqXfXOxpFh
pdJWZvQnQGK44moC6o5O7nKqb8P394t7naB+T9g7pJHxFkiEUA7Hy06c9IQuY3hI
pnF1cUsgCKWDKIm0VFWwxo1gZJkviCrLVMrRuaKHHlXXoVYqA3Hdqkg9bUX8BoDv
uGggHV/Xm2+XBX7IiEjJua5YLu2QDXbObUif7BoIpcrineFZhuPnZ3C/cKRDXsC2
Fr/9UbfHwGoxDoMEc4B1NZEQWrUKd0b6Gy/PEVMfnBnX94SAYkoVrzKoZQC9C3tn
hNJi5+nLchc5z/cl6mWUvx9m6KCfrVe2rrUy6jW7Vu9Mol7zENcVyktNbwREVT74
ibOiN92wLkzTo1psAkU0IwyxAwV7Ee4s6qC26zyF2ceIr95zsmVGqfWx6/OVwglA
itOIPTIrixMxVcaPdzaTEFZ/u7KjodXiXPyOLA6OdZ6SEwL0blPEn3ewsuG5oFit
m893S2pQZ5ElMTfhaGDsCUzCHDpfKHXMGECCHVff59tfJxF3LGEoTTm3/9yo/9jl
cX/PDiaGEySbq7Ktc6+tThtWd9TpnR8vfjSa/E1SJm1ZxPnv3Ra0reM1jAs9oIxm
JAg5FIGyNSW1yH2kVgjLsYxJXq0EoGD5DpE24kp0LLnMDtk03Cgpwwz0RC8nML7/
TnFwu1lhzTQWbYxz6hoKZYS68yOdHl/mmTlc9XqWZbkpgRtAF9CXcLMUEr7Uh8I7
jASVQXMMRjU/FI8ZpCMiQOOYkXhFKoyjk+wbjdjR+vAKNyt2884pKrWQbhbo8x4E
F6WX9uSiC9aJzZQFREYiBZKKyHPC+WBPracy2Jd6Vr206PYbtC+364gYERtRAQON
gyyr8eahuIwjhNUw2c6znFbai3oDjnndhAGnrH1gj9Bd6yq5lCdcPF8nsZz0rWAL
/3/dPKwMZ9WfeUizZwUeeIXd8CiuBqpGVyYg0EeNV+nrmBlz64j0dLA+m+Ah6CW5
zaht7wDwoypeaCym2STc+3lcpbSQuqlgKErfDRaL2yqiQy6FkhAcqv51ZwyYwXRv
l7yHL7Rr7nRDnTkOt5Mkwjr5P5p+dQ3mutvEOJT82nNMQVJ7rUjznFV7amYjiX2f
BfwWA1GeOjfOes2puMT2GIHYkfSIlYtiKgskCN155X64a6QCc7qCT0GEZrPWaMUX
1IOA0Qp+eFXNRU2NUGeUX4JuvfC3SY9EwjZm0ea1IldWhLNPnU2YLuu1/fmflFH6
CitRvkgcDryRQmnAxnRwRdmVVoeAEZ9Su4YJGPlu1C501o4CB9LPhB+IHr2lEOlc
C8G3y4IebC+6DSNJPWO+POXaGZxYfxVYsRrEqYLzYsBXqysWbm2biGgD142O6nbo
UbWKaELEhfhoPcjDnURsHqIeFOYb2dQacj6S4lxOAmPI+0uqsQ3QcONZUWhsFGFX
WcDW2fmGUFv6oNRXFWHP7NoIYHZC+e+UVAkWQDvGrEeiYf8szccLB7Zt5VV99M51
atqmHqwxeiTr+K6Ek+cZUWMskhj75ovn4JS/svIX/OPf3kl0xqsCw+fd4M4Rphnz
XfRevM61gyJ3Ty6aUSITNgwupgSV9uo4R6dvKvqwS9R4MZz0kOIF3oIXRG1BcgbI
miMZD4CTAMRVUh+lK1jh7btqrOCYlZQg2g0TnMpR4kgzXDdTWWtLPLlGn213zF1c
uUHamjJyeRMR6dPIS9OWado/PIaaFNDUv9E4oY2M2yY9Cf9bC74o8psfbUF/RNkS
seIVB+iMTt8a4XX0JQo4YA+bwb7q7cXS+n0U+A8xRNk+UHmVZwLPbQgV4NmL7biL
A8renIAn/GxHqJf2PL98TlQ8X0fkxayeHLqydLDR2lpfse7KEIt7aEI25xiJjuHU
C3qRurdH1b9qGgPdGpTIUd2Tjbh8GI8+FwOQ442F6hQQbGbLGazy8IgVqtJJFbPO
N6GVSXZC1iIzQ+KjX8vk87yH5tTKi9oE55bPZaCLpcJQ+1HY9KDVGM2IgYv1RZgz
PrI7UYM6cBveYwxCMK1tL+1N1WxZ7f/E6oEhv39P3LxZTEIjcuSaPI8clxZs//Xd
uhB2qUIbcPGG6kg7ET7LK/nSs1smHlsBHqktAJIGRlBEr38fD7VPtq5xQHQLyKwS
bwlWyy11+dGlWOyJ41d7fv9of1xhzr7nSKDd9Kp8+DKoSVyJ26joli3iGMIliI6F
4KBlYJAUGVQBKa9j499AdUcHS3IHX8fVgTBj9HjGawWk3LdiqiBouV6umPEmKY42
LYX2G0KMlnusWVv0LNEWMaQG3KzfPEK+U40FNvIeeMSET/X8b4u2zZLV1F5HcNtd
mMczQWmIkLusrEgaJcQEWs+dDn2dEJaFMEiv5L1cJjtam/xz64FK3vf9tAXEVNDm
Pmn0Pv74D/Tc5nfcUhYR0qbYF8Y66KXh9BLf0DszqWr2rLGbKECMBGYiUPJp97u6
PJNsc+MMkUGkrPDu72uVRLGkc7HdRzWBUI5GUiUxLr/3sMMDxh1HBLV9sPkz75QP
GpLIOTcTUTc4TJHLEkq0WNkpeFJT2BJ+D2dIEzQy9Q65ecNv0GUacPxWHTBifpze
PdhqJux2Cb3ElfZqwGxE7HNWc56v1ow2f45cZQ5ZAioyNeCyxwG80eKKd4UffUK8
3t8OK71ntjOJCnD825UwVRgAbVnciCxgEcYvMld7QqLHD2ZUpU/MTiMt0W94OLnS
yycUH9xiriZJ+gQLj1f8Jab0150s9HCooZJIB8fdMXZuSgC3oiVH/iSZFhisLmvo
COA9vyBqsUGdeMbaDYWf5tuu3WJ1doup38ao7yTZyreqEAB/d4qc+aeK110pgWcd
Vi+HgdxBu3nuLqw2pJduo977O/Oql5L638JSKMS0PbTpN02DhntsUZjXo2VBeLkY
qL5BWtg2RW2RE8W4xRdHNjheSbPR453t1+puSqCwcyzesy46dUThzK2+oNdnQF+z
xEwTS9Z0qZmbhxI2XrOMTfTn5+NeTw+uP7infUpGTpszzv5QIUxt4rrFXiuQoLEl
pdL0QvcuRxH2Pkz69z7L8cFSr5BFfHIAk/546vhOFJwMbEUEU40YcjosMx5JqrJu
Y3ZTGig1fRsDvn+uIJES4C8sYrI20haSLNOc+PlyIDsAX3SjxmAQjhPZ2bchfGNX
QnVwS0jXO/sNIvWOCs1GHfc03sKB2GZwoLs4lR/oMue8OBCBEYpmEVl6AQn09oB3
+ChyDFu7IukmWDSSVEljyuKR3eTR+G3exInswrz0xEajno8/SWl4bgcuBV/dvklo
kJeqNM8Un9bjdTXFZ6Pynrsr02ijGRkK4sfbG0FklVr4fTb3MGNVx80qhfEKhMBh
SdbK6icUfgzsxUohqm4Q9FNT62nlGS7pVyKlAjvEOIZCVEJLhYHafNcTyA+fovjq
1ItUVXqx73RzggwrrDDoXMeDUPPODgR9qJpOn5zz9ETzwsVN/XB+xU0plA+Sw55I
H+Rc2s8H+ewXRkhbZydbTg5cJwBHIy5N6D0TIPMVs6Fo3hklCo832aOc9DgYUOwa
dcXIS8EzVu/HaSZfM6B0HRaFV8AbvRwbjcsGSTEfF+niHdum50NduXjeeYZWSekB
dCOrRti4gTGLZ7EWAq4fcAnaMI+yun5EvlbgS8Txfoibq+Yx2MKrtUu9yvoBDal9
cIh1Je5i36Q3KCI8K+0u/65ARmcK67Wnydojv3SoCXw6GqPiRgMUbz/H08JGjKkI
xDk3JqhOGwzLz7YAo2IZWybrgobCJHH9x6jN1jTvhBSerdB8FpQ+lbcpsOihHab8
vvLXi0qz41+Sg+msVAMwzy4UysjSxeE0IOsASJMjWKJ98Gs/j8zGIcJpIMtkZUJm
MnBSUj9JyGNKXGwAvO6SOgIf4zcJBR7YgQhVpkVGHUuC1sVDoliZ46l2EhFFU82u
CrMPoN7+q74E5roFCwQH5A40ShY8xaklow46qPLKyHPPmsz+TiN/6lU6kstowiXC
PNo5/gBSYiPEcooXWSS/1JojczlnDxdj+SuvFE/p4LI5z8MlMFx0+6WzZ2YPmRVb
pK1Obolvnub2jdVG1n24f170LBb/u/fcXvt58BDE1uLIMAEj/ol91ywHB7MkrW1o
PLTXkuS5O4V/VF6P4/atoCiXBnr9rc0eGUXPlIRv5WYh00vvNLmgmPzxqyd26Qbu
v0kv6CqtJUBOU7L654kSmNPNkFqv42jcw1WSEqQ+izrI1FhbNa8Z+C3gkYdhD/HG
B3VMqu7k4HtjwLQzj1hPOJ9lcIZKvrkjyIzzEdB9eHJCIKbzH5fRLWvVR7NQuYZ7
8Tk5pus2IRMB9Mv6fqXE5Zpcrd+UjQMBbopRrvyqYPyugyT4R6VYtoOC0TkTgd9j
dOWyPnDNehzASqvEGD2NSVPJ8mq4NxUNBW9R/rsypbQjxAnbUdO31dJOAh9bzT9q
+8xJCsn37T3znSCg/iZx+mDc6gTQIE0BwOp3yD7MhuUdzOqmY5nRMfUq5INZmGAi
HnKJJO8qznkfhXJngiHDYV+M6FT+h7l92f5970IwFj6YDkzAOoTI58sn1kwxj0dJ
Ez/eD6jUyIZn+NTkCM6lWJQGRt5SUj2UkdXBL3yFWbVG7693uRChGQ8O8HvhEKt6
CvzLRmoigncQJZNCZio4hH+PuFH4rhFAPT0hmiZxBSqG/ysoe1ZxD/blchKE7yci
1m7daJ0qrZz2RtDpZOtn7WalD2j372fyQrpvXEm0HpWUl0dZF8A5nuyWagV8pBd6
Zf8IzXUcuCTd7BKtFXBgiG62+ZGJjhPN5A+0sPYyleu9zwu1a+6QD9jxGQ3A0zYp
KNwhwWbeWTkkH1O6W+xh9WmoMB47qFRl+l6rQX6DoDFWgKHqZVjxIDxsbIaoyBxX
8H+h4aKH3TySR5mVxqyZM5etJ/kr/hE00lg7D4OOA4tQ8O9C9AE7sslOHtw6EA3A
f65m59sAUww1YSHLGHi9Z1RlzM9ByhaCT5fk6xML8Fs+sNUMjq7cyhXcnXzpVBlw
d/gMEhPqretRxzjrW0W+u0eWf9b3mfGN53YzRMGOElB1N4qa9UIDlrE06ZCpRWcQ
sqG8u5JLyv09azBUkOBenflwjfhm3+IZbylwLq7noslJzp7PLKYKmA3I7VbAl2l+
nfuMv4J4XAOWm/pqS2XVKfGOp+4MtbonOndf8P8SeM2IeXhycAxgP+GUDuvdn9MR
AZpNVTmIgtOHXXuHhhWwKe+n+GS0R0flZ9mUAu0aW+RJwtGC4mJH7IkVrW5I0jaL
k9pGJoBFQZcu/eP4u8K8qiB05PBkB6K0lSgksRBl9cKGyjCWW97SUuaVjADpDO6q
9y1938FJ7G/fwKcl+kYPwKPb1YhF23lmJLL5zSNQTI2NpvlMDE3+dA2nOD3HHnOC
uPrmR8YdNyIRWDnj4GUx8TB+hQLLppFQGkghkO98WIZegwCmTs5yFoJ1DusgOzIK
bm0W646MnC2nGNK/Y70JNAMJUtK7/NuiUzHV3tnkeLvevPHnfLxa1M/vyxrSoUeh
G0jP4wj+NLRemS9YI561lJXlesYLhleM1bSPi3avoVzhBJAWSTyEXln67LAhiMmK
Fj2rq3SINx6hHDIbgxNvMFR1Q3eN8flpGU1laZ8SEMP/hcq+DvNWPcpbat9noD98
NNvKLfDSRaKdVXaqKLp3VpcoEC6+aQ9pUyH5mVtzTElJk45HA7eIO04TbPKOq4Te
XjyDeu4+e3hnoeLZP32rnX7Em+57Hi8YRGxAVCHH85xA/I/Yxbtm3EzJyun1cYHi
uBoCLXuiwu4IueC/7o1EpYCuEpZnDUB6BU0kYFm2pNbDdTb83WuIwSYqY+1pSA81
JJQnw3LzzmKuqlb5guKsoOxqrv+rLAy+raMd4EN9I8/LOlBvrUCakWAXnR57xzzG
tCXyoFi2Sp9H59kj0FZA+i75XkkZfMOtAapzunKYEVeVuC2cShrrLBORx49NZ3+5
gezMkC+eiy77bzJkpF/qF8zq8SFvccEanLgKVaww22LcqTBClInSiFgBYX8/8H//
DIwvUnCsgp/bFwx7Xc0gDzbposoqyPc7BYZzmECIQXHMD0EWoA31JarFRtWsthc9
vkRf7X9aVYun83DHs5oDBiJRI94xcZw+kB/EhWdc3r0gwwW3soh0Jdpa3O/DqqSx
gvU8MDZLVv/cvtaZmXE91FHuEhdyZvwSyEqL22YZoQcc3BLQl3O5chbS0SEN/zVV
WNqL200GAFFryZSkdC6RpD+9OOPYBijNZtLYTdjuACr9GUu/FFVB3SrNh4v+/5rk
fQ8NFO8wNvknv8ofwG33pXyCGRM2Q+DGnRt2dMoGGGouAifqBsvfRpGU8kJ0X5mC
aQgp5WPjWwXsFZxAv7ZS/N+XcyHLKfhZ0Da4YvrTgYfJ7BQ0MSk7n1AncfXQzlIz
WdTLpdjii+1qJLGWmSLPeMjqqpwgbmHee//yGWItAjT2qpiorySsabUShV8sJk9c
cHQnqhIVbokzTyU8ZwYjCeDKFV3EjfW8R1PXbpjwOhcSYob27D+YS6ykyLUSI6w4
yUnzyjMYsQQOGCegXVWuyr3ZHSiV3S/yYAkvK+G8Cf42RwRGaPQWBRRA/qsAZC3c
eEyDA3nIwYM5DRSS1fBOKyIr7NWzYSiVJZyQrRsNiFhPR9/y/Hcpta2wKr/J1xBo
X4wW9IBz373LEbZp/mHK3vrIvaeHa47y6Tj5ZiDDu1n0/ShBugNIMk4NfsdsBZa4
94BWH92hs0kiMb3cpG66J6ZZozHsYSavoXlJr5quwkjFmA7WVhSEN2okz+6S5Qsv
4Ptb4NBcjQCTpTLRwzeWLFEekMXI26d9Cr3GdFMf1qNwxkZwPcw5z1DVfqcNDNU+
gGOmkrZy9UGPycRt5q7DMHYX1ftnUia+WVs3rv1uKzHu1AHAJYBeOMB2QdKnEWB3
GeE91SadK76Zx9OV69XDwb5jx2UhOfUDKuCpGVNGS7NNx39lkt8HUkgQ8hQtm/DV
FyAmUkP4Zlqs2vtUbUF216lSG06HS3ox0VTZzFJZGXQDidHeI112HyRQ6eK2tuQ3
WV4RRQM+sw9RCr7AmgU8JAgfXdefFT/NuDySecMr7HHLgPZxJJ8ZjSPWvEFsRiFc
/yjvc/CzNLKiFK3kmirTwBYaEWowQOfGjIsEn+zug7WlikTTIFwSouvqb+MGKZkr
BUoWKeLKimEa0zO6zO0J6BFHgb3sjwXAWYeUzQ7Vx+b3UME2nb2LNK35dX7zcG2W
NaOhU5SHC63SS9T5F3cBkUKIs2l70Rw5yzh84GYhXw4SAB+6zRIr+7QuS+lnx+2F
r61dKV65BtMao8wDXyifXcf4K3AndfoePETgH4RX7RVdGeoXGnGW16cKEH60Xz+x
v5lK7Wb1fOrAl1t+1KOlZ+nebAxYdvCaKtFv5er30rClb4JVo2SiZR1YnxneyXy6
+35b/UJUCApRbrFsV75fyKPpXemzwam6qRqk0JFdAzzNWPOkylEFAulXV7T8G9Se
HSS2dNSz5nRUsgJqWDwP/v/SHvDY9vlYvvv6FmcpjTyRWre4EHEPFLQIIQ3MsYOT
Ji7ybZ/7CBxmNvQP4hwDsucwHI1ztAwYWcLhKZ753OtdpH349cQRKri+oPovvMx+
HuxsZxhDHcpXm/pkcaRRd1Y/LDurbAEeiPbEhrJ8BGtIZrkiD5EdZzEvqQZlpnw4
+iZkqy+12ZCflfcj3DyLhxDIvlimwV9hDsbHeXur03gxoM3k2YFFgTU/m7HQi3sR
xdVPOMKPrMwQDddVism/lXaYMPwTf+d0Rm4JAGentbu4+CU7d/QzNmWLLT/lZwHK
CaV6PHAbjJbiuxxrIVW+XzFhomEFPrHD8O/UcN1pc6aunpEL265r0VJyhuC5BQgb
HjP2Mr8WduUSvwgan2c9fFtO+r0Aw38JiSWrHNZwH5C4nPjwRjsR6jEU80foRkAi
ES6QrNrM3zMkpI6LMVBms4kQWbyFOzWQS92dQvYjgyI9oruSmpgssLhhRPCll4pM
3g/tHwp55nBoi/b+Z11x4rgfMmU3rhRvxgQwK8WDvID2KMRMxoYeJPodBbiNp5iP
YyC6iegOXDDPQrevVnU0rNdp9tp+/nIgogFfnUkoOXu+kok735/LEN2QpDa5AeXJ
k+5pcteXSjltH9wWf/mt0A9vawrmDV/oIC24821lznJN2/8yAXSp06AyReBnztF4
SmlUclcu9Ga1tpng31x68tSdd+ZHdNfSbdF3USxZLeXl7c4SrZ6jc+o2Ju1ZF1y8
PYT+s7DAfy3Mw4wAh7Hubtjb+Xr+fRiO3X0fGai1TwPrVlz9X6xE9vuGyq778y1i
PPU0T9syUiTd73Tv8KA7196n2zcWeRNfPsjnD/QVkFZSweJ6H6GzTZVPGR8Qn/Oo
xNWbjMizS3S9N1eORnb9T9VzEcm2+uf6TwrdfUWC6MKw2SgSm7PVvydTSjXqd5Tv
UnPP9ut48ILsLTucKwDzGTqWMV1PRN6jka34ocJU0XVfxYjeXyWZPpZLpmPjJFV6
WdPtUZ9/ap/mcu3/fs56PG8AwIx32ViiYFQ57DvtQMqUPKperg0kRWTuHc/FajF1
n+QIoVDghVnyK9PjFOSWyxymR0AoJTiQg9yK7B+QNN035lXzogLU2hiJp2SDAGl1
jbXHXzm7upGsNhzsWu6VPM0gtfL3KBYpMB9P2pBk4XfhXDkJWOlu4tiudI+jZphY
9w1eh8GoJmarNdmDzFYkjV8OT0mEy9BJgY/D6/fLZXimdCTpG1juruVp/UzRn5D7
5SI/EnwT76bgFscFtTsOpkxg6YM3yDa4DErjImKNJnENbPr8iE5/wE5HVUHsdQqm
GWT25cRNUHAXar4ED23ClwizLaM3KK/s84cdcLR0Xv1b4LTaLJvav9aU1QbItuij
BDoY2R7e17DmUF/WA9NogoGJY/eE9IrUwQuYHC1Ufs2HwDHlz9tt3vlexrLuuQKR
0zmPn7JDZ2GSnuMMSWJ0aZeDk+YAk4yHrxXTWa/T/s4h022bQKez6T35CMhHJdG3
w3Wnqc8UbIDjLiYmV2ugdT2x6JbTpVlGarjC3ZU12Rs2qbJ8VyVEBe/LLjBntLMF
mxo5BsrA5z9UbgIMVdw013l0GMipGwEDZwKom60hj4D+A4xJhJ6U40UaYq+2Ua7P
EYnMsFT5hVBV75+FIdMLhFT1lYXTd8oa1zqO8PS+a8wQMown3nKia0GGGAT2kRZq
V7Zeyon+GtJyxsNtmlfmSzr2G34i1DOVK3jd8BZHik16ogTG436N8e6zeidDqXYC
32cKpD9FkNl6vDnUFJfNQ05+WRN/xf7qFs8WtKC+CugqnJolxZ8oORby0sh0v4Dc
/UIGVWtFxZE5cqhDGx93dHSFo/+9MMYYbtR1m9IO1v0qq2UE7BsjqX/86mbAtjCo
622qoVZBfu2lkcaOu2QPT1kL/niQnBqqCKrPXMsf57NfaTQ0sAWdeuoYaGqyMVzm
DL5fAJdGoWG9MlyN5b2mS9IldJ9mYc8O1fgl2wx7J6b7fP5QEJeHEeOFH0L8AIgM
fjWLXk562aGO3wjECPb7zt06R04PNR6lR24zKJO/8af+MtZCrToNK5zCFpGg/9dD
5DBqXaEBgfBCMdDBkWCyLapmn4dO7h/IcrUb3vHmELPmJIRUT7EOLgYNY2Rm40iq
5KCtzkaP7+bnrSdNK3kyMy5+E/sE7J3Y5kTmIYG4dW4QNm2zdsfba9iR1eaHSNKc
iVBWslP36rxLCEBpN6CE5iNvSfOBAR+UhExFsd4KBZVSbIhLGV12uG83kR20xE4l
OpmbOUxFqCowD4GdwivH9WReP4O96Xd81FM+ULTXiWroV//8l8HWAEMh9D0TsaTg
KBS+7MAxFpvjB0slEIyJU6MyaXe3FGYUm0KX2gX5sPknyxYZziwhMNtHcW2J260d
9hZoQseuZTNhAZTHLfCwGXQz6diP0OjgQdK2cIl4dx/yFntxwwakAbhOLMCwJkwb
eMtWyjsfp8VN9w3ldt8YsHs1vJgOQqwKkJhxiY2UhHlLiLGFeS8l7s26+/TlbzKG
mdYEXpQ4L5Bb0/Rrn0kp2ospUGWxp+jYPhcx+W82uJGYYqHf6e7zdcoMGrrt8P8o
SZKE85jsW3VYvxH+mCr/yZo6fTAx6JJDy3Gl66eKRh3ISbu4EF0wJgHmfmDkFV5c
R7Iqjg1R5Eoc+NO3Tb4GnFsAzVXJwpZhu46CeR1+pp67AERVyrE/iPY5dPQoiUPj
LbCthBqhsE1S7r5nt/uBOXto3cXjjrPnCrGmekBBcdy3X9HtImuG0FlWnV5LNddf
5XSI6VxNdOySwYLmgMFzC8s+srsjwClsThyK7fpO3sGo+ELt3Q/Fi54d0xkXgJ/+
JE/L4Aino/R9Ej3EALGMOzYK2J/xgO2NM3KrM7LlTiev4cUyw9c52yMGGwYyhjbM
G5OCLczNANSmDY39opkYzMQ2hGt6VcFKULlzhW7wKCAGdqOVW/8ur5HLTdc2VPR3
Jl9zp9l0+0HzCBgY1QYFxsmWWgpbhGzvNel7ioxMaPgv7Y7PWKH/4xDP1fMem/aI
Ij1qNqikVJZ7eigC3rGcRrsFBbVR3f6f4e8Qb0Gx81Yti+pBINZxbYZIBiVY+EKV
CAgAD78RNn15ytDk4yAvcL87j1xufqFXhOD1z9OgqCwfxeS4k5PVcTx7pyD4ML3h
Uk9oJBsgtfyY0Smtw4dcnVzY4BbppjdYqrzcdVXKl4maVpkzqJ+jKXusWvc0vVdF
N3x1ocxo7YJPuPs64LIt7WaVqoAsOwhcrvHRycAw8wXfxJgXv7sXOAmS1mPWfZcX
w8dJSGwjkq1c5O8CHYGMdgTTRIY90fPwTPbKii/64PE2WjPKSUZ6Kq78dJbT0b9i
bXc4L39xa7ias5XOpzvGLKfYwnNlVqdA9l9+hOcL3GyIYmLlf7FecfLlxbf56idj
2aFqlxmtyskJYjYf9J1KZ66OeKTHzS9nAEJmrCFsEUTR9HrsAUFUVZD7kHTow+Tb
/IbR7kZdfe1cguAlyn8AYsXGn/NKC2nWP29NrQ6fVdMYH/9a3BHU84k9Skm1yOwO
G2M4pqnokg/99/d1Muo3TL1W73RXQbIY/2KsRciNqMaKKaae2gfbAw+2sKLmv6kC
+7Qyruq2z9yQi0gw3Bg7Zdcb7YK/EeZzw9nw5Mo+9tsZcnz7QRwPEOG0XA40eniT
GAUB2uEG5d4nJaNEMxCUTqt1ujoE0NFQskjhMzSUI+X35TYxiPeFXRbOW+z56qAA
+hA82gdLs1owtkaL7Gvhwf09ucciiit4hla7GKdumLcEjCMQPBFTXx4IA7nyh6pB
vj1tAYhFGxxZpCiHWn9pnnWKUPX75h92EcfJCP+SrEs0ddCRmyC4gUSC4E4pu8jY
eqPrB2DvO+FOinnLKBYb8Ubz2lJSIK8O/oUYyMugI/jbJ006/7ALRbp4hHhkvK9W
xtBWU21aemotcTIBPSMVWMTm9FRjW4Lsp2MduvCZao8XawSV1qjBr0uvGc8vp3d2
sC+W/oli2BiMh3bsigCXVlNVJC94S7AVvGc+SnzVjhoM/pQWGerzn46OKACIlIQd
wz5zAy+lg6b6CycqFa2xGASrvP4CA+ic5nw1rmxRHb04tSgTCm4n9z1h9uOaywHk
KMPdqlDdeNAC8Z36nh83p8E4HSLSEdOt2JkgXsX3kYfu8Kkp1Fk4pNXOEim8f/ks
H5bwT5kvzIR9eXfFQo7ssaJyAZresWYCFUdpWYz2bDl1crBK8/GfrNqT2gRcCDdM
MJdmuZG1eUC/+69TFxPpK6EMMxljNciXFfhRZ0jCTmkNgJIfk3LfesEdejjc6edC
XMbudk2reNEtu6e3XdwrqZXLjE+ymwFzhj2sbX5UV9+ZC8eGTmeYWnyDdp+I+LwN
tdBetyY0vwDYXrfPBq4FlwqKy8xLEQO3LDBX5fmTA13nIy1pvOR0a2U08uCvTrN5
ayGPuCEJxQ11+KJ0hjgDznd7DYRQ84OUU/uAwH9QpkvDEov+uVukClPXoxzlgiIz
1+zOijrfg+pq1MTr1h9VXFil5j+fx8HlVUcxR0+8yvd9zpRnUsF2yagfvuvodn9U
YWyXzZqAyt0SyCBCGsbeWOc7vAvp11nJqfKeK97a0Fl7W/PdvHh+QszUEmKoEuvu
VvTa3Ns7Ajvl0x6+YaQRVWqsFKbebDR5+CRB6kRcwDYSADU25PeggphElNkBm3rp
Tc7JC25kfm2EwAKaRs28iB53WGlWdJxDkJin7RWs8MMAJr8qaumL09Bm311pxOT2
M+Jhg+uO9hJs3stlMuGatFWzyvvvW53f79nTo9VSC/bUoE/JAWcRpatEo/bd2ILF
erLcdly3K8eqScCZeUU8I2HN8GrlO8bM5zO/sfwRZMhwhKegjPMa2tAN+oG+0TNz
F037CqPTdV5pGCwHqoPjTjDIUPWRPvvJMNK++h+Cv4+LkxburXvsp93wpUeKzQY4
dwmvM5X7MkauJuZzwuhasGM6JLvq9X5GDOLMWCVD0IgN++f1vuzzWTqBhox0Z/E2
TtnhOHSM7VEDNMOSmTh5OVX7+0kg65Xwd/KbvzijNfmNHqPTT16bXZ7UAtOdHvfE
FUEBYryjfz2mMQdZHH9AuOmlPTWHDc1DZx2FDKGHefQbQ0Fqpo7rgm+Ldvblekn8
Fs+XHypZxD8yCUAW8jPbt3gR8Ao6U5SzevtAZpUVkjolCl2gQNx12ySbz2dRJ+9q
FRx0dMwUc/A8DK3EkzKJJCBT/e8yRGQoqPu0pOjrb2py6h8QRxHgdEnH2klDOz34
ijn0eTJEzJwXLEG0XJi/GhDs/PCSDZLAp2eyhRC+S/1mhFY5AmlcYtPzzVH48y2B
vQuICZo6TOqDuAi4PZOlW51YsV5MPAI+2iqC0ixckyzVuEH8L5bh3P/3im3rhfyR
i6MEvbH3gWzJqtHHYqenpgRQjS0eWFoB7I2YNk4F7zthD/sO26mMZBbgIMFyKfxq
Yf4UNM/O2tV8iTDsvYIZnp2krG7GFPodVlrEr4xoOkOlbmtV5TgwiL4nPeI5H6Gi
WmFKmp1PNasR/+YfwY1U9EtBJH4f5Bu+Cx8CbQScxZCqF8ZpCXMZZuzaXY2U1eSu
Ix0RE1VExkkunl7xJubndmTePBxlahHP+FLY8O/vK3xjxFytNw3cyg9UZRjM8vbf
J/U3bEQcDp0NPVlz4427bAah/bNR3OlV4JgcFn5P+pvDvngHt6DOtQrM1hrbeeif
hVTDDK+X3/1Fre0ALWrnhLPv7VbGD3Zvn5gihiuatcd/HPhIr62MB2enIGoQqBSf
HsN63p6CZatIPpnLXUZIvq2acJr5RceKYlaTw390SdtKUSbH0njpGw7qOzqknNVA
f1Vt66nXjqqUCaBOrFKZAzCGz0sS814WrzFZueAYyrCjbNh9hO94vPS5tCvpLvGn
pBxF/z7zDldIKvwLvjfJsvrAJ7Y0acPudHEh5yeLbBdN9cTBf8YDvj5fbcQWyPFx
PjDmUay16ITfDlg7CL70sEnaljTH/1AaoI7y4/9NGIFnNAh5FDaawGpUarSzd2Sh
cXbiQp3C2ckWh48M2+lUeqPQcnWIelr5PwafMAr0OZVtTSs/6Ov/2hTBQUtT0TWJ
f2660nDgnaY6ubbEwfLV6mxGLcpUuv4bQbND6qyjJRY5bxFx4axNPEQwB2GgsDpE
ND5rvGXPz+7uYOdRLtdMNL+b7zTBTqb39s+ra/nLbBP/onWmUWZ7D36AYW/UiSdC
i2cbPQhvAjwE1LOu1vJ7jQIMNqwfsw2JELTWB3uxuUQT5kRHnvsLVjwhklD+gQjm
ZfCVkzGQyxSIA4Upp0RxM5pwOdStSCE2BbROitTdmaVxBb3esttvh5xq4jzfPdM6
Y2daoCgx0mneElKGlp/Lbr0/0b3VKj1SDkQsQk8qMNmxiTcx5KKCWyMOJUdnvoV3
+h5jl3Izt+1CZZpFiIPgteUlLu4S2YtWs2MdVhuVwT8mZ6sS6Y+E7r6JqxEgMOuU
pDXI3DfTqTCmee1H3WxntW2oHSGL0uhg1WB8nA+ESQc/ZxEaWJcrB7jcMDdFLold
yIfv8TkyovO4P7IYJJ6d+UYVleU5Kk1fHXHSPyBy9sZ9XNFY7KLm4ah3r/4+0z/3
KqtOFgbUTMhnzftTZPir3Uv2hv9Uh9AtdFTHK3VCBWKmJT1WOg3ClZAfmAS0U/Ru
ityxdk0Mxwr3V2uZ2NhZ3owhRg5FFhUXYSzeWioY17qwqw76aTD0uW20Mt8lz+3/
NtQAef4AngGV+IElturQT7EmCsV71iy+uT4bQpOjOD2I+PtYCx8sJ6OwUu21UADZ
zw2WQknUkjiFqlLSmybmyX+h43T19aTYEllKMr/11nnO+pQE+j77W9PYlO0iU2ZS
n6BGZd4MhYmrLGVUTAFF6H0fAawslzYGd1XXA6ha8HtIcfgmyctFFfV5PUqxhc4M
aRs0XqlLL68G9nWTeePkvllMX9GCNertXyjsLjYkHUq7hPBRu4T7m+YptNHs4KP8
2nBX5BBZEEirRYQQFx+F1JMVE2JxLB+OreZiRZ8RMC0lLR34S/PmCtfz0OBZQB5+
PKazMatg/nU6YfQZpUlqGpuZH8Cj2cmjPQfQjgpGOOzc+xsxM/INe6j8hS9/VKKg
hBktPaDEXGAxZAUNMiBHmmmO0Qxp2pMjuc1TuH0AMOlizkVV0pfbQEcgwsKTYOtN
Ek9+hffeYo8TWKd5BCTVy3xvYJy8o0uAVroHXC1TdTZykoysQgeEVrjHZqVn69xF
nxET15ml/8vPvWNgeyg3moj7MafTi/mTxsCeM/q06eTzlw4Ia+gufqJVXrj/vljx
YqZZN8iNS8Qx8X9YsVlk3VPyAAWwANpjs0edAUG80gZYHdKvLAGGy3r4wAkSxfcj
jvLF61769DHW3boczA+8411TLNqkR3BUPGoqxGsumXJQxs1N5YQ4C0vU2AJFb3ps
J4c7UrbM9RIQODub4ZYoOqZeIae4AoaOr4W4aH4xX4fM8/t05WQzDK9PkOd99mcz
kkRSA7EoAV88YwmkS+NXWAnJ+h4hPH1j3Zaz9DKllhiI6hzrTQGoRl5qtrI6c1jb
IUsM6jUfwj00L2UyZcH1QSbc9AbWV5Rkq9EpHxNnlLuvRJm/prAqmglsSX3lDkNJ
IHNU9WaHxwTcMIDsSbY5TEbHysKYe8jkJM1p2UVPpDajsiOqN/XzEm9os86GTL+k
jLz0bgOw3rcjRvh3gtMNrGHXNI6YzeSIQlNWwUNG/9JFy+miU1cryk/MHV38BlFm
pCoXajHWuqzFYBdCo1CVfYpQbdynqIDWUYVcKwPewEzkRt25pfaJG8FtJ/Ff2jYi
/8WqBDWYR2gW4QpBZStvTVFDQHwe3or6OmMRMiQnxKoSArfe/uXJzBczETAZvI4f
MrO1JeKp9WvlZ4wZKzV4TP5p/l42Pd8akzOAiW6bKRXG9BwUC8DMlJ2pykISqhtt
BWI+ED+LJVtNyap/4eBjXajHvf9c5HQQxLNElsxQGeP3WZssfDVr9RQI01eK4jdA
/YCP2Ni0GT1S2xhoV0E2b65Nx31iocbWUw+ZE3CRIsPO8DOCZ9mJRq3BqKDpgNGl
wF7MCvKTlFWA04w2XDq6dnteJa1O5jeiCHQhIVE7jgfU3CSfc3RtmmbhxpiiMVoe
818H9apOt8xnNJpVjBXqt5MaCz/oHsBXeUXfZFTncfWJ2tbAYZVfXeOuc4LGEH4L
aZ9/KcXSGJRQT4SZhxYq2YlmbZkgSJbzEbXLB5X/MyC2ZAoOoSS55RGq8v360OnI
+UACsFWPAFo07V/K9+1B/rWquQ1VH3UQAptO1UTh+58YsI+9RyPPrUbwZIWaGZfu
KX9QAREEfuFNUQqcW3smhRToCdnJpsnx2pIc9TvNuVIZtCsT973YsnQbmYdUe8/g
sPqUoW6n8ocK5m4IK1yfpxNhWQ1T02JiRoVrNnn7OKYZRGKETcHwHLGjmhHdztgx
o8EV5cpZ3Ul4GBj463NLsqbNBG+bARUsSI/hZ4wz0AhHP2LA38e7h2AT6YfHfNRZ
SUmVdBtL4S6s4bJOsTg+6UlNXEfeGW9urR2nuzdyW4x/aYcmtMQCr83WAKiZtwEY
a/rRrSs8bEiDuWezlxCFEUCI17njw7VBIc1D4mQSgLVN1nTfTy1UTFfvczxQFhLS
MNauOMurXGzAyh4b3dv/sNRgn8t9cAL2Jykph27NKwwy4qxbzAm/yMiOV1MM8w41
6u/86sxR3ALjyGRcwXkGcKKziygA8tq6Mdlq3riNh8KeQiPo+H5jWOCUo+rZoARr
CP5tqAarWR5GZ2j/53doOv9FBaOdABWlJ5JdZNmjiNbKiSVp1viH8gCnHFu+d5eK
BhwlGJcvzDXcrP0xIO4a/6aKuowXr1hAt6NbN0Nh9iaKzfqCq3RXhqt0DIyYp5Kt
vr2pi/pydxNH+6XQtPMyUZ5Xc/vle2luiQNQ4BX4DQ91wNYFOSLxbjrd9qXqNOd0
DrUlIoOKrXU21yCc0ws8zqhJ7yvk+h4lZRSsDLGs3/GIvckf+w4ubg/KAvDQfWCr
PAhLMl03uOeIVi6HzKjjPqCJ4h3MQNa82uDabd5+koWblT8WU2Rz+77K0ZyEmron
pY3QpxsZGoXisDtYSSE6zJD4FSRyvUjuMnId+s/+fj/IIFCLTAXhTLkLcd7zhMG3
A69hvPUJkdT6c8My3n9rfOeGNmDuOX/vchud0lebHZusq2D+Hhc/8Kj/pEOw/Nej
IJw44aJ6QW1N2M3qb0g1TPhI+P05dp/pSNmSP9CwRgi0LX7B6Wa/WX2lhGkU2z0P
5mKw6M3i2lDsDNLexsGPXTZl5cyGv66jk67SEaplmdtS6k4/QJCVDtZfEj4SewcD
Zkk8eL0lI9qgacifv1lb75VdyobulkPjTZNZmSLler1yr56we8C7VZcWSLvGLiEX
QauwLTttb0qg96E0u7Rx7jN9Y222NkF2DTdVSE0o0c4hRjnzq9Rogky2Ignf7SlU
fXJmBMRlEnTOeRo2DFu73uH/LC6hc+tCJfPyfKIwYm4JCL5NqmyiWHzwgjAp01fi
yatYIXzSZQsK7BYXt4ul80u44g4EL/x/xkF+9UvTITqzQbkfTWlAP/i8YgJYqJpO
cFYYF4EJd4Qtau0I/18DieBbZ+3fTSiE9OHawQgfGTA/yKN2i/waWI/YakyLndfr
P4yGBbv60TmjncHLwr0aZdhqz420fF0FeDR3RTKuZYILLup8P9zq2he5IagKOJ/s
BI5SxeM9/l/kBe2/hN1RIHgM4SUt2NUQlBLYjBuou7YpkEIzBjEF86t/WoUAvraf
cAOlvycN5D/N1BtsxkYYseof7PffmnAcKkDEC5Y0kgPz8+Pv+LYs5xglEhqgUTkt
wCwp8mXWSlNycAvwmgN23VeCtsz4NAOtf2Sxx3ChSyCAnwQ+fOsQiGKpZlCrnjhk
zB7oO9pet8EozBSxP+OSlkiGklST1E0GTYl8/wbzMDYPftuXtoG0/tYXwoo7l693
gZzlMjcaYc9NOC8F0cEx0IA53pwRLdGhNVtv4nY8w3ClqemEMznhvit/5EkQJqzp
Rln7ilrHgqx8fbGdskXfWL0GjtT5nUAfhs8cww+JyVk62VlOQufbHEq22kaGKXvV
etlBxAjHd9h1WIx+AQIiMtrE+uASGTDe9z6Eup4PKNJ8RHOufEcyKeblK4NK5/wV
XjnUM9tmRsGHyFv3fQBNz0PmWIoOEOyfHYfK/hgCBl0bT9ib3PBHx9Zuu6qKhmlL
6yJ+3bY7gL+IfyQA76lEz2bzuwLKSrdo7KcIJdV2Zu2UVR0IKMwImZoX9/wjPrwV
70cDrs//3gWLlJOtfZHeY+bIH/fNiGVai2Do669+F1goCPhbnPf/Edtt2b0539wG
jdoRjBq4yss09Zw/08Zp4jXUY/AbuFnNa4Mf4DbFEyH2DqAU8fZU9a8XRqwgih0n
+nY+haBcXjFgAH46F956njPXa8oU2GnqswiB1hROT0fdTB+A7HYXo/HUos8kL+58
AarK278i5KF4Pcumh5U9NT4Cvcbwlt+eRQXaxvEyM6vVjfngun0QH2J3uR1BdG0F
NIFXHLxUJP5kCIxLpFjKNHPKs41hcobTXk3XfeWv+kvHEpZPsEv/2ZC/a+0wQbko
smo5ox03poZuHk84KUFZIj9Fpkp63MgWjL+kWWglON3Igf8m97pSKmsJCvoACA11
A7nQbdz6Vk0QAvymLoE/tH60K8P8+lDHK0OpPBOmNWjgDNDze69KkVXOAxKt20rQ
L6i+PrJySfndOSLYCtNsJXBv2WIIgQIRGH9jwFXP8ydkXrZEFmhelbm0lj6wWcI2
PqslRjtbpydVLh7cwItJeU8vIWQLkQJBRS5qdd1ONh/b24Ix8n5wpdhqn2oPMDfl
8eRQY4qJBcXgREaa1ETzXHtT/0HRDzYgqA2P6y4v/m9Uhei5Urx9CFf4ukkrb9y1
VFcUwnjIYjcxlk9G7mPpDoBxQS23OopCk614DKLCmwCAahJ2floNVhpKIFZ6ZIjx
yHdxKmCBwicjM1evvIgFtDCmaGvVvzOku1pcZqccwSURGbypXZancFQscHca2+bd
yy/WOSh9rBT5tJyk/+eXddVRSrAUYz/mGS1AUUT79vdIlRNcRiDZnPeF0d87vbsm
HRnXrpyGH/PwlgADmdkNIRPZin3n9i8z++V9RLsI4XvbHsgpJ8sg06Mc6Wb1+szS
0ucre8GJbhYPzqyvu6VBKwG1hMPl637pWhRLGJNmona7TO3p60ntlr3WrXC9YVWl
QOSnDi/akdiAUMNZslUv83s+woRTeepAeXBKHTcQGCY5y+3a91lHXwUK9fTfx/lY
vDX0YnvR0DmcEJvX+Ov0CYYQ0mp3T92+Ubeu2YHK/uSfiTKJukPkgkeRigs/shYS
aWPleofasNjVE8MUJuOXRyEJeQ+Oao+Ik4YiqO2ZMtY7lVMv85flum9+viNVfow5
nqZcc+zrrhgOl3PeBV0gMhAie8JYN3y16VmL34H3Ol6xU3GifM1i4zTvCzB7zxCI
l+VLiVXzeuLkQXsNy2ZalkJCFHBDDgtz4jT8uHzwKW/V7DtPVScYZANs+FIlWOS1
jiE7jPr85YrALRQZn39xtn0O4ja3E90OcogpqkGaxGZaEF5NJZagPuQcntZE40zl
/JfBVzA/JXa5m4VmC6keM8UNgx3rgM9Fu0vEfl57UUZo//8CDQFP68DIgVUpU3pX
yx9gbhemosYgjuVyRp8/ueQsMstfhjfw6uyHoIl0JVzC1Agio0clQXjVsLwNMwuU
oIROBOxoFcRAgbz60ogAGNN8+tOis9WKAYtY02gJnVd9runR+N0iOVoS07Utl1h/
oQvqY5gXXXlJseBpwBktZbifoHcjlWjWF6QQ/Ux1t3ITq0ghm5gt0bMY+ZS74oiT
ArCQA+zD6PIfg5X5K5uBlcb6rDpD5UR96vgpgqSDXPMvuBheoHal2a01V9bFIuge
wP7i1STCWdhQj01HAs9vkJUWV7tdtqmHNk4haAw54/UutT4dH4Xi60iugPrwiO/4
+LB2McydE5KmUgCwLGtfIOfgWyEkyJHj53YkZ3eoBLC18hdU1M8FZKrdjyJ9BY8I
RinkAvukMswYgbEUBbYgG7m3iAd6lw+ft5Xq9tPXP76UZ+StUbQ+Mu8lx2wMmCfF
sdkBC4TC31szfjtiyLq0U4qR8q+REuRrZJQia67gh3ju87lW9KTr0vUzsxJwW8Ci
R0sRPZbYvUlAuZPU3MTEwnPxU8/p/LHjYe0c8wcHivMIiTJYbKNvWHYKHOUmv7vV
BOPPN9KrHJOXPSDlMhDP7J/OAjTGayY8+adb/WSGQ72dBwdC0w9g0AR4qoa1pP6q
LfD5hqv0D4qaz+MQ6LmsSR6KfUwdbAqr+QdxhZlHfMuIO9qRut0DSvAFZ83ABZSv
bUMSN7koXXvFomM6kvpq/87zrXfTeexVPPS4vPoPjLHLs1DI5YQ6kx/Ko3G09pKb
ippaFTA9LEuFQtk9nXtuTx9JVjIev6UAjaMuJTqaAreRrxbFSa0XpCiMGy6yrFbI
DndHPQzkgZIzbHoa4gLJXJgCUKmMFkqqwpwOvWuF1vQxgcFHcOoEpzQAt3EFWyhN
QosBwhRppHMMnTlzDSbY8tDVOffbQFM9NhdtxqI0PCpKovjaxbljg46/E4ZJdg4t
9TDfROtQQvU+k3My+25GDrV0wRh1jmVMKBefCoaPHhPna7rh8Dwp/PtEN61JIvTv
vOSyK9wrJ1dKbpv9UFpbqAQR1xHglz3GlLhSWWVB+ZipVF26AXAnA5+xA7sc8PEk
3RdQ8TJ7CjoL1gwpv2q40tZJlJDNNx1g2oubFAIoMdyiyf5NN5fZWjlyl0t1OpaJ
HiKTDpKUHyMQOTYAcM61p1wnH8ebTZJOfRXCZISDu2N/uP6B+8LTD3pgy+0xag54
TdT0NFZ/UzVBN9VN/Qmq5hz9FYCIueRBvMM6v0tGK8i/UMB0c3d7KGRQMSLG3gEy
PQ8cwNEJG5aOWPA2qm9N2rsBLNf9w60rVwgTYThafscAQhRhkxkABaX3BQVgT0tw
pPfarPW0/UFZS7rT8YAdkrS+iFqgw/G2wzuauMvrS5ZEZSdsMOTJVVe9uwH8KMWz
iyzZTtmjtQ7fJuM0bzurJdxndvTbyTzkQ4VtLomK/LLt9T8FWTTLBaDQtDm5/j2G
yhXLFrzPsUyO1HlJaJdC7dDqq6IYHTGBqharunQOCW0cb7E5tPb8THzxYVBfx1II
RbuvmEV7K3uxd0BJV9qrffiT4Hewer/vfTC1C7Qkk3xOo6WbDHjwC+mOEqq9yIFF
lbpJOymJASd0wu2EwDigo+yhvSaMyd0eJ+ri3pg8WhdqTjR/+LDfpVYn18njQN3x
R7E1KsKohkeoHftW9NCo4t0Ep4MVteO120x6P4n/sELPMLfGLF7G5gBs3tbLmS/J
xAZJ2smiMCQoAgqZjpDWWxD09bEFKEL0j3OlMgu3B4u2pk1cRizxtV7dBmN7nlz/
ZEFOsWYdjVDCLao6lSMBINpKKG51Ig1pPK7UMtNtvU4wjJeDrmFkZep2L4RGtZ4e
IxALpm1C4Ny0hPj1+dqM/Riz5l2gtBcrnlUkiYqL8pXMTNO7bAIrPEJelzamseS/
Cdoc8D+d94bNPvHA124CKEGxanHSpVuuuRgXD3PtGp4q5XvKdyOPNNQHIuKI4VTg
bu9sfzLP68hd7OBgImrXI/Dx6Bf06ACREGPUMzpU596NJkMCJYR/bTIMTAV/5Ukv
rOJv9+BiLPFKg5dLnNjxSyLnZ2aMhAoaHx+gx0vDtfLrXEtkAbSKs4jviXPLYYWr
b1yFVS0tDT0n4DiKBS5nslvtKYxlf2HO62W791d7qDG2tKjRwPqDqL8lGIfkDahp
c/uLThSuaaIm80LswyYT1kYs20A9kqsTxkDpTCdj8+G51eolqYTunopgeK9UdVyW
NRpikQzqOfS7h1Lv9YeCWgYSQ6BOqeVXSJnI7ACNYn5WRUY5RgnoF7IMl/wh4rm5
Wdg2wxVz+hb6QXOnU7EhAGCzADjNCKKf9r/bsHx1QeR454e3lm/8cAKBKwmw1PL3
N3q4G0AO44cIkSY94Y0xcptUbeMyTSY2AeHY5UcdRtNDKsd1GSNcx7vKkps0OJI8
4ahlOCw7CaIDS0FZqeTUPeR6JMpaKD2HpagrDEMr2gEcxbEMFCFMcLbH0ViWoMvU
RfSQ9EnM5nogH+fCsxKvRk/IijUWPnmYQtLnYIrbVz4xT8PcCXIpTMagc7v769TC
X88HVNoideUd85vVPwvTO5AwLjxWVyt3fNbQ8Gg2ByRGG1VScmRPR7VNxDqraXcm
aPMnjY+w/8j9EeUJwtcubvjU17KqeqX09s/5VWxw8POBcir80URsLKJUBrMQy4lv
lMrioxTebl9z0hXJlmBasAX6bn+qrOLM7p83wIbmM5N/fGnJieq8bYXX0jEKAYc3
N4u4ozhzSn9Vob1Bw6tZ3GmTnKoTUzuzUCDMvyex0+1sk/imomBW74Av4gm9j3qG
s4IL7WnfECDivxDVUPp9tMOh/5YIPwkUWTgWuQ2DkKTQFRqSUBHBqJvpwf84rOdw
MpqkK9AuA8aQkEJs9vAZrcNy+mRJWoyorEHuWHCoWEmWePndQ/guQ3RFcRMXK9uA
K8SQSMrCaXCGR/QInjOKy96ID6HMutkaqR6KH49kuHdwRAGUfi4jTOlhSmdoH5h5
mz5W78wt4IsJr8HVBBTJ2J8kmND1wy9MjO0Q8SWgZh/K5mY50jJTk947h86rHyhc
4l+Mk30KL5LweTNhSv5N5GOKaC2aqd1Col5wGB9ExKX/sm+eSRtmChi9QvUkZwG1
6K4GhUZjKexKWIIbmBoG48MBZgBnPo3UcccaKDslyUPgACSrJSE16ea6keJTAajZ
bnoQV4SP0cUW5oPKJHUiHwRhAexYyXIDr7c+EKBTqeUggdWRvS/slZHdz9FxJu+T
sJKTwjU05J7rAaXYTk63wiPUlI7vgChn4fC8fywnAM2E+s9rjTqY5cOTpP/Pu+HA
xJcMkDd4w1EyCNpLZQ60l/wWDvhPv1oFiO5P3gyrbaltxTVaSfbIa2VUg+so/az0
IQLaYzICliB4ey8TdAjukpjXKcDlf6dixrAWP9lQIuCfqLh61Yiw7W3TjCygHyvn
oA19dIJ1eiG2vsYeyQAT4FW8s1LsPZgQpDVDOEUHUgfyfzSBbtwwxBUorsLe5ULx
cxqAJ7SeVbLWgFCI8exbgdxilEAIqElUjuINyTTR7on/+GT3BnHwlF25x8iqSsyz
DMVMsObmJBrn+x2EqbwsmgjrVbdJjlo4O53IKwj+w/UnZBgrkU6sC9cPc8GNiNFQ
XlBdUK6p2DoGy5I+PlBWuLDoIbEOIiVhnS8VMb8xNTUxAUD9qnICDHPbviCccAXV
afF6wsUdZ4aChiOimYYLuYl9EJRJlgzeadj2+o3TX2Gt8iek1uuiCcuDD+CJorFI
LeGL/gIsaWT7YjIJpF12Lxvpl2XKb2CQN10Y7O6K7BSNReHwXPD9pp/bhulk9hUg
7U2XF1Hu9VklqnQDCDMlaOjvpAjYAJ6kK4OMp47mx4ml8WgQtBG89gFMFGrfnAd8
VAVQ0bQlnZopCOf0MtORaQjGvqz5w19496Rpof3r4Eo61gGvx3rwVaMMNUP/o+TD
7xfNuV/5oyNberIut0Q4h8KI4ks2dm2vyiYIgYw/MnWhxFI4ioVyDyCs59K9XBSU
BbnvGH0lYD2Gr3YhH9auf0ruH2BNVw7oASvzRjD+yK5/3MQpvvE1jD5K/xHPn1Wi
vLSk71ytqqb0nOwzBLcmJK1tcDgb3LntLItwZqqXexnYmBNXNuXhbbo4nYWIHwOJ
owf11ANcaqNgluVPTgxdWxaH24J1y0et645Njrb3eBupTjJGjELnZeYde/yy24YU
Ysf+CWsUPH6j3sqARgXPLtnEboWz72Yj9iqsm8hTKN0atuW7NH6rK+GtQMBl2EO8
WWVT3SKLWm3jvrE7uQrL09zoF81nLuQOPIQcYl9lHKMhGQMc/9hEGZsckivUJkI6
oglvUJuCkWh74TAfCxgCJ3cRAbLtpiFYwQgLnrdYWIdyU1npqN4erTGY+No4IHwg
POjaVhQaG1r9EOwdmYcrHrOqQ93X8QSduY5hYgXgqx9fDf3urPusQEbT3GRNznwm
zPgm3EnHrQBgaK9qs2esTCpgL0JQGXkRgMn40UVbuTEHIVvgQpyJeY4/b1B831jz
76ZBe6tT8L/uom57UIlTA7E/+G8HsMUV/+ryFXbFg1f7f32k/zWjFO5MsGg6ZeCQ
T3ycAY5UdrN63fwHtrARQJqf2+VfQPo++t6Co/KisYOqsVvEjvfsc8e5c65gKH38
Ngzk65mwfcwL1dCLVgdMsm2sPyIIHbEVNjXR1mHGcfMZyRGp0pniUzZhiBoQrMTJ
hrLGfGMen2tlaI55qBwf+MKLIMYHRfyhXTmeudBTMZa/mI8ikbcYv0iSftKTMsR0
9VgsjmWtUk+MBEgBVP4EDrZxH4VlIO8POra7NAgi7vNiDMszjhuAK+IdircBzd5P
E01jPfnhpe5D2RIFLCWARxOOXZu2T/58YF24DYikawKlQ6QmO5VGOL1tJJ/zOfNY
Ea8xFjOFiK5yJDFKpuOYdgsrUp8NoUV/83iaAzGiZXauEVo5pK8ivd/pxiL03b4+
q7AQYlTMBxAB92IW9WxAqvL7B4KWDl6LVQ1KuebImhwlj9fKkeecszFxCIEYl5li
c5adP2pDCtn0JTocOSSN3SLv5LaeINebaZrBBOqbSfcXBwkBYw3feNZQKJI0OznK
jW16zwnzRWaoAvSxyxwkNr6I1LMeE3yS8kiDU1iRniYIr3FdeopzSFpqeB2zjKw3
Z4WHbIhMbJ7NjiywCSgn8qyjVuvjoct7e3dheZj+CmnS/eu7iuYMWFHIToZ3ZZS3
he0ZEokct1vGzrzx/mstXjI6BD1jdUZzGFZRw7VKCGuoStPItqaTuTRoc/egg/jg
Yq+CIL8HlleJoDvIxbzG2qGaOwaym2Vayc+1OKiOuksSj/qZZXqt4+9Pdo06WP00
azSu8PKv9RA5rjfcTTzPpRpWdkYkjEPWplSyQgsg1443EGOctV5qxstEmWsZVNdC
ULQZHw1pqfPSWTThuU46zBKJt6JF+hRnLCdOuX/GH54ZSJIDt1HPILYL8P+1u2c4
3gqnmlxedrYbDGMBBhJ70YQgqbSqmLDsE3pIxscJ2f8lmNtbfHEMdWlNcKUge9Ax
tkyArdzrSx+clPMYVjf6Ru0IVOM0UYz2PC8ntztSvocDIecmQeVwIlsTNZrxoqRl
BcfIt4YRI1fa3OTJF2MBTgy74V2XJsM1lwZ993NJR3rsngMG/gC0QT5M1r8WIOkd
PzgwOzjAWDGuzq/e9Ld/AEcWI7iM5QuK56pnZ/d4ujj45PrMhO5d8DBJkAbNJnW4
k4EdaBvG7qfWN2cr3MjfJ7VuuPtMaSp+/3cyUBDKlXDCh4wWvJG1l1zKyWa+wpmi
/khA3tyjahRznzlDAZwwgABsJHenjIH+wBY4IqRArbYT25E16LogQAMw2OQleuQU
+jHo10LaIQixF++RbBhR6Ydn+wO0YmeQ+ZeQKvb0Ka7tolbB8WQYC+VIuQ2z0DkA
waPBkB8adjuMoO2cTAQCgo9t/ywAarBvyLeMHV445eEVYwowa/I4S5o8VUsMWx9N
OU92j1/rmcV0TuvU3JzfndVHt1kM9UV522gI7z0OrQcrFHF2SpfT7gLnNZs0ImID
9iGv5B3BAW+7gXOcnojQ3ciSzFqjalT0JarzpdZ5tP1d1LnLSmSv7ykKQ3K2Lyea
aaBkFhR5PPPkajW9CTbi2gV0AX3FAhOpHzsj5NYnggXfsBcGcRQXLbT5STMa6mp6
PNSAp5pGK39eljs+gdKGsFM976C+zE4Xh+DGshm852rC8c5W49QyMGwL4p0vqCvg
T7Q4QDtOV+BMjASViXtgCb8NMGCH/pMaIWWzCjiWkGSDU0q90pAc9X8SyHGuT7nf
zK109lKJI+/Q68AUatulD2UlBfvlsVwQuQRL9Db1WmoOXycLekRaHESyP0FOqfwk
U4GrlkMlGqpzspUcJ6OEy7NlIv8SdWv650bXytEqRNLmPdi+zyd0BwIkh5vyjyhS
6HvoSObae9kTWRLDjTOMY0M7QyfZ32kAVwQpyuxvKo8OuzQsp7jVaIylT1ycFJY9
QSvwDt9IiHh+3HqcMq+U/YWqO/6jP8gyP3+uQhXjAjrmdmMtuVd4U5RPm2bBtzHn
8Kq0x24cm4mA8/7axmskm9XgIxgiUBMEvOtpAop9eBuxtoyksduqTUFbEAC7Vp/G
NWRX6Xd4Wd+Yt5+kgSdQJFER1itMb/lwuKxcF1emEj4nILriU2kJN+BtLSUi1HFu
3tE28CEAoS+wP08NTsux01aEwMq0dv6GQT5c/6RSWuCLUclF6aRpKUfhvVAo+XRu
IuZsx05vU+6XijX/VHc9eRrGCdIEvp7pxaQRZdIx1Sfh1Lq6OzP/ZiMr0+XvT3RW
B88LWD87CFhCUSXFtaC/2LhADB5S7yr/xWxRziTg90Gc9b6PNG63guwLh7fXuEyX
oLRSU8Vpcw7P2JROWvCVUOgwwjnObSWkMlewJ+mjXWfBvJMaisUVb7hn1H0f8hs+
FaDjSi+9LFdgm84oe+4B2UOcDH1YVTwRWBYILz9VKQKVUhQBDF6hqLYvpt82dpN+
27L8jRO0E4PfYS6TY2nci1sNlA4S3aRITkSGhSg22/JIgbxrDikUD2HrMpVu2pbw
TMw9FBXIJV4C4msVEgiBRsQ4U7PxcuvCndx+sWLZK7m3tChi5FxBE+Cy+HaNuNSC
SY2FBpmcvCiHo1UqedIVGNmKG3lsSB7x4zrbHf6tpafU0RYVXrFUiDhnNTCgMycz
3TlfxQgZi6zJPVnPHGQM/zxc54JO5WZbNExbNEq0JzyEH/7STU0HVwZ06Z6aEXUu
LX1habX+c4qrCGn9afBZ0QSIhFmDbp6IgmlGk7e7pQfmJRaOFxSA9wcf+CBKyYaQ
YgalsgeXbdg5iKNbfZWmD59LftEu58MQZv1SrEE/EP/O8YcTlOKPILFUzIQdDpYL
bj6o+BF3LJ8AMTbQ6hxtc0LwBOOcFgdRlFW8SQEcT/bIwSD4awXXBVPWdiz6oWSu
QmK4hAeTcN3goJT8BV2y5t6MIYeK1XC9ZB4o23CPuZPZJufUUr59P1GG25BN4/qU
8Sm8XBpjNq6mD6fIWnulziu37VQJYKDR418ISGbSVrJi5JW39WixnFYn06O07EaA
g577xZryQvY2mq1m+xCeWLYZ7kT0gAUofQ2wn9g8MXdD377lRVOcCBPJiKwD8hYM
O7ZHdLRTd4z6vuUYhTgFOdiW8IrvpCJsq2gOgm/9Bfom6NLa8jISVIKnPYbuu0fM
70LtCa34R7kwYxEPjf0z9oK7SFpFsxkszO+3F+ld5Y/9ZGI4+AYDciP3XPZquiBH
IyGx0M5pOBYhtAhfKlnoJ0uBwkJTGxXTTVseKD/Nj9oMNOn/ITgPkWcMZ+m7NmFJ
BMpC6MDCTJwc/uDzQRtGGBnKjORUsiH3HKH/2FuUym2u+9DDNzpmc6pdN71fLHlI
eFCmAxn7QchrDL+WOyV9+wl5z6JJ6odfMst+upuzP1dqDlzstiF69YW5XHUz42Ps
2rzQxbM3IlWkD7N/myI0JOJOfkQURl/ibaroh3RQ1DxMxSqLB9RtgeBDsEMpKx3q
NHd+XpbLR+tFcCVFz68oV33M+fh4flqHGRGv+JdT/Gj6aSlEaO66SHLGOL66NntH
7UN7i9+T6Bo+NtHEijCQBL6/gCvlhmnHnpfEau2rD22K1cWupjJ9z0+MS9pJG2m0
JmJ2f34YuOigdIduLEEHgqLVpuQF96LFb0Fd5EpAMCL+MnDUwx98rNuGjpZFCu0S
vpdxWWYG1pNjAogHUdhJ5SR+l90cYOi8El+Wk/8MZMqiaAusFOVW1NOeNT9F0SrT
yGILz71h7BzDFly4hN6gLtyOA+8BbCOLB/PfOg5IEYeqgxnw/wWiA/uZOoJ8Gg0G
bHcpv+NAKNoXZCl+/aMlzHYQlrVlac09Myem4Q+J5YuNScllXcxJEOxviVVCVLCD
o9Lg10MXMAevEPu6UepnnkjyWV/ueMjrYnYDDZNP0CkG/PaAtCnLYHe88HEiog6Q
Num3evYr29hereG9xthLnfNR6CFrawiX8dhuTEETXBWF56nHXa4+LN6TN++V4pWI
MQPzaqHrowCj/q4ij1kbz0dNL93gsEvyVm6LQOEVugaAjZZ73ctOdxdEyt6tChGS
BjWunB6aBkCcJtOGh2xjLsmn1T3oLmY4jDTVjR5ELe1SZMDfvYzRfUGUkXxe8lAv
dNwj/97ht1I9uqkXZ9NtygSbO0/P8ywWsnk6HkEAiAgY118ItswK5U7DRlIuzI2J
vfVBWKEE4Z4kNuUnqDrOI3w8MJ6Xp/tKOkfc5q9faEKGr9THm/BIJILyQV7MaCwh
yhucQ0w5rfOwWeZBqJgMV8xkdC+QijX7RzgMaCgHMfRy76c80hQ+AQz9a8bDPFZO
esbamR+nBbeuMD4sCZcuGEqXIF/WWYCibbRmGlsZcLsQa1+6b0Ef5MUl2kGGbWqp
k7KRpcuQXVtSJ2Kt0RnUU+aebR+vfq4G1wFKSr4UfOv7/HWtCzKBqklKSTfnrjgo
gXX4rgycxVWMMVcOWFG4viRKmNL4PeFOeveKccrI3SKW1PoZ90/cZI+kMU93/Oap
zp0K/DmFhS4vMVtFKDWu9A0fFnsGqs7XjzHgKTMD5sREQC/hBPdemuSImLPBA0rp
CfewpNVVDdUDKSMKlYAPjYAnlBtx7T3sfbBzz3BuM9NIz6j2cWXVBT89wnr2rde/
uDyrw789shk/6jpsfW+DOOffs0G9iyPqktIo5OJOnfUT2PpjNM0x93sAs9iCJ0iS
sb1s2y9lIxwjSojTw2g4Bv1dM6R+EoUzv9wC79rGn+wknyBrvasvaGgpSg+YGoSV
2Y8eZ4WbSjnblDrWhv7Er0NBu2C6UC/DrDKaeCUmVQZA5/PRFVWMvfaezLOOSKJm
cKg55VlLrCHeTgTITmjegRFP4CxviUc3DMG7wH77Zvcj/7GBUpMKuqTlD8lNR2dX
KhUuU7AwccnLlb/EpjlMfTp7RbJ3uWjiP+bLnw3rLc6G3a+XuqiTLJZ0V+bLk0LB
DK8Jx9qrmWI/EX3qRb0QZfCdnge4kv7jMYq5MAUQTgwzzuHlcUZ55Mdbnk4qrsiv
UhXqGY9n6icHFBWguWQX6UsxGweudxZEJJxTR9JgKqT0snZMuVLWvAl6CCefeeog
7yAMBWYxAxvLrEuwKj56ftTCZfGSOyDV5RhL9BXVMNXGCVn8idKO8Ktus0A558IJ
Yg0zjJvjPAHw6vDMGtU93vay9ZXJTHZJEmnN6xl5F5G+ZeV+ZwRzejA0Phjhwriy
PUz/5+7AmFQ3zDpKuVRPZRQLo7mRnn0iE4hCE7Igoe1Dx0/mv0pWGpGrVfAUwzbY
hgjYq8QI9caqk22CzmEG0ZpcMlZ9lNd3u0MDvUTur7RMQWYM9wXxLEuDbxafJcBb
JtHsxoO3WtPtQ2E8HcmNjdkbSli65HJBzLI4jQLpqw9ksQhmMT4QZqt16GcIaC+A
T+GgYv6xQDh1v6xx5RwCuLW2Yl+TSPwBVPZqed3eL7WsxxXCkalV5H81VvAWtJr2
gGKq/Ad6iehphO8mmYcple9a1ApPpEWu+9mDgXdmKVLc9AOUGy44jw3Hu7Dw0OaT
IhM/W5vSD0VBPbKpJI5gGNHipHKs0P6anYroXUOKOCL7t67ZFf9MNQZ8Jxrd+UOI
VbbQeF1+JsEqk8VGUHGRXia2dV6dFYPRzaIlwgauvXiicTM5lVn1n77sDShKppMe
AduV6fOOQDSsKY5aKzr0NhAldHXIS1QPcaOfx+u2HEjVMG+hmOIwjWKUof8LSMH1
BluSCHk057NDMotoNVLyOYi6NWI/sn8dZFeABVvJu4b/JtRdZ4tbdeO3HdwRWgRp
ZXVqQAPMK9NrY713SNJZDfmS8P7Niirj8OBLAtpDqWO0AkmcBy5RQSbeNEvoCNEt
hZGS93ehIRXw60+d/UT+qE/67etSy+HgtlNPXDhdOo2fhXRol3Cq+X1ImjPLHkQM
PdKLC+vFCdw1qidNDvlHkdgGYKmkvYsDo9sW9YyshEjUMGCUssUi4Oq0jIOIQIRH
hKV4YxWgj0oO7Pi38maVQlOF7c2zq5TgcoSN20Bg6SZPygQEqy/0tcvDx8H1Ith1
oBVxtrLRbOSwfi1zIXZQkiiBEk1O/atYiTZU9ZxtsH0cVsjJjCPlQ/ZZawDO4ZSI
AkwgKb6Vgc9NwkAIKbGVH+3JXDWS+gUfCR9iHJHlstmi4nKgFChdaWC+z5BRObnK
HhAzUKHvMoCahx70zx597bMbaqtbSJnvBgGH5N1eg6QwvXaELnLLkE3xqs7e2jqK
z1cRig0eWro0v78CWUPZ2pBAa/Dxi/BXxgOV8wSgTzZVRva7hKbPy3Yk38DIX3uK
A6UXF6Ft5FxVuFU6vMNcfYV0SowMeLB/ZVIbbzbAW3wFYwE9DYcOoFXwJn2w+gz0
sTg4jVuBhF1bhfxQ2/qUKoRT4/d5t2UChRb3itzHCGcW2G9yZ3XGxxXE5iIqaNIn
sjReH3pz6iahe/1ZqemjFSwHcwo/snuhgpJjpXO5J2K+My3g2GifGMNuRe7iNTYE
IuUjGjPfZZyeUXMoTQLt6eZCGoYgQO42a6Zymzr+bVCsvmsQwNrX3KM80G/FqpSh
QSysaVvXYMFoCyTuR6mnJOAsSpleZvg+93djEptUPEKyKZOA8Ei3ez3pU68mscek
s8/087z/bHbAB0Je36PfEqlA7dZ9x2qubXzGGuit+rjCIMyYMabnvnJbLgav3AYk
Nhig30LDj3SXRBRk2m+kEx56OrMjtSeqGUw0MEqFXKDRhVr0dRhbj2fwmD7N1oBm
cg1DfZrQFWCVGAAYHHnPYoqvSVc1uQKrk9zkYtoAsZB3mEh647YDiysCg7S/Csde
Cd9KViD0M4dAdTKte0Vbd+EH0nIScVK2CtgmFoCYhOH4dGd2Aycs3weMJErJXsqs
OYbwnPZmQFwgx02aMQLx1VovFGMBFZ1k0+mrboGBWjUQv4DExqXdLUCoNxcOf0K/
DtJAilDmc1g2skJv3tgXXYJ84RGJMiBT6PtYy54hl48ET2FAwCFl9FfuYg8VwXJw
zpTUTtKkSyRpwvfCo3esFQtn1F7hDAsvL3yMpZ/99gkeXT/CKS+djMUYIUYNmgs3
stLp+saAXS2Otv8U1HpoUOdT1BplMZEcLf/KUIMGMp4xMOstljereVWXVN0Xpv4s
629b6Ay8hrOAyEmbfR8lWXKN0D69pV8Lq/yOlAH8hNChQIDl+6sooFMdwj4TnoaH
j+Jwsfzd5bKuqiEPoGNazv98zWA9zwnXLfZquBXPSizv79+AoFNQeT6XrVZlWlVB
u6nFTFNIejrgyKzEjD9jAnZ8BObqYOwPjDHq/zX8DauccyNGC7QSxtrsO/VIXYSH
evwK7hTDJfztYu4dsIcPcnGzlJ+Q7diknJ2glmqEVOmvxyxjRHJ8qQtk1iK73Cfv
ppQhjuszakgQPyWwlAvHg6jRlcZlyyVf9tAv3Kg27dzsNr2NJtRYDJXt+w5k9rAE
67pfHV8WTGF+PlfwcrrUCI9ajjmojwGwF6CpRl2a26lC1o1o7pg6eMBxludM8/9m
V4UQrjs0dHa5b6bfrkROdMPc3OcQ5TFwv7rXScYDMG1UkLCM8q9tx4NOZ8OOw/mJ
G33QYcOBXELa4nfSa3KNSC6Zi405mnUxQKi2+0XHiFRnA2CBFMixyeDv4VYfLOS+
iYXxuB70u7ivAYEUSIbQSxSAD9cwKEXN5QBYyJhEeRZn9Ak34+lbjjaT1a3aj7DK
o90WyGO7VM/Jfta92ccEjlLXLT+Ri96Pzo7LofCnrOr8iEjeHz0/EUofPYSY0OAt
p7ZuVq/ijr1xYyY8vay3VXapqt0ubi6C+6mfrfK/nsL5KTjNBhtrNs0J5dTQ4gka
YUloyyeJxHX6m/BhaekFqp3FKn3L9k7LCdt6Dr30Dabr+3WeMItruiJRe9+9pten
8uy6ekCx4M3xktzfH9Z9xp3T4xAgkJjmdBe/H6R/WzTaVQyhIkjpRfaavV45WvDP
FYRTlDgPOYvxf69occ7Im2T1UeMiUb5GIN7TXsX1p3/1bVkl3FWwm3XmEulSpIfS
VhbMZeQPlFhwV3mld0PvKaTHggEs5y8Pi4ORRfCFoyfxLclxHFS4xfGuLiMoRcgR
/FUVUjv1CClzHtCsR0dzKT9u0x6E/dHVVGHX7ILjLxE+AMGkG+RRVyrQkN7TccQy
Opp7pdcIuGOVc1mwYoRNn6AgZtWMGb+IWqlj5zw2rJ4Q/T4KJ+/a42p59LO+/IGZ
0HKvTJQWTFEQNaFqlNJlp6zh2oUWrwbxpXBd+MEgSLs3/tW8tkVfW/T8rA4xZY95
PnA3SoE4+tzYonwS0k5AfF5rTD+ApUDNkZqQI/Poe5S7GTOude//31VTs8EnsWOd
VVgIEP1Qd9rWUqXM2YsbhNsbNy1PnU/ZHwrwJJtXpsJmr+Ef56V90svcm4kCXpnT
CCnbRpiYOccXv1lN6FHtg8gFHloyIIVA+zSxMsqUCvuOHmaNkrAuWbQnZx4GVxy+
f3r78RfyTIhhdV7xNG2qHT8asmQPLcz3mjkCM5nAd3sBhD3N/WzgGKCvIwMqOmD3
5B6016rB0R4R6Q3y+6HQ+XoBw+ueaPc2DL9s3XAjbVQYYkYgADtA/4dGip5P9aVV
GTCHBqRzm0XerjCkHYIXIxVjUtWZw984f8WWmN0ww8/AXZ+Zk4xsutF5wCTnEcDI
ZuOsVwTSarxoB3K7ih9q0HHptc+e5Te6UyK5YuInkIEOl13ZI/KsmtYpQ1MldcbQ
AMhGvxkMb95dkVLV594vo4bBMxXCOim2H4zGZM/PsVBqg7cOYBBVTs8va8jvz/J6
r4RN9gLkGo1bj+5PKxqahlrddC3G8/UVyHweSbTZxVaU5fb8eXcxM2s/omkRw1e+
oSneso9StizAXc/fD6JyFIPF9xtuZSXpwfeeO9Ic3tJIedrF3XzrEULgFXregDt6
vQs6kaSSUqW4G1T488z7NEwZB0r3Ow3EBJFCBm94J9ehDuzHKAvRTbqVBZWIiIuL
eC8m4k6t7PpVRMcyf8G2o3tUbgkeTX26ehc6ohYcfXUPJqOj4CnCUmrB2MQqUowv
Tnq8CpKaqzVIOfX+FISUaxXeZhD5W+Ac4SsLfYLO15tsGAKcbQ+25OfjCIFn6XKq
J0qrH2qmzDWc+86w9vWf+3bowWJrBw21K/7WUL6/cRg3g9vZe2aL37H0RA5ZlxGh
YSPAje2zaVmnD+EJVucYABZvQAv8l9Uhft6jqcUiPPPNySukTGd6epMXPlNHULzR
TnIY4EPnrgAY6US++REBzd/Q/LRNHm2qIVjo1ybM7jzuE0TXXFG3ygxDJ4v6w3ww
hYUm10NSK4MlJvrdQZXGhBiM+LHH2VUrKnYW/lqunOaCQ5vpqkpwRLD6RMS/n34o
6sDPuL5/qmB2vkF4QPfCGw5Qi1CdG/SqehEj/w5MlW2KY0wlTja7tPU9I8IejtTy
sZw/WNN5vRjSQF01x3ZD4cIhlrVxIdHu4lBFdixRJPpCXhSRjJvjT1nJD+dtudQn
KFZD1VCj2LORFi5t4IBsDVTTrLikmitLfork54Ja7z6avEa5Mwwvmt9UFccgFm5u
2BihdO21S0X5LluRUiKnW5+2OHIbIQ7olboB2ZjYNKoszwr8NbNW9jksR6yMX55j
xDxtjj8XZD/qmbNfWLCZY/ua/dw3YVN7qh3Wm9xqbOtSEUqJFjrBiwyv7wylCPJC
VO+lGlUFRK0wdGyOyz3m+nR1jupfGYvXcDnTNV8mAnHUgtArCFYqMCUxdWCp7zxV
JzFotnr7+LqTOcJFv1TtCYkh99oLTN00fpbuskywaYPrguXfKpO7tJRYeikXITco
eLVI4NYQtEuJ1LPGax+Plnv9kvA4U4qy37WCXkBpxHPFf9css+CJZ99+cS2sZxIm
O+T9Xh9KSn+mXG/1tlCqkdALs1d31tbr9a0accahMZHBb/z94DouqlbFdEhOLPJy
oKdwvqz+58MxtbewQEK+0/m+5TIoz/a/okPe27cO36R/iyC3iNk/A/JRZIRmWhWV
9RthlFsDCBN4/A0CbmfntejMEikYAgt3cgfoSC038XJBdjwQCsR4GxOdcsgudn4t
BsOd01FF8h7mYbwx2BczQrcldOIVyjrdDSbnX4eDu/XW/NEE5SsjLl+QWCvo1cR7
Ft/LPEOKqL8GHOF90sYai9NJyrAROlqma7zKMbLHr54kCsb7WQPZqONRJLH5LSmN
Wna5WJPtncJJ01Oc6rW2SEpwzqFRzDo2Lu9HCfaYwSbiofq3g6MqH0GsXbKmSbZX
XTVRE72PToruygc0AJX7b2/C0+NliR/u0fSIL/Tmr0DNPKD5NOBtunekBa0/t256
nDC1ACK/kNzr5W9ObZ2kHRdq+1YCoOVK4PygjYjE3bbrua0gCEHoPi8zKUaAgM1I
OJi8sDSBVwE3gDxYNCtvaSrbsabNfrLs8e7YgCm4k/FOwxMFVq5/DETUfVwFImWQ
4l+goXaixgMZ2SYEisLKCqedtbNXzVrCloBwkjBDuP7NtXrLnomn8ZFiATcjamSe
5X9MGZSDGpM4slFiKRNUfITqxvCvtGosQ+rK34TN0Rpvm+d9upsmtlaMU7Mm3iFG
xN3cCbW38oAvWwmgJ402lS1+MUDdxPu4ulHxvx/mkUOnY9JgDRMvH4JYDCaQfFhW
7ngC+zsZevML6dDDNRemom2Ssg7qpWcoRq24C7Lds6BIan2DDqDMqwXEdmdZH34v
Gcaxk//XVFY2x2kziPvbVca5N/ExB0GeyEpO3XXDW7RtJ+SFX9rRnU2fWS6iIkLb
+GbAjJILczIqOg5v6MJUFe3deX18B4wWJPSGyR/qZIhNbBFfAiGf2axUGpWykK+H
YpqzMcM6OFTlB3LkSEAXmQnmfzTU5kElvp4advIqaBMowllBeibSvgkqZdMfgytf
Uy0ZiPJ3178R1bHRc8y/zrM63CRaYwjgGmVEvRM5iFCb9WWO4JF1G/TPivrg+kc4
7sTmBtBBvSbcrP9DQkPb2YF1Mukmjzs5Zcdn8jmX3BA1b43wMVNXBFG0zBfLILRh
IwaLyzboEeOBnEXIz7hJZn85XV0AlPKHbqNFM3bKg/DfEiqBo6J3QlHg8ucJ90V9
Wtprkv88J/iXjLVEUj+QYY2PGV941H3AMOlcf7L9GQKERlO42L5lShvAkPi/MWaa
F3MzDtaEKyBrZfAiVPNoWE5tmcTL4GpwCBFAPAo6IaacP6bE6BlgAFQPueNN2/mD
9xEwQNNmEhhUDv8EOp3p9JYzAvNwQ+kS5dCLn/CNeMBntdsErT3SPKNlf+qp4mgY
6JDFsSlCzd0WmKybJ7SIMcc86iHqObOPQ863XvOkVwcLqTnO3TenRf1m5RlM9ayh
HGNKgnADxmxr0Ms95B406igXY/8UYf8ij63Y96TMQpANB1ipr5uDwiqMSR4BtgDW
cA+T9nR/gDW8pKLo1++yR0UvYPO5opHys0hvtZ8YMsQdikIKIYN2ByRngAo6+twB
3M34p48RdSGo7LSuBcxqMc2LHS+0rvXXkcGfYVmkate80qqUK5jv+JlX9ISSHfCf
5tJ/ltC+lAWVkkllY+Cmp+lh/2EqohL4sFgOxIzavdcQrIi8tHMGrCVq+hqx60EN
4BAOxQ6L1y65f/mXH99f552EeczoYuVagjoB4mtfGO+OA9QY0+TdYNJHNa+NTKqm
sm/VDITL9H1GlNxtnNsVe6o2Qi1LuiEV4OB5C58cITQfhZXS1XpmFVdepYjAuNdn
ForHrfI8PBxgLwD5NeYy5wNpXTJpR3WcwS1QHzxgxDOAzRI5s3BR8i3MNgWFVMDj
se8z7HkSQRmLIvQZwcgmt3/jNmmFVt2568A8dEMezINjStUKnhBYQDhb42YVnHgl
4FbQj+YvRvs0HpadW+SHp8fkgo7Xf7HKjtPXjrZJz05A1wPxY15SV1hLk3DCpMbS
tAdhTcjOnNAlAMBkk8Na3xmpvF0voXbGlfOcTLYoQZX6h5gCo0pSDh7YK4FWoDiy
n/5kx9IGo6Mh53z9AqNGxW6lxVmEkQt+4HrtAF2/6nbXebIS3Bu8uPg8BIbBgzvq
k2J1s+C+KpbbYFmlpsohPU+cXWqQRs2NHlqImoicikqncbvBvHD4pqz7T/8qTQ6J
vUmF8BG0zRXpc/T367VRxr2wT1IilwoJSMi4+S+4S55ItNoYeAuaBBICWTvVFhOQ
A9P19R9q38RvLci89hmXVrqKmDmlHRasPQK3vJ7c/0gFofxW4gbgDznUptVeIxKY
/O6Y+PmTuevfAbJO2CznCcSVJqIRkF4mT5z/bXeq1qP2seunE9waezrluCP9jF/2
+0/VPArVtHF8Zgbwy3kQpKOub2rNcGmwZ8r35Q+ukv9nw62obUH9diijtbF/fbff
2764+gfmNLTrLEae60hzUG/vfjK+epRuO2jHOF0yBe6Tr2LBiJIOmGeG7M/bA47x
hnFM/IaXAOYJHIUDaIXe3e2eGO4wTwMq538Hqib8Zstb4S3i51hMqeYsyiflDIq0
LSL1d8V+9vezD6Sg99OzoMI/H02vwltjsppBOVodvfXQL09SnrP0o1kMqL2pxfvG
kKhMiNP+TV/TU+DbKc5Rg+R1FFgg22oWFiplzJBf2O++m1iaxQRe2RgKmg9C4mMd
AZ9BzY/VR9s8wIJKe+tNptHD5adDbc8G+WQXy99tcMQ3GVi5yowgNX3jpUMMClev
9FTKLYIOAGFVnf36bQ9R5f5UoJ4fKJAkjJEElGpw5C5jp78bw/mwY4CIztQx8PVd
tPdEGUyffVqwb1aPDOCsOINMa1WEhtxbc7v6HJiuIq4kiz3G/g4Ylq6eGBqIiSqF
jBi1bYcZ5cKahUFIv9f4GeS1RICqtpgwLj8RGUq0sV+RPZnQFeRmajSAjjTaNcMo
vga+e8y5XPctse+wjXO5qs7vRRAe8ftLYBka3uuvCXBgm3fhIiVs3QekXSYAOcip
hhMwtU66pDLStnHLm14TqNwzMBg+QysD7czoii5iHvUA06OaO8ggOhNAZByuUDm4
LKXAXfa7VW5XxqLdzolpccT3y2smnO9KRPflRkpwKW6vr3P0BnE6/wV4L06HcaWa
QVoyKCFqeleg1CuJeokIE/426MZrp634tZcRBJolR1sC3AFojG65X1TbZVlNFELt
s7S5shFXSi4vCo8atMX3PNSA4vlHOpRfnzKgVbdFI4fCB8DP3SVjBFfSDfnoR5eh
bQ7yCufE62i6/2Ata0Hqpl1FYoa4D/tU7R2iRzuQuZY5ltw8Hr5NUAIEn0qsmntP
BeVkHZEiDMRE9yg9JGHu+S7GnGdIjqlIoUiMyj+tVbI30T5xvjXobxoK92cLgLe/
kbVs5yerB9c7U8WPDJE8FlxivyUiWbYMahi1oRMveezfeeqjEKfE/fzOEgfuVzvu
EXGtoMHGlXPEVb6a16bT0uPurQx7oT3VFdvjGK2nHOty+Uj0EmBbqFFD3IO3hxQw
PGi8bbFb+ia3B3rDZWecjtWSBeAhO6nSvkxLWaawUx1nvM54CJBXG732Tozdb1Yu
OR6IzCi4Fu4KKovrK0JFBmv3GsIgBrW18qLnsLjtUGYw7gOwJiD/1Yr3IEW7HkTQ
1yHwnjOCr9eiNL7FOFtNzLNwKKdza1ycjleUzD9v4TBYH3uYHrBEjqKCtJ1mY/n1
wJxWpEGBkkRv9xg6xGWI7/NDLp152lASzA1EnadNTg7nchRhwZT4ALqLW9eQp5co
D67OejAonbDzmIZLRoaaqV024AqmEsyV+wI69obtdsDRMKJcmlEZF79EtSemQKqY
wErdH54RBWRnk1qCvhVH96yTN/Y5hdfP9PKJHscVcl746M8C6ypWx3tXwWImkMDz
90b5yZVpszGWhU89Gi08aa9TAHielBrRm3Y+DEdfVLmAuY/cVgU67oXacTWf9cHW
3jGdpcBCnZ1hyFGVdNNAnyvR3sLfkthKvBNz41ONrBLStVe7z6Om/myNHS1g7RxP
KvBiZoh2IiR2+utzffT8oPZHCdB5cRfkXsvwhpbYyqAl0Pm15siExm+8ejldduob
5qlq8EqBjJhwWj8LaQbagzfJBt++uIeN7CTXhccOunPkFivjuKh9CVo//MOXA0j+
UslQt4Ub9sWLqU8GCg0R/0X1Ya1EcqsW7ECiBzit68G1/q8fcKTHKmlNgYs5L7Xo
166LcymV9BUQ9yBPGw5IHg8R5zuw3cBZDN4d/OLPaSTfZlHOPngqLE1MPbQTy+rK
qcDCcwAgZgM8M5Sll0vQcVXtEVoRiNcALUZNX7LQ3/RmKEyXfeLsdRW4O/YVVe7v
cdYPFPBA+NJPtHoUx9FfovPgi6NmEp4Hy2YRE3imow/K/UkoytdAPQbQIDfLeYvC
c85V+cUAgI+kRqPfJHEfmLnF3K1xY3qxmrF++NgcCG5v2XFJS1w07wLpCeNidKsv
aL4keBSJRnp1WNSWrSpOoakmq3hXglbv3oAufM2bvpB9t5+Uw1W7IuSZcKY2NbYX
AK2krWH0/EHRRaXsoGFQ98WnDrr1VGPeLybB8p4tu7Pv0F2gyi203uJlAX9033Qk
yRWId6yib4CbPzN840BEfKW6d8Cdj78DKH5FtrwGc7vJfKyEOdXJ4Hf8seYDiPLN
Tx9I2of96vSmywODkBFT6Kjvv89mePK9BG3IcMaXzDGZ1HDZ0bXwU8qDgf5ctDyh
ZtHcNp7p7RAEDuoawUJtcy5KeRAyQEcRPqnRwVnlwyJ9wRRUqX4wlsdQ9dZoABPR
xRZOYUv51CgdPnR4WJPUwW2fJ/zlhuDE6UgD5P8LFiA3FhtQWUK1tC7SWEr9GWFJ
oS16ORRXuuxRiBtSA6V5cJqS33epLkSPhKGQaw5SmWF9XP/vLEjL6LoTUqXCqw+f
ojLMS4NvBGkNwUPTiRP2RiQrCw/7WzyrlfXTh8eR775DS0jQtS4yLKJPcL28i1eA
xx4ta4MgPXwAM6toLIkedwq1zySVSyB73x6RMJbiJ9a4fy50FI3txioUfkzGxjff
MXxU1/Fuskiyf9DyX18CaxNxKEpOgIfAy/ywBsTkELHkzr/8OnF+ugKfoCu24sYm
lPLXT/KWz7rQRj2lMvOVplz+kzXaVaL+3H7Xuubl0YbvZegn0nBj5wkJV/alTQ6f
c7pdOJRYabNaMJaozijoHeQKr2RxFsx8ls8s60GHC6NBRuKs35IQyCNymgmpmVSJ
f8zxPC7uFa91Dbnp/DDOQzwb+CXyLm70mpxAlDtyDzWd1Hz5C9uWVvs6XGKiqmWy
pwoBq6rpAJnJGOMyhIMcxky7H2kpEm6C5MtpIw1Ci9kFNOlxN3LUvBMt329oOK+T
Dg7zlDsTaxFJ1fPuJ8zHYc7Os494uIarSi5MRkaTbTIOErPPR7Poeh/LqySEI1BP
aCWiLz7o+z7/RxnAUTHKuVPo+Npnwq6YJGY3uTgSs4csEHOMQCBWXfZB8XgxJ5g/
VBKwAjfx4CWtwc+6WyxHGgzCKJ7xIUhZoA2whxLo3KGFqyU+dbC68MyDJbWbo48F
kIA3HpC0QbZKKXIPQh7t+xCvsrPjNWxVTmsKRwDc1qcmaeYIc64mIZjj7EpJcYba
2XU1Jwy68plhXLaQ5xxEYKRyZ0C2pvBZfOBSClXFeA6nyD5gytqotaK0lt/xOJYI
RaOAeJpGWh4IM7LjbVEB3/2ER/9M5mgpFUiL+Swumaidw5Yo3YdCGDolXDzPDBsb
ZvrGDOJgPl4XF/dl1UXBQdq402ObfjkayUZwCh5yVidjC8vM/VWVI8bldWkdGD0T
nwCEfQKsQ6f2Xo6yI0SKZos7otq9W2wGEKVYZN1GUnrJA+7s5VX7PXOgyrS6tpei
DoimS8ie+hNmhpfNsbcwzW3uzmd5alml9DLVXXwyVxOxouKOXyMp4Zn28fE6HYrR
fKXEFd37WGWwPV4B2pI5fh3FT6TF55y+dYeWbhSat3NCh1ozYQKLpDxcCGlOYiF1
BSY3BvoTWuG4SRxI5IBjKkGDo9ljgNz+tfUA+c6AJTcuqQr6oCcauWjJARRcvChW
nGextq8tobg4/wJ0dbcvA2WY6gFtuxjTlS6F1kAD3IcoxtSAniIzyNXOJ+OrYSi5
Mqc5+2tkNyUmEU9PRPm0QgA0d+W6mO7lSUVBhNa3/7vogO6yfy4b3+aCAqaoALnB
rs7/hhVZvZEXTI2TJzyuEDVkbBt+17CdHhQGY6fGeeWFS0MxPh83zsbKatejYC+d
a8HkGq5l5c60dcdZ6sp6rtbFMFyeJ4xAKbhmV0c4V0iZCsp69O8zh6V/nLhv6QDu
ov5EZi6kCvMc3dveVpJL4dleULZaQPaqgESPf56euKIP7jeNl1DslXohFOah5cJY
m8vRJESuuzUcy4wvojFTQIrYbSd89HyfYv8r7Ewn/OUG6ifQzmT7kLueDayV/Pd+
1gzx7y3bbc6e5CcGdRjqCbagN8IONXS5bT0Dy5ejdJBxYL3xknIoSAR99DTm+6i/
SVlVOtfiq5lmcMPBCMXqDEAz26vHn7YiOAhB1wR0ioTgVen02UHptNvG1vv0oToK
U5rPeHtCWSECgvQwstXXGSeQWtRTBIaaxWIW4DgRlBderlrpBwSihhJYUVeS/q0v
nj6Sg02sPzWoIm6JbhLpW8+LsUA1xtgUs+Gq3BlklInh0OLrh/J+qHjBgNsvZ2Le
30ObCzHRZ1m5gW/lh/Lg8o//ty97oY8lcL9CWQFYylml7mPwBHaMmczsxbhlvYw/
azkI5WG3z6ugJcWkYwcxR0/deXqTAZ85m6ai9MHmmbiWKso33sdWL1cbzGd+82aR
3J6hXZywWsTWd/vMYJx9WCl8TZ5ny5aIQULgS8apokv3VrFFM7PgqjUrdSm3fyPd
U7ULvmJZecTFb8LzCzqa/8sigE2b3aDlPvfGlNyTYjuZmFgIz7HuQ/G3ocLocwmR
QAebC7dt4joUjnfbFu6AEu//wlFw6yGrtegWLAtrgivtLNfC8mYOR6nFw1OTGoea
Vd+dtPGFiGtgUmYP1KPcxVWcl9H2Wqj0y8FXE7tIDQ5UEugx+ga+HsJPewvf3Jij
Mq4OOPAQa2ARKI/ss4IDDoRm97y17BgIeMdOi44OD84sRk/Gyb6mflkw3jcPT9vY
pq+IYgrKfHS/hjjv5St68PoU/IGk14Q4RjsnMPaYZkay1Dk4YKzFJ/AgvLgSwrOy
t+5vwf9Vs0OBpd/cIY1MGo6Axl2ovhJHZ0jXUd2BmkPt722+4GnDV9JU8pVOdiPC
Z2oFCN8uHrKbP/2AJLuW0nCteWpGJ42zHJy8giRPQlUPKbtKfJhqawhK5v4FJpYA
a7uWfAXhux6FSkmrzTuU2mW52rLH0nPcZfhhVqNJgDLBC6zTI0kMnc6Yp1nMoqve
GherFoaSXhiJhCToQQV3UMCAi9cSdbmfUYQf/1xwZOCFVB8TgL+b2lyLXrLOodJ2
EAaibR8tx78g7y1rzDfhp/96sWaaNdJkOmgTJvGTcVbIhXb0SYlVQ1PCs7AA8MEP
8Skdta5YqgaR+em7hOO1nynAIAdNecWZ8naXsIwFpKW6UGkYmMB6iTynWuZvS6xG
/JYaDSbhBLZqo8PXO8LOP860o7nicmZ1r7Wob7LobbRrgCGsqCqNXaxqPGuiUldg
Ix8uyuIbWkMOImeAx1w97r7T9uaEYA0HkjZDcPrmv1BH3+baldJHGhZRxEqZpCoP
jQF83jHdYSd5Ajbce3E6FUh/JeufmaOZvqPsxCgD/yGBX87m/tV1p7W5IPKWio/C
sPJfZXigTAGL1zGWLNsIjH+0S15k/xh+jJdS2VWwST62WVvn9dvKsqNj+dr2h+4t
8+fbPuAFz6gAtPTpKety0SNr4RnmklXv4PlhZHoKeG2MXnTDgfvJWYYtaOoB++G6
PBc8qh94CHF7KIteS8+z3EG9Ru/PM+zhg0Y30PRn8zwXZvnID7kABxi3x3pip5ti
vfJft0aRrzO812jScL7nchIcst1bFvHV814AtZGkaZIWPk+kTm/I9OWKaTRoa3c4
gE9l6VRiakYZu69RPvwO3V3b/oX9wDSERP07NWMQ4KZcFSEJFAbXjDN7mAWH9BQF
YmHU5j5s0elFzmZ3XQbx79M9CQJLMzAUhjAqKly++LR9GFlqtV9eMdD/HAaRyzjD
Mi+eT8VsLKBGN6bzkAa1pdefKRAuHoy28Ph65YIw9RZeG8BSXbRYli15SZ8a0Go6
Zlpvun5J7+tq1FsYVxYJnROLM0BgY/aByxT4s06LnldmhQChAzVP+k2Tz+bAkpmr
kJBl3yGu0wwOFkSC3iGvMVA7zgRln6/s9KFsfR/7sHJM2n/zvvQYH4UN+waF44m8
EvQ4RKcKV1+wSewZXtcSMZDfA64MAEc32E3WIz0TTjyyUTKYKrj+GrMcC2Tr3+7i
oCmYNOMKyluwOGW5h0WtOXDkyX4x4CP5eHzrNZ8FfIZAIBlhivm4E8Pw/9iDsnQb
8k1/OHGAmWIXlazUilTdMwD9Yo/yqGvySnXbVr2iNavDMm3Kxmr27H51y4nCoRSx
0XlIpVWoMrGHkMSeKMkZJqOb7B32YwrI923s3l5Dx93SRvBLoYHBuDCWyt/irylf
CDrebQRMPiwwJ4/mgDKTCl84F48eHcrXgmZaljy/Ekfy+mpB+qLU8SdzKd5Yikcg
r+EG/wHLuAjM3vHaI/Z0wxsqBvJ152WrSJMe8Q6CqosdYitat6CqcauuKJ2gdLUA
dlLb8LtGsGeBih1hAztHtYBO0HKzEtKNXxhF/mjzQiUN2a3QBatLHyMIvbH6+FuJ
twEdDphS+qRItUR+aTH/s/JQEkwBZctVbq/A+Nf/NWkcZvORjWNdnzaLdTIMTCxh
IlQYhvbErE6i6cgRvNgoHfjgLbrgIYGngrwyQ0kydmbD21v/p43ND7rmeJ5tybIT
hXu4F+uHFPgwNjAPigPT37loWL+B/Lt8Ws3DoPhpLdii7QvOd+NFByXG2oX31lGE
yAbjipFEUntC1Mjz8KdzAQzdkT4vCoW/FIGU0dd1GmFZOGLuzrxY6jQQL24MzcTY
iRXkF/Av7KNSVz+n9QklM9KSBuKHsDkzWUId7QGyaq/hCxa+9uBPpcmEjBD/LirW
lbbhVakLwUVgwYQswKDn4Df0g3ELvaMT3BUTuc0Jxe+B3mbieu2Y/Y52Fzv3NNLy
KicD3y+zJA7IYEux+/mapUFWT52XdYN4cTBil7GQbWgoAdFa6Y4RB2wvK2hBiH9I
dQPOs8yZ6Tn4XPFzKH1FB54LJ6c6K222EMlkO8jgVBmCbeoDHCgvpCFQQVFAqW4m
MCoEM2tnLHhvkbW1iFA+D23xGNdSH00zs1omwBOV+93d3VTHIeNTGTibc4D0bzU7
Is+sURizyudFNcXzU5gKFdpsm+iyWCA2B8hR9I4wQrv5vLFIW7nMrBxDD2ksYlHF
zO9dmVsmjg5vtcG2rZmOPZnDQQsk2B22rv/J3jKl/c3QOMbdbwclY+emh7+t8iFZ
B2RO7T6UR667eKs5IjNs44Wqgs0BIWsvJDkuYKWNMtabL/KMHNueSIeEW0E/1PuX
/zU58ScxmtsW2P6GORvh0qrCcs26oFwa5YWcJK4zjudwzHJiD/621PyLaaDNdw4a
kOf/RqAfMPIAnmRa1eDYtGOTzplWE0OAi1+S45JOW8FfkJBJP4FaH5tC0mW2PtrC
BvzZXCqtYdeHKIBe7nK9R2CFTLc37yTmw4OnzjOerU3iywQgAk+8I1KwS1E133R7
dwzJ6/7cp91Io7b28KC/THMf5raS+qmJcYxpIPmC+F5WyiiTMYhXEIK65CtomWVn
tDxO2ww6oMITljmTtiNZOq1iPauKA00Q4RR9rLuWOXu9WYB7CPDut04uJFWa+gCj
NDF7ycOUzVdKP2eaZW0y4+VAbzCox+gSad0O4Bw5nWFvbPQ3tGsy+RPh8Ztnm9Wv
v4Ip2uJR3Ti/yFk5QLD9Wa6cVTt92rxwro1NkPViYcsvCxEl3VdRUREpg/tw4kMf
61k1Brp96K0ZRVb2IZandz/S6Wvzg2ETCzHE9QF+hHY08Qx2CRbpvroqSYm3Vk0d
W8+6t8k3y6tLK/Dij+KvuZlO8N3VHuVsA3ZV4JfT7nTI/9dEmXR1rPzXNqLTcfDb
OWc74z8PPUKrL1foU4JIGdTRhAGS8C3QqdjbFQvDCHWW5kItbUdig7cl19jUAAt1
4923s4G/1kXMBpgfjCd3scFyodFYZSIz3t/ccJ0JxIakbQEZOP4rEUoh/4kiE8vJ
3mGrqRDM6Wljrymi7pofizJ0FilQb4eQBdp6t7mKgFyFa4ePdjcJSQkAMFWnEfu6
tEZZzbrLRYYSixAM0TVe37HUYsv4q66vhnPIibWlC3j3v4FMtN4NFFrG19QH0bT4
F/rGGQWZCjX7gly850x46ms/4CJPP6K69SV1kkUj71Ly30QjDyko25JPUy8lzUzD
LN1+uaKcfMdMcD0qulUuFPHApaacEEVL0s4YtyUrOquadhxhHwe2s+3n070UYAum
TWyqyAzwboMTx54s6dYepr27Cf2+GMmBHgyrJwSnh3UoLgvap3t0IRlXA91UtxuI
p9+TymozdPgsI9xHGbAuAzqSMmCndhnDuyRC3pG5M5vwnodALLpgFCXxerJKBvMe
XE38Q52fKwRCpiZ4jXh/Qk6jw+AGKEG/cT+lITqR5iLXXrT/y8tj3+oamKOgl6P1
o1ngsqhFbr1G1bii7lAoVHnQgNcVCmeqWgW8Y3vPMSjL5Cz0jyRdr4LiNns40I3d
kFlho0OlFY4aBANyFpudX3kWwv2ndJGhcuyjKtuHaEXyRW6/vQWQsks+xJYt9gAE
Rg0PpIwvAlRbhP+++XiLoD4stxhCpE3pUpx5UpHgFElK6P741LAcviJbEqaSU/BE
QppqYhHT5Vdyr1w0IrUr65I1JUOdCYNcl9iq7vZPcmioSqqZuoJimbXnN0RsxNTL
GLpeTMgYvlK0ihEOl0T8VH6Dn5dNxr/O2pEV9wyQaOi5v6lW/BezU8DMszF2rhb+
nZbH/bolD6vI3inM8xlPTdYL9K4EFFObNxNMutObbxv7lIzDBVo/Au0nc1a0tWoK
RRsR+lal5UeFWBG7CRHn1vST3dcElDu+kd1CUMJfOQTncb0lCCQMBjxmfHFKZnx8
kRmfl8fd2tZpyCPSGiFGfBTo39YLRSekWtV/yw71rqhxshQoyOu3KePd8l2jMkpY
HBKK+YNuJmLPQIYUr9e5IEXhmw6y+bsl5Qx3BxaSBUgSqft0u08bMV5us8rhj/Jm
GcYYd3qYJXzDy+mNAVTGxi3zLrq1Z7tJF5eR3oVllDcZ/8zrJIVRgdsQOqYkI5AO
N8mWV8mAJuvqlTxiRkWhUIZ2xFyOdj1cLVtG20HnKiSZKh/CbzIXbRiM7A+GUylY
MZ6I2tTF2jbF69U4af+Q8VlHvaNc2qpqZb7lodAFvm2IuViBfbE49omHpa5kEZXd
0asH4GbDHTyHxuJeVEEUdG2gz5G/GYM31B1H9HxxruNoWSeikJ7T6Yrq8Heog/KO
RQML5U2Q5o5zzcXRgGiC7pm7tSTLDi4mWB8IYWcVUZwI5SAnuFObtX6FhF/v3jJz
h5jGKYaI/I6QS58/HcbDI9fALT8F4EwiIcsVsRz5Cv1eZ1p0VMT4mhLhpl1u1eYF
y/Ab2mofLeSTePKZnM1t2c2GAxx1/eaLyFkDXaEqM1R2H5ukLHViObI7D0oh2YL8
6ICBEZfivueCa2AhSgQ5h6Pf6KmU6VPzMnK546qR3OredjA9ykAggjI/nKMhZZvb
CSBRKVXIccS8685CslDGZgGjvyJxQaNVrsnfSiYynKLj3AB9Dq56wy366hyvMiV8
ZPdYWkthEWC0/zOSbQXbYhxBy3tgubXKleWsloVa7CZTygrS+lHfX7mz3+w9AboO
DNftH/cT9k2L+R36z4Mhh+69+w3UfLEe+0r+M9YKZ3gfVJTUWAh9AT6ZLQZIJ54b
iiNxrdFMn0B5pULpj0UqTmkmYAO2e+uCl0eSSPPBFxGBM39B+Rb89uZiw21VntHj
hGnwGZdzazLgiD9nX02SVeztsJJXM9R2NK1bTACUtjGR2dKutirMK3HyVfamVrQA
ekWmLZpmEdlD/M6ZtSFSr0J/kJezHm9eeGh1/TOud7OBmSf6+H0FmqBNtRNkzaZP
CPTQn9z/uQErtVCG0oF5ocNOdC4sg/nlEplm9D2Qae58aY5/uJ69jL1JcfasTLfS
2KveEBuzXXSBZkb5E/G6fzYux8IS2QtdwA0gvf+1AxxpaJxJ/0ReGN4qVCPpRFzq
NnngMEILoAO3PatJxKseyypIcbFMIfxXGpBO6gPOzlZshYHvCxx1VeP9AXLn6GX/
/cmd+au2NasbfAJ2+P7D6aMFz2xGgdnQ7/Pw7uXzmTcvY+yr0v4DJq78sdp9U/kA
CC/0kadb47Cm/ShqK6w6Vws21PWptOiyC/zNuUhaoHbPZ2qnKcHl6qDUI7abOjhu
7wGARfV0EM1gNO2JD8cMGLhTmXhlkTvYP+4m3wj2bZzhq3FsHCwfr0Zhixd6VQes
IdQ12+C4KomVtMcxu/yNvIxYFO4lPDKdN9QDF6dHtnydR76Te0vZ6VKOnYW2tO1A
dNZLIxmpw/WC/CUVXkhPl/J2EY+vQ5BgBQIL4CG/YT9x0b8Q/yAmYlMnHBJHGrig
4D4IKjgkoytr0Ua9jDdhJ/VG57YzY5dRCT0pWrXdp1GkA8q9/fYJlpEA7fNcgLx3
DI3KXmPteH9rIJMAegpZWeimaHH4a9uQc65WbAmCHeRy1M64Cxu1B16fr5YZzkfM
lKqSiUiaTjYMpD+34Fn+GLiQk/Xq1m+s5Wf0Y2HtQC0HliXvtuHuqGCZ+ygHKmrt
jtjCjPDEVYrvXzz7vyPIVGPe+OaA4Bhpwyu4ejnvw+X3oNEYoUkUDeat7w6gXOTD
KVF6/SJVCfhmc3d6iaLv4aQRcpXUOlWkoydZKFbcFVtrppttiAW9wViJC82PU5V5
eu+yC69Mr0GBWIptd9JWLWXHoBMBz/MTfghH5N+C1AjUWcVSr/pjN8bGFUl6TzYD
rO/78N10Lso6GqeOHGrOqxNkYEC4Rq4Mo5iSw3of1VPU1uznm/GcAbEbWq//UI6Z
pKoZcpIhv+O8g9Rle/mWW2euRz5nLT0GBXhETqakQ2YcT3yrJqSqNOQ3d+wKDxMW
ASr/vLuDSaz0LwcwXYXxLUvLrtq4oCPum0HvQnYKl4iotP+3r4Bwge4QX0nQ7jAU
WSgh4D3gUh2feN7RS/jiYKnIg8LahP1fJTOByfBfZCsrsSbKv+E2WKD0rp7vvxsN
vgisxTfTzW+8SXcfIsFM3iR4EVu6iq4mv/ZXHXSwyXjpvmFhCAUSuC6jZJXC7IEE
mw2dNoOqYKeapCcuolm766sTh9TQbX91CFOjT2bhTOfbby12DxG/ISfsr3U4Gea+
68qhiZnzNJtfEgincAcApcFOP6tWVQrYosrJXLJPk6i+OojDNsgXVX9mUHfA1F2o
xFN8VQInKETA5KvM3rDuzik86ltAol440peA2Kz04M2PjHZAyv/dFCbr/zJ0knwT
yHxjbF7G7G4Lz6HPCUPDDSD6ggf4e5f+P7tfHpX4HR/nU0B8V/GWWy9SojUZwSfz
OgRSUNcNCZ5c1rFHA+gu8Q+gt8wldgdngm4L/CbF3ZsiWxUYnEyVuLnfJ4X6+Nkj
mOhdA2lBVMtN9t14J8k8DL4n3AsGOJRFNyTrZmBuiXByt7hN68JLrq8wHhCJ+SLq
7olc3I6pDilXWbppQG84DiiKyMIB2HpgR2fGu8bTvoXZ+pFRfD1t669NaLV/b/UF
uAdQCiNs856Pys6ErhUOhMjzQv/CIJUwRqYu9q64L2hri1Bglq6XoPNHvyDhgowk
5KjZL2XAfq/QmIPs7noaY8I7f8wB7gz/+s5cdsVM67/sfs4rVuC0lGbF8Bapryz4
WC4aRv0Ue9ASEwPCcob9Q8Dsg6oRaqhrdZevittDQWrk4RxAYGtnQfQdX4qscLQm
DW2YPvAWzoQJNzhtKbGwuoG14OyYwycSU1EloL39SCama87V5tQrsqCy3mGGk8IS
B5BBmkx9G3Pm7eYZe/NUmTMf6A6u4A6riZXD28qant4/aUgorzJYft/j/ZNJTVll
G3S8CTkl5Tc6cDP1yBnode4xRtv/m8Jf+fbFzdTFFtYc+RFw/Xy06eCThx6cRGlF
1P+lBvPP5lvMx5xRv+N1ihpysVEmY4wCHoOWztIBWT3OICw7q4+TrSwEE+qGz/b3
UeJyykoxth+G41tBnUiESxrlctKwMqUouyjK5rzCQIM7l8mt/UtP74LOsltcQbQ3
mx1XMzLKN1WrKK7wWVZRdHEEEnTVcF46eL9Hadk17QheGwGUNF8Mc7mZmjqSwRV8
4loqjY9Hvr2xHj/Mc+mkd2844oLJqfrVlShzk9ibpI4k0TXiH4uY2Pz42ehPxDNE
FkUpRtXNy8f9+eNqlhdA8M8NIe9svyzBxqCs+qB/UnqTLXgFxJ8CW4cmIKhJRB41
WvJIRGGKrnIJvl3iJKoEqfuCA+CANq3CliL8i7+vSSywa7PszduDX8CysdPU3aEh
OftAFNKzrr+eIADefSLNXrVN+8nkGtJ9WRphNbbutePJqzaA6r1Qrtti3mSJA6cu
rUlxpitJLT9405mKZ+JnJoIyqHdKEPrUmCxNCqN2zpxy9ptjgToGzwZ42fxUiAOB
peIuNWbvMEFZ1cy4eLyKIPLniB7Tz83bVNP5BbBINeG8EDk64+m1K0RjOrttZo+S
/q9AvcSb8mRlhe4u2kHvyW4a1IlfV/27YJSNdwmBRRdRfAwcXVm1m0PSw/lx/oes
h+wnZT7pSC3zho+3/xDcJARVAO/276iy2Vz+UFcqfM33ypy5TyHnNwGUIOTqLqMP
i7JKUTNj+cUzPJXQfUwNMb8IZ1zlZ3Rnu3UlAsJsQaNa2IUoG0CvCIeNOe1BJMXr
/l0ynbEBge3fhUNaofQzWKTEUetgYlT6kAszORvg8slIGqYHa7Df5/6ygiBhvXo5
Ia4PGNk96lMxGiKTxRaT1epXMw3hwiF0e9/lX4TKSmutbgWtR+K8hLuDQqvIIaSm
QrL0u3LPNgYm3BwutV8Tiqrr6Ezaua7oA5p8f4d9pYngbkA2L+DPl01G3YrQ4cyw
aepsajp9jF3ocFYvhjmsLQ8QdgPBnMPXfq5LK111UVKskUsbgt2+fHoWK/3dKkvd
QFPmh/EW7httc/Rw96JvcyO2OrIyNVbmPDG4jL0qW1u6a2Am5mozXPh3ELo7WvKt
wjIU+3Z3F/kY92uWHSgeJg66cu34HeOBVwUEPLjib+IIHQ3NzMxtdKj7NzCsr0nO
tYl7p4TC7bFp5+sb6UIcKGq32/t+6T6+W9anEu5w9iXFy0qcse+aJW2Di3BR4eBH
da89SHTq4cAjAfCzHkUEykl3Di53fsSEpWrZeA+j8GQoXHP2xDtqw7tOExGC6K7b
Nbe5n38YVhc+V1pSqfOARHSBL7kbI7+WIHhmvzkEXi4j8x4zmW5BoA0WMskffBH7
4wbOFviMQDgx1iXT896aC9m1p/N/Sz4a+swPGvPyN0/pJ8siJ03qCCWWRrb1iZXs
qZfZvyK03RVjt9YgoZBQ9GotJlQFmA9TdO/qvVWqSl8a4jZtmAYaxRItIwec4AAW
88ALbZ6gfjPaoGZTMI5F4IXJNfXyk+KevQ4cKoqexyp4nnwyeJ+578xmtaicAQfH
9CJy7pffPboLi5APzePVt3fwkyf+BD8jgZ97j0TYRM7hVNsn3nfCAKo80CvAWFAK
H2qhFscCa7itzIfUEAqL9DYRAQT214U5iQUmWlvdMcjN3eIDc/03j1gyknwHlC/K
fyNB5AqZdYfQBlnr3OeWdTe+rLrIP74rHnpdAeMPPXiTyMdMBrWDAUIo4eeE8j4n
fxG+CO+TSSeJGcyuqY8DhrimMZ/7OC9NrHQcp7hB8uJUSqKdJqtVf5NYs5n3yHsq
6K0ktUKEDK2TCv6z8wS/00DID7o0KEqWECCw9wzOc9dTtn3anfJ7RwbYxncsGcrU
31574lEf74OxWf/YUH2AzpJGn4ff7op1xzYQHuT68lAFNDUt0eyqaJcAAuzmJiH6
tHQ/1rn7QbP+HxTMIcWQQ/nat+TmmYWgMy5KwFhK0sDgnXoMsg7SY0hCUB9kNg7F
eEBtm2xsdkbz4eialwblzsFoNF9LHOUiuPl8uob3RwgLtn8piNK0BbbLb7DUwUo3
KnfWN81yiU0i7mivjJfnzYJRY9N2cdg9kbo5GChw7BgQzmlrZeVaY7QYxRk55BWp
L6pPrQ4WCTsruQgqy183E3GMhymVE7PzuICvxEu06bbMd2TOg3k0zpjQ5ROkJxdx
q362p4HqRMc2amofvZ/s1Dg05C/KqEGyqnHnQyiOEA/n+D5t8K/Jahyd8XC37kdL
YSFMChC0KdZwBkLnc5Y8kikobe/KDKpKETEEUj9OeJBRvI6v1baXnMnTxiH04JwN
2/4XG9xlN92gtrASD8kXImQb1nGJ7h9AM8lFDBFHtw8Nd7EoF4CCd4Qll1sJhx5T
hcHCLwjBdzIrtyi5CzJwc0FYuRvhGKXTWwBE7fkQcooED0NadJyRnxfG6eZMD/c6
4HmGMpsLPbUGPafbAJP8DeQ2Gx0Q/sUF5rfmBZA1AcensQydgX46YC4VOmHGuotI
PeCz63UECHHsl3TJdUCqDXMlaKgELgo9WI9pSW6Z4WN9UPk/e69EFzbLvg/GASGd
kNywknp0e9VHz9dzflq/FOcCUhzeL7sbQWs4hIiDYEhAOFP6YE/CakO/XmqEqMDP
PN+N7qEmNn1vnHsHiVZ/utwbQHDQ8xqC7NFTUla7x+KuWMt+itUjc3pEN1jjxoLr
fgzxsAY1KmhlZ0QqVqQXZ+E4xEQbFpkb3Kj01CLr9cnzeURqGmLjO0LWIRyaI08F
B05yna+wl+kCoFXEbSaV7Xxl2pI/WLfTbfHAszZaV0+L/QoHzp937yP6zpU2FeI2
F52V5PUcsJy17ekHdQGMKsJg1Thp8JgdGRSsNZ4qSTknDb+Co00Z3A30+UUBKoRb
0A9SiYLKpWKUJZ9r4Urjl2i3b7ey6UOi76qiFjSR1InY+aa4+VR2R7wnCuBp1KHN
2izfeiV2IW6BZ37f02ZZr9AvbxtNlkbLScOWT3cLX9cIZUlnq4OQOB1C9Rf8xRFP
C7o8pZjMJ+Am6JtK8+IDy3EZmANe+7nomH8KVVZuspWi3XxLjauj83MXDtgmo/XJ
LFO5IXKFyYKBE2n6IoV0v0JHrNTW2fFE2yXXIzoXCTnlvT+yq7xnunn7HlCxZCgz
1sQKqLcYYP+XCY9rDdt6XShLXvv3MqDqfCa05nou4tzFhBNHB2eeZLcwb+SS4Jn8
HInJbVGSj201Wt9ri0N1IEj8zGIwooR1MB3EQwy2Dw68sqEDxWDCaVFCQW0NX3Ei
iqBokyDuG2NzPuOCo8Qw5oqN6sHBjARONkn6frq5pK8Ubczpl0hNKSOor4vMdlRt
d/7y4tlRnbiuif/55nWeWo+zzZmnPAvscvbRNqynp6sRtjBxkaPL0XCjWmU+9SJn
sNBu/hhmHcDoReK0+l8kDxdHAJPLZGFBg6hYkIUtV5f4y4VlxxMRS0Ov/eOCmNY/
BowmQzw+niIxEwMZCOeHUbAy1Mkt7LZ9vkwR2sGS+29N9eOE1S0bR2JnflDHYMW7
L7R84ReW7gIzMc6QW9ta6kBsiULzYEVm8qG5+/DRrEZlq4FQEevX/+MT5noYFO8P
VLmpYr97aJuvgHn/LOC4B4C040JSIrR4hjxe+PirgTVpv+G75rBb9oTr3jaQ5yUW
WhX5KQV0EyyNULLusqpe/6Dhw97Xa5/Y0Jo9rMUpYEPHA9uzeuDhGbdUw+K/SJ+d
7xy+3ofBe4YFj36MWhPG5IG4B9UhFWfd09EoQKWVie30kcrFh3dF8/TTTawkkq0p
BHBdRawdm/ToH18F7+4PUSwwYe+Djfs88J1EwTvCmhw1nJ7OLprHu8b7czC7H0Yf
apYGIe11xcBvrbRwlROnLPsqiNLoayKiCA64FFdNJtdUeWRSeVzrcElkzeASK4i0
Ab0kdd0mow/C2wr7SdklX9KOTtsznjtDGUpSUhopJZmki8q5ilqDEyulwoNvgu7G
5Fu+1XwB+IuqdaCCyxiS5oBnWjIEhw05O4cLqkL3vU5fJ3w6QANlu3MBUIxfxEZ0
bBYlydVwMdx+9MTNxiz5ju+1a85YuvQyn3kzAgOC7YWW8Q2V4zDOeKvBfdcIVnKy
RioLlsnuRk5mQBRcO45VtpR4oPBXKyWLdXVlgGLtkqen5ZABlzdCNn9q1x8vl8kc
C0xMNeOzQQrc/HGPUd+hUest3Rv4j/SyncQM3iW34wzV6i8uDn5vumGrZDDtnljB
yC9QKvy4rJbrlQXOR4JjyhdWaXjf+/e7J2CtCPzvm2e+WpwrLkw83umjMiznYcpq
/3i/QKjg0mSc/QqU60CjBiL8/UjR1bDKZa4V+fpw88BRLn0rJEYyItSGqb6jOWEk
FXpgi0C3qofQa+p7CvbIDbOd/R9BU8GDvMisxfDWX9dSfANzwLWHEgCH8wqtVkRh
kbzuP+XXT0CxXyIuPQkBQi0ogQrMEjaf2d9L8oufk1CukisgLyvQn5/0emwq8z+x
/fhgCkv+Y4CNpyni7WPSvpkAroYvIcAJlWHBo2Rv3fBRVtGpYCIxKXDc+UhpmzDn
cDterYV6oW3AdD2nAvweIy4P0J4B2XAbFGwrxphTkYP1CV/t4h9v3BC+sMTQmq0K
3SX/RmasjtXGzIwjJODYD4k1S8nfCAMhZGh4ReckbTTGU3j+qp6TA08nTX8F22AF
m+kT0BZSGq/SfKQwMvuYMy+sGO1uxdGnA+CCCAGiDyQ74wsPetSjrl0hnCtpqDQn
6JRqO9UIGNiAkjHHZC7HxTJy+5T0kfY9xeNog16R/8S90esySHUHQ/sCCpNkqMRd
T3WHEXKmeo3inXAyI6Ht6+UksnRlCrrykhMd65w+IZbDS4Fyx6zl9VvBDV9nNOfz
gpXoO/kN+ji6B3fY3Y2mqW0Oz7r+SdC7eNK4yeVOODaauaUb9Fd/Hh/ZyIsNiUj7
EQIFgFv994jz2qr+cwXZ6Lrohk4XYg5vp6ePe+UKFK1oHw+XdCKe24cXIyleQRff
rdlJ59RyhqY6X3UlU+kixM0a7oaNK06Lpg7p9H0wrYdBcOhKTIQQ+0Usw4meVX5k
J5tD9nDyvOk5NfAGSjFJuxWCiDotCvidvIhiMJCtQ665FzYe4DHda/GZGV/Y1I8Z
DnIXhXOVyiZngQzhRpjk5juHQBy8Ba3UjIRZbXqByhCElZxlf0L34zZOpfD+f+Pk
jRsRItvkLYvKTeSbG7ALpS7L7AqmDTPNDlqvYi9HmM3Lg9a+szopAHQBG+yMANnT
AlxTU1fhBDs4wez6rbNetAVlBAd4V7tUTL6gyo8FWnrKk1hzT8p+2t69NWWkLTpx
R6wWXmW8eFxq0tsdgWfxmDBoUIvcSsmdbvM5TQk5N0rVlanCl+ci2nTpdApk7bpK
7dVihCVON3dj2iayu2sD1FXvzEkLuLSMQfxkb4/RcyLhlhFidWx7qrIvRPU4NZ2a
y1GCs0vHisDqfF2Vs5W5K6GKMC0l+u8s+fKYfawocc6kPlcB3U4vY4LGI3TCF4r5
fPqgSvBTC3yA5LIySqmh2VEVozg0tckXLPzEupwMiaQUsIKhvGYSCcQb1bf45sGm
gk+qOxLpQ/EI0iARUElffC62uzr0W2toxDit8vczASlwXanFeaPod82OtZ/LnXE7
SOzWWobextQ015svJi5mQVH98aV1u9FDvoPHiGdeFA6cgBev38NueKo5FKXlCXfO
lqmuaPnxKeeUEqicQ2ImooqjejtOv6Q7fuL2xXGNwbUCM9QY8W0Cg/t2p4jGbuZV
MYdVUp1fmK6RrnVwDfgpfpj7xKrk829G2vz3CO6EcSrMIC0IfxYFNPyNBfhr4aim
dCVQnrQ5kzr5WsBpxepPnFDjkZeXXPHzSP/0KJCQlqkegoQodWjxxe0YlpioTa5Y
c6nH5EMFnyKUs9VJIdEpdskgt6qgE++KvuHGyHZSsRkIVQJs0TXclFWc93Ilenkq
+nRcsDxiJ5ok+wv30JP+BexRHDUJruDIRiE9BOFBtSozSRYBU+1kuODPa3sG1aGO
HN4GpwQ+O6hTUx3RYZid0NoCF/CLtg38qY3LKzGEDpEcR+NMKW45gsnmRY5276/X
J6sfiQtu+k4tbCDMlwyIwBSvDzj/XfBksXZHK2B0btHlvLVmXqyPrUqInnNCFN9x
bbTikYEOp1bjOXugY/zKFDcjMxw4NRIttmFBXST7Dx5fYCZhaw5d/QpxJUMmue5/
h54qDeRP4xjL7vPeoZWCeJ62QI9MAlLLLZaXpDy6LcjTBodwoAfT8Aijm1uqNS+b
+P52C+8elCUZX3gMn4ximNZwzSpVRFXfDeEhONjaO25O3c9eqhKg8HYmRfRbfO5p
Iy2Dc+J1iz4ZS647mL14OA3CRylk3wxw3+VYSeU6W/oR7K2LQJ9ZcXM5XVGNTp9A
iXaANmLgHsO6dLvLntJN3Ou/7GxkHfUlY85m7413Igz5yCUKrv1NBhhDBUNuZTq4
EbSEIEyMFXRprbcy8UpeaUZSNHb/woCtFNuwBepL+1SbztOh3wOgiuz/9jiMcGs/
GE/sL/PqCUXnrCJzUEPnyI/IRLPVcoePFOjIj472Q3dn29sBTCzDoBX/Y0hS0JvY
lNg7bE4s8AJxLmaDuruE7E/mfUE09h62SFD7DY+yZhRCl7yt3h1uI1pRGRghUUa0
GOvMTerITAStWN7o1Ji0zK9wyElUI5mFoCP9kg0HavNyU5RE87l4Bf6f+f2pKpf4
R1gsG97g2xoOJ/93nQEftrNK6FrkFi9RvmumFx71AnRI89GZItb26lMBQw1v3bgU
YesD9qB44YB35l1gtU3czcOXH6qKsoXEMZPMjxKWe5YD4ZpQpBIROVkuyVO4QNCI
DBhYbIpVapBJvuv9dxLl64qA6UEOUOEi7X9p70gJ17N80xQ7Mg09ZOVdNv73p+Mb
KxnQjxOnGexZfw+WYB/ipAVNdgBfHu2zoqs3cPBdhqCNJpXahEaC6iyLs13qMufN
QRbN3NpFiJHkGhqLnd80A6OE2WNzdOGk6cNvY5puR+b2iPtDz2iMMhM9OeLmoB8c
YujpGv7joav1o6LJtlw3rZZ11ule9Hq044RRfnBa/bdIp4rCdAoSdjaNLCPSHUmJ
len2wvDcQqbsWcd6FosVdVMFG9apYXX0W/fYiIRvTqdCCuMWEaIADMxlu3lWF+LB
3p69+g9Y8tDqKMw0gnp08ZM8vrRKYF8vtMdaGy82yMDx72CNIfNqsVjkwYOUg++F
pBB9XWPGGyL2yyF/aPYpul79sCsT5Z/hbooBWQtE6hMi+9pTEgYKaZgn10RuxolM
QjK/ocfVUmOtJr1YpxGHp4mlXuFRRiTjNsM+a8ccSx8nAlSsQ9Y3W/PaT4ZZMNqi
da3gTxrLCS7OxqzobV6rPrOGGoGKphlZexmT7fRMVxUSEgabKaRMnirWXUmcsIIN
f//Mgk523nkqZvby8M3IqjDLc2sYnHBydsBevGwdcpBTtxznhKtI7BHv4Rr5m2XI
u09sNVC/vjbuMvD82VTbDEn0pauoWe2UhRNlGIt8L9vwHOp4unmWokRD7s5DNAY6
2NmA/dUpRfyhUg7MB5hDFgsB0Q42D0hKTRA2eyxUHsGT5uYkFy0yWtsW+UM77fLU
PqAHhUXCYwGtcE/Z56o+VgVuzU/+O9UPrT/tUrlAqL55mj/28uUHAof0GeQngopn
I2wzKBjJadAa3g9lmxA62YPXnXFcu2EIMfD4cZGMutc0JYcTolRahEi081hGlizs
ZUgznKdjgRDY9ncPxEV8hQl/8krDznR9cvJTJYmoG9/tunwJ40Ufr8ft76/4T9l7
w2tlpFZ8lypSMAi+3oc78LgxpPSDf0HJm8mbVKt96pXt43IuVq+nGmAai9kAQVBU
XKwN+vcJOvHNX6Z7bnyx0ubLp7C9auepKNKLxclox8POUSSf2HBSqyzLXNk20oZv
a+robcIJH+JOWyrCEpB6q0SRu2F04V45EKoBHnzGZpzslXroLIBBX3EAO2WdkIn4
FzKkT7MyPLfQADpOM1P68NmojBza48CTO1guYF+ufr7mPyZMMJEpXt1UkzP57amm
2u0ontMRf1hiHhgkBAFwHTKFVJyzpui+FGEr4zH1fz33v278GcaQwMz+VhGmGzs8
Tij30Ud1+P4ztMhKwGLzdXlkCJloypOYVIMSEV9zZSP6bOomzmS8z2z6zi4HKCIn
u4p/pw8YrwxAyG0Kiw3pQbse9ydM8tK40pJlaiKP+nj0Fubm0XtaL0DDrHSCcCUp
Pbca8qDnGbRl5SvofJHWFg9h5pM4qQSNc5Q6Q+r2tfTTcxPM2tvaEan4RUoCa+jJ
OlylI5sDq/y3YvkPH90ERytcOyIBp4Pf+lBtUp5OXkIh0GeUite7vETXrpLSXvZv
WfIFP1WWZs/UPAmb9CGpBLXSdDAjeIEFUZ7aROeEQgzcwy2OBElwksKULT3vH0zT
5Z71iLUiNnBhQFU5BDCDp2dvhje2KRRmKcN4IK/7W80diKgqQy2K5cuaatthfneG
9+NDm7ZetMDtRAh9Ja1G2zp5sLyKjxCH7PN3iGbOJCLb5v9eUsCxow0XM2m/IIRY
2lE5s0qUmIfLtXJsqdsBh44MpPMlCKX0TSMMEmDyNDvFSm972uObG39kPJ2MtFyv
Ox4511kIHXxexZfXxPMS8xuZN+TCSWGNr9RXFnkkMbAx/g12UocDDUd4JyO2nOS9
epqGp3cC8+MojlUALnzizPwHRRzCG9mkk24UkIX8+ihSguqSJjPVA5iKVS2teS8I
qtLfTWchQAa0ffaoAfjCh/yZ+m8Yowvwjvfa6hWDGLa2rVaJmv3ZrcFXDQGBUunm
FdOwf7hnv+4DTbBM0vG3ZLDUnqDXfMio52PKNZvmFCJUYYk+yhGDJ4A4+x7T4fkF
bdJnjsTZQnNtlrEI1okgPinmRN9YyHXHuPdPtQI+iVw0tcel3uSuLAyRNyMpWjWk
jFD6O1ZErohRacAXCk0okL2BfxRo5zkLv6/6B1d2g4+//9HWOh4hDizAx/ampcom
4EvYs5P8jAQLcInkVb6GDTlvRfAgctXShw0YdV28Y4h5uESto5rB0j6+jIPgnXoo
zMo+XTROJlSKTofCxCOYBe2Tjjhr5nPMkG4lYy+Aae4wq5ciGE5RrtqOLDbUgEZJ
c1PC2sQRwT0Z//XOLs/acE6Hf0J1gW+Z9Ny/Aq5nY1JRK/sQsWIPgQQjTvgppQ0a
H5kj5t5nq69tEz4Sbpvfv+gOLoJK33xqsAKAo4RJMRDW50wXwpoCr9lyJuBbVqRA
WZNjovfPA30auDVR30PHPUiBN+25s9m6tl/xvqIOIlaOmTWv+pzgio5hD/5z0ETK
y+6BK9aXhRF/HOB/qs079TORFMMfok4IkMKEdCIz6/d2KINucPsaSvYnUePcy3w6
NHApdqTWQ2hF4dqTyy3k/NnLbbonAo29wXE44ULN428yCelm3KXKVgf47P/3AeYG
F0OVdcKtnarY8TlMDKDdgUVB3QtSoy6fxR1KPEgppr7BzoZJR+p9KKwxeynuu+yV
7ZkYmlwJVVX0LPYSWQGtni4Y6fW2FI3DI8zwLJVqYpr/ZTOM/rnBYvO1A2e902R5
hm3lhVoiNJEYcGAlZHccmXlh8oxaWBI0Lb+K5816GIVbnyX6SCm3k2+acOHyKM2O
A7R0O7Yx7A7rNfjD+a9Jy7hJ5JmWJoRCukgWKIeeYpOUtGkaVNztm1UnwAwC4qn6
dbYNgB1g9Yschprzwmqf3eRsYpyQBLv5jitTVNP+RmLFpJtaxr6rmD5EBkiX8KVm
SE1iKQf7DjBQlvuPGJuAqqduwkRlRx3naBMkNwBnq3ECtl1O3aemR9C8yHMpgn0F
LOaeA98euzIlnzqp9T1sTCpVALsuCHWEfysNhMHnyY/sr+5t8gWjcbdW7pxZjDC0
72plFvapqUJgbjIsW36fHYQpH5GQiz7XGjqXcIdc9Fr5sVsCigzNI8rfm5ePWjXx
aJ8mWEhr/VP50rc/n0m8NLjut6wVkEP8/2IPUS28RNmaVh5Ublu6egVaYDjdAid9
1fEX0+07H5yFucFCft9RdLW/JenEoH6s2X8MYbDe8RIfuDm6NPHTmQlzob2x9TEt
+mBU16ckARsZ1RG9z4Xp6Dv0WKc8xFiiq+DGJ/D7RLQge3uvjaOEAWuiEjsLjoTq
Znx9OWAO70KhlnQV1SLdXiQwdLZb9u4iX5IZK18H4cXWeOe4Pw89nlJyZyPehZLK
CZ7NEsuFC9oM+mR3/QbYWORe7xCl69+aSgF0axigAa5Zad8IP26dq1TWZxA0QDmJ
QLN85uOiMnfjMksB8BOfyeJHQFAD9SEihHU/JtHsRNhVlobjhaVfZxOF3RYbZl+L
j7op6PYuTsd7rDV4N9pN/VMHS4oMQHsK4gGFu5+usmh+w8USGcb3pfAZAii0bgb7
GHKe/8supy0eb7gOsUcXd85lEn1CKrOgpoGbGmIOfLp14bZcvk7bKmKifxX2tgMA
RGabJyDAWK0kopktseAkBSjIIrOVC25ftX9gudKUj3GlSEzJTEFzadeRY4CfiZmz
JVrmG/vTEcQn14303cH4lnLz5oAycrx0+mjlV3KgCEw8F1PWNN+hdfwMlDQN+Mg1
FdF49t1vvHL4v7tLTObrVs5+dpAD5AUKc6r64viIDf0nkVeJ/+4EH8fQY9K7z0AS
Bql6WyriPilZ/M82i31YNJUUI+FluIxo56D327cDJH27mAys0ZvJpJTTJ2xEnSn0
St1J6nSqhML+fCrTNwzuFCGULKqjOtDzppGRB5kxQec+FpqmBKNa9MB+ceFvCm3M
ygp0qYI4SiAK95i1V1AbDQ+KSR2ioNX6DZfw+uA2ulqCq126o6VPqtxrW93i8qPU
5VpBoVvNGQbmoVR9UImTGQujyXK3Vw8AouzY/13mWRXIi3GWnNdDH+N7pRDdDZ6u
yN92UiIW8oCnKz2vlArjH/2YyLzg68xmPOkT04XiEQ043DKFQIl8e0JkIdztYPvj
WJPQRqhoIR4IceUejuybIxcBIaXctvjvAVrZee4Aapov1aX5+Lp+dnQtsh9SMVCn
RRG+shXqkcaxHoNSphv62swyCDl+jb9Ml2Zi9Xvwi6uJvT8Z1iOqUUrmXc2ZZEnb
6QNQVkwbJm+zZIOJ4iDRHKT6HkDi5IJMziTYmk4BCHyxrQi3epkRXxOi3g7+PkUp
hev6jwH5eCz1wbXg9sa6GVUpwpQsbO4eLJuVrgrhINTXb5gFzunxvYQqXkF54IYN
+KAOvQWuLK7zc44Z0gUFkheMfYn8gZW9FXvkZkFwgk7fZ7ELU8Wz5EJOH8vKgU33
Rc8Ar0+yeuGCsM7vnpgCXVBAgvEmsCrO5SSunL+u7rSeO+f6b+QhYgE129gG2q6t
evwOHtmc2BpXTMqm382PsJTWztqfS6jh4Y/MVxtQclpq/tW3lpvjJV8/bT/MCceq
1agFM+BhjIflAPOHRbx0T8bFyoiAevXeign0LRKNiOhFt9mrYAaxgbaRHBXCKBs5
7qqAHsGy04r+NNzB06P7WZlerFg5Rk4JZP7E3KiepDtwfjl8kh2dFA8NidiWM05t
+bpP3F+EdWAkLaUfl8FjsTPYcBzLif6Eyede6zoujpoZGU3SRzOqYsyxoLxtahDb
lKqrK2FzolyIzZ5U9U9uePGO7ps4Kr9ypzHjPioLwr7/ldX6Fvp9IcObF8VD8eAk
dKBjcwvszEbTaToYh0HVIy9H6EUg1sj5C2PpU0UbEZMa3TRYvELBRQ6Z7m3E0S9h
DVKsxFx7tMQpkw06P1BYDyuNVa/dXGs4qtBRsiCThRliza+mmqm1ORPkg4Zezj1p
UUjWsmwpRYIo5bFYDJeNa46S+qDkv4OEaiGR1F7KDjgZuDd5p33NvTFMO6ABLyrL
EtFLE06lJustH0IRE48x8/LrA/X0zpAYfz2DKojfBCFBukK02CIr9Gyc7Np0X7UT
rkd5wS4dlbl01DWjKBWcRHtKdnEayyQF/XmlCxx1tPmLF4CH1W6yGhYYAhBwlC6I
bKs5TmiNtgG9t9sb1vVJvq0a/zrTkCWtE/KnajgzirHXgjU+DxOFKCjwGshGJ88a
fyuFOBHKhYuCD3J9emPiKTUE16QCG4Zs2lrqUZWrpqMjrC6ubPIaAV7xXJbqrmTM
w9wd3lc1fWPj1VrJLVkm/tngR3it+QwjPqKimkxbx4MfefMYK3SFzLrBAqK4ZNZz
mi4lGi1ZR5y4VdfY5o85gDyIiSQwIf0LRXnbpigH5u9Iiv0pEWXuw67NAbhojFY2
pVLvfiSVEozJ22S2H9LPghssQ+KRijmtD9KBuxQWORRqkZNw13RzMEwG+fdkImMd
DhSgvo738uRPeLlowtcNxWsSUZohjfUfuYwbcDkTRik0d+tHpxcD742+zN6y0viu
Dyd+JpmgbWNcnzLYMMiTQXekUkTWoEwELqQLK9hVWOgiAOAqygbu12zBT25LtXHj
hZZDmLVc0zMZk1kedE2AApJInTuW0N97iF+WUu6mUW2AiUmrz15gIfbtjQs7TEk5
42yJaKZCK2GfdohaOJRyugZQyY55r1dqmBJgdIeAXaD7hrI+GRoVF6wBSfQkEhkK
WOIjwxUtgrFc+V1lwj5eGu6bS1Mp0XVe+Sd/sdYOztfZ833wO6hyvZvFU0TRWnxh
4Nr/qDtf6aFgR/FhA+06moNEciehKeKypMESjw7/240vKO5TGD9RTvIsizCl5N1s
NVrgYCekwHTHdxCOzOBkIl/5GWlX14YtR6uhnVl1dx12NJl8F+wZdZcWPwoL0Qw8
/5y0eI/P9i1S5q2cxxqZb0oB/Zy6pjWDLvnAdtoqiVI+fp2Qk9/COJuaT5SR01KB
oGGguFwN9JIDsNDySMYZIZ2TUElCf9BQSUTfwp1AUE4NOIoqyDVD14+F45U0cCCY
sVP4E1g33vYh+zb1rD8pwlBFQ7arLnST805gFwqtv3BqcH4Iaa9KetFXzAJ3dhrS
LzlhrzeU8DkGP5xtYEXZ+4d1jXPiRw7pp//LESae8oWZpivqIZ6MuZjQmE9VYJYf
c9R68xALVxwoI0QWj6pA+WiXDHnaV61bSFDO+flVdFu0x0QmXyOMts5lsopjsdkf
LiXs0/VR63LRmPRdqQDdEa01sDsizBt9Ib0jUQXZDLBX7dvdmNT3AtrBCpy8ky+I
2ntGoXfHIngJrHg/Y0Rov4T4dZnekRnkELBu4XTR+UhzpUt38dAyWwt3LKH0N/dm
aJslk2UPrTIpdujl7ScKwQ5Kk6tWGXBkSY7NsyDs/0MWd3JauwPycsDmhL4TY/Ie
xve/9Li8pm95ZAY+kojbeumbWUp0iWRs7vweSuppf476HJ+bmv/SrgJJlm/uigTQ
N0diiiEPghVXOJOxuFDuzyfsnEWlyZLfZp3UOo/VFB4v+vy/1JRYkdxZ8us1cvTv
+f2zbG29nJJ0lUWNUddo87hmVDKBBx1EmODOJLu0QcvUZvsEkKnibyjYrhNzjAnR
GrWQd7jU7G/rKV5PHulMRDyioKir9XhjaftC+cq/yvkURjlJdSm7eGxRMf1rgICi
jfOSBqW4UwAqKMpxB8YlZ01ul43TbWAh9BfkEmUXNPJp/PuTY0Dc0P4JcOxUD69A
bcUBobhWaFAqoy/Z7GvmwpoQxRiTovxtUKOmgMuvesX/TN9JqwfR0aKagl3G/a64
ufEfBc68K0wHJdm7l7KbzlUJWvULaWfbeC00Y2ESwh4RJSl0ITTg7Ssv6YYQMIHH
2hg5nnygo/1aR4bQeQ//lRgY7VNmh9RmTMTlg3dL4MsdRvToPMvmqfyXjJergjPC
NWs3uIJlqcaLRZ2ABpYC7xKC//bvOIJqMeWbzuXFTgitnd9xdAkGCHq6FM3c4CoU
ExBtydRXDDA1Wa3GqCk0Zlq1yvNtZEIrs0vRxqs0hMeBBocaYvrnsawngqzHmKpT
BNptnYJH/z5rO3DzxDGKGGiPw5ZrqtTlp4PsfsfHKlj0+0dz+wMEPU55dsNqD2Ft
DK6kNc1Ioz0UdpbV5Obx+0PKEVHH+dAPLgzo4TBUCccWIQIDMkO5HB6MI5DHkv2D
srAtRzoWpHToFYq7d6vVP+U/od+tzogklVksCU34EVA2JWp6sMEFWvhFkFRoHLmz
5+HVH1HNu7Rm0TuFFe1AILyEI0EDHHs1lkIZoCfMcq5JlI4P0bDCpYSdN2uyR/mp
SkW+GS/a8no1XFa5zdBTktI4oGNdXwnJcwZOB0BjUcDtD6qVw/qjBZSO60h2gKws
wpMyl5MiiD18aSl1EjDltDRiN97bZidIlDVSJNLSiH4jim/sDTLeC7e8N/4KzhBM
CqGxmGIe4RjmDbrVQfEjjgMPHjvtzgoJVTjSrF7esAaq+WA5GwU6SfkSSnFo9SY4
tR11VqY/GSuP5iXEXwmQCgaVSOu6NCPLmGJOlg+08bkJFsjf38AT3wlrKNWjUOhC
JmIT1AfHQrFqBzvUNSZVCGKXuzSnkJEyyGWkxUhWsCPwOaXlfKS3Ij8zy+aB/oU5
REAXSqvC12hT1NWb/btxFL/ywHv3cRHf2F7xVA6nUC+0UiwcmzN13vILCJE2xz7k
+eS0FGW6RljptHsqcHb5rbC+pIGFxBLMgX33Qn4kxJbjRgnPZWzii0EO+Od5cXyj
AA12b0OEdRjuufzWKwTGSQnq7onpfdLE6AUuyO9usnBD6+Fu808alV2nI9FXGhcS
6ZQZZzuh0aT4RUi8G1flJ7bK85EktSnBqZF2m3balnuAwdhSX5p6sZWF6jKGEQO1
DL1+5hOVgjmCgppwxOTlx5MFukXU4cQSxYLcE1SEl52etUTNOT0+sc8arTj3rsDL
YFLZymSmMa+qxtI0k7nNHm++Dj3zs/9X+aAiRxLQWMnUiiaoLkOOdO6xubJupGTI
04FmOwpNo3GL19ltAkuGZk28LNT2FDhGkkIpINnEYnQU2x1IV1M3B9L3vVHkz4TP
hm1vSJqKxIQ/8EowHt5zAcbDdtEuwJeG9rGFnLpuzzy8+c+wS2encjqzBrmKYPYQ
7IPaLRRAJrA/xBKMfAVm0nZ/bWrLgmi0zS4ADl6GyvMyOUvMzsAt63t4cUy1YgE5
V1d0qp+2OglcZnClMAW4UjqSqD6jL5/JCIKtyTkYTXI7U4pE+EITe2g2Hf/ovWo6
9adQF0XMxSAGxAGZK9c/JQMIu9c8FzcKxq/OTRLTzVHP6lzwspeujcZ+wbrI1gR/
3P6V+0mQrxdPi9sDJ5FKATdNIaFMGHi3Xxf8/tlDwKVAhIIUs0pxjBV2MrAq1AJ9
M9UumXr/Q4Qm6Do3ZjjqZwiAnJOd2DPy6NCZH68zGMQl5NULgw34tIO6M7nCSZmb
Cwxpm6su8LgKAGtF+3PdnutEhiUIf+J9YdR2Tq0wtAzspchW+NMVAcu0LU+Mpin0
ya/tDIeMq+L+b/Yv9v9C9VKrEYLEk7kuFHjETgR5mEuOel8x5AzsOAMaPYWEKsn9
NwujwRpOFXPoa/woH9uU4FBj4uS3NIRQK9EjrEpj6woAOJMuPqUfmkc3yJRzCIqB
ZqydobCcHva6kY+o2Uyiol2p+n8IDr0vrg9z1cKibKzMSCbVabWdSIEKkG4tKu1C
HG1HgIqw2LcbAVaD/1GDzoDuT9Z3G8Ldc9iSfm5whR6uIEfOB0GpQEITy60YfRT5
y5k1tK+wbsyo2m5car9xB8M3u43/qPcNNKZLXOzzKZrQa2O2nYbYer68qsyFobAJ
lEXN4e04YojoKMsSAqoAFJe2ZTTDhTklT8NVGqEp+ojNiBjbqZPy2DzY2F0ayYTa
wuvtvZq79jfKOkRH/wQRYwjAcuRZ/pn0aFrkNjiuLspe8x0s11B/CQP1RxUXXYFj
5GrljOLMEN9k5pgMEg58zEfiTvcqsGtrb0/v2GgXLgxrHMkvxlqtPZh0pmd3TsQk
0nZVrUhTvqhJCoWyollUQ02YVDdxVCw6rP0azA2S7GJCa9M+Ly2oI8MNWTVi6i6h
CWwjZzjVELN4h8EjGvTemFn8Q1qy7HpypluvgaAl6AypKdGjN1VgO0o3ZD8b2NBQ
GZb5ZWAh4busSoeghGDHj3Efw99jBZCSaL1U275+E3g4zOF7fx7cst8S0uMlTlNM
QXCwhEs1XXJT+8Bajz7YQnQ78FBKnbsTnX/KA1HtJslbnw8CXtGFre6Y8aswel6j
LeMrjORHzhVuQQ8PizRDcCrQ4VoqmzWsa/fr9Z7lxSuRrolGIm1TLwyD4uUViFEx
9ThKwvBw0o/DTzyECiNpDos+RN8xRuoCkkkOYpiu4ntXe85uENvcQ4MgCKwvkbVO
mERTbh6wiCUWpqL5vy+PzhIoVyyetswv5SwK5XdVK+tyMZzajrSGpgUz/MseDKEc
jXFlLVJVnpboQtvp7vK+gBLuytOyO6OB0Y20K1tdGtVGNVRKwoVDC92rJdgAe4Mp
JiN0flqkfEAb7Ldba3mBasKpqeVWxa5icbPeMlWAttlMexTHts8hCm19wfmQr4am
YUONvNVofZQoM1ujmOf4nSDkuDZrQ51UMY8+r76jFkgbQTKod0zrHqkb+4yG4rGj
JpcP1PskMQqjLxj1uCvQLxmyUd4qsuWXogQoijX33soNclmD/QVh6imu2zacatJ6
RnePP3/SnsR3erMfovLCb4pWdPQ1KZIb2Jqo5eSmnno7Dh+HKzhrklnewpu+bJHo
ej3OqXumSuPgd33WvFLH3/TZmfdIEDSTK6WOUzg70YjBpko7I9yECWnBcwxgGZn/
dpYcRx+eZoGwAIrSYVZsEQ685chQU44OTSs8iNt7FUyx3R8dr7luDDdALy4f9gsf
BQsMOfe1fOTbMfw6qISnQGaUAdbMU0Fw2WWXOmwkqmTedXcr2T1HANumO3Se9MKj
4JxyPrqlV8IwkhbLOMhBa1OAzeq3iW87Ex46YQpDzHcCJH0uUPMGiORbf6ksFjg5
PXNaAXVQIOxxtMRuGM1/UJ7bpDG+rNnoYV9hCYS5E1fOnhIV5ef1jGWX6JVpSFvG
NWIkXXUosoxSPbFUD4KlsSrxleLIjvSk8wXLtXjK3sILa28n0vcF81CZA3lUrpEy
BRs5ZGaGm6WKwrhhLc0cvlMNXuK/UsoTJmwmXH0D68SmeFpS+/TC6TJZklJWltY+
Ht5SIIMf2hNHdWqyhQlEfYqV0rW17TRhBCoOz1revdE=
`protect END_PROTECTED
