`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xCFzu3UUGkTLb63FygnTlAsfqg3cm0dNDRrmovVTHd70KhajoXQTYuKXPhXUA5oE
d86zx+yjNnoFRtlge2ixo8o6IhmCWc2Fbp1CgltsmOFzwgvpVHmh6jITbR5qRUDI
5jEy6OlprUhdxuZ4C3zBIDat/AdmWxquk/TBlXUvgGw2TC1k4HAXKXWCw3tYeH84
THsVTZC5ap3QZAIypAahKQRL/VcGZqVLKsTqBGNCEd94TgJjd7j9tfO2k5l+mvt0
dGG9eLhNWpCSeLxNEnhnRAif5aIG3oBpYLhgdfqFfUZ4iEyAu/pQLHhSh5VaNr74
v75Y229CeOQJuQp1Ty6eB5iw3+vB7iptAFXNSfKr/CzUbSqEFWMsy2XqHjA53qV5
WAHik+jTrNEw+h+vHFmla/TV1AHqFe7DnHCoRVHZUpyfpNNLfPYQA+AzhGf4jI2u
BPhy1tWbsXhr3nKmr7RfOHvZ7fE6NhquXw09QwDDALNvifz9IBWAPxQKTqUwF6eX
3q7a0sJB7fvCwTtLKF4UXKQYScNHVHZ0jpRSrPQ6srCfr+KhOJ6R0lnkt7M1FJxz
9HmicwuV/KeGljBuYnF21Cpgzoxza+X0imgNpPD9xKr9k1GRoEku7I5QaKq0osb1
s69dqHWzYUOpVSMjN5XtJTVr8ECZPBAni3PiValmFhniiJL2zsP+gVpr0FEBNK8j
macCtuKrMCeEBb6SkjcerqeHCLzLF2SxuvwLmnq99bx+5KxZY5j0nQPB5ZklQ+ov
Wjxr40EN/S2omtjxJ4QU/DBsl5FkLkPNKD+t3Phj5xrwjS0RhDwzZr5n+Wy4KhnA
oEjb4j7ezi6vvu9Dh9c/1Mu99XDxK9IDCupxtbjmuW3X2aEGRj/fx1MQB0twjomn
5hka8kTxNS1YcQ0+Riz7qrIgayOrUrtFbWvmfrBlDJBywKMsG8GgS/Byr89RJe35
Ea5ebbJUiP6BGmYKDr09leQqie6z1UQ0EvWk/Nt8dkKvxsI92zi/uWFDghfzeY9U
k0lcPOVS3Feay/5NYohbX2Ve5yv4/SjcLSttl2513fJDEd32gp3dT15H2cT3gTmg
wWVxZ7DZFORcqlPS0xu3JqVM8UFLUXqTShGaaQuNjE7inTkn7VdX1NYd45kPJ1QP
qR0VwbENVlLvNBQXB2AcuOGqLx2v2Owi4Ls2GWeHs8nF9tLeAJCJURUUBzzKw2ko
cToKkCaIzOFSMNDSsU4YHwso3ZvRXV2G+taHaXnIzcoMTZQvpDQTIjmrwecy1igv
I/3j2IPfGnp8FQm6QJqpmntoLKlC0U8B02T1xbuwUQU0r7T8yvziOQsyclwBSeZT
cNa8bkKzNO2zfb155o1XsBZBwueRzXZhtsJUNw9A4FpdkYgnwa/Yc6PD1nrBCsA+
VFWz2SrXMeUp8mLpRGYIq5kl0alFpVITLk0H7ZEo64G5CEsV/l/eDwxmQpawS9r5
VrTmnJm7dfq3qCEbS35SSUR8g8Pv7KfNlLV96FgKwCAe6q83UcLRbXWzzZh81Gqp
nJ3Owwhk2lMnGz9E/lnLJsYUIMmdfQdbjFDdh5+CHWfu5a1oGljxPm7dgiRG3nFZ
bYeN4BPccEkkqR7tGRkkK4MvcF/15Ca5qX1dcKQ7swPwvVQjhfK+Y5j63P8lpyVG
MTLh9myMclHLte52FCSet5DePFZ7+Cd62nze3QlWZGcWNxFUGDZ8lmVDQ2w9vPxo
u90PUkb/KLTXj6Et2tyL9Q3G49+qqQMeo+QquBgecoe8ND3/oxM8OhQwq1A34/kT
9itNBo5w8kxmGsF3T64h0XSyJMolkoFsG8j8wIm0KzBNjO3hKyqz1JpCBwKvi+tJ
1hdM8F0lIfsdxzKFXl1vsuAH2fqHOQTR08qR+Ae2AlRdzrnGDHFfNVRP2JSWzdTi
rGSvCv9eCENtBboeopUiJYJZe/Zet0kDbI9dYic/mvTTaZ0Ra5Q0dyg7gsDjGW35
4CHARnmpzGdPmB10GVJMOa68O01tp5HTTT5p40mrWpc9DBm4ITNYbuzbqNGW/3wE
4QHvLn5oT2WoUqhSOwD1iAC3NAmO+uuBKWD3/EnLImtV6sEwXurZJd23hK3HSGbJ
X7jjrqUHPHuASHKtqKFb7ULDzqPL7UoP896M2A7d6t37BazWNl7gIt3HiQGMSYuv
b7+iAe+bujI5+DcX4HUfxDIeFKNA8Ai7Q6eyHeIfcuQ=
`protect END_PROTECTED
