`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PQK6W9aqj1IRTrrCjv/rfmmWtrm1hQ9gTqFFvvvimSHksOU90z5AAjRKrOszZ/Jg
aMRPDsFZY/iXICmu9mH6O1rfuS5gRo6hwkUfBG/slyARIBnB23ezGIJZVx0fjC5g
Apu2yGxpVyld5YOEllWvggK84+ZuMQMNTTE/MXgszXVcwAXWMR5TF4Ffp3T8FYvT
MRU/cdpD8n2KKG1QlkXpA1T3Lj0blJExGcnEV6FT1XZiC0vFy8p0RPk3cyUpLmRw
t/dE/VesR4rrC6psz0nkafqDPuHBnA5rBC1L5faNW2qimGoGZBgAena2UCn6lOEm
f6M5GbKXLJp/qzIiameRo1F3TVNd/oKGiBgBnaG1lWgWR1+maKpho8YgD+Xbt54h
QFF9t4Oam7pDqYUo/9kbZFUlEEBFiwjggfT8RhmgzBWTkpgYXR68wi7cLVwhQ09n
gxagAp/r7BGdpworeXWndP6j7egklxKts0vLgtZRSnl1dsRUCfYVJW3eXXCPpiUX
QOdMCdj19KEQJliUbOLd9xYPz+3muFORU9ICK3wID2bo711DsFKBsQKUqLXkcl/5
26lFd0ftDSQj6KfTVxjudaHy9iuUNYPx3I0npTZOq45FwctOzN1Xie29riJ/lPVZ
Ti02ONnQmLJcQvlK88DkzqISOk7Agu9sA/maC86XGmg/JFd4T2Lgf93ecbNTPNXK
bjdp7vEpJTb4Ff6POYjRSXgjfjRQi2JEVQpfYQdiTSpkWquAdgZy2Ft9En7KpSm2
jAhhnMkqA/FZcCYegBuppvdH4czyJdCAjSHG1S6uXRbJJ/3yMrpdcKd/xiTCT7j4
qW6q1bd0+ymFScc8Q78XJi/LRtt9+fQN/9hAKWxQ3ZhJUK4VsKjNBnH6NmGZFrub
Ti+Ja5dPo/vTIBgfx0cJ9U2ihoVl0/DMHtDd5/Z9lBeoewWyVJrr++AYvXRmxhip
aiVHOovQWQ2K93YEp2Bo6ytXsSCTd8pXhqgPy3sSCqB0zIuhrxiUuRsUZdySErTM
EfLuCenZVHcFHM/HBOsWmhxmXEVF3f5ChJpbHvNITPagtxNQdqvIxCWHOderJPdo
haWIsu0Y8hWnAA4TFt3Phc7MBwbiLE2b5XS4XRVD6ffZN7kYfbBlhcltr9dNJnni
62fWGS2ICaG/xQOwsEvEQWSmG4+s8A9Cfczxu+93+Jv6G7GG65nxDX/t539r5qO1
Ks6zqzyj2HPUUWQQB3lwIoJ5RWhOQsWljWXGjn6E1vA2pvtMfbaFU0m56FqITSPg
SGHdZeo07keqAG4x7oSV8UaL7+BLPXbqRqlyTseoEDWuUP2HfL9hKBkZgnQesDe2
OGFL5K+h83DRiEClgT1Oo4A2BCgjzGKXPFe/dCp8XN2vDIpxMtN8EnFK5lOasxwB
1We0TNB+oJKbZzJcY0SYu/Z9YhQpXNA5LrzUocoAlVBKygrrSgs1uyE/PDFyb05+
sJypN9yv7H1HK38i4lTlauUeJPO0k0X0VP9VEiKg++xBkCXpb5lN97s04KP3ABgu
yLWn99Yd3Tq/rhb+P6TFaxbDaiMPavpsXXreHGkqoQcu6qIepLQKpdSLLLEnohAG
nhzUjThVV1mtYmT7eaq86W8Miv8yDh5V4KzkezXXTbVzvjN65PrqGKSnsG8dF6kF
I//B/vKxt9qzn/2StuUUAMWYz7L5CVY7sskI+opGYXW5snTFXbK9ZBZLiLisYDFp
bShuc5iYs5W8yNGSPrMHDa+5uAf1pxtqC2CrZVrN6QZjvAlVUWnIQl1HdN6FF3qG
P5TG0IT8LqQDNICjP0ZmDl755zaGlS7QuxekB2+hZs/1lLizMIsdTWXWVOYlolnY
RISXoiC+MZAWI4huyCHvd1g+ltdv0kIaZjXhxNUJQcuuyvADLnWtWU0iGVCgu3c/
2t4zpzOaEgbw7HxNtYPmpD6pN2Y8NeIv+84nwGjUDjiJh3D8AbV5vzuNxonU/lAq
X9kAP6CxzkK1bF0kqTKpJTwtqE/t1XbcAYrnJfQBAtExaQbSke8NaNQkUvUc21cV
5UFx2pApVoVfy/1TyTws35voT7cfF+zEtCgF3R+Mfwn9qLqwk6YkgQepQFdXZFUY
yJ9RkncZXIb4TKj3Afv/OCjDHkhB1gbHjO9ciTSxR5exkLVUTcAuBJBmc6TNCGoi
0/0fKWcO/y7nu78ROHBpbSbuK1cdEIAab0QYyPjoo5gpSj8WXPMLSW+7uVS2fwu+
MoVnUrBEugUUHoAxiqb87dO3sAF9OcWP3NgabfUhxWkbuKwsXSn/nAPolynXjC5R
hrgZdSmVQ7sAdpzz2D+Nu5IJFFlvGzhX0HdaerZKMSCIIf6tao2KaFFQLv68S9UP
/pyD0292ESJ/gp3WAN/BCK1EAbXf7eOqTizm+k7GVu/r2hIEii6LQmNzTrh2L1wH
bdVAzxpplOfRfQBsXSL7v0QT9Pa2IMnUrFemWAkQ4os18AuCcaHUKGAW5JU6VLLN
ye+3WO28sTOzIfyT/UArKLZIWemfnvW9ap8lNaDBa23+HAcRrl7rm559Snj9eiWO
8PYN5aHKauFSruP9Lh0ty1+x7QihD9TrcusbJ18aUOiKWemkj6CU1t8QMr8d1jUH
ntKhJ6kf7uYjBFR+kuYSlu1glLiPQPZL6mMTWD6JWmgx1KVIJpxtVLQlPt/MxIYD
efj1ANvifrcRIUyz4jaEs0YX6g/QtjtfnyjvfvbjqmxihHAPWlH14KPJaJtqWiYV
iRqvEBYv4okgK9C00KFU3hfmvK6HaG1Kj+1HQGEoeQQSHMtXDBl9wx57Fk4a6tFy
P+jNwmIkgWaeZsZHrREIjiYnWVXVxT2mu53vPWb6AkSRaYtcuSn8YNBjuZajBS1g
uyekI4QCivRaU9RoXGQePvo5xfvy9xb+AG/sz60VEL1k7BeoW15Hs/6kuW3ERqS+
e8355GMlAb9Ru7yEYhZKLxZzKD7bLD7bTQ6uyzLGy5XiXy4AIKcKCnh+vDbsqN5t
8otBb0YeN+IiCQxRWL/1QSME+MXdZCHBIm25C3Q+cxBpF9KrQSpxbHnw8OlDdTUh
OvXNInesTauj2lnmZnsZO44q3W5MtSDXrE9vax0sAsD8O1VP6PbXwHsGS9xXaYCd
WxzskdQvNe0tqfnERmZSTsv6VmE79Jtynuk9Ngwam73jlKHqNO8LX9OWLcwrB97C
99FGI1S4LJGvFkf9VPal5ELA8VD+wGVy/2rEGr/z2CwR6dLpR3JopDj6p4oycu0R
bQ8VLq0xm51EczKEnyeS5+IJOIdr0bsFexRJDVfmJaQdX/lTzRjDgjbcj3oJ8T9f
6MHd+0gYH0nCEpyGl+tXL9qnX9q7ZT3ANe7gm2He5H0TX1cch2zRBu84sLYI0YZK
SckEuacfAA7x4DQ7+gICsnQ63NM/v6pxMvrMxqsSs+8sWj5rY5MDgDH1TV3m7eBc
XZ0WrLv+XPR0+A+z2IzUpo1Do9HhE9McIqFZMMyEuUcYCavkOis8h7BDxlradVbX
VG8kchP8iUEGWuT9jOYMvuAr487gFfOIj+aaJhKmwXanqalWg7lAXvmIhKmfAFPw
QiGiSmCHl6SKssmZcW5hZz0LoqlVu9GyypfJhgK4r9N9l3Il89lKPd2G3HvEmz2r
Trmw3NA0Y+fWbetA+H8F/3NVEuZiusZiptQwZWCSeH9kBIwCzPQEPSwyJy/kZeLo
lyuCXrWEX3Cdl5vREDk93GDRo73d04RYPls6+1qekAXtR3HB1lL59mCATITIhx5C
berylnv5SfAIEuNScPNPNJniKnrqsVkR6i4sS1YIBIJDRLTHpeKqHe2I4dXBQ0i7
e6gYsb/19YiT5/gvAM//lKVfn5xeTIYR0L9efYoECTiB+pWawSGSqWLRNT7ADyOE
jgNuwMgwZBr1+CbNN7aHN0QmbTbZd524FDw8ysICggMrKVMtPwV3z3idlBt8HrSx
O3VftgHmpLYzE++NFy7UeNnaztQfkEMytsvKkkP9W/ILLB1sYw9OtUdhppoeFB9N
MeEFFjk0O+J6rAdctfu2J5GMjkxbbzFr9LMbn/ajnS2s9VYyvsFgcER+Sx4fJBMM
rIvfX8Kz0cwCsrB28gfBhXLLmIvRhfwudNkRNz13hNHKcKI3Xi5z7Dk7YLTtQvu3
4e7HRw2AlWfP/s6cm/H9KUmt3HAEUeaifDUBcDR6HsCXx8TptH902AVy02k6sU3s
lwAUZkJnlLCnxbJ7tPpXrJ1mZcGh2OURe1uw7qD7BwyYSmbZS/ZSG4hT2lc1scIA
0/RTNIByXwk32puJbGKqYiiDk/uemZX7Qg8k+bKFzBETmAHtCMCd/RyLdpEWzvDs
FwxgLPieGxqZ2CNtHIhIWsVcRFpqICaB4vOo4VpByA33DG1wh3u8TSuY6CZzHcks
KdoSC9trF+NgwiFRp7Tk07hWeeSFLe4ArUiJlpZ+euL3cIYI+fwDek31BbJke0fq
z5RrqmE0tRYUsZEn5oPBBsmDu3Qp49Z9/HPsxBPC/MRelSH4SJ81WKpVQdFi41BI
LUgu81zoz2/9oFPkqEQRiHriay3UhY9MEkqkNL2hfoyFlZufRKu3G05eQFjHkkW0
VUjoa5kHSNJtDsAhNG8Ts9ik/AMqY9EVFowQ72/R2SZApVQNx45znMksrzQb2MKM
J419aD8MjvrrltTfNBPWai/VLCnGAoyqgH85qqSyivRyBgxUiuR8PRDMlP3K8zTn
5TnDrLG2kBXXSKBoti231iOpjPw6YKkGDkVS2HSjIi3RxygKW4hEzGP0WbWhqpfZ
3KDyeCsEN7XmCkRMUZ4WnU6mTn51FekL57ZxzwHM/hofe9ADr52VVtMJQ0hcT1Z+
oq5muCV1AdIcM3RA//O7kI7vnhUEDeSummA/EyWcZtEQGuO5BnJnVWcHl2WGdeOw
QFmdizm/UW6iCkIZ/9bqQ/BuNlCeV0JzDSJbUeaP3qlliSOQljM9D/ETXVeRQkz9
fYdUPoD6ItAzC3NXk4g3IgIW47xXfLOii0yH7Mkq86f2+B1BBTN2yBp+4qYGqE7S
c1/CvccmQMqWmWhg3ZEbHsEnlfFIYETFX0ZGBQ2Z8aOA0HA0TPL5LcU4BJHWUQ9A
eHd3v5izJsZz2KhXAH3lDTrFoAfL1Cxi3OklxYUI03eZPLPVRdDRe0qwFOEhQcLe
HRx1PsH8UP5ww5+SvHx58DQ4pMieOiEPCHp0R6Bs1s2EW2LxWH03uFjvaJY5ev4f
HegWaS8fzLMYQ7SmjdgFy+L4QmP9zZOfLj/o+Hza62nwpZKCvgVMDQMfWloS2f99
NDQSukJZiPtUiCmt+6LpLtwQ12ss6PozMqAkSstJL5AAMW5J5FzaQJHHjDZypTtP
IG3j2kX8W5w082Vsvm6jATCzhYQfUJdkTRGBn2jiUSsM6HWjtmqTzHxAZ5KHMpYl
KDNM0vDOigf16QIpXYsJkGViOOCy1zoVOUIC5v7kNTFVa+buKfUXXOLyADcy2/Zl
mkaIUGS9Psu58g2Y/27QtFWl3ugLj0MZQb5ecYOpjQ0Ez5nMmsJ+9fNYBhvgjh+W
QxzStlpqY3eHDUuBVNDPihqZztEQ4crVNIYbmNqDVw13O+T8lb5gzo3l+Q3hzg3/
H+fjqUYZk1ocgC5fj66Z54HKLVYUCpTS2j/vvu8kHEV3lmekgSsnKVVz6vNCEi9t
g0zM6FO/8Cxgnwwi7cmZLAH9hVJldpX53bubDeUjxjTAY8e83NYxwuhVauU/wmtF
8wxamZwpiEAx0V1VvD6DS0H04gzQ+TmmuDKxb/+NTUgaAh+VZQ9XlgYTKSZRddf4
IklxMNw0V3WIFJlMzhzZ9nQANERAXtPvgKYC5Jj/4ZUvD4R1ksCz9INKkFq9dK/B
WPVOJ1zeZLQj71iZIRF1/kydPs3vsEitNOQ9gS4IdXZ3VTyjdQCCoqdxCuoqYl8z
J33xirwBhqq8/Cfyx9IKj8BKpEYRngkVRjqsehwK2b6LZ5F7hOFarPtTNRhBLlqz
+dRHtdi2nA7WMFbCH/JWyGKLD1KtP08pC9fKgLyIFRICP7OJ4DEiJLchxSO5fYpQ
VicvnbKRtAwV1Yt7JO4+EGNCFgT1XJh1r8f5ccIDuboUR6oqvS6/ZbMCGJYZLetm
WNqxspUIhXqUdzNI780kooXa+jt1sjyJnxtyW9xQ1LDsCSQfoq9/P/POcsSZJIwS
2qoWZuY3wGLdUsgvIAE4OeCPS655mHY0SWJ5yYmI8KxJNVC9iPuOV9cVGWck2a/N
CRjP5lkxCnZ/uhJcLty0t7Rm4uqeadpMYdsS0jKIf5QNT90dHSIPUolEoWqXQQRe
eV7/ix7/+ytmyzpvz+Vtv/5SHti1wATwXSwaRAbh8OxF0+7JHz9EPmkK2DCJa/Wj
nu7TthqkV7sxm9Ghi9lHiqKrLZTnhD2KuA1SWeLYC3C9u/kPhzVHKiM/5R+4GfJA
UPlWfQtK4N1OyamyDiPFCqaDU4PCfsuCZ/EiAK80fAJpvXFDd4SY4PGBwvhL1WqS
u69llZuSf+ntq7R4WrjjyRbtmsXowyy+QYdpghm3He7bqKMthxcKCRtiGCLCroOq
XUZAjvZz1o7XuClnbviBN/B+RU46lXJrOfclmv9DfKZtSbZS5XAftKvFZzFvbBKB
q8Cwxjgi57jOMitCtIac83Mh5O5UcEaSZx9J3FwD/S2UlPEjvqGOmWXslUNO4jjR
24TdGSZHYNGX22QVLM/BCdNZCg+LrXYCdxF6B7nXjzDERhX5DNNi1vU1FPThhYjN
f0WIqHYmWylqimzgY0AwYIEayvygq2J5p9qDb/jpzeHAtDVUkR2Kzm+D4SgFGjMX
`protect END_PROTECTED
