`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7Xi+mcP0OnFia02qRamPnkqJ+z2L9mzPGBnEFAXHDtQu+Nx1sxr+pQDEb18skQz
BsDNp0KCEx/BiPFjMKUotnGx0OjfbuIQ+ny4QlIpVp/CFE27oF+iIOXH8z68E6M3
ROHYa4MsQ9PnqcKYn8Z5xILqIdJx08PpftJJ97BJjV84hVf7D0sHH1wyGbXBCbFE
q8+6gpJoDP9EshGLoNkX9bWzB2duOjst4XORL4bTGbB1vbCRrISL0PkDC0MgxZJB
qImrGj92r0pPkBV0X542AgFDrFlHipLnp8ffa/WpjmqH8ITMVU2B0195T5iX/bqg
2Gp+gVE/qAH9thdT0AZMHbzZOFne2LlHNHFi3+vQF5huXoDVVO42/BkW/cNCYwDT
/hwcPGPk4nBlVm2He8VHKT7Zl677fAUnoxwq7EvZbwCANjjSCrv69tEaPOHvLHLb
DQiin5utZuCfxaFyqFiw0/fiXTFq43x+W+8HuCIs2klUM+zxTsyTLSJ+Fq+Ukw+f
GxhzMRIsTI4SwkTX+7RP15S52xEKBcBelugDJyh3q/Vf2xKzTzbarV81/fmg9qvM
UXLsQEUo4QdDHzmpzEQb5M5MDdL63f1999OXVhS8w0hQhnHik+9bUTWdF8YawZvd
8j6yVS4EBOd0/AJcuSFcusHYm9Hfb9Q01wsRI9yZfUU=
`protect END_PROTECTED
