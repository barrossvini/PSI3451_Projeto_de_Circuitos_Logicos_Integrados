`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8CyBpmrpZw/vSnCOCyK9L9oGxy0hnhAH5RNLQy2DhHhF27aXVJi+2t3QC0riCqHf
sPnNGJAYxLMGNfXQ80f0EmnOYCw/hHkKky470v/h1QMa0A79PC0f4U1WiE6EZ8EN
iW429RyZ9DE7DgYZoS9I1uJI564Tsopi1LVEBTwB+MVckqA+JtEIj+zMBc7cm7cH
DsuyQ3YWZMikGwBnvbM8oaPvkZ6BH7OQvqYnbM9efyLglnBc6BCIjhFRVsjgxQQG
Y4zNQ8xgTtN8IvtvKwsK6HpsdHk7ujgaDf0AF99oCmxu+n1wbMXaSwgM/ns9vzg+
jXG+Dttx+rNbD+iyCYjcY3WTvYInl2B8gAVD+Eiy8ZXZ2XLmc8dYua9dby3+I7yz
YnEdm6CY03HLfHwH4ln+Fj99yILAZtS20/7RkSrbW6w8ZGGAi+BtHkUAR0FCbIY8
z2GtS9U3UxIKOaISjh5VSnoIRhkL1/Rhv6y9NCmRO7HSXDOn/vlkFcw/ocFKI+/s
kd1o9huG8jP/CYq2/mX+PsBtCAr96AK+rZ9TdOYO9o8r7fpufMdnDWmLNKb1vsUZ
/GbgjXRuFGDh4G2n7CKPVE+JqCLAVJ6HVVTXutYMlTSb75BtgoE74o3NgVIIYAQ2
LExlAkQydA1RKKhmOh+lpWNz67IEdRcHH9lnC9F1+Q+KId1KeYugVld2t2DUuvho
oDWVp5ZcdMcX9b9WAtP7xWKy0u8L1JaeNY6yBuLA514yeOdCTLSFsSwEAjRzdw1u
8qH9YGsBSInfI0/qtbtAaGM+H9JtUGMQ58/hThwg/sOQx/a8zCSj6fRF+BMcK8cN
VR8irKG4v0pXNnwQQcNUMLHHFM1AuDAsQua8FkD9/i7/Paav8MNBi5dfBZdFn7ez
89j+treEOe/SDnsmM65Xn2nGUzGne8/MzEGqYAvVTT0VfucCfXa1D1knoHCvfM5i
5UFHBbA7eAvbiqIRBfyA0vqJ51R70mRcpqgy56NQyJTYsoZVWCE0mPbg2sza5jYw
NZaSYnqpYL+aWyoq2K8nYACzxuWt7Z5OlmKP1MNTuDXByD0ylFO3HOMCj4y4Uoqs
LSdKy7tLWqH9enNpMNrA9Cg67Ri86fF1Fa5Yt1rdrKs4CKX2peXbdZ4BIAILiQ4k
YF92pf4kF8DII1pVSTq4Ef5AgJrhIuWwz6/OiGfKSnvHdwEMSVh57IM3sMqDICAP
WCYFbB7Ja8zDELXkUk3dyQ4ntdn1A8WQjXpcfcucbVLGEiMUVJNoyNrDq3blfKzY
qKNayV+FkiI8fhrY58d4ab1389n7Dpn1LUb0RuQLEpofT18yGxIik1mLpJXI4y2S
bIon5k3zU1S2P9sZ2V+AcPmS3FWTxtKqba7ovI8pjSEevtBvQH6n18UnLN+i9mgM
vVstUVO/SOrZ63mCOKuvVuDTwrceNO8ag45tB2+/AnJXmKTEy+C88i5Le/AZxhuK
BFOmAvUyiqv1K1hsxTYHRArzVUcV2q4bIaiqrhaqlwcjxWoXqQRRJAG/122tTrrm
LVoAHLs3pA+maMI4cqLyOrvBgSAl0YTdI2FUvmHXUFT2J8KdCiguKevGj41q6/CY
UDc0HM8U5cpeOB13AlpNHJ41bzWTBlAFFos+bn/xwTD/plj8p1vVEuIWPU5eMfWE
GAWjrVXdonhH7DV+5bhZozzeFEHDAvKJAcu8rtKITOEwTPf1WPJek/NrwJ+ipDYC
oRh+e5XOMZPkXD2kABFJrZlw8cTUpQgs3ijCO9vqDxBhQJl6Mkho0dLov2iTlQO2
jIPj/LyawtNA2wdpZUUfDu1X6qozQhdylx/sOjfDinnucWKYB/UWVf811KI6XUsS
DFhkFFRZ9Me/bs+WA+8v4+/0+d2fC50uKgleyJX0q/0ZL0luttGpbm7URLWBcFMr
eHd1brrrJOOw6/QYz5C3jFej5fqOSw5itxoXuHjrNUKmK19Os6U+hV99CGSfSJEG
Ue+ZRsTDZKKVJJ9UOV3QrzwIps7iApgsxDaxJzYQ8iZVwOHdrGHs9q55+sW1KlaR
Zp2dhKpHPKw9a89qEEy90hFUciSWOu9sNpazrjKJeXxrQrDViahq4dqWl2caOy1r
+LSBnzTw9Gn5gIT78XLK9H4oabRnTCjRViP7cTf1Qj2h6W0ywFVBZAloYSfWc1SG
rKDjZG99cHYpZ8t4W5vSrmjmgAzlIMtA+Q1064cxj0UP94pVvaR7qSQQrvSbCWN1
eu2fYCCCjhr3Suz2VqKAD6YBdg6xUgAkujhnO7MrGokkpnh1U9XCL/Tc3BCci8XF
Q32NaOIMHShALykmSFRVNCTBQT+dVrdXAQ0/e7Oskq98VFLHHxY5NBtOLINf/3ru
UQUJ26tNDdfOKVzU2Z8bPAFN2x+vFPfry+HxYkayD7TcfOHv8gVPCE3ppsxDFjv8
sHFmwGcbLPIIR6Rbn5XuvKzik9YNvWsD+z1AAI+SCPvPC1bWAo8mRaF51zGykVOQ
ICV5Bef4y5Wx0+7BrItF3Q==
`protect END_PROTECTED
