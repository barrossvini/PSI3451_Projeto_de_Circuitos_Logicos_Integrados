`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8HX4c4V5U5Lt80wnGzSJqeygtrB76TKWeIWMuiCW15WqieECvHqQyeJyhnxslV4
i8QOWmOKV3vYvQ5g49yUWU9DJ6diNSzXwY3wXC0AbozsGG0MnWPoVW5lWmXr5Vvd
HXZxWmhpz5yjYfIWA1D67yy23WQ0UDyfGwWkO4m5wASCsMQEPB3qsOgXh5hc/KdN
`protect END_PROTECTED
