`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QPCmNUTKiq+5QTka3VYlR88Dr9ZImHo40m3x5Ps1ltD/mx0pNhIfzSudfc2Aa1AW
QvD/NkqwQvfudc/9SNV0YXdgeXgVZDIuyhSq6XfnakReFtBx4kNReT/b2b3AD0Nn
JeEcd4WT59dpdOwrOB6KISk+8IuO5Sf2xS38b5bDfznZNIT1MWnIjCsvM9bgHCz5
02HsqgK1syWiSk9aI5kqlTUvfsxPV3a2F4RKzGu8havkhmcQRJAjArokKIVCNLKY
5/04z+vzptq8k+NHIxRfi0x8/UEpQLQJNHkdjkwp+cekxd5QxvUDNdyrArVpTpvx
oitSocbZzRrUrVedzh9KJwd64Qul5eb1FuM9K6RCf38sDI35mzd9t55B3/IPDcBU
9cg7aKXOqAzVPGdwipNJ73YPoT0QhmLeVFD7qSfnRw/wJij5Os7b6vO+npQ7jXgD
sn9kSjYdbWCehn5A7KLgww==
`protect END_PROTECTED
