`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kMTuokYdg9/tWWvZzTF87Y78nNOlxnkhwFElz2MaXpfgtNU67So3QktWiXz2TEVD
p8aPmMXA8iRoz0e4aq82KWKwei0iD0zRbYQ+j6VfdWYkicSyapxsMDCFi1CGfn+s
LpCJw0tSfPtrEeOVfXzwE9dslyYJUNd74zhd7pvSEJ6jzpAcloGhK8bvTiI0qc6o
FnGDQcpBWpzta04K2gubGvlKfTfz3PbcnMjS6D9JyK6fPZmPlxaFKhIl7t/FWF0z
h2z4Qdl+xhjZMxN9D2aSnZQKvABV2iGKE+O/UGnNXHq5OaqTBNUcSuzRjZtqKFwh
FtKmK6HcDjO+QpR0w+eaWkoJsamjIOsJP4tTahwpkdzOdfbWHezArjbtk1ybFwvl
k1gn6ZdZISY2PjxH8SJHf/4FpkoXBWRxpRmt6m9g3GYhznJTjWjICBAIRxLk/vUI
fqPlHPVq71Y22zrP83dqYYCILdigiDmnjTtBmuNcupCzoo5flgmS20A0SELY7uPB
UOeKNdEUjiYp4DUuY6ZvqGspnaSmUYdx02zJgDzSLD4mTXvvFOnLKCGcMblSsHGI
OUdRQWz9vxffDCULESeY/8c99NVM+UFEgLsF7oaV0mV5yZwfspBC1qEqT7aXiqEL
8h2Jpc8AfnOMnpjqOw8A2KHFhIcYpU5ZmCJoyDYTk0mk4dja7d6GDjxd9TgtqCrt
o7uoIqZoH9eSaXT2H8/Q30x2De+B4o/9XpDlvTC8C1vfRintjbNlFIFEvG/ITVf6
sdV2qFdHOa929ALrbvDdwtPR8cRzCnkLAlf3muLCSovG6hqm8MMKkUohODGB8xBv
zuKyGqt+D/dekfZAfSAZN294e3sPGB2UGOVGNPZKI4O5y9B24hAGYFV2OKVTgs1v
qy29ds+JvnT89mkqRXd4XOEA/j6zZ4qVlPG+k+Je9DBUycCFB2S1sSteW/HQTvPP
XXUERoyqm3M0u2kNjGjo5fyFxJyzFnFVV7EueBkbQjXbWwp5PSohirWdKzoUaR7p
qimxrZD4zciXJnLLNkmVoHVNxw8+4UWGE2V3n6gIaVALFdKsWFwtHQshsNShp4En
crVYk0TbtIiYUrRhe2ZYVQZKL8MjiZBp8YJ+JbMS4O0fh1wCo8OVxMM9fCyEydMM
ZQkP1BbIUoUEMfQRxStYck/vq9RB6ac3yR8NLH6wT1oeRZ0PPTvugA+uauN6EXcd
x0dSKhpy+JyML2szve2ud76cYJ2Ujwb4AHswtfQID0ay5bL5StrntHs6f1QChXxP
nFCsVS2aZC4t7rw3aT9CTVmbRBFoqgj2VLE8LvTppOUPA3sGeSVvHN372k8DhuCw
uOUlmugJtsnCqsUwJ/ED+nshszJduqNn5MXUzHDTsdLi3Lf61CJM4UeV6egaKeC+
6+ij/TGUfZx9DxTuJ1vRk3dkMphoywMzb7N/zHc3qHE5p2VCN8299ohN1ggqJrPF
SDZUeVLTOwdn9ss+0t0Zfij4zunskVPrJ5TF11E7fVuNNcF3LwXunb47E7bxR7Tr
wxVopG3QxpS5pS/8ecA2e+AyB/7YX9Im5mWeStc6bGvEmd9VBy5P7F0aXYXSzS3t
UR0/SRjWCsv0M6pw9TESgqAy6lUN+jckX7n3WDHc6ZaEM9HRrBXR1fssF31xlqFg
BVL4CUMh1CwSDF5xigeh60ONRNPTyLNQ7TMzJIPXbeMjTX23MyFQrb1gX6UJEtL1
mNZ5TbxxVXQR6D5Ot9yz6CWp0yxfYwd+glESDY5spzqHGMS+5pFqvKByAqi9PQeo
aoSPEBJa+fMcUgE6LxTTCIc12U/8J9nN8m2pYXFwg62JE7nYZDBTZ/hrxyxzs7a+
C7UUwFdU48ZgWwXzPe2VKoAF2EGBz0zhxSIIaLDLKzrzZWATwti1dbVx9wwMhBgV
Sco2I1ferlImXrayrXwK6NHwC7Wc5wEumPsLK26Qf6fq+f3mEMHIYEWuMi/HP1XS
1irnwar1b/QUR5AEZG0E1uJF50sMd2TZ10cCx9i83bcPUhHT5PiyfX8FmIzUvQ8e
3jwJsQnwv6jOezhsGZK3z4QOQeBEQITu299To9cj04Xmb+1CvXEy+jrEngPwO71U
zdPvDhkBRh5iWuZQyXLMn3uptldjmSbdxgELf3QscpL5JGfIOHPIABijfobDlkOB
GXBCCbVCoUYqYfYZr8uzJ751gGONKZezQni5yzmTHWPNTjh0FZAqAhEoss2xpDY7
vmo40zu7aOrEt1evTsy4AJSv94JFMbvnTundvRtXiYiNZD0ju3vn8XBC+sIgxskd
IqLFA4qeiElRQjTL2tzH1zHD9MIpeP6ZfaUSpYVMUADxIpqdlTE8mN0RqNEvvDqO
tg/xA7IVcuY9L9nw1/NewMzjKgkhk27wODJpRQpQDhhXtOD1HxzK1x5mXSyA3Et8
XwqWuiSODjwYSa+CBFyarg7WY3GTZlNjwUePYv6cng172azxPmOI+ryR2kowrxwP
MExv0QHuBRazYaxfg363QguEZASwU/tYY6xE1xdUM2K3AafvMztyWy9hjolnt6cX
wLh16gEIfx071l87Otv0IRt58KG+gfnQkb85n0D2DfMU8OnTuORJwQIcBXHuYG8W
6MBzdmnq3pR6vcm8qrTBrYHptHqPzZlyo3UtDqd8l9SRxy8j4VcVWH6uaFEfx68j
c/41g5O8Dse62RnOlJZMnYzrJm9TdZrOfa0e/aD+AXX6uDP5M3CRhRA9LV1yk7FF
djRfAdIlkuAUVEGhgjUUancGUBmMBEIKmejYmnHfLd3+lVbQt0huwOcuFxZSwczi
HYDdpCaR9/mZkmd9thLQpPwuYgsynB+K6joG2Q1szg9KTTL/JipVh8I+QUPVwWDm
TYHIqrehCxMsgjUmF0lVZrNQiwm2ieIcoluqft/EIivsG4jhepGSB1qw3K/WIptg
QqPiKDatkCOwAtd0+XisJcp54kECgtFh5mhN4XLy+06HMyhADHjLqCCpSnY+IRm4
so1b0J0SGotR2ywQuW8gYcGru3n5yTaV9dZ08AK6pM63FHXbwhPljuYuTx5tNv7n
OiO8qDyPJYJ7HeghyrKu5OqlN1xm7O2Gp1jPdkoWv/DrDEkxoZVuOAQIuoJWkw77
ZaXtFjT5wACaTtru0uNDGyYM6C7S3XjM9k6PJRnjFpJGkQ5MewvrKed96yEyhFXG
fvx+SsiLjFsP8rPqu7Ev+7MEMsuWmH2LluKOq2jh7mQkwa45qdz8k+nYdAOH98kU
7GsDi20F7Y9JWOEZ9stwt2sdImPMPTgKxZ0TdFUz4AXSc8eUyABHhrS5X+HFlnik
KRNNzz32E2H4LmO5kfK55ao1z6IiVBIc6F/3g2xba2qOq/xGo5l4S4NfWcNH1kxl
JH8Ah9qZlfN+rSUEgUX7GEsW2tDUFyTgRt4Y5wJzbvL5BJjghdWDdl4BC3NRKD/P
h/meElzisSkDHHmBFWKOdFrq1YbD7vSexzZEWiDGWH4vT/PJ2U3QgUEVArDBIFWr
kCSjESKNCE7JVEt8enWJS6SZxTld8HPIJhhv3sP3luVstDOvym2d2GGsJqtO7uYs
JvFnN2XdoY/6pIFwVdwAbwE+obvq/+FzUGw4LYrL5R3oA5mXAaPols/eMwg5IZ9E
ECTTk0zl5fzlk1dOz1Ug7b4ggPph1YEGY57iZ6hjNuG2at6Sf59QDyZ0g9L0mcnC
0Ctvjo3V3uDhbazSLQJ4K/5ZBq9ks1N68Wgvbwghl1jReI0PIQc6pI2GEIH2lGUD
Dkdf5+nqy5GfXoPtCM8Qv3x8AulhiF6bRPQ2SxQlhGHz5K03hpy1lluhKwcn1+ry
IBwiB+F8UtlNtObIHrJ7qHnQpAg/DSbpkMG/ETSwjo4TIwiEJi5Msj903YyEfj5p
89KChOysE1ZmoktUonpYHEEUKtttjB9tB9PGE7/CASXzmCcZM6PROJ9DtdajYqfY
p8OAjcIVrSNUTPnVHk/g1hNM+XD30YxDTWYC3UnNuoll8v/S1HpAO1QEnJXcRQlo
vE0tZqhOkyIoAWGXxSuqkl4KvVZbxAto3lMhF+nv37pcnlMgvF/ievNFUmKh+6v4
L0zPwd7plggzrMVnA8bCzUxiJfOc9oyk6VnAt+lKne/gmvvO227T0p5mU9CGbhUm
Cjp768GtWQieQ5ZXab8JxG877HIl5vsfwOfr6GFAtdGffoep/PF8JA/h9pd6k6mo
fFCLf8fRJwpFGNhaLMFe0vF/7FIydz2+Kkijn+mkPbzwDlj5tLp7f9ADHr6d56gs
kyXg+VoeT+gS6nmpr1tHVocDq+QePG0efMZVmn/ueFzpBmZbFcpXfsSSragZAq0S
zQeFGBkXbJgtgUV19AubV0/OC+jYGUNDKpdaJdzwp8nGp3ScYIHOw+LEnzmalAmj
aJxCWJApJFNxFlV91arU6GbXJK18yxal1w6s4D5xl6ngC8ZnfMuu62vi+foK6ecV
BFQG7wyMMq7Tg9Cg1PcXEspmJ5Cjz6opHIG0qkH5pyiOY3xoFhVLoi3pam7LQ+94
TE2mhuETm7/kXKbBBeVu7W3jNP8ruZNltoLFJTuERGWbs11G5wIsEyk+8ZO12zEk
XF4B1rIDz44Z3g/C5GegQ8pm/ZhWWo7FrOfpL0SfEg4k1WoEZyqASjfxNH/NOrnS
x4Vr/4cCIcxRrmJ4rlQUJZQ9efYHXFBxGY4xe908hVanUuUXSvFMR/v5dGkDzWYm
CHDQlnAvj+XGKMdg4W+JJDTRm/VGpDDkcZVLzCicvt25niNgYjNvdFVpySa5reeT
dzLLKWtSK89mxBSWrfqTLks6posmxc1rITnU6E+RKlLwFKFbV3hQMAplXFBMuac3
ODajNWqU6+Tbmve3X+ol0C5mFuD5cMj5kUcFxi/MGqk3jnoi68NjBb4Qe12E7Zoi
DSGpjScSn+Wj0atMONwzSWcZMHcxSwA/Y/x+LuXBui8zYekvhNGdMurNBiQD7qmF
VwLPXKIT5cz0d12WVtrU2hAKH2UX3N/rOFbMlcbQJq785Iqvq7eqigRbK/mI1ZXe
61qfEj9ZE+pqyjo1feHp/fllNgvY8d6ZaPt2nkJxBmJiz30d+/KG27sw0WpFQMIX
Ru9TQDCLlJ83rpjrLASRdDjgIAbu8pFzHC13dFYBeGueUx2cxkQ53aqBNVxFnDsX
cTgX2p54VWYyKeHkKC9m6DN94lyfCA2wh12whUZ4HgTH6cjYLxsuNsOEGG4LttJ0
PMIvoyml888D6VNEboVFOfgYyWrZcqdvjK5uH11jDWhbqvPhoMNL4YqxirUzgSzm
W2igShWgb86PoXzeVc0x5ylkTbloawEakiYguMJBFvZmPMXEhtNhA7tpmZ91Lyz2
CuOwAjmTvyF5iNI7CYC/69EmfdJfymbxIGQBrZy4HRwTP/TJc8SBWSmH6Z1pU26o
5tQno03iz5G/bp+D2b+prDG2iQCFYrKNk5f8pkRhrm/xRdRM4tfhm0C6lavLqsF8
fcuVz/AcT3q6QwTSp4EqOTDAWyyQ5VCXSOzeLBrsCsXsWXkvDaqo7ykV8LLadV7E
VPldsB5LwzdeokCVN13zoEuPX9M4HgDkO66vvV4Sn29HyLgVRbaSamGee3pk8VT8
E56tA8CFdCZ1u3qsYwwAdPdBh5f17anxCMJWkHE3cs0+pf2I7DwZjH3POl5c46je
svrPrpseYPHu1YswZydlTas4qj3GfUWnOjNCfmprXpkXnYITJVUzl2Aj1Mby0Kb4
DoFL/TIczk+gXvQaZx2SoNXHHEi66Y9y1dKoVjxd0SbN6sjbS8GCQKXOiL39pDMF
+RYDYPm7SAoY2+6xsGrEqvEKkrcKHQ2yLGa/kxzVYBqp5H6ni0T7dF0XSX3bdhyh
njd4/+qoln2PVZIXTUjcewrFUjLru5qM3A20DuZaXI9pJKxkYtZKRfB6ZyIUTnrv
DQmn3nJkTApFGbOP3H67pCD901AKLGrUOec/2Tlus0+pW8IiiV1Qv1LB8/S583g/
WTND8hxj8tRe3uMMxZTPWHlFZ2fLocOVd20CXT/IILgb9HOxMl658EPl4hbJ+/4w
HJ5GOiaF5DXhOQK8rJNadiO/1cyVDxKlpBED6sTUfDDwBdhj0TckJLYHY6AcnBhc
IyaDRICuWbnbnNP+4XvHKm3apaUcYBwHdd71iN0O2Jjta0ywKvEk/523FKVWVO+A
YZEZLC2wFqISW6vIPuQHl8q1jXRBqfnBs4vrtnQN5rJ+Q5bjWcwCcEZEJKa4SQkY
aLXg8o4SoalPSG9dJ4HGb6Wj1GotPqnFaH6TNyIOKhaxXGx2PIFPsdFHA1dkp4Zd
kX02gugItXmyiaoLS6wWqiM6U+5+hlg2Cm7heJE70VA1+MUoQZtf0a/rDa0hWHZ8
dqgf4crTvCVViMggm4mYlc1y/zxIaNAswLc+WJLqTbtr3xrxQataHTiCvsg81RvM
Lp2vwjN45cgrIfx7HadjFfkv74J/1gdd7S2B+CxJpjwnhIlBHZjl/sLen5IX8NCl
gmMhCj7Vx5ElTrGAGRnRp6gFBmhCv350eO2dxPrFOg7XS1Z7itYXGOcYBmlg3SBs
P7y7jZLlvEY0OcNcEpMwRNa4Uk4K+I2QWPG0hQKSW64g6eko/rDD3mvpGzk91WAW
OSECxZnUACJVh/NlpNsjTCm+Qp+V615ym40gqHnrQ2atrbX2dDsn8ErWB0I0osKA
d2EOUryUf3FAkM499ulpgHmj9FayN74c7GUhq5cBdVbHa4KvNnVD3JwmCb1hQPel
eD9IDa6ck1OApnlTGYPHnMxclKFuHgZNTA5+Gn7X/TqxqpRlq/BJHzqr6VJKInWm
AsjvwXcS4s93JSTss8mh6UlLLr3pVRG5b+unZsPZe6Vs39wEuuf2SVzKJ3QqKISh
tqmXQg39Lbj9TlcOjnBKIIkfY9vYUpQKpKLC23deIvmZNtt+tmUHSNT2jNkhIrN2
AXpGOkGAcvcgQLTD2GVnpSf+NQXtaqrlTOaTjM02j6UmEATWa4Rpohqi7sfj4F8F
Rx979x5NRLKQUod/oWhRNBrqWCP60/rxAsAQwpLE1zCllE6j9nlJLNk90xU4r0Qz
ucgpNAoInNEpzHYGzulJoOi5ou1a0XWt3T+G0cvKXDmlP2Ci+CFBSC08/tiaS1Dn
K4DtuzXoOJ1a5unaDst7vU6Ig+sK1NSErz8TOBtuyKAgTv3Pr9UAP39QNOLJ4xKa
awA168+IHfFL2/fuIq3cfK1Pysj1QTpEEpd7QmHaJhE=
`protect END_PROTECTED
