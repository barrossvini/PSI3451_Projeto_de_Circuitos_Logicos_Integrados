`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eNkbarWwrTrAnIWMvgPpKBkEwELqeYewYA0HXwtSj7rDpVq0AJLdiPiXm752EH8R
hDF+iA33ozG68pZqcZbWUqFgr+MPXOOv+ePtFEhGx9grqyo96nwpoEChYZSgWB5w
qL4we7VOAZvsJuXMrtEMis9z6wrVhPrjOWO3Ed02sf3XqItJRA2NTG4EFEefiYE4
1LShJa9ilHSXL7N0ZB7fTgLNkOm8hCG1rQb6bL5AymBDB4xGfCcd/oDP6OgCENoi
mfCbODF49JO9VDLGrhgHdKdANRzJ3SbNou9lwxOLBMUTMXPGA6uPT+qlOT5Gjwkg
c3cP+MuRNlOWp1jpnFg8p6FSEiK42huJJzjrsgoJ0i7rxEcIVyVUnnxNxxsKBmEJ
WiAy/xspopOZWRGZo6eWevgjXqwtrOFQqS03lnmiKPYYBRaOIvKmoaRUFrDuVrWc
iUBp5FJOwdpvu9RZMtZlfwPIl49ggOqL2Rs9b697/d6mWZMR5FiszCDBP9ExPHxq
g+GKP/x5iYN6Hnsna3/3qCkEW/ZzKvqy9FErwzgosiXxEAYLektOZl7wUQM4dP0C
694EhR9b7YhZTFKx3ojXQpJuAmY9JTd0jVTGjMMqhfSHmhTE33/D8IwcMDggnv8T
kOtGZhZQD06tp/ZnRtiqIh1O7wPGhlA1GNHm/d//2B6xh1P/g0Uk5Axkp/70q7o1
4cD+cyezSyWkCwOPPXgOFNZCw1fH/sGckYQyNTi15wefRIIg7uX92YgkWM+Djifb
f0Eab6bdA4lX8rHJXKYsQ2YVO0xPfphgskAQybgq3fsjwhVv+4CNpFHoQW2n7lGP
9iTJxjZihYfCGo6MuahsVZFOevl/h8FoCehoj3qO4yZgAOeCcGvwPeyRlWizSCbi
/jkDawjr9u3fBGPWg8Nb+PexCM1a0ePZ257Xbjj1sBJjNsBjeKjdQ849MND5seca
7i3mvzTOsm/9BvUGQGx7ysPDZeRkPoRiI+2HPA4WuRtw3VwYG7+XFAkI3ha8sNqO
87bq49iDXQImk8J663wNeN2wZ4bNyqQtIpXMrQeIyTU5mqWAipLKiPgdSQUDACVO
M+x6VbfCZUCv6ojfRMqh54+fS9bsGPGq1qS9q0Bn8oWwixioYJMrC8USbp2q/LZ5
2CnUSe5nc7ku/sp83AyTaLcAeGUWbHBuOzuL+wHPpJWHbPQ6oIj3P1fbNfD6swFn
JBM1tR6Xc8JN1KoTl+6+YjNhqg1IpA6a8lx6k2xSrFhNUoUBJ+VnbaHXQHRlKx9o
QX2hyuS//pf2PCQpCA83lQlM0jO7paAUp8NJhzqys2pNJoBSX5t9Sr0EnW/NuH/m
1OOmEqGS1SkC0xfYTA7MNZOnMScHJ+zdiSk9ZMJ1J6FOgkyd9tq/8GroXp2daYJ6
ogJTBgwdstuNYsLnWep2NNt1b+4T1OQTaXCv5Lq5VCnVFAie61VGB5AaEJvuanSd
NkfC9hJ5TmVh/KjhM3kJ/rKvH9qrRFeChbUM8wL6zM9kYSGrFJzOCFDhTW/RVzql
WKZ8+YqRk9WgUZ81Ew7ctPHaEYUH9TSsQpGUJ2zbjHvYydXE5BWicc0yppwoAwPU
n06a9cwpx4EvZALlLmfbWI55rDey00iUD0DaSf51Fm+zpuZoUqjnKqFdWvvzC7XV
rqH+OXI36UFKh8dxtu/8etRUciUwUFa8yTpKt12ssmuOyz2wmBJqezY35eH6nJ6m
jDmmsKLqA/apIiLDjwWs04/o5A/8hrXSR4aUJy+L3RvaVfZFMtt77fh+KZYaeqI6
qFfKaAhaRN+3ST4LRxvZltTITO0enk6QZRfzQes9Z6WRA+TEO/RZH9zir7/SCS0P
vBg0FTRpSb0LgTgL/InQFsuC0vUXA0x+j/ssTJtNNO19/Bda73zbRKo4YXnCCbZA
xOFIUEvn8vtONbh+uKqw1yakHVIdY+jOrDFDrou9Qoc4hm+QaVn2z995lKzmfF82
5o7FwHJSoKlwPUSnpWptm81EvhDbanljmqTm1bLQyF3GaHgcsYn3WZVZATBPmTJZ
oFt+VQlV3vGRfniPkEuPgXVazLkPUOlHu4K1avmAjDV3j2IcWyPaNV83C/kDDWfD
xQvwlNcca+2euoHjHDkDnmizhOEBdt4vY8OvkvKMVMC3Ujx5mRNtP9Ju+iBJBe71
RUpD09tBXuOd0nal+ApyFF7OEN+LYu1mehq9d9I9gPzBODotNfQFwoUNT3Nx/dJ7
9VeJthJj9vZ7ekJ24ilodPEQGyc8ETYd36kdsfW/RfCSkaXwjPsLtVdzDBz34pku
Er6GcHq+W4pSTyiK7Dquzel6ny3qGAu19z04tJiyCZqR1F837uHRZEb3380QXGHn
cw5Bxi+maNA6043yYz/bx+rML/oE0OyQr1Y7Ay4T4CQ5J+YfeBDzFTdTcNTmTgnr
PfKQ5TgUXXfu5yxZetZU2HNrI7pyIGLCA4O1pN7ZGWISWOD6emay08VfD8BmvVIn
B7cahqveOC/rg8DcSy7W2J6iNQ3uTotUsxMfB5S9eKrWSn+0lJmzf58PG4guIARV
+OOlIczdSkNUh3WlzD+4yJ2N/2Jee5KhusG4WyqsiCSmcyIe4kTNO8tqPAVHkHLp
UfsSrNB2DddBRKZYTqdejJVA4PKxnwrn4Fuvc4Hcx9qyviELiEvYscQ08Ep/kaNF
2uAY5ERjWhBQQRsg8BvLlrOPV/oxgcwX/nI3/d+mVCFIsUqU4gMeDPTe5GVsR1DV
+NRTkzdph9V2awaJ+p67u5neXsiHQiIA+lODPiPKIhNoNpqzlGvpg2vf7dewTOsM
o9vWO07NndKLOrBcCECk53oLa6v0+WUaqiSavlIJsdmreaTOGw0XupEL2ItzNIBC
qoAa7Dgls5vc88TYETSYaIizC3vGo5QSYkVWWJ4JNyIOWtBlv3kxH3muUA88XVIA
EszEQzBfS8KFjfNQ4hDtCpfPCrT1ybU+IMhs7gGZl+8lJEHWsoEh4pJp1BmmshBX
0UvtIaPVvwf10/6gNbjG++5R9LzFDgDTfXoubts2S0oYpY4h9MrHs66Kbkv9Uc8/
vzVZwHxsKgZXzMoysp4TwDN5pb0oDrFQEPh/kAjjrUowxVAfMDgvpGWCRJoxLux6
Q/UpWKgmAEkJTKBEKRNnwnKpoi/zZkXGm6SMRGF7m1VQFemPVhOR6SYHERnqooF8
eHSliN+cnXxRdB5rTLvc+tCu/ZKcIxqY4L4XxGXa+0NF0WcfVVYULP2Oqs+CjDWv
0nzC04J1sqcNfw7banOJ/L6X5mozgLgnz5bdf2EGw3JZ/eyD9A/QOFVmxlrcgEDw
2yDY4XHlHUWsLTikEhPh8R7biROTC/iJVvjl76s6cd+b5l0R3dJuzQXK0Ez1YZMD
0luZr/a4Vw/lu+sk+rRnCJc6RwSuM3MEjabdhzo2dYMzP0lHjUhxWMBbb/PwYLo8
9ZvC30jW5s8u628M58EAzp1J4ZlIAxyRpsV0VBGUccY=
`protect END_PROTECTED
