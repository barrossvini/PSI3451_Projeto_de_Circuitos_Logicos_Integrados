`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3zh1I3PPtCrXJxjdTewlZsu0mlnXIAfEb95w7pzak3gZ2XChQMv9JKIJpZJvpgEB
h1wj7cgo6g0/OZTNps0HM7vWOdCiwV0P4OREN8aR7wsNfuqVR5hfGRrYbSvvWi/H
QsKwxO1Jgdc2/LNgf/tNiGHILculULphxtot1G5v+WPQPi1ZTYPUUzD19JQH+HsQ
ejgIOcJ0tOdrfFj7bdqZ9twvxd+O1505A+RYnovbGFeo/roTZ2x8qblr6WnKLczb
RDL5CBtzlHTVRz17bwGF60yHym297pDp0KcHBlt0uDaELq/5bQGmq0n8+RA6b+Y6
OrldiB27Axd4M5thiglAQlOUdGG3a2DpLKjt1oq+TkM0sBR1ob+6oAXcD+mzRqg0
6JU0CvWlXPrhM9xKAUrXbuW5xexx7PNweGXxFACVK6T1TM4a3kWMmBOn9VuyDWzi
wUqS2wgFFrey0tRfRk18nZ+LUjwTBqSkezxGAXuM5NWNnr3JrSs+bTiREu4DiF+6
a9ExczF6mGmqCkPRVHKr3z8h21ZQ+/WTu8SAnMbUs9K/PoGswjDYZkrrqn3s4jeW
VHeJdycUxe3sRDKe8xkPnyiGXS8ubaTMNty8rFv10vZzHE3XaGcRSJoRmQLRWC83
ILGOuFLpkl48bBv5pVkG6Usxp1fpzqRZljc5F6uUf9zuVorUl+/kfg5dlC0nOBe7
XPQBTHOVgTuQfWQ+AYn95U/1Gmg0Z1Hm3JBTM0h8Vc/uL9pVYi/yB+sWZLmpnUoJ
mg/Hbq1Fobg8icI7D1qeFNa5qlKTexqI8SdfR0ajdhkjDwlRTpQk2OciPdi1JnZm
5Pavfywm0nL+rk/MdBrxgOVsjI0WDcKW5EY1WjADNvu4Efv90rUX7hgPdXb/olDo
pR8PtVsn9iBpgqYHMfM9Gm/cvPv+n68XUxwgMpXgLdt6EpXuLfAXdOSVdTlWyAm5
P3NRtUadaBcXOXSzdyT6ECpHqnla+qdrcl4DrDrgxAxR8uvXzYOnCjENxblelMx1
Tk0tMp/cuMSza+ag3r2sIWdl6bo9nhCqrGq5l+QkF5Js2FDo5qLMXoZL1fA34RtS
ljiTdP96CGW20sS5V7GsfVOIfRWXgk4WW+YrzDYFVwSPJYqTYVM1mNEH2ClspJq1
i42Kj2aV55n6RVJxGcaNHAou+gjeJm/n2arLgVl9rvVtDmYKuQsO1UA4FCct2H9c
1Qb3yDV9ULiWMJijGuj88Ef7SBHTgTjb4bhYzqVn5Rb8Qc8Om2iJgz+irn+bMUlB
BCEaldtvUBlXtvFya3dDeKf76rT6kZ7NBKXtfJdhVPWvO2P4r1TtlAUgjfYG+5L1
FTrpBarvq08f3t/2wbezY6HIfWdRswBI1YO+8avZOuKq9TVQofubK+LiidXCQraJ
c8sldjxX/VvwTPtDaU0baBk4mvD8DoOq8K6sSAG+ew01A9jD+Iw2Sgw+g8iZbQbQ
lLd/KfsDCjSHl3e4nmZpDX78KiAnM9qH2epeaQ9pUzLIAPQs9NrPnxkDut+h+Kb5
K8W5E0kT4BYvA8gwVkp0CA4/BHId7tKBAcYxDk1+hogz2dBK9yQWGNCIUZhTrCdy
kV5+duvet2yFWCzYQ/mDa6P/Ic4lkXQEKzzE140Ar9VOBPZmwNFaGpt4VLUwG8oK
GS+yAmyFijwfKUf8WCY7GjHrBDtUShtmnSNl7m37RSPqqjGLKozlNapiJQGXAUHZ
7KqXQPA6YvH0zbu9oIluSFJN1Aznj/TxsTU+j8JJA2yr+nBjR/Bp6gl8uY7UwkCb
J+MXMdUzNXx4AMFgWQJCxXHPHXUR9mnSO4DO6BbJzzorQd38Evq34EZtxFaIi7+C
nVi5zRdDBH0lJzHvw/hw6qzuJrMYPnblIZe+dXKyGwu7Vs4jE+giz71F2hE3DE9u
DtM4rIyP0pl4+eSQYbk+UMpjtgDGOgdfWOC31LW+5clgH1s2uiwkfWwcAjQNJClZ
aM8GDtZfW8r8T1fHATfc6ZP2IainLKjQs6tBpHmoFQRbHIHBZ+evPQg9r3MDJ5Hk
cHv7IQcSOr+Cd5FYGTCDRbwb4pHlPY9JuWY8CllQ7h8/4NI3LmXQLgFHbAfUYTwo
vlXZwkJIO8I/TGTlRI/hBl4BDZ9PdsZ89IvUaUKiBQxW4es30lwjAPJzKDDEUAtc
eFAC+6uApcNosRWuLY2oLe8UlBMnamZ6wfzIjXPmYBq2HghbyenkDpU5+JMzgS63
guBkJbNWL6tdN2fCxzEvtYwuGDxlUymSvwvbV+InTzj6BO9RhZOsEMfBMhOUzxQP
tWV/6NUyUMrxz4NE5QD2dw==
`protect END_PROTECTED
