`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TIUxIldYRnuMX711+8wIZl0ukazwwstXHI/l2riUhukEbf35r3QK97QKONUWKAkB
8wSVBcdDshuWS3wHoo9GeF22RvjCjoi8NnaDJMeQ9L9+fjefVqspxKh2UejaATly
K66fHIwOuLT2sRg0D/D8KMh6JaT188ZluekUAsAtEF5kR9MChfuDKiLTMg4dZK2u
mCRQxfdi6Q/EOIFG6xOWrO/JTZJexwW3Nz8RYIQGk1srj1oP6y0QbosS73V8ib5p
C06SJI3J9BYyqpm9xk8OTfnVj1hhRQt/SQXtVtwnJHsJqgW7k3wIwE9zK279T8p6
JL75Uvi9enQARzYSExmhIIdwm6FUpznHC8SzzTvjQX1GEvmNgRIwSztWZrx3XhZX
GYzyUxOiAyySmwWyM4BPtFNdOTTnMhcG+4a3ewj062219XxeFJ1Ml8MDarF2ERIf
KsFgFgDhCkCCTp4v2Aid3cYcCZXz62wtAjOWmGQBpW3SVVCtBxpdtXs7f6hWTkgl
f+81R/iW+FgAqbzsu4OTs7sXrJQgL87n6KLXNuCvr8dI00CPc28sXuOjVLNoBqU1
zVmmKTXDxzRRLgei0RR2uf+DU+qMnt6fsoWYLGBnq3M4KrWd6LFrdIL8JDZfyhtJ
HJVYDAP++IsbY8gE616CFMuNqy7ApcG92RyrDL2IcgDtrpqc/Gl/3Wdam5LgswVG
jhpDDWj45ETsXPYWgoGKyrsSY5zOAjwH4d7J5hMVuq3DvlWaLlS9fGJvvg4RhZlM
KgPq2F6iaxvtKNcNAsZ/1bIAVF72dt3eQC68i9XITkZnQwWSVWDAD3aag0mM6WyR
nuLj9zbtew4XR3C9VsuEu+MI3EIPDGt8OXptP/QnzDTi+yFO/ke0cDyVRYvJo5Ct
x1mUNHyxG6fQSS3oXg3nqik76qZSO8wlF+riNRUgsrcrJ7lemTOblc/UATEEau1q
9LsvZIDWSfIX71T3dt9Xnf8Q3g0PHuWCO00PnrMpMxfe/JuZ1jHr8o4sGnLbAWO0
fZRbdTKwePDjwXCRJ2zNzwL7V3QEaIEy2V1qryUz9QG5YexqPytKoZ2qikSz42kd
bC0LAWG6nhVoK0/+US1GLLLx/OIkYDZHco77VJ2pZgjjDu/1VRfTit4j8MI8xNzf
LIyCzTtR7CoEZsAQGPS+bXdIQgWB2KOmsjFj7TigW1YHlxoC9X/3ZGMRQ87w9BfF
UNH/YkO+bCP4l5vcox1osVNsOoKoIdypHIO/NZ53afPh9Yiitzp8wQ1iZFCTQ5uQ
mLc9KPGU+v9tnyDs9kvn6rrUeI52GWXyWf3wferMsPAtV7zvH4T0/Rk9CuMMmfgd
Utdvv3LMkAkWUVRvdeaw0okA8TVBx0drEucGIjfUmSFa1q6QCSIPU+00ZTLejHxG
zoFxG55YpGoXs2Bk7srZBPqBV8+B74Fl08/B89GuDdr4DuUifHmrL4KKhCeIPLLp
WJYRvSVoL8C9ehVSjPMonf93t63rO1Cfbmtd6bOHt6C8vmd4nrjt4ojmm5fYPWkH
sonWQBpaL58vCYeLV0UAXo7i6QS43Xl5qlbBQT/Fr3tgktmDhd8Bpy/6EsBEWJBZ
c3XLhKLgPTcI8ANehPLzQU//QtZAEczAHEIfNyo5Jmpf3Z6n2p1iJQVTk0alAdMl
HAhGaJGOXRDHYoFjfw+fD1coWIKjQ+GIjLL0J4OgmRQNsntgJEdDy/zN2LONyCJV
taiEdrv1CxQUtKCesPqG+epGcz7ZRebpQVtsA64VzevP3m22m9FgVQN3J4w5YLbe
/N+gH9IWJP9ifpWja8/ld3zEZFk4+n0lWGfVymKQ8MRSH/Ag6W5poBpErzQ68N7I
SrI89pWThz9xgN/RBgmuldmbJV8YP8K+OCCsmuQau2zCZqaj9y6ggBQt0t3G5Nz6
dimABCVtuNH2c2kda7BSjWVUdJwW1YiL4mmC7y38cYUL/yB3ZwFoY6IIv5Etb0iZ
uh8IBLVuIyOwqN+XFNOryzsIixYAgog83J9SiCbM4dRj7q17lNYVahcGa7FJnbt2
Iraew8j4M5yC0PD6d7qopBYV9VW6N8BuChH8C7PX1PDiG7itQI0/nnKqk6lzmdbS
XEPtRmGQWS5AL2yn4nqkVXVUY3sf2nfTZbgmZV7W2N2eJR+QYlYjOA19LRps9gQg
ovNarQbfHZkXjFOG406bh2Kk9epRtjlQ6oJAFqzIg+3kSEC4FoB5HhkrbsbverfT
ByTKGXp+0AED8i6wpmDCtw/AD4E18QFM+4Osv/lJULqpy6SE9H0XFVyl2zNf0eEz
KQF+Y+7aBs3nRDE7J7dvsibILrYYifVF7bMEjg8UqhzlC26KGMNq4BRV4/5uuNuQ
d12vtva0XcE3fSjgOTohNJiOXYu75fCesFP/+IinNJZMigURBBPwS4kAgRYvRTvz
aBnASo7G9ROhSWVVobi6h3RtjwtfEB/mGWaXFxuhp3GH7ranjM4eAbpfJ7jUQiIW
IvO3JUVgylBsv53Iay/DSQwpsAuXxBehyaQ2ew3dXfnirsH/Tjx4jhVH6JYWQKOl
QsYuvtCDPeSZog0QOWCStlbRXQRnYMdqLqRVRIjeoFMV+Mm+wgZTZArODyQqMgOq
QhxW3ppzeAr6DjLfjgHHS9AFw3wUly27J6mA1XIKrPTur3kikqnXxAnDtEoCzvCl
v/IlE1tTIr0QB7nLgPfzvksb71oRwRZ8oYp4vp8ge1PSIapMFQPP2khDx9A8yI/L
Z0rXBBBGPbGcTA2YYhzUxJto0Lv6toLeZk0T8FIvtdYK5wFraTYrEZr4a1oB8f9Y
2yBOR3MkFCaWbevgzZ7O8ifDsdJx/+gkdaJc6cyIbCyC2udn2szCnO7blRl13mP2
uiJF7doUx/NwGYSM8keFIwUQnn4pOL6irZySLwE+OFzNaaoxmI46dQeKiuK0vF+E
sl/TC0RLJ2nB7DT25mUwDsxPUmeLcAAZstfNW/o30SgxCatqMbE0GCpcOlaSEE6u
IJPCZVgVi6C1ubqQB0grKX5IUUxDcktLu/y14E/deEMUDiP/npmPO+aWanLqhYj9
rnYgITI2kMkN3FoZ0O1kxIxFXM2J6P2yNMxldfOivrfsQjlN0masggST+tI3f729
8XNvbs8AoHXLzG1a02YUsbhcy5YizWvXb18N7EgFw9LZczpHg1H/NYMxSfrOKBWO
YCun17IbKxCXtU0eF0LufVPcyZY5oNcj/AW2VVWINN+91wygJorDWNjUNBarBM3d
JMtUvPzN0190AOUP41jy+cJxc9g47HXtdxKEM1CKMzjZKpz3F3D/x6EJby5KjT/e
KWTCoIi6tTwdby2nbUTT+PqtlV0EYA1fWjeChVwinKhAaXKZ151RX/MViOR7Sqwl
sAAHKQwfjq8daRWFFwlClyXf7bSTRvMqHxT5avkV2yjy1W2T/W1wEp+36AUnKAOV
AOV0RjLyWJ2TBpGkUA1mcc75zpWjJrCeryWsLkPuIW49DYukypHvKBuhUqspsQX2
GfvLqJhLyoumLy99F3a2ouIHpaqLj0NRSG0EcMIR9bla2wd4Snuqu2DrEjLCxXg7
CAWOFJIQfJv8V+YMlWdammgoCyC+8nx27hpVoJEjHMio30zIirqs50999F51L48L
IEyDmMtqwiNt93hm5I96PBsEEHPSdeWswjmIQYTzsH71uNaDAWABzXZhnvRIcLl4
Lul9c3u+TgnZWYAtkq5Qm4YR5iBKGdDKc/pWo3pWavLhgbSoYgv4V67ec/UBtmi0
Fv2d+To5hRfoBTmSecsOf5jgV9mN7AV2OWqbAGCCFfBympqyUulPCi4iqqSdOZG0
Usgseby+TChGC8wPxmGPITB1TwucCqOrjLCZSDbwOt7LvsFgQo8CaW69yDCNRNTG
LVv1gJNq//zm534Zz8HU+5xlmpMa6P8lqn5/EdaAKG9d/tFXPf1SG3MSfNkscSPj
Exzrc4mEla3dQunoYAy5wqgFIAxb2dFEPF2nelpdVgSUNmAuN0kmX/qcjGiL9hdM
AOy/QmvH/dvI1BjbCrz1rQuqIo0gIyxDivkydo6tjkU3UhLL+TBzd3Oqe2lhMhi9
L+aBKtSdVhD8mkqmQ0mK0gCZqGFTLb0WMTMct50X/Gh7fCCdNyDlmdxKyEXHklvZ
/uiAWUpRSZqUOJKg/Plw8dwz9NTmKd+2rRENvwyIXofrRbXdfj/qW81bFD8KHGiw
mfHgrxoEj7FPk9p8ABRE+PphlRBkZMED2NmT9DhezsKCpqWu1zlInMzweviOh7YP
VhV1mjS13LqWCJE15tnfQuJ5F4ic6HEAX80Rs7VFkxtB4a4ZxM9pWTNswdK4JIo0
5j4/QrjqHaSTSsQsuTgbzNF4hes9iojFf596rptrJLhxH9TZ7886o5hon2CbnPet
xSE2PAEDNQ0vTFXF9V7F0tXe+E4H9eDMBMAAgjAtJmhxweloJbCL8G6g3i59gyux
ROsJ3VMZPYl4Mdp5+y4nWwfiQcfh877lmej58YMR9AwNcCrtKov5aVVTchF4YmuQ
LQYkgGeiWc9RjjXUIToQDzjB9zte752qMWhU8O5RIBLykWV32TVYh8a1yyRZzD8x
G+4U0o4vsM57cJpqRPEegjuy/IZa1AwYPckYwqtzQk31AF/CqBTIGS5/CPLhpyRE
vVW1j4osoZ2XnikH1L7lw298gIJHH0uJsmStx8Bg5sdn4/p1+NntxurydJjo/DIH
mWCla4TAwV3jl/rQn8FlkGlvD8tv7ihOh35A9eJPASWjxLZ39MvZ4kwlT6bsLjya
ApFJG58XgIqfHD2FZfl656Ru7SWHe2X0Do9NahJblwrenFrN8UzNM8tG3k15g46G
oEX8+CXIWjE4/IeqUQQvnekGl+Tz4mibJ86OLUX0A6X/R8ta4m2ytKclG+B7QWOo
+lm7pWjMKiQdu17lXIr+aLKr0g2omlDzAkrjW5RfnbAxqs1TboqTP1P9VL9phTdw
Twkv8c+Tf/mltn/GHcimBRqbCWAX/SEWqiFQjPR7ZW9D7yIT8YwAUNKQA0KUcg7Y
f1iw0kxV/99CKppOO+7fYDbyAkEI2BXHN46U0f37pyVPU0nH6RrI9Cu1L/y8FT3b
ZOHyi/0/iOaJ/f9PaGRWIrWdHqVk9MweTgbGen+tzLLsHUwjZTJlsMAnv842lUw/
8RZSNcUc+qpmmnhCxiNLD2R1Oybuibndt7uS4zzRlt4yBTkARfyBqaxByt5b7bpg
o8LXFPOrVm+MdoRKNjRbC2+o76B/v+zUGuDKibww6BsEbZPVAIUhYb1k3bvgi/lQ
6Q3nFgD2dWYz/xqFT/m6SryAAlr9JgfnmYv6QieZ0GKsi012hYXYCA6j2WQKwP5H
MgsnrXsOFrU84daXZ6n6z3JkRmBPgglxHFwvTUGBx67d9V8sgXjNtrJKuJ0RnETM
JvIcweFmmYtXegIXbgukuM+pYvussbEFXQKq9IkNQat6HvB9ikGcHFY0IhwdVbxy
BXUEODY7PIIGEiKwpyn7qRhpDAUiV1jjS3AfVieoZfWMvENzBboITcJ+39MYZ3Dg
XY9ZpXMElF3cRh4uoHK7Uj2qyZH9HWzH5XMBVn819Yp7LX4KA3xIS61u3ggzTn77
Sf7FXPyEV7w3InfnGA4M6TLBYIzaqsU23C17vT58oFFdSg5VyqZRRhaHxP5tl5K3
YRgiZ+w7M5hSqQ1zkCYlEE436jGKodleqPcxIaqE00s8Ioj4qx7KLNwojosgvd7J
ESdFX7jrpRi8rQGvqro+0DRFU1RU2+B3+8dAb61CDqyNB9SHHR6k6HjQ7w/b+XwH
HFsBk9n1aPbQY1rmnLIf5NOaUKyyOjRwHxZxKIyx3z/K7c7AmuDSQWc/WBCFTBe1
h/fy2YJ3gsAIqvfnM36t4XeRmxAS93IjnhjE+vs2bZbVupjICZ2mVZmeqn4DIRIA
XRF2Rce4x0B46b7zlJM8w/Fc97MYMXYT1/EbUqQEUlzJwKXk9AZHl2Qrq6w7Ab+2
lNYoyIC4b3SnTVUEo897hT1IAhAw52RHRaz9NbrcTiMCwpIh3pyT0xio4qDh3C4Q
GEdpf+uGbtOhXg0B4hEDlybKXEsldU7F0cLgmct1Nk+hMZC1lW8n2Hz5fDRSIug2
coZL2THfJdp57knwLrr2jqPavs8v5ek32q/ByvpnYgkP+p5AbgNCyUoTUCTQ7Hz2
lpjA0HpnFCmbpfqX6EUkm15lXOyK4t519smTKbrkAL6Zib8ZQoYe+2675DHzDxzx
VJSkTEiXMtjBejoXTyIDB3dcpyr5LQPK9BTyy738WWryR4H2kpXSZ32ogUH85ldA
gV9Hc3pLnfn+dQy7lhnxYyLpuylD5kJ0bTuZnT4PSmMdjbyr5TFJbuSBCLhXa3wB
yiSCTPVSePLn8b5HUC41fz5sDgJJlX7MvQBTxgIQ7hHJHAqc1f9knPwOFY80owS8
Q4XzQRbEnMz3UjatSmSZwiMTjJA9ctFc1c5MwGtRcxkxtD0Oisfrc618IZGAxlo4
4wsGz+Uw/RRsmhKSj6XL92vnm4rO/U62IV4MQ0DcT9WFVDWuYQXDSuliqGdF+IqO
Mg0GJZTS6R5rHkaY2yA0xyN+/2pOfDBIB3UZ/P1/sg4T1vhvDupfARNl37859xfu
DyQRiu6hQB2RnP52HWUHPuhvrXESBF2NifyqGwdV2e4Ey7znWwUqBJrBNalg2Xln
Y309cDFtvOWMUn8yJlUFQqEpz9UZcrh9WLFgARD6hvnYt7cCx6B9TQIQx41WSzRS
JAECQCFBbouE1X5LkHNt0tf6+f90Q9fviv43STD4Uh7eeg3SudFslzEW1or0u2wY
+ZWdIC04/baWv05+ZSoSH3ztJg3XbWYQ5iOwkrcg9pR81WCh5zI4E94Mhx3/b3G4
jmG+l+fkQNBOq0YLb+5bRrhn/qzYygsxFXNPHfiEZEcPxtYwhX51Q3BZC5WNtdT+
Ev7xN6HQnD6j8XtplAkY7fxTChLUrvc/jL7QqLzxMc4e435YsdTzJT1LdOGLc5/Y
6+Qshl34Yun1zAYLlbPZVpRzbw1AgltkEvuESFO7znA3W+IEQsEKnItxM0idJj/L
qvGCTinf3pNCOaJg+mCbQ+eM28QNcNa4/mzLenW/cNW13UmiaLtW7Wooft/s8pkf
WkZHwMY8X9ulRhDMsnErHsN3VGDQb3zmr6FinSmyFmM56Iu6Z77sAUxQskY2gWO8
udAlN7VdESP5533SoF50GdCwcysgqPpULXSacZsSM5nOjdoAit0/Dwgqqe5WBRTG
GDM3c6DWXzQTdZtIB6Mfwn8Fkt+IGBfGadfpNS/B/gaGcmppIgPrhYwRBAtH9XZn
1CcYy1MifHTZ7t+kze5JteNEx03UTOpeziYB0O5/Jl4kWYOknYHk9bXnHSol/yed
KDjJo6kKQkmP8Uf0xPYAGlq6jkbpJPn8Yy+prRKbv1BTCNzjISB7F3/UEoLOukmC
eyUS7QblvnxZuIpzOozR+tHCmRaOxs257qtg0eX7IiUUdjJROU8qr5YVKL0osvSO
GRtfeWP+AkOtzHY+GazV0HQ1+EikqnS+H622GIJjEFvLJXUujSvdikGil/vAUcxG
jeMVfhjinQ2OLdDIcOjI80HGWnOVtaoF2+risznfi/cCyqWtH0H7UNYV2mdM9Mu5
V/WqlV56SEjUMqMBlJkVCbmZgi5kMa6SWmWk5QlofsLAp7lTLB9Aq2ec8Uq/XBSw
30MIUCAs7RkCPuDBiGTBoKpngSQp3v3F+FN2c/WpFkkozBr+63gqudwOm3AC7lAX
0EYAVItoOXZ907heQmRKtuXi2WhRI82t1iqhIjUDZG98FS+s7RWFviP2BJOe00Xh
a3qg6sPRT76tnUquwGENHxagSDhvB4PNQkO6vnqqUTYL00ZvHKaTQekDYh55MZyS
H+Ax/jNzq4fHA15LrnRev2G9ZNbkjZyXI+CRW56cMgF5R4a901UpZyHMMSd05qSR
fiLXK4IFciVbnnyQAk+4k8NYLn9A071wEcGgk7OgEZIjZQKUFjVpGfEqNCod/yUa
v26KwpZNOqniEn7J7V5ZJ2pE2Balo2Rkj0MSOyFUU4M8TETBhVjG7/BO4RfG5p0Z
Xjy7B5ev+WSNHl+VWjVk9hhdsVgc2UupHWrUeHc+I3QKs7I0Zo0iBMJSwAs4U0LI
lM1vvddts+zFvWLnz0VX9hlfAUwFkRP5smKBzYkdrzvSG35bLs+g+r1rnM7bkR25
XX9PD5Rs9KcPBLlHcyGsKYUKbOMPAkl8CRcg/zwpVlGnJD3s3PmZLM0u38BHXyxb
HIieBI/U/Z78kV8G2TLO1mUk9qOYKxRVKALXyb6+nIpPshD7GU5WjpFW99VlO2vk
Ucibj/XRJUeX63tymhDV33hrH5wIyPsjCBd7wogvOGbN+GLMQg7OlDiDB7jwHz+h
lP8Foks9CsBlpnyWW8qocjlYRfA7UywR1DOZp4QlrXhMx0/jM6ncKPX4VYdkaxfS
TL3SJkIIhu3YsLmVCy5GY7WKGpAYUgMd9mxIFDaW8ebpzmde3xhjXOGbK2CsSNaq
XoifE+rleF1gFCp0MWiVNkxsvXZ3ITjDw+E3X5K6m8N0ieRQ1FMuAqXN3gaDoZYA
UiPUh1RW5fgT0ujATWv6MTAii1Z+OVX7IVp0r+c8Bi7+5J96hogcfZN7rqVZZI8N
GP5asWYE6PJQd62oqpzzwsdZW9nJ4LzNkLJCAPORhYD50x0bVKyUt88zMmP1Iy5p
F6LpB9NKy62zfyb8wOQ1o0u4ivBOph9JvVLAJuGDL7GjIukw2Iuhvw1ILMB9kl1c
pfXsd049Ny6D/GO/jitySPQx5aaDcvXmCLrHhh0CAW0AAo+4rKzX6Ciq2LE0JOLK
oxdF/d0ZMupqzehGkyrfYROXgTXwfQQN9XGCoADhBA82dGwoPLfHu/qp02IOHiol
eybdrr9l3+Y5f3U9YFHJdFWWxhYB1zm1VhINeGMgpjMROnw3jc1yEZo9qiKE07rs
CFDbg3wIuO8oxsJIb/47bkFq3dxnwjCfGFm5htCez75tD7MAOSc4YvPqmGwqIezo
AoA9FTKH5l2uz0rnmcA3bEvA7q1jPyzrZAR6SfPfAN7PaEqO1RkuF8MBdfgQqunz
NQx/oS7n6WwfxR6gmP6gfEsMUzzBDu/WpXuQCc0SPyXDjtFn+4C9sc2swJIeilQU
YlY+iUMSCQwOh5DBHGnGmYwyCTkjvLu4/tTmD4fPhjVO2GCBUH9y5HEsftqttPSC
3Kz0jjXLMlJ+NbGoy6k4dZzEC8SotzaqOrc4scnhKSsEJStqVtV3jHNmBFjpTLZl
4JfQAJJj6AKa1QLHxxm7Su45qh6yWL8gmMbxNoAq/u3DENe2tk75QSv3liAoCJvt
c29IF9kJ9h6v9slfvze8u2cA+rXJJETbxG3Zw2KIXXEf/f3jVNrONud03DW2+Q9H
iC0y6srYthXJgfkee7mHEW8d5MeTvDOUB+OFXGnQmGyFVjbfDn+0SiPIyC5/xROD
N7U8uUZNtjLSZzkAyTaSJa4yiSuyG4kOWjGfgVBoOp+xJwqg4rgZUbMpkPVAilxR
4HKQIv8rroYnP78FMw0HVwK7kRyQ2E/GaiFYb1+iTnndd0bFUxQI9pj4kcFUhZF6
no2GJw8WqgFy9olQg5IEKhelDzSvk/56X+S1XuoKE7FwRJ+d6qYcdT1t3J/vL0q8
c8bMoVALGUIQ7LHTv/BwkLCWJLLzEv4O46aP1gZXzRIjA1klW69RKDps9L1oAjRJ
aYTXmUShO2j77V1Z8+45CUCyZ2VG1BfPjIzcs1+ud25aTJZK/WOgGdXfbRSD6PPs
C/jinsrp17vxgRAXUNZVbAUgZFs/x9iu/OaQ5i4oicdhAcDyBepIlSmKefLktsrd
a6QwTYAb2fDw7zU5KHDehWYEfeq4Y+im96d/PDopKHYhL8yjBx8pj+wPbHVQBU5w
7OOEvLs/Xu7+r3GxVKZECN+KaGz2g0egrnc2GfcJV3TkdOTTlQkIq3vuOcb7vdQl
bMHWKCMpagEO4L4y2NIx4f1ru6TBfO88mr+uvEQGdaRoXsAcPR7bkvkkuhKzRH7z
SQNmNOgppEZJDz8I+ixzZrXk73chYNUwVpvg3FGGUCyNeHUma6utedJFIh445TSp
mN7VYICw6dnm/3itvo835iIo5FTGrE+Q5aTScdcotOUZbs8FoNY0rCNh6kJF3K2/
O14DKzY4WIIWFtKdQ4vyIyu+j2PQlJn8ctiG9zYew15urnNpBY7lubrB9DQsaHyG
pLyzIIEdNSNSpAEbqFo0JNEWqcd4M+HtDs1k4uGwKKmJNLnWboQEFxGhO8z+zLqV
gn6IB3E4O5jAkIgehPu1Yc3zzOLIczt3kXUXoMIKUooq2QsjOg33OSCOx9JWXVLs
Md0iIJGxKVf16DIGXQ5u1X4Nvxp836tWWbE7EQOGBJavpgPKu8MrD3aXc6CvqRrI
61iprupYWg4XRPHOH5TOC8U/4c7YD1JNN6CSk60L5HjKwI102BB+4AT82ybstqJL
QRL+jJaJfQeIUE5FmtEhi2M9uVLB668gSoKZpL7r0GM/sKSFqXPzDcM6mB4Ty3px
99ZHPvksRuMjFKIHDvBiY8eCGm7nE/ld1qOu3w3nNAks4FS5go51nxCBOM8pQwq2
DG9xKxdmSPETLOwRIrnFVThPj6n14glQW+t2sLZb1XuFRzPp/Nwg8yjjMJuoBOuU
xDHlG1KdQOjfaiASlxnRRilolZd6sj99ggMNVgHq+tk5MtrXjsx3RgBxUkPrGDGn
S8GypuF0I2f56d/CNsHGB/ySUGIhBFmf3X+iEdx5hS6OjOEillmrdsG89i+aA4aq
`protect END_PROTECTED
