`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1aXo03VBRwHvUyWXocBpUa5hxZExxVdR5MKzroWwIBGlb4cEjFtkyFwRHdyUw+6B
CmdPEqOwJhlCJ2jIcLnVKDwmWWEM5xcNRfqoq4wzNiioOiq8JxWwaL4cu8XQMh5L
46wuvjMZszpN27jH8G0iL/U83Eda4CIoyBEWQJ/B8pmxM8r1mfVI2j6CmTkwzZNa
yZFWvF7ikGN/lvfGTtZTL167auH7+r7WQLiujk0LybQXaWHSEafDOCUpgWBU3Xq0
1Zu8Et52eXvvsXBnh97/Q19Iy7mPUoO9OMie1S6X179TYHqd631IXDCCpMXVbKLm
+nps/Qbe/acQI7PoMbpfD4sxMhFQXstXPkwO2xex8yqU2rZ8d5no0NV2A6lbztWd
vg5v3No77/dal0aTVh797/NPnJUsiSwbvJFSaXeNQvH5X2QvXZRLdNYiy8mr46sE
LZJlaFZ+aie2u6aCg1VD8clhFw/KkJS0fPbrWvZ0kiCcz/0dOcg8NGgZyKTd5Ppy
8fwzUKmADEU/S5IhfHggp8nVhTXBLMlq9pneQrs4mquYnQ46qIepuc8NWISUD0QE
HFVlajFd1QWkbzug0lXRImHqgwraR5NMTmeSc/CsIDH2kTfrZszQAoiZsSsW+Lpu
9+8mbLLMC5NtiLUEANGdfYoXYcF31HeCgooSAT2zRh0JrAQad081Mj9b6h/05Csh
bAukqJD6soDU5fejx1qo6iiNIaQqTWW/2iHcqJCdLMgBTz/zBDMzx9poanzfmJKO
YZU2jFGqmx6i8d1zmTABeMb08TSMzr3QqT1hUyYhDACbjMXQGakaWjAzoK02VVyK
stK6HmA1WLzUXC/az1MzphZDflPOXvINp66LEFtMvmxZ3ElHwZO+x1IfskSZFShe
qIv/Y0vrZ+1a4Lqw9VB+AOyHWSQ24vywPO2qZcR18PZW4y30bw5Ndhgm1WF46HY9
XZ7u8mPR0McAbkZSrYtifD+xltLRUGiCThILP4kBwr1b6MKhAKYYEwPwJV/Yduf1
SQ6U05jXrbmypnKGo8kUflNDqucQ9VD6otNMcJZPzHMvXhFldymI+T1oNXcirqDD
aOs0hgQ+7GfKVN4AzZZsHRaPPeK+RA01mcaRExS3s4R2F8Q8hCoJLGiNkSqethch
CtxI0E8ktLmEGHIbhsWXPGw497sKkWvbngCDiBWNyxUZy0lNnwdjyya5Zva5ZXjY
NIdW4W1/iXHuIR5H7hTLf/i+Uin2DCKywr380EGjDsl5yJiXQnbgZKa0aUTCAjzR
P6UnpqPbQWlcqFWF2H797JT/S/rjxMU070vcyb6C0qNfvRnjsXkJId4hxd4b7vkJ
wsYQkjwc/m7xFGztoetfXteucMivMG25SVUF6ykM3crdzPUHXP03YOTelt1S0WNU
xY+XTe9aGTGcTkblNGfkfZj1atTMIpArAgN/UpV5yb+N3XBan2m5BE5S+rijwB0M
gyAnbwELVJEF1YWRl/4diaXiiAbm30uMo1zOACFWrOmtsChalz3AxAQxNPbxdNv2
xQwUY4Hbr+v4sKQdxfeAmd9oyXdHqTaOsw7BWHKrJvs1liWglbNFq5zUF2zqjFox
MkutQoLU++hqVBEs9Niw5zt4l3eZO3dNy1t9UVsjzafe9sFLeovM7rOC72y48wQq
IisGYVP5DbwPfeo003hqwnLOjM0po4CGNW2lxX5NLp5UvPIZaEn/G5OKJ64PvUCE
ZLM5PjEj2hHnNMiVtwW9P+1gKgnQPXP272G2/jwQbf1io4xYj7Ff4gvUM/uWgNCk
drvcrWMALzYsGXXppII+8PueHSQKq/OHFiT1M10l+sfr0AygCxxBmkLpIcxAlEQ9
7DPWC+qsKYgzzOqihpjqgqiYR20AbnDfaL7LbupWUAGkQOsNUcBXF5bXasQZezqD
845Zon4pLuFlbfjqLyfU3+RELHEQasXRuxOG94exoG53PnQxg7gwzl2LMD2guX6G
ROQGi3+zVjTmSPIbXSCZkDIKr6CDwsFNkTddIOW2xkPUviRajqWWKoZUbaiOyfOg
jjim1xViGOMEqCOynJGS21z0SG6v3nNvC1jZBWtPcHCLmpZz2AcP0uEgUJ9+YRvL
bKYfPpNe+dx4M994uiUcAbASux+STst+xyEejEf7quTCDYdyC/ZFMua3LTfmFvFH
arhRSltudwegAsp3kR/6psRe1NGpQf+rDtlLxPCOAl8YZUIldvt8sM162rd/eEJv
nFR9BvT7YLBUd+6asFq8yn00jWhcMMQxjRxf5Q/2OEcPePsyKakR+6QtHr0JMhrW
YpjfxLpyPlVjvc1AOndG0ngfYjL2Dm7fgO6qfyQfEFCGrT7a5CmE199VUoaEM28/
PVqCpvuduIXuF4ze/M6KaOy8fBBW2Mduzp59iYrxshMI8wfLjoMc0NWe5ZhwMnTT
YThwfmb12uFw84xf5UXEoPRWbvsaw3Z8WHVKX4ivAhPNWezj60r5dcfgJfPd1moJ
9Deg3zHIRDS5BAejQOpcAZUIxFxke7IvoLu6mwOou8u2u8ai5GQMnrf5Nn1KOo+m
HKFOAeMCv/8TD50mDy5dDCkRcXlZ6Vydwphhf3F0wbDxiWHBuX4k2IiftEQUJezN
ZuNHXKXf0WTyckdsPdP1sTquqx7NPZYh8LKj2y7VRvzyuEVqTZalItNOtW1Jx3u/
J0FMkGA6kk1ChScxcQMQqIehYZ/Ge5tViEjfyJ9y0UcTJgJ7A5ttxD1mPVFyOzFP
W5DNzriEFzYkjS2z3e9rlEcCIhmfMkFB6F7TWgDk68lFQivhnqkONKR+v73OxCxb
QnKoWKkifZ71Cl1IzZ/pwU1HpPjpTc03rIxkQVo4ZdTX/D83ejOEumlLOn7y/U/0
eQhSjh1u56X6HahwHPAVoRlQO8mzHozIoeBdLz3H9uL5s/ZDNXQ54DxKWWXSe7DB
fzjDKc/z2024QDbQcBKEbNb5qpx8/SxhA/sYA+9o43xY83n7EYlzR5pqZy2d7d+S
ed/kjwzhnsH1hTElo+TXNxYcNkNdwfQQpPh5MwDaubYkHcbjrPvWlQQCmtBePtT5
lZrErUmbPBEAzaKX8VaWV3jrAzKkPWzcdzIlDr2OwrcIOZBs1eX8+26cqLsaGvny
I+Kx1hVh2DCSnwmLau9QtOvLtC/ELQSQMiGfDb5WyPMD1jzgK8ioa5eoBquwUhEB
SH4tLZzW6muL6LCQ99IxjqVWhjGZBL/hdYkzIytj1ndGmmjesWb25dH+HGN4RcT4
sGPFzWQa+vnT2hHtTK9RoF14BrHk36Gu9fW+U8tUFs7dVJ9BoM/LV2te5legoOlY
7G8FtisM6aQex0VWnRZKtEp/SrumFl33uWJNo6AIOvRA/5eJ0XLReZdbPd97HLq5
ln0G6OEJ9/c645QlnLRrkhRzBiceFeh4mlI79W2iETCkoo3GdWmqHXt7N1AVfnC4
ZGpfF6sVMyx0ujJ8YzkiucCy2j4JVbs9jFL4PW3Jq0vFxyjc3yiIulEygjVdj0ef
wKpCvRIIq0A0Ve41G1AaO1pTAAR3JkkgfjEVeK/f2Uy+IPw8AzoBs9jD9vnIGcJ7
T0VcoKqCK9rnqYLAFQ2Poe3g8Xd4n5oof88nBsoKTcavD++hXUF8t+kVXbD2Qq2F
EaBqX+8+rJ+jhur7JSZlVc33sSkAqwkGDFc1Anxj04wq3P+B5aOuVKmDseDzi38u
Tf+4SHlmixferWxxlJHKEhEhQH1Qr0G8It1jCepya1crgOob6/cyVF6BUj31PFFj
rjpad2bOz6bXF41yfuyJ4hqxnUQTSWhFZ3gBbnwM2tndHkoHypcalMqyGchMi9vC
hxTmWW6dgOkjRapUQg3K5JVjMcf8xgu5A5UrCaL3PNEvBAZPN1rIizWQSd6HEyqR
PENv0tnHlFeQ77YZUR2DXEl19gFw7OhqASH9HeyKKca5hqYDv1vz3XM4Mo9riMtr
Fi87mxPIiDipweUamBtjrK5XRkYRZvF61xT95Q9ntmgmQ5Al4jPaF6Afuq2puBXo
Qqoenu8uumYozPDZwy08lYnALHvU1I3FE4iZ8PrN8AYsAYNh1w8TEA4Ego6GeoUa
hhH5yBlGFB9u8v+DTbnWLX9zy63987zrXYXB65p3J/wz6lrPujP+lVa0hv8jDcca
Ypc9nb93+ySrxQyy+vkrFCbfE9aGjikSntm/zze4la2Lx8VkbMMGMyh6w+GHCBhW
lVG/u23ER/fzKpOleAu18q0RQRB+RXKa0x25D5rUhW581NwVioR2HS7AYKGu1Qnp
nNVI6GwI350fPLEv9yM8tlndlHNZ7ZRYVuUuBHy/qOrmxNdGLhhDPJ4dU3e7Qe5y
UfC6rhnsMv5h41034VUgB8yoafetNf+BOW7SqEQ8N22ZgHGKxbb9f0QjdWU1Vk29
CZpjB6oIpEI1SXFme8CZTcb0frytjyRUX9TXJ6a6nRJXPkuf0iepJJtnqAHLUDzJ
ndh+bx+7nIvfOjQoqwqXSu0VUBtcLJREiGZo1wZ7Gk3Ch/adQjnE2yxiImPiyt+q
YiihwU4IQU/v0t0EXSO4nV6hTsbJsb1uYOylPY4RMaYD1YikdSDafeeMi9wao0gl
3MtBP2U/yt0vFwLso1SCajQdJmm5EeuBf9jbufn2t/qGvmOjUAvBB20uSMUhJ0oO
Vs3oUhjWnClI11HHKEfnEKBLu4ckTU8Kt/KKFvLyw613QttBi+oAuO6zI55WanYn
FVM9+Ey6U6MLcE1PpeY5phaxl9sSDbn4Y2STY5LCOmBkMgbKTQr4vcdlEyjoq0cE
UQJvUZNwTEQz46Y42bkn+58C85NvFiBpZYqv8q2uOlbViyww9sok/p4Gr1NxDcCw
FHFy4sKrRRRiwvxPk8lq3ACTrSGS9/sKmC6tJfZrPYnIKqJhNpBbxGSoY8CqdCk6
ahvIB1Fe2IV03clLpV+RBW1yjRyF7cfZX9NVVJQsB3FYFUEtbce4lvZwhDjc486v
XbiNqzjnk4P/0fx/L7hX/wXBEJyt0RXG/qfXKEDl925v0UPvWXY9rOKmM0POaf3d
vD+0oOiYJa3ZHQoH/T/f8Z6eimbnOff1QWos5XNebV6spWuQJlFEaq6ckjR7mDFw
87G2+rNXRlIXirNrJUb4b6G46qN3/dPoz7HldrO9UbQrRAmYG8f5TFXynCVFDewL
QDsuVexbwo0YTHK/L5AqUVj4XWT0UTVJuAZdMq90YavqwSTgGVHsnQfv+ph8DPDz
5wKF4CtYZBRM7y6iBQg9yYXwwyKGq9Aqh8XERYvmvNV74Sjf1vFsPe+1c7IdqjLW
IkZDNiKGXeDkFzFnETXQDdgBWnIsnzOxGxZn/qfNMh9n3fd9xDBjEWjWZgI6lljP
oGTps/f0kTyYbJgWi0n6VLIufkicxnOg8JoKy9i+zdUPZSYC2z0c56giwu4kp1Rt
jKqxXvXvkb2ZRhpnKyB1Uu4Zj0VOH6JORNGdCJgqOZgAl7kKNG2et+Yg5s+nJyfh
OSVAGn/4OGyXWE095uLorZ+2y6DY79PSdsO+okoZYsfxG3OXlek4gplpzxdq6zEf
lXVLeIV7nA5JczRQn7OvWqjRSFzfN3vIlvtqao9wJ3rJqXEtHZXhXpUFYrmequmg
LAmztQQBX8JLkcRdqaUtlQ==
`protect END_PROTECTED
