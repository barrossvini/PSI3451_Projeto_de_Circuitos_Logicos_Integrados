`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NUe0m7JEmB3D9JtdJKvOL27d3hD7Zi8RpdXJq3dVH2p/OcocZL8gIL881mwMR3e/
wnyOpraTzWDcqVYEW5KrwTSKNv6x2sCX6iC+5OX8URP/5p9+PgvPJg9Htyp5RctF
ZHmpRNDm/IAGav4OSGs1SuddG9pKEKsKFM2Uh/KoAdVvI30VYR+ZGoM1E5dNlR83
KUn/SDTD0EwAZuhI+B7Q3+dWD/8YL0JLdVjjJqhd9LR83Bef9VSQsHyMKZwl/Fsa
PGMggn/05jbozTqdQJvzgydjvq1EhL6K7ySVrx6GKaiE5MFi7jWiPVkaFanH6Yo5
DEv2XpdsiXrOlnrfZwnv+QGGUlw3dDg2J5jyyLLfKNBkrDtanSxyZhVSckpF3Vse
2BPNTRo7O+V7tPNzKbrB7aIOeAGi6QZs+V45+JDEPVBSS1498OShZQx5mBHn6KM9
auKFthxDBbTeRvwUg7CiMylBQ5cxQZtSodOnvsCiREK/5+dSdYH/8omHvleL1LWs
gxEVICuF0srubVug5wdlHZmDjc7RPrv5qLu5bY38Cc2ExvPcpIJYbWx+R2GF+T5D
YAnw3FFeGcpP0G3Ebp4Es9YcSeSmsCw3StcYWKhxC83hglrUE6pO5oMaMPEdkckX
HK7jgMsAvHfBzWOZDc79y1uNOSd0pF9Lw/CILR/CffhVjCtLfdeatD2KMmI6Vn54
V2x5XOKGwIMUZSU6HixE5vuDfV1lSzC9HkjT183Ucqt6VyFbmYvmk0JjgFZ3uG0W
s+drg5Upgy9rIWJQ3aDhx0Pk2FDnIG0wP0cVqQKzSaM4K9wJLkZ3/59yTfg+zQ+K
PxgEPwOWBmcTvWLgEGb9qgfiaKetM+yxqUyd7wzx5FYq5OFS1gzNAINcOHa2kGTo
iEOnS3rohnQOwBILpi3FJOQpnJ7Y5XgeDl6ip2Vdjhei/uqK2km0IK38MIeQ4JpP
gfevnLI9hG+L9L8zDLrTmyaiA+2fGR5jA6gLRZaPrOpbbIibOxAuMGXwRaqB8TwL
HkvWgnLaI2S7SDefLdeSPQhgtWmkuSP7eLQn3xhRLScFM9xgxjDfcI9uyN5NIfUX
exUoGOeL+60aqQdXJbHgY21hov0nalZoZWvEmCrXpj6U89eyxwo2Scu3Xt2gJuhc
x3EE037uQhKBQrYi3hI4N0kIi2rkDAObU+QT+ZrLYHD9cqhiA3irCwqv/GsGEkiw
XeAEYEcZjNqVGAalpK8fBbCY5TUjMolOQ4DBNqiApMZfcdfjdpGos0i4uS9JSR3J
gP+LbhmwQR4hX7MBKZHllB7xoL1eQBJljwmAQ2dDGmc/Svh8PCYfg7VZC2hdPNMm
FYuBBAFk3TbUIC5zLvuu8d0IcIvZoUFpP7qcb+YGPOThygwRYPOGdGrN4xM4TTgx
gvHurFtHYfj8vccKZIuZbdibY+W1cl+zA8shbReKu4zTo24TtjqRtALyBtfqcew3
DGmnE7oYTZy2j+wPepUxRmrtcge9VpDnuHTfnzhBV6BRfZh3hyMUOF/i8uTK5d1G
4Syfk/Vs9ISQUW2HGHcP8sLubHeXrKhbHZXOG//ks42AUXLfrhByAcSDZmhm12P7
JGYaivUhE4rLtS+1U5SHIMp9CKfNpuN+bM2uOxCa+63v0VbDrqxVZ0y9JV23/KXx
6NEnzpT01zgvJGe9APPExX2bkRwsjCb6tY4YLUBtYgDndHhavPKuNIUlPWt7PXrp
aaGQQ9QOLoM3XWEXbUoupYjijIodJrHj0WLSZPzTtzq+el6HFR8F0jZSFou/F8yN
DCmfzOBr0TDYW2PRwkyV1+TdWn8YGQbR5kWqlu4Uyuz2xSbdaZPj04RABP2rHfZX
xpP0UNF0EpMxCmoh365Oqus6vTCtMKJ8Zm0v/Qgci3ZgLBzNSTRYBlvkGDpP0AQd
p1eKDRpfNbrCKAh2ybqq6cmxmQOwYW5CHS8TUV2n6uTPBQ17NsFfRPePG+WrWk5L
0hC9AsZFzRfApwkaZ5Bu4nnIUV39hDtOOPXZMQ1TEw50DdisMhRZO1A4jiowiQAR
ljInKyeoSLHqFinhhz8y5BiMEBWPIoYJyYYhx69BUEQCRrf0cCrZk0qPg5mBIsRw
uZB7W/IKzAEwbvTDEAIEEz7F03S2niP1X43ZC19sXxTaMpVG8XJabgpks9q9WtrF
tw1HZ49JDL6eEYConzTrYlJBOMX061zDmnbdyWsoJZwu0pelnNwAj+zzKwvZ74yb
YgrQzod9n4MP5lnV0bh/1DROtOxPXLqwVGRDq23RgMXKC6BHEC4kvlx6iYkWoai1
shclBwaJ5N0bjzaKHuLGVn169v3fZkn0ZX83H2wFJhvUya9qqJO287tZVe7LTTAt
0Q7CN+ifrk7GyiDmRkKpugEO8K+RyU6r/AqzCK1lnE1WbiOMNfOomgbpxfA9Za8G
CtMgjDfbNLsf0yleP+G0A3rZRx/umYbjJq/PntiNg2iMUDK0LrsvYWH64FB2bVXs
EOQbOyDGLAySP7n18q+CN2thUH7G37m2QSfdTYxvyVG6My4bbNwC/F2qQWz2n9nN
1CR5GIq71FR+yWVSRduQTkwPldIf5uOCLtQU8Cs+3OlRoqDH9LvbuThSv+ArWkgR
DZkfhlPI0IAe+DyjyTKIpdaEFA9zbiFHrRX7hIQaxUfFFpyhrubN+aYsrAaCyT1e
aH4uReNYfl7PyfPLSvNlyV1+ZmgQKlY0OSTa9K9/E6duUkHucZz5TYPYbBYPVGiQ
/g1Hh9b+a6P5tSMNJpnAYoZI/GCiWphg0KX/qvESn2A1xgmMads3LwpvGYYfF66Z
8+UMAZeECWj6bFevUzTW+U4LjIi4Week3pMR6A+GGnLnWxxuvDMGTwcKE0yK0AP7
d296o233U5Si0HDdNCFDnKCt47nQYpilvPkblQ6+upUzatcSQ6WZ22ZInvLHzTvi
b2tQybtXypgyNLNqHAIiiC5CN7bccNE1MuPqI3rsmRffoZ/134LVlp4wy3O8Yt7U
e/GwMA7gQ407iqe9cLTEgiqTRRJQ2dQwI6KjcGKpuI/Ug3ghAFBEglk2EU8NetcC
3tQX7vBr/5JwU302CrT/uQXB6DIFrg8PgpG4yXQIm+q1Gi1lcZQJs9dHQFVh9cwK
ePdxdtftOjCI/jkPaObYrvCMVxZmHDM9Wi3dDuMmckk78eftzySi2c6hUngPG8+G
L0Jq1ds/vpFnAe34bUzdf/UK5H/WMVuvoTHOBM2Urp+yia4E53Pz000rIbIn0mkM
Oq6wP9s8y/5qZjClWOitcJmkPMD1f+ZddIamzXXMLSr7163rivS+PVBKbZt13RDx
Gtu/Q9cbsKi3CNCW7qQ2cwkJAK2IeQvT2XdT57fZQlS9D9eQrWXdbd+z41wFMzca
gPIa9w0mf+b7VbqSvqWl5EE6P5tXfkkn/t1KgQ9XlhdEE8CYlLCGqcRk7boJ8rlt
omIZkKut19VZJKUUUCoO8VvB+zBBsQ/ZxqIqWr7ukpDhvd/4WS4Y+xUpG6eWF12q
CvzkWT7f7gCGnjebKCi2pZciurOgIxnmQsqgBMcqeG/17pxnmsa+2UyGKMIZUx3u
zyQfJA5WareL97J7nl4J0Nv/JYAlIiUbHL13GiZjRruee7Lfv7t+hR5Z8JTDVIjK
hbKfHj322nGfrT/OO75wqU73ZO9H+F1TPPpsXfGiwoppLMQwMEC9J/XAWVTjskAg
MYuYTeTr49ULfYB6MgxQfWxwFa+bc8h9yZYI214I2sPoAtqegHBrpWm4sGqH3rwX
mSdlhYnX3/sxDeLetwoUU3SDvxF9cLHlBqVhEbQ6rMBHWy6pfgFAXvKoH+P4Sdlr
Iqn95hasPpGjhPAe/GqdgCq6zZ8pPCWGiIvpOqgp9JeixHv6fBmDz7Gnz6Jc8ItK
h4ey22ybZk+8dxohuyK111ZDRmXaY73UdA+9CrWlX0f01aDJfNA8n5phyAdOMeWi
o9KkPxfmiNSbmhEK8IgD7WJQLW2E+Ggtcps2ryv5YjHRybVvxR5KDW/whXvaWqo9
puT1SmhsQkq3xVTnM+Y79JYAL2jUdLnbmKfaqPmj0ShAazQSmiCWbNOq18MiASbz
m5u9N6JNGunp/qQ+gMjxg1cdbdBSCAFUj6Y4yAl9ROIHiqgt9j5TY26DgoC4dM5L
2vAiletpkhOIOuz1DhJvPpk4anvlFazo9sQyT81L2funeGPBAKImGJc+XEEWfhYz
V7pbhEA+cG2Z03sJb8JXyku6R6pmIrHFuZLVDTHE9zD7T5Bi0dp9x45Dy/bUTMlw
nb9gJL9YUcYoEV4Kn2E79VtvaTSvRfhhIHvW7bjWqAnE1WoQpxIbxHz+HvQV+wvt
tAIjte2VVo+gWyKGmSMqZIewcLxuj5E53Xo1BJHWFUmge54DiHPKokKWKbJ6QVBG
EPQSnCYhBWeSWDeHH2n5yyXlSLXXYBtyHfbMZ53Ei6TD+pfbHWs6BlaozXeKnmcd
BEm02c6JdwDOtxB2nt8e7VTRzZ+boAS6PnHjIPCxW1WvulMLffggC0X19jZyS1TE
OFL0MCO6/QwUISgoIcm9r3MPHQk52n+49t9BgeA27M8nflDHgqGdXyWvwLPnv9Tr
C/9PK3FLZEiWEnkVZWMAc4aHalcaEk3viicRP9JaVVZ4GxZ0wLw8lmVdKEL5KLXN
zPzXJ6VfSGU+BCoNtME5Bv2Ic19Cq5twwGEGTwW926bK8RL76Fdgk6l8iyEX9ovw
1Ci8W5QNKcjqX9nu2kkfZmSo7h7GHMblqelLOvo8YBTA4NrU7lsIFUbxtbhgQqJV
zNSWlHiqbc5kueM6parww0qNyBiBZHzTIKYnOhRVh0Fk0tmhL2yKbo7iLGz/ICWL
wUhgLFeMlEKvqEIMZGAQvTItisz8CjxIYyrOQasZIDcDFtbs39LJ/rkUNXKBbqK4
cIjFCcwbtacjoHdbttM/1JQC65w1pOZSl76FfoNgZlJhq0l5LY/sIt3EFpC0Z4Zx
ICNqY1ePFlelcL/NhtxyV03u66abpakuk6HKRTZcBFKSsE/v9DLjRyXe48SR7PGn
2SwQ9ZfIGua7HD1kZ8RvoEz+zpDh41iI9dAecskc1GoCk59wXf0p02Q7xN1EHKTa
xej/S/qwqvjoz3GRZ46NfXDpgvM3Qw1BrL05BG/ZMNSN+1zITaTrsd7e0iSLbxqi
Myf1XsF+fArIpaXE0UzZiPoh4GHvVoQBoLgWOJg6A61KjG25/r+e5TWjcWWoFh/O
0j/w8gE74pHyK+HBoAMefT7Sap5FzpIt2Dx1Vsfm4KU21AerYsUc+X4Y+ja/65Ss
VFAbCNOefKFQO/c6Ko+KLhd+W+Qwlv2w/AILFRxfbMhgMQwnvumXoFqzz9Lsmeht
Q9ofbIxd7awufLGVVr7cQIzGW9URlqXpf2fKqAi6GNTZWD0KJGAcK4NOUyVL2RWc
I9lsJzfUhPbeQwscegwUBmm3xka/uHzJeBQb32HRZR49QlFiiHrLCkFIFlX76DQm
Hbq1Mj549nGi2VgQoLMbqpNLb5SuxVZyMKy4X2oIS0oZl8dIoRWP+DKnrMa5EwIX
9gaO+GhBzj+mURrTISQlCSc05C6sIXXd1x5Xw4fJhl1dqP9lEknkxukqIf0k8QYV
hJjSlWk7mn/5RQxSpSQG9dUoKV6Nua/GsTIh3kmnvom6l9FhgZjeHGnD7sTiXUnc
+v0ITI8p+XW0zzA9rN9slKpyPoDpZIwN1M52hAh+9DXhUIDqH8IVzr8S+6i4yU2V
e1kaMSlw0MA/lCEd6k8lKt7EuZsFit2OBQq0B43z1fmQtAmfKjp9TtZTAnPCVxqm
ZJp8TIEGNvh7XfvuoXuzlX8XpRA0c12T1xoVBMBB0R6LC/dD8cKWG+UAhTlsJL1J
89UfQRbiVP+AfitNrNKapgFYfRgrOOp2ZRPJYWjUPtMbshx64f+zoBMwqxxIXw9c
tDAfr5oGbK4Fg8EZLlAj0nzgAox4HtdOv1UfZYGR1Ht/voKRM29+ZcjiIBvWlYAB
e9YbXvyQUGQBfbbkFH2uBsEvFC5SD8MXJkOI0UcGF8n5zQOEd1f5JasQVvbOyB7E
WAMc2RFnTY5J0MSChrAdQiVj6SQV49G5aLWMfEjhC1iSlijKcifUkAO4KPeqm1Yf
M435mMIHHuAhufWtiTeZ5celhakg3SyETNmAi0Y6k12WF32TKMQZd9o4BtkiZRBl
Kke1BV0nSzrXbxQV5J8tsZY2a5wiCCO0lkY9taumEmpH634rXyT+sbkv/K+q3/p0
uHegIwKZDjGUl6f+ZGP5IAoEixT+rpTPXs+da3Z0MsXoPEgH6uClPROeahnqi/C1
JQeD2tX0Mpb7gjPGZJ5SWHxjjesFIvYd4/jEzQsV4Gx75aucSHyU2cdUlnKJintC
Ytsi7cvBm0qJ9/4qL4uBQFu3nn5+a48OJCRvwBy3jxaz3QF6cxQBUwTGK6TrvvDP
7L5ywUlH5OqOWzD/8bjQVJ11K/iGOPPdhGxUH9yBsmEOgR2MWoI7PbvdSJROtyRS
OxgkDaugfdiO2EepTfh+Hkra6KFGd2ZGlnRlnfzxnZlWDH1jNLjIHOiX00Y8U05x
ZaKIaFOf/7ACwodjI+Cl+VLEh8ZS/5Aa5sQuItGUE7FFSYTORJAZIIPQ7BCjudir
6DBt6t7KxiAiV7ZrckKK0Ca3lJXJ3y21532fHAOjVCea6fVTyoNUg7U9qBFnVnrb
Tv3TJPhXIr8y15RYJ3RGU/86NxOpVK8y4orOoM0FtJymg7qPoE3vWAKIw0nWlexJ
4a/ckTVqartpbh/LcQYzJiCz/6G90w4XkjPajqKpg79FyXj8OkYGGLylIN3CiqqJ
Ihtwve7Gibsjp5yGjpfHJhSwxfxtDXiy4MqSnk+wSGrIrVty889ojz6DSwM6AFs5
B/WfG9VIohlPwrYD17zTSX/rzZKd30zaKrIFZ1fLs6mqa+wG3vRoic1ukr/gRuL8
/0whhuOwJrValqPumSAYluO2FP8Ue9KP93dUoB+T52lHD8uoba61dxJzbjQqOJDO
Rer/01imZZrkFaMtesVX6oH39cRttXbwXdH44wo3Y72HKgLw2ZRL7jnlF25CPyBc
AEx2iRxPTjGv0Fp/M0tKN14lTTVtbzVBd/I/SWDntVolGUi2ZHfuWhpVYfkm256k
OdBESOWaMW296IO+1/sYj7I40QydFEOcSb3C45GlCVNHh6Xvd2rIbF51X1WTdIiY
aAnUQXnj+gPKVITimrOykvXBwL+fhN0YpDMx6v1CuFy0v5ftm6Oz7tPH04z6GXta
1+3AAwIJVjZWxlLMmSY9bkcwl8rUDS/CfEFbAPbDgEbRux0NPLBxcF6ind5G3fMJ
ADAE7ssoqM65slT23y6aPaagoNZSUB39wAf9JlBcLyQLfuQFTvx3VfMeo9yWtyYP
+vdB+dK3DaLjOB7mn03sYkZb0FLJl4cDrDuoDbU/+RE43oBDc1NEYoKUuIt285b8
1NN6HeazGPxfhvvWrZ+GhGUB8TaCyRg8+O19/jeBJLL5H/JO5U6fh8sicXCBM27Y
QMJrBEGqVXgFrmqXiMNlRluHR6KnTuNHnoVO4PXdpAbFBhtm6bg7M3zsjV7D4Qfd
m/4WJQUQQRbT5BIeR4lyRRnAv2GQzuALLwbyrVn6Wec/bPv6xPQSyd0nSBWXN2cj
bTqWaG8LgdIMS1MfvTRrgrXVqVaUiPrNLvrDxT5dz3zribhbW5iBGty34Tnfn14n
axHOHp2PHz0p86AD1XDw5ZTWKk9utsHR8Dcz3IqXOxNDYnTBmKPBmHQPVDgxSPVG
J8XzHvEASrsqPyAtBx86My7p6vzir90IDD4KyiHztfz61/m87JyT8Ve46iwnAOV6
zwFMFIRVwPc2JHYOc7Q3P2MXM1AblXOwyHoEnzT32rPBYogYSGeu5GMF6KybQGtW
hoEvaIVowRM8O2jbfl+FcEUJqPyKsMCGfTNK5m4v41i9bVDDmEc1eg0JgZiirLBz
hf9fB3PgNmFiQMYXOadcyBLaQ1e4agcQr2XHE9szngkaJjB1SYf4J22B/DNxy7xJ
CMDHY/J6LPE30jmDFDOj/7vFBXdU95/UxFgh5OiWBGhIcR5zkDKJwJHaQDTxFquq
b1wrRYkBtDfq6+k3Ph85qeI/nqj2eEZfiX92UGIgnsVPjA6yn0S2Dbt4UqXXEclE
TkwiFdDrlLGsAYHivNoVjWmuPHMz9HXxC/zh+wyW9UsPVErv+FcbobLMm89eKp59
ZFiPnGSFhBrdB1it5743ob5bCXImqiw6/o7UscL7gaknqOOuWGm6TACxN2P61zJ1
r90TgTvW2cn96gM7+VAS/kVq32PbxfVrbCByTkKu7FruqAXbikOWjy4GqcP03pWD
5yW3ocDS301OaLooedBL/NoCoMUPgKpb2YWfc5morP6QUEnyZOhZCpCAzauvzsgD
/rMJNcV2X1eyq9RpODuaoC75UKy4qxpVUIXIDWKLcSdBoWlX6mto2jkxiFKToggr
C8+5Y1TBHL4tJiuYhBdLj0pxdhKfrqhj+P3Cd9pqa6x0a8tBGxh/Mw9DFN+iDmPy
n02/yQM/YEiSdJ0CI43IDK83o2OprepjBBAJW8J5UBzhWA/EPB+cgBNql6Z6YiBt
GzX4v6/86BhQE3M2Kytcc0sxIAFeDI8Ysj2OlzpBEuGf4lFnMdmAsvgUzX0YmdG7
nANvfT5N23Ijen/B5osj310VDVbvvFZ1lxbCEy6Tj4dtf6BBkz5/6IrskgbRj1Gj
oZX9hYmEILyYlqNGaZ9815XV7j+pAcVYnnJ1Axlp3Ox8U+iI5eV3BVXJlWagocOn
vTOE+S8zLpo3PmrLvLQucHxuduZjgZ4Sd7h2nXB4QCY3AQrsSf6sJJCnxR8jn2ul
wSO1EK76oN1n/m2BfgMlyVyeD1BD2D81QJXuZRPF/rwVkbrlxbVfa3PoXPsEde2b
2CbNbF2n4ewsJdHX8mgyYbxlPzW3fD4ZksnRSm6xh8NK8NoH+uRJG3iLjTDOx5X5
KodIcC6/bvVLCHa6Q2JS8vvrV7T6aOJVCDxgYLJCDlwNM2S/pxM5HzpcKg5dUDOW
LZPTqRWiSPho1fbu040O0uIFOxc3X2Lyc9ev84yg3lFMxAg2Ta7zCAIQ0wxabQIR
HWWqBscE+jU7eXpgM2LYDCQ3AIc04Kquo/SaB8M7OvT2t0wpMTUclHHFGUfgV7eZ
2rko6bz2qT2MCgOabOSVM6ECBM3mlX5/IP8DiOC9VYoOctET8EmG07BTu1IN2xez
eUwhl+NWw1ZOwGv49hk162pRn3rKC8O0avUhZpj7XSmNUmmLFguq8Tm7+II2yp+8
y++P3byUbj9iYfEqJH47pXNuJ6NM7RlmVqgqxNRQhtDFMB5tsz2nf/RJ1qAjx8wr
zJMbAZJQAWGhf4Uad16hBOOg3Z9sVOz/p7Zx5hO/xmThXKj0UbHLK8EWxK6ZPUot
mxzSdTT7FZ/6nxDecHpnEZ3PnAtGzow8eylTx6L1BNqHNKPzu0Lf8eAHwwOhKGTJ
uaMdY+bZ74LD+6xlj9RZbJqamZamUhe1lIdi5IiQTWl+Pt0QK4SJ3qgZilr9+B4U
37euVQhsjU8KieLx5CCkuOnTZY3LE9nTFki5RI0bhACKHZHpvD1f5Dr0dmFBj3Ja
XInzcZYU0xXQVCSxPe+dPTQM8TyEZ5CpTfIMAp19pRtSgzzLlDas1F0ej+gpNN3h
ynv2tK76vJblBo6oLWZCOKTp5W7OZehRcEdICVu18XJj77zolXGpzxZoURxrALKG
c7M1hOgWgLmAIterwx3ia0ijbZDk90+MFbjO62Faviuuno0ln3JrtyQXxknXS2vb
B7LL0kLldyCmwPB72BIVNkNVDlolKO4TmmqnuYvjPIUhvkkuus9bvXKAKsPNRUVw
kh4u7iPO+KYOhN2psHXSGHVo9Xk867vNodRFQqAbHCJavGfZVd5x6SnYrS9TiNd2
wrSPndJ+2Try+wGTO69+cLDRyvZvNGyUFmz5pJVjmn+SAjuT9rDkaWI8nKtB5kVS
nGavm4PSS6q0GdElEtMWY9RUGDiV2ffIqpASEi42B95FQXz6VuO2Ejryt6K6vZr4
1QeG3wNsvuO/QCH+44B9H27lcwimrly5xWVPUnSRz1K6UoYvI4h+vref6OvCK3QH
BCTfFcaveHWJ2HOMv1GKO7LjoHwlRJMgLjG1kQ4inOii3AeK9BTIZqclMT5eMLw3
ets2IJVbeZTm/QhMszpcWB56j0zRwuT/dW6JECLx4Xwi5wegjeY31+jac2Y8mczL
kZjADDNo4ZhzmJCmfxfc1MmKQcxbuOk1sgBLlZi+GcKJ0Js59WdYqdNnyRwmTZCb
On0FUA/9t3mO3GL/TIOzPXS5Snu+0SJc7QfDNMKHc+kCBbJqHnDHAuKhJYt6+4pB
nWmz+87ZuTa1nE5FX9cKh29xErLzA68paI1782Xojn8gMtU9s7InqA4nqLCrpj5B
qJZU6TM15cXoiqKMboSbtRVd6PABjEBd7fnZXlMktTQXjbHiPOw97gUqIR92ynDM
x8HVNAmWcX34pf6sMm1t4lBYq6a/V99pDWOwgt3NoOPLwNHOCFz0ULby322p9dCx
PlWhv63UNjgpDIWUoGCB2MHgee+p997MJqXCbUO+Jaf1xYTz6Bxi9wNQczYHspRu
gtQmLxIdVkHpo/XVpNSrzz+EMS5OtF0lMHdjFoy+yEo+iZj1iHN/HUnMPGsc42mJ
WowsqGf8L2ByLYOGOFCDpxZPfYtE/fXlXa9ddzkJAe5frL5OfJk9WX9Mr0+c5HQe
O1MhvQzcj31GHeD012/Njur8PdoV1OlVRIq2y1iiVy8psFFflOeOxSbkQP/Cxvvp
zwsHOxDaTWm9jw9Xvh3mVDImaeDQ/BNQ0M6H8L69aTtE2ovDRkN7Votoe9TZGvj1
SfcmUteNWvtwsgk/YXeid+V9TFySKH0UOiW4MWRE8/huP20PkNJr5fC93jEqMmWT
eoIWK0jbTnxB5tlYMRbpDIf+fnk/qC+Uigzj+roys33nTnf7jMcNPh6dMlPBgGl/
AmdnPj2i37yH1xNAs2OVjbb/tK/vSMGT2/u/8BT2xelFRdzrtmivPgu6uQbXP1Fn
PWe5RvJmq4LtZD3NjrMui2J55BR8oZnO1VO01KzHme5oD7FXu6Q0xMnPCBas0f7u
C58AEUkHTipo1hKYbRHedN3sG9dp5qXw8AAyLBL/K7KbIXGqyjRQArflomzJWI4l
xxJ5nv8qRuG9Wv2RFXGEyS6R1XQ/ABH4Jm8/625Oj+/vyKk+AhKTGgZ6BW4aiT+n
515VP9FnIIziITMCEm1SKR3KuT8ba+XBijWUetFZsILNru960mmtr7UO8obLioPi
BkCeQeDl3E42muzwIhtm8PAImkaGGKDrKMKN68Y8n3fMrSdM+FcDvCymanVuskhJ
PEkqIsKuPLjIFplKJL31UJYjls9eD+l0M4CbszWyDGJIOi50tAcgTr2mRW/oSiGG
W0Z2USHgmQDqXeOFuAU/1K9Yt07IBVvVROvGwbEAGd3MZ5EM+sIIfa3L4OrbJ7lD
U1IaOOd27bBng28aRRx7D63sBtBt9+tjTPc8M9yHxp16eAzAsslspoD+oBG3Lpyi
J1wxS24mByamAqcp/9kxDNx4VMEc04FIeSmJOJ4mJCR9I7tMOGixA/wNt6ebP1Il
pnoUaDtl/oL+FhBYOllsjSSdT/tZIP0eNJtyXatmuGEOeVQuoX/0vQBnG+lnmSQD
tk+8G0HgYiHhH6QvUQDRLG4Pf8jcbu6QFI1kKEhufBf4Rf3ud7GdREk8txb2ndms
ObCDctAdnzJuIIVm6z6Ajp03d9bdwct9t4/tzJrMf5dVmk2TBgANhE/Gscc5Pejc
xffUCuTohwaEYBNXVyWJr2DYvlEOkEPInUTR873EgzSRnhEsCRQCq6mvW0pLjoJG
x1j6iX5V58vcw0Z+vYEz7cgvJ0u/eMpWbmbegdIWnnUzxes2rK48PJcipUuOdZns
WBMZSEyMh5waFUn2nFdoNUnjYOI3ONvjetTdGNcLzNZfZMDKxJxTM1/tgWNcUjtJ
xw4Wg7qfj022RUs/H5QO810EH3ho/CwSnFXxK9vmQTj59TyRyWWpZY6qa4Qa0jwb
WNpXb1w0iwdwTJpSTVDqc63mt0PSnX/Dqz5PG7UAnMPo5d00FFrp1QzYEKuWpkxB
7oGhiFFFSUheP9+4OyMS4QrqcZAkVvproIPlo9VK1ixeNbGc9X9fklS8g1YeKL1A
ZBuq8UO3gJ6l3OIb5qsFNgkYDzBTGZU9ew9A5f6s8jf5e4j4RO6dMheizaLCyGxI
Notw285qGjuzQ/Ymexpc/vObuYXdQs7P3abZuY+zfVdv1iD0oX05oA5eYRP27hMS
xL6FNd7yYLV8D9FehflOIupQdwDyYsNYfr9eM4SZSVfFEzY9JDKpS8a3m7xtrvri
wCwU+zIi6h4eQuSzAKVd4Iozsf0OotIxst4FAZDb8Sxs8cFZNIp9LLxsvB4ageXZ
jsUiBo4YFzS8ztAwoqdooy9C6L6+yV9z5Ly7vKZ0EwykgzJR0Mrr+I9zCJVtQS12
5VcyFENsYCGLFFiN9f3tfBEz9y5rrZQlJH1pc1B30bglhftoLlR6uKf7XC49FUp/
8p1roD6h1CRZyvWGbjJqgxolzKRXGgC7CEXT7A4gsXD5dWfUlItJg79QEhRtKnP7
KiajnJdm5p3mI/sbvEox+twvx4KxZCepwokt1vZNrYz+EtPlPBGSdorNUHjAf+tk
e3AHBV71Pi34l7eKHTIH6QqMNCOlAv7hjTCReQxUQHqfOh7a7IfiV7shmH/n52u3
N7l+8uj9sw8xY4yaEKbNBu2ST2ocT0bGml4BhAqQRzUAxnY2Z9Z41oh7+flBcP0b
b3Wz+gY1qROyofbf7YUwHTWLeeH2zVanMdpcHdyx2j6T49d+VHAXb3mmua8U0OF3
/Yr5bb7B1ERRT3c3IkvyBC3PQaqcHwKL4wyE2MhaPal2BsdM7n9foFUac7CAEycg
teicZkMLXeVI6TzqOZbuHz+YWteu1Y28hiAsQIw8AE7WNdUm7hly6Q3iCbCtf63l
LWyItWUIu3WXyjZjmx+uPdkJdKhgbtgFpqKyKBO2toFqYgEHSvtwH4PpQEZPIpSO
60BUq72bOv2N2FTtAv8p4zNCeRR6cpSikrg/xHAyER5T/a6shVsGFKhebbGWzZii
`protect END_PROTECTED
