`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Er6G3R/VwFK4YZzBkWyFdx3wEgEqmxuITAT9O8QXRj3y0KcEF1vNWfT5x06XTKcl
uSSfYXpjE4VfoKH1opNmVindzS8/Esfx4BPGrE4KvTPaqu65H0Rd+HHhlHEBXtdY
GqBTni3xQUnjuW4AzTjuiaGQ1UsZqHI92zU8ISUw/ZaALHc/rTf0u6gkvqsqORWb
B34lpb33H3xxnTUelzdSDIIPyR3WTSKv6PyHbn7d4MhHW38DKRoI+L0AytDBz9EE
vb3+pebeV0V7Etb5MvvfEAJ8WgFSnD+AmLY92R+7sdVGFNdmhsZRMOhmObmKk0/I
2GQ9C343rLaj40CcHrwJXICxOfbiNIl3Y9P20z/tSKIIsQVyh6sigtUmX2sDJ05K
3ih22AsV1Sq9gmRkktYbSd4kzeNCx8/k0dQEIGrJ3RUf2rgOd89ZveW83iz8JuW6
d/ASu/pg8mACu4FX27K2n5vMAaarH3hyFhIU0PFDVfOK6u15uBDyl05kUMrdMYJX
9KPPIrhOg0fj7Y1dzLiH+eEcl6DIgJJRVCPKxFhbeSJsfdIAF6BKWgBBbvy+zlcF
JKYKiAqKggW2Df7XCc+ItWJaLAoiGz8z1V5FkzahZ9Jjl+djqtJ+mHPCN1oH5cQ9
5v0ZLqd28bYyaQqCuIgffTEhR9FFoqYarHyM4rwmE0ZC/caCwp+MS81m5EYqIioh
lRLheg13p+BGsekZWRZfax0h4lHe4FmJCV4yuD5PJkPPdWCaYEI75nsTgk0xWJcO
0/9W4L9UtlSYNuP6xB0YReskfDXw9IXTI29FkypGW2KI4900TPhmu8fdY6GDXA3u
vPM6/aqyPJgEu1Gbhz766oak/Vehh/M+IB9NLtdZJek=
`protect END_PROTECTED
