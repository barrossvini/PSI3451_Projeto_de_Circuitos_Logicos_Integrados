`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9xWD0muo7Baw1Krb0kAf+lncN13k5zU3PtONALb/9VtsRRCIEiBPd2PGfTv9sAxg
gWR8B24TWm55+G+Yf1Kv43L/h+yqcLsINywEEGwA0H+Bo3oyJm2DIZSbdnwrzXD/
okjQvE360lUHKFPmwjfkXePrXPJIC1XY+DvBYQISLODlzIqL+5NheYoLf45QotLu
WOKifVRb10Fe8ayj2QCxDYl/gVfrces5lOrCKF/xf4N9qSuOHyGo7Dg54t13fSGL
sXu+hkMTnDHAvIDvGBFqvhNmPR6m1mQqeLO7+CSUyT2QSB0N4aAupSmHSiycYTf2
7GIKPG3BU90giUxyB0AqYLxDh8VuEyoIK5lSlfM86rWKPfap7eInScom4aN+wEXU
6W7X/2/3cGpLyoUCq3gIomB0wUWo4Ql55yVy7EALVxpcpQV+0FXtKYlXjckG2TDI
`protect END_PROTECTED
