`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g39rPLlLs0xMZGIG+HNHQRPNMTzXyrjFfMyqv8U6iZYvjwrmP4RthiInmiYaiXCR
61HOkAwWREdpnqsDHp8JUuBaEPj+G/69kkqCySXiwskhd3VeWfY0aCCYcpClymbu
4wingfl8Ha6qKamorLEU3zSHG3gqNaBSJ8XZ50W9DiVhW7x8lYeU/ktdvXQeXwno
qKwWkgES6HGvKN2Erin8WfFQ98Wr6vAsiDr+tn9Ng77cgxtQEXBoKfuqsxAxa0EC
GDYau1K1ccnr2wWkbL0ilkmQuV/3tOiBrCuhkK8AA8/odEdUWmOWxX8rhgueobR8
aHu5tCic1ib7+OyvXKvWCR+2lUklN90XHxLNLyrUEtCrnELj2LUQDlnWSfFKDkkQ
Jd81/2WX/n67o9Zdy2C4XyXMTwXoW/Vx0a7Ajq6vYC07xslDouqF3aT6nnGFfwN4
S0+ZAOEP3wNdwyEETfCDRLnaG3iJo8Mhes+BPtclXcYrYNdM+uyUN1JZ91UXlYh7
Ub4I+NBFVQOhFXWkkEhKyYWstLcJhhpJu3WByogGUaNWV/1vrEo8E/Wtq4j7QTde
WzHQN/Cwi7UHEvjaGClaK2GpJj6LlWqqTt41/TLA2okx/XSk+W61I79Uh70/cC18
z4AKMnTTKPTyRf/anz0zqY0KbbLG+Ch1c15NI0HMwb9FHENvzNmH1Tk/CQxnQu0Z
Ojy/sU1/HQWAD7N+8RKmUequqRt+B9U0qFT2XFg/2nNhgZQabuQSjC25/bp4vmvW
V54+89g3It4ZBBnm4s2COaf7v1Noxj2H/dcP68lGonngbSQnzaI8u1ea29ipAY45
IXiTWQzdFvxlV63WWDQhaDDhWdWiEN3pTEhYNsm0Bg/WYXy/jx2gK1S61swd36yC
Jz8GKiNvP0pn3QvLVilmJKNI+DDB3Fijba4KLqqdhDpt/UZPDYlX2Sa2bF1UKPLD
12Hy0ckyTCltI53bruHVbC28x7ZnWUg0oM7UeBEgCkgu9Zjq+n/UFYE10JeAut3R
hejxDyXOcAqiNSUc7vttjOamAqcgaw3/OW0DYA1zVwizD6Gb0XAQhOMTkxXdIf0v
K2dzM8RZm9SiCkZzC/wz93Zb0Fv3DUT9cyelU7MpWu+nK+flB0iLbmAhza9dhRsW
ExcHZ4AXNh/OadnG3PMMM5EWlI26wm/cWqh1TpabAbnWPXyOEuu+3N41xJnZ4p1R
qW+Tjhv3JJJsOBI3cz+dFGZIhDMPz/dlIR1pRhVJzAtbksemHuLSUvpE/efEs6JS
KWOB2ai7aIH0385IlVIVi69q705J9Aom6JTMhxQbDIIUBNoziuSe8BYzp6h3CSit
y6HJLkVH6kePbbR3UyMzX7M+NXYR3Pj+2PfXov/UIVuH/KMv1K2UgXXv1DTBL+hQ
I1ivdDSuiPipaIgmNRAXTAaGrVfhcHS7OtKYu5WIL8Ixkj+3B6QkBPPS5+rsoaIV
uoXp7HC+nzKPqFHyhdDITe0Ix59iHLZEAd7oMdJ2UgtQgraj41v4WQRyBxtgWUiC
/J30S/uIQH5VhMIeiYeYARJaMPHNLfoZ1vL81RpNrHtpF+U2eMX6ub5Q9hWuZ8vX
KdAM8Cs7MouDxt4Fq0adtdSBDU4vBLT/y7YpJmGmBYM78TYHmjKaN1mE8YSngbYg
zyevGCbzcZgMpfgwxWck0YAdQ+hPknk/E++YPhsUQzSZnHhgNRSk3mHRuIZatgHi
HTNoASQWXVoMb1NFbl607bi4tBUCREfbWrnbL9RIBbPesoMhASl3AbfxwQhgtWox
ywz7saqp/PYiE1XERfJ7PyjpGObuwxexeXOU/gM1WD/5WjaaQfmQUeWM5IReox4M
e8An6Ct+6pCY2xGWBELicYcKK+grTyqvjrdBQPcOhK2ACckx4z++bbBBQCI+wfn8
L92D0TySf08xdBlkxRLWaghA+LKY2dWa3rK9dBZtLmA4iScaKxc9IxScTSCupS49
z9H/u+nRsuZJV1Nupz6j4zfo678V70bl5XZRhgUDn5wuht99J2QHyREJNUC42l+4
NIwHunVnkyUMRro56NLJRQS6byQ0n6xIUJ5vejwhoit1DK/H4o7pOEyzmvRLg+3c
UdVIR6wBBryIX7JlQu1ApfhtlERfDLfMbv4x+XUTfv4mqNmYoIy0DRNbGxSGN9wh
J6OH8o+i9Ys5Cfis9iirMQufG2AVgt9GLGpOC6gz4cJ/Lx1Kt8iFCedgU/+BnbOI
LQL/wEeUHnx2nIg2LVHw1JLQTkQfTxsSfg+BoT6XMVRfhPYNjDHcB8ECpf6wK1rk
rm9aU9ebELwK5qoed1R2202y1/+pdVnm36YZx4F+5l0sh6fJXRXLncgmAEG3Op7X
Exoq3nZPdS6o+DXxB++FYtPgRlZSLuciUfira2NK2OmTkJlsSps9igGUPkzHadOg
AywWjmszcnWwzw7OEIHqnlXdgMehkvp6TvezlIFDK4h8yYKFZ0mnPxfgKsk1JQVM
gJds78x9JjtQeOXOHTRU1lpJCG4bMoP4oZwo3Hdtp/fDSaxY2NWQm3s83T2FX0SI
Frxvm0XqKSHpP0Suc6VAcHDEpn0k0SvUMb24EkwAwEgxnC+Dc5yo94g8UiMfBVNH
TG1bDYzL++Bc1wlhj7K3mW2UarOZ9bOAn9YOK8g2yJML33fLB1k7/1o/47z5zLr2
Y1Mv3d0kY/Er87UqtEFJRqtXuROrTCcRqCLWAemt7LEQhin1WsRfnbsVz5c3deyP
Q+tT5OUjlOBdwZaDufbdjhsdG3HMRvxtQRhLcKwFZwxs64zM9IZ10yREov2FHnYw
4VVGUr3YRiR0jLScp7AGg8XOk6uoTFTVz9uglE0tOqU4sBtL6/LN5lrnit9g6ye5
JeM1T2dZdo1w9Nu2QSNOAd42jQXQoLEq7pMHmtes6M7U55O24BGizuLICWo+qWtN
NPqU7WOurpmeDxJ69DkFApM++WjQOcVIOHLT3Y1ra5yARB85YDJplZkq1xOUvyUj
epeKaxY2vHPX32Z4QtJvN76t1a5HQHHmlvt9LsE/z/q5ciYMVeKpz5zNeBzqhdCc
IO3mM4Wz+NJHuvkYUZQVoq/zQDGnSFVj5R2h8J0a8ZM1KXUSkQusqhR0F8Lmhq+d
IbZwgPHir7nawJXDdKBtcTgQ+muGQgaplGLl0tT1AcWoM4fGH7LkKqQiKwQuzG1o
fVm6Q7wffTPAjr9PFunJVvD+dlCzWGvQn2WMl1i3KEyJ+KcDveNGbYtoenVKVyBp
BXX93/jSWHe/T/5R+Tc8pxpvwB80bz6Tvq5brmLZ5NJLO8843tOgYl98CRgWgEvY
QqRDXjR6dgk+uchfVjbohJeQTZFP8KLwZK9Y1/loI/uDyLqhJmmYxCYU53yp13ai
ZQ+kA7hyh8Jn79PldHyAmFoAQF46wlXvlfTy9sX+uIYULJiVmgMzLtDRu10evOo/
NDeiJXJpDR5dufQxtppiPCBG98G7fbLugrm48ic1oFyCOKwkRhxgLf9dQpxxivGy
GbT8aEnowjdTplEmp8G45aow4VQmwDldCONGTZ9s2u1RACRpBVTmh4AQBT5EnTiZ
Br9mxe9vs2WgijhsmgT+r4GMrYRFsulCcBSBefvduBobBwrmTvqWRZ/4VhFQKsjO
yUVrtiHF7tMWi01EqZCin+CYwj8IuITurLgK2ef/3eKlVNredtC6XhqAY/tYQ/zY
YlgHrHPn11ph6TVfvNXX5zZJiDMGSF35/RULRaUXajh70PB2xwhNpWG8h1QnrdUm
C8HVouZNIt06tNLW+EK1kzyL9o/H4QGcPoSyZkqRyeSGNX+/h/kz1KYY66Dq7mg0
aMKrt5ZuppUniPS0AGZdMRdvqyPV2xl/5PsQXNlyLv/LpaV5vgE/wwFf5AJmappn
KN5s+gQoRD23yoKknWVXC2Rg59Fi2Bi0/16PGB/w9OCV5Z4N1maXO1DDyUkL9Pjr
/q71JkbNwVeIxbqLpAHHJH4M66m23CIlqnSlanbY3RB37XoI758nvMqWQPHJMftW
HkP5oitXRw3atjvykg/ZaKbPn4GbeiMnn32IEwom2yZZkLRxfHMHKPigfoGzSN2H
d+SHejA2iFYBGAL7YMuOcKChL4Sg2QExytgjqdrEBGhk2RKMTmjBQceyRj9Gv6F5
EY5do/MGH+yrRGQn2htAVGy+UNl/CHo4w+1mLnavoQmNKl60HgH55tY5KFUUPHfe
7sIydkAYBSKCvNF7Q0ei0cfvt9trFWPJj30zzYqfiBIYx284XQO92Zkds10JG2Pn
D1iVSiJUPGUZBh61XAEK8cpbDaGB5FtHybLHWef6F5sYJvgjKQ7rqqfdL5LD9QgN
Rx2jexAswbchFIW99WZrt5JCat4ntTFcCd1HO6o56rdE18JUYozl61uhXpx1mxuz
3HgawDgk93R4fHrfdf14Q2im/qvxTttIa/RviP5CqvODGUN4bU7v1ny/eK1Gvpda
s9YVTGWXrbiJ1b9sAptHVxCJFJTv8Z7FgQDCBWUbFDPt7jNjUKyvoS1/uOii9SpY
XW8BgkMtIoKG4H8xIpJgr+wEqdcCMkyaVIQ1tSC3QSVfQcLUJOGZLIM7Vmrxl3yG
ydxwJ/Rb32MLCIfdfMW8fSHOaBd/B95C+/WEBqIQC2VVlqmXeOkLyQaBs/rs8DqN
lG7jaDNvRm5E4cLesFV01dGKacqq7RJEoTh/s/BtxSGtA/uXBvMmKZHLwD9NAa/v
bbfCfzZzSzxVI/nGyXEHGQNnbgTdb+OJtbQScfbHjE2x6UPMeUL24oXdW/DCV0R7
lDd0K7PBTfBFQgekx9c0y9d5wSy9p9BFXBB27HgfDKXmyvllHkrfHamod2nqmMnY
D8NvDBWbo12ybUyykvVzox0vS88HQcASJgjSt7uvoDsvYsGM00Y822txxfmHnulz
Qz7a4+JfOij0HORaD5WI5fneLX7xl4YQkFt5kqJZ6dg=
`protect END_PROTECTED
