`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VfE96v7Y+qHT1Ds+bAp4zu7SsDGNp8dYKXiL/rNp/c2NcPCuoLl0ueyRUyln+/fh
NbyT37uNEg+KlP91KJSTLC71FEpZFnJnYCeR8To1rxtsONUAUc8amTgx+34rn5OY
hTJW0CLXk37rZSog6nSNcPoEfSExccD1KrJghn/w8PpnWlqS61nyoFgXvMUKXOpQ
KshZ3HqjJ0SsNdM+6hRDZzBgpMOll1MX6iyClZnyya6C5mZX8HThL+Wouxxo7E7w
KzJyYfZwFq4kN3rFSWCd7DSsetT80tgDNN4ZMX4RpeXEUciQDo+oETn8MnxXRmfE
c7HiGW/gLoS8DBcBnIABoTFVTGu3/HiN/K1Dffc7iFlkTyVk7o6ZkCVgJ+hPK6+y
1elp9HD0dQMQL78YgDSQIp49x8GoFIWoGjJvR92xTOuv9+BoI15WclR19RKySCIT
n7x353TsBLTNgAboK93okUUk+FRq5Wyly0fqkV3vwmeFjYvCB5ypwCuQobXQqHu2
p3lOJfAXwYWvoxo9DlmR+GFdwDKxHB+fNjfvlma8yAxZ56S1kjwCCOthKtsKVZpA
RJyGayO5UcO9lj2+cXKIRM80e3DfqgjQil3gDoCXNSbalFl8+CMFBS7flv7vma9s
Mu3anFp18y/0Hf3nqn1D9YZftUMbjUjLwQmTpe/joE0DYlGScFnMsSxCTDbpxNv/
76Gp5DutVItw15QOgREkgIKBaciFm50MQuJaNUDmCYhufNVqZQ3QBKed0F0VeppC
gsAhYr8jfCv70mM4+INxKZ06OUO1amMLwfqMidzSYaZUsENqjABGlJx0cWkrm5ga
gx0TcM5BzBHgMBMNwRpaZG4b3LZ7jwQjgZUmnUKH0BPEjV3T2GrjI5aP2Qp73iW4
8QUH7+jH71rEXVRh7U2g8awcZWtXOM6TEUPQo4B+dgTqZeUQg/sWgPAGUiN9yIsN
ufMxj26Pbl9D3yJjb1rgGiGs3+AHUDr0gADMC90CcfuMW+olzXyW3d8qbrhYvYlM
kxrLCFuzzIAMpcn03okvrDeH24rkM2ewiuSmBSKAN+0LGHxNDbSFv822ldiP6cvH
bN3QLRs6ymNXIfv7fQJFqMGM/L4zS4gDWEIpef3k32Tjpo6z5wx53T5sUrFyR+tp
0DIRJPjMSpscK6/Vp3rUKNNJ9WxMQ1zL/XbK2irIiUfNRMETuji6Y6k8U5CODJ8C
8QwuMwS4okPIv+J3VURsc9dJhJ8kNKpANfpSbUg3Uxa7UNg423SqGLloqEJJNLdJ
D+LYvnDWId/p3GXMBd+bHnkOaT4sa3jkwsM/FcYdgqq6Kw+6C+j0MhVhDfyygauj
iGUDT66emmfvYSLpoR8IRLTbydBnbkViCHTilDnD5GA2bIw2uoc3dep1pUfNqbef
sBTCBH6q6+X5C/3tY7DZ8ZuaM7mvVIZclnIca/KDtmTaHgiryW1vd8Vc6yihD2X6
0VCArZNps7pOHKPd6g7Re5PtXFAtFnHpk+U1heZLPCEMQKhcyNcECdBMUYNwOF6/
3lhjOGk0cieb3KRCjb/chV6cmoIjFPE4SaS0m/b6SttLgDDo0ojjx5+1FuK+DmSs
D5xqo3d3rG9+hAVztLoB/UenbOt09gQDNqfP/7m8m9/lbCpyzmbeyIZ2tF3qlpTK
/Vdxyw+F57FiNv+5eLusi7PQx5ViyMdGq9zMDpLC+cO4WJjRRkUs085x/5NKk0KY
BaCjSLg9aZBoGxO6t39dJ9G0Cx2le9KZ/Iieox/jodBsHbsXe7dWTkriH4cW+AmA
hlNevWols9jrP/5Lk2Ll41ztqN/gchP+eATM2OOLFqER9dbxH+AoRkS7k0aNKrAG
eRoaGAXmfeqX0GwT4sDkoK1GL8VjNbDrzzL4cU4kuSk/22DOdANTRYaXOhxzmjV4
H1eWu+s83pwHF8RkRpqf3tZyt3NSQXBT2MCCA4NB7mQJ9LPYvDNuwa/aXvoqSg8a
TvtTX+FNT6J6/V4ydtfP1PinFwWrs55bc95s8SjahvwpXN9gEyysl+odcSr91+A+
VgjYyndK/JWa6l0/FdU7oRYVzWENHwcrHve9NJUfBWi9OGFcvYSIy3UNaC/TLOTH
BJrNeJB9H5tEWE6c2sLMfzzcUXFHdmVdrvaG8PKKHXsR1KxzXPr+Px3bYtDVGvWH
ZKgRWoK8PzPnnCyv6oe25DYBnD4q4A4v56rYU5csS6EOWQLw+9IKOuro9HGUac6N
yw3qKJEgjej2l8JRvlwB3kXFt3++C7OTMwyWVRByCio2Yg1uNbf6/s8U06qGYBFe
vnpfLwM/8lXjcUh59EUjpVYLgNn5duUAO0mmpzg7TQaYYGYYhd+DvKEVzszVCDTP
ABzyCijRgjzwgFdfvufI2tGEfgBEA7AX0Y6HI2YKGLXKxaG6pnDAr2KFAtj4O03+
MZ76vL6uwaI6nDOYvNXZpp7jV6TfKzZPBRd4trvIL2/GW2v5gdI4pW50Ic2Y1zX6
QSYBO4v3suDDUiedMItY9TLm+CTIl6FCMiud2x1x+/MyXtT3ZrGoHrtT1rWoNw8G
f6qYBvtAYctFgF9TA/ZKNdT1nVC2JiwH0Vta64usM5RYIlzzDPphpJfniQ1iGyIj
6RYMbYtZA1U9xyzVcd2agGYLIA565o1xXmC8mTIzJn2M7TSapAvJ432xpWfQN2+S
+IH4s51f3/TAT49e8QAnBkm0BH81J/nU2zeZ8FCk7l6RnRMj1dLEliIUZLzDnZTl
ziwHJSlS4vWUYNIa0Cf8NPnaBxg/XdI140nVnh/IBqzbTO8dWsJ8MIe63IrqPZye
qN/FJ7XrKpXsskauQWscKh/Co/03YU9KZAH88b+Mb67Bi52f0pzhyLQBrvwCEJgt
EZRuG12+ap2LovmAClv1y+v2LFf6pN2kH+FVMJ/M4vxyClxhwsUzj+0pLK493MZu
YjCITcEcweO9Q/Pl4ux2nqF650NoFbx4tG6yD+eg60WcMcnZuuOzLSoLgRTiXq9p
30/MagUFfKPRB+43OybsM06GcMKEcBnjYW9g3K5VFcHMlhD3oUe+MvpmeZLJvgSg
2ZsEkNHuvHnfQh19DEa/BYnW8imOH1+deioF/M6BBISpZcmWgwXCeGzYM9LuidkW
cE8pmsjgtx4fywK8lhxKSkYCuk42vhXgxmufgZdJpIbNL/dnaYf+mrNjPBp/vMxr
3OcQhIcjMHPB+eJRc77isskyoF0pqHqlxTIK7HgwymE+qUrBdYD8Mc+ZdUZTREwP
VXZBWOVsZlNRq3sbQSqVFwBxjukOcMlNI8Nax0mCrtvTs9CdRxKfCXsnx1QG9NNw
fFE05FNxkMoOLLlfg3DxCnW30e2N9M8f50LCT7Knjzrtg1kA+TEyMPZUAXD5ZzHz
MSifn2TblXnRJGKwJUX/4WHshOpXsd5nsZzZdQXkvfY2IhKfXI/Xyvg7y/AASyXz
d2O0TCNY5maW2cNYJmnikAMqT3pCv1XBDbpOTwnIu+2cjWUvTmnyHIro2aUO1i5E
PhO1J4TwqsnGWwcZYetwV5QqAnROi0rFZxTK17Aevru/3TBTpsol365fSaBmMxB0
6h4GuIX9ijepJHwSVCMBox67snMgnnHJNWzaQmTjwnXgBQz/q2AvuRFo3ydwR+2R
ZT+dnOdqb2UfFKV6dniptj3OchUdZDwGvT57u58kONHEWkWpJaNGSDjDtpbZj63u
Ac9nosvTVRVhvAmtD0kKIB7tLRlhaMT6IKQVO+0Nz46neIKaJMm/EbJCjq+8FtKG
KzQltvWCQiYGgP8ohdDnJr4AtqG3Hj0e5V3ilqrGFM/R4NlKg7CEes+zMEqfpubB
syZjSpVvjnoM3OH1x4DHLxHaVTmNZuPZpzglr0VqX497uaQ3QhmTclXt+ITwhWxu
aCJFiSvhG7hopxGS0JCM5bkg6303MzXSIevdatcrciMzuZfUnRx2H6eMtSk5JkkD
UPyOEL/TkyfDTv7UOrwzjNoLu72dLAH+3tNhvCoNNmQ07Tpunc64iuuw1sFj5Omc
Bi62tcg49NkrF2EeIZ01/vrcRRhHkO0pahAafpJueRhnTyamvqs01TJlyPwEXpmn
kMFWOocFBDEqBBAtXUrTPwa7OCkTnOG1x/9G+o3MmTgaYPpbSr7Gwj1uOxs1kYGV
0ENGn+ptS0J2qeh623vbJD8S6mLI0Du6f1yv/CS3E2IyjXPOrQ7qsqo1E+1SR9FK
1CZigNX3kSB2dIekpQWjcTr0ECWUrGHhzWiSlegkGfi1Xo5zACkJx0LkLxnqUmL6
DGelD8D3zsciLsytaun1eAWyLDOaVGuoq7bR7dYF5IQ4Se3TSwrTo4kYwQBd+Crp
ShHLPaBsc88ZiwvSw8Pdulq7JaXTJIUEprlGacP1M8R6BLZy6CCQInImqQe6FZBV
l7YiMOBAS+CwAZO6V2KqqoCzwbfETLhfzLaj4UI/QSuVa9ZOx++75DLmxoUKsCaT
/32p2b3/b8A5xIWeZRK//qwNCAk58QyUSs+eV7+2rsfVCe5EWwEqi6qhQ/hrWoxh
7hxttPL4rtTWOXPAJ30mR2NLjph2ru8dfqHoxLXpXsA2gj74qtrkZsFBSZZUPmpy
K1epoKN1vOHjG41CO+QiUOOWAQj1pQhFGXo81YV7EoN+q1iylouzMYP85p/a04Vv
zqZ5NukYgW71jKR+3IW0cQCdL9cmy/mdtW1WO+qWaOxaxMmlKcM2LPH53XAqMcFw
gg57QH1p1eW/LBkHZH7f+2LjvWMftj33G0u8uslIjMFcBCut5iXYlIuxTlljHrqb
pKYxBTHey6okkf3C3lvrcDhJtWDqdGm252G1Ccs+1V2aIm5PcutQK07e0bo7eDXf
d4ivLOszaX5qb3y7872ACwfHzaLsGAe1eUl0RkJCYFsJoM1GHDEjv5diXfcLbNFU
x5EsFbTqAmaVlYagpM0WPsEbM3prTsa+m5wNIR7EEvzvNd0j8msfDENeHoXq6xxK
3YHKbwAuYDip7Roe8jsWWcyn+I6HQiotLhQvn+pQ4q7zV6zODyM/nUNQDj4cbAuJ
xgh4Y22uCS/LljTST5J65uk0u9VTwER8aHCZizARiOaSpAQgZ04AY9yc94jyWveM
uZAFpN3Cm8FSWw5qGvBCr21BlH0jbP2pF9PtceQ8qHhV/Q1FtdkjLODD7u66Xz88
CBFTrmH9W6Pes2lLIY+BI1YQ7W2YocXL5/5+MECWe109F8XYcfvjlu+BONEs4x0c
Im1TH/JW8QJWk0eqFlxpDVfkoo9xbNAI2SpLoXr8Gz2xa0sLoR8+VzcbEOxE/IfT
hTxT8DHWXjDPX32ZVIuxppowUz1Phio7q60qOEd3uU4SgUxpzVRb74xl4KaXy03Q
9aXBrFFfS8HcP+a2j8fdpqlJmAYUqeSPhNerWEUWHBPsroIhRFb/AKPMthkrqSYw
qj4nXZgg+eIH2nPYdxMtGrZj6fZ+yo+E92lpPFmJiToQPs5hqrjqodyfSjeaUroY
RMm7rrTlwaLr7gSrnm5GtrZRjtvbxWNiIcm8oj3Dn4i8FoxLFM9TiHmXsQUue3aZ
ibZDdyLnNEU2WhW2R3WNjXr12VueleAXYvARbZojWXrNhKO8hmXd4Gx4CWpDUhkE
KaLOcd+JJksqL9J7/ZCB4KZ3gQpaIkBvkVbRv8JY6Q1BUomhE0kMejx1XJT9oG/B
4rs2f1Yywsr7j/ERnNubuOm8KfebiBxHFntBCAzbTonj0Iha1hOq8hHvYqLLATJd
AglWenS6HjgS1ghCTp083MdDwRMNtux+6b3jr9r0RckEU/o9sTXDq0qDc+TB3YrO
0Xkv3xSEZs27ie7rq+si0OL3n4ce+F72nfcRs5iu8SaTtslsd+rbjAFrFwEiWsNL
cMtGjJOiaH6PSzslK2lCGD4Xl3ToIbNwC0HkXcy3qx785jjkwSpw1zxVSNr0ljwA
TtBY3KdhSNZMH3dWnCDhBFrEVSEeQtVx57zp4lXkcgi1ON8bFrY7tOMelv2wTZ4+
f7i0xctrCQxdm5WP8exc5nrW8u22km4atM2pGx1zuYCuq6dy2xC4qEOHd8fnFKsK
Le3hz12qg+hcZcIeo8W6UZ3p2Yng3ig0IL/ICt9KOo9lpSHVkwBA9gvUcRAXKJEq
xy+qvwyQh2H2sodICCDK1C9jCssRZbOv2Tt/lNOfNAA0voIqXvhorFOk2VdY+IpR
EahM+pIUooFzKKze27EyRoSVK/zasEhT1EPyacHfp+ka2BlsNfu8l0IxO54svSaN
TpYStC/9bpisXgCCVigBCPK4Mkcou+4Iacxl52e4j86RB1KbAMmcl1ZKKgchs+hQ
wN14dS82AlefssieNd/uJuqp3QCvCry1PbefEet1HHIjEpNT1M+SF7SDtHBRo9W6
PcsNQYdZmVqIXJ+UJVON314kGFwhzQN2AYnxzHYwyuXZeZLYkie2HGFK7vh4XvQF
V8NJZ5ACuZrqQZfTJyybszie4581XZT0ZvV2u64MsbW+q/3504OEXroYMoK4Lq94
uxl3QbfNxm4M+hUXuULIcOEpwgPITrB36zWCX5dEIlZgOR//4gx9O+WOn6Ww0kdJ
A2iO6JGV4jdNdM1t1aMl8QXbYrq/cjin09mKWgT5bkxbT48oH9C/6Tl1ZHkNRcje
0OVc6qw5WaMGPBoF4Ux/efmkLXHPoUR+pT01TliwZNf1o7DmuyV3rN1IhB9sCGZ0
VzBw7VT2lVjfwp2z/PsIDRty6jprKXCpubE5Zu74hmBX/MbdP25p/BIlJuHeza1N
E9TuMzMCeb/EBSHOXXsraNzEAC67+5bvj9xWrUmehoDI24sv0OF2nBtPviDjxbeQ
ogypgWnyTlMdAK9s85ECtQBj2UtURBMkxI1l2lcpZJzIBbfJD5SM3WxRhXdkSC71
FtwrSUTA/ZTEuFExxwuuW+qija6rKEVQ0IjookQLcXzT4HdBulgvmffOTWzCsc8J
0hKuMmJ5CWmefZOCtKbscUHkPW3PCGscKBFR0iIWFCU1faT+fnbd5f7A685ckRav
faEDKRPmw9fYVdtBf79a5AaVCs/O3fbxOArdPIVbEU9hs2hSu4M6YgrReM5A+O6s
8eZYFx9nr1wPTzl6IaP0kfmjCSvBXTlzzuDK4t4SUh7YuDH7mOGOA+0sw0b8eheM
iqmTYxe88hU2kWtNc+TdHbnmGgNsi5LxJ1DSYmvrp9iEqTHwpTf0wnBffNzX1BGB
sHJaUQYuqZXOBjgOOQMPXdmgpBzll1fPqAK4r3VPuHB/PYPT2R9Mo2Y/iL/u8VBy
oDJ3m0A4xNy3EuhvLEul7yH6V4Vh9gGj3neTJfToq5M+BTrugHIXe5Bu9pEjuyyg
kM98aUUNyXJuEXZYXqGIdY16XeYtawbYPWMG6KfwcjIwYlLwbbDx/gxlL7FZAAZe
VXEIdquUksHw9JVePwMwr8TWJ8TjD0YbY8YPdr3H/pK9v6wPpqGHp31XDv7Yjf69
C31QRRnyFJZ7DAx/uC5Q3OtpBzdglsR1dnoogEwdvEZaW1qTYD8ufzojjf5D0FpJ
C3oSerPNUZwulcfmMJdv1LzgmCcT4XE2O1dtBWy1X/iSk8J7L+4ppLandmTNvKx9
xr8ajbNMrBiSD514oWTATSTEFIkq/YNphfQC9LE+c8jsGQHAZ67E8+iKmGa7aNp6
oOewNiJsNZkH9hmJ674RscbyQM3ItN5vsVPF7ZHM57j0+lTj/zYHBokg5b4o3t8z
92rMe6CNEObcRrmRzC5sJjVB8H/p5JqeNn3n2A0zFqs06SS5ckJ+y+eg5hlL86nW
hMW6mZx9E+pjF5voKMn69f2vFZ8Hko8igaFhOIPSxLUdEnOYU7Mr5BqQr8PVAyT9
8ZOYdPca4Art7Ty2jS+SGJpCiNrx5gHVpE4S3yhP/ZeibAxap9/UJY18pzunGhqN
bDljOS8PkGKTwT4MajFPNAOkg0ZRlHo7OfRq9x+qmPSdjtqv/6Vb4qJvhR5hHJQF
tRo7NcSTQUhSccHWondClDM/kBUx97B07CGSGRHpEptgQuJUTqQAaWShwYy1LFgi
RtUFJMCg4eY2i+7DXpvVG5p/pE4uSnfv7Ly01QusbU59G+lpMKGmRDhtvgxoRDmj
opcROwoeg8yfy9mf8JSTjoVCsOaDo2ewe/8TS6/jpZxqtTY1frYiJcYwmgY4fKFI
0d//NIWee95OhuZaWr6cTqoxBxOV396MRBKLfJgjTYWWJPY5c3M0ndvn4IOCS1/I
gpXSzqt0t4EDo2WQ+df0EW/MizQt/IjhXoYK+mM3muRNlEwwZmcygaE27oFieDKe
5cY5jXq5CuCuyRIzSok2Ne2IcHdQRs+k7Rp6PNMNSmpaNdGkwInXR0v5AdnlZ2tc
Hrt5VcjlFPy+JYS7FQ8qC7n+3gFscldAdlRyRRYDlS71q+SpMHl4KWcq7DWFjGhG
sotGjTk6mq79D8b/m9+VIfvNBgfsvBJiOo7VaN/oqiBG+s3zvvcNTTnylM9wuyHt
9BufxxH/z9lLFbONOHcXnPXRZpHevLYxvjpB8HY7ekv+j8Y2Zq6WzsBVww8PHvv0
LQlFFosnCfhm5cFdCp0Tlw1alAsjIMmUh7VzwMoS7JkrpdhMFZV4cDXi4kpH9bay
2MeLS+eE+wfcruwFiiC14ozN1MUMhFvJQ4DcTvVpj6XOkhxBmrx0ZlcsYS/2E5WI
pKKiS0QEkBg6B5ehfac/iaQ0WrpbEYTvjq7qwyeDWSzIEg5jEfHUclaXqC6QQRX2
FQEoq0HpdKbB++NPyRgL1kBklqiwJP5gxq9nBxDanyWffmChkLg26H+wv5L3Ofpw
ACCaH0HeL6bXjfSC34BzJcuo5VwkBOms6LrqQqgwIBLdA8nix90XEsRcAe3eAqBu
a7M4PFv0uF9VodgRQJ6F56jDfODiK3qw7KUL02KmeCOQT3Y2DLTmiTxrLgj/Hz0y
EGzkscD7KqdS81rfD+0Zd8Vphx8bn3fOyePf7MIzdGL2oKgB2HakZ5FdoXN/TzeG
QBr8MxpiHLrcMSD3ji3Ke/SaghxpgEBuT6mXeavJxGRTzsqlAiiJEO4Ss1Xg6Mto
ylLFQYaWU8jbcaRxsdFlA3hsePNE0rkb/u4ArKcn5ImfZTNpPGd674GFrvjr4Pvc
lUv7NiKqo4b2XBa+hXSSE3RoAr3Niy4hToglHDylqzB6ROol71rfI2Ga5Zo1uwtR
92KLYGA9XqXcM78TdR9KVXIKPcQMeiPHlHx46k9wpJeRn3VF2w3XQOUTkAESbjks
XHa1Yfa5KU+FLlG1Tf62pTZQzJxmd44iv9cnsvquHu1WU5y2jQhwiizrl4cyEj6z
GV5zhnSg980ko3Cz3YhUaRl3hUU8WzEejO8t96gItTqU0pPFrtGpdexM7OFN4il3
eCXAbJt59HFxl3XF08lR6BilaHyiFRzVrzqb8uIoChl1Z1htiDcNZo9K8V50HnjO
2crWAImKCFtAabdJAoXLBcOcsi06sQP5JAGSfniJ/BuY6PIeOPk7ohc66oyAlJwb
WdE7MquSoep2KLswD2uyhJesR10BFAUaTBRNUT/42ty8vOMQuCHOAKf34oDOZInr
SzVVUIoAFc+KbfiMLptuXWzGQel3ugfyGHJosUXCGZ1GNY0rBGIY5O0nX5B2+tVJ
VSfYihvODkBDq1l41PNtWreyQQqwjsACG8W3pANP76iitCkyXsKUKVZzt5XMf+MN
gVJ4yGK9bRXBbqZ79T5IotXdgpJh7EqeM+65DyXKel7jnguEqq+8pOyLM5jpyZuN
RKj6N6LbaqXguAmiVVkcnwgY4lWxGabkm18k1ZKnDWC4dWsnj913AdsUcypSNH4i
ZAh7Jhsy0vGKqtbrkTUuF6jGsIPaIk8opkYyHEAghXLoolBLVfRaf6xCPrLeauBk
Hh3dW06BaZcJvi+sEo8JiX72xn1Pnk1G+nNfRmmB7W9gaZ6sQEEapZGvFABGkbdE
hjtH31kCZO/JULnp9gggCpaeejmZUjW8B7AhLlrXP9tMHvgOh0+QtVZz31Fjuo5n
D3MZ7XXubIz7eP3OWkdMfpPwFJ4+fgqUW1DTZxWT79PoDDL33jTHtN1ZLugW1Gj/
wmw6avp5Q7nQlAeEsmqaCBkUr6iDnG0Zk2NOSpcqaiB746y3yaXzI2RE90I2gGHw
sKryjvdU8izjT8hMps4xEbQuW5gqAj+Ui2kx4SAQaD9TEIMKb1DBJwu/6fdt1lCL
8786ZuqRILmUqHpTagZtq994uPSNxxjFqHGmERlYSi6awCJwbmNWWUsDgfLH7vZz
RrvaYBWtFU6VrfsB2VFOiGmGu9+b6wJcYEF3zKVDCb+/95eKbOt4wcnbikr5ebss
MH6d9Ff06z0tqSMhFD3pxCihqYsvEWh4dLYHHkQB128zZpOPuYtSKgYcPtjnVfiX
TeFo4HAHpMQtRF0pud5WtnSuX/zax2mU/e1hIKUU06KgYCM51YNIJl7EOBYwVCIl
ZFiEeJ6ruct0V6XC413EcYHeiB79LmIW98SRNcP7XQFM3RPaHfr4rIjRWNn8nzs6
HRTkRa58mRK688ayO+WNoDJ/FTKfTGFbdGJvxP5DH8RCTXv78uhQmxhaHa5csLKX
3c4G7jRC5TbGM9bBS/5CAPNmPuoNwyEo2lfSQN1Jv+TyZW30gXpttjZ3qr9WYbtg
N6jsID+cwRvcCAkCOVG7w0XFxu/AsceC7ajJbnXLY3R2V2/6GFKnjFZO6wMlfEAq
KCpoMfaRPCD0PSU2ateZk0r4tudt7ntQqGwuOH74gurllnw6EkXBtq8jFMM1s1H+
pbwWZ1qP0EIt7qCdgZ+uABdc5MwQL9gG0MXBdVfkAfFJZDML/1e1dXnVCZFqk1/l
w/mjcvvCWFTQ7IHFyeocmDWLs1eGQALFd8XBpAWu7P9RNni3igsTAFpqK1DGfv1i
c/cBPZWFsdEiuuI3A80Egdnsgl0hPS7De6+xSbcrBFUUBm9+DtIcV7JfWHLjlYB+
eO5Nh6Cc13ugbzJH6oFeuUm2ArMQSc2KnIkv/wPQ9VxgvIJXdbBVF2/G6riAfZwb
dPYgPggXxLxaURPkFahpKvRjKnFedSCvdoRBlDLu8YMbMEXuAIqZQU58tFspeHnr
lEnD/Wti0efqDiFNY8bdluDgrP7HkKY24K75YEgevOdgisA6n/EB3y8NLgUKE2Py
zHrxMLRfeKBWBIirHbN3zqf+NFWtovTWqc9q+nxK5614ZV4zOqi0KrCoBCruBIW1
JVUdPYot89i2c1Ha9dGbPNUqcCE14IgQ5DGAJUEitlvKYstnb6sYmXO0/KHCPz+7
bJWHbnmwO/RQbxHSzEbj4XkAkln17hGlhmD17jx5SalYNQjYISoKeG8JdYE/STht
1Hv+pvgjc/ZZ3YZb884DBa4HDXahnQLvW5HvRT2EGgVZotyU6qWgYLOPgQbaphDq
CDV5/vcZWEUvyxh8zgkgqhCx2QaJzkyK33Ed0T9vyRiCEJP5xc6ncr+fMwow7Ujm
fWjWCfK3Be20Ta9jpixoaLCwy7vXPmOcoU/gbjp6yvtgHTBMeldlLb4Wwy/+DP6y
PUCWGg24ioq1FggO4FIFDRWcV4upG+eWo3i41jbzeixBizJPOgrSbd6ToMZio5Rw
Xi1BdHpvph+5fenahRXlQ1PthBV3uanTYtxgywnH7tWQMcKQu1YdIBwl5QC4RZZY
+eQW6+UKcKdfudCGfsm4AMbpbbNv6Zy1Du2+Ie64G1mji057j8Tqn7G/k7ioUe6/
pmwLbAnozdNZf0E1WTmZvfGl3G8ny82S9sGod4oO0g1IxlqtPcEOyc2yJzHr9ozE
7ct5FGdKfKsmHKxQPfangaf7K7nK7n0eOaNLvRp4JIWP8mi+r9XtTSKtpgUP7gS8
sJ6Y3/Pnc+pzlH8QuH5zGkTeXL0ngcUl3848nbuDzD+iWBE5FtMK5/G3gq07PST6
oEYKAKQE/5oNWaIwwMJEqKkDV8NAP7XdiFPqqbpM2w4wcwf0WO7sRST1hTaT0UMX
GQ8PgIO+syP532oEXcvUiLb0PLTOvn0gQ5TGxZq2yKSTHRduRK0FmmjBhHLNf0Hk
oQzvsoAV1n42/CKsmaSzgWhZt8CV0t6sAS3n6nXFQs5+Gys/+tvld1Ioj3l+RZII
zDHGV232DNSAqjo1yKiFIMiJIJSjESvhQ/7vdNyniu2VFDMfLyUWNOzoJJLqDFZV
bnSuz7YqZsCACC+iONG9t1n4mnK6JGCdBqyzEE6t7GsJWUcfkKnEquajWtEEI10S
+U5DPyq0CiEp8gj2B4Grs0UgYD9LmgYwoln0iL2tlgSzUiE6mOqqBtvrr3r334TU
u/0lFE+PT5uyQn7rcZGIL7R0Ci02o9kic+3KsJFch8VCfUCCExyYUJjCw2vVfdcf
UpcXcyUCqG0QzcP46q0A1nKNcCLMK+XZy9fYA8TEvzh34rViocoYYCKn0Ys9mgx5
prSsZsR3OgET+KpMd8gmPFfOgL8jSEJosC3fGzVFB2YDKYabuE4Mrl5XyymODY0/
SIYtDz2q6T3n9geOdD/BIw08Ga3ttJyEGEg2CNYH4vZX7cnPb5U0Uv6gLciaZkJp
Lv8oo8beA0hupZCJnHsnzd9YxfQ6mkBPgd6WsFbVX8ivZNwPcWoYoFxXtWJN67Hd
n3Zc7Vfaz98QYfmzcDmgsqNuq2TrLEmf7BcoUJiB+eJTzXjZh8i5tM80rDWtOJsf
wuzlJjB098xvhkVFMIbR7Fz6PftugLS3Vq+HG3T8i58UelyLuSncn4PHAP1zELHt
gVFS45r1/JmuAqvgRUhxuyKJjawTf9DA6l3yvhYt+U+NDH2LmIWxOmzN6W48nPQB
IxFLARK8j6MHz4FjyWk/wdmzrmMbZZuFj9bu9B8bMSbB7aZNkXOLJRXutiLKZ5Kf
Z2sWQ4T1Z0MFBbSAB+tAncbj48XiPn7hrqLP0KwAR4zAMGhBZsTqqG1YLiw8x+WV
doa1USRadKBRTXciL2UGVM4soHGpR6jWORqWQ4315j2gl1r7TU9PeSVD5jqpCiYH
EH8gEts6alvptLwPUrFR/8+2CIimzuyBiuGu93stndSz2rxt/YeJhgbUskx4ie44
37uhjhOzF2i5BIvozPYY7zfc9YFayRg0RI7b7GUKAjf3+IhUfgOmnlOT4PbP889b
lXJJT5KwMBjy0L7zoMi/e54sYDuwNe851bbOoKhl7yZVSgL7nDQHehv1vrZ8Tvhd
Pt/TMkAkH9RHYTpkExDAkqSs9AuJNG/tz7hl967KE8RbAawM3kaiDKOdGrCEXU6g
n7uEExQlwjW8D8PNJllhY0x4Nf3UvKi6ycSw7X6uhWdY3FMm2ccf5p87eWlGAg4s
xPTKcsB9APwSZCbh58YOQQH2E3xVoEkj4InASPf4YkuGVnARpq9I/ThGrwyqg08q
6kEkxC/sG+5AhpSjqJ2ZoMlD/BNjTwn+mMrSvQKs+8RZ4sMnBIyRZeX4swsjcmIM
a8/vgZ94vViwCitsIlcGmOeIl//I15A3dlV4lfXnNLpRsfNXopMjqRBS9Rj8oFCX
4h25TiTuZVEdSvIq2uuNRcawCGUJ+3rhZNes7f1J9nMTHWfaT9ZPjGXN/VmHMgau
5mDZk/wTtqsr9hkRtXKbCuRTqo5vE7enuZv9UOR7kfthQOvTcX8sj/7uCscgaNDA
A73vSfOnu4k1rOUttxDz30eXHn9/FXVqe/Jl1inoR3lit71+xOTNxsSqRJgnDTGV
fLbHCv12DoM+21+nPd9tWJDOEIgb7mPRMFsmelVHwb6TU4NizVJAVBYnd9+3ruyA
8d4FKm6CRFb8A79ARxCuzkWRYsmkv19pq7wXM0L7s+2ucZ3E5VBhTt03NM0V5uL8
ucggU80fx0z71QvpFUrN0Bv+iBxWUryyxh4Vpczv5iP/pUNdwRXQXKwyUYO3Ls1p
+HmqLQgNqztK6LKDou3M8gf/U/UmOA9g+P+YR3guWFsVmZWbyz5cBGAtb+h4ISsi
aRhmDy3jPqFvWAYIlQ7TYTPL/ii2M94mgrqSUbFkIpzThv67u/74f3XuEMJXD3NG
suJed6iofpccHglTDK2Hhdl+GZXvm2zjmfo0jnDjSAbWnaZl5aYWY4SzPBalRgGG
1yp3RJCdw9odncUHUJJbpY0O0rgOR6kA84/L96yPxlyB5jAGOKs+JUj8AhBlASuR
4ndSYHjj0kBeZ411sPytRPtREgEoGtTlrwKe2MtdKIFKpxIMARLRI4B7XrNhoB5S
Tm/oSpwI5qgY73RayyRNP7eznPAh6Jzq2KlZa/i24zE/dZZUEgGgtFEd3aRzXeb+
opuBiIXvdzXi4jL67nHxGfBTMN8Sqm6Wvury2pGo8isFNdFFdkG/g2ElMs7Mq9I4
OsBbfJUks9hFI2UuUuHY1rZpPaNRkzXsd+XR+pjQXEZYrCBJtZKCL1istTY2vurJ
bS9oHHfUWlOxfarssoNWVfQQFvt70Ao+KTiSwRaMl/5/wVT5j4WHfp7neMaA2JOM
uNHL6XpuRXKfOS866kpGDDmfGDr9/XMDltioeMHlUHOdqB0hCThLyEw9HNjvYcpb
LJqLLn1lFILuUK8Kh4PltcYTBhNjmGh3GUJ1ZPm63Hsz9vIupHkbnvN8G4W3DB/c
YfjFx5j+/MEHf1+8d1ibR6mt15FrWn6OQJeAGJK1sP0lFoOOB47ivFOG354ES4R1
3lOSWAHlTGIfZMcjginARx4m6oFcFZ8AR5bl/tJk94TD0XfAItEIotyA9jSPJyZ0
3PBDOeFDb5+VFNMglcsnRysaEFbG8VciMHaC8zuxbb+v///1w0NDZrGfWMhZ6YC3
Vm9VyeoqIaNHoGn518uMWbFWaWcUywh1idhOEfmjLCV0Dv4eYQvCidc9+5J1x3/w
wx9n8U2koEE0LZKobbK2jUVbGxyzCz4V1Gkto5pAVpw8jLjTdMYMgxoeUv+oOaGG
iX88FyQ7cwbsuHrWos5Xibn+pGz8zkQhCa0/V/je4lwzlIvVLQj4YPiSSL4AuePw
okUWpBWsWTpEUAEcIj8g81+d3hnSbYqQcP+dpCzn6DZ6L2NZzR057bakxM0qhX70
HLBq+dXSZLj3F/bNiEL2NMS3jMi1834zzyspGjLDpdGYMNLo9n5smpuqn74nLfsP
tkhZJyRLJbcXNw3PkxLSSkZ9L10V93f0iJ9AIpFRDRummtnivnVYdpjQydu35hm0
txB8LjwGd4Ect6fD6QCGlm9SjEZHytQl3QkcrGFZ1yjhWK6bVKOPIi1t21O0bbXq
gfq2ZILBVLXTLPcXdWQaohMO+K8GaM4rl3cYPJRVpuYmrtDlO7Wp1Qm4UZ+2KEzA
en0j9WaPYvsGmPAx7YRUhgTb8xgp+1s+1arBde1AjS8j08gPRLxxzBCn2S/3TcW8
SkQRszmpqVAPe7mdlcG2Xa8LP6iTPo/0AOqtCraurODTY0WiOMKzdAG1sfTPDH3q
3fo562xoE1G/m9CrgAGBIW6HmmINhlAh4V9ZtWk0Pxd5THJa2VhnCf/PaCqalkXm
BfEwQpVgegg5zcC0R7YJWKoEYRb1wqFkDY/wddIBJCE8Uf8a3uw9d65eKRHmshGO
FHr4oGANPfBCJMyi6GOtXTh97+9VDHHtR6hSWM8DsxalQkfy4njoqWaNgA8NUDIM
Co1nKjuMv3qnQQDkwOfqXuszn4KVQSyWL4Kws/aJWGzTzVi7aN9t2zT1i0VT11JZ
Ya9Ye9/2PqpiE32EZl2GqC7pJCQiYKcRcDaCS7DeWCoOO5hoX8TOkz6VncmsFnbv
iTcWYQrdhHY8OdqpqMwpVaFS1+SrKlKoz3v7PCkb+z6X7XIrBR5JQVaTdkZ163J4
GK9/a//56jumI37W7J6jmRYkzIRG2ELLAEwB2Io4jqYEleiR/Qej4Q8dC7dABzrT
2pW4BPPRMqL/jAHA2AwGKRICmj4yBK0B9OwsrEJI+U1JxVTjyGczZ3ykyg17qnDh
0psYp8r3Y+WapImgjD6Uw36JD1A0jdmpbr64pSLHkO2L1bIuGRXVB8eqlR9baOss
VEZ77YEEQQA3hENax7FowUjAWIdVX8ufbACINIs19B5s8615E3Yx53O0rTzKnW0B
dVdqxRvcUExkDGse+Fe++sqOq4TyphB4CCtDfig1H779f+YFXoclI+7k4lMr16PJ
60EEL0XKhB9OUFRlmBdbEGr6UZ2KS5CSpB/kvNwufM4QPVLJ8PnFhRtuPS84QKZK
DZMguoAOIEF9+frH6yBgkmcmGi6S1eJkh//wTpoc/9+FlXzE0nENEb4pQD0NFNk6
0ZAMBtaskpO8r6npGSApxv5+uM2oYKHGpeS0F+7bTvJ6Uk6BA14GbXAuFw0md3Ed
5ymrbROHR/EOZ8byDnW98OxfSjZfmCZPTJK+xkpInxwZEMSfThu31DSywe7JiGH1
lH0fjw0B+WKroKExwZwj1p+tBn+IZ/J9W2e23xOypCF4rPFY01m3X7RN7nmRhMy7
EF/96P4yOEWeHPZ9n/xF33wfRLy5zutrLPz3mghcux50E2bkqQM43iige3ggQaeG
zcW4oFnZw9z2A7FQTeXWHjE3gohjWflHmd5+uUTv2Ew9EqU7UCv6bFX4xLE6UdWY
oxXCQSl5Fd2Wrtp6YTQ23YasETuT371AWOYfmfhfERVDhfWaHE1Ndlv7kgJI4jMs
czbhFzyuWQSJq7RCZmDHp73HUnx6+TBWSHhJMSGnlIK0oAndXUl1XC/KBB3IFXo5
kuZ1vNg35dRAwjI2Vvma8MzbpZnThBLOcqFi6802oev/zoSNqfd2Kyb4FtEADVdr
5xdqtoydytaK2tDDeC4E+wCwfX2UPDGG9l+GnLx18kVqLIU3W9fwCN9e9qsBtCG3
m3AoPnynhiIpkXgvKJyV8ZPl8BmTuk76Sf0NveqOZ2FUia/qQ19HUjydqVf1Wxsv
UgFo5gkcTmZ1d7d+Yu40do2NjOr+Uf1qnBpR0b0GHIdhDlM43y5vKhrSFXXl+rjE
uI7p1u6r3+4KAenJLDJPNgCc65EvYDN5dnGa9IMJrDu4TEuFJSmpCu3rtsY98RyV
R9sG3ykINZ6Fm1Aznw1KhUGTwb3AQl3nXYCWzdu4E2cU52jrWgMEsMaXuK9E2dxC
UEso/mBwxI0ZTpqreel3YV7UFHW/QJW+mIJ32dBKs7PQvo3foajb5zLt0e88bEGE
L+70d472UPhfnan07VLSBsrYAWb9++MBQcokzj41YoOqii3l8/HHiTgM4elFNFr0
6Hw92YQiGpcwGzw2HQBURIfoAUoQ8dl30+Y0/GkQT0QNo1u+D4LMoVV6zEflPDok
hgg3dAUnvHxnkpe2Pl+di4/gWlCi2pnzz8tFJZD5kYTseqqYfvA16aF7zqFbimiw
fWYwPwUdgGIv5QQ95glidaouUC3moPLnASsnDxDcKqaXyESAKajit9zxLsQA4bWC
32H05CeFHW9MEBwKgHjot2vUCPkeXg19K3dnsHM8ouxB1yKJe/8KKdYbDG+uOwLD
U53dm/IR9jZLQi67s7Y1pj93P69U0EKhgHOjRcrKsg9GlIqLVJamXerQhH3+vHOX
m0yiOQrssPIKpssVvTG1E6vGHAW48bxNaC42Q6uLeuCzGeTQ0XbACjfPwaW5pSNB
TtbOU+rf2v8CS85H9pVONuaysQsI15bblT0ZbhsCr7oKtrn+MlfeNTK7BnBmMWB0
3TDcYqHRE9nj0PhRWz1TevTf/MtNMEW8YtdULOkQKwO33KWdstkmph1SsGBT7S1F
1wAdcPnPhsY6HrMCFLfW7IJQ5giZx8xiLfx0RZFsRy2AdZaun6APYSoSclw7qqhe
H+h6VNNSpAMQTjwI+5/a4cqHTPzirsgBn9SK4EUhx3u6qRjM+X7AcV1wqUnheymm
cxpvR5IXqgWvFlFyueUlUGjKwbd9L0l2S98RTsb7wsbIQgv8bSfeSXqmOdbqT8j7
GYg+9p5yX9bis1kTtECuxjEopXnpCcgVlglCFcBKcPaGkZZhKAtucJ6ECKMyT57a
JVVzkSF50/Dvb1w8OkpzMdDAo+jZAAFXL7oqDLB7HJ/JuAFyf2w8L6p7DSphM/ds
ZBeh8dKw6E7UQL2EMw7b86XEn8zSMaTtQQb8QwtAvaTDxO4wjmlptHdDrji3lVhr
rkwmFOY/9s+LP0zhIwBhXd7JdXm7M7+0s0TtYKsAfZY2e7lPrOzbvuTfeVOWfe4w
+cIJwgu3l2mrzrC3/qU81rHzrDbMdwntLGgCFKzKibq4CiefbSNMcM8pfatLRhcR
hfByiP/1s6XspadBuvvgoWXaJmGmsSjnC3rpUmzzfTA3KzdouGIH4AdzCdMZriCZ
WT/4gJpVVXNYBq+SIxplZSRGy8vziEH2M1gO0BmotKgAiiqKjNMe/TFy9JMAeGGG
lqKDW/7F1rQRpua+ALhJZQbfsZDTyfgHlstJcY0jKgkU5j0qoovkLyR1fuSJDxXA
KZS7WQFm0oxGjXuYrwF7H2nFn4+vIJBoZ8j3O/K8KiTUQfFL+3+ceAzKxTUW2MNg
ogj5AMq0jN0rALFl6IWTWo57Giwizv8YWEqx45zxEeNxkxn+IBIITZpw3NUu8ZRj
q/66LRWofnV6EGAy7SnRoP8GAdxE1vT02THcW3goVXfJrAWyXkjsBIOx0Q+OwEQ5
eO+6FO+rFtwDL0c/jxXlTlw966IIf6s7G1kvC015E560HEPvQdUyv5MgIopjv3y3
u6MRE/EIC+WB+4/XB9mAZWAApI1b/juxiee4XT9XqGr7rLqnbAf4IRQl0qB2E0Vq
pYhNn/owVrL7Cbb5oNCUmPJJAKDKZ1ZXw1Q/+3Z+BhKyuDET8dRbDTY/ssn6kD7D
HTbHI1uvldsvt1e8u3nLF1g4SV/KICCxRND3Ac2WCDkazmYWwCYpUbFo82vZ34I9
jy1F5O+QxNyHwxtENPXtwz6XJ1zjauOgw/7jFOhwFrOS6o1bA4Xqdlz7he8RD9bq
kgQlzyCzY5+ZjBsXPS0IJPOa20KNucHPbClZ0wFj+cWJ5LoS03/pHs1IW3M2ZG3L
zdIyNg2XSbhJ4nnqRWQJ1OU8tOA7m7r8Vv+ooS9dTt//pyva7HHNim0HAM/EJxLr
cJiWb/I2J9/nDp5Z+XfxiWBc5jvDFJgcFl2Hkx+l4DFzENUbITovITCQblk158dj
rA52W7OA/zxFPAaPRQCcoI9pbb1E7x+2tzWNUpgA9GvvX86f4dzF2YRN0ybhMzTO
YCgN1zu4zQyi+S7NgYuSHjtTnD/k/wnoq4y3IGe3uU0ajjhQ73mKPgDZJsSIy3rt
ha181TZB98fZ4ovffaJNoX/RloXHLUXuexXgA6Kie/AWwUXRqZltNsutzs1kgmuq
pWNHgJAn1KwMhabcFkMT/lNNjc7Y5DRZp0DCKhTiPnY3N4+L2yODbRXwjvQ2a59f
B7+WaTTI6p3qjqgOQ//Vmb/uizx9M+Sc0KruuzSfeC5gBWwM67x8R18KGcLyjUP3
WmKyqUSUc39jTJkBkuJqF1cay2nMHYYgOXtZB7QM6W6mrPTV97aBGpW/ptrCvDFQ
rKZr1/8vCZqCIIIs8cuyQ8tG9TnFgYIoT9n8TeWziDZDQAWNILWvCxU/WdcDEATz
Q7S4leFzbCp8gDWkjHyXrTflI5uoXMeEBvZVzXBIuLiuqHYw2dpBqKI5XIZeS/lG
K6Tv7a4V9EGurLXngfUWwyV2KnINAT0wqGnPcoOCgbXCREP2SiakYYuQnK+9cK/v
g9icVb8RQCsA/wxth7Ya8WrWABecAKinJp/9oXL8RFyZEJ53AiNNgy4asWQ7w/M9
HRMJmhSoF9Pq2q84fK22VKZL7BBtqWnzvZXBZOVsC146pPbGMBOFvzgKDUGUK42s
+5ggZDRBobwkQmo5v+eKHFEayMKFRVQPgAZKrZoLSl5xBYNqDkXYAa36L9eNAamP
5nRkYJeMmRUcAdIqhwJlfJoaM/mWXz3pJsqYgHHNEywpY+Z51Srhux4ymWm5KC87
8zYxBKTggM6mcv7F5Qb9FWft7E8wqvVQ/5u83bPHMDPqJyNYUTXt803jtQucSYMk
yhuxSRO+iW6Cruy1mMtXa9nnWrc982zBAQyfcrsBzOeHDMNpb7RrFxJczzYZcQsG
XI7hFFK0f+6fYtywmguY+2y3vVppXleqdwCCC3tykGsxWV1V8rQWqMJFaMayT6YB
P6tW9Xwg7Kw7Igqn3J3oO+d4d716fQ9AErYDNKPkSPr2i491gK5dE6kVjiL6qlAf
YJzyMlgDqTY8I/aLKVsIbVX1GOIAO33OHtTeVpxWwVXyRAImiK5Yv9PbRG8j87ht
ei26VQfNWqhXwhJWRVGYEy842jutDjBxLAfxUJFnK2GmV2wf9rINcKb0bDwHVFoL
3thLt7UuUPYTtJgYo6ywZBISDrUjB9cCOzNE+ScL950gjjoy9O7/5X8eJQrNijsi
QSu9Ilfqjj+tshTQVMbXppm6Yos+MAfWVrQgcEp1yPNJ6Ybf1kTdaL5JTmn3YKPd
WOZTWDB++fIjYmTYfyuzv1kfL4IArHQZhB2uxAvfVGjgS0XrDTeaEQZuVFVBMx6d
+2oOkyTzn4435/iAkcMiBo8AsuuQweT3yA+YxKKKMVzeJjOizrQ4S8ZgCtnhp/qb
ajOmJdwuY8nGn9EDVtcYQ1Ek3GY6gDxo3xqXsgiUe1KGLMbK/dtesbkgYRC18FbL
Qo5FKmLCbuSBIn94Bo3wr4shZ3/SHSLUJbtGzopmy36UWbxgnHj+C3bC/ADHn5Hy
qEhJryvgF4rKJrYWWYghexb571UyW5mpkWha73khVR1fP+8QvDL4TTsOTyOAu5VO
Fup2wB20x9o7dyUn6zuFvlCUU7Yxj64s0RoWrzwvQuqJ4CTgK+xssob8ag8AmQl1
mRJYCNR8xjMm1wat8sQS0mHbUTb3epugneEbJ8+PX1r4O25cx9uv7DulogvlCWwY
i6sa7uV9rE6+o6vDgO0dfjZEPwsw7qM1dgqWTXi2f/tdtHw8lwnEVDJb3ex+Blo4
ng6kvEc5LEMdDVUxpRP9XJWPQc7TAs3egtvWwtWiNuhSf9Y6df+4s4+IWBoAqs1T
E0CXaYTzuHVRmMuVbBS2RvY5SJLMX1rBg566YrvPPIXYfJnrSgqiXKMHBCbQ+PcD
wMqgCPLA0BCvfqorSXGhyVOkhTTGzyydGaiI13JL4I+pMGlUZ+Vd4qrDq47UUqB/
EhU9papF+zmu5l0tbb1lHDnio1GZWT1NqOtHB+qTpuX0UX5+ICSVlyk9ed5Pqyfs
pSWPL5btkeyA9VEacLrD/jmyXzVEEtgfHcoliUG+Nl1z87AGW5cgHWa/MKJxIoo/
o4NBuGQwMpIghTnesvwzHSrsSUpA48YYQ/fnPc7BnpYxAy7hX2IGQ0EyOn8J5DaG
kDi26v4xaU0mpEkxY6ctwfACp6uZfpVcqWOh7jHNHswrwUGlEJqwag6aw6P1Ii3T
e8+CNkcJ+xJRAel0TTvb2cdS+jOiFuHIxVhcsXhMLpfzLEYrPhyfPXHkLrnwTZNf
Cvl+hn+jf4ru2Eupyofs2Yzu7X/sR2whmFgD5BBdYHGTiaYqrMBOdevWQv7dEt2b
vTrcztZ07lcrro5+ylIs3z9Zul18IQ2CtZ68O80lcdVUUOBzfHCL6SjwXa6Ih3MB
c0NDW5+DtSG29qnoLufu/Trt6n10nqxtathMOwjVECZoKZRWTMFVKBwSAkP//G69
nJwMOz9a0QAwaqLySuZZ6wQgcN+ZX4CHnW9IhC0VvGFrEsU95Ng0vK9pKAW0dafB
9Q4xxORszbMWjuzL6heRO0hQ8rXNbSDdB45Z54Ja3dDjgv9LUG4zfQ4VNY3u3X9/
Wf2+u4CGeb5k0g3VJwk9hLHHi9+Zo4v+gjWi/Pm6E58xuJvFK4rgo5RrRtIyVQ1b
bTbEiGRApHf8QIhMqFsTbhNhsck4knBPEMZ16Gh+SAhZQyYwRFrRUfoqalqlyXy7
lGvnXbwO/HETNUs8nKpvrQjRFQjmWzy5CltjKbQ8Ln+2knxqb8o2T/fNQo6FojuK
9RpeYi38QCT/iZEJl8uB2/5VW+8Lk+iFK6ZuA8YEV9Cf7pk2u+pGUN2hE5ngF1KI
YhnrmB98hU449igWl6O7fQy8hD6RdtqjLKd1Jd+7ThUsFpg0gMisqrAkMMuTkGjn
+c0XCf9A+Pq91R+vPVXQObUOE+V7Z6f3MTyUReQYrsIETw+HzoWiChZJq3ej188U
kse2TYaF5BOhEWXP/NACI/zZJMCtzSb8I2Oe2f03eEYkROzFxh2EmIy08Rr907GR
O4SYnuQq/nF7078xYyKN/9uOe/oeVOvvq67ZepFfYsIHLKmeJREYs3ibk7m0ckCt
gq3jY1I5zyzfyT8Hnwur6S/xntbmG5Ga0dz2tZnjSLIBYuj7DyoQTt8Tb+HwKdtZ
ivoqvvdjCiTo5rFj4+FOS+BKtklSpaKVbAdkUPEoME2zcaSI39rBHPXjp6cGmMOT
nyskaVziXQsJki6zdHvO01+qLVF02KEieb7WsCwyYYX5BTMdWms4EAU7wSRawH6G
Inrtlwsv2kr+sCRi0av+UusjiG0X8T7Q4Nd1J7vQXVq/bA90miyRGr1yWtlpi4Cb
NMToq1ZabFICGpOtIN+tKoHpCS4GYkxfjEmAzpNBUumOJN2FzP+aj8dJCi+BjF4J
/TG6ETl4ElKB1JhwgFsYfm3drvT7V1YTxap7BQPyD3puYO/Oip/pnEyhdLQYwMyv
Gl3GLVeNSj7dn5eSZ1nkVe0xAfdaFKFNqaazXKBcEOF93xwhc6d8I92CSCC7ug5S
A+BlByMIg/pRwtol3l2w0vjgu/NOFQPxCh8TMV8jfIy4eGExiApyzPHH8lfnrnhY
y3MuAKCcaRcwfS4NtuftmaPr4pMAIvltaWV4IuNk2fpOOO3w7tGzt7IAYwG3E4nb
cAMhFLkThznbqwmrPqv4fctG+MIVQ0ZoC3vJ8G2mQ0Irp0LH4wqduD0U1EkFRWr+
eE8z0pWqpX+G29+uIpmUfgO4o90idRPo5+/QVGVyrR7/87A3tYun0gsRMGJgCcqj
Qga8GgoSduMui+KB5lQtztyeRhM99GuiHHYqZuHu+8Vv3I8ckhP1frm3cSEPKW93
rnkc2PXOFsi0taePzmRFPVqeMUl6OfrbvK+alkksblDH1mXOgbSNRXhYrI+1J7vB
yXmhCT3Fr808HQetMT8VJSUbnHWVLnNRB2hC73gbs0cupWkYWkEtnAvWLQINN+WH
k8KIiuTd0bXSAiAp83hLbKXDtuQV78B2QD+qqcJf0lrB8/lRV2MmloDBoX9c7YPf
h0EMTaXAIJ/SCSM6TVk9MtaYHJ9pMS+ZfqAERL4oa1sdX/+G1SXp2H/drplv8Tda
tJ5XHNpgqvooUCTDUHPci9/bBNXlDS7zJBWS64dbMPCWcyJyPTRinOGoaVgslCHU
3Jz2Mex2HTjgmyDpgXEL7rl3sg3R3TFGFgtDPdRp89WjfecmvkEdoEO4ZaF9UwzM
7ub9tugzlcMKCI88g/P9ARXW+IdRF4Ej9cCxcyvSI0TZ0ias32a87sM5amavo3WK
h09+e5EJpCKwJAUwFCgmyV9JuGjf93Taf7snJzKikGRdlIOvWYb21EideN8X9GHJ
QMdciRYKSl9Ib5Gtw+g0NTAu5p/sKI3BqbAzZ06KyLzScKPwEqVW0ST2Uv4pQk1e
mrtOZM7u8QnGcFsREnwBPH+ZZK23drgbN84qfoE1/ju+RYakOifutxm6cR6dkGIn
2ke79FEYGrZ2i7OSWfg+8PQIik7XqslFNk41Z4t3FsYQdJZ38BoKDDV5C49nQ8W8
gDXRYFXAvBSaOJSoj7Z42gOZhVDb3iy1y2TFgUG8NqwwZs3XBLrgvc9VEdshN2aq
3szy7plQQTyXxRPJTbMbhW3TvSo7UqYG+CyRRBPGCqINThNDajFSVwxbOtaq9MmM
nuGXvnwIJS1PP+JdalWeSL/+M81iVIq0R4EK8iUbvKT4wGiCStVyVc+VfAKAY2Ge
jtfN4TljrWO9C/+wLBiE7Jmwx3QVXQ7wyx7E33rIVa9otSW3g7S3xv5NhzmGdFpz
483hEww78zJp/w1A3fZ2ifM6c1swdvjNZZYoqoIxdJ3+UipjKh+10txRxMNvJ963
dBcHuPDaMdyxF9matmwDZe4tMFfiRCOakvCG3TbhJKeLOSvj+3LLGEwv4vtA/P1n
02s5E939eJhpiQRs6OJcQ0S9uOQRYWhlwTPLy1Pj4jRFPMV8UCLDir9HmxQI34Br
IqR7i+DtWHI38g9QzyvIhiEwWU8eMSeiyNM3Bkl+HK2Xi/nv0KAUPwoVQrpLyU/b
Bo/p3miIokLmFe5m524CbG8TJu7TrBxJzKCPYLQ9WwNQOqe7Wo+fIfwhIQgUmoWk
iyylKHHS3dlSi1x7aJDyx+iqBVZak0fj7aT85HpRVyjQSuNk9RNTFgqWHhpZ57wY
M4sdUEK78rm75VDoTyEAwsKH4u6E3ucQZN5MvN3wLoNaVDE6u1AOqHp9yW2jHmML
ibDONYDs/7KQ3sMPC4FJ2OIXr+3+VdAqq31uJedK2tiQG71JdBexxVkWpRY6hAoa
NMjG0IF06v1QxL0DlH54hsBOrrCxZlxS+yTmF4LKtReKjPBGMTNaKYXFwU2rOG5F
+FPcMigduiOeMpCgCrLgq1uYOdVcdybXlM8N5H+zK/OG3N4O55dXvBIKPYNzq7lj
hXIQFXbrs/ktt4HO/fNszsiw0AWsk+SvCXN70zc03ef8qu7p+g7ZaIovYet0m1FD
htNxD7Kw6SE/Cp0/xizyhkqllAMWlrDHTxGqLJRt+aezUjUBQaNTlcOmFHDD6xx0
vCjK8VBiY+bll6ClPwaQoItQ7tIvaU7c6i9p2k22ZkEb2tk/A+YagUn7t+w0dt3S
SXLo5i6pfBt3h5IxzSuuDofBR/Hj2ATr4tJjIB4RkLBq8H6z4clXHw44EAfx8NLN
9HV80ujy2Mt0/rQREAurDFWrUL4YpXHoZ1CVyBJjeaIsHM6Ak6Ql4/Lri7KO2g0E
4FcVrTYfxzx/VwnxQtdoWIdAOZ6IizYq9MbKDVswSPm6YKfOb1zvRam+/DXjiAvC
XlH2eyZg/YcMt1LpcY0ABwLoRTZMKITawa9tZcZBTtKN+lP4NUCahHp1nsUJCcD7
3t0ihXvwKvh1//mh9vTtHWUbQws7AoLbcW1K9/vYLrUJXxeJ6MaAYZNPCKFcBw1j
33N631ZPvwErcG6pGLRWoEjaTKO+l4FUCtC+YIlYOGgXKpyOyiFn4Bmp+GbQ+NIJ
j+QtIBaoeWf+oR6L8cLoU5T11CMWKeyJUV7i84830wlUa7BLgT3wmV45wIv2byJ5
CsjrZiNcwvI/xN34tl4GXn44BiqeXxZL+4pU85gQsKWv/yGxCoXiGC0CQ+eFrhLq
cMMdh0LQahlXBohpjhKVrF0/b2kOQcZHCpoWwB4a1WM1Eo3Y/YAVqpWz3nL49waK
lfpfeoOzg3p83Mk3lwsGSyzUndzQOZH9wQJi9dja3A5Ik8ciwrutC20mtN8wQ18k
GfasL0phFd+BYnTiiwsUtEfrvxZ38GuTUGQKpL8G5NjZ/jE5uuRaKU2PWLWGlY7C
XOlmfv+9bGXnxEqenaJ9dQ+OpSgg6YvqEfhhva6YFTFeqYbBuWQ5RRfNeBf+D+Ni
zBgPmfaFiURPDUcMjJHhkdHuOeAJ/ElkhPIbS00aB73zPzmsXELYa1tmrLokiVqi
ZMT/wdbEUMLzQIrTzOGAWaumX5v7XgLFEzmWoaK3OJ647NXDlf69HGeXanMJZHqJ
9K7kI9AIZGXPAEroaeNWze3ziBuGCoTapYWOiLqef6tSPMhtKbP8dPiO9Htz1BPr
OARa+8gMRf3fiJd5ErDUi8Xxf+higcbim6N6KRpwM5HgAp8Qvb7nDKkd5cd3Ylnz
v78Cc407P/t/0046BofSjS6M996BrNbn/zczSlr76a++zQ6kacG+dFpxrZQLilo4
ZVYPq4ER9Ng+cnd1xYHFkwnWTsUT6mbq1jdwQoGhUML8XKHYIpo9P7m/0veB99cm
llh6MakUVxBXrkfDbxR6Ey9DxBIoGXnpNGH8HQLNDEnALpMHLqFld+FZbgd+FV39
hBG21BZY29ItBFWgWCGA5g/JoAK6MEoFBv8/oi8tnBLLBTL4QCG8k9Z47bovxB8U
vbobxYb6omrE/NZmnK9rnxQpl9lw/QxfF+XoPtgCW6zd8tLI7+DjcLizSleggEwT
og8+B2YeiYBH1kfioacbWZq5e+Ba9w2g3I1STHbml+vVYd9RP3tlw7ZWfKiKsnqZ
4EhLo9njugT0SjieKVhP7scVwMsdSMsnmQZn/PZs5hdQbNNED8zpEY6qkjg8Kzwd
IrKjZ1BUeP4wyRQHWDcR0ilLCgjFRwrpv8M9WurCa9BOE1tQPRJ4Cfut5JWtSf7Y
Ild6bCUXfOECc+ChSITYqA5UI8YRAAAmVM1QPGzFVJ8JF6GJQu9XDxo0T75rkSxq
xog4KAckys6bGqfs0CS1mawtfSMHg/BC9i6677BEHrPVQ4QJh9XSotSnmdznh1PQ
iyg6i/Yf224Qf/36v3/dc9JWupVPFwDTxJIIHwae94zK5TxutYnfx5RiWa1bhwo9
5pVWnMhb6CfXIOEMEcd5WEnwuAT4Ev6EOlt+yshHlzQqq1g2i1jB4M+fjiKryTFg
IwKAtAgQFLYgB3TZ8tv9dsRCG2NCtFelW9PHpxRkIWzkpv9R9PBGsxxKiUsZShxX
9iHf3WAvPOvdPktdInjIuaIZpMXsAZ9DSw2OcCxxjF9VT/1eegr+YYyrBVGJ9wjE
1wyndKvnXGAY3ypuVmauVMTXh/PWaUhNCXj6qoo7nNAIx2NDKGHtFJkFnI4moNhh
jXmZNOR9GtbqlovWdvO0ImDy5yvqPWlxQrO5aEHtiKvMSxLky4BM/PIiK4ZZ2UxG
OpI8Pm2iOw4dNO9r3uHEvSgHM3U0AIy7TAuYHFN6lz/fefFEKONPx0a3ujEqGBxI
fAlg5IBJxOFS9wGnd3SDMaEqauCR73yl8YIT0i/XcxBg6GlBXWbT8kcIx4Kg8z0T
OQPfy02T5aEcZOLcKd58ezAsy6xj77euHpyU/dIuy7JtcHqYuEsHHp63By1eZwkj
xyA00EAMF3Hc5q4ayUs/2A5YcUhPQd+wgtijRJFQ94BF/4tHagWo9uUjYuEbsWFQ
KfqGhe7u8VZm5YFNIGVQvmd22ec9mOtqQyi8KyWWGI+avL3ouRWDMAeQhKkd718E
AzcfzD11PD1WumVpe7v9+WnTfR2Gx/OvbU15QVTycmiIgEzodmscyG9CqUbXPNJu
pABuc748auSSPEJyXUNaNQ2YzGgwnBsEvD5cnXSx126spVasfjQajQdPyxQduaEZ
DSwx4pWDExf7FUjKa/sj6V1+d04r63EOvlH8VmuVFVPb51dwnX899g2S2Vpuusxt
yLV4Ti7nrCdyRGB9z1IPAYQGxyRDztR80fJsprV5sURups/iO7nFrOs3NODaa+Cc
LsFsKByg5DMS9lwUYBzyvWSHAokDpvsWs/Rmy5+qekuviBZczAnaSfsPCnzBADCA
m+DAE4+6ex02GL5pmRjHCsSAgVo4A5uDzasZgoyFP1KcqV0JgrBaitpL/Dt38b8l
aQE+Ypgusqi7lwsqZzm/paj6HlSIZD7MpKn7QBMwn7yOwvF2J/2cp2MjOffb43BR
6nnvlm34Q+UW/+vecNvOIj3FNGUR1yNiqMA8+B0HyOfdixKM4W0NtUVbcubke5ZW
dADI5AF8+2OBpt8eHxKs/nOycT9d7RIfHkqIwOgMZnXDmWZOLjpnzzrEwcLgHcjg
cBkmalcaEyAQnApBHP3iXLXNFuFBUAIMu2ILyRBOQ3WeIqLoV9VWTLL7bVOWcFtg
SpGPAafvoFksDvNjLgmgCReJKYknE/XqQbD47hkctHPDFIU5Li95jSgCTtiy47h9
F3jzQY8krekzoVxsomTfA16PScAFAlGd8era5z5SIxlcQHCyYQXSiLLADOpADR0R
NMQaz7dFym/ZEbhy95s/auSeTSCEsqbkygO9VRVBAFBpsLn5HYa2jyT79CZYkcd1
dKUlyTqt1Fw/mskkYL3E8k2QF2jRgnRMNcvO7PmretsE4dIqGheJ7Pcmoigf5x+4
RxgyFu2d6ukNGK6byn/TGdyUKt5Dtsb+6QBvskJwS/EbidXdEPwYzBs7wESbLViD
DhqWl0A1hGGaKHMV0PnPFeBzAocWuqyF/mPRa/1rBktHd7GL0RT2wFV6r4oV05YA
cBc1zo9HYvZ5KY1l2pn8bJL8T7l3ORa6O/XLYn/DMqt6FuA2rDTvAZvlFVqm3w+m
sMrO0OgRqWYUVvmLg3Zg4Z1kMErGhWHM0yMnmmSHAEsic+bicq6zSwyw0Ieus1kn
iwtWEWhQQLsONI9SjQjnD0bHtBmSkoxuxnIm0cP7R504hYtxDNhjJ4koq9QbiuAw
gFYpIX0awPIssX4PQyxZNsP4gwNWgA5fsRPBrIQUopY9D2gG8PbqO9V5JBbbPrqm
6qjUZ46nkFE00Jd9WRN7FVNGsRQIFMlsjM4HnVsQirXQZvQ/31mSG0M7WsXaZ4bM
plMbPY2iB4BoKfxth3lmFyusGJHc6XrOQzAnzcbThz9GWN6//BVuYqdN5lnXEMSo
NHR0apsMGyo8hUFWGPBxoNlkXf3f0SkCcjEDDmt70bHTefNufLh7rjnouTrUTbHZ
YtTrCG65shhXX012/ZimpMGQK8a6euamD+ddxsYquYowV6tZGWHM5DnhPZeo31CF
h9HfzXdlqFRvBwjtwJsl465IPJrUWSVLl66ZJNaA0X3tjpVS997XT2B/zQbGjtu/
LwP84bmNdV6OSqDO6oMTals0ZDruH+PtJOvF/GkJsyRSoqftriHEPiOqZ8l7tjmR
IcLOir2H+QHunkmcgZkULBxo015LwvOm16qga5xrO5WzSleDRxdzr/3QK7Hna+fi
QUOUniuv3+kr0VctnhO/3b/DmcCHrCnVs5aYcGeoQrGlDrgx7aNpMo0iRi8i4XUU
3pcYmFb1lAVD8rcd/Z0C5qVpnv8uk2FsnTA965uQbQw/zkrVPhb2gZd6xGhteUS0
5qAucUF0bwiJ+oaPrjAk9tpiuX/dqMIUs3CXtVR2uZPf12GBeSU3gISms/uRvSTH
g0sbevWhtSExFZZZG6gNOZJxHWfNewIiILnOppQZyz2JIfXtDXIDU9WqTl8lG00B
9Pzl0jpo7+E6YG9ELvz77fMOxLD8tZ/+d0jOnhloEQ+CKk4kHKGe0obvLyY3pr3k
97FK4Pr4bXdc/8d5MNyFff+iMtTgvK/zR2Zk6zWIiZCJ7wazvIQnxw69uV0n3Eta
XIamvSZ8IHktBpxwurXJ4uBcJTOZrhs61hFZtBkRlIVdjMGEE755yVj5uDpoGi8A
ewCW0rnsAxUV5eeByJIzl0SUaXCHnGdTpFrvHRH6ice63HtGVaPms9ZTb0j54/ca
WHbzCFQoAqV7vCIBJMXL/7EkBc/CZ8CLyGZYQ4irGpG6OOxbUs9pfB1K7+jlX1ZO
271OH0YV0sE37yLAqgef/XwftsWn25L6/UNNktwPPWS08lpeqZWDXwtHUNX5oMGK
qNX3Bs+2yDaKNcFf5UK4sv9WTQlpc1Ibw6K+edb2z9zcLse/tJzebwKFrKUPykb2
zR0wr+RBDeXXIkn4sAV9BbAwtXaH0JOA0wjIa61PsDTsGlSgFdyXly5PMFh1VBXt
4ibSMCtKSU+G6mGTSpsxe/QDK226L5N0N4hN/+KBL/mUiNvWmFatNymhfHBP/l98
NwdmxU4s+U/O57dQctYRP26JZJsngs6WjRz0k12MbeU7p3iI4NUbvXlH/ft+TjEB
hULp4iDcvakCugVopYY2lvA3SonDOfwJz8nLcf9vO/BCVwwmwciaZM+1jATO+zJS
+IlUQDGgIr+lO2YUvdMPiM/w9uxh02hj6pPaCRpoYobYglubuXhhqKcwERYiR0kP
yIp989C40E+5xINRTaD/EXRsL9kche9GbxDV5n1wvAEDIfNklAauZ6eOKlrVK7nH
ZqYBRZkfk+Y5f+oi7729+6Dd//3j3fQuEom/ySUjWLXYf6Q5VvRCuJ3JWNyjY5lW
pzTCIT5A99hHa7J61q8RTeCPJssSMCtwZOZezB7YSRSXJxyIWSGAAKDH4lqgRpUN
YW4eocHzrIJrT30Ut+IRdzFJMu05nQFNDQNqzPDVJGd6m4MCPX+Xo9cR3AEoPTqB
UIDXvt4zrDZEV5btvag7Zh1mA1JUkwLmrAuW5UYgALAXjV7xiwnDtCba77IUSVNc
BSHZA3mcb5BD/HOa/z4coVrVhHIUIRImbw0TDMtHXbIb754YsjoJMVYSCArXObaL
DNlywkKc6uSn2XiOD+j/w2DBrq8RR2MI4IepdUh+KyUfr57tHVeNZLuhu2B3ki4c
GLZD9j0BQM8ygo98C64OQHsy/tVcNkQmTnegg6rcrq5F2JlNchahtSG6pMhR1anx
+kAepv2bNJ0iYbg1sd8pZkc20PvNyJ3YARxLK9infJmR5q9jezh9TkrWRR97xHbf
ktlwIbMEYLm7H9zDkd/Z2q4Fn6txM0S6vMCPQUsh1mN7QZ21fNurTTa3ixVY+ova
g7dD8RZ6Vnc6aTKnpiPxBsRO79Iq+bWOtFKY/8vUOA3MEFBrTl9nKLyhPagaKXp5
8dvePWYfUfFd2LHquSO9XuxOzTBVEn4tcJ2kvMQw3E+JELjrkHn1VmI8sc2JUM3F
3sQaB3hTTYWYrn5b0ybvRiSsUu7M94SDPWSljHDS1GM9p2+AoyiMMJtxwuiq36Oz
p1Ia3QvRrwqqEwKDsYa0qa0R+SZtzhj/f872kENUs9nOIujUNzDNCgViQGn0WTjb
TgiyvEFIwSjP24iBNXZ5XUUXMjhjiMIyvvKEgs16hKZDSUGt0jxzW5bnEVyd4gkV
WiH12MyBKfMi25N1jsYylp4+NynfZnC+cXIMCPCodUd+WjBceeMsJ/hROaB95pSS
FcRM72lzXfFfiTuX71kIbVoNtLKQmlJUnPIRMRhbW0OXyzH8MY2CaKMPY7v6DPpP
mg5u+uyUaCG/o5nv48BOs4tovDvcIF+BM84hzNA9VKGnQZs+JuYP0WRwvoO3zvhk
C21SmlylGVsSZ8FvXYEIAeSySt/lAwTrlZ4KhdOU3PsymGgG2STyYi5h9DRWJU2A
FcNztHTMQ9zHV47TX+Jc1mdfhoJw0GNwMhcj2NuU2HblFaM//tnnfrimUW7LcFOg
CejuermbQuqsaKBb6bCsZF9RF9P5mKFiKQi3OPGGmmS5QCOrJTZOwQcwJXddvtec
83I5RyJ55FSdEUpCWf5V+ckQM/jPry4ShbFWLT78LUbn3XWsEfTaehA1kcMjYWWY
MV91+RUT6fjnZW1qMH4WEhm5nRb7zfQpSHeZa6/XIubjOvDGZ84Hr1OjYJL4xiLS
GSTiz9OqfyJC4uCZ/mSwz6B7R/xcmyYZKOTL0o8bAXWY9NYQn+9rrCVy/ZJKzJQA
AtEvAgVp7kBMaVt5sPNDUVIaoBZSfr70mvlFYl0szFLHnHUPd+na5sUSj0TC1CM+
ZPMJtomwP+wx7BXh5wwpKAkIzIkISSatJ+rp1DHQAEcPpDZ8zj08HC67FOo19jhX
q0UO1Fnl32q/YHrQvIAJD9z59i5DJWAgwyFIQaVCO9OdcL4XelKbKA7DpkN01tQz
jzl7N29WFAhjgXmWxK8aLZQOcz0PF+RdeWu3JBRz04r8a7xoffZKzkdH18g+pUbo
Hvh/b+w85ShJMJKjzjDRB5RrEuNo0fW//qJA/yvuAmhYavaPPnsksOGO6eS4t87H
sPevA0v9/T+i9797G5ZeFqeG/ihlVYtxvzn2iW323/GJAJEadk5Tj7mHkwKHt8O+
czVFdr2ihBcTXMG32Lw7xX7TE7DLxugZ+yqSOuuF6gC/77DaF69aoebbVGmRnXLH
hknp+R2Hv7QnJeafGtynXSqwkKRJ4bWyS0o0IYVBPZaWWkLa92EWWpRnUgVhHsjW
p7dDb4ebN2ypALQw5WDfounG7LwNj0bcGqE2uxCOL14Y4A56Ge+tcvf6zbfBMA1/
3HDDSPLejLupejYx2YThCo19DJhFGi5qiB74V2KywuxPeHagPXkv4FZPy2rOOUAF
EPW2P+02A1dEQYp5hHDryt4TZJpSVmWO9MR0WmCBu+XCMUSPSMtFBBmQod2w+lCt
FcWe4CXyNVT5JwuSWVwE9r0jRvxqmnykKyO+uGQS9K2I6EV14nxJTMrlLkxsvwKc
BHr/ODpHjtSAhaG+wU7Tqn0EGBC+xRnPBsBRAWt585Zc3au3D26LKsblBr2xzE1i
Wzw/+8jM9Nb9lnmVMTRVnQ39gSW8Hl0DvYllRDrS9634noRxuApUdck2OzkHgKEv
hu9kRcwmtVl1BRGojQa3p0mZXP99Ui1SvP3OcFPgYB1ZWl7U4gcxXhKyBiA5S95m
+X/YApBm5yRyMgJY7hw4Jej4N+KuGZn+QzYjdEelpBmIKMTheAswlxTMqoSIpjP/
pkQ3DK8N+WEauXP+0nsrFyzH5JgU8BhAiSobqDM0gbAJ/wyV8/l3ye9dcWDFtpYE
ol5aQDzi82fLMSJLFuIdt4vuXQeigIjhljkWXfcZB4uUvXvFxh+dRHeLGX74VJts
8Ppo9fxSNf6gf/yd15aMMSt1dBeaHsv5eoDMZ8N0NnpDrwNwuvO6XvbIrOC/0LrW
tSD6udVH13Cj80BQl32WJCAj0a2xsXdWebN4IMN4LM4Lukll1E8oubd0uUD/sCzG
J3BvpJf7WAGxlnyeRLVbovDOfZPsbwkgUr+OzlI2bYQ6lp2PA6CgYl9XVQaso+7g
6kmOoANslM5Cui6ZoS5Q7R+S6EGTsJx7D7DkoVUWcPvsIT2jzvHbspyQYNgxDTbM
8fzq7pzTLOWF2zBG5QeN42bwCRDLwwqzUqroZkiHx8UWn+FVDu8KocrC/CAWByL4
BEWUDu62YEw6V+fjo6yF/JJd4EDzoSewSYQworxKfWJS52qpOhrvlgZEJGGjVbrh
2cnZmQiOJM2n4GhvGCyDwb0XrIfT2F1BaYd0foNIIOz4usVt8Ea/plMyr/Fx/PSl
hZwEHPumEhqRCvZubhZ9WH/e3t+1AP1GJYo33r2O7jKzV5reZVgOeWrHU/pwBq/x
Fy4jreo9gqjFofLXWX34kjGNpWXcL3df2I2HvGADPbKRDTVRgQGRbD1V8Dx8gxVp
tAecQWunFD2sgKWI7FR/ZwvuUwNWN6NQTF5l9HDevGrf3FKyZUe65peIvAXvtqUT
CVSyJHePE0Ge4WAe7tGMnKecBn8f/bYehoRHsxASf5WBYhS922lf5EGb/4GyZZzj
P0FrH2UJWS+6a+3NpSULite/WeB5TisQrHbxZ/YlgKoIqQkS2pRP/M/hTLPvp9ch
bP16I6JrA5HDuUxshurEdYrbkRfmXr4/GehkXaJJJIYyXPRRn7lQTTrmSfJqNo5R
RH6D3lKafdiEFOxAGJNNODXA27eaeOvaAcs/tavCjrGnNYbofT8NSBwTJRffGm0F
AkaZrEIBQ1LS9sHTxhMnyB5pzY5SS/4mxo645l+kvuKhauNL3TM36NUjt4/S36Cz
upwZrKfdpeeQKUIGfPsL9lyFXfNvtjDLXAX8JQHvs4YwQ+uRvLFbcH6nbtOXp3AL
MOFNZFwA8BeoTaSFbkDE5ERhFxuV5M8kTsXBJldyN2TCjjowX0RgU/QBW2JRpRvy
/gj2CC7rHtHw65wSWjNy/Aw316AO4nVOLN4xZb3St/EbgKDPLKjb8mlCRpFM44Q6
li05ww/zOiTjKfuBjYb5zvWoxg9nneEaewtSuG7vuEZdcBqgp/b+6iuH3yJT/I3v
C7BN4JS/XQtjUbRfKzVhUz8XDr2lwR6iF6yonHeSxwFSkssLzf/9yoX9Apa9KPiS
lcoqshGTlzsgYffmIwplYbeGRXgMSctrf7MpnxfatAM7XmAvoXdn52c92q0g+05Z
0xyR17M0tPfeLezPGd0CflQcXiZxJ6rrpVqFe4VxKC/Bpa6phVcMfliADSuxgPE5
FLW3rBsuxyl4lCQuF19PPJLESaZwqIWBLWH7EbQuvV29uW05n+1jL2/+OliEja9Z
ub4/SpOdRzbBAZdL+eFyDKZw0enoF7glIATlI1tnnLauTZg8lDsIfUMjVT8JvQIv
r9L6BlhnRsv0l8hb5/aOkARowP1aKnh/GJIwz6wILnCXq/ychfiEKbxxgWxileZ3
PEVqGNUonVvxOXjJZqI8Rj+uIcUS1wh4hj1sddY5lkcZMoUM1mw0BKtt9FpRX71Y
XUBhmJirszY9zu9Msd7/AHpr3KgF/M3L7yZpyCRAzQaR43yHpmtIBxKcJAwaWZ5O
pN+wkiGYOEclc6GJDykDjfZc6yCtoiw5uoaID4FfTviAKyC04cUqYvjf0VVoX0sG
7tQfcV39oaG6P+e9zEYSYTZ7unc8ODXWHj/XC7CV/NMc4DdawiP4EZbX87Wc+E0q
KiLNXL9n3kOWHA4UFOYiFaZ6QZPnlRXA+vqbJXvZrghsMYVUJ718UULtBq1egyWM
BsrDh3jvJjW/+sQCPHF1ERQVyDm+WcfagHzy+A11DD4pwiKIcYZCzdPd1+buxNhF
od586O8TlhplF33O87SRQE8MNzskL8MH5AmPJxuSiHAdYMoAYQJgyuJN2YSSXVuf
fQqUH1Fm03HT1V/Z71l7XU1UpLxtM0JBtsKpTqyJsrHCcoFuUdzeObzfqwrPfz1y
MU+xOfuac3cC95Gn47ncx/VUevzIQsuRCVrrqa3KEwAp4sMylyPRqWzaPOv5P3bW
THLHzW/ylVsEzvWL3GtdD/oCPFLESHq24dD+pRLP4y55ZG149fNYIhPLMEdXBy2s
mR8lH812E4jw260YnF0eoiEhORAmE3W3cWTFLnZJIvzyHSRJgRgWelUjk9zPJykh
poKU/IUj2OJ01iSJcyZAIr+vaMAL/ku2pMnm0eWkatx/WF5s/U87Y9T6mSuxcjuV
EQIDlIZQUaBmOCMBNxxHpO4w4SjNhKaRShXp8xbrZN4KS5SfaZW8FsjThuM1C+nv
CqgdmhC3K+XIw7i6FLOCiFs7NBU1A/hj8V5I5o9sHojMJVcdJTcFSuid63Eot5Ej
5Ct22IwDi1Sl7bT66aI91meQcZX5VnhYm5ZUpsW7gn+DurxQDHI5YqK9g5YO/B23
x/9QuQ184a8QVAvfBKZwtAOAZk+NSgugh7Z4XuZ6gjFSdAlCoiXBXbjQZ7fwKiuI
x+q9BZhR5tp8Hib8nJa4fXlq8WZakI9HfbIlKZEQmosHoC2lXR8Q0S2H/Y26/gBd
pwW3vofr+RNyhBj8RYjGmqF1jMt9doqjONfDGX9tabwREJt04Dj13hIaMFEMOnKM
T4zt/Tp/F0gU+wfeI6K1eD4rAsHzs8ecQnAY7lOk7qPj1GJYvpuwarR79sFvKZcm
uzVv1SYQRnF+/p+PDUVQXa5g7najc/J1XvwaWcmz5ej56tECpgiF/FqggziamHUQ
trZs3kztqMwur5Y1TjX9I81qcF2ohMv1hwzG3H9aQxZSOeyNMJa6GUqioJsyZ3h1
FrL1s+A/y4ogD0pwOa178go5aFYdhzq/ARtCNDHIqCaGXrjulu11XbdJCMXrfDDF
4A/N/y35UarbOPZV9mvdwB5btam6jpnCdP7FXxGjJDRORojIF2Ry27qA6+mnCkD9
Z+5BnfrO/fk9rTHLdgqBFhap7spuWXSUX0ERIQrQAVGZf7xDVqmeVEoECjaxCIC5
Q/BZNJ97qdVS0QSzBuauIIuwkQkYFpfm2H5K8oS3Uw9e82BjpnwOQEi3A9oIEstq
UA30Ecy3MeHGppc9qebNJwziaDD79ahyFq+30Em9g1gxyhaN+KGUBYHM2zgIluth
O1H0zIGrqrzFuZhro2WBLDiFFYDCH8+cEHHjwM8ICXBQty+txjIxnwlLHHSfdWBd
6dZXoh1aXryL9IvFqZxiVv39UqXLkZwTE7TDliL/xQ10d7YrftY0b0Gy9eJjD4Jd
sOTmi6nNpoMOi/ckaDJtpnDfu3c5lyWSgfGjk1hMO6sZzA/PtyLY30ctsVLz38Km
o/5weMeZfx3HHVk2majbKzp8x/zcUiV+d/ybq7zmBc8dB+FrlrJC1cnnpOLuNV5K
HemzHOmSIiw++kFjtybcgXQDpz1WAU8wrKg2tXEEDwgt8ySY29mw1Kf4SnVW5uQu
KXhC7Lt3bg7lNlciD7G152WZLZxeYPkIWbH71+6LDbmWxztVASNgZ+AbL1FkFivF
zvDbikKqNqIGY3wc67He3XKIX7aXICcYPhs16aBaryjYoTqCzxHRzfBd/U0+UmVv
jjhnZ7ZQ71rOJiMnahuXzeU+8QQ1sCe72sL8SWHsRPd5rZdnop62PKcP0kSbPnNi
5bbBnubFiAhh1IFLbj8e899rpl+ZiWEPxK/3BgZPTWx5Afic6vATOSqAPkG+IU3G
Gufa+m6mz5SHOvTP8/5bdFnrjaz3QBtGT43Xq/OlHZhqwZ9ITiXt2aDYs2DFJ7kM
ApTroZkR4ShXGxZeuEy1pR5Rs7aSPo8N3M6ENBAUsYC1V6r4XywG//Pf3CU6Ok+H
BSi3s2IiA4osfqN9BuSyw4v5M98YnFa1pdwMCCad03YsqOtsugHBFIjd4Mj7nAph
AK3Ik+wJVlP1uqjvNTnQb/tj626M8Pce8LmzVs10Vtsih6uJBAbfEL9tu3HtvlCe
O5SFS0f+wwuTZH0dQ16rTCkjvSrocsD0dhhAfV2poUxVaikfgtD3L9aH29CHnPRg
cnyp845kTVRKUjFgcFFMA/uz71iTIh+rfC+ITXy780NorlKdP98tGi6sXOc24KFu
oX/gGrsxAlzQ2wGMuVYVGEPxGZ14OWVFSHEkhrRYe93BBjBUBjdwYtURFI7iYGFa
iDTGyWMloU9d52+kM6WF1X5YfcfRCeVoizjipCEp3HzLYFm1oOpMm9M47nJ8nDlb
/RJQrSt2Q+eAQ3gaTDDgi0SBO7ei4wLlbRWlnudS0qPlg25NV1ict2+4KcgEaKtu
uAl4UFUeOUDEozHQasnJrMwR3IY/SCdzBW76bZHcOHR+HYNB+QxBFr06V4sb9A5a
TW8VnVg/oygibwW/qcq8wMcEnfNxiTATQUjx4+ERK9oNIMGWEMMEQEviMC56xVmD
xES8YwrPLzIkY1ecCCMhrzbeSZyyYUJvQ52oVQX23GepY5/riguPdcQlVjvvhdOj
EddZemEkkkbgNXpZ/2KfsUTniA9WqcWI0qt0zVFOpCo8o3UAC/crefoGEEBODFv0
8hoH/qhS9LuNQCqxMai8CHMPYo99h2fjEYWJZYKw/jrRBA5elp9fjnaN5tnG32Hk
E2RhejOxwUnv7Pf5S2mHtaM+Ne3trJjgehGcTlFNfYdRVs6veyv+N1KWqMZFNQC5
Gu8CnU7A5DA0ZcZWAFtAug0oH/6YPyfACy911furDbLWRya4ztJZ0RjCl7nIQ5Ia
g2Q1HeZrFQEvRdlPL1Q8xAfHHtt3HopTy0oGJ+0sYHEtBrSicEAaT9pm9DunDjCI
eahfREt2rkZY8t71xHSaUr/PED6ruBjn6DGV7QADOAtCi77HtGvBZ93QaV/KUUnd
kF7nMNafXOrTNUvFqYY9Zdk1uxN0Q2WLLAT+W5C2VnCkubQ0NBXXNVALb9Pb3rgW
m4rnPx+lJJOmq3v7gtP68fWXwH8sCKVFfyVdwbUaKWgYcLwAebGoa8agd3kek8no
ea6zQVHVBQWSfRNAquEcPO9W0AmvhagFexlmShqfttLYItFqp9f900tCXvk8qhkg
pssU5kNB9g+RmhXEfKXQtug67OeF4bVOu0TqbEqTiyd1NC/loOem+SuwFT6omF+U
pgPQElqO/F+OB2iG4+P+TOI+5jwBnNuCr/u23QuQ3LTYbdE8HYiqhU+s3BMj5npO
h+hrHai6JF+WPV6N12OWM2pH427aVvHMx9KXdGr6B/QirmVXkwhd9KrLSJO1kXSI
hNZxGQok+t4E7ZuHMmFNkcecaqrafDm1/9iPTPHnCGG0Imdp4xq39y1b16lY5sSy
1cxwGelivOzIkLGuGMDe2Tkb6v6Ns2NYHnKVD5bmkQKlUl0T5RFfqzgnXxxORiwg
3iGL7euX68p7lLSDjZaMFXHhBHtE5s9KlV2NgRKdOGHbGwBlH+YowUGDo0hIku44
UehpkxxgblwcTqGWHZQot9XCzIhprXOMuwtNEyoaFDFnOoliYZvPfEvsr/5FZf9j
jfchIJfQbRqByoey7rznZ3WOeaQaK80soEIcuXy3fwmop4/kTQfDTU2ijYtw+bsN
1+AhiXgHH5ePU6cH0xoKBPw26w0vZmwltMeEfMpkvIZWDO2t+jEAs1rG8qfdVSdj
LCjkvlL8YU+EF7q3RADVLlTdiy5XIFsIu7875e9B66Mgi7WyG6Ik1DqZXo3Mn9vj
sw7Y91XcYZdi/4gHiQrICFxwB0FEgEfd5HN6xbn5JZYX7TlwS6QioiQx21cHsPBt
E+oKznb8lZr8TMKV8zsXnmxW3YJ0VmBRNKkXBxJDmtOFpP4LWBSbq1TqcvrOD+9u
q9oaI5lIA8jLGTFxO20XE++V3xIo1OTkgbiYuZYpwtSEa8LfxBqOFT0Q0+shT1Kx
QlUKrLDHKdm6ifn+J0mK3GtfJdQDmoiKl+HzXbqkKV7+WSQGKyseOoqEILnUMCqI
DZRbYX/xlZIY37wcBo9T3BtUWOyS+lfQbWT7FlocdcVF7zKKdhi2A6UllS3VZET8
jrXL3qKHjY7sQa8B984/HV7TbGaaUB9yj+eHdaQX3gfHBM0ccQqOt4fvQOkAZW0S
GIXGtcQ+gyE1J/08zYf3njw4ngoHHqxD2U7wSpLSlm0gp4WN3+Ds4k5kmPAj8R5a
hpqor1DS3koh8oQWT3nj1NA63zHz/W4ZXeoANcC5hcXVhUHnpmkmqpJpy1MDyOSa
qq+yfTdSO/XthEHcFGBAr7fPQ9OPA6e3PDZH0yPVddED7KjYCue/dPgRLFYESXjR
NlC2ZVOdnEgXmr298u6bqQjsI5hoa67YMNfTjps5yzlsO/uwAKT7/1Pdty8ZJJa5
GW51HYLlWLMAh93takTUNkaSyJdKnGruKnVsongCH7IC3bZnyCx9S7FAoK751zMo
lQ1C95OPHTFF4tN2ty60IT4xdywSBfFasKi+d2ZIb9JrWExm8blIFu3EieAV5JiU
0ou63fMEHArkbJtuOKb+s2WTVl/0yOzKgDLWIv2gJTR/4RX55uprOgjmiuWE0R8j
vuodW6ypZY+OqM2mq+J1UC5rVi0wBu4JZmNCjP81t0Ex+rv+HWE9E4rojiWlxFr+
wKsgV+Dnaq8Wn0f37xfMC8QYufYDa10MfQlQwibnSxajQsbY+OqLeZYSCBUsT7Ge
3J1TgsDZfrzdvwfJZY6ymNsnVeVJHOQdqA+C2De1RkuAOu0V3UjckFoPD7q8WBpc
1qpSxKspuda57KFCYlmzLpPeJi7IY4+L4QDkY98Z3CLyzYFSEGTRzdf4VuZQ393W
V5e4UhrkR3lGIXOT5hVN+3EQ17LzSfrG/6O4QvQZC60kPGIK2SWS1Li04wgoBgkZ
lkyMeRPGnnQmoMte+dLy7Oeug56Yg3rnv+8UVhmq1emEk1+WT4zXrx9cFnKyYozR
E2Lp06dIPuxlyLheQ0F/PEL5T2pOJfSNAJ8R3Com5a+bgsOaq3kR6PU/L1DjbLi9
BozawtU6wZS7bo5DvzG4S7P8jk+B5IafuzT8uHzZBxPyBz3el5L6PS4zficJ3R77
4L4N/e7wsArH0vp9s8bOn1VMR35JAPltJWKKTkcbHm5H4Fee5jBkx6uIJaKF4VOI
IVAKYC4XLe9Qz4hq3pQHyFe6wxMbor0IMmannaOe42YFeAc44UsZsVlZZTMSI/K+
RXFgJQXOCC8Hnb8gClsk43OXsHr+HxVr/tMwULHzHVV48xeP5os5KJGAMpnZbMB5
7cLmEGFmF2/fnqI9aU9VEXUX22GFzbBfiI4fwHTqYtaHrmEbIuRDycY84H3KJi7b
298l5NYX89OoBON2yRlrDHfSJKif5C92nw7v8B7DBBr6dU112JUJ9n5+PMgdeHoa
sGeIri+NCDbX/JBw1HKn24fi/xj9xO7b1RK6P5EyE0oPj2PEjVEcdCiCYAFOg7bn
FfmeSboOiJWlvA1fqfNoKLm/bQ84SpgNHfhIufBhWbcGqyFAJrAyUeguWgE20/+s
hmb27MRbxWUaC8mIrG4OShegtD5hC2ye69S9uKCIYWVSjXk86F+sRX8lHqjR4T0l
RmcIexQjSeBsulqZ+ZR0Dh06ssRlHf/NROP8yQfIh7UAvxv8qbnAWbjL6dA/YA6y
uajsw2rn6FsQpTeHCvaArSw7/dYBp98fVT88MeRbodlKx36nqYi3lxwyZIEOtwhp
gRex5XcfX4rt+qamuAykVmb3LlNzjXmYQMZdcONo9eNjSqztamITpTLt1XP5itGz
x998OSfTGmEzSqo0UAG3BlfBrgTuiqand/siPjgrTIr0P7CM/qaDX2eWkJIMhKcK
y/O3a+v2fY4DPDNYvBFzEp5/QFcHMN+zAa2rp8Ch5wrsRNOGLoDgpETFAi9j//60
TVJDFBrHeNzASSpMKZ/SMvYHXplrborxrToJtotukXwULG+ULbBHBVu2b+w8iGcz
lf7WC9tw84fGz3vhz22qVgJUrWz30f7ivnwr8avAijZ5vt1X/oMPE6qZNpht/Iwl
N7TAZsfZYgRKoh+H/YFE7gaF/3szfKnmZX/Rioa+GVR7Y4be72/xXnBtZMU6sYYn
CzCTvVknQcOh+w3ypA5dquPnlFehDfT9UYFNiqeJMILn6wuAs9UvjBNk5cS/HawO
5igByfDK40tO+hoKFFJHWI8LK+zM+y+QfjAfKzUYgO6YzvYlgpDf65WWMc5da2dl
08att4BzbVObxISFwjGDvhY9c9T8zEq9ZBFrYfg735qdGD+me59Cal0PLj4F4FSR
9lj8l1ZRDhMJrOcaZ3VL7kfHVe8/EommS3BQQCq+mBN/5Z7NpECHnVms8MckAQEs
EELeh2wLPEV93m7DXHzGTNTmC51Bw+YrMteeKIfCVfMj6haDAD7rSVzZKh1tSMyy
6LO4GQeHP3KeR3WeWdZXGAT8xtjze1BxHIH0Hb6qcWQ1X5K/XA6bz8+6bvKZV4kS
DJ5dkKaGzkz0pJIz50ZHVoYy6Y0xZEJG57AgsuYNT9+lC2un196TZzVDdnpFn2GI
46IJ4AnZ9uTKXLd/6kuRoE/8FR8wDiPwI824mnve1Q4hzbDzmafnS4p3We7RWe5v
E699DSraaylnLGAo+ltc5i19HsDdRbpMMFP13o2cJFn6LwiviQ8WI4gQLbc3+25F
Kcr0GdGF0U8WjXH6CSJ8c8OmVcEWxUKchMMnGXhuiK7x9V/hcxrxl8COQ9bNMm70
TXMS0MvAdhXZv0m+JKcPhJjGLeWKDY2B8KVP1WocuOPBBtErCeiTDRYkPJI5cd98
zQt2TSt0R3dDQuo767HdeCxCT33/mbL6H7qCJTeBu2XWw35yMftsgADoXH5Ua3lR
C40OXN7OpMV2zVPPDxvUEjAhzLqS8E3vuPv9LKnavNFe1yG8nKlPwa5i1LyckSVq
SVh9y7zTPSUjbBOsKmZeLENgfpCJm9WQf8qJ2+nV9WAGB7kK61Ao+xmH63V7rbZA
c/kNkHHIwqg7e9UwH6zHXK/SDh62gI4Zi5OmM/uo2u8l8FP5PrTDdQDVOiRgomq/
kCl+ybaH8kQxq+vFP7dYpCMN+hbfZ59pP0H+YswhwmHyvcDZ8Nlqhdu87q6nACcR
MtDFmyNj/Khq2QUrs6hC6UVkzrPVIPFbI5vBcZaLReCe3HHfxjRZHZigGWxuKGIa
2b8oX0NO9q6G/l2oQucQA+Rgi8bb6Qp2pmSku84VhE908JmPWpfxOVEWQaeWa+BZ
vdBjzUV2T2Lcnos449A/QVQO4i2DhCurqmnJ/DNbAWLPcaHJqC5D4bNCfaaoiACB
gms/rDXf4QWpM/03lAop7Mt0ClcaHLFw9MZadG8+P33GiVcrPqKrTnxYuv8bEZIf
YtJyJ70Ra9qlH++CRN8CVmlOpieVLHBDMcFSyuOCM+z/1kK1CV/qOgwucyaA/9pg
hrxUlYZmHX/8n3XIvSpV0+YkqRN3tFwxw7RJE0tD3H8y/AlE5Wo+mKM/0ru6FlFU
eQIRvg3ORoIA3tmCiJhUXgRz+xs3VNNbyFW5LT6Uhd/GxPhUso5K/IuyR5pdMPu3
R6+2eB/psniYycHo3NjphFqE+kN5KaQc0q9W/dQZ2eNnAClFW/HVfKCFye8rXaPl
5vIkbrL7bsHAFGkm638Xn5IU7L/w90MtvaPQVQYzk9+1ev8cH9a5WnpCtvYg36CE
aYVGzMIJ51CqtyZZBP/1UaiGx1t/C8Wr6C/vtYBXmewFuaEbJ9/myzTPiAh9NgBt
Imwql1rDZme3pygSfSyjqv8lUbBEZdh7XfodzIOMefickFFG70EQDgb5OvA7z04t
WWcYltag5l9dOEdaUTEqQ/QRfu7RP6aRPM4AsikFa03IJsLaoKXeqpzhm57onm98
xKdAQ4ZjHYwnkJFP5nGifnCqvIacOvIKquXd36vv7uL71LijjxKv3men9wJYXDI+
7LGQ8fBqqcX9Hh9yHDkVy+KJ0zOyHCQzjbnreqfOhm9Ll8isZGrW52YhYt9csOdO
yh2odwZkV2TbHwg7XCLoyQveIsX6mFFwCTMUDkFpBWsVQ/jH6zugX5E2N0E+Gitp
Y9Sm5OH2xIBpkyg7Qe2sYqeB3FSWopslwzXD2+GZEAXNnpHMO4keyHGbO9rKeq4D
vt6emEHbZVHzDJkb7f2z/2WaePE0PTo3I9J3Q3lN/03rB2YblJ+YN81OPghn3rQV
qroFbenlE+mVF1c5o+bQPXpUuf7lU2wu1A0kzKkM0mp5Fm9Lt2MyDlLjHkgpV+Bc
QJeqPCJORRa+X00qzSKfYrfSW8cDpFKyCajYrlir28xc1vsc8QMPZFkCZgOwlkW3
UZJnPm5k5WUvWm0qqBFxXE7M3Ha2tzOGc6s1ZVE04cJoaKUK8MMMb4gvqBjMMk1+
tnYmnJx2IE2zeP7yaUBmOxZ9/rrDRijQOSXyl9z7y5ocTcKgOxWUf5EHXfNXeikQ
7DNmvQi7hFvh+3A6nCEILAJms/5PCNdXNfw/btUaGYYEmda52/HvOCg+IZreUmSr
XMm5VfDaTnP0JZgbu2DlnEd63EfvOQfUbjlEFmMLUkJI6XbBDgoIYolo4VT+DuS+
1VyDuAMAxuerPDURlcdQoSllnv2XG/iBKV3q7cXYUj2xoUr0GUbZ8WE9pWe1v/Y7
Sdq/k9+BIlWVvx/IDrQbYOmbkIEOCXCQOE6kc1MinjiGq7LM3v67QgzjO2+njwsz
jUc/Q5aSxKGYuEnGv95q2xmlimB0jZN9mQS15BfVFKCPpIQMA15fYNEFJG93suhZ
wpLajPiFARx9+vkHZhKa8okYJBTeL7oV5ON39itPIRkFVWKyVYJI+zcGYzdSCTIJ
sFdf6Gp3y9mo9tNKH+GG/OPNnEn5d/c5bLuyUpE66wd455hXgC8ejjZDjrmTYFQI
8X6qVhHfPCtp3iZCtzJPpdzNxJQaVyYqUya6S5G26r3eT6Z78IDyavhgXfHwI54M
kLOzvnGQbp8ZAzSc8yNSLOwcWFLvOyA8cHKZJJ4FeErPx/LWPrkaFZcK99vjOHGZ
kdW6EOm8Ydzmyc8dML45N9ZRnCLD5GG6hQ54MlxCoo0tRIUnnONIrvRSHRxMQsFG
ciOgv9YRoBSCuC2ci9/7+W+J8/BavAkNFKw9eWgyXqFisuW94bXe3qgclD51aYUm
7ZlGWBB0PXyb5tT9oYezAOb/EGADWBRswxvGa07Ccq09yXkuXcTsRDtDZXmLEyQw
RnezDd41GFCN2WshwzvPDiCSAX/bYl3gfTxpWLdPyH1WqYGDG2t9sBZxSvb9bqlm
ExkKR2gfkYuJXZk/XqZmDySdwDGKu3+zEs4bbIdgz8TJzZlNt2UPemF1ItmWOBbl
PbCCu9bZkloHLOXq8RMQYrMPWc1hScwdbD39GqqqCyKR1gXgYn9/4ysgnjoKe72V
6AV1Xt2SrmUbKgd6JW4/5mC5+W2/+gtXV1p9CIwfNwrPCL9uhohdkmmHsIZh4eje
SUO7nsBWlqB7MfoTJGa6MhPutNkEVMclh/Or7vVC90fmsttzb2WruSmmvF/O7us+
BgKXcAymSI0iCd+C0TbbN5qKVZOHh9M1GYIplAcvrX1klDUY6SUkmdZlh6BS7GPr
ZZPZxkZfzwEHAnQAGPpyIPKudNmXWNBhh3Bi3ciQQigDLcvpEhdH6Lp9GNIvRHRT
BG0r+IomNJh/mxm0d8Uz6muVSyyVgJCZNSqDg7wMGMWXLCgvMqHZgoxLqf8Wh7W8
+QzLcu2bCIESY/4EYI+VpqbOBNPO0ykWqCU+Et49LvMyirCDD9J17ts/xqtfhk1B
0pwDv5GMTtfG5aZIQ1rcPPcROYzIvWUKKgdL69Mn6GUFnAfRui0I1c9ptZ1Y8Pl0
IPqGa2uhkCenrYmfQc3vIwXj5jdftEGkPcY58+lQCD98ScjnENPbnesBS+efb+Wl
etaMcvdHTuidC++ZjWUCr4FMk4mbrrcOla/DwYQkQNOs2c9OKHetfeqGYUE4usP+
PCgy7yqFZs5IOVGPBD/tDSx3wmWQnU1DLpYTIf/AP/HqPo0oqUj+rfT2kPMpQx8E
3KKoGg0W6/J1NXmaopQDZ0vxWb7X8XcSunnPRdBFKpOlLTqilpw4zmK/8Vo7eqlK
JoRgUZHfa128lIQgACHHa6Zb+iaht0wilgrFuG7+UQJ0iPLTL7jBpbQ9J5Wp7EuW
q6R4wpK/4us8b6th9iDkQSwc/P14HzQay5mGp53rxJMvaXsuXBzakp0pQTEadG01
24RQi4zqd/Res8S5yxmj5g1MDLUsMeL/zQ6A7vqOdaR3gQ+bM9kO8ezESjpaNUBu
wSag3SEoiJus7FcOUFoRCRJIFYmwK10WkmOBtEsWitxvA61sXXrUvusT35g5RQHq
fvdV6B+wGYvNqemqinvIZMQK5TFkzbDiHiUlW5+GNAai+pDkPHh/r+IHLE4pazu+
GDbRdQS/ibNkIgBig53sRiAcy+yC8B8yXLLQDlZVG+H66yoSqn6T/W1HT4egVPDY
1bJIoK/k9qF9VEiVgrFRUuO+21sl+Oknq2a2Qt0C1QLG1T7BWXeR/3plECnYFgfA
U8WgPfX+dIcFy7Rpnt9ick03qGTYcGWpZZ/EdHbLSZYq+zvDIBVw5N3m6jMDa3h+
ottkTaln2Acb2IJ1p6S4RDJ1L7HTIAV1V72I0mqjRi3dtc3SAQZ60qYG+IkU+KCa
u9ztWyX/QKMmK3p1mNDJLcGoKrF07KsZe1PFjL0qcGus2T1LDAIM8KNJ0oNRKCR7
snqp1kzIev6m5n/xgMBnWqJ+/tM+UBJNJgkncOI++FVQA+e7Oz4AQFjylUagE435
hfDzAMCqq0H1Z9+FE20Tv923hiPZebmhza6+uvSAWdBVPNF20GwkcFvZJ8u3N41x
YHMOafK3y5SqwSaBSIlLakBFegAnvkMv4eu760ze8gzRd8ZLdm7DzZTe/MDSXnOD
qHs9i8qHN8uiNB0lsbOgv9nyWFH128uqP2A3bZ/BaYnxnQMTP/ZwOQVw9tj7EO+X
YVxtrbqzwI7tIUR9AuRRgcZbDwKyoGmbNnm9Muk2lt/09kwVarHW/R8HvdQ9vwcv
Yuy1rFCZZQZ+ERzQa6Xv3LeIsIC1PDgOoZqlRRxRHFV0/mqp4gMpJon8CoK3YON7
JXSklU6iowDH/5b7TqzmIX15IIS2We+EjRU0yU93/NkwOy++RXgfuQVyyk0REH2H
J061Wcj2CqUooaHcrWPHX40GZmyR+Ez1ot6GHplUidbPztvh/zXhddGZ74K6Km8y
rG5tfKDjss5fpMSkXuxu+q+d+ARiLGZU3K4pzmoCNB9d6eFs23xpZHa+ljkt6QWY
ph7gMEWxTAppd5D7MpmAu64eDaHIALHb8ka20P7D+un4ggd3fkrCrq8HImrKl1Jz
RuD0Y8J8WSE++xOIh/fhIYJqN5yGdDrpGqBYiGvZd73WK0rniCXT/1o8fQiE/TAI
dQ92Ils0wM0JmIy0wMOJvbCzu0XMyWBtZ4bKuTkV+c2+kkNHhNBYrY7fZR1apSg9
nSrfnZ4P0utnjYdc9nOrtk1Lsop5St2zkcWuF0CFZt7BlLujZ7P861Xte1/4eA2V
S6BTRLFnhuYEp+jiKQWhY4g18xNloRk8G576TSZgvOTvnuG4SB6eZO6yUJ4kYVi8
oOXWPoGvcaESCiCAIDhw2AuzbEu3v9KhaFD62E+b2AyWZQR0Ag6QLh3NogzmtZ/7
ComkQoGbgGide5WF3LMNMtR71tNFxl0P/ZV3s+369AkRJCYu/qdi8uApGkkE5b8j
TpeftGkZCa+yHOWoeQBLOKtBcsGH+S51vG6R51MuIgk5qlfuxM0zbEMNeAT2crx9
Q63AjFn//30PLWjpo4QSnBoIZq6EXlI0yQTTRowqyxcsKb1eFf0sEqo4oirgucqm
H0vKvpSV8p1Aa74iwL5y+ktsTgNoQyTPjB3p4fkEF6+tR76gSY4sRiH26gzC+aUy
xxSre7hC4PXV+DELZoIBHUK/j0YVFPVgb7B/fQfz6USHUWoAlODpH63gF6FaFjNM
omz+kVmQIsomFFhQf8KDSv48173S/steUfV27C0TP4wzVkeSXDGM9yFP+gO5nF5V
7XF4JuYQsfCc3dztlrdkCHhPrDf2QxkfXW3wOUmzzuKNJ4V9W+8xOFd2Yp89jsn9
2aPBhq76Pbicb+OVnIjgmaTSt8qq4jVUeGgLjB4lYGzUzqeGqPqJg1CpghBlFRW1
dmSazyUWrFR/9BXxXcrz2MeP7vQd0r0kn1qbKjj/uhVgkaHWwr1aSp899UWBTT5C
0gb5CA5eAVM0ui9JFZc5Qjfv2VdiaLUTQJq2q036i5UN6tbH90cNe6RZ6TIUBpwv
x9Oe/zUDB8XInA47kRxUvNPN1XFQAyvuTQcDO8QTzm6UHeODEJSpC6Sl52Q2flqq
CIifjaGrr4QeRvt2ohr0dXG9hZSUXU/mDhXKWYyPstoVt+jaVNq9BIJ5MnrfSLea
kIrTMu5Q1EcGWFrBkGO+oHV/Ic1N8YyhhxY39GMi5FRDr9DdZkPLp3X6kZ96ou9a
laVIQRJ3ah0FQ5Zp5WoTe/DPe7ZaD8s1KJ6YIh+edTPWq0sjhu/7Kmeg9eSaCxFy
snr72cj+Ug402u71Ag/HqAWU0i8VWLQnrjTVVnfGUefCZVG8t1hwof5GFkmmogSw
XCaZ3kPmyc+gr1I2zkuHUq26FEjfdqNugPGTCcyXfjET8kTjRYeGXu6c8Ka3R2GY
6rykXb1YUKtNAFAFGA4NvECL4JSqZMEMDkQTlr0nRt20+esITt0sLZj4dC2d8Tp0
fNqTAEeBnru78dBMo3qWiiVZDHv/OzV1YgmDuci+F5LOYZZYj0FefHS5SfQPO0ep
Khd5l8zdpilx4yF/y7phYugflm/NctqpRZgFS5RTerZ4EYoRz45F34SZ5kAn96HK
Ei+PCP1O9JNNHl1a8CL4PdkapC5yFMeSLGqNjpanblrjoKRNetNabp5Z6/FZmkEx
PBQSEdKVIvPRafQd6LfAZ9jK2yX5GPoXxF0FIBKC4oUhC29tW3cZuwVzmDYvhnzx
0+e2cn5kwUDUDYT+5hnoQ/WqQ5XjKVtZf4L0WXl2hR24DADvzdsH76nC8Jt8FRpV
CGevnOqN5iOlZNYr6P5by10/JveqSPc2nhKNk2aFPUdsOvYAo6qD5Oxi8z+lWqmd
WCzVRyRiYiT3W9kZrs38kFt+RpQfSBshS9Mq0Yd6tEKmJ4fb2AxbVq3yP5yqx2NN
XU76REmtH+r+1vWKcOwlXeCFHPlVCIVBej5LVd+wcWyMIvLvKlz5Thoa5JvbWp/i
MKkU02lyK+xCRP9pSeTahdd2mBOwiZIFgojAuNA7ImMf+wRYj10FtScAUwPzEXTD
t2foOoaJTSxFoM+BsjWj0fhiANWFXvLqBjU3xkxcTOFgtigbowMzHUUySWo4BTsU
UGfT4ftjiHH8HC6w9X39r/1B//HZZrCuODA+JWNXWwcb62aHtmN/NmuRdyuNRjl1
2wc5v7vTdCYUwwk+ZctSNncKVk8AKL9u0f8amWffLJpksA8PyQkmubrpIu1RmAFU
HXTXGukHwkTltgS5i0Iytb8dH2Vhk4MFDAXXO5T/8xyru4ygzFuJrR3bgFhPkXty
b6tpV2YGq9Jz7rPkkfVbVJ0la7kWT0um+pk0jWQONFyRB/uLsicsmHAS7wnak4VE
EKvcxSK+GGljJ8Gi3ohNh1tZm6T/ZqDXwDr5WRECxBcnecjBDQbN1GlJ7js2eNWe
HTjzH6EDuxPUH7N1w1Zd/cszgmprWCDbXo4tatvsPrLUi7K8h7xEf0e9t7QV8WFh
gjdE0c7sickTHabsJG2r3T2dUgFqWV0o8Oauzl+XraFGGkyOzOfMeeu9Nzix40sJ
F/I4beX6A90AZD4Q/FyCcNubGAywa9dH9WS2i8uzmKm0NpA6OLOw1pLX3WclnO3i
dkNgXP89mwd8Sx/h/g81ym6p26WPJ+grl+gYV8Xn1wUSFUDS6lONJ+WJReUi+eFP
PRi3SPB0hzarsxW6JokTVH5GXzAv/6iuwds2ufGvIFx3rQCmuCDU5PR1IrdDIpr7
UVsTDZt7T08TopQUj3TM+r7jBtRcwt4skRK9H4YpKSeUXyPhYCRukvxXP7fepKkg
zaYX/jZj416maUlWIW0No2t7u0lr8wSglm7Q4tMfkV4EeR0BPd92nxHirBH19DE4
qM3B0luzqRgofCi9R7qescdqlmRniwIyQ/gGvX51jmHZHj0CQbG0afKP2mLZBTNW
Le7tP3FltPfAVV3i81bh7YYU6Ki5/cRZxujPcCrnnz1G8npO1rZ1W+FbXN1MJtu9
AKbrt9sH77D9STCWv3v/VJV01VTf2UEnJySrF2d8QQYZS08IUTQm6Z71kYaXQt+v
pUZbXBc5HC5uRAvk36sr5WOY8DJUhHTl3iW79aY00qUUqsfGP4CKjzaXMoVOtaTZ
853WY5qAmeMTaxAJ3xt3JQhuhkQfPr5s1I5E66vsuLYdFZeQ3R0GMMKPjqQzr+yo
9OlbNnkBCigsukbIqfNAMnoeLfdYJTpLJeOVIRvQ6rNp1wWplCPjDKhbmb9jL0ti
dOMBWgjVguTEyFkSdUCZZWiF48hzY5QXIQBFekZRQcOIjiT1SVs6NwXO4T3+Juab
LCjt0ojLES2kgXpW+KzOtrfG3imzwizDPw9mcqti24IDVeIXPdWfd+kdfDnGXhoh
T0AGkFcxUgo+/LMw5U85fJEg2pisi1Ehcf2VnN00rhBRBFt1dGZZtA2C9guu21fB
cB8MswdszMh2ND6m6MvkcpLkmlWwBSww3Q6/rJ24YSvMjG744x7zQVKSet/fHYsd
CeDBK5z7tmFJm3Y/bNfMeJ9lnsaf54/xarj++DQ+G2K7cNStUKqVweYwQP6r98bb
zNgypxjk8ErLkNMXeQaAEfSgvgyP7y4VAH3VGNzM65kSSDdn8AZfnrzhCOjifFY7
Dxq+5Kni9KaTFepqMrBJk49uwdKtWicdKo1TgbX5Jp43ZP4bTTOfOafYVzPGkrQW
CK7HCBbTXJev1bR15wAEt/UTDbkbzm9LWPtko8yhOkyAGpkDM2VSDooRGUzvSdZl
2fWXsO/Hbl0VT0eJdIJ/FFnLrndd8ZlXczpJKuWjowF7ICg90DsqZOi5Z/RmauvY
V4v3aV093GgesqmaaPe5mHi5TURu14zmKiKwTQuWfrMMIgUUf6ldCJ1UUcr6Zd9E
nsi4fOLuHxEiBnDI/QMVrKEoQcZQTWoPzbVqog6RV9+c0KtK3NNM3eY299UykXN3
1i+QvaF2hu+RUGAEEWw2ir2GGgHcUC09tfQ9r/bWDL0q99IO79ZtBPzAHP5FpC9N
eCqyLF1acafzVgTuJGMUkjxGgd3RXYKQiZkSWmD+Kzjb9XyLT83KDoj1nOyr6Tme
S4MTNs3a0ADwM85DqFYPCNFs8a1aVMvBLwMQC6K1nNnPidM42uwOLQUrcQn/PXPZ
iOKx9nhZ+t9cXq5423rTdZl00UAAOfaeRBbWmdh+CZ4mXuyngFOgBf6oiSdeDKMR
IbvvQcwqEMtb2x7MU/B2zQNy7Q6rl0gISWB06Jwpr37YDVt1c5iLK5yO45Si2hW5
j24YM28H3bTca1BwRIjzPJrR0Zop81OVcqOU4/r6PJbYnhAj5Iuzg2kPf28Xu5z5
j/K+Z+ZFajsnE8fP/c6POWB2zwdBWAshQM+kdwMrLtD1eYMukqKv8GTS3TSUq3ru
er8P0CyVhXgGZBOqW+t3D5Ec++mmNh/+00/huK3OUN9dAV4iV3uUxY2EHHY4mrmk
Il/RMmHfksUEBdWDhrqyP6nSPrsxMnJDu3UikbkDLONUapfMJ5jKVx70pBwqdgoB
OpI2W90zDa7pKBSb+J7FMxOvWfd1+efZ/fg5jxxYbSkoq7cIZ2P+652uyXKTQGbB
LuhUy829owV+aAFeBcZBhUV5X9zDHO81RDzKqprujpGl3AaPzI6RT5g1hC1woVfM
4irmqkT2Awiu7PTPmW5ZzprO/O7d0bjx92XsMCC+tITYnKx8Q8pVuw7b0Kz7t/+i
9SkpYQdEsp65XlpTKbZTbo2Tg9oYEak+jA0qJ20Q/53ZKnGDLaYyoNJKsEsaXznA
T3mTyAlrBh7KTqkoEim0C8qlkhQ9ZHXG70Py7d1Cq5z89MgxB1xtEwtFzTV+p48Y
4KmYIJtAIC3tAkh7+YTsoQUSJITnaa+eLFiKx0pKecpdAW7ILwrsWMtLeEq7vjr3
Ung9cG7z1prByEKWbCRqTpiePnqKbZ7zxeWjTus/flKD7pyc8ZIFwDGUc0dtV03I
vw5ypraP5BzJrf1/SRxyVzWILIJRD54PAKRcIZ0VOwg9qeqgy8A/beywFQWGjPRW
7rPi6Mkhwk0jzmjmfK/IHxe0QuNvTtvvHAEPYAGhaSkekLnMSxAOdn8AZnuFFLZf
fW8OBrx2xCWIGn+UNwZHmKYS43Rd23LVBTnrrX8g3fDMrI2s/SUam92hsnDuUyN4
XxwIaUPJ1FnW0OdDM8mFBKl02uFbVITpR4a7vy7nd4GeLy8jhZiRExbh2ju2H2tv
vkhPtSYSCrYiuvNOIKV98Po9g6vNayDdqxxZ7stdUhRO1Sidot0UgLvLNXhpa86+
kcPHE3kvNo2kcioC5qELH0RoWRMNwIdIlZc4gMbvhEPMhcUijrgwBdm++mOL1mHp
o3dC8uhhlMbiXjooN20UvEuRAocx2KJddNuE+ZrQcCXG2hV4rYIvbQvbMRxLBIOU
ky/MTMp2W2GZuMPbmbpQ0BIwhQkLBx52u/M2ZnkmWem2+IZuntt/phX7s2c6cnRI
JBTNVeC4by634TUoU/ZSqo4so4nTatTA1EAAeituJVEFjs4pH7gTz9t3arwnnFmv
CMjCp46TvlTC7ZimbvegFa9dUEP6XXhbJ/Na1VG94AFkaYFJiavh5JkI2YsZbzDt
Q9zBlbCpKtQLA6RzJtdnTdchKP9vObi5m/U6+vOnjY4oHzqvL9VpNy0s6zXlmw0E
S/kdk3/adUNi+IVLF4d7S8ZPHT/px0bUQPdZ6VrdsqSPYSbnp0jEznH6tBCzkSJp
t4iQvXSkZFRE+Z0RGehH0vCAa428f9Zn0ohE5VS/qbkpEj7B45Jso4GyUzAyeMqk
4gwXCQWoPjoAZ+pwBnkzovdmpSDlumfcg6ciX71cRY9z1gh/Q2cG3aAegaBbcukh
/w9RwH/tnDm17CFz3/Ua/KNdqyPljHPyQwE3NKbc3rccvTQyuG99I7xvVCVFTaJ3
6mx1ZBa45Gy5ZBKteDVfw8bo2JjMRr2ti4D0MikhDBRexgAphargBO5aeXGeQ6jc
nxKtg43/J0ULFt5v+lKa2aW8EynHxf58gQsYk6C+hRUsQ2y3MUe8uXwD2STswzIG
5RZKqcuQ42tr3bayxBw78SZ+twkOzyZl43YVAvZpKU0wd3qatWlcSyG2ZkcwGo7A
JVTc6L40+yv3ERVDDWSWzmkPA9wZnWJOo74BVtV8BfIcaefNzHp6xSDomrFvTLjn
RjsL0RyE4EVcsv/zq9CitOViXzOZTxxYjin53FHiSgR1YV59lTzpy/wrc7C46aLg
a27hVjdMLXXLGxnb9pHVIxfRq2wcias21qCsQGh8NHJ1miu9IQyE12jz+TlO9Wps
MQBGMrPgg9fExjgdA3X7TllIngOWHYfm6MscO/Y5ZH+dSIXuSzvQSfK4wPuU4CkS
JRbkP3Rf5PGURa6ltSAbd/XoRbenHg1ed/XbM/eTylD1Qk4FvtgifBhX4SZ9oDOF
2jUNV/HLxrj41srwrmSmKFJsIxEcEH+q/DjupzSVg/75LBYSdRkcQLY7Ne0COwrn
6reo9a4PTo2sJBZ+K5LeMML9QT5Cl/JdFujybjW8eAvHLirCq96GI4Xc53B44Tk6
6PX36Q/BE1+wsmi2VF2TlhsF5N2aLa8ZncVXyKdCD8gL6RflCFCAn04Q0DYP/7cc
qWozRbIUtYU80npXTSsaZafD4eBEgZmBn5BrS3ft3XhNVlOV2ovBEMFy1bdCAsS1
Kts/tTiHtG+4Bu/AdkhrbRPhM0Y+tQXPPv1T0iyPSEPg/j7VZSRVlb0k/wO1VXjY
h6aR/BKaIcnaQOLIwuHSBfde8eyDqguGh0WsUnfMi87YS7MOX77hPPbuoO68I52Z
kyn6lDvhmUIWjGF7xOfHJ2JUKC9Wh/0K7orivs99R1M6OIoFa1g5IkxxMOsGllmu
djZPM+w1UybjeWl3KPD0v+5A+65B9JyruX43zjfhzh6HRFfaHt7X7P1UfoDeT8l9
6JGN/0tuwT3Bvlri0EFslVhXGKPDUBAsQxo0Gis7DHl+3oUjjcKWEqYKuzay6fcR
bcGjH/AQ7QBzS9js6JvRRLf3hvkXbgrRdx8qqe4epBZNbYQGDZ3txxhmLW+/Xp1p
GF/XPLmYNzNJlBj02vfd857vqgBAjpnLWsjnakvORuyZra7zQWvgt9QOOZIHrRXC
47lR8BcQ02NanvPTl36BHLxyK0DcmsjNuzRaAZPFbhLuyAhhuKEJoSR5M/iZORBg
uVsl7Bys/Nw4Jx5Auxzp/rbK/SzNAK2MHFzRj90tc9cbXKC9swTQGnmJbLQItWQl
DZYP+xSZTiKwQRZcNdQ8UvFr9AdfyCwmfK7e4NQSRVIDoCRVdDVB3BUmI7V+H+O0
Ea0/pbWg13wSvMk5FCHUByG7KI7MPbX0aNuZVA6Di75uJ1EL136s3qcCqcmMVhAi
7p0bgFQPOPPsYkBeHa7TE5WTYLZ3JF/ZcWH3DO1C5JH66d+yRCJ8reTG5NfJgVUZ
Je4nbVtPMgsbV4HgazCNCXqWrtcantVZCiZMnluyYqL42p4ho9GHUEqnam/i9lE1
CtRsebAnLN7DpbDfQ1Z+I2U2TrxdAFt4Knma5TBuHDs8fLhxv9tco6zxA/Qpp58+
c7q3aj0UZLdYXvO9IjN21PtjWkft3ZiMUVW2S+XPi1qWQ6SpyICtFxVNI0c8DTRG
Ux0f5kXfWhlF0xUAGdg6ZJQP8eJC9CpNTz/8iLdukdPY/Ae3jSXRui4frWMkEgly
lKo/8tDWjeLgjK9+bfV3VB2Ct/s5kOrnoSFIsnonl9QZCLQFk9HIDiD4OX5dzuRm
BaDG9xyBh5rtKM3Uhuj1qIIMmPstubCi7dD8bcj5+g8huB3MJXtCJSw/9gyFx9dX
IxpPOWGBcdgoT1HTfKbnMVWGNDbyaqHx/VuPxnycpBM7jyqFDakfmhFvJGwl4+js
UUzJWd8dembUugmTmT2e+xNzOclDebxcHheBex3d6KIna0e86Ck9gwFa1IX45hb/
C9++C+q57yekKY7IU7oZ7klnChtiQd89KPmE3wVDtFFVGEAoquKwv6IUr3FNvkcz
p/bLZwmLKueNkvg0nBXu7Hm3E7N/rUxqCAh9WxAopSXeoluYT0ciNmbVlw2DyKuL
7p1JFJSH6B9TW2c9Dc9PA4JPE/EHWH+7G4feVxJnVamlDeBvaPr7Y2VhLjFOZ2nh
/a6BDF5o0QzUvT9HQr1BeqjRK7eG1q7Mzwz3uiwBcfAUIPcPjdSGP+N0H7HwTyKn
3VSLRS+hgnM0xq2epIT8iow697WBDYCmIk+ENkkQlZ5sdEiDjj7ovdQJEJvxJgKL
+xJBx/2fylvUcWHHz1HCj87zpg9bdFlplOfRyIypS6h51snMtj6EThjf5sPZ98m5
i3Mk+EI6CULEIRGccX+olIUuJ58PouPJEJWwasGqU+N+dDYl88+znyZX6Hr95Hwx
dKk0oDXWFLCJCuSVOwdAU6dN4UI2sVCjhObThrdxHzZ9i3w+UMJ5FHX2ylYyh5TV
uz1pXIoz/e2fUHymucF1HvKyCoTC2pRS5uAQaseisuP9cYM05Yejtf07I3WeUJx+
GOKMADnuPY2oKSjBUpOIdyEuZ6LGqYoVT87viU+e1xrou2xUwqS+wFEJZgj5xag6
q+9Z53O7nkSXytX+aL9PwIaLFDPi6xhFFdKoXoY/zddWYqSg8PkPXcupjLfY0E3d
00cporio6Zn3+sfkY1GUZbjNau7BMGpWzIoe8cf2+c2twEufVznS7dz52kKT90T1
ZNxylS/of4EvOm9wMG03awwXtt4aikc0OpsCa1Pon5S2W4BE9GSDdjVgUwAlhAct
UDScimJjT0JcuJcTOSVl7Em8Ke1xkhgUN5pB4aBr9ABCdCtvbyKnZ8G1jVGVtMS+
ZQmxGsqS0IQixZfQpHkwjXL6C5StU5fKuMrYhiZlvQnwcYyrd+wjydptXWkdt0g7
CC9iS58+rFM6y0ADS/IMdDUbPPKfB4/pZvnPDMLCouQ++cytI0M5Qg50/mLIuT7L
GJufh+HH9UWMQGl5+QNWR8R3eT0Ln3BKI3i8Pm2jqoS8AbPMOeUo9b2m9Iy4aIcX
H8wTB9l8cH9PmjZKJf2Gq4hYJ3dTA2YGWz8e6Ecivo+2kuxKCIhBbZtBTaXVTpUD
3i5VJUNeZ1OYVJuamEwpF06pXmRjENstLV88r4hC4GjdCiQjSyFQ7Cg8vlkhkV/u
kKmw4bWtaTFldslfQzBKpiPyF673Pkg4ng7ng6fth2HLswNsa523pOVA9L+KhzaI
aNKwhiicOCBpdF7zBehxmfKZAuiO+Zlntuy7w4aiPSlTSP5NTYHXOm9WnOct+CbU
9GgVX/7qJavz1W3vovi3YerrLQ5ucGBWB5EzRx8OH4kdfRlKAtyE+X9QLo9NwFl5
wlHH84Efvb5MSClQTRvAVhBNhOB4R03NNHCFISXQFVFA/gRhytnuw/noNcxjFsIy
x27CCvr6Fo/mc6wbEiEvRqkghFMY4JPVFlWxKK94WcYeELKhgxuH7LtclBpuowpP
zLntuRFem6t+PY4zXa/zNOXaTUD+iz6RQHbKBR4n3zoz0uKy5SnLoT7sPWhmDIpk
nYXu52i0REiUavQZCn9Al9VB/Fj8NlrASvSup3NMICnUizlnSBqAGHSdiSigOuYa
NyiYyZuJSHlLnhJvdQZ1AF6EfAQ9y873PWDDatqpMZMo0Sur+2duzs+7U0kqchDU
sZRIxb/dyZCH3MrbSBxW313CgozMJom5yA37PdbHqYoPOS8cEj87u3VmmjHyZnPz
/zm2b7ffrA4aPX9SngGyZP5aEK1xc5r0KgtROCRYdCveNFOuNhOHhJc/Zv+VkqVG
IAxPt6DLWYVCxcse/WPapsjU63tG9WD4uzP1g4UMj2lJdzXRtWpuwFaBS5A6Nj+h
EgP1jFiLG2ohc9GfsnGldya9/uJu09+/RSlifpHHkrRCP7qLyI8b5MrAubkCM1FY
NE0LYrq00aTA8t5aa8UEdRttIdiPqsp5clfeFUqn+zv9J21wJwjUuMe7oGqDFCI7
HitTut2cw76k8OYQbAX8N3Wg+6wwK1/WauzV/VC+RlFmR0KCPzoCC8Nt/zrZK59Y
zBjKATQ0CaUOILnz0kPiUiLqllPn5Z73MOdMFiLbeMOSFJpnItxMvUOGwpVxLoIS
mYfAzwO5UQTEaHpdNsK6wISZAGxYWpqCEOqmeMFmyEvV/gC+ocAjZ9Z5HWWjg7g0
jNdj1AmXjSg4kiX0tE0PirxTqir4CjfbAsjqag0ckBvWb1tFlr+HbxXGMF2P1U0P
yYb/nE9CjnQXAACfT/t68ZHdlGLof64Svf61JDOg6gd922b3LlxLmYzTYXLbTqgI
Syb6TWcSQ2c9MxWEcu+dEpyoLbHgXa9hcA0JY89Rvwaph7wW2VjEAFn9pjwEKHIB
5a/kh9SBUgAUHT2RyMtQVtP+992d9H5fYfH+4QUDVDOferXi2YayQ/1kO1w38oiT
qezDOGZCd7/2TQhCDsoh2eU86PZnZExgOpTMqHtaqCIr/A8YfqcNEiggeaDUNYWo
aqBTuoz6yKLUe6bNpE+Wj6/I0GEQAin3Y64gWi/5Noy3eiGFaRy3Fqpi67Qc38xl
QHSlRHw09dgUDYJxDrBOc7+8zLvcSM9slVjOUaVO+JBFLsMkp27WRTdkRIMWXzRt
b3L3Xw3OtIN7UyFWGmqhLS8CbhVcDmNkHVc2OFSITuW+OEeCjeqkcbM+E2tNRNXq
gT8l/X8+SrM8EQlm1WNC/2oobGtYSLidnUnNKdUS7nBhaVwK3Tx4XJxDqOIX3IvW
HQD4Shx1ujNLuIDSu/jTI9REy9R2E9LSdy1ZIOp8ms1BcfdJtvq+p6l1HVJtTUBr
jXSf86gDhWVnINTPVfrA64Q0sBq8XYvy1CwvbUrE8J5zHyeOb4Yd30VhlOG1G0VJ
lTh9wkR81bwolODjk2fLnGQrT2Ltn36UxfzaRKp/kKBpNfCuDpDtyFaifR3o+hsw
Y4xhLLYm0nJmA+gI6viTRbN4Wv6wTm2g+H5cDyLfs76vQ8rI2NdvFvgJ4Kw/OvRg
f4AMrNsYLI1fdK4namdBv1Mc4Ni9U6FnSdYgVk12gMeYwScp2FIakhjpr4maUooF
1iN8gN2oyChe+fSHGeUodsFiPtUsRauktudAgB3th0pFz0uthY5djZa8SZX0QdF4
cMmi4PHfOZnmMC0irZXrlzXZDkCvmoeZGRMXGNirUb1cXzUrF9kVx22CNvw1WW/f
lGvBu5FDOpP1t/Ma7RhaF9QkXKNXxQLXxjAKPcQhHS4jTRyy6IYtRETFrV5hisoM
v9NPhqO0GHdS6hiH2ADLwDj1N+oqxyThJBoELrsmQzLlSKvr1E4JfiIrdNduPQ2A
7hWX2dUigmScY5PL6khX5ZSgNmKj+igz5N/8aTpk+lhoRutADP2+SjpP6yBn5LBt
CUuKkDF6CHNRPlJLRtgempd3eFy6fOhmFzaCw6iHiNKI4a9OZ7YwLvgS2TFRSIPP
ZUR6YL2apb7kittWtHEFv5lLB/0+eD2UF3SkoaH7LhM3wG7yGd0wCB0Mp7MGZ437
5Ak1KEWD9XHBlKT22Qx0b+wr5o3pZ4cDFXcDQu1VfO/hw/fOD83GT3WsnvNFnbCE
ki+kB1ImSKUAcu5ZkZwh7+db0CPyNbk0gdyICRjewCVwSmQAUfDVjw6bOhnybWVp
Sw7aADrcAXm08/L7e+aB2d7JI/ET1TQhFrf0mi8yp6PEJw5djn3kfyT311poNgmi
XEa+u9gukEdLU21Qw16zpGtGuXLE+zlrJvDzW9buiqlS5cNy1FoYbZU/VdUBmKEo
PTruxIqrBihQZNIONorA5RGyKREDDpOqnxYuAknIFuR8LEK29RW5y9RAnx0f9B8A
YcbrVy0rvm8Wr1/F6Vp0F23P+8hdliYPs+ncn3jXCyS89XYlqk4G73PmMNOMO0Tl
wu4xWug2qm77cEwaeCWT812wtJCxk/f1x0R0DPraCIa0oW9P0uclDcdOS8VFvGiW
7geeEGX13KTrhwrBMKiA4cDq0sUdVWdwY1YiDefOjloqIXg3nfd5d+BbjekngwAZ
+/FbU3n/NhqjMIS4XgiM59dU0ZdXXghtUIy4qtchRgtmqLmNb5m5yNa5YqBpmMfn
43gqX010mnLuXyslToDidgxqFOmZQkt1WmW81c/fIXEpdg4VONgHIlioN5yvRXfe
ZXRjFhuXUoR5Abr6YO3rcvY2DfLx7fxMsEnmNv96DFPLRPZLrqTX20iA04YiT1Lf
cJz1WKz0dLr6b07DWLz+HHibHkhsgKImhWDnwm7yUaJOerxvru19lq9jvyrrmvyB
ECd9aFPiRKGaAph/pimnWHIaO4IVzakdN2S0I8b5w+UvGEyCB4+34lTvKkN6hsG7
/i5qPdCTxwnSE9acVXHaQDTfKgLDH86hVfbTLUIMappLHeBQ7a9PVwlUEagC0PIW
3UgyGul3WGGJaQXWRb1ldiuY2Ekic4Tr4I0kX9LjHgK93qWz1riXt4m4US/+zsTE
ilxSPz/G9EOoIT0gewWYH8ITeTRd8fFJoc799fNvBTHgP3aPwAkC07uyaxizUBVf
pDFNzJXN+u5CZWvIxj2PreuWcHhh18T5hPEhieKghVG8MrTejiMTIvB37nKazbi8
bAsygjmZL9snSJRWcjh19+aedoVPlzEAR93p1JgD6dLSeocQfw53OVwwYf8Gq8p/
x++cspCBmnRQ5CjCVTGX+KTCobmbs14pIBlG1cTLaUSH8AChuBJLC80gLAERNPjT
Kp9uIRqeTn2AwwKwpT+hYzCOJueIStD+AmPKB1XRK4RUPYbR7ZF/oNN153v8idfa
Cbas3IJTaWwrXSlJtvM2w/9INeVKXFfFvbEo56GoEHAX/FRTd2Qwh69OTMvn5nNu
Oi1iqZPaBpOn8+QsYDI+05tAc2zDvvbhyWXX4bR51PKivIJFWgGjiIaG1feebxAE
TKx+6yvg+dHkCMGl9GdZ/ItRUet55QnJgtrdffZUTHO84PyguHxmWWXEMIzNG4o7
U2WFqepEJ6tKwtAKdK+fSTz8+PTe7k9H9FiwtvESiADl/hqUNeomMNWQ5IqdwYAW
cbywXrkp0nX2vea7Y3OD7JnlBzubyFNXcGKj09IgmPKtJGMOuLMlT1Qq4f9ruEOR
IZEu1tEMs/lRH0GpD94y+BDC03wno2sR3uyK6QRRWemfpa5UoXeRLHB6TlcqFo6y
ZFpgyLGUdscou/+7C91TuBsYtzSPwPsFZUVu4fQfWyYV4j/RTrWzcV7kF9261/G0
6JDglmSV3TpIAKEa4zhjHoehll/HKURNWy+yWAP6AInZLpnrzSQG+Ao0ytBb38wx
MrQ9mFh02jiRiB+xKlOcw/J+n5p9OMpe1mMwJkuVus+5dfDzmtzrbW+1yQ2MpJGR
AG5OLLFTSiV8tO/fUk3sRds1sgqI5Qdr/XD5dpX+vRy8oOYsB7Z23ZpCc0X0fylh
izCGa5tkKCfSs9zIkqQrYO+fAZBJ4cgah6lAKOuq98qrFq1PFzn4tw8uCdRgK22R
ooP7pzwkYXzerjjtGiw27V9CM7oBp3VYMuAza4HhFccvD8xyayz+ZKV2aR3qxMFG
ubhU1KjgBli2tW/uqyZldgaT+35rs06wPdlgVuZ4+fgcFjf7wOdOy7cprFr27iAR
EncxHil3mDH2T+LpxdMxQOF0GWLj/2kQSkvlybfpwaYbIK01m7js4/cFFq072uTH
Pd8mS3zSPvYj8aGfgvjgIO5o1yGUOrKO0n57r3+EF7gNz7kohfCFIqNOZdOdiwVd
YwDcafrS5yx7o1b+cl9bibqrXNnRvkrAvHqIQZcHXuL5a1PRF4xhy9nqDMds7Gna
qrI+faiOU9yoPz8m5+uY7WXaEF3JG/snJ7VDZW7Dz6FLp7fdW7u5E6zChq8y96k9
kK28v8Llgf43c6RtJsFZJx0eN+JX+sz2CU/MZHAFRS2WNEsOnJR1j00YQxPrjEkN
k5Q0HSldJ4oqlFsK3pQJH0r0aXxTjG938EimKjAyKl4tKG4OjnlY1PDVTeMLcv92
DJWvg9j9QKoGvAgMijGk9eKbOf/vjsMavtBwKoDvMuAWQ2XAw/DmwGn1E84LrY+p
4ki0Ffm1X4qNFF2l1cRP1uhbp6rECo/2lu+6i4lpRYdKXW3gYXt9IS9OGaW0mu7M
2PQC8JOVt9dmWCc/QR+QjWmYZaFHCCDLrgLK3baeVe6RJEbqXAQj5OXkS8BkuF8y
Pka1s6lK0qS5zK0adcnTzgkeOzXUsdtpTYBBK00KMT/c63ydjMBEp1wFEkXGhqve
hCZy2M75/U+BTnjOgK8uj4RjhNHIFxb3XCatBmncAh+R6g/J4EkavU9iBdMXiBQ6
7NaC4KVOqFS4HTqihCnSqzOGxyRU+Xmtv1uudTZMWKBWt3fXNHIhVa9t9eHbLz32
xVRGASqCUsfknpHfPicp+W5zqbIoqUn93UTJ7ddwjfBq4wt5iUJWNM7unIhO5AF1
XLaK5x7f1+fQXEdymI/eL+GKdP2sJmW1tzoTZGdjSqeih/txz5vhEneqHjG+s/tY
YFOxqe7i1lMBfQmp4Au0ZNSPjpBriuDx1EcNHYoUeytMLFfimzpRL/bt06k7kRQi
W7krXZN/FJxRUWesVEJzYnQiQz12RdA50BW9AyQOZRtery873N02C0Tb2YHWrLRF
iLZlhB9oGgdzfmT1WCvZBWmmfk866UQvBriX6UAuFjT1QgLFKE+JMbpFnEgjblE4
pOd0aSRv+W+SqLCTaCM7jEv9yGXQ1ujHp/1vp1XBRXn/eoJw598oxWFRgh2AzaRN
iLJsLfNUeDWUUWwfogzcXmniV7pD6XZSueqxoCkNEmiwRv0+bDSl++0GjQdXSb/3
Wl5AmG6XEize9nF2b0oNMi/qa0C+LwRR6I7rgTKpOdNaighvLQrPe6VfiKQe0Yjf
YqbHO93G5sK3RUy2ZWapndOr6/emlvxCMExq4gz1vcBmoeeuByGzGa8iGfiHV3ZO
gJI79/7XsAn0eXeQ1Ay9euGmUKTCIPJg6sH2Cg+kY/Ww2vqbn3VdfUW6YIl7xIKP
kbTohmqD77Xe/KDxs9/of42Sw1ttTbLo/Nvij6uV2uAkq5+Xao+9ZCBjUZK/ZGUU
VMQkjvka8EYZXQzN+J4d1Vwy5eZ5f25qx1dOc+2ktU0x+tAX8TNuNJQ+mR1aMVE9
ppNMQjWELbibY5TkzXtSCkUebjqDsfismoYvWYqi6/I+7/7W6KuoR/WXQVUk32Kp
BgFPuE+e9PhcU6A1UTVLKurZGN+0qpGH8g+FrApV2qv66VcHZXRDT3M6RSp2hffJ
2qCLvyHMdTp3nesqLiEEyFP4jNenX9tGuJ7+NNg2tosDii3/lbUrj5qnWOzv+WVT
vnxA7Che0hGq3QMGrN6Z0idi8W3i47PTfBWsuVW/6r+WCi2t5v9iEwt2rtdHPASr
ajUX3hNRmc7q2MNxZUH5DiNQ0uMLiBgL5s5EDuHhdVaknvqlDnZIoQBHIgAMnah6
rvCst+IqAcShLgopyZ9Bf/g+QyLBmq1wNuWqvDeqBlVjspOM6yvkwys0XyFESy8f
HnJzJ3mkj/mNb5kIB2M9w959zOMoD8n2+/nlrtKRGBu98wnQI0JDY00QOvQR+RaK
nozaGhQQQLZkkMwTJpY4hbcHVlPqMnPV/pRdkwm/1KbzdC24vsAdum4lGC3gPcIo
3ch4fhy8BY448fvjai0pXposmvVhyVERMSgB6w80b4YoFVxLDG75rucAhg5BnQvS
tIOtkZf2+Z+isPWAllG2bD1n5iFwKSE8gkNX/6EspXTVCj7NqlmaD257M6ZwnQjF
TIOtRuhVKyuiOD+qBU685RdKspweq3L1YtVfGhqgZH7iWmcrM4US47tPGkKCIez1
NsxTJwq7kw9NmVisgudrMg8/7oeF+alCyzB1mK8LmA62tR3CjSuTjHwnbeqfGfOt
DLJ7BdYlPhRrlPhT4/5BkxKTPQuvQ/fGQDiHhoS1lD6SVCzJQZ8PCUJ1EbcqpD7X
MUwFWnAwJ2lyMMlxbyiGNpfDnaeMpJEUSm4guVy4b0U/1+gcUi9fgLfUcyGpxq1i
HhLW4IaebVAfKfJ/behHcWzIeFTS5+HuTw2Eye6eSWt+dzHXx69qRa7AAwZUKtRe
svO+VmQ//xqeExPo/EGEZaJC3tPYt/zZcvjLh1X1nO8eLROLB4TRvlJ0S6/SwwYv
03CJhPTHkOJQR/TApyIx76Oso5oWc4lPS2kwcuMciD0zizaf/O0tvE77PB1I73bu
yOzYcL6AY+8FeGSLnzS2oqaf90W/I1VPP/d/36xpkATxOH1sYLbgJQYyyM1JgJux
OoFiTPdYdwEZC2eM0L15m9+Tnz11nTzC2x1QKB742htaRhdcEYaZ+uwcvnnp6ggg
fMWDweHIZ9QeR6/Z9MasR77v0RvB67s2xJ0QdD/b8O10tR/tQO4FVBRs8RPH7EcZ
tmffk7IIPYKHF4k873m69iE0BW6RL/s+LXrkorLd+iRak3Hph8ZOyuLFhG9uSLsE
Y5jxGPVu2saudVN8TYOKba+x61/CBne2Ou8hL/NshaHw0MQSt/01+LNoI3AqF1Oz
QAT2B59iqzELn9uJz4aG2CDWu79ZD15rC5HCQgwO5YSkRY1mkH2xEXdIHHKIJ/wC
imqz2f+u/RT1kuU5BTVlUswoPwzk1Eln5py7PQjnSKv+KqtS6OgJWNdH8F+WALnW
fBaRP1o2yreSv22VGXyVrb0wC9P0WpYjj8EVKGpkS1Dk4nZ9CRviMvt+se8Z6GOq
Af4PCUTB/xCTTGG3ULYVLOOZAPOpvWnuMDzbgDbrN56XqMzyGEI9lFS6Nh/bwW+9
KYjypEd++WHEV6a3Ac8xHpP0tzvW1qDa+8aJOF50m7ZMsOMRGhkSCLKlsznyy1k8
fASzs4MAOOj6ykuepBjZlP5MYVWpkAiHPx2/vRQ6mIIo1xkrpqSnztnElP3uJFCm
GBQ+aujm3sp+p8FmlWwhJ2a4HMViELVALM/H8nUUTnUw3Uj/xesY77XQvsfmaDrW
f2EJjYaMiyU7tlqj0W0eZS1bbh/qSy/rY98R4aMypq5p0tGvFAgrmmm58K+1kG+B
1a+iwQ3lZZ+SSOiEeIHBLZiIxD3kZFOSvfOPaCliv33cAiFGt9BECZb2cTNtd0WW
MzvxBczFoYMT6+3Y1hXs+koiNyv8yaJVakDHa25h0MkTrWQ7oUY225paynccmVZR
ipiQhhTs3wm2Xjc1T7QPnSK5VYQK/Mjk9JjMhvH5zIkZemQnFN8xPGtXrpXk1z0L
WmK+0iJMnnMkfPXGZXhakpOI6EiKhmag8NODZVOQip5TmWqe2DgmYnfi9t8bYx+C
VrM9KjogwMSQj78gKsj6uTkqiyyfuFjG99aHCiPqyRw5yO/4mYEx8RpXQ7NQvucD
Rf+hjvA7UDQPu+OVp5XziPyk2AG2sgmyNsiPcBk53nCnvfjcS7K3oii/gREBRe8L
mFxICQispXiJSbOPAkWV6tnY9OYD/IKqViWBo4Z47umUsgyDg+4SWvDeY322pHy+
f5nRuC11kpnYXiUhcf2awpJYTrBspTsTN9ALQ4mp5A1/sGRw9siymvzmQbdiZ3gH
80AmbH6DO4yOWrJ/4v492YDc4OTzdGy3tNlp2LhYdAFTNNIS7MXx6ZCkEjh5X9r5
RndriBg9eeHGt+5tPVpqxp+o2dIwmL37SHQdY0UKx7G9SVC1znjFhRRBDea8IfC8
5SDNNXvigMAbcNvnRuyhXt/RB5vMXbmf/SNC8WFqgv/UROFwXa5S28JibFk6nRX0
SoaLf0NY0BRI+MxI6srLlpTbLnWNcGXJunbT2+3gMlQebCDzbX0fO1eLdnLH03MH
mX0GstwgakHNpWU4ECLFFJ9JWo4XhBzJq7++HqshN3xWJnrIhnluCfcLnkGQ24Ex
IOdysf4egQ6OkzCUtLpj7kngzZgcKzHDn588ePzJ9WmCxlKGE3c7qv/F6ok0AvVv
3X3Zh8HZ+EyrkzySIOokDxz9c+ezi3n3vKm3fD2KTZBHjyxU3H/RNnUTiPQIMRZy
cqW8sZbmMrAqMEgcS4IX9zs+hEy+wxTaI7zJXQboucvXsMTsMNsFfpkxVzUAj5ba
e9wBNJwtRAJLVTSLW0bgsRIZKM4PIDTZIH6AhnFoneQOhbfPQ2QUw5OF7MiS4nyk
XQMUwRxtDTxBuE8KDSWYOYAkYntcBTIi+A8RmEACQgs54ODUk8WMJEusX/JjWApz
mpBhGZjqZuztkNzEu+LK9XoPMK7xjYyw9JNYSAzgO1TqB84cNOlpxETieGKcLMPz
VX6awkS+elHLQoZLs9InoSyC73LXAxIRzMe2EhHXspgMuJJnUiwokCkA+zFANpfN
rWU/Ltm4Q62D9pR6pBw1lxdLleVE52nnHpbR4m3emg8z8udyQ4z/wrBxNdoJ8xyY
3Do7Ac4X+9rlg0AsbkIoXE51uMvUIHpPQgvwuKOttzSnnzAWXE8mdJWCIQ9jyfS2
IyDcmGZVNlcNktsNoo6AYrmD/fzA6xKPcfISGOtQoZJPQJ+mB0UXnMDTXatflmcH
Ya3IrzXrCeSMiATQY2vsa0JZPgbgRIAc8CP/O6CUMj7R3yrrIPOimp+Xc7xUwIch
mcnBFE5wosIqeQqB/P9wfPS1cvpDTFn0dzG8hNt7NIOpAtayPKUzsiS0vtdj+lir
N/pXBtLbcc02u5JhHzAAqFNC8JVAtSRhKaXyOXBsDsA0uYbgaYRleBVQQF45ju5a
wGywKZGARoi3B4rCzUvJ5ghliKUt4/xrjl3CJqavb2ibhEBEwOJnGSSUiFb22AN7
WEDbXNes/OT8kYsTV8hmO7Vw92pniRIGNrt+g9XOqQO2QhcSHjjF02+u2DJ0z3qU
TZyvDNmHZXVgjstQi5idIwsCuxekWvFPe11otlib+NP5qdHRoCbCyAlCVa8zitIH
rDxRvOit5oF92tQS7GnniIScz19M1TT8RuN5/D7GjbAI21Fg+SrElcoOwCQoKcHX
/9wKi5DQWa6/T3hIhhZCXdJ+eCPiBPo9hyExLvEqp7br1x86w2TnXq4b0wrpbX9b
gbh8zfmmfy/0jNvkrd9UPWJvj30yiv5055IbEB+/yesFgO1ScQPN1tmIYdd9djtD
SSr4gmhoSIAmMKuMNLK9+mZu1vYA97kpmyElX0yeBrbYmKqlOmBR1/b0vR8MfUtL
p25WY/bmykVECjTU/R9/TlAlM8AvsUBHx/FmZYsVrwfnIBiCc81TdKTd/9Ex0SU0
/fx702hAvqiL8Rr1Dob4rB+i/hqTKikp1JtzGI/uHGB3T6OPTdMJThRfeAGdqeGn
xM7GLYbAhy52uEFlSzsomLEmAkDfOBWIdaFbBTKJT7OOuiID36WE47x6cA6Dozza
RHb0JBxIpUWR/xl0vNAI9cBIQG2uqtkbY2snxcvVLds4aYz7Ad2vPnoX6hVXSdfh
/cESnQOGKDGx1AMToG3eYgnxA0ojQoYO1H1OIoGZ9zJoN8Kz5pooqGsJ5RA9In6X
8ooeorEq5hZlMhaJFXYMfgperw862zKe6sPbkm6EpgQqi7Shvw1HsFk2ofDr1wgi
ctf0pPRwh2WY8xqJcicP3R5055ORkjOSiDVgMje9TlkErmUnrFbnpmz7+lAVbiST
Y91g5p/BCywVv3x7/5wlduj20bLCgFGeKP5NNPb4Ja0m17dPokVxFHQsyGfpnG3q
afi7IA449c4lflXPItiyjv63z5/b/1SKiNeXBZIeKTl7NM4c7u6pxdKKxgXsVtP2
1FLWgb7AVB3757SOwfb777+RmVlhj27cKFQgOHR6NMdnaa6VaCBexn6jn70EtUPS
hCQLrbZ7RQI7MztpabODP0pos128wOE+mkwzxEZgcdwri7yUJqGsS/wUXWeA0eZd
wtQSa03ykAaq4BTRevDtBIjAXcqRyx0MImfnqkM5r0kaJIqJOr7WppDuPCMO84Ev
EL1Jakz3L44dT3ZXRWWg0HgpXLzTRq2TvOBJeKSaPSBTB5gXagQvnTH52XMyVUVx
1GobxZX1to+L6F95Bp2v6VjomV9d5huPYMfQPjYGeLXE87TPMI+M22fROwHCNppG
6CafqyHnKl/OezlexEH9AdlSzZQaoAbCq4Ti2x4nl2At0Cg1kFamwDMEYnegWAi5
CiaGuCA8Ued70ycNFdrnD9aglnUdELIziraZs4lSIoiup+BOBFPCLvbx+/vQ223X
m7Y4+ANfqL1FXEBZA2k9D1dysWdxFvm1Ge2ie1ugq/H1PCOeHLcdfp8FjDzUdwyc
LpUGnKpbd7oW+AygaSn8v9eXd47KC2hgxPcPf/RtYTZzR8uKXc7lx1o6VpWS4JFT
sUT1y99SSx8hCXhhoX8s7/2bHR8mdAzP4nH38Fy6cDwIrcF/a+QZdVvztHqrvZ1g
+r2j4sgs5jglRnLCRVVReXM9eAPT+K1xU9e4K8m3zMI4jVbEC6PkoAoGNKz7Tn3b
J0/hxT6YoUzTfywylejqhd9tscQceErgWP0CSEBT20TDo6R1SL3PQhXxwZCRoAAD
wT2CJnUwdl4Ooqv2jz2n+JaY1v64f6wQMHV+xmy4gWwYkGnjFh82q5QZmkw50BXS
IkVD2XqAl0xiOSpqrSDxV6yq79KqlVvxod1403nFlEisA5Fjhc9zkQChUrHrK2iW
gmTBIzO2Ejwt+siiYvVrM4SMHuu1kZyJAsoPI0n1TGUHrnnuQcUxoEdTwRrRpPwa
gdbz6VVrQJ2rkiBl/WmvvV5nRHvNsUz0hFjkzbi5PeuWbVp0PhbfL7gjzQCzNbVr
w8IgQgDTQe0oZEJG1p8n0QO82Rh8e5j1lP6n3Vs6LvWljM0LHuahZEjGKJWNVxo3
gJkWqwVyN4QxZWIWk/0uJljVUemnKx00dkHpgweJHaXXNfxN3uXhPueHYXuEGbL/
Zm/viQ2Q1mYsfd9NIzn0kOea8+5mVKt0ddy3x7B1ZrI/BSUF4AAMPusekKug1c6d
xNkpQ0Fjl/DdikNNle5lLrxSg0qhP0IzBnAKKOw1egTvOjwRkAykTGeLUFiTzf2V
6vCnxEE6FMmxKojoQ/xy8vAysGUoPw05/TXcnnhtmgqeEasvPYODS3p/WiHY8ZRM
cMHYAtHDR8PnSpvqiMa2gNmwQG+EVufOrozuVJDCaX5Op52ltdB6tAGRDXTBKp5m
DaRv3FdAd5XX8Vy35nYhstxUlHWdN1Y40Y2P2W6Otk9KorD2P9mNFDb2KAPVlq2D
D1CDS/YLw0+BduVNRWfGD8v2c09AkKnppBbRbQLtsv+mZJ5UvYt/nbHhSiVPACrI
2BedT2PjEbB3Bx0Y7yJp9lXo0ZsV6m+kinP3Jkj3xNOVCa/eQbocMA3MQ5QNPsYB
pg1bkNCtWnW6kO1iKqdKvN8Y22AcUVYVQ1hmbXT0RwlLiF/F+Fr40svshJGWbhWJ
mzFKTP23L3O518N6lCpRhfJswyq9umEdCPxTNFmppo24scv9z/lbGuyaaMuGvcqf
iCjP6XgGATvOpfTZ/0wM7aCE1tKhMmeX1bkJwNoPS3JIPT1D/Zh4R4RWBwNJj4kT
PQT5b29F+VHn2vw65oEJMcJTzooy8kEKbMudbrpNiZTN45NRP3FxiwSUSuZiTeA/
WGa0/+PCp8XQEawhFGJc9O9wqNP3DiR7q1tsCoqhR/NeomNfnMM8c8GT/lqlEYyn
e5umEbOb9sofbs/8+BnaQ0pe06H040JuN93nS3jFYYbrUQY8NTpUwYPvMmjOXrFJ
KR9rZnrqD9Twawky9Uspyu0TRB0MYh9RQjkn7wBFuOs47JFs8hKZdFOvaPC8K9LH
Bc05DR9ANymHdvLFhyv1ooSc8Iug8pLRt0iblOgtOXUuKzEEdow+1OybDYpnFmkr
9Md7B02auNguWOnvxBpCUsjzVfMLD2cSeXYPWtzfHzH5yDVSg0qc7U0grspE4a7S
rbj9M8cSGbGwlSPA8DIbgHqib7T+fmN5LTC9Dz/cID7akH9p5BspcTeWCZaW3BjR
f4p2DTVQ9nhrYhD04ddgYHDDyFWkXSwijV8zjbfkLyLrGnfPmFqYW3+1zl/jYIYV
otbdWRr98bg2hpyc0dN/PK2DG8UQuJfWY3xdR4Jz8ebZ9YxJCK0wdGjp7n7w/kBf
lxGgUEuWmihFi+0R1L+7MJnvEMohY68MKOjW8zb2V1dyB0fM+nJSPD219NC//xqV
OlvgMLyzUzuDTkW4HlbHG8Kv2cieVvzDagWA0huWi1wmLMo9BRO/krF38tTzQWi4
XNKVwtQZ7xfWkIa1/1MUG86gjcSZUJs1RLxNk+k2W79asdu2I727Yn/JY8ArqnUW
QyTzEKDI6ieTnHuhmWfcN/5xiTQ/fLvjdi8kAUM0m2+1ySWixG1IaWklQVgFv/sx
qn7+IFWlQGijPsJSus/9DIuxfzO4qEiogD/Za8rl4WUAagrYzhsMSSionmmNhKl7
AGEsonMO9aFAxn17M3IodRY23C0eSPesK46f11gTHl/ZM0t8D5FHepKzBOdv0wR4
2syJHlyJUFGkwgCr8v/FCU7OuntW4I6aSo92/ytnuUbMafRXZWltc8oHlKdl4h5j
YygQyOYR9wIRFQw04Zrwi/L0OyekYG2TlN4v39Ox1soVANfc5N1qtrj2VBcS8tPC
JW6gVlATUUL9jzkD/JZdBFjDsi9X2UiFi4tVJi8/+UlIa7gNaCDJ8uTWqp71MJKu
V6p7osIORXF2RBbTdzOv7XKTGU8HLDivcCaHiLonWN7tc/odkEAgQLpJClhz3oql
1pIgIvDtJ7XqLmg3S1Bhh3NArM/TlxLXMfYlY1tuArO6MkdatT+YQZquomxcuCnZ
K5u02mX3nBE59FpeaUkPtCh62ZkViodnWu7R8TydHqjUqJfwNauBFge+F4pnmBfr
CSrUph+2krviMNzlDveARdYZZZ8QtIoM+0XFBX7nO7LN3+vXGvcbnlC7D+uru1QS
tGlAOXjTGawNpF+AWdhxln6Ne3CneIEOUgxyzvBg5r6JkbisSlUD8akGFp5Mua40
hdMZVEp+aqWy4tSNkGwbkmbv+YV8rieotNQAiDlOaixA8wXekwZSxcy7mnxxjJ5Y
vIt0INnZaI/9n8sC0kpVuiEqlxOj42yHzHakgCR+2gZXNjWUY+8LeHLW0Pq4TSaM
4wpXFCBE8KOSVL0t8IpMHTy7W1Zdm2XUHaTpB3QZFcaFu0zMWevC5KEmg/I3fgyL
bYKb/TSDXBs27QSNtZLh2+VBKAvQR9LfFaNao45Wvks7QsM97s7hN3HIUbA+TOZt
pzEVRbCkL1aVVGLBXnoSABSGOfEkqrf69z720HSth6EStgJyesQ3OMnLqrDP14EH
HUdA0NTCYAqG+R3YCfSu4KIUpcujB0d8oy0JjD86/sjuLA9xZ1gxPFRICQkNE1mk
gVJqTI8BSxoIAoywqJJ7jr+pSI5zhbC2kdmRg3ZRWSMRBKM/6Cnpa8LmgkLPR++5
zND9agDLe8E/8UngwwnMkc6CQr7zmT7cbvFr8KHsS4Jof4R5VJCuIW8lSx3jW/ry
4TDEuTC1pdj8qR45EJFpBM8IltnCGTD+uDYr1IumZ5/z5PVE9vWgb/1gvFq9W8ad
TMFuaMS8x5LaGE3lFvlpTCWVEVnE403XxhviTyWwmM1BQPE2KOlO06UzPXtaoGQG
Ay11DMgVMqh+YYAF0KwY9kc+w3E0DP73DEAMrZmSQ2LPuyYrPJpSe4WDtjqA/ols
HT++K52+vEoQ/ObWckxw9nMQutn9gakgEFtUYSLGmOrvk5P3efoOGRPwT8Fl3Wcl
Bh3fpoEodkdGuj5PL/cGYyQXvdprInXHm/aRWSjGCdvmHhz+xLkBt52XZ/5s9dbG
QFb95KOYEXd8/FNswduDtVrU+ZITXn9lnSspPi78ZDDA0mcu7fFMmegyAcvMTN/m
UtwcNKSpI5SOYplLLuVK9MDrmcqSOWi4sl+Z0xfMihWdLj7NKntQSXFyKQ/+QLZ6
ThrCDvfiElIoYRF0dqQWxXPGrgJJIdpwoa87zVPcG+dEtGn+Wbb0vlgNE59z9kd/
r6hiAPEc5fEEOC3jyNREAKQMlGSUsR0TEHBbKCwPyiO+0TJC9HgU2MaGtsZuQA9j
GWcoSQN5rCfYoRqyAHVEXs0ngQLiW5PJ5et8WMCHMl4w46UkRhUjtHgKaQPw27yC
rnS2oi6amJ30offYxp7czzhsuyOTMH/B41fAc0rqmqzpoBYTRP/B7czCCSKjAsHz
yJmVI+TMh7PYNPX5YCjKKF2XM420Enl8OBaKPYMFAliH3RRqhyUUHsMfp2ULC4e+
VK4G78X/F3XSe2Z11SejpbDHl9i4VAeIHU1eXXYp5qgEF5OG62oxLwCtF8AmvnrW
AZ3wNtRHcNH4ugjIOI3P2MncuLpqgA6l4tDdh3cputtMxSP8TvfKvPFYlxCnLz6M
bY2il/Z8hlORP3ddUuK5VMxTngWG5N1z/wMKGfkTfLkZu3rupVHY74/QrMqeynzC
nb6mWU/EpBF9un7zeCiDGoe68jN3lIRmsMNEJ9AEwbZAI8j42TqsfZdOgYrvrVkj
mfSCPnVSCrp+o9m8rXvCZK7VBYAUI79EgBrXHbtncx1HFOkzRAkff53V95HHCeSa
Ehyqzb7jUd8nnzu+pC5q6WZiO22DxrUxKHN+6BLW48aArWR4+dMV75hC6En8l8j5
VnBV36OGhc2WcjfVzW6xoZuSIBZAJy6oIKyRhCPjGaKPN3PtadQcHiubg4cgzLOp
jrHJEatnCPjIxiqCjjk+oTwSJbKE2WTEkBioEYvYu4v0PPkrSIksFIlVL6p8WFK+
nTMStqlj6P1IHzS2pKaBQnwBSHvJL0fwPn87jfzPE5O1IVeon4pm5cwRol+fkhcR
Jh8FC1G8UZoWewOkR40iqjIeS0wdMgjhfoxPIlzxi6ZD3s8mX+CN6W+zVmrycefC
reXEvxj1S50PgdBjf6ByoPFeKQ1S/F4gYaCwlpgHaKQCmL84q9wGvcayNbWRa3Yg
BbwehUMQ42OsERpGFL+soH5fvew5BOcA79TX4ZfsFbC/DzegIUBJyugGdZsYubJT
HxNQ+KBOvyPsB/kKsBhJXjTyoAL/AIbbNh3dbLTKSZsIzukh7eHZHCN3+8XawMVY
QWkirnVvlCdFQsKl1giu+mupNoadNGliTMKJtslYt2T40U7u+dQHpadgdUHzd6/Z
/te++ujVwwxIEpCBbSKuZce1Xpg7iGherXOOKH+6jMxG5WfVUesBc7+YxhTGIGtT
Zkaxejh2Shf+oFwLqrVlmGDXkfv8gTlwugDSWOWpclOJKJKAbdDZhj9pl9rJx0z+
0N/aJ5M71lARm3roRP0Wwee+B8ASghU1hXkqVI6pV3NqN8m74NaeFHlsJzkO1GKN
NmgOrS0bUx55TkEGW7K/6fLwEBhBJD9f4UZGG/lmD1G1wCw3SJv6IXH1kx0+57NU
0Vm6EMeHg5xJEQTIPzoo6JX51FxU0VCRFVIZqbkJaqkS4PZvoZoALyi1eHbwKfCm
cu9s1IOafhxX3UclaXwqBxL6Q+GZ8NsDOGYOW3fbrGV5ZgjnHDX3s6ijaIfUhwVP
OgwETjyGZltKM7DgRLsu5/9IwLXrOdXYPAiBBTW8f2rt+/NFp7V6z7pE6raaJlWp
K4y1e8/70XXD8fumtw53fhmd73iU7omW+B5FSBxyJLQ6XlFypmV/lMfGC6SkHmw7
vMB091yJeuqNygdPht/y/eoKWBllio46ww746ZgI8OaG/umnJCjET+c43/z87/IZ
sxuFIPMs6d3dJ/eNsT8kgW64t1nB4ZASk6xsCT5B07qPTh/ZeH4TPrh59iSg243G
pOiC9zvjt7GrEwQZneyXpGMWSAYoqdu8X7cAij3aIEVsQlA3W5FspwZjSk9YIVsq
fxcDex+rELEhYGW6NdNg54Fa2Gnv1k1HFccmRvcVkjAI/YiU+USM7FfSnxGDfAIx
U6DQZim2O5E19Ho7FC1KevBjUQ9DlBG6+XHWO3lCcaopLNHmuUWZ1559SgIH9AEC
pURvUnOcKTlCBv+bSqpZAckF6LSBfehmoLMjTF5QME6Z1BG8iWcKyApSGr0eHmq+
PBFCYovyjPtg9vqrWR8rcahLh1Q3UDR3YrUnV0mdwxOuHj/cXejDPzyPOmZziTuQ
9L9BLNEfjV5KuWa19EDyo0QXN13REP/NrdHddHKfcbrb3xblhTg8xQxadH9jAtcU
MZ6v+XZR3maG9vP4OnfCJLnXnwL54Pw1NDluqOH87llkL5x0x+alEO2vqGl/I7NT
0VdGuDBHnL8e3H0+Qh+xpkgu4A3TN5emDYvsZ605A4atxi54suabJL2tkfNUca3U
3YcQgMQzk4AVQhNTV1x5OdzGMpEnbtAI9NTrktoBtL/rN+mIxV1CwtYtS+rUbg4R
/bwhWKZ4JCh844cGJUVPxdr30pH2UYG57qtS4s2Gr27TYIoOnZBSjMCWIu+Klo4F
nnqQRaSpvQ/7y1FkLRogf//kO6b7uEDAPydNaGDSBh0Ks4jrr1er7DoGtvvJ+AwR
vwwACa8sutgl8bUW3G4aynwvkvsjV5FM+0oUkqzgZvHFUyn+lQTmcGtuuDAPLsvp
KhIxKZWDO/pfJTd9YoglehmliXVJsJcm1yppVJvYMDliFRNeLXEWgLm6xT+AF7ZS
5qMnHlpF0/MSgL0G/wc0IHg+YaoMOUYAML3Ee4GwPvsstJPyZtO/vVgNIbq0RAO8
Sbb8BmceUv8wpdws3Y2SiSpEOcPqyxBktf2cPpAfp5ND3yVe7zsv2dCV59vkIf7o
QHu4umRWUpb1QCVTmfhp/Rgme3b6TKpjhD7NHU7tJfh106tw9UP4eACSENXRJM9Q
R3LKVUQCxomkN01dlxkIxDjiEa1Cs/WsTkAwJX9HmDcciM21ZRCcJ+po6eWtMZzR
RVXMw5R4KEPfPZpqObduuQw3T7PvVT+22UDQ/Q4FgbqmjxnuS4MyJgVw1XwvaaTn
qa1Ulq8ORZSEZzdzXU6xkLDK/JqmA1EfV3JVAlKqyQEQxFJbOjmGSQxWc2O7dEbP
k79mdPgM+Hg3RaMNdloiC6AaKmVvkDgxPTUy9+/HnpLntIAtxQB3G1j6ulx6dMS0
t+44t8Zu+zBsEWoZj0BzC5c8QwBG8Akz9J/XsFGyU00GvcqS8v9Vx3mFkiYpU5Dv
VztG8BbRHHQzM/96x7B3iwFupSzIj1/2LCXjrPBq3cN1jMOEJqvDluaNXGFZUjrF
IOJP6H9NAipopyMXEPAAbeDrZlaR9MoSSQgXo5E2pYDYikGpv5C0nMbgnuoU7nml
vn7hsd9WPAr9vzZKUuZkm69Eyp3ANz1p7q2a9lSz4a3CS/pgMC+hfmOkpdiEF90b
+hTi0xmWAmf1Bhfp8mktfUMRTe253PiZngY7LBqLsNbEUlmDP4HsuDNghD0/SWvU
3cyZ6ihnnPyPAsnBglAbat6cF9jYoU4P/nsZQ1NHzSz5wfh4+oao9uEIbqOxBuIu
wWqdSDjx2MwyTRav0OG049+b9KNXLqiMFapwN76UTOP73xMOj2Z+fmr7D0wuc5Ig
DhiEP9JYgtgZ4NP5bsebPo2K4S9PaQ9SRNKwN9rQOGCPnwEYKiCRj+Lim9GkzsJy
LsJPSU/Mz4VsrxXLVKE9vWpdC6DK+Qz1oN/qZ+4SD3S2UfeIOr+kFD+HJca6ll0I
Z+9Ez9mVmrB33FNzmtCIID7jzH5LAaDM7ndTjm6HJCdAxNe4xVlAo9bQ3P2QtEAR
/qRrVpl3WkXcueeS88MUSv/1f4ixG/ay/yklcMA9tQBuDErLS/xg/0sPw7My6IPX
Z0j2YotMcY8FohkhNW0/quXTYtaGOU1DrZEp+/04tj40N2m1pzoyAFrsefB1dF3c
N+qrZHDYli6jvFjYkpe8zxJV+IjCZD3Cn1jLSLKHfO+akfiEi7bSWxG5B8SOzl8m
Zsm1FDE6DcsZkNT2EXCb3SVQJwSoY1dLMxuDZb7hMQxSoj58LZ+cCfVxuUSvrnJR
c0C1bJ6rR6uVhdtGppGISzkkMibK8j0W8vU30i2OYIbIvWB/8b1kCdg4HMvEJdDJ
iBMUGToWM/+/yhwP5vVmoNtywitjQ8RXmbzAvID4PM+EMJzIbCVMW5LDXyY41dbF
pbsrOsdHfPIj5oDUg6Xc3ef14lo0w8oAF1JhvhgWAkFHg48JJsxdxIg8rWxKOIBo
jnVck/vPBJmnAt0xuAqNCW7WGGkIOaioy9GdYgHmUT/1RAGt80Dz/m09EbgL8WAJ
foeIyXFKYdxnusz4/lB+VRlncSFoBcHJIGzdGE0Mi2khrgscUKzSDlhg6FuxbbEk
5QZuxxv5AkLEfVXMglId+GhUHzOpc9T26d6NpfM9OeX1uA4COX4XU4/BhhBhvT7O
qYimM6mB4J7GXz0EhisLABihLHBc2EFTrw+etZUXGI9gh6DOtLo0ifOFh6dxMhWQ
CBrrWVZU/901SLHtTYOtlU6HuLr+97pkW+CWVd019fSw65sOM2vrAdQqhUfEeklo
PKA+e+NmylnT7qLxif1c110sGN4OtY7jL/Shmfm60bNeXu53picX55Ao3Xo0f40k
c3MbCKupzjqMWY0iBn4Z5RprdnLNcyo5xqHpX3WO/+9XVKjRNhaAf8Hv1d6gHDgX
QDyRkhhiMJzeoYCFdsjybxQ4H1EH5CU27cKSWyKWVwpulbNCChyPEPLY1uMT8/c8
HwjCF3Vj33eYbaJG9PZA+7p15mc2f/YiOecTNqeBfvJY6SNK1KdVeCNdcdEulbCI
6R63uqPx0KAqeExHGehg72xFbFbjkO5kc0LExTaK0zhGcWCKFWvmeJxF4IiXfKsD
qRPzPoZd651j+GmHk8G5ZrnOSIVYK3E3Vfat2n5dhMZ9N4SOb7bzwB4AHnGTiJyp
ONGXQ5Xh+SETJVakKEKE5oq9mgM6n6az5Y26Q5aWFqrKIzoXC049E8biNEyS4NNP
p7gRtcB9WXo1IuOvgfTwDQYlLe46gJVqBzVW50DO+rsnCwJvIuLE4P5RPd141tTB
iRKsjjCaiyjICAVmAvYLH7qMKDObf00rMzd0bxjPomvStDx1OUqz4Pw8J4whHsKq
NNKRbrr9RfyidNmBhISEQE7IzHaHuGK/9UQerbDxFoeCIXWqmZuSDidyL91vF0cE
OGBbuwc5ZkQxywDWt2tyXPHZN3tJy6i7HZBD0oyS7B8hO06squMxSoYRdVXih9QQ
0rg2uS1cqYLlma36gDNHvtnHnl9WNol4dI5DjPaL2lVHwcOFYrozmxtUb6JEibGw
f+gDKDqvYApwWHasQ+uiJ2CB6QCMaWFpHD2peICwzkiyYzc1pDCBUkCBVjlnpnTp
XWS2YuO1HXrXRto+5PsqcPiw571bwHoj4Q4EQUW3PER+fGiUiaPWcnpz/kmkp3k+
upuL5jChgpS1z2EA9LRRojjx5ES76wguY3wfS0uNBIsVWcfa9YVeQH3oVm5wROUz
r8T6V27Ztty6bbi84zDRURS13cf+wpZLa9+fYXKhQsgDqAvbaUPt9huF+4ruavQl
IW6fkaA5L2nbwx1x4y/iYNcSPIsKXiThrHJyw76OiO2Z+TG4Zdje7wgTFdcFk45A
y9z8A/25Ofwaz35JRaiGKse6a0PkbiQ44CnY0NDj8uRxLrOORH6mYSWip6TBNrMH
ub4dpOgPX8uBB0dy/gR3zDT/0jCgf4pWKTpGjjDAe0AaSBHy36jtjyUbiBCLl+oN
HwuOY7/i2on8Aq7KTEGXeRb7NU54X2sV+1pmWmejUP11XCgHp1JyZm6GEp3BG6jo
hQp8S8hwTYFXFqoDRI2YyNQmOILBm8Kzv77HjTF8BZCIDgrzJ5LoYPm5M6gGHbE2
LKjQ62ykXGld6V8QTWyXFx3K7xbVSdRuVg0kfw0zQ801JzD6YXaRFWo88Y5hyP7l
HteYZpxTdA8ahj/SWndioKXCJmYLjfUS1iGDKzIh/rboxGKqH5PCgNhDkCiXkTAg
JkW6htOs87PSWGdqQrLEXmTwRoA48QcWOMl+imaT1zzet3Fw/5jESnMLnyaywsy6
a6DVNk7pJs3O1gPGO1et7/59/qroDlzqaKQFepHDN7DPGwYLHTtJboINOMoT4gaj
RGsdT7EMoc3Q5msB1qAYuhDKjXeyC1zT37zoUXzyPq/7nu1z8ON5sn67VkwRnTna
3xi/LLLyal0TFcC/85vIcaIb0/j2bXY7nLCCEHatjHohCe9OZ++jqCsD3o/rolAV
TmtCi4AhCqiBYRLzJRLEMMaGL2Vo+5K2WHtrHpSks/DBE+uwjeckMrdl2jbZA490
2H9QVK3qKYm1JVD2LxMdPky7DQ1t8PKGEoTDD3RZ+0czId2Xzcxp/KvztYfabvIu
CQDliL7GiWg84a3qa7Ya6r24hYNNRpoj7V+HnlBVxJJ3Xi+xTFFwoY9UAVar2nbp
ajfEpsKjveBCsZGlbmOXG3DTpgkHCPeBd4Lq3CZzgzfq+OId2x1o+7CFPOU1xZMP
N6s3IdFZ/TeJcn9CLUpkN8/7tC61XZ8KEW9ff1bzJwHVXU1wwQ7egV9ktpt7fAd3
UbEIcGsVRRmoQ/4alqkRbTf2m72aHFkeCkc5VJTS/U5YjiZk2+8GSUwXfZlE2ORj
+GltxRnvqtFlEememZeG6tpMO8QFEMfvC5p5rhHeuMxLN+ez30aEfwDLx6qq+FCR
s3CdYDHFqIQ/TDYP18ulEtkXQ6vbBYU10G0Lt8Xi832yZ6gr1huPe+5NBL7T0cMs
Dr7l6OLQcH+9BgC1fRIgvtG8tg1Ci6FfHwMn4zouneQv2uCVxNxzMgZYvdvE8iUh
Dugn//PLPrgVz0duk7ZcOT0bfSj4kbje0grZ4adR4kBAtZYmTTQybcxXSo8RDY1G
LX2ES7hiMCvXNr+YvTnvh/338PayVyoeC5vp4vD7X2wbT5nEQ7N6+QZHAoUYp9tU
D2J/DnznwXXt0XIHTQpBqp+SaryKdVW/PK2cavFurb+R7THNJi+MPduUzOXMytpJ
rtIBX9LoZ/9UzH2EOlLMidw+leN51b/pCGRfAdIYL6xKTaLSvF6YZBQOJxH+ZWCp
djrj5BJNkgeQ3bGftWcu8nSqacyNfiLGgH/OZNvQJkmWk5UKMl7bcc/sWDZZ7qH0
rVji97xpc4xIDrtkdsG8NiRDN3frqCcInTIqxrckOgsI8KBCC8sPBE9BuBZ49lDb
ZoCjGZcQRyeotp9QJ07Lg1DGWtvecLBIE45hTDwBCA0b5+5pi4tAuAjhzd0AU10v
0/6xm39p5iPyTW6zVuk0EZmsPEXFtvNINe6Z4ezYyJmxKGvwr68vrY4pDlMwKjZH
zh6INui+iO/b73tzJEGUPxgJ792sMcdG7BCG/x3bS2WuW/0OJBJ1Fa2hXrrqIdoI
c1lk2FCx3BGqvglLaUmA2dAByj8RffC+Fk+CjMImMmCg/n4Dpdv3klNbhnRPTfp2
UV8OiLKi8Zc68+KlAbsSyrfA87+cxmCJpg7E//aczXw7htz2tOisVYYEUQf1kuaB
T4vQD6rJ91NpK3rPihvsJWbvn6I/AJHwV+L3KildkKzNEWsY5zbwTT1YN0ui8ezb
wSOEsG3yZMwb63VTOVMqrti7IIH3Q2FfgqL9kZzgAUWHLFsrV2nQ2WuZBtsqav2I
9NzbT50Q7cva3osfiLusvJ4a0YN5/y3b0ANX7DDb7x/OLIGHEZVLgDADoW5V1wJ+
L0KQsbLvIOEOyHPqY3QK/QTou42bPamYRP4qrQovOM0hgcnyxiJ+2gGmAS6f57hm
pKbG2jVJYCnDQ5fLPpKVryqq0MbxywKFPwrcuh22SUEHp9MTI5oAylTPqv173GXc
PS2v+4CaanfUjBYZdEmjhfVrb5ImUzRV5NjKVCshDGNONgppUEiaZ8jJgQyAf+ns
vBOHKVlN0buf6y9Ol/QN9rHt4RxUCY1kOLhAyL32SgDW/wl6n1D/DolkxFc6iDd+
YB3C5OE3oPxxlQuCVMsQn3Tb5vygw3n2RfNSfqipj0gx0FcS0We6ExqT50pgYKsT
+kPuYL3rvK3pgqc5e0/CUJGv5+eYveRlLQIEER6yvvClr2toocXMJqlW4s0Cm01N
I+kMcMS7+8UlHQUClPxWOfiHzn2+jYh+3OgvuGjhyBNxAqhjJEC6IpijG/XupqK+
I9Is2dc6TUxPIrxkSmn6+oHhnftxLJi8Cby3yT08XftYKQAq/qAsFEheG+HkDHVb
DyuX+PSVse8ox+h8n4PpywHuCpwmiG3Xfza6etRWNhbfmeK0Qe1RhgQSzkHw1c3o
bbaZBgFVO1ZB0YQTxYXlYjKTuR9BRn1qDpN1juQdkflhGvh+jiwEgp8Bc0L3JuD+
K9QbusIevgBLrW0ApdRPcpcAjWKEsx6JXs7U1dgKyoJlS+8flcA6AOuV7MtAsn4Y
h8gqAgNjLAPe6DCOpXrKHKs3b6aNi035RDewyur4bQJaxLCPcavGtW7E412ijh9Q
OcM0r5VUdIXjKr9abodKE/4uHGOmwca67w4ySqjkWI7NUx4zxkXxZ07bKB5QK1Xz
pNk9RLHPIshEcsBrx83usF1sL2KL5fVK0Oy9Zjf3x/I13282mU9QOYT6ooubhoCj
6bEPAj0cL+In41Ckas+CpxaK0X/ax/ggI3Cx9wE/NTNhpeuNceJXOOrVYR7t5rGy
Xz8i/FJBtUjUFIhroP5z8NM3pBvGDDx+EI+ax1lsypbaNp/SeMarEc0TkshCAJrE
88lA3NVwmAAWrgJ4yJC4BN++6d2ao9XMaJ73a0p9sxAD09jQ1j3n+vA+jVEmoamP
ivUAGgvK5uZsbVdKx8EqU7i23JN1r0j3MpGHgymSKC0pwkXJZ3u8zjDH7nsC6nen
U9YGTmOHDsM5GVMcBQCYo7O8n5csi9uiejicuRNBgop+xQzwbsFUibP0p+If83FB
5HqX+J4nSRwJByHBmDa9qgZC1+kUoBDW1uj2BTKvNWypoik1crmLmaCAISuki93p
iT29mR3tNpNc+w5oyjIf8ZnJmIxfHMlHfprd6hZ9mzBYdftZF8i0vZY7gNmLWshP
F+2riKoZXkuPfs0tM1KoKIEtZaSDz+/MNGdBJBV1NY3xodx2iUfWZYc0jw/ERwbR
hFWvmLDn6WkNOky9Y/91pwh/OfM4+wknZ79vup8x1JQ4ndN3WGzOWHxGD7snJ70/
wQsikB1AfZk7odly4ZZhcKeEnoNFBqggC4l+zCPgRHrgAroUcGprq5KPrsOB8LC9
InEtmg36dzO1hAAhTzaa9KsQm4XQ/RstZhIkVxwKfeDSgNz0ftVKPAKbu7MxXUEm
RdwHpLU6gN/xu76uO2Qy2BbEJiMzXYg+2TvtnxjkBTarPrfboM4BhpCzveZ7l06I
/Irod1/9fd7APK0dXyyqPIOO4xLrCBa10IDnB6V2S0deeJZyLyYFFqs5+eLk8IrT
X4wYb462AwGXb7s3tc+eSyCX2Pl1E+33V9qAWWuHdUGrioaQG7DTCyM+9ahTe3WU
hfeBpAUi0prkTuRYCLitIYVIvzgxQfRAvntnYQirSc1grJWADvv5KSg0SHXcdFeX
zgQvTkzUF1wYWQz2gHGMPiUiM+OqNVnsrOiWbfc/14eq7eEMfcmU5GfrVQeHo66G
bbQszDUTwBmJ65ghkvBPPiYdxUU1c0I/1zWqxGQVlyt0M8C177bm/Feq3cE72isg
JTNxKb52n06/CCt9kMhYTwFnB9OrnKLxLY6LmDM5Y+Xt1S1fqA0KAipy/cI/4c6v
K83Zv9cMmiSSsYIWXIgpAbvpF4FK3fzZuCs4aP6l+4cCDViEh0mygZAk04vhjrXJ
PpSxUYZZlWIivwziF9aY0eHHEK+fv7m0qvJsyMKHfhoI7AQ3JyD9odM32/Hoyh4b
U6ZAHQhMachQnxjhvFAxX+a8GfzEmGBOEqxGrajjXV1iona8RqhN+sXugvlPZM2W
ynLiQ7wCxU7CR+6hf1zZlXQP0v5jOItNpyoQ8NSlD3qtKehEcWzWhD8j5Y/v77ur
LZPK7hELibxfeWPDtO2192GixSgnSOo8RYyIFUceZ+H3ycLmG9lHFxn1v+z/93PB
O3afvROXM4eni4WE0wmvkJv7GCC0zxtxziJB8GLcMB6Ans0yAZm7Xeuh2BBIXEOr
ywF2hh4hd5mdrX6/uU6hnA3F9rm0zNXrCwzQEmRqaRC+9IMbMe0jQtifL9yRAnis
ZOWd6aVENNbJGsbzoEee2Gshsjcxj16ywhLDI7fVee8SdYYe2jkkMHmttZJ9hkXE
s1P/NTka9AoCit6xi8tmqHm3LRprmKYuDKJS4DX6PxyxxasjmWXJ2jIu584hdA83
jRSRsUrqH7iQuymQNtWi2ye3XMTcgRbO6KWoYBiWtHBKqgAAjBdzZ9OnCr2srsQF
EHTLKzyYJoo67ST7Jq268ZwlBzG1eqdBEP20G/gy7XwP+4pvXG0m5OsJpQ9hHZYw
Ud9ofP+Nx9CSp3T4n1srmAYGbJmqJ6jNK0pqlqmOB3aZE9oTLQ0EBxslA0umQY+5
TfztSfofZDfXbBV/PuqsxjYakHI1Ul2EDGvjfaXYJ619Mm/kMazG/hfMRzisKTP5
dm+aMd9ZVlplDqU/gAriVrWtfmctNw6a0ve67956BzzhUF5JVENmNHIGkRGcAsce
qmmjmW3/GEbdF/wccURW7DmPExkQEDbQYWcCxhIl7UTw0zohpdA3PC8Jh5+KysGn
bbg+JTXJ398ck4Mg82rpUCBD2CObuH2iHUL+UgB12xajrjZ3MocyWKcGkRaaV+Df
NX2J3bWp+JZxYuNp14LO8AnNo+R7zojvmImslWphEwP7ah7MR6qiQO7tEHnx7XIi
583fVN8xLLgpVuTAEKkHzRlg+G69wQYVG4ELghVYP0Re2yEcKhH3nrZJlv0GM35M
9hHgBfu7NqjML9sTh6gZrbkqib0zEEZ8ebmjDMfEG5W+uIXDJuUouT8RbeQyBaMS
Mga823ggiGSHaU3SJY+yaYgRx5JfQQy8f9rPwJEfuu+O71dijxNeTsDpigPFroo+
sBU5eRJyy0lpn8Tng5/8nl7ZM1iwqoAm0JkbXhggKN5UzUQWN99JPiTvkFvSPDDD
TeR+1qv/RgC0sJtatUrcD36Cmysuou6JH0jLvVNyAE1YgaolwBiTu9Xe6IEYGgQ/
E5VK5eNnOxX45LA+6Kr9L541+RjtJwMHkuFDAFuLP5nVCWQ9v5IZ92RdmiYHQpqw
Aq54rklW8xE5oBSm3qOzhf2V4/fX8J507IjtCr2KqA9BkhOxDdmp/74v4+MIssmg
pOAmDlECWndtuagri8NMPNvjQIl8t8i8HOspi0igcS8833JI3TfqeYj+feSWo80m
7yJoo5j6yCBoAiUArU+/CH/3vv85Sh6CURS8MiL2c7W+gFoaH/IPZMog+9H49TDU
fSBRAjFEmHd71ZWqKUhXnQcQq7JetyLdf0YGu78Ho1Di/XBWKbXPUKCIxh8+PfZq
+NZZrhXdJcEdwllMdym8bPaqNQvw6thu2p4fumzNTWbwJU00eL3naVkaYufqXDNx
rbxo5fB19uJh2Vc3MSxz/WrJtBYzpYULsbybgu26Xf0b8Xjr4z4c0W7E/nxj5X85
XhHw9zBc69cZOWn27IGdMK7j5rrmT0VYYyMre4OvporYO+/Q89wZZNfYBoXyjRFA
7NyuQeDHmkE+2v7xx1HjaPrVAavJobuFpjtEybmP0zyb6iFdB2n0crPj8sOZGsAi
JfC3RrosBKP7mCor2fub0pZepDpDdTttSEL50Gp3yBAfwyC6sKVOObtvNSjJLAqS
36SY1mmSJspd3KbNYiBY44Z1JDtZz1tnXpRgqx424fQ7QqgjAsaufPu3i9pKC3RM
0eKPMigmrPtjarwxhToehI6Gz7gp40LUC2Hf7jpc9JCV3BFFtwN2dN7rKxWiX1XH
Qn7GDK2AEZMNZAkGE3RNZppiTNhzmsPAYGU3vhLFzWJVHZFMp8EYu5XsuBleAJDe
XGgE9EbThLnGArsaRWuYKIgcyGQvdG4V22PG3q44vFcrd6n9Owky/QX+DtH06FOs
9iqfrxYcVhgR59/7mG8mcN9wFLBTSbnNAYIm4XRjNqtuT274CH0MY0/y9NZRriqQ
qfZRRhlvz9dPyvwzE3ZJrpYsHH+laAt1vJLLjbxpf/GoUvnDHi9D/ushlsuctrlz
JcBCK6boqlC+rl0rnvfBRoOybHy8MijUyZ7fqtWqBaioqZg1NISOvOoi8rKyTjax
BW2wy0pk6i3hAxN3QOgM9KAQw0VNYe9kjZNiZZpMFD3GxxhNk+/ymY6ivOJYkCk9
F4Ml5/3Y7DvybkXRMJS1rfHTaiCXZWfEFy6FhwSdIDSrf0q/Ouuwk0PiEjswHeIw
2y51siih5nSozHEaGAglJuNUlQdTNm0tlboZu0xiQOpuNsPQj2QknS4qi+iKrQ8A
Z6gtqiHPmdAXSrkAAKxBINxlzWao++0gUtjPdfAgYvct6urQ5ZW93+PKty1kBcge
NKRpOX4qDQ1D5WYJOZqfPONYNUXBNMBU55U1WjTsPXcGs/LRlpiY3cRsvTYO2YTX
EpjE8KUxlHcG4ZbzRABIbCq3vPfSOhQqzNS1rOdjoawbCl1lLllkwnyojCHZomT2
E99dAcRj4RMUfkAUm2+aiMoxPvoKfsay0e88dugA2nU+ZsUPlGpcjSEoPf1Fol1B
4wNwimdmQIm2U73jRu4GZK3rePzipco+1Zh0Si1UIIXRxzmv5kXa6T559ovc4dkh
+OvMr8SPRjdCRQ1vUUxE7AsG76azE2us9E4D2FplkcPIdW+QffX5iuIwvbwEJt93
f/PoFXsKY2TXqUxTRwSXJBqar1OsSeSi2AdG3lnhyY4tpAXlbYX20OUcD48UF/dv
pKekic8zFZk64dZMVjIrZSUzNZY1RQIQdV74fapR8PLtijyQZ1OQ2rar/w+yG+pk
9wP9wdnUXWhLDDc7j8TQqmXIyVXkCwzxLJYk7ER3anYwtc5jW4Ahh2+UmMVuZrYe
f2FnYs9UyHO58ltxUOCKUPqa8LQ8GgaZ4w7L6hG0Tx4Anpb9xFUEQDL/zyEUVngH
4dQpeS/n4BsqlKVJ2LsKrPV64rrmRFU2d/Du3PJ0+UlvaTluld+FLDVMxtLTzFIw
0nnKy2ah3WrtURRTWr/G5OE1W6eX3J1vGVC1AYxFrjz/lBXfz9aUrFQS1GlxwilY
04pEe+HsW5gd1kADC8sfEerzq1xwbE+499n/dPI5VKGK+3Qu5Y1EAWyazvRZIZg0
oeTInrglCZnRmuvMwFEqEhm5eD8KPhZKhAKQQ/QC4iuf1RMpmEBKcoVwvqHrFfm9
thQbJkjUzz22CtFpN9wel2rRdmxPOANhl6EW6065iIMLlnWNnRir1c2o8Qr955gd
4wQk3ahmze7QLIiK/YsNd94wW1eaZ1LMmQypvT+PzmGCIwToTJtw4kwOYSvP7fTw
LhBhPkU0F3PuKW6HNJp+UrObP9nMo3jjm9ZPy91YZKfD2V4ySsd30xUIXMoFc9S6
Pxj58X93mNMoCanlo1SfkbgQts3Cu6ghaX92O4AdcGi2a6tKzUzybiYOXpLHWg53
GHv4OwwptyHzXZtvhtHm/n4lXwCaXIyLNA29a1o+Tu5i6iml8LqauvYmD8zTtbnJ
9dK1GJiUOx+nqARxJSUcsyl1Bf3F/uWHfzuWf4lQWYyMtYZIZUv1mUB6r079qZQC
dY6TTYtmSfuDdFjUnlpYHG0jDuf/ulmhzQVzNoJtWXQJPFPv/eh4omlGLs10LwCc
3uoPVrbvNFum1ACu187p0vo610eOayYZB8MWqyh1w2+4uXuedBVLz7aC5+YTpuVA
Y2Wnz8ksg8vfbwf3rpqu6uK6K00RGxGexMK5R+rzwtU7KhRN0wSvvAwkQ3dnNop9
2f7argnXVA6pbP2THyp6af8A4iaa6lU+ho+u3t9nwaY1EnGUMUgcok1MQGuJH8sA
brhPyt7kL7LeJAvWXDz3mlZ5Tu1IEgvNe3CSbQJeQXtW35O1VrmBD7XNbYKQma98
x5Cpapj5fSc5LxSjhFo6pG2KwmZURV0oeD5589FiOvIbkVSThbIuyOR0s29j1ZkJ
CVUC3cPuOXM+7foaY3mV/D/3zMnZ7vvwIaiejDzS24v+gwUQgNhLCQPo9CfxccRd
4Ow8TN0PO/Sr9XSzaUMYOeV7AFlYdUoaWzuH4WLRFxWv1VAkoNekS0sMQGeiBzkU
yByUsYgrToC4Pjov6VsY6P75+O9VwyvJgYSdI1+yomazaNfBz7d+YEjESx5XADVl
1Avcew/4KvAQ+ckoJ/j0Hd/YNuPizy+ncprUV/0WIOACR7XA9v19wNrydbTCE27S
HkvI6MlLfT4IOfZeSY/jI/swpmq8PUZR3Xl44Df90FldJlGaoRpkZD30Sw0299iD
f0SLE764AZzzfQ7xbFtRzL0wfS1VJ960HLKL25poDI+g3Lzt1rddAXcjJKp+htDE
ilUVCDgiVWKh4/DuE6g9xK06C1z3daDiHYcUDNz8dWPxH/lEGfTaFi6wQ3YBjIyx
RhnJpZrlA4jx+RyUr4zhL/s7QlFJOWj7lzDxD/NOBrsPi7Agd1Y/smwAVLvkJuNX
41d2sOmCTwBdVJxYy5vIDJfODrcJh8/8sUIZhc+vlAtL84iL88cbkGeV13UpSDSN
UDoA+c73dV/poT9YoIOwJJRzyE6XfZh9XtMcxWVI6mMACyy9L6VDNlGCJEmwo7wZ
HnJj52AFzbE/GWUMWow6lSrwnIFDa9S2iBy9DdfjBomfozV+vF7/ofuosJX46Wdr
ejEpVCOjVEH8frlh1Ww1cggvvTe5jsHfw5Nn1sVdR5lx/PEwkj1fpP5gxMHEDH/w
DBLa4HwHJmUVhxYMK8dBhW0FM+bJtsHGsNkZj8Ccn3bhamRQUB2tLFsks5wpF9kA
Y1PqlOhLPskNPRlgm6SWoIzWb2aHmdLoxPngo4fz/i2DhXgLF2Bnl8omChTda/vO
43rBigD+9Ig5/iAMiAimyKkCoJcMaSuq94cMd/sOycxrtkMVY3YFQIpO/1dXAmza
ftMGYQ+LwDw8v0bE+wjscGO4lcRg0LFANijlaqi9xTJ6lFUL4PlJo8R+WT0EsgEq
TomOjDPITP9nS0EaKCrDdau89h2pEdwLCi0etaUa2DiagGX0/k1X7z31mGPZczw4
kAVcAFikeLXxyq78CQMh4Wj35LivNIuxNwnbNCxnPLs+B0pooy6eVjZNHjHYI+Cu
qMQ/7dk7xW7hyFLXeJz/Us9RWpSLenG92Bw5pU6TEgI+54SyLOoLSueM4KFJ/XgH
SZXccMpRu/72wK5N+A0jxTDTVJQqDqxJK80/ZohUmoXcb/0vto/tcZvd5ojkceHK
ME5bpWlcKag8s4tcUylR+TDX5GPbwKgfK4rT/AHQLmq8DwPPkG9LTalh6SYBsEAt
wi342pAVDbDtanNBNpbaad1EyILZAi5xgtSyxdH19smi53cAVm9NV+n6WYp8oAbN
cj8WCTnrEonf9VjHolwgHidmICC3mCa8f/AAfB49Dw+xMKjAqa2zj+BFW/PCmVCd
NlFp50UOYr/53BLHCFBMSKTVK53vXGJmDIbqmWtTiBNAgK66XIT6l1/SsBYXHy8h
QFUYx5IscR2pw7jI+96SpqYAWXxgLoZPauTH1KwcNEN2ldmfrAfKcfHMP3BnXAXB
EELAnv++Gs3HijCui0sDUfpY+bX68Q9TKaB1CLkOT6hRrsdhVc0AHJh1HrVcu4c0
SmL4hfxRUjD2YmKEi8SiTkDQIko4vqQTXnQt45OV63IMB96unv/gKVWUINrmbXmM
39fn6TPzdHwzZD3JHMtqYHavqiVKu8yGxD1ev2ZuiFBKWBCeGYjOBr+0D70pNoee
Q3zIBBmDE6oAXFC1pWZ3DHLsNcNRBzs8iRufCRGVOGrKxDMRS1EoF+4gld4Yi05g
jp0JRRQxGHi+jnOsRN1JvS16WaBFaQo/DJMrdULDB/x8uwq3GtbXZ0ZUwF0Cd1lx
hjAr2kho+eqZQqDNL+T+P6JZdhoQFcWPl7QImPdJTzCsJ9ut8U2urmiuv0fJ2bxu
pLDHIjBe5j3ndcQ68SBe/KO8FeVG81RzmMC6boZjGQKiwtN0D62mcmHUOeAvBDnQ
lLyXoQrKE+jNn6WPrl8EpX0OmqaEdnflZ0rDNtegk3SmUIZz//LxxhrKm5/+zh2m
SVQ0LGEK/Elf/1HA/ji+xR4awc17q5uMt2oOMMCPUo8tPskK4Zos3Rb6lEeRJcqm
JXlfMRxGOTEuVpS/e/u/YNIgocQWJ46oK3hFRsI8Xya+IKdWOLfmot3FEfG0kpZr
9lY9EvX6zMmujrWYnIvDaq3W2eNH0lleeZz1+QoHEzTErSVNE8N1WrTsLyWfqCi9
cYpb3eAy3EyZPT5/rz0PFW5oVcrJhOuuSzydja2eOcsvSyd3ZXjzzQonLWcbadhi
35pctn2gIwCr1VQgQlhih69LR327KvL8e/LfyqpUzGKfGlAf4EiVHgVvYFutSNLB
kSP17+QXywfXpVT9U7wUgsVecddYl3hgATZK5eldrZ4taG4k10ZRy6oOKnPk3Jdv
jQrW5FvgwYrWWpG99nKin4oi6EB3RYLd+dizKyKB4L6cmpdgfCbUgSW+mn1VNTIj
0Qu4grkVIMZulyqlznX8/WNlkzQNJflGgkp1pavjAfgKRpGFU6IL9QxElNQCudnw
Niw8eMf/swTBOLcwZWGjuhDiFJPNk99p6hIxMS/h0FexzoJHijHk92CMliZtTOfI
lS1eISQ4jFeqQ6CnRrY+EcXdlo0gh1A6ZEUkHYBHj+umy/UKfSN6Fq0utvcuww6d
tfyCmvLirNj2CYXzwD/7uwIBRku2hUP1JCCDwFylmk16q8kwWWOLA8Y9SbPca1Nr
UUA25M9OgdSTb2Nao/c+NrbPeNHW4hNMkMNVDryx7CD10j0eHm5m9Gj150T/Suwc
FNx2Ud1GNfwVf6E8J1sf17AKUhGRxeUwaR0FeiQjuyLNf3Pe03fgsWzvEJFQnots
+cAyIGXcmIlYBmZ6FgQQ9o6FHkDjiHKtSFFVjG8dWZlk7V5CkFUycAgVWojUWnlw
1IEa05dTH892IhQzXoEcMIKd2qGOVO3M4y97G+7k8P3E/5b/KAxcXFaoNB9cSnle
LF6v98+r4lNuM2Oz2sqiVaM5KlKsxvqshsbiVBmgUFGkuWHrmWfueimo3yndUVAW
BjRN2WguTdjBa/loLoni/bVZ5MX0zUBK+1YG1HDi7+d5rZeofylkAKk92mwltDEJ
tg7jKtFhQCWzAuJYrm+a96f/5QPV+VGJZGMQSdy+GACERz3scNhSqR3xG5kmJZsj
NO5aRhK8eVQdfDCk+ty/ApDm6cBM8D19UZzSQRoVyCXsmyWGbXA2IV3T274RbseA
slOX9uPkIsX6TCS7UkqizhCxfNriBlavjQZKg4gqXenIQBKYOWgCYBrvUXADBJgS
ROeIs1rS7+hnAr1VtD6yf80lkDJc785KC9w6nf2z8dFdR77N/n1wpExN2M/hjKvA
M5DjI0EY7YW9+veuwWlF6buxZUrltQBbtloB7+N/bqc0dtiuhZ3V52ARMCHzBonC
Gsa+Mh50DGq5IADyig7QFNWOwuL3cqppc3KANtYk1TKsq4nG7N15+v/7J8fBYzUb
fXVqR7bjsg/rcxzYyNWnCCqMgunSu8z7J6QYtFahcIOi9cj4A1+YF1XVqOPGfvXY
8kPeyU+jmV3GEfo85CA4NPPiMvjNKBGkfFammly4dpdE4RUa9NlUq8E6GEgB3V4i
2K+ZjkCCNCn4u9OMCaRHRxUhaZYLDvlYz0NozG/eZFANWeDUrXwshTTSC2bkAJvo
CW5/TuA01pa+54prlVyM1K+h7454EH8xAP1/ICauFjS+4ODsXerkY6jF1o5wb39p
oVvBdaBJve5SmyRyMaAq44dn81m1cqi3UlLhjJJH05E5+fUU5BnoD4Tx1vOGmFWZ
3ihPrr+P/NUnS3c2VfYpsbuJMnF+9BzLDrdAinSAXR2+Dg9ORyepoUTwCkqnjC6b
mhbPWGwkQO++ZyxZiLvjozlMTJKG1iVCxo4H9Iw9LRS97eOSCJQp3rwX3LBatZ53
vxBxsUOYafjJkMpPgSfR+f9/M4zUI+fwZgtsedpKCQLU4UVouQQZd8pUCHNnEmwB
ifZ2vhdW7pbALqU+RNOwC2PBw8IS0DX1TGNA5vtFNi6aQQejgsRfeTZkX3UOfXdm
2w9f/l4V5mxJXtyRarNFMQ5u8ZZxXBEw2WlB0A2RIjq1bbRqHTwbG8K1C951BMl1
kYYrmpP0+iGh3uaffjlRSfsbAPjgg4kuW1n3+QhyY1dKR7aBi5L9zY1xPVDKaF12
M1ynihsvRk6gxK1dewI4dKx0vR//PqCSWsyhlyfNDjEFhUX7GOVIsmInLLd6A9eZ
XmyYTYOVgP70Fh78pQzQos78CHHjTHsgzZEdBlOjuUtuAYMBqWxinD/2xV8n7SYE
FjIWWJbEXqCDFVpYniZwVPsK64xBPHNjw928MRN+VGxtFsXVjFTDcOXhl3g+3Ysn
S6Vcdk05g53vvfzbRFGKtY5aThB2gZzAjZyUddMuZq64ZmvZTzua0VDyx33vO/RN
SFSnTDyFpLn+9hj8+iRVlFUvm+f0t7LU4xII/ONfizkEOU+dX2gqd6HF4tv1A/v7
nf2q++eWCITfTluG4Ig9CLUef5gb9wQdsxvmZZqDb+rBylqBstqngOXhIq+EmF4t
6rsGiSeTSbklJwgneklYBHQpiF4wZ8Hw3e178kv0vbUYzcDdV+Z1DAPCamO7kzcq
FOvTgcS4vq/Gwjk8crSEl/vJXH1r3e5L0U+oo0eni6GvQyrX9gA09YBA7GpZ7rpH
UYTiWErmt2fziDAihptQgC/lLkCdpERFm5ne6tUL4pG8fjS7tLFzTV/T2v3RE1Dw
AgxNYNsXmK5trPRQAuwBPdfW6DLSZ/4gbldFMgb2OdJxT2aSY+s2lhgY7v15j6nC
iS4BjlDvkp42xClM8lMm0NH8C3Fuovk33GDzjud2+Jj3cRzRCYQDfbqglFLXtfUO
6bKa2cf4SUXSw6g4/UBzC9PYdMq3BOFE00A8aDHVtyHTLIXKxG74H0j3R5R8b+sY
Jr4B1w+OLEUgASs2mkx9+OK1GhGuMVyIaUc5baEPM+y7HF4erBOrH5BduhlkaGdO
pMssbpXuZWNBIIlmsqJhhvin//UqDBt5/tg+0kPEDb01utYtxN5aFl2Obu/ZGCoB
Z5R4TRbdOnGP80cfeePbJw/oAlvkPNZWjrxg/myQzNAosu+TtCvfkWYCj2O88jeH
siq0JpY+St+6eme+vzAsxgE4noG/7kkEwKpkxC+2uhv39qEGAcBU4LgHKA4Mqk0j
uv+jnu316MGAV6C49mrxnBuySGiESP3fUn41akQYsvnh2fPLdCKK73oceLcLzwvZ
fZ1Og0/7TxLHvocE1Yo1EHBp4M/nNh13gLL5l+LWMIs2DGsuFaMYvQ7uZtYrIwcf
sXXrKeX0goPfa6ngCVpzFNSbQ/QExzItTox0x/Dt+6ABuHv0ZuV4FLED9AHwnmOQ
AOAAs94QVD68m12zPiiH8TQJB2BG++ieNudfPUaD8DY4RZrvLDXozZ01I9f7+Xks
q/rJ11UvJsOzchW7O6puaeeS1B1KmdSf3qCnrsYTiZweKm9ntEJD7u339MQ4Y9nV
G9sAMxF2ppk4Od/BdeKkmdOTdPuBsB3mjCBDvJ5ZXiQkeu7fKY73Hyc3BTSJTc4k
mpN3SJlwuwERs3PBAGAdzwdQEN1QegM0ucCMLdf70edFvsClFMLEIU51ENsCIdC8
l92RoFPuj0Wag8aXKmy+ACFiqRtulYw2ntgUuIn+SebvkJCcZIzivULI/QHxt+qN
unw7LHBSyD0c0JH9mln6PXI8nWsF6uY/q3l2Rz/ietNtvA1qvH3mOHBbKSxZoRRC
e1gxtl4qinrVFewSCW8LX6zG7BJ37qhEokPlWKFxb6N6B+bWmSHmiWjEqSJG/pFp
d8RUgZ6bnytAIwX848D1PzhZRaUGxOH7z0rV6ag/gr6GkzE5K5asr2DxXJaUGg1o
E7E+92NtN4mAXi44aCuftFI4sAMZlUWhNtQ0d8EcoaGWanqD3ANBIDY6TLIKG/OT
8JW0qiUobbI4oWAj5mIe7m3Venja0R3WGH+MIXzNHJFNADTyT8TlhAAHvCzGFXi/
kErnXDKRWxoE9UDeg1MtztcTilFC0j+YuQ3d9LSrt4CA7dB59BYAY8n3haVXujtL
j1ZultiHoem+9qm1gCwwUbQVuWjEh9D08kWHDx+1UfemEFogHfJIFdBtGdDng36e
LcZCr6rPI7HUJOlXqbi/EgvKR4hn5gJnXEE/h8hdB2x5X3S6sd5ScSZygtO+pVH1
k/Jg4Zr+Dvm15X9UiASbA320u8P6bL9Ale8oJNfyMN9T/3Sp47B3k6F5KwM7SvQ0
dl20u45vpIS4PFMxVSmRYitLCAOKyDF7sLmyFgK9SOfJRPl1EgFnlld8IFwenRCT
WnxkvRVUx8re3p4ItgrmoW7JAj1qAfhTgfKxxeiuLwrbrMN7DhCyW33q6HGWeMYD
+eULdxn7chppKyjUTAF0ZW9Tect1Rw4MaI2tq3+Kxo7j83jCAv2i/iWL0gMq30vx
WEFEPs7K1AO1lprmo9vzizRHPsLoC8oq65gHwig5qg+GsgVxNGXvaGi+LqGvBpYr
UIUxZXEFyZ7wTEOqSX9qXMJap9d7L1iPWhHhj1/dEGM97UpUOwGeOKXRCGpbVjn4
Bm7eO3RJ/kzN+b4DnJmck6oValPTAzzAT1ivsUyBob/BCOy0hVkURLpxhoEshK4K
Jb1MgIyGMrgoA9vV7pZXn+slZd3CRsWkBDymzMxRvbrsz7lMscQPlqYHU+FtlEYI
RJDBwxXj51WdKEfnd4CqCcfO2kfOklyuIpP7lWzu6uVPzqwwc6ST4C1lVzSnAGsP
JotXo0eyXKFfsOOze1mjbG9YqDoTC0U6hcvdIim6mJ8Smtcp6UXit3MbCbcAjEsI
jO1K1Jg6hUloE1msjOuUNtQ02i0rovSo9cLzXT0/2R7CVuGNYpi6j1lapjiMmTBC
pG1bpf7+pS33/jsmfOpoghStjnnVRFRxRmonenGhJrd47bVL2hPff6wAqNPBhNHr
6vCgkRp1Hreez+2vbLhodfNjoTAMCqaajlCo9jzBTvvDsDBzeKhuRkU3J874RlOc
d5Vdw0AT8jtY9fvPVW8wO6A676qBa6iN+P+KxRHydnkybYfaUYoZ6Gw0mleM3EpF
MHOmvmSBAJQyFdylvEGdsrdFO1V9SwZz4j0lMrnSmapVo8fxSsBEVDxVsNkeBEGD
B2FB/rSPN5KqYM9a/N4VBaALVmr9eKFHGm9KKlkVrVfxjdXCjNzD7etg72nsMzl+
c5hvH/FR5SrmKFE5sz18QiFU9uLzi1zIDFoEJ3tT78MOFTViDVMpFL3Ig2CJUsb7
yCb/IiYtyiTaMgTVnV9e/7bqfCgPzGc6w9qC7m4UkXgFhEXvLa4zsuCO9ZZ2VRdb
bOE2A5uVFTKAov9pjizZpBvJdbZIDuWoA50bE/QONe6uBO5fMNUVrqknS3R26nan
i8P2ces0Eai0p4ok1JKFP7wSf1z8PDq0SkjacFiYmaSZXrwNiN8lp2L066Jub9bU
h2debzZ7VVGO3XBN8ji8cVJTvoxVCqbdLQCen6bi0XjtVIB107lT4OmijtxuZ1wm
BXWWccXyhFQGMAq/rITSgVdvXVEnxeTmkpnx1No4ZB8OS+9MxMq6DyaUV123JBGA
bqWGTGa+5iTy/jGkxZWwKnHSY1XBVGKYJGR1VGP7KPMDfC5pOZ91+pfQ4WO+GJWI
o8kmYz5WBNsK4WF0guUgfgRWvIy42t9cS9et2/xhW+Fw0ALaTbpd11/XnZwhA66u
O5HyhH4kKw0WDVQgsQbuRScpL63hBKfFdZ3hnWwqAWe5lnwp9PqysRVBITLidFQ8
VDzlmtfqX+ptuQyrs5Cbv2PNaI8DzM6wFw3wI6dLO5mbs3dsO8Wng2rjJE1LRQD7
7Z8o/9Nosuib3sR2s0rgQWqM4h+ecyhcatdY8OSSx7yLGspPXn3TnKOL3vQs5H6p
dmNa3b2iIQJbFKuYKBaqykgzvxED/tyXC3UFk0c3GHNWiu4AhKkJVg/dxUUu8xEn
DdPqCPB8k+V8vUEbiDIaYeAgFkCWhu84+HZG8AtIB+rjy3DDkltlvzGPg+DBbyVJ
5RNkJoy/hypxPP4U/HTM2D9yrVHqWJ78ojguX+ikdV7MvMFMdfr7qY1miOYuiAEk
puVXHZjpxxYJ6K2rOsjJWyxoVnXbEqmSTtVQUlk+vTPvfoYY34pJfu24j0lR+AMH
C5ajnLsmwS56+HjvQ6Qh6pP1rtWq3q6nAEygSErObWFVZAhNVl/xKiRxLGOo0ntR
lTgC8pu7PyppUyYyx8BDhrTVfAX+mwNMRkFowez2+J3X382aOcmWF7a3z3QcB/VQ
USCzapDJO4VFetJKML2BFWGROGYShQ+y6Ahyvs20mhpVWNYPj0IGgrS3nFSiMTYQ
ITePfKpafT7WUd0PDs7AfPIGnHu3MFqO8t7YUvw+EWq2hlWOfjlitHqNy3w9Wu1V
9Nula0ugH3d9oQ3UM0ZRLgrGPML46xh26WktEeyHaob1P0HsfKfVONFbE84bYghk
hXw3ApGW1DWN2YgOJpT5bRAYqhzhQMEVLSPUHoRkzT+UnH37vOoUlya3MC8bnhyz
/bcpfnmvCrPWp2tAioTwlpLwnAttP+pQOPBxjHf/6PJkRMkTsvwVXapOYv6hvr9w
w/c9A1xddIDs6s3dDcTNhvRQ5NtKpRWg7d3Ozl1SwJF8tPoP5kOFt0gCA9r0yhre
F5zer7O2tDsQAixLMxlSOy7gOn9U2BJPBV2V/WgBCUh6Pu2EehgChtc0LHPIfMpa
lmf16RswNzxD0uYmicigf2GAEUYEvngLvIGtde13Ue7O1sugpoj1Eog3Kk0REV6R
XGFvogJAxZWuSBc9gz2GZWFSn2RJVcW99myhoM7jUcg+bRljRVNKQUXagb2r+QAh
f9yNDudX0uBEaf/81pXPPlotWrisS6/a5x3r2xwaiEb4b3FbEnB1lmlVAhGvBukv
b4K5kbXdmtUvQCkOkWbPQfXqiBpJj9ccBLj0Y5lVf8GjCQQJ8XJq4Z70ERH4sOqi
ZIkdy+MBQL3MO/LsADC1k/qVpjdsnE1UaorblkqZk9DmPV9CFMNnToFWCiEVYQUv
W1zgCrRJWGFbrtv8YiXSDkhwg7ILfXOQkJdm1IMT2tjyNjiKmM8p9KxFimMitIiH
w4IADP0Eq0Wew8MdzxLV+JyTLCiNYlnjc6xry1TCNMOB+a7kcN32Wdfzu4l4dRDo
z8Hh6yF9lsO9uvRuXIRz6qNrZpO3TKPcmVNAxhfk+Jn5yWg7MPDUZ5oqbdX4Irdp
Vv+8ZodC9EKP9nTDOTDFNf/H9CCyZaTzfVBAeSMN76QdV0aP/Bn9+qKJbHINl2SA
CienafdVujaLvlkRyXR9o7uaO7ebi59iNgs9R38Vk9MJg5zaxVfZ2UuE3byQRd/E
n+Onf5kuZWceekZyxlChcOUSbVvDUZKkWDs0UwzoZfXyBEdyGuSTzFpzjxIdIEvh
A69tS01/79Ta9pQ6O8fPh5lsRSTWzOftBCmoicc4dAc0naq9xEO7Ttzly+odZqKf
Se2aRDaf3Ohv5hj61qP0rVcfj8Km1ObwKGmf+/3Qt/01c6iMCqN2oH4Bv7fUJSqR
VJbtYad2BeQfcM8JqXuyPv7VJw+txNo27l2PispqT0l38rt+w2IdhYMN78j+jWLl
QGwbhUdeCvF7cVzVM66fqmQ2WDZldTtfd45O6Zzv/3+UvJzD7TKMtbVqZm8QBN73
2SqKs+P7b/lFi37UiZAvKVjouJCWpnhkrYsXTWAofeFYKVeMj99frB9wJ4M7jRBt
A53twmYmAcOHG650qaT10J4ac7LM+9kh2OBb8Hd2q644Zf9SJVMRovhyuEazNPQh
hUXZ0DIp4hDZXVnH4sPpDlQ9+vdUxqnmJcCJSgCpjXofr1JJpPFf+6Sf/Zdi6o6z
bMnpPNz+G+EBnrJPNuYb+VievOpUtvYMq6mYE5Rc8rIIMN7wAFmsLrwPn8UhDKEL
6T2StZbSQnPNZnfQ9ijzYlQu49PNaC2kEjm0+c6LM8tMqQ5SOUzxOZXiildLiK0s
PGMMrsYsuVM/jRZ+PHBj8sU/efOZWyUYRVzpoduNPz/Ndg1trGZJnA2vShoC2+gU
1ITZMid4q/2XL+oU7SXHc+bN2qTb+vFt6zvW14kcilvPKY/pdWSTuke2QB3Jh9GT
qbiiwqBzsi8QnpruTMJqwUK8DgNuGS+UnDY7DjkGIK3gUPjsUbnTG5+n7K1L7K5D
jdFJoiwRlmhRihwbM9O1IR9uFzhbyY6erftZDbB+L8EgeQQTODcvptDiKfr6+sdo
S8sNS1fdv4miBFuqCiMO5WZXCIMocwR6De78wt6P2KucIQzUjIZqjmNbURF1tsqQ
2Og8rVO+wfQEnlfSjeiy+EzOItCWsLhid6Sv4AXmTckEKBRDpC3zpa6dCF670uMi
3vLK7QYMEm6zsIdTBag7aGnwi++o9RbkQa1ji2ON9LV/szEZj3ii0jCtHqe516Sg
eI9Wc1peksmF0Zwnk1u4cpK+4ZPCwjI/WSFFPxJ5CnaMo1+ORmqklxOseRB3Min7
ZKKeiDyu9u4W50yyfVui29mCw9FMemoNNAtveQsiu/EvK7oxUmMPK3uiLBqjPGqo
I2Z05zpiM42MI/fn1vohEqE/HoIDOC9SMPI7HouzMVSYAX8ERhpo5Lgt/Lbf9iAX
7F5ZMwoBNANCmKrE4Vs9zkn68noLyR/aLuAEU/oZfiqWPfwEvmo/m0riUFMD+UB7
OpbSjF5ib49vYhujXCq0BTFfniy9hcLZ0Xc4GcV/vzFl66aOguXSzZxCsoasRk4o
cccmi+rxkqQ7tlrbJ96rZDKXAD/kpyvg2qmCyHSgsHYTcCfp0ZPM3k5eMKxnf7UO
tmEH+TSSapel0pIKyN6BwNAPngSg6gHbzjd+Ulx7jwPCN16LfVBw1TRL2w3H2Yhc
bhNq8R9uekf3yL5EGomh2UzxxDAgLbpJrdhEzuLTFFrceAC0BH+wy36JdRVLD0ih
MHMTNNL74DmnONZU3/E9lrEU+deoes4kfyRAA/qZbGzM/tCwfg4vSYEF/0+gmwym
BEKEQoL0DM9Oj/h454OWwmpKFo/4aX0GODhcjQNsCxVL4NnIvNyDCKmY9DuKEhLc
1mStfdd2uoRYRjlQwzWzgimCb/0c80gEZPgwZvv1K4jay3FvGgtcRvGfQ0ZL0qyH
SK6TFslSRmVbpCADduNLI/CM731SaG4X2TEtzMnetoddIR2Fg4MV46SJ8WAHjMl1
h+Xwg0Q0nKbOcTrFi5PphTCFDNMLLuCoo8cekmAVr3yXgPuQ4TyIUvTdJFJ/peJs
Pu7LBNmf8bhwCd3oWLga5SFtBrASFZYTCDUBDH/8bX8nTRP+drQtZN0wu184Ppvt
2XUnNobwtsycXk0HvZpAV7uwaZxMljpb74RbqT9X/UlhlS4jYarZacf9ECWjJG2x
0niFHEy8nxlffq9jQLjU4lowOPhOJHUqlppvvhkRnQ+ybyOHq44uMyZ4CqLLXwEr
/BIAps+6hunpaMwuaHXNoAKCgpmSEwd5CNX9kAGFg1iYDXmW48kbc+vYdPX7ENBt
rvRQ4HerOuacZkdYPSK4GhYcPj+z/t29ntAuoc6LH9QAn6pe6Tkg/TRAVClDq2Qr
f6il/2YtmKQ9aWraummbXyJPMAkXb1tsZ1SnWUDS1/f9eQV6LTaZFmsRvOswiPJq
1qwpD1OofCWczd1n6EJidQyglfDcewcqK+m8VBJc9w1/zKvvTISdWpYSzFi2CEHe
mXFycYNVd8lWCAImywoe4OtsUgaNbj/Zh8KmjitY5EFWjvqZSieTAEOwyjw9hE1x
C/eJ79vLYCReNFGHR8/FwgUY1lxfr8LlbO2D/HsC3pqsZCGe7ooc7/09hEp9Ump8
+xthJw2YZ9fi3onkpdorN6NsmgVhYQRleS46HpGBzZ0DlbOUt4Ae3WyUTa9HNKbe
1PSsvvU0fxLKkgZfNi4+0uJjeVqUSUCkIyNX/n8HLOMigzg0jbyhzzCkk90aiUUR
DyWD0cSc3cUaxiwQG+yQi4WZXfLjsZxnRbqB3AOmbIorOoYNCmpFopv/KILR562F
2rrIhlbyuiqt8Pyc0un7WVCL9lI8hJp76w1KLxvocEVnVzg9HLBsu+jMT0aIyxjJ
B8HlN4dsSf2+AzKZW+OieuQ2Xvh4h9PTb/VooW5V7M0R5xgAnGicPFCE+JLb6Wae
OL7SJFXdjcxBrCkXqGqeE002L6Ez5k3KivyUcHcCuU8hYW+jeojb6/C1OJtixQm6
uOx1SYkCpyi3R4v2hijUJGJuNhVl17uSYGgA3yYVdrkrlZNWYg1GDkV7hwCFZMgG
SZmRwqFko/2AeVB6jA0qHSDf1eESBfUIXclCMhUWHb3kJLvz/OwJ2QIqABeamF98
L2WbTonIp7ICaMiYZ6f/tKrfcFzaog4I3WTiFg9zzZt6vdnpEPhm87uW6fuMWZc/
uHAE/58yLOmUJ/jOF2liaYwra9f2gCXHdYXpow7OtwcdnBkU/6lQyBi5tcmJopM/
2O9fUhueAUFdWi1xiI07T5u7rBpp+Y4/7XeAgP7gzdj9V/n9KMu9tsWRdWKq2npe
+PmU9rwsa9lq+n8kXrEN7+yOKf2yNdjbpz/V9Qg/lMgTpqKexmtVvx8DN4O4fnoD
8MfnteK6s/2dOsRhN0jiJ4WDdDemDXHiZ9f/W1eF2dZZCNSQ9wy+2fO4fplbHZJA
Z8dZ8Akjw8i44LJKhgpoPrIxBZPAJf+LKOT7FgF6TFmIXRmf2tQyxNP5hSGrp638
Qc3fSgk8XPkh0LuFEJrNCJ+7aHkkIIibTq9fScIFJy46EjyLX9JMGeCbXonIZtIC
DtA2qXEJSgjKKgXV/5bIqAkuPSd2teOCzYCWDAzaE855j5wqydMR/xJc11Nh1blq
CJr78hx1ukSUJb90449KLZ5jm+WN1LFG859oMePH+2dsL4GHanHSFS7h3Rxp23l5
hzeHw5yNjCPvjbFB+6wacTRt3A81EIkBjoSbsTNMQLE2JkZjgOR/43QlVDzBjELC
xfvVvHQ/Trn1eqlaeq3Owa1P01DSi0B30WUrxSV4rRk6/Y4MUvO3UtuYOuG6xFW3
rKUcbxRFCPfoB25aipYMM7Xvs0I3ZnQcs9EOaLnqB81Ui6PTdN8AAye6D8JTkstA
f+NrjpkcD+Vz+vc6Bac4RfhfkjUlWvbJjT7rRdecBt4pK1+UFaf6jlFlzMkA5P4x
XjJaZBGgJMBU0dkwsSA6jV5u95vXYSV5mkl8lEQBb1fq4akpjGlRBtZ5S+2/PoxY
zPlzCcfcQobSTM4CVEWDay8/zcrQoh0ki81mTql4+Mo82SsQJKyIOydv24YA3xAG
4qLb1JUsgqUdiWy4H6TZBCHocIOaYYsudA0I+jreqlGqxHAFIQZTcaCYDCt8zwn+
ZHYIo7jSM5nzS9ZAcrSXei8jIWmarud47+enb6ELjxu81AHdL8QMH2MLqHDDXj4n
4I2xRyQBet7sjbecCHVDls08dpHQYOljQ75TSjjW5HoTWGfCEWOAuDp0sRPrldeD
rx0rZfFbI+BtCEwy8nUJrR8M1fMqZqJtUTp0f2mnpLda9WQ4Tn7tVlMA0pu/XkgZ
2VL3wLcvFyIrAxu0A3qfWvRfa1s6ihcXUXayn72Q8VfVUagMR2RPMqI/w7aqu+7l
ykh6R72APWj2EkaCPNwVAFwlhkeGkkwNOmM+B0Mz1yj95v3oNRRESCnqujjVd2Lp
Y9CReD5bwMc342D1vW9DA/muOR2OTpc+S9LGoJqXjInDPGjBS+NUaXKP2bTCzUFo
97M60mt1pMhk8PaYXz0vngcWbgYtQTanzWnb6CGWRqmIO7rH9XUcduEGvQJSk0mu
VM9gFmhwA2ZFhlgihmBb1asx+Uc1B+ePggpSTwxqrn7wUb2XA4VTlPdMOT/7kXGh
S5dqjPTU0Ubzc9LxaFf5KoJoS1hWDlVYk9H7wOznoMfCxhoqTtKjbIKr91yELvuH
P4D2KGo3en3cEutPJzaTpDnXI5yARETZFrB3V36SNVhth3v3RRFF4UUEERvCKu5w
siUdydUlsOHj4RobfYTZ6WzxsK8qSzLsPMIQTI5jzWLgeppffivWxqnSMlPYuSiL
hLev9+B6+mfVRmeEcK7fGGX1anSdobgngxEHeTYwI5GtvnbGAbcyDMxKOXKU/vAC
wMFwRMdtu6lgGL3HziHBgMQxFA2Nh+lPskDk6MlulaprME7ttO11+ihw0MfhcoJE
DOM7r6e9xzKoChUuS7sBp1CamhQ/VGWI16nQQsjcfYZMIIkYiMY4+zbSE4Y/rJaF
5jpRP8egzNyxfbjoFcts4MBLIGrDa305y2OUOGLGTt1dm9kQgnwTtxJ5FZnBEH/0
iBj4hJLobb8tVTgeh167EOI0Ir5K6H9ZxZppDnZNY2LMKoAgbInANW6ZJvf1nv7u
I42opOh0iaPYUFPuanXU0OylHSdP5rC8DKTKBgdi4RnQRrCx/BPbQnUpx/bw0kCW
yygdku7hOySXfkrMtuHqeMw+5O03iXXCBKLnE6UPN1vJF4i4h9Zf/Kyu3JKGip7W
PAcQtrQw7LzV5XZ/Vptl4x0C6kV6iAY+FGUkw9L7bXCdDqY5ri6ESLuoHDiSaX4e
WT9Tv7Sv9fpusCtFi0OtaunGUwcAIUhRGGwk5X+KGHnP+vpKIzeXnk0ih5Hg6otZ
zLzYJmeBGKXfSDkBD4k6yjy52UoQVft0SL1e8SpIl03avor5HTbpR60NGf8aw/LS
Mq0L9GwxZv9XKPK4QkECXtVDuQraR5Aw2H3D/cnoA1nf1zTsKqz0rw0zYxBtLjzu
/wrut7wUkchnKwCagWcOjnixTMdq7o30doSxGodWfqTUBhFwBO4aiQ7kPGSLsuUw
6GxJ1IraK99xfDbzXHCBR/fPKPxwv/4rJ+7BhxiTeg5UdOVrRKq7UdoY2Hy0hJdD
0Wa5YIfyIr1iPk2pA5leqXAUHHG+0Zb88xXsp7v2CGStrC7fG/xqvQ9B2cXQdHZe
zjIE1PWxwWDx0n//DNaIENFPqoW6s+QPOPSaWU6zlp1hNquW//u+AC6Rk3qVZ1BI
B+z24rKTOzlFyZK1Eut3N7oYq2gNhvRz6NDnAMZLK/izdjfNXolwmxGZemA89ebg
2KHE7Fl9GW5m7/i17O0jx/0+gDfYj7v2SSCTvDm3rRCsUnh8Do/7aLmy6muUcqJw
zdIthHg7WT8V9pMy5UwWprk5R58UiO5HyN8HxlFgFn18TXwEXRrlWuoMMgwJ8DXF
Vc4vXP3mHlsAiE3LJGYZyLCRSL2vu/P9iP14hPU3zM6R6+OKzSTZCrjG4tXNJCEW
HWmO6I8LG8SFyibsF+U6Wt/CZoCm6JMVEMUuPooIzqI9W+z7XLyoZ5DiR2nOXifV
pexODSGWQjmlou+17yHvfBpEgIUIVUGNPDIyrlMdPg8mq/ugy7ZEIHy6vIVTNtLT
OXqbO/EvEt6NUSmj1nUJ0sKQ6K0tg1VrgiAFBLx+5nO1DlVVoMnr5cRgiYMLybag
KPALuK7thUpZcCiRhcH8K/Hin1eAN7+6fuaOi/KBl7W4kf/LaIF2+VmZk5eh5JLS
i7Vwo3eaM9WbNolSjlU4zPtuJrF3V0yf6/f862x/gXACoNL3+9cePvjD3MgO5HnS
G7fJjvIPODZ2teOzagB+0Na2UTZupsdiMijqBz1ZOoBKXluCHcj8ElHdIHAOK4iX
QyQjNzrrB2zZ4qP0oOwaMEVMgwtJPIifmAzLfBiPwKsLn4iYo7oy+xrt/OGC9vN4
zBN78ZX3I6DqEd8AJuTIaeGhuviXFU1/csvWYdxYd5bctz9+3k5hZbpUcblb5LEO
rdN8AKjEszjEZsOZfk2Rxz2PHVJR9+osw3lnYiNtXXPXRtbdYYO6vOk8c9Jarof3
zfUxZ+HQxLDHRGcaD4ykeOvmzxnIXddO4hfQtFx90xZPYcJUxY9VKhMuy06YQWWk
J3/v4BehkmuBxADfq7PIB/QxX2ujQ3XegRT9vP9PJgwLzI6G2nmiXblmnrDrtVO2
pp86asfwtQvYZu91be3dNfSgKxv+uoMSiVLrvdGdXettInu48xAyFjU1MRc8HtPC
a98HLNzgh4uT3Us40sV9g1ryx96XxB6M65FiyQKHy5FGTCtJUa0TSrl84iGTbgPv
xtTl36Y3PrLR9oJF4X6AY05ZevbUgbNz1URRB3YpY1aVxIX8t5Sfuf9i0q7X5GLA
QN03hXl22MMT5GvmBOinJOjcLkUm3NTm7DGe+Yx58fpQ9BlRFEUu44q5/bY1LMZS
z0j8WUFkf4jwTxB5mza7pHR5leYNvjYo5+P3YcXOwEEHJU8ys1RaJJoW0QUgrN1V
1UsGdj2LBzl90jihuTfbKf3OUFvym4sQKzSeaFl6VDN4F0uS15Xhvmx83cG4JdOG
+vacdze54h7bfL8CSm/6ggqgRl3Lm976kW0u6lDxLJzG0C1LTm858kR2DEWRmRcT
KXjvHArRqkujXxh99B8wB6qYE8NqFvIdcCuM3tPdAnyh+rgvOLcFv1XsZv08Azbk
wFW/E6a5b+n/MQ7oIt9sAPSN6bqiK2KnF8HyUNOMFPCKjKklZ0rLd66EJi3LoprQ
iCNpJqdTof3RfI7Og7TOniG/RIcHtsAlSyZQnEb50sXeFkZOuvnKyMI73vYEoqwV
PL+bV4/qyNpG7YCEZrPMJ81KpSad9iYU9TliYBsbwQbq/Nxj9feUUXS8UqKwprVX
+OtMT9TXNNNqe9WOM+mRFBz1FKH5ZVjRZpg4ar+qWBKTJklexmqmOpnwUkDNPu23
2sBXE0FluQ5eW8uQwfIxp/a9FkWEfcy22LDii+fybIagboyzGK0YJRodoFwzZG+/
XBI/0Fm6UrGmissAvKswI57V0AINBA6NJBFWvTZ0FRDS+mk5WOxukuzvb7l68rhH
RmRrnagDooF2dhsuHqCArVAcuSa6Q3VO2l95rix/E1c7PaK0Wojixd3QKcCKWjC7
VmaZLQesqUeiXHtVkdNPFddJyCicpCuKP/wbHbHk1ZjTffy+omux9/NaGZORwarX
BYabCzDRZgCG39HKK5XmAoVrJDtxPmgjglWK8cmmD73Yl2XkezC5Y24NS8jBt+bH
8Rlfiae5mLpCqFByATQfbLEa/0X3sxg8dWhsu/Jl6NNvq15T0otfS89Yjr86V0J4
p+z/FKExogT/AcH3P2eBKWJ7S8LFExnMKlAvp0uqTujBsSBT4+mRAk2vf3Ecc3J1
PRWFj0mrlz7qQL/bTh2H+Kh3N79JZ+z9sR6k7kkKG4OpnoKx0H4puBBx3t0DurPZ
VMtXAKSD26Fctv77DIzf/paqNRY2N+5eCSX57cKzYvUzmYrH/gRQYZ2hbMSqYwqB
aJC3bsiS3eaAj1ffG0xmhyFwU2MPT3m8GwXMOy7cMPQRUq57IWl/dkAx6h/CQM0B
GRGfDovwE885qq2PmTQOlwBCDWseWc2g2SYO6a83xYG3jrF/K1at8duyLf2WMmWV
FIdjhldPcfbtG7zDOaDer/9CnNXdDIPtwCkjfY4XtrGW8vkOEIdZFcbRF1qV0u4H
t6B9r4YLqE/upz6BQu2Ejpqw/Ame/MIp522uwYKC9qPrd1T+QkFPaWcVjgdVuoXi
IqVbMQxdEyLi7ucfD5QiJqlpeHPm6D0gu7PiVHI+d5/F9LMlHIBOMIU/stIy2mVm
9e9lgQc3zSdb5DRbV/5iT0+6HxaEEuMdRToYR6BJCWR3rAG/xqGTnmTKuG2iZLi2
lqM3KA4kwRgr3yNzTrAngf0gJ66NBEBnhkoEYxob9LxPzXU2PUIwm1eXrBf1qpHc
K1OXKOJ5yG5Ry9gWgkGi/rpmkAHIIME8fRksnVa1t46+SA1d6rh87YRL4JWH+hcM
MpYlj6TGglO8lDZ8f5ciETEn92Y6AnLSHvWQqu5CUbOeb4SXa9kIK0OeBluwT5Hw
qAgMh16WJ6kZHSB2e97z/G7/Tgwbb2WFf6Zfl+Z/8oi3YBQWKkWMitwY5y3bK/o9
2/ISBKRjKUmAMH8hq9GiO0kx1GSzm+/G48+GV5h1GgynwEohoHoCzdrmK8dAVXWZ
XX3xvkQCypxKir5blH8dpE2uefWgpTy1ocg4X0TVlveuw8SnNu8WEcvwWK6O1JRB
gnkWv3vBpDWDLMA0KXMSZu0S9vrqt5mW6+jlizZ8xt/rSUHl2etI5oDPGZwWNcAv
ck8vqcSKlEFhJSkRyy0qFx8Ze/ViMPGFnoM6jvaUyq3+Xxo04x871Kpf9MQVyMfS
Luf+o4M2x/bq25iHNjJIhZOEHDcwyFyiB3SUPo8GY6OPpGmgOZZlur9hVQQblQ5L
Q3OrKm9MRi+uWQhPsO4P2P0TGqKch7Xz1RL2mrRVkXvjoFa1Fs8Tzk9uqPn4PPGd
kqBbta5xCBiQUk9lin49ipHHvnoDkWukdiYBkOtTQRObfzfKE898/zrUdYOTVdRs
UcGZCdYVzuwMczi8VILfcHjXzPpgIKSDgQExAvtXQiKsg4/TWjcN9af90c4IiGe4
T2+3XdP1fOv0qM/re87U10yqukAmgV+ofosjF6F1xf3/npJf0ulRDX9w5Sz/ogul
cTahJjQjDxsZFczItaKJuKazXp6eQWTHiHN9y+/b5Gyhrp4BIHCq6I6c6NWqmagQ
xS+BH7mdWrsEtylZBiH9CVinwsuGLmOA6TkQVeD6EypDAgMr59W6XGNVUzfZ4F29
g+ZEiwdCM/kKXCEc/lHAPciR3p7N7MEEpArD/KUsY6OYkLKgBVcJQ9NQKTAefO4p
v4AhEUiYV38E4JVjFp1NoaEG4+A07uhp32R3o+E5s7OKzvRPw1mxJQNJjfkV3Fo5
rzQymeqN4nFi+WFwlbNDvhpE1pz6SAZSMtRrorqcNCa/syyWTF5F1WPcJj1xOICm
nfyWZibPQkJF4OYyv4HtqVaIL8Ap9/WIrciOS8p6TlR1l16PD5DviJJGii4BFkRG
yAPrBNxKYPC8pX/Hln7ahXAk0rfqVPJtNYorJ0qxSS5vCAmtArIrQxG4T/SG66s7
ZceF3Freptg6NWRIYo6yar8NL9lOiPh/ipI1jQmG7HnJcG431prB4a8hpGhSyRon
2ZzFHQwPJBllx5sy7MncxOM/Dl3E7eCvmsW4FLC3RjKCJl7UeS5pzVJfnIUEQ/Iq
NPsFIT7Ejyi/Fjc/+ofBtCqvvGi+Io47Oaq2sW4z0+TtQXPJYUl3JznCoACY1X9u
4FlT7me7gn6alhkR/EUUeb/YlLnuTc8BVGoqOBnoZI1kg8XGA0IfrHcy/3eqcVPr
A4jhBlLT5C4w4eYks5Zz4rfXHCn1toy1+0Oyrjqxk92xI7DPMbtJ4HBUYBfIQlt9
mCAFW5g8vcKgpL1JYTV4UJ/g56hNRr+UiJzsxMtSsVz7s4aw6pNRbplcqpdFvl2U
0Oez8EClXjxCfduDbCTTcDGiZWxPLWj1s/zeXTRF7XjwMA4xA++8tgvsXrybW8AQ
V9eDZoLlVUT4oIS3LD8sPJKMU8+TH01zQKr6b4fIVwyhem8KRtjQSlXUbGF9hp52
rINJjQMTsQ/7pO3WcQK5uhhJgZ3cLWpZvV+0eEtVJHTQKcRelt8sLwmX03gSem2u
DPeRBPD0twZNy3y500x5+gOc/0IMQnmtpfGD+949zKT61y4HaBc1wGaFelUPLGku
aARA5E6Ow1qrl9G+mOmbEG3xw+sfOT2+EHEhlK2lGQpWaM0Di8/2hw7M0wX2e6t7
3rAvDXS+SeZyh6ie2SkV0hSvXdAyBsQIoeX4sQCEw+SytrWmvy0gcoj0S9nGQ4k3
v26xFpVlxy64LsyoIi4sO9ciRYoOfQTGQKoXxukW6M+wn3ejizvErDxr5nSzqkhl
T+45nM1Es4w2wqw/CmQjKzFUWrHdwcvlXKjZkY8PSqZYBnMAeztIPCZdoyl6ZIyn
au3n2vysc4FVSs17tGKaDYiMYeo8835l3g+Ql8LM7iTQIiJPcd/rBH6KpYNZASC9
z7VvFRwCartKXMEIVvHDwlm9dwOnq/rEeAaBBB2w7Ntz4Zp5BzH8AKs2mqh04kDl
nWwd+u1/gfY1ld2RWNfNVJFrRg4vl6Db2Z9kmACbXxF5xHcg8CEd/tRAB4B7A3O5
PdaL8Ss7dJbMAGQKcdGww6Z9zfXW1Hd2S5KLQeI3S0dQmg6K9E5xunXjTX4vCb2R
4KqFkI2LycvlK8yY0kwKZL95XD/Z78wd/NOdTZzKbO4U9bQeFWUIl5mVKAW0nUxh
HiYGNRv+PE4bsVjxTev2HQvDXM4x6gtfiql72XuG5ytSzf4B++sSOkvt9h4bP3Dg
af19o0J9U4+Vv8LYNiRp//ay/PAPSwC/H5hBauguR8cundY6aPhWXl8fLWGjAtkw
Jck3xopZf105oPzfDjoHwN1IoRp0DXrq0k5f4U2NY2rdgXHaA6giDjtSdE7niSva
uTAbTu0kVjKk8DtJVAr1fv1xD5bD9aIIt2lNTEg/Zb3h6GzNHl7WzAZpK/TKkYAz
b1ZDYS1IvZjVuWAc6FomCAPYl2uXj/rLVZFWGMwUmAQ7udkksQ/q1pqEWyYLwyKl
bvyWsp9Pige9+NYd6+bol3+VODj+MaYwBsSTggWFPRjz/R+G07mbaoekKxhokdck
9OkboYpEsceICGOCKA90RgX/ntOF8GEe3QjIokog7QkAmM+PTDkgG1WH3hKgfvSu
MObNo7G0gxgd1kSn2HBVIz/oYfLA6Pp16eaIWkc3vy0cFwl3S4tOngUgaBTeG/7V
JRYQLZAgvSzs+XgcUOPIF0Uw+n/qDjMJgtTWNioqmP3EVmwJp7DXsrP/ne1b9838
UyWMPdrws+/SNuKk/jUcEhqdDxctGW2sOBtiTByumV03mh/GgPa27RAN8B9zkPNO
iTh+mUXwWn/VxlNvg/UkM8xG2I2QrTZ9TIklXJNTYxkM4/luzk4B2HXFCmuIo1Op
duOxUVtBjQZ2XmH0PAymE8joEfdKXn4XZwHfcBMMocDUAuRzWbPDIR1EzWl1E46R
h0FcCNlFLPPSEaX7fJyEDlf083KKf7xn6Nz6CyOKrPLERTZMRpG89S0tyCrkZymM
bVAzrbjRjd6AtJG6touWfSAm7PC6CoVd7P6d2pMFhxq16NLfgFdZYbr/4+nletsy
1sHhOAqCtB1otzhR3zNV2wcOXdr8Zn3I82lMGXqlNCOfHjXVaEJGVqu1Cq5KU0C7
xXZOXL4I5p9i7GJneeVLkGkDJ8n1En2kymJ0wJVV2wESqWPkgD9gSh/BVMWdr5lH
veHzLowIsJ4oU667zvLAqDfXtsMCw4CUxfVZm31rxhoVVPFXd7DZKH8cTqIU2Z2K
Ftrxo8e0DbFXMi4U8cAvev/i4zJYWDBTvKOpacqQPbcz6tulOJkgvSiv0ubldbL+
xoAzm7jskORawu+OmGwcCHuyHZuB9pqnG+0JVb7Z3EZsXnU5grfDzrISbvrBKzDf
sAXbO2FBCEZgxm7vocC6rEsIb5v2uelx/vEIKQJz85l0UvuPBxSDcc+0gTTtZDw9
ljPNcGjf+xd6Ws+3cxpjV1ZqslrVv0S8806pkVKPGOZNzdVVCDtktR3Mn4asda5L
/np1QX+cntnAgvtx15fBCSs/w6SdV4vUsASX10qh8f7c+y1M5bmfDQnFikPY4l4o
gNYTIqEmjKBa0xBb9yx9Fjp/2JvFT8gB/Sn5NdS0gn2tAHPdckRHoFvGbPq+dsiR
Qth6xdQOT7ZfN/2OX7Zb+tW4D3zu8rpDLQ/X0KIRAJlgiAFu3G8+LJ59udv01ZuJ
Vd5PPuw4+9Vfsxamlh2u/C2g64FQxU5zOOqL+6gpECeyRCuH39aonOg0TsS2AWPh
+TJkGgClcruTxWI4/cPCV95U589v2bYiVH5wkSev24ZoZKvOM7K5ckYl1KlJOHrm
6YRt2aMAe3FFXwJW5DUNmMPs+lkw0mSKTNrZGGLloFTn+u6HkAWgLnEl16nahIUo
Uu9sjgZCAxjrbOv14vCp5cmRmtDHuJ0dg9U7W/XrXUk0Tw3pzyd02Fcpv69Qcu2C
M69RLU+/mR7LATi3ZgTR9OZo1oqhVml0KtrT0nR6RxuRHnkE0f7VEZpubQ+8ARjh
qzSO6Z5dF0zxm68I2ppgaAByDSXB7k8OKl4hktgHY/dVjd+fZ23jEwCbg78xbzSw
ogq/LAzPJxw/F9RyR4Nf+ipjz1DbNjYrqLdsQdgv9TRRsCKCL7/2LQFq40zG/2JJ
JfqRvwzIeYnfQ0hMGqi3sPt7ofh3v8KZ9urPHBRe2elAwRZi4WVbo9Xr0V7qGvS1
ebhwcR8QEdZpD84YtpwICoaN8Wnq4yPNuiN07d5XU9Vz6hXljlYyJzexZNgxfQvk
43zib/9RYD392woQnIjv2EL3ZDygVc1uwQUq6U4PxJpCOoL1TjIvUrOhFyDFbZF6
9znlVUktSTHnJJf/r9ND+s9fkWh5SXUKHCDY0VzbwjYd71KCBTcUSFyvSTd87SDj
lbDfUlpJ5WW7hskhETHM1V1fID69CE/DHfv0f+PEpHFDQg23vUy1WQDBl0Z48yrp
Tztf0vZF0L3C46q7OKIkReFCCAiklibq7Lms58Vlgkso4L9v8Vbyya9zxL/w+R9c
o56QTh8yQxgNlsDsU/H6P4u4Wc9h8cxYjhgGQKS2fg4e6ltJakaA70QezvVP/Sb0
SUs5Sewui1F4OCEwto+RWBBUxcXMtU1OMptMFDzVWd1jW3R+/9bpVDgwYRrZD6JC
heujjPdkAaWFYU9XcGVktanEsLgQmpa8Arq2vzv2lxEA7U3ltyjOeVyWHIlP2RlL
yq9c4mNrZcmb28ITM/Bwy33nDqiwH1NTow8S58pwOq7EqQqqSm5m+gqxqRiq7MiO
hcWnM5ehA94P3emIfrX6dWK75ot1Fe+oZgfc8SLXErSPuRjW/vE3QZ4GIh0ozTPG
JKabTP+xwgunfSpOx/k2wwX/tXg21sJ1n199vPdtkWYoJib+qSud7FviazvXrYWe
6AHH+FZb7bp+4sH4kT2/eTKJmWqCLAKTSO4C7XWLjx0Fm+kPgm0ijBmip5+TH/nc
b8LxzJD041vQ9XnGc6l7KxToVS3MVR/3nEJjzualDKfLygXobi2coqLWl52aq6QL
PAxDxSUr4vs73T/rV9EzUjLsgopIwMnQpnokCAmxPJkPlbNcatvAVImRUfWzF13w
nbufau9U/IUD+COXv5AJuyep572jyq4cQP1YIY52T77NiRCxT1v3tKVbMNNURu99
GirOIP55JraCoL3lL3rEdlHoQJDz/BZgl5Gc+mFbEqyRZCUSR7071bx/NnwUjes7
DvwzhB+SdZ+nFPbnzmYPEa/vWaEym26mnyCAhzrnbt694O3l47ELOsof45pH0aUS
3RMx9ve3mmTDPVPKb1PZfz9dds84OEbu/Cd1wYlo3jR9afcrFpnQGPR99xU3DEht
Lfatm5BGZIhfXYWAbxgNH7nuMdO+BWzHZnug3q2ApS6TSkYBYutvMSYzVZIjxOaA
6hgX8+Iz3i5XyVjv2LnDL2YE5FXTovA3a3cd4hrUkaHND/DPgjCtSa6+5zvhItqb
efTrGgHQJfjcbra5smWpO2/YjZLtC3s5V3EkGC7/36cP+zE1R19IhQcHdLQxkwfT
EBlVgyd0+xHOfe+Hw8S1kgH/3/EW9a+PJDFLgFDxMP2PvVY2Cn4BGo7AGseZZf3z
4O3fIbnCj/hDXAzLEGAtP6VDFrvgLvF08BJRESBGpfJ4IPnDBT3egQCdeOyq3A4a
1e2SPidXN75alGsLij/etmE7anLwXLEkbQzajKZz+FuIwSTi4Z+uTNsydZx6MFDH
BF2gdpVpU0Adg2xUWROrV7e99dA7GaxiD2JaUaA/PXDinAecufiikjXiN7yvzGcd
t70+Sneiw2ubSnZBqO12OR7vDBePb+Dx1+EbzZwV1ddgiN2VTM+INDF8WibDdUio
PmLRjhWPbJXNr+W84yOaKopINVzGFCvMS3uauvpQ7Zugd6ZrBUwZMlHQsAAAjpra
8rA+N7PGsrPJPyf05CfmJx+oiu1kVVUAEv1EfkaQqc4+ngsvRA/NDF8Lf4kaMqbj
X7KCTmSB9IaG5PPCLNim3lLsUu3AhFwZLhZtcN5CQDI9oKB4aYGBbFDw0prBvMtq
13onk9USgI2AoqqoQhQqvXYSCEhmUO6QMwbz6DwCPCXlMarP5oqioaUV9hPwXuHx
3pejWmvQ0mlB/knaRMRPx+zi4wRTWFjsg1vP8cfF1fp87zYoPyeduLj5B5zMlvhA
Y1EBtvkxDrKhJzNvFcYEo4jQ8SxGdy3C9EzpQ3A6V2zrItpwtQ3ORHNy2Voi7JD0
7Os+QF9XMNEZy+1GCARHJnI5SWQJTIF+fAEJ+p9871PLVXImfBde3l1B9DESuQQR
7Y0Ja/BUR1RH8mdLLvTR6bfmVLZJbdEaR9XL/CBilghUkqdvy2DT3l4YIkHaCzl7
g3ggSjEcVyVTQfnhB1GfD4AHjMSGBUPxu/GUUU/DSQcu6PFoRDKkeVWq7l97E3dw
3BsyAcADUhrOFjG4aPdQzWXS4QcEmVukgKEzgXnQTIp+Mk6HU1RZbjHgaOwfZAJR
gPbFwGnkm+MohkO6XhUKXnSXmh723faXykhdtDVG5PmqLQVFqQi+N0zrC7VTwGcf
osJ4vO1L5MwgppmEvLqm5Eo8bHvkM9zb8I1wQvwoyE3WzdEVS58jFyfrR/NoCMPT
cW40Ka3eBIS6Sl2OLhtX7/RlZbDYBpdQVvv5XRpDoEWF6dlrzDzTQqAJNFzzgaLY
C/UiIyQHViswmLjuONIy2xQNxghtj/MKZVe2FhtDeMMcbKPwQE00Oia8zT446Tam
kArutWkKvmSefVRw1FJYD3TjkkwpQVIZN+ZPDGAt8LEKFFdWWwxQ3YSRGjB2pooE
7tgj8Bja8+CO4P8Bketk0NNvduwhL2OPKl8U2OR3uMNmDECj3Pc434O6mduhxXVm
zIL0tf3qC1ZNEcc0ZDUqpSpC8XIcneweYaTAJROeLbEXPUpU7RFN7Ptkn/1+qJyR
Y+db6vK1ASqRadwWalxUvo1VxF798cYAdEiGRMNM+ztH+vUWHgnhtH3HnQvNLYWZ
E8tSeKh2zi7/UgR5WMi3Nyjl9thYEJ1HnXgKgBJMPIl40K42+rpHOl8RY5VbMTrU
IodZd3SYX+uybJNSYqtBMuP+edu7YLnl8DOFJTFnLjecgkkLQ9D8zU1z/sgvRFjq
dnRe3GWmaKvcqrrqlxQgwabXOUU1F6LtYCQCF38kttL7xHX4GDQn0epgaie7DWzk
d3vl1u+DpIAL60dujZml+hRc5RjENRP5ugp3uePC89air0mtvIhFH8fg/frn/5gj
+c/BiY9ZWIYEEKxuGukB6kR47gsL8jgwix5hPR8nU7bn9qHx30XyhgQS314Yeery
ALP/iXDcdlLVu7v3XIw1YmQYg8Izzx16ZXy+srk/et36H4ZMrGwzTJdYLPD64Tx5
T/G6LJv8XDNLYDQgZdJMxwch2ASPrdOg8L5Srqy4ZafLRntXfyb70g+HJnl54Iuo
FmO/n7vCDbi/eTMzWbcRoeAw869YEkAue1qz9yrnD8QTL8z8opwyfV65OoTaEsLV
h+mjmvgE0eor/PcnAZzphC8FQ27w6jfqvu4ANiFCBBXQlMpaHGa7oQpcKrgcvYWg
sBV4wSjuCuX7owpookxgA9cnqxpKlpspgqQXhGagdV5SLREnyrTBU53rp7NW0zNf
k6/aV9Nl8pMlS8DJG4P6nCjaQmxUpS6Wo8jtP0VVUgJkOQ9eIbmkMG+E6mqpl08F
dOSumg1MV8od6oOdHX9pTMvqqd7Ab5NB9gHKQ5JhVeeHqxc6UrVsnj0FrHwSX1M0
d6EEYWCUXtzJVnBRxG/Mw5naI9RYTEiX+kFzSoxwvVOD/hhCX2trz6xP1B8imTXU
Mzt2DXNDELJhve7jzXXhnLhH+mLeE8jsJq9pPTRKKxDKLAY5zEJjgm9WJzWPK2yw
9meJLznt+UOYnPLFAhjZPptZdblIYIiZsbfKAWaquwb98768EImdVRMDZf7oYS8W
tG7Sh+JH1l+T8Wio060xKDv/wECE9KaLIqtE3jadDqexZVWeNno6F8SoZJiz5c1H
keBuOsDRTjkWJgdiC3+jKRAlTS8xYdLMFzVkFXpSkX5IdZEvsUe0hD9osQOEXKlD
zcbao11pv0g0TQinLOfKDzFlJvxqiWjmfCiYb/+B49jr9F+d0C4YmvE7N2GGooL+
x1QxpUFKh1wQWFyYGqU0KgBpI1LLDtLc7U2Ho+tMFjSCWNvcCi2z0BTSnK4a4pSv
NMaIgupOhfQDqBtiZ0CYqTvtpfWHGBsFarLEDn2Vt8/Lg1Z9A8pVzuyDif7NPDfL
xNuzPTd762sKU5oBVIuWWBGbVI5wPS8dTrXEQS7+15Ya+s3Yizt4IIBLsKF6D64e
Vqio9wNLe2IgxUWf9BkyxTHKEuVWXbo9qTRLcfNO4oGC5bQicqNeBCp44F4qeaC0
HY6po32+fw7++sIE2veEZVHwhH27mwzxMLRI+pqasNF6vBKSXCrJTnsUuDI7m+mv
18eG5ALAk+dG52iRJSiDNF52XHrnGjYX6G7FmGUKBRzgD6HIvU0Q6Hf7/wMPKZhx
p9Vrk1fNotKu3SS45XyUwTKA1KHrpq3XQP+z3JLZCMPwYv7n71zIBOHYM4d10V41
ZpPWQJYbw8d3vMHgpWqDy3EzriiUuls9J+fPJNYjobhunG87Lph8/re63oiWsfiA
ZopYJ5a0UWE++bs8onl6BJfcuTc+DgXBBl7n/ZyLYWyWYz4PrTDoXSfTCsnKyXrq
ARQ7ZAVDRAlB4Dkm/2CNxHDlNqkY8t3zzrpyqWBW0oBE9Hkj1Mv3yTzYqZp5FAXS
YaYlo5t8SnUJtvZF30mQ8QsXg7tk/3HV/9GH2K0qmOWBWb2js5BuzDsEMqeQRmH2
Vol0epmc6586IyfgX+Ssqgk2cOyyqr8YSbqnEnJV64zembC78F0gT1o9RZ+nPv9B
EJPufJ2PExY4uSb2jUh5RbfqcZAxoJIicxh4MdtK3OCkgxoXt9hq8EgWVQVGo+LN
AN1opNxzwRhbezC6M2ZTCcFlK2/PfqVG+JBrJ2k3GigAeoSYSQzyPB1qm1tdQUwq
AT8clxdDdbKdav1xEvkprtQ+E6+ve/mnIiuUUkaMgk2p32b9rRI6edenfwuI1E/L
51Iv2BUNLMfisyBvSiR919E5x/67f6J5UBhalQpAJDaNHFW9hylnpXTi3GADOqlm
9vyE+wNg2NMcvqw9dPBm+POaWvEUkhUddw1+2D6eZv6J2qQSySmmDIv31SnomuHx
QRPtnHNiNyKmaftdDpo5rUIWv2gALbK1z1W47/y4eBTRkOs8SMwZ4983vfMTasZA
CDvyxi6FqgpkzqnUv1VTtcVo/VeeXiMml1OsH4pVNuHyPhYqXNcSFaxGW9rQgzQM
6mZ4J/xvvuBHMmMUMqarxccfGN8gu3ouOYdKzjhFBXK9WDPhs6u7b9A4jHtl46/T
RtkQ3Y3Lu2McTG+IN0czyhyhN1ytV0fGrTya9nd4DqmO6RCBAUeYjrkmsgGzhLPs
XFnQRHOKARFMnVxhXyqqc2uPxLHN9gsrvI3tqQWbJziGWAeHbwzyiNJCsWTR61D2
92hrCO4v4J8bpaPMGshQJpiEXTDx8xLNDBsnGnjr+zM0S4HuRKIoeTGz+12ADn7z
vM2hGRRfKBEzd0ZsC+EI8miLRASuGMQax02scvxRVOC+oBTXgLEJQJQ++l8acmjB
RCK1NRRNOThzUy94woMYCWD9srKb0Jk1h1jMNXF0iXhZX/KessoIV70FG3T1fc+j
a0fuVAvbi3ODC73OWleTSMsZbygk+UR1VC6qfwzVAbA7tD/8wKTJece5Ky3NpDdA
Zxf7Pm7Pp8eHPQ79dEcNP0sEk3DVZJagjajLLNTnwXjFIRej8hqaS3pxgi/irpGq
Mj9u3j99Jka25hIHiQWKZr+wQGaGdBMfwPyJ5p55OPu4kE8Oe2O1I1n5gv3cdEuI
cJ7YdxrcIUFma4fKJ4sUWodi1TB3LJTUYKdNvTCEQIj8UTjOqW1Dv1epn0Q5E3PX
NNGV50VzbAkH+KoOxmdMOezZTV8RYhEd0ZAp12LFlYc92BGcsUqGyubJtE87a+5Y
LbOOCJGmVC5ZNGo8NPFVmBv1hUg8Q88vXDOrLD2z71CuHchBsKJtuIagUXtjZQYm
OelDiUsCyiMRdnpulUtqHLmgAUhi1OPpGav/RK2XAVJ5+vSdhIzUBRwwP2bPwY2B
zyoyTw263H6WgPxjs2r1oN2ZXQdKNsdAf8pZIySvmiPKQH4BHv83XgAAXnMCh9tV
7kXncP+8uoWPcr41uXbRiXajPogHfDnXqnXYPSJAJuF9CvO1dnGfcsYMWt9jifDn
5cbij6HusrJOqfqlbmmkSAli/n7Cg+1ejgi6QDFaUnJUllNwhz+Oi/4WnPOPqHwA
pjiTRNV8Zp2wfbNsKtsMLQoJTJxqpoQE72iEQ2nX6n2OjpTp7xEUmJx4d0rb75Iv
ofnaot8FE0kwqd9XfEifjKQG7fKx/riByBnhtAyzk0pOoRvHKhI8BUy1IFUylL9J
xh+bU1SM0dQ1iFsGiFRRjJ2Qd1LTm6BPHSb41hl5FGUUAF2497UocX66/6Wby8Ph
jQYwGXXwqiOxKP2P3GH5FY6jHXOT99h5+gHZCoUpgsFCTBHn255e2rtnXf/mxRfz
WZkAS/5rbWL/TrR+gRqzCj5uzJoyFW5fK4qrl9ltqlJnxNsSCjeN50Pxm4x641Vx
/6VW1xEwuGgFMarURBLEblHpI/lKzPB15qTLhdSBE214OfEmsWcaEEEVXq5syut2
1LPOPwOn1IZ9blZ4KkHkseFIkuB0GjgsjA5PdRTyJ/fxJtLA4Nc618YJsFEAbFo3
PHH7SgjfqN/noGMWHp+Q2jgVvM9iJzknjZ3KIx83W84BaH37ULasdlO22RHBcG16
eHjACy3tWwJ9orgfmrxzwXuKs+cMaQZ1oYdN//vqHZEutwr/COY14QMQJC9jEvbf
geAqhkM8Z23DNK0T0hlVJMB6FbcBvarBKc/ZUV+A8Ojlwk2tBbx6sZMgiwYi/fun
vUV24wKQ3g8cRpFDPJk3zBWYC5/6mZiI7+Jbu1+RtwuBvYke3h86LajN+vscJuFD
F9ONUrUYJhMFHPbvDEnQoIdichKHbTT2VixqeppVi5nQ/DjRhiN/pLMFyWWnQINE
AET188b4f7jPE70yZvFjnkpEkEiBe6PbtzrL0w5yRnM+S3/cJ1YIiZopmFZ6kdi0
Ya/E0fegCm2l5bsZFdDXmkJcWeKt8vJWXlDX+ac1Th71iQDX6Seg8fMxne/H42Rz
1zy+2ToT2zWDvLyUxWKWfBQW3+DMStOwB5c3tdY94m67NtPcPQ9L76f5yZhrNKsx
OtFEvRGwehIXq6jX4a+hAhlp70B8jAwgnt4I/V/Cc4TAAf26v7GR6uUcZC/5Aux7
0e/f8f6IdKELv9GqNgWqmApXC3ne6dQS5aTgsFm53F96npmRSxeLsIhw7sjkuj+r
Fdo5MZR9GvjjeU7Dkn+yS2lzTqWYyZj0gcvnqp72KYIlfM/M0x2JlqTqsJoS99YD
DLGXpYYmdpnXthpU+tmn7jnjZ9DqP17Msl3pO+9HJJ2x34396uAXrCmD1IJ2RB1I
Fa7nytfqUnSpXdUC0TfPZ7ZnDnSXxduH6yO+mQplURdrjxWKb9ISeDEw75dOlUbw
LJadXWxy/iX05P+0OR73dJ38ITZZ1FvnwPA9urIxL6UO90KDcU5pSCcFQ+YS3BVt
cvGj1Sa3De1JwACZCIClDHYgNXy/TU1W0UyZ5xF1FIUeVlxTxmvf0yd64hlN3Uew
t+wjKuGKiSmZdfmEreqRI8VyCM+BzMBSyC/DI6dwwCgySpxWFCVuxff1X7HqopR2
EPW+/XCwSFod020QcjtOxDiFsiyig+Ckpl5oEFkKz/QxF44IODw5EXpD/Q33WDbi
/zr7TNMRhRRRu1bXkP6DPEWx/Kl+KOtE2Ji4xqcdpwgkmHT+nTOBElCEil2VZbBG
ycIrDp1hx2xlWyAiYkerPNUm6UcM9SrYsFvnSCOPoQtEp6lXsWcCOS1MlLT+KOVS
8k5S19gmMse+5J8Oldnif4IpvJpcvF5cJLCU4DUvl5F0JGCaucISXNnGusnbou2y
NA8f/FcB2yiSDZ5YajuqGTS3l1GPgTWjyeKoAn/mPGrKyRBfNBy0PvTrmAGiioZr
OWGRkyOTNUONjPLaCjH1MMtFjkWJYQPWXMtBr+tcdmEKT7I1KLgj/9ct1mNKDp6c
2K6/+Ln4Ksf29pGxq85v9RkGeQb5+wNZqFaiAYVS6tIrmVn/uM/mZY/5mzGFNNW9
AZV+fWUm5kHayvNFDsaMlPnVgEeY33dtZcKoeW6Higz4xU6KZa2aOYF1l3axLtAB
U1VaW3SPoq+yNBphWeV+XUIixZfdDkVttG902dGJa/sap4mWsOxuVkJcdq3xsik0
bV6S2iPy366Yh8ehuPhyD/NNm0WAzv00GHN0R5kYhwnhwztc6xCdoDg3sPdKpEjo
p4wn3TaL0iNXKNVg3MLWtAC14DnR9gRmoE6L6ach5B+sYwpa/5fBaD2w1wW5FbX+
mROV6Pbg2OyEPO9C+VswwKtleHCBhUeJrW6ovbddhBtB87sFk9d+4fcDzIPRcB+a
xrKm+5agCrggLoSSCAUOUGVChuilQW4QyWE6dgxoqh33lKnkBybiO9Gms0YICYmQ
U03KFN7LU6Ba4oxB0qZ509ucFWJ0UarHptvMVYB9Q8UrG8WJjbmGqRxj3691sfTa
9MSf8umQfSFVnOVo/WdwRO9WZElnyJBHhoGWvXzy/3RKnJ87GO+UbBkV57WxrtBt
3OMT3X7PalLx8YfLh27jqrL7Gn9pE8F4DJi9pnoUb6AscavmxqUa0wRPMlG5gNxJ
A6+EOLRP89e6WNVCVfCYrbzBmYW/hVB3MVaoGdx8zBVYOx85Z1cbAWMj6gtulL+6
KcDQ3p/qz+2bERaO61p34pLw9zVnXeG1evotvhpl4mmOluRuVvgLYs1KjavfpjWh
d5IFxShC3KpcmiIeKxYzmvFhhDWGOA4ZLKAKjcYK2zl6eWoFBp0Xf/WWlRrnoAK2
xkP/nvz7CWkgK28p67Vv16l4c3KUAs6xUeUoQbliLX0n8WKKzljttYPOZwirKbVG
8YpcVtd0xPAshw+a+ZoO7AhyJFcsuSSIb/pBC5sh/vzMY2xw8dm80ku6AsKDUK0H
+Eqv72H5azonaOIPqft0lrtBiX8i5Kz+2R7JaHuTa3nmvV5qIKRj9bU5aimeVX/J
ka7OD/dyM2M1mkzuplwBGQ8SoObheWlhsK/P4MnTuYwKDVJgrTIRfft6WSFtsLJ8
Z8A69va7Sz0BxaUiOa/VCVXrC+eKv1b92/EX16z7y5YhKkWlQFtC/CNxKBw49JgD
MvNvuFMsMhAkKjuUSuy6vDmXA+0fwRxbc8qsmbA4f6Ate0TDZY+6TTmifsYgiyiT
C2TtDYk/J0ZMZOPy1AjuOosgEbUrnwdpsTuJnWSpUhW17r28twI9pSQ/3VSlIWYf
s5dXbiK7mMNuWjSjsQmiTXSJh2OwQUfHPvHaG6tjFndGnJTf143P/iG0qlsM1KJ8
wD7YpX8HO+VOtOrKs1N6eCO4GX/LuoR79LRPXhD7KmvoFKuQugYxliH5QM7FGAr5
VA6ABWM5SQaqYhKUkMfH2vdTPCOAR/eC7C43WfZRr2vcgzWm4XMsU3iDtuhw+NTb
+960YEvlplZ/KWDCPankEDaviBjziXoVaZAK+mu2nS4FEIXoUg6f2+5BbvH9gN1s
wlACWYwDRfWECXYY0K1hGtYvpyQsHsDnF+/K3mgqxrHvWOpJVMu5CK8rNZq7c61M
0ak/mDPybIkt7oNbTkpSMY+bXeJoIWOAaJOGL4qRbHx7w+tdKDWhyLx++hpiRYeq
yt+PDmlY0Q/SMd6DiB4Z5bgHUc78/jRRhqi2AdY7j4Qt/mgop739rgB97CWIKcV/
xH4KJOnWmmm6Y1Aouu9uFDBNNxGh5CbkJr06yFNQUYA4PuDA6X6XsKPn6H8j4xR4
nVKVNFEfyIeDoA/pqbzTmJNTo3bJ4joCCrtjSTMfPVirKkPhuediZeKNWOhU1zJf
eN4T+n8PYDsf0IjIGFeKl/pDJTMxp5jJEhKP9plZ1k8fe2QcRdb15GB6Zju48T6r
YZStRAphinMKtseKrhiQWw2sYjm9Bkcmhh5nhtkpYWmWyZNCYTEUfXK0piOfqGrH
dsAWrQaJbV3lLAqRqqxn2qwxRWvY5q6aZGbyDf1bdX3uCv0rY19cnS2AyTRBu8DM
rZvq4zsYcoXKyXCsQUFxGzTZckRqyryXN6fbwi6ZkGOrS+FO4mt2fxiO0hIJYbRh
SNVqlr1467xUu2Yvs6RwgO39oP9FeQinwYu7xYGy/61i87b5n9lE5ENOsLI6KLTV
fqmS503LUrTf601YGN5TykNh3MeaQmmp2uJEpUqt85TAH4TOpq+87HVQ66+IbYkx
S7p4w8YiUvm5ecPILBAbeaIBDSHOOGNwQlFgBfpdGx1FeYCnzc7dk7kEE1KA5mCm
AM0MqunfNq/f8tVak0Ay5p4+UmXchhr8PpJy19zl2f7fhywCDlWsmRXX1TLlP9eI
he5LLImFAR5d1/DO4hFmElDZEGEH6lIITQ78zTsOg0x5lTS3oTuW0fyBS4vYSsew
hc3T1w6EKVN1hMSSdeRzZw9kiXm6yfVO8yo0gDubSldUIkgh5klg9ZN37ptqqWxj
9fc3psCl05MqA/Xw+37iKCBXFh9Xp8Fzs0LBPxb0+qnYxusEp6z0Z6+r6f30p3QZ
6rxKNUMGTAWYgakzq/4oeyOw49VKC3DL3MMTJtV2BiOQmyLC4OIsE8qjGc5pBUK7
/iDgmUNEk9OCshYkKRUaeGrSDN07LXZLRYWEkeGOBbVPzJ8MSD7EklEWNxpGJ3RB
iHtpRAyrUojXcfIPG6/hCoLUVzJdCDjfRjS8hFTOFNuxVXID2y3ukPl7FPhxSDQw
BiWha7tMrMNaa2ACswezfaGzb71Mc2EGHKkp67m1aL8bLmI7aW0HF81+AK9dUTS8
5bxlfTOamW/eWENJbX80B8LNoNN96R0CeZNbhGTAWIgIs52xsdA9a7rrTHKWio8X
d8MEGUTGZeZhYianNcUfjGgngm3wN8dmBvWKQ4Xpt9hfoGrQozUjHFHtbsPjqHaQ
aadaRBno3+q7zEwss6GAEaCxoNr0t+znciEGmHBPbARHkK0lXbEMZh8KUGBCV0zQ
0TRxLDsjPnYfgru37wVbNswGAvvbPfltc+NG+1ZiTeo3pU8Ryf6Hdje+7C52yOKg
xHiinPu7DytLAKvnp+yh74CFeR+6kR7ZB90Jyz0Usj8QmCuNQYVMDCld9kCs7xhz
yn4XPutrepbPgJhGpxwe0TNSNITPQmiDV/7M8w1RPbQcbRIACUfCHISECL176QLn
rvrBQ2UBJXmutDwcbxFZAoA+8rx5LCEa6KxL09GFcBpGUcmsWWf7eH0MnsGI5eG/
u7nxn2kOruluhCMMcKQYi9i/bzUCvUNVN22uYuGY8RfPZ0hh4FLEu788Yt0RMH6A
2rzkqNp3p+2ej7WNy6bFNREyJ5qvepnNlylxEYGuxjNLxwgNYufU6W1LclA+Uq1/
1U2JUOSVul67+TjsU1rlJpD2tMYVxFvzuuSTplqkK1exYnD6lZSqYZ8XGEdcVTNH
8hi1tXuE2/5G+FNx6NzhrIog/O7HbiRS/hQDZxs4TbGE/SgVc8xniEsIugSDOlsW
mYD8AeU3WdUYqIFwNyL+Tw+3qFnPIostohB1E9rVvWTiRphHyNPoOhixZoLAUJHM
nNOUvlfFFtOTpw3K6j/3fiHAzRI/vVAJ5NMsrg4cbY/L2EOqaM+vJ4wGGXJCdCIS
IMtsf7UTbycHT3zf16VYLVTkcwiExWcrlFyJaevOte6kS8YZ7ALZCHCnw6LgivNZ
YSaD8gNozHRaIBUcE4IFtDQMF32HsSnS3TsuE0e2eJ6H6fwA4B+TghvCgZM48ZzQ
uUuRnqJVB+SdlktMyMZsdpLEWhHZKXHj4zJXqckkBRPuuOO7rGxs3CR4fXJb2JHB
fZOWppreyNFSr575dyDh4gsyxQi/pI41sz3w/LaM19sN0ewvsHtC6NqHqb2Cn8Qf
MO3iBsY7sUKxHMOH+Qxc9D7hB0tuPvE3ZNxt32XtxKa4H6PQ9REsVBnLAM12Dm6e
3cdUgxu/PjGWIbEP5woMJXeA/ugBHIk/uAbk2x5+rSpSGI7bZMGsQJ/MTpsfXQi5
V/azLDSmf9KFHTDNiVkirRvrtbDzQOt4BbWyeqnk1ihK7Lvde6ooog8yr8XcUd8j
2T6IAqkZy9Zt3eUnKdfBvsY1ft+0iZfNkBKyB1IaYix8N5SvvEM7+K6n/B9cR/5R
J2am+k1lmC+DklgN8JCfEHmJnDUdKD2Momv4MoJ6AqCgWeawYgowD4yf5k0OILfL
LtiI8H9op50DnUMx3gO9uZDwdAYjGpGkF9XAcb9J+PXMrPh5z8rR7BTuoCC56ekP
XJE5DsgxBkLs8PQUzMzmquADxTCKifkglY4TE3ej5XnoR44DhZgCHDHDzalrQFaw
TEZ4JSM5rDeyBULQ0PUd9H+ZMYxzjzA2w0PMAhRB28OOx+qI8lJWzX5MNdvtAwND
Vc1gMA0Bqbv+beq9YEvpL/naVAJVeTh5FF4x+AW/B0vbDGxsRsD/s2q9oq+S4X7v
MoZmGUOTK1VA4wbkgXy8RqqmSipm8nnNEFXHDbrSpyKVl6ZbGs5YZ3IyRkcyMDhF
POlfk0+cC120qunThK+k1m/VjPRSx76k1MnjsdoifxvYf6ycd7Vqmb8mFLrUCoa6
0iVN5SeB2OWCRWsNVYj/nCWfOi+coumXvmiDzZ2FGObyRSwslb954VoWOYX/aIu5
c878ZFkN5QNshN5l6oo9q61RT1AHi4PGDFDmlvjlxD9z3iiGpsFMDWiCTPBza8vL
AtUTSt3Yo1sjbDt0Fc5vTPWDeym08R94Nlp94WkC/lI4Gk7hfd/Je2lrwV/xRpeJ
bMHht6L62bW+n925bXqu1AekX6IqHYsWN8LE+ztbJDZTFtLuKreGAsY5S9UEQ795
RJQ1Q5c0s21FdLPcWJ6XrGKWaGZOoVpIeToUUQxMBnrgSsb4UiDDcgaUDKhXwl7y
sWdddmZn1mY9YWE92JzUzFtE4ovUmENXvKBy+yBGvV5kSuVC2g1D7eoaH3TIyOXL
OJ81X150QPcIAVBo5mzFHYnwLEijbuB3Ikp3bg4W7lO4WwcU/mrQBzZIDos61R/k
as4bv+VMSlIk97WVn096AMCl46257OARIDb4kQASbnQD4QpgmB3Qyzf9yxcEEt6x
dx5lU52FJfomX9Z+GyqxCGP190iC06X+uykWAtkfD16D1OKhtyqunIdOU90ZQEej
QJy8rw088ezxzoZd5E7WFXLjRoIzNuHp4OUUKzYmNQ3rB8N6DTBPn1BkIfc09ubB
C8ft0MC4FPbeM0lU57cHEKw4SGm3QEVQR+cCVh0ZSjJZbLI8xr0ChFRlK5rb1qhH
+7I8sxAmgEihFFaNrpiUNm/auIfbd3YulFhxzKqp9MyXDcotKsT5Cbb1bGffLutc
5i9F4gi4G53otpdN7Rmuf54qdGYZ8xKYWQvPXO8dMRHX+qRsUyqcrsX3iXBfexPK
avZW6cr5yLxJqBefNKKTArEQqCU/69xGTiKYY3OkOpsCBjllAYF9nNnSHVPhDNzP
IKv+zNk9lmqeW3bDvfDnkYqNAjpoiTsq2dxueuaxGi3A7wRrvU+cz+vLBREBxqEA
iUeI/rtB4su7EjruY4ALvXSVhgetU4alImeWB9/GJ3LOu33WPAwX1My2ch80A9yq
r7FaBmXY5GuaNbtf/XUXpEX9gizwqG7DuX9+prNUa+Wor20RArYZdmBUdg+vlJtH
6Tus4H3KsbQhQyU+4MLyq0PJ5MkCjzs6unk/ebl4Bz41pZFrBVh6ttwX/rwxQ4uO
bW+7DArbeX52IiBarLmxlCJEsoTogajwBWLCUu8mJ5O1KxXuweyT54uZApqkUDFL
pdKQQXTryQ4F+UuJluw64yYlQqYcyG4L3gHMEU6CSNyBWA19yQoUgHdIzZ8X2KCM
rZCTYiGrNJLnCAEUsNdxRSdLFiG70XniCseal1N/LJbX3Vp4GvdRUXRyD/d6i6zL
I5IlmfPQ3RJiB9apF32kiCzfGoi1F2vY4kREbLkETDvYd/RxxiK7bUKn/ptfEWQ3
sAFeXNpX1zGzKGRXUM1ZjeWJNeIo3EP4Ef+spJHnc6Q+Dw8wpntnm8IalOd6WFw/
eITf3CQuY4k1M7KP++17GpA3bMz9MSHkIAZG3YSK1EWiVlFH/ue2cQsKTUePloaJ
VUakCBusg1k8sMrZqakysRPjem6dk4zJCoLHaFD9Zmo99YAw/muDqZztJVQreGtn
DwtNQuxIqDn3FeQTBXYX90kw7gZbBm6ZTsjvauqn2oiMcDSsNhAoCBxWdd5DgquG
itZzUbhMr0hGEgaEBIhxg1Es4sdon48XVTT074ZcBfVag/czZWGGFfUeXoyHHLzt
oJ/yAnNHAF/P1d9Zc5yG15f9PSPhZ6k6k9/gs2T/Hz7XYXBI2ewJsPBG5kYuZt1o
Jw2pHEDMtldLLui+Gb8dVJOs1lIW1OgwwnL33QXVI6kf3gcMjdmH5C8vBApy8Qkf
mcg1DzvlqdUT+my35vUoLlHHsiosEhqIOJe2CvEG2D+IKcID3WBB3/Hw3uPQj2ry
0SpgesjOeffesAeygP3MC6oFjrzT7H/zQVActuPwtNIC0RaAWx1955DrSJvCyj5n
OjXYjMC5CWhbcFQdZeQDaBrxIMLhqqu2+t/ddwAjv6xnmU+mDiB4DHX57hkiosej
4rLd+rHsFju/ENaD+mzjJQzQ9Xc5DkR6CYYF3a6JQ4UmPWh+Up+YXCZPzSajwWYW
1D+Yx3cs8z8fwRLOb9QwXyxJs5ocoP7weBDK1xup9TchbU2coU7Szd+qIAA1cBxf
YOHjsob/e9WyecOlKjJaQ1v03wkbXa05UGCzNv9umHl6sZQKrJvfAe1QnPdAnFZE
n8eMlux+t1vjw64qVrpQCwmiG+6jdcRdrOlIljLGpaz8eRohL+nxW7zG6XhythiJ
N6I06ehiDjNvpauUf1/4CjrBfjXMJo866IxPINEdyINzeB1/bKo5CB6gLwt4735v
IkelkW9YsdXfa36R0j/tdo9sBSqO/56YKcMek8zK/U+16fcgIfeJhc2o75fDjpRM
aM4D/fgfeosQROmsQn5xEuBbhNcYaclIf8imAjcS9jaDjpTmRMiRH9QGVLMoX0+w
gvGO0CibIrxs9KhZ48NoNZEIMK3JeVCSv+xLDx1zPavrhcfEkT4C2YdvQtRmwDnu
w3wrWO8cIzkP5mwv2NWb2vpSIcAhi79B2ysintkfWgIgklXfpadpXUI3eWRehwJV
gfYSYvpDEQJsK5Llm3OI6s8N9V2W1clhXq3VYdJ5pk9SXkSL9xDPiDcTDowdQ5h6
mTvyDd+y+iEM1jJrlDXHg18hqumIHPZ5gOnR9Pozk35i3EArXS56hzuoBnXdE1vj
JJL6WBBv0jvDPuL6+5vm9dbygajNYRcUWEQWvJxnsjOmMNJU3QcUrFMg5rL+6vBV
B2/Mv/W5B3hg8plZd4qZQ/SFjNHPlm/90i8NIuqN3PTGGP53D5/eewryzBAb878k
mgIS9ahWH5JG3GX9AR+QXNNSIfgUfgJo2g17mSV3fbdUiqRiyeEdxiBhiKJTiPs0
Dr6Btn0uTGgjCabwRjR+EdZhTrfHkLcl0YBQYX3+Qexv/0ZM0ZrZVgwnXk1JJ8Xc
8nNUV6hVb40o/mKDAIJD+aXlZrN2tMZpRC4fY32dSVXZ7UUYtD6rfwXskmRcjPlu
Y2OkvJvjkEDzsphcNnRQJSMZdmRh2sklkkkwKY1ZuRSctSZripiLYU/GYTFeEkSd
d6B8xKJFKuRZvoIN2D3UiNyA3SfgLw+eJj0IeCkNBszsjq1ocBKdVjlnY/mJEmwt
whMAygqQ+EDXJGLQOdwcBwbpnMHynp8J0yPHCYW41ekmWlzsa7vAL9egvI4yaJDz
xZErcrQerYfri3hC0uvg/9CcEqLRXxm6ggxmFeFv9pRWK1kUSogoENGKBLw7R4mJ
r3+RwbrubKB9fz1iua13EGWW6EpunblIpZLMyQ2H9BkRkDApB0lfABhCyeHEOpIr
akTEguruPbwqw8IEZgFtk9RKPC/1d+W1mbsCP/W7j4YFZpPNksRWoAqiZHvqsIx4
asuY38sCynt6JHSfcMvmVq8PCjGM6GLzeMGQdkOKQxCxTnTAZkrxhYOV4lQad+i2
HXkkUSRVYIO093tLQV17XiA6WnGEFOX9D8CX+K8K4wfmZa+/RRTzG9O/TVtUGBl+
zwWxZa5HBG2CrTKz0ZVNNXhbyysZKmqWbvHgeWhuu7qPANyy+QdyJj/1/KMPqyRh
4/fsWCTEMeFIVr5o2wU2FGqyqkDkCtFYvW3abI2ZMBOSgW6uETvE7kBhH4i+eBNH
WKz9L9mO5+3r8KDikFOa6EjeNivuYEZNmAnSePb7wzbWaL/XIoHqQrIFqyCriXMY
ggqs2FSsXVKUtOzqRMrGJbUDIisu1a5uW94S+oHENRqauNtk4ojYX5hUQHWU7w1Y
D0aMap3OO8JY406QRsj4hVKOaHfQFH6mLpWFHvKBraRlIfVXJFvzaD5U3sJ29kZ8
cAhb/+gkidch/8CfPdVCOCiVTh5OjEBhYvJo+Jc2x8pRp+IgjFvYMQgNl+t1Twgs
kJk5c4m3hL5OoUAGEdsZCOkhzyoMO5r9vWTP1ew1GRFGCkhoTfoqe8I/Z2Fzq1ng
AlKS94j23K3ksrw47BhXIdYsBQn6CAhDp4Heo/bH3I4b5MrA7vlc5ZG61L2wamZE
KmFvoDBJYg9H4C6fQi8F/vQJh24sHT9njDjWAp1Di83y3PxPrKWJSTktDG0GeZBf
xCuYwYEMQpaFFrkpiLwcUOsW+EqWCxSzb5EInisE1SmwHG+hMKvkgU+2qkfnYBo0
/wzgnVjGldq2cRMCMFObgNwmDm5dQbx/xsVfpCsw8b1D327Bd4bItI33GNEa/ySy
P/5FMLwwj1Efg3n5Umi9JG5hsZ01B213Ho4WrZpLGjwXMwprioftQKJtKyRwogmr
azE2yGi2v0XpsAD1/FPkvg1kulrbX4VlU9CeJoefmpznLZXXswELED3amFMPiPFL
A1X18tpJtuqmP9QiOivLj2hOPMPhIqHnoYPg82aqMRj/0YToRR7GStxW4QGbK9Ys
LtAegVkhe4pwyHguBlYgF1ZoOJbs4XOSQDcOT5NwL92b+3bz/fTAvzm4Ok8R0aZU
IWgHLzLzgVhcQdPivnGJS3OAHf2ErtTrMiD3x5oHosWRlLSjx+Pkc0e5s8yyjQeK
W5HqpOuCJ9nc6BZbYOYqDnVicWi8rCiUHMIa3F/1cZYNo5LyjQ/x4IXl9Ajd7RRu
Y1HiOYDjVi/0S3uDdgQ78DUxXGcOpl5BU/ExvpXoukdHyXlFWUnpst0iegiGcsEb
p+e5by8lTR7XfEIQrAu6TAYe6zKbcaRe4PT8ZnCrp+92GgI8RaZF9Sdhad5iOZbq
CY8Pfz9vl0v/hRMtRKgw7O93ARJON0+9WrhH6B/Y8/P8e3liqTU6KS9s1sPgbxF6
RNG2MHLoyN5/omZELS4GKWR8dKLSSsL3aes3ukFPD/ePM2qxTnGSp4tuHTANs7pt
/+aYHrr5zmK8piB8mSvGM0JGBVlQq33ePEr3PYGZDAtIRfiUfXDE84OGruPyxS0g
AK+pqABJWqEO/of0zqcrAwPoIInm28d78KJKNeoi61KnBUMtUPOf3p+c3tvP0ZWW
0BHdj7MqTfnDVwrRWRY7FVYFPKAlBanAz0hsSfc4mcLOjL8R0QsLvp284aBSXSqA
tU+LXVJNGgIhvgNw/PBL4YdbM7hLdtLc1msFVjrFgs6g3wCRECZwq5vd6f+HipWz
lbu9yhM+tYRi3ghnj0a1HwkwAFwLj804dhsquYYfwQ/dFC86pSnJnmhK5l57MHui
IQCs28bbAY7wUBZsn8N7sWtelQ+y7gBXSyV32ltOfx+vIfxLsxFh3ZBXjQtnshtf
Akqm01h+XakEPMV7mbuQlkMfpViJHZgKxnMEXTM5/210u5DZOep2xahoOWtClrwc
UyMgk5AYU686OXq3LZzOOCzDy5CanAdcRx6AYq+Op+Bu1gsGe9AUFq6p38mo9qnW
VCLOaDjutwUBgCetqZtGJ3zPeYp4L5lyVahKnY3NHzb8z5pLKh9a1vMCr9oruIED
N8tEhZRhXvjLqjFNrsOkzBanLLpTCsMKoDkmfKf+uPDOJsjDu4YE6UWfpPs8+G2B
BqRLaACIVio8E+GAcfSPXQy3ZM+6tsAaQd6svUdRyuWxFjD2jd+zGtpWHJqBUmc7
GdLQopt4WhZB0USqM+UcvWZX2De23Pdxub/7gMohO1rnOTXPeH1JL95GEbSBNlTv
2TKtOzGQVt0F9fNglfUocJqwoXGOaIqKXaZai1+LxLcN9MIfmozh2R2YXZdhsJug
J9Spb79vhez1qY0ImNwoP9iRdDO1YUrSHnOraMB8/LNNgJkn8PzqzTEr67a28NXb
tnjBPzqBJArtl8suPDUBAdAkmvhZzxxQ4RsQXANEu2/cOizknBbuRWM5QT02L/9F
+ChPKwmkVoECG1yHfHvW5ng+2S4rHs8cAH0BAiYSNPEYq4oA9EKJSIOklqfgWkqq
ipPEcIJGBAr4Xugqn04PTk+G+0H0YBOfSYv41DodQdG2FNh/ZSxPzKN/1mhS1Frp
/VyhhfMn9FQg8dvsTPOLfDBmECVFxw1AAU3T7ICXgtisXqpInW5MIvTBVYAh70va
wplrVjmqBEvHenpKnz2dDoDkUiKm5JdDy84cHBJKbQ5tmbnOD8qtrdAejcyAO3Fx
QygXEEGoXGtsCy6l+jD+9gCpYQD0wATyrIFlH15qDMAIoAMxcXeRU5HwmRunlRTU
VCbdi3oQKw+e6zKYb6EgB50M4+n4QO5iObyAzEODcbLfKf2esoAXb+TeCgv6cTEr
v6h5cAFs3oYBF1gO5k8UbYY8Fdo2TISFVBhHuwQYA6n8lTBkKAjE8JQcMI4at4qi
4XL0XeXXR24AtTThoz+pClVLVwrSK0cmDo/wvFT/X6UyYOmoj3viRbtehzyNjHKH
HFzjPuizK7ehKFDjoR8zn3jZUaM0r7gJhJwrJfcaH660l90e/YvWqZT6VQtC/8Qk
1+06nlObKHrw51kqIy6wECBhxwTi8uPSrV39e1EJmfMJQZ82R1wyZfOTJpr0asJx
GIoBgXbHbemXvVtBtQazBXUuiF4d0R031KDe7rwwMxfUjhy75N4sW9/eAxDpD5YM
E/o8SuajN77mNY2YA/fJKDCd8kY8JzTiJXsZN6epxMaGfaX0SXHTuEaq0PErMI8/
7TCJrc89b3vALYZk39LuixOz7f1uGwa6Rk+plSWJPZkPQkfnzUivi89DubYiQJAS
hCpU08AKM8Ouli3Inc5L+dV2ajGtKygDSAwUelk3ntWcZ3Vx/FavwzZH7ap5jpFf
k9ZLGxMx1W47jWD9qGa/E/ob9V0TDARZ8FZDk/nnExAhV5DkoH/kxMK/P6dZDICb
+FB9qM7t9bmfLJADDzEnwgXJ5Tv3kEkpwtivfa0DgdJvO/IRIoMQ/5YO/19H6SWO
6kJh6MJecklr6k7t8zwtxfELOECsGHh5MQW7v/3e5Kj+4u71qKcQ3cg2/3+7tdVL
5riuLFOHF7wkk8ltmDVpHJTTT24HpjckOAAOdU+cGhX3peR/QwEOXPMMdNIaWbKJ
S/lmDlEvKJTcWCfdDM/PGFoz5QOyg1pGsvoHpY5RN4S7C9INmzanU/pqNyn5UlR7
hM9oabZ74qnnEc9cJNPvUxSgN3Fq3fSnfjRbdIcxqskKqvbiKAQ5BRZtlYzbmcXf
oKgO5N+qsIVWraRnhUa7cQEgbjwAwIQTC6Yjegs2c8QbkCnMUvng7pFVeWPziS27
yc+NrAZ7yUmm0acQsWWljKBtkdDmO7aoIiSn1bOOoNHcdzeP3JZb5Gw41RoNJ5/7
5+dnBOxxg887aIFU3SSAEH+6tgHKuO/7ZrMgX2jfosP7iWaQ974RXg3Bd1Ow+4qT
Bi2otxYQVocl+Rx9GH8SEllWcC1cJbW7nvh22yTUkK7u78cZHFra9HTKNw10l8xu
QOstIXZcLTJOoGfIK80hZjFl5keUHIslGif8BXXSmbo3SPiI66cSgvwRRXzQU4Dk
xN851DcdBIV0TcmzDeYbJLUtSEw9yVgQoohCZ6uGbAnGHkDbsEbpM6mBGdArhUsp
SBD2ZGNpqr45rR+JjqLwqF5FAafp+gEsjJx/ISI8OyVOHKdryaZTicw/5XJ1AG7j
pFJXlgJQ49nHz3PaBYFc//wkBTLCA/aAbI+H30EAJ3ekssoAqCJyERvAxrA2sQMP
Lv2GXenDG/K2IVlW6cJa5Tv+SMOfPXPiL40GoP3ZNKW/4GZ0UY3W1XlxQepJwSzD
/nkgAP2tLDLkKs4xoCmW2TSagvXUgD/gvt6IrNpccq72A9aNtQ9B1+QplosClo3j
8NmpY8IjsDyzVtWxzFqgcNB2RslMSGPPEQLFxVjdvm9LVq8+Aexnh0irUTxFtWP3
pz6o+mbCCt398f5ECSJ/vt6jGF2e+W5Mt2mFfDXlDWpTA4kFcui6oJBKBcpFHHSF
o85KOccXEvqkdtRImNA0JsSy9jyxkoq2rrKrT40mjCdzDb0CwNNyEai813DBo5WB
7TLqUYyPphxbSMaSoAIamZaEXfFcjowiGzXYXA2cGBB59InWHr1yDG/6kM1ThPTq
VQsqhDGKCfr31gzOGyNSWVLMdYuVIk3akCW/EiPVoamSXH8/4lkcqBV4XipbUhXp
6CqdfmnqY3MKVfVL5QkXf+XCf2KNsdwvj3CnjQgCrR9g/7tJyGWb0PthyiAxF3hs
EPutY0ThDlaLhCSK9oCBOk/flk7eRWsiEMQ9GPxVf9Spiv+40O5bOaZVPWey6uZ1
vulDOTZawvxu1xLLwPwh+eLJNFxG+qozMFSbFwKshOtfEbWZ8T5nMHV3/KV0ZMWO
XX6uVfth0+uQpMatBPnhWhqPgdJrh4xWCKB0CGXJ0chZuV0xPySnZA3WB/wR//wj
nWfczbkNUCuer681B2tDCQQ7BL9Nw0Yih3NJHvVjmVbxhSAFWt4f16zxq/f6ZNpq
1mZZ5jq//pwn+/1pfkRfI4npXUgMAYzJGgIOj3d6Et+LVNgx5+AZkaUcjdSYMOZH
fxeeyhTaHJenxnwaIeNWTHp3MIm9kQNWwiNlsridNQYojM3YhJZq1gxBc3kGumb3
im6/BCFeRiL753Le1SjOXWIYyaSaZz5Dko8wg1axTQ2eojNNBgDlIZ82QX9Y5Zdj
HDCARWSOAmKSvoWfStgJbq4xrcDy/nojKCPDSB6ZdpQBagqXVqDthZmwkRiOmEfU
l7PANoV4my1Gj8/QKxMUOleRMmSE7IU5hqfQUt8ws3UpwE61ujVBVCk0nwo0BxyT
3YaulWLxlZInp2ctnA2AVW+IJVX7NAzpid2ncrueIm/kpUckW6+xnBTGZZb5SZLF
ZewbWO8W2KoTPZvzXFTNEDyfR65xwAOcXbCNxqVGhark8Erv7tXlNevRp3AISnl6
o1rT4z5IJ8Grffo5cyEaFxtmQWjTzZ07LBf0CklaeXZ8XACTlXLEYWKKqN7qCV+T
oGINJZVcHJ5W0xdlixpTFSSosLWNn4RapMAWe1fMAoLbeSunf1bESNWcvm77MxWB
6M+5wDMoHkgNPm1uTJqRTWKxw4tl70qCoQ/CA6nqoIBKnEZYC6Ngzr6l6MMUU3YY
0ajWcYcgyIkaNCPMyRp3ALo9kAOX5evG1tmevwlJgPgCsGJXMZMa7ptvoJUMX67A
II/TD2L/jS4vQGVWKBMjfpjdm1Dr1ESBTWle0b6pEnyPI7EE2+DP41YmdvLhLGD5
bU0uOEMugaidhaBIr5mlrA6QV/SblVw+SO8woNQjo1BgnB3rxg2+Dfn/WyfAHPV8
nGjqQg+TypCSUWxZJ6yXBg9HfoRIl5+rhh/C/Rs4YuRY0jCwOWSFMRHa5M0ITwyL
HVA7AFWd8jc+hw57UlIgSRyhMqpvj7LK+ciDBtMlJjcwTkh/soeWxGALVqCJd60t
uPYWMO1uxt6Owsqfhjt/A/OtwHctoMxCsAlHuJ3H4S0Eb7o47z5SB1O1v4/LY6z0
lmPM6y+T1sf/5cQjXNDdwNKyK6boSZnvhwTRX/dkZ+NA43YMlumNhbgamaZ3+dIw
8t0VLboFnKuATgMSSVsj6OlgMxKgMouC8Vhl9uTPg3EwsQt+9fc86EzhWgeQ/Ula
Igw5Gx/cLnDIq0jAbZ5gnABcS9eELw3KQ44gt9wrTB7MeOs/GB28eTszbbQoHNkN
vKz2n71K6rbk7yCNNwoq2votN7SnlAZ7VW2+fpa8btQde0yVRK6qc3kr1TQFu/xp
0KO7ihgKsVq5FjeMHZmItq7Rd+yXmVMsv+dJkU6scqNrxnCKaAr6f/52/e8i9e0c
ENxGXmlbnFc3chv9SSes3gN9vyu2qFvMaLOOQF83oqYHnOqzL/Nhgtpv2FXRIyUK
JWjiKj2wIISVNERn94D3JMEw7C2ipaNVmeWIbwlELTpZSoBTPgXLIA+TUtdYwbtB
TcGnPe5ynHgEl46qRH6ZcIgDSU0vExZ0n82svFa7A9R7G+1RVU4JJPtG/JbjUsTG
NTb1ZWuR2Nkhc7QU2AlTNiaWNioagu23/ekOE4+tN0u/6MM/l+80068vwlDMOy9+
2QZmYiIcj6OBjOnO6Q1cc4t9s+HuQCUOBSXznCIW+IttAMHtD1Kt8/4nfrSv4HlD
TWR8RlBugjUvMJ7i/TuLGUYeZN1OhePohzJ+ADsr70mRR1YHw5b2q4N2UIZcYhoY
+WFRqOldtrN/OaUvLsZVX4YXCQB0N+Ka5/DGiaz5LasTj2zY1iqNo6dHjH6nJnrF
cUhn4cJK/bnRaIpZyG1cu8IbrKDoiGKvv+S1s7R801qMfggjVbnG5+l9087JCaU6
rWxwHP0jfLY+3L0X+4301te+VWzm2HcCUuvMq+bmkAf0Pmt80IEZ23FpDRVH/lL+
frXTCnZXfQE1lAHeA/uxK4cjYJQlrxDPeE78JfYD58wjbkW4RNObTzjXEjCAO4/c
rh2W/P9WAUNLYviP+1on2U09p4Kv9m0gMQC+c09eqP9NKGoS+p20zYNKgmRK9I5q
4f+kEAsUEkJRKMxzemQUkyEkuLDVvTVlPZIH+MnYLCZ6B1ZFfLIiEkW6vZV+4HPw
e7AXECS9w0NAvDLPhnszSDuAt7JacoeSL5z9PPz1XZD2lbt6hh4T+MBv6k0UkRPR
v5KioBi8ULnZd+T3F/Srr60ka0amtTuSaq6lOsV1Gmy2bBcbQ+exfeqlnbP0/f67
V6W1RyF2GOrJOXJBhBsi7hVHT7K7EpmPgl1iEvjXNrasYivGW5pOfS26UpboFN30
tmIDqQeL/8mll5F7sl+U8cjdRzKu5GKXnx/W5vv+j6TsjIpM0B9f/9IxQK8HzdRS
dmNWnVvpzEmzwh2vlPZk2HOxKeJk8QyG7aobjiHt8pEdPtbJ1cNB4njJe82NpA19
DtAeFPVBhDwzZ3R7VRdXBdRgvQN4xiJl7FUa2p1OdlCztQ21fnmWhGK4yiYZeV4c
yHndTNz/AzMl+UibqZuUGwT8r5afDwS2FvmHf1kIddS/7ogE5ljSrykmciBRer31
FFd/txRLUi9g9hkrfapZLxBRUmz+7TCMInbabrYdEpSUaZ4kIq++xPl1TmArMaFV
cNnTSp402UhjNgvDkUkPh1hsI/VdDCIkON1g9iUsVpVLcmA63K5u9AP6/PpYm5yE
RW9BBVifUOmHQH8sUOg/Gonxhg0gatdIGxXCPUviWzjxSbiAeFmB6/Ct0Hp/zwX0
WpQ/FKPwB2xPdvFOyMQDphwGmZ2ge9wqOnkO3PX1sGS3mX5EAs6Mleo1BafSrz3j
tXeFn1Mjx5Au2g+XNVWKG7I0EBbpQjX3lH9HYH6HYG0nLeEEoAsXv3QlMRy2/TwV
syYouiuWc0wsitUngVwxHMhmDJlIG6dsowBKoHAKHcfiJxdm+udv1X3+iNx1uNkI
eThdnYMHkuKyWLqKtocGIUt0HGy3bfxaRVW6iJD8HXMgQ2WPMByRWsRkZdILk34G
RRGXm4jN8k7rqnv8vFY4Fdhpi2H1uwpYLB4RdZF2ejeLMRJRG4VdMy3GtqNm0sHK
jPftdtxOwIXy9HfY7RhIEnO//6+YQqqP9TB9pZrmkp4plp9iVO6yGqfF8koQNsTn
EDk9bC9lpofgoqFEt/lYjKEYp2jXFWQ8z0/LaVx74dUsegrVckt149GCDuogHcJ7
fM0AYQHB2CMkRqyu5/ch2NMeorS5gBXbyOQjz3G1VuOdRmv/eL3O7hqbUZVlr8VD
Gh+zb32mBE0QRPzhbUR5VTfPlwc17REoxdeCzsRq5UVXrvOQY05d4HybkEKGlN22
/g9BcKWzNeFdVlYU/LHITnML/WW4V3mx1Vw/JHi+IsaMhwPa2nSWeMbxFgK5sZ4K
UtfaAgn8+x4/03ZS/RSxcA8k6J5X0xaiwgeL0h2/ijV1l4ne7jZP9PhIDe7S7wJs
+fQK3fvycF3sfWcq8VgPFBLfKrcJTukCTHVJD+BXzykHv47ytnF8PIYgiU1/Zg9+
Kxa2IbV7ufxtnmslRowW7xfqug4qI2+PJ/D9HGru7SWaPXp5c2COLvGPrfbJG58Z
89nIIl3EaVdw36u52PeLnzQm3XaGNIIraKga+/F2PTdXSRlek9DtNubN1m4gxpfp
KVBP/T/iuGXBfWzXXCYeleOwswh+FEZ+cx8Uq4aY2lI3t2atVo4fDZVPf9WL8EM/
aUrJNl9BS63fwj3jwXnpOZp+lnJDjUMHvavWgtRo/tLXojQNT+95bw0AJC5Vxy5T
+wcc4Z9rY//8YfNUyXeOkxolbj5w52AStV8S8DDnZ270Y+2NFnv87IyyXSL7ZvTE
O3cp7b9PQs/pV+0sWw0r0rbNUrFDhXe8oHykvnxtm+zy+e8NsGFz/2U7RK0stgEG
6MQuaxenbpC+uzD6MGiNbfmJfVaKE4eCRKUTCuj5rM/RKhSzjR7NKBg67yXMdemC
YkdZqi8PHDhLw0KQyE2dbcIrIXcen7KvMGGy2ZepDc1Qtwkg6IXVtzFpyOfLyEjR
DZlOb1vaV1DATHHt8MLCd1lfsPGncqfTY/P3jvgAh5vWisuAW3suq0Hxc4dxehWp
wLkG6y2hTC9CMHVn2ZQTenNXnw7LpXsZleLxR5fhFuX4iS2c2HJb7MZxY6Q4gy6M
b97bHda56leHtC24JEJUSb8uFoqzZwRb/C687Co9ZKzMEAdv7mw0wU1uoq7NG+GV
+Dxtqon+Qsr+FsJzLGnTz/GmcFhvuNtAoxTWsHg5WH8d5j4SYR3eHlxPES4DJC7D
/XbnUzX5MpUo9MTYkhAvGac6CcF8NGfRrbGYTLktXXhCD2F8YtpGYV+Xsvsyx2cD
BEh1NAIy0yQpo7CXFNH5ULe9zQfssT/kRiWkxAnhU80DX3JGDplcY+Vlb7qI0o/X
IeaSpxMGdqVUshwk0vVwQIrvSjjm4QruqSAnQHLfItCjv4ETpNoL0yRYG10LnEV9
q+JpzZo6E5TeNuAX33yLp03lPkz93tnvsufZbf8a2i5up4GTG7clqDbcCAzx4SSm
6Gnl+VzlsEyn3Op9a81AyhmGwRt3DocoXm5mv6SmO9wPl6j4uJXIHWajSL/0d13T
P8ktTmuegDtlukoxiURNYq35jfx9Kd+KZ/YVC19yOQ1ipB7VIHDfC5ZaC7T04s6z
do/kLO0c8s1kO9yBbOFirIVGpXuoFTSnJyCheA5gfmThfxB8wO6BH95rHqGoPgXY
WTyUz4BakV+Yd8TgeRh8p3NDKSoT3ocM+n8vitEwPLKyMGPS4JP/SkYJ6yXyN2Cy
uPQJGfqLsNhiJMBOInQ+h3/EF/RpV0aGu70bhCE3G99XUn1ZJtZccqRLroRXErpl
XmOONr819h8saWyWMLOkiTABfJVlSoIk7TtMAABtio8javLBy0dwtrWQspcXCJDN
JhwSUxTmrLB/AioMnjipTZB55NI19QUtOZrpTOXH9qG8Vqd4j/7orZtO0oYfkZ8A
d8yqja6ULqcIdfEdCSZAt8t4GJ3WZaok+WJS/7GF2i3ysAN2YZOFpxAMZwiI5eCQ
ib3a6SS7AW9toW4qRbYJe0cd9zekjl2t944PieLowWNgYO32cM7vRgikvNL9L02+
slTIdR3wxg107dcm8dzxnA7E6at5lKYkcT69bxdbjxXS2YMrYxWJhi3OAC3xMG3+
K2zSM1c6/kC+ojuxVwBH4InGEvvHR/vyZIcgjcDORP9YoxK1bbqTkvnTw3izechf
y5RRv3zK4HopXUGVpeoOrps3UEC2b6sf6ECkCZkwx3LmQ5ZrPVR41g1rRJKKwj4E
ar76Vz9fDX5RJSTx1KtUOJbSOxnQ5G9XWcwFxMqbZuI1FK6PGH/+7p0wqaWyaa+q
M7yGPGCeJzQXzGA0rxSJl68HeemRIDMOx2747NnIfA5kVSdYYDI9MGETeJuZEcIX
2BLHem7No6B4bm96xNPb8xy4TidJxHxp/G6tDmlx+nHws2W0fga8Dc5CeVnaiGVx
AfaZ8HAXbcDuUUbx4EK9wIY9b8ui12/afSAdjUzcGwEXOiUynAUT3jEnLiFoJfnk
AHMEhbxbul/WgdrorX5Fx+NMCKNjtWFKjZ6J1hmoKgMT4mvTX5JeyBYFB5hwz6jG
FoMt2wb+k1yIMvSO5rvbENR4Oj7SB7W0wQ6+a8ifPaK5gb0VpKaYlOTS16o/rmbl
xLPQHXeycwZQq9BYEYXbk5N6OOIjpnp5HOGHOcDRIT1hhlNPxmAawrzbww0ClMsr
1tF78Zjpi+8jjCgg2sCx4zhCeYKxxF5JjZP0bf3ocJdZhwpmRHfkZ17pUrTTCcrQ
TnJepswDeJ/9NW1/x6BVijYayGlBmYJ8hpciOWtx8Sp8tvxT6Xh3DD8Bn6ruFnEQ
hnpDgrhsQr2PQInvZZPzBSriWh1j/r31YpCjCsLVR1i8bUvVLwByKV7CdudM5jbN
ClCrBvMalPNiVkSzjT3PbCiJ702DeG2BP9fg9+PflBD5zDy1DJl8PZvYKTBj9wFm
uxF77Bh031SsqyVJhNDRCrv1jS9ZNKdxmUCn/UjHELj3lG/RtVJadTCCM3L6CbYx
3mpGodx+imvLyVWl3aaYQspkPsp+pkkpi6S7yDKFnftNTIzqgrzf91rdl4HnlTXw
mRrX6tceRTeX0FAoJbGBoSdd7nuBaVztEzj497dVcWRILlUxaxfi2gdetZQ/Po5n
pJTwGl0jA8GcrUrnDSSFr1UsdTbjM66rWiFtimDATy8uNkR1OnTNpVUI+pfakWbf
upYf58fPJmLkKJ6VHGGgKzh3EcRT0EQAkOgqcygh5vvTIZaA08vzYUCcIDDFUzCW
3MfD65/1sxztF3GqAoFt18YbynHn6gNuygSD5HwVHEahStew1vaA2yFvbz950kqE
qghCrQmFCr101V7sWDpzqwfTMw0yX5oi2bhYpn92KpBFVeiMR4TS8qjCJHxzMpXe
SU9/l0EM3dFVBe2RokyCXMUAYF97NEYZreSc2Tc82FxmAK4O6W1ITovCFGW5REel
YsYx4FDQ5Ab3dw4dj8fJq2oMywjd14yofQIR6OFvFwZQyWCL5H1ABnyqu7BQkgAG
Cyi9uWWa7uWATwjvgm5aKjzgWGg/iFgGh8w2AsxynBkMvVQkPoMZo/u4o7mZBMtx
Ra3QPxbdi4NVdkLcnuczT9bhWFZIN/pT35FQeg1BAsX5OzlQ905N9vleN5WbtQ9R
QRYbP5/FhNEzqLAWlHF9EmbFLFNr14526LVmhrTp/BGfAPFP4CzmmBYWTyKClooU
x+4Vy5+5o9OfufgF91NTLSy+5y66nAQH+EAxkfI3em0PTSmrH2ZsmDOh5s/uIHES
vzKcQurFFmFzhazTxVBboMOCBWAa3KlRjvScK2e+dVxtRIFcoD0O+1Y8HvN18lAw
N6R4bMW8qaPn5hPYafAIeRsHiB/ulSw701iweps+EUDki5BYzpKtsE6pOAct2CIs
ER6IDFD0kBvB9eRKjjHjF9FgYf16N7QFCWexH/wDRAWe3xIG9lfX1zuqUrPQds+c
eCR8sIZJ+TqnGR4G4qIISEbBKSl61tDdS3wQ2Pt+i+ZeV7lzs/BpqwqfJphhtRkV
IfduVx90XWhni31Omp7M6z3AcXJiO67BYeWO84xAsVDnoTlQSOD/Y0AmyaWxJiqT
2z4ukFZzhtkEUmuELgMttLlLqiNaXOef0cRGxaALDcP1kJ7sQ6nFlsndsgB0JOde
I0/3Ck0Bpjtc3v0RfhwYupqCX6n1BidSwP2B6RfysrlgY/M9/IkfCvDfjDMUUr9o
yyvKrxAmdOxqDYcI4EtdE8QuYVPhNlF/jUnE0B8fhh1WZH/Vezb4GmwKCZjd936N
usue49qxvYNHx6Qce+QP35wrnGSTfO3VRkv9+mjxod/mcu7nwwi3H6tQnKUG4BDu
P4sHEmpRCzNruc3iF6z7qARCv7ldZ9sBs+SYC+i32Pnaw3LqmbGxEAMt0puy8VhI
ip/HlsuC6j7Ruw7JStsYjJkORmvnXWiYQ2mWfC4dI8p28hHWCdEVrwkyzErd1QMS
QgOyanPuCmxQJ55unmM20WusZNgWUPKpK+gPQ+BGDVlZMej+kRdhvWEHS2GobI2S
YYo+6ejH+FfdTfQf/yYP0C+LAR4E7mHUZJTOLhp5ydENFfqzm64XSL3NdOl1q1jx
qBSNFI0Tcc6y8qMcVzueV2R677H0n8Ls2gzEmeQm0Vobv6NWyCpYMqM8q1Xtw1FJ
gYRUxXizTyqgy21tH4MoeynkoYP9kWN/1Eov40ywSKgmLVVGnsr4tJiHfw7ah/i/
vLolU9MfB8TTaEoyX3kXRMyhsxmn415xeqB9TU5QGSwtdw1dcULHV3t5EmvFi6FK
9LyaDJan0FOlWuOKKfuLfOua1NtFytFi+pyyAIuz5N6iQgKric4B2yAVA/gGK4RU
Wk+JuLVMFccilx/kUnitTx+azdiP24jAvURoR2Eff1qpvXaO9qdoaitpBdjZE0lI
pxegAuva7QdWOaHlh8+6OcBQSCMG6KUi9VoCn1bbeO1Oikuk53SCb7a7M6i8ra0x
27GeaIQxISSnTCW6Kl1tvWpPmxzQUlfDMRFxbC2ImAk52xY9TLiEw4PG/VJR6zbz
92a7LnyM6U4x+64mq143k35CCyyeIlpIsGFZsYSYbHjGDV5UNyRx8fBBiAlZM6XQ
DuEEZeeLOmVzfCcvsgaWFuKRTyoDZN2fJhCcJm0DkFKQC6nWN1V5IXjxxnSCE5Gz
0JgrH81hBKAblFQX+Engnue9a9vnqj7NK5wSAbm4E1m3s86SRca1TRd8AmFsFXsF
20umPZnnxGHwzag/51+uXQGwxUsMof0TV4MGXW3+6yorvnbrl1DlOwJX0O2hJm79
JH1NPIc2lap+BW28fiO3KtFJhT23tnlDgwf4W+UZRGXlJHLmDMSz3UwijaI9GdoZ
XRXGB1nyJJCs0WbRawHKJVlp3+mRhSjmQZ33GyI5rvHn+rg3usMNsZXw7iLyPw7y
ND7fJEp8EygoLnODugvmimivwiPZPcnHTU3+HEvgKRbRZTCrJpWnX9dO9yoisJ0D
7cZ+BYuRE3bnnKLhX8JFK3JNmlAggTq7BFbdlnpYD7LbYmV+0R8rVGpJQaFowBSH
OmCiX9CsCZcnU8Hb+Pei9gW1PulcX5JjMruluL+asZ2w4+1pdhuDmbEmYq3yuJs4
BJ4okPIjxQygxTHYOAnxGCL4j845RHK0UuQN85e6A97k1C/uh5FCdgNx7dqAK5HM
HdmcZ8+AL5lUMErfdzai1ji4jcpFMtAqKgX2+RvAy1pNUT7NhIP1JMlBWnGLmEGr
bK5nMc8iVVPZpL8ISw+aH/fxoFk0DffX4XTU6J6eZgZMLB+L/CXU0gkJb06aXXtQ
cOoaLYww/cCIntvd7AiBnHHjXW27xf03nyCkZ5q7a9fdNL7FKoBc7jr4x1IQyN0x
6vMMK/bBTa5eibKeGp33a16OGMsPPL5jaLmPtZdiCwf4dwN2AdHcDxag5cOleIxz
Bld4U8uIcTmK9sljaa6RBKx5SF/pxnwTgWTggw4OGVx2aePszPxDSUoUIIo8DihQ
AIWSxB3dY56XzceVGnPihJIk58lwog5EunD1VjNJEw+/39KLvMJsWy3jveAIiFgq
oLBe+dHeLtpP2H1HsOmxQAiY7VyCK0F9FsWVuNqKfM7ViGbB7cu2fzMwoQsHt8sW
NwLQhotUe+6l4fMUPpeL5cftb1wNjhe345R4zsqXtMM/ajp15rp+Y7Gxpqc/u8yG
6O+AlPdM4SVRtmIU0kFZ+dz0YuSWp1pD9GstiMVP4uR5SWpvwqc0GcPR5cUiQWFZ
RKCI8iAACchoPH0Qfod3t1V2u8ajLTRUaHy6RB8TLRKIlHVsEQnDzX6dNnDYKNfj
FBay2GsPX+X8m/eOzpcn33FnLEhV5h+KuYGw6pviGEpQ0rIXYRE0oFOj9Rd/C5Sw
ah0NgJ4XDadR/rUGrEwSVtLlqAnunC/ptfxwoWM8DFGanH0NRMmzHLJIX6nUaUrK
NoMYXFtWi1ClnXJ+oYFzhyB+0E9mW+in7rvqXsKRAs6Jjv1Mrgy/cC5RcFejxRdh
bjhTLMRCMDnhPSmeZ/1byZ86ZPX7KBNTczqxrlLnsYlS/thw79T7jAwfVvYzxcpn
ibsC5iyiRHo3IOJWyIxZGrxZMGUofPsLz+zmY3iLYPfuq6xHXhmIPs5h+nNka5za
ejIAqK0OKJY7xQ1ck0PjhxQuF17dJ1R6rpKCLXaCamGC9a0zz/xnhgukvZKZjL5N
4u/x+W4vijkSKDly1oq7Pn8ypVQryM5v9hH9OrYWA4tZR/x+8nT8x4CprWriPztt
cBHxz2pBPwOpT8KETj9baORpvW1LUf9tn8ok5QufWZhHK9uBzYK0kCifYwu51mJs
V6KETRzKtIZ7tlbUk1eTbaZd/21dXTL9D0gHOoP/IrX2WwUSVzd94SAhyL5LwfAz
QonRLaw5dbLCs9cb6RptUHmOkGDkpjnKV0eibzItgN3JBlhKfSYxrs1V4kKbMf8z
3nxxdYFRfMdcXGxkaO9YFvFvZOSgE5Np7eyiA4ecBUc4OpAt0TJThtsRdOFy7f6z
mX9cZZhyvOyrT/GmC3rcNYJA2+f9YmjDZ7qYhaIzUjlV0ogSDoXoZSrX3dQB+Bke
J8pDT894LTARFznosAFfPwXwppt8NrqCIGODOnCVz2e/I7FCCaiQqRsTGd4UD4iD
MQGhyMcZNn9H3ID5QAZ/LMyBG1RSe6rfJm4glx9OC1gAi7R7/eutNv0yL6OYTYET
hm1Hyp1Xkpsk/6Ded2wQLfiakbzPx+kVPSfLbA+E3lulbytOMwySInoMG2yxOjB6
9c1kvuh9nUCm8Sm+ga6iOB3QvQoGX3Cl1jlFJ1Np+Jn6AtAMqNdFp3Pl3SJcO+1E
qhy/eqRMKvyjXcL7/bFddFjdZX6jyoeGaee1ki6b7TNQ4TofObZoAFGSvg2zexfp
Xun8YHinXcBelftGK3xWjLMCWS/F+jobmwSxvaFPROWk8H8suiyegmfBX6mipxpC
eykoGBxNkEpuuPRuLzDnf8hihYa8gzChTBT2A+3DpmiK4ZJuS9FRt0Jl0HnwM+0a
fzgomuhd779VZX6t+t46MPJ05xqw5X59H9wM0aAX7sPL9WP4u0msPG6B+rmSSgTS
D4L0g2EyIYbQUv99zcI688mN8FyXyERQAd2WHnlwavuZF5EeVPhJN/FWDDnrOFW/
LwmRoQTiS1JhZXBwZkknsZC0Xg/KQ49Iq4dBqtNlLJyB2ikH4n338AHfwY+zoKtg
fd65ol8XJjpas2PaPh4mKztx29AAWdiykEE3yKqVCmGC0UDgeDqTa5S0AWMmq3dJ
bvh2ZV5TpRYNje1kG6t4iRMho3kwvBlSlj2DTaw54IrhmaI4/yw4Y5P8SPSfNTrA
wHcVQvDWvWLREfho10EeA1XwXsWeC11+gJEAF749xiyrdKGA3GvBmeGWsXGvonAn
3fuxwUEXgUZFQrZgWvUsKtXX3kXJxzAKW/mfAKbbnjvixGoMTw39z9RM/WUbJdnG
YFd6Jo7EOgTzZOmqgtzWo//sPhFNn95TMRbMomn2GMUjX2teiKon0S6VT8SgG9H+
kYGoI/Fxb+r4v3nMH24XTf1GtvaRsHEIlU6XK+opEECAzEsGU2H1ckVL9PqHCCmP
gd9xgrfMl3ZM1s3toPoxJtmXb7HtXuDmMTjnYx7eXhAxLNZugLZydr51mRZzCBIm
KOCgTNR48Pd+mixXeLCwZuAJdEizOLxZijgjIIreg1fgObGth/DJDhGTA7v1oduh
VXqk0fJB7KGsPHeIkdZ2GM+qHxyWeCr/jFEHNe1cjWpBAvvlT0OsRNE1LpgFBxXi
0v3VmJ9RXcTh0JuYHbzcOvEXNyJqqiro046IOp6nS1X5DnKWXQC/UNxeSsj9EbHl
+kvlB1rMOb2W5aWq1Cd8Jab2PUNWNaRmv8hg1EV5QAhEk0KSVJen7eUkzGQhGrkl
n/qigyte7tXZrE9IbOi81exrZ6/a87Oxh48Snd6R7SmyKRgou/Bgm0NQjTTAMaKI
5GHnrKuaBA6+NDJxEg9AeRNlXvv7WLbc4uRHCZSa9YJj6kOrl4zjSE+cZiszlx93
2Z5HJhK+HQ8vhn96Mmp2kHYSULYeK/G/xR97vRjwxIrCs1nlohsZHk/lv0rkvnGB
nRRWXc2cFW0sE8D18c6AWhdhq3MrNmaOYdneFgDYWoJ7gTM+bXehnaQZwgfZdSjJ
dbm/4aVBGKWaAdULU3VtvNd8FxEdVkdCl1YpQYkydmD5d6dNFKH8Dj2P7ddvJBfD
YdPqW9z+fYp2CVUMiI20BZZFpEY+wVHsobDR3Dy+uLVazKsLFOYocTtO2l1Uv5Zm
1K6SBx7LEZeznAH0uRvotajMcGO+JAzeNtLighqM+hbxP88+CnP1bcazyFHHTUXt
GGuE5cW6TzhszeMdZtAPucD1Ms826c6ZasRFxrOdM5VcKPvGck8PgMVfR6EQUCcf
u4nVnvYGTHRMJrcKK2Bxps1IOvEWfSjaSrhX2hpdNR55o6MViDGvJRC4Qsaago4m
4n6WinfP/ttOQntM7Ejg5rqkmsp1lkHT841YEM08Q1mBSvowyewUdGUPFhB7+W61
ZgJCE79EXuOoKmGTEWKeanFe2o7VG6RprfEF00xTl62+d/XDbPD5tYn+HHUyU6S6
Y8xKLO45MzB2WBBXROTOlKPb73pcgrA5BhsfeeVv2D4Cc9ze1X9HC2g8aC+PPPEj
fo9tu/yTiWGb8KOGhE4hbIN2c7KeegBwaXKqfSQvYZRZbN1exBzIfypA+ARIPoSc
8RB6ZxPL9pOw8zeKb6vmYH1BWMeYcaPHKjU5DIOMcgPTjuU9UAKxKf6JEbELtyZm
FIf2dx5TtuZe6cbT3V1bTZr00V9K7wKTaccoXtOSftIVYq/7usbkZx9WzaX1LxuN
fA+OFuZN7ysVA228IN3d50ViqEBSrqOSVeoJSIBVfbjqJSCPzcaPU1NU6SAY6FqF
fYLB+lF/kGIxbIvdFeL+QbEQdy95GciOb5l8SFgdeG/sIAIi0UUpoYrWMSja0grx
5EKoAm3R6LrdX+JNBxHVOrdNU2TFZXZRgs4cvc0SakGBuLx/YJlFOdTb6caHe2bU
bJ+IpLQw+n58y+DsHarVeJ2ekyZ+1ocuwZgeNYO3bB6uRiPT6J45LnHUhMJGkelN
LLndIPsFbVIZ2LjU/02Tm/YUQymItTKYjjCaBSQ7+IQEz/4zkTNVz7RjcK9QGDsn
2eGbT+4VE7q3y2NhsfZka2F+VQ27qgBVTyLw4vxtnxWLHNTWBaITtZ+9nHAqkVSD
xfY5bD5cPeo8BTldnSA8Mw2rRJ+rlAMqT4z8GocCrgUGFh9y1KoiWiutNaKKfjpo
RY9XOSJIeMhfgEgVt/1i0n8un3JGNWgIsOAviMSlIkTn3nLSn/NJnxF01rtP4MK4
6L3AtK2/Hu+O9JdFL/qOKl0yOS+8om4w4TnQiexhLi7kc/RVpqcphezCfZQxOoFe
MgxTA+9En3VD8DZracY5Ujjc5jAh4UFsI2mkUeB0KhmvsICX3nWmBjvPb1+swLlo
7662XlarGUIXnAteOpccdQ7uVfHZtCgE5YNt7XxQ2Bgx0PZatT+R7MB5O2pXskZt
DVyRgEonwL6AxYktcTmO3gv21PKfk62mm+aVbbDoh7YVN9OVkNWmcSyBQJCTN2Y4
nFn5fVrsmP5gXQxrQNnwFaCvbNB/luWSvss2uuXbhYoCrOqOAjq15twGka/ZGKnk
Ryan3r3SFR9LQ3ngbcsRWZS3472EFMWoWjaMjfG6tDf3NgiTvKvhexy1Y7ZQutEH
LhTr86/ckfgRG3ePR1lMZVCaSYWC9WKKYREGLZIXERS0NeU3TiJjEPrB3ZuZ3mVZ
iaYM9V8bSKiti2/6pQIQWiqfgzF3NuAxwOaxun0BjJqIJ0ShLRAwQvnAIoHUvIPL
XKeoMAzWsS/QXYyIn7UCEQI6SK7VcWrXTahL2T8rCUr073wzY+2Qv3bq6uYorVjE
1rz9zSVrmqOitQU0NM0LLTGIAVIMDuh6ZlHPELzgTJKVIFjyHYPAZHAcUqOB1JN8
7FqwizkdnsxV+U5YH7qnBKx/8jWUHvcZ4YR3Xll71TAl7ZInn3G83Ip6xJ7hJWCv
TBQypI5l9jDCqPToGDFZ4ELxdfXzRabwgysqLNV4L4gsK2t7sXxgbRJxoXi2TSRF
C9IcO9T8385fpUTcFeuM6EV8kqYsuUTJwDk/Ln72ZV8mPJSi5wnVC489zS2SRYo2
qAa3NINaNUIKGA7GI7ZYIejmOHgrYvTelFCRCoK/rlmNoYu/CWbTLMPKYKPx70Dh
G0jcz7jPOmG4vcxUXvhR5TCBheIxIJfLg9BQi0VMvvBomVJrU6eHsr1Mr+UwMFqX
sixl8DUR7oYB0aM1IiB5NdofwLBpBKCnqvFwlcqa3ZxrBdoCysDL0mUk4VsdOP5l
ChREspKDbHx/0MV+CTCed9lelTz20QDGUeZ2U7uW53yFiNJuOXD9QrZOABL3YMcl
3+huoylmg/kI7e3C2myw5VoR8XfxOmIj4DIHLvHFX1EhqJWFy/5XBsDzRwZg3K0S
KoPcqCtdVQGSFsyj0QGH2E8BUlZCxD2gin+KCOSK79KckFKf8dkpOjCr3hA9j3aV
tsBhgL3WIMzRCds3DovVnjVqi+S+xb47adillceR7UyiTJtvP71G7GXG0pPAG1TJ
MdcblFo8ERr7r1nPUNe7O2yZKyfKJFSZgdw0tH6RUdp3lXeH7voM/A+dk1DOzkFy
OnYKWjV/z6+fpwI6JPmsJVZY49B3dohV6KwNx3EcRt9tZNRvasSNwcZYjJFYW6HR
L9bZCfdrTGxLymlj7g4ADvV3SOmv0IB7kzchWtGODW3Kny+Pjm6lr6qm9HwdxVCV
Mb1PuMPKm7XfQOHaoO9KDHm773lRGwSSj7QqHEkIR4TyOSxq5pm1/yUGUvmS226v
rZrjb3Hcuzao1OxkKVimv8CkcQbFcJw8EZIcqEBPcdC+vflVWbXuEy6+TCvYEwGt
kQ9HqSVKb2bBIJ0EV35XIZ246Lv50CNUEpbohSNaIRzvY/teFtyDe6Frc6N7EK6Q
AI63UrtgXCSwpeKPUTc0hgwMDtNdWNIwSC6JPE1YY1fb8YlH4Zac7llF1L6WvXg+
vamNk/bAQXqG2x6slkQd31/KVTKyxxdCoh5bFzH/Qdl+aow+88yIhQKaOwpFmZYv
0vO+D+/g2iszzEza2AJVZco63a9f+/lK3nVwFRtxQp4Qhvvf7YRtJsGlaIhXE2tL
rJB8103PDIQKcBuO/b2PnocFx4ptCXicYBxEuWq54c7Q+GveEkgBgs3qaJFeLG8C
DDnH26yUFw4BzgNlcRxiQ+QLR2clGFzZP7RYe+MAndoZoum/cceec4aKMxzSQuIg
r4ZTEUGEyNXKfGOvhAmLLItUBDzl40vLhIPcLN3PujQ6FbsBsMlcPD11Lg6puYSI
etHRbFCvt5R3xfWZc1LNEtqKeLW+nKIMWEdGctCAkOBQXfPQFcXCfa45NurERh4R
44MAfhhaq5XkUucI7b2dodQbF963o9JlP8bRwLXFb1fShm5uqwq3BSEtR7WpgMqf
QxCx0SfZRd4cJq26yZcaeA3Z9ZWUemBqeWR50pE1bzbd/z0gF/aw6nbpcLd/Mm4W
s+D1XTiOf6NpXOnC0PN1L7srsicOm+tv2mPHYyxjLkKumAi7BSI54pPzoLTUfioY
cEM0cmeLAmAq7LdJPtQCA23MfM4VQT6F4dRNeU599WcqiRMZFzVwhcoHoZ7FPIH1
ZcshZ/lchenOnoipSjONtSWXzRsWgAPtvwyTO6ZgkmsaR2Fq4Pn4n21mKYtajua/
Tsqu95IugizgmG658GhEEX4BguB2//EDrGyb7Ja1SxCt064Du49OxxE6ASAFnK1K
oG/BF1byWytlNQb5Jdz4F+Tu2GjqK6A716aXdsNU7Q5ODbZqs49cbLRUprLmAG12
vmKquM97zcSJasgP4WDvOJSgv0Mu+I/3VGFNXJsSXys0slm3Y7L4uTLJP9imYCjt
SB+bd1LgRpHvtWJeZTbXakf8EL7y81gakPIchddztwoeJQQTr99Q31UVE3CNhneQ
iA/px1fnVv+d6t0AbR64/n0s5yFGGA4lHxp7/H3zXTR2kgqFDwgGomBaRw9ua7VJ
tIPMWEIVWBE40l4CUNJ5SSAK4RLiRPeeS9VloyVNKzr1j1cd6swCDBoU0Mum0lE0
27G5eMEfJMJX/IHkBvJ9y8CNcj4L/fVKL9gWHKXI8mD1aYGLY5Vj6yVbpVxlqB78
ra3Ra2VlFXYtWxQF/rpb+t9yJrUYPFvVN4y2zaxEB4ImscRAQRoloCDnHSyThOhE
5azAVBywjanPyrguu7bvItWQv67Bu5RI+89csPCiW3G/v/NHDZAE2FC7h+QOBc9y
Bnsu12LTDCEnvOOk6pDNeuX0IQzUckWje310MOCA0bhOiN+8SpDY551ulBpbqih+
orjhBya6yqn2mx3OgFsV5ruWSUYullz1xzDKGpU6lnn1j22vkw5f59XFFcDU6A11
w8fTtGZcvzPtrA67JoRl1i6q3m/W83MVUB4gMpatWLNm0y9a1PIHaXA3nuQAx7Vg
n3EkndX2uAV2FnGV9hKJORVcqiPCE+MHrdzMIispko5qvqrz+bCxfHKK4jfga6q+
WogHmDTCJ/sRb9kv9bRE6MFabQXJK85HJWGdw3mXe95RRkFFWSRB3xVX1jCyVtT9
3+SrADp4MWs22H3EBNGca/OJc7CrAcxevdFpGgVHqcCK9Z9e61VWdc/oNwQgGFAv
1mbrg1/rj9aBBe+pzgnzoEo4CCwhwwvf0kC7FWj5ySfLPlAoFO5uy29Zg1C4sapH
P08OxpZZnYPXdiup5iNAQtPO/fNLWHme+5g6lk+fUy/IyCaIbashm9gNbPg/kKKT
glQJyvARyndwuPkGNDzQUWC+bgYuH2/9a7+ExOOFsPRgy5r/5sJX29QF1wdHZ1XM
rLHjz3GKeF/3aOA5v5cNlbqaSYGnowz+elm+1/mgxyHIGT9YAHFayDFyZ+4zKI9E
YmSsATMTlvgns4VXQgn0puYEJEOxdA55XxuqsrvTTstOYqwA/TYHzc2J5As1psfg
TIcvSPKzt2gBw5w6cT0DNwVlPu/8IurwNjhmaq7TrmCAQBg6vXz6VdAFq6S+1OSF
AvRS/yV9jgjTQN7sxYSeGQoizbGI5Ei45xhxe5MIQtjibEceghcKUxSYj5mMth7x
uZ5RUfFHMR+QfG2vqle7jh5sz08DK8EICvC/1VndrbzMESSzcr2DR7w7+tCfScL5
zXJhrnRLTQEQkUDoZFQyF5jUVxzw2XAyp1lbPqOLU+xIL0k8Tqb9Kcfqs4akxlD3
yYWSVyTCzV7gvnSrbD+UoAFxIHNFLH9Y1O+epkDnp/cv8fa16CkBbuSqlGHWc7rT
N9Iwl8dTgaozUQCg75mNIAJd3f6W0FziQMuZsz3ewU4AaXuCwhrcb91qBFv3ZGiY
2uwFOIXrA/pXdFMpXYHrql+G185BaH/yzuoXbtWLdR1PMZh1DgTOktKgYTX4biQg
LpSuKophi1+kkLh/ZNvknZ/km9V0eB/fPEpuYCw/zUD9X6faDiHL+gcbREqmGZaM
SnavrwPGRSecJOPdjb/uSrdRu9CuBLo7uZ1x+byFkpFMxtZSATJHqCPu4Yte8wXt
XSj2ruwNep50m7q2wJQeZaSRoPOow/6P2nqFrMugUzjV4FR89HCopCCyN70aLQgB
z3FKvFSfMkxgGwmmAB5foovbScihVU+N/Oa/ujNIidCPOCPW15lgfato+oNOT9p+
CbAWXaX4f372Hy6nnurl68w7pITyCXHUBYONU/HWxcMWuZnKwmIRNeCk8p0SiMZd
fqcmUWRgeC7fvvgXyH8RPmJQw5r/svh7Yn0sjdoVMRjhPwIft/EDkwcJnKY7j9tO
wSpLziVYMO7d1xvCL/ERIukf3e+Iycg9UMaVEiQFWZFAk3loM2iSQx4Xlkzwg3wQ
KWnX6Auo/X8V+og+h7PjsOTSUgs80LV8nrcnXVwipDuUm3QJ5k3U88gvvTpcLoYF
3LSRPybSM2YdmN3rJWmUasHC2G+Lm+x9LnvKuubAvG0W8eKW6D/HxvYvHgueIRDu
fS3s7iPU6fedrNTd0y8C1sKSJRIIF8KGUKzYNAbOjdTEvFqCR0ROBKxo3ZqPxToT
rpk/neA92/C40r8BTCVNShiynDk25KDNXC+CC3gVFK3vkPqhtEWKeM3eTcD+B08s
i1ry4wuW1Ghx7CPmw/v1gEvjyNrdA3FtblWqfo5RMrCokL8fwgd3BS2p7gvEoxI8
NlssIDYyJaXqeOCH5ZdYpPRHLje8zEdwJ2H6NYmsSJpGFlQWOClfMCDQQKcRuq0g
GwvRAiL3yWSW7a7Z4q4m7/cSE6UWZD+SzeFAXwRKU4cO86InvA7M3PLwNoDENseN
MPVIRPzDGHWOP7VyYdkOXrXshWOMS1Onp+NEuBWDf6VJYpLnZQKbU7r8VKs/6PNJ
cJ5nRxhv67dAcTrMi7RGdVarpYekWjwMYrdB7jZq+aUL8NkGUquJF7j/EdxTn9vp
6+5je4K9d4TL4maXzj8NfyqKhfk0QWua60vsCEJGpZHkUF1nL+KljGFsTqRIsP/0
TFh/osaUiEE1b63tDIc237qNRdE8RruKOQeWYseQKN7b/Lt9V/1aSTCukCAeN97R
hhoxLiaiPBdL+VcnUsoUUhtohyM3YzmUxx4d/kE90dshX8upr0BarjExVG1D8XB1
Do6Gm44QeP8hKBnRQHNAQqpT6bB1JYtaGu6VkyUgHOP86NeK7OzhwLqLTt3yh95r
wb7k2gvPZJ65HjUsa5WXTT9ZLeplybQJO0jQMeqmIfSZS3DrV9BxoE1jZYwgaoiV
wUQplHg5/aZbOOOxvqpIl1Sh/pzm87S1kwnnC/Lvy9fngUXUp6cZmhkuJ68xPCuw
OjRziJQOSoB4wvULdVJ6ADvoJdTb0cxPJbjDklqn9zWFo/a4GAiSdUh9y0BZQ8aF
rUGu2/kt2SAkIj7AP9Ols+tgS91tOT6rpxq3R2AaQBAq4ubC/XLvPuHE2ZtugTJD
RUZLf6FtbG+Frt3AH0KXhw9hM/j00qE++tqG1h81zfuH2HAVO9EiaGXZnAMquM0q
7MJvEP+99+7KEM/Nqw92Q+cpieqgR8e5vkIpiOgCvOEWRNGZi/J2PUS/c/Y1xe4y
Eq4vonn1XZ3nnscbhovSyb2ZpbqXw91Som6yzjkLaEDpBsC/g3DBYColek5yRgnU
FQlHGHaw2u+JrICToDMqUMmARXhNsKL/j4l+UE9PRgsMCx8eWqD3ONJ1PB6DAppO
0Q6eRwiAxhm7bm8vVnD3N/eCYBbTL+wjll2c2kgzpjNwhVwsViskFjf54ryVlX0B
8+J2td/D+U4mKVfA+MFczI1s/4GsLhu6rDmWQK+fB8nvBj29gqNhxujkQzEQ+4ae
F5fRa2w6feCsTBrzMbpCbgsoUe9cZO/X/v7xaIjPqZHK81dXMP9To3kPSfFE+JXE
aFTTE5KvJqfQ5XNmljk4U7QfeSJxbbRA9NqwcMI3ie8ZKH8Yy4NunzE2xeBouf3O
uc9Ni1z91ZjNjKL+R146wLdOY+m7YY4G+i8dgIHpZeSGnQNqZMUvYJ8ubdgAJJcb
zNkpLImcUtp02RnR65/QCt1raxqkZh7T7Rz30W5i7BTqjrAsuPrRbDuwBlDFI6EJ
FFSO3jdGmDBy+Lj0816BJuqQ3l/dP/gyciwWGdRgrsz6KtxQSgoJC9YdN0w8Z+nJ
fBduf2gvqNCBXeCixD3ePcOj/fvJFNHvtrC9BFi/wgsViClu7Zd8PZ6TtORvGO2E
zxtGIeKfXITtoAyno6DMx4V9aaW/Dkf6wBNSiG9nJkp+GcGRcNvH6QPQTKaNcnxG
9ydIdwdMn1/SqEVFS+KTkHFKT3JtmglZEZE+0WWk3kTh2pcRQbmtrZDV2RXcMsaL
X1ghrTigtiT4mE06YWPDVNWiKHqUh3iFwL2d0Ft5WjOxt/qENHhBOcMruMrb3pHW
eDMt4D7edVy/Lq2+s4zSWRZYgILNG1QsjbbHXtUHvraQrbwrkEY6mPHiZ3LOUE+E
IUXqUk4QIajeuvYYB+OcpaombUzzbQUyiQYWlpZQRuWNYjFIn81bUrJvrex9BOkz
v5W5XaJDI19DEnjwuwoXQfkvg9FHGDHFdQDZJ2izaTCOZPPKIXwStJKe11m/vYjc
ze2WWEFhIe9QS1fjax5AxzFtJ/6wY2xvV6dg2s0+OipLEv2hzQiYGNZ9a0NCQRm4
SY1i4fDKUVxmOkfYMQJGStOQWDGEBtRVebqPOXy7DpR7jkEhkzYzE26Ap2B1tCdj
BvtiXJssvH2i/4PuUlli5HdMECRsPYcsCd60gEido3/+UJDBfM6EqFqz1ufBqWz/
OSBfKRvq9vwiPs2sfBvKvdR2/uJWDKD5XnljsgeazRrrImRreN1WQUzzzfIKIB1v
e2rcjp8bTS0UtiBCZI8cw1Yvx3UJBBNKOc/UhOFzSg503MorEFmOENg0iN5tI000
ZC6zEfkk1B4oTrp60Pc8Vpkevif8UswMWnVrJNsfQ62Ojz7kre3KBaxD+Limsd7y
Q9RAQo+Teombhjag6kZjlidl7Vu/CW5tvqFidtbYw70Ho7rVlSieU8hX7Ie6fmnS
I6m0iEwVygpjnAbmww5XKa7KDx03KkbdDGVnmnOkKAsVu24gRicrmoN1U1/W3ZKZ
HZ/lj5bAww2Ha+0Hag5L+EEN/9JlqWgonXFwnthruYtP2We4lyQxwSPypVmOE4D/
sYtAsrl3SnkA2nzJZqOkfIIU4uV3KmYrFSMRrSg7DMqANewFrEqkZzXxIBRKvd32
ebFML5/SCCkrlkHyikWI8Xl25KMVTe36IJuWOr9Frr0WnEREBX4yYLY7TZoQAMlU
7TalyR+UF5jJ0Z4y+biVbF3uHSqWqAPVcl2kGImKiZyoQWp7kj9RLABKHtCsZIFj
YqYgcP2SdQ06weqkyxCKPPFw97oYxpIhPffyTEOmolrjYYWFYsJujILf9DDBIhbn
71X3DNhieHAUkza5w2G18rwGtFMh/FhhBRVEpeLsCoTRqsN1q500vJH2YjYFTUhT
5Fk15FDv2rPVhQEoL4ppkhn9UO76Z7P4aaGUcmO4qsz6UdBsq/+sJ5h2X+wl9QP5
KAsYygs1r4lZVLF1BfOxLX9rL8ZHpdbUeoFLCQxhKMRKX1cAzUIM+U+VwYEUtRyR
9DU5o84ml+XrhLYfU4Xy4jMWiZyhj+QJWdFraOnSJh4PG1YsuByMimbQKgrakF3u
A9/fBegVdkD6QRN0XjHUiK0+YLlIOZawKKR5BJz1ooHun7NbIuPsHY2OhIixlFYV
HGQxTAD+/TuTBxMUw/WXVZnCcNkc5UEarTq3mFo7KuRKHXD/I3pmcj85YG2JseX9
Bji4TMX4zdVwaviE3KnEQs9Xf5mJ6RidN46cI10PsA5KuOUhTCbFCYLjQ6/85i2W
t3MHBLZH1iH1NhuACzKUsh5ObexjV+UVKPqDmF13E/00ROWYfNwiKluBWek7BrpY
lhw2HcE0pEqVJ162BzN2blI5Q6wcPILFiul771mwegQkvZqEU4BU3SskQyrNlRyB
/7ZjdDG8FTJAxCvJ5OH3DGN6OhXkr3/Iat5Q4WM0Q/PyDh8e9IrtqFEd/Ncktrgm
EKK5NzrnB4+fi6w58UrJ6EpOIidUzClaVy/zQSYtypLN7xH/ManFGeCgcKtpM7C5
RgfpfZAprXdnzGGH40NbVbyhnChNX9rBYijYIcWixiLH+aSSXKT8tRvVyE/E0Yw0
cBVqm+iSaM2xQ3Jt1mqWer5yIwFy2dI2Y5tBMvuuWgl8xLVBk2DEWggF2/oOxaPs
WGkvx9Zvzr72VTNul7WKEqW+yraJ5Rtt3haIcQfMyV/2o0+FqebVARQD0ciBsoKu
1MYa7SUSn5MlRxx5BnctElpOegFRFkcVriPC6vN/HKVfFUVvejBg43peOvK2meu6
SG+LUAISmDjMEs5P8P0+8fp6xaU7ftZ8GL9+gsfkWvjaOF14v97XZ3DjBhpF6cC/
EbrOLmSUAH73pI5Xe7QQkthodaYL1xAU2X1y1g8PYfKH68d/Dtcz/o1mXOZyLcQb
rmKl3ygw6Fcu7RDETVMgAqBULMZ2e59KStTShCg6ODcS/soQb4ldQyWOo9th2CbR
utScnhflyTX8ZKYB/0y8T6ECAH82mnMOS/nfMnK4EGgJGlbeWXP3ZbVIF3UvWaEU
Sm/B+bQFf0+J+8nz8tUb6e2ZOvqawVbobDSYko9vyoAxo4KrT1XLFwSyoHvOwtQS
gAfieyt/B0Wfm18vDlbVCEfT96+Bp+/PoLPla3aSMgsEHsMx/yEopWDCvlrpRmO2
5vGlC8QLWrMNdDkNm1mb83Zrt5oIMlhnloUzW5BiCtVm+4UsygTNHGYmQxu+TODo
6MLEPkfo1uyphBrTE/XMrHcpIIaUqyp4K3uEBokeHbW7SiNWo5l/Yv1l+0973LCV
ZP0s9Z9QuKeITxXBJindn2NQrGPa8SIjFU9y4CZTJhrqS/+8HDArGMwyWPHhvczT
mJHs7zMMY1JN7J+hVV7ivKyYFSp7O9yTvISGZAUtuJ0alXLRPAZcaR3xB2b6BMFZ
GyrDU/8uSb2LSmZafJEKtmhlGy4ZL1SoXFpityh0t/pnpCRNaVpQY4qjGYLfjTpT
exnNylyLQU9gzsqGjS18qwRjdyqGeUyNkX2ylaTzg6h3cPa+q1LxMg9WxqC743f3
DjHrgm3oxZhiUIVIbmCRyhyHws/O4vXSvYBkRShB76gea3CgtA4YpJ7V2khRUkH/
kC/TnlbxdO/RukbYGM1RyRwEw0QNC0lO5fHz2Kvbaa8/SpylRcmZHfy6IikpOvr0
rXOuv5vongdDLbxhbjW6jkPvCylXAioGQFDCfsyIR38oGHoQ7HFeRIRRpwHwVWNf
kvIzGBL+2Er28bE40oCx7luulcBvjT541v+/WNaFspid7ff1FmTXcIHki5QN6hBy
4W/Q+Z0oM7UQMgfHbCgu2/xgpkTIhpQ/FurN2aZ4le1Pu5a/Gd1VAiBYo9+Ks1IA
vNuCAYA927XUqgdimIj2A3WNI1vmSRexQLxTWdwBrcSyxk8hVeMCfs/a3P9mKJNp
B15+pLROfss98nKXk7k4nDRH0YX/PRTvyKaI9q3vCdgF8f6eKfJ9ZKD5cl8l3c6i
wnB0UKt8cvgMA9K0igblRYoKry9tA11gJeNof8Zv3ZIu8WxfhCmcOyrAJOTaEBKL
bT/M+FDOiPu83zrXRlJ4ZVpL86bG7lMQDvG6Ubg2OYJhYvtaBWlHJp8oP8PDxYFf
cYtsFPSomZCZdSBXhcsaHX42SOJ7B6Vj1Wa95pzEybVDOIZ2KEibq/Hk/FvAHTyo
f85tIKXh8djXZkLBcrBCVVwIGhU/XbtAwVpq0mwMVTc1fjT7Pj889TUexsvseZg8
7G1f79fUyPTAIhS9zVp3rpjCbwzV+X7qJ9Gd62drpmYBrRBXH4oYckw1JxIyWCMz
P/knL2poXiK8ZhPGaLgmWVtRkDdSEI/2x3NMUyyiEWEgxpq1gdtRz0/sAMUTM3xv
rTBd98D4jK8Jz0195aavht9ofnvAzF6c2qo1+gntWsjyeNnfRyr2Mu8+oBctGScE
DxOHiNMJu1Na3p6Sv1wJkU2/T+3fBUexiEv4fO0VjjN1o9dY9lpkHp0wbR9HWoO3
ZQArw6lphzys3Y6N/gZw6KTQA71F0uIvbuqkQnElOCYakKaTVk0fsYNdO91CVPpW
coFLpOf2+XvOP2T/oPX7BV7Td+CWysefElgYcENsnzH1Mc0MlAplLumfgo7ndLHU
gW+/p76QGSBKn4oy4OkJD3jPzVjH7OtL3vg83/9oBoix25evhwqg/fDgn39vBjwx
P3I0gVB1YGcq3OBXF6nxXl54Dvn5c1pgfJCKFCdLxoCfLUpQ+WiN1SH2PCA7YM9O
6DuQSUdr02egeryZHJV0eG7aIdJNsUqg47YyOQVEb0f4MkSadepO+iyQYmYE9iA+
nyb2IXlYCEXiByYvKrBCUR2J2OyuUlxAckoreexJrYDBGvbBHwkyHxEzcs/nefe9
iHS9lfAvsjgiiHQ1JsXRwDlsVKLRp98L39XTtm8kRG9DUb3nbxKb3yA+OY/kADXv
YaDZXHOWlsI5Mm3sR4ppi9NTE9/POXm4Gpado7i5b+KAWmynjiOsM/y+PHX432i8
0LAYJM86mzhaUFtQ0rSEdEjC8X7rfTKGSw730sEakDEAsJ9VAVkyTKhiBdKlLzT1
j+26lGUv646RAW2KmCCjQSweMPS4exNybvZYiTfwTD4lIt6v2L+GZSQipck1oYih
wDYlhuNhXwURqqFjf026ao3VVpd2z61SsprteOV+SFLBdC/bRk7ClnxLiFvgAqai
+BIPfDWHkU+D6e76FpTLN0vahyTVAZIwjijpkJFsK1bToC1XjwLXSC7uKS6SxJ9Y
jrkz9OEunbK+pYbwwLpns2rBRIsBQW5fUn6qVgqJKJxKEPHP3IKCMSaMwcowT21z
cTlmVgzvoYBbcNyds2WauWUwGZpTxHsx3zXWXdWNHFIqQTS0U/fgjzqY+slmq11p
ajlxqoEHvOtieFd35AIJ2mJppf7ZaYg0H3YFn0pnPrdehxtlN6E+f50bIxqORAne
UKeUx9+sp3bsAJuuvWADr7uvN5bxLF0fHMwmz5qkFn1yFyqh0g4SPecfUyuk75rn
UUXPZBcPz4vJoN9rVysGkw+hMKY4dN00G0hhA1LZF9rbWeqNZLeV8L8n/VjNLbbQ
SsoDCwimVpKN+L762VhFRkfznyUagckbZOi1Aas+aeoakkbrm09D8MDE/8ZBKEaI
7jxShWRjtV5KFWtn1tNAvBo1H/FWMKpfz8+PV5Y/GSR8IURAGOmJ2zfrXZktRTea
0wUGzjwlRUjh37RMAySRdxNkaksJw7pM7kDc2K7IZnc8q4oWxKaDeLm52GawDrWx
aHVAih9FLgPEyO1/9SBuo13yoGsFQAaZpqlSgzWIU0wurKDRHdtm4AZDMRKgv4JB
Ep9Jzkp3246SkhQFmYNeyx10upzXh7N0D1xmBKQYuAegzatPIXira1+LoyQy6ePb
1nh/xxW3yKHM49EEy4xLCbT8CFcOGjQz8xFN7MqfL2BgLslK6iImx1rkAPss2eOh
WyX6yJQ2FRrjskr3ZRSefk2QlOOiQ9ecI0EhCZcw5iuF8nPl46rGTT9Kuac4yp1Y
gb113LqEIstftFRjmaBCr7MNQw5DpqvJUK/CILvVYpujdQOWdELDakdDnnrUUM99
JQIVy0ilyObaAcYwLMJEpBj83RhskExgpqqMnuGCULXHsPXXd3FauVdKjXiY0Okf
AaIWIocVpxSjlo3krUrqMHDWqk+4noOxXjR/xiZdgt38GonNCDVoCKQy+yuVwR0a
um+H6p+uPZnj1leJNwLHfdZklXnY0GXpMfQ9wyE46E/qMECU9CSpEExTVO/zJ1pN
PFu/qyDBHJ+vOqsyijs/qONPUlpXRDff+02elf8fYIHU5dqa6a4Q3KR2/HVkI8AP
e8DFWR9nZ+OxOMbd1YEGV06YDi1Qk6kG9nWGvdye9Vhieou1yxO6kCva9iXL+Ngl
roQMeTHQG+++2AFsFxbEs/7FxWYsKZsTnhwy0fclVat366FOjO4FCHDYCG0uY1e6
ImguYE7qgpKcRc8N4QyTfSRmzgZ3/ro2OZHnEolYRJPJSp0QEwGxz5HH4z6qFI3I
Ds7i7RrHhCNj9YrX5XU6asb0JUB9OuH5ItREqJhF++zQv2yHxP6gXMbuTAxfmvZ0
rB6xN22C8aEmx6ujVkn9p5WwlCrnij+29sco4yum1K7yR70ltW8v43PMM15fFH/U
+4iOF6vyW9jt+MlVme+BJsC2EpPD+t+iZXDKIqWeHWQqNxyPIce3h1X0OqciLpve
RMbqZyetALP7MJQNz/qiLjP1JU/qx8e8JYajNIEshzHSmtjxVsMNt2IMLd7RdUyL
nCR0VkL8C//jLJ+pOXtvGgqULZ2qe6o5yWKYE/nxJyiB3Nmp1BKwcTsoBD4aeNOp
YG3T/OwyjzUan2LpRlPEniNnkPNE80hlhXWRuCS8RV2UHAxoz1uz3oOFbhERIQMM
LHnTkDkiHZjTa1swCgHUsunmCAE6paiu0AvgvGdHnY00YsvWpbeytoK3ObldMcYJ
mPPCxt8g8ZTrFpZUtMJWbaufJqsc6QHJL8YWFC110ZnkEtSoeGI9sPOOVaXp3joT
Xi9HMKe1iPcaAI1uC57lbLhVVspPvDCLHxVzyp09E37NxSvHNfNJseuPrpci1wFE
05gVQO0BoJMRLb8dViQNIBmAQICDRKP0pZdg06z4Jov/6H/Je9yy6YNxiECzz0Y/
zqhuTYF6OLX6MpaA6uZSZxYmEShKkl8ZpC6oHtR+2URxmpPRUbAEydpGYz6hkyru
dofnSrutMIALgkk5uV+9Yp0eKuYO4ofLT9V/AJylPlNgIZBhm4+CMOxLl4EXI9Z2
EBhnZ/5ERtsNP8hgbWo5UcEfcmYt6uLD0q5Nzv1PWgydvHcsLGRYr5tSGyTbaEsX
F9fI0aOfX4L1QUDbBEjoaUu7Qk3y0uE1lPKDfwy4nuqdNPaVBw8T85mqkdXp9E2A
GGIYUGL91PYm3XSzAv4zlC+Db3xueob70rhxcaF/k/Q+oPaf4fL1BPL2Fz+u58Zo
Nufylqp3HDgQpBYR+8JoYWPbE8pDvUuyD/iZSBOwcq1V/2uPl4q+ZQi/rWcrieKm
7CgVnSHryQQ6RaRbO/8W36Mn1Gt2KpoN9Hv+X42osvHx2trLZf2x9T2mmZZ9UdQe
2nT3ToW5sLzv2nlYZbgtDYfFWwczszKIrYeoZBDE7GZJ2G83zmRIH8plnt9W0JaZ
fUi9uuM8c2bjfa0v8GIGjXKo3gRx/LknbtPI5cxL8HiUwLGp7gg1FX+WDt46ASf8
wf5uVAAoSNw0ano19L5ncd5eZsUGlfvNPiSZ3iHNhCfXu3KZrhQdA6SNwKOH7aOr
/ij8pLtZ8CbVYc8n0+I2kMcNdCKmGeHC36sgfbJif1g0hQClXkaWELE+AUtydPKs
tDVPrI3Z/AoAwfPxtMdCgtDrV05iawobxJIarDkvcxLKtQKcTqKdt9xl7FE2njoS
LuaV25rhXGg6YEbuft8hyLW8WbM97WaWkhODeZmVQr2xyW9s0V9xoKHECUV+51WD
nHEX0I43zVac+2iY4CNW7d0hIeXE7FPOkskINVMiyOI0rwsL+Q3/ubvEOMHZnWLX
Fn4ApogMcFn1k4jRXXR0WFTPX1OouQgy1UOWpNCQryISz9HHDVBZP5HyPHDC0G/I
WKqX9RNAmHy8Pt0Lqbd23Ou0BQ7s6j7QH/n/Jvvn0U/SV903EfGQXfP4Jmew2bAq
ZF0EBWbTLMreVej5eCckwuz/nki7JMTfUbq+rZE0M3DcUaUxgrM+x+qZ92LA3YNe
lq6wr6QQ3ZSUz/9LYCthltUujx8FBr87CglucIwVPAN4xYfhVXXNWpkzXOzaGM5e
q2+9hIFMLifTtryqYdXhNCDFs/PLU7y5SzhbaQ3qArfi6zRVXJI3VU9BCkcLlwe5
Zu7bgjzIOMiW9bjWXwi4uQwTkQiujpKjXx9z4Qdma3BtXVXqdW8Fd9/8PaEvNmYH
y3+4/PVCerD7qzjrNpzqKhvunkWWZkcHTMUh0Y+cfxE/RkOdqm6u2zy9s7/4u6VY
l4q/vZ96EscGku/Bmb/eFYQvAz8uA/mICi1QUkJeBTJTUxMfC+S04FBPGmA1C9tj
ZvxK/Tx2WpXxC3ZMf7Ken8C4eVV5h6LygaqoVqF5GvV3vLuIn5JsnUU+Y2frfOSh
eZJO9Cf1uuRKbDwRNuRmeA/3pnVXTTRG27PPjiC1M/cPI2ye6y4AO9HkmV2hQA6J
Wpw+Z/7iM3LdDNSRqrXTqgx02KBsQLjsn+Vz0UcDlWRzATmHG7BKQcll+b9USXrk
6f+Nbf9nQshjmjdYZy8IM02PVDV3sNVFRRbE1VVk3NKz46Oev2KYlTejTqfzlxgo
Yw+BBk9JRMYf6ebD1VEUQQYrzRGOk0SltkMpL6f0e+rvwCmp2xJqp5lnqR+AV7M0
TFeDfV956yY9SkFYRjKMPMCkKsj4eoul5kKasQp3XTZMJLihmXUtP49A00xvxaTp
k+PuXkcSXTfXQQC5ZaEiPo7VdsK+Ejk/yfzI5cBdv6vvCWB5HKujWgt27nc0kRMG
dHkiq4hr3aBmrBuxXcQza7CpQoHsE7KL25aMow2S2W3AKlNHredJitRfs28Sr1On
Pt9qX6Xaz3vJqOlsirB2taLH+3dAwOWgE9gfCLqJF6auDY6JIfmre0LAT0Vn6KW5
VzAcBdf/2Iu1iI5tv/9nseWiY2UITibxuw9HuXiHjeaHPxxJwocpYylzU9xYAi/+
Bt7qqJ9RBmgc4cSCBzxaAlHicinfzLJCTMHWN3rCfTo/LKf8ZAttyGYyM1GPCmOc
51BxEWYZ3ptkewrKzUChe6q6p1L3QcF5D7UkieFhpSa9fH2onWucwaTOpJn+SWZA
bVHG5TUTk+D+w2gXIrtSU7QEwzDPCTVZPe8jNd4rNG8VczY1Cfo/MKc73/7v5+pP
/vrdXnpWF6OAI/43bH4IrWMWiSLHi9RxC3gbxNkhIFEG7L6V6liqzvFWOzofUrtm
YCCpE3Wc+HITfkHkqe5pTG38jj6raHuYB32fLUD80min3R/kSY4gAvCry7RbixVk
izfpiT7o6WZwuv2e8qfDPl+XvW5yesesdIoL+GY7qC6QVyGusNblJr56WsO2LO8u
cP5idAnEH2SXVD78Cnh/gStVkizghMVIqMbl7pmugN/kwfqw0RMPBHAW08jJW+3k
kdWvpDmzHNKFSa8bqgxqytouY3b8hw+2TmdVDv9MiHpZRYCtZL3cUbFACHh3YpjW
93AoSJdLFvB4t25m1comWuEzWJGjG7AlL2ku0vxyOtaW04im+5dGucTM1sF+oqyb
CdrLt3TCYN9k9Ih51/bSwJphUKhNPwyyu6J0F+G0n6abWjsSap2Vo09I02uzbk41
b4rpyQqcz+4/34nT1U0N9RIJX+0abm/6VNWjjuNCDdMjCsx5mr8Y4KlPQKUvhGBe
mleYCZULgodGYJzSAKyTKX8TH93g7fm2q5/yn+T/II8JkAdr78aJECzCU58qK9b7
R95MRVaIuBzbnM/HyCGM+6re/g+xnq86v1yYRR1BI2zFZubQ0JQOQrkk3ApVJVlr
cDQPw8cGWfk21J87miGP+26WymdgrLozWCnSQF93awNH6MzI48q3zWZjkNQyAGZr
OXMXf5aSYpWX2IZjz37KaEHdjcSER0mBJ/N6TVZFrhorelZA5xW0Tlo5P09Ia+Om
VV4TNvZK+UZrjdLtf7LtrpoTDtfYreW+XUJ1HhIRfCTu0phCq0U0hNDEFRxqXfK4
MElHqjpEfaaEcDwIXYKZft110UMZfClBnBijXmhX0ME4TspYKd2zS7ZOs6jRCHCQ
RkK38BFzblwl5ROG+OsNE2cOFJDPhrYw/ZmzScfZrHZem17GhO+2cG0QcW01DXJ/
ucpZvXN37/RwQ1PauI6P4tOTFqFQ5bC+62phvcXqb0lLd9PKQswZXl5sNvixOpw7
N7W119MBbHCUdpPcmtA84zisEW1OlyngCmF/EVefLs3yB2IKJiHvPZk5Pzw4ONiF
t/XlhYdx8TVOSHnoNp6wRqftk0A/QT0CSfKsblA0DbYFX+DH6NWxAbP8euyIhjKM
XHjQtufy2wocOJ+fEStt1cVEHZn8tMiAe4jTGncHJFstbBqBTikqF3meYHxVBBvW
sPXbziJuHOmRpTpcR/0NYcpNzPFzv/dPnwcLeqhxghUIU5rzSPzDCLtbrgjl/qDB
4BW9k5GBQfsHutLKzCvpHOfUGY58MdzUfYza56xvHOOyhQet1VBwxMvuljqW4/di
UmQAvU9tDyFRSRJqG13leJlhf8wgyEQtb4ooGgX+AZ4mUkMLrPNIvrIyi2EHLyeO
7c7FntiUUk4dxfymW0wNixZVf8jMbKurSFmovn1IobHCPkQAOU4hupPpcJ6/nnfY
BbJ8QvaZzpc6oxMPRdjCc0F3rArfJhArXKbGooQhoOKvTzToZVEUyHMsgwkTZSTu
7sWo1RLE08tAEgJ5EiszgbjsNmmpgXNxmO8Em0CsnV0BxSiTC2Hit1PhP//450Lb
m+D98KNPie5vHN893M3ikta/QggbfLkHMAazZi8gDJxBJ2RgPzMsWu3WpKDF6fcy
KIVnGiUqH6gsGa/lJYnlpuGfgpXD+bHc/+kA0QND1YVZyI1DIq3yQcDcbmYclVfL
ilXF+IIVxSsBq+g5iBxaYXdWhYlkxNyo+Uh4uesvdVGARaW2Q6gIVXZkEZvDutns
DgtsAj5qwTon/ownZp3cMuE4tN7OXQPSk+DFm0alUVoV+3cXRDgxy8oZcO/TSvCS
YQ6VsCX17jgbtPPwG3xlv7cWW3vcDE1R6QAYwy3cHj51Nu3lI23hUwJOmpbJb/6h
pfkNkYFVYR3YYBhgfWjjR4VKQEivGmoYcIRK2LxtTonR7enw5GbIEygLd6LdBBf3
fF3P081pin+bNqt3USVlCqxwLjSNlWNV6Ht9nxuVt2RK19kg+Nf65O+ADX0k9NwU
iS49y7dn72yBN8F7wF/kwrSFVgT4SkzO/Lm8RQkfS3IUbrRxbT4acJqaV5rTVhc7
GnolydYB+O0WRVLJhxvPmfiRtuJMzHmT5lb4nmFZ7hvx73D8Vg3Zd0FoGmGzzLh3
GBHT0QjiFeluVE5z/4ww6ma2xpGbrgPcG7IFk1o0N8FudBz3lf4od2BlcEmze7lb
vpXkvuGEjm06hPuuodrCZ5rrnHiq2kyI4KC5Jo55at61tUbe8qIKyU2/pwTFWKDV
j99e9qL9XYRAIfJMsZ7WZJr0RHWsAcCruwlE3vNb4MZ9REyGzV9/qLYYya7WtrZz
i79xKqKVYYORX+NaXSaeQmPZjFiWuQXL1NdRDC/DpN/yPSfQEgF941XnbnBH8WDr
q9EtyGmD/1wrSMVvN6AerH/f5LAc9eeK/mqPE+S5sJmduW6o3if0bjSnRxPyWi/5
6YKGfatgrysxVpYzF7uX4aUBxmz+n3KUmKSeTiEFOekJJ9sOfcvJ6nldtPykBRny
MSIxNNJglkLyMBUCODHtBv90Z3lNjYvwjXvV3NGBjAzSthbfiX1Nj/YYWBaqWBfj
JX6E95ORfQIpSHmWpeUFfNeYrF6q6vxU06emJ5v/IPwcqTfkCnZTgjP7+6q9aX4k
/RgByMMVwrRsGH8vNhBvfk6ZkJBE+zd+HlJS2CX/l/Pn/n2azr8VUCa65BuQpsky
1YlRWD8ptOuTHW1mMBffQJMe6VXr8gdlOZuk7zwuHDHfcg6TZSP+oSNG81BNmfud
y18xgQQXuQCnCJdPaU+N1uoIFSaDdVMDswDdvT8WBbMED5tZfmM/N1KrM+/2h+Yx
nZN06Cdok1fgGJNs6YbdCuM/g+f3m6SaikWJ71rEmdlBzon5hy0YEhOrtofjsPIK
tv5RRrR1Ryt/Yc5M6q9n29S11qSaJZ9RFBmc/VOPzsQLQsu3/XAE2DJcps7V2Kc8
QbsC9AIemHMztkMzcwpCwhMPuzxs7iZ23wgEgtwLisRq9zeGlN02fSjEwIGj6Un2
YxLFrJLEq+G8lfwrRGU0FFhBiLmwkcfoQvt6713uyqZyytBQdmgw3irfmZx71mz2
8zOdd+7GTolMfLmKK/Z/SYaO8+nkqSyV0Os0LLrMTZk+gMUQzO6YtViZhkwdVVnJ
Qm8Vq6TZT/293DnfiDzLE0vRXOpvRTnAks9ZZymHDLmKN74GqKbB2Z8kxN50BVAw
zX9fhnTC+L4TxP4g7VvXxcFfK0HKn7tbuVmEw9ioxknjSHc7Ju40U0Kt78k1imIb
h1HSbOhdrNhURwY/kSMFtnj8GvdV6emyMLUrELYbFDPn5ZkC3+JGDFqrWi8yDCoX
xLOQzpvRKf6P9DZxvw1ujO0mjsR6T8voP6mA57DtAIiQ02GvJqxaOt3rNPedMP9C
tVrD0Gmyv8gpQmHC12RtkQn74kMW3/i4RGuVZnM/hHA5OH8Uyf1ahFKSO7NoqCux
6KV/FOrBa7XxLxndPc5kVlroPrCW8AnkwaOz0YuT9cqkLj/zOJU6HBloMBcHPEkz
2KAxHZCTCLPAp6BUGyzA4NXZAhhQe70Ja/ui7zbL+9wulAXz2VeNghoudGfeFGZD
B8AxVwTRgcv/CQz504QHxlw73Mo+1aW55rl1HX7Zg6UaxTVQ/Y43g/ZhSP3L4QK9
5kmSY8Tm55YmFcO/8D9coPfLh0fQBrXuB2IeJSrbTEk4LSJ4udsK1/d6w/bdIxij
zRZ7EtGyqgequp0la5OXW6xuw+nPLzMkqNB8zptXEX4i6AqU0HS+g+9IPvlVK2A2
nOjI0NfL5DIKMxVlSOfaYFnWef/LDK9Qvr3OOfg2xuXyWo2tuK0qfbfGbwg7lUnE
szOKX0gifb0RBZSATBEhf82dvXJlvfzyCogWRxuOVDUqmhq92Gb+DeDWiWu2MqdY
4/9iMeigvUvKbxKmhtpsgeH76L9fnnkp1jyp3pQbR0yyT9J+zqPK3xsg9J5Z3EfQ
D5ElqnMSHpfCWOPlsPbZ/czelzGVX1xIIRHLjoDK8XPCSF7nYAQEuhszGsQRDoRI
CUdseICn7T4t+iS+lEj7Tlvn7uDrh6cCu1UWUHgmvXUOVWqcHuFIV01XaMCVP2so
llm+QWUuaGRiGrwCrLDgdNrDKxS2FWDX4y03/xhrX8KGm1yymdOMxrcmoYWBcmlI
v0TQswn3RGLY/gYy6qxalR7hfE+0WcJZenBLRhZ1VpfN3ZWc3Qo9+lpJn7u4Y885
MEoCYNDXf4BfvcqqAy19BZxyi6tdK3opjjqjmdvc+jXOEFQcTAcnVfrNJPzSQGIj
v5Mbm+1gXK3mGgQrtiC5mM04qjXg+xASBaaouyuK1+XeRPbT4CsMD0V3nGl6sFOM
6fSlK7xf4hT3i0/3T6sC7ZaSZejxQHl9rS9ZOojTMigOI5b4E7KmiYj+LCEiKiZ1
XJ5Mp7V48oMWWt6Yo25GgQgslpElODl5xrQdQ20YI5MV4SQEDOOBr7xjnCgy7xHP
ckv6dnkkiGpU5KyW0a0/jnYcST0lkllwt2LTbp5iWMA5J6f+HzHJ/FaDrdmq2vZu
LCktA/9zEco0hsZRKgBOSWpRcBSOD9U8aXQNv51zea7xp6e90FMrI3oqsdKEXUVh
3dUfACfgBkPuzLGrub3Pmxd4ZBan4xjItcjhiDWyWRpgLwqKD0Y07L6KZy0mQWPR
qczRQ5/gPWuZtiLYufIUQ0bLi2W7i9qncQcENhUjsQ+5e6GQXrlLxOXLUpvs27lV
By2yw3uTiQwQlswfLfcSHxXd2/HhW33aHqkG9lVU5Z7Uk6VPWQIICIvLr+DK7nLf
HS6NDIm3vrpVuPAtlhFuA+WJ/qXshZsh72Qg+3e0+54I9ErKdLTt1DFlbG3DhxsK
jKlPBOFCVHbBULn6K8RAcHSJ7tal7oJdrpkrdMaoPYre4LXE2esHvjBnn1pocsK7
KnSR9HsveL1lTIZwsZqjrxY0wHuzS8fW/8kyzbLyst2hZ+AX7mcBohfbQpidReKB
McAqw19pAXB2StDtp3foXEiCI7Of0eIRtzMuBDlwhIX9S2bRrt52hVM0Nji5VPEf
gBGXpBtFMsjr0WJPxWUELm/Ds6ZjvV3kZ+duQapa4/zuwZ56Bwd+LMDHcAkYLB2a
MY5Ap7EHSz2AUheTFChCMQmfFzKhbk44d102Yp+F2y4H4nhS2BtfjF3yGQgr47d4
ozrOdUZ3T7JGTsUSAedNdjMpfU3lHh8DeU87dz55BtH2UZS2zhmRw4ghLxb7Fb9+
Apx/TkMNHLyEn65dBHkifA0Sn2pyLNB4Pi9KeG9uc/neRkcPMVSVG+HyWTj2DvHn
0Mf/kyK9ckllUv96fa4DYGcE/c0x7Bvsyei+GPED4q+pu7hxmqWaG9iFFoqHmVY6
FvajBEDbqCP8eu7P8zMjo393IG/g07W5GwrYCbFb0pJcHFgVrfHDhB+HIkqywVuF
m5nWGaoiEFUl6T++9BRT5zzvsGAaG/ZEIqs+VrIVh7T4NQSAnN623siljzFj4cBW
AAwaWphot72W6Q6YnaWllJzoN6Jy5/SyEbDUGeafYFnCvqeohy01rmQdQbB23tbj
w3be4DnNQ9+kbNE0+jp1Ehhga0qVw6HGEoZ2YIKRzOAIGv7QzKWp+QO3Q0+LruY9
XiBnwpvRLazWIAXfCndWZPyetvEln/o0me+euy8hEZfkQQPYsxD1Db91ifmPbSRL
qJGR+WdtiL0aoWlOUwRBqK8G8QCEzYhgq6r5wYy5Cim1reAugR9ZwMmqloO7+w5T
W6uUPLY69cIwIp0HhvEix4ZyJb+r7xD8w2S0MFG9sgOWD9+kBoWYOCVixgww+Z7V
W6HajGwofs8y9HnYNVAydOCeHOm14srPucCxXMXmRieRrGQBShor8oCfEb8wz5nd
hBV+g6u+5IDK77rrMo769si+AZ7ALgOHX+8rg6pmjy6xBvTHOUpVp3RtlhdCFu22
PI+8CWsdrXRnYuZjGtm1pAtih2Anng+Uq50hT49IREo5d7q/kwja+3DjMeKzyw7o
pmrDmCbibpBf9I6Z/USiEWJZbg5MluF4uRdE8OH9o14apnhGrcwJoD1dUtZ/0p3O
I4IIxp9EIjx6JNk8CQBd9hGkCz/7FUkNI/k2Xr9ss7FCJJ7/oBdR3hqO2Q9kamNy
aOcxBV7dyck9VIGxsrhFnIo66t8qgHIXdMPw1UisRck35lziocXYy1EgdSXLao4P
Q7BVRdFJ8UqZiFSKLAISFBjbdb5agu/+7z+TdY6d8mahoclWA9n/ShJ1oohj/jc5
CMHQRZKEdzVnp5iEq8F1UIpEyhP5Ay+H5SBgTQV0DZoSLAUKXBlFuQi+vU6VBHFD
zOaLtc6f1fj71aSEi/HNk4xr6bzZ2yzyvakjX1JYjJnyavcSiJZFYB6K+ZqxoplD
mLIsvXp2f4jVNNQFs1ZISDkIxM3286tu/7jSQ7F/29o0xLYUqou4Qk+T7seHTymE
1qnOTIw0G6WO1j+Kv3bvnjnyJ9uV2nV6B1XoaTdRnVkVW4/s7fsMau8hfVH3lha/
/l/LFwt1w9pluaalerNpKaXXNm+TBwyhRJU+04T2g0YQPkPKMmQLM7gkboqRcbky
FvPOGOGkqEr5amCHlVEZeqR0J3PnpjtE20bSEmz2iiuEzu/r2BAUGx3L96hMvFlw
L4JECdeKW7CGJ/iWb5bRaimmJvwqHaptZIOr45EtHHCcnodDBLGhWH6zSxDyDKNP
UjKCkc02oQkRIH4hsdHiNHHyIxuJ/FiNdlN2QihHEeHA5yLbZXVr1lHepe5MXcDf
nBju+Dtd6RtTk40dwW8j9fmF6701Q5GQxFrS4dyCaF54JjpOx1h+yPfGEn+GB9SQ
dF6ian5H0zS1vAzxRjBH8V9N/3R/vIEj8n2C+MRM8b1+7RuStE9RxuFS67xthj30
Nu4sfp+aU29UvOqW/oQFyBTQZ+zFT2oT+QyZEjpymXAYD0kXOO4TQuLaBBkaviEq
y2bYqbywiBp9t/BacpL9BKKt36Kf6yt9ML+2slc2OsyrNH8tqezRZVO1b78nXmvh
BcyZ9RO8LED6K7a/VOzyaeXISN5FV2twBDvWwiMxuxNyDoW9Te/J8W1ri70uF5dw
H5joU1YXGyGAVeMvCbITQJCA4xmUTEG0ZYS1bmGlnunmQg7MWKhRGi3LU+R3KcuA
YPcF1ywYXVFe/HAeSwJzzyeakhbcj/tzJQ2t9FrsP9JCPUm5cuUBTKI0FYLDh344
TOs85hgDydIzxFc5HJJCbbZM+rku/DaZv2dvMSRBN9a1otH8R16m9mAbzx8+e9Dg
7wZjBS+mk3wIdGJa9ehMQb69ls5dnMTLcXcZ+mQUahthLr9K2kRMX4Nsc+9gNRYC
Zj3DbDj4cydTDHIsOeyBeS4QDmxHiT3tLX1MiwMejloOShLc17s+NIYWsE3sJwqa
3WAW3P2YNozF4AzT0lDABZYUOkl14ga5wHAyhNQ1FcYvqwkZmMSbhdIlrWgUv2+/
1Vdw1Zxx3z7HzqTXfbu15Uth1i7AC1WgwC3WaLDDTUS4Kb2Bq2iGBi65GfLUOKEH
VfUsURu7SWhJIg/Q1xiMI3PyUiIkk7Pn7CUaUc0mhyR49JDl+TdI93MElZwFeuXD
k6tCyy0mekD4mZl1dgX1thIt3Zl7jipJPLrecgG1DzMn5aymBCXvQujEItdEN55G
pvta5VTTEF3ir5sVY33WY5zhfNvYeLIfCvBbtZLewxx2WclRrS84HuNpecZehtto
fVlvd5BrQGeN3DGFgTemukByC5+0eIjJfGV31zVxEbNOxkTGqsisvcQr7x+GivSU
/N13qfvqshRJaq+EhWG1s3uTSvhpfoG5mGpfpxw2SUPuU71/wkT91Kb/yowsByfH
Ka6dzT7b3+Gm12DLNqIrn6nnmPU+CXhlUD+l1EGVy2UOtTJhqvcrlDBkqaVIL0sy
2kY/fQ6pPROwMTbFhIULsNdLX8M8E1m9Uq+7ZSPDuBWcGP3ikzUNR/MuiUctBic6
sjQKCZdcAnC7aEZy/xhi3bLdbMk8b4nPNPNf67rVj/yXpiO/VYyXyYnUXvpfMZlv
eegVJBDFpGp2hMuR17r2lI//1kTDjT4Qedw6e9+N4O9S0tlCradtLOUKhDYkKaF6
lXBn5Wv3Ib1dBniHY17mZD6FfeyZPM97YzCPWfqZ9LCCDUw+Our+ycT1g9AshpV5
OAG/bAHAcegm7Su2I8EXlmQbsmiojUcDye5iXlQCNJjj1CmW6Qq56QY9YFQJBEUI
4eKU3BJboG/3CJVD3QdDwPnpxWFAOtkOK4yXDnQiqBzUp2jrI4pVIIfUZGHSI7Li
JcolV5Ew1ibLp7irYkAvwo7bZoTJXpgpHl82JPr5OfjvS6ujKBmLgpUHx0dkNoOX
0pit6obt6LTOWRfVndY3MpQIQrIg5BiYhswUK/58kXW5n/lF8GFrzZe/5JrK05//
X4vWVp6rQq7nhzBuJDYmDlnyc4MI6KaN9Koclv4eLqHT3qc2i4O3SYS5F8sDSBLO
FgTz45FBfZzrd1KHS5iN3i0ouOLVCo++JUJj08Fi/i30LqcKIwNf7YPUJ16gBbEA
n+irB+Sru3AZQ1fXDtdmxi0PcbpdxQLxs3dQLPYARWnpcoaRxzY3cYeF73LKFxNb
72sO+b7K4adLpZUy3JVbAr+DhpAT8ZYUnU3vTdI14cKasAPRTpETV6R26wVuKFUb
PeoeCcOj9WNaR75YLa5pV5qPrhI7IUPaOiIt9pltY0rFH5YiUNbCW5NC9z9AN19S
RamYr2ilEWMuZr99cgems6uqGsi319XdoYOPAb9SX5EAISYCP3akZSBIXU7b68X9
xgHUiLAwwv3sPX92o0ODXC79kj/kwwjSpBF+wS7TGB11XrB5p70cCkecLtPOhc/b
OHkQsuDQ31MFW6izgUCJi9bglwFEmSTV9fj0L++lnStVfpKFCLAfEwp2zE5UVPfD
bTY0uXBjVDuH0GInByOSyVkhlLwEVIskNAcnfyjIxoMW/pHYHPkknPzDQ14xl8Eq
FAjdcyf1Xoh+gT7JhY9mgeeNpogHZwTExVKKpz1u/5lcp6YlM6WG6kQfzC2cdRD6
WSnc0s0EGJ6J54lnQRGNTJxR9zpN5BGzfgsid4saDp3ax/i5WZgV8T2f1GBALPjo
FrGj2PSb52rkxUR5kU3SuG0WclURJBhDu7zfj+E83Iduh3947BGH4TLr+bq19Bw/
YdNmzJVHMrmBvXX1Y7p1GIlIIlxzDRfGLdUjzlZrPaUG5MqJajF7jmILUNUaM3oV
czKluabWpL6ygsVqpPtT4zonzkICsGcIAqbAQ85SKl8ntEid2WxYRUemk87mKBHf
KxUUJAAsd/11sdx/U753MRGNC6aVHjKN1jxfS0Nv3qQ3Gt+PpsnbbkK2lYLdsGil
/dOfo7bjKHn/Ukhbw7ILM1cMhbkAR82OcWLPuuCfZQ1s6dFDNsppRer5Vo2GjXoR
ZzMB/69Bg82i2+2f/Y7ImEjNlm12JJVkbGAV5XCCxS7VBcWzR11LO8pCbvY2QdNq
IGV/HW1bhUb8SJpwW/nc9WSZtUTEflmZZZc1B/6p1yvPr7n6LCGstzux9jt2ZZP9
IPPkJ6b08pJiDvO9k2aDpVxIBuzu1o/CzV3ecC26yrB0+cxc+P5kE6lDuWAvnSuD
gnu8cIIHunPuyNKFVnx+owMqjBpuJCBA413OuXnd3bk+YZPQ5kLByF5WD6XDg8Lu
zpyETV4GZ7vHIUl3zj/5EaK2NqGmhTkghOPsoHii96rk2aARW9+yuuBazv0GIm/b
Q7X5PLT5bNC3E4ALQKFwJSNref6oB8J5JOflNE6diFMIxyvBJ5eMFmd5t4yeBN4N
qNNMIGt9YzIhzXr/cPUZImLL+rgrgGyoFgvzWEbinrzgYjPdZnd6724LLkBKjZKA
oRBRAjnnjuT0UH32vizv/tEnQP8j2si3aylGaTrmz2o0sSliHtNu69RLon92ZaqX
5j1sjd5hGD97WMPXXYaAk2vKtsP2mdAe4a3XeJj71L3KmZaOt0haoCyeEaHoUyxn
6WMR/0Q/5e4ogUNxcjfIZhLunw7rCOUQZ7k8PaMzydMglrg+/7gqU31EWYP+QYwo
z/xEYgQZdgtYB//RFktYDq1SJ4vOb1kFMBRamSFKQqqr76WwkkNiNaHJEFIrDjr2
ZoMB+AIz3hisVkRgmHAam478SlIlocM9nZ8SU7SmN4bHdb6qOH5r7rEJGnbfxaOe
zT3wGSNArYhdfHS7nXarar385ieBYarK4HPo2vBXVlkAHEWBNl6HfzP7E3bhsrmT
GBziJkTtXLkmUFJOAKWAkpnKxPVx7ARs6idZGHN6gUK9Zvafj7UH/mFHuLUwysLF
awhsBiwFqCIaSrog+DUhmlSJdR3xLymV+hgtHVkPh/Kuh73mKWagEn/Ebp81i/2D
apy/JDKUcRfkbN/jDrRDylD+Rv0jWKggn9/Nmc+AJUIVF9itolf04gVHd8PlPitW
Ml04DMwIonQRqUejM5PEQcoAdDNQbqpZUrhn64lTfTxwjY7GTAL48W2TNsy2GGYo
2mxz0b2hg/IWbTW5hy0O69xnOWmPsM35hoIZgPemlZSI4nwOWamnI3YJsxKmDimE
jRNFI+FzbJvVvcotKNeYoliMTSv+vjD1NTWdigcWMaQhZbAQQhhnSeJ8uSX9dc3F
oFpxIFnhpaIxg65iudMx2aGifghYSrw4F0UHr9/9itwBynORhQg47onUJ+6+jHM9
DWxj+UHOrgMSbjdP8Hllt+cN6vsoPzhFZa34l/37owJ/7MIkBVqZ41jCOGsBkKWm
lRBq/wp0XTl+A1fX7WBMTeqdavr3uEHPuX+deAzptUmd7TchwfkTtqlBECB+GeIp
NU9GBwX/SxROP13S/5RmeDdPmgpTX2sn6CPr7epCEQDf48lYfRPBvxu8D+Iiundt
0QFg9pzsJV0+nCV3e4sUup0oXCdD2P5KVfooktosZUfsT9smxg4G8/PadrS2V/i6
h1TbuaA+01w/H+RHvz2cCu4odBuQx56dHhk6IJydBTdPWV9lVz+Cg9rDcVoT/PZ3
2WN6teJ8Q9+thruEwdatu4VRsGmHate945OTBANsriQCvAie/u4fmTGrLWnLxnfZ
CvBViLxUEKTtLaMNvNgGUHGNbkk8fPNan3oJDBcUX5FmWnzgFPC/eOgVB4M5sXRP
Gepl03YWY/CBUd+DuoAbWUjHr4Z8G5c7kD2rQaVFh/JzCzRAx64aQPyQCRBOb+eI
+TaVCC136KYgNmmy8Xk6VbRvp6LqjOvFWHsDEVPKgYB8ivQjlsBSvXvcvHQvXLKF
86Ktb8xBFTYL+bJQevuQJ9xEu45I/Q0XfusgnjIurqeDBEWRCuw8WHGfcchk7lTs
3Fd3nYkpGEnBeKPh4d9GiCicwP24xQBpT5b6mdzw7Jpn1hvNTIOSwSYGAUZ2FMRt
TAnEuUVOSR81JNBcCj9v/QKm4NwE4uz2XQjFSykwCjODfJTu6MreC3AOWqTjtHiL
0KyCZt9DMLzaqVrxJhPWlWscZ9KDB0khGA/XYVYDcn1vbGgk3UBGHR8P5jjHUe9o
ahoyKigadIsPI7GOfOX6DQc1i5kXBDujdyjzTY8EXegGki7NXN8EUN7PUfI5gElQ
uzabsddvUlX7lbR6Cj5LTCfci2aaD5TixH+7Q6OKWyu7J9S06isOEKiH5NuZEoiZ
XeKCkmdavN+SXZ7Vs4zrwan/d301FJmAOOtwMQN+incz4fx311ITtSiwMkzQ1muh
84wAoCnTjTdrS7xJMnmm0/uVTxkT2HpqaDoLpNKsT/WlG+pzCXOPGlcos1zB4ncg
knvC6xUy8ZCLpr3whX8HN09Nc2BR4Lqlwzm4DtHwGo+lmXdpCG8J3pIAemYtmTwZ
6uFHQwaXSX1FHeXOMllh8FkYZlwWgVW7Cb/rIIDqdYeLCi+dsUkxotJkViqRX3Rf
7dfadvQzjkraygAkytd3bAQTCfhfYmmMn/LkixlzLcBQiJeA46WYo1zLgHYq7rEw
h4/4VxxCjNasVqapD4VOfXInhW8zvCk4/7t0hVfuxVr3X4yDbYZAKkzfXHlPYEoK
DCagLxciMuAvsF38qA+lqmuB7YXprcLlJlC/63DnwbItS25IKqf5u4IdIFlRZY/A
S1ZKjmxFDf++KrX9ze8wEnsu778zxrkgcJz4DIQso1jRNicTzQ9UvX6jSbfltviE
qn4DBGEtgOcGMorERbhDRG2ojpfgdS39W5ZQwJkHhWJvsQywFEsVUr1KrEIMktpI
5Qs51Idty/WKJEhUB/dfPdCurI8/tWP4RuuZx4LKFFv8qIqgLETDL7JQSOcKpKHw
aNcAIMkGl6yhEHZkUBsFbmB/qTsZOHc6B4JPS/9FrM0Ws3ZbVXc+sWyXn0BM8myE
0VU6vGqjxnlRfemQdhBjt0p3nCck5oYB2ra63mi6G/lUYBL+DusYI1w508dG0Est
QDRomjCVX7tJ9OvNh6qy5h6/1aZHGYaIKYdu5rS0ArmbL5Ksl8ks+9p/QVcZx3m8
1JDGEWYT9QliKQjg+f9oagpMcgb/ZRRTyvHpL2l1XNQHiDHqnAaAmR6yeBycJ7an
W/x/GhCxcASOQrcbk1DiYmUkgzFU8jJhJKy7NG7EoKr74HN6KHN9GB2Y1Kh4c3Gr
P0838UWXpmin+bRMBdBjyEAPSAOzbR/jbc5nx+zgGplZvd89jEvcBD2hndhJB9FK
s1eee/I4FHSdI+iC+5v7lPvC+pdWOsOwZpJEgHlPJrUiU6SCbHCDK5FW3F+5J/NX
NTTXpGYM4MmTlJJs6TQ+8BSfBJRjvhZ6kPSGSn5qsg1/s4egJ561pdgwJakalDfu
QdkJq0oECdk3uWQjeFQzcBkrAJFkh81Xi/fn1Ntbkjpo5wJgn0uqmDYC4zLEtFEo
W8BjWMFvcQA88j7RMvFQAhDVHpqoaLkz1WYYiBzAryXgBNs/kMLcArN6cUNwICmr
08vwaghwcaRz0epaF4SsK0x7Os8dBbt51lmypBqx9XJoZzTR/Mpb3bSMxJdBtkNz
malystBhViJ6auPtgtZpm8Cp2wkbhiFcNSZEcbrstcDRrQnykdD+VdTtnizSh6vg
YHSLSS/DkzMqA8BNn8Qmfa+tlFAw40oAYK2YoVZZ92PgQvnuis/cLZTtkYt9eeTC
Rs+/ZrJJrbrT6IM09nPD76ebz5dRSRmTxO2LocN91L5CPpq1PB4nGnMM6ijr6ig9
jypUKyzAj5oxHLf/X8zDjIXLCKo59XoazALDqdxBWAGhXR/eVYXCP9jLi/f1Cf9W
CdYaHCJIpwOBAChRWM4dD49mCoqkC2AmpYX877nf+RdxY2V2NEHQ5HUEPWe5TFwQ
IvbgVtRu3vIFB0/gPbMn7mPBikLdeZiUMl55E/feF51tvbdHabbM56nr2lDEX8l9
OG3zxcIu7fHSwBaqz89HcmM9graVKRKHyJ/JId5lpM8DG3Ne/74z8uj9BnAnwO6O
5/95EnGgJkOr6g7PtKavb45MduB2NdImjNUyRELDN1FiIG1JFKGhVPhIL754WoZ4
ziW8EDLnzpOLXbIO96o2CJ9jchWh0Mca7j4G9xbpLEEP0cJHbGMpJ4ozMICBpXqY
n5hcSAGxkSVz8qZKeYovAgrzwHiAFVh6VWTs5iKfUhiI83HprnOnCHI4fZTXBKKh
ZGeJYC8PSGuoTEs2uKXqlJSXgEd+qFfkybfHhy70XpWmlDgtADt7bZxsvOTnM33o
0sNtkmjlA2ZyreRwK5lo3C41FXup/9fEj20ICg5Nx/9VO3lBfnl6NB2We1m+c+HG
zxdThurpo7DohAogqZ2ZrjJf6bC03lYQ0lzKK07H7kyadR5zpWmx/D2ILGh0K8at
XG/cOW5vvKFwQKPaAJB7xr2g7ZimV9nLW9yiOnpwHVXMVJwRSZqW/6OMRT/zDK/B
aQslhH5QDtgyJqsDtM22PrLSBeqyoyNaYEQVCSHD8SFBbRKbkPnuwHPuA9LwUi6d
CjAQNKlzJcUnLwC2cgyNVEDnPw1/dUSzEUtt+EvKbWIfP3fCcPnjUtBOhHzTyVbi
5+ayR37ks7w3dUe+XxiK68rUc/Nd8kmwPBK9NijrXP/6u3+5OlLzAHucnGoLuDX5
mixtM5i/Lo8zmfqlix7S5oEmMymo28eqyBTBXHMuxu+8xVtE/30ko5loQD99QkhC
ESqMK2Mq5MXHoVD1q+zzlFop7yrSNz+wqxChVN2OyMAVBfBU8cV81gNlXgEXmdVM
jutUSdwLYK6rcz+gIpvgRwqdM3auKGDGpx8knIPHuBjH6ob52hSGDDI7Mw1rxc8n
DPN4euG5w8mvd4swgjhj3aSNbvo1rr/WWtMvpf4PVk8E0MV5BSdUmlxYiCslAtbu
iusNZpShcuOcUCJrppedXsLnQfESV8MsyEepSOGaI1HFxk8RDzeKE47l+vOzjN1T
3OGSJHhgxTt3HhWIbe92ORYKb4ehOhyGvwBGOLkmXW7J6CYufFhUAUiBG6qRRgSS
g3mTi/QwjxrVHlGL0JA30BBt0eBp3ftBF4aCHac5T/aCr3UKcMtT4V0osW6gyNrY
4JheS4kCHVC2e2aZlCz7T5UTHUQngYn/WpgVA7qRuKkbeOdoC4k7FxPg21pIB10Z
1ihCU8TfnGLxn+hFP3/FyxVKgxUI6OvRIZ3qUHkko7TxU3MJEM1vCUvicHkBhamD
r7U4Wx2qvNAFQO+InN18slNV5oEyw9MWFOpPXivlZDOxhG0MrTZzpG9U1kqjeeae
RZAD3XO72NTzkp2qlCMEiBEA7EkIuyjs2T16J9R5JOHy4M4MNgWOuVefpVbWE4xK
8dlQ8QYf3o7MX9X36Lyt03AkllODLjscpMwwGrKRdDDCns2WiiuDTn/ab1tQpbch
TYlUdy8ZKbKi9ulqwJ+pmJtviIKXBBMakqWiKlto0g6d+NvUePvJalwYw5ZLOC8z
1Uubitk9exWiXfzE+o9xw4pWwzGfDk76jdOgWzt/1YkSFrVB3MUrftwWipO9G06T
41WrG4gv1Gm1FZ/JfieHNzeYleum2wleQhWp8Pq1tQaUjRv61CeU/f9+vDPJ/yN6
h9CSOsZ8BWPjeI+jBBpQxWAWQwB6fyRULKVxEucBvLGggdyVOcbitcqZaX+IA1dW
c+UHXBgLy/cqHJUy8OOUK4aSloFJGHETBmOVNzD+L7rmmEL9W0zVcW5j492fVjnQ
wR1ZZKDGAGkCIaRViFwixpvtCIiUj6stzh64Te20Pudxp2BnVFk771/9VlqVuUET
y8x9nNlKgXtESPdNkAHrCjkR9F7pF2HaHnrVcJBx3+WaM4PzzVMVFslw+QUkuXTn
zQppP3hZfRhq0m2XpIVncm18Ysl96Lrmu7W4MN+sY+wxmkfVfnZVeQKsRPbFRWhv
C8y6PT6d360KurQ0hiyEy6oz/JORFFMTuguCywHHufNWc6dVdhlrsKHit6tzHw1K
srpgZgNP/ZCYVH3S5Nfc7I4jOi37oOeNH1LOaGi03ksiPPmScKma9SNPhRmK5cng
Wuaqh/aw4Ji9f9dvCnWJDjK7FNjqKJe1qbX5Aek2uiz0XCy5uFB7Mgb22MVFLeId
4q9+dzdf7K6ua8oAQi4gUpSM/oM481NE+c9F9Ph6GX0nc1jidJ39td8T4+B9dwzM
ANZeEfdwWx9Fhh+VN9yodLF7OHLSuMu76SBsEfOz1TWarkgoHhmP7bCgpEBl5s6s
2wj4pB+ZHorhRQR2IkQJPgmFtj7kHdmWFPZKJpstnTU8rFH5N8dODQp/u4qk+Oz9
9+K5PFkQmfpX6nftl2rBaJGvKAuTy6poTsn2fxwAJ85q4/94y3eYYcEj2it1Yzex
xgMBe7FqEDr0tQQ/meaE5h40xgmK3qdvyWgrhS8xgtK00KUyG7y07mYQCqyDasdS
ocSLlSqmwgz1+5xg96/39sdj8QIGUaehT5Btwsx195MOvI7fn/EB2gv/lt34DPXY
B0OW5i4D0hO8sNeJwWdgphm+LRNLJ0pRnGpHfdBSGIh+0qXAbTfDNthVgIdHz8oe
7OjLvFcwGsaLvzSkyfdt+cPiI5w0g0lwUX4p+MHrMOQYHZiHJR+p+OzvDZ28rPRU
yOhV37io9KhpKVm9FaBfKWD0DH+XXfbEKJR+ihK8r+uNghG1lroOy8UIfnqu77qR
3loeP87geoIuBqgTOxwE7GjWs2EzcHjc/ZcdQ5+zf+DV64UXkI5mlDLYrXT20CmD
1LsV2MePPCtVgSwm1qYaji0NNRuLwi4757TBim1lJDSVkOWeMPjTa7R0TcGg8QGr
qaiII5I8+y7/Y0EXr74OlnwQWaro/Ck/hy8gjdMXpHJbpJ71NlweXNYM6noevg5Y
7pCD2oi+fF3PF7s6/NXb5D5ov1V0SQRuFXLv/BcrOQ2TUvnm+szkXZGwwMZgj0nq
41FLb1Z7pePRGIOAjkOrPRbpTt+/gVCKDoqtHYlkw4GZpro86GK0Eht5ppqXMhtg
VnHaKlis6TeBfxayRGDdh1WH6cuPRdajg8Gfm2VPExz7Klug8HOKzWD+zZ+inOZn
KT4obRPYj0U0wj1Zw1uoLnVFpKt+8MUBksjRKGs0AqdG6UQiFCDqDEN+JYquQoaS
HPEMWRo82n9LdHy2HorVQD0hdwbuHO5+kdHTuO+VpV3duIdt1IO1Eif6iB2FmqZE
5Yubv2c8QZiMBtTN8UtTrvysUZt8ZnhYisGSSdy9vH09+nx2r5vYt1lAQPVI2V2X
lsM1vz1XM+URJS6wOUutVdRmzaVf5TiRUoEHkARjvrh4iAeeQ3iuccXPXAZ+ZQxT
bMqSqboq4SnAiB6Iu3V6buPOi6zLDfYfw5q4+wu80RgJk+mJmPvNBNfrIQ/jT78B
tup55E9S1xzMxlPxLJmjvs53aaGbPLuo/cPhsflY05CTGtoDFPS9HiTzamkmQ7UQ
tUDVFNAvaHBPYq5F8MLhi6eErnMrCQsIV6GSCg3mamgq4fFtZyvD/iEf4N1PZC0k
h5qRDFKKG+47+0tJZkr5Q4gMXwgg8SOsQr7HJjeqOGtfW7rIk/FlLkdcp1bTlnz9
HQrn/uYwfZHcE23RJcYN+itg+Nb1R4qvwkBW+A8+wyL1k2qA9LS9CJSH0St2PoZe
/DKUr16xi1goO0xpd7EV+r372OimzygP5HQcsJxvw0FksTGxITBZHyL65TdgHmdM
rQNoqaiNcRy8HXjgyA2XrPziiF8HVKre9Xrf37beb7Soecrgruw6KVf5ADIOHYS7
0AYCLX49NycCIDVPpKdos2saZnrjJ80y3Ejvz4b/07kyQ7icz8ydEsMXJn6Bx1Fm
UQmtFjvy85sVOyAek+eg7hKbVfuWxWj1A/5U9vv5KXiY1ly6dpGVEeJRPKOkuVMw
u42YJStNG9VvmnDkxBQOyra1Hzp2jjQoROxW9pNBTd4IZEr+DIL3xL/SkaC8ENW+
uFaGHm7hQQAYnqZ5hoNajqve/BrQuYLiz4oxvW+XBv3K4hnSRgrkzkltSV3Na20z
s6Rm/J+Wygz7OL3Ui7AwoL/P8QFnSw0PyHMCq8KBLlPRiN2nfMPvkLEJzADuIiRN
cjob0lUnh/R1GhB6WEUY2KvQjsX6T6JsI3QAapVkFraxnfbXK+3qwrrXKg1ESq8A
xVK/JfnLpUz9MdiO4sdkK/GHXs/6Og0bQvQApF5eBSR3JiV6syR9zAZ1AqCLYG06
aJajkNN61jkWZia1lSO1mGG+zlxfVokhM7FUGnDadpjkVGVVaHBWpI1V3/uCQKcS
XthvEEg7Z9EHqjljPAdYQo2s4YMszeOcTwOTPgEG7hTZMGZZB/KtPQIJjjBhka3+
5jyGjciZPxAF1dKWKFUXJqNwlR0PGx7gfIDbLEUpcRL8iVOOTaHPUb8K+FUgfeL1
w9AvrZAtvkU/QJF9RlSp7vMAsjPUkg95b6b/udin26GBFzIDFqpyVASQtKwqp17D
3rCuwzAhOb1//VxJjjeyOchcmhL2dZJIPXHhx6juuGhz6dv9Y1LI9XB4JDYo8uol
BmGctF0mrwFdtWHBTV1ec7Y/J+4StGpqTbgKS+169xZtG0W8FnRiUryKI2KJfLiJ
e7eay04Mk6r7wxJ9g1px9RiWqiVsCdK6nJAELFrPCA5HdGxh1kuVREHUaBdeEcdo
R8Kq80yaaxqMiQVANJZqfAvu9xrj0YItBI2UKzf/05Lw/2vKycKU3DBIkgRDCzOp
Q1+zyOxaKx466AzLRlnZ24Sh+/7NyikpgVK13T7F++EVQwc0mVqHU4swpUC3leJE
p2FoflxEJMOW7TFQTuwx33cHJgGMmZBrskmj1FWStYMfrIZ/9jm2EEfPa7CL7CQk
uPdiA/bP9Ypih3KmydbMuVVP+JaO3/dCPehRHG5B4b9hw7sZR8JaLIyhukwfz7g5
J98Ls4FuB7AuNCXbXsg0kyhQeoh0G6DuvJqQT7BXHi5r9T/9cckxz7tluh+uqnJ4
NuHZJyvhIRQQ5+VbPANMxKM0rgHngtI8zu1hs6LijWqR293tZmIOD8W6JASC+k0y
Tjnk6gP/H5eeUwTkZTWclA6WQ7rV3TH7bBhPtyd+mwkPhzyEMRLTVaM12spvvewX
ZXT+V1j5Uf4sACpoSGU99OQbzZfGCqtGLsP5D+Yu0MVQKEj1W5HM41+wDd3HJpNB
G2z9zi112gnm4JvsqE7C92j1qEb1z5ichlA0SUC7Rh1sjOo+OooKk2dR6n0Jf03a
6qlBZb7pKxdbsS6zax0nN+Z05+c//OAT8LbSLlbwcq1O1JOdLQPd2xoKjkVsM9rI
N5TJqcviGJeeG5tQF9UNPB36anj0rD0RZZZuT5L+Y95Le4ldcow2xnWNeIHXwdcV
ddLomObYVOzmH+ZO0Rfz+YMmbFFjBDooJIreulkz4jENExIZqtgL89R2txsXYHW0
bqH8qnQZFlkXxF+M0ds5upoil8N9AsmoQT/z+xo8sDDZ53Gn5v46gUS/lB83oAhh
w+S3mKUDy8NEMLqb+dOonKqeswr83HMxniTq8Q7YC6P58TyP7FQZmo/rpCfYIKT6
WeWzuGgzDpgrX3AKQ0qWLWrgzZX1SkXkDJJTfTanwqFUdigibCPkntXx9DpGS6wS
eBe6ypovffC6Vy343N0SZfKvZsfUAD2en3ufUJSyJXep/Ge7zD4a3FDrS/2svzW1
ZYsvfTUH233dK98oHMY9DYOtct7/c41FNd979p8J/pg7ujUkf62NYkzf8Ymjj54o
Je8gqx9YosKaySpmUT2ownXhd1EmiYdZQpBy1PWL7TT4K7PA45XwWaBztpJfX/cB
Ywkfp0OBdmdpiAyd6MlNKYgTwkmqD3OzsQNaRkxtFIqx+SzbO0VjD4DoPyz3nQKj
mS96s7sWHUPDV4GNCRSYACqyp+DcGMtTfEGXruwljcXHyTJTORskcRBfeW2TMB72
aHZoeJkrdXtPB47pAh3grdxh7Z0hnd/0C+LenfyZ/YAXdvcXQathvFgIaYZ7fNUG
wbEw3IYHBREPlcQ/HVnOaxwmR38/immjRCXnPor+RujgfQVilIKetvXGC/VESl0q
6AgsnbZY9nCz2bU6mErv1k8DE5pp5ijE3Cat10ymnFGi51h6+I+WuSQA3tEHQN+0
/QP683XRljQ65CPs2Lh+Ox33KVE/tGgtRVxNfCBcMwAuvLDxOSoWxhDSZkntje2/
UEAfWEQK/FlI+wunAVHc+FjyS2QLSk0DdqdhRAVhSRAPZ+OBgoGQ0UDR78Blqnzj
ACeXl3rMSYxKmQMddcnbVKsyA06lqANjv2DxwhkycMJXWdUO4V3fIQvkkmbKlB8P
6BSr9yllfGcczyuArvz4vQLM3uehDB471UVyyMGzfYLfIkvcZNC7jxaHynOfnrLo
lwIUW2HY8FLA5amKWrJi5XAv01qn9FyrQhb2MkhQuvbzCM+E+GlDBXgcMtcoHnI7
78/0iljjmgsM32BVmhZEkEHB+INiquILIFOqTUyHVKURxursi0RgUoPgIxw04wld
QizU3QzTRloXac/jDPtChlZZSHXHdtavV5+fpvttetv0arqPXJYpP6hI2mGV6MqX
NNtfCfuzOKb1H4QiLEoyPMlBI/M4DhU5yLRZPREuZvNhz2jSROsuEHR3EcvY1r0u
6HD4SJrSPZK8qjnXWAzpg/hFdfROKrSoi31R1ByI/ZYc7BRwsPNHLAHlh9ycZugI
d0NspQMzPscVIM5g6J+mXLhEp14YeD+tB9dI65U24RmptxwgDdiuJZA49ejwBHpP
IOTrrJCVvlVUK5mpQQR68axRZ+W6GwmVnfoOSD7eQFlvltEzKgWXRUAStnDcFzZj
ShrHHsU/2Yim8MywZelYWNRj2hlHTh6KQ/blwnvW0mNzjtcaU9Uf8ygPwVzkagO5
j9NURy4ETUvkYlBxGAsJDyyP3esDriuw/kBAHfnuxUqjBdhs4vopANgRZM7HzWu4
9CzxPgP1IIw7exOAXBJ0fakytJ6ayaxmG0Ru+hI1J033hblQwgN5g7DlYsimSEhc
igaz9C5IsTQZx2M03+VrfZdkfE4dA3wSSvFdpOtyO/8ya708aIZpK942yh8X8XAd
PlvW/KwJfwNUlG+nXPVkLkSSsk/ycds1myvr1gJgkMWCBqEs6ujAiAmG3lu+49WT
O8FT0rPuh2CgnZiYohOxYOymhErHUYIK6SaC/ksPnlISH1DmmrC5lDcSKXfuEM3i
R0y86gA3n8SGT4pZbaAdm1G+2xaT9KybuTNl/JI0eBbWW0Pvl+dYwcKDu0wUn03V
ruM7ML8j1H0atDJT2U4kdGv7MhL7ILOb0SXjNHRMfjO/8L3yS2BTegCKMsz7xLed
DvUr2edMUIgxjTB0RQwJewK0Ag7Ts9rOx8uCrDOvMCB1W2VcB/yVtUi61xGE3qgH
8GSA/Fzoo0x+n3J9QH6Ooh2WoYLNLd9Zl8kUdTNpK2QTh9rSp4GLZ/R/mXVeqp5S
blJJR52ubz57kDf0ynlMvhjW2bGkZckj8Z8TgeaGklH/bfjuZnQxrKK/7rMGcQUF
belTjGcFHArS6MHeY98UYo5Xd9H+Q0L+OOzC3dz21m3Nqo4wcnr8ZM59yp79SAAU
Xl0uaJFVvsmsPrzrx7m13gps/q+gQjVWBrc2fsQ3eCFLfcieCkawliK2XyK0UTAk
uIWoIoS/Oz7z1GHr3K1e4b5kp1fmrRnBhdRij+m8SIbUAImw+rGkkroYuF23MRh3
UVnxkqHxkD4/Sam02uRTI0U6Mc5s+isQEDI9hBtkhqFTqw71A9V3TmgyJ/8G4WQa
7Vo/OMsMmUUJYKmJfgioe4AlhRWURJnLiUfoJJ8x0yhBNNZCF7MoAuSMeprkIFkm
jbnT+S9sYHjykUZzA40oumNoKouERQXPhzG5+U/fpgc/Bdab+b0wiwTrnuR3I7Gn
ehK6rOkvgVXaZSBcm9akzfwhzLgiMWlXkZ74rsVXc5edpQ0YzqyHkCSPiSg1IOQW
kS4IORkjAIUqod5eoqdkV0QYG8QrW6n9Xk4a7eM3KRglAY7/4lUqDz3eavOqZlqo
N21SYS0djfcvTIxHUK8/TwhiPXIvvJCjh9YRsEHknHjVdjCfOUI9dhibM9fnNpp5
s0MInc/wbaEI8IC1xJlKcz8nUwxkQhoIWYw/Y/8OFbbnOifcgAw4KXFduZQCD/PP
PhUyTQuxI2mgZYP/vUY1A70mgn9wqyRzWSvFQ4i1xjJ8WIQv8cW2NOKVrgh9jxtl
AE4zPcZ22jclmG/uYy+ESG6W6KXiSMV9hhmDG9OepAvNwp+zA3Dkk8Q1lTHdJA2x
eI+SqUC7XpcHwgB6EoPJlwql9aLjoOm6feVjNbeLyp9IpTA3niqwCQc0G7d+ep+9
mDS2pivuds9hvoVbzM2ZhSmcTb6xehoZcBWRExynNfS2ipQyl7kRzRTgv3H1nsh0
PayEDVr/qh2sWbeBd0qOlgMGEIJoHc6r40hITFPkXltMjFxgzBAnBwJwym74NCFK
SYPA/LSPUBf/2BF9LNcA0/NHukyQgtO1BycF0JU9mv0O2LG3TcdgbLIJliZRA/tT
wm7BWd2RN0d07sz8/t+djt0mkmpyGwPMF6aSyPmiq1ddFlfZrVord/wJ0fSted1H
AIm35ihGEXO7vmUK//FXbHMIbGnV4p5Bd0P8CtmtaP+BCwnTkooZFX9rhwnOIFfi
nofWGBJNaPnsVYKC2IHJEqs3OpkHW2d4b9hI0IyZ3ms1TdG+fzQxcp1aOUpbtV6R
aa8hXYBrZuHw4OzwwX3XgJwcGE34G9Z2haaE+wHzCjd5htImcpVTjQN3I82hn9+e
cRg87ntzDbo7uZDkFJRH7/Y7wOl7simHF1x0CKxVHJ0F5bQm+AzmMGRdVDfFjyG5
ne9mvf7VqxxDcshp1t0ox/q0EqJrvNdqE2AMT897WTB9Ld3KO9TzMoORW5KWcQTA
zgOf65asETHpOcGbMBvXIKeSVcFjrwfBHnPm49R8DEZw4AL58MDSL8uHjRdulEmS
QXuPm9aPZCoT953dtM4xxNhZx9w4b7/hkG2c6KKMhDhXFOyHtNfp8RZZHhv/4xCv
ZBbFYSN86ULrm7sYUaDHmai7luGTLj7ZBdZABG6v5KWb9fUDRXV2ZA3oLJZJjdIj
NIItC3OxmOXR5VzdIGkaqJiotmxb0QlTIqrA1X0vl+dD2T1M9FMtAsdYd+RFtKEN
CGoc6dI31JvxjXTPqINYJODpChs651Ms4IqrM9hr9HJ5VtRWkh1s+6+M3wJAoET8
VxCVQ++9ohzFdnIFinDpEzMbftOiUb+0drT1M++C4FHR0dhu6kc85QllwaohvUiY
9Uy7V3hCihc+zB1LY0KvVmoN5fhIBba3U5d2H7quLCMu7gEBGb/xbCVNFeIR5D54
+80jUs6Az2DBXOQUkdosf2dbyyjWp8G9Pk9A1nyclysU/YBWsll7AsiNvd9XiSie
Tl/IQzD8DqDOGCafZQ8RAuMxUXxOiWsJ1MLx2sOrUw9H/tmxE7GLz3GvRJTHWB7D
95s6eAVa/HyFYgvXoJ5M1Y84GWTj1WO5u9w/MxGFidjel/3uZYiApOxVL01VCApN
GvwDZvtfiiuUGNcU63fdX5+NX93/sCwJH25TS/wfixZ+QAk2a9dTKmUdDjW3CUgW
5+IYM898bNWRPx6rRzMowZXVKksISbbwMC1Sk2BUTcb3Cq+BTvZd6vp/BQWpC+NO
Y+NXw/OEnxGfrepERJum0H4wS2yFAMWZqJhET7BSFEbh9/50IsZkI06tXvbsaUq2
dXzAA7VJjh1ZBxB9p/QxMl4uaioSdLP+OC1xe/4eyFb+VBPjNDJgTTLHYGp27dAp
4P4CRsp7ems3DZC6z7Nt80JfJ1m/1cmSiwr/PgxD/8m5L/VGrlfn0gNZLCwMqgtp
zo9rNoin0FUXMtvuWFgG6yw5pB3okxjn6HdJhLg8yEsECr+Bg94F8JmsaSedHJc/
Ip2BW2jmqJoRLHHPnXMIDIniojDAAJ5JWOcs+1pKyGRC4FLqDi5ieznuIkBv+BbX
FMpmlNB8FX6T2Sa9ezVAcffD8jIQ4+d4QcQRrtmZ4bGTTNs7tUReBGqBph3kmXY0
rGwOltb3wBvdMtngwrO7AKIMwBDbq2UuRAzIKFn7Uy3vzsagbjeIo01aum2zhkHH
d1c0H+KeVP6c1hUCAHSYrOoQ+lNo9kJ/koG7Vt7s3CpTdx5x5a2P+d3ZeYjKXKhV
8GQcAA4B8DVWoiqgnTVWCE+1sNxDlK52cT00900DcM7MBOv4wRR08WLI5PZomtWv
H1Cq1XqLn+M/sWsLNEY3Lnk/r3mzEoNAwNJIuMz74r/qolZA5Gcmp1P3XBQ4OBA6
EmQ3zdYaQ0P0dIlnDk/A+IlRwTQnrIlJO3lN9BHoD8GE29Ju7Z/toSWK9j62AAPu
MW7bJRYjjHmP2eirrT5t7Ph5agZB/lDYcSQ08//AfY22aCxfmhU1Qcr3IXaNtDqx
loqp908o8ckw7uUB5c0S0DE535su+3SS/US3C/ABkB26Al1/gxA1ult39JpqKTfC
B9YCwMML/akr/IaKWuYZz5UFW14dD2CbJMIn+CYzW7tdpJHgvEX2GsanHBexYf0f
MCSNUZBC0XVaRSK202GsTSgoDIcJUQKrg3nmzT/ii+BUL5rtRTakGNGG1hGJvlyQ
g4fcO6Cfss/MinPPwJ+JkLdeD5G4S3/W/7SgWH8Nt5OsXHHQdMH/9dzZ+qJpUYDf
DfN00HEfFBqU3nn4/7vNzyztzpyVrcs+gSxcbzhMOvti4b6iJrZxId3QPgNRsdzE
ilZj+4IFDavALB8mq23OyAlnC2kLdMYYk/KXygS16LW1G0LqJzIbFYXpVkiZB6mU
CYAFT5Zs5jYImFNGmlfMfOwHGbDdJ9We0BNkl7tqsSyol0fMRXxNOnZAgolmPu0P
m2zEfwlcAFpmqNflcfjRN7F7VzZ/NIs0SPd6IXaPhazeAbjYPMRMgs7G8nmSl0/C
9eh9BXBT2h/gIFOipTr+zi7kf6O9wT+3yMYNDDkOOn/FnHxLXdlaK9h57Xpu8lfW
IXYuLzHyVQIe7ONT10rdDw0dRsY/ku3ENRPHZcOa/8g0SNxGoFotVLtkMBqi5wJE
PN/mkT06vL4KpQeAhvu2DGxkjkphs3QuIn9H/ZDZl43qXDB4xLjo5W17m22pdYWH
caBXa2UJnArL/slO7uy64XyKdscyPuL7fcwPNQWLR+ngyeZC4khz1YQjagOssBba
blDBNZUoyP1NqdiO6VC4Odob7qWuW4Azit3ITOuH08JIOSEdCZ0prUcTMWvUxJ8l
7AFF4kDg7KpG79RT9LVx/Rb+j1zboNqHrMoEfxzu+4Dm28+1i2trqsUzIURzYX2H
HeGIG4PjT9zg5GwY06MwT/v4Y2f0vpfNYjl63rT2Z50RYfbw5pZZ1xvVxgEH6uS0
8Ek1mCMVUYRJ7OMqfnY/4BA7FHR3yfU2ZqfFK0JOWsfdSMfGDdRzzDxJ08w2x3wZ
yvP4JFYCRVdE2HUIq7+4//6qLMk2FOfbMeNfDkq9Ys5cTCW7V9a1nYFWGDo7P86x
dnSq+wwMSjE6xqBzBGrRM/JsJBi1DMlzhftw44i3nEEC0Y+rF1RHr8x4cAv8mIQt
o7m8smzG4ImrP/2Hh/bzy5rk5qTWnC9F+oYh/U7wb52zkNRxSMyJXKzZ+ekcYq9n
ueXNcWaiyPbtXnYOyOD4KsWI8+4OcVw0IP2TW2aK1R5sR36Uog3GMMLLezkApM1Y
X18VM/KxOeJXaaaM/TwtMkCH5GWRxYH7TwxNQjtI81jl2Hdo2yhirpPczpbilQlE
8wtCeIGCjpGThgTITa0jYtQ4GLgPz0hriMyUuA9KFkeQt1AD+5Lbd+UQrz2UbpCp
/DS8pJsYQH2ya5lICQ56uHBMgEAj0MpvMchTRXptbP8gNo++IJAP3xqeDrN9oq+z
2MVDArCt2Ki09xHCt152q9Cfg0wh9N1OtUBHdfm3YsWg/UKItGTA256XUDUCKSU/
ck35XQW4bAutb12+TQuR2nLV71jK7fILRjOru9NTUbTn7p/dljuivFSsOeWUf6Ea
lbcddIgW4ejFHe8wUdI7tuqIzPWutZ9tjW7UjhikNLPO+dIAn54inq5vf/SE3ink
nj+fVcSVy5A6uOP6+a3XWQlbyojBuG92vhS77IOYXAmfJ0VWgG5M6xYvF+gVvpyi
4dBZgQhUvxxUi1VPh3aM8CL6MVY4karZ3bL+XCiws5tGKKWstaVFLihQ8kfB7yr+
YlqUbtRiLikX5xXC0uuBnenX/PkFsOdmbaOdbJ3X83Ac86uDyTF5f+yvg4lAYi00
EUtvWHV9acKoUx79QIieVrvgHV94P3xSOzoAGFhX1dl/cqdGZHT3W2zjKCbFCDNk
oIlm0TxCawbMxOtvS0LRQzFYxHE76m2FZfrQNJSVl8JGklNpM64Ivq/TyfnE0ZUH
aFtd/EWy/xfOTRk/zPCDR+Htv+DabaKCw2q8Hs/oJF9cEBwd8mpApCIOpCW99aS+
BVMQQ48Gdm55OHbGQgWExK32MFYVcTwJW7iHgbZTPjXVS9fH30tbV3E6qJjLhxOq
zoCm2Ijlm416iG7eSx9KNstJmksTr1Cnm84EnCYDsVq3ML0vKVEKqho0g7lkRKtF
Bxcw9d3zC2hAzgTWgjhvtHM6vvjah1ZjcaPW2DI6Py8I19j7iDX4916owpOY8pb9
RX6m65nhLVqDp2bPFokWz3sZKCJ5V/GPW5JBd+yWLp2UjprkG4rpefrNA77b2y6g
rW1+YUXh71epLnX8bOXO2kYz6SSdivotXtfwmuRQfb2XR9eAgE43F++ttL7gYNxl
qR3DoozNUWTO6XX+R5nx6uWcMFLp68muVpsMrSf2NHZAA7FWSRQRSg4s5v9LSR6D
U2SLoAnigdtC83aM0SeNSj/hYq35NvfxUs/P3mX4u+mcrR14cUtiG0U5MXcsBDVi
UdxL/EjqXCkrhw77uUHBGTrwbtV1V3zOD4BC219f9eEkkJHQm9lAsxZJA19q7Ikz
HEqkxl5FBPMxTY0V5ltd7HKFIvA7IxSKpNqlsSxwv+NmM3gMxsriXCjE5L79144u
fRcqVTMbFq6hWVWx8XDFPmuDsmldFnutSByUiuI6ObahpbeIFHA5euKVH58W0Lqh
ctk7K0mPqVf1oqCtz4KanepmTjpWed2RaMKUROCZArOcAZFoC3oCffa2CNsLrIsm
OyebVOKWbVEJCX2HcVZ95XbxglhbM17M2WvlzHY71vhnd9SrXQuRW7LwMxljsKoC
Xm79zmqxUQYEId+3BQzNPtRbqP2SWZjpW7j/Dk0nzqQCmNoPs91oQiQPfwhpTAVJ
cHvsxzzm+djJZ8NJ3M+4SSn6h1pl7kH4giTwqQ48bZCHVFb4vznAIIgdsPWPUjz/
v7kadwaMBuHRbexqtwYVPEo0/itBEkQQlonZnwW9q9sFm+IjYpXIudEoL6jMRCG2
RNBCGq8G4OJWcgYJ2FgH7ioYDXHGW0biaxs7PdlRutXp7BOeOOzKvy0EdW1FwSv4
Jw5U+NB3SUOc+bK5tkR8FOk1M/24+isbBnMiwSIVkc9zHxLvf9SAW3mqxMcYwZp5
MAvNDalQAh47a1QYlMAL/tden0IjJfPHcOGEDG+ew2hfRfrf9G79Wemtve2oq+L3
Mg5VfYRN4DFWMqd9NiI777DEnO70TZWEfw/zM91UplGPG4epgCS6ouHc0ajAqrn/
kPQgrOp/NUPm73f4X4rjjqCEd44uhWPw/90xVCauopZRQdjQTa0gXWcBC9Myd5/K
37MfK0O0IopMQ+B1JsKNTWyAZ1x63/VGMicysgb3xOFi9vY3OEx/zlJuoFb9GxqD
RMXpsPbAP1ninIhtukhK9oZgSxO9LgsECNpUe5PpGpaDuUejKyO+Im/Wdcl+rr9x
VwdzHH2HIMb11ZtFd/SiPmY0W/zi7WveIsRX0ZOdurVYYz2NSuQp0deh1lAGM5b0
FXyRL5y5dQ4u3nSpC4SC5nVse1KeheDwhyZu2ucKmqQMErM2PRBFmSPCkButZhQo
xN1IZS5e2CXJ2cDShmH6bcff6cP3y4+gqxt8ziJlFTOCuNo0kz+HbmpkqNnlJ4PK
KqZ3wy1Bkv9tHgreD0SlNHEegakJqx9QhZwQpqrwRgsT7AeRQXlnbKaVWB4fCmjo
Mgdr9pTQyUbeFzO41mCuNd/7+f1QGg7jgqD+pAnxpjdUmFHwyfM+LKTFilNVuUui
uOrvfQ1rFiGKYkx5yRSI8m/CGZP1odq8eRUkm02sqRkfVmHJMSrjPAwYKCyUruGd
F39VmswXKzlF1uIF3RhtjC4GGk7+5x4QOVQyQJiZ63kQ2Nl1qAVwKwQkiIR6z4Vw
5VJC3vqZqNnsq+bpFs23hilVicmvV+1U9g4CxoIFeT1PMlpivJl9Do2GBgA7Ynjv
iz5SOommvIfOlCvUYWAmk47VpQCqoPE/TXkqLMtCPnP94KuSUUXTKYSQWqbT7ej0
eIqOJYCKY5Nwg4idwAeDt1ffY7jlJ1ddi9sx9TORrv6pmWSweP8exnQ5K5O4odwb
rzLq5F3MZyAV/HdKr+lOBbscuFgweCtjeaiF0vz2u+VtbboUONFoSSu6JAeLRpwa
88m7Ed158JwoD8N+f46yk68MNckfl+tvRuZbgocsFFf7Gv1JfoiKOQ+qGmUIE71a
Ov3ULVkxwXRlxv1WB44BMLenMSolpmJ+G8WxhoypecYF/zLLpwM7+6Ahcb8Ddrz7
EscgTnu93mhFoTYmkiK89M6tZD/Jwvazd/i7lP5tUJOr4ncf42hsr0WgjO8cDfdw
obg0jIewRESGxlvfep2If0XqGgGlb6CdZ07DaaLohGpQuSud6FGWwxOolkoLI5YV
pMtmc5U9V/MvPUgAr22hMnNy/50IISyqySO8ticG5s7u/alLB+37zj6GD2etMgzk
JPTCQ8EXGPVqeGKzOOB8pPDo61jzZn9a3l4sBzsBdlmJ7ClMBj1FLNw5eKFDo9Hn
Q5IkPKALs4cexEgJNE85SqkpxYd3oTlY401OBO4LZ5Y1RiBUFHo2BlolR1iOsrsL
iwgHc6SO1oYU+nNECqRfulFnzdwmfoDiJj2w6WPpzdFuNXc5ScLkFwr1xL3lf+Q3
yt36lOt6kC9iVNtgl3nijBZ9w9lkBB26TM+juPzYHBkomq79b6fFqMaFO0ccnIJ4
RDyfNJPzLhb34l30NeoxiEecRfU9Uwx/T6wc8M/A4CkWRwfjGR1CSykxWasR/gKd
i+5SFk6skD8TAihaHwNevKSfDIbg4vBMEcuGYiNyhznxOHjMSTteclK4DtWT4XHS
1ZChsXxlxQ9NSOB0pqtnCyqmplDENaSjeGswqxJMaw6kzFJHxdgakuUBmTxRSKYP
+N1Qx7idSshKD2c4pGtArhMWEdSLKWSnhNlgieU8aRv1HsPCHI19CK/Ul8mZk2lS
KFCHTZvMUHyv+608Jrb5cEr7mptD671ZX8ny4Vx+Y4Oo15HMQwXUSIDIGffi+Uwt
LX4rVOVwHQx6WkMbjH6yeKf6bbrYzCNR4RSiAIDQyhOWsrZ8Nw+9JHaAZreNLIis
VNRE2MsL3dwyYSKqJQNEXDzsXdZyAeLyl4+Y5WmTGOqlQoPPOT3rKZODzt/OKeem
gGaSKgFzle6T9myevwdFDqzUYoTUsxaH7JHlT/8WRy6VZ6yNLXIibFWydaJ/rpo3
DLcoTKR0EhfzKXFpvvsQ0U1vVYKs13f+Q6OGyIqSgqJ+isZ7r7+uOseDiHdSV5gn
dxjOK6XvUDCceMxSWXhXorNaKR5sJruFQWMsM9u51K80eUPLkdhk4LsMIUZLDKPG
jBxbJSUS7NkVjAIyUE2x5vURjBuo5fERyII8E0ElMnbriUfd//69CdoxZoGrBmr5
jRgiO3IzX1kQwPZgjCeOM/xUzkK8Nshi0etovDnxgsGXhzsosVtoZ/HhjUu1Tj68
S9kBuTTwYyHOlWo2TX/oSoWsXVb7Klt6tzFKZ//lIe+huvCRSOzcJOeV3i0sg25y
8bDb8VcvBLk2tPVb2r4kc7bE0nn8e/9BIKiWqMcwLy+8PrMiSKCeUHh1iqD7fEr/
ep5eZUbZneICEsdJ6ZLDixDWP0FkPKHJ45TLmCbtb6ys92mc+a5BNmW8r6kF24mK
CTgHS0tz80wh4M+CXLtO5obxZg56kX4dYOdEy22g2vb9dtHawVYyCdxD/mo2eqMF
VVPHLVN7uk9iu6w0gzkNd422aP4S4gy4gQ2cBFnTCvMCgmKR+QaqLorW0ScgfmW6
ZbqTcAaueAwXN9K72cB0fXXRkLSxFC/9QecFl1arhwbACtSL3tSfxbrizTF1z4IO
mSqytUOvGEkNQpUftY2t/XB5NTdzQqPyGAssKTNSCm9LvwtMQgxprXdTzROEZMX0
40WZrslLKDXntGDta3WGpEnhecHYEttVQvVp+rqRHmo=
`protect END_PROTECTED
