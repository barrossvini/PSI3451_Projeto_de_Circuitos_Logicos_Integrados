`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+j9LDk8ctli1uGXJmVTxR1GlxQ0AbrYDE+K1nhXAHtM8prnj5ZLhMmhUAnNwE9sV
NZweIgcXU9Z6Tl0MvxOf3TXhq1gy7wBINB5VvQVlXIFMIuCce8GPi1SU3gT/zofU
RDrjmuhtRL7Ss/p80uuQLOLMdHBHIyVZipDNJ8iDKVoa1hliwddUo0MpAVSiHGCi
`protect END_PROTECTED
