`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mjtzkvn71DKP2gQte5jaDzVAhX0BGi5GH+eTj+lqtQ9Sb1t+HYPlXroa2Ze8C0z7
f0CsXKE7xnqaTuaz1k1IWVSYtIi8qVeXEDvGSoZbljynz1KPMdGNbYbGDpBYMICY
3j+duM8R8yXc+OkXE2ji6jvtdUdbfWW+m5fDY7cNL6ppALU/YJNUVkqGTFl9oPJ0
hfQteV04WiAHLs0K4JvkUKidOOO/P/N4ENZ7Lite4JK72PN6ZAsaDMBy7vOa7RCa
GQj3MyTBm7FtdPa9dG2CO8BrBF2hL22gd4X4DGU4SjbFq95YUuf4pjTPrEg2RvHn
PV+a6JccyQtAASnbS92zTW6Hdd7v86t1oPhA3OaV4VIUKktfp7fwmOEkf2z9Nc4/
Y9q+3QfA7J9mR7kOBgLWZ5RfKbO66PAvhk+ukqEWZ2/4xL2skJppgKmlyEQf89sa
mbIkCVk9LfmXuLp2668Y+g0xImXAgFGfdfy7HPFKpjSx7jZantr4gu4mvp2FOKRc
q8R5uP8fKNTYNLAq6+zS5eKlxl6z7KyBNz2+/t7xQmg=
`protect END_PROTECTED
