`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3MyFHyKwUcmjFqHfPGw6TO8PPQQ/QlzniFS/loy78ZLhEe8jRBP62hBVjLsLsQef
Rj+ODbIN86uuJdvGF83K2TEKQLzvFTzqtpsRI5N5HAN2gCGDh4GuPndkdLxjAGiC
OROcdMQANZCIa2z4McsbvSi7kMciwFVj2Bs/N9JC7NmOpCvEc4r7qpP8aaqjCkkf
2zmRW2OVnD10wMXLi47DwR0CWKQ0yQUlqNJyIaflW7cazsthA1teecszvIzMprQM
iwvutWbz61pWKdyC75IAawy5X3rFJJq2WOmy8t+gUT8pKEA/ZbhBLwkvJxp4/CLr
QKCFjAeNZ4KUEUcPzv1RM8Y5A9x9E/PvGWd//rnDclB7f3DcVLDKX8f++OxV+VZv
2VXaJEQZT22AZIYZbl5dJhR3JA63dlw6/e8SL23csiXZorqUqe7XuX1MkxzYh1Tb
hLDmhh6y/oisXyPIbbCtNFqmzBgDQev5NbA+FnYEHoy3kv6aF/uOq7RP/ZVMxWa7
CYphU3hAp+3Qd6irSEHADOl97MXXrfkoQ7ReTVpDHiBF7dLyhuncJYQnIMGcBlLX
sacDSI7IwrbcjP2y1ISEm8p4GrzuyOGPC6iasZ8xAyHIPo0tLheZCA93foF6wuQc
unuUsTrSF8btS/OAmVRgxuNqR79aKasFzUiUciF0bjzX7+ZMavoCcAeuggzIDc5L
dz9x/TdHj0aDGIfw481Dkjmi0XFTyq5zgYFLGW31mCnPV/yJkD8nGY8hcy9C7wIF
cqeu+7VhueXTqP30LrUhNl9IyEtnEgsDFjxMHP0/cWOgNGAXEPmdKtlI0GaMTq2O
3VNSSBOYvCf/YpjGR0ygviLJ1BVQnGcYEnAvkyzK8VeUH0gWEsyLO74sSK6g68+L
24h5+A1XGrxmBw13sYPX7dSfwiurUkCO2vSdMx1Jw8M=
`protect END_PROTECTED
