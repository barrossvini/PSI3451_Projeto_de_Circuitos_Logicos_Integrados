`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A7bzUu7QwxNF3aKagUHCTiIPtRDSFAC14WULBtsuYG9M8/qu00bN8UqgHteMPju1
3YRGSgnpdj6wJ61UjuGCSjq+CqyM9Nbvm/M0u34cT7TV98O1xQQ68sYnAnZTJy0p
awoKPeDGPCSsT9gvi+XzbWrGrXiHx0Iou7PnvqoCtFbcanc/wg2LifnfhsXr/+T+
QNpv7/3jHUARBswKfVElvJMIKJMs/xL7EuO70Ptnx43JyJbc5nFx22TgZWJiKMBM
gq4zWb7SBfIPrjNO3Iyz7kk+lemTUD894dB54dwLhuol/9zWWqvU3d4LCmDaYrN5
rryuoqsmHzlDX9PfDB5hi1P1uSah1fbblm+K3az9opHkVcSXtTbN2GuChJtIKkW/
M8zLAZUts4cRD/qeSCbu8EkJfuzuWYswO+FanlH0itlZqSutEDERehTE3N/OXx6x
poL5unTAZRT6J50p3WrfGvw2wPcAPXLw2SExcVr6ZrNAdc7XzuyFaEXCLZSdkrWu
5AVgvMeFdQGkyYKh4a3HkwgfM1MFqkeCaFZMpYSlJBFp+GnH7D2lB5L7L6tJXaAl
+OuxiTPkL9T0oNnb+QefeIsYTSrY5U3yxAnBdqHzPUKAl1F//FAtU1J6XBx4pQiY
/6v2lj0TAVwEubq5+MX9q4g52fF5L4SNsDgs0ELtWx2PGPz7zP/qFU8Ysqai3yAu
VWI2UqRhWenw4HCRJhq7Y4IS+PYHryqH41Kp2Y/HkenrhtrgQgltdqN1sP1i8VXG
wWO/ZwHBjkRcghsbDD7fAA03I7g7UOzIntwfKT7JWn8PvyOUJD0bDwKwVnAkOqmE
`protect END_PROTECTED
