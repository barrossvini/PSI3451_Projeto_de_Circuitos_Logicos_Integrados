`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rIBth2HVfPYPfbsrZxyAybGjTJlVg3ViGFELvxw6wJUYB1d9vDTZt4D0LdVH9n3k
/THpI9SS0mgFwdXYxHdk13OVNi/gWg4R5HG54zQdMQiyOz6HcM46beignYZIq1ZR
u6mjv5G6AzmPkm71FK3dOADEg4iK3Xt2pGs1T6U+/XSqvFuU1BSWqCWqj21M+bzs
j/N27kTipdmIHEWi8kSnwzTYtWxtb/v9lt9G6HNaVg2y7oLb9qPTPKn9GAAjbSl8
8gPH7QruZiWMfhwhfSE27EWZjG2VIsk28oa8DB5xA8bqtNGCVuQQ60fAQvB1LTP8
eHPH7TJmYyMTight9tZJ805o4kPJZpXdkf5ZkoEUKmjcDZvzH9dtRFFo2JmKJYYB
vML8eIxawteWHQ1icszmd4mQ3uLOa46F6U6ISnfLFPCLWDvan/O0p3iEx73qNUSi
Ut4fz7Tuw+VopAKMI87bRuNwycp3lphUEY0tFKAwN7E5ijoubmOcfx5YYSL0sqh7
V9exWOpUlQOnXiHdqQ6RMIHLVQG8DWotMdAfWmdN87x72PGiehLAha5FglQvLKIZ
imu5mEiEnxVN1HKOlyoi3STO/5ACKCF1tostrb8cFTrO3GDpztdH4a8z92+fg8i1
n3zgEKLgslt2LJCl+aVzrFMARogGaIYO9/vusVPR/2bXVmACmiexReUfGeQw3jm6
L/aDbdNMGHk1xHnKFL8Z9lP388uFmIAnWMO6jFpDILpV+56xhyzpyPkT1urMtnjw
gPc9VWWD6JTGCQXs43rZmDbF4iwYn9PA2j2I5VQdjMIb+gyfFfsBhxIzqJx60vNN
dFNM61rjT3A9SpbYp9LJ0DpaP/+Cc0pdSd80rBc5T1xgWzXeUdWcpfQBToOhWwFo
fyFtUDHTZBXeqska7XPXFIna2Cw66oys8NwPpmRCj+p8amEAwibmMelEigvq7Vtm
ugSQnLG4li6NnJ/qqSTXosu+i2xpGJFzwGMK/BBliSiTgwEHx51WCFfV3XksHX3N
F0+IKp1b+C0URWe6vGoezFtXu+tKQH5uRiLVAkEPx+raL3ywzHwxZfR8mF72123T
Mz6nTGoWgDoGT6wZ651gkUPZYP+DBGo0UUEHXNyQ2DmMRVI7JiGZxgRJAaBhXYRt
ehzLTH+bBIVjRRbeXIIGNMXV81Xnn0YcNhWbfBvbN+Lk4zsO5Ki3ozWN/zTb2B6J
56axHvFJyDOxFjkZNy5x2KDrWtjJkzFVPyxafEZB9DISkvUibmhd0W3UGbWJ2cID
ErRmzgpnOc2dbaVoSMNTQ8Ulf4z3fYCNIrXAwpgNf5tkWUYwPZuld2V0x9H/erhv
/gdnfqwV1ZNs20vXksnkRGu7A8ZCzK6Kf2AjXv8G4BExsV/rX+hhSxtbdnu2qXMV
3mqkUa3mwE0xRgGOZR19g/HJ5aC9nPDXYtQdCtAdz/g0iBdUqaMen8yMOSGhlBF7
vsB4ljEio8JTW+61ZVXQXA==
`protect END_PROTECTED
