`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NXMoiO00jK39XV/oOpcrNLBR7JCRtcY3Zp27wtPmF1oDmdrUGcqBS8P31/BF8OTi
4gPBXRcHXI5m9MbJj/uPfB5e9YLfVASR6VPRbAnaPttl9fNCfCxm7fJ6eRptF6Sx
hflolUNbVY/TqQStHcop1qVog9v+BbRCB2rWs7lRwHVT7fBboR8STwVearmFoXAI
pii/FaSY9IdEcLdyrKj38u0gdIPqiRRvOLS2941Szw/GJ/EULcbcY0+00WGU1Ugw
AAQP2k9zR98TlxJFq+ISJdI6L9hCVVwDaM83x8PjLIrTZLv2KTbSMjh9nodx3K9T
dbKKy+r2Nu0yyzNbqpwDcUvz2aXz0FPIhz9xpZAeDzvZvQ0ymgVrmUjhgN2grYJk
ZrQdq5ieIsb+aZxGPAPrTMRzKzIZS3SFBxE85gFgImPc5hmlovUjvPVNb1bcKLrp
XTQGaKelmnfupNbFHxwSn7M9ivCTZj6Qiu7YYwxs66GdJfCAE+ltLWb/QeFFoh7G
AaVN4+IonCRhacPmPyUK/lExnv9P1R55Oic7MM7kfaDRwWcu+AniopNrdqVGzNQD
0u4Jfi1/HCOPMdINwnxPFrdpqwqASknibqzW0zUzcr3MiMpspFOm19oJrLlU+wMu
YWRsVhFsBxR/nObzScWeqWfXnBafyNF0uuxm6p3/QUd+zpAxYsCG5psGQ1uthEgh
/E5oVMqTyz92tvBei3tgMEeDt6ZuTge56s7D3zXOnjZMjTKbssTj/1b/0uu9MDlY
+JfVIJqo+yoO7j9T7ACvK6QUUal9U1ESuTIG3XsX4Ufh6jWDnKEJ0iqig1xZDPS1
Kyj5ZRHr3a/1tZyY9WQaEdQJvCGy0zNmJX8Pjc2tJe7p56SAUV130cflzR3dYj81
8/Dw++6dwFm4o7Uegvi4HHS8DwAtyxHQVu+7d4OeourzT2hMo4oel+4D4vLeqOBS
/0p2BxGAVmiXxGUHI5/YsyTPu0GsJjsbMldzJpN/trdgSqQkrHo58neAe0EHRILn
7XbmFMiEiLNl3MHfo08zL29evRNEJbAou8MQiMkPxvu6J3di0S7fHLwbak1g8o14
AsVwZJ1kb7ix8yEzP8OLrrmoPjNM5WSFKF+vBxbQbMOuo7QvYfO/NZsfMsRLgLPJ
uXId7pRb8QPtuW1VXCvfWQqwqVqndmOYz6UYvRpHQCn9gK5zSMyMHUnhqSboI4vz
UBtfSfpVF0dPNrgOMgPdfQpVgRelfPVsDbe00BNDoUj41SLWTvBMbGgySlfh98A7
CDWPe9TBhtp9BN1YpSoYao2tDX1KlB6v0Qe0asYTGwLkV7/+YTDudUzLVvue3OlD
gktq+rWvTyRg/iuRNmx7xI/kMRCMiX4V7pcamJ0qtkzFy6WAYLDnwLLxZ76yPpbc
sIL+UveGHb/NI6ZppU8PnWprTFRu/mvZH2hWsv9xzp+gJCboo87RbjyRGxih631i
Wjf23P0e2OtOe+cSPvunuF2saLI2wEhAUph41+IeDN73tJ/TKrKN4Vs9B49i2cr0
tSGJ4wa04YeS1smLeDd9daLUECHn+1nuAmG8ReDd2uW/8NZ6t8ByyJCeZZUtX0NR
yQkfRfJqm+wLZXtDJGYQZvrvQdpoHKafzAmwlma3xhLkyMUR/cH+HiP6b/cistxF
vAYUnXjpf4qs3PxiJwoieipvZD8t65FLSKknFDnsUHY1+prUeZkdJC04FplubzOA
OmFGj4IDQGuaUlhjkUVIIZ/jk6TKI0p0DLP53maFXsE=
`protect END_PROTECTED
