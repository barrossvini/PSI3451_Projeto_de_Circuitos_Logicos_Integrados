`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KtGU+ijYGRdbAvXBlnBcKPq4glXMNPPQ1A1PQoaZH+QXyZU+MREi9KbH8il9JIGD
pbLnWu5FDx8+gzki7clkpq+Cm3357apM8Ddi5G24+Hkv2+ZEJqwTB1707AtF5thi
EISHT0/hThnBNqRa5lTg1Trxbk06LTuvpQpE+WGr9uniJZzxdFFFqcDl3Y9l2pGC
XFnFhX3haY9rA4gURWSaaKgIUjiZGNTkpH9137VX5162JkgjS8j44fh8irPU9neh
tAD1z6RsSpOmo/gaeuNkkT5agqLHS9O7l4xmjWKAZF48BTCOZWwLHFUyZsFuJGL0
plfVXjwlISats3U67AepQnVkJXgaqz9veRiAw4uG9t++IlLoaP2lnDqvvHcKHARh
Ywf7+w+PRsAruFn2plR6Z5r5fJ2uq3pKQF6TX+OPlG6PDGZTyJK8DzQMw9iGECkv
kwD4PDSHf4ZTa4V1R+Y+YCxnKblyuBKIFuSWlntgufRFfkyNkLnUwQSGd0ivFlZg
XfpLViQoqIH3BUksfG35E4zyrBQ5fydZ7CUc3Bq3wZvt5YvCa8Qp/StG7piM6WyO
J8j2UbUHW+jQ9x3KnBAJfYHc/wrdvnhMrwa611Ds5z7xyDh+mCwN0mh8ebob3aNr
1VKOOrX+69gNPnL4ychjEXweayeh3TZnCpruT2z45kPTfom/RK+sAubzNYe585y7
jFirrP5ZL46PjOVEROGZtZx/Vvn+rYlMyZaEW1To3DDFXVpRpr304hLRiDS4pYm3
Z11AzpfYF05lOSOyKYh6fosW+SQIAaTfOWbLyyLTlc+yeoiQg+qh45srL72ABKM4
bdhKuzF1xnVVregVpFZOMYSzaSuKNG1p9HLL5FeNFczjibToVDuk0OSMuBhJIJBQ
LExHX5EIWT0oluFGemb1mlfGGhTOE09SKbC2CkzWITVYOkupTkWAKB8INNmPEJTN
+VqKSjhs8WB6BsRmcfjmH0B8ZXV6fhiCarpE6mKT6TfGWCeGIkiKsjV+EbtFUSOP
HD1sq4iUw/TnZhxIDYGR9rXbmtANewQoaHb6b7k5LWQJb1wrhmuEIXMoZoU4QcfQ
dgWrXARU6szTCss9/BugvuFfI+MsauEqPnZzAkgOMaANf4SphrCGD3b6W7XGOvwP
rN99JmY9dmIpBQVUqwuteQ==
`protect END_PROTECTED
