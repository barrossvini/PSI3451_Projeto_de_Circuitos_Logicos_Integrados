`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
esGOX0N2HUSObiSo5ZNlAoQN24PurUc56mt/flnwYYimSbtxqZYXBSKxEYROpwk8
0VMFq30vbgf/6tfDMuRnaaKamkU1i0M4Qe00N9Sa+2Xt688SrGwAFfkvJ1rSbKtg
cs1xSTdndFd5Zo3FOHShprTbTOvjFWF1s0/M1mrkVDq3YDBSxBzbrtmiyrFcnLAl
IarJwFtN+3uaYOf5kA7ztZGqxSUQd/Ih5ffwOGWDSKw5yM7Ne/SMK0yVyZenq6n3
HzMqlPofYsMxH7YeTQVaICJPDJGAzSkTKrZFHGX09YqcDK3IpkPBLImDtHt/ZrKX
dpZwGDJXcCQuo39la5tXtZMIGobQJb5sZTr4ITsB1IXPakWc3R2iGo7dLCXvPm6r
UoZ3//PqURva4lrl2FFKYRMoTrN7xrkh+WOK0TPZVlHpRwSNISsORlVoRpGFt95V
UjL/Jo4w/I0iza6KkYbN59n7jGt7MxPkKmH2kcYfbCEA0bW0SS6CA0n5NrGKy19i
8LB+H6bkHLaSJlJpa9jMrXqPG6I4FzFIqwHMyFNzhdKf5ETCMtGM+sFdmwwtgHI6
TimCMd8HSt1RdOPCMDaXPr4Vuj/7IDEj8n47vkazSsciy6z83pc28C2esuxstW4G
aXYSD7MsQBko5MYkZf4Nzw==
`protect END_PROTECTED
