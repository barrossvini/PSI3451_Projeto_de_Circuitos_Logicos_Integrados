`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MAPCgeOmmzEADjSH63UBQiysawGCA/V4GElCgTgEIflVU983dGTLwps8IxsZgJbj
io1fPJmDcZXzMdb3dzJhjQh42ppHCoB5syQwi6SmvoC3Ot2mreeyYEKFIpXlTr0r
wH84+tA67FZgGGFRo6l3Sg0DPa+VbdqMKz+8NM6WF6GQmaIxmEL6B/LdudfZXO9p
XLRDdG30ptstVup1gaCyTfjpadRk3lJMqUsOqJA/kd0P7S+nNSM4N2eqzVMoLXCL
xKHMMLnt7rUYRPsHN3anGn7ku+Sv7NxkVW5ZIBBNMdXRi+PbmeIwpUawNOP4TnMw
7IaBOen8ry2pW3jKfNpxtyCHZXyuCXgkOqSr+4KV38IM+lkbyylppBjP5yQYa/zr
tEFpn4tep2iux60M4dAOY3a9KRbXLw+Za7UYotLT8xlYSuhzXRUFVBL7mnSorspe
TwD0AnvHEPps3globId7VHhq9juFLx3wgTM0y2cJBPd3Gpe0QwKBeJr6k+De6bJI
gGxoV4kGWgOBCBMFIJMMcQ==
`protect END_PROTECTED
