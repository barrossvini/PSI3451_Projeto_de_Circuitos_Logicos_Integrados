`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UtL6K8cVnVVYtw8jkX+234N1Kp7AGkcwGtxRcVK9pXJbMuM8Ct55N1XrrIZRgBx4
QoT3lkO9myKXG65XJHH25OuzqH4BT75Zv+0wRt8pHg5iVx98NIKED+BwuPl0d0N5
+gNcoNYSpc2AycLSt2G+42RccnEyn7nt6l0nyIagEdvERRh6wEEgHtnvpSV75rLI
RKwWzivtgYpHyV1lKm2cXlHFqN3rgXXG6zWmK5cJc8+RcEbK0ih5ulzLhHwIXelE
KAig9G1A4R2k2CvNm8L/LUWtH0wjdxKgtyrSJ2BB1FvyPI88YapTfpsk/RUi11QX
Tl+TcdqelRozTUHdnJIkrVc1aPqNcY5rnltY19AV8wj8ep0zOPa5hy6KlnzAM8Qn
e6m0ysKbf3E/7bVJuGis0XvQK2yPhCec1FGWraiKzS1+5eKsTy9WJUmSMmrGivDY
ejFEeQuY2GAu6HakvM5kDVf7/bPssdAQ8Uej0sx1ZIW7Hf9Ns9H1Th+1JA9e7+u5
eKEgqZFRnhv+tjSIGuRI60LSM3oNjDyCscpAWJ5tyL4HrKabwtopSiJCZ2fzKdED
TH56Ui1GJv4rHzHPGMIzvtTGo6D1URksOmd+O9OsLzobJegTCd3Q/thXtyLwKxDn
JyRfZJgONIFd9lpCF/w1Lz2FtVjIYsQpn7Tdbr6Z/xMFHJm+VP16exOlvFoq/kwd
ssBTIKGPIep0pMasHD6fZOEs3MfxcsMGDmm+PjoBzDrC/CXCHRUKst1p5X6tap8b
EvxXlzeKdeQZ1xa6KZG8VhQFso8NCoo30bqSTOpY32dJ6Xt3QyKx8HPsyzCGqjh0
I7h2uTG20rRGOWcuEtXcm/fTFlZCzEfEcHCCvbArew3+5v0mm3+Wsbjqijtr1CZZ
5JW92HKnHrH2tad4PJEh3ohY/B3Rd7KUCOasQCav99KDvsdX7Ps6KptxxA5lNsg2
Z46i1eMIJ+EDSbe69xddJdQMlUN3vcNLrT2V0SkVXwIz1p8XW+a+CcKEH5tfbyXQ
ftA2rgpmCPL0GO57hkTH4jiOzAqCC32pCtLBq5kqiYYh0kXyE7csFdosrzMgNEIS
i2Y9lZe9Bc5uuWrx2USYRR9lsRdI8MQB0kDZjAL6WS1qbYfkXZzKlmI7AeaPiIvK
2BuWdRKzeUZ2VOV0HLhUVQYIH+/vZ/NIzoq6ITqX6hwaXHMNW/X44bgrKIQCD1Uy
eQxYo59SL3w0/+Tak23xYTND7c2KGxjevw493eteAFrJRELd9fLXJ5T+bQY5niAF
xspy87Sm0vrvlworYIaE12yV0KsWtWSrKHR8PDcYPdO5/dgGUyu6tJ+9Zc1/ziS+
msRT8hXfjJPoe1CbYmW0c0tfuZQqYTA+0qiKKC58eA/95DTbs5QI5niAvPOj3DDW
kpCnI1aw+7vHUFUVvZdmU//p7sho8mhtTuE6GkKB+m79fNBtuaUF7vO4NQ98bLpe
m541OANxXyJTdrNaEmmOEnO0mWNBP/69uZj69od+0upKYbGI80Z90/VLH4wHk3AS
bvvTUzApJkzmfze37/IhhkR3kl20fs+4lP+KdmnIr7QuJnAC2n/8FjRLptLAM30e
/83yWxVkfpCTLm7fqFZL1DBprZAnYwJ00tGgri4KacUvl/H/KDtZNKccy72KqGex
2PETFtCvxFgPlSZnJgLzeL5bptF3MeeZlcNiDtz7Mo4k3CmICJwdXAHnj5nwECBJ
A+u9waIZMUZNjknChuoSUhSCfxnZJQzGkIyWcaKG0bi5WUX11Bx4PbupjoD97g2n
bcg50BBqnMmT3t2zmLcRaH9VAi/t+YV4uTH/DrYMu1EmG/7aXsR5Vw+b6nGnlZg1
nhzW8ttlWqwgxh7fVK3BQtOZOwqZ4V078vQ+2eJLihYpc6XkbfHibLbdmbfbe7oV
FLoDhZAgkOpTImJjDUyGiAzJ9Qk74Q43/hp9Fype3mzfV1OOyDenK4oNv4mH43DW
NysdKmlu0/MIRKsKbQLVmYliXBE87wvwJ9/IcQL8KWkyPhWB5OyFfJoPl1rtk4DI
IRGzhexbxv0xcQgShPAprisu8ljnwwPOBiXcZ/hqhSDNbCaq6VDIYE3xHdrgXXu4
/DrZxn6XET+45K+spqke1QBKkguzEqD8wdablvQOifpWZ9VxUf2ZmnZXIIZl13lO
lJZLwNORISY13tKdURsuNxk1cLpi0PxsWioz8LrTfXHouHT1BUytNBEBMyMxZPMW
9HdKaSmeZYmlxFuHj+ex5q4hpR+lDNC9lM4uMwOOGi1f4ZzSwPLswOr/Tgh4dVn+
VaJ0+TjPP9Fp11HLuX9SeaJMAQC638tx3DSqAOQEFJzSsqJMMzigaCXXomn6Gf2z
jI4VXuIdCA3rvu3z+MN4ARVUwDMQNJ+igYItWjt4ch+S9S8cRzp+J99Qtb9vg+eq
hDkHBv1XvsnAxsSSbCCo7J3xR7tBAG0CThPaVlXP4xKQdy1ttOHDZaB5hqN6p6QP
YXdEihbgv9Qledx4LuMVOV4zhQc8rc+beNHLyDMTOsT6F/8H3a6aUCrzJeJ+kAt6
TzGaFlO5BT0SSwBL+up/HP5DKzZsSOK05Dpfb8UjUzHUYwizJDHiDp2AQkxmso9L
mjiNPzTwGSEHoSDb221Sp9BdR6c+c8N+1+Fd2q2JHMkyUUeVUbSkOrgaWczyYNOI
bsAbc9dFM3s2+LVkpmLqJQQqqazyvH/Wxp1Nbm2BQZZclP1BC7ubAKFYOsDij4tM
3vD35vAiBeP88hdgR58IXsb6mL/4sX8teCIJXI9D7LT6o55x5JUhsNzCoSKW3V+N
2HREDmDfvveK5d6MtJ33hUnb/zJK353IFt9No8AvV13t/7dnITlqX5KcTArGtT5v
HRBWR/Kec3OT7mKeNHKzJlmqakae/TJdDfpOvJoZok82hVu0J1mC3Xj2jtRfNhMR
tqVGNlndzNjCaufNF1pziJSwYKARBSsgpJjN0ZgaVR/3YBi+VQPIaY/6pXBM1kXh
DT51tOWAlkxsjYxvGvAOsit8kkWqQUynUoKueNI/cTkypdHJ9os9dCEjafX8mnOK
7JOCVtioQSz/4z16oMhGqin2ka0ZOM7ktKyQ7XAui5wM6xDgZx/1CdqL4SMUspM0
V9IqdHTNixI8WOg4rN9h0VeLvQ97sCfXVJtFs05Uds1bhGD11UdkAwsRk3OVuleu
m/xkb4ukZvWHqlqHVH2zXRXkV9mz/UdrF6eO8vxozM28IvM6kmDrtOvCjXFZxv7E
w92d/EqLWfsaZxf8rUlcgh6Z+DwILN4xsIt8sYCOxWOEXvykDPbJ0J0buOvTQ3gk
RohcvwCBTGeG7sAr/uXoI0WIYueLGXBI9MqPzZyPeHbi7vyUtd1ygvh8HrDbNxDA
fAQX1bsLd/t1Ilb5xH9KLvQZMDQFpMqurNZejzrWUM+iFq1S+7eHeMQ748aQgjcL
v1HtSTHtmklPTV7457fxzobZxleAgFTNS52nRK5Sz50YhvWB2gRB5IjhX7C6cFhA
8j1xG7KtS16YDg8cq3Cl8B358rKvMCZkQAKI1V+7kVDMEZhjDvIoPWRpaANuLJsr
PYVt+nw/OYgS6n7oCYJ1FBee8TgG/O+ceWPaFuwMfhLBsrJxSmZkd9x1FNC5UzEC
Y5XF1/b1HSbKZ7T4BGS5OUo1NB96gNZ5G1zMaG0gnoXL35CrJU9FMqAvKvCG8Bp6
bDQQ52oL7k1S6AqL5VS9UYpVp132InSGV5JvFVIaflSNumFzCsh50pWmXJAWS8Tj
NsdlDATnJwARe3cJN63B2VyveaNXMX7ZcqNkUpXU8iepXrFawskUwuCZq71x2Ewd
eHvTR4nT0H5yXo2xHz6Mn9CFBYvQ20U5YtFpFTsJ6iYkdqARl5KiylQQJRz8vcf1
brhqG2XqsHwUmYlW8OLvIPYc847DR04zGFAIQUuen4DHKIbyKC0u+1/wMyKrtuCy
+zg6lKtZ6/ycFbnJ5G7hFwwJAMD0WTl/4UZrP0H3OxWZaODBMbVriwk1T4H4fkK9
Vlm7xlg9q367l7IlMO4rSbjyIYkIveTlTzZvExQVcPDK7T9S98iiN70+Pjhdj2BI
0Sj2F1KkRyCYIatadmRJqkRGL/JTuf40wiJngkjSxdm0f1gt9io0a1WLesldZujy
cPQk+5N4DBpnLQ6T148KRaw8gn5Ez3Q1bd2/MuJ69UZkn4cKzC8PfuAJ3WbZujc6
rMI/sbfEPz3hkaIkNILkqF9XF89K5iI6Uw+6Om8QBauVp9FWlt5qma8K8Zh0A88D
pF0OIYdcavYjsyjAC9d2mEFq19O/jlkGorbktTY0ed88zBF9j0JmXjFZgojur/yo
m+K3V4o0Cs8aQf+DXWCMMi6LFECMisvMEqA0qIhVI1TsOCDWjZu3izgzXxgm18Tr
qJ3dCYiembSqfCQuCragpQUUu/o0sVdU6q3u4PjG05bRRVdhWZuzB7YrYIYq8StS
wSQ9gySYhUkYAn32Jh9dvr4uPdJcieMJX4AClxNd2ZGYr/fQOqBFUfZGbPsb1kTx
fkb1PkvkT9+syZYdBNGgtU7K17jUzkmoI0eD3VspFfa2TohnkC+lvtF99cmra97d
umQ21eQRF58m9NvkKrhBvTsyKIgz3XPugdExg8lXlg0AvnpqT2JsWjqHYJv3UOpr
4ZQvqQnFWinQ4LmyT9TXPXys44Ek+fqn3yMTHCmEa4Aaki6/sNQlrxTUWVqhsn6K
KRIxQaYFFWcv2OL2zwmowbBHsjS2HqRmPv5c7iCNTx999TCyG3yQ1f0UFg9aL3EW
wNVTcU0LuTVOPWsZp0LV7a1xB1xAsk/q5XTILxxMwKZ5r7VhROwss6qUyfEu05IS
woHbgb71aW73XsLnBU/1HO/l65KOyRVmGyoC73LV125dITYIseVGWF5vBjGMYk3t
WpLho6OFSxHs+lt5fo3UB8JA4aUWyNsUpYQ1M8RWb8czDIK8HR1HWF25OLgfMx9I
q/m5ceiXkkfNWkVtaHBEhzD+XnOaqLZN90mo7/AAIiZmDt5jGurizw7lJPaOSBCU
K3F7LOuFm6HNF3GZFwKQGMh0OVHYfhaKLtVG/jALyGMGMpLKYNwjQum58ouPSC2U
DCu+FwbUN+3ZrixMfiT0FsgHlZ1/5Hnme9jbMMOBRGBehdvrL3hcu05FrhK4j8C2
duRtTSpuuWP/QXuN/x5bOIvrfVxywoTqUBtwHSfdx+ZcAoPQW/Cf1NTi1ek7CWgr
yhhim04x4gk64inmVU1pCPg2xrbBXP6Ny2/hukZ7Ou73EBDQoJxFoxt6Zqcv3z9U
iJ9l5TzKMij89z2N9TmGyG5453fkHIwkA4qD6RV+VqDFOTJ2Oo6qC8tEvJIH5UYM
dRq0bFoU5kEOc2vucJuUyDTfq1Yu39i4SfPG8XBX5uwzaFxMrFtdJavS3OBIttNI
X5E3vU7PW+FkZzv61z50M9wSI0CDSoazk2oBu0tblNj8FNjcU8r3uj192j2vAHgW
BN7OchSkixk//wNe8/KYaqSziM/2T7uDC2YtkKIurO+x3oXxmN8DHo+mcvYNPUyh
3J0Y2i6KwindhAZU2jgk7Zx9bUr7P/2fav3Gk9aQ2fovCcD/B8NkT+v3YDEvSxHV
7xLu68WUyv3Ut4HzQFW5Ntd90L1Ds3rXK8+OvSyVqtcnaQHWxyYl2z3/LHLNd4Gz
QkrLY36va+nW8GPpImSWlm5qw52R0bqFN/8hGNe9Md97DrgSFwOOjzpFK9oWUwL/
qHJ8VdqZn/5TQN4p4DV8aovMXVBDtZJmVAbmw/wwqtlC65euxPPwaJwj3t2LgVpm
cDV1jsQOkDmwvDSLKL/t5E07aJ52pvIVex9ZJdtOgaggcbK0UuBgoDO7JbAowKMC
1bNMnK2K+pvWib8cSDPdUX3EaJWkymKZFJJaGpGbY8hDSnadZ+E+ILNaJL+GnNMk
wv+K3yco3lxFmwnhEx+VmshM1WhB6XO50Pz5cEbMM5IUVRZw/goLAamYuizPTbuC
lxuJ6/gecKzFqlauq6FfnlNzqpwElpQwQ5sNOlbioxneAPOWlW0VmLerN2qp9lB3
TYwVy/NRfT5GoQrAj9qDKgHXxjOnKdEK2uI94CA5OrtBfKiaDwcD3z9xuszF11vp
eZAv21ahiySMDduuX3Ewxp0pz8tA3wVvCUq4dQutRWMoFtI0sSeE6G9FFH452eHn
ZpBpvtSJl4/T5OFkYAi7rqE7QBGoh7pSjN53Z2gbmmIbDx99JzR4D3yVWL8MG8Yz
W3BRvotvQmPIYe1H87qQkD6kp+qzY4wKvDli33YEqcOIYoKdqPCH5tjKPhQEXDby
ALksnlT7ds7Psjud18W2T7kngWTrQJKLOyrIhVtdXKHPOMh8WA+17Zm6iEG05Ftn
EjB8kwr3izpd4NBjOsCAseNGGsyjMYImjxNYjLiIvCxTFgwJypuAef1D/CZAUpZl
V3wWwWJYcJiWzH0+WvYxoSbgQrZfbu5V5flwyux1RacZHmnbHTulJeROoOgC9ztW
ZMSP7XSi9n/aGIQEypILcc0hnGeEiA6fwNUDBSvUHdlOVWC6K2p8TK4cTQoCielW
KdwW2CEbjFXlPWR/10qU9mAKINWdm7ym10iY+BndlwbtXRjKy52MDNkoMnmcnXkm
f7uo1rT6u5FDEz+1owvPWAQSPfWkb8NpBdma4soTgvUU920ZnKZy/mLSNlIio+2k
Pp7cf7wLOufChXjKAJElw3UkUnU5YKYSNqmIUl7ERQZF/B8r6wiT5/oEFLTMOP2M
pQjBJd3trKdBwrnvkrefY/JftQXvbO4BAdXCJ0Re/yjU+aqFb3sIEkS7rDsJpIiS
gpvCWpWx4ELWVAbfypSON/MYbzbk0K7bLp3skk/gSIhrbYV/8UWZGbYAYtpD+MhS
Cb/+cy1RqjKVTQW2BysSzLFx0S3rmS2dp8bGlxahlbSFwRjjPD1jMtTHNkkaxRXU
5rGDvZANr1RmUvJBosfJKGJfCx7cay+27Q1zNPLKXrOLIKJtC4WPYceNY4rSpB1P
0TsX5jq+ao4ff9Y4AB++gZEZypTaWn4xFIUaEXtGKkY6Z/kE54O6vHn+RzsManXf
X4LbX5d9bTpsv9bwa0G2qfLbIGg/WmS7EGslsgoZHEfSBtH9VZhka69xtPx5GkGA
1WkCZGpFzZlDcCq6gCKxQZ5QT+KoVFpWIE/chVnHtIvpatiyta1+fApnjT1RtDF5
fx9p+7yN8MCKXo1C209D63KAhZ7MDL46ROpSO7faX+4u02NNxO97JcuEHR46DX5m
aymC4XE/V2v7cCT1AuhBAtEL2JkcJRFXb41IQN01rUN15lmMKSH4OHfc8ckAoVkq
aGBGjGLk/zXCc+PVocLeJa4NZLaOMO96kCLbL+QOdLWj4NCTh5ireQbLx+pvGcrk
3pdJl4rfLoaCi+C0pWihXozCyYpeA0N/dGy6qgAhzCX726rd0hMv1HEi3kQZAgbJ
MWOwBiw9GhOFQzx7O0BPLilztvtz3xAzLCmoedUGC11tMVHPMZ3bTlC4ojmFwpif
A+0TrzaCi5V4AnE/WP3OarjCeflvo9M6jXnki76SOMFJS6tcEg6DMOn8GrlvvtbH
iNi0v2BBNOLdUj8ZVuiShgFc4OApNojQwEYWxu8KPjN7LyHMNKN9wh/0Yz2rmTdi
KN1oAkq68w2cr//PcW223Whn0UcqyckE71DgjSdRK67fzDngYCmgI5NasXro8FI3
Mj+iRB0loJrHWWp4S/SB7u09zYuN3SV0SZNz9dt7NzaafH7A0XLcScXd2dEtI5Lr
u5/SJFOQxEu8Y+Cz8kJDPiYaesVSv1S+37dLPcXii6VqWUKiQ0uXzDKnmYHRals4
iY/3N1988lJ6cKo8Mgs01B62RJHXY3gE+snMC6IhCTo5s21EO0rajgeY0p/gYIRB
k717ibGF/heO57UuScdb2btcGVURGDd0I+JFkQuzQhLJx5ThRRHaaJiVxAu9GYnB
S+sQhg3gRvFAL/uitl+R0f3ipZKbEy5dKDvIN3JzO1HuHyahTZyeRqf1nx7V56ad
MgiezlkS4R4yQ4hYJvSQMrqbnWeePfZ39YngL8JYJBWzdVt6fviirIeWTm8u6f5z
Q4bUgSsHrpYuO0dsS0eBe2QS7pIfLw8myOMamIC1nZ8t5Hc2Bna5eVWUgcIMiZz3
cRtdBn1gc+vE1MVe17x1h0ALNyGB1nFLgcMGI5bSTlS7/YtcTXcAJXmF29X4BaPB
1xSVY3okCXgM9L7Y6JFtPauYC6Kw8PZyR514FEU1CDaJif+vx+ghXDsZSbgItWa+
XkZ9JlfsiYK847Z1uaEo4nmWD1eJPIdVwqvsdCf3LVYQZVy7P9+LVcTXER/PKuqc
I1FFn5Zge0cE7JRIFgv1uL5CdMG64f0SNISG7Ps89MNAQO8d6jYgGkgdzfQzvLpn
SzcDpToGPzdR3ENTnr8U7101wFDanQemm08mX6X2LdmCLPhWruo1Jg7aRVzz+HFO
o/PogxHgfF4oJIgYGimAUFQ/CwNIYHJam4ZcYtMk9UJebJt/edsRSvh15lapy0FA
nenX2Ew8ofOhFKoOba0e5rpZXmOdpHBOMQs2XHXrTYCbErVJcffeLPtzqCM3NpPj
iwtWtpJTj1CWyhhcpX8Wq7IsG8s9zd4ce+5WEgtpa9lHIc/jruJ3+5C617zbl86v
wl86hfBuwpPhe/61QdOcTe0Utvm9tDx2FtIanYaMu6NzG60f9VytyY9LeUqZ5agb
KgE+302BRKoRLQYamfTX9IildcNE0qY5rpuNR5YblwFTZLo3Kvh++vWwtlFFNUmy
l3fVdbkSQJ4ZC24nQmjOwM87pyzb4oMNCKGQJX5W1s2WCzsWKFHk8oQwhFALT/hC
fi58+i3Ry89VUbYBkn6nbpEGI0viF6wF8B/SObRRRzEJxJBCKNggP0VrBaqglE5R
QEycA7BJWh3RE8jReG38UZug6KOrEPvcEP+LrDBip/SMG/AiaFWQ8QrFE9htjZ1C
k9jKmFqfCydXGRj4t+pkB93UDNXEmeJngJDZpIGb4HnWt/P1hKV4whzmCuCqwo7S
01Xhf9U+RaDZxYlV4b29f+f4wHgmIppr+ShSTVO45YKFDQ71O7Q7acsedffxA85P
NVZzT42KZm6VB+RJzBjQn8XnvWzXSdpzkKMwhi2XXyfKV76vcQvS1D8gOdg37m80
GYvyWck2Or98gLz5IkxYUKTEvS/lingtsdwX0Fj3FR5H92rlEy/j3mPM3nKzvmui
Nm8vN/9l1LOi8gjG4kFZer1LIabBrcU8lF1nvf8IXeuJNWramM5OEiKPl3lUqWAK
y2iLZ0jHl5WfmsSWpo8Mdh/NBfeudU3vMTNH/MtI3P2iDW2RUD+eSvRjKKY/eU9g
Hj0e2EvZXB+PxbfXfkw3N0OOG4SKpZQoiX9Ol0eeYHgGmRW/dX11UTRnpvsh0khj
SsfPVG8QFSXTp9WCLjCVqYO0/mRCrSXszCAXEgUNQxnTOtkFUDRHUOKoejMxunwG
3NGZZz5g8nrFV4EHqugagKnJUX8SEx24wUMNkWHrBqRGfGu0yZzHLtmL438JpB3w
gMzZumTaXETgtsxGNDcSCid81LwLrs4iqlhJEXcjUm+2ncuT54nQD6sqCdbSkfwL
sgNdGtxzq0eGaiQIVgwg7zh2pdQ2dRFulCol3VLhcJPJV+RrLiMFQuotavvjXy33
3g2OqMyJC2toYIdfC3eglOwRiybJPnXye98ML+ogLULVt6fDXPWNwcCErB2JhFiH
d2ZAcRhebfvIza3e9OUgD/0NEm4auWKnqcINkv02i3SiAt6j7glG/LSMpKd4wU6b
VNAD1GI4IaSEZl3UzLUTELibEJ25GQ9Ywt9RMdPMnACwncFnSmnrH4hLOqAcHkdN
+XAc1onOc3t65VJzZMTzuUhSbPiG4Zd0edVsN8qtnlpZbuTrhNjJj7jlth5Nut2q
TImdYGEwdNFOmV1wLPG3E9s1YYT78mNYSwgT1fqxMCkSxi32HRwNF/2t1R2X8lh9
g9ZmethKlWnUh2KYUujYLg2nSE7XTqi2/XbatkQFynejA7/I95/Jm0mzW+MaTPIr
BxTj1lpoQKzS1gzet+NOcUJX9crgwNuIwyD1dyM8l1rI8WdG+y5+wUeed5ljCpxp
4Foent44WgSaS+umVriUOY14lXMWhyZAf5GNqCHYTK029AjFPDxurrPZSWkqkzV0
IG5DOE98W8x91fN1s2zltyk7b4lq1z6eFt//JliOqUlZvxcJ2taQht7Vp9bjAr4L
BRhQ1Gqkmg1NnrKPudxYZvqISibw7mPN3gqEUcFUisiEsjnKpSY4JsU40odh1Myo
nHQmWGLCk/R+RRUq0BdYNPN8DoJIqoeApMAvkDU4drCQHfdG/Fzkm8gmUYl67bzZ
Tsa9Hmm1LjBtCabLyS/N/WR7/aEBp5mVyORR6JzNhBQRLRHnl+ZSmV1Q5NVN8z/r
ncRE51Ok3fdAOD+9/nkcJo/cc9WQ9V0bMOyVkzluuCv8Rfw4IM03Rzq3nJjfCFKU
ZjS192yZa/n3SIfCGnn8dM3gGhn8tjUIW/uxOlu8V/qxhEP4K9A4mFroHPPAO3g2
E2NToa1BkgeOsVdwUGeziDedpLBw6l+YHlM/yUmKXlpxkJ7OaGvd/MKyF2j3XrXs
lBMI/25E6MRt78FYHaDk5Ai1hMpHjou2RH+/PtmEKEDVrRd4OSbOjs9aOrCeuC8O
9YpqPkT/YfTv5MHNSVyB5OB7yZK+cvhQrWSVPxrIVCTzmvhz92XW+LdfSKJjyFOX
C058CiE6mjlKJbeUZxjGNOT2wVakdpiy4gDE46v0unnvZAxK9F/srZ+7jqevmj6j
`protect END_PROTECTED
