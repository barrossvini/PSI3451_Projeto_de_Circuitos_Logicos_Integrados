`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XgUJ/3vNQR1fDK332QKdaeNEnfzaaAcLwD8ccLmxbQIZWTJ7n3u0/UScfdORdn/Y
QN0pr9H80NTZdn8QLk/lOqgTTRx6g+k/ISua2jqe4HXaWrTIWGILUOsrToRmqYkx
04zCj7F273JyuDUnkRPnO1Yp/yjI8Z+E2SicdEoiAGbViWnkbubpRpKCwSAn5IvJ
vYCgcH9AKaMXvQVOqdSwTXhl/R6zL5xifjFQihW4Sb/LFW6tmKHcUvtv31c4kodG
YDAUfEG6A5IsyBCADyruDcxitVVixN62P3tQRip7gSfOsvAvMvilclynaUpcZKc8
EDgv49Kgfv3aat3MyARitaCRjqfEp1Zt9NziVILYGsyrDT1Y+sfRihF3/Tw2mfUO
m+RUIgXuqt7MvSbUSziMOtWVX73oqA+E4B/JN3rI3ny+PIdDsypMlkzOMCZgTmQa
Qd1ncFRLI72BzBb//bNwM00kDYZc9FS+Ojp2stHEtbLxXwgUvFY7XO8JIMBxscAq
tPm9Wih6eTaecGbbvd2KARBbSu32srUvuX/IOXjD9TBMqHOKVYqDg+06W5j1cTXF
cA5z5CPVuRmr3dhd0VtZC/554IgQMHELtD+z7mh2d2cF0J85QUiFmRqrLrZWfKv+
vnpN/1t/PxSgjwEEhNb8fFs73LW4m0PGMOjxZv2s6g35LOnJM4pQi8HxdoxM5f8Y
VdrxNGEBxTgTVrYkjdVMrHDayUuX3q+yqTVRCjc6mgPCoR6wnuw0JTSWoXBlxSr7
8jMpuMlbQbS8HF5rTzvtYVNsqFnkBJxdBZaORZuPmL6ch/K4+F/LKRzouxQFJIBL
j4bUrHSipTdh9xfGDTCMOjhqc66RsynH30SNf9oQKPKI7U+vwdOTZs5ooOqoEW+R
9Obl2xkPERUq7sZ20lnhoocnhK8EiPtBlS8GA6dOP73U0lr0fw+4XOl74zXd0zJr
gGuBvedtJJOcozt621eHn74+lMOOwXI+aGaScZlnJGxa4P8dW0Cha0PCnXRqtAR9
GTqLyRvOHz9T/fa/2+gRlt7t9B34hIxRsLR5Z+nlS8aFvUmuTQccDtPm0tryJsln
WASpdn1r0TLtF/32LsqWN5WRPZ/eLwZB+OIxeORVi7glMQnLujMKwPNVO4FQEgTj
4OthE0ztddVZCcQtH7v9O+OXfX/KfKzeEg/TYiW4LDDvk2sgSJloOQ93y5nNGF0j
RSaYVQ9QpI+1S2xEHSUrjjc10y8B6j76MWnX4/AyxQ6Dw+Cc3nUSs7FFEupgismz
`protect END_PROTECTED
