`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C1spEIz9nt21z2C6BF2SHcQM0yEy0aUbYWH0bCdChprqaJ2v4Vg8nir5GOC3SSey
wyZCz9EeYw2i5X/cxi+eHaEbeFrwrXtU3Aam/LkrQIvgqccWB6GPa/DEwkOK8JBI
4MdU+hK5HFECsh/khKidW67q1GxErgaE7fhJ68jifkyJDXmMJXuiRXYVvYvCyhrx
3Fp5exAV/rPLLUfxNMBoYKGaT6VucCqJuR2XmXp+l9hmeY5G9ArF5yu+J2tEpCN9
TldMAw+7a8GQmdRi92dLORBsVBrVS3OajrCddRUE4+gcgX1bQlXjbRxp7DpWCnK0
aYYgHr/wrYxrjy0kLMN7o0yjck8JEa8IlSx6vL0TOyZ9UyLapIUNYY0ku+7rPTnW
DfR26wz62nTokOoNoXD3WwxNQ32quhXZSw2bJf6gOjQ4IZiejjQgBUm30wkzZHPJ
NHsr29KGfLjXTliHvOXoRiefxI3wBVyG8MPMzOljtp0iLtYoeDqqLAYqqv6CMquc
N+5XkhqnESDyA1O3A3BqHqU+4HXsc9oEC9GxRJr6CAuBHLlmVaMFykNNY315IYNB
OTkxZqd00NiOXbF4/9++a1eW9tB7Sus4WIJR6Yb0SfKEb6uS6BoEQBqCNhKaYZYl
9iL1CujZRArltuWev6rLA8w/SeDQdL1mdLLwcPOq3Sq+qjCvQcV5ry4Ep5aRSVru
NeR71O3hYiFewSEDp7e4e+0nYxEozGmRAYc+L8qYbMeokF6nr9jvguf6GyIjMiY5
wshAkjCI2oVmNmI+hXEf1YwU+SsXMFQDZfPWUSkXMs+PTR7DcR52WXhd7XlykaGm
+NiqJqSXf2Ia46lLf3qVsKeTNsTygAlpfLbCE9gW91lOD+/A9IkUPu7g+nRXMDdl
UbP9xpI8yxVS4xOEJ2Y3eJUSi3UP2eZgvZOu7D9QNrZygnKxHUGPh2mGsl8EOgeT
xBuF4tbwJTsR5LlbiWX7LzdF6WdIzE+p3JSC3wuROuMAQmiu4Q2z1lyUgrdsv9MG
/HGfUp6ix56ma69f4w99OCZ9JMwnhDGZUC9v19YkqnZhA2YW/xBBLxVRokk8Gf85
roW/5XlHrWiepHMzmidd2515pDCqSitMHxkp55y1C3mKCJYBRYDHDOZ6QjGLy/m0
IGguYKehKZ07TLwe4ByEklRSx3I2apOOzSZ3YOMxI8SeEe/uOhtEkZVBQTflXhm2
6MyKoJRM42GwZiTqYaLQNlfCle0zNI9HVdT6DKUyFNQx3McutT1Pg+Fp+3O5rus7
gkLKiYOq2tCKFRnoZbl57FtXV+L6PJ2weVzsdczxH0u+QgKuhNaCGchse9BssDFy
jXV+QQpaPUl+ilRW+DRLc5P4uw8rnk7j9zn62P6lAqpnNgG4b0y40laJBu4p/dgW
HXumMfISJbDVCH3d//CCQOVTloLhXxGChXeF2hgq/yGJP5ORk+s33pOiOOsupt1I
8W/KY0ThdAb17qLY24agIid5gETTinViULO4O54PSSTYFzmCPuctjddicjduFABI
XFqJcmY5UmjrC65GQFFd9mZBpaw5vPzu+NhXZCxLq4kXX7ZQraI4pT2TdE6GXoi2
bLH2bX8dgMWO8dqHBhOdXy/qA8isefCJEzUAWrjIBSAFWn9nA7fB2QU2X79WpzrF
zwbDdMBOEf36rRSEyhIOpN0Fj96zgzXG2WOE1M9P4BV+Vdip7drJ11X1BzCk1CAS
N61PL5223nwrCnrKAPbPBHP+MWkMl87yvo7CuTWxFdQUDQAGyYlh48U/o8leIUqu
xl21Gf0J1UtFs50XGoJlBTLjgDORBJ0FsFycLdo2hN7RsjrDa/jcRuYjMvGIevK7
gprGn279ezNQp708o6npc0lMcFW/yfPoXr3gjPUUjzJhXw62Bv6vn0YmQoUZcmGc
Hpwp2avJDcBaYmaqgMBFPQADkUiyQh763gXlHFzM6eiPodzGPWxRK2vpk6m8sut1
4XdIrpazBXp9JkWED4kK6B7w7OqdWD9r6nZuW4xO5szxmmdXCmJXOVqZ8b44icAO
yTZYme7CvYoyrRKJjtg4Y2+6+mJEfylITUEF6IBPu+UzFtxQnyG0jvFvYI6YxcfL
azYWY7xgi3695fSfOunux5i7/Terx3tYo9s7NC/LnbpH1qR3HSdhQV/XTD78W8gs
4MbRyVhEvBvCmI6FcuOui5tCm2daUfAGbE0JeYwqoMHFKsP+PGrKpzDl+nWyn4Aq
TYDHtM/QsrqYIJxmefoJFCWY7mx5bfP6shYrRxrFGg/3GbWQNjAKsPGPZSE4azmb
FjSjrJF62rRAINjri//ShQKDLydwtDjeNU5kQG1GAtm+Ot+IbfY/GPfEcsxj02v6
tlFRpl7Ri9HfBwg83SlrULa4zGWS/2UbZhONDTilaGd8oXifjSY4rpMPycjCnGut
Q3oDZ8yrfOIwqfmAY4CclIEtEQo1a5yg3GGcG+Jof6VGrsI3Xtp2zuJUWrpdUd0S
JWbW6Q+BklT3Ot1psNusCMbbRd26EOJH6LpvctKLsc3IcoQ019+Am8bMNGTGh3ix
EA1lzEV5Eyl1c7PehpavMm9YTwGvSk3qfjVUqhwbQ+LedEVcb3w9UzPuPB0XHFPZ
cWamiv1/ujOeNNgHVfnT2gd26UkrkHNldPkv5nMCsEtdCBB+5sULzZWn/e33EOkd
qfKZ+EAouPgBe1lFc6X1hAOFLbi9Sb2xuWisUUUEAF0RseQ+0FrUNxv+rkIrBwDh
rJL7E2oeUUi31Cx0WfVAiz4A8FyxlB2m5FfzbOHfZoNt/V1Z8MMNxtXZQAWSi5Gf
h46/wVk8kZe61ahaD2fvT24QgGmkGGwxzlOUnaH6t703GQUO0/0My6Ucxw2ziVhq
Ucux4SbWz1xQ4OFqxYwZdPVbmqNmxQ2S1KxwPx4BS3oV6VHGNegOWm6ZA0xUkaXR
cT5NQ71FysKB5PrfSgNSMiB1GDm30DMhwUyqBJtu3mcoyanwD8L6zkhfUBQBMfJq
oEmSZ6f+m62ymwin1uVAICWDTp69FrmpgTqqh78r1Zz0u43sVhexPJ2WlSdOHfHZ
IEWkAI6eHTSDaC8AlodxN11Ef2zvYgN9EXzW0GelrJ4I3TbrmjE1U2SfsqJ3J37L
Za7icvwKTPxpdTYNbAF/kAmY2gREana08NotgdqJg3fE7DVFXTHzLtW0Q4xqyhGx
3kU/EjWJiRB1LylFdxB8HyJKWvaRfVBukE/9mSPjnoSN9jeDSEBUg65nTGtQjPSe
aKcvjA7H/s5SRPHqlHLb7eQ8jY9Waoe5Mnwkbn1ZzDVCXJ/9dU5fKJwBRwYwhI/8
WWBoRzy9neRaIQzQczVZu+waOEwHNvVCDBdV/zUlAJjMCD4XXXR1beqW+PCarBLa
IIiGXAV6vu5461fPEAhwAelJAENy4ulQ6Le4UxsoPOKJL9+iZSWwtFHWja4bafkD
OSxAP0ACmt5uY4QtUfC0AJcoIBM8FYwy4/O5BE5W5hzLYklNgadAsEC5vzx5Wvjs
ZqCzL6WE9Oum2sqhAdTHrxe+urdnAX/yUn7P5oR4ck6IkDEBbR/6EZ1wXnwlmGpl
omHpTudCyEF1PwvVPrz5kZSfqn5bFPC3RiPh6Ex8Zl4975VxsqyjW4PcpL6bBoGv
l05s6aYdTEkGz/3HT8uQ4fnwU1REQFTCScjBgkqk66T2c6IidqsNvr2N6QDA3DuF
wqphauophP7OMBP3Givf6da7Lp4+I6qoiFoioyAF6U2vhQCV70i3jGJjKvWdPa36
CO8LEL0CRJoIq6QAzkWAz7JADOiPJpLNN/j2JxjqNzfzZ2MimERHmZjj9NWebSuK
BYxot5Kla13E0sZbk5XglkOEByruHCxeDeP+2WaobY+JC1YLZYGADFvtd/h8h4L9
NIDGU5GIyCYZuPo637wpRh/qmNi8DNeFVSZ8HnQtlM7P3QhdK2DCDn9vm/sgPMQ0
CuCNccGzCTPoEyolzMr/YTUXmY4Tc5MAdlV8Zidg9UNjI53kofuBkjAqkScvYDTx
7OX3/SWgHAOQ8sGdwqGH0/sm7WTtZm7HHz3+x6a5chG5bOwzI06N6QWKFop88QqA
5NJXsHt3mjJ3+D2HS71CbOWx893frPkihIVM5QxZt809kr+jHu0wudMp3rkWDc/q
yNr2pBJEbjD4gWd/4U9EU+dUgShL5+uGVKw+4VglWNHt5FyoAp+toQILa0+6inAW
zGKZS9ZSrOzdMXUX9S4dfzIXd72q/oLkfXsu5BHmfut1HrMSdyAXWT2ZInkmO1B8
wGsh0zafLNHJs56Opz65kqpHWvBpJxKvHsn5CSLBU/1rv7aX7RbAfehZMWTRkV4+
27tT94qiCeXcbiP26TFlhe/JPDMJ90uKE7Qn1UwjeT1raKW8Irku/6zirs9ebtxu
Sxhjdb/GAOHZ7Ncc1xVy+nxWkDCwwI3OLkJCWKuQ7f2CbJ8dERPqmduGdYI34OFa
HQNK3DfJBuKLbZ59YxO88fVZy3kJRYiH7kqymRLri7fDEj0QYe7FM+3XQNxk4BDR
pywteJ9BX8JOcR3kHNArpPxQ35kYfveyDDfnyYKbUC98n+pgPH+V4aTzpCOCsGuW
aa9fUVEVI8jE9lV6sODRJM2LICoTCQePtAZ8gx4qGYwfP0DZqJdqybMpjkugGxKr
YbjKbPmvVFLxGQU8CwsWxMU/al0hxcdqXlDhf1E1QPoU+k2xL4hlsJyr4gLgL6rQ
KjuyWkegTVwNtZnzJDruxhBVbfLAiAUjZJv8Svx93doJnR8dMyCTMI/ZpZKYTvnY
0n9e63TTbLgoAjoRHNVIo3YW1QGSxFmATqnr7wVvH5TACj6qEnHc1RWaDtPqHhyG
mHgnUDRJWSteCFrMIjSzo0NSvCLIc0MNUgkK3nzUsRGB6jTGsj+5J7Sqe0feeopI
d4ABwWExOdmE+pLXyF+BSDxybFLyHAKQyDRmmGGLu36GfJCchS8hzXG312R07Kmw
i6Vsi+ST2HWGzWTQscN2jd/EUVZmA9LXpM2eF9lLkjYE8utC0TPRsR5bt0ce0XcI
gD0yJmNBgz4JKcUD+5VSswoawR2JRahqEZdsAMHHEKy4+FPsnBLb4lOJVOJ/+EGw
iS+gX8wzQb6CRaWP2iM8VJCjD6wDV+BBbmJGP7r2Rg9QzMuQ5zilt1shNQesJ/8T
Lad2BmelcERdC2pmHWMmuUB16B0PSl5ggIw0k2hsPUsyKHbncXzKAOSdJgxwen1B
S3moU0/p7VHZJ2k2gall463ow/6nddtF3lVOFLfFzaqcTikQMXQK1Kw9+HZHbnu/
oP39ANwoyfvPOFDKY45zD1PH79k0SY2YDBWP8ntDu2U1acffn7dkUWVDe5lGYYCy
8zPkHQcaEEtPzjp5YV3oxmjdlaMR67cvjdswU1BXw52LRxGFcGytmPWHVk+cipCQ
vyThk+o8bLRoAaZFEtGCmtZysEI9NfF1D1szgR51q2wbwE2h5HN3NDWwGsvJ0gm5
YcufdxEKUeKD4uhlbIBDE9jIMTCEYSPeESX8/4zjZyjkJfWZwV+qSg3M+rko8AQq
RoqtlpyQRQPqX2y73eoQIZd825n5bTwyAVY+0RY0okK6mYLHpvoVoxemJyftWwBf
T5AZx1sWjm3lhw2lMZyfbotuhVdY20Luh7RefFNCEjsLfZLS4Bf2LkhRryvCjxUp
wiwFRmZN3ahAdWiO8H2G6kIvX1GYkhwPxKk5zZV0lKrSfalf26gJ0PAfRkkysTd3
+dELQlMWcjmvF4gF5yEt2TKwRehRmyInmnHuIwX6x8gSDB3Gft/j84fAYT5zE0Up
uVJhaY0/vOd5tg+c80UN5Rs2qsL8wU4ZHRFikwBbwRG0qJnjSxuunmi9S3iUMd1j
FBOPNJjNuhUUr4JZHwiqcyOLgQi8DgisxdK9b5oR719lVam8h0OWlxWTBS8LeFGH
wmKrCOaz/JuCtPHDRtGjnB6vg7CJR+spNzFZ8GFLaO6icKL0eh1DSGxogcyfpCUt
Y2VPzqX2kzoozrEArESpw7LS+Pi6yJ/2yG67hYxZKCYV1wKe5iovXQJjNwJPzbmT
xq9hxA6GrCK26Vj7SiI4HOqRWpBYHxuLcAJFD3Jmp1Oe8GjzldpVB1vLJXlpspu8
lAEuj8XNNoye6ZSuIqEOn27tNi72qX79RlU+Kq2msDTWOPBh/hGvja9MCDhrLHuu
LAt7biQM/Kh5BtoCaosC7zlt5sA9p1xz1pIE2fw+da7iB3pH1l1J5340d8h3/Vdi
M43ghb5vvzv8tEAzPph35GHReCIzpQFk99EDgS/HDHNRGUXWistV/VSCh2yZ19Sj
9EByMDkeKSeBIgR/DYQim5f9hg43BZdUUDH4zgCdXXXpmYQ2rfOpVW3HJ4pXG3qj
aeAD/sCMCvcDPcc64lPXG+pP7D6XmGjlyKpXibe8Ml8s9foMNcBH8KYFtir4DZAD
/xPWed+sp1X8cYY80zrd9C4sk1bNXkzzLZRww+rNX/FXShW4PgW9c5chhwxU67Ed
x40jVL9xkhSAZFcJaBFClfbPWpwiiN5Rt0eDDeZBsnVozXzjtYiLCDLRWFLw+tx7
k9ND1N+QY9H87N6OwoL5YJwI3qIJsO36ZA7FIsav4+V38yaKl3Q+6eZm5BfjAYbW
6zIOOkR3P4dQVgjkgSgn+j6mbjX8eoP/Zl8ncEkEUsHOJCoo4uam3AjgHnxyVjo3
Zp8QY99lTYWlDUbrV+bTpgWBZ9Knkl/OCBwVIeFaU2icuA4neYJJGkujuSrHqfaB
gMwa4DRRrL0lXPpMQ58HJ/OUfaZLP3wCnqeMef5nH/7yBjUowPvN2Ks2qPUXOGDV
QkTBwAxm7/avwF9YE0fzUt6Z22GruIAD+njQiJXjOTNsSKQqeyxodEPMO3NNtZi7
Turt5QNRDTpvyn7LcCgw/dAJY9h520zZ3P4l+KxcoEKmYXV44JusQR9fG80jrxQi
7LZkBbGZfccwkD+NQ/UBpOZyWlcbKNRfZRfXkMEbKCXoUh6br8CTdnn5cJ2wWPFy
8KYxFsMizEJQY2kHlpMYX/gk9MuEdqBeFmOr6+7zPA1cLaITNScxtc7kE4GNRr6g
yLDKVaodDe+y5d5719iEJWr8HmmE5nrCAinCBHd24SArq/NxRS1tXba0WDAhxGNM
+X2s/PXJuuIk8HLRkRnr989AcyJCONysCQtm6DI2bQVRv8RAy76EWu1NAu7XqBwA
H7T1LO1BD3/+nss92yc0J8GcoxfXSLegJl+3tB/16koW39N+CSawRrnA/WuXkbXZ
cnXuxkvk+fmbwPj6+NigqcrxGv/CXoFltYUHtk5BxrEJ451tCZ1M1qIv61ChWxS2
K5qcoEKoPHUJzNBfvgbxreMM5PO+Qwtnzo2lMmLxPbBlk6plC9TwMK7upUE50rXy
ROaAWkPFn0OTHpVzQbizhmB8QHm2r/t6+vTDSR2OywOXE6nTpVBRDQv2PvIiw6TF
D8UCi3ktRrGCLeZtzylFjHjWDAvLtnuc21OGRe8MhLQ1Nn338ZjcDa8CUdTbM970
RY6YnJB0B3I83ukumXSCuTrMACSXyXxAd5T5K+fXZY9aMoIoessER/+O956MhAcf
EBzh5VWOQ5SywtjmCXd34WOhaKsfs2wXlMfdaU+XVTHmUpBBIVwZC4xt3a/tlS5C
INoORP87Z3DQsND7bhkkEhRW1SkY6xgnE6aoXeQtFGbVj4uKlegFLIyVgba0CGB9
ek0nBBxdIjObEPifBlssK24vEaayweJKhZXD4mLM1kYTeox7G374rJ9UurjjL0O9
D+YrsJKM5hLFrt6TbeWxGGSCRAevWASfdV+g98rfxbykOSB4qTkszvs4dSBpORns
RNYqKliUCly1Dkgqgjy1jwnbpTrKNKLU4ml/XF8eR4ckqbI88F+OpQJ/la7r995u
XAgG08q8YdzYcmTeKPlBlIxUgYrtPmQHJcOzaPQcFEXBJvaujJAKag5vs89iQWK+
oOVgA6whHGX4ofjySwN1IpUJ+obIQoLYJ/v1H4A2JSz2CUXcUhinWtFGasCiIhVM
wqwVgne8VIGRcd7FbcFhCiY/idrIFiA8OKwVs+Lzs4j1QaCZpphlyEBhsS/XnKBQ
QoL9vzY9pDGV1GLnB2nZMp4F4bvsKCZ+Sg2hbBilIJhcdCK93JrsoJRhKQmjdOjp
/8M/qtnuzmmA4JhZZlGuG2dLljS4dVxJmr2SMzGLoYphBcZQOEviq64znNLor7rW
1yItd3RtpL3vbtxubApJZJzxVd46oGpHx8TpKyVyM8+DI8brOUN+bcOU5vPStXTk
hbZde9XgeyELqSH3ajgAlSlFpDca2u4SaFcX3NfcNjk1JbAtJ1L2RvJD2qA/JYCM
PcC5XEEC/9t2m9wSilWDirakDrQG38yUX1FViaZF+zdw6U58UF16OKnWKpZhpRoW
KThdf/YWNO1EIpAF68aNhXCWnmE1S5gom3t+sXkpVJDDZyQX5Ft+5/vDA1HQZIUP
PREWB+kOkKKxLw6YMfjfy7tDrT65E+E9QDpLhA7oINlJi4OdtCoj4CEyE+AWzmcz
OTFKeAhrdVTlCRv05jYWOaF5foyyayvNOyjQSSm8VzXS2EbH9EfVobIZxbUDMhMl
pgU8S3awZfBaT3Jt8X9EYmkiAZWZniNoSIaIsnrta75HHSH3J4B+d8NmDZSNegF7
0NLbnGa1hoDKykPhl/yC/HtI+660zf7ov9HUgZRbBCNuLwlGN4HOI8MmsyfkHegc
lptUDk3SpS4zq2wmJd+YgKeulT17DvpV4zfkCamnUGgbbu/0vwBkp7Q9G5+6p33O
o2iO1+YSJl+Qh5+CsilEA7zLQ80VPW1O+xfXJoKwaYYATqtjUbyuMJuX9TdYMKsh
XDmlM9qj+afud1H//f8Nc+yO1rWDM31imVevaHGRbtlSyWqZHeF7QJ4cj6HjVR3G
cEFP+xb37XKzUS6b3Vq6celpGEwrpLPVblJQiHwZGDlj85BfuUif4kNxOFbGOEz9
rAwx07lI0kdkPuRZfjiIFtanOYc/wEslt6/zw1Za/hempwB8Vpn4nPvTkpxVYDML
XYIJakLPJA/St2gDKVA45Fhiw+V5oumdelYfqb2k2sFx1Y2368aQB3Xj6lkGuQpI
XsDUgDcozSdihsa3qXUArYcxtbTgmMM+Vzoniv6JbEZWL8MlJWxErZIBvF+1e+4r
oH715vV2AGOZf0YTXO/ZomXqHZaRGqWMutAZn442VajF9RYNnyWw9EHj3aIltCY/
GTOOVU4U06zB7dU54UyS2xPevmU5lckIhMkWJgbEdPaU5HM1UHlwxJvR0yTBA4Fq
I6eWJ2CkLbawg1zPgdbKrVtnGOrRsZzXuiIYiyqwG+AzvQ3HUjmd4maemDtvRnyf
G5nawR1qkr8GETEfmPSGmQBKw8ntHYuo3Ztd9GJ09ePuXQKu1ZJKRzAXMsuB54cL
4S4rWjIY4EUyHTX8nygy1+vj6/xH0YfoITfJG5zJMdMyCAGXIQJf02aAagMBmZD/
jAa0LAX5y507eETSxOjVGcsStHvSLM1MRg/AKf7XtD3uWvu053ywDQXyEapZ8a1o
QgjYKxw21ZuMhauIcDS2UWIwmou9SlNn532iKaJoJN9/ilyV69aPNeSVSr4B1Zis
GvevmtfcT1LM9td7G1KMwqWZR5FUbOV9AZp5vtZ/eSNdJdLHZAAZueKYpJIOZW8X
8JVcbjKLb6zCvTIaugv0mZ3nj2KDi6jvts+X6yY4kecunA4W0h+ETyClmBcDL0tB
f9QwO74J/KxZta9dRFkbZ/yTh7tuHbAwUAl+NPn/9PB+m4rg42oq3O+4nKnhcWru
FJ93RlskhA21vkseb/kRWPMMoQ2pf0JVaynoSShcFyaAj+Jsy8oCB6V9Xi9/iU38
AaBy3z8WNqmh0BxNqlbpJJOvxcTSXcx+9vTpMI99EK+enKkLd/moC5y2Zp6b8hPw
KgP20RhGyLQQois1JtNkGKueCJIP9P34xsp/pxr2dJ8jQ/03ZXBkCwa9EM0DcgdS
ZYbtKzQkuvnsW4FKkm68d4cvjseGRGSB53lk68TV84xizfopltlWVZV1TIRU7/iL
JX03BdEBi3rpO7vYA+slB6W/SQ0bbpTRddT2n6HoICp7/ZaVbSwp3FFAAEUeLHKO
6RWeke+Kj3NQ6SYz0aw0xyeKwbfnC3QZLjxNSW3XQxDI/BYyqvRpqq3yH7/pAt+g
RtPLUNbHRotpPce6BjSU3rxNjDTubVuBdPaXx/EmbxH3j9Uj57wQmJyClOv+N/9d
AlaXE/jo7OWmg9iAXdmm4Han0vIpCGzBJZQ0nFBIqXEn8/aY9XJMQbI/o1CJN5GP
Z6TgiBWxmvwgCESyeTlIvt9sZ5aoCDXJd//cvpT5z0uBPNEydI4Ai1lv4sVBx9TD
UZx/XebIRWpm7LLrfOWgtH28GOLjKUQxBS7AO5vFM0/iXfdi1VmlFHizCCEJsp5n
2npvf0fU/Rr1Y6KrIQJozETXfHPPZyF+qAC75UjP3VifJrgqTkOvf2Gz2PoYAlfs
sFSUZiHKPRkVQ/WihlrxTV45GCuOFavaa6emUp3++COW6DltAENfozvh0H00XIFT
BmcZszjy7REJvtHf1dJgi2SrIbgCaymlZTkL6Vnu3kKCswPzim/yPJiNA3LQV4zk
4N1QYX+EeEZz+4hHm45O3gzZx7ApsEeXcqAxv0UXS1/FqwG4pja/QRCZ4r3yxLlm
nBbrWLYGS4xTPVX5ug2/M1RcCA1Cxr0YirzacSF0MrCv6hfIRXCtywRMT8POB3Xy
pWSsrfhGKDxUSq9sWaN+AbhtCQrpV21QCm8YsT5tb0TH6nKvS+XlS3ZXZhWfQLI4
yGeiHw6nHNKshazRN238K1AuR6kveQIJ1bOzTrsR/NsIbxCKB7snK3jnqUmPPg/2
Ejhw7muV8N6dbLhKfEqdRrS5sZ1emgnXlqovNSy4mf0m4pdgfOJH2L9H0+HwwX88
J0i9JDj7mrb18RLnunv3SSGWh0aABH5ePB8fQOfmyZx+Ew39jJs3L0jA1weBEjbX
RU0ewJZS6ZPvBVLhTc+eKVt3ALG545+KUr7DwQ1z0pxpYSOSA1Zpplb2ljXoTwnY
ura35KKeqMSjxkHb1SZcdJhy4FXDy+57ofw2wRHZ9LuKkHDygLLfS1lC340lspVC
G8kdWs+6SfHipe5NJv4ven44x63L4cagoKm/A6rs8oRislBiuLd90rX/GfzxvYd/
gfNIA/duU+T2wqhmvgSUj1PTgP728kg+qRdu/qw7lFsL4iKZkveYKxr8eK86nmAm
ybaZAcELGQuXhjjigqLBCudZ7A64fBYv0yKZvl1AOX3g5zzgnCgL+/MEHQGCArm3
OOqH4yuuymyas4tVi5dz+j/H0w4O+hG/J3mbbx9Tg3Afhc1PaBYrB7IRtog3JO5y
W+z8UGXF/U6mgMYfnNPn1Aa87s7tSBwIIh7/uTRLQaXHqRmOrZGIo443rMoYhqdJ
l4tZ5bHzCe/N2I4bKB1nG9nUMyiCKtKUBNXw6kYmYaaHB879PnWq9OGdX3qsEYSb
dJOYWFOwZXPp0ik0QnVqUxTyQ0KPDsDWvK1cnnorw6vFLCixgbgQazWDkqRYMrHJ
NFewI3PkpQGIldJqMSv/ER1+F/EFfMhcM1Hz30JVMjs3u4pvM/C+HFlUQ4zZCJ2B
T+wwBlOj4o8BVnxePySRaSq1RRT+g6z7OUWHwXwZy5BhVanqw4Ie/mof8SKQEeBX
tezuoQYiZYShweo9yfeGD3vkeQJEBu4sZdNfPhzirdG77Bgx57F9/8ti7iR7okRI
3LP/NT0T4ww/Oad7vBo16pU6l2PkB9FnqtQ34LNiaW+QxDAoOC6srksylQH4pNMP
g+3eaz8YKOwcTqipP2du4Y3JK5Z77lfjme+Wq5NKV8R/Od18ygdEPIwsIp6fzdyo
hiz1lTwdSDhyhQWkIfOTZrNaqXt0/KhxAb56c48UxxlhBxJG5qqFZmCFokRAC8Bc
y/tUMCRt0CgWZUEIOewqhdiXpPZyaCImRBR0bC+oJN9HSsWdudI+P9fYpPqWCgEL
2abcMmyGxFzqjeEnzNpWpLYzw6ZglczyVM5KnCS9A2yd65wNxJZGWQXO/ayGij9W
tiXWujbXahdGijSSkksPBGqyyGntp6aeotl2Br/4mEXqRAv5allHtC9xJb8jbo9l
1gm14Nc3dSDs4ZbjNBNAbe8Zu9TJmNfBp/snJHHI+GggnXf2/HAoo39X1QyKHp7l
YtKshnOakbkyrBzKlpkGsPkc4GddFlKikSNyuUYrAu8zCgpRebWy+6g2qqkKE0wF
4zL7JZuLqQSWuK0ksbRB3aIbfVFR7axlSn+FXqfTqnq+yI9HyDUP3OnMqMKCgx9r
B7Z3P9k9SDuUjBDdonmAESDSM6OBHl2SizmHJR5MFeK98vh8lk+75Nz7Ez7SygUc
wPwhTryMTqQaDbnzRdhcluCh2OHoUesg79jBugx8Wpll/O9axcL3WU13GfGODxjX
lA8hyTQVkPAVp4EX+D1WQ5JV2qYExuadZ3rAb7ACCHHcPDUI8t58yA8sDrpZetA9
JMb2qeXxVK0O/1NTtjh5DM86vecduadgpU3zLKz4GQpVl3OVtCbQdzjgVfcIbD5M
Kr7lDiolFYxhjLnVUDORSQf+GWKPxatRt1OQrQfQ5o+Vd/jMOGY43ep8ACW0xuT4
q4rg14sK7JIUEerPOli1JzcH8IYQAkHS5IvGLjFig6VU+E+2epy8rdB+tOekPL8x
LSbMsWkE1VBSwPhDShk82SIuQuj4U8Kpx350ALPpHjILsGYE1hDdifLbNQOXXKRn
gQInQg09oh5FCSLctl978hHthRUVsNCC3zSFrfYekKTkeVi7sqApW+/7zoR3Gspr
fV/U41Oa31g7/iCu8X3dffp3u8ZSdAybsCyFNgvhjqlQ0JzD2sv1Zg96EoQkK4/7
WA72KIvYk47QehQDlnL+3/lVSAJg5N6tNpSNnjuTFIUVwffLOKqFmkDfpzW129rG
M7ciyAI+R9RMQoA+nH8i2NfKZM1ibkmFbAD9LVSiFRFsyvMQVLJdbbzzXaEMnCD8
eEZI4M2RJZCWf+JUSwCufQUAIvwsJpAWrhPPuE9AHl39AVAwyLQqNYWOq0xcnFul
WeDsR66aOJlNScA2a4CkyKVUpJ4c2Q2vkvAzoW7wRJdCjIHqBBbMrTZF6afEF1os
yX+oBvN4OplC0s9vrK2h2iRUKdaJhKZSqx+Ayu+R6tSpDHk1bhSu9tBD4DZ1yyWZ
GSgt6xtY4yQJVYvgLA915STyPQVdy4h62L4Z13FgHAXi/MvVs1RPvCUwNM8ZttYy
zhPyTJZL7ud4vRmAyDWoqJqyoZiUvWq5O5k3q1Jm/OO7pMzPpQT8vn2B4gBRE9ue
9VPJyXNcNoK0AQqrQLE9dN/vtvDpDD09EUmc9i9GCphL1Cku79kBC+77ecAvnMsS
XpNK8xI3Z6ihCRUZh6FTF6JHEH4bH3gVyv7f0Q5tVLzwpRGJoV1gD3nKg9cP+SUK
dJxXdDhHwOvzXRGU5YtH5LmrPvg0/L6IxpMBu+j/u7p+QdLotPpncuKOB227q2t6
sDW1UAlrxsAaUSIEWPt7ELgxmurxNrhg83DJh1LAGFLtiWYIJHTgflODR5QU/fqn
+D8dQNSe2e1F5SnLhugdkvOEfnqY/AbBMxM2pLG0si5PMuromRq/i2oY5eVWoA76
NxRne5vUG/C8s2SIp5xVmLiGu4DROKAE4/kqM1ci6Qc7Z9Niy7ZvDc7OF+dMLpla
T4Nb3DJlIg6Y/Kl4kL6s7G4ogZVyEHf6aPhjESeXx3y6kS5EnKdT2Nx2U7kKd01c
eWPfKOQiUToswmsbCDCWazJu4wry/4AjXlAFzfaYQ/KksHWm/eyqy2OYyqJFDRVq
qDQPlICYTGPz1nddXvR1qbw3q1S7PIIb734TOJVPqZD/MA6SwBKP7kMyCqp5XaU2
BDRD92bjgwQx7t1W0KLlRt36d+aB1lOyZmKmfrv/EQoA3pUB+wKiFR0zLzZmiV2p
UReUIENazrHasHE/UcZaQK2PorhMTPD0TsfFMryotBqUTIwdIYOdsy6Mcz+0e/DU
PAi12HQwYXBqnDSAPc6citRxP/J9w2dzpCEJvU+sV2X0CvYdgI/W+sIJvA/G40Mf
NElSELvZOENta6yYoUVjcjWlq4Ws9OrcJBppy7rTmb5yOt+NU0PK0F9wF8/pgOJd
A3fmla/lpcoCu7TDEpALZqHIfYFjJ1OMy0ak3yn1zt6BsLwtfxbibSuAeIiuRu+k
pVE0H980iDl35nMvxt6jNXO57f31FvK/W52MCM5zk4W0TMKBtRoHxpraHcBC3O1n
cRskQ223Xmp950Zc1QfCUBRXD7o7H5lg1SYEGZ3r67XOpK+McTD6Fw60U/Vj8KIS
QHdwg/WKXoaZGULM9tjVdslCE/6zMi3Z+AL9SpZe6agfCqnW4TaYYS2lU9soKPJw
w4RyI/wI2WISp4kUtCcBGLETFp7acERs2TUU7BSa2Be6bZhS+yHejMwznymzaW1x
xdWfeqpcf2Y1VY09MbjRbeGbKZlu3b4GUHdHpyURKXhDtKdX68nJtWEY2wrUBm5Y
ww037QgTzsHCOKAPxZtgH03VD59j1m89cO9hYmtQoDjzQHfJDLU49qLeXMa5EiEy
B6CUS/4jPb4cU7A8jvVAejVEUXjUILsLc9fnAqC6Qjrzh1qqNbV2mNG0cJOPZsk4
hGFfk6HGR8QXlnng9wdBlYMe1MGGcDWLL7BEFZUoMIrqqw4dFgEdTwmZebDXx1Im
i9vkb2IAvq61za6FsfGYXeZwCNCXvYTPTNL9ZNoAa3l0+gY3P2yM71QxstvTfU/4
8gTX4tadhUKo1kOOddFxihLHfvj4E8SmnPvJHwtzMwj1QsjuW3DQMpD/xaBq3Kjb
tkrIBRw8804hAoAy77Z4OfzyMZCW5xFZDC/PGJ4Z463/tKYiYWxOM8t9UMDqm4pH
AFAWjhUhE3v+SqVczNJPLcL/6voro06iRnPzEru2r7qBc0/e+TpU375fY20Uopjh
L7QQsOza8mOPAm6w62xYlLL98WH0ujflFfWHixt+I9uVcxmk2EI0tF/B8MdRDm89
3NGohU+T6lmliwNRBgIE6NPhgt1jQtYlJzgGLwA4EOtyKNv8cyiE8vZPxiMQY66z
H5sfwxHFxNC5sOC4tb1N/GvdebLsLhfbWl/5F7N3bqBiIt+ncdk1t1WaChC6mc+n
uCYG/kHMPE8NFuy9DytVuP1euhWS/dOq11jZkH2WDF9PDPIVGVnqaGS5TYbOuYRX
FKinFrIa27bGLu+cfLJQr0uCBYcikmSPFp2LJmw1qHW2VTGlK/Kx90NbH5spKSw6
jxsQLCHrN+BCBxqZ0lQI858/oU5HEeX1cILlorAXQIiy7QY5+eHgfocNTtaq1QRd
73GANGTJIjL2gAATqtWBKN5jmR18KZXJkQn+KODgS+JrpXZAOycsxaL8KSjXRQUd
7Z+EuIV3LqS8PGR2h6K0BQJ6vJDqYUwNSUnNzMLRo+Dz7ht/FsX1tF8obJZ9aBb2
hTV83Kq+4VXb/wGxboWmcgp/znTBPsJFsjqD0IdYBywecc8pvxBQo5pCqbX5Qcva
9RG6rlGSVqmzRvSiDQ/F/d8w22VSC1Rrl/Fg+cY1UpaOBuAb2aQ4Vc2jnTxYlNgK
rZflhYLxJDjuRTuoNqm5kGh/cQfIc36ZvmtV8q+n3RIDWQLf8QRdhic6M6g9k+pN
JLKT/1O6iwafuYNeUxkg/wqP9WE3S1ISYqOcZi23+JTmyyG4iAMmuOklCVpDwZZ9
m2GVitQsVhoEwv5SbuGt+z5HWQYEi0jvT9v9uU0jNC8PnX/MQzdQXvtN2xWsmB+r
uISqmKen9n2GVgTzfpgwg5EQ99bLIjEsAccUdXFigQmjEx256579ETXImrBGzyk6
v0PqKg6Cg2xlyLDOL2FghtQ8S+0CAaB5dufYch4gQdxO4x0z9jQfbvUGESPbHzTC
MO1RD1Nu9cf09pV5u2AeJdlpCdVcwQMVXMWOsyCN1kxqUjYmTClQq3ryNde96Grh
I2p8WpYhgWyiI1K/ksVygy5m9X5YcyXma2JcjYy9B6+2yXSpkpSOUl91VAuLztEk
vLhjQ64cvdF5mselGLMeqDZdOkG72PugQMRS7OQvK3HQlvMkovqNaxo63+0Pu4Oc
mVWD3WJjaY5DJTzNyoXwlOIeJ86i0NyuigoTePzLIEOPxbbCPaisaxfbAkr7nAcv
lSmcg8/vtIa9T8gDeCVtr5VKihO8zvGU/SoaHO05ru4aMrKfrCy2NRA8MqKVdW14
fZ5ZonQVyv/USur5yv8ZhsKl5PlEmIJTIRHcT/sUB1ClVJPXElbveslhuIqT8BO5
TGI9dYj39swsfeKz1Q9Nz4dReXGXK+jd5dJcp8wWbSnyBE3xKPpxFKSK1j/fwuv7
xlbxXgVFg3RntLRMlfGLslhEPIv1vifWjNEnjuZ30eysFGNzMKFd/vBEy/5O5Bp+
PZ7DxbT2IaT7i5t4Jgx3tupIULFxkU15MDiMjc0Vdebh5pg+xIA3z5OLVQ+DxQRt
7yiuxS0fHHjOOcQHYkIYnrqx/j0byHmg5a1jo/3PyxNrLa+06PxtKiao2p2uoi0x
0JS8rBoSBrcII2q1/ZPmTIih/QOZwNEVjMiCB6afaKwnv+FQDoJjyoIlzO9697o5
v+YZHGOr5146v9dad4WlwzdsWntcmg3EF3b/UowixM+olOmVggAZYWcdigFYD/tZ
XVej7eTxo3LXSdNDhLbiAuL1/2hrIDc1me4Qb4gDyvPWG4ERM42C/Dbfukek2Pz1
MjyMQDQPbo4V4LO8n0jGkxjXtdmzeI70Ve7jdZUv19JXjyG3/rXFxBBLoLx5GoFB
M9pqt2dhHicrrEH3d8rlkpjNrUWzuwtFtMfD6mUjjjBWdEP6H/DX/42dbMjzzcFQ
N8/sJEdp8tSH1lMt64jgTIp/9VSzynfIi9lDdq0sjm+CLORBwUwY197fy/EELrOs
7rgPuA7I6ArjArOUxhnJ4HYFYts/t39WXJlYHXSLTIVyhLTaXsviyhEfMjkOoYIE
P3m/jZqus4L8W4kX+jrSUJePMaz+Qx5I3Es8be9Q/7qGP4uoZ1ZJtK+7OC7ZUuXi
CqnzYUZn7d/dMFM17HrMMXjngjEBFpGJ3CnmuCcCYafm0fibFavAAtu1A+AJJRvC
iN+rhpjN+1DJSQ5a/nvKqEe9Hqm6unN7t1UYrw3UYYJpbTvtueS5XxB2J1VAfxSd
w/pPyPI4+82wbbUbfvqjhZrj5YceUJS6DIhE4apaPOJPd5WaXDqmsKKk/1GRuDPs
o32Hyy68zMtK9Ykzbua/ejv80efWBcKHa2hmgiKaxik+dws6WNsmo2dCWChC2DlL
/Db1C+Vy+GjnYdQJC22MpMQgDw2Vr4d2ddonOSkjaUm+c12eoTOukrs+iXwDMjXb
38X2E5of9M0BWjCbh7ntP1RLVlfGt9IibsyVxmVROWyy46yWfnBCbkFn0UDg7GQL
X38TbckJn52Jh7Xp8fooet3OYzKEK6JKwSva0jF9rj/xN/V+lDSjWZmGGs925Sum
c4iBqaP0IeFJF8HaHG2y6S5eZtbYLPu11uAKrzISnRYbeu+MQeevbwAtT2JdrWDc
Z8O//rYX8DenRYbyKImTzw7up45AbT0lFazH+uKXlRe1rKElI0xAnGtt0LFpjm9J
F6Ybk8Kibf/o0A+EPATCmOCfmfjuOL/o5zSh75o+7Bhdrd/NRNYOm7NXOPsSGuTx
kIYQHD76CnNa5tU9uxl/UX6updTw/ff+KDhjUGCtIPq1aSge/hlVgE2tPfMlPEaZ
OXhUtsjKlWT+jVNzdbj4ywsUYG7kGA4LPqmRrAWvnpS+H0yIsUBbGaB7XlI1MlRN
Xq9kECuJa3xZ4XrH+id1F9LXCD3k7QoRBJ+YTTa22BQdaAJquWWI/NvyD/W/sThN
SPDcsgviVxVj1fWv1duZHx7aIQ6wK3AfRqLuZEChXDy7PbdGOQGBwDvV9u93KOvO
09aWvqWpHyLiCSsNqV1uF18F52JX/OO13KKtSXtOgqPR1DqdiIVwEyB3CmN4tLD4
x05F84aKMDvK2CYlRndbiOxm8HdeG5WEczRTY/1P+lF5YgXDHwI06Pt54Bq514Qm
5FTlP5pBbKZIrSZfW7+CEWHEpNcCwUe4sVMWRFI1zvlkh0AINQrAa122OrH+z03C
kjI0xJa5x7lYF3RxCgEcAYgJXjbca3HuxPbHAsDHZqIG2yb/CQky+TH5G+YeJdUE
MpuXR0QHccevh9l0Em4F0GnJ9qIKEWqin7fCDzntKNstlZFjncw5hI3AOCrot4UM
crQ355qg+2lfQQN75ASQXFGdvH8q3Q0Pv0PjCs39T7+mgL9zPV9xP9Zdgcg+ZREr
Au6ME6G0NNBnxwu2c8+5MYrBXsaaXtUU4kyK0XeDj+ZsYBZ1CDIS/fPh9MciP+zE
asVyN8VlbN0GsluaLxzZQ25B8XQL1WmJZWI2fVd3HHckeixxFPLZ1LcVygUPxdc3
kg33QuRh/HgPw98QKilyOA18qBNxguw4SdsTfjhelkSeBfi8H2/PCTlpuUZ1FdPQ
l7twYKkWs9ND7qeW9PSXnW8FTt+HtGxlqUe+YAVFwt0Em2gGUcdi0Vx/fL6ptjYQ
iorod3QUs8fu5nZhoafom4aL+L+sVQPqwvh2yKOAqZT3OimOAyVHqIwcCyrIqyA2
Lcj2gVkIKDXVqVWNGwF53oSZ7XY6LI9QrQfjMQdEcyFvf7F7gnq2LnCDMuW0hmUl
cWJryWPc4hlwVX7pIU7enHRin/qRpIZGCXMcn9TYiTPxpzjThkD1jdxtmdSm8l2g
oQFbaD5rLUBo5oZc6PsmhwYvxLxAc1J3f6grP6pbBBqG2pYSW34WoU4H8MtDfggl
efLbVvGqTkSRMI+aS4Ahx1BxiiV2ERRvL9VSP1LImCxh+v/wKnmq6UXa3M3iLfAS
qCxwlqObvPEXdoBJ9FrhOsvd3jQIQsbPJ2GE/q+J1iTqebAlIfzGv/R4ohT95Ctv
lyFrMbBvgGqR6o8A6ucz8v8FEFgCKPTSSBG+Y2SRLl8em5nws2uzihXIW9Daybmg
3YS6xztsBMM2gujd624l3erOFUY691Qd/RY99eFnuUGGUkPNZJ3V9iQDg0MU0r2c
8U2V9A5fiavHvAoX5uLHNlxBH2YOZ/BPOtwN3dUCxp4g/u5Uu1oqTSgm1aNvXpPa
j97j3mF7QE5cfo4nlm7XV++fzZh0vUVnxdPXlfxN8NsDoXBLg8NEJ5E7ESg5syDa
darahSsi/VjB7dwZ98b82iFP5wecXaRgWzVN69qhh9KzZNUcv1cUPc0jcBads6qs
Y71CQVWd2UsnhqSelrVEcAU3Pg6VACw/qV2L8QloSa+BmcHy120foYwuZaE40o7V
df4kzFbeQugac8J+gjiON7CRPk5uDt6RAWcu6IyqK95AQ5avEYQlr1eFpT9+S7St
9lWgUNgXTiOt6WVNFNG1FfRTl5ofItY01NXu3FDfbTytYtPFhQkk7t1YK1JRqWtj
blp5xsc+3NYUjb4+ZkCtwmI8GV4Sclo3U4AbCJl1RlhCz2Q64VbOQiWra+GylT/W
/8FCu+Rj6WYdv2kNdHCZtVc5Oj42dMtgm8dk83s3PdsjwNfzGhgDsuRbxCWwGO3X
reuqfday5Jk6VXziJPk7UcGRP2H6/aHZ2niKxkG8Ijq594OLfVG/Dy8/mgW+1Tnc
f7ZrD9ZyYHqBkTgLarl01DgJgO4fW+1T4kX7K2wIMC8l0D5QAkitTt+gRpZZX5GL
Ufu2TDplIdZnCn42a03aKyX+q3TNNNTbPyKLCh7mRUNDp2vrlF5OHyS70eERDy+n
sZbYiK2QogmHkFlNrvAF/+L7xP9YZWDhhRm0BBR+OZg1nW2uh/Zf/HIHrnHwDfhf
LlHS5MrYUFzTU6fFFl/himtbm+EdosgrHsqDvnzN4znie64Up8wsmta8hcW3xonW
E73gejRcjTTgTLTYJ41a2R4tvR5PnnM/KFK62eto57b5I2VJc1jkveuGIguv/lEA
0ObiBQmbrbiIX4tgAed3PT/rd1j/yzGPDicfUhTXJa6gCYD3guK5h90Usl6u75R3
x2jaB6/dNT47ZDNZrb79j5MuF+dcmO/3VNjpFfgPIsXOUniNLytrk4LPVZ3wlGon
E+GyDAYxhLl9bgG75/7rdIo8MyhHja5ACmoBdysH9hAGMaANzbITD/JTEhipzyxh
x5le6FJApDVilbiHa0JDZJlsAsoeyFUq1IWgDqOvvT0toReBmLt2W7O4ck0pUIxn
99RDqoBU7tV/ioehKPjsPpokr1noR43l7ycK2FYYd5NkqGNlXrDoSvqVXc9Gbf+q
7StHAz/Pw+JvSPtqgu3VTCHCKiSbOq8gaEPhn054j3Y2EndaLnlxRxCqzQ/Am0Em
6pWK/dP7NQdRXZwZxQB8FkxgpKXeLGwOkH2TMXvk6ZWfaIgV0YVwbE7rreD4Qbrx
4oSAX50cJDtn1fx5zET/Y7XTgu0j18J8FsRyJWPECVsX/SKYINzNUa3OPPklJQzX
auICPIlltmBjZlLoRWsfWUTCwMgjTNANJXk+G6nQF6ChrOexIctOehecjJen4BuE
8v34KVTUITOOcfk/sbe1f7itXvUSX/D2D2GlPISHQgPtjljN7OlEprwRALoqOiDr
MwQAJabKo/YP2yoI99HM30cCiNwde/6/wt7Pav22zrH3D6wlgAgmIviBaGKY82Tr
2ifgANy5V5n7E5yJHxw1o7mwBdQrNYf9wMSg0N2fM7h1pyaX+Zj31e1uUA4xlgR/
dUaIqqFgs5EZnQx+VV6vrRlufwB6pjQbHRoBU8dDRRjszmd4PkoeFcexlo9iv3O9
YLxif5gDDZDi9AX4i4uxpXRxyA8nCGnVFIl7ey1ZxMxjLtibYxUfGm0ioMcd70af
s/LJH9cHIwSzMpMzVyzjVDtx6Esoj2VFqtsH1/GoNVi0d/IRlg/mj1vI1qZi29rV
hs4HPgU73VXEYZ1JrShu4ou4KRA8WnOIZrrxbzuqDxARuaB3ZcwGXXyKNGfxZb05
9urZKOq0v//8AvfmXotiVbeLmT9qY7d+sbW5zRbLE0YUuRXaBuwGS5ICPeEzDzp1
Gg0Yrdkof2q3HHuYSQ2qqorL7ku2iM9G9yq+KJ4mVxp9jZl9NWPDTvAshmiDXYJe
LQdAFFy4MqC5u3Nf0PKD4LE2BriKGAmseDexCaP1pGrfZeuQlMYWtSU4OkhUVMAH
e62WECIxSHn6zyQ90/y9qDAVatyTPHLmPn9Vp/nfK8kkBMQp9J7kauJyhumfGqKc
BzQntXKU6DPIQBsM8XvPgarK4LaiDubgZuKvOwNrjBcMcQgjBFzvItH/OIHCyQLD
oSBp6cRAQPOeTrZxBhO+tkofnVWDnnh9WcSh6SHTINnuajfjrGXkH1WVOvgjyfdP
jTPmYDN4TAniAMg9DJwcVTAo/Nu4nIJjkFO4BIFUGW9tvdBb8HT8/VO/eHO1apEr
ExVtYUb9ceEnlgBRHvd1jFTdYVdAcRGiXPgq9xc2aycdMNdX+TPP6nMTRnwo1Zdu
UnX1n21Cghq4rnDfBgeUHfmDJPTG8A8yUxq8cvzT6JUcwoyI7FhtePnLAN+YnJTf
nwcYD71MT8AB7CqGlsu+qYVzr9ZeXs1Q0yaZRe+QUiTneNfdxhbGtWxprPpVV+B6
N/JKSMeaO5xGQPebv3G6tU0l7a9/JEvPQOBoL1CrjDZHS0o5Xem+aqEhuZ2/LxhM
LKUq/t//CBPqGdV5iz+4fm7K7LLXHMHKu4WDZiGrWPUyFohsTBSMD5Irj1gCr7eO
WQAeg/nd3jmYrR+3FSeqa6SGFDKB2rEBPBKZjvZhmItIGh4bgntWC/D/X2gN5daU
WBGul7LCnL5s0fHLf6Yv6+uXqcZJRF2NR07o78b7eCOo6qBCwGOWhD82Yx6VBKmC
D57v8+79EttI3r+WO+fXBdgp+v67auVr+UoAFFt+YKypoMKRIoBtv7msQWSfRT04
N+m4uX8N7HGUnT52cXwJSl+ug5noe6lqcjZI8/1kvmk5PktpK4fg7QKRarhXgLJk
1N1sdXUN7a5u9MCq4Xp56spjfZ+7w8GC7gIIHgqoULnok6zuaBPRwmRgO8najil+
x5HGwEzCKLXrh01iqVl+TRcgFZ+8Lvv+2YJ8F+dWUt6GE3MES0fZIf3y03FItGYL
J1XHZGMYb3KF+WyK28IEHEpyBjRhKst6UpKfDg2IGzN5ZVYsPaWC3SlP4qOLps5B
bTjpYPRD6Zy8Ge/pYYglLhVeol5VvOEmyM0zK4GwW5Xt9KwfYQn5qAlOFHvl0RWJ
vJVqOpS8AV678/Dp8s2ylGTooFfBgqiJvVcHV7S3P4azifT9O9AyatXJ9Sf6F7Xm
38LdrI3BnWHOSzXJoi9u899jQeVoTN4YWRV1sU1TBlf2SW9aAfAqJJ85HS5THJUE
7eIo/18tQzZtyB5o+CSgeahrlQgGDtrR4RbL5eq2wRMEo1v+k5GFvRKfj6QGhqtD
ndeKRgvaijieM+4lwWr1OfnOOXlv4d9Cjiebhwk0G+/zWaApTcRUw+5m7JSo/Y8b
52xI1v+/BgtMCOjY4X+AExPGUIbv39Z/XNbcQ6oD3USaVLufOESDbZlHDwH4Oh+m
j3oj1Gc+CTHgHVMHCvosVN8WzXCmb/TohC5+2QAmJYJDKjraOH2FQKQJvljTdS+/
54Ey8BiLJf7jUgtx9xbhPJbJNVVScqFdjpNEJSVGWGxtY1aJOH8M0+RQzrqssQGs
DBU3eYZBYNUZCYqX+IPS4pVnChgLLUY2SUhpjQEjVZlmorYApjfwbsXQIDfYdpDy
kDkef3N2lxgU3PLuHN/PEyMUntB80420DwdfcRM5wqlKeCH1/T5Jmc2s6uW7MiRK
n3gw6w/Dlth76NQgRIZm/dAEVW7ABD8pX48Vm2ss/MAVCnf8QbkBEJmIy+cErWTC
0Q7mCUS/BGdTOEpFvji0RFwh5c7slp8hRF2xqPDt3hp80bs7hxxrB++UgQtYTIWw
UlhsVZQ4HpIsWXL4rHAw+aohFSsx0gHNkvUBQFO6E2xHaGzsfodD7TJtfJ1B1jCd
5aGLY3V0HGXK5xZS5ZuI0bFOyqHzSV9KYsIdMskZMOb7oVZKxZ6ihsapiSl/3F52
hd+8AwzdRctxIDNKvCMgJy14ZmwaLbPWXEUZMZkJkZrwUM3/3cxPqegcC+o2XKj/
70XCfXbqIco41V4FFXfqBWwBtM4bWOuPXFMi56/E/4IgscaZ8nNf8ce+LYoFkK/W
coeOsjjfLUH9rhBZwCXMPSFxOKhtCDuBRDvdvPT6H1JeGi74s24P+sOTCQTAFlSI
6r3KxuKkFb6+uQKqy1BvGCP8pduBTjelsW3vamgSHEWKhvkI3aVd+18OqAKku1dl
4el2LFCDO2YnxRjAfNgJhJO09eL0KhpOEaG7f+uUOWyZAJEPXj74qDmV/97RXRS/
bWTXbliHirWRMBEq0ltcDuUc6VSPFMNsH0zk2x67vS1H5hSJCoslEdlmsIPQrqtl
8RUOf8+I7JE72kh61h0XedsTG/f9wY8NEo8oxDn1n9ebLPJKPpGlLwd+J9Bydd9N
6tjDgyuq53QRs0C8tNwmTqT6SIgSc6j/KH5l37Vo+X08N7ZA3en9SlXtMt1hkBPl
ipmEoIvUkBF650pdPsWJHxtPlaebm871ioFg8EUbZvCkniFk0BjU31pxaCbZCtN+
mV9wpmSzNhr4j8GuPtT4z7XUHrnMvKA+LRjdF9nCiS5w1CqrazNNLtoaAUFkyPsd
O/yY30J0EzAjfClNb8I2h5H3YHS82nxcGuZ7gr/gB/dq9HmF57nexYEFo6byTyU0
yMsJi372Ws6RgLJEPQNFDHGvRnSiLWpLwvMAfmWoslXWE4giGYggBpeDXDKeiUws
zKSyMhROlQ+nxpokf8y4MIMW/QDCnnDgdeepqdT9oUblHS7ZMldrOaBFHP+17Or0
XU4oFSt0Hni/Q3iziowgbHoVtrseCccONN8Yc//CHHdGIQxiANtI0lHLcD/jZ6fz
Jced+IMDW8F/SO9fLhamJz8ufh+5udw8J9S21pdeTRxPqSim++LVPOAsCu1iuKfl
2bOq6lfLahovzrgatoj1/CTryH/WiPYsL+H9CUpVdiMeYzSNtFIhnl4hCaLpUTyM
wZqjobO6Y19bO13RMx1AEnCUfK0fh+AiDeiwhjk3s00vZCxHzh+buZCqXiyGvGQF
BkRIpd1Bj3T0YmwGipObO8vXyKLCAMyWKWOFrkpuC+ss6JjOOBfyI4wLOaH1HjvQ
AniJ7216E2xaQBsmcwH8KtRofBbt4vamVTlhkBRMt0Qau2/42ujSLD9US0da3sGH
l47cNXihlfAkgH6SCy6nwc+z6hMqSclepEH97d0uMPj7TfE2GUHuE6EB6PgTFbWa
4Fh4qHQc/c8PyaEkF7aYkVrmKtDeEusWGBAK4FyNHxXPJZcqU+qWrcWTUWMo20Xw
FoQhKgyIg/D2C6FGHa7na/NS6m6uhBU8mSSzrOZ/etIEgagjyXu1e62V1kZ/evQP
AIEbi2fH9G7BojEt19UOQWzua8qxFU2DG+zi+/JLLvR4Qks29FWmm7fYyLG90SBZ
UEpkbGnPj+IO1V6vhY10rULO2ZgzG3qFzhnAC/efBQ5rceKoelYPpESbGevHhbCQ
JSlHwe+t2LPD9wYW5gzlY222pZvj6DMx7pf8LrlMIm/B3HzdyIfn+fkpVL3xLzMI
sWAZ+PDMJSeaHdDaw556HDQBvqpH6QxN7YAY/kCauah6DXM+xGYRtnbMG00KwMIf
9VzG/GaPJIcPpxxJ0AcxPspOwpjsuvo62Rgz7eVljIL/42/kQdkfOQNN8/pWFxUd
En5LIpqOvw8++CVi2Zom8rHyJ90kC4PBMwmBprXVsvoL3Jv45tJeI97a4xZlCwYP
3z0aMBEY05limOGVsBk7tEem26J3uFqn7O0b15UhCyKQ4dWtyfQgJ3XTZMsJjp5o
Obhro8Hy1XcEukts6iYW9rOInJJUYg/1XqwaBfdeYqKvfvXkpjVkvK3wayA2nwQk
8Y6IrUmQhFmLc8tJlfPZ7eM8zizRLjQHqk3RAipVNjzo1Aay6LB9M4xHUF4G0QSD
30zaXBfaT0PmYlLCkCl3LgUtFJgrDnUBHha+sSYU0hWnKaCO0ZWSsdnWwSqI2Gyo
vhLfh9MyPDpUTJjA/J0H9Z+DvT1C2lnlI6ikmyw/tDzMGoeaVOXi/ZiqEpvOmbjJ
NPSBBOLVDcFppwqxIMpFyP4jnC+PNdzVb/6miggZNf9RyNVjEyxM1PSOxzPNzxGY
Tj+DozMGNXMJiFbv0TZW6B4OtNpRBPgUKtPHQ5MW8IJzx3kzscLz86uXQIAuvDiJ
WuEefZ0llP+AouVcicqwGEjbPIIM1mqLebgIIK+lpjkweujwzalXOzHnYjrzHAbX
O9YSVwz0ROron9X1Wqoxd1X6nymTV9yyaPmzyXywSCzdFJbl0m+g8L1ztIIChRUk
y9PYil1mBHBvn8AH+kXAqugRjZbs5X8C10wsG/+Tv0rB18Wmk+oztBjlZVuNcyyb
MTSBOz935CJJ5IK2Ya7TZLB6dLctPQnusNdJmw2IvW/fz3i1asbqEw7AsC+Q1D1w
IZjTmpGwTLvxuEsN0gjnqx9xyRFIS1uT1wKGtBUaeCo6QfS27LWjPScOb0LtZj6z
bJZ7sK6cSpyfnblxDQZ7VX+r2iz95Uy5397VTLFGy5310VV9dMeiUZuiF8YLcXJP
25ukkMs62Z0WOPWj4XwBpJWKlm1TfN0qEUKf6ycVBsR5SrVbvFxeCxDECidHwH7W
wFEmriWykaco26/xqcUBcF5F/Peooo+RDa9MjTU5jqY6ZN0nbpFW9NCfFnGSYv/S
uLdVvi8/CmCHu4k5B5YnuLLfdLkMjBdJ500bCt1ljOIqJYsQsGK2kNFdwNI8nMjg
cUGS6YR/a8odqPN6YcqgYPwBfYF0EA8F0mUsjBTp5pJCYr3x8pPoyMMv5EAbSA0l
lixB9nZTpZqr4km7+P/6xFlOlMagPHqk7hKTCbvGurDXM3u/XHQ9rI1G+lAwmL3J
Aour8mXTssA2tyZo1fu7Xasb61s8jCg+4VusM32V6M0D8eH4P+rIqj/TGQOC+Rnp
/4SdOZLsNk0O5U3Zp/JDgI4vgDLRPr7A11Lc6PBckuG9TwHxNvEeAKJOtXv+ZITU
HgiGqXsvTHq8jlcEYv5KB74dwDKMYjoMN6n6Hqc3cC+Uq/wimEJKRwJytKYc6Wa7
y+N7bYwE75T4E3iCpeagqNXUrOcSpAcBXL250AH21zdpGZjZxZCmRgtiBsKRdNBu
YUHs3iDMNWpDQKAXWI/vzvqdHhQfVCgErUEkoCbrgROyKesnQqQ7Q0XNi50Knqde
WNIEBDu4IpeTQ9CdNoLxP7mFNhb3iUjEy5wRJrn6XbPVrDkpVvTkj9QmC8rex//H
76EYPiY/WAFOJE6KdPRE2k8855sEAdCKbvRevZVLHKPQbLtsALLJYRxfeQjVJA36
mzhm+lql4kGUcrpXD8Z0LMMHbIk1Jw+0XcC7oicder/Yu3ASV8ZrDDzbXaEtoOVd
80LLHTR7eHZKr0nQ1WCpYWZNSQvD1gCuXaeX7TCMPPnU9Nc2ymeklDYcA8oWn/iV
vTrNl1dru6Ydm+4dlmASbq16bDnTf8CmRqSmvZ2Bbug8+/m+lzxwltMD15BDwLhp
8tu2jicY6JMNnZuY0x4s3eDcNJ7wf5bKf/tO9LOMSN6kY01DlFzu95IoXySy7N95
wgsZSSKY6NA4Y4Q95M+NIenob9ILcR7chE5v7PZ8ssOr9nXoaXIQ8ZIVmSLk8XLe
109CVvAhYqIE/YACIWDlgncS17N9NaVGt3Oc3XUPQKjauL5opQfTbBTmVx2r+tSp
ois7B8RD9aJNfTHKbtUcNVEgpPGXgt2mWDlHIeAyLtCi03j4jAIEm6A86XdaQQUk
BcF0hgOY2aCo32dqBMhInNETxOTnpyyJAoJ9ddtISJGTWk+iDBqjRgbhEYDlmDiB
Ua7pxpxxIaUDEciS3CLGs7QrPH5q+qWbi/7gb9iVw5idDz3pRqug1+U4c4ygjKut
kOsW5Ps9anNW3Zwd7+9VyqyCEtWpuSvZGoIy57zgTn/Al1FPGAxVWUYRtaYXSTSw
4+kTH9qGpusDQQH87VlhgFwnuV+oQVZ0YZNGcB4/VwOdKqtaJ0ABj40TyP5Mm0Yu
u1jzVWMCHsNZCMPOoa5qSI6MEE5nyRXCJ1eK7NW5NNYtCFhxCoZ9GkHivnkbi22K
AujeNcnvqxJQHXyR2+B/AFT3ndfPbjdIDlOmFomzoHyhB8XQh5IsJDqcaV/rbaNh
9owUz6wi3b7bU0mk28hKpzNdTuwYcv7gij/RwtDe3TYxDfievH9FTAu+VeY40PrY
aMvv74koavOxynfXcv1zP6GCffqKknmydrsYQUpyoie9dD/TqtT9S0KFQ+zT7BuV
oURKacQGyIMV0YroKsooZFJEhbUXUuuP/FmxurczRQHhBPDxzkcYcwyLu1PI3V4G
Z25f+m05OL4hYz5TYEtuAND1iz9HQ3kDQn5odYiWeZuhV3QZCwHcdXg8iOq5f29b
VBRElDa7rrdYKftSsijb+Tf74jjypi0UKI2tmUvn67JXRQmLMCQOEN4WxwNi2of7
67pnPAvZ5O076zVJwr4eI2Dmktj3XadATN6URkypB6v/7XKmkW/bA3TK7io53PoI
M6B+IyoGQbhHNOOJwcmfAfpiS4tuMM1rlVQAQ3OyZ4sGoU3zel/knwTWrhIcJ06h
Bl8yRpepzcWgAAmSK3jdHd7za52OIpwW8g1AKUCjXdEoulAOjj2NMQDV4Jt1Ktfn
BFWeXUa43eKlPpjI2Q3EK/a1jnMMN7K935VAWPUuh5P2UKpUovAPhAMnxWEkgoez
bnvKqZualcyUSgvNYwtu4vvzLET8qiI1XvZNkksD0ZQj43JcVNIPSW9oyulzhB3x
xMmZsHER/HmnHFUOH33XqI4sFBI0eHmOYi8RBqzi2GfZZREayqKP8Y9xDxCqoFoG
/ITtuQdVZA7CiDK6Aj8aLt55V6u1bDVHsMVWjl7gqIT9gXLda9XokkTj30TmDchf
mVQd33pdpDeuHlslD0yXge+txVU36X7OP6kSHLOyKkraHHsoXGnLzdgcCKxrV5fs
IHSs7d1V2pWrnujNLuoXlgsdEqC7f/+akLN34Li8vo+YHXk3gWNR5UHjuJrCqJ5h
ej76PHN/Iu/8S5ToMLfNQ86J0n/UfgnkSci+13YQ9J+Y1PZIblrQSjIlOe5EvZCz
PS6/LNUPsJW9QW579TFBBC5t9876ThiK2aaBwBzW51PYoczcpxkJJwaEwW5iRiSX
gzQ1KqSDQPfUXGp0aPGadEJLStFtir3Oj+XIoJr2mtKK+q+HqaAenetlGoL6tfSa
Te95nqgpr27+v0FdRm+76GuxAror3my9sU0o1cLNhO9woEJaviq5DlWYjCpCaFoU
uCc0/y1QnUbveji/bCrdqkVgum/GAah7lGlBoNaCFc6FQjaJtEDxp8scWASofc3k
dPYlgHUKdEmO8kzot71k/uDkbg5NV9vz+chyxzfA3luW9wc97k95bOgKswrIAV8t
1IHssTJktivzP51ngIGDK/eRQ+lDGu6CBpwgt887Cao2p8dyVOX32uiMgZ8PHsBo
EqhMHhge4reWjRmAFjktA3KkthXMOYjgZy3HXeOd6r4XMIcXI/3OBgkW3IXtpW0A
HGkoY8V0NWiKDqPJmixSd0QP4JINupvq3NsiLoj1RLj9V0GaOuWl0NtccC3M7ULD
Ifebdw3IBl18+eQno390fwYszmwWkQW2J5F/un0we5eA2SYEpht6fonUUw4ORq9G
GurVluFMpkHCiP9Hu1+SzJsbK7EzyNmcAIisRzOixRe4v17R7dDMCPcrR165f7GJ
Gfyes2lM72KPB6bNtKIuU2WzCzDXh//bE3JuDTPbPuO1Fh2T+F9Hvw1zZctfeYhP
l6Sx2FAifjnYrm+kgdA7iRpSnPK/msCuUYmXFuNBz0ZzVNmtYzBTeVVpesCiKq0S
xSQXNSPrLmV56XrjzGGNj31ZXbpfIlKtDZM7MEB/aMf2OPSTtDTkD5+2oWZsuW++
ikc65cF95fhPVB+pknSKFq22vbkzgaQ5bUmK4L4g95h5lZT1vlEEZTmcvpzoJFbq
LziERJW+Queo4Q9tcFiPa0z6EA7S6XmqDUuAPJZRmvAy+WgJByPByEbR6DL576Iu
RcIRIYkK12g3sxAOJ2oMTfVSrxJkGwnacR0OrznDylLzAPqtbAPB6d8NdbuqR3Jv
+HhlIw1Co70GiREyMOCAPLL+iV6gHyqmbB5pM3K1VXeT07YJl/tC4aDpKFyfnpSj
akBhSCYPYUXXqPrQ41+rkYBKXfzQovRMKcNFG3UpeujN+qFHkoXdXUvRj4GVkGqu
p1qRm9B6AUbDaN4dZg0bhXUQz0Stb0DFwTGvqXjGlPnQJQIOuv13zsO5XChCYIKP
mGjH/rWGNmrnyp7H0JVMyifyYDaVeUIzUdGPLDCr5dWjCTyFE/KaqT9tyuC4Pq5D
b+lg6wS7th2eYaLaQn2QzNOTUFdlQgJPZq1P9TXmppbdVtXgMLt70pRvdJoP0DCs
KGuOb7Cn9y3jylRhjdBU/kIrjXLiMWX5HqpY3SJNvJUwyIb9xhQR0A8PvuUaIADx
OZRXN4cR3HwDWEpFSUyQbx9A/qxo3U8fRuGhR0AxkFMyphwkPzuPf5dSBVxPCZV0
Uo9Q8o0GpWZwSMtbbmRwfzzfqUqW+1YKsfWsZjJB1aBG83Jw+GhBingeBCbFen7E
ih44aXmYs+fweGGPR/mUDN+GXQ2cViD3V7npJqATpzc9wpQqgXSofQOUUmUSTs9k
jxyL8B03+fUNyu7ZA5gqu6LGU+Pbk/C794U/UoJj9iy9RLB0XJQWozNzLLiLUBpC
r6Up9D0/a+nVxXOLxd+qc6+Alge/iWU2UeIoa199Y64vQcIPiqL/zgCeTK/QJe0E
gEugEi7IAZ4FO6jZQu9u1lDzB/PbpZBcX79uAysboTOLIhF/jefJZBDZBBaeMQRn
xwzcdAmFOAcoJsdWqnvrQVsH96bX5UIxpdr7TrXVoFDJcXpu5CSwTwcmTK2dIrGM
EOLwm1jL9o7/nC3HzdRTJXqHkxTMYCL5MAjOzVkzHMUxv8t6oVm1rdUNs1PYWgps
4kEHVVLj6PwuJgleri/P/pmymvS7Na887WS7n1YHaMcMxCbi6Kf4fUtXJTjefQ/W
p/2Dy7k3872nsQVsJdimKnL0abi2JMRcq//TNPZavsbgzyAHzbmZihon8E4v91QG
uIYBOpyJdCK1KsliQt1IQdSyct8g47PN5vcHg6+PmFdfXCiK+wtGU/hbHLnn/8Z/
naQ6IFojlGQ9t298ZeyHDEFrPsJdcTZ2q3Eo1MAHrR/YaCDcfpovb6n7rmR6NeNq
vhmKNYC/YEl9UtkTh8AkpVf0AlxIec9vjNDNCxaA5eVIPXI7w5vt4pFFvP8RYbPl
RiT6CS90fa7HyI9AJnCr57vuzxHs89IN5bM60FIDlERiXxLGrdtc724M0lKWegiQ
UzIB76ZfqOc6cMUDKRcqCTL2iSBq94FLP1FUm0cOZqE8QjS1Tui8FtFTIiyzYuIJ
8j8nsH5Xz/JDYuOARE+jhumZ+jWOWd8B31QPYVfFJN1XjP9FlXR24PdKGvIQukNj
QNY4AsgwFYv8AA8WMVCQ7tSdsNoTUa/H+js6mlNRqMfDOeCrU9cM2rSWsHQscDnw
yiQTkH2b0F8K2nZRv7oI0UJr6JvxUxL/jI05fsBnhY6Gq0LMhMI5BSWpdE6Ns9S3
xd4DsYnHS8axKy+v9kWt/nyFMK9SCtDM/D9K7Am8RGEcVw4D/ttqUNsqwrMWEFIS
AzpP6+ovwv1ce2nLzTA7cCfiWyQqW2dDfascn61BR3bqknNas2lmce/XKkaIGSDT
CIjjqIZcrlYpcgrkS5dxmkTxB5Nto/3wZUve3GD3mG1+cO/dVoIPnp09vuSNR2tQ
nTflBiG/PMcZjUAPNkZh1q4YwDHdORtdXlU+DqQIy+j/61BE7yEScqvLFqbhxkSC
MHTY9Y2l5HW8cC0xbKvDyKUzsklvjwUo3tL5Ad3aAk56vgpD/ovGr0w8osBWzGzy
NuFthh2hJiAU0ardYz+NbK05O2wAmQ9WlIaBo42fu9kMbnhJwRnayl8aFcBhkTsF
T36ZA/ug3UhP5Aeay4GTOFeI5YDoA5EPnfgSbqguR/BpIBd6e/Pbi/oLTISfe1GB
fMMxTJQSvNR5smXNlghYUbro+RCim0EbhtwjRMDbggBVYFAKZEDdfScUJcVO4WLF
mB7a1Q3ODuxl+6PchBjXhTcG2EG94v9HmqXWtVNtiEyQ96uxgmavsU9TUFHbpOqo
kNQ589L2FQHKr8hxZMs36Z8ZkdxeZNwgggs0ILSy2tXatQRFeQSQv4e4rk0/RntA
cP0GM+AnxlwWpRF4pOJPfxBtOpX7RrSInU/o7YGrGvXDXFiQz7/v1qKjdhuvFuMm
NdyALuiMfNMzh6WVg65ne0UrGvyF86OTBRK0NIIe2dwB8CYWWatdximh5WpRcL38
CDJnLWWgB48Ip3YK7Ib8YicJwSRoG5fbmBW9KG9JfPIdOHBdrgGi9b7VcG+0oX8c
7UN4ZTiO1srJxeL4hHO4fyV6FaGhWPWgQWFr2Y3IGG9ljOUN33qxPLnHUBdf27kv
whPjz7wQx37wByPgHdDaETcX64GiIOwemWC1BJBaCHiqCXIyk9o11+L5YCX5BQP/
8TL664iEFbnhBeOs/A+ecjC8oMU5bg6JVZohUYkYwoVeIJToAfphcgtXjCgy5z1K
XYe6U+0yn1QEQlvujqgZeODR8IdMJ8tScU18yRy/SQjfddEXdFHsIoZvqT8/w+CY
GospIGk8dEYk6pkr2Wav/QD26czSX4gmoyNfB81lvzLmLKsYQZR/eDcaVc/QYyzB
luYwZl34Dbf3TsVWMBLmZnwQcdYV672W7LLsLIQZpqErWz/nqeCbfwmjpTZECseR
8IBMTKNRdRQ6AtGvj1A0bTSTTEBKvbZ0VSWe5gIiyAfDfAC7ukHg3N3FUxST2neH
DMXIJ5EljVlkIqTfowYbn9/8DrhPefparpuQWTukfRMqthXrj+bPwc3ZSJ3rq2QZ
6EPDHFRfMRu9NZ63XJm/mRS7rL82gMjLvxbvySMc/kPFtl8kN5vz6pnzkbswx9xk
Y9TkvgG/5RSxyI42zDjcrqVLyQzBOF4CzASd26YDtq2JXqlpJ0/s/FnfJD7d5GZd
ZYDtnCQr+TQviwc8XT8TB8aNTkgjlDmYqAy7Ny/alLY8bnJPpDUZoTDvgtvsh163
WpVW8iIKaD2BDXlWBEy59sO9fxPJ7iursWSZCiYb3gVncGoVw9mq1IKvWJhfkXkb
p8zxvCJ3W5KQtdw7r7yNL3fV87KXTqaHPKCbHII81UVd7l1JB+V8n0l3hK5eYp2d
xLaPTN1BbUSKzlfwTRQITPlsWSyd/ebNYQ5OmOgmjgnE5zy6I++MzWHLFs/nBVVP
0iBok2PFbmXWLA7LsLuwvRvOxq0DtKLPPv9j2KxSwdbbWE45Zf70/I0ZXMmFkPDV
2sVFMnoCefss9Q+5OhASR1opAz58puSpDkQpDgKE28MfR5hVQ5ZrcrBiIE6CiBc0
y7SMRi4z1qI3kvrrDqDp2ujrRbr/ih+f4EWiIBqgryX99lwl5FF8y1LFJLYgxpjZ
tBIufb0xXBp1BAPDHUkuwiKPwi5vkJ+yU6J+HEIvnzA/LvxneTlQKRai8Tz55pOX
0AmeAVo3/2MGNwnaWp0tGIDp3+Vo2WDrgLF6tsZ3N8V7liOE+qT1F5OjCB/3YsZG
1Mj6Fi/9wcedGDzOZ/JTqHinSuk7ciKXP9PGikmKy5kvdhvXERQJgExCRMPdxyb6
xparxho0x7dDBQhYF86ljPcUZnlN+995o8sAf8d99G12aMszlVHLbwpTzQZ2pg1x
l6f+IajMQhDehRnPF+P4ENLvro8jdlq3SSBFqnag/x+7yScBCC/ogSr9mHnjiUAR
CGySuTla7fH//7KyoGtb4RAOE5PlBD98ba9ZibPjuUw67l3NPeYbARsFc0TjkVLa
OjUY5PSC8cv4H9NCCaU6cI63kkrwZXFxgmtIzihlROM2oXMahwtLvR//1GdRHHtx
OXncBs3ryzUwWb8NDz7rzzx7fm/4v233L8rYPQp2JZWlfuWqo4tNwbOXXvdIm3O1
QxBaCUoEBoUMBnxhwUOQioiE3Lf6nFKuhRNRi4JLvHKKTiUdcFpS52JD2UgWFmkL
44It/CTq567irIXi5eVypKNhM2m51EHQqkmPWYZEw/iz0NtJlCOzhVlYOUV3CEL9
mJ6iLOR4h8R7ROcXkD8qvh0NkuHa8FgfQ+v7wrfY2CUM+dJpXmjpKRBuC0IHlUsP
iV4tsFWDFGwBb0pPS0IiwiZN3FtzjFl8xs5UzXimGLZy1AkUZU9eGt8Dafms7Dpo
RmYty7edDc7g7FoTmWS/GvoY6P4Ch0hsmJxPHl/+t3oBYtTKPnaptyVTY03bVCqQ
dIXks6BPGsmALiAii6V0btohoqAesOOqF14ymo2Y2emjwwXFuMPV1SolQ4PGd2he
E/s0CBrdNug1GnMfd260Z1QPQdbR6TyfmJj3JsJOkvf1Yjd905eBM3WCd8Jo4iVG
nmqP4/ozojm8DS8wdquh3+dV46ZfpOOSSLe/dn4+LOleEu/sC1/jO9F9DO/ZZ2Tz
i0RL0eB8AZ6A8mq1pe66pSQ/gGAl5RgqZlCcsZU7H5XVJXMzSLTmGkAI+m679QJM
XhZavJcZ7POhreqvsnlIEP3XT5C/MkAFPrZWSQXRIimpnEWEK1f+BtEhUCmtrbyJ
4EfPoBMSTzbQ4vkiEUJmTP2/GVFfhNjRSWLoqgi0Uf0dz4lzmgzDeTUqxd/ZjpmU
v5ampL42BaM7StcCKXcWjCHJENlzJcAH+q9KAKB17a9YBvMAaZUfQpvX4E7sO9oi
qvgZOqA4DKiKbOGjnkSAZS80haGpXw0wzfqDD2uyvlU7HP1iPPi0TlinLHJWJTs5
COjcilQqB6TKfa8f4b7xCz9KYGj07GQryJqDZdee0aKYzdr/RFL9ZbQMimy0GJtz
YPK7edsUq8UY8wwUsDlkL4+zDPxdT3emlMA3JzhwwWD3B/17qG6Z1RZdKPKcuxrT
FbUinyX3uWwTWlsWWWqQ6nqvkeqQoEqGz+/jMKZgY4eJxorCQl5yec+1CL03Kic/
YFFv3dFAWN19o/r46hVXB5h+3qaEMko7VgNg1PKjRN+63eXjOfQomKQlqKbOcR+n
q9OiwOH+ty10WzmkJy3RWLr+ZJ12BGggV3/oXlh9ZTzLlqXLYWTf+CrFL6qgLy9a
iW1HjZemOfMRoF3GbG96CLl7Onu/5jrMZ7XFHXTY7wH0hPSgj74/2fVi9Y6RQ57H
37B7sP7J1YPOqNBZhMkAuPweADtVxOEfI0o3IPYFq5jVWsbZiO5GamlNz0lC68EN
D+ynHwqVACdpiQYa5D0JzqAynO/84uMm7dOPf0jX0/t0NFblhIhctbV3aRNW1NKZ
xFMcoODDbLVMyqEGgAI275/U5JtEtuKMSEw/f9iF9VeyIZNyEQGLJJ3PhXFm/H6D
UThmRyrJQEx5+FjA7GVskp/IZu2lV2qTdnVHtrvgXbKOCzW7HxP8Zdg6EHGn4sDf
JECLZwqelJ0lu7n1zm+qmmVoPsIquZx5b/9gl4BjoW754mZqCfusBk7IYKaMpVst
WFlLvd//gpRsWgKQkvFof0hdttNSjddMLuwtIYc56EWD3OAkDpofYS+c0Aey0ita
o0/9cIoODVOg5owTD4Nw2QrEhtEFq4XnEowrrw9qGYWW7nsmWSigZ4/lZLSSeIDn
UhhxFE14lzr5kEtSXA0l+47c9hT4BYiqCfK8R25+fNK/V7i1ML4uxO3hTS/gIFml
yLS32rLupDRqEbG9xA9We5ATIXpTIeovap/pd2OsyjVhEV88zaducDgJX9uZMTMe
BRvmQPqhdB5PlugIPx4lVAbmfINcEwHtVUyJaxswfrLJEGloZULhO1tTUpYTKaKS
z45GHhrj8BspGErvZ623j/pxNsOWjbqTn4kEczrvcSzuB91UCqNIK1dCCGaVnlh0
sFlO9tviK0PoDWbQdb6ubcARzNu3bhNOFOI+U2k6zRGo2oX+8WaVvMQQ0ruSPTOD
zYwzFxVnAJDNRBm3AjDaekP/S8OlY1LUrMpcrBPHPoHlAUYOzuqPwh4YH4GxleER
mMfhk1QBy9jSGycL8tL3NiBzec8brchKX7paaQlV5N+S+dVuJFCwVBq/SlhcCkce
qe6zeABI7AdYiXYgluq+LtDqRCz1tnEscWEMbC9Tkl1s9zGVu/LGnJS+QJP3oDnY
jcvJxaa24JchUwDSZoao41ofqJ8Ku1Ng9guIVNq/24nu6J0AxWoX+iDGUDE2D1Vp
+d22z+2eK8Hdiyoc2sUEDyrbpYe92hdkKmRcSpHHUwFsdVm0HH+DsOYiY4+DBgeQ
UIKYNdJRD74w7zWrbBCaFdbZakVJ8/7DE7jseElAtlF0YS3d38f8yUYLJVNiqSLF
7AE6pe+dCZ6Q8n0kXxg1+DS0LQ/Bn3AIOwD0U2pmrUWTStRb03xkOf6wieqffWcH
dYzKzfqsBLW9B09gakxZiStZgNc7aayaGihNZvllfU8PVVUqZiruXmtlHhWvMku4
kCja+0jpWWRp6+a88QuhBbpRYPsiDIf7DtInr5WFkSbNShg8g7E9EuVPzNg0iJ+2
N1U669HRZ7g9Lh0ItO7kplRdNrbPvsuMbxzKzZ+4hQCMr0cZrOr/4l3OfzVgTc3B
TevTbG9BE22rfPZgk2ywRyfzcwbnCgechCnW0J32KqvEBKwn7MHj7ze3GQnhKrve
IRpNY3WMiBOXV+osFHr2l6sd3TmZc1zUpFCuLSDDqWLn27RkUpl0QTiChGEA65Bc
Iw9F55/4M3CCD26BbVJMmtZpsXlGk/k7lxGUmQoxbprPNf+7Uhwr2ogd7XP6IF6v
9b5KDIEGz7YFztC5W6pobRFrXqj9ryd85m++KMNBlSoB12dYzx0+FNNnKm0J7mOI
L7DE1ajWwikLbmfoukEyS9VwrOs5imRfSLX6f5Fkp16AhXoyPcefUuhE+tpbbiy8
IqgsltC6r4RIlmM0xt0tzkkUHo/qaAE3LhZ0HMlcluCANbemLNQGmCwmaCg/X/nf
sJxdWIdOZOR0ga3+V4I2xvvU6gPGVIlzZm9grwKpb5wfLZ7jPP+ivseNI67g8K9+
2aEFiHuTALZsfKkbw7f3rqvUtYpmU9bFsRI+OdSUDELD7Fv7Xd+tMM8sV/8bp1h9
G4VJH83bPUmbuivRMUZcuZXxg16BQmrsJ8xguRgWwWeHZS7M5Ydm60WnHxOWgzQa
+SR5IRoCmbaztpiE3WrZYcxO+xInSrNuoSTpeg490LVK+RtM1V7BwTrfxoEvPw6l
0bA/pZizjj7Po++gQlIp1z8bi8c3R1INpj3yZ7fo/GRk8quN9sBNnh0XJm9KcT7M
sjnqiOxMVr9+j6iES0t0eVjL83XcSxtrVIvvL0h6ns0PJrZiz6RZdPVkPgZo/N6l
LfjPR6UD32FkNWzaAcBRMw/f/BwoJzqa8EeYQi7lHj607XbUcK/X3gdRKZP2mRF6
BOGZdfMiR4yJGCe+OiqQIHTje04dXanZ5cME2hlA2vwkaUAGKiX3P3zDUmpmJrep
WDTnkzCIrDgc3TPjO8JsYVc70fFAUDmklg3BYO7+KKIigEuVofYzuU7d613keuUp
9RMq9yxRQE/ESIQDlAZW6Ic7bDZ6Flss8KphyAim0ZYHxIWjO2VwN778haCOQO0U
7H1WWzWp7YopxmJwCkozOjULyxjwH3V/hbiun4sCOwblC4kwqhpv05kAEwU9aOma
daiM7lvSMVEIeRmqqUEz4atBvBbeS8cWzUw/E5DSCrUkUiHRA+5YhogI/dq/iUyO
UcjlZS0+gixyvsJT/wBDDe31XfqlS4YqyIt1B+cNf/1prmsdj05Ae70TBz9WjHix
s/kjUivCgKQ87pIno/EFZiAT/ameWrRZh73nTQj5hXAFC7JVRw+YdQz+XHkCPVcj
0/HuyVzaJTJxxNRf4wxcfTklO6OhDMP7DVz5X120dCgkxwakp5WMDNHE/GxxBg6y
cMY5zYniR44Cv0FMu8s+QdT0GPTW16gugwu46VkcW5avV8g9p7FBTRdUN0uFNdtX
nxA6sfMNsXJPR15gFCumpMkBSCD4/yvwV9e0VwNXgBLfTUvb52l7PjmY/4omcDRt
RU2IC/jx2oZ0H8oXAcYndGuFO1HTDJN4GzML8h0s+AWO6TiKWrNtMO/cJRGUPhNE
FkwJJUrgzE4rf9FDVTVS2rjIbsqTiz5VJKU5UfGA4VN/MmBd42YHn4T+BeUiNPOV
VrGIc/sCBdk4z4UMOfpU1NFPhau4lt8u/lbMwiQvKuTRnSd3LWVf5lEgiw75TVLw
ogJ+11Mo4hK5tOBBdX2PEZbav+5o0SJx5Z1uMJOyG+XsxKkrc710PXgloG01HtDc
yzBAaING0WEGsvDKGGbXFoeAVRmMUq56C3U4u9ffLLGQ03PJ6XQOCQ6JW1pgplBQ
6EHLyzO1F2oPfdNy/ezR29lPZ6SdgSRW+GDU5U4CInRu8vB7AbE5Lo9NtSK2Kl2e
ss7ALRFr3uoG81GHbTRPzdoiis8/fP8FAbQw6AXr8woG25b9ykVS71Zduf1tI+CJ
Ox2mzonZ2WWLafgDwuFrKsoWXXIlzNiRE4EwtQV35ZNhu+MwdQor+zpIvC1cbf/j
zE6Ay5AQj92BX8OXqIO0y4JTuLJ5hfWGxZqneJ9/jSw5g6/YULg29aVTKQnbzR/v
UhfXeiTGqGWg4+tMijp6MOpu3J7zxVgxveJ5Dodbq5CkyW+ceqbfsxmAChrWK76/
9yloQVb1LTlWb09DeJ3+A9/zppUzkB3T1PermpMUQDlJmu1DGXG2uDezJZRyoIVq
wjVZC6q6qDwE+KcnnWuLlDTKkYVw44YQ0VCbkZnRyitEH9Gea93V3hOU5XOaZGtF
obnVks7CL9NCCIjXw6hOdKEihsUauo+Pu8XVPRcmrjrUBPNCBrHZaJh5aLtlVXtx
Pf6w/4JIY+4Xgg95o3e7ZvdfoJJH+7IVejEjTUAQTaTM39jkicCfMCQR4sYN3yS0
sl9qATV0P8ztz/IAIwYOKy0Tn8/k5t15R67X64PuH8OkW2UE8y8GMANmYkEylGSd
hRrtivUPsJhD0cu2H8jo8uVu/teU62SxYoPoq6D+3o33YmKaPX3yEP425ajNeoIG
bu+aJe9qmrEnPmylucs2VeiVfF4egDZZs+v8uz7uRxAtI7ieQt1oE3lODPD25HFW
uAyKtuzAfFMKOCrmD66c7HI44m+ZCFoxPcKTDubfwMVl6fZKYg2JrnhI+5/63B84
ZNjfHhyFyjgRcqTdcVhIDX/iaBE16m781BoHepYo+z4FaWFOKhkUVWW7jF3gLylR
SQVZKe4+ShXGe3K9bfvmWpDkSBGIcqd1Mf6pTF6rJWMPqHcSyiOJ3IpdjrCoMc0+
TXVtPVrxBXyRunwP6PMka6cGWdn50tt8dQHPbBVjMVaAwNyxC+kgkH4tjLJwC88R
5GOwK2g93c3ZiU/PLpczRKYx7TspMh5Cl7UKT3XdzulIx9EpvW0LQG8Ei4cl9Oh4
5dDJBakiRS4jLHlLMVPusu4dQSQ3S4/4HOb+OudtKsdQMEgFy+ktoCRkBJs+NOkh
cCN5rBSuLXVS4b7cmJoS0RMLnF/96s5b7v0ty/nbV8zVqY2WAkgPm8AkvaP1KI+D
+SfRD3dSguibTxF2ujZTH+WYL4z+kVH8jhPFJso+f7UUuKJK8Zg+LcWQAZD9GrGK
FaIu0ecGsaUIUet2cAslgXJuhoTvAQqbSyn6kTZQQo9nRS2Z5R8AV5fn8zLo5SqQ
u+7nMkeAHiH+Xo8oW9BDy4TEGvXeuFnW/6tsXRy7SLbAwm0z+ydFIHvrtv9mICbK
WpDqIkSdIPc860bzIe+tiWCWWDZd3E6xLYs2vB0BLIIedQK41DxD5wRX78OodFeE
MwurSdx+LmDFCocW7IAhfm3uBDeLun18aKnGUJsHD33WMnt7Fbf+ciWqfXck89V5
Dl3HcCihnriyZe3Htp2ZN1pJKyrFsglFmTdd+6U+TMt1vVuPsR3h2jkLHt7LF5sh
rbpCZoNMG5A7OwroaZgltt4+ROtAkUtyBGyfGDT9YYAEXFD13LUvqkDwV0CfJcPl
gO1zEpBJ0yrX6FCIKdydzk8RVUPq631G6C64pSb7YC/ll7aGjkbDba+KpICR8hHy
PuzhL5CR7YrCiX99Tkrn6Xan+VSZLadpq0uBMMOJGblrQ8eObW5Ql9qc47MouJIw
F84kcWWXKlv4clxPt48ZpE3EWRUfYktdIkNVS0FLJzejOj+lDw6RywRLeKdp5F8o
dfoMc1fnzZXQBVQDFQ2wSW5ksv8NWPgr683skmck5rgejWcT93IRHQOJt0n1PJ4a
lDQ7dVIvExoR/diEpINJwXc+IpYCb1XiJIKg4ZZLI++Ad3kBL1UVUxmJgZCvvipu
82Coeto4/RYEQ5mCAgPp1Y7FoRMOushOw928Prtn89QmwWFavP1oOZv0fxaGZqsn
wSd8s2+0XDf11araLtk6y0a5/V6qnI2hJ04smUnnA3LaYjPGWMaOS5AzIEoFWR14
BVtLWJRbRGDN8c7a78VzJ1NUgpKMsYB0Eufq+4m7R02W6vyUDKX2J29SPvX+Ll9w
hDDw1OdJ1NU716BNwdkWvCCaJ5E2X3EvIGsT8ciqwWqSn/aMqKA+Ft0ljipJG9kq
GfkILO2XD1T1YhcMnZnydD5fk6q9u0EzMnxrEd5XyQmu5HHPFGPumyVgso/5RJnW
KTlP+tCizH435mHzXvf6nXz+gCPBt2lo4TGlGAxyjz2EtP52+bj5xofGiYbImoPG
UV8pVTsaYdnx5wt+SK5WpR+r19XKbrwQsgq1KfSbHDayfJVICW58nOV9WIdNYnsE
/yzOwkr6XqEut5xoH4h1Ib4Muk839S6Y7wGJhvZ1G3y5fD/Hw1aXng+kzq9ALYq2
CJpxLxzLyQHf7EeTwnZ4f1gJAHHcXqt2CnWXXaeFS7SwCS2RkW+hPASWH0q9ibWx
YUdntJ201LRnpHsVt5vxDmioo/kSchvSjjE19yCVb9OY8lwgAUQS0DJf2B+Hkgab
2sZ2Xtiqw5HEUB/52w8XWKluNCuwEb1xVoOn5kda02IuIcSJngMAYsoP5tLDVHPM
1B2mK1mF6AYSPFx3CJtaddTFhvMSp4ROodOHTiwQMiLNX0lyxJmJc4U2tTJaDGAG
RKyqZ589iyn/kJDi0SLfznzaGgy6Y8O7anKXGAVqanbMZsUw5YFqHkCyBvsrH5QZ
l11yGP21jt4DLeC3NTyi7/Vht7TvaxQ/i+Ti9YAQ1yt/urd+0sfAE/KX38XWaA1s
omKX1NwpywIbbO7hKMUF/L8wiOw6aXWBLq+CbGAaQDNkdG3AmuisYTAn9bntMwaB
+RKfPAimQf3JXsxaQRg+X8SQnN+O8O6+EcmZp+/C6yUvsk4A8LMTJC3OmFHl9Moa
tQOE1X+EzqYF7mPkRtXq8S1tDFypAnTKPHu7vOyyVoMzwXxc2bhgikY2asmvmZdW
1dtdvjIwkd+JAtU058sgdcLo7K4QGQpHYvfBWq0pJ9tNuamA9cmWryCYYokzQsKp
ufPOE4fzyTiBFl/AKzjwKJ2m7VO5/Mr/4mKeW16SkM4r1HwvdOt+9sqL1t/4+i0c
DP28RV4U/PXe1T98mZ5i0emGjhZ2cSSHuF59MQn7IB8+uN+kDLUBdk6GxRwnGAEK
2oJmkbPdmzeFsMfBa25wV9+Bh2VGKuaFM2P1tUd5ky0+gGFmvdncC/YgL9MusMCU
Cv5TcHZ8N5WeXSLbC+5JYITJB6JAlcaAh6q0RZExyiVtVmSf0JGbDAhKA7xymuF6
Kdml8hR7FIRzGpo34L9uGM13wwTw7Qu0eQSBUjKa/LO3mbfL9YUKkxemLX0oiwxv
+DfVAc0jJpy8ny/ZESbv7r2MvwovL5JEwYY1hqr0oqIQKDi7rA3RfDwUqPU6RUiy
Fg8u0OvRj6cYKcl+H6eFp34UWxWiDeYCvT9vzACAEb9A5+pEQVAbW1mdc9t7ysfn
z17tb/K36VmfOFnie1pFRxQYV/KSKSVaoDPnypcPFpCLn60IhWPYh5LhtJL2sc/d
j0vpx3HThKF4OvNXskLFIRIgtmgO9EImz/lRdcH5qIXKc8mue8iO5+1T/IxO5OaN
5C6Fs6fQhNRdJbiFdRZRxU1ckA2Vvu3+fQ+3rKKV5M41QvjxytRrOrYVy6Suj0Jn
vDp9KOYZldZy+/MJ/qsO65WnMbjLIjnPmuXB7lz+F+58ebm7kJSQKlKLLWIiSNtB
QRJp1/u3hV7B17rskEHT8aGsJOdtB+KbFNyJcra6oCTuBC2Z5IPirAtgLUc4Qe4j
iE4XlLWRE+Lwq+uXiaoyV+qwtoftXUPNTSoPbvmpew5xK9f6Iybcd50vWAMxfcQ8
KD435AZR9o9HcCqMPWGcba8aFHbbreq/C/7evT6ATdCqyYqRUP7YJEUV096NVXQo
a4Z+ZiM6rNHBk+g3x2/f/5r73sGkVERExbBBGpgj1YHsVcaWD7lVqwf6L2sLzcbr
uotvIvucA/IiYp+SecvXpdxRN/cmnl/QPoFVadcGtiAF/2xZ/0vAQy+yPpnD3nRt
BmiAVUoqwUHM+VNYWrBMXh9t7BrXbL0XWN3EFRryOSfRDs6T2EMzXg9bB6NM/UVF
4k0J5aGU1jGsbNnZWsaL/oUbAcs6UAW9WQhGPCS5ue+bgIePJ+f91ffNKlIQiics
rTpJ3Zo5tCQe+RBphRGZ/Ma98632JIEY+U+9yzbz+M4BYUnLLjC7Dh6sZpTdeBsw
d8zx/13uuLeqO240O6ZQpJHH438pt65XB6MV9/dmXZ0GA3kV3FumdjIlUVIzEl7j
br8kcx+1oNpmcqaJ7CWhPPWGKlBljhj5lb1GaEzRVW/05Ij3ANPmAhZCwypPRFqz
WqZJgPN1NchAXxSSP/36979H1+OWv+knXqUHvsthE8I7cKrATusWL3oXeaajv99i
u0FMwTpLdmDN555PB8s2Lj8rRoZ81Ctjsgd6hizojNQ2KhSuPYu3RqC5YomlPOXO
fneq6wh5x4uTQnsqwyOhrVL7wGLdu3iBmj0ZE7mW5cJlozECl0A0zmnoAGY2bboJ
HNg3LCALnk9Yi5PpJjDQ1BKGhUY0eToxhOLx2WQU7iLPcd6N3WLlA1IPHS7gn7QP
9cmreRjL+VwdSNOnHaxr6LxWQScDzqK7vBBTyblW7Rvv1246idRVOXMPmXH0A++9
m7tXJPGALwRwpRejPGkM+j21NQ7VYcsFmhz725JRWjdhxA1mlq+vbnuKe3h+W93W
e6IKvm4vxkDKCFKbRNh46CRPZaQCGh8JQWm6syM8MsvXVpuCkWZOTVX+8X1rPQCq
Z5p2IzE9i278URBAQGmn2mfAYlA5MABff6Ay/Z9rC0jZOkJvWZjUB6dfsQDaZfja
8BAdqlyOmyhQdNZEYYcRPASew98BSGG8+lHVtlD9+opsju4zaPfoRQ7iRKx2T9V6
EYV+cYvTSHqKHTbnVe5Uk+huHugl9VdlaDg9gLttXK1mxUHaSt5lyPP4+OvnAMgs
hKM0HIViR9n0akWa+ZBinaGlTBzDdWL7M5B2/XIjNtKrSXiZUPKdwm7tOVHQokpc
jwnsTgmbdgzm7Hm7OxYDXO1s8iQOQpEUjsE29BvBXtz+YZV8DuD1pVi34l2nX9TN
SZh9p+MaJqafCHPm4OQL4nPrRviNKCTuRHrevIH49szOYy4Rwlz7I9y3j8d8YoXT
0gmOulFiymVS54dq2djR+kYjJH91wMtLz8yDxAkuObJMA9xE79uDXu9zIRCCrMhF
bUm0I3dWoDIlWdCdnhBOo3punQD/pqtVsuu3lypPJYjnRRjMqE/Jn373iv0mTHxk
0iPMo0CtkGcsFaD5kg6Yv2TGjYm+BpyW79rRCkxys2icc80Udz+F8HA7f/yD39f2
vFjypqgNReD8RRS9SXkspmhnIqg8RlhkrqVg0NaXWRMmXJ2f5wVyVUVJUV1wi/7J
rlfT6ehCFwFn+JxPIvfPbGev5lhXXToUEXuyzOqukqxz+oDT8aaRvdr5x483tNhO
TRu7enTSvOxSHvcxy1oi42ublUiGGxNZT0MJfQXoxfgLTxltmnOqgDJBTq5N3bQq
k3V9steeW+nO3VVXo2OMWvROpZrYJF2eJQZTBFqnuroomXRE3H6kfw0IagvPCHXO
QTsPmbUV6msZ5VjzGJ0M8Z9BA8FLAevjyNcghjq3eVc5kNn5c0eIymKi4MsMmles
b4AiH0w6/vgW6Y994FJVRaeLcysdeP7dPLhv+SJ7BhTHBDxllWqkuSRaWrlqAjck
iT6cEKnKXUvfwxw9Og8usJkvwwU3vXeSdupuwCCH3MWXBKgEKkJr+9o9ZnaEa/d6
ez0U7FLrtB3E+XNOZTjAktjqECEoGJI0w+H/womh53HHJ8ic12aXlPyWJYS9T89f
T0gC1cuKTeQB40d6LwiAB7n2N8xF85D5UTOFhhN1TvP0GNLw1kIADNJVNade0M1X
iJZbHvvfEkayWof9j8uJ5bHh00U51W+MZPjdRMsq/KcfiBxmd/HZHpc9WOTU421V
7BZdh8lXRgN1qMLoadsQEO446tFZxdlvNNSXUxlho3qIHVKrYiBiByl1MnXcgDAv
eC5rrEqTA1pFxHdrHT0qN4JkihXqM0NxtbXZQvq1jcwt1vJFDHzGSwQscAzDOfH+
p3x3llZxS3F/x1Uwtrmfn+jauAezXnvVHNAtn8E0QcXbbSz5jpO5ROukDtdq5LnD
GVjMJnyFr6Fpdxmu07Fl5LnKggf3vlUdxNBybU8qYfB6FIe9mzoJrJF8dvfi4IOe
qhBtf5JJ/Hpk1Ouk/OuY7VJuMFHuifPcj2+C8yGCyDKPjS8Kd+9j9E2lJ5eTCmDc
jh/8a7qYssqrAw4FPZugzIsVg6z3qi0m8g7vhi7spT8KKqcCnTXXfpAHw4Jn8ENH
6qhiPS8m4kQ3kvD1gy3gar8nGTCgioxpBaYVnIGGouTpTriWXqPtlyaAu9Gt4cvO
qdiaI84/gkJwdRATvYmcrzgel4K0LzlRYx79Zjo/s0tsaJVM2oEVBNh3+tjMLOwk
9j/CAjovh7/ELT5yMVxWdeE0XEu+2uaXVstONWaiyKdf60ocYv8FE9Xq+o2L0Bph
ctyo3599BlJePN3qdbWNW5/3lXNf9BEmGG6EG15w2cNYHStHFhhTJcYSscFn9TBG
UvA2qcF4UpzteJ+bz+SnbLsT6whsVnioXywrVyzkhpR3JHQEJH89sOb/uoNxy+l/
u9O6JY+9rOjRtaiIn1InMpaVaq5MUWe94s8QKEMjuMCKK1KfsxDAltzJ4ebEoykt
WSgP+ujm2T/Yjh77Po1m4xedAdBOWXofOsHkNMj2VmyGjWF0dxqrc/FOAK7348d9
HOAzmxhguUHMADF4sn2sKUqVdBIwwZMNGShizEUg9FXKAefCDfO5KKoehowvQ6KG
uPFe8zX1AFcKErr9H957WnWAYkRO6/oeW60cwaCPcTSI5SkgEfbC9v9wuB8HReAZ
T6uCWqVW9ire9Fmj6ewC798+1Fhr/MIgVmclUxwgOYroLTR+4xvjGvutPhCHNLDf
Her/d659EtEby2WOOHikorDxBDc2WXBzt1YnVfMIaGaJCZcpkxKwpQcj1CwGOZkU
x9Eh9HNU0T+dWT9V9CgNufY6ES4F9VgoZFcRTzC8micsc8RbmN9pDXHZaokyuMmA
Ujxgk5eYH9YKN60ZO2K824OnOzi+sZ0RlYsnNdt62Qu1gnNYPhrpDvsRqXI0QhBG
U+Cp70NrCtZ+8/YyHDCPa/VfBeh9C6JxvSEK3XtI7+rkV7m5Q1RS0bw7WTP5AaAl
8G24rF3ujzWJee1Yf7WTns58csXsjSAXe+91ApsxOvVQotQM0t1LGptL6kJjth+0
NmbkGJEBvwoZB9mP2cPcEA9LI6C8zyhIeo776gsGTfyoq1+i0tCXB1iwQA99J6ui
3Yyb6z8H277dLHmLTM/fJJLg29Kg6IIACpmZbeHVUwBy7JK142TcEm+4Uc0jJef5
Tw7csQuwRX76GjGywcJeY5gJV88kP/dItKiikOkjg1UAnyXRh5w8wjDVHQrw44My
n0G0xccftazlIo03uFnVJqy1fOVxu2sTNhUkA54rLCIirKO0jF6U/Bjc39X0rklH
GTjMaXv5Ok4wsDV7E8aXWRRYfxBOF6jBV1qWxD9Bg+5/LvHiLT9pdfjJYOAOdEOH
KyqqZlNpkQdncmLa4hDuAX0vriq14NmQrPQZGq88VUpHGV470gudiFOsoybTgqPx
0mESeG1Mcjc3KxgsLCLIVExx0BEs395Cl2yjTc3kiXyTC+Zu0NKOrCb/sThj5xDu
pS6nm8NeVMBa8r3fViY9Ug1xuX7sC5IaXHx/DDVcP07Zpsnw6Nmvyse0G9Bcxqxl
kNbFG6SI6xDSn0XLZm4qjAN3uJyKMIFAOOy98psFsIzp1siuO2T8ug4zMpMvNikE
WfEE2hAg325QrWDNeb81FnWVoq+gDNxJpygEgG6FhfliBOOURnqK3P6mN1M2WNko
65awmPkev7bFQPALzsK9tkbpFEGVX9NMX3J5/Z7bWPnhZqvJceshNeP1x4QUEZce
nrrwPfOayvMIViOv8Co4OeHyxMqnA/xxsigZ/uMB+F20ZISn0/RubcED+V+4yT8s
bPg3e+cQ4CckSybiykLbe1LhT1dNpfF7UGeTJilTywKfAM6f47n2DQAALsE9i+z1
6g6FEP9IwaTCgyQpyloGaUjgz2ae7mufL9ajToOuTa4YsK7MgjKSvxfjvjtXc/Re
ygDFB0y8blz55PU3uCKnJtk/Bro3DXZ9FNvAbjHsQs51IFfWqeBKq00LCGplz5pI
CIn+4G9CotdnkZbIjZtH/pMQJTVWLlyBDJleWl8ufARPEA2ustF4fqVJ9J4nEkVQ
EaMJcPgSukH0sm37HiOLBaBK/EIV8nagnmG3Yl12DYs27h7cuHXKz8pu+eQlOJH9
9Xvt++MvHn5L+ucPJ4V8xVcufHjwL/T98lRyVvsKSb2fToe5A+JRGCvZMpW5l6pE
6tkryQsTVHwGLzPFMxLnEfrlVCwOJbTSY/TQnyZAxSyt+WqvAimSElprpGzcBBml
VfCn+d0u0VKq+zdkcx+iOYh39atl04i/nuv0QX1dXUrvKqr02P10ZhsM33EkIpFc
bJ/uv5cJO32fT1g2I8OpjP6IXHHjFq7xJj1zzKUUnBZ3Y/wiL5sTxaG7eppVv/bu
Xt1n8AGHWNIqjUaZgxth/k3FitjAh7Hqpcxf2cewLDBqnjWNTj5k3VotW4jySiis
pelvntOYsaA12Vthq6mAoYdFyEle3jU9Yn/6iUWmzvEZyenkgiqspvnmW2Zjg25Y
mYfC/uAXHuy3piLU4bn1TDWML407Q7mtrIBS7kwCVlCvvXkG1iBJpYCcm1QTO6Ii
fJcW8JMlZh6Fym4Ndm4xAy2KfMVdsIi90O0RdObSIYYJPuc84lsKywrXEor0/3vW
LC69mV0dczRcupH0/qVoWcFaSWHywQ1hBVUxmHbu3utKVhrYt7LcuDnOrkoC9FNv
hMEEAZshF8Ha4HHNCIQUxI+jOJT7tt0e1HqLoc+LG13zmfhBiyftW74Dtkn9bKmf
wgPm35pTcLHu4nWXn19Y9oL4WQqUol42JIs9oChXGD+TO4tlCDMphA4CFjT7NOpZ
Q3ybWg6R7VtXqzEXkrNz7/RVMjGsMFBY9uh0EKKq9d60Kk+paq6uWebixUZGTKho
IUjAtM4gbjlikad/nw5Oo/4j2xQ/ZIIn9d8je5ojR9afilndKFUpE6Z0zhAXCaGQ
wlcfmUkrCttaXYu5frZt+pTFRAseFn+a61SBZ61EFBTJ8zsnWf+PbqhEk4vqQsoN
sGCDrGsnsV+fUepMzLc3IggZYaiQO7iKfBOsAsqywePFSI0OHDRYNhv6tQLWUwZ5
tmO46ecLczhPQPZgqys9j45SjynXaT9ld1DJv4Gxicr9+ACqnKVCKsDnK9foelGq
+v1zzItjMRNliMgrRzcnhsBGjkvlHN+4cdOV+F0gwInxfxb9rAD3KjxT4Eh3Fehx
HE+EhwZR+KPWYNfqvFH1sWUfc3Eody6Y1shLFsUNdrCpDqqngoXKUCiAdax9pikn
t8GMNqqc4Wkg5si2tlyUumlOOlJYdeh8XS/kklNGp/1UVNK6qTYOrnSA1AuPbb2/
n9M8EKWr2EzkegZlzObGMmVUJ/Njj1eJr4xVz/TtGBKkf3Qpwa5E8xdNlPwdZ+H8
iQ6399XU5V+BWlILN+wj6TtCfEEwYqwN4l0JyuPHB3s9iSMqKNf1rxClRXrGakU6
fgoV8SGVKS5MHsR+maZgcFrqx3EgxMBV0AAuhWfSl1x1FSmgsRGvsB/3jywylTFx
hqritaO9yPaM45UPfa3aMR93FRFaaLf+C3gy+8V06VKPemu8ZcdNN9ZwnX/OR0By
XoewJk6sX5ZcCCXSkwoCeCoYSppCBBP2bfDz2OZlD1sl+45X+QU6ignWCcYMDcuA
LiXxGvSIjP6GaSaB57cShjHgZW623KvoeiPY5xGbKQBof4azOoKEKNPeDCAxarvA
6q/VUYefCSPUoWqtIGMCBi1bgXRvQaN+KthKvSW3esMt77NlectmYdmtwcdlBjLz
jrwZNUCxLayrj/M1JtaE80TvuiS+k1NIml2yrp+9pG/AVUu/iVzMyJ588S/AHt0I
fGb1e54cM9vTMHajtKu2DynArvNXMVv5KWSGEZzyJ3K3YMFV+ISajJHsSVtoIbCc
FFuDfxEn/Vsxf53cOy5ukwwBKoAjMbN+AQ4WnalGEe0CF46BFNUeDhl67XArnMpT
0Id1iqEalqFecG7CDYP5JzoRYwN76mGx+0SJfz1Fuok59OHRIX4koXUL4QU7zpni
yxPtV9q0WkfJvNVYJT4t22NkGv9Ua7yvDtOsI9ZzThk05Th+YOlutWlnEW9/eKbD
owOCsjrTrcEZymK0tQ0PMXi4RGmZD4f1/W0OMEgVL3iJQVUdHwK0ERPf3eQX2Wv4
WkXherBKdeaftCuCTQxows/ZDG72mKYPs5lhYcI790whJ+iVM9gOViSUv+Yd/cWB
tyjtvdDmdJhLLkvhpaKrlOXZc6nK7C3YcG7tUkNGKCphkWXRy2SRO9rXzTsHcC5Y
Aq4slOoPWeHqRQ8pNsN5Xedel/FTiyilZ8MCMm+LwMYNQKwuJX/5omXnY+/d4Cl2
vlrbqnm9pO8/H13IvRHfaADlXQZQF/nmfqCv3U3mxQ9LewrAQ3yiZvM66YYHLpRb
rL6tJZVtt/1rBfKaDmTaPzIgvGWKw7xc7n6LBqDj0Nj6sGDBF3vKUo3DHHcJfe5I
YMuUw60R2KZOdH+5mFjAzCtn+kLISpkVcV7Rjec70wI/Sqnjxyhz8xxScdRe6WmW
XW69Tqp4eXrrl6hnWBX3Tj66BEaaORt5SDiZcn+/wMI/+wwGkta37kWufwfCT1ev
Pkxz1tPrte1teFpSNAXh0m9gtNqCMisNitU1PIh7HCinWqlVfgV8n27+1Cl12oWX
VAWEJQyzThxhItOtrDntoR5fMw7UjUy9zNdocAKyhrUNB+rlCOwDD/tcOnfvRJWY
K3TGJGd6r4HP70SnZxNujS76I68gTXHGduEuE7ehHd1Mhzkd5PYYsy062T0ykHWn
BL7pb3EvuAmDIeHSvl6XQzg55HLhc85WfR2HlHYz7ypBC+evTEWjtQBMJnHiXvZ+
HEiMmCO3XKSs4BLO4XLdvDMMyesc28TmeIXvEfjDmXbpmsfqwenCbeFkFmgxcvO9
ALTRqAiTR7RxY4EtBLaWGExYMj0lsneAIQsLzE0UFiBJsx2KHiVjSLCmSfCQad1L
JxV8/gSEnJmMfykHAVqMyRiJHIThqiUdyiKdunKJUbPypYhuKv0IOMoNagtXfKg3
VbTpOVcwgHqn0Db2uuRRB5wPw0i9IxECx01g2RSX0H9LioPUi8SP7Ls3USSK7a3b
NrznSG5ufo16cgvx8UiU2tPb4jNztLGFIzBQIucRfovgC1/bTyj+fLeh9YUv3y2t
PsdWWunkFUV0+0rN2M2saCpjR7UG3jdH3Qkk71REDgTKKJQAHRXypRe8XRHU0sML
bKp4Ku+I/IKDKMOPgffOYOmE1UaUL04ygc9S7BUKKqKcJekPSVPoRy3HYxXxWEvj
MIub4SP7hXdUGY0iTMhTkqtvx9mNBBaQ1/oezNH3px+MXQhuRDb1Psmbn7pU6kEI
jmQr67WYqivsaUVTHiGacso9A4M+1Hl/EIEszLHKuR8i9ag9/4qXGIZ1IfupGBqH
slCggX3vY6JCbgG3aHgnzyJsuZeWvDEnjUIiCLeziImWakJ34wWIspgbJhfyJqlP
dxYpeG0OcP70VfbgKEASB2qNKvyF9B00btxRA7kat4d+K6YkVnMGLa+lHlCbziZD
VXvpPmEzFZ+RWNqWk0CfOam/JF75oafs0dAXWnk+gw3KTjxce8Wcx48FQoYJncP5
ppFdUSKF3re1+NTOcZMKQCNPEEr8YaORlkYwN/CkCQRfYADMaSveVAjbUpKlv2No
Had1wk9gXmk6q1+9eyXQCkMsdGMVrobtnyCFYVkQtco07fxjBeo298Seu2QKf/Qg
djUxXPWkhR49p17tMgboN8KK4f/V6pE9qfy5FGHo6NJfRTyL+xQFQ+Cme6GWacpz
xq/F/ADIlwhStqhlRsyMk+rpWd/Z0ZonWnQrIpPLVhcms2e6fC7ZFYoS3kiWFCjF
T/q1inCWUhr+m4ZYHcESJCpkjfTpBGzFKSm9boAp0C6fpD502HA8XGOIDeEHrqnu
DaVFG4RMt4xWsVHbHlD1ldvoRTzljWbS7gtnxuJ/Xkv2PQCTo3w4dZNDeGj+1Nma
ZvK/aa86sgcdICsKiCevE0tsLTa+4howayas56FFFjwXvdVamOOmwm9r3lpL+yhx
sk3zDhh7uDhAd1SwH43p3g57vvcrS6tPW1t8p8RD5ynK+hHkUe9LgCd4+V+LhGkA
hGomcLkC4J30Uj2y7HhykPu3pXjAjc9sx3CJmkPT+iqlx8/W7dyVreqcm5BLY/zI
RVmGZKirbnXVqVtHVj5ECBAqkgyfRKNWJhgwagKuXhhMlagtAURvh5ZnLrdi6+0k
MLkXl6ew756AdBs52gSSRJh5NOoSFgO9kz4rPf+Z2tsWl4lyjviYSc5zZNBwhwzK
2wVDS3XN8dHRjkziQKUSb9gBljSm8RHPURwdY2mrgjHLmRefm8CVcKE5ZTOotgHx
Qxmlo8lNJGU1NAfXgF80lMJ80J4DNSkedYPrsme8cz65bjv1cyvfV8Byo/9909DP
UL1751iypGtTD0wG7qPVFOE0ZkruTTTplCC1hg4nXGR2x/f00YX7zUoB6h4OwbzB
I4zJKmReG9sl9JKIwb52BL0o2vStMhF4XpoHtCSrde57QFK30OfWcJMBbk4zznoZ
kjf0hxDSgqnbuSdmHxQjQAtPLkV9yaRLcuob7pHkdx+WV0paaMWrVUCmijV60DcU
vSzYVRH5C/jSlstdg5tmrdDsJRSGyN9cddqCkt6svLkYyavblS2ivvDqyXel5XCo
hant7yWh++ypuEXWH6838IN/6bQiyuvL25rEgcTJGiH+0FK67/sseK1PI2lTJfhx
Jh7DhsTXb6rU7qqivJ3TMRuLHJIU82r7tk+4jE1axJkNDrJ8nhG2fMBstNblSGUm
DYBFgN8dBbAYveYHI0N+dwVDeCxJJiSUd4laTDzEETZ2GzxJPbEpvmLlPHRFlu4x
q1ThjQddB0eXflH2CTQFM4+yeXurxPwv7cpz++ZIl4IUcAm/ZpFLD5YeCuS1+1Xq
RycRRpSd2AErQBiGo60eABv/24SHpbbiaBBvTiRy+Zu15pl8mGjMyPWiJ7fZ06tI
FtlMYKhdH0P8Isaz2nec6VR7Waxn68xOMfXHpwgS7TtbNnzlsG2GZaFhVntJhLha
Pcc4F7eQkVKFJ2TYl5ct+sDXWhAaV3nm00WakHeEkUR1+9rWMPpRhj066n28eEQ6
tzNowfpnt/QckjsVit4brIBzTCKwZzSqdv8shlHi+2JJ7VQguclDASmb5D8+Hzd7
KZi9y/UaWO17Ukb/L07goLS5NmsmQlcpxs60fO8ZZpqbzRH3kRmrHySsE9RqIDv8
Mmda11rKSPZWx58MNDWce37lzsZIeOT+m/K3xRMezHpRoX9lwqPClUEVtxuIFG+i
Lcy7xNIzmZHoL8RI2JLcchhBXTlKtInbpI7Me61fOdhavsnIl/sOvQtiUN1XOkqW
ORYG6yRsvMuhQ0eohhzrdeY6q7FAO2mkEpFtaoRX6zL/l6dKLVclzykHWp9cFUh+
PnRKk2Xu33e8A/jfSVarPRP4JwGn5PMDMKYp2C+ADn0K9E+UFciXOH902CYtR7x1
lYocSCYIsmkXvI+AC+nj2IGfAgkBrpF3qstZh+Vjo2f3Z00NrsPnarxQf+TNFPcG
BCS3NPHeI4jD5LTxilUv84ee6sWeqaB6d4okyWhH/dmb8ANNGm/8b4AuFJAdB38t
m/B3bnTd0aZ/GtTYP/CXhoKwLjkc9gRD8MBIjiVEQmWxX4j2/v0XvFeyMVIiWLL1
cCc++JfcO/hU9nH9XEASURGAOwRbn4f1ySbAbDi32r1wzNUJDWqpIWm61PM01bAI
hiuD3m5BLWSeqm199D+CuD+e7pKsnC552R+b6mXBC9ehNWquEhKd/OPz2+wp4a6r
SvXhWbUT1oXtdY6iaB97Lj/4w7/7LbwVsPeAwh8kH5QJ9sa5eqEdHLk6PZXGhwqB
S7Wx+RTGm+MYVUQ/uPl9yq7QkiBPoINcjuDamY7b88n838uWMl8VSLhRzl55V56C
YWITAeWvEwsJR9eeNwCbinRjfiZVqPKpQyGI73MEbDAHLSiXeu3h4j1/WL89ngOl
X2iao+F8yImIQeMANtQyJ6H/2r1mjsXxbSlBYV63KLwrDOwbvguVrDrp+8+Xe3H6
hrTLmJZYp0NhrSCnfeLbVwy1H2PgWgI7d801l8kgyNuYRI86C5fWJUBs+o2/n/2j
LjlTMuPfOovMHAmoqPHh5WSYKoQQReuOqt+nA8td0XM+Uy0SZNChb8jG0BPXval1
A92kteyEzCVgaNq+I2xkOudoLM/HOA3DhWTXb68sSl60zIlvSmP7LLPbyEmV0e+2
tnYXccKQ0xKlft0dQtCdhbCSfT6ASLJVJYUj4DoAhNOvRKQhVvUXgM9yspoebujv
NpjXkM8MQtDVl5jWsCZzrm+tLn3Jb/f88gdy+y+Mwchdw8lUEoKGKlqS+EySNE4z
SVD3WJwF11wA4fN5ncU59GjiuSLrxmuWrzrT8XheYkMfDMyPQUws7vy2Zvfom1CH
3jwnQS4yl++o2uf4+lDwLEWAY4ViPcsSm0Nl3HI4bBJqlSH+M3rOjLMoInHGG+IJ
fz5SAfWAGpHk/VhDKGj8/xtg/4hK2RYchCxKvPywfnvJkfIFDGC/uEK4Cq1lhzIl
kN53qKIXp/dlZbdppqj026RNvwJ29FMYuoGuXpSc9xI0gvdbGkWqkBM7v+ENrDXL
k3LOTT5JwuKAXHvBq8MWWQ+XWXl3/0vpMz2zjEL4ZBi7PjED5jIc9pe/fhTiZkiP
guFWVPLf9EoxMg+TLaLA9FbqQz37T1itp/56gMKGlpV5mdcGABgguGsz6m7rr5BW
0KYPQEkRugwMG1TTLubehGl3GY3uxbbMB8yOXrTNVwQ41tRjhbqqIpnyF2FIfQre
l+KW8vL3guH8LNUDz1Vh86akwrM9nIRs6lKrbio1M/C6VVSxidTmT3udQlvKLWB5
XFOEc9TFTr0zKQAOcd/PMELz8a1/B6hYPD9WBCQ5gmdaEKKhZ5yHA1WyLBbVFvZs
jbfsHNk1hmTuXTRIOpEgOQyvfX8CNw8Fc/U3c9WXrUQJ0lL9Y1OB0J9M5xxGkAZg
G97zaZroelejKKJCK8xevR0r5V2PbG1tXfvQTr0f+Ei4FgadzeDbWVo6ih6Vz8zG
XM75mPhMe7QScHxVAM6dV8j9JV01rUITRRvB3KIeh1gSjLirxFrZsCSOL6wa39Rd
vAthI3oKQYOm1nOz0tDmreZGjjD7tpwXe2Rh+CGO9nH5cTf4GWXRqs9TdM2atlyz
+1wHUmiDU2+9zhrEnCP9EdS8HKCBIRIWIeSV993GfCAU0WcnGMVr1IYByEMRrWXe
mUn8AlmyHwsnGm6oCt7h2nZ7p/E5TzWO4CCkIObz2vey2wTlP58NLnv0nJI2OKeA
/lmLOkXm4qCliBxwskJmPX+/X7JKkxl4NQbi/T3h8eSQQSHsj2aQScWhYT7tJ/6L
qgAPvesT+m/6AXnigZb8p2iTN2GVeYecYTom049PE359adGJly99qDfvjcYj8tHj
crQmmN7uLslNns+C4Qi5+Nt2XSif1SccToGrdubbHuAOsxthBpcW1EAaUDvKMX79
TaC+nMIWZqahx9vyk5vIXXRP2JKGk+Znp7KapD4iUXbsh8vApAXQME+S8APwtYIt
QLXWVpMR3GYHIyUP+PJlGeahZw9imDJRlKgvpc9H2wS3gF0KUULR4rQnY+Thbas9
1OtnNNnZUDOI/fQIK3k6PFgA5j8kllxp0flAy4foSqftMPRcQ5K65nVOtCkYDRDj
ELW7M51nXScSDo0RxWC8sKzvC7edFmA5uNG/faZeR7Vuv10A599JpoQtJA3JG2EM
9DE4Bnpy2bvY3H1WDJtPBL+FN9NCVJWdHcvOFc3/Hmk6DHpwaYatviga0fIh4mvg
ZTI2N02POGcKlIP5Qq8CfrlWxn7GAiy6pafJULgnerXeKlgDOOsD5NLh9LPbgf5Y
zDCfaWhJHv+4BZjknQsjuA/XuHvlpn/hD80SeoErA6nC++2OlMAL0xBsGsrDx1V7
LH44qJooDQ+Vp35rXD5EjK2KK5NPMDajWtg+CQL4hnLIquehM6fReqp3TO+UUdyJ
ZG/XyDG0k54KTTIMnyuQkY6Drd17LENcy0l8Jjd04rgEyE2u6k3V4f0YuS/c7nIW
TKzgYtSgDDqd7EnS4ytWwHoVu17TmyikFYWxuSBkxptL4a3gdVlDiKt7r/pefpwE
TyBF27dUhzi15Jphzg9igDE7myK64pAkApfv8fghnGfOVvLpQUivqgruOITu/Urj
XAPGA6jj6Z5VaPI9zRNMqojnCoSu9raLNIcvswHm3QzwmsFOgYxlE+tP3gjwP+9i
+C13wpyBMTibc1T7uNXvRqflPvQwMkqo5R9ZNRzMN9Hx8xOZTMi3njv1+2FYoY0X
QdP9A8Afd+Nx/JX0xgARSrWolP/K+hDu1ArSFUSejM9RH0U0YUKa4B4upEpkZTAU
4XPta2qop1WhCTdmCPhpo3CPyGq7/hiK8W2VBOeX5+8HYgX60DdpK5tRoUMX0pCr
POD3Si9TEOQ+/N4GCCa8swtGDi8Wtogy1HEehK48LlseqCxQNKD9gDHLY5NUaLmr
Xr/gu1n5XanmOC9XPnR3oihP7PuQj7CPE5zZ3mMBT790iHQyBdrmTBd0DO5TzNrR
mmMytR/zXYZZ/KDQUOoHegvEjJyM3beu76GRESAsAV4+LAAAOb5SV99oGJMRJiGL
m0+m4POjtBN6ZuUhoZW8I+cdcndeZCpH6+g/DLgjsD0Ljrxy4DqEZsR/MtIa1EoQ
eWGhOhc0qMwIWziOKDvWnvMccNfuLNFNv2r9yxTAoaH0med++Ywyxeee1Ax/rMAL
yTlHPAJb5/yIIJncqwlDQJsnHwcKAEt3Ig0DI9xiS284FyOCLrW2RcYrWLblXyzE
5WHyUgb16MxrMgoQBRtsuH3RpzTo90H/5GNQph1IrbVmRwHofF6MSnhbDBXBaamC
B4/09UQ6VqnVF986iL6cDMfpHWggvIR8omP1hgfwZmlF135PxiM2NjyXEB7l54zH
u9hlqRLFMiumx6acPB1rbZNHM/7GxUnwno+I1FqWOzOte5m5+RBJzI7jM+7u0zNG
ZR/JnbVdZ2dSbL41BcT1k/TGeOWJkoZyG1z8nAjfa4xmStRiymnRQRD2m0uoK5IB
xIF2NrC1+tWBYdY6nzZAS9BOLwf0uF3o6hwwajc+412hr6r4jgNGAHI6o7lJkGAF
vhEGr/5kBmHR8l3dgq1RBtiQuztS08tJplr8XR38gOtwDrtW3oRaLHFdyvPIVGYI
vO0ppD24u8Ysjyimj498Gdtmp9nUth/mQQSRELzbSRCR8C/cGuqVGzsBqE7UB2vE
aGWDaNzb63tTNmkveXUj0zulzVXSd6ggfwUpno7mtdcFsbYEz/f/4dwzf9OhzW67
7P2Eaalm52evzU8C+//Gj3cm8d4dmAaHnlLwe9HNf14RzYcu1nTCIKx8yhTuuZG0
FaB9iey2+ym3Tkogu1safxC38hN120li1SufPS1znmFzoYQ3fl6RrX7FJKXHIHR4
zUb5bMHCMum1FQbmsLRcmlSE0hoq94vNe6IWpPzNd+RaBOUEAKh3eTq26Pa6reV5
IixrJJn+yuhvf4LzNwhJ4taOsrcV+3IOpH4UhZ/p1o8Tas4imemKk/YekRMe+iI9
7HJFPYylkAn7lbG+SZq6eGpeA3dFuSCccR4dJWRT1mAYkG4pdFr7Hs8LdROiK4/g
2WDare2GXizO7XAsqJczmxcUgkIuyVboEMCQRpr+LOf0ooj+40xKKj0mK+WCi23P
l1AFpXrxGZd+SQv0u6vabJgCxqE8FU4O7jrpezBY3Xn4hb8GybVLZccH1qJwMym2
ocHumug5GNIr5CnSJ8cH7ZkmkREnF1fx+bhO4Cb19XCcxfNtZoH6GC7BFdhgC0Zh
m0HgGi3PNZjSxiQNq9+nYtpMxzFKyjF9zRQIQdAa+101QRgMtBe8tscXpL4LQSqk
/X7Y00AsEs/UzHpx3mz1FBind9ZY7vS106VSsP+eo2u1cG5gu01ObzOo7JPj+DGx
b+QDaCTrg+oqLBocxJLY7z8tAwp+f9ixyEHmZuAQ4+uAFRlB6DYAXHoxSzTuPQCT
apViEoxZjmfP7qMX2W0a1yx/oKToYFxLW2zqZRb+oFhGriqnbwVn8B5Idq52T48Z
2suMLG0YYk8KMtT7klum4XfQtgMhKas57+lpq4+JkGkKUE2XVxYmvvfGCBBGfOQA
StSp5xDWoQcjqqAOxTO6uISbFg+hPt2hxCOOOhy0fcLzQMgIFtgP3nK8mxyFe/uP
tozVonzIkwSNLG19e0fRXmGDfoXS0y+a9THMfoiomuXXh3RKxI5Dah/GPqbaGC24
N5uXNyViXWjc8vJ0eu+WyaPwz1tcqw9Wt2H2XytWXyj3ABIpbQ5pB9HBjjya0xRJ
ZMfmz3zpKwS7KWlAqcspzS/p6puVGbp0efVXHJSBK1CJUWNjacG7f52l5x/CHY0i
JpScQQOpwfBnCEktlJtTa1IKoLLTtvlRsbDaVuwvbBp6cF+jtBOldt/0e7MjQE/J
QXnoXL89KdTtlMfIFVPqwi7LXSEtPJIV1eqoKvnuPYw5FitCATyFByma6V43PSKu
aPscr89DXl/QeoIM3jwMB41h0SU1Uh21JJ6p7WG7r3wdp+5PAppXmjSM7hT0mbm1
j7nhnJyVv/4wV5To+1yOwah41f6gcdI+F4kF8CMPouIEtJitQNpfjA457vV357vO
H+hi/L1NuDlsCTzXZiJobetqDElvu27uRhSCwaOuiWG2FrR0IScebNSC/BaSoj7y
1sjbGmefjR2X8utxd/4gfQ2I4xLO2FzrSxGKeRrenCqNygDF0lxvjhc11JZSOtzf
EW1IUoPlZ2lMsrGnAkTXuByMttC9s9L/k4j1Il96oZ64mcFGjiUtBdxoKcBMAypD
pYkYeq6rqp6gk1xwG5Ruk2xlFS8QHeXb8kkZTfnET1x2NTER+YLYyCRJ8gGIez35
CJpwij0EdUffi+CcMnefaEJV5ad2YKj4NQl9zQM02F6Gv5edpDt0kz/YGCJSgGMw
6SWq2Qx3EmIqR0eqc+5a5rOuydroiXE1PgVHnNxwSMmfB+wvfXJ5mHb3fPeJxPYw
E264U/v7lNMe4Edlfuyh5es2clCfwVLhvzmdcWAK+BssKDI0ZcdDu7MQ1Yufxcrs
yJ5x7X13UEHBrGYlNvscj0rySFFn7SxswHCLc8bZLOnwOycGtt/HlwpjK3D/8vrM
SclfSm8lTP+8jKDubl6u2UtYOW58z7jfYOm5xePnFuVApUs4ginhBilxrLTZ/6fn
mKhRr3yJ3LyaZSft/pfe7HYlsqahwQyeelnnaXsdV5IPlSVX0r/DPqoWR6jTqqZF
17WiJKRfLRk0sKrbm7uZZk2QvnsIAoFLBFAMVGs2dnzvvJsVR1Ti4LOz/Xm8v4wk
EFClHYwnUbiBe6AWaXAr3mwjSkDtqf2f5tb1iabPLURZLYNVMOShG3jNgida3OxF
zzIveEmXMXwM19ExUPoiLyLrjcIjLv7b4VoCLcGJZPArxaZr3memF4+xoZu99aka
3CMKLVc8Ve5VuZgs3D5MeC0f35xOUL9IOi7pNu9ttN4iL1boJ4nEdcLS48aZRZRX
r8moe06wioQvO20KL/TZ37p6xLBW65ccYGnbVwUfnS6xfMYbeeUT0ytWY1g9kb1b
KigbUuoU32TLfwpyC2OmDCnGMz0DhWskt4FIyZaudWywXJPzH8rdIATCyCxYOdW1
cLT3X/SkLa0Z/MZCb7iSxZ2v5Ha04j0r1VgwkzeAcVyVGXEUFwvzV+kTF4AWiGGh
N90KpAe+TnIvQHpCuFv7vvlkOufxIYOiftLbNDcWMicSuiXSAz4NHlqr9LwlniHT
RhQ45KqD5Zjc8Ujzvl5HUxlvUoDt4fa14E04w9mpXhQu/NxwFYcVpsTO7QVgXWu6
cy/Ep0ZI7Ynzb0gf/vt8iWVTXsQKGDhUw7RBu0bM2hmUeh/7N6OjgofKdsyi9O4F
c8lzk9N1dfNjxb6wKDxo6mRxz14YwXCrLg6To3IgcuGcA0z4qamkrLmf77eKLi0H
Ba/PmCrjSzpNPdqeAUybxV8WDUAlt091vaoXzZBCIBexS34ngE3oPGr3tCcDjC7W
UO8TrezdbHY+57ZOa4T+hJRTTPYxndX+0mmnCiCCUxEJJq/8swUuw2IqhpbJmQug
qC+W3FuzcR7M9VqbVcVHyQIZk2VS+9/IDwWs8MAwty5zh9jgwtvlew6LbJVo2nzx
W299Y2UBrsTWaHSk2/REVNk956bp41i9fm78daSgkG0AmHBLJ8mOrCGRBe/IE+pk
zGwNvcc839QBhEIjghGXJn+G/NonrcYNSNOmRUhbYC38FsJ60kaR0POG3JEnlE8h
UBxhB5kHuxJ9zGVJESeuxQ7DIkC5JoljuQK54DMMkeXdLSgKbWL3jgpISt3KyaPZ
dMjY50SNFCHKpd8cFpJx5KHhyntfgmxMwpOtDEkb5KPbk6WbLBxVNJoE+YHCqba+
i9HquGD8jOoyNkJR8m0HjSeIf3nUaooiIyhdCNZG345b49U9grWvdQFivQglX7ED
SAQJflnDU6il11zfZK8SejxYb1Zhfv1GnbS91iYaPt56ESJ9pRDpGEXLtnCTPI3z
QatRp2WDu+megRitF59qrDnBQ+dDe5KKWWDo2BDginZtHdljxxTsl3TI/qFA0xFR
HSU7vdBaYsQm8iwI5N/IgctqwvVVOGWhcBYI307scq/xhrPqjam/nK7O179pAYQy
idBu29n+K7N9SbLZmzeCrZEGOJDamA9QZkkmVbdMnf59uyarGY46HPEDH1+MTGMR
uWyWyF1oflfSmql09HP8/L4B6t2PMmSrlSoTeuf1xrK7C74DzOuKcYvysfo8Mywd
Z2eq471fQ9Kv0o98QxoqUvpZSQ8JdmXBWgal1k39vcUBxOnsL5/EqZ2XEqI2Lqkf
Nmy2EuaT3ojJWt3e3tEe0/67ntfTBnccPHgmaZKCAWI9I7s+ZxVuhkRqJB95tlgB
zRed/zBbnSJoseILzCjukO5xytaYkv1hXonMYq+Hosk+yd36o0JCAxSyXJQDOXoZ
qF7q26itO1wYCPnsZeOdtAG3sKtivPbC1pQAxdbnVx8M6W5WfEFdCyrGGgvaEnBR
G9HzBoTnHG5vWhaE3Vxyvq+IwclAE/TDXxG41GYwLoqqD7yZz9b9cHR5UDi9awEh
OqJ+ZxBG5hIRWnUMh+57Fw3kKJ4NksmLDQ1OgFFZpT234EXM+U4P79LaB4qULIs/
qRBGUCjTNdQ9acYZd1N7dwcyrpLA9Hd5HeOf6C9ax+DaHLgkBgywIsFuVl70m+vV
YLYkbHR8b4bQerGvubw9dwrp1h3b/JIfJtDBtLd66W6n+RUCelZ/71+68o5Jc6uZ
Hb437RemyissZ+HzBAjSwUgGPqSfGDAm2IDy+SuzJEDtZ/tgXaIfCpWGpyNFM2xG
/jCSLsXvy8ZZ6ReQcNmo5KzXyNuryXe+W3CWOkl8cPfoGiC3St5baqWXx+qjXK/K
a6C8pOtMycDwknC6YVtwo2h5QHllbE32qWiQzjuLMNeMfDaA3YdYx42EntKI3oEN
rSarvnrf+mMY5OAcVGqNk0OX45KsvaRBZqtCRsneukZT76URgNAp5fkJmxEvsNtA
sJuQ9I+L26PVFRuiaFkRUe2t01fHWJ7fKGlncg0RaXER0d5tssLlq0AJdFeyAubs
+4tvP097l7htCx1/ZuMqhP2IT6gbbQyQOrX5yMr8drxn7bmUU3ObVxlMTUBqJsp1
BHXkAQEBmrtDSCd9T9OznpJc4Heh9rfajWvIEMQ0Q+DI5Yi3EOUWzSQV/HuL3J7Q
y7KevzQql0GA81ZAhxdy10ltsoC+GY7X7K2ohZ2YAt9SPyph8ZAHXusWhlwk44w5
nwGD+OsKCrh4pofi5l0UHQznCyny/qBydDgJtmaJ0NB2QbPecbsHw5XFYzNnyaGa
O+Yxo6MNkzFZMUhNcuvdEBuxs2TX5YZKrUvmOFcp2xJjVFxkZJIfXsc4yCstUJRF
7HugBb54lD6tr1c9vvv+kzpGzBt6oWgH+ufc+Xw4Ro5Su0Hxh9ZJVcoO7Wh+dmXT
ITb3JriCXhwyrsft+oimPDRjYE2d1cldl0hyobYgvR4vfXSxV5wypi8kRmUjQjl6
SL6tXsuVoHiUpR81U3tOzdlf0osMWeBdh/3Zz0wVj5adzp1bf9lORLKIJ+hrr0Ey
ryWkpqXgpyHndKKQd1EnWKeZEgLJcRb8Olcyc6twr90RgWQePALgG5a4hZq3FnA6
pXI2TpQaVLxBRgpAFQlf7l/mUjV/CcsOIC7GTWqNohRj4kgukKLWdwdWQQnP383/
IYWg0vR+qosFEMSx0d7BwBXMBcI0zZhhLL8tfviieOMeepnR1p9XjKelvgFWVGF2
gOhzrLiCqs/KjU+wzyGGgNSzwlh2hfAUpKjfiAPUCp5/pSpi9Xrotjzyojb1PxnX
xE9tHRkWidn2pylPB3S0qTxiC1JOWX9qvdVMjlWFnJRvA0gjyNW6LNt/fGYTu9fP
GAZ8IQQXueLFD3UGPpGql9EzgoCNnTKFM+G6wUsweTIbzIKoU/v/uVYqklwfDRi1
mEr8t7OzV2nLWlQ8PVNuWurmI184wCu3BNi8bK0o0UD1lRGf/A2mk6p5EWstGDC0
Oyljwydp7M2RnWIQeyCe5Oj84D4WS2mUez/xqBtEna/Bzlro8KBFoJewyvNB184J
+mWWlfrWwU38aa7ySkdwDYT6VZ1oOKwGqHG6b2fdkwPaR16z9ap4p89gBsYFByRH
Lh0V49WGtJyn3h/wZMtUtj1sZiq7bagSc2xsgsAP6eLoFx1vLX1fu8nE/mrps7o7
vVSEOyzB2xaZIReQiE85OJgMLdVU8SR/xzFHUTu5KjReIm7hfoos1LNPSrl3zibg
g7aamZ+oLMmfRx/fQPZcNrqY7Dz6pl5muei50TcwhCpYkv7Aw1U02WGsofHMAIRd
2J2v4+SMudH2YkAH2xvZfI2gBTPO6us++2b/iKChE998PD++sD2OJhyHWkOt5S5Y
BKHd30HrjSp/sq2rQcPnP6JNbd1moSzeuVJ8nGDsGH8B0Qmr8n9PfDCO2Wbx35EB
YzifNpqMwb2C2PHKWidXmnF2tEjn+nDSpvUSI2SRvOmTuPoiA3bienw/C2/OhwPP
WZnxgBpuaNxZFx6HhFI3GECD5mz7Ic0d8JxSeJqWeeqxspgS+jBR3MPgP7vaIiGw
O+0bTDv9ci9YJNHSVGpyi81ln8PjYycKfjp32EiCpiqt/kUcpLQgqK84PwwZ5E4i
hwRsgBEV74ozjruK2aacWPbMPJPVTrydhZAlBVS9e1byMJEoKJOTTEjBIcQ1j4oN
W7aN+MEbEc6I75uqmNeHhv2hZuSwhsxzzYXMi8AEzTV07pFYb4NB94Hwr1Agz16n
eBv6dRt2AgTwEYL5Rdje2zOl3khFOo5UmY1YzqnwGMqKUZRYBv72F6KDWkvtsv81
EdYsMAM5AdcuFUmXfCjw2SIuX1JpDyKfIHhje3jp/xPq6YZtDL5Rtgl1j13Q4Oam
zfRxhe7Gk3Fn/ZU+OB0Q3BQYtdWCS7YM06M75drLTjR7vzkJFjHZeQXlvVmh5skK
+e+wy285SRNFu+HMjmBFDNTee3Dm8uh9bsOxN8tjrA7nFAwW4TEW5P7zegUjN5yq
aA4rlVTjN9MXY1jO9Z/+niyG4IPWs8fPckELM/bHt8W9/bONICQ3MSejefK9MLmq
UbGCxEqn8Soih6JDZUCuEqP+9NEy6+ZPBv8Fs9j9+A3Ewdo62yo88RXFzgGHNCrF
wckfNsWfjwoBflrnCL4SmhO2QbffPVQ8PWSidjMKUgmXLDSe0/2ke7UC5o7V32iN
H26pRRVYAWYVfm85pknc05q0cMGIzno/vKAY+x4Llew8tP4bELt7gALy4PPoT64P
yF58Zkix1DoK9Cq0NylfN4ag5xas58iiWRtVec/wLuWJ+dBSVM94xNI4jVdgZHu2
F2q14q9Hl4jxtWDBkbf+fV/euMErV49d/d8JEAWJbwTQaMmf7R++s/giLZxZZWOx
Z+75nbKQG8mTtdrFjGwlsyXy/gv4bmb+0A5ZJjNh5M8/uDuxgh5K6vUfygUXShB7
2O1QjB2pb51kTwRep1Ziqku7YDYao1DbYfdf9Gh2hgEZVfTJA0uHmIKds1n6jnTu
HrUxsn64TAcgOtn9uahP1OqbaR/ddJUgs3j04nxLq50FKQnjFm21Vrbdfkp9G0Vm
jq4cBQkHh6RpwKQuAv2rboxW6FIiLAgcTFa0HMfK/0eKB6mlnpTTY1IE0zX9nQsF
EReW5lONXM3FjS2NPK22BAsSDTngTAyxmSucS+JXALWrieUiwFH/DKP49AgZqdVe
X/dtkNcPityCnNDboVw/AI7Y0Db5YAAXP5pdKEh7v1ILQWm5LxRt53DdR81s+FFJ
GFNTVraUyNvZ79aittvXAutu2eMZx9c7sYr5a117SgmNscsOHVLZQQ2EqVzeck04
zUcidHgFQ2PYnGHiKj6rZKBji5ftpIdCD8nwnpkIg2FgDgfPUVbIBqYdLdWlpke1
1CQdpTMNZKD5hlFxCfE4QdWfTZX0SjqlqPB3ucrFvYtcbCV2Qvl9WlrTvRSARX8H
q7GYu7szrzn0jRvwC3R/QijDZM98TpPQd0vWpt8kAFsZ8f2NqlKiNPg2H1iKGguA
Rp1QI+VEn3XNz6Vhr9Y/c6F5ZR1lO7ZOmv6Cfq4AbarhagQw3N5T1DX7CYmErnqm
wzqIsgr/h47GURIjbRq/U5HnuvORVi5+Es95H6TkhcVUm1WosOdkX6ugVYFXjMW0
4Jt7XsWZlwFZ6hD1s35EF/4/a2mvc3FU2c3oTnazIoIBw0O+6uRMW9vxBhpccgHc
EQTu2fmt8UC7XWsTte4J6ncRuOV8sbd/zP/fL3AVwRy9S9EMXeO1YJo/XSCQUFtW
aA1Rna5u/OJmfalilLRRYsb7yYb122Klr0p8SQZ7C5FGy/S/umkfzGfvC6hPfxPr
IUuOSQD8+0t5S6+oFGfRdwOsi0PgkX13mt11eGfuyhGozSCGwXswW6kbMt5BjQM0
427bE6EYX6oArjGbaJfSY/B/dzR3ud4B/Mlj/q5U1j8y4oUftmP8pjgzEl7cu2SN
EQe66W36LzwIyMjI3EWm9q8nePn5/Fy0+Dx/BIgFq/4jIiAQ/7mcp2zQ2u4O6oT9
wCUEJ9X8CnQRCZsKXuizgNsKnNX0uv4rS6KaQLKs+04pvJccEkDiMVvpeD0nK+TG
o2abqlXTIIrZuuacq9SqfvLg0PQifNX7+F89LfrEj0jZFjrdREZ7OYtC7gbFNnvw
Or6XUlwU02SCNrSUd3I/JpJB/O3T+F1XA0kxTBT/3WNc03FVx6PzAYJU+sMW5gZ4
usOMk5ShI9T+515lY9PE9brTzofeE7Jm1/BLCD+fimIOj63of+LKRWVsHKM2J7ex
bmrcaD1qke+ig7HX+ApREOdX5eLlDnseoeAEBUhY3UKr/18tAwl6YF/8w/YZWcKI
fpBHCeNp4ry0eDJumCE2GE0MFKjXTnckG3jE0/tVfJy3Vy7xYogx7zWd1BaeMHlH
32ygofh3mKtuY1mCD6FjAazZjGlpFjU46hcbyNEebr3K8yFJQ/tN/XEm7tXDa6TF
ZRWqQuFBIBGXoT605+sFMsaoxvJcrNMnVl5YOy2wb3sKJl/2LMvLcCsFk1ZPGd0M
TI0LKZRl/L8lSI/0x/3Zil24J+aSfK0PC0XSxJofDkwl4JJGQimPTMgGPV1XsrNi
ME5nI0yZ1TqWrwQTLyviN4hjhuMHVKsokPjkF2DbPQ/LJ9pIuDHvybgt/lCglxjD
r/fGDoFvNtQj7UGF6P4i+RPB1GusX6SxHh28R7Lo5c/jY6jNignCqBaZ9AMN86fj
LZUopy84c5XM7lFxyCfFuAQd0Q9G35kZWN+SHzkdgNOrUMTuYe/xS/BK8mAgu2E9
vcmKB2IEfTPTQ3um3eADqf01F2oRhHH3CjcZuvtytsNGLHSDugSsoXHs6yA6c8W9
mVyNR3plySPjhIF3ey1K7A+DdHFXxyVzuiNQLGhhKhLqbKWzOAaGxAV1JdQS74N0
ogJ3QmasgKsb6CYoYWHxNVYjF9YXv4jOGzzQHGlst95g7MQbontpNWaIzdmStDIl
buTxppCTwx7K8Net/Fl45PbcdLTLo3vnGZiGfu0w6LxxNIosjR/iXx3L9pvG0PPH
1l5/wnbHd/BvQPXrw7WtAiTjSd1JAIPdvzLSK8b8sgV4wudmg7+5ddy2eIo20xTV
3Dm2EhzX5qP5wkSrc33m42SJe+tBguK/+WeTzZyCVbE2Wkbva7pWJeFCffbMansl
lI42ZS1WUDRtMI9qNrd73tVUNaMOmKJYZDpB9i306Qp3DU7VgmHfvJySRzbMb8nh
S/0aXq//H8jmy87hMREuaQpnJL4nhTkuYYJg0Cs0SJskjbQ6KQvBc3BMpvgOTmcY
WQ1DhB9/lYnU69WpLXISQ5lyXQfQqHkMcuAuDa74MV25ADcS6crt3eclut8fMaSy
kzKP+4U3Z/ebGeIBSc3hkBkBbNLwGkSLRNQiGFwxG6h4bsKccCnJVv0zpq9EEMx8
KZLHtWi9j/kCjUZszWB3ogzeLNFW8tFbKnDLGELwfA7BiZ5kVGO6ZH8PL+WsQb72
lbE5/w2GkP313e7yMr/tqAwmQnRmaMvPTl7ebYm6w2rraqItwDlZ22jIN+RZOEqT
1cgywF74h+uetcmebuD3ZFxlcHXwZDdFhzOd1jtQQp0UZBXlJm3H2N6fK53rd/eB
ZDX+w6hccBqLH9QhAaLKMgmkIxGsXp+ZsCDLcqAt41DGV/CBcnrtGVKXsN14zfAw
qYohVI8ZNY2q+O6ckCAOsqof9P3eWciOR+NQDP3B6xvyGu8UNc6O4LsxJHU/oSRR
/qa/UQNNiBZV8N6cjnkAuh38TWOhQo1ZY9q3z13vY0cUOevTIyVxrPe3IZw7xwUM
5T2ONS0FPWCQRYWEF5RxipPdXOdigjDrTJ7bZhTstlR4nswL2HYoP3U+G/YLOgFS
O+ptUGmXbLdEm800yCx/m+okJGSEzAi6m5CF9b6S+2dixi5g67v/TwssWVpLU463
WiNXpsJrttZ5XQ1j99kl2XqV5sH5bOORScrK0s+oQK35abBKstHjbC/G78m/96nn
EO9Bjs14sB5Y2zF4aw6GrrDnj1NTyUGb6IGc5i02AKPXxe7H2DaV1po+evGNyLv1
vk/u3Y4IBZXs9iPl+EfsShlMbzth1ni1HjjHMDdxqgSgUAQCwgKJ9mXVKZdKLXwl
A7F4tL2h6MheEvy1VCKTXHxyRF+D2R4nAAEzNdkfkMe32ZBxsh/xowqlk6VQwP35
21uJiYkGocajBJ2AKzQzLjIwT3zng2rPmG2fKPJLL+QY7cSn2ro14DPbcZ/W8wog
S40PuT6APVj8UL/FFihT+1wI62p7R+XSVv5sgnbChTgUSSgMlazl0KrwjwFQn8Sx
MuC2zXoQ/svgjMoTciOQBqIYattf/b9FRZeiMj/MFCl1PBaLfB2X2Q2+gHg+VWJb
lMyzNrDXPGEh9f5XDGSdoqySIGewhD3XsqLo0jzIUIuk+Z3CePAZP7n/pokQu2pm
mDobkM8CzqrwO12G3/ALomcQPJEflJEuwvYyxoizirXt4ZYUm5HvRORdYFpkS1LY
XDLMKhdG8o/WaXWpJrAFBAdqHu7rdKCBHK9/OCfDs/Y3aEyMIQnFYjwEmqP0+Emv
pLhjvDSUJt5yFEbn2AYSOhIdI9kwWsJKwaZjMvN/r3C5sFXKvGYHU6XOBjNXsKhq
xeMXmSLwQdcOtQO8E1QFMz/E5bu/kpWTY/3kMO/MeSUvvsyC/WWBjYqThIj7b3jj
23bjPIyTTZbHNUcAVrBKGicLqlXQZzCOTTAAYBFaqdK5G2mjukQJEDX0p925nM6M
VDExURi3twpT8AXh008U2AcA3KXm8qo8c8QN2ecgwCTAXUOFd6HU+jzy1xfQFz91
v2Sx+M4a/HTXNShPRGVaJ4UfQ427vWd8p67yCvBHzsuliv7eY3M82RKfRdBYCd7b
19D1I91fCeVCVIaSLaZhbXQIC07kz5chJ0VfhXsYoAXrz5hxvkPDzmADQ4iJd9xi
vOvYMZvD0LI1y/WO2EuNqHNMhMStV0glx1iWyShY3F1HfVWV7zQxGeiuSpI2rqfR
dfgJzAKcbupbUdhgPldmkn4W+/GXdDziGSk6sj1OJybVHtI3BlhNZMANAOqiIfqJ
BKQpWBUrF9zFHpUQeJWXodB/7BCDcV07td0PSMJSo5FVvt4pQRd3kUGysJu/QlkG
C7bNxBft93Vw8emgQIkhVYhjDydEaaqFLPfgSQQuhtS5za0YIjwcWScoyAYDqnzK
gjbu7VHEiGcJBQucz2egH7WHWYbv9rxY38fT1a415+PuO2H1U+pB+USFLQSf84Z0
XZjQKZqj0NwO+9fPhVXlGbzrzqmavGeK5a+cfT9wPz6GWL93R4EdXz/KSmiYvmPa
/GRPULdo3JDdfXzdfAmbGZASaClXBk402eLH34bSYE4yETQl/4LL9myH2u/LVxFb
SFae1X3kVsZ3T2NnBz/6eZaE913DXQRr1R7/5n40/xqOEtzd/V7HH/BuwJ2fnoPT
wzkXb4YT03tYyylsfeZmuKr35Pe5l74r8vYaxmN5DFE5hytlF6CSxmYjVF9dPP0S
gV9YCLh8zKz1rRxqt6yjNfww6Sw5ZOt8HN0N6uA/ETgoXQYpYwOq/VbWrFAPuW8S
pOtNepPjD7Zd9p38E39U4Wk5dCbqhlVN9k85mmOxMgR1p/Q2jTcf7eeVDC24hkmk
Yuzl/8Y94nYhlwXyFDIOrz49YextFrY29Iji30mSgTlNhPrn2joXMa4QhQB6etXt
aImZLjxXgCu9Sz5pYDvn2HQAi/Z3O1GQlxskpbXOPQcc6L+rzVXdXWTYVYmtzuhe
slSZ8AsHojnUWIovtlomUlspKJGNfgUyKrO6TWStJCkVMr+H+GxtkuapAlmxNCqk
tze9HccLCM92ecOgHcq4Cbyw0FVe2FrvdGI2MuZ8V1tup8jiRNus5Ec07ljhMZ2T
TUitD0hTEFqcfNTMx2MTME4GeNJYqt/MdRY4Tsbl0E4oem90neJSHnoeqAGfx2QX
msHgtuBBkVb88YOWFJ9TkPHXQwxnN6EmzBUwowCF/3pF6+8cgqn6dRG0+OT9hs9y
zUws0t7SwLaPdHm9TdGCpui8kq2vH5Vvv5t/gjNlFZ7qXmwTcWChG1ruxowxsFEX
sLnCWaUMV2Vdfo/HIXDNHcdCup1WyJfAy3rg5WE5FSi+E106Z1trWajAPbt0aXy9
feUbBzQUGfgCWLPLBa2qDEekXQkfx9yG3G5yZLpqcNsMq/R3KTeqLKaJjlMfxdi5
gtYbWAATKbozcQM5kdFeYz7/64cyDhicHkAsudBBiFBDGpkwgjF/uVPxSSrKMl4O
/aLLAIjPW4FClP3g4s/46Fyu01pYGd9A2ct8RFhOJaoJIPJFtMvzFSdcb0DtIY4k
gYNDyfWlQEjsiGqgeMVnHsX7l4/QxhTBOCJYPfmVzoUcY8Y52BvlLJo7BQr6u8tv
X6eLp5QpjXmQZC8Q9gL7y0IA51scyGhCcj5RgUwSeF+kbp6cpcdyKO8SahPbIOjp
UOxjxPEkh1ZQMgRFLueFB/mnc0bc/nnEuRShViJD3rxL8q1EPlx2lWPNyYO0T6r5
uWKh4IP2BG6w5+uRMHbob0JPuhNp9VvBMjntG+twc+UZCJFQpyprQfmziOy3bpRh
+jcIdHDdfUkteHp0ZUqfpfRPDSWmT+yUQPAvifxC3s39ym8ENFKAygHv+cZjLQw3
4jlP58CjWuINnQsBnIR1434p6Ksi3l9yHZltM7QFMnFTLDwiHTU/pScSkQNhRygb
eWvczWvQ3dImWv3OqIlnuJcYf7WhQjgyxN37aJ2XVIdPpmPBn3pnSj7pLV/cp5vm
PZiEsiYLRpba/ury+zwg+dfEEA9cPm5vbbqmQ8OQjajsatTjX3XSz17CvupDvTgv
Dex/CtiOiWd/25Tg9Jmj13JZPT8LiONLeDUob2/OJ4t/RFKiNsuyNzoPMVOe0DB2
O8asoxxqQkSbaUHyMYlwAHBXQPGArinwQ6Nrr2rR5cj0n7QRc2CEfIV6xY+8WO4Y
FDhgdPDo/ZjXcBbONOzEfNyphGgNgyqYoWZgGyoVebL2O+/SmSvJjqwQFVH9Fkqb
wzXZqltW6xqGUbp7e0I+PmA/4KaQlKGPEV6ZuitI2SRhHtJVA1ttNsFpme7y0a0J
KHX81HLUuJrj1p66QPRl4Fe5aSrBvc0DRVcKVZrBxP/+ofqEpNc1xy9gfn7u0y8C
jJXLvLHeqlRWziS8omNCxir4LUobum8dgIvmnVHAp8yq9bae1SZEwES6GME+x/sZ
kY4kPDkVVSmCUU/V/1ROjfx74NK09Ajk3qVqfMuglgzlaqLpq9J8BEytGF9UVKbL
1hykbX/JRNbEm61zEl+lhkBxo3FWgriRT+7RpyaGOu++EOGVpHsvyF/o9RdklgIH
/UjYYNpbeVWd006sLxPNHnRpWHlaNfQAfVAMN5Nvx3tMiQEOJycoCHZveIRLOijo
FIe7RSc+QWYbs4F6aZLi7kWgDG9d9XzHFrB6alDnCzltdoR9SsmeToNbTUcJyGt+
BCynXfHcgD7yjKizItQEKLIbNjrX4a9ZhDVczEGAnW1/5Lde3LM5Ugeir8DyqJsb
5jjWHtW+85wWDFkQ3c/d6pV8/XUQegSv9yCLMe51ykieRFLiuGNwMc8K2NOBroBO
Da9nkVL0aw6IFT9/wQxr5Kwwxzxk/ysW69QezjfZ+7LeRIoDscLUOl3DWM1QsJdZ
Ux7Co+YZAmb48Y52Jy34EBfL7YwU4/LLQ9VzF6UycsBLtZselp3WU4ePMoBUrAQ0
93osSMjqYjH7U2Zh/8+ANqAJbslWyqeFoaNANhsZ38XTWpsIPLqjwUWvrCg68WAI
KtMBsOmyqks4asgPSXpW4Cz3LeZGjP9pyEyYnJ51Ng5iwAJx8JWQN6uwQG82paR6
Tz3YArPkiOvpG16CxeBmhytJo2/wByr+6kfBQHRQ5eol5QRHvX9sqLG1DBufG613
Gh8+1gRICr0+5I8yIPIuCFQQbCQZFuA+ADU+2ZrR0mJibfVWqwYl8xsIK2uquyns
HGHHEPc20/1VctTdm5Ta/EUyVe+3kaZkdg7qXL7XJfgpeXT/pH6UsmSPCjg3MvFa
Kg5a9H8pFmPWYxxnPq04Rpp2ElP8ROVpfuKrLpj1gkvGV9uyOubQS9KDfCPvKqs4
cUOybYrksEfqu9YHXB8ViOIB6d6/WmCiSMsl9LHgq4RbqVRZklnoJ00GRa9XgWdE
jQUfvb6gFjcSfDf/znj0g4KFU8r/hvGI/6jKBxBN1iwpQnd4gdjKPdTFBsz4otQ9
Xu3wf0DsvY+g43LUhD/H+231/HmhtARE8es9W2iIEAW68q6cK8VK5XjG7eeiF5TB
4IBrLjnmPMXAshuevbLdvrI6SwQhvGmCyuF52lJOoZzjOfOiDZ2jy/8TrW0AjVS1
kh1DHtbfT+eRdsfnkhdg7c7QFxjAU6BViZiSzu7S0xluXxV2J2n7zKs9J1H1B6IT
GtuFZXw1lJZleXZecax7jAeoPjcBtzXdYvVpm1EidWDrpOUs9NKl4OLZvh/1wBK2
hSkZ4f9TV10bl0cXHqgTEuD6XHxrMWyWjGJgCoyIGwDK80Omtcp3FwZah782qYms
11wdacfSU+k5TPFwU0lajy2M3j5c8XE0Ep2Repc4yHCDIX0eY4JgfhU5xy85m94V
qgbHojXLr9ub28C32oU/kyjTEwQRqKRUepOAh6EkVxqDVYiEj1HQMZBufDN2uKs0
d5FCFORCFpMe8uemVIcXSMbYZcExqgehdgWE8D9r31BZ4DMXxVF+sA3Lgq7FQoH4
EBpxiXLsEPGcycWLRbKcjb2wNMwq9BDIYh0Cj2BvVyDReO4CNYSzseCxb7zFbQht
mM3HRWwGZAuOmJdANuB6xMTMjEVUZvq0FNLQJpTOQ3hlhArPe3/e+Ld9a+Oq6Lbj
Ph/F7CavcblrI6Nmqp6xuCJvrRUka+2AZnyoEAYc59IUN8wAJcmPUvKXiDhhLcvE
hafdMQcuNzQCxL6oct0p9sN9Z0KppCP4KSLnufYBJj3+wWUdi3RxXI/uCMFGFBhK
81yv2Kv7rYVBRVNW6D5g799Bg64LpEhwvbkFim33oOIXyKxrNMozknmIzeEc2ELN
83sdlQ6Mm/TpSf81X7ZF4cZc9M3LI/SlL+l7nFgVVIvFn6in57l49VlQH+OptdYx
mKym9XLINfW0zrPXO+sdqX/8lS4jZmRfqknPWSizsj366TfsMEZS+wLcSqUf7/1b
OX4EreO/7ViLGkFf2wbUSj6WHmMvOQkPKVAX2O6L/A3NXig6dUbyVDPdND/rOS3A
1OtxEVUEAk6wttr/a5ASiHVsPJvTFjPzUPX2rQEb/LkVK4GKezCINInTPmgL3byA
qYQK0ExfPa6KCQkCMmrJsJ0X56Jw0xq+N9kTTk06zhEv5jfY96akDSmB4wzYGZ6f
skNPGYLl9GiJDTRWJe56qt3JIuCY0WKvItYK0I/EHu4ZmAttnVhVoTsj2p2dCpPG
9DqWVz939daHkysW85W+M3k00HU4aM3J7nVL5DB9RgaddW5fOo3leXDcBH8miaHd
/TMvpoj+vxg7bqBbPhqxXrDs9aiaB4NnAj9KghNSt+r9/C/hPYRBWb2qc5HaQI2N
m+HcOqVLGnlQ5tkSv/FbKkagAUSPITHUzWqwEIYu1Pb2hBssE2bd/g7pjJV4lNBg
hV5oaComkS/Usjk1wgLmtNkyifzOknW0LpL8l9ZAYI9zNl0Fw9Yv3NStMfmV/Ljj
UltkfNFjAa8jM/hqyJNILoK/80DS6klkY23ATkXzwLDbNmM1O57twLMPIAavHZVq
ezZLVx66E2jDh3fSlUbhx1YBavlUKadLCSPj0OfkItjkV8zlaBq90TlhgTUVkEXz
E21JNK6qaZYFnYkGMq8rev5FYEmPTxIKmMHYz/fab20qWJb8TJ1+zsQKXtA0erGn
j1OpWKDtErK6XxMJN2Q/BFzTIztKZczF88a0cqDZVRoKgoP0kKS8LJexS4zQg7EP
/G96uWs3RFRyEU4KGXXO1ECPz63oEgm3eDKl9hFqAzp6uMbPEZPGDdaikVvtlmNg
XBmDW9gX2uGsczXiHZD0GhseJXgdzV7sTCi8vmn26JWcVmRI78YoUvrDAvjqmrol
JzK8y0xshOAojWbO/Bh6Q7HzXkSFYN/UsSvfP+78rEpvwJwdB2gQbdhFpTOwuwLW
AzPatB4UWpySYHX4CPguSgcOn6tun8y0ghOkALu+re4x3alq9ssqFITQAC0Lvvfd
HrIF7g9xiItCQkXeip1PZ1U/P7HycJG0EoT+wqe1Ono+7mRRvmCULB1CT4XVgWNv
qN18ZlzlLWrrU0q602dqYXb4TyGwTZyo0jG7ITYYg/Nm2QdhHAbO491gqqf51M36
rc0+sw69UB6HmYOClb29t3lk1PjgoFFdt1NI8MS4jw8AawQe9AB+g5wA7dJiW+RR
uWeyv9yi2zSpQrDAow4ZIvDxYk/SOgwe7Dqu6bd5H+7lMh+5UElCzvlH2Jm1CJiY
ZQNiBRW2HQuThRdH8iW3yexDAOFZ7udaqoYTVwrk6bBFahSM1kZpY4O6dLIDl4u9
BAPCFFvVLzIjpRYpZAsMzwnrJSleJNB98bKyWpAAxalqiNQBfh+PQyQRpuY3NeYn
q9fw41S55P/vLp3sbBVOuEOVUfAK5d0IxD+ImRb1eZ8EyKDfLQi+VAoYiP53zyld
HG9DIvC4fz8vojhjkrcBxVGVqQaF2raO+2tWgYorJ8EtT0Ij/6HU5MQnNcxTjjox
JDxCoH9yMIyFOjr7O/V8ZfD3CtBF6GiHbiOv6z0Qgm2GVJs+dDV8a/CPLqJVE3NG
K62hhd23rVbPWfHpeIy/AwFUM6crFj5FJwugSyGGUmO52BHVktp6RE9JKa0pVmKu
gRTrXxR4mfKOyFsgNxF6/gXNqN4qHoxQg8irU0M/VkbyAfd2s6GOX6B20UeUIK4I
6XSXnPTeM/uwu4WoTFreN+Emot02/wOTGuf3TB2Kf7kRX2h4K94HazDZ/cPSUhQ8
WnK5fwsSiZZ3jC8YJLMtTQ6Ubm9hIo2jEdhY9nRUfrE4TkTJjxX9r77RMnajpIE5
/AfqEeS2npW2cp1MIfrhHuos+cbnadpeSTKEWNFVxBSSPEFvFmPJov30haBFa3Vl
IrhIAi4ROfMPIFd0/Wc96a9IprnFBXOVgWQGjmRjsDstMUdl6D/8kyWU9HbpYrmO
D93TDwKFHsBkYDIyJAq/oEU9PMw5q7sTmLjIi4eJ3o6fEQ+kTu5owOkgC8YJ/8uC
0uVtD2jYfyT6nvS7QBnW3EFmxCEd9iCJ687d0NhoEyDRF/uvlW+5v3evQ97BFBVj
X1WBqk1METNKhX4WDcvQLAH8tVdTbi+NSc8rji/eOkWr1seumLfSuYll4Eq1GL69
u8gFfIY15O+fLBUEwkMvQMANRDPKYSSFbSiGmtHiqCT/DZd2sD2DRb82NMPs47dT
vid2Jr4knmE+yPGGchbGoI3sX/OZqEmTrUOe5Ep8yvO9WnL8EBO6tXwl9zTwNlGw
vwvgLuWVawBXoLZzM06irbklXsMCaNyaWClUUF6qohEPC/hy9DBnYkOTEikPXY2q
GKF7KpKnunhaXwGYXgKRqCnpSdJBgV5d23L3ynYmZx9Pm9L5xkieFcpHJ0BraL8V
DqoLAqGrE52b7z0jZjSyKCbgaU6g9DBQADdX4bc+I6d+lM5IPBqJl9nuhQCsj5J4
0xsArJobPbxJ741Mbh1RTrba42XCHCuvTxe421ys6uWjtMCFdhJxmZ0vC8kEPEy4
8+pws+1hZLkz4KgTY3/7lXAxB5bwXgnjPL2I0gp/lHE=
`protect END_PROTECTED
