`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u2XZm42AFP7KKtbak+vz9rfNPux+vYuMxBwvblrIwlzQW4f6OGYhmqbJprdY/ahP
timxdUCg3++LMt47p5fuF00TNa/UmIUwifZ+PYkPKD6XA9gqtCLm58DdkvUcm5ax
mNDSuYXhC2i3PCB6rZ0ttuN1BT8wWkY1TpAYLrc+oAWb3bI801PGiM8nfi5ZWVuD
RslHSe6vdeN7UELtoFh1Ymm6cKxLHLOjw+rTGUxAd4CDriIvU3vrSToTMcZwwU9S
Tam1YxFe38/z894e0Wp38FLGvdCvChFFitsk8xII1MxnTGCIPYKXWzFfXiGkFrJA
pdwxsTmJmkFmlYQ8i+96YhZHI98G6emu410tsogVZW33hskuC+4SehBV28tRneXz
rxf1SKJDS3hlFtXSGF6iCabdHV5MKJMghSjA+0oIl5dea+0kDvrrlVRR3nGOMTIn
/DlgDHWKWS9bv+QPp0GYJmTHj5Sv9OcatwzI4do6N7qaDoaoOebcc3TCuzL/P1rg
Q7cMa6Jnrq7UIWNzLyiMIs5X9owk/jUQI3W0UI8EaIMIOuXQPM37Ngma/E7TWDUk
8835Qo1NFxUEtIjj5n4czvACq439dM2xHra7oVwEIkwRxa5GtbmutydTNSZ3tMmt
IH0e3VEUuCpjlea2TaqVacJ1gul5hYN14tBhFDo7aoKU+hKvXe4peG2qMcWr95jY
mNF2Rpsr8KzKi1iE+wtd8EAmXRm9xqGvxHJdLfvJOSKkj77rd3GpVXFHaXIr3JIf
pBcV6lQEhT0ABFgMPiNFEQV7zAGuOCZBPCSi+3fSuxzoEJLjJmWFXBcXCikZLUkr
w9nm/ZlVu8+1TDcIKxrMeQ==
`protect END_PROTECTED
