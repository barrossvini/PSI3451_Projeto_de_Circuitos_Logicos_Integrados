`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXvg89CP2W65UN0IUu0GGYwPJ2hBQIQhfKDdxQ1IUq06UMlUxfL9h6hUhGdp8B54
wsViIQW1PbnlybqhXzCkeeww/QJw2A546B+rVEYeKM3nEBflZ3DudDE87Kk0CqoF
viFEVgnrRGqtzFUzRwZ9jZ2a6SINfKDWDKVm0sK5x5ZR+g2OkNI4IxsekWinJGEX
JkUDGft3bmmZkdIVR6fj8EcwE+t3s4Kc9w29yhG3JaNehT0Uj4bz8jmBaSKF5iz7
MeB1VKt39e+XO4+zFp3oNvd+485bzy0Bpi7qrRL6Zjqv3Im1gaGRrgIgYGIPfLUV
RErQmgK/dlrqeQNuwj1cesMpzktGGzQmid2j5s6JS2FMrF/AMu4w9R+cmaTrdAzh
xSyXewPRuywSGKbZa/qprH61goLUaLYRddoOxW8WcxgUlNyCr9A+Vw0tRZFNjMKS
+mMjbprgngHROPnD4UZvwcIeu0HwcYV4wmfWz237vTwRVsOCt4+0eY5R8qEtJzkg
iP71xXaWHBt/8TT0XtsRT1A1xkCurAt+ayISRKOJ3ac=
`protect END_PROTECTED
