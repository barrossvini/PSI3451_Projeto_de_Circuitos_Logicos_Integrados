`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LvqHs8L02FoiRhmV7nCqfQrxm7HYcpww/HkwALlcf/kM1xILaLHrsBWrObxt9v76
6aOx94/W/hYwdi3LQiim8QVh1WDi/Hk3mhRrJg5hD5uJR39be4QqNZwZEytu8JkJ
2IPhTcPdqgX6J3izzNuOzgzgBUq6jxhTbApeBp41UkoEv/THmmwh5Ja/1uchHR9J
NrN7/dtyUoWKV1qBKvHTuoX72uPEhTZCoWmRDAw8FGsOYnKKryCqeC3Pdv1uairD
qTHXn1Za/ZtnCNVCBEvg3tJ00XI9QMUzdMtIaks3N06LUou+aAyayXEdupa44hnp
z2chW9CSiPMmm25IKNId8vmf4qr7fAvoiXOQelCkK462XwAxFFJl3dS/wtIigWs7
YjYLK1bv+VZDMBnu0daa0riLFNJ0vkNw/2f3QCoNk2+EblT6Mo8BJD7U51E+5FaT
SfibUVmVhbDCvkM810MgOe6K6IZcqsV+l6YjAeWALumCyi2SOMtyqQKaXdhkBUC2
3a+4RMDJNS2eixogHwj5GDneyOnwoM3RWT/kDiacFro6we6q4TSGI8Erqm0LDo6A
IvD0KeIPne5OjrfOTu23STWjeTiVt8h/K2DCHWxbm2D/yHWR5ZeX+YH8ycHP6G04
MB1xjGgVgOuAWGuyPz3WkDned2l8+45GD3JPkywEc4SG2uKdXFmWwUoRPJ1L5zej
Qc3fs0gK/4P47AlFmjI4p5vxhu10FCgTCEhfOvnbFNL/Uyq679dCY8ytW4nayaXu
4SVKVBtZHo04iTwbE0Rl1Va6PJlePXw4tqIL7Cm3TfGI0LI9E98swfkhfgjLb4k0
xggSjqfSnjMnGu1d5BNs86Hjg9mx1haBv0bM5x1lvrqmZ4PJIhrMzqtfY0kC8pev
9waPSOEYNIqadicFCG3++PevQSBWa6KM5oencYg5FOGaSVhTnqlRm6C1au13SBjD
PgdypbJOwlVDCesOTn0lSPq7LTmv2fmqnurSBWH3jAlmWnYzCnWIob3uH2ZEf0Fo
G9xAmce8MllIenZdkp3R0j99EMq+E+igI2RsI1p/4C5S+MdRcKnjCLwZHV8OwllC
Wobx68VXIo6iuBXYOKcIWuUQLoICfxBlAELXWjcGEjDbhIPure1Di7/ehOo18HTx
6rG/0X2lfAm7YwbhH8DSOn/KGNsnd4B0LEpr0GY3fjTMWjb7kRsQ5iqCQMjQXM0B
XGOntQPNc8L7DrmvfRCwhCGSn96X8MojomafMzmlwESdmFHeCMD7PVohfIlR2tTP
KH7YDkVSeEvUgSt21NkcDia3J0Acy7w+PaXEyu4FOvmCBGGXLCJQJT2skkFzTtcy
h/NjfFGJ0YB1+Q0+uqh0xnrY67sh42liKh1JAuf22vdHCL+02m9q0pRvNwWsEYWZ
6o2/Y4UoYiB3y1HFtykEc9wqcFNxiCxJca1mfkxydzfqZFhlF/oXtnT4UcfL4TUk
NzAKJ8sKVTZ5QWIE30umPsYx9J7Yt1fd1FRzE5muEpIuQDIh66JYSbe/+kSPZ+fK
eu777R7l6CoyNnmyIv9Nd4e5QhkbNdqj1MKYVg7r1gsSo1FxGiNXamSuM4yI8Y/2
/2v4DUo7abBt/1mK9yjTKy93qJthWSk/nuPcBPepGcL9WyKgi6T7zpwvOu8+FN4x
dltyJ5wbpMD619lzJSTVRhDV0CgvFi4DNXw83qx0EG9Ozyqs72B2VGmwq/dDnGOW
VS/bhcMydqQdEkIPh1S0mg==
`protect END_PROTECTED
