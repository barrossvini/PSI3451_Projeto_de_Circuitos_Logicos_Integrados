`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mDbc6SRBXtx41w2WgDCl9QNSBL9Ddn3DL17ffWTCHaSTHDREMBFuiDUFJAgnfnYb
m5SaoyXg6vHxNXrO9CV7tpP974ukT38l8iOa7Ay9Sa/X8OlMDc+bWRBY696EY6vY
zONcsuXFcqBQ51mC3uE0NT09DnvccKH9DeXL6Y8Z+Zx61FwQ4Qn0HSvfR4c5i3dj
aFSjTqDjYm4e/l5GeQcEHMKV+0MzHagQ0ZohosTNNEEV58qY1E4GTl6/CpgQaxLg
Fa/p36dzK4c1yjUJEdsA8nppI+S368azp/XxGW/8Y5LpmQhtQmuzkg41Fx+B3TYI
tim70kF0r3S9UJ0Tt2aFvilmQqFJtYat//X9CaTVe/eiTTu5jIKJ4STnZbU7UN7F
LD7a+Q1evm0SiDCom9YxSAKhNP2ZMW3ruMiPU6nP1ihj8/tCVJtAVury7W7nV060
80oORCx06i7mr3hj8ITOXcLSIMtfMmziwvFTzkn0Ce2cAnilyDjEHdbGw0kE9cHQ
acXJmx7cw5R7izjMH9V/OPG8xqHPx3x96ieyu1+SYHxPfH9U52Ps+H0IQf/g1iRI
4zi0/EapcPsxQiVQ3tiETZ1sJyh03rmu501XtrMulyWT47bgP9S4IG2zO0hRm55T
7s7WgdoUrnx9560QdFzNhzNM0k5vsjgPwLdPUGQb0JRZQqYuSL1JxOxA9az+mgvM
OxxF15tpTvc041k2PyrmrInAq/37TeyBbLLSgRcj1ROadsa2XH52zPG6hdZVnzeJ
7Z4pMqlotSbpHomJUJjn3cz3wx4ldQ01JlTzG4e6FrJiG0MczGYp4hYakf110VmL
Ry+CISGAwj8hxICB999STDincTUTV1I3FuvErWdZ6ngkDBuG7fFRGoeIjw78bep8
K2f4WrGRb68RD3z3US6xIHgHrojLqX5gxy3yIcqp/BjEvQWhugMaeqcvcL9VuZXg
UjHsfkXju1kjka8LFDzydh8YsYPxcsCYhxuvKF0KmAZRKlUDKDcEYacsutBpthsD
OMgk8QX48dCMYU6VtZpthOW9Voo0+RI2EpJCZrWlCGeaWMxmmz0Ua+hB4WA9bjgh
EN2Ol4mZqITnPEyYqvfl/9Rb7WmZ050hBcps8o6pSjBZd4lSc+K7ZNESYt22tLk3
fjnAY6lyJnmMw1DHLPGPncl8KLe6X6s9XkdZjRuX7GqWTf1+uR7KbfSkkBbH6swb
R6OvJdhE84pXrNsaaHzZ4SQY1QtWmfQmbhcl6kVFGkMsI/pUVXPkwMzKG1jte943
f23tjuVSMwW20iWQtVxcJqMw4DGY67SQNb1wYj8fVoE71m3ETzPnX93ZdEgQ30WS
pp2J9C6uviFFhy9zhUktB9/G85n/s+Q3AeKU4qpAOSk=
`protect END_PROTECTED
