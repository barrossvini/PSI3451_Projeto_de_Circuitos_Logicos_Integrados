`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mdD4yWRW5d4/T/8MOu4EvAORJ/dvyofOGLj77vsJfZRgBT8BKYT87xVcHrceqkPk
fgcQVqu8ujFPeSkQ7H8ZGTEbLtKb9+yQvnofG411Bf3qLKBQgSgb2baI/FV8bYVL
/2skB1vJ98woeg5DYKv1hXg1adXQCivay9pUQj9GFivBOx+Jq5rLlhh81Nr4+mn7
K+YM8X7sUsrBmYApGgpwJ2pzllOvYG++2wNpDN/SW3ho4I+X1z8O+p3o+EUmwGLH
Rtzf4CEIFduAqRm+CbPwvL47mzJWSdmWnb5TR+OJ+0LaFwocXw1ZLG9P0ga2yYjZ
d9gSZHijTRnrn3nuvzfp52H6ulwkQg8xa9JDubg34daqwf+815NlIB+3tL1QODD7
+NaJxuevBoFTYPtgzZJIvfQS1OXsUO7CHoIMacvh24k6TYjN0MCJ1lQR8Y2EvF8X
QtKjaNzL7jWHuxNcO3jbt8QnGxDyZg/IqLMfIBnZwzmsT/zo7iAuBeT8onDFtE2o
NBo7ksj0e26/joa5CZKsMyc2F4F3rNWZ4LD4hfwFPKOAplR7DXMHh4lX1AgoHpm4
XOqntJtieMO0I5iPNUbGQZXpUdPuY/PEYgn4Mg3M0h41Tobb/lKNaorvC6r0vx0Q
jHDWjb2PAamccTv4h91LQfH5qPjE+56TB2ZZpil/ziUBvIf1q8aayQN0N6C3UC2e
akwV0kh2vOKnesvP7nI1pBlWDl+FCij4thi0m5+A31aUxrhWJ1oziOo2oLtbn1FM
kpFJXOS0GAwuaR3Fx7gu2jsGBSW0VJQMzhrKjz9BPgVPc9dX9idFRFEn2AqVm0EM
IADxSaYjDx8v011+KpggGqw2r/GxlFkkQg/hr/xBJ08=
`protect END_PROTECTED
