`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nQgAbayPW+PDzaOJD6DWQTW44GNq0hkRYzleFlSuFo9O7Xigchdmvcv/iw02jT8/
5sxCiMzcd8IxJxm8ocJdkmvIOuCzUSr/8TpFRVxNzKcQQSw1UairV7Km61Zl/pT2
CKpyvyVTPB7snP3AsuJEnQQV9Id5twf5uH4X4/EcHMi1MuKmCPh2pippYC+euO+z
6zpfG35VxprTYKIMUfbtRvnN8131ZVoZOA/eq7qSGDQgiri8R6UM5QTNprYLx4Jf
53AWt/zZBvakG6crmEwaHWdoxkC81PKP2unkp26ezqaWKhkrAPyJcKJUfj6yhbAr
13JQzv6pp8hFiEsBOJhGDbaryIQv427yvpKQGDZS14JlCFf8UjhLrmJmbn/T6Tfs
I2IMGa8hCaGxzculOxPnKjEMTjcttPHJPUkc2JWRGBCaSgatusMBg8HAKq46vfsW
AUFFtFfFNw/wxpQHEEThkSRh6SQ3Q0RFYR8ajxwpMwy1F1qLZUNuAGkbsrEpNd9C
ho9M+RuKaVzw4ud7OV/K4llkNRhCEC58ukwxCMdmiABv/Ue5Cw06vw8PSDkcNPH4
Hyee0FKwtj9LGk8iS6zBj/63x+VS+v5MPS47dxfxtRuosZDWC18OpyHMgqTzJdG5
Mc2HKEv3Z1elMFXlnCL8r4owZTtiYFdwfOguy6AMBUExSUAutLnuVUiaWhpViy7F
TA7HS+ByBh0L16CTyE0p+oJh28GXqCqajJbMWMt2iVKWu/BQTtKK1yvXwKpScwVO
78Y103lIG6ehAMTikRxN2sKVlzwnGiH/sYyIkrlmEqdPuYEVVPaBXa1YVdQudOwu
hJw0ZFXjak56RW7gFRvaij2Mi9G/5HmO72nlttWKVkofHfKF1ap2mgHgsyWdRGlP
zvEOypohkgxtg/kqLscKf5AHSRhiLofqCMFI596V4XwshGL4XmaF8FauXZv6RYJG
98l+6I9wdOsravY+TN2EB6hrwcCDQJmNcUY0IDbtp/RQZmCR758raaP/kasaUlf8
eIyXZ1kti8GkA45IOTDyIilJH9RHJBYJz8+p87YVILc1NNf2hEJeu13QF8bxhw7I
PPOaWkPAutFQTqidz4N0cOIj7YTL7K3s5T+VCfIRPLaO4DzQ9QLB/CP2go0jOUYa
qYYE6LKr77yWawPeOoCWr8jLOLl8W6kWhVvoPfpCyhSisH+XFGAQbwUF0lfb7dTZ
WTcu6FQnr6umoGAB1zgNySsy73Gs7t7jhWBZ3KWpNm2EVUOgf9nu5eXbsREn9BVB
`protect END_PROTECTED
