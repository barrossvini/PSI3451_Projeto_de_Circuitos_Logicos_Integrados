`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yTC/sIijB9Etv8pWJGtabyQM4w3E5et+XeH9dD0rnyiJAdZnkoMpKXQ/SnPh/1g4
dM6u5JgREchHNBEYhCRxlNSgAcxpaCYn9g6dL7GfK1LeVYfuk574S6t0tJX6Sam8
OY76C3Heblk0CO95jwDTW6AsRuKYjLMK8jsJdr63HskiYeK2VXQ6itWyUexdiJjI
RIBRLAzUPEqelRxvMCzsuJHIuAqZrnzwC/Z0eayEDoz7dNWGw46oQNhhh+qDSf01
MKK+z2p3DuuN50tNfqq3sg6Sf2z93bgLxDQVYqCCob0Pat/C4I/pdEtylxR3anEo
YiKWe/xYu0zeWwASra7/TUWKmwQyetIjCkgwrEzoNMC8jX6VKsJ+1NFV41V4tiNA
LKy3LM/4lFwUsAq83b2vxVPfIH20GgTQ9o4ECy6K2Doh+FGnnrVjXoK1LvVWhqMk
N90KDaBElGMfEKnpCDPuJh9eUGPxUHgBFMiQHZfrfwjmQ76Tyc/RXd8tLVQZnr8E
Dk0ynVgFwd+5nE1raHfFLtaYwh1i3Dk9qnXV5hCqVEv8GXm7/3kiSE95W7ihr4XM
fKDtZl3i+Rh/Q6lj9GaORchvgV9VCuU0F2yOMw8qloi1TrrtZWt5tjEIO1NWyXsW
urYHD6AM3+FS1lAB/QMXASHfs8dN/1rHKbLv3rm9SNyqJEAc0j/oX7qIIclkEKg6
oPIcEVZ4OqT7ZXTzPoo7X0GF3dLoVRoxzIA7hybtuywRuWjTOgLXF+I+vtlSEa7R
rq8VtQkeUID8qJlE2ZHKs7KMjNHrI7rhP/GXLA9js/EkjjcA2+LtF56X0F4Jb46I
rOiX4v24H3gU2Jqkdhg56S+1jVitDbN9GelBYcOzaGcNoR7KhMBzoR1ErK4tVakn
Zf9qWHeTH9/02BDTg/Cwx5y1fFZ1I06knEwhbNj09NbAxgjgkxq7e6MkvcYOnXnn
F2GTYmTUspFG9g2HVAgLXKFm9zu4esojm5H0SAtKtZkQ8rrlPimEcsr92kxfh4oK
JNkQU5Vnbff7UKRM8X2oIIRRsM7dLLJzETH5NHOQbTr7/o6uKYNgWmKPa0z7Qkbt
0T92+t6SLibTe7gF0ZfnLWLVjVwqad/Mzn9Cik3SMRv5MEJZ/5BmVNMLESyOJhVS
zgONVrPzK9Nh8tgUBnVJqJnNa1JijbRdngfBJlLFCaLtlyA//Y5I3W/K205l6njp
Fmf9I5kVTuTHyI6Kqz7LZSbKC1rULENsARyMg0bR390rMZFlQ/tShrgArsy9MU9v
yfYbhnanIjsClgyEgo+2Qapmr1xPNpifQnANouCShgsbDgRscJPOf0LZ6G4HxZ/n
cfq40X+qD1YKmq4LJrCynjwhneMAbEuGyf+QJ8xTFD11aWpykZUfewQIlsfYH5V+
44/l8+qS96wrlAjJ42fn+TqaxVZ6ZT5kZimHzQEQQ2W7+aobfoo+LjX4JTsimKBc
9+qhP7NGHVsN726d9KqzvwJ6FUJvbWvO9+Z/5BsmAuznmPAhHyyYrKOM+nV+/qTC
gU/M606M0zVYy+yUqqmmhi6x4Dx4chfLruGbza99cuMk6ynBxFSLgu6yF5lTs6iP
svCcqo3dYZfPOQpeuC4jhVYNBAjffhSJJmSxZqORPHu3mg1OizMUVS2HRvS3UM2+
vT6niofWXMntA+iEJSkFMxghLM64E4csURyC6EYyZAkoDcux/57CoxMsqjMPZ3Wx
lK7JYm53nNsZv2okKzdeiAR9pLbnpnkdsKwWZh0EM744/lYJNBBJ3vG/cgO3F26y
mUHzyKSoC+Q9d9c7U52R4FuJprai/T+g4/paO6+evTBX2au2FF+Uyv+2dHS3Qmwg
1sG9PWfwZEMmER7D/3eFw7xj8wsvgSx30oL6Vf6z+gGNyPmRWujulCK71MnAqcmy
98mdEYFBZAkZ6siSLDpbPCWc0h0F9okaTZtOXK240y3EmUzSJ/BI3WbY5JX5OKnu
wZZo8xhRm+BROEu85hFLYryHgPssLKyOp4ndUBHfGP3e4Zh5TRNE5A+41cBbTFSr
8Cs0ViVttOoPb4HDKUKFf9bihDaWRwMr4FgD9TBL6ThoWjWgFt/Ii1hziCZO9AWC
Tuls+ovdyl5Fo0xMNEaCxXUwtsO0Ory4PpORQT+/Pmac+tz1Ue5lYUFgE0qhuYAU
CTmWEF4dC10OGy4VgNSspHia4vLYf9ngzPqcIWClZxj1lFrx50BjBHGejSuSWRzY
vZ9lyHKnKVDvdPCqsjT1DcO2v8Tiz+/Lb2v6srrzX++p+7ulK3GPOy/800V148be
Aux7zLV55w02lbqNCB7fW2So50U76x/lOZLlY5v/LpH9wHslG545u9AXvRpxdfYM
RVPgzcVaHxPhJl/pvVyrA2dQpi28j30p1Vyfo+ILz/TcU2fluFo8BK1JIRRzgx3h
f6PQNy5Wf6c8OQgGsSgKc6BFGldHx1u02pqZHmVqe09R6xR0ATSG1qgTkeWnd3xe
yvUCP6G9gZy42mnmd9a/FPecILERMur18fLZZhNTbTwOQSx9VgcI3PB6AkePfp0u
+UIekWAgp51IezwR1VZ346ItAQm/SZGVJYtdNFF3gUBnB0lF60UA0GkiK/VCt0Tm
nCCtMDuJlXPXKw4+ZI6xHiEaaOl6dfp2FSK2wwT/uED6Ce/xzN0uT4CawzIZJqnk
glo0MT51k/h7OQ0USbVRzuxdJ45xxjHa1xHVyZRtO2vBDnSDMj+WXUXwAb6hDraT
ndPzzhSGqpjOmtkbxj7br57JouN988Oi94CbQDHZrC4kA1x50QQPIEXdJyYTWeSN
h43B/Rv3fgnovrxKGnqjnCd8hti2mXIUwWqGdBY6T2KXyB/1xzFAIJcO/6bF7bxi
2Q/PkFL0+4Xl5ysxqEC7fDPGp7TqUA2lrOmQLSeBq0VExlZEktm2xJh2PC7QIux1
ScBSsVVF8K2wOpwfzA7e9PIKLZblfV5c2DLTpMXjtrWrLk5DkovDjf7tB/sctyrP
VrS5kaHRL8YzJDOpYpckCwUrAGdtKOWOYg09JKtXt+PW2s4yaEeq892AwzVbiF9V
UHk7mkSUSIbaeh6jPFQE6Lf2ftkzFJq57LAi2uDm0GB/HvYLnbTibAnRfKRBNE+M
DiMnHG8e4mQyopQpTNbfvRQhvLnGn73WfFvlmFcN6b33PgqBkwLUV0OiVwWuy1V9
do4mFBc+xpROZDMN/m8b7iWonTm9LFPyIgkVeC8igsULgkGDWZ+rU7dcXuW0Z8Os
w/dj467w5t3O8UZGqQcHBH4rmDlMiQfnfRsXI0wkOX+ENQz6nS3OsNXYknbECIBc
1Q8TW9y4bInJyzVju8zpXH/HFcNNWsmAvkihK8oBCcChIvMXjyqP4Iage4tSmnmM
K2R3Jqql7LYFQl8q5VHER9WcjlNV05/L+Vc6tAvZwdSW1r62p74aRKu67Mu1aaOy
Y8+0Lx780BPfZbFN18d1eg==
`protect END_PROTECTED
