`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zvD7kfb91SmnOxs+5FIoQF5Je2EFcpgDFNdrgJBZB0mZ7Dbfq5S6gWVZMK08vaLF
zX4UJPv+ib5VdihGv01Jz8fCYNQbh+O14HPPajVKYUExiGJDKRSoTBgKtQLoGAyp
I9RMdGWttadqc8pZ2wsPI1dRaYN2N4toD1rqMWJJmqyW4FyfiKgP0WCh0px3GkwG
el9ABy6ckSIIHb8qK+Cpbn+RqlDQOKciv4DS0Yfki3TtGkKleqankQfobi9Rq0x+
ppKzZHXpRoqfFbtOpbKYQwn5G+MdOhkmX6SngqaOLwwppsZYcW3ctm7Ea83ssYXo
JXYv70ZOw6AXSRipBS7smjsEMvgMCIWdv2yrqA5LNY9kP11x6KS9G+4d/9XcWYb3
+U/uNwWmZG7DLBYOSzjzFtwZqU3bGCXZEDrIsZYOWJqoZ7UIAosQgqGatFYef7r7
wSWDMT+wdRNuwRbmCBDwyvOM4v94OA6B9jAfIRTYCMs0sfea1czLCmhCX6Ds48Ey
RfENXGex4YY0gxzusn+1xvYDipTfGQ++bV9rQLz6Ogj0FM+Es4EfWKmtKbyytwlU
RaEbMZfOvgAcDTT42+Cv4+xKe4gW0Eh7NPUrKWMtbA+ogqG0gazwNdbqPpNluKTX
2FuVMglgQ9Qci4OjRwrR1g==
`protect END_PROTECTED
