`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+GUN8lGRlXqGxB2fn9E7UPqK5jzlUncxnyvD6fRY1+qtO86pWebjVRwuPztvNwNO
NsPDFXmriZXbPC92FMYnV6Okv/QTo4NZmh6GrJ5qTSRzhpzmutyCwOlwIPvIwPdM
w7BT0lKdtponCWnFutLLjb4jGR9s6QhQjEoQMlhLi6l70Lusi/Kb3SK7hT9kd9eg
UifH/6boahYflkhQ03DdtRWzNkKMMaw265tSJzZ99EtkishZ01F5tnBe71zBeaqR
bIjIh39lYqvcPLJvleXEo107WVHK77WAz5zW4qlJ0RhA7VO5xpjJXBWrZRKfd/r+
EnV0uZecQS0biQYGdr7/4PLOAJkyo3AsddFpLzP563nm/TsAQTR5SDNEu2RRLF9X
kYX8zA8OiauFtpLVEfBV49jEEJuNjxMI7QF7LyixG1RpaRIevVUFEQlgSGU/nzTR
wThDsj4N8+fZAHv6LKIhCgXGzqC4x8h8p0uWJTniq71OW5rILONauCz63nSETcw4
2J+jmzxKOPCS+MVIePFhVdqw3WWmFEghBVl3mPRZKQU9BVcYUJNBRQLZn7Bvvj9e
srmS7wzTCnoya1CjcxgoY3PtM6iDHd5fL3qjeJ0bprsaNOezlXU/+OY6Toa1CK0D
MN8W2oVHFFKjLA+Qu8nGQlb+oc9m9mQuNu33eUr1MKG76VUjGWAav/Akzv4cycNC
Li8FKVDQpDkrpFNi6zUZAVSbiGwtU0fKPcFpiS3866Bmtanql/bAI8Ak7Leh6Z4p
`protect END_PROTECTED
