`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DD7Fyg/gTtk+2Gk6n8UU2sPDOK5xTDJKSRN1/Cn26joky5PhIBgVsMPvQBPrBb2E
6ISAljzJto57Tb5Wa91o0cC9acDimJvgjPH/IJRl+HxH5TPopRhmuecFEl/9YrUu
agLaqQTlW0giIVafP6I3nzQdIGEX2zpCukmyar8xwGVuwO5ajZh924i+LpB1Jxmv
eVcgCUeM1YG8HqS6vCKiNesAfZHKqX7JOg5GgDigEa/EmKhw7DMl2h0xaQLhr0DM
sn+jmoPB+eD+mUZEgOQVMtVpfsUy1ac0fhJVn41UlUeMNjghFbXzjI2ECgq807N9
JF0YNVtj1tOPmapSPYrZPDQcFahQeBOvJVAm5jUsAL9lKd6RFvrrS7EbhMtJPJ5k
sSZz+k21l0+9AX5948NrjpIpK9nf8pGKCrBmRFCcbtdRn1j71LhFzCQZM6dg0PVe
Ur7QYykxrgTcewo7vY5KxqtM1/VR4O16tPyBEblEVhoVq7KxeGhulm70lcDSLPwu
BzihN4/JWV+qkQS8aUwlnfhSw7TPwE0uyv/aShLjwyAS1BHFYZeHAdu7uufptEFL
im1bQaZwDeTYIRsqYkHn2D/QskKCEdCGSGOpE70i1aJxfld7q6YAfqkdHAoPNqAf
q8dNigA9jPRu4MX9te0vyR9pDppkIbsJ3N1VjIMJuTzI0xw8pF4a2wqsVpe2M9NJ
9yUB2zs/AlXmrMbjwsdEKp9eRX3np28BpQ+wAubvp6U+DLaCBl9liV6weKhx3LTk
Xwje9s1vhDXbWxl968G9f/6m+EQhTBY4YOTAqDXNBfY7WIgnpi97FlNQ2L2b6NrP
9Pvb7UPUeUjf3MqxyqzaDvVGKE2SNFcaZQYYD1/J0zegXwYP9I80M6aHDlYjjqFW
zfuhCd+CpBSlBoIxJntoga3rxesp38xGBPHoW/19I9sac7uk/44L0pmvziSQ9dnI
HFRCpWwEm+ocuhVasjIZjRjk1rtVaAwjSr4FIUMqtOh+gzAEQ0e2BaqM1C3i9rQZ
+AC/TK/WC3rgGQ6bxnSuFIhFckRPruY955JttG/q7mRlkMGgX84TnCT34BHO8l4G
PLa64IccNwjeGTNd8EGQx5gBLAITLq3IKLBarMhQwRekzFgOi5Ecq5QkE3swBCE2
66TFGF1pb3suDtb3uBUoa1o8sfr19xZz34dgV5PL11zsszOSpdQKuj4AlgQ1gf59
g3OuiI2/XTb49808GOCKm8Im1Y2zlZT9oBoCtGihUJOBFu8ah8zCpKQtfx4yxcyJ
3yC1CbW7CoyXtlHk7XiFkBtyBCRUr6x+7TD6vmX9vV1BxLogIl9yubImh4a2lojt
DB5qSGuhTmXlj2RdNjevAE8tWF2vx6to3lxKQ3wkDj6LNenneYejBF5hc5Z8M/bI
Fwa7ZtSbs7AP2ZI718pwxYdsDSwQrk2cA+qKavS2nYHCTYMdiIfoXkgn8Aiwy/Dq
Y+dTD4wDmASSz7ZfnKDDg+DZrhrZb6M1GfWDms6CjjDGO/L/IjfnFZn2aBHAU9J4
v6Yi9yGpkx/9VzXRCB461r0dN0VqeNFtkUi2ehmflwC0zN5GsWPo/DyzsAppZoKT
wZq8zt3hew7RVzwtJZTQPJHhKmPa8gVzhMsTQ1aT+4tcnuWlK4RTH5ZO5TI6m6hZ
cBY2kgl/d3qqtfBB/6lxstPQqLnwvj7QXmU86VUmFDcSr3MQSiiXq1HNyN3BoJce
ON2RgMY+oy8E7eAav2C77QiSkJ2C0HdZYTpaFswEQelCxTdrC3trOv6UFi4vFE1w
Ixa1cVZ+z2XHw4dqqWhvQT29r3QxqrMawjYCzQqJxIzriTXc++1E4JN3qfOetIzO
ehJwPFTMYEl4u4lG5NmaCCZiNLrKJSFoLAANXZKPfar9vooa4d8WaFUPB6NrdVGd
tiRBa9eBGEFRDyFuR8MIZBaSc5GcafFBsLUQT7BA14xQ9OwNZJd1gJgf6BBhsvF/
fr+vni7dxZ8Je8uWyP0FO72sJq2hQKEyD0W2ZdZ8F82SrplKIr5UOcT1707Hxu4N
IORRfioFxJlQC45muyJmDVNPFf8dxT3nhbciNGS7k+TdDbnawAMIOqQU1MBXGKur
0VmhVFfQA5VbTtbzHML6qqV1kubhDCYWB9c0XqgdWQnFB9R7/+F02ZcPHC73+L3v
h3pDkKQ2cH8JiCTb2kDDIM57YS7wLj/OQPokNQZSgyu72aMN168Yyi2jfDkWLxQu
VKMLU/Zw1GbUpRGvNki1eswrM6XGb9/lFkKkWKyDesHoK2et0uvqu+5nsP7REXfB
BXCh51V6I6AP15cEYdIu5klihQKrUiKh4DQoE+W6PAgQj0mhStDcVT8giCtWeyWg
VghsY00esjcs5FYiwaleBC3fT/7dlkhBcZhO8cKWVSM+UYZb23FdOc6+u4xpCybH
vIXu6y5ZSNy3vDlCmlBMGQN6ySh4d6voVWu8z8phhA1DPCnS6dwklyI2GHQ813qo
nhWeJlBOkK0a77zLMAKpCO0NO2/IucW30MRQz2XKqfmhZWA8mFO8vxSM+grmaVYq
QUEA5ythyqFyTSTPNWwJ5A+6+rEyQ4y2OnB948XA40syVWjmu8lR9EJrKWr+eUSW
65dR1mFgZjFPALVJ+/Q0j6Q0QJJK+LMHwVClsADyBvIl3qp3pzxaS8ZRmOhTEoud
OzqjLBgr4wlHLAV2O9/lMgyj5zaHTT0/FZGf54QVvr8Kr1ZygajjBjM2gifgUyRv
w9or2Q8nq1Cy+QpbMtm66oxFBcyA1DU6nnAW8t3pDDo21N5WC23BB6dBD4ykGSgL
ry/Ii6kZYn870eahCQuRbk68rCVgXfqyUuaY9x+Y+zBf3jjsRBJuHYtLyfujFKQN
K+gzV1XEDfosLskZ0yDI6qVLVAn/3Ehh8lE4btH6GrkkuEmLECPMyQUQM2GkOtF0
jaxx8pU68z+5ES1uUqGPVbCq/247hEDvgxOJ2YRRe5l8xDdMA1gu2JLDbEPePVaY
JMKNizqN/kX8mCocLxnWztU8Q/H0xZ6LXmp1w7lwSBJepPyaA5rr6hNHBYAm2SLK
BJpBOtQ++F8w1MgDyj+1dxRrLBB0hG3cmwQxoyPEmexKhZ73Uhse+xwzLzqAoahQ
BwfJBhw7VUUMzWOEseJ5gHU1aKYWyforC5VwMotH2bThVNZSdqW6qON5vdyayltd
V2ewRBPzSxDs7v/YFDPEvaOMHGtD5N0wj9QE/9l90crrdHLkVwE4TByI0ieis2n0
Gv02VJfqSf3AJ5Ch1MKD2xykNOaCgm5DXK8/TPM+eUWKWGrTxlGAQL+iCWheY4yT
SV2SjktjxOFyF5kfxuNt+l8V5jegaAXqVOsl5+TVEZhbysQgnSdE0TyNZFqW7/3F
y6SqqYub86roEZtgUTxN+eGDjYuLnLP8ksD9rPpb8FCCGXPZa4Ajbt0OQNCSOvwd
snwyGExXuWUOHYEgrGKVWt//7JItZP4ws5jDahm0nAq3LIKqI9uwZSkD1J6Dq43i
Q5d/AsqdkIzcXmOaft3PxnAgXAad9Z2g5YczHqBfhNNRXecV0ePRdtoVcbsCH9Fq
q/nDu9UPDIX2wzyuP+3/wyPQ1sRaBcezkbBbQ3Kv/9JGrUH97Uu9UnPCASavq1pM
yAoPn+9XCo5qDGu7vuKUcA==
`protect END_PROTECTED
