`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KdqCxA91fJgBO6MGPIqUddRgUlgVVpnfzC3sEajFzA5FMWrZT26jOnSseFL9xnhT
22KPq3D5UjunfWdgD3n3H0HXXKISMLL1Rs9Ym6AOQ901POx28OELHx7vfzAwilNT
rSqHdPvUvZxTkKDzTggyplTThLd3YxIsSPXy+Oqmo1Mj7y1wTrgfaqweX6paKgXT
tp0nn9wKy5RxJOIygL5PtXR/zIKpDStULgxUl1sVFUr9i615sykR8u08IvC/4d0z
P56HFHOdthAIgPPYqp+ja7rpPeBwRvdMNIYBvLcR18PAmKMrhcj68Lg8ICd1BjeJ
0GdAt3kzHZGY0lPJ64b/3YqAkX/06doDVQN+Akn/Lg7Y1CM5Rr9nojjriatdUH9L
14MnQzkFPCpnLjOafgaA4xDiC7YZ4rp4pAVY3hJZRW1SaMh0baeIuo64jbHLhC6Y
5rJx2KwRLDqZRllZ5c1smwkphmksmyPTRi2+rQkrYA2qSePgVMNBKb21udmVXsEf
eVI5opdZTDbeDW8SE2LJ7SVsTCCfySyrNye82Vz0nb+lELeix424L5Naj6zgeV8p
p/JEVis5EQjTxDvMcH6Rt5IEuxuxzFaJ66eUNBge0HQpcXBagMtugqvlLkb1IhMf
lMvJiqi44iJm4K14jEmhF8ABU4z2IMMuHmXRDn6T+0zaTI+Z8/WAkcwtzHxLoa6C
fMGJ41HPBPR5W5h8aMu4A2205HQj1wCQyQQnfLEbPms3g0syK7Eo0rpeWzMX3ZCe
Cg0OyTTdWINRKDuMDtWKC+HuJDBSmPNWDlONHl0Hs6e+fQZsaekoGUgzFfLAQxdp
E6JOLDtnAXZIhSiPpEVXHQHyDjzzy/CG2b43IZ/o4fefx6KHi/iUT113mUlz8c+r
hbv2KzxQEjb3xu8n3agGX8WECOK4a7hFAE1zL/Rw/mSc6z6cx9JLvGK9q0kBtUgn
/MvIyMNDk+4r3874wEMRFBUCCMCWlV9glQn/DMFWWZsABXidYt8yl8XTtsawumyN
HVN/S/BCMAqQFdcWwrK//mPmniF/LG45phwRnPs2zPDNZtH3996Srnb9u4oRW4+R
8ZljjowDO7XTnPr3lOy1ombLtR+fFAz7pf+qVmXcy2ptqMDguBbvtjVkAzS7tMux
NiGKQ4Oxf1Vb3YgH5ifQLzCzLqnNtwPxsIRkkIOVW7BDeI9DoDAvjEmsNQngdwej
Cj2iSDnjlRrdg9isoidSHRHu2cCu+sVsVztxsb5rq/NY8ccJqR7IkIjiWVyiuo0S
C5OxvcIUW6qUezDlXFwAmX0TdBDUU/amOatoCBsvngZpAGnCnfLL5RluPhOKMUKA
/Bruxs1V/pG6BUvE+fvazVu3Qvh6Vzl/xHzn5jfPGtaENZqlxJp3AzMBif0trThi
el99nm605MoaNm37kQXmzMmhWCtbrobp34pO595Ik/g/+UZDVYLJy8jaEpQEGkbb
+dxs5R460bnd/7ritmQrVltLcaNetBhcCG7lgRyEcEURcasxhiB9yjx9qwjgFYzX
QfjUvitO6Uqq2IE5xaic+tdoL15Be6LtuOBnC4T2inhpA7+MotA4EHh9za18db2T
oTV30X8irg+Q9F5C5zFYZJVVwutfJy4DbbISPQVJ40I/3JvkbqNQd7gYMtWVIG5Q
47DPEB5ApzM9xzm493CRpZPL4Rfbk//Yn/CN9ZQ3jkRadchsN1lbVzxUyhcs8Khz
d6cggKWy9+4U57QZOjHtyEAlzXPKid6gEQnr/N4e2CoMWkYvWOUGQafukaBcbpOt
sRGEmspyCXW/iuMsxhUYgaYf8J7uFThzzpo2mXCq2cI9eLyUshad7qFygoPjP5GP
aIM/BtwMayDcqJIw69m4oAOHshzK+U7FjXK/zvbNgyLgpxM7L87y6AQRlPpykzWl
fIlWgvjRQ2F8v3xKs45yAAUGcFK11cRChaJOU3EcDf8aS5Wd6Drg0erilL6ZEDeo
6Vcrhjkvz5Iq0WI211aCZLn2RWtByBDEvab6WzX4/wSImD4mGyMn0u/vSZ5uGvav
oh5VAVdlDllAy3912O97evJEWaNLnItSlF22xhC4pdaju9LZXh8cfSFV1F85a9/e
dobP5ov9HDdxadnguGTcigrVznYA9DqnFsQGYrsxkPBkJoDl6sD1/ouImik4X86X
W7D5+DQ86WkuyBKo+WuzDhdtrVjtTv+zeKCicEnAlKkv+Pi0sDj1nBCODDsjkm43
5BaqegVTcc2dUrbTqXjkEOzOJcRaB9tl259+yGVxCE99u8wzpwToRX+DCYZm/sgT
t7vBrhkRLalqIQ5aa2Yw2K+rNEOSjubZ4lcbua7VVTzRxMoCoZ/2OWXILNk0x2Ec
TGt9581Cs0bwRvW9j0hJS2Aa5JK+pMl6vrjTP9f/rbC42WoAZasOHc4CI/kbxQyM
X4LRIFJDaupjVwCvHK6lkdvGyW4Tss/uSgLleEkanAGB9ruSdg70CgTJjXrChy0Y
O0JLaH6tx9OvXC8TktQJe48T1KTylDW1C+sAG/jdbUEpzaUNqHsg4ctxFOGw5kQx
MVIRnR/3lLcgCOucagCilUPQ+0bA9gyR6atNzDHDp9gPqQ1/5u63X2SFfRIYXM5X
urgpeXramGrseJ8ROVQ1L0LvFoRfcTrufC4gu8kqRLIqH3UzNOIzYJkKHVU9H3Pv
5CmBy/ak/01/V/9JUQsj5ewHIIKDzQ2kHUFWTg1JUlKvF3WFmVwRI+nP7OTE51S2
6+8fDse1tVjrVB0zc3NTgXGq26gZFKOeDbzlPvnD0pxYm5tkHrf1eaInInevX+Ul
qX1cB6mEMl7BVlPzbvX/w5a9W6x65RY/kcwPBJORmmAaw8Pvkm4goJv521agFpr8
HjV9Z6TOmrUKf3mYm5m/csh8om1W/NT7+tMHXhMpA9T3YaiQDWu9HZ2Efr/8BbTQ
iilhbNridetTAYY8qY1WuLi1H+LIivgBTADUczu8wP5i7uMio7+CwSeDvv9ZqsFl
EZZ9WM+MhIxT+uLi82NxUNrhWa4Gq0y6UHovgzH08990WjDkZ4j+ZlaWWgedW7+o
rIo4YDAp01NruuX0LDCIS0AL3LOBTGWMjqAP5q5PK7hHKkUgpJ9PUuC+aJs7I8pX
JpWJtm15jZ9YojmZ6REIzqTvSZMZQ+/S+aAuOXtZUhNJHU7G7se5iV4TZm/XYIoo
wSLZq3ZBEKhjTDgZ30STLZNwN+ezS0aP4ZRz+a02wDEVloNDB29cCZebfkiWC3HJ
TiVXO8qDv4a2SVO4O85cyPWBjbYcfO4/w8JGkSUJqVXtYNkaR+aAJHEoLktueE/A
eoXDMVfBOjDyoYKqwIUS40NqhReNrSTaYnmvOhStUZ7tABiEbRjh/mh71t97dlvh
V/Q9eIlhZprZNewydyvhsVJqw40VTiJAal0QxorDvLJlyJcBbMlg1SUwtESSF0xb
EGuml7hGj+r843xqhfsGkUoPNc4WM4BDs9P7bjxRfB2rdD22V/uZ8KhV6Ta1a0sz
SOpK3MI4LVRtPQ1qux6x0pYcTtrp42smToQ2JHhROYZ1fYsaYGzNWjZC/PP5nYqG
ADNOUpi2jV3CDT/ocCyyzT+fsMkkSL9nKICcIM/Z/qvDJ9yI3pXEsp6Ph9NYE5li
7RivcrL7gr7Kt8qVxbLEUJS5TxZIcSdvSVRNyexcGX3nsfdBUT1R6sT7u/fypoGv
5HVHxtB/u0mtyk8lbM4/biZGcGZQKc9VmJcNIoc/tWQGOnKdMUv0Oz2TgYkaAyAN
3vsuO1aC/d4UeZauX+aUAYOXUH7zPBzi5ygx1pPez04nKKjX2qTebZJSoxy+nKQG
uJ/Ph3fnELkTgHktNlxzXSsQNESt6oYRij4WobbJ5R2PFXIPTY9IcYxcshkySo2U
REvhZ45x+4M11dg02+d3QSI/tLBBhTMQC+Hjn+No24b0xv3G7cxr8jc02Qet+WxH
pj0KLgpz2QsKe7Co9PCOixNdq5Wah3gxUfT2CARtclNtLtqO0Ibs4f9XX6Bm/OS9
Cl1hbzQlOLgf/733RZwdZ7WZThTaTbVZg3/ZrANCTcdidoUeWyAEqrpXZH1JMBoe
B2XrjEHVDiRhJ2OYlIS2wXcJZWGBYSux59vyTGo2pLNmYSBW3T0cmnukSKqxR4gq
SfXreyGBFKgPZNX/lbrRMZsQxblyU3Oc3+W3ZlWKhi173pQQ+ixfhstzCXfL5JN2
DtBMfBa36NDADsANprOgFFwOIeJqU7UJyJtZ2XAEVUVdRPiN53GkVm2Q0/8H5K7f
yK3cTXbyS37YHLjsplHdMjepvH2+rRniApmj5AGXi3R+cIOT4hqxRb80nn+3W2X7
eO+IRpnW4dF2HaUo6BiJg2ao9uoCV4Z+Gml7HDlIPeU/5FLvJPT9K/z4Em/sBuvy
m5C+PM574xVzeyMEuBzitxfm/z4R4ITP6xyAhN1HAwIA6UdNW1b2NBeuIVeUsxA5
0nvxa34jMOanf5iPwr/VqrCuWw6bDHybAtklqyfSh/QXnrC6Uf4V0eaGxwGyABtU
vEN3pbd/MAVvf9K9rJ82AZ6vHmTL7iyWOfuQS5KXies5KNt6ygPb7roaQxtJ0IvJ
7spblBlaqhFDjzswk/DlHEmOwUXiwqwOLTKpLqjBMn3I1xz+VYcxYpDpM5YPQBkh
kl3Yv6cgg3Rs85uAULIVKIfSdo/GF/fjIEkfCWzc7Y2/dWBfDQLtlhFoA9VPBhUQ
POqDqyKuSjHLvkqZKaNAtprkhCLQXLlGDIR5U3xwiqG0UiRF1wK+kMFQmaxABMvU
XSy6522pCO8SpzDh4Sy8qgEEkD0m5GnfFx/JTLth3e35giUyDtbYCiHD8ob+WS5e
wbSGHeRXHOk7ru5qZgqW1PCAx7QqrLF4bnYIeRGLPurETrH0Tk0lj2kBffMgy/JV
uCUlhZqEnJqT553XSSTQld2JFMGcTlzLmLA4DMLCBdYsETe50xrDJMj/7Tybk9r+
BBDbvxLGIDEUBqGRLBzvcvJcmRpaj2qz/W6ia6BaBU/iEDScfXKmW8l4R01+3pJZ
3TMKA/KMKuMc/ur53jrkDnvG9TdVdAx8/aQ5KyiL58v3wgMMlBo2XuRQxRxx+B6Y
sjvQNa2JLfCKl+2WULCPY9V/2J7gW1lAiUTTHKIKYAGqJqJTjOFWRzK7ZXNvKtFp
cZpSEF8WayxFXxh6oj1lBxjFEHC9uLb05Rm/dDq/YOBm+Cm3aamGMBtF+MNg0mKd
cAr051iOeZZ5L1WBzfwVhoBCYv5x0bmzp1HFty3bprMmJwj26TY2ZjOSZN6BXVTP
0VyrWXqT5fIQwB4d2uD8dFCzYZ4tSzj0D7EXV4XiENoZxO3dtTDrsFf914sqqRWf
cZksSA6RClxvYsDfdA/lgLEw+xuk0dlE/KrkHOxGynwHhueiBVtyBjN+OKlqm05n
1DlaS+UiTWuU1VQOevG/0Bcy1RU7imK92v3T5EFKo3LmlnY0wPaJjozV/4IbkY0N
J9S0/ge2sdMKtfRXP/FC/I5NVPBuNraOl8MFowpIQAQ+XkRbFsVC+KWoTlEwg2IA
wVQT/3Gu/XbQTxeMQ8XQST6xUW0taiIfD8yJ/kgbiK079AUTupS+hMjzseBN7x9m
ePgnVsR0AF+ZKCTpOzwYsJUZt40KMfVWntm1xLlm6avzhT2JRw3AeTIWOntHegGd
axg56DPH7WPZc7XR3XVjdN3h9ZxyzohUObWXLC+S07MTF9XrFjJbdl2oIAs5lvVh
ELYr7cL0x+MxtchRc//5upyk7bZEhmX+R6lYs4A/gZAyj1hgB3wlEXooae5MWdHf
Q+p0lkDIMs6vIqq9ygGHYgC5l0ymu4wWhArhuKpC7OhWL9VKmeNd8hpYR4alL4e3
uLzTzpQd9OsnhxtByFfC3W8mENMxNNWiSkqiRs+2b7Wa6yE2vzG/sKk0RrXUPQ2v
a9MjAj4JUcNr1pt8VMNi6tfFe7RFqcnrkiLXgTmoOAjDbNYO62SBgmabBMwWqgMq
IxYl8+z6iXSHhple49xoCDNWWim/XKqPOTUAXNif0JLhUHnLsTP30NKr2z4WP5v6
Dj4BKJerSu1VQAhvaagSv4YuDIsc62P7bMWMZ8S3ZrSJ05bG66BvZ0v4rtuKB3UZ
aNku8PJnsKckOZdojq8mym6WLpfa/HnMjctPy02xePon5uB4RYzXgUPRueEFdtIL
h45OCMpkKEASZILLKPwLGfBVruJEE0uFE3IkTQAZZSJOqYoIofL/hlW0ifbn6nUQ
sblZR5Bo0igCb1preFZL4puOEvnZ/dtYatTFCHL8GN/RwgPj28hal/ZwoWzUIhSu
N4KwDGLub1UO8RJbQuT1P8xPgBTEcHCQ6mYw15DgiY6JA7MwCCp0HOPKVs5S53Wc
u8nOjKQbwgjG9oRhlBO7DHw4cDArXxAg/HKXN89F9GUE3WpFw8VfYqXQhnIWUhg3
CQKsntmqckqlipgDrpqg2VgQ/WnoCkpkbmPY5O717iurDPqmCv8tonyK1OH7nFk8
DxBQ8WgJIwMy5ufpKlU9DlCUF58jXKjFCq3bLxm2i97GWzXD3C7Ej/fUicILeP7l
SaGe4CUF7gXLRKcG1kY9S/Lqy7p6/Cb4CCggFgZ1fO1HK+jsbTKu3eSg1jJiqBVX
s4kBk6lb9P+UusnIuhFidujmAz+OKo3lFCAd7a5dPo4gmbYGRjJqS6a6V8+XTaFk
hRQyJO0ICVGkb7qpKtRQJWr2RF6rKv2qGGEnv+0QXWKCH3CTF3FXIF1o5lCpdYwr
xSwqmiTn1hV4ejxYXVxQdF8mWlZKlpnImyQIX4DAk53FE0jXeDT0iZmbTZ82zFX/
oqGe6S1z+zAnjS2MKQ+8b0vXs/TDPoSFJI6cne1+NmHQzxqYKH95L1MK97i4KMVK
P+ZHPjrxMRzxtne5QjM2yzSpYCafxt4R07z2asFLh0gXbch4gayCzx/tgcUfe8A4
mdwKIYoUGFNA/B92yudbQ3HSUVIq6zXWRzTR8TXoKRVntj3hDk46KuhODHR3b+sv
tP2zwe/qqFaNUnKr2ijcs1nPyaUPBCcYT1vKNBeU+2B+5u2couDeEVO2sadampPS
bG7b8JhtcAtf1cpxUkhOmG2RY6i6pdqrz+a3K/zQ6xYmWrgd11NP3esBsjjLPpQ3
1K/4PVWC/EPzfcEeke1kX4W2iKa6iQq/QLLngrE3o7LDQWdmNamf6M3S5Zng7G5f
uQ0sBJj5D2hz6ADVNsy7G65nWIsqMN48t+RrUkOCAJwbSgi2XCSvurWjZpLprl4G
5l4x2TCJZ8L6Pqin1w4K/7skcRLANGvGaoswhWbKhnZVz2Yrb0oSIUAJOO5cLd/S
u78wZhmoCDe/Rk4JsvYmdhFsDFTRc45bi87IWFoxzAspdwEVLs9VZMihRqSfx2ZQ
dQlWLxeNHE1pk4sSfNinySkVsSLQK7x7DCJoVzkoBemi6q4xsIHzsLJpC7KPiakP
ZAbQ89+8I4pzAMVXBz+BiHJL2IIcqLp8MTqKTF21WjN5wpJ8fDJsbKdubzi2Hj8l
NPFAEJUXE702krh4FyZ/QPkfD8jItwSznN0CPzXdlLjCYiEPUlpFAW5Ybmg6CinS
13wIZZmJJitblIvVSVPjc9n1rat/XRqHf3bo7XgmYZhcOwYkR/ln9xLBY6/t5tAy
p+9RGW5xBFkdyStHk2GkcBKDbcufoziV7N+RcTXj3/d3Gjk/S2g3UUsjHyIMEtOs
s0ZPH2hEUv7V1yYtfrzEmlaY8w3C6HdV2xLf76tTHWcN1O1H8bGTB4OYyaNSe8dj
d+jhtlTa45PtF7rm0MSQr8UAGqRLBu1gWTYi3Trv5vkCWDaxErjmO8IeEiYB7fXc
/Uhkfv6rhV8sVKejFTSGk/rbngIPDkqv3k1iJnq7/vxuatJ//QWq3FtkK6esjqtt
fxENsqGWA2i0YffDv7ERLJAXUtLPlvWSE8QVqz4RQaNlWwliKE3Jnr5ue5EFCAgs
w/F9+ht6++jmuJRbRuDluPToVAaEaIGcvq1sUAhbQvUUEbZQ32RsOrEXwZgVxoWd
r0tYxjFY37GfTCnoS0ZswYHdUdBw3MQSfxtB3H7ncMRbuRefF4j+DXXYyz1dAFG1
KFq8G48HppVKcgo2FG0nEE7ThmxaJNwPtsS9Iz9xfrfeifZvCjI/IxRrWE2QGgg8
seY2+Xe2UHyh/9lyPh+YDNAsWK/5xiNF4KkUj7Kfsq9qZwHP/U1e1tWXX0W+dv28
mcapDYLgx0fQS8Dz/n5eDiK44cQBsc3L+6ddYdx3RS5Hw0xs5OGJc2JeLn/Y7BTV
2h1titmo9osYTkLRuxR/5nAOsid+BQv1Q9ze7SxjJ42SVsA3qv2kCiWlBxB7pwvj
uHGpkBI8NcTHxXwWC0XNV9Ase3gajNQuJL+HCRLT73ElwKu0jhxIIf4tBP2GZKzz
FPBPOZ+Q3Wsg/wSc4saviVewhbtk5QSymSJVrAd83OVR1HFDFKZU/4nc5Ks/mk0x
tz1fpw63nXvyje/yTuIRiFWsz33mTRUsLn8Gtwk6LtesuNBbjOGK+cEj0+Lw2PLB
DSubCmsZaQe7MjY9BOVRXxiLDm+7hrXNL0WQny56g9lIlA54H4eultcmYQ9E2Tbl
PEtwolYcAIl9ZrlwROXgBEP3tSQwpi31SuUKDkDKhHZZTfG9PUMQhlhi88S7P+BU
dfpfKv+nX8JrkQEQElwLv5mbTv2vfG/GuY2TKeu5+nz/sO0JUAIQ3OtJsVx2Y+uq
4b3jmiw8ggiOaqtmOHF2xOzmVaqdD2LaAI9YDXzfjr88JGeWQavjOA9cmUvyb21P
p5S2P8fHjpWLI+7pqdUrXOTNADXNJDlnHzQqQT8s0CYpDqh67MjCvr2vL5naFgZP
FphK4I/pb7eK3EXWOScAU3HKki+f5ywDrH4NA4T01duTBmWqM4EAF3yc5CYbh8Qf
Ha1X6+l3YgOUAE3CrcOJPT5wurbpjlxDgYAiBPge455UReOVD5UKQIvpZxxUzeTL
RNj93te6sZeOm64zR9+hvzmys/+OB+6vpM9V+/Spjpe+yli5Ovxi8uakuRJk8BVa
a0zw97s+dQam/YFTYgTy5NFs7QGpYsR5QyhlWWKZrYYrQdkpWg7KzQQniW66gUMh
wDq2ZT1vtAM65T1uQZctwCr5FSnR3MrHIHEr5EJehPcLhPBw4mMQRJUG0VyqPCgk
JgFo8kNFxyuCaD5EGl8E+Cj00l3j2PNmJO2IQYkiDTQJxGoxfOgi05PUYuYmRre5
f7FTlQ8YwI1XmrtcVFrr9710oesLhHpjhV8HwMCSdO7xeJbbJ+7uE9o3eCJh915w
4CnAb35/jboKmvt1n7nZwtxCPRAIzc7ev+ByWw2YA2X3ovd3z2ELhQFHLFNRY7xD
lke2cq5+VRuHWRgx+X/CUvlJbDQvsH+acOk/za1b7dt34hly/vsLrE7w7FmL4h/Q
gVuxSsBh1jiw03DOdFeNsCzKqtnw6grZwkP5c2fwOZlDS2VsH23OP2sIvh+guIju
Pay9yWeaNl1e3q50uxdKIcuuH+L96UgJZ6qKo4v21OpPWOmJp0+umHB9xVDv3EHM
fezMJhnPazpD0WYriZPDrx5d0EElEQJkAEgNio3d/D5sKjzOTxqD/D5dDhTqz+A8
/asknjy/E7/CheuUuwKGlGQroX4JGV8jcgAc/HCrmzIl5qKk5DcqArgBwQ/Y4Rn9
cEG8SKFw8VxzcjhvZdSpARNQHGLjw683QnxeL7HiPjVMgzkvBy06ZRnb9wYAwfYX
kMCbXkFs0XRoObee2jEaN/TTyxx8E9PqNs61vxlBrLWF1GtZYSE0dmYUhj8b0Q4+
q05mBwEfW/Zw01Nd384L5wyMxtWqqveFzVSr92FTPcx6pCCr84fDDeB/i7YFLRBN
d4kJpvOsuPQ6Geibg9qfoqWFhaIlaLyhfWLqVLt9A6EnRT30poREvQMVvgYVZzpu
4HCPQyc1Nxa4KOa1NlW20/UJDXviU2+0yvBqwS6scsM0T+GnPwPCRrRUvyI2ND71
LLhZyMYe+66kr15tCZt5S5i6ZSpmRAUTNVi5fDTDhuJHiOvjj+P0gPTJJEyXTdxO
qeosGyroxC6AtJttgN1f0fISiORt5LupdYK0BptUfqOkxN5OHtsQPwVVC8tVSym6
+ZIkq3g8uljHAnqWryiaqbH0a/vAeqTZDxaUiBHnGcmDW/fleLl+vU+VUuVn1BVX
+nb+qbRaw8iiZw27LT4GvQmk5RX2MibK6WqURqH8bn2WnwnJrYUvMLRos5I74hec
4aMld+QyEW9zJeon4Kw7Qvligc/RL7kpa6BFJV86/6O83Zi0lIgmz0DyGNL8jaTg
Prg7gw/0ejrmwXCvQWixTA4oC5Oen9EfE20F9EWe/13J7OKA67R0LUk5J/ABvXIA
DYJk7PawfVtbLtuhhEatSMkvUmZv1blXL4mkl0bXXT8+LueDtAyt95owA0+g1PIH
aFuNnl87GeSvWkgD797QCKEUHidJzA39dBH5ocz+oh/fgMTbOa6i+lxNHwb1QEUO
ZHqJ0E4W09in/4n8sanLZdm804XpOoDX7bhgGsEt3aShyb6/078zMyLBr6beTmyE
5tnGlXDHnCZb/HGSlvHgG/PW4VdNP1BaHgJDfExvr74ZZyk+Q5oQfjxgOyk9ZMHj
ZpWsd4S45mRpJJ9L3m4i+MfD1DTVraEYmHOdL3U8Xnvm3wBSS9LKScyEXu/XvUI4
Wm2GRvpQYXHqI9F2rowtGH17y0NWOhmuawTQPH+oPO1sK1e95dxROMgeFTovBlGG
HPsTN5Lj46w2duMIHNOH1zFvHx/1b7lRS54BksZK2hH3osTe4ohdVa/zVX+SJG4k
Qzsp5bQvnZRif5kLAju8oDmxW0tbazE8XSfIW8N5GjNskj5KdEMgynI9I4KlGzi3
1hGcFftIqzGJng3aSBTVP3oa7y6o5KIkNHTVx6Cyc8NVjL1youuqNqT3OVqSBoMk
nWXQn6HsSNgr88YIIaIcJ9d1ZLkyK/QNzHcXzs15bEzEnVDWQTZO7iZ3PTzPPfj1
Plz0+mCm2ZkSJzFJ/ehR5gmE6VJTYLE7PMbakimtX+ev2dgHaxEm5ntjT01Tk5d2
kJuj+IBftyiodjwxjqLaBdC1Kc0axDuXcGQHo6Hr44vPVv+3tbqZ0dTntjRyYuqB
tmryFjxqp7Op1vqTr2/+CQiK3FiTaqjDLj3Esx6mJLvvAFfUuQOuMNxtE2Pg9+yJ
k+kbd09i/5p0LT8mAAK237ZhWVxFoiY6qokQQ4XkF639oQ9g8iY/H2zfVb7/EH09
xkqjpGg5M2LAclj7c7QceHgsifnFDK4w3wIVYyK3jzGuNvSsi69dfM/93B65YJMz
FFIu+28jsFmh8xyHcnQ+0adSE1+lSLEl3/Rny/Li5LQ74LrI+OgfC9+j0EuJytvT
8/zV1t38Nh/dXZs3zYEPHOLpCIHEL4zNLXDBkl2W5rpMkiVqWkwa8l9mKpPvoMaj
6b7yNJHMZPH9y2S+GI5UDCyxaplzd2WJZyz5G8ZEo2iiwQQLp9SjJ2DO9sE0navP
nX7tCgXmr3jZntCnd6aKMmD1uTcfPYeMmO6W0bjHafGUAywgVLZoALP7+x1sKv6Q
kw6XngQpwVsWoDv4RAv4QnMpSlazS6cCxvpd7J/FJ6cbPuuRWohNHxVO5q3Ty8a/
BbZB+uGzaEEff8fb0Z4sJOOslBV2B18wgWrkT4mHUa/buP7i1lLFCCYAl0mfc5EQ
2FNVyqrLYYjIiiGAz3Lo34vQnCzKT8e4rwLUmU+IDIM5qzAIiCr5yRXpH9wTzDQ2
8Uu9Bc1e7TK1XbHt/nO9JBINfzKk2j6a1P9DOgKHwSJGGT5cQXKDNY/3cPLrhaGN
54tWbNJWDLjqATH6ZA1/hRCWVsUNLT7ckeBrip/2+hAkiSpxjMku0CaIoIUn5rxT
w964a/l68wmk35BPCdY7VAp0rPKlJYPFKE1jFfALT8y0LpcBwFH3IBpliI2aoySK
HLu47t4pz0RsIFG9DlUrOOrPnch023HUYqp/vA8m4IbKI+Zz7NkLCHPXEoKFD01Y
stFQNMo/e71RcuzXF3/Cn8vKeqGwMWmP4bmHuLtWz46wnqbu9KEctDS8nz6Cl4c7
YLV3f5cb7Se+fRSauf94RLZ4qMzZ9USQ3aDBpAyj+BgTpXUl0x0es7RQn0XX/whq
VqlemirMd3w52HrVKyiTEserc356Er0d7wajM6Ny7fCnKIVjhbkiWZm24mn6FyeT
PapZozRk2xeHjCHnFqOaWs4LjoMPKAMtopQLr7T8BYGtMaBDfYzQxn1iMQiqmVLp
hV4r2Thf5xTW/TRlCC2ormsalH8j2D0DmNhQTx/oDdPfeeNbi3nEV7mqZBgcu5Xs
8hiehu+y5ADuxrNQacS3EBvEHmfDytIyzbD1tJzUXBKGu2vS2xwug2jt+S2ISJAv
fXEeNbOhJhUpdK8ba+ygDRo48rwiC59V+0IPue+RjUfCUToD47Tith2qt8+/vYk0
NVq2wf4IKdDzyQDGcVXscMFvWvGqsF1ZXw72gA9suKcsICNq4VsIgSPGgKyQX89e
G4ZwGJ1EjlIbBN3jauSZeZIzfB1j+VKiXpnd8gsGL70O73cEpkCHfFdh3x9J6OdM
CweqqZPyCa2FzaKeVnIc2gjWLJZRmd+N11xRaiEH6Ftgv6YV0zDP6916dhTgJnmL
wcvcl5wmo+3DEeGCkbLA/KYwdE2Y8+ur6UwIeLkC8hDmvoaD+YOuNNSJZ+T7tDnR
r6ZeMW3bI2pCO3U/3vb95WzGt1eQxUxa43FypSQzcfZci6YwtK91YTsXrq9e/05C
5QafILUJTXtTK6BeMyE7zq8Niq8Wim0S/P57xm3y+aFl8qXKvQC5z+qV55hLCkmR
JtL+doyHyQZ7FY54z/74aa/LJlcImzUrQpqS4hr+0PM9HWsaJHYV1c8+nApl6Hse
NARfRgfBe47V5W6ZxdJraSPxWpWf43an/3X9/DUKx/g1nDuOZghi+8j8fVKXlv5h
VADsXRSTD4CkanK7mJg1uXw/rAlLcrrP6s2+ziUHz71By7CX31LPwZulAW8ec8/8
cjEDzfeGr1p/g5UFZxgvOGle5gYAQ/7Vv8r0zDMulFhoJI+WxhDw3aNe6LTdkv2I
QhoWa2ybKrjRLCgDkBzA/tnT+gliDt+39UactM2XL9orJI1lOMXoCnu7gRSEHw67
6NXKYzHLlU733PUi1xbjRrt7H1amGHTaDTV0MmP2dS5gbPpCbDxsG2GDUBWjC27f
Cjde7ZzCj0fa7wHP/YWu8CUjvscswOeI7uQK/0MzfLWqYsIXKEsCTSe/2DMQKNmF
ocsu3cWcxfJ09f39+5mHM+Z/Oz3C9fVE7iBns4IprvVdBR+LT3uafb5X+FUVi8IY
JersHv9EcNL8PODA1ggb57UBg/BuQa+9CdC5dK4VaBpBR8EVJB/KU5sreqB84f7C
CM8HXzxu2RRPigtdrY4AZloPJq0+CyAfB97VtlVKv9CCxbKDJqNJgTBIQJW9U1P4
zwSmWOYQ3Jo5rhWKch2k4ebX01Kv5nDYhl3wLr8oPhHdX7/qEPs9NNxHQ/LTA2hu
sBV+/tyWtb1lIfGCAO8X4z15bR8i2mbpDiT0ItNlHFFzFOteVipp7MwxwnRbLWG1
gSQ2zCx0Th9ukG1UFw8DF2JBX16Qyh9otftfg2dIN90dbtg0Xio9CfYzIDLqwVty
x1U4bw3y/+NwiZVxFHXKY7LEzw3ga0nJa876cU3iK3ydiBKXwUvxOoGHcEvPkeqc
Zf/1k37eM1io5k+tnR4Ck//DlkGn0CfG41EmltMZcAoKe0caCZKPmzWWEEWoE5As
wQIHcKMT91LT+RSf0b0XLUiAE7T7OjjGGHEf89/ysCe767L1VL7GwfisFIko1vaI
GY2O07+KZEsa1dhYZsi1tIQskRTUGpmFoXMfBgglXRstw/uun1ULYIYzeOr0rYEm
a55aKgMAH2oRgeYS+r8HmOrZl74kd4pnVoAgSA+zjUoQelJllHr1RlCckm20jygZ
g/XWohkjcFoCt7tfkuow2Eb8qBj4myGRqwT8aX6Y0Izeu1U7tap11tn4+BsGRWCC
nNMjO0ealc3iJSlnXlWMD+OzxBqc/s/Qfcx/o/ZvDPQOH/UWJTnmpeDl44PcpZl9
UFVsCW+lKChU+qKy6ba1KaURwonoG/Uv4JCbDLr5f6nALh2mq9fWDE4TGJ4bkuPL
TLwgpg7on5CzGE6qUAaX7mRhGuIBAJ/GNyo/RIsZa1QpSC3I6O8oZheQuCDzxuk7
7Sr3OUdYksLnv6es9oxETd2uRt059rIs7yHX2VOb/VvcMnlLjzKkD5SgV9EIASXI
2mPfOtx2uN8rSLlmttGkzng7x02//++V38RoD29uXgt3+3gfBuSbBsD5iOTEwi8j
gnKJIF/SwGQyzzKpVuBFXqrQ0d31YSAztZkIYx6xWyvkk8tj5t8HZ/5y+CIRaYMM
FaNu4dJ7jASQF9vfs3rW6L4CF5BBSjeCA3uacwfLlasuV6SsUX7kXsvl9d47Z9LS
MiPdW1dASdh7RuRQ92bgdTnqn58xxtM1PXjUWfsc76ILrzmEfGBCbOv5/3+GfyCY
TXU0ldCOlTAgB26uzXddvM0joOttUxRhFfr+1ta9D8pDXQYc9pJSkdwW+JY55QXc
lre1zzBvI2JL9g21UtvycpL6fdX3/8sCrsLZT3kZatrSF9wQJv7hzrxdGNSpGAB4
VGMH1SBgPnTQpupSpGp9RdUGcJpthZftwquIZxCpGjJuciRWOvcPvifE1uV8TefE
F+Rg563LgVDWQ38D4679AnIBpnsVxxTbmuTK5ON/ixYoZ9Qhwp1PrCIpQ4CtnlVH
NTtTIZAAiKH/MltXERfug9FMbLUs7IDxDPYtEZ5LO9udUs7o3vAun6X48b9XBADV
DOgTqDZzQGskxA8z61CVuMOHYM6e6nAMfliXp4PVkSLDj+Qzy305T7ewJjZ6r5lj
ImPLtSeY2VvipMWxyWoePM1LvAXiE8GdqtnrwdwNYJZcRAXACFqXj6eQ2X0KAevm
+aE6zPtOhQSkn6mjaqsylACaSrZweJZIgT12MvVQRGMvaYpGMc60mbvkJlM786SC
66sR7Xzuj0rmZI5mE7OXMYM1DR/hyhRULePFxy1n20itpXE9jGg69x/b1sFOQwQ2
yOLU7ndREsaoMZx//goFJMIfhJppeuTBSrKMB12ZmEBheXSPBOWHJJ+Jfks1nxhC
1f+fo25vcFr28L+O4UWP9S9iOiJ06GRZybQBRC+WWuAcqFHCY1vXOpNCl7lgwAf6
QKO06ei2sEmfkdY6monzaw4lvpEQZn2diYdSxJ7UAY9GbpJj7Rxzufu27jJb9rku
0e5wf+VAML4uAbdEHSavfikkXWGMzYUIS0oFpDPvoyeeimjVbRrezA0xjSTZNJOF
j3XpO79vJM1j0WlpN7zaiYku1M52FjPdVO7xrLKlmzhckljeNScdfotD/Tmd4i++
H92QU/pyOLmoSsb0tTU7Gv+RS6R1NKVSBmQsQT4eN3YWml+3I6E07W+DOBQmJKPa
nmnq/kUT+/mm6RHHMRuHESucU4hbDPHP3u9KK1itcjrus6ajUQwC0OQ2Z0oqc+8v
n91CSFeghjRe3BryDn+Nq+ZTAJM+j49IxLP4I+u7+uPpmXhXjTDSgAtDrF/zy8h5
dJ29mgng3KCSAWncT4hqmYRyVWgM67sPYBA46WeZ+1oOaZDaUyljXuhHIf/li+7f
nhkGrzKi8woxoNM9frO4ErJl6YxwZVARNtXHmxQiEAIzHM6WkhA3IFDPgeQHuSoc
k0UZ+j00bEKyANwQ3FPeAYK1lINRKpoJzddTgwxow1H/+rM1+kfb2UHqzUkwEA31
aFb8O7E7pO1yFqNpheMLSUaOK/Cjg17A08yyI3HRbgRtEZgHEf7y9W6aB019WZ5O
wtc/ozuo+mgGo2d57KvRoaKkAyjpvl1erUw51zWeOTqV2tJZ2iaeGAsBWjP9w3P1
eJVvqO35kV0jxH1TLkG6kKmLmzXncZGUamIibG9h6VMgcRMxXTIeiLD+oLA1JL4P
wY01FRohFEgiUaIpIA/dJtgRwtBsxRrVP4NSI71JhuduY0JvOI9yyN3ZmVev3HdM
Gn6aKwzbHbhnKtKuMkk9MazGdSmPc/DF1Kd8byY3nA3ti4Fzix64lo8Zjg6wItS+
rvv7K+Ag09zOtK2qJcNgr5rl4HcWiFyAJwdBz9wmGeBVrUErSIwMSZgUUN2FRYx+
uL8L7ncUqQqoWhm13Sgr54kb8Pdv/zJ6y2gzGc7+JZsOjX7fqxTErAW30/JQ4acZ
YPkw052fYLJGFgN2t0LTWI4IO1gxZZJfRBD/e8MI+iUhOlbtiPutDgWOrVF2vVxK
xoevF8R9npV+jmoyfnTAGV7CNDLPmfurff0DHQNor2ZAG36g0G3TxIDmjFDupcB9
RFrcY7eQnTJRyW0G+OIAF9Fdu1TlIpwR1tX6WIbcN082Lt57uVhaW/A3MDMpEBl0
sSIwi3IcFxaOHZL349frm1o+cqwaeL0WCw5Z9rJkw3l3eBV8RPK5nGFF4j4YIaUD
rOI8wkqC63PzpjX8QR/gS4lvt9WEZEl6MScubZLCEzb/jKomcih30Qn2RpkrQEYO
mb1yKkqh6/8t0GESLsUaIWm2lE92HQoDoYx7Ngvz8jPzfk3CZANWXaWMoMBKpD7i
cZXqstu0eq+1yvMpTm6gRVrmjrEm2C4iFyuSd01+85AJGBl/W6pzrKQYImORBIJX
9Z395GuYLX2YEhjc8/Wdtjws4/vwjO7AMFU8DOBNpLZWSL4O0kP8ENGAhNrAzESz
Pqrwb7TAexMXnRduAd42kR688x28/bPM6cpW2YpBH4p3FIDc+J+b6V3JbEToLCGj
u3X619HZlCNLhyCPO1tfK+2Mc7QDcBaezgtEOr55lUdfH5JjVMxWU1aYpz2agcDU
VH7HjYQI9TDtl1X46XJ1B5EYHGUZVYIkt0vefemTLaqsywc98O8wqWsmlpbJRBHq
sfycMOh5UqR3DEIiy/G0TpusneuPx/88Wpypr+B+H6SHZxPHalmxQi7RDEc9ys9P
ZPJ7uUKm/gxtBsj5/nLMGqMQYC/ADWZpSr9xjPaf4o9OQmcOpQ2r+0pai/5VSM6m
pkMoCyCSktBNWQG90alNRVetCXd+ivKvu29mfj1ohr6fUuGmaS/sU6a511Ef3Nzv
J/AO7TCz5iv0ZbpRnt/5fxcSG2FI6MY/CVzknBUe2NWHf055dnDlEq0A+m8EFhW8
/coL5TT6y0Uhv3k4Jzwl3glfGZOzpWxvi451PCbcKOSeLqtYZWFSMC+z3khNySp2
CNAeWIaMGvjnZ7FQkEwGL59YIBA3qHHZhZRwya8OjUaLDniJrTZbl9EfWoKN5P9L
/vQRJhKW24EMuCWEfqmU47rzkJln+7TCeJ8jEeGo2mbkqHUAwwaPcYSHjmlIYbAy
cJZZvNeCxtQw7+NO8FBU/7pa/eIcUhFA2Hx8qQIVJaENMb7r/SMYgCya+q/3znwv
feYz3JnbGY8eXDJg9RqWjb5qTwMNdaW9831Di8B203Kc9RLra0YTVXa0iLsYfW27
mwy4ZSl4Y5sb50lRZkP05zoj1cWKEGJYPhEezqh6MvmtOB7gw/wIq1r3IhKs3vZz
4xlf6PLfjAsisdLCAtTvIg/9DKRmrKfMOrWANQg0r/Dw10aeq31hY7M7MyigqvZK
2kCiN+Z/77dx69ZEzTHR30JfkZZtL0/euic/T7R8ESTrGb7lF3fMbGnPvmya+NC3
c1/XsOulFtidZcbV6INaz+UOWvNCcKRxA6mRQjZZnK+YToAOysMkMkLj4ZEuf6BB
QQdgVLZEQ25/plUYdROqtzNbuzd+X5eR10iPQmcWEeDoiuLqt5Xb1fakd9TldI4F
jdRJBGqKchZkJmih/NjUrWuTjdEUWCkohuubCeFlPtDjg6+4xyBgJjTChp8O953R
EAOtFlwaJT6qZqp6356b40Bhjf6pgkuwnMFd49PdHB/QjZmTySy8qr2L5KMoCE4S
B35taN1l1Fo3PI6Ef07LNQtWbbcnN3Jj6tEd7Y6nqluzQi05XVUY7R/a9ksTZD+7
VtgEhs8U1hjeQS///jFeAa9thnD02s4KYMYfGxWsWcSyLBdFZvHt/fXTEOyFSpBu
SoW7N79DeDtTn9G1UELdzn/1GkhVUutNgU4Hp637/YXUUIUcVU6vjLX6s2RRkmm0
JPdv0vqeWCFX7LXhLv0h9cPzj8v/NxsnuwX/hSy4bNaz/eXZzhD7hZFvtkxSv5Lg
BG7m+NVCjCPTzjat85aQ33OIFCWOfibj7uzK2XGtK8DQQZa6J+SrVCOWCElusTnz
/RsrBzKmNxJKKKPYDp17Le+8WrE6StV/fXzDB/9fG1B8fu5Hdsc3qDlj80XYhwZX
MJjAbCIGHnWljUva9ctokLb/kVSdBtxF3V7cbEJdNGthJTrO2OKbI/gSLBHIza9Z
eNQqK/ZkcI+SoPB1bRSpeI2URFnp+vKpzrNvrbEH0yQoPEMNquOIrUmgZ9HtyqeE
WZ17gNksqKT+bjn+ppEpnMm8LBxsETS5+RS6g24yTOOb6MsdxT9kHSOiw9cBaRGI
T7lOfOVPGdMGILNE8l+rqIreYm8t7Mhtg6Gpyj7v4469rKma/bOSpEc/R9sUy0oh
AHyJ2ieFR1kUCwo5mwC1k6fgPC/qz5tHd4uR/QsHz/w+0cM/LOzDDaLvGfQ9xYOW
7RZrXi2Et+fJOn9dquaxAdatnLjmGWk3dvMreGqJu6imEnyKn7Svz3V1+/X5X1e6
+XzOZbRcrI8eMupjYJuKs5xettqFJiYsNjodpc4j8zSGnIlt5jhfA4HKv/HyRLl5
2ajN2K+A14deOdIO/665Dtn6LMADjQJxx9EJ+DwnRNA4O2ExUbCf6OZuI2sA/frI
C9dVxvGvrEkFdSGf1oPBlqk3blTF9IDwWWz9aRMz+lvQAQ+z/smvenlm5k/A/BF+
Fa/laooUH1vQcH/P9PLnKAG5V3+9/WguHgsUQEpTtjCMYM0ElZicRJFB0NdN+gXA
AsD/9Lvg5XUEB3k6r0eLtYrJTLX5obZufh+jlOAMso3I+Rfl7KzG7eyiJWM4Epl5
eTsZQ0xRcry3i3LjEZRJnM0lcNQXUE6ybA2nB2iT1ew2QgQB8s3wxa+LVFIyLgDP
aCs6MSLU9kNaMRytfNWD7Nn9IBctqPix6IKwu8fYivWs//0VtYUDVZS5q0vs1MVE
JoeVV2OzZg/Gb/ZC1ZPm6Ps3ZfbRvS7wrtLeXk4iVJZ3uMKQX7fhU+IAmUNsSqUS
wsiGVsEE1IuDkq8J4/p4vNMgwsgD0hpGpDN5UCh47OnR0ou0PJ1A0QAOav76onPv
yyiHh3oVkwt8Jj0nj0mFg/um/ravFw2OYSSJO3XwZxQno00qum+vMDZ7536scu+1
+MOIIrRE+HYDs0z1Ef57Vw7NQZSgZtwkBOz61ma2kN/KXB0gLCqNYrwdFW6eDwCW
rKnNkjB/BZAuhoB3YLcxpLBaDJsB2N+j6nuR3l138d5IioCRxooLdeAo+qR99g/i
bgRMHoa17S2g1UGCCrD4ZfAQ1RQBVAyrr2ehRogQxQ1a/3WUDpXnF5sC0kkSgjkI
FzP5WqpjN4VVyWQa40hddX4N21lkBwLDJMfMzEzqUTrUHHI2hU/uEfmNLYfScFfG
SCw/kWigjKz6yqX/pcEP+wPqj19ZVj0z5xOI7sv86CIqBz8lF9ec/cCSPPl3Sc3b
BecQV5bXbDSlwk6cOmfotgDTmKw2uvJVPBSgrmfRyXg46c8oYVsnlCHAkc2TNvhX
tL3gAEaTQmckMPCGpgO7eYjE/uvT8+J8Ffv3WGZj18auppM/9nR0CyKsOZSEY2lt
QPUOXJ/R0IqLEzWCmjC/33G6k9yOn1v4isP3NOLNVunXy2Jr1dK+EOLJkzUcJ5YE
o4lDu7m/Cv6KiqYx8QTCfrfM/CrEEBF6FTaWNRn9ouoUcSqTiM6mXjM96jEzUuHT
8yK27s3OQZwKnJ/taMDE5rsHt1BSFglmx1FcSndDEtX46dfcwFxQxlldDLPRLzbV
QrfdvccgZyChwrzgk+71Zzd14t7fXuTsFZbHZ1rpxiVyVbk+SIgZgEIoAMw/NUlr
+BKWymmJQBoy/GI3+mjXCJAck3CbBydH1OGt99rFiOPObEeav2ZzA7Ha7ohGrYRv
IzSmuv6AmMPR6SWJUz9YgrLbrzjqyrfZJMgcGQ61uL9ErcRDepSwlr66rOmtoW4K
zV4LjzNLFBRtMqugmthKb1bTsvHwsnHVStVpEcwnTdCy5VRkP0px5EJmzvzjihf3
b1W515O5lEOhaI/P8VDB80SEwpIVrSkteRnfugh3iLTWXN+fh7FY5R14HIY6oM9w
WwXDYhVaCnqhAdFHR4iHKxRst16+RU1mIRaEpPcLBWeGUtYFI37elzhiFfZtqVan
yKThvrHSpGNLVMTx8bKPjeGADGy98TF5WbdnSzlSPGlANMvVetaOVs8rKb4T6OS4
1kvXwoqiICqam2RnB4KcqkMJe6pnKAYKOcxv/Ks0Og0xLiH5rEeYkPNmNPtXamwR
krnjNDT9bQyeW68bfoIxotzdkXmFt9fzhy0EMnkEUgN1I8QQqq6SaC8SwEVdvf0c
bud+nkgnvoAmBjFrqDmvayQSoWzOlfBblEK7qtgepHmxOefwdR4VHYBX9daJ7U50
iJaP7DROTAPCyxPvqM6IMLXxokuHvmFQqL1FTe/BHKn4KpfA7HZFoqBy4bdtaPxn
nI3PGKKl0WwnCIFNtJUjtUrcWccNsXpRIUDYF/WfS4H9890cFtu62NQvg/I8oBEA
X3EkCEG3rkF2t3WSnG/DEFP13bZ9kdf6u8XYFTnlssZzIxAD5N49rQ+GHUuAwdFj
C/RQgRI6+txuPNNVt2Wlsj/NuC3MkO5HEjLUWw5diAdCkINPN6abIhH80cz0L2bM
dfuG/B7m+efpDcNp7nPgCKBdq4TAlfD1fi7c01sC7d4pOkbF5Rkmse77Dm0BUQYl
RtKdU72UtCg7PypPR/1rhMDe6/x0scAOmv6PSv/ej/6bpiKMbXhyVO1y4QZSYrRh
3YJaf76Vh2BU1G8/TDI6O+ZFDO0NRRwAbHtnhyIDaRXLIKjmYITJV2WHJgHwjZ87
0lkcAAyje+ThshDOU8A6E5s0OPNpeQNgu5MIfPJHRALRo/H+9N6mDk/kJdG3nDEd
eCZLmTF6OaKbLybHK7Y6ch/l+Rqrqq6W/p23Ef974BRyuGdhxRV0Yabxf7ZH3BjT
flMmJirPUcrT+eHgOcwk7n1x8laXvFQpvq1wQELwm45VqI04ONch3LQEnieSe/kP
+pzr9ZMveHQnB6TS2DaeStGq9kT8kIw1byk/AgV+Wg/JsCArQFpHJrG25pW80wNx
hmXVLMX83zuGM4/dG4Myp3pPeViR/hXJz4e5GbFM50q48bHWhMR7yrRgbBGJBL5+
ivEA8I7TOmkpLdU84qXL9NqetjeriPt7IfLrdL1Kzkc63ufsir68195+Ah+xYCM1
JdLM111DhWvaplZk5u6MwSmkVHbepBbgVozD4KYxT0XzscG4Ii8uvyH734WYwJGn
N6T+FHpLoIEwpzipodQeURmGCg25YU0cVuXxYnZwFX8QwXvX8cC/CoKCbI2dI0Yw
c33aw7K0gaIEkJlTJlDlDSNw3gnijwCIhPyZehEs2lYLP5Z7wJBeYP8WHlLHSz4R
VDOgjRH0DiXeW4ulQXr//h6m44oIiIfk5MYXp96w+yiFmpcIHJrrmwUCR9Rk6rRJ
/hlXLdILbtsV6o6pSFxCAny/L9zs5edfEW4Nv88onxD/V2x2gXkWenOBpl3KP+Pg
BpFIdniFDWuf3I/Sv4Kp1+CGz7au732ueD8o5ekVKWZx9MohCW1vyZyZTubG2yAF
xILxWY+EuytkAp/BdeII6JZLbHLIfnWxI3MhgnrFrOnxvmFyoQkeIThh45f4arLH
KKxgQmcKTDAgzbDk9bxyrn+gHiU2UJd0N0xraBos2XpeRfuLLudDqWfon9kXipg1
yCc3E0vaRrZIbLsvcEtI4FALyf8AyA0pDNgaFoXQ6QbcjlshWieCcmmEiOhkx3je
I4WTzUXUAiqxBi6NzIDX9PGJ/pTI6Q3FCyfvzZsiyika0g+vK+YMv4BQwgDqNqaa
/Xs+It9sibSXjjTEGSC0kPIcI366TX9sZzJRcPQqc6S7xcGA8wbTSSMLOsySzyg9
Op99n3nAIQ6UonBZgQcjCz/URIc6HX1PwjZmYD354qhfBXlPMPHh9urzjO7HR26W
D9KYzGJOD3LCy8ShNQgNHdNkvvZfSeQhdw3BMgkSGjeMRKND9ipIksOiRe3+WAAE
DYK+VAWSTdFuykJTrLu1nOYFgbTv8nt++XUfhDaQsgARPtG5qZayxAu86XJlAnpv
Q3eNBpQphH+BYNiPilWqweS7Syab9fnmw3dw5gE2Lzs4oEn+TKGguHYfuQn0W7zf
omDtc0gBVq9AP5Eb6IfqzfSxazf9JYrKDfGZNsfKolBauty6hJUVM3BppXUXrq1U
mEqJy01kF6WP3tgJDZvnOwgcuCynApxTKBtjyKLF5E0KJaBm9cVtDqtIrWSkS8iA
ewYKRGC9MAa0sTnz0dY8AdFVUoDuB195+unXLToWh432mrmdQ2x/ems8QG+yexwA
QCiakryuYiFUchh45xHi63yFjdHZmdiXHRaQYsed/bMZPl3uewjjUZsJnjRJ/peS
Cb4MZHmbX3uTszmLwAeXz8kNRyrGXOaewcYEyNz7nx0WqJ1nI66ZZDvS+m99g06K
IcNmVynFMHpCPNBjAyoiyYlooymIOv1kqXY3BM7YzgHfPhxEcVlPDW0NTYWmoLzo
2//EuYAEp4Sfu8Wpj+HVV7EIOe9rUDPLSVO6DgwpTnLKG9aThNy2bpAhQYCOBPTN
NVbDVWUyTajovj9E4f+MGCQAly6uf2r1fBjK6i+d/hkkoyVYPrXM9xnXOw0sqXtu
wYzv10nepSQ9FZBfT6LdUwP+Jm0T4IaJDipKC1m7VllvOuuRBJ6f4Z3F0RO80cjg
k0ARZxw5cvdl1RreIuFxlwvr+Iz5pIosRmzD7ruprGM3L3DNhEeV5oNrvD8wEL3r
MJ7oD8cw0ZXx2KR+ykSo7GvqfckhRVFCIzJOMko5kdehfXyRcTVJhlogXdRH/Jux
RvWiGmhC6BjzBezFId/oNPsHPhugI06JQXp261u61pZ4ilkAiQhNhBD1UswCCCNu
uM6E6qRcm5eyOvPVY5KSiPYH4jxt3/RdhZ7hSfzp8jWNXTT56x8hw1AXePi25B+0
rOZy7Y684rZ+itsYH6MArtalfvPrU51SiBkKR90hqPHkxPFim9eKwFq1v7MW2egB
ZV0v8J3FXAvF1ynyRPCQ8kMEgVrDLuEzNKcz5KjOfzh7PgPoi4SJVusayp1Y+3WI
WGgLw5Hz9NMAJUugIfCAkIWtuuL9wuKf7R0lA5lsEvt3bwLL+EUXPn/Z9tKazRrs
6rj1FTz3/m4pAt9UM2KZTi9AGP5z5b7EjqgccrjwPTsJAZ3/mqXBmQZfiPfpQUsU
vHRl4/ogm9A5Q5RCD1jCd+Y5xeOe938uD6f+yzGdFvgpf6UYj3fKpshn1CNcq4zM
rFwzN3B6tf+9PnQAGU/CT7+CCb5Qae9U84Cf7j9vTQeDnq8uSEMUqr/mKQ8e+xJK
1EE3dVJ0mF99SOIWLUY2clgtH5uDmvZaE8FL35ChZCTaZuLXQeJtcpGRdhyMEsFh
9IleZrFtDapPrlYcFkEANMkPoaNnxh8nAvyw2F5lojei+nOdr5UAt+xIDU0J7d/i
ud+Rv4oc8NzF08wxjHdUmVM/HjUmxtBy4LlktXqdSKryYFwmmmcYhqT84G3ZGWMh
ROHplHkfUT4vpkxuFsB220zjUay8rFtDsa2/uNjNLYy6X+ZZIVwUMs44iQO8+pkP
7Rkf7edoTCYqV0NeYK2mYyG00gcIdBNGTB93a5EKFBqUdMpAasfcyXXhuyKZkVYn
3h7V8hFcF64UuT35bNabQofKnaUrCs9W1iTHMWXDLfbBRBnhLtLBuyVzdpstnZLa
XuVN0XHanXya3oPJupLZVr8VMiHBLsw4iGLeSC+Nr8RYlzU8hqJR/0O7AXs4g8go
lc2fnJZO2MLkMfI7VJUzgXThuPgQGYMV9bUizphcVyb1pUSkk19e8H/miC3gM9Mu
urudjf1B54xlJAYQ/b4FJMU3+wkdagWQBa3ECQ7VPi2ykBp7CQWeNLXK0knzmbgr
XGEp7ghoHo2DgoOQjeUrq4EbUOJxdwd5hdCJHy31zYtfsgTO4bvKdrK+S5h8+K5p
sWSLSgTn1WwtfEFHbXesOvGmdp7j8qfsYfymbRcOi74czpuz+SYFf5gxC3cNMHjJ
FU8DRLbLLtCKt///SN7jHhafpgqMigcLMOL3v3fU1wcCDZdqwIHaI0JERMDlwlYi
pg1JTThnPvxN7GKZ75hsoQK7Xglagv4wiNJsalJxyg+jmvojsTIRBWyFC5FljdlK
LBQ1z6d8ee30qcqkkj3GI+I1dMUkq3LDXw1ChGDn/QOtaBVkAxzV09QZVYE2ojV7
Hjqh6dJUI6pgm3qdMNaK0fp0o/U/uM7WXVvktcX/MnbavhqxMcfA5V2gr0vMOG0F
bD0uw/2Tyw8V2QfPQgg2t25KhBBwMMllrVGCBSXWp6RIbc5nnX7JRdpIghqVTKxk
DuLcCCBps1hJ31bYQ6NWmp82p7jXzLQbJ8Z+7KTIc2QizVD39vuhCt7lv7zPv6OR
CnIgEIX1w0WTeSX5mdlBmXaRjc1vXSFz97Agj+w2rrZpegCN6rMRsgqY6gECkJTl
zGzNEDP9svi5yLDsvVYCAso8vFlPT0lNUp4gBn/Gy3+MkPCuemuNEim0yzXjnj9G
LHyvPY146SAWvDOuyLyAop4/g7OHzcy19aK5wLnxGzAlsKy83bohEqFDN0bk5WSE
5LE02PpeqjRuOR8NT3OcZ5C+IdlPSJZv3S7aOjhwc0F0Goh7KlJpCWySOA2ssyc5
wKE7lqDkQn0cAtWxd47d+oB2I4STbstM2AtOYDbD6LV+/g6RSUXWz/GG+TmcFlaP
vPt5jsq/g3hakEILUI0+A9kiHJZ52SvgyOLZBkm56BJ8opYyXqer55R/18P8ueJb
FgX6yGHtUd4jOHUlDUtYUs65/JQFmXGQOKPXmxdz/EL8s9IggoUmpUI2TyqpftEp
o62XNNsGclBNF3Kg2MdksInXiE++06xyveXQ/+vEtJrtInmLeI+yH8R4sYf8Dht5
oEfe/UAHFbh8bphx+2Eh5fOIGY9DSNCivRxMqxHryuM7xr6nmZf1AhYlcSbcmey2
d+PE8WcKmptKkt6VLghPN3r9P/ZygwzLBeBOxydBOTqHIMkDDD9ZsLqDpGSQ/IKC
FE9fbpg6rpTBuTAc7gePmeDPEZeZP4RyIxytxPcNEpKa3gNrfq6YCZzD55jrOmZv
PAfOA658Yd5WXhKaL3c1qvNyE0akdk1W7M4Ae0nfrrXKJVn8bn7N2RoWlH6xnfaO
wyVt3wq8cBcvJNHw0GQCRNEuemxkEk5gh/gPbPMyVRcBpeK45ufJv/GJ9HL122Zi
gWRc5pqk3SYktYMtOsb4ZtBoR7o84mz/cYKgzJyjk73OD+mRXMYUJ0YqAPs5T17v
bCBwEc8mjj+GdXtezVTdZMwW4WqqYulCJccbEm8Hb3+yBtbPcgqpmNp/UZ6tsoQA
akWTpSTstjPKozOQEPiEFoJxQv9I3u/rlmnPbReQFu7cxX4f6i2RIyGeliXieZAm
Fpp1niXqcSX0Unf7GDHDadjNJ3+hkgpj6kerEMKAR/93N0F+8tS4DiayN3leJdt9
9ACbzVqOLBXUayPcoCOUG+3RqYxGF5WL8ZOxCkZbEwoLaq/BTPtNxTi5WNiT7cX7
nqp1Uia6PESbDjJh5yfzRIMd8fBZI7y45rCLmiYWcXwisvWGBbav8jxmMw9C0ola
u6Zhxfb5gHa8Hm+wW/+RGp0jiqDr2ETq1O9Km+46J+vewft9AysspQiCP7GeoYcP
VWXniRWctrgxDb2rV2a5SRQ+76vGJDpHvBwdNAldYIUC7bHtV2vaNalU/GkvlLHn
I8bIZW1aaDjJmy/yXQBkok8Rk5S1f6REcVOSV+t5IAJg1a7Xnn2kiCy5Q6mKv+zc
pmzN1+hVGrqAB09TIQ8DNtiiL5vLhXRT3zA/vZM1EIPB+2z0oVZe+7Tv0m25dB8t
g9UpHZtBaiwedaRQ9UcAJmyGcqXWFDgPhE0CYngjU98HgrKBSI/5jiQyKVYUaYhh
u8haA7h0DiHMDB68NI/YqBubClvAn3/Xr0VLit8HdhbcoMENKZSXSDe0LCvaQy/b
Ll6G+11G7rnxJssxPGvoMWE1fcbx+0SnKyBX/A29/2ppw7FgheZuj7lOR3RzAsA4
N/efv109LYq9R5DyfFLzgFDPvRec7s9FkVRgocwRYczJO87qi9GBK/fHQ2O5te73
TzKS5vJcw5BAIrQt0rKIJBUXnEg6amkPbgj+Ldcj7UqiRpr0ecUymIsEuawQKiIH
HBwfnk88I65qZZxD9CU/0XaYdbEiOxv76AUjWVcwakNfXDEoD3P/btJclzL8m7yC
NWn0an9Xp3JlT0Lv3rcxYD20YS4ur9FLgz0epsXoSrr90MVsYthWQF408BOgVYzs
x83glenMlrTQ3wk8ZU6QCWp9uiNBpiHftsD3wC+sbL55VeOoj7p6J1JiT94Fj4yg
dSFTmXKTayfmcvR/lVZhU2lrXRubXKzL1j0nI/qlcqnGihm7cBBGWO4fCE5/h7TO
xJRfXj7jeDYnzXQNk/Khz/V+P5QPWHytrHN6Kc8peZIrazEO7+1hN52TMphDZJBt
fBPYTx3qjErt2cIEqsqjq7CM2noP6qUqLtv7Kp3c1uDYGhiKsnEnAxbJdenMKnmh
66Eg4YNwRkIougvWW4u1nh1j2qaSG52KXcOCePYxW2eYxPeHEzh1OfO2Yrhze5Gk
+oKkTCd2e10z45VuUhFnGPLFwnaHEgYVQ0BIVmBnzxDc5jLsISYTlyzmJ3guILpg
NW6nKnxIYupyZpLb5XVC9MvfT+dLU8DDDIG8qeR5138LRGOlUZoV1EnjA4IxWSjh
c9GsWxhFw20x7Plr4jaVESJCoMccb9dulGpU9tlODpGLGK1k8NWEPSGbFAHulqh7
5nKkBm+HxDvPRUAkkGAwl4NilBGrxM4V/uwNSY+oPHBwslU9qCQ8s+lixcV/5EE4
GdHU2E16W0q+uK1+zozhFxoIRkPr+jD4HjFTCSUJCH/0ChkPdgYQI2A0tQHltkkL
mnYMzBGMhdRRAmUc+CIqpbsy6rQApPkPFknGLddXqq6owNuy9EXtXxfWAvPvkPjK
AU5Cb0F0l1GObsTrSMk2vNiGeLprCZF/GRAYhQd7wERsThwq13xMravaRyqCnfWT
DAYCXIAF6f8ZiFwLQbeQBMAPAb1c1f5diI1hd9aAHi1jdSK7fC4mpObcz63N+ysn
FEqDCGAXMIU0MWTNapDb9blKcv+jJHmNLbh5K1J1grQLtsSVaQQT8UO6phdF+oY0
G/mtgzv0kD430C9QJas2ll59G7FvHAXSPIqfKpn5psuyGdqwZPTfd/gkxbubfc2J
ZrQm75qFLEDKcLt1dgjSDbKpQVZonVAQryRC30q9BFeUXUyNm4Xtf6ou04/0ig2u
o9hSTmgCHvczZDN9NUSPTJOIRz+k37WY4Nb+O7iPgSc+m4E0sbYu+d1fVNep3Jg6
HPVG5oeYuLtolNPE1qVl80SEhGotR6X9WT3xdHmoMqx16M0SOOJYSeqsVROTnfGh
1XLzcFnLKoUUaac5vfbCvnQ5P2mODVSCGS1GQl1S+Iq6DSOLS8qE/L7ynraEciHs
UO21lp0OX2HROdDriHYBbEKFfkLw7B6PF5OxlFgp6mtil7sA4XIaPZcT356S/YqR
NWTfBMaAfr33bGLuBc+PNJ5WXRREorRa7yq6rUBdXCJpldPGi698dLjGsyaQTBAm
g0r1ElQeS22COmDFDwbzetg4gcynK7Ui8KfoOGljZ3KUZoR8UAzUox7q/zQZhzAo
UfOgMJJZJ5rOQpRazhylkzZB52CoLxm2Of0NFkqw1EFY6ay2AD8bchLSx89Cyk5d
FbvzZVKBZ0A5yEk+1BFIJqVqqTmRiIBhWcEMom3l6ZgoU6F7QHhH82hWPaSvj0Ez
cLztwzpSgbSQa0S3rmHDP5VAYZpVguarAP6BtURC9tFSRZyJJz5fEr+6VEPmdQzh
AjXPMowarXM/6PFHLZq/Le9q5BB8HlW9kcBxTdF/iKJ2cmOQVXvKzGpTy6nB/cjL
yqXMozE3iJFVIHrPlTUrkrAsGBjsG+mTyi4/W1NLxT5YSjvdJnpAUVWoAOs+Q2Hx
UDrcQPOim2bXQGxVDS1FE0A6lhFXpjeMfkstyuQHZY0/kdQUVXLB21jsi8qJ3hsm
EB8DO9BPhrV43ohmdrgoV0RifcNolvX1mhqxGsiOJwPbbMX2HrY1DyL9CSPRxRzw
IXe192RejV7OHNt9gKteJRaCU0cDh5aFs5h6SFaNJYxRZZAwKk7T0ost43rw+On4
EX8DMG0iRGBzpdJ5ZyNG37yPNyt8KVGcqUrZvxS6CxK2EJdhImX4XRrfBeDa3ebl
NK8ozN/BBlcbiYZ9fEh5pJkslkUpzYTFvW4NxQhIhj7Y5f3j7BTrwwgjHmyK8gch
aBk/6qDmToO0cT7smTlJMEHNqlsLFG2z/RMjUpUk06dmw763mClYAJUmNst3umFK
NXVJxgzAqaB0Br0c9l91ZUDOlG7bwXQ9xw3iAPkrAMhlBSKfVyFmnjX88qgSwUwE
857YClrS8ZCjN1TNyxyIfOLIkeY6uleDdf8ETHZPr4yrNemVHK7HGKERxqwhqR70
UfUYg5wRcpMmjcIPYrWjRLgWvrMUWfrOYq8cqJf6lMFa1PjhKOGkbg6TYWyoelVw
rx4gIf4OPwKKG889IctM6n6NLyWHhYYHauicAdfpcpVJxLyvXVMO7IGuuWa3wi0z
GDgm4rrgauee2jvXUJJUu7kIlmK94BEs0vaSGOG1OjvMKdcrRwzTLzpFUAO5JBJF
EFEcP7JybY2DWcMxKkUh6Oc+kyHwg8d/Nzj0h7gMVHRsPVq45+ZYbhjSt32TZxqE
NC7ZRTN9/kGnV7c9XpDFUxyFAG8/ZlmDczW7CCc+B15U486dQvrQABHAeBJDqWDq
ZV8snlm4t9uMvVzTe/vbOyaxSVwU6h/6lfmEs+A9Hz8kT+P2fCkl1YlRvnxg9jTI
VSOUZFPCNJ0FgxVH5oJBDAO3tmuc9Uum2zPiNacoM+0fuXi8psFapPV+u/l0F89D
ZY6UoDoTqxQFdr9X7hxD9YzP+tr7n8Ih7GV8RzlVug9mlbcJFrzheU1yR3Oan1Av
wKIUZUiOzd1gn+b4D4VM11fPhGasQIS/r2JeG+AIC/P59MrMnko4m72F3qY0uH67
jb1WkgHDarIigUhz0oZbS1e4BrjZwSYHtwaYMu595KK7cs1doe/BawX6YYkT6Cz7
J0r+iiuKNJEUPjxGmdl8FIEn75HgnvoO+1s09440kaj3a84bmVg37K5PRodZYJJX
WKNRKEGLImrFSaSOHvdVlxFHz+LkIXAy1Mq48LEqbl2cT0FFGm6G6vKReBLkCdrq
ELO1SixL1necgEA+UPVlHB54oUImWLyQ7yr6u5KxZXe430lJFj7clV/LVTZnt4iL
pW87H3cuZRQGg3ZRUnFeqEtx/b3wUutBecBCuByc/6QV/Xt1qEUcqOkHgyr/DOfy
DHVHAPhk/XC4XM1yXbDa9dznSVCNX6Tma8evq1mrQ1wfYbQzfgMqpBhq3O3t5k0x
yYBg+W44v2dHJRsW1mj6DGeEWr3+wr7JyDGJBCH4XHAjFf+MnA/9MLDDgKEbi7vk
EVZg1LJS5xC3WdSzrEkoMxiDBEnk1SjuT4d1Kjqa7W+E7cmhfECq0HtTXTIBdtK5
GWrNcD2XX3k9xSirfseTW90OIRL9rZxwwY2HCQ0qjgNAupu3vTyAcNwlA+clAEm/
6H2z0kq+2Sh7JWVRiWm7TD7V5tsJ2CXYaaBBwH55Bn13mjqLP+2u4dm9sEpBF5yK
LTB8GohhYQqfZykNx8oruLvA5NWMrnYSxbGmX3rVfRP/8p6uqhCtg/Doh95Dz8rH
RGbB5bclo1yZUd8JkT8AjcnHVpk05n8aEadOamZyFawEyN66GL5cJpsAKEO4/4wt
LeYg2LtFx30SSA81R6fRY3Jj6Xey61XOd+xNUwThI8oIvcIV+G12tKKoDmUOkKtU
3Ctmh/egPOD6ADNXAkx/R4n9dB+vTJfGd9kirwFTzhW0cRGX7BfphlQF1meoqjn/
YDZQTtLhbuWiDVGgekBgbObq4LdsaldNJ6Ipd1wP5J8ad7O4pdXMso5awCFqb6Kr
jEA4plZPChruHmjdBpaUomVcG0AOiCGHaVhxkYtqfmOAFzwng0EoAqTaW9c30kUl
D+6NUdlM8r2+MsUeZPeejz12MniYEisclbhCa9MihhEFuZsR2be39o5YKVOcxrMF
lY1AZKnsuNNBY4/AuoQ7EUXuRLQR2B/4FdBpnb8Z53jWyVMzg+fCPNL+xdIeJJdG
iPIAaJ2VUx1pLHPLz0MjST6pg36+H1+AeOIBP1cDxs5fVpjIQqHNo3r46ZfZDpmZ
0Dze6Ss6CZP2t0jvHXzHVoL/8AhJpjWPf1EqYuuAlkjADtaYqgVCUvPLAaXbypTs
EFOza4Txru6vNciY1kOqGJfD9/iDcKbjbqNEAFii4+qNoPmEr/YvZVs8Tc4DxRmD
tOHBOhAKD7o/5uykpyemnjXyPuZuPOX5i1ihg+WywdTWwieZUtsUe7aFn5dnUZTc
9qkYkjh9mPJH4nRL7dSRW/yT4FahEmOf5rMaUVrWWGBXgnlSGNkFevsvbHB/aaa9
TJGIZStMnOD+4PHHwRJKDHxX4Fekv2mvxqnquXDb6W21Ts0LuaszL41dmEMTP0NZ
1hCiGjqwVRf0rGy27V4m44VUFN+25ax/ST8TB+2EgBYwJ7AC/9hEH5n7rYRXQ52C
CQZZmFHoKm6AoE1PQQMLD5OKZtR5FiEZ4LcYkmdJEB1CerG8gIq8pLe9baHB8pCa
nt51aw9KIOMjnNi1iJeupGJjXrBAjNEfgvWX37FXPGZaTm8PmQjHgv/B5EKdkDU8
BsyzuJy3AB7oj2QXNS2bvT3eJL0zMmzVqRoUGSj1+Eo1rHG9ET0OrM+XM7cd3SSN
rIHXEso5/9uZwrvBnVCPqZ7N4MRoF320viNDcTlHRNag5Z2vB1Mog4qxLQ449GIK
E1yTSZIZWAvEtZYjVXxW1EW061Q1nneQZsFXUHBdzwxMUOsboehfOmxnoqVPZPHV
7WeW/8t+QM745bOkIjPEW51/M6GSwmLqp2x+sa1gZUQByEeNv/FzQz/f1YggR4j5
7bDpDKqiSqsaCMsu9bBsT6LCNiVJTynfcITKqtUsMWGwDpz8R9k1JIOIMYNNSkpy
I1DqNQno9v/jRVWcBTaHpmkfZsPGCKz5Of1Q6ckMN3p7AK1cAJJO8hcfa3RQmFTQ
yOeL79YVloELrlDpU6I3SRl6Z6oi78J5xs/GmLhB4+4rIMN3HmRqZ9F2s8LSlS9G
rPCoE/zTCA9i2Zdb7hJEpW9GMH3gHoPZb/If9hAbMIDSTXG8cYBbCXRVninFdp6q
ttYupvh9SD+hctOIkXkp9G7rWB2xBpreJE/rQuTcKgk9iIvEzhyG0wwR9TS0o5Qt
AbKMcsqS9hTg1DOr/Unj/8iR9tziI9BvZ/X9HsnMVoCDgRmLQhZ3g2Obzty6SAIt
7EEWPBLUyuYMPlEXV2Nu0l+ye2dUkCT7uNxZHzGUkL8QsR3drIaiIOJsLmV5fPv7
qgEsrqwHOggc7xUvKoXpRl5vE7iAqd1ALSVT+rLz9YC32YkO5Mv8UqPYOcpHVvTQ
o8EV8TnwYOJZjam67iYlynBZpj9e35BT7u+kxXp8MPl1FItpa18pGwTMPmqjoBRj
vuVo8bYO/tQ6xh05lIJ6NlR6IIPKisvQPocSqJaFyHmzEknpa1gmsjCYGiCKaNoR
Mek51tPkbHAOLtBz1kJRzcnBKbcWou3vB9Z7Tr6KYR69RnZL3QetzVPTs2p8/uzT
SEKNX5/e6w7lKLwMrr+rrq+ddHmlHLyJIZadzjewhZBT8hrbogvew2s+AhmjVO34
Uw1ybuUR22uCSDUVkDern7IFRRwSPliE/h6vIRJbhKl8Iev9GWqIs3h+wfBOfsD9
yjDtQ1boG0AWwAsQw7lSW/tUhLg2o1FiX46j77Qp8fUMCSKjRWfI+1AvuaCp5mvE
J6wFP8HMdu6t/YMl2S2PmUvAjyLutmQyeDrtZyAg5gjDioAyLag/gE76KZii+DX7
w+DMXFXh94u1s+fv+5Npm9lnTJkOQUmAxh5hQLygEP1cCXiJXsWTsMZJAX83dZO2
vur9mFJNi3iZ/QqIfRb3ONmsifWA1zqaRxd8KA3lTwV8jYT9VLQ03UzkUdzLbGHQ
lG9Fu4po+qzNYSUG8dystMZkRMhcO6Yeqfre6sLq/h5R0pSYhM5SdtNeXnonArnb
IVSoED2yKzS81gsWB9doZ/FApQ6YQ35vOW8l/q5jhozxfix4dmmU5jDbHUi8D0ci
+DDPrRtRwXmOg4XF2fnQ0Cz3rjSADeRMeooMGMCAzV+QP87EkOjmJoO1Z7ZlNJTX
3xCumNCIYMOWB2ho0bh7rKmsC6EoBHR9EGADV0a2XCW85XzTSEX8PwGIGHE+k1cB
64X8FWImdjJfHUHtluMUwdjAtpFVzGT6gfDt24DpK4EGkvUPfSwgGta30PhyxoWu
Ea/iI0+2fAbfSiuDjidgx9bpMylTZjWCcIOiK7qj0qcIgD7x669ONWaQjT000l9M
yuxFL6xmlu54D3xKVjO1otAZM1HKhpcXSsDj8DY1ChwoCQq/W88x4mwVDNYkimDq
kfeYz42VIkPZc89kfk/OgtxyK+p6cd5kbkKbgFLbGHWHDhyGNanl82zcH38DriQ6
Ni18lzpyW3/csK3YfJjx66AQgk3iZyzi1B/v0whyqoSmfpDtb6mjb4J07/FDT401
9z13QXQ6/mx+kg9bsBLORlKLUAGqdrwjqM+3t0i123BQpBEbEHkaRVVgTDFL+zoo
8rP0LbC78Gai7hgU4Z8YeD2TE3R5glJOpRV+VPaSlHPt54bJxg81rXLG/JNdpOtm
hgcAnO1ElYbTWx68FKLi2k/4VpSSCS2I9CVpcc//VE6LFp6mgyVJIak8y7rRBziH
8Tqaz/3pOv3Y3l5hkIXXNHOJB8XHRktxTm2t8UHpERAzRtmYDMEgcfz/TcUqphMA
jmKWGf9j4QWfi3Jg3E6DV7Aog9vjQ1YT3NqRxFREU5IG7NL/dsbIeGTZSccEOgtt
3qb21/GZ6wGu2ew4y7yDX+y65PHwl61DbJwmSgoFftI88+rXy+2Qa3IpaFZqFGRq
k+RQkw/I+S2JLTUDkJw/boNoq07gOuhpFD4OmnqX5vUIrxV3NJSfIpRh5pbs0jw4
zLjrpaLfude5ylnvQSi74YluOiNlh1+9CG2/02UqHvRn1R/ayhdf2LKshouZ6Iuy
sITw7SEFxrNkWDiwJmZBG69UbMctVniMQUZWy5rDAzdBswNn0V9ymiQoIrbLHpG2
hfpSXFfPgLmL4v1oFFxVW72FZcBbFbrYvZ8HASnlEM0WETL7aWqK4KXBxzLT7SzY
WSnNhmO+hnzGR8R+QAIsE+zLu+XMWwlhRKyVX8/4AkG4xGjqgqrRlDCgM4NAobjN
lPDWBR8g4vnUwi6Rvc0ooV07KAnPz3oVnt5C2mVn05AvewqcdhQEnqvnSoyYUSDx
rSaIrtfcx/fonnePMAk/vpvv0Kg4I9z4ac2ePgWOuBbIbBHXA0f8gumnUnVvfsHh
F99pnBNw3i2N6/GMVV3gfjXk3JueJfEbz/c4QVXSjIC6vc/Se4Ns6hZiie74nJ6m
zLCFWVPPpoFw6TTgmwFyFqaLRDKR4vs9tH+qqI8tyTRQltSjYK27VLtKkzrddYWv
FUN2d7ScYkjQT3jYDWc8C8KT0ViY//9bOSyaqqs0bJxH/z5uDIGIf1lLLuK1c2Di
++bIK9Z1kb+DPcuJ9xxLWYRIKfxR9f0aUdmKcoU/rsF1An1kM0/Lp0nT56hW/0Gu
6taVDtBlWK/AKrM7R9GIK8zYnJO4zy0BGTtYErwYJVOLAzoV5erkYiKnsfJW0c9I
rzCIwU+VKOzGmgaRy5CLxbT37GdJCjpPdqY35XWK2Qb5Gho4rNzxOujk4QXhqZ3G
N6b9DHBo32zC0nfg88EYmi5OOARTCBqrQsuInqjyqEsqlwLfLjp329p043HW876x
0S+iHGPbDa/BbNkaceX8xDnzp8YpaCz2Ymuut1VBMuxGxqKyJjYEkmc2u1RE1B94
DVBEzqhXqyFU6uTK9FsuhKe1Jd+8SG5E5teCURbBcCJ9AN86V4fI4pFRBgiaoI1a
kIQVFQCsmG9Zkh/IblzaJ5yATf5kX+2RDzHL1FnUieg57Ke3dfcdOhy0U/l0jwYf
7NlS8PAVAZlRwnUBPptzUlCKOfmkEWmHy0UnnLMMvoVEybMpG80gPkqmc389Wt/x
+A9EsrJv8VjBQsXJN4gCB6KvrqSQlYJCKkVHzYo14blt3FmUCBKPNXI4Z28fqGFI
xafkxus8WIxllVvjdWFbpZ9KiYOq1yiG5nTtaqVV3v/QOq2BkAb/ed+7drA9/uv6
f44g8TQXTfZRXTufkcOZX2MXy5cS/9PtyMceIJ3v/VbAidu8dFSseojnlOJ0SFJV
aPN9pH5uDEAKL5eAAB29TfOhZmG/5ee2/g09PvxN5kvM+54B6AYonSy50ZNXV53c
rvYSD4YgZrYHe+Ur9xLOc1++mHw4rQM/0Xj0FW4WrIy6TJrkVR0Q3O6E4aUJH8FT
JRHvRsUsMBiw5xGJUV9ewuB63iXVg9hd5C6WZ+HBui79g8ExaveL5vKjzzoMb3Ji
uNOzo74uUK6qL6XnOHHPvrTU1DUUz+n5GyRm/jPLxrLcyClo6FcfLqUNzXZEXp3H
GUOPNRT3Is25jggBp7lyB6RsF5E6YcU6WWLEhlgtpU69At7bWGncGZe+zn86qaY2
JUvlCPuVHa/8uM2PeLi0isWAtSPY9o14SYZTyxAQC6K9IM0m2QM5SjfnnZ27tbUz
yb5yI6TgqX5FNB1SvZfph/KY3C/nM0sKwPizjpBbi3Js2ye2+nS6fy5/LQ0F2mbj
aQkmc8t/soShOC/jMjCFt+mpbMoKAfV1xofsSQJkRw8Z26ZmwwjyZuoFfORpReqQ
jjCx22POwQPyieEaNKHQnZE1PQbliD1ON3HfzxeglVFfWKlWgjCX9RJRMoi2I6up
B1nOjhpK2gF3a494BIWOTv0vb+g/mHRRKWtPI10K8EKI2Xv4EfGYl5H10gpX/FCl
5dnpbrrilrEoE/xGRk0SzZTVKWapgec51ohciUfuPrkXlpGl2RaKFdpaAuMovWWn
i5G4te62JBh9Uizv5LPSw2NoMBMKpcalZVgnSVyPj2OIbyqr2KlSGx/ggIHcARLW
QQTgOz1zro8l9l910KHNNBMBbTK4ILNEJAN7N6dTBLCzvbHz7Djbh4MoPNc0hxwT
u2dOpgUw7PYRpxyi0Gqhj76/OceY2k8TvCca81iJaWya22XDs9Bn7MUY7Z400aj4
n3C1cTogeNHfGUVxeQBSw78nrnUVv6k38L/8jfhAJzsVADxnH9B6VzobDLEVXO5Y
o0ymZ7dp6zGd7ZCVUxVTc6NMxmAw8RY/q3IjfkSo4dBnOsiG+SD95Dtn4N379/GR
M7oAiZMljnIy2gLQN7u7ysjUigxmYRRvE5ogEk3NvUCRMtHXbrnCQz3nraLILh2u
wj/q8cxuYFdKg9ORNlJ23hejcfop91d14YyiSx72AmwS4bPtyyP7GLLpH3iVEZj+
0rm9n4w+A10LFgCaj27qleP4CXNahjt1ipCJy06dNuX2K4jGfO0c3har2M6Z+t7i
mEWB6i0cquzjpwyzv0jyItq89qoUtDvX7h/LrUlvfVTM3UQMl5Je6T9E1BNxUB17
95bLPdmotTMxFJwoTFB/xgGOcFiT54yMOxAJeqcLzst16Hl2flV8uPwMoMG4mx+V
haW+yg/MOadccxLJTVTOr7IfRd5ILC5Ds5iX/iYId+22bHHrFB89lkMrlkUllU7n
cWp5PAThYoFSJcNZBbivrAAfk9gwPaGCDDeBm/JypfrQfcQje7/XPfxtJAXsf0FZ
Imb8kfMmElikK6NJJEYtIzxhtQCzeEFVxViikGGVvAaYiJtRE6J2evxt3Ygn02Rp
44N9ZvIgLHQZVPIIzhY/+7Ij4yPffjwyNhAhxXA9234nF4JrhAtFCwvrVlVaKYs7
sRyrwQAy86hNnu4yGnL+IgqTf5kG9711MwJrQrWDSS4wC8shwzqMWBf1piOarJKF
rLxnzTD/uP0de4e7OV+SP+xi6MNU3gGUVPfJHmk8Bipc+emSAhueAMdsDXtE6Jja
p7tp3Jrm4vcddCd0bkRLUUIkaqun74vJaREajHNtWGO1enuQG/yKb9QXDiklh2y5
bUPMt8jm7WWkJfDfLTwnvOYfEQZh3gkaHQpaWafruaod9B//yoF5iht/S+WVUxR5
ZQ4pn3clwBeUuoO+5QAprd0SpjSQRT98Elc9GHBLZBv8rXnDqp0f+dsyv+1K7ZyP
QvKAgIZ3bmF1tiZSgGhTbU554/DC7/rdXsrVQFy7R3Tr3AqQHKemic0XmWdsDv2x
R4YYESZ2H8fTzH4MR7q+X+nwflQsVQRGKdbX5USLxJKbYI3o++bl/WJ5vSyVU5ad
GyNUB6AURK8W5gHK2epT8niOCl/dPlflYQzLwK6Np2fbF8IaKMpTPCzh9J1ghvDA
cRObMEHNa/7Xm1zFFMzal8K7XhmBGcfTXvkGn/Qrn4YXlUdjYo2l0C263OJU/0i/
yx+pSa0DVcFpHHnCGA2ZJp5ISSgPjITCoDDiMjhUJgATaiQgcY7lmIgBJesh/DRi
qgLaD8Cn70z0lhJh0qqhnCNsH7GrreQV+2xLUE1Kwy4rvbygPce3ufjJsj0eDO3n
YArL9srU1NukxQDhu97+fZ8AO2Irx2wuP9+CTOBdhZ0A419R93tK9mzQmCKVVIAw
VZIgkKO32S6joD0TtBKzIJksu8rxs1oc6gIq9h4idF/NtIgrvhOHnuNFkxOr4yB5
Y/eEgj5ad/sN09+Do9QFSswNDQN9Na6gUjTVLOvXGaLKvnUl8B/4V8B07WnoDY4S
3iF5nyWXbGcF296m/BvV5IzLbvCXFR0bP1aHEtqADmBOeCOzXQHlQswH2KCD3lai
ao75PiyCbnds6xeTDeuM1H+DYMpeYfZkj90gLtNnKu5vizKV/heJsbUTqebhQGsU
/936Y/hCrxBRd+VVha12S6/lg3aSvYxIgubyf6A8tw6xqEyjyfCCW+Gf0aEFfFYZ
5lSW7wghAHMnKzDNMfY0Fp3roFqVsYxOKzxC7tUZwUyma/f9n6olMsuVkNClSP8g
SvN5GnauQWrrQLR1SlIguz0X+B+KO9uqv01R6kWHev/dkUxvM3i+B+AVTV6zc88r
A66bMQoBmQvHxVpQJ0y3zYJW64Nl52zcpXieObPN9jIFz7YoVW7epsE02tA3XSHD
ucdO9ZtHNUXpRcetcEL6j2yic/wz8/Owlaszw8N5e5m8aluDMIqDt/KL0+gRd0Z7
AvkgH5EePvYgqjv7PYywu08kjtSrrybNThiZ3/+MX1FOXJr8lDjh7wSmi3NYIr72
79kLZl//UJPfHSLyj6wKe8+33VGbaqP1B5fYYCRjrSECBUENn5vZk6UlEypaF8km
KHcVcOkTre7Ii4ej0pmT5LUkWGREyoPd4oQiMCXxfzkVLg39t1cgc9i03CaWBvu/
B9Q5SXJs0C0MtgqlzPB9QvdPjgNvVoc0gEzJo/JH7qlkbOBQnJbytkfkYFRcROau
r46FPWcNSLDdGsIYWJUB47HcUvWmJV7dAx+FhXwrDS7W9IQdKupiikn1GpD6Hf+m
mwvjJHsZ5yJNFR0QVJVUTTJztsOC9C4Vi3/lFLmcj7eBp9+ZwI83plCwGFv9o+rz
zbDQQUjM+WV5UXmHtBogdRPNP7n9RTJzHf8G0EMwmbnwKEcNIoII0ZN6RYyGYZ1i
aiH4OSM/9bsBiYSct4bl01kU3TkE08io74rJ2byA1HVIWg6D5p9H54Swo9Jb2+jj
Ycj5E/XyJ5cm+QT+EmXJQstoloHhnQC3/I9lr1+K4sWJzd3FsWZKO3Q7otYSF61/
iZ8Fojp0wWGELjI8+IAvrneZ+FjxVvqxSRrEZk0tYzyh5AD9vpjFTj5fdLeA2yvt
GfbLrHa2+/SnNivtNDk0lNx86IuFw83s+6zho1PpHLb0G8a7/wUwTFT+yP1ea1oI
9ho0wLY7TGbeVXIO3YaQrMJFNfad9Y1eY33rTfNbVvQmd0Lseit/WApgX7XIGql4
G/aAVxuYLI1rVLEAoUF354kyolukl0Y/DyP46JJatDqjnziMtqZIpSDkCKSFM3dN
omBaj4aeiWnPDQsSiHWdLBjCIUFBVpU4/Hc9999ZD4MlW2I3pTucW18dWNi8cSS8
lqUyKmRIrYQ8wH8UNKEFXYLLE0uSEl91rt6lTpcJ+piJhLRPg1KvdkZ47NdZp99Y
Y7WlxP7kobqvlaFNjoS3kjESGjMm5A/0rV4/0o8tnmKrpjgTETHO/nfGeys6esTg
4ueowfGSeUX5OldDrNL2htFShLVS5kuhkCDo4+jwl1l5XqvHQDgijoDwP8DUXyLQ
dBw47saNRPKWAxmsavnnhstnipl/HvgQZ+OLGs3ZBMOuuE15IokBeRcAT309iGA6
FxtU5HMqzP5hpJoYnOYUoUZ0m8p8Qu+IaD8uzrYQ1w2jo9TmJoLDh7sAsQEkKWjb
s2dcm4E7CNz89vY5Cy0KGaOeWYYeEHaHNcflBSFLsorSgp8GR8+mMUS16Wz9bWRB
oESgAbbYJDFT5eBVaZDjSqeFmXPKcqsa2ErM2GbJfgVtbrwYUGJCWA4oc5hpZ/+n
o+Nsvv6vd49PVyGF8ErbKyx/+IO2mQz3Z3YOuWHDoGpQSaudi0XZj08eo1P8e3pt
jhb9TkYha6sbWq7AP2+0RMZnVchkN088BulAY9BNfgCwlhX3xE10LzRhG0z+w19C
LcqYbOwV8ORGIWJv8voY8us6HCPUnB5+VpKRZsqvSRx3gPn0rIWAvxmZVHqpnWGU
D+7Ll9ElrlDOepliK3f9nADl548XveuZW7Yv5tXOLZmxt97gh3XuDDh0ByaQ+Qq5
moaPOTLvo35mQKyDeGaNXYiRpppnkoGKivy5EYLE2tFLA+5fzV9ojdlhGLofN1td
NOZcx55rrDqPBJ1B6IvUN3vO/dvlTs3b8wOuFmAirS7SLt12v5p6Wo1qmHdv2vYR
+9cwXpbhBuezw7vxPNSlPYbFX0904FBWuJF27OY0mRffcUs2cwHA7jqBsm5GeWLA
mmnbuuAzCCxkN6A9L5rAvsSjkhWGdjqEF2HIG/OzGrf/LGKcWCbMzEUTZYVklAwq
vgpyIRYsEyGnvgkSoDzNrJq6HkTTjbMP8z8720fz2U9m19TR17KcXFvgWBKPIvJh
R5v9fstaqEyZbr9rebh7m7S0Vs6nkwXt0+eCK68S/6/FQgTCs6i2oq4liFFHzfaC
S/+D9aLPM5ITOtMb4YWwPAlmeFlPNCBb4c+jitIQ2vB2GkfF+gCijM0cRbmgnl+d
5smqlj3wrQj3ZExSzaeh03/mVi2M+p7uVwpRXcFcBB4w+4RJCViw0YL0jjFm7aSd
1NQO5Q5nDgiWq3PkS3K9TL5SRXw/8Kyv6sztZp5QMboYbTsfHC59SZ+6BFiFWbIx
evcYvA/qPssUX8G+Dsz+IjhC6Fyn/xVfVZRnr9L4DAi+smQljrdiiJfI8giEb/Bf
sM081rIlG7pQAQOAnrFkn6ge2XxASZGiyEcVCA+DKnMzsMqELbuB05Ynsofaahvb
PfAcYAPdCcPpGgjGFc+AwiBvtlsy0Y+SxzsAiKrGIgl81TiWjJhEfkVQx63oeWu+
yVyfnprnwbUgc1tYyoXAGzJfSVEZfOspX2V1Zw63rRw3EfCTc9mTsOcDfPEObZ7m
mAh/7sBzOLG4S1or2ltIf5EUHwuWq3BlSTKLzilM3flv2UPxPP2oZz9UXWvMuIqX
yPfFqMP0c34FK3qV3uC2wiieq+08luxyItrQSYoQM2O6RTt5XErpYWZtKpLbV4nI
vtwGBvqTuRQeWMRg9d5f6RlLKaPY1MCXas3QIc3dGxx6mBm+Uaa34HI7xc+KQel6
Vdm+FD8d4NEp7CqjMwDopad7vwpUvgTaHcnenBY5B3QeUSHXLPgFlPSIwYWxFTJH
TmxzC80daarUsrwuO27C3a1TaX/SlKwl3x39O+hJwZgShOkZAmJ+idW26TE1F8Ja
APXvg1733MTi3RYac+LZ9KtXQokKeDQ+KDyXFmvUKNjgfWFcXWxZfDrDl/Su9lJX
g6yz7DfFrbQjVTWhdhjYr+a6mtFMdBd82ZkuDaZkF2AwQVyC5aJfJH0YkpLxyD4J
vvl6S+PrufpZYhjbHh0RpM2QAYlcrOJSAbAnzvkUvZXkb74KG3WY3P4PMRUdw1/p
q8c1e38Z/c33csIaZFigLsKdvWaMx06okLxBQT0F1ggP9ilRDYwRFiaCBm06GQkO
HOlJFQpFa0imODor6sUPd00INBI3+V6K1okCV2VaTdRYDmmwT+hfhgWecDOKkTIV
+NhQuVqU7DZHgWUumyfi/5QIul4/G4VE1gCs5Q6LKneDOY+aqpU3DZgHGMXHyqRz
QadbpQ4ZGf0YeKJFIbCeNOU2NjnBD6/zSM+P0tdIsdmEQff4Ko9p+sVCMA8dXezr
AqtyL1fTThRJyAll7P4/WLzgJyVDM0tZQ2S/pSX4SzThpu19nGwxIjkGws6vMH1f
972Id6i+N158xnXtqJQhY4f46plbRDzAG0WLpvrrZ57I/YZaCrsOV6H33IrXeHXt
Mcr/3gU/vCQLXvIHtzWQgCGFulpITvahiY3m45VSbsWjRsF4oGaut0+5nCgy/omy
hIDWSckrJ0bda3ZuNLDc9MLyzNkL/3MwMuyuhBlrZBu6bKvK17ZU5olzi2rzyS45
YV6y4H74jRXMI4JcS4mOpNc/YScZOnfg3rRLWfaKunZUOu5SBRqfJ6oDjAlSP/Fx
fE7MElxaTpzDMytLC+rz37TYF5SZjYL+OMij46HTAdTuUnv1g9lKaf33KS+X7BYo
1pF2hNyRyNMdVCwzVBpJ5MXYjWcO8PWb9fMEXIDvyZ/HrQMOCMTLltpqcqX0m2Pn
bkBrQ0P9W3GQcQ42pgIkwAx1rB+JlB4g8CEw/d5m2uQPwmtzh3+d1Co8fiLMic3+
BArnNw0pjwvihvtBfHSQ9IYXlJ0bnTKS69LIEj7DF31nAGN/6lPfHLi0rFgcli2K
swxbg+AkMC0e2Di4krflqufAYuErRtUCjVEi/o5AidV5PuYKZRIdYxcBigEtRVJe
dvfUm/oyLiBBLCOYSfbdfF+MB2TSCiXmSxStt4A8EOBUa7ej5p8fkaZuhcYid78w
tz4gsTEH2nLd7tl3KS8sgPCRtBoFiDW33pvEytG0ND5qZBT/MLaGWgHyoj0fgVsj
93Bxb9pYeZRcAPsQGw5uudodQ/x3ZjoFBQZh3eZcTYRB7m1TELS9Q7U+uPoK+rFE
0uojFoaFj9j/TP5PK0mvAyqs71gK0vYEZZ9NBvxBS94wzjp9MirSFmcBwE9lxLAC
BQkKIYMZCv8QO+uYMBPVfyb9BiRBUyNg5voJbYB+x5PSThktj/62kWscCSf/xUIz
zqulfx1JWXDK8DitV9JFldtt3yKLVPaD6XtwMvsTspovJdsl861O1+UHqzj17epr
npuGBad+5XUAFUJNdEy4hOw8Eaf2n4gPPN3jjcCeJzC1jKJ13BE1ByfypEvQwwvv
CeqLkOKWtjX3TleRhKBhmfiy0kpfSqfNAHzFUoHTN1hEl8fyoVAnwnE0fowIhMIc
2X2X+jDxFLOEbTlJxgG4T+lN2UQ5kN+vlyH4OBmVcoNaamyrYFC8KzaXKbzY6EGk
ai1w8pqZh5l4+5pPi8FrEFiz4mWDr38ngo4ycgtPAUhFkoh02Zkn6wNii0SmMFE1
DeF79VRVpAQ3sPGetg5RsHeX60dnSV4efsIHwM6XoYBIUABiszatTaqpHt2KCAzN
wG71clPAjRGTHsWoHxvFyDh0+P1CRHUA+7SlZaVImArtF59o4I0LI67eRmnIOS8W
W3D6qgCaYN5b3VNoCy+nq7MII7IGZKTal8wjZnxWyj03s3vdT6oWLH/4atL9JPu0
iKCBpADDxoxFV82GRRLHf63JagXv8qMaiKfBf0aUcSwO+u0IzaJsOKPyj7Yn8rCr
xqMlpEOsop7QnS7yk/txZSb2aTxAzMdJaKDYVzvqeYEAYtzMLZf3ORyXqRHfkjOQ
bKHu5CTxVX1oAKUXU5ScBOSLUbcz48aNE792R9Gdj7tCivphqmaRop9d++xBQWBj
BSJn/uJhfsZ+y+GDixS7VGFYGo3tAkFZ5TvQ0b/CVF9iz3Lcpue82FzikeunBwwi
89MuIxMonnCsEUA7CR0ubNQPwCI+O2MDOzXODSSrizvFjwYj9gOty8t+YDoabNF+
FXjUXR2Gk0+ci/uq47oVzQVFHFcSfcmG3RVYXvKOoBF7UGCW6SPyHpd/5zM8q2rG
UiZM89aZbIFooMi9E2CeEoDXVCVhtlSk6SgwNeQEbTVY4ybmPTjx8EQpcOa1Ckdl
7wDIjny0Ma2ELaSO6zAOzYAnyc63+h1/FTYAAkViGTp/j8jor8fXHoSKumVDgwpJ
1n9xJKCocMnFGhBGc5xu3ro/+sEZyk6/30D/ibs62GQRdh+EYkR0rI+ivWkJBsA2
59INI66+/bZAREPJHxxIP3dMcd5+mh81ePEWSddmE4vSPl8oKxiFMy+juFKMSDWq
VoLMKyjtbVMBXv2mOR7qm2a4Kfkl5BkY4RGIvWk65feJWqLlTghXa+apYCnYshgp
AyRpi6kEdM3dxjXDv5vYraNanP1FKqqGGeQEICb/fENP+aXQ9LP/cJcX8NCzDMsY
nGjZ4fBSxUxN9J3o5EjDz73KqL+jShXYSyko+MLfetBIzuEq08uen1/J6fVet7Bu
T3t3JvM+HfhKO19f6poGe6k6i7mObjGoOyx7w+COWeS8hZ7UlaZlMINkcZ329s6w
GQCgafFY7P320vhNmebX0N7iv0qm4HJO2eeUAAG4QE7B/SETGGO5D49l5e4ZOUyW
XkD2IW4ytqGETZQXD2upCTgauqJDG8nHUknSMYY9pvKEx73FztfN6771S+5xQ1T1
g7kzjO3S3AeUHel62pV8jCNFtlvwByy6T66tWsOxbWL8oUsRxdLuXlSTr5aQh0wW
jdhtIBm/SUOBKUaaqf0iduaSa9HjoD5EXqmY7RFFevwAB5al2GkTWO9hLvEcVqvT
JtKD8BxHNiTo2s/ENp5BYPywFisIBAcT8/rv7G7zWVYEiA4Fh5RYDF8LQXRGLjol
NuS6AGr6Q//4t0p6Qd7pku3NVvAglViBckhnCL5dApkzQC9luF2Ng1SHBoQWF3Ye
YPeuMbsItm9oP9UgRZz3vDVZ51Rc+aPiQXGawDHP/xPbxkEc2F9OUp+ZWGilnWGk
7uhIv1TWrNxXJ3VYSXRQgzysR4EGVdk58w4y2TILdYzQqhw9l0uu6AHak4iNzZPy
zDa45COsLBnBP0ugJUErqrouzfml4UEzFWaOH3lb6wkjV1rX7n33wZZGLCbyZ/zS
SOxiRs0XYQxMLKRNZdpzQHV3O9waEOsiFKkiMqSIxscwG1MpPTyRKM+TZyJ5V14N
nv0XZzTF5apcHaTD7RNnri78gG/uQN7yBhDZYBKpS+fNbIQrPA5BKPuIpYcK1gXU
tlo5cfURHV183IxeUgzh1S8B7SqUaaZW6XB1NMb7XSFNIWgSwEPvazxuKHogLBOy
cAdOXWrN8ZvD9bWhVYP98Ll6NwPuIl9uC6sQuWvaZzfljVacliixBddGVU/tR0JI
2kD3f37barX7tn3WCVbuKgPb1F6kLR/dShWT6mTAYI7LtHwQ5H6s9bcUdAqhZEmN
+YcU7uBCKL6VM9psdBhbokYA/jcub8rYL31fzh+7aDNK4RMtbIhG8SNyT/Hfo8Mk
2SfZ3ufbUqMkUk+CbB2X4u3RsJTNTWY12Nq91HxQwhJ45XVzbUgdU5BehA3uI3WQ
QWEmBKLzfR9/+6N4daJFrFyfXt/aaw3e5UZ7sfZ2+K9RY6N3YToSFy0liOf7XrDh
iI09E0SPLN7MFVETLFmv/qyhF7s/qfwehcFGf3mv/b23Nb077a01I1sYHWvphFHG
GeI/7pLsoypL/BWn9FiHRtIDV/ZEQ5BTqgzX+WJ+oSYnCUFqOpuIEy+Lb7Dd2Oml
XtsQ0Wxev2JhghOrrMXOMxos4dEDExBVzvXLz3DC7EcxItT7hcK541OuPeYAVOno
wLg4Ccv2Uni/KMIWKKZHRyXdX8LxiW6sTWoORsqllXwFNXW2oLr7oYqoOh9Erv5/
BSWrZwnj/ESHUG1VsUU0L61qx3Ez8gwfKHgXN71vuApjhU+jTqvATwP1GSG8Rdsk
3V4h7dv+cWGgxvLsvq5BMHpCDpSSW6BBS/JoH7Pfk6+fUySNMV+vuKRThMsovnHK
9UGU8/R7i4+UMyZBPULdk02M0f4Wg5HoPzRXX+6TknDZT+N2M1r6exR/ivS6EXO5
rYmXS1rjlmKV4VrgcqSFsoia/PCetKnl71hxCHWGjlHUm7/TQ0TMiiak5bO+jy2M
R/0ij+sCCTBXjo23KdauonXRrnEYbQx2m8mN2nUUnEnUDyzB1YqRCg5qaxwGvm/d
WsGX4AKFVvcTyKQn/cmNMCQvFgiDNvVMsPxjlYI+IMPBTVYF6fLVzucsDZYKV498
ebFCcoipp98TqQpuHHaIEZCdBaaNudqNoR4LlCIvUvt5dQTNZ+VtBNH76g5hdLO/
V7LQc779Te5uLoNUXELKROThxBF/uI59xpEGMIm6TYEw2TTkEIqcQi+3RHoVdefs
Mgk2uFrBijKYs+SoIRZ8YTqwfVIvxmRVLtudKb1QAlU8nRRM4yjr7xwVV/Zq8YN0
U4zEc7aFpQ6ojY5MgiEJHW60s5cO06DAVypWzGyGTRKSfWI+g++Ycxldlf24QCvK
LiiZzNC9JOg2ZgROKLOvI66DsL62T3TD+62OkjnTSAUeOfZ8HgELw6pmkSUetXO2
mU9X95mf/P6rIMUepQvRQVxs/NiVyj4fcrTqXCYv5x8EAJNhr2iMR0ICKW6XXdBO
H89hyg2C693DkqNFG8UCvl+7u0w7SJmd6zfwQVy0cO0Y+aFgFM3FUX4o5Dms2ZEl
gZIS+SV0zb06nGjEYWM92yIdiKFC3BPuT0TirGdt0DBZkBHslmxX31NJpIvQOhmr
wWXekexQT5EWsw1H+JQAU5sjLy8IJOihfmT0FVv/hSvDpP3VxkADHohBtgPRTV00
ktxOkJ/Dt0aF1mIgi6JPDkMgEVPuNAxJWU0oRGPmPv0/rbUdlyPnXuij5IFoLMve
vXLufqZloJYxDV54yqP4krq+HuVD1zqUb1nAFaxekp+e5OJpxFlwxHYf+kXfNZOB
ZMuHBBNumZaFwm2c+a9qG4RLVupre6ma0C5rMHkVdv6v5l+AsV04KoTw6OZtEHSd
Pnvk3AdlAHiX7nTGaZ+nFHWLR8/8jpTYzG1t03SH2XDqwOQBC+8WY1KYD5XxBn8D
xWFTmZ6pv0bHPfnahK+i0J06yR+YXfn2En9jUE0S7ar4uHvbHtqKeZaTPm/WJD2E
bQQZ+gVjHiSfEknLo/lWHtdVUVQdvns/juw3UYWgVBfxN2AAja/HMxlTzSZATZs9
adcXiEAaBvPnlPZAUF0y5d8oxr5Ljde6adUo4FDJZlz+hVXMKssjKepo+qqu0VM/
ZUDj4IrYpoqr3xhDyFRpLEkUb9SIrG9lcPDd4/sSid5Xb21U22Tnb/3/R896/xao
6SNcBECEXx3ubQHimYBuo3W6sn93WXDrmSoIuw+aYiEe+EJP8gpF1tsyPE3YJoO8
n+QGrKBpZxj+AMgHeegDNnSQxlpD0EdyW5rY+KEv26qPdyb39WaWjAetgssbJ6yI
7wXIL/skHwqsnv2kmUJKhZOUSRuz/JsWnfoNe4NgaxUH/Qhcy63Bfk93KyHkFy7W
LbXbjmqRNpfKPB7Pnxytu/SbebL2if4916ewE5626xD8JKX2huzUAqbBEYjBvtZt
zu1hnjsfTJ5pXlZVNqF9itA23EySURj3BTHTIRvyhOgtQJ6bxKAso6Qaap82mFlz
eLU29ECsavxl+OGMUtpw/PzBHVjHmzO4gYLLngq/xQ9Jh5l68vCNe7gASkbo/CRH
tdzZSLbuBP3+L/CliY36VE6zomTXfmKsO96YrxucfD5g7z7QV2ZhPN0XcdhgvMbL
a1ajepGr6JEvPbfoMDIcJbG9wcOjHr7mlnEFNyM7r4sIAaAoADEl9MpEDFDbIEz5
Nnha3x4U58Cl/4XCkab4mbXSyffvUsmFqvTtU5diqmGTcRwu1Hgu+QEafaK2jim/
EBBA/S8yVrqD8xjFxFdTUeT+LNmALHczgKOREwDdSlzpC7nzSdizOc58+Vbs7sI7
l7m+XAcyCx8/9kqZShtmK6ojlXNlNtCSg0DQNrUHqA2tw+Zd+Q/lYBVsaPQpoefU
vs/GEnaMa/wOhgInRYmyNPf6AZ0yNFNUK63xkFRnhOctb7FG3zK3oiq6EAk02LFg
tB//7DGxkbbPlOcSg7UnGYc1vab7Uh6boRKwSWNHoW0x867lo3NroHnsrrjLoEeJ
+5bmqSQjcCgY7izasAmAo3m/GVYogBmh4CwUMP3jId9rS70OKwG0KGipFs8dlED4
6r+IynIejgkahdUEa8IT8B0RJyMsqC1Hfbt+ldp/plsMSgezcbx6HIyNw6/YRqP3
3NZh60x6BRHbUFOKI3fbg+V7EUwWmo3U5LRsT8ZYs99AZDnkpT10NywkTvn+yV7c
/9COrlyUwxLgAHz2gudq41bm3fbhzWEn/JaiL+6ksCqYLLh28hIwqIImpm3fReE/
OIs6StW35XL6zEzAoDxGt/llL4d0pJyW+yX7nT7JHKGbLWj+yPu/bOBY8KnpL+hG
zhaB5aGr+3zQQyXku7hsAjoizePjC0PAcEOAXn2ZkCrgzMPDMxptQ10HjwlR3/Qr
hMGwaioSFJxqjpAwREYGpM+ZuiDzgXJxQ2m8r9LlpfWcRTADgNu/jWEPZcot9gMH
xqRzwZBT3i6xmvfE8LR/EXu2m78swzCFu8Cj10fAWA92XWmb2d+c2hmqNREPmPhc
trw/WY6gxOBXNgqKIsWIIf9TB2Rxmw1+fl1XVDxYTKQGf65ZYvmtL4MgaZJHrlG9
dnnGdkiUyITl7EHqcY6HTZ4OsXaxrBy9tkOQoAmO5zdPkzgtXtNNNo3sVQnrbsjo
VcgXyysnRoE/hjwbvflm2X/HnD2z9/0ZMryztGIJ1L7Nq4o2bUeczeRadEWq1Gmt
sZE2zNq2ngAgRybhT2WPX2ZiON+ZakE2C5K6qEus/8cN5RpEvbILZxAbnpm/r9md
NK0r3DwbCeVSI+L2j4M1nVYZ/kCn/mdp7ObryljQo2jd543K5cbi1PExf/twk77Y
oryJQnxftU2OJLiIl5/esUjarXYv9J3+vhb9B3BTSfm4bX/Q7MPk5VMIQRzhU9SM
XCgxHmnnh0GsIgyBo9/gUiDCw9kXPlltzTxdESSihBbDCqWcvt/uDCGMbXWHB3l6
XAKEmAxwfLrAMyKhDnegJAyJgmZc2hPzNQX0721KD4ZGgqF+5SJthOrq0POAGnvg
O7FeCkiVvJBMLJ1AEfgSq4Pnf6/8e6omuoEQtjDlL3SOUFCLCTv7kP4NVbCUdpcc
yXOPPZD1zjT/1iO4EeTG7l1CQqnEEaQ448ufY4ktkc79DOT8Tux8B3Fx9JirYL4z
nmng/BSpy6t6dtFDoBisV8tG3eavGf6F44tS8AH/rNNZjAqT5Fc43Pbsqn5LHak7
nzDNQbMZHdJZ8g1IMoYxROu+SHqWOke7eRF9zDB1o9y6GhFI6kSxR78k2Q3gmE9B
ycftvPNYSTTLPqOvyvOoZjdx61vWqV8m50M/tcQ407thugoOIQZVXg3C7KGkjAjE
NjC430J8DvH8+REHY/eoLd2unzF50ePVqftyJqm68VoU8izk+3wP1NIvUnaefoFK
HHMPZobbJJAPI2SFJ7pImNcJ8jkCq7kvhMhoZXV+aP71x0g/lTtNKE5v/JC/pzYv
ioYnCYr9ajjzXV490YJTvGqi2nQNmY6pMXj7j56ObRaDp5T3Arh0eN7cggtTR4WX
owS8Vsl8q2Sj08ipEKq4PqL3B3v5N+jGk/qhgp4gzEue78rEuh2XxY/qrkmkKmxb
17L4s/8gKjgwSzultOJmYTK+qyWOM/GOrZeQItxl4sNcAM1dB5vvVUxd9RRsiFgC
hrxm660hN4QYQv5PbEQJTyIv8lfSZWgc+5smhXdAD/L0E7EkbtlQV0ne8v1MLtcM
E+/ROLtF9BnPEoY1hY3Lclyv/QCrXiL6anBeZ5nQ9smLoq4HOF8K7ZilNqEZIIlj
Ty0VGj7nOvwy4GeRgfF91LBuvdS98rnLmpY3py8ibDUF5SIwZV9l9vKNJLUESQDX
tqsTa8byZb707jUHOwj1ZVCfHiH48WI18M/2IvGbwD+jMaDfKzFlfUUtHe36Aga+
V9VViyemejBU4gozJuoza6ZPe3WxNfn01XeeQL5dvX8KSupkqk+mVARvfdesK0yX
xPS/c9DgtL+5CI0soDDx1EjgpYYDG5R3a0PaSnSd3IN7jVDhu1AtqRCZntNI1+y4
eZbVpyfzQ56B0JqhGbkJdyTncEoDOl+n0qf8fSR0KUpllrLbhryHVY6Qd1d2AIpK
2dZpTcx3QQkKG+gVslmWYuVMwIoxOhOsIyGe1g9ytmWjAyAqK5Q4H6sv5kwrJJHb
h7xzDalCfTkv93wIWER66O1ptI2gQEpwM15VkTe17CIMhkZWOVarlF6O5hQOhx6w
2QiFM6Ei+pv62FlrWe1W0IRSGEXoIRsGLpdPIcUqUpwOdc0ylX04u1XHIpn3R5IH
1oelzckaAicCZ8YZjXS7H2z+PW9Qa0zfN2Nd10lVxYY71W2TtogfA8Y09PD6D4yw
sG7K2yR+fY3ucGWFHUbJGE4GTy65A+RmIqT7ICm02Yqb0Ez97uwhZ3rZqq86QONe
JvgbMglAN+k1G9QX4SM1Xu1qzEKPBH7c+KlNsCGuZESHDdKI4qvqdADFafchY+Y6
28e/LHjbkRrvhX4gGSUG/bP8AQitb4W7GWlPjsvfG37W8OAdAjABcH49T/lf7taH
gfujjGPwnlWTKBCt14pJosQuEidT604kKienXoQmpOenqATvAtCgR6jKLb9P9HEv
ts4/qcBRSDQp7qr4OFI7TzBcZGauA455PxEz76ViBgT5hS7NvT5KqKW57wG682ML
Yl2mzqT/HOCH2thOqWblDEein1L5h0edj22fmJTaZvxtukY4kM/IBkPexJ+1KYD8
KzeEKQURDSKgjPy8FcOjJYqkLGyNpTQpsHAWtVUmUpi+JMouwMaLYEkN8tg+XeaD
sKLubR1n4Q20DcGxc7DKiDN7wEjP8MH/iPVo7DekL2+wWXYayDBtLWsnvrAotkaI
CUmsagk8eBsdR9NeontJu0TcAFfdbci4mE/G88ZTGvhX8r62qdcA7Rppvb7aOazz
MLxcS9ZHQwFRvdSybati8icRUDF9qrHOiVF+8KHtQaASWf+B4rb1VgpQ726UTnBE
zUjSYUGsxW5UnPXazzR2Kspt9CdUigiLIP5Rn5tP38z0rOa5Qs+AZ4s7WLJLyT26
Ss0wR64Mf64BCOLCoHWe4M/y3zVkJSyV3AqnRy8c25pmgde1TUlVB9czRLCmJxEa
`protect END_PROTECTED
