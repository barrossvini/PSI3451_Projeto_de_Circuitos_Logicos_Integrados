`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HFuHZQLEtG6Zu5zyJ3oMG0TKWnnkd15pQSd14nQygScfRHhKfQUIsrOw1Aoz7e9Q
WOYU6eBzh5jxJa8KX28EJ3YfRhChdta/HpnuN5JsCynXjvSxKQaJLRV5wDMGsufm
5Eo8wFScr81x3cNIHpoEYEQ7p8twbgpncA/efeGsV+Ryonkbsq9VRgzYdEzfbdDr
192QAogUL808EUeRnr7PsijewXmxE4PLuAu+wnP7nF8ON1N0SkBSbZemZLzFglvf
E7+Il43kPMiPPTO4jGRdv/NhY99aDKWwgUu3g4IxQhQKrqDjpEcQxZv8aRmlIJ9R
ma3tdjVBaHBC5NKkkjWefSix9oiX7eSBLB/2xipcLtPMKv9B68oXGnNJSeBYRpXy
Z5DMVHmno/oc+kDyKPhUhxGGuJHB1TqCodyDSyhBqf8U1W16MEeqHSBK/l4KZAEA
NR+Ckn2zFUJr6dRTORJbTh9Pr6wQvvNfy/r81q3Nop5RI30X9e7ctdN9lGkC9POR
7fAdzLo5H+QcpGX/vAUZKbZpxObOu//cdQmCoqMyoPsly+2GoBro0b0Xixkh4zRs
NfTQgMztJ0AiTNDKRyCuxDN4N8kZPYxDDG0lLj2FoeVaKv56N0JBDPJD+F+UkJDX
6N+XP2cUfK1xwbztlki2SJMLJYsnsuBG+DDhHkbRnq+TSWdkYGu4LoIIVi7ev1FF
VwjjP7o3fuQnnHiY3APjplzo30kjTyq/Gxo+peLB3Mrxb39hRHjv0bv3VAIwuz9M
9xk4MQBV/YB5wkCkEsdqV7HLxXzGlkzkOMZPctJGBwxqoi1XCDcupEvuD4tKVxWZ
6lMYm92biEwzVOl1PRViMT7aSM4VYi8bfDErarKzhMSpunhbpvdpAcZlS88fXylX
3A+TKODweTAxqUhPzFrewgZu7lGbsyoZrvs5Eo7QqTaXvKk9K8fWiXl8u/OZ4bCB
mVEDSCEKYf4H2opFY7xL0CIkr63FqkH37RdlaHdvDH9bP6gLA0WuJGsPwNwbGzEv
ZN69Eu13xYVaEoh0mtn1O3oYiK2u4YGWBZ2EDlAQChDJnPsMfuz2X00kFfyE+7KT
V2QSp4dBXwZ4OBZyFtXKZA==
`protect END_PROTECTED
