`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q09Vpr9jj8rx2eEvH2kAEC7osVEsgu1gWNvBnqYdwShBbpniLWpC5pyI5VWdadX7
CSUNm6q33PCkSXFI/NuKfEQwRTSJ6cHwav6gaGZbyrUg9WSAg+t8/ZT96HzuB47y
37cXtwgeVKprxIiM8cR4d6HkjhcAJ+EMLR+F1gXkcdiOkh8a0ZLmly1c2Kzvbx06
YGc77t8YOOgKC2GpFjQrxmpy3a5yAr8aiXXeMWy8CU4CkVqvLG6+MpEkLMdB+rvg
yCXktkJPW7E3O3q+BQFnRV5ozuLJF3GEw3XschROzgW6FTN8RrP4VngKRoMqw0e6
/vfT0nRHqxRMAsiUnk9pcZ2KJmYsqj5zIRY7yWNxEhyFZ7xKHeC0S2hWxfGsV/wI
P+YJ0oD6DgL1dQF+7baUWil6kYYnCycJVvXM4mrdTOB0MrAQQeMmXwWeUsqUseFA
9lP/zXaZmHuHWNPyoF0WtUYixX67nIQXnJ/hhW7TZIJT3VPtrcIZtXVOn3iFjS4a
4nwjllULbLle1nQyJBd0tDmFnXw8OZzdQB2UrbBI2QMOBATUxbSqCdzmnmCYYokJ
YLEA5xW9JSpEoDW3zxWBKBao7HL7sbqKt325Qt7ZsCN/Kz8y+qGw1qq/AhlU3lVM
e4oxeYvblBkRGcBeCz4Kab71dUzT/ybORz37grfdyNVf0+8t7kizzzK9Mbo9G5Ai
sLy9tYpjII663aTXQIfApYzRa5h6HHfdrzfhPj7NI3W8N/eNSfSlI4LPrK0+3LrZ
AYGiPSe3OTRrl1OejmiT0VFmvEv6WY/xMknzp4PZKDXg5cxsw2aZuCNhykujmrUw
WMPm/3zmkHr2IBhC9p/9BidPcnyZ26QJRfQLABOH0YzTUnKOhK1Smmgdm6g3YwUc
Ot6r4zjv/WFnR1XQKt3RZjsJhzxwELQUUZ+TEqLHy4SN6eWzb03XD5lHdu5TalFD
VTsZtl3yNljCa33VkEmAP9BUh+FXoYNU8XDqfu2yf5W6GkyTSCtJ7nfdDAkQztZJ
rZQcjMFGgjZRobF3o1UVLMwLjRp2yN9Nx/etFZCYcQUlL/cyhXgnSv8xcY9ooMSv
LBdvlYTug0nzbH4vpZSlrkjkL65NcYwsO5QyWGeK9CrcEZBcg41G78LWlY6rwGtu
/xYKuD8oszgsIIqh/JqPgNhXvja5oU9JxuE2DTVFnvAzBrgKNmpm31vGAyYF/xAy
jxVAPMegBaaZQEaxCjJ5P2D53BdDk4tgUrJs0CCLl+3S9vEAAhcDoNeoszmlDNnd
nPGUVjsN18SatNQ5SoJI/oAVjtiYAMZJ8LmNcstM/w5tQ/YzVoff8uSli5FguWmf
uPiRB1SmqLrqvDxgouDf9X8WGRaQM4BCJl8JKPXqhSqRpAgLMZ25XD+I7VGnnOCQ
tBQ0+TEs9iqQien9UKGvGJo5XF9cp2DXqL2RyuiDjJ6a9oxQL73rdU62Siy2wknB
oVlhqG7IFUmqS6eeKcV+SwNIQRlj+NrIcNLXuUIeQc39nLhY0UcAnbPh+FkMlVhm
zuNAo3J4B5tIr2RlY8GJiphVL+Ac5O2U7nhIXPMpvkwFQnQruxUsiR3qc8y8G1EZ
Fkf0XkfDNIalxr2W4bNctmXpacymb6y2Wa9tgncfx9RCKXHk9/BssKOik8+hg81E
iKhKXtpiOgAnRV5V9dtCU6HErnKnrj189bgP0u12x7reXcdsn6TmtdlHYmvsUGWN
vohCwsXJ8x0/lc+vxXQka7rtPrL/w57jGP9zkX6eEhYTRtO6MeqALtiICj8A0+o+
BKHqTQGFNeYlb+yxe8A9z40mB66USYMpz6GPsWtI2vaSNWGu/o8jbKHo2xbBFGby
Ezw3LTZmk0saYPjfDG2p82PqHn2RqyAmAatGo8yhXoTDa5N4Jz8UTfmx0AIo8tUx
dbEom4o59cRo+PYGGuvsbXjGVQpp8LNpR9cJhE/1pxFhb43K8Zgsb5xpbl6ylqAx
lcyV1jWfVGZbYVbTlwQsQDGrm/XbQ114jxXqE9y1Wa37PtbJdFM4TBoTU3RCBK4X
ugozO/P3CnOIH1DdKmCqhzoVWiGQzUcP9UpqTpmYZVXk1UZQH1nfZcG6qxJAAOyf
bzS1PMHFcCN0WvkC1qtXZq3Tx+OeVrLjJYVPBodZmLWlGjrUHGcR49ysuz6AV0kJ
I3/GZTZEHdIekbhzxGx+BFc0N8zxrGPlC6bY1IrxOWB5+tzl4N+S19r5fwJSMw4Y
WUnqPVx4f7NGTmDIVdG2nWJEdgCo3e7Z53lcAaYOihBnjxZA9OeubB42tylQVAjX
l6V9qf6cagIqEqkbTJxFgyr9FSAx9R5ZeLyWhLWujMrGeaToA2brfxre89SwMHBD
KYDhm/rdWxqzx+hMv2BnoakVySBZgDBM+LEid/P4Z+LLW2173A0p/oUfjk427FI6
ftSlndWL0yxL1Wl3LMS7BME04VlFUnS4MfAnk+BGyo3rOAS+Juahsygy0nFanWoE
kvM58aTiFz7Zjj6IiG/tkyGelZ7KRfCQOj1A3SbzxdGNhhCofQvLjRfk3trAzNDg
nq9Td2h2+lc7fl5vfgbh+gCbsMDyUwyNdtLf4TAjhXVVCDkkaNIgVNrM09kc9gdl
mGpa9gmUWBbaN/uGs6dHIo+kJCNVjyCQf33UjxTP3Aa/mcoTJRWeLcxe3eCoQ7IB
jPgJ07gwYDi/hDRaPFQFE7O/kGgAHt0PIpzlOujTFMQzICDh0VeW/XCnv1WCzZR5
24bdzmh6bZU06nyL/1on6NbQBEuVT4U3BN6/22Osx/s8PgsXxBSwXtQhjwH8qAOr
lFa0syprjwS25fhdyY+XkJDdXi7qFdzUlZj4dKk83lH8r7RhKZTewd9bhySt7U2k
JtBd8e63FzB60psOp2g/ITpRfQQDdimenxafj+NzxEDW05glGOyW955bH8SBVZZG
4kMMkG/P8O/ohglS5/klBjsx4r1kZTlXYdIXwHnv7XjuNuCG5XsBJfrndx4MhYeS
i/SR2+XtpEaoq6KCyfIDFMj9LIjVF+NL27CvtWrh5jW7k8KtZiFByvDWZrXj/Vst
n8+9+pAzBh4pjIE9Lc1d5NF36n+ejEAolbd5TMi9kcIO32ttbzSgL/Qq0njQ0YZj
JfIvwCUsTE58xCT+WK+YNK2YpDWRUiIMJi6+wmHyiwdCUZcyjtJ/bBrp4Fj9P1vb
UbV81scIojFGbl8aW8c+EuuHhfYKJOR5aU+PhCLrVgzR/cQcmxab5wTcI8m5Xlpz
jV+vswYjnNWhP3MB19KkR4FSKboj/ozfmLDkWDVEbegxNx37gMJjBSbuOyWX5yRs
U7Uy1xf0mfFDK14TpsPZURi1hHYs6sRVG1xS+MlC7gDS3VVvJ32HazCbVrMTUICX
h6dwP7L8w4ZTS5Re60E6NBuklL8/BUk4wk1CAxqQvBQ0b3hGXdcjdxeVdPj9/nzC
Ax72blpxH6ZlCOfw6kxajDe5R/pWh5lLJh6mN5Y3j/1nr81aU3jnvUUMGmhrmdmW
rrONgUx81b1qDp8PjLeWwnXsHWAQTqbQQhGUbOrc3fcC3zsYm3LOQOYFe0K90Bjr
wnb1tBZR7R7bgthLIOwHVaLMOTsL4BE8ygI/FsURQTqW/mshCx3gB2sxpbnBz22/
Is+s0iBEIieqol75g6kCWhPbtdoIe9UmyfqKsPe36VRyAAOEe534lN59FoyhxcIf
T9R7R8n24SLKYHaFLLAo3EPUo+/WAVTlsRkP6yhV0jv6UN00gHZ0dORMfyoIAcfl
btfGxK9ifGO2dcC8iXVl92TUk3s4lNuKmtTshPhw05szsdzhMMRHCH9y3vzWAQNl
a2ZU8G2SOE4HKTdRVeuLqvKADswpys7XGoig9Q2OIBLShiuh6KuTOgEfRsmtCCjJ
6HaIHWVPYchR4SgRm46w7pareY1LZnyGOmbN/OY0xJId2UIeV67ZkIdyJsk6YdMH
15svFp/Dr7/HWkrs1yhozGYKbc0qNVk5sjh7tbAisX1UEUpGgts2Yi5YF6m7rQAh
sovDhIxLGyv19OkjFghNY5SZECxgSUEb2q9Mna2qMO50PnJTddgAxw2EhO3pRYp1
aj3sytjS2BfmRIinKT7YdyReRgWaPvBpHKGlIRammMcP9iWesWOMclbknygIiSUa
DQ/j9Z9WfByuAjokh29rs2hzr+Z03/UosdhqWA0f6V0PyJRbypJETMBznmCL7z++
AqRGiTYVq8PQ1kjTVCxaHhkTR/ofwKOtm6q2+gFJTasGdkJsdGO+ezThNKtLueyX
4ubezY4U2immjQi7rTk3cfQ3MvrFL9pzK6q9NKtQMbdd9FZCqayXorRxIpvBrXKV
oyEXXLYnWGEWvL9MKFqVgfT5vqgQRxOvSpYr0SlIauBbzk2kmYYepWDy9slwhlUn
qmonjbrSzkYUNRbd7YSSTR4D9c/FNpXZsOXMzCYq/9UUz0NnhgaP0y3Hef633ELe
peXjaUrrrqNiBX+bTPwwvAcS/zjfGPgr23ITXq9tSLJeKhj2sVaCX3xkBxGj1sg/
WXqZ/Jj5aAVHzw/I0XYBA61D7E2QKjwfMdxYlGDcy7mGDwNpldjoq2bgLVXM0zFk
qUPLly5809y9fSg7uyh3USMreNTtzfK0jI3IB9DSTntU2R2npht2I5SMIHczrxur
semEIWnEiK5VjY8UnqFW2LO6ZFlzN6ksNC4Vyx6HanIFhhW34IcIPtjBuzj9ymtZ
/9vrh0+56/v4OXtl2Qttl6w6nFh5MzqvOvRVw0M3oFrRyaGLYlNrQbRuNe8/Qr8Z
haSyfb2NA7NhUMIMVolxnwzt3adhGHPw7y3CM71c7gKRSzEnhoxjQQe8ICqEmH8N
aKXXH38ebVSX5K6oYvHKmbA8c4g7xwZv+iR+eWvEjnYbYNpsiqISrChOxOcArS42
mya6xRu32r4M5EbbKUMEuK/egajS0VB/KRGphRbCrFsjwJX/b9ZBNn4FkeyoEM8y
kyfgAL2oRlJvyA8WLroXmXZUKBIXC7OBIRfRIOQtC89SHkrfXrOGanoe4uy95eOK
sSqw7I4m/XN+DfdgEUaNABNNLApBndM8d2umGz3lCB3WXqR/23js/AnIxeTOwkZo
0VNdwxsUg99voiDJ4S8xwQZbJ/AP/iPtjeXxWCyeDRV/TfO4JRpCJO5YoTAM4Li+
Ns0ovIVeU92nrPBInUmhYQvLYaTfb6UYsQ2nxvvKK12pgI03LRQNEWOQiC/wB387
3f4EYwlB+w4Y5nWbWyxA7HWh6FtLwO0taMPGrPrMPHOVOGTxjXyxpAhqXUTN59Ki
gqZVjyW2u4eRxAfK7gwqi7oTxusQayUln9erJJ5wunB0pNP+6b+3Gptyeph0IP/V
J+3kg3XN3p5qtquK35UOgwAoOTwP13rF5IvfmNOID1w8mYcGS2FeJb1B+vyUCeLG
Vz5i4G87gXawaNJmq5/sy9j0Z/C++on4W77JjETS33B8AFeHI7JAIMtjRxq/f/JO
dz1cZ4jTHdoMi+ewU6RkS9APIBHZSvRhIpoI1d/g2YipW5an0ZGPTzPOvTha70N/
nAxBAOGdRm8oQ8FA3P/gzU94ZdfhbOnxrSAKSSMQsUqITcW7JfYRp2BCIp/Cgveg
lxXD2WPuHqZjMwz1zQ/9ZVXv1u5zwsVR+09kYp51nbT9nplaVtkCT4VGitml10Mj
djJyYcFO6Xh3CMKk20V7TItdKXP4nyXdd/IsjyP0Bdq/A0SJSpGRHbogcJbzv6yG
tMr5ExVQxq/7zI4KsBvL1xJm1+faQng1q516jDVzUIAf2Ck3rcwYvtXou5Podbx0
oGhPDkd+4hm22yshEyaSQE0zvhaYeshuzEBFcR0ENGePJUZpc97Sc6ewQJpH6RTh
hJqkEk0ldhGVYkelgrX9DWVWrnQyxUkqs4racFw4O++iGqDKkZ3TV40YW1zAwzcb
4B1QkrIRhquurrQx6SiAo9o+Z0ZRqwyXARFa6yUr/H/6tuGhMWzrzvsTFAEcm4v4
th3n7TNUE2q8zOwjSIEzewtS7ZkU3xfYiwgeKtD3nKLwL7IEhRudeNDrEvjScUx3
pmmppbdPuzE5ZmcuwS3sPRjDobiYIFy4z4LP9Ho3F4/xLF6PZVogbh2UD8tiSk8S
KLgxygHRkDWKZGK7Q29s/4g7tuwbEGKKNIJq37d61jZXywTWWDSDjfq0FOFcCifY
5S41Y1SswrZ/dsRNvcAyim8ZLp8P4UvJNm02/0FqDDD99J+zQ7pT5ad9TjQ7ZHDr
sduu97mjOfzKP1GjT3XZFTvJ2FnT+aRoFrk8HGkwdNtGWz9HDr9lQQH7gort1QQu
wgJHSBaDGnJ85mKjnRxVNICsM1jWwALzePDGYcbZPACXuZ6HTsa9dhzHxpKfW13a
vPjluFmApgId8XS6kHUX7QqRqxLzClCzqDiBlrMTB4zSJvzxwuHv+QlhSlZXKVqL
zr3CkxLwsBnwnExl7nULM8fAIvZdwR4kiZFT7l3DWyvQYjn4O2So+MpJSGZ/ooJy
txolCJKFfmCywEEWIb7WM1DSzow2Y75Zd2WkPs39JIlc+8VNMFuo2ykm5caDYja5
6XqCKQJmqNydwQnL+2Ykc2R4fzCPq2xYUYYxtrbzTy01ymqJrrvZNSIvf+Qa77w3
OH4hJknXK2mTVMirGCnKpvnEaBr6+cxSFA5kOykT25VjSNMQWn9U8iLK85Cg8eT2
SCODibUE3OYfjciCbm9JYj75KwWMM49STh/lEPmoPrZzsl0Tq8vCLDxxRrcazOsy
VTzTElySNw8y/9z+cQgQsdwuQ+DdAeFdLbDpMh+K4qt+N3uO/OVWO37OfMnXK3su
kYrd5ADtgg6uE3Hq1DITeOBdcczTzn9c/iF2EOl7oq1vey3VU/cH1s47tkcU+XDm
J5QMBle/g1Jci3RPqSQjg6Kk+n8G2lUT3peYRDkiepRvQPZw+vGYVQGzC1k7Clnm
viBh4rqec8fOL5pvT0wNJGCtEwUqmG7yqh3ckidCofo7ZLShtGwL6WR4PTuYzKsi
1D5BWuLeZoShlYwo9iXTo15/HcJsElXhKsxEoZZ1i7+Xw3vemvU9zovhSv0H4YIn
lPQiEn+x/iwiYEawpvAbb8jFUVkTwyUwjK2bHgV7LrT+WF9HRZsibosQVE76UT36
WAK5XWzgE78SkjZGQ/PG20d+Re7HCVh6FW7q69+yLHvN770+7DypVSRqTA8uU09R
uG6wdRv6ri31ltoogwLy/W4d61dRoTubTKR0i4Pu3+260iHi59tBjH13vtI3yVvG
fdiSMa56UCEEBi+qBjWgcdADtUmc4dlR5DpYgsrQZxIFiULHZm0K0jYBf54y8P94
8/ZSs/OCnZS4gmJsj0+AoBnMGteynuiW7z5UpC95mReRGj/x54KxldtGqXMHpool
E/tuD1ChYzVZIRZY5Zg0LziZICtKlW3SPTMdjYLH+khkEeE+VmKjUyLBTUTdwrzU
v+PLj3T+GxmjFXX551ch9sJpPxBP8u94v8t6chkIEm+M1Iy2FN2n4g8iLmnIJqhJ
LHWMJ8g1LxXfydjyHsYrI1bqde14xrxJ5CEzpa/Z1OCccSNA7Sc1Tsj/9hu9J21S
X4zJmWy/n+v/HvqXnArfSt9xX5k2/mNghrblASGZNeKvWLTI3GHvSHNnYghO4Qpz
tHA7T2dhh7Exp5VgLyj8uq1MNJtrO2SsvlUf+AowzM+80L/g83TJ3LmRYglQE3Vx
Oz9r0+GgvovRTsPR1+a0GX1WHCdWNal1Bgkgkgdb/Hqb7kJW4euTIt9oljPHlgpM
BATNTknq6hwYzIZ12To/LUdbeAyuEBEQ/zePFyyKIOd5xM5qfJRiH9/lixiV7ci7
7tj64SM8fxGOHUiwVmunacG/B176Lqg0K0N5oXrbt7HAYr5CZsph6D7GFc5pWurj
+4yDcJUT3n1r/eD1Z4w96r8sZfMDcOjR3L4XfsruM0yuL4eXwakFZfQuJJuk0Q0q
F7gyo+YEhgTc0JsoLhL15+isJ89uHYeUDF5c6bTxD/ylssfuV61SIWrNu/aXXiqe
ZgnvjqkB4xMZB2AIi0ZMx7aXl1WT/bQ1SPFjC8a9iER0qHAVltmW33BHtT33og5N
C5EYzxazaeKrYAdJQFJEQm79kYtRf5BRvKJc2RWX2uys7ymE4vBwOhHt2N3wbJgT
Px1YYI8xam9VM+RWPunGwo6oIfxVugy/3FrcmLN4vSVG2Z5Gd4TnbeuADKNkiDkL
wjTQRvJ5plISjm35NN52o4NQe7IdR+nXnyQXqix4YER9iKnm+8Dbfb9PTFVhX8my
rhVeud4dQ2cltdQeD4NaD9Ay+1d6tHuws6Q9g8P33U02XA8G5wTCwG2lWDu19oK8
FjbUTqqmlxj7HgEpAF0ImEQxDno6oASXsOaCLgJIWXVJY8Slc+NC25/PQofSR1Ek
cKCn5HNkahLOenIsELUs3oH810WCtV5X4ZxavAq2U+78spynlxqMOOyvc9zICPME
dn7CiuZUoPfDIg+uGDr7GDbDxhZfOmbjuuEKpZ3i1czXWa8Uf77kTJdUx4wJnt1+
ST62H78LBbaaAVhuXybKQAGRAuX5Db8SLOY3jbMH3EDJ4bB4l7TJ94wfsvjqyzfR
87g2DcqpguZowru4pHGBfnmdtP+q8mI0/5gauGBsPZpBE6cbMbMQLF/Wm/x/HTNK
waiaj8h6BsjQvxbyhW1N2OF4O6q/VH+Wn17rF+W2oO7bGlT/RoJBbwAEJw3t3X4U
hH1daY+/WAKykzqaGLX0n2WuOLD7NXDNUnMWv7qPw5JvL0CjlFfMqMJfv46fKibu
itqmZ0RLgBhA1cpnCT4gg0HjNnvNggIqEkPoKp8OwOocKWiBuSJA4iEFasnLuVox
BGj5u7zgUIS8P8PS437oURG9K+UVWgiwD67MnTKV1bs3a/hK6MlaZEeK9uNf8yPK
GUp+VDSwAE+zxgXBL9HTnzY717/fPpMtGz/HrM3tRnbjvYJZ5ff/bGWkoQeS83xg
KrRLUG81Yu5P5DxXyYdvOsTIYNaFD2evDXIdp/89Lbwz+mSkL7c+c1K4ZACRZl8W
xiwYk1erNNfiaBk8iYAtKMET7C1N+G4hk940xPrWxKsZ9oBnAuGLGwidKH9QctI1
m3CVCTkCombyojdjMaN8yXjMivJcE1SCGXtBAx0rqEI1DGeSa1LUGXkokYZDTuM/
ipUZLv3Ftep47f+kw2A5en2jxbVhsgBAQ2MdHYg2zZHl+IMlyQ2h37IlGtIxuZKo
aHyMTAZ0EKFe3wp3n8TsJxQihjQnU8c9h28a8Tw71bN18O9KRZ9+DbI11EM6U6LK
cx0i2fUz2lJ3KVfkl1EuX0afPx4gZM9QVzjNKOrFFHl/lQbKeSHQaJUpHQc1ignu
9+zvdZA9/fP959z4/cM1O4J8oP0Txb6DOJkR4SHkLR91P6G4b6K7hgsyBzl3dilB
DmPfzwkZAwZzidDAFJTSUWF/Xz6OuAiHRiVJ80mIDmL/zEDcOLHqsb0p5vJWKP+g
hElwSYiVebupfjUSZGkuwldISaGArdbDs92jRGe4zwcDXY+ID6SLqbBzgwhmNOZg
C40U731+DAG8n2OeFMVK/opcAtx3DJUhX+s4QPLFwZ/I6BoYTjikKy7ZTkGqcNak
NGFPKNzbr/qYGo3o14e9BmB5bc1sf4aXbYPwIw2mj4JzNpMHytrNAiZS1iiwFRa/
CE/6ymnRxD/NfOFXnBqZzWErHSnwJYjccrhWMW1o7Z3GZtJk/LMI480LEooHmAtX
PtX2m9rmLjM26Foc6ln7m0PXxFC0hwl33JPbXFyrVHp27B4u91oeqe3q2BcuGckc
MFlXAhMDW1btCCwqTwVzQmoPZKxgEvewhFrp26SmYFII4lvJk/m4hR756/VItoRQ
BFRRdiMoTbA2mfrbPPLjK2sQ4Qxb/dh+FGqdW4Vus5LPALTLFklOoLyBO4+v+J3n
iXE1WuAI2ZsEMTaOckwmWAVLfveaP20jRKD+UgFLLbtlSWwqAjLhnpUJwBkQ3S8F
oQdbxj7CYkZ56vFQXCRAz5voiEng1wokURcI1fSkoWpQ2EUcKZML6EHl4bMfOuKI
Jm9xI4zg8hj2qFBXX6vh1S2IXLQ62XkjrwGvmsN8OKXDnE5jbQCfRS5OkXLYhtWV
qIF9IcRZqoXtf6O5XTsdhGJjl8QDea/axTIvmUEkQTZkGUY5ggOHJcYsddKghJoQ
Vhy0WvToi5Pi1SUiE4ITkiFYc2Uk8w+NN8/WWi/DThCTs6OPwJtoaQHwZMaM5DHb
MYS3dzHiwgfvCtTg8Zs8nXTOPKv4gGIQm6kgHyMSlRHXDdYkhnmpYT1AQnOXCUlH
8sQfz17U28RXBaASxRznPvKy3FEcjtrtfL2oGacAEW2PbpoLueDQ560R+ZXEFl2f
8A9yov6WgpqGFzZy068g+1ide71FP4nfsb9vRymVuRfgeayMTFV+/2k1+1zCIbg9
HU9V6i6eoYbtemzJpYjqLBX+ns/th+DIKgB1i7jXGg0ctUMfHg+FkOLSIfc2NOnN
jKzQEY8SUVXgTmnmu7ijadYaWd7Wknw8fxZxWQDsnFA/G5apOosm7qJgmVkMmat8
Pk6U/VzaYobS9YrvTrdiYtiw4gCYSO2B09xCDxb5xJJkTfRTN2zmjcPhHWcjYZso
+3dM+AxXSKZM3GyF1Qos/04VK1AR6Xrc36Q2KSVvLg2vA7hhX57d5eusB/GsbQpx
OzF1qF5plss++CAX2r0MFQCv8gaUErpuaAjhXIYOqBV6HyKH27iOWgjczceeWaRb
Qi0WMGgdB0Il2b7NzvYmTC54Rg0qEsiY1pxFjk5i9zmBc6apeKg8Ty5minV19vhZ
KLlap1RR655WXhSpmix3zvCgPs0JxAUvpmQH1CvwGZx571Q1juJPXvMqxyrytwzX
kCt73pqzIceJDJbsVc6wTAFX9FlkjCZnswjk17qA0NxJZHc7+LX9Ua3Z7ktyy6qG
Hl11I9GA0/eWYpQ2K2GiBSVSuOXa6+fc4LyFf9VkDXb02Mip7qfxxPp7jzLAFsvO
p7vtC2SBL4Bl73yQd5QRQbN2jwOVoBPFTcqXNZYbNaqDJClqiRwWBTjuFBkBumlA
7j0YcstljQa8FA8PhUD7JxUrwtlRI3D5pVv23BfUYX2F8ICjfMaL9GD1c8Pjo8hR
gkcEPxriEMvRCfTlzq9rcgZKsoU0hjIzZZ3MnwEjcoUKBO5ng2h5Yu9EXdI2TcCH
NaHkQdD2C2+85rUMAlo2MMm00yMf0zS0uD1z3zy9QaUskFfIvqgsAvLhea17ruzx
29Gg0/l6p0i4yKNASPLpVAue6HQwoLuPqAGEFVj/phn2wLS4r4bkPWzBSa4eGDFR
NBvu134S8rwOXxTAcUeQOsKbRoCA5M5tT6vPN3hfR/v8Ejw3cD4RsafSnu4iDZra
vBbFAjSgb/0zuuVAK4gKelk1JSMygwymtxdufe8IJXHpA+4bH3q6INiFbmVnb86S
dr1jgEyYmZEzK35CoQi1XFd/+5vhYk/zft5X8UJXdNhggphDtaBC6Yf7zYljM2Wi
44nSoyNFk+zoUX5BYSbn9U+HHF6er6tdAnEhbHjkz0G5HgFgJqGZGcKGyaQoUYlZ
HAzOc0Xarb211iIZTVn4zk9LOJ9WZ7h24pvIX7XF42WQdnC9Z6Gal5D+/ANRygVF
wY0WjGIFCm2su4WeYK3GfcQMGXb58g3tHYXeT//dEJDACdBGyPCvZcltncld70xP
OlX2jH423tpKH0X/M5UGwumo5YXmrq/kuKgnhUjnBLcs4tJLCPYveLLwvaZmd8m3
GSISYG7SY3dquVkg2mWSwVsLNpVpV4YXW/aQbBFfqsjGX0brRZzS2H/78h2EUTmX
QRBLSvcwohyH1KaumSsK/UyjZfcq+7Ma54nq/WgkfPKF4UeSYMWgUZGO3j3SRl9U
JFH3VDibpqhfN3RDR+CmhCCNKcVgGKtktkRao2jlPS4k9UWH+XEW6AYQ3xwL6ocV
zy+FDNxBcjyMJepk8sjYYTY7asXOnsX6zJSYWIJjWY25pCS+jBPp8zC4SY031Pmn
EIAEiPbWj7IXds9d4NyiX/8wScB3pCP7Z++wJUc00bH29nMYoU52RCtrAxYO8azv
Tsu8eXpxhvJvYSjVJJ1vfCB3Zwm7haTwAeOH4011BDtjaG5AF3yLFptwb/hZQmkB
q0CMztHDB7nkWiVKN8Wqu2UfD4g1/tGpK5Mq24/5llFkt95rFr87BNQnFzGoG6uP
6g2kfFPTpcRVfk9PMBLtFZgcx8t0Utgw8BIhNbm0FrJaYDjqQaU5d0ycbH0upJvh
HZDJtPm+aZo5vNvvHnmBs+rVdWF3QYC1cXKa4Om2rHRaPdenKngBpOCM3c0x8Le6
W8DifNnv+OMmUYa0iEF4BzeqzbMoh5E5uXU+yVFvkMZPkVGgACeQgDadL5SlV54n
S/md1pPa6UJwx5uxI66wMX3EZCz5TGNtMl3zjepZ9saaMuEmB2DOTntEHH1a87Bt
10AI9Fv/PMWBcOSQrc+wt2s1PrsIcviEDZ9O8PN2rSTW3yTokfZyqPBi55T9HsqQ
+G9+F2HKg3Jaz/sn5QofbEbci/MvmyVey15d2Bh4QbrGrKrxudwL/ovf13cY8byL
8cseUl2qk8YqGqn8fiyhhV+4KswLxXIVuNp8I2TCO2d5Q1NUzaKvJMCbTxoZtFjt
1Teg8LLwZirbiamexgOXQnd8g23A8bPTiuWm40VaIN3+H8K+7POEGUkJf3Fvg+LZ
uSX8qkamufh7AsM2zX2z0c87z0pmgJz9HBkcQKwIJPJ25Ow3Fo2h66B+NZM8jAhW
OFhGM02mc4glGBa7ZyXmvo1XH2nVWR2WoclQtfGDfFfqRHFAVtnMUGSAopa+DIQ1
chfEs+dVF6BYTfvqIgfB+yvtHOnPZ2CJCsv50M2lP0T5PLIuc4bYAXgcDyTxN/u4
ANqJT1j0ZX/C+OItBEUjh0+ptxpQKFCULCuyo4yKiUdKcC65qQuJ9JDGINZAwa/1
cM8Ct7kj71lu/P1iOtojGchCtDbTDUTfs0hbMrs1dC68Y+42ciTix4IDUg9aVQR4
tRYRLuMWbcbPft0xWXHg5nWug5JPMH9L4IVYv6xHuOl3yg7Zkx532cJf1VgtNh3T
3gATP/wSrvzREoV93bLRrMUrU1kh39JgXMz07x70cNsAicAyS4auVF7JwfH/8xAm
MF73tGWFRG9N52JtFsOb4diIeXz3z3vDGnPe7gtl7867POY+eMk0akHozxfdSn9m
IxVALsyF+xyKYMVsAHGoZzeY1EQw33fvUQFb81ibVshcVbytSc3rhQYDsLSe60Tx
m1zYepv1letpAITVxB766drUZlH0RoOTBcohgOOkOYXZknGt/We3l5ujF6eiorX6
a5HdVwbURpk3B/EJWakzYKtT1kU3yfj7s2fVy3SHDZTWX1YSDlV8o9Te6kv++g2H
9un+fv0gR7oa4Vwe1qkbt4QsF/aPlRlgT8BlXn58bPUek9j5WsU53FQ5PSYEyF7Q
nhv+mTwGsZ61ilYA4O/HcUHiVJmFzg6yzmJKqnroQIlDgcEgEzUI0hEwZy6h9Wnc
mv6I7zR3zyujmkzqIBS6pdJCSKxjoaXs05qfUHBEUo2Aj2Utl1dvhyebwN9moTtK
e+O/yV2swZZKqXytDUSXeC6SyynmNKuKGLXVGUwbZOw+EvqrhNPqrcGPMQBfxsEw
hyIjxzlUuSziuq4DzOTs6PELDiLlKQcRwLkMx5QOlXZg/bS4xZuVWZ+aUYEPghjf
B4YaYAVg5Cu0U5IqlXctZqCcPC1qAOlkNZ8A9Ug7byvclPlUMXz9vDAckgVd9U/l
P26JQFIcLOCosr1pVqNevDvomTZD96t5oeZqL1Jwz2Zz0mBVx6o/QCFUuOjt5ARB
HJ5t1pvQhfTb2xGmLmHngEM3WKEknX2FE8sZPQlfpuzACr9qcHQwkXXGtetCyyTZ
NBXcrIuLS+kcdSjmAj0/HqdOXqFyJInv1A+7+xjdB3wiWjpZf/AIdYRQ43k6vsYZ
4rqEaWPokQ5B70rXW0bH5W1wc/JJmXLVXjvle/c+hW/mXKzaWA+zTGMrM9JlJxj1
BFgQhfiYB5NhPqlhWJZU+wSFheZ4ZUdZvbZxB0xuARfb9lhabkosISru4+oGzFH9
5YNJlENmSE7DGO6R1ee0P3j2poc6xngHU2lYeYq12lN7JMpwHfTrD0iQ0tQ9tDsS
ZTk/NguiZ6wubfW1gUTK+TddhvP8xav8NF2ifMBaLIi/R0LDNfUKRQBncKHumSnI
WUzrBL9nJQHbJ0HHSbOb/8k6XyLpBTpJvd2LUFMNh9qutKLA05r3Ofk710TMDgvt
cs2QXwTy28XHTq7CnhnkwQhNbi+8WeCE/ammJPOJzrR4O4pOto0ooD/YODBLnyhX
V9+zGCRS7Jz3mDf6+ZWdH1IKssgtTuSjPbaHaJTRgnwMdrmXdW8fmTSU681fOIOu
SN42FPm+F+be1EQL0gbl/4IkTi3cRs0Tiy9sIi/Nl7Kpx1djTgegZZ0QkgT7oxzw
twhj4sOz0lEmLECCMSyJVinPxBOv61pYfUMzeOrXFtYITyGP9YSUq6SCYDJH3OSZ
k0rqjUfrUjmCjDf2moeroflqaJDKO0G1oLRrjgLeZ7UcfRp5vNj6cB4Z9g9t5gMp
8c6Urb6Q5X7UzIpCO+N4O9KYxKEke3MKC5tAsKa2geUr3WyyiuA3Ah6JbSAqJg++
gm4wQxMqM6uMWhHieaJH6W7YYm6RCtP81w8XeSlTfshbrH8h+UiI4dyYPRtWEn2h
Yb7pOJKg5BlTmwGD2psZuN/gsgBoqteVfAbOmD3O/E+McZD4b2eluBlHbwfixiP+
aTkDhBPwbhvc+49Ug1/10ZhvgCNMcnOqwxWu9PNZCPVr4ON/IvcK0DXczCUVslUT
1sY8AtoEvNwjO3sZQwHrOaDQGp94OR/8iW9nhJR3drTLaSO3aW6jn1UADwA8/1q9
YwncUbbEnc8z1PrgAczcqzRBS/9IcAWdprrIvSBnPambECzLNwevROSmp/icxWLw
1o+9lXhVEgrS/CFPwMyIlC4TxDXoKiurFx0HKyqQWpQLuI3rQmSuh5IUUZpUbavM
MLHXc5ay7OCu5gVYf9fY8KuUzyF5ShiVAsvskCsYwcRG4E4uuZOHWvZ1rQFqDKZs
jmBBqJIy8MUtOncCbdeH2nTE1nIsDAyiLpr0ANbGFW9JRQfBouBknKaP7/eUDeCL
XVfO96UEi9/OViORe+yyICV2INoG09MvR1Tt6Lrw1vZORgvjx4vkmNjG4Vh3EBPR
4fN0Mzk7xaIx9a78as/7ZKJzD8GEkxcg2yh11MpYXG/4wZ5zNVP/yLvaFEX9SwDx
qb4ZvKXzjI34OQ+ZOlYgHvJ1FNagOgpIxoIkcdvU4Xyr1eDRswHE4o/BKA+AzSFX
hdCH8tExX4W6S75I9HXxysGWdi5Fu1+f/MwO0eOz4C7+dAVkqV0h3DO39PHQuRmH
7MoLpkohiTy2wk350dlMcHuEp3l4p15gsNe08FVv/890HawZ9htxs+pF8pOYMlIC
Ob2ycN8FJsoj+x6QvVVkxRYNxSrFGkvJCQJTmQDY7NaUif2KBUFxvdsD3IOXOzNL
ikxGanBQmj303dNRqH8DC4vpMyt0Hthfgf3930Zb128y+tA/U8H4q+ruRrsIQayT
ijPy7by5kgTNrt1TAbxZON4ShpmbI38kv7KERxGu/fDv2wrb5BeYqFPyYqGvYG2y
n3qB01rlh3bJ5//OBOwHVviM6ex5ZMwd3UpTbYyr3bBoXfOKLR4moFUjs5IRnus6
5XqtcWtrbjah3GRxOX2oHx7PavzQkKxnQ3XpPPWpLkrLmLX1yLt5nPGUXWtJatuT
MUIMKGbWjSqeXFQVd3nTkrUkqJEqI/aiI8J3XIM6ZyqF3h+HxKa1fceQlfoe36/0
YVG/jx5aGL03JR1fepVEiSw9n6RdPVz6j77QxpkTiakHtqR+VxhKqScIvTWDwzbR
HJ1LT5GOXf2Poh5Eq4Y31GiLvmGlbKjxqoTfM7m03oglxHPwhqWNY0w5dBtiPYma
5kZNhfQpSp6HEihFLpqvCQa6hbeR2IvgnrcjNggZb60YsXaHzWf8UH9/OwYBcU8c
a/rYcUCSXxYxsf5ON2l9y3qyfru9xC7xLySVegTDK0lhnoFB/Ej8mibPyko4gKa+
s5EDWceycBISCpfch9D/mBFGnZwPLFlfPuVMhbqWTYig94GFL49hToFqegO9u4NK
C/HQBbHdfobGkRe/ijvwHbmZfXID5nVGp6J9SodnUAqzcaAE48prnt29iWJ33m2A
SkxJPoAypAZ/x9dLqX0FCLlvtRmC0/GQ1vrsAunSZjfzpHCPjiIWZImt8fCEfOHA
+GQ41Cs58TzrVjUa1clgJTjSYxh5LRzdsZcOa2Y0IVJdZprzSTyLOeO0i/PcTJrH
pY9/+6/ORhvXOGLE/NM8MAObkZkJPbGMqdCXGJs4Z3s+cIXSSkprYtKdTnux/Fja
U6exXjMUwZqH1e+lYfNY/zOp3ebUDZhk5u/drzdbgBScDhTzib0/DbybW9Mzo4Yg
+Unxyb7m3Y1wv4uAYSI6/isJaApdDdEuTvtCBegfnU2IAvilOAFf8yo16UZeCY+E
HZz0aoQeijTMUm12TR+xsICTaV6jqB6jHQ+0muc3TfwdK1DlfC9Hih4LPeKbrNNt
lBXlfC+0XSr3AtIvwlRyyjbM3rOX63ZA8rYjErjyrfu/DAC/vmvM1VKGd6kTJFAf
ZZTYJqevwBhLFT4GVVm6LY9N1YcMwH49yQ2XAiJACozYMsUexCCHk8QuPpExxDhe
AahpDOHFyofo2PeiuCVHUPxB+I3CcDnImlLTWzjC6vQ1nTPc6Nj/Qpb/gBDpsjUT
2aK81V9mc/+xHFsNxMeG3VzhEKbG1pwZV6Pg9Y8u18bMgXu+sdqgBnVP3oXjfq7T
ntWHPljTEt5fqgVkhcMH9SrOU6/DEVLDcmO//wHnDnFgHwLjaloI4L0MP7XbuCkX
68dF01QQedYCX8SBY8etji4yQHrhyWlIC1JDfrBOc0sb5zknu53QxjaK4CXqZB4M
QVAQVPncNXsa2Cmk2xhU4XnuKCuvLVWs3smH4QB/94Gdg9ELF1kFpt39zWHLGYDN
0xS4M1OSri6moYnBYqF4LHB+m6r/R8kUmSfdxAte7TqLWAQMFMTQ5qGQO48OhUM1
KZ8XVAxzhrKtyC0exwJV9HxvBYophjaoGG9enIWQ0iYXR9d/9CuT0L4AryPK8Krm
UufzAuEq3GEdYOngM70OyfvWN4H/heBvP+khHqR1wd4TSWaT8qhwFgtEq/V+Mm7p
EclxWYKmDFo1DffHb9OB151GXO9lQG3KtdzEcJLYZ+sX6cTtJMK2j1k2DRAD55aM
fk1Mmh/RQ7xZUqPKJrn2a7Wuo1PBxICinRkPW89bTydhx0uOIfZbnIrFc41TODrd
rnVwsRwDhu4uve1rzAulOrqW/tDdid2wQeuARgsXGfwdn7QCbvK7eTEBESzJxteF
xM6tnH7Umk3cYz8wz9uGzp0SNr1WmqKaPYa2gg6e+33h6PI0TX74XcWfqThv+atV
ZV+uly8p7O6VAaVuVCss5/UMMUoDx5H+i/3hJPiEnQsYJx5DYwnMOFHMDvF+VQ17
ZrvCnXuHx8DJ2cNrn0d0q2ildp390tUwrvjY9gJFrx8D0azvrCWIhdKEU0nktM4f
A15f7T27Dk7RICvKMNTxugGni95af4AFOz/3OxLvkcbqBV2Br8o8FrI9UAzqLxDq
jHI4kd92VYKUgTl0q46s1vSxsQftvETpuVcqMsFyouPl8WCEbskX2AMGIr9T7Llf
une9Ycm2ZfQrScknx0fYwG1xcv0SZRGkI4EZTTwUL5WU1gVGs1p+UgJSmH/LwjjR
fYkaLtpeMQ6KXADtVvq0foDpcFP4HOe0JX8y3OvlRY5LL9G8uya4eaXX+wGJfyT7
YUAThqt89Rv9cOYPmUeFTeRbSm7OQvUwfr0r2TA8wU/QIKC7F5bl7Nqae42JvtIV
iOafXxSnowUV4qXpEVY6ShudkC4b8sC2hvRQopdsGrrqkXdC+qTwLpFY/J3NN0mQ
74/HvQ8ViHXboM5QiNDEMc/5s/5OHIoBhNv5ME6kHyX1foR9SlwQcrZeecaCIdwW
QCHW+iPDzxx5jbVGR6jfdEoL67odLN48ikIrm8ZmqXpDI6N9GTkvtj8i4aWtn0j8
wCYGkYw2uQkhPlpq7Z4NtnuF4QDF7uY6bTzOfnWjn7CFHmHT7EbzihlJK6xGSrAU
aTluGejvdKMB24Sksh/Umn0rpCyBrxXMO+/5RGtqvcNswRpPlZ4VRKL0gBjehdf3
Mfa1IhZrj399GlFmIro2jedz5isB0J1F832E3cTmvY/Wtk8ubbzBVXHXZztcqjFD
x8SbaCpv1O7yFla1oLxDImmoYCHduzjOlEIa2Ac+LKPPeFYvJjvljNZyq/3VVg/O
jheLf+a6klGOVEDa77nxB+RqEZ1i+79K5zcJ+/QXcw04zPsHfuMROSJcsYjrcxuM
rYjIsbmh6yMVDkNT6PqAievwRX4kq/FtoLODN+L00I4Jg8MODypvc7SwoWCumdXR
HUilQS07TGKfM7/Tw8TzgPrZMAxYlpD+Yn4AaMKhp1jJxE29sEqPPH4QpCzS8LlY
8XkOGB+LH7QdG962IA5LXmf2+sqhQpNAXxiIQUmTWn6ZF/NHzdZ6g5erCS8t47uP
S50HUzlzrbEld9nQuMp/MOO/c6VWRthTiVrTJcbKw6THABT2XhPmRF9vDN1bUjS3
nbOvPapobrDk8pigl2cjtm5r6A1oQL2VYc0IPXUqIuzMwmTBupABrojmUMwl1cLx
l6uQ/JCqPnMXbkAU8DFXsgiQ46tcwJ4sPNKT+fysDmef/yHmAcRyShBJQ8ZEQpI6
TYcqAzxLhx+qx+uRMSOY8OVH2uYjb62UaekHAIBwRVbsqB3pchM19lpip1twnWPl
+cpjaUSgU0Zq/Gy0ZAUNmxqqUao7jvAGkxB44eSrjs1D2lDkzVaUgffzM0GD00gL
VlFCVCFR3zsKzy27jN5jc3MpVvOBuEMoQoHEj8y3P1s8aTPACTsTx/ee+nzRB3El
c3C4pIf5zgbNB7wyN/rs7PrsEzh1dVJbh5oIKKsMyUtfNSfAUp6MUvcW3E2AzO8t
SQkcOgV7XAHg9xlMM5bJCcTt7+IPq540jaq0gJStq7ywtGS+d/vxQ3EYMQ6mLtR8
nNpCtObeoiSiSwWzm9BGVeFMXxtLPi1PqZo+K38+f/53oT/0o3EfUZJwW5nghoB7
r26fYiU/B1RtTbrVyr0oqg1wh+GAJwCrjMrqgznxdPl1Q9e94HjE0fW7z5CIvb2W
RRDrOPTHusMd2qGKNcQLSp2epV/O37f4MVCIx/tbNupkStV5oim+4fCyCh7x5yuA
WQZ9dMIcqjlFDm/B4c0aV9WnZYd60XO76mKFn/NyCSH1Ln9OGs0u/RX/FKZiFIjw
j5eq8JEsv+PRHmqzqfjDbtkO7cJS/2JevsFFMX6bXXWZsMRYNFbA2+OsZYAV7CMr
d7+6F6dav0gK6w4QXC+wRfkIvUxjopj+D7L+6X6ex7xdYkzdCtjLUidSh5x4X413
f2rOV6/JFIjeGKO16Zxzk4HMYb+zb4x1Ot67G9XuPnAYj5V4bSGCaaaTblP6ZxOL
hCNx5HcVw9Lv5acwPnSqsP6y2Zv+pqk8B6tblbKSfcfNdKKnP8FSzGVk2fkLbabC
MOuFb91lSWanqSfGW9v+6IuvRAQqffbgy0oImHFYlmvlDoKJhzDKflDcmHRtQa9K
B2guT/nL0hbRwOUL2sLlAva/O0BuYuUXP0qhbRXneDeU4kLuo6yunXm1pPEqqZv6
s5mT0Hp8KMv6pvhaNBdYwoJSEI5goIBn0N9ht1H2d+DieRLpsj+U7WncasgjhFrU
ui7ABN0L8VKTJAHDi5X/g4oz8vJmY5idRkr/XtY/pRU2N5bYf9S+ueg1Aiihbr0D
2JMKLUBJ5hTVcANIbRZU9PyRD8b9aAm0KpEUeB62hH7DbbHw41Xb86Ua/tpNU8GR
aL1V5NJgbuLIL00zDEygfqQF7NP6J8kDzk1LFCsHaD98OpG/coJlqToIuaXZGgud
3hQFDIVZVUMIJ1LfiawT9t+0ZbpqK4K9C7P3OBuhDqFWmoVrEPt6VxxcENkH3wm0
34vTYJqxORCXuX4ED0VSWR3HZrkcwQ/ZXH2eLwY3+LvWZfSx989xJtZjaDI0YTC7
gcpq38I9HS0MBUwcXN2pw7JFMQWLnBEyftTVOhEqbf+x9qMHyqhw2dZJ0VQOnqHk
Wj1GiO36qpNCjjiooQ7MyzmqE1cF8SEaRVwk/An+rXVymlExzWf4bcha6vNA+cGh
9wsTN6v9+Vio7njIB+PcnmNG9T5bhAfKP8EIt2Eds0qeiDB1Pn+hoJoFtdHNntQp
fCJzxrrj08f7yAvByf4mA7mSX9Iv8Rui9oQGoRiMyOd11omIE3g0SAxG4k01n7Rc
4JkGooMK6gk7B2rXqIxU7QM1bXrnS90+YdQlTEyCoBMWmefTGQjIF3ZJK58mw3UV
IqRPHEEFQKT+gcFYVq8iniw1vQxuoQmsXg005OLKoxNpBgr4tLFEPlG+YggYRPr7
aYtF4GgVmLCYpuGyWZlWbTcfXhZyCvlENxtREzybQS7UFMNHKz9nuXDZAT+4YnPP
re0cVo5kDO3pFre0pgxRMxx1JImexTb3qVSE7RJq+TAzzxV6XfF8+UMa76F8LJAm
KJKco5y0JNKqf4y79V2Tacp+7TTwfR9n5BVrKcrVzlZOSxtEtaiyj0HQe/K2OCXk
qOUK0F0iSpVdbItzKcUop7ThY2es/fhWFFnKqfEmddhwvXeX16rFx0PjVl0MwAC7
9SZQXvFVSOnhgeBy1StJlOlVtSYeStjCgSe3e//ms6Horxbv7o2caWQ1n3/OG+x8
KSOU/5rWVCNCry9P9T6dCP+IXXxf3ZIrXkVhcsW106+SC18DcRBkbzzcS2RVXIl/
N6aTfVbyhutmrKTDTvG7BgLQbG/v6RGjOGcFJHOWpOgCiO7Ry519J8l8BCMGtwq7
/XG05IdZLVO/lWBqjGVGVjcSzjQsJgotVmtqK5/5kNWYx8WhD6eV376x3my9HOro
lN8+oyEIZv9uyT5dlHHSeOJ5GDxv5YPnd3G97zA3UdocJDstwMN5CopQgc10Nz4I
NHyMogCbWT9aZRLg7NgSpNN770oStNMAGfV+ZsdZuH40rhDh0hMq4oYyONcQgLS9
hVaTiFCx5nI+eeuK3JuMD9bZ8riKZxVT0VasCGBAgQtrb6YXA97KO82g4vY56XBW
QYjFi4NazMI7Ip0qT1IOgK3p3Ls3GVfm4WGZjg1z9HCeZiIaahjKzTJWjSWIEPpd
Uf4OwWPgsa0K5gLH1Z1yflXWaSC5p2+sxYy3PNg0xKxF6MB9Kh9TwtKIuKhIc3Fv
NWe4qJin8VUjd1zgD4HM2KEV0AHbktw+AsVWQoMwmFQ06VlUk+ls3BMN5HW1WXgl
PaYqBAmB44twLPx5GQIXOvAgc/X2vmIgoWO4/IFuhhM9KijDNlSVBpbN5zCheSku
I8pXG5NiqP2Z2oExN6fcxpEj1RRsSsbkA6F7voGOQcrlYU25mCrEzMhPzgqqzuqU
tFthIC8ajos3DHAvjYVgJIbV2xqI4HQ2gfVDXHed2uo7csZh/2jPDNWmTX/gbm8/
KXNK/V4TgKGMXlD8c+jhWDR0MYYq315g2DdbWUDN5mE6xZ4Wr1gCmxl5GCjipZQb
XpcgcnnIfKwzxdtGVydi6DWRvZc24YOC72bMtprHVk2LBGc+j75JkItylqKwnXXs
mbPvz1oEmiwfJfcj1rCtbURpDKvvhcMshBVuYysxXPoHzAwt5oMjKnTNnqATfxRv
EqYD0AokjnaJHJ6zyh21TRd8DmgLDs8wXkEjI9HT8XmpYOTnqGCjGMCZNae5vDo8
rSvo0Xgn67U3lWe/5H/bn78Noc0vDDC9A35W2zoJE58KrTMZe9Yca47/Ou7WePq5
Qvd5Oo7Zw0eKEfJYVTA0qJbTr2xFk68i2DfX8ecPKlKZCjmheFtOrWFAUdn9Hemd
/HyExbu0icz8M7xuFSgXtWXdwrBpC/SFMcNs/ZFMhaRcFn2lGFoUhhNuOV8qarNE
ULJhdpk9G+songXtLrr5EdRd6iDqACbGYRuHwNgByFMYgdxxQTWOaJSkg0cSSlfN
axx2R50y0PaejJRm90etrX5YWIjIgVbiHWicKNEu8KfZuhJv8GnBYVuRWL05H4bm
wejTWNoVlsKciXWk+5Yw/ctsec3/NWfIsW39VuT7FwaYLvPvjAXy1YduT45dAzLb
e1Da+FY/JYSG3prYcBGaq6NCGznOjG5lVyxoPTIgoDl9MCtAD0WUbIbPzPeyHbY0
0lSheEZkysA5IK4QJd6C01DsJAj1wAb/aCg7Zxi1UdftVBf17tR5C/nmbims+aln
ZlSnZXDGWmTHvW0N3cr2iHWb4qytZlA3LhICEehjsTmM1l6xSbWskcqEuaf/zVl1
fD5maz6Zkslk336k/j+/imOSJ9epEymS2m/eCHscTddFSyG/ohJptHad2OPK0I+8
bOPGvKUDcJIG/3tbR6EFMLOYXaffIbI+4GkaS46uVD5Gz6G+kmeQ943zapRuHryw
THLiIrSPVS9K6treALtaXaryeSv65uy8g0Ti+BeVLPR/1BBjSpwEXlcMlwXsrx8X
Dev7nahKQ0T9ahY9Pk9RYR+lOtbUuPCKzKMnMBoKw2Y9QWLi6oHVw7PcpJMl0ixj
9JUbtlfz1uWv+A+YD2zuYt5MlKr5ZoWYblL5yJcQY9ZHhqBEiJjpcR0lnKpC+2zw
6urhVMAH+eDBV7oV4FCM4xWqXa1uohuRvroYTWMCNKDGswJ5ot9JmCXXyqpP6Jrs
+sw1oWtAopIBCgtI7KXZ3uRouNppJ+RGHa4CFpsYmVlIjwPtAfx2s2+vo+AaDXU9
eq3xJ7nYSMpzj07gUB+8xP6PVQRrYpbzRE9et1HA2zRVFVbNGD8LFDhjOkUfiF9p
BSknqxfnMuuuAJfEjYEc1e7M41H4qvx/jWt8AKvqmg224QBjQBDn3g8nn59h9jsI
PrzsfvPdM532pR878bsXWj5WcU/w3D9R+ZCLKGy45VV1bHaCfQXsFHfyFMH3TXTj
mlKAnG9JionO/0/GGR7X38ZYnj6uzCQ8ueVbvbxhvDAMhfyX9OB8scUKgVho4yUn
epjnFKe95qMqK2YzV8gZtKusBF3EBKBI4JljJep+xX26i54Lc6z2Of+coLARIoLX
uiDzbWcLa10ZNeuFcQ/BPbAd3ZtmqKm7/AGF8GFgiKQmW2J1udEL/WIzfBBkMTAG
wzWYIS5NOWBxRjL7v8G9CwsKCQegsbrTrjHBEdaflmsfyXdfM4TkDjbqN9IldtZR
quz3nZBpQelqoUtJrS8r6iYZ5PlVDIoW/x9iR5X13Va4GJkD8CTTbEDg+p2anQXD
Ynx18MU50sXeSmM0aKqD63aJydLtEPY2T3jW/knMhD/cDl8aomYEOFlfLU3nODaA
/rc/VeTF1CZS8jH5kZ7vzKRviSuH6tzCqnYtlQag2CtrkLWQL2Pu4C+mOas0RjwR
SEfQX+9ZHYtXNpOsDx8ePopAcChGh2zvjHaC3020q72PrptOe51ZX95puLmq7rGr
DhTvqGRVNRvU5U2mpy5D/tXC4PFpWZEgY4hcopEUkCGGN9Qn7MzXPSoWyUHsA8Yr
BAdL5Lvje8c2Kd0dr+SldlTiI+Q6zzOS6CpiSiIQJyJYTzlpsjar7uVR7yC+nC37
16fHEAWCyFp/RbYix1K0orOI21zlev3tCmC3ObteD2gdGNwAYqtfuCEfGiBFi6ch
I39V96x8UfETPLHuffvtdwSUCxx9vK37tXy7PAY7cgLpWyHxeym82cFZZBwKQD8S
eV0QiJGz5Xn06lO1qxx3DCYqbRLxFpTs5JQGrXrrsm0TFW303/laGpErz/Jeb/VT
DNKCOvZ+uVrCG0XXE0IbUOKVHUplXAMTP81KadhqkEYS3YXfNMGs3AfdvQAyPFlK
35Xm3lyna9rtLsZMvunfLY1iW3EXDEtdtjHNXHuq/h7VCKUGjMKEkkSN45ruSxe3
IfAbr3w3BgkvWtbiEIuh9t1yJtK0AsH1oqmuYFtbumXCXzGkehFU3x3rI9TCytxn
0DSuYujeTgtIpA7vxfXxBNUM4h0fmlX4IvmBHaJ1lioMyh9PxGQkS0T2POjUY4hM
/kgIogIFw4MEuZmuHjTJ7Ssys9tpnGuzdJV2aU7HO7GUUGEO88Rp9kexZfEQKCrI
Zk7Qly6N0TpIsfX9KwdL91/iAlZAuC0vDtV92ZuIVt2+Q9XtwMOC1wa0AQVmmu+n
59xEYsOfKRuD6EOqj1wszoP39E6pw2dNto7AhThz97nALW7PR5GKaZs3PHtAmESQ
TsUAILP0Kp77FLRgCe8rcwaYQ2DIfvixGk4xySlKgeYThDMHbv4k+iKQoKqZNdn2
j20VRj828Acb2CzlIcvfZOvHNf9TkT5cR0kkjIn1oX213GBA0ruRRTJ4F+dWic1J
Pv2uFEEGBeuMaNZlfZit9K0oqadXmuslHHajsZ6bysbD2saj2AvpAJvQBSUGXpwC
pMMXWPsRjdTOkRQBU9FFL9uREqCybpwNSLI5lBBxkODUfvlJgChDHm5z5l22UtpM
kbx83sMRvZcYdn834z0tJSspaeZntCxx2I+kF38J5wD2yW7/Q9zd8giLni+MwMjX
uf9LjBJ9FlBKI0yde10hWhnZmeSzCMZNVlrLj7pOF/qNC4RquOZsIiqvQaVnJPcm
cMr6tpMeetpi4S6756OG4CeQrcbi3gvplQ/5Mi+3IxBlN6e4tY8a4c/1/7aodCnG
mxzfP7MWxp6ZOelGvpasVz0lzaUL1F3QvMKxs1SUB772cRmq1n06PFf6hEcyt0mq
MvLS9eExuDpoHE9YviwUg5/xtfhwAHuTi968z2NGd2p5Lwkpd+mcGANP6aaI5zNN
YWd3/+TdjWVyM6RNmA/28moSHYzQL7pH6WHLY70PgiuSIwNqJi9m8QQFrnXDgAw3
T+DY4x+0GXM6McVokkONW+8mrCrV8GKz7zo2Cm4W3gnI+DfQ3xbfu/koubE+XeZg
waQd72DAlKcWIDoopU255Fqaq6dY50aedlDNZTugukveNncQ+B3atkizbAiCv88b
+GrBxLeaP7zo0F/mXTVIVezz7DpuJk4giQ8NZQYPZav+EhwOv5+/xjvqXoqSVtwK
Z0Wd26LI3L8eDy9rqXNpzkNlyR5PCBUj/MhcchGy3fQfbPjxhniJGs9kZU6jnOga
a6CTxxIwW8YC9ULbmhBSAh84LPzHcWhCXUhY10c3hsUQJNIN1kzIhOwHc8foVgT7
9BGfsaFJAl4XO7Js5XPEapPwsrvc84ovq0Whe2Q6aGNQRzWwCmdHTI7KRMGXxY4Y
kV0NWOVEV7S5zbQE5UyF6NvVrVvOeVXxt9o89ylHJy8Q4EGj/lSXm2rRW5r7dU4f
wjmUuipWd/0nwyFtx6f4tpO4/pWMBXK4SPrN3lI+tb/z2ZKHxUukw2V/hgodCxtN
NHY27n/NYC144pnLdZLNRzEQ06NSqYxw6JdMli2+wPATA6zUrGNfdq1UDhIhhcnC
HzuJWTq4TXCRuZ87GLblxlQ9xDNNIC4YyRkqXGR1PbbIuN9hkd6hpPEL9Su5bBjI
rY6w4/p7DLTA1w9PX88JXLk51K9fLx4e5F9e84asWw/Y054szCTwoq0UAh15ZbIT
barMYcNx7lpXpmkZxS9zUo1l5T3tKo5mF8dcxVj7wYXRAFQTMBqTvZwcWfID3obO
ERl4mOxUE8ZsWi+E4Jo9x0OSGZQQJOXYspbmEwsPS8xgPcthHNNEZ9wfQUIHw8oe
9nYrbucmyMevF/2W3B6cI3gFu/HPDDIJtJQCx1PYX7Kp4Hh+VKPnVwMCwm4WZdW7
ZAaKwAh4PZcYB5Tlc4HluiBLITyJ/Sve9RhxjFqn4dRLUi5c+GnCH32f1fpVOX6/
uMuaJ9DKY2HXlTbtr640r/qDY41Zsdn/3WGSUtJZ8qb9NhJcj+WWEOjcqGu4wyQm
ophS45XMs9f+KCTzUFWeYolOTZIfVoc1xWQSdlVsND8h0hTJNR1JgWh7JnrLS5Mg
hEUDGmysUtEj6GBxuet/ZdNokHzoi6CsCNq5v8CPl5NZZPFglOE8U9/X0B8+foDP
O9ZKtBmLE2A2gXT/H7gV442VMWRQmw0CJ36pMUALMjPX6lK7xgpN0Qqaq3OhHPp+
mBrtQkWErbLllmntg4RUq8qmKP4JFtFdIDinVU0AGJYI0bT/MndYjx6EvJS/nqd/
d1F0n6O4ZlDggc/XF9qQv4j80E4bSzjwAxsN2QhWahc2Z/DQCpmbiZEgJlzW2gYr
fBG0RbNFK2jrOla4sslBWI27TUeEDV0As8ECNEj7ox75NJwDRRuMNVEr+S01n/KY
ze80YCD4yxTPK43Zi4Nxb8BHQTBnbHOhaiLGt9FKDCZl0jf328BsyMzqsNklLwom
R8s7ti3bzPErNfrMsGclzSi7644OGrlHqy/JVLjtG43HxIV5/izHIEllLTiUNGeO
S7zTy2Dp4yTs25lvq9/zaftrs4a8Ppp5SlVy6CAsUNndhDGCEwYpoQarI4H5i1Tw
sc0thp1fbklaW+yH9UTB/6RyYAtZRLsZkVyfZfGLTkNO62fp2UHlATLzncCtdJAw
NqkGqz04Vr1D4qfY1fWZ03Jt/chP6KWtHO6kG8bq9AtET6FJVx2ZULUPnTCWrRzP
WMxMueOF7MkTDOmwmvYFiPpwgnEKxuDt052mJetgjxMq2bnI2Bpt9B6qU/ZmhcOT
LK+iy0VrULu1jz1TgWA8Ltrheaqm756SeiAruEGK8mM+8wWD01XIHPie2fiRMcl4
jyGMlDmeRbprOt1cRHhLCn+Oz14tLwDBgRKhP3aOHEAkOhF/xp8OC4BeMNrCUmX6
jFon7sAh4tqGWjt4SdvlBuiiTk4iRRC/pBnNsU5HEXNRbcg927wZttYOT7Ogp+kg
93VHjCOgNZT5l9YLZBpnydM/0matp9Mal7LpiXSe4f2zWNpKR9uuJuZvzERmxJeZ
xa3joHZiC0A6yAydiyPsBEN9odj1680oN2mJGx/hVneW4JDLoh8r9MkLFm0pNwPz
7XG8mWyoJznpbNtUPAJyUMCJpFD1lrtzFCw9WIQA6+iaE29glO6e5JiEDDX5Qmji
UnR+KYiFsCRVx5MIMmXH4FmuDHXzBFUgJkQTK97io1TQ4C+pcPxvYVoPOyS8opVC
YCsbjqxNzahGjzDMhCuESE0Hs4jdOWQzQ+qXs20F6fcJkQPtuM5HaAsvjnvNMU3N
jfci5ZzW2mA9RfY8W7eu/EUdpQJX1PdUhKgAheJJOMArejqpA1KMShGWs7zeDpiJ
37ZamBMW2v0Jt8QoH4f+pPfSXLAGLpP/CvYjP5t57afPNq/c0Vr206rG8rrR1Avm
viUkJxJJ3iGeDf00vkLFCaaPWnYXmH7X5ddQaSILmI7B5NUL/JQNZb4sSo83jdyu
XgVUz+1lvr/tNmtzkiIjh632vjWo/Ppe39iU0Tzum7mow+fkmFmXMyYLsJj/m5KL
LuLN8DUEK4YO6MYkJ/zcSRtmV6SLcHdxgEq4Ky/We2Y1hYYi0GVzsV5hLjYytHR+
ov/8lVq49XQ4ovhTKsNhD9SSTli8RYEnempUc40W9v5yswC7iDSytqBd1ntGgDke
a3A88aaBm65yvw1D7zg+AnS83TFHX4DL6pP/5TPC0RjaAchF7f3pgacOl0z/0btn
FyF3KeQuPXEDMFUd09Vxcee8p+Q5n6nTL03BakoLVMtTm0OG2FOw8FZmqVebcIMW
VDnxEGnT1VCIo/7ud4w4oDKuwgXH6tyzjDToeNWFeY7ZCrZ16Add7NITutp4sUW5
Me/vxFDFtuSlBmkhM2XuCE1nktHaAXU29BqtR7e60/PCTrCozkJLUVSBRBgwezQ/
GhSV3qz/55V8YYiqu88/cPX53q/q/TNSGMfUneRlWdWTQhCrD+SasSiLwJ7Z/ii0
qKevq7Cys1aa53KH7xaN1A0txfssa2ehqmEcAUfBhNIMRf7reaN40O8Kc9nwqJOk
tpj1m6FCAy0xbaPWxgrFiqxX0w2ohbts4mdxXvY1yIfWovCK7vm4rjChIU6yuv+t
WRFV5QoEB8viCoDJydohRdIK0aBQrX0galu+DxYymTsTb2xXH2fr//VgjILY6a1C
nWnL96uG5fHFFmstS/Xi9YMMNz/NpA4LE/pQdxj4h8LujwN6m/fcsTWmGYSeLCm9
uB6VX5INBDY/wrjK+ZeK1MsGRK3uABvUURjF8oEAi8lkFVsvnjnyqDC7PkWoKUx4
Nf5aiRgeyPks88YhOUG+WFBex6fdAYXp2YeaqZZvJpLw1AOs3F67VjKF4RhE9uJU
79k8Eg4Y1hSmsEE71cO0betBuw6r7/gpFw7fsiOr5RxKwAxVFEt/BBHECaSePcF+
fDCk5LR+9BjbodMqLaoV0JcO255oVJIbU0vXeRoi7WRij6oEPXhwM5xxLS5mGxIO
Xfrh23gchi+/RITGxugK//EmcK4j42B+nxPEcvUgI6bCFMDoOouBvuwP+4I62+JN
yr3Ft/ezOLrpBO5vJ++0okdwW4egf4VBb5nTMaI4JsAg8R2q8w0ufFBT7ZiPtfm3
c0X1EZ3lNGW+Rm2se8/J1rmd366PhfjfwGfiWTXMuqrJgwd47s5xxWR0G7qOnzJs
BlQaYTeblcj+FGPzurVtBsBfQGMT7J0+XxpwVhOV3wYwLYGRkfJVOZHONu2HhVIB
H92PjbG8ydkpAhzUYVJJK1bO/lYGhIetiTtbuodU62YOcwmD4DOkyEpbYi9IV8uH
wrU58HOEZ9hMd9VhbvshHmcg3tCASOl6Lu6TMf6Atc9edom4ad2gbcd38owm1Vty
Qn5AdFDacHExBTD8B6sFwi6kUcHedcTF0mdWEeyJv2T0xhXYzYbvXzhxssMzZxCq
Vcx9zpiDuGyjzPv7oOC05l0Fu52pK0ilPUlf1kzyzd2n3lkWqxZYzBKm/X9dZ74o
YH0b3JRrI0cAOndD0P6S45hK3GiUYYr2pGNfIgrglyMeBV4599ELYt4XpkAgnDZE
ShZDiE9cXIPjFXywb3XraBVuhwPEEf9NepcRoaWn+wGqzLuvftm2ZTNwx1C0afWc
3gW6em/RcNsVPuc2cdhE65kWPVbcIZM3eXU3V9vyUi5SXkKMUQk70Lz/uS2vArGF
iuw9JRmQXoNMXlBjsn77ireD/OZsY84ePx0lszpVB3O33Q5cnS6laxsq7m72FKMj
80cTdI8e91jtpsGV25imdfpyCN3dI0Z4Uzj76iWRSoQTOjeNR2hRXROnoiNAFcup
JCT8YJO/OwAR1cP9eDDdLStFhKcpDFgfGwPloI5mRYH/id+xXI0hHIpvsK5Ul0Wb
0u5BL8M/3czAg8xOt6FIY01jw3SCzJhpAyTlT82Ti4tV3Xy+6xHq+tRFFrMges97
jNvgyaMdiQhxx66HLPd+wry1d3yDjNBKWUFrEOM5YeipuC/kpz7NlAjAMCzpvxze
707Locijh9CJRjGgiMaOySKMwFTUl82DHPKmuf97h56/ZktNHTSE7aGgLyURyDH4
1kRYj4YAw6pEcIazfVdVjcT6ZV3Kim03KGtGxY3U80bdF+AibHjxMtg5bfEaNyue
D5zp+b4mkiil9yxey3YqBQG44zT5IsdqtM2AKoFFxnwG5LlKMCGe78iektlw7vWA
zBZLUyz9VBLd0H5XL/R32AxSlSqoQzhEYdsvf2oIUPKbV/OhYJBfDOUGynnPlaYC
fMcCme+oDX9jI8gfsnEFZoCBN1aoaDjsC9xwczER3LdVUk+81SMYbnbML1NUVFu1
lehRLl/g0Baol8cKvN6/hLbn+/Ijbjpui1f1Teh497oVZu8hhKASXDjguAnFKz3g
WyxT0vhUDe89WnC0r7QYYYRstgaGORN8q91j6Lv7GW2jlQa7Fm25A8oPuH5M5LX6
js0cOT++qFjBDjYBdgl6zw7vGyKZp2ZwS/DCZSbbo4zGngdxiQ8Qs8Bbgn7MURDL
lEombOSQx2snph4tVJZ5ypMxhCJ31Ti0D5Ke7M/iHDGs9qPWngII8Igi61kDIYxt
6PpsrV2fjM8wuHOgopcy8kDNRqIAZmtFJqP7tHeRxRTADC5COTNUG6jR9FQ/fu/r
ZrDuD3d2jDaVA7FqxFv4uJGQ51EZco0brI5w655BZ/jOIlUcicmEGKWMC4dLbYor
/prDCRAO239t6QWe/ry9BWiFD9IoeWokvJcBpfPGF0sUc3oZGiJklFqTyayG7ULz
kGc4RCfqW8gU9LjREMvRj/soKZ1D67nHQkWF0OLVJWjt3alVJAwY6tTEkwyXsAgB
klhrtDniNby3p+NhWdfOgp5yFKmt2aYFDj/N6qL2wF9ytaODrx3XV1woH9JEZBSG
04mY4uRq3LY/9HCD1RRP8YeULdkycT+FAXJg/OJOKpRH49Ljv/yte+kvP4l+6QVO
7f/LGnydHsUTNOrG4O2zUouPSv/XOOx8dpYiy32fH+EKhf6/KZwlQ1KBDHn9DO2q
CrZve9kLlsMkfQwkgQDlN0RpBRz+ISB9GCZqocflcgK0qugvpNPmmb7o6VKHXY6y
4RT097KIPyMjPaJzypgrqCSIisMwRXhEQEfu4vMMTs4ni+lyRaOxdA5dyZKvLj3d
019huI2gkNnW2Hhs0ElfyaolSgcDvfs5kPKWKIuQhMdwMN/RBagwNJEtxgfKiann
0/dF30Pja9bhbeLe+WNWG6Ka5IxHnyxzjes2xM0xqPoxk9SmFD+0i/m7h7AquizR
6T6EmN400+E0VRHoobEKUxdQP5JpdWT48HHjn1z4yxot022XfjPcOoi5hIQYD9EV
+MV24MW/NNZX+enfb7ivQ3iHwHe9ea4eVvbvzRRpVYAr7d0QopXnrg6E9iylvQVB
11vwWHIh7WuhuXHDnpnEC0sCdWJASVDTMZGdoe298TQdcBhnLIX1006RI+N/6kFt
ZpUbA4ujT+gfNygy7Cs+yqcNe6oUJuG8kj/uo9TFPAjpNPop7p2p3xPlLVNw7SR8
edu+9txyCmGycW6m8eKv1Rgam1uaxy1v5rwzK20NcC2508XIn2taDEpLcRTCm/RR
wxGx6ZykF0bHifJJ5ze1+02Pu2xiNatcOnHLK7RGvv7TzXU3xB/h3XXBI4Jne7yE
WJmBtpkjTCEojYtB4+8ZG3cW1Vdu75y586biyYbLP4gx8qjWbSmz1eU/iQ4N1zRS
ekbEQpFHtqVYJ9f69TC2pEmsgBTis1JQo164c1KwwogZicTTonKCXonMuiaZaB7o
zjMZ3j/1zQ4zXQoxJuaeGCsARNi1k1R+EDGGZi3fTqsv1Z4akDXXaWgeAgSLR5ej
wJfjfepkqcwZm+AWj1BBQZ8X46kCbROUllqyqI9PNUbaJP0MB5Liya1D2ae8NxXW
T1jXuZLIi8ztdy2HbEzMHR9sKe+sAmmt1967aDwwf1T/MDoRaOQix3NZkPmCSyWn
bgav+4ag/udFCkN0DKHfjpZz4T9aYFTy5+T84fCuODxBDHd70TvpCZfL58zzTdMv
3Wse18tCAVJ0f3GKaJS4e8+NDaHsyKdIk2vgzovKSjFP4dJbZ1/2urYR5G64vNQR
w0JMwy2cQIhz4/pzx2Er1T+EeAGKRyRQks+YNr7e4Bl2VVjJ7sYpm2yUxGD0eG3y
JSxJpxUuZCF3Y3ZiiRuOznjL+2GCprnSz85zBHRnEKQu3gkYLNSbm0pyLRkW6N9R
X+kzJk5uX998pZ+AXH070u5sEnnOGIeiN/+32HLac5oiCtrMk2K76s8/IWF7zntq
sSRWcmx/HE1Z+9D93/URyaRcQi5NZv8teZl8WQdBaVPMmuKgn7hUh/nTNFR4BkNq
xw6LEai3AOqV5JYJfV3CsYaFDLt3NKiilUAVG+LPqzc2Mu0v7uslvWMJKTQgwn2P
vGEqxn+VpOtalkUomvOH9YWJ9oFiY09be3lFpt5hTfyiih2pZwLxL39CBB2QIMr8
fWdngoQ4tL7bNyOJLVJR2Lbrm7Aj8Fa/akrrAyPp5SojAYsBB6Drf8V0vrBculv+
Jduu1XJOF8XaMe1naB+vKVwFclAXnL1CwHPx0AxEzaPAcsgBRzHdj0YA+V9tMFkN
eRi6RdNxHbRB8zctGwEqu7t0sS5qCX6x+/FYbsz8B+gJBU+hEli938Rw97ePagd1
6Ea8XG4EV50i0+fx+ckiw7jP8tByqc0sebQ4FzgU1OzRHl0hDyzQ1t8k0iAMbCQi
kERjqoDS3joj0T3EP7Mty7BlpACHiFOcGY4UvvHq8TIb8Msv4ZPK7HIefHNCgsP9
1ujGrwy5D3Sl95ASWl+224eHEBOtMMbBcixe5qoO/ANMWSVI8H70mf1crCqawOa7
zgnPLLxD6WfI9GUG1GRRQIcgxgKGqNUPeTmcpGqQdJJ4QbsvNocNsTHhlcBYswmg
F09SMefOjY8yv4Gn8yuVJYYm/FtmqIsZc2P1PQRozAvcHab/9jxjgGqM/gLQ+PvW
quOnOPNe0oNztkvyhlmFJFYArHcN+nsH0btvLhjCAnZ8tKMevLUChiwMGxONCVXu
AALFwwbVZO4a/ZlEIKAM5l7VELS2dqQuiqdZTnkOZ+chHna2mJu0IlSgPclGXHJW
o2dF8fUo5VZYC7Xf5xMxtrEyLRtI5cknlE3JGM/B3ErvATAYoIi4aKx3+gQ3dZaU
mEnnF+Ci3OvcWco2dIOqVT+z8ZRlfSTV81eloDbn3dkB8jlp8QyQhV1TIhiEgekF
nDrUyDad/bztbQyo1uzFnRPdXNoBMyJKLEXN+KeLEsxtfgv//5jPfz1lLLOrrxT5
ARANuUiz3ADhseY2XsOD4OidRAcjlNAgrjj1DYizxOjs8dunZsgq2Soyq585K1gS
mXZwqQ0BWBIEAliPNnY3x3+8R6dDX9Eu2Fda5/OmdZlxMALSEGZZ868ExzsaR+Zk
mRXQUmAJGsC9d55JLxVZM545TENDY2Aj7s0FpQ7NiicmDJCdJ+F6tg95w82UPH92
ysHAiREyrbY98UU0crj0GU/+5zTyvVH0T0H+2N1sy1K4DJfiLffPAMREJ+s555W+
o1VcMWAc1Gs0vK+Krcu/jJP1aHnG3jK+Ew+axc8hN6qyMa18iL8IS5SAfHkajflM
oe+BOrSoYblZ7LW277hxM+Fma/uTowx141+qnPGjE2H+Qus5XkcvP+wf32UPMvzR
AB1xEINBZpwvhovBbXrMyX/L3lVpG/ry5hGhNV6Ul8m75Uw0L/S/+2J9hYn8oZU3
TtqBzgo5T/Ybee5vqR59bld4DuUpMn5KFAtjTOmZ42ZWrtyMCwEwI8aN1idSl6bu
ybG0S4lGXlITdUAln6ebFyXmlsMY8G37aYkqZhqBslTCCNjZW6YhCj/4O/ewe1ai
3ceNTScWwlcmai/KFYpF6gVCz4bno/QPosMHRGQjU4pL8nWQN+VFSZpmiZ2kwQA8
4Tkq1qYspX5MUAmRozvdoL/q+AA+VK5r/GR2+CaODzSM/qsb8dp9qGO1oBOqpjJD
63crwWR3ty+lHCzzAYvg8H87LdpscwIAC8W1Pt+IsbZyaq1Ysz47BEe7wCbzLB6T
EpLBXa9UG57ykiu8wE/H7Ci1G66V8dHrAhGKYmWBPUKN3p4dGYzwrQ1pBiISGg0Y
BPfBtwzQ3OUhLpbyCuK/uClwDYMoqt45wnjmctMvCP7Wiv0854e0c4FpizC+Qvep
S5WpWQYiiS5UqEGi43YdYs9jwM2SnDNUjUx9yqZHeTq7vzhH3sBtCzxI6vrJc7c3
G50w+/vtaP3IHSxUlCR+E41Vj3GEK1o6b6I68lgdYT+zra1sdYqSCf/ieChqi1/5
+70Rg7frO2EAh8a16rXW9m85QtL7gqQh/97iPnWypoGBgNqKi8uGb3234CobT9Vt
dBLuRgRNelF8pTV7S2M6k67uiymTb4pc1Eec4j2NGRFKqM3YFskroek9xAHOaBPp
QKFBdDy2Cfuoq8diY9+35p+bXgpmtoAK00GdxIissDdp2CdN+HeonYdL0R+PxTTY
GJenMIe1GVq+cYQ7wjcbf+8FMElBfp4w37gqfWlItswCOG+Mil+TVGQy6qLXqvG+
DP2n3Ak44/Yp2I9LW8L3QXqtGYfNaJdAR6SakEu76oPqYkZisXT+ZKWIRaaHRHMP
tSd8Q6lNaueqTQIxJ8KjDJDdAcV0Xcrv/3EAhPQ5T7vLfVClEMNtQHzlqm3DRNYs
QF67l1Q7mMlK5XBJIsF49JCX9XzWyGrCEgw+Q02sOAc3dxZDbNr3vfRItiH3jLt7
L/6JiP1gmSa9EaY3rT2H5siw60OKVWc/DEygX+VLvKv+Ye9ZBmMOJRmvcR3RLNIA
5SjIB7oOwbun77ct7NGKCQ2pbIDhEK6+NJvA3WAS6MNHs6dGbKnMFXpsCMxUqXHe
n0efetvnnf7BB2TGHfPi9K4UmQ6z3ThJF6KRddW+83W3PZIXQWg5sZBJXyBSSB6n
vnzNtTBTa3MOadfCGBIRWhGMCyjUC38boJadHjThf48JsYv2lZoEWr2pT6KqQBMA
m+If165joW3Zq78KvGVF//YHZglOZV/uWHN5A7mnxxuGw3BLKsmn5TXkq5mNPU57
Xj+xhuiZkMcXTz1NmgqGCbO5DFmmn/DmzPq8V0JNVkfDQzqOVa1ZrkFgJLTdmMDr
He4JQRhxE39MoEK4mmJoxZmx0sPiy9MLIzMEy5Ma6T3l1C/Q5ossGh5FkfWjFbtv
TfnkfemKPrSAiYBEoit7tOVGe1LXhGIopJlTdjqN2cNc/a26L7aNCqQ8rmF30Vw6
xE/NGniiFMm/RG7FywaLrskBtrsXX4F/MEA5Ngal9mO0Ctrf0IvmGmO6A3dwC/Tl
HYPBm0X6apxJYdYi2gwAUL5NadkfLTPAss+rT3eRrVA+dpYLrLJwWOe6cEt+KnaA
0k9sZ9WWFjY1WQWfupBWMMvFDZL6O6Ewf7DOv/bF74e0bQNfXV7IUHEsmfrbDAXI
9mi2eC/NgY9EpzZK5gE7E3FsbAvW6pKKRTOp/RphcbGlJ+0XwkEonUBOjJYDsr+D
/Y1LfkIJqvehtGALUq1SPp4Xo9Mf5KTr7fyT4mZq9SVUD7zfXJLVt6SKKnAQsMox
VLa8d6QvOkf5HFoGI22NQESaqT+USdIqH6y1LvVmFcni2fO4/jswiSrV0vp+F+JU
ukduiJwyElLTCkJizmy1fYtomXzmID1LuY4zOI23FqSE9JqZQWDI7nOVblp7iem6
W/9stchJJvf9dT2YfUcOnGZ9Zoont5w32aaHL6eGkgLg9rfy1rwLeyiMdhhXGPNI
kUvTtLyq1ZdCevPwQc3HyTLsycIeClddYCzCGHCv5eL0PJsQJtswnvUTzWiC1lED
CUI2Pvqt3q+ogSBjgFXMVohhI2EeiwdqpSBJMwqp30M/2wuHcZMGCX29VZTwqJ0r
shl9xc/Waj3O9m5+FwPpREDoILp/QjbdfZ2ZU4sZajADOorbWFHKMoy2XmncQkpH
RnBov8WOKUCve2+J9pRJLxuj+gVu0BYfWfUu2HUyz8du3OT92q5ati6KJCGZkwH2
mipmvZ3JSnidhcuYC4JbeCin48dG3+YKLGLw4iSdyMWNZZI3DvoYJfM/hWGt8+fe
dfXtVfDbTJjp/1pllsnOqQunnVKqfG8J2ZWiXgLB9saRTvyBvrjGM3N8K851yrFA
vgGR2uSNNs+s9sZbdFgECewA+FWxLHUwlhFqXxZQyLotEozXAnKe37CDTMx5qKp3
nAZk2xdZ+mUOHA14neHtwPCCXPEy3KPp4687lcelYpsQYQ4SAwUTrzI83IeBVDmh
E1wQQKm+olTtjcSP8zBqDIAo5PZjsl2ZEp0YBD1AY23Jj3wjOIA+yuknRQsgL6LY
fTXtZ2iK6DUCQxf5+W+W7uGaaQSkBJbGIlDhTzUWfttbU1g/hB2wkuRyDquWUDLm
Si9rKS4pJVmLaLqaUFmzgYmUU53G5PR9hCemJoUPQt0VND4suQ6QEtpl0dOG94QZ
UF1H3L3fCNFOuqpjzYNUonEkR417h64eLrZHubfMRC6OWqtVhhSFATAb1LpehFim
Pr2zLZ2PWX1tPgIdKbK/ec5w1zTBwJXIZIFrV5TWBC5s4DjpnBAoLJdmSpIwaUB2
n9AUCbg0VgpSPcO4I+NOkBwm89w0B9MLFWf53ZLL1QmGKrgkf3QWBAacghaJBDXf
+wjVSRKvQPQ0KHdbwfs4W5mT1mkakAS4EOmxSwog7gn0X/mbNbYTnQIvj5E/NTvc
yfUodzEz4Py63SK/KlhTckBZ/doBMYd6jXOuFC51voqyNIcMbQk+dat21JhGFiBv
VxegOzxxGrqR4Hc9fkZ+HKOZPB/LhXkUN+wCpTe/d0EsmqQr5OFfpjcDKqpUrNsJ
sP6g9gniirpNX99VKw2eRSYtAxjtQcvaum7eOjd7709nnmmXIL5qSI+Nwmte+6c2
vSC9p/4+nXWHnMcB6VxK6irldMSnZzTo+QOvhFdstm5JFdc3YPN8BHJgqhq7Tyrq
jdRckymk/Hy4dDpVLTYc4Xx1zfKklxQD33fQ5dBrP/yH4oMU/PWuigq/DloKqYd+
OMSFjahiU2kYomVAXX8Dv4nfOFZ6hxUHWQZioWgSqFh2J9BrQ6sGMbow0OpISRrh
4keteQvCRTQ7ioykvQh7ablUb91WlBRnw4dTOWWjgveEVxkQOiqN/9u3D5xSAs+K
+BnwWd5LkCR4mEMgaBqrbDtokeUkM7wO0LpwT19YtvI4Ng0Uj1mR6GlTqDMBCK5v
HKKEYzBePfeyLaXMrUrREDCeYax3i7s1OPY7ZNBmBatevDRz2EUWrfrM6Ga/TlRN
QWih1V5BqZcajVmg+o1jSG8hjQjyNX9EbHx65rj8eaQ040f+CT00umsAvQX1rRwa
lJSSAauMDdiooFkCG1cNx4nlSqSOy8kur/ySKG8wSPWhzsOX9DmdU8VquUfd/exS
CryKVXc6itZqEmnzOYortm+YflNJcaADt3PNA5OjdRcOwxHTKfTTP9u5Jnzh9K9t
LeXxPqysvNSGg06hc7IDb2PCCANujGAf7L2RsXHgFTs6J5IXoCk9JVhGFg0j3vDB
/78qp++pk6P6Bnup2CTmW0q4MEECLzHyfgM0oCM/9B/ePFBSvPf4bWntkZ9QSkmq
LdveRI91bFJyugMNiFIYR9w1OQZhPQkTvmZ9//rdwUhEMAE4eF+RCU0rTFV9hD0x
8wEgMHVb1t6tf5PVQ0LjwUT5ZoOqR9ijcmVXItGAKIA+5CvRJAHxCW88PBmDpAkj
rZdhbsxhbGt01tJam4GHoG3k48z4H2fbCJZ9gEyodPe+USrSuM/QzawK6OWQdUZm
pvlzvzgT+cIiBhHgZdB1HRSEBpnk3p8cs/gUl9zZpMvKZMjqYp4FbXGpG0uap+wO
MC9A8u1FIJqb0OucIgxJUPc6RtO1aipircZkdOu6cESUj6jWvGZxko4/b6r51cx6
i37CaLdg8SzfXm3u9DuQsbv9UQ3cyFh0X+guNVY5kIY328kpP1PF+qNBnMyN5rYJ
g966Hb0fBX6KXIdInxuyHlh4IBqFjpqVC5PTWEtArlt4lTKRZUOhU6o7z+Mrv6eD
t74A7iX2onpNlEMuoUXO2yyGtl4IH+9APDja2G2CL0zsGuJwshy6OrMCVzf6dYdt
fMYgZGTsUMofm0MsjpjPjxwcgpq1vpTYBRzDcjV0v8xEDAO8DjqEjY8vU+nCceIT
K0jn5scpUsBU20Kk0eT+21A9PEA0AQDwfs3X0wF3Q82F6MSpfGLPLc8P02H/Tdyi
MV0fb0UklledarKGfAoktyL/ibo/jTNOCyBKE/O7k1r6VHXF9qsDA0rOFVZTjWvV
xQ4ziqKEL7v4e/Omyl1eGI3iH/lRbPdO9G2SOYb+x8o3+KY7iG3Z/xk5IV/E92Ob
9Dvm0NlZ34SHDtLzjM7FIfNXUJP2pSrQYGXzENrwH7z3+FQ0BVWh78PdOQV0HcV5
xrUIuxSsxaPjGBHCz22zNRZC9F9OgcyppgQoWVLJj787dPWzSOWviLsAWxKZMCPX
71bXMzvr4gfiDxLEqyF3qrCNgqv7ygEkIOwdflWdQfnoQ5eenUOGtPBrIDrkANAk
1bNXBvlEVctbUcyKD/ldzbhyOSUIwpb82SakCOp5TAC4BaHGtdRxH4/DBxqRdcx5
HOBzpaMmkj4HIbYoNYj2FvXsEiz6sLDIenJMe80zLTRtnr/1qbjb7+6tm1ErFIvi
4VCRuZWTUiHu0KS8b6Y4E3eeqI7SBUfoRVJ8qKHU14vRYh2UHw7O1kl888HSFPQA
aTjT3RXmQlOIErxkHYU9DvzV/6ixEa7KakHn1Ziy2FXmqLjb+ZZquoE8eFSZMz5Y
5RIK9ri3BK84LjNmhfKth1HQPPVeAdiFlb7G4U4VST4icHfn+Khz7WN8Su0TxP0M
RG0wd5wMv5EsuyqCg/U03opS2+ZJCDf9g2UWtB6eqfzFCINVG0+xuSb7mxbYTAho
yAqYC7fQO3uSWwPU+h1t9YvuTMBZiipgq8zdEEGxBtwQPz3IEyANw49mjP+r8bG0
RIQY8iqI2ttKkKYbvBYbqEBTpWkKAVsUG3Zh4wY9UDEH0Uc9XU8iTDNpWQrNMIUk
Row5btnUCSEX0KuvVolWEpptJZRMjZgR6UsjK5oINvAqdi14hfw2AX7+pMkuL2gP
h7Wk7Twlci3l1fsWtB+IvH28YSfcL91bgQyEAyd59gYwWCTpJ7uv7UneOkCrMOmq
MoD4sfObT3UKJ+f6VfeGVYlw4xGwCTxgszys08dZrNKd9vt7b+k44526YgZDWdHZ
ZFibqWjthSTxqfBAKm1x+kjBFBqKeUXTxxICD19ZKz3S9EMW308zldW1PiWEbYhZ
yXmkikxbfN0AEA//jQ6E/vOzNQ0P6nSRu3q6qbqrEWZM1dxJaoOMAVRONWjXLR0R
8xfL9juN5bNRczBml+hsnpxu1S11an8nA/0rq6wXJfVF6MeF5UrN0XdOhAtq1fjP
Ie31vlI3XsosYLUubm2Mr2pusR2omRq9k1HqM61DtN7SKFm+MR/73tObuAaVdaaF
UOAmLz+xdl3RFJb6z3LtcNys2xrjOHaEsWIxnnFJn9fuLfz1EiTpq5GPKrZcq9AI
wnBwQ+3NRql8RdWlNTlvMuhj/PIuL3CekYxNmQhKDtJmsTJ1bgGvOizWl/J8K/7U
vzQLRBr7c5A5wPygk11pRV0ZC7mPP9IOxyKnmaMo7W9yaaGx5HhJ87XclU5tPDAd
Sbw5EIcjCUhuL+Hg+BeGMJ5to1Ub/0bjy65czadGah/6Px+VEo2g4PmRYdSL85pY
bDD2qKtb4TD0mzClAJf9d3WBvlAEPG8oszaBHwxdxxdhFVgFIKSaRJD25LN0ETRO
LojS3KWC90lGb1Lk/paMthrDtpZ+5u0bAJxg8mmON3iliI8iRv2w2P/l6TNG2g8d
Dh+PJgDipKko1s0KaoIci5DmZ1Lfmn4LHC2j2v8saxG/iTud2WKTppXco6DgBoS3
Vad0SpUYMw9vJ6Ij58ucL3UfIIEplh9i/e00+7MMyR3U43F4vz41p6uhM6xf2rKD
XgIzeRpz3Lh4v1a7BwW6hrepDj9xTPxWhVl1H8PILyNM6G/DwN5KZAe/PxLGYsst
hsHOdM/Ex0iBDy4F50FjwHuNmrmhMeFi7ZVH2huk3xkcYaBPKflb1emSeQf4VsBo
N5KBUB/1CetogYwjFqzZvMjqiKIwWjV1jZ+38bsigRBzXKB2fvtodlsHUq7Cy4Bc
ahror+QzZ1t3gkUnh0Vb6vcjVbFFYDic0y/AKU5AvGQm0hjnJ+KLPsjVThoQeE4V
ypnDvzy5/0RfekzeJzjhgAfL9T7fVNzslI48HMNPYeB8i42Ha2e3xxkQgsfpIqDe
W9AZgAjKIu5dvd4HeZgkhez7MYma1G6kjVQQ/030MhhgziupnLKZDoHmiOZhpuTi
niKXoBZd1tGZEN/k2F+cDfIIC6j4zudIlcq7dcaltw3LigLH0NBnBWRmgr7JDuim
i/rcE6YrPZ4JJeQoAY5UfB2fDe7zLPINegHUD1SOxKO0MhH4d/1SMa0j6B2K4lRx
gc2VGRa0j9nAPCOE8a5UDvmhTbo6TkND7NeDMVBYkU4rYGrFCZUiG9UwjX5ALWXX
bSCfGVBRE3CE1crYOPZxnylsh5DBCGVRBR9NXnEavigabB4c/HvPI3fWVDaVVtxN
X+JAFeqCsiVmNJKkR9Q95IEr3htZM5sPq3CzYMDdGeEiiBqd2dwEi8n+kB4+Nnbq
ZD/zo512H8zCHJOAaNqcAx3YGt1vGWcoOmnnQT8vPGt3Zl02DO2xMz+o/EOZT12v
U1AWZB8EY+IWoNBS4nLMy18O22MTcfziUvkRscM/TkBmD9G0hqd9oZHeXpXZ8spk
TnDJbkWIK0rX7CPpgaXNv/oR+y+1vVd1arq+J/MsfqGOB/v7yF6XnXfVM7op3S45
sdGHu3vpowN3E+yS+rDH5E54WtMRNR3ILlII+GrgB9daomL/yk7bAml+lld1P9GX
4ndJQMkoK4WrpuCdUSv8MLXxjeIl6rjHQ8aBvq7QjWViyReCYTrBtwAzUgXzRfSU
jvChGTWIGE+23VIMYncv0gltdtRvxsG+cWeplq2k0vxf9iJGo0bKd4jpZGYBSAY8
NyxEHTvUCdQVDn60hCQBesD4DgGtt7GTol4lBvCJaKbZZ7fn90+glQhYBuFxbg/H
bn4LcGFph2exxUULKMZJZfiWVPckbQwdMw4/WDJtllKcqU/2tGv22ybIMV0i+a7w
cFJc/9SvF1k+NbkCm2pq8qQKoWT+kUmM0QVEEsI+MckUiIoTKYe2CElxRGiTenH+
Ove49Pedb1PRIviEaywD7pD+dQoLfoCw4S2HlmNaTWZNkJlOhHGPnlmR8hwbs2Oy
D3tQftmRpDQ1SfHFWtvDMmN0u/T8K1H/u3O9zwEh2We2NDudUlTxRedIA+VpF/CD
U6ByVn8ZIH6zMAyltgKm2uNN8hVBaFTr0ns5Fq5u8ZmRdLsEUqnDMuNvIow5kexi
HULitG2WbZKaQyn906MYBwUeaKVbAvRqE9Pd3OXakpng8sEhstjKJJ4QR4GhUm0o
ACiFFTzDMtzDPigVt0wg6HE+90mp3fYmkgFxbcPnnPnzhJ7QuINNxGa5uMK+sXMC
uUnAO7JnWosCiG0wnJIsRSdY5oD9QolULUY01jvETg7hIvjw6KWXsoTEGut5EReT
ykj5FTAPbjGrac9bgFjF0AuHyRkX+FJ5L2EPONFI5TJdJ63zux0/uHfODxXlpQpP
8P++HvruyBYkgA0X4qhORFTFjzNkYSyGMokmT7Gjr9atxqtNlOnlPrpfibc+3JIf
FSeg6FaJHBoVIZEt2K9Bw1ZyPkpwWUgTUhYcPB7Ed/0QNhmBtRqDaap/SyKPYDpf
ONnLcMhAOLIPF+kmDHMkTuW5J52z4umoJCFJTSKhw8G0hLCSAejbQDdCxOl0pnFU
InkiqpobkgRJruDSKzsESvtBm/9On7gIRijp+xZpwJ7VAwzntIApaDK1/0iQclv/
nhq4x4DoMkzUtCgX3EkABAInrYoo2+U9yTwMU1+MHTht1lAR6KTQnBVEELaDLYlH
qOoRumstU+0PLjvBpthyImpM546C+NUvqBpLhmrTAXtKk2ovtFrQ+ZyWn9StO9d2
G5cIfVLBuEft3zD0TuBvk+W7sQ9uqgOt64rDp1OmpZ4+kH92NwfLd09qazV7Rra8
niqLPVbE86GPFXjJxvagYEZCufHuqjVWkc5WXFxzq8TSAb3RV93SSgr49SGmd9jv
SjzRJiDyXkaPW3sk05HrNM9TEkNJyKlo9/R/UmmvX4xm09Ohm/BR0vpIayTwA29D
QTz7K05Inh8RRv6xD3kqDwyYRWyTWm/8S/HFhIZb8VM3Pcbyh0pQ0Cm/j84C0RMs
5lou6rxt6qYjKfRuUmLelnFFV8bDWD91mw8eknA5pkIre5IciSEpNhpPRnGJUC32
qEBIImuTkgaPbf0UhPw8quJrb6kisiXzJlcuBW2bO1SPPzx/g9dWW+7+DcoVv4xI
cYzWHm215zySbfspyeFCbOGTXc5RLX1R/NFq5cjb0Jjel1xUiupShky517nqzSzi
Rh551KBETc9MMbUeGvRMRuo7xM8W3vG4aTDx866oPQFr3efrJRf1M+rjO//DjWmv
gE2+Q24LOJD2uCjmlzOa0oKKrGs328LopCWYT6cLSWx2UWB/NMzL0N69zwf7Erfy
NmZkI1NQRxtV09Hv9IRuEZEHIm/Jnkf9MJot/Cg/6K8gGzsC/EwMrZ90s7emkqA0
29WykSwutGS+PQfu+c7Mvql/a/9WXK42oGMeVfWqGrQiPs6A+JDfcuB/zk1GMHtl
wqhqeCYddvIJcTsCfJab7Y8L0bcspSVWqKC9UqiDVyhUY337uw4LZqF/QxoB31su
jV7GIPtO8/VvLanspBq2Q8mw20NoMUDnatXKmzFURom2vnANsfTyjonhQZ5HAv7l
9l7e32Z+svboo5BY8oVp98SaT9/7tGVCUtMHYhyuYR3+UoGz/DrY0HWPhokmwepl
9WTOeybin/tWfp38rHh+4/CMv52mXZhPBqYKTac1pze8FLoWKZ79SyFKT/58l4rn
xSvIeNdkSMchGrQOn7OQngv93OBD7hzKDjGzIwERKZ2odrhM213iPmPVZxTqQtVh
podIy0zzjw7K8mgPEQmlpqkoVj+Z2Nu6KVF4TvzoEYzxg6nh8T3CI7JMT9QIdQLF
5PWHfpi5F/bMC15L11Lp89pFRm5IEaFjEK5l5+Yqr2XuDnGxR5wSClCT49Sw+XzP
qhM0C6fKEePDCF4OQ9HJoXuD9LungLKIzzoajKW12772Y/Wt0ZewFnssIqtWWEYZ
T5f57NWaDEOMqt8Xi/pNky49/rfApBXYS+6HVhsF7WWPuNRk5GPbNv1JyurIMDnL
ZwgOIqrspNfvI10Th3a8ii3L4g8f1fObyAn5u+9Vr1N8mlPIkfybm+zy53RjhAzQ
CkhQdi71nikhyVNAz+vBkcFOUAm4wGKbFsLhri5K7vg5a9kUxTvat2uC2h6IBr/e
/v6bMM9bS2gkoU42cTs1yfnEWjVCG1hA4iSqOfh/f60H8WIN8AyTsof+rhSezukM
9i+PchVh5BJAk9OwzQwSbEV5O4Se7UujOQN7SHa/aOy2vwoXWCInC2ra6wQiYVhP
MTNBy6GJ5hKpDaO2ZqHFnIjZlP8ADcVL7RN0LOgBQyfMPB+KGpL9qjj8gF6nJcoy
mmnAgIMfe3M9A5RAzIYayZunH3qRWOGn+RWKS3ZcBQ+tPtFQJaLxvA7bjvGOzJNH
74ugH7S0ZTVrzBikmhfGx25kMe/c7MxR07BMk0P3VlketsB0E+YdYPLleDgnz1Sn
Y1o+z81zVmxaDI5wpTq4yf0OYQCWcFAqj2fPSCIYiH4O/jK9GcVbm2keQtw6gyA/
lV3JLKPPagM+uDTRwYNUN4eYATbCKyjYTlRQC+ENuHxZseKsAcnPUnBxl5DLk4gl
MIau/2LpcpXenThRpsAbWLv+DZwXiq198FCgCWtkmPMHgSyEIsoRVzJt874FeO8u
Ig6xwaKCwYmQdHaTYbhnmXYJHDaWYFZffgRfVfEL23wcIIXCDPQiARBYqML34k2Z
WGpaqmA4oCfV4UBXwhM0qiLus4j5lpvuNE8kgvA5iAtq96ZEGCKWqIRntm/rt/M6
YILgCdcrR3obWmNrenOC3IEbiNTfdwsc+31tTbyJKnJdobxOaqrV9PkcfZBPZx8M
Buqd+X5qP68E3uzgDfEDOP1dls3i6yIGNm7Z6lHNjD9/l0ifAYKO5ieUFgEpzIh0
iYgG9sNf66FOpRoYfPixz2gZzGzHjEfzPIlLllDm6cGwr/cSdmJMxCth8fOMwM9J
4TlHnnaKm7yCohVwfkidr7yDfYA1Y4D62CvW3k49pneaSrsU9Ug7jjOGpo7DsC6b
Bc1yJ1wh+X+kX+1xR0YxCGF6OVa9vq7n7P4lLDnh72rttk3Whg7dhgNa/YvbKjII
CUb3blknYH49q7rlILtbAKkN8o+owbObi0kXUj91EVUPN7bmLBorISaGAqYRZnF4
cpdUW4P2/sw1fVGZ6Oy/U6SQTkFHZh84MP4iwu4u9eS4OQ1ES1FlR+4jJ0zUXezb
V5itnFV5d++ARoDDj9UOp6X0IRzEgChVvJJ0RLFb9QVKpJ4CUT76lUN4ZcroJeyQ
wJsyUn/QdVd8WyfCRWsgferMlYjb1i3YVgFpdbB7ajgWIE8DINt8OjKpE0Yt1FlG
i2YZxk94HCDeYF6eodeo2WoZxQfTYq3BfQ0kI7+CQP0CTLdC8eeOqssoLL8KhVlL
BRB5b8HlztaWWv6G+TWdrqLIqB3SOFPAT1mcsyT6+HMeVxNsnhiRec03ruRbUnBe
QASQpuBYi67uw8xDfK6z2OZp0TY1XrZDWL0f61Yp7T/566t/laTXNEng+GHjnXup
7C3bBr0FA6/bKKDLMPMoOvMsEoXTR9MClxhoNPpgQvpLkdNXo3uzWkDipp1d9Igs
w3d1y6igakhwOuNRiqHAw6bDuL/bV2jTaCWiNjzBhEPE5sVd29vcSXTxEoWakJiz
6e8jsgYuJvwLbhkbGe17ULP0sWaQGP/Lphd5XzuWGD2TeWXUC0Y3/p46SHilsmtM
iGJbzK/HF0Hsx0/jENl2z/v6gqodRFFP9qCuvumQLL1cnL+5aQjRmHo5SvwQ8vcU
ZevBcaPHIwM1l4O080SEn92ggppJToE+k+vy8X2YGYMjG7rOTIpxG+x3rqEVz7hL
ydP/K6KYqR5wJ8A/cOMvA4Qa+AomsyjEhS7i2WMl/AzM9xJ1O+Dde11JTeHu2xtn
d0+u1/E1BD0jRunfcl1eK1Wwe2Ln9i+Nh2MHFNV2vM5WJKvwAKxzVa/w27Hmp3qG
UFrWp/NBEaQA93S0j1o1SVml8ZOf/R7K5kPMZgMZpbbPVHR4qnPTwLTXU0pgrIaX
nvofkAdsY4yJ7pYUUv5mM/5wU/aadAjTfXDjHXLJQJCXyVDrZzw/RM/gK7qoUp0G
kbrq7WROASwOHAggkoyh7QwXRXjVo74ipHvfA+3eI0oYB0FaPRb+ZlkDCYIxFLFK
uR5KC4Srnj99npJaFIMzadAq/dqnVCaVTMc5435xXbkkJuDWejj54B7W608BQqHa
7pPUyyPhdVYOEFtJN6UbxoYhcYORBz16EOqSsS3JxjFJZKMrYHnTwCeXuetDiFW3
DKsUT3+cBRiqq4M1rFYzWaj3zLvbpB0jd4syZhA7i1eDIX/DfueHC4AAoP8D3HNW
d+mthL1njXNey6ZFumVa4TxLI1cg3DIfHUngcVxog5h7rJE30K6/DFDYtPgURi2m
Px0w0+G/krXFaWszmJThrE9OC8gO72fB+f/kEANSrTCQEluhf+qg3vnR/jLu8tQP
xoP7ItCTVypk2nBsbvDvCQTlE7PLzVKuqfH3KeJfucj2ac8W7XUr43xtdNiZONCG
U4Qj4lUAECwiaZAeKPRjU+SpzxWABHERlaZxVi/5iAl8vmfBd3IJIpkpX+jbr0Md
jbE6UYRgzt37+81qUAdi10Hq6FwFU0Ryr9BcZI3MgQWt8XSTyVoyBkErQPYDQj1W
C/2ryXJoUw1nRkgt9eX5h7DoefCHbgYCLsmVlRZuj8DxTb5QpcOY86J/QQxZxbT3
tiM+1xP54Riz+9QmX2o7V5w/j9xKsHIQqIU4pqDRRjAo0FsnI07yI5IcB6PWPAnQ
J/7N9woRbQJZ4L1gvPsUjzOeZOlPjV9kDW4yTivyHWcHBauSTzexq1O17oHQCIvE
921bAQK2NBqSs/0PwYYqhzaIsgTWZUgTMkJayxYQlLoqRisI2S2LxhGn14mcNzi6
kXLenSR0Vc2wTR8O/Uk/U1CEbni5PPYQ1TETWL4+Yo/f4bPDQ43lPsx2r+WTgNiN
caiRQmJeUQI9x7dZpKrL00T6qAM8LaQnnu25nokjafS7KCnY22jyINrQcYFsIO4x
risBX5TbRu2K5btoXHpotYu1uuXfznBK1YnOIpI+VS8=
`protect END_PROTECTED
