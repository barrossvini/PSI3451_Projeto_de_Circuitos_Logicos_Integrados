`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ODbgy8mPNMsU7iYGjCi3kAVT6fULdgS933ETX8sbBHVDzPsftmAxxgoZmGanA1x3
0N+70JT09358icD0GuSRmn1vusMRbGlghjY+73ITbfTilaSf5DTVzJtRJqhpFzCB
HQPXJW9k471TIKsQnUuWlgQ7saf8nqrq1JHeCQrt2mURkGiNvb1X27JdyKP1JCXC
AAxDK1XSb6aiopMZ0gCfimg4KM8pdldAwh9y4mg5TanLF81nPzk3nUp4orad4TcN
5UjPUguknx4pFJvxAYd3W6XN3X+ChVORW/D6ANFln3xpla86Ni1Dmb+JPcTSScDp
NSttVe/bFh4jvcw+Tj0eIBhtRYB8cfE0oMg6bElyau9a44HT4Vk8KsSy27PewQiE
T8fGO+9B/7xN2j512iWV4386AhTZSkAGQ23KJEJJB4nlovaiOK69md8lGgQWraCT
M8fZ/9+gb9d6Zieu6pbIlJe2jG9j76cJRscwi4LfkwRlU1oY6BIgfQ/9JOCKaEjM
ZOnlHLx3GYCFwwCUVlSGINYM5/QEBNx0YE4gmjy4qxvbgr4yoB3fR3JS3t1fLPuO
4dxOldMVWdc5N6EDQwp2Jwj0xxmc9JYaszdUfcMzK6k=
`protect END_PROTECTED
