`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HvTDgC1C5198FcyJZjgixhtFtfgWH8XNd1B+cdRe9c2pAL8WZLQsLd63e551k6NS
SlxaxspeN179FhpI9cL1h2q+lP1eXNI8dcF7t2SIBCifDdkvQEd7yG9DjmQ6+IK8
30bFCQ+xhqMOlyNSrZNwsOogGryx8bBMpa6V6a9jslMzYatZuiTPi8idcU+coa3l
eEwKFGlYMWQDzg2k60nZ+kQYCNtyezPTMSkgVQYonE3a6LVxY2xtc3JfOpD2SSCz
tzVfaLvVDBx4HjJXs5/SNcF1Pe6PwpsPBzlZFloj2otk1zM2ni4OP/ThBQrNv7GU
Zg5LbqXSxLM0jAyOO+lUCzdIB2yzWFkeWvDQPB1ztdnmH03PeYOgsAYf4u5UtMDr
UcWx3n+OSJq1Plgz36oY0EIHi4ToKuEG7IflWlJjYZjHXfP8IEmpZLeMItKQv10+
9pVHcpZxlDsy9zeFtdxFZuPMj64EC5Al1SJrSMw5xzwTzHDlQ/2/2lxy4avevSZQ
3vMbS3pZRDsNTNEMIXwrShK/yGyc8pU3VoCAm6+2b+ooldw8dozow1BZhL5/5YCp
WWW9LLRyb6lx/ORBqkC15Bf2vMmsZ9t4gpwnmch4hfA8o0yqlXjQrqpXoETsXh71
kpfdtu9ViYcGMZDA6jBJk/ZTdWv3eUmnqabEmzbKaexNeM/4qDOHrWiEW04O0COJ
LtQztY23TfGMuiEIuDjlFrAavFwPkGKSPgeUVdZkNdZ0xE21uyhjwP2x2fD2kY6l
lU9OLi5s6d4GgAl+V2rLuj61XGVPJew3QkYaLvVvVB3qikGpNEheGpu5SagGe88Q
qCdDNOT347Bjlj5SetdozoMCKMaWeqyTdmj/Sp6RtjULwxaXYMNH3rtuPpSxP1FE
c6usJX2Skgh338T4i+G4hoxNRB2GYnhPat7/EUrTdSDit1L3crOZ87GsWKle9Xfa
MusbIn2AA/f3YELhwi/C7RkU5kg1ptOHLmhxU8/R9dKnHrPI229l/rvYQE6TMrNe
GEWhy18LLbix+3tQ48X/mDsgTf+ooa/6pI6R9tVhX/DuzzsYAKN97NOmeX2ENh3v
oPY0SirpK7V05a99AYHH6cy1qZhxmHabwXZoywe4vBP2yffy2VKNFhhD9j6mHR3g
qfyVaYvmeihTGz2AvOVg3SpwkH5T0kHlrJ442hJ8tP+Q1j+Zt4rpUEUlYOca+K7h
m83zc4jx6eqpJlfvqGnhegcwsIyGharHMJ1yv59wjIl29qsvPCV3LoHbNdWR+2Ag
IfnyH+SPzTPLa/uaxvRAxBS1qws6Fwxs0Ot/dChD6YhOKToij9jSPXejVkCyHoYi
zeV3Aaj/7IliIk4eHlOfsHjgLeX4HVAFOQ1C5687d5W+41fpVcTi04oOIFgolTmn
n0unLF3q/zFbbvGiwFFMhAViV29KNhjWq0wQwAXjOH5gEdwS1RtQIZYVtlBks6uq
nr7KtqzVa5D9nisxSjtItVxceElIet2g2xeAI00xlFM1C3paYEzUwz2y+XU+wZZN
uvEJUN/EoeSFkZWcPE4Zo9KPR6eS8fDLDoald6UYaIdm/yKd+kDK4+W+S0GcR/IQ
qN5I0tyWc3kDnz5kbut6/t38o9qhAtbBWuvlAM0MQv/FJyfO2YnLqxWNua9LFf63
Gmv4agHz2eLypYpzKx+ZmwsdzfC4anmhWMzpFdTvA/4DBywPV8cZAHnWIaiNG2Xb
d6tu3ntkHTESDv8yo2O8G5VBk2A6Hj4T8YUv2HYVkOtAzf8Mk/qO+eowPfU9mE5k
e/M6WmAeWijANSXTrSzdbOtJRC0cd7JGRsj5z63t3OaAvNKdWyz/Eo+jLISltTzw
y8eSvaPhXwVYUQOr9ux6gT+hN9iLegQqqhpY1XfdgwV4hm2CBAgOYPaGz8iBFXmX
4GwCwxB6OP6GnrGfwgtMSL1Qhy/kIk4DMgm8/nnEs7Koe5/lCMcumGsqA3CSdyOK
Gx6/8S6txaLbI6d0nrfHglUerDfT21c9HAmoPSB7OC23aKn3ZCrKm5S5yfq/agae
yXFuMM3GfAkZZJtHRy7nBrR1X9WtdccVWazQxQfReh/qzev6MX755XibjCSpqlDH
gLtieDkotXu2XZ7QSgpz4zQbg8125w6TX2IXVIyiGZvTANplm2IItSXWLq1yrMEH
z3/1x0zP54ojb48nP1W2wEZ6aZtF0wHVrQfCVG/HxdC9KM5I+RV5wxa0mZZouRsa
vMqaJnHtzKzxMQxtsWsxicGgyXE5kXrejuoif2alE54dqQJsDtk65X2IrtcSErRs
uVVvV/6a4lVeOFzD/BR9vY8fqRywbxGk3cwullebywoImy4b17dBAR33OooopGIZ
H6+gKWElzNOdEIXGtahimv2aMZYY3rw1uFoqwoCZOoFDx7utz9nXIYhzvoLmwbh0
lcrSGe8H0PiUlWOIV9OvH3Eu7iQ1HlDeR5eIdrJ4FBhvuh9t/ZMk1zD0adnGjZ17
WFjgvUezt4yaoUQzyEZK89r978+Wx1+Efr4uv8IQk65lhMH35qurFRJbc1y1fU4r
pes5EbbQ1WwCm6mvBH0mIe4+RRYBhnOF785LBOPxYdosC9wjnKHeQMAfEFMfdJbi
2kkIJV3LAUZJ3OSNZmZ8abKLyzqqB/cwf6zNNgTQjj17OSb8Wvgs0H3olcM8Ri4+
lKyF162hCAxQr9KRxfOXoWItVyzvrjP/uso1hHULso2l2X4OzHzzvcj6l0UUJGkY
`protect END_PROTECTED
