`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PT3yNCXG30jc1dHagM/qLV0qxRl+g/BKjHus7ntWxtJejEkJ4wVnANAIoqAsgWdk
o2iemmiCeB9Nt05jBqc4m7d7K0QVyZ4SX3R9DyKqAiAJslkkbMBUkzQk5mx0wJJ8
KQkgV7TKTAp46wEdo4UCzSZ0FGKY0WcFBV550G6hwFM9ZVZdCZrg8H4E6k+BldWx
rF2RXCpud/ilLTN5Q+njVtlaCtLBKyXB+slCEi+y+MV+mdEPUvgS/CxKywUZfO8e
orSzvSP1EbxJ1g/HynjtVUWI4jwypE3Jn2MaHeXlhoYtDl7PDPahOQFDF9Jz8mQG
qPv0Ci/ZvFqdobyQ4aTbfqxbVwIf40DhTMPit/j5Nga34n/BRe4wUyVzWq2j2wa1
8qhvGwd7adkiI0vEb2k2gjJkiwHszXf1TAfjUm+FqSBtLSgnSAOYsMS0mKG4n5RO
eyzXbpIBL3kOKn5Lp1FNm+1rLdAo4HL4uuGeUJQbe20nYvvkFp4COy5rJxc9AHsX
3rLiwsglnhQLU2vHaFev80waaKE298jm2JH99u09+wSS17A88PNlKPBUxdPFQjc2
RqYH1N1LIigt+FL72wCvBg7i3hD5ZNEXLjWKHPDg9JMsT0+2TILnV9gm7Ygfo9re
5qqkTagw1xDEaGEV+AP7r5aAdakZZ+JI6qtVZaRjrciFJsKQGCGtpyZ3AFoBgEt/
uz0rrgyS1Q2UdCC/Dvot6US5q1Q2H1voVXTHUCxL689Yk5a5eo3isLOvHWBCTM8M
1vGLRs/9prGMZXhFty8VavEN6jjoxkLClFnfWYHToJOjZ/KnpOeuZv3xcgguLmy4
WAQataPPffnuHXN86DQTp5q93OEJcjQ01PvCGMmiRbz6ZiSLiy6VrU/RWzGZZPwl
oOXxO07M2L3KeVk9Y0s/z0cgCFH8uapKup1UxJrVF7pAf8zSZV6bh/OUsAXoJZi1
MG+zc7fCJe4pWhFj9dfYDhdmm5qF9VKhp1j3gNA6AZTJRBIw6pQBXAEWaHOeqH/a
oa6swLH4VEgvs4Pws7SQQYdOnPjrPjHPUJ43q4aBhDP+vp1N16J2zlA9q6a8gtfr
Dm8JXyKQ2DmGM3BV/JOO04RPfRVzdF96D5Qhf9bYmbMo4SzmV/U5xL4a5C8QrYIB
PjBVs5i9EyN5k9k3FKLZAnzjOlefvVHsyAdSrISRIDQGrNqhckzRm28pV9Eom/nd
Uvv09TLBbmENkS5YAi9YXhb70FV01D6+dpKuiSGXvGHlxbXzZQhcHmH+uuR1SoV2
PdznIsRTQ9jVOA9wYoPCub1WwMTOT7auz7X5RGfFA9SfhtdhAGC8Zt3Ui/1IBL1G
JcILBmVcRd6cCrLrzhma1XufOxm2I9LIGL8mANWl8xGfymcpaI0Cq52luitaCT6o
m4jYiej86puzoB97DAwvlWYVGZUlRDQ2rueBPUK2iagZuQJukRze5talczhmU4dP
OGZJgLipti4glUJLhLSxaHvJtVJN/8FzN2NHzQe7YDn3rhZXdcboQYzdc9jSS5f1
SrsiyI/MMQuvEfh7Vhq2+NlTwgmIdDtOMM3rhYyrxVB0TfoSTSlGMsK3C6AuTkPy
lOhCwgdsO8pujjZbPx6cp0tJ9Obp19KUHK/LVxz5crjTfmln13oZj/jqgZhkFqLe
0plNKPaURibWFhGFzv5TCD1njWmk807rjXDKdUJePDrumaxEqJR6MzM39QnA4+s3
GzxpdviknsI03NF3ZBrwpJFXP3tkr5JXcQ2a9hVcsyteVDh9VT0a//pHTymKcgBL
QNjCL6AAeFvaOHxDL/CxF1NcJM1I5y9BEwOORwQHTZyNxYM8vlamKOeOGMzQMsB8
MZeH/MxOZzJ8yv2EsicCiFyLKqlMzRGuo7gJKef4Uv9K9WZD6VZZ/cMAYTiCqSFB
NGnJp+Wh8oVN4rSbK6IDDXCbdkUCpv2lEJJacKweW7D6jGyGa5u9BqQxui8SYch2
Ga8Q0Gxn3xEPvsXztsA6zYuWEJdjSnHt6DDDo5TN2MdeQ/ljC08lH/0o8Yt4Hroq
hVgaot+4ZM9cKWYKns1u9z5PUBKg0Vta4sISmaKoffT1uY74vtR8SDw7EUZsQS+H
Ke51wMXJTtJ3E9NhE8FDKKxh8dEOD6juJM7ER+sfMuFCw7tDo9/ElH/qUBiopNk6
mzd1tDz0BQE64F6EYoL6oB6l0RJiZUvSLoRgnuxEmXvjB+hLQoSLkyPzgn974WR0
n1xfhhPQKXv0OM1PIJL7Fyu+NIKNd6bOlMmJft7oKS646AVlMvlK47PPmcO5umwG
NJFINWuTEJAedxhbUjzXpNzwewJnD9waWAyfrOaNLarpggnf8JEK0xj8yJ+jcioL
HdcEeq3meCR2zj9ElC/mRxzjKMAOi/+A40RJr8yzgSVbOcAaJ3VRZDUcMk8WYy9o
`protect END_PROTECTED
