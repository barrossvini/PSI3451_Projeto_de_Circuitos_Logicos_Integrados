`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2CTc1TtKDVSHkgn+8vr6UZvT8DV55uzd6FEJZIRur9AjG8Xwrm/smz6b7s7WyAbn
dEkNL4iyJ92+CLcgAFEe+0DXCBNTWMF9tvVslyZuVTFIJ36iKsIDXxincViAkDBH
BW8FAf29wiKxH2YQh2NO9ID7sw0F4mmzJ6HexfXDbCNmzXYvhhWPPUvJEArmPmsi
1chJdOjXVQtBtjZp3uAIWyGPiwalb0MKfvHmEFB8Mk0eFQoumyhEDqEUaAdeq4wC
kgaoSQFA49bWYkVhkU4xBxHUp/PCShG3yMHXZo70w2EwKjYQ/56LWYyuwBknE+6V
PDlNZoaLwpidyOIsK27j578qkmFeIZJY0vKUy2nBWa5n7Tgwn5jJAF8do+TVl3At
0KP3B3p+Pl93xrbc1MjCjmIOLqFyamwY9oK+wSGKVNyyLgTN0Ibdg5AvTKgDR3cO
d2OryOg9H73BYpltswyucr2Yi64UfmTZVWQy31WUDeuxYoHM3XZXhjhUDleiAWDX
WrgTBKHTqtTMm1XTKYvXC3NmiwOwaaeXiRdrHAOmf2QkSQQSZGAx1aJDRZiVFS6l
2bMgVAtOrmWOPKJnAmQi6VckEVS4luA2J3Rb4W3QkMc=
`protect END_PROTECTED
