`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0QZYMZ3DELXNWkPt0uQMgsZBcHtensmsiJcwpCjQiPV8nU+r256Va86HSKXRI/jm
4aOkcznqPmc/hZxqxAB8OXHkq3+8qsOj/owGF/3My6oyPt55c7XpFN8Yyd3acmKp
+8vN0FaMTTZ0TwBoQtI8CxA8NKiplD8UfFG6JI9Jj0cbVKdPkVxjYTW3lvRrx4gm
qQgWXnNEJTcjRev1uGf+E8i7A3EzCBjWqAOVT/4sJcF/sPNps3wEPUOVOYy3LIBz
NWG9BUmHjhj3uTxQ+9HT6UGmEcRg/Db1Ti4Tk/xzfgwqigPRhCcEWJf6hMe5xds2
cp1c2cED4EhyUgJO2IZRJBggbYCN7OQDg1mBqwyzMPGaXTRiEZcE7/lOov7JTyJR
W39sSEHLnnha2Uq+qiwZ85klEMKLb9fWwqhOK8kJVpSscY6NqU3Ayhb8PSd1+HBF
N2ILlIvIE2077rVf+McKSPAQmGHVDt2HuMmVNaf4pgKbVg2u/Ubh+TmoTFq1en0O
Q9xeenlLnxXuSNQet12SF7FBJr+Avn220XbUF4gAC8aSlhxMsx70ju8TUxiimy97
IjoaWNwVUcDg2awfPacEBUXlqOggScCmYf15gHAFQTPMHfZ5mwlFGNbsnUfuFTiv
I8bmZ5rxgfneqBLMHx1VQgb/AHKz+IOJkaLPKw6VjXugjj07JOQ0DUhkJQBjKJIY
S2tVRY0Gfh/2v0aqx4wlpNvECtWzHsPyFxjgaSnycu59mt4RCvIgCiMNX986DiDK
QWSRaHgNXUAMY8GpgLRJT3hLavaZqbVu8ZSsfY4xYRmI0GamSMAjV9E0Y39i+Ezi
3YDmevlP3m8RdJ56k4x2OnGXPg3szJvqNxRMnXJEo0en67uT2oCiZc4DclzkfQOI
w6uQNDFLYK0tjv4hPJ83Y0+Ytoqoiv0UaNvs/Wlxi6O/B047EDsosgYkARYbXGFx
2Mvlc+3SdlevHJSyIzap5umPzNvPAS3FPmtNRS7gNQa6YfwkRziw9J+JgyscQZXo
NYHHiKL2bJBrJo9D1Jkzna5YwxCN5DsXBVlG/5mxy4RRzX8q8/30C+rS44vJTg9U
MPuj+vmg5BgbHWejc2ULh2Uxrnzbvt5HGVFW0ocvHsWIZwbmpZ2qMUEk2qJnsGWI
zxxQjrtmZq34nmWEjBXEw1I+v1m7q7arXa29XeGYhmYOeGpy9Xh7mu2gWWySoFey
ECO6Dri92EQrEtuLPOjA/RJvlXTCvk4BNyTRWC+0jPr6DN+cdEk5Z6NcCZBpnpYT
h56dX3e30EEuG7AnFoItSnC27kZfhglRdLjJ33Xw8f0zHFym/3I6sPAdw8DofsP1
q5OUccJVYSVJiEiri6RgDI5wTdfUo9WQuYVGOGq/1+Xdz4XDQbLAqvEt3KfQ2PR7
QK2lJbPbMoKGso3iyvIgPMWTjN5a21Dva50siFYbaxTN9mkWl2GSZEB/5EkI6ZFv
yaVG7C0WVhDwCbUBRon2GHHIsHzreY0jVcnqKPwIXy4TJ78rBwnXQP2SGBlzyOAL
i6qIR3kmn/H9sPD0/jfItm6YIlALUtbK1V0na/kqVNCjb5iEBjNZa+YvFgOKTDO4
FUO/lZHc8JSNO3dvW/+poFxEmeB37D0CqolZ/4FDcM2OKFZS6g2rEM+7Li42MJs0
gZYGMuo2DHmWtUfXQkF/XVGzoWOo+NCH+g1pxjXIX2F0/hlYRhFgFvs66WOLFMh2
Ss5S/bIVkwUpsU+OfkAOJ1um6FQ1sMBjfzU0A8tF9BNwPpU+D03h0drB96EQa1sk
FZXZfxwnFoU15dS1wt9dDToJVN45gKHim+6Gv2xyPFs8I7OuqCLQg6OWGtXUGsvx
odxuSrncebkBW7O8nqIGPlrHjgLrx/O8PV1lNOI6oq1A11aDI3ZXv2cZDssTi136
`protect END_PROTECTED
