`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7HdULT/a9g0cZ4xDJNMs1Penf3NBmsNszeoNUAulYwVJ3+AuV8Qq0pDQDAbKWIAe
Vr7acdDi+N6vZBkntlPVZUzLuLsCmnia0/mAsWEsAHukBFLNL9xNUAlfeHISBKdg
IFoQt4zvINxoP5q1sYdXtuVJDtqQ2HB3Hd8iJUDCfVPvqvbLJcmSwMheHIyuDQa8
u49RC/iQRU7MWX6zEehOxsbcEi0fSYz8D45IF+elnVtDs8p3RVVoXI5C14aUcdw/
g8QFk36cnOlR1QiSrfDcgQPRIlvLS9EiKd7+8tlKf4wGWFfhLMg1If9B/JGjw3Ng
XWPLLPCMZEtCXm5z7JbAt16wkotb0s3S+z/Q8SGctvD7g/3x9PBNgh+DMdEH9FWB
QrYDmfp4rAQ7bCyKeecj3hiE/cth/bacp9vJ5n3UdVDJO6QcBHGlyTMSbbpTdyFS
5nPrSm8q38rjFr/1xSMto36cHBNtvn9clqtfsHLaQ2afBA/hA3LXwAkVVuE4s4Bu
INrT7pvuLhlJh241XOydplSoto4vSVTrBVlTnJy1l6AjtXH3MQ+g3NBqu/p5ED0Q
hMM0UscrSveuDeu1ezQWWSmho/sescj3o2MrEFJvJwusATICyXniAdehPwl11SPz
BQljpeADayYmGtiJQeknO5gc7nzZq1wpOqRExXAQgSF7hDx1TgVP75W4cNDRHUsl
VBOwJrUHqtjZHcEGyGO3y9giDm27OLnSyT/bYWIZAZFEIO1eK2OYjb50ujwL1bwI
pF7Rq2f4Qn2fCl193m6nyLKQCehdXuhuUxbdOjgPuUsgf1m8rlPxMLHeo4HR5EGW
iXf5b8fR5EB1jFBe/ljGsCTtYC39i2X+M5np2gtzTp1wqJGf25p3FD2cbJUKqxRH
m4wukGtK4QVEEqWZNvs1asvvnvLl1rEsvYD6A46AHPdADFHCS5FmfsZPAMkcJ8SN
0R0/dQFhUiWm2BzPajQuZp9EoNCNTYOEF8fZcGo1a9tUfHpuUvkyDocxn0Qtwc7+
7kWMHK90OXQAl123GbXlitI+0f0UBjJiH8GwBzulHCTg0DbSCzmHe+A1Zd0WOrat
xGnxkkHkP4k0KcQK+jCIbEKPJSNmOhf8xEIyJ3oQfR7z33oUg3GID4/g3g5z1Ixw
AuXdfCWlT8ZQWcJxUbXeIAiu5ITXMbDf5sBnK6H3QCopwMXRBASDe93FDvUE0NrJ
PvtWrCyNe/YKGcwLEgl3yQT8Hi0nOKq+3cIyowQOcYI2XA2jQwBwvOpcz9DJEkfD
lbpfjAcKNM2G/P+TiKYPbyPkh4uNuP0dXctzcDI5iDynFB6+qG+xxpewNKFdyHIV
USiR4/fg50+rvT9M91o3Wj6RE/R+uns8tFcyd2RhzFcaEHljEc2xBt+XpuXbV0mn
dEXzyV3EMJBkgaJsvfyCHHkstbvEiYaRCW1oZZvDX7m0X0CXMgBS0cADiUdbbBkv
2uPUN46UYmdlXHayykOHKTNNWkCNdVP9TKgfOVL2FLnYzHBF7tBPU9hcwZz9ulFw
GpuG8FNtsDleS36nRA2X2df2hXtYMP4spCEnH9StpwvREQPZxK0wqLRj/BEHB6TB
VRemGsg5XhXItVlQYjHDMrLkVSF3IDPyTyzq13bvwjauE05Jk2htdh464qbHWwqS
bMD+wLIzopI7pBC5nduesAIgHCyI8HymnYPpqR73csBFbSbFE+cPM0KX5z7W9Fs1
zPiEeZ6qfNFlmkJjRUfc0MxGJjxk8rUG6pfd3V09UL1opx0AnvLztwWOqT8r3BsT
zSCsMggGhtO53Ie6ziGp/YglcowOG2i+U1+zWJlm3oP4OW8ejVCnl+/v3p169otC
0rpaqclxh+O2f6Gnn99w9u425jR2L/c60uo8tmyA4yGS2bOfYd7Yw5gKuR+Dm902
XYVp9XNvwmQmy7DaSHAxGrFgjmgvugukjDmViQNKrwql2fxjkJX86BBcVW6MxSt7
jTKEXqMnEzor68qzMmh9R0f2moeJ3QgO74S+TetDqU5WFhznKtWOalMd/8mxT8nf
iK3KSuh7w44vpo9Y5w8HPm+wTf/3Z1q5s/h07tZQWbPaLopVDMPu6VewcqCTJfKv
WanYwI1zhB2vhA8OIqXvcAdzwC+Rhvj/qd0iyIy7YKwtJfLWqYI9GJ7uSd6j2TAO
7ZizkGg3jqKmQe/wJAaXA8GHITBDhy1eCQvU6MR/9pCn7v127clKcPWwYgt48MuS
UjDZMpiUEt3l9MyuWRMcuA2sxlX79CYPmpBDO6X6sF1ZApahf/gKRRV+yucxPeyl
BUkEerOBlTHGbTkO8JPAlF7vCxxwjtK7JISKWG0CjCCQCsIp2f+RYvE+uiRKPcfT
p+7j6gJ/pfo/cPG1IWmQa+VUK8wAtmZYktgUhuN6nWhkVKyU+vCWgjQ69lkx02ma
Hy5YNUPSN4pwwY/GBMH5+0566MLccpFOY9zWr1pNx3/MtdobvV5PQvLgKOjnr787
otSMb1a1zdvIn3FBtxuMx9NSUe04dsPDWD7pYiCUOtJsjO87/Q/L46bLecVyko21
xG6wuFNoWhS8A2HTpCXZhid6VH21chFvXifFbNvvPfcrtjCv3TvQU+DhLa70YG4E
DAe8x9niH5CBmDn0oe3OTjBQpF8QfWiLZlg4c5hFDZXIAARrSHl4D+noN+w0ilpp
95I82iKeI/20+njB6GZevWBxAS1XWb5kFg0ZN96LzxU9JUK65p1DTDbJEb2bppa7
ZUGcJM3vQzT21zzX131GutcyB6uqSclgvCjxyOMltlqHvKXyJPVkN8fWS3z74JYj
gBtoeO7CNzEsQFud51GUw9rDwoc5QU5+y54gejzkAL6jFaFnIIAJm7QDlUu1shjB
lhq9tjji9Cb/jIGVUQ1YITjMMzVJ8b8Hxzeb3vTHa1lCVlnql2F892IqSYp/V9Cr
pm22i9vbih3rV3F93HMNVsm8AbYUQW0f34jiiiOwALmiSIfEKB36AlfsoFHhGaAC
7AYJejM9Wlc1J234t2GrKY6/+swpIfp8p9HhBKGaNbl3BpWIBsqj1uyWo1S/cT18
jn66frIS6VFG9/HePICEZuHOfnuCM2aur1dHbDmpTiECfMj/lFciaMTCwVowUfmE
Fh7xEFFec0wu/38ghbA4AP4QuKPqGPOoaXLCW1z/+6xazx1XJP/YWgITFBVMFO6a
B4qCObVFBJwDKI23Cix84NN4y6/I4at9ef8LFGd49iUjRffRE5dg6/f5t/1Bjfoy
XyUCUCqIZ5bNG/R/HkjlES6tIobcJrAO0Yi7+nIPDhxLNp2DBIHDSU52F5G/de0m
eYhCAjrLNc8T8c1V1jmoYEjONkL882DUtH1UrPGFM/0VGmDlMMiJ/0hSrcTNamjb
j/fg6LsOMp2f3yTGSCA8/7YCz7ho7PBf/90YvUEqysUv8RpEHcHx4hksTpq2Hq9K
2WoahBI3/W9L/n3WjASz6w/JO6Dila01BcDwQavGHZOPxXxYa0WYdgW14QJ/s6rI
ju5uIXSJ3o5Fd65ueCZ1amihN+V3hHUfq8gXEdITtohWBZDsFfs7RjBT2BKbwR28
kim0TS91a5tXeMI0aC/xFbfSEPTRj7o8fgVgl9kZ86kXt6QvfYg+AL88PWFg6Qfm
65sqESaAk4PQETTiCRaqdfXXj7Dz/0puc9doZGjYEvvH6Yr44QyL3XzT9Fy2k86W
Zc7CS5krc7DwYC4wEBg41tEtW7L3loByBOcMiQC8TjEZ5+3dMIxZUPERQAPPR1zE
T4VeC5qD+5ayO3fs71bpkUclotz0CHQHKwc3uqidQIrcOw2WqnujHlpi/VLAOWMC
8xBGn1m7+bu5YZLjfzyFP6iFFXbrai+RGggUj27w8oh8UDoi6vqMPB1HQZriGFRr
tWZKSZKXxDnvZg6f0OJ154SSm2DZQXghJ6rOcuH9UQcqBfwTB9C1ItZ9eE5BoVK7
hZD6VIWnc4GeYDMGlja0xyEIN/y9mgAGqqvL5B8zAuqEcjJ06zpbpKN9emRkuaZr
git8sHd+Oi+hMUc4SG7gTWasoql3K0NsFtRl166Y1SXEgbtnB7meUunc8qugBPZA
OMsriqdHy3NWWBwL46ZNXxxmlGr3S32kX6jjpEVL8yvJ5myT1oVV/QJzMxZjCwnn
I5RhYUWLUdg4lUrPWA92ZFXQMPpJOpl5Obc6DuAcIQnjS+lVLfaYoV46Qi7V520Z
TTI3Mu3kfpwn9fAJWAca80nX/S2tmneS5aV4k7ixstToPol2RiVrC+r5Kqu1uW5O
qjM8TcnCBzrU8sAVUoEcH08bprDXiw3qajSDZtOmWuzGNYfHPpmrDPUMrGipBiei
DcaI5goNJA+A16yLLCLuth7txJv9rlG5CHAypf9DFeZP8DnoA296EdQLZpD/BpwM
GikCbcusZCEkJ+JryFpbuOyWkNTmNC+pGP2aJ9foxTFaROXiq0q4hEgjmkNxCahG
QgZkyjm8SXmKpxqGPjvLzP70sr2/a4f3/L8q1UD+URNGNEPEmSkvnZsEQGPl5Jrd
eblKdR8tVFAMBxI2gk7MVXAI6kLkl2SLidKSt9zK+iyd+SFxDeVkvIPqAi4vmbUg
qTc1chVvNrSNcsxT0Uj1hdgz7cOeDhlrlQdVN9lGeqaLZ0BaIVjvUt20I+p13yB2
XlUtJKooOCGqMvRsEcI7uk6gFdQRx+gJLcryt4S0zrYg4HXD5RgIVFdb+nM7CnWy
PvoPnlfCNHtrQCRW7BsF7ogu0QTBzq/se8VCwjdYPpsLJhuRpm2+uJFK/zini31L
3BDRdYQyVoC+IDimm6tSA3uCmo6kqHVsSu2LmAAGM4hSr3q5ae5axjWpiQw3lK/9
WyKtEEVVqSrx17QhN3rxfN+uNtpt/FqL8zmmziI1luLX+OwXneHHetJD7YzupxQe
3KJstULBfzFZKt5KK1129M2UwdE8QUii5NoX7H9PDvOrnytS0wl/I32g8uRMyFat
tbGMqXoKTSO3nmhmNS/GIGqIsHboLMkqQMxpYkNLJ7zB6Sj1rH4Q20hgvsi7zO15
4ODC5ZuNIszY59ACcEeccfSUbAvq4biuRZ7momNHOroL2p/L0wNBFCq4Cx/1D42i
/KIX5OkGymC+vGVuWBW+csRreJB+8lgYtBDz8EzJm2zw0g6tQPw8GEqEtwPlTD2i
UE36foFTE3EunHaje/ijxRNg7KV+kM7SJKSEhjrp8lTfTU+54ELT0chgStzTHt0G
F6/yZ/jRKlCYfr2vkIn0hefVImu/J8/H1IcZRL2b1WqLflkMbKZsSUGrPDGOzZtQ
dVrzk4/o5NWyINMTeO+bUiYVN6vwn1CPkX30Dx9Pu3qYBVTgR2jE+TURQNLTHRbv
40rgcgDevEspwUh14hDQctfcVATT+VQpVthKT0ERHewCaNq0nExDwAdtFuQd/YK8
owOdvL4aFf+XY5/QmtDlTzOS5eQ9qKZdimhCBjm2JBOT8IMqfEfKvj+mKc1WRhmB
89AOwNmB78OrgzcqF68Pn+n5gXxuOKMjYc+48iYoSmzOhoo6DUAXUiCMUVfQ7Df0
514DLb0EVpGZNEYAdoUizLM1JZ53FaF/QajikKHsmj9pYagaTRKvDiPvcj4O4f2/
tDY9TRzcFeZKPWZIqIGUmKw8gsWv52DocvBTZQ8D7h5Jx+ey27GkBVUPiwm9W+YJ
hz7iLFHJLdfWw+K0f4tb3FcQRhuL2OlyL5b2ELBnYjEGsCg9iaXAYLboI6F6AfLf
t8Jdf0iAbTQHSGkuvIV29rnLAJZq13vGvc8Hp6YwORWRvSboCECYYIazdi6kXll8
DY0gnnbny/C6RWeucSWRwarYQFmIPv388Ul5I+9aNIrEAv/Wf7VwrUxShMJLtgvD
RJN3pmyOHynffXZC45gnlXn1o10PRnmxgKiDjPI1kToWUnwG1IXQ/4U5bgEIxu6L
vJ/V98Bjz58NVobQLi/6CxFuyqC6Q7DcOjJ/OzWQ8XeSKXGm3xXYQcmby11PGhow
uQ06sy5v3QKdHGDdJF8pa2Ryv52JpkNhKi7gNkSdhT3hvc/u5bjmhUnEdPKifa/j
ZxjAC5dfXvcqUTaUI6/8x/7be9uwqz8lguVNe/DdiU/LjxB/68RM/Gc9G6QOQxeT
9RVezqW/s3T0Iw12u+jFGWoZVC7vYxeBd3gf3ap4yBewm5uxG+a4AenctswOMdtn
gyCc7GVyN7LTI0YuzhL8Mdx14q27ed0zfEG9bOtt9OFNoSXRwx4tUPwZ5XWa2hw5
yK0Slue421Kue+FYh3Ggmpu2KTQzDzfMoOpN1gO1gM7wScfSjjV6P6WhhSPh4Qkd
4v7/7KuQXORbM3NXPu8xWWYTe+Yt9tonTUpL0VHOtfhWRIEgFESdczyNL6+j84Kk
TP9XXmEIxOtqJXt6aO+jHIaVHz5UHHXMUFrvsYjtYAXTrcGTUKfuXg9NxtF/rjav
O7JAFfkIWZWLUp4SQ+ghsqliVJrPOqikzt+BJB7sid33Gd57107APH2r/xCT+J6D
6ZRsqMeTcLzfMHzJgwroH5kd+ua7GIA+s2VBtU9iS1hjY814lhbID+QtYD0z/+Fm
FxXRsmWXJ5Pw8X/DJ0uLwBH+pYHzYoH2VhqmQb73TtRF6miDSF2jIfShLwMpOICE
PaETWKqxEJ7+g+xHArheg3p5Jy7jkeYnrgs3i3475YGi6nD5hpCehWs8W9RqI/eD
IiuisDEGASPU8Ovtt2ODijTeIrfBKtX+m109XLSn3KJ+9AbtHigkPwDXh7zPvW39
ckZL8isT+WjDSHqVzK7IhzUf2UNJQPJS3OkvLz5g0K6VEFQHZwxL7vsWfW1yIncS
hxBSwLy26eGokfuFWDlJla6BokoV/gVC7OFOgnhtRjasPSbifXTDcr4mC0EA65HY
xVQEFAugdo4/R0jyFo6WYzB63ejD538mbdbPxeYnIkzenZ/fduNaB9sWBirSiYyq
2p1AOVEklzvdZgPFWTzvWYicRI61g3iF5V7wubH8tFrEH7XC09u1KuJErSjWhXIo
RB9AgMeq3gV3I3y60YKg4OZpJTJ7TNYFVnABd2w9A8SpAVRrciQJ+nGDCzz78lcz
nWJXG89CPCDlYlkhzz4B0Gp3oCwC9z4Bni442koPLNZF7AhOUy2Ei0D2QIyILeKK
eWYrAc162JeFmzTpesHhYoPwMiNpEhs+4TbIHqRSNBrs4ZAgNf1iPVj38Cwr6Aw9
Wr17gEcpqO6u4JIsQE1GYckFLRsVNUbxes+F8sHIy9aB3sPKLKKED4IIDGCekBGc
QI4PEQ19lTu//eKGZ3cKnER+PTKlG5p3XpKBMZUmdXEfje+mz+60XQBGqhvFQ3f4
0DlLLysddxzeOAGKUDFBIRaJgliSAnYoIVxZc6Mzd5Q5Cns3fmBu1B0OhFn+3sLL
DxFWnPOWiDrrfjlaKfpF//xJE+6nC+TQB0LDojCMpoEvUf0IR4XZk+hnGQ//OR30
6kyXb4rmZcxaPIV6stq2i9u4XJlxvTgbx7MeIRIbroA6hgwGtvkxUtUswK/j22F9
E4/Ad5/vnFXfXDvlk2iqJ2o6w3rqmr8oWz3xDm/5mN+uyoDIjqLr5V/EZo/aaU6u
E7dqqGKebjKWXMG3lLJtsljymfw7jib4v6ZvGw1+pJff/M0OSJHB+mDCJRK6lHWh
1F36dXuNv4HwaFtBnhwNKnWQaTVvhfvBcifuE1Lsxc2JYCZF6fAcBoCcAKPG5Otn
+0iyRoEMn0Td9fBgS1Yg5gTIiKjtGYsKn6NQFD7lwBzAdMjc6twmt49NGuKMSCge
kbdcHqhrTDl0S7ha9Ri0FEMkeI9m5raOoRNlviBCrD+2ZzP7+zdwh+mt+Or1sFw5
hsoOSN2Q+2dhQg08xoKp3uUQB7VXOfYctrpSkuAfNncG/lAw9Rh0+QZpcFftWeYp
z7wtUnU5yryqmb6FPQfHSBk66/YanvITATinLB0xVsmwZHQa7N1zS/ZOFgxTQ1AV
3xQMlYtQOegRyxNCOkWdwiayopdWu9XFocFjMolumXn271N/n6FZcORtx/b6lVUf
vpgZUrra6psTLSWGlff1IACkHIknkfHJMoadE+tPX4bp0Of1FqSWyicOfz7skfrj
hVBdDNRmTUQDyRcmkX/c38cBNZeeSXFISF7SnLtDO6Wvjd/L8mTmg5uBZXCNfluc
Jh446vNInDE0P0Wco3m6taKbHhc8eza4zqFdfRm1VXCQRnrgMnl1OxtU/6oTLV9+
Ao6d6de7uUKPZ27FJP9ejCan3g4OOVUMYOLRZuEXAkHiyrS250jF4fw2fhmwIpIB
bO8PxM9HaJ52f3mqlZqdI0uJRxUKVYnBtjyrRVDwR2mAOesMv2dwC5CCOdAHqIgD
qwC6ptI+SSerIfjUjCCeXpovausLMtiJB4XD19YVg+UNhmAjhulhOKhXdeQbI4no
Tqpb2JwKIPfdIHpGeMiu0+qOQYWodlIzOde4RNhCBgLdfVHz2LyOToPh8IBYMM+n
JCZ0QleiTK2KOpHR3KQS/h3DAO5nNse2q4UUdJhbmLkv8472aJ4klnJ9d/zHcFr+
cqg3yvKSoVFdtVPvMx/8KDQPuxjsx0rtFiYoET68b646wC8CS44Ahifsv8ZYDoo4
TYnbdYlwgZIPCqNcGaUQsIJVuIjTFYQF2EuvdahnTfPTnlUzW0BI2BsFufBlnQyz
XTlsc27wc1eBSc1y0v0x4LEB+muULtLCUe1qtAOd4vdaBX6BaHm7x7j97rruEvuB
8IQ5yAKbvOqAMxrtSWPPf8mUAjnPSi10jJySroakC1+D2cyZBNSSSTzU3Q7rRkBx
Eawo+KWuwDXic1G62tXMdS7KwT+j7XkCUR1iyNraWoOyomyEyEf+ADZM1ovkEWvZ
G/fSwXmDCs4uRQS8KYHyJNoPWHadPLB9FTBP5RxbQuQ+hDrgZI1BnwnbohrqYbn7
VsrFDnbqSwcOoO6V4MzoxkCtge2a3UC09EKoB2THD8FQVcDE0RqHX3WFHiSy90VN
QX8XSowzwGtNu3JREjhyZaxh5KOpvhCwRD5lCzp7+auXnQ/EtUi+FIYWctUB+nH5
4yQj6JzqvXCCi05FlhMzpW2IVndkgIJheWvK+bIy53AlrhhvsOuHIVqGEeJTnnb+
MNGyGvJYffptkqzt/Vq1GhnPnrzGWR+FiflkgcATSSSJ+oVGCdRc9BnaeaEaqsOE
zryBz1Q+N1wSQfOpT8jSBMXx28lYzaWmUEDy7GDtCczMJpfkySGQHudFup2JJCQc
7eXZCgkmF98K1CXaAMt8/WZLdcq6kwx/VNRKvNF/IzezIHBxkJVXsqBCKoiBMNWQ
5ew1zmDC33778EbKxDyGXjvIHiqpC/LKBl2MMttoKcXkZvomOKDDb09vbyrvfZlP
eG0rhi6xcsUWEogIlUUeKNmJfjF3vo4BkfeWWi0GjAH2gedT+j1XDfIAVBEKqL3b
FHfbl8g2c48pbnX3gXH+qoH2qtNchixR6aKAEbs722DTco/39BmlY712OchphDPB
YNH8weI/FSX050pmyFUCk/40z1LqTCBIacPfPmJrJrstNUUCnXNYfcSP9ub1f9Pc
rAJXsc0EFnhbwu/TLARApUQlG5x5qhZ9ZtG52roR8LrbhAAEXc7AUcHItyALOOhw
i7T2UHEc9rjlds1y8JOELqfGLIb/IGh+/yZ0DLy5uDiXC2xgQ9tt9NWgnCWw7VEm
UIhZYnGkxDQy0eUp1DsvDXr/W+wmNwiaDIWL0AK+aLtZ5PRxLRVHxDNbJjrFAKbb
q5D2t2kGfI2g9qhJ3dHv08Tvsk6K0va4Lq6LQq2DXy77c/QImxsSxQpI9KZV1xW0
yMdw/cj9Z540cRWdepkGDKdBMvbfeXrVdKH9kHisrTfZxyZXe0G+3eGsb7UQ2stV
4xQtTddqqnuMRbd8qkVxollgnwCrR25A8BJU6xl37TW6IQENn3NdyTvKCQcMsbVe
v1ynmQBxkzTWhJvY2PCekResG30sjktXfpd7rrMem4e6rJO0YFLf1KuuelKJrTn5
gZVW4IN1tAmnXLO/bqGygTJfqTkDQna6YOLoXijZ7YJpjDmxJiJ9m3jTDn3BYM1t
N4LcZ4NHBlWb6puYUrPws+NRAN+T4dciCCcV3Zu6QhOLTUoG3jBm9eDSXxzW/GWK
nowyyA0eoalCKdRv+ja2/Aou20nfOUBL2NSU0OcA+FDNtErEGByxEij+nnVBU1ZZ
yAocvbv5lA/v5OYBnKYSwZvfh6VvJ3thPRocJmraRr5j8Cvmz7ekt4f8vm+joo5H
XRWFHvR1upZCM2ObH0hvR7gauaMO+Ip4qAd+D20uH6qoZL40+2fJSpjJnOVTZ1mJ
Surw5yL/mCAYnP0CVTZKovQZ8qgrpFNXarzBwGCCt8pzkkKWnvc5iCWN+MKKQZw3
37xthlBRyEhMLVi/9/s7JprL/I/9jj8/k7YOKhYtrq+3eG2m4f0nAO88EYrjeMWO
U9jTX4hXAPzHqFpQvBJdZD66DJCBdMLUk7QawUHrKUCRJz+AnSfEsGAOYBoNb6Gn
2V+z6xHfyU3TDF+MmkR5zd5sWkJHdk9HeTMxo8pwYkIGvQoaCRdX1tgEChpkNP+u
zAekhCmlkRrednrLcEn9Gkeh5227H2SJsK4HUim4XHYD1Fi2zbKKLPxlzAlaqd1y
uARyKlaIBWou6gzLTQWm1NFOnMopwAPkAe+gteU5cUh6CsgRUWAL2DvEFpuwDCtS
XfE8xa8/0yQR1Qw+r8zKlc8CMgVMG/YyTb5KbJiB2kzZIsdbZTQ4mJcR3iCF8qf/
0l0DDvr0f0Uzi3JOyJrqyMaJ6+LDF5yyhheaKisP5GTXKMCwEfulSwI4fYeYOc26
+rUoUvH5OjWtPKzpz3QEBg3BtN7/3O8T9Yd039BHV4CaI2wBfPRPQvtV7P0iZyD8
a3/5ElozDkyig67j5S0O0F8Y/4kprC+7tF1ra8aPcBuKv0KchSgpsUirAhuqJmay
fQlcQIKhbrWpZaWYppiPije5dVm10h/8UhYuAtfCHwip2UDHasP3/MuF8+dkRFy5
7alTRZQ3doh1E4JC3958eoc+OgENZJoRnKsckn/TETX+JbtIOV0GNUUTmgkPmBPm
G3f1EwFRiFjmQZstqhcMdG/+E17Evs7JuK2CpzcYySEqv9vuj84YE1wkkqDTMFw6
48nOc7FfeTr+tIe93g7C8VTQm64JLMxCHLcL+VJIoMPxSGpctsPUqT+SOZ+M/bDY
GUC9hAamRZbi1lkCxyGCaBOyCSYjbQz4YVtW2uO+VGv70wedt5PPSebClxUQBXqg
2/9yXwkHgGQWRv+squ3VvHYS8zTN5sKpigJsr+IDBHF/YrOUl/eseCYJ9+fUxZV7
1FEtUkiaCG//JO0sdV29Eo0/Y+/MQQq1m0jfvrprL9nPkzqeJq7tTV2YDkbawEHi
jQiF35F6Nvl2P+tIByQSCGVVgo2KSFtJ6Q7OK4UVP+vvndejRcb3xEhAqwm66QaN
NcExFzkHUkoQIFZGXaGLZbgna1wvLdPwtIcsCqzYMX3QRwLqIl5nAq7oQ+Hmhctv
V/FyrBwMD0mTPO3jv+g1F9kthxFLXftEJ147ei4xpqmyMAQ0kuZciXJQuzsFpg1L
Bh1i76peKT3XdnnhINhcmZjX2usk2EOJCAaMC9RvdUzs753JzZY5w/9Lufn1JTL9
bxYTrQXTNAzvP1Gy2u/uZKy2f7C42lxZlvncf5tpzZn6lIzbkhtCSCpFoCiOObRd
xzHJPmLkasBGwjKSz63Atw/I19j5YJjDdjaJ4NDhW1v+5pbJdB36MCkgoUgPrEYb
XG1FDtMuxn9aupNAZuMro4Hwu0Rdd9F9opQac9bBy8pN6/Uxc/SvdVG2zmDd27fi
njJRHbCUXJxD8PGF1fiDpFVHFwGcLSdLfxZPBh+d5MWAv2OvT/VKGw9xQfAAiYVF
M+chI2yyjZmpJdLVion28sJ/gSAEKzpWVfzHKfWfKsqR2f6LEHQZb/I6zPgTO7IM
4UyCgKkwdW1+XgfQLSqjem2HCPtFDMOkif1UFUJ04bnhBUqCci54CKrAsSq5pfX2
hMjlJNG8Ablx7glRw6L9eiN14jnlH2Brh8tkl9UllDqgTwXZktuCgVJxVmNkxE98
FnRRXmWrGX7PCepmdohVL7Da2FJW395WS3SF4D9NF6VovwKS4MipwNztbU2nJBPp
REvKdhpbVBIONRb4xlJYvNTkjUF95FkM4k7yx1Ixp9P+LxMvoLWaKEuNjl/M6LNz
qYhaerYurF1Ba9dxW3HY3i+1mZ7YpSFJC51kbSa6pvBR0qYL/e2bFRHSOc5kkPgG
9lps3HC4mMq6ZO4sePnGqLM4lxJt0zozynB9FYXxK1JVo2N38bnCpyQenv9S0Zx+
yHayJ5n92a6cRVnwqkNSiAWKwvNNaweEy0itaxhm7ya0a9Hf2ev0Neg2m0CshMVT
7Xk+KqAyF7BNZxpPJyf2E3SXJkUrum4dE68c8Znru0S7UTsdI+69VpkhaFF1e3ad
p/p6U5pD6FO96TEnJwTkZcgkGtkuT5zxA6tHpzKpypIdZqUYPAWW7PLyo3xqRU8I
GvOhHizRTBBEZXtFY9r3VXynSk+BtQ1mnrLlkqGh4vybOvjoOUUhEQdw5R7pLbHy
1dMYrkm9sH9clG0sXOJZWR87YYlePd/PJk2s4IiFQrkFA1a5jjFjyIr1hhcAmM1F
Bp25BtsNc0vH74Im/FT/nJ8Mh6vPOU5NMXHqaHxKcysS83Y2qGqZ7Ox3kKCVnee5
0/ZGQT6S/ntwKk/Si5uG1yWZCBTaQvlcdRXe7M+ZYz4w0qsV59FM/AvwEdHYBNue
sBa16G7pFT2WhrAFuFDUgC/OSAF7oGK0E6su6wds5rg2ZcRibeEqdDsuq0gV3/T2
MgbmO8pmvduXX01yDA29dxgSi65fKN2PfL/Xi52QyvaRSnXcQnR6kEzUEbzSXGUh
TG9iKOwtE2sPwCh8j2nP8x5OkKHqCLtEy8o/w8UWqNq/S2Dh39KZwAWNDU8JMkcs
nUEmYUbam0DiKuPs30hniRC+HRAqszgoY8oZI765l3vWDT9gM3lo/6uPyuM7bz7p
4qM/J9tpigdz1ydyKrtgcFs39MN7fBMMk0ek8NzVHxEh4OG5sAH9qYpej/ZgQbkP
+T84wDy42ZMK96P9WQUsmMRYYAJLGO0bONa/Q4lG/YpTIBJ/2n4mKqgsINUyiXME
f26RLIssFYj2hNDr2KQoF1FlNUIf13boSqRp1uzlmIA9DqyAaS67EUnKMtKi13YC
vsXWB4Wk9skZwoyzas1D2ufs4xHPJi3fLBrCnUrQdZGzLMBVs+jqsH/G0XQLtJDZ
sirLrBWIxsqw+H1rMduxPCNQ2U3F6Gi83L3TAcMSMRN5TZB3cvFWbpnw8mC9e+1I
g43zeRwNPg8HNsJMYy1Ykf4sM9ki0rXVgemkY37fXBfTY8gLf2obRQjCj1Jv/KUg
a1a1wv7ZV0Md+XJK2T3Ri5VFuDobY/l6Nm9YYnOBm4pRDdl9GeM0bRnJHI7KjheF
UQpGA0h5GctmviPKbe7Mmyeau9NowqJ5r/KXJrSNj/83KMjimB8qLoUu7wW+fwfm
5dI+gi4AP6qA0KHudW182dZ6j/0M7IMbEkQpwTGXzOiqDbBR5a6IjDXUPhGXTGRr
iMU//BQUV4S1DgssOwJoVlyfYzEBH2IYeN/j47rWKOqaeBiD90YEK+YaiYOSzmsj
/IzkCD0klTsmApKRZcXyCPLnw4ql24jaW57I7HujM4MOSHdpbBO1lPUmesBd2JSK
BeCliVZKV4YZRfFEG0Jvp2Ua+alBOdAv12XY+202+y37kaSv6Z/sIc85bENgkYqW
6HhnrPX3hn0nUMDnl0ROlAGDQpCGFPt2w56F/wctk+7IuGUO6UwZJWDKRWGESy5j
4jglqYnuFhEW/+uf+qMv0odQ5zh6bihr13EDr4yLVCGDngeeOeelb8g4woNTyfUd
t9n0O0hCW23Q9UqVUhVYf9Qt02wdJ69EtWWHt66B5JUceGXZAxZpEG3cONK2zy4W
9cahXcsoLVcADX5fEBetLaPaJp2ZRoc9GihnVZFXOTIdXdbeIU+uD9gfdk3A1R19
IeqJlGIlLt1njs3BLqaij4VqxtIRahGJl8Lta0TvCmf1kjIhI+iQB4FuaGa15JNC
90bWTKG5W61cYY+lOixQC8W3+9tR54KJl8nipFS337xbshjkMuB+FWd4Cz+zUqIE
5C5BS8lfn1zibJxFOfbWEM69zhs59biIg+EoCCI9oY12896wMbuvFAb8znKX00F+
4vsBsSaO0dmAyTPpGAlK0vR7QlSPthCmcvNOiQOLmkaHi5nzm7pf6FSFM4NjG2CC
zeFESaQPcilCMw2Hm6CTYqWItbdaLjDTKOVXwtKQpY8MuiwgSPq0xP+DNwRNoZ8o
3aja/jZGjiBs6Uo3Q7zUG3qVrszegXACzP5KQtyApZMd6xbIf4nKurMrbP8jS4S8
ehZg2Dn842QJzFh+iLXtvcUVwuwpFYli2EDaSzsQp75ef7+8hNZGAcL6dykC4kXD
LHl8dvKis5myB4lHFlhd4xgmYAjNqmkKUAnt7l/O4DpOIJ31YokRMnw3mWTDu9WO
ewWNVjEB/B3E8Wwn16D+dOFJIUfu0pafcpmGfNP/LedMcUpDdqwlB1D6nVEfGo1+
KyicIKIkOYeGZTpG1F/3XS5zT2QFbXyo9ntg8VDtrLAjvp7dJzN5A14ZbnAx2wmp
lREkmoGHt4ZN9RuBXM51cWrdrJkNx1KrFU8boqGEg4BPD7aMbZaB/8df9W1lSzGN
iLXltRWo5hjtf4JkjOtYdEniyeLdumYnkkuCuNlZTRHZUUdfWi2Wvb2dF6rlTkol
cXW4S0wm5mJSy+0yxdLkgyvy3lPaDCWaRjbrobY3iw1+VY0Fb3kD6PwYoIt8DGuU
ia0H0tFtl8T5y6cprM4uh4VfA2if3Dg13seDJiPX9YfkoXKeg7kD1VW3y/HecajE
ZMo2mQoBaYQJ+yp6s0tnTijoG0XcCHQCXAWSdM+Wd60pTYRQxH6SpCXjnJkvzy8n
fQksnLAstXnIeIMcJ/vZC7O1AcS8Y8RUsJXrOTTNI4AqeBcOGLIalPnQ8necn6LM
pEcnGs0g3/tCQgzepqNh7dbN9wwCBZ1veBfckB0W7iMyvwb0EfblGmAS4gWzlo5G
N+RSsRbWk/x281BWa2u4LJ4REvzxsqPP+Sz6+9Z3i9+w4J5+9SZbd9yAA2Mv7eNY
QCMevr+FDkrHJ0QklCEVazl1x3tWDqR+pqFwLHkwhFYjS63UUlDO6zi1QBC3LUKA
hGNOyNnVogqkdmOrnPS1bZQgrpD0jXGGRWPe355B8PV+8XQhPVjM4kQobj+BLtJ6
3c9ficxjMqA1Luubb/E3KGGw6fzuR806nWv/nIN2VC7Gwv630ckTmKcWDE5NVr4T
C6AXjVeTfc0/7OItRvmzXSlnZPE3Cj8/+yzVwBDMpGmUB/DOr7QIu3JsXisKYnJC
IKfaZJ83YwzcZOrWegk7PrFO3vdzC4lt/ltH4PeTRSBfcVdBJ227l/QHXw41hmLV
fF8O9v3A66O618AORuBm3wCcW8cNi+PdjX9PgNihCf7BY1pUhqV+zICM37HtbrOw
9OAeyHFcKyueMwjjK2mAikP1Im3Eg35GbMt6DPPJfW+AL9ETsJZRcLH19UE32C2U
WCnPjnnsV53PUQSVoWZ9Ge+2VLE64304QfuMbDut8MfZ46jXLNGXOzEWoXhLXbDr
dFJ+rgjlWFOgCvGvThjgwPm1c4gtankNpdi2x440YZWhoTR4FLIIQqmvUA2enuvR
oCpYPJNNIUezXXMOV2lNxZ7Kfv5zNTReCcPNpwKrQa5Tu1WUMQrbJfG15rxrQe8A
0oP/LR4C/KXqVEsBFbMQBSqIusjho3EAsgBXWCAYSzNThfRJqMrxV6dJvQaOr9aO
OLiHKuvc6cnIUrD/DF/CLoot5qZCV7yvpvi9GWvjkT5yTt3YnCh04urchrJL4y01
mQxQIMcejPNd4PGLH02PbGxfiRZ86wToh64xCiwgVJJvY7u4SaS9I7fbYcKKI7A5
L+f4u20G0yPDHxIAQCfmlwk/xp81++B+WzEe+eNJU4QCrIeO8jfAHV4aQI0xvvlZ
fy+4mEt0ft0DTfzvmbOQLIMH0kKH7AAU8MYS7U/FJ82h7ExqqM1Ll6+CZ0lmPZ9R
YkqqNrPgZY9dwARPq3i/LgGUUkgq/DZnVjTCnuuW3qBOvJL1yv7GQTMGWw1G9sVT
D6rSw838Wf58W1jgf2KMwn0JVsPsTpYFDGyPrNlyfHFtmWMm2QS5TcsYEOdg2jVj
l62Ux64ct3r4v3Ix1GV8bvmR6G1iHP4lBUeNVEODWYddsLC9YxfqLmhdLLGN7lun
6u1k/3hl/XqjOUPZm5C6xF/sx60tmBKrlRETSzdKPRVuAFjDy3IOmWNuqUDJ+N1b
XeeUZFQk+95ziTGadp/pYkl2CuGgaJ4AIOdTsr8xCRiF9AOgbsrYDpfco0yrL8PI
W9cZCqCV8Gupys0oa/ogR/RYh6xIozpW9Sll1+dllTmUkqBAKxXd40XqiThC4QKn
pkvYL/CsFuQ4G6nUCXzbwiBfL5EEv+d+fqfcBqiPG4yt+nt9cbVYDtVIib+Be88B
FRGvBxZxAegQ35rL/s8jkT41VnbJpAFPbIaktGIFNv9u+/vQeJAf70hHRGNGPfhT
QEJns8uMT2Vuyw7CkdBdDd6qx1YIXdrHXTcLgES16qXau9jgPLOxst5cGsv1Qmm4
bwnaUgTdTZXxvHVLD5kujC2wCNHm2St23ePEfGgz4504sRSLZDB93n72MVPZ1j7f
yK3nsY0r6xJEUy8wONXZAvzWZQOE/dM2WiuIcQK0QIHsyTwsAAbg5Hx8OfspNFQ0
JZEFBmadTgvjrJoXAeCUKRPNhZlx76hmK3y0GD1sMF+kzTsIaippDFt8x+8FOWp0
ExcS8OmPYjsVFicK6iq8kwlrUwH+ZiUgSIrh8yMYck9QWHtTslli7pNQnNqC2Pw4
wKQtEceJ3YMdFefiNQYDqWdedCC4Clh+vnua564LcMJR6vO40A4SmSPD+wp2EwJg
rNa5qCY8o5zk6xAkcMzh0C2YLptFHYCVsOZGEBDUfX1Lat0Du9jT6t2PQ2kmVS2i
qkldiE5YkMx2m6JRThSMegvz7jr7AADhk2u4mjdHy7BuhGRLnSRYI75S6NWt6TD6
UTWWFTrhupN5InK2B6Nxa9c7s/Ayd7MLl91YM+l9SOrGMg5j65RV1uzhzqjmYOkD
Gh+3nnHsg1kjwoKoQnxDZ9preHZWwVh0e0/NdW0fCKhsz1UT7Ie9CnM3Dnruiy/0
KeweMvuWRLpbyNfaH7soHYgxDnFMJjeiInxS4K6irbldH3RAKuCIJZyL9OVIfsQm
jCI2wVYloT4gAEqLrJJA+HyWqNxOmGxL+PiSf7JC7GOesPvWIvpVp2OdHAygo6+E
z96yVx5qk2TwJJOjGiqrQ3asZEJ4DKeOtGWGR4GIs5YqevLR8rtCWmeJKf4vEBLt
l3CqLDmrdA6vodxq5P4EUJ1HAgUo4vPG9uunVN+aOUYkdGtHdPFV8MaarNWwKyl0
Ieq91ghmX9Yke9T2pl6JGIBB5V1NgUtEn9YLchwozHrh+DwDLxo03utSGySBHL0M
lM1XkUzPeRQWiR6OWvMzOdIlMBTtGBF9+/FyA5P6Ar7kW/BELVvYKaZ+xCyh/K4+
DdbDiLqaZzcRzxD2l4pzhmuQFQo2YNAQ8ZdbIUKTryZlmVYAJ/X3X2HoASBUlSQz
+n1G7o7M65cEi5yJ75fDyDpErJDUGyH2rtYeicIIwXOSpss0Xf0Q9UboxbJErj2e
Y+YB25BWtnOfEEYGBW6//O5bDJwJFrItBbXqMojcqYFwpI/ePh40Ney0YlGGM/ea
9EYLLlM7a19iJ3KOu7Xdk6pzW8HKxcPASWUdHhHBfYWuo4GUhZffNCrycxD5ZchZ
YZyjUHvdZGiASIp3FeXJ+bbx/jvonv5x+izT5BHC+5wy09j3um2kb+jwAaxqtxjZ
Jdi8fssOG8pQsuSHOkkOkXrbvpueEQKbQc6KIMpt8164D7VQxEUm9c6ePcGulhEE
m+k/xu24n0bFTkl9GilMzf9a/lmNb3iL/mdgN7LW7L7D/fk0fH9GRc+EqD7KUx0j
AyR0jjrb9UfRcPYa/cKPuxDFZ5XUAfPT+3J6cODBXXZM1CvjasafgXiIMoHVIeWr
pUM1B7CmCVcXCJ8hdOsdQ9dAaAYQSOxdq0Uzf6f5akN3sjLymhQqZo3K/IyyZTrU
804yAih9ImA3N5ausmUuDu/B6c5C2y3uYqKlpDwcKQ3ufZJAAoB+dusi/remNRfd
hMMrgrulnu+TKukTxTu5kc9klKf1zt+Zo50gLCnmAxTaWYrXKmfLmgUPSRPENa4U
ZsB6DKkNVIUK8iRpmRI2fGJT0Y5m0s/xuV1p5vlky0hwZOq3W7++O89O1jCx2xxe
vFGWTyppkcoYTL56HiQkE8q0xXZmYimru4iyyKctmCsT/9jLYw1cY6RCxfzrUQdv
zQmdUGm0UKSnOYJaWRCA8IlP2q5zrL56amj+NVheM7Lkwq11j2zQ9XOy/OfX0/9/
GwPk6eduq2fohcr3saIjEJ35Y5LHgD6TVTQx3TYycqhSVluF27nT5TBZ+RJjtCgD
VwKwicCGvwr5Os/exeBe3lmy5pjCRF24U8y5NkLGtCggv6GofJmRxL2rex1mbQcR
dMbFA0o+228zcoaUmUyx28/8PLLAdOZuIJtevbbMe4i9B99sp1C+1aO3RlzdruQP
zjQ2zsDpbY8I5iEBdCJNQB90BtgXKuIIJZbivcvC+MJUMTEkMtghoefthYifIIb0
xjqZlt+cwQK6o/mhOpRDA8PYbVgPXRvGt0Jn2tbLBHSaqizs8Yopn0Ih+OAlbgFI
gGquTO+SU+JHbU0gWkHv9K3pLSUkVG6i7CvxyIHlK1N3akW4HXcF6RHQXqhFxS3K
hCffo480EbPEG1IhWVgNWOEwrFgeqRGkwxPMeFbwErypuc85rGQgkCtOkTJPQ4+4
6CWUVwZLs+l503KbEJzVEcW5p/jNa98mQXGJ5FGbZK6guXcbO6q+AqwE3cGPVwk5
L+tVPZbeajKlqvxznX2x9Z2//3na3OzCQc5f2uAwv5Z6Y1YdLghjbrn9r0cFy3Xu
pPHBqQV3GtMvANo9D+3hupVacMK4DeU7/B+bXWwD0bojNB/+K/sn+HBxDTRBmr9d
K7VMS06t3kLbhJ2iBWJdEZX1RDdkxcNw32zWiLuSnbTyw05QMjlftV1SPqhi33R+
46RBN3E2BQ1AOVej1Uve0oZVg7D2/Yg6IlujgrNvoCL+pQ30JdSZdqu08qNj1kWb
bLkYkpyeGBOmBgTsYzm/OSGN5YJeP4Hf2PV/J9qwDP+BQTDMFGhAotVkV/yBrvE5
y6sqOVmim4TKan82kCchWfrip4qzxfBWqR+tIcZ9tjCTowmmXhi6YGLRoD2l3u9C
IL2VjXkzQF/XaXPS1wDvUlmoKmKlJLk/WAQHSBJ8sLFg+MDyxeDYrl4aJ2PYOgeG
n2TCEx80YjbNEHYNoct4iKt1RXA+7ggc4f06pUtn2Wcfo9WkpQdZESFIPrzxb5yR
LKkKMuVQlOva2nO4nnSl4g/qoTK3V0fV7tAhyUabYNV+vcMEnPzKJ8wfGK62d58h
VlmUM29mjuF9IH6NAmEddqRuxr69i22gsO61SSfqAfPfyjT8xCpsG7wm3Rik6T/+
0l772UQwnB5jJRhSAmxMz+Nlk73MB+dJqe2vxJLO09rZaVFFquLo7ZrTXTE/IQXQ
Emp03FLpusD8GxRKaNElX3HbCJce3MjXwzuUwQvhi295HB+l+Ks+e2YN6pIqw60G
D8Ge5UaxZflsThx1xwG8DApKV+bDlOxZQV5OGzi1HGkw5kaQzkeTAzWZprRKlyvk
IlbXPPP6IuPXRelsAYA4lQ4VZS86TCIAGMUroSGiVNPrjhfqdRyDDvz6J2yrNyJy
PAwdE+3JAQtDJI4jRIrdq+cPuQsyC0VljtmKE5N3pF+zJF23RWFKxPvCViBiT1WX
OzpQz9nAUPFB5uQlGqTJWDlOJCz3fuV7Zq8MiHAsRLqxmWIphMvP4gSCrm8RQbbi
WNPEdgBeMOLmqye8thyzGOY3m566Hic6Cc9zk/F9lZkN0AkNb36kPNs8jdgFeWYV
E5I1NihoLmyiYNdjTSHyQltEMLgdxozZ3x9/wlujfN0INSwleH5iNuxubL893mRH
BCYlCftI3JZkwGfWOefPQJQULnzzGsrNfxm4Q147T6vvq/7rZ5vm8ip5MjKiaDLT
v/FkBu2u9p4gbbqnjPx9SVuzsz45q+FkxWzxM33Bw5jL8dFPaNPOP1mKy7e6Umac
CjbaSiWwk8TLQnLLQC9qWSkLaejP3SdR4zFOI1nekqJGYmCWrTiUyiQ7TEQGRkeD
zuHtN4V+iIjuPNy5CG/AtWuHv0RKlZG5AKu2Qz97aJN+j5l2lhIXXtbeRpWolR0o
Eaiq4SYNRcdv/m2zF3QYRbxhL0dd9/IdHGhpJMCUZdBHkK0jlDxYA4DnBYXxh/KD
CoavIQl1luliGWXkMV4swH3vFu8J2lOLFA653IQxOeSDsjUlqdgIdGBaHzPo66Lb
ZzwqnMqtBf8sxkalcUjdZBASIALmF7iLFkA2bVjRuNvJ/VaKSo43OFwGoalM7ONv
51vSSW7HrInsQaBZzydBg6F4GTyvJWPiISxvias3fMo8POOEYFcCnbwZnSTFs14z
GbiRL4fdbMI89S6q+mwT/QV2+mQTJdhHH1+6x7g9P0xQW9ma1WMxna36913GDdu5
VKaURNdOSqA0fr1tsfRb0rWNvGfu3HRU/L3jye6pvhSGyz9RBbHJ3/+8KaczGQTy
eRmLnQqoMtK2SJ0QK9p9zEbQ/5MelZtDxmgCM2JiCu1ByERZAi1V2o3rkvF8ZGbg
OtgmY7nakujs4RnNY7rwFtdAnjjcIW1yR+ynNRDd5L7KWvT4DhYv8BPMThxrDkcY
OHY02pl95Qys7tCYzNS4sTMPveojRqzvX6B4LUm4GrIUvHx8Lt4+XVGcMi7iJgEg
zbc8uPbGja+3XAN/RDRy6YcWDdBAD46d2BC8GGYKFXU7LX5IHkfqnO0pCo4X5hlN
0FC1HFpEhFHa2mZLTq1F3QKm13FOBTBkopAHWDtYy0d4JKlmGq9JuSs3X/sB2Kah
a9/B24WQ05y6tWm00iTL2SL1jAy3Wbo/ZsGowXNtHRQnO7Vw/sc45/e3uA2Dq68J
hkpv3DirMNyu0BDptLI2nLLfNGxHcyz0gmsEbDuQacUhEFDXYrOFAd1IwgwAShMQ
2qrQYeg3gfSxR3SCALtYcRvwhjiajeDlaw2drVHb6tW/m/GlP5GdU++IYpqRrtQJ
tFbPil78SmnCDFv5Jqvd/VLeeUT2RaKA1eO2NJCowCWsY2EscBtUmA/ku3qcHSX4
U5yhNqzq54h6Zuz2lg5yXXcdBISD35uUlbJKIjWgc+zrVkSzq7TwFG6q16WDWHmH
THRtSFuCGctOZuOGfCOaxRtYUgfBRe9G1oTgfWVW6Zqlar+rKuktK32QvF/2VzL/
eRHtzRG3OTIDOgu8tKpgzQW9nnXS6bgTC9xotAMTMS/eUGZ7CnZ3KjyN2zCPNQc6
Ba+LYSoT0Q1Iu+ptKc/2a9Qhy2zmDszpPuhDOu4vJUgPaQyDnr9F89SMcj6YGB/D
tP6JV7hQJ/FtafjZRFYXOOz0E5MgDAypblzFJlPU2HGObA1n19FNxfaBBUS/bT8L
tC1CPHx3SHJq3Brhs+HUHWrFWNtOE1cdeaLjSU6OC3QezymQabnncy5NeBE9VWfr
1UufgBq2qXR0nDDxQHLC5CdnDbUJWfO9skkZkbjGe1HCosJjURauwkDORPOxCKp0
xX23aFu7Ltct61YPcGnXHYMrKrMCbxsX+HzNQ8cs9uFpghYD5BY62uwDz95CsMGY
tcdm8RK8kcwyFxfUoDQ4273yjo9kCM/7VQL+E6XpLgGibgcbHzMZR1snU+s6Gjp+
DP4evzPqMdA8PJsail+COvhA5FtkTRPaZ8RqNpAnUkdqCccbLktJncbFUt1dJ+Np
llgcV0fH8WM4lxBqZVRPBLBhgb+fiUKbx1r/3eDjdUvMSbIc/nvObL50dgbcK6LP
x9vFwZd9J+9QkJFKtwnTfoj3PW5h1hgwB9KQbm9k1TKb2m07n20wC88/nJtfRP/H
1jpzeakLAOTBQLbZPyLMbIStD+9klQtW4IbTQ2LTm4A9Hdg2W5U3mQoG5rbD0vYJ
YA+dukXIGSNBw6pK+IR6U5PfFinI6R+ZX9+UY40tS3T+R4ggv1wXHJdT/0wE6IRC
kYBWjOsafeX8oGCeSukOY2Jk/AGeOKaFpbZbc1f7fXjVGYxuQYcO9zcfQI3o7RNE
hG/Ff8f2BZeoWYgbJjp4p6V3/TxvcAGnSoS/x1ZZZWsQHAxVLG37mMA600YuDqhJ
KAgtAQFCFUvwseAkXnrAe+UB+1g1UAv21N2xZhNspHI376K2zrUYHIitgJIsPgV/
foXlzz4xCxDlsPCxrB9eIBde6eFBpsooxFt7f584iOEVUw38ICPm8o1vPyeiEFmv
lVVh5DHkx/5ziwKrd467kR1CUUylVKeHfoR/9gYY48ohA7GA+IEX2uEVEigy3mxS
vkHVZRKxjbqzdefxoR7kVgzdTTOh2tO7xyWGzIVlSbSd1EQ1sVLbZcqoMEEDd3sl
5SUb4WDmhiXLGVHr33uEwWDNHyBAKkpRDS6kv5ORz8gbjVZ9H0FBhj/7xbJ0/FCQ
7iLLHWUUx9mDAHwsnIZ8ydtp3rC9avUJYYVo+DKBiU9k/ojMGbWU41xhp4B/Uvi6
fgT4vG/j2UKJzgIX98QS8fJCAcZVi4+3aAFMkMDcKokLHcG77jGswManPns6+c3M
Iqz8dNANqgz42gdEJ1XrjMqg2FVQ2MGyqlpz3VfpVWs+/b/QwR41+xCcWyob+msp
ZViLT1rCRIVrceg1FrgwVh4oSqPuHXtyr91Wo3CEwPH0Ygsb4otb4LELrbglkRmO
WehHa9+yv2Aa3TEkNPxd6Mf06ywVtJin3YQcdggMjZBzqi3wTs2tWHcVLrqvroWr
g6BtzbtAEY4sJ1ABgpntSDkn7tx8oH3uwWQeP8nAgu500ebA+uMimPLTR+o+8TSa
z8zefuJUIk85LHJdYdzYo5jnlYLalo2jE5I/41xYLgv8yL/NbdXQMWakZYXeDHWH
wJrXYHDrA5Lu86My3bp1ORy7iGdS6knUTmCO8gIlnJ06SgRF63yY6jvC5wPp9VvM
hIJYtDixjJOZaYWaXyQbo3gUJ5ExcsIYIVCox2ZkpBEi/FkFqExjLp6mknkdGm8w
g6QJ56qv+jN1mUcpsk8KVz4UGIx4UPlLVvp430xgn0ZvASssOY0Y0OBNLfn1pBG0
Xf/Z6buTFTVF/yhslXb4MKqPG1JjSEdndP/l1A89TYTjQEjXGHn/jEidZo8V9VxI
fvr/5AVRHZpZfHIuyggvE0o4+Un6iGD3wPGP+Enmr1z4jsvs375k29QeOi5aTx+4
Zpx3Enh+pij+dF/SQuBGEELQ/18OrMEIO3EMCIaX0gqpv1zBPve+JTGIogndhOt8
u76VqeG/bGiVuV2OB1rza17nRHAcW1Auv9zoIGnWJVYqN8UusZnSrBTLAqt2PnA4
bmaKTkoh9ECWklO7pgk7sPqZaznvOmkl6N7q5+LCyzjWObyqhbBbAxUSxrHoiufs
9d4YXWrb9LpomjurbNLMLZgjCwGC46wRivVaHsVJ0ZdPpTOHaZJd7SQXazvojR6+
KnqhIROCD46H20J4k8ITFnVJOrxR82VsUUfBD9SsaP13/hX/Pu3GVwWaG5CP3vbp
0/6Mm22G3+IFoRaZBjkJlN37vzcKLLf/TrYnk/wHKqLE0SlYN+Q6MNe44cOxcZ0c
vmlfYpwzYeSK9/IA84tcScRXH0x7v7XjWW/NAapDZHkxVPMCSf43794F1n7rFmYL
XXfS2XEkjGF8e8MnJkGtEsy9VtDyUGZ0kWD5+X/XXq36hXYgXQv66ypl6CYKV6Q4
9MpLp3RHPbg89dw8oactOvLW9e3z8UNY9W3nSjyzIVpIgNnilZ9K/qqBvVIjzhOK
e++2s6+8Hg4AuduKQa8TyXN4LlMx9wwpzlAoyVOsNMWlEIcE34zQ3AWgYl3wQZiX
9RSvw3EnKACis7nr8c24VW/bpwcNuXdrWeownPLWYJ8zeomoslaSu3vYAtN6q+53
X/3c2ck8plwTSObVNUANp+mNJLhFLJMBabebdSn/ORBnaRgI5ClKNwYREIyzKnV2
Kybx4OYqripA5wu6sbSUSEjmFInq3IR0+Xxatd2mSwn6VT2Z2sR1jFDxBAa9c15m
ZLdit8EqbwcZ/pjmloU9kJcCZjRc4+Ok/IqFop+VczGdNlgkUFQmLAPCcxKAz9+Q
6014jGYyUrfM5APHfnLc93wIJfP+EIruoQ/9uXqPbbEwNqIgsYfHNI4Fa2Ep8Dn0
0GuED1fKY4l2+7XdDSuQ2RxY6BcPDya/lXfX0Co/y1Jiq2/sRi1pgGqFcLR4FndW
5Ju5D2LZNutkFCxsddSbvEqgnZGHTzBY3XmCcUIQCENRDuAbS3pDhub3Sfd6IqH2
4kJr+VG0INPd/jfs7LoVJ3wm2Y2x7j1qWl4zW4fkuRKSj+mXrtBedfuLuF4wW68d
KilQlSusFnGeKzI71C/VZXZ8uNilyBsYsROWpRUK/k1VGtOl/w+Vb7cYgLZrxAdU
MYesg4JCk19TmRo6UQ0qcVIBWKGLxU2VvGlK38T2Gr/Ty3QCz6ysWARgXxDhsvug
gZiSm1nAAYAF/HyD2V9vPGhKsolVNbmZCFW5ymGxyQQAZxC6H1S6jC8yfJEKeGRl
ALwr9zTi7R5olDyzYxqlpSWwc971KXJMc2n5/yNSY1AaUfThpBA42MxLT+/7ab6U
VPJoOanZTj7DwK0iHdaxEmfmNYn6dGHSOoRcvEIJyyD3YxCa5jnl2zUsYXfNk1y6
ozHxevf1h73ogSldueg6Huq/SScmFpCAOtwdRjR8zDUmYfTPPRuDD4ReI+nJ16qV
mTNL9nlgpm7xkvw5epXPDQMPZAP3J06Qm7HrjT09bpTyOGqBXbv3ANiQv9xXzh2e
VMEQbsWcRrPgiYkJFNf/1RwkQq45r0gBBmLcyTMbxiDTT1X/XmkgNDgX1HlxhAQE
OxWp0KHYxwJvvpJz2o5liMXtG3J07vXXq3NOHjopW9kin2mZjbBSEB6FrIBJRixb
jNB0Y/qm/Q+Ws0lMlCQtGWRzWEqkyellfCP10EJ1o9+HSbBtfEC6NEHUVjg1w3ZP
4TT3Kb+UDztIMDWWAjIg7c6tReHmQOsDp2I4VRoXISzCOgbsxKz/EHVIEF2d2ez7
4yoo6vpxr0FRBEd9QgG+zt0+cbBOqnHuo2xwrtckp/bFMvIXtbKdHNLHzlj0TDtr
2ewXzM12rmgiXZ3x0aO+I5BHPQt3sRt3LDP6Wvk7bXFe+tfAPA8FaDJpWo/v/97j
Kch60+fgCC8IV6fMWkA4bGD00jG8PBii2vQNBORQR0113Ajpf2LD12qbxgLHeUgh
qNJXFObmHE/5Wn+YFwjvAtokJfIGVyoNqJ8DCuzDTjduO0R+tUwRuKElCdEm0Xzb
0GH2P6qF72IuUNB9UrvA9NF3ePqCbxiXbe7e4dVvj9s3QGQbkJt2rcy45lgrgnVf
5HsNjcatTcmiDQlnSQCJoyINBe57WjENhUS7M+OI5ltVcXbF0KDlC4/4lCxVDpxi
qhYXYsNojVP8R625gl5Ls/jx+/gogB8hfT3uJqNi7ASOv9wyeJTkymCF65TYbsSk
JPJvB43w3Q8H2ilXuZ0tmNDzwch2OHQvo9cSkVgJcEttatreYh8u6OwVEeoveQW4
XOm2/VEB4GDaseb75T4VFIYES72XvXQkStXD25ZI9BDCxeJKc1ZUJMb/w2VvIVfw
6rU6nK8APd8xhClfzds8LgfUstUg3XIzlFQu1lkY0+OzePuVyt9qx3KGJy/ArXCR
SZcVHt86j3G0XBMG3nsROSFhc5PDRaRMmL90jzj+U3YmOMsT68hxfpZXDMAY1bis
zIGNGZ5bgKUSNuMVUNH47PZr1KsYojzf/4KvKrY6JK/hiOZug5kQLBfb/jws/OIz
uk5a9ZxzKO+xAlddKzcpbKAwmbAiEoYLsGiRdLW6qj0w8+g2QGioBoDu95x8tGxS
z17hf/XamFtHfIoI8l0Ck1ZlCCh0Zp+o57lpK/68i5E8RxbbB9g4adIknJm7G/fF
MlGACwxPzLqP1b/1YCfhEWccfWmBCDoHAnyRGDNTphEIs7FLMK0cVBd4lu9hE3mI
ypG0iwEO6BkNlE+DbBMGAPbVyWAXml+1rsC2gvYpLuP9tfKHyNF2l0aq5kH4kyLS
eO79sJDtcu1iobUIuLMpK/wKgvEfuFgn+/zZSzTzF1i8uVXBAbsUqNMDn1VOcauu
te6kiFCrdq87bK7rdOftnGkr7amJhCWSy6AtnBOB4IKGDwgyayGHgzBQYhbLhlBb
YrrqZw5cutmWrp36iIFrGPzuk0vwkZaOekqNY4T1r7dqxRSyCer0LXdiKFqH5c3F
Yg5oPXEwTs4wXzqzltU6rWlwwbD6x9fyR/9mcp0zmjtLL0lILqvkOa6goTx6s9Ur
qjyGzppB7QPD2psWWErXKLN35QmScfzJHNq2sVF1tEvmkXkcncS4S9YfX4N+hk5j
84prWXm1JbvxQLLqVjN7sgNxHckeuvROjU/Aa5YR0q3kL0a9sXn+e4v6dQbzSIsA
WNAvgq4mz5HmU38DwIxhiN+1HZusXe/fm8R2CNgReqlZLmUrqyNu/wkVeB05+V91
xwnticITjptZ9GQ/nzb89ebsZnran/T/MV54cOu2dIcQgkqTtcF19yP2Ydc72e2d
S4+iyORYN2o3iP4BoQi4y2jxRqLRH8wBUKEl6n30cNJhdXJsITblpgwVLCawsL35
5qGM+FNq7MJieMc93C+7M6fKq7TwRKFW0olAMPi+txKxDPKdS/RdJYSxbw8JX7zT
SDMUxQf/Di+HVKNFPw0si6iWAb6skhJfntQmPUVNIUFsxcKytDYi2FRLrn2WLiT5
fjE4LJ8PanmP/7pvXF8x9sG8xvHk/b+6+3QrVUeqBeN3NLmL6uBONmisw+wyGkLh
x5roybNbC6VSiAi2JZuuHEwuUaPo9FRhNkLKGeusVu+XZsSK1UWQLSUV2SF0OYkn
6D2yd4LZTTnvuPw/ovMkPOh6VOaiN+CdWvWyXMk+Q3p98BQ3NyUU76yyPJyycfQd
7YS6xRyg6Jd8hDzAQMOidDa8SE1ldH54zFNVZ+/oMI7oAdCPBrr4GsHUlc9ggTDK
drv/1jBCdaWex0yRIdVMooBIm/wb0ndcQZzBd4sHJSuQZCx94fuQYkYL+09r6o1K
Oom4cLgcwRUIQGWgEjSPrxpzZSzwVwm46Z3Pbg9NPaQL87kEGlh8EqFBgQ77JUhP
XDTmNhT803imkhegBCHjA3CDlrKB6Vs4x3JMFaQq/PurgKL2F6nIAmCN5wDJh4i/
DoU/ylCN2L8qU6IkbqrCCDqhlrf466NU5mm0cEfFNtW66RH8ZRDDSTwz66suZXRC
e7IVWcB/TQhJdc7B54LDiSWQDw2SM+DUauBfGEGmdWjiFYuDdzoD4g+nk8UsBryX
oPUBqlCFyI9iPtBDpvMHgJiRDPKRYrXrWtwBSlvOaBoaQuDE2eiVJ969wMZZf0Ke
4wUTRtdrN8Ys4hESC3yJfHjIRSAoVZD+KWWJt1Ao1VUaZIMotKfj0JaFMY8+Ljas
RWywh/BDHYJ3xZUiQY6o71jTN3Pn8ZPDOFwBF1Dgw4o3EuDL+lmR9QI405OVq8C5
ohSi47kFUaSxsrNk0Q0fx+VubE0FkBnGYEhwDKy8f3mjcCzBkZEDZW0V0GG644VH
XwlLtOFxs7XHyfEcQXZ2IIGDoDtGQfd692kcCRAMS1+ImMXt111AL2R/IK/UQjC8
2spcoRU6xcbAn8zX/Q5VvpWQl63/UsQAGcXKcxMuf7rWaEc83DU+KMgZ9UHgqm40
+9ZiASzyIHABnncNSh04LUhIapZrSmVHB2TZDY3KCnVxVw2CaP/t9Z51Tz6/rK7x
LosWD9b2++DdkaqHCXgK6C/7D6ErAyZE7Yhy5zrkoEHodredERtnVnvRnVctdBv/
91xUqLYbS1S7hSmEUrE6IKWiQQ1Qpu5DfqWCzpc879LSjoKyrwDNQoVxOlpzEfHM
5t6muG4g/3pdJZuY8hAht/JrvIJT3QNDh8C+p5ktoLfmHIci6sijZy6867zmxnk3
XiH2z1KJXNmlcoJfuWEuPvWPDh7uUIU7gsfUIn2DWvbxWdtefS/f3k1uAywdVkSF
PKAgvHQbPsmGHT1tBVXSzw79b/snTJY4LJB4/oJmJmdwie1vm6TwxIkBR3jfH4/l
+OXjF0sHxBixiNO5/UJLmfbcZvmIz9j0q3ji7GsiI+5XIBLP+m7j8+vCewH8A2y+
11/9tXh53FFRDUfAbTtdKo47+eYlXH1hwewpTrJUXtOTuJCP7CfW7Q6ZiGpz6hNl
g6qa2Xcsynl8t5AhPP3+k89jHJ1vdMcfva6S9wjbMCyWuE2EOrj+8wSLf2vlM8OS
agU2QwqpMDe+hzn7G12xr2Tl5rIRrRQFTFrEFxTkBlL6i03rs/SireZmWvFZ8Kof
nBj4Gba5nn6bO/Ixog8THhRUmVeQMnNYgkXfo3rN/RPUDJs5mA9IdhYHElIcdlEm
KYdsZiXdVsmbmsl/UiXlg2Z1syZ8HrMMLE/XsMxhCeGmsEkn5oLvKWcs7XueGrhQ
4ZCPEholetJIcnAuRappXxf3HC3vspUMUZliP4rXhcQY3yjmBeSD4Myc99W5tYrL
Sf9uLRQ76lCoR4Ak8XDsucxqBXEjEk7qRjyl6XIzLif+yl1zdYfW1rrl/n+NsnMB
WYyur2znvcimMCZikNmDmGb8DmkPxu3wnSzqTKxtOexkgcUtyNOVOTmTXevMq53t
MKMpuCy68/Lzi7iBwV5qKJIX6oAICdRxiVx7HXBySDsQLAUqQ/u24rN+G1+UdbKG
kmRMuu8ZL5B/lp4OdwEUjkHwonA2m5OIDzmF8aGji7bOXJ+rgQPmWc40jrGgFOTB
0Ev7ZjcEnqZs+MvAxFxGYDI549xS97tjed/MmrI8QkXfkwUJkaUqjIhOSHFu75Xj
rep14EYI2qAzfV46wtPSfdHGFwyy09C0lCysqnY1LQE6WDYmZyMqRQj1qtNkpVOi
aovVibS9WYPT9+QYzuetVr8cgUXnVqttGefT8ubxbkJNTeOsvq0EQSfflt8AsySO
7gQuGi8N/VsMHIfzaYDiloyKiPoZ9PZ1oF+dKdq1+6KN9kL2bMxttgGfVA8rxf2o
EGzi4KoFl9eaKzjySuBQnEAavOCn6WiyjXMGY8dEQMDNsAl43FzL55p3RJAQqH+v
wemjJN1B976knKIeBiJQ3G7grGdKg1kYSSKPpCWPgwqHq32gGyDbjLEqyK61M2EX
jR73a8BGeh2hdtDAaEm9XeilsZdvIUxFomgxlWTGmnlvsluBcpaqmirT7UX6NQjX
GqQhOHLGory+952BiML+UakOKPTmub083jyLsUvFiyex5iKWwVche1dl8ZaakU45
wbsRMZ4lQk1dXbSB+0SWDYHT2P9vowjp6fA3kK7XisZ1tEcGDGjC/f9zSxLDzDE1
4m1cM9gjJoh+K1BWHGckQNs1JKvB1vAhr7EIg5LfQ0uECEk7//erQxTQgPN0cZqF
R9nBU18DhT8iQNrrkXy2NvrXxC3YqGz14/Q8QryjRIATQ4eVKhU1Jz4vg+3I5AgG
NKF+wi4DtdnNRFE5cRPfYBEosr0RFJxjdkw+0SAjE77lO9DQ8ZZtY5dEaom4qp90
d6aYynTF+djl56aIoPy+WIA1QcuMxLw5Jb/y8L2tien8dl3HIGlZiQ8mjVFbYYQn
voB+SSKmq45oqAqNvhxvXNINTp2R66jKrWS1eFPwYClTYMXDf/KxcYkum5obLjj+
HFeXZnILpaQAK5213slF5RgOlf6OaPcfRg9o0/QNrF993dRTlfWpK8F8r4gdLic5
WpwV9oyHHvu6HF6JTZu8ibjmZdlHK4/gtoJmKnuKSJ13zUCIanpbcJOaRKL1MNR9
Wn2S1Ji+oXxsofXaZ4S3xgkyOO3PL0Z6FC+nEvK+n3k6L9BfUz93jsBAXLf8YeVD
oiHzpIrhmVQZCQgq4GG5zPatILQif+iJbsD+i99tsya+phgpUxQzUB19mWUmHQqW
SACicDYMkHFuCvyl5Be3o+tAWELiXH9uZGbBw4JQ+D+aw6U21qrNB84MdBlS1LH5
TPbiTePpgHKx5swfyBQlQ3t6K8kV6h3LCaVfC3+zpIu2vkfRvfGLOzV5oE0nVmYb
whfOs1EdTbUTMPa1u43121xCF6haYPsVI78Y6AoyNq48rZ0zLITDNKp7BvZl9ZGP
8g4TWSg+rzZzqJPSmqk4Sd7WlW6IpIXb2lLpgsxsMOqriJXbshkr2ocVa4QDXlKe
1QC8VTz4+sEGctFJVMvtIU7DqstpcxALngww8Z3po8zUqUoOkHKP9W4OASkB7ZlU
mS47QJhXNesrPjRLPIi1PctyW9SBPpE0cFYyD7+S1ORen3dRrIoMSrzRj7Ntx88Z
zf+YtjAghCLF7IUUOMlwAq+dxnV6qRBm2xJ0dZBsOkpUxhcFwaftr8OeXMzyh7BX
Rahurq4TN84TRY/NOa1T8OtSGNSnV2U+Ub1MGjvM5hU09brFA4q6EjHdvaGItf7b
cj2TNvF5ORNTOwi0OjoW8Ylpdb+gLWEeYZcbFaVimStiLfQEqE89Z9vsUbdRl6YN
SvnPKUaLUCgEC3nUObwSKCbZjYCCfPGfpdwHGkAhYmyLj3THajHWHn585JhzECz6
KaAOvrEDwnSNHB2BtHuGnQeKJ45f8L2iFFAw1vFbM8yaBoZVRis5DlK5jfr7ItCW
YaKIQ5pwwmr8iMiD8kRV1/meqgnzXANyDxzj+gK9qH7/3H2J2Sm9GqbpCPlM70sO
A33gHxuplr2mooZKnDAeIxDzi6/VfHm/7KpjH+ZNhfIwsHpFgD92fYOHU3z/0tOU
zKdlGHp3ngsHWfhyMsSfIMx4rxeNF4bsnABdv5p6xHOX/ShkcB6ucVn1/JCTKqf/
zAHkDvfhrS8Y74z1gRswgR+33v6Zt0x/OVpi3ZG0NcfDTLrmQimnFhvKd82RG8Kk
XNzja8Z/pkF23a2hGLl2zuTeUNs36kxIWnOBnxJylwXxe+xWqmuexc2TZ7WTO88M
378XKWI0nSAZwpEckKOTKStrG0V3YJSZ/R5MqW16Ish8swHCoU6XzB+b9F0XUVI3
KQgs73l3Fp5Ikhn/6f8tYCVq7vXgGhl6qNHqMwbpopoIbNnjaW/IM4aboO2SISBU
m5I6ZMYQ4PvhZNPS9t/Chf6LKuLHii/xufMBRQk+atNIvRLEgDSiewGmTTKxkQrX
6QMxaZjByscnKhlMc9FGGWrvhsqRdG4eBzOBR4DgD4HeD5pFv6iJEXvwW4DUrhEw
+8eojaJC7C3jaXHdFSOv0EDVFibYtLEqH3t9YRToblcJscVzHFYEf4EPgDBs10ZX
SMu8E+h5jSeZEtwA4zHRhmkUfkZ7tzn3H//MEqkgVkC6Amkka5TMF2UsW5Mph08E
ijoq03EN7FI4i7wUtXJzofVf7qqUh6sGO4MCgLryynrX9Fyj4jHLgbGO/fPE352g
XzYG0Qw9T7jViZ9cUoGmWMVfDo7JVPidurafmePa/was0gaUGSXkxMT8JuM/zdh3
9f7VrT2hRtso3ESmXn3xCgK6/OAD3ekzaTgQgKkQFKrTlCznIaJWnE3YDkI7YP+w
+JG04K+Os4t4arhN6Iu51zp4uKmX7eASZ4KflWI2kpJtEbifALKZXQ7VVEvIdIW9
dAxhhD9pcwWFg4j5PLSzQv6/giCPjq3vmyk/hQSULfFleMCg40dG2z5l3nT9L8Zm
xIs7/uabVU0nGjBskkzRDU27OU3o4fg3YY1nkRMMKBeQFnHyV5k6VQ0kU5wqQaFw
9Am6OApqBCe1Lyfoz4OyvP7PI0P05RKVKkfxdIxMbJqBPtt6cuTdiHe5hul4r75o
+NVgyV7umL5b2wvLYPj4PhBhASpwwHPext+0n0fnvy9rWZa1PQuNXlRh7qkMeVG5
GCWqFhEmRTWq3XDqsMp2wCvTmPFDkjA09Jn1rxxGPFX3TrK2rt9iJuib4Hdnb2Sk
sZlXLUR7lFvWvb7gSeyfF325ESYwrPSC3eXkkWv/5pWDhtwlEQQ7fZMGqXqiFLQ6
TVtX6hMmDqbCna2pTXC6XrhYCtzpcZYASG/96KRSF0vB2dy2XwiuYndxk9YnmYTo
EfVV2dqWbx1V76v2l4YQvbJp9i3EOY9kroFfbtubEdutF9JO3DAijYlKHaQplBqx
kKZe+cjaKXc8Lhod3ZQju5ARPGx50wvcAFrwT0tt2jrLqrybJaJV+l6zh9Me4EZw
LYRT5ZW/T2jDWWE4k+0e/agl99d46pxGG3CzDchfpMP9pF+KNIayxMsmKTNFLLw8
8L7DHh+uGhJ5/ZMeQGBlE7sZB8+oftm2N9XEdDuP6ztN9a5ig0eXEotRv+KbptPT
LR+Rd8Rs8RehaZZUDPfMeYjn5Cyn0c9X/Bj68HotR4tpeJqc2OwFJgUq3UK+kzOT
OjS5V30C0ri0DPKnShhk5GThUkKi4Nz22tWYKkcNceaOee9aUCd7OzTOSaKoFNIL
M9L2h1IaTaFAfmnU+m5yNAZT/s08or/F1r7/WsO2XYlIFdgCG6bLILedqqwkcCMG
jE3ueNcBWYbUXd989e2yfFpEmXwS3FRnqB21tvX5aCR3Y33VfZmnFInhGC2Y5qu9
0eya6AvbZDgm0W+LttvZOsqzx63Hi2QjoHq9JwjmMwXRwcIYs45CgZxdrIlinO70
wx7ZaLDHBRpVb03f9+plnR0tw5imcK9Fi4lFu3au5voPFBGLBbgN4pm58AO9qjSQ
QYe5Rt6n0VRWLfdxwknVDNxhIwwSCrk3PHDEAGz0pxLFaPsE3eRMvtyYwPw/+udd
ZnlJZPYYRUakpbH4WCa5PWiEogaWZmDun6lnb6ROoDHxOraA9OaDc+UoqxBf+0jZ
9brZBTT2/tnFnbfds4rZe9ptovAJipPMKqifAARwGutvdxGsExROuOwKvLvinoD4
wd/ciYQWUspbQ3VxGB1EOWpl6WfD1p6jpjg1G6cmO1aHZ/+JLobCs0pJ0MWDsHmN
pdDXUKQUgMRbMvF+Erb1b8DfJdX4AcMLb3jOn1OE062inU2gZsDULZ7oZHq+4/DN
qyjdTxD3xsDKz+ORjBvCKEd9T4S7dc0/9ye2rAZhYVOYZNEM7nLFIhVf2fiUVn/f
i63o59+HCB39U1xM6OBNujkHVwFki8+MayAE6il3/84526AkAUI4KCWKTTc48sj3
a2vajEhn+Hdz0LigZUMZqb4Fq61fhCHRis694kIHRSazecSqq4QQsAuPsRfg2sOF
E7gSTkzJ2wsZUZmDbLwu+wBDynS8M4B4Jc9HqpM6yzSylQwI4MnCQH5t3N82wnaU
1Dw8HbE3cwJeItjvUv5TQS5oq9Yy6gw5KU99484/f5eyHxXkSVElr7jzXTXU8NEL
0arSDPZboR8itho6AmuVJl0/P/WiPj+ECMtL+LQVE7/VF7gKMm+B+iegQiitfG9u
Nb8TiVV12k+xkKCPa4DNlAXLMnGHYHWY9eeoJB0tPsf+3vu101EcUa6lWuaoj0cd
ADGkUAxB3qTBnQecfafurkqg2Yy/6h5IiXKJOGZWnnvOZGiiXxO6+dL06tzzXA+Q
DOz8FLKVRDvOB4Twjl2yUQKtJgtb37nWWpw5zu51e6hMJZ1oIonGg9//pmyoTm9K
PJo88Sa7oX5TIN7ILQjOXldQWxEZZD8In/06GvkPqP2LFZV7fVltHptWWnpAVUdv
ObuWHHAE0rLd0U6MqeVm2IJK+eST8rFPyc3se5GpFzUlC8g5ZHChdUOFzz5ZTKXV
3Sjh1AJ0LJByOyef866PDBhkoEydFOYkCFJfkYGr4QxIhGnqX3ZiD+kbj9qbGVIc
lsTW2MsL09vvZZrvCSv+3q7KHdNK0z4mbZF/ALDpu4D+xVSzQL22IFghEM+jNw1l
b6wjHTptcd34S5hwQta5ZnF/bJ1VQ8APhT33P3w/RDNXPrP0nn1C/tmkuoaTg8aa
bLiSrYT3ANg8EtPTSI1NUlCVQ5imcBuDCPSh/HCfd1ztgwTvGthFKli9wzi0dOkZ
fQXDq38/9HUFKWVMd7DFpbuOcjqfvxoIujoSR3s4+dGwJ1KoRTnCTHJu3FBxlwnm
o3ZR0eViLjo6rShsYuj+507DNH1AEBQvKfjzTY/tr4ruzox4YedIP8pA8jP1ozY1
U7YMrWEsb5+5VSx8gH8nQ3pOJLcRyZzajDtGOVRuE+j4YrhDlbtn9vK0rMPfp8r+
RAq3pZVlRnwlQGRSDpIK+7/mzhdnEPSDmr63wJjPY3rJ6XL2JOHhNdr8rGPMY7Od
b+YGo9vIYS9YiT01DDLfaImueL/z4Wrc5WqJRA1/gAs0FPkcuGqr7VxpxiznV6QO
gKgKgl1dOldERtV7Tzdge6Lc7aiyszKJwuKJ6qo2iY2oFb0JujVJsLZt3Yh5bRVe
HDG3fScUGRSPfVblSqVPCEy10dP/RQa/8YlONV8e5XDSsiCvb7qWE3M70suZ/m41
RTbRJ5KIobUR5QcNd+bN9OAy8rHfVuoWQGAHWj4I7CMz9v3brrYkEkvE2IZZ6jUH
SgtSAZmPVhNUP0irk4gihWHjcHEQnIfY2teE79r/PFr8p90M+O9+QObvzl7VI8DB
buS3HzUF/kap4eenEIie9mqOu7Nfp+JuI5bxhLs0XhNdEmbpY67W29wQLRxhg8R0
Xy7ABXaHkmiGFJrLHugHL5A+6kjbaZmf0wK8QsD7+dcYjB20LkKoIWYgo2tV9tbN
b0WUxlH1GVkW81VU7QnrtBlmjexCKZFmPa4Ttcb8/aSttr8j1UM3HEZYxnJyRMQ6
nYNRSj9K8CBKN+W0nGWBZ0YDtV8PK0sSQo6OI62lZinHpVDUVCtgzILZP0ASQ8p7
NW/qufnohciyoK+2awfAIEoGlSCk2lD9RplgsCPqziAKqJauIXM3bubcjqqGgAOr
osGO+r/joXaatkhCRpX6Nse8S54lHc1rHhIuxl6VqbZ7kuawEkHvLdEjm+5Vwzsb
2klumj35NDb6wqr/IRY79jrDmu0a7rHDyd6t1HsMMBYQOU3BvbsQVI782zIL4c+Q
GoASH0InA4dZiSW1F30eeO8y5G+i6JyIzSbgPNgBWE/2b2ta+V0LoGqhlCTX0MV5
yNYVJ6MM5KmLbsVr7mPHtYoz112ZyHUtKgtImHp6W835nzpPf5OCi2bv6aEWAOVy
Z5gwUKawJvMHe9Q0w+w4j3v0NBU4lG0cHE+vjJNwiUgNGaUIyn6Y0vd8a3daAqZl
QzkGeQ+LR0Yozst9AnzN77AEkeSi27/x4fMA9bgNuXfkQNkljaD8B1iBBXBEHtWK
+a6FupXupiNzg9utOSjaPHxfxcTONIsS9E6dLVP8GTSkN1z9Xd14M19pdb8jqawZ
HKvNEvoqqcmSQ9XgCI3RqFu+9x6riklIisgj/S1jS4qybko8SRsN3j9f9qQ0uclo
PjvC9rvVqXnQlrHpNvxuvmagpDRMMDp2mosKdXzfCPyqLWthpDbP6K3rLoQDk7QV
3vfLMCJCcTK6X6OcXnPr7KS92ffxuU5ehrFSTCgr0iWohhCC4bY3Tu0cA0zKamq+
1Bbygxq7U88VyeO5c2PkR78xCFm3cyis2y/AAmsk8sUmMbbPwaf8eKZq3CHN3BTS
Or0DdMds/3c/mCkzMdncIP3FM4Mw9Ayu+NwAwvlSG02xe1p5kDvCvxj5mwLAYwO3
eGLuR9Y3EvYmQEVVWl9x9K9MC5h1561Gamlj6K3kBHkpHiUVmWlB0Yw+GCclzEzx
okpPc3GqjxrAac9FuqJ7gW1q3cWlThADNg0qlQalPZlzBD4Jily0t9HGz60BlHlH
oRagEP3kD3xdG/o96ip+vt3WoF90hKMpSzlqjT5uXnwJBJsp+e4qH5txEA84s2fT
HBjqvQm0iXZokYRhOEqqXbuMG/F+iTjCmmOV4sKJhhnTlx7E9uBFyxQMDRHzbjJG
AINoX/8WuBMwmuMo3xN1QpgMGTAJvg2PIpDn7kcw3aCt+3fiEgFHe7A75zRyTTZX
fFI4HRBdCISAR8BsPHV+bqwSMcS7IU8ceumIuBIdhS3uf0OdwouZvGzpIOcps4ln
J/ECUWU4eicVcfJD0LyiEDnO1fYrf5EnUlbLF+BANiJi6TfkWz761GVW1cxKxBE3
iMQ37zJL7QRsujXTNon7Uh6kKaDcBiw9RDq5k8uqCusrDWGnEwHVbFL/+GE8MNxH
OL1zDMuGvFLJvlH24phrCqxN05T0ana3Mof/kNUVEC3fUMo4j0TXvM2Bd7HlxH9Z
gJQ3Y2BR+hTwfU+rfh2rewizB2MkbSk+SM2LaO9MmhvNpuXxH+12PHPrWv8S3Y8/
D5WkV/YChcwLMCQffdUBnIs/5wlazrlxFmnhnkR32mc62fLzHHqcn7rYeTBx31/l
ZnmIOlxIUZbUo2YVxVcaDu2IKe8vJhFLzPy6moI1fzgvUBEvjYn2vKR8NASJ+Jrn
SYBsvaKTx6Az8pyNIdjbRZtfQXFAZuS4Gk1Lyx59zhwGVZI3unJeKQ4V2SECxbzv
9u481a6DjJX+ZwFbsb0nzNbHkmoKWkXnm5SjlBLpPf2PQqYPNllwzx2uX7P3L6lP
+JVEZv9JGUxYnLiPqt5uods6A7399ofAnxQOn5h9WBlabA9TBbhyih2NO4ua3jTd
8wW8cD9/Yp9F62qO99+2ngkJim3qzGJFaS+FuEL2jwg1g3ACwAvTzjft+770jhxR
eAj1S8qgu+XEZ+8/KGeyvDp4ffVp16Hwcm84wh2mNeyJMv0uumiDtyOHB5CrNJxO
1XSfJ3FbreRGlx8dGakLgaPfxmHu/nZffm7ySRxMBkjDr052kHFigV+F7YMDVicP
mVEqSiaYkXq8JzpCf4jEwzkyv44uOvTOpmFPatO9+Z+3RdzBMb1PaPGiINS1DI0i
p1D3OHEkZw9jFfOjrY9DUSX7tLxFPd8QRevRshpfFuHhsPFM8HfUrDPSUW0B6NLM
UBNIdSXZdafkKTFY1rJzJusYlBj5XprwG0+MStyfdmb5Bdi1Wj7tBbToY6gHn5UV
hCkFo0PfARJOlrlLBbkL2MC076zJJv8XIaol1sbZzvF6MjYuj3eH7gc4F5bXtpaw
q2mjxibeWDNS5uVVspsnvx/q4+WBo3jXY7qChFK8/2deCUDMVS7Pfwic0LPgIyXz
6pskFsj/uzXQ1FDvl6E6LU/+L3LtKf9mSDBxy0SKR4eJbk1ethuyy7EjN+iPUO6S
T/Wo6tyAkhmuXN3api2hJAk8OIiB/69VvEl3NZas/R+t6HvMA1lAODknl4BintNn
+e/8FRdaELCygA1BaLHt6itS2q2DxMB8321ffKbZDdqiJpgrZH6vFeGljpm+AmiV
lTPt9CVUeCjtFmexxqM4RmMQFtt5iaEv5+z1boR6ApEoRsTS7+g9lJnrBN8IRoO/
X0FcUOp8FHAwYBJzkkKYJh3jWdSQmJBEkZmH6h3qMeREWYKKT8ouwRsd0dBFJLv2
JcBpQyZiRHs/CVFgL7jciip/MuyjHke5gLIYWy8STXe/PcxImPMdLdmbiA212YvM
bn9qvLkZbDpeSfI72bF5KkP6R6fB5CBsSH78RG+EGqX79TfWm6/e4C83/8uniPTe
7RuQjXa1nkHqnpUYCmeuFy6Uw9wo9YiUkmF8f7aeHz+9m2ixPX7Z7IxMPDdVfxc7
O4m3ILbGR/SCXfTkh1jxiysKPhUGnENdVFaEvVCiFserDXfUhyKR++Ui49gFoMU0
3hMWgnObJfLjxcNAa2wDdv/lwKpmHGzUd5wbBtS84G09OW/lnyrObWIlPfXMBCg0
CEDC/nSNr4oB9dLFbvmX61Re5hShKdF2AqePLBCOh4ssi6GwYnKE+426d2zxZEu/
FzCkRu+jvRUHK/uWj4u4V0dW3e9f3ox/Xqzzy5xCuYPiupDLe1FFL2V4IyfsAt6s
Re4s7NTdZA9WO5QQEOAFyATUBX76+D7ZR7wN6Wbkm0/Fyf0V3/VQAOpqKu1Az95K
G6ENb1L16lyGP/He/C6hRh51EwNrcotfQnzygaHj6/ph+AidYmjBKSyHaPYIVDg2
HgEYGd/UfX4kKTB2YRSC3g4I3xEf5+0BchHXrMduebvC68i9pN/n26hc4ltXcqYF
WGYjyVKY0+fhsja3fi5GnWWlddM7lpeIw23tHBnkmwujstPVSNL3XFRaLTl1BGW1
f0L8gTfgoNrrGYP9JhQwBcTZdF9szL5zosw81RknP/0DT60Ce92ncMLeYdesBvt9
hmlvGfyw98lGX6ZN4HyPBM92BQizC7AGsGUYJrjuIFnDwHEiCwUDOg78kQEYrMsv
fHFLjdP+KsQB0O6HD+2vQ2V4HaC4wbpzp3ODZfXuxkQVLibpmXjxn7gwPEKyqot7
IngSHKezcq39Aes7oscmx5pJcIt+onTQXPC75m7s6gduxw9LzLECh7voeaWcilPF
l66OR81PBkTQgriEGiIvb+CDYa0MoeEdrHvt14gWH6WJnnf7cdD7kM5c3pBrFFl1
hfEC4ZBGLjDEcR8ilP0zC7GqbWm/3ho8wFimWkMVQlc68SqVOT6u6G8cSuSaXQKL
q+NfVDVSgTO8rEOA3ZmX0R53aXWKq6qZx21xqtxZ+LKS0T/3AnhEltm08j7mGKyJ
UQDxFLBmQSt0Ywq0ZvZJgFD+j+eiC3vq3BFJFie4HppuGoydsL2pVutDFDiJMuVF
6ble5zzykswhOW4QMbhkI1pR4y9NpXJC/xCAq/dXStNBOoCPBlcV7JBMAgltv1Xu
LSY+hKq7JfVAmHAzuI8VPXQ0q6vxHANKTEjhnt76+EABuGpXKyGQC12clRdqTl6I
gHVBi/onlAuJxNjckfkpfr8yKwqPy4LDIlBgYgL7mrj8Xgll9TDM2ZycCuTH2tR7
zsw6qh9QTDbyHmZJrCZNk7K+3zyvB73Fr9xP5hpjS/APBpmU5n7q1bNG8Mj7JdyF
zFkmIV8efJNts98nPTQCp2kQ7tVXZME4rOa6QVjI4begfqsYAArI1zvB8pK/K6gb
SWxcKOxSBH0AouPiJMPfqNqVUAfLZdK8uJ3Kh5yH74QI1RBQml75LaJ+H9jqqviI
fHW9+KEUoWY5cOcv9PnPktMT/vz9bk2WwV7l/dKz8I++/KTHfwnHUuEQ0tqXZFns
CMbMlnt3v1fKNu16m9QWm6d+JoRJ3lhLbPNOh4rPp4dDZi9bWx4t4pUatKPQVs2e
O21a6sL5cS+LRfDPXwYTWSgo8zrp9L2Y3dZxHnmx345zoUySLx4Up7Hj/xvv6nbt
JA+X61JZDo9BGFuDsdYtA/C3AOszbZB5xxAx2ys335FUPKQfpOCAUbH8bx1xzHh1
xMS/QbMrE8cQFyCrkfJ/TBVr5Pa3nbqTgHPb3M4O0J3qf0BmEDe1fRF1/AeSoQk4
yZ0TLkFM5/dlICUVyK0n9KaPi7bjlMYyw8u6+tNeDx5y2SYN7ePfBgqfybM6MZZc
+g4lxrSNLCnDyUDB+jPaLW+1RGzfA51M+MdAaYDxv9CGG30NuuB6aM2NoWHFx20C
wsSwBVmsk73EabXeJ6BMyIgT7tE9NakMwsR/awBkVCX9ALlmKjmaGicx9gmhX9kh
qwLo80jHhz/V1z470o8e10ldv5viL76iJCu2kYId957c1hxtKVsY2ZZm48iel6WN
bD7oR3hjWavl3PWPiOviMntpLZfnIwddkjVVmokaAIpK5iSGyv0JYcUeo9/gKp6b
GeWBRE4tLoDQ69X5SEuPVwvm/f+SNx7F8nwwVMAEnQjYksZAfJoQKyDXTjRjuhp8
l30x5yarZ4582jYcwdP+qcj5L0YOX6M1FnhnzVqJOYPe632MszyNAXEMrkgTFrp2
9h7LOyp5Goem7UHw454YbBNB5eHOa0ObVYyqE7cYiWNPfhAohs6DfXh7z+foO0kd
epSi/xSV+UoIC3S/tqPUl90W7nELaoypfB5cZKj+LdQcAZGVXjH3S8aBPg4oGqIL
kPRf7fhzQnhQYQMZunZ8+UciM2EWQNec07mYY87GrQSF+VX3vH+dHcrxayKzvTJw
8M7j5z/TIMdGKaMrWuxBSiL35W+Gt4Qvs0P+7lSeySX7p35JdvX3bFuVZNoLyRMw
tvfJ5MG/qhjXfp2yvHVxjdUCMDKmxpzgtJFHudcvNQQMymFwnYfsGLlU4796B2Rx
hKuLE62/ZHmbMixV1GeHmWH8SOTJvO/YBVyHQztygSJBeO7URK5wOl+nAdnbXhhD
Al5dFsLnR42kk4bl2qO4We1wCuFz9lL6ju2Di95PK0Zk//VhHipydMMn5Aa7v9W2
WZm8vVTCMstMF7WG8gWuaKlt5ERbXsM2QyStWmgL39UNneNbGBPnSpdDKq8JOgNO
HB4kfI7+PXCvGE9qENhjOGD5EKGAnyMjBYnJB+iJdSL0GofBYuslxsJIZF9musOb
k6yRATUres7ejJTaANgj30oRXBd4O6uz9Z6AZxMI3QKUbc+F0mhd3ciDvPh5ClKN
UghfrchUHkG4F6uOrwXroD3otlPNFElF0roLbX51UhdrhTnT8nf386U+uZ/m5u2U
swCqiiGu/03hBwrmtJncuU59QDutmNXolcCKjWZwtU64R3fXJedz5pBWcPSuu9jO
6Vt3rPaGLGALZrAa7ozN6V3qHPClQBCelwzM0TxiYAw14OJJD1K2so6tr4PdXd8o
zIzwv7WaSlptiKCZ225yP3PUcWJ06kZgZ7lSYG0OPw0f3nT8iDcDCLsy2q2OCJ1E
wdpGku+sNyVRDgDndUZbSrCfNH6Nf69Wyt5AnxLbbOKk0ZfOVVPqC168ZNir8d1d
IixvRul4KtPeYrhn4GN0U3xODP7aSlHTY696/4lYoDYGOMNJJc0bHf70Fb6FY00l
b7IfYwyJ1v9Rj5tHVP6lCsDQ2xl2ehUaUbMchCUtE+kWngHXcoAIgN6g0HMBD6qS
hgIXBs/qgQCA6kC34IuXLpDKsjWju/GVsL5Bibl8g80Z03KrPdSBgSpIevlwaepF
w8qiAtMsuB9VVsQY4OjfRT3zJV+bV5KyERjrFjgc59ZGTm7w1/aiLSZ648M/47WK
APOsETrFuMnzoVyOsVrMl4tZiBE5wQO5QFZoeeHB4smDZb/4gRn1FIeNzK6ZT9np
7vz7lQlXyRFeRyHS2v+eE2WEhPjF36tGs1ZzMSFux6ebfFbYzKpzcrA6tDISv6xf
Ft7hX4pXAX8l6p9naS6VJkhYAnULIPINaV7jfalQoZwgAWq7KI96wLjI7UKYtjXG
fgWp7Ij7d+3jJDVi5fkZqg4kdEN5CqGyteXmvur7SKyBhduN6Uh6UfCTpR1wGIz3
JilvalXHjBolx6J90Yxour+LHq6CNkQQudjshKFQMOQ4SfMMICAbxq59lOSP/T3z
XYYKRL6JIGK9Hf+X2PKGsDYOEBqX5ox/pu69GAQOkWmCQDunnnde7TSqSjFXSLNY
7leqBy4/7WPuo263PvRSh2YtOp0oNVbCfp7wdXxYI/QrMS8Y47cTpPIP99QtxLWS
P2jyQGM26uHSix2M5gUmzCb63lARyQ5b/+Yts9cCS9TFMyw64pbeKOAIJupQ4pQH
KCqcQMxbjBZUaX7t4vRv0/2/zQ5cr4AZ9tm0iEXO+gFZ3iko1QVUZbIo6HvPEF1L
KYFiDtLoCSydvy7FiqUY1RFDO6MD+E6LIpe/KM+8uXfhjwsELCb2CQX5xX3wpBiQ
YPTBNIFfislKFpzTN1ziMocKepV9Fm890voXkRZ/fKE6vZU6rUoqtIdU+W9i61QO
d7D72zmyO/JGf6LokJ7YQbFALzwk+6+c0MVnTnN7BHNxOU130Trsv1Nvn2jgBhO0
xL7qbF4O7o0qoWZQ6aA4tHGCjxOFlM/t4ATXWfxwD0rAatyRDzWfmTFJl1NgatDM
Cgrxvfq+Hbrtm3JkU2y4bnZXO4/pCUqBQi1fbDcf3kobAgrp73KW43Sv+gcIEh7t
86naFD06T+kch86raZVq3m8CyO5vInlvex/09XK8tBBH50qEQ9jx55wD9bUrsTsn
sVvJvkx1O2RWIP8ECqRB3QBeKi9X419b1KU4Hl2IC9E+dMQoriqNDAvxJECNu3UP
sPtGDC88UIscNoy1DoWCWyBqEnB3HHAbkEJGa3r08H8J+c3y9eAD2xz0LLvn2cih
nLTVE6QPIqVFH8l234ctvm/9/sHhgR7FJSnJv4fsB/bKEtbTz9ZTOmxLiYt0iNJC
qwRtN6qq7MMcOwpIcL969oM09un5juWBLvUTOPFVauAc3VaQXqAxmSRcDK9FgnMm
HQKmLps0gueNbzfFqo6gpH8IB2L/YwJznZXHgF50OxdKt+tAX9J2Z3kmkX9ki46Z
kByPbZlRb8pJysn0ZvkIuL8UXNcVrEOd3BsfFLutiRnOiqGvrxwWaXTAf7Vz+prT
tLKeVDkTI8sx2NP72lm4TuLdCt35I2NPFxOEcvHcCY4ycEaFJZJznRI/F3gx4uXi
riTnQaVQXM/NFoCqkfwRKrH/MZbpBkxs/0q+MCHMnAlraRRVbggoMoRVVy8SstWF
52diqd4Vk/fz7r11xbGtcJOdE/S1cTSmIVwKeo16RKJT6byw9inWpEzUzUNQ75/L
gkXaIgw06hzPzXE6hslkVKD5jigpGwQ1VJLh0ESQq5vvNKm0YX5I8eEyUxW12ajE
9fVim9topSEMuva9gy9dIgEWrKH0DkRJLkPUU4sNL/xcJC6Z6Kp/dv2VJYwhHcpe
JWw/HPASwCHZXe/WeYIc68NypX+o3CmYg62Sgs63Dd6QzNRt7BvRNJQ+QERQR2fS
/xo/dRoF2DqA84aSemjFC1rliVFN81399bbKgI4p7plb9F5VorwE3vMD2R6LmNCJ
J0GdrkWI9MqDq6bUJerOynML5pcw1GjadTOopgcvuOsdV7WWLwIWduW1UJw0JOzr
0/OLkEq1A09dGSRz/m38LbnzLVa5giIrT5lvJC1HwA9Umj0m4KfPTnnxHEPThRJv
+wMo5B+L+AD1+y68A/QCKBKmKoixHe+ziOhNDymiInHroa2OKZh3PKueSCcMsJN5
Hh+bEoum3B+B2IlVoJGoxuvJsCKsdsTdygQ9mw+Y9DyMyX3Ywt0zPcPxhZWuRFNq
jevsGYGX6BgdMdaXYdA8gs3kCIJr8PIACvCANdePMCea0Rvg1sy0PS6s9n7SsdQb
BBelj28qnhXUUA3C2pbpa8O4WzifKjxoVGVbszR0PO9UPdBB3avvFKDVIVxI0ZSb
Qc4NO5fmrBC1BTM4hOlV6LG5VYwUOsHpMKrzvxGK2hJaxxPYDROB78TJEZUdMIDz
gyzG5GVGALZRiYoZ0e5pdJm5U5FZrpu42DG3h5M5eVWJKX8sPpimL+2J28pMEAzF
JXEot/OB6vAYVqeYXMXpFO6eozGYJsvYcIdvt2JWy1o+G5XO/0Uif/j8K/ogJ8yo
HGimXRL3TYYGqobh9XO2H4nRlUlECKgPfNqxtjhpRocvdLTV8A6TCAIRILdWkZrg
mbr2Sm3pahVAfy+uW6a8n45jG3AzhQO/uxy6yNtUkb99kBJ9RScGrWBfr9DT3ZsK
RiX/mp0Ts+CYY6GDEBFcm69frYxJy3bwz24UUONMNalL/YvbAqFDsnHoakkLMem4
jpHUxEgdXtgOkde2aII7ioA5fg0OdXHuJHL4OfntZ6lxvWLgXtSDTYmXS7amPUnm
/2tENoZq9e1ZN23/lM1bWKJm8WTMKBzrr3RPzQl5GtwlV/i4L86BtUkDinHrHq7O
ULuJcOs19DaZ6MKd98mOM14l8im0m1J52Qki88rfWDBA29Vbl7dIiX10Q4qK76Cp
WU28PqPeBLqUg/RxFK3CKtN7Df2CwU0zcwKshOd5uTXMHccX+hvSTMzWxCF+NES9
YcvpX8IGEpYGDmaWqd7llEhCDCWWaNR5E437jaeLlRUxc1LGNo4UFgVJqT54SzZd
AMp2SFeQ3Afe49W+kxDsNU+ioXv3pFjs1WH57Kp4j5zFXCAGYUJ9EV/0eRtush2N
9sYzOZRAQbYKU5qqoVOwsMtiO7S677OStOcxdcMaTbgV19Xpbmt7aTrg+Yc2x6+x
BYeb4VTFqbNm4xWiFO6SwAEQs8vsVZ8PZowQLFTnCSW2mR1rq0gOOU83toJcLYVX
GkIAMlfIjGck1Zxeb85NgLt3uT43tr1J2Oc6CXlluCuP2au4iPEPqcs4UaAAUKF9
c/x0pqhbpv3ctvOZQCWnntNufTHQrft55DexZMcmNr+EYsG8zaJRibFBH0vSI6m3
OjPBgf4w1/SW9RJ+T0bJnvyifkXZukafejBmPDQjM7w6bGCruaTwcuiMXKv2h5nA
jGZiqQqyXYQaBP6Q11bCeAKrY4mplwOIAYYYhRffrRQXq+g76OqxvVPO9ph8c3iA
FjuqklPQKCW+Pnu/rzEIT0NZTM+jKyh0L277JVxAhQXfnNWxdAAOUnINRMp54Oxg
fBmvKmrqZUqfjQJNL5PMuKHG27Z6OKh0PwHr2mNbVhGHcCL20kXAVMb6/yZRgnZm
N+t1yo7kNdEzryidgGjSQ2RsMP4M+zOGpyb+Y5gsDIsuM+bycAeoTHW0EM6oLY9G
4I77G/f2D4Ht6br3Zp53JAoTJ7Ohipuskj/FQdwsollkRJV6qo6IefQAkw+wgbLg
apjwF4DL8VL7exsYTLAoDhPbjbu5ZyWkWTEdfdFjm+cBSMnh5FUgwiFgZNdw4vQe
DCuIzWQcEX0u1op0BJoWic9d8ExXZibKCCyPi66yRJ5Wpa/95Q4wXS1v8rQx9vmo
nErNgonnwl/nQhM9Y2JPGUd1PPKO04XD3EtR6RK71XAlUqQJtETOcFCRPOasv2b4
vGTRLa+fMtW/QiNpD+xLsIrRRIdwDfcWSuO1CisXib+c2RBuRkUnQUg61DVumyx+
CtWjUz0jJhng2a9viXg+iHPPg1Qb5APTCw5Prhy+gSMZtK+57Ceu0gYJ1DVT6Auy
zczglV23WOQjJ8e9hUrehSK9+2HSHXkndK3FCnOE2S5PcHawXwEoJWixK6m2SCIG
tRaWQu/rsr+FED/ePTEPoE2L1G64AVvtADeC5YL2yP1mp8qIra2A8prqS9rQ2oFG
Ej3LbVZ5EkX8UkB5F9NNRU4FDrbI/d5TzpBQHJStPR4+Or6PD4oeiOmBTjlX78ve
eE+c8TXLJMmrd8FuDPAA+kZKD3BzqDXcQVD8w2if5BMtZlXzswlFrRUcBf70roi4
kjatRVLTc4EQNNxihf20R1esy/hfWybd+fyAcVIgpbNNl6IUx0TXzTREBxqIrRsR
s9BmHvMA/GSdJuIfkiWUwzAVTJRtX2JZ8Cl7zaqlJ9BKa7MgwJYZ0ktVoasbCIJk
Vfyqk/vaJDOwTMfzUoFR8NZtoIUK5YE5Z+akXMmadFGzr3bbqLJ6jicPHm7+koXm
/P9hP85J4a0XRqb3tDVJ7b1RioMSJhDAxCl9h4ZciYJK9T0fZJ3wUTEjdaLw1HiS
kxX6ezFLe6rID4ZS7IFszBDkF7pScve3xUI6kqYRmIUynTG6Y+5bTaXqfodzMtVx
uWvrEhDsCTdlEyl7diFAfNROTvmGlHiwy/pkEcYnf9tKpqK7JqCtZZW+H+XTao1B
NV6QBUWHOre8rdZs4jz3+kO2Ed5d6H1aaInw6ts3K2Hh4SLqZhoPrjaQt/UQMbZa
I69gSCbB8wzoaIudCSGRx7E32pwjVK7PikdhWTn25/dD5rGyoGo5iyo21fLzmmfN
Cu+C/924jHoRNSeVScg10wQ/ZmohsT16GxDDiOmgl63jy+CU8Mtj/CyG/htK7xXn
th+QUjuY0YheS7n0mXCobHM5jw5hpFGVoiwPOC9pe/z1A4KaGobI8jtQXAJBUqh0
m16TyFLEbdVH3JWFyCP1Uvd7hrFOdLg21BVJWZC7LHSkkLzbpSwbSVWauq3XYIzo
vLDMddYDDMw7ceJCEZCXX9qIzM+z35jQOiFnf5McHjU/3A4ODjXvelimVKQNYjWd
B46s9BpAWzX3h1kBQapZOmqlaKVta2oMS0QmbyKWij7UdYSk7BC+AQi666oIK4Kb
MXaWFiJQ76jL6DmcHOPEcHYzFakoMlAOf94gqD5yIqPlU0N5t1Wwk3OylAWJsm0V
5b5WriYCNyotYa1awngCXpDJqV6in0TzZFOqeKsNHC1cz235XzMXUk+awH6PmJOb
QyZgYEk14aSj63IRys+hdNL/6o8EANf03tHbDYSLnmLXoi1xKn9ARY4hrhArjGyE
Y3GKcWKgRapmz+O54RqFyjtfNx4bd0Er7RWEDS9t7bDMcP7CJS5vZU1g7oIkPoWs
911rZgiwp9om4th36LpBQiBJdCY+nCN6WaMEbnT+NEuLIY5/eDUhWyvhgG/wHPUT
wv8pYeeshcaQ4BLt7IgFe0BxW+I/BXyDjQLfHwiJy2lnG9hj74e5dpSu4GXesaoT
TooL3cgGXAbcSKJBah1sQj966LFThR9x+m3miVQ+lkQyFyHFVCTcTp0ec0693Oth
LklhRl/Y5RU/jdOio9uc5hxFZcyBJw/J4MUHiL8kM0IewfYuS210kDIiPtc5XW1j
YiJ7/rsxzxsoOL4V0VMLAlPXt0o3CY56Zdpt9NtQOOQ7/Rz9o7mvCcAVD0x8vjGY
uQoBrU67qthtkVOSr6y8B4krSahaTxKYolWRP+0AKLiHbB4EgSpuSYXjovhav0aX
W8AvPb8EzbEI4n5oglf1xNLNLdI+AYv5cO/0GFJPOyaWTYRt7KxSq/JPw0xWKNFX
fkt2E14DKqUq0sYkM7YTcQmYqV9ZmHnY6NYiKf58RVPsz8NGjxP5B4kYb7BPcdld
06zoSrwxvrZZQip1+xOVtq1bwpZZh8Lshmmf5UzH4MFYLycVnxhqxVNpNuE4/SEN
YUJ3lNUJlnE6nX95X6tCj3JhEkrs1RqFFSd+gYuTHW6x2MbEXFb/V/Q1YN1mVpBy
DYkmD6atoHMBZmJ2FLdA+kTQ/QT+zAgGnO7rgA3eFZqPwsVwgyouIZWUZqOFpImA
nQHn800ai3tmpjVEgGyfxlyFZL6XT0BSVwOT23AyOTxkNFCJvtvcCp6+WRhR6SyT
d1dkiGQ4oE4hIFa3fLy9lX9jOzSIQOMQzcoNMoMmtW6ye5O8c0upL0vOhNqgi/dS
HkVg94q6MNOlj6QCTugfbqVGkiTqoE2EsmomQG7wIMR0CItsLg1E1KluiuCw5QVe
vKhS9TRIHlqWfzuB5IfXOK3yOTLzDdZW0XDreqxIm8iAlfJPHPPBfrz5vYaZRM6I
W9KWVBIk7TzjyM+LXhu2hk55c/QUNezsghnMji3EoogLQ6QPurxLxNGzNzmwCkF4
T/KD1DyQINH65Xqh5oLa9EZyPGVBPFqN58yfZhHbAMsoLMO0uOModFSO4csxpbaY
S74UBx+yGEvh3U9Ik+UHoQlvULid8W5Xu74BjtM3BOE5qUUXxFu9FyGCXvPdSor3
Y/XV5E/7KWTIPJQbKNrj/LVlHuOSsp8S5WmaQzs5oxXMsZaXC1MO5kyhLW7cJ2s/
zgt7MI4MA9OABYqa9Q+NBkb3tsAYxDE2iDUs6LJNzWsIS+Wg08HE7yEJjij5p1/G
LvPj7ZR7QQmdGBV/KYHDM76sD7/jUt1mMQp7jcAdxA7ANVxpqKGpVzZbmjtrryOZ
FHG0Mqqy3+T2L081Ou0rUSe+FBL1NlYLkJFHvcFcANsSFgJcNY92iOuWPIIVYsN9
X/H8xdnBx5h58mR1MWKF3zESQ3xo8zzRM6PGKINn9P1KLoVJTyt4x0djSVwJpifb
Uc3mAL9Qk22WcG/BOChMSj9LsgLHcyG+ftbmtXfIe+Pf+zCZ52zXFWiPfBAZdbpV
iitf3xxDYqCPxEojaae2m35++MRFJsOlDWr5QMwlkOBodpFhWwQUO+63Tj++8rGk
lb0sHh6JepUIkLrNwPTWETth9A1Mr9UycMU/Tm2VmLzmJB8Wxd2AGLlsIn1RiZBE
Ezqdsq9JP/TRricD38vGyX6ts18PnfLfbyG+osbyK0H/PDZgmidSM5/lBwku4Wgq
YEOhBQHjTXBDVAYo/k/GRNy69vWO43LATvkH6pYhvGjiR0aLdSQpe398TCTrZzIK
+m6BxSKeHWZKcagf9/druIGWqrSZmyY3hbb58pC1uoVs+o9HM5QqscMZ+rMuUsEL
lUFL7tX1yeWoZb+kBJ1W4gdeviWscZsKsYBpH/CRmuaqr15lcq6Tg0J3adR7DaM5
MaV5D4YX74dMcjxcn4R1Lyc4WfR2kMfN3iLzj5phyIr5kfuNupMNTT1BPwCj67Vl
4aFFQi1dgPYl2fY1q8ACSA/UJfVUJlwhDZfXZcoKm762YzhMe6ctCVfbzm6xDM25
bHkUWPp0Mji+pShJm/y1KKbIuZ9p9AJyQNqLw+O4j6X1bc9p76ZsKapzNb1gVCb2
35W9qUAyogYrVT7FNMrf+BE+1wNDFY2OY4joxyWUdkENmwGj2puBAeGmoRNI8/1s
NGP+QzTGIVJsHaJP2V513NQ3E8u48nx5KHqqA9eIFVFNlsSKYzrlsKV8DjXITRQd
Xqt35Nx/DSAfu+GWAql6G7/YeAKipndiwfr3R3o0okUnYQ0JBMtosbpUHlfAhY0b
I6R8B5ebm9z9nUmwuuPz2txoFWVyKufsfbdf3gEQ/vM29/DWeuFYcZnTueIAH74x
mJCY7fMx0oKo4deuvAhnn/hvwuqJ8GjXetI0wVT5OSmfZ6KJOCk+GqFrGBj8RQ29
QKCB2MEY2+0iEHZTEyALD3yETNJH9XZBqC5Lz6XyydpV2zO8XpS9rh1RGgHf6mQG
wSxNy5wXUX0iaZku6LIi0N2RmBeUYU+FQAwIMSZwzsKeu/a4F6lqEr8Ws/SnPjY9
V/QHcNYfGrgQPFk3QJTbFo05OSLmzzJ23PqQ2+lxRzejTWlSNdXy2m+qNAVqom9P
Bt80Pot8hAO/ZF8SkvdBknIQlbogtVrdioMt1PaskP1DWlIZrT4YrDSxghaIn5OS
0uu2UoKk23EGfahdU9K/RExlrRG51TO3KmlvLpSDl+J0pLiGjGENPYzogpIXNeSK
og5/hUc62s5GOvg3iEW9vNlTdGMMBCkppnytJLimUAhzvQeSwqeQFCKZ8vCDoPgh
3Yi9TpCI3pniFYy+sghBBHzgvOelPFFzoijkKTonBTvyZL4DGVLOZEMU9Z/dM3tp
ARX87yBXma47XO9eFnblbEWU1qoNF1tA+/Ut/NZI6/KKoSvYzs8AU6HWyeV3jVJd
iUT2H0VYj1Y1zofSMvFnCOkN1zFvRe6Ra7XOiOsk3LI5zT4+sLZEO3Bw8LJxhX68
awawrFiAGgSojhia0Pw3aza04em8GiANWaF8r5pkgfOiN5LFDmnaeHkBVbsjK0S0
z0Qd2cAQbK73JPjCJbPBVgss24ASxtzIWjmkJDzWatLhIUz0sOFra9ljzY6xg93j
oiWWbXS+FiiH4Z6rpaDGxOwChfZzBLDzyeBzz+1XT9iTLxUODGp51XdSmuKG0L5m
7458su2PQiyge17tPwOjTd9HZAK/1f2CBNIoQ0lEhSgTRYVDxlV3RkEI18nn4k6u
Y5BuIhnhl4vkgPEbdZ0L2cwShgGegh2UX05p6nLWJiZ8hyJvb+2oaLAtZTNpx59Q
zELzjTKIiFNQZUsTW+1Dj2C/7C0Qn4tagpgc9sADVRKaC972oRxhw0DSe09WkRQC
L1baLhpE8RW2iOo0jE3EXI7InHmKaU4FYFy/nc1mbXrnWmBOLai4JcHbBPxFxMRm
Gmd7FWYNVMuZRFMPUy2SdVvcPNJmQYsflW+DznpCMPQmfjd3SYubwXrPchnekURZ
6LX5NX664n0VLAJEvbu5m5qr/4Wt8cdGmM5s7PXSQSobuGEhxmHrF4WaO7c14IAD
MoP7DH76zcFTWujx/REN4Blbtv8pvFBHcyczeLbKsLFPzOkdMVWGKH/rmupDyOov
1yjEXLJ+j0vh1BAvU7+oUuuJ1OsZqdZwBZBS/LeCiVI6mVXEpVYStQ3lT/1cJ3OC
I0hGGmGeG3LgG1mZIwVjaAhQrrwWjir/4PfpIqRAetsZ2cWX56fuEWcccnwT3IV+
I6ol0wI7GZ5vA9nZyeFKXQw32JSTLl+A0bj772h10jk8xNSoWT+0s9L30Rj0+4St
Ri7UCZDcj5H6HYd0cZTzpsmfmx0Rj8LRtKuDyGB+OpxTob8md9zrNDGLxz61E0Kr
csukmbzWRLeBngBV99FlDx0+4VzGpM5lWQDNDtKXLrodI3QIAJiVVk5ChxuMKhO2
pLqnEf2dBAvUOTGIDenQNu9s9IWyoKrm2QxixJYpS8UQG+yEaXSxu3AjtFUmmMi4
hEZI3vQ9WpczVB6ftC5Q9rytBTCOkfPO6tTGkoLtdiZMd2JRYoS1iCs6PEMDAm7W
XI31vHlLtW3TdAqN9b0HEM5y0bVfv3U07qfIesRAzbHYfdg/rV2vJzYS3lqH6Oy7
dvzJQvmopCFJOYPSPJMERp+KG/EXj+rRIaYntn4VjS0hf9ACyLekarWhAoEzGc3G
288mTTHEhTcnzE4TalEgVHPXI9vOpr7fcI4o7gtaWzUhS44AtBYSdXNcfUXLNsYh
HPjzRcowq9jXls8bRDOPItozcU4d1G7Vawcd1amwzsK+LH8nR7JIdiTWXI4AQ36I
wLpjSwHIRHc1Sikli5xjVTwDg/Uvj1aiBELhXW/ay6k9/5zUH1ndEN8A+GQvaOaL
6clk/Hx/gibdwpjO/7/z9KDcRMBdX1FzApeq4k3j0GD/tj6LPsI0n/PaFuf224gK
M/gsj8QJFMF28tGmeBSd56/HHshtpJmAftSeTlPNvDfsLwn9nLzuLiOuBUFmBJZ9
zsFsVusyn0K/Fj+Ez1NB3374T9mwpeoAn/2ZDMUFnSfUlRcgWkLG5Oh07EyrgH/1
DKqeB3UVBPremwLQZGnTBAJ10F4Akz/XxbblW9rn0Jga+pWLY5B/0I9ZCUIRtqfq
sPKEPTAGWqpTnFrT4Hlvk4KTGbbx4JwshRkgsrn5MzSaslp4L6+jOl8t6ghckn4A
QtFfbjhPKraJnG6cuLCsJtnktXMjhwslsIyMm8ZpqSsl1q2lxhgXdPZvNC46czUO
eVozZFheVeQtFRrjyamdkH4AR92WgV645ncBlN130DBHz9j4mFovVIjh5VsNaKyK
x6oXyx2VFa14AdRFjUx2qhuQyBcYD6RV9965Wx3paueo8b1ZUsQdeFWfaWUL3OfU
G0DcYjY+qX88qWHBlG9ykF3h9hZNbBKhz+4nMpIxjKt3uRB+kJgp3nLGloYAcmOp
y3MsYnHJt9POx1h3ozrErk+Pfyhte5Lhf/fikV7e32rKekiEaB2QrYqkaBusi18C
u68Mz2rnckkqOSTNQREHQXXIm2CD00/ZxNxpUhdPKhkfskKwwseMVAzcz/B16EvK
jPNNinZrv81Qe6iOLF7FNLphf3MP9Ig/P7f5jB34eXw6rHxWqRUNKey/YLmTa0g4
LpKR5O+vEYxddCGdCviXH8lFBiNvywfjwFiM6H61iTXV1EIxYw9BgkigMH6NBQ2b
SfN/8+i1VZPu8G1/jg7Lwm1oLnWr4KdsEFHeJrUQu9WBX4XWxJHH3AaUFt6AawF6
tpyaUBEDRuxykxe6iULGNbfDJcTZ+YXzNDIUi7gKztjApD2KLu1FCrGmjseWjSks
WIEWhQHEMv8aD9Cn9MNFI1Tn6GnRC53RjNriH0JgEd6URbFNRVYfMXExqzLoxRyB
xXbXibfcPl2Z+2kOAKAax/UFG3MO3QhWFI+mokdNuftsIwRtZ0d7hlY7aREaiYpG
Lu1Fngx+psa+hfP92hPVZQ/HOeQYCpSt4HOwiJluFigjSyPgEB7+Jy1Y1AXbJTPZ
L596JSwvRhdkf6QTxgbczuyH8aV/k5fNedMSzmMibyeGjH/HQ7FHUO2MtLh4AuT1
5ewwLHra0G4cxWK6Xle4kk4/4sC1heK6Td3uYYU1f4Ge135rhHPM1oXCowjnQI0S
7IZGoImijw4c0U5xU6Z2TSqWqh8uJR88rAWWShozTms3bXTH1E5JJM0m38OOBRJQ
aQGe7hteAXbo/qXFtK+js63y5T6MhM1CKJ4mj9VzQWmyMrCJrzwS65GEZJ5rCRCo
JMXx9zWIsd+CMlcIH3Z4/md7AdWXE6w+FcjIF2uybkbOdGGop5KSKY4hpVj0VpCY
j8MlUWuTe7y2RYMQcUyMSWGoO1S+d7YhU8TGkMyGJKzPeNx3JzTy30rOFuqzQGPI
ZUt+PTgit1SVQyuoGpT1+JoWSs00TtVgEA4UaIEMa3udezv4cnVBdsRSPOiYYwWY
aEgaV4xHBB+YBm0hh4vHCRx+pd9OVSLTZb/CuX5Q4nqzHlVG2teSk3yJ/m0/SCAo
SykAGLhCqo1+MM2AbRTnhUf/kKNErqe1A033+WwLyS7Qy02/wyHO8EB/NHHF5PE6
DZyGy5Auu6yvkZyC2cozH7bKBFpEb+Nhm/tqdYCky3n1N+pfcj7Og3j5nCT8Lel3
pVAny17wNoao134bq1YGpb80lhc7WVjjR4/Y/aDLBJqJES2ePFQQ2tl5RkUcKpVs
VANUzW+9pKK1GTQDSA1W3I7W49sR8u2Va4XvhlHkFyYsZGs0i/YI3dffawZ61A6L
F4PIqN3a0PakvBd5RQUnZwDoZNM5opGZC/M1tPG9AYAQeS9b7UrIDE5wBGOCiXrd
5HqsfYiS0FEHEWWr7kM0yiWUQ8ipFEOIoEN6mhoJRSOFlD3SitPymz1N55zrai48
gRvWp4v6QgwT/y1B1LaTRmywjkNw5/Yc11T3Zdc/ABbybHL9jt6LNVGdpX2U3h7e
3fdLYcUSU0vap2GD7i2Liw35Bqyzs1d7jxMLj9tWTvmX2uwRml3VsfMJyN42zI5q
AueYhGDLrDoW3eJYVsy0JYpgyrSPXo1mLh+/zhhBLwOqxAPSqq1avysi31DrrBb8
UIgXoGBIgDqyNsjUfLng2ss1q5WGnKc0icAUUGEa7vj4aqDQTwbgsotoT0v4/3Lr
Ef2w8ueW7Svvt1ojOuODbAH+3kiGerh6lz66mqnqbCYcy1tT25P5/92Kfrfc2AjP
z2+nmve+XfW5ChLSP5cDMIHDhDVn+P/hcbQczJa5ss5a06/5Lb1Jxsf9Z09EHcX3
Q2jbR46aY70yMx8zYvUGzY2qvVtMMP2gQB+x+yWK5DXFtuFW1tX73zprPJ4ONsXB
FSS0zm4Tzl2wqIxHQLsKRRhvnZzkSlqjgb9VML+gXq+eNxAeqvodiQFEK/6P2zex
XH906+G/nqeiyYCBjJGzyw2VI6XkISsKTyE8aD0PITJDlcmTf5LM8y+ApWT4BS4d
LRzRjBK6qcQ/PbzTqjRPrhUk4isyscY5CZ9vvRQYFjpdJ5sshZMvvIsmkMgxu35+
2oUaCEUd70vhVzAewFeaePgN1YJ8fTkMtZRY2oXOnoiGuyPiaeI0KmpmVHEWfpyy
oE2BzChSNMbNNztYFcWixXJLofKCA9aGnrGsqW+/34ankgt9yVSYhDEG7J3Ij6Px
yciGY6glLLiQ0zh7c4dIkr4giEyD6b4g7FkOZqg3lFL1DuW7I2SwHIQXbfnvRioj
valsDaGVdbo4ztcrBT/ZA348XJzT6I+n0TWCol3y3Ugi8wAeWfq1Gus64v68vErj
pgAsBt2a3KUQ+V24inDPKPBaHYaNxAwVg25W9M1GjNY7Xf1gnY/QAuaEuDI9S11I
QFDc4VNyUQvy/OGsHYrlHoVZq7wCFw3agUEaKFq9/AvNIPSuRl5/7kKqkfWdg9Mr
AgB8t+hmAhULMn/mnnTrI3dCcqJuleMwSuMtGPOL/R4PRkULjRdDD14PeVQbRLMS
qsL/iMqAs7mUgAGSGkWiDTH1MNTDYeRR+l6mvXVSrNwv6NiL0NG8AvMoHharTjCy
B9zcj32TgmtZ5SEP0yvaGbgVCnYw8gUBjBINSKbbQtsLh3xYi4kRBdtfJN1k+UUa
r4kARhCAwDhsYY6SCg+0X+QnLAJW6wdNO8kPDZgbvsIZvuib88E6icI6DDNMIokH
H5OHFsa5lacH+J7kTnZnRdX7vz1HAM+KEVpk+C0MyqcJbwVAx2lDksBrLnnza0fi
BeJnxZYUXjQww3a/KG0AQGiyO02qezpT8pB5rTkq/GLUyZzDfy+cflKPPaM6EV4j
gG9Xl6x0LkLNLDsBLIFyJrNjr1M9sSDCzWlsB/IGOS5ScVMDDx9BMS7QSjHNigCF
rZIMn8xWwmNcFWDOO9Nafy7p17PSzp4KHc4i4L05Sgn026hlbO/egIszbyM4DKwY
hj81585jzoNNEIEMQmTZ7pHAwvYobLdg5H+PDsIdvBIclFGTQ3kMJd5oGA79Ykyp
JuikjRg4i8Zc0+8I1/uWLthOOgxKwm31ZcB1vkhmpA4uZdoylCDapWQ5mfy7h8TJ
XTaNGlHKiwuCtEpc8oPbH769J1RvKzXfZuav9W+eGrOcBPZ/XPxv3ZEKURAzlsek
Pcbtqedg0ixTmHrRz3UJAYqmrhs7altiosXn0fZPzazR+PlQw+2c28yMt5hZW7Rb
mpblVLFcfAKxImDaqpu3CRwt1hmhivWDUq25+3Vr3JjPuga1zNFTwEG+fvTpNjOV
R7c01+tizJVSoISsVXDbNe72tTzOEdfRJWxes2E6hjLXtbdnEg/T9iJ70Y7+altP
+EtIvInfEcN2+EFjIqcLkxGuYmg+EgxGAL2omqSo/8g5ZmrtA+t87iedO5Ko34wI
41JaV4ch3hXMVOGp1YYP25sMzdyPP4/mGyFMt2YewxE3fEEsIdo5APF/EbecOcdr
jJdx83xqrTBC85/Ro+PGlslUBRlCM15Jc0XBTjtvROrisiPE8Kfmo9mvEMHgaiN+
7GuIMC8mx5rhOnRivbAtXqyUIE7hybzTg+65G1ab2EzcBhaNpHx2q+rPNH1uqoFF
efHPbnvb394srAfLIV1Tzf/OnS9B+2M3D/mwSIblxpev0P3wcINZdsmqrjRkgfAv
LXmYlwN02CAvuXmS+Ngi0bTNsh70m3M0WmXHAqoei+VKZOjF0nDCTwGoX5qW78ax
wFli5gcwwJnHWc1X12LZx9YLMq1UofK3avykLLP9HfHxOjj0Cfjmx6l+lJgk7WkA
Syj7jVzhOiJzUrnKv5b4xbavWYzlhTPG0AwN/v1isdCQzQ8lHsYqL4wuA/4S0pcA
YPLWPxAAgw/wElZSiBBTM18qLB37Ay5OSQus3yGVbeG/SWKmNxLSLZt+4RUW4RFm
0c9avm69FYCrLfCPrz5s82dsuhE8Ved0RnFajrRu2ELvSSIV7ijOGduDo/Rp+bPo
r/Gu4kLQSWYdlk8I2ndCePdZzHfGc+ENXslGcQCobf06r85n1S8MKIT1jMK5W0gg
a5i/NZX2BY+roWf0g973rdoRjGtGXm8EcZAsdSGRy+4uovLxzNlXZqD1zg/CqEMw
7N2c5NJGOjdc2xtiJDfFYd9ccaxWLpbjRgIxHZfuokYui3Hom0DWsq87aNxxZ478
ZNjwBWCLgaUyfywfW9FgU43xCCHO/gNCwnJC4AdW4ZE9Ymn+eZl/MUEjnTeh2cBI
egnxJXA6iMgh6Lg8JHw8UeOW6xIh1wGtISW9mqVKK7rt9LIydUICJoly0+TGQSiQ
UcySnsUmTZYBv+ltnBSirwqimndHSRmdHxuBOvpzR6+BEcHwAciN2nG/j1+MN7eU
sWAucfOH/7ae9axpvQcMu9BZJZZaMIlFoKfqUGlkUfIeS7821liTLhTmS7eC6RsX
yC35L68RGG4J/PwvQioUhjECHkbwpFd8+35bn4Iv15TePHp1+sqQap83YeYF1R4X
Te3oKLyCC0h8Xeuhs9OJYW7+hdmPIct/QDqOWgMGeHGGH2UMOabUi2luaiMw3xji
pkY/vhzmwwPgrfq1PAlsrla2hNjbm3hlG1lzASR6OEp8vx7gvTWmXMIk/OOqaj5P
xsyGoPTTRr+0sctoDbUbjFC/uUbpy9O2XigQidRJ24YfyjmXAXGwCx+ZPfIfcykA
A20RlxqA5EFgMGIPsrax55RRtJfH/T3AsPXfNCVO1aK3SMhtJEVIiNrU+KuyAkoS
672pnrPP89krd+UqV9C6PVzj9hs7a39gLmHSfgiBC+l9rDWFbt5KHgulca8nJLIK
h2bg7KNMuD/3qAfuEd1gdcXGY71If/7XXvvoZOFWubz/u24IotJdd+DnvfxHWHEi
/JQCEr/5sHKQhYmN/xa1uacm3v5CWMqWmDofONTf2z1d+BDzN8Ud45FbdDGPhJxM
V1xCJHhTwCW7zay6dN0zM2Pfvuo4C0AZJCmmy8cj3mi32QKG5qy4PnfLar6AP3L3
WwOHDs+ep5O2KjnRTNV5g8VOmQHRTn+opDwYwjQDNq1K69geelutkdUR+q2/BOBJ
D9IMnfLJU0CtusE0Wyo8ifr6Mh0/obIu/ft1EP+DMBfJNJK5648nJYr0JzHdi8kU
HizQvbJ6JJ/yu9U/YOa0OoSWC6nZL215Zw4WAiFublLjHUKA9hwI2A6P04DxExEg
YzvzMIeJFY9EIHq7/LKkJsY4KrkUClMJEE6Z4anOoAC6DUaUbhNBlScPvG3bBjzE
wmgjqwujiLQX6/gFeUjW8KmhVbHf+f3BRfmiFOFFai4dtgv7kiHPdy3CS8BlkckY
wyC11wK0NxoybI0WDBpaWT+T46Bhjj39ew5mZkgRqTfXqWB8RdhDdfbi5Ky8L0mA
nsXf5eq5fiEJ3/3yX1JcJ/4sef5Fz+7SS3XGEbP6E5BxB8pjqxoo2s2gwXp8N9pp
5B1sGUAjPkLZ6iU42g1WQSy/mFaW4X4nQXo/43yj75NB5xlwxv4RCG2A7EkLHzXU
A+pP0DVpTx2nEysEjquueEq80U02bdO0vO9fCKJXnW+L/8LkDBS0O0uVgZ5BtnUu
5ltx57ATyYBTP+739SyyGO0yEZ4CN6IRfMuRBWVUKsy5jbIS49ScnoVC+wuM0YFt
8Jaot6SZ0zYuf3oFMnLVoS8oGtnIIqR6AjFzFtT858Q34uQbsr3U+jGA24cjH/y6
8K6RVZoEqU0wrbm+ZvDvcnbGT7n69xOyVBolVIgi9I3jyd/7Op06nF8aeyGox51Q
gYHkItTkzY5YAPuycOZGa4zyBoRObs4YuxlGDpyhV9lUZRkb/s+Y+GYnZBYkjOjC
psO3kARgYz+I6rnqFvWvulh58Rdrors+S2Ixsd6wO8bEBIOGaLk2UokTc1X0FE3t
1wqTxSkYZT71+TFB7I4dC+vH7oggK83KISPLCyY3FJkNak6TNIVDOap3U2O+C7j9
vecID9EtzjKnZqc/v5KpZLWUkEvmtl+RUsE0Sewcp59+0qpk+0L0QGvbxR7HSCrN
QxfAcIaLmJy4j32IxfhTIrW2MTHghggsMRXEElC1BUrVDdvZD3SJvStMl1AjDGWi
zSijqxVXmo/O1Jrpvl9D+wzCaHLqx/LPBxCQcSfQknrLSjsrDPpTtNgozfaeA5Eq
/i2te7dM9xY7o/E3s9ZAPty01QhU92f0UK1BiLZzi2YH1zrGTL0HkLNQ+MTQzY8A
tSCk7yp4uezZLJqA9c+VdQSz5jXyG+MNtFKSNsxOs4NLlyGB/3B7Cqlf425ZeLXA
51txLd0dmJBf+g8e462DkWnVKspmKBCIARoz5kiXVuX5IzU8J2jb9MRKDQp4+jw2
HwhnvaSKcH5RZUOshSKHIntriaYPZOtdoVVuc97Dq4tkhBnEnaqxp88M3QRXSS/Y
7NssNzU/3eqfwkfwt5XZFkUvwor2+c9pnxbEnX1zclwzZRK2BGLrV8ux2aSQ363i
3kWCkpLUYFKzf8qAr7TO64cQoQztus1Av1/3wMwBkdghKwE7EMCV1uyOF4gwIFzo
hOt9xXLb69+nnqrvGCdHhPnUn2vvoDZKcLOCPy3Redr++i/uwtR/1QhhBuGH1qQg
dgHWDJ80XnQ15hL2JTscyIstHU8qY0xhua0iYRdFxeBSmPKJ/6j6zHQLZTz8qggi
xd987zN/tbxN4kIXg1P7+utIPNiwErwSfZcQsKbS7aPPpOqCHqWnvml9Zpp1mLUc
jeu4BwNN94uu5yXZoUwBSD+2o6eCrIMQM/fRNXYXPwlvymnupRFMhmgWoroyY370
GvN1D5zqOSbkCRP9733Gyzz8TlytSNCf8F0KJ68kgsoAsEbf5Lc1OHO61+HDS1wJ
pVlumt9ls+CHdyLKHuWqiiXbCBnZzQKPNd+5WL/jvniTnKz83upGkwLy1dH0faJ8
GWk53Vkjm4ajjg7FxT9qIjdy7D91+P4/vMWOZFpveqyuh5P55clrYqNiIQMEsr8P
VLDs+1F4c7zypEXLGndTZ1/aanDRF8MnS2qPj6OBDJ/4jnPdcGMKds/mb79MXi2O
hIGUoDZXsxego8ZRktcADipXi4GcV6wUZzA9iYJkYzvJtsJARq/Og7iMH3/XqO7v
9MHio28sUgHSXlExn5X8Es9ilA/21wFLPAo9QCVuqSKbdzyKVRTN11/IWL0wT6ua
f7YMkE0UznFjv0hoA5EYyjsaJlqiN3Dk2aLvI5d9uYnfb+cUnuyZiqoimTEcaa6r
wNp1CzeDj3xgg/qb9hG270yxp/LllWvN2Jn1lfOdWzfdGI+6F4VkQiAqIYI7V2nx
eQhTW3oqHHReIVmJJzFg/DrCEdX7S8P7BL/DZJVb2UrJKIqSrrciIsquf6ZVclSP
sMMhL+55cHD3rZWnKcUuXk/TkQW6OAZw04/f+UHy1Yj6HGto469nlSHJ4FIwT9H+
eIt0chn1uPv/yLEszb9/CVOJCQ77zO4kNdFSXryFG2awrlEvbxKOhF72J3FI5rvJ
n4vrIuVkXD1H49s9MROR/2DNkHzznLU6OCqP+D10lEW6BNvtVkumd1ue7F1XaJ5n
EVdXazg2fdXM7ZualSoqdcKgi6/WvUZH5qvbwgcL/Pcs4zbSmh2h5PhwkrWESRmp
l8X9N7xuS5eiW66tjiP62QEk9a2RIy91R4Yj3xUm+S4WrElp3QTEAaIgeSgZsUNt
wTBYI9vjBPQ0Drg7qzEOreFbDJydjHFNZSYk1Y3keXUz0EdseKgAHNasFN/Phsk9
e7nnGSbHRs+lfk1csUmPv04XKjh7SgCb8xd9kUasSmAvx39aHunGNJTu+O772awt
yvpjYFcIxk0RG1URa9+FVHBg7I5hnPGYFfNgomuZQmuL0XtaXCIK9EfEOUmBwoOF
V/qW0VoLF9rHtY+x1yQnzHYqv/1nB8Y8ZdNKjvmcDUbgm51z2hGI1WgVZP0U01rU
RbcQNPYu4cgRg4J3o1oo9rN+lC30Okw25kEnES7bPkY3diBji8SuZHoLfA1emY1y
ToLM/oKI0qzXa3DXsPyfVfKcNRe7JUu+a9tFYkKGHHr+Gw3OVabtzAUiYYZYTCyt
NmjBFiepArc6/ANQWy9zZWpDz5DBjSmg3ZZloGo/ylqqjcUCSRD8qW+qXVifrFp6
xe1PCLutoZIMWiiSPppRSBYKsFaQgKm4+QL9f28vphurQM2wMH/7kTgtIfnPW1vN
qQCngtPmQKcoT6tk5LOhM8ksHcgxyImCwmmBD1OcCtL+0pile+FkoTtk8sRUMnau
IxqZdCNKPpUC3FPzYaYz0JyntNgCD5XBiegP1m+vW+IcmInbhHl6zQzPrWY5tiEt
l6HubisC26ylNI60HnjrckIS+pCB4KWHEsTtrjeaL66t7Qg0SqFExxfdK7CblwGV
zi2OXHdg+U3cMYILPQ49iPo+pU43HMj33X7zlVMqgIBoT3wIjNdXYB5JNibBSjMa
WuYAf4r+yMd+p+d20HRwn9lBDW/n5wrBszwjvAL/o2jtmUwPxFv09S2RBJlCU4Gd
lbeSOSJf4wtbPchM7nJQ2D22+13ZZjk1broXN2RFBhplDVGTBZvw2xuER8pIT/RW
DVhDYu7b7jTWJ82AXWO4eBQs2zxWwBQSF0L7u5xOXCiL18xDlExxdJ5Lx/rWOVph
DZKf2Ur4CMbHQSIctB2UzrbPCqVAe+i2TQJ0rWs6p37yG20yxKtDBBgILe4yoOWJ
vQA/fN5/JFFfcYE9JR8VjRXK/g8KfFg0Ch8DxEpKO0BtR14R7Ik5iuUs9xFYW4f4
DTe6OtmoIOmWv9+r9K/fyv+1o6EFDbPVCnn9YVGZ6xb5T2XWTi3SGhkkbVjZkcS1
pMsYfDLyAPmsNmw5bkF+Ol094iDgsGJs2B9aHlNAF6YurJMuu2XWEwxIY97Loi06
X7CeiAdzY0gsmBFXrz7sXZfEzETwKk1jY0HOqBo7aJ21j8DsGwL2W9dfEDlA4fPI
Ln2+5EnGun/dO2t0bfqrkYmX/52X0ucM+su+Ugs5YTQgaMxuFrkSEqFhlNuCpq++
gGb2ekQyUELnhYuLH+DdT+4pugxAFRgFEoXXZY6NHahQK19H1E+4giVZGlL7yTIQ
rJvhCUV9LR+Q2KjhDxU7WkfxHkkgfCimgXX55evuzOkmWeJCz+evCxXiUEC1c5+6
hOM5RJ32Tv4j4EMGR+2/jKLAbV7PdOBkLKrQ/HIuYqV1WMhlo+fn+2JFHrmsk1jT
FPM/LFiSWry1PmyRJHgfS0ebEEKA/Ij1kCptFgwWY4fvwrz1xkjMjux2WD6GR8Rr
CeinC1NFZ85m793Ng02VWCRbTPwl2TTSXkBhFq4yvOdsRG/T+JedOF+zKx+ACyJi
qtWXXLvKDSDuaxMsgZ394S1Pnh733yGDwtKKEl6/1pAigH1mUbyJk3l+g9DKo5FI
oQnD1AZwIbi1M8/D+QEmZmVnuQu91BUyArHEcAg9cGYZyl6r7CqiB4gIR4aAhHYJ
g5P5OURIk9hlpxuehuaF6vyO0MHl+NXr7vfyjq3B3tC0DfZVucaFLV1WGCrVTr72
8YMFu9DJKAui3lZexeu62bjoIj51en/m1RoUOq/NPB+skY/0GAA5j5JiCecPRJx5
5V0cI7TQBYh88N1Yqx8LXiG54cGkysey1r81FpFHPLh2tw/qbdFlBwrh68rNG4qL
7IpS+G4+7eBbz1VodBbhGjIwZd22scyDTwtDUyciE12LSR53uYCI4N2OZOA53q+y
5YXxDDnx/61txyOTcGnxO7tq1xp3PoZ50xWeNHqyBhipBoXAzt3LyYoNty435ZAW
SI6HG9anoq5ASImD1z8ggLZRL1avEeELLJjYN3VmaFIQMimCPhQlipn0OEKTwCXP
KVw0kn3X3KKeCj2RuxOm9gORi/fix40WhtfMk/pnbvjiCR6H8pBRkr/enSUVGvap
vBEaVmWMUhs0DU7iTOY6pQMOKK3OLaqInpKgtGtn+6CUFWPBqnUxatLFBDkDerod
HIoGZlAK1tcgog4kVi1h7+/tR67zZxigif/c7tl0J7VTpGgDfHcIT9cKNnWC01gJ
LmTCbLNp7ynHIK99Ly8/egG+8scbf+wM77MBpQtpX4QbmRfDOe83hmmeSk/EhikQ
Q60MGlVbKCLvCt2qU1IK4xaAyDI57NFDde3r3oj/jzqvVVUfQgOVqbk57z3CMqDM
qmUJfO5kzlPxSZA5o/g1O2jL7MPmgVWztK6/bl3ipBrgiYtSp7RYUZ5yrA8RA6p5
rbqQxEUluplxGXBtruPFB9kUXPNFqRrvrJS2b4IFNXEpocpSdN/AZLb7TPN80+3y
5eCOQh5X5bbebLYWTIMk9ruka6H6Zhcs3CDG4J6RdAL8yNIwjyE/ACoTr3PRGlHm
F1Ks8NZP00GDh0qQHm3FCO1OFA8KwBlbFAaTSQFmKfr+s4P5fB1QCcljB/pL6vXV
KwoiXSFgG2fKfjstv5fc9//ev82Z7f1WnXMltEwfumbKRzH7yP+jfDmtybbHZjDx
KquuSK7YgeerctLb36aNN8jTkmwc/aLa5emOcIDU5cSX08FSdthUQvrMRXF49xna
jkhxsMEBujkksB9IgBSxvzfl/19dbr9b29i+GC0WN0bRfSnql9Wbxd/2jP+f1jn/
sUNs8A/CJ/g/V9M+9ycpD8XbhaPVrBiin2JPqQBJCn9pc/NzimwBS71FJABZw2ai
/bom2GcZl98qw8CrNQcSOPYlelgEKum3R/YM0fYBMf2tgdfqQUbpqAMGxIICS6Wu
uykrrquh9pbsEj67IdGLTfvXHjzqlyY5bEqs/W1hVmJWECu2fm2kdw/qDKcypDlR
6393oz0NwAgkRaXH1AS5aaB3H9mdy+z5TrR3k5tkl0T12AiuXRJt9B8vB2YFaIe/
RnnbL54BjA1ZxzqxQbQqaaEf1s1SfpZtaQoJ0g5wzqJfkbiW3qAx70iKAE+D+/ly
tc0USFycybxArCSTheCpBRYvRmpqToaYjAz5rQOjlxVa5WXfFOun31AF+Xx6/AO/
1CaC7dK541IL+h2SlnLolrETHtkL1lAFcJBMn3vgcJIN2SJlPsK7eP+Kpm0T8kHv
wc8yIJ0tPXXEzcJ6eFmyeskQLaS60AhWWTBqshXn1IFRUdl5/+m/cpPBbVrdhOu8
d7vv5/PMcNsbT/6OoiVzJTLAtOAROT2XsjW/sHYfxjsoJ1+pF0T/1ZL6AbZwi01y
Prx4s+Bh0LvuPqScamP63eIFsBhmTtxdAWagF3WcqNu1lVIlvJ45JZbeHnK4J8TT
UkRCtrSnxnaIB2P29Ep+W4THisSz4JdcjZNz0YuyyhvkX9S9NKxiPeVXhYaqgYf2
hvvDjV4t4cgqvSSqc9bVrKVTYx0CwtwZVnb/e+Pmw33yMMlAXQMc24ICM4U9vLpk
d/yxU3aBOl3hdaYgrWKUBQ5QNNCHFmNuLsWvLbVchRgvkWs5PdRj+a+iR5sj6AaS
L57Oi0pF9yQhSkjW7XG4Vt97fitqBlJRiaVrRKnWYYinPCe7GFGqtfDAy1WV1wS/
OUNQKTSCZNoHp3b6OwdGpetADoYDkyT5EIbr2hffgZTDUL7XY3yTut8mgmrfER33
Sd5j/Os8PdMoT8ct2a2GLCzgC/N6cJJkswweW8rfEe7y2uAqzh3k7Pc4ys1M489e
pnXFT/6wBnGoUajGYYpNCDVhLXOznU366jTk42VGaU1C7GIMelr0gWe/Tv7pzXpR
lIWshYW9DsPTi4oz6XYlC61cBsmeF8Gpuyre/0WiHAAapBH2wztWhwEkpDpET5pC
5jPl9W+XbWCmmL/8gnSqxJQ96bv9Oa547KZI+BWHewaK1/8wmiNEgBfSjchKFz3j
u90lwCIv1/O5Qf2CvWjjmSBRdJMiLK38BEI0AIpHbdNTrmSAGrlpzI+axaeanF6Q
gtQ/LyuO+COI9IDguA6BuMnOUE2U8CjT/Yjf1kojPxSc1qeF89wPLwjVC1dSt97H
NAI8PB13ZwvUX3q6+d+U6/tM43l8Re/x0wWY4Ott5xyhyeYhW+wO3Aewe76QmsNU
uCzB/zwkEk60P0mOrQFf2noic0d+CkUdmh1Dapb66/E4v1w4dovjKE9jor2rG48O
AIHNvPGpSNqRDDek7G4XSvOP758Pyo66B6cQlfxfTr5e3gu2WIskAPnr5viHyxuB
3Y2y8wFACBIOl96W96K/B41/7U1P9rzQdQZDcAhBDm/9dVui1e0Rz/rlMnfgnFDn
z86xS+1hkyLuRmjliPBn91D7+lzVgZJ8Qj6N+mKkU2mZXL6OLhQ8Q6q8IsoR7erQ
Fcd7CcuHm2zUo/dDBwrRK4u/I1UV2aVOg11X5TQZZgq1B9yIDJ6RsnTnrpzDLDAN
BS2Hr7dkAIz7nOFOQ6Q8q3GHiv2XmUw0UQJUWQP7XaigPtidt/WDB7T7/efQWux+
JHMsOjFLwfI6UCPl0LxOnWZSCWtMGafgYQFKUh3eVYezCS1PupMFQtpQfuXNT97J
xi+2GoMS3FwPx6LFukskcVRc5LzjxlEuIDYAPcOq34rT9UJAD2G/1cYp+ieIc9F1
bxLjDx1vdgLBHeePYBSP/6gxNbjSvkpftE+0f519eQMHvNKTsURgTeJtbcf5lBaj
rJlTWIZmQ/VSxUHNpMCnHZp1sxYXs7rVi2yrwu5KdEvM/uYwb9znFfmUM3L8aeGT
sWzgfB3UDFDLwnFZztX0sC5YiBA4VFbOjpdyjjfARmqjLKukwypZSnuiZ07LWWeJ
gMNae/iojB9FTbo08dlonUR2We4+kkvny7MzrXNOSIVoIjF9FVfGzLCwJejP1ZpU
hagwsN0k7PuYA0/U2c5psVMb7pw5hMSGBrQ05pxkMH9rePZK8HRdlKI2oN0wuxxB
YDaq3uiVY9Ll5VPQQQE2Lj/sKw5eQe+riFUSHSLgzy92n+YEwWzyfOo3BMiCmO4h
DlT4UN0Y5Ftmm1EX4mi3xsdng86dRip5oWObQt130vTD4TMRebZwIW+pQ9zQH8W5
EA7RyDmZIThv6IVQ3i1KPhqf258VekR2fsl4BeflZyqHqRPjtyXeFRZhJZie49zT
DPiR/RnAvDF/cwvnbtP8UojfzMjoAN7ZT3vJ/rEbhNIswK+dG/PslmaOEZ2Xb5Xv
8PlzA2FeVdJdCR/r+cXkz4xMDlzUjpk6liPRAgbhNTplic96h5V50XO8LnnpQ6ls
vhHY4SZQ7pQdEzFsy+ki5bTOUCFMCtwL2+n4lLgn+XFDELNsbpHe9Kqe7EgoeYz0
QbiNPFPDuwQQUO4tWXrA9N0kAUCUDjfJgmSvmcaYUkKVzG3szEUq6A4r4VjxtJFx
+e+DGbbSgnSkoweJk9GG8uHuKsGq7lBQ6U06dp3iqmjPoZ1uOQqOSgm3ZYzgHj9c
xnmc8uqjBCAdR4hA3H0evGvFJAbWnMK/hQ5iKh+I29hNB5kf7Rd+vk+sGlEq45jz
ZNnr4ORj5Cdkx9kkSLGziR84v5Htl3JF+lM5BBbt2nuKBawgJoSXcERImO1oiQ7p
infpArZ92GUZCUMDQB57LWY3GipwNcJGaCZhZk8Vv76Oxhdex1PdcP4IVB409vLO
0axKtIAOsj9JbN46E7h+gcuOmU6u84p6in2sND3hOswYhylpJf7kZ43xz9LjZayk
UnSIqA0Jdt+dCfulkTdUh2/qsNkIbWNgXgCicj3vYVJM7brEQpuRhxq3MKTiVQgO
GwuYYhQqMrir+O390oudyZXmxY+eXcI/XbFYubaVY9ybmwFJUVDANfXGjMO8SjrB
dk+yb8H1vzu+P7Q1ePs6FriVOJEIEc3eZuJ+lnGR+pzfmv7ZO83FcB94hZK9nnyc
uC/eT8x1oqotZMIYOGWVvGdR03lj3It12wSvuuUYCKNdZE3K3K6MgAZCx0YVTuOp
awVOSEO8qOk8aVw+B4K0vMz5XQM+XS7ZcNn4hf6FusrK5nnsrW/tSGCM9lFEa/n9
yCMISTi0Fg3hVYeS8Yt3ZGevUVywy57JpAdQjpK01v4mNZLkEyCmt+B2zHZ4I/WA
pjwQXUmU9Gk0xrqI5N7r7TWlW00Agz9ESVRhHOyciP6a/BjerDEh8XsGDbBoNyp/
ntrxFHLtTktaiOVM24UDqXAMWdyRH5rTMkUd3hnPDWRycSyfsdhlVudEOYbBodP3
IZ2PJwwYZ7F5itEB/8bzHwbsHbMB3aI1k5pkKQgPd3SQH/eAV9GskQSIBXLlfNqi
hhnUz7U4bQgSTc9gtcsOJIMSTQHlJPecJmgOEvgzR6rq3//XpM40MQe/g7KadopV
Gr4+bBvjR0EdMejpofVturfOcFrSxzVve1Ld6qS+UHMJBQcofBHdv7NBCXK+ZrIS
TDFvQeCOY/Pv+xY7sYJ8WooBBogg/0pm4H7CdSADU6CWvLIZLmHwJGN1YZJDHqMi
uHgEwf/tWh7otA12dK9Kz9rlDm/7ROhGhTh1NzQP8nef5X6/0tTyvnQlaWYynNuL
QovqC9KqAQPs8yRU0OUuGjkXvQkgdl9WQ0lAtS33QcY2G0siEVGCjpcIl1S4Ot1P
UtJ5SMVGfXrZWqvk2URDpdW922VaM/H/+WPyoGfvt2R5wMhv82PzRs2q0W97uATl
VnTygZmSYfTNOH2PT6OB45c/ofu91PytSjhqk5U9/PWV9ruYz3fe65PsjKNfhl5x
btlroNdsxoDpUuF4CAJ968HMc3K7FwbBIA42ac4vHfvcys878/ZBidCsvDvb9cH4
hs+h0dkwoI3wA54mDaJ4L378jvR8pE1S4xlQjS+fqz1oi7wsF21by5xad8nigqLX
8uQ9lRwhwlu9vi1LX9sCbyAbtr1iHZx7aUo0Gj70CRNjfvOuqsMnzNxxeNd++kjN
rOsH+VSUngQsULG+c37LRPjEoqEGjbhBpwQKB1oGt3AWUVqU03J7N6a2RwJ0ss+J
To8tLhthAgvSiPMrGcjNgq51TFRlRUrpaSRY2lXWRW3YOLw4VnqP6Fl6v+q33ueu
YA9rv4/Ifz89y2DQei7LyRSQmtTf8LQYoAD2QGYN1qU2cx6JvdewhdKRILwDiG/X
2FS00jPmqy/G5dHnoQrHZXAqsyxhsfGyRxHLRNgmUW9vwMwr8uBrAmQnrAEclbDO
wVLkLolIi2YEZZw8qZBsoW+IZJX5U4eybkyN6t1F/QcV3wPbGWdksLAI1bFSUezu
/PBORu+SXzsoGEyXxbvAL8a70WdOfuzTa/9W73vOta/spuB73JD6trXRrT7CDAJw
rUF8TvruTeC5UcmqnYM/pLdRnDWRKCtukJysqEoqkmIforaCU4NzzTXMTkF9sAsc
AKcpaB5J6d0JIvXEN4E+nhcLjHye5o2N4qY+uNdTGlQQdFjnoNXix8QUIF7llNBu
uNckTTT5gYFMS6kNC9h44FOPHDri7eW4J/7WOQvHxPjSN/K3WZGDGYyiLimskEmk
CQr9objcUyuRf6F4fl52niMmbhoS9HBhngKHFRLm9uDFjhZow11yRJV1NPYOJASh
DcLpe2iuaSidKglixgvZxep7a0jf73tC96z8x4ZJRlOKeew5GGArXe1mZysKGNys
RuSmYhWC8fDBUkBcjrhE+ATKz5P1MCFnT0zaEsh7kCWlrJMAcU4Uqf70/uGVGg4y
4mE4eQyVHGn/ba9vMIy8WRudR8VNmtHWhslRl+B1+FzbmYpYLmz+pDGNV+sZVFAw
o3b/Np333FTC1RRgxOneWPd/4dxtienr91btaiX9Ft2+R2pojdYd4x6xPWTRVfUo
SFu/DZaDhCeSANuhfIdGNTKL+CW9oXB0O64FYWiH5oOPQsbuZMuTea8IM4V/ByV4
Tjfa8Q0I8DKtvzwHILYG1w294Z3a5Ee28XaaGvBBuh0NWOJzKR95zLZOvq4Z10Qn
FosCprMvci1jmbOPYpq7Jkbrh51WHcbquKMQX8o2s/fByKYjw8HkJekjhj3y9Zf7
eKq6bVkfYDfWqxQQGAidK3lB+muT9FtDzponIiTESCjlQxdSwrIJ3fFm1SqIMkR3
ai0DGn3IkaiPtslziPL+Lsve75P38fB+HKUoaiq7qFWuybV+BBUtYbXVVPQGVKbO
mtZGuXdb+65iximngbU6u1TuK8qfrzxu9iLCM0UwXkRroMOqmAmLsRgYN6qLywpD
gAlKmVNI44KmUzU4iKivzHXOhZaCJ0Z1MZ/vEEDygMe8gjmXwY/yt1Us725RyDXR
mlAEYkdL4JIzgQlHFmmWfDuDDDHH/x+BbESSU+8BxXCPitqbLMEf+eCAHaVCRlIu
gWxa+LlAShy/QPBic6in4qGDMZ6pTC7/q65GCv+uxl/9CkANGFeckWwSsY4xyEjR
dRs9ErxDahB0I3KT6MJtYKAVVxJaiz+fnK/vugSYC/ha04VO0KAvSGViRzUfijQK
CK5PqalqHbni7mucAmbr6Szwnwr42kRyX9sTFzk40nQfE5n/SqwtiLQUH0hSMAb2
awDmOVGFhHYlIZMH1xoztLASs8Fp8QlZLcfh5Cw6YHhAbIuqUiLFnsm0CPNEibDw
+aBWLDkNvr7gd7clFoEBiAn3vZdpWl8TJk0e6J3I6tgqqo5/8SzSA67dzXA7C9qO
M7nby6eS8577A6c+egMst/v5DUJd32ZREQqhvanu3yO40J2DXLlJgJrtPOEjwsE9
pzVMvuPPWDNQw2ZYsrQDUohgXEs8sFV5LxfCB1pbmR90byHSvVlcSycww4xlVAP9
3w33ae9QUT/LuDrqewv9QHYuWShdDYzf2EHvcWvkDn6vHkuCnzdxPe/i5Q4DE9wk
nPI1clTAPuTe6UXP11FNSY+mCQRYQA04nC6usgNrOqXbbdXoIS/Vt/okr8snUNhK
1F6kkbBLf69UMJiuJ+LWYOEIgSYzbydC+0xrMFclWx+p/3NLIDqMNbwb6s6SKLr2
q0BrTfC3PcF4nzJuV0SG5+E5GTpxoNRG5aDAeG7smT7+BnoL/XrJ5UbuTzKhvWZ0
rTCsANd+p/phwPUz2ik6HLWcZJu6KWKBAFFeDZ9xGQbeg7Og4Q00Iy+pWzyWCDRL
FPt9824aWkxNh+oV2ADVbvKLFopPm2OjiIi5BrJ5WHBVDdeEQnTH6dPaH4GJE5Fc
80kezouGAtEiRzkriL4ELkA4DTkuqP/GafXzPOHdD2tFHqGNC0TfQlAofr0Lb+YZ
rwTpfdP7jebrSnK+SQFkovKLI4Buw10tAOLVAQj/6tH1Xtn0OZcoaEGI42B9tbF8
71xvODqZ1W7BKYvRmTa3gVJhCZaAksxnoYwIlntLULr5Yo6uuwo9tEHqMyQqvcW8
rH9be80/htsiB+Yaig3HrEzROd0wDELrilRrVrAtVWp6aSNMenUO8pK908uCoUTz
XxJyuX53FVYPGCI767oL7HI/IPBPnnqxHuulKSmhxXEbQWya235uXksFI3jOVWg+
gLRUYEpuHrCTjuBPQcq+wgDz8f+rqJl37kusM3ZdbppVd3Dp4C4tmGwxXGVa/eM7
3t8rDqPhizl+530NHUhSTfHHRa3DCJjEDznA4ZB3/eoHkrKbs4O3VJZDzxgiLbpy
pa2ntpUHfvg+TtUwF5HAtAe/7XFK/CxZ5HV/mdvMAlNgt9IXFkubnY0xznJgOuwy
7zfXZ7h1KFigTbXmfrHppx5ru1LRilGupt7y7begd1mBSP1HsIeYT8Bkywgn0Efl
quAT6xAAYflkuQfe+EUwUrxgXbIGwUVQ3jV9pnLj61YqXxdHKbXUoUUPqUjjEb6M
lKyOQMyUn0Z7BcdtiYE/wFhQ1pWeUcxN7s00VrSOUGpG2AuhoApCuTksGAPkd0uA
tNFdTRiUWA7mMmd65q0lDrbc1wtqd/c3tWmDvvc8Dci6tGLJDY460pbnl4tpnvAE
hAF6pZ5ifGbFZ1NBiKEE3NmHscfirXmhZ5763IKkzEm4czMSDMDwBgNI5mlk1aCJ
GtnwsQkYlYDxodGDRmLw6IkH3W5IsvUYPYsF/ZYxvuCZz3ksc5aN6mRvVKRxMUH7
0S9+/H7X48eBd5VfQVNmyk6enyWmEDwAArrHqe/NPYkk2Uur9RN2Pv1qD+AE7b9E
FcHmXnr0aakcnyq7JzSsHNkLaAgulFJF3mwBaZkvy3OoLeLl5OJB7fbS57QCl1cP
08WwPfgRtH+A2hm8YOqWXhSJA7nTQKgrs4WXSMhxeXq71QVF58KlERxjPP/liRy+
Kz7ITy21XtPGb40YwJjwUoSR7EojZjb2Aaswty76wYBKhzUhP60F2c0R0neOYucf
I0gTmvHsJAk9yeIg4SYzpGzrIV820GMAFtjCsCHfIcR2JTkUdJZdgYKtq3DNyL/e
WbuMiExiABCK5SIcF7+MaLdIeh+TIQ2w9XjqTt1oElymn44Gn2dO7MXRKWpbWiwx
C2NPsSd6ddlRFa9Cia+f2Z5bin/X36KO/OyQFprJR0UejvoQ6QyjqR60lYrlT0hq
6agq3frudBD0wtHN/H7OVf557KkgT3m0y/3w4DM5Kfl2VqzpOsRQS6RvgzbojI6C
5bmJZ+u9AOTPMu5b46gCVl84Dk0zMvlchO60Vg9NU4+o+OT2rYzqq4Q8jFyhJXal
rcNNNxCCN7iNipOM5x8JpH8+OY/5m5ZVF0PXxeyX7EToVLZ//hLhl+WBtXEZEg1N
lM1piVMUkPaueEqgG3ytAgEryNiB2T8dgq0a2dtVDPL9s6Tf8e9TL4HK7zhBqGjh
1nv8+6XTInif3qAxkltuW92iT8aSn5y11cySl96YBQfy2Dzdd9Oo3ar9kJCGtbV8
Dol1atx8Yk7QTv/1bJJl1D9VLsEUAnrr8P4ZVT241j3oEQnWyEXQRWbvenKr8CVE
4mt7ubGx/9Cv3uPSLG8YwDHQ6yFeqIqYCxWKROer/Safx6HkobNbTxyor5Q+k5hV
4SXsC0bWgVaf/kVjd8itD0TdC2CdSJ6nMw7mj97C6cnhk/w5OIlL+cvZ2kROLlK2
TRjqUoos8qU4T/+hrCe84G6HAcpClHyqtZyBCu95byJdnw98/Wvf2l5SVsQAhW76
eFlprDL5JX70x2862F1YQ8TLMhlZykRJO1l2VwxQ+CURfiOxOWJHsMCKjrOgpMy0
t7PYsx32eZ6uX/mWpgbRJ29AxvPNqQxeSLLtTccPrqQyTTLQAPkOJEMDZ2Hvf5OF
AW6TnJnORi29Ts1Z+QI2JpK7Kl96iQpPskow/l1F/QTHoOoXa34rcSoZRlZ6X84T
mGdwiDeODdUqMMwg4a+BiVTpH3vOdZ0Eq7XN1wKYNuPX+rLKpeJpfmrqyaG6w3d2
el6P5dwgaLS3AYLn30HG6XoF5YVsjrsDAfdwKRfO7EJ7uYMBrFHTVe8dGH3BtgqJ
hHdg20SaBFtJjoFQb2XbF6Zoed1gzofAVbJnVFvNOc2zvfVWgyaj3ajIM6FUYmgy
LVnp+XGZv1mT4jzZUG5PUIEekuQNIuiXYm3pp8PExLAha64Bw5dVxkleMii2mFwH
T301mfzPMaaezQmNSTB6it0e7tmZBUhz0w3HDft5qF5F8pMWyMik6Uzcm+jzMNST
8mLC13cg61nqRYPD/KiqN66Es7A3PAxuVCrYsWW7je6LJOlqnnqtkVYm4Nufehav
jnLKLWHDVZlt8Kmjo2NT6ZnnX7jniLGvvdDFu8VhCkdehmKCANLvA6OCDfl51ukh
Ev3nnq7GgT5UetmlTCrXlgevW9NWlJgSBa5BINaWVT4BuNK0Fh/zHTek3pxtrjaw
S+Yqx+h1Cqfq7HinSOugST69t3xbmE9h4f8YrNIzL8FLkigdwPdGNWj8tIA6lIBW
pGUkfzi25fqrXe1L8CvdiZGDZu/qUgBJlL770gmTefPFjTgNHpqa+O6CP1RVi2aE
RdYEHuUI9tQ4pL1/AbbKa1mPGfuUz9D1MawEEsO0LWdxpd7jvVJdjkFaXJ6PlCoo
+sIIx1sGOqaf6gLTqetUGB060otveats49s3uSmpzHbxVxu/EOkPsyPBZ4bSBJyH
oBMQVrX+KrJtU7IxGYKsB9QqdJR4XI8PI9Kuk3KCFotIR/8q8WV8fXUeITuPrVen
a1OHApLCs4rMm7O8z4Ft30tFWTN93zdJlIBUMAWwTfyZWDWlXrtv0bOMgWIPNy1f
WEYh+aXSAbU15eoWsqvRP3D+OnAKzH6pk2ftINBRlUZMLx1ZDyMTAVW7rxtFQinA
vfcjK44Zb1Kwzd3dkCU0lfCpvyv05P1DJaVrQ+J0BKjtnYkWglNXHuVKsnmQThsc
hP5AKyd6tuFytZ4p1q07uipqUFmZ1bE4HHVvvUvGIh9N6A74gM3yJb5KX1bRNXka
YLKQBpj5UTdAgDXWTWEb6A11dQb7V8CNIapLbiYROdMX6Lw2J9HSLxCHK13BxOo1
WJdPPz6nqZg5ZfyvB9jxNhVTndq3oCodhTYuRZNAeQrk+Vp5X7XNSnZjwpyE8FHd
xGqkcrWGbjW8kIIKoyKI619XN3E/WNq9gvtyfVfiO4yPR/h0hpr2Q8VTEjvRTthc
N+bSK07LPM/FUjwkcV48LJADJdgoeojs+QJH8Z+mt50oehDbmegrwrzjHPJFb10C
nyzqFODx4fNV20Ih1PYkMiyNJJPraxsyOmBQE+ECaHEM/gUOGM+0QjEQsyt0jzVV
KSoU/StYwGN9HgkR1wNsaFZmQdIyCNTJwMk86j3DUI5yeelt7hv6OZ7PdyMGbCzz
S/LkF4YwlP1l9+xxy713FFk1ARQYJJPNLOvd3TVHcSZiKV64xPE4Enc7uFfRkTzl
lCoQrJdkVo7frAyw/jo12W32NxEPAiyVZJxJTpw69btEtZt8RIaywuGcziWoEBN8
kNW1aJvTuwp3nFq/hrcYYkpEs+dx/9+XZPRoujX++wk5+IdqW1A5aeb2aOkINkql
VgsXKNol5adr6F2GepEMaCaUKGQBVIvbWGr4c13nc4EEewCmz1bRJKrvzDJtJeJK
n/xPpOOIYySwmOhgtVQuaDZ/ckUUD2WCEfDVI8uZral/kSupls5+FbAHuOIlldCR
K2p/r4VNZJ/GAUP3JNJe61iCsFA/rzkP5yrELZFRU81AYEvjTOX8qdoz9nv7r/vS
nx6FZAR8rDqZTuFUEuWk8Ih6LXF1KDxOfevTAQUsFQ6pV9CaAuwDBchhGm+a1p64
SBvTmWtCLN09vl2ESCQTloIQAyK4VlKcpeU1RKwTd1jyIScfdJWosLrLeaYFuBgK
sKZhaj/sWUqAdGoJD2+WdAVMv/zSyQy4x+tGCYNJ8sCCKO1fyLfmPKJtjhLYCTbW
JSkTL1C27ZwDD+U0gwSo1NAIhlVv2sQrxDnIUt7Ryc0bYeLJFzHTkbq1+Vt/E8Ko
KJ7GDNgDAwmj1PhEdL5ul1h6AxYbKtW4nsAoxYDZK2dwb22oO3GwDp0Li1wopFPF
TQqdDYOZIxpYhlTRX+gtjUEKdW93sKSwtLkdpAs+BIzluCGupcAOjgkM35mfOWC6
IpmrQP/SzdgNE97A5WDMcNv5xchN5MWNyClQ/gL6JZguxtY9GGiEpscUk6yBoZMD
VlytBITvbMnSuewVIyBO/7CiGGgArPUVYsGHbCAYDxbu3dXVcly5NV5CwM+SfRjj
qWXY3s9BAlxnnprjel5BXso3iIJoHEISmFqku9+vcg8EnKyB3ZP0i0DElPiE2md7
jXvP+qEfA3y3eBfvFsqDher3ana6Rs3p+k3eJnk3ABs=
`protect END_PROTECTED
