`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CbqbryKh0HK2EttbV/OVjzjAFbVnTbxKP6g/vOGo6DyXjccE/mdSODYFg4sf5LrL
SYOQeBOM/u/d1xFtFXN1WJ8n5Q+CtKVVjSXV4SrdE7BFgZVu1HoK4YIdPqsCJEmN
x6iJhvH2bY3t2jNYfuFE3YH1j4JrCSmkWI2MLRAoIX3APqU0bGgzVWy7dU8r1pIw
Ll0BODimhPZQ7KYI/dmG/SNc9YSBKzMsJSO7mv24FDrQvPdWZKqbgMJwEbylsQ5M
LU1EwuCMSQKEbFWTQeJN3n+F6EsnamtSwU3A/37ggIIUynmI57qc6ZhRO7pBXAdP
AtiXSCoG65yKNL4jroizyNv9usqTi6VmGwSFuafjNBaI7tAkwHcZby+Yo/fxAffz
aCwYZrjWZgE8a5f8apOuKdwY/WEC398N9qaNPirk5S+7ixEAfU/40ixxChkRzZMF
pZpkg+ryJ0e6uOT3qxtNt5R+z2wrRwtd4CUwkVP6mwD3lLmLzHZ88OD5NdunGtfB
d7IC3PsFPw4Mg07VXZAUi6OuM28YPyW/E37UB/ZmKfqR3oNQRROzOe06n4cn4lH3
N9ab4J1P0M1wsY9HvKTAwjuX4+KffmHGTJQuMy7pGZSDel++TGRqXTwWp3H8Dov9
rRJGq+QXDQc9xqRb/bOjr9Q2Xtm16wcZAUQPFnCe4KxZ2U+5Huqy3vC/FGneeYKY
IBmbV0p7CAmPepeYRjbsOmxe/C9RtZeL8iSfhHeaOIWxTPPIfmko3aorCn+QZ7Mt
eLY4xpT6VX68TKaWGIugzJoaHz2gaZHhclch+H9udOFJDyLe2smae4lffKUER5HU
z/sNqjvf/nJhiuzAvM5eEhvGXoHQrxqETK3KI/VvrzwoDsFEUtRjJFejaBOVyzHL
OqG0hhfYZjodwNuEDzBfb25vhWLbllS8BPmrXxZk/B/k8kN2PkvuOIH50UIUK7gV
v0HR28j1Q+GA0pdOwJyIS2cmGs+49uPEj6PIgkaNscfZlyhWJcIskcpCuPIwv9uh
g8PDhqzkrKWVzXrSNZKKPQgWFTwUSRMV/GbTqEhZ+DZNt4f0embBD78F8x5kHv2S
WaFnNWvZZK1u8z9byGsBqMYkzc8Gj9iz6q7qc8kZ9uBkMU4WKqENBqGJPiQChjYw
`protect END_PROTECTED
