`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xYGM7Nma+yXQHYmBz4MKrjrB+qUDtyPAyg4F/QnXu7upkT0TCUqT36pC5QpGNlOg
aXrWFNJbH51i4C4k91Js1BSB5SmsRfc3e/kv/bu0306Cz3R2rplR4euruAOMpWY2
El078065P2pkvcxd9Y8BAY2SAjrNUzXaebI2+J9HlDQ8obkQv9K5wdDZZf/4l64U
I2X/pEXAikdrmWRHWsVhKKTK8lIXqfi28+Vr+dXGQjPS+J95Yu23gyBs9adprZ7w
IjZUAcdpJInEYzIl9g8cT95w10bqLul83thfvj2MqhrHlRqYZD0YjeCoP4wXP/N9
EHR462jWge8NxwBZhemxEGkrQqoktaEafSlWr8hagUK1U2r9x4jGrCLfgEkE1Ta9
h50JUkRdHa8o9xkeBcUSZe62QI3SjPFFRTTXdOfJ74TVQ1wASQ6vkO7jot/pkWcl
7+8fUXFztHOaIqNqo17bJxYZSyr4GTDFdSfxf/EdgIz0UyEGcBVHyWvL+2bxnWT2
e8iyAOtdksZcaMrPeEFf0noU3Qd1RNZTma9fZJW8UmZt//1jGFtPBzYvSIm5VRYE
Jrvjy8wFmrD5bDKRuD3V5lrRvyhSoZ5Oypg7TY0IkIFMimOJvaEfGc9T6tyuMjAk
FJgKr5MjILhS/A6J/1M3VadORdNbAn4WPtFnTFPryLyKZ/ba+ZfyCHPLBijMCzY2
/Osc/RtK33n1av8emgaF+8vjiARiTnUIA+34B6y/Xl9WU/gWjBx3cWDcIFhCiGxE
Q0tfgTNQ842JKpw97CzizPNHutT2DfD6/s04BzMbIFL+bUonsw3/xCLrp5nbirow
+QLjsZzYvZc6192ltDJCct6FcNJJakfaGZSJGM6oinxTmAtq35Mr9au0Vf6LYQbo
Bap70brWG6VcCfJTJ9COssbGeKHNJoU73Wg0Umfyrr2FUALR0lj2JPbUUqCKn0Lz
UaN3ahLtCxyNEiNVhvpuOTUeduuzgk74Kw0KgJ9RZ2k7SQmcbY1beM0uByl6CcsF
zFRV77koEO+D5uV4Vsc1fugENePjvzDXsl1/KcJgoQGZ86gMYF92a5LNSXcDhHug
Zzk4nk6DPxhp/gb2njzKuuv7AgVgXRNSEHWaNonC0m+N/gSfZK4kuKTCQGtpbqJW
Jj9dbUKjZ/8WN8eLEMSW7TPmZikkqdPE/Y/LpALZGEZkcNE1RTu2u9YreqMFq3+y
naPyLJ/I6PFKEbBhS0V5iwK8qtkpyoPB9tueWtk7jcDkYK4QHhAdT3muIX4EDYVM
YZb+o9mSPNxU1MP8rZuP6VzOgo6Gq/L8fHxTxE2Z0278rh22LTvwvHPDFExCUYuT
HYlerGQoKUH0vxCbsehSE7qnPQw3gYUHwZ2OX0x4U5QAco4aKNTvTx/80tWmHQbn
WOrdxb/gGCOO0nQpudjL8yATJ9h5OcadyoVDyipj/0i8Id84oaE8/ymp3twyjfGZ
F7OVe6ABvmxkeqXtwZj8vXfTJCGPar5q7N1r4CPTBUQMmsOl9X1s8R4J+OSV4ArA
1ey2F0gP4XcoQd7GHZTdnXpmjqNn2ZZMarsNeOv7FTWa1nwDHTRWQSke3O4Hj77s
kD1JakBRpdjcjIJTZ+6fRTDJoQpXAJVsBV0Jr2Ea/z2A8N3weIdgWW0IJrVnMfNd
WoQGBqGw06+37yD5d7GiktEUQ4Oe2QHd6+vKsGTeXQjMKc8FV/EKzWBSR0G9px79
Mq7GIemaQhFI6QGsmaMAd9JVZhMSHBo7XMbp5dJku0s2XbPnMwKJZRhRSjn5w+RV
tOXKnA3NSRdPm4OeRck20YKnsiswkfHVi0uH4LPe1pE=
`protect END_PROTECTED
