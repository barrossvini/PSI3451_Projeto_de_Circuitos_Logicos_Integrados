`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f4oXQTT+PWzg3Bv6BJIve18DZEu0E6qxKua8XSsOJ4EP4dvFz8RA2VuD+fXLJxw6
EgW+/QUAlA+mtxaeYoQddmCzNyHXsM/7+6FcIEEUN8CYsWoMLhYlRBpxRytzqCFA
Bg4GMty3N9hcIYPwB2IVjjq2v43+L0mRRWYB8ASrW/1reb3zbpL/RokjCalvQfy6
4+9E7kv0RjFyWNKB4HK9v4iVg7PWI58MiHo3jzBEJXhTOi8xNgbVDFuz8FO/llYu
SM/wWjzND8+d3fa9TwmVBv/34xocXmJS/usVduGMAY6OQAEIuG1HDcZUdgfcL9Nf
4M0qYnNTA8r0lrtkx0TlruL/hZ9GEo7BFELecfdSNV61DO28zl8I6BtgUFu8kE0c
yV8y3s+sQzTR18gz59SwD1OjYqkJsH9dDHFZNwhREHg7lo6SDPkY2wvrUDBi0hAx
r/wRiq5h9rNiH+L+bjeHP/4y20FP1OxsQwV/Dkwkip6q/u1njZIIIUPG2UrC6wtu
XXdPQiGMx352KeeketHL6AYe/Tz4ROjdWsEYOb0+wMOttkOT19pHUGn9QHi8dlQX
l3oob5GtxGv9NtlEDTBaV5jckNSp9kW7lc3IHdz0zEnnjrh5ss+gib7CJbc5Usy8
cG9fIRR76gUxg0WT2KWvyavsJW64NgmhjGMD61PI6/ZlqsgJ/xiUeYz1tcal0O5u
KFAelL5O6XjR1CZWnVmTQRCNKgPZyOTPNeiZAxzM0UbG3lkFf84r9mlycalCxtLP
6rKc+WAMc7OaSnK6a9LciJIhvnx34P0K6W2SPBZQF6jGEEL1KQQjlCucgVIiwnjs
TogdaYBaG2cH8LlhCjsbnMIQt9Uy4yY7n1WIBhr2n/sHSfuOxi3MmHIWjU6IHO60
pTFGQbLT1hPhVguyS6LS74pqJ2vAk0uSEaYBeKihCqeE6Dnli5BUJfb60CDqY0zJ
ZkZEGupQLjQiLdRXXt6w16r9B1Kbku5rZiM3o5+Ctzy7Y8XCgEmTC11fx/Q8jVw+
lmgW3gjoIPKhiXiHkM0m5Bd4rYdcO2EO81yHdJnmnnxzFYNHz1RD/dfl3TL/W49M
syJn6/awB5UG+gUx63J4/ATET68mLwbLxxyvWYYPHSTHHXPmv7+CCqqm5Q6k1kHd
Sh0qN6ZvPRSafkuVbfE3gw==
`protect END_PROTECTED
