`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B87J7V1o2b4Zr1apCAHY4OhmXAvk6o8KyrZV7vjY/u6N5wx/itmUAao/UV5NJmFR
VGg3JnREVVRgBQlV2UkCwDJ4Ers4EGq/DgqlxVxsmogWrUFZVWFdp/VyEHzMJANk
F+G928E7nqGWakxj56j2GICJIGOaq+XAh0/+gFtlQeXoyGRDvccW2PYuCPEpMzZ3
ogwF+M2dvtElzp/IUbJ3NqClY0BKwFATSBXIwP4Svs0VuelPOProaujcelExtXw8
4bWO6rcC/VYm5769Nx7siMHn3w0rsvGa6pvvjFkckaH0fw1BWgAzalbAB7rc4k7+
blfn8zcgBpnpLu054SO+o3lgcAFG4r9qjley/nQuKVUV2u3LJsV3Fd1j1ALzB1zD
MG7He74e+r+mSWK2l9my0KDlaWwq0SeqG8CBhkU1DOHGL0ogNSMYTexibKSNuwSQ
mlG/rDiyu9PIOTE4zLnyctddqDHYnGRLefYROBaP1jpfeBcKA0M1nIoGzno4ze2I
2elRctwLUEfNzg3OpBsKbAzsP0M27xF/aJE3UCnommqmB48X0uRlYw7Vr788hdRC
sPFBGI9SNcoa0eAm5zYMHW7M/9oEQX8yZejhhZUX5rue1niqMGZdqCshdf6SB191
h6hrC+mqVHoaykFiz/6BlClAvXBI0hkITDwW0shpB++9Fj0vhGNUfs5iHGXtk6OW
1fyl9kwm5q1J1PFRt563aQuG0jw9bNwzrXqtWDlbgUD5xl+UuhfuoMSiQVHJfcas
cvmc4/hbZBJIcung7WWdztnuUkYSnE5/MkNm/YysLpUVs2tS1szDgtaZOTdVe0TL
1fWJE1jv9ELVIgXhGkx9OJWdqV2Z8fAtczsxeHqa7Cdbua+BU/zyHazqbaBgXNeM
07N1InOG+p8M+91YwBlEkXWdE6xsfEk9QNsDtjvcjlJjb5zv7JCVlVFU0QB5Jn6K
EtAiD4x+PV7F+xDqf4CmFhwZv/lZl88Q9iC9gOvTtFiwv7rBPIpb4HIt9sonC9dA
li9UWyYBxHLRvUleoFdD3+/leqjLSa2ONSpQUdQ5LKUzxOwDDu9MJz/f++FXwu8L
xPVrLn+CbvGbTs+9Ny6sl1M5lCgBjVkimd0JbBDVA1JpGWRjZMC39h+ceAMkhHhB
lfJA6Ofne973C5pmBgPG+XcDZgqBQ9BpQrtzrnRq08GmZau0SWAcSpx0iPoHMzpE
0eg+Of3huJ1mCPS80YJKdh7vWANiPU43tv6vtS9KFvBMsxWHHcgML0iQyS4Yx/zN
xzP/xGlBFBTqPGEs6wf1q+gjjGZyCm01lzfiXgM/UFzdRSqTbJ/QHhADsg9uR2TP
wFyhVbBOq/ZK3aHOihQM2GtsaIXkP3lXMg8tgc5ZzFC496B+eEmuzcop9xFm6dYw
wnnlQdkk4Z0Kpw+5QqLEZcEpVEZ/H9e2xiPfErYrstMdHTRO8IcghZ+n8VxunIRP
h9o0a94SCnD6PSldVfO1lK4Qb8u4QTQeuVeMWNDFkGPfwjVPDFAaGMkJkYYKefku
dOlT1EqTbzTWkuUDm2N9chy49FJLuxQ1mmsGeLQ8tkiFLTWGrXlfh57GfbNCXmba
VCxPvLeSeqgaTi5SLwyt5Ru9ou58+D9ozWBMKzTCf2qCWL/zLEq3Pw/zMmPBQZ2A
FAhAOGNkzknV56siR7WUjmca9wWTwIXENA7f35ruH/ecvKOG66xMEPnn10ux1iki
3uqGyn9HytvuzxvBXIcnOiP31nM1nxWngADGKp67yMEY3BLehHpQ/909l8rZPQeo
xsQNhDGUlMtbGPxwvgngUs+r868xFt9g/LYazhLwWCuc/nZyybOokUvh80TR7HUs
wQJ47fIi5aanIdbysEPOSwftldIWqY+Nc87alqEYzXQD1mbIVqxu03efA/+hRy+6
0JVSUOGCP4LYhB3/78PV8yDdKPxwoiHXg1P5GAbVOo+jsiLEKTOc/eakkla8T1k1
scQbXBWQTi4j8wmIVrJfuk6uNI8JHS5Lyq0ALl0XawDicKL5H0HOVJrCVxfzxC9V
3kwRpRrG25J91la8G5H8E+IRD5jGaMdOM/+c6BKpx3wT4Xv3lSIB/G25IbW+cmF9
Dg9oRq1hirAE783qcq51aSGdw/YLD+17cji/KlVDuJjNGLtGzb/VPxXf4l7qoJVJ
k9tJvLtWD13VLNpgL9sDsujn6ZNkv/efB/deALIpmtl/AJjxV1dkSeg10qjWKngx
0R4CjvGMcQPvUC0VIoVcQKF25E+jqmdUS4957cwXdFraFSgw303uHA8pBb52msFG
TtH3U0Q7chvwb0vln+6CPlUH8VdmtXVK7lfZ+Kr+dN+vUGrFhdTUQuJ3GVjUkgwt
jG3MOkzT5UWLeMY5JM2wspnI4YBiEqWK0VXQLSu45PzuZPeLQ3MyUfLubCcTc9nf
c9BQrUm2H5hW/BN1oPX6/+YdnDZIDJGKBf9eY2didYbDXoC7uyXdyQ//DvWW97OY
wTSWEROHeaNfaykl+gxbmaxvhY7UEMcvHRoSuEarPulGAJrnHuqKusK64GDQTUGG
YQggi5ZJj3WBWSSd8qp8va0/zxWdZFDylbPIpr0bcisx4LshPFp+4MF8akvdJOQs
/5dEbElZ3oD+sT7N8hA8ncC4FfU5tJyF8bpE8h2YvlNwfEABFvoxdgz6+SQDdTCx
2x0nnzSXvHB/9cr3LrZDvL8PGC+lnRrSE8KX12ytGeSH6vIyMtFYxCMnP3aPpyHW
cC4rnmrT1tj1MlKtL3ln6morInvGVTEIlOohgl0EF5gAO5c2vHHtY5wervGPeRfN
Q7sEq4zUTmU2DsTTZUkiOap4gWfXMgFtppCKWBlfZjsUxCBKNaSOxBpdefrACPPO
Dx3bDhdAcqpWjrmfIRJdsk7Mv7CyHUR/NRAy80fuxnnONBH3Pczhn00QG9a3SN3A
zbdbf3nTswD1rTNY65mEZyXaa0gyHKZ6VW6wKAc1G/WUiYN5YX+e5NXIKkC/4sEu
fX6avai/fZrrikYBZ5B0i4epN5W16NH0zu/5M60DRRNCVQKjFiInQZzu7m2vhS3Y
bQnE1/GhAn5xnYqjt0YSeSqx0rJm3h6TuWFk/ydhsAjQX0/O8h5PLJ+UHRoK/x6s
Ae2W7qSUrqaQi0wNMd0ZLLJEQQCy1jxqd4h4pQXzx0V2nRSW9c6cagPkQNkl4HlK
R5scZPmGMXgiOAQCMDBXH/ivuq6UxDeUDwmGgrG3TAbkZ7tUSfCrbjrqRVD3KVMB
N75HcRchThws1YFGapOg2i7lV2tnuNdZJz5r9y91tusM/j6NKaPK1Fu0XiA0YCBC
ToEnq0funRfvkSEOHbY/NzzUcVoXqAXd7ZKnlWQ4K2xIT6wZJ96no40c9hJCm3gE
bJgkJthMVFY2Wi4R4EPh+qKJNJppFHbuUgspdUhey3m6HbMkEDhc9T7WfNF1a8wn
G8iyfNxjWB57utY7XYCsNwqA5X/jrOY0kCCUzjWwdQwvcd/rjJJvSABx2lm/e9vA
Y5vpkq93hGUewOYDFPgSCMgMw22TyWb/ejhw85Kb0r9opPgEDkBIsm768R0SQYfX
62kWG6sS7OEjmUvkrYD3m8Y+HM1MKJnN1Go8CKqZFzrEcmoqJBO189vcw9PCr8fD
4eHAnd2fH0BrxH70w0j4EuqQ3dKV+qZ89fnh8k7+y6KpdTlrKW9pSi7cD0/g5taW
GRvBSA1VPFrcwtwMKOSt7f2kXaSdLN0rirMBUx0Z3yjGg2cO3MgayIDdEnV276LH
wygyDWRF5VEzdKnK7eS8rccGBb2H6tTmwU5kcI41by6gcD0Je0Q5VA/oRItf9F13
25VHdAXJxB0DB7APu6urITdjVFJ/hF+sIlXvdeYfVwktLJonePMwZ4BSWlrJP55A
52sUbTN+8flXzvfF8iDP/o5igCANjWZN95qO4DPjsCEQIrVohJeZMdufzYCEc2Kq
O615f3yc7gEvsAzKP3TNXvBMq9YTIs4Ki9YmV0aPkoUNEy8Ahw10P6ChSarOeEvx
M8iMlr9qbz4ZWlRSrvHqsh+W4O0t3PetvZxkEwVRP/HNyUf+2SBEws5/TNVzRL9F
n02uiNY/NUNszffAF9fekU2F64Rwy5AiXySgvI2mlLUN7DgHJFke2Tw1LuEn0jAd
S2mX/ODEtmybO6ktVYYtd+8troE4jQ2SoalobRN9TY5ax+/ahN64aS4/51At6YUf
qahQW0i25j2vToGcbJC5pJu7ZjhwWOHE+BT+R0yMBJbbVo4pl0YrjP0IGTYPltZh
imDu5kmIfwboNgCssgLAv2rJ2i4pHfb6dcBtRuwm033/Epe0c0wuFBA682+Vh4mo
0JvF1e6CnY+5p5l5vyNM6aHePrkC6kjlrvcmJgH73HbXHks2SWFTMyJNB54E2JSS
+4KClHcU1bc6hzx19dW4QUccq8VFe4RYn/hJP1EizQ4KJdi0IBnXpKBCJWkH3Rww
aonpS07WZeQlcOGTMPqlqIXjdORdQEa307JvRu0HlUMaIB6hdznA+r+aRc2RyxUX
9SeWzdrAQoxwysc2MzVpj3DatXn3OE/A2Zzw9t4ua/LfrHaioBmjIdlJlfCkaJri
ktK6H24EtVNEd5ld1TwSfYDRAScG+h2UXE172bLY4J66Mtj4Xw2tXgWeTJ6gjlUC
clP9kYG1Hl/J6EYNLJl7f3dFtSc+WmB9gALZ4AbbPF6+h9C0UQEEywWWlu2Sb14k
aBhQaC53NFWZCSnnYkkhx7UGlBVvMUPImTc5oAXkiyJF61VXmPX2Hw4P4wR9TlE7
BQERIIMWp3HnA39WenHGQGQAUju3Pzn23LMt+wGMlNr6TmZs6jm0Dt7+cuIvpKYA
13xxn3sBy4tRGoTy53G1oXmlBREBUoaImRaQ0FZwUb9H8HviLLOmZimDmowSO0Rg
rwbO0sklai43ocmLD2WpwvNvc0ymPnPvLo3n9kR5LF0KTe1fA/q7jqpXpRBxx+PV
4kiaUT/e6xavZNeY49tTDXWuADe7hbdYC5UNwwm/alafy+Biuhgw5ou4Dg2ynGuS
a5C68qk2gie4rREju3A0WDLZm8SJjy5s2CdDD8PFcaqPoozB2sSVzUOHV0TaI6rb
D+OfgPNnO6hXUsk7dMt5k2p/y7GNDgLKndRENH/juELWZ668ausSybIbElqRoXuB
dSa0yJu81FBTr14M0DrmAV5yUa97XZu8BrFGYy3zD+SUB9J7Nlx4SQIUpdrKPDsu
CsoJH+iYXmnuQZH22qqzeA==
`protect END_PROTECTED
