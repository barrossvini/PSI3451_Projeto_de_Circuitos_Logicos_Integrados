`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
36koiLISnq7+pz+gOPY+qvsBIgMMuDlP12zA+a1zaHgfmQzayLH0Seu4GmsGkZUM
pYeZTBCcT/T7tfDZNNFHu+E0OKWanQeRXYZmpqRby+IEIi74raQQLZrnC1anlc49
smd//slqn5Ts5ff8GA1ifUWg8TuSHvz+ihdzLUQx2ai9i6fl688Q+cHKVc5gkr+m
GTbdKU4nkvzbbmChTYstBdtRXW0mq5LT9Tp/6lmkcreUUk60Qg5JDTTbW2yKK/bz
syYb9AqwpfoXMOujPMavqfiFz5bLPm82Hfc9gtXCHS5982fcGSwSYnGBI/gDxr3A
vSZd5R/jhK8APSHApMiRgyH89U10gEUd+J6Ck8ifkofigQYfzSfVveTpa2jzAdTK
Kt0NXicCd063CxXl1zhcg6A8JvZwJNCwHUOJa99KTRmLIQR9YoYCVYgGkhckwCFG
O3FUXgaDFI0r6DkXJVWEoSpyuPCr3S4nfIL32JvbqcyEofMnSM+M/g7hF4A3+BRB
d5e2E3jxb3eCrK1z/k1VWdByVGMbAitRfigv/yOFFiqVhpjbpTvPjSnSaCzd3oT4
7sHKIU5cqJa+GASQgNYxQUiS4amoBq1r6Hx51dUVRFKxxJaMsM3JbnjJHO8B2ZHC
wEMw41VRh1IAnOq1hjSSGW16Gpoj6IvqBmDYBiRde3dyk8gqtKLQ3LFhEEurxtzq
`protect END_PROTECTED
