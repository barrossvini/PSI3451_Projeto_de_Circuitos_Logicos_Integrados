`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ls8khX/iV+1KMQ1h/P7ZM2W0hosu9tcSsj82F5LVTStlJlrpfP0RBlGjouAfF6kD
M+++qceC9S2n5inAfrbiW0GGTXVEOSfdEkWZvDTPC9QFeTiOaS5kXpC23vqTjra7
ssqkIRfM3ZmiE8tgbGajWD2xQ1WlZmXC40Hj26DmLhdptKH4D84fTex/Tna+ws+m
yBOdcDbFvYdGTFgRliSlQCvTDiVk9Dtjxa1qo1D+IhUQ1x1r8yO7suCn8rrJZgq9
ASnu2knFH69IzB3078EGjGXhM/KsIuAtiWcKMtxjq9K/rmlEk/Yxu/OTg71XVuBr
bvYRBity+g4vq+fH/C3pP8WzB6FxCDwimJXzepV6ul/BGBCqd1LZ51wuf3S2SBt5
MU9I04SNJuVVdbGmS+76prdai2mDMVnmrcPtGqWmTdpw/PYdrquxF1RKEBe6l90X
5/Qfmv8R3SPqZX2cZ0EKjHGBiSDgg7YfHS1JsCIb25dtNrBGbcgUibYEYs7M6jTS
cqtaKqTZxyPVNXC38dIlU8zqkGtx38i2g+xA3wRewyzuXhwc8oicOAUot6CjueG5
TRFCWLMOG+GJruP6aMi2YF8Grs+SjmuKO9cKpxEQMHa6E7KBuXlyEQA2mktlVii2
8vG/S0LXhnhYfvmPCb8tulYZR9uWdkyWc4/HFckbV9psI8QScF5XYfG2YMSuXF22
VkMCMu9n7pliIR9HPLBAQg/S50UXdfAZakQU+iRMfz6JTHxtY/yfe77A+uOHOZB0
SFCs36Pq+CiwCS6a0T8UbPcoIeNaGekHArntCFOuJsUsa8q4h3vQ8bHUFVHEGhtr
93WdCDaETCASn2JImlVLmn07dqMurYxDcBi8LRB0PJ8JPdFrOm4edv6E+a0G7E8l
5okdhot77myKbjRojo+m8Cp41WZV2Eigr384sRyAJBSVMyjsivSqqEYFEE07Lk5H
qbO7iv/HCsxv+KWwsLmIBetvDXoinLmmLR5SUBfPEj0ezue0fUUu9NZesDVJ2VUG
CoUIW7ZNciOa5L3MAG+YWq+yC6JD2OeGlMm4cFXG6sdw8qREH7Y2shCia/eo1vLg
nmA2se2b3BoMsGtUIcNQNu7ohwsVJQIrZyhT2T7tGkvv56Y4IrirfMU2D/3q1PqO
kN7Opsx9brrliD619evGN22vyNOsHnfMghLAUoTnm0Z/MKRvoYuCP8HxRu7z6w9o
xoGzK/lJMSIWFjYrv3jb80OP8yjhc11IISAqETWuc793jNY90ii6KxrqoSQ+myPS
xIPcGIRCLciT4Rjk/ct5iz+azh07dSw3Dr9JvrBRlq4SLpCPeucDVh/EM+WH7RXE
fmwhS0L4cPuiOkoxKl7Ch3Awj8UyZ/oprg+xUuD+dM5jaUJXwLCtoKcnkQRree2m
jwssWSYsWY8YnyB9SmQ/nLs5Bqw30ahyavohpM6WT2hOPewsZa4XypHF616etB3d
RBF/52q3Ui2sjG76yr1orZlgvHHKuAfxAFYB9uxO59jX4VA5wNgcNRFA3B0RsQFN
evhhklbsy519J3h8srlPBqSQk1Lnlq7mG6Xidsy9rCRE3DVeQCjcUIg9zPV1mtty
YwanTwFgcYmDn2rXh8/rHAO/Bi4NJWeMPf40drKD5cwXfSWpxS46T8fZ10Y61QFf
z/VEbuJQ5T3d0uwXXAxSFH7asxb53LhXNMmASTPpWVkloqx9mC37fcudF13hj0Yu
tcD7R+c7u3Zu+iSA8XFxBO+zKRTL9eZq09cW14hxwFNFZLkhc5C4PiiH0LljktQa
MgAxJrAfRkJAeg6W8Dmx1OZQCZGh5wwUrxSOLiUOyF2aMmnPmPYQoKxsFWQjb8pR
l+lTb/xFN6ePOKe+fS/EYQBAaFlkklw06Kt6hK/0Dnfokq1S4GhOWen+K0pJlJQX
MpKYa32gy6+ViProJuzmErwngu+0dhuUiKRMkIcbe1EJ2jv7NtieCpeTGSL+0twV
uaxYoljUuC22ue9W7uQbQ1CUuIh9dhhsCqSWL2scwPSiN99FJRCfrzHXEwKMLbma
WOHKzY0XAijeQBTcIlMqSF3eF1FK6WDKKl55qVyp0gnoODWKO/YuJHA7Ktyj3fk6
ptxTNilq7njdgiMbhY2snxaifUtKn0rHCV23sS1I0jQwBoBBX2axoYuXiP+/lCSL
a4qZrfM2ly1gjGw/P9nW1sbsF0LMJ+jZWLBo6vqIsv9bmT302g0uIpxDegt7JSJ0
KmP5aIEDbXNPsSohHLDV3PrZvs1FRNl+tQbGQAx4zLYXlJkOy/15KVUp9IVHYs8O
JwkLMiElNsv/aGS/6l34ww==
`protect END_PROTECTED
