`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2doyjXsWirffRjuJoB0lSeaPfn5izNeoWCD5iEgGd7vYJjafQ1v1BGzMW8bm3Ek
G7eIK5PQ+OLRihosFPew2XpduJWCeztErMfqoMiG2Rt7Hic9X4EyLfbl7UO3kb1d
5kxHoUxh7CHtsFs8lfwbdLJj0OWxd5ANlqIETIBuvCsp55DLu7QurfIFa20o7bAl
6r9u532qmZJnoxyeYQuuY5AxhBsyzcwYGr8exX3Kl30Sftma1LlLOF0MH8Qbg9QN
TQ4VXZFGa/mxxpmSKnCFAhmT+plknYc875+7KuibwrIP/+ris7uZx0c/FL07bG5z
jcTLueTty7Sx9ogmM2/9bPd1qaDqIykf7NPZdtNxNXZJmbfwSMS7NVYLVlWxBo0W
BcoaFhsZiEP1pXg2ztXuZc7QNsTIJf+J0s45l7fxd4QeMwh33VP7Csdmven1wqyE
SQGLMG7dhnZP3Poad06UXAAxFMSIoTiPBId6Z5qkpEgCwfKV0moYSurJYprhlFb9
NDKusfFxpfjgWvef4rMgbP8j3fIiycTWhLaiO440XMFpiLI3dscpkVJ9XBz0LV0Z
7PbFUGC/34yr1qdDzadX5U3DpLvYNcNGo2ASCVzpIdMsSMm2c43yafft/MtxbBcR
Bh658colmp0ycKpI28vcB91ZPzfesRHF+EBg5EGkfXFQuvE2Ms3+5r0oDor19HTw
T+9Y4ksYzOkaUYKBYwab2Ir7XRkkLHrXmjcdRqxm5pn5jpfkTXQfWBx4ywbWJoPF
u0N4Dh1MlkRfpiNMyhIaz7vUaK7jIFpjaWm9TjSgD2zJdBDbvHlSpIqiFjiodsWT
NlTK19yhvgiV/ewkJKhxvNBspvAptWH3v0tyGaK9AVfTtLwKAg8vl5HotiFiPhih
q/nIhvMPmqMKMxYKwP+69kgqdMYL8LWUacX/l/gQCiHnmxfUogDGCaaMxQzfQjbf
98eTcax/UBc8ZWjpQ4Muvw2qJf2qNNpcmp4ZdXr6jH84ZfKDnjoLivIOM1oq4II/
fs5gggTH3bs4KDZgahXmH8ohcqZWl7wOeorsxCmVYtFVwG6x8yHLkFCLCSr//AcR
yQPQJv8DLuNv5rMEDTvW6uC91Lt1Q6ILh+EB7SOnB3PC4Rm2z1RzsNvDw4ZM43k2
1tLriHejOrILFxsUUi//kKARbBj47wcM1//dEOWelMPjgLBHxGjnxtxn7iixzX3R
IyMERfouobOme0Pii+fFIBRTXkEbqscJGZF2oQo37fkRpdn2pIM82mj9oL0zmhqv
85kghg0TPHGt1d+AOUDxZWv8/GuhYrLrtmKC/13VOlDqnPGL43se3nsDz4ztlLjW
zG4lidfGKvYoDOWOghzUQxkL5ENFLIsXYrPlf4FkL47OuwsD91Oi1pfhtCz4YudY
rEMX6XZZVseQcOMJwA0Y4HZGusO0eZIy8C/lU0umlspwG5AwquhoeEKPaMlXrKyX
qYURHR5FVdBhgKhgtekvIdXStEL7y3uWjIpivNhNhYmf06H2B7pqZBYfrqot44NU
3cMXgXCYMrg8Ltk4fb4BoDGuGmINr/bbX/t3rt3+vgndK5uBa4OSPrI24oMDHq+7
m4fD/j+Q9ier1V1FnBzImdItQAWY+LSo6z5URj/0X9KyZM5i5oP4mKLBxthBkHKP
tstMX2HK8nM/gnZHntcSM3nwyfvQpa7D5Tjyk1oKjHgj4zLJmQmPbAfeKyVulPvU
GVPTnuZ82WkkRI58yV22E6JCQ093vaLcFALkfYAyANrrSJkUn8Gq61XpWPEfKql8
WWtacNZkwknaHan0Ajs4FxeaRAn45S4CkZF1/XMi/7Mj3CNcGg6DgM76+EpIfKQW
p/c7Jr8i2XHse7yVfA230wubmHgCJYkEkllyhBWfqC3vnUMgTzreVyOyzCtkXk5V
/163XmPcJgip1GpDj3w2jBJ/ZyxEn3031L7SPYhqMFFN0tB2vGwKJyirtgCkXTYr
oOQMnMF85VRD7IO0Gwf8Jpp+55645u5DAMTDP/ro7kvLMMYJpYXbsd2De4EO+hR4
WtbnEyB48nIhEShpDmqzw8sicgcmNEz6rqYbjKwthjah13eBBKWO7w4Go6S4Z368
tumJoCeToK1QbnFDaLw+o9L1XU9sIAfWNQTCC2T0CCI5SIFOIMvItqdDNU/BpD5n
5akK9oLsjFX5CyWZfWm8sVXDt1XavHAku0Tk+zLJowXiIhKiT/K58kdx7UwButrI
QCj+XelcPiavTMimc5yvWfWrSGMU45MUs3y2+bF7kYCYGctCmhhNq92Lgxr03Ek7
hTHnh3vauXGTeL3lPth7JTr2QXZIMGZTlbIfYwougBbuM2gsT5Iia8ofOWQNkSgV
uCEtxdPuMvCE0bJdgGd2mY/YBpp9f1euylFoqXbfiNoCALkuDUykOAGKwaZomtI3
xWaiqbX0Hueqpoeo8vv8V6JdqOQQUK0VpQEcjAIMK54YuodvxhpgBWBWKltWEGhR
H5xxu1JosBIVZkKxJgCjD5FwgtnZwjBTjCaYby0L24OZHsz2S8/Eg39p72eT4WRU
sPddlViPsGeUjRPq6+Ixi+NI3d44TwKjirkrhRXynSVf2Ok3j5nMFeAspX1NAGU7
AeW8BGhGJnf5Bb0R92YPlvBChsvWsgcpffGtp94RZjrSPpcAXwoqqlHuAZvJY5po
gmdTpHUwC9UUJYR4xhA/QdptncYPzFHRmMvpko2I/WyiOJku71qYeA/fexasZZ/Y
IEsZnowj9Xe6unFgZ/ppS9p9Wcbz466OBocchpGVSQ7AE+7LqHOM5EQgAlg3Rl1x
fLXs69uYAmZqhUXFyZU7HUNbYbIwHOPhsItL1K7b9EMTrBWhmeaKcsAKXHUqK0ks
kAz+bD6QzcJvK9ZRu/vjEDfnpmopYAsmMmRcSMdsmVOOFEXgIy4umyL3tgGipzc+
E9NlA8xgne61I2gf0iezJDzj6t+KtMj3iEgp+PSQjGTyaU8M/MAlaaGWJVxno2p9
84oEGA6M0OcFdpeLiO1vbGNKcOpnnNxRG8JjkrQP7jF+QOLcBj2yTl1TO8LEf0ef
x1/AmDy/mL9aLNqOO/1O4NH6SvC+KS2uU7z3kLMa4nAbZjpOZaE87b0aniEeCZrI
bB+YTXMgb3pQaSa3hIAHAtBcbAeMH6AP1eGZ7dyS1Dg59oBD4A8b3zmECVnzxT02
vO2kWewpgc+gcyG2J5ncK+OSpH0Ou7TT3ykgBXvsRVVp21aAcUDkEH75R1M0Z0vW
W4NKygaExkeozIrF8F8PeVCdOu4lbGZZQmjY+nEHnUmhEkPD8zxioCMJEj7TLnPB
UJiLFcKQitDWPul45MT7WV9GDP02LZs1XIPOookm2z5P8n+pW4LHyQ5pjnkd+YFr
OKwMhbohZmpktJGdvxdnR9AWAoJZwMyjmB41lWcvZLlkDZvyvy4HaN0IPCMgrUVB
cWSaeo1GCl7Fnjx4rEvHHQ7GpLd85li0KouX1Tr+LsQizdS918dzeFRDyIY0hLof
PIOzp5nXeJbXmG+XXNFD8XQUoUi3Xr3bEFuDdRHfP7DgyE3YCfTGC5aCc/44wqmx
RoqQXPL9289yO+5O8vrVA/1XACPmxiGxyBQuqn4hooFEuSmbGuIBPAbVOWraYkDM
tZrML4vcLXB5AnfNslC2phBpfAnjau6CKv5TtMTYxhtrPlPoDbLMoRTS1nw0IBfI
OEKj6GivF6WMcTWvG+jCB/80TQ8lbGLw5rF+RAxIqhO82Gq703yXMQHQ71tmDLus
fd/RdjnAl7a8E6hXoOSj1Y61k25QrrlqFe4mXnlUiuKj8Jb39MWDJFKKMFQzvbty
cChtEky6LiQPocgqyiOTng1azpuMn65Y8uLprNnDPkVDhyOnicwg6BryKzz3u6n5
WhuoCJTFY+T71DyuYOqZZzloIgXmkaCABFVq6L1sgweGNOfta3O0QNi++9EbcgSL
r4AWA1cIRgTIx/kDkbNMWkfRdc6t4oDu7LAcddlFT0fi+Hdu9uPHM85qKyM2Tn2m
3S6UWHaVUxZtHGPoV6r6NhqexO0Z5BHjN+BTXQsMqNT67qhkmtlWSDRIZpXTaXda
66e7G58TG8pX5tGlUWVbzVFMZ5t+b0C0tClI1ST58vA/IySepKJrcPAVL4bFwG69
sVLky5i0C7V0kkm2DNZ1D5JnHwqkKuKhUzBUGd1imgRTAuWk5NONGtjgpG/MzhjQ
mbOskfEERqouhInZtIQ+JSVmQqv2fBDVRAI5OSYWjLYhJiXuAWF22Zs2A8aZ/FX7
VUFrqSHVTXuim3xtwNv6Kmt3w3RTW8W2dF3/OsU8sKk9j37fcD/16mBPJ3Xy78Zx
64yxaI7PYsX9+ij6wIbwRYcN4W+HNzO4hmYG6y8GgXWD9LMyTQiUdNktSXVr7GIS
60hk4vjJ22vBCANR5ZwaD+YAlqMYwwSeY/CI1SfHcd1O+Gy1GiTCM+xF0+PXpI/4
v54iyULWR2Qn8mUdvzoym/XTUWamIvUN/q/ulBTjuGMhQhbQjRJJMJcHcnVknI5V
WgLvoZsZLkXuN8WOt+g1kQ==
`protect END_PROTECTED
