`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fdOeQpQL47zFXf5rrdibhmUnv26OpiE94pF5LDAU9rA9cE36RhmnmtjuZTRA1ame
I/NsZxe0JW1cLk6qXVTCjGGY3OTYRNXs0Mg/5kad3NyXG8EN3UDbQC15GgdUlz7H
0N/DaUwEDjSssgg2tbjwTD5ZiB1MyuD4LB69AdqDKLSqO5B8MjdBQRuXsJibwT/H
PjdPA6NaXvb0rbg0uDuZLpVvz9Bo/2yhnnG/Fyj60IUiP4U3dyx/cdIeCJ3+rc6u
VsYU/7AY3Gw5C7heXCY6YoeD8sFmjijDe1M3rftkzL39Ozbsu0cyg4YXQJCz1HaY
oDfWRFuA5qXgeJk3KJdMzRF7+I1WGvBxgfDBzzTa7gg7rZgTtVNiGQd4qMu8wKEs
jicwPeWJhVl6cEysjlUA2l56OR4hTaD0/OyyHciNeqYCR6IOcwk1j6j3+sqsEtQR
q50F0jTc+LuQ5LHA4kIYSSO5T1FeMfz7O4YNJXhOboBOL1yyVasrZWrrWHrO52ne
071rQdA9A/b0epZ66U3q4dy7d4pf6ErQ+KnHHagpqTW6Mj3lWRXHmGql8RpO6pID
TK2XKYtDo9IwCnkTZK6Doq6umMRFvNkILv/WXD46JGMuKfVG79r7EE/M2Kd6uHCQ
cjFgwXb+o7h5wfCKDV22G41635OnnqPtZ6CzaMaJqS+TA81YK3iJTrqJQ5eGclXG
bSlXrSVAyiYsT3p/LIIDIWEK8VUoEe5IZJafmygte4/0ZdwUk47AIAWhHvupc7j5
LEzw2IZsTJSY9Rs2nI1GNuhpC/csrNEeHS5wsaYEEjsX7DwNRn0a0+W/5eAWsFkr
TcZAM7FVrGh6T0G+HpVekQTc/w6cbdgnzpN0Im3GLc7LTcOfAW+iXvPlncfLusIG
Kjy1bp2eOgFiKcBelK/Qg1br5kOyK54d93QY5GQWCVU+ORz41qSqbk2BEnVn/q+g
h13WfRtes4o1LzDuu6eBdYoAWjI4EJB21vtGuOfyCGVrpLXKK4IuV2U4eXkE0uog
LTBproQMtrMoCUecSHaDnObK8kn0mLGVg6wJCq++9YSWrBOQbULNBfx9GysquOvl
cj7D4/PutQovaXk/lhKqKYgUpYE04A0tx6PcCE4wQoy3l5nBkrDvy3F4y4vwiLvV
+R1ZzJB0h7r3CTYnONHjWpk3eUvD4g7RHLEk4gQxMMwwhu9MuqqzBRBRQU2Snusq
5F+NGScaFtzpp7+CbWzMW7NyhW8hbYxoUYlS4uorXn4P5wrJx1PXwMCIVDrpq0e7
y2hQF9ZLscdXvj8dUVXwRSR87SsbGRvR4JOJirMqaKkGA9FeepQ7Y6AigDR0zKax
0GFSDH2RpKgZSJjHDqgFJAtjryF72w15aXbLSbyyDrwj4oE6AYVIdxLTfs/mcv87
yjDctAVM9CRScNoVti4OGjNWJuw7W3ld+P1Nwn/9arVRNqPcYH/iAvIgr8aA0PMx
MYuPnTSDp5w358iYQpGdJ8xcxCVKV23CJb5KuRIeOSo=
`protect END_PROTECTED
