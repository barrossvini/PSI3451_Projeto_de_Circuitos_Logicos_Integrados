`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bvqGZ8+uSsM9E6dja+ZWNIYRXIwZXq73Wy04mRTuekQdSJn8EReigQc6cL2NGqpk
cFDmKenb2cT0JAlw7PHs8gGAbh3NxV1eYy9KxZ06voNgBrYf8tA+j8bCf7t08OT4
ta060RpXfAFH+I44fV5cWR/zZ+jzl3LCCMo80pp0ixmzDNOqbPfYUpX9sEYgXUXK
ROiP9gUtlGLEJ70vwwhnRlGqDaor0SlpSWuJe8hR3biCN8qlmLlvvIiUyDcmIjmX
4ukcw4OHOEpxIEk1PLpP8mduhqRuW070L3ibhcLbyMvd1odTofne/yVpcDoTIAqq
K2I9KlPOr0gPSQyRjKSR0p496IBwfOk0Af9gYUS4wBDO9HmDOcC0lu+sIJ8EBmJb
NOrtdVg+GbUwi4VNraKt8YUctLnpdjZrW4+TWJMNLZ+gFPGOQMwpvvXyzuP5Ls1W
nxclBmUgkLW1KwQZgzBQEFE0ygorH2LKJOGLi+G31unkibM2ciythcTzK++H3waL
x2zlxk6kny0GtyI7t0Mbx8+iRwqT64PFXKr6J9ooeJvEFhq3wOf8Q5Y27acUVWpC
u18NqnCzH//RFsnzJ/SiObrd1foeiDgFAvcQy+cwZ8lueKfZbPvqrgH6nu2hJ1b/
Bw80hadPlzZrBLW/bf5YBhImyoO7MO+ePVn4x16/7GTCupY1vIMoxN16ePOZGFT1
dBHN4MPQwin4J2f+6Jn9iGGYMXJp/WBZoWX0dMGVAAvYQmYt0L7yRIEitP0WfhIf
gYbPvWsGfBi99eL3JFPfLVisEwFwKCdABD6UtkpoTnR6qQfTqF5nfs2K/CRXD8ii
t5N0GExTo619hIs7hfM2lk6NjdrjIFPuuvPRZofBWYJkVOA8kARUKhvKA1eEOfQ6
oWL2r5LikHzpqRoXZNH4Bv/vCGh3aIc2VoOONlKm4rztq9bzbue29FEMFj3lw2Zg
U4jLMNcWbilFkIX/dcOThFRgJnaDI665P866vqJbpE4kYDx/1kTr+vnRh7gPSubA
L9rVJIWh4pTpn8YnQpAfcmGVLs9ssSl4ZpB16JyDeFg0Ce0Q69iDNnm0fyqEgp4F
aqGExgZMH56eIYn7Deetd36ReC+o4A3HBt8Hr35LRDYE2lyY3Luas/OaDxtBeCGC
7SuberPWII7PNs1ZfZ2/huTqPkh6Ekg+Bm6e7OiOsaxOhOyqBMap8zwXfwiFv3FX
6EVsVnGu+TFTXfj7J6tJJ0V+CHwz/p6kZ1Y5KmuvU/yySwu43eWwFF1zzN6Kw6Af
UghwRBKIV4/BDM0anAEyboTsYDqHMTtDwXzQ0zZKJDGabzaQInwCs3pN+wUbPW8B
ZsIu8oyXjiQ9Mgx50NQeafPKIj0LhdhmB9Cw/KB3HlgfSboqQ7YvUcMa1jBqeWte
LhkBNDa6EvmpHiPBrSF2nvACRhzEwBkJADsdHfbl/4MzLsnLlBdQ0kGFqunseY31
`protect END_PROTECTED
