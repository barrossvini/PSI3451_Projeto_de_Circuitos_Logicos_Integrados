`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PvpVPSX9COg91mYb+w+T27i2Fp70vDj6S92lG+GTLuBJ/nm8AJyr17rP/qnQtjPm
uAEla1raIoXRiX24FtzvRnA04mqS8MtfdEjRxDujlRxHX3YB+4ZvZPcuC7QwQrJJ
Wm8vW0ticBEpo1rkoGTbBs8x60YqwIP7ycnas6mN8/YqeMBYfzESFReIfUDJE1ty
EZQP5wRDZ3f/RysOZIjY69guJNNOi8r/FHGULU3+25mztXAgeWDTfUzg2fTtcVdw
Zs75pVkmRLOxJMK9GeIDIRIU9KrYSvQyHM3g817Enj48Ikh3SqMwHETuSFWkLR7h
NH/IH8YlRyndZQ03A7ntOTtPXgZ6JQ1VtZy6uAN3Ylog9oLHb2Ml6++kkeSQCUCw
8bHxHAxwag10U6Vy69V79DqkZT4RIadw3cRZygWB4sGx+ZpVBsIWa7GUhNDgLyEE
SzZ2CGi2rQtqAeEx7y0c3bxfJ5PP4eVTcIh94uzBmJNEoyMFbP/okNhHrJSELkTG
FAwqILX/Q+pB+O5Z2H4vtjbAc2tjpJP2XwcWF0VMWczVXXov52sjL3RyHW7SFq4I
aMl8gD0GhAlEBrvnI5qW1iWRg7Hcl32lqTkHV+QqKcoS9qMGp6CYDizCSE67EAHR
UdQmv/R0NJtB8H694LrqGEvb1HS11tNYQxAEZYuCtb/Q7g0Rnwb4HH53Ugltee7v
y8PTHwUmKmugbXxeP+8BIgKv53vopS2xjp23/9IZGQLsrlhfAa8v4+uTdZYSfivk
3VPHQLuJAnyCEdaVfFCLGkY88gIZ1cugsF0ACYv/nIbbpyQ5Ji4PfLLSANquT/0N
abvIwxwHV/eyeyfZdvgGsgvO1VoATJxiKOuBmgkIDGnr2Mq2HTzjt678MHCocUmc
aRGdHylLvTWZZByV3mRBrxBuxcoE3on5S3ZXbWKY3kCPJ0gxWAniWtIkk6O+KaSz
J09t0Moopw11x4JJ5WLjMMzdDHUzpcVDEO/UfVro7hn8l5W6Lz+00KJM9+ZSd3nE
pUO9FR44dY+XbRRgRqTqTrWuMN3HnpxVocRtas13oe2rA1Hw5DOF0KKRr9evKiGy
1KUWFgukIhSW/Y7RoSxKZ5X7mi9w95XWaHL9BtCq24jWys3ZuCseGRFBMyCXYnUR
VSthg2cJfrP+bfVohMq1L8RKLvkfFGSsjGacIknW4QcoT2WrVwK07AlLz+yUgizX
QKGg6iO9DCcEl+ZdHIsuY9gQj2dHy9gH+k1grvlCc7YtjVWjG82NZBlFCa+VlwgI
s7fSQ64nZW2qR56LxVhQ1KxMHG0yfjO0kLGaMpLR9RJxoLb8PsE0SObkeG/iQaRJ
DgPJgRyLkC9rcplUPFzhmm97Jh3T2Ihxe+tCD386wII0dCH24xWeJgA7407Md574
OKdXIBNQGBrqJH/gwS+6qbl2gatqgqDNLs6BIObZbHJt/0V1bz6IsSxcXIaTEfoG
xzuhQeyqUOnCjuc8kIMk+Oz/wG7Knbzc+HpUoOZhh4KP8EbLoQaQUdehqlloIQ53
Rje2pOUJl3QNePDskjLfNoJzP5YJEgwFBV7HfcLe910YnSZkHXbAhpVD33K94dAZ
+lK7w/MWgv2oeo4IUs0uc+LdxasqIR+LEcrWBFr40jsVgw3JMYsdO8eaSMAfVNzp
vdw7tbSexUL/TG2znKILuJd1ZwltgBDmsQENwiwMeH54ltTHSgYw+MT0jOZf3glk
y7QC6n1fWk363mz7y706mHw1cxsV1z+X0m11RK3hzaXcHJ1iX4Ds0uMjO5Q3jsdO
MOVLnUtyIPePGUN+WkfRXzpYWbShjekWf5SCdwzbX9aySL6SxETFz0hmaXzuZG3K
0Ab8XtJmyg7L+gBlKGesPaHtU6Rh5IZJyRtOxTu8iqkSATulXem1L/C//u7vlAit
wLIzEDmjHugzLR6ldxjJ/Qn10NoDEMYn6veqil6NtLvRunF96GpsR4lyf6UtuOhK
rUx9lwdseho0vnD5EDJt4sX7KYVUj07Kx6u06aGNnK1w0d2LK/1EiO1c0YcGH7Z3
dJPSvQ8ehFp6Rf0TfizeHwYVf3qRM7KKPhsHb5lPAD1ms+tffiQOnQ2JUjJJtVDw
JOGX57iPmmA33VXzURS+trQjJFt1pH2ODZhmrvI5lCzHM7cUd6+5HEp6gRBCzmWn
eQx6LnK1o9xU6uR4JXoOfScwGTz6S9Pg37hX0b4gbmO641bt4pfomDqpppAspBjn
/ubGd0b4KJiMuNWNTVYQDN/HPXlZIq/qUyRskVXIcbqbIc8fhAV8ZM/op7+yRNP2
mfQZge5O3GheoQxDBmvmPL/nH4celOYPce4NU/KbIw0GUasTsn4771AROjw4s+Gv
WNyWR4QIGCLGLZkW0CjfgFxmlIxfkHioYKYrrcdJKZSVz9UwLvjslFh3iOvmCxyM
qcbc4UEqhStVULopuFSXG2ve2pujRATsQ4QMJCJe0c0F2JL+E8yfQNhTHORVfwQu
2tTEV8XRZXF7Cp1eDRId+tLSM0cULE1P3l3wTuI0GAxAZpJnI6H7ZbVfOoFfDdTf
b1H48SVEYN4B2aQHAWsFn8lUH50K2cCn75gzb0pjSXnrMKmt4I5+oyMrrXYc6R+e
uuN9iwAGfIU4rnMz4GkfWG0Ohw5DFvk+1w3KZAfGrvoe0jrGHpXuIvE4ilPJSpco
1//otS4Q3UZpB+cbsHzI3hfjWpO80Z9yJRa/tczaEk9q2vU+Rh9bkGDFWJW93taL
F0o41DYZC0bQ5JeFmzGzAN8vuPunVlrcCWQLhydcBHIDUaN/Uposqq4CVOjlvdej
9xwCFW3eNeSqjGL8psuZXPFLmzypN2fNJquCJ/rUl7LmVLEELNscW4NQXnKwS8gc
vd1CnczzkVf85QS5F45j+YSn1KOuSTsGxU95d0VgTAyWbBimru7ZWTVbbsCkhczl
oqGleIiYSfY7hrgih0ajvd0IIE0a1VMHhzUfS4jljd0f3ec20p6tpXoXRKNve2AA
hT4scLZB3uy9G2ywiwb8eRlK8DE+zTuj6fxR0Kb+KyYMZk6ekuFjZ8TyICHFAt8+
hPLqIbau/Hpazg1Wf1ujuC7Lj04lPYXfku5WfJ5ITEvZtyB992gEVNdUFTH25Oi/
U7E+/55utv+ZHkOVUTfyf0WAetBh4HJarS4rp6EA0kNtoLxzsIEd4u/Jd4PEclvo
pKwq05/YiUabfPDlvtoQXUL3O2jAtK/+Bfv4R0lMWtUppbKKp5+5u+pHr+T/GIup
jK3l7al7l3yXx3j0YQjArlNigUN7BiqM0jNAdKE7eysc2vFS3aDyN3h2POaBV9Kv
HrJK9+5C4qIJq3CJjuvJEKkyM+359ID8pGf4jyYGZ2rjgN27TNvRQiHysFaQIt9c
1tJdo7nRAXxA6QjCMdci+TgmrtM8kW63mYkXTzo5yqwgiT9gySPo7meHQgRrcszB
9FDfUfthQDJv/rmVSBGa5uaWP+NG7w9ZcGATR98Xr3dhvBfp8uMLzboblenhdTlJ
620r8ntkmI2xzfiVJt5M9TrV9uDJvzueqGxeP0XHsDjjAAMYNioLwK/LaWRTlgAJ
2F3NUnDGpoX4+q+1OGP0CJBDYOQmO9nhkuGbY00l/QGVb8h0KuKRHoR1A4jF8bkm
kUYZEw7O06wBDEHJDOEtaEid0csH6r5WTg5BfVon8Sl6f0ljkG7PtxqxFwgm7DTi
3zsOkLuoCW36FvEi7ZTRr5a8i1Bjs1e6xUY1Xr7ljzRrIafvWOue/4FXSBkbN2+5
AFwdBzHPo7flNUkYIZsBmLM7S3W/4LNqDz6W02xs+4IV9Ey6eW2t+dWwxGTbusfw
64IM/CHt/dXLOU4fai/W1JbcGD9Yjqohjcq2A+/XRmZLt72x+f4KT4f/26+cChEe
KE9TmhwAKdFDihB35bTCDImIl0rVXYIgLChrXOw2qq8+7xXssJ0oqzJvtQBqWs1S
7BQQ/NbXT343CimvVFaWfHZsT5lzYooXV7eI02NsDdpNLJWXQ6TaQqqrvHvmFFoQ
Tszo/xhRCUs4hYo7YzZhY857fHpQOrctdCP/t81qx2r67UFIt+gB7XBme3bFOqSn
EcIszq/lGNSqzJ4Z2s2cCNpTLCI+R3X+YIwIXJsMQRc9Q5RVFkclpmGhxhtga7+P
d91YDtampgaCWyTRcVyjnqR5I79nbpOcM2qmlXl/xt+zjreUv42Hk+ZVTXLg9AY4
gKt52PDmnbnFi/QXYWeD6p1E+7dekRmVUot4TP1eaXMiw2pGeRqcn8CbjXQGpuCe
neW2MlHLPW98q83QiZF0nEsC+NhPdY0FOIcQRDG3+pZfaxVGfkwZhT5jyRnN3f11
q06/dQMd3dIyNW8rSyA3VG+ugg8n9elVbTOSXglriGIweSDj4HH3gFLbx8hVeDnd
5kuZ5XwKEj3WAmPgIwHpr7BgjY8iLoSym/V1oFQl5qAHLaeQ+Aut0Mf/7kkaMBGO
mGYc1T1VUBjm/v0S9+qF6KG1GEBf95bC12UcheIGGYuKy5EUI2N1xRRXs+lfNJwY
deQZlXTatczb5b8yd7KRIqmfPzySoRoeE8xtE9+z5gELOdYkCV+3r5vMKqWhcz1/
4wKm1IEH6bOEVsoaWBbL8QgKvMfTThlfLV+KT7fNdZKxJEF5jLMJ2tA0yLjLGDZG
uVj6dUbfHlea3SYuIufPSC/kqvxseMXfHTU+z6WpUnRZo4x1UzSfKnJC8Zv7Vs7k
WIGUnjCKzSOT/bk4A5z71785dHzloI+WSl2HJyYoi5DH1Yq1Rf7kuIKj4sJfRJQ9
bc6sPA8QOk7qVfDLrT2W5Jfz1eFNffoDfI3OrDWMYRonwxpZiDKIJmeC+0/zA8fT
iChI3/VkIuw0jqo35u9ERkOAz2SYsTayZXNuu06c9S5BJeDr8lH8AYUWgQJgqxEX
ePGyDqoj4vcpxdK/Z8DAFeFTmoUJPrp69oabp8M2KRj9tF7POGDZ/L+PoKmnN7OL
MBxktER6jqLZ2VRls/r9dy1M5difQSM4PuKi0xURxSxJtj837myMaCW7CYg8KpBG
vrqr3W5yW/LJN1dIciITmW19W7e/jM3m0IyAP+fGtslQobqZgI9CRKL2iiL7d6/a
z3HSgqM9/438bMrk9JkWeLvtU828I/yFdOSKj+XFlmzLo0iYgqjDRMXQigcdm00p
SLQHXHIK1ESSdh5UfSe8WCCbbcJKNWg1kRNtCTlkaxj9N09VXm3D/11s3qj5qlIP
dRO37WJKDKm/gMZ3+xUEDhz/Zng8Tj6f0xi7dRro42pt9xpGMbkvBhAW1CjUbyFp
SAGGu6RG2Spm00PujA9Cjec6BpU31qXL2tZ3KAdt8ayi6cyKah/85mL0FnfUiuVe
zAszLKWfNPcRTU3z8txVqMBn2j3egyVgIEo0R7V70DXbC8tIFmtsGpiNyK3hkA2q
LfQD9ih3GTK7Ud6cCc9fhLTkzTjwTV2ajiJG+kBJw72+d53NAAXItWgrXK0VCcXr
oN6sH8lQC4rgesPlHDNqxpGDEXihLDc3xE6r9Be205nNm5JM+0KtfRzhl1XIc2IE
IHxlK3pzROjRc9o3X7mYMUuhbGQ/bpn2Mxdp1n04aKQ9k2kHkbSkiWbNTKKYKqJb
he7BrA0lZHXLatwKulwbnMnZY95oN0r/C8A/M5wKIElD/wLXa0v/YJONzLvX7/zQ
Fp5h7KImWOooztAatx1k7PWMyvxPn56nbArbgsHAIsUQ4wWrg18mUln8BaKpEfBR
xmzEtXIGCEAi9M9JpxsOURnbUYGIhb9MHu7ZOmiMWv8WVgPY3oKgQNGhsb7FhAG6
eJIjCExMaP/O6tyB55Orf3Mzasy8aEmCZ57bXWXqNGx3DnbEVFI5rk8XZOnEVf8F
IszXMVJZx8u4C/XdfKzq8aDlBLuoZv7PVpg7RgCCtNz8B6upMCrwE6hb0ZYmryhl
6+eLvy7vxlK5Yhtglg0jnC7IBisKvKJmbhkou+pDGPaRpTve4snUH6m/iA0HFg7t
MaM/JudBMVTIewEtwDkQpbCZvkmaY6P53dcYiqcFjBwZsdQ4dj0N2/RE6XuuVKb+
hRgp9i/yUjNejimnz/j1+3Xkan0SR4a+LsSWyRSHx/lckrh7o4xKfF0YMufAilob
dznpNw517/P8BUC94ZOTCFYYJXwjIt2C/rjKTxlyVm4dxXNDdqA/8n5TV1GHei22
mbBZHea/LyL0y7UrWkapbUQLO6rBkI7Zrl5R/akj5RLJIeKb5yn9lFdjEGgF0Wf3
5//aZRZQnc3P+FoXcfbQvnVDkKOWg46nsXe59/vJCSCAIpa9OIhvexGyG6R1krMx
3UKjlf8fWV5VBJiwNdM00/jpBtpDnB8hcxI56BvecGpPNxw7rqNZIddlWb3q7tQX
BfsJSVA4Uy8UGwXqUu/Lby2mBj9HIMrBMDKhIG4HFtyEDLXora4vWwxYVQ9gSuu/
yZQ2+6Jn0J0aThyL0zRr7glmakssNMnW2w4WucI1FfpjeeNriIAMu0/1LvM4VsOI
W4xnem86Hc7S1V0yzcGsBTgT1B23X7THVjo7svbfnM+fAghAoE3g9qbhQ3xco0q8
TUqeCM0mAlGFHI5iK88w+INxsGQ2R625o5jvCyYlZAuLjyZ2+2uzZKTeu5+Rba+4
cVhFx/ZGVeFuBEM6phVdxR4b06/D50XztX1o4B0v+suCHt9SBqr2cso2BnMTzzs4
U9YJRf2yuZ745KH9oyeD3W7GzeG4/HJOjNl7kmGPR03YqKg0tSgP8DZgW/zrjvER
6/spJpbYwVd31iWgUryc7GblyrUISw1YDI0piMPItEycIYLT3URmBWTFcozwewN/
qwga5cS+KcF4gZd3pYSXCCf8KNqgLtPrnAjyxSKx2IREPKTwbgaBPRO45BZK7u9a
HnJNGSe2BsJ5nt2xqAqP3fL94g+zz/UKuWuNi+D6zEAOYR72iFd6pzOe+ZOjSIcd
eJ0PA/xqTWuAo7oDG09hT6rRWYfea2Q/8Hf5bMdSRh+edu0uWLc1FAIelsltBRGr
26NygDtA4fjDjq8E+eApVa6OSwwb68xfrBhicegrpvvc+xuPf28y1AdJynXCfw6R
JVF84SHSNtq0LNabEn1NB6YHiAxiwsc/6N3+K8hhmT32aRw0DoG/4niH0l4H0Van
j52MiV/jgPH1J0eAwXsaJ5NMG/t7R52jiqCHHSY7YO+M4s8rF57QAvCyPw5zd9+N
3MuiWDloCrb3bnK0NDmvvtkaoCJQPX6GJW7wp6fibt5tKGDFSEDwa1iroLjkPvQp
fyk1bvXZf7v+IIFkAJEI2KmO+t6Aq3uPmSvR+P7YLMYdTdF1G7St4X9zRZTuhbCF
GDSplND3JQVwYiRRSKYeI8xNCsRr31qIlndXh09ePthNnf415LoKCOVKkp5sFwpx
ZQLWILlysFh7txy8LHOKI9ZlPngKLaB4bItpEmE/RHaVY7JgHsGI5TjTwbKuy0ZG
DOV/go5oKMR6yjc2gKan5nQTpAMU60VdCibMXFOSu8RfZLU0IjzAdAc4O8NLi4vJ
+mHxXu63J0g2UoKmxcdijbE6ddYF3kVEbymaDG9NuQ4e/BPOfVCzGIYR6V1ROCwf
Sm+x7/WDErYXZ4893vFi7jFoig5cqL78Zw0hXIiLeCLWf9KVE7kUdNq2R6DYMizi
CJSzLdLH3ztE1PQSpNQ9sQ/9FOMtWz+aAZHjNkKkiDGprn4iRh1TuAF5PLHOgLTl
kEoKaBTuyGS+6n55OS37gC4Jg2DTsEu+f0Pj0VUDt1qJmZND0GClxrIY4Fg4a6KD
KtcYoE3Pr4oIgkCGE7bo9o0AG2Aq3I21UsPvDNamRgCjhOEVVF1aP+XJZqQQ5Njw
/PhhrKH5enm94puT3UZgdSjyl2jn75wrROO9JtCUVlpk8yi48ncyr9dEOuuGFnCu
0g3Z/ism68BQYPFFKCYFYcAbthNKxCCoeN+rcNaAJAzMevb32rBlRI+OnV34IKVx
1vCxS4whgdxdOH4+OsSNlPMcJaMKcwNsvGECxG3pt4W2ggSkL0C/6E+HhOPWP1e/
/ZAcdd8ATptPRILyMZRp17CIclqCkBzhKGzqMagCoj7ehfB8Gc1uISzTTmJeRH0r
EVSrLWPMLB824PTZk9BKrgFuwAudGAUk6p3OpCOVKR54SgTIA1oWjm3yvixJ7AQb
MqTN4GlibGhYxm/J5Dsvkzwkuv3PDLJfb7Wr7n998+kyG4MdP6qpSmFGcTFQPYu3
YfBs5kigIc5pJk6EmcdhP7XptrdmmEa+PkXEsR1x2U1F1to175ltF0Tas9w/bt4a
PdHIzkMgauFQiFwjITQTfU2ydg4NHFPm3JnmWvphcvHTHazSKN2D3/2YUidAfoRZ
Zca0i5d2UUbV12RMJkvZqf3+otX0ke9woZJNFJYF+CEQALEwgpkYG8BKvxQpHngi
H+k0p7N/P9Qr3mboUiQWpMN9VVIOdhUs6/aW8azWZVj0VCPwfE/sXfVMJfYOdm/m
KgM1JofVWqxbmOWyIlbLyMu89dvIgW5Xk4/AD39/Ipg2Wz94x4bmsfy66roWkRd4
Jkw7GW/TGQaPgtRbLlvp7eH8c3zwXK/4G9rDpnIm1SzBrSX6fWyGC1tMuOLAicGy
SdPnypcniqeOPf9vWOKUw4a2Flv12wvLdB7MKE2YjQ5ZqcblxNd85rFe2RxaaJXo
/yLKcxAlYr9z7Eluw+pEg5LkWyWc/mEVJ+4LHtiPx6XmmnVoAjjPU8yuui2C4X7R
4ws1eucCMB97mrbMXSZFi3e6wwykM0r5K032GhNAm1T3DavXCwK6ZGemJL384gnk
xqdQVDm9ayjZDTM0G0FanLfV7CI6qf3HcO3isAKQi4Wc0SKYu9MLAnRhA8DLbIPe
Sv4JXmew2uxoAsOCgGrqASrNaSG17XLFVjfGNRUxkDCZk60cjDiMfUyYUSTmIKsO
WYAiYAdJAtqMF/DFrfqXrIPmWoiTs07k8ONbFDiBfwquxWMQ1phMLOoPTsTn4y3w
37V05im1JLiS4EqNWMIEYE4DNORCN/ZjH4+MPZq1GK46FPzDbC8gjpnqE8Agf/h3
+2v3ezuj0pC5TjwqlHkcUMRsAgKWaxP/u4eEoblH10mgqhJiDLn6+1NHB6vNOxNx
1dfW2ClQAOjTjTZehhX3nnUm9SlGb6icV/kwRvOb8BqPk3x/DJhDa0Q9/t9xJnx2
k2D1R5SMH4i5a7HNaj0VJ4IPYtodoV6xuYxZ+0DOLOrqnjTraLp/RN3Cm6lDSoqz
LCT5I9rU7EXR2NQrcGPAqFt912L6hjm+qC2F4OVJd0Og5d7nqmS/3tP65UoxWmU/
sK84XUOUE6xbUJmxRvSzLLnfxB203s5IYvx9zU2Ft2HKjfjWGuG5YlpuVvNnojD4
bGhTqs8zptiXPpmqtnLEkIyrb+oeo1+ZMx/s/ux2toHSrQvUDm3yibtA6jE7OPB0
qQ62exNP6hLlt69AnBX4u7mL2vlKqcTEHWmaw9Gx6X9n0DVHptOJI2m1eTexqN+l
S8OctuVP9B01CtI+I+hUtk/BdjL4JDziBvu6ARLzNi8WpOlc1+a7teqbKPQUylm4
l0Mt4vdX/datRLL3Z/dCrzWOoE7v6xZwa3h7T6ZAnxp+6jj3wLoYU8VvOQqbXfum
0lz+J+yVed7DgHIfYXgI+RwDhxelCkDskY4WIyMtalmKWEJ5CP7Jonlvf4aWw0I/
vhx518ayA2+FPefUtlM9DZN/YMNh8zxnoRcDeEPnOp51ATaVMDJf73j7bDlUQ3jB
UK3XrmCcBkKnlRcsirbnHwYT1RUnH3itEayOBzcclmHHod/v6T0AdkdF8ogorHne
YcTWka/YXlj6T8BMptt1MqMRvPK1l0WCNAidXFjwLG7cw7lZKxUM3qP/kfiSmjc5
KOhMLS8fI2GqOG9xmZZCvDna2wKNgTZQfTip/7PY/OK0Sf9uyMek21rAIB7l6gCx
rXLCDLO+IIJBPBmfpKQLLHX3ghon/2PeeONNJZneFtqLA05Ezo0uFP4ossPN4fKy
O2YIZd3aeknEP5KKqkb1ZNCIdaAaps4z3CL3gTKQPbOhqBf2NOc3X9JWWE5YTl82
u5ltvMtVu0u2ElyFGbB6cRnGZ55VoXWFv70OgrtkPpNeYzqDC1ukbdTk5s62s4I3
gxTKkQzLSQu8YPfLsFpH1tSv+tlBB75xjY65iiyVXoRtpM3GCYnUSKnwmToxzoQl
EzErrp4hSXQyjr8WOJaFjQvJJJb51yretiBO/7f7l/4otB1GRyM+Zm+IALMobR1e
liJaV9bTcdZxZE0+wW4syZ07BRdCUjsEW6LVWQlre7bk5nTgw/nqEpzLEaAETcPP
OHPCcEcBQjAYpQn+Czjuh37zL31uTCjx2aPJVfcRU4lOZGb2pAdKBZrdWO6lhuZX
ck7ElJVC514XrT2zBUKBDCUoergESOgMwjdC63h8jiPQzwLWoRSfBFAyWCz0rwbP
OYZZUD2V0RR9xDD7y8tCa6ye6Z2qFTeusVagHdAVzA6WrpGvnuh5Z8j98djEU49U
VSzGm2RLd8mgVgZkUmxzPLEf/UZxxiYrSrOCm4rV2tYLgFsXC67Zt2U8kDx2gG5U
yDZPeUtkl4g7WIfPPZxGnEp6I5zQiWXpSGNc1ohiAXtX879yoJe7rBfMigqJmMp5
W8rt8dQTl/XNWE3pqoz8cMrUxyhP19Z3nlBxWYRDfKLF1/eca9T6jaM8C5MjFVA0
YTkalseYvACxn1j1T56vAYa81humI9CrqafBzj13cjv0CMaSZQObo9LR7sya9ofO
ujXdMUbGRxjQlj+4AgRJM/m163m70coS+lQ+iuqLc+k9IojQRnlpfg8NGoGWdfnw
yribXIQxFhQV93dBe3/pZhNzHZgI8C0D4OHPE9/2sa7k+TI5tniV9AFd1Lym7zWm
LApvQmpHyn8Uxu35vE7D/Nf+hXD3TVYjAjWjEZ6P4oIiFUVBv91lIuA0Mvip/46V
0kQt/BMSYrQDfGTfQUmwPjjy5LnkXWSSP/DWeS27JJLXjec1NXVK5A9xagNoXTTP
BBcGK/HAm12Untz21sfcbdBgMw1/gnOjIaHybmgAuekDesE1AjRTDd5Wv/zMXLEu
Pa/nCGadBZ0RuR1ZYc6afxdceCzPTFxynBBZpLqYRoYgfeVPe4mJdGCtuNKfBw0L
GNa9magVMNpYQN8uQgTyCDBjZaO0kUyQux1RiiPzrhKmaI1ppZYMdt6N9xq15gs3
82LcuyhOuQd0lEtHdlwNIFmA5wJYIxd+VeJEPwgn1e64YNyoHK3QUVvlq1GTml1/
olYtV/e2K2aimt4jR0Ux+vn3ELL2CWI1MLPw9VhZJZNcJcLnPEnlbXK0b88PfP0K
uFfBMWmidiBlp5P1GSHXTelM4R8dMwB5r6LVRZnjb3ftGSsjc+Do/Lq6qwgPtC44
a7afgQ0DQO95dk7nfM7WhqyghNMiylmdDu5zZEYxx3y91Yx28OSOsg4n1CX8rTZP
Laovb8xd4P9KmOD3jm/dIl2BpR9Yv/smzL8QaBSTqdXdIc3oNAxRBHeiJMDeJl5S
55bffBiRA9+MPsfibKYECAHEaSQJBQU6GH2HxnfT4cGZsk39nApXnF2wlaYOjBHj
+3A64eWy+zmGP0TQ6ZfmHH1kFXILWPl2unEdKFnnR+zVJfMRP/Zz3alZps7WPKI6
y9oNUJf0H3w5p6IyQLD6P1Q9amlXTpP80dbH6cuTIuts7jjwJcIHo7i81NCZUGva
8uf/K7DiObDlTVn/RIP0pJQ8c7cpT6LU8X5qteewjY9o/sSx9QF4sZPKgihPJ5K5
jJDzMHDBxxS0iek6cp2kJfXzUs0CiPAbm9VjqpoxA3TOM+5Une1Wx/WxDvUyiJ6E
aM+vM3MR7LzfNBqoBIWJj3ZOQMbhLHrHI3JSmL7OAulNW21+nRou9JN+Ue1pK85r
sATmwrAswrqF8n96uRL0qdJ70BwiA/8Twzv9XQWENZrTgsXPwtkpIgZ3vHwVTTfY
/nAoem1PY0n3IwiHfE526bylROOiYkdpBLsl4K570NbgKAa5vf34k8P6c+IIT6l/
Im1l0VhbMZE8ljfSlDtSiYVWyWZsr9mq6Y2u/IqwTAbPeU+P4mFiI9lhKos1fbuY
BRqlFHpCjbAvSaTcWkXIXJ7d/fsFSs+kOB9ZpBVXHhrjxGN3mIhhkBXvokq/Kclr
SJT0bu4gB7kI6spcJXixi25Im8ynQ94MYBDuvsNTY9QUtfS9ZhVtl2u8o4QunrDD
WSA5D6akzsNhPd1rdZcLzx+JYW9MN80Sj1XjaeWor93zqjDEdZClPQoSrWGwoiBz
m2JJYwYBkh1F/m52atB1NisLuo06Y3qhDXZ+IrM+mohRuTLGoxQ84H7MQkfw7yOI
tWaoG2mxZrMs//c37BjcMb53swfeUUVtuBz/c4C9x2Z2iTCXeUYSKePJrzF41sbQ
HDpN93t0Y8pQrzmJT/25cEdspU0GvnHH+GHWFnUPtw/fXSp3VFOHjl+Ewt1BvLaT
IjXwP5Kbj9R+kmmexO3pWiz0F+oyHor63xD3/fmVYmL6lH2fyArjrPF7fJJl1Vbc
s0qolNrKQ1lZCoY9xLjULCauT8LMGIRWVzUMBfbQq/WJfwvZ1UQBKkOr9e91lrbE
uDmuZycrb6FJp/LBW6Y38+ayNP3+795nxRAY88H742Zik/SGdxfkStHZEug798t4
XMQimZlov8FgtbjoPPi2RL4LEJ7wWzaYNtJOkHkG6P7utdfCEiM8GrML7PWC3aHI
GxbemyWX7pCO8JfxFFksoDN34AbkPOdMV+2iVCb3HF1z1wRmW4NctZGxIBr9REvv
2W3E0ZyqamICU7V+5MijRVeg0oY2yTJ8cP2y7k4YaLdZqyzSurViTcuZKU0vt4Qq
x4czJzacMSelx3niBq6lvtGKATCECuTfvjSWsh0UUTnD3FN0Asx+cTT69+9+mCI9
6qCozwFIf1wGpJzFDwuuF9zJ5aVL4mDWjZFi2omY+gSwm94sDJHFI3ArSkOsZGf6
4FkAlkPL6Cz27lY0o/NhosC8thRPAX0oocQAWmaqDzhQDk2/qr5V7sgCF9Vyazyh
p/DcLLYADvcJYsNP5LfdZDfOAaEQ9rd9eUacAaKFGH4qTBqdr346jKfOoRiLGeoX
fQ28fsdcDhJ2MfKItKBa0V4yvPhJqX1GvcSgNXBcm6pmjZF5J36nRMg719asvH8Q
+uP4fmqEa/IeVGvmzhbuEadaHJNQSn+Ad6aNoUHL2sjp4lC7+LSC4BHzJpFWz1rV
ZeB17kb64B1CsejDBZss79psGGLafHvHvv0h1sCF/Of9n++B8k43xVoUmjBluKWn
V/qQiGjeFLzXjcEeViz7wLj6pszZ8ESyXhavDivdifp1vtuKNeBmHqJBbYr1zJUf
l7ZXTjfg3D8zsJ8YxIWa0uOmbHaTnA1KWaCO8tzECNcWtnFseMyVd7FY872iI24f
tEk/fYfehK78A4N24EBIVyh65eyNiTt0XmSDNv/SBCChLXneocFh6uLlGuZzzrDG
zsjT7lLXzS/kz8N2H7fU87T+IrEY3hO8J+vAcofgQ3HnqZkFRuYbXGRrZHh4GJ5p
Egrqa05g0yTOLhRroDAzCeirWcbIZudCTvKWiZC1xCX7ycudKJRuRZChnSCLyG9r
73Sj/VJWB3XzqsTWxVGVeXSPT/K8GE9DRYcjHlD1Jur7gcp3hYLDjyCp5Q4Xl6Q8
Upfx4KoeTG5/Q+ea+HTLmspZBBOqhqZb55NlaMJuco566CG6LQRPtFq75jxGS70C
FIzjeSkOgKFQ7nSI0R+6/kgdncp5iDmlQUILRoAHlIU5Nbi05fBpgKsFZSAXtP6i
hIdmh5j8zonHsGF8Imliqxv5GCvVFMubkiKsUXL4mVdlinnxXAfUZ20+iwq6B1zV
iLrHKmFIa+VPP5pMxYNP3+zHUoY84AqztKAwJ0BQ7EAGv489dvgy8ZhKC3cxtAiD
pXneoNcFM4ltqi/Mp/enYCj6M6Ihn4SVDnlnetTYDe6UZd+xIk/xKhuPFjq2qR3S
vwkNT6mt3URlg3oNugNK5oMGcaQ0EDHT5Uuo8xnRIFn0jZ2X7icb33VYtJTMow1v
dcee6vBeFy0DaoYdv056fQhUtmH4VLeXfY+wtwnToRMCiHbmQQ5N2ia2dLrBP1NV
CClrH6IiVCMauqHy7VSlEzQBHx3/1O46mjO3Yhh95aVbCR54WgwhchOZL/L+yn7V
hHrTA+XqYniPHMrCJZe8tiFiHT4TxnMGl+3FXjDPDO9aZNTm2zYiXTqV2hIRjLJE
ggOpih6ILq32DJB3p5VI2TyB7KKXc4fw3XFquek7ISMvt+LI+pPRdml6zL/3ndLQ
ptQjdct3WP5DcIB+v19qHraloECizzl9jdDy7z2AqgmEzXJ3cDzKl98YclhQcEVN
buihBtgGGFEkaQE2yHKcQ4ovwaPd+rp8uKw6FOf6CuSgBPD0LlnO2xAM0C+ryfVm
ljW+cL5dFkdN5e/tFKrMvurO/0Sd6/e6BUZ/1iEn8+Pij6lpDj5rQeVtxkXEf6Sy
7xQ6c8aivTvJmNUfEL5Yjozl+m6Y/aL5EvgsFeveW6aIYxMvopl4Ow0eZd3g4mvS
coz3+oSgQLhkB7m/JV6DydVmuFpZI6v+rtQn/Q6jx4jQdHy6UVvUh0oDI50l0Q3i
m/BlBvaoVrwkO3dtdS/UZgIKnfc+UPP9vDsKESSln8EiQnBnMmGvzBRk9KjDnwKJ
BPqxz2aoVaPywnd+U/JLX6KXSzNdYV6/oensq2Ccmh9/0gpDoQVk0yPrX0bWuY1n
vZYXZmWYQfSGBFJrocIDqxd/1ZlON9AfuRRPHHz2r9cNam1eC8ImXv59OHLRlR8D
TgRkAvzk0fXZALRUkxxEc7bn/BDdxHeBqvgr/xHKMQXOUlchWq1RPkh6JuS3yoai
YcsQSdR9z53ZnLA9mugbyenBFPshKzfPTVeH8LT9dY8dr2ruODfjprEtIvpUmB9K
Y8viBMOU2dbV6N3OGzHM+AXkjPzGJBBlMh8PLqqC9R82d4Zo0nPZ2Tu1WHXdKRSi
97Cjal2I6X8v6Gcw12Vh9lYMtwGhCgFZPvbSnZma4X7QOUPtQK04nxM803cYzahG
HtzR6B8BMu95hRO9ZKayhkiLfy2QssMq709XTz9vxDL8hr7ndDPPXUkf2OT9NigY
11Wj1bnJhawPrSKIzfcbXYxUEH2hbokRIDtv1qk7U7zu7FZr7LmwJhivoHQycIBF
ns1HvqFB4GHhkJRjsm7mHM2YjBi/UATyfOpouZvezJZNPxv2YMcZmOgbdyBkqRKJ
yAiy1EHc4GuX+knQaJuD2h+93kYzloC/kmYejP57leE/Uh5ScWW2GI6aoqIqoDs/
+vTPQ2CkzwmD10a3KIkNH9Xh7PWeaWuvuA38fHCrdkej6BxHhmDkI54/4+kgU7JO
gmKUvvOZ3yX9ejsjuV2Ft5J/qjifGyjsedeF0qY4ABHk2YOJB71pBQuBzTeQOT71
N5hI/h30pz/sG1E5O4UTO5jdqF5HUejYMgVYxJ4cgPswW2cW8b4LCD9jp7aUwVLT
FGnwqInc+i9yzKuokK+w3bj6jVFlyaDm2rjFo8ZIx5pNJM4LM8YyDDDWXk+mUcIx
O7m0WS6HnS6VlFWW/7N3L0oZUchehmwNPSsWceoF+1lk7sbKlr7BQQnaRf+DO8Rc
+H9MUk9xF5G3S/6FY0qM+EsJnseS6L1CYLKuhPyDRTjziK/RZU/xejSF8OXWYSzF
p4unvUSX+PlDs9NW8obUus4L49fP1F1USjrckHI1IaNgG19aoB7/3JhLsr/DRTWr
l87wzUo5qhTbHUAK4GhXCl6VVeGLqRZQV36pHHKjuavodLdD9h8lG2rGshFL0Vfy
edRv+zzIg48Y/G4C9GVnaQwCtzEvesYNnS4WV2I80OHngwdolVkpCcYYmHygatZI
eYudOXb05EGFh0UdWx/cMZRPdj642ILRx8KVh5HO1Mv4fe8TMkhwiY0gynKeKHcS
MJ9P+C0M5GAmaghE23IdlDeW8QxxfeyMjebUG3IYBQpLW6PxeAB5BgyF/bRE1FJC
0ypml6lTj2IHTcDb7vrtb3uWJPoUVuONFw7FSfGDpGU5wxu+IQ7JGTzsMauNqDGY
61Okzo82LqYy1etFXub5RKV5slMfJpLGioQ33o3ARALSzKIkSHvznZbnKth58KpN
YIaI/dMipKcLj3yco/N4fn72cXwhCo+jk5buUdGYBjCeJU9VYli83a1iWXn5zg50
gcqVygqXfARrxq7kQJRF5CYnpkv+rh3K4DUTlUz0O3Y7XREcwd5FnS9cLwXCQdAf
zffa1eQUFMQjeinx757S7cpGv2jBwmu37FmlBgF5CkCyCbNfLU5p97pR/VqUCMSY
hLu7zyFSjTyW6yhsAN+/mk7jzLREGMCljY1+XIwNpL4bXNgWVHi+WSXf3QZdjE3/
NRXYVk26uEfsz8I1+KP7dCATbtRzriDYlQdfP0aPh8dzEQMh6LQLpXlPo1wFjh19
yvwBW+1X0SP1BK0q5yMrI4gIlYgDf5XvgdAAfLbJgl3fuBvrYexJtD81BkhDgrn+
cu05IUPvHzba9G9Id9X2w0AweXRZMuBTygd1dwp4ZG1Nx2ApL9qaJKTdqBBifBNo
1qdxvtHv4bXUdM8NlS2H7ZAnoPlaDAKgvP7aSU/hxvmJqUGrjh8hEc9H/PzGy7AE
TDPwrM0My0YPvzJZFBlU+fQZ2vKJhlLqB85aoJoDwNEun6h4DN+KfZ2xC8i3mKgU
IVIH20lLbngDn2VRT5TJJM1tc2fDmShMSV3FFxygTRLbUKRCub/V9H1wlwt4K97A
zj8JIbjYVDcDHKvTYNLrWsw7JsAoFwtAKNdx7hqSfCInBlF2YaH7RionFD6xExel
S7YNBXJOITA1u6L8wqXo7D4PjSJCOLCG2+OZ4QUaAx6OLp8W6edw0rBDYg3rzgLP
og6Ogd7lOX1lpoXkRfuQ3Sr/9YkKa7XvaW9Gaw4BqNtpsRl7PIETbmTzT56vVnhE
kiPd2smLYibnDHyUBqilMZpAVVuuiE0/NFoIPZ04leYLGnMKN+MucxOphXrJsKpI
8SlL/f0fCc7MOAZ2pZUSVm75uy84Q7cmNn9FdF3z0jiSo8BvD8yxAeVcKTfQ+FNV
Yi/1SbosIPk7Xk0pSIIP8pgmeJjSbE1xSn1stVKjU5P/XesWCD6U/NYtub6rFmbf
ro59qs/AKg7RXo0tOMFnJP5G0rSuwoD8EO+o6FiNYWz31ay+AcES3c3y5CmXrU6G
Q7mgQ8iZiVf5L2LSS0dHzvAkrqtRh9ktlp+P325iIqvGzLQ9US5mbcQufgdqMugd
sZBeMAKyUJg4PkxziKSaL7Q7h/Mvq2Y2z7ixQAwNJI8cyRSsk8D94SWy9UbrPxAH
/gxDSYeUgV8zp0RCuLfO2jDHPy2Umh/pF/vy69/ng0x91UvUkoGI9vFkAVZLcydk
1nWuRR9iHJxU4aO6elLN1iCgnZsfzDr9GXNcZEOd+aafh2078lR9oBW2mIYwizsc
pq2DVXFCtqJkHZu/Jw56bm5t0EEq7p0dpIR2Y8fW+jSoIgHOznb5vp60V4TKyEhp
6AxxuxvffQAeUN9NjpOIaHOYDyziBgmAIOmxxoTKmqE5E6A8CLdSuGI7NLBlfTHk
/vey4Pv3IP9SciobIQkueyirJN4tkxcx308pnCIKAoGxP3k0ckSYN4WkNUSrRXfF
CF1v5LbCi/IlgD/G1L5tVdwsDdD6NMnO+zr58ns8ATUmN1Uok/7U4eOd9B+tIT3c
Xg1zjNTnJFeOIbYc3oLRUbHixGnt2pfM65IjQzkNnJsqPdI5gEZPV6hbktWmmAC0
RpC1JhMZrWkGmu40vjPZHs/deReAyKbHCCMPsVkZzsM9ohdfGHZ1CY0ebZIdGH9/
/w0Sf+AGYesQFPZsazb7zT5z7XnHFMf2BQliI8/Oj3T2NKWMt4P7leEyBRphJDwm
PWDS11L3P0k3L4fqVOCU8jZemVsv/AlN14Ar5suMaVlBcLh6Cp6I9Z9+XB0QhhNP
i9qj0LfnDqgJSKvaOQ8RPzyMmGB8kTrFT/UghxnVRpFQk58L7Wgadp5Aey9LP7JJ
dAnjzRcqKTNlBpZ64t0Q7cUoCEfNOYX6w6Y9fhzWASrTr/OjP+MbD3l9HsjUb+iP
bLbvPmJZylXRAVACucszAP1nGW/kxj5QXQmxjVkcovi3OOzyw9Wbj9KDVo9ypKRt
IbMOqng/VM6FQrvucysUKfLEq+ZDIH0Udr+acP4n9cYbJ7S/b9gBKfP2hp9+vRnL
rY3+27U3WGIbWtdvlNlWLvcm8E/ITmtQtnTg8GrpovXeSldxL2L3xZ0gRuGJNSgT
+npcF+ie+HrK4tCL+Wf169Ucv4EF9C28prTsXF3RvT5ocBfteIxg6aCbWbUpnl7m
iPxvI25dWifC37FyLIs19TGPLh53dgdhJhMS5KDIUZLKGwz0GgpMlqeVxR1gp0bV
NewxaQOHok0zqIJiFVROnqvqXvRSF/nGzAhYPWC86zVtOZUDW4iAc23sOMHRwxGk
RA9LTYY/UFpMxJV+P24pghJrD331sDADkRG6ylDkykvc7OG66ISyhRjihPVxDXki
VqOmbspyBBoL7zjfR0lvy3/DQ1SAPSbIBjFgcJGME+NpXP7EOhjf/WUVAK/b0xFL
uGDEF391Obm+lJG1ZIipimxZvIEuFnftwmwtU5SRmuwwmrPJ63dZdjj9EBhN5vEW
wUH4EWSYAcq06oXUeVyHfacSssZs2fHBf2RJ8pvEQChlNB/uwoCz5thhyYnV8nBR
3dGOzp2FjCBOB8/FJgF3gIGIi7OSZtnY5VAkFh8hmJyq3CKII1+QnfJKkkJ3INgI
y9Da5mSIkMS3oIvuqqgom3UQhDtKbVOFavF3E3otcRUciCFhVJ7Tii0lURDhE4Mo
ndBHjqRG+tI9CKFSmzvxGR4uyvvO9mOVS25DR+Ilv3srjgwxTOlyJZl+9JkP3irP
P+1MUQ6YjH+ljQeN48p0YYDk4iQiorA84JqP3U/egPGTXlpnMg7ac8fa9NVLjwxR
LsciOhxWJEbj3A7B5mE879DHSIkgowxVsPRTzEuafmxP0DrnmvMl7mhHX1EkXZtN
VW2Iq5Zz6sk/cOsLdGQRPHPAUUegGnjctRsSx65YKQy8Vlx6vVD/ZJtzab244CZ6
SxHCBP6wwM2rlwlR17PTuaaCSDaufow9ABjqtAxNlTQUh/8ug526bpBkdU+DzDZg
+YrATVWRk0deuifN25LiGzlMkk1ghex+/hgFmlZwHZKE4Qp/XvApFVmO3Ff932bu
lEDUl+kCEMbX8ZweylQLcqWH4V6yfnSgEB82+u7Z/r13oq2V1jRUbJ4IdlbgNMkl
/0Cdpy/zXqAnpDR/viX9ZLXVnFhYCO/hEz6Tl5QtEZAdeEd0L5YEw+9PKqERNlT4
56cTyQNZxnH3jbpXRiH7VIoHVpW8Hb9hTeVsWhtGtHfBJ0YTZJrae2f4ailpGvJ0
6rFS9YHkQfERxQUKimWZycK+G8O0jBe/LdqnUndNH0lHXAQ9SYZWINR/JqTZITdw
jCcoe7w1Mo4oZaf9tlp0HMVcgrZgJ1F/B78MVDemQHc1F5HapDgQSxwyGRKIN/DL
NoHgAQ6T18VHJNBNU2BbLLCUm5WhS9/h2gQtgISrIGLtthZg38bBrclutIPG52aL
D3f1/ckY8Ls07Sa38G7PofaJDANR07DHcWoOc8j4oNqEYUhCHoI9rKQyRORK1su7
rZa7e+XY7mWm1EymxteheqezQ0hqPQucknSnKkXhWeeTkgHocgQ+vKD2lhCqeNxK
JxUfqyw9zR48dYk8doV8nZBfVkRBO9q6jGdSXb20qiR6R/NzQsaqKCDHEY4T9ACO
+52gEXe66I+kO8hHiBupUIyoetH8wm3HMrUy6xJ9LI3Q6XJKEMYcIo08tyOeibcV
Nc+ivT/EVP50t6sMFGlq0FEh2wlUolo/hGopgUdE8/SeKgD2r1BOZzyz4iiRGiT7
ZKtP7JRvk6mAumfDKntrWgwiW3/4+9k5mulsDJbLNrLNuONvNgpLrHM7s/qaITP6
/zpM1q25B0zURxOUV4g18Kaq1fr5OTxKjGzmc/QVs0xSPZp6h1wxCUzMs4e4a7tz
JRbVfxZEYSM2FmtX9r/MlBAfLIAIO7K5TOpDl2cEjnDZtOEm8XReInM2qkB4KIVG
Z1U+er3kf9nKRyP5IBDW7sRZ7/iYB+Svyn/aKQKOCFKCIgM26KiNGweav3OJeEXt
NwgJ01Aimd9Wvk34sZab2fzsqXjtitbwuwfDwV5YLUX+kq9efgeny6BwxjVg/AEK
XXQZs0CMid5sEnXrVnKv4t6lUWjPzmgz7tm1VVT4LCBYR1exrMz0YrwWHDeeJ45W
AWt3GkPzEMn2/o4K6jHxCw5gZokXXvD8zQO2NnZriNuBL6pVRzN0o6X13lqjZPSC
cCW2OWG5wJtQ/N5m6wzRPfFc8+l+0yJZ/93+S7guHE5Wnc2OPWc+qSh70ok29o3H
jk/jjZs1LTRk9D7YrsVpyi2waGi8jOfB3jmNRhrWHtowjvvtiPdObLMKSWNV8oXq
7saq0WvB4jtHOfCyTIYaBEeIfkCVfD8NvnWDfTakrKZWxGYfgl2u+gKntRFVRaK1
zw3oTQNBXGHC3aBesh5ZWsjvTW8VDzEOY+xa+l9iEQSVRkl/fxRFRWSRldzAUIpT
4pKvxeJqxuZJRMfigIrDvOPbCuYq96okQGK2FA2Arrk/TavyzduVZymuov5hUNsf
1ZFl/9cua0hTFrLErtY2j2UnAclUDfhZv+MgPw1zeX6dMGA7ivpmg0CgNdCnmMCZ
7kGWAUCp0IO5Vjfi6BKZokuBEcay8aMSc93u0ArJrK+JdS2dg3Kfvm9bjJThTCbb
ufKAfGfMNBWXh7TyhGSHVFlNKGf59YA6QARZGlUhYnPN3Xy2RRPQOCxmmVAo+JtM
/uO90eFq/SmPyJANFVQJcVUPTYOK6YEeaWazOO+VB4J1Ag8jna9jMF6ry6+k6Clr
EVQImwsL17a4FFmYHpLKHQwUxzJN8iqVrWfEMjD+7wrH4F8ff26IoTPi9RB8e5Ep
1he8DoSU6emSR/TO5ime7F2gyk+3zeL3ZIvO1qGkKEF09q1eL5dpq2rBWNRhhEib
IffTl6rTyOemW/jQJn8AInAdW4xbyHnigWniQZiYy1ZDQlnXLH1iqmI8ugV6woXM
SqA5wYfgA7gtVVJxOIXI6uCPyycynMASVnMfQiSRRWXqnnX3zGlHwltllKuuOCE+
XYXfbZvWN6eZlo1U+RMp0c7mfcysEnpc6Ek3hk+7jOqkCes9v7nXyUV83VvdzGVL
j9NqbgV0GOyNuEhj6+cY70ZxwzXGw2widssquHZmHY154t7srOYURdUTRu29vjRN
CSpaKYPTYDLQql5EX97ojx9+V8+D7pY7n6CnXPAEHSL3DStbhP7hkzw4YfSoQT3i
h23lovhk/pUDy5fygZIOZmolDqlozY1TIdRxp815HhPD47rviSItoZ1a6WzHBrFJ
2Gpk+PpV4OipvbbRlzRQtsXxbcJFB2AD7vXzwNrxDII9Md0uIp3Uu+uv2WRJSjoL
lxeVUwCo05hXfU+kX/Rdxx0uDmI6YazVWpI/0woivo8hKmjcFAEhmngGLbjzNU4e
BffVaJT82QgsYlnDVzluis4cnjsGkz9bbH66zqNqMRXGAUqXJsLu2Jvf1I+X1l+k
sgMox1CT+0vISujt1WZhSq/lF0M374QRn3iCTn7e+qftprS9shA2TgKscI1z5AEx
mB85WKGsSPrvz5duquFLU3sjSUDUBhF7XVLWYQ7eLH+es4zcPeziwwzd6G2ZW96V
odWmlPRJJWu36lCJ6SfGoswWubZeLopnRO7frTvMDLxPXUhANEbmVgSZT+zQPJFH
DolNBcRoOB+QHEb6nTbaaeq1sByZGA7GRazGlAdnejG+xygTaKBZDuLHrXihL/sF
3AIzr2zjyEPgeqyrUGnPwi2wo5wZ13Dnxy+Pl90A1m5dkT/rThLLbnnCUcMFYwVB
/bDrw9rygSnrSMSZYsGdX+lZxNhllV1JQluJqKh+vdVCA7oAKecYztnYu2JkX5GC
6hRXK/Fm1ybXcwIPbSYIGDCasUoC0B9XuzwwKWSqZtfQdZYVgHqKnEPZLSEC82l+
cwTfMrDaKps6s9lBAWRmPSEpZYqvvsVgVy3pRCiM2i/Zuk2R+Wkf+R0maU8hB/iZ
T96fllbGUY7agd5IHbDh/Ouaww+k8ghjnuyB8LlyLti8hdqphtVvxwtVj+lOEPZL
6zI8D/vk0d+sFn15b/LZDbeAzzRQxFcYAnlui8nZglBVaByHmE+Xu+B06F3rOW7E
pflK/caV8DurGHjYOYe18y7nTNAQuVwxvR353M+/MnYraKpIAdzW8SbT9wPJgD+C
/q6EoOTS7hLXsAHsmhYkV3TsyqPOWJPD9FgIelmLlavk4LWpm/HJUhHNuDeXm9pT
VAJqZrxg8fAlTIEEtdZlKIOat2gDEboe93PZTMla1twfZXLts1OirYrpLz5fHild
Rb46YIqhQh4zym/34o4mB9H9oBaqiC4wcNFmVeElhYYd/2YorQgO0px8YUejFs6J
1/OIO9D2xF7q1mGSldsNDJwRS5pxBhxaqwp8kEqVBLNRe2pSd+AwxTLxyA3kO22Z
yDklyXYl5TO7q8Gjl+3Rz1RhybCxv6P50oBKotYK419RsnA8jF0nBIV4GAR3vKdz
tAptvijQ9z11jKK7aAjRpTWgLcMeF1yekFscZPmim41wIbeMm+3zQQNj/1ckni//
SQCoiDfM6NsSanT5loWp+MfPjai8J3tO0hUHhSs9eZmv995vqM0MO1GAcehMeuyj
hGqTdSX1Qes7yBYQJrJ1QFeH25J6XdVGfdUfnCuUY4LgVBHQ1HIpQ9oSWzon85LX
UXAFBqS/g5oZVjij0FGId3jVTZqfKz8wQriBHrd/UbnDr3LhPWHM/q8cYHYKeZxM
KEuIDjPHQdbjXRyaRSCQdvl9py3HutCkmKoUC7NhZxYmu0ncB/HdDph2XF5oHlUx
aounnVvJVKMz5m4DgPemi3wLw+bbr3ywza9cKUtmOgmj+T5Z7ED/LFPxS/y55CWf
L8Cawxv2+OjZ2pyizBmgzZl14uOG93DUjdE4XD6sJwlEZhwGZ/BKwgDLVGX8jbqU
9AtslaN0n8t7gg5rsSoSYe158vo0n/OeTbHZwtIjQIT3uTH9SkZr9q5E4gXqa3lQ
2EJtHWAWowrjAqXse75opkXmaKDu7KHpVc5e10MTYdb9VSRRIYv5pR7ump1DUEiK
Eo81CFxLQPjIF8SuDWBPh5taGDuYX+Q5fTvVbYYeZXi19WxEJu95zFRpb1dTMbgI
SDxrYMkKUUbUiQYFbJZjd3ccItmYGOvqRSdJzSc8F7h24Uctpom4n2iWBwDfBRN4
sFRYeIgxizQD6zXv3NcbHaSyD6FG+4CWvb5kYBKMWr1SGox2z+0pv3D5QlB1UR8H
k7HM4x5y/SnV1UBMopfDi2BzpgS4myPCLycPE0zovz1fp/KQnZ8e0wbHlA0oh7BD
FE4CSbdt+SM637MmnstoIg4l/lY2Z5zJmsr2xeZnwQFhjGsKDsCTfko72SsGm3fH
rKTlxrnb5znxx1yV4FbhogdDtUVg8vYlEOUInUwnZ/c904L3JndK0RXBX6+VnNoV
vcOKnK5IGLrQeuzkzCBBylmquSZz6l4q/wB+LvehyB20vjs1YpM1Sqo2Kzcpbi7V
8Kafi8tnL8cdZafUa7uGLpbTM7g8iyenAEHRuSHuhro9meWlfE97+R63hNJ+vSCr
bbTWYA6bXwj6BeFblSwKGO8DjU2SToHvOpos5hsdvmblCT2XjqfQVeBuwhbUZZvo
nxvZD17MSU3d4MFv462nZv5TRmGRg8ay/g73aSIFT4tI89HtyQF3AvduDNYlwkto
QRdKn3ka7zy7NKa6VDZiRWURtY/wLx7k+7O7rsAfnr2XonoWHGey8iTjJOFX/Qnl
xWZY+GKEZThPafu4HR4qjXWgqDaunG3q8dI3Bl4pg2ZET0S3nGECIdNmZWcur/Zj
yiah1hLI8LJGi2JdMtq+hBqXcBhiOICNMnUMi33d19NpuiafBxenAY3UJnLhSreq
xKQTqd+5YtcH7Ojhd5ywKlJhI7Jo7ihN220sI4i0j8u8dIIS2xN3YtnAOwLwv2Xx
tCkLu8GXRsl0mbYyxCWatTKq2V6CR+otIrL+j5U/ZFTfropjDQGzIHQLhcbJkLl+
farldz20TEd1fGzReUWkPttLoxpOz4wG39XuJfQQJGwQLq1K8MiW3YUDjDF8iKTc
lAf8OhULmy9A4Trl6UmQNcfpTkf4Ajs73Ne8XaUOtZIc6zHJxuwbl7WK9FXWgAQl
j+SUZlBs9B3xo+kL1z47jeyha6RL09l54c/fvbxfTcojRWEIndLdIiYMV0A1R6n/
q+f5XBVcheYC5jPzdgH0DtcJAfuOq+NuUOBTsHiGNRJ+S3EJVfgYJPT36q13LJFQ
FCYxqylIT6WWur+KeROQro2sJOshDSFp4oQvlnJtNb/n5Xc8pdpUwEz3/31st6D6
fjoVb5kAzA3MxsO0YWe7b5Ka40ijGluSIsKv1TQqTL6YDyQrWyiGkPTt+wtZsaDa
UrF2SygFCJvyUIAP7zilo2bZ5ahmP4HsTUftAt+DmFHjTMOPvyeJuE+1UWsW0bs3
Ac8Hv8Tjwg54Y5ZZWh28kqfg+CamaHzE57VVtNIYcLu9Rpy022VslL8TTOdjJBJ9
OUxZftVjPiYh5ppc/18BEaP0PwnQYi+4Pk/U8MFnjOnyHuDzHdbkbeyGXP/5flrG
emuXYuKIUUe5kbhYSnnELdUyJz+u10wm8BBYkzEod1KZ7k2NpdYg+DvWjaDHh41j
nd+F/z3MGdRcLLST/sa4fvGaaIJhf/zqxbESiquMrKj8q3wIVWQimf5MKhKQ8Z8z
X9d8xOvXDmHVi7Y4CpIIYVoh29tUnu4E3HP7TJ9v5SFp8VTiqvYfdjg5hqrtJKaN
76X3869sI1Uc0zSuAWIEPFlf3GyW0xO6of5FtkBhPOMB//DiUF6dHsWgA4qMKfgG
cDB4coTKATQLPzugCtSFOphvdl/V/AVfuwoouxNJUU1a3qObz4sfMaInEF0IFbpF
TGKhPzev9X3aABhrWuNSogs2Ym9AZV2833sz1XkDwMTEzZkiR032ILDXDr5InSYs
fSbNOpWgLyJNDAzz47YFus/laUDbf9InDFhBsjuXTff1+eOJWdTwYIGrLhlO+5VY
k1+F2j1+D8VI4/uqo7MijAp3cvK3ljLvJ+26aJo42wJ0SdoDPI417hF8mbnXYQ/5
+QKPksFFHPYP9q9DGwuKjMTPe/Bh5bbmDti+3SpXR++r/RarvK+vNq7e2IhEc6V+
appRfsN+WmydRmVCS9UbJZ5SrhqhaAgcngnVdF3T8Gd1c09O1nnRr01MQC88mCRs
5FWqcc7DHcgGCMmGxUWnAIwjWUSOAOkh24eQ4GXtQrYkH/9LSzmq4boWSgl6N9uQ
EiEe7Txj345GC7zp8QR4D0HneqtF11xyYt6fCO6ntu8pt+hxojMvHdbuLuYCmS6r
0QQGxVuuSbrmIZiNEb/ErAabmecpeIylYsmRY1cerccIZQBUjGkcc1KVR5XKd9ao
NEhRMGrB58ugxZG4SCyqGPt4cmo4vplMAa8BO+Tte6MINrxsGV2MwqY/yafvqHNQ
Al+dHefiuU0wMpPe/YNsmjxK2opzqVjEnRY+E7O8BqBpl9Kz7BxVT0FYI7pc2wjU
pGSc6h3Gl9KBaqcmHl2EEt9lhW9BtQCuouqZUaoQ3wQN/zfUtM0YcVRAfJMnbrNy
45JmzoYDUx6FGDmNAw2eIItK5xoqmWVFud6G3AwU9Rqbcg1A2kLejnRoY0nerxYd
DGiyuF8v2sE3D/7Pq5Vk5uXocEkoIQFV8+kfojp+ltv4pNhwGRkdb73DljXH0Y14
lrP7hXCrPesABtevztpKlwlcbkFE6g7ynIXfI3nTDPyQgd2HdWVG/OxfPylIXURV
6JF+vgQbFbhqbgE8xExrdiVov5jC66ssEr6B/oT9EYI8XftDmqoYzS6TSGEJ8IEE
N55xt55QBO/ofvCg8+kN1uoVwwluVNhAtmhc0PnvVBjttL6dILLEAUZBPgZBNQKQ
VaPe2OluOTECvPjWwyhcw1JgJ8F8HR88xbKP8zWDEVf3/bYtYK7MkHZmohE/yNFP
vknmCCmVih6Fg77Yf9nEcSUFtHrgeJjIB779Q2+yNUQQsBz+GaISA+YUARV0rNi3
/dFxFwTjGlJLEotbXNCPfHrvE/Cqnvi0XXm/TcKFNVzYJhQXzbWmAsbOPALbWGcu
cZrXMnQFNktpl+U/LRJZp6ZSM0gFyq9ssVmvtKCQMczFgNVJUZaXQQxmdkNmZFmp
k9KkQ6Ynv8CNLYDteX+j6BZGf8Ct4BXCdbWUz6VFB/j5PqAcbDq7Ycy4yk4EE2ka
HfY1/f6GDLpyTLokykZdEA==
`protect END_PROTECTED
