`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6sLOrxbQCOk2bkXGNPer7gZlxunBvfyWq5Cj7zlcdkcRU8h/toiDuQB7A6vqNTOI
krXdVHWwh+PcmAh7TNHylcw26d2CaoBZeF0g/z2vgc1HHrzV94efe9U8XPusqlCZ
jJ60nb48qTmreqKVveBqqOc0mgLMyPxC/dJ+6BclcK1sCp8euHC1UJlJM7Nk8lKE
2b9iooOPOfToxRH51KVPxJZ878cDEAlZ0sEAnRiHfTBmJXHdzKug10IVEalDKju5
m+utD0QV7veFYiOBzBFPyQILEZgXir/zceHCR2XdQB3JPJ2XfO4waa/sQb4B37wb
GNJc2w66oIZxDqhJf7ijEf7qD6F3Xd5ujt2zQzFpXovibg0h/GWWP5fzgvUVNPzE
2vZxMtL/puXUzM6bmdW3ITmydvF6ULILFMXWkDRJcr6aKkdmXfUb6tm8saLvNv/l
o86VIupTaeuvTO2FXVzL8Jza9sQYn+U7WsKv6uD8MGbcDN8qiE1bghW1jJ2D0UdC
XNofM/pOphhw7LMO1rrb4XBlzM0CyFF+abrW5Ch2ziGrc7iiCklE6K4tYfCi8qr1
i0irZSETqrHch/yiVHRNLQTOWCQF50Q1lv5Liu23kCYIuGWIbGPUlc4uOiekQFiP
a9hUXRTFV6UAUwU8n6AFkltk/UVoQhDDfifG4TGADKXneagKSCF/9HTzp7jxTULx
o6LygEbS1gMEtB68U4TPyFKOYOzCGnnEXou0dYA9j0RLbQ7KXBWR52/sNajR/40k
skN36Q4BuXSLq9tjwxOmWZi9Cd1zmtDJCWONsCIUfNPYPykQnEuMd8O9P3RW/dNy
lS70gT0K+jxrE9JfOhGuufNLrrlTLZVeZ5tYOpdOULgyt9TFrI9DtH8gu7FlSf1E
jAq5Z3Lut+OXcR+OTvN5pk9XS+ofycnBrwcxv50uq8oCKOasb+gFiD9PBdTju1RG
U57b93DQdgyKvrJmGgv7kp4GTx5LAGXKAZGPv6Wfwq9Lhu8Z0+oalFfrwdx3jXMz
ATtbSHThzpsU5p0fn8Cf7HlE7yqpU5AC5jSvU6+QdL6FuSGiKFWjWnUHZiNE/W2X
VjE9Y+qfyR1G2mk67uERU7c0+mf8TfNuJs3tL+Rf70X3o+cbFj828AbbTchm2a/v
S4Q2QtlA90LKOE0HE1L5l1j1P9yra+ltw3qInlbDyy/4G2xtghzpPMELjjIn8gvG
RvesBnase+Tl7rBzgzkdn5OyWqQq4CehMqjww0aCstbpR6F8SztdSgG7P73RsA1S
qw+qd7czysIJUpEsZsc3qE/b881IxdyIkJyRMcSs485W5oLRI6b3RgwRqdlRKrPj
9eNkVG+Z1KByKTnh0BEhJgQaG6U6QWL1as30MDC+XLp1tGUa69bzHRU40A0XDPi5
hdQfb5VwP1DL3/7DIiQpRw==
`protect END_PROTECTED
