`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8J5DPRfaSNADNdCI5D7riYsiAJxh5J8liFl0TEgRKDQG89oQAUsCsNFS8UWtrBNO
kBNKpgXOg9Goi4JhaK17DnQyNMH1Kdb4YP4xWcg1qBo8EVGPNA0v1Vjlat67X6Bv
tO72mEI3wqWC4ofXetFe3CYiUUFajbgQDt4WzuAmhDB7gcelEzhGB+McKWsyzIMj
KTIvg8LyJW8iDYTsH+zYsI1h94nBMlYGfL2rZrhB4xRRpXb0YmTpooCemG4j0OQj
WVoixNi2s87ZQkIlvw2dJyBDUXYf24t1GYxvV8Xq8dsJajcFGSyxj9yJP741n7FP
WyI3/FYKJvsHZ982lnZEcaiNbhfDOADf0xzdvcZzm7M87hXCFlpz7rynwgtIBMGy
kBys13StQ0o3sUudXYm6t0puwHW3prsPIg+7E6SxwLzzzdloFO0221oiOblrF65g
QQ8wRBsfBGFk948P9bqcA/TNTk+W1cjlanoVAH3yL3sqyeELM7F1UmaJhNnOlqZ9
s4Tsxh8ncQTlOvDrDnDo/W3jnTipgrJQNKVjm6QyDZrMQgL1b6+vtdGa/F3JR5Tr
ySrLgL6rvN0H8Ivq58N199ukfIEvz5WtHOgHWHRdeJnG4nXBEhUM9PX9Y3Zn7PnT
d2mICf5SouitPKpQ6w9g/EsD8jSKw/XGjRlGv6ed1/yy3O9NAks+rwoHZpXiFUYP
ECagkogJvoAO+DCEliQ8T7LbqOoiURGkoGdgXGqRshLtHBa5JZOtMFEpjo1uRalQ
TYNrXKFuZI4hhqjgyylahOwj4NDNdyAYBDm0VGC0O3SBT73zExp8ODRrEWLgGpVe
8TBWg0lWl9pSLtR7EKnCL+gHjhpJcbujruETEPCGlRlkKJatJIKZUiWNOAiX3mwv
9USP/hTWkS/TZ3O2pt+TuDwZS4nQ8MMDaRtIQLen2Eq8e/GeffwtWReUqwedxyTP
9nEHMRNrWG8qQ5OdqNu+bA/Kh2+ng/FhwQE5IemEoFlGo17zfZSNxU5DHepC03Ws
uh8ArRdOKLOEqRTR1bPdo+tiZI9BTcByl+ITooensgCfZnWIfVeSHuT4zFgEuoYM
l60MFeU0MvzEgCbhAu6vzOqGFxOOQfunVVobvYREPiW1lPUlnqUmyhHaDu+5X7yk
wkmCE/i74jPO7GXgYtLQvD3niyztveUCaBnhs0w+X2IOVS8Qe591a4M385K1Ihfa
yhUnKr8sdawX2UQGCUAwqvLdAeA1FfcNG85Xv1WJihLf2RlAF2oKxaHRi77r+T2g
hTaW05hhyDUFQIGZ5FIl9KPTWp81+muMyNa9Z6etndaYp43lUj7B65KIqhKCgS0L
g0ZTI9p6SR5itdQCy/lVtGuScxzbwzu+LjMJIW08OkclkVbo1smHJhGEjdBxLyog
07PAWezyoscezst8wAsV5uzOVTHuptEO5Se3wWKatPCjcEg+Zm8qnU45JbFAaNZZ
aJihNjnWKRSjWte0oOlfxyWmuXok7DDrOvqSdYTfFc8nUD6mMQGBKB9ZladJUHPQ
TJ+f5yzURBt0bMg/t0ZpXQdsiBGoxbeSzcgu4JtiLRWNe7ULZ15P8t/COxe/aWQU
ilpFN0x9gsaU+6tOPpZUlZDy8jBuxm6emUb8ilWeXNmGJEKv9y4+pi9T8ghg7j5Y
3O/Lt/sakHwTJbEHxamJfhU8yrDzAO/Lu0r5QrwGOkaIAze8eLF4F00BeKhZBz5J
47SZxfRPq5/jB8FGMyNkSFlG74BoharC9pD6OEcxt8R9VaIouE7uSfIeFfJ1rRvv
o4pR3GXpVC09o6uVEHjs9Jysl8oiUmSp4rEN3ALg331T5piyTobpj1e4w1xWDFc5
Cd7GM27tEH4aPC5KQRw3zJAhMGBw/s969fPLcAUd2K9EWsW7CUP1bE6/bmWk7uYF
ODvPX5AXT18lEsPlGp/byPvjIkzp97G5kACadSxgQ7BmtTeQ9IpQtjsx0gLQcMnp
M9E30zsk7NK3B27P+aLs0vRiYQwQ5L2PPg0sbehRGvOBLtnTKrRThYqlNJ/ITMTe
394gyMGXVPSKnuTuB+l34Nl53bk8W+GMMxpT9r0Eef/W8tOT+gu6JanDK2FZWjst
i5IxDscw1ay/hEiGBzEHrFEpz14Q00ccW2y+i5Ot8OJtJAp1GKgJ1i/w45H/pvz8
KwWPZQ6gO03ZEaKxSuG0gDqtGdOkdmOttvVnZipR7HbI0MFdDs/So4lbR1o5j3E4
rNzsFQSoJNIQswAEf+Lb4+mHeLzeDlNkP/T9Rm7lZmosw0u9RlBXm4oTAA5//1LT
B80ehDKG7plWCfKSux1y4GAWgSk1rqnUiQxPsujBQzfeAHko86YywYODPBqZqMYb
gJbNaSAhdF3wO/Y7+7jIcQQrpYkkPXGFl25oBCxngzQY7HZdmgI4DeaU0HLr94jc
CEUkjGnhlSLdgYl3LLjIfeHP+lbFqCew9EAu/CkNboCvPOOQv/va53KtSGIHNW/m
EuogBtK5pSSeWkxe1zDfQiSr63mvKAyq78VPi4XcbT2xazjYt9O99qjZIQoDWo9s
RtgiZ9KvRRkgmmssgL7WbE4ALZ8BU0g8VcIcU6icJOl13y6rdA5q4AWFfE020KGA
rnj22nKESp9I46LFS/hjW35OZiP6r3BtzpON6ZQrLDhJ/2mawrEZ9xos/Lxfj8cl
TFxb+smmRif/IHzdp0BoUOO7ZorYmv72jIm9ccc8ZR9q90Cx3HsZyHQEaG7JyNy6
C4GAJPpBaRV+p68RgNk+MgfbhEnNy115jV7KUwtzyH/1CEawRo0kLwltytfVWwk8
kWDVcFFkE1NEnRCUspV/ttrf9pnArm4FRAhjJmObCbkGpXq2gOsY8v06m/FzDpzq
+OVZ22xRtSeicSkGSK071BYkvsHZPmegPnmi1tRQVVw=
`protect END_PROTECTED
