`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mHgCkq6qfLPnuddgM97dDKFeqhzbQDelEeCHaimthWhszk9qW1i9VsARpP7ws4J6
pIj9TRZTw3l9zo6wcehq9b+ShHxi97cNlfve0fo5/lIg7YIVRmvevUhXR7wHNReT
4bwKe7gRABQVyrGDAu5Umyf+GHDBVlSqGJvNmoJiBgKvjryYo5R6JjRtmE2WbJsC
K8OaxNlmnh0OqGxUpiypYvCQBpv+/JbkGBhPe/s5jRCqVc+6hqypi0NgohEtTGya
BqXoQEJNbXa7ovPiov4+DcPJadeFTvSBQSX6p3S4BnIUMaYQE2lPqx/uGmioo7gI
34rGbsCJnlit6Z7N/Hj0hQPGZ3kpUMrVvpuOuqVU85/2EPo4k3Xzd0rgl46oF0Vh
ojUXwY1rideKH9MtGUk1ZyZa1d6bBO7rp9iFN9U6VDePVNMTNHnoQt8na/xYCDOc
b0Wb42vAnBpXjZsKHNG5YP0W8f6xrNcvXdrk0QdAIyprc2drrzm3KGIcVe2XMLDB
Ngx3hdlsUy/OaXjFmctpEGNosrsgZIJfbpsYvl24UCxL45e28FQEjQ3Z8iWnrGkY
+a3UU93YsB7RoRGJi0Ua88a2zSaxW8nKyXKWbQx1jhYjCLlT55mOYH2x0YtcX/Xn
WjIApFTql3Bo07jDwCeDBuLgQpWiTteaDZffbRBkKyYxa3wRn2aSERCqgn4KwCgo
HmrNnmaFBimHFLKfw318gS+sx88K1ToxbOGekhKbePPepywm4BwNAOxVUXtRTRv4
uH1oJi+uZxo402qQYfyfVcnH9O2VR35TZ5isMvkATofbxEuNkskWtUkY98Z0QDNO
8Kvz/yx2GG5wz+GsREtvuwnSvhkZoLAgwEumLMIVGVyRWaBALpzO/Tpn3KhUdgVd
oAXnRgC4yjNztl9mYuQQ83kb3ANP2UL/Aj/dHHbE3vIfZNtedXue17+RVYDQszG0
RVHB+KGkt/Q9wPu4MdOtkgpN/Ob9XjDGCGxJO6rQ8Ln5/WRWyN2IaDCsiuvfDmT5
g9LLGElovMf6KqHLAMqvKspfTFVWBmIDTouB7C0ZyRTnuinAZ0uXpGzUYVlpRgfy
Nebc9Gnv0opOUHpQlcv8QPHE/z1BTH74ce0FaeSjmnt3084Nd0Ih+Cr8Z8H/mKEs
yDgzxzz3n3iTDJSESSW/jbDUln08K/421FWmJ0sqtya3g/M8l0S1C7VHFttLj55j
+fclEoOchAujn0/kc0SkUNWjpDrvYkngrXWTC31N8EPNzQ9BoI6IArL9HForJ6UG
2R280YPGqFTOHkhJYrns9zPSw7+SYbAz63s+mJu9iZehGQDz/N9HKixtVgSkeTOt
ynCuUHFARXy6E8M1xvYx/LtXO9+gNXmyAJYi7HOKs8V0xTofZ4QaHh+Vn7u5Hbkp
HMiaHTA7bM3TDtWa4ahpYr7kGHtMHmhWFn/2M+XIM2nMvfKmX1IGYgBNMNxEDA3v
bkX3EjoCuEpzL+aoKtH5BK+IoNSsdslaZExwzQH3KCtVrPVsSOQfOgOzDKPYqY9x
3v5ySpAvU5IbfQqQmrNcqt23pWtNji8NuuAtgz46PMwwZzoxpbbKm4Z5VlvJcxR0
qru3vh7QwDWL7g1RiAoCEKMap403Fp1WenSSOA2U+kiXEOADMKQzeAqrI1pOnGog
8VLgrC4OpKaU2L5DUZnYH3C72f6+JCYO2eMeyVvHZ6rFJj8F/rCYNLMh46N+Ysjs
NiFSBIeAFVnGCAReG/GtbtU/ZZhtLrwn2nYBLJHKsE4clCg415usa2/mqtbies49
BnR1w4EHbIPoJacaXO08ovXJzWW0QBGBCBkRsbfZ2mW3SVvUL7LChKhs4c0xoW4/
CcjAJTwqM4nSs60GbICi58KPDkr8LPtcXgjGhAz3Ni+tK9hXSC6tbO43YEDAqdcM
E1OnpJHJDICspURfpmWlgskvYhU/3ltcLr+ED03mwkGgq9l8u7sat1yqQfuNBknw
XZGz4ODP9fGUqVZfaC/As+0JpOddvXiAX1Ya1jup3oxnJsN7VVWk6T2qIoA2f0UI
jA5OrMJO74r0AS6pUI847wIxWlTquf8sYzQJiFBj/ebcT6n+3I0zCCOopKtFcXLg
t8ZMKtcsJmW8c3FufzSFfA7RKBvHWa0W1HQU9s7bQdERkWx249rGF/gYlFG2+G0X
nJqoOEs7RKvQS/IcBJgygx7OC3OWA5EgfIpTTUvjSVmZ+ngHuXvlH8vTUl1rXqP6
lsvuPhdSpMr8nHO3iQqRYj8trq2xu9HfB5TWfroq+8XDlyL6+gJSQXr2BlLewMH+
ei/1os9mHbMpWkkAWIeistmesp4CqHq+lS2wLGHCRomsYyuKe1zlNSwnzX8jPw0P
EhzKsjAMCAEGXmz8f5OSHFFRY/AZtYAaKulGjl4+FZoYv89TEUVIiMQgrmxwj9oA
mqSRhI8v2iwRaHum5beUCPRSHAikzS2kiGg6PJ6gpagbdk2qKOAaOXF4v0bUDL06
fi9MNIGqgon5+/tTzsQzZN+PnGbJbJX7UgnO+yIF84ighaQezwqKs0mvRTGh91zG
qIHpq2vFF3VcehUzK3Tdq1M3LWzqMIWwQxJbTM0K9oqUPyJT5uN4ouaKBNzdyDca
1/t7SehhADHz6ww4oTRyrIrpY0n8fgkt/NDfe/IhAGLQDK9DUjBzSNf1086LVdCv
QLWPoPmpJyxArdB0BKWBmRRifKg7poPdYyeJp+9fqnzQC8rW7zAZPzmRJmQ5hQyW
jKqAf09iogetsy3h96JX/h7ceqqEd7d5vO/G/ffwmb25XtaufUklQaF9EMOgUAVV
mQvqTJZiTgpZq4PJcRUiMB+a7Oik+M5+5LxZt7OiH0oaL9714lc9HIx3QhJuYS81
p6tp/bvVfsQ6WxmgCBcUOy2kZuWIPTb1lpPLfRHMKN2CRwvxFG0KSYi6ZcH8iheR
XPq6hwWD/EFhruk6BS5Fk4DxId1eqeO/gGO3EkSkB3ZAHo93YXBubMDt8udbXiOS
Y9pFDXj9NS738EhC42ta9gtH+QM25gD94IfmkgFetdqLia+FWI6IQylSzTFCFnnM
VVb32kkc/JEelz7aFZXF6UwHbkwYcPehgGZ38ikR9/JWUmYQIxd5LIOZ2Ths1OZF
wRegGsw+ijhwjLQfJLtqZPzYmRxw5A5LLXIpYvkMjwF8kcCdXxDoydWaAD9LTkaW
OiJCLMRHb3JkNYK/+HVbT+dXWBQAr6tZfz5pS5wTF3uNl45AGRdfC3JGkYSDjrtQ
8o6vbeaDghQ354RU5XEnfZBCI8fUyLQG13J7Fqwn/SYPcHA0n6snO2c0bbRTOsH9
cCrMyLBx3soGkbTMyn/qou6j9/YrL7zgPA3N2CHw0gviRnrptojfOKUeBobD7310
6qNQAHHFulOXJKNHanajSwBeLWJs2wtRjRSmlDMa4wceP//z0f6NA0GtESho1mEw
tOBCB3CPqN3qaDijYYHraLG6JslkdID16yCCVMiTLaWP5RA5kcvGW5K/TQGT7emc
tihcJAj/W5uvau21D1fb9H6ruCJhM47u10iJPSjTKTANGq6gnpquAG/Uvw08Mu58
+2XL/WrotIVC3nMT48OExUPlLhPbdlUtdPMmgONv0rikDmccEQ/jqixOTv3SXKkn
6CHsNUlW6klyazpwA0vdPhzbxzxapPAsnSV1v1CsBAwEzvp9JXwgppz6pvjW8R5C
Ua5D6/KV7IXVpW9cgNZ9iWNZRW61h2KSPEvvUzRY39ImOnwI3uJZaMgsg6JndnBp
CKKnxIQ3be6AfgIpiEViFRCsmXW4u6DsEraYDxtgdLryW6Swl+WmpR5NCyIwD4nt
vtaulIp19N2qNzxroDLP4rhuePvdlqpEtoc747NJwEIYp+Ig78I8RPsF9aIVUxWi
5mLrkU1fHkVXL0WjTOqFHeSjK2x2DlvavA45iicOH0TmD2hG2k3JB66uYQFH6Mil
m1B3eJXfvS8aeVY9R4I91u90xuPW3BsZc24Jo3kw1B0J5/R/wHvi5eF1JDL/+q3X
q5b3AiBzYGRJrhQJPt+PkeovOjxk8K2by8PMPGf50ULXzJbYfPPcvN84NHBAD9dE
7gU0svYHuBcfLndd8OVQs55CUrBgOisZLv2kLN8vCjGCy78/zHZrwbfzrCtjX9yN
ExUeNZSJ/Ai93LL8azC9tpaTzyvEZCrsD+zOLUHlr7DFo//c/Hs/q54B6qK+s/aJ
MaWuS1pw3qmKbxAqvKkjmR7fAuI0tsYeP735HbeZc7hy8WJzvp05Jhf9FtoM6fXK
khSmFZrZvj69pBrx//CEEq2qWGh1Pto8kXS9VmCFeIUhv91oQXFYiALvBjveSgZL
lIp6DVMW9riEPQrsYVSPhf3fIWO2Yr3IVtiI7/2ZTPo6//m1+wqQ2JcxuwnUmeI1
HuMZOTcodLmFhIx66S6anJ4kspHthsYsX5gxML6YgtGXtqQqTTJcm1YPAIWCBpbI
cGzDM9mLQR1qubtH4UINTT4SUOwP3hpDfEnIEWgJyh8cwXHMOp5uY7qJvz7+40si
cXyE/N7b6y/Hy9kcuw/SKZ70NpspdJ5cgxQxlmNn7Gye6R3o9HgMyg2RrARY8r9r
UJKRmgoDvC2N0ovTu4NOOV4GHDcNIZbkLDCJbilGo6jwOA51k2QHD7btFLBng6OS
VXsEuc4YIWei0Lh1vQchY/VezVHnoEu69bs/dVwwBCKpjOCf27oON+gsy0KVxlBE
w5Q6mpE2fETcz1roR3GzdIXKhGRHD+gvCKn5Nfo+GYmycsnV98r0pl4B/4SMS6N5
N3mj0ZDKeuxqJ52zLN1L6HYnVrqPQy7HBb9IMvD9f1xJXoj/EZ0elRxh29MFOJxr
dFncmJQ3Tu79hyv4Cg23dk4AN79u9GggppALBXDBJowSoXrE4kLlL39aIro576y4
/e2JSgjNV66Swl1D7I7lp1xXeEPfpjSJrk/VtWovsqMTTdG2m9R8ikzI620FI2+1
SkqZ/r/afNQn1o0KUwefJQP6TOM08P3KivPBuMvhgATeXWwB/OUibfUad+7OkaZB
kj9evJ7QD/fjsuvxntFwSHei7CKsczsjZo8IrkjvtEs9eSOqQAWTcYlkancaoAuV
gMyTw9sHo+qzRm44z0PWiwv7sgi4488GtWeoUrZf1EkYiEeUKYgTJfsBa1F3zuN5
eIfP19vKyUd1s/Z0vL/jcEzd3bBY9TTS2d4mWKh5u1860oq1HtssvqsYMIU4GR8h
hqmRlA7YwyU+0c+FsXJUcjqwnnIECoOYihJ0POYd8wRkh1a4zUYabaxpvIZTJAVu
1vF51qp/IKzdxE/St6AZFwsGf1EmLv3Vi2KcAiRUbvNj3awfS1grKy1e5Nj+o7vz
9dUZle3G7En+E+zQk62S+DMnkb0xnlpl+ZRHt8yZTRa4l0n4SGa42Z7IsD8DIvGE
/sTFEmCoLpXU4xzWVww4KDjJrly54jg4RAqOppi+z30UsMTtOXdej+YvU8emuGbX
KlC4tCbWLN8fYwo1+8l4HSxtJwyr2Pj2SP3y/+Le25fzb4eXREScCvijWi1K4ONG
0cGqFOewdBaLqGvvuO4hQS89/yAAjoZRsixZOsbSG3/QcPcsZxIbDWTFgysemtDz
vTAgVHINKRCcmN5VO93Qa8Z4+kpo/VvfKdKsbEoFiUFoYeClCdwm3Yt/oNlD1eO7
2R0NHdpmG3kpOVS1mdb2+J+BDtchiYjDnChMS2mhuwJHfp2YSPfG5w8kcvPaky4F
wd/N3ay0IOtHn8jT1VMFpsu8UaqK0Xx56EYeDN/jGBIrAUacuQZvUb1h3Bs2Orea
zhprMv8u3Z5n6A7mx+6+Hyt6jlGeSjZ9PVcP+jcIKawg8sc/ON5OUj9uQ8UpGEX1
udTifl33POvrMa01ugoNcHjlVcf9CSfIqeYlLWU27zcy1i2AfsQmpqWkSGeOChzY
C/ZszVSN+rqseWVussaCK0WDtcAaBnP2UEQt+lJi1LiJWln0+rTaB1Phx3gqjgKs
hYSum+tPXESfRwiTwDPiorZL99ppEOoCc+m3gv29VqykDgLzf7UBLiO6hyLa3UVb
HZQJjq1s1b5ciy9GY248Tk2Oiicj78WeTsJA7jI6fDYnfqtC4zpsoCvm2K0qGYJc
F/qzlEOnLugLrav4V24LeF7vf6gyvCeLzqeYf8Pj8Q/DmLMql5yxV1iTpNX/Cpwa
tHdztUdjv0HZPCOLsHTe4XXLPP7+PTigGicUb//I/ZKt7S5T9Jx91EHAOSWCjq8B
7WfVVADn80N7IZJRdSaU6+Zoa60DMHosjuNV3mzSL3kPUm7aFdQDwMTE6W8601jD
6k+JHy82ZgRsbMwzLGcHiBsT1Ny0ArM7Ip22+GkH1IoBnglzBj+Uky0kkPiFR+Xq
eoS05pSlzGjV35xUruipFbyA4IvQFMWX005Ke6WeCzVK91GufQobJMZfKH75Upm+
FVRHz7hMNR7Fh2pfXZTNzxOASQ6lGDadWuFDBf1xMqSO6IU2um1Rj+HBkDG1wxSm
5KqsOmEBdDGPagNO4qE9EPEfnuuil50C1AHU0CNPyhTdTCfrlWjoRAQPzSNhqT60
cCrKUiWUynEbMKOw1EKOu4gxnG8rKG6YAJi5UZHhSHmDzkddDFmawgPC8rucsy2w
pfYTWeeou12DzVBFoRzqkO6hsfJ/eOp+gud4kyaUGgK+ZxnvdPgtci21F7V0LehC
fpNZDvpu/MmIY5gqzQ7wiw+/AFtz14EPwxdOiSgkidpTNs4dKljKDyPzHz1GbPvu
aiB9IPq+wIeHNn/3/taT7oxWxG+dFC0QV8RI2W+dlnTmSldDBvySSIcvfu3G5mE0
ZVWr2Dob69LQJM8OFdQqi0+Jrv8tysvNATGh7cIcB1yyiX9Wgy4oqiEcIXdS1FJB
fSIwlG/aVSfM9CykBIfxBaClYw/s5Wsi2sqAIqTgtILgYtvwT3qXk4vUxbWReTfy
xlo6wEtfv5x+OlfpyVNBjuNuL5mp+Si1A0nMBfTbLRNf20cHbKPPvLe06RQe1XlV
w6LOcS0it07z9Wj/aeM0PEdusvGOC9GJYOUQ4HDt9OMvv50DsUqE4vVqdRseOtpZ
CGu3r9dhbT/beLXGnBR04K6CCHNRht+3XPsYLKbEkAHRRUBPrRQy0Mfj9/1hv6V1
Rqr95f4bogvMLDfIQPdCnen6EUXZdTdCPq90ow65sWO1wa+0wtdPkW9VYW1GLkc/
v/oLcuWcFAn82hqgkp6CEU8jbs1j0PN5vy1MBYk/hBvngKrEOmmB4BN6/01hHO6e
K8gb7/iDnucV903QNPx5aw==
`protect END_PROTECTED
