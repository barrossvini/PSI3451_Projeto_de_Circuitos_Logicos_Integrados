`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypoKbuipa9Vjd3bQPH7Nq2Pk4ShsT4LkH9XZn3/x7BVGbQzY6kDKS8WmP+0LGhqQ
K5PW56iMuiB+3iSD5Kw3cKXPpjCX1nAA9vPQqs6OD6lI5hDlaH2VI3OorOIr2qad
jfHlx7JUuF/H4dIR0vwuXPtdMtB76px6HJWMjXVeDgl4hdKbMKfhBRrJkU0IopIb
iqsSCAxYVG52ed7/Cl888GcB4R5X6PIQeaTM/L4TugXiKeYuZN+rcnWmaO/00tJz
H8C+wGGTITqS02WXLPsNdj3nmFoiCBj/vAsfaymrXSBvqKt2kcU+8y+SDPboFkAX
L9GTxYEP5wc/3asNwjNAwwtIeOj3Jj2ke5bizmA5mdIsNQcU0EYmZjErFvmgbFUD
w1v0hvJwHl8c35/Wdz+kudfPTQiY54ZFo+/gFtFCG2e7EsqUltPjlbhqP5onxMH1
P4URmIae7/f7E1TVqsKX1OP+VbUoGKVY7cw7S4G8txoUCblLLIwgvVoZm9fqYPCr
5R34rhPs2jCGZiDsCy7LaqqZ8Wc+20ZzN5ak+MlNYZA+kKW+1RzaZziVfVc9hWsH
v7tCyYe2FpHkkHlZ+Mj86iPwVT2+MidOhdxB59aHUvq5/X/jIDPuQq24igeiPBsn
nGZXXibV5ZEeXYgtZxgWA7f+ztDwQ0TsRY6+o8KuIN3dl9uiVs7uwP2kZ+5QFQZ+
WGSYHJ3ck90ODRKnt/9rsjROe4al+jd1RS7DOSnhxktllH6SrmHqH8YLd/yBFlOJ
Lo4c5wyz6vGcsUoFRe9puNrIs0H7METGP3ULh8SL5MSAYbQrpAj4KuwuIJEQ/p0+
Oe63yd9+XLczBYa+j7UL4u8eGSy2coopmGxa4Pkt5fVE5r7nWKqtjwoHXNCZm0ZH
pVehl6Rwauts+JWNWcs01t/3dW2tOsSMGh8ky6N+tdT9XaVcK6Vr0rsUc4AlraqF
9WAKVJNk9rNj2efxQSNLBttwMFZuKSLsALnlvcAnVIH0gxL21sAXJwx2wYGekmYx
tkNpVPo5yLrI0xdi3Zru6rYu3JssuCOzUTh39fFYQeH3bORKwbGUDvKgRsixZZIZ
b35Z5gG7pQlgrcDUGSsDYDX0b7w0uCqyYsRrBJGjw3nzADJ6fj2aQtbjuUL52EoK
lvxeVT7hfXz+tJbHeHv7fqIf60hRd9NEueMVFRhLQs6W4CBptIxwfVynD2nFml9x
xLJhqtxCtsMcbsF5WdTERdB7Jp/l2ZeZHwO4iiqiSI79DqjO0XatOMoaSBGjYny4
D27xgMLd8j9ebLmSiDg0ENN0RFeMAZvxZmngX1/r4uUNNpGVe+a75jYTX1ulybAl
UY5cqNjlorhyH2YnNMXFiiMmSTc2+anivy5n7vX68v1FxZJuqwEi7ykBC7ifO9se
SwN23hSRizzb+8xhHI/J4IJVCIBworWBdkYqHuOOaziP3AS3yMPT0S/OEnJFVxWf
`protect END_PROTECTED
