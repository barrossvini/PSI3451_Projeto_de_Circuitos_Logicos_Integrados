`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sy4NAYXvOgvAu1KB6rrne8nvDcg4ukaQYu0m7JTdfyNDFY4CpxHT7D/rxs5crqix
nXv+GwuaPfrKMDZAAs5ors+Yx/NYCzcObC4kAq5TE90JdyqizRXawof8Zvr2lN3B
kCoPs59ePi+8JhtM1Blj98QigoCMUQldIYzz7oGUDUXqBw7qwDliyA+o7gfcVrTR
l00ksqaT6kRamckSy2IjY4wXDdTY05VcvJmxchP6g+9z9aX644OjRsmDLWGrWZaK
YqhfavnzJMguQPTFmms7tgWiPlfBph42ndRlVU8CqpCzQXE1igqDaZKUVoXQuc+y
ghEYhS1l1VrwDoA6kzo5Kk3UR/wt26YlO12GxQ1QbLmVfDGofvM+qyIkPbJAwd3G
PI+uea3HSM6zoRvgX8/jcPyaWRlIFMAyXAhQRszICT8zcSIrqKEGPH0lzJcI4Lh8
km/7ZRC7dDNdQBdep2us0xIDz22lSpAC3l0FtFNUiwm6EZSz58Z50WBOucV32hNd
Omu9C7p2rdfvXeX6KfxoNx9nHrcLiCParDzghZyQNno7rRueVYavbPeBdQA1TR4a
1rMbG4H1VbNCWBjWk0HfMh5NY+SV4r/u8hbxlGqbXM5g4/EBnd8fGYhrmBDPzpat
V4j8+ZmbWyxlQUfMArSeMvy99skLQ6C0y8VYIWXJ3T2ObnUZtJZbxEnbuRD10QK5
dsm/7NWrvw6/nIx1CnO/nImu6wGbsnWDFhdad3Q3aiUqNt3dOSppNch33VBQ051J
RPS0T+e4yyptL1pjwjxDpBCHlPACbmx9IO4tm/SzmaYM9U4KTA3b3Qm4RuUpzqN6
tw/VjZENCVx9Saj+8sdJXb11StegrlOSfTz5S3QZHCUNxyBiM36lE9VI1v+l/cnE
s528Ua9CXdjQCaMAZ0nK5c5CvEWGwW7lp+wGBN1zOyT8anWV5hyocw0e4JyhNP1I
DgbQvw7K+mXKtPNmrkMmIw/zTLbecFlHeoQyhnUEwysPeLXYxBmdtJr3SKPvHfAX
ckbTwour1xG3sc8yc/UGG3Gm3nvwTFBtPks6RzSjuWnOzpZpC/01gPtRUsi9PuJg
YnCe3wZqbMXBiQ5ugt7Sk8OEPDVMH7tqCkXxquf6wTQ=
`protect END_PROTECTED
