`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4VmREh+pCcGIJmlj18TUX9Ie/ybLQqhzKboJKrWhhGHbuMknfoxf3MFxk1Qz2hZ
QkqRfyE3ntKrFHHaa5/cNfeCtiTqVLKFmtgzpdsCumsPjQA6BG0qFh8DDEhRUFiJ
ti8giWzep8oeDiJIc+bFCsP6TmjSN4JKgt23GaAhAHRyqiwRa3J1OrUtdtAUlQOH
mviTVi/gm9BGMHVVtu5swW2x4zrE/sl4COeTg6fQpAhkRDeI81Gg09QFV0bA2VyT
cgYESo3qiUqrb3/2ekbZNOWPcpcoK5OgWY9X0aT1R35RSBjvAM9D29S7pXBEw8JT
I6balxg7p2NW7JiWDPuotvLj/hqj2saC4U28uk3g8/xa2Se2MrTGJMkeUYAzynyQ
4CTYvjgo8Xqr19au6pE9X5Fatl8di71tv3Yz8VH8PXds69quAc9dBPJnUeIRy5jL
B6QeDqpXhJ479Oy8bsQHiOR+1sBZxEl0fH32Ju9v7X7YkMc1At/sn3nNaXdIIQez
L+y00nUq/HsXh0lMmW44Qczz+ZiRoaRC910TXvXSJ9leMtIQZXAdrTYztN6Pq7HK
+HmYwMyOa9127awFYe5AAqiRwc1dbmj8TALHCUMFN9fmA/D3AYpihgYRbaSdm7Cg
XD7KD6yTCAuCkCN3OVLKM+8CyYlv2aZ6F0w5bTa7gqDvnlrNoFKI7EzjQsC87qM0
+aAAkZJDwPYqd9X0BcxHD4Yt6f6jA8BUGR8x7z3yBEmtwsLqFEQMtgnafF77RdEH
U2s7KjBDQdmKUdBm+mLQnND3scjsn0KS1CrcGKG28+Eqio2mLPixJnjPRbWWuzn3
L+GZ/cR7TX7czUjhQqTVBqzqcrV8Y/Xfb5bFFvV/3k9H5nQ4Ghhx8Dlo9d024CqJ
IoAk94kCPBA3JbNxF4jYrWbTG/WFzAprdefwcA6SLQOBBB5VkKbrvnOUtywuldGs
M39VmXOUw8OE/Hjynd4CwnmPjdIjvJMbcliIeI9mfsRlQNQlRIMToHSWZBLU5VUs
0gl5XVGgHQJRz+fGOrbLOOSE4txQBsho1Z5L2+VGJsCXsdMDYKU44JQ5oi/XcinZ
eXwYrYUubdvFZx42x4bcAFEKRDS4t8FtT4J7ElSIqkTeeyfJ+jJAW/+TK7PdFqIL
50ZkZANxBV7pwjO6hr+LUTWkMkg8jn1xIvb6XfENCPGeQYcBSTBb+83HFZteiOfa
gFtN+Oc77Hl64fhSC8jkegFdl9wkdgaNn2cFA6f302mdJxXFTsmWtPdD/3Ml7kft
lWKT65qxrHFtCrr2bLsZrkOPVQT2YuOnVqmZYmBAww1wLKVKO4TVxsz1E4Hwghvp
ySdoQXYy2/kHLLIkKAUYdygKr74PkgDJyws6ilqQUjQNLFfzFtWbHOrpxn7pcFTx
UBNgzz9rBCd3X+rlERvDOFB6UCqHplLcJ3isAYyoLL8AJOr+62kqLKpIn9x6233t
zwdoYzMVbUDRgv73Mpv4vOzb99pM55a5rVXSSlSFv2neoWOC9rsIjQqWD3cVADH3
29eujzi4rkUdbGAZj33/YTW7/9cspuwgcFUpwrNJy58YNar9GXNBI0p2PMgteSBN
LlpZSPQ1xfNWlHRNpiX7ZtXI4v/i6Zab0Ds0DAf/4AosUt5suM3m/MSpC0tOxhd6
6rsvjU6co/6KBEfd9JvIi/cChYMGEwxnL3RGguncvVgnitir4PIdqzWJz47kzm0d
FTcSnm027Xin6sRFlFrzC741sGq0mxcxIdxOERlm1Ca93nnQnOWOHJ8FtWI9BEgV
Uwl812R59lNxHD+MZ2bSq3FmINmS0dmj8fgxN1o6fDkFiwlfrrjXf/1DiGGIzRa0
pDFnz6UGXOxqhupCvIpmU5b/lTJNB3oCXJFTpcjKKwL78qPA5i6aAk6KFmW7IJHW
EfH/2ro6MTiw81jl5QneIB6StVqtC59fsYt7SM/LiZUJpxwfj1DGOj/+1nnNgaJQ
Hs1u8di6WnBr1tet1guDp7GUTn6jCpXzSKsPj8gGIFDiqgNn0s1Rw0iiYwn+yBeJ
v3vLXiRSqQY9PNCwBe2yCGGUHzLPdm9+xW9nxYBszFW4PZo87jUygIiSX+9LwloX
/gKEBiZbC6W+ksWfY2t3NtDh7iiV/3PrxLO9xCHwCXNEy845ZgrlHOvZniikvjF2
rwEeMRR1fCJ64VD+0aTzwK/LzsEMjBgv9S7u3B7EUuoS+LPfTfj5n0V0BrkKkbp/
DfD7bZZQ1ZUcXe3pSNRRkdfnDIpYfWzdEViYeIgxKzPlsGISXbUG2x3hFFr2+9QV
qZxepfzPas6NeZOzqckC2n+5SqeeV+pfEGBhKMJCbKB0b/NjA0/O+uHFho/lc4vh
Ib89VRx6LlgRxWRewbXOlboGFFrCcmRY8ygyfZasyZ1rmILLJTj5w/6SohvjEHps
LvRHIHMtU82RP4WJ4CtErSHrFkG/82T0bBRrV5zX04mZVjD5RcqK1OVx2T0OPw2g
zV1rIMsSB7Ww+nbkcHyA+CHb0WYI3DtaX1jrS2DVa/9zOPltedXYWSZMSzTUgQSi
wsUEt2J8Id3N4ianpqcWryjHLDRHgKEBY4uKhOU490BsaKebIk6yMD0Zjd+25ZyH
A7ZtO9h0HERp0220natfoopDsYMdAfgD3817Ymq70ESS428hTG83rj3zS/knZjr3
aDdFGC1KyYvFs1yDRzJ+5iyGa7DxuMu36K5E8rt+ZkfaA0YWHrQmLpUTc3kpMCsO
EPTkq9QOWS4JYU0a/b1Zln2iPbu+ER/nXJMC5dNYVWC/VkJLz0b2hVAlUXehcSuh
aWC9MtLb47uSK68kmggf0JAIh6fnM1uPdtjeX2uyYoBjYigUdUVkWr+DgGY5nOBV
O6MiFPJsYRprBjBfQmMJ5gzK/R6Ylk9QOePHHkOcXvzygiJeerAl9Oz6zQBts0Fr
nuxBXL4dw7OpGWrzaJo3GW/AGmkj0mUYzX+gcPSyR8zwzFgjTrAetSxNyeCgRKNu
9zngkgOAlTVjryHYHl1rpwSiVYHgtcygGoW46L63bTER8G1DwjaYYwqHFn224mrM
Y+mswgvdBMjpIm3GRzdWujaAWhqXES8IGtJD4TfQSRFLKMqWO39woHUzxBGSHDJ+
iv6yCjcJ37FEr/B+E6s0/hU12Xn0rIapZJ4xx7KDPZf/CtE6O71EmbOx0sk9obdR
Vz5OFILtEP1zxRysiCLQGznADmt4u7rYjkSMA88Gb3PXL6aRpbBYE/P+iEnNpOcC
SMOoVjZFmA13H1zB+hSbyJQMFPJb2+DrXlBK5jVsTuf0hIMoYdief06cWHhBlMiJ
TbIsUbcRBdX4r5wnKGI32vGfM0IZKCSUgoHlKFPwQ3HSRGv6Zs0am4Hi3Xs1PCph
fMhVrSeHgqyD+gBuxPppTqSprMiCvzs/XfpWCWz/EUCPc18dE5JKsT8khXGo2z2s
LrVDAo/t2ti5r0mk82Q5zxies/qCWtOym4sp152iHKMd3rcOZM47EIH0Q1bByNSS
qKOUNQZgumcHZBf/LKWVf8GVOqk3RClt523lTBBHtmjHDJrNPyDwllTc7XnIGagJ
SFvyhfz2d6xBNWuEDBF1vEk3C5tXb2J2rF55yobmFFiNBupV7nqXG1UDNGKHQGk5
TSCUqrlEvhbirURcRGCDfSIye+36haW7kcttQb3AjTgaPX2Sj2g7V0qiFnGIelN8
7WOhbeLQGvLH5fLYLgMvEIupCMgY6rPIuX899FKurGKE7+LzG4IAX5xuCHJJgj8U
RpJH3OD/2pHH8jk3QjkRsB6d/C35Czo5E8XnpIN6QXvV8Hf4KCAPHCkgbQJ8NPvj
Azw1Lj5wCx4d/nkMfpL1Z04fqjgnM59MCCXW6XjyDsRqHMg50Qe+ISYpm2Mg7sTA
vfiSOs3ZHzYRby8o0Z72HA8pyO0rvOVYZTWkZCkuIEvssrT+q522/8qcux54vl6F
xsscdmKsoPRVHyJWnNvDLtI6V/oNvpEsYUQYFTtHAHwa17BgaRReO222DWpdqznF
MyIE2IXl24YKiiTmSA2RWuuha4aF/nlJVZp2Enyu0Y6A2M1x67JBx2ovzsAePoZa
tQ623Y52jZW5y+qWE0Ci4pMiwbQyD1byznGMik9IQEa7jjg+nSrNbDZu6YBcEEYh
X/kdsGC1LV7qehOqTV7hQ82zU/rWHDARnIL09K4oOojfkbaq+aKQNUw8MF9EfTBX
+i/oBetsIdw1oC7XxvwRuzJSjn4sDykOKnbXdXA5m7CpnVVQcbnMK+yy9m9XTyB5
9VV485KTAahRCm0N1lAmsztqnmUE1Xak6dLGRAQyruZ4VwYm0HH2U9pg7LmDfwAA
OYZtbIty64eFp68caREiOSOEKOE3craA9szfNQnWS/c71NBe665T07+PO5szxh6/
rqNufnCXhfPJMgfqKCTHZkgHYqviKQXw9TOJSxClVvWsCDCEw1gA4lWztANkNHlC
7cYyjfnaRWxLyoGEKRcezDRyEs5m8hTXbONDmEUK0xADpdPzUwNatm0gywBekMBV
XM0cUqEYOZguePcuNIbF91Xp/JDE32MgjJrah4awWD+i2KJEIEnkloWLnArP/NSt
EBe15yg0aMjEbhYNmHQ4EkItE5AHB4tib8TPlVjGX0WOdJk4Czq0Qu+DQFDlRh/0
HwcewaqGvT+D72T2USKQnupHAbyxY9v8kdoSyHMoJX7O1sfr1IPNe+PFzU3eUEDu
DvaQUFNZSsxG3eIc+4qO9j3yCdoDEdzVLlsrT9SkYc14kKdsNEkLae/8Y1zdKWlN
LJ3uftPGssQqMo44Y7aisYlVVeikfDgcgz6MYjXp7W2HB0ItMPuOoo6wzmt1jUeN
eTZXWDzYT6MhYLpmjx2dTbg/7TiqNPICJorklX65lK36ywuxDUec0gjvqUgCJYNo
JoFA0+MaQmKToeGuXTeEuAVJU09/hK8LB4XZkanC/SO9SfH0jQKJeRrIyQ8jGgiL
ewb1rY6x/d/eGIfPH6KpUtXOL/A71Fu6vbbzXlrualseqp5vgZJCqyX7BRptZ6ln
bfkLjizqyNc7nf8zmqD1kjjIl7Ne3GV3Ze5/eJeUGdeRxnkVAc9bA4nAXkPatj58
xUkNd2k/nPoVx1G3/ptWtVxbm9TNtyGVlwMt8h4IRGR77NIjXvie1aDgWXsiVCzb
rtVGCXV+6pAN+Ab5fskPSjIUHwzKni9nwmI7dsMemkOwdTzYl4Iek/qnsEi5rxgG
CJLzLFKOfCWiay6RcWCxaaOhlJIajbQz0p++znsUTruBcpY+9Igo0GGAMJVIEAwb
RPggy/Ub4TDQHVMY28rm9Ezgg7f5Zao1dsNiDLJe3aa71G5+NsEXQPUB/ZEcvIqt
G9twaylVPzuseOBerqPTiYigCKKa83+89xHZNLgGICxBCfTvgN3urNeJaW4xSYLU
IyYyCtN7TtG32TmZNsd1MUE0qHTKJM4TAy9WWgdosJh9lRjk7RvtTFYu6benzM0i
ChrVWRAxQ4IBlRFCva++YTw97U2H4MQ7VfCSWmDA3WXoBPdAgeIVzd0kacJWcdrD
ulKhex+nEgtzUMDY4bgF6OegIwGXx+paRQQnjYk5djFqhqXhNT/HiwOMEjsFR5PO
OhIdV4IC8h4zKoJwfX7tmme8ufrGdZ7AJmoQAuJEPEHNKdY2+NxAl0wzLTncxVog
2ZFErBSKUP0ZseReP3jrbQPahPG8jvsDobW55ifvLEYWzs1UBmTJpC2HTQRmmUgQ
DIrQOuTbvNoheOm5E3AwYqfe2hazWS9ew2/pTp9fgILm4Z2v7vS8vA9QTNxFSVAh
WXyxZpp1RGoZ1AViZIfvxfRl/A5gA1SPjg+lW3rq/4L14/fs2vI7Pfr+oMCyxjja
IDMWVGDGz+yMJ1ZOjetXk4Q0vXhc0rLpWDVUvD9nM/bJQWWYJYRY8yu8ex016HOn
eXP+6jVfAYMFkcdjtbuNn7qs9qSbc9oDAffZhwXWw88RTUGumeFjndWwvdGTkcCk
FhktbMOj+9klD5fx0f6f4TNLwbqgFdzNlhrqBzX1v19Qd1gryXtKyG2QqTa29dx0
VJpPdH5mkXHBbwmRi9QXC7KixfPWck79lcmjY+Tvgq+KCZrjAQLoonhguFMU8lyC
X1iwS8MXfa74AdLGghe2DtDaNlXZSZn3DFx3m/QOHT5woa0cGtfPIvBnuYLn/n9i
VSx3y1WZmNjVUsQdTGKGc9U2jS5N++3GEK1JzDHSXryRO2/FDmWrisrxWISo0dPj
IESb83v0bJTxrqhEWYigkREQxSJBr9s4ADE12NyuOsnUItS6ML5GSQX7gU3B97qF
/PNZuNUSuUw6r3Xfl0pOGRlTlIgCBJV6RhElSkz9WZ0nHVmrjGdevYDak8rlviSV
pNWO7CHGPexH1pEOLy7ZmdRfsMZd1xnLPqJOtmk/Dnli6w3LZ5nGuMcE+AWQ+m1t
AS/XlgJ0zBAgBbw3w8csWPWSOxMzblqpykf1nPHmG4BWzbDPJ1gb/lUgwAqIflDE
xNzE9O2uiLOGVdr7wW2Hgrow5GU1kPiF0mctYMvMxQowUa4Dsr/2wf5QVza9qeGa
//BuH6i2GU+XGC07Ali+TogbFXMW/mTsTfWAxklxCBpe/U0wCQtqrnouNm+cRHbX
5O4+SuaOCYYrUlytgFS9y8IY54EpGSD/W6/fSElTkU+CPpMHx+6KPQJ9RROu50fo
nql/7cISoC6cU0yhLNjp376iwyHiuBUGilA3Jc76twQID28D0bRpBKbLt7Fqm0SF
r0DWMkVFl3k51Nq5Bh63WbYfJChFToe6AGmbRTZIGtAxk9ti/4QnszBwRE93FN9n
O+5EKiWDHrldhgTvBdZTBdqmBRWc0BtlPBAvP2OFIn+BbU0jMdgisC+iR1DqUhxY
g5759JAHrTbqDHNXMkjNUMJFI3f/5q8eohpY1v+jATTciIcrCY5MvRlZ3Nye+QEG
l+V38cgjt7E+nIUfthZFIbT6se61PXcaU+/YsIRDhnMUL1eWeDxbHwGpeKiP27tc
/Kvtz6//QoKV21xwe5UXfJIYRNfnaHjExP99xOCZNvXsWA3Qiep/Muh46MgM77s1
ngMkEppB1DCDxp3ZQ44DJHIebt3NFa2vCUt9UKMacdovZWbgqFk/x+zYkTaHW1LH
fBNMB7SlJEKBx9UVwlNia8aYykB0jQcuZHQ/8scCvvDZCPiNe/oz28flM01M46AH
ziMMrPMN4+sZAxgF+4Z5J3sypUOOo2utkCQoU7oyKuGY0LDbzgGhGmuUajWQ8u8a
DhCaYU7CeerQng9gxPBd2A5Qw8elAjd3wJ8cBeCqdyFXAFaAUglK6YjbIAYp3vHZ
3qn1QmII9bHT5Xny5rrGvMydHcSaOlvYP+lU7CSdXLZ7Qw8/3sxss+0I7BTnPcOu
7j21xAwkukkoxnJf00i6ZS9fjErE5VJcvLNYivQumhnWhEAWJjCPsxsKWqxxFMyH
7amK7OmEcxz50LK7bhFTcV55gg+t9IFILmJuTP9+noIUcnFCpBdXUZhbYl9ZKWrH
PUkPB5nee7mA+Ll10BYJ3SY56hpW8TjwgbdJaj3tqub9zHhwz15I1tOqQDfXTUy2
a3R+i+dHCOFWTG5IsQ0mWgYU2zpjT6OAxC8SsRi9wAx4QQ9LEq0nfTNOnNp1SiH0
8D+SBUeguHua2EAy0VOXj80bU88vbaSm2kpA5YlEzB1qdtixXRJCjSlXonA4LDfW
jE+XFbeyOSGTZ8u033sPf/1a91h8C5p4mbsM17TxEO2yYIPAuPUe2kmBwFNTZ5ak
Mk4oHzdFWbHnuvblWC8zHT5EtuNM7YTXF3v8Cv+vnBj09ScJ1wBzyW4HDhyprmYB
8JqBcSmjnt2rqdFFYn80n90xqZQwGnYJag/AmtZzcC2vPtCflWO6HOuyqY2XLrKD
Hdr8Rd1+jZqpvPQoYAJO0QGV/LnPrUWmlhvUrGlHEUMcczh7wHndLWlViVrPWc4Q
B7Yz1v/pUym73B2LGTIyseuBCFQglCZbIrvtKQeaOBpvcHQ06wzyqFIrEeskPDZW
+I8R5wt32nslsRd+3NsNlpVaFQ1IHIYArsGaTRb5GLOOTZqtk1gjZ4SXeFEC7wPi
vZeo/mMWVEWmAEFMaT6jhBbgg32No+bPsMJeTKQujYHbzucjOuHEJcEG2RcGyK89
YJj8nZQ///jToqoLyzqbvlWaDgbkpjNZtZ6/CuAecPq0Nt5HRiqVpUWgsx64jZF+
9cpsXKaSSRHmdQubp7TS605wepSx1BEbKcCMcFgfEYsksSDdP3JX9BOqD8MnuSwb
e1qd8toGbAL4amvDLXPiSwAFtzvuNttE84FeHsNxY5UOql0kjDHOf55+Dije32qC
LsRhYOS9luTd3Ny1pvEFqjdNmV1Fs/1jxIp2CewKVpHgQGjLBaAtwqJgZSWOlfaC
VRgyfoZP+p5USbLLPmrRkPY4uDCGFlcF0vShlvR1xFhN7gjAG4fuKuIBp1oxq9ZO
hOP/uzUKy+3kN6JHKw0p5ocu+kQMdyXhtfkyH7O16+7Ps7vxAVr1iI/LlwQzTQN1
QM8C2gBroT9ipYaqVTYa7ibZGj3TfyqAhsayQ2a88XGHzCscKvjDs2iwY4uffnF+
HDdGOAM/1Zzkq25QAdTmUT+wr6VFtYApz8kHqnFk5FzPUE3BwEc03BATRLbCAmsO
PfNNlVW0G261yv9rrw10P/8piFzXPIdPZdgFDhDegagai406fSrT8H96D0KDJBvk
y0W5Mh/TQrcXOOHNLLyM5/Y2qwMM1dGBqkfNN34wY3DfFCy4RDvfso6lf4i3cztU
Nz8KmNTlkFsL8IUQk3wAU4WCp58tzbYLoGm4hz52l5eMk30YM19/pykTZZJiiUVg
X1NNLLIyQOpdBKLgEhOv+qn1EetQM4wkPdJq0+DkaUSDQSd5X1/c2Yz7SZgxU4FB
43oSQ18uth6AhHm0GxpuPtkL5thX41jBFLm8twYjAIjgxQpirW3o46e14C9e4Okj
iPBFJPwBcaxZAqULdDB3z0IHFUJ+x0i0DQD2TWwEhGCP0oa1sq2oNkHHMfN9qnqx
ox/79MmdV8alQNlChw7aM93yI1SFZOBFKledPUN4uYcUFXAJN3JSL9x0t5bI+gaD
11ktEwK5ICZX+HofuFI7nSBpPcMbkCgOCGHT5512cNp40ntph5Uwtu0t6ruKJ1hz
bTNpZo+HtylYOwz9ctryKL4l7weC2i+Z5nnoQnAvTpfPrkXmI6CTvT0AjEuUSksn
1ENNkHSCol11VzkqEN5V3rwRUqgvNyX/+e1penowhx1mHpwgaozwOx339uOLDCIv
+98NtDURZGRd58a2PcCI6CH0XlvbZCOr9Lyxy+e6YZhDFNvmsV2FVbBXluR+hSqV
Y05hVYX6KFmWZc8qJ1wK9BhaDZOlqkJ5e99G06ni17WtsnouNWAysz6m7k0+dV78
4xj0uhtNfvDF+ozTSN9YinzbC3d5/IDFDqr6UhnxtnDaSg8j0zS0adsmIjLikMaq
VZcO9+tZf7gKyf3+ldNv+xtOGkWvNvDLCSb1tdd9deldQ39D/Fj7PnlWPRm+dvV5
KfB2+OuV0D6zWRdbqgMs+3lbBg3hRKICwdLDLzC18QdiTejgFPlX9KdD4G26T+N5
rxA1JF7o+ZyJ+ouZYC7ayasydqTEGHsvUtmm9Qrq0v8KqUw25hzy8SHJW0XIvcmR
Bxqa6rtUME5fCBNup236+DkI8JKX2j8D6DwkRecUe/FgMWuQX0JAZYDNzgbJYFCG
UXbdw1XaOIOv0oJxggsnbmv8SBoos1Vu2e/MRaa1VHPDaIyjcwS9GbCSldKVPg3+
ArSVzSjT23FSmDckqBPJwfVXTafQv8Rq1CREUMSZatGKnsueHW8x6BnEI/Q2unnJ
46nqY1Dop/U2X9Kd09YSGnSO65U4onmMFmyn36vJ7opP+QPp3sS4LDOapwGY9/St
+MGgYBGNTg2zAsDUv9n/Ka5LT7Txk5nYiHjjrsXSyX08M2JHHF+trYQMUV+ultt5
Jqx8Nbkj0Cqyhs/Wy6FQRF1/mymst8sEl4IM2uIQ2y5mb5NEWl8wwl1et6loEyzx
9roIfcDzegWqDwFOKUxBnJIHch6yrxe34manp6nEGxYSA28t+HBJ32AyhGEopnN+
bKF+gWatarw174jrUMBcsAywVQl9h++yNj4b52+gURSe7sBBrD3OQH8/F+MfGOS5
MW2O0apM3ovsc3rvizsGS69X+Wzs246SmPtaWfIfmmJNx9oKjnsF5y7rZCtHjtD/
qf7jXOEyAcmfFxi8lcV2tdMqgPYUoEZ0BA8J2GedFC36vtc+cntP8Xe4UdkSvlDa
uyuCn1Ju4e76GvQzB3xP07iGCd2QH9Od+B4PL/BquQuymWOFLmuApC6He0tFGDJp
RV9SmSov8pG4r2Bb2pvYs7oDraCw0HAVxLhfln403ZBLSEVCkEQaYBAZTnbPVPkQ
rTiSnmHxNylc2bI0c2E0Kk8ig76LFgcyikKJn1RwoKcivV/ya9wE8MZQXRIAkUFR
iCjCSfgLRNTAgdQdC6FJr8EUEDCczpOMyq1sGMn7bCTRYwgmuzI7C09lsPYfB6Gw
USbrBbdhU380imW7mTVJEjKjcUxnHsKfVSy/IjdNJ4ot3Jdi0LzwDSkEpQoVY99a
thiU1m6RvlxjANHgpItqZp25nupPNT/uToTnuNXKV75QFxlVhb6OMSWv8ND6OgoY
VKpEvK00AOiwLRJY52e+VlgYwGeOBAX0vP2xybR1AcmvN/7HduGLFAxsdgq+F8OA
Pij/jQx5WQY3kMuxGXYddVqXjsRO+YqqNdOLm56vP5YVb9wzUiLJmtVSOfNon2Wy
s/XYKMZdkJ1A5ncxlE6rozz3fA8wWzya269mrMAWRLAXNtVkMHc6DLh7IKqm2QYU
yZ/LMouXj+JyEjdSEpv6HLM44ywnciM5SSmsX/x6zEgyRdcDo+j9YzJb/v8VpHYP
hHHfOgmvUSuPXk6AbGYtwb9bcI6LNDV9TX70jwtHR9uk2AKyAXSpAKYyM7qbCgS7
sK+i97IrgYqKRdC/1PSlLonfdVMei0HUDe3ZtGq3n+5RW2z1ROarTyeiUDl19Zgv
Hblp3e0iJKdqYks7vdeGE2RE0wulILHY0JhDPLks7/gWewpb1v8/EHMTAaqDZxJs
PvFFyblV/rouNdwjk+eazpb+qoHlEb0TqOXU9qy490qxrodN8fKue1mPzPSgv4zI
HvA7vrQ5WeQ3hJWeb7jqGKLA/lfX6yiYv4Naq7853rNJeaf7nkWxcpJz2gOXy/of
fleXVQYbkr0ZthKPrO1HT0uZkKvCNuF/n55KZvM6KtJBu8UmXKCxp8n9l2weFV4U
YpaSPieK4X35O2dHMxclaFITH9y+58wlP7Svadd7/cdHqny6z0Om29zGBEzRTeqH
eDSe4lXur8k7WMugxfJR+zMzlsovpZJOkp1cVwQd+1HYIwVikxdVVBLXUMd0SrlY
DDmn+omEvhDWkdY3xsNVjusqFvW3SEeaL1Al0utKB4i2cp47g+CbmCiqJD/xz3Sp
mIw4B8Wl11ZQETT20oD4Iyj/lpLbuh6Oi3J7QctHCRxnVQRHYXTKA+B09/GuM5U1
rcW1HEdJKlb5m1pAVU+a1sYsxqtV0d+/ww01deCWjKTGsjZDFQyoEgGeU8hlWEsa
hOx/FsWQbPGk5Y5adSMIBaIbBIQ8yX+a/sQ4bYkbm+7ZPC6jLqQFtG1Y+mDyqHtl
j5MQ9vCy+skoZAK4FIj6HZBUxEzgBlKIm4BFKq4SMQktmtvAIjO5FlvUc+FgrBKG
3ADdkHzvCvYtmUp5arRkHXQ7Rf3gt11JN9GPLJLyCE5ADnEduxOWG8+iD9pwZVTL
S5rV+GDuSKLPUvfQ37Q/YfKqxED2VIqHayhG0m/gdiRbfzHvqIVUx47Cz/oDd0Wq
kzghrnItWBsAW7SoKN+6FbmhMODULe1/+At7axaMO43/PKzb8hnp1rLXNQJbWSwV
C3wyYOIxfxSBdSHM2sLmvhaRlJiEMIu5xxQHsDtXJEmNmVZd3UghokqAD0+5iFVp
x/fAsZ5pYmbJVfzxmOi03J5VqycVKH+Iyz6RxernebrB2uR3rEWvMJkwefZOZN67
mtCJj5a16i3U4TIZBAqGwS+s2oEo10Q1/qRxpjPT+MlGOUGA/nOScGqkyzsLna6i
i9IvyXwJMXdKWUzVC6/Q6NiJB9B7NQvn6nOpA8B9NsRue5W0ap86WgHrV4gOtxcI
twMc194nyjBIhgKogOJnipHU/3dv3kySStA03NEYExuAMc852vNrzXdQa0WhEE4B
JBYOUIQIHk+VTLsPXZlAkHeg73hhVVHqBB7eRCvE2Ql7Ch9QVWYiqAopC8rNx0Jw
G/ASJtyNmAUHLKnLw9Gxl7OJaER152AUgaaynQVNu7fgRrgRF9gQFnsx8+TiiSSa
XeqF9H48JSATEDx9njsHFQDD9derzezA3iA5yRsKhK/cEAdpuUUk80GXABQlY76/
H/VVqHih0ptnTMFgH8zkvl2SjBMWLyqXCWENxL9dQbMqk/Ftf8IF0TLXQV1krP67
167sJPSaK0fyOLP4imuw7EwPDb/GW9zloAb1QyGMzLKlaElfIreB/josrFub2ZZl
Xr8IsJwL3gc4abUjzUQkFC3fl1/FbJJj2XlkznIbdnYSxmogtWF+wFJb+ex+S+Zr
07UYGekI7BnAUkFWVx5podiIyTFuvf/ZpkQz4IEcl4wdSXAUFvgXKjZasmBNkaDx
alpCDSNia4Y3PSrllo/eurjphGCT2tXMc1j2/WYmclNB+qJMES5d2w7jjyU03VTm
vzk1/N8GwgxM3mQuksQ7VozGWMXoE7sD9e7jbYX9z+ADymwr/wcQDihqCchonjw5
xOIFK150CPqAT94KJIlSlO/PCfPZc2pFXP1F/hqzU0ubD1euifcALpIkqorJtFgF
z6J8aWkH+CblWGZwln5N+sKfNsv9gfkyi6kzh/e4UUNyxDugZrdMmscD6jiDjxR8
EoBpZOvwJuBsz3f009RsbA6P/C0nwkZ299xksFueY9famtB7FIAyGyh+W5CDh57K
vs4FI9QnPz141WFfgzKq/ubd3gJ2n7JoNcl5m//5olJno+8Idu1kSrSZtu382Hn0
+UHeQk0cpLzMEjOMJnmSkzLsGOt1sNAYp7hLBnMyBsdjMSWZM0QZaR1Dwx7Mvbv0
3L7BPL+XGB9hbdf0XOlcYW0xR2WulBRinM546B5s9v1D+c5jAKp2cuweRLzWQQce
r0LWSLwkwuNgxNW9Ak835A==
`protect END_PROTECTED
