`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJBi3TK170gQKJPQjpSV3ArnK/lHj13FvlRgFCw0H7Z/FKQNjlQIFKL9no2gJarN
33wdR3GpRl5Ui5vkEx0lztE1xAMJzqqAy8pJLnWtFt3GAhzKSlyWvhyO64pgVEjp
7X9iHIhxwSSSbal6MsnOAAP9ftdo/qe+Fxr6oO6ZQ9v8nts2o/y59m1S5dEaPNE/
7Qqe+5ggAJAbEkkfMhNVmG4dlNgACDWJVv2pddscgrdTC/2Xp3JGwzxQYsXlm33P
ScQdMMl8bpHc27RB/pjnuADcqNbA3KUTGkUcJv/R+SUHdN3cK5J4in35ANu1wT/q
HGMos/Kh9SrWFKGAYGX8JZXu+pEfeVAS3mwF1+ZiquVQh6+1NInTeWdxeRQo5k34
yYTQSXuzB9dD56snv9DvaG239IIMXWBpmKrWRbvH7oqg1xWRGhnPmbEoXQXl0U35
HLAVQRP5GC/b0j6RxPZf31iUAzXaDYhEzpMsplewg8Rmy/zX/mnGS/E5h30Zh/Kd
3uBhERfaDiuQrSantLVWl5wv+qSzM51oHb7yqCfoO0uSV7wfxHJkkbIWB6UgYCus
E37lleoV2uAM7PRIJhHZ3PZ5qZx55wndRoD6P4cYStSTawJLgTMsscjqd7PlyTeE
8vUGHCzGL35zIKy61GUWH9akIwXjYUqpGkFwt0Alk4gwkpQekb0GhkmPYmNXV6EF
1e9jDqsyyCW4LI8qYwXzj8FFJr2Q9M34Zg9E4AMlzJNReFS1lpmy9x2yeAVxZ/YT
Xr/cNr36UMRqc71nqSC3v+FDiBAJMoEP5Gt9SUa5yFzyHIKhHAU2JSf+ViakC0SX
JUWePYtJgbIYQtK8Sl7gWb8VqEBoM9aSdyPpjz5Tfj8jXgwcR4kiIy7hR0EMxpnF
jFcUdJm7Yw8/VEspfW4wVtFNvvb9nD6hwVMIfSRI2USr0SZW6pXM/iyeHZAwrTkt
6AuZo7OwWILtTl9JobGdbU0imOiV5Pxf2XXkoZAmMxTNbidR8ZuuPNt6uLMd1a5a
Dntrq8RwwSw/AYr+6eVpy4nLbapWGD1aH9XWsV5quNr5okolVxXCHTRCEQQg8uTW
CY/fJGv8iXlC1nNZfTIifMco4uvTWycjj0y6AaFWCi0Q32HhNBJ9ojqhVzokjgI7
dDQbunLq4BmTFRFInt2LlrdQrHdNPA/HZJwVp51e9FdV+IEhIjxgnUbUu44G6J2l
n3/59F9kCunm4aZsZzF12tgqrbaF/FgbgGeY0P+FEjU+ilwIlX+g4tY4lTohu4ck
rUWA97GkiJ5tj8xor8hsUma1t0Pg2QcNvD9nYf8vzD6Wky9Kjg56xLJ/YJwbnHjS
HJyjmX4otgHWrGEqrlx9DWXv4yCOIwQ//jtt3lEJ8UIRdOvc4ZKuCGT44ShQdQW4
kdE+anacQan8XrkmA3baIdNV/JTS5a+9ihTu/n0tKDHYigmsVmgt0Cj7nTotb9E2
jmH5b6+eARebJGcjbzRnDnYyGac7/OX37RgHChuIPL2z8TNanmUmgwUq3vxGC/WX
aTx1C5wp7ZkEedUcNMreoVRvh0Ig8AWUJ1id8KesJXZI6DYoWLacq2XdhtzEncCG
R9HXi6HgXIdGWOpS+WAe7JXy2Cs5+0p4tnafrGWuU+8=
`protect END_PROTECTED
