`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BtGO48BobeGgL4xASaArrqorjSdGHCgkhMYkTraz7+DCoNmg3KRW3AT7h7PixeCN
2h6c0kZfqyho233JUCyzPizSP96EVZeoGoxKYT5Z3mlxWCs48wY8DWAF7mzl19bs
H7YwHJyABrB6pmfkNN1Gn10cMifUzwSUfAOVBL482FqJVGjZlsUYCTXz33mv9IX9
m4g0iBNilHLGWbGH1zsO45dSI8SSTHZVrUJ/d/0bhkEhHBXEE0rxDpjE4QY9T6HI
9av/BRu2RTaFIbJ3QRjqvdQG7ksdajvOHwoNu5RYLQ31c1dWR9qJsKE8GyAWpBWC
YrbKehTLo5f0lKcVlSf56lSQkSmpGvIcrLUvz4phTbKWvlmnfsQ2FxkTmCWOdL3M
`protect END_PROTECTED
