`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4hrbmSFn/yay/GkV3WCpZiJn5JYv56otUoiJFe13g8xb4CYmYZETlKfab0ubUaxd
aiwKYM1N9VweYiGp3hB03pBGd1BfqG1/qEZmyHvLG9kJVYtflCbhGPFbipHjBAv2
lbg2jXwh5DffOh2w3AobuZNkck9yEjQmeHf75C7vL/97XKaCzqFUuHb/DinygiLi
OV2y+/oOnrVfuDG1Ms4mkehcVawAArIAo1Oi7ChNR0yEtVWf7kRR5WVUkHJ5ijnP
y4dArvps6qtYasFGhC5ufbypSAV9H8jRIviyMhkzyNHQBgMnD4VxNqX0lt5iUujN
T0ADZSeQWxacf3gs3Uuh6GH2UfCH9CC6N88sj6Q4lXjgnr6doH+TTDA/luT0V5w6
r2KUNIfFaPVVXojWt4wwvRZimuBtsApI7y8asnRgs02qNMnjRZGYhgymVNZkn+Bh
N9Oz4M8bZdPEMBLNqMGulalqqHvalKtG/gIfpBzTk3RYliBzmv3er9nb/7+CGiE1
Jzh+19RisU4EUE/oUeH1ovZRwMwc8js9s7u7YwuwQeIaw+VgVisdWjzvzV20wFi/
AsQxrdmu5zpbPB+VzlRSz7n3qa3VC+gEKwn3D1w63sYHFalNlc3EGRMi+4cVAAZo
ysfTkdG+dt0xrY3ns5oXQxbw/KdUaDCP8jNGUVTdvOE6TXa8EKcvkzMnvkK5PNxY
Zq9CrvBWw60d+rETbN9xYyQOUMOuoATmDA5vQdM5+P4CS127wXeTfyu+89Q5OWiy
gu1+4vbqwR1h7Vsw2UEn5wW2e21/A8qETiVb0uEVtXWqxhykjespn7etdKf0YgCs
sa9s0Dect9K6O50GxukEVZA9gf2l3g2wGc5qQinGJn8e1Jn9eEJkMi8Eg7ox+rSr
5hke0O6ZLcTX2gK+remIzOkXwUQ2Im9c1FFaVnmWq0u0ZlyXRBAw5kEZYp/zuznR
CJj9lx2ZMC/G/E5LsZKG4ovPrr2ZiNPAyB2UX80zfXdOsVT+4h8pXOnxfFjcrxOM
ePnOEnq2XRO6sgfCYrPnP71C8lrsLfyMzxYrpMzKEVORZdW3bNk04AhThyTmxWFf
T1t/fO7EsmNOwV9Rm3Jv+DurYOHPbvmUGg26Hc2QkXR0l3Aay576rzFEitKfcBK5
r2sm+kEWzdDBh5/LorgooB/t1N3saDcjbySd7/e7zUUotJnf8OVUWjR+lcPb1tpS
yWkva1aA+d4jzBVRHSKVadir2SHT2IC83DcHPHBo8y52DQY3TT595jN5+QfhAaKO
JKkYvXlVq8CFQNBPxe8t9FjrI2iZ6aKJI53WdGv8mxxX0aFEeMx39lwl2z+jAz6P
Nl6+P1sryXUYZOJgKMjVSks/QibbAkDJGVBcZWCgGY7VzaX4KBkxOOYtkpOCDcIk
wbeg27l3qkhtMtnZk6Rt7U122XT3pAFCMPN69pWGXJbZhuzXjTtyUp0q/mztbN2F
RvI7bREgZWWd5owu5fHZ4ppzuChMv6DBCpJ8whxJFq+pZoeZMXu5ig7mx4LfULMW
`protect END_PROTECTED
