`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mRB0mg4wrDPu62E6RHQgjIAuXg4ehtwG7mcyKA0zeB8zNVRG7MgEY0JQwHSlQ1AV
N9hBl9A99X7vND6rZCxS9SXB7cGcmrPNDjM/MSxkEPvmQq4/sYPKsMSfnGczZWdx
etTpD5ZcGirBCoHSDJKUklNK/grw6XFnwxTGn+Qx2hH2OR0RthSL1ri+1EzZlMfv
eG2Wyi5x/CL4ZM0hGCIh47j5vKErFUY2xPwAHZzkEHStOoLwXL3VAjyr0ttUvWWS
8t4ttT6mLANlxj00G09brzjfldY/Kzz+Im0T7Q6/DCT/LjB1ygMwVapE8oE1JXu8
PPbn+jxsYl5uA+UkWYjd7Uc5yPzcn3+Qy1ebaM7ULOxui7A2f9NgEK1Pt9lwJoQU
MTpdSITsxWaLZY1alP7ascj3JaFovAwdpovS2PLwPP1W2I5nE5TiVZuTJTu4LSA7
l+XNm8Ygj1kSFZbpiBAATocizaXR2ELmCw1V4Qa/RtLzNHxwTaPtt3Teqm2XydwN
8WWV4TZyPNGTeM+0eJ5LOW1qHXb9UdqR9kRhGgHBE+e1UAd7s/cINW4ndvpieECr
/T1PzGIgbMmJ5SXgdxJBNKD5/hPnz8NGmL5jN3HnvJiYhEWgitwXaIkYQ1jpHix7
A/qUkEGTKdwVg8LTbPL/hnRl1wJ/a9DuX/YlAHx+O5KQaVcY79ellwerRowQTNF7
fBT6MgTj7rq2y2i2y663Xn5+2l0JKm2CrI2//rpjug+uaQU0Ia5t3fY9Vtwf+PLK
LY1r32On9bO5ZkQw1Pi1mStt5tDRebAwOp9kiDb81BwI21DUb0HLEYulGOVfDH2B
+J/PT+vcS+inR4pu4Bub290M1lun/vSqUaGdhUEy/CQuVxRiOdTi61VmxMOLi4We
uNEbuFSo7f8SOzT6cDN36NAIUZ/Bk+DzCOnqqoEE1Mi5jbU+UVx7lwRf0DVctzFi
5ldbebDL6nVjdzP+tyNVpHjIYGVkJhnft4Sp2fDNd9oqcflog1WchR6tSxIZNN2p
IeTqS87nPw2LUEvbFdTPNc5z5dPBm6PCR1mw8HS6VR4oNnmmNmuQRYdwzpswCrSS
Kw1ZCV7JCmKFhjT13NnpN+Evbk06X7DMmOiNLXfiDkHzZkplwgpDqCBCOP+Os4IH
N7zuQZZcDI0KVCxoEGoHFr/lkaooulvvfkJWfajAPzXVu+NcLN0JgC1JBuVQL8D6
77uzMgIIb/mFRtbVo/OquQ==
`protect END_PROTECTED
