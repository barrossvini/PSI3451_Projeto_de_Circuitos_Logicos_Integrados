`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2UU98smuaaWUdAJ9YIbAKNI4YE1t9p7+cpwAOHSLk6/bzceXyTqErMGk5FNiDNGJ
BKYOXfcqQKlSMMpjTWUR7axUpAWycQPydklmS+oscG6W9J119uSsdN44ujjqJZuv
JvA2ohswmFEf8gTGLtmpukEECBQGiYDanTF22oJMpB3dqYBnC+Z+rCv1Kwh9hzb2
ZVIQlVRfztJeOLEnuf3qvvgWtjv8gkuKKhFVH30qcA0XUECZlak+VdZTAmp95BB5
KifKbuAgwR5Crfj+SLM7BUugLqOG+LuZSVaI8hLlSKvL7y4X8Irnj+HowKNe/vIp
y2DZ4oGpppt4fO2SofRpDzUjIIyCZyKd35X7kT9tHyCnXmiNfUmWoLrfPT6wUIZ5
VXUCJdFp4oGLjZ1UFxECkXSeWjELYFFHu9fm5HiqynKkXiJzkdEMSfcjfJxtzZeK
l8MtPJGcR4agL7Q8OH7h8usQPmCunmnVteuqTAECjyWb5fLntkx0NcL9hwqr5CEw
DUlg4+V1ncfgm0Z8wGm42/xeISmwqX40b8hkPc+W3c5/9m8GbHHvvoIa4ebPfZ7T
MXvC0PKsM5KBIvjW33gNHA==
`protect END_PROTECTED
