`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
43SXcg2CK7t9tO4mZN8+wZWXPvC1WK1WpFjMQD6eOFuRy/9NZNB0BgYNqeaDEvdj
LaaZ3wyyXuaLFhWgEEzsiTvtHz/CZu6zSfLcQspmO/Cmp1/KjYB5rNvF/VfSgGZJ
3uEKGPe2UAGeVWTYpr88akD8Zh7dP83vJWzgGxB0OXJ/WHINbux9ammp0EjLn+9o
9N8kzdOBfD9vwaU+huj+8t3wsyZtlSg7IAC2T9Q9pGah7gQDrsk6H5NltTEPlM+s
IHD7n1w07n8lGwHcb35W69D91KslFUE0y2TPnfifJcMk6a5XrpVcZLOBTCHcvwgR
ixYPGGF82JTaGBW0m5ZgbfqQQi80ZbCFqRVU9j9Mby+8tuiTVCLtw5FEKG0jU6vY
sFJeEwPH0gFYqTe1qE7ZZU4pqzXJGt8AqqT5gerDtGBGChZTFQoHgmGI6ysULdkQ
QreZaPK0jB5Sr870dHtVLIERv3hEFC2BqxJfSH1h0PpOssId6Fkt6SD3rQ71GYOu
ub0kC3fkJ0Wtm00F79r3ISO2hseWXu/YxVlk15Vgu3ng80+5HZWpqmoo/fUczanY
P8bRdFuD3L/Al8lGWCpvGxO2YU0LkNVE6xtRah2JxJFT7nCJiI/NKZDUYhEqAA9i
IsYjI9JdAqtyR9e3XOKZhxcQARaGbzVNDadauYc3An/PPMaQl729meFzC6DTUyUY
ThjBjO0vpjE+woHs7ajR3nvup+tdjoqbQRw5N4QPSej43u6A1653nYWMuGwbdDWa
meqh/n3PMVFG1qlwhK7sg/YONIaPshCUDQGKgdO5frL1U9t6D+Vn8F4/U7JukfxD
LUVmHa6eb8mYLsFtBLKabBr1eoot32z9AXJ0Q+DAoskDZ36Xmf8GT8+GLIG9dT8t
9o3Tkhfut8zB1my1ToD8BLucbSLqCDb89NZlXGJhBmIib4ySgb152stk4h97aBHF
9vOpQMfx52ATWiFCcAdZM2Tse8QQG9LjYRNM5SY+Tj4ElH5p76eWvr/MErXHDKUQ
Vn7GfAxSenDivNUJ5/BmICHG40AH1AaJnoQkKdGJ6iQnhe7eZirIYs0ApsCI9Llj
OXET8n5Ta1wVmsNi52rnYujClphKqEsCLdD67bPrx3+ZuLEYYb2affPmuPbHTQ11
tp+nRdbJ5SiOFNrCRKz2Gkl6XpIKbJ2tAzwLbzYrgY2B09GXY42cO1dn+DjNQzyB
nusdYqUzYKQOdfDmasodVYBYCBodZwMEIQ9mt2yE6ySXcRd3a+TqbIULCVocX7vA
99iB0hm006B6jzuy2vCRLIZcPJW5WfUU+l3PwoerIUwRwtOXPS+Daj/EHxCCrJyq
xFA565FBoNXemNpkNXOrc35TqWtL3Hd1D8cAImGmhZXMZL56QoePk6xxRy6UpfND
trbffQFRZi3ZVUMuin1nvj9o6b9yDF4ENTg1SU/X42jkp/VRoxd2uC19tqawmy32
GhyVDchGbODbjZs+DqLj/oZ4Gsk+fJG8sBZ7Hh2aoK/6E3C5vTmgkJKjV8rR1PsW
Ht0Q6ALkdsXjrxG3Tyq9gBBc0ka2gL6A6s9jhnNWIDBND1C3JwA+ZE2Fu/OlqX2I
WqkHuaX7bFmHYLgsQWsSmr4+y4cj2VxPyniwiTv4QJYe13qMVYe6XZk7PZMWwTOQ
BLXw2waYlute/2AU77l8OtdaUXhDZc1I6JCgVLCynIIZI/ooJ28g9irpqnS9a7ws
dXfbTOsPKaJPqUXi1VvgPMKc43itH6hQG8RAr6x0XHFM0/hePex/QdKsZxpT7RmK
x8EFG4n2BrvTAPWem59r5OKUF1+zGNtEkljIEgb9EebYdxQSsPAthnfRP/gJT15O
ctPdz2rfPyIMFnvA8UiwdAc81vrbtvhTmOrlyhMzI7tzSTSFMYUy6e1TiZCcN9+B
VrS8J4ETo+CNF9Q0wIB3NgirsfYHVIRDOIjV5oHSTPlfM7bzG0CijrrXDMEPGx69
ETbsN1QiKxYcPSRh1KEswTOY0nyU8u4GAacFIpN4Fps/nGZZYD98KM1dnMalHBfH
W1xdIatxYyv95VuhIbkqtkwKeP+s88Y63pR3Hs9zFI3Gabm1Sm1Tjq+HGuO3QBl/
J95XjocqBL5XOO9JWULH/yocHeUTKksOlSxC/srIC26SrYmFNNUNnz9ImpLmOGr6
toX6SS0/NDQ25w08GoiFa3a27Lb6ghyxfKtdrb9yIS4kZGSMJA+uuqoMPzOdfSG9
Xuo87RmDJsXecSJ9My0cI97Q8h/VQzkwRIa4kaXQQdV7aOgWfCpv+2EB+ygWTzrT
CnNONNMVAQRBa5zKHz/4F6HsrUyG3/7z0SepwPcUWGxljESZjgK0wio9PpN1Akjh
AK9rwubg8YZjNb9BfUGhNhbKaohAa4KUB4IJteUS1A3lX0dZ+d7TApOkzB/tJ/Rs
/X6vQFi5R6JCJcL4Pgv/aSBeElAmpzj1xaM2kACSphrlsbH3+5QjHfWZCNNyiZ5C
MIJDVT/GQ/+ehfxIcnm1bfElI9gBLB7CrqMzHBw3mV/96myAUudVCfqwyrzI5Trb
wVqywDOhG5iZxm8hxfYqqt82k37IhZGdDu0Yu6zO09Y/2lR9ybitVzSGeVfA5Lal
BKL506qOVB1hk+jf1JXWxFhhAwf1tUEs8snF7WZGzcdHfM1V/xbx+86MM/1C9x7o
YxJJQbi/krb2tyx0h7ZwYvb1Li+PUWmClq5Iw254+tBLumKt0+x2eTwVxHyyC/uV
xtB0vjf7JYVwFlGVfqZkaJR+GO7ij/d+jGYi9tgupjAuZGRkn98PyFpNFQpT5QhW
PC0dY7ds2RHqUPCb74K9c5ELBJAFgpETEUzmuAFQLS0/O9Spi52rW7ffPgK5ztaT
AZavcRksQ/CKbHrSoEg7cgQaQAHS5kqQtr/wreCcyNm8vkh6Towt9UJWrmzhT8Vh
s/aspPX+mOAO+HLq2uAhpfGl/IIqCHHkvV9oPXqlP6z7TzkPaVXr4pjnQo2hTVLy
3IFxgMVI60zolaQHaKv20edxCLax4InRIUvRkYn1cFnDLSawmeiDFLKSECbu4sFN
OxE3y8TDXNM4UV+1Qb6FR763arDwlrSncYS17EVR4XkmHiD8Clq8E7360e2o/GLs
wrpnCacP4TV5z3OpvBJ1WMi5JjiCSregGUtafYv0vmpVtexyMGyoii1oIBx1RB+f
3VaMSmG2vpKyUXOg6PDFVLhHO0nMgAMyD0LW9v1TfC/3IExApcRH/zRmq3B60Bxh
+XvL53ReC+g2ARDGcaVhHVB5XAiFq+nRB/19ukhuD9LB7XBJXanJVwbvUjcjlki/
5k1R3qDyyPkD53uLKBvHqBV0IUh9uUSKg/RGUitMX8bSaQ2og2a5fdFDToy6MkfD
bgTVHVmLLN4TROhqsRBc/WsKL0vDBWC1IRVOojekxAinTvKgKEJxt+cueD494BG+
PdyPCXuhPUuUGssAko9Q8MN548owq4p8ykdiLqWdhOYnLm53+B1OVWC8zU3jx9nA
F1GD0Qbbn/nI1fhdpDXHhwsdbvcTHn2+JyR07TQ/FcocjzL5d5Paj3Yw7t9EBStt
LqGJic0ztRY+M5O1o0kZXOoguoZespPX3x8qa05XKCabWwmEKjM151plvgoohAxK
y94j/EL4u39wJjgvGA0vh87Fma+TwcHvrB85kT+D3vqh7wy8UHD/4TzB9CAWL0Vw
Pf6J0Xev/l5rGKZmOfiG4cu1ipAx0FIMjZSUorrJKSwEsmhmHGky3UoKd0UorFW0
bs4rdNTp+RFJJ6k+AV8+UKtJ7kX9R+Nes/tHxHyieoUGvhQRfmN71jEh4iWb8RjU
bcSGU0gNUadq/6FxwMfdj3BicKVt2215goHbfF3uZ197Z0H8PLgVS/n7KD3WG8RC
6DGCpUAGohhyLX73faGYBtY07KYaam8MmbylcY2IRkEOfPttsytU9Hjt5mHtNQnv
ElNAKANz1i6sAido5WBVlFld+Q2CjjkFF2AYs0vI9QgPD6S0HykTNI7PxPmCwEo+
E4L+8GCh8lnblEsZvUf+QOlIlV7baifOMtlCqpBwermTusi3LN7V6YYW1EFnBMFu
qr16QuNXF59oM/bulj6bX7gMFLuQNN8VTzLygHkTb3MeDZNoe6uvCHHpm/Do5guW
1DqeXAIt07zosx07le35fRC4f9wyZHse9TpwdzGApmHuBHWSupJLMw/prEnrtZIu
E9FJlQq7ELsr24Kt71qtCMXXDu45jlQSQeCABah/EWnwuhie/1gL1Rba0uiARHe7
hN7ehvLBK9wPfsHsCU0sD79zroz0a/J2uEtiOUJI4dUtvYDPzhh0gWJsdWghZw71
gGTNedgbG7FyryvlSjeAGTNr03jjKZ3k2TYhy2/YWQ9ivwr0V8vZALoFTnE7GeUm
vuL3MXMCejt4iLg/FvgNzWKBaBHjrYqCaENiFherfZkZJEOvq+j9PHAzzsENAoCK
B4co/OS8GniVNAt5zMK5cmRPDUfJwjoIHSMHAI6EQKsnAsfOiPmxcgx0NZ4dQ7gE
4UkF2Cg8mA3FgOtOaPXr93Roa7eHfCp7KVqc0BORTnI6df5zuEJ6z1jCs3E0o53+
`protect END_PROTECTED
