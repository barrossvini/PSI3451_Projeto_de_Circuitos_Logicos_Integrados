`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lOS7P89zb5FpAEeFXYecdvtIQ6fWDdwPmslWpIzNq+8JI9zj9FcQrsZEL79rBLZU
1BkHcfKUhdnI1Qf4p2H14PkLQ92cK+36LJnGoQKSK+/d/ziHKfSO4r258iw1UVQT
XmWOdeWTRU19ilpvL7SwihNssNN8Awi6eO+T1Th6/kUM9GETtwrLks5f5825Ww06
w7B8nL6n3qBW+C9p7S0s6PXt2DoIJsU8+pXjKWh+X57O1etjDmTBAHx43Am2Keeq
k79xjF+z9HmQv6Wf3ZOhi9lSCMEsQHh8XUVN66H71FvpqypJaTmemXvPuxaVEM3l
crFAsmbM0M27MJNr7xKKkdEFIXNiX7Vq/MKobaT7pzKUSH/bkiA/W4wrzVVzllAr
J08o3BUyqKt/Zi9cfYIo1yJ1OiCeAO20JBrzrXxflz0UkyJLYAF+mcOkqibelPKH
YwhD39aHF1V64/bB1/hBRc4xAPNomRhaPJaQxsx3t64NKZQ6WPdSBTlULl/J1gJV
HJPZxUSK2wvvDV5mfUBMNVWH8tvvTKKjdkQ74Sv3EO0r2Rwd2e6V5bVg17EA5gm7
7C0HN0UBPZ42v3Va3g8FLQotJ2uq99dSCZuQoDVHBRaJVBSU2stSVzMdA3Erp4gQ
PP2V1pVve3ivvSqnv3hg+O0l04cTX2YM/oARb+fDVlNkW4KKnfOwR0Pt555OuBGf
y7F815leyKHI0TykURhHsglCPH7LDnJ0LRPQxFp8QcNu2d5Z/lpvz67EareLdT2o
gWiz7QPjLqmy+NXqJ4YQLRrPI1Uwgc6UhUNglhfspc9AJc5+dngbRFvWcKb90RvP
JMVcR6uvpgBPR3vvE12iNcZsRR4GzVKiNAcKC+PJb3o0Mv1SdS5kTawPCT7GrrQF
wQXxNBD/4oAA8hdWjc7xZo/f2B6392Bx+sm4bH1gG6oPDEZm9xjocrDywAhZU2WK
2Ne9gHxH27Y1xnKxbfbUXAv4ELegSvW/oE9Pzd5Il95Zh8juxzTVjoqXYqTuiuX+
2beuOSJWzEnvLb3VBYBBU/QarCX1YdKytbRMPdRut1wn0sHprPem8idCLhVhAjhy
hNDSaCKoj0zwpoHIzOKFDx3yXOIqLg6Zkq/ogBohcJdtOubo0Lu1MAElPQeZPuJx
/7Ggk6lbzJycZcuua/rodc3bGXueeEan/z0CxZ6LMbWEwq9WbTW3jvJlLUxsg4Ke
IeqIPe+ggycl5cjkOZP2FDmOBGkec0fLlN/8FD5rswa3FECmWQOCiMuma557TH47
8rIYhGHGe6XifwAMKNImB9lLyB7uEnd8x/yPsVlJDAr5xMStyHZ0NakMD4CEczmg
yZ3+YYG8l56aUo1eH+014dXbzLIqqHHuQnX4OkWOFeXBtcUfZh88Ldwfc45unxXy
+KT5vl7WxNrLqyGdyo18EpmZrM8N8MES5pu8p79C1dGC55LnsyhHVBHz10wxQ19a
F6iy8GZOqp1DNwAv3z9+izOcgB0K83DAV2ew2fk1rNgGZlNa1DJ7bT9ZfuLtlSuc
tO+kfu8n8vPdCXqiSKnviCXZy1/bokpLZv/4+VPYxuLr3wOqu+RxzzKMuytLJsly
h75EA+i8lBjYcSUfihtGXjy+Mld9zPh/7u9erlqiOnD2dpsd0ZAfAEk5y2Z/oxLI
hSQTYqEjr67Vv1Oz3pinUOp7DvexieUDv4by1elDaiLs9zIlovYwfB8QfYZWTofY
P2jXARyS8VbageMa7lkP0z8i0Dc/613PyLWSdvyxo6RWqCKKOIU1ibg7QFLgZ4Ct
tRXy6DVdHWEEq6Y5DxEsy/SHzAK57f5ro9aJIwYE+dbX/Y//vuU1b/PXLuND11vR
vxBPhDdszh1HC0le2IaLhSDRrHXVCL52uB69lFelwel2gnV+2ydqOxi6bGR+bJ5K
8MoEPaHA7LR2gK0Xhv7Vk7VhEE//aT0bZK2qbgtnyUjdpGRuIV2EUVkgReGgrx2m
4P/uozU1haCJ51lrwcrlz2eh7BKNxqdSbtPRV3s7dyNXshh0kWxcKR4DdE2WHgK4
/7MbFPKFttoJixTBAPPpqWoB/cJR5HBdQBIOj3BnyYgz1vVlPWxzTVfCWnNXQf5N
D7HHhcGy4UhS4vKUJRSqMT+ZxiF1SW+MJu8JUFusEyHtlpvhSGGw7vg/jnJ5vWqS
AqmHsWKAqjsDw1huZl6qyn478racpHQonsZVuoV3/lSOXilR7vMP0pwLBuxE6lp6
45v3KxG9T936rMP9DQIOOujMtqVaXjwouoXERRa5zCEtuQFTJ2/ZM9YWnzvATtDK
GY0+IdWagvlCloBeFZLo89dIe3taT7ufdO1OEoVP3MxaPJ6diUFLwOGPlXIwR0UY
6Tjgm2vBrkaOIyfZFfW3cwaz3HTfIBe4HQ5baRm2+SDXHmWODfZN2/XhBvMf6vEQ
RTBe5K5i4MZrzz11/HUjeSVdHTQoaZkK6eGuR53p+kqxNboNVrE2msWsr8TgP1vB
n8m8qtwuzjNgTXvwQdhCRZU41Hdz/IbqGvCBUcEY26FT8opD1n71Lp733QjJy7rZ
y0rqMizpQDTwgv1d6MtgLzdi40t/k5IgRhtSImjM+Bbwf4xQx7JQvknXj/iM3BUW
lqGhkqyRbu4sF/ocyZLqhSegpRYwXdbxJpI+p7oM20c8fhiPlKvne/TvzoLnVUjv
VaQj/t8LmloOX+UZ4tbg7zMHtrn9VDAZM4GB7Kggovy7TQAAJnwVxTRHAUnYkCx9
Bpnrn2fiGJFo7fCPGH6JEbZmgtsHppVHHUG3/v63ZLz8Dm9/LKHEZFoc9fHCUaPl
TdufXUpT0GxjDVsgjdpl+qe2c+/klzA5NkUQkdyzSy0mk96L6it5xVHawHB6+768
H/ljIcxc5ndiNibA4i4tQ+8cv4ftYzlvgA0OYUG9tbtiXL0ndSx8gXAHI84kpJFS
YX46MBe2wXU0vd/nr6LDUJEo4q6h9Jz19BGniYXjnISf8/o6lICYQP6Ljoj2T3R3
NUU3BRWqmnRSObnebvgbdT2CFGfJB3p7+7up3vrl/aXtlkvLWmzWtetAsMX9Hgb4
zUrmXdyIWhQPn4GnK4qNp5XfgTJM9WIlmdrdBwIUyfIrXfKF+XCGhD6PDqpSjf3y
S31bn/7ElyYVoTtvOCJpeh/ettR6+gCuJWWZkDlswYXtc9SV1CD/0cyZ0+LI1Gsv
LB0UsCGfAu40LgvojYLyQrcJwzUwY1qKJqlVtQd1tMBVy3l14IiGKvYfq3hMUYcq
YGSsBr0AxIcxeG15DAlefyt1EXoQsuKL4LXpTyY0TAQ4l5GpmwQvhE2EJQqOYXCh
LupSDXK4NTk5vuF/kD/TdQtvWrQIgFkcgHzWDCmRNmxU60d7JpvLzn7qdiz74Bal
Up8mchBts2N8OfTseViD6IiVwk0e2Zt2PVWcQQkE/YAXCpyI9iONut1u+VaR2TN8
r7VxgPxZH+NoluuwHxMWY1JlYZuu1APFym3pAEvQdwR1KY99XX0LbFvCXGknzmIf
r2g7HAMTlB556TtbBHW3nueh8cB4UmQXKlxaL/Sb4+VjbarRAVFc+rFQ9NINEfjU
5SAAMMEfaj4BfBySiv0JMKa5l5G/7Sq0te9IKwojRZILT/zULe0/xmvO8R/qxmTf
eAIPTCc2Ef+MRIdSVRo9qtRWh1OxtRjCjj2b3z9LgP+JzQFIoveXfLK0BQb+gUem
2HMUU15MSfItG7CmAEJWkMlE9wXGMmBBfqfT6B760i1FwFnDO6cFFvN246p0jl+h
0aClFfEPJehSIp4W5vi/6qIcLlb9FrSiFWnKvJb/WLWHNyebZViGOjzTXbw+h+QH
Jf8PxoNTwM2BiFgF/EIuEHbToxk52iCXIk2sk3/okJSxehPSFZX4mjOO3GctV1cy
Mrq0nf7BRGTnn8eW4OmHaxL9H7/65zgJWFP5gGiG6aQ0unh5CEZj4KZJCe61u5Zg
QUTeDMn16te2f1c+8ajT6eGwuMe+gU3FaJhzhZklIBBSnDClEs9t+91qE7adTZYJ
T2Y/G5rVAjfXHTJNyRKu8edAw++tf5grTdayY64+Cs+UP8/MXUatcGXxSo3SRJGP
KbdVKQMJZAO/uA9bSjN5lVjGM+XqTjcdrYIjXEdlskP8ETI+3mxQsb9FoRwZiorW
1SWZBRneVbL6gjjq2LbZB7aJlUYawguI/xGQKnSCxpRZAIUWAUaRB7qgzjmrZqFs
Dd6sFTLSddRzKf1WXklCFWL5Z2/DAiPVhw+a3+1Q7Vqx9Qux4cb+/rCYhTjjL+lT
9orXObvGSKv5OqqoeaWlOaF0V4PDB4VcJ7C7ULwNhrccJO60WWrmKwOFbJdxUPfG
T06lUB4vrGeZ/LHYTLtdHk3BSRhwKei4/HcArFRFv5PiiZsaMpYHH0K+4eqTFGGN
3qJ4uZgQ8GHUqory1NUhXQRwgCg3XQJxc1IVNFdstH8t6rw5z74G0aIdlH0RVOE1
3tfI0UoVqEOFE2SVhLZuArg4vX4M5t99GgArzSgihK0jfkJ1lKvxmR+FplqtJxZ9
KZ+nqrrcN+5/gO800DSrXPLioyZEyTJZpoylZeAFc0XLfcBID+4+px01xIgujFcU
xpvdp4u1mPVfZxwJsG0GInqViDW4+AZ0pArhxKu455q8g9rhsazfOg36sJJy07c6
QKkAVl8aOeOzsbxZGduo02oo3shqP+7+7ctJ9V20jQ5Q24tlte2pAwz2CxQXetfH
RM2syEDf32Ty7TKALS7ccSAhB4P1RYgeNoNwfABUZnvD/oZJT5t50uhXD8rdTh1a
z3TrBPpQM2CMxotgNI5o/b5mhG8D4ELqrMoi3UPa24vbs2g/jZqXcEQQ4uH9ICTS
ouI8oce0AlGi0yNssAKTfWACH60N+6beS6PBHkeX8T853wwisuYe6zH760dhXlcZ
nyc4LdlMwkMq/k6N7NT63CmXcJNdP/JjEt+aupfvlbhIsQ4zNF7hcNCIuTRseiB5
IvAR2IjRCc7/qU0XtzVDmxU2yKJkGwYigHZfGzvlJ6BLUfD80S0CN9MOm9CAvXcb
bLDGyV4Ylt3V+KAnvXjQsuZpwDeiV4Tr9eeHjLBKiHq6PdfqxbtWNfQ3yExJdGfv
krTN4oojuhkJIBiiTXsh2T8M/1sa1ToU5ovjKEuD16Ovwau92Kgar9DVSZNxa24A
U8YJj4MSPuZBae106QwEoGx7o+lNFRV+Uq5A0XOC9YwECv2Qt21VbL5vkDUSzjtP
VBh3HKR7m+VN9jFWRadv3L0pheg0vQ/lbCLZgK0PhfKV8jN8PIXzNwE6daftefEK
C7hS41irMK6U6bAHvPP5KCmU0JLMBbGi8zB0rxpIU1aXI+Iit88Hb0zO97u4PZYc
rlDaa3uX6D8W3dllpmp58UmlAco7z8vq45NXWf4898WboYhD1xTFe67XIguVJzQF
jNbey+BRX/VkbS+AzwHoXBxIZpHO8sQFj3Hra6TqUIjiDKN75kPiq8I4+mdtW/z+
zC5A5Rq4SUCBH5eOhcuzUYElnOZUl231stuseGvm/tnAZWzEm0YCcex4JNPA41B9
iX7alVqeN/hKUOET26lQRVv0+OPwxkZL4/4/Ikyw6lmwWwcQa1a1zueAFcaKlEaf
8kkaKr0BsiZpw8i6DCO4aeH+1UToZA9GrOJXnKMFeYKiTo6+b+GttT+J/gR1nlI3
mw4tSXWqe2qfHpYenvgi4liDRV8GTBRdvWgJVMBBTvo5rNkU22S7Kl0JrVhEl6Sx
/HHPmJxyWjCjmii5TDWbwZtEcIJ4F/cDKyLX2oq8ETWVR96KDslJF48jh1pPst0A
/QBvqnsbMRPxvGe3X+Bf/ABS63lZhrMYEx5oUrD8WZY1Qk5VJsRY1NstKKjQSyZl
txVAHB+lamYVCUAU6sctdSC0Ws4ksWowZpKro3vNiZXjqarmKrpzwtEO3Pv766s3
MHr+p0yZz0i2nn2TlYfoQkiVaS1PsJIzVfE/OKgbTlKuNWncgIZGJjuMz38uth+E
CKaa79S5xw/TVGuhYGALr4y6PF3G20PmRpkYAh+KUuV4u6OJvob6JaSky3+M7g2N
TXj8Q+IpsR6as06jYZuUc2ssXyMyVqxo7a+6pr/mVmrlLgFC8qY0FZ+UY1c8BLve
/wQmhGI+DAgPNRBswqMryCBDRr63hO0UyaaP0FN9mR+qjCyiksTtvsZNU/U9eHd5
k4WYCPTYb0L9J+TDDzk4IMNw9LcaC3HprlE1ZwyUwnRFJFg84B0lFRErbSTK/oRR
4tagJrbKM+ZQCV7FC0WqhdiL+GMl9fXevb79sHleW1q103OmO7ffmmLhAMNL8wtT
FqyCuESmJ3pwmTL6Bnr2iIOhaQwJEL4QKNto3UXR3zhjIs4RDsLRQwkyYq0209T7
/UDl4ebdATPuD6aSh2GUVJr68jMhcolJEODEyHWy1RXw7PyZnlT3SDQxmzD4FMkN
HGFFnbYyX2iyltqHx+18KNZjq5+PK5ZECBkhgwYAePT56gScZWLpkacJ3ghelKJQ
U2QAJS1i7Bb4XM7vV7hePtuWsYuh1Y5/TSl31jao2cER5YJa9ILdtvG/cQksER/F
rAWTqtSI3Q5NRF8/XoXDrh6OhAMtXRU2Qv0xf+vFdRuwd+EMGsChc3j5PahRaPMG
JBDGmGooAiJyrMiu7e6jrERhgrh8hJb36g7JuWP38jJSuWf5RPHl5OR/VwkxKQCk
U5Lxwh93ETwYITaq9hRQORU3CgZXG+C+q4DL47mQeAWsZb678IArRoo5GSkKOEHV
EoPHHaXNcxI0VKH09ISf+4rKYM35RNHQjtPkgLJYrVlXvtFXNZVzh9sFt7ATPtME
6Siixzy+sNT0i30EFXjBSmhQ7DkccJodMQTh3ah+gQx6nLQwxukzY3KE7wUPHB90
vmeVpc+SKrxCOOF+0MXiuw0nZm/sAOvf7MraDixv6kCcb6KafHAkZWY2DC1CjCa+
1tiW9PUBVQmEfIpWNCXvlBT/yeJHCY8jvIVynt2vWjNKcfW2HOQdc42wj6bwM+4y
dXM996GQMRmJiIUTmhf5iN5SpDJvZMH56/Ve/X5dIiA7+QrwcEZ1TkbsJpM2gHit
CX4oVxje/BHoe5KoTXu2b9sPo0pmzRy5718X19S3dL1MYKATQAnzvS12GOzlGUYZ
betEaSSSAhcXdjI5Wwc7gSXTaVOVNLl9Lw9ygazeSKukM83kkesEg2aWDh1jW+E8
iw3v2tv830wcS67wTXanWs1CQXsp1SkYa6SG9nasL/WvESXzEQk5Z5qB0rgCJfnX
ScMskg73+Pkestn7pZrB0emPkiY6Bd/YFlElM+PivfYfTvTl7AM62rrYJhryNGPp
hGJH1cQjEsbWA5JsBxpK7b57GVnL5Rg4oGx0aIJy/3x6bewU4HvyxCkwLFgxRvTI
agrSRRNuCVeLt+MAW+lxHYDnGt4YDiJwqOGw+povYo2K09LEFY0L/N9L9+kpi4+D
5E1gVtmnnzJ6Yc8hCSvucRuz14bWCOSvYr3HDRUm5yu4RqmzNZyPntqefrIeQ8iE
hoPxH9DzMV7MObswKta6JL9lbjAJYLaLxr/lmdX8oQ/Y9cep5T71j4BdLjs4vsw7
Q9NqAf696cSEnKPTbpnYDPDlGk1ogiQNk+6dNHWH2frYjS5/TtYzXeTc6YqfO+vM
SSaxZKoI/iwrGYZt5C1GK7DIRxjEuxKB3sUDTvjJhfyNDqq5f45bCz+R1qQCLhBD
qAxsfeGyyayIdhVsxBEE6N9PFg/i3lWTZe0ZA/HdgydSRIhRxz3Tx2FUTnshQ1LY
HAwqEEJuqDqLFTwf5LKlG9BllqQ2xlEMvAsBlSCa1eEBkVUI8pQJ4AHuQDD84KRa
OcbPi1jqaCanJ13z8ybYdFmZCoIYokWeyOaTcM4pxdqvLfUhiE5JovkQFCiVrGHI
6qeM003jZq3+xZ1KsYr86yD3ckUto+PMFW9IfNWFHdUCGCSrYfJDlErmt3Gzi6jE
Qky0vRuhzIG6bXfJjfubNWRmranJpDeOzwSEtTv1kzL1+8KZ3LQmy7ShlZsMVVil
Sa88YeFMNx+LU7ICdslz06vrQMXgkxjMpI3NDsN3nwu/DQTUaID72YIFM1q4nJIB
/ylyrVfvXiN1GANKrgoHa1Etw4+UNS47JvElDckTTfOD97nFYgdCeURNKIBBHFuk
xlwIDcpjPHn6+u58h2JlwOnfDu0T6+sLx+xZaNg2FYV7dkI4bptNfW+4eOnJ0RhE
vcyPOXE72td2Ps/wPXEmcVg/76jXyR7UNWjoX7RHG2dGdimhvD3hTFrOw28FYDWY
C4WESfprjyLHUi17EC5IwRIEcXO26kTBlCYSnsyJMoCoWSDBOQ5cIUYLabCBt3t+
Q2H/AyJWKhmGIj+h6zG/oCupUdB3WedKm7fHwWFf48z5oG2o60xbGzmHmmx7EN8o
ivBav4eyKf+miEf2KQopFVvUSZWwLB5IQ5vKOgsIUxByBC5JhCS9a2ym9VTzOq9x
RgPQDmJ4H3rl86Jn1NMaDPca8SFlX+HR+/OK/qfB+21RPoh3XGikct19OKWNvIS7
2tqcGjeQYsPULqsnCkphWBuw3cfS03DMbymgDpxdBT4zt1BSxfBMH1uzlaqehuER
58d+Rjl9hCGYOSgWWdnhwT5U3vOIPrScuZSUAJJcezfrzIztpAkJMn+Danj01VlF
vGJPbBtxcXd5a5IPRTILbZmGvRY/PxvcAS1MyKhSOaklmiHwhBrXI7MkitIa6ck4
zG8F/ksKe/znyv1CNoEyK2y93x4A0xFN13RFparF8zCxMwlYBCfTl7Q/roKnhfiY
EZmMXeMiUFMtQmgDQLH5j56gGfNPJZtj0DI4C85dxgH1TdQphSKJgotok9+Lpy3m
hCf2Ux+PiPXWoEbwW7zIb52ajNsWA6hxztJszJMU77WpFl912vJefl4RyRgORG0R
fTtxFgvBFA1QqsXD+ggqVb2VirSNdq4c2H9Z1a3VIJXpyXgAsXA4VhCFyKix1i7S
vvJTwgAtvQj9tu+deqfgD/Obl6aNQ0Z+ESc0SlayggNASqNTbvABev3c5ntDfJD4
UxDSn7f0R34JywwD7ci0jqXQA5kbRYLWxJ5g0fH5MGtJsvwoc8wHcBWYiNr/pCk1
VmddvtOXSXCHF8mpANFPO5XoQ7sFUT8D/Z18QuMAKexn0wms4ucos1jsJBF/2CBQ
cgAC/LAVsUOfcCKcQs2ihpNy+CPJswxV8iF+fnCtKRQzqV0KLFhPDfijmsPloQJD
Bx+6pWCcsxZyIrTYD3S+AJBdfwkvPaOi5dwrRpFDoHUwlQpUjHsESX8eRd0Vf+1T
rLXjWKjglRIOBzK8QznYDX6/cZ5ivk2SoIemfbiYcud3sOLttumTgpLMDMFQHDWj
jiH7QWfq4NvpYBplxe78+lPozTZjQdZUFPNWBVNd9/8E5gfy/28rkn5F2eM9MXS6
iCdGWEHX0CsU82UcbIzP1m8U0Ljjt/YGB5SNQI0zKFWrCz/g6CAORTlY6zV8wmJ3
U8kLD7XPa/VkOgyGt22TenS+BPp3n2WtuD1vbdSpU+mbsOrVhZiNrfyFVTZqmRdr
4Oml388XZUlFgdt2WrBErUSR0/wgJiCj+9AEQRB5WdOrIae57aI04NNhv1vn/tUb
JVKZ2I22Y8P1oanHfIXhTAQurYpivkDV7nI3Vvo/Bp81oA5uHUj27j/+Yh83tYA2
4cBcRGpIbD+KA7Me4afYOBZs4qVb965oKxdVbRCRJWoES1aIH5p4Z5mz7ykYglN/
Le6ovcMmW8hyDcMHt582ffa5jgmJURr31YVgw3RXsrwaK6zCXeFaBm1HAsaaeSPX
bZIb0jWrxQXiwihs3e00IfbisvtzJZ0iIS00j8ILku2lFrFe3LAArhkp9ludfuaW
uLSd8ydflV1ASu0YZjB38QsgFWOaaDy4qN/s8uiFDxpg8nsZfDsTju8Xcr8c20Iu
JLfBq6ya5B+AsPtKugcbuiCyzfUuBsJKYBpsoWmkDeIM8DE8Y5B2VB4z+pTytXeq
ppGfYMAQVysUlqXtT3vY2Xg5GXXnDb9J1Obcbu/U4cNSC4Cc/75YlfQVkoEZecso
ny25KD+lKwCEzdf7xpSM1go/Kyd6uOGej1gpUD57lKhpjlsG5gafmJJPFuz/qa3s
FgPcAh8Kwi+Wok01EPh76rQTBdxal67hed/xQZfW9F4oeo68vAKWJscUusnWnFi3
h0Vjp4yYb6aRCrubn7EcKmsQSqNXjPI0LkKQRrgHzGeUFEJzRydKKsqKIqlo2vF1
4bdrmw7bSv5kX3CuSv8vhWPMcxFK6ABoWbk5Dgm4tkTha3XTDhISLDW1Imcpe6+8
Dk2SqFVcgqlsM9jr3q+CxQrnhP571FKt89uXWrNMcMmOdcPf/Yj+FJUxMooVrMxX
skQf1s4Ml3ZyuLdjvINQtKfQHe41GiK1YavtnnQFNfUAp5dCURNdh6ynBC6n8kXh
6SYDUtDj3t0gSdNTHhq2uBad1RDAVXw34pOLHrHDarmaSY2nSxLLZPEYGbxicWHF
Fn+TobIV0R9u1eG2qGZpn43N4h+nVCWhoTLj8hEgZdAiVMkWddbdusRv3+WYzar1
sTlH0xghQvPgErEBPJPdvdV+sjo3KzxfFliT9xqSAqzDVVbLdDhTzGHziOIf8nX7
NlDKF8v/XIcPddxqmSyfplsgTl3QV/bvbflcNmYRnE3RrdNlDHL+Qp1n7h7XbEl8
jTFnHc1PK4/0Vrgh65n6KDnOqXSnzk/WqlaB00zC59duu1225+4fEIeR4I/kHHDz
h+gr7E0H401e8VFzuGJUH4e+EORcFIOPk+PKpXrjzvRgTBqTY4wLgvBzLwu47ouW
RlwJtdGlCSGtqO+DQknLh6zqni25yqUgL0QiZs3H4Ls8X0rufS5TDa0tZeT3Y+Kg
4tUzPpzT6CWz+WQtIdG0wj7featEm6SpfphOq6/NXih7WTsu5EITb6slubeKXmUt
lSflGyAqjvcJ8Vu7a6MRM+CiWyX0vB8c2rHQE8tFl8Aqa06QQpADugHeUPzaSLqB
RgLT8mNzpJOfntqwMEBB0UGV/DCmGqaJ0SKYW13s1J4LFwj3M9kyfhuGH7r5idCw
DXMPniST1V+qvou5Y7e8H266Wqr2r52UUC6eT7RrRxAKvMLYc6e+9msBn0md1x5R
MbaUSP8VwvTQURJoo2CPoNXOD3OQ7XMJm7/JLzwCejBSge+3QeHOMEmtjTHtN4rz
k8J/LDwmMgJxWu8r/WTrBzYni782Ji8Yu+T5C8UTuAdaf46uwzJK+zP+8dxAVJz7
pEDsgQFj3MM/R7IyjIwwQqrAJ0N2AQ2KGIqesNGpSMORVvG0R0lBvQVrJ3omIGWS
84Y8VEIDqsLWn9WxCUIajCqH2EWfZ2NwYnIPWkqRSrhbEZ5+008UYGH9ycVtDLsO
lJpFxviBgJ9HPNrGHjwt3RXqqqXNYgyRg31Of1LLLcqAamHDA88nSFrDto6xGaN9
whTYAbwaXC+4wtg51J/AIy+geFNqeDcGzn+QnzopvJwK2Gbrr/BDpiFASF5Mp73V
BlTKU8t8OG1uGQCFsNyya8SxdtXp2jfvKkW2SZYHBdXLobiTEik7KqO/AbiUiJnX
a6zFoAxyWR+ig2fnRx5pVdK4+vT5BnzeEfWWUNHujcldJ6QzMwOBvYYHUU7/Q1pB
4PyXtT6nyY6EKGlIrqvHiCkh/akrwvznxGl0cJbmhRRzZ1h79+KHKAL49V1FWMk7
pgP1Xdoz0xM9pKuut9BOotMrF5FNaJ+jMqyfJ1EpXqN0b1zK2HOJnsdJ9h8haoX1
YuofsuY9XTe/qlVahSTeECNLcZRLfWrJmwPyPlLugLCb6vp1NGVdSswoY1B+10IK
HfgrrFOVuo94fs0htRbCB/mfIKGYj2y2LTYLIKaqCVSDrKhsJB7RXqoixskF8Z0c
TbxI4zGqeHQhNZF+3Berunsh/bWvwQWyIBnxFBLPbacarK4/Pq5AKO3on0J7f3td
1fXUK6Nt1WezCwbDBf6WFtPov7t39DObV9yyjoO1+jrHLycnIvu56INIrUDsersk
g2hD4Fxh6nP0ifvCa1v5ZQN+51q+1/QWkc403SrtWYmvIi1vMtSyGcpFrx7tTYuf
U8taf7PD1MLdw48jp6JtOXW+9Oj+825bofWmDdCu0wwi8fuXH+U+s1moXLRI3yCF
bV8skrk3zoGFVw5Byg8r3RE+Bng1ywDKp/419d9//VY5YqLj99N39rdvk+jXsjqg
7vxBY5ufi/M7dMmEJxSDuYDuL5rUxWbBbNXswWhFPkN5f1TuWIDZnLMASdt6vt6I
9EFo7s2lIdSmREfxmmSsYa+qWh5hWBCoLspwD7BvIqmlKqxAfDoQMe8sHDqIRnm0
xOVD9TdNMKXf/+TkOFLuKE7ji32Ddr62/7SsIIK1YOYuL+aM3jyyNbsArISmKdi1
yPeaHuO2QXQTc0dxJIa7cHg7o8z7J92y0apljV0tuMnPpI/WJOoYd/i5fppYNyvY
kKA81SmczF1fsyDcmatCGucBiFPofdLMcYIbo/CWXseFXn1IUCMdcXHzLjC5ap/S
lFBbcE8/5rHVLG5D5nHzrF2NMKbAi2Mm9N6eUVkqmGVjGx5YMChLTyiLNh8Xd6fB
zb1EgQhZAi8GtfAFC+PftmO31uiJLnAKSOi5+M/OXrA8aqZvYmTExj1J7UyM/Ixz
W0squDxrXz9WGAdfGKrpEDoiYKShCdZ1wVNcVf1CPnP4UJ54+ZqSemeoTFT3zmHP
9F+/ogYyxZVynZ0quhOxl6lcawmF5g/7Q6rV4afOMp5lL+OFw3nF6/BJoV2TLdao
1yDaVf8wm/APx1kCoTok/Z0Tcav6TJe2nIiyxJ6zKXNSgW2Xb5OSsAkLKS83QobN
SIpPZvVdwZ6oOqKHiIzalWIzuSUxBIvWxUq5J63PLRN0Bkfpu3aKWdRkuej6G+kY
7hvI/ZmYPDL42Jb0jGEiUnGlC3AcIFcNISfL9Un8ky/oK23FIJbOjYIyz2Sl2Tvg
SHsabnyJ0UFul9+G1W8A9Z5Mnj040EdbrKtQdTVjQOh/oUKf0GzOXO/jyI5sCeIu
xSyvz650v1R0PoUjvcGOAsh8+xkK/cdbcNqvgcL1p7ek9fcrF9x9i4g3zRPRqEdk
ZWxWwHjsZRZNJhyoUMmkjKCVIC+AToZH2rCY5/jsmgPgweVXXtWUgJwIOWIky9Cg
kUSyfjyU9FU0EwKDLVV+U5zywyEtlmakPrRKnyX/VT+Y0yGNiaJqo7XXBFqTNtpm
UYRe+xlkAg4uisws1HKikF+SPXgCRoagXWLoJ8bZKurktdJsxRqwvLYiMdhJ7hQ1
PDo8bY1gstg8XWMp5tHKy7w40gP2ZYcQGBXSvD0PmKHj7w7s6mPaPJ+8B6zUHiRq
sTxed5GkxpDkwqrdwa/ugi+T4i/8qvMvygnGq6frdE1eV/5AAW5XPcQYGdOJeDdU
BbuxieW8cdhCAuwfgcgeOZhxIdtiO/OxPrwEsjZWZ7abh7arWgfDAP64SEwWuwf0
ubxI1a1b3j3J4Ek+rcSsBvbexo6jWzy9O4HMHz3/L4h/EgevISNeEHfvkxKcAEsE
BTdm6QKT46LptMgbHkcj8WK5HW5rzGXExZMmMbGd52ZnMzo6Ky5crwlp43TC/DND
c/Wm99htwNgpIv2PaSBeWmD4j3NqlPyAAh2UrWeZN+SfunH0kUnLbonSJrUyjUZR
A9piZKP9041LxaWT9vDPs9TcEYFvy+ei0f+Ql6+7HFBtvSutoPeuszEfUwkHq7Kd
X7OhNR3cTPBJnGe+Arxfb6Y44cdbtZxfPPSETRgIFi1A4oeFN4b5BztRA8XsYwI0
FXegxup/PvliOYqftuOEwgsLHfD0k48g/qAj8g1U0zczcI223f0Pcx2TYJmWfNrN
Iq57khE3RLobEsXOXv7z0bTlFLIO0eQ4Ug0fu4BSTPJDXM5kn9C+L1JzwYnBghRB
HeWmQVemFiENkoY4kQD5G1cXr11TTw6KiF+6/WoBXKVkeWtyZB9+yUZ+3ZTBmidq
Wx0e1IorWdLz20nuxJStqliEabb11Bro7vX5kufMsYumbJx6abVHf7BM6PpkWBjv
cVfXl8zgKvTb1KDNJKnZXSMcqK3agSCeNExa2uDQeT/wdg5pkPLh/FF4G1RPFyFU
8z2X7yKfy88OOOFt0dGk7I7mlIU6ex5dynPoT5oJaPxAxDaBhbWhsZLdokVmCnpM
QaCfQcRl9S/XilZaLX/x5Hx8elSC78vzLId7l7HF4Zm2Q1Af7YilN9cCt6pR6+tk
+EPeY/VCUep9tzRjvsD2jk0OObedHOU4qQ/PG9s1QZJgsWb5hjEVfAz39D6u64yI
Hblx2g7ewSSrWthuXFr1wvrcDbnxdc5nN/BExmFjx2Z/GkrWK32S6MifAn26Bb/m
uuWzES8FFnCoWyIrp6aYKR5X6myTdgb2qZx1ayz7tLGhVFjlv05eSk5MB0LVG8mC
oi8Ftsohyzlghyyx9vEx7EiqevouyQCjfr/w5Cbk6ckWiUI5ET6LsvKnfXjo2sVz
PrjrXsFtXCL8KugOc8t9o9HpHSUjW5LwL6mESKtLyXhpqR7Mng4Oyt97SPM+rm1W
TBan+RlUJtpYggycEfr6U89qx3SVgyfFI5/Y0Aaq05I+hL2ot8BU29nFr4w4sv6s
4qt+TlzmvqJ7x2/pZHmXl0JLc/4BtYKHmwMLikTqWnrUZ9WmzyjnQTH1gVG2anWH
BdxkfIkkGQ2n4d8d8pdgC2tK067g4Rqgd796xs8zLmuSV2ceMP/WU7hJvxyiA21Y
P3aLePRcr4RasopV/PuZg+OfbvxfJTUM8AS0jfhlwj1t5ZoX5zqxJasaSySUIyqe
UhKmNFZlEXA6DathiAmKKVEi6VRrlbrFxhsIx4q/BiKSKeMIaKM8JTvjhPVGZUEz
4ho3mz5w+LBfjnwFBF54Q9bJYh2WN5rOsAly7hyyO2CNlHA3OCpGX+OcBYrnMA4d
iWnYZ1JQYhXhnfRmMc12+M7yN/sbX8e1RRGcRoE8KDNsI5WnLQdfHC5dwb/AFbi9
G51cn3apmROxg6VnoBhIa3P3tpzt90lUvKZnAod0UR8jQBbJzi7qYzmKPncxFvEq
G6/Kliv+N8+Qe+LKCQQ4fxEAfN1zybEw4xoH7qBtQKYbur9AI1Y8XicSM3sdCM9T
ffM7z9iRNA+cnLtd7ZL9+wId9vKKIJn3uhc3NK9h1oHrQHLsqXNbGMg7z6O2crBb
wHALZ3skw+xS0PMlclWjsOOmrJIznyVDBbnKJ4EWqE/xgZ++YF3eQSKPO54R1Ji/
LRhnb42eUxO/oz2BAGpzy3MzWU7+Xgw1V2Rxg4oPeBLqXOgCzw6lbOgQu5nNkkQL
q63xOubyFwNoAZDy9E0ujuGENg8HatiolGMueA3of5tCoM30R+3JPyoYuURrugIu
UKy21q91Y0vcmr+d35sTqkB1y2mjK86K2ZB+SwzdEGg47p6iGVge2I41Syv9bw+1
SmUcC6MHI2tY5tQL6XInVPa3J7Qx/gVRd56fdxM57DqjKRMPFgD39cenMbf3XHfo
qvsMx44WRWaPW5tdNLwH0nVwEEwLwAC3C95bhF89uajHPHsjMKdL3gns9etA+H1Z
iMWyX1iNjoCNZAD1jzbgdvwRUhTi1wEIxaTguWkUoLfL8+AT8eGwIvzJPVGS7AYc
vLNNqQ2F5dKePWTENclhpiEd28Xcr9rqJvbrit0cietfgfrmE9OhYBsevZ3rdPru
8fntQ7/tuNxXeDulEV3yjKIiGX94AV/eK/vRaI1fKXFRqZQ9zTLmn/Qh+M7KBuqp
MCx5sdway+5iio3//PzoZGcujVLcjMofhfk07lsIcp4PKB4K5pvHmXsEZPWwPv0H
WdUUoOd2Xj8briwoTgXfS/jtHDUaPqcsX5TQM8Rh/TbLnzTjaPDUpI8Hptnqtwqa
gqFmfulAlnnh5feTbV6Cun8MXsNW42wj6Qf/qbi6QfkCzpCo+ggrV+HJvtgChl5T
AEWQpKkp05uOOco4wL5cj+35sRtBWlFDMm5af2ejcRhvQhgAyJCPxLHRheDftR2z
tqaJ6O9Vnmtyye+RYc3ucRu/FW3wJVfHp85WbbhghmGsEvWc1tNRUmmjaIQYZtmw
7RQYwY3UZ6WiTfDZcm8lNkMNdHtC6+YxnGAA4zOGmRA4wE0HiMgw76diq3Vc/8JW
8KDAXPc2T/iU2Boq+JZfCXkdWFcVpCssbu7ZqeR/YFI/ZB0q9LmvCPG+XpNectX+
PoaG2BEVHXLNd+Syc+vm/Xqe8G1d8pktcUEkRr/7eTDZqdWTbLYma52i+GAqoMzm
RsErxqtKKNCZeOGIpJWnLYbc48gBSW7Y+5kfqAtOE2b9dQJi9/ttSfdsWypKPdB0
RXAby1rALIXUm24CkyRj5GJtv9TXCesndkYVGxCpbrhaVLokyF1XsaIQqy8EoDJh
ddmbPrh9Lsi2afqJhYIsD+F6hACwe52X1tqqhpHCTFMD/NTfq8pPcYAHgVsvvbdT
icQre6k8dQGTl6EGX/bz5j8NqQi8e+zRW0pC9guN7v2Sm3/w4T6LqHxZdGWV3Ljj
qpybWB/EWghxPx58f9CGKVGSSwWblG6gUSBafMQgqJG5FbyBRzyATcnoEQsZfDEx
Oc5nf/6ATVOOw3z95e7tr4FFts9PPH3ibknts74H9hvIlD+U1J8YWoJq/03+TtCS
Qw7TzwXkKL9a35pate1KiCEzuuESVCFtxkO8ze7uhm19tJOWKKp9XitACm3Aeazs
xOP77TF+d4myq8NFur6CYynqWKX/dDM7Xpri8RN/CArSF2oHDOp1DWY+26thqTWy
ihSXZlx8jAldNFTb4Qi2P6e0nC5SGDeWKnAZxZ3KpB1LwHenPOuCq4GpKqBt58zq
BdJKkPVcU1TI5t59bjNEq1tWix+93pO1czlJYQShfxdOpZgbli7Q5KeT8geoHqPV
ySCjTzNPzzzCQOf01/kyUgOxxLZRguUmdcumILX5LT9jcEfoNfSgR680N00SfA89
sJ83HHT0UZ6VthP/pkSG1RCc1LWdlIyXImJGrFV7kcyojAyX79wYSvT90LhEbQrp
r/IkM1cLOfod/INu0J60pDqrmAQcyR7fds2hhKpGbwIpvPV/NBnQjTKY8wYOC94W
luyALAshsPJBmfC3tOzE/WoFakTnCN6prh214LgdjYAiSOTX2COcjBVDGQVd0yQg
UWICOkHb2p07ZSOdOaYxZ5Fm5cAX6/girhFrZXgBTj4J/MLzquXU0XTzVnPMSK+w
gR+0+J609Cr4qvFG6GR8cwFLd1qHNj6bBanDy7L6D/wHKPuG8YcU1ApYctXOi4eq
SxEFVmO795uB6PYD7sfTTtOENg9m3Ub2GpFfpNgt/qJ7fqqKyU5WA7jcdaD6GaQZ
OeGB6WoLfWTbyMMsYH1mWri3UWXVZtrFYrn8XhB4V5YoZHmgEmcZDyksS7kzc2GW
TtlBoTOWVxjPZe03eyyd0iTOODaXg9IYNb+jHSamdk8KkRi0KN2TR+o2Tux8UzKz
7iJiwrFfEugVZLQPXBbN37OAhLpSb69ClV+cl6snKKgJPPeKD0lrJwXakxoBEQnQ
igKs+otk/wTYO0HGbZDj6bbfSa/IOyUTrNuQXBULgwS8uMofTEyf/oE6Bch3V8pa
vz3DHF3hRWfESKS4zYFY0PIeXmkQRwpbCaRhNEdkX5/LDr07iz0KZrdmaP6zP0Nr
gcuuI1qYqxurL0w7o8CAfnw6E8+cgqRsIP8AfKYMpby//4oviUTJUthutQbs9VB8
lA+9ZPD8xVdWh/0AwtrM49SEW8+/59KahO0hMyHxhRGxBr9bEpG+UBNsQmHX57h1
a7RJZyvxSQpVzq6Vh3q38aCg8WuFM1ila5E4cOesA5Qf6iOOjBKGMPHsQ/wc/bXb
1zgA2EdeC95IUEfS5r386mLyD2evhe+xFZMi8Rn0JmrdjJ1ePBqFU7ugJfPS7HN3
WhdHrJg41FmOtZhidwp0V8jY2evTVHEq3UzOpEyCIUFRP86y2RkCUZUYSG1OQTUv
z6MFDRrxy0LWos4Eyk+MZHY4U4Vj++/r2z7IeYt7Giudjx8SIGetz0KRsIX42bFh
0TwgylUTqfb2eS1AejvZJQn5/1WOm1Ggraivz4c9B0Du5EAHMPUWTmHHhOPptam3
gsGqrsjww2XLwd8K6Dca0zlZJQOd6pZJPgQr18AjzBz7racZ5oetiHBan+VsZh0/
F/1ZrRckwvt5wlWjiJ2EJYSstDpTBWWcxzbM047bT4jWi192EybNjCVpBQGfPoK8
9eYlriI3z/HsP500G7R+VvvZVkSHoQG6gme7UGnvoDqE1IATLS/Rx2fCo0PUG2uw
1IogD98NrsGd3i9eB/6+3F5yYv9cdGic8pMZlvKsYlcNtqGeCMJcx5MmaiuCjg1o
a5ASI8O20ROP4pCRApY6h2O3JnLHzMGlqQ2gGDDjNNML3aaO6hywdZg+QmSturoE
ilrUIBBnYAkh/5VQW0DN02rby+t8XvO5E8KGtx7sPjVSHR35HCI4HMBwjdhx2/GI
eomS9sbChXkOLcfovYX3cPnSoXQ/FHeiGTDo8fT0/OuMC7MLLWDObjSKx2AIEGwG
7I2/Am+kVxVV//zYdMqC9KRUuWQXaJEKpVS0pStOtGp4HKPxnybFzET9fFDDflDu
ciK9VUTx0CRcE3NLr/dDHmw8YZoe+t5o+fcWqr18G7RUiUlX9SpQBN/mRINyoNmI
GEiBNaiuBEAh0ljPTFma3ky4H5ts8DpRclFCKzWondxADDkkZPQGBWq+pBRJs9DK
oLiHDBxm9R8GDlthRKPoJsGx0XvXFrU2JekCSltBxLEEh1iYU0GvNAC6PjcqMxAN
tMrZbKK4GLy8JqQvv8QnQPec5Z8sadugOW1fgJrlPrWbcVDPrsMvb0SwSB3VZTCt
9rwzUUACWkisMLYG2HbNsM+4qtwXEh6DdnZKOLjyixi4WygIAM3QkpFUyGotpnLe
6sb9MmzPRoIXh5l9PFuQPnQRW3sqX/QjWWQ+GYtit+jVAbjasMxb+kxmXaEOnke+
mHrTdmsZ8ASaXyGb9io2oly51P8zLLw7Ykvc1kU9dbIRjp8V1YDJJortbIIQsKrG
2dSJP08oOchyvrIx21qzd0rj2jwjpM88fvRDg3++gk+WNR1GCYOkJDiGnU/JAPsd
0aJH8YRgBZUwbfDMxeiZ6L7+3C2CH4AIfxZtdAQL3GtUhifxavfxIzxX5HnV3ph9
llsKJJ5dB+86GEmHc19uwfQVcSR2eAqCIK0eaATojurwcYNR5hrO2wOJaO+LWyZE
9Z8KohIQrUvCM18OglHqTJYwQP2g7367naXZewJyuvU3HCDE68c4SRaXWwdO9M9z
/hb9fV5O0sj500uT5PDh3Ojq87u1295VAS9apw+rknnFlFlmmJ2Zh/rZpSXPJhn9
yz7zV2B5Jv189i8whM3FqWV2UxrBhcO00gRGqtykOcPVpCdbtq+eHWVB04nUJqgO
jAyGvCFgkT7TcrE+TS0YIFWW3sXNVVunM2p7hNmuN7Kc1gllO2P+7u41lt48lwib
6bUrTij1r9XC9bRULSd8bsAS5WF/VaNtL2+3WuhYlVHquGsiiplR5BAsqckjMpeM
9Www4MOW2y5C3Y4CjGMTJZ52fgPuc2KRjw4h9U2ADz2Som+pK7fVC9UfoesAbbGj
AKszGXRWeVI8GRpACyzcxaN8gk7NZI8BRZECJDk0DZB84LxU7I4Rl2tYJWfjXdwJ
ihrhZKRVieGw0UwwYllTqCArWMoCy9fWrhz2VwQD5Ukmaw2xek82PIVamW25LroH
SuUHQjfUP5P5RqjcdY+CcgRQt20CbrPmgOz2CXrVKzWv9CotQ7x/8CwGk4J7ZCYT
p2h0ivYnG79U4uLGdYL5K6EjEZ7hF920e/yKxfNBOIzHkEht4oUw18TSchS21wsR
jNjtmgEF3LKxvF+nYi1DXhKgsIquczwdtsNdwD7ILQT/1DgJ7Ncl4d40S54pcTUH
A4S5zKwaBhr8KI9nCNL/3EzQg8wiussOMDV1k9uOTHWjGyD/bIipTygHWfo2dESV
DmMWxvu8jrFXtmRpIQg4+YkeBBGnD2jQT7L63WAZ7x3gPmNMkhzwZm/MTE/sPQAG
ma0k+AJPxFzP8sU9W7Vox0wlSz8NbrGMS5qu7FSoTo5uUgEjDqU2Ulg+R0ObITJ2
HQrhWWiK+r9EXznrt5A+Z4A05MhXs579cYbaX3nRz6Lw4rR85JmRIiPhpgEs+qcO
2bAq4iOPMV2jwXiirfp0u5l8JfRSJheQEP8bB8aVFFl6CEX/gK8owU45/LZN9u9P
tD9Y4s3jN+2K+ycGZFc44M6MKmHAoI7gppQIxsufvrT+kfpzaGJy2GziUNjeBySm
ATLCT38g1EDuzuY7CrqdS54bltU/LhixyC2uCVXYFaYvUaJ8/xkezSwjrna9wiiU
IwsZGOYtun2PAVv2yRs/guE6BPd/g6d4K2+hxKu0FlOE247E4RvOgEvm6gkZnmOC
h0N+XPwMbeaZzPuMlFhlqHs7wvx40641QIc10XGc3dqOmj5rxdSCzlfvw7a80hfg
/j1wZjT+Wi24ASFR+CyLLmSjItYsfR+NOn2DK3K3gFAi71Ve5f7dEu4q4MN+DhYg
RICXXPwPSO7QxoLYa4PKWh8QyI2/QDQ4BaDspaOBkz/hLKIitIor0VLqoY7/xfGg
35NRVHBi4860MDWfqUe8NmCcpTXzDRloR/h83BXPO+cGKRsGOtHDCX80HBSaDZaL
mC3NNnJFQqIqwQ71LucnWe2czB9vaRx6rABZ5Xq4LHyV9cjEfuMHQlFcgcYwLMHr
krE86LKcz2CIclDVbfLnCjgcNsrIoVrbaQH/4ieKCxCD7j5mulbzq2Db+gjLlpfB
NYKrYo7+Fy0rJot/utxyy4oiPkN7k9unwTCtXfo7Wp6mtz2vwclnlmPSmVZpOWgb
cKK/vLaFw47DTy7fJ8wXvGMV/Hc7qhDYgOdKGrZExfzef0Fh3XOgfIpyTK2C6tZK
eqB6CuefgaozBQv+UsME6jdYBr2UWOlryl98JXkQ38YL5ql1T3cFBuT0PAkrgisB
Hn5X5azi+4l3TWaieVnYygwDIw4nwfBPqEYeM2xJI0KmrN7cxITfNCJGwxzlEcOy
w7om1cqlOAtVGkiNMM3Y9UsKNWevtR4nNxBitpVCMjSPHiUMfNyn5zcslXjzCTmp
OXhDi6GwPZz7CL/cEmHROTD8EGCIwBH4P2gdviltFtPYkGGT7ESCUjdlerlqcCFW
jleC0Kh5UnOeUpngXdNjzsLLOXZ1i6WIUHhcolX80DhEMBYOjCemhNm3oBb8Lwsu
fhqUjsdoZWcglTTG3iei8ZPKOI3YQ/aRuFU5m4n4XbGtNGqNMrNiW75drfjSlr1c
77Lewgeb9lWjfZJ9gATB2JW7xZQilnKepALIVtQEPH56WDYZYt7khVkX/geqNF82
L/H4aiqOZsparwAN7JDC54+0pJ5XNuE6oYvgEdQVwg+bU4HPtunLIm5uWmQTlDvY
WJPUHGSwuxUiayHqG6Ugy4wcCajuXtpEb179nNeBuMwPVYa7kYXFRc73xiAytvfi
UrbY9mTHGVdFPOhyFsY5dpno7VpSP9O5lUqjY8VSqkJPZ7LuTmPUmSJzhLTiV5mP
helLruxabQDPq6KwILa5Eu4mwieV3UmypD8hp5eF1/q+9faJC+VgL6r6z9EvqB4L
LJy13gZxacJILJzoxNqeyvTBjpszOH+Ea6fCx49PzxB8qhE0x1AiGseyLvqdoaAZ
O+8OH1JLdOCF+ja7J56Q/RDZELjCTqY+Vetx5fEiH06gsPSBrl7yHNDs36KhyjPw
1KZR0uEgAzOOT/WrkBc0rP5hcIbsujaxA/8udTgAFhMJxZ3bMl1Vrt47G6LJWuTz
QqEAiTlTZu/TMcUDyOLwNLfcXyLaWS2/dd0B+jwqUJvJ6I0wwHC48ybaIMaczl6p
Cwk3St+lECUHs6Jk2tgnSObilrTO7/Drn8ITGW2xOjf2Jn2T8ctaYIF3CYNVHIfd
RcMGn1myaufbxKur1S7uLRjmV+9DycxNp8FSe2xfAUTAQDm5lgudexy4Hj/ma1yw
GqOJ/oj+V8n5jbDdCZ6hSLcyR0+QFH5///SmiAfUuVLl2j1Q/TusIAvAtVfxZIUy
dEkuz27nw3lOqSWV0fz5BAARY/ex+zbnYx7qPg6PnwUfzdtRis84pdYwHK0gckWw
10LsIDyr57ezNClWyuUzPROwHoaTPYflyyY88m/ePtTfsjmhznsKmlTjjaFR59K2
lEFLbG9pRLIGmKls2aEddEb7DQjihD+E7N9K1XuArpEx+BVWZ/6Xq2FlQ5GPUD2X
prHTIDVco2TNMdKtqBRPSytjr2cHan4xqOxU+VLqe1R6Ffc5Hik74rDoCqXH0G9q
mAi/Fhj/L1Ny1KdXIQqO3kfK4KKZItzv7ex4sOiEwRWfsX+rR/il4li16kr6s4TH
w3WjM8GEnUTk68D+tJaEUg3Tb8twEO8yM53AbdlTyIcmPWIZyMpKeJWpUvI/qiSG
Kx7jvwhOlG8Cp3giv+C+OgjUYhkSElKKZuu6ROaHE9WC/AXdu53NmWsZQdgdt2sK
JLONo/jQkegsd5DJ2AaF9LiQzMr9vs3TGwUzE2LaBdR26KafVYp6JFZWytKPHNVh
5Kli66zGQJnab435VVcov6KoBrSDkazQEVYfUp/uimnpH+yJlvelXtPZsL6tWWLZ
eUgfxYOVGYdA+ZZz80GTFCyawYIkuM3WGwt/3PRPEcw2/H9fMD1VTr5RTHQU76np
ltm1hjcme6xtL2D7Mv1NcE8XaTEtiSkhXaLe0cPnxIwli2CwoRJjoRBMqzdgiGdS
tZUh7tuQfyFyKfEbc824lZpF86sd7IE93uwNFXj3317khz7szuEn7xM/vnbHC5HA
o2nTb4OYntzfomP2fJZnxSJfVvktzyxdJ7pv1Q/IcO98qR+WAPZmFlqpZhXIu0e+
xmcCGg+69ZdKticEvSidXkatpu/GZWRwurz0tvY3dQKrpmnEdGqQD+tvDF0OICnF
FxYP6l9V/DztX5Fp5wvKMpOSliIPrHpFo0jyooP8VlRhNnVZkj7pZfTOUZ1rS8Ch
m5SIWs3CEHpQAJLnwH+hiRBY7v1LgyJ1Dze5Oon1aq7lukEAJ8BeonBJ2a8xBIK7
leu61o6Lw9Q+N+kzoR+B3Snc/M9+D9DqYT+YNsdF8KRlYBReBLPptZTbp2SG+mMC
WTMommkF03eaKVMyL1gCPMfMMBThtL10/TxgBUqB5WvSbmCGRC5ydk8Kmj+L0/XY
Zcw2fjanTzXc6n+EbJF8D2DHQ76lKLcc8LaaxQVykZ/VZ0hRSDEK9PMk+oWWjPoK
gZWAVEwRJjZfuSo/E7irC6/UCbT7PN81WWT6reEAicdH6RTJBOqv7ZGxAzhE98Ol
gMIgp4m9QN1wFO94BcVfgP9X16Q2h3pXqF8/mGamMOE38qFGMG0GeP5D0Gro3TqV
dFni7Yxq3LljY5t4lk4vY9smSfkAQf3n4ks7tiRDu9ueaNVVU3+Tj9A2AsNMypdH
95PbYPShwJ0M+Np+VVlgolR+qTqVJTPgYZYxoAGUsk7ibeFqIBlZv4kCgm9idxO0
mVFES2LozQ84CjwgnuHYyU1WwfiGa23Om4ZUcXo4sxVPgRU9xQUGsFPaSkdtMywK
LM51sDtXk2BcJcZASRYRVtSrrjmLPpPTik/vA0/COkfBQAQhKSKs4W2gcGlpmTQx
Laz6/nTDwufJ+zj0pP8XEp1lX1l4ZHssI/Ul2T45X5OUv4MMV05HzD22Ly9zZeyG
EWs1rmkdXTNr1aXF9VpmT2YXjd7fVP6dOytK9gIjsn/ZhUFwW2QSGrZIGvmkmtG6
b9C39D82GGUurt9m8C37Cq/C+HVfXoWPfqybmwusnnASoq/Yj6e7jLcoNa+i0mMf
ivcGrOFMABFXxqH/i/k9X6zu8xCiVDw7HJBksVwm5RNo+LPl4+/bkWTeXnbdeVhK
1Xyqsf+x9MgKNrXU/A5dKqCiLuertnlU1ue9EPg20T88Sgpy8VLijt0vX/Zzrt6w
CRtbsSoVb4IL4GoQuMym/nvFh3XtZU0oFnoos09icfPpztb3/5WrouYjWpAEpRoU
VZdTsKWFJhXYrTE+XTnRNgEAVK9Nht65LYGH+oSCiA2LQ6aiYyD7UT4kSu3Mtmb1
sWN+R9LPMlOcFaG8RZwjCG/LjUF2jU1TSg1spd7Z2KKRcqDGI2A7JJlFTVOfsCqj
Y3SBoubYfxZCRDhcczPTQA2TS+DzOYskucZkBqFV01fJBapaBCN1r2UOWq0zcKnQ
QaocN9ie5C6+RG29c8J61dKPImv+R9zIuVRMEgbNKd/0hWkb9wro076MJyuHbZ2g
L9ulLeHTRnTNPjXCQxs3dQi1nE6DhT6561Z3mPfN1XOevA3hKa7acKl+1atMbfav
oqW+HrV8JancRMUvFPN65rWl2ZKbbAz3vN3fQMyR9kzFBvTKPEZAZSgxr0ptxaqR
mf325+R50C1nwjxoj2MsoGl3IVDFvYyT95NgBBmdFaKjxkME+RDVqjFrPwQjo/Rl
eAuBGBAc2lpcTjcOGO091qG6msVDWBpD/JViXsgxydDqcz0COny8XlJRw3MSDy5d
JfiVroANbgKqowU9y3ZRKsFcdWSZY+dSeuLMDlH/AfiJXJS6miVhoVHbfkdjRAV1
2FvrcjMGbPCA/y49WQBZgqYSev86w5U3Iltf03+QMgiNWn4wl5kiz596/ewKNpmu
hle+dt7pZc4zk44LxViDTt9VFvOyK3yyLJqzggLKPzXocr2PMy/K3cc9COH3hXHm
0kEq3Y9LTMwi5LrAq3R82SG/E+LesxFO48bWxwgOx4ISbf0pYLajm9LzC0ol1Kfb
dQfIcEldVTT5GRSid+L7F9GmP0bGg4l9I2mDkG13zQoQbPiA2RFTaZSGfXts265i
UM9dXIL1yL0qzsWC+QjDM8HIn22EvG3VxPeLf4gEMq6jAR5xi9cnPyZ2QVys8EJT
Wh2KTEXlwQF3DwKkM0vIA8B4QysI6q2LwGpg17Zkovo4317XXbJUgRXQ04ad6DPe
M985d9Xx5REsm7Ms+srT0s+S3MDueFHepfdi6q8LkSffqwyoKNOTsKVK3Ryz5yGU
wWULclqup08BgA++ihieT4QWcCCoEMVtFyBMzUVx2M5iIB7512M4hwgQM50Fnd/S
OVUXQoXBNmtXumNSONUt49jBcnxrv+Lh3Ukqa/uuojm0TySKGXoM5nCNvXtg4ap3
34/0I9vMk7yKeJb+yZaj0q8s8Uc6uUWM4/m5RbZ7ro/5J/m49gccOVWzBr5+ftF9
2FXpdCEtf3QSWOeLzfQjgalRqGZXl+U/4ExuxF5fgR/4xRiQas7E0KWSIOwOr4PG
vn/4HEV3n8WEV2Oc9qvqGSCd5qbx8CKzr3PzS6pOIm0r8ptMq1jVkTsheVOjEjAf
6yR238r3y9npEQCyNIxDzMYlYFoDTRnL6n2BwadPOLypbsSigIO68SrmCi6ExqOD
ahaETyuZYH9jy9SllTAzIEUResEbtgwzfgr7NqPgxOMC5PyNozmIJEsPGgW+ftzE
qOW2eY4fJ6gfjgHQkWU+iEVxHd4DJruzj087IooIZkMOJJOAMpV2SMtq1o+QtCvH
/562Sk72+0eEuxd0YV9wmfT6XCR2w1DeWSbXd9+3AeW1EAbCra8afUSUoj84DdMm
e6WYRcgwJIqlRzE9eVmpZ7F08vCMM7vDX3ccn9Jdc7HN1a3PpHmywS0M4yuRmUx1
dOhsk+CjYNm1h8bSqsp9j+wfYfJTygriCC9/hAVyPd8mHztbQ9510D+zoAujA3RK
/j8PZFZVJv8ImkT9H9cHE/9/i6DjNLmO94p2pp9A//9nzZ1RYf9eB6LekVnYOQri
cSjkEDsAES/DkJMRQryxx59UyyyVvPgAPSiFjpUeNgVkYRBfDrrJH/qm2qaCH5De
/Bqq/9Zw70maFkAVxiE6NhjJrtVVoUtDfnOw2zUYVNndi9wqxQJD3FCG+otbEyUZ
EMYAvPBDtG53k7NIGiHd7IoApdbOmU5aWEmbUGkrfUritDo6lYkwf/JOobFY7zlT
avrYT+4OJt0Ae1umIHoO3wOaaW+hnp6vHbL9TI5PGa1ThO71wj6Bz32N99Wj4bYt
LVeiDJF3zDH44Wae/9ko/7uSDQ6LStnwr35Asrw0h5XZEMCScLohCjO3nL0A9mJR
TsU5kpPLm+gMzpimm6kjOH1CDQhmN3Nc+VUY5ykosOCZqUf0VrGBqXS5gL6M2DaE
bvnBavBQWT6+61yr+nNAnUfXzWaicP9zdkGFaz8JqGbY+jQYpG51gYq11OE+FD/+
RJ9U5LINkDaS1u4WAC7sWljc3HAvwfWpfY5JOxVzfdDIzjkzMXrc21Wp6+0sYCmI
ZrngiJZrtTCnBf6GtKlxS/GOGRSg/00KQwVAOq3SJgorTu3Fz8YiaXzrNnRCGV+G
DfqxiZwX9B2eiE7AqeIcOoU1zZlF4N5JliOay3Lb2r7gBLZanZ3NrO1I515tWY61
j1EXNqJrtLjBSBsDYqxIFsTsK+x0FFOhn2RswuPvhIgA6wdlO7a//tgMyexQVezd
ZpJtUmU/8Gww0NYIykJZk2jAMneLIFAu8DinSQLZVX/754jEh2BlSrG/0QZXelY+
cR01DLxE0yU5T/G5t7dtmUf4Z4QLkf4ukxXnhz4PHNN4X3elWE2m03Zn//3lXCkR
9xtBwGuUsrgB4r+zKo1AkXSF69eXjOS6ZCIBNete8/OrNI6cHQmZmUM6olrV1FWV
DtG+DXnclGJaMrwaxuvkq+SYCR8IAPY+12nAUF3W49urZBOqG64k79z2Aox0uP3E
KT5I87ZjGB+1oMRT4/J3e42PPNH70Cu3S7VNl/ZeNizYYw0Pp9p0L6/4DJacq/qV
oxEzhEJZYPAtMP1rzTjtKNjxTAofbzSnrIsuSYlkpZdCyjBpVl6kVi4M4e0ANTJH
mlLjn3KaOOaTIdh6v40qjo5jMKKvaewV+aMCrKJzTWbe5XsnM2ZL0dGHkVx1pn/C
E1huQl2eQgK92E8XPO2BEj88YKVRcmguCG+Qwuj7GNaTwcCZjS/9oULive+NYmHL
RkGzfisvWb0ySoIweyXGJ4Pw48gA5S/ETODIwTgwVr8J/1vlwaf7NH5e/CiOoMd9
qfB/X85EEgEwEDouHlMvp9yrgLQPpvQNWGoyxXqZ8pUC7DFKyV7b1aX2SGbmzAyQ
ykD8Fyf3DM0vxQwsHumYsPVBvKIS4sy3NmNF+giWTw0FkAInG24vSNs/U92ylXQs
TrZ1eJwSjWtdXgUHtk84g6N0xyIFvx5EcD5+LSgq47TM7yi4+ZP6Yv/wbLY1LUfK
P1rSSt2i8iK5X33P2h0bmDFbwy3k3ZWnwxgVqK13khe56koKEBmQW2XLfrg9pDNx
e8cOxTB1fHdc+ssAZoCPVZWMdyIyhkIeOxZ/J3HYFOLm0Wv+SSI0DCSFrcAyavip
3SBLorbXP8H0a7BoSrDIjeG1dbVinTvewlDm3F1TWdOITlxa9lpYR7STmefubFyQ
LGSP8R4L5ojQM8hvbeQwnC4zJT50wB7lEDSY1unXOGIZ+Wno6K7NzjUjN/Lo1NXM
bEO2V9YHSLD/ayxoLl19JZ27+KYx3oOwOiVmDoAIV5WUOoE6QMlB5g08UAcVpQbw
6mFPBh1LR4dMI+l2wYmEpSDhpGfYKZJCTmYDXTopLUdrq+f4ylhsUxMWU8ZOf6Ug
m+7oO1rfd6uINj+F4aJMENpiAd2l8GCxki2IsMPy5pbZNQgf7aigCK02LXAGCGK7
cw+TvSE1r1/gWy0Mz0V0cXR5sHbOgUx0VUBP06tiKBVYRmW4eLI3qGtyN23cgRli
Pd4I6uzYAyTVWmMXxn+yjMCgVApa0MvcwuQ6jajBaLpU05uWoldC4/8lgH2gMbF7
hxMlh5OGLUB/wccaf45BmzQY4AK2STUr2qwxi8UZhTtKdP7indkX0DgECUoXArPB
ivezd13jmeIbqco+ap7NXeUyFmkpmhK5uzct1399UooqowAMndOF1F3oB4TUXbtf
7BX9OuEvmwFdkLZLxgglWprsm9rttmZxfJYyXIG6bMkrPyyxS9yxj8z+utn42iJM
sVGNEqh1j7J4xy9lGWGvE7cgj0xuL8/eYxV3Uvxqw4e5daAgjjdUxQb7K8Jl2WZs
ZM9XsI9jMWKiQs5a4knccIgQHaHQ8Lt+gjEmOJ/NJgHD0eB2UOwhuHtlq41HhEla
CS156bBNxkuuRgY1CcfAdZG2BJctr6QnAG7qtKNELj723Y2Ir3ikjhFCeGMfnY2C
LKitbyCORCb+kFQkAwBe5hY8eLDqzvnZ+O0SSdG8rK96stt8u1V6bWKOEuXNdOXc
QbwY6zKAoJWLObcju3A9N/K9qKH7HGAQCpTlA7u+dHVHMUjSECGz49CJzqBYhNk1
Qin7Io5Hl09pDIxXyIwE6Zok9fJIToP+YqyS8Zjdr6gjnLX8zQtf/EvrZgsEcnXD
u4om3YTbvcbmxJ3WioE/N+sMulN694BUO0+cnZk3XX9wXoQaWHmpD3ShZw5GMvLo
XSnIl+pFhdH//bMRxWsNrbSi9Qia06knVs79tqePQG48eT6yqodDbNIzXPu4g2R1
eiVnOyEhMimdiny37XdZCle4OXyiq0XozpEp/Bu8HlCoFW/V1lc4+b3mMzlgkUtL
6ar/MNcvl0ZevBDutGIn7sKYrZBbFCxEefxoYbwc+c0dl020dkDnkMf3qQScwZoi
mXr4fKUpveXiT7IwMnLUyKHwBb0suqRmw3ZkFIqsUjGAOB0r+Er50EGlkI4NYaWg
FroY8J9vE6hRCzh5ZNyYLiK14DrPr201gaTxgGuUTZoWwv7NnXCijBgCwVKj/QOI
MC56vKZh1r4vJEuqZTsASMdvbNwksG8mAIAd731nFmm5lo3BSFpgDcl76OvjfgH1
1a2JcJlCKmkR4bJ0glgMIKyPEyD+PCvVfTEhuTdnFMHRG5ZTAoK0K/YfQ7nqSEZO
l1XOdaU3r8RbQPuFeTSJ5B1/cvYcvShXWC8ZpBl4l/WA62T4MTTaeomPsChYdYZq
Ykoz6Ggk2VClbBNbe6A/YPXLWs+sf9aKoWfcU8QJkOMe/2OUVPjFWOlqxR6YZpvs
9FYayBEVodZ/KJClR1Mf8YYUFCzdwZOde8nZ8aRs717l4RHK+hL5eOpINpE28dCH
a36L4P0Wv92RrzAAo7nyin349mIf91xRPKtjibbiv+UoHnx6zVwU79AmexKLIhFq
AqJ8mTuRkXWZD9VHY8AEphsQ2VzPM0WOlJs5j0f1EGTIW1heMz4TAn2fRw+lVa5J
Hx/sDPJPZwBCMufwa3Wdn2AgWTUD9s07w/XoSXv3ddExFQbcIfmbP1jiBeW4ThBT
q1wUrqMhLHsKUz5FjcF1lObbK6Ay4pWxBJrmZbn/D6KVnicLiNNMQAUUxDBmdjEp
RQo97d49bdX94xkLel5+9X8kSyIXD82rd1RcwTtaNl/yaI2yiQ4kEiAHdnMUlzM6
N1ukwzl5MFpgCHlH1hYQEFXjKQoa7eA3ZwR1sqcpRetvFJ7hnVl+7VsWM8fhYkoB
YjSpO+t+haBH3eAyqIziWNiVMeuFf46q7MFeG0uhtF8lkgFR3eQ4qT+1ap10khDC
HPi6EhrR+acG9zI8aIzovE5pro3p/tDXV63yJgjrfSBCzzpqvhnvDt/ghcBnHwZ3
xKohiIC15mY1I/o4oQ/YhsCgXr83PaNZMxWdVFMJ0KWskw4tTo5ryWBycsDhRY+W
vqs5YbN31GucTP/jnbhdN37Q0BwSDMOEzgBvVuS6i9sP6j/0SxZOv4XGYm8qSHiX
I3ukCHzCLYP1DYanCCTizJ/eT4aL3PuFGUUzijWBhoHbNnlvV/QD/NF7GaryTgVg
DAE+QrjDi+wdA/rnxuLx3OyNJMbiyZnHEtruEzP39nKk1rGy516sx/c+RbB3VwJF
9iZwEQDVg0R10Foqzyne9JUfZPkEANcAGJuAghjym4m35bEJqu+YlG6x/wpVh0UV
wGidacmpx0IVFQx68SKzoZmxcxETTsBfB/PFY/dHmILY1d+D5Z9n1i6gvrNt5xIh
cIwihBIZZg+SIkEoGsGix6eKpUFH1uIqXsUdt+OluUSQ10z6DmSXLnMx1F4FmoME
zPd8N8XpMmAk+UoeHbT6sbAuFVHetXUeqg3c+89GRyu0gMTPb8Kc0K8d48d9mqN6
qPpatEQFE+NUrWJ5WzZ2pE4SQQ22vxNO+ZUOppuXDYfDRlO5CJhLFD2ND/pFSyDj
k6EARWW/IL+Lq9mAUIOuuWGneBa+MIEt1L6QqSYxAuOMWz6GopUUHTYk6BWUpHaR
mzB3cj0zc6rTEInCE0p9zk6BSK3xlnGiwRvqzuQPG8xL1Xo46nqh3V7YZnFHRtTP
NgAAF+sFtUwUhPe0+iv3QavybXJ/QkF8DUEewxEga0G4qgBu6VDLxXgFmsE0W/oD
sBz9MbnHeI/JYRjeXUu1FDYPid9vCddCUP2Y/UJ+OFGPsth5VG8fOjxACRXlxWgo
ydL17xuI9kk/igs68ZSewsvSD473hCJGwaJsfNGwro/WPE6R2mZ2fb1Xe/L38AjH
IQDrG27o7WbRPxzl9y1mU+r75qLm5/OCarkkEdMez4v2K5rWkPd4lLXSNYMOvb9c
DdFXWzmA66oeL475X8QagtKX6nwb/mikLRFInQQf1lUlSuo51sUMrJl+T+f4jLKv
VsVk4I76iGcFra1g+bp4kgA3dsFHFHPTehPPdkFz4vRwaMCxjbzW4LMfYlqPSeIe
57ZqF+fAvkamH4BbQsx4PIUu21sI423dgHZP+yZ24zQbSd6UzLjlySbW4kiZonlM
CPYZb9D1W6jSOdm+71eyl0827mVPFLNYWfj1FefpohkPePJ7eRgqpsLS/zDg3il6
FYozOZZ37QykGnSQTs6gt0a5mjS1TNg/6lsf/qG3mjho81U/Td1XSt6ThzEeFK7r
79iW3HzV7QmdfioIpXxjwH7Zv3fskUUIlkR27b4VfTWCHLDDBG4PLairJ70IZ6dY
EJJfOaXPT3CBQtOoD6swfDgkPNheVJ6Hn+vwTSRH4LV9kVbZmawtthcWl/Cejqi9
pFhxFvH3iofm9Gawl1FhcmPnlKABSqp6doNqDa2RJpddh7dYhx9Gke+7z0yYt8YS
999lqPU3twRIUJcpi/Zs2/CusB4qHICi1OmNBeompHbI0Akw+sqE3AaSkGtXajPS
q1ZpJ6sOBmqIkUdY6NsqsfxH8pus6Z5ItzdIt8iZEUZVxo0bO64IoyHoAMJG/AXz
QdRmI9rZ0LIPs6i9pJq6aKSrf//c8o+sgwG6qiM8QnS/y5DtjhmfIg/RyAcW25mZ
na+2l9aGraB0dRT7WLZThCqKdNFEgEpUQKZVxb3JsgdQRbWUhCpG/z6pwvMhlZy3
7iHf7uZdHpwnwlhSbD529e4BRx7rdUL5MjeMReMSy5ZjuuQVEmr3kLXmW+nAq8qF
A8kK1t1SxOWhL9PRUYYT37FsbLJLJyzo4hEQEL8ctiWhmxfM8ja1e7kyeLcDKHgF
C0ZsVwyvMef1b0nTFTPzg6Myo7/cOjkZSNAtSAXEHDlSbCwUfPaCbRbP69NpWO6r
Fw+C6AUU6B1CVLizPY+yW+YYpOG/11HqDrXAIEQSgA/tpnJ7HW5RVEGAJSnhGsy6
vv4Denr5lCK2pf/TuXS4fVVILIwcIsNcn58vA1u89jVQ3GtbRo/0BIyR8adVHX1S
5NN3ielORlPyvIyp3bDElaY7k/yvAYdeqNOOzCinjArNudI2fi6xWz5qd/XkSAon
0vPTNDk5QdaxIzlfc7Nqzu4Bp3L1slIeLw5vdZP5o0MlM9nKHsxhg23ezoTJbH0I
gJuezVsOdoo3gNkQhc8peiISKDeLJvEQ3m0dGhxvSFlYIKGzx3OjuBQBu/nUSNSY
iKNlRFHKCiz/XAhsJbecmEXT4FgfnowD41InlmPAJgJsa53zgwCDWv7Gp6Zq0gTf
9ysVNy+f1TTDihDlfX19dJw0o+KKpmetwSKVNTSHm3tFeHq7YMeSBmlj5dhDSXt0
gn/7br1ToszCcDgYrBKdNRUubn76TTisB6aufprmCvY8/CZv0ooUVB/q3Eug9+Wd
p8ckfRz5ygT4rD/IJ52g6hBDDqQuF2HwmrEO37eum/itKQoOYXmOKUCXpgmW2U3c
Cb0AcaRw3iO9RD0nxWp/nLtwH6W5X53JdgLk3gMdQ+v6XaivpD9Lpqjicp5grW8K
0TbtCqBzQxCOapNaFV9axDbukN5vsId6joQIw01Pv9yHAcCtoiy19DBziiTbOFnB
NS1lu7h2nov+wREIjYGUX6zXA79tfkO8+k1MtZR9BlXdU5rYa0/Outyj0M8wlyzV
fIxYumBkLWrEp1aKxhRSrA05hJ4wMDbEFQqZLVaC6QWThSKRaywXbYFh5cBfn0iC
/EKHa8pV2tsGdCZn4mYImNip4AFApuuq30RWxivDuqKF+aqZWH93KHPow7Dh9VAS
RtKw592UNKhulO42bnocODHrc2C8Llk+w4cVY9mGl25LQLvvL/fMkgXBEp1w6t3r
1iHXDqs6iCAG07Q9aCxnqu1UHYIk1SMuhqRIvYSOK9XJwENEX0yCu5sQxMhg7A5I
AhndGp8lVfKgKeb3klVgsYnyI4R7LEOc/aRyIeu295f/iMck2cJexT8ubBYPL3ZZ
7tytSr2PMaKaQoITHdPosZJjE+wnFJ3FWuxhZLBCLyGFJ9d8ecxzhXl0qApCm0dO
SAbckQuwh7YluGcn7iiXkPuZA0bstlS2IYdANUz07+dT3QwmSc323fuXNSjTWsPB
09Cb3S8XY3u1DackSxixoMzNdhjPalW2VxLUKTvCzLPqdQjco2NgksHJY5O7IO3C
LY5k0bHd2zyJTfpKFXEjsbVN8wrOyam1QXr0m5Bvwq9USR3DjJ8erz757+NaHPYV
IlNJpCYpDr6bTj0gW79m4D13hu5SA0fvQseFDlj19dBqtbWspx4UbECShxULs5I1
gVNg8JsCAoUmrcgFvQX+RFkyvQbxeM1Dr/4uurBVoL5Yye+whV+BoZC93l1ld8C4
JYKwJkkI3KI9BFCifNr6Qw0KdRFJI7bd1UEgo+IggDew+LfgPMlJgaycOc4F2WnL
LgpaMKeMfTKW14ZSVnJRJ7Uebu/QEVj4d59JgEx0pigkUrbxCwGwG4KOuXySFIUn
a8LTkX5tIls3PUIDSRwnzMQ1c+mRGQe0bzHG8qv7bc/p8DJ9YkFkhWUvatMS/WoP
4zPNq4lroZz4wbaCqeyn5f05pWJ6AsSDM7+xBL756gSE5wHFz6b8+ROtSZKBV7Dn
UtcMDcZ0Ff19GHCh7TKlW7SDRw/1EvEVzf7akOiolstAlrlm93OK7BqnRwj42s47
E/9pP+dsz5rszVLCyFXQkyFnwX7oGEXUKsIKnLhNqOxjJcaiQ6c2oeXWdlFOKFAT
T6rj0PMgZNW24NwFEL+HmaE4YZRM1L+Aius2gq8GmJut6bEN34uCJAjr4y28WoPv
ym3IMaoHido7203te7pAXOX2TGXBy92ycFaP3ve4eHhtux/lFIAK5rG9rDAym8OE
OGDYiV7d9+beDWfvSgvoFZXeJIUlqwX2smtYk9x+2vre5Nsyjs+M032FYDJVhJXu
MQsBxjymxAeWyOztSoq3WijU9tDgyeg6OaDKFamw0LAbaa6cGDMPV8h2C60B7msv
7E0sJmZimmnH8t2zfFveidcDo6IphvJM5KIXVr99JkumwJZp6GCpqCy0mgqn3yGT
u3SUcCqJe4iyHWALlSZlZhTuGIScm2M7fxUGEjMe9xs7YlEfqcz8Oh32y5JsE0kJ
OY0fz7nOsniK9xmNgoPj1LSpCmwv19b4cpAtMxfFnTgt4n/SO44BW5+OrxIACKru
Uoy/Rf8w+7n9y/z76yYeeBeMfX2uV6TBJEmZsasHHM937CLdWImoQkHV7q2+Sq9t
AQB+n0B21glsc+91mDjkUbhZRNlLjqbnmBIZVZK3GmxM+VepeXoQI23rTxq0gR5k
kH/05erPrnPQdKsTnNBRH2ydFEqHEejxWhshlcU1DU7qup21Zr+H8nt8YXbeHV7K
LUnw8OMarf0S7TXkDk0gC4ELaMc0x0mc8YtR3zX9qtJmgQSszp5vMd10njR54wDU
pLD7l1z7WghuwTTe22nn/hQ/QQ22a5x66I6M8GcWeUQAy6CArYRAWJ1J8ul4xmsv
gcz0sHWAUwuzuhWhS8DkpDqq9cGb/hgnUYZzCY7NxVTDwbuqxkn3OIwdztCowDMt
cBFUnITFCE46NjF0qLtCfilVJPsXbN9HcZl0EF036cVKd521bFTkfCIn4Kldym+4
Hu5cQelF27mejjzUiBrvHRR691OVEnj6l0m2Navd043fxyJfdUmp0TKuA3bZ6VQy
KKGzG2DWwOT1+y1/yy0AN0VkYB7907iePa4Bc8YDwnKnnhdRI3ZmRc5iHVTjFXSE
0iThhEPSAC3z11TgWCL+EWkGExUOmrYe6+i/yo5+LCE7uGawEvrTGZaOE90oQ8o1
wf0DdGxHOGdFGSyIwSWHlPxzWTDRDjEFR0hBH7gIzPeyE18wQmVI5ZN1CskwPH1z
jFGTxEy3+70YnIdyl2OhqIem2zneKiyrSCl7EisYpzG0/04/IoVNGESBPuRCtnk6
yQJJth3zWZEc2KYM2zvlUEhPcXE9yx7I6b1N9DEAUHFIyc+Q5rlxl2ccUWqL9O+I
Av+R4WrCNvkUsBIqRVp5Z7J+UohD53bOytBxvpC50KclrzBpIiB6xP1OjUgFbZLW
1bh8HPbH8m0KnLJ7t1wD0mO0JNBiH9ePd8xqRhGBcrVgrP8X67h4/hnY5Z283G7s
c2z6l6obja20AxGyaUKwjCjMT0feOGDcPs8W/rS3c8LXQUim5XL+PmTIR2KWRU5F
cqaTdfz9XN1jdZYj6FyxhhXpaisMeVDq539iPIXsT0YZn3QP8tPZFV2ZH07QqqpY
Kjs/YTMpD/I9tp7nThy5zG1SfLsPtjJ4Q7h8GnXMtYk7qSxbGX9nsZWzg6i5joy0
t1e398SQXtg1ccsIi0hwz8F5DruaH7YWO7KuUYo6YWbojE7DUagSLyIqESKotUAp
5KZ86TucAGGjJd7A8bczPVBXXf4PiN0Zw0iZqYFcoE9VPqKZ7RQLwakau46S4gnH
S3Tfc6YD5LiPW1w/SNrahrcl7nsqEGHW7E9KWxXFI1V1iNrxK2+pFukASzAzeofZ
1xKipJdVtSptGgra8sDq3kA8zSyMHEOFmEZfOozwqg+pMa2s+QfNcpVIgjdpUtm8
bjH2beRiAj01k1XsYHGJzBm3HS4MVMY7+LZ4koYvjq63NXvspmPHdoD1TID7fPYv
cQXwsk18aND786TTZjEolz7MnrfEhFRuxueMMr3XnCsh085Ym32Wv1RnHAEJOwFU
/2GoJVDwXrMknGlhNUrFI9D6AQxFp7YGZ3A8Lyrvi80hTNjs6omHtI6s4uT+smKj
diZtbQ9SFgTU31R6eIkPsfy5fgtcwDMfMM3yT5I4010zboqODkTqBvsdZd65YCPw
oW0OqFSxmzekBiSnECwTsNlLO0tYGOTZL9o3j5chBMOdI/DbGe57SylxLYT+eXtC
eKdIWb66eyBGbHqBvMmrf8pjCOFYV54Xr6gGefhVnxPqhgf7PYHM5OPO53TX7u/K
084fx/qTZbGJIc2/orRjJF9qlxFcsU+kWycEhUKE1AkNczqA3Z/8Hdo80057mFKn
wtVGhtVH1dHBT8lg6PdjaAUeLS2ZonvKNN42spwcK2wL2+wHIinUw4GrS11EPpqG
a4L3y3u29Dx+cAHhxDoOvvqBrUQLx+N7GuWEijxk+k8xMC3DHS9cU/Lv/wEqWoYk
B3prV3mW8AqqWlCt8hIgbeAQe1auwxmjGQjMPQnFGvjLpHctGCJnwgDYjqZUgGTA
Q0IcVgiCgV7DRTbFFwVoTAbYtuik1jUnJiEBO3vLdCinWYciwoOrbmXpbm5K/XQ2
cCsvuJrkuA7sHB8CVWE6CjmX4of6leh7y94ttRtqdJWWjWBjJ+0Wr7KX+T00p+OL
aD2bPOzcDoI9RWwhsxILTHqDNazgMOs6zcEKMdy7zv0Uhf/yGdvf8x6vVvd8Eg7Z
jmxseD34A+qdHsq94tZKgY/mWyqDhqYeSjopeavpZ9ZAqGqZb6gBNudvRpoEOkLN
E3XWtrbpI7aD8+82ZiT6cJ1Ot7nKZtNqpNyrbtNZM0B5Q8+9p84XTnv83+lVJYXe
RhWF17cCqS8gAY1jNYzCbgc9RTr71HTccBtJhzZ5SeyN7ButniDtW4uLywUIhHnM
tgRXKj01g433XwsvSCXqyxJRnDxmIv20fhnJu/alfy5cjTbJONw251AlcqcieIDZ
svId17FET90448odzPohKJ8NKzg84dXQGt/1nQLqFaSGqfZQKlo1oI3A7OfewySf
Gv5fb3s7zEMmtiSdG6vxLz0MSA7eYNn8SdDEf+SJz8xrNkiflVj/DbDUxnuG9HwD
xsXOXPuDZd/VP7GRZ3eMBMd/+qp+bBlZxbNnwRSLWIlG6sEp8y7uLRV5ZaGGTfRC
bldYVpPjMIHiPAyGhPVKdX3isw8TPzZTtar4qjxGNOLKgA0cXmrPFG66ZdIGtnQG
1B/mmVhtjp7VGGWhD1UNdGOzLezsR0jQUXQa47xUKA5sssJQ+YIgWMSS2OkNVRha
IIH/W+LZ8SxsrPAHQlIsg/VWKevXk/RnoUXdrfzcxexv8NMmtOc/V4XGaxtCn1Ul
YHIoxvRjHCLd/v/DFxEbx1hRlyVpVjvPqQRwcw7LidRXP/JRcNmdMxh5dUVUYYwI
odR2fHfU4MGKb1ioDHthHrVzGDnN+MhmFsEq66pNEMqfNaokkB8s0+9WbQxzEhdc
bOsCzCTND7iwIMBkhOAkcU9+gSwivVU36wUaQdYdoJRYtzXlXrdIH3V5M/hKhAI7
5TNA/odNObeqGyhqkve32V+aXuzTBWu/y5n2B87Nf3GQ3Luwi4lxpe6J4dKMnziG
vAFrXU13sV6vnLs2bB9tsc2s0PK6vDGT0XKa6gMBLU9mTqEhVaTSklALlUAhKvFK
qnRkOsPik6J+JtZyFHyI0rV1NO6MXvgvYygbBpmnJY7QLYrybc2JguIA0FwU1ZFj
RJmlbdQkhpCcb0eL/bBR2BO4KfNHeZL+pTIRqyIckMxQjH9BmxiGrHueaoW4GR+G
O2xjUiLOl3U51Tm9wh0CZmuq4bCcXbr0STm3dFkwZIJ1QrgWI/s9nYXXDXHFIFGj
5/MNwMzCj8L/h3npqLcn+T1KpA30a93gZlwdH6l5LJwIFmI4PetWUiVrCQCqr4iT
CI41jzpTBRgOeaJoxZoFAp+9rzdRpUJvhnzZAOCqvC3RGkdzg69IoRxJYtznXo3P
U6D/DsPrbtkW13M/7wwh9bsiVvmPO70he1P2zrA1rgC+qrg2Ss642gOo25On70gd
zlP3LaQu9N3V+Mjt7wNGlr9iANhoZ714nFFE6kCSy5JsiMsljXS8/mNxg7NeslOJ
T8ldhQI3apyQnjvP7oZJyX4rtP7v29jUgays0m4gIB3mZ+PfKfWNVwfCxDTgr8j7
PEUVb5RcHRBAGIfRKwibkQm2gopx3XknVeYwoaRVXPkwYYEaBxyxfPjyH11ANaZF
EgMG06a+826xJGTOW3YtnHCMB4+o/c18kIZw0Jfme0Bw0ZpOym8XXMCEo8GvcYOY
NBvO7u1zETYetGfsAPf3KwKVLLBCYAieIFiEIDvBSdiBmesfT1GE6llsKPd4jFr/
iqs4Vg7/HIkPa7RK7wN1wXsSapho6HwTBp4APsTHE6px2cjVVwNwU5bLntXvD9mG
1ljuiliyi7Cx10lnILuf9JyaUYXMN8JbCkG2pVSGm5eZQK2jdQw0Um9YO1ycSpSS
LTnkLcT2xouNQsQs35OqWoksiiTtz3sRP3sTDyhcz1QQtMoT4oX0B2PmjhB3w+CL
jdyHnMxET76ZGImRm6d6xfmosNeiSfg74njEn8KaxqanyYKszr0lJHi+av+Gamki
EdkmWs9Pc0YJRBLk0BUOSmT0tCuxdXww1XoMAGl0chwnucT20zrkpDq8f5YwW0hU
W9bUIb9//DViunoUZ05V+/gx3LqUhtUauZE0olVifs2FyPSivgVxhwyBAz4aONZC
M18FNm3OeFIEtYUgADUjWaEE3j37VXmVvxhr13dvL7GoX1ZltKGv8mK3/7w8qnEm
XEHsVQkorGP33UTtju3+GVb9VGeAY9ZSisHbmY1VwiNMMS63+pGTiotXjtdOIzEb
7VIYGB4/2kMRZ+2FUdDZMGFspEWbs7kdHIPUi73pQsmXRUfG2ifxHKBBNjcZfWUp
QHSVlYknvs1GSlvsylDnazwQSAUoBFdoY/nfc95iJlfNOjBxeyxPD9e+FsK6QHSa
adTmy5gy41VWaYhoWsuEhcNJlE56eXuj4YGi/tq7WCdtsOAt8EbEcN0ACLES5VE0
R6OtWrrKpUvrC9VVw87P1dQMFrljj1rICEuL7Oxi6sUOcI92GTEbMXBDRqMtJxay
0RY/X2LM33pfhvLzRtYRB1p4wX8yk1cmPFVG37278Xhru/1L0LBPyMIb34EF1XfZ
mEVEikD5Ay4T494WSQt6UEpJyL5AlPGcgFmbudaRBMq0GX8O3ZffCwgmpyIkzpl8
uouNzFpRI2hnQ4ikQeKmz8ZA2URrAO6aGkqCp/YgqhOBW14CrjWjt5YaROVU5MPu
Y9kw6sPdl2iks8+tnwxbZE6oRgk+e4LCVSC7i+Sbjf9N3BWcou7G2YLw68y8WGDC
UKHJZ44d7IdjZKGSOKeWuZwSoE3EadznEtyNP1jacNcnJkm34WK/uwfHyaAX3eZl
1zOIs0lS1S8v6LFhy2bnJs/B+AZvHrqJMdNHbkXL1HHBZ7h2rjdbAjWo9mmB7oAg
l8xTAq1t5/txZmzgwEdXRq0ZE9h0taINh169lwNWQ1sYYgPfdCPylZ43dzMZq1L7
NPj+36JRsQZiG5WVaiH//T3Z55nW3soyyaKA8zg2ZnTZJ8UghEZHm00zHc7ReoCd
9Cf5GJsdcvEtESbrc8ug2rnNY+VIDy5SyZql6wR6wDKIs3e3Mn+sOk0tjne9Wk4F
xksfCT1PQ3dtGfL2/r7Vf8Xedf/zt7d/+7+EHS1RmslDwfkBFlF8oJwp0r64wlQR
yxjkHYiG8C9xBQNdPsm8DC3zGAFtF4sTf4LMOiRhRWuG9KgEsZlgA4xcnNRQKzxI
`protect END_PROTECTED
