`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qn3jO1jOjgFxl0OZ4N60DMbxpUyUx3v8pBVwEo418j2pJUmgocrLAjc7syY4x6hj
iLIkGZ+rOgAjCeYngrAeCSwcvvnvT2MLb64o6uX6IF+UCROQ9V+yMpSzTmJJoZ6e
hI8wFQ56EPPstnZl2wbJB+YsP4Kcmzy58GNNYF25x4zwml7ZkXbBiP4K6xJFKFOl
pEwCGv+xTJYgiOrZbIOUcnJeevNUCFHpxEPJp4jPVds5injm/gBZTAsEHfQz7TzH
0oOHS8b2pJkUaLLKdqlzlUqIGBTMfG7OgENvn3EOgcmUmUbRNMdr1XVjnm/1N80e
bPL6FgLs2VlIVxlabM2yTB15P0G5oTcorZzPHL1f/8VeSzfj6ZzxHcLa7TVGbQVE
kGbVvP/yB9k/Eso6eSdYMYxkoJuJgQxjtjHzzsK3p0qft2LtisxlFnemK8jFAfFd
Xa06aJxm+2Rx5xKGLSKeTRPcQ/nr56lxrZ2mQMl//ip4xVfzZXOW17pU4XE4X9He
6CtTZtv8QUbx90oUtAVIlfASpOtlyjRBI0KQzPXMrjqHfZHbUzK+cH9elnwV8CuC
J7QaPJy8VS9eQrmOv0kE3OW6hu5dds9oSFYNE0/YFZnTggWa3ALDc5ef3AtYA602
bj+/BV8rmE7sjCbl/HqJkHILOceLT+U4JVTdCRmSX+THLGSwd6zAHbvFKbd8qOEU
W4cnPJk+OsuaDI8I+kzmB2l2oaiFtoZRGQccM+Q4E1ImVZWqOJ01plmFVRusZDvF
2YAOSPQowKk+BfzTFQIy+0qwM04rYVvjEnQSO4Wh0MscTxFcCoECiVgJO+ehCp+Q
FvTG/9KCwJPXl+tIfqfRNUmnqpj3WEWov1ALHvI/qBrCm0qnwVrW4V+sAn67AHXN
wvGB0znTbelbul8/WAnbKHJa/kLFeuissAVtX+l+L/VyJqcHF25/SfvAJM/QYufS
Dj886MLv+Y775Rc3J26diN7c0mStsKFX75PJFISnHA14Cj59BR+9zkkYdQui1lze
Hj7ciD5Nm/fF0dbktqwYwcu7iJIo5w+TKQSWB2+1uKLImo3zH356DN83NVG8X9Ou
7Y1n0r2S1gQYhdyueIZ0GdcpuN9bGtLMjRokbjSfZOT8MU/xNb356Zk2mVh0Fi6Q
Yn5mNqzgLacJf2cAcw92Y/rmbeWLCNsgE6SQaLLXe5FO2DFhGRf38m93QDbo+UO+
i0FNJXbZau4mxnMAWgHC7K8BWTvfTvGX35URQnZZbxTHemS43GhXGHAsm7mZLENG
dhDhd0jGimiSWPM+LHnkXM1wdmHmsqjnDS094/aOtUTnJAuVgkI+Y5Utp68FpVU4
QbgeNYQzC3/7gCLNUQqg1GMUNMb6ylYQAKwf+eIYQm8BENGvUJOfBvWDBD4nJE89
a2n2sCCidLOSgEQQFjR4StS5CXd2qU9g0w3wOJWZlLdKiHf8dwXkpRpTU3zlwaWt
S0rpxw9Q0JhKygx7j7ZpiE9Y4ALhDKc5PZo+eX045sb58TmvjALQr8zxu49+fPen
TYoozFG4jnsrNQ5LcdhN4tyPuxeKhG7Fnu2b21CXjuRhNUl7pBWkiZEMHse+7SY/
Yw7nx8GNLZFGwpftPCxJM8c+I95TEhrgpcrtwAr1QvAzpC1C4GrxMm1dIRn95o3b
CqIiT8ihouoNwl0bS78zgc/OLUgNt8ttc5I0ruqEwmO9L2jy1pZJ4+2vLKRM+NUL
5Ph0lcYJ63uqHr5Rti/1/4Z4jOavyOVdq3PTiMQSNi2KmjzA0u1UJzdGMIk7YNFz
X/CaSkga1GAxYrdMXX9s2DTRzK/KgcJE8gLRuaYW0CRSxkMzgqrilDGCoqUMcYSj
Eyv2Dj2u/apLnUVsj6TrRC5rF32Y52yptEZ2pq8bzHDjZcTGN62Xjr1wAflOiC/G
oM7E1aIfz+1xsoQUu6ADksN70Qc3LtG62WGlZruJcJWsou+YBdnEjGSVSPeO4gSs
uWIabozY8I2hMb6B/nTLH3tCuAoy9npNl6e73+w7Yu5/vLJkQsTyIBNg2p+ZW9N5
hthX4njvFrPTjAoqo4IgRkuFEFUXIf0P5yS71m/Qf3nEiCG9Ylbe893JmXa+2nyR
UlD5l9N4xeut6R8OH/z60e4pAwAtut6qNz0yXKQiN1Du6rPAsh0G+Z3TXlC9aEAh
720KdeHArT4pWHO3F5oxTt96GX8dCkleRpMg4KkLJh7nA11BM8QXNgslF6pZYCOJ
dOMQ9JkkN41snjwJhw+7RF3sQ975TMoiJfTu4gDbBwg1UnORnByN7N3j9ht6ddyi
MRAV4dmqfUpNA3EiIpN70AOk6Xk7bskC+KI1zg00Qpm2FgK2hhODxmvg6614VKn+
lvQQkry3oj1LRhFUmXmUS+LAndXbFQ+KuIgp0luo9y0m0uPv69pCcLl0fYLWiqIV
L8i2z2YVaCjolknb78JaGbkD30aegR51bnsV7S5XY/0NPNqF//zlhrU93AkXEfzu
BUWexHMuP5mZL1Djy2XFGQyZ3ua3O++FqpZfk1FJfV6wh3UiF4cDEUDffP97bvWT
C2XnYuoqB8vktbnvkYUdsmy4F+kHErowZcdIfG+Kz9ymXRLLA/poNrpTnVjXmMYA
QUGfozwa22zNmKJ0lDwTjpdM7QsAjNtxvfSdXxJ0Msi7EttunW3l6FbTRKJGJTPg
srNebRXCxxlyXBtQK5Ampcw3Oeov2eOjt78pdleWl3unCt1YHT772WxQljO4fHWO
RgX/50PymJPdeAnBJ/SJY6E5bjEW6l2FxznnFMuK1o81/MShBcRhjLZfgJ60kNQ8
VP8wCtUsUOC/SpK34QOjbx3QXrQHvqSqqfupNuxRJO8azFu/wsERQVJDBzgh+ppP
jSLFBtQvt3NaYEvR/UO8Lvzigk0zow6nrhILyY/we4xhbZwcBOpvnCAnwhkYQhQZ
2S8bS3Z5eyXHwYxKSz6/YgNFnvGuZooKIAyHqbnsP+1BuiesA39IwYo4IZQIKoM6
a+hUks3rbTa+iGFIMjxk4oPvAadsH+iyZRFdOUhJUbQSZjwlry/upAHyM4rwDo6W
9lLH57sqCybXlQ1qZk65gbQRYDRTUI39riKo94I3z9bGsoTTWkwcJr4bV297Pnbp
jTR3tcfuPlGQ9tAY+016sn79AIc/OUHHO9FkevlJS3R5bGq1uvS4e/aWMgHxyYFG
SECYBgt5na5hAwYOHdX8YYflv/uURIvlaoO0SJ4BOQt+Gx0Ee05L4LM3hee+mZj5
Kw5kItPa+Tpe9vnfqwgdjHs3pdyN5P3XWDE0djnYKPMBpLn1b/dk8cPt87nTSgqY
vusSQawtQ53aYz3Om0bw/2OFPapP2bMWTdLwT1RxHq7DyTInyOlyRFOjCr50rwF2
tXCw3N8nyLgxzGxWkl5QV5AjlZkHhgD2XC4O7JRMobCZOkCUL2efIU4nJVIpeaup
z43V0Oj6MS9SCSr0u4CeH1euB6mssno5tlMngpM1Hr34Jl2VI5pHqwVRXWmqDRDm
PdXB1LcB9dkfd8KgW5yQ2JCC7rvJOsM2qnnw7g8MLT2iVz0zetp1uQU16ceLskRz
lgSUmuSNe+Ru7DFSmej8CtYhe5UXc0fdIM6430csMa8JL3dH1NayyBT12787x+yG
t5gvWtteiST1zUPpHf5P9YKNITtKAJYFvXpQKCQ9XrRaHXfNNybRD9RGfHX2gfOm
MG6ktCOa4G4v2NxoXSJHwjYc9gvhs+1RXBcibXYnTNf+tAzNnx1YIBEOIz9kanUA
OEptxcCyl//KRVgAZJMT7lbyLmQfLUlF5uWxMiUGLtnlOLLpjLU+RDUOiAdqmVrF
8kNkIVppH1wipgs8Uvw+vOivv1dKqU41uTyb8GAHiKOEAogUITwZfynOXR1Lhiwd
iTeWuLlNwRmtCgEV+5UlpSKJJNmO1OtvREINP+KB7WchOfGQKIuD6pQqtpbZMrNB
isRfTK4Kr03WzHmYHZyozQ9MFX158/dVM+g4njDdY25ECxkL7+f+5aJnioZ8i4yy
iZ/10OwjSRU1RV/pk3SgQoJx9kZ2Bjf/wGE86xBaivXJ2yhki1VHH8B34wW2GhAr
pvLDH4oatyaIFFaArw29mIO4YUUPhbDHmLavPHhiWVdhf5THMH3stLTVsZOJcMIO
opWKv3hqBjQ3TTxBpKyrrGf1FYQJ17v1gC+ZdiTeQvlKxILvPEH7F2vOeDWV3Eva
5zdh9fGPcZuiVSwa1IoHbAQ019uMFUTbSNbs2K4L4/XpW9RhhzWsePlbU0uW+wk9
CugMZKiwK5dsX/lQ8QAc8cgTKlSSY3e//x20AxL/1if9oVJNQkzlzjL///VlNDGs
wfs7g+3pW+dnJF8s7K5m6McPONFedqEnL4Pzk3u+vjuvUiNF2qNpYxwj/aVeWRiL
y6mscYS14Lx+pl8+506JtA4gyqBCicQ042pFphRznmSU2E5UvUnePiYkjEdn8tl4
I9SzzyfDmGs5x+AJhib9zyIwgEEvTPgN4rKmqzzM8KAg5ED3rFemU8noyf8ogGz5
j18sVt0bdr6ApAu7vlrxYd3KMkykRWaErv/v4oRL5aSQtvIdh61kRYYZornGXfIz
Vbqt+RXyEzh4G3LW7yCTMhP9YNjzCV9ZVU+l5LETNWgscrHAKwkhWakBkXt/3/rf
f1QvA7A4bGQWB4ObvLHN2ZOiEl4bcaMF8oaYEY2ERW4aMT0Qk2AAXAYSomlsj14R
cT35idhddBFVUbzagFkGkZfBS8s815YLwGvDJILYot7BcaHv5q/DlHAWsFDAeg8/
YLlVTq+Rf77S30OJi8PM2RP5MV1VgpR1yBweeOMcI6qP+i8jXjyflr+hh7QxrtPx
pYf600EcoaF8xKURmLwhAUKtFFwlmFsnSNnBv3Cm5cLrSWVhgZIq2l70R+zgoYul
NBu9rIoJDR28xtz/bMG17zNULiK81x3+t0ng/x+Ofo9RdOBuVmZ1EtrzfJi7Zlfb
D+WpatZNKHJ7d/5KvGpFVUrRQFDSHtYFcVXjiKBC8eJcqgxi1rpdRh5z0FdYJZf1
an9wLy0gU9uSKWuVQ/ruVaVznC8Tj5589cHnOJbAjzZMWWolJVKh4uzVKoeB1YaA
ykwtlxonMjnE7bG8NIOcGHHh/Wk/d1tCgTxe7uKIAgjNJnBPtNhPUDAa/eniFAAJ
7YgrdNHlMKl/9QOQpdmTwVwXYuIOE5BeTyOB7tZxQwJDO6JDNlCsjxwIbIPiCKGU
20ziBxF2Nq8JtJqWK7SAnDIGXGZF2jv+kAZCzcRs9x9T/qe5pZR5/+27/TYZYxXm
YEQ4qTKhxP5ROdZl63WJh8lp7np/N+B/HogTyBTb44CSRAsaxtWnGl2g3iVSLNTG
+Rv7Q9/mucGhw/rMjlE048iESaSOmQ64LiMOHlt2MJKQlp7Axz6L9uN7DdJdpS5+
n5CeEBptqU1DtEWHA+XKZaO6CRJneCzazxp7V5y1P1fG5wjB4BEAhWbkk6+SWJiw
e8OsSJggW7nPETUyUEvPPrg8+l+GFHPKggS15fjsMzXwjRA2MVvOQbHT9PF8ZSbP
oVqv8V0+a198yYiU1TUZiakE+AK1hO8s0CoftVS4JxOsVW+O+GCyGDVYAoKqb8G/
d1oMj/bMxVObow3keKrss16rSPjyK18ahP4ZmoOpAmF1OuhqnsKSWDN3wxTCzYOh
NNcBqvXCBbebhnNRijk66uy79o78zGvok/0y4NAk8REA4geQ38CWawZ6wRqMvnKo
AFIHCPhPvvMYu4xeSXlI3ZmQscnojM2LYoweWcy6eBjyP6jyCPQYLomVwSbIwj27
EB2VXKtpF+6Azi5pXfY5tz04i7t0wzZA1bv8CC8Zy80ik57ydIaSIOO7FegLFDLj
Rfa47EblbX9O6I0ZLIfW1bYu8TSV41jn/zidi1VGhyK9F1SFKuwgNk6SEULn+W/f
uG2muXr7mXbzI9CRv6l5DEixOBgrDjtg+Q/DNJb84bfwPsYuAvtP12omPDRMFI+R
3w4eyRdi2oNnAUmskFr47h7n+lToa8ZGePLilKU1SQjkK1L81wYml6mJwk14wny6
k9wLGR8KF76vNnbK8qUEw7qQyjDwfiSj8UfACG0yarc9F3i0bSC+A3Zi6SDPz9FL
K1gvwko7EfcJSlb4IKmdg+EJVNoAZXA8uj8xrNVJojoZf4XAicwOwGO5H9WLgbXb
9J7mb/JPjZSh3xkEZ1CeT0saWIpYEtMgpjSYfrxHAvLZsq+X51MyAQJfsFUVI2zE
D7TjevV0GPWDOcn296W9eaKhNEOHaSt1IOrfLNZtPFMuem5lhOe03G/EOBk1ZLCI
sl7ODff+MsXVrJV1bEk1VcjwNQ+H+Q4Mg6IKVRushMpP/K/p8RRhbFP2py3bYfwg
xDtwotF6fev/jXAky2RWYjYcjcanRQAF+oEAmtxLLp9ypZf22nt/VgSlhaU3UIfz
y0HZ964U6QowI+6dMHJhIVXKFi7NJdIqoVVag4avwx86UE4O+v2QeuENcIb4JrTf
J3k7ggxq7w6P2Spwc0QdeWUF+wifzNpMCiqEyMvh+CRmHHFUIuUNKC01k7FIjDaE
eXKV32G0gBB2PwgCpK51AiZKQUUyYhK+I/upENj/lIM1fwRfm4Ecg6qhFl95a6pK
8XxBb3UcbUx9+uTFFvV9UmlQBxmr4sZ3bqCJmcrEtpysiQwD64C7KMlsroXWnLcG
VsjPKEjVS0mw7JFi7vXrrbruy48oYBrhir5eQ/BzzmQquQGI5W3IvHxUg4dFaJfp
4JuTjwkLvSvPejjsg+aisdTcnrRPM6ZiGPmzrfhjmAcIFrkf+DRkn96xpNyTowzQ
OPVA0DeyDggW3xR8jRwDyoSxw/QYV1xxptmeB1QukQKU7XXy6e7U754HNOvk6kLB
+/1MiW2UQoNNuKPNSwZCHmUxzPgATyELyKv+3dPHobCQ534IIv/IlGcRFt3v4bSd
KwAmr+HW/vTgJuRC9TyUB9ZnCG+5NK8zCq3IkQCCUc245QSTt6Nq3yv/InOCxmf2
eUaQ50oL04QimIK3EqDg0usCFU2dul9i3Mh8eeaBe4qa4aRJSkJVWlFk5O+nAfZf
T3QKU8OZiM1irPHnFcEL1ahHzMr9T+JwDTVqKgqLlu57G+o87ncBOssp06Q43AFK
w9Te1zU0hVDv6vuqCpRrbSDK90oXekPiE2j5gEW5835+cWNFxLdWMADSZAYmgnZa
aSvyndaaK15Q+telT76mOudSwiuXEEJJImPU9xpE2lS2KRMo8R7sS6ksjnOMU5Dy
KZ4nxsgGkCiELxbZuypl2ecNDRnlCpiUtQHQLPc0HrbFzUW3FxFjmz6QR0j2XOZz
q6sSEqL0Vkcb2Nd9wsvc4s/mzobfZiLUnt8w/3lIXr9K36VUL/2LbdRAQL5QqsNz
YfLeteMI429N8C7tuiPlnuNzx9orLoTH0L1x40aYf/JfLEJphsRid39kDcK2M7KO
5ZW3E1RbWuTSXVmoUwvOPXCiWoaTbCm/YoNLewm0CcLuZCqurRcqLo/WQvSmqJT3
dLgV0ZwGoUn7MB78mhAQUqnJEAXOdf5Si7JRxqQfnJkv7iuHiq/bKFvxQ9QBUTr4
C+qHpEJs5N54BmeirQ/yo8o/EwoH0TFqNqKaSpW7lZ/lq3vqX8UFHvBFIOIPpBHW
fgytVy/dnIk4w7HGeK3dE3chcIoPuSHGIRm/VHnZQk3dXxSfhhMGBvJTkc0yFBFB
cXCS9WkJ1KCS/wVEsGmcJjkVzJUPqjq+9mwgbx9MjL6aWnVP7n6NdfFCZfPFXldk
TKoNNBN7MQXbkzrAKdunUwyw7EAQedXA0yU9bLzUAaUpG0v/feSE8J23NSOZHa82
eXfdJlkAtwrseG6lsMNSBgzfMofbcl3ZK0UmPJVh52yJ39+k1pZYb+otBPc6AygM
L57i/KXLliiku5sQ/p0zaIeYjaVh+I4p8bjFo9OWz2UvpPSAZMfkfnSGTfc36P8+
pACZ4YxPU9sANGw7Tb4jUsHMVDr2htx4gFU1J5Js+Hwn2W4vBYPa5pDUUCeqQH37
SHIQ1pKA0HdI9tnQ1SFb9wU3dd7MTGyuy61Z5bRHEvSzBD7erPUwnjgP9vharMlV
jF/8jrXYTuXKUWZkX+z/F8YCnuClltFK8YezTmV40s8FYHy1uMgfF2zONHZ0NPyc
uP11c4RcFDbiUobsuCkYQ1pVOtctsUqaqoPQz44f+lLIYILMEU4A3HT2yPXVQh25
7YjRKglBWp0cKOGrTCCRcJWwJ5AlnIih1Nlpi6OeuSQA/PWSY+eTKg1BqJJU55C1
12kRKPfVITRq1tlakJb+Rxw4uL+8aDSWdlpMibTEJazaE9ocghi8yJ4NOVlDfF+y
g76PbWCbAtmnacgme4Xlco3yX0PO9O/Jub3a6sreaZUrmV+tE4j7FWAWgIJga5zG
WLYkq2+jEA2Te5/5nM+9WXvMvMQDR5f/wdP7sg3m5S9dFKo9r/wfGje53xAyN5Xb
uYOR9DlBH4y/IF6JzRaOVkRBLkBTS71PA93z5hVKgFrZbWy/sYiy5XiQ/vN1JeBl
vwKOmrc4TjXqjkej2RFvfsP8w2S38/h+FjtYIre1lbm0/w6H4xi0KhUMNs06Uflm
bSyb7ZBifOFneDkNkvgpwupVBW3SmsBi/jwASZBHdDh7txZqtGCkoK7gVSf1Q573
TmjAuWLOQDqlQZpf46epNpH0VIb9E2TCCTmcYKJQxGgUUf4wBNRLK203+dKnovjN
3VKtKu7RwBoRdmLFmANA3Jutgo905TyqhgaiBw0FjhKUeYEhtPxk+dmxUuuOexmN
fex5Nqqqn7TGj9NeFYgE/YdrJuwqhSJYXy8T4Wk19h9FsP8hEOw5Uea18/IBJZWB
fIg+nZHj6oAbTJVmwnyob0w9VsgN4ZFWhkazMMD1MflkLOfISbEyMQv8nyT5Sl08
X7DWbrociRyBgdtY/HSvTBIRmxX1zyY4J2a4KNNLvLqx3phsy67YTc0U0UjlVLlf
wbnOjxZIkb51hOsDUPZ+ugiDmetvwDQSLvnSJZD5538mGeH++DpqR91BSEUF4l+E
YvkKGdX7A2YAAJFoCsCJezbOlTvuryF1qWm1ZwDl7VIbCC7XBi5LtWcrDNTT2VT6
Cn60Ny/V4LrMZt8LYelMuDdIN48oLXvuMANyY5J4KV3zJJ/9taPwVddCLhXsejfZ
FSPB+YfDQvj/nMQWDmPj8VZbAcbCbbTHjO6e3x3343ihkJerxZgABJlIu7aI4Mlk
FDqla1Gzllein4meMiu7wCx8G5Tv4NfYUpq8hlH/7yIcHGyMm8Veo8M4OHNnrn0t
m+b9Mbb3OT3D4lcA9JQL7LHZe3DoEBEu6RfZ8PRHe3VfkakXN9J42dNHwZ0XFH+n
Z8ZkQCrGHI78DxzNc2sblEUkgx9o0t98kNsH1PSmdqJK5+krZ/1//bWHkJo572HQ
6K0q0IOUOvAPGsF5OEHxtGL6fJY2C88yJcm247Dce64hjcgtEctnLsD2FdBuoN+6
jxp1Sb6CH/6i7vMY8VG8Z2u9Nr4oqRcxnZ0xEG5uQwO4h16C+Y/mZSP82kXUID6J
snAVruFDxiqonEGaculeuJjtR7FbRFRQ9cigRji1genParT+UF5ant2qvp8jz9Tf
roAe+dh3wAID+3keDmgHiL4Yik9IJ+gXVz84pIsMO75I0/JUdl86P6uaDuLm5lkU
Nl6uc/+SWMxKQkj8J+xeOw6kFcGk1j1uszSU+SXjE6xmdKDmUxqVEufc1M/NmykV
qC39rHbmWdbogcUOecbS7JVgP/oeBuCYt2eNzLBVlxCYZlhkNJnSm3/DKlWVEong
HmvNh9wuURC1ITC1wPmcAyhPW5qOjTt/muXBD9mqlw0BlOKMnb78sarX3ozKeC8s
DFfsdGwh+ErYN9o0Sf/zTfMScNzboyu7LzOoTptaPPjfsM508DpM4dJitOrx0hXp
h2ESf8tcHfZeMeb+u/RP0lii3I57jJHAreK4VVlZTTakERFEa7jJTwIner+T6ohZ
4sQJkJQQo2Vfyb4BXmvbSlaAnu+zT+zJYI5qcAKn2MCxi16VXUCbLw/8l9GAE/pA
AiptKx90Xq0Du8j64s6sHnyvptkqBowY0w0syqAm4UwsQOK7ZhnZjppGgHsTTHRg
IB7cEPMGDmfoINhb/lkQToxWwmapZ/jWqfyXqoZn/+SHyfpRdFqvEq/RUfjilX1D
emK+Dy9hVHNzM8JDyIMfeyuctAledUcm4ttw0RwDCV9zmb6T9ql4uh7CE+zwfs0M
05GeoO0Bxe1IN78MnD2rAN3oP9W41oE7Z1C6NP+/PUiRGjHtcBfhBH0K5354io/O
o8t5rfzJx2prLRxFweIuJiLX3lFxnfQicTykt44By/lZXSPn7ZOVI3sHy6v7WvPk
mkdJt1FuTtDWuA2aSRt0F4j3Ysml58nic1qZsXz1zJeL6FBre1/gjXRVIoU00Dn6
Dwb8w57Xm/Jfo3+OhwJPtauNieQxf53pDdvQRGoPwbUrf6wgu0IcSDBs6XHSjLoZ
FTGJgMRpYR2jfF6HFxNojGKCj5lSH0zX4Qg7mW04tdEM+uktafG5aCzGjTqC2pB9
YIXkC0SOK1QE9+MMXRKjxLlX9ngSb90A1BbirheIeLcDJZ07R0NQcLZPv+w+i7OK
PnXWwSPunnA6fyHfvmmr5/m4wi/+dUIGPUwy8X8Ds/OlgUHvwnB7wBwsRgY3uQFY
gBaaNKe5fyVN6yydqbAj2snLOJoHEpQEkYXe3TkQ3mf/FVDxtMYlQPmkNXzZB5Xp
o3/ZES5HdkQD+XSFuhr3Gf+Jbhv7tKczg08V4xn88W2LOcQ0q77IwmymaVuiu1Uw
PHNMS2hHm1pndHswRUeiuMIiceq2R9Rhr820S0yLvL1RFWhKja/Hq2ZrXroRsIbE
m3RJdJgH8XXLXEsOPRrPNCdGR56xiEIh0uC55MrdvC3ponuPIXG+W8CcoEa7qNy8
j6zECba8KjDXZDa96tHgjUp0mkFSmpImDLEEqAyDKJmQCZ/FvMckgHpTjTxw7lzF
VhVMRoMaZw1XuFNZGI+9XzFi/7hjTwzRAFHYZyMe5Twd+NquxOZyFJAP7KzVuwsA
OQS9trVo13Ov57qWuszvmRLHzkApMpXNalGVhQh8ZT32J9ywxG71wG9qjYppt6IN
49p+tu2a0IyGwoPRKGPWvNAXh9J3u4BzVn1gYmmJwE6UwLfRb3uX9f0t/R0Bh96p
7RwOujXB5XbfMGBIw+nlq0KZYC/LTX83Ed89dK2YVGh7BHN7NZuVYr298YnABcDl
UoYJP8PV0tXi5o+jjuhGMiJzDfiqDjHGVInCc+qHSF9k6ExofPVco+jAh6mM+rjD
XJEaCgHWoDaHK6PgdiODC2jk2IPtje2k+9aIDRbTTV2eLLWoJOh/NW67hMzSM4gc
JkQpiAAVfZXtgkXOKhq8czHY2chE2ZYlmRboKcwBbSGIjgoQ3Cbau+OqGHyiSK1V
3PCkbcxS+x2cjri8RhM6gRXdXAsjv316gyDYbnYfMduBTgBr+Gw4XB6eu2/l069t
aiAxx2eWrhEb+6TWMPsM7nU+NkW+m6pHGtBKmKOwD0wPjn6dFKTYOAuxeg/wNOy4
fMXvzpR5DU9Uk3Pe2qQkrnINpODlJWqbNSrxT3+jkq752BIgMnLmqzOFvvf3bmI1
htyMwzj51Q7Dpm6gsTwUxxXeqxKk3/zgxsusnaX/npkUkSMRNW2FJbTBZ+xit9dJ
qtqcFPrb8tjzSLZsGYHbBygrDneXZPh1Cpm4boCxJ6OCeqT0AioatdZB+HArU3c2
SLxFrOljc02OrFjXQMHXwKXLV8F5/dy9tZqOFbjj6VYMy7ryxzrf8KurAzoOvnYm
buWVuM9OtgLvZUegRcqMrHx0tXP2TEDfjvteuneQVX9l2bxGdBU+V1NG1XC9Jj6E
6FoYN91x9/paMrN2JwW5w7boXSmcrG8EfYt8hHI6bFR8iOfdP/aq9P8V80xvGJn/
CnhcAa8on//Ak0UxZfBA7i5OVTTH4M3HHHBaXPDpuEDPRj1VTTsVhbFGHmH/PxrX
SlIYv3sKJ2YDnA5yn7hjQD/p71YrJv+WgCt/PuBdnpXPDQVp/gM7eTdFfp6ynFEQ
1YqVzHoR3z5zix7MbXBuSwt689TkkHbUaA5/6flvMHeO1jN8AUEvBOqrnnJcHccK
jacpq4Zn8au1rCzsykKPAZ5qMdYPyppvJrH1RnJnS9YDjuaD3OxmrOv6eJcJ/LYz
ZsCAr2FRCdZrbwol8709HVfGKE/x3Ra9l7SpYqrExW3BDQgKQeBXzw6XpT9mapQ6
cYXfjtIK8EQD4wUEN5LXMWaBdRcP/OCNxqm1RTL+W3yal3yHljh+vpGgzVNLdd43
LTVH+aFxojWiNTgQrQ+XyegPSRP/3ToJYwuqOa5Rzdo+LSUGTH9np+jmcKlDJDo5
TKPfh6em9C4eYtgsuB7k546TNT02PHW/tQ2+NYFhRQg=
`protect END_PROTECTED
