`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0zXEYhH2B2HsY7Zmc6gnEgDBYSFxcfcG5+PDtNjFWn3+gfDaF4rW7v8zW6cqkD4p
KFYFlbKOyaRtZSXVTmYFFScuKks2X4oE1OzFfCt221e+wS6qIjTud+yDGPWHrCCT
qCXa+8WDA5gJZRjQiK4mBlw9JI1PtovXrZZJx/d9V2e8A2FE+tzTWk778Mlg3ifL
EyNFu0ucPhJUBaLolo3BiFnWH6PN0E4XesylfigxNHOeUujifAMAju/kvgEXdp1K
TCmttZwEw941Mm+oN7wxqAQNUD64kbmR641G1EqowuXodml7OpU5812utZNwcOQ3
Itej5wRcWJRgZD3EOgbURIEF0LmtY83wzPaCdhie5yMWKJow5+eUBMmGY6EvV2Bi
xBnAI6RDaKqzLZuyiaYRIoXxWics8lnKTRn6CkSkrrL3E/8WegrS7qeFHZewlfv6
9dmY+0byttcWWwyJ4mwPZFDzq1xRRGa6Y4GZZ8yEyMW3D/7LrsDgVEY4FNfKudn6
vW8Jcp+OG9xGh6ReYkDHMYQTX1v3E2pfDZJ8DOeRVE17w9rpfeBB5uSxc1khRTz1
aAbOxm3P/L6gy6M/+0u/kHhBmPDAl0NAbkCP9iACocXKbaYs/xHjW472iONlFi9D
Cg5dkDGa4YPd/vWr78LVoKPgMzEq2IyC1ZAnCVPzj/S6+4fe+JZnizuCr7U6nh6N
atpRrP+dAr5BTY1MHC35xR3UhI+E/C1aQKZsXxXvlce4u97AUjXUD9RKFClFq1Rr
BIaaNJp11E121vAQF1UgIW1eyAvq8LOqjufoDOvClfJqv3oit8QeLcAVy/7M5br5
`protect END_PROTECTED
