`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ALeGnZnHD4uBKq+SN99HvYAxDQ6uuS7vCldv6X0YNhcI9eWpgB1zi0XB+gbwk0Y3
TuFByEFv0L6vec5XazzIw71ZNhQ2rPg1xxCMDhQIqd6ZSSKSCsCi7KYFoWe1udVE
sjJy81WFpX9ur9aCYb/Mf/h4Jj68LL9GqdFkWZ4Uwf4qzY1xIsylNdjd6hHjeZl4
z0/KOvn8BHwh1RNvXY1zsz3SL4005EVGIZ9vbwc2zA0VTzlwF4WTFiNVdJ0+G8jk
CzGl+EKHRXMzDB/4X3eHSn7B8898Wm13RVc+nsjdrcBfTiZIlCUIWLWbaOJaUisG
hWgRTFRbTLJra03eo2SHIA7yNrNrTATJTdfcq1Sw8cb0nsU+E4vU//A8o6uIy16w
H7IQe+QZwvu0cWQ1Jd+Tvh1meAongWA1RdEejaFH1cVTKzGT4ubT9qfH7212fOIK
AakDq3lHRqM9arnv2ApV4yanvcnrda4USDAito5AJrVcUZe4QXOzOXXi2ErGLdiS
7fDc0hNztP42VN3LRprGZYPgSQSlxmmCeS02lax32OZb5haeeM1k6EEbhkLAzzR5
jeVJLodsigPuIOd5y3U0clXdNpnBD7Av4bwCbpA7n32fFjKxrmK9LbaaxHqI6Gxc
NR9GLqtKL5nppIgMACm8lP1dpE9r38WWLUf7oWB1ZBPtTtjYG8xVcMyZnetbsAV9
ZALfet7WsTK4v1SUDf9QrO8KqXBKm/neu6WPVz+LLi8OMVzkpmPTN1qCBjpJnB/M
5+/KpzsYylE9HHrxPrRKKDPlbkXmpSu6ljvaKcSAvGJJVtZeIv3SPcMUQoPQrSFM
SwqQjPBX52MXve/M+VWZkIsJYpX72ejHp0PRDd5S9ylv3GwkExuGzVhk5dF+rWUB
indSGWFE8yGYp1MB+duTdXfByTkgxhYu5tJp4fU5XmG9TKwmQkULO3OcolxQ+0Gr
vqgMA+wd3vlxFCJfG7SZr8cn0w7ySNYVndDmXcIJHDPVEt9W83bDYHdH5u97Xi6P
4T58gazFB93QJkMdmkTeDlAxemtR2hPR5KABiSuzNeuDhC2mLYQDKa+FB9FjAsBH
35r4WdjdfLYlaVpMFQjx8g==
`protect END_PROTECTED
