`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
06PS8zEyFsH1a6NLSshjXXAlhwdQ1sce27PFEH7IihgBbbTW7ofkn4tHNjrOuPzS
xPzxBt1D7knfKP0h7DRIjmcQHzXZS3vO8K6Yv0p8dcsMskhijoksZpZhkfOfo9g5
vFEveLOsds0uRzx0tgen32XZPvGEKazeacv8zKSVO3jBbuXMvWrjgzEiDad3BCfQ
7P5ufUBIwtpW48bNo4CJiaTUTUNZhMPXYM/9fclfAfx8fk1ywqceL7B6jQYpO7an
2X7dsCQxPh9qIOPFFOdY0GLAS/rVw6vdUcPAO/EFpLQbDMZGko1ZuPLzv+RpM4UR
ug+BTrv538nH2U+58uE0DGZZy8C9aeTaKiMT+ScThtelUxnD4Y8dBHwRFSG8k9Oy
qsBHOhiUM3Gv/I9AadUcVrWscVr0KgL2zFu1Q+zLX22wAD2g7IDF4DvkDr8VioS+
a9WnpfJPoFQz++inRzJ9ncyhypNOvQeiuaIwgiooV3gXV9e7jTKuFkGpjVsilbK/
FURVOwBi/Gy1qD19IAIMxrZipLeZm9xnIl21Dd9VTOEVV/y11JrLzWTiitqgbFNH
jlkjw2pd2ThRw9MxtNs6vLYCyLgDgJJw84xAF8DAcJAmp5VdMdvGp5TVSF6MVzjb
zy19raLCR7zpgya1h6XFScUJhLnPtVub5zaX7r2NVN91n+ljxtFzB34DIG2Bj4FZ
7Q88YPoZ5Zdd+ZnUGwrunwiEeFe6FPLyOtpAbcJbF3fMsbpP1RjvPzwYlH3QyJ+/
BjzQOc4WB5ZxmnA/DjAPMMJm2C/3dE0nJPbOlNMeoZveoB/v1bqqZeIf+xnBEBT+
spWEm8zX2BfdqEU3K+LtdVQKtGNBjz/AYAqJQ4SY2Zl8Bt7m4fbt+XTjikEAXgrk
uma8z8N/a9+BqyQKGXFYwvkW0Ts+g0X2ecN5qBI60rtJBKgyOndsX/HBTEBeQnlh
PR6PnItiQ7YDGbcT8KhJA9af8jvjSyK6vE992HIXDm1QOGKvWLuTYDaCBZE/ZpDw
GB8WnesZYFp/8oqyis++GMNNn/NvdsrZQyj8SsedGILu2xYf55sBbXXFMWzGrOZ3
FF/reO6iuAMQK+qRZ0z7QrjUYbkkD6l+jo16BB6FN26JjmP8QuxXQTNhkIEauYv8
dOj6Rspq49SGpxiCZv3ZI0AcIuTpu55E5Az0odXz/TcmY1DGfTQCJ1MxPDz5qWFG
403juMhaSRkmkofCVbORIWYzWQxPai4ACvmwlDAzl78d8ovyW/jfcdsrYG7StI0b
kgncsn+Ph4zpxqi5DeNwm8+A/njiCcEJvFX5Bp7hZznpvDnp1TBVqptiKVeUKrAp
c9I1tGCesTSqDCJN6wSR8qeOFGOeTNe79jwlseIP1AybkNd4rN7dBWGeIZ/6mwPT
PEvBknOMhJoP1FuSBHhG3rZvTzLDFufut5zXDFaQMoCCl93IQzRDAuG22Z00qIHe
6aUEV1tjBTD/6ehmquPlENXtdbDH1HKIHrRPIcxSu5q5i7BBQoo2KMjPQO73D0uz
Yn5V6jzN651alloPY3e4pugnluDsGN7Q7x0hl/gN35KBtBQVPi4WvWxTHhM1YKjq
HZr+DJ2xR0AAC3CgacpoADevQLw9c+c/IH2nPVM5Ka21eULb/5hRMzKn57xyQ4ZD
R06Cktq1xMQxx8BuhK6shYcN5GWTR3N5okuJbWHKh8pjq7AYw2hHe50PV+BBRHSx
QljtWZIzVozyWFygj2UdTmxreG79oIGITbaXMuu3lCF9bg2rQUw9wZrs/xDdXNza
NK6UyDI5cwmguT0nAPPILHjSMZomtDVU7DhpIZNp53S7ky4N47VkCnxWqnV4SPYp
MUArAkHzmw7SWPyK+BhllX4lNC6CQwHObuOKNvQL9/fyV3zt6C4uekZUZyyKb2az
Iwm5lHw2usJcXXj6GlklXsxT57X25pvUCn45X3G/J3jIreHoYdhI5ESyBZd1EwMT
zEf6hiKigPLK6Jm3TJhE8NPhD6PVG+Df1lUFDYJ7MN0rtJWqEuHhcbc7xV5yzizS
ctrR1Z9Rbl1z7gXw6p7ImpClbDFp2oGbBgUga83ARV9jWFRtxt5p92bLoojHVdBT
WDV1IHsvKyhMvYNzYRoq0RMclD5wIjzheyQqfV15U6Et3NkCDYonkDSKvRVwPf2E
7wfnCAXa9rYojIP8s2Iht5IbOmCU/Bau89yMccak/JgrJA9IV0kznoPYW4Cgx7p0
t8mDLJrH57X5SIqBIdkRF9zBSrywXth2ASiebA4GJqyf6kmNeiWgLhaZUaGBfyCp
/76jR0FqgwtPVwj13QHfM1okD8t9+tN5zkVk3x0g4sUN1g4eO9bY1eJ8VMJMdtAE
DWwNVM6oFtA+CSeTsUGU4wDk6DC6pPO3qDNuZoUH06VDu80OOxzb0seNcjxRZ6xN
MSxyTYl4bndoUPi2/YjAu0EnJFcc1VlNMhppdQKT9v9ldrMiC0TjuCoUiU1avBh3
VHKt0CKy0uDHdcZcAviAH1hgPLGvl1jP8txDNWQ2rm5knbklyqVdCxzOztIpJ0fq
8xK7Wh7HQSKQTYJTN13GbndJtoqooeasT/UGI0GMI+ieaGPKR8ODGflCpDCGvke7
OHmBLlxLYomnm1ZJYLJAc6vjldRY7UCwG7kly+yIIwoCnIrmJ5NE3QTFNkVF8wE6
9Yql2bBkqxUlt+wNgDNP1fVYpdc8tUWg+i1eAQ4Kui0KIRcZsRVA3zgOZe03Xnss
rz0tN0X8vTfKvhyKsvj2+GYHn6QZAsAavrYu0/YVUZfpMd5xivkx+j8KVnJT1jmr
mMq+2WanEwwlGaIt/Iql2U/PmEJtVwPwe4dMN4FoPe+erLIPf4TKlao5KQq7nxG0
rw2W84Hc2VJuBda1QC3Jk+eD6oQjo5iNt1mfmP1VcAilaaBgu9frAz3FgHKIjoXT
Ah4cjk3AlqnHCYkm/UJC1mZxTdT+il2lF1L0gnBClAQgDfV9j3hWmp/vyZWLkQJ/
pLljiEr1X92RVLJIb9otiuZEfIdHCkTNvIakzInbsSzwCfbHpsJeUbGiIs1cQUev
2dOqdnzyGqjs7IP04dF64pXvs7krT0/PaPGzzOiue2oa1JqOE1kswi8cZCGXRuiv
CsOYhchdKHfYvuUSYN2wSyiGWUIBPVaz6eqfqzr/+fS1LK0YiOOE5m0kJOPCYngS
BP44ZQ/PWx7xzDfXMWVZy48Y96GZ6+fmyD3RmPuOsjrtOGl8XYMY1Rml5F5JSsY5
KlJ9dqaM2S89BqV+yeoDqNZRnTRO5PU+qv/tI7DQm/+ob07TuNxahAqB6TgVjNGF
CldoydIPSUaoQi23Fk9XqV4JK1VGdSUKjiX+HKsNmal2CpXwe5ZtHXNydA259j1z
o2SDcDxdlW1B8NqG5NKhuziqtb5af5L15PMJCIBeKc2WxptJsxlusIiClCuzaEVX
keqJL8mxsLenzZvMoPYYTdlvkRyOly2oWGU/gSWutC1DJhO06b+jA7qFog5ELRFj
EQheSAnrhP9VdnlWe4d6sFDP3Qs4uD/68CvCeSmRRq0cZ+ZqOAOqyl23F092hwqj
buAoo6N12alenvRtt2JTlpCw0+y4X+3rIujvTOk6s+Eh5zbPIYgxAVSTF9vEa1d0
WO4DkHYu3S0ZLIn3y5yM7hNr2JhHH5L21yrbPVbYLrS9nowhBThgpZoSr41xmaRu
22wQNIykYOkBXVwxRDS+m47N8AvzilJjLE9JZ1juiCLdf2OqA6DRl2Lz2q20i8Ej
GThm0qK/sCVs/sr0bU8LDelL9RIzn2TrXZH8WyAZdvKBOX0eTBabVf6ppTWOnpGz
Jp9RbwfoBUkKKAE/J/01IKv7c8nW7oe5eC1lPiA0DXIO62gkqrfGzc0Cs/X0P95g
sEwVx1drs+dVfJXKmf2jaisAyPv32BUkcumeU33nMgJpc/Ta/O/SXtS2Z8Aoz/6R
2Q9eKPMt87AvjeAUiGT78U+9g5O3iSLCwhMCFkkLH0YSKtGPPrnuTFF5mcdd37mM
NosiAuWT9Nt8YujOWbQJxsRvYTVQA11hsuQhMUEU0WvNbumtjyRtGQI0UF9UKbsC
dJGCgn/xoj7yh0l4X1MGZSGLPlowHA6ztdvPaggCUddx0E4M8Z64PPjY8/KoJC9o
6k85K9TcdyogBlcedvUIWXoTPwKHCcnShbb+TdM5BPbwPWYKrPiJZ9ZQV1DoHJoU
A0jUjfi4c5RWsGsvbKFCObo64JZdiRWQL9tuyuFGVpLWRI6rpEh40nNkRdGITkCT
Oly0FEUv4ysUamzPpCnl72WwZMh5jMoHyeoM9/YqXoF5xtWrPrLs2/QLdA0rraVq
CB4bWCnlRX+mKIEYE0OfPcajwOl3KA0xSG3ZxOX5K72N43Q7X1CGcI38okv0T30u
g/xblL0mQcCJkZ3BNX7RRvGgVgKmmi9TzgAdWlMaBYKchD/XW1N+9tyB06132uNB
Xj3r/b6dAK5p+QRSmKicdC0cmcRz8xTqgMahRYojgjv71Nbn/NdsufDCVfgRDK7y
95FOXPkSFoKLbWiasp/pc4/EIN9I8K8lDPHpiJESVXijAqVXscoFpIKgubu3szRV
iw26piK7v9KKKfyrH8THiw==
`protect END_PROTECTED
