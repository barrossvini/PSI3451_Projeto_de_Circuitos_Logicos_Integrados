`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zUsOs1Q55vajR/96QjPIaoQlzAQJMyoDYV177/HmvD58qjEK7XO5x6712StI4v9y
sVxk3e9Cyjrcmc7x0JuAOzpgS7J8xgPmShQ2L+acrhuoKU/CNMteTPkfcyhDXN4s
ZVhuQsUpf44rsVYRBRYkbFZQ1ipXOEwVaqPJk1ZDGCw05QnVE8cOKij19XMGPfAd
63jtgPniTZe9gg4YcmgnLwCyKMzwPyrGHFCqRRudWqUDX24a4sZAIzqaIOfWv4tI
hI0LYozWtb/gZsiAcONJG8oPF6TNME20nYI65sKvyLFZOfrHy8Ro637JDyxR2kdw
LymuguP+pkMwgo3Ro1WIdGyYFFxaiWx3noU5ybrAMWmO8VkQec/8x4T2S0+5CgXm
014ucOuME3duOx+PbNCz1ivkAThouorwyJutgDIbuYSX5ZBJTJ9ZUMWM652RvFc9
roMw80hHrTUiYa+eHkL1ujyxfAz8vuBnSwHr76+kV5fPROfIVvyP9qv70FBRUphd
Q2Tg4VULzyjA6iFss8pxgmk5J/0UyKD6Ir3TVFxZoX2cio6/4KyMlL7asseTH5l3
UPA/kWiOKBydrELAI0Wy4Kgz0gNDv6fa4fF7TSJG9+rPqcHNKSgLTJWTB/rJsZpn
XeV4+kjIA7yzW35xzHdt7Fflmx11riA54ICD0xgFcBfSp5FI69AAIgsByADLu3n4
waNGQorD4CkzidjnBxoLHELlQwHscuuZDyPS1tAC3pUOxZOs/ZBE7RUuw5SrFI3H
B2ov11y0AybfkhY8TXgRZgUB8RAC3enI0AiMTYOX/Ehh2J18vBiKDVUHIOuCZFwu
5Yf/Tuk5NSwo2CHwHxOIllW6X2addurkKtJTaK8xASDOvqCfixUiAFQ9QS446yZh
XA1BpgSjy+Oh8/e38AEvBNNTimvc3J9CfSfBdhMCFszvfzmlIXZipvggaB2mCF+u
cdh+htFgVYW8DnSUNWQBI0SjGNwz7lRnvHp7vv5WmxLCxwNeHiGUWXp0cV3BnoSz
3qLATx+mbQHK2mPJ/o/zPsH7o09dE+eoTLlNxKv4L2Nxy6/M/EX/RVIpg1m/wqSI
ilmyRTn4aSagA93USUW+ipaJ6l7bYxkDkqgQnfrYuTDNZAQNIYEm2t5krTWPBE4w
Y1MbUVuQnCjv6mQWIe3gpIonRituCZ9CUpQCNC2WFhOy+ySp8sblNItTW1UlcNmP
XTXBVI7RubXuSKQE2sIngFRW5NYgeNhXcPLGeODVlhgPMVi84eDnliFJXHRisJRO
3tP2Cqtb3z6exB0Ebxic2YfsHD6NL+L8quhCKFIKlsPrZJ7+pEkBqreQXPpKiEu5
rkcBmvI2WLaAsY/Yb94rSGZ2GZmC67JiLgPZQKD7nAX+YyYUZYmGAzA7VYydKagg
77KQYZDRTBTB/jAL75pu9WV/n9LqHkpC5l6bVl+Goj5bwqwr64r8zJtaLBR26DSP
wIyViuD7Dp6PY+z1hKgTSjbGdmWqr3XY250JDsghAJV+anf5NqxfMaPByXolyzcW
gvD7X06Yktut4oIKEryW/zlWQaadJQoo1Sw6ovTGYak=
`protect END_PROTECTED
