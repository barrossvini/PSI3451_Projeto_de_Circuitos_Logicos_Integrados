`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9uq7EFR9b+RCRhKBY/E2uwHQyF1FlM73OHc21O3Rui6U7oP3+umL/1sUO6y3f2+n
b3tvoOdSqn2+UdpKsAvWRHvUcBvKJHbTfjUJmvekaL2PnRPX10djmcgbjAxfqDo+
vlHuZU7xQJ1NZ8EAUBmuLxuZZM+odky9DlZISpH4vqoBEpWCf2xs3efMtYg0K58F
jCdIjL7So0T5J4uPq1lxvw9rSl9PqNf9APxfcbMcMYbd/22mJzkyX3ho4QQRO9X2
zbEZgaoSLZwkogbj9go7XUUNgl3iNupHIdDlTapsz5wfJeeEqDwhoUHT5wS+0jXH
0RYY6oYBlf/VSAAPFfHScv3kts8ytRdoeRGLU6O5qbrhs3/1bs8zgxfAWd/Ts3Df
0xlTsBXNyh15R7pKMYL8BTuSSiCR/wrur1Z59S6bv6x1Sz3g8JomJ+RCXegjqEn9
RH7DUMlKQ7S9MmU+jGy0eqC1dquf8+BUaAF1oU8EpoTpIgZ3kRUCA4rMm9CrvyWA
cbGwO8EcALCLOjvuxzaWqY5NZzOeChyeeglzuuFo+i3t0tGC+voERLnDmDC5jvC/
`protect END_PROTECTED
