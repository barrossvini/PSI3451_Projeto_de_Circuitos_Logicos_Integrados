`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
29I4FmOAmqRCEeUobdHIDLPyIDHgY+FU57dK6FPOkUih5hkV0fbJS6dLWTF/kYpw
p9ydVfRnbUNBF0srtIMnobtwMi2EmEM1oUv9OJi9e2U6Puk3fzttx7KY67HRWAjK
4XB424s+JF/N7O5knca6uJCMEoubOxc7YqQv+e8VNnRv7j0cWwRpnZs896pAX9Xc
1rBiwKdvzzOaN4E1aZK3w8jFTAD6uC7sUFOlyvv2Fjxqs0QBspu1IsxywBCKq4mK
cTGIx0uSTXRtrBhTqnRroxycH02GeX2n0BOQ2JMVsKIeoo5rhj3+EozPMjynqFDe
ybFONmfIj2MwQZeC9R/zxHGuIFQts35AYLc2U8blesyV0RO258t68D3YI59p+s/X
5vDRedMZ6K7ZM1vfmUeettrNOFWK3bhtCU3g+UZWggoZR4IN0h50SZlVHwxfzx7s
Rdpbj1GNWe0VAcxaKZLppaF8XUdfw/g47Z0uCAlFKgzACQ5S9eSiwK6X5c6zSJD7
YTR/ilYnY8UnzawCx3eVHsAaum5qwrnQPg/ffyOm8wtcby+K6lEmK23tslqRkMdA
H8tADVID3PgiTt5X+M16vB3XrCweu6GvOGBGn2GcSQ1FCcBFESAI76jcUfvDcTXj
beNW7P1cIgxSI1bDkebxVWxOcEjZG8jNm5yDyWs2hOaE4ikq16w0+zLLfHjRDjmT
16kaGl8CrQTFd2RrOsqD01MDLTISe8XbwDh4+6JubfAIUT2M7Yu+LcipLKySW7Aw
ymcXea69L604weStsfT6R9gEAnH/JHs+toZLyDXIz8cZydVIDY8i64zqTDGr//uN
Jye1fdg3RcW+oWeqx9vrWn+c8D/agGXJHm3zlF6VGzvdw+vSZxsJUIg8/ib5MUmH
vYJsiDT6ZVReOYYkChPho8Vx5IR/CD16o3GSzgsQp+0CmmhCMSq8qSiplivhW3/R
kDMJ60qeUTIk8W9WOail112EQ8sbdJRQsSkPUrUEx9Xr7JAJdLOPqXkzZ4naTXsn
nQjez3f4cWYcz4AJ28jfQQ3d3fQ1a7LCb7QnWGwlvZaesbXzdU+EzbWX4UeJVxYs
5OhVA38n+WnSgEGGDYt4GPffanRPR5N6/VZBREMiSTSMWyz7oo6zyeiw6I4UsvI2
gkBkNA7MQ0x/7goPp5SmfjCCmrfsRUfnj4PoC/CwbMhWZ3Ead1BCR1foQ/wXOFT2
QbETmNNOAA3yuF/qnn9srCPx8vUL7laHpuxiRKk3PvefLvEpEhzODahmPtnds++7
2wcBh0Atb5V705JQKlEwCKbYIkw8oYrVdEk6f3a+R2bGIsGaECiC8YbHkBRQ8PWf
9oNRpiLIitNl1x3AWpbJYSRM22HpyYVSVV0CsBgR/obB9qDLo7ErTo9Kbg8bGUNv
4YNQe4h5Td9K8qz4w2dSnF114S+k699XpZ1bTVWdjC3Fw99UlixImVpr7n/RXBcw
hJQ751SwGr3udHl2BgD6Ouh2va/eO4lsQCkcNv3GFSff6vT6IJmiQAMSwkRO+54Y
rs5Oz9D2TcuGBvAY6QRfZspMrIRfEKf4HpYTSS1SHSrXUnMWRI9PRisysHrZgoh6
iN0QcLsYXnwNfx1fSvIsUEooCc4KiEXX5kX3c3i4d66tfIZqpNdYPjbsUSFzRUqm
EDdMDwwSasS+DgLg1an5NnIwLv3GIju/fg8pqM/RePAno/9Utt5GBOECtEhBYg5O
1wHHlCL+w9ufVjYMb1cAFN0Uh8mj60xB4XLjGOqhq16z/wxnRkf7BRS8to3ZkwYS
tsRFi4l5tY+j1opVLD2YpNolTmUXV6SgaJmgUsbmCD7cUbnwzQiUFyc2CW/y5h3+
4TWmCJvc/Kf/1IjqmBcIs2ENvs3f0CPWjHlPZQLL0eW0GonyZ9YJnhRVTy9/od+n
xkWCW3gyXxUOnQOaMewnVSWhwLHdrTPg538scqOGBmOVkI9e4PdCq/wtArF3WhWq
jpv4u8YZiIXlK5cFZWuvN8OmkE4koaL8qT0+PkYkj0ViGlcAbDVx3/wluNGiNh6p
gJ2G9zBNTVVEmH+nCh/SEW/dXEIq/ku3BqeO7Ifw1QLTMRbKVStEPY6UuQXmweMM
OkVREKVsZy7YKkPKfgbOtq2dOoG/oi+vo+YHS0OoykeOvxpW4ykTRbmm4RvKMCpn
WZMhZosKbj1yqyoOOY0d0suQ7nxPLrEX/d6sKO4EWzvDCtvZNmg+bOJKse87mTDn
y77iG2VBs1A8KlfTP6JhgZJYGHyWTF/SGPlmuDP1thmVeoq3cTV+A5z/RcCMgeaO
j12ZAeE4MxQDQE47t4KJ7VPeRkncdxTiRuwWx4haVwVpEh75U9kbAK3uQ4Nb4vp1
CWuHkpJr8e5fGSqkkVN6kg==
`protect END_PROTECTED
