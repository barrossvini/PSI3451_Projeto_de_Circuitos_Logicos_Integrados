`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rNqLeAKLyUEMM8IqWqPJ+HBqsLyb0xSb/7EvGnZoQKFFxdvZH5coFg10TCuhlwvx
EDHk6TWggBMZkd/9R3kd+MooXQgNnIFGWn9r+Mh2+qZoRPqknZVxz9pF+IKDzIN3
uOnaaZofqXdv5U+VkKMPXDkA1c1MDc37lCXABSlZOH7UMBXeiGnYpAMqBuJcsqLg
JzuKsu+SN0pefzYwuA79Btk3BhfpDN5EqeZ611iL6zAz5JilyOxNnC/6eeEuXaHb
4CQHfp+mnq8gFnoRQK/DG57XWxQ3GAdOsI1MkPkG+LJWVEBqRJPe0c8N+8FSivgK
TQHASpOPB7CrtJOnEWYJEQ==
`protect END_PROTECTED
