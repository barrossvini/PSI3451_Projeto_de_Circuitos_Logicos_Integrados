`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Hh+duQbPRTTRhgiVaHjrw9wW5Kou5XlQt63WF4Ov4YeZILCFxB1LY7Jk+VJei8j
1sOIFYz+Ybv2pjQHGs7HO742el0rW0xlM3GX+l2GgSLiAoLCQ6ttM6+L5rLUm/K4
nyWgPXj6HDvQvdEl2ScMAwd75I4DQrU2eTtK+powQaJnrNYyfxe64KDAj88uc3Tb
THVA4v/7yq9nwIuS/9rBJqy+oI65LHgN9LTvgAVM/wYiUo/nn2iXnvWioFFQp3Wg
eC7F7ipXdHMC80Z6VigKOq6h5iuRRfxfO6L+9uEYNwWdhoFZTeo2jQTm2y8sAT4w
wv7TfPrY5ZAU5jut4HpKsllOS5hNM/h3eFP+kZWoJtTcZjXU9o9YIPUk/3dlgZko
jh9Rn4cau6vZXMaeTj2ozyPSJ/N66cquCOsUZ8ooHYznMA2u/3K4QQE7RgtMcCPQ
QMtmiUel4uD3MKSbhs2pvUfkn5RZY8taGFvpc1EQToh/fqwtDA8YB3LMoP6TB6LJ
VSmNHmQ73AzJ2QOzsIwjAbvqx9Vx1IlRZB/xPnNUy0pcy+Y4UUVADaba3HrfX7hS
dMwn7xkcVhqAlxUjJwlKodYx7ifIiGBw1oUAIipDwAoi07j6NquimDxORGLXwRfB
2b1o4vPQCULlIWhAFizyAfjxE6sD4Qh86P2bAXaJD5jGmrLo4aX2rBPU5nWGGcPK
Tmw4Jr5/4dmSRCa4G6CNuAHC4MH8U3mHVc7GdeQqjrL9NC1MpbMJFM+QuCzecX7B
JvbguOnXFKsJQjsOVYJ/n1nJ479Wp7Ovp8b71kDfrvE8zxYMHEBUvfj4d5+ekAS/
hoqx70FljIMc9XUvPVC95NsBTAMLmlAsSG+zFiHpFDOam5GoQ5Ed7ORrfJrcFVOl
c9EqiwL2vFOXMef8s4OUGCPzBZynkmCp//q05yGaJwE=
`protect END_PROTECTED
