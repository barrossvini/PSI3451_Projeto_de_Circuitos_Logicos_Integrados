`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
175YRJ+ZdNHzeNPkx9UQiw0kKkIxx/9OaxuKC1s9ORr0b7+45tGJcNtvFGd1X8w0
eJG2OgsosX21byU/JefEzPihNPQ4EPBt1+0NJ9FWZ4clENzDut76cP/m8jZdhXkW
aK5167LKsCTfIeaLUqUvBCOp7J+i57+M4sLwPiJbWg1swqYpM9TQW90JwXWY9PkS
P4w0Q7DWOWbk0WFFlWuaQQ==
`protect END_PROTECTED
