`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4suNnM52hTwpPi8EeT5w237dZW0BQVaQtGRbMkBGtMfQ3jwRTQc5u9ARefXeK1pR
PL35hLoIFF6cfCaubcLScTw1L9L3THYZOnWLUwjndj0bP24y4DUbGlEvQKEBAQrZ
K/9lcDR1UTtdtTlQAoEomkw3lfHOxZnFkbh9OdCKBIsewf+Y0RYSRu3dBy76LZbj
BfKoqmHOHtNSg4aYahKRwYMJKPQBZTi6P1Y09NudPo78lQj3DOlq6J6TVsEtcSkm
qnD5qswjE/GdmITYbeFNlAHkCDhMFBCyI919Evt7vtJXdeKyAk6Q3PEWehtSbrrV
DioDYmpoV3oTtGNxjVPnsYuVIeyWChlKqvis3+6zr1dw/bpRVrmyhH7HvMPonIWR
cdsWs+1CH5brU7VkVT+3St4r626cFGn91UIjz7tXLDmDBCvL1RDr+FcBzG0ZIxU6
KqWc6uG6telUAjeWFag30zqISDMBoe9uuip5eyl0bbLxfWRfwhLwNd4QqzCbbm5d
vXoqr23rXx2jFIPlAdjQiHY5zHLUaUh+YGnGwnqWHsdequBm+5oONnxZTiz0tGCi
e1jO41DyOzN0sV+mrhEMyI8S8JuQtfsmqE/4BX6y7EFIfFLibBEw7WJz9Ks6BP9G
27A0Pmuga9oEh0UtU+oXyi2gyuB5Uz4e4erjQMTZRStb6lm7M0o369m7eQQLkEFq
OPsBhW46TIFhkdVcf73VI7MExcisEBEfEtkz5KZn3ZwxTA/p8qKkjVcvbp4UOVZK
VQTv4XJtkD2i6hj0EVApxpbUUsseWKvH8fH0B+akRtDIdfiR1wZ3DH9OI3ZhUZAc
5r+pXFX1iKLZsl2jVBcrunNTwap/DX2pt3uyYBuvVBeUDdTYb6kbJvablr+uN7Tn
DkyAhAwjBdABKR7krqKEZP6ou6goLakwE+VErCmTCKNSxwCceTyk7i3rg1G1Cshp
+kNF5C2hzuX/lOcb1WLQET4/ga0kqp78qKUfeNymkCmW0lHahgA+j1iOpmgGiq7i
F3NwCZ1IDegbe5K0dlqx9Pl3pciYbgb30soimWG3+9WVB+RARLjjuj615td0RDR7
an2fxftW/0vtjttNf4xRqwx+LvGaEYp82wqbBN3aitB9qi3WRHNMu2zS8jrFVpM+
Kt2VGeA6n3Dj/KHDuRMe8qZ5rHw2NR+55ROvkdIg0v/aEt81q3VbEZ8laFLGC0E+
Dyu725KCqz4Z2SFY3kfWGxJvZqlW2lO7Iwx8P90IHust/+5zjnI5pFwdBhOPeoWt
QG48NiHa3O7D4Rk8wJHpFH7PrpUf0oPtmChn8riwkIYe8WeOl99+gekasTY7VfBU
aB6+9+J9EANfnxK/Eu2l/218DmUB82b77C+3AjZ2fP5OYH9/oC4Nu6Peh18btJBX
DZ4mkpGDJh3QUPX8gS1MpFkPDb38t46EjuK7h3w+KZCP+dcOY/XA2ZW54WYN1E/0
vnASIKPD+DDDBirotXqux/9+lpU5V76WbiL02vM/cOf2NqdEoW9bSXjrr+j+ymom
okwWNL1w5eMPfaTHhdNajU2qb9SMLTHvJaTL+qtqg3UbJZe1cwMbm9yyiupre3gb
/vGmlPUuJ/49MInXEl9xHu0jZbL1xBrYa1CkuabOP+FfZKCN1/3zL8W/NLDNWgTn
+21Dshtm7wbWdyQt+ShK5jRFI3gvL8kswNZDm44BFTAgPpKsGC4Ia4jLHDnWliUS
2UHZ9djLHNkVllbtBFaSAH/rS9o5nVwiNArZleaa1+WyxO0GCrsbIKsn2jc9K0Th
eM/cgpCFXLD3bwJ7E1+QiYX+TsR0VYn/7JlUEjZI71IxrYya3nYG+wYMMOUSQChD
BPinBw11X5oXkzf+sE6T4kpBYq/kTqua+I8eziDSKew0nuewip0WfxtdjoeheY9W
e/odn27SZ759GSz0s3TY7BcwnuZiONfucqw0b7jkkPancatRjHLyNhmZ74FKrYRx
rBeCbamK2JSIMe2Gi88gatb85Iy0OLNCzO+GJicnc20hxLF1cbxV+ETLBgkVQJvW
KwgVnhf7ozMrgnMbvR1FhbQSUzYUweHEBPypoq8gMs8zKw1dl02cEBClapRL6FEm
P0Vl/3+oQbEdxfpidke9uVTWvtCTfnnFR4F3Ds7x5fNyJ3JQhNSxJ/yAfOh8v/IS
ire9lAvZSfwDVpSwJ4EwoiSw9cc7FtCT5CcDh50/o26eA6peCXCZCM1dgjvQRRoU
7CRI4IJkMVLj2SQIm1gr7ZjI0KDd35/G25oAEgB0iMzMZlETfqQcwZ0zaMG1K+w4
5PtdbU/Wjrp47nEtI7CF513+lt9h3wRf9W5d6R3kYwiom14giRKICV9D29c/hkMp
LHd4jiSeuDXDFOKtuJvKNRHURC6ddUa/Hw9aaZzVK8Ko5M/zQeiG0hzmm1hqZnnR
2UpbJWtUEa/Z+Llf1DiT7ikLDNyDGfhLHPrzEoS9Ik17TjFzwhSE7I+x5ZPAq/lF
LSQ2nISF+znUpE5hzg7rLVOwEC3emXu2vHBUEtdvl/D7UN38lp5mCeOUsop34x2h
dO0Nxd0PX5lSK0hrHRIZTHVewwiJsGQK1resCDLlw+U11bijyi7kD2JUEPBEF3aj
jVTxZy6LNJmz0ArCqgwMHRA+DXe6LN9VQP98mkyw3+1348BTLzpkYaIanGAqX0RN
PFGKzDxkGqLMwSi6R6v9fIykQpUuFIDyyU0VwP5m3D7v9RxwJ+DRYNk6slX89+c+
g6nLa8X+ivWfobIvjysDru2AS7WD/gDYZzPJdMyTG/Cdx+RARrPCt3ZrNYhC5o84
a0OM/ozJfuvudBsO51iLvjzlItsZrWXFlh8IP8lHhWtqtUHXwLlz7V3becDmrZUY
QobHmeepK9j0B+Hubg1tx2Knw0TlHr2Fktb9SYP4etAA1qbnT5R6wyOgLOv1JgpY
DE1ZpKL+Q7XZzqnKcGrD9KtAQxeFLE8glmnki+GSNmmBTS4BR2l65TtwljAVCavU
7XCYVF7rUt9D1KOf8YfAZOb3xGBYnCEayPiW35Kl20IGRkb8gb6eD04eDnvOxsgZ
a9sfGYObYKK9gPNurN68iWwOBjEErGcXrgoCspEjXv9PgqhXBpWXdOUlkTwflAKF
o0jpR3cJZRyEGa/X5ucEx6LEFutzl3ovYqqy+5FQPxyPV2UmruMg9Fl90ZL/y1HJ
qNsY5JiMXKlOHKBmXKbK+NG+cdVvYCntE/y1TxM1Uifdb6b613+ZGciDYwy9dtFR
3Ua/Qrxbw2R6WVnOJCvpkj8e6rbZc5+NVtXzzfHdAja9k8x9wQYeMaNwJST27I9G
Dg2FHHo9tmd6DU6B1uYTJP5sXDWD9mpAQ8sFW9XaOwb6g1f7mVUlP32i6776UFSU
H1tEEKlyUhuK2E6xHB7fLKU7/pB8nHbvyGzdW1GwUQqhsri9Flm/TsDMmFPDQ4r0
v7BCyX2nohmpOoadR9c2+vLyqFc2LhRZaMC8N14n805RoJvzN5H53w5aTjFhAKAB
uCXCJHZh1pYT+dfMy80i1EEbR02EmQqJ3EWaOmTSAr7j0KtsjbMaDVCBQgYM0PVk
7paJzN8AcZ+1UmOehgUmwjsZtpt1LgVpZhmhM4Jq+ViuHCb4WWpFpDwJqoEBtx9H
s78BRZvwx1t8gBqjSDyhFjZu/sncY3fkkuLeSyN3YqctURiJIi4g48z9ktK6FUf4
kQlDbcbqzO2h0F3elNXFCyc8egwg8mytlm0LjZUWv/yvQamWqQP3QA3BzC5sWNUV
cElQmkabR9ZWS71XvgKD/8amvXMGYeh0MM3c389rMucYV1MNjYfmvUtVCtQCqhBj
YUu+ozOs5rK03ChmD7qXwoYt7z+H/rWHNfjVUhKesZqWPB4e98iXolu2tsBlzpRk
NAqsC3jm09qVVlg87QHT3pVPauQUxx+Dyhk19K/81r6762mAifgIiM9iTuLxy4oz
KeUk1tNU1bKMxKBFAygKzzRMKH5xrGL+pg3COwzlJckQL70xAOMIFS4tOGnTRCcJ
IyCveSLSqnq6aTokY0AuDyVq/Kqtlz3UeHB2CFlsTw0LH8gTmeEL0XTbIEsb7MxB
lkUEdySm467g33egon2AF1WfVKeB99ULZJYlj7YQuoe3UC/iGfw0QQ0+LSntX2I8
qdSsMGCVTkLEnFz6r+zC6+TpzwshJRx2e8GWL4Ofub91YyBvWYrZDGiWBh4axEgG
2ZAQdRBpKu/lI28v4u9Bm6I0v5I3jT0HJPSFkuJr+gxZxW/Vvi5FwzpALQOaMsUg
pv+tagHo+734CyGrtZav7V/RXnMw3pOd9tvT0e15TzNJ+6OaTh0JKFKZoctoMg2K
BoPj2k++l+GP0lOPfx0zZrn/esmcFv86VjVWy2G8FWdn5P9KJw9rEd0Kkmmy7U4e
ImS53BzB6bv6aUyzPhTk1Lub1K22ZqrIWUAA+g47TrHwxIurnvHdkZlECdUT6OuG
Td/U3rWvqURREbrwXMLtkTjbYoxanXmf3q5Sp/uDW9SRJcz28i6ozYgrY4avIWBY
jH6AxJeLvkEJGMoTBb0Eg0vl/Um9/+ZXyRXENDd/+OS3xlXuRTW2Ip5ldUYCcp66
gtuIhB+W65aeyPFnVkRGWxC+tDDUDIqMiCVIIsEm2SH3PaZBQYGl7CIXzXZUYsnY
nnN8QhnilQ4OWbx4uEkAjQX0uKLWi3xf1bG9ULg8trHGn5dC9EfJAuxmBhqe9S7e
U6pYV+61skjtaogXp9tBcnYW2nSXXRMGjcIlUCRbfw0gXIt/GctmOBFxizEIk+aw
A1unr9Z856f6LY//ur+T0EqVPRvQlcuvnUKlGuiTW7nDIfq9dBE4GUGG7Amp4Xuv
M+os4G6UsBKg11e+F5oTSa4K9meWZLb0+eCOGxg+u+G64J5WZ/Xi/Ca80Sy6+fyd
NwUeL4O9RZm++A9jJaqKs6forOX1K64p79DkvD0rXWXv/O1IpoqJQRCYcWrAxonz
JKeU6h0gk9D7C5iYqIpPJ4YlKv5/+qBVOrwCy2oh66+7QSKEem5N2NKP70tN6sRN
MnvhKgIGiCMHXJEifPVxQumuR9Og4Zcfzz1Ko7YhRmbXFYKslLw9CVmYJBqO+oS+
zEzjs2K2BOwjKRLEnHWc+pYvrFU1Nmo+OZZNz1dfsvV9JeDFmxQwTcLKryyZcUR5
FlL8H0WWWvPnp0GThlDdrdpUKhl8Xpgm0AT1TsQr3kjW//bADDjXa4A++KgDKzm1
UT9EWu24KxT06OwoeFQjDey+UUc217awDL6eOC566r9Pk7w+EFy9gafXBieVzeQY
GOS8veHHPnKcBH+6hy1vPbcwwAvGNoEBkgOk2OyhnQt1kxocSSnRuP8X3SlGxKS9
uFiPWgMr+L1eojmRm5eeut3rWDFid5PRGxNAm25ezwBdYp7Crs66x5+Ap3mwv0jY
YpjAshvk+XZ6A9xL0t/Ec+AljuIVwkAlqbV5ZhOHRq9JlF/A8ArY6MHw8CY7N/cF
CkVqpOK1KNqm9vFmdg4OEvQo4tu3PHc031mqJ5xV3tkTgSZ2nYQu+SsE2tcl9OQg
HCTxlrV2hkV2M6W8xGg9Jiu1Xew5i24uR7DNQY+8QsYPHzEHJF3yT9rYC+o23APn
np2o7MMuE1k8wrxVDHc6jR5rzdfUux5R7101Gt/AyPWIMJHCmgwtSeTftiaAQbrY
pmiQP/bI7dJc6cALPnozUzwJA8JsHMJ+e6zSl+v++AR2Qu1pcJEyE1DwpOgHFpvU
5zl0u/G2rGHkG/Dn5XHJJNFusmlQHoeOn4E3GRGkLzS87y7CrkOUR+ujpmr/9Z2q
24T/C0djDY9MnpyzGmQ2Mn3dcoJu7bAotqY8ifgsrEYIQMrYJVM5PsQoFTgL0inC
fEq9Nhmqcqo8CU/UdzVq0o6/yYgDK994ZgH8FLVz7ft7s6zRseciVFMrXdviF7t0
oCGNn0AjBGcOulPn1P0YYq27f3t3Wl/xvfoEVDDjDCIMRz7RFAcsG04WzIlcb4ej
U7EpHpx8OTSyi75S6WDqPMsdcFR9YqlzjkOA2GwJAtfPaTcPE+QejVOOTGXkxMZV
68oDmrR0zKKhGptadFdaSjlXJhcm3V35pQYXDH709Eqk55fafqMX35GglTY6jA2J
0FDvxRajTWDSD5yJgXG7y4phUWqebGbLGNwrPYom9e4frTvvRN/S3/+IDk0HYXPM
WjCyp1QWyHHAcxxQQwHbIRqm6M/cQ9adopcc27+95oU7gzkafu5GQ0v2QMyyZY5q
RWGosiGxirZK7tZQ869i6Xtj1ahYoNzKVCkJvKSMgSViPy3sMvDJM9MSERCzx5bh
Sqt4JXV0q+E30hZ1Kc33E4SI1+2rnAAo1CpiGVtqk+w8VbrB8fREiV9oubM6v2d6
6v1AsTicxwks85P6jEfgeeHM2M+j19Iug+5h3GHXf/U6/Eef8QJvY0e42QVYvoOi
cyW5ng4Hn+2UzGjxr5UcqcFLR2V9uu+DVTFcGL+7JJRsUyNPiuo+OuyPt+RpGX4T
S4uWF+gCiAqI2le5suRjEgSYytVgu44esdev4VyRGZ9GXaByBqvNDYcslTAEadl9
zzNG55nLWIoh79+LC75O2ETJb3mtbNYI9bMctcHewp9Ta4k2NpL6hOaYrXLddLEK
bf+nR6+R+bUasqjoBM/snA0mfUD/HGJ3NPwrcc+emPFB1FqNNy0CHttAOLJ8qIX7
jy3jG2U7sQ/P6g3R/9rgfh0HdhHnG6y88PPzlfW9aFsh0wnZ4wr4P30WYGbhXFyS
g8/xrQdvGJnsRaMk1i+u7N+AvFeS4rXer2OL3ok0X9SWQPPTv353BYgQFFXUVaRL
2XWQPqKK+I2Ur/LbwpGG6dC8JDybRftZhzaxzqBQT2P1D4N4rh8bf6lR5iRRCABj
1ECwWr2Hu9Rg2mjQ3YFPQZHEtIaFbZLuCxUSAxWRlei1OnuNV+p08/+jCzz37BvR
8Zvv+cqvOX4oovzVKlMuqgVIQWbLG86Zari25NmY59oNuphyoE5gtuqwPHnixPVo
fuO87EcnxOW14oifgJuSaZaSLnAiOAEdSC/iMh0t+Mn4gISZeT5vXG3R8qQSNIj6
oNAeEmChuZmJFb6YSHZs4dChrcoMM8tunvNzC76sixkEbl7Kg+vSzzrAjJcQEkDm
oBv1PjUV+POR6XsUD4mV6zZ0IExZq4tPXQj2ReISbNHr/S4XNXKgqAdgm5lbvcDR
0KYaZiw/Xox+pLlRjaiKI/J1y1YVoPLqsdezPplqZHmjC2swx8cbI4rBajkPWQqS
hJwC4VbX0+7vZ8MUR32EKr440q9Y7sxJ4HwEpTyxJ+opETc1SCvnPS8WbdWTlXvn
YplOzk7Jj9iG4R0rN2zvo2t2WVER6yrtYUz6UjN057+5l/GHOnEtwmaaGsqlZlAJ
3hERm5PS8j7z4ZXdgy4CO5Ktuay0gt1TTrG8IGPOSQHmLY7d5ddo0DbYk9Ua/LxV
TC13LONTagWfyzAT8XuUW6kPfsk/JzE9Tz9E6HA52UQ+HwzXufrS712r1/vtqPvt
Eh+QgESSEDTcwAE5fMHqgr/xBy4K7/3EP63ZHzwn+/eg7hkffz87xnMoPNOrDC/H
2GRLlr1VR7AjpTJGZPNu9/xpHPBeYr6AOe7+YzMWa0fOg978s5+Sq90GtApU/xuG
9iaegdJzV/LwKwZfyGeifHcbgME66AHehOnP1bD+TRD7XtWBfN1K0MrcwcSgRz4C
A3o0rmMOgwWjKQES2RVNLcieXmE9myPz0hmQ8WxtMACxh4g2kLoXjR8LI78Jb9Oi
zpWSl4gluIO5MrmmOcKS2PAzoelfkwGJ1Z+1pq6x8GbszFur318BpBRY9IQb532S
5zErKhijqck1Ws6WvHICDA9T9E4pDL/sUy6MyVBfj23HJZ80kV8x08msBeWgwp4K
UwMYSnvQTo1GJbcTPaR+MznwIYH1QAAhtqWTX6titkMH9NmM4jpxRtv4J7cqavcE
vWPmZ2ZFrPpmqYAksU4onzartyZyvGWTMuZF6hYwt/w86gbzOZS+F0RqvvR6nMIh
XAFvz2Rz6RtmZEkJerc+1B/cLazbpLYi9NA4D4+MMs9iUVub46dAY3LfugKLui19
zZUj8SLTIXFWNVMCcmuqrWjnhIqxsZA160DOv94O3L3Jh2cPQrXAr0ria7zqURE8
IemupZcv7rJGVBzQXrdHSNLvi7y21hnKyCn8fXzSa9UvODLJpacwXGppMWJCspZH
qDSiVyZSMOj33O0qoD9EnJDzMnOSkxIhZ04xLjQok7yTQtzCeKeiwM2SqNuFiDXu
kIq3h2PmpZj4duqqNZibTdB5TILjZUZkdZtIOjzWxvseWfUyWW9N0EYMfeBEMs3G
1hiX0aYXJSRmPhD07GjrmZhGjYJ3YOrrm/gELQ/1hIPXZE49w1xMYwoUSPQk0B6Q
yuFbLjcAamg1WF4b3c9KisbMS/dyYGcJzCM3252iXYmBN9DrPjr1OVRBdNZrsxJJ
sJ/LyqucHF+gx1XK3wtuvefAoyrLaVlnCDbZp0bDQI9hFRebx/HtGbjhrrpA2+Ug
xdij6jL+i7Jgn2q/VJ2ikw47vBDjz/ttXFEHtccsDlJHaWyFzrIztu/OsnChNt+g
5xDD5+/bcnVpEB0UmIV7u0p2eEX6vUHSU5vfxFoefWFrziKYBXOEwQ955+crybbX
E8cBmnxztQEN8wN6VPrCRL/AaxWk/zGTpTVzA/ybL7mEz+rW2IX2Hea3xy6cBg6n
Fk6TNgSAsQqAYhqtNXnFqww805TyEBH8WzD0rjGtApoOgUWHpmX4UoGn1+nc0XtK
X8YuMk16VuNvmfE7fEDGH0huXOxyVgdmGXs92asFgENfmCNV1TIS4G8QbNOrjqXO
X6MKTkG2kp/EF9kjc4m5MPw/mo5bU1/yYxFg3yh6DM75lKG5goj51QBqTA5cOwvN
mhsTbA4KMV9qWkUnf9rV1Yc8Q2rxQKqp/SJZSVrmmdOXgUYdKAyapdEOFU2T/JVC
wxl4ZwXCGWkASSBDrcRnOkweEThMBJ7wt/ujPn4heexsqF4KRZwAxJW7lwNmsxRv
MDw0nGJ5s9qivyn0dHhfvgRKaznYuMXcCBYUQZTdeZ4GXSwafb/WCL37UD6jA9zZ
SZULJCb0cedzb6wjoeBhb7cJNpRfTf0TJGDtIVHWePQ+lC+oult1RL/tfmmnKMtW
IIfamJ8G/zub/yaam4wmWu9bOsN7VK4ncqboDCP/4Jdf1wko9frGUmA8ayYVNkgY
Odn4fd7mSppwKQo37nwdrMPSO0Jy5Uw04QWq8b215BW7PI8ul7wDSvUndm44QK1o
77R4gPU82UT4clnTC7U9LqMI/Flin6GBNK3/2hgloXCX90GNTPdv0cDhmLvOoXww
nY7EVfH3nSSCF+D73nUX4NShE+3nAZqk/QFJZ+/ft1ShTgV7HpQuGVGH60TpIyho
j+mlMG/rxj6xNOIczVdcCjXncoDam4cswReJ3Ud5f5/LVVgXmxcX7Sk7qJiuKDVb
iA9zMYXKG4itw2u8uLhSYR4vW5vIE6KdbQHeaqU+NCgGspdWv/iYBoh2U6Bi7X/v
967lRt8lBjXMjHelqi6TuEFkWGxCXQUZ00qwkBd0wr+36FGV9h3IH57A5cX7s9nX
meNYJCYPIPnonjNcJpIxpu8icUysr89HnjqDqJJCmNNKKqmIg6ynERUn6jCOX1QY
4/1RsSooydFwUcyH8x1cvcnmJ4mdxQdaTaOQhudBJZdO+82w7Z4VXL0O6TWw6coA
o82Jxmt5uINIU45APKkZw3R7glohdGh18wPgsxKkIwBNoiaFLx1jPVWM6tQKZjBS
4ctAgj7B/e19+zCNsvaCQbuzBoZ8fGs41audoauyRG+130JlH3UXHordWChA+NYs
QIMlzzGRMBKtwprkumxqQNiRV1Uma6453mTitdgN0OkmnF1waGFpSz6Bug1JM+cf
cCyMhsSIt7foI0ROupjku7zbP0bhmkb3LAE1G6HUk6/ng72Hn6tCrkW7LmPbkSeg
KEvFQGw0KhEYZYfC15BwHZHafllyYEZtmprps463WXutNqR9sbC5QMgzC8ikpLP9
8W+6Quo2yq1oiMSAETDRn0JL2QtgXMyD/C+agtEzQtirN+j+yjswblRQB3jKXHQ6
SJKbi1Rjuinct6bvLR0m5jadKnpgEsFbw7H3B+PUxM8ubFeMxapuACq8upjbN/Xk
l8l1dQDKdNBs61PUm8lQnMbxOiBIcX9nWefWVFqswRpCVgdBhtpu+FISWIsHy4WH
McTwuf/i5FlkhpRl0I5dm3KAqoI14dampVOjtY9OLfmGRnRd9ct+lctlxi1Wc/T5
SY2iCfI3eMH+V9Scao6dSwt5Z3fjUDzrUX6twsHdp88VRW3Yv2ZotlTLHsXCoMn7
aU0oUqqB5xX2Qv138UFbbcsqAD5hXGEqmNy23T3gr9cRzbp+UOkfsAuOLxfBntFJ
mCvpDDXhQCId80eODkBpz5axnn2y1JRCyxA7gHDrwo+jlfPGAi7e7P4XQflrkAon
i6hLdpn3gCg+F+C18Kl4wagbeYXHKwycWu+GMIafXQ04jQlOo5Bll2Ic/MOMt++v
QKr0jrhhAZUHeVdu7T/OF1nsdHSuVzu2wh77bsP19czzzgiz1jWkPITFcw9jCs72
CJCjrVcrfPzpbU5TmtGDLJVKTp8akryWvISKpLZMJh1812fCF5ig9IzHcbbWOPez
1ybK0uVlYVZoJTrppRC4OhpuRzjFsirkv/229sj/yBfhDC6jw7xdXD9oGQz14zQS
XEyrxyvqX61bhayr+vM+kAwW2G5JlV+Ske8KBI6VwTpMIOv5w++aNu8e80KQp0TE
SS/WjTIRBPgElhBOh5r3QB5CRkuBhm0cpl4qrm7QUxzXrWfrtd8eKVMiHT2sxqU1
vN2X3q5asm8LNiia25m0xwSulM1g+ypeuPytcElyIhBHuswcrlS49QCzcGOY2fhU
KKcimGkhd0uJ071UzR78egkHtbHO3+TS/gDts4SNwuCfrA74KDwe7U+jBhALtvvy
WffiUkEHlF73/eqNUNROo5slUjyCrc6NwoQj+Wiu/+JNuAlbuikHBLtCBv0iJlhX
o6k7WK1+ytofAgpALVTv+OZp6qCK3CqtkOc8oYRBhgmaTikw/DqJ8v6zmVdRRhmT
2eB8mGcLVZYlCTBZv2DCAgtOT1d0k3RLK8ZqOCcbpHFdUreAo38S78FcYuQKXg5o
a1dssnSPCs5Ko/pokQX/dk9ocJ76JuX8ZgtWzxJGuNwW8p2TDA2erNzIYJMPnBU/
eMim/JOfa2peF9LUpyS9HcKyDLhy7MzBFtuCn9eFaU/Iud5/mtxg6pOa/d2hmO3G
HcoY85r3snGM99P2oSoybSRsDMOi4loUpFP6oS0L6jxbNOE+rZcCEDYvdDMFSc1v
HeFluIGR4xDTTR4kw2u4frAlf/adVkfBi0J03X0+WAsmT4/vfVn0ceRX8XbIEsVf
774yenFjhkOhS3c6OZXfCeyrCZjS7oufKT4aKAN6ALGUfWnwOH3uG6t7xfNdjYLb
zoPreks3pKlaoowD/7p9SdLvNYwdYK8GcsqrzlVJxAxrrKSJuk2PSvVnlnME3QVh
eN1fW2R4+mAl3yrIf5DSMk6M8dKQximIXcLS8mQiQFviJIyYLTH0JEssD0kDjiPh
VUI8jP5zpSrq4RA1PoqKa+hIsbvTF0dIJlutwiOMWai9e4u9ocVDzmfEOnmaBxNh
iW09Hi7jfGmzoeCEHBjnLn39tyE2ntGNxoc7Yc4XoU5u5KzIwtjnnz5kzfMkzcor
K8idc4VVw0fesFlTo55ZPxvqiC4oaB4itdZHkUc5tcZchPK0lUwpgOxT74dJ0X+D
/iP96SwBMJPS8rdmzE24y/WdzuIcszOGXWmv0Uu9MEIyVuIOEepDW9ZpvZ1VGNcU
H2yrOX642F05X3LH2Y3Jvfy+wFUTnBM3PlIPLNuDsN81gpvsZrv05Akzeia82MRZ
LtQKtmxIOwYlwfKLRqPmtIHS5X21UwrByswm5o8KUrvKgDx317s+vHmn7XYlzJit
EvmMe5cfjcFl8HQORAXCoI9TKo76SeHC6Z6v9JDa3Dmmu4T5USx59fc9pfprzSgP
8DiFdtzXKyjQpJENDpNSiK31vZk5ipzEDozdQ2IKUc/PHHNbLaQQ/ifG8cPPbQZH
4ysPAhzkABpo3lJMSr8mGodHww9PDL1mHb5owFknWA/TJcSSbzC+p/88WWqP/05I
VkSelEoIm9gzrtEmee4jmWDHwetTmf2cL7RdTnFATJqIMnWnSGspte9kn37TIDd/
7YsrlvZCO7jL8uaWrXDF8NT6ZZNDggGU16gE8So2Innr2BWZXmSNE/Ep2a0DGSlr
AGLFa1oAoJL3urYL8OV1IXyd9aKWF1kxbJImDikiHmMWRECBdRTJW7bN4DzUGoc4
5ykR1e9t4H1eB+5A2DzRBeZ3a2MjQrrCsFY2lNVMPTjrDBs3Ua8Yw6TVdD8xh0GH
yxXpVJJ/qIh8IwEQrkmbleSDq6XV+p4h16VnnANCj5DgRf3QxMNvFT8pAabTvaC5
mH+Kaj1ZtFOCtQ7sfi8ukcgKwIgULkWRi067cPU2GQFRR95qnhQ8GmYooomj3jWP
cMsK9Vjt79Pr7kBCn5x3CPlsQ1uQy1ywGck39gtK5JqCAGVHxletPSjtp3VviOTY
h01ppRo8RH6CfWL3L4Z5R7YXgCdOHF1WWKs8tdBVUwENbZxKYcmiIi4kIAQUoFlu
n9PKmMZAmMy+kaRw0oZtRmFY4PSQjCkhO8jmwYrwl5Xnbc4Iysa2Q2kp4H2XT7Xp
/eRCYL6uzOTANL051lqfse2/ZjETvmazYp5tY2bzO5ekDwm1xD9VAtc4TQkz8Y67
486J92McQaqaEXPbFvb4VY2T3YCSPgG5PX4lm9Ozaz5uBjQhrALsZ7Lpeppok4WU
4HDKwakuTpskumXpRJXven0evXbn5Nfe8f/EwjzF64eFJmrJ+L8p8g+WPJzoYW0U
nIz3NRvV9uTJqLv94qsE1CiUM+89OmhoqG9j8CwZS+ovolTQYXWTU4yfb3hm7w6e
XQKaPok1t64Gwv840kFGeeTQfypJCqN4kqfnD/A1sYKgSTVuOQXRj6nF3kbRm5k9
hfAnMC7/KHdPsjWNQQSzrHimh0BuIHUyxicAlICkHUhDe+biZUA99/WaqS9yK9cc
u7vTEmtSxUaoY3LPGjHUrAQO/Xkb0h8N5YHFa2/BXCES5EaF48d9NbldfrFsA8pW
ZYZcMmwO51u5esOXQFtgRK25mVesGsnEtyueWhTXc5fgDB/P38TeRuclnTkMVsyT
UdyB3XPK1snFf2IQQq8UqiEHzcXt1PaX4O7qgPrAUhkUL7+zLid4mv2KsIlADgEP
FChDgrqxJuHmBw2wg2aRLImMe5xvLFHrm/Tw4z5wsssqk1AG7BHgRf0ybt5yM8Hh
c64WACABJotoDn1/jWTOewvlQYKV6XcHGl26/aCGHEpaIH6UBLZ3SxNLCJ/asnWp
gfj4wJinapbGy7oPhR042QwAlNVqn7BDsm1zU8fGO0RE21n/89umrtnmuvCv5OkZ
8dWXRgdk1BOHyR/JY+xbWhhRHfLigXAHhamTe2hlFBYm2GEtMjf5Tw6tEwHiehyl
j17YEp0o3nFHpRUzsHCpyyojDZM/Az33VWV7s4uM9A3r7TPBV1GHPpaBxeVfhBsx
Ndhuvjf6N8T4lE/oAOZIMxwDDp18TnMIxbnoO1xF+ecPPAwIgthqoWRt+0xBzfu0
UfGudJxj6GDZUNk11fDztISPNmF0kSm10XJNd2b0lZVebnE3E+zhsQ/EZdC8m2Df
GeVqps/2L1OPD4A10cCHERKtGBv/6YKpJDO/L5dD2OKa5b+shxjJNg+CtkZAXL/s
2TCVsG/oJSt8NwgoYQaKtsmB1EHxuBa5rAbYZoRrfMv7IIFo8fkZD4XimWsiMLtg
W8idFri41CZ5d3gXIsdAbULZR4GT6Z4JTgnsu2JFGK1lpaTqbmTCkxN7Zz8T2Bhk
DXNrmtqh7/jJgrzCsRGoq/6fMeOPiIJu/Ce5vyKheyUXkod8MA8TsnHAHkW5TzUf
UKGXkGB22xIv8e/V80FYMlT7uObDh2DashaJMfW0ECwVolzchgnYQBCoGa3OOJrM
s89afINV+NsQmbJ+YpaH63nBIaD7R3drj3qmtu+RvdU5uMYEp3Lb0k7Zum0d9Btq
WBqr18Qf83QCdUbBJeVjJUKABYJVplUuzaKiCpEDN7UVW1Wr+v7htTw5oEZhq7LA
O8of73wE/eYsTD6tda/G4xxDdOQm7Swd6oetWRwxbsq2Oxn5Y6WQlAZoNXtCnCFK
FhpwEpg+pPEeuQTjQATojaygQYHEstIGOW6jgQmTR3FyVKJqkRdjKuU7qfrS7O+r
c1cNegM0pvdqZ9OWUzgFy2JJZQGbyT04T5lHnQY6PQBsym/afImzut+LGvo95Hhb
WE2hUEaIWYYZzhF00pqGTo27+aUkDnl1GXXuad5lGOX/P6dYbrcUUDDvN/MOufoe
dzxDLUHvvr9t65ExucF2XZD0zFVU6jp1Z2nponQUMO0dz+zREjbA6Iw+wTXhOEVA
uzSjHMh98VZTqcuIX2aQvd6LcDaC/CAd5k/MqLtIxvKJhrC/8lwywkO2Mh3LTNfL
38NKDyra43KNxCS2AGg3aOsBXqNA+KWCzI9HTFkNLQ6wx6HUcCtVEVlol/ZDt8fr
KY9xuKsqdath/s5L3ef7ay2eh4jPR3air0Djdw37iffDZNQdzbGy1fCqrVdUYRVS
3iOWgUrJd6kWvoGkDEUFBsvdd8CrHjKXO0nl3R5kVU+uf981gQgurtu2vK6/XWNI
xKBJ04YIQ4UH3lf07hQecCoy9zTucyR0R63U6zBYlwssGpbH+bJ3zHTFvadRFQIp
v3oHE5p2lF9YJtWfe8qSbntn38Kn5b6yCb2JkBnAZBdxfYUA+KfV8D/BoRcrRGO8
8HyIXEpQcfZw49W7QIHcyWbQIpCi1cpO/fKFwC6+o60dqu3rB0tiRnIfPBKUgxNS
sJ4qudXQywMU7D7AUPT4OTc0D8Z3B4AryhxIfAmkohXav2w/8nLEBfcKnP8YHm2s
ih6wb7Y5J0TzjEXZhgqbc7ifJ8ucupnFueImCY2dr9mlvpawR/RjBdDsSM4I3HCu
CckBhKmPXmF/JxOThU3UKyAooC44Yukb7u0p/jDzrOtIs1eAuQb+d9seAzXLHIAI
icoUdhHq6S5JP3K73fZ9HOMTF6C9spCNvQlPCNIPm7CeUycL5Om0hJPYVdJCauSK
vbSbhdeuY/LUkzhit0EzqxNboiCfjH9pxE75qyl3kIMPImd6ecy3nqbztDN5rp4u
jVHwcJEKN3Bge1Bdv+l0xMV8ihVoUdG4lZf0Gkc8B7nV15Va4O5vO+CbMDDNuKZ2
F4DKgpDDJWY/GEOT4MwBJVBfH5hC9cHI81b/b1FGNmWPO/aBZBk/uNDIaqiVwXHB
V5T/OJUDuiBuAzBDQeZBBZwTaQgNbvTNi4P1Wod3HYR61I1fSS9Wv9j1S3RYW3R0
VtapQm0mBrtmdaiCBhiYA0krnLwuK9YIKyL21WAprnVWcs9/gGxsUrewsF5Gw9uk
xPOjL6YbyZ12bTc0gUOeABdBdk68r6CiRC+7opBVOhQ=
`protect END_PROTECTED
