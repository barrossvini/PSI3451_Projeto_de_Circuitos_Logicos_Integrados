`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rasXyuKCWXgknE0/b/wy15CHHDwd9UGa5kMLd8xjEQb1DbOcwg+ib4BjIKcRTkcr
jGqwEDvMP541B/hnGh513hUvTCytXmsabJPjVFgX1JYRgC49f+/fXcMHTLDE6Jf5
A8Zx1VkahsLrg3mB9AS8eyg0tWjAqnhPDFS0amtrKoST/GWfzxZApik/b5wWo2am
Iom99nqnBZlsyH3EtFqDWWWCF57cZkb+gyMQD5Lh6+HOlXkgJXavs81J9oBkPdNO
kxbRvbGwIZoxOAbdd1fCbrqla15FTR4vTBFp40BZzWuMqylBiHY4nl2UpNb1skZL
PdE/zG+cFLbRvDTPBeqPWFCjjtNKJV1eonbn2WHO9F7nRvfAefXx8xo0HIb5DZTO
Gofaf+ToMO3oY60az2xUzjQn+F/6LsEG1shRbqTKJTPY5uOh5J9FLa7qiFhwEwnJ
NeBi/iHXAAGzfb/bfRi1IBl+hV5IVK99JIGRbK6arRB0738nMuou8kq1rJq8h3LW
iieZI+n/ZieEWZw0B945m1eGFGKBZjn55TzkOOj+cwRI5IkI7x68EOsPjxGY+N+r
0ekMtilmLnqRisB371F6ENKsO5izt1T16b3WP7lVPUZ8dZfmyVjmR/dE4Wjl0ndY
56YlHEUsjDdkoIMc64WthB7BQo32R+9ty/rHWf+eCdMruk3criK4Zpxxj5Uzd/U3
uMNVuwA9jfmTekly37fMP1LiPLe3uTr8sSNGQai4aFRwNDxKzHbiP7JqdjL5e3SF
eATU233GMPN8JrZVtYKcmrlRDookSy1xOHPNxzqogs8aU0sFjhzRIym5D5qF+XmJ
aVlEVaXF30UbdIQYkybiiTBgk+06lz2stck2axyAC5vr548YxT06bxABIrhTgHCp
mlb/cfb02XjcRmUpgkDdsAspwbsbrfBEQTvB6FP0bVtou4R4tvyWIZopOU42OcfD
yrE5q2WwgGGdtoVpUUweRVGGRG58wKsJeDItoYVCBBVwPxm6pIuzZZ0gRozNQDkM
Moyknzd2s+rNVTPOYwEjMm00/UPEGVWy6hMAVNQhpQ4SqEP7dEGA5F557FJNTPe4
gMoaQ7hdYiG2ZoKRfzwcYPjVxwGCdWCvFoi/EXbE7YvWsv634m3X2ss3mtYW0jbE
mQgIkt0ctsZnLar0sTSdP7GPgDGZFJsJguYUExPs+qN2h3rAhKliA+/K77UuswHZ
vAg1MXVDh3utd8xMCgcpodRU6mMCh2KlZ6zRdrKuE1DrpMfaI2T1rIHifP4lTZDK
W57T+I8eCQ46N7sO5lm2KqL3WcqUiK38AYdh1mPqX3q7AZxfB/SqFXAIO38EFVph
/hDbTSKbulLb2/TbNFxBtDeBz+zQ6EhVO8WCjUYaBhfCwEh3vPCr5A6L40UeFbbm
laJur60u9h0uyeXxqviyJs8nO03z/il4DfQx8GZCcS/HbMxKSrluBwjuvHnQYsPH
0VhcFkLCmCJBCLg6IZMScyH4fPyjgopAJu4E2La/3pTbmf5CkhuWTEmVUTtpnsfh
RG7JXxSwMYZN1xM3WbK06NKU9lB1aOFT7I5T3IUI144BXllO0zZIpdIu+92IaPh5
smtp9+rfUswrwGGQV+8VR+IzEoyrhJ5odvZnRKuD8y9drMn18zj86HYmbVxJIf39
iWydbDVPYZEST/y2bKIcUiLXmVztg1SbCzvwI3JEEfURwpCT4/kKcH6o3Meo10sq
l9uSuXMMxuHSde3t4tn10SKGQeltr62K2iXSE6adHds5nJvMDn3rZOnVEE0MQBL/
5CjrpjD1UZf4qz7+CgNPddaDLr3a2PZrJp9Cjd7v5NKJeZoF1VloSpXSHOp3esI5
opmpnsqDicjNKmwzMoJWoEH5VHVC866g92GDCSCHheyQSduOKSeSAfZmLNZbW118
nmcoO18XkokHhKF9EIJfFG7LLWnqJTxKBbAqDBMROfUVW5XzotU+x4yFxNbHl6E8
pCIMiSutZddizLlQ1GuFiJmG79e5WmDzxL/j9kGD2sJvnepGMQQ1/ufdQ0dZ5DZB
b3Cs1qcooMG2ZLeoi1fzUbS7O6KFasMlnabJ1c1NS0838cnTB0jYiazyWMNDa/9G
R9N0AVkI0o17OhHbzO6HDS9UwBJnx6J6BO4OINvva0GgKShELWWLictWtVNtn1qS
GQYfgXQeK055yJHOeIOJTTB9a3ghwtoRPq7KN9bGq6W69rUPH+ZhrxMgyryCoIPh
TCXrs2cl3I6jy+F4jhjmqxXihBYMkRr5y2Va4W7gB7RQOY39MxRD2jW/IiZXODHT
L4tgHmUapm/IJnQKqYgDbJBka0joCnQ7aJg86/ouIymeQKTsQbeHauJsFNYqpzUH
QR5Bb/pGllxMsqJXjhlaU3UJHCUYUmY56PSIFfjqVU/dGRIn9ZgX7f3yr7ZbRiwV
SUu7K61/+IqajkRjnaHYJH6NZwS94pgBu1sEoxWc3GWdpzyi6cBJJHCEIPsYvhXS
qTNJ8g+kdfm/iiJsBInOI6kHD81GW8quqDnZLWZb9fizNIAe/1dqqbN2JXazXG1d
B43ThqvAKcvqQAZEwpc37nIvEc7cLhcxpI1i933PyR7Tf32VFHuevNWUboODAELd
6TxUuYjemhPexGSFyIPCIZ2qIpYZMMcGrMaw01MzJbmtsUS0N+XAosDf5tEZk30P
1u4U9+vyUBf81tI2hy616GguAMB+DCuocabVjFFSp0ACRfBr9LXcv3vriC34BjES
l44C3DUvNq3Iy3OI2aHk4MSVRf1ZjQELO8wDbg8kIu5RiItMM5yHuakm7z6IIFU2
f7ZLuhd9oEdfLlO1RYhnwNdH1rOxYmE3sSLkLe8kquuGau5BY35zRJmWE9yiY69X
TcB7TQ2c53y5udcBzG1gPFRmqHPHghWRqMBdvg3d8cfzehuwr+wYyyPpQXYPSfET
z7Pl/jsrtxQs2bmbh20kPFU7G3P0d8tuTK3zkZ8Zc80JtfCB9b2ym2YuoBbEP+4C
DKfWA4quxysAsZ37L2GA60QTG/tPkqKTTW1QWBlU6ODH//lzKzNbiqdBHqDixbqi
n3Bihk8AIRh4qlCBbJxWccwJfeSTudWjxA1MWVleM327bkVyuJRn2nKhSOwEh73K
D0gkqzUhND5iXcOf/Wi9yIwVAyu297D040xGIiz55eiirp0RbiMg/LK32kk7d5vo
pDkvsBdBBU4floNNkDdulHNa/2ThDTp0/KQ5h5tXqE3NsbaXvbk5D2f3EqQx6RiC
U3KIR/TAj88ok/jVNzmXvGoe0R13DQPAdjULTarbuEO6VVJW1ZEB1clvqvjrHCDv
cQnXhnsgccbA6UNr4AWuXeqRF2lMMWrCRmHWye7LukxIcr4Ysh8iIeVw7Fe3wGB1
+6pSSTvLoOqj4oJf8lOZa4eRixNMpkYXEoTPNJ8EKK6oE34gL+RkL1z2TE8ZUN8U
VYK0mXgfGvv/PTjXxoshIRiMivBARYnC2yTiHmpg9fEE/Ga2MURNccDiLrAE0Yiw
k9LdZMUd4MCRbjJtmB6q+X2pnMLXo7IOt0gONIARrQKEjHFk6FTY9jw0KNM3b++E
wzGHUk92N8XUKhfLVwO1OC5julva0p44f/z1up8F46oBb+vKn/72VzqyFdcnzetL
86RTwRqfoDnNAktSFXOm2YQmbz6Ni+lSep1Dnj7ukl0HR0VgY7kS45W8gIctNUWQ
zwDmJLxppeYq2tE3oQiGCHZ/WDHFv56qtzo3uDxaQVj7jjgq71+IfJvi8roI61HX
PDFc6TcrqLGu7gkuiNGKQ1pLOx0TcpHkNxhZV2EAgb/O11uxEXglX2LDnE8RPsId
d+OxhEP07mfX+N3ANak2a+XmOqMAuAT3/QCKOPsRERRTQkdH0RKK8hBaQA+h+HBk
3j6QF3xxfwWaSsJ8r1qNsPAtif02ag/ioHVpB6MwpkmQdUEoGa7PN4H8O+1zqfqM
P+Z156PtBEF4DyqTXdjmyNtRRBa49S8ZcDJXENa4wCeX98xNcHZKKdtoXb2Jcmas
Z8ZeKdEN3//sqeEdkP+WVb/9uWRn0NKlC3NApsnfxqIPt3Bq6vklUpHnuOIfRVtp
zSEQQw+nX5QD+eX78uJ5LaP5ZxHNmdwZ6PIR4UPDqLzLEUpyRWfdDzJFMmTuJ8E+
rXcliitw9rm1TcYHMs/YzXY2VrUR9gv/L8Rwi+YzRg8kn4Ci/iOq8+y6OG9o2afn
GhUHEQBkPLgHlgqWYwAZDhDUE8v/bw0F4g+BE+bi42lTbtvGzF/HWrfBZP3kJEDv
X+OSpnXdg9g9YEtub+F/6Dy1gmzknVOHerGvVLaw34MqQ/uvOwBd/+tPDZCP2nEA
hVDfl5HAeRc4muHJI/nugkSKkAPvHpQjbkAVMWitT+8GuAAOSL0qIA6i/P1Xd071
2aqw0WNO8z9lJslpJnM7b4rsHYENu3ohSU5HJjP7agQ/3npSj0naqu3hYKCCZLsY
fr3I7WzZbyga3dn7t/KgKn17aX86EFDCIN5RgFmJBl6RXJxHUT+i7mCEZH7o6WHJ
b0sU0l5EGBTVFXZ6GiZctKItmvbZIDH8Vz75yv2CnbT5joVhjCTfTHi/P7dUpJWV
Co+j9qkatPfSnoPQxh5lKO6IRcObswMo9zeVhKO5r7GKJ4vlMag2f4hYzpSFiUWb
q2h/4+wIwcPnhaKSkwlI8JVCh55wSGT0B0F4iFV1fE24R5oub5a+hvoJDWxotDoB
imIPY6dQkVLRQLmqQMo/DzTSf8Ct1bNad5n7l+cEoeUErjGrQy8QbPkRRWM/QLYA
L8NlxWInK3bJZSafrpwaER2x3FYMQb0Hvy8jn27mgfTfpu6bmDDZk0iPn6YD06da
Lh+F938Bf0SojqyPERWkNtMFC6SaLWLXonFvwJYGVmtuEEQsAAoeqj7u9jd2OixT
zGJdVl6PURZODuSfL6OMtFqrJueQRCXlYXzKT4x1FyxLyr137tGGA1kb9SXaH4Ya
S27U71kYLl20Nm3NSf8x3N+LBzDLUDvc+iQPKRcLsOmHzabfI6fn1ZkwxoJwT9eG
x+4XfVmYTm8sRN9thtOOsREehgAZ/yIXcylJ6mBBysMiZt4rmLS8f84kaSHYRVEa
pVwVsXrmKFt6sN0ZjMvRPUzykt5XgEIgwGzHG6J2qOxNn4pu7KbFpRUUPxigwO+h
njXxdH0BkYbnS7zxfoB+RoyjY/YrF/6Esi2siZUyChZ2/FyzG8Dj5VBZMSHOL5JA
VfFrE45NS95X8iAwb1yh4x8ffVO4Gi2Tddn5Ou39+5f9LIVidQF6avr07V+8W/Xr
gQ+uxpXXGYr7s8gXNU5Uj243D5CMLAMQR6JauTYEjKDVjKNHdj5hFL4xsuog/GQj
+44qleJKz3E2yoT0/3zQV07s/l89LQyc+b83Uey1wy5Jg5wJj3kHzrFUecDrQt9/
HpQI+/DUuRu7AUl8zKchSedurQlsK4Td+4VgQaH/z3/qr4qetxakeSjF+86trhxj
oetK1s3kUqeMDjB1JhSGFknRKyyOskDXjUp3J5dguEXgzH+xbD9gdlgv8DdoX2vT
9QIM/OHi3c7ZSm+TbSXm+bDro9lBFyCX5vlhKsCajtJBtf+MNwBgxHufYOVoqO+d
8pl6IMDgXqRWty3jYb6U8W2+6GHlNupyW/8wcwu1taJ71atk7DeopXR0x2JJ/BsA
Q7XVvAMzDfLpqQNOah78YRupk4E0Eln/mUnoUXb6zrigJ/m4tdvff2deSmuYAPaQ
K6WG5tfv7/KGe/vFGEyc0EUlbz1i6p3EMZNgU5zbAQzuiX9NBmCgpZCYAZBRymxE
e+pXFPwQAP4B6C6YYAdh6aA0Jzg8zp9bWPlovwPnG9nn96ecrXN8rezPTN/vFEjz
ZGVPXacBBisWNdSVxmi3LtzNq4UXn35h8dnNdbRvRPOX7bSlPPfWfTIWpdQbfzMy
UfJEVG83us3sOqQH9f/Nt0pr8+g8ktR+Eyj9Hzw38VzoB6mL0XUAcfN/E2xQV1TM
z1zgVl6xp27qCRdUVh9pqcltFYY/LQHl+Cr9+zCHPpWG7KCdLzjrHJ6kUwVWaq5r
WYArld9TOtvK1HT1mRQTg9NCCUfLMcqrWhkzjxhqGMNTS5H1j3IvwqCebc3sikmm
ivfCOzHsOPbFU/QAHmXI6k3gud+bTGdQ7iBEbb0zlgBEJRCmWej0toIm5j795FTU
FTajQZtF1KRAFj4+/z1WLXy2tE28M1Yola/g4UBhEu9+HLPvCXAf3xpz4tL1DSjK
4JorhFCWzpCxTb/JeKMpmh1AOL/HZnR72kmDIFXE+8VoklQI6dKs4FPjUnGzqDXv
LZ9JyUvm5sJi1Wa3n+bkaq7aAj7lR5z8gmbEuW62yAq5XhNGE05sxiBEGbcu1qU1
tFtQMWtFfoUhgS23a0iQ2yOuwwDJrJNRHbi8A96fZbqXtnbK7dW0kGEAwg5+hYhW
hlZcq0lvKTu9Ktyfd6zd2PSTuasiVVNZLKosN8UvW2dfd4Q1COUfrZiPyXMxWlH3
9I7txHDDyXCF/T8lQ5JBaUJkBMBU7CmKyGtu/cthFkcOb61EAnzo6Oy27MXCzhNv
c+c0Bjet1cZKUSGG8zk/kKmroSiPdiGthmQaolXHHP5rLItnzh2sZ5h/1yyAGUeW
qj9c2n2U6BgvDCXDlpOEVA8mz+sLcN3yILp+rN+8BUMP5GwW3GZAfqF/JTb9IARv
lOH6fMwV4My96Q8k6YvlWI2Ohl4MA0J7D3CZMTMx+4OT5L0st08ZsaPKjy2M2GMM
N6ZpLTT28I9UZj4vgcN5kSKYB40eT86yf74Zilh2BByrR2Hc39lft1D9KkChegvg
u1h8HVmO6A/ljri0e8tYexf9OYSlk1jpF0B116XKWS+RhG4i4XcSa+I8COCoXMZk
kz5XfW0ToL2XwWj+fMXoPoLUR+BkRBZkAU8FpF+RoMt8+7+h13iNG1lA9r1V3AC5
mjzFTkXJey4Tns47C5JtaAs3CAleOnFWR+WgmEpDdtVMxYm4/yPm7temErRBwLv3
leo5OpyMOUOdv2awLYngu3Lz4mGazeUBGY609fSN8VVQIQU/B3XtL4YoG55jNdus
NwDZOTeubl4Rb1Z29m9VuBxt5zI3XGFgGy/2/R/a+EL5yKbv+v619aYXAo9hUst+
Ue0A86Oc/6d5JFOwvizDhe7GkhTm3FmHow9sVrrVcIue68HM8XyTAZ9jNlLPh1lf
cMAqn8idSQryRhbwoSG1ND+/utU/WDimMsq5ta1zSQxmRaZol9D59frFcJ4Lr+Cn
QJY1wOvTRhKNgvXratXDycoFGev0NHKH3N5IGK2OdPMQg6+xpPttSjfKj7/Z/4aw
qoTVkxxP7yClwd+GL1609mHdOPbo0iQYQU/naViHmmqLa5nllxcHBdASkOHm7Wvv
13Ijdgrw5DJE5mMOUU4z9DFOcwIqSH1f+AEEBVbpERl1ve/MWz5Vyfpjkw/8FLP5
ZKwdA7U/r3pCjpbOEXcFJO/lywZRSwR9ln28V4pWMdb+JKqo7Jj/js2E2VUdPX/J
CGUkkRubmDkFopFk0/I0c6YZxiOkTTOVC2NjYsfudv5LagxEs6nucxgz4xaaA7ip
sKH3nXrggFK1lDOtjNm6Pp/DMLTgIkbJPb6bmXj/Iy+FHUHjI0cZ1fYf1JEOX9u4
F2aBLmkFtyoZBpcjNsT+LP+i0QYoGeMsFHUvn3qgkXDz49gTYk3+fr8HHaoXuayW
pfH4vmNvY+Tkmvb51n5a2b0liG+Odedd9chh8XhqHtHj0hi519Hsv25h/Wn41h7P
VsgtR2ZMLaL/+P4gsPC7oL8+0U9/5+KCJK/UJ2BHBWIpYPqoqJiRZ7s/E6LLhUv6
Ji0bkXZLP/2BGcT8yyTiiBCVwZQ+Baa7D8lR9on/8d1cbk57GTbvbrPuOcgzQwXM
zvRRc1IeUWY9BWGYcZCg+jFNAlTmrmzf8Kf/u63I4UVVosnGyAD06zVZhMuzeqfb
INAsnXZC/utv0NwjeIzFiugIG9uDOQfv1OVInvdjTYJril+cjtLPyYwaQkQ1FnzD
lb5wSf2XPRelQyg4hb4sMMic2tCZQDckKoZ7/9axjOZiobpxvEgJrczCPRvBVr7Q
sq32IMEqXs59sZTIimVFBrhd5iyG1tyTW1/vo/+n1eMT+jtw/O1yQSCuA5aYDEfk
I+od6GpUvhE939bB8T00tDA1Y7KxmEbDcTkxCUOEL3ydIcmt7JwZFiWCS4n660NV
xQxHNSQpl0FuC6IUhxHOrRswzL/+w+s5LBtmBhVroBMEyLx2rT+TW1KtXaTe4AB6
4gDZBzV9nrvg2sFrV7bvsqP9pX+1GEsFjHCtWA/MLKndTIAJEHYBZCPPdMs2e6gv
Iw7MtRSGsz/IrjEf3Eo4N8OCCMvLC+YWPF9iFLSBUkM9tJ2VQyIM1GGB36QD5hca
rTWx6Vv7LRBKHRkz/DbIl2TA4hICRM2HNmudnGdejqfIUGOLqaZS7flRV7Efx2xA
GplcVeMYh1MUm/ta6Rhg/d4BTsDbLVZuXdFlCluhZMeK0XhJVmID9tGc0Y0w/3xJ
ji9g+FhBAf0GH0Qf05ApHMrEXteirJFTbknUekQ7tEnsIZRLRRWseuCdHt8i2214
//FdqAFX4ANKokB3sc7lGfTHRj7l/fUxvDz6NUWva5DmrcnHHL3r1TXO2iLl5Tdu
MS+iaZMAiMRZ8jZ/GwVFv7k0wOERAM7YK1y7mSJh2SaBjg73aUbvFJK2w+v9Fj22
Y1S/bsxBN4caDk/0VUESWgeJWOwaXNyj0VgvXGwiQ3qE3C9HvW+jOmnHkOIi2Ebk
X70V5L9rr5wo9g0tb68iX8grwFlVCeRrm7YUmDbn7AKZ+swWzxfROTCHvij+a9wQ
FvOl/wXRdxbId9o9Nu59C9KbQ8Imihps77bbzvWZW3O27A6CJtmsN5xGEMBsBTw7
7sDvnoB4ivUp+gJ/+u/FYTI47KYLhSAAu0z3c7bxLb0W0AsuGM9wOufvbBrqTY66
pPnVSSIyw2p1mrgFXFWnOW2a6HdeYOt7J06JP/pgc44qXyShmYxSBGBYijfd0lV+
8IV6kkzbULdnK/V527IOEW0dnPOgBcEiwvcR8UT5ToVsWGs4gMPFI1ZTS5/a9x+J
rEPGtrCviOP+YCLMjZPCDm9O/8iGhRKZE/xpP+eAsZuathlLXnldJlcPb7KCyMvu
6sRzC9qOwt2vtI6VspsTEQDz1alS6qnxGWlhSVtRxO9CVA+2mPWpbRUSRx4f9aht
9F1FXXpdOJFZH548B27DV4ae4clRsjrJQ3LY5WyuPBmVzui0NAkBVO8bs8N2U2P6
+Zswa7QBL3HnZIf80AmKWozjQdAd8CM7/cfWRK5glXhV34Q/sWBxUsXfl8mckFJ2
pvBw1VHeT1zWyhb2zObhdXYsx7zIE+0Ek8ISCQin1MSjs7yYORcuZd2pRvDjW9DT
bUQHQrxlj2osvNxTt/dIho80gH/vcDlPfF039N/LlUlEm1rMwNuK2orEhvj0iOt/
wmtZrGSE39GfX9mKGIvNiiq8w9S1aYzdS6H6gCjIR68tJxbmKVUTUnheLYR0e6DV
xxVZ8QikGaTTBleiAd+ohnsMcjENNb7i+OtT7DrzqQo1WPne9shkB8ca44IH2bIv
Shw5JWDofWJ9Rpe1rizu3kCT1fzrOkdQgFsgjAyelFdgvqAjwSHiE8MDKG9fbJPm
RqIdDL8n66OtDbnsfubQn8UgBZXk6vEED7ST8yUeaWP/uxYMvfGrXhW/2ZB3dbHi
aX6/qNhOaGXITdKfc+fXl83AeJUvIGWgbQ8dyiznA8B60vE0/+5nEudnxLyw1Dbz
Ql+XyO79HKUGr4KZUeL++ETVP7m/tN/crZiN+WO4tTCc9tekjAN6OB/Ef1bahpTr
FdCaMweXuQ0vJB8/QDWLtRmxhKOwZx6f7kt76UCgVRQRldCT3WulYUxMVao0ntJA
1ar2boggOtEB2vYZ840DNELVuNTiONH0ECOZkTNG/c8njou++iJqUyFw5yjs0zMX
YvonQFbIweT/pRH/nOKxq+K+UVLERAJmhC33i0YD2nltgcQ5tUWDaeHv2FiBFEDq
llMQdNGzpt0ogZ58AnvAFDrfHUNnIfrBNqH+KinAjpKfuSIsoVQZni+0dtHqcjex
qGB7VQZZA0L6DPI23xeb10BYQ47lnoM7PG4LQ+bmw2+kCIgmxAMEnonfKxQyvGYJ
QZoMrpzp6mxR94iLWhZbhwZx7ki8mz0eYBT/kPPSSR1SRzv6vYFdVLepf8f0yVeo
RffuzeHJ027tDxe8TFSeaqrX7Xwzlk0wUUubt1tb8HKtPYakowrMfmrI2lzyTfH9
GcuR2uhxkEHT4EAT7NSvs3gJwxgNUA+UsjjFReS5URyDYz5iJS9EKMv/eQL/vEZ5
r+9cTwqSW8tCSZx9mdUJA5VXnrePFqsshz0U/Ok5b3dkNm9GoSeMp2fY9Fjj5gAc
HwbVdjZiw+MzCLGej7Yv53Efpx4GKeaxLrB0pJwsbP4Z7d0QQ1KfKkA5fpwnlSRe
jqTIKjXUiaoZlmd/8cDrv0qklM6el9Rr00m+lk9fF3IL8YPnywSRUFdXLP9w7IHU
myddrK7I+sYA89bZOnI/EIsGtybxjSQb5OMf0baykFuZ4ZkVqlztxaItICKMtASY
cQSreKUvRS5rOQ3p2AP4h/GjV0eji2vc4JGsYbbrQ0yHeA6yQUYRwam9lM4QRCNC
fdxgwaH6oGvsCvtmn8HOZUWGh1/oSxaX0GmLklAeS4HFrTsDfOaMTK6AE9R6Syy/
vwnIn9dbfn+z+gYeIL+C0CpfrnkOmH/5Okdcrsim5//FpkplkVXuTEstZ3oIIVws
xuD6xFHfIMoA3xUHCQzw6ClYG1wW/4vP+JzKglot4h7JMKV4PifKoZilrxRUCnnQ
GX25itgnUydA831m+pNiX2brLCe8BoJYPE5djK+h2ZgAHZxdaQ8ZAdGHg3XE8Lvq
ugsI190W7XRUXPGTMp+AHYRX9QzHxXQIOAQ8gnreAdmBQTJtyOhN6gqQVe0KoMoQ
qcK61sRNgepMAubzy59VeNH4d1D74qX1m8kbJFzNuvr4FDw2dJbR3Y51y1hg/x+A
6EdK0GzI9OMwqYzHhq5t9vsFCTrMOpyrIzuDk2dQZBruwSAzi8xxsThKrFIRYuKW
Jd2VQ9hRuGQzJrCa6LQdIt9k1/8EXC1zZILG6bqnzC5dMqHPh09ArUABOI4ZNkC6
4KrtD6t0SkidjvAFWufEhNwmQH40an6x3ovcrVkjRbU0e9+FR8ce0HzbolkvNsxj
luZ6VwujG+oXHQBEtQvasQach+sKeUk96FC5i3x3l8EIK2thC2e5Fe1uA2DeFSUq
0JrPsTtHtxHpi13SXEXgitE6ADl+iEVH6cHmIOMTPwfZdjEnH9VQ6byFYNnrShV/
Y0PivjrBfWYDj/5P4vl/D2YSGsewQeTOEMJilaC74Yh56ohfS5gpnVgb0uqLbbF5
u5ubTO1c5uvw1SOq0/hWsaxDaNTAboj7OxuaWfW8RTQPQaO5byIc+ApiLDY6knrc
t3oDhKvo8vW3sR7WOYbA1TWnKTSAwCCDH8u4FWgcnbmll+RUwOsClP3hQ7JoQ7WP
qopi5B+Mbm90Otg62MOdjOpcWCyLixqA5LcFcEgk1GQ6/PXDY2nu5JSxZokKH8JI
a7z1+kn1Jcz99KwFYMkGjbRTnnsmuSGUA5T4PBOQs46+DnknpW0cG7hYrr9mpJeJ
uZqs/NBneWHf7dBu8XGZdeY0gdJnoesf7Nnqws6hGwVi0igwD49WHSIbv8anr1dI
bKQXrNASfaDMiAI8RplKDpOic5DxweF/zpMs5q9Yi9z6h+2mSQHFU3Ay5B/W5Uv2
9Tdi+1BsjhpyeXcMxDoK4z+VBvzQvzGg/TyZ6faHamQw1IU7RkJDlKxKLeWy3cQe
HXoJrOevk7jUUhsA4JOuU6u1GzFLIPQ2YA7FerJLIB0NYlqVFxckj45GtiE6qdVd
Hief9t4nHRpifCfsNcpRPaWDbj0T95X+x/LtxYXOwETYrtZSR6c9sIMgsuyekuX1
dIVkGxywIwaG7ew/1jW5lEDrA+VclvUonx9TiIja40Giv0g1TC6b0mTzj0dvRHt1
vVaVIntVGDsmCxtu/F2TJGUzCD48tXbxjuI+t/JGfioVUjisvsd9fbip2u8m+cuv
z9svPLQjDHqUFZu3Grdstlsg8sB5kACARssfgNfr3vmcb3CC+YXPszXk6GuOJ8Pb
HwBeMEt+I5fnH9Ja42sDWAIFu8BEOV/4mFxg7U/uEGG8th3c2smtAB9U9Qfm1qSA
rVqTMAjaxcwhglrHwCwZex7JPYrzeJHlxhPYe+MRDxHwgIlOCyWxSezDHX8e0ifc
M2zlW0qVKh4t+q3ZmwZUVwTTh9GeUErJiI5Xq1wMxVc0GeTzMvfMGIgifD8EZoh1
1C7gWg2Cvmikn3EY9kJbiEHbxx3fJAv3DmCL5fvHihfAvGmJBSd39/So09bUpDhm
5ex+3sOLZfDGwZpiK29jDE49oSqB+55qhxLiCDQ1qUPj0JSTk0GiwI9iJsDy+wew
SR2Q/Vxk9HmeHno6Rkdp1KddXOVAUSqmGDOKKwPoAYuLe5c+KAOMXDCwsY1zlD6W
rDFHRJSKRHQjdzFIW2lmSM+2KIsmjuCZeVAWF44y9pjOz/v3TjjCvrtKMcL+/non
aSiMarvVV7COKxwgO7CIPDq9RBsMQMSd65DbAyM0bCmiUmCmIT+A2IyPAfcLjaPQ
lh4ioKVjYvtX6rb6HWGHSz4JKEzRjTUyIx6eOjV8+ZHez19thaWlkN5UNTih8GT7
45jCSUqCS1VpxcPHkZqNZXUs5PpiupEd/vFNLSR+DwEkx+6TdBFDDTTD3roFFmJT
Nw6VOZ8PzyrzI0nzn5S/Br6CYd1DXG4MzW/2+WuVlcUGSThREvAoFBlKbUGdm2Od
W1OE5g3Z556RW1lJmT+UnSAXwnwol4NGnv6QTo7s9CZe884w1d9YM7oEV01EbUsH
9Jpfq2wyp1hcNv5Bd/xGpNKvVHad6gECVi1wtockaAmneiTmG0h4RRq6ynyKImq1
5MBF14/j1GPnLymM3pnuwNGdXxgukZ5yVbL4J0gvg//QhvHVL/9gPipWTXPyfIkR
ZeC7peu91Ho7R7qHL0kNZ1/171vfIEhkddMxfp2OXA44lgrbjaIqQPczCUkuiJF2
bNpdRjmjwqjiZ9oy1pPf/orvXxTazmht3MlkQhpnBFhBFl44vcPdzI1g7MXFmEAo
nLRwzNZvE3U2cB+zsmVa5XWsQU24e8xW5wmsFX+qgkwk459KDWSgL7oLARVUh0ob
8NAcu71c3A12xmR6PJp+iuRmpHtTq3ECpZB/nb7M7WEMW4aJs4syEaDHx2ZrGEZe
nKJj8PLV5g2vOaKp2VY+Sa50BGzvhtMNM6h+Ztn3vpPR1mWCB+Maf+2t2VO5nkcO
Eku89DRozSaP8Ak9Y7H7TKuoiZ/L9hSr4s9hnEWs0mrPI+TufIGFMCv23Ijt2C9Q
QlutW5DLgGLIwKo0/DMllub4Ftbskzx9zUCw8ZdabpGbSSM71/8xOzIcVwImeym4
80l5oXFnivrhPqWGD/JyYdlrsDdhOJrrmy4tkfD8f7nRMxf59v1yXiw4eligpCpR
twEGCPVFbtZyBYLOzno6ffA1rkulQzAbYjyDvQBjYEhD1RJA7igMQRXrdRWwLKIo
O8biFBimgvln7ywaZh2786wF4pm9ddUqbFW4IGA77D8d94YNdAWfHleIHATxef5t
L2Jp65uP6/JxD9zeAKyNXqCt5w8aRVbgnQhu7Et6ImkeuWEdMHmw6en2LdivBXIE
/H1sNH8506WLAZh/i+QdTvxQIksHm6pjm4p54Kq9S0T8Ew3ab/PlBwqCoGgvl6uU
cl8VqUSnH/mlbv3x8KqG6CC3eXc+SU9z8BMcxx870C+XeEnLEsDCRHVJVCQJtAGc
IIN+68DTzscYQpLG8xisRJPxYqX70cVBzTBKR8+1WjWOwkn5e4jvE7SMbO2zd+1l
gFCAsL9FMEpO3F5yUbihblHK695nVc4ulchO9lmJWrp9zVkcAWF/+t9GYOXJfd4K
PNwjpCocAznKmCyRlnW7rsv/bvqsJtTSPSyVZFoXM1xKhVbt36f0lqNACPATVUVe
RokVWMlej2i+QZGuYSAm6h6zlG5Db3OJbHqLKJ8WXEOhPO5npobYliL1N9cL+g8H
ESwC1TXN/SeoGK5eyB0MVwZR6Uq8rd/4g8DEnEMEaHKr088mA65uVWpCCAvrneM7
OoE5syzHwPHbUV+oAflTzCN10xEwFj86eUDkVrHzcPwBuJO9xN3CZd2bCRFSTifd
WJCs2Ei8RH/ozHuORpveqMzFJK33RrO3kAFpmiFtn6JAP1GXyF5IAOSFBGnjZRki
M31QWA2iXqCFn7aRyeQFxYY31IQ270yNnTTVXkEGMfJnFu99nL4UpRQr76FjMv9o
wFMfsKf1DjarSFiUJCJsOMyHH59ouHM10q+exgDl0T25U7VjnmewJHlproGUgZbS
ufeIv/kDqT9n0d7UnGrrOysCdd8NYMqREjpvvALx9/C7MesPY0TkjWV3yM4aBKti
fAe2WlEHkrB81JQGx1luopYX+pqnBcdVvD/9u5lL7PF7ogAx2rvvpEvJZDkSGwW5
0HL6N508IGds0bTgjy0bZihl3DGDiJSPuDlk/Lm7oJivRpA25Uskj81JRJVZIZd5
a+bGs5YsickgUzn4+u5Kxq9nWDFHQ4mTd/LJUAQqtoeOK5cuASa0EOh7TjxIgXaM
AcTTXSdCqrhUfRsrsyUfiTVjn0ALX7JbMhKLXYcOsxCOOdO/vNRinQQcZtErSl07
AWEiNXT0ae0tRcQk/Z6Lxk2qz2YfXhWCjbaA9aXtpxIxsuxoKI7i/WIFJ/iXIsjs
6JEX21U0xUo9X59UtI4znMa/8plD0aE1lIDM8/Z40S3mroMf/qneLYC5AFHQbVtN
UQAndV7Yfz70GsWaQdqGNt6dpartPJLPAG9STaelRz7X18AkxoUMORStqZWIg2La
qnQ22xanjn/x1W2EpxZAth8U+yyziePrNDkXK5G6fYiN+nXQBjEIJyBGX6qApvvk
FFePDDyAVoqQ5HeEiKRDhx7D7VV/Ul7omxowXmjqKPR0GWwNJVZ6HkutUH+Dnkcv
6/aO++BGyI0vDy8P8o+uB6ia8FaOVSYql9k83ldkhk9arb76MhJ6TSz9oFyMdiVh
FtD5eVhxJZzlBTSnEiCXRLzQCTfDRYVvIASzNykxbityoMll7AdKZITpa6X3vPea
KkBaLp5/a/is2Zl1Ml37yXH4D8wzHV3LYiLmbWfRHUvu3BuNuIaQxmMZ6e+6ueuC
e4eMVplZE/bqMimTWCW2FkXg00egz9mGyQ3v9ZNTSjy2LKTVIdfVtC32IKE2fhyS
BTkWAimcQO+Tnf0OYZPb9SkbLI0KItyU6soq+M68sSsQ4ip24qkBbPeM0s5B0hOW
qWeP0lOFymW6pfyfiLpBBCVRWGb3OsqMB5g6hHGXqZHNEAgFidvIAl4ZRlRr3ofQ
KAI2ZNzm1Amtuz/6vjVTCXlxS6bMn1/Sw3vFmWsI0U4kYuD5bVyAiOzKbIKB6bz2
E9RMmgmqp+/0kzAg1sfWRQ2CdqyoVapVGZly4qTupT1dN4chvpi+IqBpLUxk71Xd
w1amLmjKdFzLUKtEVySXXqU5REt8TYCrWCXQ+ZE9uFq67Qm7kgwd7Oc41yXrcl14
uoap6+j6YscXGoDYzcSG0a/XPayYqoKRWA5YlZ46+pE+rzjgXsU0MpOm0lDIkoxd
jIM7mHBlhN7rlAx0Ax+cpFZPLOF/QNJaOHDbgJV7k/Ch01Q39GeFskGBIo7m5ndm
0dJ26eSL33OQfa2UicF71hbkwR+kYrgydodIy9DoAEmB64K8Q4VRij/XM4xpK2+R
mVMxrtn3CHDKzKbSlEcrXbHRSVwpUWrvDptjBAifrDTD7rOo46f1mr5JrFoeLda6
XaA59HnCcB/sgmDqw7zrV1aR0NCbfoUbS41LB9Ns8u094p0BiSJM6oyUZiSlHY4/
VI9lAG2UDI6LS1L0ygY6by3yQ569CLf8/I3l9CyA56BK1WjuUrTpjs2AILMc9k7d
P/Zv2KL3QN11bVeTRZSOO/GeMYpYy1zCg3QradqRR52VyMknmJqBPcl/kpIKKd15
x1MRGhpKbnJXcsYeAoNMk1vfJNER1P72kqt1z2O/cNv8kF2BCuCILS+O19k+3zY8
ec7Gdn+gguXayOzl9aU2tz6iHi4019ZSCSRruCWAC4cuZ15Yf92gD4gqix1Z+VhN
JGJ9vVuFek3zdKigxpkbhF/0kAPY1zJ0ojqNkNawfeo7rCktjaHn0SA8JTMxAY+U
BiRuOLmkZqLr4LRNspqsU/ous/Vb0asEkt2isYxkhsS2IL3dNM7GAk7jndWvRvQ2
v18LlB0bqQjfUMKhUosPWU0UGlGt9yM7vQeq2JCQStoHyxJAGoPfjjb2ZbipXWcw
nbb/vQxkYuw3xG2Hfen6u4VXi3vucEfw+3VeoOeZdkpjs6/jrS5T0tY3bcBcozRk
lCP6anMJ/5tnmknY+XoZ7SX9jlLfDsiw3dmdKW/bc+Kj55NcGqNHb9t+DCpPJrwu
IGEY+jPsZxzBPp0gv9TDxdrab/rT/9tdI1MRYp6xWUS4joAxYF9B26+EXFS6Rnwo
RK027cc04nuu9D6BijVXTsn0H3n+GH2WxuT6PY9AQje6j1VHYa2r+w2HOWXHOs0k
9i+FKa9sFcVCBH72t96KazTQoC3IJPiWzucLhlf67pwn9jLRCBOlBm1SFylYBK1P
UY7YNSjctMsXqRjaM4MzNNClzxz8at5h30k6+dN3MhfiWSyD3cH8kFx0wvWrMdPB
mGg38TYtGwYROMn/I5LQTbOm65LSftRG2P+lZeiEdo8SBIgB5dEAI1nIF0JrH07R
TjOMuAmvDF3czEoOupODAhkTI6z/hAFcpYW5CnVdFRWfHOzPnP8y6x2zBxzfGVFL
u9ysxx/L8ij/CPmOJNqjfp5IE5StPLwwyUnCzwkeXAKUbuvIdFXFDtEdMBs68iuq
Euk7ExsmpjGAxCC4UXyS8WJswafUW8MC/QfeJeOiTL0vFnvPMslEGjgCQMk1nCyW
6AXr6mmPy0T/Wel+1ealtpkrIaKQR9E+06aLpp2oLxNIq492zj2c872BMpkKlnaW
W06Qf+YuEu+FLNvLNoNNCwYmNGLFButKecgHrT7+bl2YdXd/zY5WWb0MLNRuFjEi
rRYod3qKatNof5lX3xHvdTr47Q/aoG3EBy52TjBwr/PKt177FA2dLbF3TFzhDeIW
xhz/qaEWzvbb7Y7DPnmb5M0e3Zu4MSxLXuL5FU49OVYSpAwCmDYUZetfUGR3/9nl
2xMKFSu/wJ5sC1pr366X1EdPdYpwN4EvVGMczV6DhWw06r97yynLgmMLg4GLfCnc
B2+JHDd85EfJrUQZYdwpPjGTDbQjOv7Taeuu5m5enrCMY1Ki2WRh3bEeViAncoAc
6A0NYUl46dtL4Zo6KhAq2e9dfHAe9aHtwJb0GMXZ8XmskzBSDSKvROQgPEMkocFf
WRPyNG/F44PDybm/BjPA3ezodgl7x82CqvTCaCSGcxZCgrWvojnNnz9Kp5EGLXY5
fbXMqNm98YHF4/lfgZmrHU+1ukXPTnT//Ai6g4JO7KwSB6/fis0H7gqwdxrE4C2n
zSrcVCMHt3NWcgcnXP249gTDuR/UyvvKPThsOFsjf3lbMz+soboIagyrbWYT7wsl
O87KmNFPYKpnn6YW2SNy7+5Dm3tpH5veire8FPtXewdClaw3W85FODs+3QvF7wDw
J8Oo5AV62sCCQ0xDKeCwdt9do7t8YMKzurr+Xlx6/I8Cza8B2i4tR4MX+pTqZAFS
buxGm3RUEc9OZj+1FwvtJsPiniZ+d47xirpmD7C/VPgn2OjgE72VkiS7WfIlkadY
pL2ywQui8npW+4MizcD69DqNU8/RjZD0zntucpjIkM9mLqhy6V1ArNjHrpEfJ/4A
SwBrq6n6wyFzfMrhKnuWXC2Nh0nGIFVeAszthxHUzJkgCx8g08Azmyu3cbbxg44q
oXHxL1ZjPcWsOwjnIL4jYEjUSfzgVXvOtQ1rWzH+D7qAF9TuK0GZ4uDNaNnKMoFV
oaPKGp4unxN2DAyLgkZ7kiDthbxg+ABiDCbwLprbg7hCwibfEUUL/ng69y5BZ5wT
CK6aDKrGe/C5McsPC6B8zeonZzfhyhqatB5KjiNbDcsxJ2V0HRMnmVfwimCCIn0e
H9IxYMT/5CB6+v4x2mMgHhkWZ8J+msU1c2dM1Eum8RCogN3AJNgc+jC8RlinDkjV
TA6m+ZH+Sfvkm2aUsRZ3ULZEMRVIdJRjmGge7O6FIxUzp2kgS45UZa3mmyxUupaU
aYbzLeHkRGkLuBPfociIFnrL8uD1yTYZ5mRLCHJs/8HOU12uUY/kgoo3qFRhlBp5
IeoSYBaeZEGNvKrfjdCESfCXtCtTJd4/Zz8qfbyugDTDMcXD/R5oobUoeu1NRmP1
keVxNN7ULshbJaWilvB01O3INbMipAAeG5tLcQh5lY0UMbbG07Ked4MfN8t2Cwtk
EYfGz0/ITtoD+XfmJ3ZAU2JCPmR/mCoP1ET/jLpWuUmTBSaG29cP+eUS/VSctSYX
mERNRfFgth2pa/SycDFC/cJuEDY7ZcL2h+m/8xpizBbMqzqKS1JJw69x0Dujk8JK
yFO+T3M7km1+DDpIfP2sPVH5PebqXvWUZ0dsBUzInZcKfv6IwNhKU477x6LfVsOd
dYDIrNphY7CFUFItcBq/TBV0shzYsCaphMzAko9GT7xJaQOkzjqKJeq+rmr1OUXk
fzStk9nj7LTj7/MMad+TPlTwP84ojdCwB5Nk8r4LtxnsAHIhFf/39aQQRlOvaUzM
XELM/5yktDm3eVXjzDPPg6F4943VoQhIPifrL5YvUM9QTNQur6LXwmWzJ7yyXINp
u7cjsKVuZKNKdDt8ypGlH1rr3LFlx91Ze5xHyEXCCT3ZZD0gmXM56KpwC26RjeBa
OHObEeqQVkwT7xkv5iXeCbi/fHccjdqA1AwQ6pUs0VXycF/rRM1wOOY+kcUuYdP1
A/8DhL6dobJSHTMqzGlJSzNBPrTJki9mq2x1TmwS4njkGuWxdT7J6VGVM80QtY1U
qRhIvFHrKLCjaWob4c0Ll45G6JmEe1wVNj1ohkGHuECR7rO17YI35sxH/cvrJOem
oe37Vp3lk0dOa/wuuBg1fsg10VLKusWn2mI4SNf1C+bE4FJ8ao4vNqtMnevT60YG
THtKXWQti/8xypaWwEttqpLTf3EVT5xC8cqRurQTjADm3xJasl7SE0PObpwkjp2Y
Sq7kXUC42/zxb/d8oT7JFsm5HWSwF+QCpDgkRknFQEK4XTu5yRIMJaRZJNgwQZOa
W/FfF1lYeQZQxUEQY4uFJc86YlfTmvH3k+orfOkBk0nPTgvaxfDVtYOi6rh5NQSI
5y0XuFCApNkxPYAEwJsRr74hIBL15ALOS4StOA/TkEbDpG+1ESLDNNcuA4ZzWpl0
QxliRrsxYgHNxb6i2AtjGOLb1CPuivjTrw03dqAAH6owLYoOqTIdrV7zZBRlF+0O
D0pOroYmyvWMJgNpdFuJ2eJBOK7xd/qO1WDHTuUaTFinhB5lmPd+MkkjcQgctrtF
BxfGrXmxQPvkMwYqQxLqGslcBf2wQ0FrFCmjEot91y8Ns0KMH4U6o/OplfQE3Xuh
rrgtUW3yOmhZ/f7NutOkWXWcZYc49Snm1j4wb6FBCpAXjf+YbcjNcP/OX1C3hk+S
t5cnhIcx6auggdJKvbjUYuWb700fyF90hNfsBt13OtGPmigXXpKKvbb+dgoHUsEX
DgDHygvmaZSWsGpZSXzlVR8E7D7jw33noNibkiv8AqeNYfO4YSlmk2/tFQLclMdc
kjih+DgY2xbkEC4/g/FYcUurpSmiF/6XAdVEI9CxkDuIVSJbIurfxkdcN7cmDIRW
JqhP398tKqL1R5E32O2PWDtge04JFgKJ7ZYV7jI8Jl/1dL14VC1pxtTMO9KcN6Ue
SWhOrOxVOgXX1QzvUe1m1lXcwi7nkxxajyCC1wtXUV3k2QqTYUwiz3eYGoO2X44R
Wx4/7d7W+8e9G2+1+LTCyoAlBlN6xrmZxfjuntzUsaLKs2Alyb0IDqmKMeydG/vu
7U6KpiXfWBeDoydeUUmW7AZEmyTf1QQ8YGNRalMjbRQfl8+z/+ZQCuM1UsrxzO4d
iCJg0/vLkeKT/CYn5DI9X/CBWgN/IQokBRhlAUPaex7h+CmHi8zIS46na4BtQzm2
LkR9YVb3djwOiciZftPvfuvVnU5168akeiYp6LmP7aIoWZHr71xk9uwGV3Nmv4AF
tDK5Yol/+MQneGG/8nVrmsg26KRTnKonAZaKT0LaM8hQ1UvFesiYr6tqMDGFQFjb
abYxXM0oPAg6SVWF6pgxdkYnfZPb8UFl+5fD2fLUu8C+WXqdiLBpxLOGMDRc9xMV
d62toiCmJyLRZdTBJ1lLwKd3qLIksSB15q2wlhoY/xRu2I7H/9Lugw4HfhhvGdSu
56FnCp+rF5o5ibeo4Y4AHYDCLHmX15q/WWipRQUYsmAKE1srC5v7tixCd4jsam96
ePKclK8avB6bErnGT7qbiAxAkrfnpOYbMnjy3Z7Ehcw4KMyMmT+0vU39RCH+V4tz
ZbdibHI6rwbKIH0RPnRgXUD/gD4qRbCB4/SnGbbSLO78FLI/CovR8PdunhwAg5V6
ueQoe9XEDuGo3doOBPRgodToLZsnhsc7DFLkruyZjF/ExX9jnONfyEIRXbehBsNK
PiiH5/BmLx8pFuazKnZZvJlTq06x5lVPnS8KvgiYNUTVmTr+7++3NHlVza6fv0gn
GhrZYHw51h4++jlHJb+EoajltEytXLQ3+q0yw/pE9pmQcdmXrRMd8xDzCk5vY1MC
dxlMWNgd5mlmbQHw7J/s6SKZECUokETcWohZ2srEdXjuQD2QRzDBFr/pZwfVMZV0
rj8QqZgT0ceyuaqhul/ziY7ukyu3dZaIMrddSYDb6tnC9qiLaD2qctRrEh3svYIE
ZaSBdQbkLluAfNwKup7uSI/hoylDkFL/FWoAHb15JOaX45odchZrx6Ge+PIqtIJs
1W26QeLtzeWUZR6KzB9Fbflx/GerxmljQN3pmzAJ6IEkssqHnAkRx0dOJu5ygxuz
mV5MS9knbxPpbKDs5tiBxdcT6v5OAsKDDoGGK1kqCswn+aeb3x1D/lRNmU1rpyZ2
LuaWj+vqpQC1Kv8sH+bXT5NwOQ5whUUBIkatLjyWoE0ehqACvDu3KzPOX4D4qQlY
QH3U2ZmuQepErNDRQh4zIFfmfHt+DbjotHSf+3mp1qrUYcIrAagQpwv0vZQOflY9
uriOAPAK5xBMwGZm8PkPo84kbb9vWq8k5vH/vHfgP5vouo9iqnUmTvTQ7+0h0Syd
KNUP2SgGStzfcBrK4J2wK1A1HmRrOaF0RiMHhmpdtX6r1GlWgr9T33My4jS9EoyS
iWKNzotKHaW6pQuSdjK3TquQtfzn7O7QFo71qNq0JLR5ZOnmFBCdxSTIeii3HUBb
3JZ91HQ+ylJhc6ZvFX6qHTCPyR6/9PSKVm8YHHsaP5xDoLHaGClDoVOt9ZNesp/B
55xzMKibeNHiiKOJqP8J/QA/yepy4QexvdJfQN1GFKTr9dTFDDCYqaxA0UsNKy2I
RjeFweOTFzbh0e/xepSZt+KFi7B7bLP9rM2rBZtuz9VHmkwV6AXwhTNHXMb7IzXJ
pqyiiI29vK7MuL92xh/vs8jIKnNfKDbELbswdPj4VGD0katdaZD1VNvp3DqJK6Dl
BYJ0XNRNmMn5nRbuEjLUeVggvuCi5FlWr2MyRjmzdozf7B5utLoB4Cid3U8zXasT
RwlAzeQmK0LuaN1UIlwQDvYSSZGAjxxQSuUcbMtLw8HzLWLI7IsfSa2jMSUI0OvY
nW/KwXyZlSR3cO+ffu8Y/Vb+ijKgliX31SAEJCm8Fz4dhbU36qbY6+Jy4vSvifze
f/WetVo8+gTlZMGDIHTTeUXEgjZyrgOYG+KChqU9aQVKBiVnLDOW4OZQbldoVPXx
Xc6j+7Gkdl08Gvoph9C7kpiVtiF9pHSHY2zSN0sRd2WvrZhp5zWhP2LaVwBrWXN0
50Qr+gsxHeZTaBi2FZQXEEcMSeZj75M+TKjDJUBRRiq7xcJfZlyLZrFrKTwkhFkd
+ghJAvrKxVz/IdaJtNCNDGPBa3mS+0ordZMP3kckGsK0q4FEU5ZdpQS3TGvGgV34
gU5T98e+R0DPGbG83k9MvoTwVWdfQELdI0zZ+sHNQ6XOUi9XXHN7QCJOc9rV7w2v
t5MsMOZyV+qebn7xsjvjOTUHvU85G1QpnBNXCPRbsGQEj4t3V+p0PEiIplEchCfV
lUuzHklnID9DVqXcRyCpkZ/+iKf48f2ppe3QcJ40K+AzwxiEtcDt04eLiSfobTsu
WZAX3sTYLAJ52RxXsH1BfAhymQIxVkgtNEuoQFooN4UFSRbb09hjwz7SHA/E6SRi
H+aTyBrWlfWpCFVrBq8gyYBg/M3LPAddNetLGsbLs4iy0e2DUcveTOxVsDQG+iaq
KMk46xmwivJ5bbyw5j965c9PAs1xhA0HAthBCmJeO3SX78woN8v3oyLLoO9dgo1a
T1aG3/j8M86b3swaj2DJVyywX1dGu2vlPsdMI++sbP/3qQc1oLkd9o/9Lq8NdmqQ
BFO95wE9IlDFstTvyXtsIvoHboQDEq5NPig66Thh5dL60BOxIf639ugxrw6mdW4X
RsHoyzxE7xR/cqGGfEpD+dI3rFpVQAL7CwTkWFa1GjPO5XMY2N/fHuJaxSqPhhyX
zk+DCUKNRP6dH7xWRKxzHq3oWerlZ+qm6HON8aDSRY8T4FIofykbJD2Fb51kNhEZ
BBsJTLReu/c6vfLLMsFuOAXTLrpZoylj73vXPqv8UgeGJJaoFZ9CMSzxKSijEK9E
tFFI7BfhxagzbeetE96FNgeZ/qf5Ih8mRO6tgv0szDu6sNFbkJVWEZRumwWHVS7N
d4ZwxACEbtVlzKVVDCQLosegCT4GW2uHQy1QTHy7NyFZJn57WDyxjj8GU57o5PDQ
0sluBDyBPi5xBRH4vI6SUz16VlrR5//fbZix4UQojIeBo78K5UKJFcjgMlQs0VWH
8JnPE7phtLHcqrrvH70F0+RihXlxxTAtxGEgv89B/7LjOd3shycsZ/gaCyQBcTXW
EGUDbDMie76o9EjMyUDRjnW6SZi9YA24GHHTyEfoDGh/c5ty4UdB0YlR3Vs/D5Hk
4Y46MHcrFIWFT4Cii7Hn49pC+WEWguIVB9gWQj7UbvqF16+mK2CkKy+NsbdzzFWE
30HTiM8N4XWu0cKg+OxXpnvg3KDjbgagb42brGpjIQ3suUL+cy0HJZHRjzOeyd8L
zOLP3ZTdaYzCqpJuWCp2Ur0GezN+uty7sgp//xePMGpQPN2i+qLbaiKDjXtCklUz
+e2GQa+OVuK9m5668Ofm4J4uaK7tBGBVkKvKbagujXjoIBf6MikFCPoT0Hvkr0kL
Ab/5tkoBPfbly6Xx8S22V3ehuVzIW44BFFQexssLHFTGWjhyh463WKwPeqU6oisK
7s+yQoxj2tnyxYjRPRPDzlFasQV1znl5Zeqmm68nrc4NgwEd5HuxhAXkCMqrYSEH
YmHfwOqdFM1u4tl8yR2MvXqWNzkVhNgOqq0P8Z/LpKIJmyBDxoUu8CuvqLXl0lvA
6hgS2pk7S5JjrbJPtGURvb9qTMLwSzjH5dYiSab6I5WbzHA/vXTVpiWphMXkQtfF
n7VtqCEJcXH/2MLIMY3tzrZ3dX7POXG83gCE083cZPNyWFiiBs5gWj+/3FuPoIRz
Ox72C/pSLlIo+6qAYuKJIqvdB1aOslgVX5P+QHvqiDfGSTekXpZboJubmudGFQ3G
IPGLj2aWwUlUtSeZSJrpwPOTQJuE85CyWKTnOsnzpRHRITl2S40CBexLcgdfe64Y
lGsn41TRLx40y0Nr1/Dj+wL9tkHcJkxn8hcuoiOMW6dhWOsG54o+azfSnMx5u9oo
rJviLzhstAjP5RK9UwpEmRought7D/ISp2qkwG0X6yqWTWrezTcJ26nNDRDaqvTl
0W6ZmeUdI4xWSRQylQnWu2D+7aOFk3ZptBFT7zWtJA1QXEcY8K19DCxzMFuSwjvH
dHsAlrKxgvSpeamGcuP574jzg+46UpeFI/Usq06XpzC2ps8S7MHu872+9H79LD6s
XhY0EexgmCM/rBxx/sYDL8N4hVO9j23GgKmxeSVCX0+9AJOBc1nwIuk5ejqluODI
Kd4sxhg89lLWybtnuCKEGLWtkqol+N+uvn5n/62HU2tu1+9qVi+ZuFV+wdCA9V00
a1RsI1Z43u0mCTqZcyYQTE8BkcA5iASUL0n1UBDauLyM5f6vL5esMrR9KPMkMfZI
vyEv1myMkFRnfEIq/RLgtm1VDH4ogHZlVJ0nicl4tk1tUpg+Xtf7I0EYh8Tyicxc
kEXq/QGniMhyRkemxb+voZpzkLWuULAr8Mk7Wan/Ykfn4mEdgANrFTrxBF7Uib8x
iI8XV1YMIeI6WQ9OExfPRKhpaXQh2skJSsqkeKMrsYD+PP1ZIEa0hA0xxvxXaiUZ
yWhAN97NLde38GYA75cuIHeZSWEuFEj8C2SRbxgsdyqSi7z2JcQUjS/BD2NMOefX
hMr595d0ENYQQmtt3kgQELnceEgCWJyIFbkhYk2BuuPEQyzmkgvn9YTLOYb93zPk
JsogLV5v0ZC9hjE4VTXq9MRZl1joLV3HKxuoFoItzBrFwIXp0472Nx26WdzgUhaM
2A6g11BS4LixptOvfkMghQRLazoI1eyoNdUG1Lm6wBbX32KMPFvxqfYSFKB+CTSk
uTveFJfXuP0WUnErpWnMdQBdF+X4TXAhi2qTl8FwI0UY8+lACozt2mAGJ0/UYr1J
bqxhZvHDBxEKxRfJ0BHZKXqITRdwRiNdJvXlvmmr4H9k5mwuev27nJt8dKf6Cioa
FQUjRiKi0/1KqB3dDE3IgrnyUCC+EpFQsM3Icym+0a9jEIUcdMmo1Qjjk1gRa7yv
1VlXSa09RqbnMSYcO+JC0PJ74F1W2wHqvxcHAh6ml+bwl05GqXI7d3yELSuFlr4j
WCda6aqtDZTQox+CmM0BGl3cdie3wDEZuZ3wNhBRgOEKobAmQuwVSL2zAV3cvlzH
0YOzvpu9Ox8c3y+jJcpfBhiwrdWcw9IgHikCWCTXUocq1XH4x1Gw6X3V4LK/wDFL
0MB4medD1WqgPFLPMEp/zHBPdXZvphATmw/3pl9eh6MM9BLaCBbSEXV8eK76zIrp
tzNVL0Cz/VyPyGiWsCHBtVPPHCwedwwGRKHJdeOBV2LC19jny4yryew47fBY4ym7
kIgwO88VWdsWSj3dPJ0Oc0zi0Fqivd7jfNmhpHOO2pPBkvD0YfM750A0coLMHggv
IiQrDhiGuciwmzr97SpstAsTuEuKxG4osmtrlvX4Ebn/acobt1Kxt55pLo/C5jxD
1i7AoMMhEijG/zXcsHkK1TI9uyURRQKr2sOOQBndsnNqFK8lvF8WNHD4QgiJmJTf
yBfxSlulfo6H0vRmQgjlfn25TCIvPHNnZLJtg/jUeYph5aZW7r+WL/X4zfd4a5yF
Hfd9iTqKcrPK59st2fsRQ9qiEtf/19XJNjBzt5k0TCr7jpnEUL9OzKDWsb4f6FTD
89C9Vdl8MiW2HQd1LzAis8CbirhhUNvnp0AUlhX6HSR1Vsa8LDP4cll+y6l967iU
IurTzKORCfcPb7C8rqeOeZ4nAlYLlTA2I6Kn9WNxB3FQGEXLEIg8oLbMmHkIWxV2
/JSKFFrY8qJdadOvcQj1t2S414G4/g1GHZZrJGMNAfJ3vuvqm3ZHHosZZKm4Asvy
H1piEVjH+TggfGd0caX3jsIZSDtPj9JQzrF+E/VbjZm8Zy0JEbijJhp18Q6NdiTb
LL5rFiq0+oX7tOyWYlKvLlEYBypmbZlezy27oqamvv/BcYVslYntKuIYWMVQX+HX
VXepd6qK9B8zdL2UfFhv/EEq7CfWdliXuiNsNFAtcPE6bxIRku2+HZxC+mR/V6xZ
0mykuYsc9OSoPN8lilDzdZXb/T6rQ83hRQNKgjLSmMN1uo5w6JRh2gVc1ul6qOwh
1OXsDzYG5YxrxJYJQ752zGGiA1E5ppEI0f1PylkWUsZGorMxTY9KU9u1xatdiQ+z
ZChfMS5yOo5aslNGWXdmYBDSrurzdax62l9jhZ2unVYRSZQ3rwFap5G2fs9ziwUT
W3AanCmG3LhI0Dd+crRhQXJJnDaBg/E9XVXhZha1Wn6T0CuOcQQHYUDWIlruFnM9
hYpFDbgzbWjMG9PiATJzL501RCEhBjJVjLTA+J5mg5P0aY2CpDjnt/FTCagaeodx
nMfdbGxq0xMt6/xPTVQ8ppQCjaRwL6IfyMqOP2hcpLwBVDdaLcfdKEze4/jXidoP
BUs3e54KF4ao6tdtrEATvtEK2uN/a494GfdQIutExQ74ogPu00CJup/jJyCRimn2
xcGmaP+12TNT6GcmdO3ETik0pbOqeWhVAK6jT/7Wx0h0Rqqv5QCDS4PWdaGg7YyF
Qq8Rux3gYhzUrlZNxr7+9rdZ0q3hvTVwbqYTToBFSl8pEY6fGXzERnqQ9FS8wOhA
Bl/eehAIj5OX+71rzgB02zhS1vj7Ye3hCqEol8xYdJtWeHU0DhT4fH4+SkykI1gj
4VwtV0xa9138uXwg1m4fvJcjaV28UUnEKYQbi48YA6S+d3qMvQtgvjKa3fDVJoSu
yOgbqU7gnnKUznbiwRqO7kDSpzZgSyD0QudljHIukg/PEsLVx97zgmzQ02bR4JCl
X0SWcrLell/Ll8GQdpXWfRGR4A91G/OWJKDL59RbZd+fCfVgU7Asz9QSZHSp5Z87
j8izxI4CvoKVy6eQIwxQub7RXGkyohf5OwvfM646K9O6D4cE1Vq9nKwEWZvKGsIc
HWBZgPy3rm7LTqcpnWqMaVR9zl/cumRtCfhlzqTm04cRWma8RWDyooNss84im1l7
XLVpL2gLeatWmPBTU9gNm7oyyYVMli9KmmUpy1b1oOjmYYtimnJkjxQ/JGD5iV0H
FXDKbLKsi0qjeK+g8hqm5wwRUUYa+SUyBcm16rhHAHnzIQV3y2YpIn9/CVRZaUKZ
KEKKT9vuWQ/rMTwi2BFtmwGIXZ6S4ryi71dbR3o0k7GprQtgSY7+jBYnsSWKT6og
Hpd28oxJ2DK59xSVATt3dnA+XkdgGHpF2gnotz5rcHXnGlwYeCfULI9PZGRerSJ3
5tAisy+6F/MbyKHrnu9EJ0k+uSvMcF8BhhXEvK2vPiJkjkxnIan6V1Q1ZfiBqGr1
9AidBVu2+eaLTzeaUYMexh31NYlIjMGRHyT5OFmKQSDdtRZC9/QqhEuxp6Why1ZQ
Q2PKBj23/RdQ1dJdHedcAdZtlHY8USvi2inXGGogGiJ+J1RRZu+Dto1AwCcbhkMe
v7dAMBP0PTdVXm/N2JQHXq2FktwQHWmAzXgFLbLVm1Yv3rgxer9Bd0tdCDh92etT
RdbqEsmHXz4IMsC0SJ+hS6Cr/7iS8hSwlp2uKZG9DWOnFcs8Iaffv8+pcz8er6aD
YVKuKSsYWrPtscrJwmoeyEBqoL0SGzyZ8ESu4d11d33thiSFE5RU27Kh25cTzXkB
d+L3hxDYvHFEyk8vAOqly/ffjasEhBULhAuxHRMCxMD0cK/VPUb6TOvY4zySZVaM
4lu6qML/qbbva3SC0Z6PHF9mwxNjpBmANf8efwbYl7Uqi0AvijSksIrJu31WbgkG
M6GzavPmn0u0tPqfhtI+qHFo0m1seqZXki3rSxy/mIFJ4w/xVD+zVXK1Oq9Hb+It
8qrLfI7uV+zledVrXzqYjiONoV6DSb1ZjeuOjq4PQ1Y8KtFwE82j/9U8NdQK6fb8
WnxVBBrRT5XWDc4+SCp1Ut+sxxR74DfAXjpCjXtTGZvUULgjqG4IJ2mjHkvChw80
jPiPrgog7Orua/mL2SnVYNsNbnIfgspltQu6r5wxLf7UXd1NeQQDjd+6Ocw+WHou
n73aIlS72/+xaaYUhc/FwMUtPU03GHTv1cr7jrSjZIR6OnU7frFQw2NjMStWYzy0
+mJpgdr09tSmn2YYktr4eNYox54KuSLb24ZK+oPSg1mcflbEvr/djKsnLoIjT7VR
U9wTGn+TbwTV7vsrvw3K1anaVf8NDhHVW6CsLJP2FDpCFw0mLbkaw4WI8RQuQUxi
wFSklCEut5QU61c54HySru5Z3aO94jmJmuNS8KFy6qN5KwfYhNXdrpc2FxdHWmG6
HAMYwHqC4GyrGdPSkqEsudd8RIc7EzuriyaQkTZGt7qyHB0MksLp6FaRqosBImzx
mRKcR501fBaxy7jUoWflyPCFiBGvdyVRltr6sqfU6/9ke7RGPtHa8bwk/fEn17Jf
CaNUaB34zw7KCkMqsLH87KFhQvWv3uQNs2kcY4gDr7zGT/PTT81aqzVfZCqjaY2x
zBy8aupwYFyOK8JbsXl7+KJB3vZA8z3H+A+BIgbm6ZtMrpHnv1h2po1WigX2Jzo2
aff1jWjpzRGLuWzh7TNs30N1MRWGdaeA4GUwomDeqUJ5BnLxghs4SOf6t4OnexPC
UguzCQYmagt+GFnIgcIv7QLmR5yeNFIAWzoo+kBBQ6ThaHoBUcuEMjP7HQzEpeEP
any5KIKeWVuH1v3L43pQn3tDIaPctAqbqrCKgwe/HterNVkci7S8D3exMi3IKQcG
drjvHqV0ktLX8VLmihmPvf7Trrv0cpqI8WN81rqKF1Fv5GKXpLmL1no6MEEB6muU
1bctDqUBTuQ5pu2yb1WhEFOAWrllJeytc0f7U17buuoXUYih9KgLSdMbH7TARceM
Gq9UX83gvke4XSXDmkpL1ZtQAefwvem1NcUwbTjViJfE4dIEM2QScnfV0036sqIn
eW+gMXy/bOFFONz+P5PIodMcU0dfdI1hqsxvoi6wYv5tORdR55Ow7IrspfAKm0zq
4PlQVtcCYWDwQcfmfxVW/8cVqPRFdRNJH4D+TDXg+WEOdiuCibTh0ul2wUkqk13n
W1KTL39DiZfG6SgHG1zTDnkat71fG9EEbu1lhctUh9cgDtws0qgw0EvYJiXAfrhB
IeYmVAjsjeUn1x/OZTttIMYDAPb9ZXEHP0VJpeXT6P43VobzBq2d+HQSmu8W6fpm
MEcCe77nxpiGMjywkT6/cdnobPZoIMdq38hdRWbbOFpi0qsJoY6YRO4aHi+MiUld
9JCX8evoMdJuY5NW+GRqXEe71I4yYCZBoDGMeMOVIXcij9z/s9gtPgMyKKn9e+de
+5MKsPo/WbDfAm711s5Thxc75t/jT9a7lVxhtunJH6kCmw5FiLWo5fRdfJaSxL51
zg76JkJj9cbIW9BK53zY28S28WBGYjelGFm/2ytDlj/4BlqWV34t+gy/cCGg/pG+
Xsb3woAStzCZVwYmr72bnwchrGDHF1stj0tEYMUmz6MGjPhSAG8LLvIIhkiS6qcG
9yYvdVWEwpJPgTwOsJab6Gb2nP1sIWl/sWJpNbBplIARsobZ479QQ2BmPb5jvdjo
XnoJgGSugb+adu72eq4/cdNqITNcKIhXKJVq90MCYDKb18KvwnghLVGyH6jOH8XD
EimOB+GVTiZmWO+yGm/0B+PKwggfoPFxeyh5OwiwCcEjUmUwZRlAUZRSlz6x0sve
5uv/mRkfd9qQemw8gq2bLSBOBvLx8mHAVOw3bPtkylzLV+aAq3L0+83BVZCVXXCa
wqWEscKJDwz6/pn+6TvQpx7CkJ2GrAqcQ6dIEb4/37p0/c0WPpiHU2js+ns5v8hI
ARLKBX5+oPrcKo+MgIS+wDVuqANSii7SzVnLZFk3TMNo7pILBmngvRG20IGHLpdD
2qwNPHz9x+Iv0ckGMeuOu8hSuFyf7psOdtOb0MqBWeqNhZN7htPOVNUJXv/xPNKJ
FWKwsDXbGwNEpJprK/WxPeahpwgH+BMALE7D8DlVPO1AK5YnYIQOj0bZQRolI5G6
S70dXNHr7n3n/HymIkjez0wY7xYNQvrNIRAG/fg4xC1YdLc2YleHd/yLNolyzer7
6Si5QebB44CWGFNFrvChT0Zk6+npXBQDG9EXM7irDSOuVYqyw82GgsVMA70wcOBe
ZW+Z3e0I1aBvEvytKh9nm/xvFu/jZM1En7NafZXwxVtZUQzUQnQ44sFlJNOvot9+
eoZ8MiNH7eoZibRGkbXyCReZSv3Obx/lKixC/tLZk+enfq59rXiL7QhImyn1tv5x
JRCgph6RvCki/LiA/x4eMLsHjVVjpub2ekEzB19MRlubo758CXyW8xN0Ed1s1jZk
shmpaZgziC4mveG9LOBAYwPADQNb2CZgB0PYlDO72FvmaFfaAU+j5WrHEPaDx4ay
rE3BuZg78Ow22DiX1iZ0pWR29gulBOpj2gAL2rZAA2D/iRiBT8ObuqqBavCrCEnk
Rl73hCzaxr/xtPdsUrFD+DjysMsoiY6RDzldeN6N2fFLkp3qOZu2O7RTxPs+eFdl
2p/Gt1GMeIBQLdRjTD8Ygkn/CKzeBCaMFaIcrhGqdRqa2ERyjXpu3N2GN5r3K5g2
o83BdVZ3M1JBKJzQ8ohGGKmxohCW5ybcgO2ST1Yv2bYJupPL2Nnf6nga3QHXbth2
PK1IV22u2YRlQ0gPXlvqt51Le8bkqIs//xZTDtToJDRsxFPfi8z4gmxwZ+BZ6POq
rrLWqIbQLIhX2h4l5o5vvuXId/wRpmqr10LiQPG43ID8v8u6ivRcKHMJCNeFRsGg
EBhciJctUboh67XgAbJZ0Zvf3YOoCltNANfEd4Sp6cQZGXd4menwwYT8huq6ho+2
C/K+Qv0vkbWp3jG5gRD77nq+TfDLSt7EiSMbwjFnDPXOdS91Ow6kFgYhsHfNZ8GZ
pX0O25l9ywYl/4CEzEM1mEAcRir9m2prhsmcxy5tRtwZCclhWqmokc8W7noyxI81
uyxh7JqDgMITQZOPp7kADB63KsflOtsmpnJ+2RfoQT8h3rEAJpvgxuEDgGEEQCIQ
4Jt1dLrYCpMk9WvBUZodJhvluSYTK3AAq4gs9I+qfE4k2NO9QUJhwfSoi1B4TkG2
+9o00DIT20LUzHhey+lM5bU2SF9h+c/uD6+NSjr58Ns2eOVMxjv/TsxWI5tbuDvY
HjnQJNbC/5EeznTrqTg+vi4bM+ujfkOs1xg8LSqYF3bl3ANTdZ5a6Mi19AGOUfIV
X+LJlBo7tQsLoAifF7K0DnbPinqCFU6Y/BsFwVeEci+wvkvckyeeE2x4JUXLw0Bt
GkSIfAFeuAgnjeqXVeZMwSrJYsbGHrDJO/G9tWMUR94LcmUXjbFOncyG54mjQ/lX
VQFSXtpm+0JbniIlpkf9P8+rY6JFh0DiqepE1zJjTUu7k8I0wiOqKP4obXknM7nY
jOCAXE9sG6N+b2WYB1Rir41z2F5JujqbGotmBICIVpGSXSB4mUz397EYqZzCKOWa
tmDDjP+8HPHjhnqhwdeRT1ZdRUXae8820zqBsvXd8cSep3A21Vnd8ox4WyIeivXU
/5IWn83bpC9ZChIXFH7JTAzfWys07xPMd9GwMqdUc6PyhdeQdu3B1stofVuE6rbW
J85jGtcj8mTpDP5QXFDiDSKUYfkJ/ZVR0s18cBA7g1eJ4KMpG1pkJBGyCTTXjjiT
wBEVZdFvKTjeGW5XJZu586Dqaj6iYG2I54ao0vAryu6dA8xk+sfm0dRyXStcOG6Z
ViDpt5NRI3KYC5Urr9TAV6HdAmPfKUGXEy9FS95xxTSFi6TgBT/upRe25wxxest1
cQOH7O2/3Vywex1hL4EhvwW3/pHwRTKA+XcpIcuDW8EtPUwjUl7z+0nnRCHDjtD6
4pGiU8lw2hhiUEseJ0eS+mGbG+oU4hDnaHjIMhKYB3kL3YrbfN2IWLinU9a+7+bG
vIon2ezK1bOZKD3rZa1eJM7xrOngIUO6+hVmZ3mo8TOzq77R+r5CXdI5wcKu4rD9
IArfCVIPjrgQ7daLv5NXSwyLTLHHO2DkDYQE1MoGdSMmAEsvgmw1gR4GvYYM8Fpf
PhjNrweNh4HL7whLo8lpdk3GT8TGoOeWuzehbVziaVsIGujqlu1sTGIvjnLWPAqm
CHTOnS96U8UK+Vym1K3jBl5x8oB7CscxZBhfERn4rBmJ7RUli9IPM3Hi9cl8+iQ1
6Vv+WFwTKsF+z3ThHlezxmHPJ1jfn892U5sCJCu0oI4hvyi1vYzDdo+ebC/xAYTv
FCf/XVRPpRmhjdsO/mZFwN+UhphP1taNKB9tKBL0ZYtjCHROTxUqoDsUFxQhrAdR
M16w+ZF8uAcwTSJKQab6XoaebJlDFVUpxcTtnks9flRjcHN+sABgcc6tqQYQ8ssr
cvxFoYJt1hVvYYK6AYbXoLCKQ/MH7ZJFNhLV0mDS500LB9bq3yExDZj0Gl4CRFT9
sKM5wBAnmPR69mUQNN83BmXdQ4MBtSBGbqGc+sRmIGWUcEtF2RSCZR0OQjmN0NNb
RCzu6/4P6uwUvz6wkvZjg45+b2EWg/0GXr7CFq5HU8zT06CrmGGagNrCySUvwwco
cMfUgiLm6fDGiBamwnO3FXRzJNXTPMuyvJ5u6oNo9XjLrD1igOeoyA8lbpW6j6xt
xcpcDh6kMdZBUP86XA9nAwyi6An7YgBOK3zdFKBmf4ALdby5UrNz3EKodr+XUdhE
r3r79GYjoqWmZ5KFsSwI1XcXEsaMV9EHVj2BHOrXpA/FI5L5gAtUajsCBJ6MfG59
2wJ/vzhsQboIbL3QVIR3xXo3sxd5/Lsi9Utk7i2VTdsdzAxg5V/J5ml8XkuDJFWc
VC8RFAYNKFbFF0yWyCorBTVVn/LsXD/NeL9szPkP7FEOXGExRQCrD5hznCyI7VS6
x5nC01XTLSxM/l+toAdY1A2f8xTJ6NwoeoR2kN0xQ0qCtWQTNngXAtolf6LmHJeR
iFSDtKkYaw2DMGBLBFEFl1GyOKVMlTng/kNBWWi6IROVnmLI4wYKUh/2dxp+QVqq
68W1gJO13CFzE3gKPY5izeAMf720GE+sTbYv/oCmCAGSoNY33wkDdOyW/gESaz8J
esqdnQ/Y0lUd2edST+caPVqjeuf2E0xY+fiNQQwxVtuyUVPYQPQVoWBYpStThXRl
N5AoWO1t7qIDP45PbbwKgBuLtd3pgVKFy4ngUQhm1a0o8x9hsw/an2TFoeKGIlmR
dlkhvAA9u6jG7+JKCXsKixe/HozferDEHNSPclBOGtPEGEqU6D84ElXDQ83cLe/l
C5iy1u/maZFVHshxX8Axf2u0SWudhoZ/p9TyoU4vklKGlA2xeAjvjsrSftce+FPB
yiN6vLOsNF/YDzuZpiDvzIbKzYpwwJzl1S8PwE/Jkw3JPn5aJlneDPWezD4tD99L
DBzBoqNVfLlnqvoavsvIrMTBsnOm+GDuC9EJhghFNQGSzgbR113IQ6JvJ0oCulT1
iqbKE/r7OfOJzWStW5cZMFoc3/+XMZSkWnG+9bDj3Pqfaaq7OWQHT4pG6ZVfP1c5
wHU+p9lj7YIeOUdZyDtw1QHNUnvQX2FzMFHomCuquPrjTB63S3HI4mRm1w/SWoO1
ccBtiD+9jTHfSungmNXi8qLLRQwzrX8mxL5W19xEuR1FKqAXb+KTW1RAqqeWM7FE
byFKnMpuIVMZ/DkKh90lYYDaStOQm2Hsi8t2/VAvGG7lV4YGltI6D72a+3GYOdoo
zMxp/U2bAlVHtCt+D6WqEz7JS+d+kvL9fgBa0zst74i4LsHHXxfzh+7bsIYr4Lyw
dP0GucDJPA3xiVEkx0Te4QEEp1eeK6/AaTC018AfHs9PyZWGqINzD5U0tKDo79jU
L6IRSdBBZFklOvzMLPzxr4LbE8Yx3odN0Vo+jvLzri+hoMc1KUWvJrOcPmC/2I/X
J6eGaUWhPEj/xeljwuUClLcUBjQB8TWCiAaL/l5HCMi3PrwXBGMYKSTYEKuPNfce
bHABgozBbMcy7chnsOtpe9VRWL4tTxdYmyIo9OPKgxBIacLHbWiJSem3KCJt6HSr
boq6kHzKPthmq9aZHDGnFzcB0k66Zoo40POezze53BA8qQSfZKUAI3WnFEVFq5V4
PoxMvzfRPJc/tnbtUJgL1cLRpvLLrhWCZHyFgqEj89NyGd9ZWs11lCbBEkNBwht6
RlwQBvdhOuDfSc+C+eA69wCCBO0+zmMe2szTRinKV6VH5j+8Ul5Bj5iI5KZ/is68
YZ+F7dawHfVomFnPrz5UHCBB7/rcC3T1ogNJJ/ixqD5alChwO99MHBsMjgj82chJ
X1vck4duJ+fRWgkGmqhynd5JqJObpdydJlY0jYXq2HC+AqarqM/o3v2R5X3hdoY1
BnLUKgSjo+57vk8wOnDsNse7Epu/IgHsG3Lq4mvuN1GPwzv/L7lPaGTF6A3NGPBP
9uosB851WW5xDazKQqPkAPKEQzvVbgJmmQErl7GhmOXth+2btaaYpptdI+vRjxqg
+5xzTAodA3tPMKaNEH/YHPuedDAi/S3LrbVIHaWoo3H5zBY0ZKXEpnUmfFN4xJ/f
r84hnmN2/lhJg4vgykB6cf/an4cTbAZLhcyNit7q+YoFQzF6LQxxI1tiJcJebJli
3KolZh7KepWqrOjLD9TBiqzjSjwFon1N0YF+yEvSmXTva/sizXzxFT+tA4KofFin
AqQYqBg41BbW5FtUMhRmBF746saM3/ifiNX7oqeHJRD7et+vhFEKCEryytI0hvs6
hdn8t5DGtSMgXigkXBfat9bRbC37jcUQQC3Y3zRH8i4D+6I3buIeK+vXfAAoN2Ou
5gC49K1omNr1laiQPlHuWw7JAWcG+sN+aOtEagTTuuuvqzRKIN/cH1RAWwJI6/Ms
UQq1pIwDbeq2PQOe5DSkE76mYD0e9/GmUe9J9hV4a6HxDMMBSRSzvhb1urSBhLjd
6KwCNDiP/pcvN5gx6IESWfDSMsGKHfnLKPb+pOxqJqiX5FUxNIqHy1oxwerkaEyU
11Q4E0DaztRQzJ3SeqgyguXflxp2JraFmHooMryMM31PO+5MhkUVmtpXM26vO3gv
7m46WDyLNMwyBIS0DH42aqHqCzN24E/3XtDeNGzM9fGBmGoUDBrfHyXYCre8t/Zi
vjWjCLcNjXqfHKFD/AQoJRcv0Sifa3q3blMgBLkwSvHBr0GRvFpPYUq8Rv64WkIM
WkuAxOAXwfr7l7ZWU+OpGQGEk9QGKLikJjWF5DwyNacEGYBzgaARJ90zyiBwYmKr
JXDCQQD+MbcK3r5NNWM1gGJqp0eFhBWyd5MKKo/6nO2Sms/szzL2jut6cDzzxS3y
Ihevgxg1wNGN6aM5nxDzBJe0jfj9ou4BbPK8+OybppbqTvbr98uk7MBfGeeBcdA8
Dn1hICM+WuqVdRE+JopFysB58/Oz3xhveqh9hlz8mezqSifGK5Tg7Oj9rdRsb89W
t0eLUDaK1202COBadqsV7a05C5onyv1R8z91J5b1y/stu5ssVpGZoYcwVB0zrV/l
RR9hFGHjlhUv0oB3pF0/JdZW4xzOVBveo/5UgUNUpBuj8tWXuhaiqvSMHHhZ2pNS
4DH/JsphINrufT2Ew3vH0hyJigkx1AY8crmzWjH4ixa6nATzjvnwC4NHn+sqH8w/
jv+QGkWfQcYMnIWoJDGbETpWDIH3pCCsCZSzx60oFZ9EC3eDSgS2rHTn3EA1aToj
eBElj6uTuNTA5FC/8kI8uinxZS+/MJbZu2zLMSuWMjf0QyIUDSRWVeM94UFq9ybR
Jm3lUn7m9NCLHF3jYyw3VJGoNLWjSci9NQt3DePEjA8t1cjt9wf5C5bN2g7ZeBZi
A5GPedjwQyCMHb25KB2Gjm2KGEkblHwiSWvkz79nuF2bm22hbo8EjnInuSJBgpBt
ypVYB2wHgUU/FcOsIuacwg4atXpMxo5SPCXkH6cU7WaIs/9lygT5jytCfho035Os
xifDwDJIQaZaAv7s4F1T6bLMMd2daMldzFvmJff4rPh+lY58VeTv5WVXxrSit/QF
u5UPEAPxNvtqHpI2FCoP5ofNWUvIJxVnvdDowL8J8epV1tMXEuMVRINx3wlr+wKk
iH68S3/orvq6pUqyspFCc45jnsF/1w0V7SzfMeeMIX++g2NcBAfdXPYuNAHKHC5u
odvFjvQlSu441wY4k5e3OL/CxuanHqBEoFaApN+QoEWoVsIFIDwxiYeLGnyLb8Pr
6wozrwtE+mmJU/NyUJmGd/b8Xue/7YIhbOe3IseXFpAKKefodvjVepxa4fLNnR9H
6CE1V9R/O/qiWnVVKcAW/cqwI0CEaLX5Do3dFW6eWn3pPfUZ1bY2uT+gLpNoecAl
eGKq4+Af/E5QI/Us+V/Iq4O7cWiLMbuBynOj0gw3db51nmxRvXszmZQNpitaaA6r
wZU17dm2CC7Rr/If0o5fXUDuvbO8qemzhzpYk7NOkD3U7qgUueIKQDlrrVl3SYGo
eh1tN5p1yhx71AAL/GV4pKDintR8/wXEOn64+L2sWfkvKxlVq0FY7z4xGbcwM8Rg
NTnU5y0OJZOc+OT9HOWKHLp1xWm3TNlkeBcr54ueFdwYObDYhuQvnV64z4ENANxm
tvI6G1yiXkkRmqkvF0SZKinSPXaHWuVOdOqKofBqqE4KwYAzLWzTvFigD8bDsGfJ
kmjS9jcEy96kvD0YjtO6NFMh6wF3giZo74fO+Il3Ov0zsDiHKwETKLg64bUUizdD
1/BA5wTcTtYSeKhb6nwkp65kX73r0hrZ3E5g9AJKZgAQfKOVGBdxkEoOw7A1B/8p
sLLWrbAKMEGpe70QbSK0uhGmp2jAKxmoyruVtUh7gorFN9Be/ln/0H7cJDMFXs4w
bDOnF9vmjmHH1dV1AaGci6cxRjW1LRkRv1xUgoFVfDN0DG//zaVjUQ9LvxsxGAdJ
ONMQ5qKBIwsq9AKcYKByvX0mG9Bdmhr2HmVqCfx45iMCfprPNaarpORuPtdLHL5W
yjE74WKDHRGZQswqeZ/f9eWk4VxKDdFhZCHRbjXZlKVmC5GxmfxLnW8ZMeEm9ngs
WDXASadynIffQqE5dau0j6Ps5XkzTMbNwbaWW803F/wM/8ys395l/6NLeFCpJO3U
8vA8Sgg5ws2r3O/Hjrudaho4ilXc8Ptkhf6wQDkJdUKnlT4GSVsNSyli9CwHFsAU
8sHhpa8glOE3AxvOR2OMIYrJ4tthY1p0fI7tS7wzYnGk1KWshbsXJeaotFSWtklz
nLH7WMrNojxFUrGHL8bVaMW9XVwcgN5R30nqkgzngFxQWGojyZA+zZjIayLfrp/z
UVrW5b2cgUrQyM85RQShewrHu9JMWUz0tWeSvq5a6k6f9X2jigIBKrEdio6dhzJS
/VkuZoOY7ysWUilHlQBNkPJ4vSZh0XaRM3KjzyLPEC/av8y5sjaM88wuvLYqJO0Y
KAYy5nKtON/p79vgvN73e+dci9VClEm3l7BnrmJQqBNT6/RpVyR5xSEE1+B5U2Hw
SSnKS/gEBC4pfQF0UGaQnbbKhR8BSA3mh4Gte6KWY7KMUzaCXAzuHo7YhczHVvIq
+pgmm6ZhWlcwWUUXvoeud35RD4CsGg39393n6xREFloFuLzkmcCiMM4Ia1dOEk1N
oUlBEOhOV1DwXdTDsALIIc8R0hlfxN/MrVfVHOUZ7aH8cRWnae890xxw9SVTDPcu
LIoSDgWPhng6PySbun+SGcPAkrlKL3G+npv1/M7X1ioE28CD7Wn0zuOTgaSlHJlt
iHdjuSGQU7rVvVljKBqXDjBg8ucbUrZHZvWATbnogZsEwKoHI4Qc+sLyeWiv5bl3
e2mwp9CevEH9Z6XsL/tW+zyzbwl2T+D7REf2EBMv6JHP4TsN6G/Tm/pcgqXeyZnX
KasJGUVvQMXhad0LNH2OAvGRXzwXmUBup+q9M0FGBTa0DbeSDh2f+jxEVogZwHUz
4xXd97Xle7xuXdTnHGTzwyConTPpJ6AeQDynvOomJ0SSNTVPy6fkU3YdPafzmtef
nEkoKCjKO4fyoCubLKfWjGuBaMT867N5D81GKEanxc7hs+r2mIu1wmGK/XP+4BTv
J7AqJOrm0XED3e5hXrfQJVlX5JCMRH6daiT0e/2JiXlLGcIHn9mIYtExiqetG66+
XSzWaiSX8NUpTtTkgi21CYdkEjInCeta7pjVSHAlgBeZ+x+6hvEY8zgbdjNpVQsr
vXbbFZhz1UcTW4+zpg/BSxgHE5oRM8bvU2NFnc6SehRj2Fq7+YNoaUXMqpcve6N6
9/xfnKsmnCJFjU0QBeZm9JBWllqIOLar3mJRQwrPdWkkGS/UvRhIfCYDbQRKEA/7
l4oZOZR++WgajgnI94zMZtGeVDYzTMzi3CUTlfPbLGDBeBhqmklvdCAejXmf7pB4
frUVkRR2Wr02IdyM3X2d782vjLJsBCfqYBl2MCQe61WyL82iUEpANlneQCdGMd+w
gIm7voo3EVgKqWb1S40jDzlpW1Yslhf9LQGB6xo0wfQkZny3i16L7RLj/8EdDruD
uo/waGBWZX290Sd/6Z1HuxkZ5nNisTe8hLMKe2qocuzHRTtfeZ+gpq1rzHsBEfpQ
Ov6DEr0/hCMYFT+YwkvCwYZ0/t9/uItcR7RPO7U7dmW0PEdQG3APaloha743VUVS
1E10yEyCdz2tvMrmHI7mzChaOy07V/vmFHJDn7N87VK0Vn16KtWRhS9kbNuO3juw
Uv5HEeh6/R9Iz3dTRh0o7JDSojIMSoFgKFPHmH3WDbWW/pAhEXzm3NM92hk4zowh
HCKBAsmGAnYFXPixnAOG6s4163ZjXqxuey3lP+SJRiszmN7NTAcJORy7vWBmqVWw
tFr1/aQXTfMR7DB3hm8zWGUdrBK1Msc5GCdt1J6E5UVYa9sYHHdrUmoV5PKLe0eB
U2uUBRVX6d0KI62/duwTeMRbG1lpsDkM0sXm8xq/ViYzC79ybBt6UEpxU/mZWcTg
2TS3/tl+f+iqtOE/2GW8aaP16dqzXe+vAym3+FRlVB5456qmjNC1XkVJUR0QtOva
ksDx7NnR7w/nqBBBa3DxngW1v3iBY4Icrb4yDUvIVs8r3ghqPrV6jUiOe7k1/gbc
/Q5nGCwo7JmYYiOXRKU+IAjWdwf5O7zHUkxcR0H3Yv+N5+yW5nWXOW57Y5fYe1i5
DYtA7altuR7ENHgHj1EZU1Sxh2sOntXaiC9TEJTopRarMbbnhuns7W1AqJDJn9QC
LYHGmba0QFs37mEPw8I0WqBHYDUSVE9VBivew/0BNrLGFYPM3MzQTyvj8mlbTBli
5Ucif+aSb8udxgnDBcepY9pTXyIG1wNywbpJJO6JuM5Lzh8+hFm6K4T0Te1tZz6/
g/+UwpX+FxVxxSkGTQuuF5pKC/iom/MLG64AYkOoMGeytuCPtnuI7GQgfpd5mXu1
HzVp5P+VcUtps8DhCHa9prZLN3CN75qoPuNWAEdIcV1aDR7v6emDNMBfsPNe16mg
8dVmAlfCYHtCm87U7uyndCxDXMz7StRDggJSFAQJp2kf6dxT2/t3jdLysxNKavh3
PemWutgky77suegKCJgeZXA1DhG55Srxsy8BC1SicMdYnDFc9OwDitS0Wwk5cWCp
HkavMG/XX9R0RKRrPZZtNSMSp2LBNfWW6ajicM2KoLdKA+FzdpOm0x8HCWXfMdOv
x1QEEGHGnXed5Yip+jt+9X0tN9PE/zCzqMqPWfMW1tmhcUEA0NuSyWIMdkD38I87
JSk4qEzUhcEUMTniqk07KpKROUK7ucGL43O2k7KG3Uo4iyYYhNH/GQ4BAc3LV9EM
PZ1UtVeifQXl8F7l3920QqeguwNmnTL2BP856w8WZwYOe3XH8pFDtIVO4T5+QY4Q
ykmMU/+kE8jgJY0Hoos+Xq0rA4QMlBgki8hDPkKmrPUEaRFD2VpvJr+iXjxouTXT
fXixxaiYqNERNc52liNsMwDMqx3e8SBGXCjBwjUwIFAvjP4LJ6h3IcXSIYkOuZTb
MCtGf2pjnO+oQQu9aKkOcQR+mCANIwQI6n3asvXhVti/K3pXryIjPE57BdlLJMz3
5J7NgJVLoXM1rYlq1r8gnJvgKD6dOLZPwUb/ndTsBnL0pHtQ8o4kk47yUo48AgFa
9wZRpY+Wr7Cjto5ZEg+TAcOMrJ0rk7yPptuZJiJa+aKA+aCxM2QftqNF3WlXyBig
BjMcygsAUM+hsuy/tUUF4skUJDV2QGdeQpcZc2RZg/+jb8lmuGbkKlIZTPbG91gx
GD8d/8OdCQtvywQQ4I7x2+JX44DEW+xwJI7fPV+u6OJshd+Xmtdmu0KIis6OGKlP
VgHahv0CNbM4O0rhq8rZr2ahT9POgmqQgNdSLJw010arxq1I9lMqZJ2ZO8IyWbsj
iYwaqtoOrQSB8rB2IqP38ugQ7MTchVF4PInUqhfP1WQjE5bGbujNMVDi1ahQ0DHl
L28ua3cLv+ORlP2OcWRoTQBvNSMLsmttd27vv0+8TcjK8UewceVQEHs1WXs8oTjZ
GVQZk/SiyHb+/lxN6YjEPrIrtOqmFmLRFmTOcOqHC9FAJ8VDPK/LpADTDxOUpxVw
c7wCtPrcEKvT33lCPgnNIAZOjV5tvAGTU6F+I2zvy85D5RLijDgtBoGgjuNZB5F4
OHvNwl5WH1/i5NrxyiRR/w8vB6EVAUqemAvYmCFB7yCPaXnyAOwxnrObWi+MHAUq
Ba2UalUlVPLBeZUfN1LQZzxdwFDOmLkbsiv7lDmWy9sKg2NXesyZmdCbc2nJCRT6
gz8sqAvNTzn8hy/Sail/aXjyYta8lYzdPiupUmIS4CuZPz0DqyHblumhx9UqyLGV
ZGtfcMssrYC/3a6VTkFZmNkf8oTbW9yNd/EZcJDw4mQLSLI9Es9y+Y6r5WQBF5QF
5TvZwR/1bM6a44m0fXyLp+TjvMmxqUOExvuy9pGz0j+TtkS/Rc2sl/ii2AEsvrfk
QqL7rhRe+A0v7gu69QlgbW0DMNl1OKXELwWyiqPFz0sUhdXLgPIJ9Dhvid3W7lFd
6x7NJ3DraQJ67147xuyyyL7v6j6YMIrF7z0KOcSlhOYGLQFuKfhHAJRSxlO5k7mU
bxUDMYLC2NJxo0r2Ut18vTe/5gG/YzVhEfEE6uTCFmJQ6VAWiBhuf6ULbcu2H7de
ZmDFSpEqZ5rCLv/dTzlRojjHg2i3DAlowx/qoOKP6GEpMwqLoiKs4+tv96L5XcdH
bxfCBsYlvYacLkOnHr70xP/EQZgUnJcwp9ANrhvYywxAqtQA06iZWfdVCW9vMPdF
ADL4eHZJNL1TRicUfvmIn2rdKubrVrjsaBTEoeIm0B9V2R84DeOEdaVyP16hG1gT
swLgYESGtG1U0S2Fk7KtsQyJ012hb3g7/IT50z6tC6keAtIZ+h7XaqB0A3zsbSeC
UTR4eK8xKRV4h3D0cQgx5RuwzlEk6YydQxPl14SHhi1NjaINPKa/rChoWczoSEal
e7rQqdOVg2EkjyNH52cX4X0HkWenwCEWV0TGLnJx2RMqBL0IrWBvY/t5352X/pqz
M7bvssJkKvagkWvbDMWrwHEPpoFoZItcTpVPVY2qdM40SllxJyxe2Z4zagZn2GsF
WALGoso69jxLjyS4qZhamM21kuA1Hyr0yueenf4z4BPhx0li+ZLIXokGrZgaEHbv
NP13mKVNm/fTsaJLBFwlK9CrJUfash0TeheJkohfcaK5bMN0fHhliT3orGdzuAuJ
jvugrfHxj5Ap//0jMm7Dm6Yfd5dgiKm1upkL67hk2748eOv0afuvw7YKWSHPzU7q
ePihSOOI08EoB3FUrATuzjXyMBS5XEzcSpPQYSCbq2HeE7FIlx1gXbOUn2FaF2/o
HRckiEoUTWSZv7LlWe8NMM6mxquCoSHPB4kV8pA+CZVsSo53d76ZC2D1KAnoRj8w
2syzz4GG2LnpnSrutHcj6TQZ7tXdXUe0C9jSA/9hF6kj7QHfa+2zBGe5DAi5wVUx
rUxfC65+KdWDv93yCK7zXwt5ak2scQS0RtYllmfiaYPJI1wuZN/nBJ5sX960xOQy
FwDtXf8wi4iF8PIGoT0VlgpELIO6sBGKzEv/yPLaVOC7XKLxT/Y871w0vCxWgdmo
oc+ie4dBZcoXq7ysgx4V1Wf+xdIJFrLFhYqxIXOvMF/Ic6PocN5XlunYgGqdDFBy
Oxrk827+vZcRg8albAr6PoX8OmbWnIWpwqIncX1bTliL/Yb84k7S91gl/jEpAAWt
kNGrZryrlGU/fiHxNxTruGMqOCc/y42q0QjNhfkeFx6oozCZscTpRcBK8WrQe/D2
kf33uOSzyK68hRHniVDxus0bvONmZhQTP35Wm9WN47KFV7zyFY9UWslY9tGBbhS+
cUZUGKlhveyXQy/R6uOEpWresMRBN+moqM1Xwxiat7KV4QpO+coXVpJck7gTVoD8
kM2m2QuKtXeuwMZTxV3+kR+U3XqCx5Grc5GwnqoSAcWMSDBhfnmEHbNB0YJy6QDS
QIvXpwlQ1napeFPuzg5puNV+VM6LYoPpDWBZQt5dMEWnocHhmBgq0H7mas/y36xO
PsBVw1tCXCbwLRrvaaVT/C8e1B3a08QuyN6Uu92S6gHlo6t+Kbxdr5jRJ2konneh
dUxrDcdZrOyWxNsWVD448PPxSxtYwXbxeL2Y7yAHeZCd6aeQibqGYZnGPAz2eN2G
FKUNGLZMHOt82X15xDnkCeZVrM1Qh9ur2GWyK+ZsGGRnNEC8jAyE1utT6J5dtQ6D
MqR6zIV0c/irNkg94cJZE7VMLmksaUutxEeFAtjcfwPmiVPor5TfPMUWXRCCWLzJ
634JeLMc5ylhufiClT4ikYvehiMyZRtUVvZy4JtQxsFC9FZuTeU2wt65qa6dRD03
M1GFZfFIqGQ5mT9PGbIr8dMrumaNC5dWhcjBDLiE55fD1ADQ5TcUsNZmIZb9Ew4v
zve/PHWEPmDyQ+y1ZkZTI+1BwADYBk9MlRYobUHnhfzvo33++yEMBh+viiElAOYV
K4t3fuKRn6m0tpGY0KDUdfrZZkgYeokN0xn0UfGe80tDxX2ycfSGzQcYHF8+8QHT
vGEjm5P01JfFk7LDHjKeNy3zKP1o6qE5Elq+qYRMxwhgduyo6kvS3xbhvJ0Q88XZ
QZAgfJADeepYW3Y7oWFHb1OXm6c/2tvkrpT14rIyCB8+r+YVMsI7N8hEjUhZVGsY
2LW840sjoG2jxO9gBh/ctZwDFqUObq0CNG8xzpF6lBXVixuxWKEFdSETqrOMARFI
vNANjkZKbv6EBC5uJFmaPy5vdrAltOoPr7dmUWbK/PaniX8mhnZCutj8v5oQr7D2
KO0FWVXc7CG/vpTWuHU2DGPG6fUd/hAH1rfbSSc2UtBifPEIaMP3iTPkcHU0y4lG
BAOgvtO7+GXYP0hMEXANFW0huTs/F1r9Hh7GM7dAlV9D7xmxETAFPuGhNtv8BtSq
WlNq2TgXqUqEfVwXMKF8bNhVLgn/QGpWrbvXGeobrndu9UUFhcncUQo5BONvZPA5
uKH4abXxfserqT413IFGiVohOtZB/pX5rTLCWkVQSXLWMMAU0iLanHRq4v4j/5kF
Voe3Jouj3tDOdLKBz+vhpYcP2dnQxTbV3500u6m3eAsGqdDDnlmjDSEXRikQttdy
fDtyTFwulBgRH6XmybrRY95O++1vl9U9aqW2D7jmC6Xk3o0DxN1vnliDqRu+K7UG
NZ8Rrb37pr0xwOk2qAhXYZ7NsYSYLewWeINN8no/uAxRPxvCvKXHnOH4dE0wBm3M
XQLYlQZOhed2ffLNPy7JwX4ppQF5blGGF2YdGyof3fuND+/p0QNHIzlEv7fs+LMw
IJinJUgqSQjFIEI7o1l2Bq0+1mXBeqr42hKijYdjm15tH5D86+is4XwTH1qiyY8+
t/M9LuuO8T4USRsHgoBuLz4JLQ8X481n/0KtFsV20/bCC9qrqCtQZ9dqfPOU6rnl
iNDvaEqeOVr9RaUMpbwIPKEg49zIVvOvN+JR1sESUdrhGpA5mN9+p92sHo/8zMKr
ApJJrWJBokr0WYh+bT/j/x1PMtaJdcwJFWXaLXFt+c/C2XH3mqLGj2BWKt07++ud
NaFAsPycbNaYDyqxTAySsNItJbxAqVAE+5WArShPerLEt3bp5uHrN9hz+DVCXok4
2erPkRC7ZrRZlaq487YEMBqG1ecvssr0qPULH45UPVQAtMErFLisrfPQTgvj8Gw8
6Pl3+8kQibEpIwqVOur9EHnggWnaKwUq5Q2Qis0Wk8+WMpWjdDsov0tCEayEO0fc
aHlxJGQjzNi9lW15LvvEDOjDWDcampc1rDGyJhLPRhPFVMeC4FFtpx2Cs2OH7sUu
98JoKedwTCmarMgnntSwAAKkCK0LIVnx94rBj7lVKyUMdn+MeX7MbIUnLTcohWGF
7acKmaG081ZaaviKCmiGUp78cZFe1sYZ26pG4wKaGu2ATBfTuwibdUmcHTz0Pj0q
WTTKgWJttHZIxzhgD+i+SuZ1jE4Lew8DvFV6e5t4wRAd9o8Ai0YGZeMOTWwte2AL
nUl3e/YspYDpmoSDw7zb3ucgvSnUq6PUInNVV3B23dfdD6Dp0fDSD61rr2ZT7MVA
n+fHO1K9qzka+V9oqTd+9ZX8HsIBMbbELbCTFsvhxkhfwjTL8RFExVZBTIU5PRDP
VHPMXAxvedgu52iQF+ccQgWBGOyUAG/GRggv5sgrfRyGr1m6iLapZd0eS2kwI4At
z5oCM1qZEKHCW2qJSFKZXr6hLcSswEKgZO9so+PPtRXsSm+zRzvhBb2byf4pxlxh
zGmB5lWh/d75RGZYNFkW1G6R+x0yHh8ZNvKKofoTTb0YKTXHS5s/sCV0zXMjwXn5
H2f8zc6ftW24WaSpoJONS/6oh+vpqCLm2DWzXGstVngOVFLUPipK+sLRroq4opQR
vdQyAdiVgXsu2A2XR9MsXonu/b8tnZiP/KExq4aj7Ek2BLu+ljm1r+Jrc/1NB3iI
2rZsE5OIvYCw99oSfazSbJjK1AKEGcJ5x00rtJd4gFYkKJc3mRdJOCKYhfmCHNON
XVvO8jGfh6mIv3Wt+xVuVi5CIy64r2qPqb+8tIRj+mvbMmTKENOmAnX/n9ZdCsh2
c2pHYb3N059AYd15rObR9bzyxVO7IktjZFUieyElLgw2Z3DmL6RbRqP70Jh+HvGN
OHK8VSXDhFH6xxxkJdpbA1ERM7nUFujTpdOzV/FIW4y/vJWP1osGsmZSM1ZtdQq8
1Db9gy9ucw847QrZ8sakbSFAEwauXD8u2kBDKzV/IDBO71b9JSj/IoDlsRpF+2ED
vYTyiwTXsdXzNmYngYP1tE5iJ2ikA/6zdlhqjCJrzZV6J5OKpGyGn5t4JNig2EUB
MBUxEgDG/TVJ5JkMZQbAQf1XGpZkEu0IPb68IHd5wIOR4Qn2VmT61keXEr8HZAS7
feePbusBwS6OxmH9iOTajilFCi2w5HgKcP0P3PkrRfIkmnPMiJKtvLffbstqtgli
toCoECo79a5f16wtBx7SonUxLi91LMHpezJeJeSSvbg7HOnDvnrcdLZQqoBXEl1R
bAO9iIFksBF9vd+/X7J0JzD0LJSNUgOcJnT0WLO0nvNn4LdZsRpGuwPTm4Us2J9g
KK4wBGhGI2LDHJqXp+Pv6rLywDR6QmTFFSd3SDGa34jwK8tIxxR/iV4QZMZe/Q7l
Wuo7HbTslUKz3iABY0QjihQdikfzsckafyHgtZSfj55UoudHJHNwI49VXdhWFn0p
o0XbmVF1HmGtgfByNH/2pS3VIHFu/dX9/Gqscx9peqK5yZytYPww2lqlbrsIUHGo
0LqrJZ65uMVFBnR7D5oZL8WX9QNIlAgvGiJvz7nGd1a4m3rytIAumV9pbBXJsYah
Celniz7fmx8AR3DlNJAg7yt74kP+8UsFQNXTo11TB5MpSWvivmjpZ5kIuLkWGvZv
YxvhpeJjK05YR1tXA7a8mBYWrODIyO8Pe+lE3FBBh3id06viZY6ftXVjrgYETi+o
Ee33p8IsJmV5lhyvOoaV8DuERtVmmDvBoP9skawkSkJmkJuXHfxLFnIF8DfJfLxN
RyaYH8dzprqZIp4hYCMQsPpB9OeFdQTGpVX2GpiBEPXM1Fk8ewmvr1aK7YDtkpTv
CizVG0tmI8RRaqRGNn3bjODq+zehGXZNjRaLBwoydlZWnYoW7P8h1WtFbL7lNvK2
LO9Z66YCyj5qvpmYyT6U1ZcDCU9CbQTx5AEyRsZNsI/r39hE6L2UUoZykecKJDA7
mOKE8RKupSn0elczPAvAL0txYloMU0+d5OUsknQooLEMxIaOOsARAOGqInRYrGU8
hnGpYiEvY4kPZeAv0DFrqlLsX/+qOZ/U3dSau8J+9djfYwhZz6S2DdL66DaP5wS+
wzq4DIo/3nkKfkTExdiXZvOeLy7KXmEU5Eih7I7xAKwosBSiLD4GOUOrf5W615qC
TjH64d2FgV+41o2qrkovqlGYSOUG+YI1KzKaQ1RHtOyvB63QCAGf7POhch00Mf0W
ZSjQI8mFXxMqahdYSNZIieqcQgfKbYe0K4ik9vSglt9yr5JHXmHVPMsMVZa9djw5
kxWaFhwJS2sS2EJz7k0HC7EYzTnGfF9CIf4Apz4DvlAdixfybg8LqH2TxU69rJcr
aP8np0g746Sfo2EuxbmLKJk9DJ/J2iy/gI+e6eelyVlmABruUgSlvmF/XRmQ+d9s
7O06gsIB09mqFUFkL5WohfC7hIY6/nqxJh5fqnrdjzuWf4aoS9iTDxGvU1MivhQ8
KJwBfNcdX53UZOwduyPozcdT/wciVKLUCGlfmA440Vh1IV4+A99dXUupgc+ZeaUN
eJJRLY9cdyRb1I+l4VLSigpKOLDjstxXOzNPhbHSAF9R/Jswv4a9J3cGkcvErCSN
3S0SglHQTdFNpFiP7umUaQVTVGmDzNnBB1uUhFPesySLOt8Dl+nyn0XZNiPvw+jj
JYKZ6gYmnvTAoiGmQM2lmaPjcUH0pvqyNam0HzNk+Y3BmiNtfl+JvWhlUKkoj5OI
mztiHf/96O+/fPygRQy5tpg27JssHmKW5rJJhT4+ZQgHgD/rppAqRzv5QK6Yhb3v
WKoVtlj6L3wiL4jS2M+kTFCh/u5IWl6ayAHYQM/Djk7YVGfEFj6D/YvR9h6jVYyB
Wlox+3AOM8ccGx9OBlo7RF+hXeFhujpEc3azgRpYVzyjiVgXQWu5eAtunZB9HmFV
UwvMArbqdUhYHPYx9vus/U1UialVqV4RY/sKUvfFm+L274fJWpzWvxU3DZMk7cxT
E0GDo608SLOsPOBn/vP29yF1/gRXbZnHjb4D88+Tbs3eMDMeQAM4OXOWyTb0+43e
C6EJuOvsrI5IvDvlONx31v4zreVb7MlXrny7f6i8H1KNtjyNG8Y03Zvsb1b9Z9cd
sXUQQ5f2nQdsz5E480XAiII4exyKVRecaEZc3ERZAjqeEPx8oPA0ZHT0YMmsl24O
7iJftJZtwrfsaOXXaZGWlK4aY3uK/7sFAR/9p16jMO/0blll4vJ7VEFBU557+0Qc
xFxR0vZoDOBP0DJzFtwZ0mMk1XoW2Qmg+90l4MsbCH0QWZD595lmyOaCzu6vmeEe
4tUGr4+nm04eJlYqN4PGuzvOEyHRKaXlVBLHmRLRk7M5KNeXm/F6vFoQPvw9/kYh
luOErLdDBN/S/k+tprAaLipeIF4H4H6+GB/RqhVsjipQ+hB8Gn85rEWyiCOip42v
viQ3JpfEbNKBzwIbhtvdGMqrNBDNl1h5Y6FQ/Mp4R0wJvj3GfQEmnqzbPLeb3nbE
U37Tey5W81ZehEClu/d41MzPpR6ijEzFrRtrK5OgZjPevhsihYyKrCsyiEmuKLYS
b0ieGhu1f42A9rFTAIo+aJ+hWAe3ox4+4MunrQqCM46UwJ8hvFJsBF9rhsUAeroS
jErDLL6tOq7LTnGRJdZhfYS7fuzSqAppX+LqsaUELpLMcQyc7G4p+nV7jwdIR7S/
l0s6NG4Voe8DwqgCr+kqM2GKCwoTcdY6Y2zXnN0t05P8JDjnizadYQZ7trMvMDHQ
YbPjfJGWntc3cPrOQlWrHpnnE7+Q7rOhQ07vHc70qjNASFrkzMMKxa0Oajc38Gxi
aODWe2CVuyrejjx55ZdpNdspC9LuUQG/ZfvEIj7MyRzuBX3YDE5AeQ82PUZca8g3
OZc1RDLpIgoSlWQ64aGBJ34SQ1Pqtj9WNJnojKNPymzlKI00WfovYjGw2NpuhnOl
i+LycUBhr42N3ykgbkhybzMzbgirLxP5l7UcSKJWi16OIp7wM1eyg3nt/W6W1IdH
aeIU0u1FuxfNl/sDP0TVKyQz+jB7JpQ8kDfrQHlnpyfTWJAdCqi0X12Csular7M+
NRJ1MaBLEGjwDKNECy+NVoGaB5llcMbHzxm5GQmEGTZnWKx1CSpaPlJb5orwosOo
ZmjcEuHfyKlykJOAeRsLTvnhmsLfsw9uBhgibdmM+YRzCMOajaccrktZYNvf0cGH
h9K2CtS90mgXYZloX+ILwq437bCTeBbCELM77iYi5Oumhuza3gnt4u3fl6fzxqjm
nRJKdoYzkF4PBJn1eQwa2RcYE/O8NJJoeGyYDjig48eVxQ6EQAubQPQ1DYRIymDh
k6Tg2/nrQv9nWgjuYH/YrHkz8iVbrnbpowhClFPHyM+bylJGmeBpkRLsQ3ynvSDx
H/e5ZmM+GGyhPKzqrdQZFuSNgtnT3cs0mN7HcapX9cmBzupGbjLolmQD1o/MezA2
PlJcnKUihWJWb6KAiWHVmYuipJlyfdjmoCXoXvHKKvM1Novd+hXlFxtgeI2iJwzB
IGKncV/IcoPw448i5iwqkH4GNyxDfvu8woxxo7+isHp3y1KqE2rVwKLqJR9+vLmP
oGUnCyAE5dh6uMGocOHQIrU7W3PvKA7Wj4eioYrdohbfG13GIEMn2nsLVoTc30R4
74LiO+N24efInB70rA6XAtMLJPUU8bfrymsJ3gyKCztS7B20EJYqEp5XY1iqlhWQ
AiTSlL9ZGoLj70OxvL7+ph4g2Ki768dVtLVMy3shSR7sgx0l5Md85BbilKS6ff4k
EBOr12008foNfbprbv/g1Q7eI7nhaKQP1zI1blHytgl8XPMFK3XX2WdWmTDq+Xq1
DdiZIcVVydNNBO+Z/sS1cIWfNuTzkSRJNFp1uuv3Bzt5H1IqKxjPEECWHBBhTuPO
W0yYkt81nB41sf5z9d/qfjzbYjZ3JJaUWZm1JDJGBQTQDxprWmCcPAZJR0TsLf+6
MsRMJWZD7OZ+EP9VmCbyfadXVQ2zo3FzDsPpFw4tZV/RFn9w2ZtoxNg8KsAuO1Ja
DyNJGbcxYSyWkBXzzgJyYcoyeUnrBsRshU5cXoR37nyRfzAX8ZOsCQIAYgm21EX0
QW+zna5nly+do0ulQ+F36+5vDZ84Uh/zLWWyLSb39fclpUSgK+dhAocG7kVCsS/j
C1YVcD9w4CML4sCJqJww0Ee5e/iQmD6scbw8Q/2j8bdFewZzeBRNp5M9zxuDpAv8
GI9M+gcy1ASRGgIdT1VVZpm801vENAEGPaogJGEsMDg7D3SC5jiID51HwId+sPKO
VCnsb2OEt9pa2moA+izQWR907kp3eK8fXuz3XB+t69/rLTqo8s8yNOkbq4ml3EWQ
MstJ+I0BQ/xtmg64rq2j6L0f/ztCKEdTZdntOAxwMNcHLeub7v7T42LAq4F5TQgf
FceYB9Jp9IOrR7e0RJ5kwoN/CPh58oEL/fd5pNRIk9HhOfgVilKd9pTKe2VFf21C
ICP7Tt583QStS8NkVR7NEeqUlkey+1Ww1DNh1YXhvyOEP3PJsxFCYDyj/AjFBJbL
as8B9V7jW8xTSNSSTS8zq88CDl1AEfrANmpDvxhBttQ6GwwZibXcvAD1aKFB+jMo
XmcM3lwH1yZYvbEAFsJqRNbrJktnLapHrq9oGVJRItYQHnVx3xmoktpt/+Mch9UP
JykY+oIYVwgeP11uWbJT7m7Uhsm+nI7YLBpi+I93zhepIAnUNwDNULw1PdGKMse7
3+SuAUvhoKukJUIpmOFIlAB8G0zn6Fq0nsi5ycDSincCLJuK6EN8YziptP6+nnbt
`protect END_PROTECTED
