`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ux8mnrneyQH8vgewgxQ4bUFBXjAWBKRVYmoxoZK6UvIhDnjwLnh+wn1BdJn+C8QR
fdgFHKiVXK4F/VeSIaMJcDBBQwn6QYp64hIysCR55RDKhD2do87VAq8UK/cYGbnG
Osiuymd2tKQOlOqwPW4sCt/omwob1DpCWbvUj6INvZxCc7WUSztVB+fLNIGxXw7T
Kw/6DroPyINXpLAK9j+livf8IxbJ3MQcSCz4TI9VuoN/jgyGpXnMsZ32oZqr/f8q
uK5uTXvg4iyw6rRfLiZrNmyybuafhFz164BZfLD5WDGDl1gCukbV5CUfOQFilNvY
NLyqfc+Z2hK1hWaalGk0PLzZzW0HR7SsfmWJF8bPtbDB+cr89aVRaNbk4balxnyr
WKwMKTCgLidECSvPQGOlVIx7Qu+0Bu+TVbH2GSP+EpUrDbCHhyMXzWfWAht7u63b
1vW3sbT3mFzUKP43meev5uBQM+ayAhgn8QTmY+titKo662RYRmz1C0nv8XfBEz5r
uU2gTUn8EaRMii7Z+vUAhM0Hdq6doChLBmbQoHJwd0OrTCwJW4dReY2ktv2RQqoZ
gDbvzJ12GmD3Leh18JN/VvT8qr1zftksgDSToAGXN70nrnU0sJb4ykn7CDH6AIrU
+i3msfy5rDThhCh1MrIfn0whT+5D74TGe1QcGA70cGICx02PbMu5Wk9ZPwUsaIYs
YfXjNZOQRrGa4ZaNwRXA9HWY14DjXgrN7g4v5jHkxU708lWNzn4mgpZIkTfr0tKx
Ex/B77GarLvjLvO7NfEPz05LiXDwRCjvjiQGo8TEU9zRmDbMtnhoUvbsTf5m5cfH
uYH7ordku6vKAsDfL+FnLtMoziiBUHo9jm56Al2knLs8lDW8nDao+w+yd0VD4Aju
qggQcyOP9i//HA7Zj28Q9yO3nfGcSRZe24m9PJgahjaVHiZU5RL4d4buReVEMOi0
`protect END_PROTECTED
