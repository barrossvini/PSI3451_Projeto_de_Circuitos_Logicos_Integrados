`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X9MJQU2S5IRIg5tzir8ByD86CbmfDzGTpvmcPYF7OtQBDSNuZrhIyUVAJ2gYuwBl
cw8u72wG/PdZQtewWwL5Xystai9sHOv+WPKKxxv5ozV7ndUpa4gVEihEos//IdxL
kziwafeBwfYOamdvWO94tkHZduGvvCAAxn3k2zEBKqqEc7ZZQeonmr64dJBv+8LL
QNH4V3yxLALJHbeURf8thjRKtjaaWV57cffq360wDz+zheMDwEfRONPkkUyqmcVO
nn7a5LFsR8z8nqDip7oe27Dy3OhhBWW/7PEzf1HhRhifPxPNTI3+TPNxbFvs495N
kdiBkdNQ9S0fFSkvPeiF45vafaGiE/sJxJTC1WyunfxoQ3ofKKxJm9Z3xhk5j0Ja
qjAVdVAJ8U+wN0z7M21759ZZBMYa2HTzQatzOdcOmR737VW/khu7uPcGJKd98CSf
ZbYe1VIZMaTI99iwBvi7Gyus/74XQzSOvJ7ls2p9xaUJNWWRBPwMdg+5KQhysvdZ
FDisWl6XK7srnB5G8xBdtRqVSA7M0zXIh9y2bPNvqB2qn0OTCtCVkP86bKRjNs4M
j/yYhHkCSEdt/KC30BO9s0d6f5fszd+S88kcEi+aj0072Rhx6++EWZ7S8EYVrEn6
t8Zi6UztKbWqzpfKaCwTUUkeFacu0hZaom43uS0XicY/9wa6KoeZh7PjnfuXjBI7
BRprE4i0NJkTrRVdpFUcZcQtOd1dVgZhVn5ohrMQLEZ5KmaC5ssvyT1ZCrVrarmG
/LaS2EU0iqHHQcdgUmyudstH3z9rIzlzf/Yf7xSQjVNeu91ioRzR7o4YtvcozA9D
ZO6TJFNnoC9rokD8hzNdMg==
`protect END_PROTECTED
