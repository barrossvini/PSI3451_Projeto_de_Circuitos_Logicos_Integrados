`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dtrbRIJt31+RNoxoXWBmhN6GilXZ4xryNukKp2SbfZEoDYIBnJG0w1i8VFGg0w2I
Fg9jTxNIwqMmGOHCGgFVrikRINo5vyT5podvSIwm2Vhtr4x4egohK1rjO1yBgyiX
zdDh2oZeGr3zcs7dWa6C+lsddjvQYBTCj+5ca40yQaPVD+K3aTRW7y4qyL2Rd4CJ
kfLSiCRUsBpo1Q3NCIvok0AlgMfL/MMz3/PXJ3tQMZetjdP5Yt/3so99OGQHP6d9
F5ntG/ZsGWH/vF1BfAKGhemGiR6YPINP8UyKJloovPmIsJ1MS7AJ0LbjHlZ++B1D
DEdkyRnnFpgoMj5ZzWbub/zAAECrsbF086IrTzMbYvrGpysdVKA1cNQKXodyaWNh
DZdJ2FW5BJSM+lMOVMLRZ1RTM0K7XOPTEaQF9buOCXlG9bqSL+VEGpbw+rO9Ufbl
lmvz6f3BhyUlLEzv4lgYXtbX3SsMOijazeg2eleZkSmiUcTTiHvpbPn56RLwXeHB
BJHYtW2z1Ac4lMUScXLrsbF6iSo13uRvQGfeMhwM4Od5SIGJfIDHEq2vChBCwJxq
ABOWBxKxvfJ6dpCJsH0fd49Z1gZKhdSv2KqjbvKTl0nxLj8snp59jTsY++93b7DB
zFLs5f9CfzGvBWUqvsMzGUgw9lEvuBxK8dcA6nMvzSIa2g3MkjK8z0fBwbl/ta34
GrAbsICQizPbxjfB3sCimXeTGnrg/vY6rTbLzSqbtbC/u1n4GAFPtYPVJ+ZSs87n
MHawiUbbJA2ZqnfXHOdPjU35/keit6P/wj4+xK45lUxdqWMtPfmlbSiQlOg7J+1j
GG5yX44o1nqQXARwr1qq/qT7f9LDgpEzdhpRKd1m/P2/K/NJeZre6in8kHBOvd0C
DVVOlF+eV7vLKeHGDFoP5aZnqlrIuzgAGgmtCmHsTp6+DmYJSwQBbl1xSTn9z7rB
TKWue7/3wgmgS12oNQKRXkG7oPA26+4o0zKafYmylL9hQPEzd3PXHwFAYzlXxbx2
dYfQLBkunk4u7eLZxXPn1OyynhFQN3cLj5Tl15G42eKRMjJn6fwK5cFl5MbyO4Yi
vMy/ukeEy1nkWwpYeZtbqlnSycOtDIBwmQa+fZFH51AjeoydTh7ZCaP7KNmKCcfm
ZA+guW1f34zc3Qtdsr8zN+PxVglJP6lqM7M3zDM1F6TgkphI98BgfAcj5KI+nzlE
joiqRd1aLrrC5QTT7+N14xaiwsmutpxIL1BVwSrzB/2q/h3JgxA3t2wTD2nWnG7I
LqK59P9nLq6m9ZoIJjIjgtGP5C9FnInkTO8vZE7GRLjIVHUPzGm0fW34QI3OmCfM
afj55nTMgbzSBzPBEhDtNm8335kpZ8JZ4rUY1R8FC2oZZl6GVPD93ssUIHjQibSO
BGQ1TE4NOy+B7CAK3d4428rs2B3mjdfnVu2sb9ksSkazIWBkvvCBdx5DHvuvkG2y
qTDGHCiN0eqTq1ugY6B1F8HTj8xPzSThphmI/+1qG2DYVf5OWhRb1y9uGkKvfo+O
i41bJLm/5gf+ybMIKLxfshje/CNW/bC0eV5hpoPf7sm+OEJDthK8+gSh8VazhyMA
3XA3LfqUe0G6uWntr72F4qZWeRaKDpo9hkGCSVSrMuQtpo4aTbiCAJt6VthePyFY
KXIN/js6dBOhKmrkGliBmXSil8XHDVPjuxP/EnOtxfxfYG2khxmcMVSJ5ZJOHSI6
wocBuwEyWDywAOHL+D1c9EKQryVg/5MHRSGaotNsS69Q3yG4COHRbuHuIWo4QLya
ih/pSt60lt5F4uydOEJmSfnRjVN6hPS+VK38Swdta8M=
`protect END_PROTECTED
