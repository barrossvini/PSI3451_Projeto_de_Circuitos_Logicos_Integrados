`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XbqzlCu8ZUajIFpCP9hlEibFCLArlmw2VENsyh9U5MPstxl9QgKegmN8nwOo10Et
ql8vfx6a00/Mmv41VWX5m4yBhgZPoSS4dV+emkJaklaIlppHckZmv18wue/hfY8m
aEHq3ISZGq5KiiP0TvE8Qp8zkvrfycyV2cgN0B9byLC8NcJ8PLx6oVqLODtkJffY
LEODorL7zq5boBvlyW0xWUWNqRIW1HTKytvu05OI3pSW8NCcVKTl650lHLK9HMjr
W/f+pArKntbpMt7AUGJVAruitvhcz8nfwO14AC6JV8SlI9R3O4XJ5N649VW4YO09
dN3ezH4VoQRSeWChS1utwg40iEf/462Arj+qgJs9tHaIHd6XMAGCbKXbIeSL91Mg
7x2R/NBm28iV4w3vbndSNrSWL4E/HkQxrP3Zm8v95s3yrFgk+9fW+r1fSX52NWlb
ygSAUvOEnd0GuEopsbc9eOqYebAsE8tRo1JA2aLurswSSx52JQEVI0uhtqGhB4Kv
gLZQDE2TSd6yDB1VCwFVXmAEyYTwAN7j6fcZ0G1JERbTuU4VvDZslPOnDj1CPDhq
g67fLSwhD1s1duShK8y5OkuS2GHV09oQsCB8o5RrpIlX/bWqsb13BcniuSrXkf9C
tTKXnouLarckQDoSSpalGSxYn/X1T4wRsBRyORIqDYFQvERNFLzH+ZiPT7T2Q4bs
/bBTfXzf0mgSjOSyqaL3MdZuanfNoVoi404k9GKHGZKoOwUcwkv/5UT7/pR35oAt
govocC5R7v7FT/vEzwaiqKyaXG2utO04dWY+wZuJpBBb5ba1Hi4C5LYlZ+QBc8yb
XDK0uBc+NufKFvvzhWXow8Of/uw+tV2RyjRbR7RAeXLVbVcIIe806i4HPeRZ01Iz
jz77R3ZaJc1g9tjCezm3TSCTLTe8/2phbeIR8bHm5X7UGj3vHWsctCShnU4ldL75
W7lftrIhPqYyuR0d+jeHbYbLUax+R558gNyDFFFr8tniu+e3twQLgsd6GdRNV8Xu
tnpCuMCLOi+K3U/FMwVq1FJi/ltdfFSFNlMCS/+My1jR2zKL+SQZ69e1jg+KmSfd
lIKd59jBEtbd+dKZI2VpcoqDGDwfkvzYt0CdfVUniSl/M+B6GcUc1QfQV/aUz6+S
2Up2G4BECh1WOFOJE86n4JOg1m9dhSYiDxMRrMElFIITTjrcMTb1ZLaa7bi6IMa9
xfIHfPW7LWY4UBO62B3Scoq8YgdVkSb6SDra+jPv4NVGTnmEc73nypIumg1Wfqr2
YThCLZDQ2ncbsPfrxihHQ2KEfdXGjQyph9rQCm48fL8gF0nW0K1rOO9HHaIxoxI5
ul4Rfi+YF+s+iT/mhfLmo5KNmLTGRbMaRVeeOTWX3QlyHMk13luxLFl/QcQG0Haf
v8oaguEVTf8WC3lKkmqpumJS47LYR7CeflKhwESblPfv3Y8sv6Q/a+vO/Okr8M6u
sBanDwiiWaERgF1iGMpAsWKiFJjtopJ9MZfcstpxkhzt4VkbWd8C44ElIi8OO/0O
jeb/YL1EjUeB/BugsuHQkNPF7x4DzNzHCriMUibuPs2mb37AIhRBD3i1xdCkFtxu
mjhXbdEHYswcqC3mfshDzGUaqsgGYv9WufhjqGGGjEHphX6BVAJhFScxmcSq4nmq
iafIl4Xp/fIf5meaRUl2DoHr+pigBzYSIv1frAf1yZ27KT726mnahgaQxc7DSyTP
2tezWwFv2K2inO+OvjYYghgeMcconNifPFAFzM0o/QA8SqXk73Tgft2p1ZD+oRKl
3K83RhoK26Wyo3JRvzhMyG3jzvtq0HiXDNYMm+U2V/LyKAIYcL6LzmDBahVDhgsD
iUi81Qulljh3/RgozRRlawl6fXkzWihFCIWSrPpvn27uM5wGgKZpZpjHUDMNvxON
4A4ViRo8L8mVzCIJc7pVyUZc1Y/uX0/vHvAYWR65tFwrtn+9ZyCHJz0LEDnI3aCp
tv059nVDAkuaMIPeusHKaWQO5Kmf7nzhL3+RBVoMyK4pTUygdexmrwqimePtYLth
BpHQWZqlGeHpeaAKYKLfL8FCswFjgIrMv87tWqqROD5xkCQiIPyIv/tqnKQfAVvF
BoJlu5QAKMN6GtmiKmv9GFXvRRzpKuzDZOr65Q9WcyZCfdUQtqXgXpf38b695oLp
/p1lZq3fBEas7SFww9xGICr1VTKtfGp+ws8vplAZ/wGJRA8ZsOhhOJRHl4TwHfNh
NeWr/956B2cgK71nIV0xxQyz9f6PuCo1t1pGadyXpwHz4nuGqhwiAArSXm/3Njb8
3hEpNhBAhAr0ZXKAiO8xTu0928v0mwZEnEk5Po4Q5A+hcop6FVCKB+r3tCEoF8h1
p8TNxarD5iZRdAx/PYvEdgxA3QbmVi2qeeWzAw/boxQgEoH/qlv1Pg+jteQqRc2j
jfHJUy4gXwH7uY9ToAGLhcU7eqokh6LQEhGMpQA00Kdh8fAMrDItfug5c5FlFl+R
I2KSHRWx3BD4jKsl+eq5Y7uu/M5dmqPeK3MmK+NJ6vdeFIMbCgHJ3B2VRbd7Acq/
zYheQhWa4VHUjC3voaEKWDNKCWP4QVBWFhuuyvOJH72EiYDzeGmQHEAp5WiP5AZB
DYeeiZlDHU1HpBVoUJuasxH5B3bHlYo7hXXrhatbM1gDUWfBns2j81DHqm7E0hEL
24iIddqSRyCfr+gtYyLqfUlXW2/S0WoYvGD0SHSuH8464znIMl4FLHl3zcE8RcsO
gZ2zqNpaTIqe1SbL2JP6PaCcipATTfLZQOo/t142muo1fs5RkL+E6XptAC1IfvAi
w8s7wD/vvu8ej6XtYpcXX0p7qH2gi5c3OhXM9KJQqBEf0SpURZ6GE4pPq37Zz9Ht
1FMPYDHGQQHQbJdGeenkovtAvdlFaVpIGlWHf/0IZ9d9G2GEL8+wMOmunMg8I6Nt
3ClBXI80jXiWAinJgjZdpwdP5MgBc43mHe+LQirnhDurOZhzWXzwspdIUa4Pe+0Q
NpxEPxwJ3L7rSa/Aii/J2sV59gGMUHsQpRAE+k4FNJp450LmbW+iJGGYGWaWKi50
PZEpXLJCPsOWODqY6lnZHASK7a7XU8Zlb4NoNZQ8NIk+fgpUHiEsgNau5yktu318
dii+8ysncAhWqZFqUXWrnzZJufsCBO0HoSymXJyC9kIo8j8LuE1XO+quVJgnCcRO
q8r/QhuNe4YLJjLDsVFgsCSyCbiCalbTgiEjOK0fD2tM69nmR/fPD/0YX0WHIWhf
EvClCxFdTxuHRnhBTrcg1AoFJ51g+jj6KVQkcwj2Y2qfAU9C78MH5Xuq9uBjWgwS
Gb2N36NwdxQWEptoVjL7yPqT+uX74gZpUtrUm14ntBVIWDKf3gOp6f/2JVJMnMkC
gbiU/gEljuX+gU3F/Pae1DTLWMkO8usNtuGpTyDUN99MEGvX/xmCBcSul7LU+/UA
WrcDXKOKTSPVhpIJu1bC6m8Bcbax5vTUIwRvZxUPrbxYUDCd6j0rYiCD7jMhKx2e
wylclFtLWhl8N3aMh0k8vF3cbSyPAY01so5onsRZoeBl8Y1Ytto4dvOJd+CVWFH/
Un3j+8sygnLanTwTDSj+2a10ZWxb/IiskMqnmd8h7FzDb7FFmJbNiRPam0cYDvt/
OHRoj/Ubop3+XvIm3o94kKlmFk9mdA4dO7PB66FTg4Q188npiojoCjpVt6rIkk93
iTmdij2q7a4kQwYjAQTb5mT2KH6NNg/opARG1q1Q88MoVuUtizFZ6s2fR97/66Dg
urYGCfNfxDmbfjUVnpF2BvejMZjP6GkCmBfig/UYXOnhzL4WPzcx3erO+8FKQIKu
OMZSFGVCLm6hkRqUtPy4O2A3mPojPq1KEhagpeGqBmwVrHHz/mteehi/bsAipOih
CFXMiR+IXA9aZqPmArezhSBomR+oXaxudT3WfZabVFS15PcIpWwcgao7Uvr7yiyu
X4Y7cm/LlKV85u1u6YFZE82CywRBW+FGNJGJsS1GxKFIN+9ceEuo9Hkzyw1mvAXf
m83ENZCqZwsMphaZHyaZNlrjJ982rNhb8STKRXgLw7BpQm+TTbhj3uipBO1OU3YE
8XRcg28U250BhD1wqvvyowdKMpykhFbSE5l2uYsfF8Cnt0VQ66IjgedrVCIqUaGX
M2pUgYN/BEu89FEaI4qNrDgAHUGswr+FaqX2Pop6XhwTx5j0gZkY1NXFPZ6QQ45+
N5enSEPzG+IqguKhyMWnD3Uq1E04xqLE09OwonjHoUBVWhEDIb/YnzhRBxRST0uL
2UTBXHZKAhw55uAvaXiz4nLPbyJVycZ1oeL39V0tu1j1NPX/nINrN+dVO5Sw7ybE
XvLoHxMi7ZeabvSqNixpma0Rv+D3fo0lzDyVWdmls/kqyMEgja8k5ZD1a7eyuqLg
/R9x5udu+7DW4u7CgxXG4lkONw2JTltKCEfDblJDiDLwEUdSRrPpv1V6AHpZ66H9
CPyPYn2SWDUNcLxc/YcgfLpx88Pckr4vUQOytSgRAT++uvpTe9FCVGOipyF0pd+T
dbuvMd5m2DsnyVRjOjEHZ3+gUFVLoRFf3xoJvklSGN5WVWbauXrn3H1AzAmxsST7
eyPt/ghxaDsTFxf1UK9SAll740sqh9Mnw05BALYhcC5ddDBZ3MaXmXiF7GXI1PQl
qFUDPERw4oC1t8LUxJfx7h6oi7Bx/nN2DIlyW3ixx2QTcKd7eFgEpe8E24TvOnMo
aWjM3Xl7kxm/6pYo3ioGbYzA+EWlt1K596GiC8Bm0sZaHcwiNgVh8JVaLIA0sSlu
6wXC6w/7gWX7FMYAIpcpD/lFHzWoXomam8VvHUK1jXGQj6fOxUr297z+SGBk2pYU
R4tD96sJ3bwWg2keDy8bXA5HBGAh6VhHW8LY+lwS7RG297ngh9uYrERDZN1SAzC/
wCTnHsGZGtJUPWj4E/TrhF45UUwglGjcstILioIYcrFTGQJV1A9VtZAQ8hl4PB0h
IMs+PouXtnJ20yn3+8A5Dd/8SLHWAOL7LMJxv+Odz5A/qNC8kkLVm/uS+x2zmRMl
hTXH8nQjB8hgqz0OXzlLqRGKPUD57W8J03GeVPfUXtRTy00/xDMp2RgoA9UEM2i8
61srswyvI2Nbtz38UStSkS1UzwoXd+9QuQMyQWemtluCs4UPGsJT/YpRuBJOlQ9h
voGXO9Kv0bE/lmIS5MVikeHb4TcZoPbll2GfDXO3MC8IzI+ByjM+dJjasIZnpISK
0y49ofcZM2YUhJHL0mjWCC4IS3TBn/Xuv2+Z1blKVG1r6t2dF2pAQVWbwJ+ifTXS
DTBlYxWuy2VSpuGSxvfV0M8hYeWr/W6wcSQ33vbtNuaP2odCQ9mumXGzgUY/MRIT
hJQAYZcYk5oh6Q13qKbC8TwYgAtrMK87Y7+554js6bZlmnZlbvtqjbD40kR/0N7Z
/1y2an3vLDHkWhUkB5Khew9pBtnbTusloX/YDh0jGjRwbReIZgifOyuKZQSPNsbF
hG+HlzlrgX4U/rzQrYnUqLSQ3qxcCh1nBr6NFMGvhCGmcEyiuIPDslwYR65bEgeO
tNYzFfORe3eg4F6LpV4SUogpYJY6pE3lBMfpgq/UWbdgMUXuLo321Q/fO8kdeVQt
03AllzBzAMX9qTSaIFvfGco8TbP3J5QW+ZqaNpvwBmkPQ50dwwZxf7u0nZXhzqXX
ePYQYgC8NUqleZMvgnhSOZHwYFBE7GGFOPX8ERnsx7mQ0SLmFdO0ErkIJbdvuqCh
2H8v9EuvzoryMrcmoK+amEzc8bRUQWtvcQhTic/7+oul5K2krLN0P5vqBC/2bmyc
Ntgx445v1W+b8XGulr+01En69YHZEjnoMQeoAettGA5cpcVYdmQ2n891sul6MmS+
Xpck858Dm/tt78/sFZCLaoi1l2HBpmXYDoqF+ncv1ECpVuRhRmX0SiLMKgEP52T5
H+8sAuBQlUtJXcqr0yXF39lz4GDIggukdamSdiVMWRj8cQmQ/AqOyU8eq+7eHDBN
mEzKOETRg0Q6dwubdWly0XKp9OUKvfGpQsONq0ZNckLKMrItE/vt2KHB4HKN47X8
fDninlVcnrcnk8qASuWPgm5zUtc7tb8A9GoDb2fbfSrfUsc9CiescVaffq8qcmLv
/PmNTCW/YrGPi9eR9t6Es5G3yI9s8JRBrzqOUKZSr3A18mxNYmTLKacviesbccJy
RG+KjtQnByTwbtKtLuc2B82tqiu81Z+iGkBNWDsZW9VCm4ZlrANOO3qKv1R6dwCe
NavxOpYlknDcAhqtLi0qA40ueJOC/6pofK7ehh2RdBWWlYhacu+PflxhiHuup8dF
MAnE8ZgCzU1AExtJdniNYRhei6khhUeoe4hzr4tZRm8KLb9MDb6Uk7nB4j6EJqPj
tImyz5eEfOt9c21sd+uwLugFlJliQcm9qY6NpFQxrhszy/g305m9FT4L4I9gb+KB
JYvjPFt7Ba3twIU1ByBEDWDTbkx3aYX0QHH7kzlyh5UDxM5PrRO9IROGbfGJVGDA
HAfbIha6qFT8IOusu913M4xvlgNQyHaidOnqJbBY6IyLUdqFw0vx/dZ5KExbADUS
WhF36Bg/C3boOx7v1F+3TgId667IRtoO6KW+GUjjBeJibJy6JtoMm00TJ1HWwZL5
oR+GQ8OA3RiJIiI6VFS8LeJMs3nH/0X2H1mm+m9HY078pStma7lPXYvLqfrQI3Gu
Jfk9USGMbI4YlIXzb3vp0CiezB5+Yosn7Ac/CYGT7ajZsj9yUDkYWeMutr1Xi3nD
/twMm0RAMrYfyXCcFS4DGFK+toZkhRY+uZhZ+xUBiWgih/FGnqBNCDySI+vYBteT
oj/J8XWb0a3whNipWuialy17TUsMjLQBBTCxEsDx6UgtTBavuMICB70LKCmUCr60
cbhed+NlVl7SQ6wKVbb4jeQPM4P2JaOrNmBb33TIjO8QEAsSyBK21/wdFlC5RL9H
qlZ8jjLvdiljwd+BrMmiH30rUjg+eTSSgUIYA/soQ37sjn4f0vo7mm8HyKiAlcrG
e7BNXeY9KofRwJD+b1FW1ZFIYdjtQdejWT1mU8/edhmIztE7LiCO/YakwXHccMIg
LDLFTZhZyzutnqTzz3qijik8Kn4cPvKXKfZTxcFZ0KXlHXCRCvpeXhMEF1i0pkKg
AhS/TYHCNjehFGJ+49PgnMiQFZ8mmuYEgSibwcjmriR6KUgYRkccM4fmMc66UG2E
c3lIE3U5XLyHZSZNU/0IfsCaLPeTtev8iLcRV54pEdCT1jygr6slPs77KkhbdS/H
jivxaW5f0G4r6atIz7oCGt5kK6sa6WQAHO956weYuHqE6j8303fkDP3LI9Yyay3f
ovjgdNfDGdCKRrDJ/zt+NgM8JrhNQ1/2Sy6vlBVuxKWuDaGXCAShFkHD1KcN9JYd
jVrWDUTNdhQmN4naMd5Xm/aag78/1lcEVvv7c0M5DzLEHN2VUPbMZryOTKlGA82r
IisaHiVpJWOZUuPWB2CVeKS7JIPV/F2t5JgVWSsehtjm7OM8vt41IA2H+TWO8bow
+QSUqkvWh4DSDIsyhMssKAF94XK9CGroBbpA97fcnSXq/nhhwI36pvQ1ERZdLP9c
kTXUi5F07YASd/XasBlochvA4omnqRZ7KkiHVuLo88Sqw2sT9q215o2Rndcy6uUq
d/75bAEuOqZYk2MvpRHA8BUmckj2+Cm4ljdRS5Bn4rYW3yxNXAYvqx0PVF5LyW2w
xb340ZjaNbF+9DLUx1DgKv6+N5hlWqRdITaoziWz0fw3p88KOA334thnFAXgbeaR
sl1yDtC2E8WcZ12AAmOUckT9+8zIQzXbwDYGKDj5z7130bHDjyPuCtyrObpd3nAk
vB9agQGSmz5CeNXh2daKlF5jmV204KAGG9OG6fPJZoF9lpKxbiOSO//3GiwwylVp
WNhxtTQtGk15kYIjVyfuhN6ehm1N5RP4xuqPMVpW2z7NUFVd8AX/LSpV3HeHhvih
Et3+mEF0Y3oyX318ZFhOVNLIW1rUI1ajq6vI/e/52S3f2go4LNgjw5PHqUUj46dc
Cas3SaPCe0G+f/IVpZ6epaIFq4XsycDVj/PAhXv3REXqOAECkf4ANSaMRQ2MGh5Y
sX9yLewNOGXdbAl7OUD2cRhLIVB3t39wu6RImK5M8w3sFKBL9pdEvAc0rOiuyrcZ
a4qqFgUuaw4qVifb88bfx1Vxn/zVbEklOHmo/yL8mNz2xM7yNCqjIywdauUR4ScH
xUv+TxXx3CODaX9Kmv4Eb8DWt+PXtbAA2FSGSIKpNhU6cnyLMVjQF8sUpKNZyeKN
/q21WuP1Owet/co+MRx6mpo940/KPbguigse/qID2j3e2leK8FeFqAX6AS++3gZe
ete/447HBeBbrXenaQM3L+R2RVyLTmbukAPOAo9WHd7XretknlpNxuNinEQvD2mm
YjxiOLPisAb81LLDkt8SqRonE+yCCJrBgaIRixLIQ9KTfiR4R1GBKc3dWoNLLfX1
iAeqZSaBbmqYZSfslbDTwCEUoBQGNxCsfk6IDRiM8hEpOEwNMRfw6iD+gY6dlJhQ
tZqZgBeO+UbE/0NkiKFT7ja4bK2OB8vWRmCFz6e8UrRuPyGI82g3CNobqbFfTfHa
lmAzW0nD0KwmhSFO4EtNz7WusPSPQPTpgOLcHLzvEppDSWcESvxiR2kTiZF61dZF
SlGT2Taul/uf+/gBbebbdCGWCFTDyrh1bCj7THW4537OsgRnkL68BLnftQDCq79F
dwsRH7x1/qYBwZtcfVHzNpyM6us1/HjcnL/hHSbMC00E07grQFxhjxx/QxEPCz2a
QQDPpkWE8B48F0RQIUkeE8nNO5VnI+ICA36VYYY/yzclvCUZ1wezV0HqYwynrV0Y
R3M6vyb3saYHXauniiyYDukZlC5hPL7EDSbOY1NGPuqifwxIKXvnbO+XZIn57cWD
5F0ZHKu31qC1+/sGFAljMotJsP8FbQOUU2qtBhDIAu7v+/KT18gORSKY4zWDAVIb
LJvlxsVRJbJ3MWp+PAnTtycJOpTZT0kMkfAHKjYNFjmLpAQb0u+TzyqkV2nCdsdv
bJmYGXr5SKgsbe3llVrMbAdsoub9khHGzIYMEseB0wc/8XtF91L+uqaUSKICZptO
tjU4JejFiS51DgrKTL4HvWf6GTjxU+gdC9jt3SMwI2tXExIN0Xix4vcNT2+27DFb
DyATSCBOFF5vQ/1bd++diNbsGkHTlw7X/xO/1UuW50FbnBlpaMFFQca9/kZMGwnx
EdRnw04aX2h/JfaVw6m98UBLRXdohFH9ymX5qGNsLUlbueXo7S5hMWx+0AnVLvjm
ZOnMT1f+byKrL301n93MkfyMWDB8t/jrWvJxh2WKYDFNgYNAxA+bEPVrKAVLeK1l
pcc1afyjOLidCJfk+EdxgA8Xqx0OlgTfPDm6cfArOpjvI1D9nLZui3EMS0kn5o//
NTzg6ZxJ2zhLuNBEnAVtov2KlqR66grE9t6fMhniBDcJ6+9uwe4+KG5+4a1YXIk+
P0mx2Pnv2yOURVPT+baldrcQeGfJYKBdXd9OMDvE3d0vljxC35fLW85c2zv/oI3p
8XBFqNBx4EFlQBt1VB9NRPSs2h4BBpjZZ1BNh8NFh6lKrbdnfOtXSLcRIWAHyOiL
xx8rrveXLszizNLdtkMsGFQS1JnMwCS6lscRiJvCZ476YLuF9V+OtQJW9vO+gOiV
DrnpTL4IyU9BBI9yFoGMeTJgC9/qNaPkyJbmLBUyGK9FGNLFsircLoM6iOjfRzBu
lMrDDwtEb4oQjqcGh2gEXvYedfNq6rMTKhbxZspCUv32P7zrI218dFt1L4DS0U21
AjmSUNe5KM3QSh0UTOgtvN+vNRxjr+v+Xzogi2L74XC1JYK9dcobyWkrhNqC32rb
SdUhEb8qq7pRpSOJkBrS6KHnXCpD4W/9+qrlGvzYLSg7bCtya0iLARAYQjNkOMSy
kJC29Aqgx5L5/MKfd4M8QvJ3Y8cwFpptgUCfDFzm1H7cbDMlXKZlYUUoW1ERcW+s
jvPwX3HSAR7x0dD04YgsLf8hKkLyu/BTnG2/l19BMQOQxIF6FfDVLwjrq80A2Jji
7/mOZZdkh02VeqgtlYv7clSHDm6jB97Dq9m6UAibiT3JA3/JbpsZ31CBU7SeGgBL
cS7svN1CaS6NPDZxx89FkGnqg9dEZov1l/43/Fl7qNmres0RtBKoN89RIDThtfyL
OUiNi0OVKqyOvQPTuUHw89jMo0smUbzudoj4ig2njeqaIUpr3x4GNDputB9TJHs8
VTZqvx0vOzdF9p48uVq1Syr0kHGWUGQ8bzkedN/d5mSJQnwuKgQNYjogOl6aNsF5
ocH9DKhbKqyYvJx54MfgnX1KQ3gFKCAB2q2lJB7hhC15xbT0rTUn6XI8bRp7esGo
Ahsh1R5YG/CXRPrXE4+3P/3HUiL2a/idBXveJUWKCJtnCamiZN55hIP3vdTFjdQ0
9mepRtmiwrW2d4+7JnZCIxQfiP7TJ3T396XvXgrO6Q4YayCrcLHPRp0F8an2bNQA
inCShcujMy1XwBvnrg+yvrydTrjLCdNPlEHeapePorJXChK8/NHKKmBYby8tr3+T
qQUy/m08yAZ80uhwatMTToFteTEGGZEcQH+YhKM3L/lDpOPwL8GrY4VIsx5mDjXL
YE5YO+fNXYv5qosh2V3dwMBxhv9Ym39wFr6U9Qi2qPX72XKWY/WCTFmxBaXqIzH6
Fsr4Q+RjOk0WllD8JVra9lQKn74MvQbo0rHf6Ch2hv4PZsYJxGQ6nl9MvwrBRhf3
Kb0zYecKDhg/4eif3U1Jo8I5JSN2ZiMUbrJM/vXQFEJ4VrSnX0HZFkM1nFfTU7DS
zC/y0dhkljo+duZtyc3x4WIFDV3LL5Adh+ofHopecTcUgkZgGTitHMLtNWFlSwGJ
fx8QxjtEtYKH1AvEXRDwfMxMqgS+VxBYR5xBhZ5JJ5VAXZuWaDVUGN07Vv2oAdAY
pTnFItDp1Bb16J/MjV2C2SojNzCUJVrR/lCv1hSh3nyW5gvBYNxXXCRdk4Xgd7+K
s+Gk6N47vH9YXBcfCDU/m3lvKCsfCiGeb/HylKmnTZqyk+82Qxt3BDKQA1l02Tav
l4wfGTBOTMjisHSxWSi9+2paruy78ZDDkAjpYhwDeP3GzbvAFtPhd8wQxRuv9Kj7
ytkE0NrWt0LW5Cu7t8o4mmO3fTxM1fsICF9v3Yuett7GfC6AB5Q7+wbz3FSR6/om
XVZRLelhvgJz/VIhw1P5LJV1sLAG+PPKjNtv9WbN6vQnlK/3B4tRAnq0XwiJT1si
r2AnqoCHIwwLA6191VDXLs4d0wb++GprAIj2zRO0tjJJtFUkj7kCEEA7I93d4Lkr
NgQKr4mamIMZcHodyJpdDh1qnQ0BY4PDGvb/oE9TCiQNLMNiH1itSchDd40NB8KU
NcMUCVrn2d/4EU9IVC58Pv6+BB0yuyEytuBpV2rKDHbnTuDXhmNkPM+RJIvr8jNr
2PELcd56OYYbpejWQwxtg8szRxYR+auzhiIgVbKW8MQ8KHckUTyuIpqfx09PN6L8
wsnwpwrL+4AOgcb9sC5vJhZAryiqN4ppZhp2h0BVmiHK5gyUndB+WxJbzFfIX2YQ
teuOKXwH5BdHYNLjY4l9zuG1py8bZ19U3unGgI8Dj3ktURblrewNNeZYtAmDTgFt
lJ5rggO8CpxqwIofjIMgVIajdzcQ/1ahSFVv7yzRPlWPhTyCMZaPVLMQoFraFH93
vJP/DPTfUDs1RawOTTj+cH5UXEy3yGcgMSBfmcZsH72po3SnU/UuMSEc0SMKM//d
859NFzlTQWZgA77Yfwd0YCNvxWXBwiiN2V2w7sY1WzLjE1yXBjOWCy75cXNaiPoz
JIXJPp84eQGSuVeYgXbvjjcAfk/jmfoAZDuuCQCJLuSq0rJRf+siXUjkqrpHYeRL
b5BCFY1xpJ2573tGVTZKA9GwgNQtKuLVeUDxnA+u8kgxEONy/pm5aCykbuykukcR
a60QqC9ihITPeYgqcbYe0Yq7RuvASTwdqIAjAHsbMHc+nxAvhcbpmr8pZ53jUKvU
7KQcsxMyGccMT9V8UesfrQ/J2avu7qrhxHP9FpxA9t4e0S5h6sS0SV1xzDyP+JMr
GPqxbL4O3NaNCseYnwcW3NoTGDXckkLMQzftHa+xqhsS2hommqLXUolrRmJUu/9I
v3A5C4KWM2tMK3y3h0wrtDGCuVS21xg7pJGpzF3zNxj08VRXQ2WDcZrIadmhZLNi
vTeynG4+TIdbhJa/Wy5hbt00qQ43+WwLAjxlbhwJm+hC4ntYGIVD1md2g/J24lFO
pcx1wpAsa0ngtyK6KkbeGYrdWI0q+ymg49BCwlQ2mRi8egJjPZnE8B8U5tXnWrUB
dcG7Wn1pXdeme7rp2GmFs5BSyPXjfWhNe82oEEc6b9j+Op9d9CzCHwnvlS6waf+d
XF9mwaXXjEAwdQVCnKpAXA1lUeauAw6HALVpj0jtrSi86wmxUOEpJfZK5ci5bRNU
4MOyrJnZUAatAh9A1IQVdEEpzwmDfPLUZmeQHxTrO4Ke7DqpZqmPRZy4hBBMf4dp
1HREdPpoqiGglfMpwDkSQJ0PJZ4sA00PdVCKRX0QEqz/32L5jXF2Mjwi5MsRYLy6
AbKioXuTzeeFjimm0rZ7iZJYgd3r6t3s+pQFpurwWpMvaE32lquz9ZcghUdCGJ/k
JiDAQvkn1rHSwXXT0ia5u6IZYC3Mzz8RVxxgQFRc7zjOe1dC3JjpaptQIXNNy+W0
3jKQrXiB+j1s7Fx57mdIoAbtUBZudPPi3rIChUakCneccJcEw2Rj4rBKiH/Lq1xs
Brgt76Cz+GNSaKCRq3VpwLrIOOL1ocS3ISdHiyf8mHcE+T57JTVfphB2wi67jwaB
nNSJ8V8b93pSnauVO4f/Mw2DYCjS/D4IETxNxdQIMyesKtPbdBMvqQMoTEXNIlO6
B8p3H1RLq1/TtLppwXGcSrcOisCygrIVMTfXq2y1CcBeCI9iiC/vbjW76fixn7QC
xjLe5GcjYFgz8EPj+p9WTSNBe3FZscuJkC0KEBKOIH/Owh9LmhQWl6YMTP0VfvGJ
6Ag+Z9PLIViCA0vPFSdYHTyS9gbdhZI2g1tjXP1K8lM0pPUv4IUs9ZTCPh4MqMJH
3N9eKpWsiVstc5hWWANgHd+guwaaQEKlmAiuwxROSdtAOqxA6CDIVTJUPVW4fgK2
GChUd4Plbpaw+Q1vvbuUvbgzCJ91zSzvR5hLSoKUWCrWvFCPzZPP2+ZJoSAmtHzr
gfDFUi9slY77OcWrJ5Sfl19hWKW5U3Oe6XQIXEVLrBb1qBsPhKy5M9Y5GMIMDTsU
9ks7DEHQWnaI/krSe+GCkpbBvPmUiSTdwogPHtDc33/ZTbsbtVI58ez2PMTWEqjI
mLUxfmNXqdZ9rOMCv/0GlT3Tgv/2bW8k+QL9pzZzKELXaLjyBAQ0AoN822ME8Y+R
Mc7YixOhrkOHuSMB7kZF6pjytCekUhkybzGrUpAkaurwG/fftAN8NhNxPqyZBTMd
+dlOPeEp/kU9Q3Top3jp3dKQ5KbbmZu8a13nKaybvX2GHdPRHOetzgZtpytu2O4b
SaOqrfeDfqrvhkNpb/wIfAEIpUVrERr+ephxc5ZiEZOBkew3klw/BLEWMLzIPL1O
OKdhyEfrQ1bGFVhfDBEaPOPyeCd8DzdMY5UcGfrP7VbNDtbVgTeENAT2D4TPsrYX
kgG+VfcMLHEyA6b6JE9ZpvhJMnx581FEZxCDHISQKCEUwt87Cxa+xLulPHDg9/AO
tCx4bhJq6o2lTfqB6VXS5Jp4fba5PjhQueRTGrowbx/lfMVNw9qc9StBx9pEyX/+
NyBGcwKGrPxS5hbAD6ZseKFH3+DgwCExtMV0SGgCxBrxzxJIv0wVMUtGjNWJQKbv
mfuP21HHyvC008uDjACHN2UnfvCiNcdavHUrlIV1AOkjH19CnordNkX8y13cPpmf
8icAsuvcLHu3kzJcDj+JHEpsbM/SCPUaHWwY67M2H2LPOuQBNGpC0wLy08xX2/kU
pc4Z5/VGPPQ5CmlqHQSJcSvxb5sptVcLh4H1YbXOohd0XcO4t2guxjbLJCFGjcrB
4xgPH3qoI83JO+SBN0gkD7TCoaREX+TuEFu3DjusbZcgmxDXrL95QmH64GNdCqNO
L0NOKGnfGDQqPthGD8rTQ5mOqguJEQ/mRY2og+HjmFFWH8RJa6Ujs9HGpNytCNRM
F3wmALhFjTZEG9LPYTTXNK2XT3tU+pM6tTL6hEzCQdT956ahUKuzKnji6Pq96fxb
DdZGj70cT4LyHc2EomLxdUuf+sfVemOOZ1PHS0VBcHT2gDhT4F1nPYpXC60kpPQ8
yzf+JdgTQcWigiQTpuq3gMQj8LO4ktsJGRVQ+P/PmFPeMFKmIjtHUCW6iSaTvjFg
tOOp0eIBx0N2WkHwvnEOX1CqlBnnohbk0SUA/juKQMjgOf8hjWPuBiu++t3oi8Ws
Mky8s3XyiNvgxLVIEaNYdWt+MGOUCKecQ/yNr3RnOwdtReYSu1ZfLdiw+utju7Br
C6V9A6G4OrG7XRZ+GRC3FinjmMDbXduUIGiMX77/RNmPjcxbiIUFGnVPdbixY2/6
Fo0VdG0uuxfgSSsZRT3pqcTl+TIfAsyJEnROwid4vHRIrKU1eWJFGqMQ/sfFQKM1
FbqitqswvPzsMsEfBGDqkOxmNFxq8+rDXbHNI3RZw3qeGA2gfcjTrm5Cb6UCDCl4
w/ZbDGGkhBFGi6aZjyLgPqw8+OHroFg24j/FtDuy5zcKt33NoaIzowmtFJ+KvbNy
auzrpyZQfFM5pAn1+pDCBUqHtvEHxJL6ORyDfx8ICc6mxMpLoI/y2GR8yu8C24El
3VaFwgNcItEtDJydiFJwqA4M3c1FgMN0pzKqc3fARikjHrh6e3+MPj3cxBzl6dSq
yb8mXpuAsMBh0BcCG5TjGRuODFBx2UIV+5E4KJiAvyRxaxqN6JhXrx5EmuQd0sc3
hHRYQvzzhrlmlBXNcUYUQL8NwHXkAH001CRIOycZghd9mh6aP/P6+u2Pbr38QXUm
YZ0g1vS9nojz+ggdjxjrIPenUqbcpWcA0hwJUt0KhiTouCGwcBCTwCS0zIhVZ+xs
OtBAmM9K4WTU4v1PB6v7FLYqQU1Kkbl+vfztCrgbZ9AQoNBYJX5CPQ1WMvumltaX
9uCBMo622bvoQT/T6YImujppXf1tUgqfxypVWlNUA8UvtF1fu1Tit/SXgQBCC7Te
PM/r7XSqHVXSP+3HvkEDsSdFTcZ2b1F71LoX2hn35ros1EzRSI/1YfG+9xjPS9Zk
h6wr2FkMKK/AWBGARUQSsWa3diZf9mpiwAw0xrR80oPqZtPSIpH+3T1rLQS/2IHr
8hfyf7FcTfOHIvJ42Uj1UddYX88GFy+hN4YbUX4qmYbxQerABdUODFMu00LjD8Qi
uxmlbFEy/Hc48XSKaPi/jwh2InfloeKALpdM37MVUPVxievM35mBcKd/EzV6wMNE
is+kffbgpQF1a7WvfmXD3k0HaOoD4Is+DIB72IomonEdbIVTlW1kLMMKTpvBI+p3
In2W2OGeIC/ZWLV5LL9TjvEqnU+oY1/W8DBI/CB+TZGinlPx7x+fzDR/QOIdIUUh
C+ecT7tzC/A/id5uvJ2apBrJx8wpX/9DfPNw2oA35Th1zL47r2m2TdbOkPUTPni/
+2V/FqylEh31oLiD6PlQoYLOSOqVBspb3D4RgC7Awk3Md7rC3U6zjxUo+PYXDWLz
y6M4f5pyGSRFcZYcSj5UID0eVmbFEcPFbu7GunGePYs8MPTIe15xVoKgd+y7gxYK
NjMdLVzQDNXxgNUaQTW1UartkA+FwvHHkz7CaVKc7R9qnd11rD1kXS7ra0e7VCig
KS26mKpJFV2o6nPWDQ1XYzVnnzef+VIgV0DxDTyYP88j5p4SRm7wY4+fbq1k6JST
s8sYvXW2xThtvyoqf2AMvMz1lj04+YCJ3p0UzMf7UCBBKiFjOPLB98W8vNqB4hb1
jjTx6wLCBkMwXaMQc/Sl37XunMY95RzoMZ2d0uF3LBzMUqmoqqnxEniwfXVmQyRV
ImTDCkuK50dDT4QS7dvFKIR2ZOhwwo0bQfFhCwxDeq0cJtuAceujWZN+lMX1TRW8
dMpjFyzPSXbADnTIFhCIITwU/Qh8J24rKla7U9uCyZRclIaFAQdkQ7MJ6tzJfEX6
vEtUwSWLsZ2fM3SuKe3JXJof6FowvA32fzCy8MLURBKozZGEE0U8Q4YinJmRtJov
fWLPQkpnu35bpp3cJZUR9cnuQzQMCHnAt2dMedmKzfz4bQXxxXXtYstkBaPTpU7D
5CD3tvPBwT36zCmg6oGzslDTlJPhUiDhmPVl2mRP4H3eZglYa9efJ1cQ3o9jMaUY
FekXs8w6oFZbiEw2ywjlu6nRO5vqetQNvs6mJDhWZb379+xJpbJo3zOrWsMNNj5R
1k9yGBQVKm/3Ii4wcarf+tLq6jgjtcqQvXmvdQpxduu7gooL64PIk72zZ06pS2Wp
vxaxCp81G2upS7cCQpGFDOqBLMNchuyHK4xUiQ7IVF5d7mej5DVsNdWzXZhMyGpz
BWFgv79BvfMG9wveL28/gMfVmvlEcKnl6aJbN0VYu3M3VOa5eAAxNn1YtG2tL4UF
V1dSja+YdDC4MnOV5kbuLYwPS1gIn9SZDQ3tVjFMNQipzjYFqSTLjAq4cHIjEpD6
Ej3OJUaBXSzwFRIilFBgrBXYn5OLsmyU4aLZKphbKsHqP5WqqCASh5pdAfGS3SFs
Xn681eQGfGVAIQBcuiyMIRb/HxYIoOsvo2e102/NmCx0KRJVj/obrO8gBEmvmHb9
LiIJhaGjTE4d9PR/wW88146W6JYsF6gcItSfNEQFOKmbpLUAFq70MAgIp+SsCu94
5qqAc5vLjvsimQndpcc9nYk5e00rZshr60vQxbhskN0ab4qdKV8q8ySQ6OxrlJvP
VUsPhEcaeQhs4OI28zzQQtiehcZax7dFE7bCCeSAKKo+mVgPiiI0n12hCI63dXoO
1/na7/MFAMXmFZGMmGs933CBYte+A0FVuZy3esCh3a+69RWHF0nV0JFr6bU+ShVD
AVjJ07xGGw8ka2ymx1dsMDYutv2ZlElFav0x5kdLDxBLW3NHU3ruYj0ZPCPGYObB
R8Az4I7u+Gmw6LQ9g8dWajgQt4te/fw7bsUEQxR0PFCgwm3iIoLbEoGPHXysjj4m
8jpnbWF/CRrfvBLm6Czio+Ss+jH9qSgSeBf9XrmdFeZJasXPiVHGFpNLFBuMnai+
aWkr0Uqm+c31h4vdUHi8PtCUp6gXyO/T13Mb/IzSUIPkj/AH96yOhMLi3Iz0ZP6J
ppcO7ZXN6n6PYhnUgoqdYnntkR7aT8n040ZFLxNaxnHtBLwWRw28nBrYGvoN/ZHu
BRUEofgpZABJgogw7ejnOqBTjJEqD+Qg29fpijefJtk/WY8NaRRkPOA7HSm7hfeh
g3F2qNUDM+KBkBY8Jy/dyWQ5m6Ny7AqiLwgKM0wu9msLZ4OaZX3gHMBNW3Z3sqa9
kf9OMFEZRfFZkNuMjVdTLN/reMm5M0myZWOkoHk4adg8mveARNK3Xa/u0YSEz8Qp
U4doGRpwLjTb05GHPQYzONzKepVe+FH9ikKRFNCTNlBdU85Fit75zI+F7ORnnm6Y
fTeojepRcjJNN8bugb3D1J2pN0FyvUNfs0PFn73ntvya95UpPaCfaLWcl7W1M4Xa
E87Vpbei7rT//tiqs8YLroBtA50c0OEIuUCvZvrInHwRWFH84BbYhsOCqv1ueOaI
qrVW16CTz+ipxPFAm0g9LtgaTfu+UNfq7xTimAkFfJ6W0f5idEaPzZz5x06oVel4
Sta9LbaTFWkIoxRoyOk+biCqNuY6X3FZQQBX868jSPeG54OQBVdGf3cd7KE4u48V
CZLflWEO0bL3KPfeFb+K13Bs/qDxma9th7BGOnFzM45Z0gJIzrxZXDyt/SxneH3P
R8xg+15rUSfHx9FtQ91p65eoVtBtiKjZQAzmtc1dHSrOtEcG/IHY2XHRvtxhNH3Q
6InYngTVDk4DgWDQhFOPYsOB+uZQqE2pmFC+P8/ebUjPvaYKlogOOFCdn1+LpTCP
/dOndIfhrYsV9Zt1ZzJGmQkdSCgGzLDQTxEtjSXULmTBXf1OwuCo2FVCb3PfIyOE
0HBZXadjs7UVs4kVvoI30JC+Zn/1r1zMAYxeAiQgPnGhz9U4hdJUc/2sk+oRD+MD
wsgmXZ/2Gnpejly7+zXZwwI7qLH7LKB2k3MRr0d4Gn6DE/k3MaVr45TsEPMCFwtx
ZnrNtn+wibcrtPWCyEU5l5EtN6qdEakEpAzUG97Y3RMoFZS9WBJeveLzZ/VuZVpc
OdA4lIeBRUnaH6JpvU28QTm8WnCxlo0m3BvKwKZL50b41UnNAkmRDlo6O8qFMpmM
JmwE2xrj6Cvkm/FjueFEmRgb3ki5F9xK07dIUQFfidE1uq+CAtXVKuKVDTnTka/C
cCECWT4Z/9T9pB0q+NwLLqmdiZA9SrlxWryUw4pgHXQYvN0LjAeoHMOcTEDD6UcA
sL1jBGG/YOQsGKVmCsO4I2K+c7z6avbiVl4l/mOLwPVGcHpHZ79s2JO2o+R3aFLN
tKVwaITqF0Z9Ei+owCO6sGGJir36VV0PT2d9vvc30Kbqs1DEa6WfSaaEPFjjEjUV
UNb4/ICr7E+JHrdaP0kTc9+EL4e3xsbeh+piktR28btnPPyOugOeI7LTt7zLr2co
beBIVvqhqqVqSo1sZOdIte8VNMtRvphyZ1UDopN5NXLHJVMHUBfv1x3AO7i72F3H
lsLIAdg5a5308YhqnChbtQso54459fVTxjHk5ciZ++aK3mH1eYZirzXjz2NnISm9
00GHEQaqW3bEA7e/jbjE7NLNmxF7G8rAmK3Moe0d8BX46cMyM09DJURhs3X8zI4H
zfl5tAnM7HMN5/Ug+PCyUUeHn4Tt+MPaqeP/qizK6Zk2hED0Slw9vD6IaSe9LX3f
RTkDw+hVTcBfsor7lz9eZ1RVd4XF/sOnqGlX4kSmzpnL7Sk6bZLvgA6MYPmgah6A
IB0tLILS8Sb9dsAcaEWLB7k0qMOBcLtHqoTj9QoPnmDEDjZvJDnOaNucVuaSrtSK
tdPHV5tlc/7x0misZcZOp6j8se3YXtor4UXxsLeajdaaOv7/7dM+wfcQmpuexGsK
c3zINLyduOtFBi6gU1BWG4P/7syy6L5aJ62xtDHBwK5XS8FRvJvCXzFksEWndCBx
PkDh7Ba/4MP0Pi8bOrtteg/6p+4S9YHVmEZYfbEFUilMDcuZiJcySeL82Zo2mQSf
ETWJk+BVVEhYPlFWoGMMYkJe3dZjum5/AJPTS/h1ZhWt8YBjLRN9hXgOb73DgYRR
am9qp6dxdg5azhiyWGO6a99+nWStlsDxU34Pk3p8FlJHuftWtlrfemz6zDa73Hjk
bsCw28Y7MgcG21uIo9FoG+TXjd3GDDh9SDobwBKODvXXZOOQO+lLtqc6SAOjVCG3
2Z2+oOziLG1d9hdbPR0czeHiMRoGenf4SNmlmzkicsQlcUVnk4ubdu+btPO5enrW
ESdq+tKltsZgyTt434YcBqvqtDl/SXvWxnQ1JNdrN6IPAe5oRBBRBvRMY3LCRyPF
waokO2NKqacffyKLHhXVCnZJHGVmIILME7JsUBc8qwXrUeeLZSi8185mjce00PeU
Kyzp3ClavdcqRBbgl3Y1tK4CiVksyOzKiqKCTCEmqIb/OTrF8k/khCqqfBnH5nS8
GA3RDmnVJwBQIe+WFarG2QkaxVKuFFUCHxwZ8y/CY3936SO3Rj+V4oI6ndPNZE8G
P+ScGfqPijpoUcnr61BavyOYvZWC5WUiWCTc/fYldZ62N5XOxDKKQ03FioPcEvUi
/GAMhfD7J8Kt0PY1Oki2wcxu5ohNqyiWR3ecoWwDhIuYU1O6y+29TJan7snKwU8l
kjq7btSrrKl0icei5DM10fKgkcLIsxrNSRuFi6VpQaLSXX3KNHLoh15CslTI6jxN
+mn6/DGupaK0TjFDQ13cx5ecLj++F2m7xT1eyx+szMqzYSkSW4dWwCX3Z8hMV3pg
dWMnXl0Urd9VTEBi3/vEyq60l/ZoQuiGE+uky5gL1bM/NCVx3Xk57Fp/ZQXF2ODv
3Tvhv4EZDe5P+fMLmA1s0FskEwZg+2ustL2uIhuPkmN2ki9qVjQTqYYDAvmmj8VC
P7DijMU8MvU8FGfYZ2vg42xBDMb7Rb0o1G4w3DyjXhC2T7EkDJRbILQj4PLU60gF
NWXrUb5fWUuJN/09zC3MLpHAl6kHrA3PAQNfU8vPv0laH7xatsnIEnsaEWRCqhz7
JFdWuPvKc2claykdgSlhNGzZ/aY46vUMSUHJj8FzXPPD5ccOvp69VjdRLBm4vxIM
LnIbh4TC4XSWMeUgruVp1+0Lp+hRZor6weDvmDP8Rvod+5fZriuYjXjA/aAbjnsK
/7ioEF1CTZ91ElWm6y1hi/DoQRNjVqrRRDDRL1v0xX1dJkeGrjXrcdiBPNkSwiI9
u77X9GfdpejHbvCGs7EO+Noa3A1U/+LgQIAY0TE5/gSmOp5uVQwF3yfQ84UszNwh
Nu4WZ3/KKreSEp/+O8CBIn7CDulgaTxpgEZ++Szfspg09ziAg0rvIL6Qf58uRuew
isdzR2Sw9+U2kzvAwr7is0hdwINRNbJqz2reYoWgef/UP6bkxnOHZQBdHK0jWT9V
/5x68eMZxITGu9d2cSd+HEJXDFMYA4w2kSIdSEHBlASQ429bjl1kwgFgE633gbW2
Mtm1dC+Aj4dfy9cJWcJK9YiBUJYIJYPcWw1McWrkU4bYIEHjoWJP14nXroPK4zsF
9PL9tSyzswLxYFvQJOjjCocytRni6sY5YlAFGHHe+nZkwumikqbkVBmi3+gEwi8K
bbdf4CWOVG7emzrfQ/kjzKKvU/QQMgoTtzVl9gZZQPZR+jGI+Adc6qioBm5fX0ic
HwZ3t7YFTElcKDJDeRkktdqKFfs3M/MfGd5YH+ZSkfnGpS7N8Op2b6EOYheBsdUO
6F6Vg/TCTNy8zUWzRwdEN7l2j1elmjHeZGdS5gr8PEOcfAKTCiPjoCSoUYEsHU7H
U9BplQDEbambXqePU+WMnr238wLVdPFZLCLNJWsIHowMGzJz9CBrPPiQy/EYTVNH
rSlHbNZ4ugCHTuJePqpX9yCFYtsf8IpXf0Tfjs572bv0ifVSLZuGLOdQajir2Tzg
5H4BWHe85wMfxkzquCgH1AQwS+H/UzMj7nmAGN6zdYGaMSBdDdPc0lbk6obcPljO
6gKLLhGzkvjUG8OCzySOxty4VTSK2tbwhQSequxlv5XSUavO5pruZzrMz8E/ryLA
WbEJWAoaY2L2b2eS3Uy05rTJ9dWQDSR+MVib3VjMbODfweUK6TNol9Eq/Jf3EIDD
M40+9uCbIl3YEsTLlcGgEiFmdNaGKAIjh2Vj8jpDSM6DUzRgrpRAuapsGKMPXrlF
CCIrIc5fLOD+dq81v4ey/aQ0vb2zCl+DYh/nIupSUCEp8+kG5v7nAY3y98X/RhZ3
x1G1VEX0CHTVWK/jPwKzhVNrQ4IV0lLiooP5kpLQhLbsNH3g3SirXDaphO0m7M/5
sw6zK3A3kq4yjtHn7sYItvFAIaWgi/FeYR5bE2VcjjDuAQ5uRJQ7BxDzkEyp+z1a
pddR+tf5qwSx4Yu7Rygzf6Splx7LOGz50Dd0L2AHa76Ym1ZPUkxsy8V+12aghnaR
rj3BkHDSuvGCJeNajwJXjwn0aLsz33LDTZsqKDarusLWZDnd2xjfRpNvS+YvrJOM
x0altoxxkZRCEx2qyMwp8coqzAbdUKhcBMv1KKthDijyuU8Rxzbv+031Gax6/Izg
Np+i1d/SY7QxJRH4yXU7OIuZjUCCGnNQklyc6f8hM2adrFeq+Rd85CPPgEcTwDoI
u6j1ie3QaIctMrd7Tzd3bhdY1snO8N06JLpvqkVbIprgdKtKfKKvPWn5QEOdd6bL
rQ+E9a4vTDWrIkWrDr09tYDjYRyNDhl4WNix8TnOOzebndqpUt4MoceNbumDP45N
0+SVX94B437fw7JSHZrTmnc2VGvquReckkGtCrLlxJY58W7d8WWqQPMBk0727vuP
GyUjCZRVZKm3iMhaBaAZ5v28vL4M0nhk7Ay4t/hp7wiOrpWUy4nbWr99CErjRRSn
Y6Iax+8iIrkW+oLf3k/pe18qPzP8rReyZBbnT/BYCBIMd8l4yX9XBKB7ydayeJ/g
JuoV4L0Gm3rz38oVYA3msELuIIH0/zCPGq+ho+RuyMewSdplTLYy+QQRNd+BVLZg
VY4RHHLCit8yt/E1oFL7bU2xNt4vAuyBTcQbwWUE/saX01uBBwBfUSiKN7hJRPMQ
/dLYG4WNQQz8YlNYAfEsSmmFJpYK3uY+V1NBFb6D8Hriy66HRduv4fQCX+DTU80Z
bKWYnxsN82Ve37mBercMcD/07f47KBgExHsl7xr4f7J+gfw4t3ZvuIup0wfuIWVC
M6XO2Sq+ehiOK/+EMJDUGUjlyiKiyMX9nZ7VpNp7hORoHmpK44M9bXqeX98x0INu
wCgwZRAq1JPxD/d2AoY4lSqatEzafyUNSlAL9JExBpA5ImeqeeolIXPZ4+esY+8r
wM22xewR20y8GQ+aabNJKLmfS8IkdhOu1W+NuYiM047vM5M1WiuNfMKrY2CiG7JL
R0q31m+4M9w+0lOYeGKPn2T8NICZRDV/AJvWYV9YpHvbhbhxP3POLlXrPHZYiDIr
YjxCCdGrU+xpFwmv4OwsQLKxb+0J/xDNPSRLtlblzq8eplXgftRonEg3RGcTIadh
bzzUYKvH4Q4bQ6x2kw+mit3q+1g7b3zaCcb7TvIVdqcgK3kQa9WS0SeG8PDO2H/V
NlQwHz1HbFS4P7thQVqrTpPjGb62tzRjNxmrlNGgNKaJZR1YeYaGOolG/sG9xLRt
OvdP6luo+YXdBlaSkYbo1vZwogtn74dSeGMjNjo9xQ8bjBJPDczbFYeVWW+2HAyn
xUxQp61nAkGbFDlvBnk9NKPnHFmms4usYerWpQEb6l9Eqs6rjvZ9c2kD8zGPcCsC
bGO1pfejZg/Q3watlRrzxblHh9lm2VVflZa+3kAb92QFLi6e+0al86oylFsYtG/r
mEMSvYmb/ffA0wAFBHhfKZ7FOE46UGhLo67c+GLQeKDqn14gCQeU/rkJyPiNHLt/
JmZ7ZOB+Cb1D7MHp3Zk+0mdI0FooU/klkvONsyD2eDPEOhl7uS/1bnQmgqvPh3PY
ecyQDnleYsOcNlzhgkOyyagyo5Q81Af8/iX3q1Di6UlZfkPDqHSbwdovGluKNC/p
KPQYealUKW30ODD7esLp4eHj2ngHLoRLYSAgkMfYFBgmvQ0ROcUzJwExqCJruDdD
gJXMr1pm0E2z9pHtD9bugqjH/oAUSqXfq6fcNau5cYHkYw7tKwTQ3uXyUNp3JMyE
bO+VBtCGx2F974xD1IsTyZFdPwu5lauCDiofV/znyQWosNBpcu656PGdBaNHutOF
WL2E+dhqnUffoKmu6sgPW3KwFJeCs3zTxwwJflUzMTaEzkPWHuuKYZ4U2XW9QwrA
jcuLbGyo2PedAYODpCusFUqd3G5B+811Tj6511qykTCbwtRl0lJWVBFK+xyQdDiJ
YrRIHHg1fDaCmNwfqdzF0pINs9RJIK1OqpwrZ+ZHn8nx8OOLRsfIwOj3UyQN8uOX
DiGZflfYrsoetK1MaF79veySNmzMYOZRE+X6Op0YoQSXti4pfuZhoP3O3h5BwwCv
/nO8nJZq5zl+NnO5RJjqd15XPALizHSCPuBWAg/FxzhATrJ3V6IgbrhgoYTr7ENi
OXnfnXXqrbfwMrIhRw05duEkQ4HQ6brjleRTng9LAduIymUeByacY4/Wx1v+dOyl
BqaUM2PTwRij0SPSGrhagjgrjbQQKP/TOWu14a66OihvR1Gr2LXRuMOIZRi/dBQl
Qjybaq1R2CQQnABmkFHNnjHfxTPkUxfrjcYQ6NyYXR5nD7yp8u31NVevP720uYvZ
cULVFrVjS09iQecW37nZNeDLuxnLrSazstXystk2Hx+8VcENXc/4O6J5nIrAc+kb
8SRQsjV3VzVDpnqOkK74zugSnlMMLYVwqnd3BxHVlUyJH90cN5Yl1UCGUHexdkGN
hXKbnVZo594/VAz0b+ovxFEB1X1ASgIt+Dh2bVDUoUibevmFvE4Y+jk42xdSwMfP
T+QhJB3l5CoJibvV5MMcwYY4+IIkATElq0vS9ScL0TztT7qNh0K/rfQlXVH4RaUw
K8qVUzUHh8mBwIQMOLsSyDUWS4xXPXm866SENOUABjQ+EmMRpWsrQEdhGb1DQKQC
GDeLsU+ijO2xAGoDj1IpEu8a/LnKV+Xp6SmdGLiD0N6g8UXZwX13+46Sg7DHIify
n77UFILh6XMIzkaYsLi2PALf68TqR8i46eqxM/CrsLJ62E55Maedo2aspSmF7G3I
jU9/yvVSBSAYVdEK3UD/snPFQoPj2hJ+957WlGuzTrX1pHcnnSzQLKdTq6o08hea
kZWoIv997pS8k0zBf59WoUG14aAVsXnwgtJiTABR3aZg/lANrGaNecfgJK/57g5x
oBXu6PoOgiGpGqNgzqwe/4rurTUYRCRSyPRM9hMbLP6KcRWdf7DCx1FniMAYV2al
WDTZNBvfdcK/iO/MHGcec32xO+mIJpyCKp8mlBhac1Gf8O02E8SXelIzLN6kbEeA
0xiUs+nvPkWDxQ49CMEVvKRZL5dBMiW3/cRvsxFMMNLIT28yLe+qndCkecbbyiPm
hZpf40x8wir6XsLv55jyNQdJl2/1LdzjbiOuo0ymKII3IaYe3i9h9hul2MphD9Tq
l+pOFjN7DtPUlRyq9z3m4U/vj2MX8nv0dQmOewKamw06yoa71bYJ3bRpVfHl+eLW
OIYpQaGhsGwHvtmQRqQ919m8RgFJw1RdFxg8OSfgBqitxYIzgmxStnY4JnKzaiLv
gpKrwtidUYEgMmmCYT69v3KoIStzEcZZGn+9WXRepFKR8jBnmEL+jHApTt0NgARI
WNnY4CbNTZBzrlyyS0EA47TsZoNdQI5OLL6SguXvq6hj0/DdWefW/JfdCf5aQ/Be
1VXOyobrkOM2/XwFxcSamQpiH6F3D5beHdBPBsvL13/kdLzjLtujAnb0QD2f4C1L
usOEL4ysgFElKodUVQVcQ8MXpoUPa/vYxt+r8hM5OiEcX1J+Hdx1EcmJ1y0gfL0X
ZJ+gAtYMR3zFpW7kWMZvgIUqBBguGk4CDIHl8RhbQxoxoNmDKeazfCu7LoC5glmp
OqZ82nJTMnQDvhtaf4cedF8/VIw/sZWMphWOB7fN8aLaNEu8sFgsMog0PhYDaEvp
dWh4QqRzyY6l5vEkLobbOYbbfFaFcNFOLteaj3/Oy0NqjMwRX++EMV9B8sceXzdb
pjgGLZyk0A03VkWlXejMzvSFJf1tJ8qGXnoBjzbaopQ75Rv+Qg7qo5oOM8mJwbw+
nj/2atTA7dD4Q4uVVa/GTP8CP8eZrHqUV2RstEhMXsW8ueV1K7gmuu719mRbY8ai
tSCRNYbipYuuD4pSQk1qOiTcP/3rzup1MkxtQCvDaoOl13T90pXUiZLDZSQCg4xs
s/iqZF93VeCruGhlFA/GpvRIvIVv2pQ3no3k5C9jxNlxFcaZDXaC4PjTF5V8SqkK
ZDOlpTBqFhSDKFLx+0x1SSVaM8aIHgnNjnwmFmOYEkiNngQl6517KlXgc/4HFphA
yLCkMOCFG5Z2XQkE6rULED4hUjc9lqhWeYfRtgylvhUOPBAqMqLzkv/EJB893q+B
z5UU74Ab8TcgqJdInGy5+6SV/JIk7kfTXReUP5OXWjE4SDGbPweyIg4nUdJH7CkH
5I8fLWrO/MiSTpm3g57aEwwtjHT4uP0jWIDsSbfwUg5xRbJjfVDN+XfDYaD30s6k
1xY7xP/j9Rpfh87anXIJsf3w7NsXxvn13+NnBSRd9+H97+npruX5iyxf0A2CJCDx
1BoEM4mzKRlfTFw44M8EmZfJODlsw+/8xWuRkIV8DuSk6Tl8IpW8hz7HVtE9VH32
B1f9L72Rq6qiH8tmDSIBfUi1xRecy7YK0jneT+dj6ZhfnZNtaxtlhUsdMwBiYe/+
kshycJeLQeS0fQLB2HCiKzyu1heLVBztRqi4iOPF0urCMOzbu9oR41aw6o4sq4s1
BR0yGJ0tdyVLL0fHp8kdtryEsGdEcyaqdKLQGl9uX/AjtNIrClx79HI0xwg8jFkx
DyKqOSVLKepJRjfvcgsh6BrOBu67V+JiSWpGCL/ybNPqHveyATvgnIzgzlMRqt3v
Lz2rj2qmBGIXDVdqwPLB1j4jPdHw5RpP3e8xVz+OFiLkBzgwyM7pzVBG/GSnxSdI
PeB06Dla7vItCl98yqRmk/+yhDEtMTSgst73awYzve7ORD1vYwXYFSjFPJTJQXe1
adTnTU38IhNjQJTYz3g/aJNmWDkpcMblhwWLgWisSKscYOdpbAyPuRYmZnBDZil0
e5ZzlpC5XetsQdHrhQZ/Y3H07FE66U1OwVywmEFEGrzFtfq01fgfl5SP5k9LUgL5
avTEUOgODiQJwfqvnkFXEiMLwKgRDS8cfPpACEEqAJ3E2N7a6qehoKo+Nu0FlWUd
MyvT6U9HsrRS+xRplxCutG18D6GM6yWZDzrkknvEKvHp4k/boz59hrnJAzlK9dH4
7JxpXbMnu9qXxZhQJbF4rP1+BxQMwIwdLBV18oqF+6/03TzDdkz7m9g6ASLVpE4S
0tlrdI+2v4eJ7S67Fn2N87wPVxkUABa1T5/lpE2ICcQqrxGiMzVS/HwL0taNSK33
bM8yr2K2t30eZckxrQfsUOe/M5DL+qEudJXxNqwELCdlxqmH5ahWwxnEI6gBZvJY
2UcSd2A8GjnQC6H0itA2dxSW2OXMxr4zHfxiyrhgjDrslIBfFaPUrn8Lhr84dbvY
Fvkponb7jxFrLPi4MJkeJPRFS/0LOX3pJlvBNFbx6KXC1iv50VUpJ6W2xY0qSWsp
SYDUfuxWIssdOu9vet59193hw7LiUXniIcYDqhi972RhXWhRTCX5Z3y+Lj9sWNIx
ocelcJpZy6j1kxwBsfHO1egZok6qEOYpjnbI6pk71jvGBzOy0EgwQmIhlFX+ygm5
BsAXsdEdIjzTi76n5K/d6+k3XzGIYTc2rhMzc1jrtzwlwphjiz1qbLzTXPwIihb8
vBj6fYAkoF6VmUkypMk77zpqj5m9Hg308hOysgwkxGg3hhTEBNLqwr8xxYLaWmze
D7hU2IfBRxNa2iCoHEBnsYmfMB8n7JzkNzB95MA3NRUD0DS1ZLupmGZBMNyFZT/l
NfF4iHLgswO26sHk8Gspbk6hMeyKvkMWc7spteG4L3OKYRm8YF8CyifO8G+szvAc
HvDKKe/ifdHBL4ntdGJ5FhfE9lOhHRSnpiKW0cPaptuYxw1oBR6RllXu3Ke3gLYN
Xv0T3hsC1visUHy21twrK+7FeaBgpDrh9QBD7HWvcRqXEE5y0Q7zhbRDYzfWQ1e9
VlMSdvbNUtl+0YNejHF4f4EBHqWe7niTCZpoCXF1NrBQNtJhztJcaEC72Vfz0Ul1
tyltgu2/d9c1doO83PHGLwW8fdZzRGGykIFTpc3Gfq3qDJb/F7ALRg+Fq0f/vJx7
uIkNCQ1Z2K35453x4uz3ZS7PzgeSeP39i3iZWgDpwh2LcgWZ6NNrh+8GPXI2VOum
/QI4Bj02mYuTe3kFgXoXpmHGZtfvrBO2jyO4uA/lymSQXSC4aq++n+8KDoKWRbBQ
P/EXhslJaiTaoekT+/wD8JMgI2g789EzOXVCTpF0d2/O7TxLAi8980OAD+1HRcS9
VNixO2jO8PvtqvFYcLO2i97ZIbKNxTeEEnbAg+b4eqDJrUDppp+OS7TxezHJJ/Tp
ktNB9Xw4y2P36FY6Go3qf575XjgdKVtHJl4mxus3my/+5LTd73xn2mAYC4nFWv+y
8S8PlY/NWyghudmEwRrT4AZEUZuemLiB0W7kDVgJrYbGkU1B81+Mv8gWOdgI0F7e
t1NhVd4/wR6kBmV1VzQSB3Bc+lYyXcFQ9DKl2XXWlha/VtxbUijlE4aVah+Evtqb
DWrH+JUw4oMZZIpbVYEiiSJOscTwbZf8pA2584KlUKbaWvyoS/5kAjkb6eAPf5Xu
HlAJmqx5UvJTJMsj5vTFyclTHDrcq6JDQmGNbZGnqDyOjb9/qrir/3Hp6KFpaD/J
X9fDvLw1XIWuF+0A78IHuiGloKa/ttHQI5Tea/s5DVw2lUt3H7BylYLHBTk0ptxc
7kgQU7dRE3luHB2pgiFVpGPLjNN1klbVRrqgDwXVzxjYxRnhWkeaV9u/VILn2sCW
FYe2Wn1N9maNg0a/89tuIVUxq5zQgA+HbISo/h247SnMZsP0Mk/DcPG+JYudrCev
w0rqg9ajn3Z3KgPgEXddZQsIfhIeI7NdwW8jlYxc5GkBwKqXmtF33eh+lhi0+sI8
rFeojEPRDO6WUfoC+IOlXxXW51wvlAQ3/CJkZiM6ZMcQ0qEjKcvmae9NOzzfUdx8
vpsaL1Gc8+SxgnYHORXymk92LLGqnUllz5C4n35O98SYAd3jH3DQScEY8HnCDRLm
sKdeDREkWv2iMigW4utmkymOocoK88pcFQ+mEZW/zzDqLuDFrRUjxUZgj4sB2kpi
fqoKzylvFt7PdxRGjLdtYXeSAGQWoDFuFS85baXYyiQKoxP0IpMRoKqLT/vHAS0H
ofMhUrJM55Pf8YhcgVXeaUIjzIgR226M5FcPn6C3L/Bhos8w/k1FplddnpS715nP
1zJKv0mTx5vSBOz9qxhQROx1j08GRktiVLWfRkQGHQHafs5rw39RESL6wlDnklrm
trxHafeQ3+wwOi1ZGQlG3wHh0rtKp2E/R88M/814rrdux1NQvcOdvlnWUjOIA8ny
WsTRG7AgYBMzQ5wAramllc8vtrB2TQORnitC5DCD3dRnyLj7l/P7tzgtkc9k1lPQ
7AovL8QCPz/U2XONY8A6Gp2plbJG3PBhNUAYML0v3irnIvcDLCSOjdmB7cEhwe/F
tMEMPsFMMLBXjzJg6w4t5kt2OyVcNWVYgISc/vVQsUsexrGUtaP2HhEcy5mSQbeR
MOlIpYAmNd/6qmDVT64WaHV9VDdfLXyqwbLg6mMGzyCbtknEfJXz2m8tm6CCZFTr
zYrTtTcQOtyHS09aqunoFVvJ98I4VZjw1yUUnF68v89cH8CcZTPAT+0iGZHd8kMx
wcleUyjkYdt3shK4FpbHMf9T7VQTyhe84s6XjyOR/dvApugB2L7IYF3EqRPq3ZqL
LfT1YAk9K4KNEV2xekhqROQqNTU1F+6HVkILtK3b2NSazQ9SnX8NUVQWF0Gh/Lja
Me+DzdtgxCCVhTso74DiV+8uhypa+abzfK7ND2n+w2T0fi96UwvS2tugE/hswzNd
KWe6R8DGIjaxSbabMjDUZ8AKUTDvGdB/uqy9Vqqbq+IN6xNBOjkLFaVG/c/tegMN
pud3Q1XqzMc1gmvjaXrdQOqEPoWD7KV8B96u0hKXXrHOLdKAr8ygdR9KHj6Kylan
WQp9i0heMz6BjLN0Becfrz1lrTyUCzp2JRWStD7Fawk4Ew031o2mgwg5X4LeI7fd
Ioej4JLSiVo1qq4onxWTFhZuhfzoOP09Ln6RCYgstZAAnj1tyABfvKIy1/J1qjc4
7utrk6EISeUcmn6KoGnnwEF6lJEhmo4DhvXk7FZ8g3GdL8B9sQZd6LR5Frq9VowZ
dR2Gg8m9yvo6wZBPzQ1678aFd1JjcZp56NwgKLQvTlxUybpd66SI2E3f3JO7ekjt
BRfwkldKyzBydSnyeQ9Xzq9DNrw8kHKpQDF+dHxVC8V2LepC95tt4coNNtW8yjdy
J5Jqj1+RuJke4/j76xM76iOquVU1ADpaYNo/pfhkVDntCdtWg7Z9boLlrnQMFq/i
qiLzd+9IJlpdNmlv3OWuXH6KFdI/l9R1tbV+IV1LriRZKWXNFrnV2HyHCexzFHHZ
KPGtHS9YRv/RDCA9+JpR/k7F9jOWymK+A4JthV3T4BnoIvTO1vKgcFUUMvfwkTUY
E53Ve+3bOPcXgjtvb2ieiAuCiYdRbnf5/P9hobJy1vTtyEPSN4JA7rTwl8Kf1z3u
Q5rTOLRzKoW/K/7QCxFO2chsAUDRluGCaVBORz2DhpyclczRE+vQcGus6G8scs6G
VCzz4SsXj3SlSj/8w82q8LoIeHx0q2kS6qT1pkL4sXXJVs02IaiPOztlushXncFv
Qype8I7YHCE2IBcXjCT7c0fNbF0c6iLNx/mrdO6dacPc3fE5gMVyVSrybrfOS6mu
SWXMeM7Tu/okpZaYb0PdTZ/yURRg2lPFLqmdgX7O7oq1wHCKFhctYgY6kbQYPRzi
D7ynEGmDJi2AfeLv716/lZ8sAidi302DAuuU0u2MNp2n6puzcDSIVc4eE/kkKO1F
ZBeK4oKH8YkCmGVuIvDF+G2HCLcEToMj2X/p07YyDkR8uyceC1YhYfvVOr9bpH/W
078USH+JVlNuWHHpZCHIJqfIVszqWHTFvGgo8wHmVTN0LX3dWOKgAr4sc9VBRh80
jZEkMy3g0xhvgwOtvbCBdDXXolc8lJTmHbcwmUA8t3np7Z9hgLdwnK4QzDY/kUQ2
Rrw/hiX2atZlXIsr7BYGSLBXMGFY/p9p9TPwxZh/4M/C33hPDTg7LV0vJlps2OId
Ke15KKJ4DyFG1T4+WP+z3CJUwJdj024wDDQZ0D+v4OlibooLAXv6pKSSa9mHUjEs
eLuPuaaRivQyxLVXG2bGl1lR4lY6gEggclgkqlbMHAcq06ui4ojfCwK67WPRbUeM
aYP5Is4o2WysSCL4V9jtHLF2aPUl9mm2mR5OeBZqFu8kSqDvQrx/mA0TxaQxsn2G
0gOAj0HLMHlX+LSY9QErbj4aApTtCh/wlySB8vZi5KqoTqd0O7KRBS4gsXMw+HPL
xMJhNciAM9/Aw5ozgamrgqZSc2RPGYXkNwkLErD4hl/V/3uMS9ER75icNKzS/rkt
aZHshMAIFn/Q7EpHNbdydGGAZN/KsIcNEeTQU8A8Do/m5M61M3dw4FbHTSn0lAcZ
ph/rVR1M/lc+8Jo1k7EXAZ5SzwtMPzDa944ffdSM92RXUctM5lwMELABKUttvBl1
rLpn5vUze4PA2DH+2JsbIB3I2nit9ivRwuxPoUel69VirsRlN98TLOC1KBrHbVVB
/vRZMXt8TCb6uyl07uKo4bovrAlVwbIesy1iKynnMiNjn2lBwFfaGAXGmI/fWeSW
WSgy+O9fyhSbCI13b7hNG09qWPSTw1WtUMN3OlXYNzrYVAPiPOvRypgzJa1NEl1b
n25jYxcOD6VGnotttg5PNpilVsRiq4e5cx9IPHGLqGM6BMrAf4rWbsywd6/ypHCO
nYp5KFkBs4mSd+3iHwQfGyEPvQZ8zGmSeZxYEzsMBv6H7FQh/QwdNJrNYfffEiVk
9KcZRM2SkNwADT1gn37jlyemKVbCMi4WwkAUx6kbt2gRwvDLjyEaT49q82+vKdFD
DO/CVvS1LRs/2xn3pI5K2+JEA26SwSBRGWyQlRCyeLgtHRaiFPFWRXONdpOGUkK3
uFbIznPKFsW7uFDqp/aJBRyuO4OSYiCSv6LUAn78kIKGOWNCyNA3zUhgZOWOK0rh
oJcyVHBj7lpa76njfAMHfbPwoa0tElBd1tyzhmbO8IRFvB4qKT1ufsarIYYYzeMG
22RGdaUR4yEMHo2bktGl+P+BEzDtKgUe94biM/sP1UO2Juv/K0grHY17QqQqfsNX
xLvvVKG8QaxvjK30Aib62D/TwAHb68BG9cfTDQeajPA4aHXocdfGno4cg6vOPJcs
/gDUOLmxbIRX0vcHttS9RIofh/MzpPqsJyuKsiBxOYZgPwuVDhcTZQYdkfuCd9bM
lHj+BiyzNr6gu0fnHKjSPaXuWmURO4J3UFfwmjOq7X+y9Uz8/3C+SKfpmTIKPnYC
UJWb9b5+filmAnAogmDLh3z15ZjPWOLYp2Qg89a3vCWkWHPLu3rv2onu+ltbYHpC
HKTgqJRiuKtHcUO+xxEF3oAz64+W0xGhEkxWF8h8KgcdnAq0flog/e1aMEet4dFL
Waqe+GwN3p63fUYJ5DKzqh3tccQHuXjDQ2XCQ1zEM+S79JFuaf/vROKu58bn1lGz
eIcIylrJJpmtR9z7Fcij+31/+Uy6AGxvDPLYAKSwI/9wHXWGilCKHVLzFGzz2L3b
qEDF92czWW8ajITqxeJMzAGSpLvUA0fGOEAMSRA/LSSjzOOV7AfEtYSCuXHg7m5i
4xO6QYiwmJrJJg1qglunOcZWif2lTdz2VgciZgHdkDaHQuMo0IZxQZSauqJe5XGH
j6UoLcv7IjtBwVPVt1QKFhz6aLFS7rcpaQd98qm3Tmd0Wex0Y5rmZEMh1z0ayuz9
ueSWbUX6KDPnZ/0mFvl+xZ5OoSaJ3zyoaDQQ7SQ7MXK5BEap4Yqqoj9riOjjM6DK
iAgDoAzPjbana2lx7oXCsZAvSSuu4VNzhmcLkRivR6GcyzYPdkMOYdEgqvjBNeIP
sWjInkoH3mhdXwqKuVmz6K5ywZ9VF0wc8sNhLyv+8TETmZZ2oPWzfeUWKQF354iP
i9a+0XGAuGaKNYX6KI5nifsq51BtN9qSxVHmYtZ4LboDaeDC0VzZuuMLFKTLNCkA
PWWF9l6dhLXkPgPmiYUdy9zEW0i1Gws9lCdGJuNtfl7aZxjyCQwyHHHCDU93cm6b
6YkAls/cGM1XE5OAz1nvMItLR1eCJXVzelM50lUQ7de00Sn0J78iD9kSTHRpsDQ3
GqAtnXWcfzNmE16UL5H/9jLRmxC3D3SQV47FZQSB+mPbji6WbXLRYUhR/eTpgTmm
Iy3bwgDYcx0QwdtXfDQUwaE+6f5rKyNW9vAWfb739erCKZU8EGNkVokGw4I2litm
tqM4uJq3MzGGrhcRKaTmOJLAHmUP0oj0SbkcwFtI9E67h7rlzVloZQH8MHQtApFm
vTUanRy/bz1KuEYjQ47nDP6RAXG0Tk+bMBCLSseB6mffAeVMfeg9hhS97UzeXKKg
1W/c3af/wY2KIxCQisUT16Bfgokbpfz/7kmyLIYRM2UrhJ4LaEFBiBOwurMqn0fS
2BNl+dm6Ouu5UUlbwChk2ssCB0MUQYBBvSpYacLhkwmnHsZUdU1iOHriyK8ga9Wp
bXtcE0icD3CWCNwbqG4QozQIz990GcFi/8vS0tOLv1x0amzDYYxFb1lVcp33wWxR
gxn2yQ2FafKpFW5kqcJOg6+LpMjGM411K7mAhZsh71yq7ueMs+KR1RUTtlzdlKby
qktbLxwd5gS/4Rutddp1uauPV//pDJQzxOnQx1yitiQRYsKwqutMJCGVBrRiJbgb
gkck/HCnkYvhwh2oWH+uw+0Yk6Dq3Ijo2Ez7aNORHLaF44ljG+EUuJCe/Q3VDosp
VU/jVdDPASXEA2XPsncLptm2T8t32CdFjJUBwp8nb81bGvU3gc2UxmTl8NOauVn4
IwngJljHnGICUN+Tc/bG06H6hBjh6QPG3Wb2NFWI7Ad3rMNlNUiQgS5Th7SYL4wx
cUdmTwVTW44EK55gR9ufLTrNW02pKWZ70joUB+MH951DQ+VH6FOopL0QxzfqGs07
L33SGtiXbqYMO8y8H7mTLZmUPbUhZ1ec3wT5TmdJvdRiQ0IJA/jxZCk7vMdbw1Tf
K0Mr9/OjP5QRMfp4fdbX++Q4jTUxGFY0riSzw8QIoXl5MQuPLhbTnfEBuPjEVNp7
6oWS/9fWu5KqoZ+DF/LTu92/fqnFlv4SnUsTVHnJ3FvXVoDk4h+GT9OYAiBjy1su
I6DPpzNlWPugliUAh9NnQUzq4/nfzbM6fTHErZW8NU2CK6tSliEQW6t1WRPIIuB7
CExWJdWFLrolSADH0PewL5BEluH8vcqp9gqEe1rjrdELFImWGDjKCDAPkuQ6N1Or
gunwlL5D103Zy9Y5P6eOtCvMZGhP4uPiL8+GC0ZChxoGWfTN/9AZgqoeqIH9lOCV
y/Ws2k1SLrdZdno0PiYRkW3lYmffn5jJv2FcNidAglv9bm3X41jYnrgbUeuWnC4S
Qk4VLI/RvGmOFfYXCTPmyVzGa2HfqRMwsp31EdQunMIlTETRG8FRI7z3p8k4ndJ2
DoDP1h1TaWWfkgBx+gY3EaCCDfvSb4f9gRU+mitSUp3pixoveG6xUL+zTJV5wz2J
385yKjl+y3GHnbf5fPrygT5Vd7wTHnIyBmzbQU2vmvb63ySX5GxF/HLMihUYrFUx
0FGTZoWVXqGNlj5ZY5h59eCmqI8hE0Z7v/qJSvDHAuKkuMkqVdSPotBNJA1HYQlr
iIUGHmHUELOT78mi7EMgGyMOhIVyfsF/+Vxw3IoCCgS+8MlN6iH/TFkLfAqsTFbL
C55BkhqERbvuCXoQzgUMktmZtXX8/TFjNufqR+HBtYXXdnKjca0aqPnGgpMFFB2i
i4kJRtbJgp4NNC8H6N/W6ircfFYK7DMRV6N+LCKjWmX6mEUACHAnT1jCKCLpNuAo
leD70qhFcAS07DwB0fyD08ICWTI/eW1mM62bU8pEg7m06tj/APfOk1Mm134JrwPL
YW9HH4WZH3nTnAUJba6L6EuZMea7I4ocu6yUTFef6lei68DSIy1UHOBzwY7MeC7x
rCMK3kzq2kD4q/Nzc3No9pjgPAv7aYzJY2iU8QEr49Jr4Yd1dKsvNgxSsWr6DDQk
o/K5DpYv+v/az3aDbIzo2fvPQgYY1mWkR6r1xEDVthnTLDZlAKOxBB6JTd7EEKxS
iJso2KQGjPCgb8gYikJnWbakOuin0llxo/Co4ADFv4nUYxUNX/ZCD+H9PtHfihqh
5EhQ0d0Tb2ktITv4pXsNzU6lgadwPiE/AK8NfOBmY3trNetVIOQloOq2gRKtFvq/
DG0fr26BNzQqdTpDR61IH6EEa2pK833OPWDH6TY408rUOKVV8qiK0N8DlXzQ80Hl
XyGKqwKUPFQhoLKcr7zncUtrokl2V/U5UtgL+8n3hRiIw9aNCbmRpV+Cg/MmJFoT
3H9RFa1f4H8Z0JvDvKMDZAxwUsQsYSeStdC8eCkELW6ZSmberiq1M/LCbQa0bbum
bJ4LNZaQvBH1BHInK8V36boFMtI+nuN4dbiWA7gYdXQERLSTREMo4Z5xCTu22HlG
OsHR68yITIZkv+1TKxw2SD3DFVR4ys/xAk+UKdAgQD0AM0af+HUfRsD8bibGJDf8
qyoXqHFbyzDhJYvWAHXhfHACqUEfQ3Wq5m0T33LCWnDzZ9z32bz8QIxxnY9yve02
SFjFASBe9coffBCSHsEqS9ymLYRJxInxvgtaop14l0FDGmnm3B9IhHwwJkCFCImd
3o32OvnsguFx6D2xxOu6uGespu1BYHjtSopQpJpbwovZME1m/C+Cr46ZqXPbTjFm
2mZARlP58oZsgnCHGCejMLJEuER4w3jc3eBJzYNhTNnk0JYg3ouLb1ETAan4aHVE
w9bLDUl4S4snpsozo1P7bm5UV7JQTcqNgX+Lg7vdiQuWRMIi8PobGWs1yaSea7/w
dsaJcPQomG0s57PvcE2VeYeX80pC7HSeZLmEDcU6Jre1akflN1M7hhQLGDiftW0m
WkwKLNpGLhXlKuCuw6sTl39r68z1iJFqevNAoGY153OaliCjZO6DltJ2Y59WaM/m
JKF0EgPLj3Jea2XIIldphHPhVd5+2jndc3bzI8+4Sn+m9sJfbLNIBOWPCZifjlOn
KUcwRdUspdCT6bh+isyYm8Qp5mAL8kDrGKImIGlxPYhpzjWID2ebABf/eWzJ93i3
gkrEt2t9P8hLBm5OV5FaKaoE7Y8eIuLhpSJLlTsp3QcZzbKsYYq8u61I5FrlOklS
xES32rE0ZWLFZoOIK9qVxkZsJRxhjlp+cMtjaE0sxr1gPj+srVcv+icjH02pQXsk
NBpK8DKZ4ZZNtOgNq8wZoxfgBWEl5mVSsUc2rtTiZ0Tn82jxXlsekr5peMioulCi
AQ3hpRzNjlnybDPg64AkbE4G8iPEVdkTmvo6ZmQqrhNVCWkBTU8nRwD5632TNWAa
tcrZLEXAybT153sx2mDyOYlP89j0GwljRy5VJ4d0PLTDkyW7kr/2vz3/Yty54+YZ
QSEmeTXbk+O219NxzRL/sq6n6qODUbbkLF04SSF6OsfLIo+nd2ME6H1Yr1HTBPkC
+Y9yErpttzRjlY4creWu25xOUQhjyOjggBe8RiH3c0yGicQwMhOa689vv/uzgm0O
FoWti4ZoV2WJhKuMLbz6bgXCpyMcaS0rS1Jt37qXXxauRBFfvKHfs0Zg99cIsBhB
kiTAL/yU/bN5Xx+f5FohKG3JOuxQWeuMZ2KAeOjAILntZxcpLHCMR06KDvk3LWvx
5X9HBp0lduo+MColXZG7w6t0ui5bkeV3fz2/EuskyToBaTxr/l/xe3xAAEHIbfQX
KcSmNSZip8x1xPIz2FbbepB0jb8mIJgHyn5+n9U+U9W6zPNiH8mIAfuWrkvYH9g+
HuQ6CtCRrJoOBKGLvoFrPNw/YIB/8+Gddz8ILSd9sovWnkuXhdgBaJqh4PHZuZU2
PgqGHSJ3nGJH8bVkIK3VXsbSoiSUvCFahtgA6X6wYMEDuu8wepzgEp8Lgb3uEwA/
3LQnEFng48x0GGBs6nEkIfhWAW545mVuIu/3zs3TkQkd+GzUp3d1yGoCERX1631V
pS+w7iiw4GlUqBPmqAcvht6wsrVebuK2DymbzpORPlqqro70fTXbKKOkxNJTiQpN
v+L7xDIIhpj9CeNJB68Vq+CEDlxenZmCbQ4dsnTvb9F0pml+NV1YzVEP6/y6uxgq
JBaJvCPZ3Y3mwB+9BCve2pUtGVcsmyhq410gM3Rk2DMmqOLpNjAV9H6TPo9+nYSg
PckwXLZmn/ksAEIfJnQxYeJEwrj0a+Yp7BZkS50SCmdTwWJJp6Xragck3j54LWdl
7waW9h2jmovn2PuuLfkavqqvlqYOVVbyg+xJ71sbXnh8EQcgFghVKyHVOOutbnMo
bR9C+CLC+0Aw3A4dt8QUVIK9vsyRnKgD/GaKagSBDk3S8oKz83DxjmGlrcwNADmA
4AJPAr7uIL7fWfywOlVmJu415ztwtwgJK4dZWnzZiSM2W/WrbhUFnQ9yZMvFLJf8
P0dF2g4E/DVS7/e0eBKyoeaUkPDwF3tQVgU15eI2wMMa1zTT5YV6eEyq7LX2NId/
/XI7JOcXopqsfe2QlpfaTcN6RcNORpHNM29Ch816AXk67h9gTin2rSVbLkfP02dD
oVRLTdCB2f0M4hyHBH5d30ZviBUKUQIjU4x86AAkA3lNaiqgGIHbdmQhJwJDBjN1
T8zBNhhNWU+wWyRLeUz+D1FQKCyMSqa0RP6RwuPXPBF4vz4PuT1QCuXyRrcWVOzY
xKvGrbn3k7Mo96jgnRUtN9KrM3f234Gs+Igfg7eH2Le/FS0KJB6WpalSvxHz7LJf
nvO17RgMTgGUi77RgRxddUlLM6P7pwshzUr93VHsFGH4g7Y+QTHt/2UelbLt9w8M
mvG1pihzl6vMdHoyp35gg7XYk6zfQaGfDSis0Yr7a0HSKj13i251K1Sq5jf1Kxi0
qxsA4XTcZLbfot3N+V7Wk7H8Pfj8TFZ42Tt06xtLIO2bKgiBEy1Pmfuqxzna2/8i
uvMNtrivpPagMsu3Hj4+hv0Le+LkUFlva5Tv7h+pyC/aooTSEwsfGZB8RZh/mnqk
SqqUXRr4uhlC9/MVp6CAiDzcecaalJ7MTAOtXgPpwGmQN0jZGSpyBbTLAxtjPOGf
HyEx0yRW6NZuxpcUNL2PnYQ4KSK4cW3DUA2hYdvKb16aYIaGILMYbDDlD+L9A6sS
oVEXTcKkCa9AKYw4onFm3Y2t2LMwxI/61iQj9F2mF6x5ADUoFY2NcTuBpNWYgPmY
2kfDjK7TDBgjR17XrF7VdUvn15Mr0kcSWtybxXiio2we69Ow2uVy5mLlQ8HG6ptW
aVdRrP9+KLN64NDlqu+4rBbgXusF4p5WdQbPvo9J5W597Y+BREeVTad3EtMTuwne
mtUUF8NWZXpDvQRN0P1N2LdI/VXHtBu0L3PRMIn+URVpbO11Ix3gVup2344ZMrpG
9c1j+PwzCeQgUPe2PBgO4oYA1Yoz2bvxjZP5GpJHrPLLfhPnuoQhMGzHmmozOyNS
1w/YEELPGW3jZvx+/nfhryGGK4igry2w4FftImcF7lpJJlIMZ4PhnBPU/42cTKor
AsI0zUT/zhSULm/69yCjr+yLVXQ6Lb+opj7DdQHAmeGkTnpohMWNAc3z9d9FbcGE
f4qzif7HWRqJ5RVmR7N9PN6jgWwrmHxXnqJ1KkosJ/wmvYupi5C9OwgTVy0/nJvV
SMrDKAtdT5cDnHJ1NFTVWPp/7bLySENGiuYycu8ftLdtt2bYNVMr/JCBlhxds3Nj
Hqcb8FO3Ci/Q/WU/ePvBMvxmKSpO9Z7WxoQWGefcnc3BG8YEnep3S1g79UnaUIRd
0XEVksUHR9pSyPgObTOATNXE4hhIkif9BLU8Nn6cLKqjpQhc1cnwTNihdCzO7Nmq
Ol8T3ycgbhAMaH9LF96Kxbs9icyh9e0I0jQJowXDF7Z8g2RscEfUo/YFPl0vFHu3
fkONtIUFB30F2WXPZfaq1YXGnb9aKc0DbX4wvwlgFjQ+0TEfW+zWUGTU9Mx69LBq
swoTZlQLsRK1yUef5dTXfbV1VwWW/GDCpw/R+zRj1tx7mYQ60T4Yl5zGDPikigkK
KNGNXZBfiAlpmA1d4wfFJGnRFf1fEQyQfR9tI8BTYX9TIRpMihhG7+jKrJl8+HL3
YXBv1wBmgSJ6blVzucQ+50tP63sLMA3IfHglp1jeFJbrGWUeFdAuPjrH6udn6tpY
mjDWW2ibVR2N0LSbWda5+3l2QfryEqx/8Wkm6YB+53MfHakrZS3kiz5hU1BRjTEw
uvhvxrfn11A3lv5a4pYTqN8S5TDt/SKDOR70AoLlZokixxLY848+snQVCkJyH9pz
IdIZEWMA8WhvViFSqy/e4tWHLGXU+sOtfnEb9Yi+42B0LnJfzsKJ790BGyVQ1aDX
F/3NEp/zkJ4TkQH5dfSTb3TmN6ryDfJzoNYauO/yoqPc9P6O4lbersZ955wAHekM
5hqjUQct28WKJBRtPvxfgppu85L0DAWd5YhYwNlbEGLoIp0FCEjEDLAgfDFkohiQ
yt/hpc1PeMS0R0rz2TdyrXtyyZGOUlXlp4bQskyKhi2lfG/fiWXwO1gDRKRcbZSs
UE78D6E6070klvl4V6bVys8XiK16QM76rIGHXfCHh6wjmNdwtGijf7bal5czWg/J
lr6ITY3gfdSBa7sim0K38D5KM63aq8VUkNTxpUXnxorP1P4q6xl0/DxAsbdLoKNh
tAmmUWslnBI8tLDInTwN5F3S8zwe6FS2kA/QmFe0J25TRdJeUdrB+ho1H85RS1wr
L1gF0GNTZvfsdl8ZoFptVh3Q6gtH/e2M8A6WJjdf0g0UOAojhLTpLFbrK7hn9wzT
DO0h5o8/VoB24T8QvfVVilWZtbQ45Rjes30B7gctJhmUIwXU+Zn6duoyeEOjElHT
VewgYkx0zEfi5wil4RVkV5gjQLcbxahSnR/oYzfCiOpHw6NvsDozheV3/hvK2C38
iZ0ClL4lRHI9flUmAcWJhbrmPxBqqnmAp6EQmn+z6eL1KYMihJsVGk/3LKuQrPbV
fGNbFPYXN/ybGL3DlA9TB4DRLk6GcocFvwdEv3ejTVGiJ3osxuLO7lcM5SCIFm8T
oJ00tMRe7Q7Ec5FsM/r8r3EBhxJYY6A65pcaR31E16c1klOy+nVyVc5v2U3BA7vM
5vN9kPINCFqXs6bp6+dJ+O6/rgMGEE359tWOJuRXBUzTnxtn+lnoLbyJnO2HML80
u1jSZOSkhIRfaFotCfSSrnXadnuVe80LVHB9QXNl12lSuSRn/rWrPIwxFSAW2N2L
TY3niOuwUwKuZ1xLGT8jAlpjdc3WLvRyQW/KV77AFQe8iEAQYvkF9Xbp34dhvXFx
JZAkM7xKq6Fq/GM5tMMQjV+VMTBYeOl2skPNxjXX0V0qmrpb1lyJ0s3dbiDJ+dXc
XcbBX1locHbM3VNVAfTYv0H+VneW33u5gb9hYafeqWupo1d/uLmy1VlfOG6b5p3H
F/32zVAb7o3/JT2TnimX+Wk22eTw40p69w0yjagfTs2Hs6AE/53T/F5sJjqMGjIq
zWzw+BAragMDjlVQr1SRDPICUpIDiKLSJ7jhKjufgagEPIfs6VYlpukGQUwtnyEN
5G+hixSjq5cY1TF7QHx2rLNgfejepHkIS++WHBzSXQkCEdIFYRZvz4FhMsD2pHH0
OnyuBicdqtkIZoXqx/m/4EQYO+BwLoRykX166AN9ssqByKDu263hspM0dq6yA1Uw
/7YpdJVkruhpHdPBdEyX/BUJBpUBhTFCkbZtOTy0k8O5rHZ6kiE6hm7Mo3UaxfXs
+7KO/1PssAMP94EbjeU5M0oZDzzw0vjKQmnWAQfqFH5KIeo6d9vbOi34CkIYDi6t
KYR2UqMO24X6p3ToTwqOzgTb1t6GzMAam7LtEfYcn9BBdtBg+4fuG5x4KqvH8CTZ
J4V9uzmhuLVgW0P1b6PoM5GCu0NsauZ6xlFDRWLE1iZAfDl+2TQoRgidVddRal9p
K5rNWswwGbxO8yIW1NFaq0+qVwFGiwbWLPbgFyMEk89tCZAiduKaAVSvphk5hmsx
rs1lDvQt29OTlbpHEc4yGOwbwZsumzjNDZ4iFcDNEpVh2Q9Nq6eG3vpeAXsTbq5W
d/bV8GhLInWxtMmi2Yub6A+bvL0/Tyms2Hd3WWgRmhlaTamwQl+t2VtwDaOm82Vn
9A0zt/sltxjfAyFGalFh0oItbdPHKhkgVQITroDEudke2YopKtPxGBMkL6POQnFv
oMO2Q4yIWt7dway1+vGTIFYgl/u31deTFma5Q2Qz5urJZQ8hEOLQ3tnZ7YX9RVKo
x6PsmgOdgEXonsxltmFwV2izQqSzyb7CGVxHWw04N857CSWFtqb/tN7ZOffXcLzT
C55eeQMZeC9bxWSt7hAGVFAJ+n/+dg+x3IOZmF3qUd2l/QZITIqF8bKpoks0amBR
dxynmZdWBhhQlhR9W5FXZy8kC5hZKWc40K7zAjKkCugPpAWXk6JKmFBAzecm8Tnt
zYol1NhrzhWv9Apxj/n5wsPTAR9wyhMfyf/bji0x1ZnCZ89X+EpsgmksFeGvsF+t
xlpSGzP7eWFGZcgl5DYuUrZVfaDZuiWVEuNPzsNK4cyulA1nGSeb/jM/LTqRSxXX
RNZgzWvvI+qgP6fSNsrNtf8ROxy6x/fLc9S+SwgIGc3OKk8w8ddnEdkbl3ggv9TP
Ib238u66I3DI4u0WbipH9MzXn4U/8GF7uJj9NkvtQw4tU3zIHpjTG9C7yAhShNoC
eTOO5kIHY0P3ydrky/q82/fa6JfS9ha+d4EaGPJ+1n3TTyZgoSgr/egQMsMTC9vz
X+R8uv/ELE4vucqvtF3XSs3VWb3lYZ3RM+If79tpjeO9RJ0glwncBXFdzDe43bvL
i958w/Eio2GZTUzyCSkzGP8gQBTvnF/lqwVtCG7SRVKtsSw5xG5RAKRmK4A5X+cC
JBGWqrXMAYntGxFLOs+O3n3diMIU7inb/qr8md+PcR6f5VM7SL1ESH2cGmyXaAB5
9UXX7Qh/1OZU+kjHcK59IyCgEjKsNL6ZShIseBXrxfAUG8i8RqFBeIcuKDfRwEmX
HT/aii4Kim8miWc8h4VmvDQkxGnt+yUNdIvR/ewq5RaTVgU7I42jaD3u7gxxOS/H
x6Y42+fnHIfsnkP0I684M7txOSXdlKMEROj9mf6r8oRCQjNs7s3b4GVh/rl/mZOR
krlQTo13DBDjNScF2jc8GyW06TFWovgrndKYWsjvIIzxaC2iTCkl2C3hklq/VJPS
hXBdBDDTjKyiCpy1V3ql/eXDQO21zWMjWXE6o3w3g+J80rTP62/0bL2etPj8L8qf
b2RFoLicKsX2698bhQ74ib4yL4OYLl25FgMXOmb4CTR3MSLxT2sWFPIM4zsPzwU5
JXsaSY3gAunqrfR1u/h2VQIDXMAHQElN5jxrCmqTGmxj5Z5pyNXwQJXy8IUrH6P0
+MCXg8ov93ZBW78QFzbzPp8ILLhM3oA5RzwYtV5m2v3H1pwUdJ5nwrZSzAr0yVgm
q/N5G6ToJV4okWSDlyEJsppKROs8g4M4WWuImPKPGwsVr1hpkVIWPMtrrixlRrnK
s0QxiZmC69/bTE0QlZgj1oBPD7sN28tghP55F9Ipk9niP6BT2Sox5pjd50+vcypx
9KLa6/JU5fRZV/XbpVD7XC/u4iwmIvUoRpsl9tOYh5+UfRUkmIg+tJqJ+wdXmNSj
UGg3pfejH0zWXXugWH6gjdTFCc9prAxb4S0h6mgkScbwywITzIS2iN1lLfaClnSs
1tSagCyu76mjPml3rWotSg4zBrCRoCSsyT2adf/WsP9wLc9oKmNCw0FzDNjDY7Hs
FBmSsxJ8Ur0G24PDz2JdMlA26y7nHJk1Cro48J24KjVjO8HYeSPxEmL/lnt0NosM
FjIhON9Bmx11BFzhlBDxD4IvHX7NXWU4cF64hchOSj8OnnFOWuXDwVYyddFrjqWo
7ADd+jKKQe59LZRdvJhq+qxrwCX2zQCzFU/vvara74vezJn/2prBDIbKmFq+JLZK
PdWcnGxNNMa1oXpeOI1KpUY5W9kZ02L5GyDEHoX84lEfejL1DCJLiuBxlmWjSmZF
asPEe3V3s8HbEcERg9CGza9WQUSmgGKBfZM6W4UvdtUt3OlV5VGYa8YPFwaSKXII
BWGnA9dFbpCphE3/MUlWxlyhpgAugucWf4KjTm2JdByVjKcIgyETLIXLpRRQ6LW3
RFvd8acMHzcpmmeyIrDaJrjKZIqDq3MKJhefpgviiNabk0py7X8zE6U9jreAGybO
rp2KgBMnAxY+a7dnsA1EaJWPVPnPPGitZrlw8bkXQ6DDmOYslC5dP0hwTHPstMML
FWyWFulAtBV8Nsr9lb8nzfqphCytJ+6ldYfa6zkov4FaSYMs81L2u+81cuAeDA6p
YTs4hlp/rdwrjS1VN5Uuaxc23TVwJktmtATm5ljLPbxewZZE0yKsHnCyQ2xnjkvr
W1+O5nWE4Bi0NVSCpXvhK0lM1S++8zYq8IgIYLvOc8mVxhhggeYxy0Qh9Skr0r3+
tCL7ik2b8LU3PDXJbEFboQB0kMToBWuPUdExi2UgjlzukyKt2WiFuP03qZ1qa86M
yk4v5c339N1wpVh1YDkVwxUyshlQ11Ow4rcbiDtrWa9c7WJjqmwhm3KvBuEAZMlV
s8Axn7pNhOXK32YGAsOhIfueDVZgpQ4nirKE8rG12BWNr6G53D/hg0d60DGzX8t6
RtXomSHvYoaKsGpwPP9eHC8JRkO7YU0wOhy8kGFaOLxiumLlPh6qGR1e5oAz2Snx
46rMPr5ccjJx5KbvlKsNzVGMHZq/mReRDFehreCXgjhH4IHbEzsyxp/y6q6HHDtp
fgwsKf9XxIDfhzWHdVaQCZlgr35VeIeDHdWbgvYBd/3PwfMwbM/wrPJNT9UDnoFp
rOfGKJxWmQvz51SJFEUlI3EYLDjJkH852yTExY1kl1lbag9R10o0maSOr+Sl9Jfg
P6YU8oTKQ8xJYd1jpN5CFTrCCfQRRcJJjHjjuMvFZ1f5ICjsdEww+AqJ43QP6iA7
Ajoe4lt1Z+r9xH2TnXBE3MGD2s8ugEb94/6zp8deQntUr8v2oGfcE4PVGPMf5272
pLJcTN/M8IoN0UeOE16m5+GDn8L0xwG4WjVlGQNrRSA132OK1YIAr08VbC+N2zsX
KPeq7udPMTWT8MH0+dLkHOui4adPkRO2Tz4ZzNx1s8mblTf7++XlptYhSwQFSLP6
eTTh6Fwr20c6fkT0Qr5vNC0mcFmI6arrdblc4AZD9N1wy752LU7+XN2ulTD05iHy
4RzkqKjOypFAuGWLcqkSfEpmdJnNXVqZVKNSqEOnwIhjcVwdPKSK3pcFxJ/hDEWq
ZECTGIm8vCPVD5uKRQTYzQEM25HGvq4VxRZX248jl1P3AVafj4MNV5YCajMQauLQ
oS+a/Ip+AePEvkXZoMZbO8R8nbjTtlWF3hEr0x1bzCoIYM7zHFGrfVzlggFa0ZXX
hw9sVmhhol8bHcmpv/v1XuAtqzK5qv9UWVrTpJ2NX4ZTc9gVPufLOUuhv30AMVMM
4FWMeJVirDUFZTVkvV6AzhxNsDMftEKZc6nn0ez+Em87PWNJYaIallB6BMTEdFYx
HyhW/uwCd8VnGdjjCQP1h8ckNBvHYw1cyNbh1rpWv0FoN1Pc8lM/wIzppCGroGbA
yfp72b1Xa6aP+7PqRdaOFm5ZjKw9Pm00WbuDyoJBJ3oMG9xY2zOYjrfJZJo3PKKQ
s81c7dqFthhVRpBRj8uBkKQDW2KmbkUKbOKSRgewY2ioGu8F6Q/LO7R7fco1YafK
QzeoTqILeIlrvA1pn2aNTDrvoNzcqHfCIyGTrzH85xFI/51DnThkfTKnmsvETNE+
MsWfY02Y/P0o5rYduKkzIFZ+YprM5S86RQd5Cx3f4dVqnNpO30C+XVT4wl4zaApx
qa16uXPC9x+/6gYGq3yJ46WTLgQI+R1jCrwXiXsF6ENnJTWGBZH4VUvBSxaLoxvL
h/+PiJr/Pxfa/TM93c7sJvqfO8H3a9y6oAXfkyr3ZrrlVgL6lUCWYvf4YzQ3GqgX
C2ryNlA6iylgrOQ3LBmXZrLlUPsXcILZKUjN4q1RNQMX77FUFX6X8g7RGy7gtJpq
LCji5M0ozx1rz4r/F5wzFfWp71dQ/hpuJmh8M4VzNJk7HYCzHhirvQEw8XiGtAYL
veR1t+jOSuOtRdAVxt0mND/wWUuQucMnt/Lc8jrOe3K9ui+dkL/bcafu4JcxRd8T
RCGt5tGdoZ2WoRO11D2MSOP7qk0EoGRumNLMfvmDkmXRxXVHIVL9iA4WGM9PC2lM
Rb6R4Qs+oi4Ev/HXqpOnrHRATzTw6mB9acwGWZRDYMSkpDz1LQfsy0qK9bamSKHW
4MRAd7pRI31MtspPF1Iqb86XSH2jotsQ3B8sQpH4hBLJZhBBip7jzLBesRfU3SFS
btVTZ0iq92KML1Jfh/jdAP9JVqg8ut9oF9qdxchqOgiJTez5v3B2zR2mk0EF66hX
vyAC+D5mCrPtdnH/FgeazVwtCm+im/TxahhKWWi8QPZrrTfV4sLTWnKZ40NlFBeQ
boB53xc7y0Rp/NzUZQQSRRX+Ykz5F2VdFvjvVzNVntRhwptHh1kUnGO0tqPMFwdq
ceT9rhd1iPXV19MH6KOm8v341QA70cvh8e/5cydP+y8Fpxi4e2xbBcgo6cDvFovO
xmpXdetTFxWE9J2se/SD7powx8zeHCoeRpSzFr2FjKOixYdNmXNWq4Y2CwQpb50J
BWv+Ll67KMd4jeQX3BJ7/KIHTfdhIgxor0gQuPj3Z5lTu90re+nJtozAROCck+lY
C2zNFenuramBKQAB9eMaARCAuac5fa5wxupEPBVLd282sPBkyq3PQT7TEW+5lF+C
v8b5AG12E8hb990RuD8RPGWHDAtVMdCufHXHAXfTNBMkWJpDRcqt9NSN+amUHp4L
aQpvjbIX7OHR+w6cIVIzUXdYMtma8cNMmf/4Xc34t14qwJgzhMsXFAJ2OgMcZtJL
xACr/GmnDv6qI6PtW12cX0PlAenuqAdGcZhsLEaKSO6KtMc9dpi+8Lu0SkpPyZxA
WKo9K6NNmB/3KMHMaiOyv72yR3LynimJNsDIrkq4BzmFFIBGima3+jUUUG4HoxCK
aYf1Z8+5Xe0R9tJ0yYTC4S2BvJ9IpnZWhgf80/Xf4ibnzQ647g2+lR0dYqEaGPVR
YRhep9BXk0+t6khJ1VsQng92whrNt0bNjI8JKTe4Hbdi95tvbynoh1uupDr6xWeC
XNj/vUuw53wW0tUTARA8riVhkyqxYZxSdm/WpMkV3DAPTUcSYrxkzkWCkv2VbaWK
woLnRW2BPc/DGZKRKlh0GGqTpaL0+eEro3eGlzocEYUJ44ej5CUq/G+JJHPmubSW
A3uXPz8i86ne7iT1yQInfzFglYOUro9FqqbJPmfhj16gBs85oIa2A9IcP+W7chge
g12iw4sajB96sERG9Sz5na0JzDwDjOx5zfmJqbiPnSzR3p0yqptA/L1yNE1Hg3pI
m6RJD/Xb61w1C/kyVyjusTn9JG63kaCBIfd8ATz+YtlizeSA/8zVjoVnR8UVHhdL
GAy9onGjLqk2N8YnbxjCMe2K04KA1q3F5EUucHQKq95Xodw3I/PUHIg7xb3b9aOg
h+/sxYfHhFQh3U8OgM6XFRSGtQaDF0FrvB7T/MQxWB97bfU1PzpYLOwcjtzLEttM
Du5cz2RJ8mH+vl7AeaXAsRq7OfkBLsyoECaQvJRKPTJ0uuVJNHlWmjUkUueWmHOj
coeuiG4xS/8AKDy+UsJJGiWHbskOYgoeVtlWrtJed87dgTnpPpxrmI9dxvEQD2SF
W+Fwd8J+c/J3JPPAAqxeegT2qnEmUDJta43KEm5fxlD/c1fwrH0K/EKBeL8xjex7
P/f+25IdpgO4JYCzAyBipUhP8ASjRG9De0EYmR1esl9e7WjFINcym+m/8iYnO+BY
ndp6fWJbN/avOXCDkP2b8fio10jVbcD/fV/o3btBcsD9odf0IzSTEeTu58F7KVu2
pk5zr/Cq5WOegh9hK7DOTsTwPSZY6dQEsdADr9pU+1wLVhNz78sEu/Snx+pgxUlH
oZ4TFcJmqAKBUBB1GRUC7hrQ5K2wguVo/HZ2whSuprLdAFd1mSNhgQSvSH8aQsh/
kV8uwgXhX9kPztH30nTN91XeN4u8ePl2Bn3Lf0ablSciLq2rEV6qGCl+8tjesmOp
4Qenm1uNaMmtyfc7E4QowD09dD+yxpt87er7IX4Xq2zuExPW2vyRPZ+PXpaUYEh0
VX0tZI5FFNlZWWBaEuSgczSQIcv24imajxQuGTU61IKUMQHXjVGtaZP0cC/NHVzZ
2WQ2rJeAw2tpJ1aiXZKfEo6eWumRCLFPcKW36rmNGJ1yhBNvdpnYfiGxP61/lJme
d+L21en+tNqUpQfJgcNZPoJr3ObI1Layzcn8mcAkfJQPmHcoAim3jMYQb/m1cJrn
M5LplUhhtd+TnoMi0yp9FPDPUYA8tvOr+OZwB6BqiNUvz/0SYmm6p//+2vwkdG7n
sE7uWH2TdeDtXhQmRa/Jq2/safiyXV3W7QzZYAmPhb3rZqoFGA5iwNxGwt//VZ9K
xrc3+a1TbPkKSJxFgyrVoaITghyg2lqZxPMpnikH/5iM+yrTmEDTevrfp2bCR/tz
zuIKfuVBmGiXxHzvCq5mUGBH8+E7m8Yd/h4pePyWh6Unv46RYUIug0PgwbOHDtKS
24caVAaf8aD+9Or/WYP/rutDrrcuzds+vjPzj/x50FG7K2qNCiY2f7/XeF0K14os
ZJlcgD7QIWujxy4Q1XKvQSPcsqKoNacNa0gcmNdsqYBu3bhpT3sGDxiNGFb18jEn
RB8PAGO+YMZfuwVfnkRppFQuDETHBmiG2uR0VJFA4BNdTgs0miEvVN1XrFJzIyZd
cEtohEEnmetzPbdPmS+RDhv4QJSHziLq2Dws+/2b5rT8CWzcNrymim4FWRqc+1p+
2ecNSCo2G2Dw1E2SGQEhhj6joQMmSOxEBjlaR8LOKRZu85jIhPGSPOvrkctjA1DP
e/5ffZaMXwFL65t8StpLtmHJvwIJl4bqzZcXgYKtd3h0cuQRCpKAAgY4/TICVJTg
5k3qpZmV0R8qQNqTdiP+GWS0epsiiRJnKhf0MaWtXY1QmLlX3l18APBkZuZQynar
dTXqZz99hbSv7OdK5mKt+2evQuOkX5fHheXcl1xtv9qqBX1/ZXQlAS94FnkwPUYQ
67oPJCtKaZ0d315/iadAFwVRIBG9fIFSpf9H4DVI8ka8GFYgq/rUGuqcObC8HOa4
HU4ECAkJ+Gh1oplHeGhOiFcQBJIR8gNMV1J4o47YIb+91oKOCIoAvyV7eSFz4DwX
xnShYoGJXAs8WlYG/LULgCNa91mWusghHzywDNkcx+4cQ/dafkyE2HTGu68eK5Tb
G6aMVr+VnsmxEhOoWXjZU+nUz1v5lV/a5La+3AzOD4MqsEE7Joq8r9VFYRzkFnD/
9Sk51PsUbZqPt8B2c/7YlGPeJmQgi2L44/QB1nld6pDxxgsTlZMChKQ5V+U0Vpxm
wPHaNFpugHMxPSg3ddejmUaPMCF4eIOvm74JipUCM9iGu8zz4Hm5FbbMiHlVuL/v
zF2CXsLwjr5SZB+fFSltyiocp5WDvQYEbW9gc/bkRFL51zzR8GPSc7gjmBmz8Ldl
tuWwLTSi33wH99cXXznaA+xy7JybDOTsKM6EN0IHGIqoRkIahNyp4S8HFRvu+rCY
kqcnq5EqfhHshtLUoQdOJLOsXoFVOPMDP7R3Df5+ruX7r7jPksEnV4KUPqnJSovh
rmldSb7tshfhnLUrjecLHTASH0VcwbskQIseVFWvqIq2uZTwWB4cZTUf/gpkhuea
LxnIKMRP6i3JALGgWeWHXdkf57LyFfO46dh+wDyAkmJF/3Go76LTxPs8XHWDzZuH
vYU0G04y1ojVIIi7dmrzzEf1wdElAVKYh48vKk1OOu1qU1n6E/rzzb4Ay37M3q8q
aE0QAqjN3qHWKvryZ4ANlbrZYTmS2OJ1eCEh0UuUXG53PXS/JTdXNwVneUARYUwL
5JfIddpXcmYDSe1JbWNYsAgGGo8Y6FXh8Hd9MbVkJSrAm1T4oKIM6EJHyyMJ01IN
lG4/bVZAiR5OLlJKKrD1kCpyOGETTnnmv/fpoYqZ5hf8G4siAPaOXtY32From7lT
1z3fU6NUbKi8/hm/FQr/294iklAu4vDonWJYgwKshQ35IwjsVC6vuaax/BgD1ZJc
S5KfDbEcRC7vn+uCiLqNm+M3RpbEmVklc+D1LOoEtJjUaefWniCxzH/EjPdlgsRR
C7wC8CUIVpuS5IT7zcArtoOwbplHrDwkcP9VaKqE4Ib/LDDE9uSXhsEe30CXn2wL
zaOLAzeqqrfmWbQHpDTFFK+R/FCgg4ug+p/o8YsxVdCv8esGHSX2+jV8VQNyAI/H
3zJgGmiUkvs9vPGerCJVoBUK7eq+8tOxBvmYMGB0vJO0FpkCusZ4hTdQlNWHVdmT
XOShk+4kFQLhMuISrqYxNp4/pnvyRP7F8Hxb7lAa4ZfHpFQ5hVzVL+z9G4yIMA7+
+CDNMbGzxjN2QKCLzTTkucnXRub4q4+5JGbvTVFzxT99DovxthbznVh93xtdggGt
NNOCNYM15mGFS2RWCGV8HoDN0a2M5P5UC81DlRs1VtXSYBknAj1qRn3MuQSdxSWG
XRxpEm7WT/lnyjDCQCVdJFdHQOfB4cvJTVBAhMvbkK1yMI4Rrew2yODKu1sS9Gaa
vqfNWJWPIc4zIRYU97NygDuRc+dYnEKKZv36Pyt8mfXDh2lBqwWJv4BmWy+FTBYr
o3JxS3qiDKMIagx2ZMOSTWheMrMvktqMNzPN3BXOBzBsmMvPba3QHhFM+iOeBZSP
d9BoaTXxN51R7qCSXtbY1CI0i3QtqmD6qwz7W+HSFUzyqywHb8sXCLSVBiheQcs0
gKVq80rdDyXZrs7fFl7wQVMdaPykJhnB7/qUBf8FkvjwwZl1+GH/C40pUHySSac2
IKjH2ZHB5zyxXjmoqJ8wqJOJLdtKelTL5AgODUeEqxqtT58VrjEewkOeQ6sUTE8W
1EIVonF5kkrgqI3fBTiiVKx/gc5QklZn+pK0OsT6SHA6Wi2+BAz/LhQrLHgMOdL8
3QtQQ1JUzteVsns35Rl97sAyF/Rg90ZTXocWHeEgI9VSlUsHRiWO2m631ri6Dk/q
mADj271jVgEzcijlFYxntrXxAH8nzwcGi6GV2R7VxCxK0CutlaXgD5bun3W6JeLI
IWS8x+7dRXI5FqtDk6U7V4BkcFLBaL40bfbSdnI3+VSLZKyjESHnDrlpZmQmIC/9
V4I/Q73Rb3q0g/OFyM0Y+0wz8lD0/+UZcgdnj9y5ZQvmNWrlAgCIleb759OrBY8H
h+Sy0qDbZ5BQysi/rwZzrMQETyppQeOos+Y0+jIKKlfdCz8FUhWIcwYq8K3C+IgJ
pbGVwElbdGbVSOv9xxI2rGsbG7D+SSeBvHDUL7+dC2/BwmRALVMWIuzonVxHlyxE
IbpVOF37ts8KiMzC4OIwmuQ/gPhVN1btIn+c8m7eEx1ewNQ4nhhNlrXSp0/IcBkQ
gJysFMiNOFUJXGlAqXf3bjJmafCTmsX+6U5eSIh8h4u7FX4SKboDS0LPKvQhmlYr
RRcfW+kFg4fD4c2E5w9Rbvwvx/0fVewp53+/qBHQBAB3rK5Ackcrilp3oV/nCaLs
AU14/IupbfsvKpyCeDOY6vKPo1AyXkBgjEtAYNrwSHzjVQIlaQ7fAWWDZl6jSWty
gH7ZSDcB3cODOSzuOzRbMm+/Qo9lKC5ssSU47Cmcp70a83mOK8i8T5QmNCC5KokL
0V8CzqOfGYr5h6FGQK2GcO+Fi0IE8Q67nztG2FqzfVIRP2jImLbOvTksWfrPKDlD
2cxqiwCmePJV3qm0unGIq7qGGcQdzGKeE6jUvsX+dkNxOW5RrmvOpsx7hiq3DGN1
n4SnXRjnEjil4XB7aGVd0DXhhJ2n3sJtbzfWDCKqSNIhRgaVOuW71AvfEnZmymwR
/dq5/mzzbh22zJRAqfNlIM6+dGxvHuxpXl0TtKBQJO1ehTRBTmutnYHHm9Yr03NN
zTApCQ94a/0vfcveyaQStP6tEV7Slf3GewcG6VM2eE1cM15/2tCYPWE0w7orc/MP
PQALk2VIETAqeksJ8Pq6uWT40bxhe/jpNIF07DPeFHP8mQX8vh0qRmrVPzsfi5/4
lprICn5c5cIPeOyrdtK9hr/pAYNzxAd9n6QRs/zPQyzzSaBe/1C84XjuhxLPbgCk
q4L3elsnQH6C786rVocta3HL0J4d6DQtBZzETazfAT8O/Ydksb01U21ps4tjzGFe
/GsWkgFROzPqGaS1Aoq31kEaSPnyjldFQvrPonVc63vjpstE5/haJtD6B5Eeeien
JzD7DFoQ5zXWXYUREBo+sQSG6t7KrlctExiCJYB9SBwR0o7YSbv+mjqBJ+p4WZcr
S3Pn4OcwNKiOAc1xFv+VozsuxS+09ao97EsvaWs3CJgn6O2dvtl5GIEfEmRukrHH
IZxD7LwEsdpMCwMO6o6uHm4UkAOnx0YQeAKHXLsPzVq7qz2PBygoQen9YgL096+F
RjQNygYS43u9L10+U8vWath/vheRpEbzYmQuCbUvIjnp/GZOQ52IfrDbFMSlzqOo
ar43ACF4rOoDSmWozCOBv8giNZ1tdTkZFSoCLceSiXnJApD2Bz71gZZFab9ksfWu
EDlVLzuOvXhvoyOCeK3NIvfmiFjzQ45Wb8bA0DLLi2iiBn94qODoO9FXpKijKxUB
Q2ZeHbG4MAQzfxVNQBg6K+L/YfoiKBs0+IpJqy1E6qGTKUlqrs+aw3FMMCr5jxKh
jhgc2OmQ/bgZYSSPF4LT6Cw8GpOKvB213O9J4IXBy2tWESXsLt/8NRZQdEmfysiR
PuVuS07BUpJ1AuX3rhW3PxJ816bylFHt4wTfXbZ0da8Vky3I9AVbqNvnMgoY9bq6
2opMGRVVRmdc3jfePDYJr6fiyQBQ8MJqEMGLZR1Gj28by48brt1XTmwHujDsgT83
1RqxShdcuHzU5QzjIJ5HQv+8K8j3mBFjvXskCK0xkqorx3/k2ukLRbFDMkv4pGrO
LYBD7rP2E9CYX0QI7tFJBosmGhcG/rPl6wLxi4Q9jaYNSxHc8LAcA7H8+5qTg2vg
Qbd3j6K1txtBpyHqwVjd5pSiMSgr6oITnD4J060qbkt22byNTaNcusqernBSlIFJ
KOZshd/o+xIBSgYAc15m1WDMRifCzboCN5BjNuYL5hq7lEfWoxWOi7ae1hdc3h1H
6HOBtEf5wRxSYmtwBHlLIhOG3aFKfel488H2idvGlU3vuHTsnhjtXTzm0msB4iN8
fCwHC+LVodfN5sSBNEnc0ZekfuWj8jm/K4gH/p0rmMBGReTrMN0V8NXX2WEWu3Y3
+sBQTnGoMoZswtxihi3u1mmt6N+2Ddz08ftsyCa4URrZXxHtbqkzyO6Wr3nD1jpY
wMmq4jFOAmgXb2yfq+E8z0AyHGOZ7SLscA3nJ8UQBUSqjxFJqbRoM342cjmu4v3x
9UyJEoRrfh8sTs48cFopE0/WPku7a0SCI/7e1OvqiqC8MSvZ+dcewoYAneUx4yDA
LFJPTsIGxUbpNbX83R9a7G+0DQv+LZDd+qWsA9r1mFc/57vk2Ek1N4j1YVU2s5H2
TuelkswvvHdtjLn/w/C6NMDTflxyuLu24/u9gTiENwH0v5c7ym5Rk+UnHs8aAv20
O8UXEggiAj4WWi0NfU60AnRIzcPN6SD41ZWPyYbs1wE/ssrAyHI5CzL0EMa7BYPu
ITSuOp4j8mBDwZP3walVAseESEQQB1zhb2q9Tvto/6gK/YThbloBXpdQL1Re3iVb
nTvNnNERGCqdRspM1p67UccV5JzBPt91HMh7XERopz8RuwSTn7cIXoX9saB0Ey1M
rFGn4LrsVanwM252j+IOJ0PcRl6op+juY4JA/QqQxhXZG3fi3ncg07S9F+As5NtT
o/Mq/PW8PVXIrvURMVQ1LhCR3YXVXpjam+gT98uMNKXZTtNIerW+M8VLBuknmwtM
keTRl4/laddB48AnnRqfV4dzkCIhnsCZhW6j77SUZaSQcFDBNeMox7UNaPe3OMj8
IZGAK92vdhsAm6jsRooQ3kaH9Yu6aCItzfpsGcK6K5/CPJMXscJFkzCpbRsFmWNf
Sxp2I66DZ+xBB0522CeuYLTKQ+Ej1Nln8pEEKggAdG3RAsIbNFp32RanS6nDWs77
cvISPZSP9cUSDrq6C4D3ilAniV/as+tcyDfm6DTDzyhtF6RKWn9fQOtMfSt8Vgoi
n9uLywFCiIw3/tW9Yj+dyM2c/H/L5tkT9/TTS1D+P/APp89s49UcaPVOC9FevYLF
MfennoFd9iBZirLihFkil515O8pDBOkos1aAjBEvGFxPIh2uhu2KBsZxu9NUQ3xU
aC7S3LZ2kkv/4px4InoZ+dxtx4nHnciDyCZh6+TVukGlTcFTGqLDsJ6nwpzZX5Tf
3ccR9NjAFfzUT0f6InVnddD64nIIV9abkFNpYHF8ZDYb2igYFaOyE0rmDD+hi/I4
ujJ6w3gCjcfSb5gv729h61nMCuTN3PXGzwGoOiaIm911K5sr4iBk4cL0TjG70TZ+
oCh2QgpKMbU0jijjrFxstsiP/rhlnHQNUy3ZW7k+oTUHJoLDgNlKEMZcl1KSj3aG
DnGg0x2Qd8ehzSN0iaXrPL69MnH8NBNq6HWv55JTuMQdf/DesQxrkG+dSSh2qix1
1G20f1A3ptfr0jgfGBxJDICVS2ufxcl/jx0KF2byKqnVaC/m9B+09HgX/jLbRZtf
gg6mWeLyA4QSMLcIVWpRGGsIgTBhCKXIqrKh1EhblHoLbN5N450xKrbsuDf71Xyt
SEbS9gq6zEb8OKLI7iLg5TQ5XyTJC/9+gp6JbKY33CPh+h2pWF2GP65r/xkD+ZeL
+xR2WPxw1l3oWZNA4X0EaOkV8A3gP1NdyWiL8jvqgaBUy8Cu3M2qU73azxCHAoJz
nyh6lRNrS9/9R6jyKnRzOGuwpy6uzpbs/GpyP7YRk2Bo3Ohd7xENUEY7ApYqTYT6
mQ+/nsWlfF5FMUz1646CHCkv93bbge8az5b07dw34hbiwKGRsp0uZjY7vwWZ/Krz
cToE2fI1ezYjs8qPppa8AzCMRk1hyCYg8Pk4UZL38v7Jhl3XgfFewhPM1HqL5rlK
h5sryGCsIL6zll2hLvM4icmrimux5jkvD6d2IEQPi7+K8gVYI4m1/1eMMOCfCuy5
4b0nnnNNvh6uuXSGYIpGnPteCZTnDxEJEVdLuJD1UYr4nsqK96rrEZDSJR87GLcZ
5nxK+OHCxsSZJd7c1TlJD79fXqAudL0+iAFBXaWwr/RiSwyp6k5W7MBpXSa4j2WC
NwsXIYbZ44V7oVJS/QhC5jFGuPsOhA8OVDTbtvq8q8hSn24HaRBWBGb3NMdhBm3s
wMkhT1gtiyfySJFCBc3XXTyZm0leFlXP5LcbWGVEtjmIb32RKzf2I25H7r1mu2Zx
fZl0IYtpvGEsr5I3sKwXt8eudMV9K1Qy9Eh90Mx0cjx0elsEiNQgE4RTDMQI8SxE
yrzGZ3mbBRwAvy1R2IrG9su2TvL9LpTy1you2VAUQ4b/T4nKpTbUF3xa7dl2a64e
Kbw9j6sVMjfewF9iHqqSI8iMW652MXyxk+hji9W+shGX3mPrXmGJqModoDfDLxyM
sZlvh8vC9Bp/0UHcTKvigY9AX9o9y3fnlVnNBDQR9FAfMOAbv+zLrUXc9i8krR05
jlPWOuXKKWw4Rl519sGWkRlpYAAoUQJjWafAPAK0rXXC3bctTJxee4BKHrF8sBIJ
uIphLarLfj/CqqBizTBcZ2hBh2ZmuSt3iJcRRjeiLZf884XXyykHC6WgMALZoCFf
wXn2KKaJmrqyavXqaZOf/+BuJgKsZeOqJH40vpD7tviht9nwCnt+FEhweZi7cAwr
EZyO2rZCZwqPZT9+WlCx7tQ9Q8MR5Fe867mgyuWR5bIVDqWlcQOf/ZPdZVsfgUqe
/xeHUKzrSHEO/i7AR0qdCaOTihFY+0j6cuZVnrO4gLy6l44z1SN8vN/B7va0no4Q
N53t3awiaiVMfk5+uPuT1stx6JiNqj6Gpox/i3NdgmvpbjXMxpm6a7ea9RXLy+qD
xYz0o2yDYfgNllTmAG8VYzEApdD9W3b4N1nESKLEfEEBSTz4vktyMJ7+T/i2LLY2
TFdJWd2Qa0fMe3yS20do/g/ilAZmYuwwp6utTyDjfnMYmJtuS8i9KEzOrxlPOcM1
O4Nd5ySG+/JYHqkicvW7zyRwHQx1MjUqXVtXRZl4+/ZWkKcgJXtirvOP36h9vyMt
IuZhI73hgfOTh2uFff5WTSR3EqPe7rZopxcj6pl9I5SWGA5S0e7a1piY1H4J+tY+
CU0Ka1gpdTHg9lvuGNE7MMiNhergsjKZZFbR15p68E1OEMF/VsP46vhT3JCPPAKl
SWn3BFlifXcMF5GDcKw6XMe2cL18Q4p08Wp8QE6wgifNNu8ONNg1H1EVcKSUh8VY
yXLO+4/ORTYL7ttGY/VGyLBQnePjmJF/l+MFA1KrF9Ix74ydLi13mftXL5HDQCSO
u/9kdUIwKMhBanQJgyqEFIRSHB6xQ66KOgITxjwSl43y61TgcOWyTbT/wuvZ3m8t
amYIvxExpjljXFv8fbc3gMULTV2iYMgs7Fi8nP78QB8maqBJ//6IudNOkUkxlhXu
4JBvMNVkH5AdNZW+2WjjchK0EWmHqTTRadWuwxWhojyzumTGffvQD2SqzhdSJma9
dcS4OzAx/aD64Kj1zNoWoiZxi4xejB5LyxLD6gNOgYSWjWoWgK/Zo5+6F+qVL4tf
sTuvWeE9W5dmR4Sp3v4sbn079+k9F+HJxdGhEI3P4MuvR7Vu/IYPkn276fK1VYSJ
SxlDaMvsRkyau+pcuHc6oGaQ9dE6YGAbXfldnAJTR/jtYtunfZZ7MpFuRK6xRCT4
a1WF5dXn7eRgKJV1G4z5bjQCHuLiQFs0jnFjmwdCcZmeO2gQ1cLd1A044LoL/b6T
STyIgwTF4WKl9uqSehMZbDM4ZTX3xw+HCeICyJepRITD+zeEJeUTFjByQeWX/TZs
j/OxGFRWCHOqEHHfAAjQFrg1jvBjsWgXDslGBllf1838n5p4/nk4sUpk9Qv8F83j
zCtCQG3hURkAkC9fZ7QZ1RUoptl3n530aauyWc1CaJ3CJqiwC2MiYdyJ3HHUdWKZ
XiC/vNJ0k0+SaCBOL41rpHNnsuVxF5HWTQGN5LDLer2ji1Blwoocg0DqGKbPEvvN
Lf5YEgylD6n1VM/FDu1CGQV0YLeQjVvB/6+8o1AGcDrqigky/28EqnV5nScitywu
foMVtY+l5qoevx0njRV1hEtihcntZ/ckn/429zaXyIuwkWSn1lh8PwEx900AOFbX
x5LzxdFTrwHqSEgwE4qG6LNRkjXBM0h6x9Prgtun/ZzsWNv6GkLecgIYOkeWytRb
P2gw77Y61HaUrzBE+Fc0EctPar6zAVE8O+kGcHYFsRWZd/TSdG4P8oTOZDKPrmNq
wlHKJfUiS2/hPSGWgzy6BuQjD+RRwIOp6/5lWBOouF9y0eFSRbQa6xeoXeYPYV09
H5mYk4/+DmLa4QwKWxokJEUaDzlQE4YT5YQgpNQcVXEJ0MioiMoTJLg47Msnnc4w
34qEEQ1eFSIP8Vnt4jRCHpjaR0zq3u5jqp1cLQNkgzuQUdcpthjZhcwInr8Sy40B
TaJVZW5CDi6JL2KLxvg6+9aos4pupyB152FrUMnbMXj3HGmZpkWDwVhfX4ZXREA1
YR/FCkaF71mRYgL4iROpeEKcsMRGJNhdLXmv3fN5vehQg8vLToHBZ0glAJ1YHR1a
jVeJc0zjPwJL8q8OMpIO+IAWuCGW0Tcu6gAcZxT6vsKvbBzzVyhPvE2dkuydFCQT
vDKrPD1+JDC/BIe+ym6EIJFFahBmIc9v04hZGKZIhkbLeFYrnejlrH6hww724VjP
fjVTuz8t7eodAaL15E94V38MecTxLKkDQBJIOimmklJTa1VfWFVWifYAbCAMMve4
j2w3Ig3fr0fUoiK+N/WkbmrHzkERXn80e9vWTEMKuX9FbK6cu7LBHXfhNtfM4SMQ
8uRqSynwcWU1wmP1IcxS8112AY3kEVRE7CfSB4JJDOxvC3u/v2HLZ8kVz0mJT4Z8
Pga3fYc9+0fHlV1Xic2rUZGzqRx9S3wxQJFPFZgoiLBkEAnraj1X+DwLKAPj9rpI
29LttVaI8ioInJb1FcSE2nPny4yg+y7H72w2P7Byb0nM/dZo81u4WOhebdXavnIS
u+BtfUB1I96JjwvOVWdAUH16w6QepOSH++PWSIsz/oY/jdrbvsmsIrkB92h6JZ/p
6jpp7uS+DURvzpUbN5FV8OEaiNmkaxeTN+we8OlO0Vi4eUDDzIfmwHmMnWj8je2T
/NFRuYV0d14ViZDJhIFizHW1Cm+1zhkd182EufjRV26JucdIuXlA2YeCWtJt9Z3J
WGY6HCkqqZOPrLxiSvmk5iCymxuMgWHVoSKPkEYq5b7RAU2+iD3JEeSTArlMgVak
RtWa4nk0YGCWERW5Xpecl/ZFtQplcb24XXeE4BA4c/d9U3T0/iNogx8ivlUptM+V
G4/lvDBCERB+DwRhnby52eztXyFbmm14eryn4fvTvh45GLDq6fuywqglW18AjMdn
j31iTkfEM1sEp5WhlSepc6fed7mnh1/vBYRRdH85fYtRR1vULo7KSFw6EwY1/Fb/
Ck1MDsw/xjEicFZ8veefxJ1BSq7mQS6u3fuiM6or6CpwQlK5/DaGLiMhWjCs/VP8
gVTRqNtcByqwX13Bcn+/QTbL5Xx4NbAt9WIA36npWasaJmD7L9d/Vgr29xUxbZIK
7KrQSJ9O44LAHclBbUatc2vf215vOwgGufh7A9aB8L4t4JWUSMFRD3G+f/QTh2oR
XExSlOHzMtlk2IDGjOwKLc8HwTKAlmdGSx2JQ84L94IMtA5ii/6Q48Tkp1JlzHXo
bjj854pdZxe9aEdEYnTGfi3baOsTt0TkU4j0JAB5QM1k5eSj9nN7ETGia9r8puYf
Fai6Pukh1xSmslS8+LuT+owcFHoPab/CjK8L1oBcWOwqRJ55b9S4Bd28aaG2aAFJ
RuT98EFayRqlRmjBdsH6BGz1NO7ijs3JifJHNiU8Klrln4suXvqcdxjLZb/EQqCE
E7yaS4egcqtcEFOEe40zfMyaBCOp+b1paQYI9Zzz6Jw2b3SsXxTXLtiw8owCEhh7
JSbwRg+ZRPK5pyP8uRClcGHDOq/XMIw/wzgZo69ZAugvcwyTqPBZcaW4oKTA6ywc
Jn2o4xJNYB8UYM/wmYzbsE9fD7/niAcNSc5IKb4wU6XZ1nlJJFKDEkVp6hva3COS
xnvr0pkKtbihZ/Bm9RROZ4UmRq4+d5VN/E1I28hYXSI//sfuprE/aXJGkYnHG/PM
Su9JBynE3aVMMkHm/kOBPrr/APiogIXRhE51vViphxP+VavqsF86JbY1QNry7UeP
hWM6C2+tnrasiLZuWZJF4mOwpHgFpMgmPhsze9Ad21qgdP68jN2uMybbZldfUg9K
kHgWunXyx7ioOXwZUV/wyZ47scdzCTdFmjWUJkbsfvyhd4ebfuk+Npns32MtJcHd
EExnH1JQun4/WecXGEebqFHMXJHF9amF/sbbHhekXdFvreLcfEuYGV/nNF6yPIiN
J98HrxLok28oz7/8Bein4x5QB0W47IDhxnK4j9frt1pqA2uMWEAzPsZH2NRizjS/
1UWEHtwr2/a1Nm9MYaubmYNHa2SOqXcALqT3GsVUoOSu3LV1l9zZv5mFr+rNbPY7
ug+5AU0Qbay0wb1ONd+ciyposJRkTlElR/yqLYYenqWEnx9nMIr2Dux+epkenvxH
ceC75j4NrSfvLyuuyr7emciBH38HqyAF/RWYkxZyL7IRr0iq76B0MaDxU4bUpPG1
IeAP3NmVc6aAlz0piAmwFP7GUQKElrEkn0mYrEgr2kB/lNdcFtvV7ZhTpR7MdEmq
utd2kFbs6wvhAuR6X+oCoNUvbGNwcE2BmYrnFyhJnN2dDgakpiWiAZ8t/dSkHRbl
/eK1OYnURqW1GhEVhRcLX3s623UIAhfvNuYHRjQtmJuzNpIuiJnWz6xQDruYwB2s
oQpuMMTwhRmOHVR1c4GC5yw/nijQoQmQVoxEwzAmYHpIn+mPK5Y6zJOekzNp9oM0
IqTC8QPlPDqTzT/Jf1NcUVi2Q9CfH1wDvYQqp9kPYCL9IdmypRMLOKMqwP38SXyQ
DE2naaFN6T7RArsw9q9mTJsGF6VptJmvJdC5gaWixrJp+XUsC477K9TI+MU4FMiz
11+66fGI5eCiG+EX16xAMB/kuRBLzoeaM/ynBFnloR/0cVseAPAkoPPmqY5gC9TW
HXUXCt5FElcWgy05yj2PkofuSXTJ2y44Owzdgxv6NLjcZr/SePyX6/wEJlCgmPJs
nK8oekQ3gj7QctH2M2t73Ua+8msQo9mDxhyzYL6LIXyoVEaqZ+FuDOwuZZtxz3Hg
h4UvkPxU5OM6QdUVvx4FYfRWcC+p7eF5mVcYvkdF3k/TCEcqtcslgCns6HY05lNa
VlohjMFQgxM7+NsiSrMHiY/fBoZIl79BeYujN7kN/Pfo/0IlPnEFd6+fM4MDMEhS
lL/izGClzqQYOL6B9rJJU1iNsoVXLI6KqUMYMC2GDFwxWhqAWjnALFRecEBC4Tac
d91oS9jfP+NwVPtuIHURvakDOqj2LWqDrvcTLpf85jj0LXIRJLe59h2AdI2ELdW1
saT0Y60r/2D8spRR4l5F4X8OFq9juUTv4L9nqKvmShidjIH3JsSuD3EjvCFI7EYq
Kzd947bKOa8YTGvV7AxQVa7gBR8Ob2IXDsZsdVXayj7yBLd1E/KDDFeaG35HXGxZ
Br1Pom0b/cPQicGx3XNhxnJ7zZ3S+I5SvOLvQA/BViOCXpndk7s9iDX86I3y5tyZ
6UYRd+6ES1+8I5UjPrQjwR58t3b8mMARF01waT9GVTVo5sFD0AvuBF5TGuDsogcY
TJrHL5w4AysAagYqcK2DxABD0ovI+cIW8ZPl879rUUI/FI35Vcj1ywW/DajVTAm5
3465PKfjPQ2YaF1ZUDKyC8g+t4L8ogsti56E7EwJ0N11k5mp2k2ZWSBnkd9izw9c
JUsMajmN7SKOwAEhKYf5FMWr+xbTQBzQ1t11rfbCACpBqiF/1s5WFvTHTllCLH3a
Pl444hN9RI4FfZA7oXXe/1yKqF1Xis3TrTl6ohjmyfiyqChASEpoIewTNGCreJVw
Mdr2Fa3n2x3UThmZ1IhkMYxPVL7PhZZJ29D59QjROlOAX+GOOy/FWYla4pDmZ8YF
vaBm0mr6gXfQA1Wkc5KXjVLfnCdOs8f1nTZGsMq1zLFVhbP3UCRmoDyNLxwYCUw2
2xwiboTyVPvxqenoubQrlvncXg7W6ZcCv+E6YdV9GWcPzlIWMtAyV56+bS6KNOkj
tpUYRHMiP/hSIB3gsScEmkc4vlxRAirlcRg+aVeJcAHRCbDn+KBvo1cizHSvnJ8n
LiUpmUlD39+RZPtrPdSSqOk5saYM1oEs80CAfe57lO0ewou+XwAIi+96PtPN0IbO
hfwuDob42bq+UFQY/6/Ai71IMf4AIn+nMAsTQyCYMc7sXmcFOsHTIkT77TCil8Zv
uekJvaowz2YkpvG8aNfPaY9x4sz+BQezET+dMVglZseOG7n1PNL4M0VlD8DVXh2y
HrnmzXCw1SG6brEi6S9l3/LkXbQjzOjkDYQ5N9aGKCyaT3wQmKrVuDdSG3pYbfS3
jAgABMh39wZUQcdRW4e2hTTUjH74piCPS7pHFRRc0aodl+ci2PI281w/mZ9QITUX
Odt//3SRgOxx17AOn5eAJ3KR5+mcJFTBBt8NdXA29hfr9vGZEOytbYV8B2WQ27sP
Jk7ZdnB6lARXIBGZ2SW8VxrHG2ZSDDCJWUsenogwotgzgYFBSN11qOBQ8JmzZsnH
Lj5ozSo57Iy5tbkVG3VkreCvsmFelQZKLOGR4zWSIBnsbv7UvOG6eivdVOpVMENm
lz/sfX8s+AoGsBKEWBYeQtrCV9Qkuv7msXOAh0chCqPQ4O1eljk2KBLj5FEtkSv/
SemMu6K2wPckAsHB94nIs2/oGgMwefaKhkoQDaOgbLv1iSiw5QpCS/y6k51yBAEL
0UfLOPu1AkmyyOFdoJoKvi3cM5fp1zRfb7vilTh3F2egEPI5zFPPO8zDzw4ZNmlD
fOjl5VYz612G2j146fFfuOi9zEoZLSYA/lMEDfJdxlJhApOiTMXmLGBy8I9wIFsp
zM9aCs5vlFTh71ROIP5uqbGIg3cARSje2FUBknhO3NFdrsrzp2pS2XxUNTcHhWaJ
Gfh8Eq62CdODom8kbh/JVo1Ia/hBVappinOdIzErW7StsDcvMggMU7XrkF3ojdvl
9xmOlR9mVYnHKBvVI5yZrbMYpP68xI4zSnzHM3Y0tIKqsYTIG54U+pMHItGpHuaQ
THy1y1ZSWbAVpkUNxRrm18PnseNM7NgqESkar/YCY2tsjRWcutXf9IDXDfDJLNUH
agA36aj7Sn3mp7r7vhZOyG5u0IlqPYUYp/ayjAuhOKAzGcrAmRQg3m2RmGskwAnW
XLX0Hn3D0YuRu2LwecUqQOzFLsSBzF0twXntGLEVHkEwWsf1JnE62DRVD/KQB3l+
sRLGh0n5nhKgSkGFiXgnglPbtYo9+s8QfsoQDiWJro+jmc3ial1Bs+gmDm7iAzVu
Bjc+M8qcSPSO7vcL1VQQRn+1R0YpbkgYOuB4o1KXo6jQuZRCElAQmBssUoSkF/1a
0uD9nl2DzNqp+5tWF9Anm+JohKkdGmmp+9t03kGwHlUAYswdberkPjLOAa5PQr9t
W7ZEsYL5tBxYfB5a0i0giPrLeIETvW4h9eM+5rxooekdNYgrDCpoRvcchHDHYQma
l2ryg0jOwF3udV9Rt9QZwnoIW6QmyMKo4JXGBptyMmw1kbEWkOcAg6CyoxtKupSD
GaTSZ6Y8ZQsg0Eapl9ZNDLq6pXAZLfL1F7z4J9JMR1W/gKUeqeSpTYdhauyOl0NH
wubWzhCDL3Yjs7fLr1LHbH/UC3U/tUswgZ549vxgLXrJkOWh0bdVfxObbIdjIO41
DjxTZVsUwY19255MkTthXlv0jivJrfqAqgxlLIRQ04SsgolG2HDs7019mij4336k
ZbxGdSaX1jlNDeXEKd8nCdf1+4mHxyBLVG174Pra4qveMv5rCfXcH5CNST1UvlcF
XWd4o0xUSO1JZhaxu6blYoS5nN11uYhu9wcoJ7ZN/26zlXMtg7QSRmIbC0QBGLLi
ZCQAkX0fq/23B+IHT9mA5sWMMJKp4/z9Vtxnn5hndO9MIslNlpeYA8yB4huAF+Ys
E/GfXsPsYVSiFId300X6c7qc390GzvCrfjnsnNDApAk/bHL0kEcXYzgu7Av+7qmq
Z2TPt0DwN6s8GEkMKOalfd78WkTrSU+pExjebqTqrBT8IRZeaN9UNRscyMWj93Di
xTZLmDoPhnApFaXZ+U2out/fi/5qk4GDZueXyUCeO4OStwCJKkle0kjrPC7rLPDj
3aOTbx9ZiuofkkZS0xoqOwISosCknVQzTT8/8xDJHwIEjB1GyC44AgWrknmhQKql
ZQMtnCS7pASSJuSxY4WjZX4f4LVTY+NplgvM4yKJETjl2kRuYuXCnSMl9d+5zNPU
3G9BW1Am/u1OfRWf80XcG5QfS8MpfSEPPvzl26Aun9H14mnlOJlZ+BobCEgCtoLX
41Snvchrja0KtK45yWVSvmrYJ03+UDaK45QR8CRCw1M11bg+L+CvxY0ekrjPq9Yn
FDd54zX6CaOxzf6PwXAellSfSR6pgBglIeZ26FCOCGmYWCgKoPyZOT8oE/KIXopP
cIi95jGkL6ICNNnKkdaDm+bCEt1s8gbHrrk9R5hXrFKGGkuiv3dPqIz2FAq1nn4e
ltO7bHR627VYwA96ajJxdk+yf/Kv91J81BqtROolbgBobBiMvru9YM9F1IKkcOfT
weeEOybhuCMjvKB4PqWx9DW20j9fcHbhFwEEK8J6bkD4hd33dQBeWxsiENwOKDiD
gbsatbqIZXPO9kQal/cGkXVZPWuRTcNDnq+pdnvdShmwz0Khf7O2pFPD7KLOo6p1
trJGI6o6V31kXWjC49WrzAK2/CO0MypcjtDIJItEO/n9j9yTP9b2fmFvku5B9kGr
5JJTRVCnK23vofz+mT9lRC+JbfQDCOyxPOsvtQJLXuXvNYIePFdvfpq+FWfpF4Kc
FHbjU/QTwI9BMQut8e9ZdK3ySb+gnv6W4GU/FWpXiDGbhGfV95IEMIwqR6z9K7hW
xn5O68F3BbGq2qseY45fWuCTa0/GeT5fSvdV8dYLo/+zZ5Wv7Epm9pKq8DiOl+Gm
toyiaWre6hwjWfcPA6Te0CyQmkfa8htpJIsirj9RtdCCMGMcEQz115rGQIZLTPUS
RTpctsyymbcO4ZKgFUsrB4bjL7XQfZr7bd7ijaKviUPHWOmplgWYGyY6aGTnhP2n
nJR0XsswtzU+Z8FbNB0M11u9aSrMKYzZ+RjndbhN59stIQcPlOVYEIxgqbnodr9S
7XCNNQfoVOQI8Z+oprJpnCMk+dpd0vEAbmy8Y/eteef3+RKRJbJJKLHAhGIaReXg
KrlYfvPepuZU5MMT5ozmAnMQpf9uIgu0nkI9nKsdzxIW0KERi1BjSc0eOagH70u8
J+ob9EfZLeZG5d2JLbawqkHDJCr+7WRwGZ7SgbNZM1xb468Yneh745wD+aH4X3Gl
kp9yzJz5yFjPoIVSRdjBZ0aRZi7tV7k7MKiqTiGZaWDvie0lsZ+w6vMFW67i41Hd
F93Uu+b/cyyeai5/Pzxj3dzGnzbRHTiPcDAQ0xEMEbH6WWAmAM8TYb3hIn4l4wtA
LQmqfOlNEFJLpQzAp7v2C1r7OHKCzWbQJGvXz+BDR9ZgaKiBSirv97zXMW/1wykl
PEyeq3dUbnZzfk7OUqGBaxxMwyJaZW1/lQ3e0TXLdWg/s7bfQYijHNOHWXlUOhHq
GHQINoy63Y/e3LOtUyPv3lNwMnYzrx0vwuqPrcb86RcdLb02FkkIMx1SRzV64Ta9
RJzo4KCCtZuSJXRdIF2Qx4N/+UCZRF7lC52FSMbG3SxcZvuvk0CTcgSeIwt0PSKs
Fk6LwBzZ5CqKzoDVGH+tKT9h+tY8GwGJV8yirORNLCcyX2f/pwyFRC1f/UNPPCB3
F09JKcozmJxZYbycpCkpG8fT0YiNzaKtwQ5TojJwtu0t8Q/cguvDHL3mFRDFwNHu
5UsnnNgH5ZnSSb8tjJb6YeUXXVqTyJurx4uFP59zJT3L97XUa6rP9Tefrsg5vSKa
GAFrRI3P09dwqeDhlPVgr4ugZ4rfHIl1FaX40SLcrwlAVAZt/CklLf2AuNavhUq8
eBnxAYugtClzvlKSnNhB9WpwGOBC43NTc/5RpanSNNcrMIXf5KhCqe4dEfhxWGRv
w1fK42v0Iis097asW3UoL1o77shRbuD7DG+lvM1hQmxRmzhqM/94m0gD8+hWC3j2
X5d6xCoJ/wKApEPexGHnGrmzaEITm8Hb6Cxx5ysS512zTxWBoT1NG3tq6XAWEp36
0JzKFyVpK+x7mg8bqC7VRPTofhLEwqUKLhANq8A/Jk2wPCQI18/nM8fGxQcM1Zn6
7YTl/3fmdeDfxy/iPRakqqn7+xCDCk1MaDp+D0kbSavNJ/2YaPntIvODMWOffxns
L3aqDjzATUMYxOR/op0doaLrYk7sxDYx0ALxKcL/9q40yx2wlnNJ+JLGLtOikhQE
Bkp6gga4Bzx7+JZS2B5SfTH7Hf50XbZ3byoSNB3xwuOlKBXMiNdyEs+8NMtNchRD
sObkO8KJf8AfEJcb9UV2SlIxJJQga/wu1N/yMvQLMv2ES+LgClhzGSkoW88BI1tb
XwqauhLsgZl3khP+mI4D1W2M+Owfc8p+OoBILKHVD12ahEEd5mQoOFou4e7Z/dFi
56YUq5acpMk7lYbpOiLJoZLshPAngK3qPFZT/pH8nMGEtyMF4pULyTJodbKEJ9Lp
XzYZ50j8xbjm6oDw7EQw9b0QNh+5HqqQoyIruFOg+nzjdezUkJxQcqdtKtxMSK8Q
Yrseq7Xoc7/r2rwd0kGJ9qqlavreet62c1fk5C9e4L80PT5668lRj8IwABZ9rmfm
OjWYTYyKOIZXa355tcJA7xuk6avA99tf4SOnmKq2meM4K9CQ1OqXsf1jQTJST2oy
Ua5sgsQBZ629gjWuIQujKE5yZE+05IeR+0fPmWm/s1rqDOAROBRI5l/3wR3SCw17
lZwVhlXCVes+D7ALs32nZvyARABOdEKeJMPUTR2XmrjwAzuH2axDd+3ryrKWI6U+
ShKv0S6uhdIX/W+qWNXjyIJB60ojMNVjftEkn2a865xj4lBGUs3zzrlN6CqYZGxX
gOZ3W5aWi/tInEQBBzRxuHRKq7c35BUNGkT8CrwrlLbxPSo6/mJkXzk4NuM0zKK8
EcTj9VoNykXBf7n8yznVI+wtJV0lIfbRmKXs6dPsvkwkc0vqJpbZK7ko6gWyP3v4
WLd2bSs5Xiaxv0vuLW0CpsoR0Eqvdm1Dlh3HUmnkbotrxGY7UdixzpsKmNIzx4Z+
G/HYFVwE2u83PwQXdzTl2g8dYCzSPOKiYwIzc15kdcfkKXc5GuKkVV9mS6Wpr90Q
vuye3K0LdDgPR0EB8Alj+hzIgEcGeKgbdlzEOs6EhZKaIwqy0eY+gZwfu0ZMi/YN
WuYd5hiBRAQeF9DgRuL2v+N3XYM0pxTfJ7wyNzaNQqZzsM0JopFTGdCivdr5YDSn
gn1O2DGbeP+H64N1iBSyWGeX2AomoZ9t6SeoHpGJZtryZTyiCZ1gbSg54MpXqqPz
aBtMav9c5yPR2QLPR9RtQDYc2KKA+8R9bpGfKstz1Iu/RGyaX+YELvXeRwRvRCzJ
pYllMtvQN2z3srot9JoXD69TR/bkEF+GMcsYYQF6Y4GnE2cMUEVNWiGXZRaFn2xt
mOFpW48dlD+khRUE2rD6WmFHMQHpuna7HkbJp9PZKlahGJ+NkQPAfxrGLXf3cWTK
9wrUtIssIl5BjKYIAqMafBjlymGTPaGn6zYDT3HhUImZOl733VGa0MlR1Za/HJWb
WpxV/ZT9xYHC/D7RUsZv6PhMAzQumSdD7llcg3iGUqlFbnQthd56DjXNrnq8acqB
EmTKTbCLs0y0yBcHtt45zB7E/5gCuzRPuO1/stDPwMwacc/JqTD/Juy1uibTB1AF
lGdGzeOia9RgSHz+B9Do7yfvUJLAOWPqh2ufBcfyuNgmxT8p4e+gT0JJclajDx4x
MoNNizc/fRmzzZaQMJRHGgY7dkHk5+ckIM8/Lm7a5WwwpsST3tDTzDvqb52HsT39
Awl6BVl4IY+ywsgPLiuBXchC66STnJL65JvDLpaCK0iDzxYC2vLHC21EXWVjk4e5
pn5x6NC+0zIqQY3AGEc9Q5necBfEvdRf9XhHuwNmQ2Thah6Fb+t68s5r4buoBybX
VR1tHZHd7guK69fY/7PB56/IIYqOt7DXP+skqWEd1cWuiJqHBjrwFvHDqMgnaLq/
cf6a2okEprqUHcZxdHu/EvLO5fh5i77IYQI8nkeJ7Ebo02ECtdvMWs/kZt3zNLyo
ApJvhm8Fu6/4fDSW/xw0UesG03Mp01hGWs0Af1yPahu1Ks9Nfuup7c9ePpeGNvBT
VKtEIxcqhc7Fn6taaFGEKVVoXHRcKfB9Mo8nMwlTKBq3VpqdWPUuEYMYlBNcNLXR
WfYwE9YG1pLus/OoREgiGmkJc0MbOclUov6s7Gm66Xk10wYmjOnZMg13WGGDDF1/
pSVDeMqnows+6foTF0o3B5qjyPFEHV5oC7JvZOCGgu/2l6CnM2EDRIi71Kgex49b
y0hZKzKLBEGgXDUxfMmhq9lKpmMRsgsU7sKioiHJmExP+YX8VoFdvlbLKo8xDEid
M4K4VW+KPldfh3S7Gf8tmgVVFLV6oX8W3WX9PzJO0sZUqFb75oRYq1szqE3pavWS
bUW8hqSJWiPU8R9lGWak22utVwPeL2qw2kuy+zjEHmCG1+X4PON2Cuw7fw/SDYpH
2iTA2hvup6SnrO74W4X8747gT8+NjE4WoOZ679Ndvd3YdRPS0/GuKiD5BDvux5ba
0i1+Gp+xJn21+XrJo5hWdLqLEUJ74fkuqwzGbTC413/QfnPaMFQ6QHdE0RIaZofQ
K/IRo6SPSrRe81lmRy9HZzntHuCHKrJwQS+J8SBTru3NsSyz0pOuFohJV4fFTplW
51332uRA5uL470bl3D95kXPXCoPm/m0nQsFGuHMHiCvpE1Qhy7Qwa69V1ruCAuUe
XXKv/qwsrYdrPdTQDxjPE3eoQUc2jUhRFS+Jr9l1Vr450ijM6KWdrEILgl/qqhmd
qniyS4f0G5+SAHrrcwu1fD7P0RwmhTSpBC4nHLd3WO/c0L88HJ0aZ2X8cERSpIi4
032Cl4KlxU20UFyAkcFunY8+cpQT/hOdc4id42QCRV/yb2SGn6ZFKPPsk28EAyye
Xh4b3PdvAjauhtWOLN8X7B4EqprFV4xzVlAY3odoeRtehvF2nWsFrW8Yl4dgIUDF
FMz+ijrGU/Ba34ETFIUnzn4vtx/u566TmG4nfBcfg7ZHeUYUaYQ00CKgPncR6XX0
egHrExLcy1j+zciHJzVlEcmXrol3E9JWpERWLl1AO0kas+zmDtwR2F1qcbyUDJp/
1TDOVEvTj09/elXWe2WH4jkxpZFbSbm9A824AHQJmfV9G2MaSLMQo61rVP+snx1/
Sb4Cgv8oTGYKDX7CTD3OfjPQ/0L/et94oj0/RJvwxW0fyafl0L9OeJrETPB2xUOG
CnYNoeBCYyB0DwJ+QFUit3im2YaRWlqKWfau2GKUIXgV26Zo7dJ3CNuLFK8VkKff
2t2bpJjLbQujfdSTZgPcL4QH+TyuaWQHyuP8ISlNU/KWfoe8N/HK08Qe/rJltRyY
pxZSXGguYe9H+4UZlwxeMhAlJJp7WZ4UBA6cZLaB0Ja6OA6f5YINW5NwsHnV30aR
BY88CqPBdQpZ8/pbeBYSidTtMuYFY/fXD9NvRoRQsRrZO9H1LBq8+qgSXdoTKWwH
rwdu+AAlFsvi89Qy54TW+Q2bvMKLPzeeB36yeDcoyUudp5gxNkQwqhrikvdI//Ub
uJqezY05kYmK46paBUQviszaLhOLl8Zs4NN9GvK6pbhlQq43ZH2hpb4LaJwUcuaT
qdkJRFpzdTM/pFrHkaeL3Ev9wvJ6Fj34/EnWMrCkaKCLnNtJJWB0EbOiV5bjsKcB
yngGKhxLc2LAjXjF4vBZ5ezoqCApXCuErcd2E5CKtGbS/FzZBCgDSvx2ZbZlHHxM
4DZ4FU6V9GllRpTFZSAi+hxHlxzIHTDaVmhiDVZ8i8j1PSP1m/mGNdshiDJfMmmN
gcWUOJ4/LocjtUQgvzBXwJnkizZqBWFw0pnDFf1kJyH9V6tfBBCl0LxFDtKXB4mJ
not0XAkB5MF+EUeXHCD8/yxm081CBltsfuE/pWRqFLdI272zHz+yrZ7YFNVqjkEs
GGVrPrivwdGPiBV6OxIPlrAvSgcncYGFw7/Wfy7iSqtn1yccIOXLdTuw0dyPgJLN
+wM5ukhLui/IoM1pdPe7pJ5oKegX8TLGkmEwk1qLnIZBOxAntZn4qdRhu4i2B30m
Q+VHGo1wh35ll5AqQzvIGVMnbcNSdZu3BUZWChfI9Ksq5lAl8xxdGwggPovuo03F
6B5ooiU1zf7zisPbDJm7hhKr2sBJliwmS43VEyxsqAqatTOcK+to8EnsdlBBjFgO
n/qwXIbnQhn1/HmHPodFFD623u2XYBercF/msfyIUX9gTYHY33b52F7UWI+Yqw7H
zUwK2+nKE9ex7C1vZrue6alb8puus5Li30jHnQK7hTwhVcZnCh7DTiDz9In0kBPL
t/WNkWVYfyUC8YinL8mlaJpe+2zdQ3BqJto9gqM5w8lp3CrKLvbZQXEX5Rhwdjma
1TmKzIf3I9K2frZuOoTcP8eYj9qameYKAMutKNaSNH7YRdm78JgdQGCZG4ghKs5y
meJlyYzyAwgY1+3f86nB3WNpGdg59s1dMkWlt9QZOFtuS+iy8vXx9kDonNfbP0yJ
Bt1NVz4Rlc1LD3xDrziFehenAsiSe+Yb2YVvuM9h97OXYS+Ltmwsknl6q0Cl/aA6
8dU3brVm4wvSp/ov/k9LsKJdn27lMzuZmyvNZJablNoA4IgZRUO/QylQFegzwEhZ
IMZiYxUqNUn+Xr3XBLo/r1ynGi/Uuf4/MOfsVk+1+8zDJvNGin1Gy62nAiKnyQqE
P/GrnzXM4OIalMRTOEPIlOpUcGdN/vzp0XZpYAH7ZdF/+PuJvmNh0ept1QWhKvh5
yRByJ3bFTSgSPa/tJTOjjR1p+JWUc9/8DuoR8b34cfZTDVtEv2NmrhqjJcSMUvAG
T0uvZgNPJFyMYk7Hv8jkfKEtKk/mLpfQhfIuqSzBezHopbFvgcIYp4uCZ1gOhKP7
JMiAxRCROsr5jS8FD8SpUr7qHja/eByeu72nDqexDcYMA2rdo1fMYF/fbDvKxeE7
yb/Y/Oc6G/zfIaZmJC9xj9HOzZ/M+XvcM8d9+6zyFwUK9FZRZM/vJOM7i8GMeu3y
wIkuMCaU9d/8Waylc1tDh3QcZ9srz8BRMIwysZiNN5tpaD/ThlBC3Aj0XqkSe7RG
zpNXAZ8boDMw0vp+ATsZnTBCmM9iJK1u0Nxp+D1lSutmDk9eDS3ipR3QQXe7NxKf
/BX+pyanTu4n3Fz4oyF91ApFMvKYY3sfM+Ij+eznLyQh6qUh9kSMmpqW571gRujn
m/M0rjX86JpIOP0GRCYdyxvHmGqa/kYNoT2D8TIAeKJ6GSPBMh3x0ysv5ySl7ahw
aa/SoBTImfop3BjsFM7Z0ZujHfeKKfn4ivJlGDGkkBEGnvJmGPV7DRNi8MD5Dp+K
hJYNAJb3LfU5DEki7k8cXCiqr060pPOQbepyVyWuPxA/BkXC/M+QJlnsmQSIVmwA
Ct+6qoRlkcFrVmnyyf1AHUtmmXYw994Y0aPV+Tbzro4hgahmxqToQLJYlzlATi+4
VUWOvAKLyxZc1X3JD7DNhMBBDuyDsxAossQurA1dExYUOOt54/8dHB6eVgOzqkNL
kLkU8JgPnBRJzN9YkcvX+RwsV6sV2eeoKzq0n3Z/g6UFHaj+3tBwg6f8qbEIFRnB
jD//Wn7LL+Epnwsd94HRVkkLHu+GAL666jWB0YSB1v2fKTLrlqALhfHWJSClMJIX
liCuXZW+e/CiDgyNguuCs3SaZzIFp4BizUsDTrRDXohgxS/aBUB6n14oMjVE4ltF
1oUhaCJ0y8KVPZviiwr0IPAY5+my+3lEIeOXcqIP1SyzlHOR6wL3HATKqG1dkWks
ymEvhu71bklxCVi9Qu0XUXQEiAsXpy3RsqIDMxvpLwbUVaOYCxzGHV7Q+5YVvuda
6NGx4Cvn7MMljzgj83f7VwGa+wko4AjiC8S26wXp103GCe7iVK6uu8nWdrp8OcJX
OVKbbccmvxEx0TmIXEsaTo920MTLA4lilzS86O1xoDFZrE7+kKRhj0rc4yEbjIzU
NP8Ry6f0sJ2Wv4vn/04+PXo/ePPOtgiOn9UAu5uk/o0Ih4WphpYhH7XvmVG7717m
yvLaq++LvpHx0qxf8NsdrLPXDOaoobjpD2LwL4JkKLOjMlW6fhzHnnPhA9DdQx/4
O6hNKupZg16W+Nrg1BC279HAnTis6JU57EbvXsV33PPC9vYtxtPP59Z2jPzMu7hx
LUl5VvDdQ4uDZLZtcrfscAWWqm/WAiDGpiw5MtBE6qpNa54GlUPJ5wY8X+pm04gR
gi0Yc0K1lerLCWw7WLore2u3pkQXESJ9PNLxRI7VJ2bisabkpQTDYp+OfVKH8+Hv
zqX1Nhmiu48w2HUOWF3NNwXdMh99rjd1bmx+rPemMg+N9G0oXLUFkcyT5qyjGzR0
Bq5ZcBaykJXavcbA6RYFPq2K/jDY9j9N92i5aC7XGD+4Y9JP6u/M2HZDq4Th3HRH
+NpQgVPPTPY2ByIXBQwuYPCMTGJRbIOyJDs/95apTKuHEX0SAFFDyggO44O2sB6R
lkMlZ6xwbFQfFn4tE2TUg+J90NVUkh3TOz4pxfSXBtqhuIkMUyWLBZJPancQc5gk
fYRJqOY4oagVxhhiX4gZLxtoMMXplo3193G+2EfXKg1PxZSgGl8RTIkKOdFJD+Ih
9UWTmR2ch5EcYv9icDLbxZ7k0zzWAhTxavdYLIzIpS/Rw5N89Sih5Gxn+Jsm1mYH
izpha+6gqwAlnXxE3VpcNDTh1dQGZQ0N2LFE961C+OmBgKd8tsvPXeDQ6wRDX72p
qQHv3dv85SyGYVBkzg0EBmt/KwnWZVJbczjdSIOfvDepDpXY0QIu9isFKdvrC9aw
WsK5a6U07lcUPNf6ZgYadi1Ng+bgobAe0NePfLyOpuCJjsxLrPyfNMPo11XZZSAk
5+4WJFA45MIsyECQ6ypgXnj/xVQq1QENVDp7C+rk1mmelSLCCfqXiD0pikRqDk7e
DBdyt1mSVFVuPYUcLfgLxq/LfQbQ0OxK4MbdLmEMEYnPIlVShfut3TCUN0yX8uKv
e62knKGEFC3O1jL2YCtfzR9+w2Z/ifkLZxWoQd0/h66hT7lUdP4uYtLyRGO63xVB
vGOey0mH/M98HRQV7y/vW2W9qoNeBSE+QF17ZNXl4tXQuWuDoeux0DwhV8DPlI6q
e6kjO8jHBkaBB7y6s0d6GFPkqUVJpPCZXnXQNnAlds9+p5ZuW0pjh9Bfv9Ndn6wv
R1SGKYSZbPnMZg6KF4GimbSJE/7BSU8/1CL1ptu4iV0u0Q8A6btR4ZZSGQPqiXpa
lZeR5hOHkKQ8Y/VQbJ4LrzVCGPYXoarl8qyVgCf3R5fuVXZseJ6G2+lR6Y3dT2qa
G+zIghQLXlBDugMvkjJqunzkd5ADELPrN7Cn/6ffHEewLqYbHLGR1EhSx2Jb7i2z
2DhaGYhYV4JsyTTT+TAxTG+umy1IqKOBbPT3QGxcGakDilwTEe/Wzmy6kO+JvM3O
vXictbGluDWytsOlZWhXhV9Sfidw7J6NESigMfug7R9TRCfv/P8cdTFNC9N+KwHi
GLMn2S6HNhJij2vgDyCIOEc/L8boAzmu+FUsR01AsroSQHH3s5gDqgPAk4SsjFDJ
DsZ8zFhDJ+EAnNtScF+YuFM/pSwzJfY98C5oz15mbO8aQISibCWNR2njIVMA3Tep
W8V+Z+vVFONCEx00skGMP9cxM4c/yb6bnL0oY9wyMHMIZr2uyt3ibO2ycmWLaUw8
3S5WBtbnMTgS6FjTF9RwMIrkBw7UmZbpTf9MVS0PJ+KSJmrbJUgtI0shm4TjDHaR
nPRIbdYvCknFjm8k+nwT4tEurVAGAMXR5w3XtpGCuvxcJt26Te3xllg/8tzV0ymG
eYGl5CHfBYthBQ+1F1dEzT99/wGipd04iAVMpfdysxF76OzFkDQN0nHiEk6Lh3b7
IsBbCQ/4mf3e1jZCQgIdKFVpLXDEOJ+qye5JefsQHBDRGmA/DZ7S23RMv+AKqRgE
gE2BAhHXrMz1RgrltgNrBYvHn8ibKesYjP4Ncylida6yrvCtbFVUWT/DIK+pEbsP
ZtMqdD6f+H75GVBMSDgPrGRU6n1lK0wLuv2B3GEGJuW90PVfhuJsonFJt02WzmKV
C5zAhbYaZBzWAceBU0PKDm0nMjVkRkS8NG39S86cECAWFEoC+iV90tcebZzxVzse
+pkidNGoqAAwGxzugn9EhaGlEdLcrp8BBZNxjnUiS3vF31D/OwNby3IZDcOoin1S
daD6ldZWczxQexPqPYXVNjIE1k/ISF3I0GbzKyyolo7NijHcbfooTprPrJ04KBtC
+L2Tz0YLDkmzX+Gp1y90qs0h5EEkbFroBFMYnzWV1Lcp0Lfl7ZWtOnqkZ7cxNOJ2
6yqdM8RXcUfdFA5Pur+dLuGaUqF949Nw/rtAGrhvnjmO4oxnZlKsR/UXt3qgQoBw
IO9CVuo2fR5SkcZFbnJaOPgl4hKBN5skCSVgKilsRSOr5zGg0N/c5KL2xGkLZe6q
NztVvktX6TvetLNNDDpfWGydYUAHtPt3CFt122juzxQeiUfqLZQqP+p1pRTC4z+H
jn6Xqs0/xCI39IONeq1IsTUcJur8EN6t1DFhW+F/OmeH87lIkLbqpNIi5IYeCMtz
hrS5LMXqpi0GhFjGs3LI+aPSICg/cgxiRFAUX4vWV40hqg3DamWSqOd8xgseOZQR
qetajrkhjU/mpPwz6dNYVcCCht6xP0yLbjnUvjo6kYAVmdBaIO1Xus73vm9hrraD
YLcRSq2isR1WAZbCUc7I+zhDHS1G+k3gNQR/WhO+785pm/L62TZi8UBPss6T9d8I
f+ImDLrg+UA2eyykG5H8BLk3l9pGY5X9570XET2KBIA=
`protect END_PROTECTED
