`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ODb7n18LGMT8f2Z6h3uZ8fvv2/tFU3MTNYIlLRl+OwGTQAKMFM8Zg0hNoqWRE2Mj
2kEGIiX1A53W5vtFon/016xT6XunMRYPH/Af6IDkAHEg5v90hpXL7jdjtU/eHD78
8zO0gsW8LUCNb8vCKhnPXKrgzJk7IPh9hFltMf+U8DrMNsjtbfdLNOT0JD61S1t9
CdVE9LZm0AHZABXoiFvd9oehbr0YGF2xLFdiOwNcU9jMEuT1spq7iOrY4vDjuWkC
2AJRVrWfl9/jyzS1GTQtVjKda2tkQ6WNL6MkVGE1BbltbV3p1N3RIvEMUojfBdvl
WHm9DQPzfaND3eQX8Gw8WZJ2p35v9+x3BZoMy9UYxV8z5YoYrvvLsQUf0TxHvBF0
GIgHxjQUrZa8zoHETIKVijCLPlapkVpZ1bkpGjOMCGAdC2LM5YbTOM+on6r83M8t
B/HufGy2uJCnJyl5SBTBlqyfP6E42K8HYrXbGs5wCOpf8gbdfVEq52xIk66GdVMU
KOwEcpaob2aeBlAO707J1UvcZZF5BrU+AbOUTa6nYAd2gGBDiYPUC8wlS3IBoQjM
F/lI9OjUXLz/QEZ+STTzGEeHaZdPljsLqb3IvyeC/UCZixSMKOFkqurwYuP54keU
HMbeyqqMO3UR2rR/MCcuAwYBAe4oN4gwdvWcaxxCP0ZSe3SW5AmKzufqCAFslOjm
/YHjnRDtT5shje6kdFV/nqBpP2e+FbLWigFqMPRJJcNnUeS6yg3oPDhF5KvkrMl1
rNdvm4i9Dn82wXLIt+JpIzJMB1woPzrwBsExnufMkraiEtbAR6lBQJhTw0gTldxd
H7gltqdTnSI57RonduhzmzvHCQ78vq/XWC+O9ds4N51XFUt8N6ms3/Cv4ML2pT5/
GOrO++qHa1TjWig6px9E+VBF2dIRGE8ihkJuVwJfrijRMDem9yqzGi/axgRcySJy
vX6FcAkdde8ug/SFR2IuIno/Vf2kxVQTaNKHcW9Q+1j0CpEQFe6nDx16iuu4fMnH
RVFvXvkBxCwIfV07haVEyizGm0LqlECbTR5DLUl/coszSdj/D5frOQ7Ze3Wy6mG0
iaQlROx6se/e/MzBsFbmsojsAeboIoHoEGQnuPww5a+xtqyvFE7Oznz8bQ97PRat
tIjUaEMEyOOwAF/esfOHlYai56UUMdlbeFa1H8ngH29yaAI78/6auaEbmMR9zrqN
+L8wP+2LrriQhByt+Z7NR+9CmCquNpjWI8XtPRyPxqM=
`protect END_PROTECTED
