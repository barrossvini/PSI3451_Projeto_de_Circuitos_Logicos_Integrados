`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wNlzNdmvY1baFSQZZxYmOkly4nxiwociBzIjujv/SrJ5KWRqNVhJon0p4CrijKPu
LlE9Y+otoXTIz/KE1GYfPpti1h9iU4avCN8v2/2Bsx6eBHTXV7FzM1F6PX8rLa2P
eP5MISPAJWKzB4YkPV6pE7ewoKAFTKRdaukZPifW3gm92ugF/tmjLJQJsdj/OiHk
3wt77oJcwboGLxyKlb75zMh5PffvGXIxYNYxhluwsT70iSAGHfG2fDeyjQ17zQ4T
Tn7D6wESYWSZ2IdCEexnAX4DeBS5FzYYpzYrF1k8HLA4HzADacZALTNGQ1MxFGxW
tHwNYVzOGAXeDq35HJCOyn9yuS/ClST7/oDwvIQsA2IZVI1l6k0SpX3ZI0tBWsMb
fnDkQgTxlWZ3VocXV/BeZ5yafcw9inKuiZmzq46HRpqPB710BaMQAeozpiDbRHXk
eiqRQ5cYZVtKEMdSy/4n+XVpJKUbOwuX0IKTSkVTuTzllokniGRhJgNY3ZO7vl9X
gYIo4ki0vNL79k5VDHsFkuzt1JqVtu/Cvv6UgkUclivpy8cF8myzz7B6GWL0a7a9
/sdZRjhWpvC79yj6BHAtnEPXUALYTWhCK6YE3TiaPPTCOHAdcy7G84oLq0UGGPj8
MX1q7aFvAZ2FXFBdarIsQ7we/xKVQ8pz14RgZsiJCO9PvVxQ3cwVeBP1d/RoXaMz
p6NUusYD/bAyvPozMQeK7GU6m/p72j25OobODBLHJTXcwTGlP15Z8B41ezJ2OH2e
cMIpsFu8POpJ6TzzKwI63Q==
`protect END_PROTECTED
