`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3fHtk7C1K+PUAY2n+vfsU3TNCIHfzoP3iuG4i8MEJoceKFh6LSKCQkwApAODnqZf
4hn0Ex/B5AUTyIqaJctmIVkDdRDL6F8HIi0B2w7sb8VF0u9BvCJZYfkTJ50l10Sc
zs9Ym62zQOaL4KozR11Nn70NwG0Bp75NvBCsaIMpkKFnfsbj9uaZCsm/Yh34BkzT
AZtH0/suzedVg8QhdYcseBtZKLYj/I04dJJx5xf9uzNkBrv+HOrQIzaouPxONiHD
OSX2YzBdN6/byJnGyG3kkM7B8bS+RKpHniT8XhUtb2P166ZGLI4ncePnrB7HooPK
1bxELlCj2DCH/ga9l66Zyf4l4BJO5f3qAl586Y+byPPjiEf4zHN7tiMannVNw/RR
pSlfWk/0ZJOaAkUpQ24rwGDl9CvdIFNiEYbT9tdcNEfe8Xdpeb1W51rsG7QxtwnT
vYQLEMFbREngpWp8jSvxbuZqNLycN+sfmE8KRIUXUyyj8ZlV32+QPi5zSDfD5hlK
o/VmHVJhSm6iMfJ4sxKcJyoEKzFDxS13Qog0r9k7bzIG/Hkcf/zo6UhDjzSU5YV7
l/i0azabJrDZ3UgQVty7sIy/UWp6nTdI7WaMUS82TK9NvldEEoJaNc+/O+O+7m0g
tVYUR1XAe+MKPT/amr2LAqXzKXFXIi0KMWmNvIows6wxu+l1xIEOEiHCNz2oUb8D
YVE1qaAp9JTelk40coiehzrJE/aTUmdpVgQShg4QjPw=
`protect END_PROTECTED
