`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kd84RUTgTKaanKaYBLrWcfApa/b3Ee/dal1d1sVo+RxRCZ6M6A+QdKnzW94E9BbF
407Nod7NTp83MxJgqZXblfCgihd7OvTAeLzyR3l+VESAMlr5/wqOVhCU1iIvk099
NoS+UZs+CEjELOhig/jcJW4Ft7ZPTXR3+ay3y0FO3p86qvVR4WOrC40N4I481Zpb
dXhmzpvsnSN5LNrn1UNSbNfQdUScW8/0DMq6Ed3eskgAHMmHTDqolAV/RbQWA0oG
AWMgeS063Pn/+MIuM1ZyA0rUCu0sCwGmV2BQxee4Fjf0TIMMXGbBDKLIusBRH4ZN
hL+p9kYRRRTAnKnuLnrYQovVIOgL5MCteDMoa0C/EY0A/GMCM4fzkWbxmULd+eNC
0YyL0tPwTogP08j1RO74e3X51IXyjRrqLeAv2qrjD1rPl5sXgS0XJNOzIWw5DpDB
ycrVVecgfkcjOtGYNgbPaqqKlE7snDX50tO2c/drNn6S1zFX/+BJUTDR4BthG7fc
iXvVikkW8/x/C0INn+ZUDrVf2NBFLth7+MgJpejJBzoIOp1pXTA+vfTzYlLJ+nMs
1q9zNFEr0gqfQcs4sqWiHHuEqNbqDFI+bX2hbfY0RiUxq8wj47VOy+rCSIkP6SqD
hxQAvXe606pebX5Wm5444XiSS1d8i4KZ6F/4r0htmSpmz8/kAN00Rv6TrjUPjVvh
tmia3u7pwpioTA/CzWVEb/QJwvSbdw0za2vdhHJ5PNIw1SVvBTBF+8NcQOunuKun
zY96jZQLBeWzRvzQJ+pgeVjo+3ygKAIcvsDhI+V2b98fL0WtWkGC7WMszp781UUh
ExdnYGNDFRAFXPbUzB0ZD88+W9IpUEHBKZuuFr+QWlXxiEmD2otiKLbPdlCg+fga
YoxtCVOfcLVyCvJbmJ+QwpjYh5HRRUGHbcBvdKAypvZSEWzvxWx+CaoBH68CFtmA
9jI7tjAxj6WiuM6V2CO7I3SkYkmsCWFirI8W5mQePzPCmxMeRbXEmR6ytTyDORHE
77pL5LvLswbyumRqamj4kfPp0cUCTJaYXfMX5QTiFZQ20Vr8tOrgf1/urE0ubgV/
11f82mKjcBFdzIzsASSQdg4EfXE6J93Hkfvr5bcVIwytPy8h2i3j5xomDLfUY4TN
UQ8PaZlPSdlm23K9O7gq8Rt1s/O1d+bMyw3HAZvIPh5ok5t53y1ikpCYJkqsS3Mw
yG7G2chjlBfxfWOMaLHoHACh7tSyzm+KPDmRZN3P/aZcZSjgIc1luSTYNHG6/o4q
5vNsrMdcrM3o8Slmpta+hrN4b1hwrwfcIIOtJS3dw/QehR0skMW7Q2JE1vk3FDrd
Q0tDdqeBDQE1hvXQEEtsDBdwy4Wt2zAk31S+YCOHZwltw1vKgyaq1o5kiLZfREvD
7WvOTrNMlaRcMtFvES+XjWGhExNB9vYtrwH89JStKZlMTHpo37ZpZIW2DtcjcnsK
Qai8bjPz6BY0f6fZiNy5VWXoOtM8/x/6PUbUiAa0c5w=
`protect END_PROTECTED
