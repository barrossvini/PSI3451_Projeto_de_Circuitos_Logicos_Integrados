`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mfV8R1Nyhh2o24A4mvcn0/nbHZz8zEKFwceiHy4wzeGqtuzemj2QQ9BGZZKGYYN0
ujhFUV1WEGCJ7BzlQPe6PBpvhAow1noWbL4JdwazKXNwZdIpaL1KA4BCuJI7OxMj
+Csu86ry2Tvs6XHGRxMTT5mIlfyokbMwoV135i4fXUzmjATWFMjPwy4pKrqcQjz8
tONo4OlcJ9Dij++vsgnVOT8Lvk1XgMa9OOQJzD6/lxmSR0dvHdS7PNcWAefV+Zb/
DpjgMxUeNtkhT9CSIQBqetLsfhdnva/a7ERiGV7L3xGQ52/LCf4Q3AG4owsOKPjg
fCxTSknnhLdzhdeRTt31e041slqSjklpSlyJxb9pxMBq+Pi38dkDJ8K4z5vcFTaI
Dc1n3B1IlIV9v4nY5BTVmucN/GFRVtV7DtUQNpGsQQPdIHQsYU1xHHT+F08jxyNY
hZdwHcAfCnAhAQwtAqZx+AFViHzJPGkSKDN8k8g8pZHvZt8o+b9Vj3uc95quCvMI
8lKYwN4XIpag8Gv7J+zi/qsuuWMyGEynABLLOSbEnIBLz42WV9KPUGyg6ORE6OwJ
ZgW8GqrZa3X9iRjLpB1qVFXu0wy11W/ppdoIby2IZoDl3QEtrp+T9mnSRiGI14uJ
IaAD2DP8WLz4AZwBJMUksGqlK9RpkvBqwiWm0q3B23jA1V3erwv7te+77CFunvyM
qM0dE8JoSIME1XBoPzO8RgXsSWKTy+zn3sFdJljFSTar0RJYwgi6Jz4T8yubO2PH
dk7p4VDIbO+KScvTVZS7o3Pm1VNN1knpZMNnIXfz5BgjZI8aFrDVjFq4+YNqIacU
Qv1IJamoGDQLuhWZqba7lgkNP9HJIUbIHxV2oheWmls3ObpFRu1MBRnEiibzIk5J
I66ertITloYw7rAM5RKvlOFrXacbr1mxOcFy6sODCtw8UM2OKwhPhX3hbRTcnvl7
GRNyCeHlU3w8xmVPDg2b3fHm1F10Rsxm7KwR2G+z8GuJc61wyoairNH3oHRFDH76
+6WB2pzlz2mGZuLTAUiO508eMcLhG/Z6Pt8v2SNNu/vOdEuK0EB5V3QZbV2WOtQ/
O8W9hMUDBRLvkjWD2M45PPNjy1x0jlbC7FFXNZrZMd2AEUr1/2PJ/jqUXn9uSqYY
Vp6I94fI02MSfToJHmsnaBNrYDB6StCQ8Nu593eR7EdH9F8CDHK1CX8UutZgbR5s
exY6czcXTnKtp6h5lHxVPMh8+SUrQ9X0AAuSPkBArPgb6gQF1IsEmalJ4Qc8m+6k
`protect END_PROTECTED
