`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/bOT+WkBXTbu/6EKt/c85dg2ToQKBCqk+l3uoNLpq2z+yj63rStuf2D6Kn/xqZP
84rKUF/yZ5AK9b72YDodZWiZR6nzImdYmnx/iWIKfOmMKNPugefpTcnuruzKeWri
SPJbe7x3VeShGBtNJ9tPOtkB4K9Utnkcy5KhIc5af4nyju/TcgQVzLg8FXjKCKjq
d6YWTn4pXa0TjtWrtYMm7/nexy1iLg7Ow1ygdYvwRLN1564C/PAH49ranJ8ZD21S
iFFbs6gR2trhTmwTxzr3uS0ycPSHhAW6KMKVnYq7zxB9oHCgKTXt9OxD1n708oZ6
4hv8QdICijKu2z8SQt3TCufIMHdSzWmB9Llp2IBzClYfQMVR2s3ZIm/TolgO6PwI
Um5kt+uEitb1EhsdpeWxB2hCSCErd1HA12AKAwRqGySN8edhdr28XrwKhirPdtoS
sAsaXUyZ438uENa68h4KVPKvsu+npAOPepvHrc0xFYslvwk862z5nBnJ4bdLWl2H
xcIXE0iDjI1xmPozPxc/Ns+ntbK8FpuG1UE2suLnmgZHRYFASRtQQAna7UVjeNHI
LZlpoq8qHR9WO4MrhAfyox0eReLuoIaszuXIrB77KlQxBzbU4jbCXLPCQZwqzfLb
PC0P0cNtrD0I9eEHgdN2O7Q5ctLUsbk7BGEQg4iIpbmokmobD2xbc2g8bAUPlB0h
zSdpaQlQzaneQUDmf7BzPW3NgylsiG9PjPo3MXQ8nEA=
`protect END_PROTECTED
