`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PGNn5KB29Q0vNhvdt0JSProGChvMHglA42r0zwT6TShj5fP308e1UI+KBrmhnR7b
Uo3xOFk5BDxBdtYQ8s2OghQP4gCrVkFhyxuliO4N2MNpici2OCRJCQBknNB50CYT
2cdrTC/R8o2urGJktjgqbsKg4lLh4T/0fz6xgRFz9p1Ulw7r3QSPQlaYuDPzRbNM
SELNFVZImTD4K7/uQsnEtY3vEqJEfyqFo54sm3v5vBa74Vi/qu9KHhwls19l9GuF
+mMPngnxwt8Z+xwkWFXck7PEDt4+w4rh0QqzrQElVTyn/j7+fI/bGh96mfEo3EOr
/zCntxztXdfcl6fUDBFTliI41KShZ0IM5GbcNcidzAyBBV1n0IzrJwV+Qc5KHcmw
iefwDrsrhP6R9jJwiW/ze7QyIxsY11TLw8tRK5LMu/gN1no757zc0wZQWRMg2rf5
fGeVVbDDTFRuQpb0vVgM7dAozOXzw5eUi4lNA5ZkdVt91Ma9n8KpwZzNEi6t7CxA
OsvrsnU9rN0+GkXj7vjpr+Z6K5tZKzuz1Lf+E/Guh7wSbU9uluQyHXFJ1KPzZWw6
rjqAaxl808iv89gE/hX0Bs4DBFZJYi3SDk6ZkhgLw0GqE8f6rRegwFBDgRQ5ib4s
u4Xih/p8qcuA7RIT33BAwMdFl4v13FE4+P/p+9xwoFCn1mole38sqJUWg27eUOiQ
maQ1pDIn4ttzwWH18UXBsB9VPCE+rU3KjnQV9GQoEWBVM2+ihf9F6njS9LW0WaI8
0EpVILKlXzac3759LfScnBkC9l2kfTQrSPU8rfk2MVwA69XE5uKIffwN3p7FtpoF
hMC6XHnmYc4g9UULi79eFYZGSRkA7BGIzWWAHSnoDpR15eHaPM1yUcPd4IUjy/CK
kZr6hQC84ADE7yYc+KiRFHJr+hvF5fyTdss89GE14/OurK3I00uZBunhAiJ5uVsC
l/BMuXu2Xa7nt4HIAIQ5SRz4TUb7CLh1mmmDGkjDKvpLkBUqcVVC0lLHaA0u4E5n
E6AvBJfSTooeb+6MwRR/mzxGVVdtxucoJQ1rKyVmX622AqApjYeAGlDzb0aNZnaE
nWSwyqcIN686pyx81gsPtFztl1JIqj7riocOL2GpCL9lDCGfrVDwNuPBkuoj0CeM
ivqVRZmNhvkl+v1GS/0jbHGtj6+DqwrMV+DQyIFi/dtHjIUDviTMehHcziwCLd26
+kaNuskdFEV5PromsEvUk3nwO/FO47kR5QzqIP/C4PfhO1+Bg76zLhFliL94G0P0
N7ozL1xWfigL0qTm+txva7FIeKFMtNzOjB0Q3bn7cuLsvzeowhpt+Q+eeqjvQvvG
rKHFAXygn4h5h3VBn3R8mBcnNc0lNAoHjFnFDLE1Px9Hy2KaQMsVVfIHBcmr1fx/
ZziT5rvW/1S+rKtE2aZdsriVVNRvZ8AcEBGbS32oN4CQ9NUk4MdrHVK44uzvkPSq
viC/vKSGYXvV03Bzdiv50n4VIE3Xa7ib/whzWJ9LAGx7syUUcCNaZVbbecooELxP
2nMQ/elS9oBvuZ2l9UruWUgk3keHRS9BVtNpVNj8ACUdS6UBQY3Cx00jT7HOQmmq
W8kG4DJdIyObM9FMe9VQ93SpE33slrUAourta1nHnKrdKKMqqLih+uHdgbEYJDCn
+96eyG/44eg+Kt8TKdusrudMwSdT7ZAa3qeoPOJ9XJKv9qoKPbNg730crkJKWe6q
8UM6Tq0QLHpaqqitTgVLdKFRwyMMD8AH7zYmgILZvU0taamgIlNN+XkOpSYyjIMG
SCi1vi3RcEG9jLmV1pT60p0tVmDUrPYNIJzt5fQwAOeuRk2gRrotmp4FZy9ml8BR
nbBOzZfPi5TVduNSIgLKE+2zymEYe7aLHgCDSEb3HPxawAO1LpaJxRYXXIrtpmgQ
qMOvglCb6BTfRxFvJeN8hhV3TRHyBnYgbFKopuoCsMUL5uSJUMdGUYB088MYDDao
ITKOazx/UVTNt5P08g7v/joDv8Chd/GPISAMfoKQcb366sI/Z8NMXYsRf194jQW1
EhOVDBLrPKmEi+7ZFJEIax+A7dzqx5F6CBoT2hXuhWMDHp2zRQGiOduomF9nu+dH
tRjdoc9IJXbr3b4W6oEqzVVGXl1cXzyEa4vgUEZQI/0p5+lCt23wGXxtJD2MN85o
4x4mciQolRfIBJ+ikLTbvwaYezfz/eNNuFOSY1xnisQCdxB6BrBMlQmyZXTqozVX
kotp+4Fk9eZcch9fE8v+iKYc5YcSOUpldfv5EfpsXB4s1UOLdF0lCvqIsN39Otij
42iO8OPuL6hY74gxDbprw+GAtyeMcJFAI4EbzxSRbS3l/Nd6WnkG3vPU/eLydORc
Dwau38i/OmGH7tOWsyuU7kg4cfHEku59LSKmJeE6zB6xFjR74v2A9RAwK60ExFC3
gFf2QsOFAhper70mjKhP/h2hPL2VCcnyuOkRnHHe1p3xQzyzQPH4awc+2+9YP34F
inbNP9DmD8FOAWdlVS4oXBkM+DdcchFTBKhuQOQEZzq1+EmIuREdpnn213ruO8Z3
A3Rp+QE21tBABOkjUCpJttZJ01OIN6F8fXuiVOb7GdZdWDQ+dQkIKvm3ZK/ApfoF
27s5k1AyPQWIwwr1msYE5j3yBaygSPxiAaoec5jN5wpc+cIWy9XoBBx2LeMbjX2x
YaBQkpU9Y7AyTZvXiDLVm5FuiHy84nhe1VkMffShEWAgy6en326NpRw3xoXjJjwx
kZa4g4omIDYAKbA//R/SjMfc75ysQUzpCi972WMMJughEXZ45jgIzR9M3G0h0ReH
oAH/JpNmImhhkBJ+jakkoCFFMlIc/MCfBo5H5/acw2qezGdOseNiieBGsD1n0c70
ilV0sBicUOOyTgrk5AzvC/QITYXrvwe76c0t+HrmzzvWtZ3ouja2dbIikJN/qevD
ZOEq3m5O/bJ9HkUPMmwhtjqMJzH1k73peQ1XTDmSWhz16i9WzyRLL040OIJR6Y1s
UaTKX5mltdIKjoYsjHUh5P9PbIOH2WpgePGHjOQ6tdImiAvLBA1azmEHt6mnyv7Z
EtPOHYgE7Gobvao83PZzVB8dhgomL21rjthvJDoInsS7X+G6SU0acK1UlrVtNX7j
tXm8dP50ZSRD3GydZ3ceO7FK5Vl3cVcwHLYzvX5aLwt7Od14G3GftO9s98sW8MO6
F9JEqFoKpcrt7z9YU2PctuNRvN96DuMrKG8S194UVFsW0M8mxF0crLfp5xRsoKEz
DB4T4op6vDh6n8fpcHSVJw9aI9f/FyEKZl1bUJFwtUPAlHRRxkT0b8aoik03b7pT
kSvQYvX0GjCMs0YtqPdivtybaY5j150EWbaCsuihV7StpxFFyQXpOhSdQiIAwIE8
rj8Mt9iKTdok3m9e/QIhfpQG+eaLoEyTreE9ArwEXb+4YYkBd8dDVfCEvQJ/d3Mt
VukDdAk2/s2AHTS+XschUjEKPHc5zvuwgsxpLloBsNWHmXzLpO2nCB1Gm11Jc2Cu
cZDtq8kKN0dCKSsbMz0hdSj7P+pIRFtpNKNOCzOi7gBdB//op9rmzu1V5VgTqjgG
USS3rGxVRuAmrlw84rIipEm/dOYJmU4Q5lYZOSaytWfAXJ7fVqxB53oFRemWU6cE
gM+nMaRxvrs8XUYCIZgowA5iNy6hbD34sVRkl2iI2KyjGSJt9nkKtXszIj8V8iDz
aM1gS2LX2Thtmts0oXB/5ncT7jRDSFEOfaYcLJWKhO4YuKhFC46TINw8xAF5bR8y
zWe3lXFy9/I2zlMbRfbVIQJzQLLxvIqhAo3IsHp/DJtIuMpoYwRyge2sKBehf6m+
3M+EZaLngpxiLNVG90JhURBOq7SOyHSBrZJFwqkWFIzIX/JqQ0AsgtKVpCuCVzQ0
mdZMHdkiKJVvNRl7o0+AJQZ+EEtJUO+3cVP+EEko9nVQUKp4VOfuekYTGZMP7w8X
unSaS0Cw1XkntaGBPwFOYPDpCfvNTUpn3q6j+X2RfREEhSqVQlcI0pOlUrXas0Kk
bw/n7ZE/qNjMH1XkPY7fZ+tui29qBEcWPGFHEvOle0DLS96rOjoASeflVQsXdpiH
IicW90tCIs1a5keXLjg5gWk7VKdjcw7sISZTub7k5RT8eG2iHfdRzHi1jJhBq6/o
xyk+4DhPpLN537AHQId1qzXpyRlfcrmo1jqakJrNtx4VCTdWu+HRZO0iypAGOX6Y
qCayZgoY2F2Mdih32St325bel8Dr3D7eIcBh9hbtM2MuguFFWknss7ArrgAS973l
kwECMp50TMXvysQFsRi7C3NVknlQWq6xFBEdo3BET6KEoFJlnC9BgIgEDYSZ35Sj
/55+8gmTTHtB7vQehLNE6ZZHPpIgZ/HLiFvxKbGRrCLkgD7lLa8Mxu5Juz2ggpCR
wopddiGS3eIh2nJSpO2b8YDqI6IoLiHatENOLf709jjBgUv5dhcJedm4hhbElAdF
sEMgcOXgkqvl9+Y6vJL7Yez5VDVy6iKVlISV1nmPIKeLXrOG+61gT3BxIvEGYNZ9
Th8SOtpNeUaUEfUF8b4ww50vhZqir8OXGRjM0BrTST0Rd68qn8UGQCmt7XdxXkPs
XrPuEPHE0UTN0ZkdO6vVebmWonxLvTIF8g6PKlO6jFexZz+65cCtTD4TZwRl+Vo9
E1f30uc9/jd13lHyJL8NMLGqPOaLtFSii2SCe63SyQQ2AJaejw2rB0LALj71Ulr9
BIRUKPDOeZnPVL/n+DSjyWV/eb0CmtOUCc7EJrrZ2vmEkEl5sv8QgDeKO1yTkJOU
WAPcOOpjW6iVHKajLL0/S8wpyNryOwMSwW9LOXXQ8E5Bi+4FFhGJe+s3Zp1kmWJp
ebvE2y3UTEla9LrhIpWymUHYUGiq3kHS4FdxnSb66SzfvyhV+6WvFbcYQUqPaWhr
AaQsc612hRbFxKanVhTEt7+b9OKXeHCz8fY1HJVvRoB+szHlPvMenT1gIb+SGhTG
RXBz8spgRz+ahKdv/zqQQJJ+wFBh4xt6qUbNgePxZhsO80dPrdom6sJrWGwZauoV
R7Y3nm7OYFPCZkKxOSsOKA==
`protect END_PROTECTED
