`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hPHODA7Xw8xSylC89xGzlQEz96b0j2NYRLHRqQISjCcS5ixO+RkLW2QFRDPY7Kpv
IO7W9KUx+fRs0MP59MNwH7yFliotvbPge2nobVqCNP2QOdYLbV2ZEgYKT9Assl8C
Mo7iTTFR0X2cO60Hbc+cDo9pYptZAT4UL+ISl0ga3KCeRlvXmAS0/Z9Dn3KbZAS+
192Gwc/hmBq57R5CxTmUmmHW309sicMQJM0DqBafl6DwPzPJAIBAGTKXcHAazdLC
rA8d1saqTQKhGZY03RW5oRaM5lodN+8aGStoCSoP1V6PIz5FlZmpO6PhN1wPLjpr
0xbGyim48jC0lQBQtkW0s0qN9uM6BfLRQLnLcNwMBs+LpzbqLxwqj2Z3Mephm+jj
wqfOtxZvSMTgUdxSpu9F5DeljPAQjy8eRAeyhOa5LWexU4yjnYeegfAVBMO96In5
eWi1L8ZmophupaYmkU/tc0GqtbU2P4ctyxgC2UPutRVmL/tRhoFXHmcwLzIjQ4Qa
BiYvYpi0f0Ag4bM2P7TIEqEgqvDK/wihFXrc4jVp8ttmc2lPoXPXS6gq5Tpj3CUu
22Sjwg6U5zqv3G7ChO2bjE+A/VTNPMEPhPvkIw3XlztlmlkgAQ/Gi19EL0wDrKoo
Cfc7DivyX083dfv14RKAlzlAreLrYNXYcqyzuC9GK2/n2lfJp+v2kmaWjcIVfOoM
9w6G91RCOEvQD6rfquUQpqmm5HHX2PG+qHy/GSTaLIY2WTwq9OhuxB6Jzl3jWbXq
XQ3gm+dFIaAAzQrI9Al3jIvB8zgDNF2+/V4dwP1dJR6EEYRpy2bhfZ3GQVuvqmUp
/QReap9S4L0VQcVOWpZWMuTqFMEyBExRfzUUh2JEPRcQzxYtkg5akmXqaNYB31lb
pfo2nnVeACvguUW3n7Bl11ebw1bf8x7nAh1OEcEh34wCAStmvzPRjS/PHad1VjSl
cQetc5dR9PJ9Lr1dtjRc/Cp4zRQezxOqHUnnbgS/67tHJFDkd58BBPy4NYQ0z65E
6nbseqamNgYwu6Bv/Vui6xt63K7p793P8oMJB3IGAw/+s76i6FX9iyGKyyfhy8Mi
LIwOxvD17//dTS+OCLmxkrAXZPgzJDEd4bs0NwfCJG06042V5jsjGgVouhGEpzgh
YCnY3r6xGtoP5AtYF8R1ICd1Y8+cS12ZffFIyuLxlVf2/l9B3bzzAR5b704TIqCd
wuxoJNMGpU2WyLCp/8RT+CYkNEQdrPPsfCdqFl1VOpWvj8J23CXZVthyf1585M5U
`protect END_PROTECTED
