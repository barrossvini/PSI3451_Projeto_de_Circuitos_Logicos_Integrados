`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xxro/xxBp77WZLst2whbXMIAgyLzeowuDR5ZFnIMbLqiaVwEUCyNMjdRfm/gZ1Vh
57wr0wAjW4mI56kAoxKdKk8Y7Fw1g7HjJyAt9cDRem8UOQnIwda6lSug99gKe2yp
2uL66NsBpm0IWfY88nGlmORQaRi+1HrQ+XUqkw3ZLTGwLUTZ1YGkS3DIgli1+RDu
p/qBGy8zuEIB1yddhPAHZJwLpF5AwpZJf6Lqy6mcIz5u1ojbMDk3r0NlAzMZiz7j
8mA8YnxG6lfLoU2NsaktP+642e8NWSd9FFgy9YFuFFVoTxHowpyZrfU9wTQ1UqWL
SywcW9n/k4C6iPLuzfZmS19Ql31a6lQ8G9GA/zig1ySHcfGJNIwlHYfVQT+BszBl
ZhZuFf/Xpcn/TwumMBMJhbvwwxF386oUhpU3C65JUcyWXBLz9oEzD3IcoX+bdXks
I6qRQeMXggO8Jb0jRbWbBE647WWTZQE/LK4dwahHXv9scr3X6V71hCG8kOU1XbAt
mf1Zl43KXdGzz4J7eYTBx9fHLMXBEmEuQXxYFVpfrGyXBySeBzb+xmbEr/wsJWbY
ofXFp7lchEL9fNIH6731PkBYhaXyc7yGQUZCJ2JRLhiksY20IHUkRNB6mWUam7e7
hLEkldIcz3IP/HqSaDbeu1QcguaFPP+2czMH+2rejl07M2srwF9UxcVfz5pyLibJ
XMmimKN9db0JSF2/uQVkawBzhPNHULVK+/9tSvoz8zGsrgGXrE0nQ3TD1GqmA98S
eFRggZkD8JRoOcvcMi3sATaR3atWrGCJA26lhbaDg3+EqEkIgk5Nkbj5gW5+D1xG
VIiQlB4qdO4Xa4lM/5jpky1JuL02h5xRr6jM7AuVt7IWKxz8ucrhFI1CwPZvZzHh
/tGdHfSuZ2cxFTfr6+7LGfJt7XT6fDmUGxnRd3HRWBNoywyl3C77WR+qfyu37T82
SOP43ln5H1lon68XDcRGqduua3izbx0sgtmwxK8E2DkFh5rvWMBLvZfH2WrhjZeq
LbJ5COoWllUW9WQjVEJjK+xPDZRqsquvMVcNeqHNNglWnTxcBuFKuz/3mBtup14d
vPtSswKIC3J2trXOCIj0/3/DnzRXTCwDqpXRn2N+StQzcijGpR6bCInYc9W2KnSZ
TcLNPy3hKqD/nHT+aa2QY5tCfu4KoBadUMZsCNFH+8oMoYaqCiWPzjuK6RYILiNh
MmXSCrnFLL8+5OScgJGO1b6kubCc81S72/9wb9J4qcd3N0jJP/2onEMp0PzUXzxC
UPzzXHd3iqBUK8qhF3lY/vMBWvsffibYkVTD8g225L6C7rejV2tkUou1Bx3hueqe
yMHIWxFXwXpyArU1yylur4NO0CVIQXQ9Teh4REzm6gC62QRI4piCRzRNDJWWOf+c
MuvjgBqHn4N8HSS2C9z5wNNVgb1oZGFTOPoPro5uzdBv7UsxKw5e0B+OkagzCjDn
hcQGwBvZKE4QKfqtcYTJ9yJee+F5oPMFuGAuRWruNXfYIuyj42GRczah7+DvXWLn
kiT+F5q7bvDn7/a+b5Um2dkPZlrtTaZmqGUgKA2w4M/BmFd43DweguTW0u+qshuo
dsK1xDDJffaGBuTx6fvNbo0JNoPhOk5E/LjOdrvbE+bgRo5GGmoRFomRfz8Gd9Q7
9D4aaFekrgeXCg/6P+EqN2/3fUQpMWu0a3C+tRjirMDsjI+JegJ4kgNxtF1bTzVD
`protect END_PROTECTED
