`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dEjWveWx5jHczILnaYiK/8aBS53LEQLXPQtaNDdP3KjkjiiCU0WjGqNEtt1DfrMK
JXQ+/fZb6BoqoNTpV4/kmPoTuEnqQTWokwmIX6CLSxovmPjBxwXMM1qlVjAZ5SiK
wmCrR2IxiTs79D8dA3cMms07xvxMT8zkeIzzmoEcRDoVglztWPUdpDuKRIOyVwN0
G/GJ7grTT6QiF+5eyiSJ4oTpWgdbFnvVayj4JGy0+5c9iRJvP2/QQf85oporbHuh
aaKEMTFWUeybaRTDpNDeX129EEnN5uCWwU89vDnPFQJZ5JUbiOPVGEQWY/SfgMyt
z1UJ8s6+kJNz5w6UL0e9MtXbw2EjgU+5w2X7su36UZyN98jlXZuETf+ibCdh8y4R
5HsMOrw2yepKwGJis79KrZ7Xf3xqk/nV9kZzvtmErpY1fys2twrWUa9WIp8LOt+z
VOxwkp6suX062LIiBJhNCxZmUG/jwi6OK2PDs7zU2Mrcz4597V44VXHtqmc6KMfN
K6tZCtoroF6VnM4/Eu861VOwZL2HBB1gjFzbUeGGautyEk/UilM0utel9XSqn3XO
NEO+H178ziGdoXBPwRVU6OUFX0Gm/QvcO7wgCOrI3cMqCCufGUVTNsV4PkxLxts+
aJubLZpip1CcLNZKIHyJWzZguQhh9hhaBi8YM0hHzd8ThtcWy+BCQOKEezZpzbnk
1XQ4IQT+Mm2/fHBOEDqeIULLBn+VDGzg8GliWc8IsNxMuC5pBkgb/F9wkM703wI0
`protect END_PROTECTED
