`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gnOJ+IEP5d1TWWQNrujNPX2Xubo54rpu68q01AD3f9gPppSWcqwFWoLXiFT0cSfG
6MzowCY3loVwtqTQ1v2WPMCMjwBoDYi3yb0btpTlBGDQc6SckCCn+89yfgxwRU/Y
VaIagasI6WD5vNUYS9t3LmK1S4GvzAiY3ISIC7lxYheobpWh+pQkY0bocvgE1MQN
cceUztBNqnWIzzJEqhXp5fkY89Vw5WvdIrbfiSkadpQ8oezE69SIjFsA8H6fZ3vt
dDdwX/oTLYeYvM2Gb6bS33KNaVurepesBQvwBZfjSOSh2jnlrr5lrlgYJrow/0Ad
qLrvifUvN06um0I2qVYYI2XS1NugoGrwmlylC0M8AyhxE0n9wAVXI0WzKBGonzVD
yEM/wwLWRLKivreDjcM/gSP6M4RIQbR/I5wY/Q0tvtDShlOvYDREkF+um8+qTld4
yXG2hzOE+N8ywQy7hBcz78x4/6XputnZeSE+z1L3aXpyYYlB3tHNzrzXqL9Th4Ke
bYmjH3nvycov3Sx5GfzVzlRoHkEpGU7Xt7UDgzv2FIyUtZ59yUks0p0U0Oguscl+
6De10NB97XBTPDtLn+5eOwvp1PZxxx5H80gh6uWXCzHCWB13MOfegx3W8XecCF1O
CchByTegQRLl23ZzCARyYyvQcEVAXnwjhQQTeM8ZuktAD3QyNlv0duXpV+ERAMUe
STzfclfs5heQJNnqNOqv79L6PK2UnRU2OY9eieFsW16eIJ6NpwPaJJW3uLf11o76
97cUT0I4OfeZ3EVZEskQUQrB14SGMT49Jxt7fyLCLAPQA0VTmXiG+Q3JUHlhfVon
pHi8ZIO5CP4NdLhUhJh+gAP8ciXpdIMwEuqWm0wJLbKxKNFXjw0HJXX+Xva4J8fA
HzrAj51UkWxwSfRlee10ioRiazvJufvfLHN7AI+xv7eojMG0UmfxRxyZx0/66s9y
wqB5GV690qdtVTu7en206cQPTZgQ/XmxqW/yioIS91/mOjY1b6PJE0YPb8rsQIoa
oOAAhxDzS+PYGZI38UAT2gEDGg2FEfgqBrsm7h4A2c2kxSFuBhdle+igJOfpgG1r
9w1NdJBQMYKXAui68SnNLI1TGLLPX1R784OEjpFxCLNOIhJriOHOyhnUyR6j9AUT
HGq9d/QNkDYcK+K5MxGSe7u7KSQVMGg0DajX9aKJWahpaRMpfO+g9aSEoT74avNO
rSDHDaPAAepaRMVrNFI6JNI0tgjDwDMLiCV2fBAkwjGGvsTKt9/9rDOU3imK7th/
`protect END_PROTECTED
