`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4HJnGhwv9ogqYUcmH3UT4tj1+nNPt6bC2n1fnq68jW4IAIQAaVZI+ihE/HBYhDdm
e0I7BszsUdrxUQdmmCM73qonf0Uyq0JR8PFM1t4dfykfrxll1qYMt1uE+MYqLV//
M5xinXEjIpLztsITTOJOOYaDUmJp8WTVX+4vhbw0gcGTrcb3GV/7RZr2HHgisN/o
GwHlctWo+ePxMXwsMzcpez9apxz8zMAn8SgdGI0frK/++axNQxj4s5lxwt9aV0Vq
XRZGXJu4Gn4pqt5lOJQk6ZR0kFKpBjFzTCQVXywGqSzix5RK1O4wcGv3K6fzCOwl
FC1hKbbhwSTs3StKb6BDr6XWZ9XaRmfcpfTkGgxl5gov96cD2Xlxj7KjWoRQIb56
vkZmZxkuzYuQ8JTwfysKZ1mGvS4dqRGBudcmzkylUL0MI9ULlWxF8I0TDSgHBmyT
cWXFq/Kp59KcR86435GXkgdwvibp+nBsMKTUxugbCDg7Nv8YM11IJmQkAm7xiecF
pg1CP+jCmg9gqvX0KwmdGI0JJI4kcor2ZIBe65Lk0REbU1ASP7fMG5xICbUiyt8N
vEuS/ExTMCGrB86QVqEkDeHeyuIVPOcypx/ijaeXUE6Wy4kaFeSHXDhr4RFl0YvA
Q3GMAvPQjBzly4rS0U8+sptXQSwZjjqkANOSpVWTAIxV3sa5hEO28hEyK/9c2pS2
xrI9cTmRnUZO+xFTeqDcZ/R6s9careDhOIP4uZ6ZfFRenGE5zLK3fvDxbfWUDuED
xb4nEdkOMRwcljb9sCiMBbZMIbVjdc0VMK7X6ku6EKZznRJxHZRfvUVdU6UCBhjx
lqcvfyyzq1oQ2ZpobKKYU0jKcEQjV3N6ZFmSClInZZQ=
`protect END_PROTECTED
