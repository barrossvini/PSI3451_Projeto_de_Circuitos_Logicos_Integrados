`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
49Brr0HjvQwwYXlXvBHKeHab+MgItOeftnOIh9fVyi5HOA+oRpkLDQ8dyQjsqRgf
x8Zo9vw6DTRBKfHUAL0UwDULk7sxIgPU8zipNQ2ERlY4KNwj6NLr4ym+eN5OL2ep
AavHy/iYuJiCPh1XXe7bru8+m0wVemqMaS9ed+kANT8JaVe7mvCbR0ne8ELYzXmL
U4Q9aYHRHz4P7gBeCn7GkRl2JsXyr+vcmPovjE/FRStYCbkrsyZiZ5K4ONTg/CNL
p83ktpdFQ45qEk5uHRN3q4Un80mEyNwXOT9Ucxhwies1Um9oxhx6qNnrUBRXaGFt
N0gi3fltif9KXY51cPZx8R8VRrJcd2KuvavwHSjrUuuiSTu0XuQRRTy3BSYTQKl7
YkFKsQ+XiWnfxRxcQAjCAQ==
`protect END_PROTECTED
