`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3kCv31J+fEXiedu9Op0SsZz5bJAUofXTnIZXdtXoyI4/P8czYPn8xbhcIUOCGZ/c
pXIKkXo3puCKPKS7g8kUnfUl20G70GPQIzBFCIQvdUAW+KBvCGwIH8rBABgavJVV
SL8PqxUV+tAFN5VLQpuGhl11khdsEizmMVwri7ga1zBX9OpsECWEIcDAjgt7RsFU
pW3kV+3j2018WMsFO0reJMEjgVhPh17jFIntfwxRGbnMWIcEpUsRN95S6vyZUoQh
91lT7zYOZkW0ZdsF/rGdxIvtH7gTjFRJa8XsXGohs6mRtTp/eXNKG9YxulJnqFtu
EK3NCQvb6Da6FTrBTaeqZuQAlQspv0HD+eECKHjpaitOnu7FsxonPpvDo/QXwQKA
OVDZLHCSlmQ/nLns47ZIUvGfcIO7Q6SEWPP6+ng1dAQHQs/FyTwN41E9Foxh/YR0
u7qCUQSH0iM/qVqtm9lU5iswA6E/Q5iz54xweB1J7nEBGkBaEOcdIVsA0g4HQ37P
YBHH2y7FfWkTech5cxtEIr7tevgth43tTSl8MXg27Kzh+lKTT3UWAYMXxRsH1OlD
XjmeyOZD683xabONocWeM+vGgvsbca7Rgek2oI15aRxgisgWQ7wpm0FHma2UQW5L
r9zlo58kcWcA13Cfq3Y6GbqgzdCPG4Mc52yj4Gpx5Y9Tlie8bXiuRHiOasAOD7C0
uqKviib5jUn9wJtzfEWE04XKcfBZEFkcW+0sBP9rEzJqnQX5wW+WU4pVzqmrJEw7
UswlWPsm3medfn6pw1CqJJVmhNmBF1CuhcTaDdrJOLhZDRfADM2Ek9kGzA9QXOF2
4gywUoB+7A3UK128s9o+XXUYx4E5zah1zOA6zhy7fb7DCVDcO2V5KxPvs8/6xE8g
qG6rPqzs4IQqhdCoNL4bfA+DpFzC19Hxg6qQo9lGiB9g1kan/9SrHf+SYFs0VvNP
U0iFxwRBI6jX3cqgDGqIequf0Re0ZaUky+PVXFofuAO+EjWeWymczqSQ/38d5Jpe
wsYjLakQeruHy+MusIfXrKdIUoBr23kzAK4KiJIzZfKsHK6gS3hkCoSMkuW1vAVv
hl1tZskwYaqExwzdZ3M8rGaBsYsGCwfnuhV2koko8Ywxa5CddOrX7pT20qWm8INZ
L74t7DIz0bHzmhBGBxshc60x1YHTgbfsv/IwAqQKCDXRel726LVvxHv8Xp2XHJxR
KfVXpHbkZGZDKpqUI1WyMGDphT5asR4NBexBpJ+P6EBwlXAv+2m3Jlv2+a1CwNdh
sVuHIMCXDQijwGiVbVez86DyP3eAjUmGg39OCXpxmO7rfgac/KB4d0bTdqPF6Q+1
+gSZtRaY7oCjmixpupD0Q5BtaHpM3RdIJdenHDOv6e69SC181y0f3ihFmqMSpqlH
6hO7aA2LXp0pj4aoZB483cUPH6Ps/f5iV8iv3NVC8yt+C0rTSk+quXrLmGnrsC5H
o1ANFx74lmjgpN1nE0o42QRKaM6GcJJpYVolZ2SYqzhisOSm5oKu1pNWg5yAt1Q1
Ej1Qo8CMTmsX9+OD0ePYicuS+F1+nkFLP3zVqRg6Qrb5MTsYZPt9P531EgtfdoOW
`protect END_PROTECTED
