`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5OLIC13Zwb+RKl95gUa5qS/0Qnd9NSmZpM4dtcj4lJFHamEfRPSAiGneItzvgZvI
JOTj7P733sbZoo8z3YlO5J2+wZHxLpvOOoXze+ZH3uvtDSxu7GNvfp+c7VOn+9bN
BkApi4WDYvtv9RqttONoReat73+6VOkeRM3FQ2VbvSOpDff51XFFOvBHPYxRCaHN
s6MoctrFtOXMUQn0cgowJhSrcF4CQIQe/8Gz0fxewwmyi6/xEZBNEXPwovOmcV1z
/eHtvCy6xyHMoM4e8At/sA/LE/BXF+YEvFW6GujuRelN99yLqDslNttG0h0rz6aj
+Zi0K2EXsLJiB2p4QvsxUatRu5R2kIWn66H18GjBwwpZWwPkaqbVVFJIpaQlUXN2
BIsQJajkLUC612FxzaBawFuJhci5IK7eJ2Jo12wwutjjds2lxwN3RH0l66lJNpd9
qGCNPxlbjv9uhzc7KfJaK1Q00pKWm74E2APBx1TlxpquKvJqDp2xyRoRRuNufwmN
UnBuU/guWZla1+uvBSaVNjQM9XJqqkUiVujrBA5+LSe2dq4pWpuw9EeydijYuuw/
0CRMPLqMbhjsfM0BzqWnKtFQ0JKy32v4ljVn4x7hKcNudAAxUGCs7OXKpw59Ug3I
xlyu39Jf6zP5aegJnOuFh8IkEMBbsk3f/Kgd+jb8Tlv84pfFeCi5uZI8kujJYPED
lEncmmDrHY1GSYynHvoxWyoxpBeYWKvSDMooYUP7eywkKEkwOqCRz8MScMokcCEP
Uxl+gVFUhCc/3YveqOuvFd0WDBlhdOMZ52dZh5Zc+eNHLgHGxH2c2wOcfG82EUX8
Bs8y9ClCu7A/V/1zyz6+SQHjQCbCwbUGDOPctwINM4y3RYEBaDbJWShkzIiQDU62
N5FwFzk8Fd//3pPdtWb22+Rzlo3nYxNLDM/5RaCS5NtjhNJpW2TBK1km9+eL1+cR
k2PZT9Rv4q9WH3PHvxEpAVksC34RPtbQnT5T/GhrrxKGaLoA1/tzCKSEukW7DEc7
Q3VxwD6/lAI2Zq299HTalmH/lGpYUVeUXPmTCMSr6r9/R4S1bWVKA8H22UxP1Adf
N14aqdbiAZ/OKs4FAvasDKIfUqv9uxAjw3HbA4GxD/y/ISuuv/X+HjehuP8kJoWJ
O/V91Xgfu6nWDv0msbm89rSWfCZb5Pgbs8DLvPBBcHUgfXAOs/s44z4scDP/xS2T
GzO3KEP+1zQcz3qix/FmOY/hLd+81rxHbiz8kqTBaICEhYTs1swakh+qknVggd1k
/b8T2IKWSpHirWFD/hE3YM3RraDD2IYw4CInTaRPBJgeGOajB/LeRDaPct5/Wi/b
a/gTz+/Tn54dqLmwEyAJHRi3oMZIYOR40o5RpLLKdPUNRDS7npCaqAF+2Q+Bd7We
ISaNG2LbyXXPm8Zf+7M/Z2vbFdDloVagxlSRnuem5r9QTha+Y9O0Rnhg8TMAPpwB
gSlBt2y8tVKmKhKHJ0XYOWo92uHMWee+n8LYKuz0+knha/uMcjBcoenI2QORPTk5
fGDatOp+CNF0Ys6AYeqIsQ==
`protect END_PROTECTED
