`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TlJN0GCUzSupdcE1gHGETEERXWRyaSdULtGJ6hN4Obr6F75tqJ4jeiRFpvS8cuTG
EabWuMRIzBysXsxMjmTzsmhqqsC/ae10AN29T/FLrQF3m/0k8xn2igTzHmTd0WOc
ImiYudZFzWAqIyZDpnk5qyALqGbQpFqPKrmAA2mmp7q0m+o/EU1Qe6wbJKdjpRRo
EE9aBQ+wpv5eEMMJ2xpoRnMfGCUNGsvnMNpNwa8dLqXgswlaElQKprLrGPwrvsPI
nXZDSzn+LOIAIRpEnAHmQcBKN2Mkfmv5tJ9TsvLx90agqCSYzotSgwCcNKnZKt3Q
T38iycH3CGfh3/TW7YkrG9OmG4dglrqbSO78rK1W5Ygb/e649DPhlno478ISgPiO
8Iiv/5hzeBGWcaS6PlhmGMGyREbjYIv2lGxaHhYgqrPWWk+IMQjU70R2+dWzJz0d
TuruHi8J3EHm8AjlsdQeK+yiyzEok6RecwRGIWOpOtw3dLWVCROVYjkGgu9EHn8Y
yExkOMJH4t2E/GlHamkFHb0+ATTdQVH1bT3U6+BYs0pzpb/iQG/SDWsenIFy9Kxp
e16Yd9sYplfBmXf/zOsIHGLvtkQiW0PJg1qbn3Kt8lNdhQQbnPrx8L/qoSXOgwX4
u4j3d/8c129IwTBfX5dPlCz/15IhGNOLVltHdV/EMwfK2JvoSHlb6CrrxQ36SFkA
0qzGXPjljw/8JhQGdbXb4B7kr/OMM0q2wgEWIE2BQZmPUD2VyB9tQRxwmaoYtyYq
FlS/m9eIFyY9Z8HlVzY8DrXG148Jgv8NKEXdXBAx0RyvRVzHcJoxKJwlHv93LwJ3
LjGcko0gv0Wb36n2M10Rh5lP4jauPv3Ew5RAcLDpl/XmVw2kbzXIZviyxP10lk2f
5Wc6Qw4k5kimuvZeC86ZZb4pF4SzJUkcT/jDzmgSLO2Ioe2gGPqUzO2VkeOHg7iO
a3dKrj7XWQSM2GUWInF7RrYER5gRSlRxzjRX2zDsn8K0jV9EOio9qCFWXxrVmWOs
Ts+ZfJNg31UKQRWcqbXUHM/RrB34ETnm/vVLP+pEj7RXMHYlbrbWOAHq5N6RHoq2
Eexrw48okroHlccgSZ3nyKtQIM2kLFpH2cLCLn2IVRrDgRol7IhgfOFiBvX2YEtJ
L6TEtpSIvBvrtTqdz2DSQM+XwXU6AFYJjJMr84mqVQFSRH/M7TUy/uLsX8sez6l4
F6RPZVxboBdKAIczxM2EKig5zDzGoLi458dvqLxYZpYv1mod7KCT55Zm+3DGM1dL
edYY3WBR4RtART+YmsPqJtztN1MEEnV2CQhFC+smaBRHAys7yRsus6vDV1Qs1/8B
c1e1EmKorS1HERYrsz0xgtgef/Xz9PMsx5/rKZ9IkJkg7+eBtRkWaGf1femgorsw
CwTm3LlPL5Zb5zAOxTo9HpBXOaMmd06EXWlfNmiDMSOP9RrLEDJja0rBv48zE4xO
MHZ0ZfCuozdYzVsNhwZqvx6bT65t9yPHc+L8d42/o6ID0dswcPtnOC77qgG7Xc76
MPLfriK81md+1sYlN4uKFQucmfj2oDYH1/DM7ma+rICqcFgf5Lujm4hGRs+rhpYf
dciqwvXZVD48TtCkJQfy5SO9OXC3Q9WpfXBE1sjXOsdm8LlYdwq1SuPARNpJPJKh
CljD6aCYnUnsn/orxbg3aOswKVMcS+rfoZVezTkmR2JRz+j//H0BdE+YiT9NsQS0
o74fGmquWswY5Cx29JM+8CctcjThFOV9ufNYqqljtCNw/y4BDCTLgWQMP6pXx/rs
AbnQJQCETD3S2WgaAh+0G1YFB8Nql896BLvRXAkjFj9u9yy6wDI5EX8o9JydgzNJ
ST4gRkGxdI6U1jU2ORAnujQFpm+JdnwPe0xXwXgK+j5Nal14E592zTzQe9Ovdg15
cLYadwGVHwIx3VhYKKm3ANJWCi33GUxA/rXXadhejORG3G2MugZwIPmpEeMgpZj/
r4hdqiQWbSipI4xYbFTjcu2VgC0EhbVp9MY/nTHVY2LJFLVGv/b4O9rqfY/oazTE
OqKd6NBKPkZvwkcV9QfyNvrjsdd8tYZhKH16FDhE60n5kctKKw5FPLUylbfn1C5F
7bxOOVXu8BkrTBZRwmRzhgXJElZo3/2oTSX/hVwkNDM/ZP82NKGR71eC6EaCM8JN
smOOGP19G18eZJDO9jTqiDpSaGTrsLtaMW3sKdJzPXvudj5ZBhEnR861oMNAbWeF
uLJkHJLddCiMic0lE3H6SRcUAjxiPCfKzKkXsO9uftqxwRnvY+0HkFfE6pYQLWTF
+TpJ8D8UJRmuxSxUqvnPGItgQ1/Y7ozgVn5MxCFNFA5IhKIJ7q4u1bP+RrVCGQ58
5WBLzUE+ZdA/l3m7L8pAy0sAx7eMb2cAPm3v0trOMQlD9cnuk8SwtppMhCRVluBr
4z1MsyAvyTHrbXCB0X1mSXduuz3szl3DB8UuRgAySFnWDCw5qxVDG1SVoQxMjF6P
BNhSyhpxNTZrg8URn5lO7jFVZ+QjUwyZGRX6l6VKdikaRFfc88S5nuZQ7aRX53NZ
aVPTHrDEyleGeB9r4VQF/14TyCvCAo6DivfuDWaxLvdMsIXNqRKWtXe0Ycs8TF17
knXHQGwWqJ9b47ZvTGKftgep3NGflqrbauMUFxo7d5H/Htif5JdGzmh8SAYWg8Fu
cloY/KObode6pRwmxdm1ZIVGkDQNgsT885JpjePSUxBSyQ3sZIZ4ORj6pVLiunXk
NdLCOSWKvMqFm6tJXOjrfOnUl/8COw8FHpcCXwa0z+nBs5Q3VHZPnkQjG8M9fyFA
+Ivanghu8Boqlg5PftIgVy+SdMqgkCCLqSXUHjb48ip09MrQ5P+Zm6j9VznUSp6Z
anv26RLKPLDjfOEaaLzCEraaK7GtcNphoCCvcGpRrp76PpjoAW9zvitMKIcf4Fqy
32tjLZEJnAKZ1PItcUwuwXACi6/PzJtc7yC1RSADzQPpnGRISgxia3Rxfk3LcMLO
AMNiD4BENl8I/kbmojyBoWV6+gMtFLv0YlZNc3l8R2QCxHoPOuhvOEoY7K6jx68k
aE93hLr3NX+nQgX1wkFF9lOf41DfKAR8fU+f7ScV9+VCoCZsJ4+Rcd57XYPP96BU
1+yZPggf92Pe/TVghn1yElMJd7VE7xOkEyq/4UE3Bmp3+KvH7tkKwv35BYC2Ugof
eB7cU9DhhXKBTEnR7t4nINlO03C+KQk1wLftpk/yNWcI3N7tBRrccmPJfTns8ZED
jfGhIuOKf86wgi18q/1ViIxOyIFeNr2d6s/sOGuuvL8/GCrI61+UMMu1LOR2OsNn
DFR2y069ZPSGnjwYP5Xw9Z3WqiumaKJdhH1XXVHAoKnk5BjpFlP8adyZwd4F0MBL
D8tRRQdvfC41sLO0FB28FrKQgV9lhg4f3FecKiewV6rSVpDfWGAYRvSMIC7m5vQc
XLVUGMn168JUBvcfKFhhKuw7eidPk0gfONEurE6PekIWazAFgMlCTZw76btb3fM7
PGwAXK4XWuNLQXvbdmh8Xp8+/dQErsM8c74bqY10KNIRRPS8/MJpoRVbk/pAUm9g
qCuXmb7SCXgkJFFi676kNM9m5m9yKz8s437ltS6LWtwoQyNV4NWuqzrUFpmq0Uxg
RCYgQIv0X6536GSj1slZTb0gqcDiqsX0czqIISvbj/yE0WhUktD5IPFfDqbYCRK0
1jXKVu1rFYL7eL7IlKu83mEZy2PxPdtGvMwzBTy0Q8rmb4EAsOC+fw/jYgGdnM8L
PuUG4XQ1dbvbxuQ4zQCX5vhNYX6Ld/w/lLQCCAaBV6HXXYKQsrAcDW3WOhGn0lDW
ImPlDuRmmzEqIgC3nM+L3HCXX4x7TMoM6CiANBcyj4xflSGqkaaLVknJnVM54p4b
ImnLuuAWF6ToMjRN0rIvaLIRqrnJdI2pWKudknJjPlVH8BavzZ2uPj6BaAWAqi1F
tt1U/90/NGnNaODkXUjH2SFkj8QtFFMzm9U3SUSWBQz3jTon1neIdfqr904udmv2
GehkYApggiHy4jLWMmOWKI5TnOtYyUYAZCyzW5kUhL7fB8V4prHTatjdX1ayca5R
wMLhL3VEqFeX/7gru+1PpgqSAqOPNJXV9Q51xtiZY2CbTgddgdFtJvTZ2/CqMlHD
0DzYQxOr7+61gWwWi/dx0Xx/sHULja9TRTpueW0CO0nrPdgybRNoaV0fgCgHYMF4
FSp3/xVe1DA6sEjgDNnpUVLlpYqxo5DNddw0atfdfT4VRqiL1QHOwPQcODcxqyQP
MDxXE30jeBfVX55yScyLfBN1fb9qKRU0vD0ckNn1p616tqarLoKNRENpECD/8oud
cuEiyGgC/4Bf6UBVyn3HIq/Bu8P8NLvFhVZTQlAWYXIR5nGZqAd1O9cpUk+LEjgx
G1rFKKGpfrJuRRfuE6z9yWQo1/k7dxHBYGtwxkvOMozYtFv5ZPKGea3BOkRnZSE0
HKTDIrthO90s3ChYsIL1V1UdClfwR1otMV3wooQUcEQb8IGQz2tgxRlOvICxOkhp
CqCJHQZ3aRMkzB/bEb577673JMtAyYostebiUHB6Vq/mdJU+E4cx1wxfnAZGrMz9
AngSDc0bfZ1m+6MczHXm6oSEG7JB0zuNYQIykVutAWycRHT9EQe1Z97Avoq4p0lU
e5RCPzSkum3IBCFuIymXL06ukRpTqDASHh+x87doTOGsr+5dg5HAUVX6Ypi21XhF
3Dn2izDfFf1cDUiSAbjtbZKe1nki2ZmAeiQrxJPbdlEJMY9rEmJf5CCwW/icUAi3
vomi5zVpVAMT/z6hjmT7gHGW4sYse4lJnP8vTsf6oqolGxZNB+pm1Stf7UoyeDVq
vEw/6PHJp2Zp9uoqVPa7yu3DAZYWqjydxc8Iq2EvlOG0sjxIelouUyrRLgvav1Zz
Jfih5EfeUJ7qmeqb8z5QtoWJTbO7CoJIRI6YI2SDJmcsmdFVLSZyGxXpHWqC59Ln
GSUliPe6GU12KpNOBVdDHWlBdEKItw7diaYgWgz960Ha5lM3JRsCz98boUa2X5fR
7joEYrheA9kXjaG2lG6QIGydblRRv021sG+bZjhDffdjjlLNoRL/j6QKYQ5K311A
0JNgpYxEMQ/XlkqjxL63OVP2tZu7GgU+6z5xX6Efic1i1vuhR8YMDMOeR2tlwPZy
5+H/36m1oUYEIiEkttGdo1rPIuJanL5evcGzCM1MSeOK9vaPM48vH2Z+lVQ1fhca
v+oUBbhoUNNJwMBLAl093J9O7HTLLI1e/ZI5e2T2sQtGNgN5fSAy7amWdHAk/lhD
KyZvfYBMQHIuygpQTcdEUP7uqJ3S7cP1KS/Fuvw7BurMTx0BssBk+BEq1CvwH5sw
wQljcqrSnaH0esbw8ZZNpqCYmI0KHdH2i912a0IR790wnpCiaJxgHR+KL3VY1/hT
rS1UpsZsUZKkK32DapP+IzemyDo933F6/1UnBvNgIcsxfwYgBABe2eplfkvkoWqw
wNaGSiL0jn69il6ubCEIk34vmvnqPenRGCwVFQ/Zmd1zLfL7v8Tyon2LWcCJ0s5L
nB/T28nEawKZ2rdPfj4vTFzYHkfgEnOznzoXSi7nHH7a+I2JhwBdjJsRk7edNyY2
zjD05Iia2hwCK/MiQvtzxYynaFxmbwZrtp+6atHOtopUAcfY+YvHgRR14TO1RcOc
DfzBM3R8tuxUPzd5bMfkMeAFdkvNNMsnaPDY/vTAOsOETBTUi6q4HAGw32ESqzWL
4BU4BstE6bCBPcBQQpDipjHiMKQ+ETV2VgPWWgDN4xQ+lsX9PP5nsdjQLDzm9+29
JBXaq/IMEPMf2dkY9LBgk+c3k/pbsZv/yDBN60mHpeg7dV8swMznAu87PxqBCMKE
8PN3zj+6gdepRVpCTcw7TXDMKbljZgeifxCS8xbTikb/HA1jLyV33TrhhxjdwWE2
UrIT4YuZ5Kn1pzUkt0DO8rKnmx7G3ado5rBKLvx5IS8YiHLNS3UPRst37AGI4swr
pt2/Xhvawx1yIW+zNyrQHNaZFJmy7pYRe5j5vuS3VM2pZ+BjuEOUK3meZuJGhqgK
bBUbpkzW988jaDJSgrPkl6qZnhYlvM7O3H5A97B07FJk6JhWmayWlrhQ2fLlhAbR
cjmATPCePSyxl280vnL9GaZE29bk9EZOtmnoqg5M1ZoVG/mRG3PMHwWsCWzpGFQG
+/D+3ZxqmeukN1GbqLKirq5XIVlBxYFT/Fs5lxhUT+CtKvZ7oZRPrz0fP75uJsWJ
dUIbt235BeTRYfCaZXwS+Eug421KgWZ+Q05Fz+vl/FpAKf0jv44xDrcmVpZyNaut
uc9xAOKRPVyvtzMXisizBLM5f4G4iIlcGZcUW4hIRUroD48+2H7mvkWhwegI+B29
jStO1rqtz2StxqQko6kLEuA/PV4QgZAD8Ci91CzBApLx+kKbZsarpVW822hHLoet
dZ93ytwL7iLDdZkqTczs2/ANj+JyOpbDi3T71sAirR5hx3RPTvecBzRGwooRi614
pllGsdkefYRwB90mEsMF48UZL3ruoT1aGdtFr+L3wM3/cZKLlQZGSHPPQL96qxyV
1bIZ7Myqk9PWVILbOXYSiIiySnZK3JyoOO3QxfYMGXT5cRtkNrCOnww0eyq131Lx
uWvF6jiNQRsQa0eFjfJg+00SvDEeigEndg4skJ575JJREBVrrLHH0sHf7B36L+hm
4j+Xsvs3/aTnEAVPMsWWrTSxe/1GzmMSuYk7PEF0BuN6R1AFl3jWSkJpLb1H+025
hlHgwpBTQ1lF8xhPdsEsf/UkHoi26XgJey6oeBTDytLIYmWSxxeqKjwWAgAbdMGX
eE5rOf/xBK8SufsQtt9N2dU8ifz9kSbvO3Pow/mGYsjQ/jk5OEHRQhUuVwT7RP1x
8J2wpLuzhgz86KYmSzNv/nPbbuUpsfaUNqnMrIYxwUK3DmCwi7U4X14EOSFHrter
W9yotw2knkQhaCpgvN4Knc518xSZf8p88RON9vpmao4UrGHu314CIHCgBvbKA4zF
qEGQX9+/YloOeOgU49qGJTJAHbWgfMPudr1vvoTNEN464n8C9AcJphuKcetr+uA3
8ku+Ot9t2B5HR++39Lekx261bqCjRCghWKlmaO24bagwUwNXVyb26zfWX0+hhaye
Rlf1XSo5gGAOcapaBljITHRQ3gLM8ZCMeBWoDCmmBbWM6lM2CzarD4jPUiQ6rugd
x6FboRJbHxoXZbmIiQRu3BpSc5hXgVzsvtU4+Xh1Xgf1PRlZpTXe8mE9/Yk6g8np
AIzpjkTo0bQRi7fStGdzuJsQTyXPiLtI08euswaTauVvHSqFbTb1oh+qbpEBJar4
uohBk/dOUub/S6zz/Y2y05P+5DXbnbDU1lo4368dMeO9abCm4RfhL+0I3gYMAf45
08H3w8/1ocvwcEcc2ab28WSUS2yXzdR/eu4ibfGaI6Vmo+h+xP7zOCcQOX9e9x7N
Oi1AHCJ7KXbzQ9QweH+xm28IhlztSJgxOK5sGmiShlQgnbm9IyMmmXibajUT/UR2
tsg6ZdHW+XEed854E93l1nvp6P6xugmGILE7Rx3Q0k7Pje/oQX/6YleBSzZyW519
nM5BpDoMvPbyPFW+ZDwSXvplcjviQ8v0xSxPFqSE9fM7Jj18LTMFWDQa+/MNDIWD
bsvFYQxLiEL2//UDBJNFCa1bJH/eiuVNH+5H3AaraBzKw43W2lwXTac7pbpz/oX/
/U3E/tGd+mDBjNXwpyq65JIeZXhHduO3+B45FzpjMlo6O1RCcXUqI3lgydNsUpLR
ZG5wdyu5KFqP9V83kxITrhijHRhXn5ThJBZCBcl7chJ1dLHdkde19Wg+X7eeWAPC
/9FQnFU06p8VL9ojAjIYLU7Q4NBZzluzRFHzmi4tRS93cA6YWPdrNSr2actvuvyV
gD47mend7R92G7AScoxkYZ8Rbq9cxpmSMQ1Qc5+hchyAkQmi0a0Dz8E98O4VeyEG
2wGkr5vx7Rpe1afKeRng/CUzo8lfM/NEERMMVTV2kNziEn26xuh8q6mCIIKLqcEa
Ww0+7MdK77KitNr7uLCYG1+0WtR3REs0xVu+uFMrwa6CVba5cH8IL8rn0Mm+Ubxs
4sKiMSD9eWTdvfdC8m/xVEPre6aKPmlO9hRPs2+ig0p7iy0vViUYyKREplqbypyk
C/E8Tq2iYigNtHTQoTPMuTXdK2x73DCWs8Z8g5rOVAaCQnbkga3KZ2QloTQ9LaNQ
2M3GMdFKICC8eLVQ2qpX2KEaBxJdR+vSS6GmSfTw+HZ2fITlq7pn8RraFyMeg7aa
+S9CC8DOkeAQW/dI7kJnZy47m+70zMTe1la0BQVlQlSPtVpI/06EkfPqW2JGfbD/
Yxn2pk0L+6WwSFs+THwtfdzqusWshIaT/Z+evE4fmUjE7FGTUf7OrAuUmBsjGP6Y
J0hsPCiN+8vUBrzpaS6TxHAEYehhuWzWDig6NmXWvX3TTDY1q1XEz4l8wOcwS7GM
fbRTF3jpsI5BBd2SIZrhO9jAt2tne7/Nfz3H5f91/T38qR1AfS1iZh73g0a50qaC
yg2itjN5PXikwKn4vfP9RoGQ6Nm+1Q9b5O4UzOkWCatfjrgMI/QpOsGH4xn5DakC
LdM9gNYoI7zk2nL2LudAbKW8NqoDjQfFoBYkputvzRf52KIUqgYpqJyZv5rMNDFg
s860gaeGXwv2jZiTJ3sajnuJyOfmw5R+OYVdmLDIeGz/TVS9JKzb2rYE40lwEjES
bsS6dd+N+MsiNbHVvLRbkyzjjaEXzpLcDRu9aZYzmk8R+LHuQkzVbxfga8cYKyJF
07zLYe0yg5qlrG3a5sqF8tRSBsfbOF9RvN/5iHFRtfIbsaRt+WPrZdvnavvviZua
3/x1AJVb32pBJGoiIteNAZ170YoG8ftI+dJ8nt1xfhUkKncmvno2PIaiKkyAzOzC
EeoMmC8uNHDaDAcs9WXpncoPy166JSvM2t2CYKDUJqn/KvTQ7jvUe3iYCCrPSf4e
PuLciyZlZSR4aUP4d9M1PdcSOu8Kv84jvGc8KrYfU2s8ub6Oq5CRyHBVYS1CxdHL
qSoJ9nX1rlXw7bbFpB8JFOWDTYJKR+01zVpmTDA4T1n/cYSPVKQzjNLGWaXA/1ma
nPo+UXScz9t4dWjIRfhhgRbdT6uOM4X0kpGf1NPQKTTVGmJ9uj/ixF6b8/3UbGGY
dUaG6FJSVjswZew5CQGcxMGNmDkfxKaluMcDIGYpAVHVYkBydXwSmtfei9favLEm
XvkjoIbKSogJXa605zZHsTy86aGQopNCqWPH4fD9tEyofCBsdM5/CekDfgv80rbM
JzcA84hOExPdmx9CAyhsPQYPojIFQbgWolsfOrTKKykIdbOcN3zB4EiCJztqmtya
b85fIfXi9+JLQx3kVoLAp+iwO6I5HfB+9SeLl92W6D66OXVo3AZtv/3q3KcpdFza
BLf+ZTCbKUtzZqr2riqSt0Ez7GOowHbbAcqPW/rpK/msTZdYUfdo05WopOpha8Id
i2Bc6L6GsxVqAUWYurjOjeZ7ci3BAIcTsh4PRSBauMfqkmXj20ErOYB1hqi5JOyx
DGyeAP2vKj7BW5DY+KWQVyZA8qg5UHGDiiYL3PRmqgvTuKWErXOQS3sMnuZTyYLS
/HlIDoET8fw5bzZLeoMI4DBA/erjK/dPfnkCLG81PyXjVJ2YunGWh8zyWOwtIhg1
UUS5dnOGw7UWHp9/1ZiQY63+RUQdGSTjTyqb/PZ9GTqa3rC2Q+jTDRqjoeaPF6oF
zBPt55yaRnFyJnwX9fHGBDhaqX/ARAHtjuVI+82RPKprt4Kl3Whcs+SOFsdfX/+f
w3o0kqWelsCElUWDUqasVQmclj7NoD1m0eMHQjB5fJQMcVninCkfShKBz7Esnmn2
Va56y7ukQZLXDWQkYRX72F6h1oCtd9HJNwgbYNlV/Qe7w2FHxsedmuWj/xfxelpR
TDRDlvP7598ZEsiJwofH1VSwALDwqwzZAkDW/hjM/XKFyXoyUn3QZgss0GcRBbbn
lX0o3//DADqSgbV/bb2UGBL0sk7pcIJQoc+NPBC6Ixj93XkYlliKXu8Zg4hfM86M
8ZXV5vTU5tlpK9KA4zzJZKYbfU3pUOlUP8Ymgq6LuOLnZAqXsXgJvw9ewMqjhp/0
yVJqvseNfsnGqPMueSlBrtq8q4WCXypOf4T4BmC0bs/18XGmawquCQLvwZW6pbFL
vnV2G6BC9dIBLy2L1SI3KfbPeLq6tMBB1hTL8/BF0BXnbz6IwBgN8L/lCQxJxq1o
1iXf6h8cCVomEeXErz5Et2tvXImp9YZxaJCsQD+g1sS0MWm+rXiNXH8Io9lH7Rb3
NejPQG/tIYD/w6DH7mYyU+lgoQEfiDQykJjA/lE3TasUPa40yoAYwYVzVmDRWo+H
wesCY9jfJY/YGk8qEE8p+MALmayF6dOfUDMI7at8rOWArGZkT9wqPRWm2QjqiNFW
mz4UoI0X08qpZKCskmj9TVLztYAAh3kMXPyu+vBvcXq6BQM1N0jXaU1hbDypJnNO
MJrbZiNEt6QNGIJUtEZDNzbp/gn+gQC6xXgC2EP/YioAH5Va5DIn98Umuzs2koAE
PUEuavZW+Di27rdaDJSo/nBdzyeHG3h0pf0cwSBbDmXkZdp5F82tqHkCk6PwP1HL
uzIl+eiOsfunUllfotzCKmnlqAMuLFntwJf6DSndROEUVsVAhzdlevlHF6jkr5oC
XdxfqKchknOWonlY+6iqsiXrhAQp0V7ZDLiU4GSOtRdNjH+0iPe9X6DNaS0XXSnV
D6veurFcQD/rBVSPRlOjMooNE3mVZFm2CaW/FiqQH8Sloek5r9SjAq/5qKnIJ6It
Q15WkckfdhQvv0SSwTP/gNBafyazFtnkLGI+VfovGuFpTEyX3MSOeagEHwjAxLSR
G110t6fBpxBaFr/dAjPCQjrjlp09pTbrBlcRpEjOaRn8WhiNkRfWIR4ruZaNBo0o
vom9tchxFp8D74iTndr4Cut5m+9lK1H42WqhYO+adhbMvtjyN1qVTS9ylWi834km
dI8MFO3CsfQo4sP4SgRFhJt5Iw7vEeqtfsDUJYD6kMfJzBhZbtrILMSe2HHan59y
cjjsNbUC2ku97bx4mpcJnTqXTFr+DTLVqXHcN5Bk/qON2zivbPyJk6G+8cF671GA
m8flVefkXdgq+GSWIoye0qjq26Aqw4GjjVF909sbGXARSzgorrIk9orrK3qOADTn
GjrqKqOMWjfT73PBDV0zOIkYr8UkIHOjrXhn2cc+iPJihR3x96enzcwXW802TpHW
M+NWnZQ8cZMG7YQcWXWzURf+U9rLQ/Sz8lx2ERxCt2JlAxVB76QxiK950+xvwRq+
4vb/38BS015h6SxX7Oov/mZnViYvFKXBrsyuKeIGpCdZqlRfVUrEi/e5C9rXpJgG
dJUZK4PQyrXiLCikuolO2ShnNWgYRvvRH5MWs+ZNjNpD+uHhR0rmgwsdVsGOVcK3
Xgrzi8crqFnCWCsY2Mz+hxq+8duN+hQQFbmlmhVRww2jpYAmJ5PVQBFUL0PmjQ0H
T4QhPjBWmgoVRsg5lHkrpKEyb0VjxuAB459n4DplvOjcxj7nenM+kbHN8fSciKW7
//W/t5SfKXoMPML2lOeVKIfzL+ypAyK2kur/aAQyw2CzwgcCA/H2ihdD4jlYojYB
WkIUJ2F1U5cHBRz++8RRvzp5WSevy6xgL7UltvVeZgp5X5PilkftJXy9To0Yjfqe
HvjAeudMTX7MF3AEBuNO+pN8iMPnMFlIoWR+86TsllhrvrwMzA6kdSeiGtNEnpZA
xHvKfhhE+agYZKxo0bue0yRM4A5Q+z7DghakR8eOIepqszrGWniBVOABnZpA4xgn
F2bXrVHKcxUylPIa1lMRIShFyhwU683on6bz3NHTWTpMF5GnGkiwKlel3axq+Bzh
Di5R0rHWcaQwvums7vcoif0683UbdUm8iVtHjMD6BhPt1BKWLTEAtQ/3IT8UMyhN
cX9DNdGHhNN9eb998e55RUl9aIzosd4H/YmVxn4cm+V0xl4Si51VTVKGF9WMXNAm
HAJFppDiJB6h9JxmvsVEoO0RNoSPX1QQFgcWlYFbU94ieLB1j3PpbDsaKIhC2sjJ
zR4OGJ+fLf6HElctVoPofHaPqceHa++EpoJe6oh6W4DHtl+bwfrYD4SaX7PGrr3o
6cfbmuFllHu9aR6aYUvgrw4SpRfc/wCZi+seWH0gUpxuR4kIcAEU9M5AV35IAMlB
DdSO5A9CPe5NWvWPsKA+Fe9M8nr53Fnz3vV7QN23jJ5+44oLNZplLRXq3ZLDFz1V
iN/UCbWbogPYwtq7J2wGpB61BQx3DUlBv421sq149IrhPhBfwhs4xvHQg57N1MQV
294Mr3BNfE0ZCn9HSpmu/i5VwW9MRTUya1Y2DZZV71T1Ahyc4XFkLimcJ0Vq1yJA
Mo3ewiSERAhCbk2uL8IURVp+8BdPE25+heUG+2voC7j6gSfa4874y75+p2Hphpkl
EmhJcv0ZNDwXeF5YyDh+rDokBKO4tJqVn8i5rBDZxfMVelfc2628Z7FHN9mrhabX
vw67in65UtLFFfVzX+Uv+fY0CGzy+94AuQdBIPPwrtgDpN79v33Co0XOyvQvBQ8s
UYoXQktxnVE4wUGMGzCPWtkeX67VudM2ePnp4Ir4qwvEWCd3NzrB62xN1UQJn6hV
EjjlvGmIUw5tCGJpqmdbqXNgVaAg/E8kHrTnJGNZX+gyyf2P0gwkHU0G1rz838Ok
IAIzFOMrD/RnPTc1eo2CpL+9UHolK5+CvMGRtlrylDCFH2A/jww6gawGGQBestQ/
qajjtUC+vMM1+nBITAuYntq4p9uOkRgLOmv6FYDvoEIxpr+g6Ax9Ze4kRRWVr3zL
SREjjSLycVerRRqo03fZxfotSPU8gA1cYorRwVhqi43CzfCzd/ug4O9CqW9Pys71
LDRQSKOmE1t8ecJfum1nFE490p3gEciM1F0/Qt1hRurdeqJ5gAae1SQ0tV8d9jun
ra3xdjXsSG6Q1dDaLlI27bHFxOjwVDhLS+qiHVfzKKc7WiGi/g4Lgl+vomveGYRa
beKk89xi3iXKN+Yluvrmt9CtduWWCP6Kj9mnxPcNkVmCFK83rTtkzhyiCpRQsJfy
+4GrC9iGf3dJVro+TGdntfb/g6ClQn35obfxEepGlL39uzqx6IOLezIG09lqiM9t
abhasCynpC7uI1ZEQHFgWhHTXupgLDBLMj/VGJWmu5gztCsrOD2K9z0xOxl8ocCk
0pmwRdT88xBufbcSNZu2r5j4VNW1PfnxmCn9ZC10zEYtwV04CL+oLG2yB3SXFZdR
c7GIcGk729Bo7xqnHGJGA1altNxbNNQxUMdyfjqtq7Fgs1vLXvN+m4GSAF1xIPlD
OxZPEzlXsE96zEKRRC0dthFDHj4TeAKPfjM+qWa5C9zZ8YzstYvPzMszqfHIRpu0
CJiYMTwhMvHrY6dpPgsSkTKLunURzUhcMhG4ueaZftpA9uokra8yNu4A6PMFOT4w
gIZSgxA+u/x9PiEE0DEaBZYs7WlI5/9YrjxlG81FatqNFbVKIGEzxA5xdh5jK4hi
di0naW93d/z2kztCR80yoFuca01Mh0tcyidtdsFQ4xA4cclcPh37mcbYJo2+0mr7
tUs4l/inIC4pvhEWjV0XI5kGGLeG3tnHjyIsgd0GgfIBMtYNNW2eB/uqwO5Ss0Cn
UdroCq7oYf965z3YFYF8eZ1Y/NVIzRL8hqCXvdDPHFCM3W10tD2jRxoodtpgAdwl
p0TS+i1bTvi8vk6rHXTmzV0oXqSIaj80INE/hJk55N5YzxK/PYTobiWLQEIlhCpU
dAu3Bu9M7ZJDDk2yIClMWe9OB2Z2e0W22HmwK9EZxNdVO24r3hbAU7ElV+6XC/Fl
Hz2dCvgXtiidvu1DTHB+SnYgCLjhkKNQOY6wvVSnveqRK9P3mM1MKmtB/K7SMmDn
AkZYBgFyU8pSYOUZ1lMynP1xcGtCrWEchQIxDEZ1XwXLOabLntNw8XXy+6HtDy8O
ZV3SToZacsmalv3Z1igMN/x0AYSokFtT3wFkFEzzI+sg8Qp33ho1QfykD460AkJX
HZGm8hu7G11Ds9hqZu93qybjYaAtAlgqxzkj//ZFaO1Cd5SXHYz2/Yt/CqElsbDG
Bq/SJ5ZbGDKqogCqwRfATR4SnT+DXGGYDdIhIPVHLQ3K8ZoKfuY0PzVEs38D7Fj3
pbjmGch6b7LAKg0aRpkolTq9jF+NBOFes+r0EFsm/TMGIbaUx3eF6RqBfvGylbIL
BGl4w9MGSCQHjtLG9px3cYVYn6s7PZFmyVmht5UdcWmB7MhBsJs17Fo8okw6FrDz
HekWznMZ+3YVadyECKbno6pvEQ+NO5xWXTBTVhGSu4tFB3Upqn9cstFfRwHU4zwE
liYxDMZw1N0E4fQlYP9JMdBWGpJ9Ed0MZEhiPP8nq7RjOB5sAWgbANGAHSGM20qh
DGDoBDL355Kf7joazIfMCXwCMbmHJ+k/zQAlZ4JrfNGrXExjfzq6Ddfc3yvTK8N5
o57IoXNgSRXlN/BIxzJHTdF7WbZIB05s8BdpnYrptgxiYkuYmbHveEF899WX2aJZ
HHjDQBRLW15R0kQp9Az49JTDvegw3Ux02IRBi4wjv60cOFHvwzSf4ipTswqSsQHW
5zOW+VAa6vsNs/dPi3ywQ++1iq/SRg66KzkMfpcS+9mV7TJfVt1pyIoP7C5hhc9P
ZsAMuKBhI4T664wd7oinmwEW9Ex5WtVCswGd6wHbe0yDl+WAQevN6iAvH3d52D1G
DtMnEdRHeFa19PoUdwQKmCNnfXvd2BKWsTpKqTdl/bSHRy3FukC+2svgzuFdFEG+
WiuGtAEPaBMBnShVtipg4hQ+4iJn1afveHJm80/9sPFpbhQ/LPyP+twAK+c3lLRK
VxW0CITOp08teTtLPF+KkmKjcKK+jVirqTN0P5FLO+DCDcBTV18mUYnlYdoh3t1y
lQnS3mcvHkccbW8II1wRqJYk7LMecxJABcV4XAP6RlLqkG42i27GMGX5IEvLAOJ2
GcnEfjm9lJqBMrX2FhyAmcjzvTjs8xPF8iJeB0yIMkN3JNRBkWtaA5MxAN44jXkw
WdWBsV26lEkP3NFmkFPAEXAhITpXyxf+kNagOkvFS4JQoPpyZ350/8sLPZuevNJZ
HNks9/AeSeuLTevOX+FBYrWptYl4sGbgED7/4y77qZBNiU/s0ObfkU2AZBtZe28Z
nCru0f5I6ESOHU4J48JLl11D7lXgobs6Nihj/QoIOczqzcVXsWr7PfLVeWdu30xQ
Jf1MBHnMyhIONlUoP+PWH9VZsglDw8vfakYx8fgBTmxc99H+48CryT61+G8jrAbk
cXmQ4E4Iah6CwnVe74GiBFms1GiD46RrSEIfpf4ZeGcovX038KoVpRWWSBxPX2ux
tGCpfgKChwtVDcvwyrhAcOAw7Y1PXm6fP3/wRdU/X1MZ0BzldvvtdGFlvQDZLLsk
64JY7vwa49W3of4gM78IHvYrgrvk+P6bf+hpfGY9cfKXuwSYttmoPbcaFVR0GTC0
RjAVeTH4ChdlgYqUfvY6U/FApG+jwBlIyQMhV4igX/M3+Kz6wSR4aCwutKTGR7jW
RlGuQJJKNu+/m1Y96Xz+M02A6jOyKya0fPrmV9NEb4++jr0lfo4a3MciMoEc55kA
ZqniK//9G2COaHGGQSFHmzmPonQozcXRc6TPVuag6JyBSFDQzNNUmBTmXrXEKiLg
GzW0DIqUQm24kUhagAnYPnKr7fEBjctQKbj2dqyX4FEMJXixiRFYD2JifF3Nsd3l
EHJ8d1j1DTwjq+QRb8oEf8vc4TQBwCAu0h9UwErXcsM+j4rUs40hXUl/oa2mm/6M
Wybsoil64s4EqzpcM5yGcBFZxWnul+NcujPi7Wb4RlIS2z3m4uVDi5ULyAufZrZM
frWL+9dsGv6dHwpKs+5/z12sDUt/IFcC4DVdQRGzoC6amrqZPTbKlb8lz9mHbDod
53dWeOdjtFfdKrs6xQwHfwn9nWrO/xva6Lvk6nWspYH9BVIFTvuM01qGbsBRr2iG
1UqPqG/UFmP2C1HrEcmoLI6HJmcPxji//AEpfJN9hSKAaypMW57WNMWxLpSa6++i
jlbETTHPE4ozYgQpF1eiOcSl2hMwpkQ2Fnf/9tbercH15L3BLKy6CSWj/BEb6IZz
qjE4EDs32zcDytveKsPkYhfvgamBI/rlaCxs8YqTgpcZnzw3yQjs/cRwywOtnOkg
Z17iCv4Npjd3Cu2+YP8SmMnCnov/VvhArN5md2LdXZPYwHETPdvmqWo6NzF4FHnL
hlg6AkNIJU6si7Af3ZPB5AnmyDRL1YzeCVqHwNZSqwLS35PcT+XwcCH11kpYTptd
6SCGisSThn1mJ+PIYAjK/th17Pxcdpt6VFkuusA1zruNsq+p5c/LOACkznR7OmS4
8AwNB9BU57a08x+GpLsb+NWeklo5QXv0U3DDMHmwDw7xa0HYFv4LEDnWFhNQ6s4c
QsqFCa7K9VSomHGobKvMqmIGiHClVjpiSgdoe77YLVqC2S5yuh/0QK5BdlGcdqWh
u3xPGLhhwo8pFvoaHRdE4YwHnEJ63yFiKExPUeqnfxpuI2ZKU4Bay//e4b8kadPU
Gm8J2ClZDw8l8YgjiaB8Dzsc+c7yXFgl8bhGCd9uULjBOMHxRXNPlAv8E2oiyT3C
vIyezBtMr8Be0oDYdJBD6vC3PRbmwuHc2qz5hEPl0hO+y2U1gzoivUmGbmGDR4Hz
64fKnroVi4+Uqogiwq9Cjifq0KUV2c9k9GvIrDYit+AO+Lcquyjg769uNfaxSaYy
e8GILihzskk1u2e0H408neM/Z2iWMOPkXkxjbzMZf9cBy8UXUyLLaOY7G5cLm5lA
6HQu0wkfOJAcORydYbQvUTqtnU/SLKpYSvzSBj6c1YQHz+/n34Tyr1+UmtwIMhjf
oyz6/5ELrp0X2/aokZyDLSIHeu7T42xoZGxHBdc/TmbdDxo4/dHh1bCmRqZsU/Rx
QTvi/IOstBEFctrREEOOGQCvszVeM9hxMgoETvtVNgwM3/4Lo+KUMWiTWCwqqKxO
p87BjBlGNMjDIbj//7uID+nB/uXYcxlNnEIILJIfgTQxUj4Cs0f5N5c9JHbEpJhu
1SaFe4Sdo/mRiVf1lIa0UunBnE4K3BhRBEElhrRs1ESi0shLoCRwQ4g0W5uaaeZI
7QmTYaiPUm1OvTIrrIAoXjIbMnz1z2gi2GcLEhGjiqLviWX/3NQEmRyvp7iUaVho
atCCb6OJLpg5Tkwv3gLVR5K/EdLk7ZNrFhpwQbRf8UZSZu4xlZAeTPAar4pv/NH5
HKbCNf/eK+HRHDYSAEDEBzoFmp5a2EQ150vMPW6efZrJfzRzPQGm13SjtRZQa0bc
Qal3L1HVSZdLg/gh1opT7QtBl80d9wyRrm+bp9TIt2bi3w2LTA9M5AbJ/bSdyISv
X/9AzvJOC0f+x8Y8F5VR0frSJjZqaZlC8Q0vyuI3ZOuffyze+o7TeC/vvMOOYfWC
npCVHb6xur+rouOS96giT8uTprurZrxbqWc0vWU/XHLL5AaHOLMPn3w25Dwc7+ja
iGVEcDQweZ6fQpSZNovd3BkIAgYqS97A3AwmU85gcSn19h96uLRWtTlE3ADMLpdd
lltaz7HgTb8Q+05rGCuRVTT0UjSaZZtD9JUMqKkVNs7VtEeBejVuKvY/TMhKItLN
l2U0nxns2Y6akjAuOHMHP0gl1I6463BZUksh3rGOBtdXvgBlcnLS5LgYWt4PRsDS
LdgdqXk8cZKDzaMyGBYJmOQDh7lKNsWqI8zW9qeogF61BEz//th6bABoPLE0bxt0
jbBIrdaOybplvVFd8hSg8hmHjtMgiVNacWKtH2PJR6vEruZ0Nq1wu1IClBAZiFwf
AYhPi3ZdB6wFAOKifKmdLr27emA3uLN9BhU+DpNULTg7aw5ehT1uGj2h1cgvf+Fm
QcmVm/JQPdV7gC3z7TmCbRZ0KbCSEQOR1x6LxCyofOfWY+2eJmNjEvpoNMXsyd18
Z7xVvC3ioHx3aStCUUtq6hR3xNL5wP9vnbcQIGioFsbRDU3XynTSDEI2/KHnex78
ht0+wrqQ442GlKFzA33OfJpx6hTVqlkOL9pD1IqoPc9CioWn69xrC4VTk8Ghd1D5
GbYlLoinvgXf69aSBKCeJOTk/CYnvk666qnOhquLy71R05zGCz8VU6L+tLI9iQxr
cylc1QTYFWsEIQSKD2z5EAojbZt9XODxphmnKCM981yuuR9izN+FIZ/TMxn0cxcc
SNQ3J4OLwtNz2JOXRr+ToO19pvq8hYoZq0kZ/TP+et50T6WirSX7pjN/LczfMkkq
DnZM30owE5EpWTNHUraH6lk+pXtWnb1Cj+n5IczvsZKXEM5hrQVIOgPFaAmbX8lI
VH6aVyOdl+J7TcvxwUavUlXmi9Qp7DgdvNEPlworK1HXdrN29kIuwu43D81Zt239
+nMCEpbhsWHwactdFzpwcAxp38GZo2M7nqv8rImV6JyEjKFPmyTPo2VI9ttYVQIt
ywzfpcK2WS65TF9FR/DLaR73uwYnmrthz0QExw9IfGgTyd5OZRfR8jCdLtDl3q0h
INCg8aQ7aIK9QstJ800lw1CyZggeidqDr3xUXvgDmvgcU6J7ich2Lk/As6Bl/75l
uJso2Hlu6zmMJqYLgkt5X3BkUa6pgW4t87xEU0YjruggcKXqj/hdY/BmAj+AZTrH
rGNhdJEWUV6INIrbU7CjcxedxcHUeIyuS4Arh2wWfKyPpRDUAEjqMCz9YL+neqSA
VvujRBcB3k8xQ2BlYdNsP9oOepTq0jtIh/DJo5QLM07OGMYs0RUGOhql2zi0boYS
mEArc6jx/uFOPXi46sHj4sCUT/SNhZs8CQpIm37leQQ1z+EWNeSGB6cjWXRAQpxb
BTcjQ0kIld10Zpy12ZzBP4/G/NTbybpjZii29nueLgze3capH2cdaBkkaoAYXlLF
c+vrpJniei9291Hy+DDmxw0Puj9B9iGK7FCIVsNWkMu/+JcNO1VZbcG5Entwn/Ws
N+Fjgh+BtN+MZLozfv4GlaG16wg3nKuDiEh5jUX+BpeQ1F0wULpI2ZMUdpEczt0P
Tc3biC59wzeC83KYglcB2HOzyIUFh1nb6C9NyPFsg/SPSJhicBOhxFEoRAjyNkm3
ITK5TV6xP+9116ZjFq5YOwzzLbLqQ0ij895sbBeK05oMbCXVoHYDMGWwctTIHuUT
Nk4pdsN39rGk60cl8vijRyXF8GkTIdkJcErLRUmDddXyJBJYlBUU2DC6nNlzLaN2
pQFjYdDFu7msp9r5x1ptDEnUZkO4ZS1usctp9MNZq6H6+QCchQuvIzkBS+AjoKpg
OnrFv+RLcBT2W+EnrBERzpnnQJejLgMfP/LbhaMM2lfUqv+7X93nz6eWKIeEZH87
C8rPgz5ZrcoFoQ3se6sg4AVeMsb4x1uDMZj0Fjokr2eix3chbAKPwa+zwG4SLcMq
ippDUzUocNRVQ6fPtQRRI9TYtNobQQZT5TAxPmNEpIDMR8md5JO3FT/N+nFTwqwd
yPYcl2eqjE9WT0U6XDtigT61bl/9qPaoxVtcA6ew3VQx/lb29K+0/0TP3p4zmQLP
k79SY+WMJwfmxZdpsM0akkjE7QjOzMAxH36pZUPXxW7QLknCNQoU0bdkuekTYaID
JvNZEyG1+bh8Xm7tn624+Mp/QBlu38ONXnF/qYt48p/EuVnHYpG7Is69tH+l73tA
CTtVE/+5vCUtGnKWTXzk3tp6ys4Qp7q+Vryejqa3PqK+SEjGPBWCDNVQ1HrFN1vT
Od8bIVO5v4jgc+akjykm7rkC9rh+sbGPGXfBB9+F+N+CezTOX5EGsy7Qb/e5nXRn
ChsbGC+9MVO4KqdCpKaNtOpkP3BvebyA95prYa/wDOPEPPeJDSnT2j4Dg6t4T7i8
qyVO4Dd30cDXMWx7kImiQJjA/xrqouXAHr7Vum/s0melDLjhJubTh5hgk3MpNn0c
AfPaCjQq3ab7R/OZXtHk0Asm8xBkLc57LqsiCHzcjXmb+j+nUzfJ1ls097U3zPjb
gQz3TPDvdh/AgpZfLvTqyxtXFYAhCsjwnlBG5d8K7zUdzt2At0puMpKO4VzAlBXp
sSIehNtHETWD/UM7p7RKiXYLqBatgO6yMbRgcw81vBhswNMtT9+L8JaAmYmgr23C
L/OzUguNWey2TAkYE1UtUBR9kvRvWFvi+FJ+9IDmPLp3jJMV8kJEqjxzwSjBZjYl
FBkLi7C+yoLtALabXioz4dFNds+VOm9wQwyl0s1tHQBeMaBqFfsnnRZka4YOkMMO
E1e90G79yfBg34byc16FPsSZmTQzTNIafxNyoo1rNhZdL8nTlvxe/Rr3FURctUdc
WZyvWW4st3p6rGbjrShdOB3MqgpWti07bg3+jkm4QEb/acZJuo5KQkXu4mAXmD02
p0IBOS9BZwSm2KrOeeGHQ7jGxCOew404DbsvGVUVm8KS4iei5/pOKNXW8IxZDzAd
sixT5a4MZAVRtYBcHGQgvOXVWwUPsiedlRylJGz76UPrBCiJF7al5BWIcH1/J5Wx
mPJxXhCcU2vGKhi1qaTCs+vpzMdbyNU5WRRWdurr2B0yHbYDLkorsaEc9SfhTBdv
sikn9eLNeSVklWI3UhxFi3qtkA5mjB0nc2PzKeWFvFBQiAj9Iem2edQjJQ8nZjR3
15vgHxdXPqJ7ngbVugZf81kb1IQ/Xxgskh57oIg3OhiV7M0Be1752YBe1kkAZy9f
6lCqAE89w87ANOKktBIToosVlgZX9U+Cm9goC7dPQSmccKtQGuF2iWlheCCN2C43
USwTTWA0fwZsHRBXRxkbyUJuBIOitVEbhRhPdecWRkacHh3RvPvrRhu8HrRwLapD
UeYMH9TTJYJI7mT9vQbhp4SKT8sWmISmsIkuH+LPf7zCauckj/pwhy/J+i8xE3CB
BtOT+RkC1WXPjFFb/Gwwan3kKAf47PTx98fF39UKUCyvS6tRUP0o/f2Ku6ihCPmj
B/EygrJ+4LCqLCfDq8XSB8z0bF6VZNLNzNbovzzKPvvj5FWRu3Q14COJHisY6abK
xKytH3SLq86/pc0OyKXOOq25QPunGhlmrn42X1TtoF3uDBa2w6mJ5v4jAaVEJ2UI
iVchnMPNfTfKqtLwaNSd/8OABxxekSErZHSHpgyuGUQjooRuy5JuVl6ln+1g5cDf
cmuoYBWcvc2uEe4NsFfMaAkVhlUCL7MfMr1rLAi7MQGg7DGzUltPaQVlQu/F+PJH
YKy5MbHHgPcs1b8nvZG0FFd6y4w1IwZpWjQokmLpWVeEWDUGMogZVbt/ELhkt2RQ
BfUxzegP3RXALRQwuk4lg2Ls2JK5WEembA5v8rzA4V6WVuRM5lBCCoEpAhlX7wGP
1P1CTTATfhfTvKkUYimOzyKcPGLe/dv2Vgx4Vxgq4hRSqpE5ZC9cVc3pp8VvNuJl
tnd5SPSlQFfNnib6vm18YtoVGLdWe891OE2vWlHXErLX1jGL1sbDEGdwXP5rEXC+
Xg5gnSNxQoMTgqmVQnJeDHD/cGYKnZbh+xDHw+3MEM5E7JivfeP45k1MdGk/2Tqt
G7D3B+NGLKebANEFi328CyyovCcUKejJzzklnM2WxGo0o0nUAmU4TJzhkCDx4Abz
gNXuzGR621+hNC6/t3PdONksHxYMczg+OD2XzMr3r9XA3vW6fN0+cKo5UQkHxVT4
f/ko7Gv+/8xk608GljMn2Y+A+6vFnT2mTqzGZfQuIWACn0UGJMfwAD14+002e4nL
Vo0aBDlYSGY5vQYOvDePCHhR/BDGKuK5SXpXQo7WVWrBf/eRzirWECjKp0l1+USe
DRpjpG32gpAxh43jY0xlwSZLbj3rs8d6L3+mHLQWlSGDdMO7wQ+BSuTWK59bGiV8
ZyFoDAyYjvEvZ3p5KbNg3VK2OmsnwGhHbey+a/WGFEa6oMaS4tnWq8O9QoKmKbTw
0NZ6j3wWhyEh9vStoc7kqy6i8D1oJ51gXVhyfyj+QFg8WPCGowLAoOGB19vpCn0l
jnuGMfP4IFno37GBogXH0T5sUSvWXIIM3PQM4GrlNV+0AhMQpg1a6CtB7gNaLcyI
yL/wtmH6VVgMikdNEeTWxXt8jwo6A0400SKAWhhL3FctlKeIhSHKfKaOeW7hRtwO
BOGU9Q38x68ij1igQvZWbnS2w6msco5Q7zKeKhzzePWYmvHCUFzpCyrNjajMe/WV
ubkYy7scrfK9yi0ONjMuoVkIu4dlw/Krxlgf8Shzx3HiJekGj7IKJp51XngmA5Cj
qitMlmTNtYQKemS5pKTsquP2ADuPKRS2d0ZEw7xC6rAP+m1qXgnORuDYwU4h+UzL
qvqMQugiJg5BH0kJG2Sme30Y7rVXdcjmJ4rdZzI8Hw3thpSmUX+3ZLPVR1Ni9jcx
VnTwDfysMMdpns2qyVhvILc+VUE1Nujp5ZAU8iSe0J0SVg8NnTVlji1M1KsdyAYq
8lmQUtHWvF0IB0cnGTksP98Htc4P8N+Snf1u7lc5WOkvFn6P0AhrY7nhghoAhKr7
IVShjMwLPPIRRBLh/K2nRJhTiJ59jIKIWhNPbcGwTa5rVFtzwkWsSWckvO+AZP1k
1ML9so0aQThY0aF9NqUzKUMDvcn/2W+8NYr8eNo9xHRE9pbv43srmJ28bve+3dZe
AF6G7J3s+iLiKBkjAsY7Mzen1Q/n/cZ2UdqgDp/Xs53NnFUgW1x1Wa553vyoKdgA
vA8hHaV6asAbiv3dxGxDccD2DDDQz0KH2f/V2g/nZ4WmIm1qNIf7oA/nBECIfD8Z
DDH3GnHMusfFFzP5iY+w8dD9v+PmZN+gj8q/KzPdWYrf73tHs6GY6KOpf3ZhaHtU
dg30xddLYjKxwgtv5W/DwKn5Ue6NSNNKqiGpO9kNSEqJFqilaxX9u8x9DiewEApa
d/8JTnsQFQL9AJl4CzfXxy02A8KZO48eJQtluDL7f4xZd5CMmtzFipbtmc83M4MP
ZdYThpoZgH1ljyQgTbrNmdq+FG61Mr8zDKDF4S0KbmBKyQfAD4lAR6ujfpAVPYYC
4GxNfSAP8VRqzLuTJnqsWOwhnjnYJGH4bwWqaIdXm59IUUwYD9psNL662W+UDzOA
dI8lIBiiYmEix3TFoapeApz3e1GJ5d7dmqicKLa0hOiCRKAmT3uZzuRpYQ5dbzBT
qHhLoGsgSNIPPSTIS/4MFE10MdXBF9vbJ/mNXeENw8G6NVOMZlOimJWtLToc+vOq
XDkzaxfzyXWezrL1+H9zHx8reQItW0wJYjiR4b6V5Ap7lP97d9l8mjR07oYwaOsE
CuTgEEnxPuK9oOfp6twhLFdTrUg84vLqgyUpzsiy5iHhH6v4BTVDFgS56RQeCQXG
TqYUAGDFBSH2QP8WYcsgW4mtaD0thHCaHGtzN2rsS2y2dq2HcpoOIou5RI+wPhQZ
vztzOoPJwXiiwmgnV2wXgQCooUbjiDmbmxqlT8WAAs9kWWuM7uUoHxtQ9zV8FyF/
5x1pTtahk3MIhCRd32qqxk9NkhPQL93KiShAcjhdNLPcF5PI1Yi7K1oxRMEyQkUE
k6E2fl50f/dbSEZzPQd3iMNU5HLSzWvtSPek8wjEwQXncVsN3LZecFpveahr56Tq
3D0+7dzmbZAPM2smEk3KFkf9lcCN7mpUCE6jsxam2j2jlQKY8jtjJ5WoU6qayOHz
cjVEZkbPGOMInjMshwVVIy03mATutsw4vv2fsWlj1JXMPPTbNCEVGx6IvN54KxZ/
wn8gEiRO6ZFSROosKVUDH3Q7rEAfBssHyDJKUkI7jf6IOU2pKPu5wgPIMoQQ3fVo
2F1tkh3VBAHv01JrlQa3oIn/QpDIzWmp9rFhKTAxcLMhmVuuIQYj5cIUwvSv5pAs
qaNDBQNy393+GSJoa3f/J3O/SfQCfgmys7VS4RxfQ1yDmbBBK88v7sfrxKgKHOMH
2cq/sFKSEaMTXBLyJJ94KVDzgaU4Z8dlGfGCksd+lewnprPKb1hoeMZIIimbvjy4
PSSEjzP63u0odTEVDjOQkUCbZ7Ktl/Te9baWh0+x3oIkVCaXuA4BbnXnwR3IhXZi
LmxyolzJJy5Bm3x0PTFVUG1thA+yyKdLw6LTVofVDOGday/3TVpN1MzYRHQutL8w
bIdgxaw1uxrhUQtw+WZfwQ1YB9O5AHqIkHnlve5zIh+kGqtTImnORF/luft56Anu
bbScP2BHu6LG4jubYYyEuFZ4aYjfmYPIi7KQqyvbTndK53r+3esRr/YLcxVIRq+I
Z40P9X/8ww6nuwrUtvh2xm6eyJWGt4fnkmYmyWag1Wa641Zourx4sC+g+F5buHNM
uqY3/xYf2eoBvrvy/g14kgWVzdMQPNn/i0HjR1nyPkbiMMp6GcFh3Yvnwl/3cyrX
BqxQ+sWz0Rj1O+xI7/K7+Zglc6GeMSS1LmYJxGwq42ayAjT0d1etpBEplwN5FCPX
ebcAkf17FKVsvsZUvYoZAIy57u//cUhgeApIllCOYj15C//YY3XcZ+yU/u3UTa3A
jIXIDZ/46mxB2tIuKIPWuAmAAyi72MIAmO19P+Y5V7mfWlad0UGTELXuEtFfpn/Z
vY+IMFT/gm/PNzXfNc29JNe1xgDz5FbWK7VNB4KEYOjQnWmqFUoOBUvsn7iauH2g
4jg8by4duhLZEnBhcFWBfeJtxNCvrp9wg22+nB0mCDEb30hLPArhrutKbD5xNXYi
OnRv+LUw286ZCfXH5nIT7haOAkOYCQwnR/RyvpHZC3+fIWwuXE569w+X2oNpxFA3
5omC53A9RwKopgsdOrsoeuhSVFmDAK/IRwrAWt3EpMhzSPw00FsXb+xOcnrCEWnL
S+wT/87vUXE6tVN03H0K0fwjHwUeOiN6AYGsLgdP6pHtJOCOabnBpWWwhxhCn0P6
ohgSLsi7jOuOibRRzF0Ztmtlh4jPa4kfnGAfq1JyZWKJjZzAFNjRgQ1Cgz/SI6mx
ovinMrhQBccZva2b3F6/u4qs2VcfVLbR8nv/sVV61IOGlzvGxqi3/vpO4vMc5tRR
ukBy1K1Vks2quzrYrVshPfDPNVXTrQ0qJwHAuEfPIutZvbFmYegzpxFfj5yRi/nd
ZkHbfDd9qlg+wFwz4G9ScdzLIbviGvxs9kqno2Btc1LS0zrwjZOxUDFx2GUOZTt6
T/Y6OnzQMWU1zJsq3Xn+ku292s9hAXHTdzkrkZFwT2HJiaXwgCWyTeyI8wgP4KxG
/Vxed+wCXYPv7dyOTZTNrs3NgsvIiqPJQnpMzE5r5c09QXCNS85owEp9ctWmu3CC
Nc5dO2Nl101eqAWIO6BYGyaeWwn9Vmz0q5ZgsIcrzed1VRGdH4kcqp6ASqP0iIGy
Gs1mfbQvFmS6I/rCmvMpwPG82gH2zUEJ/ekU3/qYVoMfhaKy64A0g31034VUmUNB
zTX+Jr4rklwrT7p1rnJ8uUq/yv4mMDy71eolsSj6I+n+vrpR/l+dqN1HoAW4hKMI
FA7rXihF5MHiAMF5Z/nkvNnywtoyb+v5unT7vtxIZ6lARlSQAl0xrPHm+qKXsx0C
tDX9KZpevW1qOLVx7DbX5BX32b6scFs85xPd2ocdIjYt/3tTK7gFkWkqWQ3F7XC3
19LKULHNXstWYu34jaWEc77MkbrhAl9X7a702P7XztE4P44dFaOImeVA+V0ERFC+
LFZgAYaHHXoe7n1TGTUS7qs48I4OSl7FKqpWqRdXNiS14k/X4X7LyXetbnmS1SQX
1vzEIImJ/j9wMQny5yEVaQ6eTVGB1f2XGAQxg0YS5ZlPPaXr1BcCrtropUf0gMHD
0CwBLsApIE+bykr+8lD6vFoRS7h/x/nuxfAJ16xXnq15RQV4dMYZC6xnwVeJ/jrh
j1+b3akEhjFkEodC2U/MGAXDRsnoVMEbdp838yQ8s8aQIJqRF95yHiW8AGqIl7aS
58FRr6Nq4ZOF2oMD6pfs9bNHUkYjCAhB33xRENbc+i23KuKIRL+XELV3tLFV7yRd
XboJymmxlXR/a5CXCxt5s/3bG2r8H3neUVtWNs9sAXnOa+lLcNjSlScN1ZGEBfs9
U1snkxAR0r3O+q2g5odDs8AbkjDgpzpBid4qR7UGXHIE7uSHEfXP/NLDaALytgZ/
hXzvqt8n7PoCTPtY3gvtzJIC7XBpkxe0HKfKmqXzsLh794seys+rlVyCiQc+TDvI
+ZpEXE1/u33n9aUmbm7psUGCjDTugIgLvN7/UdSxVHcajwdiiB3l2i3UdiPsyuE3
j+YSwEOOqyWWyRw5Zpbe79M4/0t/jTi3fH5XnJ2RSys5FSiJgpA+1GJFaWO4Knmg
jJPE+8R3sbpnFj31ps/7pEMBt8n7MJQC6EZQRHBHrojj2IROzhe5mDNx/ZKBlEB/
N4B22XuSmwuGFgKG+DeVk7Ma9h5/qWJP4GTgVea/qjEl4FEon179bjf1YY8ZLI3l
I13ofZgzhZAHj6EhoJRKsSxXSUnBueJN/OtBUIoSB+oIvs6n8iSnCuDP9wmI98oL
c0/WTXOti73XjasTQNy9AP5jwSfgNQSLHH5Kk7eX8eB4F+W+tf60EtZNDip3jY9e
qeS7ZdqSzhtPVDnrHSCGgxaUXCkfi/T0kpAamXhALXA+b2heQ2o7Klmfct25KGF2
Iv1elxPZHWzw4XaVDsQZI4aYAvoKwDAeDl/HI/Cs3SYsur/17im/eimTWRvAKqed
v0Lf1wxNklYxodYt9oukh65s2H++t51MOVikQv6a2jSxirGook6ocwIX69YSymIl
8PHaxy8eWtN00yQy3PtmEczMpsrIQ9BDIAsYbp4V2UVihxtiY2wqZvr93Ad5mS7v
b97MiFaAm8l2ULUlMzLZGuUwdJuGP85Pj2mbWenHX9hbWWx9g44BCu9KEHRmjTOF
7DihEMHcNyrLCd8ieSS+B1FozUWVbzC4hF4mKNLmOTGUUkAySiNY661NP3jBP+81
j5xd25eVGQ2WIuzAM8tIzczOneiIeLRF+OzVrmSkcIAV8i7/y6hIZW+Y9sa9FGiF
nCzRMQbOX/9G0KLVRMltLJq9gtYOwYWljPPQOIBAboq2Fu9lvEVzjDJ99JZoGT9W
Sd5M5PLPcA+yEUfpubStY3ZxcDdvXOn0qldh8znJ7hACJr2T7Lpw/vzfNcMgc0lk
WRQfY7HylVTmVwbBx44+pX0lpCkcWOY3HffoJ2Wp/42He2RSnSkFNe9WHU45k/xn
19qXC6ejgUPLSx4le9HiHo4om0qGlbhWv0z4bI70QcvdeIgkW8jtV1Be+YkV+RPk
2c2EOQTEV0oSxZPhu8dTGRKLtoOcgvqR1omznYmtLjDQm8MQqgtq7IDvRb6xZleP
qSECs+iVU20pIVtM7wRvjXUA5ii4GWULr6vC0bdMZjf2fU0yr4Dv+mNr5FB4AEfB
57LdReUhKD2ER1oFmvm1emLdI4qT4Jcg6RXzzapck8sdeHddgIJeeqOCMAItMbff
EZhh3hU4Ydl/UIVMDH+SaGgvGyoBxbQwBMOuAJtze1+6rGXdir1EAjFrezJ4eDrp
hSFx4WGFGvbgVZPZllBqnqZlYx+g7TMcXp90NqqytNcLXaYQNIObV1hP3F4pGgT3
tZlmhfpqd571h//bo7VCrThU0lx8qB9NpuwqFog5dbv7tXX9E8xTS8hMQAFC6lDz
WYdx18rlB/tYUrxNI+AfocdB9EMXa1kTb6NIfehmtHRDgRBTAM4mQiun6cpUqrlH
SQLFVV2zOyqj8YxZ+KAdiLmxNynSScIa2+S148fDiBhXjK9zsj6+lbF1tM6xS4lP
Fm5tmMgDLQFGATshhMNLOXPLCvendz8wDjSgtfIvqQTliImHck3UOryhCPnl9IK8
xWqb6Nc9yd7C7YnDh2PA8PGRkQ5bb5wFSCUMLqMWX+Yl28LTN9M2ePcJ4dk1ol30
Jr2FxrQFbBQ5b7S+l5IOlpWfBYkSMegwwJ+ZvNhYA7hj2tg7H8X41CJA2bWCtqV5
M7pJTmZ0SMKSf13LykGUgW81YmOtIu+hHvUwIeBSF0krkG93U1EkW8iLTW9S4cxq
tmthFinbTF8yXxz4jGiilLWhS6SCXZ3k0ZRTAQaL+a0fJnEPVylnaWL59pXceEDJ
D1zr+G3uv8rBtFocM4N6qHYg6QRCXNxgT/8ih/P2mpEQWHuhbD5ulXMBU+C94bJN
41hOteZlqI0/iZQb6mDhRrLxE6SWU34N4lWvskwzelsEf84yu9WV+yQjSv9C6VUK
4u52mCd6OagPiPRQkdykEPAN7iKWqxVgBeZmSgEjakDODiQ+52iO+w6MJolVuRwK
IU8ATzrZmNA89R1eZUzsAtj40qAogihShAgR/wYch/di2g2HhNPyOckh+GDoMD6Z
TwplPcIS0w5WrYMU2IsqZN+yfOuSjlKjIusfhWveF4dL5l1Hay1R2Ix+Sqeirj0D
REEcVoVXzUX+Xp2MCdZJtBdPWgmwaCmlzfPD5j+uLfPhukoDh4ngns5J56iOgAzN
yrINC+1ll6n2d0GSA7yrpKSRRarwYnGRs2GcFbDmqMo+5mZwEKOUNyrTXWkq1qG8
r53mkdkTIZcgxrsmPQznffCfPebO05fAOXixQvWr5PustiIW9pPKK+RLW15QRS8G
Y+lfpXT3cvpca/kTwZiwpocFk8oKysnFUITwMzRGWleMdy+KD84VFzoszm5pFgTN
0XgoqGZ2f4FjbbSqp8VVEwoAuo0uraJQO2AAR09NavEKy29ugT0A7a1diIk5pN1C
KsMvvy8do+baz2fDGs1oTHuktnvviC6OGxcjZDmq9vyO7b58lYDldR75sdrg/X3T
P7Q8J3tQmk9Re6HF1PbR0mRHmnvU+V8OogmUYTq40h4qaVAo81AS0Uoe3Fq0+T/+
//W2uNyPjbZyesC7sznTCmTSUzylZREjy1MKabfhofK9UgGtJ3OdK3zZFYyylfU2
L7Gq43sOamcYz4Lr+dX7L3BnS9XvuwxMiTCL5/wFK2cZsxNhT1Jzw/AXMsWyfhiK
aTNiQGkn4RmTGvT9EQexTtHlJ4WdPiEBggsrvI9v/OLxjrqBpSKbjMDo+jyn1LhJ
EamV30taaScpJYHNgscs7pjLxQ1yh5/VJLO1befnlIya0FsDCJeVa6pfKXMUSM4t
9906vyooSXzkCBfLjmMbqdOwa8nJd1uOxfTYLbP63kOHlo/+qESggNkgt4pEK4yr
9ed2d1i4sTBPfNAnin6nrPdbqVOeVhXd3y6THIwnHA+84pW/xEpjZAGLisguqp1q
FWoBVnueV7n7dHp3I995MfV2+ACZshzCcw0Vbrp9YPYYwDaZspbC4wBSKmvqXxJn
d5BtJ62XZwgYMVvwoM//pCR2BMgc2Z36c8iEYaAIdRBhcZDA0KHoGjTfI4GH3gfm
gnhJq/WskNrREnV/s+gtg0+5NWKNOc8tWnS7p46WLz497RtLPujQ9E0X1BYKUNhL
BPyWd9MmDznl/ZRDyIiBpSQk0hDmDmOP1QNM7E9REodCUeBo1KdCo72pboHSe1Bx
b4I3BcnjJjySR21Pz3Mg+wxAM/r0aiR4pGegSg7sKMXAm0umsCqpdIPDDhEqnkSn
mqkCQ90u38Kzijh1EGYKHIqdzsrZQQjYUXfL1ASQ2ax3XYCjOMq+3th5cSqUzQXk
azvOTb1u8z9xparnn+Ztnz954QyxIXxMKXVdx/tZ/1T77OfwCrTZXEW4EP13Wh/v
biAaCxK0BMtaD6q7BIVEfeWeCGooHLIEhQ+0q+pDmNkEDG+m1lMPm4MFO28y0EB5
e2pB86LbCWbVpqQMCpBKEGRfWxvgzphGk9Gi6/L+yAJDcnWuUTD43XdKOxvT1HD1
nXW8oH1Q3PGYov5kvKqvwmDr7PPyI46oZto1ruOS5U5870c0DPl78A62DggEmBML
U29FRsVSEdRZUcHQe/wUmcO0izlHWm7xky08MWaNmiJUAdHWSXeIGg4n6gmQrrhB
lyV+pVNqeuFePnIXmNmC6JZLPyymGY0XwQB82a2AJPue5QA+Jl+QbPxCogIkStOk
C9gF+EXQ84W5ERgEzmteFRxhg/TgjM+sSCMPILv0H00UyA8fWT0dEXMZ3YzdktJ9
eAy328zyQJc/InaPfAcmBCfZLZvRl3EV/jDDqNCT7cMKOsS5KqQzu/HRqwOj8/Ev
dQOy3jd/2ipXotOSuRpyHEz1Po1ufHF+YdgFkC/8N4EjQLDIGLUp7vqS9/jesj30
owN/bdnbK/J/E18RAWNPghpDnP2soYitj6Eb3JTOCiu8wVtazkqrXCaU9HTF1/sV
KkklrTsitbpraTvSI3nBPvHWtht0qNlV3ds2xAsAqtuPKFfBHperjOEPhQU6lfgO
ZK8YZqej9zZGNwuHv1AC1DaxLDMoCUgKxjGx5aG5aiJJklt6N5GrCnzVixnl3crK
VCZN0gaEGJUsGgCk1wMOsC+4OZWDRFKduYB3z1Xgvploip1JmNwADnMNO5K0Ze8q
LihodJo5CvFqOngrsGU9E0DZScQa/v1D225ZU46GouGbmZzy2uLaMV7Zd5WY7Szh
2BxrHy8ZFxAHJevHAr6rA+L1blIMVXURfb63U2jv3AUepWAEQOkTZpLQbw4fEFmL
N++uSMjl4B6aPXlQFpmiZhV7ecf4rLEV/ZGa5UPj5X+/fxqjA0H129dg7hWw9jqq
/ckKmSkaWH/Q6suJAmFEY6Qp0hPJ3tIpCuqGYDHlpVe2MWyar8adaTwlujo44VcQ
hictZkN1anbjBLHNf6F7T4M579Zt9hfKAImXB1Wa9Sk4lXQC7uoHM16DyzJqvF6H
DOml5emZLlVzGuWwabVebDWWCnSCZ/g2THdVd/X1wHxYH5Qq36xDUg+exwKj9i2t
38N2cXK6ty938QCk8OFjF+5CiuLUlrEjknnG9A1luIxo4Pe1ENbatuqAX/TRY+Hu
aPhNpbyYYJjL9gu+UK6Dbpjj9dD0OoFxAfFNQP8r+0LeniH5mPhCLrNEVYrFQcgV
JwAhl1jDM0Yq9eDdtZAU/7+1Rjy0ZlpqTIsrzjqKZbjHfaaBk2ayS6NVwNpl/71q
dn4IJ9NyTiOqL6oX7BuChfsj6poAdCtuyclmaq9hSnjBEERhESxOG3gY0YmgkByk
3+O3xOFx66Y1gEAjjiu1YGZAq9HIlBavOa3v7bcAM1w6ZApOd42WAhi+NMdUKYfl
mCIogZ3jBQAQk71iEyGTs1I/lslScxJRxja3bG5Cm6ZS5wTLFPmBLF5y4MYuHv8Q
qVO6BYQKgIj43ROTVeWYpKOJkyxI/lCAKro4m3J4H7dg4R0BG1/cDx3Hi0bGtIVS
kuDZUFUI/+lciMOH4I2r1pyKNpiTWkknCYBV9xHLZL8lgQbbvBuYM8s1YBdw3gkB
KlKGaLGi9RBdjkhNYD21FPSGVtf5Q1VadBYmwPf+P0qr62k8rS56YhBgc31DdUeA
A908pRuC3dPnpoPbF/+L0lDppifOudm/IA6dnDnx0AQ08mRCnIKXKt9IQvU4xucr
492BdSKOhupeHKkCj1X2ioPvhHzWk2JHw8c4jlNaNiaVKgQG5q2WZxB+6pa6QMvg
rbkrAhyJ6/KisvecrxcGkBwWy6ioa1gBLwrqnjrtwbpsBXjD7hbd2A21VTJ8rKKC
ncmsuHgLP0zCFkSHc6km0QYRQLlVD0c6C32ZSecjts7LbC7/tRCOk9nolFlCzknC
VKw+5aiuj4xXqVvlSsdjqcK0Mit6wtqSKA5YETguEwGsG8BoP+xr/G9MS00LbdFP
aMNgXiJmkNKRV4gKNjjE9WCxj75fqYFaFqziGFag65DnC5Z1Cl9Xn+5uGFxK00/u
OrrvnOjwfCk5tvSyL8JZuao4U+0nPvppkPXA66sM39wiqpuegl2ZlkrmFKpkN7G3
X73P+JoCsld+S6U6Fmx7T+4fXRy6362XpyH8lki9X4BX5Q1iwuVkitArVKDhYYQY
WU3lldm/cSxwaVSO+6gQpWbOBDcx9du6UQO8cvbksKMmdxSK6BLytalgcS9ECTrh
Nee1DuXaBUPerh3j+in5wXnM8CoCK/wLvoqd42NbErgfO+ptuyf8cs1deWSg9rYB
PNyAdotmrlE0QpZJOttWyV0ci/+z+5K0dyq/ksw3PlEHxrPGdQ07xdHX36nEHp9U
iJjH9JvH0+tXnKBi41hPdZTGLooBP/ETz5DB0sYCrHmuTDhc9jO5OhBH4Fn8E+QP
5Zt1oKvdAYRzYKKk8FD2m0E2a2NEYi3rPiSkkYOQlquMxpRl1YPbkTTQLixzHQh0
zO6CBcmTktRweCnz6gztjA99o5GlHv56jc7vWsvSr+Yd3UZ/IKxjENdQzmmUWBd4
aXSX/zbrol3Yyr6wlDXKs+RcR+IYrtmNlkpp0nrjcvcmc6zWKBpu/rd1cciQ+HbT
KCg0wHKbly7nO2HFHlxWyXj1Lx5aYGjmun7I1QakkkBskvKj63II7P1/bknq/QtX
pXcGhN22iPdNKt+nMkhmLa5dIFEAGbOJmt84Z7XEbCfXM9UN9f4kVMMjyftRQQfD
qFPPgG6lnQwGXIMMmU0g6M9arfg4qfw+KSa+5btlx2kaFs4v2pV9G6SyktEtdrXQ
JJz+1WuqLSOYR9bLCB+rPfRWJDPQ7hGoWpiNIqGaQaTDrmYohfl6+sQhc4c2XkJp
MFILjKpYM/voClhdGi104gVYFvULZqewDIXBJnqwk+OPSneBXiNsm1g8lkNWoWJs
xIh87WngNBEPimvoDSGe7a32i0gMH87LAti693ky3gRi8HEyT5rvzlvxo97M70rv
ej95Ehst7GRsv7lGrv3W5bI1RuKF8KlTbYBQzVVIY96Wh12dvDuRcpMGfF2Zazn6
uGwVcX8HxQR81IwXpyyKjsPEjOKeZOiZJ5YpkDqzpRPV6lm/fmWRfZPbcBol+odj
8sxFQdtyYkIXKb2wYU4mW8PD7Lmz/o626/bCc7EL+oCEnd12oOCw8ZW+EDMPcqbu
WOA+4sPchD+XUCExng2tTUx6Sb62ynlqmmaVkqotrrjB9q/G+ovP/fFQ5bHoYMSv
/KwCQrHw2OX1PhJRuIzdw63sLW63sW/3NoNjktOqYcc8dgBghAeeL4xwVv2G8RSi
afNcNu1ks5ZLmgnZX5By3hBNq1AN0whVG+EmmAaq5icAnidllbl8HqYa/OcLpfKS
BfJnMVtRTAjWHWJNBzNh3HbGfixtsWyMHZ9/fVq0OFgkJkGfbq36HM4UvV6jsTq1
Hlp9vT0n9X9etJhdt813ULPeHcIrSJiY49I23LUW3v6Jc1ZSjsTEgC1aZpvL3jyk
IGeKNpeD4X5DsSw51lsNed28TP5fCXZ+LS0Qj1QGUvo/aCxzsoEV2m3iLAtJmob0
NGCCW1Nj7A1JujJLKBgEPjZAsntX8PM5uUYQYE0buThSN321pcE8rzzgOqz/xQsr
f40dKlIfhSKgChqEc++qaw36g1XOs+vCM2GkdShlxVKhNdUIkVmp7dCnfNFgK/4f
VlWBwydVJYibKsDiarpPExZ9+PWCxKJXy2Q1vQmVKebctGsfU1WK2LSM3c+2FPdp
ePFvp1DC+ymmRYnGjvQM/u4ES0mVZywmZlHvzMfc3nS07dqVE1EZCETspzGWK1NR
PSZFZo+loXrSTHHSltbXXA2U4QK2FTUhPy5hcCTySW1aumux0LIrvlIbXh4Nq7vx
KxAa8phIVd01yYo3hx3vLIZbXplKfI7CLWYAj9RFlbBn6h7d0ZyAbugNSN7thJGt
rkN2kVJ/IsswyG3YpSCELdeCY08op4AF8rrNIzLH1bHTez6IeMjdc0yk9RF96Fml
vjQZVMe3Us13LQk08BVtsrrv5UaBFJ7P3oQoJ3Mzm+gYSPPDk53FAvd1h6Rw/8wx
hJvaaYZWpPOM41BfyqPWD39d7VuykV5XRIESVpOaEC9JhiyypxmE9+12ufJyWDNv
UyElg58+/fznSsLKFziIchhAbUyAzkcJ3cEyQSa+F1KsR1W2/F/kj18UPv2zKCja
OGRyWBvv9/7w6NlWSLCPo/0CjypdFTtycAM9bYDQ8K/05nsrJCY+CRTEl5Tota2E
jHiY+PmbegSwTgyVk6WhqX9nKv7zkMKFD3NLYHbXs+NwtcaUQ9zZMgvkpo/FNgb6
DR7esDLyjUU9qUbYDa2zVp0acvfx5SJ9WRAee2D/Zj015UDgafOvtGdNqSWkCQ9k
kc9iXD1hqvK4RrHqxnLEXoIlXjdOQUlKfz0sIIqTlzJmk6wYGDxiCdJv3SQhHyaV
qlM1Wi+rB8ttRB+6THhFKFX+VURHSfwIi8Cz/5vfEy4a/WI6svAifrAc1x7nkTSV
NI2MqCJMrWxADTP63Om/kEkzmw3hlMtr0GXUQXKkO+oWQaGQNqko1MrAYA8UuVL6
d8ZeV2UPmKnQ+DLV4dHb7jhzdpBOmvE1F2OHQH3yNIaSIBw88gH3Zs4KON9dJ3uF
jT6C2U4mMxG+JZT7mbtv0zzKWuvLOiXsHCZY7LNdTPyTtb5dybEedZCuUwoBhseR
eeodZhKVOCQkCC7aT25bctsg5FQA2WNXJNau5UAZLVxsyBVFYKPj4+T/3Dhu05Wr
lNl6tcIhV61oKok+e/1ZPa100BIuRHDjjMrHvTbpvSg3jfSPCDB31e4gNS267jdS
TjDBx2irr/rLCDMsN6WgDxq5+NhsR+1jWDMMfYH4E6L6fTrbxImsQbce2utrMeFi
Y9g9Akq5+drZIxPQVAhT5neXYPGToTxKpW+oeFvY9yLEVWudH7LyNPIbMESJvC80
/qhibbm5ADsB8HHsy3DMJUlcUHaTaalxlsQTsLImvPy0I1JgTq4fPZAbE68g1Yv5
3545wNUnzGx78a6AwHMCTybT2svlB4LBj1CkkuRqRZnhoCzB6br74St8HFEyNI+8
Tm7vUEA1BW8+v4dMn6igq065swFSEceBbFE26fm4ptMB3RzYUiHFDTWwhBWI8Y2c
2KtvVIrrxEZC2v41xSQA/KlLYQpe3qoneDxc9vI6fAX2EkpUfy7p2+ANI45UR3Ws
IZus10/rdq6rrQhcwWpwKwB8LmtQcbt7RaipKVBSBFfXPSIu64tbKMkBnR6zhJNn
++GpIx3m+lJycVLOFNnAguvN3CbpUwGCLsVWf3YJAxZum7b8J9fVceRwymC/3pHM
spuDbLoSMXmvE20xZt5CrNT0yum44ZwVdVNLaIrMDFh1u+1/fWKTlh4jlVJoFucB
p1tE7vZ4YjhwH/EkNThzD51i4tfRJPaXmiF5upe4nvSoJe9vUA7X1dPLNI0slf56
5ajUgLrzw6riyWDnrFtH0adsxGtc4cbmgLnNq3hqPTIVBSbtwLn2nPTdwpa8PfWQ
oRvUwRsMFxQCrXlfMe0dtux2p4qIIebXJKWmjSas72hb2OM1B4rnXjaQ1/z4zf/z
p11yaNQxoNKBT+lb9aNHD801IuEpkOvbQLW5Xt+SrfS/NPldb+Ol7O1PvMw9cwyv
FqDnmIizLZ3L8CpCaq2vfLQu+8alE+TQ9jhIAga5nrPEftz93yHrm5zH79UpWICT
IjsTK2UVYsIIH72lOcrPWPI53WlrK6HrsGuV6nqaU/y9VGFy2xjHJ7SxyE2n/zJW
tJoZ46wKJM2XQf/ou4jLwmhjpRyHY6vSeVDQ9IjATKjo01VwuWXRljW4U0LCYUwm
x1JEz9JCqrdEz+nAsx1jueVWKLCXkt6qSNVdLAkFCEiulf2PEFAfLqXOrjn+Gwxy
E0VK2C7K4mlYm+KRUHo3/gPOgerAhp5MwdlRIErwL7Kv46WGLEo9jJcWttiuhQqS
4iWwKPudvfQsbdaISpLNDDsfQZg7Mj8cLegVA016MzkS4RbcyfKsxfNykUCkjexA
2fT/jQIG5ga859VwpPdyldtmU2TUDD4I1Nq1Qi5wfvxmmQHQDWKjzHmliIG649XJ
5h5fGLsxgG5ZxPR618csuIpywvc6jzLjfxafHNgRBZuY83kdIDELUHWHU8tmiLxO
2k5+v+tvlOlw9XO8/p6AjAl5IKysgrVU9EK0IhR6UsgopSqCX7HHyaYe0TTE4oB3
9M+03ZVXWVBENkVpKBg57VZWOFjmfCHQoSWCjJypZxpz1hZ+//sf2TFXiAOvOgt4
pYMrKsLHoumEFDzPYnN6ujh6k1xh6rRsq6joQoTLeg49ScDXGJNU4SOmk5B0ROEy
M0dDT4RgPTWLxfZ6SaiKQRQUn6yY7Jgm4RCAjq3I9p5Mf+KEMxGMx0bth/i1Xouy
pwoAV7Y5MtWqEKtQ8xTbMcnKqsKy8KHmRvBS2+6otxrSNwky6sBkZzWEYGxyvZXG
aLWHBD8L7WL5ZO+3sbvgKyy7qn7LKbbJQW8ZfX7DenwSBjWqf+tzNOt9z9KT4Hch
bZ3p9Qmc3B+IUu4ZArLNvK6kcbZaN4Q7hmgF1uzTVIYL0//uLwjThh9jQp4ld+9X
qpnWiqZQAjEk/X6krzhC82MEAwi4sz2eyF0uDY1M7sfVSJQUa5e35MTfWbuLfCec
DKJpGaQ859OCg9xF6jpF3btUMR/SS1S+95JxTwJtPTuA8RzJZzhFBVVBCaAsEALn
P/sHyk+80Ue2FHuDyaBnbqoMWM4d0pn6j0ktTRp1tIGqbDrywwXv1t0ag2nOhCga
Y4g6zTqT49LwfpGT0uBejK1An1YLk+RMqeJ97AGt13lcv+A1VFhiDjuhjjIXRi21
/LinCqoJe4RaUJYpNrRlh2cH7OqNPWOw9fFi7g5pPU/qj4i3Gld6YkaPfcXoEev8
yW3uBIU1qkQ+K6GVVnFvXSd9/bhETDMDfbbPRkd4VFuMoZf1Np90sIXCvJK+ypRB
P/keiyRAUoysZgGM7kuJ34V4LI09Fh64ST1wvph0LzjnyVNBQIhdKcIxLjifWOKd
HXI4LksbZ1F46lce2moiyhBTuvrCRZKDC4JOcAg9JrDfKc/xvAZdSf8nIxjPiYp1
eh0DLpLsMsZkWRdBAflDXcFQR3//fRzQGQsH72a+efRjgIJITch2gBAm0UwksnJd
isHZc2FGL2xkSrPfjSguVTexZ+AysZgLe4nHcSALha932l6/Q8wxWRD3WinXtV9v
3o8hFTypQkLyPYtNYCv0zysMqB/lrxwu1B+Q+AEd82nyNqSBwBOI1a+ZxhOhwQso
dDF8dsfaK1g2cDDb4j12JEOe4rq6G3Je8RncLCIrxIFAz5QLjvUVg+Cn87HnbQCI
308dT5a0KzzoNTt0sF6V4DWfIFF0srmv3ZRj6oEaQILME2rEdfevp4BUnMRE42VB
qS8+3hj+1z5vdhfmkVzxSEKJeEFuhIlNa0dCUVm31hDU5m2walZgPDpnb5MfQdfZ
BJJmGxw+m19fVXitTrW//jv4C+4IP0glHG3ooxUEkDXS+Raqpgt/juUsBMYUm1eB
kfs3Ae+Rx0MQMUmT+YHE13zvtXxI8O+JuuPoqwIBhjVVuoQXYK3etiHXH0+t6MJm
5szCw7DSSk1tNIcSIw4PPGlxNQhPV4mBhqtgmUAOUMjr17LXUFbM+9LWPYuJaIEb
ta6I+6z1ub31e4RAyI6baEydwd/8WGI4YH3C0E9o4nIH+wpAw/NfVvjNMtIq/BA6
lmN4CxuHPNRPwlS8sLbEHnw95WLKZTai5yxmnPT5lgOY/T4tZxLrdc5DErK/Vktt
01PlcIPZBZwyTPgmIue1rouxCHZAGO/VvkHsmvDpyARs0+E80oANcCmchkZ3LgmM
HnNFKLAZim5/Q5XmfajPLgmXn9LxZ3RG3UL/YB+uyqdSyxeOwE8bvFRbfnxDGVPr
8+YRtVXD6OOQi8hwCQk6BlAJQrFfREP/ExTr+8cblqDfW5GkkO0W6cWv0OhyGqsp
LUol00q7A2OLDlQbWpv3RcrBXSKhGW6hczl2BBHVtNY29dDLWr5cSGahH5nu/Hh9
uIWk7N8okn2QS3RhSgbrzEwuaniLZb/uG3/WaKPmUyt3L/fN6t9xrja/1WZwvdTc
q2EGFSfT5Q9zAckqTp8rm+nH/3EUd3N2yJYEKX5q0eLePPaI+Jp7fmqwS4Xy6/Wq
eKump78ijl/kGrvEKnWebkKkWzwuKA2Rhp2Qloyuq2PS9Day8Nv0pH84peNDACmt
Vx5DNn9KmLT3SKK+vv1rB9iPoPJlqbUBN9yJmub5hDO/yA0iNM3KK5J9E3HNXynP
ZLVIarshNhCr8n082mL+vRYNv0dZ5fTHVeUaSy27HOcd1EnyVAJmemW3FIM8HRVK
/lp3U1sTB7CocjqImcS5LqXrPwb3N6lVxeke61gsKfvpzTkMyfLK6f6tRN+CU5+o
XmSoVdaJCtICHTvCuYcsEowf7ksomwZXNskQqeSl5rotAn4B4mfl9thSw41c8wfs
x5fL1Tx1VHu0/LZhkYx0GdiTt4QdxREQCqQSVgkJ2cZpSIICnUC6abE+fiji3dqo
FABGG1xYyQuNaQZM9GWXa1is6TWEk5+9Zd3/JO15iXo629kWfMN8EJdXZAZQF2tF
IJD1BOTQ4Gv4CPVEE+Jag5gJvFjKWEyh4b91RMzKO2tKZAUsvdy0qeF4n06VFX2s
v0tLCC6A8gpGtDai3IMxg6JSoLsxKNb4P06mOITKYUKrjDIgflnsEtgrqLP+N48q
zZvkVxnj/UFUs3AD8e4G9EK9hMPyrBULhgPjENQp6ZcLPw21PbG0uN8oopOpH+vX
X7vzhNJI9TUAmEuufpLya1BtDGUrp8OGeA1jeNkA/EE/oIpWrHDg7sQevp/uXYYl
v4t7WrWfXqD+qpMcRnKI419ODwl3cHuEtvFj3bK5nSLkI25+//Y3T5uiBkUvY3sn
10QTgqyNbxfH7st932UvK3FZTSCXwiqhefVvtuTxnhljjLWpX/EYNV6D3E4UxkL6
ECJtTPZPRA8k0d/2EaSamehJ/mm4EAn6jvOV400ThLSv2nL27StpD3jCt+EQZX8I
oXdjuaDF/Hj65xVteyqJ/Urf0OfsC9r/JjBHVS8QawK/YJORLLutsN0CASD/ZcE3
zU/i1Gzf4H/XtNoChtp1AaFqsBJ+ZnLFcAIz44VktemXkD3TFcfpyc1BVfoZoGJ/
b11/9n6OJlu++8QutZLrBWi/RdEJRo8tt6QecrjIqILrmCFQxue9YZEZkK1UWRo1
VMNpKn811IqPMlrvhxBzThzqWEMEHw1+oDlXccd0rgoxeW1k5xEc/WqQpBCC0i72
B2LvXTtPkxtVfROvzyAMe0MQfQDx6f35PwLOKVtkhheWfhd40uMJ3NVri+LScuS3
V7F3o3lYNkaSIA/XKEMDQ4xeU0peDIGHiUi8PN6JHYVv3FjXldbON8Wp1CjFCjU0
amcl7U+oGBHAn1+HmeBEIBZu6GPF7a2Oxo0Teq5v3PvDPbC42xu4nenaFWdCwd8L
tsQCA1ytJQz/1GdokRByRalqfE/DngfwM/+1umFbKfxz9ZOccmwrT1Pjzif7bSo3
UCdA47ghmBUfvFCYGbgNcmDqBnpn4KcVvgnqXSTyNj3Fe9s1/JX5K2KFaT200aLr
21kS+mMj1pfSzDWl3Ynq1c5B5DdYHyvUgqGvD7hIpaDkhRjQHX80jeyiV1085X2D
hPH23+bGEaSuX/WJJNRRuDAkcZWEllyqHtNsWe+D3koAePye79kOYhCbX2xb1jyZ
+epOVnZEFY1enKCvswWRY+4sf9BBs9HjQ9qvuBvsVsWmuRwz9thRZEdiTjFfilG+
pGcpadinl2eevBon/tiS2UQQjDwWN5uC9uGr7j4Xqm+QPvAqcSuHs7HYRv1pw6xH
QHXbbJWoWxAif1bvq8JuoOA94K1yJcZPmA97WMu9XBfSfv8hf71JzBvimzSdk99M
xiedRPYXMqdz2JWF1YEJsRk88z8v2SnZX0tw2y9HZbL/Cw4q0OGXiwdm/pzggVzC
1YkIy2XFDudp5nOqYX3KYEb1vlsXDj/Ov6tWvJb4FVKHx9gp/da+EGmtE8kTAYQ1
XWP2g4nkuyyHMULaIhKqJeTDj+yBKlZxu+yBvjF8grEo9W4QCvPmlzrcCS6ExZAe
lfbD8sCMcdVl8kBvEJ1K1zzYkN8Az7f94nE9K54QoSUXoviBPrdpbxja0N1dcy0W
YKg82nRDsb5I94fd3LfVH19jpmeMEwq1SqttqdgHojSdC9m5hqjL4NT9mMeVUrk9
jWJOZa16djRklGRcDAKi+HfmHYNCRbNMY1yOqxGeXjtKn5yZZfSncvimMol5pTT5
7C1qSTFGKojVByrzHRyedr9FfSOJmAbZfA1FN4INmyzi6w6gGy+2OggL6B340+7a
C1L0YVZdk0baNpuKUdFWPa5Z6PKEpCZMQBcLOQmDpnUTav1I25ifYTAW2CU80dXG
XSLHHB+HKRrj8xBlrFzdOfm9sxP0EQFeg1vZgV+pjJrADhhAp3cGB7Kg2AIUoGp1
M/+OxgGVnG9hbVeAGTNei4pX4Be5ZerTkEkcK5lqldJcVYd8Yn6sw3dbeAl3r56s
OTkgpVvfiGsMemMKHW8k9Om8edhYhhlv731n8lLeOEcCxv4Cj1BXXZsSkQgkpLqD
Kd8++zpDsnPDP5v1NkmEorLl9XdGtZq4O4xXHZe7YC6PuEV6JpYe94GTEeZggWRG
Btnk9wphLyloP9f59oeFS3P5G+cnS9yZEb/BMuqlNLGzDZt9yvf/A348ax+78bde
//uOEIlHzPZr/lILcvj72AAlVceokGryOxxFkn4KLafUMwmQMEh5U0fP5VWdE6Le
ebdNlLy9MNX4bCeSLhj3o3QpZQ7hGgZZUf2QQvYt9Oht8es0VQmdVDfZXZ/z8G7f
7yi6JG0hwd2PmRb+n3fnglX9gm2603JmDyvdpoKeOg+/zgc+lUO3OqBUsNdpKE+D
rPjyP3QSJC5g7K16EyHw1yXJoE580A/XfwGKyUCg5a09lZfsUOSb5BeDXCcxQ4/P
7gg5LomC6USdkoiF9CpYV00sorRMG6kldB/B3eE9ELxqiXwzmnHGlmY3xQVcVCgE
85K+HphZDnQeKNJyrpHdln+6ZLH8sLJHmSVuqhDEVsMXcDgtW7S8Ln4fwk84xcVV
DChFsywqhB50BqY1m6gVtrYBxZgnqj8/aMyQcdooZC/GSJVr1PipY0S9MgGepBrR
Ki7ZOLpaVvL7t24ZitfcGpNEr6wbpiCpNVRWZCum41ysQPf4M5ZzUGghll5l1VG2
KkvMBrTqSmEzNfQt3eEWYbuo1R6uk6H3Brcix2cO3K2qJID5PFJjNlrFtJGob4jh
PRbron0knxIaXCgjdiX6sGq89+UAxLVMJOMMdnobi/4ERQghQ9XrD8opv6/s0LXU
wyxJU0fdXkd+xiYwhJm78NAP6V5DZvS5DPFuZ80eY1WlzQEQfzoFj0qt+0/4J+kM
autKMgMYTMx+D5h4/5boTdt7XloJWg1r6btO7LY1WYlHA3vMze0ePF/zzC/xSWlP
huE0/q2fWl4p9c6qtn0b80ibNWbn0ld/Tj57Knu93AceCylyVYQmhZtwNsOgy8Ty
I2cmMtve4khMDWGPK40ZshFx0CWZ8+6QcX5awDYOxDb2OEFvgC7AqV9w7arVoGlo
nF6pGzegcqsdGHoXdF0kspSZ6PKesqm61fumRxNvHqaPaivkkPIKLKrxyyekbVZ8
k7AVGiAAUdMAu83NAfCy5xGr0TvpDQLcsjc1lsn8DXovKGZa19cwVrUwgwhpfBYj
JLSQZ1FOKjCw1ZqyFO/zpL1EwR69s97S9KHaRYno166LAOTbheSo9uv5QOncYqhp
VC9Wd2Z+aVPHBtq8i68Gct3Le1mV0RhuoIg9L3jPlVW34dmIrGMTBAQrdZoNv8Au
dyL/h3OFwe6qQdb0NFaC4AMa5aRLDqgcO4FtJ5jxhNijWvaxswkFNKShBGTq2KaB
d+jwP70fHM5kKUoF7WR0Z+khJSZ7Ay1MYFX5FwWjfw72tY9W4X+As3kZj8IT3sFy
PsfzPO61mQd2izRAsGXDt4gbg3SdpmQTzeeuNEjM13SbF+ZwkwB50+1zCf8cJDxz
9Dmjmdqn19gz7z0a+qZDF9AE6rk0htx69MvjrfKTLyIsFJ+jYmPcxCqtIXnCrCJV
TwlBqzf9ZzVqnP1ojUUqPE74BIaj12f/GIlpYIrQMV2OwQNy+OTDphPVbkzx8WVL
tifqQaBFuhURYtQY8IWOpDhfCCsummbfBZhyxeUQaKtgRIyY8fG0EXt6a7h3cTG+
/l7KL2I9GA2xlUfowTtIGwkDkJoAqD3nvc0oJKewYDRV1atAhrUKra0aqr5qk7Ch
JKeZsRZX3sqghamB9i6zJRL0r/xZysmkoJzb1VgTdTmhGR67z/yi0y8fG2gP2jzK
6w3cVrcWH0MeERJaqRp/Ex/YS1T8Aky28ZMenI4VUXT+ZzE2Tii/yvk9zmbOENZB
mDgfam4tWb0s6KMddIMU6f8PAQIccidUVyCYJCm+13lGSz5XFD2luUEap47Eyj10
bHVkV0XtaDTJMn8Jy9Oj/PmSFfsz5TOICp7hIPOFEgaOX5KcSqIG4rlLlmzitlta
59wpcN6r2xP2bbMyZgdnDP90ZwdTH2zMG651ICdKWJu/w+AR4xLpRyuI9ax6Agpv
ZsjiTZQbejiA1CJNHBoAu+xnAr0ey79dz9x/EHEN7im7J5SeWiCmfBaBhSLg4kzE
JO6Ti7hIGqXOyJTTHivXqUdw16UAMjizfZCW8ruejd5ATDhndrPATuFqYM9BPZL9
kyhtVNz/qNE85WzdcI406hTS7IisNBaSwnd4EauuB4tvEygev4PdQWu7AHJLGVxM
EoXfmGIE38g4jBzmdbpw0iOaG2pt/ah9XVKqnS17vdM4CEVb0iQ6C0JB3rNa+Csk
ndTi/xSTQmjsiQFNd8APhf70dFHPI+5OKC6A0lnEoBPBaRtT22Lz2a8alU5mPkSs
lHfGo87vwhOQX9KH6eGezI3KfdDCqv4oXb/3YHkTRCB6pmzH3tQOCpH9A0GOCatE
4hN9WKAhceGUlz2u11YJBd7Mi0eWHNNLOWwmoYBLpu5o0mvaYwjti8d0aabVczIX
IjmwFi2LdVXRk6RfBWi/7NnIHx8SDqBH869dn8y2evGiDInrK4MpUXKjvALZ+vVY
1jSNx7ByKgtkikNaRDGfWSKYm1CjiQynQ9OvW/xQtRvFqv/9kWT0lpAeoPl82H/2
eiH6dvfcbVzToNqa7GW3au0VLyFAPBsZgjLVF2sL4YIkOvNB6Pju4j1tY63b05qK
l8jwALs5e1mls0RrYBBdltEtF0hFQI3VcbPwL346KDArb5jxC1eIB3VbAVHpXKh3
apaWjflq5VNZvMG9eBbGvnHOjaOav/v5SH3Wzy6XTbd35qrgQ4jUXLBcVlBkVB0g
Yfh9xM7/RUAw3j5Y0azo3pkbo60qQwVjJxWNcDCCownoGp3nVARTkNI04rZqr8ou
fIKqNCFFYxSqsacH3/oSIWfgFVN7w855h9m7ZoW2cpkFyO5piOsDMm38gtms+Hx7
r2w11+1SRxEDIjgyfdDJoSpdjg556upNCCnnA48HaxfvEI3s3bWjCxiriLcNTSre
669w+6k1aDu37MiwIzpyQ3fZKEbAgMWEfQODu8eZSWJAtO3ZmlxX7A57gKSKACOs
eg0CAvwDCxA/rh/cs8nmbgYVoSC7aDDnN+JXwXW7SqQKhx9VIkzn5/dtzvcsGh8B
k5LFveffaWFKdniewjTlMUrgrrylpBl1J69yH9fTVhcL/2e5HTtLV7cVfbJbx8Wx
ST0FdnV+8/bpy6VzSiltOYg9hejXqi254Mm2XaySbqkcLgTad/lo6sTxU0zjg0oH
AQzTFoiGXoyph7AIDWVuSU7S1e3aFIH6UEzC+65rtZwHGRzEzszgUV7NhPAf+rur
AgyJmvGD1rZdXVXi0HBm0Z7oVCMI+jBTDlTmA2v8BlfjHGTEJ8NKpHU6QQj4PwiK
VJEDl1L+rY2/rfyHmXkKI3t9au9sFEDPOK1wMBgwj7G/yMHuM/+e+mDDzT2TXZtp
Vb9qaeYTCjUVbtBmIhCBXxfuBNtPzIZw1OReEsx/IGeUEpS87yPFCZik+tb2dLyO
T5b4xkcypFotoJwrlGO9ogWiuZ5SMn2pK5jO5nlZzAEBL7/V4mqnHvgwvCiKGeYC
IJsuulVnwR2vkQ03RFYPidwE7fUIVKqMmDFPK6W/y0iJDEV3VDDNs2hN6KscGAjk
x1kx7JztQaTg+kIJSeCn20ph0jY/hNb/FnOfR5/DOCqP6hBKvdnsabhUB6xDOCKE
SDlUqh1nc3U7Iv8NqGew95okM017F7x+iO5OjwpACqA/th59kZTA8nUfSY5qq4Zi
r/a3g5aTcGySEzJSQiq4gEKqBwGuN6znfPk02tb6g7BzMNpuUrW3kgwdOoGq2C2t
nRorSkt5L9RthehjNNfks6uH9+N+sS+3R0NYd1jaDytFq+eP9q9xTDnuc+33KkU1
ZXtQGiaveBdM6CBt7nobZ5R/J8VQLqH6JYumv3dTfHfFdSDMLONa8KY8jXL0Z2Va
6aZTZNtRqeogqR0nAKvw2CnOy95+bgYZi595C2cDKjhEngXquhJpzH0NAWmpPzqr
bpV/7fgKuZNOnf2vAm3+ohBBSj0vhEJPRbK4rSvOkXKcBmS6cmQS4QuTn7n3XpIw
ZqoAJIV2LhUuxTt14hNEognrRvABC+vLklyGTiGGByiDEfbOvwOE/H/Jxq6Ye8U1
81617oHJwEMHWRQbyRmlyH+1fYDfbeMZf3abRO2tRAcQ7ekADivraNHKv4mxLH2G
fJW2GmA/vPSyEhAHySNZbNoVDi1dH89HrWOyxghkfAfLHdesrLEJBE4SJ6CphX9q
nINxmOueXEwQvPrcLQL1BOh6s975C5bX4e18UaWKSIjObpOcHeEhnanuK+L3udav
ZMLVvVmJ9Qe8uejf7JMnV6kgb6HZcEv9xxMZeDSYRceOjMaJGA34Cp9Op4XdXEe9
Krhnxd1qVm5M0chlXriRKrcFhkADTac7IEsI9Pq88M87PTjGYcjpGBitr6E+YajR
Sfr7H5TdgN3CZpzv7yAMYhzw9wEzbk0qim8u7J+ldjZl9TMQi0b8SXWXXIy8Y15I
zyqU4g4ZjCTb7to0QPwfZXULG9ODX3FlWwGIDkfdkrFXveDVmUpdTemzkxKf7gs5
KNTpa5gX+OA3CXHdtBPDDm+pt71kPwYSpR+V+WtddOzEFH56tbBMpF+hNLqO67ZT
aJf1lYggHKpRdrDYUysr10H8AW7yIbngYTUh8oUyjGY8LfJLm9wT3oTL1vc/FRSJ
+aBvQJvmEu9RAkw4fOPoiRjm7AKOrETNIgTdawvSfvKPFvJi14/EYCqm7PWxByO7
C+UBIfSIC6xl/p+Zo9NnYlm4Vw7l8Y51uGGFf17oWna29yj3xzubipzIaqjoms/U
wfUHqwMVvytc0lPr6+478X8mvQuu3i712JW8YdFfdP08+TmP9YqzC7j1t5L8j1mw
GgoDOAAYfSxIZW/VDsE6Lz7HRE+rwzPNXReslyKoKq0ayqrbF3LWHDrek9JoAnpy
9k3GWBbwjyd9NBl4oDyljkM3oVtxKojdtPSyxbQGrp4oJpk5JoIbR1bInSRRV2oV
rUnQ8JYGyhhL5VTJjXSWOvw5peIfq+lc86df3do9uxFvEueptpLNDA77hIFlTDzD
2FChFxUzROuSfajS9VlH+5B5ImlSfPNYI/ZtsoST2Pa+ppHFV5HjO3dVay4Pe0Te
N0LCoY4FtMYOKClv9AOnW3QEx+4azA0SUslBBj9AWGIcGBNw0kAgjaizI+gQgtja
Y7SuyrUkDjYfsrPFGRKKmsgrAKbtpFbg/h1LxUH7XNaloahzAQV22GnYHflGrAtv
1sVEsKWFOatrm2Q2xq20JLoMNUv3HzvwbRmV0pAF3hnCWp62bxXHQEWakJ5b1w9C
D9jtQv4hOJ22VUtzzmbz6Gn80v5C+OW9kcIKjYJ6/mGCFPXsze3hpzSsTKkV3U2d
uVoL6kIfCN9ZQBrk8yRFXrCPThkM+xaoYgDX/czruc3adiv0xyinygg3CUXWAWEI
KguX8tvNtyxzsx1JPr1/wBaZDW6WFRjnHqfO0+HdAwU01mcffsrgFCgE//2by2IH
MGbX0Eq17CDxISOtTogm0zuu8mqiOEO2lOhi5TaGImJNNcj/V38lmc7Wh0mQIrO/
l0eBAJHKiPTbaYd3fxNAi0li65eDlzFCQ07lHGwzKSNF4obnmVnXYJhlXLB1RBfb
3jILN10KWx6bZHG6knJ1EO6TbaMDycWJy0+3iAZb1TKlgRUHiEyO6gB615asEy7e
0ehtpTu9oN77Xr/E5B1i9KYaIRHNO42icGu0/dmhaVqRNhJixhkTNXqf3Q6xhQGE
V1z3Y9jMxOtkuGQJ79NDRCVg4wGbycDaTEUSbPl9vBndHQjoNynI+SG9WigGZ813
K52Nh/OPCBgdv2lXflcb9NstFu8Q5GS66f1V4kcMnbLKvLIjzc3PLxvsGdCPxOxE
lQIQ/I4LSOrjhX8//i+Yfzio5aQZbsg/5eEtiXUEQY3yxMj6O0uxlJTMLYMDjd0e
LppWGEUr6cZvYSCwjLC1IReR9fBJnCDGU2bRBhGDVi9UxRvUjiMQwCMrKgLE9h9i
E/uDDa3vJ1i/drFJlv9P8wjiXykvC4c2HQMv8tj9NikCTtGDG855w5oD4FZnHcRM
LFz7KarwYKFnyfAZq5sCo8l5r0t+67RBhKZ50Iyvast6hTKvlKub4DY37654ZzZv
CiOuqqIYt/vrwEjflNSSxEseHQ5tB6DaMWNSjZ4mWaXYlvYbY3PJfdmupi7ctcSt
2KJQiXkklTKwUSmVNngr53LLfaQie909uG2u048DgExkidmhPsN0yJQD7a/6djlp
mChPoH13DB1Q0ZE6PXBa2EUp9Z3VrnH4TXSUhku4nxWhXUP17thbPL2FRUEVx+uS
GBrr2muLSfgJNFG8vZ5EdcBW9OqS4gNupy98QYNZAAngPdRa27VWGsbHjXm9HUrf
/EaYtn6tpecinGOPPhJ2Imv32Yne8BOzNPmLIONJrhZpFu2NaDlMfyDhuxu8DCGz
maHK9grRdsZZzVEPZMiB5CTs5RqUTISR5zQFbShxBK8aThvY70tnzNxy+5ZSeyBU
YY+nnvfsnsOGZ+InrSMy3CN8cYVgo6O39vuWmSpJ08htpC/3r6p05mq3ctBet87L
GDoq/EeyBmKHQNaRyX/sE5KDnnAst/5EkWqo1AVp6ituAUWaLyVzf/o7EJGN6LnG
q2PiL4dbjuw93fwMEgQ/Rqs5EQ8/X8WDS+r67WSrLMUt804Y/w372FdnRZz451FH
uMRrEiopv0UzY+PlXI9HFuZLYc7IgV+wt9Ncumxh9jR16Nk8W56XehiMxsVDq6dK
Mv3qVrCqVNr4qmq/Pb8nfy3XeLNFiseFfhp8evEri4gFPllfSBIWQs0xqPSAk9xG
pZw5p+uDWLmWKch7kUpS1XwSzQi+yoAbcMxTtcZA0ZpUVBSQWsErYORXd/nHrMBr
L0e2Fo2wJXJgOwMb6rZVqUKjtrceQTxefmAdYrHxesHuelQg5IO3khJiKZZ1bcSk
JIjJ4+Ff+hv3adht5eEike7Upe7V1+B+4ZOPdG7W3F39joqeoptegTarDyoW7SqL
AjPFdfNhUnwGlZwzT0FLFWwglnEgNi0F+aOZKMhP5cWI2EtRH2gI/2JNyR+wNybQ
EEU5yL4RCx9/0owjJsc2TcTzMutCNQx5QvRX7xRb1WwSGOTnm+7KTfXcW9ipk4cL
yWSjP+1EXzO7gCZkBioVLDsejv4p0/DVMYt/cBmMTdT1oNiblsXXXKR3Cvl88btG
T5OiTIrFtMD4lA27Ze22EYHx94wJhk8a6XkK61NNVuTlIkFw2o0gA+b3yctMqydV
6xOXr3n+rxZP4h++XqAW8BdrjkK08YJBbk6MSo7vgYivyc6cx2BvssFsf9mawIuc
iYlfTNYLX9dGjW3FpYczVBlaDXO3ahcWIeqlHHTtJqkyW5uhlX4srhZRmsCxWiyS
Trk9Og1Z7QkaFcQBiutQL+RZ+PeR2ZWqsYWoM4RWa2P58Y74/mvpmkXVEaVyPL1F
+bxWIgxuaY/0nrLSSd2aGcpQe4qYtlR0LHwy5a+cKhJKFCbUfX6BRXXrQJ31Han/
8SjKiPGCVdYyp0wHpsk9AfDsBUrjPEH+bZ2huGhZPe3sX0fw/Pjr3j5bPleGBJjj
rqHpjJKgPk6kfIQPCIRs0iBc2OgYyID8OMLnzfajQB+Jzb/iGwuj7J4RQVhmXKkZ
o0dj+ZJOQvf4nkNrxKsUyFbB1JLSYiuN9bCDnaosbkNSJ1ilG4bhavAGqjWE3658
zz2DUCXHGwPrY6XHG4Y06kFEbcjuCEU/1XBFXpOl/04WwMk/RHvrvgelGw//WRfl
SewKxY7h02cBaX2OU7S4t359pUWFgZd14ail44ZH9vhcTRm1W6TMiEWFdC7Z7K1p
zCkDpO9Tvhkt4EAQeNZ7vctqz7sxffyT2nHfr72+ic/HCnE55yL8ZJslTTfrczBW
AqGxs9gwuiHRPU3Irm5U/LXZMvfz6z1Ac06Ut++2bsLM/RArQJ4RPydDvwVJkcUB
dZ249fKZSIzZTy04y2cezW6aTV98Vch51Er/fOVbuuIsPLzrtO1IFwcLyoU//u93
OKQUPlza6CkMcRMxKJibXmo7CXNyaWTSajELKNHqvkl0iS/fqBsmgMWxRR2n9oQ9
P3LUp9lMG1mLe4SEW+D6rr/8tGS7R69YwLwBeetEKBPMWiTvuxRGRXySoYbKKgPS
JXKBzeHrGXJpPLy2lQjuiibaZMBA540HqpXOgJygkj7XbUT2s9gDKoTNrXOd3UVk
9cDCQ/Yk9BQOyVkaDXaqZdjhbbq4uO1B+ZsOq7ntIvNYOPJ59VJYTjnJZZ/Gogt6
YiEYGnT9iCV04ETS9307/16czKK1eLyXSqzOArgwN2ZGM4jur6Eb3ZxnbOIt5V21
HEhRzIIpOslWa01BcX108y7BtA9R9yCZDD9j1E0tu8QZdcJk3chhN/skWDY545wT
OayKflfJPRZUvaPOoDSM/M6PyU7ZSg3n0YUGqUmizSLn42Am92jkWLg9G669VW57
KOs/zzk4+2JByGpS9z34bywbmA8+7YtZ54neBpcNMrdf+m4boz/Wqo0+/hmvzytd
vvULwVKuV5C6Wbs9PLMqXu5QVtO/Kra35fxHGgo8bPcw23EUBB3aYwywK6GBfqiT
m87/KYbI44M+yZSN1FTtHZnBDGO8MqKmTWWuDw6C802qeWCPhOtrngJaokGezXPo
7euYcfgdn45TE6hwy+Sugv6m+On2AkalQ2rn7k33s7hABG29J7DUXvnruRK9+MUr
wBOwiihY6ws9JkN+GXH8PCC8n2tLth4FZcIiLvqmy9rHbxo8DbOg8j9KM4XLwT03
jfiMRpGskKI06EcZjCv9ZeZTHxGfKM/yR3X6sacwc9QFRHzH7S05yewlkbRVMlDz
dJ/x5UVZ182de4z/NwS8F1H48uUP7sVULdIHDH3Wcujjw+bQSzNd9wH9rSZoHByr
/AHT2Q1RTsCUF7EcX2y42DqbKYIE0QxVpX1YpKfUDxElvqQZKX0AYFEnPfs6jvyB
5LHXa4ByT3Lqrcc+e1fC6D6FMPNxNc3SPOoIj9Cw/44SRrDDHM6yWoKLoJ0lul5W
32JAu3ZITz0wpRXgwlP2ep1ZjGCp0YJ4h+pKcrKVpo+uPIaiP5ZQqtscSndOHUGK
UdSX7+gah5ZAv7qaU0VSv4CALGv3557Vbioe/ufp6jx/qO84OJgR/Qefi5I/NYwe
8yJDpy955ufiWyswQLCuc4KnHqErSx+el+mZYAAdSKKgZGbfaerMs9/qGU8waaQR
0LHkfyhvDVXOlsDDcQOTP3697oCMT9WXBBMY1woCCVN83F11GpkZNAloU0BTMP0x
U7i904yqfqClumYZM3wrWigKdVPT2AuwP9S+CKMRax1IhwukPSl4fmazdl+rItmO
s5CVDS/ndujy/vQTxKaH1sAhVHdgmpqK1liGAcN5qjBhiBagEQrzLwELj+o3kxBb
HUrA0V/k8rTPuvDQm5+1YB8bMqqMp8LqqgR9ImhRr7twqBey4k21TrKdcfDyDP0m
wcjLHazsoaN884LA1yqvyk01N9v39Q8AoHvm8Fzq/NojWfSHLxAg5SIEQk9CPPii
V8fBzwLwtBlClJUlnMmvrFIJQx3MmAtjjBwTLi8IFnPqs6yO6LeoroyXFsBbolK/
wx3K1gAfekrpujFhM+Zj7CL+8uXz/FqmL7vJCWWlTudOKWA4DqazAr+pexoZVnbQ
JkXdB5Q9aGtwyed/jPyERevHF+nqWI+u5BnFQMc4jBMKfLoqk8deWJywsStFPVnb
4yqfWRGuBNpwnoDR1fO9v1RwyNPJR7p3mnxLz1VFNqAItzOeU2R45dtveT9wsVeI
tTNqfM+EXuojJf2ixJqvJPtLDqvi2JcCmxh4mZh2hTsfEUSx5xQvZfd1IUiO0wwn
K2BEHi0oMBJucGQrMGCrMflXzSAJg+tPcFgJ5QovwuEJAYTM1ctVAojPq8Pso+O6
wmuJPhcXVfU5IjSZjZVEDXz+cO9Qx+UaxjeqYyrNQvdfXCSQ7FwaT+9c3L57Vq+H
J+hQSkB4yOMuAEACcs5FAVL7TrxBiW+Jz3eTTOdPDUd+wGnS5yzYjAkWiIgq4ka1
227L4HnvxuBV63lcRSRarg4IlaDe1kCavTDiRzC0KsPakf3vwbZuyMSQw18IoPiA
3K4txoPiF9BboTcqQ+oqB+ckIm0jmzDoPMplCysefT1pc37sQn3N/WCLJ+2XtIf1
mppqBzi2j3kmQW+lT5ZeY4a4G8Mi5Ctokul7W3B/aPOsV+ydzsLnO+pFe7ej8WXZ
5PxXThv1M+rAxcZJezI5MpysrUSzIHtekKw9PPwMwPI07yUk2fbH2cDcMHMDPW+T
TusuaYVRjitFgfbHBi136bAo25Bf/z6jVeb9pBFgj7WikOnLqIjgfAtcy0i0K9M+
T/RO1Ox4Xc/IZRUSjbPHcPLeBael5NEx7SyNOr0wbnMvMcPUQUVdQlkHqbTtXSwD
neL9S6/4ZBGVzi4hG1JSeb9k+C27CeuP70Wjf8WYmoBiPoIJOshRlXOZ2aTiekAu
FO8ANEj9QA9obfbsl6CnasmiE3OjvxfCBG7TmCwzXQVyw5s9bcPOU4mxsR7NDQcp
wHgJSQrWu+cMWISgMnUZsNyqiKGL8HhvrcfjXm6TaT2CBCruY3Yr/l7I59udf0+4
hj80vCzg5z4l76FIiZXbUdF1lUD1I/VyJWUioaKfcf5HNxkoYTHTPVANqTmnRSc4
cgKoajWZVBeGKTWYtnuEAUP+9h3oY1O4I4b52vVl1yaylUIK8u1aIkBhmbWTSY4e
cDXbe00I8l7rdBgBYQMwKq9NMXzK2eMJy4ChMKrf9vfbQG2HcYhUKC6x7Tn5BzMh
aWEYbhXk4rEieb07eczfc8JdNwAqt79B7CuF1AWMsMVTgfZITdTniwslZwJ1SQ6z
XGILbtmvH5zOuXWpEpOldNLVrh8SXkkRQZpWEiZrW0P52dCkVJq0P3yoqAfGCHFH
OeM+Z64ZzE5zSNrxEJNeZDfifaowS9D9ZJQMuW+J+4F4O5/ji/6MlmGQkU2sNQxU
+LJCtubNNQgG0ejQn3X+yhfrHHWdu4UFA/6WmJUpRV6zSF2AAc9JQoudqtrl9vpm
QYKLLnOpvFVco05ayfxVGnLqMflfvy6R3FjeT/aSQRlTsxTFKSpIDvxBsMT+WnMe
dNBHsRRfru/lLmWQRLZJ7L59U3+K5UR6cjoHTb5ZPm03Y18WEjl9bbyX1swc3RWh
wI+73BMjOOT3Ueo9UE5vHdrf9PYFAwN0x6p4Jvp2/DyEI586jP0MpRQgEqGF7MO/
ltJBrNAFonl84Wi0nS1RWiTGk6ng0bW4SYsaLTjxtdW5K1r6VAJ2vELSQfayZM92
HYXVkVbfR9v66lAo3SfST+Mdj6Bom/tPGQKgGALZgJ7iGHbvDjcfz6RS9nCR2jWA
bcL0Ig14o5XctuQgZrj7QD2Wt6xEv9+HeL57HmwggejRz9SMSIdNO74khC/XsRU9
JZVWitZqefSWuS+QyLHUzH15dkkJY4yr4ErNR9LFyzkq+dJUs+A0+v/Z1MJhIInU
8m8DpiDOZwBw7Wp4LQpRO2lKpyyJ04YDt1QD0v1PVxuRneu1NQ8UUIs8J2fpdSa0
JN0rrKW5bUwx1qmY7IwgD9U5UdQVczjW/ky8r2U5I7KuNhyKgi2PvNt24wqv3Vqq
4nqb0kf3xjJMHQk+tDpNIqVtGJ4mTd4gvC409lt3uWREAp0tO1VFlObx6Gdqjlzn
Hgje2CvADrDyozVSn+PJ8/YsXujMFhyQ+4Bq7Rhh3hbb72/zNMGq7x3Mpb+gX/nR
0Ns/UoEKb0nEL/+Pp/OYHtsDIvQEh9re9DuZusBVA4prWXOCQM6H99XPZyd7WLyj
hVI4jVM984QTuwqNy74qlUgmFRk6SYYUJcnzWW7o3tX6pTgytavKgindyRXL2BgT
dTa2zFt6xgMXwxjQagOf7hfG0OSdGXXF/dIJLs+zoax7drVQWGVZ8IhnSgPBKQON
0ygJj/weRdKykm5r6ioTbDhVa/9wC3rEjbUv9J/qxfpFBmbI1FxqFzKeBckj7DTZ
+Zg6LXZ3GIKV6GzrYy3xBwXBL/qeSS0AAZHi6WcypZiwvonfIy+IWWrugMMl+FbU
0PvlJ3Q1VGykJbW5Ci2GV9/jAr/lJsumEvAOJUrgQIWpTQlPjRrdtW+wNdtmNCxL
qaL9K+0vp3eG/yDUd1LAASjcqUsvXCdxuwKBMGULazBpd9LgdbZCepyxPsCRu9VB
WUbE2If8zYXWFXLgF4G3BAOPzZYSoXdQQ4flQqoym+flQeaG6DuKCzD02CoQwkDP
Dl8yDZt+YcrRnEoeOIyVD/rH3zKPuwlsZdM2tcyPDbgb3D6e0uX9uo65MJwGL1m5
g4eck/hr8s1jKVrAtC9QL2Msg1MyEV6Ii0l/xeFwK1AZoQEY3rgLvJAppOpdFyzI
w69IhKHncVOOpJFgJgOHZvR46y5iFdpekd7ATDPydhMogpx8dI1+vfzpltl1zhzP
BydXTjG85syC2HpubwQqni2yMSmmqf32uXTw7tTgZaclHjeEZ9iPDooD/7yUXwJs
sxJr4XuKpIiPpPRkwnq2lR0KVMIax5Es9SUHwdOQoY8gpO+GNUiowi5dsCcbvvcJ
c7KH3SCdhJI/J21huwc63Fz8uIFZh7J74lMBLAk3B7fJIUe/gZcM0CjgeSoKureF
s3acesqpzStuLcKew80waaxFT1C5reQj2nl2K3jbsgaK6PQeYg4o+kIDnIjMTRnB
4MHDYLoiRy673cKbCCbhbOR2LLue6u8+Hlse70n6Tz6M+e4Gjp0F097lR80WzCER
syVmIMuOLKJeqciygUwqhmpT/0MRhQ5J7CzpNzVnTfjCg7V+tHAtXUthuQ89JDah
eyllcup3iVY3oIWTz54mf1HCeLFOUU+oTyMU2RqbbzBw6Wt22Biq+Exkzy+oqA+V
2x2v+zuE/vvDUDtWoKeZekDXE9KqhUdWJ9BniEN00LrpEa+voNY8tffj/sQbdAjg
JlrM6bEHU8fDSLBOmXGe8Ev0XTQXR7xtoWvvQv/+Dy2Vdw38xtJVOIBEA4PTWeAp
M2d8DcV4F/UqxIzNS86L9DGYA54MFcnppzAdsb1zfdG48KIXFas7rLsT+xp5j+P5
+Pv8WxOsIZwVbjog6B5QamlKrIFM99YthnqraWKaNgCXMHCqElMhGZe66WH/izwz
zvaXkpaxCamOhbC3X1h2S+doaN4LR26nHTVz2dgWNE5qVelVWFcEdNptfu8QB4P1
l67npHu7sFlk9NFyYBjd7X4tT2WDouvQV/1BjYE0w2FxvadQJQBM1stlhknviz8n
JnB21rUiQFg0SNBp/fl1dOYrIBaDbkN7f01MTkB3WrOZ/HPIEFWAEL1qofGJKahl
F0pmennftpNYNKi4Rd9sy40FDGnq6h0qOfCiOeUJBrPikopz+6336ZzAMAtMwpJN
3oZ667W16zy3rrf3TYOu1l7VODfHnetHzia6Avp0oRFKsqqiFYn9X620QqAMpOL2
VM5KXuEWald5KJVHLAK/fZLokha+ItUL+pztaAxnTIqXXJE0cpyS3Jdign4tmWNF
ZSmn36/Yj40LoxpApGaSB0RkcELMipLWGnQ4B1TeXlUmORXzA29opflydF1OwW72
Lu9vb0fMVlS7g4NWPF+ABkW06NCmd1n0JMIpklqz7+E5i3vDNHTLWK844WhOnfc2
q59K8TRnemwLgiMuq2dKcv5oy8Iv7QdPtUOfDdBvYdZRRrT+go8WFD5qJSie2kfQ
cdK+f/EZB9N0JJRI/ZBDlTq3HfQ4pQIxcTz/hbqraWQodOsApQCUQ956mhqFXfcJ
5mjWULlLgOzvEoLqohg+fNI7U2ORNTP31j40O72yX0Nxi5XJS4jToGqMkDf1QCFZ
zpeRVN4iTNyNClGm1UI9mvQIOch9VMf5N92DIFnbHF9iGCi74V0s2FObKkW3tHcr
DoV78KhxdXZjsithdH0aI8bTh5tzA95atKxknv/F3EwQSJGQwoAhwNuMI+DUacA+
exA7dlM29srdjGqFFy6EGGW40GbUf78x+vR4+NwOGzvusKnvwMglGx64EoWBjHVS
7Dr3+RD1774mVIt4KuGMj9UdVTtpvZenoHcW5cyy5AHw1ygpS6LFrEdW/vj2I6so
ifJZs8EEg9xW+gWNAkQvZqoW27wv5QE4RyeH63MZ0p1YG7BmytSFFcsLUxONeqpB
Z7KdsiSK87JCbtipo9cZHPnbuy0MQfCH0hrLO1ghjB88z9OBb+lX0nbIlwLe3Xav
J9kdvgvEeHLAJd9OSnrngZAgzCMTlnQWHKeFJvvFv6BDmeQyIKIjDe3ApcoVvk/O
1eSugi/AQ80APyoVVCYvZehueYpdcgCfoMfhn6gZyvQIhXIJvc7MdHVw96zU7rkJ
t0JnmeHkxNB/YyHopHCHGYD+bqS75bRpD58yBC7Lw4RwgVlzAlbyzolFlKzWSrTE
+tjgxeeoNIhnWp1zeUH8zMAzZi0J5BoM2kwBEsWVgaqAUp3/nTFgFivWVBRZLi7+
xzgY/Kg1k3h/4BMKvd7mf/QH5KaKkRn6Pv/KjkWNkYIU0lUj1TWsTPXDXQ215kTQ
Fgx/M1QVav7IwOWWKOWiANuc4YMizP4SSgOefV3BJvyhkJPW2CizC3kMEWKiAmRy
yN1kUl8Hvtze1RE7qazJ291mpNNeIj7tBaeD+0qDbSosce8z94ut44em2anKCsJo
Cjqh1kQfZgpUP3lcuVK5nG/TG1f+drKtogKaCnwhk/4FZRv9aM95xwGUeTr/qNpr
BpNS5kU/eiWinSG0zhqae+nq+HvsNnRxALZloe5gPzgN8ysNbLq14MpyFZwURnwV
QeP/JtZ9yCdHZtR6nFA5HMgDx/W5ifcMzWWUnvga5kfuzZOhSYFkKxfN4LvUQXLi
kmDUpeLEd3PZHPFkSFKqUppau0HYoJTRKSHJyrwVRX9pNZb4PLysz9NkuGnE1v3S
Mndh8kqx40mVdjDwrDdCA0fYuIFdgEYlVpEPWqdnIhXdwNwq9K+LayAy4LV+y2k8
mzVQSR9q3aSAwaFf4djlQNASg4/2dwUkolOXuzkMm+AvvkYgS0ZlBiYTMIzAU4bM
3k6VpjiSemUeU3HDY+tevio+xftHY0AM7TtSUK9HgLwwhQpL6wA+1B1o/6BkDjh9
f/Tl1Sz6Hi/bk1meci2XXbUYZceuKEdm+8jxjAPpi36b2DxcL0X0OHH2gR3oNKnJ
WySdiI16mzgBvu3ACiOdTdRxA8fK+XH6zR+tj3KsT8n20VNb5kpA4PUS5hruJlzT
vTdrEtAaTv4cG9PavgYbwMvThWQUBBABc7Kx4FDENP5TRnPMrEeoKFCe32yxX/wJ
5ThniZqsC5OYxfI+2PMCE5ospdxtfcMf5Wl5igmnfYNobxP4eJPPaHFo1Lji9u7l
qLQ7R5uVh5nVVlDQDlnfSGoM5eL9oyAoLDF+PZyqBsglanebcYtLbelIhNOcvL7a
2Lp6Vt4ccFTDeWzr8Msfft7YhGaRpnKbVOORx5QQFtlN2Ng4Vwh0uw+okfHJ9ua0
KgQW4GgNe0t0jhF1MyPitJdHhg/G7jjusSuy3VmfiqSa4pTX8kTocTDzK1TFKpow
3snwjMlzz1iEZqvCVFLtbGXqTIPR/bUco7KoRvLWg5XdcnRhH6jeCmmhIE6YIs9Z
Hbrp2dfJyTg/M5bivQTvk5EvoNtsh0o34Sw0xqDZWZO+Uk79RVZh/tk+HQSHvl1W
cW+olR3PWq1rQ7Wdo1mnlkkUmS/L47wAB01ztzgOGqz93mRvOmnpiN5o0sZlGRrh
oCKsgSLXhoFhDA8YDzCgviZYK44GpsFpCHE7Uqh0HW0HZyeXAcXmfcWQaLJKSJoQ
V4JnuBVbfG9dbj2iiUoVwNeHrHzkRJ4zLkOKhxQQGvSq78oiuEthxTt3N2UYqNln
x6wRAe6lB6vFIWAmkmQmya5+LgmJo6SYsKk3+ETGUhbHY3O22PO7U55hq4P0Wb++
ZWkogLu+LHhd3c4mkyZRoI5cRl++gbvn6Bovvm0s69p1XK7KF5Z9GznNHoz5VTdH
7cU4aT5T0xxeggR8h/OH3hh3wYgwuqsUMWl5lKGo6gVoP3LifgiUuLrBCfdZ/TEz
11YqjXTdvVyrGcFAbAbHAMDI+W2jKBGGm614p4GnPy+ROHJ5YRmpnyESS2/M+482
mAzdT5aCt4VYTKCdOMMCq7XO96kmh6nV5FNDuuAT1BE+6xWR2GSfo0hXqjvhnRV8
rX4nbbAQdekktJVsJCbeE5CnMASoxv0LwcCYJW4F2JSqVVGcpvssZva5CpMr1tt3
iFmrOg2qInq3BvBJ1kFuBpAzRgSxjze97qHMkmhNzF5sv27Z0YgpJYE8vTrhdx2B
Y263lxq3m2Jn+2Ilm1WdRCQhPDlGLnjFL0f0R24bCHK5ZZ+dMJCQfZ933b/tfxFG
ZBDMdPi7cg4htWBiSmkie1jHaxkxlVKEjMPaeeGiqaV+hI8i8gxkPiwtEnobgYxb
2WeNNThYAGTG1YL8de9jfXlkot1DS0hZAv9ADAxnanFRRf7PrqrE1kTMJDtQf8EN
pRBBJN3mEBRBg5aJbehiO/YGOTPDB2y7utVmEfgcPjpolEWLz/8xqAN02deqcz3O
78a2F5CVGeQfpbqvljJb/Ot52j2psvg2Gz9XM0QlEhx8kaUZ/gkFlpHNUBwrU0Z/
Vs267Z3hM76+2hEJfa64RQJ5h1fRpUF5EZK98QSHb8f2C967TRTazUnIx7jtNiT1
qsCeu6+KfV1Czk7amY5IkaGSCR19zanSy+ALL5aP8O9xExKh8gw6vVm16ydlVu21
65MjOf2Lw4iArxqtbBc8+rAL82kgpzHNC993cgjNDozGQQxGEARkAZCv8EdeQWJG
lsnFd+3ePEYosDB2uT0bSzaVROibQ4eUJSX4tZBJCj9XogBYF3eUWUksZGTvVkKy
8mJiXia09smFHTFkvr/hcicRPoT6I/hwAC7jZxQJZXFAcaddc95KXTeYj9ZfSVrJ
xwpl+olwtK62QP6CdfS5P1JM1x8H68tWQ+Ojb7RR371fPz1ItpVA+aTd9yyzlE7n
y/nCkJI8igLDuNJrO5XIinDtDhjcgGtXAhyuk2FIxYaBwEAiIO8kigErEIixIRAA
GPE332cus4x9K/oNjfx2bTtkvrDA9bbkXw7SCgaGm8xOyL8rA44Cu0J+jZhIzJZi
iP2lGiS3XTzOkT4E2ij81vHTeWJDSVNEGR+Ws1hO9g+H8QMq2QIX9EHCET1cgbHe
ckjSEUYXtz/SFSEvbGUIFBCR2p9lIPbHEaN8Z4QPs5rb4+Jc6gc/4SDKFkV9YM0S
f8YszdiTjTB7wzQYjUhoMsN6St+sjnDds267iMuxw9ux8Hpo4iLx/gAoBE5E+vQu
2HYwWR75J9x/Pon0sbSprY8BXb2UnaMEp+II8Y8ou/HI27EywztCn0AxKk+Nk0Ee
sUC5NGP7oPo9Flp677pzlW0+P2OMBjjNWabeU19FFonB83fIeCeHO46HHqUuLF+M
qk+/1GU2eHbzaY5HeWk0tM0R+vtlBw5VhLo4M8rLVpoLywqQLpOiDe7L+AODYQM7
6kYrZIlkXjQnFDuglllQLZAkN+u1WTeyg2sEesk+NcjYa355aRosFFAvBtlp0dMr
E6LzH71EkmJaFM4cai7vovFVkPi5c8ZELdT+x1n+yR2mS82ixbOlztoHMJf6Q9i4
mOBt+TRzHGgkgbv+MTG1b/WIDTQ61tNmQJSeFytX8b6BIx9RmA8FFTUPm359fF1w
SbDaISmYKwNyASY6e+CXMpd6SgsaurD7THJA5LKjAN+q7/PPbSOHyuGLPcRQLfA/
mjHgKxeNbRonc7QIZ+JiUR1KEDsUzdG45/3UKY26oBRh8k4iSOS8L69Y5nQFzDum
thbh6GshdY7Klvqr6TuCkw/m4hPYc2aqgTOCToyEAcPdqTuAJiEJSNDuytCMCjr2
azTVa8Nva/mb07ZF0MzPxHrLsxsJ0LOZ4gI/vBuTUpqbNkFGUy/Ee7RcfFVcQWos
/zyxqO3PoGFh5b6YY8nRjJXSzNmWD7Tn0MJhFzKVUsbpcZdaX7EU5gr7vXduNgqP
q5byxsvL+3kEqxH1C4aKFK0hfNLblhFLXX4Whf7JsRIsLuK/riCxJZiSnG8Ljttz
Dc1IPix1POo0/jkdYmhTSZf2MjrKEFyJcUAFWLM84juxzcuRYJfM61bmqFoKKykh
Ez+ranXMm41/YTgRDBzmb+d5dvK9BWE59er26jsVapRcOf+PYwjPItlkLe5WY7Ey
3/gk1o2LyIOa5eS8Ih6y2OtMS2/1ZLnlgjbpjyKIocDDGUmT/XhZBUq/n+7ugo3O
STfonYZnSjxz6/IeRNxacQ1rsA8q5qDPtqF9sdrzXCeo7ulJEHF4FypZfCSoDFXT
qUXIsYYdmToHT7bMK8DQHmHvJnI46qAm7+kD4992UCNsJeTTboL+WnCJrbA1JCaf
VMPeAPuT46XiwZGEKpn+KmXctENWo7lQdatTzCTcxDuQbQD1mn6wixGcP85h+XUR
qi827dd+YuXB0vI4FHKjC89g+jVnxwKH4dt8bZHy3ZlrJqXjrcrjQ8rd0+LTkHur
DBnlZj/nC1+o91mikA3GHMmJcwuj66Zjwlo0bGGVqV+ZbYgUmEUg+Empr2C+ABvW
koGEsQ/+zO2ZzOvk/LkpdUTwquFjksJ+d7HH4Yzanze4f402aDjfM63tQ/QtYwe8
d39W9vMmFRoeOszffzRbyeU6S11VX8ypzFDX0Wqfmeb+NNRZZGgBSGXW3goljsjX
pzz5eVIKJUfHILepsVHN7ytPVk5w0DwrCBHpP8WdUViSoYLIUFrN+zruMyzmxxE0
CQojF00TwSkYOkmCeEzTSX3xDPT9sJC20bu54IWOeKy4l5Q/yqSiNgZt/nx1CvPY
ZyJCGYRArUGdgXI9JnmyrFIVYCn9wxixiH2ZgUcAiG/pL1ShhJCfZt2BfROTCvR2
FKA2GAFYit85FAUPYDQrCXBotmmYCK6t+qyZyaliuPNRcB3v+HdoY1KHK6yVc0Dz
3dUyuCNX0LM9HhyTLpVsjnS1AcKVwcFBLtFiiP79XJiQ5Z5/eM8KgMLsHrRf1wWK
N76pqmbbXt+uFZ1R03p+/NlCiKJmCYlIRAIp2GBedZqaqbnE+PUZLV5LwrmJkzbd
uDtcDjgIrK5+/pfhHXg3p5Q1L4hclrcRlcCax2wTdvJUPCyEs8As2cJlHYZoVWNY
bw2E7/CUH7zCXgOA36tyEpk8t4wpLqSNEwgU4SR2EV0GKd4ocYcH+oBk+5GGen/d
r8UeHeVNdQuoJ5c5eYtKQMv/6zPxWZXkKNyAjdnAKopb23jXTOiM69uJfjjxKfhF
N41VILixXNWOi5le9NsSxmrBfyWiKT/MhF0hwVKQ3ZdVeDjNiWeJk2PXqUqeAWK9
3i/nzwuY07yw6x1eyyKvpCcYcPRsHZEyPzNdUXJ3gdxzfxC6YALif/G8+TW5ePXc
9UkkSFL1dp2VmNM4Oyjq+qq8X4ZHNGW7e6zLX4COiISIbhxg0sgO79FNbdQFkna5
QQH+AQKrM2bIKIJrlPqGr2zLoqbTad9c6EA80fTIjW/1LqObD1uFDJWk4fLlL0yZ
whKP7xk2M68AmcsMkk+Iu57Th9lpujKozbxLbvkjdvENasEhW25Ml+3YWmzvQ4AY
qdnCGhwnLecoBHx/RyENSTlXxntvx4iN1GcQ4aXoCmSWzzg8ajUGLM5MQUQ9o+J6
+s7u3DfEdAbJ1tM6Ym6Xj9FsScS/o76djRuB5gai7ozigoye1f0YbbttEy/NI1mb
frRif1/luoZatYJMNtEoiCKUKFgLX/POTO/41S1Br035UUGJTpfA5SroPbjZGhlq
1nmgM0Kbeff9KIq80JLbd95vaLbfYddwQTesFwtV/W6kN2eWOB7Ql+yxZMK3IYwN
Qwub1GaOxAdZHkvejsZMNSKjmGs2Gml1sYwL5d1/joUWGsZVkcnCrJ9TglwQ/61Z
j1r7VDklV1w0FnimRxOSTQVwPRNDQSuw1gDy85CwN9SZRxY+9zUC0NyE0b483RXY
eHbZ63s88+SHagxA0weEHrEizbXsn6TddTtBDuQ5zUtJ2cg36vlQm2084jPm2DNd
GR5fxA3meRlmWWBiwBTP3a/j9tU3EbFKRAA0CzHtfAN+4J34PR1k0HdwM71bJ2bi
+0FRbZnsPbVSIdHk7GSTlWqYNgI8j8PBgY3hBIzC3OMcUT9XPKnANPWAFrz3ishk
ev6ulZdWhhiN4AOhi6vejovZOdf3RCtc2NvEzjfvHWuQb4IvVXMiwEDkfL2TePBx
EJ9EifNRU72U1IWxGxueDToFZsG3oETZ3Uz/xwmOwQYTde6VL24ehJJ8tVrnCclC
oFjRfajfuhEJe+CIUl3hhf3Jqs3hn8hirlqy0v6bOD29jNFwGt8idRqD3SLDiYRI
e+HsObZnC2BWeSJph9np/aCxzNLW9AMoMmgttutsCxd7/GyUDC/x26Ih70RjApwD
nD0DCg4EOwpJ+s+b88hgWR+TGrj4zRn++ZcKTTkXw0YCyWpftX59w7aPf4x7Dvci
95YtOnjQjqm5DXBURESX/fiSpm7m5ZeCIRfZoxqnjCMnWztqGl1PVT3DKt3S2j2m
u5pT9BXxvfT+1pokoo/mEr6Zn/t/yPBfl8l9w/M+86pBNILY+Syxu5drKKxE7mnk
qoOiJQcbnNdjq99HKjr4ZNwvbdVD4pgd3dbo9jRp04rqTKZ72FQx3R3LXIewLWb8
EbtochPJWeY3iXxyLyy9lNQEZ3HTuDheDVxbeqkG8rkZytYQv9UG7+wiwMezIApO
yCrLTBnC24Hb18AW9Ni8NwlesjW45MVD7ERxEYLgCfbpBUDrBOfWg7A4epuy29V9
uIqMfl7Qe8S80JsWBbI2ABs16cCLpM9WgsbBEzR50VYNedeO9sQUHpiFZoshcQL0
3ZZtOWGrOYMQxrRiqOQAFn7DVIWLCChnrZi0bv0xfgaE+sJyAugHdq0BLOoEB0tZ
s7XYJ0Hyh6iAOjhN3O5RlUL7hU+LYvcjfUN8x3M0knK4O7Xi1EzODkZd/THaKgzL
zRKjn79t0lEi88Wm73heJoS25tO2GpQBhCIMeQOz5B1wa/vRe/u1TObvhJ4DceL6
9u6EZyJsXTIcXoP9QlleDB7V67MNutGaxrkeMFJEM1Vw/kmOETJhe4D8/b7naGyu
E6oBx2GAnc/RomKJ7WWdWGYfom0yLJkDK2EAneLpJ10EPLpHYWn4JI+jHgIUC4SB
Ikn+p27F8+7spJme9xZVzulz6QXqutJZFs+xRr7uam/jnOzJnVlRgqSmS5Le1S8k
B3KXFloQ53NseHxKjNmWcqIvjlunbaOMZe9cUDXmbp55xfiYCAMEk9WV0YKQW7JQ
2JIwbcUPRZF9O8Tb6VYPnKUaVo2uIIVgwsKAObq8HpXhY+tYY9ME1ugnPE4nAcxB
ZgW0yUl1MskhacESPiqHQ1IjhBWBCx9eK6Qx91eZbLxiVqH6KVXYkr/ussiMadR2
baHWxvsEeObAaGmYvMKJNcMe/5VcHZ0KlyPdpnjuT2r78Ffz+jsbf+rU8uuBqnya
6eeRkeKCVGndSrf7Co/NAV7qVHx2XLm6zqGpYX0BSodyvZYCiJbEnpB07VHoRCZO
yrxx5so60Ykgbo6QPVycpKMwlc43XMC38RymqKg3BjRmPDiS8s1fXqPBI3WR/XeK
bJqYP6AyfyfJ+c7WhR81cdrX/TBgvVOvevUlfpNP4JTjU3NwrcOHpdDzLyAlT5kh
x+VZDb5UknbcyNmr4w3a9x1wZ8KWUYgdBeYYCiKmnvk2mT9mP4gN5hcg9GKdn1+o
Xhm/rLc/zKb8u7WlZDy4K/RwXBNOeRL85g8eLgqZwoD316+kx0/2ruhL3QoXQuQS
BrLmvC0CUzFE26KCKdtbXTgaGzlnftO0GYkd+bngA33bh85DcsjXfYK45ZPSOPe/
wCmbiSVQCsGg5Y96Y+BsSmFoPuIgfoRiXB8F4/P42U5De1IUCaSZ355aCE6REmp5
41P3t2MsgDYBtN3G9YdgoSxC/e2OVMwLng+i8JD6TofC9M+c8Q1sFw3bHpPTBm4J
M6i06nLxJJu1A2VDasqTabuZFQA7KQQ9lBJeU4LIWoQdKDB67iimeVgcgj1Y0Ljv
fDjqeBiX1APFuYEjuEwpXheP2jcBNOlk+4tD4W8F4w4ioO7mUsiKoIT00nosnfSm
nAD1lC20lUHkENsenUOm9QgArW/H+EGwfj4o3Io5GXThd/2+p0jXn5rm4afizPaK
qoMqWZL0zYMqEf7Jx+qqRU5kuxqE7xsbWPYkNU5FH98E16le7QnQnk1wt2Zz6Bt+
VPpWRZ0uQdUZpNcMivGPERks0q9UBY2rn3lkPSOdmJERRUxOiq69M4CHPRXa8vU3
LLkbxH30DQMAPqxc0ut7tr7OGamE7qEi3BUW0yhz5Ju8+Vzgrn6cNKo0HQNVMFX/
yeVFE4+Q14YgFYTXF8owiPn5Lx6V3l2UxKdRXQ2rvVPLI/qRycAdhnTxStF642pK
PXj7ZBuul+RHr4ZUT1nW/4O/A5QdRh+zyq+B+h0jwTp7o2daJhc0T0OQFDfqMrSi
DZtlBozS6Mhd0prKelnEM53oUr0ODPhCRxmkzV+Ex/txcxZ/dVboxqB+vrteYoLJ
gBZGeS2UsPDoHdW+/jlVo8RhRVre18heV1+x9c8KQt7i3RoYR/Ajh9jGvJ0Zrw5D
FfM006TVCWF0txhB2zcdZ2sBurg4eNB0eB8HMzZ8EOzaOYXPQjfSb/6QQxL+D/fK
dUPv/pZ11zma0PNjFt8WJ7dWxJ5n+5mkoyZs1cu/zVk/68mmU+vlB2DltW7PgjR6
moPapjcTqTOD78YdNWRKXOd2oDhPX6AjA+Zh3xq8WmSabj6EceKUYqSAUREi61Du
XubN+EDZC6vXYgHMOinSyrnmQBO5oR+SoxBY2LVISk020sbqFpoUZu1wdnLHmlGZ
ysE8DxdVhN07erdRPSjCFPuO5uE/sP71Tpif+p4JWVKwtxGkrF7DGQJval7Jhx3e
fIj9D993mTYF1nh2aAuptPJNQgFxyNNe8VvOqzsc7lGvnb5VvcplMnJ7T3vUrPlf
YMSAfjdMOQSgCe8VYgKEzn55OIOz+uAau6DgSQF5lIP1/tHN7SgQ+0mIW93MUOHX
iQ6mccLcRfrk9WNenC3/zvagF2RKLmeOJQavpTVuQJn3pB/xdPKgFD0TBXQCI1rT
KBLeTpMFdurJNR2i5mHOhaM//8Dek/tqptpxoSEcBljvlZ3dZ/1D1CriYrjsLqo3
0nAoAQ4tex6A8ucQT56TLqD9svLt9Dgy3+tCclhsYnDhxMOySGEx4LrpD4efoymT
Koi2F39+1bNY85CUK8bhDK425MbLfmVTVVhk9pr6YtHH9dXEx26AM/6Gyn/qyFGC
oWK9kt6RxzQTa5SUb9VwQ6DbB+igCUjYbGhZ2vM+30EWoW15KJ/rxKJQQs08TqHO
MmGalBS4m/tjgtQ7PFHxwcGjV5P5EKHy+0UnbS00jpzAqYx+n6sa1LC+xQs+ZIjM
dPW8nu2sumXENayXHYg2PAsCgX6XjFm8IdVEfgLBkmFFJKplwp8L8mmSXSqV5bWP
rqmzmBAUs7+mzaC75aKs+HVS19hCtzsk9Z6xC9CXhrArYVv1IM04SYHsqYNqFCWO
EmBG1jxdq2rz3NyJXXqXlH00Ho+oRwmh9qE44y001i64ndqsus9rJYgUnCtT0nSg
xRa5Lj1B+pa/PewQmUqvzCs1gxNxTToR+rZzqErhjrlP41vRXElrs2M8CLMHRapo
wJnhF8rGV8kt8zNoSSF8bZU+I+1ZVb+CdjmEiWfyvb/USd9z8tOj8AXRy4KwAVnL
mKBx0aLeDZy2iLlGmIV8/tTWD7bcsphYdAaezNC87zHnIJUykmk78levBsYMIM/Y
4Y32Eib/ewUUYHCGA/XHKnhFKpJqR6iEs+kMZzKcph8z8EL35XTYj1BjE5QZW7Lm
fBpLf07dHAQYvEANSe/k5Ohi7dcBebokIC1+gsJ6zZhhbpMJPkygNPPVjYHMMapr
dKFydd73kHoz4WF74eWDDkr7k71tVeAczGF1hegj0BWjEUTxvvjewr8kThyYGqI7
JLGhdYQ+bJ5zAQWOUsA/ZZIjXdWfwvvuwH9Pj/m91WBRKcjCPoSTo32RJaugWFXb
11RKSTsnzpyfZOljQJqxCZ6KBQ5D4/ae30UOp5N6h1C7CVb63TjXXmJKyZBu+8mK
VzpdPAu6VdJprKhxqBo0KorrJS+vFWBUdJja+XvSBy+OguS7r1UgXuG77zS2qQFX
AnUot7p+JCvqhSzHWMdcpJed3lzuL5k7gYcvLxLVUmZNtEnCh5u2NQ8Uc0y48hdB
CcL/FjErHTxPTxTHzqYGhbUTWAwq0imc4pTZFz7ULGqlDppyXYAZo2qidCfZYfEu
psRmUOyVhfaaP08a6U6vxfPptkuGLCyxo/E3nLhDuBd9nJntvsAqB9sz2uR3Ow2W
WMCYlze0bcmxtiaAme71MlkM6LWel2Twt4ksDvLwGkpMkxKXMHxKnsvGWfCMrvF7
Lh1n1b83lm8VR7QdcsaMJ4OwP18krm5ZLwQDrvzkcvk12s99q3BdxKId0F6xUEzY
Z8aN4wC17FYuGYV1GMyzdes+9takEGIfCaupbc3NYY/RhWnqUxv956Tf46sNsPVQ
tI1cLumBmctKqiOuKlfspqrqf1GBqa2Wji2lkSj4jOwqQtBZsfN6cRqyHLsmH7Gg
sCm6HwBFYgNgFBhVCS2miJMH30tjQYBABjpIubpTmAIVC6ZWnDNmhUhPvzl1OAFr
03SF8Lx7btPwmPZqenZ41j1ztV5rAp0yRpCCyAHMlOBWWyZanGY/Yy4HSgSOlARR
aolfp1gd0sQoEP+af/XNtgJaJmEGw+CeDSbKxKGSTTPwTCym12Pja9Ai0Ww784/Q
+tFoia5cucTCZsjZB4YYr9XE+/fVgfAlmJmajNO9rAPMttp3Dy7vxZlgnktpNx25
EudpesXMcwOpchzSL0WzpKefzsc8ejUclauPDbcRg40YEXjBT6vTW0EXrn72ReAe
sjttqZPXzrognaYs/x7GXuv+GERP+2CAM18fMNH4g3/K1rnLFhPNaF5WL+W541PD
DFESar1Gtuan+cOFuuwTNlrXmBk75YztO6k1R8gtrlloYNOd8EVR6185trC5hQeH
7jKB4j1gnEfJ2JTKXo981ZjbnV4b++qcHuactP4Lq8CPmbaP+bPnBVqsK8mmYhJ1
hqBl17ONZDkPdIH5dXoEVuyRW0mFW9Ti28CUsT5M19V8poXjyqAq2R9SePW1awbg
6lejtarGuX4CxIDnQE8TvWhjPadWOMKE+CIhqSERtl+WjlarOo5Cf/fMoFWFBtri
5QSrexWlp1n8g3rlUe+bYePba2mv5qKP/M8VrqoSfTqDhB7b9dbC7B0kGKPVjWv8
LOxov+nwBeVcxBlYdlzLE7JNeIqwPaDAyE9Ae5bq7HDoX2dQql+a8pGs/nVG1qa1
uMtCk3XElzZyY7HK+mycvqy1GvIycIuXL4L+cZL0qCkWUGT8juja+GdkBwEazCRw
UP3uSq1qg8yUWLnQWDIiehZPDo2NnV+4g/KUsSy+KeubuuC47VBuqcvTrObJ406m
H4qQT2Pu6DsF801dwdmsb36fWJJPTUiY5Udc5xDWrSoDI7m58NSWbhCEGD1MK7yZ
CUD89qTebQDwbRhy3Ekf/ema2h2iMO98aVCwnMosBo8aCmdWhmljcOheSI7X99W3
xQa321R2ced9NzIfunh4rwP9fLzjFpjcep4CGUKDVshxMPFdXQTy9F6kHXZNJeGn
v6+GU0mSgm3OytyoWk+d54we14tFzFnb+PzrDFRAHgtPAs4UPJNDf7p/BwJgxRQ5
OXtSuVppLYW1i1AtvFL1NcauWf0xNVBUs1nZG0OfkJlpmylJYF1tFiP5H8Taagf2
UiUQMNgFht8rXZt/XcbSzJCluRlM1mjUVKPOlcZhbZMSOjy62ni8/wonEBcvd3ST
Mi9WZTOFlPHRM2k9hwngCTp+oVpTgW1o3ksIz354u+Qh+pbi7X3zljeC587QkymQ
h7JAs3N2UVL1fj7GJpWdNOVI62nZ7ABGElLNtkJ1hBtGtr/0LdiX57va+oNFt9HT
TWcF70W6iewPWGiqxdrj/0K1NdZlqG5we9k1Iuj4YICd5/ReEsmeEn4HRVvXh+Xv
fElQNkG7thql1axB6wFACs5IyQOOlULUEklzbDqn4+N4q036lQnzzJk+FprFbh+K
8s0BOAJkTQnerOPM9de/29BZZx7t0NbImOGLGTbffE2kcZbRjL72JDHNytDkTi0H
3sJSYIhpM/qxXxCOwmNGhCM7zw+2IzEba/+caupLrRNodwlpEF/4RiPP87dn/I4E
qHSYmNct/d8IW002+n7KprTc45/KLHuyHTzLSGHTbexL0OJB9AoANpQsP2/VGWB5
7C372dmVjy9pbVFdre3G0GOfe/mdUrnQGCuRcJ3vgx7sSB2clObziC1C9OtDjDVn
vAmfKakjYMYdGplGxH2X1g+QGiz2QK57fkYuP4AMfEk5svIDdd7RvZYGROVleiuJ
KtovaomXpV9vlrLilJW0v86msh2a9uWRq6zfj3h2p3TE8ZnZtgcI+fturoUYR4NW
MZM6QwikifEj+WfqTtl7k7WWIAfEOrH0PmXfo5JYExbdxYv44Z4zfqJltWacgiWh
xzARVNeRF00TLNflxe59xN5R2RK/tUfwuRFj2zGMyybgG3r34glwNZWVx5pNIL1i
iokBotycPlLSeUO2TT6ReKYmnkItbFmqq5a3lFEiuOBB9Ax10AS2/eZCN+dL4HYa
h0glqcrm2F/t8suVINiiX0BuM0YoOaL5xZg7KQh6vkOJcNX728x8WHWbIvnvfwQ9
8RJW+mz+9M+HPg1KeAwhJ8u21527SfaqiLbAH4yB9KGbhQApw0hW9i1oB6/SFVks
1U3aP78PfU9OfLST83s1JYCLqISprEHMnO+p83oTrbrcATZCMsL3SDtjq7M7RcNj
+E/n0qtMwG9lREyp3fd8nny87j/uz+hMCo9jlAwdrAt88sTFWulIwfM9zpuW7yqN
mdJ1ltds3D1/tPX8ZHRlHiOH0Ym1FQMc2ULruvWEme8hjNzN632pwqiPoisgskse
iBOzjzvjcu4EROG53vfcsKwOweB/7uo5QiOhrTF0JAh5GkI9KWS1d5q7XBb6lWL4
7lAdhsFisqtFCQNznxqCiAeynbczG/3CB/u7cc5wVary2NH6k0alatMzzL6uSWkl
j3xUDzv2hl1c63p82Aw/s/bw/gYJRkZzoNwBw+ULFlNTM78qkMDCFO38Xnw+01Ly
CulBjUVVckLSk43akZfqehDaddY8de0KIWiInBve0s2/5rvG6SVGUZQd8RSqcTM8
vPY0C5BfAptDZSacbwcKnhFUM9p60mc6FsKLn3LhIJCV9likJVwKUJaEOVF//ZYc
8epugIYGMM5EzumWp9GDf9bEQ4XiGOS6lHpMj9OO8qeSIc2mLLYEpqT7ia8QuJ3Y
yFJhd6PES+7Vyb5L/lIoY2dKJYltRvH+FDVWZrVkGFBoLQ4aCqmTal7ejWsrdDMi
MAWkNJBAwDMObLRcd+TxvSPyQhCq6X1D+inRE3JAguLIxy6KjKrU7G9wGreyVruR
88jaDnDM6vrYJnDQ0giu0kIGZRZQbDuvSwU739KxHi0zJHlYvj8D+LvNkR91dbl4
VHUqDYIe2SEHQLr81lChDUUvk3Hullur4xV3HjNo5E318s5Rx7Mp+CfDs+uaRiER
Rns7VY4ChUCTAC3+0RiUqsNzl/1VbG52MSeVnqjKkzgEQCNY/nb2FokEqk6udi/V
esskMxU2MjTjg9XX6V6w4Et0acki10QgtbB6VEX+7avLE73+sgvPMY/tZrXb/pO4
l+GBtTSwn05LamStg6bhgnIyAGs523NL2obFMxNJv3bGfia/otLdnruYubV+elLQ
v/pda2Gp0TeE/FxL9lLUoyghwcCLwn+lkW0BjshGlb/4CJ5DgnGawmNuELCCbaU6
ouTYDVb4dsd0/UxnBR1KkSdnimBtuI2xovPMSRM5ClWfRgvuceg2LceCMEztHz97
kP/CrUZngETKXnJw7PtQjpUKgUCSu9/F9F22ov/pjQytd17D/nFqYp16sAL9u+X0
tToRL8I9wa2tWk0eoAU9n++AX5AmcHJorydnvY7yp3FjyMLWxLx8vj8qluN0QQRn
Nw3AeKF9+VD9lGtRAUZcQy6ZvyzlxGd4cOGpnKmJUjjzozujiRFS85n1rsBqPMFn
gLcBmGoJayEeQNcyYuE6yD5sP1KqaMCXnIT8wIo1yZyKvmNRaUEoVgRvSPNsxR4I
my1l8Y61OrFb1J6umEH/Gjl/C7VISUydn0FEwbg9dWTs3HegWEEXaw/ZJ4DN6YpI
fTploA+Vk/FBt/CCB6sT+F1ymCxik+EjQ3hhzNJDFp2Gs51NzhRy7Z/qQJld5Skz
zdSzWUImX+Pd57cDT9g6xPGrhUsVm1d6DBSpOkP88fTM/BxLPz7ZptHXe0qQNLHc
9T5ZQGhcW/+95b7BeTMcJUB+OmVKyt3SADzLpLL9UVZTgYOBMOMlWHR/4pEpXnl5
eiLqnkdGI7vz3M2F/NQdqQdzoSNVsbgMZg2EW89Gc7LCnE8oHz/l5xhfy77ZyaH5
0JgqjvYP/9EaXaP9VLzHITSRfr4i65QQzowhvDvnln+cRC9HavIO0eqnYpMS/7iv
TBcLC5WQqJ0hP6H97n4jsOFAC/YEAHxVktMSLuBU9deMWQfyK6BFLhnL/j7ETqet
Lw+UDZJVrdLhXs4XI2bNIqQuUhYBmGYhO9d52d9VvmVg4THZhcb/LwtAheHw0Sxp
TizbyGcXFOcLAROFXdaSDMDHXMzgvDctfVn97C1sCus01mdSTbL/ecYBfsftv6Jk
/Mh4R7E1la2dssGTMU3pA/B/Tqw3/ECiYwwxdPpXALUf+xstDiodkO4s0f1a8Ivx
OW3OtwFz4SbkaOj84XEKtSGiMQvZLTps8Na4b7A/tv9rtpn8Myl4aUHTFeLlaugR
HFRAgQM2IyCPUBi67cKkSUbja1Yf3G08hjHPnOrvdbZetqptRvjmVLpbUUDV2me4
vLtye9IbkEcBmBHFByXFVbB/593XQsIksWsj4vfF537RrtxTEUgnfRnJ6IotOsl6
C4GsdIiq+96b6USwLaBHZ5TKjm+mHmEq/Vaet8SHfCxq1f588tC1MGfvQv+1iWfa
DtqBP3Vjkd9CXiFRFrrQXQUM6iqH6Iq1ztDXMTAAbExeX4KjEIM/ubfoJtNiGY31
RI6vVJryCe0CTiP1ApuO9BmirwNkG9yWqwwtIY9OZxQNbH85ZicD0cNdFA55yqgY
Byutooo+tmGV5EppEAF0egASMkqe2C1LRxAt8a1u/JUGY/n0qzn08qt3Z56a39XV
Ye/DNc9ypl9G8CSvVAaFaNGm5rlzqF3QvpLvXUV40x4r6LT40Jh+2P9Hq9F9m8wy
a6GdKE3AN7i1uMuDFY+h4C/BKUiQvGBbgyrFG5/xrxdfkMIfSPuaxm1VdKKJ5tX7
apLGQF10EzStBz+ITfuQ2fcsJAVt7dSbBKzC/5trIwFVlEgE9YgEHod/RW9o10vf
0p/qZkuDS1gY9bib03AdMbGEijGNqWmGGzMDXfOnx3in1Y1rQobNqj+K7ws7+7Z3
4cG1bSd6aLEGRIOOvlgFH557V0vDvo+wX7AR3RTfdtjxwFTfgXAorGRYitfeGhQz
FyLCwkQhZpcrrmjl3KEJf+9ij9yWZvE2aG/DKa0JeFLKLj5mE+Sqo/NX44XZJPpt
6dggzaYoBvglWevJNKZEURHKQCXdLlCJTIfBNoEtjsx4sty0OXs1owWyZwfSzgpl
tR4/GBrc5c7jXLVQKaNl+EY1BcPtB7DeLlwFtE45rGRCKR8Svz4gQ1wofckY6ilQ
3iXql0hW4TYn/v8Z+qN7krByPQOEmpgZJDnyMoDPuRMzwc2pFOUAxu0jQ03dDo6h
HE3pjQmM3dIybAaTi1yMJRsjdboL0AweFsIoIUPu1r4ZBwYQrD9v4yFSJUbICOFu
IQBfaJK65K76t9HnW/WKOQQrb5WTrDVudZPSGZgkoLYl/NQ6mtiuBPbHG2bxq0dV
RSGtLP8hxjQ52hWuqA65acH4Dxa4FiWl8dRW+1i9xLn4094I87NzB7Ljvs1YOsNw
zz8dbGi1cUtCvYjYeZkITmrl3lRecz0SpNO9mkEyodbYYD2ts+cTyCAbHFoSgbTp
e9gjDaBRf8KFA9DP7ewglDaGVj9JDwY5SLcUrGgpOwaK6WYGvksHD6smL1SUSqSm
Gub0aaWN4bj4WfSzT7wlGU6lDXEE6IeHRRitYvrIQCq5tp7JNE2/T8xfLEBs/h4U
1irVezp7QujJtXXoXGA06QZOmrglBuUn5fJpVWFADFmlRM55QZV/cPaPBGZ4BQ2e
Beh3Rd9GHsQA41/m2h99RVj+vk4Q8SmGmRwZBvffLQTDAlr47SiRA/ljaZGPV/HH
Pq5TG6O57v9SFtQcF9xiQva1cvp0EEtCBlejQ3l1YCrMDHIs9cBXUrXHFaVvTYlT
YlqFqbv2T9WV5d1ObGVIJAG9V6VjL5hvVsjhBkSwAyyPEJfBB+n1tyyKMB1orUaW
d7PKTeWyjMbDJ5vIp7rF6hy2K8vlCJSF6EAcy9A3Zwp6mPrfnSPgaPXXNt5tx5mY
r8PCWSvCdMXc2CN0kRIIYVh8CCyGBw2OUD7stWXUdUN7OKrKhM8J+9tTDuYHV8jw
NSxCbxhh/5j7O6T08KYPHl4Yz4Te5RASb1ZpKCBhTU7G/rhiTVWHaYhK1gCSUGTG
Fq9UqmGwh+78/bgjkY5r/bC2Th1NjtDMRkz4OeUnvrc8beh3xOEiztpFg9feQNvT
tHOmfKiiJTBe0cXywfcFH5gM5J5UnbM7wjqkRdnik2fgmGr5GXn7YP3U2e7Ribjl
389VVlI6qRVsOy2MHOegCyZQMOFqHaeJTwtrZ+RPupF1IG67xngupxFJ3sF1yrml
Hyy7+hyIeUiAdfwxEoNlv/bMEnc+ZSFS5M8gurq4fqw3PBjOKxKUyfs+BRSdReCl
HLIsFrRwc5DDomMha+HPq8jQkfcN0NiqAVFrWtaed2R6No7N3bH/jd20YFDA1OrD
kHNEAiGwmn7h048mCDcaJzCMRh6qOE1JycvO2/7cgidJsF6SaW9UARnNGGngRAoa
HL7dAXz7Gk18pov1pRpRDBLeopQnHDGsg1k1pFwY6cYq0OsLxR16kSHEexDR5T6D
QjuaxY5e8hK3xT3XsY6e3qH/vkJm8e0vQglp71+xPMSz/N3USrqqm68/FAkTT+og
YYCxDWoZc3anW3++H8sq031HknGxW9Q5fxXKC70CesEgzTMEoHuGOAmPhUlImDHc
zwAFLMwrVInSleUO/iQcPMzPQ40qmWcagi4zAohpb09uaZwwPRUDE6DJD67ccZAM
AuSH0NCkdt+xIaqwAoeQaV8Md9LzTnu/zw/ACQSEKnR8GedquQzpDshO9t9JKVlS
pFo9JoPoBqe7/0iHBl9wSZ8Gm42Br+ln446mXqGFkW1RBdS0HH4dHVzBzFISZA5c
VTKCX/fKQ23rsTz7nheWtFDqh/6ihe3oNY+yaHOLCllIHrRddXAbkuTyrVxCu0Bc
ZIVDguHnav7fKVXFvaYyVUdp4OSrP3rKAdZVrXFYykRGIq8jHOX0jUcdRK6ub5ZG
JvgGIupJke2UFWRYHywVG/HenarIxmrG5WrW9WQuAENRo5RVxhb5pySyOz/C+f93
fxQYJaq0FKKYJOITfeKDaPZ6aiCLv+dthYOgRY8vpw+b/ahAPj6vWJtUMdTxcbOl
INe7Vog7eUfpcePmWKdUv3dSk2PXEySk8zwTMEFM6IWkGKEFYn0BuH0WDMEhllKS
Hrrau8Wqp/DkgYlNm0l2XHBf32sjo+h+Qaa/j4FFcCKe3ohl+U60OFahdPUEgMeF
rf02R6LQlEQWK4WFrqzfVxupcrDN+QsewuZkRyPEZ44freKH7PyfyktpkatvmcYB
CGGzenm9sLWaTZKfGw8asuaCnUaGssLuM4mvxxm1Pa1DUN6skSjFheMpQNjV9ZpM
gH7nfUDVYAdKzFsXpTnmyb6y+uEV11e5OTtbZfMGD/P+OeerohGIQrKWayM5Itle
3rfI+I8HA5riFVtCK2avUWVncY0sarmW4jwh9QtqujbcxOkwDnuXM8C2yxUvetgs
2Zk7MxEIHS55UGKGbqMYndbCAy9tnz1TXowd/bxwgm8pwjpskGcjIdRtB26HYSaF
EZA80opYwHv74pWhxYrH1/Taay/ZiGXCgnPBh8yWv+mQX0QW9PpEehI0mRn0RbSZ
3BImaFB7nX6IqF8kK9vrfXQijEOMPOo79PzEc8PkJs6ZkQNCx4IgCnr7BS0rNRCK
iWHtIOWE73mSV1UtXfaT+wFiDBf0YGclI9WSTeJChODmk69HMBhx5oswy6nMAqnL
CSk+9Weq8K+jy72zV82uAKVXBHmz4Agkzt8MOqeLe2j7RFrPKpoY51yLPh0A2SfS
dt+iog96ibaO+wmd7d0FR0UHV+MMAXV7TPXFBhovN7qdSGhhXl+EpVoOElNQbLyZ
f/6Ev9AsambSkwlTe8Cf2MPXywYyMyr/zMyVtcNBBRKt80LO7fneOgHq7JV8S/FK
tBaSlMzPuiQuFtW6RtecUtyIV0I7XjTNmfeiZ5dW+XPBEulDPngCa7GQcKduje6G
vXf7dWHB1wazMyrfUZskgXVUH1Lhj/dCidLV6gdDLEORdJAGESbabbrw4Jt1FXey
HS9BG2drNJPYrjoHYqCQ6d4LKCOKiQI32psZp2rQEGaeD15QAfoDG4EP4ZLSRbf5
AyHsYPXey0xAiUbnKgzlnNwQmRV8skTH/kcKGHy7P+YlmXULWFaJ6ATTlYlUqs3S
T9nXklSXpqO3TIx1g9AR09RKJjqEZgXTldLm0WO3S7B4bEVCO+293sm1v4XLXEsp
ZP0oB3wRKjPaKB/hJ7MQU+dFJhyuc8WIkrcBlq9m9QEUgFiFs++F258n3FFmU9TG
Qi/jqUqeNth7hq01GFvtRX/QSno3IXyodA9AzNiWfYOS371miReFJXBV6k+qGQnO
SHBxJNqLQQMfJ/tGVydhHnLhjp63nIlrJthQtkRi3/ebP0XJFhpV6ujx1nJPkODq
5/wCxDWR4OuWcQ9muT+4N7YJPJhp5R59b9Eo2Exd/tovVWpmUzySFSa5EePVGTHh
NULOt1uZ/kPKc41bMu0VKnufAitC0ZvkXgNpgga9WQTE1nwHb/tRAUyZTaomDU2Z
7XzWxLXBPmdJPJH0+RZCN7Z8WVYCAlT6YS8HNMiA+OFvpDv1EWPs2sTdFSgP6Cs+
tECn5XR4kiks9zdU8uSXxl99nDsPfshdKELlHdXDrEOA8TjBwac/KPTJR+mo/fWq
nBI0vlZyugz4CR07IVKVVUh5ql6oKS+BLVCjSt4DDdTJDI7CN+OE34VWXSgD90KO
F1+iEoTUZ2RQEEgs5uSvP32TaUiuU6KQJ9Gl+WKn8UFURMXoFoWMrti0J+1TB5r5
4C+LUet4+mfZoaNNlVy8UIC3KNfCTMp27nkqRNTMh6Em1B/U5NKK1rEIpqMmf9j9
7qzLNwFTpRt9u8Z1k9tc45+JcF1WKv5KxcErALAyX9eKuv29QqJvbII5k/3NzjKA
p8aUpb/imng/IH/Nf1/x5SNktPpQzRfWCsCpl0NRL5zBuKGhwX3LwgAHz3fUWeWB
OzHjMeZCirR08/8Ckbq1mG3Zdh8E8r5I+dH3dkssnBhMGMEilZIOXHmEsR1Ps75N
KQ+tXLE88KUOGEgyYlT7pYv1KaZsLq30OCH04ljb8bX7pOd2HbXM25AwUfRMbaU0
+gHIOoW4fJCMCmu2l71JcOxolkHgNguiipXjYl9fa3ZuDtVKn0VFtJJ2bnEWhstv
IorJqxkBqEWlBheGBuCEwrSPgliBaAgavvfAJ9OSW3rSQhRc+lNIQaMjofysxX8g
bmIA6oiPr0Md8uRN0f51645edJqaXxRpih0NUPTNR09buFKZBAQfwzG3JCZMfWV8
ryxZ/udtDuMErvNNeWv9re0lb6+ZkWLxzE3wF3aDrl+/MuJHTRyXuri4p1x0/LNK
bdrg0Z2WyzYa/ch6UHl4MfL9Gr2HOjIQXZ4B/EOm8ln938hjdG97g3RAo202xfYR
MZWOJkqbg07LypHlzYrl8bIlX7TR2DdWpV+gRyIb26KWPXOE57brdyp4gdBT+mMC
cnodEmv5vAYYk5xNlic7Q3Ea/2aGW/CppHIfGvOTIOcuyWb3E7IKBaSmwyQJif7c
Ymyh0yzqJkFEJQj0OJ0/Em0YliGXEAz5uwY5Z4jPHtIth93Vofebs6DiTFdAec5x
0wjCtY/DfONq0bSFUQ4GNeqIGP2t64069iATqXntUjEgLMyfibDtbMSfr799hSZH
H6Bi6P5wI16zLVJyrYm1HLwVGTXXyRb/alSgc8mxtTyF/vZTUjY8W8G9LXinM4Cd
h8hm9B/gbOHXd2U4aSKBD1myPMi5b2KEYsQCM7K+UJshwNDWoVEtNSGBl6N2Gp13
6XrR70LmtS3r5c/d8lrH6Jao8c/0aoUNghU3FI9F9g+/tf0okRXoBWff8Tty2Cn+
VI2wscjcIr3ryRlaBJyLhdk8MUrl8QK56FneYU+rrosQeDqi35AXhW/I9L4QEigR
DNLPdtOvpOOKShOp2ezUS9SE+3iduL5EE9+1HDbQQD06e7/OFTyD34GuHfHA7dJq
l3PKprE5VS64q/yz55U5+pGcYYd7iW4uTSB1VCItGOkJKJ6hy722OMit331tnYrB
GLovpIdKHR3v2+xr2GoiEiw4yU99X1jhx89z7n+3zbOaPBgKO9quERibZWBN9udS
EAdHUh1fRmcvracFmCGN/tLzOQjZCCPp2RHjSgBmks0HDMH0q/lEBPQvLbAyiA/o
V+H9xvnhEdbG5qJFJ15SeOqOdxJs8V4hy07YLHJ/ZcSwFQUM49zCEtAKbbawf0P1
0pTpAC4KG0zpslvFZMdz25S78TOqqQJLSNfrdomqjL7xy2/mmR1r5+ZHrNl8bKOi
twlLlm+XndEiDUGE/grEu/Bz9RJoeYGGYoWS6ngah20+2MwDledrVQNxIGhBfEJd
DMW1NcNOulOlkjpIjbgrtXo5nmttPjatX7yyNCxmYR9ao/n5kY+6THdKVoMJbDMb
iNjLc+JKXrhvTQchk5Q62qSuemJZHUySz44twZdKrdyjslU60kdFA+5M0qqm3btu
9FAgJzzHwM5lKgi49eS+Yh+gsehzfg5cXI7hfkI45QDT0rFmme1a2okx9e7/nHYV
gN5DWvmPPDSG67LiIBKYVx8DK4mjOp+9XwqJuSJRjvso2q8upsKwVAML9brMPHRW
keJMVdK/JdPLgJ/ujum3L9Qss/ixeAtv8sIb5piVtYdt2cSd6IHzulYK8csAqlaJ
mG1GkpwjM7Tx+Go0pG4ZkbWRq+GLiQ3a0yxgW031x4rHWHEtLEOBlKbzlQK/Z5X3
lFiSXJt1HW+MnNuCIu99Jq9Hwu1Qr2eOgjafoI8nCpultBMl1IQ01lj34BteaaPK
vpyA771nWKUaTIkXEPzgK9rf+7dvo4cwd6m9ic5xoKjsQORqjTZPlL18e53pWxXx
3Zi/6tsaTm8In7b9oDIBv8sm0gb8baDsiRtpMVA/Gp3lYBgVxQPCQKSCJk0jsfgM
wtxkPheUL5z5n+lGFlG9U1080aTqfnYbneEQEmUE3HvRjINOK2GPUop1kTXoGgME
dAV72MALPFGL3i118jNNQM+lviF8y2qgeet/4yP+tQ/2NzuQEfxlVLhZwpYayKIN
uN7fr057g5huz82ahNvmHTrGWB5ClS41pi/Z0cfdGdbh0p9Up3izfXHzSTmUH5Wy
4nemBwDbi/5hLP+viL30eAIPdUAZhKNTSiHMa7vu1eXWQz670CP2ZCKGeNAJluBR
3AcQHqqvU35TQPXieq6eOXjA8OheOtHTrPBIYzOYmVgYv0JMK0c1+e3O2b92D7W8
n89wKXaYe5dTvk2cWJkG6h8Le+82fUlPRfbxRWMaAj9pxrKfwLakGVFDrlyKAPwy
H3voAiIzkOc8pkGLF5xzilwg8tbsm2II/oX7AH6qYANkx6iCAKsGNSUDvHngBLYP
4XC56MvklnRp89zWq8ssmM5o4eOa6c20I9xj5pvPX9+yPQKL/zciDqs7ejh0eOuQ
J0C2b2DCzGz8JFOWK0NEUEG0vPN40ap1wjXP++GqzDXKWquvSXiH7OKvhyFEijpU
uQZpXjhpGb4a64nxjBPvgiPsYZcw8rarc0Ddc8TnLS6wxvVh2TpgvB2MjOR+xiVl
u/O71QprTX1Zf1QZ6oNexQ5f3zBJ1jwiCAKmDRjGmXS76pX9byfp8WTgiPfoOtlf
sEfH13GtCBeMgZK+IyVPfscoe2AJnqjbSfaGkNf18xb0uf+WxChrFpg7cT17t3lK
FDXYF4zERW0WwVz7crfAoT0Y3dEsVa6AEMU3LZsZvjeSazAslBG7CEe5WmUaUgHw
T8gkGjaGC8PK6UMlctJNUAJHoeUUesrkRIYyuiNEXeV3emdIz4EmpgvuSwDIuzGN
NT9dZILDiDUEoLfIvXB43mk/YvKo6AoSTGWDbzBlgW+xLRr4JB7onx0ud+EKGG24
sbIsUXjiVJ7hDRzE6/6CZbU2JBFHfxV/9+Andca1Hc97S1aByUVAQMnDF3zW3ebi
nuSRO512uNdJBa4/vrvz0dFLjNl3Y1A5Rmc3JQJPd4VOcHeY3PSBkC6V+Gjeuouh
TqWrCHglrcQGA53OZNRsZpN1LcOwsZfiilqbmdgQyX4bxq9LZ9bxbrqb40AR0KC3
PvrvwuGDhyT9pAIkSrEo8wgqEJFpAv+Q6qOwTaAyRISsA6JvizI9bOXp+klDFh1j
Uml3ROuFQPFOZwy1Z08g3xM3FvrbNgsvEcD1Gc2211QfmAla+C1CjxSSNopbDmsy
KpwWvrX9DSFu6x4sCbs/dCNyzButC+G6nn9qY8prWcwARluSRXztpgnFYiPqFNjM
RClWrHoZSqC6Gd6tMsc6ipCfQ6idnhxUYFor1UuCgiX7Vb5tCMJLYzF1/D3b8YB/
qFcKkVrj1YgG51EswJvvqasvklFATxI07oT2EFz3QDG8Ne6WIc2EonIW+A/0fWT9
CJK8dDaog+UZHA9QTjhizLqbAzzAZU4METJC3cifIWfMreLuyRz4zC0CjooEZKeT
4IUADeo7WW3S/sXrB/KfeTcCZXhOENMY4zJ8fmGYpvp0S0XcKF7L4a7nDlO3MrvW
+Jnt9Zhw19VEM++sW1q5+xydXBATxTWYErLL1bS4x4Yu0wR5uDkBUzoBOITEIraM
KfRCE4+xCjLDhZI3cg9RZ72veiOZqXvCBgiIH3PeczQqg6jIwZxCJybu3WON0SY3
uoGKei8+7HYYMXDr24XLUolFIyz8KVTtNtyISNTGMoAHMEi7QQWVZgava22juBI9
QSC4FytWIwIK8toIpXnCdPtbiuE2XdZr2l3ZeQmwdQXDaQz6Rljch3pC3UiYkhD+
ah9EptUoMUqdIQ99EyaZ22kNW313cZtK36xmvQqSMPey50/95E1lnjd3hU6HbLfM
H6mmCiq/7slfw/KtmRCpfdiaMeyK72+nhO92QV9xRZBzoIPO6u6wSN6fBNnwrHFt
O2XokgtoMINyM03kUQ7IW+37CaxxQsosHgW8Q0rqUhc5dsF5ryDaU4gyhEzRxc5C
7CgHPeONiju91PS+M5NSoHInE4JUzeeSm6KFhIdGnTppnkWAQFnVQMe9g2+YK+aA
2p+qjez2lO/gupf2rB2dExk6nOhrI8KErF1aVVdagCqL32wtf2z1f3aH7DoFjG3v
RPtgAugKuV44Kk9Q2x3LMZmXErrHYCEdXsJWr5d7RkDxAaIs91vITkJle+4O12Xe
L1EX4LQBqU8Q9l9vCRdqJejfXuQ0A4WqvW+ayyhAt5B+t2IE/Ql9vfA2ZGvqzIIN
yhuxTZ1BrG6cQST3r3d4eS+tOk9GajHEjWDeq1ml4+luEd4dxnI7X7lp5Gszxnid
uaeJfvUldPWIBOLY+OxRT10nF4IGvk2MczgEhvPKwNW2aNYcQy+3Fbcsu2c45wlr
wf/9JABZJyXM8fAe5Un4u3PuXZQe8F4io77xDibCtfvBfjcKoDkeHmUk3/Z6Dsop
ckNzbzYS+TQ7XKQfzVYX1+Sp5jiyPjwUV+ZuDV3eUEMu14hV8op4BF2E/uVICtit
uNbhl4Dy2KuujLg0LiXrW0Tk5HlCHOzHTMxhOz6k8x0eKo/PiqjpsakWwXsVjm40
LzWbc5V6A/YVW4ytC4y41ZZY1sG18E8HDV2mcnN2kW0JD7klOaaS1NigldK8C/Os
4Xh/eVhZRG7xQWN4HcSsRpZRF7t5W9br5Be21mpUy72P1gyvparrJXQHLfZSsSCq
KzpATkRwcCm3ektv5eXvr4a986K7GBXkA7ojMUOSTxPHtW0LKpoHSbg0EpAfWCzu
O99goqdZok1QvY2kiUMl/+OzyLgsHPTi77RYCVBLlysvZ/4FFnFZ3KK3kU6/oRAL
DfGoCj8xYEvUx8tGf9/b6ihG2Bw8v/+mGZhmtNc7guHrF0HVo6R1ubA1SGY5s4IU
3Ol3uLI3s7zlVfsKzllAV5yZvw19o0RbDm2LTVqBsHd7fG5th8ItpVDTUzC+DZf2
JXmxYjqT2pLzacoCROjt0SDnvVaVdyXCmTTIAmNkX9EJPR3+n5awQGSUPoxia6R/
iFpGBxRM3QqoipGnGAwh0x0atnyk3k2kcNJO9YlsOzZlRpOIZlSHxDzA8Sc0J6OO
SlVqDzfPilRgKECn4StQ73UM3ViwslZrmLVeEfB9Zp/Z6YdDREhp0NAdgQrYOzWk
TXu0RUp/8ghrOoEAM5k1TMvAsQAJhWmPOaRMb98dV4vBr3fW9GEBv2EY1AkXWWdL
a7SPVG8YbspoUJTQrNmWi8e2gw5R0n3TZkR26+Z1C1XfyY6BSGeBG+EyjPpiZkLW
Rx+UzIo80nilUEGKJg88au8QenaSPQiUGGqFweCRcpoKZ3NG0Tt8vKMF2RPlNBS/
3hv0sU1+gJZ3GiJPMlyltaF5h0qa8xklz/g7gapHm3NJvsrzmLMrwIZvthSz9clp
JBW3VvqhwzJWqlDKkIGZ4Z+D3H7Z+XXAuLXU3A4r+Eb0JqsB/u3g/Yzno493W/xC
fx+J0qgjCXjioR71tnMeinpHImZDc53N6b1oukjOGm797D3CJm5sOHomLOuW4afM
fZKmU36zEqn/erxw6SkLWXiOsbCbRRHRVNuXEGlLhTKeEoY2/YOLeDUjHMrLtyh2
Bs6TweRHjYp3l7KBc8VO9RdPoyppzZXfZJz1D/HiBP98QuIfgVghnHKy7XcVEjys
HQs/eK/gZsOREwVvbaoRlXO8V8ke/ex4NctLD4zMHX5poK1hBVJj2TuKlV4YLe5h
bm+V1r9QtKkeBR03VfPpdBkQs1zfE4w2LfCuXzLOu5+7seIPD2pw+UZUUxGHnpum
D8/ckihc2ImN2hDt+WrRwruP3EHJMHWNeJU6tXBCiDZd6HugcFlzr0PmnM7KWYZc
1SOHVgBfyygPoNogJnVA96EOvJsmvcdgmM/lUEP7YEvVTsEkxIqoQac608p6o6LR
96r19DUPhVQNj/hc+Dthh0mmfQiG5lhQkvj0LAxZRE8jQZT3PfZEDnJqP5wiVOe9
byxbMVnCPCJGFuUyMX4MmZiuAOw0N6kgU2JSc/lVU0Q9/50dryNOkPJjgvrNsXk7
kznmVwZuTVDVDkMBtl2aJMWmEOGiZMemv7+xN8hJQ1HagRbN8ZifykvB40bejFHo
VaykLlpTg2QjTbtAcXgXYqI4pb3w5fZMvrqrPn8Fc3yuqUlIIlAx/Y15RIbpCH+W
YoLjm2p0BGU1n4i9F8DuNker35ItWJ95hGD1zkHM/FZcAHrLEjXbhmhJoKbQuZGy
V8zl0/iD1wYaFiy4a5pHC5uymwU4LQR6cWZKlgfu1gfWHp58Ip92E05hUpGGbmNR
+Oy61DcYybm5HjHLAEWp5SXj/V0Yn0HkztR4bgWG48c1gRBdYJVv74RkeoKXFCYL
dnZr+TUC4lDctWqRjnovNCi2WYfdCCQlgG2hA+cIcg0tMg90LqkSTVtun9ss07uo
jHceHopmUfGcdH9rfEUQTxjhSSfYKFXzJgaDF+5AxUMl/sk/LJtVUD72n4IyQ5Dx
5LzfcUw9ZxkHjKjHZyb+JuzbpsOCZpg1W3xpXq09WXg/Exit/A3HPSeK9B8D4szk
0ziorIL04/Q8ke5C78LrlXgE5QGK84S4MPA2a32ILNI3tjwdUwH1ti2kvfboienl
zQT/pKmqPeWFT3e7qAUewarfJfyJOKVRB83snxiBMgRyqliCjfQKXkfRvStsB1eD
ps8q4MVkbunF/CCNDlGl/xy3xM60qnNts3PE4nJqN7upag0MkuanCX4mUjAf41o2
9EtRfXvfZNj6rV7DzOMfDZ8Pmi8saZ+FWd29vdaLvzjmxeC5LbhEetJ0uGkyny4F
+AK7J1vl0fNmbSJABCB8ImbjwtH2elUQeUHwjznx0ZI9rVM7OqwoQLoiGn/L61Jp
V3E98E7GmTf9O9n+QhBCfJTlChu2H46e0j+kQkOT18D287zQEA6949JR9PyB08sg
GRJ3rgGuyt9U9NdbVZWoNoZYdf47E/SrhCwRr5WlU8rRWmQ/0FGmPBYmmn49nqly
04jeHgwiO7vCOcFVi07IJFTk4ZO8qkQmBaZjuQzgJmG4T5Wt80QKiUWfd4ovHCeR
eQvcfTcXUHzNpxBXl18l06Wg/0IgSCN6RBjCh/sl5a8Yr1+p14sY+PSkA9vKhSRl
DqOckOkhd7EsRddJQ1K0LOr6nJ4NGzPrILx3E7zXNqN/d7SQQZpMPStIMidMQV2S
wrC9lKCeCGUpRcxFDIJii7VQLqe+xF86IE9lwCKnu4CkrBTP003tSy8vbmsAmXBK
R1TvrcwjFfBtt3UMVI4fk5RybmzK6TkIZGuV8MSeGymWTzLSJoaCYf3tTAfg1FBf
ZdvKPUF5uUeh/wxVKA5eajF4YaCGT5paVs5rfhpNqi/p7wCpED/4RqS03pQfPc1T
zFqB0TTVS+LNIf/W3nEnZd7gVrCuGGFBl8DkGxssdftAS1P95MbB51A16/XDrqq1
JFWKhngAEbHh6rc8nMUPrdDd0Vq7rYN+vnjJvAPRF0xcXW0WVwH2N5ZDpER7IinL
9CpxxQ4VG148FrKzlMmb7qS5tn/VLV3NIz+Opbgttz71sdW5/FhCDWU/Y0yrQUkk
Q1wW12ekAPFuw+xd2F7eq9RHbg5O+RZvIYPZQEqIgZZaiBHGVRemLGBTES+ldTuA
5pWxvQcXEulDBo0MedTPGiu6V61iMI0I4776BMCTWKR4s+WCmPJRNddsGP4NafyT
GgWNgm7eggEwUriSlTRt+OwvgVRHVqVai2S73V8I54PgKhvB3Xlft3yHjHVUrAei
GFQNAZL4jxBo3bJsG1diZ0N/nye9Aa14GeDLnGTZ7dnfV9IRdVuXuMC1FkYlLSMU
hU2b30320Ki/u0tlGGvOmQIKV3LfMahX8Vv279Hif1PWMq7s+oS/gVPw2UpZnjN5
c0oPMnJpFQbmc4gpqpPLXwhR1HYsT5piLHoORYCzXZvrSFgXni0N3DS9+rCTb4PJ
BYzoDkp0HkAO/SrKQMHBv4zkFTaNZnR/N0QJSqV7YtJP6SHU+hmhnltoTCtPNeqt
92XAI6e7c9dwEsieXTWeU9fRijUadOsR3y4yEPSoqAJmCdOhm/56Vied3rJZZ6+p
GZ6ubOod7iuSTvlWJ5JsJUEER7ihKq6Bxy4RUEK8c+dCOVbqS06jM2cjyyE2GSB3
9S6L2tbvazCQd2pHo44WOa134IlT7axY+th5GEXC56AuzmlwpEdqmwbozMlGaUK5
6cgkJk76lPbG0NEQOGuMIlZGEFKLSIH2MobN2wDoXyrDEe08F/1WQIv5A3nghyXm
wi+PldGcYHSc1+o61PBJPAMNxzH9ghki4wfEEY1H93pDDTEVZAoZFqn0D887BBYz
hT9jL7NtDBPFaN+HBF/rudrFaA48uNcFVlpssjtpPHUVAne7M7xkREengtgarxzU
/MNq8DZqn7BFgN6eKvtfyD1g/+Tjp9IVKgaz4K378vx/YVkI1chDMdxoX90F8EQY
VksJ7iUy1Ul/si0RtShd/Ftm/U2fnBzum+pgvvTToP3rqlZInL1Ru8HbyZeTbXUS
giPUqVBEeOtjM2WZWCxpEvLMKEGSYg9ZrW9VizfzYXaRbeelBWHSmW1e3LPIJlmt
CYR1j51Kagw7oew/OwYWErvj0hgusL93F2buxv7FgWTC8o0u5hBSUSA9He+s1sKq
OlWPb91p3yTC9wxmwkFIJRtwbOBKu7OdUown1OSkVQpjBgr7vLELaVyLvW4jpuHR
DKLoJPL4fpoK6JcQtlMvdd/3hQQoQjWS1XEORMB6x107zepwJA+hgnpjBgq1dTsF
+YkBbZb5qK2mJaaIha3vVe6dOPkZsy/rk8Zrom/3Wv1VhB5hRNdq+fbOnVIf28QI
2ZioZXzJLtNRf1GA8XQfdGQ3/Sye5nFKVb4Y78jiMhtiCsmIq+Eo8YFLEk/7yqSM
hHEd08OgsiprBAx0oNxejfSrSIrIfBXHiouuxyqH9P2nxL4r6lappUSRL6v1HK/p
F1AYA8twmu7cRGwU6eBbqr1LdjrrnTxOLyZzNOtQjX1ybTbhNEd6frAlfn4lpn5S
NKruWVa+JoWKovB8lAr95hua0kYcd5PNkr6MaJC+J6QN78BdYRvVulTUTjms1dbn
jCXIq70GmTobxv8k/Eur2l2WzgL5LTjXzVG02hR3rSteAdf1vWc+qMHbGOpyCaqe
SrnOmsx+vSnaXjJ3fyVitYrx8kSIu6muHw4Dyjo6odKstCoosOGWeMKDv9JBjHTW
fBlSJrL0HQ8U0kSt9s09zeyPQgP2OWUz9p2ZtrETIEEINlLsZ0m3cZAjDNWqyT/M
BoKY5GvwsaFGB5JqWEka2hoyrG0EUr4UZF6mc8EEJATPIsyYR9Y9yQKwM9kXz12q
3BSlYD0JHZUVMxzKACN95Dbay8yyHLoSheo9xQ3/96tmBw8Yk/WQeaI7DHq2dwGn
+V9bC7UKGe+vdXdce/pyEHwICr3RGWPyumfmIyUXeICHkMohY7Bbz2XD1bFEmV1g
vFxTIJpappb9l1qqILMd5Cs9TQvC1UeifNfToenYJJZ4sOjZgMRCbUMwfANgwIqV
2JLnX4LfOjDj0xK9uJlFERYOH+u+VIAinyQqArnKhVjT2PKrg+J1gM5NBgXlj6wD
K5ZZYpxEdkBYRMDvnkVLqEfcmwgyh9S+GdNpJjR9RRj4UKpou/YZBLSeByV68PMn
VMaA9xIbxzMd/3KkRJSUdKzr5YICQ+OgLSYdeo8OxKBLIDgp6W7uilydypYCoAPZ
p1x23glJh8mkpfiUgJjcMgXIMfchD/RGuja5ipOc+hn+y4N84dt65dRcPQ6viwUx
W+qdZ09Z5FUeuH2BOX7aW7iu/4Of6pZRN3DgPxvHMaO1C2YuGwQd+wKL7HAyUAsu
7CugQIF2+8w41AHuEsRsIH/edhZyH5989f7h5TSdu3ZRu9al8yxSCyETsSPWeXy/
BkpMM0e5g8ZaMlVLqhjemXrG73lN97T6BOA/YqPg4VQISXVaTliKTZJqAiXE6HbR
I1pqEQ7JeQZIIBTfTYQz1jbkOhPebLfWpI0UOoCPO4hall3C9UpDnenjBIRtvuuI
w57z3/KC/x/vfg5X7DF9dDa+KkWipwqZgyn7bOWOK28JrQKcC6/pBHTEjfKBI12f
ZCZplN6k/6RDqJNbgvawjdNc8/9joiE/vfCH8WbKm8cO+OHvdE3t1Fv42rgn6BU6
CoAVCqS/ZUpRI6saBjXhzhxQLsngVWbtD38XCJPx4hKG/24L5w+BKL1Z+pTk0EO1
4MaERF8uFm9/bcZrmB0nC/viNNiYQZIz4v2PgQ/0DwmXOiEFWGmRJujTU9KcUlpa
tEjH0zGiYudanCFEIrytTaRVuSikP1LPAd16hutVxQCAI0sUpCt3nBCQJ8Sbt6de
EqidE2TFT893FWCYdy2QHmz6h0/g3oE/qAaD33mr7VHo2ywT2mEDUPQ54b5/aSEb
XIy0S0C2yJSVfQabFNOiy18/jIhEMwT7eVn6Fky7WURtETE6GMwM+6cjCVuaQnvY
txMCXcfY/HQEyQSYWyEtspOd5Ta42xIfxkRWQV5FPxvyhNdlgqSGNbPZmmFmYNIX
fgtpm2ngXNVrRVfLkxFP9fSx8Aj/NOCTpwd2iUoo6f1T089PVHsNBhgMg3Dlk7bF
HDV5xnoh4sWv2cnQgSug8lS9cRD7KAyCSzrGHU4IfM1FOX16BrIsON9iB3R7V3me
mBTfMzj3li5Zh8VYZst5dyobh7eSwz1wmR6seqo+FGBvl+IRTKjpiXP37kh+5JAr
fcg0fyHPKdYXTAjL6b5IosisumCPrUkYllZLlUt09MlfJOSdrk7tE3iTk1XiFAJp
386DViC2QmdNImSDplMQLDC28wlAykz/UPDTmg1VBYz0MSTL4uCwvxugF8eNrl9f
aDo1bTxF6LD1oTusBkcq8qarMGq7aa/GCfeMihK5hBqr/Lmrj99owKgE1xIerd3o
3HIqFxUzz8mCNeGOI+6NZVfw+pvCTRp0/Pr3sryMJp5lhLNFW2XJ65hHJxWGq6my
b5B6/jTQJ0cUlKRCQXO9/G1i3+xojgVrRFkjPBcVigqSwhu3PQsii7HIoxN2ksBw
L61BDENecf48+awh9VyOol9jPaii+yPno05vsScx2gyBACgSBwmeG5i3O+a9G4i4
Hwcrm3U+tfTOvGLyrO/rTqq8YfgvPw99qf9nBDfWRm835v8hujRyH17bxQ/Ei9R1
O75qhEdfNiC5R8TyRnVZO8rUFiwOaIM2MLqcGjvvtoWE7+hJlEsL84ocnu9Tqno3
VrbnF9ywULczsAUUfoeMY1RW/d82gG3pbMvviPRi26Os2j+hSNVtGLxHw3U1FiCi
PUjpZjYJcHaJkzTI6LWVRMVu1Ee9tEw0/TFQznu4d3N4/ZAIkouT73vEhH8u7PB+
6ektzAOo5eDx42D1As9sFVigjCEAln25g4tnx96lTu8qQNJs3r0XIbJ+kGerldf4
u7yYefYSH8otc4aLgCnbPRJ4FI+zHrfTJ+ClIhbhUFvTNxsU3Ooj6y5+X6bW4npf
qOcbJqMROg/qsZwBNpccwm3o2YIrApi2OCT+rWnMrv6sH5LeqA+BJ73S2NAYu8wi
FTcGGyAtD7oV0FFhDKRwrFvOh7rvuSPMktol5MrbGcXIjxT/FIpxPSu9IvYATpeU
7Lq8GbS3aR3mGQjcvE7BGcGpqREA0XgDt8NZPjqIoXdnFn4v6uIsDqsg9ucPBhVi
OamPfOg/AW4hYDOPa2pxtqI2bYGSh+GMb89mOaBKKPltBkadeVbzw9JBhCyK8zZg
Tf5MA3s90YA07JSTTC0qduNP0RURkBahOdHriiZEFgjzBj45HoxVHhS5vvTmfgtT
r+dv3/sM6P/rF9PwMQ/J19nVFv26kfl8rfFztJrAON7s7ZmoYMpxCnLC5y6wMCoV
ZeBNVUiKxQ3xKmfFO/klQOYYWQ2Ig7blh77iTt74cD1VbPdKLmVco7hRV97RwMp+
VTgTHG59+8DrnfHyqScxFLl8TnQRx+zpw3oSqqT1yyFCgD6v6cSSlPdYQ2/dwQ0r
dECA5tnb6oSnd6Y2IHE6DC9lhjR9TOohjrdBckH+2LUe90qCRmjhY2dpFVbFdSn/
P7d8YlH3kljyBVx7Oa4U3Vy4Cg7kyHnnOG9QBYIGJgCNAx/WtxLs2CxNyY7c9oFY
Mg+EQHmeUz6Fr0c/O45Ojy8KFy7J029WEteMl4r0PLHHfsFfau6UVLWUQ9bK0euv
E2CjA7yaWPHMyGXNyqj3TS7MFaGmKJpN8SDdMWNYjK0ZEPy8hOJ7jGUP9995+nX4
HkhdgtSHmr6W8HJZ+jR03LQve0QITt2zh48+TAZVnPiKFm6HJ04BgQ0gkGQbJuAa
ND+FQQqb6IDd7Rbg3+MWGRWSTNYDLK2lvrUnyqvaBxlEMQH0iWcRZOzHktZvqJ8A
4v0hz96AXAoldzaZGjQWDkIbDx1YNm0aw9k8GO0HJ6dCePYW9vyLcSTLaGGH/kwa
4Mo03VS0VrTwsmUMdQQW2e/IoxKczWNqpijXvESQneZVNE54QsL0gnHUkN+MIsPo
XL81mHR006E4GREKD/6V+wn+bPKRuT3JiYwiG+qQG2E8PXSe7B1yyO1FFBpqIY6w
gXcXS09b77MhELYpe9jK9+2R8QClPqRIUZV0qb6viLfkcMiGOG0wIj1c7OdIQ9xZ
faRyKbUan1deYaomKrp6F5vxK79z94mmfz95pka+D5yxjBMQqPS7GASVJ2RB1BcE
jtZVpkR12chiSD4EZZt6tpM/co0vrdVLnVnKM8enXoJuO3OUhJKbDkslW9X83hl7
QB5LNcn2vJ7C8ouFd8fPicab5+bKbzrCp6gXa6podJiCbviyolO0kwwAqz0CtKTP
CqyDqO81bE2MhRqqlp+F0B5K0L2bkv9jSwsl6fq0fzpNVwrRoqKtA4TRdqxCbCvd
VfhFR2wzXEvawXa4Eawo+fjOUmmnJYlmL8SG5Os7r1TLelVMJ6HbTO1SE8CESGvJ
SDqr2EaMDwgddA6NTxqE/mQMn6IQrP+rJh7x75ugZuEHgTI+nubCptFOyIo2Z9OT
o5AwwfNgIXNsf9acylcTSX7Ow7jdjk3Mrj8/tu5N3qfA4USqV7pph0EdlwTUKo6K
/ZFD3P9oQ2R2OaL3CdTMXmgsfDC492OnfyvOoTPN/oAjYTseORXqjPtIH4rMSRIH
nTSU5pejb0pBsAKbBp4wIQLhlK32JnV4XxS5QgK2FjskSK4vtN+POebK/5EVlHm5
d1CmHS7CFjT3jT3du2UeAbdghAR8dOrDKeHKH1L+eqYMI0ujAcsEDLloEtQtsLOk
CPiWeudsGYzwqX9Qw/+qEg5yjqf2sNuxQL107QA6KtRtuBJgn3+7N5XHPj5n+DT4
iCOm8VjcIBpvfGA4GPpD29I9XIkBLCMxWTMwxnRh3X/Ff4+cVFEJVlcN5lo5mMdv
hlGaUqVacu/4z8Dvghs8DpSd5Y1eYRvms94L9pm9LlDhUrv+InhLVpRoT0t8grMs
mavfXQjBi1EZg6jUMoO4saD1sLvVQm7+CrkKW0IP2n1pGLLVMXXuI4zBmG0NZxOM
KV8zhZvQ9eQRnxBHVsz/N3hqXy431w+D6xxgSZFQUL/k0/VBPSElBRtQDASvAigh
jrZVbKtIvY/PWHOcWZlQehL2DXWufto7iCZhCZeuz6PnomHGNii96AWrTR+/Bkff
QnW70KBOr1NU2TtEPB4iKIxWLHmjYAq2bXyct67ZimlzdbJKLXfbioI4zcuB6i6e
euW9KyjIzucAtQNuio5VgyVvenVhnNwK6sBSXcjqNE6aHKo/HOkyQWUTkovkrOXO
ORvdQx/zHsRiNJHrpUu1nkV6ZvIoPkrzZ1DLM3AL5zDwbmxyacoWMgCl7urZxZNS
FrDNkFJg4Inz1eXhj6/MZziMMLrxtm3OmGVTDnpFFuDFr++uyGK7gC5f/1nEdMuQ
Fdq3xJJ77eiF9yn9sT27TpFfpQDQbHQsLjsPBjxIcLIzHRtyY5FowbabCYMycPRT
c84Ut8+Bz915JHbLOx+AolNVm4Pd3U9jwiV/bxxEIkReI7QORMTFOelctGBZ3CMx
pFBu22XaCBV40pDVg72/BkvwAo6qb5eZ7NlNRFsZB43USdLHU9+jca4XJj85A3aM
0HEzQoUpYsoca5hh4+xiszgxKS/HvaPjTbrCTHjtxwh/smJrzYhJ3qKqxIvwksUG
1/UVW//5wHau341judWSR1MBaA5WscWAWpyFk8SGrOa+naW10bGIKFHOZfjW4Urs
spo4b8KXNmtxG469VfwpWH7Vw3H1tHLMv5FttsAEUTHhIhl4ua28XtGUUt/klVPO
KwBs+qMJiQBdkjLCggA4nlZSff78rMa6yhweYVs/J/+GYklOKCkHIcKqmijfhj2W
7Mussgfaxno2/Pu0r+bVf2qtb0XIKG6Y2Ze71wNqiA+pGhPZtOuE9AwraGacgreo
n2PQdFNVZEKlq6t1tng2Vc6oSZARrDWmQwNFjkV6c1aAD2vxed/Tp+g3OruMXowr
bArB4jmIRQLJ1k8sBq8UWcBUfoQEq/LwpBJzqhlu8YHfKBXVZk+Bv6Vq8SdWG/iA
oWUQRYMvBKRtSQo2/tQht3+Q/uJ0BxKv9GG5G2oj2yTKXX2fqHRiFIE8RJBkL4uM
RsVRV6VuhmBOO1XSlYjR+m7p/J97M1o9WfEOSPhEoRZRppP8z0CYgM8WrHkWfVUc
+EFyWph5iYEEvTVKAjqFJIovWu8OtgiffeMqRRIAwEpB4NR2/6/0ynCBsUZlUsRk
jdZyZwYV1UDsg82TfCCRTF/Cv8JCOAO5mlwsuCLEIYFLDB14bkZlpphgZvQ2wV5e
ojTKyPcZmYReKgeYTtRrmxVXo9o96xlJmlINWZMv00sm991SZqjkGVyEMX5icmRp
PVZYkdSzYEye4ThLUI51k0/UCgSfPp9rQ6nzlBJKgmkEqLyPWBRZOzyAHgGhfCZZ
vhMthoCdLf8ytI66Q4P3pb5su2l7HH8RBJ4RETY6U9uROCh3Nwc2IHQFrW0icd38
x0z1SpbSEvdGcKNP/WLEJ4gVtyRGzc+n0PvALLKUIJsWyDtkd1KHeTE4otK5guIQ
pkyMbsCKwitXzbmCjZGS+IkvMCyE+BkE3yoDwsHp9Aes10iO3CZOn3yDrGpFnnzc
wBG3XrwcJ8vau4wRdYfjpOnMS7PWvikNTEVZ08QRcmzwPZZFydUscienwkCCZ7v8
0tKMb2j+nwVBePPcbFqiS3ARit6D2vmWCwLhq93L9QEmu09+J4MaDCEMhjydFe0U
5oQi9oFzKg0N+gbfxAD9iUAyQYjjgSPUxzptAfphTjgKewOUpGwKfea98j8XujIb
x6FPdv+oCrQwCwzHS9DGVWCHBIOe0sKtprMa+DRVul7OzbGALjGeHo80RY06Rnwc
VxiPv8lhfTTb8ciFSi7neCtfmgKvKi9jxbWkt7GpAa/MXXKjwmmiIDRUXZ8rnEU+
rHTTHklE8s4p40hT6byf+bgSR2InGUghq2QEM42AtlQXuB+/HyS9gk7NEv6A6u0i
nHMuiig0fgK6CBxZCXkdHyUqD7vSCYMC8GMirGYtbb6pqdfxNxxzllIR3w0GrSxl
/QVBR5vgyBWyPea5iaYgqPm6RRwgasdSx4wvCXl1GtDiCzxVPhaOiVyQEuFbhACG
lSR1MqmvSgM0zxsATUYKODvOizd+EIikWVnR8SergcrWljhSWyacWKV5V1h7tyd2
PzfS/ZQuD3E+tWK3eL6vghm8bbWqqUCwjoBPpd2I7U8dUCkXmxcwJOXR2LMiKENZ
vXyWyaYC8sPNT28p2skEzO4TQji/fKqbYkVS/V4SnDpAq7lvo0mB9mt032ny7U2w
9OQRadBhPJ/6r5muuywCZBZsNmwUe7+OoHI2Mz+wpIMImiv7qj6N/Vo7WCdbsbNv
Bg51u96HYWDHLeJdi2mw/405waHQK1VtmN+SMA+etV0j8+R3x+QnDjcRm7lLpXGV
BRf4YdSkb4GVbu29W/7lEhAJ2Nt9DnYjTpWUCAh4OUUE7qPGCMbZ3QKBOJ1LOP9V
mAKdkklxzd0x38f6zQqSGLQd5+ePDfC7asVwkUftMVX2ttu2/Z428TGx3nPUIlTe
qzr8NELpjg9JwNy4VaTyLUPDrnNjMrIUnttL5NJ1l0p/ZXUa0iNjJi+eK/G5UHHP
S4KwR/ta6pnC3Yn2KDt7JcXpJrreFC4lHf3qhB12BmkItD12JkbURS5PR+ft7A0H
a2NaIGxRpeO4tjEqECCUlwq1dpfTW/xDEaKC9reDtbxnxmwQ8nA4KGElQA79Rhkr
iR7yjJ92ZiJbZu+A+TsPslhQ/dYKBLKrgz3diIYJmWh04b0p/fDUNdCWpJInntnT
FRnD99KHrSvwNPjzz8yeu0QC5AEyDuGXOloQsO7jazakFTrt0QD7Uig8PpWFraMb
KHAaesNi7varDj4wDBzKzFiyvONakfH8NI4o9CQO2vrMx00PIC/zsjyZzvw96Opc
AD4uQ8jBYlllcxxRAAaUk2h5XErNKsDQa1RpsoAogJ5gH/MNIjWozX9i4mvbHjUb
al7JYBOFxEBNjY5fEdwSTrczZcz2riskS8YeG9nKXbTWFe2H1PE3EjtG4i0jBNfk
rjz8z0ADMLm3FnOSoXXBUgGHCGUuviXoxwESeChs0SHxsjUT/MIb3byQt2B3UTtR
e8lvGFZnJ+KKz5HP7tG+hV9UztjzHLVVOxXlQDcK78vopU2ndbiaVr9L6LBnTDcv
7qhYu9ygjdkckaLhg5Gp4MAd6DcciZVT9yZ7bKeNWIMU9XFZryrVFQorw7Wwvk3y
ZIjFkzZLToa5s+UlaW1eTPnAdbkDBJCjfXYDjrKD117pimnoN7VW4/dAKru3vV63
ZVJuL2SvUtg8A+FtbvoBwyvgkupMeGOetpz2JYIimtzFnqB1cTLYFNl+KJLNAkfs
l1Y8AjGRSx2qYGGh5X/XrBk2MTKznVq//nODGl6txN84YPo5Vh4QRMF72L8K0HTs
MAwSxwSEOyzPN72IYnG1Ci13niZdqq8U6zA/N8A/aYOhye5VhmJMbW5H1TvFzr46
oXl6MUKAtGop9pF2Ke8dDS2CahTeXKVXp93+nuC1D2PCmbgZmnd9b12gfnU5M00Y
Ey1JhCzlfrRUXQvHg/ZOLzwm+Cg6UObQiqmpH0AcdHErW8wZplvyf8MVc+waDiU7
2Or/MgIAPTxHXFluXVyS5KWDY8sciXnrVElpmfjT5fbPA/pwzo7QSXcOl9mpiSrW
kCFmVpvQlEBRmDl/Z/cqtdEDEm6dtjL+x3RYfDJF49mRTqkl2vt5oD9IK/NXTxyn
8CI/610bHw8cDzXbEMcJAHgE7f+h6a8cXiz5gzCCrKMzJTPSKMNoefBs2n2DL0mt
eEqbJUbiTO6UwssYy+LHWErbuCwX+OlFy1kI0a0jzB0EiD1JlyY+TshHbYTTYwVJ
d2khs/L/RM5TLf6BKnwvkfLJsqeHQViHkR7MdpFCz5Je4ir3+lif9wAC9sBiYjLt
5TYZeoIIU0mRO7k4cqt0eqSGe0u1aYJOymEnijfsPHwwB2mUvAoL1PdWOVZ9kU+R
d1gNIb9OnPReA2/mv98jvtuI1VMS14R7evwrbQ6lIWoZ8YerVs9i9ql8QB6/wAj9
WbTs7og/NaExzeWo8SpTHQFPNQMWQ4/oXLy5p1aD5Nlu2ZPkKsEjbXCNBJ6xrZg5
H7eDNZV4tnNXMqgFt84PAo+GxYvlqISaJYuFNPxiA5jx7E7m+exZhpiPpBDqxFcH
1p3cZI1jlJMuIpTZU8orJX+crPxeln+bQhaOt7QfzsFr52cAabDgCLzQ0rrR4ZG2
k9petD9Yc0bByjQQu67ro6fM89Ub+4rJovLmnbBK7CDHkre35GqP6Nfwlpu3FTn0
vq84qaO5c1/IKd5RFCAuSwalC36Rxx3BuQXcTI02i+8s2+DrR4yw+G6gtLrwmBHn
PMymaqh0s8dquDFMk8PkCbNiZqoLqrZMbSdbMjhPIkB5pPQbjarpJFpoeMTHc0V5
KBZ2tJeHTuweoh/YiZE/ojfd/4HDmBWvvSBcIe8Y65voaZUM+DJH7IZpOnNGC7XM
bG90Ob/GNqKZoQdVCZLVklCPb3KgUmI3510IJkFlrjxeAeqkjnkhdkoVaPIsoyZM
6CT/RKs3kq/UGzslEbvCd0o4F57rdKTWfgSY1k6dproZCELCKP/4dSTS8gIPfYx/
rVoto38epQXsaAvAtCi6l/f7SSfVEdQvcju/x1PAz9qFg226n67xPle2NVFctAM9
HmBs7izY02BwOL9i6Wj5rwbv6+qf7/M4NgbWYcbuYNg+mLLmx8H8lE8QeH6u0oqo
UJdvtfZZDz3NFHViDXv0et55reUv1NZfjjyKDTc8GuW1btbt8QQldv1hmhnL2CTB
/dp6vtSmE8MhgtOi058K3MuVH6JrABISK+Wax3elBDNv+o84KTXj1yVcyHQSJjRl
Uyb1n6K0tqoIR2e4Xi2nfKkr1vaVYkIdSLA+4E1A/A66d/pYeXHCus+NFqzYmsG0
S9LVvdvQ5FJ1C4drLu5J5ncSbWvVBvQu068mdJyXy2dCjjdTJdHvLPuh90r9usrl
Ict7Linr48UdvaiUUFkrLFZLcEe+bKDxcrneN0Ptg97px2R4Qt+d7zedBYMkRV4f
ut7wSvD9fv2YK0SCnUeE0eh6hqF9ipPlpIi/pKgiT6YDSTOVqC57pGx+bJaJaKdP
T555SxXLygHIdV/0uwjIS5T4Lx8DXxOaYA6DFcQA+TEUUMAfjDbtsJTZSDQuDBcZ
hXktdqNscFvHN4Cwljk2nts77eQffO6zPslerA9//cnS3xSn8b4feAusa9x9bUyd
wLvHcUIu/0CBFTszPLFwhqj/mTp58o9+bejaPLQXJJ45ADDTyIDq37/PF9+hS+L9
oXfYOFvSH26vTTpDrDO9Uhobi0yuHlmqhbNXJeH3xguo9cSkEYU1M2zXgrvJVRjo
`protect END_PROTECTED
