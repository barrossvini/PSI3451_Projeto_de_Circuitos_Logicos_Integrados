`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hHsDDoqGWQL5BzIy7AwnVkKQA2nflgH9t4xZaKimMeEvgFSKxAiOxqeH4s+q2no9
cC9PZ83Oqb8hheRdHWuN95GUz7nyz1wNoo6uVyXjq19YbVoLWNYx2+TOLFJIoy0D
Q4xfzGVd8tihKcnuEFzjv5BojpugNStLwQsu8wWL2Wjal0S4g1zuAnVDf3fkzGjC
4R/GSfGx6VohHZBAF7xigTHiVUSdPULNdDOCaeaz1V8N8RyF4qMq834+4c03TavS
hI5iJtKHBEtj4ZMmZmRYoXMyS9GHMh6+pSIRfmRi355OGncATzJO6HA6wXx50O+7
6v4vtgEZ+AcMds8EMdDCn4qh0FdW4c/HuYM+DXyOL4C+KBTmcL6NU61ay3tgILB0
h92sgINnHLJVZW2FcFy+es/q0rap/Nd0roO4ZxwCFeN5d3laCfWg3byMta8CkE3p
3PU1j4ijPfRjqgYDgb7EVmNP/2Te15qdq2TgD5HjIFNAC/b77/WRB3r8X2jX4ykJ
/2ilPvXGQz4E4Ts+VOLacUgh5JFuI3uQUhMwCk0t733yFtDyTEbnrGOBVlyxXXWI
Ry1nR13th+7yhnjctFZALhWoNvuewq7F2duIuPFL3lyVfwfbFNMpqEKOX2n1HDyO
Oqim1hXi5gHp/dhxBSnuwtq8ZDP7kbC40laIeTLFkJy7IqbTk20vSOVCKTg2zail
qSQhizMVnlatx00mEtpZIibpHfPZPJGj4gRcug1kAkUu4UvDFKW2VNpn1u28jzRY
IkoTmut8NOgVvWrsDvjsV/v3V6zCSbEs5uxJIwJFLqUniG6C087x4O1r+8tlF5cI
ekVB0JAmImHsSEc+qyCRwMiahr7b8q96JVTWWlCnNAm4i4UwmDD8HdYmAsNR2CAj
CwPyON4ty2FgucOPfwNkP1dJYZcxcnGTcdaWVrYJ6q8bbxpoxRcUwSOwLqJigBqc
/vJDPqHXJyAuvIzkfyho6tKAFg0ummGCGjeFOWpcoMjUMEJrpN0JluCkcQn+wEQF
eU4PYrbRIZbmzZU6Y+fq3jd8Uh+khCfIqx+/0eeYTJaBZk/NX6Uc1lq9A8hHAHYM
dR/pEnIM52NSWnMmYBBN4FU7JjeyVIhqox/DH3SC9UK8Zljq2FfCrqsj+tCelqfd
`protect END_PROTECTED
