`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Q/2kFDBR4FiVE2FaF/5WlQUiif4NV986U23nPixQSpFk0z3Dd89hDm4+7mCmXZn
rOiFbbK6Dy0sFTFFT3TuKwUygWMbKsJa4o19VRP+hOvgjv2yADYSEKZxDrorQz/k
7w0kZuzz+bJCzWAwKIqWztYg9a3/GVz1zV46Ugig7+GtmnLngi+eUdMWf7j2xH65
9bcvmkVDG6faXjn8H4uokVlaijYrd6yuRkPS8nbnhI6Mvdg3pF27iuPh4NP55gXy
1PExD9zyr/nxe1fcsdUgMAWNatPGhp/n8AHIML9/dUaF7xCAJ2EW4z/WA9xK5a9l
EEvYfVVUkIKB7hdupRLWCJ3nHudnjVdgJByHxj8YwJ/5OO7a1TKgILhyGAGngf3i
DfxjIvJTcm3tjOn16oeepx0ZUmsV8LMZ1VGE5K0lDLS5Mcv5sg1LrlhhHx1wbHCQ
L1fRS8Ydid7ENCFH3J6rZbxV2l41/LFS73l07OvzgiHHVbc8XueCNyIta1UtGKAi
yBF8vg72HJB3WFAgqlz2n34ABtJx1JU4QIGiZyhwkpd564iVKPjfSTgH0URl7+YL
mYsOWM/rCphMb0UobovY/bVNYvUJylXOxi1WtQwt2Bgp7KvLYNEGhsripyyGeTqQ
5NjEg3jDrMDwCfhPoriz0CzdOOWuddj6KdszDK7Vv8WYM6yEEd4sYNtHnDFCwbtD
s4hAptTHO6pqHz2e/uLFPMVmAT6sK68fUi7GXg9cGKCYsZKzFw2g6e+V93UfgjAF
OXPT4EpQl6S6lve/O2NMapYgjNzSR4oGgP0KO0hUv+k82Jxi6fIgfHo4vBdfFLsK
3LP/qTXWOp064qD0T42vor6qh0D2RrfLLGtg+kFtEmjIECrIEA3U7aLfFdeaQSA8
2vUQBHZmAaQU3G7pVNb+GVbnQZCxIrZXkipjyz6ldxNxWhoDX2718ZkO8+3d4zVH
`protect END_PROTECTED
