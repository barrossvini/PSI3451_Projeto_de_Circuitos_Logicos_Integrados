`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJNrDkRyXcrE+vMGxJ6ZUomDyCQ1AfM9KhO+n6Qv6/Y09Agtz3FKIsogAJ0bE/tz
khg5e4djjgDDtiyK4R5rN6Fyg+MyQ1gVdN1WDwrBnbYiGOksjFG03Y0ZTNUBJ7fR
Q6xpaVNxxi8DSVZhvz1Twy66315DSxNAxMagqYLXajTJpFA3FgEhelQ0T08X7NRi
CoZBThpCtuEpLf4UFQPtAd+kg2if7IGxFdNGoGMj7Wa4STJ0eGaBqhv3s0Rp8Z8c
MINKuL3PEmUD54CDAcsPxUXxdxB3YbkYjJ4iFzYYqevCoYWAKkJCvI2Al+vlJeXT
hEfis1mhfq7pPofC5Ls23FdrHJo9bx0cecYDZg9+2ftXYDrAG2ZQZz33tc7TaPnN
M7j38OuR6oDqWwCPbF+EXwmt1HDWHlD5BgfZGNWDx7JHrRXqSMup9ecB8GqllbPh
bS6v2PnSuED0fJLoT1PFsXMQMMe5hK9XhZsEtKdu1JnfWa+uLZgxFj8jx07GKHfP
Q6uzvceIFx4MqaP/8/OHyJiZMorq2HH7+OHwy9Emxzg=
`protect END_PROTECTED
