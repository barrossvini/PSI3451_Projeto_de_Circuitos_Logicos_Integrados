`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z8/NhEbSY0Pkkk5XMB+JnA3SGdA7wUMh233pmymRNOPtWadsVMysdetxNiXNCBYE
ep8FhHhXZF3XgiyM1i6tGzl0D1QPkqG7TafgDb3Cco0RkiGgoNqYwUdjvlXrban7
kTLyRt25MCh47wdeI9rdiKnay09jXYbKrvfuoJjQzE6Q7s8/BAgLZYZtFJFRZhyp
5dmLOfG2+72AFQJucNR1jVw4BA9Z44Sf9JgzfLuTixI5uCK7fht0hOo3QBGiekY2
5+CP7DYAlAOWNPy2/cZJ1t8NuvEo/lldj+JbM/xmarFRfK692/POULDiat/hXxe5
pWEBKOG0ZOx4L27mh1zSjptxZbceuslCQvUkDrmFJe3V0S7eUP7mgQtzTrFTBIX/
MKp5U1UKaP+0KYRqo65HQZE09zeBO/kmZETF9pguJXx1+nyB/QmuNssCH3TcOmnJ
I6PbVH5ODBX1YfzlmrBmMElRy2DHT+YaWYtXmGnREP6qmOPpK1OqTDrAMT86QFgt
Z+Em+GVxrmyZfHUcw6u0EG0gKXc1eV39rNgP/RJRyBuGMNF5JYefvfvq9BNORy8s
ptoQ8FxsTWeZCqizU869rKBBEh5J+Uqst6AJ1312xU3QGPP5SeHY8x3aUW+a98se
GAsU7t4B3YlyK4SwMYXDm081MEPYFQkv3rieQXMSecLxySyUElDO1f5M0opskoKs
ujJ1xPWJOkafzRzTI7PFCWtrNFY/X65hBymC3llFHFd7ZetQoxPHpBjkJb+JV1x7
4l1rIoMwaWuDzgZB3CoN6/FSPF0CfVPq50F077JKM+2yThC22rrssHwbUaLnA/f7
3EALX0+HcGtKp3tcQa84FFDht3KEnGQoC8mQ35rllBOCr+Ki597GKODe2oUFQDVy
F8KwfVS19/+dbRv5t/aOVPsm/SZDH86NKKDoCd/UQHF52ZxuNBtPY1Ar67wTSVl9
G21g6rT9Tjn52zMIT9wpgDCFS7PYwRX+IuCDB7IPH9JT/C8m63Vi8GJ19OAmQBTb
`protect END_PROTECTED
