`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YUlIAH3cFxl4KoUeQNB2FDevPjc0ADdVtN06JhJUUOrVPPWKx0WNAZZGMSi6GlQi
qO8oASRpC+tF0r+dLqN8DjPdaX/uu8LvJMugPkiO0ASYmcLcuHmF0Xj+Nv6xl9qJ
qs1jOpZLNF3a/KTT7lQqhByt3Ofoga4Yj9wIi+o6viqA2cpK3Sq1m4KE3iGRXfrI
24qGx9BZbhU2g1jNbOBBinGif5KZC15PoSOqSv+DQGEfmDPZYFOlSZzwFIYTZZHi
QIkmAmxOLLBfKCDbXDL+gRdFWmygj92Cw/UCHzFSlLD9oOdVWnqvIiXkvR3OQiTK
WFwar9tq2Do4WsOLuW92jyfY7JbKm/0uxt+xg/Gu1izKXwzAd980nWYCeWz8no4q
F0MsDiuxVdHOiqdlud1WRCA3uHcR4OgDc3POc6zcxTAPIKezdO+2CvrIvjAZRFX2
VTGHIN9HfOb0dtNPQPlt4SEz/f2F4nZYj/WPmg3Dfx7kyclp8X9bLxaD94luQkz3
vXSfjRTVKgj0Nrrkl58+d9Ni5PpsrUAW/I3jbpMxjiO906Z4fqx4Iu4kXF5q8ejH
Zwv4/4/65ixOBpXQ5Os9AmrAIQYhh4yhvqCQmOeBt9nhOQlOn6V/2lOjZK309qQ0
tZrMnLXogIG7r05MtOpzMW/CozSm+voo2riF5Z5ZfL9uOxjki5Hn8oWwxsG/AhD5
YXBSsPr+n45hXNaPzGIp5yyNCoEdzozfJXg33etxeUi6ze0hfKP/fs7yLlLDdzNl
lXMMMCNLHfVSMqS+1wnGK88kY7rdgUWr5QqtjGMWfcW7C8+UPAM/aFhtpKOiHAr1
oGossE4l4cKP6sleBzbKgWRziNYYqDNK3sdJsTbsXYN/ipt1BA3UFltZKAmcnLF0
6VAYXFAWdzGoeImsrlNfHd5U6nio3eCNQIWqJLE23ZQOkewBdJywZ9OHtSpVVaz0
`protect END_PROTECTED
