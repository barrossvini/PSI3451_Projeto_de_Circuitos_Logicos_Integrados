`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KgfnCgWzLPBz9xDPawcMbb8FUffTRsxbF/GYYutnFepn+7uJp11f668EnOZAlVYn
+OQaHmdVVq6ovoKsGUaZlqcq037F13orAPj8MSuf9/nR8+6YJmQvuvorP96L8Y9G
ahG+CL1wnRWt9Fdbdf4reRJU7zeeNToiCRe8jtjLDuirfXMzmqhfQbV9qaN3ktOr
n68iGlVwPDYHikRglE7TRxrXiHrT+FvCMoVnxWDUHiXonpY9R63UlUBeaLOSYFTJ
pi0/pWIUJZKRfVfE/bl+RvAbAF5vVwhJtJGHzu4DxJU6wcSYgAAsgKIpXaUtSaP2
Fv3BZXD5XJjJcdCMnORKrIem2YRYkKc14WxnLy/hdQAr9Rc81+aoDYZn6movyWxP
04V4hVhNJ6TGW/ZbjDwZyoMasNvSeGK2EoA7V1ffpQlz6LQf82ushjOgAdM4X4i+
IbKJSJ+nWjIR241WWCQgjSQ+nHPLkfuc121IaFoH5qAqLOHnsoLCCezOYpAaKuTF
4pYxVVuwKV+lI8fqe5L4bbgbwyIpUDdLCmG6BFBnTQVp2YLIb+OMewMFZZGV4j0/
b7DUUAERt+gop3ugtBVhRGWBnrv+uE6fiwk8+lZclTiNbXCMU2+jxnF3XQoiKrVX
qaIILFYBjoG4fBhWCSyXpUUNiMTRfztQQ4uAdE4TxPA/penziIyR+vDPqV2fxeoY
nYn6UFrbdm2VZwDAkcXununWixr3DisXJDMPeHJFW9yNCXWy1k4FgIl8+8wpnfjE
3lX3S1yiHPiIQZ2sxt2AAqpJZHjDfGRygr3hO4gLux+gVQIsLW6d3elLX2shmAcd
cbveoKwvQW+NM/caGyHpNItIQ+77kXTJXZMsioy9elG9MbLOAA2iKgTYkNzEFuK9
KpWuLlyVEJ+MUW6iV50eVLtMoTmoyrapG4rsVh/a1ZNbDLmIsZXckkB+EgzesSNY
Z5gjAl0v5fQYLkfoBrJAdBJOZs68WmHeweRLnEQhjCobovwEf5VP7ZXxDFcjaBLf
5cYtbbS2l52EP6JP+p12x5FiuwKQ4bwRcQjhi2DCtkksZDz4x4EbOwn3rFV+k+EY
/DDvCtszybPln3fEj3A3A5yCCCp5gDyvlqIxpcBRzeczhht6fvgAn9taslqFucdj
KaiGd2QN7MBO0EjtUe1wRs7F4p/Z6LmtjI29XwG+/mSjnr7KaoQ7DX/H88gIlTT/
IBK9rJKm58Zs4LRx4uv41Ax06xLCCpebMEsLk+KR5p6TtOknTf8gaNkWLKnJVz8h
UhcyMIVKuEpGrNBJJ4cahq1ta3EROwH1e/8/3sxMPVDN9/0lbkQRO5XqTBLzl8Bu
5a+lvOdS/TZnAm5lycaMAQVaHVqdF9vx2RsDxIOJd0qfHFRs5+UgepV4ERl+cl4x
sAylhs8uH8RP68wJH7d3A4A1xidUMDmLKSF6cpC8Qtt387kWGeFadiB2gzkcEzLh
x5IBFDIwc9bT4tngjLfyhBgcCLqPdY9ArSwJbgr/7cyv4egnWoXRcCl7rNa1bhTB
Ne7cxyGndhRlfehoNM1JMMvpDsnCNsN7xiQEwFdE/oSOLzFZzgXmw9BxIanzUfQh
26WuoCxYOxLbF2cCSH2JX2/Qv54UMoRCVQ6rT5uNP+Sz5H9u8eyrxZIZLS2YQ5l0
kaj4Fi32DpGigK1RhrfiBZbx4oXa94IXfMvHRHvv33D2HsAhjaSGOixiNpMSiZkv
T3faQ+/o2MkTjGmn9kWf7taPNOCVX3vLAonChUZRMN5HpmUgsXUQFLsXuvKR30gU
eH2MjFn7wLtkqB+87PYLWGHRhe1LhwShmVczFNwM/I69sLtaZ6X6W4pGr9Psvnzz
CvvuU13/i8fMoIMF0yuIOxe9gjPNtHRrhaJevG2JSjmJC+9/KtMJTa1RL3HtaAw8
DpHDDL3kB6WnDYPLf7P3jQhbHqluG1Yd57xN0auoCjKnPbHSxU2lTQS0+Pn2KupF
DVjWalUMaKNFnbaQLl9bzkY5SDewBHiiwZXULNRCiyz7ZeBtJqxjiqH/+zNRDh0E
LErIDiGI77AJ8pJPAui4kuuc2xIwfaJGsnuXkW38JJKXlMXwASHWi2RAPNuad7Im
F2BoyuOM2jiNOzX5Ufm305/pa1taAG7AJkM91iweS5qMb6cO/6mKNoXTFoIvVLyE
HejrUCK+zVsL4dks1gcO1c0f9x9SyBq0K+zObPxRm0109/emMZFd+S/5s4fyVY1K
ThvGohWdGDA0EcBF8V4mS8Z540aVEEQElOKZfX6zk1qI+KVlnBKxiVZweis+D45l
cXhZ82s3rKumlHExBg1npbSGj3AQ3IU+AOD7ybM3r8HMzCBeIcW0RJ89KRUZvg98
cLvpw2fZKNZP5+TY5Typ6MFJwjXvhk//08m+JaADxvytHTAaiyROVairDXMuyh6k
hqiQsN9xFSCEmFs6E64XoO2XwcI9n1YP0Qc5OghNoSiuoa/IEif4rcxEI6LBRfMk
5bUrF9kTNBJ/oB0wE4it++1J+uQT6MqIBVOv0Q0uYFCI5gymUZz/JVnOClJXaQty
H7UwCh8OIwvEh7g7Yg61CkNoZL+DzPD/Nd8lxWK8f4FZfkLdmJsdTO8EW4WRHWL4
XJBhTs6RZiig6JsgEDamPX6p/cnS9lhmtxcnsGxkNkCl7S8hsonbcpZxEFEr12sn
Qvc/29PtpHwkrzNxDN7UOz8JMWqCFRTWG2IffmPlnspwWdTqbJOLSDLfsldUM4Sy
A9xLcQ2GB8wZNbLuUq8+hZfKytKGe4mjsu8gHU1mc448zT9U0i5L6VC6c94tMstg
qKKwgCkLnFw8HdEq0k14v521S3Z24LqCVEaFAeWnOsZ67Yb44BX9Vryo2Dwasbq6
whIFS9qMik9E1eXgjlM03r8AA6uia2b9+MJZU+y0paf45qOfpqKFw1yaQBg0wvyh
w5nnr7iZqZLaiInSLES9uYKWbeldC286T48BD0AXwBNqP1fmnLSvWNhi+Oq8lUdC
EsOgnBIZIGIyX0yj5pLnpVXMCxd4RGBk4wYCJ5sPnixu6GPZKCbr9K8ISwK0dzzN
hh1AMTj8IPxye5X02zJZWzAi91ApbOAQcGb8aMQpCE4kUboiqUvsZRM8SadWyazf
BrD5ElpS7gKWyS6/8Li9exjDClA19m5/gKJiXSw3wlzYNWWWolcJKDyyi3RUwpaB
B8pmehIU9CIJIvJz2FB0XziqH+/hJ5Sr6hhNWmKZnIr67dNxZy2JgkCcuCm/t59S
nTzprsbGTzjeSkvWkzfxDfNl93FaostCB03qbQ+34yXfDUoRnC9f7icZMIaac1qr
4RhePoGgj1z1ZkoE9f3C10gYTcDlp4Z+f9AiGCHoTzOWZk8D8aywR4+Yhb6j/h7K
9Edq67jPIyZkr8DQK3xMkhVC97BRCLJK7VzWu8LnNYqGKvVhkCAM7XYaEgqcUZ7s
mU8yhDnKM05jhZqec5lLJMOaFFkrEARip2sUxCUyHG/ajOyh0HyfEUXwwjTOnvUE
wjq00gFtAqsWi9qxcK8zXl2T9jrwpEAul71VigZJijLBsEMJWcRLFOS08LYM+Gtx
m3b2JfbGqn5UgyXqYAheEd+Hc/CWx/adUGP7VynwaXZ5gOLrO1G8JLqS80CKOhcQ
F5pre8qM9P1+oikVedDrEAq4hERuNwtCa8eqx8JnW17PQ1tIExslGlB5gfqr4D38
01By1xKo1hiC8Q1O0VhT+ZO8MLJlQtsQrR7EboSW6P6rVPjedo/UHXResS1AJMnZ
Vme5/0A3fMp1B4gqHTLmQm9/9yPng+6siCXzie6wvcj5U6UoIsePCq5aTug+SxRH
Zn+7ZtlzjeIzxOe5zw0tg5I4FSzkJHg8PxxQCIFqltekVNoBdv/+t3/xuid6q9n2
lNzMb5e+Kmm6pZXnJ6m83T4nWtN3E/M7JqgTT8N4CKSmFBP3xRBNELs5lRAJU8+J
az0Mr4h2vDj+nPZyk2VpOm+Qn6+fIrMo7kR8bL/uARbR2adGwdgHG/HgoZNmhbAe
ekALOXocyJABrAPWQVRJPaEuMU8vSaqMl3iMuyd6lKiDvSdCTHQAFAeSsZWXnmjz
FHG+3c+IbK8gXBsVICVKrvNT/48PUqGxDvyKZSPR2IPc7IYenx7VRdkpTmo3Ce19
5A4josj0+FsJnyJrODqavHsuSkSti1+tXM5R9prLd1oM71JnWwnACGp4dj6HOsjw
B4LuwCDUFn5QCYrdm9TWYsW7q/IRRz/LXwvgBqtXDaLXSAYJja/Ip5I9HzwBqobl
aGtQF0RkdI338lxsjmX3H7nl6HJdKh89xUpOoF4Ed1HbvmEVDa0SE9z0+0sW53Gm
5mRHTcmWIbyh0ZHqqi+Hgw6MTlShLHOhKLG6SuncG5bh5PtkUSCmlBVYuAu4aMKw
xEEoJh3S3zaBoRl9/Y9elLcQxUybTdELYikj9iIZBBiRxrYqwQdMmDAC9IalBf2X
qXiLpsYBGqsX1Oe3Cz305iQhenMLc0teRkFOgAxiRdnnFZCo5IrVK6/QfFTWn1Ma
SFi55WXb5ztmAvDPB3FkuxxyFJmsFmEPqlVHKGDd0v9ubQoIMdTUWQ0S8n/+Xrfb
O0CntIwm6iIhY6O7LIdF5rT1qwvy+qV9gi3L3g96Dskpyzz7h83FJDXlplNgInYp
4ZoNPRZJ1jq62gybVqScfcBVTUd0KDjcOSO0V/87Q4ocDOTkqGDyr7Z2KNrHhMcv
fgUyB9pIKfHNa81OF4YnAtYVy76POhV4gLCw/tM5bEXBp/q72gxZZcBkBaVDrjZC
mlcbIFl0hNAUkbWfbJnvjMO8gpD1fkSU7waNbbQFyBcty3P0UAMv4+00xmMqU3bK
8U5ogUuZrLWjVKcfuPgp4n+gUOCb4Uxz7eqradqpCJrhinO3lnMw0qh5u98OobVh
twDANfGV8TPOxd/shlEoWVH+xjRinEVtsZGVtvFfA8YgPqx2Kp0U4shonR7Oj7AO
hNvyCN84REr0rUU3AFRtt94NC1Ql/pCoOWD0ZC5K6B6sC6TTpWtTUM3XGVt0y9EE
dfYqlP+7tfexQ01pFeJb044Yf5fzh6HXYRvRfVFVAxaOrQU3qAfRkCjvDyaIxjWd
2gVY6TNkvlYL1iI79eV+cPjVsJCE3gMZShcb/yowiyVe6320tsGosafHqc9b3fS3
AdpM0lhv3Sx0jYduAvP/ybPCYoc0U7Tk4Z8w3X3BkNtZieVJHRmlQgK97eVzV5l+
zOzCWhPwHUEcMmzSdxwS4TmVAplxsP+6rN0BdI+M5ypaVX8rPYCZDh1PvrxMZwAn
JIvCd6YOPhDrJIDq0T8ayzbt+p/uPxqDAkqbM/7ZLA8p3oaNkJHU9KB97pYqeS7L
qv/VwkNoGRbsrMP1u4z0i9NcfcCv6r7iKqqWGhwJ6Ncyk+hwFgDqL/JoqvVvPBwM
BaS1IgsvTG20gvxut7YLbKpJTNg3LxSfoprD6/QErzjJigBsFkTzHM0EYoqbf2/Z
xn9jgYf4oexu3auSdBRGllHMAXuLvaDjl6BeR/VSLPGlZuf49XkTfH42j9ys8bEe
BGav1iYzUPWjpSJVXto4kjnojEVcD0LxTsK+H2fgM2kmqHvPTiYPr1qhEOtGfxEX
DSzHVXzWPOHAyYr6DYsJfnOL+mBQrtHtzoKaGn3svM5f36T6mVCpdSvXpmuYlhz5
/vrcfmI+N7YMCxqry4ozTC/Jb07ApBuazKlKGALRR7Y1L+UZBG+56wxnBfWX79l6
CO6NtZWfZY7oKDw31gWFXh7Ll1F00QMDySSrKSTWD9DXfN13jT0X1PIuHPUk7ixF
iYpEObktRlNgfjbuywA6KwFZKPvdpSwDIkKE4AAkljgds/jU1kefVJLpxdRNlybl
Zux7PgHdVDSVvdlTbQs1kP1A6WKXeg9w5Ez8MVyis0WbHjkKvD/JU1F0gObO7sis
UKjNLp7TRvykK1UOpX5EL1jKnq3v06+SVHvl0uvus3upIvb74NKSZGuOkpqIVzlM
WuyAiYuiwF7eGwkFdRuNfAS4TdjefyZjolWP6zOg3YJ5J+NL3JWxN2tiyUuwyorj
xwstwLvCNSt3t00s7dRq4unRUz7Y+ykgJDyCvZq5RAHROG6YB/Vy0K4BUU88gGU/
UcxsvAimNiHKy1vhK3sXO5OxmCqR9qxFBvnM6hUl1pD488GeTysdjSjeW9zv/FQI
Yaf6+AC5vyKO7qwFS4NLhPR/tMwmC7oKV7NbT0oo4zja61U8OuFbmvv6cjEbU6XX
Kw6IGdVf693J3zYvYe+Mk5rZj14VbF5z/0sKrrvEqVVFkE4AwqBGURjswQdEZbc7
1e3Sq/YzUfzEL0kVSz063ER7CpwB8p93qyjpoWVOAgECMtSFcrdruNbocePPtUIu
rSGZFK4Leg+vmV7//j5UaVu35jSHD091zMNCMCLCBI2OMIKb/a+2lOOkfLN7xUQr
InZAlFr8kS75aKZkgVAn9YrVghL2I5A4Zeo1YGgonKMk6M79mJQZa5mPrDLM8lqr
RS3G3AA9eXqMHvoL8HlhPlzVA3KWmB9weFHFdwsUETus2AVXaj7YQA44U5oGpCm1
41Tp6GRlWEPlb3ZFjVrycQbJcR1HjHCMbvqExVexW1+l3v9yvBcXtoKuLmMmCWTr
uJTJC41CPKdYZzTotVnw6V4fL6UGTPJBoBA8zQUX413S8YsAv+RAaBnYEuEivcBb
pz+41qvB/BdvwraiMURTg7O0zrlyNKsq6+X1PNY2lN/zKTQsF0F5b0KHERcLmcEd
Pr2j5oczP9puFdbiKuUE4xQ/Bs8UcoCihpyUP9QSJVf7+eQRDX6EtkLgKiNg72Wz
1H3oqrv2Ow5ySMa9PUHhZj5lCaidtk3IWlTNU0puHQaPTflFB+pMkEsuqIOo4rwl
7uSjx6fum7XsMByURjoo/QuzhQkrQpDLaKtB/PnFfTmJtPfl5F4zOUi+73sMcivT
2cpbZNe4gsDZxREK9jM1XEujXJtVWnAl/T5lx6m0vKaNP2CCAz5sNrY8u981EBYr
uw5cQFLAp7HfRul3B+VZMNjmc2jg5fAg6jDyGxcdfcJxcLvAeQBcJkdYwFmeIraG
+/GULa+X99CofO8yt0kIx3PtSWFDbmYMIqoK9bL4ah8oyRUmeeN7zPcZQPfbH74g
xtlgXwMqOy0u2fEx3VLXnRfr7p5gQ55WnryKg7z1xdZZoxBobOXFAOQ2+fnvQ1dd
lf49xxxb+vGLx5cV2tOXG2krjryI+G5kyrWS2zRdgb3Yw4YtMhjLEiSeDXZdY+kl
ntOO9Ol0CdQfhr5LGHaTEMm3btHyHdUYuizrrWBHseF4TysbbE4bVW33LkCOoDHk
ANJtmTEOSEP5Mtr5t/fxn7AscbQkS0kvnhnKdl3DsdDl7E2C/DCtc028Uq8aSbxQ
JOjmZKAzihjpKzqJclyi5xCuHXV4MHPLczp9EBubdeQHV3xFGOnDZna8R22XcWeT
uWtr00rpvkSS7DauwIG0daeRy2Y4KnuG3GN6TEF/K+oVLjpjzguxNkawg8d8noy6
gpMxHPe+r2vy4DCCn0wV2G2T5Vmn0WG8N6Ft3wa3quKt93T3/pHIcKczNXE/BXcf
pm81qstlC+LmtlJ6V+56ivAVEouBDV+MPlj75cvd3zv72T3/ciDh+TPya6kKIvUO
2x8odBW07g+TD+dfsZCDeoAGgV0IG/eYrOHZYh/IYT7b+NYwx3qSxRzi14v0XtAS
BB4EVawq767It4j2iHEhAzO4MATGyD/ydaiwmzUp1+btkoxonwf4Ybjqx0H2OzX7
OzLS1zSScwZsQaEvuvPWsMedUg1CMYivQg8oc2B/cka+OA9x7rrvvc0ITVDJalyZ
DMXeyIWwx4H79I/fqDVwxVNwZPet83lL5+qYuE8gbotyI8nSRtQfYcGXF3L/WZV2
pUtBO3KHfsxLjf5CpezQoTDj3wIHyqtX3OtSw0nIiqhyvipBe+dLRSqQX3qRIEpy
L/U6Le1CVsotazWljpCGBqjS5YZcQJaA5D+K8Gw5eioPL7xLZfmTBl+Wcq8XT4C4
0ebBxhqxSmmy6dFvz4qlBwN0gYCmBw4rB9j9Z9Ch9tzZq6TRuQEwsc0yvnGI03dp
yhnSlbvXbowbX9CemKddW4eHUonl+eGzxg6qfnXQ52YMhXT/HqPWLCJSpYIDIuIa
zCmIwOWEaYKsUqkgaIG1A8nABhdcPB1b6WxVhdHGMVjrVxaij3jl4TCRjpxWXvfL
PYDfTbh9eBhtrA/HDr0T99tPc5QGQ7Gl8/ROTDs3ecL2hvMR1Iwa/tIbqHQnjkpP
lm+OcTMi2Ark5FrNjfswcJrfZlxyFXl2JufI7qMQylpbsSs1TR8t2VBGJEH7WO7r
2m0o1HJggM+KfsllSFJtVrjKpME1kCaYqzAEkWVbYW03Uq2JUdArixhZEojDXoW7
04BYK8n0ZtIdmQWOz6mqVreb5O9r4hjNZSpvgTl85qWwQvQ4Q6/sUMluJXS4OJPs
xpxwsDkuMfx/4X5vR7trxAXw1Syg4Ekc56yTAGSlHkE4tpxIUY/C4pd5LTCzUFId
EeO1j2HsBSvbDZdClXtRWo495z4O/ntw6E4ik2JBamhuFrTTEy3sP0gnNqVw759Z
XPD7c0yexwkzdjotEf9/Y+ODltckIo5OSHP7LMhX/2pX6Avarg5shachyC4WEKsD
xaxA5WntWb7g10Cyp3q/+ljRRvuDVtB03cgtlk7n6IT999XNbW4BTiuvCZZJKhAF
3bvuCwLHhvSAzsnaf3FCGLbyIF/YSKBzwG5cXyKyqwpqwFmUO3WXk08efXYSZcnx
eH78R79xDyQUdUNxXCbb6jKf7CUZV61Mj/IC8ogJMhe30Xwlj5HA7J2upc8U+Wp7
ahMT5COqcfjIPAhlIKb6Rho9gVLc/C6TGXB7bRer4WVd2KtIAp2OPJ8LdpmBl+UM
+LJHWGYBY1p2uTaqyxjy0Gj17rvC6HXY9RXzvxwqasNENEiMGw69KCf+G29KEJKQ
IZyAXH+SnUte57DotDEt0cZPK88uJdtMCfl/LcTSCBLm/rHoNsSPQdogyviU9Lh3
V1nP9MQYewU3qK2g9QpPoR1CqYO0MLABJjbV1GsbZx1RBMaS63nHhyib99E/VO7Z
VaeB+rpSJinAyAr17OA2/PAjcBVxz0fdxhrsDZnxaIwTGpw6Rhj14MeNkuVmMswF
LVYGsdOOnUZu2YSrVFF63sJltwGiq3p2Y/M8l86RRYVv/lVGz8juSTqMSbT33Ziv
BtDLqK64Rc80n5Yj27lSlFooz2AMX01+iVI2DjppRD3FqOZGHNak1iN5FZ7FmBcy
RrSs3xwtS/NTo29MUaXg7GFFx1LO9h5PU16cRA2l0Z44eTHkNjbLCEVXnVXHJiwf
Is0L11RrmBYP04oE/3+TPlNhp9Lb9VCnSmb68yrT7EygOny1hNETu17AC/vWpkGv
mMZcyplyCMK8VV3TpqQRr3hnwJLpakRw7uNrtesQBd5gcEpiplgvqQvmkWrX/zrP
g2aqnoKFYCvnQzZRgNYj/RjUdBXKbM5Cg5qUAy010LfopKLgKRvAP24zGwDdz0mw
mlxmwfyKZGyCInJnzuz8vM3F0bJ178hUEjzpn+3I79n/Sx7RfwI1Q9oMxDVLlctf
b+Vl9nzO3HbDrl+aqhKVp9rZxhDHKfN6v+pc0kgQKf3U9KGXdTS+vIzCaMQcRdSC
+1ZjRz77GRNnSjeLLXe1fuffEaHoqBkBzQ2XetA2euPCg+dai2ra1Ln4dV5uYHfO
14d65HYu+5Ix8xginh+iIsvsrkeyf2tJ/d4DwnLWjQV32UZ8FR7338wDtchytVQi
R+AsiGFxX23hrniK0hmozSdmFgVAiZ5a/TDvkdHPus7yyOPmwPy2cWdM281FJyPz
ddofxupJSA3x6w7EnAvn9XlR7OvU44xJVTTq44axwb1y4iyhjsXL3c9DHGe8G3rU
hcOoTx4qKCAZJQiW1B+24PTmmBCYHOFgqj1q0M8+T4It4WDn2qRXR0GN+9cPGn/B
zHDiCC09Qu72e4tya8396HdGJC9tozFvsmNPNAgd2HBpaKRAVqz3Edn1DT6zM4ec
xx9Wn7/tffL2gumSKCYfMy3lelSHALrwC2VqW5ZdWjEgikLsuCA/UoOnLWi5qxGk
SYzUqgD99DSVoATCj6fZo2gz/h4ZuAs+GtPTg2xW2rn81Elkz+AoHn8w33hAqnNx
XNSksPJOPib0vEWAQ8kA00G9mrAhJJ9cif6jDcxh2+Psgg2xfj853ED9O4CzSZdH
KWUDqmIHOkkdy0bh3ux/H9X7yx0HpfmLA/FB7AG+YZv3EIBxs1JIclkVu10az8iX
A0RPpNF4A4kueS0fyuRJIQbOrTr6FPsnhyxNS8CwrPn9dx/E5BGgI7lMACrMXXXq
JX0HIz7TvdGJtkn8kzRQhuTEJbLqOOIehMDHoJvlf9KupZSCH2IWt5qndVjLR++L
/hE01813YwnU34MdnLVVgPz5Yll2o1MvXrnhUR3o9ux8K7S6W83w8KjzcAWqBY0E
BQKvPVkxUeCVujt1342RVGg6CwX4oCTyGPIN6hlbBNLr3zkGbcy8rmsjD1fXRFhu
/comKkzRqzYK992NUeSrXdggK4ExiJ30iEwp40XBNsT4hALxGsdtitRQnzopVn24
wQwgAOsC6RSDI5S36J2xuR8T73ncAKbmXWdoG6DApX48ZK89nb/3oyGYsDoaNsWf
2mu1jkIm94QMLl74TeEVzLvZ877oQFjkw+AjdfvypUOVbYCnleE1lexIRxlrrPuI
gM9DADYQnWyM+yPrH50oKdYns1I/ceeJ1/ZxnnPgBEw8xS+0F9jdCK+ID5A90UuR
RpMpbHq+mCb7EdE0O/qFsu7dOHGivaRpWqTXPtxCDr2+vQVZmipwFov+G8MU9QIp
0kERUNVlSAW8uiZ71WOWIqth6jkHW4qCTa96bReq5c7t+Vs0oj3aXIXzEgjl3o1o
rzlp9mq/b59jKhSYMWgOBveptG+5KdoJZTi0TgruqAGG7fQ4VH7GEQdx/Rb8+GW5
Z/GJTTKEEjYUOkyDD3AM9n2Zji70vh3dEg2mLTgHGNNxu3EqTSDWL1jadU4R/WhC
ff+Dy+elpfuLryPiVnX4skjRzk/t4Lebmk1omN+621/qWhBAzHBRTuka0UzxvCOC
zkajNKU1bVLu36o1nk6VmCxTm2+SLNugELyBzQoWDNjtRkXo8I4Hjk7OJwDhCPTg
d/x/G0Q20AGovnG5N1mqx/cFNPBtXKdJyggJinnk4UEigU3R/AGCPLzFlpGxoU2v
Gc6xFRxHZLWwv4u35ao+0bAwOb0sKDyWvm0+e6IZZHhTHcdIGwS7hQ83pwDLR6cR
NQzSZxogF3HLXvfnZJcxXn2stw1SjrumghTuEiNimhXk+qC9JIPtaugY/6QEDLeV
XJ0qy8ORCykTU9zAxzTaEohDFx06TI7YxS55zkTMH1iU46SBh6vImKugQ1hxwY7P
sfuHYZXhQHGUqPpZ1xsmAEY9XVjjwbb/r8mfu4fYC8osnJGNn/GHKQJEQS5tjb0+
96HXPtzEOVC8isC0NUJxsTd7gFDCdOBeQ67cH9+2gPDQh1zvOnkeh12x9o2mYLNo
+/bqD+NInFPU/ucjSbHDClP97uiqJZ3k344p+mYSxBt+27ADAZ9UwF4sQHRMNtME
OHmZnctY0YoFMl3o4+0zYX0LTk4z2W0/PN6mtVc6VPKm4Xr6QqsTvh+KyoiQp9X/
vKfpS/ScwRC0IQClJQwNvr5j2ykcBpNnYMniq07t54Zq+3EbmARY0U8zaLFmHrNF
yqN1sAm68GEmgXp6fnHPTaGCYY+kQ2biCIc0ogMXCeGOZJmurxn++SdylmhJdqjv
UzTCz/mPpVPzXg0pnC9VU881X8i4m6/vhUQgJd1LYhIW/Ph7Kv8XB7GPJIcL6BBP
a/6GaUPNqAqOPqMfysg/s4B5+cYAj8s50eeQMMZz6iOv5GZbVPWub1lVuWZH5DQ7
G9FEnazo+ru9j4axGcSbZ4iXl9UtrAm6c4fDAltVT23gTk3GBTXtkdojMXG71a6q
Jz0TMFMVmQLIs/qgAkjPsw94GdY+XDBTf+xB84DalockYzRY3BT/zomQE1rH6sND
E05TseZcIy4jqvmnuomh/3I6prnPAu361a9Dd8LlRvS51YWVKX4TpSLqLY11LDw+
Nm8TexBipMfOReNLrYQji6DCUxB5zv4BeAX7lWb4/oiKhelKNkAD/QHJb98G1ENy
tMJZLvnTj+aoyQs6MoFcoL3ZFPdm77oO6mB/ghGz6CnP8znHfJ0OhX7uw1fb88uz
hZdVRkUPf0gTkfZ5JqSVs/OxTigfUOHRN+T7EF46l6+1V+RjYhBmPLKH0mjdgd88
tqO7N7pnDfVIlk4X/woatY6nkmlWUMCX9NK2wLHvvfTyLQSFKi4uPp9OO24Pp8g9
UvlZyx/3AUlP1Z2J5ZxrfmfYwIEp6p/+Nt6wrokvo4oppbmE3avo4bQ6ONbXCpP1
32LhGHxq1FuqHGd7rHH/h2PqZQbGQ0vxs7l9aM1TBihhr8/C1yLH2Of7DQCH/j36
FkWU3e4B1tPAt9Vxd8nwuAM/VzTxUIY5aY3v7DiGO+0ubK60DX0wpGUvoDR/7gze
tbDVkKudFX+bFVGByPOnWaz+6xpBwB0vl8kr8X6UB9xV198AXdBvVB4AeRIWDIC1
I+IAGVBd4O3YmNfuimHXgRcOMqnuvIB9CaTDcySaA2DdoKd4EZiJCqVRKIpSGYF8
OUS6EjnPQSSbX2hjoYdJx8gc+qK2N5EPcWbC4xzT4aR8tGNSuUNEQIa7sYSZj8n2
/03+E0CY1ny5rTgXYxvSRj6O5jaOjjcsTtO1gU70TuP4CbONDXpWObxrjDdXMDIU
bLbN/IoHD4DVbF4WexP0OMMzJ6SyCGfCfc0O2zFkatyaj6CVkQ9gEm9PKq044df4
sADJzpXK+OOPdeLhChpiP0ZtMQrejt00cLBpAsi1mW1p9t4kDQYRQdzH1Q8d6V1l
unM9F2GRDz0+XVHDjrShwQtdjPuxPUrrIFngnhLVynxM/SJSr83SOZDffZiBn+94
yn9rIjKuZlAu0f2AMtpxW9DwwJ4HaaFdSxGZ3C4+C0dV5+94AqwsN//niH5GXML2
EcvPfMyIsGYf4HEk+0So3r1ikKqrEKM0xBvAbSXUuBhwaa91JRGEa8AKiITWEB5H
jlNBCPKs2FB+S+q89kVKj41M7ljiYzTajJ80nPYaDCfLDAcbGqonS2xQCAjbO0IA
GjfISHh0ENoB0qbAaZGB9wAQO+U9dQKuCIk0+PclIPws833GZtxXw2AJojIXY8kM
lDEaPdHLMBjOv4LxtV6vSp21bkHXYJOY6ykpYPK6aqz+IOh1evWWfACnk8sAgCkI
lfpFz4OL3pzp1sWLMHAY+DgT9NBS480B7j4KCsTUkz5GwjjK+z/cSmmq8dCcowqT
KgBuzAAgsg1yl/dyABbd8vmbTIayj2yRe2jFhD16vEx3UhsUpdsmHDZVgJQoWZ0T
tHPr5yAp0dImFfn4LkgidB+C2H8t6RZdtjKHbjqgtRRh54Cwfhj2Wa+88YLdrGNz
glsbfpYpM1q7wEySqn4fNujrNWQ9AOXoveREgKzbWMNi/zmz1cpytjNwJcUhPXWQ
+0qkPqXlIYqPJIYOgfbsBd31OXaY8d+WgpEITXmzP6i8C5RgcMkJz4/vLvZq+z4R
WDA4OD6RhD8SnXJ4tJ4F92Mz63bEACD3KbxRGRuUIA7BimgmRiih0uXxRLcnpYYd
BAQ2FuhesWqmnEh/LZRviMSRRJyQVkfV2fErIH0ss4M/Q/cfibvvhro/3e8OST+w
iaJfnFyg5ZPS4Sce4xnrAXSCsPJ4YEc0VsEW8mDTDh503pUckEplLrXewFqRzuQr
S0CEk/uMBxqVTfomK1SHQgEqbwVqT5zS5TZuwbXWNaKQ6f2g1aiC/6WiZxsz+siJ
sxi82rMPjuX7PbmKnVI0c687jwSHCJ3CrcCVXphKzYXNVULl2jZaINYNpQIYacCJ
6LYypz0IQO0f1TrLNXobnbCwdn3KLYW/bMheAD9TwdiJ9f6MnVtN7hB5J9ImDueB
/fgfdaMVulqLkSbfaVTzxiJFXVIRQAFyiyaxY4xZDkAHUesDzdgMJltmpfYmchlg
EHyLxZyBZ/3t68afscdb9S/y/qGePuNh+kIM7ag3zPJtgSKQ3UdlH6by5Rk7AnxE
gqUtRynSB3GeJ6Y4CziJXiSrdRwCc3NXGKC5TxI2DG0jFjCrEvARbdNnXuHJxz0Q
qa8qXJl2j5P0Z3EkROxiE2EVsitePEqemafFjQ/cezFXNAYpkYHnvdncs6sqhDnx
RWg134DNdLUdB/Aznkj8uCoaBL9nrmk12tA+84MtN6doG9tATydH8H4ZcCyye/1o
8mD2LDMprDk6trK9knss6iHbAITT66CLg8wpvT6AkR8k6oCAjQkLmSvi9V/Q2eUh
NtDw6EhmJa7zm5dyyQgbRxBc3jwTJgBWqRCwmppg9vNN2R7WUhQ29gUfCGJx2hCl
J40J6IrrGRnWPZjA8Jh1Cx2/xPEFybtyj/fybP+KOtIM5J6uYbJUguppJVJtV/AI
f6iEkTxPUwSv+f5ofSYXxrESIIPMbr8/Za2aBmtfISx4LBUcDUwKaVwPSLYWNJ4C
2FK87WVeCdWO5wNDEzvnS85LSvg1vQP9ko3fkiORnWkg+OriTA1zvVcTh6rGx4Ry
P9ZEtJ4eAQPHsYTOWS4oQZ4EqlKLJb5Jw3OnR1ht3dPyRS54tgMgRqiZYwx8Qyfq
TVtqNlADHObFJOB1VNwLJmnWggsyLnDcFObZZPN6gbJjRvaoNfhhxlpQebZkEXls
aFPfVl5Y+JWcw8PunCj9rGjj/sLMYrkzn5B2qLao3wVIeUBWBUYLxmbMir/P2Y/y
hJUCojfjVsy7nqP0Ztzhuel9aCOvXqAy7+XlYk/VdMxdINz3FBooKDJswuFK4tP+
Y4WRt/s6dStVtIr6dAdG/q1bEEGVar8y/TcaxNXa4IGf1qg2taSyjJOGvNEkT8YE
mU661WqlCU4K+hQrzI6KmLNVhNqcnRfZZsEPFfqzr2brvc/1NuJQ22qLnV3ijqD0
EO96tfckZM9UhKuEIrX/JZJrErOhYRGNud+zZLhZ/s1AIFqBZFwpL+VzOB8RHq+0
bTVV2Zqz4MO8onFnx90/OCOZOUt6sc8ycBvJOiRCsYI6bUVvYpX+Y1qi/GXmqq55
wHLGaePHHDs6rj6dKdm6J55WKeuAhtZ5H7XNRqmWqFPhL/dyeS07XkLZcUMoS1bT
XVSgiaoj+z/VWpkXRJGuUS5FKI4hpYBPwS6esPdPWdi7xWUYobiZmay4OoDkWalm
2Am1dt+iuK2WF7J4CkPZCEkYi1WhkrjOFAeVSeeGVZUfjsCU2+rvWMj2EyN5XABA
WdMEeUmV5eIYfxMzWk7vstNyiwxixjGzO8M/7kYPlngM8M6nCKLwogcU4LxbdAKQ
muCCAAvNPHWGS9Skwhp2+wsMxzJooEj8ESE87+90rJbskMLDC2h0bd8NFHGnzJTF
G2bTHii8KWiT28/4Sg89Gp7CIj9JHfGNcs41f46AdkhDVN0J7twckbSNXmiPsqe8
xctPdGPAi5zefu/S5hvUV3wHw79l44jIqYjgUV7w/Rd1npRF6XBdeGDDmDvReZDV
DW2mbeh4SnAFmZRs7QaPuSl/+9VzWygonVCP+uSIl5qMTWfKw/ZMpeF95fUppNRj
eVKzeMiNpCBH7MTECn/09PSOQ64pppNJDqWqzYKt4yqmUWD8uQIExrFfODk0GOrz
4mGk16IczhPXTJMvgEui7/3P06kMzLu8V/zYnUbVQgpoqfgOzcVQAoMhgkbxXhdF
3EQpYKgPScscJQXdY4Wbs9wD/LRJO/TOdQpKCFx4N1fmSAMHIzKM8gULVPqTcYQr
08zQ4TzxwdvpIZhayoIlHHFlb+3wtZzM9xQ8R4tcIZ3qaAHut50+eBJrD00mljHR
43AivllILCOeIoFUvTVhsaWUHmx76N62lGxlxlIlcbCFfWwTIRAN7UsLo8csZrF8
NZLPhetnlLgwvDmrhaGsrOD19b+NPyIYCe14mR5zK3BHJvqmwW1w9FZ5s6bENM63
H39wU/x3Jn9YSF4ZUJW9V8tGN+BeNF9gZpwpN6aI0b+GzTG4Se0OJI5Gz5xtg25v
SZ2VBimv0AZfALOdJW/jM78CN9tRpJEJupw/kWiqLLgcRX1so4wsbP/+Yb1O1GHF
URwimkCadsK9PSoUs1irejteLpD7UdmUuD4+BIPiL5PXd/9U7frKupZKfCq4qu8u
SVXKT4pzzIB0Z7fYswanracjABB6aP8VnVGTJkpQSx++5KncvIHRzmIIqJTf4p7F
xZmW/EB4IEyw6/vuFDR/DhNyYAiT5Afa7A+qc8cUFm1ofeLXAIeWevzeStRJroOA
OiUYAuHtbdzYuFQY6ovgmtxykI+ryjCp7Za/WG4tEgYgNBEJkpPYVHO/k1sDfjj5
VVeVvwvqXjho2kZJPa8UHRHpAtsxuQXCJv/4s4zSpGzX/D5yDjJd110Q4bsF9NAX
6s00syAE2UFreEdSEgVMeKyCM8nTLkonOO5VFcPxvMwUWw6ywYviMUAjkTPlF0uH
fSC7Gkr+A6CUoEtNtPY3C/2Lnk1/CRgrvyKYMgCUYVmyLpNzL59d3N0/4kQcOfCL
MbwheYb5tGaG4gHcBqBpgzuJXDbeVMMeQXdRGPoBF/XLVZEP1AW2ccOROVzJ5AnI
DlOlI04QVGIVqsUgugiel3MuAvBoytCZHGkrsBVmKWuB29oD8EAh9IIYKLb8ZRpp
9u0nlxuszYbGiySpGybODes2YIlIox4daBjgmkSo+0o74euBUOstmJ19unwvdNHE
UR8UPHGWAF0LtiouA+KWCVvUCUJa1TNOVYEG1IROSuBOA7smKJlZNwCkbwQjndZ7
gNThsha0k4yGzp2JHeen/JBKwQW+BijoE0nhN6fojLOogbfJGu+nYv+VrToQB3H1
vPo+vJV+ZRtfEHowrj5j3t0ukA3YPRrW2UiFGXNRaZj9HA9026cDJMPDVQkP020t
wXxIx+mRrEJp1vLAaTRqZLF85sVURoHl8kage8zF2j7vgJpitd5FpGLvxp6HqoIH
p2XdKsaC1FIuFtYc7fktmM4CJNbEZXuiXFgv4ObJ4vwqVQXB7DkW/0LMHxh6lK+g
5jXZmwy03QGxOQC7QxJJr1dY5AqDAtvGvsnS/2zcVzCgYQLZajAOXHTDHA2ZtIih
dgt7bU4nH/UKpV8RgZTOGJ20FkQZ4ha14wG1nWvCB2nbplh7RddpgT5vcnlLvuj4
bwzfMMjBImLwNJPLO8AxRYI2o2qRwD0+eZ/OfLp856TPp2dpep0BaxhJuK9UP7SQ
hwTRGcIb5tGHWg63CkwEs4X53srZR/dFpwljaj+V9a9/DAIa1l+T9t7Uq8OjzazS
4qe4sjaU65LefQgHXjjw6QEkM/oSRSURuWbWVkai76OG5LaGPCmlRKWvyMBnICHQ
xNIgvLZ6OtYRxpJbigIKV+6UhXH4BqS4EvV1Q5giqCum3/JVgBY3doczGgdx49zD
k+RD0tash0AG39KrIGzUP5eoVgUQxRZkVpZcRJSG9XJm+uP3PjCgrlriJqhKKNKN
lPA9S9HHmg8zmZYpdEP8Ov2R63cuxUGrqXvAWaW9S/YFTjD2GjPPdxCx20rz9yY1
KFGoXO0nWfw6trYSp/njLUr7meaGNZ8fSBZqPZ7xG43kAzd+khp/dLrnqlDHzFnf
cMo4GNzh9XQS27+o/QXY444YCU6oeOzKVVy1l0ojfa/E5w/4uEmz7aNWBuhDB2nn
UP9gnCZY15c8CDOrEqe3EHbSG65PtHLuuKrMkjWGiDgtOv4tAEiNiUGx3AX1HTRQ
bf4kp6h3afZC+N7GpfvjSrJVlgCorWFPx6J4Yelp9Gr4xPgdxYLY5DDPMrN54n9S
Mfgz5d5H45RtKBo5SsO5PhlI321aHUZNFnt3jVTrWLhk3q8JGetWpmVydNBW/qXy
7dgkzfryVKfIUBrIgx4gt1+mJTcRI5Joq3+aGGEZU9CbC+C4VEJw0pOaod3hgkUH
Im5hzD1bXmILPKjomE8FaQaTIDCSCTsmxVFiZlH/9PNohVUZMBJgxTycWXlhlxcx
VdgR5EIdKrnZOCN85FNn7qX5zYogTJ7G4x28utPH+zq430yrvPlb1rVBCndYhSha
cWEnrBwL2+i/koSvOaFNdQj7uKXMs1fi7LuDuU2czsZbd6qv3vpMgDJNQGNCf5xy
HFOiqsT28N/HkEaI+16xUcqfF+7KjVO9H8pJqsf0rBLlP+uCzmp5zV1jtiLdbgdS
1pOmZlmakpPsoWaM4/OEP9iqaCwwNCngEiZGOZYgabSGmD8AEF6qMYmpigcVW0DI
aYwS7aRV23V/KAw+WDYaptEwNlcRaFDtd/mF7TRrNYMoThDlNU1oUWwf0hhrNFtL
7go2fFKErB1Hctp67Bii6ICAfvAs7AVr3eccyKNXdsjv4nDI3N0RsBTMusDC+mo6
TPPUZlsZbJ1v4P0wVUa7P+PHMwe+TImDLDXyphFe84DY5W0PHN/Hr2E8F0AHYLrh
s9EsPFojpXXmA9K1WVL/l/6glMpx5kg4LD0KurPDo6LQrYD5PqXdr9OZ7+Y0Wzaq
94MlMt3ccs0aXMsHGM7Qjvca6TU0ztui4OieCf2ys2/gVniQW8C8K3I0XpbxNSI/
l6fcXDOjdg0hRlNbT66eC/dF0oSzSsop44IWaAF+S7j0HolWllP9mkdf986ZdPvV
uPcw5FXvZAJMOeveP6De+elyW7GO2COpDnBFUdKzPKugQOM/ZkjGdkm8AsH1xkz/
MhXZWH/6HFZEjMJ3RPSzRFPVtjvqJbAENUnxj+s3REojcg5mcG3CvQ7jx+xj/quN
3acc4OG/8rCcvLwbjs8X8QPsftjMb8j/pY34YmL/VEetV0yJzYZk0ErhN4okENug
XihxDMV2R5lNoTTIm2IQ0tHmtyTbj0O0V/DyOg/igytksNKl8H0eyiAljJFKqEeH
tpCARf4yX5ZyUV5IGMWSYAROTbnFyDkbjdkUqp4f2StL2v3vnebBJjNGxoddBnYk
4vdXwediGhu8TWxYjQ0JJtTl7KMDcRvL9PYPZP+bIKU7FRGAQasJWuLyF0XFjAFy
JEIFJt0nxypQ2FNaWNnBNS8Dmujm4OD/FujVBP6kDAYPDVaPR2msi5fzV/fhDeAF
BxpoV0VQzNXxE2a4MumfmEcl5xNYLaMPdiIBcOrwl3BN/KUuMeIf90G3oGH0t/Uq
18xgPI9Ganv01i9gNNL+5LLmL0wCydLmWZIgrxG74itBfH2AWt/IRlVRAlxXU2zb
/x5Xy1AxnLy4gZsfKgDcnpqzM8VzNxanLmevMw+YGmDoVBPk6+E3FKP2jo5+ZffG
eW3vZxEABn/DbQzhs8euMVeBwgHXdSRSbW9SKdMK47bvJrmuMw2unUB7h2Rh4kjl
pW1BSzmAFh+jxv/gMY5b37H4V6E5JszUf/ZTDbDU/Va0nvGSR07szpmDmY0vJQas
9PnS4KeKFypdjw1ysAn0X3uUhxXJ6hRSXGw8dt8Nf7DPFvub/7z5RBU2p9qQhCDY
ZWVwX3gYWzYkUBrIFH8Qmy+77pWCFcSHPzUH+O0xeKNfMjiRmhDKF4uBtz02+9D9
weQOAErVhF2DdOpGtsBkTxbDvNe79NJzTyeASOMTMtZi+J0D2X+jm1C7B+N8UVX7
UGiNiFnVYlACqFcb/O2Sr7ZuI5GfYjj3MLtvM3ejrSjof9vEZHLTTcnG/Dxj2lPG
5cTMChpVW4rbUqP9bspkKA8Np+EmWAolojn4YgbxTHZCnoAiE+CvLWAsrRa2AiM0
c1uMujPj7c6JnI8JsTU9HPEo9nXpW0fB9yCDVL/3K9crT8SAftlIXKx61TPIqCvC
kAq9YNSnNa4r2t/6t+JQY2R33t4Wgk2D0e3y0ROsdT6k1XModCxLbw5YlUNFQV9n
SN2BlXqTY9d5EGSpLCxLXFDAKgqvKa6Cr0QCXUnRxeYBXfbjjAg/eLriPGblgui8
GvmQhzNnmQxCfw9dQF3KLQyoNVALj3SOs3H8loOS9it1Vwy4VZkjSURUUlsNJJU0
JEB4XvirEVv2F8EJX+ColBuexFHrcU2Jm+BZBpF6iFcFf3u+buDzUwZq0bzRrPnq
IOT2DSaNMogzu1A00RG6FPXlI3O3Ax7TbmNNabGpqPgQ2Rdb9GLdX06B3566hQVO
cCuoDvc6NyN1SxEEzrNT/R5wfSy01TxwHNxQC9HQpZvqQpCVTiijQPg6m0leTgMY
ASoKfzf7/1uDxaSs0Y4T9qcQMUwZ8NmRtSDqerl0xj/KO+XjppQCYzZwUxF/Tk99
+/MCEas2ify2drZcxEYmbD2cx4AsPveJ6t2Pxv68Mle0n4lHGfZuw66v409o/2Wr
kduFW5J3armyZHYr4n60rl2CFPP5S8x4vhwYn9Al2xO4NHPIngCww3iFnpf5XXpR
Z94XuCFrFn7YZrOjTwSBRKKjOMk+raq9Y5gYLRfqnj6oH872j6s9vt2VaxHh8/Wm
9xTKaYaP27iy6mt+4aussUhnWePlzTytgMvFcTTSSszS0hBS4ZfAgqILBQpmZ7Tu
GMnPRk8oVq2WHkhJfRyp3Z9B94t2yCW7Nhu45fvdyLOUbMGvl/uRDgLtur17KUO8
kkX6MqTYxW7BUH8Wff++pDvENCxP5JssfyJRKUC3BUFYzOB2VnYHDCJ6k1B8k6Yl
bQ9kMMzxThp2Et44yP1Nnk45PPFYbV5h8GS2+R0qYfNilv/l51a6J7sd2Sqrb9qh
+5Jvk1kSPlslKHqjH8HeMs8YplrVCgOlEaka+rshf1YT/ySUNPYCUt5hnEICx7j8
UO8lPrAxy0v/Go6aI5uoyakeAHmFxzRjfKhZNQmhqUOlXEwazWfsjoQG4fHcr6PC
G4xNq95YK2c5bbcBoYqfBgZBwtVsOKzTtADxY6qnm/1zm2B79N09jUbBTlB7CZPd
rrMiiBegPYCcq8zMm8ybGw1K01dUacrvaUtJBl4CGLSe1dFBIbRVI7sx1USJodMK
xORUSuGLWHj9jplke5eK6JBZjtt0LOSwG+raGgCsoecjl+RCaYflfwqCzIznXI7I
7QbTvT5aEuSPJGA9DjZqN4riDnhB4fzuuxIptlkpinfW1sug4MWmuXBeEUdgUdzL
Vb/mTGA20z9nsChMh+uIOgbhzO3ubMYzOWweotMEz/t1bO6L/OF/o2vjCPQFhsRq
uyPErPZFJ+WhrOV+6ZRLJsDusn8ZoEnFhbbrE0/0iifAgDCE7r8l7jEDcTxvPfxn
dtlMr3EVmiooNkGehfmWqKLRxZQVyPi6CPDrsJ3W1Iv13bqYFFWjrWrEKBaRvdQN
yBAd1aTVEdfljADEUPBDD+eVRVNnB0lQVyVaW22+Yy1hopqk1B93+qboFSwObRZT
MXVJPVaJ67czeg8LOSd4i0d+8Tt+Eyd1XjerPpt7DZg19a+gBEywrcA6bC4SNjg4
kUgiouCqYQMWf4IdpgK7ahqOywD7tB29sz1I54I8B8ZVGaclGAeW/SFeVcXdfynU
2ToV9QZj3CboXAbXabQ5PKdEe+GeupU1ADMsqOSOEiJ9zjcfUzGSda2xwAs2ptOl
fZn68Ep3OSayQYNAV+j98cacfA8S2wxOkF55NJu1RKpBulrn77SzU2Rj2vPwI6s0
f2QSN9T7kRQKQI3dPNvr3CaoYsYQ1a0z69CqTIG44xN7NRZlExvpkjm6lzjuX0rz
9+ZTXJKdgHmOfmOJH9EM3HrC5hO+K5JfSZUlejmBSdDHK6K2+vbkCOM+OTNh4q9D
Mqy2D/t2hY2GhNCo7p8q0ehotVxtPMeyjNtOFbAwOt2RPbuSMVnM4TEzE572tvV/
NSktgm2247fV6GMMWO4FSjV7HDA4wDBGOf5I2hJxOV+gIChJUuaVooNE+Pvfh5ei
6xu7YRcsP0HRSu+eQOJOw3SUSoXiuTYWR4dBrK4GqMGthDdM4zXSRKWmSRB8EY/M
IRsQXXBFLQkxGyZ5PDGaN2jCzpe18FzvO3zKTkQxJLG9jj3bCQvIcugXlvNNSIcd
KKYfBBnjdlzuNh8aMIpbXNih0soWpx5Yar/WK/oAJrG4m2DVPhAA6IncHffBd9DS
UXcda7sbxDX+/UyPfrn+IoHSgKsIwpdgjtK24nat7YyLDSm4UWMcYrnMs6PWgJyt
YA1NbQIPsM66iTGZlTDKcKeX8p+AY9mTuXhYgfEQqZqqmY5VmzlyRo6a6+Q2c/q0
1KxhNMbwVZuMc4PyblQoPTkBGpWxED4zEkSvgy/U5suEREtRrwPl1tt3qnfZCwED
S1SvUef+y7DoLTfdEjU+dfYfh2NK2EwTFanG87zwLaEZLC3GLBvMLYmn04Gy0kVw
tDBTJtg2nnO9W7uf4J74aybPwWr9M+HO02FZq1TiUFm5qwd4IVCf/oaOEo3fxl7A
xsAu/1UVdOBcb2dsbi7lGQe6ynKvkTigNCNdFBqDPhzqN/gvnqlNWosf+iTrIVdp
131FEQh0s0AhWeFoLEGIKijfggkNwf9sG6tgjo+sV0EEQd3thec9+yvLNXk9GpjH
u+hSgcHVMwb9CkkbRmys0sn8wvUFjSaMLvjaTvU/SU7X9rlp2Q6c4Lo9QnxS/bO4
O73zrHQgZCME+7QMwVALj9dqbGJM1VZJ9+pUObiW4+03xOdtK/RKHiE4T3kHWfhm
JfMkKYxTaZ9E4rbHL+5c1VSD0UitQZoe/80UTs4N+kJEq5hC6Ve96F9BpdhpZr+U
YK1X2ROw1RGUsAth4FDO5i7INvD4+MWO3fwt3QSx0G5koaXvVuSuaaemwYJ85MFZ
JmV3bjb4QC8aAl9Uw7qAk4QCKEwb/t7+gPYFzAswxVn3oB5xZryzH1LMWzl/9G1T
aS08RhbHfZ2L4o+F0XOg1SfTh8Jder99O6/gjP7JHfXz7XCT4jzyxY+CVfKnoc0k
rLL37Tww5TMU/uO3LbMphLvGQSKB/7ZdrhABWHFVWQ+ycK+lqTOxGUGyJBwAz9pY
/COi2MedMjeX/wvEI/YT5QsFwGyQTKHLs2daE/kGMvPYHrraUHFTnVtqr/t1V0Hn
VuGXOwBfl6g5BzLV5dk33Ie9BcDxqIQNigg88CIPL8xvuPN/2B9VBiOrRvDHk+t/
r3KKHni5i4tFoiKmLo30eLh8C7yLpMEJyxGcgPg6shL+Zg/3+tqqoOKbnrUCIteL
tyqklDcH1y5S516EgYUylSVD6WzA74fAqP9S0qbaVcTHoxqD8aAmgS6+v3CqCg89
jwoEtZGIQB+Xv6f/18wfPO93FxW2or8kVe7oQH9tDFf0stZza78fot7cL+IbcLCJ
o5EZjcYsJUY3uuNqU6TwTnnFp2Xn+2HbrLOFB5vkVW+CqQ2uv7AOn/zpNimSNAXd
W7mun5nHbhfIRgAMDvY+fxYasFsS5uBKnANFQQiU6zi8USRTlcsHwUs1WnwjdMir
MDKO6jnRZb7TB7dtSKV6otSGtTbPuS1koCdVG+S3hFQS9ffK9dJXqiheS9wuZgUr
dwI0rnLfDj97U6CGLTPVGXsSJx2DlXFpykT+8/7iWJ5AHUoSv4Vbp+mDh+iCrcqb
khbzXuOxYzmT5JTamTL8EowpAoTm8nq2aSgQwddSbZ2cqCCbrIh0vDkviCpfrF3+
RZy+JYvEXz6Qbef1W+Q8y9fLX5qb7DeX50kG6lQyLimnR8hT2ddoJqDRCC0duJZj
lOm9sA0vje6LkC4TYxV6G2aja1bxluSajkPYMPgy5VBs0COVVpmYCF3h6KRa83hv
lNwSkSHqBomE2ODI6ZECpQLIMpwMF7Objd3RHZaAGEk6VT2oPR0pZjKBfMRjSsZM
wds2ZCyadGXKU9dPfOqXHV+IHtRyYOxA7Q+HakYrRdhZEo1MrBH6r9h/uS3L8tQ9
oHtVHJr3dti4hZsEhKjDrBh746D5yjce0xCJDXiM9IOrApI7UfPwKGJSAOlbXnyE
jLfauVCGKPtLit/xWd8WCbwzQMVNi4m1U0QP0Z6s6GpRbu+dEaRLMmf6lp3l67+1
npMgQcjjxyKgHDzwmNS35iIPDP+934STOkVocZ/gSIrFXeYQa+Q5TbFLSeQJ06V9
wgBwgzWp8XrpTUGet149Shl4w1uutbrKRK1BSlzVlG3Bg2cM00knP+kVwahduKyQ
GMCcacuNbF6ytMeRjSqaImfxOWsPhnFD63eBtd4D3AXfRpxEk+2WrgTNVdmZNpjs
+ZGfcqvvgbi+Ux5tYfPK6mgA94SV7T5Sp3sZz6AuuCrbJYJ8UddDeKmREc4RE6jw
civKX5NtF+Vj9L//GryEkNExUBkcXQNyez9/Qx3Ow5mE0Fi2Z0BP0QkRnYQsMARV
/vW44WCD09dqAZqW6pJIJF1LoJzh0lDM36qvhgIB6bstsRJKhc3attg8G0PnFD1y
Lywq7mbt5kPt17z371jCWday1oDrfvDMM6FBN3vvj/Da/xDxLCl/CG9oL52kB87y
dqEOCK9SQ9NdJWu84W8NKekiK0+uhn4vNAaKGVl5ABgzkD/25GcZR1wAHGuGQM0y
wSPcdT7XOooofFMQKBrBjn6IFQiRl/Nd9nFLyJjTkP7vFXKg9i7aslHo+GX2Rcd2
E5Q1CX5sE5SUAp9YAgVFSUgcZcIM5ftzT6DLHQtBJ4NlCTRIym3+SmYiKVp90Ojz
992EoRTN8s0K7lOsFjcQtHCUSrK0SJtbbtWLtJdUylqdc2kvxyCHCl6e90WTLBoj
UAC4VSqjCnCWHw/X6e9b5x9XQUfu/f+m1kTGGaeFmCRj4dfds3p/E3TUibkz/0Jj
ILfbPpJEyaOLRwc54LRaNGvDZg9WAa/6KnEHZH9NMOqIvV8LXLlecve1QPwzjj6v
yKmDtaguvk7c5Ymnx51GsNhQ/IY6QUKhgji4cKZNwvNJlV8torzevcVfnAgUK/R2
i1E6ivt8p1Zs3cN8qgszCVfvVvXV0QVWGUY62UlfZTANoJXlv2qU3i5+RVjAF/gi
G4bOlzLMu4hvgrIUvfWSaDxODwBzRdQVlMxo/UKmVOa7U5yT9fxAu+i7THTJmt+D
beWFDqRHTzWCyCwUTx+fcJoT6pikkiHKNJcBHyPVpjwhLaJFknyw0CzMPyU/sPUd
J6y8iHLOS8kmQxTdCAt5q3ovGE4mQGXqRbdJ5bX5XYSlrM7iOL45cWFhaYx6OXAH
QmUNfawGfiqy7rYdaAfMjawkMbAPeDO9hk/3Myzj10oQ85DCDC93AWJZr13F7KiE
m/Ry7Nqr8A+UUbECJVcQFvTx1hPB9phgQVMw2MiQ/SBNBwVS0HIrFNCbLL9DvL/E
Rq0o/0wJOI5wN6ahsTRWhkwIALoeISU2SkJdhS84jAjBn4AHmyOhNlT+rCpoUPNQ
slu+N+s7fdwdso8M/jtnWl/WV6SZqqfJarMqwAxXq0abuyEXVsn10+og09MTUa2P
2V8S76oE5V6EVO9nQ57ObJu6M8hUAZ11NuLI7UWta0KSAtjFRTv84HSRfPgeQoVi
uVzsypLOwV7hU6/3RQqWOwyzinx+eESz2yyqNFPAVQ5JJgHKlWbPllVcRdB4IpDN
aoje+bhtoWh1v7kaQgq8WpbNh8O66lPEp65HLKalSChNzHyrpfGkDu4UIJtc3xMI
xv7aTfyXQttacupJXGAsPtVyrbDdugT3YXZjGLWrN+svP6BelAyZjxqsLXHxzeJX
6IYH3aHmVbt2RaxHOTOZE/bQo37yWXUDymUY3T4axWv7RNkZfO3YiG1Z5Q6pVaCA
ppfbV8ye+uNMOTz4LSXxYSod+sCXH8u0538WZHdMz8e1+ztHiP5uOeI4VpA41yYJ
XyE+skGi83fL8oHhPHAna6t3Smlajzw28krsr5f3iGCejY6II+FGeuaEPb6SeSKq
U4RSqxjE2FlRJjN1wuBrvnyRSJRfyICSst6eQfIQ0GBvmtoHXJ/rXJUxXz+XX2WV
exn3Pv/gxI1XvfN4x/h0F6mGMfbsFbbBHl7QXAlF5N1zXIoggRHmOEHOBvbg6GsC
66tnPg6PY24ADIIR6LbyqKdnpyDbPa/F8u77a+O8wvIsZ6i0FCBxr8HG84ThQq5Z
M47+6jokLai4auvEiOHsT8TmUmLm6KYrC1nNgmlJVFc5VmJAOTKKxSg13YAAvENW
VqdyE/GYqmQLmNlqH9wR1r3ltzAa2nkhhd5F70GLZDLXyCIsXdeRQpTRs8ypg97k
Q1ORbOSF8od8vFq6Nui6sbwKqQbggBF1zGH0Gxl8pT76w4c+DhHe51OM8hRc5AxB
EW40A2P2zDnI2dQ9vpaG12vbQdyXIFJbh/d8SA3hTWwf2/QhBACFcJThGBG7okHS
4/VR+8xd6Wu3StItNQME/PyxwhnI4MvKjM6qRiFfblFgPlZfTdoLE2PwqY+aW0vQ
QajUQvD4A/5xFODOmSAOnfRLf3/QSfxmBnFLZ3oxmLIurHutkXIZdxqiUb5uuhuN
XVcXIY/9JijYeQkRfDQam9L0/aSKJD6Pj6CoUcYO7XkstZ4ufcBJc+/C57Z1LBdg
CK4xIPVJyuB0O/LrVWKpf2+Qi2G5T03gxWb684ITVhA7SYu19lWXno7K8mMtmKJy
ZepG/weqnAlAA0pGaJDoPm1Y6TsrCt189e3mS5H9YH8dw2zvLAWq9ozoE8gXwV6s
FxP/yfmg93aMm8aFsTj+sloT3V6cDtPRKI249I4EMbfiKDkkjsum4+i6hKFkijgC
PlmGMTFTOMO+UOUc6r4i/J5pAdxUWU3K9Jhwa/xVUkElb4XWXxo0HI8t0QZ47C3N
A9J7k2ktQz069109IWQ0blbZrsihtCONJqd/kYor8ZetHFMT1CpP5N0z2IYrhLYp
P0dalcOvp8xOIc0qtvY3VMHUy8XH2kNR6RwJk79wRE6UbxPQ25YrT39Gna+2DteM
nPagkdtLvwtUphDvHc9tBUONHvWpTSkCIdb9PF/UC0N16id4cOkjbXd6nHEbLyBK
Cr6lSgUQvUosagM7c7Efs3nAXLnuZArPQ4+0aB3w4OXReB+Rd4WfLSVrjmqVo4Kr
TvJzGWLfdtXZF0YtrBqGSl0XcDWKCUiYXYpYDWEwbrpT7JuGJaB52/O6UdtbkFwq
psa9I3wMj7kxNyVoUkOAeULqT7a+HJ7zHpg9h1S5HVhKTQCO92SZIZuuk8ArlzKo
hx28DxP/6qVib/vSqtEWkTljOy0mIIHQjN2P7OMn1IphIH1b1IAKKA1heQ2aw/e5
0U5HM/mCF260HPWOrz0c6uzeNbKd0u2xTGM9aPe+0+yBExvtIYgmhcv49+1T2Oy4
0NbChGIYf9lueL2gFAUxycaUBNSkHgeHYENBsUcyHdq3OPGsBTh7dLUoA1PYhES7
T3mGP5XsWLEih6mzLicIs2XAfe4tmAzKZ0yCeFWbiqbywxGJsJrPfHlkw7H2rkwh
7Sz3UbkOe1sJV5Fr8vhJTLfMya6tDw2H89wDMa9SMRr7sV2fn3vENfbLGuvalyUz
A/uvQ8Zxl185JfKdUMMplN4STH5q/vzd5ks2NZpK0WQ7OtxU7kbinyxQlfqo6is1
n6rIeGBQ/L1hWO86P7LcrRiezTa+ysc56Zud8xaecn0paL6Byk0lKV5EkRKn7SiI
K945g37eeqBZAvBuIKAm4dBjVTxiP+HW+9o00Q8amrg8TQwKkgCctqkRqIMAWM9I
IBl7NMCm8nRrqw31NYogaFLA58wmYDyZCwBHPgvZlF+j52OSxlDQF2mxeZpoDfSX
grdZeHD4DZPX1rT55mYF1jfZ4JgjCtZotXi5ade9PTQyX50C3bysXSyDX+MNS6np
rVMIzQdjUJ+dDp2bFf5Wm2YCmq4mwEN+jQ922HG5k/VtV6RVgezZ7Amm6325Oj47
DFt9Iw5VW4iKeVL5Y4eZj6dDHW4pSvoWyfhYQxsmOjNEJyvtwfpF+MsZzyYS6nMU
C5qK+Bcks6Kgy/t+2UqG8MR7q/3QDwd3jRsfUgZ21kdy12I/Lr679mdp3xiy4YMm
BHg3yxLL6iT9a1+zMXyyHzZc9Ju8mucV5uLIZtHTtWmRO/Zy7p748c1QvihzbLA+
53SGxQcedMRcye1n7sWdBzUnd3D1GRNPK+GG8hmm6ajdy0BaraaavxsGkGk1XI6s
lffJYzFQnH6G03Oxtqxtq+Rsp5p2k+3IOSPIW3/tOgfnSBScjoAmOfXHU7biPGaZ
lWBy6aDp7Msh2aFUeekIcEWoY8ip9pXCGNUj5vnSXFsDq9sR6Ai0PZzuEBAaZgYf
9tqGplUApoQr2osQwz98j4uHNspWo6aJUU5ix1aVAhJ7wjS3udx2ZzlzizjX7rjO
XbsDaMsvjmySnrFrLteQhon317XDmZsR2iFQJiP02zS5gzr4642F52Xvu+CirDcf
SyQFUCnSQQOGrCcMGFl08DnjcoUJKKRc1tc2sslKPYz96v6hPHmSY6J6PZrtTQy6
10B7dYwpYsan8hcfTObPxyPpUc2JgG9Zz3Ti8UG6LB3TxOFfyZaOI8QhlrfRKi3z
tKrksxwgAfHuU/7Bi6kaC2BsZObFWc72A9H+mKHoLUvKgApc2l4d2h/GNQqyA+tD
fvi5vGDllPK2NdQvO9QhxCPKBTKeevKUvMdtDVd0Njo9+DbpVUqOMzm0oxc+ZKMt
390MrOxrwYQKstVRXMbyegvd13NExQ+wCxzVqj1fJ1S9HxYcpe2+El1PDfOWPahl
Ezw06OD46Ir5VADYaJUWgHX9W+1gBy/c6MBsfCxM2LVf1cUKFg0nSFA92ltiu1ql
fAdZDSZbjYQdfrnKMVSQkzdAQJ7hcswbYeGsU8rC/6wqhSt3RI52KumlKpMWo2HJ
kcxfGNLw8Pfj5s/gjJTg7NWPSoGyyzw1yS2FvTahJ8noxyGXdUqKBzXLYg231mCp
0l0x9ixQDA+s4E8OsidrBNTliljE5He7P1E1w6iPnH7fyEwGyEd/3HST0pWmEZZf
EHF93KEUOAkB2VAY/nLP0F+yLVEPN77dPY+2N7HZjwAJAtyh2ZuTH6INafn7ldYO
R4eVh3YO7vKkPdllrW/JPZgp46CBML/bljag839Z7gzAUVN4dGuhDFNDPSGnDNFi
6ta41TdxyfwQcWyBAjPNj3dCKIJPU+drtH8MjCMJqxFKrwxUdCYcv3c4Ggqtctt/
e5/ltp916QEjCSgiBd8DrWGMJG6zo/oe9dH7YoNT4Xn8giB8XcglEou51RAHWt4A
LiQCjSa3dqsY7RJKeQyVAKPKipChQxdChgdA58Bev0wYCls86vuEmCUmhP1nL8il
Ly6W87ib2l/mw4DlwBnjrYXaRIeQyn86Oo2QbK9Cv5OH3zhBNA8bxLyHoqjkeryJ
vMAXCWe2FXckmVa5NWNkVboNea2VQbDKrenUQ2XPTiWIYMDDbhTiPYDNV0VzecGG
eSku060erS4MfbeyZ+Dt/tijRqoZNDLNfq2qhZLaawWq+SR8dUWj13elFFLsot7q
yrz2K5psXb6ztzWsR8TsG3EAo8hQkKygTHEzG+xRRbqZFYyrHtU2LXWHQ0Kp7yXF
Ye77wpnJ90syAtZovUNKNTEYFWSQIvfAkiqtzjc4kGxvRRddmyR3d1isu3kKRuA9
pLk0lvJJAzZGvWId1hxyC/ZKz4BQUlGne2kstnNDZ7wBSB9C+EemmRiaJGo55fRR
ZSrONV8ayQg9J5bdeBI2ZYzEijQCLXXNhTOtAQRU3s83qyvkmA2dBvrv6qI7pbjz
L/4DFBaC1My/b21FyXlZavNn/80Xnc2Fpkp5JbRHZghDoTbQqKT13aiUhDxH2mvr
ZBht6OQoSsWs4ux4f7Ggado3W5u2oFm6xk1huNg5dlGIG1ilZ0AjR/TRXCoINZAR
ftQYHKqy/nAJspkK0kJ/+oC5mdR9HSFoIY7qKE+38cazuvGEdgvTC43zq6zY5YCY
uNbYSgB418ZQA/AzXdDqtQDOh4nkGptXNffv7MPbiN2Jc+6+BRZTJEIHTRHGlAzK
95FtIlIO82VZ76QgJs+a1q8XYG20HFqKipBAnG2RWhW8B+2/Pnk2Q8gxmw3V68UF
yTRmyl3Wyka486LUMUi5bGk5irJHvGbKomTPYtL1xPXvFqtSbeQ9YWwkTPU8jOxB
QSJjIKm74KiOPNqqvVrk9W62OR0By+TO6iAq6Nn2kIWZFi2vI3aCl1lTIJlH8qDY
S30Uha7V/f50lNsqCS7OkzjTFP5JCuWR5Gn7JlK7EZ77wLMwtFom/A+nbpFFjyiE
gmN1joTcMaY/MlNk11ZmV0b2Z5lRQ6qehxF8UZLP1YkD/eGDiL3D2kAZq2yTKOd6
rTgnSuC6+p26Rvmq8+o6t2lG0EdM0PQtHB8BGUpM1C7eV1qkDLxoFACu+AsTUBRW
KrmpssbtARq8/zr2PAy+50dyI4ZN71i1ePyelFX4/+mn+ogxeqQfEadcGtpUFVLR
3HF7gxooZ940QX96/9cJJQD6DjF+muqc5CNg7o6ATIKGN06vHBWC1PMQFSj6Tppp
uYIZ5A1fPPnO94EOYWSKxwkj9/aYNgeGVdXghK50CR1WOPFMWf+C1kOfgRb53luK
kWKLOHaWcbWqicKeeJfHGzHX0RxnRTMe+XdxqdmYEKECijnkuS8v+XmvafqMBOLa
phsWJe7HkDX4IgzwE2zbQ8/DFhCE13SH7BNftLfyzBYPZ1iZFxTgA59V3K93SSkK
6NGlplXEHYeJ9sJLNWwDaFHmFKkXLzOx9TDalyjhjoM6tR3/wSCQ03+06CSaDgXW
0LnGdCu6e+HDvSa8GrMKyfO9xymVVb7zDTOwXG4kBFPtm8nOhfkdxFwmujRgPqve
qHb5ZcMd5bsm6RPw+yW/Bj/HuQep42C9SxUGvg/u1d1E7G4ibUgQHoZUVlXx0tSr
ofPxcBJwxXkoOxk5bcChUCaw3N3OoVXwS8cDZRrBQnTU4KGBOJ6x1uJBGcNyM3IG
kzkvTtxC/RlfQvTHy3E16OkNbAnLRrUeMQkc4Ak+shntqPDbyYXL66SHSfGg/Yeb
u8EIyalkl6hInB9D/ufJztMyrMe435mypOFdglP+bupOqBZTOGv3U3jQQQDs+FCg
PLNuuUdJ+672v5gYMzaPctDSvV8xPj2rOR1JBYUi0xSQnlgfVlpbdM5EULF3yPdt
lIwSQMqstfsJE6KOe9NBlfj10rTFz4rG49ftJhSKOH0yV8aLwr2L4ynDIkaZifRy
t01LG77vVIDyFWvW/2EBVnWfUR49YwNiy5PrEBgLODYciTksnf8WDLOeKwklkhtq
QtB7yv2UNdksrBM3vZgm8mBCQIE/mNN9EpX7GtQK7RC2Sz6nxZSgMqwfz9EotTAA
qbkZaSLYk1nNSR9re619zlRsyWDjwSTA6zVa4ekgixM1/rCjRSDqfrndjN5m1TOL
aIBCwqDv0vd5P0raL+hJP496h5baNv0imXuec9nOGj7RsvTC5Lmn+WBVPbCSiflj
9bvGzsEMZi7qk0XQ7JNGaHMYOAvAAw00ZRtorUxIZgMRYxWsq0Orimf+ppBnRGA3
fSbktGuCFZUBtyMBrYVf/bXyOQXJH4NoWEyCeG1xw7p0Xm4gJLi1EVqPAUh5N+1u
AdcXtVp5z5F7ttIIOPZ7eoD/1+8pjYpeYjeQZ1+GVGhzJ3eCg0r6cIjhnFJjxgRX
pb1/9WLtN5rL6jC9pSBJp5QIQOiZ8jyWKwsWRXT1XdBHlKNSsIfF6QY1Y4WwPBxZ
w6VGppX1VcRyxD+LTArH1kg/zybtARoqghhOdp9YouF+JzzEI2AW2HvNgkXpJZvK
Id/w1Q16ZzTuGLfswshd8eVj0A+p6saF+yNFK4ZRM2Cca1dvXkIOlHq1F6/74g7K
96fPHHygQrzQGPubonxLFFXgboRJwoPppAwo5WInUZBpNPvPIXwqnnC052IVZL+e
IgL64QHeDP4tFq9Z/QXLzNw+Z/n3IDF59kuwokNPP03MszaFJGoWtIlZinS2MjKk
LyExZc+xd/X0iLJ2MoTz/aUviYPcsPq0rbbL3SYKlS6Xhdn0AXpN0ithFUoEETDW
nwDXS8a6Q+oMRHxCErfCFve/MSydG8D/tlAXzy/iVTy657UJMhBKyTianOwX5Bbi
d0n0RcZrRIMjmNJ0q9XOHBWol76XOaMFEb7Ley4Nw23mDze4mDna6KnQhA2jHBbb
n+nWIPdr5JlQW0oO0WToOL6CbrywxBhOty9lsAn6JZtexiPEJQG1q7lWCLO3nYbY
O8sNZbxss4x4iS/pXPfVovZIjk/QuqLU8ZODXBBCHLAkeZ9eo79Dd1pRqt/CmcDZ
UVJ0XSuRgtF2If6J8YJhCygXjr2O2anAjggQTevJ55r2GXu0/B06u+BQMSxKafJI
fwPSlAtFQQsdvB69bseZlSoe8bN/96BvinCAis6oQp/2mHhA+IOX7Uj2Rz/klp2Y
sp/1fG5jMf3+DK7OMGsZyoqJbG+AXzS1xcbW7od3ZqJ1cvjgcR+m9xg810U3zmqD
ZCNqFuo7eyl1bOamNrFbPJ6NUL7XuTnsVhSFGZiKYUR2EjhL9Vo6SiNDEcSFMxgQ
9My4Km3DchW/aO47OjvMQiacZSs+12WgRmtmCbqLE+FKfN8lP8O1wMnHpsCyrQNu
Txl35V+C0H2Ri+FSTqOT3CBLzrd6WwU2XcOkvDZh9jbwFziZtbqBLcn9ozvDGYEq
A3xpb3RWQujfTTvc45gRbCdGthRA9RKF8o6R++i0h8Hn2vQCzdUxAcKqz8x0tKkJ
YSclEyckdqE6pPmqs6JZpCYfJWA92nrQuUzHoPMgcQAUHjtIR0h8wCxyBdwBBLAL
ZXG5z0eIki5pmfQiTBnzWXSxIrvqnL2uRS8kCph7TMgvUXiYAEAERTIZ0AN8OhQ9
5HBdWIl3EpWGd8Lu1X0QO2f+wUYj+HbmILYnGF51bt6pnWYJsb6t4xtt0sWDU1G5
n52eY7pfntkF+DY/BUZq7NbgBKVMGzvrNuTXYqJNn9lEiYxUizBBzrGBjq7iol5K
s4xU8xzf8tnFSKvAJMbOjbTm2EB0tIqwG9cC95RGpd61SiBt4XWfJxzAJB/WjHrf
LjyNLVOXVA2GxfbC+wx92waQREhPTTB1RhtaTt6DclLKxQyNmyCBIatkJyXpeCAF
4bv5narM/p1VY2wcmsuA3MZirO0lH6o5m7EKTFauxRtWmjnD388/r6W5Tr8JHPmb
K55uM97MFGmYxCVFhJG0445n7k1HkYdE/wQdd44meaOnBbwJoyOQmbcG/iU6bKkQ
pUQYVis3m+vz2JhBTzVioH9EhWSV6NMXON0CeWqOeaJ6hnYQTlH6frs4NKRgci8B
ALTS5hR9hct2UsUqIUWLqT+9YFdiq5yFfcoUBnPjb+2t9g/ds2PEbnis3e4+VCtC
qm96GB3cP8sP4+ldTbLFY8VQrImG6LFJms8c45S+rGM7EIwaWMX4mfclocWIuQAy
XmkvOLGcFrINbDy+VWEnBciCuM2fcMpN8eTz/0p3umpR+SOSPF6T9j/exOGDx8pO
U/v7G+shuM01N+fGyORtW4z3Z4qwhAT8q0AtcDnC9zZZuCCD601SwYyBCdkwvq5F
KJljEAZ6cH+dxK4Jtr9qYptqk7VxuLirMofznrfOIDtQDWsfySKHc83O9rgZNxOB
voC+CicGetxnCA94VxnGlP9q05aWP8nkQgNXLvs4UOyoMug1v+0XRIG0xhH+WVtu
7iFj0OpAJcifFQFDeDq/4kFf09i0QP5kDPQtM4btKR709/L6BdoOZfHZlESRFInE
YY5BoZZtVp/RLEJJHzRv4DTSMzHtHYrHi8Y9eugErj8hxe44J8zMrtIHeZ1vDVIh
Fra1XCwdxOby2wTHW3rHPIG9Hq43wAYNWl5W6r4qAIt498oDv5TKGRNRXMsn/hb0
+s+JEyzQI/t/T895s4LAGdMxvtBxB7tWkKSfS0fHeJtmb3bMUbMP0TEHqkPSQF2m
oNeaGerk0kdFY5EvRidoRKKSBan3y/3dIPlZSilE5nnHANQ/5qOBhAo5YWZzlsjt
jCumlOYdH6wBejKO/0SBoruWWJyCigLj47QzF6xYEWSaQmZ9i1uwzXnjvdc6qhj/
+h4veGeVngGo0d02Q/kw+5gLY3FlrT7wEp+Y/yfBNseBiMC3EjRrc/rinTZTgj2i
WIp4IyGNL779XMvsk5VqcJK2O7DLkkSioBu3Ckg/at8tkE8JGhfBJAJAMIezPoPi
2slkv5Hn/3UaC8lU1jjXJvA5N2S0BIOGc6nynKp0Wfkoj/U5OgxfLXnCwWJgINVv
jvvQgTCjXaDhPCz8WqbaRiGE/9+Fzvy5MaPd6WLvQxP18U3rtt+pWn+bwVFr0Vkk
litTiOUwvS0hkg7+rqXImNfpnGe6nozvt/qGCpcQfxuOjnrMQfdGRsWgn0bDuCBD
RXyKkZG4Nnj3e8WdJmzXZOdxCYqUaQwCvAqMJEWRIwVf+PUDjn/1LA2D3sykqoMD
piUxD39ILADTSr8r67bhbCgpBWwrgu9GabqZ9kYiaOT/OjTQDMXomCqpcL5wKSzR
NclwTv9bYuroI9uI26RQfMmvTpanAOuuIT03bPfgQAm5EycTGR83KDI6glzVmaMp
BTHOVUtA5LUqAQfKOEEGoHJzDOELQ0N9t/lPrPDKQEBxocSoRLH6VVrM0Ri/rf7R
Z4saHv54zv9El4+5PoiByKYC3kulwSqbQzD62X3y7Y9tR0Px2DDxPggKSE+O+qZY
qfdqoO00pCUkfj1cWHkI8v9NpsHyz8uEUkAsTWkiS3Hk3NT00bmRYgJ+5l1dr7aZ
bsO+UnJJlrEmZ/q7F7+5GiZTcSj1d9Vrk5CZMwmRTUMlEcsV6fERMHndjQF29T5K
MaaqUSAJXPHVMvhnaaqPW+PyM88oDMTjr6pWqsSDmna7biMuNxMaH/voPflY+cai
lzvQbf815S7fRpQctWrUvB5TlBRv6noSPfecSNpDQq1QTN8zz2Q02fzYt5NB1oVt
A80qQapksLEmZNJABN565pRWPiRy2lwUl5Bb+lH4IEOZkV3Oc71w9WzQ7fbRFsan
dTc7XuzeC/TMG1QOMy4qVPFsKFpf9aZRj3o/n707hMvu+WiHdsBdQX97JoxixIO1
aSxhp3F2m6A9U/9MxpKlwlpLAFrKjN9DrY3FfAVvYqWADWLHGJmQg5ZgsJYM6uP0
ENRVBf90r+4kWx2tjCyudb23uybMXQIFfNRHfKXr09B5DOaLwLxAoAzUwxFEtvFV
7CRZpxZMnuXsaGO3hVCZ04MibDYlNnfQyj4YL8Yslme9/I6Alay6HLeAQAHh5e8r
/uUrvXbhxWnlUZmT83cBK4Nvist7UroyG/tINsSVZFlh4JmTxOJ1zMbwbwcdxJHm
BVNziRzT+kHN1KxYUhNWZf19zb8nGdB/orCTj2+BvqmL41B2eBdOB53lwJedzQg1
UdNOisGq7H/9oXeN/Sic9pobved4eJUSkUxwYwtqEotBLOtL4GiEhVZZZBLYXSUx
i2kosYFl2zGSG+yRTkq4y/E/ZYHJUPLuGvYuLmswGEgEntjrZ8XWDjpYZrvbGqdV
j+vkN2SP5lXvNFLBFFs0wYpy5BvcM3H+gztQvJlaNuSxORox5U4/kuEBauow2gLJ
vZBeQ8SjRpOEIP6NJVMthIBAkMVVS6vQKzpfUTTnNqOxwa1aTxTPcBBBzPZM4hn4
Nfk/QTXw5LN9lG4zyUHRxcSLOMo2nz+OLtpmdPnslCYiTsYREqwCVQ5vSSD8+FkA
xWaJemqgbvRfjT/GwF84sW6Q8Du5h55+dc5GTH6PbZ9d5Pa2cT8F5ze5SiU/r+8o
4kHqQBjKipZ0pEzBmp22oAi5KP15mJA1aS7xba960DWc6npd7cxQ5hePtp5EUJ84
EL9UyKbc2+MeVE0K/Gmr5+xjTmu85seDNwtGRUlMJGGuePGfxVdDTAPbyDUiOeJM
V8xb1wv3JheQ+/Y898Bpnuon1QO2dAdnO6jXIt858qOhPf0aWVrWAfi0ikvUJ7jS
ZuLQhihM1h+x2ZC+bOJRsn2o+PBrtzeQpJ1bFtkcKXJ/iwjkQzbskRlMuBuhqrZ+
MKVDAqO0QJaJB8W59Dr0TPQHEJDNh+sIWT+4ja4WJFr9clJzIvlsAYQ+3pvHDCnN
Q8CJOzzz1Jtg9sLdqI2nnHdEpRwyjsT6T4qb5MI2rPkwiaIbhdI3JazginJWpzbO
VAE+ucfuKojq8ECAwsNzhMoPJgP3kFGvdfew1W9TX5E4G4XOyHSNfCjfbKnV4+SJ
hwj+aFi3kDSg0geNI75ScUekly3Evl0EM2CZMDS+2OkE5/lhCha5B+gr6z5ftUOF
dsR4tGuaddooEeUQ34SrFzIc7o4VOEVU63mG+XA+x71PS29tGmXzjnYsz3b5xTCU
dImwlXPXKk07VCecBr5yISlFnXOIM4LDYmp6BwqHirJ0RNilZOJnR8lK3A/OgeNB
xLWa9kK9M9z3E/so4x3sYNF02V/o4o3NgVCMK60mEenv1MsZz9x03eDFS1r/aQn4
1ak1s28bAHODa2xjFZnivraVeS/QUWyNhVRj8UjVOy5O4wJZFZDlfRYAXcJEgvvK
1j3dLRN3Z9BeedLoHtpHTAk7JCTihgWHFA+m8imj33VG59R4VjmcKM8xA46o8uzr
YtE0dd9fxHxUn3Civv/Fa0EYY6JPqRN+g0qco8NfSZC/fvmSvYbRtQLxV6EPZdHe
kfSulYfVEjrgeXt1yI6NA3rmU1gIsjlyjcEgs/c1Ihs/ISr9zb9qsCwsbbJZDMuk
RcGaslzInlR3b/zuQ9Gept8b7WW2/ZzYoCzxaIVhExlv9QaBX2QbGO9OwWOz32wq
pi8jeAM1a8GJk1ko6VrciAAefi3xL7BwSz2vIr1FqUeUPF3/ZwYgCTx64iRtRoWr
R5lhXCeuLjJhbw+Z8O76Wcks10UsgTpNY/cljwB9XJQDVWeGaxK6bK4tz/YmrN2C
8Aa+017iXoE+EXOtlJP6YEvIyI2VUzWIztzwTFt162t5wZErs1NONJ0gwT/cCX7E
VwUmnPFhBD/HHnMCPdgEKl1MjVinghigIA/rDrBCzt8/HpsQwNh2JkrYhBXaGl3U
Juyd08mwQCHt8///y+ukc7AsLYA/RU8TvMFbo/ePXThYQHUuX5Es0QDHvTzFI2Xn
tR2oAYVjZZ+K1ZbtXg5KeutYC0RbrquM9+2ygKom+EkNQw2sFDOTspPPoMpVxE8X
Ee8l/+Wdd243ysTYkvyHgDOb5+kVVNiSkIxXiuIb0NHki3wy3h/6r20lZ+Q0tV5v
QQM+rOetpP7v3VmFIZlNBtSoeVy74Uj4P8l4z5/1gYVBkxgbxmWQ0IVuB1xYsPrw
W3f3dGif69Un+PiYwzCByEKqJfXFvDVO//ZnL0sbyQsPT0ZFgN7c8VFMkc3vZitH
UKWimNZfW6IfBHwGGqJA5DMvpZSYmdtSnFthFnVGk/z1FARs2GbCFKCywfLiLVyT
wXfAajr6bHXliAjNJPN7xD5UvVhP27RaHYabQR1Cp/yUEK8Ifk0J1WRN3F3Ooy/y
jA0iZvcTqOMBAz882nD8ASfrcCthTk9Wz4Xmqg2BOHvSxusPrGUt+g2XbUrzzlZW
LIwzMtCrcBl4B2+Re6ri85tVDzAceDuBltRYyFpzKKBg11sh2KjqISnZ4G3kdtLV
356xhi05P7ZM8LCVOD1o2eCHDGXG6rG3hX8ai5sq5sjZx8zztHdAP72ubCIdDXty
2FnhL5NS+d9iAiguzuGZU6M0ewK9SjVHWAmPAoio+4tSwzsGo+5RwoxM1yIWLkR5
0P1BOn9Wmtl6/ZJESoxA1sCoEOcH5wIcK+D7O2Xc1KKoXg0BpK+0hSEPUmZ3GhDg
BsQeQS7W1YX9ztrV92pmYkvwh0z4NjsNRBMyGPXRgUb9B/79MDiqFM1VOOmEOU4B
iuOeXt6zzamPMqWgArLdX/d1n+HBQdl0o2dNTmcgsA8wng1NycQX7q+BiWIRhnXv
/JMD7V7ip6xe7wxix6Ghf3RbFd0Ajd9b1/o+RbjUssOM98cjqzBGRrXf05dagayz
WMn0tF0bMProKMp1BkFI9sCab2dhwhTgyfpa7Ne6IwC3Z6FgqUaEdB5jXAuL10Xl
2xTJZxf8k93RUbXqq7AQiM0ixI7ZeCOACZLoO0bRDdf2N1F3UzJl7ll33YreFEOr
9be2FZyXKpBS8pdtUfeh8AbJBDmmt+8766z/ivqUDiI77DGOLlaWvGghRD+BBHhk
Axy3Vnb5fTlhaT96uRnyAiQCEsjnVoGyJEYWQSskLX5gI4zaAqpFJEINOmCndF7A
lKoVrfCgCNLA5gcX2FY1xAg8TjK6RShBossmdvrD1T/BGhHN+DOW8AXCqgs9hSav
bYMCqquP68WGhMmgpmNGA2hyciTVB9gXXBlXwbUeyxoXEHwucvCR+YtMQ/VTAYGt
2fuxq2ssPiejlnN9YKLnnZ9uC8UE55Esr2OH1lckmPX+v3gnePWNKZO8RqtS5+A+
3PRHKtCjcfjNXzneokLHJ7h5ldrxMfOSE/cFYaKAluTRkT/l2OyWAz/iq5Bg3tPC
6QWWvfeTbVPdMlRVSVejKBz73DJyIh+Y8o4J21suzMbusAcpW9iJ0lWCBYqdSnPn
2cmIgwmS2TzhZwhB6sOBGR0ZFRtcXY5Vysu9XtEEnQu81AE+NHcTPU/svF7NLVBL
0QqJguaXMFAIJDB6r0q5RIEqXRUvXYGcxUJhthr/xjnfl6yXnAmRmDmKGb8bbLvJ
+EZYqPi6x1IzjPou0nspBPWB6nz6ndeVIF/uLeQiw8tSFLReNsC6bILhsYNW6BxJ
Em7L4PND4avXW2XMJ0TmmJeH0SZgoLY5J3Duc+VDV5+ytpLNZdoEf4cbYS9k3oZ7
Dcz4vaewU2iaik6SCi9qIAlu0oXiJYYUcZCEtwnsmBXuNJg86VC11cTl4CDOOI/A
19pXylN0/SU3saX8S2OmzldUOG5OmgYvQfePIgoMoyUqTkuWMCrohueYej8gx+fb
P4Yh+fBvGtzIvZVghE/mlQO0pykX/p23m0xsWv7QjgBrfx6RsRuoTPTCXbdVsKhp
FsKZ2gBsxg9J9Fcquisc3zm6K2SOx3a0TBJbjsts85iXNpCzr32xn0wgl3bdIYJo
4ka0JJkH8W4drpOL5N0LvtzM98cxQD9ucMubMfIZmrmab4fGVxAYtDNUkWc6uGGz
Urnk7GbbdXDT0CbXkHcmQ9Rc+Oh9yYmIu+S+GVGDMANxF/les5xMrQjTo7rQ8hDf
MRw8jLeE4peqxGR7zIrjJp2p1GmTgaDJ2ywo3f1d9oLbq/B+CeieqkJxcI9BKHE6
00u846q5MIhl+uNO5n7ysvrgzP8uN9EGq/uCAVdwumcYmpx8/A+lbWcD2dX/b/it
3H+im2rOdrMWHPONDu/UeNbhUedirov/nYgqaorXJEbS8kiJyDHXU7ndABZ/fyBh
+M89lh5IlYaYbXVB6Qy+pti6BthAwE8p071efHORFC6ZI31QkZ9ZyNQgnhVprezy
mfS6bizl99lbHVP8x0r91MGdREqjoQl++iXVZ3JV9/4WBy58DcyH1vEEvnTp9oIH
KOXCuUZw+Fg1x9aNHlyE7CZcyhX6zSmLfhGiJxc4QZEzIgqb1bO737eSVWxfhP9M
Bmtnd6lZk0cQHOBYyA0nt7yfigi75kYysDt/qoo8MW2I04bLZrlklwcXZ9slwH5e
7XYk+e97TMKVuPIb98r7YcXiTpHJYho28rbAT0CrRd8XPyVzjgzuFDb3TUm2iY/x
2sI1dhUpkkpbdltQuxd08nDFUJa155oNveyM8b/wKz2i4VncPu9dOSKOzS0C7KQQ
N3cXdrp+IFFotTNYSYWnUTgghZPdFdNcHJJf7IT1xyqM3OHZH2SVhH6XEaI0NFhm
ZLCm5oqHn83eKMBXmEtJkbYoobshQQ8RJEgpWoPvgerFmGeGJxsRv6xfOM3qHdaU
iXNyQVLWHM4c3xadR8lzBjA5TMao/+IwhizahYDzEWOZDl7Qlg1YhuVCTrmbQTCD
Fv8eqvYdaqJXUjVbCXeEWqfTP6ij9M2Budqg9fGdOKFmBmIKW9XZ00COukl0CKjf
+tRt9gTWSUDC98vRzcloRy4nQABZLTf1Krs07fr1QG67i9zliOXQKOiz18KOlxNL
prGSO/St0VNAQUa7h1M2eVv3VubBijIDBdBgJwkUJWqEtB+Nl/FU9SL5i6C52+gn
YuCPGG4vaGRZHufNYw+TS8I0b9LHr9OBtMzlvO4gvAR5BwYoGsU73ECBxVdSNVCE
VPdOfi7c2HHHqOYrisMGq1jJkcgrruPcSTK8pHpFNYRANWaisjSXoLKsCHISUT5X
PU9ymNSVnQQstseTwP608ygzShYeTtCeT7Y7lQfs+Fk7nMWFh7ef54VEh3OuW/Ro
pjlA1l7AMVkqFLWANP61kjqUK+ILIM/DM9TJIcO2cxv6rDZwyjCfl985moWqAWpe
ADGgZAIzB44YBnQSF/M1eVeoo47cM0SYIzT06cHSegxHeL8MUNsKY/yTweVukSWX
6snLUD0MW8+so3ka93Ewap1DLHczxwh8j2YK9958hQpn/bsfX6YgPB/1YdOELINI
IGrpdm1Td7iLKhYNuXI/3epg768k8CKCj52S7HgkDWejaAcIX0N9rEdMhQo428w+
yjXfzsIrbbdTlYe/vkCHUtr7ifrfqLGK8LLEh4Dkzewl0tAq9CV0rnhZzi4URALC
C5u9SRSY6SxEjpDnUAZdipIZQUzPG1i50A8uiKa87cWxALV15CZhsStTbCuMEOhF
YK0VPANy2oErcnvSN3O/e+rSxrDlY0zdn5//gxyj+Qn3V1APUlg9wIrY7wrrg2SO
RCnRZkta3/S4iWtT8edWoLgyUDb1Mvu0sty4qGaVPORBImHSB7BQFcMz5zSt7eLO
4JJo3vxhKBDG0TTpWu/3oWxbCVsfSkTzIc+k+8vmnAD5EIXm24hrl60SxvydlNAI
ZoCXDwFzbRzaLsfMO/9xYIOjC+qxuSR9BLuu/jT2XZKWVhU5++oCXclJZ2GYVqpB
1ULTlQlHJleaBQfWzjDL1owzKs3hU84p3JGqzMx9bQ6H4cSdp/AL56v8ktBwi5id
v/HgXwKgjxrt0uQUsKMi7ggdxtzoTxlRKE9dtAASnTgIYCto+ijMTL8mIf/rc+4D
HBMi7zWveX03q9BFNEaBKmz3YzOgQ1UYeXJRhNhNdLqU3dobvNQIH3HS1uYrawJ9
tz81cx7+SLZMSD1eLd5oeG7PSIYmtExSJWUIkAbf37xbAH/vREK4SERS0XX8pDdU
FkNiZNkUgbxdg8cnrppKrWv6xmNYWDjjBokQA2eMO25nRUUVHjEZ6UDgiObD+FYi
D1+Prx9n410jNRDtNkAdKGuY1oQvja7KicMuEBPfebRpYqUf11PrjuFlZE9Ep42R
WQNeHL7n/5K5/dCkcgZk3lPlQjj/QpKWqvB9JZZEXhPghKeVcZ/HzO0xW6+raF3k
OVtPgpAWHjp57TgTwEul19Bps7FiQ7a7bBjAXnmsG34kEoo2zlPy3pzYxxjgs6oO
DwyTO2GE9zPXsMYmJM8R9i/zbh2Iy8Sw4lw3tJSMC/pvc2H5hUMw0v8FEi873tJx
y+8l8BTEwu4oYp4aptvhUTe8AGcxtbXTfHWr1xHV8ERfqBhRQyvwixKJMv6HhdBT
XdXe6pWoSDfecvb2WLFn5aoJm4wG2tssXdLo3L1XB2skMMdziwmBVjKdRpVH60MX
AQX1TbTMUtgeIc0pO8i3gj98qUeSmhzDiVnpoSWA9rmbskmexgPnKYTvlO6A/vaw
nFhfUSP/Lh+N3kOl7cVcl5t0pydbFiXwe4fAgo61I9hhumg2D47/clQ+SfJqnHc+
UBY6pQlDc8EjzTlRri5LZUpNjWN6NoLC3v9AJfiCRWmmiJdcOUa8dZj2AB4tn24A
jrUJhCc9iuP+812xVF+wZAkm+d3j5NHFdb6qI7FnQnvlBPivnf2BtbIvCGINNOiq
oOoO78WqVOIYmcnAOHY+Uw3ntWpRlXM4kdMtvWpWecDrdwfZ3AB3ILpCTUyns6nT
1lpUA8205HlO3LPlSxV6/sB6ZLi3zByI0euhhvvMniQHipb4v86UMzpmVRlYv73m
VMsHLB8pdHsk/ZgU7wF347yv4bwHpp2tg0P7ESbKigvW4AuqqMi63kywRuAvmdfC
nnHS4Y9yxhsO9x/u3dJQwslSSSC+2YsD85Xl7W3pYj3aAIomTe49KyTfmusty03t
5R3tiT9Lmpq4uc42Nkn/t3n+AzChMDa2raL31ALTVyLZg2oACBzrIYmesQkR5Ii2
3m5UO5WxPPA1DaxGnrwVD1Gbo4TrB5ZE7cUVQUWwlFbz+UcVShmPX1pNJAFnvMm2
svI2MgNuy5leVxKIXkT4VqEgF8RDZp9u6AvIgkO68KecU7prHHsTx0QwIHWhaqe8
zKy1OUUXKl00vyaQm2T6s3w3IeFHNiFSknmtTTjpgvN4Bc2UoCCaZEzZJKDEfoK+
BLetxd8+/jgBD+leaCyUv5ck8xaWDWZUHPxpaHqyHpzct2rMUgfygo78WNKYms65
wPgbjWJjTbvA1MUlvFDOfgYFPJPNydk6wrgw/4W/T0jjCpekNto7URgfBnzGrEjd
gUbTEKIEa+lbXVWfoqxB8qj99sKK1uniehUXVhlM2bKOK/qgIJxON8IvGt18Xont
D3yINpOuX9UpNL2NUjuUHcBQ0pqYVR49EI1HkDfkKyKivvHiXT7dDJXWqk/8CBYa
RazF7xc4akkPG5gGRnnjvxSmDAy7iywONC5xPM6R5+XrXpseygM4YJEt2F2xE45n
SAITu944nq2g9QkF9QEdGr5+qqqudn03rSDL3rcTCiEQXjZgWdRRuiwf0F3Yxxuq
S/1OluFtUqCNvoZtW3Z84zznwszhX1arvX9tJE1T2b4rrwoRxDEEVjtuCpJ3BIyL
JVQEqRcSbCsuqKraBVR41CyjxcAZJBTsxr8xmjA30Jo69hEyRDih25NDqKcCffhy
HYuOzYSoyrZMN9NBZvgGHRAKy3Uxh4JLz7i/uQ5YLaAY6FkleoLP5bkL0Shk0a8q
pX6bZFB4cF/toxF0frFBU7fB8n5yKHsvbGXOoo8JQRx8PBtfNOTQr5g+9MH/baUh
5WNAlaOrJZ0Uwgvj2DelNdDM6mS1yMHwg9GXF44XY4+jWjGPN4yzz1kRLW09EaFN
HeLibemRN1WNmKhnyBphVIz7VSl7JLS/l/SH0uxf8kkuKu6GqGWmph0NWV0uV2PO
4c2XFy0kuFpDnDtJRHHWkUyLZx2C1wGbfmovkG7btXe3t6VNg5IM2uhLt8iUEgG8
RnvSbzTqAE9u9mbgGj/iz19PPNovqzvyQ4CNcHYiZ7v7MBHmi8jmscqvR+as38Hl
ZKWwbRqflnqB7gxN/K8BGLhxErT/89UISXK4HowjPj4UXLF0BVkYxzNB1ucCZphe
646r4lkEtp54M/SMDvJPDdKULakXx8HJz0E4nfJr8WMoy+0MmBNS9if+2xJ3+tMR
RJ/+ZiCcMLDDizcMNLmLMg7UYxMvgHJoFFBI84idxbBxffznIL6VXUBn+6n7vplo
SAfpPdBC1n0WDOLllzzVhqothrr5UQi8yCBleQZkx7ZeHOzLqPOjlNnvWkvVgzXY
ApzMf7SFJetppLY0e95g9FJjLRqSIN1f5NYk5cWF9GcJ4U43sUvGWpdqSZfqOmkZ
dZxS1jWaHyLBRqNHYrZ2VbLh5r0h3dMRgX6fmnFb0wgr4iOG7UvtMGZ3uIjFQzC0
A2QzjRoNLC8r4tYJBC+ou8m/w1olcOX+uxDcri2oeM5IeWBBprl0J6b3Km0xZyzk
rfyePmg2Ye7h/tv0fkE4av9AS9hY6z126FAZpbJGjVA5KJnl9DiapFgK/GncDZrD
ryVl5XZ1kU0rX4BOqZq8mUNuaWydU13ybYedsCD9dON0lUrQomIc+ZxU4K6BjkHg
wWoE28+yMiZ1MSWuXC/aISd0a7pOfqk8U+zVgWm0P6mjpK55HPp8oe6tB1cdygol
WqIOzl/Q89Pzmks0yLreBD92nFRFMw/EMM0R5SlZF8iujyC2xiByNLPlJSbvaVdr
6uDay6C7VN8WH5sREzRQhdF/U5l9MVte8Dim/SR1PqK2DjOiXlmewpJHP+Y5K8Zh
7sSmCcdLTh9FH2uA2+J7CUKAgPcwVCuR5fy2juuhq5RovwRt41APbkofJmud1Hfv
x9BXyDHiH+gpibmuHimyiYBMXUM/IHuJJAxFRlTlVzenrrX4x5YMEVrlRK6OV5+0
oGx1hcQl2sCJNKhjgazHbKLM8nPcFPnKBIaE6P5A1EsmiEkrUYy5JyaAy/ti3+0V
JuzBxqBCl13s3LISHpwSOCGnaHrKygz7ygJQvUMbtipnfeOWzXjdrswnScJsp199
9jTCIg38Hnzfy4m+CiQAQ7cbRS24B4HR/QJVO84GGjUIRW/65ZmIli1nCVKbAbcp
ObBsdpwDchtjoJzxJT4ZVe15C9icJQt3gyWM1S4i9cA829P3Vx8m+0Wt+mT3kqrx
UFZ4OS+iZBK/rygClhQ3Ixnj561KmTfTIa/vvHQJbtZsUCOmT0XTfuk9rsHHWKLz
UFckv2TlPehOleCKLZp1jTxg8QFeiL7gPW0tTEZQbjGsVNxbB9NU6WRM1PoLfo5g
o4JseUTg7XsCWygKmEVVz6OlfLGUKqaWRczPO2N2mD2MiH6YmQW1MEPXUhiI0Lil
NmqTW20oKHTBDY1VH6BW7KhCzvU6VFTzDb1833DDjdFf4w1WFbeBvyDrcx87+0Tc
dj/W9b2kZmrmgjArSNmjbC4rpcp+9st6HBeq7ddCL1ma2RtvWpotiATJjbIb93gG
uhEEeCGQG2XUpsxV0d8fn3SqlHUsB8DBEXUASu+b6RzT7DD4P89gCs/QdoC41ftE
xeGYcoMYWPtB1oHEg5HjocR9dUEmp4ngR3eE3btQ5i2ib8W/HKiqg3orbFrHzIyq
a6F+yr2a6bEfzomTrYiidLfooOZBg4PfSjw+rYBPF1+3ZUCIEHXfpA6aVjsN2kUP
Q1bXTRSACYr0YSZuClcFbB2mzWOLv2fonVSdifY4+PSU8I+BaHDkGCVHZZ6p4B5b
6zBmHGMSK2xlbMVbOk/qDzlCdczlz0z1yDf82s+jay4geRifu9Qty0L4+38PtsJz
s7PPpho9Jea90bA27SfxVJ9jVPK0PkzFNMJysRaMCxXzs1WkgHsl73EhW17Cy8y4
Qvd7bHplmv+exc4Ui7cVMAWGUbEpeKOm4sX9lyB5ozhLKtSxPYXFkg6qaj5WhV+g
8pTiOM/ytTqSXIckajpyqAZanxVaN6pJkbqSxD2GWUMyl9SDGPVjIAskf/YnGr6/
EDMK5AgSZu36+ifXxX0nASTFNZM2pdPthmYLMzGyNzM8lSIJP+HTmElkfiep+Q1p
7TVg+gjv6oNyT5BU1iIMnl+Kwmu9wxpFBdKPq3HpwnOCQMLaYgDW3ThnZQfd+/wA
llBdh6ITQAOh5r6GUEhnafLx0SsY06AH19dcKXJkH8T7KFOzV0ZVFNkGxsn3ZD6a
u1JjfIo05Jn0xT3twaZcu89dZn5NAmGg2RMHdf1O4h+ffqowLB31AiSxtGYfVM2V
b6R2WhvH42y0pbUXocVVHVrqrDzeLtI/X+UjQ3Ptkl5PNPqkR3UVw3Bgr0oeWFv7
QUpiE4SJzMxC95OXgBhM9lGRS6TsnWLi1gw0gHUra123ORpKVJKmGypIke24+ZsX
4iaYylccXtWPolPjvXidQiZE897RcF2odd0ZW8UwpJAmMwNWGyVGzRhJMjhVmzsJ
9klocYSlOMSCgoDKuSrpSSEgBzXeepHJMWJ5eTNfjj3LfSa2kM3sI/aIK3HW61io
iQrzw2hOaRI/d227JZqNqYra2Cy79CX82nE927JtNIEHcEpaTMyRLsV/MpUmEAxx
RQ42ArGb3AgE68Qh0jehEYH/gl0tb48017wcWr0PvrAniyoR038ZrvmuipmOBRpj
jy6vD0W7E7HJ+GeEp5lQQIAPi4yknxsp6VEwweAgiL8jLPwursDcJENxOjAVunI5
Pkpb6UFYRrIhCp4CLNkl4UgQEMfzm1Zgz/fyDbMFWpt5dW6DlNvB1LC+U0fequ8V
orl0LuA7lh7+NXweB7grtuHKWXGWh3rOiVwUaRGNWxQ=
`protect END_PROTECTED
