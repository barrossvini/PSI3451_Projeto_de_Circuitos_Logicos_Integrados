`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lf+ONJohvon1Aihf8KRUaRWS/068uxU2BELXinJWtL4DP20FeWtaUf7Ye1Kh1KXh
XKLUzJgz64JPQkM/zueOyXFLfJMcJXk2PQeRI3f+DMDieztX4r+tyjTEfkyNxZhY
gQvllJL+w7CPArcqm0E9wf8GPqPiOhpDB+XrUU4Q6sMZKpldCN83GioPHAehEKyZ
x5mP3/HL46MxbCCsPMcseG0zHqYFrUfLn3/ij+NnzS+4a6WET4XdaT0y6aaHdd4I
UystJ1tcChwyZAtVILDTsM2AVH+g40r92uZmBz9Tktpi/oumQ1WQAoqTr+nP7SEm
GzOStSzMVWkV/6HsEqp4+iLXMGdcEgOkZZsZle7EB6FtxXmtlQIDy0C+L6v/Tn31
rH0EZmJ3b4NbOpFpOwfmYAxgDrFiAu9Irr7TuI17v/PJIdfn0TqS4IQrRKw6zn5N
QU33StedtsU4tQj1fYEKrxPmMGpRIWT9n+4NGXKUA2IJPBhdptMJqlGmngsdmdyN
4X9UcJGEgnjDQqTM6x8hxkYS0ybFR5eiYcyEdHl8mpuPy6lcH/BTBCCYRIY/67wq
dWhKbKVrmsyBP52IaW8hW0XxximZulDUw5t5zPFvAJQrDL+8EkZa1D1elraLt/uM
QdAZ0YWPxZsFMrtGf/WUJrEjRS6p4EDXXbHgcObDTJ1dREqqU3ZNsiNqcRdtF12b
6oEwfZo1nSArENbsrkiuw7lk0k11+qry5JL/a05pO4BCjOZaSwv0UvHT6RYkOg6x
kZMTIB/0fg1NmtHsIj7XRGo5n8uCWB6JKvkPUis3TZy41ORtlN/vNos5MG8hphtN
PQmdiP+cAgpW+yQ4VRinzV8M0f4iG+3zX/xE82SAcBIENyTdfZUydWCol0AQD0Hf
7+ySbpgyNN6pe6iFbza/Bfd/Us0av4HYjyNyQ9y1FEmi/td3LOkzAyRLQoZTEDdD
PJh57Dy2M2zossBCOCO3zUK3pNZYm3DWYW3i9KJiKzpjdOuWrkKgx+vkRviw42nZ
6ZnRk+eFJTjF0fZLQMp7qBR5Ividr7smvzQk6mE8OxE9kiDu4QEIfNWy5eHG5Eq+
L3BB4RWo0rp9IVk/pNfZad9bWnNVviVxSGhefDoU+xx3JXC+6RwuygmDpjBi03AP
BV8AC2FHxRypJyrYi89w/xI5jYLQ4yFAJQTrV+KziWcKnsrAi4PkEo/B4ILG7af6
wAQ4M1a/GdHAhH2tvFupSnkZXA+ggqnk2LkY2COA8TVg/6pzGgp0ikDnoJGkg47N
RN7B/VMtQADRGr3XtNOZ+rSh1ZgyFbQ51POFdqcDWLHj7ZmHULbksmhVvE8gFC+6
QaoDJfhk/OFqZEq6TQT6e+au1XrVSHntzSJg6ZfUpGRfm2pzDzIlRU+yQyiOkPK4
x0KE091Qsw2F0yMZVVwpLWEhziP53J5taMZQEGlZekoWW4CDwxg2YCEfGkotoKoP
JZzYgFo0B/89zPXJYDBrxEuZE0pSs9yIcGUetg61NzErhZpkE1Z9JYKEdDDfgIvR
q6/wVYWwECjfT6+7KTdMd9QlIk2NRlFqiJERy3gl8ZEnpqLzj5XoYBrnjMEoa3YS
nZY+Lo/v532HbsBjCzoh3ThyeR0fjC+/ZWYsT26wS7MW5heuCe45CZBBYiCA3jOq
OSUXKcx3fa0HMYfGwSKTTZU4Xx6esBimKcJMt1tPm9w42LlMGiAw7tikwYNHdkk2
c95vYejRHQ6XY4/w9dbJoGq7XzITu46vwvEKwrHmcYtkAC4gmLUK/OqTrm5yYy3H
`protect END_PROTECTED
