`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3lLJvayf96Ql0XwlMZPYiQHS4q+D9g8lFb+WF5Zo6bL/AZ23olsOmcvofUgOUEfb
jxutXIgfJ8sBRoLmaHo6HiLEH/LeDZFT1CQT78ZmRnL5qwtWqzr1Drnr2THI1jAB
5vbnQwnAc3xfTgpZ5RM/0/IVgyF2G3pKmHOxAWRk4mAnnoMhkwNUWpxTe4GaNLVz
s2LPPQGpk997YxyK106ChOeobwDd3c6s3ri2c8mxfPgTP+cpy2HCfcGjunYSDXA7
uxJpWlzrCTGemTY41npe8kx71nUPDEQKaCQw3Fpf74oWMzLri4jUySSWdGk0acSa
BHNWhdarOo2bAqhgw7XELxK7JiQrWM+MCMnyCJ/PLlL2FbCwMZ/vd611D+4y/8rE
4z69geJXPQwOJoxXrc1X/tA03e2gly7MJXD/Be2z0xxu+iKRuNaaT/x8qgAiqrtr
hR01gXnQjzqeV29ABtHoL1ZOcLVPkRFcobvLHURrk9+g4v1/PAIC+UqOoI1v/8BY
jaWmE2LnZM2seSnqfRprY5PG7nFHx/+0lLUzVKE3nDmgZUKwHLAoLG0Flumtrw88
3qXMYaH6pKHagyNUoCZzSr1dxjnzDJg9D0MwXAQPk7x4a+58a13b9BXEH2RY2F3G
K/WBwp4+Ghjex51yc+2etvSLh9Qynr4HMhB2HQk3em/JC0xX18eXv8xPXOk2qXEm
us7MKTOTwYnOsZxgqbQNOGllpU0ewIVoStHf3kGz1gRNQoWm8rNbD3dkSVcjg3Jg
jj5DaUicHZQkGjcDuWSaO3eGdfP/BuSTpfteHubPvM70JHfowRdokwglZ1s8y+8m
ydtKi0hqVoNIhSV5CuiRtAo3sfHf8jOdID4a0J0pl63mM71d6cIECGDVxnuqCjgI
`protect END_PROTECTED
