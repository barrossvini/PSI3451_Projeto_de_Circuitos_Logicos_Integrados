`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oJdm2Q0kk+4HhuD96Od6jcToGxdaJTlySmYNcDa9GKjgODO8JzPNNliOv1/csGYB
YV8+GN26XnizMHTPF7EfP+o+/jB0k85dIqhfmmiSpC9Xyy739bHYSQoyE7GV4iOF
zBuI1mgtT6QrF4wrRptvnjyygabAs4TYw/foHO7/jwF3JlcGo22Kwbc0ziyVwPA4
43f9SPT47G2kp7AqJsyPgBIZm9bzEF/q6RFrEL2LYWqGwQNYEBfnQBQWgY66ud7C
qlXqSEszqQWOxa2iV/Jaw4VK6Ce82VJYU+K6h+cMlcMmLo9aEcvw8LW5jejS8AAy
Tpa02sggrIbLS586GAvGGEubufzV6TAZ71SP0yG2g06eWv8cCs622kwOAkFVOQqO
k32wnJgOxDK3yj09C3ZyERxSOZVdrBe0iiYe1MOxQthWqdneOtyFfd4fKAXHARQp
lryQ0jpybMBRbCth2gsjs2q1Mf3/aLqldSoAwQ4HCXnFUpnwMXe9OcLGVqyg//MX
15L+rQEw6pDm2a+HxOojpP3U0dO5Y6MWzKDwRnDc79zm3jxM/SKkvwqiKK/aVgiJ
8Bb1181aLpFJHdnZ9+DOMoiwIO1foIquKzjuUrRfAnXNYMJdA/85NN0vmHguA9L9
OgsNiTmWiSNejE8a11izMb67WaF9mHXc8e3TR97gcXrcluYkmufabjKQ1456/GJd
/YkBr/SQF0M3Bc4vwk/eZ0/s3oay5VEYttYJHGdVECsWcAI7aTgJzLEiFmJtlQRo
kL77crjL7hIx3pTvwwVjnq4Jr8rywK/OohrJxp66VjncEwMC6IQ4jZ62Su5nbqke
dhHu2nYnoyK7VvugRU/DyjL2PFrLQjj5mDUF03YFZiaRS0LlPnaHhm+KMz/Qe9M3
w5zT+0HJSE5xbtS9loccjfG5rJvQgAf+qKuldm7qy0KiOyFTjDNV0bJY5hgXo4oY
RkaRb3tjkuXhpOsWK6IJZhx/X3UjNe8eZzr3M+4oCiHUy8oDXAbYsDsRsjL9syN9
Zc4Mf9Wc5ILRPbgR/CnhAUU+QcedxzuCQpfmZ4zZw8oPBcDKI/Z/w3l8TMpoyNe+
bCJ1dgDpbxmGZNA00CKaFRzDBQqJkH4huH+qB5F25DDCJ16YgKO+UMu+XpRa5pMF
c9I7O9cEH0/1bhTAWZ+OlaHAmDmq6eJfB7EHy/SUMkBkyvmJGcd3p2jFIz+rxk12
K/v4afUu7LJ9rZd0mc/aNyUVUZh+/a7MkMee3OMhRWftmyBgUE5Hp04cFr8aKCID
JT8PyqYj//b6g9S47Ysy1/mg3v3K2TPVvuEs+lEsZj4zFLoY4KnJU4f3IaX3YCzs
jTjm3izdXU/8isk7j0n1URdtupLyoJVMmRgAyhUnxzNup+3u9/HbDlQ3HIDplD0T
7zBoqceP8pF1JquvcH2N27M/ml2XSP0Fna9jF4sW/2InEA+Cngplosy/8DhulWX3
PO3frXy2fDtOYfNUXaOMAtMjCLIFKml1idAJXha7VEueEJv75bNKyBXJ/0bdaCfv
+4WpYppYcWDaVmMVIF2z8U6Qc72Z+KFMUQ6lnR9xY087ZL4EK5Flnpfc7i6NBPa3
1Ki1PB5KdKtHDTJ0oEHubRHaI1Rq10CWU6+MZGyiEgAFqs9M69M0HVYRuGKjbzk2
pWzXPd6lWqEVAqoPyKCDnmCjULttye+iFJjTBljfswEmWofUhKDq4rYvUKO3cf2D
HPHeLBnk+J64lIbRgo5H0v5we8VnvXkC6okJOasdsQrwRJyiuY1NjLBT++t+y6N2
Pa9XX9Nybsd7WU7Zmq1VuxmZfglFgXPHdKTtGbSwpuRP/Oow47466t5lCyyYSmrg
p2bNZ2ElaMSIef7oGZuS51M07AZr6L8lJzP3dgJqsRVa+zFProQTXOF8oQaIkd2V
x+ik4E6h1z6TCJN6WHcCRPtjPFt4tCWJg9bykAv4bWBbnJN/EkbSZGpKiKvcEbyl
rixzZVxBF69qx+dAkW495fz1I5juQjS0sY5jy2yxafJGWpANoASbOkWTYdRppOPI
FAbWBN4hGfttbBgpxUjll4/Uvi9+g0k9VQ7dlWceL4jqhczyI7VHRs7NzrQE+xlH
jTiKqLEB3+ttFqF43Z1u6wuHs75+KPxeEN19cdHT2VxnmcFbRSU99w9ZUIc4dgB2
rHKa1e7bd4Owb/pKCn9XUmjm3CQFFqQMqb2VH+IAovloj0uG03BLhFMjOxzO+aXM
LAQoDDaM2JCCNDoQuyT/pdAy9NyXA2X+8Hu9cXhx2udQwsoSvw+u+LCHwtw8AGmk
PgAssMdK5GTTidDZpBu6veA+Tu3usEkf5SUOWaoEvwfSBEBDPK52PJbVnvSIhz9W
z/wVPN6MRDiM8GdadW4GBoIS3ovwpAi3Kl5RPXvTWLNgvjzPq7lfujTQZp1aC0Rn
TKSoVVAKff3BtNl0tTBqriH9u6JK3V1HFKHMHi4xmGUf0sq6eEoakGKbGtwG9/zu
IsEZVb7l4kjtuJRGwpD5sXMx+f07T0PqCwoS4uBO6MCshKWA0VZ37ERb1dywYjtD
eTLIklUB9suY8xzdX40QtVld2QUs98QB8WMTj2PRWNJdCGLtRHZSJvUfA8J3DPGA
0aJvpqkQGsGY9nyOkP466TkLn0S6TgyRq4ulBpWdyeMMQEZGE6ucWxZf99Unxa8S
ER0KO50ajhj04bXxgTEXrpRjHQ9IJAL2t9IpS65NppuaeogxJF9UR1u2zAR+zz/G
OhUkCESQH0wGbnS6W2IOxuNrGLVrgni7rHquxvp/VFaSsLicxpYdyCm1DU6L9CKy
sxPUGJQK5sjRWMrG2iX60KTLmUXcDqoF1lHKd9fEWOAebcMrNEn3M65IseIfRVSq
1hQWo2Me0wqeSA5aZDywBFGftt+NHwL/0lumYU8Xi3Njds8j9mvz2SMU0g0rPSd9
T68Wz4nzV2fraWEeB06eO1mKEXGDBYcmC0s7qF1KI2vJz9HLmdjubXW7FDSMobEB
8ed1VnDvrKtKOFsFurzk21gntTuyWfqF+i5djWuv6KL7/+3ZBiVJhv13Q8sGBVr8
AyscPb9tP+yDPseog9iSM7XsAn7NCzeQbzMWnrBL27ek3oIAULwl0eojBCHfCabW
cDBKstNYiWSf8KZ31Fl5XxtmvVZnoRvoy95oHJLLVpm3x35k4MnzTLQ8etHAQBAA
WF6OzQvyA4Go8YQfulobh9gYfnGR651/B6BKiM15CQtknYk99S2935oKqoDF59dP
7nDqxJt/OSg7m9U+/y45+ctlz7PIwDjRuzzIN/QowYHMqdIloqCPKQ03jHKH829H
d9BveP2+vMmF/l03hKxHoAv1AV5ZUxtmjFUKHowHpVx5NmBySGUzdBm88yHzEuuE
yUKNMTjNkE4fCzRLcGCseNG6Hjn2evRd08HxxEg5glhwL7m59e4w6Vv28jz6mpq9
cb4TtiIiYia5YvAPuSEcmpcBpNuS0WQ66Tm2dAvUdcp5G/ybm4lvlVIGvtvQvhs7
JzIkvZ88EcY2lV+hBcg+46SLmKcPfkF7PfebxaWcjvf8wc6gWIxsJaj4gkZyCTT4
ons3LYyis7rG6pxBL0XpNX+3THojviqgLPAi34EOsFCz3TmlqZCQ5ihC+2U6EBXg
Uic6A9mcCPcxjKfLIHCo79jVqxEXLOyU8M0ZUrsyYAW4lIKDCJZ2Gf5awb7WoMAJ
co1EgWhnW3FCF5Gomkwk/WnH2+qM/wHlTbhILwwrcmC+Jp+bpMU0krjTlRTNuzUg
CXlMDUx212KGbFPB09qTFes6YVRp4ctdh2xGRJ+EV8OTOVCYG5QxP40WFTgalljr
XSDX6kZeYtj9awNjOqiQ0wbOzK1gL0S5nvDwu8qCuobw2FSZkY7LHPxb+M0eyXNW
hXcV+M9ZBjXHUIUm2cMbHjAUjlBBWMyIDiA5Izv5TSq5zT/aKq/2b6jSMrIW52mW
ULktNn/qzNeq7fZr/KvzzlnGZgYTBZAF8gBqBLvGecO8bq+gpO6x5oyBrgtBLmFA
rSWJrxVkJ6/609VKAclXa9vTf+l0JKw6kPI2YE5JMF5PVSO+F2fG8tDdf2BeZJzJ
Oa4AKinklakOWLl1hvZooTS578a+/62U8rXTXA10i/YdmtJwdH2HZDf7piX1GMhq
OPB2R1aKmdoY0rhZTcMlbc2DhBH/A8Skl0EmJAfMAgby948Fqzrj814JfTiAF4nn
xSQtmE1+rdWnKAruRTAOULkC2m++VGWLOLedpx+AV8wjFfibKJaWuiWa67wx0ZZD
ckFgCaNzQPytf9vmFZ/WG4ADShdil6YPLXqb/dIgjbJdsFAW/RYYNsWko52qotJ9
YpkEwjw0+PLndw5rSjlSUFWSSe4UcGyDOa5jcKLHk3FOuxRqTgJdIVUufoV9Ah+F
5mJtcdW8705D2MrsIiK6lLfkCtd00UsTiJL04EZXL6vPuZo9ptvEW9yDDlJS3//q
FCWChNyJlZeTFmRhRSLUJxfUwK/LBXceYESlSXzrOl7G4mFPWzKnSjGbee0h1z4l
DIsi9aNM47Rva1ReUERhM7TeibMdkBC0NkcUsP6PSxxwMiE6hNoluSp2usFsWtOe
lwz6xmlr638clEClcJWGV8+ch5sVZJ5irfSuYQZ1meBoNuEgV4BzskP4ThQ+0x4r
Ucs5+wgYad7kWMiRyFJAMoJAwRw4li971xjHE5nvmpyBr1B815LKOgf1h20T2aOL
8IiZ/ip47+Tyere+kGfdU6W5kS1pf7L1o3dFGmXpQjaeWnLfUxSr7Pyw2XRtPWUk
AqTL8l7rn11BfL37vtimoLz4KdTU/lJbTMXEPIVqYTein6gZRafXUHeSWYyiGPm0
6I75jtUWL1SR559w5dff60JR3nx6i5aN9u1gvjE1Oqql85vIqyWj36qc8snf5VM1
73o5376/JyNeP+5CM6HdB4T3ypM5O4YHvVz/+mXJxAeKZEB7eZZcRJq8A59TPwhz
cXfaXFioEVQMfVZWPKx3kRVTeNxvdmUVIe5KHChyRkg3dvv1KMGsaC/HW8f9amjf
kmOfOWQm9Oyp7AE4o8KPOF7BGkByn31X9wNuSDOU8RUAunxCHJHxXnojfN9sCTJG
qEvhndPs/VkJyag+IJLNy9i9rVb+Di+JoLLcyFQnY5S/+NyYeyfXKPHyBHB7YMss
1qgPuntZTunVB1UPI9cEAkpsQ04QtdBQqqTC4312Cgd++pbW0NimGgCpe3Lzi9E/
yA8M6sbnmA2Prie2ustC8lnP4h5EbtqSYsdEFzw9BXDldniW68sZmHUjg23sjLb8
KEbxm/Nh15OjooeXZpd4oRn8Zx+AOSdCMGq7tWsF2WzgBuF7kRxR2A+sxPVYg1ps
1mruntSL1VUUwvX6pT89qmz8/eqol7va09WsnlCAmjSoTGELjasUqBrNqI/eoLHr
b7Ex4fN+ahwqtHHoA+JESRvnutn153svAL1wdc7C/EWF2f8UsNeREHR+YI+YUvdV
aCP96UwYwPcr9BGBGJDOEALiWsf3s4PZfZCPRTvtnSJjciCSJck5mAlmtmbINbSG
oh7+6Tjse0y89HG+cVLueuSKrEfUJvcym2nbOYZ3eYhOqP7eET1VmkxavD6WugZX
uO0vu6IC0O9Vo6pQ3BLU3V8+Ob4R+VeQ9XdL5KfTjGKFesrCaOwYUY6a0i900L1b
LmUfNvF74sdbBs5572ce16pr9v9deI8mHyfl4nR0BtIB2hI+RK7Dr2CzILhsyPNp
Hbx4GfgjANScVi2xACEXowfXD9T1ZOa5j1hIGgaoBwn14jJPZhoA4AP68P/rj6vr
4IG267dpHVbR+FSC/5wv5hEzyzBj3qSvXsG2Exuu/c/jv/D7JGsLfS61Jp66SNH1
KzyBwfdv03o0QGqDyeuNY5fY3wjSbpfgO/uigNzFIijDNkeOAGWlvXMzTKiVCRhT
csT6hLigTSK7StamUK2JnGxO1AK/ATxnZLSNm6hl3nYyrZz9OhZQu7p6PUD2l7QT
kgmjslRFStVMwTRFl17bbwZx6Kl7YgZRjELEEw3TRs8JgpWKX4eDX9yccJWCalUQ
+jJIH8lD9L/dJJ9wmUTzq9DLkls5lJEj52Hpn5AB+FFtwP/7aUeIvkT5hCTgczLf
4WH+5ZAqoqMl5IFXohEFrwfTuDtAu0NTIqIlnFTZCbtbvUfCE/OWRoTqwj/tXc1n
NrVQUgJJ5JkrRXABwNpq6ref0h+KqK9Ak1AYaBftDJj1vvqPbMWV/4tsMllmJblX
l1AjYHTEKBG0TTBdRbOg7UIbEmb++hyNfOfQqF6QUUqo7srNZXASZ8jKRJR3Hwkr
Sg0IF3BRtfcssKWVogJsQBR7da/nF9mQ7etesGkrbHZ1SOpqVqhzb/84vdmTzTlP
xg+JX693QLPDUkHlhjGpPILTZKCLrR+f3XeAnveW4WqkXEDZZr+u2XLOdHX2Mv7W
+KyEYrZaFwjGpKPVKY2xxDoSr+zNsEwiyvSzcez2KlBGCHJMuu8U7mIE9ssXugzv
DQwAdx80zc4uP7tQnK1eB/5uZuVMqLMG8yG2YfWFaRZJkKmeb3UouzTBX9kPvIAs
E7jf1whThikumSoeoEPjYVJQQ1n9ugG2l1RwtHjsiFkPRQurB2/GBWUf/9oUB9oU
EGKgPVaJpwbHjRPgZsPBS2uV/Pp7vNRQ/a1lO4QVgq9HWIcGiWea9Ss2qwUrx455
wl0/Mcrm/MLizwXGFfZtH9C/dAERREmdvH629t9ptpS0vLZhsosmLCwGS9nYGjfS
WBwf9ET7OSwBcj9YGQ4RsOC2TCmZOagtI8skquzU9zydhJTCTqclMPO+5H0cpzPN
uSBblTSyaR2IgaB2ezAMlZRcOoTeBMt6TMct0XdsnsltrqMuxlUZjURI+0g7n1aE
Mq1bdqwOlebSFeIoY1tQE3REdBzLBu2uEIqd8MTl1xd/ZmidC6DsY85wFS90udzH
P54A8rU5tiV2aosk+o/X5A0GVGzSrZR6vMl8XHrQWYX4v8U4WkyfKz7RzLdq8PdK
J7UGD+bXTWSHbSCUCccx8PjIX9TSYV8b4WHmRff+PuOG+gDdi7s/F1wE3fy1tUFc
9Ro+qeRykOuOCKFX07+tMgwCYIHBciy/9zjJpvr+J9WRMBzQpkY9ONRGBFR0NTll
8KyzEyxfBFLkMMImz7ka0AuP+vIPk6qeM164+FSThgfHQrA48EDmFbAFTJ+vnYVS
Zu1vIhTHG9kYWsYIpYf+tsyVHJM/eIy2T3ekxKIzVtwhC6spMgN9PxnzyKWLuvjz
NJocNyyW3K5ql6xPWJqfTZkEwFBjxDxHiVNP+Kf39qHsyssVySm98JCwA+pwGX0+
40IRS4LZDH9d5UZyzUwTpduuZD75eDDsSNaFKVMnaii1G029HbHyBr+qfGNs2C20
70OeY1GvcbazKF66g15HLAvQOmT7mEF4YMkmtgHo5jpSrlKs3DP3jdv/OX3FYnUy
3IGm+5/G2bx3TgH8/aRUniazw1frbNk54XM4X4QDTrbWq+FwwdJwX7LV3q7tnUDN
RcuS4eIF7jBaiiakGKaMrvUBFN/8FV4SlIG6cEem2DI9fOrau3VqnK0ByH5QVMza
cqTePRU+FDx7+PH6dOAgQxf5EGr11UYxYBCRQ83SJFVhxU+vEZNCPpzFmMuwTziW
OhX2CX5z7Fhg63VHN/cGphT6iHqGbgqgkHKWxBgbQR39v2X11yT3qfsSqT/uysjY
yHfjBCmdB5K66AkHF0egTiScwgsSG/i7+7sS1M7BSDCDINswjF4ZZJjym+hy1G53
mA+xIEfLtzD9GISPmX8UEkcC8zlRjwEgHiteSrs/G05XCg9S0V0QSxzmhLCMosWk
ImifyqfUrnGIppeTRPwMqoacfWcsyg+qTIp1nxXeRzV79zKY8fmmXWclNzQ1PZ07
JQsa8+ios0IapFF945g7YZd/V6YnezxvjOLc9a4zU3QPDt1EUXRoinu431CMOWeo
72pIyILSKlG+N036mfHm8oRptHi1m3Bike+2XG0pB6LCVHean4H9ilrY05wF/77s
I+m3hBRJEoOI83cQh8E2BhpOioDntE0wNsnmMYltaWNGiTbbByxI9l/Hv/EZZXL4
vsNGU07FfS6sDgZ8SG3C/gCvN0sQljxxcbG/9XQy5qOR/FKAiLU60wdwZcSYC8pU
ip+xns+/e8mnTWT93mGr3adx+bVIA0R83qrMIPsSthPvlmCnqXDCXjm+h/kvOGgx
RDtn5Sb8nrApv88HGUCosu4h7XiSlS94Yf3M+HaMAgDuN9HDlV7tPuIqL2uy/Tr2
18RoT3pZ/9ziIiIle1aRK+WomZTPW62u87yFQ9vMKfYa5EiOEuAXWbnaF2uVn3mM
lZeU1pnKd2Ydb0za0d0YgrT/Xu+buZZjEYxU7EQc7Q5nNA/TFEmcV2fTWAVfVPeM
u48bouEz1/PMtqgNK70M6yNLAzVEOIBR28Z3DmAiwqjlQKiRwLVYmY72oG04ptS+
4uRAC0tnUfwkZPcW+3AcYar0z2YlAbeN7zpNRRBi55ZvbZbp1Y3fc13gFBsZm76P
TMKGZ2/BwzQh1COmEV7ttFy/YlZp3/xMcB/dCIkOWxuLM/Dlx1ND33BfHnoSpBdN
znHspG/507Ak/0SilpcZjkrcdhFSvV4y7bFYULVZTD7HGkTS6LkO4krgdAjxcg0a
KsNMkODKqs9qbJ7yT132ZC2/DHj86aDpL94GI1IlTI1ls0pldt5kScu3PV/LdIeK
RwYVtIR45qosli9iNp17LtQwMnbQ3CDBh6TmenHFCqqbue95jBm/8D1n+5CjZQXF
Sx8BRjf5ixfVJKhfjJP4iSkHtDcCdHXiGdG5Cplm5coraCWX5xuCHwRURaVhmxDs
SVAs6htPU//jMsyHZod+rgeDMNXM+6FYEgVJOaqFRR7cqnbt2HJRsr/yXDfyvitK
N9i5RgqQkLLkIbFgRimBkQ+6pGj2CjUoK060oOLM0wdh0GUoEsl8t1rJBijXuDZD
dDEYoAhKHuO0gE9xVOku8VztgrCviyxJMj5uTKkNfqS6aD8SIQdcBCL+9O3zAOLy
j4nVJABzxEgsfwfeCbl1+P+J2Pv8nJK+0GH7ks89nFynt3AtpW9uWwfYhd73L74P
7+2Fya5YD0+L2Z6XA4PTTgxg5c+mPRb+Xf0hup43MomnK9fpUU+hHRBHD9lanxCH
GvAEuSPgC9gjnh6abQExQFreIIF73JqN8Vci5TAZnekQkGge10ILA/F8pUBtR5Wm
NZKSrUIiw2YlrHeY1ULcN2jiIfyuqQ6YwFCuhX3hOEHMU/es/lImH3k0PRRZlx9V
CoEZx5Ag5RFI/WMijjd373liB9/uJTpfoF+cuOmuy+EUTI8BfzwvgaHCPdrk5Kl8
ItzF+nouoF5Dw9MiaBdTpCwWqg15/UahnFEs+xMyuvjpBEw2AU2dE1kUBCHrdLeS
5Ob2bXt71Yl5p3ggQFzg7uBryyL7zA4mxDaVySSjLagHohdZiajX3qQc5PHypxGZ
433So2dtvwDCWRqUmdhZ2fOok6B5Y8jOqaWQ4gXTZfHXDT1PFczEza4l1elE0B+M
F/nUMG/Um8NhXnlES7VvXvqFgB40a0lIbapOpkTW/xHwvtdpYd4gPABWiM8xb+N4
MPq7PiWu7CAtD4Y4jvRTKlDtZl65ZDeQXk4giHDmx8vSpnree+lrZRo8LvVN0P1z
0LLhQIpqAAZ05w9187J78XECIQG9+OWEsU0Sh7Yj37rIrSuyN30gLPv9wVGUUWoU
4aNtSmq6h9hMbYR748FR9hTC3bAArUntSI8NCMNE30URK4g2SwjOo5ARHfovXW7J
NpoaR24Kxtpo4iKHcAUjK68GOpTJYgvWbubxV86/xyv1UrJXtfIxtWrwBfye2WI1
4gA28KOR19xjQt2EJCmPta3gihVDzYUmkJKkKTKVP7SFDtksCqj4a/5zrUhxMHGU
No6nJj9FIbQvESfng8yOdhbkzMk43BxoRVsFLOb8tXgJ/t2tEqVLvEQTZAs81J3c
2cp+aLlUhqKr5GiKfwHk3uJWnso1P6KCIO9tO3P8nINMg+CEY1RnKVXxuKhiNFyp
j51sexwTtjIwKOu0Vy5TbKy+pEAki+Yqg9vL+VpUK6rRDInNnwMhG04De6HYT3uv
jsrsijxUGPjDktb6UO4Hunr3WhslFSGMDmMmGAtuphboTcr3OEJtjS3RULIAsYed
4z9RQ4l+DPwYs/1eJj3F54UIcdiNDTIPeCOzu/MI89BVYLedXJWxwX7xqklkEUJD
q2iLzIg3LCz5csUVaiV6/EGsiy+w58XLkGoa4DOamFGlpXxJlfAoy3qY6RZOxqzB
kX+kW2YciaVgGWzUDe5Syp6kLp4rV4nPwU3V+BzYvzqHl8G7aFZAIPgeAzvNKRJ5
FvhSq+7rxomQiPzGBibDrj0bBwdh0YgF1o7J+laOde6MjofcCrkdpuDbYecKBshP
GYlXU3N6kOH92KgkY+tiAEyZv6ooG1ZotL11sBeTTO4HPdxxJSdUO2J6jT4YkY+4
VSWrnCHIJ+Ip+6CwK9YPxnYPerxdgjqiEdlBBcYkmh6odSqtvX6Ato8g4Lr+ZFpV
5BAoDMI5rmo+AOR5BtF/uM5fAQyHLw3et7xY6K8jrPPNjWDUwVawHQbQM2P+9bGX
W6NL9Cos48/NE9gJojpNEK3a91LYMSB0Nl1eGimlWd3f93oqvBekhFH0oO4kEeR6
P8VIpn3ymxrCeAZEu0tWqXxTpIDmc5eo+Rud7UFk8msfUSYGRnDvUn+Hv3ffDtwI
GA2yZBxJMi3I0cztre/QE9qUHYm9sTgITYpGA1uIBwpyY13qn6bJgk7ogaLZXjfu
6WNLK+6fe/UW0bNin9cu2Mg6gu4Q9tk6TCc0KaljUS9V9aaQ7DMPqvAG/ii8sJ9+
NzBo5z+n8IuiWbVXLtMvkxXogJp2flLNtPAJh8dualKDkiX+GSyB8HPeOsJ52/Ko
13Gz0ucSRZ/SGSVjsSSgVG0iaObOMfIDGB79SFzB/NKxV1iGa8iWDW3WPofPMeMn
fe0pVmjEyNoJnDGkGC4CX8TMcPgwpNxCzLkPLh9dUgNazi4IYl641RhIyBXc8EZR
1TvOY2ttJa8196IeipFKuYOR+MvIgOPT2AJv+Zd54PgZDo4dq3PK0zPy/J9MHRjn
jibDlyR79PWzOgeoQ6VspGHiFai/+j8XCjcQ4MdNZ0T4B7913OHjHuUrLTonB0RU
AjuvtdkZ/ngeB0FF1wUtEU3ErauQViFcUireQMQf53cLN5IDpeSjVesLXt3qrhrK
1Olqgw6JmG4xttoP8lC5uemfS3lo8W6NjxvPjCbpvD7S001CQhVWZJf+dIxYBdkk
Ps0fX7BX+PyZTYdiQiOSDt3WELR/v2FsPynq9Vmx1g/5BGI3uitb+he18rfb/Xo0
NCcywCg1GGPGciKBLr/0/4QUPVfyQPiSOz0gzNFaSGX41Q8RagRLEugW4nFyBQdy
oXaBs4F7oNFx5XkeasNOTZy9RH4evO3wQIp5AJJQLoZ72YKpivkALURL/xvDu9vc
Q5SJ2ncYnGY/R1n1PE5GmnTmFvgER8psBu6v2YtZvrLaanLmTOug4BFN5XqDva+b
PFptVuI9ZVl3O98Nw3q+vdUEypHXzcFsv3B+D52YCsYUeE3FJHEB+IPj6a6BxaXL
Ff8Saq2MBEqrxJAPbljUIcR/9biyx9VesVBIN/1tHTbLYroEnFJaxP5ZHPGTT7du
cVC+CdAbik6tbAeZvm6qTuq5P5bV9WttT+iAbIfcmJLpNKETXJ70BDE86odt9wwL
PM8BNX61dVPkjJfzUxzLhNoD0j+blu7G+RWaQm9CkG4ycuEco2q3RIYvrKVxgNhR
6i0j8H3RTWD+SToJ7eMUoCw2S1VUXyfaSGSh4ilAPXeOIOCkqDoIcIryJjC0+pCX
8LEnpYJtumRcSd5xwQhz6d1gvHBJ8WcPzCdq89F8MRaKlGuI5YK2Tp6NzefaAyta
2oNd0+PcF/LdHyK2y4NTx6BvwshT6IfOp+pw36FIIWwsl1nt2kv4GwvtmwBhV3Nl
HcVy8NhMCYLHTXU2lsgFRPT2ChusqYvjXIqQvynzewdq5DQVh4rdkrTVtU1RTc8R
+RP+d2Prv2cjImEUnZh4mn/Jd4d1jNOFkxowRjOLqez+HzntQhFpvfd8AIUopaSQ
slWof6+49+RtUz27UtHMAivuD7vFSdEZcVDpevUN54Q8+L2UGrZe0m65V6UTsSZU
tDiBpvOF7H4hWQrEzmpT58sacW7KG184tIZKxcuGoEq7vs3Lz+zRCrDj8s6xR0ow
+9ELnq2X57MIPR32jQChDG5FHWxYHX2FgoRXGdT73sRzfgAIF/U8yoJq9G/VCC6W
8Up88Jk9gIFxrgtbaZ0nPq/G21RUy0pH9gbJMbnw9zEn+nQda65UXBonZ2WkEICU
ob619ScazjjDZEC3IeCtiO9s8YzDtOs0GF3FcqQC0DKynI/jQsKm+2PdlbFTyjeY
nAkHhIfX+f5ozfJryw2w21Iaddlfou6gLM0UHSqchthOSpRHcRPeDGMTje8+iyU+
+/oA+BxHoXxkEpfQS1mZuSWvN7yLdtNG3g6fY9UqF2VMnWykweme1vxR3A82Mr/w
sSziO/t7mMl5x4dgZAwzZLmHGkjYuzsWGz51Qo8gnICvL96Ppm5ISpmrRyKiaiPN
skzJHOtaT6bfktlsp8IPjWvS5A34hJBR8V8ZoqWjSgfacyeJwz6J5o7aci78kFpC
lsmAWl/XO1oYUxXSdhQkxe6oNj4fKK5EnMAfIFAFlaBjbVOWBE5jcKm4jAT+WFTd
D1kgdfyy4JiGstd29dPPggtyqezsE70Hgmz4z2ow3mPs2eTDw+ttNabt40EJGdfX
4nBBejGvQtUAZEX6tb3QfTvPhC3eNWtYQETL4VDSbgBtaSy0UEm+FDYvHqfh+Kvv
AxAEz7EWyn4s9dGmhLzU8cn0jnLY4p9ilfv9/P9Tm5a7ODhuluNGe3FNTxI1JGEx
7ybH7XfUB7lPwmLwTZXZCBBWfWg3RDmmygiEKOCW9HFKNfUwogjNqWyyBK+ARVuo
HtGAvCwd8F/JBhbNyQ+Pamkr7wrbMZAzif36kXFxQIeTJYQG5PqLlVta6y6Xnct/
UrPP4hLxx/svoGCoKZWG8IGKwJ1YPbYqkSGtY+hP8o2Vn8Y8iNRzBrnhy00rshHj
b7Ifj7AXWc50fRwOXMwkByljGCYIkaj+wk0Hs579JZyinrHoRbgZaPwwF/ZcI1T5
HGqON4NTdHtSbDVIjTDlc60KccyBuEzG7dIu5Hmb8Gx8uiOrz4G16JDt4zjf1ZhO
M2GArkzyIk05S3VRdvQ53UGmg8WkWvlueNgxEBMMeUy0t9ffwIBBLoVcxyLlTOKz
dNukSdA2zNUzdyRL6D8TtOv5yvEM5LniDv03RXHq8e/HykavGkwgwz6xDBi+G+rJ
dNemJDll72HV575ru/bHqeppDqkEEZbduUBmvKGx0U3ZmFyuOefoPpVUwSvUQyw3
UOLRRGO+Vwhq9bhSx/VgAcpld7u3bPaIqDQvhM4e7fYkcDbjuK87dliJ6HHSY/6u
ABvCLa4J4ucpmauEwY/Zi0H6P772vgrdKKQtSs2iTPaFjX82BJTG1XiX/mFWiGQh
kU/SFG3dXxoEzDmi6N6MCRyE1LhzCIaXqMZFQQ0qJaxs0ERxkOzv/QT1JYD+0dXX
L8kubP+P5VrS9v2Tjwp0q0NZ0fJY7XDB3jFWz+0/3zykqlz/0BtuIgUl4z4oXd6B
UsYYf2RQoEyoihktNRmEa9ZQxIK5grgUPEA0EV9vj0g7sW4JUltLmCQZxvWKvc5b
eGkgHAliPQSMKkDVk8T4HRJZu2upSuH/1blG58oZYMYylNFoP2dQQShdVLFf8i6U
nl0z2ySrBtor25eMAr4XhWm8TRtgXoUT8UFVG4QWsjj2CzNT3PckXoS14zRKJkLT
FyNtdtOyupJ7IhswUyw+6WpuhGX3nixvUBIDrz2Zw3ocffE0dS9st9c/Arp0qAvx
Jx9oxI0YWqNQyemCoznwxHtq2OIvkJDeNIAuRjOIv9soC9EO9hP74ax0LZJNVlsV
RZswQ96uRIqQEZOe1eQlDVEekRl8xAikLB1y9IylsbjMI3tP/kU0cL392Y2TzN1z
hvfYvj/eruuGGXRdhFrK5DgDmZJVuwwH2vfkco7twiuQqiA9eu1Y0I84uGqJ36EW
LgPaXxH3wQEImNqS7/addqcs/RgxrYGQBSSgJuB73eMzGexCS3TLxcpNAl4SAFM9
do+Cz4iqKOgDUESO9rXEMM0SVuTn0oui2ny6EjBRZHxv++X4XCyqrPYQdlQJs+7Z
IrdmE9g68WEWtyIGrz6qwSVokKSjT+43QgJa6uh04xOTkCc1tuhOQg9bnw0NncZx
LiAnrIeeRWTCRZ393MOZDkd/g02+CwQ8NClmmXY+ZojdOTKirCs0Uw7Sq0WUtrm1
IAOlVGSMbRO1SV400XPdtjQa7XP4jG2Z0ouORW/dzGjISEVA4T/FMhoT6GLSA71n
zAg1Jv0R/NaWKo825CZr7TOpLtPIBWuDuCxbFJ8HNiROcnWFru6HlB9KpaLBddGH
OX47RjZBXzObWgLcjHlf3o/biLVntEu2/iiaBBrbaU2byOLEBBz88LbqO9l0mGHV
/BqLWvbA4hnSzO02hzGSD7bCdNEOT88m6lVRtk3XrxdFLuIZdRej6eFsE8girkkM
lzM9umTEhpIu7wMC72pUhxC93Sv8QrogoPApfi4eFlP8ZF5NAKlwXbapC6TR740o
5n4Req6IXGYpWaRa9YhivVuUZ7iwMfg2kpxq59fUawGGicBeotC4FBf7NN8lMn2n
Pu+DR/B2feXnIleFpeZoqoyWVPRp/W21sGueDVCsemC1hrBY1CDoFzkAKZ2FcZA8
mv9p/ZQwnt5x+3N1PPUWWa5sbvLLkZxVhjkKftwIsbuas8FM/XG9kH+YX6xY0ZJI
be2oF6EoaVo02p7b0MmMI9jSnIGUbh519QCkLIAm4UubXO3dJHJEWYViR6s2Gwao
iAE0iAkrX9/h4Wf8Kv0HT95LBgZMwEo/7SZhUDlYfJsO4g4bEiAtMqz2po6KtjFO
Z/tctOruklG2UmLoD9opBfULKJ1XINcuop+ib8u88aQ96RhYObU8qaCWMOfV6uDv
f0WbHZgOtgp7Et03FtuaFAASXFuiVY5KH+ojBVSLUeIT9u1eug/kh6SO3nWeitnq
guAT7LF7w/+XbiLY/DEIaqQ7aV7Aye1znYX4E1A39HpoVM0aYoaFP0p5l8H/eb9b
uieLcO1NFBt9oYD8WmbNRGat3OImHUlX+O9wQ5nKUigspEqKMaRMVlPaAoSGYBup
4tGSqNNNazO7jaF9Fi782KIZUA0aukd38gdGSZIenJKkvFooi4t3Vdebbp4ooMtG
PGnJj89PXLjmHPK0voeNUaA5hbifDgil41+3GfCB5ad4As7aII2Lngvia8MNueTi
vVbzhlubVJCCXmMD1ZOfTSJ6AXnGZWrBJgz+LNoucG7LtHEggiYfm93dZJOhAAP/
9V/xtwg6PQCLVJeY1GVAffxEcIyitZU4Zs7rt76U5bmmL9qhfi4gYLcyVjHGPXGo
4Ufbk14gUFMddXp2816XXAeeCtDAergGWwNTYvhtxl9Q/FhTKKpvo04puII5rmPx
66B9jPgj1nnphh7Ylwt10mnSh44Hd2AJf/jdjNavEnNM5Df6Cas+p3DnOMq2bYV/
lPrS4dXQn8TMN5bs90Tc/AwK++BG+cm+58k7ecZtgcdAVVKAZsuGPbwV1ljIXJHR
0ctTVCaJ+qJPIjOwtTI87egvtZRi3n2ppztlGwGvYFJku6Uy1YsDxVmbdmOGh13z
eFTH8tHLsXkyCjAM/cONy+Bkz0i5hnYeA63COHV1pf4mTpiA1HZmIMaN99BM+/sE
8/fQQeLQWjDV6XSNoUGsWa4WpuP9l2Lh3u9UBhYD5GROB1zovM2PSZw+0eSpEUBc
m6kcttPzVUX6by6UbKRax37RRW5y86o3UEYyTu8Xo1y/SsxAPvxTJisWS4wNVyfp
GNKObcMDmFW89XKiGOkzl90hZIxyhrGo+2CSF08e+u8guTbnSf75e5EM9ntNSQtn
brKsHEorXZcYIA4nzSfEAK6mwWWRRTk4kQmtA3U7iRCT5aEnqXz6xPOMP04dZ9sW
9ykIdquoG6AvfCxMczSwtE/nbyGJ2L62bHP9AQaSbY3jbBFiRC49AIWZLJoB0xHX
9elNNSxwVyaqCiGUm1/LVTlNGBqDJ23Cuync/K7xhP4ZOU3YuS6zKyw7FUwQ8f+C
Q66lruOMyN55pSJSRYMuYaIQQKeIOk3Xy/sCFCy1fsU7uPzwthGjK1fxZyJ5VJr/
ouPOhkxGdqCejTgJUwbyeEzZhX2UIp07YPw4m/SrxRUBhp6HYeq9vtoXzrF9Ze6S
ZYAJeecSITqWBHo3N6xzHAPOali9/xMUkjVsBdkUnPJgO9OEeK3KzdraCv2HkK9f
7iLzaYU9nzUUFbdhlHq5bHrI5YvnzrahoMLTKDmAq+/P9WrLcGFRwBXYT7noaXBD
h7xAXk4u64JbQ++lg6IsP5u4k4UVcOsq8UWKHtpIn9Dpd7SAG5B6VX5SP5q8y/t1
L9jMvUvezeSTwMLvLQnvKwPFfHKJX0mDRTCJXv01iXSTw1k69MMXPWJDCr/Ie1Uy
6o5lGC2+TdC15oU8DXniIinb6SXklvAZOekzCuA5pFkR5+pCcv/mxqX1/Hy13/uB
AZqmv0VbRbgMB9UscvXGGAU4rB2St6jNc+zXKN82FXoCHSeS6ZEzh2tz5fdj4EIB
avJtSNpeS8OV67knnLYXu22ZPc2MlHrqxoihO9a0nqpdvJBScAX4zwYOS7yUvwPr
rmKDmYIf5KSVXAVzY61444LQ6teS5p3VQMCLH7Dqi2IrqfNGIzjDGsviJWPuBhMd
s1fSIh6Zd1RZAnqztwNTmNHSRlZvfiwcoiW8sqCAjbL5LHNC9gusepUtlkvi9KfM
2DvCdn8Y1iUTTfG/YOdBYSiacBwvuYrCb+NgjGKYZqSyg4y3r3nfULqRdDUAxHbT
BZPqd3ax39qLoNC5ekSKKnuW0m1XBAFrmRxLYU0o7SDC2tR5JD8C+3iDf9i3isMJ
5IVNkfASVMHC4Gq2ajYhExyKM057j4KPp0h6VylVygVFMwxMEmLblCw1/w4xGuyR
VLw6Dh1LOZZryOnWGzgg08twJNm994wy2OHYUjBx4LZikbbHOPllKyr936n4xsMm
G13IK9zJif/1mYlHQz95tkDFYP9c0QqpuUMWxshDp5AVzu0+g2lu81VAPDso6XlG
rg7yzTdhsRLXU/B1BSTxI8aO7fHR03Sv2DeeLJ/cXrTRGVek192oemyhsfnuH0Zp
zCh7Hk056/U3WxS1/M/Cwy+Z9dv1OPkT1SBRHpG6VQrDAOaoHuZp6S4BKB42obdr
YC9ahFSBeLnO5zaZtNsXEZeoP0WtS0kj1GjJwMQH9v++P7BRSv7opL1UZKuRG8LK
qPIH7BOL3UVRVtxayFGs9RNo5F+LvRdzTvWX5CcPJH1c+3p/FsfxmH/RqTWuWywZ
PUVni7XiwZacTl/Jq4yxfhsknYyuaz8xI9Bf3dMn+I2NzSCu7kP0c1s10/DuZggx
HaJ3BwheXJcuLO4XEvwoh8A4JQHayYB/we7Zh8hqjKna2GVt2OiqcAa6vcG3w/Ep
y8BfRzcETMvLWVpyy8CBUpru6964ynriaTamxSM/1fuwRzah7r6e3IQbPxexZ+vQ
QENh/yWF2kSm8GKJpiLQxdldu0YKHWMoAQa9l7a1wGz5k+5gLiMDr9qe6MX5QKTp
YnXofrzlzPeE9mnxJQccNNy2mkrRRJD+ZwSWDiOSCvKGaf4db7KL/cIjDeenrROG
q6GqKgCHdnHfkhme0+0IETgPCLT0wL+4gMn9JCi/jVTNMcQbnM+VPA0gsi+K/qBe
1jNw8kp9Q+tTekr1nJGRf7D8l+zoHqoOoS6CbDC4LPfVTY3/4pDEhl9GYYEkLmIh
3pQ/uj8EMXTeyAy3xgAB00jijA/BshiXgQtLLQbXuj7jyjUEcmZpqCHNfXsKPD5p
ZxIOr1HfhpY2bBePN5JXdYESem0FVyu6R+a27tBCCULukf1YdxAg9msz5sJD84Hx
wWjTwfYoOrzMm0edRgtWfQcSrPujIo+QKtcANxsiip1/JjwQDXPu7INDm80pbcEm
XaFtmpA+3rGW11JFjzZSnI5sfI2hZ8R+48pGLxo+FwHy7BrxmqpkRoNR2+RoLp1X
6fGi82Fd82ooWNFAt58r38aHGSQLW+0l3VGIK8zzgzH/Lo6Y0/J0EHqmSnjGWqyb
CQOi5xl/z4cZ4eG7SNyX4dP9Jn294ZVijbv11iXd2a9J6bTqihAnYdnPMOvWk6YH
m/CcW/7jOAYzsyJxSAhD9oZUmlxzDEKCeDiE6QaciW4/LVgyIAujbbla+kUYfRMM
G8VPk250sXSDjGxRX2/bjt1WC6mPJBwT2W8MaEHVkGGz4NI5u+8seXzqP5CyTe+D
F/WYQ2nZCxoYPXGVQnOXev5qa/Q/+DJ45HzFh1DxI5TNaWg8oIQvUoA2utb4KBrS
+FYdV5gdHBWOXaXASIi6P3wm1bukMk+27dQkT9QEFwWLbWhZKgJ4Pzl+MNNt6Oey
60f/cf2Q3I6md82ds3DqRM4JFpAuAe3x1s/9hNxeUF7t9LMfcGtP6PahSFXMZwhf
1aU1/bfkjBQsm1AzzVB8KD/pJjvqBTbAn/Kr2NLVGpgcdg8L5sURbMk2iBlBGkkM
doarDsMXcmdOthRenG3rUH3Qaf3XIug9ZwBsHElw9NGQmISfYyKjb1y0XalG/+iE
uEzceNVkPmaU/Apc9F7fZWph4QKQyYXWQ16KvIHGQqiT15DkytXojpNrhkHkaX5T
b7L3K1M6V/npmy3BvjRXl/Tgk/FGqdM86nh3ESR2Q/eYweV5PYI6yRyoHOMPPZ9B
DzUHxam+con6RU6vFlsUzxCRC4fyyvUSqbFZyG0qN5rrPj1P8k5ecSYY8q/M3iDu
Zk48rz/WA77o9MJXw5X811RR99hf/t1qedObbhu2vSdtWO/LuYk8krU8GgxP9YKd
C3Hq6ZdFb2oCM1aSlOBs4oMViFHfrULV4PLUOVf8tPZ5TCVlyIZV6/58dVoFXj6q
hz3Z8ldcmRfsSj2BoMwDte59Q7d/vN6gCRjgjmNciV+BCSjrK/a6VWfACDF7iW8V
INC2qdcJpe17XXah/0Mi+StIqy7FxuPHYjVW/0r8wYHXx8B/RWbzUA6tGm4x9bEc
3pF0sbCZ8/apZ80gBt6AlOQUuEPBRCOz8TfBpOScPa8CAGS5qQz0QnN4XCWKzbxV
ME0aNw0DtDg/KbUP1JhUnbLQcDnU+TDmlel52Y3zq6s1JIPKrm8OAEQCLpr5+RLK
dRzQlHTlL7WyOUvZSmMVkkx66zUECHDS1mh9/GrAoA1fXxBmZcuKi7n5/7QsIsVR
GKh2kqiruTd4IMBlWprQTwsIx7dA4VVHiep4tjS5fNagZ0gklePzU/pf0ocUKkES
T83/t0ENOATz3nGpvS8p1po/bAl3+mtgwd3xkmh7bSjjqGB3sKXP0g1Gq9je9Q1+
hC/bLeRcJ7m0oGQ6zP+JZbt5yY0W95q2Kz9YvFfDN7cMueP6QrBdVpzARetPs5AB
Vg2xJW1PAiOn4CsGMzZAAObedL1RArY4sNvZdhZy4nDxGuu9TEAVtf+pZBHwkAbP
5gys9Ho9axoLnyffx9T8kF1erDP3NwUJw+Y5kvZCEu8ve2AbeHLSVMpjLBjyf/QH
/7CWlDW57vEX6y0b9evRkBLU3JtmSijCKAe/ucf3EmakOAXV5ysmphYKk3RNQmBE
C3IltptpxB16/1GpJJpdbVqdbQSaubmknV+sET67vDJd2UvagazMXiMSFP2HyLpV
PXb50oHaYshRLoRf1/YZeJcUoSMD9/E8DTATpM7DCTTyc+o2KNmMSDYt3yZLr+/5
LPBs17+LkqG/XZ8hWiQgaxYR8sWIa71CDS3yfmnHKdLbwLLJndtDH1KCU70y/Kew
JbhPSKd6bUXUQzgNtS9E8GbVg/lzlcxgHLe5IS4ka65KoEHx9xuu/68Ur6De6hD5
a2Y0Gh2ERF8HRZxvMh5TKNJIBE+TLg5Hqp3KK23wqhNxnqq40l4I4k2RFQtvmYGx
t2v/p4TE4PkBedsvo9AC6uQmiZddlevE4XINMtQFdZXKZHWsNyyYRuY6ov4gem23
zbSLs7xFUD7UvR6v+zHAhZ/R0BxrAxIZnkm3OKS1qq1UdGGkhJ1eET+dK77FKSju
ovFiv9D4ci9p27LdmVDYYx2pzcAJitz1DeiWYaL7izdBOHqZVpQiB7yc3MlTzk4K
OHjlUcmBfM76TYR0d6Q+WgZGlECsdTSYd0VHiNOwl7ae5uHwCow/V4BVPWD8SF8F
joTzw3FuDaPAqlBM9dE4Cp//ifixs0l0CDIMcaOnUQLbRg5CBo83ay2SD9wYGHII
QdPNgyjz74W+DzaK4yQiLYQ8XhWgBpTlqYpV6rRs2pzbfaNbKFged2qpBu1mX/3R
55oIqowaGRuiSrtOnrDRzCAdOOCyIA7B7Gn408L3iaZN912uy+B+xlm3ldRob85X
IvXofGdRmQmeRgtKw2bmNboRYeITwKVVi4WVxvxoYr5Nr0riSK9DZqFb7JVCflBb
73/n6sgrNCs50uYp+YnyKwtT08S9lHQ7C/SZScMmfR7o0dTosWsQ0fcvGE607OMV
iu5Zgnc0/OK3oMvsDXKyEMv4Ex+DRkd4bzmgPlWS+4LGV64iSbd37FNcaNGluZtB
TMhyN9hTUAXwzYMJR0AgdX6RywO9OAz85rRqTUjy4WjRfa2uYrGO7K8Qy40FpyYg
6VLd3D71cRQHRnB4jjFj3Y6UD8/85SysbnaazySXlX7hC0Y+tAo28g9yp7ADc6iS
kHKw4bkbWRCVNIgzMzCSJefMYZWWAtHwvMqhshdEjUjuQq4m+sSZjKgbTL7vDafG
NNUpNC8IaHI77sLi0vNNzNcVuH/nM1OW1JxRI7V5jRXZ/yS2Px8F/r5Z1WGa5Yog
L8sMZ3JqXHuLGzvTdohQFPFs8SYG5bTQUOTlwg549aRu0cccxI1e9yhhlNkDQp6G
E4JZnxvhXtDDk09o7KKwwFg9PG+WQZIzt2ylwFU0oJMZiamiX+FX91b2dxXTRF9A
/sNJLjyp4unEcLAeyxiEa2NAfNfa8Thnf2TyvJeH2P4JIQHf3U6AlIBbkP7luJPv
9QZzM4WFd1OLSmQHCNUi7vuSHE2MywvulMXCzE0ynOi+6qOJuKmGnpBX24/29rdd
v44OeIXlcrqfg+pu+PKaHFCqkaB78IBhd88An4AbiFFD1NBHaGW02Iukn8XI/c6/
Iso827papM9DEtOcV0JRSjwusbbGa/0J5VrMtfAE20ztY00LUoVcAz/HcjtdfBr2
rlZQg+1PfwXeqOltcYa7+18vwpLoDoFJaZ5dCuoYTIcWKzjrTBYm9hNAtU5rrMzH
6r/iJUxP8ZBij8XU4JhOZevYHavkQG0fW+sI4YraVK8Ct42qU30THph1IFyAKZMY
EWrq90zc/nO0atrW4vElCRGI/oyTS8jrA1/sVkcWKG6aXKnjl4PBUui2adqQNz0r
bPLzVT9rCjOK8o5G5duFc+wf782lYC3E1SKfVoztVZuqdRXsEBETjgZfliqCcH5O
jxPpsMtyaIrWhDjBP5zzsi4QA3C1Gi/y5B5JsjyS6n1+oLkLUoV5wRNGcU9CAmxk
0i+V2BK+ZbEvW87mrDU0Q84e42S8s/KrDR/lSrhHtVrKebofZGBBmz8ZLOx0FKXn
OpnSumylTU0rIIfxG2KzSNJ1IimHEHeMTLD+VzkrUiGJ1qIH+8oiQOCX+6Si7ClI
iqWsNR9WJWMkqC4i8d0s+GOUHjit+17Zd3vN/VQOgJJAGyTG/kyc67tPTdF7BeTJ
XmkPyQzCoJnICw1PCRUQVHPZQd/bGODjhi90vinLmfHMqCGVQ3zIBI4xmhTg0dhr
UCJ5Yv/uupPjTc/ee3t9KJ9tMhrfSsI6r3IZVWJDuuKUDZ+UhUYkexsdRJpBeiSP
YgnN9O3XoAkbKt1vGGRLzwinz/rqndQOreRBhQQSAzXyMI0lXpI9EdoIghHlPMEv
1pAKcY6KKE/pcM7Pq8Kl2oTOIRIj6h1d5C2f9YbagRr1VqknCosnZFE+yegytZr1
6mpcWQlprwySrJxOdmL8+1UriwmZ5kN3o8JSwfoswToOABWfMFF7m6YkN6lXyHNH
mR8L/FCMdyHmWfWLMQAdaaWge/5VVYttq5qaDP/4xriHBTxohFVlNqaz/SHkvORZ
VjSi7zcs99a66pWS1rCuWUnAmZTUIr8ORZhh8AEZ94GZ0zDgvXqSjcfqCAa+4upV
3bHFiWDLlmV4YvGbna46ignYIA2/Phl7lKnenZbanMTpxyqoc5FFDhfdqHsKbUF5
7dRTyzE+8fhcWwQhCRjDK54k/8YeXmAjq5YiP2ub3fxE1YZxa2Za4vlLHgOnqOEs
KTQEs+wNFFlkxE+w79IYbb8Hrd3Cy+6ecrMEACPlTnbBi/dtpxkNeWMH6wM/sg0e
G3SUzMkOVqNKq23BV/1xOp+5TE7uMj0TjBuRKbD71FOK0rdsGdLgwQniVb06eUDX
sYhwNPp09ytfuE7tbkTY0/JzAp8N+kuTY5iOK/rO27g2bZASJgvNc2+Csl9wcA/F
D8rduW+9iYg/mbMlLo59sRcwUEotxFNoj0/sVTaYWMZ58/Pe9BOQFbO4BfLKXbFE
u1QqvCSScfD1n64acQntG4RUmK7Krb7g2YRPD+3Y6+Ji7nkXKgVxmN+ur6IYKhds
zdhomsqpSuAibjDbm8eNGoRVULGeYWjwc0fjqQAqa71NCSyBCL8ntXsVEd5Y67ke
QndmSWlxwzMv2iUboRU03p+OLbpG6Ke5b46bXkFIacEUqAyKkHizCbQ6bd4BWkkz
xNk+ab/xJCYPg7/MuwTq3MD1gdh0jTdyWP8bqN7OF9YHJacNSesbcaJSTW0iLfQ6
NyB5JJdDFxrzFvl9K7JNG9VumuPs14LCBIq36Yto1zfPAJvbuqnZLd59KUHIt2j0
kI3zyHDvQSiH/E6rICpnRQErhAACP2SAd1i9ORz7aQVieRIm8iZiaJAAZvBG4UC+
LBlYBLZTDhyz2dE56TgyOx1NkJpytOJRzeu507RwAd9Ii2dDNjy0nZRIcQlRcjX4
uVsdqe0w+cVjuZHsmf7vyHESLmVFTFrbVs6F0CZb9sl5WhXy1tuxQ3nnsxw5B5qN
xye5+6dRaab2acEMuffTlpQuebsJkKq99IvQ5gn3l5T8iYvgYrA9oeIiadyrZDf2
eh7+THHxl6jfmN+jeKz70jcLiyAUH6srXwmkIr/rnkNknUjyJnUUq0V+N4HlorqS
mSl7FI5uXpnX5oOrn/XG8wUV/IRv6r7j1VjPZ1DiAhh0jKFZ8ZCTEK6RXQKqmHP9
oqm7KxDfohG19+lmzFDLcx93uFrIBrGVAC9pcaGk0HIqrCnJmI3JBFf2Pc5E5I/G
EFRYQ+gaM0SPfnuczgPicRDsozNWgrvAJaemY6+BVih/U42GWmTzIM8Of7aBLin4
j8yc3s2m81AJ0w6H69V+ciTGmIJ843RUS8bRcKGlaJgbEuBM5Z0iVS6rF5RyMAOS
ifNtTXJq6aUa3NR9XnlDrapYLgNBHO/LUgEN1f58Sz65YiEwb6suui1KAF4RCO+p
ptNj/0uGIqzkRxbjwWm5ZwtFlDXjj8J3Q9DDQt60jFCwKNP3hJGFWAT07ECdoHLM
bD+pqnR1J7nEGwumeesI/he3FTy5/GQf5R/48m2JwxcXjVAdHnJDuX9QWnyaQ5y7
c2AHABZ3szAUEMjHmi5GeeKGepP6fwZyeQ6kzlCujqnb6p5fuDA+o79Ln/2aRpOg
9+T2qOtE2J+oW0GF4Iyk467yCy/vbv1JNltSOwvox3A/JAtU+KHUKBztRGydNu+p
wIVeJo180GhP4ElgaTZlJkKLcYPlH9tF8yfozYdw0wFp5SBSrlRi59zroAXPlBxb
rNnA4IDBSseP8qRMJcnPcfVVuDvUatm+O8/nNfXbvZFnstGmcVN550GCsQgahDOw
+hio4b+xPQRqnB1phxAswpHRCpr/5N5dNV6seH/cMtUBvjXkaA+dzzgN9ZaQIORf
+kQBVR5p6Ds670lqD4Wdz9SE5dP2UqBAuaTfR3HHnIfEgqjdqtiqjjS0EQ+blv4v
eGERcZPrtLxlxwTYLq1VyBMGqlOST5oPSATLGbDMJjjD3L7xTe7Gmb6uUKysRaPD
Lji0EHZuRG7O79xJpi8dh4yE0wXX4CLaI36u7wJWVu31LTwYXOdC87wezx0/3dvA
pnNIU8vc9+7LPeUICx/D3fkAek2GPXC/si6ozJDjXnVscAvxDLOeK+AmH2OpC2rp
OEbS2/l1XMZ6fciFjCHMn1OxUyjHYiOsTqIN2s0QeI19owpXydhN/ggypE9Wx3VQ
Y5i5y9gfR8YaU6ygRG5NRMZVbCQ79yYzzWMd5G+etcIEw2Yz8DTZ51ti2QmEXnhm
zDmb0Kn81C5DCDnwoHTmauS3FLrhthSLKQtZ2cCb4KIW+OWmirr91qhB2IcGJJLs
25fDrJEKCloRXgsc2zcM5uYhJ79vi4pgRUq2OLMAI8ZqFDMe472MHG9qVxD8VZSN
GkXJ/cnDUX9xNvhzQ43sh3RTI2dWDOty8h0qLJhCwJqR3RYYPXGkaOIzK6XiHCjN
+NBPDX+lNmE0MDdBQsRy/RAmdolH45+DykuvUZN839jY3ZKAu5o5035b+NXVCvtI
iooLaLjvT9CRqJDUfqBx7LmwAfFGXM0bQvb2n+4xsl5zeKJZWMeH6qIauqmafjOu
dirXj9Y2gorGsH2Ymq4q4BVwPAMTaf+MtUgrRL60AlAVZSkVGg171Ah7ql1H54DS
Io0R35sAv8mU15VpTGfp6byII6CPUCoTo7yNHvHaPOcM5VLXij7yJocS2WpgLMcy
0uREA3AvfwrJ6/WRmXA2dYIp2QJnXv3w/A380bY4ougo5hfg/Lcif2qFW/P6WB5g
XO6NOa4lrpKmD5HzLAPlXBszYWjzDA2/z25CU3qmLEfBro/QyBWK22FeHaUtfEmj
2xTPLiRKvU5u2uF3Gc6OKnPoALLba0O9P16QnhCOYUnsvEsJYA9GNHFGWbnpoD6G
924zyRHMbnv4Dr8d9HzIqT8Hlk39vIGpMqb8TV3OvUdQpkfdvBWmOgmLOYCVjTnV
uJ99OaxXE5VZey7nwKhm1wE/YlY2Cxa8HOIgAGioJqj5OoQ+M8Om+bvnN6IHwbC6
IgmVqJZ7Wbq8nVghmQAfgni1lqML5a+n0Ae1ZjCqvtfKmIrleDduxtHn/jO0lWVx
rn2FvsWf/dj2nuZEXSWd9rTFVbgiUXMAgvla9C2lxOxzlaJj8Vbc4KIkMOtNT+K/
IchZBQz6BdEmNGtwXHpemkSJmIUf4q0MZqq44FIOTZq6XSUKlrnnxcDQZ2WRFyah
3qsQMYfM+CBJnJwasCoWRSM7VmtzXai9lVkKKshi172zpG5XohcJQqSUjPRiqQnS
bt3gJYENvkJwJkD85kGWzDWqxVe/Qnkr1FHFEivfPe5q6ZzTsOdPpcmcHhA4UuAb
Qv+u/WaGqpEQLCgijMXrqooqqgaSHk7tu0Y2D0b75q+dwm2Wf5gKpe1JA0NLCGZh
YrailiV9LVm7q7lhhyB/iu2wChnlgNd1LiwUR4ZrXglgcRICkvo2ZzYGzNb3cMKR
mIBwTdA/96Agbv9MdFdIrIcTQToUxkET3oJG7to2xUy14ssWeNC/690/nZgbOz/q
fVnlsAm+4cdGpeN+FYAZs3I6WVgbfrZZE+Scn0Rn6/bL5mt5k33/6Gr2yXVs/cSM
P+cJiJ/qFoYTfqTvamX848ZMoqkAHc5kqdaKV1xrpeczvr4yM3P7jjjWg6QHvi+W
fD6f3oxmD9ApiN0jsnwW+LbET0O00aKU8051Lj6L6ckyE/WV7F+frJs1Q34/nfEq
ZltyGFBH7IlzATeWOL3L3d3xttBlRbGFbEGXjGXOJijGMfhyTfixDJfnAa13QqBN
CvlGr/d0lq+WyTUwiHFRcX1H/urr6CQ+SHLI1DDw2KHwupBI/SePuL9CQyroo2Rl
HESsJN4cbPD+bd6qgIKyWP0IZYIMy3e9jeNUCzKKNVc9b2kcWyRdd1qnXDzR0L/O
xelxCQQDsLxdZpnGNs9a12vBLvJyM97ETKkNrL+KcaeM/fK0ndbtvyuhJA0Fgqsc
t8sdhWmR5qJItgWN1/cwTBnX+9tZC7ITBXxirdvOH/jhSxh6SXVnEXRwavk2ikql
WaeQdqnmXAhh7DWYbzQC65RvOGauoWqbRfHNeGO2OomzrqmfjV8QDo8UwgPJJ2wg
/pfh+L/s/TZuEm5BvUisbLQWQQoaRRWYMKyLJ8vR5Xo2wWJvyR5Lk8LYiPdg2XJj
4R8qjHFrZwStWHBsu6aLQ/OOISH+Yf2Z53Ho1QTWCRG5J7o3lkNiGDQbhUh1ZIHx
fs9pBUA+hVWmttlMO8GKwS02alfSCjXW1RTJbXwG5Bjmx0PhsMEaUuRywqtastfX
OqNztVikG2P0r5aM9f1NwBsHKe3DcvSmiVIISzYMCHUkAK9Mk8pIU1rnRkhLnQvO
HHcpE9UzxLTzWzC2ACKc/sjJNswytG0E+3LtoJ9/mzFFsr5hAYyEshjMbZuR0mUd
3wA0fwPp/dzIwwsbEnhUZCIeuwbSHdriU7jl+F4bdSb/JLmWGUMDbXZM+sND6Euc
N42bh2T4/QQKTu+ZBIUoeruXKRdk1gnTaHwb8+yY5UZq9t6aG9N5CF5fp498w4h2
Vx9S32IihbEDK2PYnfOnlfitASdaAcWJtYdwHYbR5GfXO/GrilPSr/GvjEFcuWXS
yTngDv08816K/BzTo3/ZEf3j+3VlbmPhBBnKz06pML51hcDiYoOsJWsYCkiqGYeh
L17rIbkryd6bvwfJKR0E+1W6tbIjPeX69qug7KwNdM8em5afHuHQ2D0hWayaZYU8
VNZ00rLOQIqY5m9ayn+9IjEqAVT9aS9cnLnVvdnuOZ79yIMhothDWhoo1wHyZHJp
cUmBroy7eJIko+rZCwM1Y8jPWKfMGYkC5TVR9B2iKv11yGDoXJr8U8Hx04eYkzLY
ZAz12+3VeyX1y2/eVEtM/t4jwrus9aqz0YBn2OHrHlwpuFI6wTHv2GIilNwaZKN4
p2eAsx4hBvE4V2Vp3hPME/D6ngpqJy0y6OV8V1iXMUfpziqHB/nGJcYgr3AwgXrz
LbTZdLJEcuKXXquSJAk9O1Hi+6PT3rbdUTzFGqtib0JRUH+GsIusKnQe6MQFfOQO
CMN59SG7IB2lWIHkEic9Mqqw9IXPWZEN6tSdPsGJnkWsrfytRpGGtk7ZSc4iljYT
6ZZZebWje3VJYYtYQDdRknlCeXufKjkLQUXey/tiwDvNkZpNlOPIKtpHP21Kqqe0
uxH0JumROEt1ohtlgBsVqb10YexQywNHRJO7buXQYf8OBSGqu2zrAfMXeTGQBcnM
Td1OtPw7ghk+TvMzoZ/MTao6VH0tcCVtlh3taM4MfZBH5h8f0bgrk4cwyESRA8+e
XpY36yi9gVHVxfSkSRh5OJVQ2tYIQvaG8VA/2yiPJyLah1gF5UVVoWuBo7J/arlq
tBIybLV2t+E5boO0VJB+sADyzGSzLusDMdHJyszun05nWVwN+S7Q678eikiCtuSO
Gcdx33/KPhV891smLtcRYlKK8bH0Fw1f4yDdV8dK66Jkl8vuomdwvbOCMaG8HSf8
Zsiu8AxFUP5rlYEAYlGfZhHKEC7E7wm00BxYC2ReHlwm+fTzWwFNY8gf+bdf4gZ3
16Xp6jd8ohUOEweAbELfumP0yOuG8GH8pe6Rhzfcyh0NaUTmxd6VrP1FCwf4aZaX
1DdEcIOk18WQa4akBJzpSgTg21ZEkk1/srQn6UiySZoagRsL5GijZUckMuArkgKs
BhTpERjXAD4+tokL9cVMpeTqa+DlpYjmXN+eYCPoBA1hjf11SRuiOyrhhF7WOwPZ
VxHmfJA/HGQpHios7/MY60jdXEsRy4Os81uAc5DnyO9pYrrmugyjIcAx7hFMrm6g
HkZf2IXfDmMtctt2Gs++NY1khSIb5oDzZVHen3xgkWpM4WZTPDS9fdlvnKGO+BGk
pFucyy45a5Q8TbvMINQdhsln3AjIMHWni3zYfDq2KzDsciKIXgx8WEGlHFAR7c44
QBGuxkHcwghXuX6l9yoe/14uhjFIoRXMix33CsHQ0voalC34HdVv+NPwk2ykqExm
M1bCDmK5ooZvWsB3dyV7GRPi1sHQw/p57GD41swngrs1IznFfOzT0S80Dd/Imwda
PUA1/hE69KTpGj0g2/hLpP3AV8XkjL6/ymhsytPbHQUDPYYJ2M9Fvhxwy6B02wFu
aduzhDejLZb0P2hi5rHZS85CmKdy7Dyu8Q1GGos7zWtxtjYtVQDbQLSWwLsG73Oz
G7bv2wB8i6rZOduClE6UCRrNo5VuLrgJA71yJCipGP1u/3JR0ZkfX2P7aOILaN0F
VzAqwjIvpchWWuzNoRUpuvZ1f54XSC35jwyCOz0b/jzBVpbxKrWw8/RncYLhtXXY
AJsPo+6MOGj2fa2HBKlYgAv5gKUWSiCCXBz+SMBFIZz/us9yYlykAdhYK+EtgneS
zrb+H8rWANr36NU1KU/SxXNLbXfGyiRO8d8KimissQ9hboFSgIVENhZBSc3WPJF3
ytk8CqiD4UBUD7mOXU14mP+rk4/MxvI+P0bFEny0W/kqzMYVf97Ce7Kb5BfJFgE/
BeGmP0gd+Y5Rs4NkblnTbIZdRCkHtXgazs7HsGddwN5T/6gFjPpOyt5/wJxfuQTu
5LROIzR6kaeNZocChPvuGY/DXnICVjZ1KCbAHbVQAvmmyMysjVjPPFWUip6uO7n1
Y6xLDeqtCBT+hTaNSmwOUdGF7ANfNdrM4iDPl9F2xJA13uU3vNXgt0Q4AWsixUrH
lG5xsEWwYGj7NaeWswVSCuDS1AclHiP8JEWxgsqQY77TW9eAiGaAiPEkxvuqyWiM
yvNJnQ4mYGywuMiSR8RDbggC7EA+6WvAL3Y74JXQ2gjLFrMLSUHi5DgwBljHK34d
0pvpEXNH6S4EOCWlSnhQf4uTxY5wwjOXOqj6oJJ9Kp8TFAL7jPsHa9QYENB9O6ZS
kL1JrP49xk7nvbCws3jYiCwW4mcm9/uWjMj9d/gZJSFzhwr2HT6ADqHfXygRKdTA
t4nJiY0l4JI68BzcxvgljHeMGEjEy0sMLxhMvac13nrTFEQOiQtLhZn9ZQo8kwwB
Z5k0GU/kwTsPyROVtD+nUfdgTxE1VKkSV+zeBNUuFvqxLE3/oRktpJ4epmG0CqkE
ITE7IalB7f3j+2tO1l+dYhvtsn11DSTySYpG8QoEzD3stNkCQfjuahDNn6Ebg/mT
G/rMSNPJ0rf84XsgvBa5WxN6PjOGKalmWCAKZGc27mjgRVLPFM1a3RkCCTJl106y
QaS5vKmEdZ4r7l9EgwoRDDWif0WRs9eXBC9lXR+HyNcLD6n7ReBiv/sy6Q68uJi6
9jwfSWvzfMkBkNuLSpDQ1mK1L841g9FvnWJRsj1udixcCIT5OtdRnO8JbDFFBaKw
/U9aFJ23ukDTJ/7Gr8/5xJ6K5zs8gXnt9ZiZEIshFgskw6yBmUGwgxAKQCvC0rou
+7oh6JOFZeS4zK286cH67M2GM1KoECgJSEWV6rqyjqhbVp2VJtNoCELp3hLCCYrp
mES9uvKgZj/ZzWP0XrBLky8uA4dFBRu4xyIbykvbA6lmmOal/ogPVCnd5vLb5XFm
MakNj5rRNkvPiuoKrwLUs9mnhvZcgdM7gwwau+Zhi0MJNxvo6oLIGZXpVi0oRAtV
NNab2YWvJt8VM+Ol9u4FPi+l8yOGv1zGlO21q0YAGesd56GiDiVPJmsAODUKX+k6
bnaP/rm27plHX+R9DaCjgY7kjEQAjnTMXNxQTcsP5pBLqB7mSWkBIRZzt7VhJJRE
bG7j6+RkmSrA1dEizxcXyd9qFXaqdXVT/dsab4u8WcfFTuVMFYuf+Yh2BqHHHpTz
e8EB0b2z7QxVX6zdnepdVXk3yfoP/oGaEoCiOXZ4rjNoZjW8oyKjUOFyQBmDCqfX
8B3/WMJNoxwd21pdPQNptn84Fav7ZgBFcgF8kQYooZ27o8Hr5uCAKyqDOS9upO0j
0vqsbM69AtmPR2Rc/LfBHe4TodhyEu9rq+Is6HTppeePGjbcxzfQwAisP5+mRgMN
ckc1C1JDueDyFU9PlDjC5Asa24v+i6kLyWqKEo8Opcy5N072SGiSTXgng1IOHB1r
ebGPA+D7fPt915F10xT55Bxa7j2B/lVjvYjvGrRJBV1o37hmWUTCb8+BRI2v3IMn
igYWNOuyUx4aIf8+RmMGQSSQxb0KK+KeOkaDKlm7o2TsjMEM+j1RM+wP0YN5syl+
y3HLLuUuxTe/WxhwGguACMAlOwwz8S/D+dtnMqAtqL4p2SBKiQCXEbwFB9RcRGkm
SDyYByqbgXMxA6KRHWEgDKcFtsap6Z8y20/eCGMoPAGl5YY6tKbMDVGEQeT2sZWC
J0/2tiJRIJfhyg5TO6Gcf7FbgSbdUOKJffiyik6UY86ER1tbCH9KbZDWCRRc+8iT
Vmf/j1V+sALig//m3zGuBhB1d5Bx8EThD5g3MOQndoG4iWjh1caMxWAxXQZBZAFx
nbzHHe0W3GiqkzeeGTq84QtkZOpjufRH93MPkPoW0gnxFCAXC4/LoMPn/hBHxNsw
vYDVdvwxvFjVzSvJ7Qxq0oMxxWa+85p/JsXjE9ASSIYst6+quq9ED8X+emBBzW0O
0J5V/BvkY96/aVGFZB+3NoW40w4yBFRZ127xlHRtWXVlubzYi/PMM4h9bQ4d7+jC
Pb45geOGZ2h1mvH2KRkScFBEOiUocjDyDKYXNnB1IvdhA2stZS1PXowmXi5m4gRB
M6bCFpHQ4ggICd/RhZ5PpsKNV1fhf+gHbkaEe4WHhUYb9w/htgivGSfUjNTtAH/X
0CUsJSm5PotRV5QDWG0uqxumeym0tUGZhWVuwgf3oyQIZCELehVJvn2+h7ugRukr
rvU3IQDorx3Y3tArRGb4E0UyRtHmnVg93vfwrc3D8oRMW2XNlAFfR3mQrg1MhlRx
wkhP9DhSIvljBCa9LdoekWNM7+00gv2bRB+urnN1XT8x9tQlIIpI9Ur7DBoR+LuD
c2L/jd3eIX8iI0450mhNA/leA9zbm9Xoc8RABHHEM65zYEHZvAH3OFtDfeLZrvdH
+1zQWgNGf7estIXULToaaH5y2qt6W8+wEIeVT6c2MhuFy4OYQkbGnIZvoTKq7ZnH
oQGpG+Jatw+2TJRg9qbtwZIKqYHEoOut73JlzVfXuUiG4iQSqjMSr3V7fcPXydVg
TyaSpafNe/D9i8yYPCxMilpL+eEWSCZMzl6Itv8EoE12E2rUw6GVcbmBbyITvAMs
82A/liMlFsNqGo+WDnGBEqzV7hIJskruilYica/16/nO9kSRvyKPflSTXN5C2PI7
asPJZGUAHbiODkeqobmrQ0iikQYOFJ3Q+lCTZPIUZKbyYaE7sHeu3Tv9X32yeOad
/ztea0gkY6kSu40vrGAAPnwuDR0eX/S/RbvDxM2WGTpBzPnycgh2SN5dALcysE9K
f6bi3m/6NUc3UquiGsq5Z4dX7zXITY4rAPxKNhr81Kf3CI6oc81JaYVyHGZoy040
5T4kowGFkVBJVPt4R6ZzdCH+Hiocs37aIK9h1RgBerk5X/eziF7S8P5xXdqNFrh2
1j5IRT/cuuOKzc10S1fNDDMeDzuqGyIfbv5xFjXSMvDDNgSqS/5BX/41R0bDE5In
wAaG2hVilleY0bcVmiF2biQj8dm+Qnr1jl06tjg8qFxTCy1DXzXMkLnGzHx1cDfj
fqQHpOLxckvm60pE8Huv85oLBPPs+0DILwrHMwSZ/6PC3Fmmx2F4GDaWc5lPM36A
MhB0FrEh+1ynuCJu6XbCejnGEDMXx4fDMhdUEh5ISe1yK2OSW6jlMA5jEGPLt/ai
yJBmyO7EdQwZvBf1oeWZnhQrd7nlGpXkvHod37oByuRWD1l6GOSE8D+Pbxu4YDZP
NBCubg5u/D4ed7J2By5UtEwLbXRpC9EqQ1WWqN1rTHEbdI4kP1b0E0YCPwVP0bwV
0Hc1trNjbL040n1G4TzAJoKV+3YKoER1BYTUtG0AlJewEkyu25jKNBt+H9+KA/or
17atkijVDRF2MxG6W1kSiy8Q/d1AJLxsiXzWaN1cjIBpPkyYImxE+k+AzUdVcMtE
OFxaIEfUwy+Q0mBWq/ly0cJ2oN6tDIKr83PD3tHtvSq7z8VcM06jowq6y6tAW2/q
UQ9vy92WjAGp0AzGMbyLauf4vd6c4g7/nm87WOo9p+VCczCdWHAkbI8p7tvNlDOw
iDIY6MdXu9h+tMGcfNIohSvGvvYjY1fqeUDxRI5Tv/R5gP29higfLJpPBUcVdS4a
pt3QFhv8KJMBxgxIZdssCmac+1nuc5iVpOTVtuaM9P/9iUJNBXe8MUlY9itm3d7r
WzP06V8hrVzF6j63Z+cDG+Z6h52Dh6ZGZmD9+NgxWSoaqbS5q4xxk8TKcLndeYSq
xb4J+Eu+fQ3Gc4xdeUb6lG9U5tLOMKGKM0I4lFhuNqMTjrwUu/vCT1AhsW+6uBjr
Wlhl/zJFHjDsm3+RRLLYyZRgE5wwzIGUJuHwgAfCn/JlMgh/KviCzvw9O2j5hL89
s12FGtCxM/iWU3N6t2WXnCgbXS+7L0TsxIRcsekLyojOr6HH521z6HGMOGPyy2qD
G/rrtx2t3XOpQQYxiG2savLpa/ydUfhJsbWTaguOX/mDZzLawSMS3R9TFmCzQ8sl
a2vFSppkoecfCNVwppXajvyO1xrdVa+FLiqUc7IuO9uUGzOwBZbTtekSzUzQ5Lz1
HxJNw9TdaQM1ytuLJ1toH/YclCf7OttYcr46ZdimounzF0bw0azaDNkBJCm0jBXx
F4ifnLhFxjXUIVe5Ybj2npAytmLrckNh7nZqyDRH7y9F7DCKXbXJbvtQL/9hl7K5
ggknYNBc46j4A3l0+nFH6quR9QkEDl1ftFzXkbFuhOacRxLZOKqTm5uTaY2CcaW0
q9kxJCnn9Zr0Meny3CJer5xQ8ZrquXW0vmmVEvRa/X4HBfvbAOgvntT2iRgD+lG1
Vk5nP6np2Z63qhVKXQtqmGY427ZN9kJHOjQ+6xqbAJd3yr/vtnBQxTl3fWEoDreh
mMmdBNckyUQH87l81nDuEVQsZCVTHxDgAGY6VnrKwQsblWLVE0YZq6xGp7z7VvzE
ROa7xsc3IEaEfq0AE8Fja+CR6ckTh7uhxGscDkNTY2BHrpjUnEZPcSgwH+TtdTLx
ETLN0syameXh7rD6iIK6ggTdqMeG6vWfy+sne5x9pUPaZovNvh/jAPOy61Cgd1FH
lR7GpMdcz5A6F1IPI0+iNEVgaKE5v48NN5zWFQJFx/v8xi6uet+iLBsg3KTH3hod
f0c/Fc10p8bebK1Hx5fqxYQ2rIETSow57LVVXs7Fb6X522TIPzBVy9n1xmTkde1s
HFNEz3BX/7/CXXlJPdyBwHoYfXNctScASphN/O2upmsx2KJBvmDTOUNLAtTCHcuD
C6/pMcfGnWQDnvheEbGeBcv3NNlNlFQpYjNV61hVYnYfSKqvSk9cKJHv9H/myl/2
SswhNAa88ir1ikTSwkdVT9d154GzpJZGQuIAvsAz7wohFAgOet5Tl14RDPVAp+At
jVberFPDAEfEiaK5ibP8QQnt2+A98NIJN5sTyWrQ0SeSCIylsCfhwIUT2jdVIMJA
tURGQhSw6TiC90ljwV/I6aiN2Item4Dq9iiwfRwh6YzX3BMNsfKZH+HTW2sE4XrU
GAw829+7Dj+nlCoddM3fF+IISnRjGwfqXJSSJ9+A53LR8YN5pw/IO5yCKpxv0q5p
XWyiWq8uaxnAhDe1cYWIXlk5RF0Ixs9lZ8dyl35g0aAZ3wZLH62oyrI0Ch/gwP7H
jwD6FKUhI2AtwSGaFj0tjtWWZNreskpFsCUCZ+fMhiCAiFlCu0b2UQsAH5Lo8hcr
2G3XdT5PYChuuFEywnyDZMRIBfTk1TDslWue+7itmX9OcOIemUl8fAMEAUFpqBXo
UG6QlxmS/NNiIwKO+Pbx4N0IHinXnVHKQFUbasGZz2BiRjAOQVuczcrfr+kWlBEv
lyBvpwVv5q5niOJjl8tsDPMyWXU7qLhDICD8cgAPo27sEeYSlUhcFLYTWXUZlngH
W1jYn8/Uy1QsHZRZl4g/WczVAfAuf9dLjS23aOPlcH/UxIfA15hJfuDKn0UbwUi5
IdpFo48KI7IMiD+MhyLFh90u7iiRAxpOlGVh9pVbEsLHncqeJJE0P6U5go+stBxM
5MYj8ClonHPAyLY2/QKAXgSnpgZuKysWIuWJFgfmYjYuka89aFjV1M+y6rm7RYOB
Hf9zHoP+6Ncqe2Z2eAGvzgk4Ow955/une/AnnkOh+hguN+9x4LKOyD8fnxkuqf3x
M4Oa7ihNTuLe/eVjUgDAibvmVGeikz5lPGj5Xyp/p/DIxkWsz8ltkj9LNErYVOW0
L6HvE4uCQMvhTkaikJnU0pxzM6uo1upsakQ9aPimMkiBLoNNSDZHXxXtYVe836fj
4oMTRIHD1+21lQcep0Q9mlQKj+v+fSyKVhqmNUnlcKR0fDD7Ky6Ch1+lVYUADH+u
fmC7Uhwv1Mt/r+KJiqN+Y/4JUsHpzzblJ+LRvK96j5dyWeiLaiy4KLwysjtdegPu
UtkJPNMnTn+I47jjT77Xa/t4Wd2QWIC1Z/3stMd9L3RBmnFmXiB65fpBq86B6oH9
p8zOQJClKqPFPb2eUSxgDCOHnDGjfUhiW5dipoOF/9cYFd1LoO22yDZaIaCxqdM0
uFgIknjBE/acqSNKWYcD2RAQ5XJSu3EjqmkKFYIUGilthXFofCTLw/s1i0/4nsX8
AkblaxKJK5t52QhPfEdNScs1tK4xl4KIkDHgTusf+3MeBAauH3Bl4mqQxPlmwV1K
Jcdk73ryQdq7sae6SWdflRNM167Kg/aeevrqE+Mqwoer53otkko9XhqwsRCZmLPx
Vrbf/sugMH+yKrKaxGSzWOb7CA46B1A1fwDCAqiqzRKKDgZaI8eLVAhoJYpXXiK7
TBoSR8FG6Sf9rh4rkwD4IOildrWl1IMOajKJLoUbrbi2jivPIjMhgxcy3r68l3sm
i8MNu1fYSbZX8H2u0/nEt4oO8KQV80wxlf0V/AcmL34oM0m0W8xEqcLjLabmXT0t
csRsdrvoMePYGU1ha6F6aZ2eIfytAK8Z32Rlo5ViGPig+dRVJDPugUpAc3TPdYiP
dtYMmuuwPtIb79lBT1RAg5ZNzHSm3zJVcQzR/NtET1aW809lQwuhZEQYObOL6NzI
y/pEQ0uXIbOzwmvrI97Tfte7CUUiNVTb3ImNd09dZIDgOGSKL7INrNcK5k6Wh+yT
lp0ixs8p5TjhlSGFZ4/FjxujFMDq3ksVdADRQnn2K9romp/dkf3RyCKIO2wePdxc
yQBkbKqMFcq2Wr1I7GTiQscgS0k4tK3f1vZprZ3H3EpctSORLyuHYnqili686GDU
TUDX2Cql9fG61M1V1hMiSkVmzEVJnamCTOUIwjGlyWegcZBKX9tUtOQAiQM5KHdG
4HwjmCnZF2Ny3JUKmMIpH7myNi+vZs74Qf0OeW7Ugq/A3sTcEmApmztIAHQcWulj
QlkYO1ibh8xmqRFw8n7sUl0mnJ++qJXnqfTCbeRjRmE3VzDMn43RK/1GeJt4k1K/
926L9cCN1/oLL1NW4ASzBtoJ0KAwWnOVVF9VvzP7fM0Hbof9nrYM6rTugMeat75b
5RSM8zfVn5kVdDmW+w2pVodIi5PXAyoCaHDb/vKthJlR3ajV8RcCm7vvpLjcJv3Y
pZr+apMZlrvFzSQ8VkScZMUomE63xB3huo49r9nCfxwJgWW4BD8DqRnfF8iHKNaN
dJkzOssLKdh4lp6h2iRtjYh1M82ItdON7TNEyGMCp7LE36EY+k7+R27CeWOdadyl
oM3Y8G8fMPWUUwNyH/86AlbpmiBkvGCT0fF/ry7AtmczZhCscfRF1k2E3Ajrofxd
RMs59GmboLkStSGK79dZXKLfmz9l0xlcEgRNOWccykDX7HuXD8acJH+YG5pNGFSR
NmRuVFNiDm+CpMEpq7R29Ub91oHkU7hQxuO2RTk2HNHbUg4fCP52cf0Rytl2t2fe
53DgAEffBbj6PQEa5YxwU7gIJReJtQU0/W+onyyVhuGUPI1FlJF6VUfVladzZTjv
LYkpSguy+kYDmJGe/I/F4PWJgHrJawdr0oY2S3z0rIwlNprYp7WxXbocQR4jYLbC
rkgzVv90mYPxsRFav47rkrHHK8fP9FxBeZKk1UDUfxfJ12UeaTHckcUU9IPNUhKh
unXpGxCE/lE2dMbp88r/Fe6X2qJYpjG+4iPRW6qWPHCpc36YOxCvmc3b6LkO2ozS
HsHJT/rPB3ZgLa6DjYEmeRM04JUy7Th4aIQbeSaaNt4pKahFIxQgQoBKHYyB32sr
m8d/FhbJbY2Bdq1HEWz8PtfiYoHm2VoIoRwWqf04VhZ53SVDIf+GZ/CaDuEpCrV4
+ad/qm1C3HsueIw2YGGymJTHqvH3cnpgZVNU9ogFlxNGQw/LSUi++LquOFKX8Orp
guyYZUEjgdtnjEKpI8C2R31QRkS1nxdHf3HyZENwjWoL1o4r4N4s0uf8VbfRsv50
+8lSVDbxLVAaUBTKft2FawEOyIh0X+o3gzdIfZywtEUF0FxCz1rngHK1DbbZYXp6
khUHmtA57uvr3RkjW1k47I57etR2Z0+g4udz/xIQL+ZrFNQqhd9I3KX1+Froc0E6
MRO9PxjCZvvhgE1YXgd/6C5HEH2MLCltos9ksScSzjX+WCVvYbPHEQ36e3xBgNIM
Pc/9HPJPeI+SIf3jROV+yn5+j22CbaxS0AvPU/t0EHd5tpnckiU/fDaT8ScfJQK9
PWcEnOLQ698YwNdakkmuetaiKtiNrYaTQ/qTtGPkEFjtTHBm13SVkYXKTksz5a/Q
4NAZoP0XLm89qBzEORVP6YCaZFjcFY0i/UHPq2HE4mZohfnKQjJWsgjjvpaZiaj1
VSug0BtE/8oQ/eWe3IPFRIRcpHQA0/6J7SfUbqc3XYACFSJ8zs4MgcXNcQhTWcg5
my6l9LPx7xZDGcFlpX9amnadRJFYi/sgP9P/LGqsybQE6WpKC6XJmb22rg2olD4B
MZee/5WNMROXLh2EUa61QiI0DyxL2Gn6R7Mfyalxm1SLJkxWuCLZBpY4PcYSokR/
j1VWD9Nit6amR7jev/p0Fqore6xl1G3OLsAHPExpwssxyccy99pW311x8L5oEvDC
XfPyca9TVOW8axk9UChtVMfQTosLzRanVoW9Maj1kKTe3wK1UK3+EgBjsT134Z1Q
EN4S+s115mk5KOZW+lADGI1jL5YYzliRp/4xy0gOXNm1wJkcJsErFjrnO/ZSwydy
o3uuecxiIv8QVldOdIZ36RY5PJSkYUNu4IC1x31i2e1Fm6Rv6I+nyhL3+EV7yhwr
p9MS2hbZlZExqbPt8zFFsMIWM9tSDO1g5JeVCbj0H14SQUPobJzPXrBL6XsbzMkt
rchnzvhggktlCK1F9rGSAUUFrjeM4g6sORPb35v8ImbQlJSqO+UKdU33cTka4ZhZ
sESjGNz6EW2LUxZRE7rtKqKdXnJBCxPM2La/CiMjae2MoG0l9/3Z1nnDAM8ho/YD
E2aR/NaRavKlpauSm2QtrGG5wZ/MR7LXxzGiTC5C/6Q0k1fAVXskSP5PyT1vG8l5
5j3GH5Nx4UqnbelpH1T9a7fEzI+xPVQGgmTiVZFQR6t/7XB3zO2Qy+OI0oCD6NK1
2/KbsAqR6ywwY/fnKZz+2TJ4H9QkeMhdRB7WUgU1LAF7I1jMVN+Ftfn2Q1ew8buu
iPRDibuxmGwCo5XpHZAw+DdHiZiQpPmJQ7XWGhuwmPkh191LqzULrksw+O8G9Blk
W66VwsAnGNdewtWvovE3/HMV10UtdE/rf9RIuQXzS4MNaUHAoHaDUwQdJw8iDURV
0ZPFfkjf1P1FFqq8deLtoo4xTtaEScQvrm86n9DbKY8JUVRsLF/g4IQ8BbM63Ls2
SXZIQLe8VX+OK3hzCf6LUCmfCvNH0ni14TKfm2Ex6h/uFA3eV81LpZ+5EIZu36ND
Xz7bCD7x+UbDh9lAWMMWdgGci9ut18/OrqYbZzpTl4vb8sLko+OXNfddn7cY3Bwv
N5wtGLt9btoJmY8cNbX+9eKJ8L9uTT3iHxezK2A/foOYi0qgwnpiJJr3GWmsGrUm
UwEUaf6nQL25zdqUq9HYtCM58Sxdvv5N6Vo0xfk4ZaVwiSbcsNCS7zlG6zuEfoJr
V2aoCmksUW/HR3973cGAvokt3A2egRo6e3+uD3yx4r6v5P37SbbxW1oz8bPHw186
nePpgl+7n+CVE9VNa6T9auZCRmyx7YxuYaKS3fTb2CPiPINbiL7TqjrwccU6EpgX
POcazVP8fsjG7GzvL9rcPgrvvqcsgq4zrJ9M0yWm9HvxKYE7CjTRSow3pbMDfR3Q
cZWF2kP0QQRhbpr/HtCqsPVR4B4qc1CNdSCG0Ry24TWdv689OrjcwXkCRgdLxS6t
GBil7XwdBVyNBa1ZVcjgcLk9Oj8GHBKtwfZ/0Fuc+uEvPJXpFf7YpSTWeTg2ncEy
8Q4/6RObVe87BlYorNGRhbaH1DULkV8VoPttd/KRgeLndZZVovi+gcV1YihyEG8N
lDnEoAhDohyeaPVytWtetbmuXe7t6RBxsmdzvVuyw6RrotHneG4Ny/IBOXbRKy/v
3mI+EWqsVsRJ8+nIXhohY5+sUEM4asoV8vFUDucVEmgy5vo+NZmPtbYYX69L5ngq
S2GiSRiPn6MHjJhmNqhrJvxUxp1yrRxVNftJylQ4iayDTX4JG9zwUEpAYa6AXEwQ
Jn5wfi8pgYZhKiU3C1a+lLIsj5EpcVFvHzHNTYPRprHwFeAnT8Z4KycebSp+yxEo
LEWJW9d+gvtB4H7ljvv7sWFhYOgeifwddnkmOgydCBHaSI/9J3jHquWkbRqN+KUF
rr+2nR/Ti3PJBD1tlhmnJ2Xq7ivqO1X0Zb3OvMEnr68mvj7YdRROhSmBLy+Qn66/
f/RMHu7cf/yIIJgQ0IDg4WCKcdLbJsAO7BMfzQsm5zUijfwkuvnywu/AUHub70yC
TQs102QaXNSvKon11NKXwFaB0Z+oU0EDmomltAU9X8RntrDaCAGRgz59rYFmiSYA
0l9Hh8rNoNZGjyB7g546aCta9WIFRhWi3l3Z7sFs/ImDXJYFvibCukgvUUEN1lTa
lqeKu+8ovM5Ap6daQKR3KvcoT5Zv9OkC/lTWV+jJcSyWeKOkMlKYzQj0tNITD4w3
RjLD9XrMAU6UPTnGNAsn0Haa/LltHorT62AjS3Ceak2QTjLCndM1QWLhEINTRHUm
/3tmUITNPy+/fWQeVH5W+0OOp4sBaUDiZtkC/Lw4x3PrIMbqNdwRI+wu5c/+SvCd
PL5PaA52Za7Z8KUdHI0q3yqjduSEtuwQRVjHaMGMIwKGvf5KMsdiha1bY/rRrIwX
Q8Bte9g3maDM31JGaZfF+dneIw+edJ2nSwVFFyMEMa/eN8/NZRTKAZtH39+N66PU
XBywXb/8Och2WpC8szxDouEoidFw3099p7RVYRxyQSTkZRSNDMaR1qwKWYqL67am
VWT3XJoVO8JPneKkoNIOoHZiVPgFhyeqRvfGL0bSbTbGgavY3T24+1hunkdt2agF
8QYvsvsbgWthFD+Kpx7xhuTYXE4Fle502oSTXVrbmHOOWtN0XP2RypfLr3w5sN8z
/NHCUfnkUMH3P86kQBw39O6O7k2vKaQZdHg6S56qVWMn+IF3u09WF/7NH/OmPjfw
8ISNytsWzXhxbsk4uVTKZXdptnpA1FH+tQw4tSD4qdoQckR4aEYUccGRE27jBTrx
TDxyne2Ezu2wk8/8BYd7jJXjBdsa/IVpc01onxFnRcEMU4Eug+a7cbX9ziis3flz
2yIzjF7pwSj8HnBk8BbocyoPWASwPuADvTsynakILan+MGdldUHXYfKcYCQv2b0i
ZcSN5szKXWNnl6YbfLBSWgEbaCJCQVMXcViNcRzaJEq3sMcsIcEsKWxtFs8G0MqL
ytfjcglV7gEvdQZtNzHwHVdC3bd2FaLCFlMQwfQMTMvdRCnWuSe69TLBKMoZrT+0
aW+op3EISqBCREWmvA1WLMxo96iyU+5sdIlMD92HRLPxJhOlYWWwAeE1pzDj8z20
6iihaAcRTCaL9zYGxy+EGaA1vcLzgTqmzwdpsm7RsaWdra7I1zOaWDFbBQVsFxki
v/SnEqXca+b453c9y/IsGA0Jp2ReBm+JBn0yvM5qJ0eJR4pTb93j8yevBXyjSuZB
aiRRfID0/jWC4cE03WHTEkLO5+mnINwD0F/AO4jwVuLyd8rFGy/AjpWyzqLlYS57
oKMD1vbKvAwtg+Qr9RHC9iskgHlgifmd0DnsS0EPWRFZ0TdX/WjGlKUoXa6esUew
sdbGtswPytf8Sqc0eO5eF6xtCQLpCMDaePPFfRHy+DrF/8AtnlKo2Ib7JJ9qbt8u
PhjRfw9nZiQrfxDTa8UZpdJdsm6fLmkYrrlgfkgVnVCPxGMmVZEDTisN2T+K4RI3
jqcz34nTcu/zCV4AxBAe/KfFZiFKTjBMynOTguEya2+XJ85idsR7f6/nuSDJ4+KD
W8AbckLJmdDTjMpsX7Ay1QOQ5I4vP5rDAemc/EIiUC09BN5DytJMpM7eui9LDt9n
wosE9vUpovG2lTkNyGKErq2zjPiKyjlvYobYc2BCiQOQcZShB3GOiIc7okEZCRRC
EnQf2j7crHclkwo3yOy+Ylqc3KLce7rVDB+6gzjexMuLW0ZqtrbgGF4cfNaTDgUC
Me9nfEy3Pz2+b8pjVcaQINGo91LLzVzeq0+a7s6lXh8VyqAfyY7CcP82NNoZ4GbE
sMtAbSw/FLZSq+2vDuZakCrH76irMuDQ4H1L8p9Rk1Q4TN89ibIK8FtUh3YKHXJo
13Nw5pD7zA8dlNuamED0I8GKlax6yOtuJ2DxqDr8Ifg4vnpUuPgl3TuxPvRes69U
uEPxc6AEm5Ot9/0VIqJfiqXlHLJQmeA+6eStwi2eMOla6jNoEiaCqdxJ4CMeXuMh
vPg42jSJSuZQVNnXQOqyNEBJtgApOuJxJR1iAtcvaoi8ehk9N0/MchYdi8C8eIAi
dEK3BvdiCMHjwj/aQim4GHfFOxicwEdWMbO0ldS7jEbbmAA4rNEWG7Xqb6PBfJJI
7v/7BAxG1SQlBd0RJHfhC7pCqUa8oOokeze3gLzN1M2oPLR3SN4Tc1cRa+bG2iNj
HhpcjYcv5d6tMsSBx3RaDW6X/cSwbCTSGu3uXceJD/l0ZN8H/BAtf6ig6bS2hmTs
DW84HOV/Xjdq9qlDMykrfZADQDXbwNanNbUOyuHAK3exg11vn2SZosXQA5iCMWc+
ZqJJosNSv09wnX16pd2wYOCWQe0jUoQWNsIfvynT5or9szRMkOV9hgjPzAUcFCUx
JjB5MoldD0+9hR+Mj9Q/N89nchBpMG1k2VTXUfkWfVqjXAcPfpG1LGZ4lE8vvQ8g
Vl3Yut7G3K3IDdj8z7EtHaHKpG/iC38ubZn4XVlaOmZHdMYVYMz5ANiE32804AQz
TIsHi8/HpV3bo7Q5pIPyZOpjrtIoxItsM2S1tqpq2Ef+9VZxUhhacJo5GXW/9YsD
y1AxRdv2eKzV8b61YmRcCm35zyF2zhDYoH3KiVPadFbCq3Uwnmd2lMYZm8Fbm6A9
6D60lVjy0JAPZvEGKI+ojnAkDxG2Bw2crm3q1BqQ2TI4DXG0xp4mrsZU4Wh8wyih
VyikX4N0OXfvcdQ2XJqxu0JqMMJdH18b0FGmWfVjlZD4ldRU2KLtedVzMbNIGxy9
3lGN5onsWoPI5YhK4i+JCUBmte5xRTU+jzODA75HTfkmzUpTr8OiYovrUIV2VgKs
9C+LC+7Dt0cjKNlAZDIrvvLYn6DOtbu2p0usgmGavnIecYh88BvGqam6IE31wqUf
lTZPKoktykbVnWqUV7AWt0Aw6TTU2Lim7h+j17OoBPHYkoK1iH39ESPDSHtDzDDL
s5vgviFtfMoveEwleFWQzMJBNK8lW3W7i34gX1VqoHSZWYPwNi9rNo/7e2IXS8zp
H07ynRkWYFWzxJ44hyA2suV51Ys4Qhmg1CMBtDkrea2InRHGZF/cdykMunrjaVpH
wmv56b2nK3/gO3heGD7YS7ZFgaS4twpd0kVqmVhriMgUQuefu5Hbtd7P1bbx/tVM
yLNocmTOCLrLjPcAZYqYz4CFqw+asOZYJKy75dX1AXDoDHwl5UOCN3e9odDINVtW
Z3+wr2xtezb8DVzTvxtZijxvWbVWa7qXHqd9d/wNU6o0jaZtV6TjVW45LTcQclCN
0dQjScPy0+OgL5eY8XlX4xwU/74U6y996bF34ueCT6g3kLimkPGt9bvJqToyNJiH
R8qx5XNMXhdyKM9jfggumQH4RZTSsNS5BUokfIZBCDtVLh6aFRFfzWSUFLlAKNDa
T/FynE7DiMsMMiFl9ViazBEMLsASIdzA69dRCnPsPThTvuiFUGa4INBRG8miYqBg
2nTZJWe88NF5a2s/otEB1/0b55ab7Ni3knlYf8rT2tNViWM2SFd4xAl3B+tH7lhf
VBYStQ/bOB1w2Y4RRkqhVUwhF16dUgrEMWqoTrqghTLe6Md2/1ZG4TjOdJAZrcom
zLz6Gf5TUNd29a8xr+hClXsYlmlTKS5UYdYVVbaytl+COc8IWys9HoCOHNx4JI4P
0Ytr5xkBGvVC2EKU2a7DF69ZCzYKz6TBI0G6hr8A9aMNNokLPYGFhWypg0qp3p+0
FkCNxzhclYR/D40PCzuwBhN9GnbBWGZbkiML49scTJsYDEkMbEeoMAGSsSmS/TT2
YG8fLH7IeM7BO6fb04rXxq82Nd5uckvZU6ovNJflqIo+DxMnR7sVfBRDzUA7Jh4F
5z3GMrosjoZLnWDjTGv4GZxjNQVI5G4ASHTFW1L3igSOI32upCY/7d/qX2lHvEmp
tPF2hilSzHXRWcAe1lOxoXZNwlsn8kXWVDts+UJoD0CpQD1cF5sLOGPfBO0xJYzk
jGgQSWFoRImeYpPTvgzLIPBi01vYNZoQB5QypuG+c3sUhj2VlhUOymIYkX3QHOnS
VETOTvkjl/9/7MfiQ8hSLQiucwnNyJ70mZ9MBsq9G+gCrOj+SdYFFhRGNQx0tyKl
dMc+OqetPox9EeIxk9NzX0OGG9wWGGv513is4kLKH89ZoNoKngWw3GgujB9ZQE8L
x59O7IlyNVBDITVE2KJNSpdoyTzRMsz+7eKgCkxr59FnfCRMm6cCixvMI/hgU8Zj
cpzILVeUdISuuNMhoFZMoTfvZOkiMUhXG3YpCooc9cbvlo+84aSfy2A1vDsIl2Yd
mckh3EfqWgvdMY7CLLabICU3L3XDcJXQRE6UTSV6wPS0UybYl1/5s4lGj8p/s0ax
iW3HSWluMRMbZUKOP7DsiZptrVcla4lPzP/YYnLqr7f724gOJ0vjYV3DHSGgcnLw
B9XOu1dniNkugopIQHogOxkihsuFbru0ySmz+9usOE2AeZKwPf1w8esm+RLepfNH
Q3OWRBGdohrc8FoCiJsY3SWqS1mBk1Qq/NhPjE1WSCQz+/TZ6dvhqOQFMVm8hhhz
okT76bUCsaliDnlA9Brod6s5K1k41Px++5HDYysHrotXxzLsnAky5xo14j+I/xRi
Q7HWqqnSyo/izzMjmqCt32mG+Acd3aQSZniLuiH1kv2/H2ZphL/I/9QNeA62SUor
APggWYR+vVvrRwl5n2hIH24zbtDo64RGdB//D7QefZ+SaDW3l4PS5XqORRp9FZeU
H4IgBPiF5lemdbo/2NOvzbk6hPc06yD8oQlChcd93WbpLeeMo6rnE+PVy4FyOPFQ
vMXAJpOUYcvwHnQLI7Gi87MUhiY3CGOjDYvkKhw7KsG4tfflrHRg7gzn2AISaRkQ
QK1a8JtdPAi4qMrCpAT8wbcBwGZAB+WIl/RMFG2fIHvji1clHJHv1k1e7fiMhBjG
qNUzJK4KQTwCtq3Aj0VpcGvN7cGI1kJrCZRb5Q+qXeVA8LAHqbRRAEL5lh4iyDTR
AvKP+3Gh2LssPvTiasoahGUT7Cbormpehb+GA9BjqYO7dzpnIQXx8btMv5DrQ9vz
BVtTGzXf0NNaOxe9C/Ubuzedkm9HkH6Yz+4GJ+CAk6SYtAM0OjV+I2ABcsXRr8K+
2d8DOzg+XrHHfzW/1xoJUSgNpIgUwABcHa732ryDh+QbgFVBJq7MXrbq8zbigsdX
bQhbB64J6ULExSiViwy92lOa2CUCvlyI6EiF82XPXIATo5/YksjGxavTFT0+sxmf
EQUVywJCx3bfhoTfTjbJq560nIoVSjiWQy0k+Gp4zdHtRQIh7oXlh7E5+uK16pkP
z2J9eTb0f+9h66ukDOFLzmDBqbNRC79kqZSorkNqUgcLRIM1xsO8zeC6pEOlG5Wa
mBxn9mr1Df1ZURYQGkRPKSnTT6Uwma+xzleLmiiIB59DUk2raaA+SS0yk4d6Ps9g
JcgoDyfduAhLNgwfzFSQDoXfN7oWRMgIBVeTo2KVjrsHd97NR4qU08wkJe5lPsPy
LxJ9xLO3aB7Zpts9Wbmz2NLPCSZ/Gq7Y/EBZyQ3hAznyYsRIFNyTXj7bv924mJ3d
+4Vjz5CrNLiDtl1Sl46xCaMXDTIWEieyTiVFQYfuaXtOJa/ZuHVWYVapDNccH8Bf
a48IJuRCSHJk9/uyTlTfqMRhf1RhLEbkG3qdrGD0FQA+ZMEhfzfAMLsEm+WHLWus
3azlRoPsN/G76JUKwE4pUWzEbeodJiUMrY1+Tl25mjGXBRcf26p9j6Gm4V1A1eVU
McAaywa2tkBXSjNKA+p9dL/tJ+GZaoB4FOxnPOP1AJ5gXMqHYf9zPaHuIH8lpeEq
SgJHvOV0lfn77IECDItlekxw8AI7JBElRn2CxT9OwbZ4ZJ0YYSU7bjdsO3PruZz2
6Vh5pVo0Vc7gEQFKPIw5/NzU6dEnJ8wPviKb00s70A0y9ePJgKxvjgG2k15QMLiR
7s2pihxs/fnbT0jtPJPlowZzTEICX8qI2uOE3853cD+hDF1QgJG9mSxtFr+erl6o
IoWzcte0QzgdiUWUdo19n1WTobM4uHq1YwjrF6R+lJs0xNeGRnZTby5MayEQs4Oc
Qq5sirc/SgsyaLLVz2Zap9IiyOsUnGHqUV65T2HBB9fNW6wCqiRtpnKy0kpn8Rj+
LtxOVsYS0NyNAwM+HZ7VgUTcPCpkz9xPa8E8SBY7XPGJprzcLwhAVzhKoIVeyVwo
02i711El8Kst4mNWo8I80ijWwLlgaoMw/mzMO0eEenGx9V1GJudkxaY3fv14tFFU
UzE+IeNdsZwexwbAJBFmBejxicDRvi3xEwC1nMf1GXOpw3v72+73JGyhHdS3ugBH
gbtF1ycTSmkE3a8Dy8IWOwkwvaQF+iASW+YUP+ObYNXNg7HAl/JAor519yg+tJAL
ms2l3dmeCrjGD+9FXHi5Pz/ZGj+8iAs+ksSPhWxTGS5D95e/4eAOekY0q0AVszRu
gL3CKVFHZLtLBX1hgQxTvXxj0aH12O5DJvToTvFc+e1NDEml4IAl31jx/A50j910
e/QkPqQhQK0sQEYNVUJvyM5hHuTYB2f7ks9DFCHdYdBbn79X2BywHDYfmCwVkSuN
6MDEVn+drqNgrOlDIxjcElZXuWIf8t+lgQ+W+FAMeOvNtKQHR83tCbrV0J3kCBQM
3GoulAVJJsUOoFaL1SdPKhsSrqyDUjDCcNnmCDD0QkimYxtuCnZVZBDWGUYInQG8
lzP0AZpYRqNSbEaGIyPjTUapxc+oObq4X2ZTvoxmvaylA5KHzF5QwrWnT1ELkJXQ
YzkElo4V953/DeHbVPagczl39hw+n3i7+z9dR2R91ZzG7P3aIOmV8F/+TK8qtPPO
6O72LbqzEHgWT4C5EYIygmIruWWid7H+XolNoXt+Pgv29buijcUKv4flTdllZC6D
4qvKxartpZ+cET91DZjMhfcSOqz5a0GZhdTTOEH9mMcaFehrFl848yc7S8CtH4pG
9PApsXhVaUoVNfDIbKHclJKHqV+XXSPHeUIBRuwDbBQ3YN06++7yhHtN+xAtVYPc
qGxomjrBkg5s1+JplNztfnBUhKFw5CdhBVVE/sjsciNp9pwJey8vUD1pcRPeSi18
NgM54UJIBXX2cCSb3uCHBQfhxSBYPnm/eNfFjyVJAe99wwiExYGk/RVGCzuIByVI
GgjXcEyiDytsIfc5s7Twqj58poRc3R6gTCghv4IF5VDSshU1H3QVbtSTMPbAHPE4
foT+jsSpwm/pPJV4X6d8tJn7j8wOk1QSAFfgIDJZfg7yytZMuzS6c0ErmZcgdQmt
EsVpR4bHEnfa29WzNDUkSUWKundYc9ULLqv9QTxhZwA/irCFtJkX7U+iT2PHt2w1
4R8EY6O361Nm0jK/iImjwjjl/rc8XreFBOu1XAKcmxkCR0SEHF8zHl6im/1T/0iP
AKrgSe61BisyCbJV6Mq5iG1pBIdv88E25vKif1lQXlkIYbSP/mWwVoB7lEQ4ptmI
i9pn6jirRaIJUnS5HuuomNfZ8G2Zp1i2mJa2v1gwFajPydLIPRgwC2T/RYv9vYcx
51EGnnLivk8xIUp4dsWRqpQn59IeWbmZh/b6dfg7N8U938btkjAV0ixmD1AeXYve
+e/yxBntX6CBLvPptvXnDA68/oy9PugUmDUqMxGsuWmCRUsL15IldMst1wGpzls7
f5tZ0jCaUnQGjkmGkPBE1NhfNVpNlJpDeYb1wUyZjuSEbdkHELjg9RKCSOlBQYy3
tigqJs5ZV46XK39HIEnb++PxZ6Cr2dVhPp4br7BuaGxQBUvGsq8NjINH/7eyCfXc
uUKR7shJIA1WdCj9nuz6+I0BX7pwjtkU7WE3jRmcvCZoNEvTdmHhZqGbyUEq6wN1
Nqkw3rWCBKS3LW0O96tj72YLT9F6VrusESDrQ6u14WdofEMEc53xA7NdHwDCM6pQ
Jv77iGEkSq8YAeerMrFdh0pWaFNJsuHm2aYYPjWr42L/1OY0fW6BLKfVLEgiIdx3
ar3PJY2WIVBVYVrq69kUzBv8GnqGtWmR7K0j4XPdtpYFOQHNMiUyLNwUB2qN/uQC
gVsl7V5C18yLGNmg5+v7RmdVQMnGOEPfT0ZhFmDA3yRvsgjhSSFwBVzwXEpe+U9A
HepT2RBX2dQUbK0LzS9+U+ljx58wMuQb76UITPbCFRaOvqRlfr8itMVyzkKTC2gW
UnqRJtwknRv2xCAQAfArE49wHBcyy/BGWTDBKb1f7+VWNLJIMKScjmvD0cKkyceg
vqOiwMGCFkn+OnBLZgSzjdfdD07LMJEpDcI9UlVAaCg5iqUnpWq6g0znW0d6VjXZ
+Nnx125XnxOdG0yPxbR59fN0QLvvPcXpIVy8bVPXe1lUw9jjEv3OTBe2QowxssBD
amMSqeeZTBc9n8bRsLaYDVKntnv2i1beEVHmrD9vbDPPYdQvVUHQySodJzLk50EC
p6i1aYwz9cMiHqtepvtLvgxOwBd6jIspt42ZppMWr58Di2Yz5UxN0tTaO6EavsRw
2KPjn1Ti6jGH15oOmu4UcRq+bCkkveslG4qS1Zy5oRK1Y7lzI8YBvZiN5nc1tiRi
W18T+o9Vat4iZfYKZ24xJlASeVpIwE+ZRHsMQT0xsYhdS1BS8W/bX1N7ugF9FHet
tvBhbEZz4E6NzQt3LizArR2zW9Gu7MFcauvzeU0vN74IFQexSIYNhjP+ag8j0kBx
2OldtkbPPEUNSpsHPfnwwqr8At1N4wASnfhRcgrJpIeNoz7wEtPATSL7sbwI4Cgx
8UDO4nn/BevT60O4MWPkyU9hMP3A8x7/OS+72KS2EMYR5ujMctDdD1wZWDmz3BQK
iGPouu2E14eEKNzXVmkkE8r0uO7kNbfa8t767F0GopRiz81zoqjeNH+xm85HIAMC
n/ldndfZowK51vWDYydhh9Zdjc1L+NLMmELH1bzeARwDha/50GqyU7yqSwTrR4Dp
R9w/zLQ8ldc7XzxB6Mn/cscihxleQBaNJveMhe41+OilG1R0GHyxevv9HaXpLoHT
5X+V5zPBy6Allcq3+lJ50Tc8MRKapoyFUO5TybJR2x5pXY5y+sOOvPkCHrMdWlat
0J3bOHBbcdQi2rgNXtKQyfYRkrYHGR88eU2WVEn3vvdmvCshTJ9UquEaPmwV5YDT
H9oYy5efllopqNKxm09qcaVWieteymcC70jKZjTDuK503ItHYZR8OpzLCBkgd+J+
X0QNRLgfCuGwdPEAGTZgGanZL5IERNWgB03fNMyypSwsVPDbceFm2AGMFDooZ+M+
A499NnD8Q4RzEirN3u2QzgGq5c7BsgoFqG70AZZNrhcXe1DcWZl2uvZybX+KZr6I
AQXoxu+bmnkMtTES+xfQJo7OQlwGp/QCWkqHwzk+9WgoEZO7A0rd4HpwWprfAKu6
kFFEfwmuZgga0TZZqNGRWeGOsTsN/l+2m8RVhgucr8b/qKEkeuglc8sLHxuhM+C8
0kVO9gBYPexzGLusEmVG9SQ99SaU5hBnr8i7MGSEiUzsnd4te+KXKII0vXrSvUOo
6QzaiQLF8VJJlucT7LPDyjPyHJTIBfrDTN5q3FH7fkALu36mwsSwH1K3tQVS+FXq
YF4q4rbF72IaumxhZ9eF3frSQ0nVtr4gsoP/fVK9sGGZGPVeuletPzy3dJZMAlTG
lHuh7mLmk281gYwykMKjrtLjOixqBJO+ilDM34dpSFeIgjlFcOgS5SrtFocdoVYK
Ms29O6TUIPu/kFBbgS13HUy6rs+BVMTzqtHN5nOnJRGKYvrVmuJtc0vQxIvzRkWz
G8ROICQGf3ZbX0whAdRbVLZ4sF18mEl9nMJhaU9k+2incqEMm+ksvanl0arGdRZG
7MDQU3NAkuCFr0P3Y47wI5dIr44G3yEVWqaNfZbMQGxS8pR+V4DiD6WywCNxQvek
s8kf6NwVqJCUxC31k1jdimVPUHE8F3JsJwBsYr3MZnjx4B+eve/TOu9qHmtTlmDs
pIrf25MTRqjTQH5o5p9u23mQtr8yqZ5TbLhqCAVNmneb1uG2P6bETfBOQLzSBDMU
1roKeVvFGorQBAmCjJDaYtldXzPG97l0pVgEa+fm9Dp6vbu4XVxOvYBHkdhTfEA4
9+XyEKzxzrcHz2qRL3SFFYeUTuOJzjMpHaVVUTN+FjfvTDYROBdtHHv2LGw9Gvw3
H/3e0/Rub4XtNpD20aQoeUvShjAuFHIqIicZtoBSqS3uhLog54dATxehSBah7YwU
X1Zs3vDEuPTB4PMvu0a89PGhHTcmxUKCWYPch8/AkBhF7U0SgqhDa4MFT60Wcfca
mKdMhcIKPMDlnGR+LTyEdPU7KF8yEIeDWUUZRuJigDNFCcd5DpT+rQT8ziySCQuk
ga/SwQi2f5KqY/t933OGaZuO9htxLb1dRIW/kBolxz6YpoRWEOqb1ZiGdj1Mu23/
m9hkGqK7GPqXlel7BQSfX6JthNxC3ROPtCSsR2/ilLNTvven0JRxP9aksjlpJUvD
1/qK7FLb9UAXOE9SEeIDovGq0qSuSc1FjIH5h2wZhMwAX+jLUlrP6FvOZTc4TzJH
Pl/MgliCd1TjXUKG5kLk+RrXWI49e7pTi2Fg/hp5Zi9sIwo9QavR4MaXwAd3yl1o
JfCfeWENlHz8Pa1FQfeUWM6L5lls229EImd7BOaIymJKGPNaZ8mSzz0IMpavbsJ5
W+nmOLTd7ouYvIBCoOBVh6NfFjwFZE4QWfpHhBQa+7O/1JOCt4rD0VVi51oLSGwX
0L2ozq4zSB8GeB5o1DFvxc7fzUeSEyTJPos33gRIUTJkiATdYTfZRiJDbS88EVrF
nJJP3W2QChJzZxgiUM7A4YybJr256YDW6F0Y1VqWpnlKhOjRjEHozpsaqRjWKlsP
1IuP478BxFWiAve7sBi8YwO+kFtCnfO8sQ+Y2YaMo3/0KJffhbfNUN466afMgGaJ
bW+xf2dLml3gb+SE1+QINSyWH79bdCIUb0V7H5msjMFuS0yn5ekwEBszUUmJihYE
YaOy8bc7YzQgT6Gh4FKqat9FJc2Yr7QbdouM8X6h6sdWNAhDQzYTfbAnUH6gCGcq
5yZGu1VbNrovMbh3NvFILOV3p1HSyKcIlixJlHSvFn4ZKD5cEsQYv0zhCA9fboml
X6DriJZv27QbTFc+Mbp+z1sPgDFJ2P0w3PdqKBppwBDgEX6JO8oYYeksEPcci/9+
kZN+fTrpU49+FDaR3Phl5SNa/FDmzKtDsqJft4h85l7CDPilaJssjp908a/HXms+
e5teiNb+JMjHBYdRzkklRF61VWrk6vCIDif9K+K4dk9tiurs/t4Lp7kFapcCw4O3
DyeBwGj53x/LGJ6tP/k1a0oaw8YkJ+jp+ooNqB/pminTWiAskLVRpa5Q8/fENdIK
C/BrPPY18gUmyolCrFnygA5pQ5XKXyUxKCD6RsEuwuzCQ3JqIjBoQ0x3lNwnw6XN
FMJmdSxnKE8L8QORAW9G2WzvS5yPF8y8Gww0eFXQWWNaRhybkMFTp+MlYbJVDSVE
ChhP9/KHxZWbq3hVFD5s9Du0jr11dAig9YfKVu0DHq7FHOY00R1szDU0/rRie4oG
2aeKl75+cbHobnUdOojxUllJ92CDRdo2LsX66XD06SpG+dW5VkFjNdd8P9D65JYT
u0KbRUSApw8NFpZ3djZ5bahbEUlaSH/p+vUzWGx3RSbVWI3rM2MBN8pnUXcv22NH
FhSkkyl7Dqoy7w6oSSsD5BM56YuLyF9CzcUkOYx2gyWEo2iWtbuoyBZ0eOfzmW6p
rrpD5+Cd48MwvAQF9/JTMYxwOQRoO6T4XfQPlJNPJruPheK8EOALeP1cXZTLdikv
9wERbp2/W+VIIvcau/JaTj0kvPC6hpfnZp4Zf1ocsTBp9zP0B8FoEF09+u2UTByZ
fBB6rEfuKPpDT5BtxSk51f35Vwz/EL/+ZXhlqEzfQhWvFuQFbibF/LYN/eSgXwZh
wop2oCKx+RJ1cZtTKmm9fesWji/AvqP1qUP0X4FrLU4iuOue8JGCidZU7wMP0HnE
iur2ZShBihHYPiIyvtNk6fXYSIom4cK9SwT8pb7ACpxZzigyialYY5joAOtHVYzi
XuWOeIIHk7jv4PINmu4nwNg1HMrUJIY/DA+UFXLcILpPTBy5aXPtGw/Z3HBbY15T
V7Bj7WRgVZYRSFkClm/4iSRYvHjKHLTdVm0gYFb8c6uBiP66MNZuaFkrC5VfR77T
WyZn/WBF6wUvFYI4+ZuKe5T/TiI3v1XjYcRd52Ops4nPYyXEW/FJL9laakgowEB+
5zZdXpdGyE2D8yjm9+w4XG6Zs5Nk90hhRQkIntdD/vMWJWLUtI4K9t6z/pIT7GnN
N2BJDaMYOGXQk00Ny1HFG1ec2fpanwNDzaVbwTMMvUGhBJS8N+RRkTXJvmD1LS4f
dvfjYw3FUzMbLERkCNqQ+u1uvi/Q7foqF9ptalC0vHpjQiQtnvaISCuql49F1vX0
UnZ3hfsY2R3DlnkZ0U2E3YUxOgNGM2XvJW+UVNB56ORNomJ8yUzl30OKJW0NJGVC
hN6qbPxKZ2Jxn6rXzemWin5Yx2ui5QxAqAGUiNg5KJNB/gEJm7jhusZnHqr0jRls
+njrAzTImQtKQ9dsDWHBSlBZaPtWZHNNwmA8tyE82yaJycyBTVHTC3YAfCumn6Yz
j4Dq8hx48PjwCACiHYrMZ4GpeBZvaf//l913NjnDnVe0hAnDhtPnF96r2DpImZL5
fOdb/8/zrrWoJfJQVdgv/e7yQF76Mn7EG4zb/hiuJXZPWNKIUBuSLSKg7A7FiT7H
f/ncJnGVnqPb640KfTASmjMHkCyCr3IioWS7vGJixmkfoaatPLc/+edgQbVWKUAj
YbeEU+s6/bDDQHHdeyWfVO5ZlgQoLnHx+VX8e3fg4DIBgkBn5uVi1NL+aPsGewfj
2f+kg6kB5MmAO8++5Yb9x+2vHMQx5f/bbiDKw/25TkcO+caxspNIN/I/dYXQdSE3
qGao+jJyVCIaxrqqx4iKcgjVDp1sh9YVvnjfFgLnNmng/CyblAPbDmLJ5MVbCPP4
lKJtnF4qTr0hx5KMb2gziwVdgFZOxO1u7UKz29iBHQKCCbUM4auCMPi86GRshAj6
RcZnRoeM/TxY4ElL1YS5ih6rSPPUXUYu70Bkrp3axGK0RKyykV8JEced3zebT+Xw
x/ylSL6p2nSY0GmccgYZjPn9dyGy4w0wF4YBIP8WVMONE5OJX7Z+0BW4Kou/O+4F
CxL/aUiXy570PtAtPW3CYxnsb024yhyF2pHbCdjyqwm25zLFdHHmZaM8ImK2Idxb
wuzMny9xLvqHKj/E+MsvbJjBp66+tnuoDNSqov7Bty6bdpVQwP6eAE3/iXy/7HCN
NJiNRro1QVikQwan6emYqY3iQrmqQltI0FxS1PG0ztiqWkZoofNbh+ciY0krsZNz
Mez3Fr2pwWi3JEcgrrnwMYWQzgfe2Fp2JpVmw1SWbpOKdc2mYtZY887T20T4OI1Y
W/dCW/mMbvYeYBEL3JT0ahBnJ3tJSj3KWzrPWcZwKjZV462gKIPPG6weUG4M7M0k
SIUh3pOB1AcKaaCFMeg6fS+o+Yr+wYAIQmJvSljMi9BSksMg4eNz2jVQs6M1PfZ1
y5F1FCsqgqseL8fZaicJNmN15pw0tLGiGjvQAT/fpxnsEPlB9uk0ZdOrfwYL0s4u
7qCLMYaS47Iau9Z6VaDvMC+/ifRs7BFV/mLocU7t9kgPf/UQzqXnobvWfsITIdKA
M1ImLap4xPJyRiTa7OTbHdjLcOammNLwqCUUQSYsIS9wly0erloKapA47LdPmoxQ
E3wI47ZPK4/oDvVvx7/k266xoaB60ptUbLUfqA4WFRn7m6qT/Xq7KzdHhDrW0Wam
OTNuZBjblyxNy7hKMiscKHur6ly8t77+9JF7zbj2blpOwKxJ4E/5gYp+oz9/xZPf
Lc3v392seWQPMg7xh70K4vEJ1wtPzSMw3Ym7cj0XNGofQwTDmPoKEh3RTmHX0VAH
z1q3SvGWRoigQkDS5Mu0Ku/dOpdXg6baHKIv6KyCN6bZgICo1Cdaz59Bi1J/kU7F
qiF7VLYCspG3GdWszfe9m0VZC1NmBmnj7cj2vy7o/9kqTeCcr9yeeMT9uzuATMnB
U9bfwyjgObVLElo7l3WszgLcJEWGtMBRUW/ecZOYd98GBnegJeIVsgB3gu3tziSA
53jVPuJjAXixgXuVaG3qetx0Tb1BWo2z3DQI5bhZi1cHpmRzLDy6/5IL0vIoQx09
9o6F6ALoqbRtAGNLr2/QRk+8qmmlIsA3biUeX8cy1OfZ6nKWpEg8zDIrcjk777sZ
KeGyL/+AIqEjMDkGP5WjMnRTmnx7W6ls72UZcPozZAoMRSNqKf4xueZ5nMR+wEhB
5Ctqd12HEM/KtnqQxByl0LHd80EMCUP/a5q33OED7i5PD8zXq1I1NDRd1a3SqkUA
h5WDVNNa5gmYYkRQ2FqCuP4Gie1ywj6wgpFTRvl57QX1ysr8mZCfFSVLbQLj2kNN
yMKihqTQWV6EU53fL8++4uogs/Tu8/QjVu5vcDFsnik7covA2PagUvbCf/TeLpM9
JfaiGHNaEcWTSGFJJRQv18F4lhv3mTEWtERSW1dCXXzmq6Om3zA09nGn1TnnW9T4
dGDw4EH8quc+w9Fw8WOZbF4vBFxfmqqK7KiYYHQ+qgpJ5vAyH/rliu5X2UrnFIX6
X4IPIsHEtocFL5aSqUWZq9pd4KCqoaiwMScoOIhnQQTbACs/I2112955d6dh2+2a
Vi3ZYrHJYPjwBpXjydbL7r4s3VP/C2mSpSiZYSAfDBEsfOk1mUAubneqdqLj7B9u
rV83oq1xauYKJ7VuFOoLOGP3y8A/l5jBqDSLrrlRBrqlW4hgf09WiryeRC9pk1oh
WXBSBhh8uYsbVLqHe9VDXRJFotSBxtqIR37s5pKVapXvL3cdCcEztQYvjuJ80Axa
A+Zbmkun9t4TA294ravi6Pi3H49JEJjK4031uwdmXXguhNNilhwKRemj3WbLqLXt
XKObBdphmNtpnrOATtqHaiw8RBuE7h6e1FbDYAzeD+LsDy1AsVC+7AfGq/tgvWte
geLjiy/Vo+mdHH++V2kFqnEF15TA+2lc6S6gXn/3iS0+NiqnpaQjbmfBOn/rLnoC
uVC2ogv8CJTj9RzJK1P8GikawNeFSAJ1ENIgO5xW2HENprbQjshFZhV3rEmsv7lR
By+Q+/SU4jINinp3nSwbY9xze97WeRTJPMdm5geWWAOEGGqpYsSTu/TuTJTE0TCQ
dkM7kr3uySVU8e6ptHjeXdS4Vvz7GbX7dW5ouFKzGlVNIWONbueL6319hw6+TB4K
eqBT6sa0UUYpZQLLcXQ02VA2BNzPMvoGgCYk85imbG2gb/E6Fi49dHCxIa7FPub6
7usonGRqymxde+4PhJNo46Slm+2rkycetoPfLsMpmLXVHTOabfTaQjBrP8C5Do6e
462pM1D7K3WU0jcQrUnfAhImg5N5RHowhfsMkgyvV6or5AQLk0Ua7aAj0g56p5gs
Dvk8x3wJ9rlwskhus0HDpD3XMIa/7UuQdaZRMUxZOGpm4E+p8vYOcQZlO09ZKAhs
iTjvJxvQe1TlwpwbA4LoGiVCN9VD8ryypVKOfXmm83oIOzbDPb3M/gstb4YYVxIZ
YhI9rsrtKthJaF6POM21mzXOVT4o/mcfsBL8MdIEaFmmdMnknWoDOyjURWGDiIg3
zj3LPPCx3QxfcNBoopoUOGKZ/rVIjLfa8E4r8ih1msn1gvTkNVfSaMV1Yj+P9Vhv
D9wDQNZHRpHvzql07oWTmUlcaFxDDc4fQhusyB/BiQnW2kxvJFdRJ5WwbMVhSpa1
VwQNQPXofxxfIaekfiaulTFUWQNrL1DyQu5+iulCbv3H+CkoK6J1/0wB80a/KJqt
o0Xnq0DFHjlVMy2FcWibK65xUofS9nyDsCwKlT/WRTNYtueCd3+hY8IDcUH6QrwZ
tAfQQmdizxshlot2w/qaI/kGD1SQvrDl2rlmn2TvoLFxmcIhPxsglPLp40l4o0gC
LMeFx+lt43F3CjfyuxfdD9Oy/CtZAqYkqcUbGK/44JcBJUraX0kHZiEu1MTurLlt
xfPTY0QuU9eCkloPW1mRXAtrzhjqZtSLtgVrETPZiSdBrOQQWcyGDQPQhEVLZBe1
soOn+BbCnD/N7dToAayIb+dI7dlzeVdj++VD38d1Z3Xp7wKh8aqaDm+CdvC6+I4N
BrNkOA4jjnhpp+2qt6i8oFi29LX7nIg1Tqpx+71bl2VRK5hMtfii0gdF0MjKpvta
Mh9g5FKXzVWCduXUklNydLNoax5QhoErDHsdHd5rHOvhwRiClPhv8SrcXR9fnVxB
4nytSKCK45CrVaCjgHfsZEJ3tvScILQIBU+jBlpS/udCBInC1lIKVLZPC0WjCxjH
/4PBzOSs+Y2LQiiJD8mXGg8U+t3RVW40N9SCw5UYMBQL0w/s4dxLSIjxAQx22r20
5bVYaNsc5VpjfC/U7zPJo9wl19koZ/+8jgbk8jKo2wCzHxM9e8gwBmY+560YLAxF
9jQmg52nw/HcYjwNLIYvizOJoEKNkvOsD1JWX6LvdslPLJOlkdtqcjRU/wagMdWk
sPNEjh679kcPu4hbxv5z2kn8+qaPAzjGlUCAZB0IlBd2v6jmjgksgMmG+vckpVP7
tYzOuErd7/bQKCCFAWIUK0TJzU7MissaL5NVFsCoVGCeUSy+DTXYTO78j3GYB5m6
oviDHqW4Q611dz2anpjS+OKSfuo2SIBEtU0YRanVpKljppRAR5XKRgU2tMOzIFwx
nQN6zN6BkBGxB5PBQSIpID0ndwrKhpqCDynG4bUILO3z/pvnJ+EGYZ8Ptv5AzvGC
+xaR+hHD0CyQWWsbakfomloX7IOB9v7BmFln+SNIk6B5Y4sdBE+0zRKNXY+6HpW2
petSgU0U2u8MYhje0TXnbFlF2nxNPP+cKvcJum1TSN/3vnDnYdFYQIHAIoCXBfJ9
1WxTfAFy3bI7nUDpaORnUFU1I/qwcPgqpAn94kcb0oLj+OCVncGMwXKVm9CiADYg
VQF3bM+QR4dlLJ3dTZHP1Zdcb5IiMK5KFAA8bOd3Rs9du+j7IjV1zzCoGJi390Tk
NLjQraAHZtpy5u0P8s7kvTLva34qjGMrUMXyDXzWJG0VAOg1nD2HE2yYb+DHnVmL
mp8BRE/KOeguf+pbYVSYHZJb2R67ZiW9krmVL4SHCkPJWRgmiHIT9zmBfiAlt322
3rdsed3XkEsrD+GbPpa7Rjvz0k8ZXPoUPvJ0LkwZWoCQcldyOaokN7QovUV2uAHn
8QUMx2Vxi4/syXHlGm01YhwUiJOObf1gJZTpnjrFRX5blnTLcB6twcH2y4OXemLS
6eiCqy7PAGkJvl++pjJtDBiSE3LX0g1lqCawax5LLN/0N/PxATMrnPIB/tcVRDsd
k7s+w4pZWeTkD/o9ZVXG1PX3jy4obRMzsINqJqs8/vZFfezrp2ItWsdzoRhQ9tmx
Q5bH0vEFCZS96/iZB2T4XyAlc0l13eL9rlZXDpc4YzMRykyFXlLlLsaGr0iiP4a9
g/vZwDuL8YBH4KHDQyHjjTly2ocb2Pa5Dul5irqNR5+Yc8+F+Nbq/wR2NUrRLAYr
irFhwalM2RFxN6LdDxU27mzZ1KT3Hr632sfZW3/ij/m71ulBFoDvXqR1nUWKl7dU
jy1WRm/Yah7hNVTYY47tvCfFdHuehNKMSkIiT8oIdKCd7eDFWlAftm+SHydNDz3W
xjxiykcGLOWQ/ElTTmg5K/ofzGT+CQ1PRM8JR9AWIUIVCadT6FO+uHo0GqKntb8R
FTMx3vmqTOO+eKPbINagCRXIvug3XCesRdr++GtzC5g0Kj+gM8x+OhGLh5TFR4Mc
yPWcwEvR8028pD2QOW7DwInHzANQcluRUylfEuozPNRvgc8SRTglX1ZjEk45MIEa
DhCEDisRAfpDe55YefKeTQpb4nftKkiTMFkNrJYfX47nJTxCYngrY6/mQfnB+yQN
Pf4eWgfo6h5hsoeRfqtj4SskmJJT+7YpFPMq6VEcjdUzThdY9IeSJedqibBLk4FO
u3J35V0sISsdd7pGeTP8ffQhBWpow6+nwgSDRCaRvrRJlJr/1xbnIAEKq9qCFOJh
HzBucRJVM0qhDLWPEaPoai7NjNQetCD/jMtVZsUl2Gc6LT6zttdiU2XpT9yK3CdD
LSp8ZSwpnHnqU6nbXoR27/5NqUiod5Uq0NpK5P+d51OWoLoWcIslnAmmXfONvTI5
gOypa1p2MzeNr4+jAsuS8FeMbLWrY2FsTaNC0JYaCSfys2+Kh3sL7msL5wgL2NPM
A6UsosZRkH8Y/9uqC0ESfdJCYTC3rb396+KFPFO538PNJO5slmipvSlCoq/in2mw
h5ZX/fi+WNcdpuvVDHmFmFIHaCYwwlly8nsuw+/DhL/t+rhGISoybqP5j7AXtXv2
TdJf11v3ZITcDdbEHQQR4unO5GrL2KEEVxPLRWefkUFzawDXf7cx/Lpf4ruuSaB+
dwolr1/JUQ/sGtI+2bYmZisZ0qyS7GQYhNRh70P5qGn+m62w2GOYoNH2dGNS97IB
YvPF1LYMZTLsw8dqyyBUK+euMbEPVU+3R74UN4zyzGH1B2beCxzd0gbnY1Q2lQXv
xRpdSZlWsk8k9KMalwl8g7e7eE5gRjgbzQc3XLL5NcFSaqoYku8xkhNudMUVjNdp
eb9Xum7+p3A/PHOr7dpdwyXQ2qL4VEGeyizdZm7B62IMyDcTOd2Oxa/A52aIInVq
PuytqACwQIsoQDViuSYI5MNkP0ZnmRx/wECFAkZMY/3pV4+57VRiwJ0uffbp8b+6
N7h95t0c0nlsnwF39L8BxmEEdB9lZlkZr3/tiXyDiIqODTtWT4vbzdchj3vCIWI/
qVVobnhWi4cfqjsDO4Q2PqZ3fAmGtA0L2a/IrZjnD89awX8lX8U9KcQqL8KW3/gq
3UH56T0CxV0eH5BkwRzar5m6gbCCr3cfYducqyR2BqOEUQlV7tYr6t27/0hrcEPr
mxjSpm+Rz7o1h1c+o7rYLwA0uOjKtPnnubipMAVE9yBVrNwnDqLRu3IJSAuUtME2
kQ0mBnK4m1h1oGUd7j9x94K/fGYEdE32uJj8XMnRzGTboGvle5ghrDtkIm5JfkwI
Eq96ppGhilj0wecOkWZhpMdTJwy04q30D0bi8yG4221WXaC7Vq3+du2vExpDm7TI
+BzkhpWGf0tjPnXk5Hy62CTQzKapmhV6LtJKruUnRCLXCZslCwQMz5K4ENwLplMl
5bkTTiux2TNW0knSqkrqPVtYfhllXDM+WNJuV/mjWTjVP5oT8FAHOBMdkRJEF+cp
Rt+tftS/D+U+VOTeMeg0Iz1jjpFDzjJpkZKH8jgx8kvJdeT9fZaizbahgKjirRc/
kyQ5BHmXFeZXLfnHv+tNlgfrT6CbBju8wndlU6C/n2dkj+R3+o0NkLitzORPifks
lqjfJiqgcrQXit5S+ogCD1JvIEKSBmD/zvm1CXz/NQk7jTl7//GYoTfob87I5HRI
xJ4fcYfeRpAwBnFT1C3sdDZ0smlxkoRdtEGAjmKKCL/IMlpw18yWwCo84siGHW3T
uT5UiUNKVxzRaNJGcNTBXjpNj092X21K9RmGxqmUMpjVjvsRBvlrUWXF8XnIhYkr
SMXrftIS6mlzgcRrNhmPCrEbFK5rGtTX0VUsLoisbdCV3wubqNNue1Lb592nP7DF
KzRFjkYlea7hPEnUN5ZkdzGclwhg6gzZtFP2fOXiDE0888P3gUpcV75ZKyBeN/qa
edNjqDy6IEsVSVDA1v8O576BKdSEOFmCATrEZfcLQF3PxKd5OjeZ4mZtrouSZ4CF
t6wHsOZyZZaD1gtiADQ0GXiukd7RwMf0XgPWRuakmQDEHBrDe3bgEc61fUWsgGpp
5XZNjDAGfDqtqmDpdXjmGkd5HWI/HkBpBR6mSoavh07ELo4kriAuN/zXYzBISCKr
TR+76rss64AGX8UE0y6BJK8WpAxwrg2TAb7kbpOmAQZn2Xie3ZBnXxN2TgF4YGo7
6wNGCQUsFXJyeb6kXmUu4XPa6W/VnPbhiW7ATZnTfpw2HmE3Ab64y1dXU/WG9qUG
WNZ81ycif1/lzWSVLiwqoJTV5d6ElXz86jKbfgeRWrPevqC4g1alLWWC2mAUdIxR
25HoYHUPir3GlsQjc3IaRsmjVI6mCEq/YFg4cSFVTQag6vrWSqjcXgyg3x0cs10g
l+vKFfeVFhwa6+IVlw+DM28EEHwYJNKgFymg5CNzZvuHbn3E0mNGMoEeoUK5GsDJ
XoLrJ5Z721R8y8QHeMdnlWsxZ+WGs9nw/MYIlwOFoK95ChK3YpKej1jQf72awpsa
obF//WYJS17gzWQKURVrURJv23TBJJ2JBq79xzpWiAcxbt/GzPbE8sQYTkDmpRMk
abgS73FWKbBQReUXkKL/eteQspJdWdN9boDHRKOe9Z38CZfdasIQc1VyWOL1OCZO
7wBd6AWGMovqAM+a40dI+YRX/igS5elvOZFJC6ct4zb0qX6HsHFmrQ+8lpHoSZRV
v6YxWlxIDaagmpU+M/xPeZvcKkAnChWyUG6Yd8jqQZIwOEfHOZerW22P4Tq2Q2xR
I4+qkLkxOTW8/zM7ECP5qUZF22GaSrCJ7Ip0VJuo1bnKQCpPZXDjZPCQ1TW+Tn3g
45uEMhqI19xWtS1Npl230SxE4Vx7aXeAUWfCNPqXcGyVDWSqv0m3aXOd8Q3Qk4w2
5xfW1V83+uRT+1urNGgnY1GDEOsAi8nKvC54tQlkTidmHNhAHNiQkx803iuwgSCt
knKBQAeJa3guYLb+Afh75i2G306D5zKc2bKNNE135aTYk3o6I0tvBUmnpQwpKHT/
E61xSYyQt0XLQB/TN6oUh+vUsz5HjgbYlQDMSQTvouqzPbHX03TNhiv7W3YbFsSs
5EDdOlcFNXRh9142UqmoqvgnHszrLf2vV5w1UvxI15Itsc7if7usa55W/fsyy2sR
CjFUmyWYTsqJ7a8JhBnylma44jUWSvkol0IRRwR5LhbNJN0vxtWnfIlMH+vjElEo
elyaFIXpqz0JThpUsKIJs/Z/Q1PhmZeWQQua6F8QO80+8nvNgwGvC5rImuEaEhIj
M0VqNMrr1ubMg3obXUNkUBcHzOQTMpg2/XyN6wKARQIpr+9Q3gyRCM08uTGv6eO6
j0apAH7dpi+zYksQyHVJSS9DOcCqXeFVfwpGrlxYeD+QgLcndwfPcyKUCZkUgWgd
eHy6vv6bSbCH69LwS+hz3/MSroK5u23gYLQM+8Rq3xM7zvU5vJOLHhxXtLZpElp4
jlzLJ0/IgsV5SQN1eOK5JPa7Yqx1/chONtb+HzUR0Dw85QTVVnhVz6vjj3HRPKOu
YZ6vnpibX0ZIcY3QM8/yfaXBxZRaZ3pU71sQ16Sm2Qw/qvWSpEYfihvTq0VRIN9T
GezhTzXL4jCaA5c+BRY1mUa3QCddXWhqITGyjsboze6xLvkcQXyljN7DJvkEatFd
oWV4/2OJN6gylZvjPf9qMryTqOXiYoz7AIKqtx0gHYlczKqiIa9DoPdLl8uthfoc
QqLf16qLbED5Fg/UoPXrvI9QjTPE8JMwa5+HG1VUrEvIqfZpjj587RQ+7yCdR/ZL
0cqXGSNvxNCJ+KPDi0i2v5vAlJojBYV2lC401l7ZysDSJzQo9x2ZHDUF0hSEdVC+
On+/culFxAma0OZ1K4Igo+cZx1wvJTMmRp9kvIukf/WquxEGZ2cZ1PJ4KhUJc2cP
CvuXG9F/VlCKeyafoorN50jh12LDSkSc8NbDqhXiippQ5MfwzoAfsfVA+tqXocz0
D1/oJoVl+aFL3VMZRLGlGBfB3w4Xj6C6TJoYZh6Yffe/HP71R/kJ1fLeXjhOQXBq
DF8wBHwqEhKl4bWi/2Jd1euAcVgRl1Wj79qGx8kutJfFexTnUZ9MBrRQCZWfQfc/
t/QRij1WR2aojYFOk0PJfH3RFGV/Ityt+bKkPrlmHuW4MH19/uqN4KL8f8lsIech
GEN5WbrIByaheq+uHflCd+Q3ZJwn+uYu7Lz2n5xS65eq9Df46l9rQCzOs2LJZIaN
T1JDr+3sNDdjycCtIOEi6qsKtoWeHEExbsDCrNIKlijfbIKYAKYUPapcqWi3rgI0
ZPK+OLCrnodcgGZLxP7Ai086iBF8O55xrdWmmxfOx5WjklBk2eRz7Q1t9nzPxVE8
wewrtAcuUkPgsGwWdY2huXaydtYBFTL8bUJSPBq1ks0tyPTu4diFIFo0wG8AzFM4
1qIjxAGCISuHck6nVX0vWx9Emwhna8hldpzOdydwCUawAj4l2vhj6isHq+Ejq6M4
2wVt3FLFVHJPIjoKACxlIyz0LvnU1qfByiNXx7g6bQr3aLlhWh/t2HzRhuDiLY53
rtQ0ZppiDSyoqPLhF9aHzHxFKa/s9zXAKHEYeytfN+1CQ/eKojupMgxYyU85W+kg
5WyAcDC555n1HMY4Bgq0HkoGMsLEOlj4W2Z/ATry5Bvep1LtjFusWcFjqxXcsl2B
8SgoOh9Ebi54qkHEVGXO3Qsuqr4G1Rmdbi9fPMUrJ3VuBv/DIPDWz9UAoOULP49E
vPXgVAd1JFJ3A06OIKteRE8Ht9nS7hFJnunJN+IWxXKiCYlhqSopdISHfASNmNUa
k0iUrw2fA1UCnCZG2wehXlZaf2N9lblGQ9OtnXz9Xm9a4AZ8FdRPvxyi9lBPzUgA
9VWzItbD00kq/6zVjsWQhB5XOfWovBh54F7YQ5lHFOgBztmX/kgXQH4z4mqPuCwu
fIHuvMY3kkQd3wA161dW87HOBqvt85gO8QJ/Q1w6fajrHGtSCQXBK/+crLgB787A
1SDW7r8KJeqCw3/HrTae6YiX1BagQ2qOKCP0j2P+o10ueewuTUU6xbdcm8KDBUnr
YL4gJBmvlr/NqW+Y6SksPZDhd7t4Qa9etiULmbvMie/dixShK9Ihym8KZU1+nvIT
HlSR5ByT1s+wpvKT4f/FEIBXetrDh93OLdD9UiPWVdj/YqjQFhSDRdQiVJClv1Nk
xhjjBMm+VhvI260aOMcOX+n/kmcpcEwVVfbmTVtWTpy6pTPkk+yaoFZcq7XqiYXZ
lyWpgC83KO6ZuSeHC6YvMe8PmfZ9Sm7rklxItHdYauzRPyjHa/bD+2kSOSpceAOU
7olOTWy/NwOMjdDDOtn2x3e7umhj8vZPuegHoZXvSI+qNrPyV3Wj6a3eVPkeL5sM
ZAYuimyEya9EIgYx5nEFMTzVxSOvLrNnWDyGdo3N/CoMHrgHop2R70oqkwpxiKN+
bwI+qSkNfTSa4mGQnm7utcFecRpL7R38/uk0u4wcNuKCdwr2lzNZxWRSVET/BRfD
TYtBZpRbt14SIc5QhIo17AzmOByF2+cUR5bw1dpG+G/3jcX8jOAt2w5J4tM1KfSR
jCsRIPYdE5WReeXyHVwY6kYguGN52u1UjfJrByJrrFFKhNl3Wj0rp3RRLMRYCsOZ
ccpu3B1tGFDi9wuf1VH0JnP2FCfvhdUUEeMoTlebi1fFTHWIuOi5JDc8yhoGr4Mg
EL/09QyjhhMK8evpyIoCWNqlSUp+8IYmleI44fR+Npn0Erjq1t2ZXssi0pZgqk/B
sBAVPzWPjoMWM6XvR4VbP+QvlCZmUGhmRxIDNm93DQKChJvT31mD4GvgvYkGBXzU
WWPlkcp8s1KuQQH3E6KBWbk8/WYbMOdZUreKkLb34mGumoqY37pBFau0jFhOjF73
lk9qdBW7MOzjRS3T2xnZbgMrf/ynjreMfYTCEuKNufH86TGnnvjBkSiqrabZri2v
5UvgA2YUHE2RkifFx/KxuXAW/o5OJctRnf44KLmTzf4/JQ+4KQOCfJ+ouXWCkZld
wMI1jMIwAAxoHVatAmGKuu7WMMoZs4LQ/GZXNSOTPy7uWGdFDN3bjD8jWYES+V76
KOEX7/dP1EEv23Qp2TFQ/1eT7b23e4NbwWw43VllnCkNrHZ/fAcZDKiGsyGJ098Z
Gy7po8fvi6zNRIDxBzQqnkHSlKJjGufQFvaqqPYyVe2g8sEslLkOmItHJP/py23/
6Ps4ZXlkbhf1xH9jcwjoRdynHuHvftI4F7d5hLWOKXlVdfSP3dgx8Uyxoka8wk6Y
9Ja7aosBYOc54Spedvenz8v4yyc2jzqf5zBkjmglGrTTQ8eOZgZFVVhYiz6ys2N0
TZG8uCEN9t4hwvGBDAxh6n6Fm0bsjOIqQg0cPA+gW23fEkC9bSVF1GsgTDb/UgGZ
AgCl2DtbwOToWWY8ym2QZo8xUK6bn++UROQ7InvjUPpuOWlmhQ84IvkQD//XAu+q
s2Co7G8iRyapZLMqR/WwXqSBv5ShFuQNeiI2WtV+V8Muc3iok+dg4mj8qzJmNmZb
dUT52NOow308bwa9pCjxpOgTyJa2tLGIb8B871Icz+v8MN9FqYMY/CBDJ14BEpe+
z6wFsk9pipwiHkXkvzWe8XqAqa81eONtFgXCkHzfo7H64LHwjoJ0i/dptFMVvuRh
RGBboLlv3w+KFr9rbCPe3nNvfVJTEwxBm6U58C97/CLW6LNwL6G1nD0QSrbgnCl0
tiieLRSmMv48iuX76PE7NS9Sy2z0lALI5bOcB+TfhHJbzKnUUowSyFeoMAlXLGbp
/rRLwPVuE9jDCTJA0TTzfJze6s58q+kwgDkWqcxTEuBnKfi9A1lVXpEN8574gglN
Q16Em/lRYARrn2S+3vVY8AIQ+pvrt007D5plUHLWw2sWr1rOUreF+ca9fqvn52Hd
oeRRLjP+yyc7zy6njtdmDsR2WVVFNFme91NTJpDO4ZTNESz4Q5kWp4kCY8Rz/EdJ
Cgf8kZnEQ1XPyJ8+PrthOY2ZNG/ODLaGbWXn2DbMkwkWrZbUQlyLYnvvxvCVhFQ8
WTbHn0uXvBbrlaB7ng8Rdm5mCcvyNg84fKdN6emAfLNh/LZW49t1Z3BbxiMbMyeO
iWlrwv6HSjy08AQO8pXV76r5XcK1JRVeOr1t+EP+qYkXeaz7wgdPjlqfLmSBxau0
6snFw3meM6idp84X6Wi9N3EGdKXUoZwp17NI3d6qfjUEqrpTND+rCnrW78UMC/Gt
zBYqiClP0IzEmN9VwC/o8UpkXkCHS8PGpsKvGVJuf0RfvD3toU7IoHhsj2dTkk2Q
c+Ls2FmZKeIxzAajbEofWYpJI0KrGqGaJTdF8FcQlVbx0sONHYDkEI9Ce6Z3zAhf
pM0oCWcUxZp6zBwr1nfTlo/gk5cylWy/c0fqO2xLqmQbqZtjLRTN3w6ffmjHuFNV
A9n7pacKjuVBvhCcFAfWNca4Xsj13UIQWFjLkRHZQKit46H6GJUxHGIDC6jM+MLQ
MELfgmIKjBZBkvFcwqytaZhU5hDduyCg0V1QXvB+9yCUfeOOJv/1f+FdR3+vT+6r
PW/vkCI7NKqHGlq/1vOKMnyBU72deN9C4suzd6yoPghPJiloXMoMVNJ1FDFaKuTe
ZImsZ0O9lY1bV+XpfRAJHS9uNdZdgzMbtBEriTLJmBmwDtnQz1xdU/sGVV7HWhOG
RTPyc68H8Yq5Nfeq+VCsYhnJuVahs0bguvriN77BrT2X+snH4zPq7QLUxKwWH4bZ
9nAz1ZrPCnyUMido72dH0rTqTxLEUXad9MimuMEYQ3iX3S11XRfoM4Sc6qoD9U0Y
Yc60W3Pe7bMABrfCb0sN+CBaxQLUbzaA4wOrMludAu2gQ25VKzgMD9rzN2bzUh4e
SY9mWOFOMJf1AungafMho/1vnVpE77OeDIkJ0HxaTGHEEEYYNtSjZPUI/yCk6Rvd
MqunYLga5rZOHnNmgep2MsRk7LvLJFyQWzPN3immHP25txh0m5paLukt4QTtUluC
fKKjJrtaAjgdj4W4WvxUc/GVaao9i5FyqQEQ9UznFQ4VVSva2ra1X75PsBiE2xs1
9lg5CdtvkUEaJwY4pxbRt5j1Sgrom8vb9PVmg3zfrd/R9tVXaoLQwWmK7zuUvdhg
/vhlAXTExGfd/1Vuw385yWdrJopVeqsVqk8CX7rSvdNlUmRGQ5R7iO3kVq+7RS/s
vqcGVw+V8Of1jAewYcdCO5OYvZi6VK4hZ1lsa/9lTGekXzJ4Wv7Z2cm6yy9pVCf3
9R45zM7kMUlDYv+L0F7A1y2rVrl/1brphUpiiQCn2GzKYvNnMX+eDFdUjv/nZj/Y
o26jAU73lAvjaGas67V58aFN7ohK+hfcjQ/7C5Lmg0JOk7BoqM0cTurSjqwopcRy
hr7FKtlG33UfAUfsdzCOCbUqHoaRGH6AlD/KYtCoIJExgCHi/UC/J/UHcdhaOuVS
+i9LEJMEBI6GjeV6zLYUtBB4rAZX2vasKc7pBkgeFxrUvjO7br+0abM+NpaeZ3p3
1dOjxjXVulVDF6pgyjj6nRyiw+sPe2iAhztRtmqIg6b+ov7H6qszZPqGN6aVTfkf
siRDEUEV71MVBxhemEfh80DWVcG293uc8UyIXPqxMYOSKXyX98tkPDnY2bXfFzZj
ydvUDf/dgJiOnFmh0XTzXEFE3tied+Z+bjk0cFKpJMElXAgV74Or43ucub4yrm9Y
PuK/Nz8HXAeWBLAC1JFCrb9WeiZtrEdyRwtycY4nTL/fHV0/BJXVEh5Kmp75uTeW
y/s8O585gqhavbmDpHW+FbWQNjkD/X8RjeDeSsUzANoYiZtyVZrmtGI06x3FUkJP
/URT+hotO2/bO8Zai35mkcuhk5Pvd7kMsPo+0kSCc9UGkAsUasGtYdoJrHZX6NCx
tt/ZunXg8uMKuSxKi+dLj0AII3jnnWp1pR0m1zGdEGnUAsv87ckJv/lwvlrJoL7/
jOVSLxBkTue4iXqJigTnBfmE0zyPaugMy71eva0DWZffvl2aubq6T/oOYUL0wxVe
PP5kd7wZJcWi5VDYReeQrzrNwXtJ8NEcSpr313vvERVG0bb+B7ueH6fmXpWgNcqh
G8fJuexKbaLNji4YjHfBTCsYlJfKW5d22IxaTmYgFTD63THBPA13QPCoI6Ohdr1m
ietHZ2iYu9dmHARDZ/Ov8k0M7Up7wLc4pGyocm1/rbOqwU/d5JeJ9G1tzxyM3RTm
eDNFwWMDh5RGdvw14cjI6UqE7Pia9Y6su7K6I8O5B4M/LUxkSVyWGLmGRS0TOJXG
261O1X1NflpV1MdTrZBfWFB+znaocwqJ7IGUORMmtdvVZQPyJp2k01Q93amcVkCW
qqFAeDY95dnt+OHnWPexv9tylK/13C6znfbsDOYzzrRZY7iSwTTwUd2PSsiktswR
WH6KfaJ9Bo9JlUiAKDS+yq2zxwKXX00lLtExYh8+Cqt8eZidIlQtKTzB9qUUvHSj
EIaK0DlNcVni+gnKiR+HoESqbUIUsXqTCx8FohsRwtIexSIgCLp+2hvb5g1UodVF
okvlhY8aoEYOw4TEqNWZxnbOjU2CKJ2Lz7P/90jozTB30OJcfsHhRdar7zd5KQbb
7MGhmf7EVqwzMloLwXCKX/NGTLyAtm796ctIhzcsv7Nm8Kwjjx5CpWq0NRuPoOLg
+N0ZGRtRiUkL0LelYwoXtT4lw1xlpUo8dXa0TLtbryT0V1JmotBhCySwfQEZqfTN
jZG+gRKmLF5JrEfl5ElHE1pZKvCR//Aq6xzN8r/1VB+RWTkyOsEZWPNMrqQQRIZV
BdtXujs4GAvpZ3PslvNj3jvUwswz6AwT+0ZHJaGxYGIOYZPUsnr81Ix9nGFnf8XM
uNGUwOS8srNJ+gDy3SEvrO7clDbYBQ0kyRfFzNvUWG7QGqScuezRUXZgn5yWOCsf
tlIMuvt8ahNxM/4bA9TkHETodhIdtbxSIhy57EZ7H4RLepCHkC+ETm0UYdQ9nD1z
yRWYlX5JWjI/dHsNBVEa6mdwHsbTVfRZBPQX3lG4d5pbnlEvc7+gExVFY9rmPdZA
Kt4QguKLKstzQJrmE49ZijicRtmRWCH52qSh0pEVnulnRmAlLqbXff9Gu+C+raB+
cZQcapnvKOPd6fDoC2AsQWra9eYAEgI5HhC0mZQCtN/T0PgShizWni0pQiY09qWu
sbuWoHVwzIW0oijDlZqg9ojDyArWnWHrzl7BO3tf1K7NtsBLxHnfD3ZJk20ZQasP
GsZPV7ve6V/JNyfKTF3G+soaHIxG+sRDjj1R2v+I804eHsk7bjsamrMjeRyoSgpr
FcYGWQeIh1kn+DGeF2rnDJwU5TH7KIqVrFtk0Te8mH1UNSZ1hSGny8Eq3pa5SxeY
oJ55t2Bs/ChD0zBqpPxCJ/Tr0H0ofD0SFVl5GLVxzTW7YkahlLipBB8/x9dSg1it
q9hSOtAbC5SPC5Nqm8WX8qzcPGtBi8Sq5qN1St0URRx0EBfoXps90XaXB0u462CD
3NFcOR260L+VPpFCmheOZE257hdPqExyeJaeVTadblkXDnNEZ5/QABunlJ9gk33U
i1Qmnu1ZoIxWOa5O4I3xrVL1kAo5l2FrzXXiJXl4N5pYWPsu4ESOYe7a/lVXOLIZ
DZsl9W07mOrbiIR2HJ12UiDF+J5UcWVXb4y3v/xS4WFfiSTXCFWrEUXiIVC5Fhdc
vgzTMdujXxmz81U1gTlTj3jDyIQK1SPTq7XGM3tfbrxrJTg6x8uigDeExCtJSDaB
4sD/hAS6ut5LDRI6EbUHIxrZa1+dSl+H4+O/Lz5PdeCWWgD3RXbbAaZ90LbeB5UB
bbJPxMtJ1L+z4nDyXuFcEQFVXDu6nqQT5q36Qr4QStO428jhOP+bh5+GURB5Iy+C
GUgVGFGFyXI91y+e6FHhFbDxuBuBLha12pO6aYoroe7T3y2+gnURXsn/1h1sdi+c
J2aW04AUFshn2PTWwvcaZTmAU/bFnJZ3exJm21cvGFfjAqW0GAz9PQQ/ZtsBH3rA
cvM3xFjR8xB4toryrW9S4/4kY8VJP68MUn3eS2U5JVHOQVrlMuZIG8L51uRyUCsq
UkRWeEaV7IJowExPEYcatnRAHGpF2hylhq7TzYT5DEVEIJdP/fQFvFLZt/46X0am
SDl2UZDwR9MQdwfSMLFnBQHrAgPFKjCKLmGwAtxnA2k/EMFGk4U3PP7ORV97BAPx
cDbPsdKoKe9HH7c4zF2Rr8XqtYqBFT4uP1klKfeXBZxGBZkTCTLOQsEG1l7lttCe
6mpc8CNYf/sssA8barXoiq/hfbgGfNEpJZToXGRcofml6mFkR0Oc8nYifXNMXzM+
ff/Z/hOpH8N4sRhbk9LkOJC46/aPNugGZVuIki0gf+MgTgg66pci58Uov3fTrQMb
GjcjNmj7kRoBCHhd9sVtuxFE8E0Lnxdvxr3VVmMndf1cY5oAGcCLhfTpgVusMlx4
AMwrsaYupkCdeoxdr5cSZ6R0c+cvYjiLzSRFIBh3s1ULoq1SfQdL6HBtSSPo0/eY
mfDlDtNV5fcS5E1IoR8New+4qgzgLWWhpkD5QYnsz+0o4DHNikIvMXJ5A6eXbLVA
BrB2OgDJ3Cr1T5yMuYJuecso1ot7KzG2XgX90TtylXYMtwqXZ+BIHDZvBkl0X34M
1glkOZdk18m8S/yGz22asV/TNwe6iTfSOe/Qfd73zA7OjvJfV3klPcnr6h2xoFYc
UgOiQvjM1brfWbmHHCXpVD6FnzE5UnEvuhM/BDSJiwmFKEmaFNOQdNLrmcflzmGE
8W4Qn1uTncioxHhUWKt34xBMpNznJozBbhCw9ghPm7eMW0X1cpThxe3GMLhFhmTc
zyuH7CDS8OdRXw+S3TX4He0qF+/0Ga+unncZl/BeB0RAnLH3qrZ0wj1o3TDqiQfO
s0JL0o6VOC+5Wx7nK5Z/yywnnSoKXI6TyzJs/en3VIyTi1tTNIzNf2nGO1NP1Uoo
hjgK6CaFk7swx9Dc1SKD2JONAicPSRnZUkfexwcCf/5xu2QRjQOuBLy4YHfRF9lm
OTJGw+A17CLU1EV450SSNrkYRtbOB1jq99N0LRgGqMQNAS+YgOb82azrkDAuliD2
P2DhV8X+bUN/yCDPJL10cg+zCT9sBMamPmep7ofsuWZ6Nk4XIltGZwreck7KitYh
cLK2Nw3QGYK/dhE/cv/Mbb2KW5QodkpsCPbOdVHLlTZGuncSVgSi4mc1cNKvRcfz
XI4SifvmQ2bpPcc5NR9L23A/hy3S2wak6QwtUFBOXkR2ed38fbsybZFjLeYomTuw
Cxjqp7grWb+Om72HVSoXvYDUupJB7F7ShdhfXMkBPjlG1Y5DTNpV8TFPTQ0PXeg+
PnKygzgIw3NC1XsIyRDcG6EF8wfIAuS4dMN6wPzD5GAgibpC6Yqbt8eAA9CaZrue
05FpiGEqtDQA1Pdyr8QZPKFDpiLXNg9wQMk2HzPCAHScVxddsI2j+uhw7IM53Aos
KlHYqj9wUIDTlQ3dbCSRXIN+et3aQ8mFDIPx77kQP05P5KrPQ+6zxzEA5Idve1sB
illl8+xMkq3z2jTZ3IdmOjuVn3IV82hWCp+nwKwj9fx4X9OPgXhO3E6NM/nDHuPA
VJk9q4SGvfa2eYaMH+UUwvwcAhWVbGo6OeEGEv7tbFvqe6ncPOsDFEhVi9lXuk8y
QXMJ9aXc2NvTgrIlYlpAi+6HGPoLxioKdIdyxTSH2RDOdRf3Ee1oauArAx7Yk7qA
QldsihniVt7FZFL/c3pZcRaauihalvYa3+wIa74XCKWJ2zwOUPYaGQ7q6RAK81vd
cJIHXgTUhCP+xF+o74MO+YlytdZwmtSm4ZJcrEi6Bx9V+b2gLQ3v9cvkkEXt5EZz
DWCDPYcTn3IZArFQtZYpR38YN7df6xIJKYFWWPG5AK89UCefOPYbnBmla5oiUqqO
z/yI8eIWtdxLJRoOGN3w+BYxTUzJOkWw+RjV0teoO4EWsExTtOm8d4G5F2hUOAI/
iOsbmVv044+7ZReVLu3s+y7baBicHLhIDEqpjNGZvRhqDjkEsqiISe4P+K778a0H
tO7LPDjAxyBGJJOfqzGF5sPXdbMZSNTrnPbQRVV8hY8qkY+FGoLoQgx97TSD56yr
CLkH6kGBKAIg4c3WNkR9W+/jxhpknxFMPvzr2aHx8QotnVcDZ4g0VUMjvTLKJ+W5
cqwPLAzaIPcmmhOQtue2FHEE7JxdkcQOVOJKbltuQUgYs9l6tRV7gTL1HjY+rH0u
88gpng36KFhqgoqFTPE80W0NPN0KXVo+cH74T1xK1rXs0X6VDfO0/LO7eYZTjqrf
7IkI0dvqP6hpMIGoDcuXHQ/mWoclOtoo0XQK22yjRG4fgaLnXAaiEPXXPZTGjZd6
0vLB3TOotJSXYFk7jga4UyQvkVbZeXWkS6JWU58ZZ7Q4yWDGAq3t6tPkkKTfTRGl
3lmyqQSllrdfChmOP8Q/zPX/XloTpk7d4+wcwbZLq6pNh74b5PGada7JnnP5+CI3
jt2OvcFznnMqVr/G33tQ7BpGPqQxDnskycSZesRGc7YmEF4e2O3uEidwXKSYbeeH
+QISK/tDe3cigaHHSVsz1sCgUvXnVe4cSVxXA2r65pzAa6o5h0RuyF6snki9JEfU
j5kSh/Z5CNTAXN98iuTy4SorLnItDlvbo6AFCsY+cN9TjN0VbNtwiPJbqk7spVbZ
SPj4wgXDZe03Nb/GkxuvbaHEScXwbdNETx6LaVPGykQTRX8oaDIGOF1slKV3l6BL
b4QHqpJvuFsj+w8UxrM3INikj+wikIPgH+UoXLfXWGSPuBeuFT/Fz3VJVDf7CsFJ
rjVxmBVyVauMzEAWlmN/+EXQN2swHiRrJcjyXyT5aR7IUWGUDSeK3irS+ZfR0Plm
M5+RWB5NduK/GMvufl+50kzG6Pe2ATB5GbBNxMD18rjCanVyVYLj7/LWfKGLQCDS
PbF+W/iSTBGw5gPgxOdJGr3rTNzw7wSTxRK5KBmZKG/A/i9QtWlyeWeJ37qPzVB3
4ycWMJMvEzH+rdtR2ggWz2pY5IIaJOsu0H1rnxx+jWIRYDnHQU8bdrd9nNlCpC6K
4ulQGGLvsq2VYJ2GqyBVCtlVFE0hvr+g/kMWdO/sr8D07/1ydOR/DukF5IXDbRDV
QuHLO+kB/yYAOmDKkwDDvaCCtQuFaC/6ej47+oxSNd87fqbLtumIDGGzh+gfnov0
Rzkbp+SIEIhH6xPnvnQYNYgOfR/QJRjCJK3Z7JPFeVcfrryUkrmDkhf22HroUyS+
PtYgM2DiUXnmUHPHB04ZnOHZgo5U9DaQ9NKQbQEignDQ2I6C8HCNsR/A0dTdvJ4Y
4qGf6a1CNIF2D3xFhNJXevuJvyto/qi0DJOOekHPpvxcWBc+zOqKoI74ILqybjKo
/HLuATwBN4AQV5K+Z1WOmTBpoUSQMZqrFtY2RJjs08nGB4O4Ez7H2TJ89EmH7f0e
CUMjaOa4rOzuS7PYM6xldnBundrnWikPztqz1csTkVtlvPYQiqGg+8orR7IZ0ROR
4urvEfhk0vbNxcxa/U93z1vPSOhdvSI4+QjJ2/4jBEYeJ686rLQTD3YZsX/1cMDC
CY5+nEp7se4Cwm8f4NT9rARGjJKi4FzuxSJ6jnwbWaWUysAjPupVTMJ4Pw/9MiV9
BtXBHgtiI7irmBlDz66h3ptWY7G8uq0SeuQZxoZcWAnHoQ85P/Bc1kp7vL48xZiK
uCKvQRaBZl2j/ifBUxX8JoVNTUv9FGp3ZzPQ8O1p/lw0jAkRkjy2wAXWOm2poL/w
Az2Zou4CMMxjMNL12dB8qbwvdOLgZy2rT9HAw8EQgWwk3IT7uhzZ/rCMRKlNzTlY
KONhyURC2ZhbE+FmgaYgiIi6wRoXX5NsOPI0UJsIZqTQ562uQpDnWwUUNBv2v+D/
u9V9VvlBYkrb0ix2uhQzj7JFb8crpDetLMFtHjYUZwk3hLv71Yoa2mrFfT118pPq
Iv5Tgb2DGu6LF4/n4sd/2R+G9MMye8dCzTAEnIwkAexNVkjw+jEJao6mKqEGC2FU
z4LjCwPPUnJvBRZj2q3GIAymh44ZwS2O+qZCVX36sFnEDxMzWOuqO+fGgwVtPLEs
xf/AXJWB0Q/QG360Yo9u9+SlHoAUZIpcaHKaHJaMaRdq8UGBs0YUuKw0LeQrwYaf
9OaJUSFIIeRcSPW4R5T2Cean2TiitLUEfQ17hwGf2M//L5ngpmgrgPlSYRpfwxwl
xoK7f8Zm7USbrrVKLbcEmLh67aFIfwrjc0bnGk3JAn4M4nvPZiszbMxVKBo/ayFX
Q51EbwBB+Cr22nr+IT97cyqG+kji3LSqc/SzWzyNEOXhKhAWKnSef+xHOJ2AWF3O
ZMRpxVmBUZuYPZNrT3DQYuGas/OeMkRfWVfQIM7rgMN3QXCg63vA6AAmgBbjkzsF
D7MMvzsA43Ksmi0pO4FGfvQM/DrA9HlxdeAdlbj+n0ceWJuIbPnW11h2p9zDGZuP
aXOF7FzsFwMVSKKzVQ6fH+0mofeGpNHvQaenuOqd1blWL6lW5LolYPUYySXS4hfK
j74ZDZBygUvXv9E8Bre77zO3ExNuFWuC1vT6SjRqr8H1uWXuLuvigv7V8kttDy1H
ViRQoL2mDFwMinoCJv8giBS16TuU1x60KXB/hhz005vIdckmGTwb210T8cI1zFUB
dPVY/QnPUgQMugp58j8708M7OtuCoIVmZ0e/CevCmVoB0Lfpmh4m9C+nEA5ufwC7
nlauWfYc4ov1iJO0wtwMd77Df4RCFaPB7lt3C7qfbzqApFdO8znIE5vlo3sAM3t1
HYMPbtdFVOnJ1rrqZ59eIk5cAXIajV09RPm20yZ9wiCOdIMRhb9nHimBazK689hT
cr2QLb58crifU5Do1leTFqhUFEPGvBUtQLOBNOFioPB9fqgFRVIZMmJFRRIJWEsc
vbMig6bdv4lqOGoGofvA/O+ToYIBuElnPMD/xaYShuUE6Yn04BnyPjqwOe2hZkaF
KtAsw1bp4ACI5bPmhg/5qPc//B9YbuTxdpe0HCghKWluVNCVTCfVywmTdGoQOLzF
uoGpO+TriK08YvCFjwEicK9//J4EW9VRwPm2fp63ezz7SlZmflcDAuw91fMTUIG5
V+W3QrhwhFp/YOU9TWRszRTadGAbSV2drAPd92FMM8U1JW4u4B+r0XiFx+ZOmIFq
u9uIbKlh7jJwCfsT2/cJHSy/nnYWEB+ZMF10ALTn74MfLRdst+cwGwSBowHkWzcp
w89GTh9ZssPVDRT2Wd3lC22eNVaynLi8KDw7Cj9mMI2VhtswPo+vtDNVtGevX0FF
dQUwFsR5I1fmIGYgEt21axVSJdUp6mzirdnAKFxUXmlUauzKyGPBlHN17I+7CojU
2th08mMI9uuXLEjmAlQVp6ak/59fm7oJiBtSV/l++srb5vQKZSav+MSt5rRXLa01
MW9gZUPUrX9s49ZKoDxk6re9KX4NmGe/XrnyN5D7vAk7tg+lsz0pVNKoh4dgw1H+
FQbgFacSL7ewuvMLozRUOitVvI6akPAEHzo53G4VwME/WgbkzPgvpkI2zcQITc21
/LpipNFNFfMHcb5JkZq8Y0SWJbTrXUKUsX7VKBoSuJPLlZcqQBl4hCpkoOC2j2YO
QhYpC9rij6sIDeYufXT9baRBPeIJ8ARqQeL+ROWs4cU1cJlljJMm2vTjrST0D5NZ
Kq3DW8x2BwlZj7zIk8lxDzQXbEWa7sB6bgRmIgwr3x9zb8GJ7wi7kYiVjdWrrmas
QTvKQ3GAbTzcTz7ua3gjNKwyHMR55KJG093/c4+deOByYJIJTU48dGGfFduw8ntR
mrXFjSFcJ4yByfSmke6R3cr4ipZ8nLM5a4DPB0ocIkJUA0sxP+a1P1CeH3E41pbX
8CVDkKw58EGvA8qursD/VvrzVVNLwdtY4TPNnjCDcEEi9feEP4pILxooRTCszW0J
p5ZCsv3TeXsqFp3OebSUgll0ZuPQ2sbun7uSifKk+FG3BfQgLx0vpqfScLc6tkKU
GvP2kj6YwmWkpdtCLIfj8jwgSa6j14OY/kvNjFfxUZwiKWBhAPRwk06cIzDEOc3A
dgveFam1B//nsJOoRiuByCQbGzDwlEMvdjIpAPokAupPyDfLfg9vcrZO8HZ82mwe
QqBf1au4Cs+BXCN7TNdVsR5hUBxHKP4jGyp12mtkG+ywe/A2IZ4bt9qDlL5y1vYi
f4KKE7H72UwM0CFAeNUwu7k4JouvkHeIZBvA350AuGZpNMSdEkqNI78Vm9ENEP6h
0nhr89iByLhsolBPrnPaYYREk2eSZ1nqWz/79ybEO9TBYmJhtRzniH1uAFszKZQo
2ok+UAnSXB1pRcIT9fBInLxsmz5l4Ij4EyhuRrfXvlJ7b2DLrSUMxVTZYNSYbxuV
iU+54reNDnSQZPyptxZ5Yyogsl5bHQs4fF8GlALMMoYs2PP9SNT77f6napm9qUui
fRBuuIiEmjWaXkGniXyxdfhzeKKjkAbDKZxFqmLzFIQnZpEvetHWRoNA3qx7ivwf
/LYbwtg8fH13o7msDBOu0bwZyb71OoIOlFmrqDAFfMNhCCogUGfMG5uY60QueguP
4HK5ZUgRPx1QwlrIj3rsMEhzaCXUDoLqiM1NpMcBdXFq7An+4PdV0btI4u5WdgZZ
h1cAyxiPxeZRuReQ/xwwFCYB5heHAXmfiRPlaOrpFL4YNT5hK6MRWshPMNywE06f
lAq/vnVJhg+JmaLgyLFEVbNnaZdYzDr7nd1hdO8QNAg0XXAIEWNFI3sK/OXQF/To
tlbaBGGekkuQlgL6XVQCUrI/7tK8CvAsPrT4vMKrG7TuXZW3QGm79UNL9rpL717o
lPlW0SceXWQWVPt9bx0wphB3NpqB69C8oC43wOtIfHUkJvlXvytzXWPH5Ees7KLt
7Sdw0+3OvfCOS4J5u/+qMGB16CP//3p95qPHgV+fkkwjs+vlHAEG3cYARursWsOT
MeABdCP/FBXI68G+/BxW89vk0J0zZSkCy8Yc9+gmHxeDz1KZv5GxymzAvBT0+gaA
KQ3GTynqddpM8uue9wWgCFwGmv8dqe0EqKKKP9RcARMLRmuwfDEp0x+LyLFVwQTb
kQuPBVRxV3vaa00t4g/xJcKbGHOJb/fo+nd5/b8Sq6FshLHHR33K7p51cmnYAfLV
5xIdQyRXSBhPPIJ4EDuvkmkIDQZqZra6jiCsma3XPJ+dmrfZfjq3LrYuoFJbh3Tq
CberBWnRx4GmbkynxtpYKuNkw7KYGHKSj2QOoNsGkhkykOwyTsnjutF7OlKa7B11
zRYCBD/eBhnKti+K+8DBYELUqusgmh/LyMfD7W6/EcKnRUNkFzEdksxUTHEmQKoi
EXRu7PC4RBPdDSDooD23MRbm8muFFLGfwl4DqtBmLR49jy82sA26QREgeCFp6a4g
Gk4l3rTY/6ktIVyD1FKG1ODiOi012oVgmhgbMhKxb8crBhL4sqQVAtf+PCkkwCgg
NiX9XwZ8pjxuxt72mBGGQGZSj3RY+v0+xAXbshEqZijbkFTqUis/yPN4rl901lTV
MIpSTNKpWZo2+EcGrM6yF6/gE/oU74JP1NILuUDVnkEQauzmGF10QI2CvOB1TN8u
gb8sOWBhn35+NdnAuw6IAQdHXX1kc0qBZGTZ7eOQk7a40agSctpE1iZI897eXPze
ZsGeIUAKXlBnCr1dNpea8Jj5P4NI9P0whPN30uYc8X+ZNs/kYiPa7h2CBjKoun9u
xjYXOpl1F+UykQMFa3kxUtbKnoNrSW1vW9W4G/YVmkTVN4RYUA3mH5ej1ue/VNmS
egoqLOaddVzw83TxkhNOsSHNCcOY/lYppBCnDxP7RHxry8Tkpkdq97LAwtkS+Phw
7oj6TV5NKei9b6RASAGJwZPc79kQIHLa2IvRSVn+en3cjreOsZh6APmsH9CQBngc
ZH2m27FZEchWHKgy3F9bMhJP2idZozzZ5IRYBineb2cq04F9EXBQ+EC3JK5BLLGi
1xH/YQ/sN3o3ybS8d/RzoBkAITcD5oX3A8X+43UlKcbqNJ1CwZclcQr8bSkPoucR
FavdYJ8OU+CqTyP3m/PhpQfUVsPw6wPTbFKNaxOCrLrKuFvUUya5QxgYUAtbMcSt
mNuSWD/8T2NTsfSphZUvh4CiPCrd9ISiPf22g4ujDqAG0cziAKlDvJmTr8EdlYRF
UY5R/k4sDuwEdli39AOhJNLAwnsCcX0Ib3JUVi4QtKeJ75JxMhVlgr2OKJ03kwO8
e8phrdx3WuvLotAxGWSdzqp89xcjfP87wlUdHZKFqH/IWVOo3Yp17la3y7Tui0NH
XyvijnB0+vDk8vDtDQqek+4d6xR/0CNxdsE7k4u6A09TGOBOf6K1kb243fypPvtX
vIaZ9tS7XX1w/+VyuoM4TfkDKbsMUrSbmMSFKXE7RCJYpu7du5PGkmTSdZfiPGdJ
AzrJwoQsGGBsrMnPXUbeuGCTIKNDsbyHQA3Kjsd0H+UMY29y33g2gub8Tdchf7TC
bEb2xGCFiZEJnnL7JanyUljYLFRjdp0in+7xZNHFWPuTXRaI1Rlj5Dmn3AkU38Da
zt71CzUfau6kjgRib21VezL5gl6rzVdW3BCL5/51/OwoH4j4ppxh6Lv3TGdtCCc7
+gFZtzkZ7JfJRUjnfmHMUF/YKL54zhEGTaTcrC5F9VWVLJCeAe+xp7NY5XHwXCRs
ubWX0DG8HzTWkVQ8jhqLwWFUJAUR9JVtfZg2966XzsIJb2ZCRslcgFiNfPxmKfWm
CkMBjgiRkStEyo72zZofsW6/nez5S2eBI/49/8pUDPs9ZaE3vwRSxxJrXwz9lmhB
FqqjsrsznmYyAo3TiJlOLvCF+FvEL0JM+lTp+fD6MMwFmCaVVP320HBY1gjnABdG
hC3EodirOzb92s9qXChXXBQ46DRq8TcCYnH/bDpweDzQG7D0mRNDwSNoaH/YkOij
LYtW0ApVV2z/tDiMrZd9t2kdKM4ixXqkE4H7R+/FUQjjhmRv77igCwf8NrdlaiTO
iY3BcStLmTTT2ZuFVmIMkxDmuaFllPTywD1o/DdMvIhoXiH1+/yddGBpmRSDtjla
4ssSkUAREBlO+AK1Ch2qfhsJW6ZBYtyeo8lh9z6BapL0wh/JoCiLgWkjuTQ4mjk8
BbdSZyl60fOwGRSmZRElJWyElwPzShDZJ/VuCAJPvKjIXpvHCSP2w6wLY+htRVEZ
f6Q+dUpcliEbNaKzV2Q8ccdhqHtjuHkuYmxpG+Km9OlPt5Ms4tskAAoikViVmFer
do9Ikavm6Yt7tcVc/rVgL0LaA4RwjKGNzrr1NGPBv2GU18PZAis7jwAJKSX/g6V/
u845qmrYm+o7xSbnGPX49ekFvJ1zdc2/RokfUYfGD9XtNFcJzK9SRYV/hVrWMHwi
OGZsvEadDsOR++hck9XUi3jxfvSNL/lBIB04q1oAJJ8LUgkCmoXp73xDSLKPt7Sg
7loa5Qi2IuhmvW4jvNeu1DxLhpwMNcj09NnevO8TVnTiazaQ5JiYh6w4BFuPs2a6
Mipu8CXNAXiD3UGZsxJ+AAKTc6lmz+eYz/uBLZHaR6036LLFLxVojJYrpvHjt3RA
isuT5eF43XgOy+QV4EAYug5FDjIBzKe/kVLfhsRzSlh5G7B4W2Z0T6u7ma3UXTz/
Iq6/T3N/m2iteixRZYP8uUjiCRBKM7RF3TQIltFPDedrdoMcDvx5iF3FLaY/AZIx
Q1uM3GVdNL7ftPMHflFGvSgLILbRoNDldfgk6Tr5GajWCqKCtcBGnD8Dwbrisu1r
/LDvema5jlDy6Z4+xMoRL4wTkA7HnwQcxjTExlWLK255ZpEhJFTbBH75YVaLt4fD
pcbgtw1GCyG8HMv9ycV59ZXTFetZzqtRTSp2rFndTrt2iN19ms6lGX8QOIEpg9ck
Hj6OVDUifwRCBAcm76k6HjkD0lmyEoUuT3qgcGbnGJen14UKtpbB4B2za1riXmZT
lEuArlBQJUMVsS+LfD1zuE7HRQTUgzFoYv4STeo/5xJWSH70yaAYFI0P1chBk41I
iGlWaBgCiYDn3VdMja1jIHF8MNaut20qK6y56lk7gnPmRnNX9pl7e6daVL/sciux
9T0YQnV6NGK/3Qx8r7JXquf3ormNmV4GvzMEPqvj0z5p9gnwYd08zupYXg3xNsur
oI7pweLMwzc7M0qjOKR+bZZXO9FHXX4BjWfmbF3Wh4LPCMBaRhiwPQdZ0orIJWrh
Br5BLaqWgjf3JmFd4ci/SQcqoGoychHPFJ8mUqBZgitUZ4JgCIVxQqZuiSELYCwf
mNtzNs7HDt8DsWgHAC4JRZYUVsOY/RGmmiFofGwM5+uq45qYbutTvt+wVbwvxhpt
mhI5iWwrlXVTc8H7ApLCiz9b6hHsN52XYYwmBtFwWlMooaXb2EsbDg+98DLC90xk
FU0RJRzlhAcoUm5/T/HGsf4uJ7NRa7GEspuM24nKwXCSnUpe3HJOUTLHNg6NThbx
L8As8XD4MH/RWdowR1RsyKiXh6J+x1j65yes0+4aKbJOObleGU8k0h21cqOnT+Wt
8KN7LlH/ZKWgmm5U0cqJ+dRgfvO0IKAkIrrHoI9Wu2tESd187ylUC3Hi5FAbIQEq
0B2ecMp8rHPmG+1E8MKe3NcKH7n1oTRwX1y07TYc4rM5d6WZaKdnskQc/oh6kJ/G
qYsv2wHFDeQOTIk36C+qanhcOSmFv9SAJXpxl0TGBJc4ZARNx4aW3Ii8l51dPlbl
chEoN9EnUmNDCl2juZ19cRWhbXhdILwTsPBTmKHR6RILUz4zLO6KE9wm8MWQfUV4
eR8o1/C2KqpOXIIRG0sDFAhiMbKYWEXk/+W6VZaIMEXGufGyG5CyJkYOiF7/1VDm
AbauVdzn8wo1r3e8x4m8X2SbE/cL+z5YmjN9GXjtuQ49S3sHCOgfcWRkwwTb7PKn
mrP+kLte33M3siZRS2VxotW6uq32rxGXLyGpW3IG1evtI2QPnF6AGKl3X9DPGXwV
Mo7vev4zGQMeLdVYpOZoNNGtZ+9brAPctoXprDIJIkwP3bROGqppPpfvIBujZZ6q
KqspqUeVxmy8skpO85O5340U9T4jhjW7K2DeMxqNLg+L/UjqE2hAWcIeGOeUpqpw
aorkA2PrzQ8umEyh+nAWsdUaZY9tcUmvtzuse0g5BU18OKSQ2gEgzAjraZ1qP5nO
EoQQCxGLGlSyKE0J1fsDnpOrR4NlE1eFjxfW80jfV04TeNkCrgdtHKGW03tv/7dp
muw9ar9oGONV/7pIyKm8nlDzVMfS0HNOmZ3qBqpAi5Y8sNSCu8aUk3a5fCDnGiuC
WwYb/E5DU94ksSoUHzLk9B9so3whdLiU+pmFRnwBQ0SWhPaYKhttCCbK8y1vanGA
uRLnCpuOi5EFh0enPxM+lbiaurf8jd4kG4QUvk80B34cuieUiVC0YBWA49SBE6IQ
6+OaEUKGu9OvKwrRcFxkJ5RWILfZ23rut51YxUub7sgtJRhfpvZ2o0C1v+W+i2Rq
OJcLYZc8LXPToizN2nKU59JZpqo87L1sxTHeoosGnfJMqsYCJkMZsP2BqX7VgFPd
MuUxHR5YF53fn2gftsl5dfIGEcoYc0QOqsSPEHn0foLr79v3Rul75gcGbQ/cub3f
hJicuSPxa8/xt2GcoxCGZ1R+nJf9xhXM81kF241IrV0EZlm3kQEI9m3I+k1UrQyD
EtAjUCUrQWARoP15Fp516KjrQx8z6jrsscb6o6DEMHQ/oNgbakgLxHH7AVO8mxCi
nBuYBk+wrnN/XNoXHmtufV65s6Ssk/XDZIYCQeNEtBdPtT0rC79AbrTBukvNZ2pP
Ws7VtBs7Y/SNwWye2FXtu8YHVhK0vunlagdzRxKyU9mEPwRGdM5ExjG/btHyyKyv
CYOWbZwMwi46FM6fPDmaZ8B1hIc3Rar2Szte0zj7CAyUVA3kPEbCo2IhH/WxWkhj
7hIHRnqGNhGhXLidZ2FQZcFsWx+W3QtZAVacf+67q2xF5PAy7ku5PuDedUeTXOd5
5zxiTK6EI9RYNt4bNI9ZsS+YxZzpH4sEbFSQt5FKJr39XUspucuhdqmH+b4FpypV
IdgJIiOK7JuXfzgRQlFFeAQGh2bnGhJZISXUbX6wfP30JCX8kw03vOueKzfgnByF
nxBOSD6Phluu5w0zsgRaLaZJo4ZTJuqdSzMQj2TXzfBYj4b6c20xMDI1Wg3xg6Pw
owLi92b3TdaPlSMDKNmTDPfLWPf5TF0sAj7O/r4PIs5RSXltvm7FrzVF4wWUrqge
zsrpsqkVwVCXe4gD/YOwscld4Tf9/8ZveRltUzVlz1PR/Wb66nWzIYysaZQkG1VN
cl61DroBrW1jKOVU4jDBKT2hzFBTWYuzdK0oF7yDbv6ozAT93uUS7H1BPS7JergR
BLkTOjJkUV6Oy50vrssO54RNDle9cO4ktCAo2iae6IIja4ic6EvH+A+wZfHTWlVk
hLdO3p4AtJNX1N0zQD/+EiPF57RhW2ImnIrHcEtDDOqDcNpTov/B7Dsh5eBHC9/4
HhDOVoUAzvDupnSslff+6VuvlziNqCnk6zo65ep9QL8duqpMvX4B6kLJAk+A28y6
r78pL7b803NuqNmlsYG1qeABp7G84GIhNg6Ln0GlBLyKOm3nqyfUgx5ul/P7KLnX
7/YrRICpx/xhZSOeapiNQ4wvidk4HVwSI+NBzprQYszsT2G0woYxpSUKEXlxD+yl
aKjUF4lDatsaqwjyzDE3MgotejB+qLa84V7lJR1UxqqL1njrDrbKzmuzUm2QcLUi
7WSjDccW8wrv9iPuYqoceWIlDFiM1yAxBRw+kcAguHzs5VDds2qd8yxuJqlqbQuN
02l2bO+rAnwaaHLNq1RfzA3v1KS7zr5oDoMPwrB9R+C2NkqwHzybFFNaq+g83WXf
x/VxHywdHed3gwE1QAtLquHSq7HGFqDgQjwZOucl1yyBMX/Ck99HijiDnar1EpLy
SKMGW2dMJbKNr7aS4MkOocGtbszyfGHhj7Pm1ofJiut0TvRK5gudSDNhozjMMNV2
EfIbMU93Y+KTKTAx3KLqpB1ptk7P0iJmT104eclSj/zwta9LIdBQA3GMOE2Z6K94
/9h/A3AaavJWXK48uT9szZjSXrAsbReVs6ZE/LitHhrjnRFPkDOZS4gHHLx6ymWD
PhmCFF3g/3EaNNoKfotV/Bk6Pq/I9qC7kQO86LUsjp++kcoOhEdQjg/7oJikCxVg
9MdR9ZrccXTbWjeYawBTD/jP9aoldSnCLEwWapcU6b00iV45PrZJQI6Mjj25Wots
H3x2vsZgyhM7LdAoKMUOwLZsOgJmq947YKfAplkjjlUOtFUEHfKRuhJ/5Qv8S+9y
8kkEgwNH7E4xHI7fRxSov1x3TCigjaxqioIKf8UaMfTh9Teo8JZzqDUpz4dh/Lma
vWCqg4PXL0mZHTHbuK6sJsYkQ9dhSKZz6THVx+o3N0qGAWyF6o23pmhrD4FfK1kl
JTgKeoBiRMxsHhQd/SQlfi45HYJ2sfkqFMAILKhvfeLJpWtgQaaSXfaTIPHdQkeU
CExzG2tQhFBlpoEn3JOUFr8kcPlCF5WUxXfBh2i1cRDwcduXWGlAumpcnrQPq8K9
zbYwuq4Uu/XF4szv5Ld3D4XS8xLgjR8Df0VDY5K22rKlUzwj2K9m2wm6tXn1ATul
7rA5ilLvSvH76xYkCbKgHhEeR0MEfg4njZ/XPfEWSUlEQgFp9Rry4tCpIJeJ+htv
H3RootY1RothW9LS8k+b4BisbAJqDXxRW992W4+yRZbi/JzNWtPh6KQksMpci4fS
+9Mb/Pbkx7TjnzCBq9/Mf7TIC9gBm5Fwx9SIkdHkOx2C/wpKNmfHhpzHZKDoAZ1k
au0CMCcb2/XfH8fB8nMGIrLZwoRKgf5MGbjjeSSQ1qGmV/FgXRrEfCmgv6BMhzSM
75svbobY6cPNUi1Xh2UWvYVjiXtaD8jUhjMXhUnnWs7UL96C0bTgJFXmNPriMux7
0H0p1zcAabFE/MXYxajaBEq1CRPrdFrCt03iheHSsEe1mr+Q9oAFcX0pyG002sgq
3cXWwEEr0GdwvmvqUTaeqXzj30jhJvexdHceeypDk+0TfdPE/aTTFwi0q1TsoA3S
vkQhoMezZBQ9F9LEwarAgK6CnksIBdgYQlIs8aBJGma5Fc1P9TTSNxZTAyoEd6Qa
zcdssjUt56rQA8RqZKaX9CPVqiixbz9P2nwBS9ihJbGT7fguHP0+tWXS8QrDl8Vs
QokpXNuXCXj+TFxwdod7/2jxUoCI2riA0z4s6c1mn8eVet4GZi6Q3vATnxgJwpN0
ohr49Ag3dgH3RSi5SjNIga25t0+NUGDKxAmW3qvFVwoy0OCGtEM+XKAmTB2T+FFv
eIp3gU76IoZLOpL/oLmRxJnNTC4K+tfM2RKzXJG7YLlvtCf+ySlXirSGf0g7Reta
FTGpX+0SkMTLx652pzlf5Hut5ZBNagfoQU6U0jQKEfRJyd/r19aELFdTRt/hX+5n
Ietog0XWPNtCtCiEJi7ymWck9pArY+h4i49lVJlqlIVIVwz6vRKTKsevV4Dv1XWa
qusFH46I4I54tJHtHs+apTGKhBNM8/vxjgKF+i9Nzr0o5TWHK1YpKJ/1BbpxaoqP
vG+UDlJx2xttpuB2tPpCQdlbUvCZJV0Atu/i7BESIIWAqbHE25mw6XnVDQ/Ecanw
rwJ+TbtCTH/xqfPc/cY/MIwNCbnHRMvhe9of5y2i0bs0YvUltRTYnfswNxsZYo7w
9V0OhcwVeh1nby4kucxW4+tCRT5JIclQZaqUCA+X1NqExP80JKnYXb0zAwMO0dPQ
voHGAjEutpDeT9knWN0rWL3Ta5UWZM/ZR508Nc/9ugqcSKLaob/b0txAbtTc45B3
sRmqACQNMtqA2X3s+SJzIay2NxLBdZ+nEvcxcEqc33/S9G0fSqhdZlk5zgz+K4Es
ht8TuikGMrSo0t4iQT8crL2v1y7X8dimVVpOk+8qV0vTEi1xRoK7fyZ0mcMqPUVI
H0h0EBlSz6hHhWhZ6DkgDAvnTXUMP7N2qZ5x2I1qgtFgYPWCvOkwH6xx8Q8MafU0
qOtaZeV0wzipkQWHBCXonU/g0MLy6MlHD+VDgatV5vXIpwNo6oz32AvHZ7E5ni5l
Le7D/7QhpXb5yJYEpE4FIff2VlAJjjozt6j/e+hPsjIm9tEaMgOF8R9Rn2kwyAS8
VVnEm7+DeywM8x/UsCYQ0YFGNsm4ElIxwnfYffXszdYT15gdC1yotpbhQsC0jBKA
vHRVg9ZP999rujNnNvz4DG249wde7CTZpW4axY2fP5QvDo62yQfLxlqmANGwLTbB
KG1XUtuVuGuV8eUR4W1BhGUsW9gkHfEH9z8m/MgesPbmAqq69y88P6PJ2aoHzXWu
zTc7xk99zfqklcm3w1bmXavqYpENCnCa3BcQoJO/TerEceKBvnevhSHORQBZk0lm
c/LPn+H+TW0+glX/XsvTS19xxIzNRcS9XMgMJYqk5flwmWp1+dmV0F0YYg9reeG2
w+hiXPuJG4JRd76/5+A2pU9N7nuJHBjUIvkOWARuxHoVWqtezFDsL9v55DjHGY2G
z133stgiw55+409LrJwNQIX/NAH1znFg8NJ65t588VTJ5qOIn7FogMyHiorA+7pR
9/ttEHZmNqMtPvjS6SvgzrEGgXKKzo1LdFiqwJIMTpXHpQOkuhencn1MB1X+h166
B1nWVkpBV6SRwRwEI2FwgqvVWrJvqCdhT4FKA5WOlHzDyvHPEPY7HrZu3P2BRF3w
JLQCem/Si35jehP+k1Wp58xFxhqzeL+t3E6QN9VlDMGFYpivZXs28jSIYpGoI3IT
AEVy6P5NXUd6YB6z+qsKIynwQ2LMgb01hI+WjM5s+oSsYh4mF66Fe0g2+S9kcZ34
rq6V97ryYdCRs5xj64c8DjWgaYvHDEcSBKGLRlrV1IxWBuIv4CN3+FFa73ehFwxQ
rKjBQqopG6Gj3lnQ16SyzP39cYcH50+uiIIzhYV5+omptc0zo6wmOw1sdre4ojb8
fWnrOu+X2tt8Sgjw49w0ko94f5y/E2sENKEIb2sBlB4T0Nh77mW1zHTplE2aM12p
JF2wxjrsS22qoA0ZAIa3Yz+zB8r6dZX7FJquxJ3ZrOJYcpOqT7c1cuKU/4sQYNnH
DNa8MN0/ajkylybPSwrdZrIbVZXkxjySnmDOBqmG5w2uoRjVVXwimnbw1+ExhrHL
xY2wgOadMTK6eAb/uzuQIZDccELN94jvdUbyhVcnMZbhg3QHHOCEQOQD1SChkgXz
Cud7YGSl7cTkcjgP8ELMpZdhM4pShNXlmEaJKT5h2haekqeLRjsS66VdS4nVjqWO
CMR98+PNi5gh4HUqUEP2R07jvhIyHuaHvB6+ithFPIasQ2Yaruw6YRDIjPtwFdmJ
MmvWdhjE9Qb0CO7vbpNb/4Zl+lYKAm5oGC0NHHcKDkG4t3HHGOxAbSF1yrlaxgdp
R+jWVjurTu/S7Qf+NVMNxT3dBLgX0j7z3UYZGMbXo4HNtOMYmMk+R22TvltuDkVB
8jntxk4XkycDHAEQvhflYNRcybQExgrP0/bQ1guUzvL9snpgM5Mu55BsibbIzetB
j2DOIHCcQ0sGVQG6oDd+nWxcsKsFJj2WcS7z+TVwsSuPWgrE71u9WPUkrYsRri53
H1GJih5HM423NaUFa8QdMx+eag62XMVPMz2hlpnQFRqkQSIS90heJR2yFQ09J6we
siHgzgr+nX6baSEVWNKQpcwt6E3qrgPf+sU9HphpSb9eHEF4gPBPZfr5Qz5Uq+KS
hSu8CdSR6mS1DVUnhL2lXRiwwbco89tusgjYyc7l9JIjKNNdnsjZmgWU9LvV51um
g0ND7WbZySfpL9mSxkqZ6Sibjq+9y6MoxYQsMTRCl7AJK/8cbUk/TAmxd879WJE8
eiwEiFIXPLsPGz9OGGCxfQ9WHpOXVbLAM8tCra3pWem+1smamqB3rpghFNhoXibK
+jmY/ojy2L3wJ3PAyioncdVmidzjb1671YHBV/vT6YOTWpV2Tptkbjh+XeyrOxED
UXSH5bU4Y89v2QrPB7a1SfXWcgxp6t4P7/yKpDT/OqlPjl6VX+w1yQLKdhWNn1wt
UDJRv7B/jscfRhuCtg8N2rglEwDR6Fe0NbehEXLpLhDt4WNtR9ZZOnbZ0bezcJOn
78/bos1UEZTgyJkHMJhICBbPONwla8oxvHr8/EFpbZNHeeer4GWhIiwmpIXeUhXC
Uu7H5CxkvhxatJZslNAWn6N3h+wPVapfVHot09keGvhTsQ58Zd2NB6NU7xE0clxa
zzHOXSxfy+L3IUOrDalE+EWhh4PNHT14IaMjjPHRvKDN71dDCpCzINX2424jzn15
V02R2aBibt+R21YGgVscvvOCJAF58O4bPAZFHRGoWuWKxOec6H+KsMikqZoYomPx
/G9DH+Y4Sn17e6gAlvlNqweN8E9BIvrRy5Wv/VqcLPbOagyYV6jf1ez1ej8AJP1U
Kc+y8bzph+E2bg9yY6dGl1F+7mxeYNR59QaPimZQTCPH+YGg3Lt3O2FmX8CaOrdu
EE+Lqn4NHtfxNAQH502fQT00ch/WGThLMtC5uhgsyOnUrEeBSIzg6RfydQsCS+jz
gjo//vAkC90YoDCFEoNJI8F+IJ/tszgZ/CmAaFEvyzKUaUbq07iqkrSmkrVzbhEN
4TctwCSZhL9VE6sk3wXyKUJPWqlxn43Oc8hOWilUE0C/3rTTiTLbPMgbX8XsxNEj
1cExYRDYT2C4gaARPBvJQOabb7CaRThf+DBcHuXtPsnoaMZN26xRt/94vq/dWa4I
k+HECLLCr3pK1IkMfZOepZ6IUbpHJ7LPGJjukZ5XbJgU7I3WTQjrXKUkAnwR2XnK
bTTBCZ+UrB0Nx9NxnTdJaxgl6S1pV3IK4aaHV4IYExP1oi+gLoCJdGZgFpfBk8Db
isWfm9uAN/Fr+sIMwkq+ojhMqF4kaH0rAbm/yGsbxw/DMC989t36cQvfMPH1CTZH
Kax5smLLcELE4mEklehyakLQzJzI9xz7OH1KUyjkdOBdU9O1KTgozmUfyVBMdHuJ
8lR8zi7HCEpPd2U2nAcR/Ic6BRvw5uX0jU+k9XwZQYAO/xRkW70TDeLUp9oXRdR9
8eycNIUC0HpX6lou+scFi83JKfZUUK2aWuxvB2qX2y0G8/c7TQyrgSr2oOgCo1SB
HxFXq24BoZQzdb7sV50yiNfSvZDi3++5zKCDfXHmuC3abQjuN1Cs9/9P1Rg2/tCE
l7TNqwvVvLETynYjZWc0VKtMIeWshZynPVmMqv8NQVkS34UJfbNP9gwMZQoJwA60
NPpSoKRaDeFIeyLy6kHFozSONEB+AvrcFssbRpuvIFfOvEssJN2ThsUJxVB16gHz
VcTYV9kpuNzGI7LO/2EIXY/6TeBkUb7svg+euB0dU5KL1O7waPs+vp4T+9PBaBD4
Aw7ET6eEa5xAwFbuRwvfR+MAV3iQQ0h770JFAsOWkolrUAvSnqqLhZN1tSrEFiDf
jA38avDbsrWIiw0rsQuotRY2LtbGSMQXpKQqSVC9j0XEF75yJ+tB+tQEU++HQKWw
pko3lvF0wl2z8+BsfAbCvMcMdn3K+YiXj6BHHQo3fwsw0zCnEY41XGnByC+rSB7I
HFS901n+T5pHMiR7LsZQPHYjT+zN+53+RqTJ3iCSOjWO8s20WGxvHTUFICqbfnWC
4pJHyJTklCM4RoF5TnSrDXMO2im79G5/a11a96IYRoMCDAhEYt2ENY5XG3PX2DSl
DHQdtEpYUalh+20MkTeUWBim6Brd/UmuwynJVrb48EFmpCQZIGiYzosYNBckdgBD
bs8/gsWjwd6KnDR50ICHA7n0XVU+ewk+TVbtQU+2OOqWgDNQX3lcuAjo5aGBA+YK
DjftCx56zFjAdm+Dr0bUp8ShNOZgg/t2rDojWJ2CI2aMuK5RSS7oejlRwjmTMU6e
G/FT2aBL0RT1flc1ciBmHaSEoAVnKb086D9qTOrOoVZuZaQzXn8WkGpILENElDwO
MkE42Hx12c+sqoBE6+TN6fnct5YOTDOl4dDu7tayrsMmkbe1nfkJpAKiGPU7QIt5
7zLa/kzIX1f0gWFdvOeIaydgz6n/HDpQetrzW29XSJ3GHMzhba+bNBbhIItYy5wu
DL5BIdY3lc+nxPhsIX4qXbsSPXgkRsEv/CB9lqbSEH464KHTOaIls7wkk7bSGCLy
OcYf893l/3+rhlieO4IgfZzcpN0/a530bJNN76sZsnOvfJwZlSboxoENN9k+1qFL
LbsZsAThn9D7z81GCYKWyCUEnYB142x3YCgQ87Hw02w/of/C55m67S0nMcnIOmUR
E1gKfrcW5gPhNLaovYaslIIFKCrVkUjQCIgfBBzE8iUa6kOb5/N4t36mz6yelpq7
aqtqWexvr4DkzWRpJS28wIDU0hTLqgd/gZyF5UQENk4HPhbrKNeRVrg3DVEitcJO
MoIWwz31iywrD+y5ErZza9WBNIFr8VybadVHjBHu5WciKYn+KoI2GXw/i64aFLtr
dtzESHzTbtktxgzIvNw3um9WvaLd0IjRc28mFOE6RwkmYx8QUKeZPSw6K3XyhvcJ
1thqOrV3iKcU7ys7Z54Oyakz/aDLU/CMwLAJ6t4pTpAUwcmreIxvPax8j6ZEzeo9
Qnb7TiRnoHFJmIrYlBuCRNsyENKgXNgbqqR2Sg12uSc85WtkSmFEz8jEfcqsrUio
WkBI91K9hdadZhGQWfEgb/vaSDlCx6CAo88Fw62gYAAH/ina086f9GHXFNHIcNmI
bPkuxXtDRZovgshDotF2zl6ka+mhBTMkqt+JR08qnUp1OZeA1/9ZMx5qVSWlC3/t
DAjxQ7dfiHH2o6jTfG2SXQi5rasiJiQM9vFenw98RI7Y+rbhVUmk7MHiLbIIHBLW
NQtL9RI74SJmpKLkXvqvGrhji9mYr7ZoolfpTDoV6v0eUUkbjpbSAXvZiIIcSott
hlrh7jhLjFqtRjF5xVKmuX5f0XWan5gbxZ6CVRAQETjHRoPNhthyXnNuhFHZpdbX
hqveHgPe4HE8APZVHMsJ/ifFlzyQw+5QDU28iZVUjnFfcvwkPqkNTaLA2VmEdBlC
GyymJH12HG/PheBS9FmrurC00u13qeGo+m5i8P3y5ORW0pAbjdr6nfe8iBhbk9iX
1w1fIo9dkUEP5jDuWJavne0l4X+o/DSlUFFNAB6YBRgPbjl0XOGIwlx7H7TZ4vav
W+2HFGzjyLHAmkLJWNB9JHDskRsNf33IGuBdSF6+OLvnr8FLwmK4uJ9BAnuDFfOI
ga6abz1ZJH+0wJqTn5gyPUY2IS9DdWNLj/qwhg+t0ptzFOqJCqSUZrogk9LptZpI
Dwld+KSaS6k4chr/dItZ8mRH9I8TvCewLMsMruGgo1eJ2R1SszRB+Sri0Ii+rmQZ
ZgauZYRqZoYv7iEKi5rgmi67N1KGoYDg5nOxEAO49V8uGdcLa6zGg5bMhkW1MmwM
W8jD2XEqXYnrmt5k1VRi37np7T5ljn8p2Mbvub6VJsZ7DzVQXQjBz5a6zAaW2oMg
UmwIQeyDnW/CS8+BAro+/w87+8wCaMB3ojvP7LFOpQ6/l6TXdhDvA4y2AfWx/mMq
3ST8tUEWXds+7WCyMc69CdofprfPNgN2czRLWv8Ulj6d/xG5dbVzkBGRpi05696b
dpvEMDDxqi2jcnIRsUIdSfzJ02wNGfSnL1/G/4dRaQSqoLXC2iqo7q3rwf9dwLM5
BC9ZlD1bjUwbK49DhM6zcRKNOKAxR0wb40Q8XTmL5dnVphACT2WuRZKqpfR9w4Ep
454MN/6i9vTWlIvv9/zUbe3fPDSXS6nKeUdwV4GSvZmPQcWYkeO2HrGRUqsK3GYm
nrbMysTjlwkhRhz6N59Y4wEVKVPvN1F6JWHLcZhDUxaaOUemkC48yhxuK0XOtDvT
3Vvozofy6iNxyaI5SWvYCxxaC1sfi6GhlJKIWfZPTfAp3YPRGTUWYiN1rzBqjjbo
H/k2T5KP+meytf1tI/y+0pAzxIJKimaPbmiuhyfDH2l4zibPbIeKgpqim8xendsd
/f3yuybeVClyBeB6JhvkLXv4Bs4kW1rPZZwwcA+6g3ztepv0kCUD4w6wBJh3zCTv
dyi6CopstzrZdeys0fjaD+FjQWqIX6WxW9EDF13uDcTpW6VA8e5NYOHZ6XbmloyP
nyjtALIz+DLnVp/oNtZTbnXJ6yS+8hsvzNAlO6UhLa8B9K7QZCLF38MwwSqyVD8V
sMGJMxPMtSBaqZbpDJxsbclwa5ZL00lySpVOdp8NXLmJiaKjX6Af8GCNLuwIb2Bg
mmAUbAKdAJcQTYTpG51KRJ2DsZd7t9Lmo8jxfN91mTJMfZrqSQUWZYC2id/aRcQk
Jreo7X3o8F5SW8WlbJoFKzfjhsM3tc4GTtg8eFP+8rjzG2Nw6+udUF1xF2q9Zz0l
k688dE5NBGS97wQg9zUgsQqVP8DmykN8bUauh2xSvda2WeMFUUUrs4wzASJfLxuX
8sdd5M7mGInpDL5/z1DbdmTBGlaq2eahiKECfGPxZT3fBxPK+kt4hSmDwJgdby67
qy2wsrqh+NeifIJshtx3Kthbmot4oV9mFgrb7oT3EiaN6Y6JC9KUVqCJcklOGNw6
m0prbrXfJj9bAZvXrzFc1w2RK5dgKDOd3zbIND1kzPEXGiQbMavccXxzr3XJkHxH
oLgQa483AT4mrLbY6jocQUO+Ct8rSN3XtJ3pYa+oGggJAoM1oDRMqbUpL/wdO5W3
hlxcplCcPVsJD4id6ycKmWftVxTdZanA5b+gJ7nmrTMxGvAQU/6P9VA5dLWjhYYJ
+O0Sgh5VanT2afdermVUoVLgk5GZDGxoMh4iob32XPLVN6rgONaZHd8VHFdvEjiJ
x41cdbSYzxJIeePJafL8Cs2aqpvlEq/D3aGioheg4nUahIOvSdA7iBZQt3InhHIU
ICl0L/bZ+Pywp+GleC718oeM54BkatKq2gZ/mtBgtyip8nvZeOvuY4giRMCbT3eY
NMAwL072tLiSuklG3llf/SrEpToHsHkF/MCg4lkdewXRqnEjVTczy9slQLbNTLwl
HKBm44lc8qmMUdBYJJMydnswWTNwNfPNv3YHgMMoC0LMv5V7t9IR52eJh9o9+iLg
D1rp5rWs4w3Y/Tby6e6SyBK/CMUFp45PAde5m4/AaxK5gJaV7UE/QG2DTpK17bK9
vdNiUdjrI5YVJI9u2IuMRcmmpg1t/2gZ3ov1G6ip8viRcwQynmkT2aAwnhpbhxXl
9Jd8CqRkkosW1gSzmM4aAXmKkgo8bAOSn7PqICVOCukRDd1NDHTS1Zl4x01Z9OjY
H7gL+lJGoLLzIxZfCeImutw6Q2FaWlusQmDG4RwdYLd6lob2PQfLMdy0BicXtA92
hEy5ju2Ap9xILx12/y1JP/ATOhhTRZLRHTrdOHrern+PX8bXGp8KkKenxUqNiMk/
cpBBOnkH3UK2nf3sTJgkCmbqrKcmj2r2Uokn2AQ7IJbASCn2PiCsodNBghZRdVEC
QRWYbdMgsvzCpXYxoz5IRC2b0wGlmGiDRSosD0UPUD59nzZo9453D3RzfA/5ZR6h
pJKZXGpsREIATl/l8U1waKmH1kxfKFT9HZkscyDQaCPbffAiXoGM3GbGoueCvpf7
aycDsS4AEKqpnUYDXXFufYnNuf98Dse5pqiATyWCvDUbvdD6i+MvZCXQXzUbaGV7
tazv5xt1H1ygjq0Ej5Zhyz4lfTxqamCKJPHprWLD66hQM7OeHhtEDmL+7baeqhoi
w4BpN/vw0NwPAcrDr0ZoHivFOpx4/tDmjqMCjJe324NqIb+52z6tU/C6mEH1HbuS
EyDCLpAWE0Saf6glsEip7uAC73b8zyQsfa42kioNNlImm1O9DTcSRhTZTWOk3rrB
Rb3oJP70iJ8qWm2xJTezB0/jgrBMCaqH/1aHj0f6hvM+aqOs7EScqa9KeeBjIEnu
UXh3CXRRkj/Duhw948OAWrcykK+v7/WftkKACvPcC1yjUkAjznSWUXpty6rUVKDB
xiVe6Zo8xcFNr95jAb6ChbuJyzZSZq5xHMroVJsbUxCUyhtVcc+ZCnwvywFSJ7Xo
ZGZby3BayeEsUosKlxAmPbOMJPuO4uEOZVL1/WfXAWX5gS8rTxgauuV6mULvLbzU
S3YdUvCQ00KXS6N42oGkAqK7s37uipddlxdrP5W0cvekIuzUXgltNBInAWImn0sB
FaE28wdaoKqW1qtPGKQZzPhjYy+56gNWhXwQx37wQ7+RtCmVlRqFNYNkpIfJqmLn
4uLhdEP/wKZonQuftUmujGA9qCJ4GhhNXIJNJ1S1/HtS/kjfKroeIpFIfx+tS6yN
71Qih5c8d7crZsUk6Bs1QcSggMQUkGYq5VKM55tvt9AZKiYoIw56LqQ7Hq+4D6f1
Q3LJi+Rjq245i3Wurm7L/6J++DsZhyI0fstfg/JzUa5nAwOTypmB23y1uWynA4EB
uh4hTs9TGdFVkou1HmW6Z3vKgtUarXt4w9ujWbxdqqqQ32IaAKXaAcMPicERyBGY
9GzRbbAFCaVWV6VGOz5xmszIjO4HvN0ZPTA39AgiA7wbLqBMwWrwJrR6A6r60LQ2
wrK4J/NQoWQvesb3BMn+MDKFF52ztnFmw7ohl8pYqTV2D8RqYGCsa1aGQKxSX0hb
Dwpv2LYEu1WDIz+GqAQ+nqA6/3ZwxCn/9sxT4MTvRjFS4VTIk3UQrts7mUlnhNdt
bLbaFWkrrIQlWIUHS/oJyxWaCZkvjju93r+qTVXT/agbbDfxqtPO0Jk6SXlo1Usi
BqOVHOz1am+5s38WD4cFgwn1SwGgN7xJtkvm9Tc/vvxyUUL1voLlfKneo6htlPGO
u64wcyXPfW//svv81qA4cdoBi1ig2iDmRF+yDjAiRpXSmGA/PT7jNWvBInzdA2r5
McjfXtGylo5EcfbLMxqxehUgNSnJCwjSQ9be0mozgaDsnQjxnGPZwLTQ0PDOxGWb
zXizpiHj05FBYqrpoJDaSVaO881/9oDIwMDpvbMDieMCp9K0ZP4XGUEUWZLBKcQP
1b8fyvcsAiJrseXRaRX9Digc1mRpt14POZvBtFUfQ3VsO4R4ptv4+ObxVLtw8H86
jSZ7alPQ+aal2l7JwA32I8rupxNEiqe5hGBxvV1f2VhXls/74cJLjBAbPj5DgRxv
VV4ko2tb3+wQz2+nL1VlOFA8y+pd8eGBxUrFA4ozjp2mNcyyDo+SEeRWT9PCiqu5
+IyV3JwX/lmTboeoELHPRptaku1AgRzEi+fKlARe8oIa5eefILjLQi1H6woquOkt
WeOBevl6Mp4sMdQ74wSr+HpQaN98Ud/tBp38A5vxxrNHGku73xTYtXO94Y/9ZyxK
G1hnD+B4rAcpd6TjoFp/S6ZyTYxZJUDCytc4B95gfuwS3qLlxU4rq9IIjksOu+1+
mlSelqGmPwz4lgugqpVtnNvRefKvq/bRS4C3RQpCxKfFNkOh3tetDyTK6WLl8xUu
4CgQMRvD5sXB620C3G96kxZsraG4evRD1DOLLfBafQPnabIhniY08V9xv193MBpx
DcsYuSE9WN9o5fJdxWu4Bkmp5uTfBFjasKYMWpFGEbvU8IdAyWNqz37gm0Jyr0q+
8A1PIV6Ip4DYeLqn9zPciHG33G2pbNKpHP6Rr3kpsnKUGi9pG+yXxeQWB9V+R6uN
k0wzRrX3dtLOC+UdVhzhYYyKLVGjoJJK2qkxWWoWA0g69mK7F0KK/T+0wqnfhanG
u5ggyWbA7fxp4SWXaF5JhSmQ+Y8NhYqg62wyC3t3m9WnyP0YcuY2ehiwltFINh1j
P9CjmcU3E+C2ze77026gW86GvjMpthoaajTrBtanuzZVIFytAN0Ryjjh3nRts+sT
jmI6KMa5iS4f/knfwNMM1cNQ7hlyazP6/f8Eu3WCgGK35AcsC1EEP3EpwD/XiaGH
OS5ggC6GR2Rq8OJSUJ+EDGfaP7ZvroNz057hCk/8RwkwlFCzsZIXyvdlva5ldX/6
cfCg6Vd4kV3bv2BIipj4OGMdF0+ORIae6267r6h7NvY1PBG3J0wEE9I22hqLNiFK
v8r4kof4Y+1YvKvGrmYsV+sBH7mX9HrP6Sy9ZT81Yor40eqaUZTQM7pHvJGdZopM
mvHVJ5I2kYnZGV/XUfML1WmwGUaYeN3eoj1o57MqYUdEiy9A8iXe5Lt3bzBochdM
ZP0qlbsiGRkRCgBqeT5NOtnE8N42+SMRee4ZomdmyOcvCPj4Bv40aQbEuFADGiH3
`protect END_PROTECTED
