`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fs9+16iz+tLzwXF1n48J7oZrHa09CsNjZ7UfV4cUe30as66cc1MG00dHbzeATgAB
RxiJIh6f6T3yZhPrCmINrtpIbb7gTgst8T1tMvJukSuDFv5j6Vi24cQgee5mVQva
fQo5Qam35MpZQ54BqFtwIpVkTseg+Wp5eRsOQUZBUxoBolm0/zQ+7ehqki5EvSNy
eltnfnq87nBIrCcuKscbA4ZBdNnh3aHTSIoiq4ot61OcmUNxT6evOtebJSqAoPWF
Xllbtudc/kieYOPBdKKvYb6ZbMUhl47cY20Y8/y4yMrCoq5yJYZT6mrskpxbB8Jx
kI9Wi1C3JsNvwqWdP9W1llFyyv7JEk1MXUfEglHZ3mQCCVLjGGbBn0yLngJBFAJ6
ljfQf+wyQFIWZqezK7OzKfG6z2yIGoQb1Q7a4wx+r+I9SbNV9uip2cOyQPEwOFu7
nXMiDxxRsnmn06lkDKxincpBORS4bHV8FChnG5jlukj1O10e2WmX5ixNJG/C/ryx
hlZQCgKK8YRQ8elzcxFSvw41eswcSa7cCAIUqRevITnafq50deAg8m4UIAN82sH5
`protect END_PROTECTED
