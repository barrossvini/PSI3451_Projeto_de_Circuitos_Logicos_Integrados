`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fL+2J6GFbrj1cNInKEWg2YMWoLpl+2t6CqmIfOxuukuB0CaNKCzMslK5HqCymsm6
5ZAih8n6dRd6u7WpHWq+zN65wMqcuPtS4yQ9Cr2f1pJKQNNjIKLvBkR/TQ4oRT+W
X35VDbwaQmNa44I1I2ZylrJqxYqi1d0XUcKkRhWQWraRCkH3BGai5FdAIORIOR9o
5ARxEtO+T/aPrSFgPH/RvxfyPK9u7j7BqghUCNarICgKEw3YyWSW8ewoly6g9mBV
a+v8Uk/MMjzY4+xlNG6Gzu0rBKqjvcqwaJT7TuG8D4rkZ8GXeJffSqfmNukAJEvj
fAYxGhv5yXaNu1HnYdF8ESrYEulHyYr0HbHVLkVCyfyA+0cUeCslu03E/2q/YIKu
4N7moCnJslAXrAVG195+mKU8aCL9RdBtjXGxVGf06iksFqRZN6pRfwqpQlMDpOrI
VDP5svrLAvevUAeKu6bDduACXjgwUrvJAW1GADzQxQBakjgnTEbpywOh0Z++vvGq
kLb9/jvuMZhqjZTnv5gco/NijlcuqWWNGlb+6URruHcy4EfAl+Dy1uWGgBstzgQO
SOmq5lYG7TiQ3FFdfgZpY39mUD7uEZNwLkS2RGTRVavyKw8kc74sE48FJHzpRZgc
pWAbOiCFqadw+MBtaT6ZyDcP58zdFha375czIjbvfOIjXtep7s7JSlmLSMNYFZb5
fPwISlYjEy/KBSN6fn3rjM0qnhbPssYwcacTJlV8ajvC8QdW9loLJKqz3AweLRnI
RhVXnIVwQcl1iH+yDtO1L9qDE8sSIlhcEfTp7k2R7lxCCntPwNbkbsgGrg7pCq92
8UZ5aL+foJ4NwNEMrmMiskGWvpbq9CdQVLI55mSvWV/Oynr3LVE46jPPPMLihn8f
Ub+xhTn65OTw1mrbCaMipX7ZvxixQa/OcGRyPNLS0/4zoQolax9WRQztB5EKK7YR
/YRafe900jRofLO7nv1eejFn4YVNDnZv1gOEpe3zFU105W9O8nsVRzEPkA7dyveh
q8/0nZoqibMek6qoEe0VXAcJXKQbetVRSsb2NhohKrPd/zLC1WNz0iBkj12+9uvQ
QkqYi/4a5S0PmayZKRlU+ML7xNmxwPwCzX+ksQJGxlIcxfN5siUH1n6M85kdIv99
LyH8iH2yyhUV7tDOLbmssljaZJkCKAPGPkkl20skU1sEOV32oN78BY0xg8DFZM6o
IqSsn+QgsBDH+11/8E3vYdfXpfzljzeS2s+hGqLhy+uQSQNh+SA8QDx5L02rNF3L
`protect END_PROTECTED
