`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IWVtsRUyUSYi8PWpPuxpijaREztubn5h4HVCAu9KJAuDc1sfIVWP6S810nLwBV2a
J7w7mAR/KlLgFt3LJrGMdYbFwB+1kBI11rMxdUa+teKjfcMPKhcbZZjX0S7kj2r0
umaryKzrWJ7ayGeMdrUTYpAyFsBJ/5J6LQGCPgiIuMpsaLMnEsFLzdRCd/UB5zXP
PJAp4ZkYwmffNRHvVGyseW7c9jAp/7hCDWYRienYgSb0BQoNpdac082L4x31Y/bO
McVAn0IGzn+M4eKkBkAZQRWi5f8jsAX/e3sou5RxGN/BInhlXVdnY0iIP9sEArP8
pPEd95V3UhFJZsXfdXHyY+5DACNYwIaLoKsXQMbc5RSSTE68wUaV4IAXgVdNUyou
anEkqaNcW6hze/j3Y3yojqBOXDPEEkVjTjlRJrOAr72rMWsgv3m2hhhaX3dZFq7K
0BrdfMexlv+4YNHwR3OhH9t74hE9Bugp2pZTSGbUMUBMjVWyWMPbJvNX2QdkRIoH
sdRzU2/kEqiQwssK76orNtY5zKmKTkNJzamfpGeOF93V4aYGMd8mo0tNH2zeo+Iu
aQaFM/YMHSa8sWvd3xjeCiRIzSDfngIJj7r1fG60gwEw+2A9Gqq5pRhwfkVelXk3
g7nyOGwmuKn3xhObKeDdbxCy4pYrQPRSgOme1ImL5KW1GVazwa7d/GtN3/UCngyu
Bbw164kSmFpPL3rHkdHKTQdoys5gizOaHvksrXWp6Fm9gWcTpqOb5itAgzlMiQ+K
QF4qbuYiKb5+d/vTZV0Z6Uux8xY/f0fS4JhKvSAdeMv8R6L9gMBd41IYJvPLMJGt
Coi8hMO0ZXGfBPki/i1X0FBsSQzXPbSAQXlaQoUZrRrgCCWOrqIMX5u4gFxbkCK7
vQxjYmhZjXLwrFhK9VMaPqez80iKRtIT8UXI0BVghW2XywOuHFYvKdg8aSzqPCoi
yUX267MqTksaB1+Ra84vDtQI0GCCYPoSQLHs6HxjKZKkCRWNb+eZsgnriq1N5pvn
3G2jNqoVON6eNB7e65B/sCByNSck/nZqpNZv9x9CCIcbtM8QkRrkk0irwC9ChPx9
qJf+ByBM2RJEefi6+YCeZVatQG1InK7vuFmT824NTBkMeFJwXKHgMPO/dFO2bpu5
UyfQU6BS42ZhaJ1zs/IwxUkG7UgIkmQ6urZXS1SU/Gye9ZP53eDqmNu/O11Fq10o
ACCHDlsQvdbCTmuwG9K4mr8/T4kFGxzyay7tHVJyPe/oCh2jM1m/XVCLgJZdW8Ia
f6PAzlo16tnH0uLC137lU69+8jK6ZWfVuksu5TlVM24yMWmNI0QDMGcBf2VdfMKd
eYY1Gm9n/dqZ1aYFqB1t1gE+2FTfkAK+l0EhLrhdXFKvJGG2KRLsB8bTY2PZdkCj
XZOZz5OpI8lfi50HLFnneaXgnD6SVM8K9u8e2ATTT7ao1hsbqSfZ99VysVfSEIeb
7AeWz60kG5+xnNUkXtBLaWNypiEldA2haZXfGxwHhfyz9SWg9LT/FTN6BTlZwJan
ZfzKHSZAirmvq6ssSUqj43CyTmAInbvIg2BRNp3ysX0JCCGh3O5nD0gQkoDk7jmg
NPsqB8Mjz61xyVVOZ4HAiSEp8VBxLOeyXky1pPUWMl0tmbOHu6AKJNBqddhlRjpT
BcBRqGuJFpUf8O0g2EHFWbGwZlSjO4QT/9sDeTjLpY+TjsK9YgZ73QSytY3stl+m
lCPS/SsDvlLR0NnzdlmtftJ+uKS/dV/Bql/iRdKGmOCo0o0rrMyvHBaqwjtMxvU8
BA3Iq/0KN6PMfAH2hwFT7iyVvlZWmeKObkygOccJfKZ+BRskni8KW9UllazlP9A0
zlTedL6+K/E2PSnCfJmM77/IR9iGQFfjqrOod9xYQYzMU7GAwefGZK+CMbUhJDLk
`protect END_PROTECTED
