`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WDIXyNzgdEJqZV5gH6/7YNUF93rkI2tY1rZADjq3ge1u/4IDT81EEdQcKAd4ttjO
nV6GPZPUueIH2HRBdzwmn2fiwm7zM5ca47o0AzSnTr/9xgVGf8s+ZxMVYueRtlyj
tb4hGPzn9P5BRDMLR5yw9E4XHkEp44cjoXhyc4dnnMvpe193D+oeBWcqfnV3pgEW
f1C0Eo6jDXZnWx28SJBMbp49lm1Fyftjb/luLPsdXjOfDUgX/eTLmzi62WzzbM29
Q4W4/ubvuqk/gCAOxof7ZG3DT2L5FiMtJfDBsR3Q5d8PiY0AuUHFVWcEzqU3883V
IN/VhB5xjMtj5oI5iHtTkRyNj3CpIgH2Yo08TZW5Q2KGqAUmydJElFcc1MYm/rsB
0Z6ePXmkh5wSi3Inc4KFlrCscV/6zaBK+IPBfx+ZslU=
`protect END_PROTECTED
