`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vjYFTuIoXLNtZ65WU4iaOswgl4B/lP/ugJ3jPvVKat0X3di8Lt69u5jyo0inXB0v
N2/zIVo3vEv3rTtEWyJQ7oLQ8kauVJnaYaGahAuQWAW7G6nEyFFS9BlMObM5zeYg
ijXvW5/kBJAO2KzLDaA7Y8l6hngWd6Hd6z31WYAA6aDF8gK1vGo+i9DEWRoUz78D
tbso4Xv42sUl50IM4eYJMsiY3dHNXymWtA4M8hDkzX96FKgJrh0rdG+OlnZA1FqT
RDGPYv8rltHF1wAn8HeXPJ5LC5m3yHwAXc4jSstPcagdTyWjgtGfTLgVazR9N2nk
5iWvzmQuvCf5nBY7PKvCfGj82XxDOCmYnFLGCOMJQa5VteTSaEdiakWIj5Ps/7OY
47xxuIWtvEJDk9QosGhxRNTkHv29Ca0G9w2EoCbuuwGQPBBmu1e8P/JF0EfeOWn7
xJN91FOwrrrpcvy17WrZtOcyf8Qo2Z+SGQG4cxBQ0BTA7lNtm7rw8ONpzEGJh3T7
vSzAQsdV9DF0ydHJC7l4lB7DgJsXCgkwOH1fz7knGnKZlRuYerveAWJQzt313HPV
uoLX2+SqhF6usNBsN8trtfgep3kfPC60O1oSq9t5K9SosCyulYUOIgf44c/nRr03
oqU/epJ4wy/s4A3nLBX/WxweWl8wtGNK+ChBR5Wn7NDH2jN66X+dlTpa9AgvGtD/
lRB6d45vA4Pe1Xeqbw5Q5MKlXAQ97gD8kPl0tv5Kc5enHwm6V1UdRCJSbIMnXVsi
TiNzBz7BobYHjHs3fxryLn9dXKsjy8zjO6VKSvw1jTLdcQq/hieoJ4sVcXB6kU/i
tmuBB+zjp/7U9gVQT8xbfcQF9fefv/+k7AWAFDcscvUlUWIAaFBYJG/l1stkHzYI
cgzcPqlGSThVQwcm62s0MiBUjKFGGTivNq2zEuejnUdtM5Dn6rtTk70K4mlxWfP0
ou8FHOKngbQvehcQwI6LO1ROY4fGBF8Zc8KZ7/S+HCWh9NoYN+QTTofIC8Qtd/8h
xdjFHm0BV2L6Wduva8X9DL3nFJ5WkRP9+YlOspdCckxOqeykBvr2w/Vv+8VkGHNc
KDL+S0vfgDPgcOOd60im7/781PWeVC73RCFDW938hBahL9L29F/H/Zw0Rk7dMugz
KRb7fXPfOFSyUJfOaEEIqVvGHdLBzEjDekOd282GIW8sLcLwqi170LAgbcBa9XQe
gLNNZII/BM/pNQGZEM1y1DjfSEA9PogUR6kDVWyBPZTEbDeweNK7CHiEbshoQT8d
tKtyjhtz09pZLG4feskPle2tXvpTDOQDpBLP+IPZWfKJAmxAA/xgvxJKTxTToPii
NNMQtyYq4vufSfmjAdPO9Frp82MdoLgyqUIEjQ2kGbd9uF0wyDtYjI8e+MK5Chu2
UHi+WejFn8fRTT4fmvRmgPHuweHx0B8SVT8fXEFUPBC+H01RNyZ7bhK3t2vAKZGT
pXyyrb+orRsCf/PGzWda8czc2S3/c8uuxlpBUjs6Qb9/i0ovESKEGnkWpaKDFKEX
kc2p+RZgoVSzQ/I5tjRHHfyLvDHSHNqwqGoXXa5Ot89r7B2UDeM9V4zEvJx1K5/N
pXi5OVvq8nGQ+XIeYWdebDOPafjTHqqkYBZ6XUZUbUXFQhk0SEKxYTEeDS1mtvpr
4r74auqN9ZLhb9ucd/zz1nDeE82uvLjF37VeWA27YtnriDWeL9Oj55od+YyErCGo
fKuLhbeWxe6puNGKmc3McXzpQpSf644QtAJIXCiVew63/wIb5Ce2R42A62RfPtRl
JVCV6vs34xVDO7I9KVzEZDiHjBgvGgQ6gdQoNmI69nP4Sg/5P4G/6b3vXwU3onkM
Q0QEgN/skKKZu7/1vP8VyjDH/wscDmkyyTppiDPvBr/4y6h97YshMZmqH9LJ7JFM
kvfSyvLrbpRQw3jNCN9WltudkF0tbAUO93eNIUDGDFED8F9FZj6lSeIYhVk29cO0
uk+FGUopVKPJ9l0wR2QLLHflsASXZ50XWdVr7++cPn5XyW74Uh9j1rVf2ECjq4zS
069qQhlcGrwMqpTPL7cQ33x7yla8hunRNLIKOSY2nK7LZMep8Q2UT/Bvzi5Iszpg
RV+pqRKGuNCGaa0u2taKHqbQDBzS1gMUHNVPuLs6xzd//kcJBTovQeqF39RAMAMX
Jud9INPL48BIHg09iIP3knB6fg6oLML8dznkecgm2RA6X9Y6BIhao3z5ZC7FA2nH
cXBYywX//YbCzKpCv7tqJ8VqMsJCuF+ktzlcJmDmW4ax2Ys3UY7rO0QhG2oDJoZC
pjtOpwFWSjdBKF735CG/IdyC62+cmUp1ZJBiaXSn+Uffthhg7ftmh4hDdbbZDAGY
FOs4+2ssqaRazNykAdgZrQJA9NaML9PxXBtSuPHGuYHRQtLkacZx1G83pk857X/Q
+UgklRNHhyHCicNp24PiyrlUn2eeptLo9IxehX8NYS3jQYAgRYNqhZkU3OnVdWs2
/BEe6Ba+DWzCp5FjfrWIhLT4XmNOYa3iZ/HVArjMxIha9guD+Ihet56lMvuznrIV
/04juRXjjHtyRpmF9UJNX/g7Tws0cBjP3v/FQm4U6hyh3SeGGUIGMgNpSz6RTmbb
lPdJjStwsGlnzyFjYq/eVLX/h9+349+VtkJuvAL2ZML2hD5malbmKFvnp5LNwHg2
brclsJLsCUW9c2JKtarHLH1YVoyEBPPY5BaY0XGT+jgHvCapLJQpehELvxiNKKrv
kWoZkrAsCu6GNOGGnlzLh7Pd7A1gw7Ip7ifVp1znd2LWCTnvuyIUwtjFEOZp2Ohj
P3XXM2QMKNnu0bn/XuzdxNgp9rrOgADHdae/RjIbOJ+EboxRsQTHvaj4002nyb6a
LEPRgrX+0mTWc7vvwgpggNFr1BuetP3ntdpXZT+iC//yZz66V8rsMl4jf+UNsi5g
ulDrzYShrv5dtyP7ecy6UxJ1HUyOoosJY/+iDIWy/XCxtvZ3Y1hsHHUamgA+ugEx
UI7kz3o5CxHUs4CkrGbFVSbIdhFhisn6Xt2F+UQvUlVebcTEbbpdsA9dgtRKAT0u
7zLbJCxfHhcLyBV/AMO1ynpOKFhDuHAvQ06fUyep+9Je2ZuiatQDfE8SiULCwc9/
TVoNeso76we48l3VkyjjHUncykZDbGdBvYqVQs/kcRFcwgW8hbtZM0+dLauYpbLb
bLra0CG7ld2uvIgXyysZigb0UM1D36Ujl0VaJ0G35tCt/3YdvSsN2+prsZADxX58
F4kKXLjcQ+uypadWxoFYObsmrm52sfaDt0mo9RXRr0F49JPIaLmN7HdxVCbrQrQV
1jKuAKLQEsRPKtC30FPp6qex9XWwyfzdNv9Bv9DiKw8vDhegKkLi+L+tBdQIbl7O
+tI2YMlCQbc2OHkaqlxNRnuQ4k/s4O+3kh2WYSq3oMlvKO99neh3xkbWvY0WYWgJ
tUAngEo/aqRYGg68rPz5x3i2YN9o0vOAF90zPS5hdRbICTydjGXC9VI0/odK+ZCg
Xse/CDgDIacY4RN1Z1CygGrFnJsnLvRAIyUzaCs7qZn4BNJBfIbSZUTijcAgpIyS
ytFo2l1zmH2POpFO/O+p5Wf9AHIUZ3G0iRs3o1hXOQMNYmDiWwz/TNtYgtuQmHLF
Fe8ccTrLyzxT96T9SkjQHcopehNuXsJHv2iomZnIEpYzsiHJY79c5vcLPlILMG1z
RMqEKFiIoWi+ZrxSpsI9QDAzE3PlaMZ2B/xn4BHXsLKNbCb0+2AeCKGzluFu1Kra
hT3diRKsaKB0tqrdSbyXYLg2GQRY4CkFrjUGIMzt8Cxde+01sZ7IW9bJo4SaaS/L
FlQMs4PndlVZcaV41cItRZjm9FAcqNnR/XTEHfKj3jNzagUxVjgvGFJjE09tFhKJ
V0X5f5SfZDqvBxlR9ZTuMxvZP7LEEs2pmk0Qd7pEINYGYycWsjSBc8cMwoR7+4tP
QLyug/5+TkseJ2565YWpsiOajrw2VexSOPWtPI+Eh/hrupeOYpkZna1z8Ljx2S3x
qLq8iu5FOuBwcpi5jBfXjrQL3w3A5EVMbYyyDlhcdyn8ZqvuPoASHigxP7WpTyFX
lQp7nCFnoP/0mIowPxHnoQBpE4YUHmvaZO880WYBWnZTSwTAbCsjmGFcscx+uaQE
wma1A56AjayFXbkqRyWNZzDYPZQLb2Gv9qrA35XyZIwdGEC3DN/4AfDV3FZ6+vml
GDFaIJBat76VeA35ivsE5NrojmBJQu/PBf26dQ2iwslW4s+9fjp47o5QY5JoCRvh
iqdVYnSQa62xKksEYQ5PujHgXg+oYOZHCfy8OiJ2PRWu42CUGPV5Cmql/5aA1FZ9
xCmv3tHlh1aR5oLHUg/fjCdUE3YzmfPGLe9kX88tg/1uSxk4VgBzFmWDeXK9uW0E
sXyEd22uQBPdKafQfsD6d12IA5fyM152KxNw+fVHs5kSE15SHbim6fWfc3S0RC55
BgZUole2ZYfnOSVSAyYFsqzf3x93d/Nuvd/pGJIT4QOJmKy3aeckdmqpC1HBQFx1
fVbxQPZMq0/KQna9GI2j8nn6OfRXZHS2ZNYkAbeoBzJmJ2J2ZgNY7lwgD9hE5oFT
oicGCF5NKAGgV/RQcgTC+yBTQqXi4BtheCGeDOKHSuUBplQL5TovdL7CRYlXIz9J
ttUyJsofaH/sAhbaYDIeLbYrMpi/JmkkE6IOhAz5+1DeUhL6LlisS67QA6AHv11t
pQFSmK6PuoxxtBJ+qCCsMBZmExdecbBSn/rTy6jhu4FmETGP+kWWAg8ErMXyqlOZ
VaLNzq6nwSwfd5Q72TFVU8Aa46ehIzew75MguqFtOboi4tjKwRSM/uuXjxdkupsL
C+bZbMdbTsbPSXJhrDd0hxXibRirfej272apfVuoeelwzEGweTbLaCBi3yPjLJFB
ieY4UybD+b5FUFn5OD9O/1oPoZ4btiWBohgPIcJKRHzF3CHpe0c1MaM9ealZzumG
CR3qy3AI/5Aqua4O+zzLxh+tCj/VNeL/BIl2A+mQPeBQpDlkJ/LEgK4oVcUGqvFE
uJpJn1AMMeSw7tBSQ4V2YFFBTTiIJIBzRiVuOt4yDubtDRk5PU1bDx2qjqtU2YRn
/JprY9O9+dWBseid1IeqNlrkMruCd2TZ8v14EbxwGYMce9AXXWAwE4lDoYZz5C/q
friBqskI/dx355sw0YvM1HcoaniPgF7vIpOsjFyU9bnncegw8r/7GudynZj0+lpj
5Kxw2rDaVynQgaeJY2P74mGo2XtPycQAqKhR9BWOS/Ixir3+GPFqvPTrQ5nXCHSd
`protect END_PROTECTED
