`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ToQB3TQ43En5TFTzN02Zf3UlmKA9G+wM6EGSBkMMR/ww7llEN2N6QvnE1ifro+xy
I1ReIHGKlqlpJg5WDjMoIpg5HM48dJXrQ4ZvE9HU8qn0/3We1NMv18Zt7elnDhlg
gh8WFYpWcCA5FpqgYQopnmavi1783k29xTS49D8tZTfAG2PRIpOHe03X4xQII08b
bh+PrMpJ2gRgUsOQfexiJanhrpgeLHQtKZpw+STQTaWx6MnM/nOtq75mmlnVF8r5
jVs9ODicOePSnXSdOojzOdENqbTQWRxVra85l+nmA0LH1nBWtdBmsaXqy59Nriz+
5Xisrpyw2tl3XRgwb24qV3kPhGcpAtNZzfcL5q0m+nsj276txhrPGKLSKiVi50NC
tjhC5FeJTA/iMAY/AqXaO+vE/g1pGoJ9vIwWAHj5I7YRtTOLPPFFOoE6igwHdDi4
ZHuMajA3YqerFdVpPNPETXZjRsQNvCCeQcQDiSegAWex1R3FIukx6j8MeF5RxDYF
/6doc5gfdCpzxvBJUpZ1K/NVmkhUFcEQ+bJLULqVK5mxhwsRYyjjV/MaDNKf/g+d
/7ijYfGyj/gGyLxQ+mRwFZaGPKO7FtmrhnSHsAt0VcaZDrqWHbavoqClKipfuWZ6
8OTrZMUR2NFPHf2yJ1xLDNFlsoPQ4m0vzsX1icWccfgE4TBE36i3Hl+5nxEo5B0m
I78SIf60KeGUovDNjkQIu1a5dNH9r1ihNbFRQOMq9Sr9ZosL76Yuttk01rPxq9ZF
EC7833bd+G3xZihc1UJqdOAc5jF0akWdQnzqWHjqC7/j292cXHzMVCwmXpBw7IVr
9yeaKTQg9xLA6ovItLdx/EXucXDF9/aBju0rhvwwUIM8AGq3VUoamwulYwyJ7M0H
6QjcKT4SY5iEmFDCuwoSYtVaITSWPjfXqMKjGbejdERIWMkt06E59uDVYMGpThnD
+yscI03e0qEVCvpbH1SeJbTI0yiMESaNk1OQAws/1Yhdm6w96V6J8YjUdRSB08bI
3kIrC/FmAuiJ+ZRJkoEoq+5EmPXnl6qIL1QGOmNh+geEBDztWrtAueHtuJt1PNod
7mvMZovLgqEeBGj72UCB9vHHut4AUN5Fke4/17j3sPjpsNQ1j2L/4Cww+T1vdFmF
TVZxeJ8fYs+93wfLAswe8378cPso0aC9bI7d/Hpx8LPfpVtRmcct0/ucBGWT9cE0
wTW3iD/fwDgFM2m5WFic8eKQPc8ocUv4xi4nHHNh/sIy6MwhnbNjZAYTeAfODpeK
EbUeoauoVdF64T3rmbAdM3YkS+U4JoJrit9AEIbvgne82ZeYrf2uNVoaxdul1O/T
G/cvBTppUhOXytJfjpvLa2LUlRfd2K5dbtGbz9MD316JGFNLccphcG6jZOvmyrtc
ybTftl5eEp8u/3KtUai3hd9rTI4XjgZvuVB8fUHpcUjd5/MUm02XJ1GOV6uwfl6I
wa0OcQVkO5P7p1CAB0k6gIMqr8ThWZuZna2jYWTpcq/X7c5NMgCWK8dqRzxuF+zx
YoEJOGDm6lMaO4kxw0HuVRjGSkB+uLYYjEB8gVecuD2Z3E3S/wdCixQnD6aR9Iox
9MUQJOFXiOHzZS5hh1/L8J3vqIwQjZbII8ex+AHOt8dWC6tIdBihM5LZ5kHLNvhi
Z/947klHVnyKwHC1DgPCxR2c+ZkKjnTQ71fBj9kQwFpW2SnF6sAhoBkdxTnGTCGw
oRipYGMiElLNgjE7DxGbJ0xZuppAEULQV47hOIVbzr6baI27GJyioCca9tJyRZrA
7rIb14SgEAMBwsOsF1XipVzBsvOp/995SiZex5jC2pdaMGMk8FwMc8yQPel6KJdZ
KGnVyW9k1DHJ96jNS2G3XqsT2kLN9Z4oQK3M126cDRrJcBJsLiYaya4YrQI0YJpL
UgBjaXpsaSyw/syFFBw95DaAv06P9NEwZWRGebc8zR9IHQl2iPNjbgW2iXH4cGJ4
P6yFO0ikdydDldwwJTXmVqpX3EeDmOiNgEsA3PKaBuKXm7N6avzB2U/DtCkmyafC
DxgyzM2H1zO6yctl3RV1DjCVk7AMBHSDN6ZB39dO5gYXaT3SWajJyKEzsbR5g7hX
rW0KuQ9Aj4VYu3PhqeomyOSxHqZzK4bwIWfEdDTP38yXm82BZ3r8i9Ty9lZqvZxt
cN1NQ3cd61TywAxxEufaS/r7nbWO+ZprQlN0DiogNufZoZrps6VNPmGsKNfhJBCa
7uZmNppE75fmia16Z41Yypd7j/oZ+rvop8eG+LyGyA0adE4JvNe7KiFoy3JOICKT
F0OzasYkLYkhHj5FDVJekAajPwHITQQdGS0MNxIT3z0lCznsicq5OHRPkYn+1M+i
/s+P4LtuXnkgteXFYsOwkA2ZzhtCeGXNYJTEAd8kIkdRu7uyYSZiBPMV4D5AgpX0
4QGDZS97vLYrSdF8HoBuWPMn6wJOQe6J8M7DzcQJDtZvH4F4AaQmwa6lYlPidb9Q
HRZy2NOwT7AmUeot+al39jaZbooDXkLDfmotJyM1u+ZfmKAPC9P/FEuUcm3bAE+g
eGsolx+dRzKJixLyhqsPtcCEftbNBrhbAnJmEsj/O4cVSUj3iRF6rj/5SluOph/C
4yI7smEhciG/8YBuxBuXu2BPxPwIy5OEui/lqHAUTI14JEXGISABkl20H816ij+f
WWmKubA0gV+utGOnSPjY6ikEgsB+p6DDvCVmrzJz+eqCRArweKrE2b+m8wnE9HkW
wKfsj1I6cExwZjE4KN5zSDRnGjL9MuhXvj/vmH8a92Ibv2BggpEsSCKioYSr9DXT
V/otmp2n/mpg8rzx9BqGl7IqWB4GMt+ZjJXFOxBlyclEVN42rYcgm1CCc17ZU//h
Wf/gq+ulrXq9Bhf7F+RDla/k0GZBcoxoJmhhXiolId8ilpvjx8DPXVIGuRhybaSr
juyeuTgNTPVyZ8/DeZmhLoYwUL80/+EmrD42iMXwUj2owKpYnSv/g5mlARl0CWW8
VecKmapqD7CaeMU/OwmAzaCWCmItD9OJSZtgFvd+8fnqulUp1STA6D6oen3ODEzb
ZfQa0FOG0TxZATlegCBZ+gHIc2FBeBCM5pXS0QxKfjTS67vcmxsjqyKgiv8XzSBM
63zHOn6zrhQGZQyTJaCtLL7YPR6kv6ak49SdqPLe3t0YpledrQ0IXLwR+r1iOJEj
Rz9z915HzY5ujAXuAJfIMmCgTV8oMrj06XUjvp5XIiqHwgHmxnif2sfbaGpirleq
oxp/vjk2b72f/goYhQsir4Fc3SbIFWZ1FYMzJC87Mv3QOk1Ua3TpGdwwO/65WUZ+
pvt3SBJxM1dAgJzc1u4HvzSTIzYqYQg3or350KOGIOG2eksq5sHmJzvXyaxYtxfw
RZXbOiW8z4ZotxU/1PQQWh0jx8aFN7UK+AWzxnFTuYXOX6DPRGhyo31mA7w9JD3E
91eL+dtVeap4neLWSriwqM7k1CR6InpN4f8ocpGnE0ugPdkAxNqTf/VkJxfYljd+
vQIxCntMWyagnGIaTIzPUSvcinuXPZHK8bJz8qVLU6AS2iOwMWXHerPxe5ZGSiyG
Rr99+MLA8z0m6KMf0p++XbjoclrUrehZXrnWsF0/SYS2Ax69H5KVng24bIu7C+fY
wsObAeTMrCpSp6JuwAsP3M2H6URg07z2eecDGhMxDtK2+2SwWRiSTmHYEKzSIAcr
8Z/mjhBH9RGywr+1KJH8k4thPfrq8eWkrkAnArG/dYN6dvDhs6z8UB3Zga9+Yf+p
B8acvFTc3DOBrnjitiIdWqM1OJRLNPNK9p9J2aNKe+73MSoTJkCXH2HXe8zOj8vB
R0poya4sXzIuyvhRu8ms342nfql41CuAtQu7ys8xe1DUVNWaeXq+6Ts46ai0p9dq
LvrId4OgumXjtbaZeCsD+kaV4ZlAppp7I75YFlamEIm6DpVNL9M7fCdY13NpkPwT
Q7c07ZSMdYnt/gyBt4F7EjBiGFUZ12rVuTDHAjCfWcJ812fECX4HNkEFCqveuplf
pRi1xjOON3V5DFp3jYdKONbrFIKbGqf7RDzDuBEYAudRDf931KjVgwoud3N5GQdk
Ks2ozSP31+3S0dlJrd+iFedoMfJGQowWaqE29iqKTOVyeewF63lWiUfkWrg+K9Hj
+5u2chCILzOKyVnStXqoj2WzHi2SPfCxkbxVB1pZCqCgCabY/e/LsrzE2eQNhMrK
dVB4E2VLNNqxwFhPSA2jmAfGuKcgTlIGVf165fP3mUk28b9s7QKHw4nhcYIwQXG7
9/O45UgexTw0ewZYXGGjKD4nD9+71J4ETaBzpvMeJQkN0ax8qIXjjF/cdwInX5Tb
oB2REn9KI0dG/gbmpNkV+yEs0WG5IUKXS2trsR8h7iuReYMen+z9q1qVrK8UKBnT
5Bb+c0IWNRthbbyVXW4/102FUQOoB4SQaATnZDwkuPM7+3s31/Fwm6+HFc7NFX4w
FBX0mGJ8WClbrIZFRN13KPhWaaqt6uPBSjn7IPo5BuS+DbeduHkbZvy8PClB+D6J
tdyhprOzy4LQe/rbwFie3OLL5cQEqh03azS2D+PhXH0gUVCc46cTMNaV2BNPxt5d
9zHpWrAoe2ZqFm5RTQtGdy6zH581npUF1wgYkMFiFlOo0NU01dnBe8JrP/x6nb5J
mhJMEgXT57QkoLXoGkb/+LEYCAzTnYsD2jg1ckjNae+q+cb6Lp4LKHkbKh0tC3nc
pOH03ot8IADO3+TOQqTHICcMBoH5jmwk0EMi04fRjhyiwI0w+uJrSWqvtdqRH4wW
JwoKsYb/ydG23Yu/W1PUYktRjWfD40NXUK3Bom0dKoXm2T4H04vMPIvKyxUMcMzW
8FpYt6IgtoM687ZiU9GzEOLJ6nz15koJeBo119U4s39IFj/BxWVxlbx++Dm0RRpF
2tzxTi2aPT0ANRw28wD/fXMYpyq+J5ECbQsNNHjrf/FiKEhdm9+T0zBWffUEGrf5
ga1PSYZ6Gx9jNcXRvzCvtCbOxZwLkeosuCdygraLCIJfivEzVE2J8ruTTnB4OL2/
m8ck7eJZ/T9w8m6eug8ogM30ugJLRpewqztJjlS1Wwq/WQvE8yXfv/oHLHjxKLrX
zwRbSe9qVKKpkXhtdPXzoNiOam2dh+Qv4U9P43zcmY9QsWl4A1QlyJQzLGjBA2Xb
ZUulM+hGC/PcqMqNGsiwbhwmFhEA+HjFTLnaf59TgbGSqV4DEpfiPVh653vI4FKX
hgt6yOoUkRtCw8a8AcsqzvdHGQKMR5KcIAtL2uKShQRNtOpIV8fEjKYGpUUV2H0X
81x/+Rqxnh94EwxVSLDo0qsYPZBUgeZ9Q4nV6Nq0Ww6Mme6qLbxEXCLOPRf5RvmR
aJ36Yv9fkyUm2JhCPKvCh5U50XnisAykwfzjKUPPQRNlkO1hq6+roiuvujWgjn/w
VbDURKN14oiVy6VI9lN/YwlngbI9RLjVygSWhjKJCbTUvdUlwEBtiNDkwrJNjFCS
ER78C8nBpZ6arMt/Mo8R5gW/XyXGIktgH95+FD8iZC9wQyWqAY1P0pMCL1glOE/z
F1IkNt1Hog5amMLt0jOfH6NHQ8wQqX7xkt3+GePvF5nHXQLEWRUeyDwwnPHcCTPl
ZP1UAipb/DhYwBin9eOhn9qCK1tMBxvYPcjS1l5F8m+134OTXH67OVcwSMdGD66P
42cVbR7ohvxcSTyu2wC9y3FtFP3XpKZrwFD2joHpJZAhM02TvS9t7tPWz892yFgX
w2W02lF1a2pH6449fJt6tlnXXTNfrtD5GdZH8kxpjuJSF2sjgNCZyPCAKhPoY0Vx
xehAEnV1p4w80rNZwFPeiE9Uzp9sFQtuJXtkZR8hLFb3kX7c1jOtYH23AVohJtK3
+eQhWwM8lGtXLm8qRyKTC3lBUEdNFqcqtn+b14M5pDCC0nYJXy1HuSdX+tNlrdYd
ygQmubDs9DuOO+3MnVLP9oCcF19f99WJ5y93VhvLwPXY41Ab0fU2u33XIpH9YJKS
0O/hnh4yRMd3rRs1DwVml8FSno4U0EvH1mXII9ASTD+0TcZcOg6dfJkAz1Px7kkC
az9gZsq5FEN3gb9tKHTJzWi25hrpnl/f7ALgJOV8/mI6h0zDyOnZb9wNsP02Siqu
oNCVBXMqSJaJcLzCV9S1XyoB5A2HrilJ4R2HWXOI44NrR6Cz2uLoztpS9zBWhYm1
BxQetSdadhHDEnvqXS/LBSs/AuV2l/WFo4QvzTvWc9bcmm2sjI/Ijg6/27JZ+B3q
4ai1lTGdNNVaEC9cOT6pqdaeAen19T9FUpWNSzf1T4HkCGRT/GocAeX+dVBNrkd2
21Q55/0igc8lzpdLcoFbKIS5eOv7iEYrXubffFEQai2D/4NOsE8afj3WaPteK2tf
eeM5Ghi5/DxcGFekfoX2siazpA1GecHwZ2LkGFQ66Zo5m8ELj6jRPtVBQMTk2X/1
NvAMRdyL5ewfHvqncaH7eOYwU1J1f5/Q6Z1Ai3MYWtEW6GNb5ly1HvZNbOm1mgDu
y/V7hSsjh7CFThwebEm0YfJthc5+ts5wwThA1eDAk1DJk9wBIJd1E5sZgQcMCkFg
G4CT2Z+HScGJVR8+ZVSz+3+EfBTGeQHaFMjQFrnLT620fskKq0NLWnCk3RidT0rM
XpjFMrtJKJnX2Zv5//QovtsXckD2J+V26jo3k1ej+I1aLDrjaO08K8TWZ41jfRC+
vm1WRaXw1AlDrf55rrJRBySnXU8Jix3RIEsUIvpAScQTdvOJJYIQvbQ8UYqPCYIE
j+npUB/F7f17FnRHqWDSjz+z4k+98DDGEtwHrKOqt9PcaJwiJthch6jGbyJrGBIn
erai+/6SDNX2JDvEmA+wyJPI/Snan5109hEnpiQipc1DDXhfBiGciSe+bcII0/3h
bnRIELgq86oYYhQRq0AD8U9LiuAKtK9HMkJcvpQq2QYFhc2JL97jskbP6jcrm+30
/xNkQCy+/90e7JJk3/IsdIAOJ66JjXbncZ3G0M5fyf3QO8gByc7ugki41UiV5G8F
EuHnlW01qCR4F1yignDkGIqjZXBj/rTrRo1VSq20fLSVo4t6Ej12Uf7+/cX7h99H
Ilnq/mGcRErtHUEwJr5Ozl+boYf+Z+9jIWanPgD/N5GKIMeNGinqBV9INMnaWnmP
HwZRsfohc9s/hSe8WL3o/beqGYVf0A70VVvfXK+LGotUS9ORtwkirbEQ9Ja5Rdmg
JO9TsiwkiSZIhWQIEQQZ8xedY87b0fAoaKZoM4RGXSmTBPzg+9z/VAThHaD/mybM
4xqUXWFqyQH9sqaczJjlkIukMrSR1wiPOhq3SZeH40xkNdumQXstshmZo9R8Gsm8
xMxN/z/TMov06uaVb0XcNN7Lt04kUOA1fbToFK7vDgpMe+9FP6itwthGqcYqgksq
vcDYdPNat2sRG+rcAF1HPnddqgmQXiGtAUr5a5L5Abq8kHB0j5m3WHXLsKzcAI8s
PfFno5FDzDRxnVzVP3/gVtpC5IWCUQEdzQTqY/K49lUg4BU79ZExQnEml2SDjydz
DOMiw8gkJqpFueZVNMdcqPa0MxKIoB0GHVAxaoUZpDMn8kgGVOw2VhVWoXrYGUfb
jKm+JLUph5cfqmMS8BGFVPcKiCwErToHZdI7ol9uEQ4TeogL4cWC+uWsjBSfRnBJ
4JyUHHR1/GC13zMH/XnooXDTeC/I8zWVhrZzZO4Is3YRDu7C1mnoYGoNsPATTdjZ
0FzAeaVuURZXPY0Dw0WgLVeeC9RlwLgD6JvZffcQKr9Gwao1VyeqpT7x03zpEepq
J2GcAHhK5L2eNVoopj5zlilXqWhxDb9v7IiAQXCIrfKuN5c/MKa6eEbQqVKWb2op
CrQakrW2994el0RCIBaIBRv2BcXDWScAbcxBvMGgghO158S2B1hcMjp9Am1RODrf
hccb+p/nnP50I+3zQGJWqgjCCafuOcWHKBa1YaSjfhrPzwf8oncGYnvfSVQQB9ah
9pX6CkI4OrSVxj32lj7QGNSLkvXw+cA99iGkbQYtKfL20C32ebbs9Iro8dvK/7aR
phuVOYA8+AjS0QmAKHzRAyx+WcL8HQe5JHY9qrayB16Iklmbp1PLg51pUxMfK9sU
O66j71bL7oiH1wczGSr4psNBPbPDXP1vZN9cD6sCqoaad9ICi+Dil67nmgrNOdz1
fw0rx/quQxbukezIcGLWairUODXGxMhHohrjz5GZo43YZuDxB+0aswMZpNkQPgxC
3X5tYJaIE2hNhwLmiEfl2Gv/5YrLNL2SSmrB0UqEPNkKf3TLHHIfu6Xe/uRO36cf
++nZyYvjZz0wtYNq1NtVUQTzCcPKKJNKmS6TM7TA6INzubdQnTJJssLV3otlB/XG
3+M1MSrJgbpRzXnP79dMfvN3L6pqEs0j6TODjbqoLjKAxMsJNA86gSPPLR5B39gl
9FsXNjAXYMRC6OHD12ymC+8L+P3ZpN/wZv2yjGSWfK5fz5WnbcykLqBxIsk0EO1y
iMqi6fd4ncuJRVjMCLm7bSukQx4LRYh3Xsz/OqbOZAWszsv3cuHxpRrn+CceZp48
r+BuOrTsSUv2dL7Lq4gNDIc8aCpckVTqpMQfkLcpc/mstrzjoY96nN6fphL9+Iru
6LbpEmtjfQRVf/3jNFkC24qKlzinriTKKblVTOcbp1rKhgPzVRRgE/UZmXodBUCA
wx+rr7F2OWoKIlE60R5CIut1HPUwLvRbWOM4nVywqDdV4wssyxHcEyKK2wGuevNi
Y6N6ZEHYQiFo1IuT1KWsbXzSFEf7SraN24f++2AUJnGj47WKzk0sHqbQLanYQjp5
9RlUicnX7vQqNfsEWWS0EO7cMYgUAKGB9PU1lw20om9g9dzaZV/kqaO/yCItw2R8
iveTlHveCuV1BKQ5YRcnl9Kb3Yiecc6XD0EvG1PNsd93/1bQsWojR/chN2Z7mMPb
CDaeF3MUXbCmj7pnIMP5QjH2VyqWCG9SdLQHASF3hqc06JwEUI9kpmQTYqVD9uAy
2eFDrAwFt+eIydcaPMmAkFkATGazonHUBiMWGALwB8b53nybiuHEU5tSuiQ/lUEf
xB/78E1VunT7BVjlJ6c+iOYigI1HyRiVtyiJ0Zv3qitNOgVTXwTMnVyHSRmr3Yfp
DtYfA00gvIfeBhYOsbtDEeJqMp59AICWuY2SnA8yifpJkJPGZnbgJi0OgtI47oXb
Q52BjHkByvfsuaxEigdrvkfMrtYkQ/qAv/ThUXC0fLBDMcaimhC2Hmx3Z7YIgHry
rGqXGfKeoMjdwGv5ykB/KPpiBkgQLLerbrmPRnOmXlttuaI2WUI2nDTFzSzw6NZx
anOGKVuqxsC8ZP6fNt7JTDzxU9dcN4hUL0A3MQmolbswTwAZx7mwJOPJcHMWYZC6
ZKLnMB/1dDsO2c6C9ea59RUgBcwa9Qf3HRVDH/cO7zbF+EtdN1nFctFQnHZHg/JK
ewPKxS2LI4uxkp2zcw/cOGQnS8VjMOaVfVznAThy5fb+I4tRcymdDtVJ7jXSRwvc
W4cnt+b9szj6UPS/PHMbdl4dbdpZcwn56ru1IKooY4uezChQY6HbPyefg+M99Hhy
Aa7Ff9j645cqi8BovCIf82eoha2rPRXOimQa15SeadZkIKcgDP9qjYka+Unl7PTc
lOOD7b2+oyqU7hs0Wg0c5zEE5I10T93+cc+xZyAq0O8YdCMbxYBeP7FJz38ykMVs
ZQE1jU0ZXr6vTeATtR59z2YElxde2KzieRU3a/XFx5ZS9L8Z14AoQQvqHXv04khN
9o7Q8NHZeYFuc5rsFH5a9u0mLogb5ka1ibXjDh58XD87AZKGKn2VK+PTPe+E/BJV
0DoZIB3RDxvsczr3mWloejGZBqOTCLgmthN99KttSIBTi86pmCQ7jWv9olr/mtKs
q69g2bFS7sNVsDARlApMisHD5HknRLnhkqnkdFA7z4QJQkffVo0vbKl3ZGnjME7k
p3W53ZLAGfgLcdMcg78mJxhojYrEpZHmGN7HbQs77N02dfd33OuJwi6hWmUR1raV
ee029V7E7B9q5cgp0A0Aj07WlreHgGF/H7MQ9CYVpczBCQAHUe34Qf/1lec4FYpH
U39EHI5BBMkym6nF/6nxd7GGQNsNIBWGfAHJogNz6P9N73y8WVtCZO/bd8H60vAz
iOv5hT9FfTv/HTkMQVrpZqmV3RaDf90IKGPmSdLw4RWRifgM3HZSZHwJk45MLIlU
BfQFZykq5s13FLPeEOQKAlCYwW9fMPjwSLvkt/wtK0q1Fp26ynkR2SJ3j+13j86l
HhFP2QfVAVDmWY0pxcyt+bhi5A7y1xZvKms+Q4x7A7JWnu3PGdOtR7iXOO1erzND
giU8iWGTcs/on1PePlzDTxTQwSDUtDu0+Dz748Kq64QQqng1yN1H5tnSUhQ2oGpy
vpyF3oa2hiD3Gp2p6pBDqbVXRp4snuvJQff/dW/MjUNEF3Tx5UUczdSf8v7d7Yge
TUYSe1DmasDIiHI0J9FDxKuzFughvpZqxw5Y6KHbiIDbpg6MCwCw0Gd3aznD7KbK
cHPBS+qVw6O/eji5khu+saG+rPBidFXsO+5Y+EjJOnW+eaqptUytsMtTqxozi6ZX
jCz3v8KnEJ/UzQj09V6C0LvAqlnSSGXly+HtU8DAllXMGSI7lzq7IzETTFiJYHUD
3Yjb8i/UqZqSIOd8rz5VvPqP+rbQpvDJhtoMpvuYng6gk1Cq8L6X/Sohr2DWw0yK
Ybqrui/hbWjCWFjSIkQLJO4QMzqbg/zx6FacuhuWz9RDPyHZsVWt8JMFZSzp6UAq
rKrDqmM8m2V2YjfjI7rZRk0Ogtkg2cAKCp4Wt9Cm0qKwz/rVY55yMkYYJQl1Q4C+
vLFR1ICJjwG4Q4zvbs8XkY98KRb3yfycGvIli0dqG61FVj5Z4NmSjP0MvRc1gMc9
fmMtdAYJunaE4Moc+wx+JyPv9ETD6ZduE1m6zE4ZOGYMqymubNYVcvG8Xd9ftBMG
fj5TaK57OhbyISAcqfnQ8nclkmnA5tqCwePRn0UMGOoicHoEMGhpgRxYVt52iMhV
8LOEVBOzvnP2B+/WVnBa5fQoBpNhhwLvDiHz5GVmobNz6npvqVSP+4r5u4IrnnJ0
01tlZeGVs85z3SLSeBBkYu+o/EYwJ39GodoXhiI8R4ANLGatNieRXtIl6qZcuA08
xXJPyOF7odK3B+Klgcwa6WTyrTAbDeDnTENc2Ct3wFdOIoLb4xXrUNM+a34/TsEg
+VQJHBs3d9L3fckQjYahiw/jLsJDCXI+EoSzHnlrTo/sDweOEFj0/UpmTpTnRXW2
ZCxEsHjJKs9gLrJAqrSwTG8skLvXik451iH2/E1wI/Qr8j4nTUKmgo6Emj9GGfaW
s041mXYa73eu8G2stC0jC1dhgRVKoxrOF9Rmdd7sh+664PaqUu6xwHnYuvm2kfhE
qLybus8KLXaR5sz+Ik3dLQwdh10/xcKfUp1+9iEWRsvCalYkydZ7uW5/40J15KEb
q4VVUNBoQGge/SbMXKePv45BMRvTMYDJxm2MOtbcEalNrfQZZOs95BsYjVkvZg5I
+jkW4Ge4DVY3zAffiaqNrIsr4UQXoyjxm96Li50ZnSbzrRQXinvyh1PzKVbGsrzt
n+Dr+iufLi9bDNUWkenpafaNUTV/vBkUbf1C1MZQIJ8lIklhbDUTfpOclrtTj6Oq
pFHjc7zXSixuL6LcBXLtksrjk3XdVOSu84PN8YhZUh6dn98NgW/vrksaKr/X8gL2
ytE1Jw3nSCFb2SYuBiEPDPW48wp0XXAmD4acehj7jsR4dP7ZrPrT6XRg24ZQ1zzR
JJc/JpZRx8JUFkJ8lAPY+Zr7xcYtzlkanMouuI8GkL6fV9HmY0a71sjMK+IqzKvW
H3xQbqfd8d6iOIfwApAoxrGPtu+5sL0WQE4RGWYyJ0Tp3Ax7fZnR5+Z8rTeLV9BM
8w5tfnwhTlttwQPv77pWEyRmG2Ehp96D5RqBfO3p5he1fuAFAe2W6AAO1fBbYbPw
EbT33/MScEjFV9P2VOqL2WvQmX2vEeAmaQsn+MlKmwfVaKFR1N4JGNuitGyCmCUs
7uunpnsCNnnKPEly8XSDALwlFc+MxcPEiy1515Mqv9GBucxOte4EbHd0feijr/nF
O0bHghPU0/NURsUmJ5apyJVzF/SsJQCviua0408lHoWNUHKDIsNVb08XdgxjqHeC
Nc4tkwCmmTtNCFGqXr7y0mYVDgEn8Y+MGkZOSZX8lHfpbY2Wtbcdp8inJWNtkemC
knTQHRPFSznU+YbWJMF82w6TeSOgAkwgNcXm0AKH9GufGmBoZeUMHBKgrRATSUPU
/pX8bewhApzkKum6cUE4C9FhX47Kr4upgJFudGg7ER83PqMQpG0Stj0zX7hafqsA
gcOaABrGPg3vLoUa5C4wowCPCbcwfvMK/UHQN4iS8y8IWqsRLEtRU7UJ4tkMOGRy
TFKXdBmrRKThrgN5XR6fF7cKqy6OpXzkKrAGPLOhd4eZhY25TXFjj9t13MvdhKyv
XXYUD8wqTHGNFNLdjZlx3zMmyT/cRdLTNnYcwOcy6j3W+tW+NFEjeyXG0kXBvOi2
/XgcFPQW7OxFS2LJ+Lz/bPNHfuWEpxFfP7zU9MEY/PFNBBKhgHgNd9/syWu9HxSk
LzrJPeenM/qPKCV4YvRN8GsQ95XVo0QrZZC/F/Dgfq/0N/WnlF9b6sxnBpEj12Jg
MDI8IZCANMhG2ifEjCh0LnyIEoIT9RRcZqUmx7BiR3Y+uoW28V0WszMDaF4Zt9r0
mlr9IIbv56zKAlE9N63Adq7eIA0OY4SUVAKFLkEZ6EbT4z7LK/dewr7NLyGScBro
VOp1rDwXrM7pElKa3kvUtXTTZw16lFC2Ful1UXG0nCsoOb5idRyJaBsBLPWcnrU3
dnjCyJcVOVG9XBjdONjjsL+NJhXGUhtEr9/Na9jhq9veWepzTvQoz8XwVv4obPFT
gsNPC5O26qRHalfWfUHEjldsKcTXntfbZzPhGvqjg3qlqicS4drOd718JNV29D6e
5AOfNBUTuCQSqJzIIURfrezaZ0yTo7L99TOQ9RjoRUALhES1TubI1vudpSCRNnV7
syDXu5cMbrBzlSwKcCbgQEoSL89Pg4wXQ8Sh21bvb7LaXapJks+dSCCC8uSIRG7I
Xck9P4MHRioIs2VTThKLTnsC4MKhpxD6tNwelj6AHe2xCbyXratQ6aTuoYukEYWY
wu2kWOhi67IuMBPKxRTrWRxKHZ2LHMK2Q3+8GSlmqERkT7xFIZsEp5um6LE+BPg3
PlmQCVL8NB+HmVB4wAY8hhyBQGE32j2GSN6YFN483n9GLmioPqkEJc/qYeNODpzl
unBz8qewVYlNZuIfLfDDkt25TbLRrfT5h6kVtLmlNGskXvBCcT/x/HS1QKjkeRPF
bADwMr0zViFePQJgJTpdLsPnCoU6gqOSbrnTkzZmigfXsnCCKobip1uW+v6blEKj
qeM7iM1cweK25j9QX+7bVGxqGUWfcSBKlBtIFCqdFtpoGoDdzuaotwTVdSAV0km3
TQO/96o1KUVhfZb7+dKJHcHeyBkZJXUZ0QIJYPujyCybz24bChWadQn6gHZuF3N7
Gh70I9nP3Gh8tIxfYjGDWnfEaLpNvFaTI8HCw0RMZ3mpZ1SxJIkJsl+51jhDTCK7
IT29iTBdFLrydyJ4kTveG2Rn3bcHXv51FTTY+o7PS+BI9FSUjheBdUHIL/H0GTy5
PZGzbDx2VcDTbHWJ4Va23vYTCuKSed8XE9H7aiLmMjbqgz5mqEqvHcU+dstP5p2O
S5XIenpxR15N+wEmV6Widopa0/1OHajPmwK1WD3z63ND4jIQT2D2yNp19s0RoCrG
E95u5E2EQB4taN3O7Oau2SkAJhtg2MtIf5Zi8gFiUBBmdtRbVtp4fO2HEqMTRfMX
e0jCH8BoHe93f2OA7HfY1kFLIJoeZ4BhAI3vciRwLp2LRPfyppi+U1MJoM3kOt9w
zDGYvpXYO0/xPRMOrLYXUtclotjf3W6ukLPsKvEuGDA8U7/So3QjocvHE7eGzL9t
yIPHodjkeH/DG/riwgic5aCpSeMtTqiQ5BzCh+Crh9Up0KcmX8AVC4ThPqdFHLkU
CEIA5zxcMetGqUflrTkWwx87SstQIzuvoLxxs7xRDGKzDitxsd8aDB0OFMalP5lL
ETiYxgPNO+ESJ5ydfEkQGRNr117PkV23leGhECPtvmdGJbBtdMQdTZq1oYbYhh6B
YDtpcT5TDkSHy8l0NTnIgMld209fc0V3+Rw/riL6BAqXDCqOuOnEB+OeBH1WsxU2
mGZgIrhM/lDa4UoBksrAo1uqZ2dEdm9GWfU/M7vTURPruxEH8ZeZscKt2dK3W7MU
tFsmBthDIgA3cAlexDV1Y7xuVaPiVHqCRckeeSWOMxQFPtii0JThIKep8RHtxeUz
7nwdbk5F5x5NAfQhoK7i4pAikL1zMFvxIcbIhI1Yjjeyo0+lC+jBn5uKCvTIYnQC
YKzNjr7gcTAy8EBpNhIriJ6B4XQtg7Z5EIx5LFM6a6CkU6intCILRtl18UZlalIY
7+fa1hk5TqqqfEkC8d6AEw3QL3yXbzxLDQdfXyOK8dd1dB4Pk/NCh9ZQkNyS1WoA
wcNbUv9pgNygi7fD+LXb4xT6d4Zp3yRBch0jpAFDPcXYTHDN3WtMt7jdv11rI1rg
TiGFkBDHAtxVzkXktwiN2NNhhDbTB9sY2jVfMKeeeSQD2Tlvyei+1rbI3mh75BgO
FRZD3wMy4/fHAWTmfCvfC4W4AdLDxcWBcPUGmWu2q5KiSt1ynEnZYPyprT2L8LPe
StGjprdDZq+AGEyBfi6oIacZNElhzGl5ck4/ucgKadY/FNRflwDAPwTimWqfM4oL
69OSdQoyDcRvKUh30e8hM7ChpZ8VPtdpd9BtkR7Z6GCIUuqte2TT5yopa23dQdb+
mGNjNie1I2lCRbpw2Q0f46AJZuDTa/pGsvFTByF9HfCGQ/W8Zp1Tp3tNnHb+afmg
cV0d2RzouG1m8cSV+baRNznZn+dfjCCYmWVVtZik/t8fMxM3tfO50243viseDCIL
KsTD2HL1v6+CJaH8L9boODp6kp5RUSjMJ1idRi1F5Hpyj5IiFF7NmYoFNLlzrebn
ja7SivVUqfKrzPzbpW40Wl4qJpa1+pt3NXgAiCuaCNNNE4AeFJcyZNUAGX0eZy2u
kk4bYcyPNpIgMZ1t4YjnyFpgnvUGEIidQeNmpYyVwv1mlezKu9ApK9FNWPVhzdJF
L+12ltAE9ekNUAv+to1vO2cdcghWkwXK8C9N2/TCFClQIxmpQb1fryLeVEPLoyJA
L1xkWiSsGWL/Y2Eqk1t33HWUXOY8PJZdADTHVmKXKI9UUToeGCZCHdGVxADoMQOn
vOZO7/HLoWPATeaeh344sltNPo/qDK/KxmWKrr/Wd8pmNHGY0Ta/s5E6EO2vWOx+
bcZx/sJk+42UD0l+fBAhnppV1OCjgRbJD+FEXEH4HXYXUk6oqU7Qc11KOkg6kk0l
8AoFyHEvsHOerB33VuJ6sdV98GrsyA39Y7Oei2VvxakIFsfF014FwIdI4d7ZesQ7
uzFW8d5FOQ7rsg396EaoqHKaBn3ZVp1Z+hptZIpP2uE+8TCHv6MHWFRBg3bRNxfl
y2fIptzFmuBljwJ9B6vcPxBOKTU8T0PioCgandedfSQCr/esRm4CZYJPydGEoDTM
nSIRSfDfWZWcIN6Vz7y5kszsz4oQptA38PvDdOeq2kOqHMerY80Q1tRa870cd+2h
1FEykHTLBYAPAG+dK40JNyk6/HZQBJDeF8K2teyznh10P6cq/G/Eav7i11dm3zWg
7/NVn+YZJvVB2VxE9ABAhKvRhVfrkGoMgdTES6vrPAoJQRIUFOyivupqrSi8xfDs
npQ23U1CyC+9R65Jzn0uD4dVK8V/nyX75+NjmazVTVdzYTP3y1KYLah4H/lhiV+g
VCvpcQYwKXi6Kd715k0RC27GWusUZNOYxIHogtW5F46p8rIqPsaZwmr2oy/ZSbbe
YvFEwjEwbKulAAVEInEnzt8U+afi7bbQTbQ49LXRm/r4SELNDf0JvPcacqXcrBJj
xNnmwr9WDEx1Qw+nvtnIZWDNp9zRE/6a3mSf6bp9rZr8LIgLyNsxha+fVh+QfRle
ZpCR0lbEr1UQ9OWqCEZFgTXA6IVEUB370Wbr1r0KAiUooHR6EOxTO7K4+4hZhHd9
Npb09PnkBb9LHsBspkuQXI6fk7u0iLbsP1WQaBUPiBhuRgOoSCb0GLncThtXNWJY
QPjCvK+K6BFjwq8+/2rkRbgeiMYBydjJpiXIECqHwa3peAyUqJl206Iv/86T3GO3
tkApEhtcbxUHcuhXsjq4YB4Yfwb1R+MSrubAe0kVkuLJJ51EyK5pxoJPLwGrFkkl
3jgRZkx/GSwEs8ful828WqRrVKHHB/4TTAnKbKJ/9a+g8ymOgc1a8oHNJNGaBPt/
8dWTFzNuT7oOjkPRThb5xuMwH3HLNolLVWGqgpdWxWlkepy+G5Xg0Y37AG/qZkSn
KcysbNsT5yYJ9Akzwo5sKNs0bJvNgjnMDMh9mqNQHpMGf92CK2LZ3sPwjW+3o06i
sQXWYGwFuuZQwBoN7v2hZHiwNdyp3Y/jFgSKFbkUHEhqFsCjsxLtUhmD6Bpel5hb
mrjPNWk0O14BJvPxG/VX5FLNKanDwhwIMhedBgjLLkwWGtpw3/436hdsge/aYj4o
6/ZZTEhuAWln/LKowLXPGSLUPh31925fE7zYg7JmHzcPpeM2SKTAdWRs4bIbLdch
4S4BnwnwXSixme547mZD8iTVL4eMyG+jrSTNMPhTlIN/o+BSEbRpQCw/LjmLF9vy
AxT3asZwzZiyyw7ZQZTPuBiecfRubwDXaK9UgPE+s5lB52olTVzAH+aFVCnnYDRU
i1E1RJtnHKVPb/Yh30IXU5qngmWpKA5CX5JP3uz3H6GzzOqhBI3+Wl041p0I1GPX
jdd+4kftdmd/SRc31BWhV0DuANx24rExV4kxg34qPZaeK07fnYEstKNUa2EveD+Q
BUm2uwHqeAHJZM4A6l2NI+VKqkMLFxaWcPSJbwAK0wtRGADG3Cph6KO0+Jywhqbu
pbZcp7TscQF2nLaCsl1xUC/0iLW8TIh8S/rRSOH62LKvKCmSUbTP9ulM/vAiaOm4
4PBHJXRfiXNiZqh3MWG0B8T8iR05fB4r7G2vT6AmEIQ9f7mF9py9bFfz8d9MpTiL
7KyVMconPqQeHoDbasDM1KSCEqU5jJTHskEz11YP+j0SEh5keYSZp/pgE5LNswUp
xCcbd46/Xdp0lhmwjx+37QA/gWu31i8b5bxRVVHXNU3EAab+z2FoPVuQtqDrvrza
mHWLC1pXoWPzKKDoYpP3/8N2uFucvA0ZtG0YEeSbOrirmw+1oyJ4xv66AWdoeJYp
kdTAHTagjf1lXsXccSYVD9v1bNYFXd5JNp4V+A0acdVwOFdyM2+ekrIulpfUcqoN
FqbcYH2xBXChf9Wx7zZm88TmKxath1tgSg48VJUsAsx1EYx6c+32WbNQlpQm3z2F
Zmja3lLo0TaJR/uSbn9smPnJ8nJbKsdp0YGubb6c8VO1aEjVqLO/aOy9yZg59Zp2
a4sJIwoky2qU4mz8IqKn/hlsZxgTVMzHACv6R0h62Ob/pAISpNAOEIIYN4OqMReV
VhUxdKjLAP9KOQ/QFfJLvJibGhVsPIXcdrIAqXZbBudAxlyvSBe8OkQBxLhqP8A5
uI0NKn526tHGqqjqLkHNFhkuqBMHstbj08WyEMj0r1HEXDE6l4phDTtIZPVwPzJC
Ah78BrKZQLaCWLCC/ZP2uZ2J03LK3cakZXXLly3f792yLl6iKdhW1+YqAe2vrFV5
6RzfCPZS3AMowzLK2ftTHiHYUJ66pmIX0NGU7+S3xVIrNF4NCXSdaa1mfj3+v8GX
jS2xAtYUIev+CQ1UF50U3BSYIaHb2SgjqOyAfM3b98RUbipY2ClS22by8CcG0Luq
waARyWKMp8X55Jaamgk52O11TKwzVizruP33EDBYQf9TgrXISauL+TIll7Od/5mU
sWYSLNDxjWdu8FixDHta+CAYfnURRprah4J2fe9kzoK1KYLxN4dAScS6sbejVxfE
u1Ut7htONjT50tkuoeohnL3I7ocJzTBnvZMToQm4x5ItBvi1F2wjwBjFbuJKKz7R
6AIezp5H7uIiYkE2tenRLhp+tLDSCHCg1GovzQKG2f7HB/DUSLfRMplxVQECvJYZ
nUjriSQkbdFbLynpxeQld0tJDfARY13RhlYevCe5PNfNZmeWMNYvMhBonO4lkI7A
cbTXddq+MJFOuoyc+pKHHfi1Lm2uZzcdzI+q4cMkstYzkn4eUPKZV+Azr/Cqo7Bs
5OIp4qUNUX5J7Me0PNPlfdlRuckvHPyK8I369R8RcSXCWm5lVzmBAhKQhoTQyAVU
l0vAB2Ne6aQ885xse+ZuYJwZLxVelzNEZySO/RkIBcMhwMb2yoWaE2AxgDCKVqYQ
ZABupuFjgesdlF/RD4L8yTARbxWVIIHsWbnBHML3Q/dCedrvOGEejtqIaD8CUNkA
auRfFnj9KV1/sLiYocaZz1OBmOV2J5I5PYfTS5FHdf7wr0JVMv6zzZsUcQ7u2W1L
7uCzOSKR3vh7XtP3F1zUrZIOyrg2t71WB+8P/qAd6EdgvjGdOclOU3XtF0stJy2R
q7G2Hc/AS9wgymsyJDVfZY4/yXrrqXEvCavxzIfFNSSt+jyF1Yl3SimvYuVJl63H
Mu5933I8uaV3fCaU34a+sQ7bA/6yjrtA56TnWNMWF57/TN6eOROsUs1bgQzHy98Z
Js4j/kSwp7dugUiUZdiklEfENtXa3Ysx7mB9CqM1xA2P7oX1X87YkADwCHy/e/Rs
tGfu1+W4N1gCmSuVcrys9SdsI94EctzsChBclHZTubVTcODmXHKH3qlFHqR1b+mQ
6excNJiPuGvSR1sVT4y6fx62IrBYdm0Qz0d68mYBR4i/R5/ZK2aDqtxbMdT0DpRF
oF7+z+umeVmcq43k3AUYi6MbXCnqIdDcuNKrdbkSUSZFhhU9whl/yqiGTKPUH1tB
NIpZqt+YSO5XQjMtDfSAt4/F8odAbJ3qehmXSxjCqQnVzG3xagEvEfAg5rYZX+9y
hgtBhWPacMm19QX4pr/vHdPXDMK+SiDzWmtsn0XKjzNUhFP6dx/AlFoiddRtf53A
Nx0looVqg4xX5BWaGXfh1iE9oyYObDlxmZNn2WLU/CUNh3/HHTnYpDEaSnM4fZlU
HDKr8QiRGD0wgEiSESX9swrUXUeF4zCUpLnjZiGGvzIEU9Z0E7amh3wcHCHPPetQ
HBuS3rVDnf3V6D6a0Wh7KJ8DfoSL2VsXJtgmoHgpZwvD3J3JnrfiMykTOf6PSxJD
ap6OqmA5Am8mvVx1M0NSjNWeVjyD5aTLqdu4vQZq56p8D5GmTyuih5i2/ki+dvSt
InF4QQXq2+KgegQqA/D+MHXPdQX46ASn8hZRIi/WOvOguDcz7UEF9mxRPCxuGoJq
J+4AARgifRgo0yJG2oanDiKcHPESUnGzf2Yw6jwr4OBXAMrhG4NZlv8M8ZQh83/I
liE5ng+e2htCt3rbX7euH5E/XYJayYkYHMnD0vM6AjqrIXAHDZgc2dgTQQ9c6u73
vQVuV/oVHT2VkX2j5+rbuTJ8O4VA63cv/IBSvvxfXZjiI1ABvv5pLB6hcwztUKit
bRAdSqJXL2RSCu7xDZnlaLlmJR/BEQFUvd+edx1gBp10W+M5ri0Bnzq1P3FfTcq3
Aj/TwpNLseZOU6vnXjzO6hmWs8WVWcIJmaPWK8j+lBSyaybljG73y6dov9MK0uT9
z/OJwmV0ehT6fpY0iUKCWWp9RQgLzUWcvDkv6NAU9A3uln474fzSqUvDaRFibWyu
lLvS+Yfb6n1ZfoYh4Kt1n5uGqBqEws6D9nk6gtydsjMwsCo1rJjcMBIDz0CDGCZy
/l6VxTztacTCU5DiFolkC5zpBTgqmpos4zlrMFRUFxFQWp2L4XsyBzrQQwTz3E5A
erO8N56ACvzmueqxfiEdOuwCD8x5EuMmz9aZfvaMbJBZHnLSBftze4ZMvCgkl6Bl
vlEcbEsuG8li0b6SfTy9q3GmIb4wsTGQEyPpuTkTEltqih1rrB7fqbetCne/Nhpd
AkkbSGRQ5nYQimvj+vuRivUYUj9h7w9NaIAYDMnyuPto6/TJg50ztw90lEyvWt/k
vzvMNBqaxZcLmzqEMcBn6NzCVTlL1bd52y9Qm0LHXWzk6knLm7BGAWsHCmq2+80F
UU8JrhAnzBlIwlXFT8QTXJypfIBbT0w5rscqPpKMqxUfWI6rbTiA1F18OyNNScpn
LQd44qvxhfYrNoP2nkpKxki0BBQElpnsyh0x8HtIOg8RJ2Ywkeb4KbLR594W4eLp
4nCTu3nUPb/Tl10XS7z6m8YiieOE4VLaknhYD6jfpy3rv8XIImfK6Xx3b86y8yOF
1ubm0hqLE02l14hrWnRXWtqSF8bemFlLKc2/YFJ26l9FgQCnNmwve1Sja+DvGALZ
XC/O86ImcvdnRZsS6cZOL3hX2NcXOHAJZyxRcU0fisdbTYxPXBnghmMSEZTYUmhw
KPro+Z/eCL5w7oafoBig+Rk83+0PDAqjhc6AqRabIeKoNc2kT0cdlOknzjli/52n
I1YkqABbPsr3jxXteF+lBOvqcBV++KDL8OAJeLSP7synbPGfCsWAkTAz64LLBRB6
gCuo3wTzDtRTaLYVduku0xvADakNmrQ4QI0b7d73CmYt9zgmGisDuQ8jPEmvvR7B
zHlG45AwAdQj9qaHz5wc+ebsEXPbM6YlW2nx02ljrPn9U7KOtIKfNXDdGQGiKfBF
cWAePXfoYEpGIVTx1NEbM8FnJFAJ68CxgOAdxs/EsPiVnI6faBoAv1J0VNirLBIv
FGt9PV7P6kB3OBHnU2jl2WnAgpWGnB6ENMa7BIWPPxK2KnG8NdNVhsH0IDJdWWPM
XspqliiCMdK0xqjgTSbJw9MNhqBJrZpHYHygyhEyxRYhz4TCuC1VGZk+pWQI8JXM
33FjynNlJfHJ3M5s8T7byGu5W+p34WThK/04jByazkLogPOBJB5NBg3Ha0uEc/m3
uhcK+Kg84DmjJzSG4vFpuVbftB4ELmrqWu8946O+uGiR+7aUfs5+mZzKlX3yDPEd
3Hk5O2ApVqf3KcgUNA0/25ZWA1wamKNUbYBDPUNsP4mCSAI5t1HLbRxS/BBcfzTr
AdYDwwi2G3GJ2gubLoBmQqUXZclmiqKXP9IhnbidIhYhlmYVTiB+vIq2RT1fYgo7
r7hZDSfqM7O0XctPIunNe2MRmyiJMM4HZx6GtGP5AePxDTM7nj80W974dXthpKpY
BJ/CYOF/9mEhJbzTMmBjNbg2F4sb9BbbVL8MaPdLPhK1lWCf8Q3L65AzTZWlpLzT
mZSvBzWK5UGI/pQhIOMqOJafOz73xi7IoeXGvJekEx7xXaupook1+M6QGV4dS44z
zCZpDhwui+vC6K3l5a5UTX0F9C62kOQdC3k9k80wZ6DoeEqbLQ3crCjqoTTrbRbl
BZjV5nJtJhKaD2FV1tpFAfkaenibJwp3hoSp+LYx90gCtoYdKwLSSdsTT/fCTW42
drvShzDvrpU0tHNkL2ayvUPgjK0QjKf1i7gZNUt5xL0RtU8HYOCE+ticE8Q0s4/C
B5qX0IcQGTO/M+i6Z7YzydTBpJAT9UyrR3VHFXwnI73hxyFGwRO7LbheKl6GXgrR
4p0mGwX1P3PlrJhNJ+L3zVkjg28aX86CE0wml4a+yqsKc8Yi0/k3Z6DUfaF+B9Qp
Q8Qhd9FyhOA7wIsH5UPFEE/lKvLzDLgkgZ4UOagRvQbVDM0n/7v3Ugg8oQA7imCH
xS1S1up2Z1pPADNXev8Xwuyw9ICQrB5gqoRUKQr1VnTZ7O491Qe9iXyFH53kQVL8
1wT7Yz2LcX2Un1u3j1Jl7Kz6nC8bRir5xwXDI5E91pi0RIsjwbT99DtKaxrgkeNe
dLF1y3Pi0OdkGKKtC5P4VqyjBOqqhV+TjPFrmaQSn1rXgatqdITrU9u5/cL/+k13
7v5sSDatrHkHIx2C169MGuVCAw1W3fdEOTgPuqxH1ws/HWhMKpl+LC0OWK8VtDLH
qnG8a8T4z0MezmNUsvAkjONL77b5iT9+rmvnQCkDwmgkykwGlUNdekMkNArwcV2/
WXOXbHy9K1oxazhVQr6+gMVTYdtUnzsxEV4GKa6Tii4qJo0C+tt2jrXia2HyCb3k
bQROn4ZEsAH50CxwJDCQdwxviu+VSMm+50pPVIAfOtDtFn/1AOA2e3/hpRcl6cBF
JkqTJ2SRHZNSXQLosXNKDEuIAZ1PssA52Kpj7GzgqnDyPMSy0b0NT6nHtJcdgKtw
8EIPWugyECK8bqUOEmWJb8aSGsb6Fet0PnIyLTSlLp0z7+TsHW3ktSmc2NypLoBI
knyEWv43HDDdRVAIbTxvY+T0C12SZQn6Vlcx9+JXQ5cSObKxr6vRIbpjF/KqrCae
YgKNM+9H0aB2CTm9J6E4X618DbXhRX8/SObx3Y7kF5zAQvUjxRB/sEhkFP8lGTZk
n8Q54dcA7NUA4yUrhPAdJUFq2L5Pfx+3DkHTJau8lasRF6DYI36kM6CxNmMBzUk2
HdcGop24ga7F5NkBHPLmh2kYULUXwKp45UUW4euMjc8lzPhjuqeat0lugrJ5PzQY
+TEdUAq/CaWcqlbDWDxpqXAdSRDB6p/Vte1CJXpPBkOvJpnPAoO5E0I7BbIkKmYw
Wx8D8Bs+g5akINLBTxMB6DXrPtrXLy0Dxk3n5M87iensNdQR8hlEZmFsvzmkrXh6
ZXzKfQdQXAb+Wi4oHMMcPGgPBtcD+Cclwr844lffVl0Cg5sKy8iuOpNb4C3GpPFr
5YPD27vDJWy872BUjOYSPq+chziebp5dFBLbNp9tWMP/qqaTiwQI7fJBiYlLMXGP
ATR8Ov6WQwaGjgaK2KTc7lW0QQbHL+LhjLsn2a9T8TtnnModhoeCgRaIKakHwRL/
fI37v1NAA6ZY+pqopJDQLhW/MmrpAUcB+/NPlRMA8ynx0x3MzFPqhcR3oNDuKaD7
Z0T0Unc6VjQTLJa2cEKS+A5Mp8QtV2HkWqyojn9xAgqiSEnVl1rJEnr6S7E03/4u
LIUSrqfZJNfNGQQgBnhrqGCOO6UAXYvS5h0iJIu8Z2QnLl7Y5eVWwYcYvMz4tvfr
B+h36hdsxqId/HvdQ+bmle4VX/b+F0ijznZAIK8FnwpOv9Mg2Q69dzlzsFLywoVT
w3TREY4fAKfnF/ztdinLwwP9bCNOpC1eCVT4XoGIPzcIvy3XSAk2hBkAIulQd2/X
XeNdF6V3DwPFlWb5guNTcVJi4TWqHo4T81pf3KYRg+aAOonTKtHg9DXOSCB0+Icm
2GOZ7T18pTiBZmYU57CUGPx4lH97GKyRHX+J2eJEXviiAEE2JVeIR9sAmXfyRRq3
SzpVvXhdTNisQ9jTAjB3AvH15/7Ytk1z6UKrOvm0txPcgQqqIpnrirW2QvmTXgO4
pHIBzPOGr2TiF6BL+nT1tN8cijsxSJNj8IsaYzMSWTGZQUZKYZoG6B4F7ah+Hvrj
Rm0oFFTSV+trmyijo9reHgAKcCkygOreJZ/6bmYWLK4hpYR0QUBL8tqwQxmiWIxd
wksf5rBKqQ04bSjPwecP6Mq2ev6ozxXQTi69ERaj9ZHoHiELi/G1qCQ7NaPoSvRS
+GBjO65alMCd60A4cavj7xPpc0VuGVXUqVQpItGUP7ISalD/LS4UgVn2hVCxsesd
ap/ovApgaPeTl32dZfljzJxzEi74Qvrtq3USqxCEMJ69/0JgHvI0EoqR54cZOfnk
fQ+a4HitQvv/r06BW2jCSzFSfs3o2asm1j4fesKgneYEuq7abxWW4Q3GW1QpUIw9
gEiTjWNqAz8CNKqYArUago+nsVHgWbPvXi5/cyXvbUVqjVx+ihhoyGzBQuWmINdi
42E68MddBEOiT+I1QCgnmUzDWFmr/MuwSW2chx4iD9gWWEm2OZB6zKHEIX25aR1B
WjwcmF4t9xuQWzrM3EYVRD2Mb/+8nYftKjMfXGI7BKvJVlXBoFe+KucXYeZBAmv8
lIWIXQKApxkAkldtJD4Ru/D5bD3AiTt2bZg9W5k4jsVhWQjRm0fY1N+BBi0ZxZNT
1Gri9cJOwt7eKzsaMFamNsps19AcNM3VyQQirEPQR5rhucrjCzg4cEfxofHN8Q+k
ZI5HJPAXhdJFyih04dZ2Gd7I9jx4H1Uy07WBw4T7wBombqoJGOogzYQ0+kJDFUSn
1tx3MiAIgxQygTBj2Uu8sA+XqxMnqDH4XcTtt6aL6RIK1dLvTUoD8GkcDeSib/q5
6ZTM3kOUleOmvFn/GIVMjLZj+zimW+JaJiMHZDwf3i2IrG1INWJNedXSS99D/mPM
vAklx3uPyM7cT/63IbEIiJTP6daD50du+dzZMbVvfcDAHH0qinQORhbfSsdLlVbc
NbM366jXARf+o/5hg3xeQ9erAkHFmrohU4MdIQJV0uhK7LuPso5eZOc8faKH9MIL
8oy0ocyIWcmHEIyu61NbnIxUsErvb2XArVVVNK3zUCoFwZBhlf5h6G5Qzbio/jea
BLIlWRZd5UzX/x76W/HwF7XadnMBzcmT4GEd6OviInuG+dj0BfYr1LvPKugx2gum
eX/eePxJHOiFENi2bpzTNK2KnsPk9o5dbf08aOe8GTgLa25BkFJ3hsD38ByUIAP0
QTVLsxsJ3sEVN3pwckVhd8C1cvUib8HwEay04nwVy8lIRKgKbkCrtnUdI72xnxWO
XqevrotBNIWyhGGgO4K9jESFTiYvd6uKM0gDnyHbVWHiV7csik0pts+rTkl+TgAX
BA9M/T4L5c9tVoXdxWF4F+StnkJVT4FIXg7e+h5wO+VLyB5DgX9/vZO5XITrAWp0
khrXxKQjDsKuWGE3hd+VIdHvV3uovQH1JN4VN4b9+THUJyMrMusOHKPXQ6m3LFQf
Bn1Q79qA1/GWTlcOmWsLYbX6Ry5Ajg4gpWuFBDvByHCDbUz7R/ALmIoR4Wpsrw9+
KLFN8AnOrzT7UPU2dVAw75VUffLvzwHTxTODBdSeG01tZOYB1E9ThzqnZPJ+V2QK
UyKuzxvhqXXGU7K7Qwv+1AQRSpRLA7Cs4yNUd8gSkW0YGSrPmFFzqwJGY2QINugC
cu1y0X1lS5QT5+x2M3BLUHxkzyDz6qvcZAL2ieaUoHpriqCzkxG0xBds7M9lemmf
SpVHTVRP5IAsrPwedPlfLrgmrAFopfPVAk/Dv/g42Vm5Kz7kQJ66ot0EPiYaDA26
ef8p8dXyFRdGu2NZdopR2W7AR+WCEhZaEFkVVKNWPKtJVktsF/va0TiCtEEuQtTi
TRNFaPl8wkBaf6DXW07AhvSuvnN+tI7GC9dsjcUoZEDEFMFpsRDoPA5Mo790smvq
Qr0+bC1/9tV2e4hE23OTp/hhhv5t1fqGSndHnLxW2qkvaGzxyGwGdCuSQW30S7aB
vKRTIPhQM4KYsX5EWjgX4s1F5Bzm/yrrp4OriM/AsqtPj3Y+cp396vBYEkzOR34t
gDyDaC5vlNaSxZHj5ry55A0FwuCa+wJw4Zo/ZHc9fmwnNu89hxfovvg7x9MR+Nbn
u8owTOw03QyaW4P021ZtVoGV62X3QfPYUYVMyyHASdIOcN9fLZRnHBQX0YnFtqJk
r2U5GUbfrx8X1okh1DSDT9tJ3bn0rUQh2sIV7waZz6CIdsLFis+9yMBh5/cCuPP9
DphnyzOPchB/N2KdS6A0RQQcGu7ebA9qCJypg7n9EjomojRuzMeo6sHGyITAu+v4
TXRdhmGhZTw5wlOdXOvwbqylZp5MtdaVCYEo9EaXIS7Bbhc5gmHOwvS4QwxuEl76
zagXFWCm8EbYx78jzMhd8x7PJiP43Eqfvg18LwIZ+gbwKdd7S385L1Sw16SQ1eAd
gqxUqELOzv0f4VUpmhPrHz84m0goKMYbyBOdxCQlHzo2Pv5X5M6XyB0QFzN5fyRm
zgR7qk8DikmEEaFesU27H7qfUX5innNPsgyVTPpc4lBB6O8MBT4Y6JlAP7Pej5Ep
4VZPwxjsZcS8gj3dCqwXXqXX3CODYRt/OjRKupaGjOmbT8h4GWiZBEQGId3XFjlw
LHaht6VkHo8L1Kh1n/5gn6FO+mfAqORtxdxk9fkcvGmv8ZXzPkdVr/zpjj01ijHk
9S0NvI94rI2ueYoj+LUs8hIGW5NRmpJZlwZf8Leh9dtBtHJkDmJgZ6LQ3Zk6MRAO
QM0zxZzy5nOKP0noBDuNQltiIQ91yM3ZzHhXxiKzm9jj0HbfsrS02vQRnPk3dRFh
JbpyqTiFzN0wJbPpq4zAsOjOLgwHvWq4IsAvdd5TXORnvJneAPjYH2MD7VqyQdPj
lH8hD2DZbWGdQUTTO50nkPeiCdSeliE0PGS2zHcSGRnSJz1MHp2mRpH2gXgwmsEE
drr6EqiJ8Pwg29I64P172zVq/xQpyz6N4t+daSy2yQuAlRbTIvBvo+CKnLXlrOqK
KnPnBiFk2Kp5ljrk/mMFJoCgfaWvc39JNTpHq7aY1ErkpjOZSJus0kdNoDlIQ0Vx
Pvy5jFFTLM9pz/sp1pHay11uzx7xaRZwL7sCEEfNg7MtA+3ZXhaFnMnvZAta0y6E
pNllcSjrKHHYfN3W3ZWj3Wxl2nvmZLrNjF0DSnY1TqZLk/sRRlNEaqZFsTbj+4sQ
JIkaTgemJYsSDDWhKq1AvAkg074OF3VT7r8ae+AEfChWPTauM9GrUTPG9QETAP2C
FvwMRxn+MrTusDB28WLhkpfAfY/3zCCgzidl0KNt2sM0yAApbiUdvcxVxqiLRxAw
i44KZfeulRiTr+f1N7yMZxrwv8XwbA7PMgwcZJ4VDYWIyWKF2xJ5lfRAvZlPwmaV
YNKtSgpr7EE53gZVX4EpcodIt0LH0bUa0H0Xj0DVK2moMa9dieGOVVgoD2J2rmTm
e3M8Lt25XKVQY269jdH1cMmyac6xEVECfe10SercKvuMyM11Dfbhim/q1PC5gGTg
pGhmheXzwnpUDseq/64SrnsRdWrb6t1clD58mg/Ky0xyshc3XKQ+v1LVXwsJZPip
Gvlcsck9m4LJtHg5TK1SEuwbQW8zmM+s4Lf5qZpxC7Qvz7QSGuhpjdEW589m8To/
Y06/NeFRLZCef+1SDKmWX/jxz6neNSyOC4PsFLD7SJ2rB+aJczgr8/awMUUi0z4O
6hIZcAspaWyIejMsLp3BXYqNLOjIGD32+PTzJpA2X1egmGnq8xpGCLDqWErZRUMc
sXjiqURTRIlBHcmQM9sH5dKNhTc1FFz6o7u9PLrlGDS13wprpnn6BGqsFr3HOawc
jRIlX0GlWOA61qwa7zlfUzfPFhu6vEaZ1b1/fy8Dur8ZD4wsq7NFUK40oP2hNT+i
iGfRvgQ9q3PnrJhRhXq/JHLI8x+BXKutmnP5T3SiL3eMPUZd3UtZZbMnLN8rMQQK
rPxFFQL2ehP/RA6xrix+wulF3uBQtThELNCBcUg0jPMexHIwayq8D21Yc8KW+Z7I
Pf25i14Vl6MVqA5xLq0pMile8b702d7rfG+PSkJXsqicsD/v87hLbHZphvJ7kgDD
Dvze9IuyFDuXXPO84cRULAqaUVGXswIYFrbCdOlU3h14Makbi7luvE2zvv3c3CNP
IDtgolDlfP+SGYSC5sQembMbcosBEcWjRDzaC8dq6DTOtJB0rrNEDMdmP4d4Y10B
htpcoVsCNyngY614Ghh0W8fmJvN6vmAwBLwteMEhQmGs826mDX6/X8viHBehQMR2
ZlTPEoieWK0ES+2A2IzcqrOtDf4IlBF418XxOJwfJrDAtEIbTXJ4hm4wXgM5nZCA
sqpM/4diJi1eae3FThRWfdWHRN6NoVczTspkEGZ5l5Ysi7Jh5YXDz6Ed9B6nEWcy
KqXDiMI4DizKdr/ms2kQBasjglGvCw0coW3Rp9OtUbxsq+I9DEUkklN8yVvGXem/
4b6dZrInq7i6eVkojEmC5o0/vc8ThFCBcS9MRd9fOnLWH61VSxnByJD1zUUYiRg4
i1QzjdEdSc+umlyee0t4uE6e+4cZD5tYihqJQosD1P45elPTFOU/Q6gVwIURzwsb
LjxVl8cEiSaGGmJlbxkV7dCIYguWHeszXJ/15RTww6ps/yRLUwFsLRdhc/zCMPMK
nlno+InG45CBqBSjl9kmYsfU5QMpB5+ubgtdX+lbft39VH2zJb8nFVKsWLsTKq3q
Pjxll6hcgpMzAI93R4OmY9BYyWU4se1L9J894grxOmwTED2sLydlGbK7UokACgr8
VhnhG9Nz2qOCorSheeizg28nm+fbK8jy70O/BQv4ugNqdjsGuQhnQptorZePqd7h
YcVsI+B5c00oLbW6uVPF9OFBIQDDlfk9+A6AD6ypuGffVHiW0L/trqAMQgnBE9oR
T1/ADsK4KXnW2UOf92oDYFpTcCn03i0bvLcmNqtDamLay3coGruICCjvRhYifO9z
Arn9JJOXnKhDb/UvQyb+03ekKaXMcTyWdYtS9MDKaPqi5CWAg5giQsntEEBsPZ3C
HcumVH1tC6JXTamwgOFztYf22VAe/uok2wUhBmpdr43QGiYPgpHuI0RAkQRXG2fb
3g3hvKY3Bgectkbi5VYOCw5MAtzL3q5RS34JwoWyLSINlb1C2p85ETH9bMqie2Nm
137Dt1qRRNx8DjPzwEbkmK5LRCMv7hckIp0IMY73Ne34svMSMqe0KB7IjVkY2nbN
YkbfFbXrQod/HEwdP8iC+eIH7FXRRI9BkiESIPW2iF92TTZy+K+b5NnCDQQeUQOX
/3ti4o51f2R33ubV09Shc95hHmH90G+Ny21FD0z+Zh3uVjbIXPEYJ4zgg97u6eTJ
Rf9yiggj1NhHU4Lxe+qep1NiS67pc+sMkFSJMYU3DinGQLVSubOkqRVyjJlYU9uS
fEq6RlaUl7Jzx60S3pSjVz+42xswNdYX9QHZ7h+Rl6n/BUcs7vrdy8astBhj1pD3
7eMkw3w876JYtM8uoYSa/mG33UiFdwokwq0agZlW31i2UUK14h8OsYeh/5pC01Y1
EplY/H7iu1niAUgdBRKfDx85twYK9kcVzRIT+Xv8QBcGddpjyVyUdbFJYWSLAF5e
jv7RSUGkBTVCmST6t+CWyypMPV68gpmKbXJQbmAJq4Yr4zxRW928igy9kRsrLdae
M1DG0suCsKAJonDjGX2oMTAwBVn9nThtMb1TjUBAhUEZ7Gpdly9UbLp/GTJV9bbt
OLmIe3df813rExsFvjev1n9sQc6XT6vMNXHffv2A2wzu3EMX5kJHRKk+vMNH1YI0
YQJcNcFIOX3+T6Ke6WoH6MVksyV/BtqfBFx0jNYkb/XfFO+nRKToK0eCXLh35k8i
Ki05lizpeOblABL1hEDKPdCPB8FR5q4l+pi+FLotfI/aAWEcIpijJUcAiUFhzSf4
m7uaQbDmESCPVtiWIxy5JXXBtshDMya0jP6SFPRA/Lwoj/F1+gP/q5XfMFpzvsan
ZnsLXTRU8O/fWTtcgACATl3q7wOAJeag5dLSor6eg39v1uSLKTTdl1RuPMvQyajY
F++l2BqoeYzBvBpB8JNnkrcsh1ctN7IbDufbKE4D+ze+RdMmefgBsKGSZSGyFjlV
933BiNKuarXqHceDfjOzMcG/OomSER9VhCutSqhFAJqwb4b4e8LeqbtvELMVJWPA
2kYiSIlZB7AYWA6Jsf8QGPK/ies/OiH4MuLfoSE9/pwBkv+fvgMCagLG9THaSLVw
ZtjlFlm0xM0WZsLDR0JEisYahKkKFl0CjkzKzv2LTu7vuyZDs4tY/3gq7//GXLLg
daMCsMWlkjT/x7lc/3/lXpYW2xgCS+kKPBajruARQoKHWzWUTr7QsGc/fZHF4fMw
krJIw3nntaSi7vezAJIWR6sDf5FBRPFusooxaV10PyJf2zrHykoI8QjqCi5Bks8w
aVYRNFaF/eY9ENG7223QsIWr3wRQjgINuHv3WcoN5AlGHznmFTafj3lfoo15fcSc
yXU+A5pnZzV6B9dqusy1QYEka/Fzngi910+vohZBHRbWJJfzPd2IdYjFe5WeMn3w
Tb+auLXcsMH76HqnCV8t8PzGWQBsSrV6uyj/Y1kfcdqn+vDpXxqIzc/oe4efdb66
2n4Jf8CcxJRO8yPmY4ERwHLyQYbALDMR3r6SxOLqGqeG+vasduoSH7n5U5PVXwoq
U7xBf0I6z7aDBU2rSuNKkdczpvFQ4qPxOxLH5OtQSiudhG9ECabbyILPrcoJAaKy
TLSAOTUYYnr7Jb6nPnVC57svC/CkWnyCWIprkMsqXHrxiJje6O0b6tyK4r1HeMkb
yLwrXt848ztyJraFAZwWGt6teQ9/+VGuEp1sNUZLtila1LXZeuvooFjwY1cgllmN
0YmYYNLbjgkxX/XWqyL/IvSgKRvyoWfyKj7Jvr1/bi2Te08MFPSaVxsrrEKGJGHN
YLIVY/QP+1h/L37zal4ebF3qJlK677BxK9dmXJKB5WrK+DOOuCSTq3g22jNmXyMy
vzNOZkdrolLJBBGlPxs+eRkFTU0hgGtwR3VYT85hN8w0KJWhAIsWuXAizu+5RcT9
PtO/5UKJ+qPf7nwe/lZRon9TtThaF0WvW9iPoeBl1ZuGqbwM3YUt/z/bFgZjjYFX
fC8ngn/5DVQxk07+L7K8rYmtwTZGoxs8tO2iYtsonLiW/w9sdZwrhfBUGa8Al+tb
os6c/1njiCSd6cfYU3TG3UUWCGKQZQcbhfFb/NRedDUPYlQvYlujX73r2TDfQYCj
fPHf9xPwo+dcA1/sf7ls/WIWQWGntDdcPwJhPoarYKP1XRjC81rL5A4E5mb/GRtg
3O2zm7kNfGb6hHbrhGF91yAnN9cDudVqGra9jCf0eFjuOROxZ+n6uXD83GQFnXsh
6BKfav9Mzt6tD6HgGQEGCSTm0xBjvdowa3vaIrSKpXNERnKQbJd7d8Zw5I0/oRjK
wGUj/AUVHN+jZXQ0H7/mT3x/833+9+oPBFqfpHHb6BSUC6+VlyDhqdKRP5cLnF1b
oOjFD1OIaKnM+P6iZjlaBgxJWIuAPvZEMdXxsA3MniAb0bBJj0+b2YqJhsmH3eQ6
AkIRyjQ5j09cpQ6fbgHkg35Grc/VXf9rmrrCq89za5G1RRPc2pmtMb49UTLA90iA
SnNaCOWMFN0ayhmQC6v9uWjIjBjyZtBpSNXWLvA/R9IAfZ4uabyi7ON2tXnkL8/9
GeXjrdSCqUQfQgWSKXXm+9LanUe30f2ASc+b9OgqXb0j7qcnlm3/d+xRfsxs56Qk
bSraypSnix9tf49M25vqHzjptTGU8exLWymvp2byJfnmLIk8VZMRl/7J/6Uby8lp
p2ZvDWztRe6a2hmCe86oxE7XVZM4X0fUyChB9jP4YVh8X6MrkMBamOzoztNvz+dY
4Clrb81C0mc2SQV83Uktr9Gs4QmZWsodReDdWSFN0V8WDFyWPkepqblUY9WvlyQf
6Qxp5+/Zy2pPBpYGVPcH7ClTr2SilnOX05dYa6KrAt5t0HXvzT8SSfqGkfX9vC5z
EO3xHbAFjbqDvAXMairhf2mLgGOqDkPqccHE0TniOMpmGxo8ccPcCOKB8r97U208
4ddlviy5wYFXmV1w2El7hXDuOLi5gP44RBlL/nIOlOcx5o/C70LWyyQGps4w1yVn
Ijxkv8Ow2zLCTWgz+BNE4VOJgy+tIp+kss/6OvWgthAXiab80byslbA/3GNwbXQE
dDhbrZCv1R2g/hg2Wf0Y6fKtnOZZo8XCjTsIkjLUbTA6hW5G5TvPgS+scA/KNTmg
nz4tDRksJRube5yyD1jqGLSnYEznSEdWU92wS6CIiopopUhauRoP3ivhmR/RWnyn
tmHVf6BkD29RPJbuOwiVoODSyckVk+S6mzxM0QF70CEz+Q+htIHZceU8vC58QaMw
Pj3AKdzjR9k4SgwjGjlRb1RNTeAgfjhapHAc5n2nAUl9zas8QX00pagc+FLFPT8/
aNUx9vRXzrmCho+oF2ochSx5/wx7X5fzT1hgTzFIEB9i9SvfpQBIeh4gbxySoz7I
uGXf8YW9a/J9w9n7hThdIPTAmO2dmwPcpHXOj+1PgZOvZqiEn3YNoKfLy+WSw8RJ
G2UUL1lCQg+ckRIdpIIiOcbgIGYAbVegvwhzT7wywyRYcqREDSTExh73gg1urI1G
XK8crNWPSxkhIBG71l+F0x+3dN9+j88OJ3jhgdVjaR9kOUprR7+QTcFDLP14uyen
9otYJK/yQOqXXbjZgEBenQFwbFGp4+ixvRvSXir/UG3qg43neJZ6O7db+iv22Ync
EzHMZtzp1y+qdokxBBDnXYHSuit2+ynrR4/0BOb7pBbfyl+gzTNyW8JqKNvvnKzC
lySS0K/sCkxEEXgujKsxxevgTK76mf3lCgal6r23jJ/vjrCHuEkHY3c3ZhwiWpsT
Yb8ZCtkgcYn9SM6b7HvtjeH/jmShNHAYCKualn2btv6wpyri20du788yh3PeeD5v
bmwT2/nYTCiAbmsSQIGd/GSnIQHg5wV0l3re/N5jtdgJcqcrvhOJtsw/ZiYFsvfX
8WocRJRrrpRGFpLNdNfOTBdlWDG4Mqa6MKbkZTGxhKne3/UbJMlyVTKWvhGxkXal
33yVBGHWZdLPisaJwe35SKT8St4YItQN+UsJGi3gAXSRB3uiZnhxN42b+7ZtJI5q
az9WZCGv2L2ctutgK3SaLCRFCYQLA1+Q9WWVtLNvpMS0fBNzOjIZh/ftag8LdbYZ
oAFtUYcQ69SqH2bJM0kKAlQh9Ow2eul3xSnLZQmocgoFjcbjEID9CHxxa8ovAPFt
A7NLXN5Ctlo4g5aW14kcnqqccBu7QDFUNkbXoKsp3QUq5hcEYbwTLdw9v6+lzn1P
VlGwOHrZ0xPiIM7JKP8EEW81FC2FrI/Y44vUef1a8FDeWBYmKr/28QQtEt6rT0rj
qAuazAHP6303qWC2eXu9KPHB81iNNFyZ1rZIYG0AnPehOmKPeeBcgt2P9nLFNYb5
i6IpZdk2D9ipUbRzJVoyb/MkYPqFZYTIeM29TPLNUn8pslOr/UPzoJI0VVlRTRIu
EpvQjou4y1n0V67aKnE6oWU0B9u0W3vB2nB/zIXBqxqoiRp9uUwNObCVNdzqCYiH
9mgi0g1Z6EuU0GL+rRnFQtccyZ62H2GPngjoMM0/qq4iQ9TWZeXxys58ZJ+Gxnco
4VupJzvyokd6m4dnYcByUfn2qODvSU9RZcUP/zSjlzzEaShZusoEGy1kCOwWLMGp
GLneZ3Nd7J2ZzmXstpB/e7gpzTg6vksYEED0LC4hDE97ZXb1d+sUb5W79OS4HVFz
Ax0qtFa4/rLZ01vL5Z90ya6upNkq4a+la7QOMN7jIPeqRa3hamsdF7IeLi2IVEee
C1tb6eN8atAFex2MIOrBu9koqNEG1cE4P7Cj9oE5QpguQpSbRUp398jfxBKBKqK/
w1tl7VEy04M5B2sFmpMtnzSLU/g0qrUz5wW+yvCXqncPlxcas33shO/W8kUOy5/8
vWdiLvuxCiOEWCXoV0nYr1nJTXSv/O7R2zTSSdBeBZ06xhnd5nJMrhGul85oaIZn
8kJ3FiOgN9G/ui/EfpFqPKKkRKVa8lAt/6pxUJQa1DgZI48VLST4n0/C74gsx82P
Y/TYJNtJmDphydNVHbdQjCoAgg8Vb9iJrcLgrepIzxOLvJPJBpPkWby1yKIyYBP3
FgvH7p27h/DxpBOzn001jAl/e1+L7kaeS73AE+z3BEm9d74wSztg/9RVsmmI1lsw
PMD+8AWtcv3q5db4wYfAZggVAlbzTv68tZRnmmhFIR0DgVZNHVIwyYvwicDXZyLJ
yLdTYAYt6pCqAZF6VKnlcQTYex9eUbrXyFeJPElyiwZemA+EDT2Awhql2VmSFT8t
0QRWOZNSboozgzn/E1OF8U0fJXBPpDr66qVK0wcPbxClw4O944e0ABYv1gJQPw2/
xhrmp0BYJ0QD9NEmFeVu4O9l5kKL1DG2plVFlOKqYXvBcoAr63D/eXJ+jFC2SmRM
G4erRjYu31MNMUH68QfXHcEccBVoeRsqDtlS8cf53gCec5qqIoZqLOqIA5xGLZjZ
QzTvfK+RFZZ1P2+RUgwEAR+swdLvUIbXe7ENnSebLxRzHSkbxDg6SwOyPSmnPb8r
gPS1xh62Fnjomzm+d0AbnnX9vy4SGtL4uUuT+9EKDQteIkseAyh4xoVhxWJpp3Z5
UaguEtqgowgOsJUkp8FSKHa4jkglSqW8fqHyNp2wteYrfRPok3g6Ph7njQS8Toi9
QPfw+nAKiAWHomHXtmGc8l5Smxvzi7vvaQZkcDZwbWO3Nz4VwtW8WT615nbYa/bL
Xu4HQ+HDuE6mMclemVqKf1zgqcEer97792bQIBxTutHbB0XWfHxnpUoyvhChkOVy
SeyF6srfxqCFNn5iZyMW9FSkdHlz+B4hvT75uSHFcutRu+xIxxeIE6pkDS9bGapf
vO39VuJVVGEYwY1kLuM1Ewt7qgcYkqlVaOImN51dKLnCxw7C66Uta4X9nnjiLYDP
6lOIzUEJlXEDWnoJDoaZgkhGrqiZB0Cv2VBo21yl3tTWYlsucNuRvNP6v8l0n9nx
vMXpecvZw9MTFIx5GgFuzDl8J43ju3rjskkexxoB6C9jSo0CZXaF/qTaJc4pTFoS
nDv2aUgP8TWc4v8Bmls6Oz+tyzqCW4ZExWl6n+xUbdzFAZu9fnxjr0q5qxKI4clb
GDD+KsakqE6l0VuEI0oAF1SIRU1w+rEtiLrXgTxhn/IE0VT8G1VI14SfjnbYZrpd
8MvJdyrUgs76/P17wjQFX3yI123GY//nLqLDRRrQe0CiNHmR0xHltYTVvKwyDj6j
eJ5XZDtqmgz2gzeGrDrU+BX1D7M5SG5aVWzUS/9CZuTWkyF9kit/F8+pVzZxAqIM
Re5XTy8TV2ryk1q3H70sI0ugZuFPaPQYNsh+JawsaC5bSTp0IfIBUcAEJOeV1uQw
LbmGcbSEiJtsYBy1rp+HfnxH3SayHzTGF3k41EVUi7ekkTpILi9+EZB99Hitzqwp
Y/F1GpDRsOa09DPKiD0u1fP7xhBPG9CAIX7HpZa8y7rljB0N9SNZQuNlZ6Dlc9NL
/zMyWASdN1lNQ6gyS67G+Ks2KOsZVxx3ESbGV+sZAf42zYFuVSLUCeG2qOO018+X
gkaCr1QCForpZ4+ZG7OmJU7dF0jCSQ2Vi3C46+KIOpjyhUIOn67wm/LqpT6rGN7H
5qgY5KNhGg/LOLhSpbwrfT2uyKYmXmK1k5c4bY3DKIbCaxNY8FGDFYEuR+Mmnqz5
U7uTvK1jtG28o6YYVdz14j93bEcGFYjfinqGXkABJezlMBxShX+P5lXKQ9poNJvd
2s9reZ5krhAXkHb0VsQIL3fyGGW6wSDsUHtW71QN9xFWed4vmoJilcw8aR3uETpY
6e+nUs+FcUTb/MK/1v6dBhXa7K9TXpCFKIeZzsqDNgzCoUFd2cufwYz8Oz9BFrQC
Ai//hpGKxBBE5pYUGmRkOv/+CrdivQUrKHP8SNHj3xFxhHhsy9qetgzkGvKSDGi3
Z2I9LY9DI2nM3q4ysp+AkQsa9QVU7Um82VCHtsMh23BseB6RfjuhWakw5KpH1nK8
HHDmHsUci8ZaJhFYgcsX08EQSlRJnCjqtAHt25tlYuT/jF6ebUCqVkIQOomqmzuu
DPPHcbiElHUuTDlZJWXWlw9miEOtqhVAWmwTneEq0Ym4W04YHs4dV1/yKTl2k3y0
/Y2vgyKLoUcINQysfoxzSOILCTYOM6EZebcv+XzxppD7KzBm1MF+2ssguKxTrnQ2
gPrBNxhPG4CHdlztkWVBoIZ3DwwD0JQ2SaXbZecPJFPZtH35QTeHCQtjTWTMKgnf
GyVEOkQlo6vJtQ3SWVmSmYNbRchAT6w/CywQpLAPmAK+QcRwRl6xly5l7727omT+
ELLMvHgiaFJdMfpdGK5FuIGjklEdSKCEMdwsDvmwd6DCBRP/QaOT8/P6SsRt0GW3
BujijVWiGc4QWn1upK8ie74EfzJ5676T+zfYDQL0RJ/wqwLGMwxcGu1ZXznGQ58i
kC0loMhaVr9afihayS0ALeaxRFfgIYdkNSpEpaOCRJzAIql0tSF8TzxKFZWwFC6L
LbXYI9c7X3j8K1ykVhKOndxNGP4HaLGJlt1ITkt+Q2w4HFaEltf/RUC91iHSAIHL
Wct9F4RdsHNWAr2QcPm0seWpBJ7nW8RoTo9H1cCsmvtvg2/oFQUKW8Bpr2XFWHEa
ABP5Py2FyFmKiLsb2+NBdK3P5ElAKqwnrbEyQZWLs+ah/2bor7ql5eEs8SCf63w0
tzfH1UUA+2PyXrk2Iga7u0sj7H+bv2ooZENo+CvzBv/K6PRCA73vIaq8v2xLPeqJ
toDmSr3SVSmef5bARhah4JmC4U5NbJL7xtHdfo47A+3b6Ot5H4Xbj3WE1AUkF3Vb
IPvc7GEIocIP8GIdA8cRkq4na3RjQfHw2fakAL32+rQvIjQ16z+aJhy3XA+KLWTU
tmvNTU5t7iewu0L03VQuW3FTo/V5jYo4ZAbDeD39h3agIAkGp1qfkVMJaKw4XHte
1NTh+PBO1Wj8LBNL6zS0/gOa49M1EhuOKXPrs1tgxMthpXODWMR6H4Bz3QjWBMUD
NGzJcDamQLoJFgUt5au29Zpb3VBay4djAegJyHLngYYE1C9B0p+OZDzy0X9zBqkZ
ab6/lllYn8wW+y4G8Rm8nowWnA0vpasUUJy+dEwfthZPV5Skca7E/o3IuIRQeUBo
udyCqWx/ha8P5+z7vRyf9BS1JDqBswG7J+N4J1vDfxC2+toAemxfT1MREIgSwkdU
eJhQ7nhig0FSWD4TM9XTWToP93BPasAorp0E2Ea4e5JrPdkfPj8OePNBUtddKx2c
mmUHqODg2h1Vp2JsFViDspcZt2Yvi2/iA6IuYhCT6c5oaiwX89Rxoqm7IbfzDNSk
OsylA7rlN/GtAxOZLFnWJZzU7/PPf2bEscchZWOV9FJnlenE7Dkg2bEzrWsWFXYi
YtsG+049MhWQz7+UNu/JuQpOSHji/JOG3cCVYyVMPDNj5ij1+o6sIDzAnZ97lu1P
z3PejSCjeoAts/fYKQLSTDZYjMgxJkd1LtkPpcnAmPoFwdJvpIzw0ltt1aP/Safo
TUCgugQoqT1tfxZ+bf6JYDl5elpspnVzvCYC10vbMolq7sfMMeUds2qwQVCAPaDP
5PSPQKad+igFpWndJ/IzuicpNTlti2xHH6SlkOrQ/D213xS8UWRChh0+VrWRm1Aw
3uaTbePwIYc0tFblvnyo+R6gpUzKwjiRu/ya/liydQTV17TuyY6oYc2uijtTWvzT
yrkBXzJTdtaMxdoPF1JMQwB6TkE7XnBzHLBantVLZM9TygmdM6BK36jNp/pe3XN1
D29oPe0InCtty9L4NDPFpeqGNbGcXAejbRJQxf0S4bPmWcuAmWRRcUcCv/LVAOU0
qttsm8c/ZORtV+ApD/2LqJCxZ3Y8uZkA1ntq0HFwydLa7hnX7PgbIrsnldKys9Un
euF0U5A5oxOhRpA+CvAuZTSC+eV0Hxht4rYgf+BySHxTkUHFWi5xQdc3/PrlXK9s
rNauQfVPXXv1HICQJW/gPWc2DMBaV+p8EUKBLbzZ+Wo0RkCJdy/fLphC5huKHjlj
jQ3xvevBfRm0a1n85lQYLgXMMky8tt12xP86eB53eVUHCSKQCcXOXfhHdTJEMNBY
IpSbyCrc51u4m636j8VxGUyTIrZr3V3zsKVo3D7Jkpi6qFtYUBdDNCpo4NxX6fOw
AuYgj1om2ZIS7ZQAzMZMkCiYZlz0qY7MMnDb/4hOjACsR1xzxhnwZ96+cT37fHsa
BpFmJoo1f2uGi+jDLz3CBmAAruLvHZZujWwENlp6YgR7JbnXw6Nc/mhMnpMDR6+8
RU68XWiLPSyfozRNBcwdycQBvReCw40qYPL3RYeCBrWs4vjQWogUlRb0VVBjFtgB
AkqotpE8b2Uwry/S64fID/LoLhXBnCe4NTVaQqkdcZY487UB3aSG1EojYLsuDoTu
G9MmCT2F59nxKOATw10Qwa1YmO9dZYu5QI6+DHFhz5P/uQk0MJ2JbsZbwvOg/UwU
c2gBdpH5GBvrZxHLQ6oAHB5Mq1tZG+NfXByzdlxUmcPvw/Yv7wYEn/2YYnV1wTyd
oZKbd0Q4VaKLBvg47MLUhNBnJAeEwAX+xYPLf0kLiqnENtqEv/BWk7q7PJSXDC43
n7ioYah9o/g56MxFkvLn9CG65VvGHQYLsi75cd39PTkGO+muw9z7NT6DQhz1SdSV
O7046neCtUaFL8IhwgFIpB0j6PfDcqcO0jkbsaGps//A9r24R4RnfDTxio3LtTdf
WnuTX1kOMt7IMwfIH2yMZVa3Ja7JfXHC3vlhQ/HkijCfPWbhviDvMvRDT2vou5sF
UaFhgLoTZXHl0Owfcl39DlWWeyZXmWbBwehcegCdOIoxW2zKqKX0SqfHKQdQd59Q
lwKwHPOuEbod67ANMmsQPAgjyLbdRAnYrce4bXWo4hv1W6fyQlVauFcZMI0MrAZN
3sygY2Xc0/9n1ltyzZj9FBw2EgfF29piQZi7EaBSDolntRW+p2y3k3wSdXkuQRmu
0r3LSNKrKz+LjKljzLz6odPim9ilKvPx7pSNNqdDVb+MPAJ359cEoN9QrKUIalYK
lj29wosW+HfkuQAygdG2JVmA+Wr7AwPufNdT5BuUuzJB5wGIjowpU3RJP2Gw8twE
YZaOkscrCO61JfxNFgpE4zqKlYOBBuABrWzienFsLctUYYF/JQ1eQCB6qzE1U5j8
sw69/+esG4F0KSNbd46w0x8fi1os+CbwAdUXLTb1NMVU/UVVHey3muym1v/Iotmg
nvBC1jKalO32Dfqb+BM7R7GTizKfFyjOl1AhXDB7omewgxb8CCtEOJ8J3lTcARNk
dY+8EV4RQIkYgOgHC8XttDRfLouxKd/C+Zy6y9HEbVWV76Ekzpi5L7YunjTVqI5L
p9JkgC92TyoFmzLZMQfbyGla98Du3ftKhiNiaFBDaBH9lkrAXoFy7/q8YYoQKvRE
Sc3GWXyT5yDA0l1zS8O1Z1If71CqVeqIG9iqA+U5dpLCCx9HqJ1CwFPz8JX7coPl
jbjarCxwaxStt/D9dj8onC8rhBpHvnwoq8BBaPOLivmitEr6/UUAsplu/vXKwCOH
woXi9Rf97yF6+Sxqq5F6VmQ37nHA+ApAvJ+aI1Z4ZVcDfyCWKsOqsVsQIfQWhAOg
EIwENhy0VcJcDllZGSkNDZTy1rEM7qdmB+PbOfVHfwvXEwC4aCd7BAewAhkvgwNz
Dsz17U1YDFIad5dPf69BR5gPoEvNacTXvOKUOiAD5eoLHAT+1GCdJ268mHLLyV8Z
LR2TBAphnrXy4FncCCP1Hw8OtWpcExMATXm5lgtNSrepBQisCG+V9KSUBBHOQyaw
j0jW33+CIp73T+Fu+AaBdyCMOx+DBef9zSyDdvOHyVYENcm7YKIvLJJqVo6HhdXm
wtlhU5DuXcLk/6qmhBV/jFGsJ8Q8Q1gnqdSruoZMii4C/M92K6+0i5aqxEaGjbT6
97hmPb47Hwo/h4foq0RZ1jbXq4+cZbaMeg2Vnr7kGTVSMBOvIGt97/JsGFdZJ37E
Y7YKtAIvPOQkn+DK1QHIChP1TJW7LkGw7+gcBIVAl6G5y2p0GEK9WWvxPPwVNXkG
mqmHmUem5snLoqdVbu/5vDN/2eNFsweaHF6dnJ/NPyzwvCp6HrPPtF48zbVJ6ceK
iHVWt4LoWbd5METDCrbd0AXXLplRBROIjsR4I79mHEYuWlBC3fvZm/fOZvShh8zA
nzzEq5Ll4TRlggffEy80TqKmvypY5FGI7zjf2TdctS1SOZRFzCp0nUz2pWFu5QSt
Jq94WkV/E9OgEcWq7QlGliVMVcmkpWDGy85RqTxv1IxNeZLN5oNQQKEBfEe1E+Qq
uy7wT8aZWs5D1CCvjYQIe1OssgyEB60w+Uj1Mui5Qzti2MW0Nl3HVRe7/2rghNNX
dwQxVaNaMCPL9g0rqDN5zL9FULJK/IWY1lQ+WAX6SMcBb5Yl1GYAMh0CctOzvxLa
src85KGCikE6LvPLD6ryAPVjnhGwCUGc96D8DyfvFeSvG9eHXelLGUMSowpCoMI6
tpyU3GMGCKILscQXfibat2egPS7O6SciiEEPrEIPE/4lYQhcUtppjhAiAIwbPhem
DPkEKwTjKftZSWrCI5b+o4fhexL5NA7T3AH+z7mF1ESPYFHEhQUsCuSQfc80LsEL
dGg/b1sfc11UAdjeMk+j1bgoMATkXf81uk0BsSKR4ajKBusMGC7GVCzlHlmE5q/m
iQW5VYbGSApT4oa2GaQ/pbImvD0K3HAd5kxLabXul5hXOghcGl6fcVSNH/wUDVXB
ATmXTnlrQ1DHRVVvSnp5H9CJERQmSN4Y+grp8vdK/n5wfdFW+jhJIuNsiaD0DD8c
3fw3X5PNKz5/ECGbwPNAgXK8INKV9/H5zlkgGcx01TyYUxZgc7eUpjEj5A7+SQq9
TUb46AZnthLeNo3DuhjvmbBlc54el/8WizLUnSgMz5JxncU/HHhZzdPqN6YnIdcs
sta9QAHTjP3pY7DYeZ7eraT1SK9qAiMi1TnsuwJqG0ujPUlv69SXpF+z02YHE3P3
P6MYSHxLrgazwp/40TpcDBkvpSBMDrVErHSHlxDzVkgAMt0IUT0/LDaaEyFtzTHV
rpRHnRsvitTRu3Z52B196FXcPWseJjZ5VtRzQ+8GGrXn7Bm7C15O5ZEaqaCdR0Sv
lM6CQ+pEd1OIBnc8GTBhlwo8MUhnHdIpJwy437ueLB6THN2b4ueXV3DREKYLvuhe
Xcv7g2u212ELutR7sIAhMr+giV75IpAgf9zIJmGPbZe7fu8xIGZOkepGWtI8HWMw
12xUGqrFmbXDsPpob77E0yfCV/OA+GxY8/NdStLB2mig/IhqhyI5nxLIaY4bM0w0
VXvcW0epIC41nTR+dNQspCMB4wxMZyloRz3/lyGr/Ub4Q7qVtMgAfWRQbgvk2kFV
EBtUlXoAMLawi3Vl36XdRoDxBV7bJMZU+TS6KPIQgOlm64HH1dfoaR0HcLAfe+xF
xs2SSY3VCaRSlh5f18Fs6R10VnY8+cB181YzF6FviXl/9G9IT0C2HhVL1KpH5pzy
7ryAQ73DnbE4RkTdmj9+RdRQx+X1x/RKVs0NSqx3/Gh+/vqCw/7QHvA5kibYDkBU
7mnhwk8HjNSkgtzzulgzEXwhJQjn9GuVLIz4CovIoW6xLDiEcWGuyRwiqYFT6hlG
APpEVKUGJG1Oe9c7pK9HxMYRStg4nhyw4cMCEVK3H4wOrh1lOc9pmJSWfD3kRTSM
u/A7F0u/oiNN8Dmlat4L4mr9kTQQBsaCAxSTPMK+i9p0XseidZRunmw88AquDcqA
cV6Oa13EXU7kJK4+mkEvL1OaN6YEIddfmTp+J1HmWnWeIlpea4yDwNZS4YOgwED2
uXPlnR1Xej5kG8rylFdnO+SIMMuF1JLA598gUkNYW5itdj6eq3Xd9Cy6GcncGd4a
a7VFfj9KFJdCU0kXeDapCURMJIRMk0hPCv4PBIjCKpKLuUHN2t7lZwWoZxhFicEp
Uko6vU4ZAaOCi+eW/pFF7SHc9sstKT0HWiKoAtdr1jTVh8sE8QRvfKN/kPq3Luok
nTXv8KOWqru9pzys8dHYXj6IOXaSgPGTmWZu4UIm6k3GaMqvyIkIi+JL/AnSCb2h
AKlmG2B4JbUuQnlKPF4ceuD6lHbwrI0wW2w+HJhUqIx8jp3Dg+QvGz41zWF9SwSh
1NlLD+5Wb4HkUTi4rzJ8Eth5ss7aZJzIHnqF42NKP6s+1+kuCuO/Mgf91rwbLxjc
zEHo0ztly4qyzrm2rVIwHQpbbvdwkzwMa+cJoyDUfmbvtosjltRUpqZzqfAWxbUR
7pP/N6oSR+8oGXzPhbtvSSUdd1s5YSg1wSKHnQR/jFwlr2Gsaz5XuWKVcqT+pyXA
clL22rqzoWsjUWC4E6Dx6n24VO44UU8hddsUVZV0c2T6bFmCfdDqeJA5JUNalS7E
JDbxycoOVvFuaGlBokt5bHo4k2W5DcEOYUtEHyvNcAnUFTsAO1P5+3aRXftCBI4S
qpadttqtW7Tb85M1MGH/BmgTwxNd2e/WDP6HN4s9/P/5oBIFphCtwExGfl3Nun+z
+f73bn7Qnj2hsYQzwbX1EYjDx/0UI1alW0mByzNQA9mGI6InhZXFuusKDAQZGnqv
WrCOUcTl8Saw9ws6MYK7/zuo9J20LnK5wvSMnRvzYFBrowxLu23vMe9MzK5TEc7O
px/gZxxvQdpJzjVUyqwGyCxrn9TX3/PCaQ8kIFcI28hJ3E0ofvoSglEUdc7wUPex
Ee9bV7V/yTInSVx1QQVg8+VmBdl61D1pn3pZvmTwEr985+wAArl0x3LjZPf3iep5
J3UraxjDXYkEpasxywjXwckhSo2bu/0KMD5GfhqosFfyr5krYbK0NlTRhARHh8io
b6vEJNXxGZKvHTa7hIHn39CqycNgdDD7MrcmfE5iMysuAAY4LI8l7Xfhy0vcmXCT
+5k7F4xJ9YryEbQa4nXiJFLGxkKAF0TSvztqHURV7KLlLlcVfk9L4UERHPI7qDtM
vn9BmbG0Isw2LP0Wszi/zWIe9wtX1keTz7J8QyHZ+2Hsjomkx+RSVRHZwdYG6rXT
dSQFOGykDNDLNQCteofjQ4nwUkzcHFjPjbBuNjs3kK3VQL9Gkv7qso2wZc1zLGif
JUSDyd5vE0KrcT51jeu9KbMvYu06hdXnCF8Gs2P9Ww/94DRQ9J94sCuljdsDNk3W
oOQZ9bZr/7H/BshBdwh92rIhEzb9+tfJAXKbtOQ9ZZe0G5JU0AfIcn3/U6rIfCXb
VCJ5k9NPkWGOgscbXer2iIJB3J2QGR5vJxKIB6q+p/yzsYly180OxNLs6+8E5rWW
/n91yoQM2s1xxaYzgOb0BCg3w9ylsalqBW6/ZzvixlvgZmBxU+TveoeWkIIZK3Wm
edMy1QRIPtjPPRPG6KVXBI6Icpbm4A8e2HOBsJRshpm0LrYdfJ0BfJWQ1A20snz6
i4y2qnBDDzY/OXAeEA9Ox203ECyKAi5uLwvxJGUltfmLrHPHj0lF2LEmzxNF5mEc
EnxtmxGR08k5ukYP2L8PRfSEt1WOQmJbKm4IOctT+Hu93gjF2R/NOzYPsSfJ/uMj
WETZbHkOk7tRE5iicZ2wh/6Qrqh0vfWCqPSDJnVZ8HF2f5L+YV6yPlGh2chY/gOL
wPTleOqFAd9zADwCiTiqhs5G/kHbRY/T7WMrzP8quG3ZqFP5yxzXg6XMO+7BnmIx
PlQjCmntHsUb5i/Bd6bbr3QisHDBFQAL9JkuQ7YCUoz+ufXuO8f4dxhy7GthQHYS
LyanaamvEIarpiuNSwbJpGk8KoG8vMX/6CvJifLiy/5xypG0xY4KExpjTzfcuq16
N6cA9XssOm9Y500aqWDZTqeazU0MgSBDiIH8Q5h/phOm/IU+PCYDb6HtYid7T4O2
vcnVca+6/FXelmiWiihmACgw0SGhOxEtwER08W2Ar7hNSyeiD9OyWqyKo+eM4oDQ
CpEer2oYehqWgjlE9+t/SEPocZNHpsNz6WWpiNf72lvUGYaR86QNIFSG/9fwHolL
//otg3FNCjKm2T4O6551Veme5UFwS+YB6j9wIMRrAL0IAzq/fsY28CwmfolWlRmq
LLgZ9TUvXu3NN0pQ8zalvCMIvjbPP3cKAbz82FYRYyqpNrIJRXnudAZRHTRKXtNb
ygMveqump6AavhW4HwUVHiTU72M2D3XPdjKK/ZGuYLPRgZnZcPERkO0aJ4Rmz2sN
SjYW4IXNAPU0XHvQ7kxh88aH6TeK3Y6EcPs+/mL97tx6K1+HHsS5Ui5H6KMWN0wD
BGZeElgg9UmXTnvichd9pn+7Bxj0BXa6F4frioOLBjaxAnuMbzYVsAuJlX2UPWNt
GRLGGrtotqhZ+uX2F+K5wA==
`protect END_PROTECTED
