`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ptzaNRuZ+PnAZ6Q/vQbP6Np9iHfBxmYSd6FvsA8UiaRCKvcepzmKondn3TOYwaup
t3RLpaH46EcetzbkcxzU6zTX7IfZc13eXCRt9OopsZ6Pu4LFI2uDAPrFLO6lj0Z5
6klEhN5N7HJ0am0Dv3a83xHMEd6P8IXxL2zFxxsqxMYFumGgDdvW4drBoE6gqVUB
tRpbEnoHY+ABoHRiDpsy4x91VNxVG9eNybLkKCk8rpkpR3mY6lTPE/0jax97vlFv
sP8oFFWqf8V0kQhG8XF429we9uLjV3kOtewu59QwJoMJIxUV3cCeAcjChAN4hhwj
1/iQN+e5cSGN8AUsm2FKhX7spJl4gJvK1LhfP180pyNh10ppM1oDZGu0giUFsT5P
3/DFytM2hhxgtuOOBMiRdgqECuhUCylj75B7s1+3qNA18RLnmwxUHoH5F87VFzCd
09VPeZTUWhzMwFNa9OLs5zWVsC/ErgYS1lnzx96SAI+lmqr1KQ7w1sOSHFG1/4Ty
KWKMjdIF15TZTCHld8FLybQDo5aod5ZKCuQ6Y49p+IW8EFFn64Oxzb0DyVv922Jr
xs5CwO9Shcp9kBbZvScnwDkXhVgvrPoB64t3DT+GDltREbw6+Z3/rLTzgeSaEedU
cm/fiJusESbGjDCRgoHm1v69Zs3AkAVeyeu8zyn3hCkx2RUlqMY1GDqq23YzYD6n
fTnqywVcCRrsLBHupAq4Ka3UGKVbuQHjP5jYn3IhmRnIRY98gbalZuyCNWpQ4+4H
faGlfI5BvOIGYyAMBfQuqXQ338d06NGbRwPsrO+Zfe2dqz8yPnuEjSHRoHQglmlO
VfnorLAutEm0njdc/JE91+v4p2pHM5P6hDdFmsFxGctsojVtcLlPnjyBTad2kGhJ
CYl/REDmhRWYJ6TYi32L/GTOnf38ltaTVBUsWh5Pqy+DaitkZClK4OqYJiIkEcI/
mTu4qj90D47LumIkRTWpiWWdqiifXxtkx1DOPwimtojHncmePVUnLGeCUP8rpRwm
zdj0HjCxkndxTYdaA2WFxzPDfuMio11Ix4/wLaonXJfFlfwh2cL2DjzQfuj0zOvf
T3ualFBZHTVH/nLt/GfJPo2tLpToHjb2iCGT+3tVGdutNDWtxNT99hgkFQY/kcsF
24I6+CTM4axlFBQqIeQPt82JcvWsj9c+hY2nicSEKU0fKchEoD3CN7EWfq+NUnnt
KBqEEqC9+c/7PglSPX0Dkchqov5tpMzGyBGfE9FjIbW0JjQwKjO/K7UPfOkBxkNW
t+I8Fa8Kj2I8P5uK5t5lxTLTLWZ4AZNLTw/TI/bemTHNekwATvi2c4YVst3BGKvy
jWwXb96A5V9U0Kvbzcg47miTU8p8wumKXbZvSyBOmWn2jLTmfDhtkolGgiwfGDAd
eMtvfymhwXf+x7DC3imPUENcIUIXa5dB4nUzslQ5eT/HYMLAsQRN4KuM1v4SHp0P
SbcjOBDA3I4INke5pHYewzx/0RgNrkcSDDyJcj/N3GDCnp6NJbjwlrGf00Nr6fZk
/Q8TaLmzQk9Hu0wLicaMB1uWQkiLfwHRrZdZnobMGruYIkM1hQMmHvrah0S4KiiB
BcHz41LU0ovU991GKOiBDKunYH6GJa46K+sElJY+sdwFybhw3NtD2TeHlMxuVq9n
e8FJxM9JEajrutJwWyYzBJ8iYddLA3ba8yxnrA35qvGvL2PZED7XIga9xFHvrrNQ
cY/4pitRgWlp5bRbRsb6EhdSPKaR9ZsdXOuNX0gh2/OjnyUrCT6iwqyicjGzPM8n
jRxZ4kMc918BSVB4R5TJtYw3XPrGN6stXiXj0oUsFB98laC1dULW6Ikc9QyPfP3o
GgoMIW7fQKOBTSJQcT0K6TCSPjVsBsKkZvgAIJp7RZRlVYKjCIZG0Lh7LlToBrKy
/XzxuLVDO3fp8SuO4f8Vvu/ZNk5mHuHIt64OyF5z9bLhAsOSEfYvJMr1GkeaH+PK
4UWrsc23bPPt00Qj5B7gaUNpAuRqZMsrTX9QckD1wQT7f+PIK8sjU29gXj1BWYol
Wu1hg/Ahm1OF8U/JUpiERqasD5NbWpoF4bFg56RWWUT7kfgMeFHjBI8lUVftyVMp
7L2wHk/Fq2U2RsCiuTTGr2lyEgne+lzQ19RuoDN6hyYJ++rd3IgtATtq5x//jR8b
KmjkV5QzDg6lIr4MTIc3z/5etCb9jaYhDqh6CtHCxi2Q0NcV0carAZEvh5OwNoVc
nGXlgWVCHnOVCJKMRz/pHHTPjEX+tz8Mh8I/KKhkPbEyYFgzAmQ95GfeVhQ0hcii
oQe3OR1YFNexY0LAq6khZSdNK7JB6ulF+qncgvobSAsIxvvO3rBX4mF8OiSW2gyt
J9md9mfC3SAuDEUVhXLDUdf2i6tucl2A+NYUDpEoMoCxtupHT9eTqN8b04GvBnSD
`protect END_PROTECTED
