`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oa1gQH4uQ4lchP9GKpMVB4N/9X4JRnyiP/lJby6RNiB7HlNX98Vech52O70l6U6T
2t5uB0XW+uNlam0lpH+1u+0Wwk5vmOvQ2MTpFy+g1clMBaYL0ExP+Cl0SlMd73ma
RPS6ncblqlc7rX7ZV+drjjYQoMiY2JNOYEJ9VxzHmhQyxW0qGseqiraOZUCYX1a9
GKsGvSYQ+nYLha87bCaQZ9MWfXXEW80bou9kLlKVhALAnWnxRxnqTEkb2Ab0X1er
q/BKs7gFLLLPqUOfys5rAm2o/mufocReWqK5aMHUvKgKPe4Ucd1Hp86y7lJpeXNw
Ydw19qG2EEWYCBLDPoCo0+5mWWvOsmkO62j1rRpPp02C7aG5osrcAcVJRYcH+1kK
YLHZlvHhW3yAl6gFu90VNcMOZ7YG1AKRgcRju6YZuP9vBtNyGrT/66l8fatSrgaa
7bmwaqDGoa0O2KnTa16S/MtHDorDhe5wsPmM0z36Vn1NVjThO4zo9SbjlrmjWxDh
VAuK103ARHUwuy9k231/VhiYf+aXI4W/I/JhzvnHnu8GKFcQ8A+qiNs7x7w2EGpc
u59UKXQb4GDsjGSzVkDNH3G4q7tuG9zzt6uIrGp6ZKMIPVYHGww0lKMsqDEq99uY
l+eBdIDZRMD3AQH5LSquPx9GTNy9vr2yZmXQ1SCAWeimF7/n3gOo1LbYyAmV2rnB
V9CqBl3u0Fse2kh+tGtuBsdZieCW4eUvxPF6S/QpFgKxl9co8P/bZdlW89RU/3/n
mTnxsLNvulDYRw7aePgpZ0Bmn3JFY9CYFJW7C80zisuPtYZ9dWZVDiRoMXGXKtzh
t0LfkarntHaTw9H+PYd8lV/s0sd8CMoq0ZgSE/Uw1E2zkpHKUvwhbrz00AdCZFO8
ksR5wO5VX33dxh0f+H7xIb22xaIxToFizhyxRmJrORk5N70n1IUKAfEQxCLeBPbR
KPHgcV4X/W8MfJszdUKFL6r92yyyORf6iPP1cvmdsQ0b/sPmagdoV1mpO4z+VtPT
VGKnNYkWDyFqfiDJA82hW9/0QUKcHE9QFfeMjJInCIq/0Nu2jBuIBUxxfvjq4OiG
dJeGZTfHmJYPAd5oszi2WWVBArk4CflMaAXGuwrES8cGXmuhGPTLBU7bIv4gW4jA
1O1RxOoa6MqhHZAZUytgS/mzxv2OIuk7JeI2l89bbEKXjJMhf7KNOV3OR/f+oOIy
3AIC5qgu0zuoeWPasciOXGV2QQke3czB6z6ewnFzwOME7nprhLLoGVtKOtZR5qCg
xxSuuW3RQ8lt/f/JQdDDpJ8yxR8lcyXCUBaOQHDK+DLEduJtXOVTYSyPeRJls3eV
5wI6cS4JJVaMJVBRIsSBSESQIzAoNf21V6uURC8xFXn+Ub/gmaQ2Rb75ky24GnGZ
0rqy14if3JUNEA+EOl6DG/jO8uWEUbM1dk881NNy+U/+BG7DhuufECCm8va7haPc
GeRdeRhDEsxC2orWqyjiLGM3JYdPJIsOBKDVAg4scIuBhK0zlh4ec5MqEOxHERQN
oGjjSctXcAweVunPSxbQgFy31rWlfhK+rql2BJuk3pzO7yu9njjyXQctwFRq70Dl
tKtO8BetQlfFUfNZyMIOdKC6ZsAq/MHUail1oFsQ+cvN9awBSnkqKWXSa42j4j+k
dZxi32CAkdmAda+zOjjchYaqnu9yc3bJyFLRTGQkxS7Ha8cDywlE9aE70G0iWscK
X6G+E6CANZao0j8v9C0avMf0Y5Fa8nChs2t8U17XDFwYqkKOdY9wfHfFyQ7iDuf3
Nfi/bsnYkOzj2jdFDo3T6HBKAclccNhxzBSi3MThy1t8vpYkLtCQ/mZ+M6Qqv5dR
469pML1NEcGn35HxXh9WgRn1m3AyurVZPb7OKuXMc4rKbTMxE7egYla0HBOA0uTW
3WTGxauAyWzJiUBlVBRozUIG6hjqpP3F8dJHy4/PBcXAzJOeniNZDR8Jrykv1RGG
uWg0ua3RQKDIeAD0Sie6Xzbb2V7Cf0mhsBOo/ByRyyRnS6houNOF3aZp3fiX5i8/
U5yf+NP1uPheLW7R5DyLBkWmGfgavNLLzeMBaG5anj88dG3QEbqRuVqtjyxMMaS/
eoqMp53I6MScjxA/ELPC9BieEO5CDqStXWo+/4TZt897/suiyfXIJm2RV+khF6J4
P1qpBnTc8ID+6nCXooZfBB5RMSZV/QQrlsiatoQEKaNgi/liTPw+Z6+FlfgTK1aL
LF0U0iInZtQNONEU4P7nhXszBjkkSl1kIrLfIFpEomWJmHkUF15SNlTB0NERHLBv
ZzJuqqdunIp89mOFr/iZIt6bHIbYpoXyGIf7XjmfSpWGlCoeT2z3kvyEh8Xy5uc4
FEyFqse+pYcyWeLRKcA0rCGcI0UW+a/PQcLjBtnlt4yk7shvGTRf79P6TGV1A3Ej
wMdyAp5K9ZtE6s/RdRrinzIOoqIVBYTBgmlAPyNeA8EPxLEdP+0QAnjQRxdBvjm8
k9kzzaFBhxQMedCSmtplom3187JVdmKsGGhVY9RbZEs00wpU3re0o4hzkDp1a3IG
G+zEd+8UHIcHo5mxdd448d/IWupmIgjsi0gZSQN/4MdUF5UBmbGgkFAangXcThZg
U2Vvqx8dmoW9L7Itcb6cBjd3+w7b1nbzg5Tyo4CUt+7QY22cujwulwCsKQn0V3ea
BEqQVW4Zu58QeDSNYTMQagwudoEJCsTEUeboXveg66aWvvbECCI0USIWao6A3L+7
c4XO3xF3wUgf5kobt0+dEcYcjY8AqH9iw5kzCMeruHaUUjfkIW8/DTMardcmPMkJ
bBn6Qjx95z5gcqiF/uoLuHk80pJw6qeWw+gl+Yiw4CNOvBrLlTOOBQERHTzvNf/s
54i/wg4XL2ukBOvBnHgLNlynnq9lnj/kpyrDdbA5UqoW3ECnbOHpZRgWBJ2DI+9e
bRnEAhBUMTqD4MSVdgVqXT1TF2AeBTVPbtxq960IhBxmo9wSV6kSxEG04YyX0mtM
IVf8rtRnXZsy9zTvVjgRMxVQBviPkUJg63g5wjolr6MuitPLrdWTXirWbfb3HNCO
DqpXE91ONv2XST4k7l4+5FRSG7gNZf+zhnuxaKLfUrNB6XmK6TRdIGFt3BLCf/ZL
GrSIQd788NqxPaiZCRN4aeSwCxzRBpGs/o2vPgfE4kRCbbvSP3xs5fekW11qaDXy
ZG0duHvR8d4rsof6JUifjWU3c4zlU/mNPWv86nXiS1rYW+k4BQkWqHOkyuBpMO4p
u3/q43ibDW8Usv20rBuX9Jc9V1zsEbNN3/zYQ3UffDmVSt4eEf8t/MtGLO/tX6X6
ECmFmeRKy8n3nEjN6iEjQZMaebIOBUTjCUNHjKMIeZAIi8zxF78My93FKhEoMrvU
7jtxwvM71qbFBhxqVK81bJN+J+UkcFeUF6Jv3IAfsGA3erIKehN4kulNgNN3fi/i
Ra4i4P30H2xFUuMrVAIkiZuxA81okkWc9f1bQnIDLBdZkRGegWsej+eWJi3A5tSK
ZDymLSUQPdAmBKHDfBcDkwW1sn9izIpByRX+YwmB6WJ2nTMSbaCmkKF41F5pEHLM
Vn9ZzTzrWLhxQMx0G3K1RXkjWiQH+IyoQoCYSteCMfRbV63H41wQcSyg9Ti8Hxjo
w+Z9i01/iT533ei1e1R57CX8y3ETGevuLd3g+jkLQ3FJBtPcWm4hZ/Xc7w3tZh7C
W9o8MjbQAuCi6LIYong/zpnXoAO50AJU8krBKFc6jXSQ8mAb9F59M6lpAmfuOGHS
8OctbU7vp+Y3k4KmYe0PQK3KuERZd9DFaiArYBfm3rpdzO3vOTdUR1YTh7Rd5aaq
yb7MAz7FYNwqS7fotKHdWf109GOj08/Dzpt21w7qsfYkpsl4+Q3QEPMOKoXlZwA5
wlmyhdPiMzVD4xMQdw5WRpHYCqeIKnTXv9+AEsHGndf9W9kJqkyhCl/oMYap0wtN
2osfdvgBSHjzyUATFskiuV5WkAQ1QQX4pH444c3HDmxPiNDMnuSwe6B8pi+6GmKe
D3aBxBoEVeE5S0yiOhsGG8r5tEjv6PoRDEzuUPajGP1x6ZCcG0exuPws8bktEzlP
iGxilWbyvH0KFEKtmbFc6klkA4V8SFqyMAJVaG0J9dkRtD6F46cdTML+BQ5T++av
AEACsaX/isC+RZ6P3eTst4498SZEO532ExEjWHvBYBiisQe7luf0FbiRWjdwJqE4
IavnRvCIg9mTY5QCF6fOEZJNtiEIEuJ0Ez2971PyO5Xj85BsgPTPQGT8MY3kL07Y
dy9012cmecJn8mS7ymgQqmUT4cKnGqrCF6mWaMnYgwLvrucr87MivndvesuJWPZw
iTdoa5hVQGbBGq0nOswZwO/VurzFPySGMwvYgtsPYlLicedmQQKdCgKEBghg48HE
69OV67R9j1b8SuiDKkQfx8unGvIMQdbRUAFsf10QN1ezzfEsAwr8cnU6qRJCsKOn
mqvrpvlyS+YLTyjtK8wC8Eq1v9ShHBZcHfAJfiMTzjMydZlHB0KEAJHZg9RVtege
1SecKry332dC31JZ0/XXGS8ziJCgqxWn2qeQvcJV9KHYEZO4Y6fsWQfT+wvBVxWk
`protect END_PROTECTED
