`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wmoe7caVE/C/ft8K2gy8KDglDB1MKBpwqS9C8k25wuYtyYgDcfSxKHmGjgRqLmoZ
UwJ3jTlu3KXzE8rCzjIpI/zlUawMbQsjCBq8tueWAzeQOmoNZMtHjjAViEZr9Qv0
YwCMrfiFN9TLQpe/a7zkIun/d9nlhc6918oyQdJnWbhvuHBPuN2ri2Tb4DBeNmJ3
aKmlKLLt8nnlNVmZOfM9GsJrXTdJb3orcUuvbPxQB+LaiVodTXkuGePdy/HybgsS
1uixMW1eL07eTVUFzV3E1E2cIOVtGWXA9FnLgJjqITSNYATW382YU3TVRVudiRL2
aP1TPadl2ffAe3gyR1UD0mc8ClOvWBGS6ymTPOCMQFON6m3kPp4BFsw6TpAKYUJ8
DheREl2oobw33Ve3n7X3ZPKlow4bIjTWKj1II5kbvinilio8MBoL26kpO+DWrhhe
PggFdOgM32A6cm0UjfqUU8I8lkQP3eU5xTp3yiYxfzHtwUPL2j+dDF5Uz72FHwNk
UZAkVU1sKtlvJgej1ev5JeUFPiZMl4eIwahWNsbcpQQzUDBQ1w+DUp+Ubcq8883U
B4Y/kBdSJP6aA/QIw1CO3pG46LQ6WxLvPmI2ljD8vitOYDW2x4wGBOaq1FArnEa/
jmhRLWxrBV7/6V8CxUu15YwUAD37hWLINWtsaw5yeQBhSisnxctu2Gnq/RgqY3Zq
VkyYbERioRDdRz6XbYRCVce0+Tz8Y+Cof7JN63duT06fVnTyNccC9CJk09nnhSxv
ifDAAkDHImSwnog4WACXuOrQ4C4UpgbDXJVWB3lFihhJTSKUAFvkO0MxmvlR6lk1
aE0cLwvzQ2BNa6uyywwEND/TTAtDXKMQO+7mQu5KLHYbhIP+Utor2SELGTYDObPJ
MOtqNETbkjh0OcLWalaU01ISCDKO+ttQKBG4uGt7/YpZUCNBUTj6M1g3rKnO3adE
T1lpXWBpx5WHBcVjp/JsHJEbZMEi7ikpcIvaPqgqW69ASqKLQH+81/YOEc4/ddT7
ugezwck9dYz2VYHJBWdcM+8Y4ZOI4L1JyLN9BPNxtM0UT6GPMfkQhPrYXygT3rCY
pplfpFQMruq42eQxxhruKyDkw56p+T4U0SK2FOiJqsOPv8fVpE1GR6iDTE4dYeLy
psaa4GqcqfWVCeZACRAmauYbGVfNiYXLba6Iv7m7fxkzkWzik2wNrE7xjrfZn9Ty
et3BgAyhS/WDGMO26eOD+4rfpGhclIQ4yTeBoCYisPt0zEt8P36eBJRmdngHv98K
MJMNIk8JbkV4QwFz7fY+4qSUHO/P5h1Rx57v62crVnazK1iloOCSfN4YF5F+zpz8
bEmTA1ZtrGpwjBQk+eFx7Lv13gF1NwnpVX918qtUpOq+5y64YyNN82p+qi74sAvc
RFj2CFWkF9mP/DBxg7v2K7mFql0hi2C9a9jChS4l767E6CBBR+pXm14g4lhpcPuE
ph56wfVqTpEWwhVH+/tH7ayRNFmHZIT0eDh9L1TApqRS/BEmVvkaHpEiRdcX5tG/
+pR80qFkmwwD5NDBeZ4xFX/qD3BErHH1uEPanz3PXl7bnkBaEDSZWdOHiq8mFT/N
3znMKOKZAoYMAFeU5frvyiQnhxxEt/ze/IgQfd6aG0EF/q3M0/M7n6t8hc3hRnMv
e8uJ+XWJu7nQ0kUNSUCczJl9BVbVO4eHQhr0NX4ETnTK6vQJYvMvFoxsomciD+J5
LFMop2IUuu998k+f9bZtscC/rFa69FJBVdiBlF9JKendlrcHNoB39hPnQRaoTKnx
EqN62w0DJXE9wBYo4n61HD84cizV2UuO7IuMEs+u9IAcgs7x8cjNpRhVfKPsqKmC
dh9mEs5nLbHtNQROJdIdb/Iu+X3eiev21deTJnM+X4puSz+dIZOZRw5MzDX8hGmP
ww0VMDSuMqDbZlL2auDxCTp9QDFc8aNTDPsvVgYuEWpbXqD4gWRAQ4MwR2tiIjdl
3Kz67/hXF5BNUjG7xmBd+CEm4vX4Q1Fk0hLukX155wocviHbx21sXoBlhViqiJDb
L4TrTF9OUKLj1pKrywTsPxLZiIY2mqWiQnv2buLhSz3tztdhSbDH1mHgQB6o6NOh
Ts6qEou1Pmr8Yb238ABaSbOE/u9Sps0krLXERrQJTXr5Askp8yEtJl6+szdT5SVC
nhJ5R20s1wB1COcqvNX9MyjZS60oqeZSWVFGXZBUPpxq5OCvVtQm1T9LBXYFzaGk
QDyu5p48PSURz0qCtQeQh0L5o0c+wTVNF4OU5XIToAwGNsE9DaBz/mUkQVFN5f93
dY4mzTbUcVXAn1VSaOLBRKGlzVlul7XWEkRDkp6DPYyDYTrWNK0NQOuDb19bUVVq
OLRLNJY+owd882equvWm5+bdjN8peOpEEzQ6ypTs5rF85HUwQ3zTPi4byGsHNl10
2vymnOrarHDdzH5UWFzmfGyB+5qtsFgsg7i+PjzUCkYSEf+FvzEpbz4w6beYW0L0
zrLLcOCzIFGvLH6Jllt7XXHMKtdvA00+GGOM7zIQdUxS+8Zl8fMZvZ8f38f9CGsU
aPAv2a829a22KrOnyZG3e7l+o/KmH8ZhPBz0rS8HFawseWUd6AqcrVnSHbl/bT5w
00yAXsRIIJBQicj+UQhG9H5L7IibwWQqDibqjEUjgWXnXzaThcRjhYSI2fEMy2u1
flKRiLfg8Z13KQvX41L83+fGuHsElCCwGWrdP8nuOXTFJTTwe3KEMI6AsZBmhLQP
v1QU1feghbSmfuw1g3nIp5vqYm3d8QIIx+oRjAZ9pGpN3zlSby0Kn7E8TmjJRUTJ
YIhfB1T7mdsgjawLnNQN74lIlp2KarMdfL0j2mZwMSZHYlCitCK3T2HEEVO8N/ol
gJvbFEtq+CwEDL+/9RmEcRLBwsWpR8QZzpqEYj0NP+VPo6VjFLKucfQARapHUF5M
0qj4lQie4Cvq7YcYpkOLfYOo1qlO+U3FDFOkZmU1ZBSredoSAxWY4Xwec0Q5Pd7L
LV6Tvrv1RgSCQtudv/5X2lRj1L1/pYYnajY21Mf/vFL+sxlkmkNyIIr+ORSFd8DK
0w+mefDVeFRtun2UnHNS1ucQ3kc1bHoDQ1hwn4cm2gGRobTDZsFaf62C8cilUp2q
ne3j6HBoHBwcb8W3/RjkfeUbdXfkgEfo6RwKbYUwe0DgFmII+QDUG5HEWD2glYaw
LYpmCy36rBwPalRFK6KWWR13sor2P0/XLQdNbX3JxfMXRKonfoD70pZJIKpnqPNS
IYJWzW0Yal+E3qFVhzkjQmtdTFDZtwdi6MmUcgFKBRM5yt6Ok4+zAM0eELz7y9YM
t8As866P4ptFY9vfDv2UYdy2FSPBUzhbCJtGQzgoJpFWpn28udljOY/jtILMcyjK
KOlq8a3TYwGObbNHS5G6wpmS+z7/IFtnTCLw4CrpF58mzSBCzkU6Kyg5xTlB6lk8
GOrDl2EmgNNSRPgbOfTwsrB3p9oXsexILQTHABt3r2/aOumL2EhKqlVnUfnsdB1G
jxft/bHxfzhdUJa2/jqZpcjpt2NYefeXv5o/a2/09BzMy63+VWGbQt0eTg9DErBU
Zvc7jzhpCWzDdh9UR5eJjvtkFt6aqPyuYNGFIpMgEwOBNzXloxqzlT84x7A/zqOI
aq8VrI29E3Jx8NJoGGT+B/7uhq1ZqOa1Bqt6nlRfIloC9ruChfto7v2bJaMW3R8S
ZAl9zLzwbQiqyVDx7LSSP8FadibKKNccZbJkHEsskwOZ3s3PLsidxWIvkOXe74bt
IMyS5GNwLlpm5ynF6lR7U52+AftbHk3PgEvsYzVXbOgcW+0yQWGr9IdC3KLSR0/1
gC4v4qz+CHhBLkNvPnaj+1cmhTSckuvqHLbj/ABwjKvaaXJbbenRijEPRa9kQLwO
7xvdayyuTK8hMZdkbbz52PY2il84LPwuG4olLhAqTIA3DjbYBplNJ9eNajD2fxGS
75dI/LAP3Tv8sQtlMBKeWhFicoQ3R+5HIFw5Jzu1DubfHLozPL8MroLf8et1H1tk
aWfZrtGSSh6Mu1xzpyXu+pnj4LN/bictckUUiufsuBpniegcsrXLVxk9Pil0tNfQ
rzQhjwd79NvsJ5Nbzmdu56iDD3zWRKNLBjdDItfiBKktkxW7zTa3k9t28xmRyYL2
777dqbSxPw8+pH3w6AO7Xn+J+sULZCL7fpiw2RETj9joxNrfnYtZlkuXN4Pw8nLY
MEDWxq7gow06g8l9YeqI+4AGUJmr6ue7VKxaSafxbzkrJAq0+cPuvfpSoA0hecid
jLucNRpmQhHhtx7dTlROBLjS9e3Z2+U93JH+nOzOrf7PG8XF43H5xHhPKWx12aDU
ZEqa3pC8VO+OxJ1aNhq4efk9jZnZhlihe+gnCiKIH09DpVQiTNmQjzwWMJHn+huj
p8SWJLJNs58GNZ3POjwjPphY3NJp/2j5VQufySb793IJPi1WP7N8X3DOP0YGIGba
29ayVnJ/mnLgPvbAvvUqqRPcIXyfaHOBNmVxqgHZzBlFcMVdKpZBuBlzdJZ+ochw
5cdnUOzn/QED9zv928EntAsNw6LDW19gc4FHWoI92r98fdxmZNrfj2NYjjGwyCrp
6unWvIR/vKLua1/74Qr+rRMoVuXMNm1fXEUIL3kSFQcoryAXo3HabDNDAZS29sle
7iuxPCFIliIdC0zOAH/iUGmSYHq7076DG4swlVzjU9Gdypgb/eMd5zH2nhQ+dl3R
BGOesxV/KlqH2ZFVcX8P9BsZaYDv/tMl8Ipz7QhWBYRIBYKDL+1Mj04vometGBPK
ZwDKjhFLVIBBSFpa1ty4o1JXzh09YCV1P0GKPQLXKUNppJRs6rzerP7XVOe+Aywx
WCZplpVNUr3urdEbuqL/h5zFOBIKblVaKMph6DymtbXXuBEwzaUivCmJ18NW2iMi
SqehCxxU3pivED/1DCksAetRyW0Q9fRmfljHgoayOt11iMXTslZ43cVFGOXfIPqQ
pJI7jCaL3EVVLTPvYNKruiNIkLvCpCxDHayHC9NNxxLycv39YKV1lf8GdMrCv2aA
6j7vHAKXrktARRHRooNoVQj7W41I+JafdU8Q/Mllyt/COmS2s8Wg6BBp7vyxeqFZ
9qIykMxzgx1GvP+fTR3Ge65vhmhQMF1hfPmttLVeatPbzaA+CG+Yv7ohSDFofme3
URcAtiWu7vLz6TYlh8deMSTnHT6RvLaq4ZWCXR4qYZqmZlAbmnGBqKTUfOR5MilL
+Vj/EhaB0xXKm7Sk+t2H8WH9r89XFPLFSy1P2lC76AJkyFTihpKUHx9vqS3popfv
s1+lrMRoL3pZfVT57E6WDkjn4QRbR4PGN4Zk8zjScTkCv3aWh2ZiPT85z7X6sTtZ
2Q4/znqRuQZqZPQx1Q3B84N9G0goJB11RHUjfOUaMOvJuCsH5rkGZtSReYQTlSta
EzEYodgIxpv/bLFfqrMzruli02fUFFQ/CPs5bdMyLwEukSHHekcn2NDzgo8JG3Sw
I8KmYgkudO7WKxJOBESVuOppG0UuDh/v6zaJdkACvi1gUi8m0zDxQJcoIG7apweb
DwSCJBJslCm+x4phmSSa6pdoyIQ9zxupmQLW7Whl+Bpvpam0tjVEHDZtqLzgS3K6
eb6hupv2MwcLzb2aiFO0JB6bm+xYmg4sTokyiycjZaL4QSJ6cLKyuiJDZpDIDvOG
bmT3Gdn06T3ZC9gv1MqSdkCerBE5A+zz7yP1Z0KQPYZEvQlL5T0gRk8EsZVtQV30
W/FWncpWqNRvyf8TOmB8jQWcO0BSsHp4hZ7hVj08Ng89Ya4O/uyZJ9twWK2XvN2Z
vbG80C5vjm2m/uXHdAVgYqr3TsrwKzi2MPEFjlR2qm4ZZ8jIZyqfq5QVUJQJ9h0k
4Fy4Ymf038pGcr+JcLqxx5UsGwGmYJLMPMWQtOx9ZXVUHKqVOvInZMLVPvL0ESx+
A9eDsN/fawnZvIdmKl1Uafdaul6uCAWQcNV3UtxrwY1HU8K1w8nVmp9/3wRnj46B
rW0SfA3X4jo1cGLTy6NHjHNoOY+yj7V10TRrcmeFLrxt4SArijyutyFKYIDTNROE
28nuujCEBo5hiOpoMdbpmo4disjJqg89v+0IbAJuyq0ImFXrBPBy2JKniLljfesW
PGChb5YXZ12RkApGSWcV48ISfNKgOw9rMyI1Is/ltWE53T+z9xCIvSavgmiRvwiA
ENDGzmdEiwKJa3ZhXONBQvqPq6kDhKe4L8XasYuRcXbnoeOjrdudcPZ73rqhIQL7
JYd4vBkshFcFQXTsq+2cTouV6RrZXqdlhq79i/zoBtkk/tuCVDNTJUxdavh+dlnL
SMq5nRZSAJKmev20r2r1Crx8kCekA7jQwj3YVwB0/pCIX8gzju/z2AXR+z20n33H
74ok+4g6N0UMM5YB7+NH9PkaU8akEgPE5NVSckcbl/WLNGK3+b7MEG3KzrbNg18q
HpOtb7+vy63PgDqqw4o2Q39uLd24z2I4hjHjgeXcpmYSCuFU51DtpbzSohxG6wgS
U5kIzXYqz+s4wFEd+G+/DLzPOTVzlwPrOr/C7s0uH0EUfiyDVNEZDB41QTs/QJCp
EK75aOpLHsQHM6EU+wl52qyVAMQj48d0837bfJR02GoIj8O3DpllY8+RiGddyHQs
KBjSZeaF54Z1E3abBu3fmqfYgp73nIiiil2C1wj/hTfNaUEB+4yXV+ktmNoGaLRH
HTTFGcd7gSa9oCdqcY29Tb04+ceClRjMWIa8y+YqlzZJnXgenbCVEREcrI3Vt1r9
P7ow4OeD6zQ+OtXk2TofMGmpiIbO5SPfsfa/pDYb2yyTxafEejB3X7ISevdIFzkV
8AM5KKnpcggo7hH9y+pWt5nY6O0EMz5JfkpujB1pCNXSc9kD7t3Kf5+n3vZQKqeH
Mk9n7TcO264KBFQtSOOvo5zaVO2FGXcCxqdoLJoOM5MNOMuLqK2pkuqdttMDCThH
7LST5rLw620gDoDPgecnboBKbcdvwL7BLt6Lb7fK+DYY2VCLrBJqYOb7NA05HgUV
+LvS4fgUjJ5itRe30QS+7lbVi4OcYQnOLYUjHlLZgdBAzLOgtGSqYQgdLTMhzRiU
UkonLPBPBI7v/txfpYRM86h4W0Q+iWsVYk9Maja3x7zXyzxKYdeq1cLwJuLIN076
kpSHcCKU/7i0rfN0SD50DpUMYzTOihF1PRe1sdT4y/p9VZg/QaqXyF7DU2e8/uqc
hutp+S7pzt4F6cNGtSFiYsxHzJrOTOE5V2ouI66Xy/vQKysaORK/5kK06WkzoTMJ
XDF4R/sMKG0dn87lt4VSK1UCHS/Zp4QbkUGrfD/zLA0DiHjcSgACACD97ThQVX1N
iozz6VRI1l1N76+SQex+es72HCQWnUCTygbba0le+Ef5jsOG8p8henU9Hx+yJW2f
FkgtHngkCdYX6n9Y5lNTRgDFJYp+hj9TCnI3IX0DmGSzXMlAwkbAADKdJswCZUT1
5ToxeHQ9fpBsbd/ngk59hyrRGa21BqFRF+KpRGC8CoUkxtBfvAaivYoN2uy6VJEq
VfRDuQ032kg9UuI6tDDgRVIibiaWhz9WeMQ1F5g89Z/jZgXSvWTfbzy9+KUW/Ude
BTD5cTE/69Nu7+VpusYG34k/mjIVAMIfa5xh/x+Rz2Mcunp9qM9SRzWwlC6vaeWo
ErXaQmeuvcYijDL8zaNW797XrAmU2fi42RE08fJle6mZACYik6lf7AlDiuu4KyhL
u3GsJuno7OzgVtV6elyb8YCbhFv/9c8JH8GVyBx9wgfS/hCli3UYEgHgOzxAVY5L
JcxwbPrKTijHDWBJb9DfBGPkyBKk1eAxCZqLjz0DBeFkjowAFMnDKvDjUU/+on38
Sp2/EeXl+u9wqPTFgWS6zeNPppJ6uDHE/2CZknX1A0VVTUkysF57a65vVp112Noe
9KHwQqZF58b4ClGrlvLclojQmZInycjPHr5dAqSnNsrhyPKHjtPqyrxOOnJOBC0E
uVCvtN/4x+y4qR6QuEBJQcwRqWQ7MC6NEDZGo5khS2MmvjYcjPjo75Ua2aNAYodh
0BfqNRhHRf9bGsW5yDvAmlAm8kEB47NW1oyBN537mPC/lolR9ilvYiB63Or/TRV1
8wkd5fVvW1IX9ywOYEeR737WgSn4cUx3/XZTfPzGyHfX+QIhD/8DmR354Jdi01su
+BG+Wa5pF8z3Hx/eL3JGmvCqbkpWd6Lv/Z6ew3miAeAvZGoUarbwZGB1QpLyrGgu
TNOTUehgo3gZUrz2/tIAXCSjGzUNGiUQraMAsqoosoCzBUoa2eT2HLNlAaQ58wZl
7hdGPPotuDFfMxNiImu2GfJedVTTgTnGT4JR9lcufI62LtnDu/pgVDvdo7D6gHV4
sySjrmEvrzd0ntzPfIJT8XE90RzD4gyYChje3Lhu4KB/ZDxcXvy4+iZKtwBkL8mG
4nPhSIIme3jk+OiA8nWoe4lkB+J9jxfYcQz2pWoVoou2y0WC58p626fnN0S4bG4P
NCwjlSTyOLHtxlD827e6/Has2XW+yJYvkPhKmk+p+sDCUVjxwq5hNDL7VCLuSV/w
/zq1bWmKWPir/f2UXoY+M7tryLoaNesE1UIPw+NRNSeKTHbG6HF3H7Hr+4KNbKWx
adsXaMJaBBiq14q7qcdwKLVvFU71gQYIbwsTBxBbM2kjEdD2Sl/glgbBehkCCH//
tlh4QNJj2OL/mzbG7fwl+YwJ7MdlfVtafwSQh5MlK8M3fTo7uHDtPASC8odQVNSs
fdCTfnQ2PM1IiIGFGdCCySfw2jC0gvpy6tY3V4qJ8HXau1itq6WEfexApPDcQAx2
MWJKyL2aAajO5O+4HsHAUv5p0F+SpVR3Md3Zd3o3k3c+Bl+3YlBsQTfxMW2xPls9
ohiJcAkEbPsPmwZXb8u61D9zB/BfevBN0OkK0toq00wEnxBxQUvA/QdEGCUXuryc
mIhffeRyDsWC/tvpXQvEXjuqO0I1Ms9Nk+g0DbeD3SUSBBwiLD7tiFNDUUgH/5sw
ic7AKGAiOXXVmreTGcYMVIeFOTy5fA/7IDyiUZnXzWZBLveaNNKF8kxCtp9n1MYA
BJRntSy+2ygmrRCx7CY28gXRv7UPZUXhGySLxkbfqH9Zbv04WjARAZ/VFnKWPidf
PEJVDnEEjxi3kInM5/W4IOMRf4kzAdroCAPAHZ/uAGSZ8jrRgtuNMTIo2XUQqh1p
6PC7fvIs7SXexhMGKcn1xArgPR6ljC52v88in+k+IfbJteJvkKhQsQ6DNaA9/qsH
2623ybwDyc9UNnXC5uZf2bDaoAJzdczlWV4PsYOBoW8nNMGtepgZz2EyIUW2Ah1S
i4ePTEqNRHQrTkCFFqavp1Kx71rGyZd0v9qbjlEhb0aDr36gLnAjpxj0pqYCcns3
mZcX6I9QX/++ki+MRx7GwLftufqgn+8rzSVQXQYhnzZSj3u+nn4zI+Pf0JNbJko3
sK3Idi8MRp2iEnvk2LH/KkxDCWfPL8YLYdlEolxmPBTJElbt0jPWSDTN/IW3IVj+
soyQK+RaDCOKb+zZoD+dYz2WSvhyRU1rsTl3+F8GH1qajr3dytESltwsh4yJHV7N
fWuwFHf4giSbnMpxLGPAzQt66SeWQybcqgtS1ADn+gmtJzX0n0AE86ZLptsxe9is
IZFPl4tWW146Iar5XZUb+J794EOk1llP0C/1ixPQvP4MjbRQTq9epZp4e4CQz7fL
56bDXUmxbMNP1ADpKoHDX+NA5aHiOXFdAnMzQYqerUdFhQA2FepOLx4BQenOdQ5y
roxReBELYG9dPd4nlTaD00x4IHJKmsx6fdMg0OLTDqCMCn52/6UPYqoePjk27M0B
tJkimJHmytAWbSh4vneKMydYMvRY77FLB9ALUPR42MJIqLLZbsoqE4RwlVMPpp2Z
tCD9GvyjhTO78ER/ps7fe0WOx3RFp8hmfKoeJqYJyFJsXSzE7jl3nc9Wz3eewyhg
VyIJL1XCzxwdVOS6jkSsqMLcApzID0QrioXXam4lNCRfSR9xx3RxIp00UK01Dh+T
3KlAAFTDwO4ofTiE3BDX+2ZrzVz1plumLH0uoV1P3V35u/HzoR84f8iyoPxOlGGs
jFZ2QvTuPrOXdhWQNAzRD3cJw+bVDvbgySoe8JM0R2Ib3qlMUlSBJRzG6lrjd3L4
QH424oW+HiMfD/58I+fASFgTrMxlEHj518V2kEvLzGQ7h31cAHXoemC0tdk0O7oc
ZhE53sawOPKeCAnoqPF0duaIY0eEK2VMa6Q/nvY2eIuww9o8VDqotmrn4Djvw6u/
UOKyEep38SiO7LCepRmdfAwh6Nl9NtLHPYZGqOEskcM8p7ULNu1ZZApphVm7TcVN
eItgqMjQX4Oka6fABzXZvrV8/X+ETUVJjkna3t6VkDW+G3ArBTY7GGEW1TuqIbTj
hsw0pdnj9M6LnyzvVNTbheDRXiLn8gkH9gEtSYfMj6Gwtbst2CTtPFQDjn8Pijkh
0SgbmjnPMFkNvfEhpG5IIaJ3fizZ9FoIXcaGMbUfbAij/iQlG6+YP25bx717pNuT
GPXWu1EiE8iaZ6Ksnu9o4Ul44a0lUdElex5HvZtVlXLVlxL+1yxrv65TE9vmIao2
Jw66WOPUqj9ooZ68rBLurywxf0p2aA8gIPHAjI7lbD4bN4iZqe5T1TJz2xHPpJaZ
a1uBVc01WE0xkjbBbQifSRHd5xpnqvapQkGxjHKrmJKVNHa5nUFBheTEd5ZQHL4K
AH1d+hSGO49hXlr0UNIEFHmZLdWuufIFS0o1Hj/lSQyUcfeAl4B9fB3g4ePjadsi
KiLPiMmuWobBb1CqKxo4KnY7QVs8mKdctVLopB1GdwXerfLgxBy60h8JY9E0uN4f
zAIQRJPYIamBiv9rAHyyUnvlslMQUSTDWLPukyXM79Z01wptN29/O03bejhtBJ3A
IRAPCBEj9zyjbqbB6+Kvy0qNGeIswMrdlwOz/EIIs4Ax7QTA9T36SDOzP1dJ7rKA
xBAJbShbN+Le+2g/ba8NJOlEtnjzZkNQBXp430Snsk4T5uA/je+V19SBZQ+/f5UN
F88H1Y/MEWjvm66tv9yqEfWM1Y4ZFKAuQXW21LGMQ4ZWP+J/VuFTZwA1qFBPUdDl
RCCiyx9mlpTTzgDrAuJdF8pta42SgPrGqIm42z0dgiGDBfEwrWB22WhgXSIfDYca
w73grAQxPSSg41I5Ytrvfu2meDo7pW7+mKBgGvQtDH1y68Uagf6FfItcvMAkvJn2
7ux4eM7zha0zpjoeBazaxlmzwQap8MQXeBH3v/jLtYR7Bby3EB8+EkbOJhiPffoj
jc5pEc7F5sXf0FBi2gC21DkuH8CJb9Dpw9fvRpf++S006CGKZf04eqowa86zO5xX
WbpWybpUdHdnP6FZ/JSvF283/2CDYWAkP7vi2sW4bqILfVnx7JxKd/EltsDpYV9s
4W2fc59nltyBT6nYYwnvJSh56pJk+BIzOksGDkSD4Z6mfk6eYTUgC9rXarNgQ6bM
eSwatJTU4otiRjNdARgg0rWU1cIcHg5L2HnyJTjOWdHzWS5piiLIsvXgRcF0r78c
ShsgTVS4KB4sLnVrJZnzB4IYuxOntjqByHzIe+9jr2L0C4IDHv1Tus3Vq2fDL+kB
PhqtnHcR0TIXvBse3TUkRoJc/I1o5uAScOKBWqCeRl3H65nlou+yWlN23kMOcuT3
NY5BQN/Uu3QJrFISU+JYCWLqd5z9S8VtNUOmaA/VDto7ynHy77yqO/2KP8X4N0nJ
AQwmehw/k55czPKoTw07REBk1wJyI289G5U0NAJSGaV2vCh6BinE6VqCnAbJ5hRJ
e3tEfVc1G7XolTJNmWcZgfAkMHqHmtXHkrG1yPuAE7++ISaLGY2kDOSmG1Z3bw+7
cunJb3QoDO3K/+O5jM1PuXKxeSkqqqmASu2YbwAqZYY5qGM8KLHdXK2Ihf8c4SYF
shPLwSzZC/IUnRjYzOnp+9ocHscASGSXIBwup5Bh95BjESHu+2mYZgHqhX4WlTTo
uBLbd/flkxpPsjKKvXVI8GckGmRAvQ/4clEk2bzLAJSoZa3yuKqyZfkc+Sdcl7eX
RySGSFkiO7pvJxPSjH7mAA1QpWXK5PS6f4diWMK4YK/WWVlI1qqc9HImSpLP5mBx
Eu1XblM34scJ+uR+wv1FjYqk+bwnNSiAUhunEJi2ITqmcmg8RHC4YVyJr63U/E47
xR4B3Id/mB/QIhrH5w3qXzCbOreldVT7BXTWV6VnAzwU4p01hVtrXoYl2JGSk5Tu
rHZEACEUJZMknjMPxWj5NB4PsmDuthniCkxfkZ82AIjPVf6SZd99eGjBvznP5Ypa
qsQ4Z8JpAWKsGQYNHECGpZGL2y0SXrv2yzYgnTEDT/CUfQrx7XQHHm3k1Uuz6Qba
ATac7OgdCjhqeYEIoY3WJ99HEbKLXo1w02z/YexT3lJBxYfPEmdkCj0WTzdsCnz4
qouaWAk+5X8JMAF6cUSQFNhmUW20LJp2gsnn0NP3UY2uuGJia+OQ/ZHs1v0Ki9ia
3l8R0SeROQFK/WHUfjZyO9PjsBSHV9OTkgZAPTaF6nGqLEYnk+IarfVgGvZm8ZAG
5PqnOVLWmfYj5UjiEnMOkpmWyjX+CjzpBdsufqAYiST8FItm4xl8PhOMrXSWq+EZ
D1kxO5csSc5ik511OKnKNEW5SVqG95+2+nhEmg7iixGfOS99wB6nQ/f3f7yVSWL8
unLdI8s1EbjSXHVsvyVweChkYRpe2+0XRaA566OoCUxyCEPw8A+Zuk6O2C/Gy8kT
Doha3EQ6txOqil36v0/8UorUZfrXgpecgbJkrk5Npt8zD7Y+Kwqjx3tLK5m5VeSE
vGSATmi465n/kLiGkRyR21Ptqrnxup5Ou78RLt61mai/+UyKgO9x0oRwHKJvfC8+
qIORmtOvSQzOZ2we0vo7mWiIWuxgLN/qW/iz+feYH7KVbuL9FUn+Xnzz2+eWeqCM
y0Fa1hcsTKfafE5THvNjZHGyRPX7mkpwB/T4/Kl15QnnQ6ptn02O7WfeUiUnpWvk
oNBB9wdyFj/c58SMGTHRdf+mppqPN9dj+g67VSG+4eEj7cIMwDi/BlqPrdilHNm6
YbRyaI3BBOc/GcsZXNjfijb80jHDcfki0zncVScsVJbU4jPOKc1IR3Kxe5YO5d5h
9bYXSPJg5848JihpN5SKihxEIX+k6b6aP+QnNk+29qRcXvPFtYSpbKvrVzfDjfNV
ViItnNX1GcNThRxaHXOPbkHxoynnSII5A7CoZN4aegMqbAKr59tMILwmP4yppth7
R5eSim/GS3AhU00uBDaF4Ge09XmhpvPYooPGMhx/LaX3Le9zG3Y0UoxsU9/cdpsX
PgFujldgLnSVs+Uzskl6gGtT8NLhmS5lieyQ2aWGPClB+aVmLb8EhKuG0vvgLM6J
+Hzn93eexsHmmZUx1zOmA1xn9tZg/qGfU/OpL3reYq6tlHlvfQlYSCFYo3kTrAKm
nVlkCEhO3I9Pe2MOA//AFT//v9qKHdbnSNzzpQXtW6aqjsV0UvzK2dgHJv+n+uNp
eGPTp7aIA8pjjKuqgMIidVRoX5pRi986YCq4LxqBd6kWhvY4GNk5C3gUQcnfi6UP
PKwTqrKn4XtKzoG6o6DRJThOm6ac1B2wLgBZH47SZZqtk+kTNFbq/VGZpW1vk4yv
h97ufftuCjGEUdVlmIYqRuZXFYrvYmQhwGEOLaEAA0j2aVYiQtwa/jRiHIkyC8ct
WO6LCz33t/Bt9e1iQdFNsPNy9rsTM+aJtkEU6TRAVBsi4S9uu+CZeOwkKHGzwlTj
lap0l+08sIf1k8IDo/5qBr91s2KlG2mrnPJfryEt6w+4wHeCmlbkduoNiDkEuFMr
1Jbn3NAKpM8wbjpUsCjGtOddsEHMQnFOa6wz6jYzR6MztpXBEg2Q8IL7H34xECfJ
lOvVJwJx+cqgOsyi352IxtYTZeBe2RhCJj7zaLqoJi62+osC3yqqb1q5HSOj2qDy
kO16sjQkMOZmusGk3LwdUdssTJ7gswvxQuBWBhdn8A4VT+jSyTrR3TgwDHFD6/Fo
ww6vud2W8YB/C7Uyr7BJh8YqhIFIdUerWA9okdsoPmJ2JkXsKhuW7CROzR7OeUGH
9Pihg6FRtfL0jokpzSqJNJWQcELGflsjluiTOX9ysSTVdWMXzodD75Lt4UlnYB+G
EzKlqJE+LNngkZcstYFp8Nlx0nB2ZXiw0qsfN0Iov/bc7NdpKQ+bnQ/rm78sNk42
VRj8bdLCAm8cdvu+i3tu8rBvawV3td3CbPT9elCJVQWj8o/lb5QsjBpvwP/zeojK
nrxOi4zJPBA8wR+iUayE/YR+k6elMBAWM10cUIDmNaQxsJ3tgw5kVGHjCmNAA8M8
l97UQra6RCyxpvdefUzGatZPcRJ88aKvzER7sZKr3a3vY1kUvg0Xd1DUJIMLOIxg
kolSdUqim0UduNzD2FfvkQWWwVC8PYwfl2OmBDpJaTes6mDIYn2F3NdGGO1FNPem
5XQR35uwTDtjiXjgmw2Hcpp+46d0fvnft0yDOL2bu2uCW5n3jt5nHeob/kcbWECc
gULDtt/J2aPRgHWhuu3rB8j9WPT2nq/+vBp0dUUBQiUx3kG1ePtLLBUGOqgKneeq
TqEST8L2j4GNswoGSth9X1GV7w8VBBpjKSmhoNt1JOp26PneS2O9knaiC8a/8wTU
f+dXgMV1EoRirg4GRQOWShL9T+QZ+HuT0MRQTutVbfvGH1CN4G572IpUKxGdQ/4/
3e9AJSAza/3Lnioq7SPb/WRU3SLFyHEQLBzQQlsLIdEDROh7lhH7cXFsda2gyakI
aeeDJEQqJDYVmn0/VGWG2opZ8/mmXdSiQugqkGGQFzn4+X5/AXB8hdSFJyWIoeaj
wxbSUjgXGKl2VC1F8rdx47ZFt/eD3PxE0YuQmK7aZHrn4lXtoChHO7HQmvXKJlES
GuE8pBuMZCmAvO+2F03RieHZvjVkIT55DlWCcovk+7cbRyNc7DRFqHjvUOG71SeK
oghE8OB2rV0BEjShdlKPI365LHiLkoyGrjwastxnQvGu5W0RDdoy/98/1B8eQdle
zGAgKQM6Qxy+kdphOB6eWirGnvbGnsE9WB3WQC4Tx06U9pU5TXoOoWHws/sz5uk5
Meh1zaFKxsJamVgxCRcNxGo7unPMktBsLCDTVxKMJZBxjXzbvLbQQZKOEvMhC0v8
LfB1MkqiAmHT4KmVizwncLTLwgQ9f6fcEoOiA7yKkNGigtR08feKrL8x4mkcpp3H
8eCZb+rSXOJZqdzuDXq5l5y9apamNQGvQ16hl7qu8mE7K7ZwoSf2pr5BfrxYeqq5
MGdQG+DMRpqhgaZ/t/29/84zNC+cXkU/Z0G9YFNNJhiqF/i6/t0m+0gO0rSpX4wP
izLOdeVActieERpmBInpr+Qh5IspaXBO/0/hHGJI+hMAwDnDu4dB69yIP6biff6T
utLJh2RiOXGfdlMOLYyEp7qEHqBSDlQDu6rI+EetfWkUqcXd2qZ6sDugyO4ZTB+Z
iT7rKCjUN/R89pdea7n/Es7drfu01O021bb20/NrP+fa/0D492xfMoVareGGAZcn
LhKe7RzVz/Zf7mSG3k2Lxu5m68AX7KQwJjIC2WVtti7BUhoQg1dYKI3P+FqCKnYV
g8BnEdGHBWBzg8Yd1cX5Y/ki5QEkg5JKDH+d8M+pg0i6I+TiesbO6300HWhAPlMl
Hm8+iQn95JdvM42xaalBOFqwAs6EEhgsPz8Q3moozVWhe6ReyT2thL03/cQGtkwg
qWEiZLoyWwoIhCE2tXMhxnJ4FRmBqfK3eKI0rmfMYfQ5gWgQCyMXXEvCujIbX/ud
XPR9mE81OHnZGHFuVTMcGoJZgppAyd7VL2NslsduN3QtZ0kkRv3YQON+ertO9PGv
kffzLA34GK15jtNtdvcseNBdRNbXUGB/zccYgimO9WSIC4x+UQHrZ+IkoVdJhACX
C5aHtPUrTw0aDmwXmASprKv9eyePGHcoVDF/IMqOTmNpB/ncGzw5MiNWiAx8Jhqb
dYP/FlygtUwF6tPWEdymHvSZG4/kdokCQxUOfpCruz1phSxxZ4NEOZ8K7TT1DB7o
N19IdzMmy5lzsvt2QV+2NZEEyvbgxK6wP7DIBQs62fp/JQ+DqPCEDaD7/aGOGSpb
hAjtf3p7NinzGadyQz+ecSHucAK5qlr4EAnX3Si8/1giSoYH8TNEx8gJAYhqihos
xWomtFxVzuAoRHIPRGeEYA67fXMwOkeq2nAcynC1/x7Ic3fe2hnWZm8w/+3wIOcp
dAzRTSzSbCDnTT+r4wIyjSY+bXHZNIwQtNjRaoupEn/NX2BKNJOawZqxyoBWC4w9
KzSp7okhWBwQAqXz/pgQmQcBjDlatEbLm7Xzo/dbTzRdPN8Rd+08w1QgM+q3mKj8
LcR9U471UnXFfUp7/L+eYy13nf69Zdc4OdPn6AaK1/Gs5AVwxZMKluSdQy0koJP5
1audP3q+qOX5/uecgazAnyvIU6S6IpbilUNR4x3keVXl2l22xurYQcSqZ/3MirCR
Erxd589Rdd+tlNyIZymjeV5kNwVz0g+qB9cWbnEooyp8imxKBtFdkKAXmmAx9qd5
I/TGdHqnFOXiZqlvsT9po9pRIRl63G24iF7w+5iF8lcYOMm5cdYjCSLeagum7WEo
3F8IE4177c6AiCLwlQO30CqH7w3j8VaV1DttUP4geonN8k0cS9xHh1MVwZDn3RHm
np5x7gffouZF86J7XnNxrk7AchAKY2Tkt+8v5WcBIt/4GM6xzYu4bo2/X0aaP/LS
bpyJCGXseaGdFVXpF3HpLLg26tiFH2ULJIg+yXXw/VNYGUcZHdhhKr530hHgb1xF
T+f8Ty5N15Q+Hp8pfZsK/hIkEIIJhsNTugacAyeIMQShYwBdVtzlLkTDGayKRrhs
YMxd5h8hfgs5jTrxOl8cylMVs+1ykhw7/v/pl0fiw56gAIyTyAPgugiBrUNJFME+
O3s52kzaiLDisabdrXVeEUSA/ML6u8IC0ciLgpj1Vqd0lrOMnPd4sKzXk3IVMbuH
N1pmU6Jg38Y0GP2twEzp9m2jaAc9+lUjfh5L4R0u+LKAI3uIVvQ3ZkORlLnDoqyc
DpN7C/iyeFU6bZws97t1ZDhrM+MujOlbEJ+bAwdZl8kmdpfL59xMUMocYCLNL/gf
BYJYPz9t3a66mXvxjt6QLQk0uY32DjXeOG+o0S8iTxA4ZMTtm38iLq6icDD4oCQ4
3py+YDHHmKt7ot1LuCTVE9ziPDnep9sI7srxXdQMJEDRs0jmBQ7hQIN8XnDnME71
Bv/Ci9rKGICnFeS6UrDVuEHjbVTAnCCOWgYjFWOd4CqtMjgcS/e2Hfr+F3C/5RZ/
8e3/Drs7l6+8MnL6aLl/Byoi3Bl0fAjllDxDuiUK3tn0mE3yVz1Y2UCFDkpHRYyT
gSJatNpj76FSjW68bqVw/5HAnoQvl8tBX9XVH6t5Qk1Cl8B2JhLfYoxsDZ10zXhG
NBZQlFPQoAcj1wwql2wYz2kjdD8R81Pxi3cvMKtBkhMkEOQo1zxOtAnHsJvk6OTi
Kt1T7/J4z43PQislxR775dwwKVouP5oqT48FWnXNhMOU9bORRBmlNGw+2VgNa9Ov
9pc0G9Ok8X0x6RtIuimX16WxhNRjkB0MXopuiE5K2SR1BwzsFyeM9H58ybACamj6
6noEgXCGbey4gf2u6YbtFoXeoiUwSmCvDyvp3H3ciIGf6c1sXM1kBIsFjYjsTWyt
11SZgxsIkH9wbB+6F4UTDi734xCPHUOGDssL/upHGvqXFpsnqALSJ/GsRdc7yUN1
QOfCSOpzDA8DMnmHZk0jE2a4BFxsWq+E3TbMsTfJBrUauDTLqzOnx2U9AUqUDEy5
LTVS34o8AVaKVODWEpoOuyLlBWAqIlNr45MOkWIIuFtcNzqwHcveADIfEWicOAZG
gVQKXuORToIzw7yTnltOyI+79CVzIOz+l4XT7wxJgyIHkYxGsMyvAEY9SRl2QKTS
gFp1STcKGQEibqBWH5xU28lK/kZEPJEhHnhX+z/cA7EelwC+/Yrbz2yZdFiD1LYW
rP0VNsfdcehdoDH1lue7mmC5lEOkw5/8vVjnptJ76vwp7Fq9Z5YoZih3d3avTNR6
D20UQ43cbakm0N7sfzrwDNF0iYUSlIBOXv1yn3DeCTB7PD44TGda7MPDAzqv92wJ
r11k8PJ2fkXNpbP0IAxRDcWTftV6ado/s9v68IZECeSwzyzhcKwXGf6YflSM5bVx
gwBDfRc7h1+DS+PvR/+XG3tPn3GLrhOuZuoA1saWjKa8XkE5sVO7GbnsV2skWU1c
BmvYdk25rN/rIl6cMJ2lio1zWor8Nm5bxXJZ+iqwvcIvfnVFLqMZ8dtFSrwIt3im
6d5HjQr6T+TF3YKfURWBP8r3mZsPAigG3YXgSRUqDsFU3VJfrNvYkVyNJ22dtyGH
B/Y0loYJTVdXaMlZsXZuNMA2zI1MK5B9eNK+K56IPHQHgreogCz0xf4O4Kke+qT+
8gQOfS9/1zg+aSKSgtyaLqC9V4EnLi1LxPKvEpJCreiXcHkwx0NV4H7h98YGtV9c
6u8ANbpLHt3YJM1wt2ABXj+EsXhY2lj/MkFzD5AolQhW7c4+yi+yS3t/SxRELmyI
AQ0xpWPoIWoAC+h6CaKxq6Z/3lIl2bM07TzVYE6La4kyMbYSlixuDhNLt40tAkZU
UZEU2BmirV/95/kwF51DQ/ocA/eQssEohUeyWB1p+736wbn9nANCoscLC/uNv2AU
y4iFX6qG+10/PGpEU5RCHk1FbFitG8vuXVAcMaxXeaxW9Tw+8/E74qWidlSrYDcA
acjcf1mfKdRGGZ6eN+rvG6CghqbZZGcuoMRostg3sliXIJMjpLgqOtjArGVZ3WHs
dSMk9mvd82pbB7Zh/bfv/bSFIubpZ4eCsalPEGVUHGyD4TwVbw8cIe+aQUjXUT3o
vkaCrVrldhFEzeSBCQre0sEWfEwHZn5nWSNhGoikGsIUGMuGkp3sqVz5YlyfJY9K
C/Y1AdWm6ISiJxvx1jwUeqX9SY2c/GcRq9wmGTmIgJ/J6BjtqJBIjSsdwfCPfcfB
n3aFc5x/6w51ksMxWgnhupokMoRzrbX8LHACBtTaTExVyAPIf0rlt7fHfyhpZ02L
tdiA7t+6M3eeyCNaI3tyXPQnOGYabKX2cCcdIcezYhOekQFnD4XsHBeLLKfjELmY
ZxQms8g82YHl+Nsiss3oRexeQH8xhYzt2hmA4dxEyU0VIVNSiKRsT8RDy8//L0zJ
jL5hoIy0pmgS9zONX3LkGaZQ1xtYX7zwJ46qY0PRL+7KPVSnZnifFJBU6KVwDSfT
SLGZyV5D771E0vh8EwfnoHwHFaH1kodK7Z1bGfS7oabOmysHgp6TFiCEzC2C4idO
J/xa9LQdT2Sxi1+x4ilXnv0UqiXo4t5Eojeb1Hnaw+64K/gHW8gNCpDV3KkzUkx9
/GQ4zBiOyLjrt7lGUFpAjHSxucHcwa+7Umbxx0JMeV8gTWkl0gJPfuQNK/4t8Xd7
qTrX5/wL+0bBWlxUHb2QH8avSwruzaZ+N+XkypyFcVcPJ8DjmGc4uaYFV04gYKFE
lLElgsYKhaxAd1BgyBr4DaRDff2UKgeNrV5/HuRtTJWJWdGUE2EdXGjzMFubA4qZ
7YTPZYeNSmjAjYT5p596etRJQLq04TdcTrBFrscnJ+/OSM/aGvhV3TXGRQrX2/4Q
jj8Hq0jtIjP7zyBomLb2KNRiTpeuq2oVcW6wSg+tEWfxnlPSPOx3AfpQL3jR/4zU
asrr63D0KRZXfDGGOMIDsYgBtIE+FijNwChjBmXYuHSwu5kuV5Aljc6GgZKPUE1E
dAuxjSeD6x5bAepXj8Qd0EeamHMTgwEiBLN21IxvLnEbYt9eI19ZTd5JtiaXxv0q
zMDFtC9hAP06q7MxxE86IYlwV3ANAqJ7ikmbRxAC4U4T/iI19poatPonQ/HjWcrZ
LkUUzY9+UPZbR4v336sWdc+B+s0PGObkD9dWByhv7vy5PGvvihkwDKDJuVHsQH4Z
am40xhsPDBmjnpYUrwd4d0IZzwL7N1de48nsWzt2yyeZ4QUncxX7TZMH44c/XsZ8
hvi4I5MrCYc7FRt+GiV0cQG/zrIXqHLTVAIofrgygBd8CPCzQuGo1Dkg/rNziRF/
h/Cj17HsHRCH8V92ZYxvWARCidFKJrd0J4jkKHidQyx5784eZo2Kb4s9ty3Azm1Y
YeHZ0Ec2i3r284UOQ9miBDaU6W5EmyFcHiLjAJcBFEWlLWvy1TpDdY5zGp1TuIOn
g0efZdHf5lNmMRBSuz0tq8sNDkziqYIsstjjrILljdXPy43PsQszQcoXIL/dgIc/
ZVusQBE8JkKExQaDdm+8l/5MXf7Gt9lG6UDkICGAy1sEkxdH+zj55wy/K98QPEsr
dKa/eDKgSOaDeNsZfUcX5n1UYSEcmx1DUYHQdMZsL4PT1UCyld6dLR0EqenTA1Ir
RbB9knJZ29Al/q5Huz7OLow2aFiSUmlUOHSAHZQuhcjXblcugfZZIEveep9vYBy8
Fr7kJWiLOpWJm1cNXC07L/TXH3zifdIm75tP6pIHj68FRbsNvqh3jGcMGBiAhY9P
yqHuY4LVOgEDWdq2g6ZwMGbKiWvQoABHmzOSQfqOuEl+kpmGFxk628bVk1C6cVAt
3564/RycCPzF2WJhUGRRSkuEac3CFXbeTmrnbWUl5UAWUbjiflNZ8+2cf7BIH5pJ
JviWHkl8w+40Jqi9lIeBp4QMeu5DVyE2xf2av8AGH1ynngqOyn5agGWRlcCDR2MQ
Pw5u6ZA3NxX2qecV/viYAzAFNDRHFdeS4mIdbS9SR5tOOHasgmpo7AKbu/vb13vb
gFcvXCaT8wmmxuPfSS0NpW2Ix1jnOmd8azCa06q8SShw6/tz17ZcACUVcbOjwxkx
wZ2GpFiem76VEHPM/1KvRgliraRdHiR0DyYofzblxEI3yi0haulc/lBPG5WJmFMQ
Smb1BziPbLVYHWlh/HULo5ROkOnt1FTtMhdpS6HCOs+FC1vFsFlvzCOnJcj9w50p
ht/cArrIS30slS5XfD5Au7BJkH5O17uZEcJ9HMWBfqdukVYrgBzRIx5kvzzGekUS
FTTSyGFEyaj9V004JajdmFfOvaCJ0oNFNI1m4axXbkrxpEb8D9NPb09PsEDZzToP
HhbRl27qczrjkuATiNogFWe+6rhFH4lfFB5IgXQGY8lfOk7ZoXJqXfnBjQYv093O
Gp8iPdU99eXOlh4HYuuu1edNjJclkmMmb07rgnG3blQp+Cs2SpAw45v5QVB/hODN
87kmRAvza97beVliHaBAZtcl7P7CLRedqMdIoJkw974QCBD6fYr368SsSw9Mk/2B
26BHMxz+7inv/A/DqAl1rRPqLONSGY5hBUiBfEOh4dUvKCkYdEUbdGwgs177j1jO
bTZz4rD1gsGTd8M9pBVE/LfkrByy9dh031bfkTy4uZx0savDZaxqi/UeCz1d2p1W
JMY9EIGBVo2Y7/pYOWfRtqQ6Fb8vKaCNP1DyBbbI3/LKAY0NIEfanXWUuLzvwQbm
wBXm23yoj/dcBwufASaC+ZZes+oZrqGAVGB51CNMhllyPux0NksMJUx/vtNtWwOo
dXdJZI7fd4V5o7VbmwhxQTE0eHzTD+xXDF02tYrA+CBeS4/qd90hurlssVUFqEbr
z2I2OqfsXOrkiwcF9p6KE471jZ0Lk9Yz8rW6eYycrhexp/Xw8Fx0bzrp5DgYMvCq
Du67HU/so0HALKQgmm6fdLHQBN1aKEzoUUCDJh9DCpdhyqGABWqp2g5q8Jr/BHfN
l+LVoWF8dr40oZn83dZBY3uHc0TVtlZe7LmFOn0ZpqiOxrcU22dbZU3BUvYmnfk5
1WQYwO3teYoct/DiXqm1y4SMQszkw75nd+F9L4JLudjoi1NOwJK5gqol3MEqhdwP
mqnSBuK2s/eju6NHjqSaNVmDZYIG9VDeeDENr9zlSjwRkfFGzHtm0AXCTYYljXcX
majnowik66SffFKEmooMPi5Y9uEA6i2qUtsSFZyp2Q1GM96TvYe3RheZYj8pb6Ia
MtJy6zcOFRQxx7JD6GaEqOkS6nY99Q4DkFr+ZWU/ZqZp9BzPTFx1rRrwHrKFhD7p
RF6HueBxGIYwT7S8DyAXmWK9xkHwN3jmBVXTm1zBBcUzAOvHQYKgT1BKyw1XmIhA
O7e44vueeZLT1b+eTXpcBqNnRRX/65oWcuqTAiTCqQAWToWz0j9ktsT3c9RKILnx
q8aixLbhqGITuuEDeiQmPsOdMgLeTCBmCl/8jqgk2KtFYnQQt58Eg1IxCVVJeNwd
NBLMek8ciB7dPtB0X9yHS0qO0HDF5wm0GMoUmwM/jjghVAZzl/XbCzZqojiDiWSL
tcuB/9rWxLARS9mtv2gzUK0SkqQOIxEAbDhv5aoG9JxBbaJ17vritPvpf3ZuWCQJ
FtWU1vifAdQdqT3gdusmTUccySODXr5hVrF9J5ZSkpX1pRtYtuit55EA2oMze1fH
ohMtf+bA86IiSZ0bOCrPr3p2FwKAY5pl9yahBErJLltRZ++hwAkW2gZ1fdjWKgtj
M4AqVUu+8GfWiJ4op9DWeKQQUp0RgZ0RPQlw0Xl1Ezk2ouMbmZeC3lD4F77/WLwB
mkl5K8o8D+i6/41JXuZly4KMCfIJGqUOMbZt4y1bZc1nLgxhjJRue1Ml9wH27hMT
734IuwK4pU0a8O6hDpmpK1ZlAxQK9Sd4z6UtvHoTR1E2GQ4Y6DtGdV3zpH4lhTQC
UWNupVdSF4NVvZYQxCWmSwdBw2cK76eRouVRrvRbDll4ryHFy8nqrbX5aL702N9/
sI07l3LiSIAKKtmHQHj59zSIEEMYsi15YSkeIE8+IRFfrDgaJf0qa1U2rkgQe3zb
EOPjARYhpciVVoim5j6pKSizVVUb3+l0H0/cQIG1JOv7MwS3bNAIPwTbP8Xuxmcq
sQ8cS7ikhariHiBSc1TEfZU2Hd+BaQdZlGkB4+Pf6W2Q3WQbvyabjqCJ9GcY3G6H
Cp5+G7aEiNEig7X5awjAoll0NLwSxXgG1oLhKZeLwsW/4TIpEWV1f2iUKrl4MeDc
E7M3C628Pa7ZPnpVdJGsdLFibL4MtlNDFmsF9/QruMRs68JOfP1K5zU+7eWNrLyY
3mvt4C6T+iglFzsdw1J/VMLk24nkjpo/9GgUDRTCpzACjmrvleVpDznR+ymPLCzn
gvZxgGNX/5jzxtcuwUdlTrRYWd6UG0ZenhB0y90juG5T+gWiPYfjZwjqP5SXvoEQ
A94azXl0itaxw7/V0v+djyfFEFgXZH4i0KpO1o15zGlIZYENw9NipZ6cdeSJ2dVq
z2X5P/xrxJzSpwU6AuRCdkDM0w2D27VRW3gxa84pEWTydc9PmX8y/iG9f4PAW26z
nYIw0Ugxoe8YppryIdvG2xz1Y2tc7tmUjNwxVlOYu4b+wNJRv63giUUu5oCF7EG0
oqk5lpKS31UZHI5KqSi0+xwT4ALQ1WIhgrVeshrsyZMVQ3ZSejlmUKpEMwcbAsN/
t9YlCearGgC1ULad2vqx2oVjM+zgD4RdxqnblcdIPVIe/FuFPFv8/+YkMm7ww7TU
pTdH9Qo48YzMcDQsZ1bFQK8HCc3AzXxk4b+YJwVIw9nDWE38cmJoP6htjRXKvp0c
RincfEMyhskfRXxAwuboek8gfXEw4PoLG463Sh3ZuuBfihH973gun7j+QEVbTYeN
rTFZcujiZlHqFyuX7496jrurg1EsG0He7gJj+HANCdADxw5OUWKj1KX/MBuZE+uN
Ku+ze0Xn3CAHYWiNnagNaXxucXByFm0+d1VqpsyCTLw5I41MoxjPg2FNUEHwSSta
A7+byqmBCQTERs63hlVvGraFn/L88/rHQCUrlbNX9Nbt/TGSbaSvBOQRMkIrvs7n
Q1i2daES5fooHAXGUAzZKr110ugugjWjcasJagBushBs2dIJTBa7EQt669UdRohU
q3sKkAiOZtL9LY94aL95lFFUSEsGPP6f0KBaov0BNC+r1Sdg6y1qY3vfZcJG4D9J
TMVWGqE8gunFsAzUF5xE6L3prKLSnW5obr3wLQwzKT4jAQJoppgdQBaekQTyqx5x
ZUs9N9Gc3kYktma6vTZRJRRubqvlW0W+TMv8/WRzq5Xfy31AwagsnGBAv9aVfusT
hm3dNidCZOy3UUgdFaywR/XyVLJyIQxc+iodAmtiSvu0Tzkoof7+AkZczbtoJE5j
0tbU9v8UEke9y6iGHPuLJZhbqUJRVX6jSGSsQnW/3xsP0p14HJ3Uhl0t/vmy1NSS
M1XT/hAL19Y5oNGH+Y8Jzrv6pQvMURrFlZQ8LUj3kPr0MqucWhzFYbf6l7YV8SRY
0KDVU9ggh/EkN6uJLi+PHrudRKGBxVKZksI2rk5i0LtV0hCu+kRT2ZHEF+XD5OHn
rgJysnxIc34MdI5cOnTavgO+bHGAWjpib+9cLNVLzEaAV78bYjKrjanJ1eSvMFdk
HCb2ha1OQmd+bFW45CKCTFf6mElrSqoE0sOiOQyaD8c3QFeNkwpr75vsqvYKRe6c
/7h3CUzvKA9jXG5PyQ1NmdRtvQMOGr9jKZ4PdAgwmeqXHSkmrDcsEm9rHpQKVg2y
bNgs4e6NEvBUU6Tn4wCi9d9Ibsy2nAFTQQFHoUNC5RqYCpnchS8bLY1epRrbQsU0
lH0Mm7QYnNNrzkLcIGZSjbL3SzArR9LExWGCvtC1dIEHMraPvYAIxpQVrFil4O4F
lvBm/bnOdyD4f7hnBDL44SpWN5q/mV/sEg2vruwS0iJ4WFJ3N2DAQtmYgXex6s4O
sWw/fbVRIq70ai1seJGqHHxOukleytEyMxub5D9Vnger2w7y+NwBQSxgsxmzQXXk
NVESKRsdaMh51wraLJvBSvJCe7y/BCJXN99XSl1T5OHRTQwqUoYkdeRnmJbJJ8GU
nrVJABF7JUrNX4tES0UvPnueCOtfGBgVdDnxKByGsHiebsKJS9KZE7+Sz+hQcVEy
HU4QMQ/tgH13aTk3KTJLA0RmhIYLmFUyFqCLOKt49GK5sU3h+KXQz9xGfzDYMBo9
RihJrU/894d6tHFps4M4+sqUSacxO8xT7QqWVQwJoyENy8eIoXg4Sqd8Bsc/0hB9
UtJHYYhsgk+hZBGyFmtZeSEWn+hiucxH3oUb2oKNZnUx2rRW56DeVAEvn6j9hlDq
SCgGOMzShB9dqqkGvCWJQrkfIiY0ARcmWdpz7Qj7IXBWG9xz0CjMC1QPyoYh9qc1
M+5K6uxL0VEW9CK+NdurvwaKb2b3u0/1rxzHHeCzgUF+mfv0yHVrl0UVvmSc9qlm
UpzpZQPJ1bNXCyO3ZpBHPmyuMRQC7taxqthJW5PHut5gL0a0h1m8O8wuElUQlDMi
3fsrF19BujxnundMFMg+RPdJbUvWJ7AzqrdM1HeUhOMdayykoyuH/LeG/cwyQk2Q
ZOqaYuMGxhFlm6wRAG8GgzrgsuEBW1RujRwMDvHm+CK6O7+vdHvtiYt3ba3IF3ia
tb9uZltrFZTx/8iJy0QsdLjXqgdIJ4OM7iUifOnQRVerJwYUr/dxqSjwM3uirQCO
oyZpRPmT9xYNkSXx4FGtH90pdfC2IxBQfEwWhDGzrhcpwuXWmtd94GlnLpdkgt/D
hGLvdBNcp7+RhJuzMBA+JTkE4I2FYmRy2lUa9S1Q1nIdNbQ/aoSClkBSrIllwiaU
H4eaFzQPJ8wxQAw1uu3olqqfDTCdi3/GNo4v7FhqlM0DyEYkwfFLriudVaUCdjvJ
7+JSEx6x80CUE3cnJvX41l197Jm+2ayz3U24iCCvn28m0TYSx4AY1L6KH0pkXYvO
zdtY7CewBtzVrk2FiNKu9bmY3PjjNzyXQc5zWXNVximVVJlBd3jvIBbTDfWuGXls
LYgAZE2ESi3CGz9wsv/PUXCe0mcQjY6gFMCG6C1845Z22cMGYrkSlr12pgsYDxg3
nweaTpg1AGkm84hcUFaK76nqvR7C/BAx2c7cgzhjaPasKodB3JSwxyUHj8KD/Unn
DY8URF8LJdRCITCCQeC2TwLGPox3wpZnj3XPCO6Z2x+GRz/Zu3TcdvdNvw3cH3bw
89tRXAKyPhnOpalp+1cQ7dvxapfhrS1seqtTqjFDYRlZ502aCKdH9LcKR8f9KfMP
3oVRPoQZBF4/ZIGqhLhINOpnFvbcxBQ/VHgJhiswRJdZFqU6GCvY/De6O0X1Wi5h
5GpMH9QpyU6IDHUW/i5b9cE5MZdnIByg/6BzNuug55YDbshrPV1bO3MSJIGKek/i
Y231QBiyaDdvVD8jKW6fwtgfdzL4QO3/Ie70kUdbT0kcxiUfVtb8VDh2R16su1SS
OmqejiXeicEYDwj0YkXWWvsH75Foe2ZATK6UCGDPpqlT7g5/xkM5Qf47jIn0S0wf
d78Ov+q7d45EC1J+dx6pGrz/ezEQKdJpxLJtIBQuhbNNkzpeqpGtVpKoUz/6pdwM
Vxgrf5Te/KpeQot0B5JsCJ7yU0gbbAWFQF67DRnlUIBGHauhzhgF4UwXZ8eqyEuN
nlDMCRODHz/AZTbCLhe3R+MztAlLGmFEjzaw7Q3/Xr5J8L3++HgqrYyUO+sXc7FH
6oU9owyHW+KrqQAvDdjL0hPrRFXMVmq/7IBSqjpxCPGXM4PELj+xR1WzEheGVjch
1u+1pm/wRu6UmgTTiTqiCYZptjfK5QLukdbaYP1Jo6mqPiCDrlONlZynmoR8x3hT
3wYnvvNikKQqk4j/vTwqR1iafHFwt0MPgnVIBXT4A2DgN5w1LsvVnPq5JLDU3GQx
uJy0IikplzhieYJokNcZflqRo1RcMrvsu9ONf/S8bO3YUiUo5GKoqaQwQQhCmOVj
tOG0LH/f843ptglBfFWdFaeD0iAfrpwkIY/nykf3c8njWK+cJhUzTQwWDYBCtTsv
M+yV7X/cCEiPrBSj8P7d0rG4KLztXAjVxBmdnT5zdVZP6P8LM7A2bmaoNTHjKfnQ
dAWtlaJRpv0bxbWLcj+eBPiB27lAidfgvyl8XIyjTwpJ9ityLELrEVN9PJELQowb
cY/Z1lrd4l690BbECok4cogYVTMq8D6417UNZy6W6cBZ0DXclfOlmiP8PC2mE5/X
jkK+WO4/ZvVNEGjwii0MYMUXIsTjIVj9TZ8YmQhsemsC/9+Oy1I35de9ejjqMWGI
F30le547pwOK2nTpd4WucCaeVYkk+XABrfhH9ubKE6hQjtc5nE9NfVmc1c8qzPE9
1NN/hM+P0fBdjkcb9FQOxpoIssThiP85gRjrsClfXSQF86RiIRF6Nrga2yR8OOhs
2CMoEKAVFda9JrZtVRPEB6pMt0v+FalIVsrUcDwareKPWDIPnoDS9wV2SAXLBXae
U/9sST1btdCkKu2TVckPLgPpD3dQtXJk7G9AdolSdYosH6piuushus4Gh1vAAzt7
0HM61TjQisFzcqZs/qHuNKu6qOlMyjEUobJpb/NmMc0DZ68B6ih12N3CTwQO6hp1
H2D3tZzADxVdY/LL+R33AhZhSP0C74mTxUtvYHy4yNLsgNNw2zXG5X9I1LnnmWVt
mgJrgUY3yw3yWDOozLStHYQT9i1DSWsAJWXFN5wo+h9kmrPnrlxoASEnRsSFq8og
JL6pBIVl3AVFDsQ9sdeywvojYcGDhGAqWr10WSnJf2x13kCyo9djugveTsEPuCnJ
14e9hRyzQjCS/PD5sHfb42jhH5sSD9c/aPBSHttBuecz3x0o7bfM7YQTvBS3y3ny
xBbLEqdUFwO6+yIMN7jTDa1RLUry1LNtyNmOU1pswmzpYEeamg4m9B8yViZU+VxV
pKkchKovFgE0UK/NJ6Bwku0BOvTU3O6Xk3VFeOTa69oW/UXS1E1nl++WPSxK2eq0
Q0NaUFM0jjNRvJMttD4Ozf/RRivB5YkT9xaV5YHSV0YfqZACWtc9giLQ72IyJ/tM
sX/PG+gXY28AyOApKcetwdAYz+ttiTfrr1gPth/N2vETz81QTsAgDowiw3Esv3gd
XsukkXgwFCjnClwFdc0EVrsGqiiXaP7OyP9KcxB1BZo/j2XPcIXGDcscwdBdpgB6
XXfIkNXc8LH6KOruXrANVIQ/G6BcOprB9TUteDMFH839T2jC1m/ERASZBTQlCwnA
JqxCAFoKdlj/4fDAcJ8LRHenps/mY2Q6x4MoUu2QchO/hTy6UkXMKP1VYYJ/p6RA
xlP8be/QeDzqGNlhh5So1y3V5V5QXB/vEH5GhTv//EkdpDxBOoR+qwRWz7Ejmhem
Lq+Q+GUz9Zw/z3T/JNXpezLMvlsN2Pn9zd+J7CFyQ4TF64IbD5dXmhE674cp0DaL
h1HzLe+zKfa4W/xU90b+oEpYD5rC1wIpcMP4blLff4hHsx5OChpNEvEI8z7XiXxi
dQ5aUpyu9fZKdXG33T1tTBjfCqfkYmMiFNAw048WLOYqIKeGxgGmiNWr95XzyB/4
eeyJYsYakmS04Q65I/bxvXBIQuNQujdy1R9S+TKHukkikYYHTMw8nRokmHDq+dhg
B8rSv0uroUrqJd1Ht73KVbcRHvYMcUFhohM+2x3AMU1beKrEanR0Y+eBemdG4ExM
r9N4vPmuAZPm43FGJwAW7nKuQsvq+vS7IgwhrAbcRq0PlmQD/ldCIK49rohNBwq3
KLmdy1PZDDJb6y7jrRB6AD4QG6SApRrz5d5vBXMvCdi3dwtsF5vU2zRviUiwGD6x
HSJRbrhgUW6VdEh5H7iOzgi6nR/mnIqsXnVXZqjFT0OXG38dzPr7PkURdIlTz9AP
5vWFXiFNX8mT0kUJNJ2umMCS4pPLk2PWdOdlrkLvszbPbHfz+yDo2MTfn5H+rYDi
qXRBRzc06BwTe2FatPNZS8MjPSF2L5BKNuMb0RIk5SXvHBFJSSBNQEw1iKWEF3rs
Q1eD4i8xfVjvtqSw6AwIfHjgd5gBXUumZkyWlUl7h5LXLCIUxnJqExXD+DTXfs/l
H1YdxqnCKxE/5CTYrfkQ+xlH+dwSdiyrEkiTowF7jV6aVm3j5znf7/ghT5HAyw7z
cTfOF0Rv93iJ9gNrU+0gE2dRlxSi6dykinScdkX4YrnUA06UCjoF6KEpxIlLyWng
o7ftivqpbJQDTP4OCYFP9CSVp3lubh4Q85Xca8d02kzabDiEbUhPqeiRdk6k7Nxv
gz5Z2wDFMS/lJ/n5z3k+jfHkvtnRDCG4tNM89iyRW65rlWLBIsIh6ULio+zs1owx
u+Uc9PKeuGPbZKH9675S1nr4+G5KdtbcJKJJGaGmg896QJD5WRBJWc98cQek57Yw
/j2TFjR1eylr8wmjSm4xW58uLlud676LrsBs+6NsBAHTIAA/Txwi+tlqu+La5ZDN
EaGB5BSNd0D5mFzbtIIsG9jl7aAn8LbyT2OumgTUDXsVI+OU8P+s4TlWyTjml4B7
bzDb8uBxnRsJIJxY8/waD1WCtaNjYwVj3nsqmNQIsVLcsaadDCd2LhvTCOaPSoEr
AavXVT6DwbhXYDS409JPuznI1tRhTxM8kaQCRDW7bNJiEh1Wl7ALfg78y1A5trhf
GL9oRCFSgsusnz4Ls3TyIbtZWTKbL/aBIysmUOmLgpXDZpWpcwO1xEfYwm4Ibdgt
phypiWGYNCh71pE3XnEvLRKRkDEjQEzJT/mBj++Alf6+bydlR44/U3cRx2l+40Rq
QBm6W2YOaPfqPOwfeePAJZPFYdfFgPL/1Q3Yi6YCz3r9DhhIiml/IZPTxrV1297M
kuZj4KbWWWjpVyC8UuX5WU26DqirQyCpoBpyApoT+gb57PVj7to/wJG/4EgrtaeL
jrO8kYIZXGhLsxY33FkwD9ehaxc6l7DuLrYboelmAdz2lSOfLYd+KFeYn709gW1A
WLeJgRf/93+inqMP8AyupAwxr24Hqbop78hSsqPGFyMCIvAy44jJgFsq+YiUxcNA
+OeH+rQXJcvGKxA+gxTxeRDALusCUNd2XVw8suAHFzwovE33M9IswR7GhUf/ZYE4
dw9FmqS0gBFGXchQObnwqoCvubTjgeJ4JUU2KbAwp6gQqMqtWRXKAZZdf5IjPUHh
154AmXYJYQG64FRLbj0Bb/XuzN3ZxvSmWCsDsNofIiCt8nGg5MjtYZOY9lMJCu3N
k2900VjCEiMdjCISqjKEgqONWo3RkIpp9I6JhpI3l7sDZIlclnJGzhgfV0ERp8fW
01kbggZBOOzMQ0HN2PZwb2zUbnqk5ibpGMI3nu+bP3XeRhfn6Nlld7vaJXXPvOBI
aO6QZcK01zdi2fzJLUqAgIgaNsjRpRAAAodS1+FjLTlfXq/zdMpvl2E6dUd252z/
H+MPahgSG8Oa0sXUKtctoCQ3g7ro6c3RpzAyqo1pZeOnw1V21zZZ71IPXQZDspoZ
JomdSrh0nuhUZJNJIC6xGTkRi6hoMG0CQXWBuvVmytT7ilC1x0wqQ27WNkqlfN9t
7KoIb1qfr8r5P433irnZ/ym4o6VpIarJb7IdvH+8SdViR5btzR5ZXB5DG7edxzWo
4RAjIjgoy6Ss7pgdOfvi9C4B8osPRVC/pHJi2FJAcemi9JHiRFg09JmmJGQ+3TLk
E+sZdWreJgwSKpjTeYTKR20iMoxvSppE0ZCwXkf+tC8tJiHK7sxGGJ01ZCRqKYIu
KVJbZbblj2bkmWfl0BQTSxQdW6B+SV6A6pex/nbLYoXjj9h/IXhUlQvg8CSa13gG
Zza0fcxMHQacM+rtDWM4jzgYQrI12PhBO00i2gdjLM5kW0aULW/rwMcKWVw4GzxL
H6WP6HaTyBzZ3MEkadYWRuwO8iHbRggpggEFZw8GRdkbe3QmwV4D62jQW0HcBpdS
WhrPm3y7BXgSY0hYQY/rKHDobJyGBupsYml1FWkor+XF1SJzr3UN4MVEH7rjK3jl
M3d4iHC5y2BZMEqfYzVEwn/4tTGfAYaG9YkwJ173oYxI+rLZhCXURynVKmcj8Ygq
3Ie65EALd61UGie2Phy0ZC2gkGgAw/SlB4vcSqwVGT9giSCgffREl00mnmlC7Ux4
QFWFBgfwYXc3BedRPpnW7lM6MyEedNXw4VC/aM2F6HWK4J0fZ8K+chNrYe4S0YVh
7DK9FxbGLVSlNHU2lUGglh5up4n0ce/qpRhX6f6waGJkbNr6dEnL6wUmUri7Gou4
OMLw5eoVmXudwvCooU1i8XRWHtUAzeuKUt4KYRuddPsPvf8Sn1lfRtcO0oE5RhNj
jdOf32KTtdldlRq3jTiAEFC8IH4kj20SgbtSQeW8G4QcsNKAQQseVBGtRNboXpvO
rOSohy/NyStcLaULqU8ZGteeu8CGS5iHBBSqc7plKio6/BriLeKSP39j08uZTnau
06BEuxAVcS8opNXkws6WSFSqFh8xlmTXgggxDtNYo8eepl60n/vDhmdAtWpuj9DK
FrLJkCtbytpUDn4F4NVygnQnhajo/JDdEC3WFUe6w8apDtDsV3njqhOYIzZDOI6m
PY/R/5Og30ofD4C/+IgiWN2dFqKPeztFNDCWzieUSKIjpqjDVCIcq3OqubLaLzRv
AwiZf1Ccj2YyWxvqQUL23BEZYG7juramkO0TMaPAX1vT7iQBMc1g82dWa7pkz5Ue
Asr9ZrT+BMfA7opAzzclYJgOxB4abe9lGG63isXCifQ/9z9c4E0Yc1U/UB6YAg/e
9QxTevbRJQvHgg2P/ttEOr1LC76KtF5dr2O7fkIXXYeCIDvifwTEerjlyebUIcni
Ni6PIKakJEePv3XMo23AXXSZ5Qwc/6EAdwXDhIxGpE3CvbBfLDhbT8JNrv54s2dh
j/acdPitEgtdz2bjnr4HAju4fDwuHdgTq0rOQ54IHScppMKlQtLPC5c0clHgOGwj
M+2bnuWspmrRn1O09PpSPNEZrKU0iz9QX+jrcpA4YBKdP5YcmQGAE7DYXbJ4nvK1
5qGaSPcDDKiib5cYqO+yNq+1dAdXIr1dB+aiaqyi/qOTNHU+dh0fZL+Tu6kjGAH0
arCen+SSTSRmBkCoM7frJEyZ507cOoMhjJYQoY1U3ZS+RzHdOdJWFfOgsxONhF9+
U/YcsldXSCMHypsB/RKiJXbwNrW4wKNgc0ZfOOzC8o4PVeubdEXBvzbzHFBh3GO0
nOdIqVkAleXRJAOuKj3nv+NRWj9i1NEF0pS9Lkf7NdyoqVuz8ZnZzGOmwJky+YPh
waLdwEmnubfkqh9j5dbYwgv33E9q8X34bCGsfXX090Nfu06g01/EP4/fu/d3x1ds
hmkQHRb7eCRZ1dWiHSvQkWyZjYYnlnpcWGFUFjP4jc6AmCKf+EqJd08BS3k1FTkU
vWhccTfLxe1jSREV/JLU+6TJ9eA1Jg3gpiaWY+sq1AIGvBIlyOJC+MjR3FlzkECN
JuAM4ImTr15gGhTgUz0AK6vvCa8J5+Z3mGDxGUfgCnXN32LNy7fOns83VwN1twQ0
PEQY9tcGJTslngzZnnUpnFriNKIKICFnwrVi8FYcFeheXimHjrJpn609VrFZTY1u
Z09ReHcE8a+E5iVYH6dlvJ967eJk/13Cj9syiKhOo+0bGnMDbfQG1nW/5qtlq43K
XW8MGMk8ft+rSI0NBkS+N8sJkh3Ll02zgpxA3Jx6uL4VYldSvfn4T7ItDtTdkKHW
UY5Hc/WcZBjB5mkhY/EU5526ACJkTz3kzqBgaxWEzoIg2mR0O0/4492giunIpBc+
wkDg+n6FPdj4aJ97iDm8X0GhaTavZFu+EGt4MUHg8CI6j1nHP4OKmf0wjx+NQPGR
JgmZZa2RqYSm75OXSn3yfogNV6PpUQC5zlxyRHuuazuQ1ECazvzQb4EEWSbn/CWM
1A0EPigyECvXzHzTSA6reP4WjIlu93TCqd6OlmPaBOu/ofYQKAyh5x+PcMFse7Tc
KFU9BCK4AdEmwUEIMUBOL3MwTLtwtySO8KrBbqOE5PHKutjEfSizB054MCYr4HGU
l1JaSK6pYXiDudLB1t+PxcramZRwJLA25Hzzr79g6smvbQLChRIaCIIrRKCDiVX/
CTslwFza0rxWgtieCWeG3nvwJACGgFDpXwb9AdEgR3K1+GPPVbfIY3Ed3PqwXdXB
8MpQmIAdHj7VyAnqmOSN5VPhrsuwqky5uVeOmwfajZkLhhd/BGRM7W8CrOp72GhX
hjgBJ00a2RN2TyWsSNAvmW0ZcSb9WgZx+iqKXO3GPzK0E753hcwPOKCYjlZ1xpCe
bNrvn5nBva+1RuFh1QR40mVacZMeRf8f/GLwXx5bu6cnwBzhbrp2BYCP8JaStjdU
d6IhqfMfOSCg3HLWG2Ejw6gOUTkkZUOee/6B4Nqk2nQGZA22cu4udP24X7S8W+K6
XqNNLTAK5kEaDEzHHKf8R1E/bJ/AnQg6kZ22GqF26Y1JzjNH84OYbvtqt1rfIQao
Wo/Iu+lWMKyZ50DKPLkqgwdszG4gcnJjNk8t166qwTePvPy1tDSYMeyGgIeDGdKN
IYlTRe4U6Ax+b3feuKSI0qGjgUomKJre63GmQL7B3GwcUl6hRXfaWwN+rrg1Z5nu
L8H/xfmJGfsJ06AUuZJeNXQkNkSO59ycPswz3+WDSpxohAIDPuuYZorVrzItBtTx
AswppabA5ypbds6oA7krHRek7qOmGegT4Bhq9MIv9MLEJj018xrp1K4p8k6e3nJ8
O4PvFaJ5t9hQqtEADDHQrd4TD71HhRb5iVt4Af0AHjFzma/7WdwrBRK+ANP+6Fn2
6IF63z8UHYfxY5Cj8JcFTu6jH7HOzokEbhfKQkydgM9Gyu7EjstN54UVMRix+Om5
HxZO8Pg2Me9Iq9AKcar+ParUwcdQEpMx+CT+dFaAO66Bu+G9qcFqetjytCwHDTfC
m1SmrYRxbphcH/K0+p4dAqa8NWYvbDhroKPYs80ZNRDcF1dMZZMzNNBD9dEIZqqG
M/DfhqrzNPT+OA9jbBRLplR1LnFihNlqIxBasEbCZwMRk5jyLJrV5sWPWgeTw+sA
MoniPsz9TXckOAUVTJB1oB9owOcf9yA/w9ZhBH5X7pWx2MY7Jzbi5cVlH6+WylJI
YL2R8P6VbCHQpNqXvDNFs8spxsjZVFT6zgdy9ighg7zlYffdiA2R0fTYylXwlc5J
m2OXPL6BA15+rP2jJbccVDp9Ylu3vpXK0wkN7RqwhFYvmKADLNGjwDnKj1sIJG03
1I3UXO5Ljl78A8fOEUjwpJY190Eo696hP6JIpB5om18Sye354bx8YdM2v7eFKzBy
8BUXQLs1Tepndb03wC8o5kTi50KMO4RfZyeslzzFKEFjTlOfUg1PXSNsgq1kcwnR
p6UwFEX3disVA1rfUB6BqAX4sOBBNvmEiVPV1tIDFGp2g7EwMyhJb0NCPvGI1n/H
nVQwhnMrEFouNmcKSxIoya2jGCaGjvB4sbNSRF+dKoAv6VpQoKnA0XsRjwdS/S0x
deBgraW7TcasWdHnYZhTbBDLKk8KPmE2vBNj6tEuq79uF8/nkrewWVfvuKBa5ho+
NuzhkveZtACtbU+j0CuYcVqTSGh1Zo4VAHsprQtPVuFaa8yM91vjHhhRIF4EIjmJ
FqFEVb6SyqxFhU9FvKZdCEC79PTHwbLrVCvr9A727xA+LU1PLfbDdCY1Tv3qPJa/
03T3G6U0XfbN+BdTRwVwQcyJEhzkoVsbUoF5urZuBwK6KMr+vebMu1rE93R9M60r
PW+p5cYFIZdRgVFuYjcBGb+6DxTiIyJDoz/f1JZ5ExGvSyG2x86qtoVEGb8pv34Y
zSv6aO6LAIG9kZouvN2kHbCtTYWNHiMrhcKC50to9dZ72Rnld3eNuFNgOEEg0PDT
V7+0u/k7kKknW7XJA4472E/iQWe7VTPgDgVWo9vJQ/YXSx2dPgOrmXy3LIYRWTd0
SURJHSieuPHxCX4A3Oqp/so7vYwNoXdGH7oVI5XxIeJ1kmDR0ftz3+zDxnjz5OUp
OLwHmaEpwWAzQIPZR5uojKEUD0u216+pi1a30pMyuyttaXXZIVJyvD6yRi7/qOXC
oxnMmqKWNo6aoS1sbeuWfECaVoX2yWXl0DXGc8Vb9d00bhxMb6E424rAJsS84QLc
f4+CMFO7RAMHalwvVX74L0pIaPrBuGvxCiMUzkuqWRkzbODHuyxXYVT4koDg8mgZ
+bZy6FKrJm7cif8YVDywn7SNwNlhooMDWe3nCSzLMrs7QkGRf6A+3NYAY70tJ4w0
gvg8q4kM0muAuWCq+zDTVyN/8jPisHJ+GY84MBZOceZkw35S0TM4Y9A3FsCzrGId
7vS0jpqhtRcW0q/XKYbjgRUU3xudK3KJoc/fUnGWAr+PGFI1WwzNzcCGLFdl0j4x
caLvXhZW5dG6PmAwPErtqlwphrSVJ/15SZyjbyuZZe9GG992YaI6ujmuR92T6sll
V4YfhCx4IibUz0DqDQ1tIuuZSvct9PKl0CdzWe3YnrJv4WnMu6v9xm860t/JSluK
ohcGKhwy2bk9lPEqjmVkRilTUh+Fr7Ppe2l7zJxcApOkGWha2mms7y4GsgcrYGhx
7DIP61H/Hr0TRMCsDVpsIz15fmbgQtm5Syr6MZ99Mm1nkoEf5E94bgqZMfxTww7A
Cvd6d0wR7TzquDoEzEqhDe8whSqCqY+eFFoJYkgXmBteS7epSbVkUG57xO/hO2s1
SasbZLC1NaPrgm57+PgDSIAu7rDhYulvt7TrAAy6M7iaWs0Krhmuwn4uoUrJ/J6K
oy17l8yqV7UtVBvgjLZJ/cSd/NcMNyitYZX3xnw6vxCJ3zgjHP1jBlPQgl+rbOCf
mNW4bSoigj+FB4G9LE0mZwIioLN82WFfTk0H6BAQcYxT4usQyqS8YTXizv/lLuZ9
xigyT9QKLtDxDgtwYdSR5imnzD3IBIrAFPaqO4z6a9+ppNQfgQrva9ct0qufJX3l
UlYsLoCOvPalm+Q5swoua690qQ/mSzOCYkubX7ifDRvgX5LdGa/oi4nEyD7+JNFB
xdp9l6xZafkHqDVfHFGKc3XKy0EtYdhZ64W2GIro4wxMxzGNBVzYbN/h3uAjczrR
J7l6Y51ARNFosprwwSmDMaI+tzugjZV+kx/PlZrDTNUF/URTTtSwTbVFrucDSomh
efHhc5UWXMryeO3WIYE8ZWNpJbu5ueU0I0FWPdpLuvRQyyB94ESlnFrwwR45X0WE
Fc6gy2JSgsIs0jOOafKyt/Lj3CvVFl0Sz0vYTVVd+gnaQ5rQjSWXBT+byNAXDP3e
JdULDvi2xuBXHyRJCsYBomSstaz4D+1CcyE6tK8UMV/WRSAH7DDVOZrsHETdSjtq
MIKCX/LESfhqUMgwaKPNKwd3myycSMYpezDygniE0A5Xb223gdaHx3wC9OHNNq8m
oSSg1twzTrbT3iciAMLEnNmJnGNOohJFrnGpI0XNC4a1slFDyrxrHFIhF1QlUhFm
4oqDSjydNLgoeakv8Elr1huV6CgPgKtRWE1wNPZ6wmqq+nwXl7g7vVGhiclZFLIN
UTXuqqjAQl5OOFrpYnBPEYs9pg2/PCeBjbKv+mjiIF2Usi08SA45e1bLIKb42zlP
aRgKn+Mjeh4P8xV/6NeEXbzgjQmnEeveJQfLoC8xGA7YaT9HsnnPL7AQSRKHI6P6
QWaO0MnvFY/b8/hsTKtJEjGkjIZSlb6mTs+7ObAYi8ViDO8OjwManac/523eSEYz
0+gt03aDbI8+uyxSdG8/YCB+EynrAnTOQekrupacyE89wPBxa2Vg0PWdYKMO7VRZ
AO8A6l8nGxmBNoYdUhjnC+OMcCastjruy/UAS1xzM/mUYiWR5z3QzXJiWG4nhv3L
3wODG976TCdSSEp7Gj8yScCXa1417AKTy2V9xxLzjalVRPoZcsiNuPN0WBGG0aKB
EX+hqqMLbase/GzJINYJt1xGG6E6xF1LNsQEyuFzJyhf1XFFIgOO94viMGrK/61U
NTB6mNLivn9NMXb2dm6GhEgSYfLzCTIRRGiXgR/TTWF/AVMII6zMHEM29TYnNMGq
Qzbsa/c/CH3g3FSP+VLDjdNHlJsbO5+smvQZo5QkRkcNI37j1Gg02U06rfyrG6An
xsb5imRfq1Ns0Rvkv2w9tJzJyxGOU3G1qaoTPjhk2P0dQI077gSnNAFQpe2fGV9O
/HoDga3H4UXyRWYn6gDeEgmWdHcLc1kdi9NrkwwbMDYk/7vAH1cZ29lyn7GKIYP0
2V186KsEFyDxopi61qugkHEZQQfFquT9pG09EU/HwQmf8AWOFzDN6oYvZyE8FxKd
cICvaNxyeuej/H20t4J+zqaqAu/zBxGY5BgpUgPZ0/VYANm5Wduh4ixclHF5XNH2
eOVECPN4sCi0BKew2aCd2LlnpMjLTQhbisxaYO4jC4LFZY/CmywyzZkViS8QcIg3
yxTovZxApYdTVOvXr3dTg3bOkkUpyDFbYnGmv73/uW1fk5U7vMUgv6UkaebvxEGI
YBhZW6uQ5/Mz/K7mKJntkNgIdKFEV1IDKBmQ+9TOzPE9xK1Yoi84j4xTD+NSkoOz
za9YaXkzgssvPWN7E3KsF7O+PPSqQJrXGiXZsEdH4FvFPANa8QABmDCt7+C7fX8e
/YXuu5unqtZfwgAIQIXm9jWcVDyZyfzRo2F81SE+3NdY/DHxzcIikDk0jQyBZp2g
lC7yHsvxfb33m6fM5OKFbmR4iEsmmSFs6PljUFXBw8sST/cG0CHJl0TQomPx4Qr1
KBDMR//Eb+xEBWt0zrufWAh1bUKoUSs+oJ9XXDSAXYCKCDfl0rL45IZZn4ztowdL
7ppp8uZ1eeXqQ2fzyTQuSl6cV84ouj2h7/NKBJalNQGPBK12CxUXSMOwOk/lznzd
fF9OaQOaYpBkhJ7UGEyqDspS1gri2Wn6xoRswmSsoDk0YHQv9S1zpy4mpR4BBE1a
ffH3ypGrZcmJLiSjJ2+0glFA/Ytl82YRaMQCsxuZ8SNs1HAgntasgYCvvXp3lArI
9KN9wfpYHFaUYl+Xd27Zsk1Fk6NjrZsaZNc5kK2m/IGVIzO1Vc9VhZMhTOK8o+ea
z/U6FDJxhPo+sqtKbzWCficA3CvI4DNOgnhEmBhuEt7iYWjbH91vnk4j6njpCe0X
JoRIDhyXMx4zKlLTZF7pCn+ayl4ccU/C2ivwlWoaR0cqTToeNvkqGCYAiaELqMsS
xh/FCjtWYkyNEVHN01t4Db3jQJZ6102iN3EvmNmfIVUdC2wFyTxD6nHcc7d9mNLO
88jiOfgxL1t7M7Om2mh/GbWa9lq+Rw4zy61FbWb+j0GyHGTH6MpsX24wJ2RlBbEJ
+EG/VhUyqvl97sJyIkDBZj/f3rkaLCFdQ8hHeHq974WYHPfiTFPsfUCELp/iGBof
1FRFesN8LsUtI9KeMH3BCPaF6rqN17N/oRrhD3OkNsyibcNm0RdzBi7NtbCMZPpN
+2QUP/tuLATcCL1afUngEggtiyTv0EyaV7g67OBezvOYLA+ayG/IG+cRI4wFNvPV
3k/I+LkMLH7iJ3aXP4mGE0nw4cKlilF1plHhYyzxpe9bC8gfvA+q1kT9ec1zQ5Pe
9AvVRWpKPdQUrEA0PFuJKHny9Sniqbg0A6U+11qgKDdsOQJfOskWcZkEnSfPNLlK
tsUYHCwM8Mjj7o2fo7+JLW2kSp8HKm7h/wAiA5HZkxza2xvw8jNzhdNZ4sGLE6Q9
PWBrRWwlCQhuOzZ888NrseIf5dDQgd/NpjqNk/Fqnu0L8YPT2rtYVS7YwZVXKybo
aHpAjnDJuYorXpsb6/A86nzBI173Wd2M1KmVKSNAZDlWw6XVU6mHDoo/ni20vZp9
lpWDrOBr9T8vQc9T4HvQvJxbPJjk8k3eeZQMANaizmS6Uxn7ELmOEUO88SR4tulp
0DmKAnR6REsmT8HcusSBjW+Ey6iTcJQggzF5KatFZP6km1uygBY76UWScYpP7ls1
4zJszuJtaUfr/anWnC2oftEgw66AoRpKysbAwoeQZPUlVb8afKsF6RtQIWcfhS1Q
kSJnZEx6y1AtwPFs15ljmKAfqf0lkt2gZIcVqTUdj3JoO7LKgaNsn8v+ci4Qe7J9
4K1ipfTlp1mCLOHm5NPdL8Ugez4C1t8Y2/KKsO25gcfkT9aDv8gr0J6Vjx5Y4M0T
6TyTerSOrp0xhwyOYDLgDwS4DL8GaibdfmXcL5L1pNCFfiJvurTqzYeM5NDnHlzA
5JPss/t/WnfFkJN1hnsI9Z7e3BR9O8ZbtRCgGrN3MtjN3RWMmZ3LzRm82AkHZiwv
lJZE4kBdJNdUlLRfiXdjKmzMOSa20Sk7NKH3zqgUx7OadaVG3ArFH1LUKqVZKC+4
ro+3XktfnbAk1dwEr0MlYJwYo4+gsWbYInp/Z7w+C0G6/sHnbufPUZ4bF1SljdTh
hCh06DNVBEtf7Qk0BiZoXZJjIvl5pjVUZVRYZAVoFyMojvddIiU16HX2V5kLWQIN
`protect END_PROTECTED
