`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B+hP01g7WBD3Zx//wpynYpUcfod/c82bnxCSrlwwMda+KSpPmdb+7U/eA997lIrf
U+3pf3x3a9B95fHcOilXLQbhUbJH58a/4V14hyFSr86yb61ehuJhwfqb5jltlUrW
jVK3DPr540uhP63xDduA9//gQVHG6dw/vfq7ln+gBjYQSOkLf1ubj3FJ6F65gGQo
i0wIkdGNKgw1d1nYZ5Hyd+B5eM6ZPoTxxyfxeCPrilYxYNIDcq/ZUdbSjEfOuOKk
O9Ou+zM0OjZ+4MFcwk5ObjvWWktMSxCnK8Ee8lM3ZwBnIfhKtO9bfAU3OMA9Gey1
d/y7Wi+6zaCCvPDLd3J66tj9ckciurTrWK1VIrZD0ZZ2phxiEe93CogepFrqcKJ+
u9PqBsABmydu15ukNYSvG2H08vw4CJk882+mByk8tkOH8/3lX/hzqogH7lycdnz1
GWIGnlCIJkp3tRmrhfMpZHGoZuz0H6eKlLshpICM6Pqe1Rn2CCQI0+YN8szFV77y
LoNPM5REJNLwRpAqEHkiozcEO2MYPRy14Y9ua5TIM8YBoEleGxFMkxRkO/5pwSZZ
xtUovln4vhWmDjfPFj3/E4pfmZ1tzFsWx7r0g1LDSEp9RgFr+NhbSPjDH8d4Nptz
RPxK253Bh4Ej+9AW+JKIPS+cZW+4PfOBbceb9s3YvgH91q+X47YEFXIvTFTzC+vV
diWkvhCNQlZOAJYkP8OfvJoXyLtsw4yBJcUGCPBaT0c=
`protect END_PROTECTED
