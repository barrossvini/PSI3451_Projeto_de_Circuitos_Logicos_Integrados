`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NCwDiVtZpHA/i9R6jHTRSjTdnReAI4yC8zLdo0LJH0gcEHhzUVM6jMpLadDN/1Ar
EIkKbL/6KWGM3yUyCK+1UxC5E7iBeEivREWEwJCbempmy1gHKrWFI3llS/A0xK74
ZHyxT8Lsp3RLY+LeNVphsfUkoPZ59IhgWmvgt2Lg4ccbGTGXdbMnWC6hRCqmIJum
1MtvHltEuAag4vDjXPEq2e5mhfvCyKcnGwTVGyEAa8mJZ9Zow7l8TaJlLiLRFTEw
QWIk06HN7jGVhWoupA1c7UtZA0EmW5erBbuSq8nu3SybRKBAtPJXC/BioMSusjsF
ouORqzm+VoxnxKSUSsUe0T79i/DIg5YHwSBvQOFrHHlpgQpnfQX3s0fK2f6sScR4
4Lk7iBdKHbMN3iZUeVnseUUJG/GWZ8cwBeUw1Eb4hbWP3+37YtlMVNdM+mvRwl2f
sxGYWBqVknzRiJuu3g/EE0E9UZBHK6EKW8M1JE22Yorn38pZ3/rgZa/2DH+6M09I
vsm06iqI8uD4qWMJnwRmcQ29Zzdfqze7z4BBbmiZou5uVVbaJRD12Cqe1r1nhd8o
6q3AoRJtkkoLGKQZFOeT1h8s9f1bWcZcI4T9PqHTNgwC3aNTHiQE153Egg7/zp9L
DTj60PtObCQsGynPQwab8jzf5fO1ImqMVKeMufpVfzp0iqSteKrVnLPOEDJbzBza
vrqWhikMqHtXZGroAmyMR7LPVd1ydWUggCmTZOD1Pk/X0f3hZqH50AVfILtgCh6d
HZ5LvBSGUTc28gVlEoAzqvruSb2O1DTvQQpV/ZziSTG4UAw1OJomZbfDGCMf8Pp8
79LW9d8ppE38ASaXVn6yFs4pg5XpaeXRD4hVg5oarUw52Jz/dkhOvyDsuYWJk8kv
RYI+ROA0Ux/+OpSa4fXr9Amujcfsk0qlilgHS4B//7tV50pbYHKXh5wi6tYIdwHu
3GKtih1PVtIOrxJWD96hVIc6YgWJ2k1F4hX4u7zYExZs7h9an1gHYFcwWBzuwsVP
f9jpcEAGVUzJyv+WGM0V1pAEp5qA2E2gI8t9pe62az06jI0NcW3NIFpPUZOyKJlg
QIvWJltkB+d1DM42PzNdxTn+wrukfVC8msz4yQIu5UJUP66Y8vt7JzY5m9bD8cSC
bLaYDEMdBTBiUv43mtA90Tjc1xoO9sBdrl+xdQk1biuZZcGv8f+HgVpI7DUZBU/S
nPT81wnGmf5MY/flPDW53RMow3KMUWiSfT5Vjx3bt08UiOLxpFZElNSW2EhxJvHx
Kc76GE6lbxrm6DEDKrGNZqqu7lRpAOejRBO/BPo8JytOwa8J4GeT1fvPwUQ4guxm
w2GGcZi8Z9SalVcB4JFcZkVFho7+4+mL/Q/kbpmv0odWKF8PZpPivYgDLVcvtX/z
mGGhNnwX8sTCbDyQqnAmcav/A5iKRQA/5ewN/7L+XOJKLvj0Yec/LmS1w6b1GnVd
pkSQ4YKFZD0g5YbsVb8UX5/3ZBh6tlKQ15Fgo5+spxFduKIomZMQjzitATBO8aeE
a9w4l+C7VuQFpcdFtDl0BdYhBratpUELyrNPwuQrf4uwJQ+VLVahq/cnrruefSFR
aErYOF5lHFd/v/e82IERuND7pS5cwpWAFjaQfsf575Oyi/1nA+ekTETOqA6F1rAC
w3czaclmYVQFRohpmo3Si53Y59OvhSGchx1CDi+Kbn71SG9Gu/KaYiRvtq1Br3g6
vlvLmIE95pvY+X+a3hNhTijoO6MSDkHiu3bsMnBgdftDC+q0w0hhEK7TUz/9WHbA
Q4beOvaGpH9B3Js0B2oMJpaUuq1Pt5biGRDOz+UECv5o0zueorD+3TNzy+Wa2JQ2
RGOwVVbYWNHldVxGneDGVA/al4yqBD+B+VYr/eyfj8JU731b0PnHtCGvGuoAQs2X
+qgzWdl8xAdX6MN+i1OB41lc8e3CseM0ozO7T5GWkckBFqG/2PAgvBI4kyoh/BWa
euiLrCmbtFPE0G7X4AQM1rvTePTz2fRbRv8tN54+Elj84K8/0IEDkmXVuK4fpHd3
p4pIHWzE8oRw0EvhlHHVgyBxIMPxN3Kgjz9IByd/sEJqyXxszCxQIyX57tkm9YqZ
dj2TyuVBd50vJ7lGPtMeHGCEE364APTDRk6Di4MswWk1FNTylTgFFRYBKdx7onef
BR0oTvNFAJ8TtqhP93xoaHHhO24rIxQc0g1YvSoxbi8VlLMV/9GvOhpMmdg3KXAV
WIC+YJT6vq98PzvMwTuaCDh4+RxUwOe5MxUvuptxMFT0Y0mzr07+yk4b7/2M7B2F
yZvdpW8ax7nFSq6bN2IfSfQCEVpNZDBMoYfgf1B7NLkbRiGeM+MGOwYM6eUfBvew
KKRgqn8rWZVHxFgqeHgjwRbQoJD0KBfpEFU6hzx8yZiUnA9EjWzFbBCJ4gAgX9uF
7wqgukMOz65sddrUU0AMyXjg6JMsT7bv2tFINIoNmC4oNd9itthFYYj47Z+VroUc
VvNAVr3zL8y72AffVlOLQR9RZt6356zzxi6paf6DH5VeEWJF/B0LUBNh2tcsTpgo
o1PRzBtP2bTStZM6+/jBX1MdXTJqSAqHn1WgNz6bZqCx3nIlvw8NKhd2N6FME0+N
nrMufThJFX5rYre5VrinpoLTCc1TWDI1o36bewoMBQsJ226GWsgKfNJ3X6oct0Ql
ZKWUk0yZ410+PzCW9lZHGL3ts451Cd+H75XwisDQD3J9u7V+k0QuOzk3zhY6FBbx
LLp85dl1CIdxoQxVFMweHzkHncRFVlcUoxO3nDUlHoIHPTxh1hhxvUzX81EOoIQq
n6cgI8hnADHk2CznPM/x7f5VQqkQfCPi3kQXpX5K3VilqUuVFDeKqGqwXt8OocAm
VzqKSbeLjcQlA+64vW0shvJyzFok0iCJcN3f6xwSO1dkClnvJA5/H2kmOwMMpw7H
F7tg680Nc+JA7dG3aUVdZzSUGOq4OTxC3LJHb22/JjOZEUpbmXuMsLfATHZSJFsI
gtzTvGHZjt/hwu3gHelxRGvc+f+4wN2yzqb/op5Ggvo6XPWGyDJEUBvMDQJUmObu
m+gRTSlq08n0vzyV0fDs55nQE6SbHgVEL0zhbIAicc4s79aWJf67v7g1NNa/hrcI
S+tfgcbntjyTMLYp4HW/ZmFi5O41A9e3bags3BjPj+kEt0mvIJfF1JXIk6apUUZB
NLkWbxPwqyoMFmnlXsMH5JWnb1DK4JPOkDcS7OO1C2u1Jv6iOkJnm9ShZB/m/bD+
3XUVM9RWymK1OX3zC223u670ngbuV++q53FvL4svtFM/SlTzWJ1ZJ9uU7cmG4J4K
6yddEDi7W0NrbIWXufLAL2gqPA1sZLPeYcXGe4L/fR82/Z2LOnqTTr2y2cL0/3nd
iNskXZVJMylchs6ZNUKbzNQPM0LfM+gd3Fhm4m1PARJFfx85iImwH0yKrLBw8ufU
3jLqYMIdJCUPpi6kw2iVD41AWK7aEOBK/3HINmo9i8kUkDeu9XpxpRJspnvOJDnS
eMM8zjqBuk2HnSA0SWiJDru4zrdkromktUklYy91Fg6Ewzmuof+scgrn3dqLfSdF
DogZXx021U0BXcPCKwamWA90zQOzX525BIgDoLBfze+KLKA9Q+YqWVb1VKN16HgU
uKTN3OrfGtv4Q9dq2kaaJPP/fK2P+MfZmHaRelehAWa+fQvdq3CL6JOQJAvC1a7l
9oYrWG689yDabtz0WxUptQloNISWZIeuseIcC5JKVwie0dQAWhrcuCSdrsipbbtc
QdDotFFPeykI4sb3CE2gfG0q2paiG2e7YqgYkgPvCWAnkvasb21EHV1IvIUIjUtn
ODeeD+LiYElHpBjASCzCmOhh434EbVlcT7iYoIePUvkNcVyWSwI76mwrzPNaZmCt
TtaxDBDUZviqONvahAdLhR46b5DHIvcpJLsYZBQk+Je5agd9v+xU+oyx5s9ycWc7
udzl/K2rto0VIKa1KHvYGJFSRvTeZisR47k8EJMQ4zTjrCmSk42Nc3zLtvIyDcod
LqWB3omjpbbQK2o391zXPDZFFY3BFJXH/thN0Ur94XJsjhK4A1BiDgfKqJsiE2iE
sNDhd8W1MN9t6G7VUj3PTJUEc1e1Vb7iMJwoIbF3B4MLgJVvnUB5f9skwDwtbW21
3NiUkiVZH/v2nUugFvv5FdNN3mE4eVmtnfWVJjs/vrEiE6RybE0zygrLZxnTv/vZ
weFKO2jdcYUYdCZq9dV3PRMITkF/NNpRymQvd4vOkCH3GW8nX/aaBqEn0bxOfq12
pMqtsq6xHULR2Pb4zB5IxGCQKngfPsriLiXQrgIuyLRKT41t4PFvWC8O7HdAkVMV
MC/eXXHjmvOp3tniFsizseXCoXtP9zCWGMIVe7UV0apiV3zA5YhWXbkXRHhQvG1J
yS1K4LrK4ZmnFc2u6lSPHuXRpXnQronIlNsnskGUiYdoTjWjrO0QjNrx9GvyJez/
IIbaYHxP5pCnAdPTEKvN2aH2hKmblrg4dS3WgbDPj8njO22gWMD8cZMLofrMDqAs
JC6hQ4j2d62CbwvChGfekon7uvKb0jPASVSWfUnEsFb/gMb/PRFsztbSh59GSAPv
wgSBjY9bnaC57zqDD2CMeY0otTH9C18ePBf2kx6bOXN73xW1HF0EK9JaMZ6i5/p2
kuldvn/35d1kvf2J9qOPaZ6oWimPLFFkPToL2n8sAWc82XXzmHOiDWp6BArU/rou
UiGrTU9nIUNXlTAv7VORA0fS4lFYNDX996tl54k7j8jNT0NEsbDU9InFNhQlf195
YbJZ6ef/wNDQ4dfpD1W0+Z4q9/m2WDrvlO/tKS3fofBnd2KTnPIKZbFm9Za1jSCT
gYNJ2CYHdDEXMyd2sJAMUzgKdp1sHhJ/l0bFDhNS7qGT8ymQvoenXdx6bfqCwEhv
XYtqwY38TghlJG3ESeYBSfzbX7m+l6DdaxaMOTrdG2A89Z3pgTO3D0bNJLSPdNrS
nDhFFngN6HxfOQcHAG8XXHKAHZMJrgpAgymaKAp+rKdRACfUWZKndtnufh1LBnbf
FVO4VVxa3TDCEsbp/cNUx1o9HZQhJ4Wd/7xgU0v8HaSofwQHtNdciVepyKq3Ai7d
wZwVJm1DS0vEmCNWKf1nQRMoLSVWU+pnQeJmQglOnRXhHGFKsq3D8Fk2F0CXnJPS
s7S0mfYHD7ccDMOipk2ow5WXU+WWvW3CL4wjjs3i8SfGvj6cZu5Ax6l5KgK7j7Up
3vp3mNJmlrymqqZf/2UsJCJRxn6Ul/FAiA8PgkDtnSJpi4OiKeVEyFWjgvSE69lW
s0jezD3nIDJQwBHauuPLjbQn5ovZGcBuF9GG+LGJj/58aXDjMYmU0d/OzHW1/47T
Q/NfkbfMd3pXJgwR597U/+1AMe9IUshslGDgvBXQ8OfbI/8XtgT5x62+9CT6gqT5
Vmgeq/8nWZjXZvVFXcPGytm8bXV0Qsr2xtGOb9CwDqQYHVFq4rl+Ld3U6GnzJfzf
X2grgQ3UhBEbbFFMB57j578zFOBxkgZxTdQ76n14RYDukj27oJ0ZNYHjpQaJOJb1
CHKw4adKAsCR7gTpF5mBC+En8YZKF6igu8yZflXeUpJPCRNgIw+z6Lpq7dNAQNBG
iH5nB7KzMtvnzD8jTvcJb/TVlio1T/QcD02uW+e45nyBNQSjKseb3JcnzPApIpDW
0OE+6nOfkBcAxJLl0evjRfum8NORVolcle/8QHjAJLEpzClZlgSrQhBsGHSrmMoA
VpWdPPzSdHDzY/F2GJqNVP/JNJ5zdPwQ5BXjOvg+cCAgjytSse+AlL1MGfVowOKO
ah5uB7M4H+Ca1dbKJbmkajdSP6wKaH84ExdFUmX7yrRc2jSopeJSeG1SsJBi+Kej
qJWfxZsSxX3TORLfcNjYO+0jthCs/JZz4BvtM0K1e/d7umNcr7ohjufTnJvyQfJu
sN2J2REEhuJ6qAAoTKlu+wzZpu2XA97by4olYqOBpbBwVSYghI3RqgwjRhbU3yLW
rQApLnnXKwMNmF/WFPlwJvAGaxjh3LZTJkBPM1rPhfclLzbxP88Qa7H5dac5cya3
G38Pw64f8rCdPtiJt4ZI5itPAQeI9lfPyoeObwOr/voyFd0WqbmPQUOWKwdV9rG7
bLniYmP3OvslmySRBOgjPNpeKgAyzkQJuADLS62tHZ6pzCiEZAznGiXKLX+DzK5G
ueih+USkM1ux4ScOpAHpI6snIUzxVApdwAzHPpqroN2JfTrEql56sfNKDuUo8jSz
vYPY7IdD1IyslHUYwt1cWBxnRy2S5woA3v/GGP7CUBz+TTZagD/xeKnB0OOCpjlR
8tZDC0zPZxydXcPMHacScEuCU5YfcXhOD9ISXlym8PZ5YM0hxPz80hTPdwvw4exm
4pH26y5xFJgs8Acm+ioBl5JVMEpO8mxXWiMh62F2sEUaGKmN+OiO54e99OpKdIyh
Ig7oEZY5phemImunD/Y6IAo+QdcECQhh2UNwX0DPn97zJDeGhH/0Oxm7z6xbflwg
yPs/fJ2jV0nsis9aHRo4YhFfuyJyOI8kdnTSGjZkWEU6I9U8Fn6dmSE/BMsB8N6X
4tqKBMOTfsGgIjIpTJ/5jXKfU/cycM0IyVVDetklyBC3NiKsvNqNa3Q+pL2jeweE
cKGJo2JENPxZYCzejR2kSBwlDv8aOtv3srdkY5hkXqOUVu/PSe/CwYkebpoJTlhs
fbVg44BN86YMyeT/JSoAcjid/CO9diDXK5QsYBn750jV/PMl9i8lhaKvAQRNHQpV
OBJz39V7pCJeUm1J48kPpM/oo5n11pqIDbrZvTpd64e0gONH3p0YisIntDRPBrOh
7P9/YWdn4SMZnkuSXXQAFHIfqb9nainMOlwnRNg2feAdXvgXcws5jbhcqAbZsRSR
/8ZTJkwYNdRZ5FSCJ6KYHzvM8K5SET98uL0fYiiC9uNxZNd2yE/nsNgBgpSjpO1p
1EagFgt30xUOKIfgpKyBpCRH4N30EBLbaC03iQ+eyRkRjf7LF4vDGhm3SDo4z6df
NEgZbyadUw/0vJCQ1Pi79CNyxxZbdi8aNf5K0fhifvvA9z8s7B4oBVGmonU70qM+
pP+oxR7vI93Cf5cvQ9YY+P8TsnfROP8g2HM0Cwk2L5Dan3YQrLRro6YvflrGD5KF
BUH8DjCQ133OXDqT0pOzxLdYiAVKg0xrzdh1ld4s3/MASzLHbLLXOPtnYNT0+JZb
rNbeI42071BCx1+4xIJV8Sw5MKFQo/UyoCD6XAlECW44KvRreRU0dGRNY2o8ur4l
AW8ugNvRpquTG97rZY0mpQ==
`protect END_PROTECTED
