`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NxpBlPv7kklTG6Rq5PLnASutqD203VO46Fl0sg5ukqp0cvpAmU0AfrY+97xqdsq0
4ZCEBsogNEGxisVPFgMlCvST/jRSHk4FJ+tS8fUkWXUEJdsiHpfIXeUtv9/yF2kw
55FAj8/UbX6Pmq7y/NDZoMYuegot3fxAzl4lXS5SZ+7y1FHqmztc+gW93V+/7Cay
o9c9dova4GuqO9acyafbuWKunTysH8xNZLy+MimAyyxUZL0swfrnQwA2SkjRLg8+
IltLeY26RfpzJz5Y3FHBfOkFFsZ9aUAaI/pAYSmSx+Ea+QVZyYPgLwhOtN/VboSF
U6WbFUK2y51J3EpvNqFXpDpFvLpL1b3t/jJ0uIgvg8s8mFlw8VGrPPj/BsiQyxEZ
MH96/0V75SHm3B8R3c9TA0gDznqRFlBQEebK+UC5TPuQ2WB0j65AYqeLA2TrhnIp
5VVna6fTNPHJjOYxQq/ixC3PwbWF1Qj6M7cZoUchETklUag5DeJPaIuYtqKRk4Fn
MDDnZQwUUrcPU8f8n0PJ/F/JK5ROo+8oWzrV87jwgjkZKMg8Ud5KXV1kE0ryr+O1
Ingz1ds5RjxM3qEhDs6U4Kcsyy1KOTjs0kNCjfOaJlmc2DeXIEJtV/K9/26s4lyd
T5U9wictLfbw/BCPmTV6iwJu2maU5Go4tGxJ6VdCKlWIELaGYPuKNAlK670jBPv3
oMdKDqfeSHxsGRP0YVuse/oZYBXqLixR1JiqcePbXh6CX4Hsz3mgwrxBQxXNCg5n
s4/H4eb2Q+8qAKlKL7QbUujAVsxWPkKEPsvFoF1/ZNxqbVW5v+oP4ZPM6S+KyZQI
XFgM9NDLU2Qe6XvGheTS2IHHmu1H2FWQlfoV8FF2df46iMRQItdLMeZ05kne6pLY
fjJJZgsj9nA/Yd1O7i+rtu2tBmgwbto9yqbX3RSr4aWJCb7SRnlZk7y/fJeOGM5f
QsAfPm7gsdqTrhikFnlbJ5PZCbTfNkWhGu9Li50KD1y+gcY3sDbdCOJdP5yIkpMP
9aiSZI+e6drMeKp2fzYllcAN/QpUAVVkuT66bjEzmBxMUc6qtf4mPz3ClgJqisN2
S3zJcSL/pt8wi6iGi3zGhv7LUhI+CNGl4IQXtuw/BXaGHnoBT9y9x7Stzy3N3nOq
w5JMOJBBSFSAs4Oyww8PNZZC8PYTpE5qKW70jA7BEvCulK72AIWLvvogwU1TK+gT
P4pI/Az4J+eaVjd18HJRnauf8T8Ry9vM/tHj6noAkpecwpC1xrCePajOoLe7p8kW
mLXP4fBpH9ClISxH/xR2U48IZdzf07YijH5j3M3+kjstDp+MypVNJcOdG9Do2IAB
fOGxbVvVRqyt3Zx1+LD9zqTcsrFHug87b22kPpZBwTUfC6C/huxfjPI8Ucic/p6Z
MW57NRHLGpllx0qF7NnZjVVvWFjR3apa8gpyLZQs0fBwe+AIeK6z5oG9u6Gxh5fc
lwsPH+P1xnOyy6bf35eEZnoDqkTVCYWL6uToxhEyxrKgL4AtGZa/QipEdpmqj3gj
EoVjnPfTPXKuiJ88RJZdeNeieY/5XyVmztRH7TUxUngHBLzOAT97gSbd5NlCFvhO
emfjCORkwFtoAVpZtjuVyYDKLugIMcu1TIEifc98anqT15O+Ain1o7jbTYdv4T5n
Ac0Jrq+Yy5zKquiwTfZzVKYpQSHTkvAV6P/7FzS4US5ar+NKHqwUF/Fi4GjNcO8+
mjmKqHO82UOytWCCwFJ6tSSN9/hXeBQ9AVaAb03w0Iqbr7NeTTvmteCdvQA2od+q
9nSYaGdTf02LdY+qgwbeNXujXxhNATXTYGIFaxDjAoHUHxZlAXVXhZcEe/oaio+2
KmDmEEVzb4yn0824t5k8gzB4MNWXc9G8rN2TLX9xYV2fpMhtrtMx9gYLmy7qz80j
mxH+RZVun3Z6C5ZUegd7SHSwS6jFHXb9Lt7DxXHdA0vVRNhtBUUdFXK1LyPKZQli
AUM6cB+Vxa1OJWZ/er8qPLuenpNVW0ZmPYT/2wqg0glF85p1tcYqw+QuQ4ckGRX7
0ccadYruP+oenZcbVJUP0H2Bfir73jiLBotVZ/eyS5DplU1MjhIKXJGmcFiF7RnZ
jcWDunS6b91XZZPEOgDfZ6Yyikf3U5ve8hHy5O/fc0MULRFMRSvkr29rZp9aCanu
JtxOkegh7I2IXeGZ/f03S2sp1KfgGSBwhkwt30i5iuJSEKzUGDsacjDLV8gJsa5X
3uXLqgmCOHTAxfkN3dhohgXde9Es0I2I+Oo7tvNg2vkgGH5lCrRLRhzG/MHuDSRz
9BIhXKSNhRpu2lESxG/jYEfh3ATCoKbNk4GVeNnVDaLizeCp4i+NNUJBk0lFKOlj
ZFYtaBQFXLDeKjX7w28Ino/OL5ePHJSqsORT88LJOPaT92KvwJEOeWlaVjWRfLHi
rcIdcBCzZ1L/tsCEvfiRm+7wRjix5k5qZJM9VSfn7t9LbnUEAd9AcWVlToLsZBdZ
nuuPhT0I9+UQN1x9m44f7zCYzFCYICyH/JlQmXlYE1nI+qxuy4cfkfgDxC/PgPfK
VPWOTvBIFT7X3oxUS+OrtESP4lKAm0ldOGfpG/adsmZM3GpvViRg4cD5UV6SpIG8
NcAveWLG4hLkG8iv2jUK1tBZQkx9R12QMh87Rpyd4wqU/cSo1qKwrxpw8SwgkF1X
b2upRzNVv/QzGW2tzvrtSS8XmgnaN7pIezEPFgg5Tx9l+qm0w9eLUIRcuN86ccib
PSzJgjtlYWluFYrpLLb+VSfk73BXY7vq6pAGwQaDNu7Fg5b2v71vZF56uPnfRjJQ
JA7lHzU8djuz//iarD0DW8CZ6te0+uv+i3I2mfKWnKVErE7tgk8ulWWEmOs9VdGI
I0VHon5iEXyfChmgIgzQqArjmp75eF2FP4fU18EzDlV950CmRTgp/SPECs2UheG4
7oZh3I7m4lF0N5dLJGnHXPxn9GaZaRGlzKl3+TGrY1zdncC5349UAIvgaIelB4as
w9wmRyFS3ZYUU26J64sewni7UAVM5ZvOUwpoUnpCeVnGxxEGPzsKgiYXM0TWjTBx
m9FlS0KGhVeCsAWFNwpm+q95U75YOVJlqcopymCALqB7/RgPohlQ5d1mYrtyHsSF
JmQa70WbcQ4+lbcbLaDDUTBXDKyzdwmmjDMdixBXof+Hs2TXoiHYWjTMCciVpp0p
Vfp+Z4pgg4ppJdCGkc147V+BdqR+8ibi0CXZ7Pmy9/F1ODk/sJUrhrQXSGF2YQIS
XNdFGoP/SgrEKm0X8qvwR3rHxOeJ2+Oac9+KFca4rpNI5pyvCAxurSwDK9I8OUyy
54k3orig6xQD0UCI+ReJu9FGF6yeCOKHvXd0Xcs4lQDWn1xTBv9Ziei2VcqSmjGx
8fNcD9xXv8fDx6fxMudWmg//PqtayjLWgpatNT4STGrO0GBnpYFJeRKpz9icd7Yq
6NiTj/IxwlI7D2zlbeSlYm935K7gbK2xohfWGsjjNpUs6iLrbDLqO3Jch1jLvtzg
Za9DeVjiAnwABtS3jAVBK31Rsw6LHHqnsH5kQMIiiNSEXTBiaQ+GvHY8TF/kXXse
vf7JwLMmFjP6eVmkJ34WLswuI1+WLFYEDmCXhTR8eMdQS47SeOVVQgUi5wBPTRJH
cF/yIawg/QxRZnj+yR3SnpKktN+76iNz22EfroSF33Jrx6Yxf6L2saEsLvyrIAEB
Ae2Ku5VQI9IDigQYYoDMdJTyAV0vmzHb8fj8oFBc4WuXQNgu4seOZJ+9j4dPJd/a
BuDvf18lIQcDpBe3eZy4Ny+3OGsPDWJ3ShAb61d068A6zDvw1lwzAFIIQkqrWmO1
imgXeZoD7d197F1TaDT2wJwdLXdCCriRBklfrnyVE9sffV2fgd7vtB/oaMFZZVbB
DRPMHZXNeNAMxdTd+1aSZqM/qKDd2K9i1096bKXQxYYRlGAInBYrjRc6rL6Bsrwn
39AFyShyt1bsQugADmFdW56w16jrWMwpbKiSbrgaywXgEtabBsVQLuS4M24NlEUN
qVD51kPgUQdFAesJVNTqBKeR5k8/JQmqM3YE5U0NLbUZbCRTvU2ROYI5VU2DP5IE
O6TGWJya9b607A0L0aS73d3oS8fsr26e+hENUFC10fPHJrofaS8ZUDJ6/XSb3z8M
TsW9c/LR5RJjepN/bbOODr4T1SWjd8xEsqgzSKFaxr9gMCHQn/dtO1gKBRtsK/vV
qQKHzpCfDCWHgw5dS48oaogcmVS89hWsUPMTuBZVmPQLCRHvFJzELfi6yKpfoD2O
X2Y3AUPjuJDHNbq5SOlPq8xXhxvjNpfDLB3v3ZGlZq+fmdjT7JnqsMybMQNaOKKu
0tuabH5utPWGeNtK42mRgZQVoFkCoT3ofPcpKDGqPl6iPrTUNqyUIBDJRYx/HK8g
H7rGI4eLFQNo7A8SteRru3Z6cjl7Xxjhvp/dmdBkZ6eqMpp566a4GQuQnVMbV5Gk
I87kj3z4QKr2OoKNFI1nDl/bzC6JUe5tz4+1Mr+E3/NbACSJAKlL/lgSB3nAIBMa
YTJR/S80A1lDQa7i1TYjHLpr0STlDRYuRBiDmMuAtNtxlFnZwIolTEvz6cWXAR6w
x9HpW/Nif+SxXxCuR+jmXVrjxNMiq6GL6GlMPy+gDfx211Z2aGYDmqCBRUvNt6F0
jWKhFRhbQwFmhOSzhnIkY7Q6QRAz36lj5WPnuYUZQA+qC8De5e1KuC/KUnRYM3mD
/k+nJjdTdi/Maz/htgCEOANYYQCSREBQCAu4YDdI2bR8gJLDwtNNZYW5tCpdCvxG
jiA2EMkA3JO1J394dgbTGvHKbr8Dh3FZOmYgwr2diHx9T6MbMFWyeIsroXEGTWou
1D44pMu71ETdGuiAmDm564hGg1XrBD4I/rqYFKykMY3rX6Lw8/jSNisg20bRQABo
h2K1+QTk+58hUGysl0Pjn+9QOAsyiYE1EkmsWy+b8wAU0UjcGFFGxLqM0X4/Agcd
MWdgkQTllnSdNy9kVGFiz3Uxja26mZt8n3On53TJT6LP8r7+32CaIykzregQXlrR
TBOxm4p4VazRFDEtslVhBV4jW5k3f9nXhARubQ10vWrJgpIkoRruz6sE8rmdwlZZ
o2XUONdjQIr4YgxBc1PUMcPpUdzaCy6TT+o1D1Z5XqHdE805WW+71ndycA4XSoAW
YqNqpYI68huKcXOH6N75Qy1V7LHho4gmilYuRqcsVwEKm5K0L2aL8oYWPzjWGTAw
aP2M7fliF1W4ELZyUFgb78BjSf7a8RWXhd4RfM3r+DejFSgzETt/tJzACLlbnGCX
duJP277ZaO8WqkEjsUw6yX6NQYesieUmqDaF4vkQ5Dz9cJmrqf5DFekeqvzcPx/l
HMr6jDYbJnrp6O0s6mT/BS+fMVHDgaHIyhTqkozZIn13DLyxlNYcyIZ5VPaImki6
jaqj0T9qofLrnJ26BHvm/INlkFkBK5noWBzMSWcJLFZ5Jyzwmypboe7TORgcX0qc
K6ZWt8bEwPvJ+Y0Ox+MpAJNTftXjfoLolVGXo7utZa9D9dfRgFq8AJKlSy5/rIW+
eJupVUFjfY7Q+1xHGNCCB4j0dMonLPu0vEFkSUWdINPlRtIuyO4gKpyCF6N9NTRI
skTy0Z3cbJllxDftk1ol7rtPKF+oghZ17sG29ZQ2f0g6Y7BTJFX+wj/02oWeKYCA
MuuXhOjPmDjflotc5Iby7dbuM6PZZR8W1peV30PtG1cPdYXwy67/wRJcCup0o58M
pFYFSIx0E8I5aZe2Hr1dLe3mackYslxPM4j4GXPpTy20NzAX3roI0o5W2ZO4ySX2
dvanXm//YbfK47eYH7HOpQc7LoGVt6Rmm/g2EoaLbj589zG3xnTn7vs//ApivYN+
N+CSjcRBKIuNppzCCvU9zwFnR/SmqpPDccuBwehWIjYJBH3DWwmLm/it0wc+hblJ
T8ZM0BDboZLDV404yDkfsfkuSqTXLdEJMc7p8yb97p6cfnyVIUY3Vse+5xfhRgNR
dHoIzcnvHkQr/79GeATGONzqwUOTVB0xF/a7YcltbLuLjQvDpPWh9lHyBZcDreXD
hiQJIicJRhDNOo2veuQirTyHn2mICg5zXOjjV6g73NM9XgRVN3xFkE4ObYNVRMFx
0VD/wyWtgvWxZ7RLZi193y183j+MKFCuTW6UYpt2jfaLAbG95HdGoYi3q7HLR0yM
sNyj8R6SzYCXCC8gSGy4x+aIvP6rpS2ZRwrSy1bDdCtBKoWEpatOAC/VK2OD4qu9
2ZW6RnICaJIHspbtY2fkhbaHYGhidbH9g4A2/RhKXbbVN8eQqDjptOrDeKIQG4zO
/+zTur159YLry6RZRn7XOQ0f19gC/NH84ow+hqWZidEMDAbwNDSmnz1Uw5+4eEMx
8JqeWG+05aLnRqwH+xVq9uFdxgg69KCr5SdTyQevfe6cOjWGM7unwAG22w+yf8R5
Yyh44osTw7sJTZ6rpBwfLCgUCvmQpzfz8R8AeuRmdwEIaeCI1tQ213UcrYahmS2W
l3KdMnqxgpIKUMhywi5c6S8ian5Y2Sy65gELuQ2Jr8udfow98HXIW96h6x8QDWKZ
VidsnpFIKhj4goAJ+t69joUR0kcf+sgYaAy3zBQWBwxC9eyeOPpQ4M6iV8JSeUK3
fJU13sKZDimyM8d0rvgVXXeuESU4kSVXPGBYi7U5Y1EVyHyA4Jg2R7YeeqUG1ZDF
Cq/pczWGAYcvNT99wK2e7hx/cWPv4v0myWmq35pnw+9DzCNwDg+KX86Q6+jFDpn9
k7R9eMEPLqqJU65CQ3tDd6sFczlkOPEnNIUO0JcHXaSoSwhdVuzmeLszKGbHqMd5
IPdYXIBMU40V0Gm/TkF471ckV2vl748mtv6IWKcWTuJ8SJHtJXkFB2ygq16Uvhxs
t4AOfH4cICb+/eCIEzr53MZQe76YNULKsh4VINp5QY6w6Sa198C5d4L1QIsRj10b
182mBi3dR3I5RGQA8006fNvI8iFuGCY0FVJpJO8jr9nzqNy6zuw6gZttId8OtM/n
d3he4HyHH1hbsFlxgT4vMDvLkc64sxuKJjTvSn20Ur4nZSrS5pP0pG3yjTEBAZI0
a039DHmAJY6+c2TfN7dTklu1/3vuOWOPWGS6Ur5w0ZR2duppJl8CoiJLro8SPYTX
2PIlmTQA3GV3B4F5h1bJL63Ev8pGgHNocNdfCuI4A7+JaVlhJKfQzs0x7p6e7/Ey
Bykg3La3bQJga2vNweDjqQdAEkQmck+YOYWUw5keCtOrUgKxGpJ4Z3rnE3j16N3y
keD6A+SbAUxeX3IB+8nCHQ==
`protect END_PROTECTED
