`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fRsz2j6dTam4fnwd0hj+0u+9z3Kmdwz4H0z+eU1sWRihuaaMx7u1Gn6mFmm+E4nC
E6tfSgBubkGswarkq9hR1HEyEEQf6gS78TB+m67ZnH+O+YQ9EWA4DctyrwuPtBZZ
U/SD7/QOULCxgfXaTjx5ncMQjDydUTj3DKSmlAmBnIYk+kwHD/iEn4e4XBhCQ+QT
2htOF9t7DtmMH/5i8eljlreMiDXUG5trKCNCPyamK66vYe/JkAc0D0YP5qldLCkQ
++N3RgRtzw1pCf2Ocd+1GiiWiKm7BkhrtlwCBHigrsZQBBX80Q/TYRMDGOgpKohl
YtuCDUOxN6gDb45sjtGzTVrf6UWsg7LtltRDXfUhjnIStP8Q253pfeYG2R9ONMsM
L7r+FWpwph2Eypck/kD0EewK/iVcuuGSejUzy2xpBOcEGGrheSLh0AybnbjhRK9f
/hPzFH0F/W+p0gIGGyDK3PIS3l09sg0HaEVhFx7DjoxDO8z2K719YpF5eNx8DOnT
`protect END_PROTECTED
