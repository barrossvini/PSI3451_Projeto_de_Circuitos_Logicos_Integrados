`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5IRKx8bv722JsgTb+ktKMIn+d+jSWdqIbDa3Mwv/+U9dpyydvGuv/5XfydIAtRJi
8YNIxis/zzvmK+6ipwAgetUXZPwDRJG/H/5qaVpKRYBms/+mDZygAGSn1+FArvVe
7b9TnYa3ciW/pb4yNLwbgN6rM6uGRH2QQgBGCqr7a8A2YtiQS+y41UmkTjDqP0vB
hx3As8aRsPHQ9CPTcf74z+pI6ftxjC5W7l7Vz41wj1vq/Y7BLR/rsTHubFfKp4SG
W0/Y6R3De/A33DifMCLtwYY9boG9E6u045H1hQwPziUmwDZXPY3abfZ4BEB0ojYd
DmzG6ZOO3TkRBazDtI8nyAZS3nOrlOGTtxadW8E1ldxz8XjYCv02zkL2RaSUtXrI
dnGyjQhmBX8m8FZbJ+XpGqi8t/qxvZoQzZIZBTgMtgEhnCmsEiKxR1VvglaLaAJx
ZMdf1o/8IlAxS27vo5O7sRSC5Y/a66THtbotep/wqDpRkG2neKgF3zegVhKd6X8D
N0WV0cfmxftvxfkTd/u0/R+Q+YXxCG5VIuzdXYghgS93mIFd4DTLxHwEcQ8iUBom
V9dY+ztr10oTiUx4eXGr1YXsg1IuzeSsUHz64SX766fO6qIuphcIRm2ZUoaQDNSK
ftRWHhahsAv3tPdXuUqYQGbbUQYRAE6/rLTobLF+qDA=
`protect END_PROTECTED
