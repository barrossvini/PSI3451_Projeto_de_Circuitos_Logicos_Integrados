`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i45cftg2oMR0bvDW8kzhbpyJfjkSRMCfRLakqg4hznjyuYbEFe1kqXCTlenrsPq0
sZOi7FUPM1w7yWfBkvNZ8YlW99bOFBs5bjcWX9cTaeL6Gycl+lP6Vi5PmcH1lxSX
+lQKGOT8kTwLK5MxiqegPAYN+ki3c8nLJIh5i0sQWBZJe3XmyJuiGLGVf1vlHX1B
dTj4RxlAFLLVAkEFRbvNsZ7UmKenNsA6xk5oiLysaPdTjMA6jikpyzJMrjPbj9S0
hcpbyixJDY79o9vVuu++eGWDFbON5DfRRtf4RDVIymfVSGCH2lvvmdEF26XgoTUS
eTGupvcy0xO+5cwuNlrvo2/Nblz+Quln7TVrYPv4la4fQ51PhiQhyR+ezzq3AmiI
Vcv2RNrfNu5GGkDlnmzfjuT4ht2xcPG4uWt1KBAGJOjm656L33Jrc9xQdtE2/z2e
/2Cx/N5oOYWD/y8jhWolRoqT6K0c1y0qz1bERHv55Dj6zeXNYlXHUEWs3SrIrD7J
nyb5mR9aC0AC7o+nv0spPYRe8vBAwWwzQeKvxXCJYwUJROhFV5fRJig22xDFkuMO
LgggMJIeExL9rwUYTKWyvo5k86KzYF1+8QYVLsQR4pvTJTBhdsehBFs4rLeSIwPb
5sSaR/Aw2oSheUDS5IML9bcP1lWFIFRgpi8OkyZDI6I++Pq8g6OrJ8k3HuTc8CAb
QHo6JCDYKdmPS7TGMtx1IGtrfuiK/4MTVPsm4htF2xdZIQNnpOnwG8nH9u71infK
WPeNnlG/Y7mHzgEQ8cvu3Tmi9pVZsYeu90IPqWQ+e/TVMgGCY70LW7DnAPty756O
4MYs6nb8ooD7SypP1pd1eVvRanY17vXE3NqVno+O3L+o4r8IEXh0FheYHZBV6LS4
6fJ5je/BfpqWPBV+9rTRgQqI4fJFc2Nml6BuJJf28dY5hZR3AbEsCpKyF5zowwyY
Mbow3sol4MhqnUoSH3c6Fn2HyMhTyzeW7yPF5beNux19k7LhnH7CRBuVzchSDEUt
V3te8FJswm59SWa5ijYwmf3TDnKm2HX39HTYHS2mNUPtWI2GJqyiybur0tuccv7D
j8kwfUE08AAFcBHniKENIXkP+x1dUtIUaz+6ULgIQp0Nos+mnVIA+Z5bECebS5fa
aNVSQDq4NGDkcL1v9X0FoAIcMI1HEWmVCh76YlGdFmAVTXU7iavB3/tA+cGmWXEt
0wrIkGrWFC3L8+IjzWOJJluhXMyZwQgI1ET+0Kb1HzJAuvJ7KiTEX3K0EHFNsEYZ
HWEA6LN9jw6R2pEwl/tE9YbECvQ1aXOG0V3yanGEs416GFddVRhPsoHlE/blEKh/
6nEe3qxX7AEQsqJimA22IXzJv4x0OZffZ+XquyUVjWE8SP+DQhAtlgHMQJjwboqv
h8gBkP4/L4wz9WUEKR59mbni1j7oosrAUa6W+CXbRqshGhxB7ULnArJim/XKg1PA
RwaASmVPncisrlz8otva9R9OQjamkxck1EnacvP1/O8ToPKUp1MzWKQJEy2Nvm6R
HpZ/PUNe642hrdn6r8oUXXj6zVYreD0UQtU3ti5E+nK7UgKttSfwELYlffUzJVk5
C7cMYecPqxwgdDm6ICvOsVGjYJO8wghXgfSXuvUW+J+Go80YeI6pOMFnjw368K5b
uJdGEX2pEZm0kFfZKwzgqxtCjD/2mUjw6v8BzJ6oL8RsomEfTdgeaNIhhuv+Nwse
pA4yy62Ks8GtqB27n9aVx3pUHvkcGqshRYWCwmfxl6W8kCZVm64c2og/a40SvSuV
8QCYFx/5SPEwd4+NVe84soDpCuAImawWbLLfbN0XbDh1t2UA9jSiMU+UkYgtfCDV
Dj8Xmw3za4IZ60UeNGX8CqUqPHl8iPdi7Rm2kGqbePpPdIfAwVMoAvqpsOXxvfw6
sIKtoiTqkwptzl+jfEHIZxTWIJgRz4PvdWzv4cL9irpjbN4RObptQkdGRwwh8alo
rHmNFxJMmXP5csin0552NEASyPw6JYS9yoiVsUHiYq96mPB5W1y19ZpAax9nBBl+
dTUG0sqfG9KljOYEq2DeFV0b24sdd0rqzLSEYJ6JAeJnLU1Mo9o8V2rBQdWR2YVa
/1K+q+2KvqOnH8rpq/5/ND9kCnOA9dm35qdEvlF1N7MPKOSPFLuC9u5DOyz+c8dE
RhnZ3wHOdRXDHgj8S2XRxiTlTqR1Rn8UO4ScoARmdQxHqQUElkTy1CQp+bVfepJh
oTcDdAZgHTV+0HIrKhNO/m+ZaYmV3eR2CWKu7tLbRRFw/m3GbcK8NQOoca1Uh+lH
dQnkFeDahRy0gwKUQ3MMHY5X25zy1lxi2Pnn2YL06H/rsG1yR7QeH4z5lqcPI3if
Ck53AMxkn+4rDCgnbG0P3IaAEqPjbVvt5uAeIAlUPdDbBaevVUqXvdGjYDyht+90
bavNTeh6mfADdU+RkyFBFA9mRl1LniA9YlLc0kVdlbOOPUH+qlr+UXuCD6qdhkPX
MHkBKpZFa/bubnBOEZpFtKMnVcVcjCosfiDbTmkTMbCPO9UBzONLmfGosLKsc83t
3g7udVlUVlowgG8X8SW8FGT3St1S32ZIEAUoKoYn6I1fUpELytusmQPQJGikscum
z9k41pJVE51qRHLocrP0GQKEBLwc8Yc6JWI+gxRv8lf19SfL+ro51mOfdVCqmtOx
yBNbFvYjH39RfE+qfWS5V/XgbACXPTcIjcCCh2WdsJkNX/JOCQUxsZSjFGuj+6rj
yYvINb8C6OV4ZbiY+Xw+lbzxhICNtZBKXrEtbsYNUiiCGh9zLfcfxEsJ+PxlVCkr
4okUOIRNP/7Ta9iC/SJ50Cza1Px8R9p8fYt1WcHg+A9UQ0Idmvt68KEdzECAxp3f
QGVMmmUs3fTo6CPvD9yeFYrPrbZAB0JcFOx1bSYKf2hLkGfr/LzUK2F/jyd0MOPz
kwsCB4V9ePH+JPyL+aQ6nmQgHfrZFYKOxJfVMmKadrJlEQfbgdzXv1whpa/aXz32
RAAtnvfov13GZHXARVnixIgeyKnshy8Vc5ZOXQCIVcVy4HuDDQzxedufy8Yxnu0E
0aO+KBdxDo9BYNqv5GRD9Y3T/eN5IiiMKymhUHDIXnbYL6Q57/DPOBon5OAOzCeq
utAkgjk2+7gHwL6qNGxqnz3z1HWlW3JVunbJ+9ZLyFoGf0GLSGAr2ixtX98oDK5L
4TsXdykYb5PHucIADRaVotDEAqt77A6o6v2kmSXkDg7WZXzcdHjlRNDMecFkmywj
pfbBBmCM62jB5rCj9XlUImb0so0hOdhf+qtVOuUtOhoWeokieyjzDnMhQ067gnc9
+s/pM04tsvoNRhWkRuqOgjnquBATdjrH6hbiougo/rtzPqvUKW6gkAroS0ys6w+Z
HEDNlKsZ3Hsi6N73Iks/e3w2i82wAz0XLvPKXAapHp5hYv9kdiHUhInAp7zM4kNd
PN5/GAc27GC8WA5Ei+ILlhhJxGAAPdRLp1CxLoBU+UL8NsWR4695vwpg7rlu/trB
pjA1zwt8+r0W+HKL5hGbXdag3eJBPezBQKMosdPV1W/iKEFlNy2niPeE98zsd8eC
5h/hrg3vuK94Nv8ds7sLPwjG4/tRAbCaYMOy6r7XAIpMRvhn4LTJfIOIm/iqpRTd
lRJWGzgShQRlK9kLNyMTIAnLf6+eOSY3pukp4pMhdqZm0cL5p01EipJJtaagkxfH
ATCuTjwPIMaJbvx5AX5Nb71T8hzekjs5VQQ5Kjc+6fHbij74HP6tTOs5x7jsD4qd
fnlrf3bkByJyTNFTRRyod5yGVk2eygcg3lBfYUilOaDV9OCWKCpOSQsi0RDAF9/r
veXMp/ZcZXbQ3Ht2su7EXsfMX4+Zk/4nhvq8ffUK3tmGQoi4oRQuJBkWoMCWb/x+
90d1x+++c1HIm5luku1gMJUx6TvtWTh9d9h+vmfL3RKNwLDDUcGA5LIqOTs4DQwj
t0TmZLYF1B4vBG0E/mNC9pH4w+0BHkv8NywD+bG0F+Y8lQ9ns79cmpKFRJvY2TI9
8dYAcbYjnATtWkmT82OIE74oi3vXykRffMYbevOrsC2dOxJZmYLRlEDrixCtUi+M
o1lgN7erxH0QUOUkGoLwNx/Cx257CQB+3mv2snri2Jzr2FXYH0I7OgSVH0SlvZFR
fXWfSFCUIoPUMK+99iJ/cO5h37Sd01zuvOoR8RobfVLXwJMcZN0o41EGt12ls9GA
HnNDO6Vq1hXxtk9SIQmD3dA8kMxSl1EfVFGpMUn+N6jOEBLreNlzFsd54Yq8mSWJ
FxWStNyMKG6yuhsJA9v0BzKpWBdIDYX1zzg/5ScPUaa1Ywa5VuApkzgNWUAyX+Iw
sbjtwgWMq5v4FZibGWnypxTydjLSxjhiyvXY4rhYPoLS+iyI8QzTMHWeOAy5Nldn
Ow4vzUvKUcSu/XNCinMUFvBB2ZDNJro+q+cezGhWAa60AyVjvGlNZDmriFe1X1ZV
XBdomLX3w2TUGsRbTnwFgIt5/sAmJgUpKUrMuaPsrjw91FCnbnLBvKrrmLSsJz/v
skighF3fF98IZSkfaJm+tsLeR/zcITROBLVP/7edSqOBQJEWUpYM0tLJ7/VVVDfc
pe7tgLaeAED1KaGQuoMCOA==
`protect END_PROTECTED
