`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jCLeyy9RX9aQEygfHjbBpSEEaaNygLFv6Kug58YHeNcz8Vj7g/n5QorXPAvp25Z
2D9Hczcw4b/4oVxwqNeDGb+46vkQbNanfHU9OtJ6I2lcElFWRFjPDBvWWXy43Fif
arfSz4VdDQOKGumqpqLXEs57X6dY2F1wCRXaxzeTZWriVJWefKQc6iltXDd8YtnV
mEIHbebOIKMIAtERgzOvYG8/OtZMH4j8fO/nnDYQrfGRUjj+i1emM7XsSA0J6iLG
4BCP2K4uBQRxdlCc0tZLdSPKulOA7VC1zg9GSDJpWWD5THHStV+asqesoSl6L1L+
ClN+iL701seEibZ0Sccq5lx6zsL2b8tmBcIphbtyseF2eGCB0iyzH1R4sX5w7Z0F
2a0/VCbSXUOxce8lMkbZbpZ9i8ydXjvjaMaLiDMYf9mbvQasdWiIRroG+LzvQ38D
Kr5hgO0AGQoEH0+AUcae5gLNPmQ1RA1Uw+aRIq0Fkzx6//QeR07QiWkFa9X5Amvh
Vd/i+IzQTl+ouIhAxF2us3YhN1pnxmFTbLNMq4I+KpWwuflxqDNL+UZLgx2dhBFV
0onU+1I9dWKxVugZ38roZF9D22mdS6h5eBLk0i5QhDTOqshLSi+dubYort8DYbmU
leTJN5XSYFrLoLvgjVZ9zzlTrMEdO09bLjVMEHlzcaJU6u/IaDF/l70VRYVfp5dC
t63koc7WakvkT2FFbvVymGi+an1B+iQX61JoyVQBGHacUYCaErmVHRCTz5jwrX2T
JygzVvqJ7beL8gNgKYoUEc37ps0PKMBbGjMwRfne58GL9mVfv0lYdpTSwB6lQCm7
rtN+U1IG468/mj1pwAP30Ts8fm/kA3mzw9OPtvTe+k5Xj/3Qef/XobYtuM3pz67k
flU1aXC7Hlp12/4SuOcDwGnrauvJwg5XJ2u0hsSNnCveEozsqBadJ7jvuH85bo4P
+VIqyK5EWPwNrG9yv/AC8me2aePWRoMz+Ftu2vX86dU/ftQehFUVNtfTLKNz0hEs
hwOV7WicvU0PhjqAvyoKXbtk+aN0Ka9mKSHolL2LCA/q1NGJl/JbnMgdFRknd9i9
2jJQcKemBQu5N6FdALQJHQLbCQZGWZ3udRBRRzP+hT2st3NqAQxqXLvXYKrseuG4
iIr3h187uubreKrvmmjqojsW4SRH1coom0QXulaJQ4PeoHGeMLX4EHxLTM9NOKM1
MTvnzh9Npwv0aNam6Tf3pWd+9FbiPzpTsKp5L/fx0/QZz3+8sP/a76NSBKdGWWME
A1cP8ffdDrpFLSy98Qx9ajuFWHrF+YtUo08EmdkYlMaPP7EaIvLTTaCNG6ao9GHH
anpymrrkJwzjLX8qQhMAg1mAE/wR48CRMGmaf+1j2SuyDskD7jl0bJzsf2l5cXNq
+/8XjiAWmh1ZPoVkWpWvWGE7PJO5A0HhIOydAcsptDuHVES8bq4MyA20GipRRpxj
ks77nasSZXJ39ABmLUDQanhX6Shj7tH0SXaXb9uCY/88BtNbnkO+dq7zgVbzLRzq
Z9yEjCmL9W79nbaYdmxALnFZKU6ibcL8sOk/WQ1A3LHD1SAhIE7mWkVOlexveeGW
RA0QF5gGv2GT1rX9V6sQjs7cjJAMvSY6r2P0kvCyNcVreFocIAAELFbV1D6PyaLg
Sw4wauDSxZQ6QdV1uLRmtnQNAeOIj8RJaiMwM+GxZ1wVtucTdX1dkp6CgYGqf777
NDe7dKWDK7PWBbu9gSPQA4x2OzpM+HcV6WlXmTn+jC7K5C9FnoLb5Pdvcki8wxj0
6YlQZvyOznZawumZW7deG5ZHZi93x1A9Q0EptFBqJW4MRas7YH/qZTwJOb+zXzsC
6ZFXRH7tLcdIJzK7Nqa57EhmF13UTRyhKAqYoiG++RfOf0N8d1l0asqFapZ4L83O
6MqRHLTEf1VMFX5Bs8osAyvf6LD25GOwdJSgh2aqy1GoNMAcvjLTaei/5h9MZQ5P
p4/jPLG+q1dvV3+dU0W+ZBM1sxdJEgYzwO22xomcuobVbOY3buQv5qIU3ZSVec+f
naEtpXsm3UGn4m2seE4+cZooGtqkmxxhbWtbdtdH48uiBoPsyaljzr/phfH1gIih
QlEeljFpk/p4p6GYnteRTR0XUbGM3pds6Jdjo5T/oBVaWoM3jHNfBxgjItYsq8V/
Tc10M9cEe4DWpgUckuN9A0c8F1VIwmhSfTY34jEEWMG4qxO96sWKqptA+lAjhwWY
zZzHm6XI1MzizUSOtxgEZ1Qsr5zU0iCqPqytMTSPkfJEnBYWL+n2Buz12upxuRNL
Ycuxi1Q6NDaq7nOyO+56WcGgEq0OvSDzvsZoj/PU4UfPlbgDVJkxSDf/Nop7I2RS
rIKqwZ1CBUL/cJ46uzpzqSQ1q5CwOyhuvRUEXeZ/rQZHKx1pfsPZLvmiXP1lFV5G
EwX8cIH0TpBbLChZt4R8o4zq5vLgk+yzNL3hUTXxvWAZK0A8CSdpTsGOY+6BmmKP
eqVQFsmT8xMxBI3KsOIhYsJK34xaT2kfYl+P6CYwrdHitM3zc4at/VcnWWppXtIp
bQ1J8XNKzocgsRoR7THNuxrQcyrfdGrQ0upJbFYrp0YFXKmd4RS/+qKgaucSLkal
3KXgpMdfXIcWfc6TFjHth8jDLk8sMSrY4k213J5YtENCKXkPnz+o6KQGqO/3VdEg
fZlIUI3KbJbfDDS0S05OxkMjky5S7JIEcQB8zvOjn+ww5bGYdHfQo82uxiUYcPCS
KUzSTY3b2ATocdMP1FyRArD/+bneKfhZgLftAS7eXRmDm5F3aQFsNI2YyBKorO5U
c1E6movZLfhHlcXWltyfRmiyTZnRYBoNkdqUC/3PZVb7d0sU+RD4C5GgWIuFvQQ7
Nl20Mh45nWgo9dTr+duQzK++fl9EWETowv1OX00ZloBY81yJIF0EHwYdvEUH8ins
Yu+MiCnSE7UrKvcknSZZCGai7c/ylqJqjpPbVl4P1BIOSm7nyL2KKhtzusTmtNHs
JifDihKVXzr9NrkXFjuwFsfAtajZnih+ppji/5EdqDUwzwoTLlAThWgAPCJNhmB4
2aJJ00dJsKRYWYAQATR2LQuVCzu6RJzjbWOOk2wJqDgM8GYFfxJpg3eGGHGTFTA3
iku3BVYRH+p+XJKrZJ8Zy1gT4SRFFRHjJyAEmJU0XeNdGDpSzpZZjDReItE29onp
KtXXVPgv4aLXTPSljmE82o0j0l931c7v3YxZ+fQEDf9sUwrT7jP24QvJMVn+GNTi
yYZ5OMUvQg/nG4OUOmVc0Q==
`protect END_PROTECTED
