`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ELQ8Ec1KlcYi9PbvHESHPBohBJTW5Ikp0dJMBdPgr8Sf90ljlxNVrimgEpuS7NDW
oQ1b8+C8gvkdWxw29HtV2+631yn0MViqZMIyJmD2ZsJUyw8/fwpRpKSHqyOBvVO1
jZa4aZBhkEwMiD9IJfmLwBfdS6wZhQZdTtr1gGyfcdZPUroWj0CrUQQ88rs4OgiP
aWmr9Xw7oxTCf3WRCjClF9B0SkFs4wFezpVGPUtOzlfyVuPVest5MlL2xpQdDB84
rNPUNL+ci408P3oMeA0gwQ87Lst4o8ffN9vn08DaNL/ZZ/s9VqtZr1B2164zfCnX
KNF2DAFS7obOwdRl51f1jAQpaDvS6P8zR2TzCcFOa3AypBvOcwC14yzKzWtjuBjn
+hWze4y+Z0dpPzEnVLgAB6SUwXvN7UhudMLGWKgoU0ULGFmiJuOka+h6WTrJBQ/2
8apdP7WMcfAOCRAp3sR16SYFot6/94bGllH6c9o1a/Wi/jSJ8VX/BFk8r+GC23zd
thyW6/OrGa3IESZImNqgFgcTeFZnicYd56XQ9YjAeL4trYlm4/CcN3GnICDB+h5r
W6uEbhTvT0VvChJu5lwYpZeqh+v1VzP5t/AKnosLJKELNhEdjVd0Rx9TXSW9olu3
KFmPjotCsMtbkKtGtZ6l5e4xhBOaKRAH4DTb6QVc47QWOs4qXV/4IGagawYarJup
zsTw1fwEJNQCirlIuIBGvInzjNMFZ3RKCqzPAJov/bRs+YuA/0Encyx8tYmMzdXh
MsSKHfwymYgN5yWWQfnI6Yqqxy/NsX2N29UqFVCZAZTOdW58d/PZGics8csXGOF/
t9gWNN3aDmkDmMCI+c9B9NS8m+1Ew8MnnWKJBba0vbUgcFnfbvg4fXFZmUpEe6yJ
IVqP0L60MmRNVfqVTKbH47pMZ2mz/HsIlGpl3EIruMVTI7o8ynP243hwVTdyb3Lb
++sFjZLnqZln0/Nbgo5innp6xBxPBfyuHC//Uu8bg1gDqBpkFQCBFW/jh3p6E8YD
CZLuqSb70D+GQy1f8FE5ja91pVcJIYtdHMhazPGUaMU+3t0v5kxsrXkJJp3vtmIr
yslWqw3Oa3d5fJGOFAwLf+jkPkWs341WdFgy7gzQirWJecxFfuXi/Ntjg+54oj+R
Xb/Jzy8bMcFNFjPClrOLNjXz7r6U7tDaKK+A6GVya4H4KlBSadGpuizZO1VtDAps
cCBCWjte6gUmEhJlNihZBQzqybJi9DcBChWGzUxtwe1QzRcdMInnesqeQrxd804l
HlW4XIrpNbzye93mSp8bnpD9w92hPSNlYNhmDQAF1K9snXfBo1ucvlCrz1XR/wFY
vXogfDn8uZU44QD0HxykHK6h9jKem70GJexSwbp12Afb1kvrJjSW9nbeXPagMqrW
8ee5z0vZnN/8OKodZTpF0LTUJArscBl3j3NCGB7Jba/dEEhctqj0NF+yRI8BImCJ
f7b1v5bGZEYezk7DOCrMJJRkEmnks8mWeeWRd8J8i+yc80Dm7GR7MbWUr4pjB+oD
3ONunlao9uSjkAnecY2wbWY+q1d4BfpMRKbQTHvRArD5HugfGLu9oXWj1M4VbToE
SeU1PKUUbcGnGOo2oqBgzica2DpbkYzri0WKRcWXvlXisuOKy1mqKsr78KyPzAO7
LFUcov4F6+HhI9VMpMxFaeHvN4q7jsan7v907YFtqof5kE5o2mZQH0lR2NnJAog6
PCcafqUeFjGFYgzNYipWj8wptSpwKQh/0raK/G8BB7HZvDroyvIK7kvu5S05Mcyj
8qIzDMWWQozAY9aDQRLiNUVquVB6yUKGeqiZCJ4n6pV2/hfnnDDRKIyoEKkioMZN
r6BjCj4A62wezYT7NIQYLDGxJk0pyVMQ1dWcPijKouugCXO0fS2snFJ1LVnou+z3
CnKBtiAIJRDZMiN8RFmP745LyZmy7XoXmx1gzVmUUIa4EToLz8aSg1XyVU/meIlc
DeO0RYkg4ux4XfO0cAr7krt4HnI3y7UKTE+6VReV9iFAptSyMC0cJOwJYEmwI7WN
WylLYobEa2dmaUxbhnFKIqJpb1aUUMraQ3DvA1/p5QjF+rv/9vUyTt38jTD14Wg1
4+JJUjdKm7LzSYVjb8UNXbjV9Pbt7uCJc/Vgr8pZqwiCpA9prts9++0P9o7PxYMW
pmT2OP6zfrFH7gKjTUq76pvFZyRHKjwKOcPSW7LcBxNMu7ZOkAh4BD+9E55bKjmG
faPAEozz0yIowQNrOXQXR2bYzmKrCH4MLeOq7N5D6eKFdhvTpd2zWyF/AFUnc8VP
8v7AM7yeNbomD6P7Z0drBp3ueXxWW36rVQwigEi5fo8vIh5TjRAkSvwSNKsukpnI
QnwO1/ZMcUdT57xDBVdklDHzlBsdSlMKY/SiN1K0JZ1FC6EvTtwRn2cnt/vLuFj+
XmLupHzNIy2Bssz/rXDr13ynVLVMFhdfBUUd/g/yfmuSC1ElU7mypmTnx7AmTckA
w2yPePz3rl4a9JWXbIZJkg8pt9+e9lhb2PZfc2gAhxJAok7cU4zOVIhHL0IF99ha
Z6MtJns0AjMWeqTNC0etcNzupj6TuFNicUuD7m4gPHSPccFrmm9UBtasJAAK77XH
AqrKTM9mzlwZ0UEha3VRZK3vQQG4gXcON0MfHkptukfpOLknGRUSlZm4Y1SpVJf7
2/JVlQZzu41kS16n/o+RlMfv4K7nxYRu+n3wtscWo6kDngjHu9e53kT/Vrn9LN6x
EQMmRFbkz5KDs7abxxvt+gwAjVpzikgcVp0d4xHoIuyS7peFvcPkaKbfehPtO5hi
odDlF6jU2f58gIfzLfBNgDoljOGijPAG/Ky++LT6bVAgiyG3g5BTrHzkpLdkDcGC
mBa5RjtD2m2eJH5I2Rfqfzjen9gaHGqMXiYgI19Iq3CgiIDpk9uVmIlfEA8NtLSF
/1uiNQw+LiPSN9lrde01Ttt9MeVaae5lfXnH6fI+gqFvhrgEPAGtjV852T7sVs7D
BVrtqZKuFMfVFBNwvsYdrPJPzGrCc7Gd/Axbc16YvysX9zofFgAznS29Hp8NIg4q
m3xZ6KqAWbzqLpd3nup2zKPFovt4uOlO6oA+eYxgswNGOEWmNORsH+21+S98uD3l
wOo0VK6EZIcw4P7Mi89NLjBAaPdyRGf+3NjEZiIQrWurdo6WcWVgMhC2qsknTsjU
gv0M4SWoocFDGneI0eyE9BrWNRXy03avxf54FTni1GJRd94G4rXDCW0lxezdhzVG
WrjX/UAj1gKyGUYz1cBlEc5uq2by5ik7OKWDK6vYEHDNtgrvg4YTuYqdx6yJgiQG
iaXKBm7iQKTMXZzYIKIL4raNZdevBQe2lYonfXPsmDQda3Tq1PWsbDQ6hY4OU/eb
Irrfp+DB9hhvwFUk67O/Z7a0APX112Yb3DLSmYCgmz5TIFPK21dhV0D6OXh6Eiqn
cW8bZ0Vs9fv1+ybpCqNKWsIFmPTeEzqr+1WH8yRG6bYnjvHTtzV9WdLD2KV3OE5J
onZLRBOHTEBB/Qc+yvf1iLlEtYUhpBDP/iAI5K60eeBs8WmwwVBMBE4ihHmHDg7/
UDqHQyd/plPDzR/+KmAt9a2g7DWrP2oGsTefgGyaKNS+fK6Uuhuyh8prnI3zb35G
H/08/ARrJCArqMRugapDYJgfPFXIZN+4sm/VHZ6NMmX74Agf5SEY2tdBDXKS5c/C
fit/6lKXyU5lE6XGLx6390x207XdGqtYtYfQNP/2x6BDbx0U97WvGFiRvExaSfn5
LSUvsnkfDaSj4V2nQ2YiwLF9LFpMfJlas/7JoOSD1th5TwkgTmx4U+FUfF4fR1Th
nf3xtWNaDBAAdnEtowzfJwIGNY3e4adOEgwIz5ukZdf8/C0TpWnJFfkNx6a/vHaX
0QKHGYKQabMaGrtUdGc6FRvuY8IhnI5VUuxv+gjsMJDOonVFS4wGkt67m8W3de6Z
0QZKj2F7X7Fx5bcQ1R2nflNUHL9PZyNMnxs+U5LhrFP+E/TMp0X7bipbiWvnHjbG
dBnblsVDDEkQCXYuKecz2Ppvm+KDk9l7CJTe0yLm90LopPxmWo1MWGrloyujMnc8
/kr07FlTWG/Wkd+7qsDAiBWCPw8WN9MZ82+gSBBqGtfGAhpCRo5zWzlhcnv3HA3R
fHsZCaOwfJSkYEcjEp0eOypGtu+Az/0UQPIoOrE4cy45Xu3cqTFWVoZCwo8g7Erb
jCn6CaR417/e8R5p3bwV8KFjufYtFjYv8rUgBozfAI9CdjCtAGI6Dc9wBznNwl0s
XePxW6+cJKJRcORhAsIXXVovpmgF2OhIfazZjbZuFaV4O44h5h6AcF5pSIVGJpDW
v9VxmfYV9sQSm9OvNQNu3qHfxLUf6Ew/ScrvjKhqCwrvUI/3TRdqyhuenWW2LAzm
yLczY5XjAS07TBvrNAj2Tlr0AN7z8zqm8boP9jxiHuMcW/R5/ZGXxz7vvz856fkI
KJSmntmbfmy0yKmUOc1dBWMTDeRju/Mx+KL9UBX4xP95D09uvhgubwGizN4LdjBz
BjOyNCFjac0qJnZLHWkUEaHAZBgYEospdgr3vtYlXPtTryHqmFjNSToXifNo9Atk
7xzRHkutg6aQTfkueOEKgOTlwYs3Fv1AjO3UTzqzC9OCurANrkCfJ4brydiGsJV1
DZn2OD2ECIDoGBlR9UUm6MKXkVbpJiC3VpdoXB6VvWaCClYXF+xwqsV0B7vL5MJs
Vy70wJBhZdDc0X2i4AIV3CBranE1OQ14ZO+RgQVm4nvC9mQtUZEtqsSRug7tsCWz
zbqKnLAmVmL4kgV7mu/DaFbtJo7dEJ35zoiFQggB5Ac8PSLyUrRF50GfXz9getPH
VlpVLmDYIAyU1Gu0+EKc/NK/bezonmsEmzk9eWmO2rCTrU29UBEAIJvLsFQIsByN
tC/s1LLVfpSBVx7rrUmoH62VrjrOjhHRDwKGwZxM8BD/na2LkdI6KY1orbtc4MW0
6CSftEVC5O38kNWkAI/u2YzxOI7oGuJuS6g0ZE2hAF5KyXkhqs4joIIaOdM8Hv6J
ikshcegee/rcYDSNQ9Tf896EFNi3AMM6MmG4oTzhKHOvz4nOnhbqm5gAYpDDtuXI
VRv7r2zoI0aOIhAtmrYLP9OIO5mzq99fCUdKBvflL4pl5KGNiv9RxRBh/RYkCDRh
7vctySF2fevSOoTtYG//C3DX2fpFjL03jwfBT/xK/nHtsoPaGdSZCeZ35TcAfMED
w6bwdshxE4bJl4vkkyVtPjqx4dAVepyZHDjX9VfQCpMdlPefX8BTGJmwzZE3BU6p
PtCeBtZWwNhQXtlnAehP6LOsxXzRxgrF6qmk0MBdyRaBzUHct+4JmTcDmwh1ahI/
OUwFiPWqNN4CBk81BRzoNayvbPN2YMQxfDntSmTukBOf5NvSn2RC1GRrizP8fBeB
Zdcq0ABSPmxkahFLlZ3SvKkG3x2v6lVNJ3SE4F4gTtCe/rZMz/Z6NMIInzaW+22c
kk/F1tAX92n4Zrrou/yDSTkVvElYEtlckVas+5MgnhbdxtmKk2oScLxJ7ung48rX
k2l0DIaE0pTbgoUmhMtbpTfcZA7W/+d8fc3084+TIgtkz3e5vZ3nsiDZeJgpwxLZ
aqB5K7MuvhOk2uZlMqnIvq2/SJw7wkMiIkMFieb7/tAA1sPm6a61wKTeDJGngnHL
zfbJ5G21SuNkTCIdZX2kZH2hOyRBfkSjA4MXiHdNE1qpk4xwDjiWDmfIZ+Tc/5SJ
fhcqCAWKrKs+fEPBAuZiBcyogF3zUnoDWoDgYRpwWkv3uQHlbbVJSfLwJWAFc5Xr
/am+3+9hHbJCd3w19T3QfMfpMU2kemp71QvvFjpjKnD4ZdoGK5bI2gSo+fJ+hy3Z
t4WBn52lpFdWLGCOXI+NUcWV+Rtu64s7mEgdXIORbnxqscAtvAs+mHjaFWFKiRQ0
UkYlSsF9l+osk2SQ5ybvW1C1e6v5kUfdYHkRaz249WdGqABEcJiCQPXhxzCjdKZV
DEnO70N60UJyvQxWRYO171wr5S2zaOolp82CHxcvDwhfozHWaSOnKsRLVsME21AM
TlWlkV4EeYGre/vQLK5Z2UiIS2GuhfvcHjvx1ZtRjDIDZQ0vaz6fPQy5dnkz8XNh
h0j4ZiqLN6GBRlHn+jV70T0wH1zsm0jSznr8KCOcLAHvkEOrRcPCm3yKJbZd0WW2
6x0VKQvWGltQgpo/AnRlNdi/shKibzLzC8uHZ5bDaXF82jz5S2DPMh3Jp08QQisH
5UCJ4DYeqHNzhzYVwI3bP62FJK1UgQBPcy6aynMeF2cd58v/ZuzJ5DKtmkGvGEVv
R5EEvlIVLOVaQ8FFVeR00ihncXcCJ4G+7SWnLr9dxnZjUaArGvXkusSBqqFL2OtV
cSPVx8oK/jqvs83eXAvdssMOjtiucuPyifMzqZvGw/Xl9M3PRV5JmUKQi5/ORK+f
fM6aO6U/fpahS0q6pLkCA5BYbMT+z66WFrNzAmqS/CSK02c0Jmg2p+aqZV8MSdnO
1JIvaZJItL3It3ifYUOj+cPo9ChYroe5V1klLmlY2/Q056uOW1xB40ILUvucR4LX
I7LVC8vIJqXt0OBHSXNpRpoX7UYIQyNyPVhFh2mnNcY46C07oIaaRSQm+zzluPz9
ZZl/PCqeQkjKATOOWGPhiW/TW62oMOqRLFjXDy7wvDT5UG3Jxdh+p3G2kF6eA8/r
/pFg+5Ald5w7cG2corUgqoJsHD5Ljte7qlAdSQMj2/i0HqXPMuCbwnuw+Wjxr2uU
Hz6ghAHRuceVahLiGUWD4Zj6ojQNGIXhNRApTM1/Hx1gbVCJGXroEljK8GtCJhFv
1getWSS4K/DDWQ3iygi09XrPDy8FEdJXXEByvjkLGpZFL54a8snSOh32DNg45HA1
S6wNZNUqgRKNQ2AqZ5D1UXAVP13FxYaq/4WI0XLkPr/EoGt+SVjuTqFzkSXL+BXa
C7VTzuC6zbFF/nOtdyao9sstqzXXkjWJGrIX2/WqNymPZWj7XvCIwywzuyLSP3hi
9xCMiMRRZdXvB79x8N190Ax22aafmtHX5S85eR2A/OoXUR8WbCjZBZK1l538yPPf
H6gZJsRcY4RDyXEs8NUGpyNpH7eEM2G2jKqVCNDRLcBWdyEK3enqG/a6xf3igbOq
XvCxlP2elkwtye5MjqG4jV/u7fPcLpMwm5J2zSOtcgk36xViqqWOlfA2PajZMj/+
BBdG7PQj3ZqiI47qIwwRlpACt1Ba0SiXGA96n6nmlMwnWT2BOI+z4yUgY2xwAnrH
vlHmoZJO9UshOh45qv4up6K26kDiH+c7l3gXsF2NOyrlfYDprVUx8BRFvOAZelMi
UOJDGPm5Xzk57dDNYZLDsIhDskruKndr0We2NZdyNprYzI75WzwHrjdWbmNV9KfR
B+0Tv8MMK4UaE+mgVZ9NWCZH0MCtdnPSTZEzuywZHAd2fguNWmLgJrVQtjDvkzgM
KsSdV9eewqU5mXb+MwPUbbrZS/qBaeGNGjyBBtT9zrPBflROq3VhPj3GoYzWqg0y
bGalXnYArDY+l2d9MZSKM+H+bBG/7Tn6g+qPpuNIniac8PgZQgb7K4Wg8q/zUl9G
6JYrZ0lyYmJBsx/rYiLBxp47p32ppaWWtKw+VEafTHrucdcD6KO9zzoPICQ8+UpO
0wvlxWMO1Rj8VYfmtdre19Kr4GIRgqqMSjhFGQv6X2/6LBy8csxAE0AJawJ+cJzx
5jfoIIlZRTqfUjnJ1bkvH/cRGkd49ssF9X9lFQxq8Rl6lC2GiHbB9z9XBgNnR64K
cDBTn+d6Kd0GhHQdKp8eLqtPHdX8GkFvdQUWlq3zE0TQIrSS79qqCl7awk4MJEzu
w/v9QIi1nRXq5NBxlnxUR0MUKHr67G0kLl8PEQvxU+ikBESA+cqOUhMY+cupt28H
Yw0GU17c/xiRNjDjaQgkThqOLJ0xm/VyYi/LXJiuGVEeIM5CHP5NflZxDuF9LxVE
0ex+QbqD+E4v8Nt4BFe1jIUuD49Kr29sXvWHbuuaRCkqQ2pV1nADlTRTjmvYE+OR
enQ5I42aL0AB40tZ4teDTX778a+/fEA1HNrDtO7Zu9M1OcQcVOYw1JBtdIw0GisX
2VY/l9dx0oD//8/ebLVCvlaqrVdA9McMEeS/PCt5MiW5SJwethv+DWnUp8mJXUKE
7GtXt4r/h9nKMRUcnx+/3vcgFwloF8jPPE+Pjm5NAvH4AiA+uflouPoZIWWhQgD2
bUjBRS0g50+Kgpzqn/fq3RnOQz4uuNZJSO6dQrpyYJU54QaCBB0bHhwi52OUvvoQ
oYGxuzePtSFwFCEMbsCrGWmeHyMCB9I5eLkhlx5TrnxGKokEvDRBCmii4AmYHBpC
Jhqev8QhDDZ5/89kUO67u/CO6aqYz9gMDtoAMLQG2l5nktGwCYPhDxHW2szEufdW
sDy3Cd1ee76rnXDwJ/v0pkCe9bjCxyh3vjKnxKO1c2fnBFmlWrz98bahThxKPHU0
t9WamANl6jEMsWgbgFjm1Z8F7pKP23+lghedCSJeLxzKCsMJYS1JqQ54RI0ZhNBL
Fu1PFxB2pM1CHJaRcTFCQ6TKZ/zJGyux3jFIMqacM9kucXSAg8Ao9qB7BdJShpaK
+6wdHoj7aIlzT0OHr1YGdBBkkP8XOZn88pPXxy/A3tJB/M59lkjHyGWcSnsF1SL7
KHCSYdGOOSEN6K0RlDpqnw/QJ71hwRionNLvYHXvbJOHjmNs0N/TP6X6R/SHvtNp
QN1ckV3FENtK0sFGt2R2Os9IibMJaXnAp7OOKPWG289WWYYr+bhDdUUDiRNMScN3
7VpIB6CyjaiYakx4OugI+akLCwLeDwZttpUFTwlJuZhgHV/pCr4dkN3SHOKH6ce7
pQuWB50SebXt1aC+PjJf7AbpRhze6eMPY8CwV8E1KnBSsEq1nEdZ+N2/rqLvyzqf
pb97rsayW57O/U3fmL9AbfsCH26gz34Y944ANDoTniVHSP2Nw/Q07cfALqLWKzqN
9FVupDWnGEQ5V/lPDLFRgylQd23tS/hekRa+2HXMezwTA5zXer3Hg2UvNraYjWUN
ixnehOeUmaG5r/4FE6pYL+zeaTDDWNx6Y2dz4e2PbYcYV0bybz1LqbANJ2voQDmC
bmc8KjZqYeC7zYoPEe7Er0XZrRaCozjsfyPan/e3xyE96VhNlUnX7OzAsOzrbSnk
2SfZX9XyYvOvpgufwrHEEsOqmiPpigey/6gWyPSvsRBlItl1GqAMCVSH0jRfalAB
hyReamWjfuDAqcTPkdrT+ulHU777VyjV3STD5AnydRVZYvOTa8dwXGbfVfW84Lr+
qSdm+5caTgvLRlZc6NzMMW7NR1HB3JFVtwHQf6GCfy7dmbujGbWZvIfwMR9U5Uri
KRHNRk0yftXA74leohg/ZpwoEqu0DbM1DueFF9NB+2LKkGUcEhPX4COwPX2BVn8I
ZSRDcjotBSfosvjzHs+OKMZNQGYwCYY6LaZhRriF+/AkVLu+wS8CGRCIY8rpEwAu
Ul3Xgy0TwzIRURDgVS6hG20UdHSWyIs9bVJvARASuTdrBoas7SCMMoCDSmCu+FlU
FuNhBvK9p/DGET2d4nXlwbXHUlwm77iUXfDLP7B9yfEHlueWNPAgn1CRKUopOav5
IxqCZEFt9p1y10NdMwRJMbfL0ZFNfQicAuJxk19Eh7YBAWTkHomNHkkjetcS0SlM
SqZSChrdR0Cf7DUqxbBOxLzrEJ29vs7I0iDhyAy5mygD5Xb+n0VGOfKyGgrAv83E
k3VFWASlhN4Dv5P7bWkGjYu/T1X+3OJT/ogyj+bDcVE87XqMZfLuHr5cy6Ouz2WB
7PMxFTlQYSWQlleJgzz6TV7cFc6WmeFRNuiU74DOIY7Epq/b8+FP3TdwhVHFLxU5
qceJayOZScpD+Jc99s8L755j1LTPXlSYiwGJ7lQVQXLeUegW4HNPDhf2ra0tJNkW
alxP4woxi81w4I9V8n4OBPxl7+teBnE3glm3UvjepcyXrAhXSwf/8DPQ4R61J7mG
MoWepLJLHl7B7N5HZIDwUe68YgmRuu+prYyTE0dCCOZgxWtSWY5SQVZ6Zae0fTUJ
tK/J+UJPy9ARFoLMvHFbQE0pEAUhV7O79QUegyXHiQiprtuv2uwcRYvMTSChUxC+
T9e/LwIdGofTKpfkOnWNl5mbcmV1jAMBj/p1u6ajHnRtxFxzl4ELZS+6P7hB2Th4
CiqSKzuvNNwlhp404hqqa9fnuU3CDXFxjAgHIO6a45jK+lKzUEl+hLtL3bl3HYsc
xxomi0yB/V6REExMTawSRRzBZFe7aOXcpcWjL//aVR5u0YzV0vsYdg+wh1RB51Bz
A9WAgIq6J3nX1638zaXc4TtZsKNflacAy8neQ0fL+cI/t+yi8nQzQfKw9ss0T2WU
ak1IuudklnHzp8k5d2YP44A1myYSpvCZDzt201iAkGGuYi9ytZf9lyZUgcQ6fT4L
MDF6qHMbZJRR0GnsjHjUwX0/XbZ8QvfSWSCpK91UZlOGVZA+8+jMny6j4QLXiQj+
z5DGlL5TUKXHI2TXhV+u/kHcl8QPF+MDEBTFqW6u2/XdOKc04buos8he3S067Z49
96+i/BeEHtHJaDSg9QuvrQJrM5kVGk4fBfkbdlOBMa7Mo9/9M5+gV4oq+HuXyOBF
FoSgw3WKFPCZJRaQGTRpwdbqOfyKW3KMzAyI/Q0KI3wS7GlocNTzq+T2oKffwQ/8
EbftHisro8rICKGOvUIdyiEjmI/AbEBC2yZUOj+490+fGkQ1m1hU9KxFia4v3n7c
G3zDqQVYjbPLOHryArNcZBWIRnSa879e1UIpBA4wBnAhPRDro7TbGOCGqcEfYthw
i+3knecrC9SMEz43ZzSuMNQpFjv42gc83udI2FabQwoLYpqM3Ukw3m24JbAE/tLb
7YgT2oRc+ipJ2dat0Y4fesDDXpev9ef7sb44xLY/UNZFlq5uPSM4b2qTX6c00xxG
QTKWty4GKuE0oGj1HHxWh5NMo6wvUTPVydX04JF/XbMvj2bkvvbVUIy/ggIVkQ/Q
N3muoE0a2YN/Nt+4LmCk+LrL9xz7ppNvAjEqIz8uyMXkzt9Bv/pLXje32QLaP7mH
ZrPcj4h6j1xMll1JjhwJmsztDwSXB3RBtt4qUNerNDfh8ixui3sGKQFqgSl6javI
fE3Tlybvu4VYGk3PaiOhu/KvG92La/6Ba8iWHrJ+7j8lQWcgoyOA/9go+7qh9tNz
tmWB1f46+m40btdtchBgstsHyzd0C1yHaVXq9nGWzYZkzkTwkymBayrFqag31Zme
mOtl1+LcBopFc/1O/Z9P3cuEJ6R/3Kc+sDhBullDAZnkAc4lj9kiArwkQEFJFN9f
cQG/Dt+9KciUVgnxWU6bnJ0se7zD30CeGgLMJsCu7e+UYwjCvLmrF91xhmduzgbO
tm8RZCbqdcAgkAYpPSV4y5jqbv+6Gzg2Y1I5mPkwK6HfUuT7VqYPlL0LhN4AFy1Z
zAe2sfxayPfYF5iL7oPM8GxnzYLnYf5iw6wXqayhBx20rHXKiBV3cVJs9E1qAzym
NXz30CY0ls6dMLLfMfOc+Lg/1WVE46EqmUS4t1MKUwhW1WceNb+RciPb1eCr0k0D
31HjhEwztzbnS8fyxA+YMx8xgFZqDfOKmiRan0Ow2PQZJrHqPQGqNmhcyzmO3mhv
GNJFJbvbkPPSliy41zgsy6rOQA/HFSNFgQlA3noghErx8mHB9cBb3GFwz8i1fgo/
veSKbgCjYo4BfWv2aAIf5uDkz9gIEActyxqsct4RfA5Uso8ZK7UOPJiE77aSfadH
wwZo3jhZlTNPbKHisvg8po7ulznJdHRBstDyi14uKT1GoAZ6wfOwtHCnkbE1DIDl
Dgg5asNa4FAqoS2swk8G8FRBivKb0udbG8KCkllBA0Rxvuz9QMQF4f965go83Utp
Hv1Xs4l0tXqHT//LuSj85M33jxjqzSCKHOLLVckwYr5mHqILoDYc4WPqiPPHlEtW
H7Ba4++Mw71GdTgRLFKKu7aPL8AmkgrElIqzHQWeAx7vgMgppG/o7auT+ZwSYZcL
ocnhsBdnXAUcPW5MEIagEd4++4ieREDB89Uz3ot/bSx+eEyuw+0h4M276Ljo4AZT
i0dEgHtbPKWQU012Tys9ByArlSYGe3jtPNhPpYb0m+SM/cnCQRSy1muVQT96/zG2
Vfd3hBwOcOSxSRtnnjSy1kU1BQfdGefDfRSVKbQJ5rfG5proUc/oPTSSknbDnqg+
LJ7+Eu/J05S4ae0aYbLcDJ2kY2p9MnH0lIdwTvgelhl5bbIjjFcbBcEJQsX/jthy
nscbhMEH19cgreDFjBwCM8x5iiBQ1w1uJm1KzujEeNdTBvBiTCAvwWxEBbqVWqpW
8gVjVhWY8omsIIM17qu/3k9vx8HZnb1XCD39S0C1AA3aGoe6kkeSUoRs+7gNBonF
MUog+GpW0x0HwFqD3jaEv/nheV5bk3FLC+pUgkr8/uaHpE3JYxvAQjc4UTusm+d/
MOg4jlSRZVYSTXOPa51Gih+XRuRR9fIN3jen0B9P1Y2qXpr03E5qN8jUDg85sRLf
y4zXbX/8j0HkolF5zJN2DXPfr3wru30Jrlfofrbz74mEx3i5elPCS9CnK3FHh81b
3EsEULko5qPM4Drxq2WmcPoB7MM1uleUfZuSkj8GKEte/kaEHWh2NQtlDY8H8200
lkp6eB03s5WmaZKrKaXSikbPvnpopDMk+6Q0cA/gHNb+mZnIv+RhzW/Ce+EOZwn0
+tkJg4VHY1S8SNn0mABn9wOvzTOcwbm6Jol1l1NH/W32+Ou5HkB/Ly15NpZ+Nrh+
V7pD7CW7fqz9Jv3ZPPfXRbbUoMxHa+Mq204MDBrjM4kOtFCxtx3nV4amSC/zOTWo
k7qtB1jcjKcP32HftFJ2SQe+8H+iUS2EPrncfiSobGwSaI898yhaaNB+ENpqOG+a
B2OMCC0cut1vtQnFenTNOi/3X/IMtxwl9cCSq42IkQJ4aH88kaRqBdKM4UHFIjuc
oohQYmbA3xzjYPhRva2gIMVa/PWc+ASqD/ihi0f8H8LyhIfQN2BNEJX0z+v4Owdx
gxxvliKdw31fDo7BpcWKIlO6+KHWh68hXf5wFWSomVt7iDSe6VxTSnf+EnXXk+Ax
t+lsqZKzpGcwHehfZPe8hV0y7xS345plpgDEnSSKfu/JOpBcNRTxgDl2IMmU8SkM
UA6Kd6wubwMnM8zpLErYDCg59gOcx8iwtflI+qQGcqEEnSsizyY4myT5LzLI7O+C
+FJY6K0nVsoVNgCiah8MgFIvxiovfT1feuawKxq9ToJW+hQl6nz6ar0zS777cpwA
gWkHaXgsnqrL+0cwiS4Y+rUZHlrcD7td2/813h8wOdUR6A1TWkUhjVSRauq7qek0
xGuvI7keCOXoHHpwFc372WPbz4QVAQPz4BoZARqDatgHoJgihRWjqKAEOcn6K4WA
iJUBzc6QT5W8AlgXTN3VxU1dsUdqrHXk2oLr8ZQmEml5OsGGrVE5QqvNE/xwZKsK
1TrFluCRGTbdU55gFLWPtYwFlhUI6V9do5PN6mMSG4mvHU0i7bc8ugiZLByE7J8X
O9Bs5ljXXTfO/6IL9kdoL94iRXr3/0tVqCNTj+2JUiCfKrNOsbLX8Gsv6I+MLehr
0kuduONmNSecoz4btAmGZLs5R4WEXYJ8u5OoriydtTCBrDua3TuCqvRECrAzQJR5
RyYQ0Xno91E5h+glDsco6Lq610Hc5U6mQKS+Ihx5/YUYsvJtSJGpod9AZA4U1P5F
FmmfD1usjVFo4B7szcuzXMyjNgH23oM6OVCfyCmkwBHM9rHlZvSIYDU574NF3o4w
fa/71MGs0vH9nL1LGBuLtBY2WGJfsdpm7MhOmpAT4IvnlAIIZkXAnwMZHGQiL3f8
AQNKcxSa0ZHw5jASDbmegR7+z7V+VEhDOGMs0WMZoPtnydfQtkLrvFyBe7L2WFyJ
ECKV+EoO+2HxCVfrF2n0wg/w22USZ8E22dkFDaH5IFwyfrTwXgiDgjeH89bmfcLK
1jRfst/VtwWUqqqAbHqJcU3xIvbZCzJhfBWir0rMcS3sU6o80MrvMUFHy/318a0Q
XtSW4F15eVDeBP/4clEuuPWOFsENnzZNt8qIoACBAdev8nGk/siESP462PBoxMmX
ICRPvBR3zFMYlB1O75N2wi/5xcURxttSXQUCPbMvC+6mx8+nKkiSeXA/dZ3yYrdx
XZUjkOaQPYG5lH4kjntxzamlD4H0H9yAjH1JXj0naJW9z+ppS9sw87j/hJF7JtcW
IWBBZs8Gh6afBe//pn1a2h2Q42Ux0+Va4JfKQcOSmmIReFHPSfp9ehfVzqm2J3Zn
D9K6UawGYIL/LAFSlqp5est2cS4nUK+CHlyYt09HEqplu3FgF+08xbJgFKu+pmKf
mi3/7qEc20ybZ05MZ/zXdQnqlXqVDIK4o5QblxYH/kqHf0BKK7Pe0KsI78U0AC4s
nr2P5VEfFTV7e/t4dsLHfuqpi3tuIAFYMelGObYiWihBzFtCq0AbqPjuKsUvWxR+
lmdKj2VVZ29iNI0ir/PQsgWHFTKyM3aEudi16VFucBowNPS5ke4AOTm1rgeDXi+i
9JkhoWk/bh+sKplgQcYKmwXkdT2KT9tr3quCydLtNfHlH+8Wc2rfn/FcLpzjImTw
Y1y/rBt0d+/D05r0eNF8qY9nH4CcHzJBuDkxdVFG1vrFxD1pVmJwtXvIrR7sJl4a
7sP1h5avo5umghXS30zhDo4byL9ucI2sQo3j2PTGpX2hLuzDuAqL0vDuMvdGo1k6
HAcHbSyCxZe2da1iJoq3DptLmFNP5fCHl87WIZOugp9h/ianWsDX7kmsz7ZQzFHh
V+xumME/cnu4xAwcq8S4bbn1usA0EMW+2+fDLAx6Daxc84KvmGXqly00UWYIqp+i
7AfigQlqERB/PoPlBPBVUnO0ek7bcuQH98vXJDrWONUaaA579gnYnt6YtcSnH1Rm
cPBv8IA/fIARO17lFTfzgUcnHPCy4Lhp2vj4ms+3mzpB8xigySFp//UjwntQDH4m
cZLi3MQ1QrfQYJGz5zIZC04/B1h6ZKLrkO2GZGriubPDYze8mbGycVWTcGNCEWfE
U/ymmQ6pze6axw6svEOKpN1iK+KEOJ1WBJ0LuzhUPPdo8NpnI2TypId8kxbFG555
X2ftQqjLlHxtrPuAYBHbzeEIMwFNNumYXjB7Zc8uBaK+64euwgpH+n3XkUZCgzk6
aDfa6kXvlk/B1JTMxGGDt5EyuyfY9n+IIZ2x6wxx+tSoJeHPp/vj0RwvLGpStTfP
oLWuvnPs+pTJLkLlI+BxINHr8PILyORGwf99s+sy90gm3hv5kB90EtKmfvCvMu7+
sBMWzcLA/geE7LpPNG043nPtki5x/jjJSi9djSPxsTRBo6exVAsBOR55BprvF1il
bwp6MIWDjsgQpj2TK6KXzu99BCjFFbytGcXSG1HZPrWDQPVsttuNj4B5UxHsqoWa
AfMqclEhHPUT+4KY0iU9cfWG5NMY8U7US3xuSblc4VzwwirJ/kXplfj5o4bintN8
Gb3UjRKZtrFg5qk9fmQGlpHAIpjc0pR1ULaIo921JHNqsqC3mstAePM6yI+GY1B6
kmaeUxnCas+xsCGGs65+sIHW1teLLR6GLet3Jb+tnDkKzhGi6BrCqhTLv0mmYZy9
0e9IPa8Kl30ZJVrcn6iVd+qPlHCPQh+GU2YZdTlJZ9kLPan40R4sz+5fmb5ZYgYJ
3Dmn6sK0+lkcCZdDJzmQkdtFdrqRSQuZmprxRwFqp8HzPBH/QT0ysx8Zh6NtPVIp
+1KiUz+AOw7Od7kYHIhcaF4Fyp1pb689ze0AGusuwqEY4abFji+3ui9zKFl3VdB7
sxuuo8MGjIdR5aMl8VjZfXDa+SLfboGnmBA9VRMznzRl099W97ounOeG26INmXb2
JwvNJXsZHyL/Uigvdpigv+1AjqSXkCI7PsA8fI+PqdEap6CoUUE6KbQ7gpnlsA7G
qqrn2HvVbekBLbxfuSmMTcWG2Saa1U1QrT9llj4P1NcyuF45Assr7J0KjK+kuQip
uY/Yp+2CFvIr6YnbJdZYiYPPM/mfnmvF/xosQ+EzQmokRzSBpPMO/6M23YDyQM2a
BjVKjb7OVEWFFsYZTLGb4dYNZ+7s/Kv6RlUk/SusE90gVrPO/2QJcovOq9CL19Oc
0U9BJr8wN/NPE16dFNZlKROEHMP/qKQulmF9/Of5+JdvHo0+l8kJ63wcaOzab8UU
+Zm0xl5VQQdcTrmPbGzeaO5hkcIPpjQEUe0RF4vI+L0hMOzsd4CyWn3+D52Zotd6
PCDjWZrNoin0CtgJNHsLciXeMctI7G7IN8Zel9k7petnGtSnoN8ipSYQhsOCIA8y
f5IqRjMkRhAk4M/05yhxko6U6h1CQSuk1pLdcg06TFrwYA4NgLC5G5zDQUY7Olhv
GfkIlTeAE2oMaZYJfsHkSr9S4M8SVnaxznh4lWBm8Mk1Vd5sRtoajl3vxo231DaY
PDHuSaY7ZKLtdIXLuQyB+H5uNsRutxH2XRbYMFjcKMUoHvTG1nrBV9BoUFBnaNhA
zgNdlQEqcc8ayIYeGDTtAbUjqC/oMZn+mS+LwJVTEP/gWHzvMhs24tVZNu6oxauZ
dNH4NXDfxxdfuPy9T2iqd0YkOgtYcJA7Uw9wyBDuH8hR5j9fG9MNkWLkz/uRy86n
hzcnXP8Et9vrlX93t0oR/UVmLnaIHgY/y/v1laOBr4/uRH3Vy1rgmW5ADS66PZbV
8Np7+kJEC8er4UayZm9U+CFnhfIbw1ntlZuk29l5s5rLjv+5DOA/BARknuqPUXGj
pu0+ZLQIsAM4V+/kb4RdwABQxacnT5pl0DYHhIqOzcj3ZC3EJhXs01nQrmVmL2Y2
5Kov1BZ3JuxYuc81FWP8KiQ2e5AWwZkFr0glQG4bx//rtt3mrXdt7LHdPNxb9UDB
cKz+T9yx5IKIsX/hmqEanEbvkAEXo/tijwwu2T+Mn66Rx0v+Hu96nctm0pWIsXat
dmZk/oFkIIm3kMQ9UVugwb//krwS+upoycWHr/hY8iQp7dMLhDuG3mhkGwO/j5Hz
bB4FAnrppfoFoDwtpVaelqBSH6jsBJT4uYaZ2oWPELYgJQ1eIJw4e3++4KzxfdaL
O12diGCO8ecG0/dw66fCmJbiZlITMOys2mlnFwAZGwAgzm6lyKnyMpLyppHJ+Ha3
ZORU432nyKJSb4awVmmsKcZINZ3L3nHGs1N8FRSK94RadmR2+MczWCEod2zJquuh
xFm6x3jGN4gq9L8biLtdFKAhViN7kYTw7pHsGOXSzV6oBcEz8IloZJZn21aPUzmP
RquEWfgAynrCVUA+JgAP0oN79xM9I+SjfXZJkWbGFu9k1F8kY9lDgyt7dV4b/zlD
7XqRAON2EBJjph06UKK5wC1dqDKDRJBphM+FJ366A8QKMTyz39C3a7YGXOI6+9Pp
PkK2aF67/rk0A+G/mKPHTRZmei9bGCncBK3DoTpXaFwmv5cRPB8z/ehe4H8kk9j1
Ez2NmIFn4PeZ+Q5DEzH+CtdTmdPUhLlquLkVQOYsTx3ETdZgC/vAPp7FJMV6S4FV
dNTEUGHSf+ON23Zlt1KJ0Ri4FQzwO5xWNv6iw1H+pkly1HcZwU/9IuV4Dezp5cDg
atxscNUEzSIvvSM3WG9d2q4RKIMiC2kkIS3gbBec3UEVV6vXbvI3EttlM9Gn4idp
0WqGZstBhFXY+RXn5B7XM6tKpJHJkn0aIljVJwb2jR7cJQuikyfvi46hITix2tik
szuDaykrAbRpvIangh5k8XuJPTb/vl7EeUEsUgFjQPpnNPgo2w/bSCU8QF5egiKZ
vJf9QWgVDDs82OEQM1dQjCXYAXUoP9KypnqtcJX8l9xHTAK7IVmTU+LEkFOaHAzy
vowRY470yqomy2J0unzubs/aGfeSVOUo/VXbtWYhxWXB9TWifuA9XuKDAD6tVpUM
JFZ9u9jh9JYjRsHISoUVQ9zn3yEHaS1fiUassXWEYQx2KNwQUcyXMXwnomGqr0nQ
70pUuAWEuvx7Z6bjensWX6nEV4Nc1ephXHNXGn2qusTcvtERE1TUD2VnrkIThbrO
6/Ijv4D0Eb+h0Bflw+pTVD1kSSAocw7kw3CyaIfRWGCsbd0h8HxCnx8v3EpcJLoh
7xVnUEdpYFGoA54LKrUi1liWqAEaPXuQvU4UjpGvn5bVvm68S21N/Ovlm4R+i1Yi
uk/x2LxzOYCk7bkcz8bYfZXAaT2Di3HfxeXIrzHpG+oxkWjVbpR6o+rz+4LAoG2h
OnkKvzNp1Dp/35wYMm9H/mmt6ppkDACG7td6zKOUsZkXCmVrB1jakzjTPzell9zF
Vdl668med81RR6DaEGuYJU4rpNkObd30QYavOtk1zLi1G6z6BxPdHgrl/XY2Lt0c
gijdlmL+h+va7R1f+Van/4j6kA8zmk/gD7e9TN/EDP6jYGLiJ+Wr6r2J04BzpoBi
2nLYjPDrlVrtZtpYOMqxE2u2ci+ueD9Po1UCYu06JkOHVBT75ja5sy2EgITUiCA/
eVqffKhIgqO1cZ+6nCFikebs9XpcF/XGgseOQPhpmJtanWXzCBGd6bW04NZofZw3
h0uxOeQU5zVL6C52DLoFS04pTxpZ9gHMR3D2MNVzYXnLH8b+NP++CG7veVQaUgcD
Y/Pt6DM0dLFA/m/hZd4y+uICwgGRECmtKqE4ljToa+DE4sKOnfRfEED7aRL9z+xa
XF/NOuuUNpblK6J5U9mZmRQBc3HeOtfei90KJ6GcmqfS+h4cPcDPVWx6WQC7S1w/
4tCK8H/2qCZZtgSOubA+ucZ8SZ8Y6TL8pPQeIbg8tB23BdZwA438tOpCtdnEptp3
bhe9ZZk4+7qZ0Gkf7zWqGuo+PVUm/WTw+r5U84P9n4xMuzhDiGaDhjuua4G3D3iQ
NUKLl6IWycz/KL1rvVeN01CJmOnQoD+Mi9kbg3NWs/D5nD89RsgTYaaiGcYa4xMP
4ZZKxLF8xFXZge0GxoNNdz1L8zE4O6CwoN1HbDo7ta7Bi9NNc8Cb8ld3+PPentsU
B2zdfKRWtRi0Da5T/Wx5MSpmRg5g7RJ8zvKwk+Iv0cwrivTiQqkM3YdyF137RgJw
XgzKCdCZcAlDRTtzE0/aNCrAoyPfPTEpFOSVisYDrOp/vJ1Cpu3VlciGJeKtYBCU
Jfr8RIY6saKn1Nm1/nO5KXavFpUrRepHlu+8oIMjgum3F7+AOZkr8qYYB4farMv6
n7HAF5qu3NamlTY6deoN9K8hhEydPFBDkRRNV/xIzAGldBDhsuCqkkjiBSmIdbmw
L2z6hc7ENSvpeSNQLnC4ebwoRSnETEQoK8mE/KE/SXOWG76KXAeYLe8jWDhUcpkG
UI7dVExAiAqqnDRRg7PHPV8G3OQx6WBulrehzlgUQK330kAsEuVtRns+RYL4z+Ul
Uwbuiw5xLpDLPBZeVCxORPnuQHBOe2D8M9hQQkXZitlrOtq1Nbv/z1xBR7ca4VMr
McgZi1ISfh/hSL6yI4eKSOrUhm1+TSkV62q5NGmUNxVtl0SQLyJWYYhwYGbQufd4
uNYJEdTP5oHZUSiNWo/yZSwBBTeNRfAHc7YmoJR4UgiTma3QNK+Fmm2MdhHHwKNC
jaCwem+hqhJ3Td8OCe3EwKKGl0/Bdn2bOZW8TYzABWlDoLNHES8J2D3srxAJrduy
Nmll3C3B8WJeyyso/twoFJuvVtsWWC4DvOL0imiDMUDenqQ76w8CMXUGqczlccFm
AsDi42/qJihzlnp208BT4yE6wyh0xIDcJWv3DWWQImowbqWuUzen2N4IBfkCzRC/
/Dx6QF8a+mGKX4t9fXr9DAWoVDf/bQSWsfxqN+twOEa7+N+iyTwH8Fob9rBOUcBG
Jm9j044BkLkB8UW9UeSEMjQVAiPSEucQeDBOFD0JWLd+cng8P13E6AmN+tPSsUtZ
2VgejUtEScUefCjwvWpvJAfpii77U84SMHZR+mDrLbrbLhohLSPrqXocSqhW+2js
PbkGeP/7uVRLTpcfbnNNm9Mrt2QA6fwwqwYHNB90oIjNRwLn7LNg8DtRxopcBPKI
gx9kZ67PSndvF4Xh4rCMS0UWExBMHmeLmnUn/tnCmGe8Ysf+F5DrWaOhk7kXQSrx
J1mf7A6s6QH8sZCoiOdceVQl/bP94ptbAEC5K/HWr4LN1FtudXnFRpCcibMVLrca
hkVg+lh8eTgQjxeK6PP1KAOWTgHFqI7gZxw2y3CXxhyPGZR3VHm4exdzYHJEGqq4
BM++SIUXazt/b8knxyUTH5A3qj+OS8SFfg665Dnrmlrc0xjEUbba+zDkJAmxinIr
E2YqVe1tB+HxvGrx7xI2MGYVO9dysJ8zbDtaArORqz4TV8eO8xIINvyBSMGTAgUb
84wrNE+hUJk4zdK65g5hPJSg5UXclEqBAFlJ/OXeD1fc4RYWAVLjAp3qBBczahRy
IlPM0sxyH45pAavnYWNRTeHFJM6titQTaUIvzampQjGSaOg68mKrfO5kS+KbGYt5
PIq9sznppGIsOPdr0h1NyayY3X9MBnOXKWpCGgRLY+eFJz4SZcKq3w8D2V4vj8Lm
EDUDCJbTQxOOkjkHZtt6zFOtKVTnAlXBJPaTgzNXRCkz8o6nblzg8/GKhFE2Yyru
YyJvpj4KcK6AJVCQzTbW2aqc/SlZ1UYP0xd3pje6fTZ74QxOxC1HjtyJRXnrxSxP
qBD96SFEj1rKBAQZ+is6v5sj4K5YMVCUB61tBpZiFJ/ToGMd/iNAiIBw0dp6tjUY
NZj6JxnshzD3vmCyW2v4K0UuMnjNOTg70tRlWZ6hqJJUq3lrdCUTXysbJar9iAHO
2qwSSp9wLzyL3cHV/0gNw6OImqLmNAI7qQrg0Mh9nEA0Rl5JjyRueQrAi/C2Fd8x
Go6/Hbi4YGaSj7HDD8LNyVYJS4dcVf7Bl+mLvZ103AbJic89xjJJcDUwwk8Bfisj
Z8xu5QX0SdhaSlbpAcAYz8UOgw96okL6cHH/bV+8hQBeMz1pvKdHCtvVhvFM0PEv
U3Y6eY9OIB+IwFhYXMpMFlMwx9Xjs+Inz2SB8Efw7aUdVX8yBTeTfoYPS1Y4fPat
JMd7S5S0T/OzUl9+Pbfwzzq5oZhK54ma6LVJDsY/os5TbDTYLiWIm/7H0gahcW3o
AAlpj0K6EexQpX1oDTYpCAmtFsKcLzbZ/m/93wH8U8cNF/6uIw2kEJu5K+3qnZGs
6ul5qhJUcgDFVqmfFzJFZrfaY4osDB75F7GMbNGbKAybm2NBhQDPFgmopnnjnJyG
RpzMxn0cUvKJY3VeXLl1hNzZdKDtru79sXO+NBRX2efODvTnV229SxKUY10J57Xn
jFwP73LueCUlJ7XZMy17ELOd5b2aI/zEHdGOqJmvSiaizWiLbto/Fmox5x2ECvA8
u/HlfUfzPwEeVrntw1SRAtFtJ68XZH4iPBUtxBgrJDf79AuVlCbNg11dcYhFCeY3
WTpi5EibX4I1Mu2Mad/oGwVvYWDBk4WTVSTlPjN6EOPsBRj49u29laXuAY8IfKMY
x2hQDtxb5dySj/Ua5+SI/es+BUDZr0/3QsnCJivJTiiySPf1PI4O7KRPtNb0TwGS
rP07cDQV+/FjEXb0HhFuXRS68+TjzapzLW184rHxus6UfgIoPL8TzNBnYqZk5fvd
1QrNTkC4Pj6yIsXW4UfBe5VvM7XjKM7YgQGtM6KyCz2T9QKaDF9/IL933IuyJhkL
JdafMUPq6BRGnvp58IUx6uuO+w0pnXsR23lgUfOlK1LoM6S1zx2nyE2VW+a2yg6W
oaJDaqmD3ZTZcw5WEEkCq3byFOK1nxIXIa2m1OgHeEUE37KenMC8mp1rmwEHGOLA
S9QBVb7PV1azjvixBPnnk/RNjWVzBVwZEvoBG5HAzqDBVyOtfP5rvnvO6R/siBDk
McgdV+ol/1hMEcv0hNMV7zzzoA4wCTtmDUCmkH8VT1qNx2r1QZjucsGFXGODab2g
F1ikLOqvLqjUbb4Z1sLcDnc8Nx1MeTDPoEDIVVXd74I0hV50qXBlv8XEOy38CSg4
rei0DmaPPSryk0WRVDphXC3ibnJfpF4FBN9CYAu9fI+nEc6RnAGVpZ41HON5UQ4r
hNgBX9niBuUxMlRy+fMBMd44Bd/dkGyk9wVosCqEnjs5WovrvZI1jeIuMobF+81A
kVDfFlauL/vqxpI9QTZ3wLTigTd/5UawlzinfOizOSDV+pHEF5JGn4v2Duj0SNa3
yu5BoJknFG4RDemGsoADqz/NdzWov36tcAA1WbXx3PKKWUW9/NlJR8X6WA03fbst
40QYKZQImMWl0pH3u9c/24uaCzMaDOg4sWvzq7ux5vLePrxmGw6UAStm7a6RvMZJ
1+wGFu8J4kRR+WZD9kLkXEsiw9QdSNbADbe6D5htI1cEHYtsKI+c+c5G7UJItDdc
u3Zckl3elQ4ijCjhEy6G8+aNqSn0DbbNCnkCB6rHJspXHxZQxYqizkRHXwROBY7k
S97/snLOu9lemVZovyJ9OJn8btl9uHXQ1ls5VF+gNynkZhF5/RMDFPzw+uMc58ti
mPzHz2ajeLH5kPcl0ZpieR9bnKcxkWblNcLSMvBFJWJcdE8ZLl8VupkiwkzE2WQ7
QAUVsOo79LR8/rCpisofsJmdcfpnnIoOLx7geExfM/GI0MaZrF4jKgAYxXiAu+DJ
zupr/vgj4cKZkKgO0dQuVO8zpddtzbE3zxXKX5c5+NtvSf0krOiGyH2n6IJb0Wrt
sHe8u9wGNmOFyrDshDQAQShBJ1If6koFcZawGAnywjhLkXiWXK0Mk4PiuL4haDLX
jg0p/bBCAtrMNXKr82TYLZG+RtsIvcLS87jcTQe8ECLpm9GxT5fTGyzV1CTDsQ+q
XZZ2WR1zVBwchFc97BM7z14eHuQYwm4EGpqMXTHDtHfJ7Um2HWdkItGGepfm5irD
L1V6ifRz85dicw8qrI2mhfvDJDTdNBsckDWisbk1Qz63icvpDyac+CNDuGs5Ua2y
3s87vz7jUJrbgC0BBhMjypWeqat3UVyz7YVcBQWLj4sPDnp+VIn0EehU+8DBzJrZ
874b7IWlCCQJyd8T2rsW2oPTnxQwj8NfV9A2Y7FXucPfC2BOXvbCd+5dFKuLW00O
myGxbh5r8XHVJUVooQ3xAiMmfHvgmOgU+hYP/+pN4c9Ar2nz7A8alHsuvEyVSj46
ijZWzBWLBIFQhTBAt5AosdZXiX+MJuoTB8BUbNSTMASdKMhsK3pbwmyKJM/ipPVt
SHb1KJVze1Aa4OGLNqDnkok05LVENU8gLaN1KjQrnfvyLTlYqTj4mBW2Tx2KaFTo
cyojH88Ck0ujMhhl9slyGPIwcO/cmBQkeo2JcNdKH++l2jHbsAOiOGnP4YZ9gQS5
oLiMhl4ZqLMQX+ciwYctAdzD0WACfQNodzwoGkkMPETlFNJP4EzDm3ArosGFp1Kq
VKQiqWecn10z07eubHfJnYGXu0Y26wts0p9FpK4UaNq9++UV+1L3hHTIlHS5g9E2
Ob4bcASb8m01/8jbl/Ppbmwu7U+uaYW9XMyFHb9//4ZmlxmXOCTDAZj/PuAktleH
Yu4Le73GVEvIGGLdOMDZr6AieBgPmuRcISoqlq4ctE1ylqOHqNq4TAo2e/DWOBRO
yf9DQN8Mh4xKgEbLaCismaMNU78n8a74NW6DXOOIM9DmMdnWiG61rxBgDv0ARTFh
WdoJkp0rAEVyyI163AlBzlaKSlI+/vWIcrfjiJIhHYYDJ+YJe6AiLdpkFalXtxOp
lpqDBQZ3c3x8LQRTK6BsTOHfsZgqpWwcyvz5ZQkqoaBrzlGPQNYrOkoILE+sx7li
O8zz7ymtY+tsoMPC5zVSVLl6HkblRDASOzdWU3Nk48FVi/RWAXp47C3s/G702ljm
R3iJoVbsfMR5LoF0HAFjghhsvoNj9t8gYyuY/BviZp082sml9HBaWcQ7kEvSYE6O
BpKujsIXe3PQHNGxco+TOlSH+6Rkvtm74Vkpf2wB7wJ0HGlsdwFPBRkgnK9SVv7I
Ngf92kDVuQAFDUY9TREe2YX1N8KeGEEj/lR4TUamXw8zV4qwGkHczN+tbkxXAVfn
i8XxYbzE8VOGjnOeRDR4CjGkPONxj0ZCX54S+/aLTit4YEf5hzjS3qmU5Cq9Z2uY
+GEyyiWftgJjIJIJC2qdzouIXqRHjINiOyD+2ye/Sg3soMUjjfO1rj/2NBCWO/E2
ZDfRzhDr+HovRlzmjIv5pPbeU0G63A1jYyHIFiBEfqXLaiLWOQx/7PuXjx4OyIPb
Vfcn2axd/KovWStmx6qn+oxGHvLWTAX8ogObh70VYnkNuVz1XbTp0g2fUalliXIn
V5BSj2QY1O3vtyOdKFOF6N7QMbsNq7Bd9AJWNYzEPDIlb1WW/zuhHTiLY4dJrGti
8/Ru/G0hvaGI6KSH/3+K8VHc2WTk1LsIaECeAHAm7YEG3Q0Sg8EZ3HUYozgVJOx+
hERE5J64yzsu7TFyV9irayVA0ColN27DecpbK54SoTqB2ZM//CnIWxmDXpTmawh2
vloUYAO+8YWjjacKYk6yEf3a/i5LfUJADDwWBwyhomPF+6ipWmdVlxfEwbGf5axS
VO1QlID285BlJr79+IiMmmWdUqX8U4bdzioHa2Vivt+QUbMjTXaQA18rAexsaFLF
2NtCdIL8w8rhkbShqfbZTYWzeXbiAkij0QhH5FOzP6uHfH7/l57t+oA99Dbafiji
DUm7Wmbbyz4OwVeuWfCceROlZFVLkA+I/hXE2DRhv3Rvw27n7mrEHe7m3SR4+tu8
kl57yYBnko97FO/1g9d5ulBnorukBOwaxR5T4D+swZv8Os5rve6cnoTxw+Q9yo56
kyoN7AE5zp6ixLnZ+crCzL+1of+B+6tyIWE9KgD74hzRv7tDfHBD+iDPgdJq5NuA
GZ4lIJ/o3XyRuXPeO6mxSVIiFk3PtB2Jzr4h9uMN5WmPyNht9a5niP3YsPSQh5Le
VJ01wZ17cSm3RexcZwuHXvYEhDAKEaBwHuwByQgFTTbJJ5qFvaZ8imZNSfzgqk3l
3CjACeLkqYoLFvIxvYndz88abAe7BIEltIaTyQMC2FxT5/0mrxGIeyekPuKQmX5s
XdzxszRVtjrKLwEHXzTfm9Q7ieILwSOa/1FXYLJ/t7yrMMaxARN39NNM3tHYWm+t
NnpR6rywT0auRRP/g2w+WhZEv1v9X+xexiCJPbLwZa4mNFyOa2sjtFCHLnlNSh1F
HZdTbsZ8+PRvBGbBzfxnxs9B71WHPmOLVklIaeBeukX7qFa1Olt/BPDdNB8VqnLe
6hqcZ7P+VSLXf4TbjGJUKfVHtQiNdPwt+N3fiFx8VJv8asEm5USWsv/D30wExgxq
w/vfL6+SXKoK8OOKq73z2PP6kjrr+QE+NBPemUH7nMa8GMPbKf59XEtEsbSemf+Q
004QKhB7njsP35DSBB+x4w9WF2uhrsVayDt1er1jh5VCdA9gk2IPAmztPqryhi+F
LME6/tJhIWGVy4V5XrnPDdlZxv13nXwQ8SdoH2vEfeoApWiDWbYLuzJmB8dnwUkV
wMSWGQPWlKdOVsRH8WYQ1k2GLBTKkIkVhr7OlMa9t3JofDu4ovqCphbT1LeCCo7H
tSgtmpp8V7McUMKrSYk6ck8t4Go65p9jSGNYH/RvUVwO2gIbWqcWZ/7Get+cN9KN
F6Fps8K7npkiu+7MuhFr93HzySOX1Xod9+oAYI2S1yq+IV9BmQmfY419q5cdeLAz
ovJL65CiLXk9uFAF46QgP5gUQqi/crjTARwxOrD0k76puwNGuKkKmJc38Mydg4dE
sAy+wTuxNfNro1s5KeEv6LwElhQ1vDUh3AgmgSjMFXGcAKJqcixiG2ZcvR21Aqxg
St2CAmKP/8OLpHJSPhiDj2tQyC8Gu7swtlU+iJXxExkiM2Ue+qDTHhmgGs/6jE0w
3bQP1nfuHKC+zfX7uDqFGoGbS6hP9k1lVGTbLUPeR0FTxUf5aDSJs5qb+n/vM6cr
qdm29LT9KEqhOtjUncA7r+tTRoyfz2cm81FSP4VBYayjC4OjPczPo2N5zS04xkYH
GwBmREyLT8paliLaIOM2SQmZiKx9usKCbIUC8meSgwuJoFtkmp/ChrR+mnz0135R
YsvxDxI8qP8+sDvxIIve8ZfX7yMMZYBwYc9oqdjG3OSnPm+3v8NBxylhGVq6S9Kl
ZoF+P887GKcqvpw9isTzorkAce2rHJs3NgfymvEXqPVisU0fsB63C7ssAZQfjdSN
uzQuAApk22HPA5lLOa3oGPMuRK1LKHkiAZgs7+IS8j8VepIRRVnFjrLO8WhfTikL
Np4JV/djih8cHdka40iJHXDgaglveyn0aRnyft49aHJSxlyrtq5t6J7pa97ObTJd
yID9j3oTr0DUdsM77msaeeTQpJ7s+wFxI9xypYwBhcp1dmbOsTDpbO90lHBjQspy
0Hn0mlcOjtFyfY0MImS65O3y2c3DV9KR/AIAieUbNyOdXzPxO+OjelZRpnNCrtmB
kOtzteEbKTZODIy1VQQ3hTAnTNLfUqtjxUWdcYgpiuxlkjfGAGsNigOIWsGoYXjR
4md6/1g3kHVHWEgV9K2uatONVUQfBRT+oLSwprzvsqw27Oo+/qBvDu65tyetkTmU
T1BGpfDKzgnOGnU9V+vmB31q1/bm7gt7uMi7p3YRlnPVX48aG8qV18BxZ0vrQDOk
eg0MGMbB2wpBnOkaNpUd+QgSszq3pbY7Cwsfb+bSUi2//NPqInDQcAH1JWTXvvdv
v7I95QSwNuOhZWzFKGKPtxtxnaFl2Am6tGAjTshMXGmDq9z66nayrBQ/0G6phatL
DqVxzL2Yqbl8mDJM3LjqnGyiLATcDuCEtGuYWcXX6fHyoI5XgyhjvU7ypGl4UBvr
C9100Mx7Dtnge8HavfMAeAmAm5ThXyd0ThcgOgvTZaaYgIpErF83erEgzcttmkbf
c95ASrtSOdHADBBos2uX5pHj+McJZHg77D3IrB3W9r9lF5Muz3FxbpkN8mHTDUAX
/mtC8g72avyU0fzPas0zOJt/QVccI9lW1hOdtXGo6Q2+YtRHjGZ4RDWBe1zNH8NQ
RKV0GxwJ3QAU9FniZYsYtgtLn1viohDlz0nmiOptAorf1outzWpkUJgrRxTfeSbR
Yn2vI/4WPLbaM2Dir3dw2Oa/7aCsfsvCSknLYVovjQPqYDD4jQOJNkxEa1ICLKlT
PX7oVubEL1frNdFXroFmGU189Uy4vPw6kyGWJEcn1E5zMMea7YE/vyYAbMTqoPfu
2MrDkiLm9CKFEThYOTedAAgHfAf5VIs/5b+Hcdy+cRB2Gdx0vQw7wKVV7FDjJJ02
/MHBOm7kGF7nxbuHdy5QApSHrEJKL2TJ0gIA7/0/byyLpVBHZBHuU3+idQj4t/Z7
dUTRsfj+Zb64SAJNa7ABaXofp3RSysVV29oEFwIGWj5AeJyLtzmS0yiBzrgnbGt2
e1HtsLrVm/kPiB8il+HA7r/Q7INApbFi1UEAlPWn86n9HQqIGufUfmyyMJR4ymv2
HQSs2/0yxz9ZZglNs5nYUsz1f3ofcltg0WlFX9JvDaevxM4lENZBWF0J2pBOv2FB
mpykZFdC81AxbAC5fwQF6IdXEj1hXQPY3eXCuzVBGkNuHTSsn7lzSwvFnkBRP3fs
MVv24eYz3lBxSA1rqfcNu0dreqfrCahS4L8G56imF4gR8H+WyHkBaXRL7hOlqZEX
IPsnjiHh2W4RcoPvC04KAcH1LKKcokHklYbWNmtZ1HnFdGwzbn7xJzh/puUGno/A
cBNB3jP92xVxmzWprDbn4zXa/WlZ8PB2pV9mFokof3K5MAaOr1MHickfoaMzqQlk
GrHUCTR5ln1pmZrMeM1xS1vY/Igt//ZuvUoPdcEBkq4tr8j6T8khdGbcw2U2REGF
xMpXjJWB7aJY5mhE8Jj/7ekQK7tL78yIqw3+JM2kT+kwNt8MWwaH2Nu2y9jhG08b
w0gRT7bGzbKuzmcfy/gjpqJwbUgKX+5xWu5NeLAGEiQCFlshqzlc+pcqXquCutjH
xz6AB6AJlsogxwiTNWzhga0aF58U4jDOliVOF6/McWg0zR55zBHai7TZvIJiSC6n
L+uauXO1NxsNgaLHcapHJItI2OJkPMZkgTqy1cXlBOxQs0+8qB9T7iiTufGD6X1P
TgrNgllDuxTAU/UsIBu5wHuJqzBpkrx+vU/DCdTgwGhXNgrhxP5BCKgUU4l5Hb6Q
eroqHLQAyvbH4Mf09W7Vf8eXGRACtrl8hIrf5pcLcd2bHPOVQ+PeDensR46auILt
BIjhf/cWRE8hSBpmefoHjhk/2BDiy3raBwKq1fYCNqkItcUBRUbnXY0WmHUM65/W
5SnKZKCq1dvUR/dpFzSPLcNPkVOa8KnSi9G3zWErWo/AV9348tKYxSS+pfnj7S/r
yj9URg3gxxtjO6tUJ909x6X4x0i6pXrFYxG2gMjmLQlvdtQni/zGEVWCnJNHNKlx
7Fx6eURSvRdD5YaRkoDuU/ANHp4QRrS0PvskkBIuajeREfUKas9iYcpn8FSwPGUZ
b6XNL0usiDiHuUlrrgmWNoo2sTdYCl5mNnyQQpZVWPeRjiCybRASP917ao3oYe/8
oG9PzSDFvq8hudeAmT/0oZVnTrxN7bmCmg0qh/i3nIAC+GNb2B43wxQ2Ux9Zb8pg
axcNyrA4a/jsrWusZ8uKb0Vck/PqBHizt574AeURcHNWpHCthuiIAo0gP1XNx2uL
7Eb4E1Jkdk3tP713OhAyVAQqVaorvCWXkMOfrkeV3eyusfweh3PBAb9IW2g266c3
EBhqrUaRGeniROWwqWCu0LiJ8yNCG564VjL9CG+dKG5RnQAE/9bw2uDmGQbOIDwl
z09n0h+hFe2kPoSPkKUQlkA/0fzO691h/SPnh9MZnaweDCpWlkx85YwoLRVCG3Tw
k/KQ7GnSII2ewt1v2wNRlqb+yCrsi+QoENUT1+SahPPEz7pJHCjS8e1KsTtvJCJE
0A+WESlSl0xYWLgcNj79Z3RX4pVe/vyagAKvzbzbkUhuP6ChI22Gmz0EBEVv0IsM
50H9UJdSD8wTwV4r9opqzcUpK+NiudSDYxxNfdXcZFfhmpV5QLuKqi8PieAVG0hf
JxtyXLZ1EI9KJgilIMyTWI0wDS1MX0ADEkC4oauvNzK4INQB7Hzck+6DG6He1MEP
5pSBJ6hKohvTRax8g0wgv5LAjZZW/PMF/o/jUAsRtsd7bN+A6dXsoj0Gt5UjTNJl
BZmquQM+qlSDhYVuqoB2Dlx0UFzuA4ktz+Jh5pRC+7uy1/TASVMD2kkFxD1jBFIF
c+02py0fvTlW0RNYls5/mRF1p+Vu2LVAdMtKTrqbt7Bszp9kXb0AX07k9LojN1N5
+muscr1d87PLXLKs4WdZc8tBTT+8mW1+cN0JFJsYnWQHeDJqOGwpGmXewLogLh0z
VmHdM8GPGXvFmkbBrSvvcX0RlMIQ04KuIfH3XP6916cRGSRW0fVc4hbHE0Xg53O5
jGyNyN7U1pkonzd/QsPoOviY+u1/wItEpa/wtMbTSQFZ5mDAHWaeW3s+oRkSVjzL
OyODQbDgiI3ndbJ7CqebA0HAVkACLLLw9qUKpm/ccL4qxaN/uOprvJUk86imMKV4
nMsjlXM2+s5m2WgTpR4ZHosUtnlISukO68wEPHg4PCXeS84gOw9/DweI+HPd+FcB
a4xHdp0p2XzZv1jETI0yuts2ufWuGMLHRZ2KK0NyXYpWU1upYqu52YJg+0PXYP+M
UMeN8MD3AVid1Oj7AfvLzUEOT6rCVi9ZA0R/cO6uc6h2TxWGd2OtB8q5tY2wjJis
WGuLdVFaEB4Zz08bf9NUNWTMldpixK4qy1TCRo+gDZeShzhjsaFTlAY+gqFk1bYx
7UGinS6l9bkvZP7x7ruFdzwOeLoAWIVaaMsb905lzZJ7iwtvso1FT0JOpTLaT7S/
JnmSmHyawVfiIosTDUv8DLd7UqFfk5AIrPZPNi+c2x7e7m7MEZUgoHI6torRt5In
3vWqoOJLnnIL3t0fsFkNa9DvE6/nOL3Yc9EEi+2/BawGiF1pFolMVi/A1bNwp9lh
kaRY6wQzFAkNqUdAJEC1YDcYnmPvU4MPF/+BvEPmsyQz9GcM9Kg5m6Xt7DKu176p
fNWKT6zbCJyvUSgkA40H28KZv61j6egM9atvW5VK11KTtEfPAevBxZJqVYoQanZs
17MJobKbORD1OINkspxjpkXnEPy1fLsL9pajUtStpZ+0Ht2ob3u4y4hscLjOVbF6
5It7xh1jFff20Zva/I/YZQrax/vNF7DOfwXBR6D/W/MKJcH0Dn8jQcpopnM8DRgI
xRTgEsCJaRIax0gkLdzKpl4sW8yJ9inNf5g1szJqpbnZ16du1Nx9VVVDZPaPgBgr
6JEWVxeTMLGzUgSZMAlK/zFcpuaU217BuwptyvpIsRXdhERffCIE7imVgcV9FUiX
mpRlqLwixzX3zvHnSKhJPCqHWfanazTEqGWgppGu6+vlmhOUkxBFCKAw1j9yiMz9
uSArybHZVDQZHu3MTZothR4ZYvyPHSOGXTqxornNQwWekY08LuTvpFAa4VdhstK2
1/lMS73k3gUsucZ4EiT2q8S5b3Z2Rk1siLaBQf/EfSaFby7Qc85vn4Z2p7bwH7Mj
EUuYXkpmGO/niVzbBdAOXBGFgYjo/6BOXN4X9sONHTJC33gB5I6Ymml5kB9f5+KN
OeXkqB+sCf+Yun5ZOCuue+EDjtpE53M0AaMdOiDUBa5+RzDcje3xRTr/kaUOE+9G
POqt5kl+oJOc2gq0Opt5JYadSoVWV2hVxLAXMkchiTXPGeKVFhmyi017+lb5729Y
expsJknZhuuChW+xfhWyxC9Pdeh14Mke8NUxKa20CT7UZsbfMzr/jjr+8+6S+rTz
QCXbxRBtGmtT0Taola6RELlmEzqXva/TTAyurHYzUKI744CgNNKyHGPYyumfKauq
AqrKihmX6r0RAzhWaf0F2w7EWAYt+oXCGL6c5oJy1frEeqNrE7yVOyBV2MxHlWj7
DetKS/wZGt7m9SyoMFxjFSxDqSsksDDMWEuScXJY6tjbCM44CLszvwxjl2Sbmzvj
2v6dqb0X1J5HKLvLVs356hcGV+PKHxG42fD10PDZK2d3XhIo0bDda3u+E6QkiEpA
0KHmW0o9y3ZqjCc2VUk1iVA3rodlaAfUNhX+Nk2kQ+OkO+Wx13dPcj17QwccJF+M
NGrAqYHWBniso7EfdqhN2QvEumFr8uOeDxV3S6KLotuP/KgtgwosCIKjExD8OPa6
P4sdZg++Gl5imLLbTzcRTtUZs5BzYDyQ3dlXdF9CkB2aZiH8OGPMW0ZH6UV2pquy
lclU06FgnobZ8pN0/SQGXqkxpCUoZ6BRaJoSQmYknvmkES/YDDJl/7qo4txL40xx
DqktRkGqYrayjp7tSh9vLeTv0IOUMm5mw+gFEZKJzK5q5uEx2ioRolYCy41B3RNn
Bz25PiciW04D9k4mdGiaAbzm72bFX9e1Scn2PUgMoamV6IJcoLjCDXLiscBHlpi2
8iOhfBfNl0n70TXlsuC5GxngcXEjMGc8B25U3YqWgwlrc/SDFaPVIJ1WGJrumNrv
Sx629fh8P9OQW9cpyjfJ6oa0zKmmmsvVL8SNKT2UgW0L8RMFFD53gp2tXupDTBLs
9C5n3+iw4nCeyJ0/z/9Q71CfIEmv+WhM3/3a/0t/51a6mTrxbCdvIWQbkpXsYvS3
+wbq7di456MSeNRe4fffEnAPkvnVOtQi0XOts7WDWwrFu+XX1JNws2LzdWyjpAqG
Ku1eRJP5Yth6XwjiyVb4kCdHDURBqy6dbBvX/5OB2DFzVV9hI0ZvX5FYnyZmyljR
deIDXn0UtFxBx0V65C/Gc6X1aWLlPr+jRJHjPuN62rTm0gA8idvt0zk4f0FpAzyW
6gtgpJ6GpEEV3cXSM7PHhfZU/T0uwOJeryDdSP8e0dxVOpQw6TPNoyVTlgwgbTLL
+1Ez044SglGHZmxjSgVH/1ykxt1nGsZ4Jbii9206bNjOrGSKmYbwmAHTIMw9gcIi
1CGk6HvNiOhpYhqKDn0TfPKBhFTgkzA98pxxQsorhq9z9Rv3I9QZzt6RoXKVEJH+
Dn/vpuqyMBCf+lXxgX4Y1XweszEBGYy9VgixIjV0l4KYnRT5fJ28xy+bbClce0iS
kuoqEjCtibKpxVA1j0+kwQZpqczzhh47J/l/iuy4UNsOjBslBSbAC8lFRaKykae0
24ndEV5zqluhKbVqL3ZhSApNx7Vgl1Q78v6TqIu71aWPSda4MXfZbVkAtwNMJYXP
QWlwifjvBg1gbsjo2zKktANE4KG1lhiXGXiT1GZ2LG8A82F5eInpkdxBxjDoTUAO
0s/WrGdYvnPDZVjiK2H3kUG2RbUL5b48ZGWpamB2otgQ1vJbyjnJl/gDLT7AQZSM
b3lC/4FTquY/gF7bNtR1FE3sUP0o50usvcly0sx3G2cdrKO13cKDfqNdF4RIZAhd
OiEVY8n8R570vWCgLRHFbQ4gIzMAHPDMc90xcNM9p7FfW5F7CykCmLaIcJP5kSl2
pD+2E5OR4F4bCTNOtRdZCeDR2N4lgiFcFySmtU10SLxgD5DvUTKEPrXTRheVkkL9
3reIA9Hq7FMl7lbcZVESsz0U57C4RcCFx6P3Nfq9AjcIU+iiKpuvKBIuHVA2NBkO
LBktqVjdTGvXXJlauWr3i0x63DZmjGEoBNyHc3Sz2Gkr+5YL6bh4jTRYHsMDYCIA
akA5qoWKzCtrJ5w5Yc+TVXzWcgpIFCGC6zAiFWJM2+b0vymeUtFW86NF9oSifnmA
oUxk+E2zNwBD0WCC8Hxg/4o6l+8tQ5pv2W/rjn7GAXyrAg42k4Gf/AWpRVED2SC9
W0fJb3wBFzoYTiaJQ8BqastFkpOOjXSPcjt0Vec4sFZxpPBvyadEUYGyA+dGgERn
hIWtGkFllgu6ASGl8v5r2D+wE0R0WuR3hj21ZyVR6O0g63wRQoUDG1guM1V3Vghz
BywR2bC5ev5ewzlFvybMgQar/tqkQXQBKXRxvkcDXFbzAraBMnrua3JTtl+luK7h
glCbT8xP1tS6mI9NtDp15LHB8fMSr1oKGQwyTPoFNTWJRsKn9/vh+6AK6qNp2RkA
rK8j/1QllB99STxwTh1IRsoYTU/H6J5aNn1j7n9x9j2I0b5ZC5EguHZHIYt4A9t0
6/HABlb7J5femjqPO1u+ybibRaahNnmtJXDNc7T+gdEJKsWlpO1i7Kn3QXFx/T/T
pI1J66+Bqinmaqlb/rpjaxfnW/jzKiWsGFnd2Qs8wDRfUVzgSPb/KrEiP4PBFND4
EYKcxyPr1SyoWgqWjJkl2DE00QBcGc1Phf264kqBzm1nfLjAUGlFAXjxvPLULlzr
GSz1gtWFhGZqf0Za/QFrSxvIm/Ub0UPeG+atW6dZCva4nyHrBv30iNO8aVsdRD9U
IsKDJCqN6wwT+oTqBmNYTu/HMA4xd2yr6qpwxsA+m1P/jan2JmVH/+/OvO5SV+j5
GllAsWXQ3Twb4MnKmYUyN69jJF7Sqq5WrC7UQqvg46503LUkdis/WbCIgjJKL8rN
dskMAVFOpViem2f/OcYeEBNGPLINU17aYr8zlS4DCZi4DUG9uuQBMCxn4Vi8ejXT
t4zQw89K9KnUwEhJplOkSl9qSxaZsdyOtF1BLUsOOILsHqWEnoicMImBvSlu1SEC
9HwsGS5oQDqIXzaWw/uhW5TEmzdLQVKU/fU/vXd1L1p3mVNxkusVNu1CKnuITSjw
WcKV0DhQBYp6O5TTzQxpmKBSDwu1P4+A5zemv41DpO5EPRL1Q/xt5irVH74frgm1
4nOVhH9hZ8q/bWWrrp1KJy56iABhnXsCvmMTGI+k29PC0jQF89a3UNLonRtobkoU
P91V0reMpgbCXy0p2sw4X5UQjUcxzfyo/CvxBYnU9y2NLtnkLRkEe45yXf+nO4PV
1P+Wh+jh5/nuM7DHGkaNtUZ2rd8klhe8WQ3nS/cX3j3EyL+bNfYHLoMbEpd03jjB
D3wPwaYnzrKQft/5gyx9Gg7QzKrBP6M2SadS13hTzwjOpuqqaF7utI1TEGThqJnh
J/Cs/YqxBGcSPQdbTq+biAudG6aF7jZtZINeT0AazWeY8JBReshoYweuF+DM2KWR
cq0RUP9t8rRzUoRCBS8VFOUwnIdU1Al03/QCpn1Plt7BwjHwz5eziRPGRh3CyXaq
4JkQ5leNlWKnRoeMRAeqxjbL+XqYiO8FytM3mAHedNtooEorcpRT2T5B9VN4QoU6
cHttYqOp/mMyATw5LmV5zt+TxlfI0c9O/VCTvfMfAO9qoMCgMuT2+t4Rm5vJ6HAn
XX9RmHvOH3zKeCK9ooUCXmrw2xtkhWLuSJhrb6YkY70Pm0gZpqFQm2tenGCKAun8
w2tGYKkeeDSJFh1X+xE1rxAl1pq8nxTrXj4uHnkRkk8Q/xSBcCJvBdItNI+coEfT
0gvBUPBWmrCp98ueIp2bd4D7EBIcP8PKZVoxjp9vVv83VnM0BpJ6xSwFJk4bkh3+
l4SN6oL8RWvvBIH4j1EJhQZVFfpg/MX0QBQ1H/Pt1wRhFaLVHraEbB7pQBKp4KhW
+pSwJ2C8WODqBPtzBc5h+FHFZnB+qYTCeMy8/P9rI+utJ+oMt4enjBXjVwMjAglP
ZA69QC4MH6ub7tQNcSf0Ogc4PZce6+FcD7u1zckOm510122FMcCtrkUzoyNVTcTw
mtz0R/SuoCFVBSyjpXru2cqtcOrE57YVOHKJJU5AKTxxK+m8xxVzPh1/TZbnLLNM
TzBi6VHJdbznFYuzILnq+iQGieMaT5vbLagWt/juy55WXeLV/7kY1RfwUrxllI2f
QxpX4sS7ttTYOMt/8iubsC/kaIE+pFGcfMbQYMh04jP0g4OvoLcBM28RjoGgV2OO
I4DMlRujGAorY4hJFgC5rQK14UrIBp3HApm4A4KNbi4Z99XL+ulxdyuQcdZR3vBz
+TMYrUBWii6B00+CJIWzCYfpoKEa2Sj7jrt59P29Na8xST6HzKNO1WEyQfZMDzlM
J+xNw1cVe6LKq5CBZouMF13dYIMYNBX4V1aWcYucvKAwDDlcRfBaiTQfjSZvjKjd
jufPw32QFbJorIV5zJYcfOGlwFJWWBE0NtoZ5nliLvtXGN63wTsZ1YJ1iN3ndOa7
afdzLEi1TEehrns+CfsC+0Jd3hNLWGdgB+057vAC9poiu2dPALAhhxHJhrr6aweg
K4y7NzQgBIW5UQU/xE2XAZsyqh3nlR0lGRhx9XTYmxp+iDKTF0SKmq7uIyV1E1UR
Mtbq8cSGAgHyOZdg/9Bk/0n0xsoxoqwf4F7Qdk1jzYnSTw8EacsItCmX4Fd8ypyV
akp1oHbfB6DVokxA4+WBmcuf4EQebRpVPiSV4Pmf3Ihr2r67XOD/I1doQVjTVeOZ
v/zZlPpf5c723lAbsBBNoIS6+/Qa3+l3k87DHd9K5xuskV3U9w5eKJHs21iplIHF
ad2pbTtEk3gyGDF4EbJ2z69ohOpbymqb3/1/7uH7bDtaisE5SeIVw1AnXAm4Lrig
pBMkGOqkjMAnO78GNKJVS1yEiZFOmUnebU37cf32Z7UK9NbZWfkFvEF/GpkTbeUD
B2FFfUu4KxPtoVsWGvfmviF9w+0y5wwJAs2ElmzLRbmgdOTlvRa3m6COeV1Gkcme
FGclc+NPIlvlq0Ojyl2pwfwbe8xYhgZ+VHGAOeToWTQ7Ym6dmpXkG8DNtHYFFW/c
l6XshjFOUf6XEdrXz0X9ZnZCS4WRijKcne1QjrZvAIsQCcFdcuNpcemjTiRx/ahn
AMTb0cpY1PHT3Lll995sryg8gEIru1karkTzlboLAcAa/bQveP292n0qYg7ao4UC
hlwQdEdEMg3DvKpYjISOHzXKq+X0mDmLkPexYaOJipmM+AVn5Ejz6l8lRTuFin1d
/NLi60mKXJyIArbqqkxrYzQer42GIbqFYroIehLTrPIar50LECisG7xNzWXLJFPv
iHGRjVCzWq3VOlRMjiG/xSATOHJT8V550VWA+QC38gviOKnXAZOrK+UI2jHNlMRR
nXUFWBVXJy6CiepT4o0WDhWdMyZtSkGZVsR9ckvsRft+jXY9qqcjV7favaYQw0Fz
uwQluT/oJ8kT5PtRTnDrNiq/v1kzUTRof3D0mRsbvwHN6ts+R07tGyuab7Ml90cl
ubc/mpu0z54q6Q5bk0gzGROXYj9DnfE11VQCIAwMLDQjSIQqz2ZQgFZQRdYADwFi
9AozeanWHQv/s11jJm3FGX8nWhmRSddeubXc4hu1ARTktQ2yYLD6kHy3D2VAFIp5
4L7Zu6W+rDd0+9mMxYWiVsHpQmVK5yrJNh1N6VfJOXj66nwA/uUAQIa6YabzDhCD
z1CqED1Lxwr5lmWo6LXcVC2TNx2gSnnalhK4uRHP9ha/Di40uQcZqt3/28/OWfCd
y3UoR2pbXEv2PL4hsOdVKLnSXM2OVKy4kqONI7TV13OqjvH31N2Gr3ekVqybLC3d
tRl/O2ChvIq3xLijT5IK1SWSvt9AbjeZDtsESj0t2tOfXsDa3ozMvQvt9ujcfB8c
UEOgs8X9ZFXPZopPQT0r5CMTa11Ry+O3lW/8BzdhiZdNotmJKAKKoYrD0hs94odT
FV7ovEbzemHQ45WQL5O8I77pAM7LQb5gSo384/DtZZAG95pvksPXWSHy1it3U8JH
FrTQhOKsTRstww6i7aEBSEbxxYvz7pRji9OIJ7XKk7q2gG7EOakQzH65PXnrDmQZ
tA3Ek5BVzeQsR3nrtiKbq7GWYOOO9cLZ6mZ1lkgdHngBAbUpR+vS3g+Y15QTp0+T
Fh/lY0raw/ucqsn6OohA70lhta0JBjbEgCq0UmjdGpojDHt0akwXSIoL1fmllMJ8
5FoVSDRUnzkcRx/OMUz52JbRh3QougY/QxXweXDMNba9Qe+pBTuOc+k/CuhiS5h/
caGhiH8b3cNC8uaF3NNSfEFb+BdEchxRNwJtWuOlOl+cbIxDJzfvB4bIcSW3v+ak
dVYoptlxG+62txFoabg2PScgI0GVjcNHmHgSyUjMxcXd3uKnhvjgjndmie1VY52/
8cbP8Bxmpu1lAqAIp87s0M0Aw0uLNr5kcFsVsVn11j4aTAGbG49O2De3v35VaH79
oDkE1eOAR6lh3OVwCm/ZjaY41Mt8sf9xsjahoEima8xQLEETwSRMLp+CA2IQ0hRq
5gtsmJzVmhe0X7jwo+LD7tiN0S27743zB4DzN13ijUSb60NeGQcDPAodeLk5/rMD
mdepK9L97UwPzyDAyjVkT/QVYiYtMkPPqPeVaCKKI+igfOrVnweo/JPWHVG5og8N
BwR2iWE5dWLJVKhlRL9Ufd5hV0F4/fr2VXP5G5Y/DahJ4mNh4qLw3s9WvAgZQHXC
OdLh8K8HBrV2q1M5Xr79kewlEVdZB2DXYG8whVInQE+6YhihhN2tCgu+yBQF7Wga
MZ2BgbwSM6M5fuTkg4ZCvrHTFL2ff2bj9/JtAFuEfiuFFwggu+VAjvtO7uDzfLxa
`protect END_PROTECTED
