`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JHguAmZrpet4RXVhYahHBk3H5SvbwANHh62lmn/8SowO0eDsXc9H+zYvxgdbqbN/
DTcOZdKpsE4JY+K7lW9NySOU8epp1yIeJ9KcsFyqsp26nANcHbFFiqGAJwPkZa3X
lrTcbknGqjsJlx0G7JlNV9DtANYJFKrIppJooCp1zEKSSG8NI+GVTHx1tYB2x6qm
aSml2afrfaek3JHVBi40gM3LMZDv96A7rqxZ3KWYZ+mot57GZVYn81kNuGodv6e1
GDfMUACanWnkrfDk4xF89whAQs4/CC/u7A5os7IZM5fVqEND6g+uat2tEy+kOCfT
wMPuO7KcuCm1Nv0dC1t8FkG69KDj+PtT5fwPvu3xHVtrrj4d1I9MzbTNmEMjK3jt
kn+LIJ4C82p7TG1q7Rlwo/ssKIySZdH6H5FRD4DNt7NuACBPiWdnStUm/CAtfeSq
7+W2jGj6HhhwDC6in5xuoS90cvWSYMbBDABWsvc4A/KCg+xcLtsIfUzrFI4B5UmG
LzU5KADXG6QB/3kYel3pNq/+kXmh5p3m/tjNBKLcflvhySesPHqpDxRqyQcFTqfQ
OV+Nua/+RUBJNO4z9PIaX+2RRJBrOunWEFR10qq9SbhDX6Yk++B9swXQzcSSFdeK
fUSeqTjVEeklqF7i69/v44rc+mvls+Gm2DNubr/SiFRw52yZpzbg4+0pxwwHZSDp
ficI0+DZeh+Ii3AIbOPDA1S2EJiEEv82juCjw8o7ncjSamsyArPRfy3yOLQRflVy
9J+JvYm3vMdoZqtbuzc61HJle95gNpIrVk0c4dTfFXCa2+6M/Dbc+jwO4EKdIU0u
1iWfIybEXXXIHT9EzTiPM6ExHdCxiDySP2Og03byyeo2wPkqkhvxig/CbfM5sev7
SYt2KvF2WRPDKbBfS+OVDzAZQW5yx3kWp/dv+Ek2iqeC2+whi52b7IT4ozR3MVVA
TvBVa1eQd0765rL//KlVQy912wIEbCnBDovFGUO2VIZMSQABUOaDah3cw6nWJwMO
MHqQns6g87q5ruNlCLC5xTMeBGCp8YF9l2LcphjechjwlOUFfUPzqahgk3j/Wdyw
7On8SX6NFS/GhPKln25RJQ==
`protect END_PROTECTED
