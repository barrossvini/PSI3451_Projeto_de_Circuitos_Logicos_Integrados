`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Aab2su9fp01DKoBazwcN65rOxI3mEBOkvysCuCBlUNxf6w+AMd7QOcKNSuZqSFq
z4qlZ/A01m7V6PvP+5Tt6g60wHv8bwLtlWSpYYNDDkMFYc217qq3aoxX22Y/aHhU
hf0Gre8m69pnILVbMmG7JLjNA1knNBCTyDrUTi48JP+5EmXoBO5YDZ/NVcX8BTx/
rmaslqtbYTFYHmGKS3Wq4vm3IVMevb0hx15405gi5EU2GWK3GHh5zIDUXqB3y9qW
21eDvERBY0IOYXBMPo0B/HzhmPkmjgK/+IMJfXgTF8NYjrhflGZd5pyJYhlwzfNx
thsy3LXluXQn/lvkoZDRBuIdpyOGmmDj0wHEoM7rF60J9CkOBY1ImoKHZ7ry5VwA
ffmXSj2xbTGIA4wc7pXce24/xBd70GKAYXZHxw16blVvjxtcLGp3APBwjq66XnA4
qbBRmKDd2DGGJ3wP3KpeENv2iQmdm4WqHXenlg0cznazU4tAXhDApfk7Qoq2e+VU
T9AnEOvHbx33y5Ffio2K8sjtcH74Zr9QibnvG4npuscooAn53KWxVscBwuLHdYtP
whFTcWQsCJR4kX+jW91Seg==
`protect END_PROTECTED
