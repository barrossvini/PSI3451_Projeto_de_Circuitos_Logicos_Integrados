`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cp9Pz8EJwOI03H923VOo0vYPxQlCzHsV8Btz2dwFS2uJVumEvgfhXZceZEJYplhu
N8DSBbqhgPCIQhSKru7oHq2TFhva6DO6gWmuTAgZFHksHbMWm8l7q3gjjQMkFxlp
XgSGyKwtLuFUMH/465+GX3GRHHBbY4QCMYzrk9WMhXmX5egd/i3mDUfZk923BVSK
um++6s/m8vPciweI6U+JQ+qQFX6+oPhKMWDxCv9AwYttpXy6RskI0CMWPeYlffdo
fghI1/sggSNxP/v1SoWvEQ==
`protect END_PROTECTED
