`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0eazXfxUjZZswQYMH/PepFfJOtjSZ+9bXUEeEPrnQQAZAuj7vW3VlU33n0GL+gw
iyj2Ja74YC/yu9RNOwVl6lzltq37yT/4FQKSFIVwNpbgCV0BOnudimjfi05cFuwA
4kXdSJGHVALkmJQB1TbQmMtZ12lsNennNObBjq2g5N3mzhSeiGvgrMB5Gkv/qT6d
drE2RzD8vzovO30K3Ic4Ogi9Wbw5jYMgQp9uOzjLzmw1ECYOHc1eqrUqglwRYD3A
OzKS5LTsUKX57/u6Jl/hXreucRDKhZp/au3VYAfdGwPLqbIIwk8h7aXgcO+Nu3YH
Gz2Z2Tq8GDI13+/COqPwi/xyFP69gyeuwyrCnjC5BF41iBNaiTLJL7Rby/FysCPz
MDljqKe/Q8R8kh9q2tcZSdq3WO0Nrdv0UlSjyHZh/9lsknp0x57Oh61RVC7uXKE/
rxLQHLEIrTZ7IQraOlzfl+m8iz+bi/mONZbZILDuTH/78ROS8Z/0dU2RYHv2TFdU
bMxGfPgRj3BkO6j0pywYH0I6KKqPbDQrEP9A2AVXa1g5CXbKmOk+mRnDVvqvEQRp
upeIgsZ1YR1tftvNCd5QT4Kkexj3ShRKMJKmZWqpO4P5YWQaQ0NKyVkibQNADMBS
EdyAc9zzfn48rJFkS0C0x2wiukCUVClYQguBstDBjVQKPKp9HHRAVuYPifDkpCFU
mze8F5FDlEr/EjlzfMg6Wj/oE9NWkt0WbPMWRogX1OZl3iQeuVpfAh49webJ1mwH
82fsA3H8LydjsEItNxs8HWsl5VYqPrTqbg/9Jdn2CPa2nzC8ntUAaRwjq5A+SeZR
NIXdX2vR7uUVyLNg5hNozDxRaOXaS4PE/dGnOHW7aHYlwaYuHv/NAHuK/bsz1BVb
wTlUwvh6zhtIFMPPgpg+2rI2v9MQgcz8jyzMpCfrjVbCTtIOG+0KR8acWvbEedm4
+nC2p5fdpYO0bTD9Kgaufa16z1/uVnEN6+7TDr4EaqsjUrTubhoRk0E5l7QLdLLA
U4yJ4o/q9LItcdl/JQtMHD4kYxVboRQPi2pC9f3itn3sOfQLcvsm4r1Mikk+NTed
cvVCU6EeV0QpHswBVSKLA1Khlvik42l55jBlIjfHBsZIu9BR+3lvkPbJvMZUAqKy
1yNFT0slRwWzgpWskOVOF8qqU83ZjPOdYPHhN8UTLWgaC8sHGNftCy1GsMwi2B+7
djHnaW19D22lz9XJZhEv+PPp+V3M3XLpy2eW/TjkjneY2vKprtYoiJu1EQQEd7r8
bJV+2r+iA5/JOguJx/znjLrpul7rAjr+CIS0XxrCkEAmJchY6uqsTnerqzX9uH0b
8ltaTwjIFL2e1p3DOpzVtrYsFfW0mYMp+I3u2OeVBYrI9hJ46c3J8fZvShYnE2NU
NOkO+eKNbJD+dh7rmbxF/pkJ94rpljhT2rn1OgldeyWfQeLWIS2+B4b01q6d3XTB
jeV6ZJ8Pql0W1ojJ1wTvaKa/368uYizyxC5sTJLhVQ6Ckq/q2hf0u5xFjEBCqrDe
wZ9PhAZHiCZQkq0ZSXUcg1KkCq+hLZ8JKSSowFMeXO21oRikc+fYjaSQo8hYfAFy
mWikH5R6g6FDoLrraehfdY0qP37Km/77zdMFFTORl6zenLAINNLbWnyFMfypcT0N
20MbPWhBVIRKjBtK6ppvL30iWX5n4fhmgWgGElTZK3ypgr33NL4o04iZpD4T/iLq
gSHRZTAMS27UEalAQQZSRbYGHig22UMwR8V2/+cuhzCycRt4U4HQNZYVzOVZ8eDk
9P2RsECGFg/8ZixEOLyuSA5IgYBsjFJmxN0UbIRF0VZT8PPaVcciOM4rVobADz9A
5vkr0H1J1I3a+r72euJw6IEbV0rs9ye2j5S0VejQiXx4szAYl1aWdJoFUp4JRZai
qxEy9JVSLgS9PUimBK4kbekh1Ixm1DTSwAaRHkhcL7+4AyNV6bzP3ZyJCO41cusm
xvQ9C0gy15RZqrUcYyK+OEAqdRsef8mhclTiedh2ObI3xT0Wsvf5Jm7DJpgJZWu5
MV0ElgoAuZnEx26wj17aiTqP6fuCOMHcipMLRnsO9Ap7JDOCMcjKMRX3RpcpVHlb
BKHMpoHAP8ednARtkXL+Fz3IisBCrRAF1Q8Rt4EYBsdQ/gcTHjuEt2hMUsJrK1hy
tFRdqoF9VMtf23DMhKvVnUq1MAk2W1Mh/oRRy0TAulXSZDWV8pbPqljENuIzlPg+
8cnd6IgjDh2+QfV/5p6NHeqRZWiNTi+khbiY/bN1rGRiAOYOqQhpyUylRz7MB/Ss
PK43UPneHKyd3xLhQCVxE1DxNcM72i73HItBa5ZN8gXOZMR/8hyvfS/DR962HWxA
xlIWnPJm8hRFgBSYSNBsb9tcEGU9rmjgYj4xpCseArc2kHAeqDOvGq2LWWy6lU4b
XJatkh4y/g69rqeGD/VTWRiNklcX7vssJDHebQ2TqcKXDWfPTvZZQmtEFccEeb/8
4mcbfuaFe5NHTfx7B9CCFg==
`protect END_PROTECTED
