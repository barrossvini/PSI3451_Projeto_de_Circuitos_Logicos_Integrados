`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bPpRmExvZevxgSMAGYqwnazpyeScQaPN+y5GSJyukl/cyHkJa+ZtPZ+9wv9Zsb3Y
7HGtn6VEXEzInq+AOJUiLcxuyUMZiXK7pSlDOM8ulEBKHta4OM08mGUfOwiAI0ZV
+kiwz/GeGJfEDWiokgXJUfjw5kZdYYlxYYS08Le/Tm7eRA0MuJYZzqom63pSJc79
wnT3aFxFfZGl5/4prMyrKhpqRn9QoL3gLwGAfc4fAbtF/+iahc1bKgxMQlRmT8tk
OWhy921rKQ6Z2Ueuh68U040RNbwuDeyVZkGlZHFsAC3sUkqgpmUATQ7sFHx+x0FR
MIbLGksn6mB3/ykHDMFpXXW2nfhHtnVUnNafuS8Oge2g+HFeWCVpK0AiJFQBCyoT
CSKRPbH5EqjRLwYo7TtB7tvt1sDBoKQw4nGtvNPpTsrGDLuUikQ5bbQSHoVFbia/
+Ici1/TCzl0yuSbqYq5jqA2pV+ekUCuQgOCmKgPZUeCu+pTqXnrkfzy7cGO6EFEB
lHAd+IQO847irKuOntgV8rklklr8wj3uWwRKFR58Gg3CgXDSXE6Jse43cE85Y7Ga
cUtWb/PwI98q9DwYvDFJJZk8KG+QBkVG9HRyluPdC7u7q3w831R9zRnCb0aFcBJj
WilQLVT2O8Svlb7LtxGjpV9Dx1JsSrAYrJiDHAe30WRkhW0Wd/ExRrFYMjSrFz15
ifxeUt82GMkToUDO7zgMHdLDkhMDQxeb3/1jgpp/ihb3D4sAABojk1D5UmbU6jv+
QWjynUPNb2IBB1c7OfdQgIxKRrGt0NblsmtvpFjB0UKSh3zWc6zMnHpEefwRYRMA
`protect END_PROTECTED
