`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lYCnz1rWj1qpJxZM0ZjttVuaqXa/Q7KS2FJdh3TQ/U1usmIsiAtdoAR8bz0tLAk4
9RF5H8cx57KDXM5xjTWpZz+BGP2XtlNnEyOuZPycTlkAQKtBPV2FJ0k6OQkCRoU5
GeBVKOCg7j+iTBBC1U8JeTDKmS0zBn9cqHF4dJY1fEIStL2MkHXgJdSDZRXNJ7rP
ApQlRssLr3F44zBk2YLnM7j7ODmDwZeWLVlGAyUl0nta4WAa6/dHjb12PJiMO1Mc
mVQkoPJ5an1mYwRHPU9SAgLy/jnlc2xavX8sAJsTITWtFAo0do9zvN6XVv4Hgobx
uocXeImp6DegFHjhFcIhkMGFvj/rKjVAMjGgbiUlogIoA00VsM39+3az1HeN7P8h
MW2YsmpQqhSviaQddaLKVW0LpeYZzfthl7nDafJqnAEQNsK2Uc10zFbjbeai5kMt
s81i5vBVYalFDPGLnqjSzVAxtn0KnRuJeI9oglL009hM2+6K/6bpIYNnPEk2N7jb
tc27Cxo0wypLqNI4tboq0bKE/vbwIjzcXMzkxfU2fs8nkGHIvjTFPMhqxx2fvq6+
mdzSNcuL+jt1DsuNz3hBLs7VSQSpE9x3Ec1VCvaufq2Dc42jPNaO+9u6rVEV0UNs
ofARj1D2F+XOOmXgnqayiuoQ1sHNGsGrDGtfKJwAKaIqDukJpnJMpx95lq0Iti2k
NpL/Lx61kbq+8Z4QKwxKakilkd2+yq6WbgIudEtdjqoSC3ZKnc/7ydhQJ4ZvSdz4
ZrXvonOk6K7cuoQGgcEozWUhvRpkf2l3q7EMjskV8sd6xYCSytCDqypuNkhB2YB/
ASuHCEQxily7n+RYoS39E2mmh6GevivrfEDhUgEVc3shjPYdGH7ZN641yde9CH1/
zlcmpUftVNaF18nzz02IzncO/KxFUpL5u58/msnfwlYyGBt1cvKg3zVwLYjfo8Fo
rnCN+wi4QOtWTGUyLX4fBngIA7y6EI0qsRhwpnaTfFt+rY9xY/7PCYAbpKFIB4Yl
teq6TIqwrqwAjjqSdBz/2yewzyXukujAZtowcoCWyYkjtuDXFuFYg76l6dmR4BbE
zI3ZAh1AloTn53+TUJJtclTKAI4fNiB7Ub93EmdIXXEc1G/pOCu7ARRm6+bizYi4
SH3P6BQ3xyLLwIeDWz0sxBH/J0obs5/GzcR21NB7KXvkqWkepxOmshqT8PjIBtou
mzTHOJjmBLf5wwpfsPC5jc7FKlHIKQ4tr+1219rY9z5jPg8xGhhaKaWtl343crHL
XueA2yIITaOuuGvwcWC+nd1qRCtk+/UFREyaWLvuoWZ01Iu9Pts6g3DAqzUDqWL1
V8kHGhjKTz3bco8BDU1GdgvBXvug7lIqNYKVLObRVKeCn7YX7HUgBIPWyHdT3i9F
9VfpcGH1tSAXTrlfP8j5eFD7EqHryDv2d1IHTGw1UwO2qftViCCD5a1hpPLvLCd2
CPGAnk/OmpRX5Gbr0nClPu6FjcWeezLD84HsE0qMSlMvlwPg4CPb+fSJ/kdpIyWl
wzk0Rt9LkYWvbtVpnSKZx0bVZArSTJlAoDfTfgT+2lCaumg1AXeNWG0jVhDh+GAP
Ps4I5mL+GLAJJHZXAROT6xb9xXo2lWcp6a7HjiDZyWBKqY8QJnTiZjQRpSU2OgiK
6xPhgMsjtsLD+qls4GbMLCVthqx5HfR9HiDG3wR/qSEqvdrPZXYYKhFLXw9XM/Fc
YQoo7MTzG5UjdjtZIgWWks9Fza5T2cTys7CeDsREW+C/7SvDFSu6ErVlc6O4AHiy
iLXh1zuFsHRJcXOO3q5Bq68sC8b7XCpF5dwi2mLAIo2Dz83IrSjgshIeMT4zQaFq
mz3DCdYRLBVqgVM1hFLnVoUh+aNiCvxEblHmzO48NxKHZk11BmihCHBFJSQlJ0PJ
ix+m4H3eyTbH/EIqPbxP7c0+Fm3fRDUeXuYvzLcM+Tn89scUo139ElVbCjSmkZ9R
h767D9FfEUHLLlP2QldzUEGXYTOf3n7jS1UmG2RVjFnhu+3UGsSoqUUCUZaCelbf
+NJ3cnM5jGa75R88HK6hOoxXJJuqwHy67fmWQgShVMUyKF4qof8fFzbrwS2C+/JS
mZPTHTBJzOyCcj35fyC4nUFqgXIRC97XmgC8tpB8sha3XIJ7WFiO4ZNACQEwJwnh
v9vVmOBt/Fv2b220fkJ2ohewdaYyeKxE8Cpk9npR+3A2fZYRc5SUOzY6pXO2LxlR
hX3IQEOoqLGieSkT2N5EHz91wKRlhx2t/IJzf4I1vQB0ZvPzmaEhyAL68slSw2EZ
BXBFbPBKWb5/NZtZ+UDlAhBaWR6Ba4EIrFILBF/DKz3Wh5XEFga9Pm+Dz5Gu50Oo
YnBlD7k4UkueBmNoRgpfJY+9REOIuDs72ko1S35vNlYQx6Ng85fBUR/WC9YnKuvb
KtDH81MV8OYShf3FVshCMVdGJic+79p8n2TyR27Fnr9MMdb5Oxlo47RaPiSmZiVS
vLsqsI+I2ZLo2RHzS8bIPIBDQ6jFsXoEegJ0bm5t4yeYOd8dYjSla8j4CB8snY1C
3YPuHcljmII7JN5P/6mDxtKk3f3hoCKO7cJn5ly5nFfggpaEUweHFm/gUn6lFiDy
8ErY9/7oF1rAyWP9daKQ7nc+XkMu1emxxsCpltgnMIy37DTJY9a8UJDUb7gcVQ04
Js3K1y2crQuB/p+FEArQhU+AEpjlhM390cS3oiHuWGNSh7ZaaOfjYVZS+olptFUx
DSCkykqVwBWQ6BvdshqKYO1H0if7LrtjJ5rK0PLzE0J0QTGYmyM2vqWTs1+GjEmC
5YxBZm92P+UIFUES7NzDuORcvBOSj+qmXPBpwgW/FOZ70WcALsIXofdCvGXTpy2d
WGeDP7M48+zHJqkivAzf7t1mFXdEdL1mnIgHmFcXOlyRZL1FYnC2y+c8nodux43o
7BrgZDEh4kvCY+sC3I6Jf03kek7KAsfFRP3Vxc6Azb4vH4qn4Io94H4oMqXJ5NSG
voCHN64xg//F3c3qPeV2y1ZqOgr+SFmONDNHbvTP58ZP3chSxLzCamRWTOX0x/Fx
RasGv/7ofwozbk8teSkf6MPp1FGhC55htmFNT/sXise3w7UCJHlxaHR6U9lfvkiI
fGQQzhWStpFaa7L6INYjz8KgZyU3oizd21E3LislTsAmONs13wArlxZ/8pTY2Tg2
caFNF5OVrw3a0FEvP8EH3sc4i0fXqoQmS6GWSWrqEFAUPbN+pH8w7/lEFsCP88i4
p9bdyGqKYhc6AL5HXeXrVKDSVNjb6gAWxF79G2lo2NTg/eb0gD9cn/itG+ra85qY
D5cxSKQJ82LgINtEnKeRsC8BMC5IwsuXopRoQ8GVgFnErpOluFg7irCqC0sB1GR5
XbZ1kGkx5cNzIGTKk2S3EaNcPz7vorWE6Y8QkiIoTNmwfY8EJZ6rxmUO0QrJClMj
H5whqdbwlaZOK9hmZxWEZBE8RL6yj5TxcmVxvLiRewhgUQxnZwCw3/isSYG6kK8V
RYDBQPnjaC40Pw1c3uXJA9w4kkwou4OH5qYkVDDlKwzXD2MyCVCbltnvCylISgxV
FZJgfcU1mezkcSKbML93vD4Pk6iPDaEAzYzT5HHyqCg2VBSZCjeswvb0S2+5OKte
ZzNgyEq1l3gJvitG9ptCIF4Jsd9lD8ETpyD5mp0420lurqjfDbVa54Fm7mgnKXoW
V1G1M7QUWnjrpjrHxXf08mDiEDzBYyKcQcBywReEDE539FFCH7ADY5iyMtcwPmdR
ovp+Kd827qjelcbJb9OVnc74mwTdaLHG7bUZ8g6ROK7TklacjZKmYr5diq+oPk+j
mXf1cvJHIVGRsC7incOwGjCk3RILLdIb/IOIkQyvR/X+4aAi/K19jFTs6M/mx9m9
k68f7xRtAhjOdZRDJAdjYYs8O3yLeapqXazM2kuDU12a9rwfXIHFRI5IEhMEO5Je
oP33sSmK7oK3h1E6jVFZv+n6JSGANu/zmBkGtfG5o0HvfD2RVCPxiClPEyPQSfns
N5u4TxZMxHYiDrILfxZ/kNmOJqqvY709AbSJ7+kPq9qKB1GjfbnSEI/3ACtKNJav
dCo6ws054myV18PykioLCv2opri6vTm6qY5wJPZbDQuYKe/yzqXhiYYnrp9UaUQP
7ChuNEVRwAnJHlRTP7O5vJfaTdxjPMDyt5kC7/XKcEg1ozMcivFdw7uw3Y0m9SOe
6zga68WO0weLkU7gGLV9qWaLmcW/v79Jwv68QLeIzTS3tI9b0mNbEcBIbqY4EwNW
xQ+SMpSHVEscBHDd1+QluuIykf/w+CzRFOGzfpry5guOOTyD7TuC8zNqhHl082yq
kWAPWh09gMqcSntHb8GqKX9/VbY9phhP9wgrrc/fbShP6Y9EDc3WW/qnACKQ1jqd
QeOq7kH/u581K1m2PKO7bNR7Jl13KhVJsuwdnJ9Fd1LI6zhDQj6BDbsZmEV+XDNV
EcwY4meqchkl3xCfk/v6wSpS7vhor0Swz7cV2lIsFjYj1FnPWhD+dDqOCmcQ/xUb
MUqetASl8OnL1lk0qmCPYzBnz9oLrnpfTaqi01svw8AHlHq+22NgSAqAlOwSeyZV
y7fMtHDEyJPO2y0/cObMIg==
`protect END_PROTECTED
