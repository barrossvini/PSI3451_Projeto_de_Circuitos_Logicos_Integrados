`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4tORzVlZbGct0nHDkqtzwlEZAqdzjkCvLrDRe104FDTRPNCAWX+J3tXiB7xxdxSF
C4AH/B0bXROEERbU4XylEFYpb3d2rOY9FySBAtBom4UOFt4xjTD9rK6HF2Mj+QJd
ukt0vDAtTLyCYXsrq8SwHk3nCNDlkNrvXoX2OU+ebs/k/CYUFlKP14UZ+DyvqQeU
faaA6Ddm/LJtYNVGo51A+0U0fwRtR5TI9ciSH3MkHXaTwpj3W2XblF+dWLorj2ol
/GZ5l4wFlZEgsBfDYOB4o2bhgv5aOTGo9QEzXAyUlhhW/Rp60EsBYH+ERqfF6fMX
xF/FVKKO86UkwfsZZEnCWTyQj5CgxbDzXBbbkz8IKSO2l+OU8f12q7eKhjKZHOWo
SjqInssDO3Rd1izqpbWsYDleWw1RWX1pWUj+J2VZLCKRShjdDjiXIq+v+7zAm95z
a1LohN/WUFL+aGnz6tByojBjn/dy0iu3COY7aDC7Xxp3o2D1CKmcrLeMvm7+mJ6D
1N51jsS9u+X9UteG2eqYrHt/1JU1+7rpr8Ecq5qBjvZAw+A/sqm6DoeSXuDuVmNv
RDjttBEW089OcdKMR5aqiQc5mNjLcPkDlSpJoucwYld6b8Fd0jWFiPhHXG3RYFde
CgkYj0l+fdc/HsTLRlobeqfn3WiL8XKrS5f6dzH8prXhEa08YCN0IzuwTdtWu80a
nBv9Nt/1aenn3E2QT4Gyv3RJ26erTTu2XD0vndAy1fI9TrCqWOmN7SskNAIHymNT
rHYeQIZ+01RAA/SvuAHDcOFNPun94lCZJsahNfhQoD+MPUqBWNc96eUe80sKCGno
1R1fUssphMvNF/BWurt/yQ==
`protect END_PROTECTED
