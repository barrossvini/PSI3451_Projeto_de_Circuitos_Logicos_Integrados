`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6jLZW6Y++CbX2yxxRF23QnW15boFOWWVRyGNpg39aVrzvESrmbhmOC4eD4bXlf6
5lVAqZbC1ilClmn3twMHFc7jpAY7sAT/e22wNqHFuQz/PLQUhKbunrFsAyZgvEtC
RduZOak0aMg0jmsadTi37EO+jB2xj4YspjF71504SJC2JO9++piEocsTLOmikQly
zl5sejdBHS3uZxBwuhmsHBLguFKt5gjA8P9EbR/QChpdygBo5KE6fcFclRIZSL7o
utLgoWILaLE+Dk1HAANM6MY+L0CdOCeMV8AHzQBMG5Rx3W79valkvLDpYnrHcwF/
cfYgp5lV6X01Nee0SWXxtQZ+uimAEJ6AN+sklYGVlmZ2vf64FXEccr78dwQaR/I0
zZnc3aPjezqz2EffRK3IaFFx1XaHZ//KkPxDFnf0gdujx8IJeeOIW09c7AWm01hV
FzrY0EHqpeEX1pmk4f2sEhEr4Nua6KyDG2Wc0S5BnHN+nsBUogr071wx78D5KiJ/
+RV0QckDk1+hSDVh1LuAEO2HLGZdxAORo9G/3nxqGNsPyVFcgfaqVBF39jc24kc9
egWnJ7DIb3ENLfyWRx7ANE+K7DK0T4Ax9lmaOdU1rmuKiaSTzTPEKxpHvVjMg7HQ
45LbndNYzH8KbD28x64lEK/pgb12cJcXeF2OEkM2vuzxDB9zOLpN1KBeVPPBEZ96
L0IS2nDp//8lQF7eO6FkmUN/iSShe2Nw6KZ45Nluui4P3jIbcBjXxmgvDto2xlqx
zdCtFUnP1lCKokBPHkxralKMy60VdDc4WL5DNEoVXPCr8KzV4oWe08Y1aKXgXgeY
YULN0vVXzncuxAC9ECmU2ZDH2zMcHOg0qvXLCrKZLMc=
`protect END_PROTECTED
