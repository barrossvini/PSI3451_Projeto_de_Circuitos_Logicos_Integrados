`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
daU50bT86n/HrWG+0wChhju7p/rI+4g+3kOJmE9Kq9yueA3GUG4on0yZ8KeuLTTP
TAJaWnLCe0Ihn37JuSclEWpkWXHncVTBD6OsGZynfM0O8gXTmxkfT5H1QgLhWb0f
ftqeN9cXVuU7mipHltY2L63uaBQHNhXjHwKVVt4XJk8D86lm6rKxSPzLRBb4W9eZ
hf7HMG5hW6S5pYfRXwOsfLoELRqKWn242PlbO4pQV94yJi7vb2c8WBMLzD1NHF6C
RUey5h9vayP6AOvDALdmlLKFBFt/w7LkrqJn5K37OOL3LAWgHfrW99YCF56Ps45V
wesgZu876WBRvaR1Qv2P2cU3Dq9inSi22X+aNjEnEkkmS7NGutJq1cirzBonMsvN
/A9kns2bg47wf7CLTsygHCgmvNaAhV84KcuPlsytcdAGaSoA8XHGtkiKkvcQrMyr
7XiIvdkNxt6sFsRemOfwyEL0s1r8riOoGum43FP5LujRJQRaRGIvz8EuMlpyQVL/
GQg/GnD+z8DZ0obCrfjY44LTqAy1IqgUJLcYtjzthr+UfCeH1GeakfVONotLV3Nb
8b7JbpNkqU5ZgKiFI84bWbBKSx3830VPIYZJhxPixgDQ43Ka1IBVYPtUPl5+1CSa
QJgI9SJ2sN1iXjKLxTD/UCzEcnz1WRO6yTENaCW4HLRQXsnNVP1LKs6+57XTwh+N
0nqhJTXd0Iq+sjepsGtec5cgClEDWRm+ZxjwHYv+YtGUUJV1ivepwRtskPhdPaLz
4Y8lm6VQasYpT0YrA3OpiZTnUg2IVysE0iqH9CayxwHUirrdLor/vLOCdWX1gWgl
AH1EIaJ64eFs6NkjaTqDW/AnpU9s8GUGSWjYCpoXYmv9QJEfeLoWThKNdDHf9hKm
`protect END_PROTECTED
