`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24N94SB2UoGG+9L5W2iHnyPznBAqNxs5grUPcqggmD+qo0/8xPRAJPvj6pIh7jax
GQcMNY7X4EGbm/0M2vj+jGBIG61ju49MI+yWhdMOwXu+RbOWLRYaVFJzt7tPDeUa
uNH+oHHkjoqicK0xwxjiX77dRR5svHWEjMyjPbFHZdhYzihEy3pRNqBaKRm/wBMV
6hfyBtrrKZ4kQyIrGhGisT3CA50QOu/YCEDGI/ocmI/meIwvcfbMrCdcGUwOz77J
4we7f5LhAMAHJ8pgmQO14ltcJCAjV0tIQGgHrS6fLT5PSfKxTnVJrB6SMNc7No9y
Ajugczc9BSLeJZ7l+1G1tmG9KG6ULM2NIhyumo8N36vrTZ8CRYTDg/SsLief+h9G
+8Vs32JsaKTv7HuNT/t5KLT6Wx45uaitogvbzC3dRTNPflynlF1sEHv8RKMgjqoK
xRirANTF5CRU+lmJ5/+GRG104x7IoWVGyv+78GZH9VDR0mAIxSa/A+ZLlyFs6UiA
5Z60deKuRedUQKzDphV6qJeWxdV1I0JKXHAjCvwOxjQnVQDeKqJQvEPj2iXznhAI
txFH1GFxcwmoq9Qa9u9Z7B8w8xtRLhT2Ect3bKe6GyoTejX32a3OxQF6nNgqUCOn
VrzJiTmy9VboTxJnMd/slIBOHLScsxfy2EH3YtnoDRGXTjoCbPJibNiT4Nk8Nm3M
+eAv9CKgu1MZDNE+AG1EcZmX4G2YglRGkyCRojuuLqzV6FhJOdSK7a1dEdDXMeO9
j5Yoo0rBIOyTx729YqZsPo7CW2Xk/5X1Iwik/bbXrMmYZgrxhZbRFXQVYPinHlbH
jizyxv/8ATqvVr6cidCSOPW9AZyzQANrlexUr1lsigoZeRgcnQhItPF8d9oI/UhL
+U8RG9ka7cn2qtzE+lH6ulGN6ca+b7X/4QVi069tu/D8k47fpNoz5HPRa9ZLkZQE
4XZ0cy4w0d6eFXkruvhokHcWjV7e2FkpWNyRAV/1wfLOO44T2637bKrRo3llOJ0+
gKigeOdDVu2sQBxQ6gRQRTmVi9aeF8EPZ1tvJsusFD1bhm1qKodhmNrCXON4hJI3
hlh7veEV80uB5ddBagqDU1Xb/lW8WMEzuSsgFUgmH0UOi9xOt054Z19u/f+JPPqw
8hvvUC3KC9BLZxZdKWwtkbIBXzz9RjcLYlsQcctTUVUHREn5tSHKMqtMIgdgoB+u
YSQmMGYtn1tXcWGLXI9xGUGw6byEYrG6x6vMGmF+Hyk=
`protect END_PROTECTED
