`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q8TPjOXaIkdHZGbdrN5EDk+PSNLYQvK5tr5/kzONltu0DFxsBcuEEvM6pWF/kskT
NF/d0xMfTEW2jjMUIWVytCpQwBtqrZYR1uAaihUNLHXZ05tUluUkY27vfVwY9oZf
BKJW88UY9FMHnz2G2sV7M3TwKb2p0SzUABVVEwSFJblPqdis5a6cFJ87UgW1PRG+
0xHkNhL3N57mPb0wXKvH1eY+fW3iwdwPm/LCOgdqMvnUuPXU1ywS2eIVij6vHLPU
PsFM7DX085V+CxLiuyTnpHhUZfAbrSVAz/bOl6ga5KiT1OAmPp8/pEcvx3vlIcCD
gjFzcbpvZHpdi9vg++fE80MaANbhcsh/z5TDB0C2EqGqPJwv7U4kZ6pixwOeRb2H
1BuHLgAKpIUGat1r8KR9JYDox/my2Q/A3avybWtnzsWCGm1pCKVONR1/5kO7j9V9
R2u5WSeI4SRlprIZV9mu9dJyvtqVjt+PpGCHeMCn6lECBHbWyFWzAqin98K4E/EG
mpTW26d/ieGgIoNp2OIbk7xL1axcIejat7feyMtV8uMMfAkXjLrNiLBHJAC356gE
svLj+u+98ysIDIJnJ9CVMECsEuiYqN97F7krn7XvyXX22S+sLP+Tgs5lUK5+DbMx
JkqVKMdaV/WOnyXOYWmnlTxzk2whwKSBvpK7kwHAxI1qdmZr2fG807cEuSS9P1DX
Ys09SBc7sLfIjHzV9Jdx+LnNm5upNNr4tRQVXJK+9ZqoA4A/0nQvDUM9jEJrd/hs
XG1i5vMoJPEZVbgp24vgYMOv6bGw5NKtZPu2nCvj/KrRswc4/pnx3x/4ZWAjlXx6
mhZ5x3ysXpgeABL/PBshm8VZ5CzBPALZWrc7kAqhXsXdIWj5JisaYZr/kuo/wRrv
PuXn+I/jkRinfVAgfEMKofrbPWOx2hfwBIdaJDgZt+5b1XComAz9dPlMe459X3Xn
Wce4zjuZDS/dL7ZMy1c7qa6NB/BMAAfe+RAPPjJR0nm21xx/XjWsc7xEqYeAhFSc
jXeKY5xDoV1MRAZO4G5Ltki3YASDxwZlesNL0yjACKtzPr99jqkffvW42BWH4qFD
tAjZS1+oUCR4PfS5EHWw5l/ZFmLkjgriC9RnyQdN6Xew5yEOzS+/ZJJeui17xok1
QBKE9uc63myIix4Tan2slJQjW1YAkiifDTG9gyqp/jVWV3RHSaq13ny4+6NQmvcO
/FhELAYc1qKYlxV3T8PeQQ==
`protect END_PROTECTED
