`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6YmUPNVk6ASG5b0jYfLPriTd1ddwTdA4J8wtUC0/3Vd4RcS7khArHx7oOw51/VRu
GpFFmJFyPfWXU3oaWx9fR2yonv2KP//f7Qi77FJi64LT9A3R3MN/nkAMN0ADTILX
xsZPaEdokhqvnvqifmUTAo6YnBtGxCDslrwTjySqn8KMVyL5ZizxG9aoNrICzPjn
kLJhpPZ1pOUOflWpF6AVjsVb+HmEmMLDGGXHqBRKVrY3t7Z0AliaBHBCvO3qgZC1
9mH5S1jMMdmIzRA1h7luETB4/A8slMsxYekykpgqLlrW4vzCFbffI45aOtlSR04u
SGB+PP5mhg0Q7/By31EB5q/M4XOt7luu+BxhTAs8ZMlNhWu1Ovo0q28OGrj46jzj
N/0uZvKCpUH0M9KknIgpm78M/VLShr58O8/3FV1jmxKjI40yBCW85PYo6b1/sNTd
QRNgYixt2XQ7/KHDwKX1P99H25S/C97HGnRtHorGIhdPlOOBMBD+D423gPHch0yR
khW/gJwfN6VaSAvp+FoVeiuMUBQYpsRea0JMliU+IPFmuJpLmBVtfDz954ASr7VP
H8TgKHArZcm8ux3g6HfG0pQB0LewlyuXmablOkCc7LWtrfSi3yZHYUrKwz8pgj6W
eS6B5gkgOf6M0kB+Oz205rzZPqsvxvJWm6Cxj6JrZuxRlkty7zPTWPA7Rw3GMqPD
cnf8ghf16eASfndqzW8CeCf5A1PINZGvxE8dT9AiYHWRLX8VHw5kelHbfvdhOPOU
RBjNemGQFKxH4jHf8GiUdZE+KgVbxt+TXMzdkOpyWwFzbR3tMZJsWUPACKN9jfFk
PX0IECZ2BunZQ6VuCvPQzdUYakQCkLCN9lswocKK8V2+3ZKDSWovfrY9sf0nZi3T
ITtkL4GwyjDnCm4Jwa9pQc5x10tbO+5PN/3h//7m0Ho2e7wP4dzTmJkoA7mnSKSG
lc7fEcWZkQUylP11aWccsMQe9ID5XDk8U0166xY0dBkpJq73qDccAv8j0T8lqsce
dx4wpAz9mvubByHSc7UshxNRHfxU0UGIHZg5rx69HIlTuZlEOVa7n5mkZFnLcB/y
fFqDP/GzkL+W31lbBUC93XwUzrk5mEA+/jcWpnb5BvLHTRpSfVCqDUNluntI3liN
BcedIrvkRBV/ILx4z0eGbjyCd0PPYC3JUrVW6lNlc+HUmUOP9p5rQT7i2QO3SZxY
0l8TJQd7bEndzf+mfOhb6w==
`protect END_PROTECTED
