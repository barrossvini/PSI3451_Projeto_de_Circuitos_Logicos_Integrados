`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y1wYdmzE/SBSHChR8nZShAJSbl06qAxR9A2mpM6Zq0XeBVdsT9GB2ECdSlYgcsFJ
46WWaFdapL7dr8UCyNO9HKRPgCkpoeoOtfItKTMg/cxjRrI2WzilY3fO9N11cOEk
SRAOiVI/f9/bg45yfgrrnmnDzvQLvX3R/CgNHoP2t9YDQ4L1eHqT0iUH67NkwjHY
qHu7yUyhnuIkvMqIEtpKKsFJH38f76N/Fkze5EJqWT1lCFVTwnz2NO2IIDUfe2dL
HNo23LOyxcqqVLaNfS79EjubYfmGBGBAdzOIf9ExyOLQ+T4aXeRSmqUlyb8CO0nh
NDfldwJhJH2oVxwrA5eeVjxoV+WhUd08aeXHbq1Nk3GlMG9JYvK7r1xKCk07ZCPB
5nEvnFDjBv1izg/xCoEP706W9cYnj2R1LrPjJFWEsXOUfJr4o4/EDVYH5O6GE8JD
VfCfGMN3jXzhDxoZ9OTAXZsYmr+CIGFZfWaQiRrv8UXTqiFx+GrWc0As0JpVTQNy
ZDnThAtJixOHrq3X1elh9d52LYKdaFl3xEaLT6n0O46IseuQtNQAAHXfHCUPUBBD
/pcpoRA+OExGywbDjfRwK8shsg5bop7sDPeLgVwHkMJHZldSCa88mXb8ZWafikcO
0KuSVv8va4Wdjzr70RfC6lK7t6oiltaPCB8q+ExNmgirYK6UvXmwDpSrSVXwoZjY
aBB3CX3I8wP+Ks4Xp7akml1znBU3/iy7QkuYshN7upxosqeZSvGspI5Z8mljgAyo
pnT3kxOv23A3iAQo7FTf2i8yNJb1SQuLzfo/pEo8snQALeysNjZi/Otrjei14rhI
d6WwmBujIDPzgO+75NqVyAWZWBBZxqqW4vxf506B8opkeT9nTGmIVwnmMScnNOhY
XhAoSsdlGiAJBk+obV6k5TyPY80AxRyU5YbXbdUQpwF1SN0uGQUZHZky7SzlF4by
HvRRZNAj3atAQJQlb5oJF/hXt0tt7MzK491yS1euTk4bQiANIa6ZgjYAqwkPfcLp
6A4GoL8yvq2NjSVRfPP/RUCtxR40fDeRh+HA1UVA5n9SNf3rsB66uSs9xawgVY8e
g+/XwDxGJMGRuFkbY9vbAzurS+oK90+hLAa8g6b5piRwyA36LkdBeaf0iVinw3xb
vKGHrnj0xHREv8cxJGRG3E+P/JmPY0t3dUMnJevE5oim53zKpP72xtFk017wzaH0
jTbtIHoTdTJNtHSC3y7ncZCLegYSrnP6sONukRRiX1fuuz6cbSCP1A2cma05MVJt
`protect END_PROTECTED
