`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/GBehalY3GnZZvCZ7J9yW10B5E6lcr1J/2xQEzGENHBzZZFmjsCTRZUT1ZBAV2Ak
gYziGiv4kJNbgtiQjOKUvkANfQ3MakLCWjm22hojq11rBX5wyjhSB5upR6XAAwwb
r/yc0ztCTw901UH3ohIoSkWbRQ2x70WAAtvMINo0ZotT/3PyJaGlbozyO7fXqXWT
7HgB1PwNKU0NUJACQTj6pSYhq66TOSkGkJpYLN6sBy0RLOHXq9uzMF31wm1sM9h+
Q82fqDIbuOl0P2aiSl7s53P3pMKHBV504xqxgkLna0aVu/DYFU54pfiJAw42b46Z
ExPn9urENDELCpYKBIUjK8YLpHZW7LWt6adc0d+tDwY8ggIZw24HaiK+2kq0Lr5E
nsCruFBb694eRFtEzdrKZMbpwtZP+vl88g9Vca/s9xIXdOE1aFxqIuQ5zxG0kfys
C3rvEojG+RRWEas+U+YepPLeKyfWfl/tK+gs/b1MzlqEOWbYZ3NH95QHm4xyns/U
4eIszQNf8AuMM0TVeXnNf6RCRMK8DnylmDjc9dJgfdvqjgzPHHHTLbL6wMzKk8AD
qD/L7y0a1VLxLYGMq7zETDh84oBz60otV+poLjaMUzgHuo5c5sMRJfUlGInnnFif
c0MVfz4r6r3loMsSZJbdppFnBzHekPxMO71VNQh9r3PHpCMb/U6eRlZ/R459V6d7
48mBPyh/C6pxloYaMtdXBR8sQtFcI/AJCMogg9DhzQo=
`protect END_PROTECTED
