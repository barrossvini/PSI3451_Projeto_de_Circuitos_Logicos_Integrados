`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lMLmPzb0yOiBwYkhqv7t6GIHSYJx1MjirRXHaX2Ymdc8pASt34tU9q8z31vgTttw
uu/6nXn4LmBl/m/9iYrb2YgGTMCN6LfEKQbSTMUe5HBiFJjNS2191OUaoDbIPGrl
K6afYlNdVcvLILdVFvEyG7zkBaQ915d0vFo+WrEzSm1OfhqO+sOXh2KAR7dFDahG
PH3un1P4y8oxxzBi9/haZp6QflsnQNeZ1JVaMwYhFEWd4qVDeLHvQ5CkxSYS6IUv
v5aijlLRdgpnIzqG40wjG8VZ+S0CwXqDLHu4Xo2rx7RNVGTa6J9LPnX9WCbvzR+j
P57ADSpdu8gi5bzVwL0U+j+AcWaZLDGQ/PrZ39MLSG/qri7uMVePzxblM7Ef2W5/
+f7Xf4mBo/+LJRg4Ep8kh1VCnv/RztuOA2s5Mp4T2uHhy3FIK8LU2kzy8pl0gW6+
cWMbyAmIpQPwUY2MZ1monkg2N4n1ppAVjRtFaUMz4p/l5NnS4f60wkOs8Ss+hVBr
zLIKasMWem0SSEIRihF1+t75H861SlyGKuukwffcAowpPaknKW/LeiMdrmu0Qx5i
xfsM6gXgfZf6mOsBSrX9SRCV3XZIrcDXIqXAR+AGbIbfYuFCvla1zDwx8HV7P/Oq
y+flKFnM+0TNkjEewNq2NpmXcklGCTbtH9kyNyhDHREpOd01JJT8U52By/97AmL9
cOIfrSzkc3vTeDd4Dry5ySti1RlcXAKv2WftaNZbRTdynHumkKnSC9kLQwJJOKCb
OBB+Id5bINxIwm1WJrm1gQffZQ+rMBF0ivGqYCLs2xhOFo+JizWv29trqLnK8ZYy
PdwvDK/KSgN0Y3n2/xXNkPkP12MipLtF1/svg1kZMGXJ7apzyPbuU0BonpV0R/4k
aMNinmaQlFO01lBJwb+H4r7/vBcz7bfcOhCTXm2EHpZaBmmgoXhGl14Zr7AEZ3Bp
ZGRHyFiO88MGguXu/coTGiPQOk+es1xHOqZ2NEp23mAvLHY7uAadflxqRO8RASxw
9y61FKIkeR+Qf+LDWAQPEyw0RuQ2d1f9TgG5mlSyfURr/eCZn8mBw317uW37ApLG
BL+x6mJeeyUBLOE449Wy2htrNlyoq9oVFXwiqgo2/foyYA6Sp28QvDwzNwJfBVt8
xFzEn6KVdgtePGY3SaNtzGO3DhXR8VnNDYWpyF2ANdTHGo6dmGIFHliwmO2f0V9F
FeKkrLgfv0LcJ4J5SNf7uHsOjn6WrL/NZ8Sq2V3CD57spkAcVEA88a5s4T3yVrpT
3T696k9xdMMlEt71LyUyjEreLWCvqgQQsksYno3rkDtjlTg5DzAW7/lypADI7lz2
6Ok2Mq0fkBhBOmvATTwsAUw/LBTnBaVMsuCuoocRUrbPlkSEi/v3IyRqE7GKzYCf
SyY3HlWJMseKsfR1Cdwk/LWWeq/rtmKvf7ox5b8gUa2ZV0l9FQrYNqlLyA25F3gd
sLTrWptWSvu4biHpDnUaOyaPYmkKG6magVeYJSeH7iUpdVevGM1Nx0uKmztdoza6
fRe4XWHexkW4e8gzDeFV0FHHniUz/PNX4O43mhQjR9CwsauhVXo09Zz6tYQYps13
9mYiBjRTrrJvskBmkDzuY2q4lobd/Cb7N5KNgG8AW80S/jnqkpLAjHZnwGFOy9Oe
groXP+Y5qT1Ci2rIBefTu716Mg5U2wASqJpemz8wkvJe/9H9uZq73BHZIiOmsHYu
sRZvSPXmf2WTuEZgDO312MHQar9JHWy2jhCTjssgPvn88jRLfvxKiGoYSuLnmEeu
bHSrTui7UPtICP/2SerAHl9l38834DGArnwB/AquV9u1O1et10WgJ1U6+3LBw1U1
R8J9bdaYhmlW59sSjH8iyJQqp5x8HZ1P83pvXQTFn94zO+W+yAy7NB3LOGeoujBe
EC+vImuBd4sYQctC/0pryFJ4voIuyrygLCcACXz6IoBl73aetDfxaXjCQxsqEXMk
Yv7t2/bb/+WryrlSt7tSYIp1iqDblOTlFNvvw9JOyCnD0aEXfBcvFSOrIGUiqpch
fwlXe3G4yyoX52raGjYgCpkRvd4mKT38WV0skR6/MYe1efhJHBWI+/M+J9BTSoIy
ei0oHb7pW/LjlRWAyzlZK23nEI6zt3+nQhDs3SJ9m60hN4/JHNsvqWjLDrDIeXlr
aR3z9YIrphm5XMJLhvkZGuOZDQWlqkhiAUkdMU8VJ9luX+iKt4P8Qt/VEcap2YWD
G//CPuw0gtmnmoJXrtTglDXLF8bnJdcaLyreIhMnSXTV9nZbUFst8UIYxEsCxaGs
wQnkIYBtvfR3ymrYmAO4S/AEsk4zY5sF/t+q2JaCCHMbccTr4AbdnuvOgXkEBmwy
4papToPCeOh2eKKVPzBjNVMEuaBr52idAKBUt0QtjlqGxP6Uck69vwPll/DEuoHp
O8KpIW+IZgn0P+w6DfFOGy0umXtvxPDbUOyLkdbhtTSIk5/Jn1iVKDTCY4ZILrfo
vcXXLZZOSzmmnHxiu8Gb91sXxcTv/8ha0cOewMKJOWGKQtP2x+FL4dnzletMewN/
VHxWUL4G/j5lomPhtCA8ktPifxmKOXK0kHhLrduhMvqzu0oa4eGdPLWJPV6bwtsx
qU2A9BIgZKNTOJo80QJlEvxs2b21gQwInyKZazIPz7eqRZuInxgYmFywYuTdsUFM
eOaS8SGwMSamn4ySX18J5ASBiU9rbsONi7M/RADfVBJ6bC2h1VYh2se9iBLo5dsm
qFiUMiTPblunJ74lAVW11aV/SuUrJaO0dT6raoolvrz4cbUOF03JopmOrypDdD1y
WqCOdBXWlttQStAATWBAIPtK2B7es+qD5TTA0qaQRXPm/DX8nCwVmGNbIH1OTcf9
+tHzPSUK2TkNObeLxd9r9+5PYh8JemzV+q/NK20KwREL5lhC32gUmpXnnFfH2kPe
pZRiJ6akF29UB7aI61FlV1v9Qi1DaJPsWHC8fzptOW4FAZgl6sNsVh21HPE4JIwn
YuzSN6+5OB+zpnbHmn+wS9qv+RvpwLQrfFSxoNxhyQOKLO4R60VJfW/g64Ijye1/
PxuB9cqKnMygSKcX062DqP1VF5fNFcf20ZRfFVmfRpR48xR+NoVuFb9r8JzSwS8a
8MH6Ezj77+0sjJ3GQIE2pYoMToFLaVF8l7+STGhYTit+aFSseY/j66IFZRp/Hdhy
WeudtejKzlRw1VaM5OEfzf7L8LDWxpE3YtEE8RIpINX2aNLsRXg2jjfTk+B/qJ4V
RSAvVI8DAYi+DjWpSJWWoKtSTLyBtaFyA7ggvsWVxZySjRrZGa7kGabbJuFsDbgz
/ytAMuTQ5/VXfM5YJ1dy76ZyMSrAHHV9N4cPwNx4Z8P1ROUh1Ui5LFiuOZKeD2ak
zQ3bttE0qaZXZ0ti6BYbvpiAho4tisizVNPHfNJpVa1ejgGq71viqfS0Rhq5IkmA
nXF6uMCNPw0KP3Vjq5K5TRGFRRlxSeIccRRMWJAn9QYcDB8VbAllBDMo4GP0whjH
S+gLet+Z4JM0mtcSlDloIVB1ym5HVvogKtf1IZQpLUyWGgC5BVHt+P+kmaf0Xian
ZeGTXK44Y2DGGz6eI1HX9ySzDakVIa+8wLvFvZbUuXZUl/jRU312ySUDMDBi9xVr
mzl/5oY97b0URTgKqXUO77bIOaXIrhIu6JirYn/Y+li3H5WLHkC8kkI/c+338olW
RkSYoyHbzk1rUWpFSk85UkLNE0IvdXcpoXcEy+3aBZgQ4xFuME0oBA8xYL/rm6xg
YcwyGMrzma0GqhLBS/Fg64Rqpu6j+LIdCqZqDAUqhxLzSSQRzJRomCQo4lV7rwJE
Sj5Jcl61fgZMwB02wrPX6hlGpl0Q6p8Xc7nW1rR/YYh5dwjcveMETGeHg+VG3fxJ
LZsU5Wh2B1BSovNkV/GxzPR+2GrAEyBDCIA4ZK0HhdzShuA8wLU+B+1Hm/JPzO08
BPmbHanfOj4lHkAvRe0CneYySKZvcq+vxq6jvG7QD1VBpV/YW19B2Uw8qkoRLQY/
0BR46qD4KSY/yYrORITQTrWe+O2435PqdhabR+1+DTt5d5jfSwJJDgFU34CqWywi
wQl2CnyP8tsZOY7IEPQ5WsRD+Gx/YK9W7BV7aCv4oOIo2gJOOV18AAYm52CTUxY0
R4b2fFJOWecI9lsc9mnWLxhQZlug8pqHecLEEAnwv1uApoWtFiXulYUbka7WEbt0
pe8SCM0hXgQ9HLGsCPzvdrAXmCSi8z7bxS5ozT6kODy8QA2z3jhHD7p2Q2OSqTTs
RNG4cjb+mSFbYvRWW+LLCj/3JNBsaO25B4+DBw9NktKWaiIswzjUjJ7ANXYl2lb4
OvF3sjlnX1oTCeYF+6V3q8Lg/irAH0RY2+kxH1VZd5S2k8nnuC4yNVeV4WraPGo8
bI0Y2cMvNRZ96HoUKd1faLxCu5stZvHfVx2TY8WxdB6/GqoEFIC0V9gnFVUkJKHy
jXlJNFqT+sNREIuK1vD0tKR0vYuzQAQP1K6bDP+OVJzAE6FehBbG103IP82E3ykK
N1cKpsMaZ11+EgRc9brtVTsrDxHnNtoVh4hX4jOosBlXCR0Cl5GVh3bA/OMHqaUm
M+p3NdEa7GGoIldngTEMICtfSlwx3jWuReLn8rIoqUHUHqrYYrethbFnGQ08iLl5
UzIcoX3bJuKdlYFMRLKfD0H9iCIFYwMeAaseFIHCbaw1TDHTWjiRxc7eUSzx8I7N
0ztDUjTrJzKT9lDXXfzqAHEzV9UA9d3IUG70+89SqPy487gKkml0aK8AeeousQnC
HUlaIPdOxy/E+sbFGcXQlV5ZaMFoUDF4h56I9YWxs4EDIAcoozJgldo7i8bc6Zf1
SEX3HXEPxoo3JUvxR86f3zkZDiAb3zB1kJL/PN6KnUHF6V5uxQuBIMNk7mvBQBm5
pFYTowV93Pn8aYf4s4hdKhYsyZhcuPD6eLqFBE86KqTVGg4To0YcfjyYLcwMxDvi
+nLxfHmZNlQYPQ/jKcG67NKSAb4j+AJjT0T4TpmCqsWaR8c46jsIU3kt1LCSFCJ1
GpW8oVEJnSDb9w5LG2WScQPH562sqKH7axhCC8Bl6bVkr5xfK66LQhfSBfEBK8BC
P62HWMA5Q5+WMFhFCYXgZwjs5SFYFr0IWS/8TXow4rKHiFMzKJRvo6n3COl4WEFY
mZdkOQGzXlTqcWBpeW3PNzFNoNzJjuAbHW/fcs57snu2Sf79eXgD8BHWlHZ+W9id
SW/2+oyWK16q1VN5b4yXtGOlg83B5BVFuoPsAPfEWGyNDZobFaYoLrfq3oaVc78E
a1x/s2607CjtVwqlOIc4bHQkbBQXwiPW7rWEVrl4G2jxhjFf+LaXlXRbCi8DRvc2
0OeTtIw2dER2p0/FYVW9Rk/YAMk6od99xLNDjEy4SeOCus+Teh9/bWsLk99yuoj9
Zq0NxgYVyB+8kRm/aNZNYXO2mcjU7y3mTA9lyMANnzdhIu/dbnqgZLdFoVRPr3qz
rZY1/y01brUCD5/qt/ISZYSS8W/cAS3HjnNfjSvx9GRhTHmj08wDAtZqkdO4v4Hv
Z0IVop0/NmlUZolSrB3074bwkG7yJzghQ1Cj9l8voEKcGyZwot1KOYxQZGIQxrFh
v8glxfTbxzuU6TRHwv0QMMLBs4V199T6YEDeIwaTTVIr5ZOyVdrXp/PtneeXvbpe
Xoq8MC6JvedtLsiMPQVdoyC5OmpixeYP8Qc03RDHoO6TrAcxcGRBKypyrNVrSxn8
JcyGx9saU7/Ls3ZL8MJD1qqpwE+Fx0YFrzvU/BKWC5lSO4hiImAXdGAdHkFTNJSs
JyTVFqk6m4vNYU+LLybIIf5PiNhN11EiBx+4/lVaa0l3Fd7WH1rVOTdCv2vAwV3G
za5AVcZQI9rSuJMR2xbRJqm8db4vsm4aJUJsrmqH5QQ7PEmRmXadR+1ys0EKFuZt
o2nNUfjmWzDvEz3PTed6jMpC7MGbo1rzER8Zq5jbq0kSLcJ5WOdZvvSkUvWkRhKI
htRCEDImycj5ntmOsLKyt4vZlxivjwCHihXY2dSTu4N3scSWPVGLE3FxB/wvqOVN
hi6+4RVx9iVH2Wv3/TviO6jo3JyM8InhxdJUjNpuecZ5v3FWzQMc0dPfsvjM1ffb
Tzt6PSnG4fG6o1Uu6f5AoFBqe9aC50PIjeVN471epXCijGmmH7sJFVrMNfDsKROn
/hyXi/YOpGkodDjEJUFC1ZXJhMwIqiclYqQodJDt+AI7mr7WUobgdP9L0dKtRaHk
qE7RGoY91s0Vpv0wf2BYqa40Fu4SHOesAOGuwnRl9XlJ9wCDYjtOSlYMp/d9hRtL
OUmVztcWaBSVNtBgFFujHC3EC2NdrfvAmYe+5X6wVUaLtYm9noguiE2JAttMNq0g
58LUOZ+iQyvqjd3AkuJaDUwpm/mi/osuQr0cK4YiUmbY9hun2V6BMNg08WdbmQB4
wXOCXLRwTSwRqWHPjswaScbnq8cksytXui0LNra6leUZ4YVyHkWtxvogoMGLuuaQ
8+OwFatjRJL2dRs9VFEw5BUxUNE7zSqGUIUZ1lVKqAWvenFfm/gUN8bbj+o+zyrq
ytea0k5qAbKJqFh07BxZnPh6v3awNPdW2wf8nkzat3010Qhjj5edCekuI04p1bRB
qRHc9UYlPpzjA7Zmja9OeXpExT8+Z3H0XhuzUVA2E5JEK8UASkenf44wYH8uQRe/
eHR7AU/YVNKeJAnp1vd6gi+qkUn0RBZZ8r+kRuWZCf/3n0/X67ekL6CPKDpt9O9W
aTni5bMBnShj7bovSx2PEHC8GR9OJiJf5wh1whkkputXokAd9h2QjljBQPAxtExP
ZWvYCw9wruXJFDz5hRoJvI3rLNN8MZYQke4tguIPMdkoXuBmMaE8aagdqcnBQOel
p5lDdSlWTp4+i+Hx3Jc4d7oLmB3/g76Mc9FL5CcknCj0UuXnPIjRuZFxPIxBJDR8
3qS9xSl8LKP1xluk0aZZZBP8rFM5F1DvKC7OLqw0Em0hY9jHwfpFE7R5f8Zt53ob
J2Av4hhuXf4Q4Pp+bSVFbgAhgIRC5WUizeaWn6hRBqZlb0FP9HAXodgzxgDUtOpf
gyDkTMEExfYYqDV3U99uRyAw43UOeoEE8iEa6y15ZMKCl3NkMkeyJusrl3DHzMKd
CzYghxKTB0OC+kBR/vYbAIkKiY5qKB7ZmbpDDY3R5C7bOxaY6wL86IHVOkBEdZzT
j5yDTBrNnE5k5JHce6wifJXMP1/d8AHbRn00Ozx3MA3aa1QwIOn6aP0m71OG4osh
nM6O+WtvtOPc2RnhkqheRMmP+3cFL7lUziFUWQYrZrMEcl6bTfVJHfmTR9Bky6K7
e2tS3dflGUMNkqbkyyg9lPiCIkDH/UBM8adk8h66HQu+yFM5Jq6pAcd/dHUW7TeO
oX0CZsooqzk1axi5KppW4Aod0ys1Wjeoj2f6BjeDxokN3RXx7VrSCZGO6VjqLuhB
u1VLwfHdMviLq+B7zPW6k25sMO4doTbHB78fhCRyuc3HW/NnhqG5UGeDWzs7bI2z
yD2vs0NrndA5EhgWsabcTEuHsHiqPnwgH1jHdR74C0KLF9cNoGJIm+/GqR4YaRUr
TEz1f/JaCasr71p+FzzymQxLg0DZRkhQFYsP0qEH0AWnEeGDfROVOO3GMD7TJbdX
HAvwv/T/tAGJvTEf8oBR66v1E7QBLbDCpedWYKqQJjeqsIxTq9NFaZHrRCigs8UE
RWNu/EBW5YsSLvXiBXnaENKc0qyQsFzV6KtZNwkkh8f2uid4HNmHy55tMzUEgYpZ
okJrHFb8EjX19enVNYUwHDQwUCXZwSOL7NTbWBAgAMECtQrz3gZUPqAFISR9xeg7
Z08Wl45vMzpug0ScnYw8b6CAQeN9P17/PBTSK75e0K5pA1+7kidLadUb6qK1fKrp
dKscvakJh179/w+cpRNDJaa0LFq+RI1uD5jXpgAk7YZfHMjhWJqOwdvCs5XFGot0
ffVvyTPs+HB8HP+Elx/aEkyWNuEjVo3NGJj1TNYRnV/ZSXkXgtKReyozg0l44meV
Uqyw0+QHlZNVN0wxH2eLq55lgNbVFYxzW8/a6uIyA6V2/XjLUPh1iBHn1xQ7xmLU
B/iW9aH1339fmAPF+DmIerZk0gejmSZ9B7WP6HW8fST2npbDRjSpX8cVuFi7pyLf
/m19YEdr6/j3GdTLCvCq9Y8s/wxl4vxsHl4+6JvtO8H1fxpAk+RmznrKvN9BYcaJ
5qBYUhSQq5Fhc4Jc1p5mh1+noIZWJp/OqLKw+FNzLDzPwOUNR1SBZk8TB8wj06uG
TSnkrCtEEAOIRqjatYIu7ShSD5+4oFg2IhTi2scQXvkvZE6emfOZaxADTF7qhpOD
8AGOGOOsxgT8JeWePyIS75KAqA0qHmyIrqN7c4Uw05UVtnoCkxblbOWlpc2L8gtH
JUKWNJCYPTS6r6MzJgWU5plqDBUcSzNp4X47iAnZPGPTgy+A1XwlyCgg5FVSBOJb
xJfhnYTY8X6En0WQPBk0iCZTSHjViy1v45EKNMZpTVaUA4VWIgEjstukK/WDuFIB
mPMKWZwdN5G6UPFj0SAFSxvIKViyS+en9mwHRQ2drXLQ1Tp3eEztk/mf7iJIO2nK
pV6l46pngsAUpgaFmDyST/QuvdAdQjxc6BXR52U9Z8y5/PzZdW//aYMCP/V6GIX5
Mj/EnPTUoP4sAUIxJHhaWdoQ9DgSI6N8UKCFpmcee9kdJO/0C/RXyvNXcnufQgCh
v/a4eE/odrvK65oJOKJ595Nk0cFrKEn6j3sNp1p3De811hyYa3+IuVWYmuCRRBMY
Zsk5JXMT9BaS9IIQ2BAL1CE+gFoxUQ+5V5raSX8TxVvJuivhOlrhKiszLE5NapSS
+Jhx0IyljfptpbqqAlCzZW+gQj+50uINesoXnKs/ayRdXW/F+PugRqb2KPz/a9dK
BfoNE6IFHwdspGKTH+Zu1AYzcASrXhdf0OU3AIttll8/C6lYr/SFjh7498lSbm0b
Zq9PmKxKyZOziZ0Mkwo7cVZepSmhD8s+f9iuIygHKIYyJoSn+x8KaK9TLjmb8Za9
e3M7MScIRfxscNAIszWQHHq3s8o4UTUvZLlP7oQmNSL4uD1is75TskRIPw/eCEGc
Znlukr6AlkQ75fWiPI8WHE9zf3pgJd4Fl84ip2zfXa4srBJF0o+yStcZSTmWSVnG
ipvts8RAJ/POEB/YSH+dzccPCDC9U9mfA3kQBkwNW+UQKYlhHNL/237dSNs6SULM
D98KFaOGq3DUL5Rhdz1oKg7lCWiXUhOhL/IC2IYMxhfjjrEcCN70Vu9KaFxobAro
cOMOV4mODODJlBPyUO2p0ketb+d0EqAJgpJjn1PAzuAxmwVwXjrYy80MK9O+Mlga
bRyJvOqLJRIYYT0e7vnbYn9u+L81hIerSO+b3Krktf1sjLQYNT52SthaUU/BaIS4
yP1TaCuK7ml0qno3daopkgYvSodjYKk0RCgSyhTANwyKQet556KIsNt6f7buwvxI
xLhAZwFx/FeFOfkHfoij9rhpefr+dof2DzD/JUg/pMOhVNwqAJwLFYqFC/bgR3dK
LbByHpXivq/IWfapseEV4vLUYjXeUPeyrMZSPU2YCen77lXaYomDi3RM+GocD41r
yrbvHiuWHlRgcxaWC5iFV67nKlrKho1Sg5eVJJvlsHtAxB8mCExPasAXw0G8j1UV
pGKM5E8rC0tddNBsH2R9qVYjTVUV32gRlXEfmtBQ5/kU4gPGKSN0ySWPzHZXqRi2
c0dBzCgCFrgF8C879Jo6GeNqFaKli0ro9QYzT9iZkFBFxfyieTHJKUpyNcZ6TZ/F
ICrxkI6L3sloaxTGeGoxvmSobHprgiGzm9FRcJnDANChkXIAVUXQ7XeCNZ9Ndptj
ju8oUIRsb4nDe30EhCqV87mSL2XNN2B2u/qcRUIV9Ve5Xm0AIysgRcFrEN7Giv9H
6ctY8EdaHbUbYwDBRcHw5LPMpPLwCkqTTi7n50QE1Q09aiNO3THBO1ZuonKRoiUY
n/SerI+Nqzt4rQbf1Oh8DuzhQ/ZKVqVfeyHus77ZIjgfL5mEN25VG9UjjrtPPLNK
Pola3TYcf1gaxzUZQnVvNLWNCq3z0xpLcGveITWXE21LLynjBTIXcg9GVA72PNBj
KfGXNHqb3UQzBrvMF+vcJxKy88xNqE6vjeYLopknfX4MuTA2LUUgt9sMeb9h8FWx
MsnZgsrYtY7B1qrXJ6tg21Iq/1WnGXTvlhxvpPU3wSmsjFt/347Sl9/D0jNp6ury
5WfyQZy8sBrz3u8cQBLQqsZ8BWPifQTYXeI5j1I145q+7da7/ZEpFSfvrncGzuxN
D0dmdik2MnNzp6xq0k4jDXrrD1+zS3e6dZ172zVlvuYgfoitGGyyrrbjpg6ipW/j
40XoXa04J9RN5Eg7b8I3Wdz4MNYlzqAj2gn/A/cpCD4zclvTLrVUfR4MPLXF3zUm
4nIJ5uvqrD+f2jjLbqU5OV2i3puGsiMf75DyPIa+m2r3MFaziYpFWft2HQnvwBkg
e2HS2s1+bg8dIIxLPIoS7aWDI6gSjClz8WM4AOYpZfUSMSx2Uyx6JLsZ9c84SrA2
axz+9lCbaytOuWahRF/HpuVsokAr9ZW7ya93j1tdVsDtiulgvXXLA7BJEoJczVmQ
Oke6NdsJeQdlIVF2ZkAcunCDmLLjQXepcp+qF9xjKPmMkHd1rsA8r3THX8ThKkNa
QUlGOxbWf+W6oUJQU1lQaY3+/GIMYpuqHMvbOKZKS5w7JORm6Pc3h0BYKE3umPN9
gKxidsvg9oYRH/c4jkQwAlZBkoCU0uVNPVMNfm+BvtXEh8W2BTW9AgY98eoEsz1o
41Tldn399X6HdDAQt5hNGjrblG4pufNW2t6+6QrINyp2vke1byLoycUugZJB2zxy
Q8qcVacXq7pcz4bmEE3yK20EpMuE6KB3P+VJ5tUuja7I7F3Fc5fIHMOSAGAJp/xl
x8PpQABnnRNwxnvFPqGhjxxA6h7eaWHbzksc8ej1Ptif3EnzB/Xhz1ADdtSwBAVt
EBE+vyFSDilsyrFSzBPIJOqTLwk7NaeShsfWQfHRahwF6sklVMYdpXZlF4BKvsTq
4VW74Bd7utaxVfB65nVh57jKrsjPNjo4VpSCHiynirDDME+M3wARCcNzO4jOmQPe
rq/dIoBOgEiCRoggI3bTd1MZ9JzqO4WgYND7sjF98j1SMU0BpbbdyB2LTYWDwhwv
eiXrx4VQNIweamj85iLFUuMCnLcWIgguG9pnA8USfpkv1F60afVrFQNgGYrtzjsc
ZhbU31sFHUnrC1gtUfZQCQ5F2kSqxmfhOywvE2TlABd61WdbtsHBs44ZtZLYxWgf
PcYGpU/uLGQZyOHv8ZYQaSU6VCAAMdur6bbmsY6bmqvoLBRv21KqH6YJPlZrfKlJ
SwgDMgNt4rqWX/V2cZkPhYT6W6qZYdkN4pW0AgeXyZWBpTYE73PvAJCR4V3sKiLo
TNHE9Wc8qn6dJmC1qgOHugD/KF/3an29kGCkVxL1W5I5cXg16R4xm/TxvX9yCD2y
5tdj2dr59vrB5C9mTx8m6VW4HApiVrJV9w/W/uQ8NjdCcHDW9qI2uxFf9iELt9w8
2S9A/4eMwKE4qq235Ku3EdHu8/eizJtZiAEbJwQ2U3l4q1M11Qu8Ynj7/gP6YbFO
ORkOfIps95ygHrzMUzq8sW6QSUxClPJfDtEOi/Fcvn9eCMfcFqIXBWxDJTCPyQML
zncSfMIDPU4hpK73JdcUa8fcKZoGh4aviLC240ATJtZufySSblPzFAA9951xE1v+
6iAPHX74HD+GBjO/0wmS2CJMbbT8H/ayRlb4mPdaCSqkDK2t6x9wR/V0TX13YKVP
Zp9zWJR6K8gGewmdtkuRzh9sWmw+yyOuPyXvzjJCaysqT7+LIX6FPf90mFW9SguD
FxUwzaUd6IlEj06FtMJaaecdFf70PfUDowAsOFQNtnv84rzd9CUy0U1yUJ5hw9rF
TvB42AGB6efIVIMlZBTOX37hpnzHAXk5W+zMNFubtfWH7AiI/sL6/zlahkIbk+z6
WyAyW2Yp0uRGFPzn2PaBQec025y8bBNGfdpLefTcKQEUv1K2wvTcKAsRhH7XFUvJ
bFDLH+qeIrGf8eI8WmzzcB9KBejvvW0XDWecX8eHdJfXKvtS5UWOS+wHZEhqWe6X
APbQoiZIR17wddfveOlNty1Zd4VdpIjc6SxwDt9ATXUfc8s2mwuSXERTKVElO1Bp
avhI2OkkKGZRVNWmzF4E0beTgRCeFVGRb17POMamPiopKkeDrjXodrECR8H65pio
q/QzclHrishvxZvFMmHultnRO4y6Unpuw8Vf5/e+A4hpCLAt5bWsYsvToiDSOUwg
vX3dCvPRRp53r48+IP+z2KcMrTpi+Er/sE/4q0fW623Ck2j6fwiqclX7NxQkQDkO
pBcuT9l3n4jwqq4/vgHmwsUPZUYkLQ6iRMvxoddsM5gOX8GykbWveSzf1AYXva83
J6OKLHbLsP7Rt4jHDLBfoe1xE6e2526xGn0QVdflvMQiZ42MDZHuAXMnoNU0S6A5
R3R8qkpeRiN49gEJOB3ijbIUfSoZjbsKbG2m8CxdC5w0t3GL6gaf34QK2aoIkNn1
2CvgCZiT0TjmUMfp+l4u8g==
`protect END_PROTECTED
