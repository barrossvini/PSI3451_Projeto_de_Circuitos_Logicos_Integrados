`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkUyVk6vQMuXEGIBrD3DIfcw2wKoEeLUC/C5heJA60hwsxmSiJwkcCJpKHSyYjVp
Q9vuIpu+lBDsP5esv7b0g1Pf3CauuIaPv/grfVNrxZ58tbBJEgYFvUjqCtmUIAJi
ZhXm7VjYd4e5wNHU1VfJ2Hh4MXsvknf6DcfIT/3pOqPT0BVxutnAAh2XZkt+EGnz
aYRFu8ea/NIykcpFM2ek9aMET7SZcN7PcR2mh+GjMULkYZb9xPcyLXvFMtz/M9Nh
FW2l2SL+6yfmWbz4b/sS8zPAllL+KDGZvWBwM1oEveUzFA6QLVRCGxFZ3C1zSQJi
bzHrOltXkDl4ul9mfPbG1yMTCe5VJ1NnGN6ZsNt+t/kmToypsUbSkNIegH7LhMoC
IrGJV8H7vuGCtCy0809D1tHD3hapsKP+ZIqqTJmnsyV8WVMmqZ5fdBraX9KFt7J2
fTmrZkUpWOwjr6ZX3bBStO4p0Re7GoT6OVE4QvwMLW1+t6ECGjBUJdPpSLffv1Ji
8WcBws5hIKwdVugiEBj6QcpvFE3q2phFYKM+vSR7RPIYu3e/kmcyEFjouRh7KDUU
8jzvUeY5EAErr9ZTzY075/L6i/6fcXa91exQJrgrwzZIy33hRaBnqKd9pip3hgJv
6CbSG4KWTks4q6uv25uJr5ilY6+CSnWxyU5kCQgvoesqjCVa0011jGM6RqjCxn+N
8XL5VhfPu5QbzEzMgD4pIEKAQnQn1TybZDTN/Q0e23qQCaIFtlSJrOmKtvm3k2jW
o1AiX+g7u3JyWqkVuJowNn8hPvjy6gwkN4PRL/4JeFWdDw9UxtWEiv91vIGAGb5K
q/n7L6EgchMwmg3fNsd6gQIOcQlXzn8q/vh23DIwuqs=
`protect END_PROTECTED
