`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lOGSzX5Q/e2OZO4t2ZDRBcNzxJ5YkmECTHAoyYl/oshFbXJthqhSQ2tOFsZs3RFR
kRxRilefFn/splpvKZpvFGVjdZzTO1E0pVkceihgtJIMNSMGuRi3bXyZNm1jMRjj
vCU9VsPtMianGmJtqBgH1B/q0FXdUZbKLm4D78kuzZG+3ugCYlc9Z2z5sy2ds45v
tv9kvy5H7CpsvuSmDs9gGzer3gG3ZjtxD/Wuat5AmOuJgLKqDv0tDRdct1xA46nA
tsI5qAb7JRgCrw4B1JXfvSElo9eEEjsZ96+IQwLYJ0ugDWZsAoy5Dxo0H+fm1p45
3uuRyyzLCyIvIrvZpMZpbJpQr36UdZzVORJXQfeN9xeeXwhbHbJ/BL2QxwYjFk09
g/f+vfKobapYYqd8OchmsF4XMOP4WQfA1Njd65+yqY0Z52CDYhHMMfncQpVzIvVQ
97++iJieO/mDIXdTe2rBtdTpoMbDK1V7nPTvUGLEprWTfuCF5mhCT+JsCJcz+bl+
qLmuiIXXEhx401XP+C+IFLL4EAp55v30Ju3edE1NqWRYhAPsfcaHritu5fOpSiyd
uFhEGk4p6kboPXzjK2XOWXgsVEwQeotQOcCBS1NlRorFme+sFt1TvmDVhK/VV9/7
5ABLxwWXufcq/B4s5EC0qqBvSYx6YPhx6Jqv1GCfRsT2hF4AM8dy+dZtexitzbYx
wLePfK8A0MlKFQ3CetzCCMm8X5hbKDUrqKrIF7/ks/6Mr1vOdS5JJfAqYUSEIRU3
3LnqaypmBjNkkBrZqluXgcwCywhEFW2IWokiQ4cX8O1CRDmEGnELihAlOlLhEnPr
oo5XrYKiH4BFVVmUwzr8fgPtN56SM/3FJ1iVtqXQQL7w1kuMDxZJKoVp5q4SSnVq
8Z2gO82hz92nihLJCa434NK+CN9qItxnu8+rRf9rgo4pGbMglCwOX/syult1xt48
XI31UbhsSHbO7n1K0OiojIvte+qwmP7/9rqYdRJgfZiBV4PoIxBr/55ETSKrzQDc
4hxDd10pDA0ddrsY8n8OVwFEBNi3bkEZnTf7wlPlj49WZx9BTVORTlwnp7t/6NME
XHhuW2LosjGJ1nyyZkz1rlG+HJY2StnjvbpU6MI+VxMHEJ+aRbs6b5B8zhgO3UCc
3PWBFUtoe5n7QahyGSfzH0Ts42avW97jCIe6TH6MYL8p0Vv22iukJP6uud3GI8pR
Oj5SVC3zKNc/lF6/LgoXQgA/7IS4i9KJGhe4nJSedJswwTmENmtisAX09FRktY6C
qsqq/6rPCkMyDchT/OE7emquUcvt8UTeGhyxLmzPT7AV4PZx+NysoISPJtB3pRdp
B34K3w95xWQPwqzazkghZTlSbnyhh6Rfzr9AV/lYiWPzhCRqqACAaAFHSLNfwHgP
nOWZICZugZdfJNjltypjnwKeTJasniDp95kr4LgRw8CMaVfPsuq0v3vTNqDFWboT
cf7Do9eG4Ppe6mYrJfIMB+EcGelvAS03ZNeH+4Q4oSg/siN3rTTtpl2Aj8n54X3n
AmHo0L8L+VqIZDLjUtVppqwyREWBEzqJXk4/3Ym9FfEzz58ofkDgboHRwZcpCNwP
8zKcxM5uvDJikaGScNuLIwVDnz4hcZ9jMkPGrYbc7qiQCn+64yjwiOmRG3ConmAU
Q8PPhg51PHl+ukOkL4wB2yZh8JxwgSbQIQ5sATXydRCa7xsBxm+CI/G4DyHFG8XU
zDn4UrF6YrJHRIb9/mYovcmlj7pCqMhNwdpunuuvt15rmghmxaeOneDO0RGIKoom
6UqaCVqt1KAWxTnShUswvygXnE4Tj7eBAFtlXy42YNdy44dXCch01c6TMk4YQ3oa
ptKwZoIc/234ojg/qixNxfzY3tRdly8Rs+9T+LflFOw/2Z7YNwpzWaOCirXVqCa/
/Sorzh+ICF5EgHYvLKXfvXOZWlOkmS0ycwnljemYZgfRUolzw0RHPMppYr4rZZaY
x74+xw3epTQCNKm8Ffibn2xGApQDk9/58UuTVRfwlMbssI/jPt9UF5Sf+WeFZo8d
MIoJCCIaQ0JR8Tx5yWMvIzDbtr2UbK4A7zw9aKhTKV5HjJ1YQQq2doq6x1VdEyer
KJoBfGljT+RLdDQtA2lxaUCmBWrxf1xNspfIENZY20df088l4S0S5e+75oxmSuNz
RmmGgdv4bzPn/Bzat/3UXcUZZBElZHX8cM83PXHtEAhUSNpBMTyT2msX1KaI0Y5f
XhfZaFn/UzXOjoqdRlliB6zCPzGas0k+60T2/U05jYu2+pY+8irUaH3varqNEfaz
COhWbOpa0e9Y16XqEzn8NEiiQ1dAUsSHqVvZftoJWWtzqVyRnPAl2OkRjAexMvaN
8L9c6V+3ud1kWq0Hu9ERZJn4Yo7ZbY/49vO49W0nfzpFUAak8/cYfRqxycahSzAe
eQrvMMuntbaiyoPd/+cbS2t3w9laLf3HJ937jAw7YYfQPmjry/h07nUJjUhUbnEu
mZKdRtJoFdzElM0sjwPbRs0isMIxGALOp0OIPaSiVz5lgnyrjaR1zH/yn7FlEyIe
XPEzy1ciRMQo6jNs1QAU7xAycraOM/I/cYukYMOvdG/GzPwv774LI1e8T72HBCw1
ifW5GEC/syAMe5VFJlw6fvPNCVDfWNAQv6CMQ1Pb+55CCX3TM8rvDFOjgIy08tzg
8l8r9xKgtOViGowmOftoNGmfrWutbCiBQ/BPjWzm5SNpzKr7dOVHmeTJc9q+Qovs
dlegE/Qdtl0ZEI0gCnVNvdTiqkGh8+ZosI+6m7Rr6PbiEwgqnOUnU21t8WKyu3Yh
6H2b8xf6UsN8YJEKQJwE8SQ8eS71L00/+1T6lSHplZPgNSVngrGYY9ZFZaLTJ8hJ
N+nJO/AYcKyIWDU1edKoRZATCXF4HD6BAFshaBMF466dQy7HAp1gLd9PpGx26SB3
rGMhFIpQMh1T68P/w4a51At/fm0klHNRyDvM3lfrBfm0MxKF3nbUbJOzOdUjh1Xm
d1JSd2yJ+bmmSd4ECmOOcFxcrF2cfHldtUazVyqKIbl1rWgbDkEuNjMLdIDTSFdn
Dhahy0TL2rgs29C6GBESG5yubhbSq3g4+OgmVN6TZCUZR7wFzwmT7Y5g0ntsg7VB
cu5nLLzXKaBv1LaiGzosH5lMZXfZ3hUyW8Yja9/aUFj/Q348pe0zeFw0R5l1268w
nZDMwRn2Jm37x3ofi9WKEpk1wN2TCxQg439cQxjX5ZwUiUHRWwbR09nme7hZBtPu
htNkUxhnJCGopsemPOlRuHkCDU8Z7gBnouJFJhnbFkzL88QlTNr0N0Kb0wTWLLpH
QzgsbLAKuKSsX4KvQ7AWcjCw9n9g8zVL+9sVKlS58QM2WslneTjrgBbQGCA5PoLr
7yI+1S4ZAI2oKlV7S5Ly0HMqHQ0r4gQ4qxre+zvWarrLrpUzmJyapydTp6z2sqB/
rq2Mg/N9Z0ybflvEzbkjD3J+W/GpzbEE16YR1SBruIcHfPd8vxpkUODPlZzzPwL/
4nD6Ww0SyZGAz69+v4Cnyh5/Dnpf7l9Fkgl9ULHpz0Rl9jK/DLQRkYRgeP3FMNdU
rKd7U8ZeHuGiDciD/trpfnbu16WR8V42xn3DcHeCA8N/Gto/qmeqCWmFjRjfexDV
gmuaJgJZ2tNxqrUilL8ERthRVMnz0TqqxFOaviGXv0sdAXr1aIAo1bOilXO8HEqB
wgh0Zlm0oY6W24gN87/0WgCPif8xtoWF9heVh0QEEHiI3dDS/LwjeYPBYhnsKDqL
FrmX4VA8GyHUWjviQLVdW9CA2F4BLkoqJyQWVpvdHyMo3J1TlNEblfpjCkTsiFzX
oaHmEuDyMqWNuumNAENqFnBN6hUqYFxFKwBMxyN1vCKjTE2kmFgv+AcYmJnm6zMg
SoVn+iyzu9gDEuoDeLfSRyDFR6Ov13ynC95KhzVAvlybKZkTAJQEUkiqySGQj0JR
CBWj9VhQVkIeONH4gVVSKYP4TTOaZdmDDVeXvmw0s9LJIgl+aOho16QIE2YRolGZ
rV+FiALF4EAbPy0PgO0ugQhz0WlZg/4t1iDJS9ZPAzdxHnKJ1uiatD+TKLiGIsRb
z2gahvvCbO9iahXC6LiKxgeHvUaR6YhAILn8+AJpZueK8vfm81XU+6T5REQcAkoh
JW3DmHXLv2uL3XdVO5c7Hb6aKd91mu8lIGSGQGEB354xJqFHax2Oo35yRuzqIj0n
h4TvSrJlFI72ALdxnRkfmC77LPB6CpWof//i66iMDIvFuBpylaSohfrb9DtfVCsr
yLMOmZUH5W0LX9jGBx3X18Yjk85+DVdMq8FC/vWoURhgMvsDAf8QjLxPn8P9gmxe
Q9QuBEsaBQDbpyYeDnAShdYvKNwWfHxPitzKnreB/8ev3QfEqLLI0xBXgkfu11LL
ucwdGtOFkL+l5pPhYGzC+kf7VeX4riDzjltyQdzcPGf5rzsP+PeNcsIIvUD+tTDw
thSpcvOOeWcM2m2gG4ZsSL0KE+8xJ//2CAu/4Wk/LLZMJut3Sk1XCRGbiFusLEHf
KSq7LJOMrHH1j7sR9w8du9n6yvAQNt3BgCdxGaVIYvVYjge7g7EoCNI7BD+Q4Fqh
qTNEr3dz45N2CbDCJRd1WY0kJIy9eEj85bLOQp4T6LkJxNWKIJ32HD1xfqfhjCrS
63ttfx47M3baSlVDJMw7ECVgItOPsr8lboGDnjjQ/byaD+spuZHzfrIzN17CxjYE
ta8x3ijZ+dRO2dOJoxn8JJZNAdlmk9RvNXg8Pp44mSO7CbFADGfnZHFoNdyo+4R4
2TsvP15jIj9TMn/HJFYeaMD+Rd2SWJy8k0d3BLoFbVFaGz1wR2ko0bxhXO9SfV/5
tavM8alz3fcvAuCNr9UAjmwseQR9dR2Zar5gad3ivST0rro8rioUnzoqVPzZ+fZI
qAR9WrNBjM9ft/AZmESEYSTmhJoCwFWtr3J2b9iRi1Tv5BtU9ylgLJkO4rXfQYY0
WiiEATroaCxJ8PYo2C5UUXsnl/KG7nFF7vnIJtXCoYO/YInnrm5lGFw2OD6F91fH
TTorUGI3g8dgZKUhbb+Go5uPfkbGPsMLLHNv4znBpPhhkx4awyJlYPmBpWdsstXV
Y56zoh/y963Ued60DNahIXL8sd4IPBl9qPwiA9FYEMl5LGtJ8yCSM22nbQgw3YkQ
dtJsKbdT6TZxirbQSeSYICinYDs914ODZSefNO1OrYWlkxK/KrQ8GhP4R9m8V0SL
ra0O5NHiY4Vmg/Nk+khjSRN7H+p4BbtS+m15mF2HvJcInrPTAXC+JEObKvd3vfZP
PGKbyDkBUC8ZiUMSGGWAdObmZnQrM/VmWTqV7Nel1lhnbQqfYNxy/To5CmxwSAt7
kpBZGwmfOb0A6AFFOXszHoPB4xw4fweuJ2qeYeWUPUll6xm6DyalPhZ+47b2FWGb
LY+VsxqBhr9VII/3gNPClSXkYKPChBB+7fqjLyboDVrA+1E3lcOFs84jrBcfMB4V
5j5BFN12IEPDHg5fs0DaWDMKj4qSdDGi5AkEx7j8gbK2ItAWG/BkEFXd2IBaSMyj
bhI8b24LxnqZT0Syiuvy1f5f4yzX/7dWaQBjj0GLxELWuu0K9QMYkFnFCGcU+Q4V
YMMwAkEVz+Dy3awOPFKhekJaij/HtpiEMxrbysAFl7B15PSahuOfITU2ff1Yyl+8
vsnU5L8Mx0N6g1RaPfjlI+zMs96bDp8ZdsyuA01Pu0LMmFcpdwahAD4AuamOjhRu
MU+JWk7OnWtcbiTJE7hnEXoqs+gPQr8B2x7zYC3YM4pfAF5zQIqJPzBG3SCDc3a8
6mzHHlXRQN7ID71VoyGEnrW3WtXcVmi+2R7nDOcie+9qI/99Q86xz5RLWNjKw/qm
DLSMJMeGby/XgmSsVfyIUygediGMRiLx6hOdVx8yiQIbwV6W+qWHxQIaUwdj2u16
AO0UPnhK746Thexpkjp07NUG/WVIq3jlWnK7/WEmzhPUdBUwFUl9R3M1M25zEbRP
gQCiu3rgBWRTu57NS0/N8cvrK+JENgJ9nUrGcG+dnHre4RZ1dQ7Iujm35rVxnnQy
3ayADNEWV0nfH/wbY11ekjrwnPE0M0L82opXqji19hiRhHBO6f4HM6aF+jvYAY3a
cI9Q4HGLUgv0Wq8xg01ieg==
`protect END_PROTECTED
