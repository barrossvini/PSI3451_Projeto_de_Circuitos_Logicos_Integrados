`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHTQrGUqQ3K0vl2XJ8cSZmmj0wcVwzADO3ptdwu7bZDEk2YdJXklRcdeKQf9ogE2
Jx3GxIGQrTSFHORlnoGvgbjmtAFSOHZy9/FMmPi4zePb7xDRJDbHtlFheYqPc2A7
Trv5G0Ejsg+6ZalBYzCepBXUpRE4LTrv7MEv4lFpv8ps70wjYqFYJSHlZimDGYek
ISAjXbppopodQHc/P/deV7CdYeh4UQ8dlnATlgNCKGqBvljJJ033Nwku1MHhrUbQ
F16cRsnoE5aBE7WOCDXkJxxu37B0JDKyGlK/pEepvqjfidDmDr4rk+Ag0THgPm/b
PNXQZrby6A1LtYs7FmiRlm7G8vaBOv2WvZcKesAULvk9Yq+eQ+qK822J+wYW2TOY
vFBIy5mkDSMs7puAFN4GjyG7SceSpx3sAcOztsE2GKTPkw/CdFJefpsqwvd62LR4
R/dsEoWlBAlmmRDtLd8sdOzYjhQjlefHVZdNO8tdlxOJX6mIaASEoTxWIl/F4Vyh
ui+uz/XkU04/J7fXv0l1+rhfc63CMUTuDEW97pUj/qG7rl+Bt37UB00qLE3GiftO
QSM04CH8oFgVFKiG7tpS/RVBIIScdyHdAeSXXf4WFF13MyhDRKrBOhEOaWY+R+Ky
XsGfgrMSZNH23vSVA4S4IIdz2qPFwFWViYchByQqB3Jev70pG8Hnkhe/ggZKhiXT
+Ha8J6VJNRtspf1qpEVlbie3dyrgEYte1dUK3ny/GB64AwCeKvJygexI+5VA1Boz
Q69cAaJIQp94UP14KIw6+VhlYbUY0myCiCcon/coLfW4ov752dhhiJ50051wALSu
QqQhRTh9ExGddw8qM/pn38xbFC4ZjfFE4xb2t9RmFiwPj8of84aucoWUxOvAyvjS
d1s+93PvfJdsyLhRWD+wBs/nGlMUTkERvxubT573gVwtcixW5RL/6iP2oCP4+yqG
VwgxNahFu8uxNCWCGWNs6Ek3j7DsfwcsjqqaGSpzWmvF8B8QPcdImHzuBX/jT68M
RQZOFNCMzGYzcKTMxp934XInzk8TSn3IG2+N16c/l8uh6JeWSZ+QkNFizFxGpBz0
l2aaDDR8lCzJ4pVzgjKrd0lDAQ6N+E1iStt4e8oan2E+og/biQ6kYA9Su4IIN8xh
XZTh5lFBTjl9FdZY3sZqz5yoT9y3yo4LeR0K8CRzGHfMqSo16nPhIYIMMafGDep0
uLDOondzH8aQertCkRisGLDOS/uOr8/G37+YtPYp9F+3smPHxw/DlTP4yEKwA7Tx
+7iXdlnHPiXlQqaq7YQosyV2YHpo9wc3/5UW4Mojat12cD0RCq3C/rZE+hBlZQvq
Hgp+Asd7D2QBr7ge1v1YJZhUxTfV6/aW3pg3fy9o6e6OcPsKfmeewv54GqV7pGkH
jzTtzYv2EhMGDlvP5rQn7MZodYxHHVD53cKuBr9lUZNIkKIYcwi0rqOPpDtRhTqS
q9Iego7g3v1y0T1cIlmm6sjFqOC8I/eEOSFWOUctbkyyBDj3llNmQ/7KEuIzSIFK
x7Di7z4mVejwRqPzAsZcVMDtkaRXxzpMhivnaF/KPcX2aqEORph2V5bKlKeiHQIQ
8kmP4FuOZpS8B37GT9e1ORXCWtFSVc8ls/uoF9jsw//25ZifiF0oqX/+1R4qA4Jd
jzf47prJwjd62qm693uEoZh0SudcHxm/w00WRxAZzkDIYjXo/GUSIZt4uphptOzm
/scmQZPJ7slK7DXkUO7f9A0iKfeZHcKUSD74VQnH24O+Ak0vCWdC+jDJBWKtnuca
`protect END_PROTECTED
