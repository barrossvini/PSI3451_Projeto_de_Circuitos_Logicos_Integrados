`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jMlX/7aAuu6TY7UrXdOn1cHs26+PzQF0jg5DAarVmnCrBzERLqA/Uhi7cGh8d1pI
zjD/iDQFRohCjfkWepX93wQ31upxH4kJgcSN5MDBAjyxfoNaku58VRyN/ERYu7yF
jiTWhJC9evWaTp+De/SMCLf5skV0h61Tp/HxDa6FtX7nL9PIB/vlFq5JlJFAAq0s
LSMZdpgqhdrDgV4hS/GUuq2SIfVx9Fj7Cl/SMRnjUeutcuoe53egpPulwk5yzVxU
a2wut42qg8WCKb6O1Qfg3CuXvuyDi2SwBfP/nSpYJ7RyusbrSmV65avBpprlv21f
repieLakbViMIltx45mwsTv43LBickS3DcQxDBs9Je2UHuSgepqX+1wMbPswewMj
amszVEp2dKlxYcuy0rd3POnA2EeazI2BnN7TeVDpr2c94hIXtYgEX+GxVJ4FIBJ9
pcJKW4XyzjOCNLf0YDVcaI5N6bcHFTnc8+Qr1jRAfhiE5JI6O+uUc7+/MjJJiXKl
6BZwAcufOIoVvNIypJANRz1Rqc952bhjbYXamnyty4ggXJk5+3wfvjg3JNn/91fs
mUUpnkleZUb5fTNd6mVEJ1M1R/80uo6+xGt4qVmSqwdk6nvfdReKy/lNObLsoAuG
VbRuuB62qPVKxd7JcDakZwqdifvES+DH+lZuViGmu6p1cwOyB56oXTK41ECKbFOs
Gaak5dJfad+5YprJgXB1tveSb+ManraP6dDfGB2QSvkh5VJEpgNd7hYbHQ8jB3TX
XkMPo1HHQ+RPUe04cjBpqwSU/VDi0e5n7JWOjVM9YPkYwjZsveTZG61eZg9AdHJa
7D8TbQhsXvqhh/1lASPCMjXa3ORoAfpBMs6MHY7puOD8fQw+cT2GxSeaTGx6PeGi
BiMfEA4Qoi9ruMkFAQQ5suSYAX+I2L0Q3v3l+VPlF83uUa4aol/M4v/Pv294aGSK
9Xwyq2bKWgL+DW2RDM3TEINrfbQxczFvV3cIpqsMuokhr+gf/Wawn+SRRRK5HFHd
ogSriT8PT0GNGrXuSEuCGKS33hZQ+23pW98ZkyT+yJsgP0Evk6xFLlOPjlXXkQt8
HknFZykJVZgLRP1R7TjJ4+d1mMsgfLYbUVqz2MpUIMpVrqvNAvufCo517qcKLTSt
18gnVGBsnReLlBtbQzrMSg==
`protect END_PROTECTED
