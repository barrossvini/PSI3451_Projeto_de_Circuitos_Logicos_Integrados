`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G0wHDiOT5ye8Z5i21I6fWO3CP2j0OVp7OKVw58pXWWxyxWtUTuVbMnptOJg5wbmo
XlY0lzq7Ey+KKcgNMM5fexZhu8eH2d6M7ZRqEq5T+MkGSx7sfRPaUB2z6yyHpkUi
Lav2c/YaReDXfK1grGb+AZNECbn+SqxS+n+U/ZiizHz/opc6eRxIdrvBC57onHLi
Nxla7KeghoIU2quQliszchESjT3vf/5wXQwYlyzQ62Zi7pyao+EyZGm9YjJ6Zn4M
QFB2etsIIWHNaIDMmGaY7fUC4bFOgtg0HxgYA4k0ulUranJ7LSuWutGFYTyIztgW
M8KnECxH1O8EtNk3T40yYRoUqB9X+2BYVQFs5VzWNQmGgLTrLLqtZHqitHtnj/+L
c52LDSaPb04a66cBBfzvPypJJCWOUpFDm95zW+beFzVyNmRcxtlfScmrTLmN0MHR
VDSyCyhc/Pij6J4821YxHY77Z4sZnqF5awbv1MPbupxzALsmkhu2/OSm+VeHM+MT
ypW7SzqvESMVKzB0jpoijFvbRqjeq7cimTmdjiFlnqaDeFrCcq8GedRfZh6GZJiC
3fTAb6BiB6/YLXiJjPrmbToWxpUgoJa6e7TMJRNu6CueCD/0zoyvd3SLFxr+GRwd
LFYf71geJMv1X81CT69KJZ8CQRUYHGaF4mV3SQBIKzWhWUePo1YaqWidIovyh0fL
9gsVXSPF7oJb36OkbDjf0ABBNgDZMWmdrH+EMOHCgC9zg9LXF6OhORTk29AjJfSV
LFmYW63k2vj9/tMuTA3p7UwJ2KiRFaZMNPJkA/0nxmSSRit+omOvj+pAp4oRsq/Q
c37tvIrl8RAgAq7yJNYO+PUZRt8BeNBpDUb9A7u+BdK612tilzJCYmy1LQlyjuj0
AK+WQFqkApL5soDd3Jqqiqn3xe2P1wDXVVPoRieyHa9idTn8S5gTWpRBlQ9Z16/e
/6dM9bmTKmh5PWHQAAVwJTvOzfOLbxFQrJSLFf0MqPBBfn2X78IjkVxi5kkgjxTn
FdyNB5+Uk8Xfy2WI4RBrN2DoL1B44s24FZoSrMNd9fV4a0GXRfKGw7Pu+56wml8U
d+jUnixyTWbcxsCAwpGHddWCgmgFlutliMMYyoh2F4Jqg08ylPfuvh+BtVVVcY36
CJd8ZpRlnxqBWxOTHXy+hVD27hLSdb1DvjE2kirmcq2eOZ4iR1oGX98JwCxOgkBS
jRVlx25fCAQFlDrTIqvDkaE5axZBRG/ga6rXuoie/E6f/MKG0Am/li0ACYVFUEYs
82/+su6PGBF5E4MIY0ZFNcKEweKd69GxYl19rIosKQo3qgi90YinjzQuHbXnYotN
2SaFkXOxTIW2JPu1InboNixWuyLNZC48uuPxsXX81RJz93J68Mdi1iuluO9Kp3lU
AYJ7UBNCPDn04P4xLcj6OyQOjvOCvXuoOlMkg6MBUUNi+NCd7CSN1pueKoKG8MwD
EjYm+p/ZApvIeeF+8QdSbKlxgOj337NqhRwxZ7lofJhWhgn3mVIzUmdinli2zTNZ
yvyWZ1DH0Ac2qqXH2j7IzmsAixz9OUtggqQyrxfOt/FSFoAqZSEB/0miUX4vsyCv
KSV8aP8n04svzdA1tYL542YN8FV0kUDr0dqkuEAHmecxbmKRlOb+FLmsjYlcVdHL
M0VR4xiyJydxuCWIR7ExaoLs/wCe6IvoMj6M3gPX3tpYB8MX8RYDedCsn1vQmrKc
wwbE1NOGyo4O14RncXnKMImZUchBjKqLWBQz6Sim992aBNlcB8pi6lMkVGsLDgz4
cUUA7bi1NckPyfHLdwk8JuTXhL2hpFCYLuk1/C582DzOsyB9U1rRlYttbE46yD7E
UdlB7fZUgG8Et5Ir6MDRT7MFhUS7kfW87IX0NfWjMYEZlDOKTf8/Yb7hXP/+r6kU
wExJqt34dW8xKdbNzaBgv4NmMBj/+TFo1obpS+JN3ZyaTN3jjdzyvTTVYVr4FM8n
DzQbpWlJdXvWBEdeCZfHJl7mnLRvhedDySBItwpmSFxMaxpsBldAokr45c4wLMUI
ggViI8IOjUjaeyufv9wbbp0YbJme3Zj+xAoFA5upSSQFTvdGThU9u2497wcGiSda
bksGOMo9zMDIRqvMTTxHBRbwe+RrsHzqT/zmz1KXwU8eFiGx1B0Fz/sNW+fWbHKe
zwAn2RC0vemeghHXKl85j0enalLbeRWDRv67cyqrjwPz3h0ktYHg38cP2xizpB2Q
Z+1HcOU1ZMhaQSMDcZUPoQBBSI95JyuPDOmjRm4ba5hYKcn0T+aZiyIs1yln+KpM
KArLwCNyDO0BLpwrfzBFa7E4hN5cMZ/oIfWsioGVyVeNq2uQhJJ6gLaKqag4bDZ6
sCU/PC1NmTtgblZVu1zRsoInK3eNPGPE9tnmO5bZwXEp8238wCu7TYUoYoxkXS5n
vgNwS1LjFAdNRLAX30ueBIAmt+du1ggJR5hFh0oYKfMBsNzm5YmisW7q4NXku6pK
0vsSuWQE2DGcM93wAjNEyeFC/o2hBrC8QlPQcOsmv6/zwphrjlfItG+B+tHS/pIL
0HR1dDvyFFXFT25SCDxS+SAg5VZc50ILRXo2zw7SJXh4fjPUEvo1kg7PoTyQc9h/
2RLW4Ta+GAzRNpnxUg7arkf17v58f+ysuzLUz7i2Tjjzuxv77csBq4+ykF2i1mDc
amZ3N4SZjS3QKjIxRN9J4c8hS0nct8Hxqn/y5F5KSjoV+YEvttNCQJtVC69ulrYR
eeafhE08GuX3ZZVu+emT2UWUTwwxU4Qg9+XykkpsGAzAQQ7LSpxBtPQ/SY+MVgrc
nAEGmM34GBqUdlCTdxXmFana8xdYhfUpAYIi6ue0S8DAVp/xOjYd2tkptMNHdGW8
3X7DQlN9LFmOkpNehwdDKF0EYhYdKd+G4gwQdRx6EyZzZHmzWs9NsG+tWu8qjwiY
V/MpAJZmB+pizlPuoh6NQr5mRCBHvVZ2stIIiZPi8Xmsy8DbDUmttrrx9JYiZ5PB
qlNYWVM/9iEx9z/kKi2KNQgE7jqG7FMzf9UKiRWpgupYs72z8Mg5ZABLrxFbvVE5
p89XK98J4yCDHCAXj1ThvARHwGyO4tGOuD0EQ6CfmXHLPBY2zR8zaXdeYJm3+oQa
xKab5XzUhJiyRLOVhcJLqnBSAAsAQ0W9mLsX3kLp+vnoVVdChxwCpkM3Z0Y9ogW2
5NeWJa5/GWg7FqLD6a8/gqKxmQGbKVKBdeM6RJQSAC9WKBrI3goHIVALAOA3BMfP
ES+sqaeq1DEoJZ+HyGuFOIuzspdNDKDNM18ZmNWC3wNfiXpKxqtC7mVqDODJPV8O
w1OLGU2hq+7L/TpJJBFI0joWnTtWImhZHmZztX2pqsqUErVpzPXC+vO37jd8eW0h
YjQIUlzEo/RzrOabvq7XLwKJlXc+wq22j+7BvNFXvINH7XH/v0MIh4wWRUPUJox0
8XRrZ4e7HCG3EmYOEeBSePI8a4MOI96JfpPDjCvCdswrbDiQOhf1Ce/xJ4FTVi1s
HkEw2jP4tBjNSiKi1dqKh5U+aue1my3nych6fuylV5dQwXLsDKF8+jancQdB48oG
ZXRN268yOctLvsD8grXsFON3Sq+LXBNpn3eevjcsad9HjEHmaJLMGCt6HqRcONNa
rmcreg3S4Xvdlowt47Q4eRRaHqZXGTrAIwzJf3M7DI7JcxMaCVYeL99j+8DpPc48
UcVBWuw1LZvAFOa3DQ+zwv59bIA2kUo/mg2XIn0GoG89QXBAdIBZQ7X5XuzhgTga
OlajNRAUNLjGgYdTW5dZo1elOjQ0YZH4XG+MBXybDWpMz0fH6L7gXNWG49MWmVON
6q/WzlUaHSQv2xPp6pyQVW+Qlt+bUMYWKbu86FqSOHIupMYuUbIz+ZXwGM+zhwHJ
hkCQbLJkvI17uZ2jRJM0bw/y0+ENqcVRWxIgeG2prx74/yV6ESwKtI9Ka2NXTO1V
soNGcY5tPnZY8aWh3wnE11GOq6l+doS6MhwIw2+pH8ou/JjRmufYMqgaui038DZe
jaKvLvjl/Ho+cFbTOV1nHqaOxEsE0qqsLjPWMRRFjldFnefoIW07uTuUsvlBym/i
DDjXrXaW08+ReOSwJo1EFwYvVR2RlYLVnchDfcFye+/yfAkZL6bVCeP6b/suDlZy
4yk4XXrZTa7u1TDckuOBPkx47KX7Bsy9xUPeADsUnq3ovxNldOI3D93maiURZXWw
pIrlL/Mo0QYnHZg/w/u/zMkW4Hnxq6uejJEr3MFLW4tgy8T/9B4dgCIu51q/rJS0
48NDMeS2ixFfYHiJrezzxjcK6m37c0CyEl8u5vPpPgtFwOCUt2jem0IW2cNsEl60
zO71yXsIHRQxEwoRLXwHCaYddL3ZfhNOWeHas+0RXQPbYNLdqrCFcbVzHSedBkoy
PHdeEP3+3sB5pxpKajBXcXfUfgKFlg6PHOw43wWXPcDPfdTEGBWRQLsbF/88MCa3
w44Hnicy0bOYkB919/NzV/AB7oc7pHWfodK7qwzDHddBb9v7YJbKxFdl72qD+yap
tPPDqlXAzgMyqu63APTqbU30xcompU8WnJLiXTbFAeq3OKkoN8/wgIDd2QUZE0xf
cjBJsUE9uz+kWK0+xDQ7SGDV+HeXtHJEvS9alwDsNVjEhBLLNlhXpKp1vUcBiNrT
tjMpXfUvYJs5GbGtpOjjD/SDWQI/1mAIOcLh0ifx3PEufsTSamyxwm54x+o7VKJg
GcxNFnNn/lNG55aLLA/vTMoT0/79+xyn0qSdiAn17vKlAI+eV1nUzTyLGWeqF9PN
+P6JUtV1frYs8af8UbRzsyPWklAE5F7B7r9DdrHAcYoNUA7CBiTKaGjo+fV4j+V2
+HT03ffrovHcub2Amvb2/GZUxUfk2JrIyoO4lhYzmnC3WyekcSBX1aF/oYit4YLa
QL/5z3OeR4PLxLMg1QTBEva6YWHhsEPCc9WvzLCKeIDxB0K6fxILHNdj5Z0511oN
jUMhEVk1/rT1PFhVxC4uPW6CxRTRuXkl0cE4IVAw006LkMw8NdC9IRe0X46TmdLs
KCIdyBKRabHSRXFkuULEIA==
`protect END_PROTECTED
