`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VB+yOGw+5SxLRSfDB6pDln9mOSY0dL5ymTYyycb2ucf2TDULY7k4kLJEgmvofDFu
2hfyhbkWzhH5Q6d5rL0bB7yqhLQ1ZB//5V2WjaVZnBhsooulJAmNTkhjunbqqZOB
8HG7DS+cHwBLNYh+vFA8KW0Z4OPCe0D6sSJNGQWXRx5CtztOXcTze0JS9YrtCPba
jr/STYR/q0rmPi5MyHvqKNrWBx3oqh+9BXDjklACQ/bqc7UDoo57IlPtP7jRgpce
4BtAW+T1s9bg3HdchWR4TGuSPb4qv4nHZ5P/Go+cBDg0mFdPMvyqI3eYHV9fiadZ
5uIy6S5t3K9VIY6cOfHnISN0MhT684tmNQXh++SfJKNGb10Pw4MhML4YtxACtBmW
5eYroT0iZsYwpLYraMHPPCImOZMc2OFsBqb4LrlEd1gYVyMC0OYHFL/UMj4iysB+
X9n9JiNkXHa4XEvnFxL8Cr0AqLD+4VvHevcyw2yU9WZjxhnoS+FcVhJYB+MkpR7n
vg52ycmCCUg1w/chGMTQZ2/M/F2kY1uyx9L5IwPPUd10YkAcXmUcKQ2pWg0Rx5+w
VTkxFBOmArH+2igPe+n/rFRUWwPpzTth89gxlojO4peNtKym7QgkG9alFDE+BW1T
fWxvbm1ZoZ0qk1rzJn/kPHNi8lqgyiodsAfaXnU1tP16Eydz2ps8fnPs2IkFNn/h
AK7SPrmueTr2pNvzapwJK6FHjSO79l/S6l+IqGt/rZ84SklSb7XdA12/P3QbADf2
iT7xsZjYt4LBcc/O1WFAsQ2O+0pvgCZlXS/MkY7vTLR+TgoihzJ3IkxLVNLJ3Jsu
6WtmBTqyFEZVTOHYbLJ3g0ozfhHI84nsE5Rb1oPKyPRa+EeWhbNP2wb0FprNpbJr
idu4dtnPJZA25yHeIbnh5kB99+JWg8O4M0Ed3xwJ+l25/E0Zicc7BhPH5KWKa9Kk
MXfrLWnwFkL1Dgrq6jCwK17Njlf0XlXUB8R88+gyHnNBWElG2TvPWvFP/30AGmk4
c4qV5MXZY9O5NKLpbTW525FcmgUS4qW85um0GI4cu190t3DqkRX71DRSsZnX5GKx
mkPPmfxxDNifYvaVXF/LM7Blk2Pn2vALn+OtCX37tqqjlj1InlsvLl0lcNFtnY8y
TPFAplJCU4gcbHBwNxMa7Kz5LBDY7M+tNQWtMYFgCxTPsDqbGqy1hKBd0DKXoZHn
t9pHobyyCkL2nSjKjCgVXp4W0RBRNB9NO5Dn6RPi06s1RB7UZBNJ06m0wkE/cfzP
I0GUJ3sSzRYyP8rTQA9gGfHUoXwIMdY2JzlTpBPDYfNLpn5uxXimVYDmPmMwBmnU
KGr25/eIIm9DExaxx3s3EQCWJulCQOzF1IBLt/qKwVmDwoDwrLvWYjSIzHzqwyij
ARbc99T6avUTEuCnqXCh7K9U9LiNRu7lDL/+2/2nR060QCAGdkd3lmsHpEz2qCzd
qAyKpTbPQD4pwNMOY1Ghul/MmzIiQkQhIQpnmEoguFKWqTKMd++RM29hpYKJP8k7
uYfgE+thFsi/th9hYtKQrUHsN/BywK+Ms1ABQ15Daacy8xUwAI8qMT1SLwLRvxBi
djv8mRbCZvg1BcFWc7HmvVRiQV0UaCNouhlBmKzl8IzMNNUM8E/FiAO8OkZIaGTC
+ISyHT9iNDKsiOb1DM50bbd1aox4pG99tpO6wMtvRAqMC/G/wjBrUmHt8oZo4yAg
NSMreU+CS//gGAqx6sAokduCByZZyUazhrpGVZIEhcX9rgeaz1tUYwcYLHO9Z9cc
pfi7dMhPmn6ojLvsI8CExfa0zUpk9Bbx17z2MfiFxMI4rsWlpu7OmgsOdKmbevDa
6f1+A52xIcgtzoXDNGBYWdt6MEd9U7m+RbrSPByuQQh8hETnMQjjuD88PGNRvDiS
FA37CC7SSVHKlDaQVotlXmTZ4YSnLIOXzDlh6/y4yGG9ncqveGbR7NTjjk4twVPI
vnpAIex+QqWJvbymDZyNNUEypGoO2jLZeBnubssWdNAqIdPy+eXkN9evTc8wahA9
sRYFG39xfXAOYPNC3FUidm5sTVl6yDSNFeXYIofN491Te1Iio9oFE7/tqgfE72v1
XQKYSupwgZO59o4VmTkyCRddGSMKygyWVahMtysK8uqlaR7xE/5XXGK7MSKjaYbm
TXfsHePmUp1mg2723LLTFNzGizXizG1gEkas+hWuxmHL3SoQQWm0wfgroTW0td+p
ntqrvCtGYN76E9j/Ko0dkuxVIIkxRk0lt+hdrp2gHtlq6g0OyKoP9M5yIVGeeomJ
JWBkc1od6aG8+L/oxe0dSXwf+WS0YVPcWklsI2swZxsRj+trIIGaq2VPHUmUBAvM
C47o7lBjX5vlGbi0REVjWpoI6tYyCss9HNPfNIIRQgnWuydDxQU3cG4fflJA8PcG
V6IJcI6azUNKN8TUbOrurTf42YoR7ZI6R8kU30A4aDPGOD/PaLfudQ4KS1sXMkJ3
MtcmEUJDtI1xJ2KllrbmtKAlSn+AyaGYN7+i3YJK1lRaJfwMbd+TtMemY8AG7gTt
d8jM+mijbuGRurQ5yhl19EEW+y/pgAJWdEKajTWc7rm2qf84pCZMvdezF8RCnqqa
q123LL1SMgCK5iBWQdor7ouJ5DWmerCyKgW/vEQzruFbNR9BFJNvyf3Y1WX7LM7K
Qn6QVA+Inl7D3vzw4p9+BErGptpZbtQ7gQ18ta1HVzCtpCpLmv3Bl+MFZGncaWMi
h5IjsL2ppG3iDmIPkhlfx2j0Rq0myHv/RdWMHNTrmBd2VDW+N9Cqh6aM71XguX6W
68J55W1q1F5M5mg/0Vh1/NDu1k9DuBO1nUFYFR9Km5Z6FT37mooWnYC+Tj9rwsCd
gJuEktqWbL5ipl+omIU9eyGGL7UfGva1mfXwilSp+8dChZy0E7cLuAW+bGLQT+6K
Os1A7UJxqerlvafQq96EahmzGAkvoQ5PsT5YR0mdnWBShPIuvfHtzT/1WODd7Z/y
aOgxwFFss3en6zLNxJqOt/SWzAEUU1vOC+1nEz+Aa6t2HjIGZx4qexLfz5yGIvI4
Rc+J82aAzjZsKlx2ttJwe1r02oerTgiQWVrvlLtT4y3d5h6ECGtn7vBgVFB32JGi
mUVg8Gank4/L8/2H8lleCrFdpKGROxzrX0E1W1tEBYGo+GDBx9fVqNIoAI0Nq7yA
ZAtH9FxXMuUS04/+1ltMKlQCLaDCHeZqq8A3A2Rz2eHmrBo47ZBxft+s3qLR3mpY
lgqgavLR310IGR2LqdGNXfdJO1rfDpBFcaQDuM32Nw2p0PtsuyCoFGFqP2uU6mYn
l0pzprvmwhFkQqcgjfIM/SemybTOGICAAzTmPB1YGIdqhZo5grsG0yWGCNf2y1C5
aJtQCXvES8GBdrrRKpsZoeP1q+qExI2UvMSXVwqPWC0hG2YDFaX9WztxQJYIUvFi
8VtJjDHxgdlnrOYaUEyajellswYP/+yDxHil5pb+GRYqLbQP/US1WUgKNyMfmOZy
QAJdpqEeizLhNdABl7RZss51rDuCXIF90xkuaf4FHghKeEwc8gVnu3Vxkw9Yy8XF
bPFQUPhkkaKAcmDDFCApXP1aUA1VuDfKS7vewK+EyCc0RIanaLiCqNRHOBTp3r+B
LctSyj1moRkpHJlBKXm0ZGKFFj+ymOgix1Gfu804ee9g4ZHycjCp+/hahGiybjoe
HE2noS06Uqde30XzrUi5H1oVLLbO/xhJJWG/tUnOJG4LOGOxbQR/8KqoE49sVn/D
msUIiDCYGpcWbeRwoatSQt0PFTXkBKL9hasZzv40t24FdFISioOvacYgJ+F4v94u
6SEldYk6lUXUxT7C3+lPo//JSN5yoGkNJeVi2CvJLZ5pSgiRqL6T/VuWKHt9UMG8
3oc0z3zec9efv0XaHsF6Wz2v1k5tCDuYxU6/F0g/dZPyOFudGfnFlt0UGEgPrO2d
mta/QNhgy38Fgbq0J1aU9o6IdTTQ4B3u07TkEcB4xc1jhskp2qYvNJ8PKSv5XIcv
14+E5uHDPopzNv5+fx8/aafiAYQ7Pn3r7jO73ib0KZQLZdN3UU3UnQumQSUACxoV
rb0sv39Uvkkb3q4outqW3yoGr4UT/FoAJu56I/UEoBJsmNeUTXF9t5nUF5s/0v3O
gDblprQ82JTY8casb6kdUTwNyadfwitQQzmjSDz2gF+spn6IvYpgqT9ZvUHNLXxP
uDYM8nqPt0FRe9R8Ce4Y0HQO1nIPkpkuIFO0ypMkVqqWtWvTQJu4Pc0CGz/NFvD8
Fq0rcGaA0BqkCMfVvsI8GcfuLwBEaAXKVv1aUy1NC8pk9P3BhwtTT8TteX3NxVwO
dbB8eYXpa6gPPX/e0O+yRBudySdalwxYWnm0/N5RcFdP3KCGlkXoI8ZxrVRFArD/
CMcgbjTKULO+0RvEGVeemi3qO1rUOjaa5if2tE+yPBoJ1mshja3lRPqIpVC+zCSc
jNmkiS3n8wJS/5drAOlN4PHxvV2AsV4WuJtd2zoiJ71P7eKJnm8Jro8yCKXP5jot
7w+fipM+Nbwezsifz4OIJmTD0ZwP4Yxdwa7Au6KPq5p6ZKRy6SGl3VM0i4gDM8J8
VQ/WIiktmLQ3Jy8sM2vwxXe9lbMEVaagxpFdX3QZLIINmigyD4IvY+UgrT87wdOr
A5+7lE1WzJ2AgYyWOxWesKgeyORkMSsvETBowbaEl21Zj8IAdIjok+ihCKpKLkg4
6r4L8EcG5J3T8UInJM4z4F9AEV/0nbJGYS1iwpaL2+AEhos5v8PdcmmG6QIqHTSM
bU+XSlcjmWJQrE/TStn8NxkWiVcccPUTkBbtlZMeWStDh6zhhziN7H3TO7C7Ogde
Wu3RRq1+OyT21+TMmwyHvj38TofRYT0r821iES5TkirdusQ3oawGChp7blDVzyY5
+1+HqTVtKFyafNndjpQIh5X5tC0wxzM1WP0zFWX+DvL71CkPPD9hgNtukSDyDBuf
1qMkSUzrUmbTnmddfxwHo33TJOOEDKmxXalxqyfCaRvp2/WhNRvntQAhN3yGSASm
qdtZNB6VSiwJ3e84exhBrbnkWUI46Zpq2Ou2Dq8RFSXYSLEYEvKQDwb2ikXs1QMF
JE0BLqiergGj7hmo/VRAU5PlH9sdD9wNAtqes01nd1Lj3EwO0lnQdgyPUyExQnFf
fKDTxPMTiT0Ubkx+yRykPHRzH5fRItfNfNuAP0t10sYi7I6OLU4Kt5KM3eKLg8B0
83rvQTDDdl/LQ58UCva55sS4xGcjZ5LlMfD0ibUu9yFks71LumjZwPtK1VxaWLgH
l794f0csm3MANUR3xAWBmet8g1CIucWRbAbCVHeZdiiLAg9yh3KFLjk3XGbt2zUd
ia2NdPJGVmxW2qdctuATFCMfN0vPXEldZsikHwK6xziueo8B0GY1/CqAxm5A3En8
YygC4Y+twoopsWYeCpSy7U9hIMFKwe3osa+oZd2LHeJMB/XuHf1K3E4H8tDxCWxP
kwOWjx1sa3InRbs2dP7qx727KKV2+9U+NywzVYSkuh+qIgpnqxOTS1APrrtAE0R/
ILdejm3BTCfUumhEzaC1TNNtGIJ2dtFxEOLkSY3NF8RaHXcOldi9nogM2vdVcRHv
9XTZSLhwxgQfwkoO18Jtv7LZhi3kesz4WKk+AUP7oDhvokfnAzWIElGLaP0ictc0
PXR75RZe28gugLIsVjrwtfRoG0dbuZUvdhC+8yR57HgEyGgTHyAice8SFibnP5j6
DeGkX3O143js1s65pPaU7J6NkW7nuLC7c9vzzANCFo3tgosRlzSSL6iSr+IPfGuS
M2q+ZxzD/LSN8VglGy+niUD6aUDI+Iu/ASTfR3m5gFDxPwInUEXd+nvKawJaOWY0
sA1cw7kfEQ3gANTy1lHlpDG4hisSB1l9FXmT8BEhSY62nSilQdw0VxP36qotD8LR
YEw7Z9bV30Dhij/IIijC7Rm3Naqsiv6LSZQGVg0MXo9QQXzMct1Hu7LIdv7OZLBc
YnZU+Ga+vScRq3lfSinCLt18FZiEQ9h9ULYWsEVi65fygz6G7hK1vz6GqAztytnz
vdWfLkqQ1fC7Wca9EPNMZ/zm9nfIf3x1bA58+sJUN300rk/LCVVul+VnhVWE02Dp
WRb/CaaGbfCAht51he5Rl5PqDN7Mqs7ysmrufppAbAi8ERKXpb6SDVTxyL5mnJZM
+STdG4PIbBqvo5JnoW/1La+y4AkMD4FQaQhXJTboSoFpxO9f3HBZj5jvk6Ij9TwY
c5VhlDS2pqM29c9oNDGg7mEN4BjX/iEfiGCus0/l75JKRebXQWCWNpEfzt6o8SIV
PzRaQiBfD7bclhqHr6IcAFJiaPtEGZSZWq+TEpNsXvdJHF18oGT4BelznkI1lyIQ
z/Rv5hEJHfWwgW4O6AsAZREexdnuY2BmOkeeMclyZlWAUfTTvlchz+Vgdc2W7VA6
82bFhan35iy55Ze6rexuNjPU14MDcKrBRMC3a8v5ZbcBOKMVO4JEL19xtiDlMvD+
UkzKJ3xLWNsLj3I0oWJoWlkIkK4sxD46ySI7ZSM1AX2vwwrgoAhkfK9PX3ouhDWm
/ZGSuVrHZotgydckWyX97WdR0bIcoyHr04ZIH5QruzyUw4eX8fUpYhTFaFm+94Ou
EL31nH9W+ScDZhAYEt+TGzN5/9Srz94h1uCYXg0JQS0Sv2CjCnonOG1JXCwOc/ql
+pDO2+M1iz4IYmuQjNr4m7m6mF5Smxkti7Z7tiLfakwfgfJdZ73xtQSqeCkSk53x
ckXeG3bjzWjh1N5EF7aPHJib9McVQc0wIaMup0ARiqMfmGDmQPUwHcWuLtzf7YVC
2he2xHvM2mceSHIMteOZMks5XMQitXhbWx5+eNPG5SJw+67ndoi9KtsieMccuhDD
dwM5YmoQRadQjqcJo+E6hE3b2QH2xdmmS5OzHLHjIh3Rxk3QRvCmNMO0LbCq15Wa
zplk2i2eZun0diAp7lHE3FtM3rCQM45t7Fqif7/W7QN2FrEC4nFt/j7IIhwlLCZL
bXwIGNVRYrILo5rp9qE6B5NdBkPDETOEAvcGq1NDQCs3BjkBxd2hHr5t08UfKdZG
8zCtvXNBMoU6b6XWpdIUYwKKNldlQAf6lKJI1aCaxbOZ9IinRrRM4Kq0wp8ZDDNm
NZDg9Icb9KUS17c9E4AC8uPZTYe+Mtak2n4Lmm1AHvg/NLuV/rMbkZIgCjCyZO/C
a78yP7QJqds2GUgI+s8kIc7teB/9XdDHICUrrKrkp4e5ZdvrOebUcwmsoz9w/BAQ
WEJvwZ7ITyI50g0Uw1lGOAD/NIvIxfYU8W3lD/hPfXveDyHKgi3Nr7BJMx6pabHs
TKID5U9Ouv9rac2pHoq/CRx2gqjifV1hWqqdeIgU4om+KwuAyZFIYmJGbeM/YXJd
fOJyz+1d1ptxiP0MrG/yvY0OcG/bW9va4E9Ixf6DJ9Tzam+2o/fwcusqijXwS9Gc
8d3i/4cDQaRJp4YpNsS1S3I/JvuwsIBUJgSRIqxyTQgij6/gljtOcYo1dx8OVMrs
X6kGRqzJd1n5VDDQeLFCnypgYKe54JTodpdsyiaP669Kf9yNNaa3JY/v673FoujI
x5LDS5cfY6FNDQAlb3eUNyNG/GdiZofBFsWOyjroo7zxlZ53vYDlq3skafM1oKZJ
oJjx3+gmTjBCjf+UMJpJ+PnAagmzWLEIcopp6sT9O0OGLf5nmkoMhVqohlM6RT2K
jo8dEEpblwcW+YmZtol5j0/9I4bngPikMr6RlnBlZZKZgOfH2aopESGA/ZwCDxtu
ubJnxesrbrcRSPQYtNuj9ASLxUPaB+OIV12yIiFmUJKN78Q+RT7dI49RJvxCNyXG
a0FyvKVGSuW8LWClXWZ0BoCQoElTCEAnWcjHjcp7KgNHmY/sJIuiKLVL7kSaJTz4
BoaKOsTf1OPspIOkXJMsfhopD/XnZdscluTuexoytNvLdWNxZYmYNNjC3+AT1XxX
n36mf2lMXZSFmc5Sw6xYJz4MNEdNYUYwWSOL7iMFVqPZL1aEDgD2cxQXbt+JyOtU
Nru04WQ7YgqZ+CAiq8ZK0aTYskGpJfhXUFrb66/MvUPi2tc+yI2JVUQfuseXQ3Kt
jlbHwtupE2DDSpPqdEXANHsHffI8vkmcjNuwFTEqcwI7O59X1dTyZYKC80PkB7FP
hGZ/z6ggQy79JOIWLaRgJaJuyOzfYaYkbOhmL2xEkSOdaUDwKPyMZGVT1CY7Yf3q
K0mTBy9+kJxgl3mL1oomUQvpxiXgod8QgqGlc8K1TEDiZtQYQCivm8PybHlzzjVE
+Q5maGSEpNek0zwAuB/XkPpeemSuatrWofrtC3lM2GivI1bixhLFwy7tVz47LIr2
lbXLea0rGSFwBLZy1Y6J+Jla0oosKsvP25pdzj4l15pMMsqEMBKpEE8UOlYCccXu
EB+lhUx9upd+4S5yoPo8R6uPLfYkE2qeM7nK2R1teMa+pTu2xKRcfoN1AZL5nDRi
fCwr4k4cDAioCyqc2sM35FYTl35G9PTLUtwHFadUrRVgiCcN1Yj+3A93FOto352K
xQWWr/K00bowKSkFBcutW2ZiotUXBP5LKxwaTzO9Dr7y+ddk5nhF4ZVMiJSkLLMc
yPS0TME5Db81uY6rAjOgG2G6OSb6y141zmMD0TzadXifDTQRFf4JuG1691oKLr3N
wxdL/+Kr8iF/mhaszLABo5gWAgyAWYJ7IbCuIJ8CAeqMp1V+aB80rckRNC1rWdrD
a8Lq7qXaV+Y+B4aiZeDJI6KS1MYfP0bvtM01YBzg5yVAbAX8WjmP5xh5isoGHz15
BC8LngIYQ8kmPzY8bM7G2AKyTW37N1arbRNONQkf87iPYgfE5Bopi3opWFOADiLg
OCPCQYsB/I3Iq1YocQPGdTkymuezr3JL1Gd8CQaKQGKvFAuoJX7zRtKHKqaq/LAk
3miq0WqkGstdepUFjF1dwQmARjcMfCAIOQw8pdQ5YgrD0YzHD/LqiYw5d0uLkWPa
4PtnqkD61PLV0jijbjomSTBQOm92+tXAeWOZRj4d5zSaFioCIe14xVEnikMaNtut
FjoYQjXf4zHM0c8jbDjUkX/uHnrKk8AJeFOdpiY/AuS0patqJh3d/kMqptERkFMN
53fA/mbTjWZLcuhNRszSXd0WXRMMXgNBFrVJnxgrHFyKpKWR3pWeEjygg/ID+NKO
EGL9R0DqU1VAPFg9jdkaO0afE14ASpk8rBdOOcgr7PtRAI6u9cybEPOS8dW1CyA7
uuPpRUddU6MA18j1OA/M+Q7WV1yz4du4461WCIMIY/KWwG8EBVTGh6sQwm88ggwW
lr9Ws6TDQwYigR2A3+3YfmpsupAvZBXXrpktcgUBBb+HRAk0RjV+czKbOFw9aokA
HplGz8uMUzdHeH7ARd8addY4U+BvnHOxhgJBwP6NJjAHxB7rw/G1KhifqiEq8Y+x
bM8MdcAR040OFwHQKDo9DGV8i4jz0zwLE79VLM/6A0zxGACCARhN87zeqfgcdbLX
1AT7mgwsdvPTlkQPbtllrASQoCr0KpGT33oggnQELP/otoUhJpcGUjzo66TkERdz
luBf7rZ7SeE1+1VAeRBixfSmfzfJm5C5ygbGs5vbAcCC38yEnvbFJIpsCtnEqToT
072/xwTA9u1pN+4mDuS6r/4Rfrcl8FwOKnyh6fZNlMBRXxtFw9mEbthw3Evn9lCz
9MQ3J7ilbM72gUMsZH+K3sSL8L0XqHB/glb+YJQ8c3W8IV2O5QA6FYWaCUPrCiEu
YKlbCzjRjJ65Pox2bBFRWgO5GeBmTTxQFI3kYIdY8ijk3/BgQbZvEJ1aTlCvPXa8
/zPMevvvALFq/xQWfth0rWg/lpqQNjP3azOIur89d/cfHZQARiTlyROXHmfL/5L5
JCWT4CuV/JJ/nbH0oxGWSkAGjXIPAsptsheA+hnNk3u2A5B1pRUVrhpSCQpcIX5b
ihgCmNn1sUbGt0xMHJl5qE9YfRUCP0oXEL7APPRZlNhKvrSAeHO94YLcc7c89Rng
X0Zv4hkgyg3YDcF+K3XI3IwJRQOIToRoKCgNPnc4Lucvc6j5Am+fl1LIZzT8w3gg
smnBVhSlqLslpx28DRE0w7ObJ5qw35gSfVm+0OCmChXNUpkGQ5STXOjjiP0t+W6/
e5O2mohIMZ4XDeOYWLjwrUuOzUFlouA4q/fmS7FUWLEbStoL9/qw/joYz3FYjh2R
8dJB72n36lRo+OeWzdQvIFxjpQ4gE3xm4IZKH+d1mrd3JLX737frSv2jsuUaEwK9
iZrPhim33OMjsNf6N5lqmyQfs+ai2jngtb04mC9TFeqPTTa6YL6xmw3m7yw/27TX
2BSxeWhS68qTbjUw57oZilXlQuVn6FRlY35eaAMotC4sRQTgpGrmrwpyhKLOknyf
o9hRwPFAzCbbCEmH4jjstrztJeMvL6TRWZMo1tc5pJkNFzHXZDA6a6JPaquer6Md
ujMJ9QqJK4O3Y2x8tgMlaXWyoMdMtOWAv3IDmeLBKPlaTw8rjYNCS2fLUnE4irFA
T6EIhMBp5LEnuy0JQzuR+CkKL0uIGUF1fPz6GrhOZPOMBQ09ccS2//b+El+MDGBT
kNiojk2Gqd0FBNtMZanKjuhkivLKsmYbeP+/Nv8vy29J83PLwE4Qs35AlVt1+hCN
FfXMKM38B1xaxIodhSsasnTvzM+b7TPdbGsx5z+y6d8m7c9CkxHGyoGczd9t+vWs
HiY/El+qdAguwzPsswO/oWht6MV3tlnQaOs5EJ0vgHYfFEOiK5Geac+uzupO3a6/
9K7YFMI4BqdNaD9OJkqh/GK0o31XnkhkwhSU+i+jeHYlmyDcAya4RvTPlGyVHQfY
k4rdVbIhWw3ALRWdK9qieH5nE1LFxihnTkOc4xfSWsTLN2gwkx42SHPzQ1CiXHY4
Ry05DuIQ4CqbaQKee5aJqVyUEgXMkXFEVkRalXp9hud8QOoCEIvm7KW2x1cUeJmb
eqdTfyPyplW3GJYGd2LCqV/dXr+SS25IjOqVhjoLoc6ias42Y0yS2VG/EdMaRwqs
15I+P/C9Ke8uLFddeK26x+BtF+6HWCTCk8C0f+wriVH5TlmRzZMy6GhmD5sEnxxD
WwLDLaxp3hdZdm6GUodvk081jtotrqJxFJk8u2mkgJaqjRlkQDCbEHx9G8mqX9bd
zC87a3sjYzG+M0X7RUcKDT11RHLw5GXO13kHxAXAR/jXk/HjPHZmRuSl9qtXpF3Y
FdRVRQNIxE+lOX2zA6d3lZKV1LaPg+0+OUGc6nMtnRXv3S6gJhoyUWMhJM98B5NS
Jh0p2TdcMsl81nIFQen2mRE4ykwAOvsO6PI5xchjjnKtR2O/m6TIWuX1KcSxdwNQ
CzPDDt0inG38jo7iZUANqfrXjo6t99sc9fxCgiFxsanZ/lzn45rnMOby049tVGMv
7AGcGdvbbiNUDvxjGRRDaiiw9aXqr/Ylqr83WEMTJm82eL5E9+0lFG8CZ8ILFEqQ
rgtiS+w9TIaH1guyvqRjXWq6c3YRr3znB2QH4GvRJ+AMvu8iZi+BfoDl/mXRY5pE
XwXP0W1YB3lmY+nyRnPaGN5zI1oLMN3m2mv9ZlWDQHBlwAi//F4B4x8kCPfXoJ4/
umGtgebDFGTAxHbCzWrBj6avpfuVa13NMf4fw+NsL4w7EntOrI0x1ZLsm7Muup4W
B9/XuoHII/7/kuX/xnpE6eOIUkFqVcBBCB6MfLGvMeosJnbGvMuU65uzwffjnb3a
bU4Kl1Yd3Emk5tGl2NtPLKdKS98Hxr0I9MuX/mkl+0ZsBMwlta8Lh3tbPnul9KWB
O1xlDRmAytWyE5yjxQcDVhMoMTOm7IMmZ0uQpBPWt5SrqkJnT84+QTPgb0ZHswzy
ZgoHZQHRYzIvgo8y5LKklY2v5IkJqeG9OT1EPVqbsIn6MRdCbz7BwrhayiWMkeNX
s4i41v9utKvBXoqBI+2w8+Ob6wySKpNPnzC0qoKl17b8xaFIKpjqW8tfTum39V+S
e1IrSGn9kF6O3DK5EAfTSGIpVQpk04+Gow+KaSzrH7KbTC5/hJ+t0GIKQOsMJDUw
mD7A94d+/pMXJwKrw5YvuyD6y29bchY7py21f0KuZYp4mozLY5fFuriCm9IBKROI
JeHI7K/S9nRzlJVj18XKV8zi8L5vqWgzhRO/MOlhFcyr70unMv9CqEB6bYlg21zp
wo1qiuIe3UO/RHOfKPSESkE6CR7nK6PtKpEqA4rnd2WjJ3CpSEVz3CvHYyk990Jy
s/xMaFYHZhsPEzG9B8vlSaPvkh4cxG5oxPY7/Tb3aTXC+dOEWNz4etjQlPAPCJOs
+pqb+0IhLfoncjo40hZpp6qg3PeRyWg2QgIfYN7hAeXH/neB1Hf0oZ2bMoJBYurA
h9NTe2xtXF5ZveO/af1GLijbFO/2/FYeQfHScY5Vli2uEu6flkmJcyIX+PUHv7IF
hmvgtS7YRbUcJzEr1mny+Z498yTqUJqqAQ08SpdFaW8MpJaBp2bBDKf6Sk8wZbj1
MAWsMx/7dqLAd4YUhm39Eq/AyoxJOijCC54yGhmxNTDlchsMez/qswsjCsJNnkJs
/wmFTsQ07IW45UqqkInVI8AprWUWZd0M4oXU0smWkemtpmugx+/Lj+Ca/0BXBNEC
ZBQf3j4yiab2aoFMT6NmTkm+i6NAXWqb4RC4ZTELa94oYhldvZlwhsnPRTvIyJ+Z
q5VHYPaYeVAqTZk+ednpOq+WrPmP5OvbtgfdBJ+s3jQsFc4Q3N4XQ+2Vdi5bH0P8
AQ6uqFS3a8WJihB3SpRO0G7WIjeYu0KZokz/3j81gLzTrLt54QFr4lt+ZB8QVO+h
ihZNv3PvY6F1wd1LDS/r/c6by1GSfLdyJcwu+T/U5NAslYiS9kMuvmgA/phT7M5q
4tbfcJak3fI+77qa6iULiu6C0vNNmNCCOfXfLoy1O0hil32CYpcX67CuriWMqNXV
e0boMqkd8eSYzFuoxODetbNiiLQksOahC4NJsWC2IMEPcZcl5GptaLHCHF2Gv05y
0COzQQGJR6fvrTgZx9VoAAvQLh0z6blQbI8eMxWgIn07VgNDUk8GwZFd8H3jt4Be
gE6VjxS4uQsCb8QB0DG2i3IqcBAQbHH1hlrn6JE/s1s0ZUoVybn3utlpH6hdTzZS
rskXorYOlfwXaChkaeAqYfqLnQH3y3Jjq+2EKoz2aM8=
`protect END_PROTECTED
