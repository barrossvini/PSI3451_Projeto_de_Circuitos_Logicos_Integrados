`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70i9f5qniBP5ik43MdDX3wwjuho8JMKXoLoDKXncpGNWOS+NNQG8T3/2/srWjqU7
FFecz4nGHh/M7SkEDo29wznXbEiQfyTuGvoDbgYQsdfrPTdrj9DW6Y4OpnKeOHNY
s9TAQWM26rxDsd0Eae+qvtVc0i3HSYOzgy1sCgDRBTJtSWQXDvCNyy91JL+izelC
5FnYFGlUSp5iB63sPKsdu+NkQVDbP5kocek8YT+PGCoVZtAASLOpmGVe/vZxgUXI
bLbPv1A+3+BcYSqcRMCWIkXL1xq3MESnEoTZMh72YeVJARoANrEXuuyfzURbWiCC
wi+wAUEmg9n3e/XkZF+bf8FZzgyPL0G2pwD4+eDloofwOX1S/OfnBhUMhv7/bidj
3hu1hEydbw44HmHczeDwyF0xMOm+brBkkBzhQE8IxxNYkwxRCBVXew4ygb0vD73f
0/FW3Dki09GgoNRUK7ncXWwj8/w0I6JXnyEB/szw6MeuU+s9FtFZCvj0635LxCSh
xQV0gqC/b5RbD+cqjosdUx6Q4inEf3zmfrhkRmJwCYXvX0tCRU2hIXs971YmgH6J
OHDACm3AFU5C9ljq2mVcw0QpdjBMvuP5iJc7xA5P/XMF9m1gQA20CRFtGR7B7naL
dBSR/XlQdcCiNtd98Y+JqVlDEmFTPjFM5aosA9GLIW68m7x3HsdDI/C4unzuBPa4
vLdFM9+wGpaCeEAyh2r+kb+fxxYE2kR3PatYqEv9Y2KpGfAv1MX/HoDtE2MY7qgU
B17jr6KzhJ7wwHEshrEj4dABtlbW8D060GlBZOot4hEnnzv6FgV4NdQT8zyHsBc4
w1tSBtjuSUbcXGWF5s3pdu1Xibvow9apBgoA8/ZkJo/5IC0AC95RsTzAwGGPqzQ1
kOcaXvUOJK6UFckr9vGwd4DZ8coNaAyHbKihZxbN7+ogVjpswyhBFbhHErH0r0Yk
ziptnJPByhKdLNpmShIm2c3oJB9Dwq8C1QvcINz6aT1bVwitMxKpePx1IqgjCBxV
AXMURLfcGk48TC+jlrvjdKekMSKNYchaWqav36abw6U53PMT3sB1ZFCLvQzZJciM
umIQRjmdyFOCl2wvLcsn0Zr1AI1G+qMpW0FpAQ5HpGOqn706+dt6SjHlvhYZTPMs
`protect END_PROTECTED
