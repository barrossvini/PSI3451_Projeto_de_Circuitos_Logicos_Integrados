`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H/SYTQfzL95FlZ/tAhqGEVR6JtUm701e6FuiVwSPX8Z6mPBa7sVL8Hxx4ozU44lk
0jAXUbxB3V0qcgsBwZtjXtDonmzNvKBPy8Fbn3KErbz20HySIxy+n+tmJuBzxCop
5W7BwsN6dSMlPkPBf2n6QXgQgwFDGwIJvEH+9g7Uc2DbTDXaGu7JwHAom5bst5sO
ywK1Bgn3SAX3tIzbPoWblEmqhhrxtAX8CJnY8ctHXxBs/0o8KrQRElPqp7nkLSA0
PrZLHNRD/lGhuW5mlSogMU8DkkpavKkNWsuzLdtp9/l1NJkISbb62Kcgjjv7zOig
pHABc6cOfFmLFEsN4S6efJh6w4676aTmwZX0FdSuwimI1HP5pQ39glOE8QljGGqC
pIkzvL8zOXIqHvORh2Suz+tULa+stfn5vXA6q173wWzmoQWjS7GxfkEBQRNMmZ3w
SJPnJ+qCKxhkxNCR20PiMMuy04Nk6DHbJP3oiY+8qDr52oTLL28WMqr59tpnMaqD
LGRyPWU6A2QFU0aD2z4BA15HGD0XZc3Aq7mOnb1T3MdKoiUCDxQmeE1Nke7RrR0E
n6z5hh7oHos3d+ror4g7xGIqEg7SVk4kvwhJldH6a3AWaryN1QTLZbqcQ8JUtGwo
4i5QHPHrStwRbJuHSa052nM2eqzcw3NGPXMidaEed/TNjDWZlXC1PDdpTYrdlwsC
kJ32gYdtlHKjc5Yx69rM72RbL4CYFks1MbB9DSj1zGGp4DeLD8Fa9+NaS3pn65g9
/zblELsyMec8DxHEjjEyJx48fTtUYFdJSlEhybtHaJTtHKGG9Ox1jz3cEsS9XYgF
SHWZ8lZiLFq/lqWYNBUgYmbYDCyVm7QXkeJgbRxntdid/b95aIFu9K6CFawrJDaF
sgm/AtccZa6bLqmoCkaUTWviBwi+PUTD8rZP8u3JuOaN27uhUBrrXSvE3SfvMsAk
2sn5bOHn998+ImhjQ6FFWw5yqs0CEvqGslidM7/mFAezzXKzAHVJRvvcEet91cyh
qdVGcsurn3Mf8PSNMJd1RgcEqLlR78/YWJQQ8FmTgoKPmMLYxEI8OzXa7shYc9T7
TV72LhRFvilU+Lj7mo+VAhzayhzqpmi3kqxL1+WF6erwHDZxBJrUGEEcdhdVJ3Ij
Qu9034OxOdlIkdFMbSxXSevMH/ro7zAvnfRhp/c93lwuoEaK4+rqM7IZfWLVzO6o
q/FD/1ZAeYsBtw7sTJL+8XF/nHJY1rHYocX13+YCffQzbjPtlu8hVLaiMC1bEw48
sDBvqfL8Ha2JPLrjFTX7TlJClRkFm0wV15nywDdJJR8iRTDdsuJ39dNBlxDhD3rq
lY7C8EBthqKt2N/8Fhss4JkqcXnN/aI2Apva/N9kDl54ReqY+/RtcX6vtWpuCWYy
Xf6auMRdPF3IP3qwoewzlyKVjwmxU3axOHplxizwUm7Pijn89P8xheEAw7Lweohr
R76kePA7uvPyYftV64cfHp+AhLkiRMCUAzFxWqCmiH2ll0LLxRWWN78x/AOtf3DQ
1OqFNp4o+ME59n5/td4eVbaJqk4w5encQ0ViKX6cGQ2L7OSaNA9XmbRY5EjdQJnU
21tDj7fQUiwoN3Nu0oIRMfCSukpLEt02IpoEIPBPYC8kmpTirZahviCntksUp5UK
qNB+yJIsNg7i8b1Rg4uFj/POGqX7GjA/nU267ScST/Yl6TeEoBx8HKeGY99mn0rz
G1X0rQaH2jx2STeU+UxFTDYk3r/hIRh2Ivt3u3hcgFkD+6TTGhazRAEFZRzjDhky
SDTBPQUUEzSBWhTn3UN1c8O8XeVkJASFZKCYeuIKNPPfG2r9W31fa8KnLQ1Okfkw
Oll9HIZ6bxhvOwvPNwk34T/4R1WWrYyoxKSQ4OtmxUhhyyEhfc/CQBUJ8akXjiqn
OdOfnjj5OfVIFRGzeyqZIhMhFcG4Y4MrbcOOK814RSWYA9YbUciUcU9UkV6JxH+k
/J2Hrx8OESAfS9dm3loTdOxihQD1Yoq3RGv1ZOZkcCjGBbm0pCY/B/zHFDH8/rh2
vsDyGO6ogKDvlfYawZezdyQ+F0abfK90lfK/y7EY2G/7feqzYXp56k26tUQysJV3
nGhoHUV9rlLfH8/60+J+VLyNCUSFePO/sZz7CJA9eoLdAUcUW7cJSV7S6JAgZ7ZA
XCAfewRsuFipGDjAmK3vrghQ5kn4EdTo3n4dhNFzqVCMNyuqtmI7zdXDWuIjWUts
SJmSxI5LMkHBUC1PcmJ1QuveCdjHdbycpbGiarrRN/gZLskvwnDwCxnaQU63YlxJ
ur2XwvMAQDVBRtRVce39gNCOIf01+Q7yTtcssvk+eMJYvh/tZPhki8D4vUTiBj4d
eyFWVDgLDgYv6Uq1m5ZtSw4DowE3vBNQFPHTjuwtBUFQ0jWqVShUCOnN9bBAx6kh
3Jq+H6XHAhiPA32yAJRoSle2YpxXmtBoO40XMcvX8MbZ5KXXg46xUSpUbfOX1nVk
5pTQrDT4w0ZW0TZauEPgSwRidxPfOjzrUWOTGBcomCZvTBV3UJuaNXtpXzwag6nK
L7zxzLLG7+NBP7DaO8slfpds/+jP8vKWAdpowagvnIa9Dz81VC4mVWx0tqG++jW1
IC78NmcPx5pyoiI2ubU4qA==
`protect END_PROTECTED
