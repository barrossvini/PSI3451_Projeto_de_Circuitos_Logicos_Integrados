`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6tS1ietSFirmOEoqPQGpA+FfUCUYBCmt0i5SyjM/68hGMINOoMeZO0RD/P/S0Z2C
gB8HAIFDjWhxGjTL0lOH71W5mt5LvWprZ3RUup4iVJvxJgnwsh195ulps/9/9Ej4
QM5HOWO7vNgWmLZlEwEAzFzIMJ2Gfh4D85nBiSVLvKGqk2h5yNauMnNddCGitIzb
9OsRuj3mDBXCpUz82YvO5cIXCzWJzCa6xQ3C0PfQzm4tC6YYdro8cJK46eBhuGbW
9nbrMvWSPe/yFC87myQAubWJ6sTnsRBHm9irYlfO8wpWlZtAvwGpeL6aHu9LAjQj
Fqcn11WmjdI5huAL5LHOBFtAjhL6mwJt8DvL+RCi6cUmfS1n4kQy3wkjxBYbmOdv
QzIC+dkK/E2mQuKuNQ7AX++/eB8ZLn7w5sKyAxGXiw3LrRfa6YUBthF1Z048UwK9
/ubPz0+6G5XdT/xlahGlPRxo2e3VjK0l3PRcDQLIxg4G26XB78quovVamc4t2O+g
WZtM3MwTWvX+p8U3oHtV8jxu0NA9u2eUheNKYBXw/ZHmA/zkdD3NKgrbJMLZfrCx
kqD14R9XtsPBcGOO4OEuYNM3S6uaYFVUpT2PmE3S7+RXHYJXk7VSLOOInDyiXyCp
yU/omYX3enuFkAzfrCGPN+8aLIslMMFzgs0Cs8kYpca0KNe7wWrL8nR9oOE+ACtr
fEGHnHKEJNKacPI7l6HH6Y+5+Xou42JnyBWAgUNKuAM9y/BEqEd9G7OleY5zuX9d
aAeqH4IEfDSTmo1NL0ZOLA4Ih6xZdDiIRa2Rc0bNGvqSld+w6Jrrmz3aZPKKIWkZ
toeJTUMCSwfFpaLEPKJSGIUSTZ3Y+pmiRBWoHm2qBC2GZrkaWBPiWI01S1u4fL+H
`protect END_PROTECTED
