`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
npo3kwlc2ReuN14wbOfv5sqbyfqilhpjidI5Y1lhYahkokoECsCudNPxZrjobugX
BPrPv+zP6sZHy4qZExBQwBudcPbvs3fWDWttiQTrbTfdOXp/kBoEhVFyFizPkQ44
fn6lSo0peVDc6cRYYaTrsBE53uI42iJaIyCHkMoCRcSiYAX6Gjx6mGMi9qMiu+PK
prHXDqPp7YlvbToy6X9ax8J07kD+x5qUv9Cc5Ddi1qxb5v0XEwOBKnOvATdWS+fc
9cR0Xxzi5rE9ERCHYvfQ7EEO6lze1ik2m5ce/nk3lBo2zZDddneD5xnGYmaPd/S6
NheCWqdavuRAeTNNPednL3qhCLOjDt+ySDQVZyjuyY5xDaQ//rmI8heMQu8BHQdD
zEjb1c3nPykTtLMb80WfGz2Tm5xVsTToyIbHjGkq56ABUDlkCNcNbsbKJPfPZput
WnIovpM92hycw0DlhSgKFQv4rsqfa2hYfD0T9H9+oqLBQjxSGw2Y9EzXSw2RIRtg
uiKuVPROGwzYbL7S4APjSHly2XpwZSsrCV/JFLLdfIPfD6R4GbvKAXuVqtwAtDpD
E+rxM8faIINoEKW0Jk6Q9RRCsAv3OZHbejfpWSgXjHT01Y+khK3n+t9r+YWYTI66
PMxzdRw13taKH6KL8IOEhcLduW9qbP1LHZhYIXsYjOtPPXpSPm7HhPXgc7dYVd+j
EBTEyENsm4gGeI1gnm1LHb7MxGBRPitar/GMJfusz3pWybIeqDhqcHKgUZtFxdQR
XElxgaoq6A/gwdMuyFVLQwmGmkFIruaD3v0gdQz23RwPcFy1d6YCGGlALTlGvijf
rVhd7NjZkrrz5nly0sD9TMPSNx0SgUui9zhlIySYOHip4wpGZb1D1fdXL1UZJVNi
/Jf60k7LEoS6XhN1l0v2F9L2GauQo5Qb+d4RmQZiKMEYYedkf32Aff3FGCsnWUZ8
KNsB1mYhZzBHW7LUYE21RM1DJxBCUWePt4jsT9PnWo1BTrPxHD+mrRUJ275kj2gA
oS1hIQ5lVy+3D9aNdP1crebHOA9EpaglZRgeEFjSU7JkiKKguj1J4Nmi3szh8vpQ
I+xaSEME539dm0oc6ptsHgjtCkjScrLJdFGOtVd1y+f1JrjdIK4lZx4uCb5dFVVq
aRuyt5KvXxfOBdyG9H1pNNRWLMBKuH9mmZPti1T6l+VrjeLDSXgb/eIR5aIcnoAW
TpLvdAvvFuuMEEEWfW3+GlTvy7eW5bkf/mlZn35XRJ2Rhs4iz7bSpcQ7xVt2m+5W
TrXbt/sqTqU4k8YaIHz0OxjvQvcrI+++DqPglbHJgn+QzKc5GfQ2zwIeeByvWcei
TOeyDALDtiSuJQm5ecOF1S8qDgpzNmBIFweHyKbjDYmqUIchvyuLKtLmtRALds0l
my0+EY6hb7Y79J0Mf87HY/+JCSEJJWpe/EjPJZzL3osTUG1zaH70DjI7CXJgcncN
GITGMrKHWQqURZXlgtAoxRRki+DBBdgmsRGCjoQaIOyRRaeJFsB//GNTsW9nPz36
Mq6ez3EZQJRbiL+uNlmNgG/iBGOBAjsoqWmRqq357T3CuXbd//F8GneYUihTC6w4
IXjKUaKIVZaLCij+RPCvXDkfsSNjJ/8pT+bPAzn6qPhD2zt5tl2SpX45VEX6nOvU
VEVDXJpmz9suxxKNdhZ/wNz6mLCNwqYrq2wwMPEzITRGRizpA95gU7dMPLbP4gc1
WmVAlnV1lEygV+T0g+Z1lWkAPulTVpNFm3u8RQymd5hu2c4K/KsqCBLj3eAEHoHk
baZo0B0LjZfPXSac3rIfbvqqMlCxBN7j6UOj2zPEmHENNlFWRtaxCGhcwMMjiL61
mpazQ8EQNGbwPTssyc6oU+B98IAZWe3nnmqYMGSybJUMCFb/9rjswwDfePubZbv6
yo33/HQTw5yLa0+BwgXnd9t4pQcSTPdE/cMW3JizNE2f3gLNOTHTFCl977WMyfpv
q8WcYMaM1fOwIbCekBT6E4qOfxN75inoDUuwbBHi9eqNf/rpSEv5Sx65AalF4vYW
UFjtjR4Njk0xDLdPGH7CKdAWDsXp3rZFbQqw776lTPIKjO9NxXctMzDwkKw/iv3W
UPwj4x3YU0WH1zQngJ3+pCTtjt8b17yp5qzjTG7FiuwjN5hajUKe0+F4OVfSXW2S
zh2tClI3VteNYxRLsQKWB8Yr8XtDkARrMy/dHKcBmE1JeqUMpOE7ZYthGRyI9M6C
GX7oYZQ8RFQjynM4Wb91Kl81kwQqxE9k9fm7bazHczX9NBrsv5TWKAVn4iwdSgrW
EnskSWJ+CL6h7Y8KlwIP3TXtSNlgAU7DqWjvoRcrWCrvXHGTHacH35ZVMETqdcKH
Hp0LFjlHkKH/uaY9rg0fVmuk1F+B6v5KNx/Yff0IP8mkxKWYtYjTBf9fpyx0QTlq
blUDtR2KNiYoJBWzHJL7t8cOtCDeBtZopqWPZlA9bZSWk99pqsyGW8M0828nyavy
AiFN7auujPebkK+ij+q9w9HaXktnoYs8HMluSuM6WxPOOyaJClmnG91rhwYCFq8h
FA5ID6pOEIDpdlBgVdygtPnyuZ/xIVfTccizB+LzgbtBHtM/PEzJNbnWdwUbjdV9
e3fhOhJDDNCuSTVqlZF95eqtcmvt7Nvgk8V2kJgrpPRUSkxbJXherv8n/3iFwOcb
bIuAiRG93lsFdICFz7eGHnoAMiz8/3Iy5wt4c9L9syfBkNpd6cZ7x5goDueXH26Q
G3nNXVy8+wA1KH/ltPgsmJSIKxzW85xySVeaWVkO4EjAEyh8Pk+r+9b/ux70voIn
cFZQ1yVumvuCglsGzpiTWpYjP0sNJxA8JU3opUHQ3pqia+W6b3pyUKIeW8mDEAYM
IfXbkfQ6RIXM5HY6SlkTca8X8i3lXnCS4Jazn21sIcuugz6mJ2R4y6jFWTzwkNWy
IEBsQXdFCr67cdGGVWxhyvvSLKz0BjPGqvYTYTcRBooS04/dM0aSXhv+ZbQbX9Ar
gHFB4b3pqVh67WE7a2w8sH3sHVwZZbnwAxSI0Z82dzOmaXdNINIPNxBrtbkNB2Q2
Ep3SJ7JvSqHU3gaV6d4DFq0O+q6j9SkrDbatLFkHtA9iOYH4nRveYa+J4V3JZasH
j26rp3q2plSvkyfduBiUxsTf8lPmoEdbkbkLkX4m/uvOy+UmOfNfUrp31Ouad0Bg
7eHVvppi5J5SLuEef3dNOT84qtwNI9kdjSsDzYEePYyAwlrIUsIVEmYHuY1qhgrf
Yes3wj4phuPe1fB+ZFwxYVruZ6u4LyN0w+/TAkRbz9S3WijJ5MbYqzS+/SDeYvBv
z2w/QEevaOjMEfRM7+gLeF1iz9VDklxhIKQwzV9NMUF4Qz2aihvyxlhdsZtZu1AV
yKlupOI3NIXeRKHh/Mr7KPUYGDMftrQusLTHp10kH2exkFdTRoW6McEz2gDfUcPx
fxEazuum38K6s5apNcSkYVY/m5+VWMNBDkZJQN3RBdg=
`protect END_PROTECTED
