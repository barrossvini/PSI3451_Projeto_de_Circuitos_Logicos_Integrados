`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/CPFGEhJMjXn7TjRjfIVUUpAPuCwUFtUZuic2nvTe4Fcjva3YPrd1ilezz1Crab
iuqqzAkUA2hOAkw6sGJ3N145K8PtRUhuDlK4T3BowaYYb3mGVDW5vGGYV/oqi7TG
/eVWvB0y6qv5sWUibdrAhv2F+8B21M7u7/iIbD/I/Aq7/s7w74bJXp774tjTc/nH
gcInJIK/Uis1zS09unJYBMqDe1FDpDuPXvFWe4/Xl6+q0NEho1KeZiNy3VnisLrd
jj2yDq+omXOTwIgS5KuKiH92BMu2QYUriS09ijA2rGZ15WTnfeKaU62dB/TfTanf
cwk1FrfdFMzO2iPqIBKBUlWwAiI+ZWchcaTIiuTluB3n4Zwh/96SwzqnCdaTmbFP
uTZilxtf65j6pzhr7siZl19zFvER5KM3heQw2cu8AiddxBUcHRtAzc1AOBswv61R
1AKkSpQosOfsCTvYwAlYLC0TjUuGwh4WMe2guQhsU646lPdJkPG5JD5ud3WWZmVP
5+CAGkdQB9ljW6o2X9VCY0x0Z7yxgxYH2ZJ8vknYGYD9/sMvZpqGe2+9BGMqcx2a
CsA9pFL4oxIz6oP87z9Lf/xZhOoDe+e5XRz9iohrtpmS/csEEKeEmi9gHNDDS23D
0ovVGp3NXBYNKSY+CV6dxTkQY9tJH4FxOKRYuI4Dm22+jKPAWsNdQ3K2hVHgKeUM
cg6HcYEWZ1pEq21rmUH2KU2vaPcMK3k6zXFSjWbFIopk+ENnBHTZ7ffYqrygLGYN
H9Zi4q8YUOIKrTyeBo8q0aGJQlHriiXkv5EuEW2o6zlgn/uMuAQdP527a4UmMG/B
klOr/kY0K7XVqKQaj5ZBi2gTHNzSJNpG/6wqBMertrjPZx1YyAe+Y854ioS5rT1O
KrXxssucsVp0m1M95ccEQ4cDjSR5BMgxKP32cuIfTZBwjNF5LJd5FtglDA4Bt0gF
a6ktH8WsIl0/74rpRFSeWrrF+MY7iFBxzfaIv4cvR0aAegMp1dqopHpSmmUw1vd8
ThWE+YUjw767dBHc10QXGQQDTGVTz+KJm+OZeG/UvtvCOnBqYMEkwXtFxM/u67Lq
NxBWSiqwO3nc8JCFpRI5agcjlYixtRBQLLTLs56A3rBP7+DiqHhnRXcY+z0innwF
544iQNDLuQAlwXQqFS3ldP0l+Srvj1Q2t0rYduBbD0VQIRKuX72mnZ5PI93n/Rac
yoyvbr9XuKtitE3iXLwupUD+DdOpnU4+o/WOlAyq28YITluJJlkZMwMdtyAMOROj
GwaKIymtUxeTHLPm/0KSikLtEA5ZbCZnv9lM5huB5Dstfq7YuU3rlsLaA7a4GzBW
qun+ZZx7k8Vb/y62X6+uI72P4xSTNBMLO1yR8oNxOJCKoT4qE/4pp745IRu8ERzl
C2Fant7BikLKe/GNff1FCyzAjF727CQLFKG6nrDjQHa+a3m0Gv33Oq3fASQZChS+
YFImLNW9xNdU9uKhBlXI1bFJRfRK1vXRZ84FcDqAUZXyBk5D5uGmhouJHegW3+NN
WZfn+GD6eO05T2AChAsuqxIzzZfFLzjnVTGtzpWatqB63Dl9e04ugGyUEhHrAzy+
jKTZe3tm/oqggLwkqCfG8K7syROF9y+TyI44Nwyfgx+uO76pn2/fq+TLerAkaK96
4ZO8MPcG7ZJaJFR8ej1fBoxwSAuboAz4mhFPDuwpQSMOBMZTLIpPoZuLM7MmJnXx
U+DRAvXw/nGlB+HuhGDyoJ5Yj6AcKV9Oefh4xNg7YpZ4tIs9QOzfocm4KBHJwQKn
wPkHy4XM6aC7NhP0iYU+LKAIbmRA3F1UmqeJdvfNlBqZ356lxaRskahJ9X1rPD/h
qKYAKqljcSEU7iLh5AtGUIjYQnXtoHc2GuVeSeYgO33Jz6XbQEZuM3ZdUTrld7vX
qGGcimZcmYzyoYNMgHL9QKnKsN2xBXuMvdALb9qAtnsu9UlKqnsD1dbkmzxfxNex
O0UlRfZVmFT5tvbcxH7dD0VSy6ShIvRDh7RdbRsXf7gJTliYWi8bH8UQt2qJ+9fe
Flc/LCHOGpVf9FE5cjnYi6cNJcpOFfY8IXyYFgpmd5P6jht8dqCBzdWfcuQaRLCK
WdRCiD4iB3slvnLrX8SYamrZKzYLiOXG7oTeYZXm8amcOheDNLg8/Jcbj54VBqgu
QXCBP37JLZqeHxFJD/9uZ7nu97BHFreS8sfp5W91WrzToLLw263JwwvL1iutMtCd
D3U3gxY3tWIxce6jCAeUqM/stpe8fP8YDLzuBfKYojBKX3DXlCImdGo01Qi3+WC6
MIAv73gXzqFPu6/rqriF+Zim/5dhjv3sTXgOXzn3R2vdHmsv4Zp55caJNmoMTAUO
sCUO36Qz0E2r1M19opSmxqdUxC0Ls2gAYVKsZ+oYyyM+cSrJlgaN7P995z/QFVEO
HfD8GmN/ZRQZr/U8aYlskViLxY43lVfe5dgPbLPXNLJEIdiuc5iWZGpLuBVPVyKR
MfSVd5fvh9ATxZdmE627o102UtE61tOctquBuMQRIb6I7ZuT11DxFWSACHzfo3bP
d4hEBb0QmvGMoyUoE1mN6ewpXPVxWSq52gm3qpUbPrq9RAFh5sNnBY0oT7EZV81M
+Lc444bz7x2yBH/Vq8709epled37IvCVHrYMw1dvao//XWJouj22GDq0bHJwP6XS
Zlt3YP3AxVM5Wo8kZQoshQzMBlJIEcKIYXzWMh8kBJGmUP7z/DuTOn2CaHJzFlzS
RjL8qFZNg0AYqd3fZedFUpBxIPdlyRqFPCFwkVxerqtrnDxPOCFd1nDXrx192eLN
CK2z0QWODyWXMnRXay/Bddd2S0hgMec7NM1QOkXJ5Yw5+hP8Jg30aXVA4iSrGJ1D
M5VopvB47BkyslUFjRR2uhV820KH8ALutuq3OqAvTcJQAMPtubEo5PgABXPIunHO
5glEkPDYizyek0W68tjO6qcbyHgMSlcjJCjnFm1jg0/LxQyrT89hRPUOfDTCZhaW
/qSifoR31dyL+kPZ0x6DqaueVI1eNMteJB3IuLvruGI5WucE7yO0nZ4B3gA9I33/
9VPosemNTMu5sutUCYX8mOasaPIO0DtPkE50XlL9/mSQL1yjPcBcPvEEvK1zIpd+
Ud1TPzOS3ulip0Pajp+Q1Ka8fZDvorrW+zZ+pEysAFdM0c3mhsNJ0+pg8TnmBfNf
DqTUgAW3JhuaTzKHObzouBJANX8BAHxaK2jLUfbmDuscoB2FgILZjtKjrzbAhPXd
zBdnKstQMKk60O1cGv2YIR1kb4O5jVAwIaYhqBfDhNegxYqEz1SbrDdd01tbP9N6
qOSeRjXMi2HkTKUg55qMWaa/xa3OOugp0EbrpLcpIIskBwBBq2qzTJGAmBocypVI
iLHIzirdbtoMpWFO7jLKkCInZWM+PF1aIDxxOshOBsQWCxD6atG8ALPCvZsN9zPV
aEvc7nIafqMJcAQh4wm5lX4Zz55ilyfA3+hbY1+MvKDbQuXdzrMVMn5XEubA8DNi
GjXV5iER4c+HWy+F7RXJGKDs3111eUHRBY/Iat+nXBTltcnFvof8cdIZi4NlWBEq
AQC+1WSYy70DXoanuoyniX9zv+REqRepCb5Xvp4MjunL84xFxiatJjclC3GZV14k
8Mazq71fMa+woIn44azDHki9UeTDYwVJMmmgJPVs338346u6klw4eYghVcl/I1lx
4OV0Pumqnp/eX+1zCjl/s/CUWFXwjPeLpzJRO9yjuZAvgKK0vjRb8BsbZAsrjp33
ndxtgmNEbmCzAABlqnfddBW6PObXNdGeEWhV3+Uys1Ec5QcBU/WurRYcEFREHGID
bTATXIf0GArxeIdCIoaYDhLIPf7QEu1YHFya9bBhds8lPc0Ffn+dqqkVTSffl5/J
z/aAbCwad0Oq3wlcUvOAusY/cNx+peEqrQNiLMxnJ70tbhl90tt2Cqc6Hot7tQNL
3WzVsnevfaUMQ8hpX6IQ7arjszZ5fT8LcjFJj/afcFlaNH3kYPqzsS96tHXHTkRh
R/97K214TP5jYIMjXRmKKGVJ+dNo7Ubyj9hseDj4Vy6cxpmqIDZDX0Ne2a/i7T2c
kemRCPV9gaaytCWfKqy7WuXdsWUM7U1Ku91NfGK5FPVQb4aDV9T0FPxyg7Eb5ge8
ifMBV+uAuiymzyS/Izs/EdusfIu6xCnJkfmnM+5JtAinIdABU8salOf4QwllXt54
iHAHFGSUa96WzLd+NSOTDCu+qw3ZEWbpirX4ify5X+34rGHkUyUEK2hDS/K0ZoZ4
OPozHqrYXDFg6xdkTdP6L3Dgy2DEiahj0mEv9kBt4MzXrU1oC4S4IBGmlzO7GRP2
DVy/VaSrBPucQe8ZmmlOXM+DX1uXH8eRf9yq7c35DVrHgCsJnBZNoZIyK/fduWWR
rzRpAcdo+SbyPybc+9h5pjf5t0/fR1jv8rfsLOt9TgDL8x6vOLC5XOiBPFssgKN7
ORVGOGK1nLkRwqaTSUpcpamuPI1aBMoY3zySXfgdSmp0ab97bwNueCPXl90Ilh+C
gw40Q1O8xUtn8Oj6UeniwmqY1TadZUYudJBTn7XHCQNWnQcmaOao7w60JmndM4ki
lG+NW4pIm20c6U3upnnEvdo+tdOywuzqfC1TWLnk6GvRvBL+0iQ1AxIED6DByTxM
KJRN6cFkPNMnYCJcxfFwPdIumyELRM0xRG08/UBXF+Vhu7/7gWAMympDvNU88Rt/
iwg796JCpkcNqWaWOx2EA2/rIhCHWkWthXS3aZArZgMLoYyhemItdf8GdmqKROB/
zKwKT+/v2J/cggCScaVmiDUM2csolok3lhfRbhdhdiUvUKLy2CAKYGBusO4GiZnQ
kx8mHUeDLvbrKEwyg4Ej6u8iFQa2ckwhYL9pNd2E/7hwZsl+bMvJkV3NvIRgdQL6
wg10VujojMQXpL40jdvv4m7Jt56B+6cb2C5pJTs5gB0hJ381WQN5mSLp5m6/mYIN
rW+9Gs18e2hE1a35VLd8nRXbLJsYesTpHjySze7RnPVZySDG8PCaatzAWpIPa/sk
Kbz7tPvW8lll22W1a1gddisg58LThpa0ghoy9/qfR+DnaSWdbIE0BxQDYXXrqiHt
RHOPb9DKv7nLiVsax34T/LsNzc8W5eRjiXcHsyJRupnQu2HOVn4KF1BIVhRLD/OH
60f+b6XGSJC79KQDn0Rh3IznSQ65H+FX2Cli0EpqqAiuVWhZ/aSNDVPHDtg6SX/a
Nxlzw9+8jOZ+H4LTLSJb3uMNQ7YDtYSxMR6U3w4UoJHSeMH2MEU6QNoWgbkHKuXN
nkmVVGdRmkFUOMIX34vgqCwxji2GUoIXlyMJAAMXGkGAmcQ5FmiCNLcqOlaV0sBZ
I56iFPioIOwU2rPkQ7tZfE3Exq6UX+ic5LMniQLXYthq6/SMzHv3TCN+IScbuwMg
Dm66sZqCUIgZKeL6Tw4hcdkatsxDJM2bLhFaXrMUNapGZHTvry/HIKXdS/Dlsqn/
22DKptqI+6sNoClpGEp4UvkT7HgjkhlUcPmd6bgmYJkTlhAwohmXJqfGX5th//pf
/MiVTKjTbe7BFgZI0k7vdBEsfKxYGlxGXnQBMblCWaXBcab3ZcAL3Z4n6EsFgbse
bYFvqdvh12s6pHCp0u5lgvk6/NtZzAFWE1k4YoQXGRi4RdGxuPih4R1iqbH7ovLK
DKWpSj0lHwZn2OTxYI8BHuMb5lrKwhJOemv5RcP/R5Kudp6wNbzVkWld8f1SjP3A
IZTVFUcZmpfvOwShvfI3RQxouviNjVjF7b61t4rgPg2UJlH5zeQH3vTYV78d/0Bn
oMIwpF0HAwZeGOTRAIalt3q6r2m9xctyaw+ypxD0j3QcnHbYbb+VmMqGxJn7ZcVi
zFuILra+jukFH3Ty6QsxzAPod3aLTtpn0bDwtlExcMDSp15rtrEBFXjTMnXhF8xt
5II5BkX+CxUFAtfNPjMUDYNYhoQCsqEbLfLBGnQTG3gT5POc+W/kibriawxDFXmb
P2urrkp0RxMkj8+g4tV3NQIWC+UbRooeygRr5MX+qKUjmGcyQcGevu8iMgbQgLDI
fkD+Ihihl/n+ii1RiEoXkJnQ3wnmyciejt9zFfqe71e9hsWS6kvneBURdhNdA4+q
Y11u+cjHHG/sYBrdFxt69A==
`protect END_PROTECTED
