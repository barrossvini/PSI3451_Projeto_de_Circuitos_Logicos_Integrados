`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16hc9nIZP4OPu2wCBd0XNJKfjpFWW4hG69xWE9GuvzY3D11AZy+Y7HWpcAPwKYIY
NhRA63mTv25QfJiyr9BuimnfmqilcNGU1I5BVgOJmIJy4qCgXCm+cHGdomCtTBdf
KgSpJ8EdKvbz6uBbSmxPajllbo4Lg+e6zyYEKFtJcc1g4YhmPDrMcd1WIZ7Y5x9s
fLNz5dXuDYhj2oxj0EUZiuiK70XTuJ73fd5EIylb/krWZd0/IHgP0DYwjOipgOJD
F15YgkCwi/pC2bg7i+yiSr7fVCEXhEyKykOFl9PI1ulQlNNe4jlJvq8JHZpTvhvX
VJ5Nx8EnOFoQHM916IUXeYw7z3FT2pQKtKcL26lNzA3cq5qADPP9aTaIcyIJjd2K
ZwgNtV4kgf+hR2aIQor9HBR9sCWntn2OMN2WqpYjR02NkCcJFgvP5RoPRftsKTRM
5lPmj4XoYOOtUi0N78Y99t4jgOe9vCEoeowQp1BHH5VFTSTpcmMW9sP1Pu58xNy/
0lAEC26mqwpOjlirtH1JLGN6kEfSVU3CZLn06up+WgahNRAHpbcP+tPv42RESrt6
CRm76NkGbo6jOr4mxrrBbEddXc+mT2iUiK8OEFoZyltjTUtOsehc6czeU+sqXDBv
8rxGvt2aDIcr8HOLZH6AbTmBhy8M7b9fmg7dbuO78KQqr/4nDpoD2fmXBVCwke6+
cxn0Zy11T018Pr1k4lDg/WZVLpelYmETEaAZnXbr6p58LxcfQTpt5T09TzxwOnzq
WoXELwXKusU4k6HaIRSirgf140BaRCLsn1QtliXaw7CTspc72Xx32wN126h3zHLw
aWFpyCkc920pJZtdZBmQWgGZGvzG4yXrOYMawh3prQA=
`protect END_PROTECTED
