`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yJzHr/HLvOJzK9w4S9mE2wjefrc/zTiXHxwYNUO8Ur2zvkJ4DHyGJ+OHmWfPNseo
W4fcB1/XhWTu5SB3kSXc+PuIvuln1OLIudzJeqgMc9j7WwC08emeLdZXRgptQUOf
JZwRQcvz31Ge4moPGp3pu5Hpym56EAmzNLDNI61URElFzTHp6mgCkZDyfCVKxc88
Ba5BbxSp2Cn1ML3G7PGOkDPdV/72xeAVSV2TH0xqbuuDHYeCdb86FZeaKJG9oJne
A++FmhmS0fGkH5/2OftvXgvhnnNnhkqTrNfR54IMF1hzaLaIAkK0TBawIZtF+ajc
qO/8Dp9qi/pJMIrz6F+dUUEuKSJYo+Uv7FUKpiSLDtpkOgP2UajayUNNQHDtECgr
75DuarSl+FVxdfVCfRAJhxkwMBqgGgmVgNf+RxqLSQvxnNC/ZhnqcBX/SziXK8xl
VT/F9W1h/4rFUsou6B+j2Rfx/fz/vuWnd0o85NOFQ802FP8nK6aVJrdDhZwWUII1
qrpmzBBUm3nVCu3f1xNo+fo3ZvhmpjdbgnXcWxhX5dFbDWv1qtHcPWiGEH1u2IFl
igClRcWTYID9bBnS12e3k+I/06no3UYvGMcJnkVjkckNcr+iJ9Ccg8Nge7AxGBM2
V65ElXAWJpeQ3AMlPFa5rKVZ1avyPxN/EolSSPdwWTC7Ykq+qPLvt7X00XeWpqVI
93fj7xJp8M74F9LRsO0cwB2J9CeAeOLSdWo9mFYcf16nCvsAl1yE+1frdGvwADrk
JtQSv/eg7h8DBH7fezkpppdaDJ3hPJ07ALIxAENusk/R/wbp/7luP1iQ3jOtqUsj
s0eyj7pCZR2Tcbia6EF4HqU5jJqBzN/rLv1wy2CvS2TMN3AgQNOltzSXQEuUSFIA
KG4k0bhLEX+6jqiOFJwrz283jgeWHLMUT9gJoOnwqBjCa8L3I3VlU5fll40gC76d
quOmauiNutjA77dQaZdIiILNaTH9i0Fkp+FeS4ZJ3RjF2882YX0PYa1ouzGEUT+o
En5BJLGzCiCs6qvPy8KjB80L58V7wQxDgbNGbvTI6+aS0dkAUq4bnZ0Ug+mKPTJw
45DsEkOraIgJjxO7jrUJZw==
`protect END_PROTECTED
