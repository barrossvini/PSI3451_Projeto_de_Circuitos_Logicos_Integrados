`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sI7dZ4Gj/Cbb+8Sp87cXbwzHpqq769LmLthl0ZQ1/0CYnhZlvtbozUu2GhgNJRrN
VE9Vafkuwb5m+ybd0cp9CLNf7UeCaAisZVXYgrJnzIPgFbRgdMiynVkjDQv3Gza/
T8XeJJ1lqN3ZLRUiNas+Fi6SKKMuZRMXAWUdnP1XlEw0L2sLsYGQsT7p6Vpu+a1d
KiCF4YJa+dgfiyg67EqevQh3Yhb/SUf05iYMWuexLDFmNozx9WpvZcqJr56RmSla
qvd6tK9KrNK6no5Q6taqBZW/tEOpUExjieWbPgfM65GXY65VlJUue4vq0GfCixU1
EwK3EYwM2lvRrSLnSWDH3XWnn2aApe+19dfn6ZgVweZlrJyMIa9ly3GLmx4E3gts
ctwLcWoRD2UD0NxAXbBWAp6No72ZbOKXTSdkmE2WRcrQRfLXSNrZ2tRRv1J42WMP
Tao5hToq8bwz8OHN6Dcdvbl0UuhWzOndADSdLlYi2E9VM6EVO66tuk05NrRjw/Hi
EWh9FuzMG+yeWlpdgO8w5Hc7xMwngeLjkJ6oLsuif5VKrXZIAtkHKd6C9ZGMvpHs
QEmkRNWXJzczOVHTs83kysi+/Oq5XlqfxbRFrcSG4js8DQyCzNx6bFDRc37/UT69
iSUK8PnMFC216Q+c5RSsMNtrYsSjixfDWG6f2vKXMweL4oR448YK1OZzLxCNpxqX
chR/0HDig3Z85josgwmCiNmdKOhQNiOQR1InqqFxBWKcoAtNQD1fw/xUIRxIxOov
UcfikiywUrjHlungCmC2K+X7yL291abfz0LlE/CZuaAKMvt8faEM9ThuufZg5eEv
IpC5+z456uDJ+tvi+FUNM/4LSuzcAkyXxu/Shq5qb8drGCaOQfjvVsgFxrvcJg7O
xPqV8cfTG5nh1LqBhqDlHZqMT0vF/oToEObSbILSPsxnrdinNRTzTalqXQIv89+o
QaLa4hTGZXoJm66VtbezBy1jsGFS6MOIu19HnPpmgIVa/ewCCelT9bZGPoHIYzOG
V9bFXNUM7jHBPTWRh2eTs0cRTZRhK0HF+03595DnvoHR8/yaFXj+xV7HmDdzgjNJ
JKIgD3ws+K1rTLnbALLoTs7ebQ8xRP8auxo5IQoYIbwLcWPA7q9rWVDo6xUaYIja
g4hcRsgQ41iplFSKGHd/ApdzIBTBUnH0iCRpVwuKNrQyap5hO2bQSpUvx9YJm2qL
CTUHXbI+wVsJRL/M4h1fDScf70ea7aklP8jhUBWltcvDFSCDkgsON9i1ZKzLnjX1
IoTMPdVCF11v5Y7rB5mDup5Sf9zd2hgZmlhJO4xiK2/E0CLOq/cCqDtwItbzcMQi
oQFxTeTeao4nKiSZar7CvhhgqO7tra84cTzwwuwzU+WApoZYJ8la9kBVsbTstR1e
A5zE2eCMQ8MS79ADM5Zhhp+0V7ngO8INEuL1bf12Kdjk8tMemHfEQzZ8E3RsMGLr
hl2zr0bXXRG4ApFBdIZ05A0qv+FS9oSbWJuKPJdAG2ceuiAdBRKi5gAbMJGMAZZ0
rFXOpvxCxnxYpE2Bbd8zZfh4KT5uf0pXh+Czc2l9t2o3hBuNEVxwI5VNn4yCyayx
tV0iFsmmgFMV1j7GH9pAPL1t39+zTw8E8UdmOd2fj8ts3nRcfbOGFbJFD3GpFekq
2vnbopkA+VRP1/O87oDhZYqCNf+HKcHo2jG7l4m/TbyMxLptX6nyC238cxo0j4ZC
qSK0fyCYHBJfxPrsLP0MlomOLMrHPRC4x+RMMhIxBKM=
`protect END_PROTECTED
