`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3nZcNq7Vx4HBa/vILG3a30pJpYO6QPnE74r40qXePiH3yGLeX0H95qpbyd9bijQf
Z8tgTwX5rJvnAzoQH2mjz6e6QSCub6v0nKUe4Zo1wTLZAjuJfBotnnO5lwjaetHd
3XUGCl6Vv7C5dUzIOSxE/6JuquZkNBpHHjQU56pI/2Wy27GZXtRMKH6FQmp7AiW1
uRl/WeoWbQLVueRjez+rn/boeQGwTmCs18v4Gs5dj8UGuH7tHSlfAEZXVu93LOa6
1Z5DYF2SChz3hspz1bSkyd6s0i08I1hkg/CQbIlRrm9lvJEoL16TXsqyx/llbW+m
vq/dJojHTJmu+iHLDtAxpHlc6ytDjCo2aWHjAI2z9K5m9y9R9/NYwQkyc03OkYNI
QOO8ZUFEOsUAfbqyEc3VipeQJAzL9fRYJDyiz+TEOH2qHL5dm/RSU8NcmWhJSdsV
iCqn2O2oTz35ERTpeREzL77u8aKQsD2FRvz9hyBhmTpKegIfKRXl8qeuXl6kWOEC
J+6jKn9Pok+V25ga/aW/o197eSs4M3YlaBr7J3tLSpo4dW2wF8yuCeOJsZgbImG7
u9eLPGveLayWR7cvwfchA3vNHYPHngYrMAac+QIusfRL/I1iPfphhKYvTBCZ4Rtv
y6WUeDqcLc9NGvNjgVO/MF7f8Ruq6BZiDRCFfuDiuhcUdHe8fzl2/6OSLHZenaj8
4cU8R57K23h9CiQuyeNqczB/BKOaLbLmUY6et8O0+71DNKvOzC9k6qZIVLmiFL5q
qY7E1sU0A/ZZIIhiaA11obMuXuQ55ipJMiPXHbql3vBcQENiYK5gnK3vhbl8Ecx2
tUeXs6qbQLX9p+X4kLLYotY9v1MfLAWphCJ6MqbBHbiSRPmD8hVyDTIGAl180VoR
`protect END_PROTECTED
