`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U68jT//ffeYAe2srJv3mMN8GKD/6NwpmT1XxrH9cHxv/BAdNPhjH/Cu0FESe+xn4
og2WYZQtmZXdfv3DcKwTOnDWv5Wk+H6GjNLFjF8UA7fgmNru7hVbWCJdZ3dRYFL4
Aa6IBl7FHvGPSf986eUQPDyzx1hS2rOtNwbuWoYmP8yLwjJJgpl7MdkCg85hLgDc
4W75uRo3BX5CwyrZbvr+TKADD9rxsRaE2gtV6kmRB9rtrsS9Q5NOaHaLWO0u5taQ
uPWKZwj8NyhnT/ekeNInEysqdmoScql4yVp3XkOL1viyugL9A6sIm3iZmKreB2lR
zjH2BS5fAQPgmjh+qr4eICxZHJ5zf+liVwhL6M5wd42mPGXCIknI1lzEIZ/ngVsJ
7fn47knDcciAfd39NOnXqDOPMBy8Zc/FtQjqsJp2fWSw4EyP7DtLqNE4kbmhx7C4
k5yxV3ZysKINl3HiK/bWdpabRf0hhwSh9RUCprB1bVOId3lEglPEbFpHTFHqLHW/
ztocsY+xnuWvvkRdtTe0l187QuMDAwSHTzY+H/690S7+XEIS/A6IhOGiuLbHXoSM
yfrHi7xA9tCf+045qrKRx7iyGbbubx4RyypB/+H2KtavstwYAwxkfatIEMDpdFPX
5N66NIPeAZkID6/fuON5d720P3QBTCAcRLNUzaXclxSKaForPHYLQYvj/+3KPEfv
ieLsS5FXwWPZ9j1Pk+egSr4n7se69mEfTPhh8VWVYzkctNF/R0pCLYPHT60N71Ku
MYk93cerImWvMu2jBJ4ojIJxyhZA965xNAqtKYeok3gSi8nxkfxGaJAfeHnkQSlP
aU+RRAMzOWs9EYyX38mJPpuJZNT4DVzd5t7eigKJ/isYbq6aPLabSwU1u+q/JOtI
xUnf56kMYUmMdP1c0lIA0Wjox3EvVTxv8WhoRunhIwnGA3LHgn7FDymYRXsz0RFl
h3kirxkeOJ2SV3b4V1CWWX/4FjVojaxJGjN8EF6WNJG86FKsb4odLbqfaSsMr3XI
QVDuKqKSpuvoSYoj7sfsSXm5+lvJKjwGan296xRctJkv/JooN+gg1WXUHE0voSYc
x6GHNf0FccTEwUf98ULl3JuTWFn/0hoSywHCPLghU6qXCAa5R2zOLD7MixSmM4XZ
6h+Tz7FZ6xvl1cVHgARKB8E2VSj8Ef5PHbxNXu8wFqePVpsE5R5iq6BKKRpUAPHq
xEb6plfpzP+8VmcT7MBJj2/EbVa4YzjdKiklnhFNb54=
`protect END_PROTECTED
