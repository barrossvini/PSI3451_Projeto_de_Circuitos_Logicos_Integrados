`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RziToDceQw635viBWtk3FroP4NAmpOH8cVtlvDuAU5uRVgBXZ6gdIaQzhlNs5xJ8
sez8o/ZIyehHyNLNVY3tWv16ieqCzuuusqKu4DutNVItB57D9NTl3xKCnE/T3jQX
J22eJR1/Cf0wrBJafnoi10eDc/jN+vLhhFrFVqsOeTk7lqXRhfhjMZHXUab3ftwY
mZ3YMFKC/hrpRbaoW0iFWbMWNcgAVcKZzQfhkltTD6dkTj2UwH8n8xACpSuMAcFD
rV4deYE3EZ6MUc3bABoEewfiTDFgCtxzuLXfVSChKlgPqPYqa7/fvxSL0EI0t5My
cWmMzq8yK+4d6ZRP2Tx087MyWtRIl5k9bYCP5p6w8aLEzWIAk80/GL1BQbGgf5f+
KEW8wVisBjK76EIn8wJ+RiICKfHmf1gT0LdhVdT28u2+w1rc2pMIPIzsaW6dMHbp
uxDep9p1MHUcqGK73EHPkj0X+Mi5p9LimLAwdyxR0cTOvFp0VhiZmEsWSnX7RrwK
eixi4aDZUNq3cJtRV/KAq2Eu+2dtIr50pYcCfQ6yUDylHsokjpPLda996MYrhIRM
l+HNtVRTUzTdgPS8ZB5sWyOoUHOrKJNeuPOrpkEQSpmTRpU4NfIMBhBbe0hwEaDY
F0xBgp6Mqdy1RNA4hazBhm7vmTl/pi7SuHnJETrW9iF1Tu3atX9oyeoIKkmMGZZc
rVzXEyzFOKkfjRX0gBdWxNbF7F6poN+h0i0tD5+fVaeMStQIId6QncqPfJMxMZAs
Ci420svGHKR8AQ/RUAxWervbRPak9nFDfAbLjwH6j7/cFOfYKCLIX9VtdhN1E6jv
f4+5XmnnLMa/xKx4xulIoJdTaDOx0dtkE2wcq6Ff4ts/YGX2hxKhK2ecc0NPCRu9
4FyVXRTK83+yTxlbdOUHT0WwLRNNCL4YAIsKBdDz1ZtIZ2DwAckUFPeVl0f1B+GB
SGwKdQH/YskVikph5VaSlsWkRCkClSJ2QgskSphxtOq+HaBk77YI0n/Pv3dccDIM
XobpvR9UKe2JlS9ZiH8NEDbAbNSNpD7zfseOVg+E4qCLd1SyKtP2wEAfyZBI70Um
aLgp0yfvKLsOct2hydzkUmeCPoPQkg+WCvJAaEs+7lnd7L/KykkRty67DDSoOER3
nvvPIqUQZtXkpegbl/oLQgq0/NEb0t+FHlu0jF3e/3zD0E/8XiFFNy3kW4B9zgVr
q2YtLRlr24hnS3EsPmAsDhfloctFDYvxJfwUv6QikUA=
`protect END_PROTECTED
