`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tk381sPybVHfdsS0hxbAqUg9wJSC30khvabfWHjHqET8prbzIEuVc1wjpC+82AyL
s5HvcBn7N44jaP6RaS6FhSbANOfby7qAyB4VQqDm1Y8Sh40UVP91cvNg6LMHK/ee
LruaINwUw93XPOtS5FjTTXBGnbGX/F0nldPOytyJViOyaHgv6I4cpE3s3zjQ8Fdy
OjmeA+UgR8YpZaS1Qx/Pa/NAMzFU0rVJu2zJylPwH9oOOV6jVlRah4M91T8cI02z
+gLisE4G+yUO6bzG9fpsbu4scEBzJ2PrJoYZjdVgl8cytFxyve4KJlccjzJsf9se
FBfdh53HlRRT/Osl93K96aqBjy4fN5SsFEGULki7Kqymgez70qTs7G3VKr8js/2o
wBrl3NUCbKV9AN/3Da18jBysJqPuvy6ELH3NctjFxQ6OmMQNmURYjXZWuosjgtXC
Vvu855gbaLeP3UsJABepusC+px4qJTcHwmBSJIQ0Wc+e7YK/zUUXc/wN0JSsuujp
y2VvrVzN3iA6ZxtatJioIPXCnbQ14gldojofT583o/LP7WcrYB4onqaZ3y2wJN3P
ZauUw1WgVjvPeR09A9MS9UEI1NJc3RAKgsSYGgt3R/6Avw5yVsd10jxwcVUbk7fh
nnzTPp/8Z/z4vAiO7TNfQqSjNboZndl0XlsiYUV3FvsiC5x6SmAm+UsV/6aLWVLj
6QUtD1ZycFRQD8xAVqQ33Y7+ngSja53QXubVQ0oczb4WOf6cAZ/RSUao2xyXCT3+
/mQEbs2t3BRaGIzskWQDvA==
`protect END_PROTECTED
