`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iMMyKi9V/OBraPICe4+cXzKZ5jpolUl50/40DGvlQaRR0P3YfcG1wsuNzMdHKZjR
weg/5Rmu/2bwz9yWKrh7mwnn/FjXkOxs1o6JdAZrfKbKpgxFgN9DUgInjU2uhkmD
poHDg7E2AjkvbjuPYdfylqvopQ1xXLOvXVJk1J1Rbp5+dbR2/o3EkYxu5PO8GpiO
pN1IDl6jzcFfyRSG5LqXyNpuzxVY0DrovqqUrwlgZaMXSIYP7hKzDSBW8Hd8f81U
Wf9dvvkv7eWzkghHGaXBC9sNT/REDLUk8aDwkV3vZwpTUgSyBoCpCxcBOJDy+Id9
NUENglH6VFLQNftX0oIHXBnZQS5SE7b39vSjzauO9W/8w9wqAZ24uIvV8h3dpDrL
V1sRrqYWdr4r17vmH2uyMKWrXNPuHKA4ehsi0vhjc5TkEunwRMbMd/YVxxJ3/qe4
CpVqgxZnsWJB2VRefT1dsF9nz3Pap6ZBgvCafaFYHuONvGQ2WCSd5QmeZaDMbX/7
uzsbhEnenitbc03e17kuy+/rdPPs+IbhD24IN65rd7IUG6yIY0awrXvl6Ld2FIxS
R5oIkDd0pDVVRDr4XcmAaiB1twFRuKgE/01V5OQpvIToQDoNW38dlMVk49+Rzg9W
c58rPoybCfwMgiVNvcP6/GU1Gu9p9bUpPBcvbul5UjOpYhjFbdNorux818V6iSd/
7+pdZbd+X7h1xKkc1dpOvY89Ag8jR3zoEBl2hDs3S62/A+/u7NxThyoGclFz3xex
apircqfQmKwixPoWxy0lPTlHX588xCHn39kxU5rsb0T7eMOmdgklsE+yFMPqlGAD
ciOcd3rwaQMxMhHPztxmseV8H2Wz2s6HJMaOzqfmksrOTfmsnt0F040LEPg3nYVp
tcu1LaOh1TMg7V+NhRvDHhgkLlQhVcElQNlg4wUquBgwbFrSfbTKAP2Df+KZIBYs
c6rbnJgb9LfgAriPKVm3EmybW7lL8Kwf+dtUYmjE82lFi3+8w6FJ4c09lTBzhzoi
kPRjklnSSarZcevvjM5vmzC6xN1b8Cn6gHhEWHY/AvoVIUdgpy4YZHpN+a1omhy0
0+pphg3m7du0vAir0zLZGNbv7bqs1KK1bMcwcKuJMlO/oTdAXaC19x9+cg+Vep5R
kCFL634dLZFW9gdPxDVYRJc3QJsW7h2L0/JkiMUl6cpOhr4burQlT7NoiaILWXHv
EkT74JibYMLpgjw0Fvri0SNyBCkQcJb/h1AFfj+MvPBHmrjPHEjiy2ZZUYEuwWwW
mYGgaZgFLNqkXReezRbjO0UHy6ab00FpSM90xRXn/nKZKnNoJpNpGLV7cfNmGxCN
cy1epyDQBbPn64VICfkunc5GV5zuzrN9XiLR4q74zG1rL9dmko9/jcHonuDUxHnQ
kBwUZo2EwinDOyArKWNb6GE1oQyC5ABSR7q+ffOcdvoXpveqVgbIUoQRKJa0lh3a
`protect END_PROTECTED
