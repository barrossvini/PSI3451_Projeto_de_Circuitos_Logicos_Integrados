`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2XIOBtzL/5wbXSp9COKpP1wIPu58H1GLR2m4DKn5utH1rCEp2I6rOhBLOtZlM837
I2y1wxhKHAw2K7vmXS/KxPvhBSX+yERCfK144hQWHQfz14ilDaupP+l84UHDxCTy
+Gia60LRhdH7wCNh97luBgVdAvE87qaMljz6MDNv8zXideVMLNe3hNePSjQOh+HE
tqX7L2hb5/6qfVXB5CeIPPFRmU68lmzi/3ywbD2bynM+E1k2ubJ0Ij0/EaYCKWX8
PRd3/b088stbtFS704lcZuBn4NiD08mugbZE7vvCwcG1/sjQq8uZVIIVf5pno1Rm
K8dxKSFCr/RhKoZsPWm7jxetPMOnSMzjc1t66GkW2kVjTJZpyAh3DsUUedNQNa8x
LkZdR/gthBs9AmXf5zx6/BiI7RpOWft1hypUdpddXrLGw7hgr7K8lgGBVARFuvQ4
0APbl6PsoHDGexoR4BaddorgZaMqHu3yJCH5V9KEnroIJRUkjO7wtWgD7FJaWZMO
OfDkOT0nBsFJqPBDL+pIHzVZ0fQUd01Oozhh77TloR/4Nge7hnYQwMYrfSibYU7i
TvNBanJChmE16AwMVnnEXYxc0vhpJQ2x9ejrvpnYIVKrNReERY5n2krByzkNifWm
`protect END_PROTECTED
