`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFeMl/jyRxjQhFAuM7iMYqiR5ijl/lsCjSaNlIPSmXUyD8bnNMsWtefkZynjCoke
5oTCf3M/fMLYWKTneceRTq3zIsbSmHDgQ3slFzLfy9MblKdSzDlPPzT6uT4VyviT
hopmroxhCh+TN+aiiL57K6P5va0o5dPSXgcGpXl5c25XH2xds7e2aGVMjijT94Kp
RT/3xdaHZ6hHBqWT46AuJO478AtYpapp4vJuhicaSGL3S9zmMsmJWezY+nRITPrn
R4r3Wlz8kSS9S1+BKVNPs7oqjHEtYQaaidStLOLrN7Z2ZcMe1t+rZwXFEjWRKEbc
Bd9m4YocAuKWxvx8+cBx0HJ8HIM9BBjDoL9toysjES2e1I13brT38WI+pHPLZtDR
GYQBdtWrRog9/y/fQ/Lsh+7u/lijYlbp+7qcvgp0NLXN9dmpiNcqVEt5Q8fah6FU
azrSOso3Bs+KGgp3ls5arLvDe7nVXid2GV8+jJTI7ZX9PYD1p9VyAZWH4ks2ntYS
y5HC6XuGSAxDCQFFqF+5wDrjwm7WT1MC5ddoaKiRDu636XpWAfxlJobUv/0P79hE
b2de1WPxuHNeq8kutHhPuPrSXF41o2mLyDRTLd9O2DjIkvneLdXJjqQLbXh6IY1m
spEMO0RRMh1pPb20AVNPY1VYuHLtWSghCc1c5hXgHTyOqXsHe1YIA9DXdquX7WRe
b5k7ILvKcRKDlXauAjK2IB+kD4z+rlHtQ54OVTv6QCF6YpAVtrueeJ+pOyxkX2S/
mKAv8bQd3sQS5hvyc4yBMme4jfTQOJpbeoxhWN0+KwSwHrR6bt66t2Gculs1HQ3y
aDf5e3KrYLoI0RbK2ccaUU+qo8OB97oHFjvoTHCPInhiBRVOaJHrc6ahoSk1hOJK
f/xfS2+i5rKjKp4VZof9ZTeuE6ggAfhiGoxS3pRiFca6qgSiKkued2bIdLm4PiGM
gdQlAGmRY6ZRkUsPPPoIlaAHwOT19ZgGPap0Gcws6jxRK0n/Jm+Pt8KC6Un3/Bu8
taH4ZdJRhfVQdCDIDRcLUsN9zwec9BkVMBj+WvwEKcuvrAbBOS0TvBAc2qG/oOL6
6c/fHpyX54jzpXj8UbuKWinZx37l5Jb9Fr/16o9NyHF2jwOkMj6x3ENqh4D2W4MP
s0WW6Eersfrv4Zx21/Q7X7acUaCAHCsp/16eVXCOjKhaxYysAaMjr9C8zNPtGhFb
M7DONnXsT6SDobVcYDbSxFp087HdmOxpL/ZzJPxPR/xOmtIYJNycqWVFBMCoYYZW
h+ztVLEr8cDZtHUX1Q7t+A/0qMvXfPYmQjj3Kk3iCoyHztXYIog+PTV17Vl1HO5K
7vO5vsXwgLKKLOxzWNN2/mANFofiKSk+tXs6U9pKMKr+lcsC3LBkOV4/lKilPbgN
Z3LwCcbAAQ1xfZNGKiUOMf86g8eMf5CqYdzTvYBMsuoC+d0el9tstBax/Ha934+O
gH9/n2HEE5YfFkkuBgLrnmQth/lyE0c7Bry+QTWCBPe7CF45DpXINermJpVlC/GY
iO5Cqnl9oQZYzqvPdGSzdhx4c0SO5yEgqOTFGua36mHN6Eqefu5Xwb+q4a2Mc96R
Zx/UssdS23w4xFNn47LUgNIo1vt86eyzrOe+wSDVv0z4SNsecTPjd0n4m4ZdbS3n
88/g74tcoP2ULc0BpgldSW12nQC5pWDfsEX59XVsEZ3pg/C7z3H0+0dBPh2gyk+4
ukkDzFugCajIkEztR6QJWA==
`protect END_PROTECTED
