`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/nPbN4fmtKFae26zYT1vPNd/zDAMOkA/bvq2FI9FWJFeDqG4ux0enEIZupQC9Qpd
ZHSw9DuWUR/P+pQsIoicqnmbhnsQEw/pv45iCAsWNIeRIp96yHX0RZa9/5B+cXoG
/hfH3E5YR/scWwM2eUvX2R22jCNBbDu/2dFmxPzo5/PMJjAGSAsmcddhpRtxQcG6
VIZ60k2x0HoOur9/Y1qoKMXcKh2k61ha4p6D8LTQFAcwQyDL5k45FKkBHwzUlwqj
s8gGv7fSrlF9iLHNkl5rs2pJx7S0B1Q61ogI62WA7BJ+pKsYIVx2yK+nfD/emqO7
HowE3P9AV8etuuXDOVnbvAn1xLO0THfygbs8pvmDzgh03OrM7SXbj2qdvoCVx3OL
HHvBODZkLgczyiUGKqvPNBVtU2nprIlp3Wed4dKbCjEyyZQSgqPOhENHNWriTOq8
SbQLCCttpsiJWE5UtupbrqH+dIvXuletri5fyeZ7HIs3nhFDDeeg+ViGgJ2lMrXo
QIouGBiih361m5lXdjgpittLEmlqHpCmICYrTP6XtBXxGNxz6KQdNdNop01kK13c
4RBmM0GyjWIQI/U/wOXJ/uHt90v2lsdqhze5Bna2GODvcK+LqFBHJ+IThO1jS0TK
z7A1Xwq/g1zSE2sJpof1HDoONhiHlqzVZC4BQ6y0q9qEu2cMMhghai0uenkI+brx
h+jl1ge+NaNKfI/GW9NlfNmpA0UG/ZdclhaStzVh6NaXpe8CV/No/RDTLI+l5+zO
9+6H90dXnGGEPw9DeFmtPqw7HG2NOnMxjdR7E7PHLGdd0DsdQhMTKsdoBvyzXG/N
eNSrFWu2YKZTrlDzz9zEzv112tNG1XjH90tLJk7IHgsFpBKvaEKzYbC7t1TAI+jK
f/iwmmBjjuOnluIgy2A8QqlCk0A0pQU0lpDeCZaCavKnJOOg6zTmMkC3oqT1adzE
oDtpiio9ewpsVv9lBUFeh/whLheNUYPT+yFQk9Eh3XbF68EKq6J3Ln4HoRepgSkG
NcXbaqcf+LTobF1sPVk3eOkw18/TI65iqkz5+V2UZo3GT56xplP4FSoQnNo2E06z
EJh3geK+fe4vUZs03E90Rej4Ew7xZUq5t1VsgSpfA8vO+zxAUy0wA6mMGFMJLlYM
P9YeSzZ7VykUf3uEB2w9MReCxGJtM3UnVYfVTh6xIuS/5JesHpL71XHTw5lGbNu3
o2Zk8c0X5xK9gltLaZgrgkFo2yLGfy8c6lzid+x2AAf7B4ZbYTtxNhsf7EoaamIT
J+Nyc1m4MihuHXz9OB43J+L33mTsVZmzzMEYWtarK0caHYJayBnPwrDdVUcsOM19
CQ0OTH9z8LFmEksicZXCudEcMiaA9h/Lp3nVP2FT5wDrrdLsEBRIcBPD22m7Bp2c
1bwNdrseALNe0YN/cABXjLY+J/APxLJjI/TyMe7FQerQTJlv/pvipHjSyWKZHRll
yzd8qSrCz9qNw6OAlwmSBxV1KxTDswm2PajBIGWmCyMvCyIDykaWbjxuq7a70j22
Am6ss8yztv7VFrnx4MdomCmpcGVYky13exwiJBt4PpYvzzixzZVQYj3lHnmaHuJy
50rICzJJdge90et6tuXBo6RC36B5r2bon97+wqW/ifA73x1KP1KF3r4Po3WR/qnX
7rq14/n0CCBJp+08djfvEY2s1ESfUA4iRaPqwCCr6tq4i0PtS3anQ6ZghE0evnUB
q40I/Xyw9EQjDlP8WPC5UdZwpUDVpcs4U+LFLUY7E1S9A5nz8WbyicmjbDKu2iV/
Pcm2kVpvGZUdp8oArjpQKCv02jFNAMwHcGCcNibGoCZ7bU7HKfk5xLW4nePU5BYx
/U+PndaBTefP5qmOkWjP+uk6/vqFTmyBkPKTfGb6PZrGo0gHoXBmHFOlNvjcmfd4
5hAokFjIfQjoP0DOVgeUwrUZ7bBriFWP+G9DQDRKS4v5zKlmEzY2GMtjmGsA5PpB
hLGtj6eWcZbYOcE6eq9vbWfNums35ge5ImNpJQrCkZvRaQUSQzVZLWdNP2An3vm1
R8Tl4n7t18EVdGa4rGvvC1Av1mZzKYoGqrq7ZBCdag3PhITE6FbCZlboO/Pnc6j6
MJvKNmgO9nuRIfmqE34KYphrm3WMUcOylIFWqhhch8lgUyj1RVaZw9RnzVtR/U6x
g58Gz8cMoNT+KhM3EIYzdTcQoPx4t3xSCAzGRVXmhnJoKCWNvmklff0AjHRomEyE
ikcWuL13wdTeUCx6uFd+JXzXj62v02ntNUhhWVgRGusQqky2yS/qyTY64V0H44Vk
x40/IJ4BmUfRH9iRPYRJSSAmw8WBk3BFelB8g2ToHqVLzsSgnsAJx/gcZdubmFaV
sXWvG9+KVPCQ0vH6ZOHlKFwLSlsVuEwTND70pMtfUmbVOfRhM9PY0KYbGlhn4Nqz
4o5MWxEruT8fpetJaGel/cw+mGVz/P8/Yw83/HTYXigrGdpwKTEmf4/dUJH+Ms1/
knEZIHZrqQDumnVZUGJv9Mu+nSez/1h/c9Sn5agpQ/cWAnJuYw1ObRMeNtQ6sMYA
+Xd8os+MpHgGFj219+AAG1vOZx8LQJlwchtafFsRF8BlWPnE9yAQbSu51WbCBMRf
F71nMQ9LQwzB9DShQYbrfCdCVGOVD7ZYTEwizxKjsHmbzM+d6Gk1qFs9m+i0tkhD
ogo4ci/KvN8221lzyor4+/C3BuaSOQZ9GUFc8CSPLagxf4WZG3onuIw2aiJsHeiX
`protect END_PROTECTED
