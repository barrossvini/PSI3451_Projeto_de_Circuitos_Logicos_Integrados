`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hb1d1m4TWw5TnHN9FU43YOthvibk5/K/fnmuueAMOJqqVGwMgpnUjusS8/MAsr+O
1WpSKzwWNYxM4yMUr6hM1PlFNJyyg0RFMfRUJAwRW1vcapkLEQa/HjTv3j2ZajQp
Wkv0GGN4w/7rK+AJghwUmYozbXQZpX570w7NjOCYeeLyPqeO2QmjxZ6Qz3lYI7ZJ
SbUT2JYWWMM6DQdWAPSw+BTl9uF0AvfkJQ7t49XNqtkhN/NAC3pT9fN2VhI31/R8
8FBLNGBkt9xP3QWkYJGZ36g+oLlPskb18T2rokNl+gC6hHkkFDsGJqSLdQM6tQ9J
dkYjfG4i1iFF1Op9DV56kDy2qGeS+lZmLbQm9a68ZUpVcNFt8ZpCl6CNyl0d6qWO
E1n7xuckfj82t9lpPbzioV4LejlKOcFWAQQLnrS97V8l8tMIIYxzdEnqUfpkUosI
3VJmt+lKrQXbpXyhIfH6sk0zqiWy8eWfv9ZhuLaTONwKgd7YR3hgN+1ZNRV2GRNB
SedImwxUJ8Z/eDP41Pbk0BSxVM4l0CnliYsu9HizfdGltKCj3q1RggZPT7D4AxXa
i4yQIe80F+Ji625c4RbliWJmPoBSKdnkPNy7XXiBJ/mC70EVs9DUe2qCBAxWSKLz
+3X/D7vdX2r/HYlqB5aGt4Zh9QAWCy00LJnfKpsba146UyNRmTmG8/R+DQa9ujf7
jVRhYbsRY0DiqYbWdP2eimA5yqpfivWBPuKmzGU1DtKlHLRsse+45p+nBr6fSjO4
FZ95G6RdEhlSx34bNYO2z4gV6VuFWVOjvAOmE5VqZxHAzjdrg2o0WNZkN/YPs2nr
j77Ju45R9X5VJ8uBGk42dfhU62LtoceRitUl1PyKNnkrngedMRvAX6DkNNo9SSPN
DZJLunMhdX3oEW688ZDB5d/+jBezGKicxXI9O008BrBex+0Lx5Hx2wrU5JLXkHhN
Nvh0AqYQeQW48k9odhL54QSnK01SB2Bdu1olcNur9t/vfH2jLd/+TOajoyM8pnay
GTy/NKsdo/TZikfQJwK8DG3UbSRCscHAPKykY60CjOwBofGKKFDNV24LPGQxmdcZ
3cL+JVTtqyuvDXfFpX+0vtSnBH5Z6B4q+t8TyEv/+Cc=
`protect END_PROTECTED
