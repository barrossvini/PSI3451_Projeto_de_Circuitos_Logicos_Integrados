`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K3z/u3y4v3fLV4jleU2Mr/72JRYLvxOpfE3ZdwhM5vlyWHVyyUGpVfSbU5V+NUow
KUKUPCKV8oEgQShTcrsUdzDnZX0AX8tlrmQ3P3Fn0FgoWavPDnRZJZlsbIOnSKcy
cMpL9lHo6bobRXZs349oLZk8nlL7KsdjLhIj4XKCLjww/YYyGOIPwUr5r31fwMao
cz2/0hM/wWHDQgjw9Qvj9W5hSrye8WIVUBYWRkGAP4CVyhL/XY01x26VDVE8ejoe
YF8DT7hfjiyjT+IOBlrRqAYcr5KdDwrmDZhk8AvmnsiS+SdRNvcLQ722qKffhnsd
7wHgW/lh5YUghsdwW7P9Xvnd0ISYaWinD4OV9j6yDUEQF57aL81C8MoL5qrTjciu
HnUWH38KNMCtBWaHAXTO5DRRQoQw8y5NBJ1UNwk84JJp58poHGfJoH8x1kSoEwVd
YyNTbzk8tgPLgWSIYqEtKDA2NRzwR+FE/RKG1HmKnh1bBY6ZdgFT0MBBYa9EkYaE
loddSVsl/atNZuYZ74TMRUNOs/4jsvGiNaRsXZavvsaxgUTsbRbjOrHc1mHl6ZuS
9thKMRGd1lnfEocxMufW+m3eLEI9sDnOYyzWAe1WQABWGUDlGIrelPGo7DmcyWdA
uxL1i6grcDVgg2xWNl9eNuVixeKFkaxE7LMhUnhALmsepZa9JcX6oOZ53yO2l3lS
nA07E3ZZGAFR7525AxOcrdqX+poKl2iv67wkpoIHP+QrddJ9Ko0UAl/dshuItaOD
DoE+1QZCWFxexgWdLOqc7ujo3TciAIL40LpDgI7WzHsfimvm6u0RqDfq5rFwU1WC
hgkw7e1U6529BQksiTngjqcU8CepuRwYmjAoisL8KG1XSX8sW2qYjySh+8ws5iyb
9F358twcdIEt8rXorNmfq+3p7XwO/n3E6yBKAqNZ0Ao/Wp2gs5kKHJvEq655W9+/
Ad49ndv7rGacxudDX/+9hw4ctJO0wJxmNnZK+YYPsxRGiyX4llCZ/aoXzSdxiDuR
f4s3smgXrxgmPyjKB6dcg5JvE2fKeB7Ljqw7rMvXzxagY6TfDfsxdN44+/TFWvmr
VtJNas+Iq/5aVWvs6Jw0w2rSk/W6J+cNa5U6+WgdskQs9o6WrBIRolR2O87ZeQTy
YMuGeP5hD8l/Aq78bbmX2PyWRQwEsCx7Kya1GtZVJT332naLeAwkj8cakduNthO1
`protect END_PROTECTED
