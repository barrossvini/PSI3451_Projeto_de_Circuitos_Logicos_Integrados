`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XALuJAUbE6pz8/W+CGsQWJedGcbAlxIfNzz7pumFpS3o5lFl8OQPxv53HJcmmNC7
8Sz5MqkGBV5BuWc7kheya64dD1b1xNdEaPUSoxowsL5bLBZ0w/KPLZzkl/pKgR7h
3lBFGYYlfa4RO+Lal4ZnxXGSpX98BVMb8fwhOt/Zw1LRfkEl9VUB4EaY8/X0EMuP
SSpcuZOlLRg239uPd2FTuKwCE4lX3Wdlq35CIaXTb/vWlLjOFDkpzQV90ESebhaA
uRO8oYoqvSJZrmhYP2hHMmF0Y7hWoYZdG95lDpcMWgp0HM2xtiqu5AtTLb3wCPk/
NuZeg2WQD2lVu4dg7UmFBVv602ISriTRADTYT1NLMMFvdsQQgVwM2tGscFNbV2YH
fV/VMGfx6JFvRBYhru1fkNLFv+FKS4yd9pMl9wQdP3QNcvZcvY3fMsfjRXLJ6RUh
TPNgbmuOCJN0LiQnNLGFpEXTbwBVE92a9lLkjY5ZiHDw/ttebHsiJeBktt8I9rcd
9tlirbJxst00drtUuBRAOfrwwhOhGVODmU4WHm8S56vXOdtREV5W30EgRsdyEH3Z
SPqzgryGRTL2/Gne1TSUo4LwTryPt4q6nnqnymTAHwEE0v8IEQoVzvBDDaTkdsVv
Qyh2+S7ezI1w8KT9GtCTBKfRuOJx+E4zug7rAxSMC84gRUFSS3lkiwFZrgeqOY1j
flm0Jyo2OfPMyMmeZcBhOtHoqieOh2YbuItludrHxOErlHY2Uf0aWpALdnV1p60R
9pUucwLPG3B3PpWma1UvDE7x5Suc1McbgvdX/qLL87PWkcbreurKGxz5Xhta93EU
w99BVdja7agGmroU6KFoNU0QwI1Pr0rTyHAITCxeja79v+unC16pTOV+AvrEnHJJ
1S25P0V6HcG8pKD+MgghayJ61JxHudTZqtUxzWbt1o/QW6YjybhsEMnSn0Pu9T+7
oUvrj9FNQizn/ofWs3KXrA5w4XIl6WdEpBNiI+1YH+EKwAmWr+V/PF9uVdWY48c6
iw3apGeOPn3Sdrfle2tTGxp+JKi6WyL/HxyhJSPr7Cck8gWNGHYvOXm+eItnzcxF
HSESIw9Zg+6cvJTNX6GgOeCeEwnfrbw0iP4PLgy9Y5vFJl07GmYm4VsLg6nTYpgq
TWJgFaKFxukm+aFBCTHRtQmVU5Zv2MPZs37EaNyG+E/e0Sfmle5TmcxOgCpsN6lg
hTTbZCn+gGY3nhznwDiQqdoh/9RGgKoOs/G8O6JSSR9E6F7SqWR3xX9pvA7qhKk7
BroKK1rtDDY09h+wKYgqRDhf0o0Abr0old68sz+zfd+PsrX2eiAfdY/P5mTUf28D
IJoyJfnz6X9fV6mIM4uYsjp2TMIYtDFyLfhu5p5pFaQQaTbggTNhGW7504JE8sRn
FUPB0emGrVCCyyqM5k8BMc1We4x2z4+s7fWRh39uECU6MX+4MRPOgW/66OwQ0Qhb
LYWNXwHQK0LtXtARe1SjYazOgTwZn5iDxx5jvDoDEz/Tz+3typZtAZnwhSxDPSK7
49OQXymIeZv3MBQ0B4P2rUGskF0Qvxc0XK/glLdwll7s6uFfpqyjQUga7+BPBxj0
O011fASd3Uuhw5hNi8VBRhW8WuJgrv5fjZ+Zb1gwTTH7srDeAMOuG3eC4calIbwP
T2//N0kqvLYK9e8wGsJ869xAZrb80VYBq3M60oxLLzwCCZKu0W2/ItahBSybIYjH
+BOahxPfz0r5O5c/3JY6JqfvtqjWadr2uiVkolvv1pmEUt1+KQfpCvDfaOg1Te+g
HZBXKM47KpiXkumQHdHxWhOVIkIMEb8cc1KmQeZvUBLYbdmCmoXNFaACoRwzF4f9
Hf8AZmSmgT6ilITb1j97YF2LCgMms1oHedGMM/Yx8QnVYGLsShOVpIG1iOmy+vE0
pCCL4R16oYn6Xc2f9JeD43cfCSCmuJZ82S8bB5wlWIwDKOfGKeJ/GKYti9E2aGy7
IhBLVFjwF3yQqo8aadwb2UFxkEoIjZYvNdGxOa+lw8cVUxPewVMlZrPwHO8fOxJz
WiiLVTlxfNhcD6ZWsZXvVShlXRSXD75JqI8rpiOe15U1GUrDQzFJX9hwDMeW9WoZ
QjZi0ketKwEMOK09MWYKhTfBIG6AmbRBP8g1GQUMRFNEwXtQW+zr6QwbTyZbKff0
4UoE+R1XcQoRyNCE+PyjImiqQQfTX+Zn3qQoB7Jq9Q9suuogpZtzhX8LjPG+61q5
EphNDcaEnDvAKFg5RGcl+Ahmqz3aUCd98dFH+KhuQrJKoUEqW4Ex75upz600s/hU
UgfWDpZ4ew0azklbGmECcl2tLi0tnvi1jGA6ZQzyqhgUUy4ss/3gRub+IN7nVxmI
s8DWNmU4+XvcjjxfJgcjDFI+y/0ccci6zBiLweLD4dx07lW0TxGXDDhAsvZkJzN9
Kk4aLKFRLEbEkxyxE+RlBlHI4gq6E28hk5fLN9SA+VmPXawHL0lsO+LZvoZnhGXM
+8eoF2C23g+PA40ip20pblqiFg0Po8KejPdSqsDT12NKAl14xI5VT90zRqsnC1sl
mQwBnGW3ACuQUVUz2w4U0K22V/Wsj924vqXzi9Yn9mhPUkbV5AglLB8wWd7mPlKS
tsESe0AJGI1PVHOxd23ZpwDAIBiYS6AyElPr7a1k6zP2WbtjGWJAwpxDcwT/9f8t
Ijpzk0VEGNgWSR3x7R9gZ69Ul60ZWTmi9kYY05/KWAw5LxQnw6RYcVtLo9Ep2d+P
ZgLHtnF9WAHuMH9SQ2OtC+d0Q3x+m4GTI25iRfacrU24tyuv4pFXf3AXANhHvbj3
XCQMCZ3YoIw6yVFd59oOvi/aqRzrgAdcaAjDr9s5fffNcHQNZTLqDoKGZlApzhQ6
fwCb0LpPreOzCs6190iIitJHYTZhsnTrNiCh3n/qKfxj9/oORiT52AaKIPXLsPLB
+b+LEWc0jIOQeNRaqZpfLWSkOnRMgI49sO75jlXbRDkQpwFCT4+H/1r4KJhlTDUi
ZpVkzC0DXXFF2/Q09JqQAzUYkP55LOuepRhrtH4qTfO6Fa4MMdfGGk9mYAJVLpug
KKf3McjE9C7Cw/wluISb/NA2dmHL7xr8IIsEO4ZjtjN60k50aQv1iJNG6h6csSnm
r4OR4cZvUijk7km3v3yJ2nL/SjmGG/0reX2BU1zs7scnSOigkoYFM8XFa6t8+e9n
5/cJqkne4XWaWhpY3K7yMk66UK/gfdnHQlF2NjbMFIIoDzI9s6UZlMxH25Zt7P/n
VtrOq7rigH6n1yxlFZ3ht7MXF9ra2RUlmWuLNnajWZZTkBcqG4no+4hgo3o0Vnpx
nrelnT+ATAwA5gm2X020IBnCtKR+zRF1LGuxZJfMxjSsQ+vOMTDgWxvtzFPFW8+h
e8Q+3g78rGyNgr+XMiuF3nBkc4Jja7VOI37EH36s3Ceh2rXVMo7tLwUvLt4Kt+v+
tKhtogqH9C3pDgzOwTfWsbYFz3eHxXJ923D6XIrmSYwp/Z4FuEsQ1wLe2QhD5bMy
Y5RbWlF2G9Bxb7hK48Xsm0tvtsQgkxy06LoKCh8A8s58B5DB5j+l/GRyrDusLqve
1+kQ1a/Vk8xlxH81nv5JNq1hOkDRL7Yb97UWFGtCHzIat0u7ZZDM1Kau2Al1MIcv
25URiWanmxbU9PGdgdUlMBYGIuwJBluuPqZ3rz/68izXcJOx1ouko5GbnrGIYhDf
/tYKETWdUlfmBC336Jqh0Oh5J67N6NiRMtgjroK92OE62rjq6dlg3GvNpojq+yXz
2t1VMq2lz765VioVjwuRIx2KAiK9UbM0YVBxRUrVm4IyCRWPzDaSEyfo3nx7YFIT
WMC4ls9Xs5T2Sktg9ZY7RACYXUr9Pmej086ZTDOntpo5sTvU98BGrvS20W/bXWcE
XPYZs4sCq9hzLWnPEkkXsIf4QgovY+U1fKBu732hU/g10+hr50i/SLywLODnWFIS
FMOj1gYnXaYvXPhczV4MWaySFwxngnUzuORpzrogsME7+qYDj6Wogr5RIOQXJ1IU
ZYcmRV4wXvvUuNr5jbik41Bv8Zy13XYyOlrPgubhtJpGGIMPucVn4ldlEa+McFZk
cW6YvVbtkjup1ejPr43O6id03nUUv6YNjIb/6GRMxegA5ox9WsBLV3/VgsOWlL53
YzZSKHWsmP0RqIgFaa+x+E1hoCvCe9XWHwAsuo6BNpkc9I4c4cMxlrdviQZyc8J+
JA7PxH08BapDlZzWLOLeoJL42WezHGqxWMx7jEYCyOrx4j9El2PdJpIILNiW7mfe
1MdpA/WLt1Ro8IoBiIAtahQsT01Y0mjNNtjfKEOrLBqLlRdhQGsWA3nw9yCoAjbg
0O7EuUNf4H91iAcBSfFE+sfaKm+RFDy8NhFDKNZjit98cbJ1suAooAklbcSRarof
TE953ZbFyf6lPc6a+EPINRr+sIn9OcdUL5onEfDb86dAZw+lfJFSMhY6K2vJpVXF
1XwFkO+dITpleIZRMFIOjGhLaBemiDwoJ0htifJsxhFHUmI4HEwG4tpk+QiV7cNP
mCqwrk0yiqLQDh2hTZLay5PG1i+5OWX3umzCw2R0kRxB97ykGgm0s9RLuX8cKupP
3bVbDmCJiIn+QI+cZiOYCRdT33ah5T+knZCh1DBLoRMc7XlbrTcG5dyFev2GV+7P
j0PXyQfTgEuiglDtI5MJU87XWFRbAy5fYlwNRbY3syIckE5dAfWwME92VWfFq4el
Jo/Nz07mMRNtxDQMIZy+9CC3sZVz42IyeBBaHkthTrbRS3L+t3a19jBezXraSQko
0vxecHWNWXXguwheAfDhskGSNXJaEWiQazra473haTTXAK/mhdNzwXDCf0Pgsg7V
nDubanu0v5GOPLy3aAB+B0tP9lRgoQL+v2oBVK8lnGmZWPWravTmj3Yzp/kVfwJc
qMxnzt9ZJ0UD4EkuNsvEwAqrmZZeCbP3eH7xpYBkycdzWMgfWreK9ut1ii/adhTC
v/otLvOK+JKDBFoAJFo84wax9fE8SeY0lXK3vnNcZqE+E2jFYNqe2cdSEqrC2vOb
0gyDQtuWkPR15rgOKfK/acbKZdF4BQufWc41jkGMoBVPrderDxATXqlEiMek80P8
NF7QVKboqjRMJ6q4F02Ik3FgU4hC/eisvpmtqGInuJgdvAXN8u9QNiKSOQGVy4wt
dqrHa9jDuY1tMugjp21lL0Ns87xRiJraEs7pd0eIWnk7MyApDAjOor9qLXVxWigU
wUX5N2+4Dkm40EKgO47zURuROzst7oDSXf+5609gXOwdfYZ38PReX/GPUOvpMEU6
j3NCAZoToy2GkXTcZceY/oHk/ZeiTayacl12vIaHo9j4/K3y4P/lVFm8/5JbQQon
Bt0LU0/9gY1zTHDR0K2R6lPz/PRSirlBaAOsAw/qSkxFs/F0NMghmEWRcSW9cqYk
YX+tFjN17LIcFIWkxvfPhdV9jR3M36WPgyZ2p7PLyWCHXqBCouEIccktgx73+/W6
q54dHUgXpf9fg/Fie8gksGUWm8jDua8VVNUpJthlnCODJSNTeXLiuS1XaSuUf8PQ
5RqU4r5Bw+hTv6rdzgymCJ+U1J6TrUeo30h2tCWqhJFiGuIx6nkXPIcSJMrloV2H
UhUyjCXCGYwRxTDittibTpLm4wqC2cJo3In2H5zHTWi7C0bX+WaGXa9FkI7662lj
KDkxhzBZFp7bTVAklz0j+qplV5E5LJqb15yXkv3TRmVlcSl+0qFksWOIQhlU7hvS
MhCx4jssY6cv4ZTOPdjnOmquGcCz4y6lPy502m8Aedy+BDINwlwGBd3laFZLlXxt
nmAFSQKdCS7sGhtRaYTiqxqhYMwfPY8/Q2SV9OQNKgm9rKLoYdNw0iFi9bBfrFEq
uSxn++7oIG8mIu7XGYcTnA1ggIrAV/VeQapNS+20c6NwoVW1T35UJhDzaTlrAQj8
SDxYaYu2dqvHJcKtDTxvgLi1U/E6rktPxj0Lx39nTMzPSk0HBj2aS7bSk52cBQ8J
Y67fNpaZLSQQbzebs+5VQ9454oaSHxp//+3yATl5JmCGMLA1Gwzw9s1gkCS8hlVn
B/QYlXquvajJAsB6mceBYfgnh/virQ7Zt+9spktT3SBfT6AYULoYx0E26laHziWX
tJXBplJ7S1fP99jMAaQLXX3dJ8NoMfcmiA552OW+5Bt0cKWsWYYjD9f0Bb8ke2Cq
vnddVY7DjAp7O2lkH9fELf466C0dPz5LkXGd5M+2dav+eI0EVneiEKnxdvwNkmGp
gzj8IkNob6bHP9OFXz9lV0dTK8QNcGNWUXUmJX2qpnlSGBIWS658ldmzjA0Ar5JB
xwXxHj/7nwvZXVBGbjEN30TTWG3MxXLpBoQOPD+Q2KyCOfwf9jYYBYA12/owdM6f
ZNobbgJkdFNgW/RA6MiawiqVKAyl2LoE66BshWFNkQiBaYE2QGSNCJriGwR1MbMz
+DFtAU2niqVl+9wcd2dt6rP4qrBmPmCMWqyTxqugFuVo0wW/abAXyDscwmLCvqgV
k9qZLb4dV1B8st5l7vyF/gyDXJdTKkt6HfvokdS+18UGo0rqG61RtmWEigsmNZYg
glRSjd8CDoM61C0I9zCCnEKxb2MvR20LptfzkkKGu1kCOFRK1qFFcuJHakO6XwGL
pugvELRfLR5ZPY/MaMabn9/W2kayo5IyK1PezPVd/uOtZR9GBaCiURWNPDE41bQz
h4VrAUlJBTjMmMIw0OslQZSFZMkaYgv/3rr9VXpowOCmcn1OoIxGridzc08FgGau
8ZJ0DP9lA1GnukKhnOOXxJ0aziv4Nqn36sW6IlkR//vG7IQ+Lu7GNugzYTWzgTKy
tSNeRjRbnlUhUeXGSmgSL/N8fRYWxN2XGLxUE2D0EfTxkevdWvDTJdXnQ7G+q5yY
BAEe1WlQwXhIik28AfXmNHJLFF1z3YrmI+/dFTNQ3fFV3CcJmBwKpttbhvWAygz5
DpoAn6cyuz2V1p7kIC7ycwK/rYwX2LAmPHsaMRHnsbxPA7beM7zTt+RnQXUn87Uc
yCnnury+AK6DtauD8Fi/svPYtj2j1/hFLmplZxlgktEqQOU7pO9GrMeFZ/L1cAsw
CcHWKm7YyoJA80zRhICcp6Jnc5A9QULvaxbCjQyXnkzyypn8mmjuwfSWDnpEAYQN
9MVWmJ4WidRZtHnb2NeP8uqWoEcZdLSmQ9dO9nVUGjuJt78Ul4pHX38yotGXOpY7
3pS1/81J6wi7kj+YYBnFgLGaSr+thvq4DwAcJP2YiVmfQwkxVwBEbC0zMxDv6Xvr
9syAhPXCUO5dAQxhW/lJawfq59Dk9aU9Pl9/Efit79DgUmeZCS4HFXPgbEdpxi3J
Xzc2lokrS3fR4oioAongfNrJJYbXM0rTKIYP0GpZYWnEq5TQ3yHqMXpbPRQk+zv+
6cti6R28hiUDgmd+N09CZpIs1Y6xHwGKFV1kgrbLB1GoW6Ab4WoIe6Ton5gUA6Zu
Q8bnUjgA1Ck2OAoyoF5u7z22skCZY+B/ZCDhWKRPfNVH+wF/XpD/8bNUPF+cRqah
HZqTnCTIg42Dge4O2fEVgVnZiG1yC6MkMF6swbCqTMfeA7TlnWa6AGIRnTh7nnGi
Oebb+BJSE0p28LfKMWv1iPmQ5q3iX0VeIBn0MiQA/bxSQy8V9QDkro9iZT03zR4k
MIhkPGDUrOsXPCyGSclVkwlDoB/NjVL7IRF/gTxI+D+oiNXbh0ekKFucCK086ShQ
URUNYvacwAQDkdWMFjzbLl7gent+6+x2OXL3m2nCihRDBET32++NiKqfb5AZMolt
JLMHmfaLR7q0VRa0dOm2RyphLi3Rfw/zAxmw7w/kYWXvb+XteCjcQQ6XZx+wxNUI
vDfj8oK7eN+5m3DDZ1Dx6SgO43QlunkkExD/b6IWPIUvcA8O+lsD4AYCDAGLimO4
VFMccXdhdyQ+blfhAMhWht+qoiJ4utFU/pEadlM+W8XlhF9Jud+5GQHV5apLqjKs
jroBiZLHBMWxYDjBG2aelHuqqeTNq5d5bd6xQJZXws4a8Oi1jDPn3vmT9dDBkbZA
3KHiMwZ/0ATj3VfZO0z7ih8BQ99g+BIqn/FvKB8L1nLDc0hEisvwB8hEvu8ARa5+
KQdPJ19U6aQNk4kijAUpLtrM4Acv8r2uRpTzXuixhctDU+GPTp+wnD0k9PA5J1Nj
g+JCV42scfcFo90qG0+r4Foldrsnr9iLJxp96fPnlC9ME5aWqV7pCJ1DhN+UYxey
j2z67EmADTs1sp7rliOznz3OF1EgurINlxFq85G1eu9l08U/U/gI8Hg86iU/4nu9
zD3QIXbtqYi8Wc2gT5VgyIWMnTVQxU+OjiPQf5qEYNc7/hSGjFoQz3JGBcYt05vk
r7z0lhiXz4kxIF86Z8M5JbJsAbN2X4BUK7WlO/+MLWucMOqDDGnP/EstTzmyKK62
j9Hi/x68gHA2Murw01ib0jmUNLE0OvPTmvjZPovwTNGyUaqSIjWRE0KVo9loqXmv
bD1RzGr/Zr3pVDOoXaZhJn4rRne8W+OHJmfDYIzPJ7Nlohu0upNSYGGkjQz3U0ox
dxo4MCdPdt7QUc6rLlrzSl0LHturigs4xikeNcSaEDNgBGS7MS2DVcs4d/xpyOMV
IThF7hp9xxs0ShxolucVUeOSNHrPqkhfklH+PC+JQhd6RxVXI8//IYP8pDEJaoHj
g70MnIrCV4AFovFfCM6EcOtAzzGCl6T1WCjVA4m3C/+BCrSacjFsDyqx5YmqQnGd
d3DS4baWthdL/1Zk7mU+bPifVhBJzR7X8/TTE81wJ1+qhxFhEQoqv9oVLSNFoFal
vE9YZIlozKTL+xcfLzQMjOOiTCVStcWvnJn/HzWVD9suhEOlvNCCc8tv2MAzOg3Z
62pReZjCW0dITO/UzIwdiDeYwfk7fHH41Z5G3KNvZ9oiCbS3f4o5zTYPgzqdyAgh
wet2LroeI+Brn1FwzMyngmC6GieSkGeauUNIKf+AkfHx535mvEWQxvM5BQ9no3t8
+LUwXLDA+RGR5Dowd+Xii+DF04wzjqcWuhFdMUaroZ0CTN1b933UcyZjUtnZv/dc
nai/b+i50QyYTJX9JojSij2I7HVp5EITIKOk5OEdxwS7TPhxiiXiGZRvIcmLxeo+
P7JsC7KvtWJD99Xugh7OVnwuJAW1lvAzm5rtH2/b+QAIt9B3WFS6I8eqrG1mYqbL
K7uI0//JgrpNnIAB7vQLZ8eMVxT7dTXp1LRCkO6lUSV9JBfSxDMP1ZAEJbt/WCrG
RBuEm16OZWfl6OqWTsHsl2K5gyEsHWZlPE9y1dp0jXNfc+Y+9Rkb4yg6DTkhbof4
vhouDlDxKW2/nXzzyv7Z9kFQcIW1fO7ozhNtqvK3v2ka7IP5yjMForyPnvq+7RML
/OhmHOI0JQGeQDV6rxohA6hx7Ah4psGuR9Z9mFtqbG8rjXZrRBOcWomWC5ht7UmT
1K3u5Sq135lqdF2oTcMqg9aw9TA63bcnQILwTMa4xLia2lCEH4oDHtGw96VkTtkX
3+GNZ/nNvs9vcVqq2f4cw/NhsFp5ysmLxqd6zOnhxAeySf15gsflsn9sLcjRerE+
xUkfgsFupr3g3hwx3/ly5c/QUUCEG5DqRsrxsvQXSs1k5Zuml2KeF6HXBiEybxd9
11LKfjiLXPi5SwmiIFQHpgW+vCNdxnz4/NWdJ7NzKKjsN0Xnf8y+fD2Xm6Kf/Vxg
7dCcNsUu27hvBX61D6Z5f3f2WhmITLN2gFAhOOg2JIKmVGhOTb9rVtl9YOzgF4Vu
JcU/NYzZH8+aEEVYFfIoKHWAJOs73ik+yQFAjdCIDegmhrZC1er8Obsx+z9ltMNd
jHQCQR25jvKW4oA8uIqGZyIDKqpXHzRaWcUrNBmkhcV0trsuwQxS5cincZ766UZ+
ZuRPuewUJ23iArCTqZu+c235RTEoNF67vXhnY4XWzv045BecS6P2EpbG9FeumQic
RQy1cbIkkvQrKeFLB7U5MxHGGpavqVwAoOAz0FGu1Jhfdt1GlGl16DvuAyVUWy1W
Dw7pFcE4wyOufufUb7wVJ73zxS7+N7TERM/Z1+jSCdsehOEGypnEV0iFQvQphf6W
1nsw0Ulfs/yQg30ySQK7kSx4q/WV1hqwj6EPhOHw6Zu6GXK6hYas1eFt/vgyzam7
Obz7x+Dwb/tInuT42nrE4CnLswiiK7d69hRndVeDI6DCV48cK9pqMeDGIoS6j2bc
uEizeqyn4KkURZqX22M5gd046pH6GpwfVYAwN5c6wAFE0dD/e013/CBt1oTMnCsv
2qUEImOtZ+ZD0y3DKjPbTl0DxYXNvo1eV3zHzHf3v4sjhmY7YWc96Zf5jKu8kWJr
ijnVdz2IBm/voXVQd/3uOhAM99gc9j+spdA9bGWxWaQivMc0EypsmXGnfYAyd3hF
/GS0K9Cf45GL0G0sRRs2c13PEtA8WEeG58Azoy7H2cmxvD23kmX1oT/ohlvaVcvG
nIfc0QfhcO7VIeps43IBYNzOsDISHuWWVwADcJ4iiX5m2U5NOc+rrizUQ/jdUU+l
G4PHPiAPdeiLQLTjyKVyDDrGLsoVUehHkcYVFSHr/Gha5rAkEDOz+JHCBZ5meVLr
Jo9y4WPbJhqdr8I7wkMS3VM7Dueyq6G8Tcsky1beD1p5okn4pfaMubEEwnqTShIu
U0dt3kBt7BSIkTqs3IZpGe5HH8n3QZUQn/q2kga7j/W8TvQEvZWtcHNMS0zUBl68
k5jRsuBgGR67o8AdILh5z+Rs4GLw5tOBBlpw5jl7tkY73GKiAI9oqWuMKDLf6kXs
0aPphQEo8iwyEGwqhw5ByjvCyafIYrJQBfvdutpQabcgq2DywcwwVBVhiUhjyT3u
De0mEUOiKWZEc6mTUvzt9Iz0D6xQSd2esys/RKyHKjyFmVNoH2Iq746ViumiOtuD
84gVk9nAwx7qT38CLsKWz5drKaADBXUKhsAFZIzXk/Z3O8DozJC+Cx5AfAqQFp0r
SuykWGi6UUUGKn2UzeDCDLLdakhSbkrvG7ECe+lL6IW7DA8lT/WwjToJeIosWUBi
RAY7pLE7N4GzC1pAMw0IkFhXfneeFmXgaGEM5ofe1q550Sb3NqPEsJRQd12M/+V4
VM8Fz7iyTeqTZY7QYGNci4S/ROCowCg9bp9p0bdWBGwPup1FXpZJ2gC0v0RKzd8R
r3QsF7rU6FcEL8xQDHGVg7q8wkYRsmTlFJhkZ38bokSXA+C2AMViLwvm3jRwUSuG
iKG/Ep5Hecv17jKPmCiHGkGKsdR+2q3E98+aEL/yWZfb8CeVXM1zewRaQbqeUJsh
n1rtmvEBSOPkDdzy2sQ1S9FVio6xxJMUtwnwVlCWLtLbz3OPaP8lAF6cPAJKAwkU
Z0FPlJ9vCBjSOndjxi9OVYdAyQFjUOOEYPo3NPdqDb+cjZOQFo5rMFuJvf++FujA
xwCUW6zN5wl1BJ1174tmBKC2WpilNqbOtzP+f+NjV/BGAbwmwDUGMwkZdgoK4D/P
if51vZsGOViOa+3x23UivXdVkhU3+gzMXKM8y9glp+MgIpq9ZCDh4pg0B3A2LB6g
JUHKeUNApT6skVbfKScYAd+KqLylTPnwa8Wxmp5tWk2a6qsRDePGEOXOjFTwW6VG
FJ8rMSyHjrRmtZ7MjHsiQffHjQweCbR88j5mwfxdLMpRHCWmBugddkw+h3ZdxUDI
NOsdiKMyj/YA5FJK3MkmhmKc4rC2YALxjOdjmqiqO4Odbg0puLspsdYzN//RDG17
3+7fIfGk7wXequBoSqZnpgH71VJ7B8ERRDE5VFr4HslqfwzNnqhePUNIBQxf2T2x
JHnpQ2i4zzQ1YycEPTTd709GX3vhKbcWRxl7bjt4qU4RxEg5VwJzM2p8LmHVdqT0
kdEqJbwVCGlyP/Nbs15Uqtxq8zumdiVKrwssrDBSPuGCNba58Wv9ihoMhIroPp4W
FUk20oqAlR5hImrKnWzl0mnbTN/YfCCkntSFqYSJ7QXqRTGvEn3RYS0qH4tClEa1
WJV8Fif0eWRgmY+t0Sjv7IMuUzssTc0q12cExuj006nbUJ03CeuDaHqIiMqDzbvg
DsWNUoR0REkHeXtx/E7cRxCu0bE+AAr1moouiKJDxsU1KuYwlOg+ZDzN/U5ipkEJ
kcvOp0TCoPKBypE6Rs9um4rhh6FqAmMdVev7bQv/bAVSUG4GA1D1iHE12gJDTdZP
9N8uLv/p3QmQRou68NtU0NpEHMDstFUEpqWQmy1lHXSEbAnfPhCw9VFvzYbNkNZL
L1INkERtRtFaquDP2HYLuGfJhyc8AMxdwh4OWsw7Ym0H5R9dcm9f2uxSmmVa1sjG
qJBmO3fCMjR273XGJfSZOYfJykPj6Z/66L4oaEbwh/eNI9zc3bAD1kqCdcohIsAY
hBeL3GqMn/Gdrv/vHIWtMxwylyLYaQ0+zeW9hc9O/f2BuEsSMubIEiw+/pQdiP1d
BKbcgWMSD5ml/pFscAZmMsAXas7Qc9JJXBp8dwAF4ZZOwiCPlz5DF6T5ViPpk8RJ
X9OmQSi7uNDZgbEgUFSLHQgJQXbul8pI7wLXtuvk3/GNba8npXyZOugglw2OjgTK
jvpr4HYbhnFJeX751ji1heeFTtZJFol3CK0ZbyEPC+0wwm6XcUbo7QNlr6F5+PtG
G+BNNquqLs1A7kfIGRnagh8lFShDNF0eQrJb8cTmjphhP0O8hHPOUq0N9OEBOeNt
E7AcNAGIbR4CYKj1GBJdDm+arYGs4/pL7oYypP/Qlt6nFbUt39ht/VpGKmszhi4W
By+HkZ1TkDbCcY9VV9Qn89UEeynZzm3UjWOiRgTpDZqeaJkFHlKBx0e57xcZCW3N
9ivPCBbpsW+cj0hgNLg0sLWkNGdFgwsz0J74ZboQ6zN+5vZT7u4EYPvr/1T8pXlY
dTgN1D1/XpfFI9tXoq1G2A7mok1Py6kBiRHSaDIEPnI6z4SyjG1oDMZ0PUozL808
5Xx0Iy5XcL/mr1K+1QXSbaSNoyXT/pNUCYM2U4gAxg7Yxkrd78bS97hhNfDQGU3B
WTGYBUlmR7ew1ANxLG8X9Szyv/LKNvqdfkDcqbLCx5jHMYvcC7d8VbGmP+8BLeFX
YSvXR6KwqAE5Y9P3yiVUqGzonNCcwgrS9x+eOdkutOcf7iRXS9HJ1GsUBulXj5t5
ldbE51bwZlZf6RjBUUlKaXTH5zEWAC3Z6OraYuMEBnU0z2ghBNyVwfTOo8iuhNeb
TI/Cz0hlFcA4e7u+hvDomCOc+3wPXKogX7CFX6j4k4UTB7fphHzRMJ15yqe1v7sp
PJ6Xcdzsy5z9O4maI/B66lpDLk5R1Y5BKrD9lJI+5KWuujN22HqW+0a0soTdshXo
YkUHvHiJqMxB1qGuG19+ieHyzxU6nwAbWUCQIBw/XnAWS5k8k9PbiwVvuZU1NXTB
ACDHwSY5ExWDllekSduRaP0qkbq/mG0y/3QVjcKSuW0vKPk7TqlVMJd7eznyR4Q3
NvNG3Gaonqej7xkwJD7TIl2hRqMLmKhHv3DRyjJlB6LXgFB8Q00xh/mVkWI0tioH
zEFshNy1jFloyNtQjtzTVqQKXhrx5lH5Yg8xtPepCTJq8CxKDUoyG2vaPiKTSuMN
2Loo7BQbCkFGC1E9PmXrC/iY1+S0PRCcv5HF7czmeIDkjMosFa6CuX3ye8OEBLn7
dpW2DMbcR0HdbtZ35wCajH01M1OiYv8kodhCAsAGPPFdj05BimG7NMGI8hUNAlYv
c+FQkw6OUADbsP3Cu3yfM3e6P8eSf5Z54SpuITv+oDdvonNqDP313SSxFV/E2/1j
sGLAykjLWrTkTsIjVHX+y+TnqyqnD8MQZIiQ5IUBNiF7a/UHn7AIPj6TEnrwYGpM
iFSwMCbe6Nni+T1O973F8Sizw8DBv84mTTr+KJoTdCmH9ZSeNa10u4Lx/Rbi/2iD
Ee1OD5W3lUVXuWneJPEj+NnkE/St1f553wFhX9FnqCirwo2aDYkGGPElah0CQOXl
+UI/Xb+g37IoMtF/Jl9cLoMg0AoickmRnN8v+NrbKAvMT1fnZfFAZ+OABVZ92zl2
PjwQ8eTwJRO0MY6fIVA6+7sVoHsu/q7lD0un5fvO6zOHSJgdIPckVgGhWkzfKmtF
fFhILiYCRyEVr91AEiNiB5jWVHVIIjBRtHsJen9WdEbox5AiiXWx8i/GxWAZPr/e
Nsfa/5s7j/PBXkIFS1gN71GeQkMf1ccs8H3gv5XsblBG1jM228y+M1Ncm1f1+29Y
DWCaGNrfppM0Ad2FarmZwYXJoYPO5j9hOJUShFyVekxVnGQrR0uORuygnZNpftx3
ev9UB1gVJZ0dckhrEZhXbsTi23OE7GfrTFGjTOzMkOHQKoX8v7JO9GSH+IeXJfrS
3fraeWMZ/W7sGb9PZPvjcyPx322bx+5kMq4fvgjoJqsnJ1MRegWmF2WCwOuiqyZ1
SVWIdHsF4vWkPS3kETreYHlmoMov8cEyAWUWo6r1q9aMdh3Qg/Gm1GzCk6Fj8XUa
EenK7TBYa76sEzyhlCUjbxZiBPAThuJJ3bcfTvBOrg3bnEKFOjf061aKsuOe3mzJ
aWJbioQJN1jyT9no1QsVC5Sd/ty7X060DPoj1mGCMxEu4IWiEKvsuCReyRKaxSl7
2LpFy8naMnLZ8eBOAxDrxlHN2CGwzdyIixNViGprDmX93tldaVHSRvg13uA2buLH
KewWsTsVns/so4YPZAsEhtWkklwm6Nos6f3jIICETds4+j5rW1n1BGVCyxfl2v+Q
/wu5Ytkhws1BkLpmACtho2RUsTXxAlY4PGXPwqDaSVsv3TSjpOV6GhLFOGoPyd6t
UKdQEvUv6inIz4yhdagnW+RzLoelkQtp8ykwG6E+xwDjxFAjLo+2qBB1LL08fu25
xa8D6Cu34mAhYM+fVpnM2o4tILVs7f9lo4OJpMu9+O8E17g1p38vEAym7zD3EsMY
5hSJrk7gLdYljmWZeHoLikF5SU4vaItjf52UZdsYiI4MMXGHgl6KhoL0QjJUqbWy
xX2L0hd8B6uzdi+m/mcfCzcXKw1KR59aAPMzBQwvXJomZ09nlCoqPIP9wXhkuDTy
PF6ChVPSW/FWXxEhKRQDTrbFtiXPi1EIs5+eNVYm9FeEenVHu58TuTouU3uu+MG4
ip1WIYpCfHnFjUuMTTpOGlCjQjyh6WHNr6lzBTetDFiyjtjdAtbuugc6jbJfHDaA
aGSb1g/a8HoiK5xhlJcSm/8YqF+ZsIzbqa4wdPYpeX3Fh4K+RPigW/p9j71xXYuw
aNN/+sbx8W1dIz1yFpsSohyy5Ec1ZtFuuEosv/miyupXlcdhAg01KGh8lsEFsmQL
6SMi4GsPLonbazUaYuIwdB9j2bbXDXcVnDE0O+q1y2VUiY5bz2EHFsd3UvJJtvYK
Bf/wfzEdC8WZ8gPQfCR9RD+l0EHmcKYlH9O0vt9IA6hK/9Af4pMmP26fxVzt02bc
2XuQ/yVuMG0bkYmJTaz1Mz51K+r3lsYDSD5MYSkJ3uXEEBLBEZGXgEljzGVMcvJn
8iL+o0GiFIuqs5dAwKIZqihJJ4XfJI3PHZy4aEkXDdHUBNaQZJxeeKUvjOmaqSly
ekd846jeXZqJw3GXBTmGsk2oS7fNqLEhYXBz/kiSeF2MeT9FB1BfXe+Q+gF7PKIb
EaclwX2vjyKFDoGtZh+ncGhxYyozw0b8tX7pqHQfKQD+AOcoiUzD1FHX+r3PLoQo
R/mJBJktpXX8F2dsDeNLe/1/4lIMApM95mGaHTxFOni7D2yTm8mKP5pxCcajcYtU
qe4nrnb5xNSddWR5NXFawFLTbyZBnwkB3OP8Lek0SMiRaVg732htm+C4wd0ZIZOH
sq+AUEtyvXVFXNYbxoauG/c9iYf+bsj6Tt+Gdae/VU9Uk7Tf6LAak2rQmjp9MnbN
VbmKQ/da/LiMsjyWw4MCRN74kCCasyj+NXJ5zgHaPZQOxVop04SDmTYN7sReSflv
4GyG2FM1j53rFbtaNAY7KaP4HkF6Wk00xxVPM7cUkBEIIOrdl/6FsISxiDmgf/s6
kfV50nvy56XQbJmZ4TsTGLaF0lvn0FM2GSBi1Dk+Uo/yZ1NxVXPcy8MwvIPoZH32
ZaPOiswlkg2TqR/exj3TWow8oKiAtixfKqabemKGPn7HFWbVbLgLIdDdeAD5udXZ
zkAo75AnGQAgX77Ilqzep9YZ2qFou+V/20ttMUXHlK765N5rK9vwqyn21PTkEBcf
kHNnS0IKptrZ3ILrkK3LCscn5IeYQ5pAmpNYoBewpSxh/I6IedleQTsKUjH8s2Sz
2fQrRoVDPv/I0XFueNrgIpbr0kUL8kJk5uq93JzfA9RQTJ+i+9YkNy9sgW31Xvi0
Tjr7+OsGH4Omf/PERrrZTceUE8dp5jfz7FfvlLvVwYlTIFmK8TwDJPBAAQhMyTWf
+mL1aiif7awx2xdXufayRaHjp7+ISS/f9ABrUtPisDd0dlyinkXXdVHrEFONQuJd
XxZKVI5/AOxiGHwLAhIrLuNAbkVHT64WuPhTCBN2p3JewOrfZQfDcLvzReunfeUe
bzx1rZXlFiiRYy17JEufPvQ2U2SkHPw6srGYkE2dbbadbhiuIPdVS4JLOv39H6+o
0o1By7njUJiUrV6/3BWZ8bcgmk0D6765xbL+j6IN6LI/lsDF3XnGjglfx4mjbj3L
CLZoHX5XopI0rS6n4G9B3V8VAm9Uq7D/NDS30KDsm0fPnfd5wlnIwJKVCPU9HA+X
ZubN/obipceDh+dNxVvaW8r0jirykJgSexz8P4doDyiujBf/w5/67CKhLwsNlWds
9iTn3nk8sPk28z+2gQ7uPRixwZd4ggtbPzb2lYfzNzCZlC4qpwqKDJOttljVDASv
MFLxI9laCrvwCX9x/tlmMZhw2mrUIr9Mtn/ZJ4WKojr/zi8nE/hTe0M4Yhou1AY1
f+41lg5IzOqEq5csIv51zb1RpzWsHXDVpW2dpjkU7arbJUzSVpCltk9kW/BbDRCv
VuY8opGqWogzK1qthYTfTL+rvlUoUb1vkVLkx+EcAxVGk90n1v4XwaqH+VrYD78m
d0R9chBBUY1C+eyhDmhCCX9tEumKVKwxumQoaHpHN5Hwo/ix06nQEgIdW4ptZeCl
EVKp/TCP3kv101sSWiAGNl5Ck1mkn+m2xVkmPYz72Llag+O97Jvdt366NvDtoShw
MJ2rECWA3B32kxl22fPBmAB/q85hikM1M8gOgqr1UqG31xcdtR2S30Ge+Yx557NT
9fPUKQsC8a7p4uzL4j8jGdKPBFosjpipKT4+NYroVJ4neOpXJ3xBMio1Sj3W2TLb
Rdj6khfAaO9fSZf4phk3o5rz4/cXlgVQexYf45v6FASungyP5UiSN1SMWrBdnGcY
eQCVYtJGbxWTLpRxzB9AjCC1plmVVttltMXf7JlLLd8wG6bj2z7xfgc1mheUNKrK
OCm2gJ39zVwjZwEfMToqjEWznGjcRodK9+iflecuFrz5WPPJRb5uRsc3dAKjp0cb
qcRg5//6PsbDFKldl38o3juCX933xR42d4b6dxl9xGude5Fz2F/J1PIB4VYYMM/D
2kYH+VU9a5hSqzB+TVi0Yz8fwzuj8B9jYTjq9SQbsMQVy6tNP++yd0DQJZ/LD7wK
unpmS6sYha99Hoy3rnmcq/V/LtmaRWZgcU6d7wUUfdefv9gmkffZ3UifdYpkWN6+
omQwLG45RpKzmY5ECF6wR3fRBTztiUX5b8yJH7+G31SLtyCy9anikgWPVpovDhaZ
w5+zdzDUhooOiz4Tze0jnqHq4yPGH1ApYeaKuala3vAPDiK25USBRjapwsnWLT5J
/NXu4ykAI6kGUcz8b7L8eQRwOQKAHnnyB/dxEYmgzx1IrMDEyK4XClAtltwvmztm
EO6JIPq0v2lvPiqkiKZ03a7EMWBOo+kFdOhglTqHcnnSJUtwhIFL8XsVDENbABUO
m2UtfkPtGeu6Qifc0uqfxBBvvif/IVsV88KiEbQD3QpUlHB1CnXqPaNDE+tMgiTM
jgrpiMfTgjaiYDx+RTfhM15LkLghFxLCbZ/YnQbMI8OiI0OvQtKiVk1z4TvkyURr
61eNC5lkEsCtepNUSkKoKgwhgfFkXikW1akHw3Ahi0IeAGjphjaklGDSVYlPdWBB
ql3NVFXH1ssz64kSuBMlgKIdEDv6KxW1/nKv8/SY+YrJCemYbjIOp52MxTAkgy8V
JdHVFaFsUzGttHf7oxv+dAPN0FLknjnPTTPh9PKBpM6OxFM5rgh8OFMmBdYFsIrG
pjM1CslJcafibtuPIaG/pD2dcwLSKmaYnLN5aCmIJ2FNpH5T9XBaJLDnCwsDI8np
MBTWBUZKb0iJxVSB6QOFPUTG8ppWN5wLWzv/RifIh0Z5ZAO4oazBbYGcpfJhoXdE
nkcFwk2+lHYMrLNwHt5eF6R/TnTANniChOjGm7vGv40tEPniH3BYpCOK1OUvT9Zz
//19j15QRKCyZ7FIQb5D7ijib5K/QzdfBxlsJZSFAHBZVfuGD/Yek0PqPm4hDHeA
M7FV8Vy/sVak8KuyXO2CEIf68QirXYjoOaNXXRn1BotuFiYbcvpccooZk7sWnR2b
7XaVemSH9u6tl1V//IGrmLXa0iiTbA4kgpYo2qBncwwVzUVqf5vqDQAwc4xedpQK
znwP+/pJH2FB2IPg3IVPZ3I75GHwDup4UncH9/3XzJN0lUIRw2ZZeTJVJcVgjeaF
xLLQApXgJF95tQSITMJesHqEVsg+5aHW+olr2Wi1vZseOR2CVfC+D1zEM2C1uN+Z
Li8uP+9fqPvcN/c6xdTaPfExyjLD9XyflpPf2iOd97W2aW1RxUXq3O9wPwJV0iD5
hq4TgwsUV0QOszOhJwjtQt+rleTKStSsEWnC4B++qhuLT46xLR0ohFMjlClttj67
i/aarpd7zjs4SDew6TZ/+Q6UXgTSGt9js5I9dVs0VGODYGgs2p+VF3el+QxKVJk6
NxCHuePv3/Ztse+4pz3YadDfJHH0nwj07QSqzFZvDgGPrJ8vawotSPQCpoYLnUqS
wju/pox2dWLNQ8Ob38twNTd6NpCnadBUtm8yNL4ZYMvMncipk0wxoa54Mz1RbFXs
Xi3/vbLHMMbhRA+pDlJAfAhjzAGBlKyHMjqjfKjhZ/0arG7ixaeHwCMexa1hIRr2
aF7Xkk3jvBEb9vbbD5qqOQJUngxxxMkLFLTrA1lhOzjL5T2Dw+QKZR0cgDM7671I
0ysIQPPXTUAK5jltAmJrBBIy2bYyQk/Va/5a1ab6zHdQ+jLlhTABYPlJVYindgXg
o/nvZjYORlNJ9hXaTC6eXTHn1kVV0m5pJ2nD2P+kRUa7Bbrku4L0mY2Vrt9LHzJR
EICIsDzR0O6eZ+qGFfqOaH9JZKBFelW6xw889WAqbZuRpUjGCosMUU8TxZtcTURk
evtuFjoirz+qTRQ2I9gvL5NfYa9I9/xgGSVGXRlMGkpMGfkC8Cuq3yQUs8j4cj2M
6E5KMaYucGxqzTmqDGl3ac8xNVcxe4ZGw3jWaotsN9uSsj7mEefOY8OUJ6DmvFW+
yDapMd8GXEVEtVSaPPEldDrTP0C89MTEqpls46NKNO1OVFEwa0T5voS6Hwozt7YZ
/5xgN9fGtxYV8DkFVvI9JF8NHm9EO9+QYJf2uWT53y0wJcOLpCxQe6jdOzEBySqY
kC0FuFO0LxqsvzHZsROOwxxGFa4Z20ELEE4WjXxBNoVHVczp7DZVGiv2mUl4/+HM
tjFJtYTt2tFCv32yagC2+mFPm9VX60zq6d5LWzC1mnyKP57keRvU1RHbFeqeKM5p
K+LW0IacHB2iSgrXtUA0Ikesoy7c/ltaLK/fwDYS4bs0mqju8qp4GBtpyvfWS8lC
ZeSGxGHCKcU1pCnb9K6F47qI2z0+JXdVw7s63qEUxO9bX7oVPJ0MM5X49gJmFpUv
HZ4zasQD3yV0hFX9AcSFhkFWxn4L/RXQjMaAO9YoWxR9AAaxmc1wDaK4cEkEk81M
m5LoUak5LuTZZzzbHEnf2HuTaRWpvyGxhLxSwvrGEymLXw5jp8241DO9fxaQu2uD
y5IDt+gayOU/dBYo3bofns16lN1K1eeBn+7V8/RNyt1YjMAA40BaIKgzaQsdQvr9
DjZ4uGMSPhDKIyZXZn/OYnKMA4OF9svxnjqFIZgkUvwWTi3iVN3c2qLOCt9obvUu
UX3doyH3hbdUUdo3BTpbiFn6+yIcUxRfWdFSJXSqMJEnl1dCp5gKP+PtSFF+4ZtS
2UfLGS1CL7/SAnYGtmfJGs2/7GcLbCFvYUwxF5Jcpx19vXG7uHblysG6/qCpnj+9
aYUIJDHY5aRGHe+NfPWLCMfyCATRfm9xL3TDSPtzLpLSzLJkbts49m+v7D2J/E89
XxPgnM+iuMDH/Jm/bOhOFvA8+uJYYHYaVPg3pGQzjBFG+Q8coGD21OJw6k3PJY8x
M5vhCH06YtNztr0lkwCwv+xn8QGrstEv/TaAjGlX3MJLafYXQe9phwTKCPuhxUwE
y4ImAxFk3c3AnGYYdA7/BeiJ2ABEjiHBzjCu5g9kpZidvHvkB6Iw9WSElHJPZLhK
HFvIDhn3tyuTnuRZRLxuPktvJww31EfkyHboQovSIdkB3HZXDlgSGPttm6VdnKDZ
+PfX7SRyDhnmZvcorgh9J/4V6HqjgBLc/nL/7Kk0FsiSlBptp0xJEaV3Ctxx6tU8
a/W7IHHmJYb0214WQmExzyoo6Ur+FwsGxLGpgFlCEqBmcsxJACqrMMT0x5WItggg
ZstPeUE/GJliW/Xa3nvqrnvN4pyBfFOyFoSKrEmTLRc+av+skgfdBNnF5C8QQHiv
PNyqReTtF9vcGV0onql6hHJ4PqiUymEzQaVYFQWTKBZmhVNElipq6aHdaLMqlv5f
WYJx+8Qt2aSeV7OPYoDQcxIOAmJn8HbE2wNT0JCzyxmhYr38N8QgZ1iCD0aULTe0
mDuZ2zNf1BUEVWTqCp83K/tTCcQgBUo+AM2tLMtmwn19C5Ymp/u2QwuBk4zclRNO
XeQ44h+xJVlsGz88m8lb9KDzw4Yed5Htk21CfjZaDYq4JU9uQTdXQqrXS3jjlEEI
N2tk1TUCnDBDAMpckB7uIstKBAgTUfCGTTsLlZI7aXA5YvkkoX5tZl8HvVKealC+
2lcky5cIR7zicQQEZW9IB6kcAyvghdQ48a644dYlcrDmdKKtpzHapATtufEQS1ma
oVY2QlXb2z0y6je7agKQSY+N/xScRzQ2m5x+8mjmHwWtDmmWxiJBc3vlU2aub7cC
ZfZgSdAiyP0xsYHtyCCTy89oxGmicsaOXPFrSDa+1yJF4GXH49gtdHIX9OkktHt4
KLxA5kXZ838S16XXtYlQ16gDsMsPaajQQ+WCqb8nYmn9TWQ5ayNDStBa81gs/aKn
3YqeMpEPdWGJgZiTLipmkB7q4JArqswDt1anuetH4DfPDz6MVD7ZFTKAEqZGA5/K
6v4Wk/hH7ya8q6bUWCalBHlY2ffm0JQhzTLPSyccbopFOzkfmE+/n7saoHNbzPXB
+QqOPEAkUa7Ll++diuEBGXVqZ28wi3c+rxTho7eAuRvMQSKB1gMkNryCScMGbR5T
3UoAhmuPUu4TTd4U/dZDZYpDUrk9xu85kxQatS/hGzrilJNx7FQQuLJtiVEA1ZvX
nUbW0Lrlfly5W0yfwFHiPo4VdLI5a8gMZDVCsCP4OAnlseYvTcmqqWojndBjrWW3
Amep0T2WrebBidvyL7qy0xkjVGwESycEf9homDX4XKyi85kyd8wIRj5XvSdPREfr
1CQlz2MtyCGbdIYFzyoxOKgI6gFAF+oHU28Q8elRY+lKnGT07MyRy4FGz0ipK9RJ
ZzAeIQe99BhetYW5KzxLkW8ihzVJl2xzoiSOHKFLxkwLVLE4Orrkf87Q/3WzShAk
vt3Vxj/34UV0u3oh+mQCZRohj7AqL2SeIVyvPjHtlagnEOpa7cpnWGe2zNZhluyQ
yCOyZoCcgmLhoF5fcvu5l71L2ZeH0WnkG4Q2fnyn57iYq1TXvfb2p90NQrpRX1uE
UPZBg2wm7JjTxioHY/vYxSO71sIOkbMmf8v6AAEQc0esPcWWG7jcix5jJmrk1Rvi
UuoDVVawlMkdXxUxgOq3EzkYLN6MpXLG5EaYt7vpPXacZZ5B+uSGI6MBW9jFv+Bs
8TJdqKZgDnuy1vIDIxOiu7nsOIIsClT878ulVLCrF/Fj9Lqqy+BrXR2pPEabO7Qk
PuSqTh8DFwZF6pC8E8+qa12spd+YzqaplRoPPopfhGy7Bm/fWdWT6fcpbkDnXTjk
antcxoOqPXnGPnMEtO+gwFdI6bK1zRmhKywIxtbki8yaUjIoGCpXuE7pVFE8Modk
ePhsgaVfI6zhN3vWXBNfGU2fBLZozIHq2T4tHW59IlkeNbdC2eY22nlevZCITElU
9/9wB1GU8p5Y5EhOQxPrlLgq/exPCo749Wd/eUAEycoySRaauIw9xw60z6y4QlLh
Gmm6NOUuU9HOxGrQwr/lf3FVkprncjO0JX+UXKkPs0LNd3K0/c5aJtPL2c39Bzsd
GwzD8LEEXDNBzvLOpMqB+KYIWTMnfR2HgA6diMudA8gB6uJqyer/3g7jWQiDIfKS
vTQRcQoYvIsavUY/9J7FHcsBmmZk+TjJNQmyQ3MwjAYgsCUbHH//Cuh3BB+fZrUl
rHXH1Vs/ya6cLVaKPMOyAwF7GChYKFdA0g2BEvrTaiGD8A2vP6edydCkvPDn3k7m
5IKEhx5AHZufU60+3bb6jp/3szj/CkEq0cbgPh42xH7ptpVXrdvNavx9s6xiQzKD
1fl78HRCtWVXEvPJIdgiue/Dd42w/iYwxARIo/5ePXEPNoCFiPu+n9I7Y51MGYoE
PUIfPG2BkS55l9R6WmFM3SCC5quJS/2ZplC2yc3GCBXKe6mV68LfeyvtEArTCla/
mDIfAjb57lTaEPDFbqsLIEZXAmX/kh4fu0gJyggFA5DMbHUPy/NaPATYJDCsV8qi
bHRpwKolB4NGGTOzqwNnLABuGflB+xwxjTKyzfCuWwmfU2yxXFRO6Z/T9+sy5Bez
unlUI5vh2Bs2wWAS8yaqQkc29fyKm7ykJRaiAtRGEAVKvZJZzz+nE57dvf7MxRKT
FnRUQvEs+Xm42iWUU+NggRHOukDM24kZ9sdtbIbDYyGrstcEwc+a1xTDjSkmbl9t
JMmnny6iHJUrYMBSteXJ2J321QcnuDn3Nj8S95zkC4TfoNawS8knHJtPS2d8oU8a
+Bn2hHcbnLS0EE2NA4ESTpoKc7SjJmeGkf5s+QdGyGO1XhH0/1+QwxYSGB9HBctm
M507wsgtP7RqLac8rE7FvNgqdq2wD0d3BpPnEro3Agm5Mjw0HYe5pBwhoZzT+8SO
CSHkM06CE542NM2IvhzDf3GLwcv+OL3Te+XMeJOogpJ71zcHjoKNOYNwRF98JBHd
Pu7OQiCg2pP4HXJUoTI9BQe9R/mBBJsnY7AriIckl/ROoPgfxz4wi7uVWlCVhUsK
jEGNN9bdS2QaNECTruxSQtIdyip/nXoQQGqI4/gHYipzZN6cY87+z7ou8X/hm/lC
Svyg/i3bCdDPfXAgvByU8i5l3W8GQIYhIOfHoo7F8IBfFrBi9lFucvR7cHebzLFB
lPT1960EXEBVOR5X31gGfZwXc2RUAja3ztIgFNCcfo/64Iy2ZRBN+eGc032PDYTy
ZnGMqk9WlWTZocxnVbHBbnHij5k1fSNKiXmXxq/ehrAAtqgLdpxO3+Tyx7KbkBLa
x3WhHPYK4hga8Ta8gV/V2AQgifJsb5a9l6N7Uh0luVM5mgvLxmSqPE+q5IkH1K4i
hSnhnBDTAMIkj8DNjf8Cw7AsI8SCFJOe6j6FmGZNyLF/PwwKuWsfE4dM/Hp7yzx8
gfoWoGfYdGsyA4b/WHGbmuL7XKDUqkgXMNCDrGu97PrOwdjmhpq41CR/rZkpB169
+nFlklP0bDhH6tE6Ze17z5ifnqPRbzNyMYCzrSNwbMOCWlN5X1zfwMe0Hku52kNI
35yCLVxyOcKz32ih9cIR7C2xICMCL/viB9GgS//vDCk6DAZKkgwucElavWmvEzH6
Idw0XpeYj/M6Ba1hNoIjbgKLN2xwgxFNJRtXen4MwGm2aYXFNrQh79dylDW1nLxK
DPT/BikT2gn38RUt+dDnMso4c+OOcAQS3cNgYj9j6trZNEpeCL1cvNPnUJ9jkCTp
ZSza8bFTN5GjtzuUaiSCmqUkgUwXcfkUJcYml1otj36f0gD0s9fRu/ZyS0fDpo91
FLOO+HDJsvhmOynYG/j2E5IF2zhHIdebj/XTxes3m23QiUkKqh2BLnSgP3hviCeo
Y8lv6hOdEZw9JrBsiiQFrPthisBzcl2CvfJvVrD2WODgfv05KqZByXkUBMDT9JP4
ye4thnikf5+SnHd0Z6TOWa7KjLObqiBmL9Wr2SQCnCSC0I+gCqb49qISSBWzRF7z
oeOpmQebsvR5b47RwcCyqlRkyReNjvoBTPLiiLNTXWAIKcC4hiSDvh7j9VXtCifj
sTyaAOM+oBBk0LbryB1q6zH6ko7s0WbAXD9bHv7d9h+cd9z0Ys846nCPhwHcgRd8
0C0EKRTrA6LfhZ4yW4SOdyVcTsJ7HGpMDBSW5ShzK91ZGesYlDn2ZMwka8Mnrg4z
u/rAGs9B0TPoiXs330t/RGDc4GtDyxTKLAfxKf1H2ViqkSIBt4Tm6KKr2XM5qE+h
nihX7nsLi+icYx9l17RGZVjf8OsA8ntwg1O9pItDGy6218la2SwKmQRBRmQ7rOrw
mvKHmndxmnhsoVPV7lMMAU32gG/WuxcPzEGXbzjLLuB2K6fdHO7EMrsZ8Imi3LLr
IYg4HML9xZybPpI4xrfCGyGQzc55aWUkhbrIPJLhXaQfo7Eu7y5D6PRmwB5dtO8F
k8KjkOrgiS+KZEume1SCjNDgfcYilOTA7jBZrXB8401wXxRfYpX8hEWOGdVFoPBV
87h9C1EM8Uq40TeaLmJK8r/rHFWAkCNLm3ohqjzjIYpwYJ/vNjYNIU8S9U1jhPft
h3m+A2VNWo2oKZUaE/alvOXjWha5xdhC8tqF6QKrEJXtx/r5jT4IMrsApk3oecYW
tqUm905/Ds3bfTvPw8KrkwHhV+Bxb3irP8H240kG0P5D19IT7wxkACM2gxxmPtR3
9VU+W0xmqjKB/AybvvbT8meBvbWGSGviovW1DvySv+EpAlIPEDzL8UOTUbNTneW4
B6aml7xweXrVDFUH1jRWYURdbwXmfYI3ynLi//LXAmqTNVhoXxOwtcYKyHMCjmRW
AvqQU1jQgxh8Tgf2+JJ1c3Hlrp4bqZYmB3zYHvT5zyz5VRC0DLxjeoJ/T9dfAvzu
NjP+CjyURAL0dJLao9Tr7afYcNt8zY/jEDY0x+MAToXS3ruinBctElB4mTEmDVaW
fkOCgex2ibUvZhtXeQoTcv+T56JJp15pPJBA+aauqblKZchEKqQMYcWpcDyodVi2
Z+FBkk1ZgQojnzBALXF4WG+ChSmt7RkKxpnuGacyz1u9BlTW7Z6jzQsVqMb4dhlk
pAcbab5GolkTJDJoiFKNREjFGGToTlIhBGd0NbywtNkvGSCVEKZYSwVY6Z1KWAWU
jGbIPihCJOMbu3wEsgAQMSNdAh2Luptb0/51a5qBjB6jgGcbfOSgZoDskRmQZY/B
FUgc9nTo4reREx+A+jUg7r1pJrUtJorZ98E/QK9f7ojnIK+6dErPks+odFh7/nq7
DjNev+I9KfataJ/WlvTqSnaLs0iRoAxb9pVAKZf++KUDNv1jmtOJZBVpDlRB03Tx
3rG3xt7jBSRekRo5F0fOvFZXPIUML06IcFPjkeN+htZUZUDFJIlzZG3Tgf1ekbhG
hIl+1/aDvS7IWyX4dFCCk4/uBjC2Ri7EzdGnPduA6pnOjS0D4sl+yCg22nm0QLZD
HgF9r/iQxKnH1Y4OQrw3ITIioC/3volofo9hKdgIj+0iIVfGIsi4jvMKxYB+l2w0
dgNcovhI8RQqo/rh18IXHGn6femRD5IUCxpSuRoHx+eCTxRLPXnvcrz1RfEpebsk
ShtHdYChDvl01tOmk/lib2zU56NRHXOPawwcwAYBZD3cFOnwO59i+nf3974bB5Dh
J02qxAijjSawFK36TPP70bWHj2wWFp5SD4DJQtdHC02xl0jI/eSbg5PvW2Awixwz
bRHkNGF0QXEhfuKu/8hY38aNLXz5A/rfo34exQ2RBbrTrW5gQP5dQLpXG5X8swMB
eqeDHskP/pBbIwXRomzkNewPolSnAvYmeP6/TNynrMtD2grxOlQ+oNtwP76Ips9B
oHKe7RHmROBqSVTRjKyQFUrwtZ4heMGvACXlXMG80kcYUGnOEfvntEsl3nqGZyjl
9WimyMxGC5lfGmDgZvMytC8yGTasA3R/2wnOYOenHVKs42ofbRPbBm1Lx19UpxA9
FN1KE1IUByHedGzAV3l2X/h9nmKA0meaGqKuTFUznOlMh5nXm89lnQvflcZJKJv6
m7O1ryWucAPIaaBOHIr4rz3R5bFwGTFT/Ah69PuVWXCrqKsLSIETFb1fGBk4S04e
PzAsQwVAbk32jhRPsZl/zkXKBqEfS7lU4a20f2jQRJtrt8/+uUUd+N+/3dbqTGuf
/edO6uBnT5F9xzAQAaqAg5viT7rRRLTbd52tf0TWpiyIa8wgzO6nH4mzNVoVv1v0
y7l+h57ynjGzVtwC6YTu+B2pPV3QyPprVeIoirmu1X7glqCpSxQ9Y1wVTtsfctLZ
oZHpYXCYi+cZHsKsK8PEPfZeF0owIJWr6/RqFjPo07LCMRp0+dsk4X+JGNhYTGif
FfUMnGspJUzjM7qWJfgm4Vp8iqAeUrMM6KMdX+PAJXvIKKOoPgPnhKQc3ZCflRFI
/2QeBVKpYCIQx19iv3fQWG46xgyq8mc2OmM81JjwR+wzmFc9B7Fmv4QKQc1qikEF
PybTKgf7TrvKF6OiOZIxa31oeunRtOO0P8DorIG1MGu261c5myDMrEHAcjvrCDv0
0kEKklcCP7Zk+7s3UK0DAbVG8CmpMbpugP9W1TypdwACz/gSIoO96iWav741eFz4
WfBQLCpYrZrp6GvyAM4Gp7W6e8KQMuTFZPCkXTUcnAN1J/1PfciA2KY35WiwMAVA
8uHJ5GZdNiCYWVhicYiclircL4h6cAfiQcZugn0y80WodD/ngyJWWwWHCOmBtS6w
LY0XJgWiqk6JwQ7i0uzqG7zX6NG0Tdcw6lvuOT4newhAZmKUKHvKcu4h7yX9B2pz
nh3iV72XATjdewiC5JzVv0qsM2WnwnuolBHEKrA6i8jiz46wQidYiFvRDzMvVu1V
8Xu6JDzknNIN8lcp/muKYzA1nBn/QTn6HeNSKjJ0K8Tt6pTq6GEVJGh1jqaMTtyR
ewBZMH7gNUauJXv7aKIy8VHhS0bN9fYvkjwisIkIeCgsWcwfNPnIh1eJgegV/TXv
Qj9g7Q91HI+NERlxgevIY2GErEHQ6ed4OGXApIGkN2hqh/i9fUbO7XyK1r2TNewc
NX3cYnTXTv9yPzwL63PhXeNIFwqCaJ9CW6VqhqXQh6ybpgENgdJPR5l4EpgYH1RB
hwgfD+66vhTIUOdfuM292tRjvHxbzQqyDoF5R5x4LNID/KChMOdiLXc2AY5DnJ59
j39RxBGSDy/dqtcdH73EaTeMNFo1AAUYp6M0HeqlOM1hbQdGgyfXt33DBc/OZnCa
ME4OR99Vco0rWp4pibqDT0wTbQ0/Y7QtNdFTI7/sOPGrq9PuxA7c6RaKYU/eEuiE
MwdHaoUXcNJ/6utZrAR6SZaK8mKY/qr5Vd0EsnuwvzEjrr89WGI/oi6Yn2oOiO03
m6KZDycXSO9vVAX8gh0OUUBYm2J2KRd52H79QyJJv3MJURSkawXvQnepj6fUA0+6
qCCDYsYQ6fUvMPnDF8DsRDP7bGh0w+EneRVJkCnly2uUnoqaxq675yzgtCgOLhe8
E3Zb/yLfBqGJfyliinpVkvzkYujLeXl38p3WlFiappB42GPNVaPz91wxGrB/4XR0
2JleWG7Cz49RR3fIyqPmboWkfRrfXVwVChgvxSEWYxVZdbmvu1MQthbw1DSozmQl
AYbAHKJUtSgz9LdJ/zg0ew8NoyeoJGUWMv1Y/NyXKhEi35MW+Fc7iw/WcHXdjZZt
FnVxjY9cqmC3PsZyBaSvKxF6AB/dXCqHrwWv19izt37ig5OhXRU1byP8FfBth7G1
exmaSd7YwJtTmE345OZMzOuVFZ1KeAGndUMK4qWyvbUB07cZWk9X49iRD6XWGOG1
elJ95VHEtLfJ2AQxQob8NcjnfMTW2xj5fRJxY8Kpe8GrH96HCPZc+4wNX0On1Rsu
zuFsVjddnAnQyltIY7qd75cwN6oQ+ezZuCfIxPnmalHl6fAk/c+tyImvsir2Ut6Q
MDwE/gA8QfTcG7oS+d1ob5T4PWPwrq3JWFFq5ORamfCRagHBP/nFI/qv27gDooNU
IKeF2tTTz8pQCMCcl9tvANWfi6poDiersX+MJV/jIKE7kefZ/8RsvW6TnHHb21hT
Y3SSdvSHC89Iyr9OdGmOh+VGlNwgnM2GBdBdHLABoVoyAqcBzGUtkTeQeusDWySO
12G8T+vRBk5bZKiq2aDnRcHKCLweQ2ehMO2Azd2MeQRFsOYPfXP0H7STqzuzZTve
QRr+l9JF2ve8kNxy7TmLGyjcowt37yXDqdNMq40AMcYPkZ/W2sNemo9CSNHJUaVm
KVhwxnLHmnNFOzOCK0/hoiUSXjLDEuAdRMjyGtKQeRGw5fpiAch8uUKM9IZG3Uug
v5pMqvJeIa/AuPPZIbT4lFZuGR9EarmpRcAw0tgVX6/6zgMx18cTsac5eULtw03f
8vPQAtVaQqjVxlDohGLPdi2DzJE2unvc15TqVKQfmBP4TQ1N12wOI6fhU5CMsQR6
NSSASO8WKmihzjcpUOcbqHOH9eFpZAVTFgxfaRkB1NAiZRmKmRyaoKd5NEaCpv24
GNiZJukq3+t9Gkdz4LePQ56VOPKZ9tPIFJ7sQ29FNBLxoAAosNSHwF15mF6lskR8
wK/lAa9RRdm1YtsE14lIGmB+DYYDXd4YYxS029sm2kDO22mxf7VktMI5Cz9bAYLH
3YDt7zF+8Z/kvjS5QlNlHOdBCZfejhnUK8XHdYpWh5+18mOWqvFEN6Pr6W5jTa5n
FzvYUzvey1B2qBi9qg6ykexwosCDkRNmu1H/lopbEQncPe3g1hrnrFA3B4nk6SqD
Td6+IN86Xqb5+t+aqanei8qU7dHyJccvZjuvoF6HfKiK7zfNlH1lVJEVcsHEiqYJ
cGJEnnjO9uPDEIuYk/tH5ZgPi2aAtyhBGH71aO5xX7CNlb3skge+lmhCLzmatDJx
RtGbPsZiGQTEuA0KXJbHWpf728WpdU+VrDuzJlGFFZKI1Ault12RwU3QEDV0xQ9Y
5h2wIrUDYLLBpzWExily8eCX5V2IShUn7F/s5Lu9A7gpcWk70RUhdky3ePA9b+vl
XcyxsvVFzR+qRVpVyGdsF/JeAE+SSl7XUNrOaeVc4n6RfmBJwF/KTEkMl/qSu3tQ
O+I4QGxNAL3ApemU0VWNIDut/EWTYfdLbuHIjxsvr2e4cvmQHp7+R59ZFggCAgih
hm+BhSx4InOA0asDAx/uha4y00s1esmbCHyMk358GHJuhnCOSxnEjty6B4v5+gx9
MhUszu2uOH8OVj8LFeHWr792VUUVrwAslufLuZ4ViJ4XlSihmtWAXBoTs8rhT/L+
uVCk37GZjis+M/sS6bN0qpKtE0/QSObWE8L/8jzNDAEUTmXVnQELJKg6C77lsaZg
meg7FNB1GNHz9wFl01QkZtiLEe9dzZKkD7VBpPKSjvmJxCi7L3vpDE8ilUxilZrv
J/kCLWm9Q/g2lccVeQUQbJc2sP+tRJ3R67HbtN6wQVKBW2ctNf/BKpdCpoxvv2UB
6s/tNvu5k3t+R4Re1yzyErhLVD3CDg7iFDyarTq1aR3zwXdi3HYFmrOXY3no6Emz
U9wBwo4MQB5aUrB3dzIc65DewJIQN0IfoRcD0OplHkXjXVtp6dU5pP1GfXZZJBGq
cLyeGmOeQreP8tgkgeQ5svkXXAgqXTcDL5Q5IXYySzMWkP5rFKxH9fktagZjOJ6p
SH50aB4CW7N4duVFQhnWsPphUzwS4P3xFDmnmPu3YRDXQ3ws2jeJ2zbuJg5TYQjX
NUkPcToX9wslLeiXS22+nJK+x7RCbVW1XhZT+cSpDyd6XAY+DFjit3VaK3tWk2ze
vkyapIsXyESwWzZnLZbuPhB77xWAih5Ba8xS+pG6bwvDIzKAQNMIXuH3B+sOK6Kg
G4yYyUm6dQSXLz12DHjUpx8f12rxDMcY+cf3KGxgOdqZPhuaVRYqCyq5TPj/fcyl
AVj+056rP8lRY6qH5jZedPcV0Hv9F10wwphXV48r0dws/fiiF/b6sHx+VxrdEQ6R
NUvgcNPGrNSj9wyLRVDzUaErDlZXsiUG2qK6nnMZW8apPhNgHdp7tMoCdkyP0VOm
ZoU69pWPZmA0nakkxhaLTxMz4gSoF4YzumTTteTciNf4A2rvkgeity7+t62FHZZX
QUwijSdeH80GVJ90MDfSMJnfWrheoBRrp8zxJHceHQ1lCQdMdaYEW06d96UtPJDV
dMm08DWRScSmAwyhqS0CNMZeFsmwSmIeqqy6IIVqxFK2ukd/P/KwMB1BR/opUONh
2sZMUhx+xDsWdYH15+ePLjstprv4r3AMvBn99Wjeiyfr58aK7jvCCsKox/57ziHs
84bcmNx9MstF4iguvVBCgKOz8iIE42vyCM+9O7yL5SrMuBN17Eb7sAWCIA4GYgOM
BThahBS0UwmfpnnypBftLOkigyP6y5bZi7jZ61W3X86dMXlDEtH3N86aCj+ha3ui
zoM+dTb2p/mm4WqzkZNopKXvLqsMOgPzW4oVj8iaWMlrr2FJTbMcr1gwDffHSBxM
HrfcDS1SQPwpGbtaYjzJi1ZMMNR50/ysxjAF/At2/IkA5rTAaHJ/NZikLcfcQvMY
6rGaeJLmUVauc9IRkY3ZSgZagovGH7/9IYv8yw2y3BkqJCPn/Go6ROp/fEcBpKN2
jvNOTd/yGHX/t8dapfO2ijZAnzWK12qBSV8tpxIL3L40YXP1Fffz1aiONtsQZ5Wb
KQf6oTdE5IR7tjWO73gNgzOUeuMXk/OzmLxu5yX+657mH4DW6oOHmeXYgLJaus7j
K3tdeXIRRexaRWBVCb7++u1LkaYRvni4rcmLFGOXCg2mlTVyQcEnmzJhwo6GJKbW
J804fTNcRATYBJkTzpzjJVQFcQwQp180FmO4pCcftZhRh55LLLPmteHSvJ/sC7ai
4V4agIoYq5EPQMEulhlUYIQkIkErcXQkAcd4pG/um8LfepY1iRKFnFfacfPydRoH
Bqm7Yb9saq33fxMB5DbwSyBPwTZlz5+9F6W6UtdjyDvohfHLWjFbMRdA5gS/URnZ
cqeJvIkALmDYzvGxe4vSoUCnWMv0oPJMbRj1D6m47pC20xkUF23Pi8b/Sp5D6lFE
pN46z5BY+QmY1yKSQTqmqLvYeEQCBAMpT3nFAT/ckjNLCs12h03aCg5WRezhJQ6b
PKmgd6h7zD0NNhk8snKKfCLmlTb4IX7HQWqJNUupDTIJnOL3HUP8n92iyEMBBktJ
iA73fiPJ6UrsdZ/zLZcqYeMhEls/1fVKMf/6xtCiX5r8vqnV3Nf/QogpOnG+hmSN
7/XPaUu+rQA5XpC1BG8PdHJ9bQjuwyfaoEhctMyItcvcnnzORKIVl/xIARlUadiF
xqmCcu6uucjahQYBWUmC0tR7HIijpdGojWDHKHHSRno5LkWRzJbnduMIQgRYwbkQ
RyNwcgm/A/5qIYzJzsGBaRehJbazytGRuw65MNmZGI1dYc5pGOYXWWHqnnEC+KJo
bzpoCyZLSEXNwrjkkh/2QWj53DDitFA3V4KAL6dXpWMqiHKa3oCWKQ0zff9bSbld
KCGVXX2PkJb135oG1BplL4n3JqlPCEcNZqn64yqR0rhslDNhGFItpa1C4nE3F6+D
eceKtPJ5Miz3ILae/1ud00m0PSOLjlY4Ika2SpGTJivTHOp1hZiA4H5bibVp6UCb
VCXJkQIVpAGQeq3ib+JPnAWbQe2VcUQhZPqFwIzbDEm60K7tsCSJRwUkyB1AsHhX
QaAAPlf7Nueo7+oJ7gHwF554n7hVOYC8mFye6klzmYUS01GyaiRslTdWqWwsSOH+
OOyeA8cAfsXmoBMuEJPvHsOFHuFFXCcAE8sGhpScjWa7XcWhuBLPDyMLH7jAjXfs
QmJzcc+zc6fOiNDD7183reOB9gD3TEypYO6mEV57iyu/1J3RJA5FzPg00P2yOulK
sYw6v5VhOZ6haQMGGp7QB4Dztx209prq1wQX69m0cgaKbsBCKtWQuc0/VX5+3I5K
bVKJN0XgDOTCkWKgdJcBmTbdHsvjKU2GehrHmvctf5Kp8aeoMFcYnUocAXBdJNXK
9qYLWMw0J0tgpsOg7ezyUSeoxIB0iY1Cor3Lo6+iItazVN54AeGA5zF1T/axEG7h
rAqIPxusoF/EdLhpxWbcAGtwbZ37oGz18bSQkEJF10ujme7Yyg/nKK2OhL3K3vHZ
9TzZqOYoyGr60MjStAisRHsck1mB0wo4pwyN9YeXMYF92BVJDw+sSC3vg18uU8I6
BkMVk5n645n7Mj8IcVblJTaetZ1JliSdocgFL9cUxCN8j4vpkHYVNBaiV7ZI3YAX
Ubg6Y8Dfy+4i7nTRb9vKt/l71Xofc9T88omNNDuhL+s42BPB/A1rA+aZ5+LuHdlG
kit5gxjJ+7xy2J1CmiImVo9qHe3ZFBsPvXvN5mhtBiiHwZY159kFsMi1GZy5ge30
0FqIwTIkT+viO7q5DrDLQNCCmLtR6QQDzR9LnjJ/fKGj1NUXHCu10brykEcENMRA
1vvoNVBM/ON4SrbIGfGWpK2ehvB4QRoJ4pA/hk+Mv7aEXJdOLCBBtlD5GvVQNttU
ZU5m1tB3WJgkuqNSoPL0ZL1UFOqrZ+qC3oxKwr54BaAnxRci9/uMr4ixHlrre+p6
wtKjbvhR3EKWv+yVv1BaurlZ4JSWOdeuABVZuTCZ3adwIYsSAC/aB2Vx8Nxm1pKp
aetbsGBboN5mm6mwoFeT64nIPure5nTqqoC8t7gOo2ylNAKvRhKdBexEhPFqO7c5
ZVBYk7CBE5NXttVp8n1lyZWVB3Jt3g3s9Rk+Y8nwn8EZHHkNLcib55BT5vbfuYxu
KdY1EXmse5QYPxCBjE7TTKXSRq3XsMgnfmV0oVR7AtH8F0xWbGOe6f8sp3bfUnyP
TUVQ09TwKBL4aoXq4HLrxt06//mc/htcBlq1oQKQaBZb4Y74VlJvwMjHqUH/mS8W
nLxZuUMuUmGfWmrIXpztCljzWPIK+URP54hBx3uL7jfJVZmBoQTKXaVUDTni4Vr/
+VHAhnk1tDs2Z4Se0HCkM92k1COdKVtQGOtcclhM3D+BnieaRgB5MKVUooq6moCN
z1Pq6qh2Rv2x5+Ya8dpuvax/LtbctRDZsU6iWG9/C+szsYjngqMznqfXO6KAIzLT
tlrSFnqJG9QPUeEVZToCsbraLf7pPROOWiifXLUVZGxX+T7eDfzpdog4sLOqy1OB
IZx2ypJjFyJVYR/yrCJaJj65AtXSn7t+hxai1DaTQUkHHEexK/4kdqkm8gQt6n3q
xym4oPNWDS8aMoLybS5RVtEzs65TaSZtYuWauN/X4vkKhWHTpQYRImFR/w4MWNCl
vrwgGW8uvoFt/bD/TIYqOC9mkPTQPqYW3oQ9bDCqbsKXhdY26E0kHtZh60FfPsZG
vHn3sbOGIo+B+2wdfuIcC+cT8Sourgu0l+7G6k1Ev71RWW8Jf90HkmBQ+Y6ee7Q1
38Jgvsyc1o+RMSYCW06guzqqo5+MUQFtl5Kl7Nc3fWT5HzUdX8rB5Y36O8b30wEd
K3TxMyR1k5ixjneuPYAishepdYJC+cIIrtSOYDdoPvu1cX6ZR6yUJqKxEwfB/IGl
Qzhg2Zh8eso5AmQkShR3Nb+xNLRfqjnJZ9oHSHiZrV/aqP9aOcBI4mszBazyXM9N
lAFv8Dz+fByVnxHem4F9GST4gpMYbkdtRxShvaNBsUuQ/teT4xme00tRSyFcPCKb
bA5xMNseV+X4nHlUY3XmvCLD3kw+KgxwLYQ7d6x054QsmqgWeDfJOVXicwAHzh7c
d+0AhB+C1duAVYNkN/LAQpbRk3hgLnajOh3lDanch6qmEGw5+ISTIiivM6h+xI0I
kLHeLqDbV5woYaUBmUh9nsbl4VHv8tFU0329XEfWQkLtNfDxhyJ/LsDL+Atk71bz
/RpTKzlwXkC4UczAGUEejlDqcb+pWSc2UqWJ9wPpdN8Snqt6YsZJ2/Bnrvfdlrb1
EeScr6pA6Q7r8wqEmpKfuGivauyLxNQ8pkiXXNv9EM6WXBmYiVG8vr+Jxyjsg0aa
j4QXQopN2qdwzK6Z6peCn/0sS7La5qls/gH/msxaUZs/tD70iqd97kIkhveOfoHm
mwiosYIbMm3k4v8VUwzTEvMBRrk6SzaRvHecg8bN1dRt9M9DBPUp0HP5Gi/DMB2X
BdEAxVSi+e/E/AqXPttydzDlvFkxq6DcytNxOPCAys4ex26+zBJc5rmWr7+rNDDe
MFn5Ma5c7Vv3UcXRTWcjpVLuRQYGmvsSPc9D8sfK2N6pd8j4JtbFv4RwFpDmJCd/
iB/mD5/47T6pNbApK/CcE7r0Dmly125tLUn3+zy4IBt3VFG16QrIXnIGj8XVuR36
wZDsXTAPUFDx2Nk1sXdWfrJrwcN8nWXTVGXk4qsZgP8Wy84sxFjXRW600W8MADWI
HvfEyZQdCkt5ldmH50mbWmfQuSWbWx7/v9rVw3vEsdSzpTKFU5jvqUOzc37BLJc4
aX1RxTzRqutWlJjEk3HsvA2/upZAAbKwV85Z0kUWtN1UBkQ28CER0jWvQbOUbXJo
Nv/dUld11OrkBoZSncSiUbGywJ6O79z7QuUHA/eHeOmXFbJ9WcgQW/cCbx2SWgmF
EqVkqBS+lpbTFf9eKupunFdZV0dj4gZJLELOtlQcXVmmx44wpQS5Iml6TASG+OI8
P7HyRli6YXWw1TiOyubQI1elWA9s4ccMf3ivYnCrpQikDMI9kJMZM7oiO3aF+A43
qygobJR6+dRDCBWeDjWMT33UBnlTo3dNfRgDxImO561hUnmqp99W6lEMpMtZarB1
ZBPikan3xutBHLLi5+nGFHbsZstrTGC+z0Cwb6DJ0laXBcs2DNe1EEcjmVJZoEs2
2yOYCp7cQeYtLgExa8sNtbF2qc1/d5HK5GG6yeAtAQzBAJqfvHnsVCKYK8GQ95Qt
5wkGH8Fm4f5EGHXM74S7KXxI81NRZLDoLRu76b4P6sxHfHbjXloeIirglfZ8sIlD
MspTIdR7lrNB2DND+SfVAR1oZ9Uh/QawEXubqMhP9K8ovSzdRjl2Gq1QhHzus2YW
SmVpcLxxNg4B7OFhYIC1ZrWfUWZIe6PANcCFrriryJXdE45Juk+GNgVZwqZG1m2I
P4lz/fxVysfxM6mCLhnG9tnKv1Tlkoy3iMaLKkxOC+cV+EMuqOn0Ngw+9AVCd49j
TKQpqDC2O190eJ4i0fVxcRMsipP98SQSwzekjbo/gV4oO5si7mwGkyMac1kdeUW1
GxE8lRma6HK8Xs/r0tsGLSorWTMttS1vJhL74kwbFaBqhMoipBh0NmBDmOFuMSEa
t5oQ2lJud5Pkf/xzO1LQrKZXqX7PbV0nxD4OIJVoEuwStW3B1T0FYKLYyphejIy/
qLuHVVC7WcShsLuKG0pG2lxNTrs4x4WdfCcU/QRB8fuk8i9agzhoRKq+4JC6PJKA
X3gAW4wDoJfNxI/GFNtA96GulDsVQNv71MvmlRWxIM4k0zcXWyHOaDJDyeGcwMiU
5V2chmyBmpw04cNaMWzlBAFbHE7i8NO9XBXQ8Y/GnGWvIjd0bElpFam6mQ4w8nKa
trObpBTmR7zErSMYjHQt1/acp4ou3AE2CgfNurtH45bSWpUNsxIK5CLpcjAl1z0J
tzDNdXwZCctPgVg54lvSR3AAxYfUFrUVdEkiBxd+tvLBpYECbAD34p+OCGEzvgI5
U9gdt3qPE6F9MmseQHI/YF8SyrX8R5j7eaaPwV/3oitmNruQleXmulsOwOX/tCLs
/fdRXlqwvLP29CVLjDaocyRKZZHOoQ9TSuv4yeFAoILLDm6/4n+HZKZ9d3TTuJUR
NWdJqXBJpiZxd+/ysn+RdLP3Tim0HyDsLSSJ/1Bh22He+81SpRvoBP6RszLJpw6S
5uPekeh6iOKVRjaUYP9vs+j3R4ASTLXtPKJB/OvfiECXy15nP0mka3yop6mWk+6d
uuwmUwqvrzYOu2i66ZtuYsOE+kfM8xD0ZQPeByMFgK3dWSznlhS1eAr9hR1+AI37
j4/ET3msfkYDKlq0+8PXif0uok4X63IrawhjaHuGfE0RQMiHilSyAQ34HInlrKWl
fjUygnRD/frQrI2I7aMWWh6xZ5SB+04slLlYq3HSeo+war8u2z6x7pGlOG9XXB9e
XuIk33yknTfNN92jNzECkLnt5dR1OjMOZEZax6fQlyKvluM+eMGe0yDNrSOr0+SN
aJpNuaSZ9yJG4ZfsK/ZLRES+bla/GspLIkifJpXUZcEVE1X7URUAVud4kmMzqCbk
4BtH7efaPov1O7LHLcimUadWTQKmUPYLJaSrkLvFcmT8PzefsTeDCZTxW7/0Yhtb
h9B4I7uYcjMXpu+/0Ai0CCpKCTMykE33KyJvsZUhJB+XJieDUMhP6oZbm9Hp/gCm
cCpnTihBXOyITVwUJt0oGQ6XcHqz4iPolEKYQLpwlAsb2mHHNrZb0wmXDshSqDgw
7K/K6kejIK09PCEpyVripE+G4IVDqy0qF8m9NoEtrYh+IhvuUcRtV70pz/1ruxUb
c7RkcNkWCHuScqNi3cWHnBryu7KV5yl8+xIuleVWeoyAU1eYkqMvrHF/O4euC2dp
ny58WXjYgzWlMX2AV1Op0PuqjScICdP7tswCELVSep7OID9n6GspHuBhQaQNNLsX
UQT3wJ6WwyvWaV8cWmRW1TiGbyJI/eOmfoifePmL8vgIOK5j0tVOkWeguUQCoZ6r
LQ3Xx7JNt8v5NnPJ8S5RKGSWjIHBiL19++zcME7wgW2o+WocnK7fYoHHfpiYopeB
OQaxAA1guCSBo7RD44x4qx+wBs7UOQpnPossUKw1J5yQJww+KJknnh8vkC1U5/PM
+jQ/BDKwjUmNwW3/oLU1RbjfqNOnRf+2v9Th30MTE1xyi33L937ep5MLIdNgE3kp
O9Bicvy5a6ag8AGvckZ8FvoBb3AV/rfAcrmeHEaDbq0sddS6F9+Hb/fnWxK3v5XJ
fEPh9Sev1kUkwLtW2jhfpHByD5rvfqlQyFVGKVtkZHkus4XWvm70YdU9UAijhGhS
OLBuhBbYd1b3ham0wgwPi+IZ75z/lQcTLuYbQPQxE6kNd6PdLbsf+eoRAl1R5gwk
wIrjMoJlAdm9QIcfuIE/mLNt+9KLsLqkhO4oIirAe8ktZq6m/gq8yscB3ziHgW9f
jxQ1r40rkCRnNVPUTc9nu5olsDwnFl+RRu4NTf+eJcLX4RmqEa5McAmaZo/Jey3e
yTZ3QPj/9lcNt4x9P7JKGn1ymr919vO2O3bAYs07rRIc/kCw2v6SUlpXN9U98Ylk
xFCOVfJtLWa535Ww8Agj5Lrjrq6L68rjuGzxhSjhS7Isgni0QUTp3hEgS7eiq2Io
4Xalvy9tM15qNGnE0jZFk0JMx4iASMG7yo9k3KR0gDy3R/7xbpjO30ruxszPZpFo
0DHgCXq2AQ0r8W4YKVTKP3itIKaR4Z2O6S4k1R2dGPBkGqDLqwQF6xsK8DTko3Ki
on7e5PbdHAB/DMugYrci7V+LD4kybqOLC1qYnmqU68sE6hkyYueJk3CezS3TWNWb
ojQdQ3jWhiwHQeF4P4kmqApNbs8HWCmK8TUK3nnfNVgGe9+SGl7dDE9V+mAhCYDB
9aQVBuHIdk/PL39bCjNLaycXU+nICRf4//yPaZc1aysQrVlWxRzYLBk93pWeRlHD
8DX9jf8iK2FLtj2vtaw03GIAYcAKqSW0D36db86CwRRJnl3Xu02MNox97C7v1PUL
LzYSzc723vS3X9ksTsn379Qq8HjqyvFcSr1YLiSJoF/iaVAuiH3tEoMepSCh84Im
i6aVB42MFvN+UADdzIN4AYcniZEJMSsCI5bkLBMqO8QVPyGoVc3uZ1B3MMhZyBGZ
vdlAyTztIEZmpSj6mGqQT3Xmk9V47Y/fd4RUiNeKdXevaV1Yy8aZ45KIzy8ILA3A
vCTlqRC6YXcueJ+dGJVqAFX4wHSeT9cxAv/oEwwlabt9E/3qBxTxe3VzZ2A1Gf1T
Y0kRlHYZ+9jYIkhfhmLs2XG4OKeey6+IEM/Cv288ebD7jBFJcUHH0hfMyQr/hhgp
FeZjv6ADl6xan5ejSwyeJ6DR08tcwN5FdVH/MbcClDyHDz5U3pka3mGSNQas7i9u
PmG5dLOr65Nb2fEVbKxfqtgGzTCmF/NACXmiFX5xUMp0QwctuPREWKX8uRidtL2g
jJyhz0a8k/56+Hn0gWMC5HkRNZ7/EgGcECtPwJEPjYAVx+h5iH8cbrdT9UivhZH/
N2BEBd+ELjJMNVm7Ehfnz5oGZowin0nUePSOZ/ZxzZEsRpVQv1AH1HhUOJ26Tvx0
KiErshButwA7fD8sM3ojvgLLg3tnE5rwTzDEXrG95EA9Cdz6FHjMCteDKs6vzi4T
wzmIbCkVlujE54MmCEMxo2ym4iSI/KdItj2CiCFOjQ336fujkRCckN93COtLCmrm
4NOdbvwWTDXBPG7Jux4PlavSPaUJXXnmKlxFc76c+p5C/EwICV7NbuuxGaVFddNf
dGzzr48+oiHmL9LxzHGroDFmsfAI0z01yzG6iBlBMcr8hSD5Ng+LyoTt9H9CV+VN
wBD3MnTjp0J6no/sDfkESXomYZQQB6NPxdBFtEEQQ4z8pdNte2mPplVUOVChej2j
Op3C+FzWjT8Gu5k6HvuGss5Qon3J86BfUdrk8oeU1krOEuQqNBzq+MEmW3j4SGEV
hq4mecEnRlodoOxTJ398ccUcHeAZoPZGgVcylF1WmxQvCOwuM5vEnQ1Qm5lmle3L
Ls5KEVP7ks7bernP1NaJhRIn0xfi/N+CIT3PZtnATh8dKq60xqR/CvioUNxIjcDG
1vKMIu4RkCGXYnaK5vfZRuKJHHwaJiibsbjKXbUVc0ZRMyGYGt/gKANrngbX7cxt
vfSZqCma2IayzoTvuoNbUJcrkjtW9lL5EymOIX0FPbfm8Fg5JrecGwmNO02BirMK
EIxRFm9CeV8nxGTs42iu9E1pdWB9XnZ9LOvm2JBk3Zd9Mvv8PhkndJjzg7uwRhA1
3QG/Hv2BY9YvMY88AEf79Ac1wz1BikobzCOSRd/hVa8sryqZGhIKDb4COrQ4848i
mMfBBaOpgdjdS9AhMJhw6zXgs2Hu1FfkKB9re9NkZCfxUhMkoDjbeUoQ4Rwtbqc5
Yi59YZavBb5+N0XmUx9L4o2eeU7ZbnhjBBpoLASZmgGhPrOD1OflJ+VZ311q8RW8
GUnA61EfALPbQKNJYjmhrElktghhHHtsznml7kmdxni7ZBGfIY7zNT+HNtvT/PZn
Ux6r08hqD908y16Cq4ikMtOIndHmL1Bg113DmplCFNCHTq3V9b1TAEtiOL6+n+vS
yXuShDF20iqrZUedDPKFOPURuHoqoJu370ev6KS/6tCsenDVIJdeCDVSgIlJrxS2
A9clk5qYs08MaKUY5TOpYxDuZ8VFBeyDgA4eSWbZEV2QoAzxy1Ynt9+I79lhRJWe
qRRwrn7GOl6uROrcEQh2nhhcM9E1f4e8wfOQfSSV0NBAUzhcL1liae4HzbFj63Zr
pCgx7dS7TK4sM8ksLqGp2KXCHlHg3WHiujQ20vXEX3X2wfHOMppF7mvQEHZ/EMad
Mc4RGDgN7TYxQqiuGondvpCq4iAkYhuaP2Bewe2CZDcOrrZ07dGwlcoU44kydqyg
1riXCo0lizMqjLcpFjcBpXIfTOfVO7FEuW2wSxBeqNsLvdj5Wk1Tafz+X6w0Y1su
nhC39YCa3oNPZDt7a6yDyWfmHCQ2FHp5KF0XfQbsPoh2FiZQbUk4p8qz7G0rqkRd
TbZuVWu+T+xWVsrOvD9ZkPglU2v8fJaZ64ob2ps9WTu97hF/ZgDLNu4lPZJojDVx
vlMSfuVFO8ngk5xtfXH+SqsZLemCKSgzvhOZg2K6eJlNIq5jP3zIU83mkSlzjEr7
D88bm2CTI60U31lXuQhHPAp8AUm+4ZEnJA2zY10b/nZKjKDxDdCQ6goXwj1KrVwm
+Hy2L2eYGL1AcQM2oQwylfgbpJmCcEOghCTdOAqrclRcTRMLNJlsh+C5dhx0V27R
gisav/JCc46lIY0+8Uw/khxw4Mh3ipjfl9jvX0L3I6cS2ks88Ymk8y9IwKimmICc
24AKMweqGHqvnrjoaTcmhP6OKX1vmv7Jn3KsT2cFF9KeFbnTuzcF40XAySlqoJ8M
yODxgQx/5LEGpOOeGF2Oh9oMEc5pJbeKMMbFOCie/geUnCKLGLk7mUKom+tlQK7t
Wc1zzxyGiwuXRl2HHAqympE61pelI6q+5shZt6f5LX4gRykAHpWvuYWb53ZKfUbs
ybfdwwVorIgOLGpt/vI5geV6Tlgy+bZaD1W1jm7x930PlEKxt5jSRYQldz+IOQu5
0PVLQT+dEqpC5Tiy18lcwCzIB6ZW2JBOTEEQjkrg2rE5EQwLKZAvcjHzlCRBuwX7
uac+ZktVQ1yZmJukWn8v9y3LkrQiHiPZlcm1cBsrL/1iHqLXlgYm6fCXAFqEzQw9
94EG24kSi4eAkPXNJ9dl6FlgGpPoh2Hm6REk8jKUGZ5AGAGJ0q1pRpI4pmCif8YU
Tw5tov86/dTMth+c1CzGWvoFE9mrm/r6yt3HYVpNyAU+N7KZhNoqkZpe8Wdmqjn8
6KSehKdXNe9CKX9vn4wNGFp3P57A257VQHEu98ydaPlMyMg4MqLNCGX/r5WEjZpy
x+NAxoyU3UEDHfNtcL+Yn0HaBkpckJOXDJ1Zy8BlzCjVBCSAs1eEgwGN6JlF79vB
Pef5cJfFCzeCLq4vzsvi8Kx/kPoLr7FoMsP9G6xcnYTzVOEfHZfrBghJ6iseSIGj
2Sep0HI3ynRS4bzv3DIlDmZYOJkCjTriwZZFripAc71SkALRIDbrRK6MReCVxpLj
+lFyMej/ua9NDUUnlsK84bpRYRD74cK2Lcr/N0uULUKUzGkHIusqRPYr0gCciuMm
YcIBaj6U+LMhLcK7TQcR3uhQOlISIZWU+7yz+y9CpB99H52NGPPYzk4mtGgiLj7H
JtF1KWgwJXbBxh9bT173nQvPc5UeyC1suBtQDlASrgYbcw7yp4iE9grUegMzGWUy
cyC6o6Wqhp6vndXrETceqMQBX8iuK4M4cl3tUhige3lJRm4KGBWv5jK5s7WnvuM8
Z0Dd4jv4U5awkbPAZ79S/jEb909psQIdECNUHLBDj4H/WttL/sgn98IbiKcLuUKs
SJ0l5J7hqpkE3pNOlpPreB3UpE3hjlh0OhjCzgGkFneHMCxuAnZf1FNnl0DphfqA
/0NImHwxwgCS/hRVVgBMAx4v+UMJjLC6J7eFWncVXgEKlLW7h/IL+v0hikuBpDum
Em8y270M4iQ8jFupWlbVkE05ypysElnkaH7EuZVZ8VnRKpwu9pB6Xmhuc/lCZdfA
vzcfCL8iYS688BhAaaBElX1x8j7p0MJlw8ZcHzKZNI7qLy2TLyUOAwrVPyc6E4o/
87nJrRad4hfsu8iHxtlTpPVrUJG2t2HiEbzUpD8dY7rkmOTIwgqJqHWT0ZYc4YFr
FFoABGI9/eTIcT3UYXNYTibPdgbtIFEuMYctWA44MpDpwypyNFFBuX8/S/Idvh8/
ykRcfNfOcvEbob7tV4m4CCccp8O07LQnzG8/+pEJqkNYtJxQ+UtYOI39RHHp7Akj
x5U/q7ays7Th4RtVmTnJpVlkp1kylcXoSk5yYNepZcPfYNk/+l4CqNV7R+RRMfPQ
V4xq5zRCcATV8c/nHinBpUu3BwGLPeUW3ylyCpTRTdzBkY3CKvCmmiAlR2az7GBz
GoIZVJyBSrth3MYXdIYhfvAg7hYvfjYwc8AjhqfIwBq7dC9n/WVe9navSWb4X2MD
jOomT46PxjJh9mj0cFKNvr8F9+JeqAHpy/rjn5EAq7XUTVSWyTte17yVB5uMGcRJ
Uebim7kAgH9VcAMMP8pjpQLR489UtcrtuVAs2I4I3mXf735y41WS7Lr1aYe7DymZ
78DQ9XKzKnQCiM3Pus6kpLm7QfwKh0BlqlOfCtWPXCVgIQG7NLkGzxpN2uvn+afJ
DRg+BIsjMqVMaGdYI7rIwdKAFVWKygxS7Gz6wqbhumKwXu4nM1dmKIu3KRAYga/D
As7tFj+1FbOHpitRCMQ9G5ThTdXQZspBZJoR0UiDmK7eq5h4WfXXhm8mr6kMP/0N
jmT9e7aDgzMZNg2hTdLiZyKHDNZNSlmmypdGxV+5u2kPILF/sHP4wDO89wR1N6dj
S3WuPEzundR3EdiJsSMUZp2Ofv36x57mcOVR5kwYyNqFFIbUImDdN3tTn+KSU/yq
K5I17y3BjeGBcT689kKtd7jSU1GADAFwplUigrapXHozGX8RPbTdsHvLv3rraBd0
UwSA0TfMSliPoVB9DE3IS79eYXTFlHlP7eAiiRWRJ5GMYmE260BhxgcKbMcCJ8DF
+BgH/keGKB5UelyFBB4plmMrzEchlrBjj0M4mWsh5Y+aIN6XvwDSWYWFDDrRwmHK
e9H95vlExRFT8ggY4OTRGQ7QLhQqrn0bRIPxsT9QOujD12vqXckg1GiGMNZG/89q
fVMScFaIB0Yi5XYqtWe5gZNff4UMueFT1Su5r6mq4wT13oCxZpZkgTvEFB8tOdS4
n0RaILyOBpe4k147plJSHACxMUKZB49NdhF8aM4ip2JkRTiVSTXM0tXBNpa8f0OG
vOEDv/WOXhqo3Uza1JCfnHkh7cGKnSNtJSPIf/ffh6emoULV/ZNcTXSeDtj2ryZ5
bboW1I8qZGyLvF9z5CJvulYQjOmD3DRwlGn9LmWtzXYer+jdUuLbdkylTr8Xzd/h
hseBFMHc208sTe4ct/L6HSg2CQPoTBpMqIlNtHSxQ/AzwGSRIm7/ibGJ3LvR9BWb
a1L/LRWFuPJt8UjKrTse2KY6x086fnZO2LAr5hoAp7Cu/EqTsLAGU41Nfx/KQGK6
shE8BqYGMky6amZM6Od1clpGch5xgZIaHhD48l7EMECgk4jes5A8hRT7vecEPzFH
SBdszz25mFSqXUIYRXGAsmC0zFOLdU0hm3qhJtDSZTvoZa2SbIEXloY+pdpcKNlb
UYLCHA2FIvinu5xnBTFPiDpAs6JkI0NQgCPpTm+YYHqPnHy3Mu2s8ORqh9vaKMuu
7zClEZL69is4X4/Auj1xKXhDpz8sYrC10M6KXCNFHHbHiue0YPrkotSq8yxUcAEZ
r5F4m7EAd9+AsfyeTZ5FAlqm+/OCEOeNgN6dtaRBAB3fswThEzdyKJnUwpHie12T
2VFBQqv/BenLpDQt7yIKCaFEMKzRY18LdXktdGwa2Wc2FZJ/fbWivKbXO3cROvkg
C398yOWSRyIG32oNRHsZElLYxlPJTxdjLvFR3TQPH0a/v2XvhvaazCySeR5+PcmA
fvq9Y+Su9iPNJMRxD3VwsFf0cklzhcfuFijc616oevY7QHDAPZUQ9F5yH+iet77r
YwuakHbU3+Uek8SorpXNk2L6jc0sr3gYwntXnjSTXawG1VSKnES+T26dN7aUOvoq
zgJ8e2AhAbLlwZ5iqiInI1m3PJ5NqEoV/P4zF/3c2avK4ASaFXPR7u7SVL/MBl1S
GV6BXOCfn0J4HSPIXcuQSS81ToqSk5ntffZvuhYs/Dz9DMakLesu2dfAJJlwGM8O
7WVM3BRtDzFJG4KBVxb92qcsOG7ijL3/Rm8yu01SvuY/iDotQIO9uh3FM+l/i+tU
jhlKb4HifMgbj4jD5PNPr+7+x8ctkQlK1BRxs7LmRwRQ1hzYYFrc2iV+mmu4QeGW
swy3w085IcZyav5FsXw9Mta+utugzbnqRqvOY1xKgiGavHQJePBYgdbh6D9pBKfl
c/pZ5025GdBWbA8q+2ZrwKhRp90BRjikFUSJWe83GGBNojcLosQ015ZplDA0JUiB
mCoH/ykru1Oqug3tXyDfBiWlPc52t1oWK6DHE4A/ct8Iv32oF7lgO1YZf9LdO+C8
J6evsUjU9vGHoxXk1zfcQ9n77FC7+4fqfON+XtQjoeMP2tT+1lBoZx0UgMSnHsN4
Wp8hRp5Toe2UrD61daDms38ITbIAscnXefypIdYYb++ia357xESuIL4nxq2ZWl+a
P+Vie6+Mi4+KtzO3Y1bdcgnNctL/4o6mfdl77/lqQgpmepM8zX8elD904M2mj9I1
s1D1gl+F8QbKD5/Jzr6we9hHv72QxnMNUUUdTRrEI08el4JJp1qpb19hatJhYBeq
NYlEyZiTmNFg3+qJVW0hnIZSLUv70IYJkGwjsoKykyy+qYa1K5FclrWKeKFyBBXi
NVGh6YWrzuiV2EWIHyT/UFbbdyZgKG/QA3/h2bzWAkVOkz9tkg+nUlfNbQ10zhsc
nNhYLWe7aZj73iYOl7/2TbpMFsE9Rfbl9STrprztncBCngKXAMC9Oc7ZSWBjI3Eo
Ei9KSWVn/wqy3XaGx0eX3l+MJwZTgmaRJU1nwi1HEzELibodXJVm0QIRr4ZHAdEq
BptoZi7msjfdg9wp5xPBVwz17BtQCbTJA1vnH1ccu4ogkE6uBXYLb1sxZKnMu3Kj
XNNGj9o+oj9iVytbin1NXKfk2g+eUWgybYSdrWO6lXUoJt7b9qucF3dY5ViTzdrj
jyTEChLg76MttgNaguCEu2eiHJ6tnkGtCYXcaswLJ8AY2xoHWaCBm0v49EoXc0p9
ZvX59v/V2d5pSF8Zw9+b0dZ+r3xXSAV21z6hMlVIbUZNvx0/8sL9V0kmStI3y2dg
bPavoeFrxzFkUg/1K7MTdwl7yLjPggBv0VcqW5m9iPYraL+UG2KXlKikKfiCBiz3
aE2MyoCuGGADmEnvoeSQg+GmaAM0pXzBcUGhY5Ypvu2YZpr1Su1FzP9xnxL1jNOo
DHD8DOn1daIXgm0cTr1vbzpwFO/m1cLVMqBP1XfF4H6EmaUu28QFk0SG4W6Nndbv
yROTiyDnCxx30Nz+Yy/32Z0D5Yg0t25DqiZkzV3uEohGiiEgywnb7mBV3fjRMv4Z
+pCYVfeRWQ9AshQOVFQ22xx7D8n5CRxD3sS20Bsm6xx/NwJuEcX2OtEooPyGDBEc
jnCGpsXskpZKHCOSLixIW8s860IHx2vwukATAJW1bqfO7dP7BFnebtTKJs54mTUF
AZx2lsPzCC4mdGxZygP5+FfvF8bFIgJGX90zuotKLdiEryMOgVXwlsUnJIogXUkB
GE6RWAIhc8cxP4PWLBhO9UJsdpfE4m1IsGYFbqXa2gdRX1OTWF+oX7vD+VmOCUC2
NtBuiUhPftU+/gUpsp71x5idtOmF9uqwQwW4lf4qvVtPrYmho0S1917Up/BLZMXL
yUYWXWzPreB6P5Dh1UW+3wVjxcDVdA0SP+bxQadW81G9Ki8fdGlUvbx1jHmb8ppG
ov7V1HjW92sVBepCTYwJII5RUcaP1vphEDfS/DiIT+YVrqHgsQY2/geNdS0JLH87
NuSYGFjSROW+WLg7AB9YKGnMK3QXRzZc6fMlWy5vzhdwQDURLDi5nKxjnHTIyzjg
OR16Xl9WLT5rnz7XzqDgj+in+qZVPNnfDgaqz648/xobG9ck4STpqiLqKlz2LzDJ
EkwKpS8FBDzfYX0jzjZfOSaIx0Cs/KWlqAAit5qi/Xp+vGYmBnPtoGzk6oqtUbVA
dNNvsXj8iGFQnewAcIi1ecDTMTHhTBtv3h7SVTJXH7rxkrFtsiRSn6R6O9nOPoed
7NpDMiciNrTkaBnmU/14Eg1goysHavOWpPo1fYzHzYk7hAQi0ruvgMihimSZo6XL
aqKnF6QlKU63zA3XQgoB2fFZLtUis45Bda/s9vKkZN6GRL1vnl3roAHgLgDfYlEB
QhlmW/Yx6OWrBqxMkn7xLiYhiVjUmPZ28H+Vpl9l2sE8MFEUq9xuS5Iom/+Qxf0N
rh6YPEM0CzzQBLzsomTTSWQALp8Ajs4kVDyJaGlLGhqQ4XCpcx7wTTshNDtOk9He
Fctd84DQcZ3PJR1hdvnDBL7gM3w6e2mKm3MGV+iul5SGJ7CoIrBZVOVACH+hqZ/9
M8jQDczGUQwgiyrOc/iMru+fyi0x+w2HnaiIBEVGiUjlQe8PoA/Emvo/YaDpUqTF
ZMhxu1QLq+K9rVyvsXpy0URbxKie5S5v+AZ9V7EYMHIpUl6qMgF27E+2fQs2BpAb
K1g80LOqleAjl1g56PKBV1TZnKUPZ0F7o09KWBs0oEar5fYS6gu1yMD2td3bsBEJ
gthyBXDHe5+N4Jt4WeqVtDog3/QmUq5iOG0M+J8ok0GjLJ+1SM4AExD2ntQyO64E
IxJ0Il9JT4uv7lP8Su/mIfbH+Uh4Y+9Dl8sNXsMeC73eCXfC9lvDYTnGZdT7xbbs
T36keztKur0Zg25NM60iUu/PyvaeXS4Q7qnVI/ftHFETvc4iSWAbFTQ1eKcQerWl
Jcvccabl2AhCu/GlafKsEo1rx4ez2WLg10rl4QQ445oy9OhqL3f/ufUHRTYp5Prg
oDmyF+Juyf+Mx0qn16wRTZga8KYq1pG2lKoCF3VOWYQ7IPFb7j4w6LZRkmnjD6cO
x7MM261y/aDTE+18wk32bbZJXh8XUBjJRSp6KX0X6uXBAHINT+5PTv49BwKQGQaS
qpY94jSyMkUc3qpx13HwUFWSLWsPfr98KhAZTvV/V3iQt8Dziu1l3e+RVkqoMEoU
XVfiokJs6WyL1YgyiNhdItJFVGcDfSx4Xgze9ZN/3nXuc0OIP1diRhQ4M7x465tq
xbx41+3t5IA89C+/4VUzcvw5BwZa5wkePLdVmu44s/OtZe6BExjPZkNEQnRNftvh
cWswRMLWKATa6FwLePtRf6iWdfVA5u8Hu6O788o/GUqckBHpvLEOgEcJgyR3eWIO
HV3KN4b+RJBJs/XuWg6zTCAUaVZUFsIusInX8bPbfIKIK6gTwpwN2jzzT9E2OV4A
3FqzNZXSXoVpggfDC8Nl7VhwY4unxXFuK9RMf/pNSPn9tpkS3tFcm1HZoq6WH4yY
rB6SHrQ5QaaLzfpuQB/JHekEhAHST2PgWQP9TxqFDO6axlszSyAQuhsYg4VloeCP
4osZhtsVzskBqYWpBKk6VWwOmUflKBij5MepQ21Uq2rUtWVIOmlq/MrPx4XP1Qfz
UJ0LmrpegrsabsKe1ZO83B0j5eJcmJrP5zDGzhOZLBZX23hw5EYPUsd+TnBz1ihC
2tcYmtLzRdQPKQvDDR6f5H16IxlyCY67+VFm5Vjh8HeiPGR4DwoJ9ZAbXlJ4ceyB
AMyoCAdQSogDzsLeaLpnZZXCKsWQpKko/o40EXoceblGnv1WSswr2L+OS0em0mnk
u78AWBkWIobTrK1ksZNaYrXo6m8sKIbRyd6v2+guiUsnLAp8glN8xxgGwlyirYqw
5xNiZT79o2VvfHg8DC1MFp0W0py6p6wNzokvqMTB0RnzCVu3MJkToP3ZI83eDhnu
iTHXMC70toBbKjdkOwW4LwPbPOO5KZoHDYliEwuFbt4ehozOnjNeSqF+cp5UFKvY
Z42NiLJPWH+wHLHDvXKvyh17eCiqPiuAeOk27+jFBoMoD77I0bDNfOSbhLqmRT3C
KCm9wqBHT2EVYP5hCasuUPlchrHAqCl2F9EuyPU7+L5MAaxOmeUspYVSgeeIDWJf
GKWXYRiQfbDpWx6Uzk3Whn7sHJx/lRnorMigJbXr0H3SMTTNOLFU974jlH4aun0F
sN/Z6Z4qgyJQgEmAVpdnG63Pxgv08r3X3qrac0Ss1z+nLYnAJUO5D6J9iFRzy3pK
4+s00flgeBLB4Tfo2jc1AhaNBGD0HR++u9OEFbPZ6h2p5QZcGQTjDtBhSvx6356D
iGbQrm6SJop9kr9OrLfwkvCqioTif1bZ8U8TuXbrmopkruME0S+WzhN6HAiqbcrU
OC+YOIriAds0F0BztM1xWv6YaKRTwqn7xUwYvSh3JbNUK793brjhn7YVq5xExtXH
TF0JaB1P68PKnfOdtfFu4x1WP+IiPUovEx5ShlimTBtznzqH16qbQwJNSgvEki+i
//7Gj9Orb8Ty7qEfSkh9s0hSd3aP5QVKPXbe3+N+3MH7gx8tgqeSHGkNuy7wAwXx
T2dfSMb1KCbjDrwNnKav7CGhoYieXzSDEnxDa09vsufDV9oM9tBa5oLTryB4vBNr
WmtrBgSn9KN9YSbl/mEPxnEDLgbuseMwAGwVPtL77cOuUdKGtAqdGf+Bb2l7qwzW
BFa9GGVdYfXxtC9FdCuEwlWp+K3zz4Hx+caPbPefWI50crW6GQkEh19BzO8mt8Fa
/Ma7VJsCy5pm0uLhcegrJm3N1HlMucKiWUJkM6xX2eSAl2oO4nogf8Iz2exyduFM
g4Wx5Uf/JJjsvMq0dBQk42I1PmkfnVo2IrVIJ31E5VPgPJUyILiYONtCMmT/dj+m
OACwvLATtHYJDZ4xsA50zb4WZTn/tNNtSUUlezk2+wU+lrfF57ZODvOwoXbltDMA
GqdFPTRrURBY9FaX4zjTRgAWjqfarqh9NJu6OvixyejiJxMnlh60uDNMoM9QrQFy
XGbIesABg8Fv04XL4b3llPnUHhgaW3vuUAN/WMAEwjfnyQOuCZaJ1SaGTNDqphJM
vszASoc7YpIzvEHBH5V9oh5Leb/dLQNcAPGs0TLXuXVIMKsuBsZj+reqIxf8f0j5
r3W50+CVVbZ2V2f8dbxmIh09d3D1Yc9O22ZOezKO7FQlo6nTSC1RVQ7Ck+PKjnJK
GOv67AturHeVWPIog2jpyODt7cJxV01LvEUgpdfAjxXBPf1Qm/BEOY0+9SOW3TH9
4ub2GmIOEZw+8l7z7Afai9XG1d1oRgGA73LbVm2HCri9LcNY2JkIqT8Bm42zFDhi
WIvDR9GW3n4KLec5To/rDgz+PqiHGsBylAd/9QK90U0pAqlzXgW0MNFSb/Y+zQap
vbnsIIasNkfY9HnP+ujOAAo1JhroM/KfG2BTNrSKjyr7L0BOFrghA9LqX+IyYiO6
cMgQJv6CMnT3SzrUeVMFbC0PsCRpZthmRIjfAThIgbSWOAcsNxl0ocIMmA71iPrQ
fqX0asrZeFhgnC3AQwkne9WTQFk/snBcx8tG+4Adge3F3vLni/j8KG2Um/SBF2eN
fqFGBSJvk3lWCPS9/mg0wKVDrX9MQul5eIJLD+V5l1JBCZiP+SAsADotvhSiyLJK
n6A4enotEUo5zxOxCndbXw3LCIZzxTmTg4aQrA2oy9u2O0dsySXvErBSsOdKO+4k
y4KVzUrpZNsPoOIle4g/PveMjRqHEKMTAIsWFAaDaZ+/unQ8Db/gd9S6h1yEih51
8zf7hz26kys96jpZ5tKaemWAREGLBju8i4C4NoGaxEOuw95QdVVPJvJdiFHMdFdk
Ikwj1kNi2/O8i733ytR1OfsQH41WMlUI0n/Pcs/f/NP5D8E0O9ZyO+SAEXlJJc9r
oJ3OWP0/j1YCwp9RxJ+BCIOteUC9EK9UQkaC//b66SUlXfvsLE8ReELb+FNWCmrk
KdgFfIVMHybWYERQhe7TW/ZE2vLocXLIxBXOPFtwdrnzeHeSz83xcb8aeIyxwYgd
JkjnFT9Tjk4mR+fKqTNkjj5lRHlnWDjyoK5bI7z/1NLw4oj8W0fhU5w0CZrS0N1r
i+jhWGgog38WIEtQ1hkITUUqWh9JEnDxBnKV0fAXbF3A8oE4Qlh9m9rEiOl14pzQ
O2lpi1INqNVnKfg6eM08mT7J1+GWG2vN/zyK7scLEtu4X0+gRjFMQAEPrW97HDZu
c3qj/PdwHrQqlOWkUfhIJrQQf7uwjRKXKx2YvNK6dbh6SVRcwbDvlxj3ZDDQ+jx6
bSH0HgCMhewQetS51lQe9IHx4TM7QAU6w2/vqjJbbN2cXpKfS3/uj0BrTv2SxgyC
sW4YpBPT+xvUfxsvU+tPZG/tbKNroFbuyc2c4I++ryYwn2nBE0Gy/5FD+G6Poqy8
iSpEzUuzalrMicWybTUHP1xzODTV7PzDIEYEo9Ml9Xo6htwVAg7rTr5w/z/WKRSr
kvcUexY0ujsm0RQGbJB2N7qB0CxbH7PGRwZUueZcvEGOiE2y25By1VnKXF/Blec5
K6GeWn07YKzV2Od7H8/lJ3eOWx7LVBnlOVjSvHWvZmpD0FBu5yMelcoW+v4NpAN2
/l2cwOFO8tmTfPTFSdM8XdQVdW22I42l0luMMWKTLRBDX1XpoXtx8gB6/oKk3vuX
FRsrPM7wYpBr+vGQN46nvRcmeJ1tuURKSQEZC9/Kszutgaycy63rxmenJxYtydzD
VLWLadr3uu9DFy66ljpWbowz0iEYDcoYpOVsuQ0MYtZ7l4au9bFWQpOeTAJB+tgu
4IF++DhDGukrXXWrThCqPSZr+bcQyc29OZYqc/wPUtvWZ4lp/o+SgRroDhjnb9Qs
S92+CzVd562uY041qrcoRsSqj6fBKuxdzWywkG0LbrIeMgU2+oTivgm9YvvxI2hs
AviPzFD5i/O91Kka2gJdy/PRoIGyNXuN+FfWgp8MFBIq5enIhSJd15nArGGHAShv
yuDEH28SWF8/AlfyXY/htEjXmRLvEX5nsb5xdn3kDeSHr9tC3Ha2P/+pGWhRtG6P
3nI6URH3E06bxCfy77dIHcSBNnOxBS0gq2wOJXDa+Q+66oK85IWUTAPL/zPaWrqM
cRbrMCSQ8iwHOMiotiyMicdpM1qOE+6RSpC+pW8FxJFh9tWkCdRVucqwL5k1V1iQ
X8IBvMTsWrpW9byvSqw0AHgte1o1FwyzxFXplRey7FkcMZ7EZMtzKBcWPJ71n3Jc
EhkEEN4pR8nvSei97h6QtSDCbdRkC+Mm5mSny2zI2By3OZE5g/ApGLjy2ZzTREG0
jVQnnz7IQio3UhNvnKHDUeoJ0YQzQ3WFhqEGqLnf6ggg9cWT50KTTxzHx3inIhsX
EyU45ZHWwJPOm4r5SVukZQxbDpBVKMRJTL0I7HblYjUy5dtG5d8MC5tApT1Lj/yY
kuy4RlzlQA7VLlU7vNPxezK77Vg6OAHs7hLh+L1V9H1C3GCTY6dhKgZ+lCg7+9n6
lDRHNYWRiGJ9V5xBfy5zMos30atq2qh5VyFEDNDDth6rov7bdtTMMeEBPmVxKDXH
HBIat7FSJUVmYqX3s3t+b/9R/FmYI3oUAbKVCXYAUlFhtrYYLNXv9eFXPAafA5ii
g/k+kZoS3uuy9qtpmCjErdcUTYjEosvUd0ISjRNXZzegUVZZc1wAY5w26pE3Tbem
7qijXhDEEU+IonYXX9lfKP+AQEv7pfTuqns1nrPONmHtQlsvUmgc7mgPWFun0Ies
Hl6+DveIAlpObM4S7JpY0fhR6TKIIJnw58MOfqFvLQEKq3aFxPCqsE9nU/qTayS0
y9yZhTqImARss/EvTGD1DVDjoj1XVPyikuttmGF1HjnOzqNEStnmqfD0UmDIpXUU
zV+6QP+69xvxX2ApE2mjHXy/MKADdVZxku42G+BVuJpZkX/dCwcPVvMLkjh3PDjD
OzwFT0dUbGu1zbiPUnaQtTRkDxrlLgnKYEFQwu4VEPUmWZ3NPY/exAmlgowYDaAa
7amwFe4JmsdGzKbTC7780wiFoNXMRF1JxQU5fc2GJSxmCoCefEwcJ6+LkIi6MLAb
CvHfxXoLt15meKOHLRqYJ3NcdE8cZHN06cJb6CAm/X0eqgBpsFtZt6Ln1fwpjMH5
qBFpKqtV43sj/Jkajc3xwRb9HmncE32p9gBsl/gVZ/DabrZxxWfVzKTo+621ESmx
a0D1mQEhUBUqhr/EXzo739ueSYMqvngKva1q+lF58P/lYalJHx+ta3qxnwAPXLEl
B7T62H4PxVq9GkPBgHPrCOxLLSWgQiZU79KppT3h0Jtehq7+JsaMWGCgVqYS3zq4
G70Qbnv/72HXYASVhS2fPN0tRDFgUqIFO+4pN3X2H0AN5oFAZiqS9NiZ544yHUj2
NdMCdIOkmfba6kQ9kgO9UBOl4fu1mND+IzHzoYuH7tk+hUd4aKis+3gJ6yK2/ps+
0PrsKT/NyfxDKwvJMajBeukHPujajjVt59mh09H3jhZThP9SqVWq9V4JZvee+Hd6
LvLAkFr75ub5QeAjKn/sglRYIxtybOV3TYbzRVMKNITcWDsD9/x5u+vFgmv4TyJ1
9vsIJlpjTmY9vv5O65GvQpBYs/ibkdi4nkSqFsF4GuQ9ZS/npdEmV3/b3JT+ry7C
UIgiU7xGBMh33Suwk2dxOysqmICtXbmB6QwC1pyXr9ghwDmHdaEgXf0nYB1ccpNz
Os+lKWDj/ABQ6Pr1Nus6+5ZIbDf+oLd5BkQWEdnFwCIMnXe9uEfPc+5r4ENy3l13
JuGoUqOcsoLOBTjlVliadd+afXWU4nXry3JQ2A2P5eG7BycUg/GS+Dqub+Yve57+
m2n8AjOxAYDVrYdwyrzZAoEuSlXow5FQFkqaK4spoVokMopkiMrtFNtzO93soJ2T
9znsEz4gEi4p90KjMky7nOARwCt6gEDaQNZrq1bRQSfv0s3ynKBYNBssyWKvYRt6
o6SOY5yZLrRWpjlaoZlIFIkQx0ZYsjfOZKm46jNq73HHjd7zEsgpCO+4/0Vagos+
OXy0UpuXkqsJaXiyYqxak5HEuTT+eMEN5UgBcKLSE1QIDqIBeSPxIPcyCa3Tv32r
2kuKPxc2tOm3aTNiXgY3jGpQTC9ThPUGTHx2xQBCBFW0YScZ9xiielP4S9ok1bT4
FLx4zriPIY9BYhVevhnrkn/PcoqpL9rNB/B/22IxgZhfDE735d46XCu4e9KWaWP1
uHzch8S3SgNNP0XpyfIBqCfaVaJBE+SFGnRmINt0AvOZenHGc7r+gER2lOLtc4Qs
2Qeot+0ReIiok57Xt5eC2cKPPFYwOR0D3D1jc/VhsidD8lRy7HUdj+R7C1rJCdV9
6upie+qPpX1V7LoK4Thi4fZczQ2OxrbkG+b2wB6I1qPL8Ek9t5rllyqToGuEjGfS
Ifl6YWsVhlplrGNb6jHgHwK6Y/IpZDTS/040PfYCo2q9pi4F3oVF0bzJL51dycnI
/K8GKCMpUS5ZuOGUq0ZqdQMSySLgWX+sEKW9ensIt3qVPwo502oIeQLLJlGcDg37
jA6AAtzZ98Z2Dh64QFTKSc/MLVcXh9GLev+bCTCF3NN6vfYmLFXjprYzLXr74cO2
xED1W9LtGgxxvgR31ZRdkBAu6gDDJV1WcXrEITfXV6L3NJdr9AM35KozduIiPZ0u
GllLPSlfutD1qhdAYY0eiiG4ScjiV6Q5pg27CLrMfQDwGYyCZjLq4HyvDA8rbCTV
vPcYSeC6nICiYHvLbkK0Z0oFS5clYzu5yE3koy72D6Z//o6hn64LB8fLL5k2Fe90
Dt4KRQlFmI41RVca2nCvf+hfV5SAThbkvlIcVApnhOLGBidLpfDqS6R4/gZpRI3q
qkPpwEc4/1cnlqBEBGZ7XAkTeyw6RtNY7lnZd4k/XgaiQQrw+xVpUmZ3dRFC9FLI
TRjrm3WvgR4d6+V5JVQdbm8cl5dxPAeX1y8lA27SH/JOXj7O1B7icvvVl8DpKIh8
fXDUQ1uMN5k0/TKQF5ZdnUxdvuoLFGaqgZwV+OC1t7UggskRPla0f4MjGEeZQJlH
2paxQgloE62tnQW7Lm8Bz+r9AjgFFYOKSopQxiTfoHssAGtTK2Hpq+f93gLCkwea
oxayuNwCPAPga46aGPfL47pKgEJ41sIiTYKWJPj141sFlezQrUmC9slAyx77mm+G
WhO7sSD2TGk9u6kQ0aCmszbuVWfUTl7krJEdaNj6zsn8QBQIBGvnlyqM9MeCksy1
dPYhrayVvTzH2UAI7Z0NodLl/qVSuOooL+3HqRScTxXdXvsSW/G9RQuY1Q5fUqhQ
TtusBT74eUNhnT6set9OLp2+wU7/degAAEnWw10s3XBcIjpunuie6eHXDcN0JX+n
/a0y0smY/oSvZuqKV96QJlzVMgrMvdKsXQQxpJ+UDSBUBJieG2bZR6IKDdpUruSa
sjFg631SakQ9vAtFTMEHJV6OkVSB6x4nKZgRx7Fc2jW6BO2B4EvNUA/5Rhu7EBk2
qeLTgvmJYoBYFrHvn/mryxdbgdHAFEIcPsrqFieBEQowz7erOFjXZ6cM5dXydna1
H/kW3pyEZ7aYY3yVUGT7bI/uezbzxOVXqfJGWionSv990IpsKmsm+44mnMOoDr0J
kTKl+Wg6Ua1bAT39FHkphJxyun0DfYqAV+QU8PKVAx2NbUO28K+BwgK/EiCx4vrm
z3xrSF+DzNF0NtyIHAEaj1i349f2qjK8FsLauCxQbM9sTBVMcA+FPotTEbm6F8EP
krZ4PMKAP7BdocObJPrbe8Q/pezmHEJ0SaCT6XTyK2DZ6+NDk5OcO1Fq6e1sSR8F
holAQ/IaCdsQlHMOzvb4FmvknTjQyEOrUWntxAQY34eRkBXqqNqC4YbulsecxyIy
GfySCao4ds2mSVwBDpBq8NWkKiCLr1lq2KwObR0aDX6wG+5eqiNxxYKoO1kciD2y
KMjWjLefl9MkQ+dXg6GOP571TznVjTEDz+iuZUeuu/4ayvg2SMem/CaiQral0CE3
orIrcEDvcaPsAJ9XNPGXfTugchue4SrxhKn0dx3SlI1ea4+FaTw/17mr+gH1zC82
pWIWCIkGIVwVsw0+GnZmgAbjJXibPmi3SKMpSKfI3p9JHp8KbYCA9bg700NSXcsD
Y3HARVwDyoZok3Sj//+yxfeIPTuSh5kUuUaibJWj/ywuZsYlC8rlqGaXGSe7c1/w
BN8/RyzQygcDoNzcQfOfPJ90e+oQuhdLYgfWKrEJ7JNybqGKM1XuIOBGv6pqVzz/
P7F34sl32VKcl459+ke2MPA0M+2OWJODMr1xOSyryVSFYLywBA6z96ciU6IMjHbN
ZLWNdvh/h7+LxJXCRNe4CJJYptpIj2XUjp/t20NlLwrQ3BdJd6obKBPg0HfmLULK
NahJi0fv3zQ63HEAyxRkGufWuoxEFb+ry5fg90CMnI4rLii+Eg7uexRGhxx+raL5
7TEMgTrD7ct/tB0V6WS8/OJ/YutL8s6cAPzyWC6DbFtV/rdx3y6U19x0XB4eane3
CPCMaefWTc+ao3G7u7rFRPwuhgxoiT+etmxjMpwXNnR9wIQ+CM/IktgoMG9yogZc
JFmhS4QYRLDSfv8LmqwwHV1A0zrR2Wp0FPdrBaeGX4XBv3QZnEEquW5hkKTqZFa5
cujvfXD3RtobGOhnW6Volhmg5SXMa+A0wJFzbJnpNyQGaGwNh6oxpVyDXX7KDP6q
6c5grGyy9YXIbTua13J4NKa6i5BIK0Qh8TCNf6LPvo5KJLHl5IZLQRfro7ttAiRx
KZPqxxe+Go847HKTuAoVS9+Wb0UC2HQdlh4jnIbaoUWv1n9SqhmYNySnvoXohVx0
y4kPWj8Jc8cXK5WK8GnG3yHa3CON1mQFL9arhHY4W6pbqSCDvkk9qmV1gctUDNBm
byYgsz5iF4d+1B8FvjJg6iZelkUYKKTzEvuY5Xfae4ydScYe6sMYL4ybm+f2lMtl
XbiW+pwrf39q/MAFfkUD0TZaqpbHOWXVfCEWgvgNCblXqT9O3Y3zbAbw+JNuJReN
CUf+HQsHbMayu7hFpp7G2UL7OL+K3ZoajYA0dykOq504mmjoxPLTGhr9RDNW582k
/41RhwKafdGUnKGwcNu3CveILk9Votaax8nEfehwONkyX0h0QJPx3QIQbTV7AfEE
8IsJZEjOipXf1t5YzOTEe/p2D/72FpBTZ8ORYJKhvbnKgyAlHgQnTHNLwavoWPRp
/rHzWIJo4/Eq0lqLnpxXchxXKmG2xYYvkJJ584PYdKkfJZ53z8ZJbnRdGdeotlJv
pGtlQuw6mrSoESsBpj8k2wqs22YPTW/QsP2OGljJ4iaUYEnSw0QZr0Ih1nyfO5cH
J8P0EzTvC3oE9MPMIDtlDmp2ex+VrnWhItXCreXLvsMuK02oFntyx0VK2cO/kFjH
ol102YOdj34WS+RH/U7FYnvpbg8Kh4UkcEFLpxQebYlj9+uGvszaR2nmGWofZ4QY
PB5ZPIB9uaqDBMQdPAVO6jR0eEM/huo4895jKKso8qGeNNROMZFFNbb9XTxh7gzr
a6a5ohI7TOwQEioT7jh9MT5tHZ5dMUwGTPfkMUuLVvYslvALyObRPpM+S4Zm4IlK
ebShe74Qbeu96pUptcWNz7kQagQmSzpj+6AhtM4OPTRSu7UTDt7j0ngRrAPS4G8N
ekvKPedfcwRV4qUIoXPJYLd5051TH3sFwscbFF3aCzrzf8BOTz25cdaNYdFzBNE4
W2Gx49g1kalBmUsifwgb3NsE8dNrNUXvrcHl//8ebPtLPlaG0+cHWMEdmEfTb90w
raMN3purYxcmKcj8rw3NmBsIct3yM9tT7Hgt3xzIw+5wM5t5tPRfnFRQRQ6C77ky
o6uxSQ/ZbFRuIfl/VFP1FNwxN8Gv8ZUm5oRMnse+MmErhpsrMOuCzU8bc5OY0W6C
wbQocqYDCR/zS1Bfl4o6AX4xnV8VaQhfOC+WRDzjHcZAvvWnfn8O4OeY6lVTu4GH
dKL8fIHKaDC4JK/Q2osJo15GHBmRjIhc9OrqewuYwT3+dBtdfTt0H37Mxqf6HFrn
4q3x1LU1G1Do0jy5wxMMV3dtQlTz58RI3BRO+Q3rQvS8xafe/FITU7J2V7Z1wx+/
CSeqQ7wDdWaF/ydI20e/ty0K+G+8ozXSvdGW7S1WV9pZeNlo8RpZyi7H+ugiMc64
2KtVoydXxcTf7x5+Eark9HnVYADBL8KVA1JXGavoO8w/ku+0JOb1V2jaZUcY8h+6
mwVireP8XfA/2yIQq5m/Y330dbShEw5w3kVpm89bj77zZgVqW4FBEP/+7tcwPW+N
LSFmOGT1pGR38kIslCrwuBg/daj5SLmrYqIriPbSUmlT/i3NGrOKdeZEZs9TPUNT
gzXWCNQSC2YdFdVclsE44wL3RaIQmj4QJ22P0Dz0xbvvO0MgKOo358TO6VsAFZqX
ZpIZbLavgPQ7TOh8IGyWtnG8J19tvGVdmsTyUtAnv7TMl1lP8PtYhGvCXGCykwyZ
3wQcRrqmsN1LxiRzg/f4of+lp9jx7g2Aye7XMU63e4ZkY6fO8d9ahjge0uIJdfIQ
CdG68NXoqmeNRyDsoxt3DaGzzhloQ88rUOdr/NQ67uqMuVuR6bDfDYH7nlxUwHny
JIFYoSvgPnp7/A2rk0PedUqRahmpZKhvy5r8hpIarr5k5rrcFpx2wDmWH6TnMopf
a+SSpW7n3HPKsxiKKIk/GsuDkiN4y1yx7hZazr03qpaDJKfjQI6pXCtEvslBgQJ4
ojqBE+TW2uXt3SrotbfPK280myNnZFsdDjnP14vSLbDOmRFN/NrKbzOriAsnOW6a
ihgyds7B4BD5Nw/YLqqRvwt9VTJos65n2/cUFuAgLTUduJ1mAVAxZCIvB1LuhfuW
7KkzDims/Ixvl4difMHtMssTro5umZFo3EcwM8DcJVz0aM3Rnd76txm5mMGY0/aS
RBkxfjjI4+PhOugy5Xw0l+kabUjpjZC2CIFJfUro910esr5irrshFvYDRw+vGoR6
0xKbJc5/TVjzHhB/cv1h9F/6r6ZAXxPXob5buY5LOiej6JzjJcoarSub7c1Spg4a
Ek0DE5SPwTaAwma77ZTgcne437ytJLNKNY2xzFbeIkVZsA1/f2E6E9i+m5N6tm1p
qxgxlXHdD197YjRf8xyjTOJA0L6aDNoQOiB8kcYsOZVk3+44LqETO1KF9CBU0XqI
9+Dcl5dFjYxR5kMxzlNfqj8olOL7JfQwIFy4u2diEhgGWeEyA/cmbwIK4PE/S7Ck
zqOc1FuVhPBJDtnZLObOXoFhHem2aUNM3OJGV/SajCX+jC3s2FWVr2byANA6cVXF
ENHmTzv7nUfAgb9PhhAR09alL8wWfPoS5/GFBUQZiFTwEytjbiEcK/9H3OklFSNs
0B3RoNkRBlUPxRtLWDAc6b1yZos6+ZnOhcRCJAiFxihBXBHcJo7nizGJn3l9BWnG
sAtfVFt5XEjghG1paiIzVzJh0hX20J+RptdUBRAf6rapAaEAPmiCV0elvP1FCHIZ
RDcDYuOixrxuDg2lMPM+SEL7ABk49ULwn8xxH5Fw8KuVNU1r5Ty+cBrdts2yi8Kj
7MKkRkIaOKLgwERSe/ve3srRQLK0IMNiY6pnH9CGh3CApxbAnr2l27yC0D0UwG9S
ZJXn0SPj0dbmBYm2Ub63RXxxFCM/1gNTZfhRSlY9Vq/3INxWPXYT3rrxsuXDvEIM
xs+m8DGtHeD4bQjqh8x5AgOpSpWtp+ciW/MJQsqTn/YG3E7ILa8++qnZgXCzvpSs
MO+HEyuQLG+cVBkP7i6i4VBOrsG3CL/hO0sK6S5FK8BjIlEHRx/nJ2JFaWBv9yYx
gdBkzL/erd+mXhN2nLNlHKW72mdkvsDYFcRXy4ujRXdB5LHtXXn7A+12isuWBYIy
9Fq09Dlnu7LgTtTRMsTbPr51Axev0MQrpCJwPvUJuOjSYfklox8M9bHqGf3O19b9
h2hI97FGmI2oBjuNV48IU8uH87QbboZBSOnuV12+z9ALMizBAgV7/deoHQcIIU05
KEdw1g1IZbVJHD1rsAKIgbLM9nNbfYP9wJrzzr5AlBEz1BDs1BcmqCjBbS2VJrYs
ZHv+YZvS8r3bbA6rOq50H15RWBfY1H8KtsE1/B/f29m7SX0kmfCmja68pVLXwT0C
5TaBMqRotTzQyACb45PqCYAsu/7MIQ5T9nHhKvGIQnZo0UMxyjrNcSwD/qdClkid
S9R4IhRfw1dtLJsfpSjl2DNCdgxTCzvWUoFR5HtyhI3TqAx49HAUijvDAk0xlUQV
/n+y607UjpuWSiyx9UcOTrrY77bXz4MpJkPDdhsdEHiPWJJX34/5AXgXE7I/Ztls
t+NRFmx8no9f54OeVJ7C94Org+RbuNp7c21NId4DOHAA8rlDffb0/EZP6M6hvcGL
txPHJq3gQ5TDhZQ37PWa7A77da8puFHLfte2VTW5ZWoxIZnVcjclPq2FBANePBDT
PMZ4lIWOcoS939NO90dz7hOUvEGe75IF3C3jR+ZS5NugerV9OLh4nOreuq6vrAvH
a8Gng/LCeMhGkjDivRiwvLs/KYzCF0jq/MuXOBIFoUlONiQNM5ZtK1je4gw4C9Fe
Dda58G0OjLTZXJeVclHXdb9vL1T9YRbKESQMvYTOFilJsXgo5AaHGLObUjpQIklP
eLAX/H8JOXTIE5ajy35YLqSuAWZlflbzblxCDwx0mog4GD7WcMQiz41ItTzOO0P7
e0mCSN54uczUysEWQ+NIui9/SzVGr7e/Hx2XYqhN6RniRHfG34BTvrqHiraEmhgF
gY9vsgVOe+cIx/SMdcW1BSsBOVNj1rzsWjMkupQbibSPbB+4bsr4MPtySwEZK0ix
sg8t1N1YiHFk8nHMwFK90IXQFf4rIqAE325uscA7IsxVxzIHW2lD1RskEKcJT+Yo
nmbBtLGRO94FNldFmof6QACXjWVMFTEU0PE9rJMjmmPwQaVo+yUzZX188ERMQigZ
+3IkQS2GfsNbE2QLFMZEYg4dMG3lPEyCuFOUs6kKplYNUJhu1iPElVwQNNCgIjXb
iFr+L+fjqhdiwW8y1iPL+5oT2gu+S5wq9F5XkrFg9oKOjP+L5WNF7YeHwwNPIWaD
j55ylQgzHpgKXxEa2E9mJPHWQA6vrmK8EzvmYwFiRhKen+QtBDE0CRnuif/Xtxtd
1zlGAV9KjAML/4pJLiNRc5L8D4sYGZp9KrCBejBAKVyIg0XgCjwe/vPY+9EBxj6i
EGRyrRQhoqY2EmM5gYFY5zDZQ4SFF0b2ZGfq1XtAxsJnoLrP3IYsKfqBq3bJ7uTF
hNKNVJKPUrDv6qG63hortNzkDsbAMxtQCeTqzNE1WP7ELRD8PuD/XpBFSYHUUdBF
SCaobsMknZz3YA2kdjsFukVH27g7QDvd6GNb7MmjtJZKpt66ryAOjVH5TX6vMJEQ
bQOTjL5QCtlVbIRbmHSuWZVfgDs2alv89xtnE0G/5o85Am20ZObTI/0Ap4wRtNC4
NZh29L4DknQEe+eXR3IfzNGZLSKSDBB0IKgJn0CnNQpkqvmJdzwbw+9bvhN1TpCD
SQNvxQqKctANQQ57AXVIF1/BSaACrf8HOI2ai1YIQHdKAiM01V/nCmEN/rqrUPGV
PAXybLex3zgbqJyw4FPvl2LyIKPEIgjzZoy1VrJc9Yn/OmDnIQlsy4QT8DzeQGt0
XAWLMWbjG0LVHyA/HlT+U5qujFEz6d79zndghqGD/jUR1zDKWwrfWk5STJ8w77qs
qNumRxURn5DPxvwyGw+x/DDUAiij8rCMWWFSnd+pIH6Xdtwp9f0nXLMtcZ3IrQ4v
UbTxe0oiU7BU4VXndc8rLTD5eiDSmSFqn9YkxUWh9ExSAlSVvtlT914X3xu0cDF+
q2Ik/NTgzj9E0DpU/Dr1fQM4/IziSLCgIKfmXpsflIlhxIAQqKrMtjax+CV4qzo1
v2LvWJeaDuL9HHCIK3A7xkMpBRSTxMgkClK3xohQ7U9zs716lfy8t5gkDgwQ5yF7
iykGTzZJOcMkOFdHHmwsIhbPXjAJGUY0rjRev+EqZLkomGtwaWFugGAiAoJyZUZf
SOuABbjXv2/s65Idjin6AVVvCyrbW48+ILsndfYIkdUM9VZJbwJxQvHsHjRN/Zhn
Lglh7wHEgRgaax6jkwj412W1p8Xtqzbao9jaWfq3f53TadFtfsw6lVfvDVNTr9bb
IxYA6REjBFkzdf0qNw3erqnYxea3ZwnQ2ICbcQMzGIiikD0xFwxkSpN3Y6T0LI/j
8OHcpznSJMRaEUO4P8Qn9TM4NIDnJxa7GtU7AUhbbNokZ6tFF6mNDC84EKl96aje
XXZwK3YBu3TPr/+motSxrgclubkFs89k8gIL5rchkWLNedP/U3AA1sr38Cb/G6R5
UUMTHUIaoFvGTITewE0j6GDGkFDcLqvkHfwRmbl2T6mnv1Fr6ol8B71NsUvpUYUD
cqd8/k4RKnkKbLxp+RndoVe7m1xpO1Zp2HCROWw+AwXkyd3LPtE+cDP9cQffGrgo
Op9M6v0dbvgtr2ix76uUsRVxfYp2QK5nH2TQMPlwB2VMiDLNDG28+MmlWeTQ9GxZ
45eHZQ2y5XGCYMOCmDa87onFNSt4OChkuHcmlgTSRu+m6W+8z+4/w0bMGKl+1kH1
hKu1E/CJJwUC5k63M4uZrVfqQBogg5OdmbUuoOs0xxip6vorMpLcPiQeaXn1956Z
hGBoadg0nXV6g9ViroI9o1n2PfBM6b/WyDlK+PHbv5HRMk3UV/N85+eptMJ/zP7E
h1WDPGT1AEcdbowI0tjtuenqCF1RnRh0CVozo3LXk791vAbw0XLuzdFs7fsMOpbb
he1dE3JOTXkMtvsYIypxjYu0TDX9VTyfehnp87EYLJyE8xENzrsExIGG1D/whQ7g
kWqaIVgo/zRM53ctq+MSexByxpmL7Hq6MfmFmGBt9MuRZ7MXRnLynF+byVwM3PpK
VGSYMFSlQypR0vCB0+B2lst6I0EC4QVhAmrT8viX4oAt6o4goBZ64c7oCnliOacd
qNKWMO0npAPsYvXGhzoljGLUdtMVZc/30wjVfZNXe1tB5dx+y81+qXUwx8bqg6pk
laSvyzt59lyfqp7uk1LVAene4P+w3GZr39GjhMH+9X+E2bBgel3H9rY9Rjd8Zt87
A+bRUMeATtPFKh1j1Omdh66kE6Lfms6RowbaN8nOThFNNHj9wCmySIm9lXtlw2qi
lwdwfMp7OJoYgzMh6/hOFtcA205yExYZXBZZrHKAm/28437ISSl2aEO0nFa3rs/1
DFs3sCRn4jOvlF7ja4lVdgVAZec44/obCg4QetxRWMHoNC/ih80quBGLbV2onf/d
MSRS3vyY6yhLAwVCdeL3JYXFqfPZKCO3emroVh/wqP0R64kRc3UBu9VSe3E5gHh+
UrGxX2TTADA6FRgn0UkXhPtGQfPhYJ/CiGcFwQMS3iOo6cfUOJVJrQBM8bPcsucc
GZbBfH2UBfDwgBMp5T5zdP+s2SJb7xrgxQig6MqzItXM+NbM06bkXbspbYteznqQ
Nnc0da9C+SSVp0fiE1Mee5L5RQrgt5m2zeqy5AVsFvrsVyasdQa+qdwl9qjTtyix
FSQLUsd0Yq25XKliNfBBZK+Y9dBnsZ0CvWJ0/KC5+bv3mlrGSJ2Wd0pOf+4c2C20
rShq8e09Gi9wpBtaa9pF+OHqdOK3L5IX/J1PclQLX0ZSneLBsdlYuWax/Ticivzs
KJIXmpbNmHCNNZ7Nyov6f4YRW5kKHSHk7AsIljAqZONxXHL9R5rsVma9GfpdS7E8
bHDraCNX+LpF0wReWwUZu9k3xFrz5MIu6RaCvGZXV88zGtdbWVfHuI7xeoPRsjfK
IeY2N+QjBohRugeqQo0f9Oy2lPkRsTDcSlAcVd2c2kdp76lqBCAUXzGJFKJ4C2OA
Q0tZHqAOOM54rhMe6PYMBTv7qWx1Rd/0X5mxRhES4TAKHy6tDu1EERulG3cZwFgg
VTXiqFdv1HKg2ax9oMCS7fuTaWSzqPL768VqzEij+onwunaFJthZgXEVcmrp1Olx
Qv8naD1yLS0iHiBwXzEUWh/S1MNZCv2FNu0kwB14mEHC7ufu1XSb16amKwz/0R5R
hI5PeRM9T34XsyaMGHCu/cxYv1lV2stNuXsDWxuRF+LIri+jw4HhsCHlhBv6Z6T4
G03t52Sa6ZaNNRX/pkupLqr9beQQF7/aOyOqZmMQbJRd/0D2X7DBMlLmxOrzrVyG
M5KcEXrcnRvu/5i5AMK5gy/rdqzCmq+bSVHcTGz5biRP9Kn046fXPwlaHt2qUGNf
TGgDAiuLdbHhP1At5LI5iB8evpcVnOLud2z4R2F9CCQQyLNb8cHkhy05vOT+5GHw
LYL4AaR+/Snk0HpugSKSN50Y9T3/dIORpamm37IFPHDxTHckoW/vlSRlU68ObPQn
PG3cFOD1MUbvcIYniUfLI0Xdqp9bjZg1Gwzve+NtN8waoDUpvpMb5Fy7HBBpl2UY
jTt6fFgZUucJm4J3If9LkH/V6fb9FuoBTcViqo8tv8Kf08brvX2Vl/1KprgsLBaD
lXl/rmN5kxdJLtip9Z/XEMlTIoGdcef/78nNBa2w3IucKgnerhq9qhHLD6oNFo1P
JOskAh9fia8CIOTcfY+JjNQGWtx+0ZQimWavqn5nJlgdShp5NCvuv5rH8B5EZf9F
QVrcxXe4nMMp8VpPIuh1K6VTg/XtFgDIk4LxOX7ZtTCq0oMFijS4kDNu6oqXXSu6
G7tvXcsapJaULy3JAHgkc3vLYkLCsjIYPbFWoqWBU/YWTkL4hvg3QGgfDUqriUNm
8/TXlmRDH4kUZ15RH91zhpwNzPfpPba4MoLGpYSNhLwzdC/phcr684CiPdFCkg/n
4cW1HR9E9j8Pcby9lhf7FXCcDhxiS7taJoPee9OmKoB5GJGf0vywOCh+SqbuvspK
kiYKQLx2nCyLgne2hK0UooPO2K0tR0R0lgLsJLGrNCgV9QzXNi33DF7OwDyWWLVa
uB1iKdrnU48TZBQOWPwIWfjzvL00pwAKK+HbNZIVROFs5vUUDj2ET+JxG51de4ds
fLY/Prp0k3EiHspK9TYDXapI46nKhY/arx8zQOcf+kQmk8DM7dmkWKgPtc7o3WEy
OsZ4LJBifyXkrN9VICAfCI3v8UbU7stJgI4Jy7vpre778J3x5hGY/gwPPLblQFJz
UA0Yu8UTgSjhzREF8UGky6GV0scFd7FHQdsRmAiQvi0L8BHuo7MOdlPkIXfJVmrV
ONgUGntsE7w/TGRM9Ey2f93s+MlNDfqE2tuqGtpJX/uxfw1G2csGXVsGx1AfhqFm
uueInvmwZ6mq4BsQsSdoV5TarW03ZRHjwlMgw67xWZYhJGcFUIBKVQdwWCmLEiHa
SsOk7IJLcdFi8bx+hcI9Zv5ST9AbWM5bx37tU9XtKyjWB1GR92qs71ltKMCbZwj2
807s6nn2tUVpRXEU69pUfZGdRfwpLlMu4rmMH1DlfMHM7R67xiaZtvCkffj18ys+
bkCUYM1kWI3IWiYQsH2C5zyn7V4aoPk/pxCfpGvc2lQc6m3bHggjsvqtGhGnQ8Kn
0LrJZeqXvJ4hGxC69pMGWli2nYGbewK4XfsN4DEMbvbsXofsXsWHkM29/mP50/Ie
f9vbhnsUwbPA0z/oPkSsimilnKjmkf1PTuvZ5dbRjn60qk1XVm0V5MWE9sc1Sd/+
YbU7ErodyBQo4V6oDCP2RTjOyV8SLCU32TylOVyZMo7YdaYlOGYN4ecAWi858wy8
IG5rm2ddnGXD+d1HuiVZyW2CFjxbLMEBymructAxUS3rGjGZb7+Geo7czBCPgNuj
t9oV1Ct2wzCqncXxYgY9MuMJCIkiLm5+p4jDjnoUbCD3qyU/Dapoupkkw9Hv5oV9
79ilwU1Ihsp9qZxjaWS4PyALkOY0ZgLl6+cRhnRvQURonM+prvZult2wvq8cWvOw
4g2m+S2xA32xDF1goGvq5drAiICy1OTgO32c86IvD+IkRqOIM3jnZolJcM8+0xAe
K5I3a0yBdjZxeVErBMaDcdAXRZfM5wLDsqn2gxokNRrFI+/s6Gv1Mc8cqRY9GZr4
quABdQBXJUBTcROHbk3KlhIuD2yuxjvQxLuOwmi8mDh8jKuk8j23SFWS9HHq5pKT
BHqva/e9Tn2z4Kal2kE4Y0LZW6TKX41nrTspJe/tpyPNIuiO87+Yv1OCFSwGNvn7
EMiGXNHBIa+GIgWpPnYm2k2Aa3l59BS2nL6cUlC5AFOqDxsLilGcL2pQ5AgSWk3f
kvKkZQu1RhahqjaYAgrlA8mTgkiX+nXl/MbNYjtT1CH+8ntx6wMz/G5eYk3nxY4n
ckdVuG+W4Za+ItclGCzkuLD56L91TKk8rpcvBP0Ka4z50HXdTl1k9twArXsU7iR1
r9ruZdFIVFZinnPx6sUeTScMRqo2b2CMVNSuMeOnX9yP9xnfLWB28jRs1qTdr2UJ
6xI1x6VtN8TLjej4EHrBl9Ab/alBht6mlsLlc3UnWQUzJyfO/acjzp8bu3yUtEZx
3Mu5vtPmXqu4ti04B3RZa16JRjEJ5eKNCDwRq2hedh/Vh3KHcQwJif/yrsfMjzxo
XsufLB8H+kTsFIuLfOygsC874rPZDT7sVK35PQ7bw+WLjPAY4BNwvqOINCs7WXsQ
/Ol6s0w1rv2aq3js1xrthrlRHSuv6pLWTokNZJlc1SHdG8wsVc9OAvmhH3lSrjOG
IqqD95ViNb3rNiE6try3Ktoe4O+aOAhubH4vJyzV+iInrg4phigJHwVxcq06zK8Q
uRaEKaPSV2oOJ7MOHB5hFh0QR02K8OnMif3mY2mxtd121l7j+4Ii4v3yi1uijIhO
YrxAq1AUrcc8gE+sl8YCk9tiq3IJvc4AuZe7Y3+EPB9D2CAzqq7fhpZ7x0B6JzsJ
p1/+wSiFbJ3dgv8LTouLDy/FqN2vyS4FQr7PhKOYynR7Wms6nT9u8sMziS+2y2+8
mrGuCs+JeXI8AbQQ0Xp7xR1eS7Cdjxmd0NlAm9CpC37LGnA9lWeIuHYRtmyTYJPJ
0SJNDvTFGhRO90oc+ZMYzgEDRD9rTXC6pC9AGNjU42RUebrYWEMWJ3UeglSejKxm
xqF4yYotXLe9HB88nB5s+thlHbBhu0NpkNLPrVLowQDkGsK4NY5DWfuL1Dml0ivX
Z0gx91IC8FiwzefPQvKvxX8xqaco5/tjLEQzyyt3d9rLlY/4WAoB3qiaOES4QIcP
+MlYgo/xmhv0q64T0SCIHhjUGW6PxIKZ4L5vOcqQU1NvZfMITz+REwTjM8o1ysDE
H1aNSJurzMYTuIfb7LlRBMD4+OczC8iACujdEjs1tj/44x9qa/nEHcAOeyB12/jF
niKHWy7GBED6tJhUYLqlXjrvjlLlQDTnkUZai0PrFwaWrPXdo0bxWy42DsUzmiB2
p1BxBqQjKj1b/icOCYsCjHs0VUyYvoTKagbH8hGbzeQ3lspEhd/FQQudXYGfz/sw
RJfg3LJLpnv5ctl4+0t4Vz5ZbgvnynQnJpLVtMWNlVj3kTm6F8l+nkQbET1A/c+7
6PAR8fbQWv7XRl4pTSebmw60m3a+RgWYxLdfoemqqQ9cbvm/jb/wlVRyTnuYTWKn
FYcfRF0XkUTureqMoV21FhqNYlRjdJ0WtWHGe4u02p5lP8G5Gak0822d4AezLjDl
QBUeAHoYzU/Rwnj4Jz0c9ItoRR/Ah01tHDUwEIjTAfvoKUshVXNvjpSePAR9kSL/
f0sFVb4JQQTYz1tK5IUVe5RD1M4zR4xALIozooSYTxzdc/JtcIxd9UNJt40g4/RD
wlScqjI+THmMM4YDXQ05RN2eOhPSnNbAAR6DFmUlW6cBCZ6KwezuAk/I4wp3YH36
Nto3OBpmw5gEItkWLfy7LYBaZMXp6FU1s4Sknsr+7gn/7rotHyEjFkyx5EhQNhXJ
Hv7irZYAOraPx4b3msfyyDlE912iUzPDDIhJL9ModJPYHIUdIHtm4Z775qIL5uIt
tMhVb8ZIHZgoGrdgRc0A+Wl5rsMW5mqnwAsRXPucR4FF1HFxgV4EhaIl6GU2TxL9
hlSY0qA0XqXtKUge1vexYBPiiSGT4BievzIVERwoqARUu/pFS1M6UW17IgWGHQSK
iUN1QPrHBO9IxOSq/dFaWKeDnQiyEWIaRYmKk01Hvo2VyuMa2QVoZ3lbfwuCfS0G
G/SKjmM9RvFig2j+Mc/J0/30ID4QVbyjVsEzoDzUfkwL6AIFGU4/jLkb5vFpS285
j4sh/skFnTXr0CxtzIUgIq98GXHiSDn1iOuebjXDezhXVG2uxFLV5Y6991B/Kez0
lPiS+aAbgqk9fyfUFb6Y26aprCblA8wHjyfykkBsH1socVqy04vAryeelF3YRSLL
5zrmOtKOCG2o21aUGjf9VQ9c4rfOaU2OSpAXA7EIFzdye/2t1YaCXYr5Gj9opdRU
OAWjYMifxJLN0i3/0fJqiKMMdUDPhIkInKthHERlafHV8OZVyA+kic6YP6LVctDI
9kdDJeFT+jfYfsUC/kDKuBBiGGslHhzYxjlORKOcakIZe2wuzgiZT5yQI13Xv+Ac
8loYZySEdBkYk20N9FWXZ21Zm9r5mN45IwFqJQTCp2ANjc9l9QF+lsD0BWvCF3HR
RhhsM6UMTqAISn3c2q5lg2u50ukPOgO5eJGy4qr31+vq85EoYbunMsL4ZdSBG8Ge
wCR4knphBF3v2bLH6uFvF3IxzBrFpkFoQBOcEOIeFxQ8zILW14nERVElGEDdjBWW
z52t7snavXNhRoPcBM3YSK3G6KooRmnpd3o+6zqQyDXHbaGmPbnkXV3XlUH4hNaN
kbrWJx0t2X3Vpna8pfKRQCIftT2BBqudB2AQrK0gY7S2O4QU2SsI6CPJCKCBvpSS
I+MImWHkqBHouNBkPfM3Dw1GQNOjWzGX1e+TDVPNMu4QA8aRopZHRKxk4BHsdxqT
O6rtxgSDrZVdeuifqDhAhDDHTbw8Z5cIXfoIXc9bRG5kf+odZNZEZ6pn053uUQHi
24mduwkzUOcZe2DcWDypzErxzaeeVgskymvnEDCdWa//EILUkyz09VLxXhkb85iT
D+mFELMZUn1B+5hDADPJN69+A9aW9KidyDAflccHF4cDFzX5PPbT2aiw+BUaKSBx
oXAlD7Qqes20Ss5HPW7pnlwKxREGAfqUX3R02XsfVIymIrFdzKuyxTwXKhlii6li
VM4gSTfxlbG/rIgTzfKX+AIC8mREgdEATM2/QTwdj6LiRfDRF2Z9MxPa3k4b+p7s
Z2kft5KAcrF0xB1LnfOIF323H1XZ0/txDHgJ9913xmciyFDKHdxQkwaPHH3M2yrH
c+rj3xYL7ihvn0piLJewz7fWdpxeUDHaEqC2QeMlosgVdOLmzaoPtoH3cOvnlgKH
vLypYPwZ72LrXClG7xp8sbc51sVe+KFAxDv0BJ6xp1IzXyR8hgQhcKGV9002dY46
orIypY2fOThL6TiSsvQQos2n53jehNdZ9kUVKoLsMF5/vSD6fOfKzJVkdkhFvyUJ
suULf60fsuUfeHMuJVj9GmnOJTDlkk4mYo6IGyWtf0L2hEGc2Ic9gtE3SWwwD434
VGeswWRDCX0YYJ6NpGO9LTH8uaFcR/gwljo4dJyIumeySq+vl9CpRbguAZdj37M8
0ySMGBydrse/I3m+whyicwMsjS+WwX+WiJsAg8+Ncyka+glqwy+tcwvHu9M/o6ii
BFTRWRPpb6GPl7cY/I/z4aaVXXIjeDb2pM3ewHVAdW/qsDK/gTsE8/jMPqO8V/hI
s+AWm69H4cmPzweWvZ8wuec3dYQGIdX2+dRQ7PBQJA9EahvbASa+5/KD7p0A+uM8
D3UgXrTgfYvrbXOP9P5mrQU9vU1+usZVzEpeKPm4n4z9GaFg+xtIiCXcPr8tIt1s
ot3ya7Cz7OPYmjKsXAmw1GfYya05ZQLj4wYLrqC83dsrroMyaQjzZGDQSD+IlexS
IIF5KHQ+qJXFFY6OEVc/5utuZ7xBpZNLSvFHiBGUFJ3KFYFALF4zD9vTpfkJeWbO
E8dqO7Yo9zY5hgkhKxaAZfrZELyNi9woF5z6pgIjMDRZvalWk0JpgKU5D5ivUHGs
xxAUkslLlvJIVyUABjXyiOo3p5A04adun5flgzxN8kCHjVbg3DJ+njq0xDbQCdYd
Z4AXhV+Aop0DP/MnToDN6mSWc2uVuDNrbzR6Z/ZoErDcG+Dv3ZnjlFXQ9vuP7Iex
MajOInqRS4ivHrKCJ/NHoz2Er195aYWt+jJUanTqahLQNAuRhNv7l+UBDHfIMDJC
8b0QjfuY7FsJZCTRhOpZHna/wyHFwp/dlnYVjTgC+wQwrjhNEhjOSmON8v6D6ZNR
jxLidd2boVR4BQoDv8Qi+0fyCwNenvT8UV8XAkbjuXMGAH5nKPQyjp+ZlmzUH5n9
F0oxG/66ps/RAxN8FtmxGa3rf29oMvmi8jKpL5OlQ8ZEdVlEOJycor11ip5kvqlL
Ie08QSnf20jR6kA760APrCd4hL1EhJSSZvubBrjP/JArXjufK02qimld4EykPlkj
FLtliZVz0EQT6Yh5j5FtEKwpxyEUm6I1/H/hdtIAKNvlFo+YNgz737XzwguuElE+
o8ZlAcK3MrdPoO4aIrXSYNoRT5fbcHQMB12Ee3gpB/a9QTT6iNDintqRHlmMcDCr
6ZfhrNRFjJDbr9myFCbN/jN1os3imF4tRuh7LzXEBCAw6N1/ziRK467mWiBYWtaK
BA6yb9pFFNxd0BQNLxzgj5CKkvS9AlOz2n2qxHHBHW3hhGpb7WSgwu8v7HOJtLRJ
/yNG/d58hF1+XYwGJ4AbSo67ktmxC+TS6ZC3ojcqcPgHZXCVfFmT+395c6lsBjmB
8fJPgM6Ms0aBQ9Oov8FFxgvMDhWDO7PTYUR2ylapCcqRSXbd5evQq0/GsVomz2Ic
LfnPeFfoxe+GWeQDHptFHjYsqRBiUKjsq2V9sxB1leWW9azlk9Ti4CDwIgSN3dbz
/GTlbcYpEvh/zTOwYlIVobj5loTmDfprpjrMNYLTXMQ4KBqutuSrDeVQT+ysfBBW
tWjE7AT/C/o/ymcFuhLYze0VBJYwK8gLt0sHqs3P170dbda8E/ao5YOj4f4mC7yZ
1iNtPxRjuQ4dRyTpHLZxDCbXbPYn+pI/DlQvAZNsQB5z0igJuWLHlzkUz/qHK28O
Zz0IMyXNHWC7YaF4b6iuZfLpRU3+Uw/j/Oe5aG+wG2ffPSeKunh2wIJegcmsVTC3
BzQVO/Kq0n7p0r1oTO9DczQR/D1RDd3WbPv0mf/X+oHff/eVcJYX+qTtkfNk7jqX
et98lZpqchei0EQBArAmjqPeMyIfX1qXDJ/WrqdfsOyROrid+Zie5ftqVPSrFmMi
IBOY9DZEHCRZZedmZ0vHTNi3uoO0W/KUL0XQhFNmhy7AmpSSDW1IGSwOaf+Ltv/X
xUDeCIcUAbTL28c7WWINleEJIJDcpq6j2Yv/G/F3O4qny2AknAi72Tl3ahBz/tN8
WGsDihJfEJZXqGBSs38sGSUXNIMbr8qvV+ljlF8ZJ4C+OsyehS8RAGn3GIsxIya7
Q24UOZjyFxXsOXQkjNtyvUeQFQd/YIrinGsIgsLbT/hhhaEh+YWCGg+wjw6uEem2
xqoviilAy6d+4oPUduObJviDlcWPTeeYW5uyew4h6h2J42fxf1j8fQMlO4CcwATS
oShFSe6VgCUj/25U3cdNf2j/nsE5/HtIQ1vg8NtuhUMlTsGfELs7azgbCt0Zh66B
nKwoJWiia8gqGMBukr0KsSMJfztW+GI4yf2RrS/ACH1xCKbgWHG5/ejDQ0X4Z2Cn
k4DQUk0uRhFZYsNokgufgOjXFA7IHqJs45RFfxMY8DOR6Q2cJfOTx/1voI2CeBos
JFCeosXjmH42rTBP8mS7NmU5IUlMgcy8mT0WDEh3MjrKSpRPWeHbsyZkyszxBZYy
exTHMvr7uCTtxznTO96w7egcib3pJxyg6/7mLlOwj88X+CbVoM9lrDmNQ4Zy+YQ7
pLqZP//X0o4NmWySyTzqmxdAj4ak4P0aw5CsCChpSE6Dv9GWC8CHrKKh5kvqIUxM
foOKVHxe1sIkDYVSYzEA09iFwZjROKNTRygVMv3QIyGpDEQzitXc+iLxAk9f9q9T
xCdq6jAxy7bxuGb8+S7lLKaynrAX2wg95ze9NddbVSci90i2sOg2RTM01MddaFw6
/ssVInokUbs8chNm3oBmicj7hgqTBm2E0FPpQvvOK1vDsLzp/QbI7NNPMXgu2YFE
O9Hdro2qHYqjjU4+++JdcmctQGnBbU3Eo7GnVdbJnPMTCvptk5FrFg6iIytcIpZl
JTw/IMnX4E0K3raAElELksxroxG6gVgdjgg0678rp0x4Zy6RzjoNI5LUmyJDj/H1
YyBruQ0SB2YxppSA+2xE1hjzqlbc4nHR10n8SWo88Id98ZlhRcpZE4sr+u9dCTjf
d2Nigiom2w+cTxR8j6Byucabj8UaFTB6yWJexowSDjWMV3F/bEteiRYsMOAT++dX
gNatgriRmtiFlUu3gyWHw95flKzcQp00CUJ+dqcBE8AcRGQvb1I9NgNDPY8lLFO2
ILoejW8TNxRcveXbuQgEi46x1keNYHFM+KWwKZhsD5F+eUHpXpwznW2v9h1FVUom
sDxBTEUkimmgQiBHdNhBWNtlJQS+tZm5XXVrBDgtPCdqxqs1PAQ4psxoxn+7rHyz
awiTA8qxEDTXXX42Iqi6uLRJEVXBHbhcLN2Ra5NwbzBeaIoFjQb8Zp7n2SeP86UU
LmuWEQRvUnfmZ6XTyOlwtEHoQQa7uzrcWjP87Meurlu7ELXusoFDNhIVAzCD2wtv
YYWuxp0KpAB1zHLcq0w/7i0ovF3zOF2vzlPz2Vlpdcw2IbgXHmCcFoUb2QsTdJoF
zeQTo5qETQrENcFb8ClceBESr8M3HMypZqVzhM8WtvWBXd1EmsnOd8Rw2vdBQ4mF
ETGy6VmAWfck5M84FrF4VbvE5RA683+kEcXKg1nXLDh2GdsYeth3KYcMB4ivv1bO
Y6JI9JHTO86eylX9ClJu5V+bzkRbd6YGGEKBrK0j872+vocXZVvO2vbXqBN0o63V
IOicugC/4rzYSbkx97uTotualQvejJ5bK/jiRW1ox51JBxVM2zXCmvPfzViMnB+h
48Mncm4+jWb1+YTSmyP36q9XsoFZKDxm3jPVBHGAUA+oVTuq3jvFB7CgJQg4xfQa
4KSzX2uE8/G6r5jDEovhH4NeEVwPgGBvV56v8Ndbvexj6yd2VtKSJ5EWtjJn8qGm
WCWVrxCrr8J4uNx3m2eIc7QFZ6TQTh2gZg/x+f3Di3rA/IOBRMYvg58TRCUh9Jb4
7fVqOPMx99rM2lJsTsgjTwAADgS2+yGalX3HbajDdVVejz5nY2kOI0UetjpAh8rD
aae/KMmLRQA893TPd19Oda71XWXCrXNbezGbgW1D/ICj1ffi5azhIFJl4FpOnGJ3
arwoyzSJ1i8SgklDuQMvCfmTC5acU48wLrSymPeS+3kaOnAh9W6qr9w4MufegiLw
E/gTO8wzycHsTTsqHwUiY1HrJ/55KAs2Q1e84gwrT1pQ1dk405gdlpcrUA211+BS
uQfQeWG3bo9hwfAbM2617yg1f3XRdtljQN6d6iC0IcZC1aPge37RSwgyiuQGtV2R
wIa0Dtt0c8jnU1yKbmQ+sUHEy8tVVe91D6xbPL/RxGApDZxt4pdDUavpUProusj8
0cYmrJoiA8Bu5RjJkB5akIovsxAV+9yUvtFqlre0e1JWUy3SxaYB+XrNqV/Ozwd+
AU+Sf2xM2JT2PlSLacaUrg7eoAJeBae0NlaGuINWVpziwlBLNUJdr1apMXEib16n
iUFhKqS2pUJTo2LMRaes+m8oLyiaWCR6VavXCgUiisBudZQ8WCxIYQ0Mhp8kpG9C
IghtistYLnh20Iq8JKmW2riMEOEmSJjttZQynN/pfQ0+D/rxUs8yKadgVt+FYzkH
UNELAKhrv7RBfmgyZQyFz+I2MTYEEuelg8vF42lBD9DTJOohFanEHq7IcbxRg1Yd
aGOhre2vXjWHUaLYglds8x3zBmT7K5GkiZnm56YIZwZXLpoMeYIehmLCDFHWzpb9
GGLo9E60AHsF3XC+V2jEM4pmBodI5EzlEK3FaSNxERKS4fmq9q7a/tzWDGYBi2t0
jlLKUpZcPaThEZUGe6kZyPi0jR/9sfyUEuAADKWF74iKwVpFy8zOFI+ECl/79r1V
ZSgaGzsA2/Nh103yN27zPXhGFzKx5JA7aJHW8LUAfy332AYujzJfXOQtoiEdJRHj
JAij2sbOJ5kwFQUoIq+tIN1Ul3+e42aaPnno0Hgu2c2t6NH5rAdeSwAmWos6EM66
KH/L0p4fSir6BMNO2BHtD4krNyXM4dBWKCgf896dSKjjYIsRKOncHtuQdqsIBXnv
NLPySxDgFTwiQ6GLXEeXgqlaXO0F7OEQo9IOVDTXLf14cFMfJkQerukkdHRieBAx
u0TvTmk9P9uRDEDWVsh6dMSjedOcUoa27Sh0P4WjchXx41btp+u+jclZm87HeAxR
Os1WskVEpgKEH4FbXXEWaZA1viifcKmdKnkgOMkCzb5CHsa5vf/mPK8v8BGoHe4v
9xY8CFQrAOORSHiDOBjjPDPOxoMOugfKXY3pgyb6UX9374UmbgwOA/8kepZoiaNO
7Rs50/dc6HwpjUV+qy96rN0LcVbYiZPkP22RhZS1rfBY4Kco7Zd4Gr0SHV196eIX
mdF2GFmIuYn5jbCfH7VOG31vMq3mOxJALshsexTMk0bwhBEkYkUP1m38WBgqQkCg
eKx7ZRgpreSbHUzq3du6VU9+r+P2xRbeOQ/nKokUpJlyIJOI42snhy17/ClV2+OF
C4U624GSV4h+S+n1MagBx+an3b62Dew89ZFHSrLLum1RN6BR8EYw+MLyKQAYyQsY
+QaY+5ZY9Z1IV0xSwKOUevOvqunXVJFYg2g3v66VD67Vqgw4EfH+dAaHjf+eYlZz
naU4VeUukiekgP3iHlD2q6AGYzy/eHCQYM0MI4is4nNdzf3KpvPAuZIXui+Yig6D
0ZX75zz14vX3V/WuTifziZIP2mkQlCJdLIj37z6wyj4qFeMWzfYX37SYHibWAqHM
o+CcLF60/oN/Hpot3+jUHqFlocvaPwxk1v9/04H6o8SndkTAyC2fw7YomUjoN1fp
raBuaGqhNKYyBxobeM7wAGiYtoal1bkK2oc35vbiqMw3g9NOpYMIBc8nwiJzI3dY
fgPp5oTCWq9m6zfNSv1SuCBuLya4RM4NlSBGmACQIovVnTgurMpNdujAMdq9tUJd
flGBPhsMGnt+n5qmm42XFNSk1zFtpY6vSJ4gBhr+8NFI3pdqHE56/EyCNBU1Oaak
jH8VGSXLfL3IT/Cj+E9rU/RuFPMI4x5sANRWxU1+pMbqmoh7DZwa4CrdwbWX94nS
KU45RJpaYnLrnKYSTgMBO0Hepc6dz0+h1W9gKz6l1W14+Y5pLHrH+M+nakMTR6Le
QFx/sWF1WP7R3in1T87rlF0gxijuX1FMkdol0EMDl6ZxQXNL1Jzq91Cvx4AEKDUX
3VXYENS62K5jRVCkO1qE/2NBEDX5flYXkduJHO4+h9v4coDcrVlPGKr8aRp3drB/
RnkzQtDIs9bYm4QPNLmch1XFb0amKdNlGZdQHSSj5Fjgwbg8nZwMX3c97USpMpGW
Rhs301Yvb+Imr1mkX4v5Dw8Nzxar+mAhdk0nw9CdEbNNTmrV/nKi27hyhHyCFL5o
o8cMWzCiGKyHq/b2LYElA7yqd2xAjaTfDqgisLGvKiub4X0wD/JbmSZhJVli0juw
C8jValp2935NLyo8vNr9VPfbuzDbM0r4TcRo5XtAOQTT0XInGwOJH2UiprogLqJE
n0UPEX5hk4sIwt/DQxlQzDa0gHP/15H0Pya50gF1SaL/ylxZgHjuZN2Wd1BMCRsV
KHWpzIEfuIU/t+0U47B/6DxJPzN9jX6QWI+GypSL3n1b0BBXV+nH9MvZFr2IaF27
lQzrjK/J+/bjoqIjsHBeui70BNbeWumj8f/Inef0v6bH18oC5g65F7/tVSr693Q0
wR7jbl8nIdFaaWqQE9SuL3pJBLlvSx9W/wBivKod1R3upffxIrNkqRghIwMjB2db
v4l38YTNboQ5+Dy0HAXm+i/xmjMU82oPyEr9UKdA6zeq9j+yYGa7pPKceea/PwLQ
6jSQYhHW3Xu4FUxPfvXemcfHc8ZF8aYcNTs3dc1+tG7gN/dyghG9b+4yI1dtdh1O
bRbgHH0A8ee5FLo8fdOqhi0Fi5U5smepR4G+a1sjyocnRy7uk9QO5rLseXWU9c9u
RxZHcF3EP0kXswk9hkBdFy+owBWrI5tYirUdm5MWu4llljQ/zfnwzZGsOtLW+bGf
CMf0b3zUhnwPrfGvoFYe0YLPUv/r/qi+JUf+8bXUXD3RIMOvbixtW4ECUkqk7yk6
6ORmUoxk3Gj3+pcme4DQEnN5g1wnO7PzRpPIwcHIJTrLH+d2ANRBL2D8L0O0uKfT
kFUsVY/1Zy3Rcu1QNPh2L30lsOCGPzADG6xNp/2aA/QVzxQag6RXlpTVyLOOLb9m
SQn+7rGYraI8gSuqkAskA7csEXVD3RDX+r7LsYR4AjsauBXXJsb1pD/pVQF6EXG8
x8EXSqRHTilnAiviTPmR9jIOVtVCaQgUqIuzx3HEenr7+KOKWX4CzgyRTAXaDL4G
i3FPlKZVnzJgCVUQaQT19Xuepc4vUvn2c2Rc4GrVYNhVs8RfpRkpwtgz5mF8ZYCW
udYvArTBiC5XuIetH+Ybegg27Z42e3NnREPZkMpLPfYtbxIlprdqCJ/L3fhn20VG
HHUdgcuXK5E0VKP8WfS9Aqt2Cn0TheVW5pzBQoQ/6vVQkGc5SbEJ51z8BVu2FC7R
kxs2pAvFE7VYdk6m4IuS5qhClYi8TZIHTHjf89y5bY7G1RywrbNxg5KXcUz5D7jY
BPdd7B7KWnG0nYN7yYgprA4hEK5v9f38K5D0lC8EOkETQHPoLcdisfaRQwr4IYte
/1rm3hTsd5jvn7XNyG4cB7jRQ63cokVXKbpSvvX/Oos10Okck8tLi19G3lfoKjoL
Uo+O6VZNjteM4loJwjOGlA2xMqfpTCAMsGhc1zq7+QoQeuJacr+RDzY+9x7cX3/y
20+yW5tKHoh8ur3FwfxuZBIu8mtfx2C0GqOuvPmhCWmgitXSH72QIuB483C8r85c
Nbu49aKWa3+kELrkQ9cVEj6FWQ1VM2449513fd8Fw5Ne2DzP7Nma4XGgjuCBppuL
4TAD1sEo+YWU1eeKSRCwnVQkT7u3eSq4KjJL/Nkho4Wh1243Xc3GN/SZ5c0VH4oF
AR0Mi+exQAzraLaFUmDG7ax1ds61dzfSKlzhwQG3IcW0FMKy5iwUfIVjgtMSEjks
0kVGgi7ka7oXX7gbzdkhjynrY/JGgoRtRHCBefvmWf0D1DesYoqByKYfAOIFhlGc
NaQuRhjS3/9sLdzXLCTsFwHp6vpPLX3MJtgstjsZ50vrrqeEFkCHY6JixVhZenl6
RBXBn3dVxH72U3Kli+YK2SLuIZx0aTIuViyD69ljzHs56SfbevGv3AaqMOpZ17BP
NTOsGAlRlNDLIPDqZ/VKUmOb90Cd8+cmayNO3rIeTMdFagBWBLNJqPtCOC+XIjQa
PtvZPVZrJENymx/eNJTsbcslwncxTqZJ9Cwb874RYbugxXD3V90cH2gK047XFVU/
Wbw1KTD4jCW73UUgwfamipr0JUZgRCtQI2AU0m6qp5W+jt6iIicue2Be4DoTVRbX
sBzqNIrvTCZwXw+ekN+AzENu9ABL1fgOPPX9ILSNDdmOG8S+wyd6GXsXH7ziip4c
klA13AyV9DH6xtJZv+eXrGFxFAw4cELKMUmHlKzamXJtXgBJOKfQhcMcaUOBwV7d
IxD+yRgQ+WpgQBDZc8cbb7G1LayxQGc8pQUfQR5SI6q92TqsK7woNIDnHQH3A/ub
GEaDgcCpT4GTWG5Qh9XOKN64SmNM5fc3WEVDGcJPZU8706LSBVuCko9QF/lK9pcp
giYKbd3+h9kQP/3+Tz5Tq9vjIx554FRXtFnwdC4R8v62qIFWrntOE43NqQAvazMK
s5nxTTlqaVO4AC/io3N2AWpaYNDABz4ixsxmhRh7/r6Qrriknu8c4Kqc42UXf6A8
X9jdrFBRucrwI4YY7GXDfGbMv96bwcMoJ+9XPDqIS+EUOE8zdYzzgvnguQ4KEZ0Z
JmO8TDbOgfAUyqrOzBaEZieMJ+/DVZNpEq5VplPi3yiRDg+5kqHW7dZwQV4UFY4N
8nPOi9bZI4QoStbxOezE2n4QP6Doc3JR03t7OyGSp+bvTUzC3Ws5saJc7WTlXCcl
JV7VLfcmKZ0AkgrdcDnWQeKaQRsFSEt258HxxlBppnNrRjVBsONgpdnN9WyGNKY8
vNXrlL+MhU6X3P3pJqHjoOW6r0w7KH0UPcmOnRRC7HPFVgTEUQe7h7pZyx5jXpkg
j36oyUgDl7TNlfjc8W3Lt1jsRZ05yeUfmjvLZ5PDSz5fFdHPyUMR+yZUEci0rRoa
n3RbP+fMk61MiQ557PE4K/RL1speeMroQcPnKN9jDeUMVtW6v8gXi4nt7Uuf8CyD
8ZVQ785k14/r323mVePXJzXu4lpfrrN5G0yVp4oXFvgRpiYpHDEgU2t5566ndS92
GGX/55/x2Sge+u6vt80Pvg4YCGbu7vCeEolTzBG5lVaQ3xh3OllJZ5KdLHxLGYaw
wA0JWsgFC+a6WMuNmoaYHCZtQp2RIkBQESMoc7i9WUtoj7JQmfzs9cVM08ls01/8
C/d5L9w8BUJHzyK5A8Q/LLDpgvrwFh8RCVo4DqHsdA1DIzgHSHL59w6vDjiYCtzi
mEch+ZZ4CqIPwkjMWkirG29TUBSc0yF9Fkah48PfJ6+XcF8qlXEbpG9Bjzn83Ucj
HkhIIo1qXqc0lRm0cA1psPWu4/Ng7fX5iPZjSOS1GW5XtSfV4gTkvTmyTDltDsl8
SzX6Yx2/I7hCWJTndgweZvAjWQncFoVfC/hKhlbbCh5j1YyKr6XqNbUvwEhx1X8m
QiROoG6JSo6p1zGXCP1NPenalwIZlcLjkHAr7TVTpbIme9PoijDCvsuiPMEdFnTp
WS49IdLamKlB3xv84vFg9SM4Zz6Uw786i6k1NGdY6mc4m9N/axVRak9bF3excFBW
Fwgy6v4bX1wy4wwO4KQ7IKUPIdR0vkqOTOvxRrG2ghTbVBtG3aXz9IyCEyfx0py2
116n+xQm3wPqUhqsksdWH4bH6cxg2cpxlsYATOxlTcAA4iu5VNXyG7k7smiudNV4
vRtvFDBW8aRHKb3UzwxO1tkM/4/3ioTdf9X9do4BEwl76IPhqD18XYRv9ic6mmcM
K1fH7PJnqfAtRDjCl50iqAa5KvPSYR80RniS37j3UTOMrQh2kG16N+35bookNf/Y
t1X5MQgH9RVVkACLq1FogIfWNtp3Aor0se5M4blopp3DKMmG5KrRuL3WkUzsmdQ4
Obj8M6eCGhUjIWBz3GzIIQWG51R/1Yz4B55W50HvHDCMM+Y4LLAbYI5OGiRAGet/
W222D+eh2CW1+qVGpYtK93aHY7V9xvuu/S3cATE5YNp5at1tpH7bAxPQLfYYYg/8
VkP4iNTyDY90ow8r1vj5nRK1DUvlTcECKWFM3mAmj/aA0gIrK4UATb4mCPFa4rtL
IiTIqWAVWjhohlj2XM7jFf6/owufnlJ1QZeDRn1fMjpLDnisAvXoO6TtnmkhbakL
2MfofOHvAYB5tQTh/kR6H/GjvSS4wqtyyR59HNaf8lFu4MJhSdASoPA8O7rRUML9
VZ8cF2YQ7CEVvA/I/HlqceCPbDchz1VkENG3ypMPZAEQ3uwUthTr2POl0byZZhEV
4qAFFior92zXenajJ6Ay2hOjTpVwkGgExx/fN9AUHVBVgtTtszkfygRzOKCDydjS
6Lavufda6FXamqp+fnFhF4TAW21DDuMFgmtZT9cV01HV5m59SVS6GHYD2YbnOkzU
hqs1nIIzQf0eYMiHJSRAf+cLi0+ibBx9rzCUwnhVxAh1yYZxYo6lGybJ2GlmwJOs
NmWEKMGWoDl3G5NJc0fDABhenvVnDa6qnUmNAM/0S/5cu5nSwahAXa1mcPpYS2EJ
lF2HZfxid+dSqM9JpurX/NOs57ePLz1ldSkwG7E6WfhLMbJLy1VYKuyOLIHDL+RA
QgHLynS/9Yyb6bCXgShTj2eQTVn7MwwJp0Bq7Yxdaogb7Rpb6HVwbiH19FlpUcsP
KV84y6YLveqAcipCvhYjqZUZuWq4iA4wt6kjCPTD4Uw3z3ltlmd37g7CxBnk9EA+
VHQ+DBPILhJyiMtFTlk7jtxYDCirm7uoLcgbEs9Q2Ogv5dy20TJX6q6LvlWkFCqz
PRHinPT9Om3iYfvcHSqr/SxDOVAbMT93epWNbp9oVqAw3BDL2uOINmvsO4JYaP4T
PSSkIUYHOiR0MfYWcUbyqT7XWNgwEpMHWilSiWQB+Blt14tU9JjOIAIJYEaKNIFI
oQWKCtp/J7VIszvpSLDwXpDRSri7XLttRM1hlrbaeyGo2OFF2ELHRbgqDv+/fmXp
EQqBS7PwryuTdhiOU+rt0laUyWsOd4mlN25dL4Oj6KiZvsn0dX0S70NetdXux4CL
fSmpUFuy7b8lPM0FAogH/NHx+9PVPluksi58QtIb0D9YPyz6tNAhxNSUkiZEumH5
tZXo1ONPRqgw6LlLdDUzAW6DjZ8i9GJeK/fqL2nAO/wyr4HSdQSD/KVOABAaHGe5
GvI+iVKjtcq6601yPYPitUTtl2tC2/fLoaNTMEezfv1bDxD8iAMV7aZ8gLwlTmfv
3za9WeSsjcy7FfB1jFA8cLjiEHhE6BJWn3zvm7BJ1VcCk+iMX158FnwALuVUqsdT
M8S8msgxi40G8Bz3oZ6N1v8WvSJEtNUZapGbVQcx0RVUsi91il1jF7ChMYHlyyVs
UB8lqOKBMnN5TeUlMDUVfbniUQFQlQtlEx5Zqtd9mjyWwMVkW7ltYPjaSwneXvwM
FGb3/RGS7hVBYxhUTas1nzOzOZKbShGWCTgEL/rULryaK9OjD5ajXvpRUtD6Dxzz
QvHg/DDp+PRl7eR4IZNglOy4CGldm6RXEQORprIIvvw+i+JyzFx20p3SUmE2qwpG
19Ce/0wvw0P93+pIXASQUfcBkIrtC5f5EdjDGLEtOP5UMCG9ZT3yJSDszYQ7Y3SW
7t3nSQxAv4B8P5cVsOe01OitCsojdqO0YXvYVEZ9+rvtrct/sPQskBUm7JimCN/v
1+dXtrp9aN8LDFi+V2ncmDyzw8pdO6D5kNhZTVN8WvIRo/oW7sHEHdZIql9pbSEw
gY0vBSj646NmsOlFOGWl9xf6MBAxQxgM9385oEP1VDuYGWXt5+5gUo1hhRjH7bKM
ujKNJQFsRGcnFAA2wW1Mh32JnYnqurJT57n9xD6Hq5vMoFEUHltu02Q+BU5nYUOv
DJAhSzLidU6ZWPn0wajdKsXGu+svO7wFQMXox/DgqVDl5L89VLBXpWk9SfmOjQLs
+ewkwTjMr5Yf+ymeKrRPbBpaC/53fRpPNWcLQs7uWMlMDYSObh1ar8EsGH85FnS4
mrV+y43JUpk6HmqTpF3/GJ/Xw/5E2h3vLdclpHSARSVCH+mOFr+6sQdPvaIIdr4a
fqnYaMAI6aHs6hCpe0si32FJ/i2PhmzcQRwKgAxHcqA/xwHLXr4zIz9Qkm7fzvQY
CJWPPXJlVYFKIRNLQJytTQpbib4D3Qa8LnxbC2tYZYaJtOAyZ4/NV0iNHxMO990M
0N1COcL+otv9kLxshVFutcLiOFhxCVrNWEAMj4oRwM7SNWV6n2+CZPzO0AbpVqnT
fEn2TEdpbm3cVYpo4tS4vT/LNsElGdwU8kXnY7vgae61337LHLia7CDK2NkhwolR
35Pcp5ctmEUw6qOLD8bovROVRtqFu7zg7R7geV5DxmOixdBnD2JSu3JpV2DfaOax
+mEvCi0bEKU242f8z+7Ob5/JJnZrcvT4qRXrnTU7pVf47I4cwXxONC7DKBR/n6CF
sfBDg+sjsFUSVS+1nI3b8Id1NrcQD6tJRJFNT+eu01GXZ938tssmUuDg6aRZAXnF
9lYUEHHeMQbN/imJwe1HzaKAVi/adEJ57/DuH6PVFB8NZ5RBWuhRhoospxNMOAAl
UoQQKNy1SjbS1k9kd4wsZusFvQzR3a2/DWDTROd6srFCbdlyqoNg25Hk/hHXvrQs
soLl+Ut0DEYWJrq0cnQK6gB1gMhqsPrbqiU9hk5cr5VLwMizX559Wfa+mVl7UaPp
R9kKXv9HrmBnT0rpM5Fn0kEn0Oy1ENgxe4wGNlFv7f/FKmJM668M8CST9bOEiwgn
Yr4/K75MS/8UMHvqMjYo+u3kDtxdwxNQAGoHc7LdDyKSUB7g+QBwMfusKsQWBuy1
qV+JjrVLmeB3JC5FPmtp+a2secGUm8NrpMpSxGXHSc+ucIweIDGx2vE+/epC/yAm
uwoyyS7d25b1fLz+MUdIIqNTmRMWD880LixtLuI4QpKQvXI67LVBWL+zvn3RX1Ky
SMjJ5o+7r7Jw7fDA3BLtl4krLor3oTVv+JvFfsZLD14ROOqVnTQx8gvxIjiBKysj
i/iYJlPlrC95L9nU9WqCNkw0nZtvdZET7ra4nMbcL/2KrFQJnxX+VxNUBij7QG9w
IRR3t+ZlmgYstaq3NiBY5URGHposT85JVJomX3Yr8x4VkH0YOMDrP08zl2JyXjTn
9NqOws7bw+jYCbOCBKf1XEQd5lY0Ye4RzPWwMGI89O0tZh6b2kZ/uUahW1AR7K3F
oUzicz6WjfpQpD5Q/fgK3zX5tw+3r1OIlk8Ti0QIHNrHi1hex/okS0bZ1yUJj1Yc
6kFpPF3hZXiArRSgHIirZMU/oBLyS2sdJLaI8RGXqeZ1PXoIR74h/W4jqzo42MQ3
j2IYGSaLUU1f9Q3C16BiXL+frV06PCrP0T1nY6zP/OU+ByntxJHmWCbef5LkTh80
1q3Pzx2QBWhZ+H4znZ6xEEpsGwRegahD9G8pvjTtO4p8EQmaXs1HYAW8TSO+LnIZ
XyvQ02Wf1KrBsvmEi8Fr4QGTV+ph7dW8jBLlI0+AX6h+dpt9nS2ccxww3KpgWd7+
SQ1jBaoHYKqt4ajJJCuQnl9ZlCg2zMUbwShn/GcZniEgEsO5SkYWBjMQpGGN6pnf
qc73h0BblZgXgAsW47KTBYi9nbaY9ufS1EdduSiKbWVFmGUlRrzAkqMrZS3Gz4Hf
6fqwx3j1hzlH8a6MdYce4DQMMwk30GITVGJRUyrET6Hiq17hnWQf/83kpiUv5FLg
lFA3JWaG7dE6AEThIftzrffGltUTYgc+lkarlJ932xyIYns4HH+z3Ue4hGObt+Xu
m26cqK9849kedW5SRDrAcTX+ceF5se3LLNPXsVlWiJTzBStuO4hNDlZoJM/gngVm
GksmvvpG0rwJvXtch/1xzoWr+a51VFmGxEgLkDxeeQBgI/go/h5MCa5+x7XmSL+6
Wip/GswYVgs1rKvwpp/hDDBdWpm4g3oCuenCYRUlb0uvYg6UJ5Fjt1uYhbBOMisi
8dN/kmPf34sGZlaV0iqcYP1PaNlSooBOr5gRxt6zLWCDcwA901zObBcVMaKzm2qP
cqShFB8iD+lf3hIdOPq1d7ZmtKS9ve+tQgZAvcobYUNzEMzoi/OVLy/6NaqLgUlz
Pl5FeialCIfxvmG3tf1Nxa+2w9B7eaPWK3KJHQwkwB7UyeP4mxfKPTTM17DA8uQI
/5dE3maHWRbTA5lYQRH7TAubyTsesDEr7a7WxdPaJSmtz79eMJQ1q8UYWy6YZODg
Oe3RXixEKSFuV0X95/voYCzLXqNSmERrU85tua+IZ1SmU7VLNFBRUid1i34B7fMZ
T5cc9t4CFehqoLhke34oHsVVRvHfMuLh5HgtaG0Wa0kGBvdvVxuRYmhxxuH/VLOW
cM/WXsCl21Zu/jjFxhQsYjkHzQSCfJmHhbpTxicYC+1GKYESQMWelMpu4bZDiunt
u4evomtUB2nvZ74pVSZcJF9y+imaJRiKfhPDKkLkhBm0rfDv6XTNhH7vRIX1xak5
oBr4F85YEy2DJw15OrtG+X/Xg6swpCdOynN3X42YgA564cPdp4H4sgpcFSEl/j1w
c2kBCNKlJuvBJxVPtG4sas/QbmAOYlyD0bTcnPdKR/8VufSxfiwawES6ofIImKEj
ai8yiHyJsmTeEREe7uQut4TxQcqi19fuA6rm6DFaUHV1uGU1cUmUk7ndW/Qo1VfF
3e2ZZmvcH700IDHVYtreeJIaeCrqDBn3SkLmQ/GzRmLf95fLoFtPoAavLg0J3PJ1
8tHzjxD1sHFzPYwRXFMrwJ/RljPrwF5hbNntD/j7akrKqqwZcNsBvTnZ8r8kREJ9
pX25886hwRDKvnf9T/upsUP/3uQCjmIbXFfDoBye3mTndE6dy96uAgX7o9FGzaf8
PYdJiTVkTwLhrlDNokrfmBQAFZG6ROPTJFvJC9QDrxfu0P3B6fpFdW6aZXRRCBJZ
ldOeoakr1g5f3mRNdETn70i00rWG90mlcD9xknTwJegxodEgoG5s/4u0r1ufTX+B
2wa2CJWsGbe6YwPqkHL20qlEvVgnUtbjnVXznUYzUO552d2v1z2cY/1pC+GTotvt
pKnfNxfDfMStfmCfJI3s9iafNP1khMdUQt+UhaN+Mws7ssJyJ0YRfCCJw1RfI3y2
/V8Mvuw/rqSkH85w0+awuGBx4bqogJIEqfcHH0Gp0EwpF/1T+3RfsPK6JIxUIlMB
hs/flDaKXlt/CK12gVsiAN8g+0t2Ov47YgEemGicQa4zdaInnGBj/zsmsq04AUF8
rzPNXt4YJTeFBnoWEhVDP9Z95v2LohwYIUjIh5OhNl7sX2raK3ZSHuqNbWlEtZMK
CPkNh8NiMMLT9oZ5I6rAF9xwOJLyisJUdBFMTlby/2HjgaSuOT6CI4zy8AC+6que
UW420SuXHV3dcNLC8Pan/f0+Q9eQYrf5vvjvoYUjhA1U9yS2MpQIags3Bez/qf99
ur7v5on1azZ2O+Ke6lFR+EpQ1YRH05hbl5qyVg9GDJWybOGrO7d90C20BpBPwiYl
9jbmbhe8cxDqEpsaUQRziDF2z3r0dmvBjV7jTfbTl1ccxADlFN774pPrjHSkflEG
ayXbY/b8w7SBAqc9O5kse5a9sKIP2SRLHxGLSeUdeUN8HVz/I/h2xgyPbzSzfpQT
R3EaUGMdB8nG+HoP6pJWzV+l7ENrx9btmC5v2gR1+kLMk6Ml9xUrvnhoUG6oqqU8
UzDr+3Y2pRuOkpboYOBf1bBjOCopgHPybLjWgsGe+bRqMIdGoLt9AhcRIA0NGasg
nGNfaJlZ0NaO0c8jv7dArqmH7qSM91Y2TtZhsm0FoVpTUJ3lbqfRlMxKJ6eO1gtY
ee3UABFAACK5E+RqJL0Ms8lfwxZJwnylvoejDsrtuIQbX1hk2HvmT8rwJCLDVYse
Hh2a4Qp9QPHp5NPmgaof233TyJHucoEB4KpIdVtT0jhD74ff7RrxmkB9PqEpNhoL
ZddYX/qMa2rmP1IRlENNjYZKlEyS2E2yupD0GPuWlLCqMYb0udpwfpBj55yDltRw
JVXDeEX2jYC6o+iLOUZ6t8af1u8cgsDK6RCguDvX2zPcryaxBG8hVDpxqEkui4JW
c+/g6VN5gJ0iQX1jYYgOlUhjgSEOT+gHPG6HZCWsl0nFDa5ZDmVOz4NDljc2J+Qp
rNDQimTYgPFUU3jyJATyQUudG//x0yPB7lqf1yrQ7nGn1rfTcYrSyxWT5brF01P7
ruEiuvaMu4GMC5Z65qDN6PjYvqwvo/XUyKX7/oC0odAa8yKxV5BKugL1PEo149SC
T538Tq9fa3BgOd3tqIfXVcXAX5UGD+o2nFMfTpqGuA4RjgJ4qZn5FNFF5H5X8Qtl
pREDUVCc5mOfe+20lVdj2Cdk+eq46ZM+RWdFXMDraAi81K1G5Tzjfs5gkg2v/4/R
h4Bn04aZHXFd9KHGzUaap4y0x2VQYXpJkPt+19XbpS9ZNiXgZMzs/9+e+KbzJdiA
ueXDzUUYFCsxpnejRmIrCa9daFw4kqukrr9Gzvm8W2zCiCSTz3eJAglDuqTaallx
XIE3IWUm5sgMIpz5Pwf+ApT5GzXLrUoHbuMMP8IsjvwTazKMspBWDazlx4eLliMQ
siLWZM290N7CJ2Xm+dI6QmwLsxbi88lCkVKTZ1bOr+2A/gxLKtm/0z5TwJiwVVB+
eFF/P+sOkgrZ9EgXx3mzdrBRFcVJeCmkY3RCQNqfYCgL8YmsPvYtE0VebsZV955o
vqtE3fIoQkK+Dd46Z+u3J9ZwWBA+CGsKwELCqcg5IJ5nqlDAiNVdfntN0Skzj7L7
y0kRLpcwvWDBfJPAO+AyStAFEK3Gl5Ap1cpb6XnFZ6cyEXuIuzmIbEarX48OJF7P
lQ7bAwUiGQRp3scWwEz9wTCDF59JJ52ExDJnegBLfLFj1DzuZk00RiX+323siGSi
QTF1AZJQMENZf/St70AvvocZv5Y8DFsDYwtoPa9lx2Tv8sOUHyXr4YS8WDXNrDmr
38reYAtJf5tOhlpz5lNIEhwlOMqwpcRJ/Xgb1N6qOFZi7woc/Ib1UqsdRYI9ZYsz
w3UoduWg0Dp0fn7kBw5UfMXyZC7zzh8Vn+fpxn912svExg2zMO9B5FMfc482Vsn1
H3sTZ1D88hepGRJMGr2b5SMClTc1hzn03BO8J93STluf8jcWofZuL3rciq2xmaRP
mHVXBIBFGkqdnaSxXtzX07YHQwponzRt0usQCjqSKUleb5oqIipHPAPQlBxBqDyf
Ysx47OfDNWC/ueGV4obZGEckR4mZkG05kHWsFBWauMeTKsz/q0UXSBW8Y78QolAX
2ZEVAtw/0guZ61Y+X9Sl/R4foJpSj8ngNw2xNiiIU1TjbqUpETKZM3r8QlHdyAeV
qkgGLSwcjAUX874x4EYdQ4VKPYv8EwKLSEs4H7wXyLRIhV4UDofZgYwMnhD5a/Ca
ZN2vL4uEnHVrHqV5dd401d1rYVi17RSsOe2y9mmS3fc0pWYKR7LiRAeheiI5XTk4
ygubnZKU5LYEgrvX4+73wSoAnkDFsVTcHwLA8ScQQPJi7xpzs992+dlACHIkKSbE
qfF6eemkzX73IA1Q+qTfhJU4sJyZ1v6XDOSejBimtNUEWW2y0DAJ361CQtEmQ4Fm
gD+DC4Xv3aC8Kkl571qdaSRBk/HjiSb/yU9Zdk4eW4s6L+33FQxV9XJDDdHyFH1M
aqmBy4I7e5gVWV+32U74W0QcvLEQWu+cES/7orAlU8bFYChCPdAioFnWUdHVpVmL
0RbGS1AQoJBWvikj1jrQgCgEVjW+y9zv90Of9mbGT0ZYIqKPlvy5/rQh27epZwBk
50R8+ehaOyMk9GjVQCQxWLsFonIYh0bXMsgO84gq2huVRGx5D6YVKp8iki5IHkH3
dlRaGz7umNq8FyCjgE5tzYdidDeL4hzXpOz+vPfmSvcvUhMJ2mYEaEEizUxFZBKM
S6HZs6gMC5PyhWV/7ALsoExPX89VXxRgqm/kmgMzAdAOiYtDZby4nK2nADoA/4BR
R7UT9Mq1f6wm/xX8gZ54eUI0+C1DMH3y2TwkgrKSs1OoG6zcqwQQLV11CFM+U6RJ
Xvyya1ZA9usj2Z+vjmHwFjqXqSulPyck6dxMa0FaSiJjHoSpqRi4Hq07eQk94S9m
MeJsy9cHzEQ72Fi8s1m0dB5ubTPTabfF9fQZtZmWG+jmCpJ0zS20uEDYqysmMFqb
K1vw53s3FZv0tRkIFDXluuYdiHREcXRDkS/hOiKSkAyqhuy9Zc55a3kbJ5i/SyPd
/ZYCuF3OL1qlTEr9pWmyESq+cyorH89OyUqpr2ypBnl1/uiQFl0Y9a4zXNeUr09V
ozFPry2CnVlHELsYIO2ny5q9vjAxb4t7VIBpRftdsPui3ZRwmSBxArQHVyEEZbSU
L9OJBQkBvb1uXoBGAaZxcMI6wJvh35XNLHttaOTnYWvmrfHDzioSL/O2XFoPXSPn
cUQNDhZcqr+2YJ5g/qd67dqxHE9j771oSIS1FMKDyq+xEido2CnX9rPi45sx9rPI
0dzslu5YoGYQkyLcdcxRuZ72YJyvaG6MTzNeC79Te+JIi68JUQkhSH7GmcpTLK0s
+j0O95WYpxFVJKsfeKJIX0VPlNoijWwzRo5QBtEzH6+otNXr6U1ZzLSduHeAXINs
nGLade/vXZ1hfNg09JEZpuJGRVxvpNFRFxStZJNB2Xo3zXCh386bP5zyIFmw0OKJ
wxb8KtvY1NsLmHL60rXp+NzvbAVxP64qEtndzX8Jdi7vsH/4lLYGJLEEStX9f4pP
HjKtrwWk3MSvlY4KeDU6Dk+0BLCl8YwtmziQRTjRWYigJoS421zKEA/QPoqEhSZT
iAVSCcStQfdWaiw670BbGb7L943axZPIU9EtWmgtZ1b2VUWlGwsFgyS9W7VpVmUf
JD/Ih3kDjEyqRvNdjQ8OgHBA79tPw1N5chr0rqcGYz+VJOVLUmOojNZG6f0p69Na
LG+RBknipDJlRSVHEQL10f98SIXfd2gVaQtyO6KflpWJnqXSBcrxRL4gsFfmy1rm
ETJSdG0yk8RL8Q1F5CNR17VQQJeoZ0vKRSc6Ogj6eFowQ6RDoTL7opbuTPKsCrPL
GrJKi/OeNH/s0WtQ9tAlAbmvY3V38ePwzTU6QgCjTb6KCWYoSVDr8LXY7PjnQjJM
gJWxq0scwEBL3f8b3eW9kGN10pW+t3Dpy0u8eFiXryHyUvZmS8FIoHwOqljlklu5
xuimSVygVn7hmNv21wacFU0+hIbqxqeQyaja63DWdH5Xv3FDrVDcM7sJrTcpS3PY
+LgOlV2P/zN83ntuj/H+FFgbxIsPZm6a8W3qerr/x38rNK97IE+FZaVeWiNnMllx
hTHHR7hiX7EkMufOwU60q9QPoyjCt7gMzwcRdW+Xi1PcJ9xRPNioQPR1tg6aYxCS
m2y5FmF3gcfVg3pknXKIEDWmciZH5jsHb1ozKfqpaQScXfT8JqPJqHxoHePsy8L8
5gdGkTDcpxVy3W4AQ0kdqY/28FPdLFX5/etsKE9QCkxw1jqi6FRKQqYQeye0UItN
35Xxm2ONE5tFjkcUof9cPaPscdICEm6gHRSfLk+9T6S02VNZr0G3DAK+SAZX4FSI
fx15G0MPYTglHoiNsc0bgxlAwyir8P9zMB9UJJeseGwGZ8gVHvQCx1Dv3cZNidG/
V5BZ3rzyR8i/isJN3PC3C9GDu/7RdyBpZC3UH1lHTWHfSHf6X+SRKEMZ20OoachO
GErQhHz16ZRAbxtsg28zDNN4d/Qbglaj8ehT/g64OgU2EaHqApvHiVHhZXOiikuR
roBbg+ywSehi/9xYG+RUv97yleCj3anAZptkrNHE3RIZdo8ctjDJUVocoExKyvs/
ovWKd4yoE8lB8SVUWSdsQ38088afoZ0ghQsB7A3yfYlJ6I4CL4c3G4F7Nfx4UYSh
a3FXUXJrIFSD8yDtnrOOCxj95Dilv+P3+QiVZGWwRKsOKd9PdxDlKS3X6xhS154f
cgVB5Q8z93rEBNrQwFXgubi4qonrc5vezDBmXcyI+ARAaqdBRp0xl2vzyV3AAyWA
udHJ01YPc3Xf46zKuFcs0rXHwJge0TM8vDq4LvUnMDMhak/CQMFQj39Jq5DMQFVb
QW0fBRZbie9KlAgbGo2+8hfdwFdKoT05m5qXOAEgXzF1ksdmj18KOpbe3hTZvujz
gBgegI9pOyQjeWF6Nh1jKiSPhUH8D+BP253IF0pVAMBGe12yXct0WqXCHidlxRgl
uk4rk5IUGE8v3YynW7vPulqq5LTcu2xco3+FVNzqhRL0B9yQLTfnzjAQoCTGgnQ9
xr5xP+vK3lF9KUZcoUpRVUmBeGCp/9UauLCqL1c/lVZVKxWEz38OzDQ/laISmhsA
uwL0izFCGt/XOJyqZT5yj5DNkH9dE6rc86iq7NHXfVnzxuifp89XAiKTlCZl1HwI
o2l1ek2KiSj24gXowvr/cdViBJVJrzaGMjmO+ogfGX1+8v6JVv7xKwlhWXkZiPjL
q26qcFrBRpe0gi7UC+kie6ODo/+a5SH3l8Tpxmm/PknvWa87ohC1lYAJFHJh8aB5
RAHbCQi0T4qxBxHQMKQRMtWsg6VrunlPOGeoQbzmgIyQ9OS72cRBDgsGWKl+xmEN
wsk9hAlrxizbzrgPrZq2vM650vOWEtExm2g/OEAIXJpzrzUkPewrpwACS/ZLwS0y
YNmu8b21snK+ohfxuPXn7IJ0/tDjysRWaTGx61kwsMVGERUl11Jujok4NUJU1X+B
RJgqCHoh7KXueUv8fAEqQP2dOK4rn8/YeAW3kCiDzBTidf368I9LBJ3CiHpg4W9o
ESHVPS19Yo35DlM6/H7dILKtGjMYrsB+6FxlV7UANbnsfXwiY748+z06CYt94f4e
94m8Fg4vZXvYYmWvtJZi6l2Hf5+IbUXlfmH4ykbZ5Rx9KVMi1+LBKaGiw9ygTI8M
M9uICEvW109qGkzvm4fBpw4hQ3Dy9LmI1WHnSC+jYn3Af8fw7RRri03Ugt1/UYmb
Q9RkTAbndaisTjDtKJgugHUjZ9N4tyLyUwexDiyTcyVTaca7KtvHKxIe54UASwVu
TXSL3wWW7JqBMQHClv4HypFXs16ZFPmP6yb/r0qEkPq/6SMYp/9BBhRFPZfLPTJ+
CI56p1056c29w01trqyMMJW3oDVNcpElS1xaUGOWHo3bEaO/PKZSlLtHSfRNYJgq
04A9O5AnTVQDwKpkLT3EjCkmkYwqs2DKWavH5MO50d5KzvJ/L7pSBHXz9/vGCbMv
bdEzfw2KRqYLuPO1GaYtCQ9gWKboUE+edoBnggh+FbjdK3rmNweKgZMPPQdSdXOJ
0enNGoC1nub3FesnwloxyZ6SvLkW/1Ixyj0XAsigk8k80o3nFjeuQj/DqQSJO0dQ
vDkPOsg/UvHsS1EaVSKC5X503F9RVkuuioy1gHZdYDNn+BDZTR9qZqvQf5dHvPw+
NARvRYbIU6D28VP91zLBj0CJYF5BFzcS/t1VEmREYxsKvKTxawBmdrFtPcslZJ2s
J/3JzeoNh7UUnaWS5Hk88ahsbODPwxj14M9QJTuWkuy8IFbUKdbGTabRYi1OPZuR
TKcSDH2y/jAckyxVZZUZhCYxJOKA/B2gu7/UN9si4cjfr9NzlIc5CK2AldV+4mY6
a2dDGLpXUMvYeqrXLXJlnRgCC2wrpfYXHgS57+A5DrIGFHuFrNdEAGKVhmwoQYd5
8KL7I3jL5OnDpwC4JKVJvlJVXulDdd7ELL3Y09LJ7BOIElYeRIfkNED3GUiJlKBU
8p/jjoqj0jPMdk50FUB1gjEbotc2VdL1zh6U+ll2bJNowb2Ste1CiVojIGOqYwCR
SBY+nZiEOVu3vLX/KO+rmOOpOo7c1oxun7zyckvAM+3u/IQUAclPwT89hyUmc5s4
h3PmmkGbzkccs7fXx7FIKGwQAMyfWbArVKDLnriC6UUrBdOeIFnkvaRkSlzz/nHx
/mu9r2MSJpn4uGApzZC1VzhekrZb6X6Bf1BMX5nIIW8bcU8wwV06XdWwvpjapY/s
qW6oL7Ko2b2Kr7pxlTBPvY6n17At9gENFf+kQJXqvyUZ9HoE6B2wJGUIKVOeaE1t
+H4XGZXxJ9o7GjMwNRkSbW839eMLtSlpYv2zQwMQ32Dq2IElrZA3HuiwHrS6awJv
zxt/K+AFfwI2Ige5B31ljJ1NQsarews1+XqFH0dY3bgSERCbq6DJUtN7O0H9FHue
KtKMabPUNoyUrj7YjPkBLQAePpM7h9eRNzQWI2GRugRFMT5eoknGR65KWRzsRNYk
z0Mghei3qG0DWaywNEB30KzihyaFKp9+O6Ezc6EbM8Y0En3CIwHIBW36eGV73mYI
iDaNdDTIIEMmule4FrqUrZfREgdK3MRqk7Qyd06/h7oW5S6ygh5nwmdIOeNK2F3x
WFGbpRLYRPzUSSgqJKojGPG0XOVraWvGjqJJZsm6ytIwqPyUKG3zv4vL5aE8wBF5
B8ofslTrmoR+Y9YyuX5FQT6e+1LsB9jh/Td/I6mKY4jBgoUiRvB3KTxMB4EPvPb2
pOlPRcKsdYgdR7FGVUPTegVnnhyzli8OLJfSLCLH2aqxNa7/GW5yfAfHyFzSmird
onS+6pWxftNpm574nJs5MdZoXl6sNfRblalC9FI5mNw01I43KVfhGDMnBAkZZEgs
MCL1Q9MvbPk+HKPu/yu+PF0VaS2KANT/pDOwb+k5NuTjH80groG2qYqdjK3GVnsM
IRLglRrZ7jS5T/abNjM0PAH3/5rUezF1Qgz3gKd3PyIanZ3Y0HxZk6zYXKaL9G5j
G3RPMkWm/zIa5XB4o2u6ghOxOY+mwpPl+B7NbSthEn4gZoKYvBcOmemtVeRM4YzV
XAiZpKM4PZPxn/L0TQnCoYbysRLg6FO66dw2sOoij9Q87I9htI5LjIICzo15SIVI
oU0iIQdSEZe++7KsPgUEO8sGPVL81WlPUOHB/yGiQAr8FaPLMmu3LkiVzzewLq6o
oX6qd61+IKWRHPjlN1hRV+PQLNFL8aa+UieuS4yuPKx+tnx3lc6pcssAVWkue068
fO4rOfKdMPkX4Tkwo8ivEoC2xkMjvk2aQILfpr8hPn/jXL0LNTsjSiQknqnI7/O4
L1r+bJF6cri60H+HqLQwTMrLJBZDFwx5GlpanMHG6U1r639F4oZ6ZhvxgCc3KNAC
aoX9QyH9RNQV0BNMNgoZkfqVptGx1DFUtVJG4MpkmkCE1yiTuE/UDDCGbx91it0m
DmiRKic35RxoTwUMnXsktYMS6LxsRYAzk2kHeCF0m8hZBn6jDx3aNiWmBhLvm4qE
ica7F7V/9pl1sKYozOoOfHJZ25jry+oulCRnypac3crhfn88mVux2UzucmA0PKbO
cwLIFYvZS7+lWE/gs8I+S9WPoLB00KjsJEqJaDH06h41QyKY/IE7eMqhFirOJ6sb
mIgpzaMZaGyPJj+wmIWNqlM9JJQK8kA23Jhrmp1vy+l3uNJtPbt6uxEvx82aolto
xtbQb8m8jgjeFyRlQM6yrnCdoBz7//4iF/Z3TZhRsZpmjJ7PMYTrn6E1UQPeTsZw
3GxsyPdhBP8wY7v0ij8JGSwVD++ThhYB/BQFGCHehyH0qXlYqOY7brGHI4sLUmdK
/BEdUZINHVux28ELWSlrAFrQMtDTzBvx8GTSej3UNjBuDWcdcmTwIeDBVaYPasIK
Cry+r8XDyaqCx5PegvkBJIkVJw12DeLNyP33dkLowaO7Btqns04O1yBxVV3ZFfxY
3w+YROXo1CIPLFGIGCV/v+ebJnoFS5TyfcKN6DyzTnnkwYhrfbmYekpbVK+QrsqR
xlV0+42DCXaxPnRX/zH8GDdut0c6cBQ8FNiapR4uBAd9AkVTSWyP13uEdqdf/p0Q
JgUFBx2AirN/nsMuAMf/STXCU5CjyK9LzCUfxy8iOdoCR+7imEEY4vOQFY1CYXd9
AITMky40pPOUYts/aH+oBCy7pKeC+3BuOLVoOKB/Hz3e7VRG3MZjf03zSJM9Stso
QX56te2K18k4OAFSfozhzYcV1T1QEZzLowAlA/S8F/VoMLYLXQPmfnPiR0opVGVF
GpOTwB6Q3iFPdTLj9Q5a0rgeJmiYA634oicJwuRpn0PVWTK0Nk0KUTKxVI6vahvs
0dwPCs/eyDysilDqBeBLNBmTg3VdzE0G22RIKwjw2oSVbcz0cOQePqAyeMSY4mKu
ijEqwby8QyOwX24R4JUNy285yDQXWUKwmUkuyqf2WUiqqP2ZQrUdQLRqC4fsFyU9
wvk4chUo6n4DdTkuXrmVdLlt9MN6VUlLuqe3QD/LPETSeG26F4eLNorM2IXumGRd
ol0cR6wYUtD2SMtW7W6F2qnHLI9PyWD09oKVEij3nMogOh9ivlyApVYCpL0D1LjT
KAT0htFsJ7uhFZONtBfGJdcUOlJRXjSzxfWc6PYFii/jm6+gBXIVWKO8aiNjuqmB
S4AzyBo7AnWyKBNSkoDodHmF5K8rZ8ZFpeNbdSeOAi7qLNjyAMFBMIomaO3tH8MY
/cQ35PXt0Hsge/z2vSjc/8gZ0HYtvUx26ZxrDg1AwMN7CgBojn3q3+j0WhX/7e2E
kRMSSPt6O8dOS8PZuzl1MweklHaAMZkfNhgVRDCtHb/MvLgcU6uTfGKj9j4MJdIE
i4PKi9QsD3u64bXn3MoszM+o2EymQ20nDzVouiQDtmILGI2Y2k/f5cq2in3umyCz
6jab5pLUCOgOkzxDAnpewDBxpYn3PdlgRrl6kD/1oQhCPuW8mrQt/vTtZjDloKyG
ByaGxqaomRtc/YByMhYr/BLT1R5smNt/MVroHsbBeBWqGT5ZgkaA1suK2UmHgvKT
Co0QmHo3e1NlfHsja9Vplvv/92YUbnOgH6l34JpIPb3nJagiVvhT10lfCmoZRGBc
2sKdUClMyksSZ1Z6QSw3s2puerVewrtDTbcx1ak4nhVVnaRbVyYGI6PBTBoLUzXA
tu4Mczt8YJL6wPXJj9u4yeerdTLL09JPuD6SKBwFJJ0h44tRVeM+R29PmlM4Nafz
OUwZrUoDSFxjhgwkZgXQWSJCK3lxWVBrTKLb/aLCgd2LW7JH5FLFvYZw/cpLBEsk
qXYHBzY7P38BHp2zhD3Toe01gBIt/4pshYTBe6kvrT09oUyO+/VlgnMCUwRwDBfx
tTflHaqIxx8ksI8vqLOZ2B1Yx1wjH84Mta2fH4+4whU04DyUgxsezMcJss+1nrPf
zZ+KdPvp3HFLDbBkOzklkVn/F43YbkQqtl5Sy8t2poPtgRcYX4htkHCrxGDfP5hR
7l3E/gofur2Imbb03p7VUeQ7aCXwxoTyY5eZ3SCfz7/mJ+5ZdMfnnfbTDkDXTfj3
X9+BWyWW+PZCSwvh6/5JePoJaW0ZkR7zIAsCF/tzB0hVLZUHUf5CfEvrLe735iWh
VO1xWDQPTSJ9pzbXkfhulM+bTb6Gh7CicwwDIJSGkK30OqpsDvfBBbXWVdMP+g7n
MNiwOKiaVWWxxOKKgUyZ4kQu4tgte/vAy1Es1peXol/BIzzuZGTLKnlzwt2wvB96
CnbU1DnLMg4tvjqf7XeNGIvO2+tcdVRP5t2GGiCOydgf/McKmlnI180dbbElqPXm
l6QK6eQEIiHoNG2dLWsg9Uwn35eUuRs7dZcMk5wiTGYlMY5urRBdwOjMkTgmTJXr
sSqtOWgHO8nL0zmkgnjYclPclIC22M4sSFpjQ1z32mHvPMQCPcyAxcDbr3V9MEha
yRmrtMY0gR2B0N0pp4ffLK5r+FWQSXQwKiXxucaPedaNDdSbs+3AZzy5cgBbrJ1C
ujDarGzRykkpaw3S5gIKthP1onKEEMRBqhrFRdenr7SoRjD4+Zsz1NeO5SxTPj76
wxl43brIz2Nuu7co9BpkEW2dCszrZTmAAgSowG6U0ieikNPCig5NTVXKLsm08ozu
NKKvWLnObUSGF/wRHJ5AihUyFqoRr44FwvsCH490j4SOCXB+w+EaUBpIUvf0EaqU
gycV9qbIT3qbYcdC9mBe1TsV2EEwhnFWD3/VORWxM6bS0f3jIPYdxg4qFy6DDNFo
llbLDEXMVKBbSk3Q6iXpa50nCz0t7MSWVng52MJJZbICbn2NWizKYpQruFfuul9i
5DESVOVdSMg3h8U2zPVixdU2OksyBQFiFHJbS401sGcu1zK/S0h2irR23pkaQmcT
NQ4ZxUuf9Y1DUiNHbrOhryD+2IGDXg+TTNOTwGwg/7hIXgiQfP8es06QEzpk0gYD
WulDbGLi14fh2r8DxhjeaV/iqZ/MCSfBECuc2fiiJ3EU+AshfQbrNY6LLUJ5RtVw
n4i6l4eex/7piMsOZb5ypzqmEFsdWVpfltskAa8+FDa22OmLxpMM6CtBFEZs5izz
mWfR0tpbQPu4mPTfWf7WpcK7RVY6EzKTZNTbIJiVgbBpCSUdWHkEB3KON/vZS0Xv
GFHaz/WtEJArg0YfyRifY+cBTUX3FfBQW7MaEO+jbQ8sv51ajnI9ukB6jWfOnXhJ
JLbZfqrJlNkmtB9H5xjOhbkwH1YKaz/xVL5cfsUn2TiJyHmnrMoU1OSBeK1OGG5g
8C7xCdpTMTPyfNBJSFU7L8dpwxshk3vv8CWQ7FbQYk1x/l6bTc2xDvvhNNwMxqDw
rYRUTYU+EjFOeO+s7h4nR9NshpYJQlegS0oKA16a1GCLHtgrEy3s2esLtbsa8yEi
g7+oJvDQmBMAFP/9EN3lrJrq2OEO2PCi3nC07SH4JRjKn4pQuhTNLyoKLsgNuTQ+
R67UbzVbnq58Xns7yl9HMxkMpQ4TwGfVBMeKuUtkz/PCMzp0KWRYFQ4L5Nxppuns
rGHErpWlh3Q1VUmtVdx7bUfZGeNK2RojB2ttCJdBcZts9HO0mqSkT7m9DIGlboCZ
pedBRQDNVwBODnGk8x4H7P+Rrj2DEpOpjnoK9tREJicNxTtqYiBX8R0LGEZNuxN+
P0zQ7bOjrDLa+IEdkACtftxvYTk3V7cCeWUs8x+aWw4hhn/mXC+RDhmhTBk2uOgF
28bnAmhYLO8DneD9abbmLel65PL9O46EJSDhGvwMspYTpz91GuRRV5+WP4RNGdgl
Y4wbqcK7R4b2i2ASzroy0xACS+08mQky9tDDbo0+qsw5+Z1h7VQ6ncwzPgPVHopa
POWEJaMEsYgRJZlbCUnGkjnyroWO1mNk2bxWtPOMbzEE42xGxLbasRM7HbdZh6yp
UZXj1FA/qqsWYI9WmT1HngAtMT04syKmHgrnRHMWFdymMaK75hJtd+7ToZnNUJ2q
oXXyRdVySfkyh8vWIu2pzzkGcr9GXf4bhlhJVHw8MHT+XVhSmYO1OY81Y8RWNTbW
+5SeUbrq4azGhKX4qUWm2iJt7fxte8AeEnfnLKH92O3TDHSN1h9Xwte7wYagIVK9
7ypkIzRpVTd1d59gnoq+2bn40igANSmXm2T+Gj6yQIJch85vW9hNkU9/FkzGiWdz
WoAJ9ENvmmdXYYmB8Xpqesm48J+MRqbJhRRb9zLGcrg11QjbQIcCSTNylrCOeuRw
FfxTr3L09A5sS7Ub1lrP7NDG0jSPjWsdQ2Upao1RMgFKQ4WEtkErnSULhCieOyXV
QLwVzRI8oU2zw8kCnWxw+riTVVhF63p1m+QCAUWzDHGW2IGNIC6TutepIBmGYiqC
A+FwnXikWrFWOIacXs0xi/68iO+W5vnapwkrx1jDASxPfs5F1BDZF9DDKd1oNTDo
YBvamuAa9KKkyaYgdw2kguwsLoTCTdC2bPm5eYcQoL5wkH3o4/IYYj5inj25WpmB
RwsYckSuBBb9qswM1e1sHcxaTdsgiH3sjEX+gSYRLMiAEwRaWjh+IrvEO/qM2zzb
OjbayvjpgPreNjlQjXDJ8m2EoRwYoj7eZkKZoAoI1gruMrqycPfD5kOAZ3NTGfwx
U/lFcfDxjC3o6AVn5joNsLI1FW9+wKs9uzhF8leEVr3xyi/V66DoYr8prsfHdr7A
JKbv9LGJni85NDDUkfpnTtMVd3LzkhbQCULCP+hXlwcWea6Ii9gxe6Xy3OurMm2k
N9kqebe9jeQbE7NWnphf+rdsdaHhlpPPMNsKx7iE4yZyVN/7qKpd+mZ87Ef2C4Zp
8k7tcMb7OdNTUxmQlBjOceC19RA3eCW+L7T/rFa0cDqthIV3rd+WpI4r0u3VxLV/
x2z3ZdxuHcDtncxcukXABl5fvMMgg4IMYqWAA9UZYVFLy+qQ/2NKVqH6Ep2EE6o4
Rv3BSka3tWhfeb2YH1LOWOj7xQkz7Xztkr0bwIqp2fG1lJp0+gHv2gg8egrmPysr
Q0FnAsN8zGQ3ceXCipGq0HQsRphSYezhHDVWkzo3DKBvP0Ce3WK0PY3WNDr9g2Vf
izUjjxM7YgD6Pab6l1t5Ak855f1uztPIaiA3SYza63gUlKLmGQt3jJESBXGxW/vq
QnEt8k8YgM0abNFz4RkvUAtWdqBXD+aTeN9Hn8YUl5ahs+iQiy7G0BM/KXaGs1zQ
Ynz85IvhlwwJgLpuE+Ih2m+/Q04dcPBaQ55CClExIntCNQx4gbyH445M7w4OlRiW
vJE3+0p+lRZljcHo4AMH62H8yvn9PiVecn34a9L/W5MioGO8C3y99+irN+dYDYoI
SBwvnFpi5mKhmUDxvLGCr0GLxTUhmLF/BaxbYinKEHEoFZjRq9RrY6vc1L/U5ZRc
iPsou6VoXV5inysBVaz6/S2HG3TE2xuCICrEbuCfkGGBtl4b9e0lgvZv6EywA604
WgSN3PSLgSwFU+xyOtYjySNH9uCqMNQ0xI//7VkOwKBMiWixKrXycmRHiTXjJ9ne
s1JqK3YVfAJKutXqjIPP4JFhCZuBgmDaCKXKvOGDDoZxcB0OJp0gDF9BnbdRDGn5
5l2Wp7fGNplhDzKHpCj/hZNKksQa8xMzA4Pe90O3wKyYVYMcUuaGB5sPaDtXadtk
cUp5mJff/82vymx/R0y8qokGOJ3KXP+2sfcidCFodriVZ0k1v7xnKY56HjkX7m6F
X2D+dPvV+jlK3WGKcRTIsiC76K4TD9HLNOn3kvCHyGSfgYbkGepOxrVGHZ5Sm3wr
br1f4YublqtnFHSue2QxN0bg3TH/4ggUEKqgiAqeWu0a3DK0wpHBNqwbxDZ9HdhB
TBpyFndcxT1eGeLmjlLgoxx85W+80CFluebbsUC9vJ4Zr9ZA4Oo/uyJp0Zq0gjgQ
ycX96STa9DYq1oB3Leoh0zsf2jaAOfh9xYgXfrq42LKo03EqXWnwb/WvXaPbu1+/
FIcxFKcPFEQaB6xp3WmxK75ZAjpQl1+ooxH8FDrnDdeGFuoVWEl5Nb2MEI2tBiSx
exBxxcvmdOEWQUdrANWNsiiJC/UM9tr38FmqnDM9Nts0+YbrPiTO8x+FMzVhhcIH
OikTKnVZ5AA+Gw34LZIpdWUq0LdePf8LnVQl4fRrAROVlRs2QADeDlV6b2+NcF5V
7FSQlnwBvEyxT4ZqUO8beCWQ0os6tz36h1Ue8CN7WFGccfHcvRh1hh7HefF4AssX
A3iyZgfwHH14x2prttGH3Da2xzMaL6kLxTFPp6oq+/vHzA0v1J2l4u2A3ZRK87iv
ljH/0/mSppTcXJubFDAddiGQ+tEhzpmp9y9y7lexD1zh1nQU8sHDiTtH1UOuT7PD
ylbiHbXru28tMmSOZ2Qhlqh6Y7T4b7nGG3WoI2OxyfpLSsPUrgHEYUyoilKFQgQI
VpK+nEczUAfU1+sawD1D6LOVzzRn6gsmR8il+jTn4RAvi0c6JMWY/pGKNkE1Lsde
W4whGwsAiba1MOxNQ9f68Hy6lp3yC5ttdFBqMsa/Gat8n1d8bGwxtdj2X3kanv+H
lhGPK07jKBoVLcLscZygrl8hwE3P1Q9IijZeOZUUHnLAoty2I29DESju0kozoqfH
T9udQCJ7yuQaxL9fga08V5b70lOz0+WJjQrHt4d6QbviYYUBlvjrP3S1Xgk1RnR1
6grzqML95F5xxBq/++EfDdCA38IgFl8T1QPvDdZU/omLMFeztzkshjfM6oUP0YcW
JkD0eH/J4wrEfqamHATOZPTa3ga6wXT4sCFe7N4M3/Sv3XrQ8weo1vdBTmtnXWbT
uKiDpnhGVz1jkKdkoSmashSa4tsmm1BSJHGAywJOTMC/4sPPB92Z+6nTRQl1VO2P
vcSaxcfr43rXfYhy/4itX0ivYGSNLBRNaaVBQuAOx/2N7q2VJ2lc6plmtQjnPk70
i0s+HLh8W3yLf9EsIcEJgTp1cgPjhts8tAA9li5pmuHWvwwi7sSLHafHJv+SWwNl
GnrK05oWVwlTV3WWrlzqdmdZmOQ7YFTyCnX6MKqkd9zppCz6w8Rt2oRJ7LfUmATN
7ORjPo6PfTLTBIRojj968MAB7P+CsBNtIe0nDAvtgDMtQlJioqgrwg/DWTVBE5xT
br46L/tNXNBnWhJce+Z6SazzU2yFLWRMhIFQKfgNGZwze/2Bfaq+pZfDmVfOu0/H
WWZDDi1urqOQYmc2IKh14oSAxuGYCn9XJcb6Zx3LIgLc9P2ZEowKeNCKOXVwRqz6
xja3TbTBBW8eqqK4kIONEkYfbpt4x2WL+t0bOtYakl8GAMEaue44F1kOD1gyGWua
+nOLEo0tRSqgzY3V9ruL745UL7NGy6eFfNYZ+IJO55+lWRgZ5xcdbJ7d7BQKSuMv
gnuQS/kEZYNmjmIqNDkfjIjUC6aR0afIKBVtF2i7Tl0LM01rFh1iB3hNlff3UdRR
fuQ7eMVIKKyYQIcBoDNUwfnxynZbxh04zEb4QJQAJGMLdHw+pVYIkdGWHE4fxBFw
/K+Hz77RQ/n6COsmgicER1EfsQEPnWr5KKj3OglzGyjQwrye0HCt0ukGAhT1prVu
94jEjvJLcVHGuLtdNov6Dow4/xdV+sRV+nPMrdCrFOWuSp16qD9Hk53+doMFHPSd
/72zqBdsFHv9rSdDCEuXL3U6skLz9PbLngPMmISPylG8cKkqUz5fKtC3dIJViQuj
FxT6fqQsYOG/pxT7tgnlOoFbvGh/QberjHb3PXir3EdH2kqUbwunnwq5v161tsaE
nJ1ViGI5TuRPJjwN++dKwFz3i6x/NtQap3QPGwGYsdggzq1WFrr+h6tLxn7AvaPd
lBr/99UNi5i41HcM4Yg2P0eUWaXWQlRJtvzbEhoWZk53yXRTCln94mJZxJf74ZCu
IFP6SI11bzXVzJb5YPzFegqSIuspYmrigJrchfiXUJd3oEw6fyUYXGLv/Q383FlY
/aMxIURO9McKORfSxDFPEc/R9Nsa12JYGhSzKNM/PQoapoVxhEofvyxd1nRxl7dR
ihiR41hlGqVx+uOnVplmGah8N6dawK12cx9D2vIEo0HYxLI8gHZKS1AJ7WwxkBrZ
5/GMP8DG1U9/PoJh0eQhTziwLsItuc4oX5l8NHaKUmG/zS1nP+8v1TvgwoawaNxp
UPrKfjIJ1xxddaAplATkMJowC0Sngu3Vy1jWK4HPFf8oODdu6vL2L6PGCdiJwJTV
oFmt2v1IFSstadqPA8dk3F3ucQXTvrxzGPZ1IeEkpnwtUttkdcAw3LxYyylt6r0z
oWlMk9nE+GVY5lFrRMoDuA69DJgddXOt99Kjr34AC2Ip7rValQCh2MDom5Cdh34q
qwR/+AfJl1VlAlOq2bUSkWQIrjqYquQg74YuBH3n+skT3dqqTs6tZQNtLrOZTh7M
n33YKJPFghm45bISpt1kl33jWqaCwfyHnJ1vYiIRW9liOjZsm3+3Cs2cOBP6upIE
hOcVzWwpsq/qhsBjpXu8Y/jKVP+wnR9JnKLb7wAwVC0TcvuFpkXxa6oPRV0GOILt
LrySFTnO7awg2HzKqerGP1UfSZDrouBz4sUKeq//Ka40xE3c6mfS9Vf8Xye8WV5T
LW4zAvaqkOleYeIVEck5Snv366tG2qWIR1TPvmgrO4eQzZsYz9xExGEFTIK1jp3l
FzPDgkZuQpRPvgkdO8wkhwKzgfwSBjEzDcmgEgbkz55WDrgDqFEHbqIxAflCj6k4
Xa8XxExaspfNCaSX7C4YzNp5VeASUmDL+dpG62rmFYSE1494Y0qNxCW/uQWUVbcn
c6VUZ6YpMqjLX0aL8GP+VvHOxswQdbnHFiWEZ1k0i+TUDMOUNI0rGZzmLwrgsX5d
dsb4DJjbjwmUml1eNTDnZxflifNKnWDovf4BjwWTA8Y6IlVrIscNGTLzyO34KGll
QH9jc7bBjle28YEqxFiALCqtBivMPfiY1NFIVdrtxb7O1tHZXIqxqL85MKXSMN91
nhnaEL1y4f7CfW0VWpQGUTFd1fuqheFy5q7CVPxdyoqCmRD0VDb9DhS3O0boKvVC
T3ZKKy+xMGTcVrJoedr++B92+OeYjS/TcMr9FOklL6P0eNn7FEr8I6tKeqMQb+XG
iZievrW6ekHE7Sno4ITKCal2B6VHEVkgMaOFQkY5DIyE1Z4NiN9dJ8cTJq3nBmJm
lc4qJ32JYWzcC3HrkF2D1Vl89PjmZYbuGuE3cfriPaiDpWQ4ijkfqrdLYEgnwINF
BprXOeDFvBr0a68AEU+Q4S8+gdqHyWzrzHJH2qATL19ffjrkZlWgmELDMdcv8yro
1xHExe7V2epe7UnWjomWbEuu72xz9rcSqFk3RRBAtQklvG4oo741E6Tk7blJRilH
JfKW8QyvFGmGttjNMPsScDJjMW6abwk6gdCz1xG0YP8padN00ToMGCgirGdODyX7
gHJRhyzYesxKkqXONKt4GMLMvozFq/cR98/pw+5yiJVr+9pQjWMYJWjuLx41Tafg
9zJEJe4JxyAwjo+ogIZCSJm9tN81kYEMF15QXspN2oPDddXFGCtwRcb10BRIqluK
Xu4/o/hzJiw5orD/GH5eNEC7Hn9H5Aqk9NZ7SIB2bdhlrDn7cwF8Bd2TvhaqRRve
NV0RPurMWy4Z+UJOkWbOsanPCzwlcooZkFrYF48uLHytWURuNZ1D28BikI9VGWbN
eJ378krFaxOKzBVCOPOQiRb3zmEQzdyHREZw0kk27iz90ZVDUZ2yFM8f2/2Y+xpe
R9r4CIaAUouWJ1ZO6k6HKBQJQKWZ4TB6fzJYYezqcy138h0AJZCQFtaLJFeIdnAI
qtaAAFggPnfIW/vLdGKQ/SeF8i7Y7T23ldEM27MHXXUY1hwQ1b7X0d9omWxm2hEh
TuykZZAHGo4MB5qyVNOyKsretYLtCxpoMq0Mh2mxocRXSa61Kg9WyOdFkwcXb2xT
n2Gl0HncKtiVLZtXsK8BpIa3mpvFLLtLB5YyZkSQVNYyZrYYtlwtGfNEOodA8HgN
jyTJUCcD4aUmlCwgMzrHBxgiXdSBcSLklfzM1kA2POA+HqdFhuX1W79radB2gvqJ
OLGq0SfsEJ4ydz5Fd4MrpemgeANPlOsH/KVquPBn4pkhnApwsxu1IfJakljM34G7
T3/1bocHahZllL982oSV8xu4Vodi+YGoX9DanfLnBCy/GXDWh6TKo8JdKn7Hpdcg
0HoLSTcr/mtCjfQwZnDAWUJdrl6/e1v63SFHgU3PzFt0Sw1Tpn3cgpqLSyep0HDV
WdGSdoEgrzJcX1WpkJHT5urZR33MdP8AfOoG+jt1YOjtDQn8yjoP8jOe4q4EmWRp
SLuDx1ETKcLfo0zHGkUJAr1ixEQPSiidti2QKLxXhf9SFLQIcQOIHFhp/wBqlhLu
VdGmWNh6RFuIv+eAWOPkRFwpF8zXDwBIb/rRZpGWY1uPDu7ZPAAmjWanRWIDRwHt
W3urN+cyHVTB1goEXKqVOPBNWF1nMdJ0w4nx3Xgq/NLevkiwzHbkUWyW8i4Y6bdH
3lvFcEZBmAL8WXg9cModoVmA6I0X7JZuxB9FcH4ZsbResEw8JsdCNYsTwmQtnF9P
U63Ip/HzUsm4rqEaEh9V0e7eJk00pbsaSoTBPDrIrK/ehZIMXfL/gxVlJkTdeaGR
B5vh5gXlPHsCLD6TMFx4cwyZ5UT0nSc/c3XDDckoQAbXKxk+CdiGfILzYmWwg9UQ
TPZwrUcGcnVeD9g4IgAV0VuSKyPkIwIyQmQkKVfF50FnHNsjZnt2T8UDAd/TsWBN
MWIXwDBvmTyV9YEkFBI59qpl3WbncwUUdTyyHuf0Tc+TcgE0TyVhCeLTGPqniwjV
OAI4giKo3RUAre8HkOSHF/G5cZKdB5i+Ll6wh2h4mjvRICcT4T/kdmg4r0yvtlss
YS2RUITDEJVTzh9ewYezPFUf6higsfGkV7adCHXwFzZ5s5QRsMQtz47RTD59WGQq
2SticioBBA12G8nmYO9yhWX/mXwPlvtno2lq3ECSccKMr/A9dYtP2d12Y3PgFDHl
sF9EY5KUwNdJ4ca5Lz02Eo9OSvdXlhiKNUtpI+CwblBQC+ZvVRU3jpYmpzDjmDSW
CQc5x2qwT/xsqxQKNJBdXz1CPiIkcxE4DDSTbS8bWMyX02keUygEXuHF2nnwBtCq
rKtK9YvXsHifePOoKYdbyzGKm47qRakSXjXNfA/CEfwuSND9PCY5petGEzfJFIsp
Jf5TJ9ntTSMpKZQLj/rqysI3VJMbs1j42T8+hudh+yUTAES0uwyHD/BHz4ZkGWqT
D+S90Sc1LpDYrIK997qSKOAxhkOraVWCgTEY/YvCRCYtwTdmRi7CNIV68ZykmMF0
UUCOwA4MdCVugoL2/1lBzFV/Uo2U0olgJqRxrT/r4M4m2LuIptmWuF//ZjnVUBsH
ff3cLHRMoY15NZFwbnCdq/VsYYQipY3A5pvvZ/OPhGxmMdMroRfdSiPNGt5KOqAp
7LKv42AT9fMGXFc7Su1jJrHV9QS63sQc8TPTKuYfdr/qrGWQCvWKtgH/M2yArTcU
BinLGNcnYynyS7D6jxihCpA5CQoV0ol2th3GNAY0YMjr4K5X9NrS5Ktk/vxT0LEv
jkRuq6HTbREBsHBlP8XPGGLV3s+TsFAJJJIKrwAddxTnsNZr6xH3KYFXMlJRxy4U
fyc8FtOcA21TKNEvsIr8Tm0bjiaHGON9957p224+dhXp0vYdZIybDfrPycOECWts
Jr7j5FbGrJO3LLnV0uOOGvVVRrmpFe6nyXhWRRyyankfHAipyBpmY8ERvnyWClt+
cBOCZ4TpPMjyi5slvgWHFZnyY+V6wcSAJqqI58Nnnb++AkMxBl2DFuK6q5D+HCQn
HhtsvRc8cCzundMpm5IipSulVOzdPfeIRBylgy0c/DluquLF+YKtKtifrkH7ySIX
QqyAJRkwqwg0XSUJwC0u82OXFcxjngorg4On4q5FqbVIiXNUzlKnTw4TmuDotlkL
A5+S9kmzW4C5/41QodbZAKZahdOye43nBD9otJnYWLpWxVOYNTYSBKv/YbEtExaj
NW9FQ9J+KfLBbKSk55QkmRIHbwYquUJIFra5EomSi9DF0DkNb9Z3DYIANvCDoY+v
WIIdTnqeh8KpSoZ+dQekJyXfBrOAcQs8enxQH0IPdF7EylidpU7dUcHcZ9LcAKrq
c5/n23x8t6oQRcKFgPwqCRiOIo8ahhHWtkil9bmylB6HU3hvlBRfkaaj6UO/XqtW
eNoSiu+dV1xoD1MY3uefxn5fJGejqlH6QQo9Th7mWOTqrSrZakUIqL43YlTrLNRa
97avICxFZB1u1ts7oXcYKCcuovp+yDFiNCceZ69QaPwCnZV/GuCbtwKnMoBeGN+W
DAfO57nq/MYGPUP+tKX4tcCk4Cx4vVZOkCkJR49ZNvbwgyCxyxyNmtmXWZ+LLYfG
tuxEftMqvh8dTG8blDnBDwkRJyFsHLTfPF5xIMnITKffg7tsNyhEq0NwsM8M4CFK
7GGLirXTy7iAceA/r6nV6V2psxMgt3dFFY3W/zS3XAveFrmPPVljl6FV1qmY8qk1
JDO6rjK2wM/85FYxNPIDFcxZ0F+LoiVBmEa5xrxLcOKl6/+i/JHs29VOlWR/72dp
pFV0Sg3DQiOuBZ/nIbcGL7siiOnnUe3yr92dALaeZs5Hs7OHWrakKkaSXkbJoxSl
7Bp74wNw8WjN42BD6e8tr6lGw96bQA7D2Yl9IODqDtRyJvbi1y8pUXPt1m+y9Vyh
xndqAGis6QTQ3eaUy3ziaKOVufixnxf8529F2VlMWvUDzGURPWMoCfcLjRfQLIYh
eiUX8cgnYunus+cPwkRcrpxiI18N//iYo+qfWixGgf4H0QHrEUzq3jRNqPZpUTuE
6yqJPBQaAUJQ+/lsEs6v34Uz7q7kRlyJ/+iwJcfAoDwV3QX8DfR1yknz0C9cTFmq
nfNFsihhRl39oOyCH+wNJ3ejhkFRx5gPWCSugMGeb8li5nndZ8EwG8Na5ynizeuJ
kmoDSserPAzdPni5l63hY+PS/8XhfmXRa1iWE1JsrOsAcHBUVHNqlBP3QG8JaXiQ
aPS+i/yQR4yI6z01455horshJKqoCniDaE55jhd7ar1i0k2wx5RfFYQH/XNzVGoU
SeUeEzWnb8ZPYT97YgJagbEGHZS+t282ZGhpEbpA/FwiRAP0QdsgrnschqzHo5Vn
itvqlR8uB2cWYVvUhMK2XiW0duOrdFI/bpTsmhDc2D4G0WjdYGLw2wIfHTuQMW1y
ZEiKJGpfkGXAMItB5nOR2/RMtSF+m7jelKU3sW9j6j+sehtGgUDZO8bSkDZ0bh+G
xXBBGGS0XKp0eGHBcL54yuyilB+P+w250R7eWoZhpIVNa0abCw2s4cW9Xafk4lOr
1btyxyGesW5Ztasb2xyrFwBKi9OhkqDnGRp4GW4nAsPFDWRMmlhRG5swjEXfSCw1
PzcCT40cT9nBoB8nCHRoASc3ZCB+i6dxuczqUvdoz3Z9Qwgeev2wC8EGDV1OyBCo
7oXyJer+/wlIqCP9E40Xoi1n+OcX8koncDFIV1viK25encqGzDpLSZWZUKRIv4FD
Y1drDvEYVvNhCPHhEvxH4Y1JESMhxa9qzUu/xZ5THdid4066uW62r/hC9xV232SI
FBi0rk0XiJq88kMLFLrSyaJGVQ6sfT3RbNkg3lD8brK5/7htYQIr2p5/Xjk7XwgP
o1k5oot+ThnuNrfR/ykv2lg52Pl53iJ74TJkZaPNs7ZX3jDfwkgtryJ/ZnRTcCwn
jM1dCc3th0zToGBfmcP1y9DZYcQlX5h9Wwr4BPoU4Iy1NKzxcxZGFs/jxGvIxhbq
B5/yQH70pbOCixImHvEVWhb7d3e0YB7o4UcrhfJJpkmOJqklowJd7O1jFKspLfyA
a/o2nr/xQ5X1JsdeNwOY3UEKTvpQ2y8yv/BFw5BNiXskNwB+1DQRMSFwA67MF6EI
WS5gyPCtIMs7mwvVIjFPW1n3tCW8qrEIq4SZkrma0vub7HUSOegujHer1pu+ypob
Tuclrv5cGpL95QE/sl36bpDq+h2MJBbDm7UtH2xm5yUTcJtJ9ECqBmPt3yxCgR2j
ojUjuJqQsT9G8iRLKc1pj8sro2JgPOSy8WyweCN+eHdgRqdwLgwubYIlNAO4H34T
gT9/wmFYiYlfyIcXa/hfia38y0BXmjPmSC37uvNpFbWVLgSmfELv9+Sbw4b3OabY
hiPapU1yisox8o9NIVpLPcFVFaUcHi6VvXJOYLNJ/ssH2yBMnp2QZPYpB20Tqqji
cgp0Kuw2afHcpeVbwyLhEjstrQ3pHeQ6+kTg6yvcK6Q57+0vN5PBDk+fBh8BCBHL
jG93sH7FRT+nejVwLgRkzHStRlz+79ZfbF0NqJpEntLAj5usu1AneaZoialWB8yw
g7yWPpjh5OV2FVPbj66t2uOavD1BR5ljXZWMU/UsgFRdRt+uH3AjS7SInMQzywPI
GObK9tWt/K5EbzIcmLeA3HyGNARNko42IqLT9eFor4lJJ65a31n+Mhy3aXE5p2FG
3nOmtaFM7c+pNr1mtK8JHudWBn6sPfD3Dd60l0L81/xXK48m/aq6c+Ao+Xaq2Ia3
AfVcfmyf9/rL2dKSI633QTA/y0UKuv2y5h0ixiVOqBFnWwjAW/tK/CKIAwX98PQt
kF8swGl2Uh9pqnNS7+OlEHD9MCbJhU/B8Z/6u7cheBRKywcW3pTgLP1P0h9ohMdD
kgyZQjFFPVgO0djwtWEgQ6lFafrXNL0wi7/dsKMC52YSDhxfbI8eUUSdklnv/6qg
5gfpu78tr4T/Pbhs3xq7WAUkLwLGt8uQyUTYY629qFCrNhRPhqznzR2kuTZmPelU
7+jUiYleUHKe6HjRPYPQo85QzWJn6Xl8qX/o7xqq1VyppqQeZcmE35vsXTSDOsM5
MxjVrVr0xbNfN1CdlgxoaLHh2cmt/veWlLFHB8W3fqt1EujQPX3b0WPSFjfJDtAA
///FuxsOZg3q3wABWlJ9MF3NWPpbVcSVcuMJRWepcqAsm6pjPC3s4Yjef5hxxerk
C0xUs3wOQLi/tuIiFup4+1fRveY6mPyZbXn4bVO1aBas/ui1J1iGNGDkrIfZiXjH
A4CfmYZevL+AnB7w84QPMKBJL1iyKZcqqX+rDPSVjTOAtHGpWq73+bQiVRlv/lc0
WEPvszsAmbofW+Cbxa/uq8j1kkhbn6O58S+F4hWcCEpCe7f6vIE58sYAfm6MHoV4
1/Z/diY76L3OwNpgqruDcjQVu1NcKvmwIDU7Pt/OgMaMbEX8yYHaUXNntXO1dMJn
M1VQhYSRzU4lR1UDdul0VrkGDo5lu7A71FGDSC7Mdd8sfNAoHgOhE2LHIafeKBfE
xffzxGJhCSp/qeAtImHj2N8vKoh1AsvWWLlETsQug+M2IqXHPWS3lA2oLJBE2gsc
ygD01ifkLwiOOLKZb2xbkfdN5mE32H1csJ4Lkfsn61y//IHmMKmqj6RCMk46JRPC
f0MYcwRrqcLYZQ/TokeThM1+EMbmSJTty/qHggvNd7IeVQjIhTlNfzM4jnfSLNPd
LN5RxZPmQr1poxsfKT6RAlzKj9pz1kXWwFdPNChVTucl6PA0GJlebKVmxpAwS8My
0tOSkV3OOi6EgbZ4Ici4rETEa+WGcH2YuTrhU/IfKkvQMlj8whVO+dwWi2tR2z2O
buKRyJmUogHbjApKZJ481NFR+r557Cajdc0ON9NRq0pUV4/hwrD9wozZm70aPABO
XrCudY65SH9tn2CtkJ0IkzRL1a7L5Pz6ORGHPURtTRk5O3KCSYyfbafU1sZNeMMh
S9q4ueTYpdGLJBLrP0tQQbp49MrgHVb9khTR28/6NhQKD0zestejuztbJsfRtCsn
tgdXFy4fa7TxTcFMvGg/6y4cgEi5jNm10IJ9viL6o/qWZt87ksR6bGPcjcPYFElc
j35haJ3PQr0iwWfiLFod+PCn+GywWO95zxKLFyH5kJzY/tFw43LcHH8cTXkRThZB
oh4ubvsedC6u5U0B8SqYFMdzy9sYBxFP27hI7Z4lhlbKcaiOXrpmJUw+KxzB1xql
P7mewcKBWTLWoOSWguc/PKiK+LEbAnnTS+xqXcjPouqvvrQ6cSxylcbtfpmA55A9
AJ1Ey13OI/ApycQJZEXdIu1ar9AWG3R91HpGtYeLhFxnYQHrkJ/7ytYG5qLfjt0c
AS1lGIP2IZ8CItGi4bdCePkP9I8EYwM2kd2eBMiieL2HlxJE3nYkZ7tvAf7OndIR
1jTX5fchHaOCc/cyEZlvIlHOrGa5v1N9utTh+kZFMO7RyzmelSiNNqO9EV/qa90V
6fcUZECyG8bq4rpcDDjf/lQiUgoE8SbxvJS1922WCf1xP2NjLqA/6L3n7nF8WTp2
FVilDNPBfaz0R72ggzXrpKDzIKab5wzOKph0G39ByCzwVndbi9zZV+92nMqVQ0GL
30FHE2+C13vFwftBnjtaOdpIbvfosZZnhWA0ID5f5n1khrK8PB4qgIzG4E5qh+5W
NI7Pj+WDEBgTAwQ2MlCkWpK1tkM5Nm9vIrRqMt83yjo+45gL4vBIDn07bf5Is049
tTaXPEDVPSlVVOBMhWxRuLmNr2G0Qg75sOCcFYNQ/Xo8wO4+QCKfwai2HZaT6W++
2hsnOi4HlcfCYheJNVdxCWOOlSv3T+/yhdTzx3LJSNklgTFxIXJ2ODi52gVS8sWU
MMGqhMjWvjEKCF7OkJp7gL3iI2TcxqmXLqWFzmTbXfmJNkIb/xLogtK3iu+VytWs
sWWW5tiVOGyEj6x6U9k4Pwgt6z9B6YSQYn5FZhIvYXkl2/795wS41ZHsz+NUPYu4
KJGTJsHGj77eTX/+EP8K/7c7MeP8Xba/EnzqGvVwwa03skSZhSS+D1AgFFaSuKYd
0XlQn5tALMsi/Z7ekcIWO9xNydDS/ERzSmyFGJzz8VFSZYnhYuclek6ZlUOyjLiP
0gjv+4Tfs3r8SbOsaFiH+nfYvY/MwHUkmxrb08negcdrvMx4W+1Xo8Zx0ObqxMNE
b53BTqb/0eSwZ2p/xTonJA3SusJcSNs5djbyBQAvdt0XsSmEsb/c7G9BH46plLYl
2F9VRqLhjbFNcCuECVj4EKh8iyYWd3aaRzqyN+J0cGHAL6jjGARKhyRFy778fzTC
vmNBVfPmg37Bgw+BxSwd9q5oXjXelDElGNlnpQf90RU9Z5HU/XQlwsXmliwK6eG5
VS7RAFz45BAcjN41cnbxsbxA7P9qPI0Y59W5JofRbk6Kwx5neMi6wTos+y2CT2uA
l3tH1G3WY0u+p7+J56QowI80YjvPnc8WBY6gTy6Pk+1icoAPjiTkvoXtZesx9aFI
H/DkhKEMeN/c+XjhgAFnMQDasDAhfy35tpdXgpNk1Fs=
`protect END_PROTECTED
