`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HuD45w7ykkG/ylvI1b3tcZDbLyua4j0I0QjNoUEKkk5ZCN6qXkzI+XDN0sFdkNo/
XQ85tvH/+/MSbEfKbI27HRLfqe7mHqTwPxUmik7hIJo7sU0/mel1ylhbmsBw+oeI
4DaZ21w0yjX5BM2b4qDh4E4jnDNuWRjVASd+3Xs1/2LtRWXEFoEJpS823el5Zi4v
hELRiIeA1O99oCv9idPiGJEVTijyQFt1QU0OToi+8+St7wyu5xBBIsnEPjMK9xfC
F+jMvRxoc/psTmq2keHm1c/InI3ge7UrM3HeQQr8JUZrm/OIAIyz5pxGHNUMpFMS
MYlZ3AV9FB7NrEm+evTtIyGI6/3w+yhMtvKChDZ0PqFdMIJt1Vb2J0p97LFkBhgx
8d/43E57vv6xQTxc4C+1qyKa6yiwbQ25smEY9MkawEHutKfMzwbWAAOrSuUtd+VB
8WeQWdcKPAnQM8ss7FLhMS0CFdyBnWBKzIvqDnjYDtPm+EKv4ENKXQuqUbs8vo/W
xgtz6wg9LS82IXwC8GKpyy3ybchO4SxxHcFF2GBXiaAjkjvKxfxN1DSjvjJl2WaW
NqpzRaS3y9qb1JwSBzz8yEBFX1dbNrWxvyZ1tmhiHUuGDAF6Fmwzwxsd/9wSgygw
xt3LuEICtrQ4V9ysxEp4MFnQLbGeFr+LNDtkdfc1OWiD8uejrgmeF/V4CYaQ2qhG
RTDJJr4SpmhYJSe0gFcZ0wmgSl8Dakwp8tti7GYMrt7kOPAsMdmnWoSXx/2VBCyD
G4LJcZ5Luuol8Y2uel0jpRmGC+fMmxw2w1DcLqKs2ve6rBUGO0mk4tYHWpRumwR3
B0KEV/PEs+m01z94+w0wNXTy/j3v+ReaoGz/MIa+PpQXG5sorQwdg9soy0xpQSPm
OjanPG25vO1+vyIB2LMYIkwgaAxt8RPhXCREFWjGzTSVSVuzctzLXvXLrjndEoHf
OfUpzI5gHl9WJAE0kvnAUzmdqHuyd7/zawWpN2L4vcwBPe0UmCnLl4ABO6Z3x31A
TSBELftNZI/0TepYWr+NJDgZUXR7x/jjMOBAjhxOq5MD2cPcOViLvQy/iiGUu5L6
jcot3fgtgoSDBOA8ozlcxIgirkX9KeOhC7r4+LsMmz+YejxOdZJl+cysPnQ9XL8S
Z2G/aK1I3kxhptgTBWONdp/talPyPkvRzwAf9B0+aXS4bzzlKWoRzvFG8+QmdxyP
7LxfpmZ2695dCa+qGQe653isHLKaLTm2ecf0GDHE0zAIdKIsqDlxZCbqz5J8JgW2
Mh0OFfz10Qyt0Nl1BY3hgvqHUug2lde9pIKgupgtrzjjZSTfdPD/VR2jZ99blS0i
xKKUaztxpCaHzbaGYqOxHSEdcvvw/h9eszkLWSSSzzDE6qD/oXGfVxB3+iokEY14
5RSo4LQCuf6+cBhh7QM0H5KoC4oaXi7TwdXyMC5Sb6ydCywJfjrk5Pi0waHAaUa8
7E+ukiTrEeYvsudr24V1GFMmHM+nT+P5mx4pKELixuvpYSDLdZwblygAHwnxhy5l
6Q8ragYg6MxeSNKaY+GQ0mh0k4m++Aq9O05UqtIE/3mEiS9mEHHjPN9lazMEiS3f
s6TCJ/ePXkTO0uzZXcd8MCvvHmE0ffU9ghRU/Vu/du3KPb2ZdBejvPEVmHFfkGeF
ZBk+lJBKgqrTFS2qjDfe04Ght6lm38aO2/GX+Tt6CT+y1Jo8cA6qK/1Mr5eM9GFW
7XKNAPpvNWVw14pwHU7jrbLFsHnU6zLjIXUiJuXtijgcmlv+tAwm+f99Ng/wiANg
IdntB51fSbE0wO8uby5AX1FRsfoXXFsrJylBgw53A37lH2MTNScukrKWr0t0bpI1
nHd7OLhPN83sx6WfGAFaOseL9isw8I0ZlElUaG8dZnEiHiotESpWM9C4kJ3Jt2U+
+0U5BZyk7HXRR9mD8yBszIwH7DvBUoanZmik3ZboBxw8kaxWlrAdqwaLq5f9Mkjt
4pTINnSww5iUexvkjIJ+9L3jRirwBHFyTJWJ/TTgSQvWxr+SHjH3cyaEZrFPGt8L
1F4B+IHRp8V7Et+aunxHLyaNyBRYCZZo0wUJHjiY1zrNHdR0tv4rjVf5lgxUvC8N
r7Vaku1rtPujhEKkT6ms2sg1Aoo7aWxSdfyy9bFrZC4bveeSt2pB8czHWGk0+DOM
YgXahxgT1h+NY+49fcihfecgqRT83iBT0ALZZcfJlBRIjwWmUTaDBK3MCccbfIlG
4RauSbLR3GhCp1Qze6UmUsBkY+sHd9xf/UVDX8CQExwdGlEnKazUAB9OR/pd+NVS
Cjxikyy+vySWPhExU9zliHoLdi+mrhwad2iWQAFQtzrjRveAYmjRN+2Oqy3wFSPP
HcU6qmvsAZwuwOCFpaLLVnK+7Emo7sg5ToLAUF9LdW7OzaUdsTN1BgT+BtFM+bM9
HnUeTDg149wTzxKe8IzxfefZlUP4tdZoO1vFDkUTIQ5vhtVhWDUJk+en9EfXx6tD
eeJnS/2VVA/n/JkNt2i016n2Zdb+IvNfPz2MNmhKEFNh7Ej09aizYQ53EJjDf7aD
I1daOJd9uKLHQOnPdBpphvsY1lMWl7CCKtYxWyKJYkowEMca6VoK4UuH9RL/R75J
+iQnQF2M2n177uSI3AvRWuAWD+paAdu/0p0h24y6HNHNMH84r4yXRsMqzCO+Yng0
eXDwcNB7M+qw1VClFFjepvQCO6iX+xcIrTawhiYn8k1eUMyDSDqmoxgBJNEQZuB9
V6wuIGagHNMyW4Kh87GRIuJ4PzqNI9tQkxtkINhLFTw5ARXuj3T/K/mJoTRFd2uw
oEAygLYnJFzYh5M7JPJHTQjV3ZJySqluUm/ngYy50CIV+hYKfHdFGd4b1K3kdtCI
baxEMlZgv2R4d4F+AxD+Dl8wz33LHplCMr243DYWlnKo0Axp6vMYgYydYOL+qIJv
lyPR1ZdRvYeKIBx3sBJvskucKqxj+it50Rx+3ZRkYKWXal30xaUumO6Kycjsi185
iRZUrw7g4iS6TDH3HllvB8qLM9ojQscR/zYX5/MU4X+RkB9I3x47uPtypVvCRpcb
/WvqTpMpSZsYOb4yRfXzcYnqVxEQcnIbv5y8jCtT7l8ErxPSCB/KF/Zez+oksdAx
Ot+3TqcPcWnqzoQAq9/VBFXE2IHAsT0Z/lKY0SNnW+UqulQO7W03N0bmEZvr0MSU
mynNCGxjDMqwcWamaVtzz/ZDJHmnfTTcBszOWPM7jts8y6jtzjDb88rjzupLej8K
e6Op9T8MftjEUUyFZZdNkXj3BMN9ILxPfgBUYvuyuwppgsxGymbLpZqWiIllhDXF
c4jZdjyEMxRVea8cJd1FTW0Br1poMD5oiZggcmPaLpf6XedmFpU4eZyrWn2dlhTc
FE8Vttk+yhVZmra3VSQyDweKtssizTEdfFrqle+yETDMV3FZEaJ1ib52CxEq3pKO
jleITWFgNaiUKt8ZWGQswU+UuiHrDhK+62WdiMte+5n9+vzwbXNkKKUQFAL04R9t
Qe0RlmVT7Tkzb72qGxt6+rHJQ5cjFWICNFjvb5qlR/zKRQIZ5kVUjvth0Y7dhsWm
62Iqysj1zgjtPKKG/FYIgMipjFkjEx019lYNBVIlFEAz8yZDU4DnyfuwhCqEjsZj
vQduICowWM7ymKBGWFgi245eNQ1+1OgijqxLHr5d8In33AhqaMQFzA6ncWJo8WI4
TrW0eO9Rd8O8OXJBQYamkj/le4lKGTalz33uGQ2yF1l8smQBpDyOBcCOtuR5rkEu
YwIVfyW7dfos+jwh2BO/8xyYFma3yDWG9v6nbFK2J8lF2ZGQDN+W2/DF3Io5g6rt
vh0VyR5nViJjnnGXaX1gKVRVCNKaTp5jhX79lPih0vfVHaYUHLvUUMIVScRIzXEy
a5at/ah/BS9ebdlScE9B9Wv8rle6X3HfmmPnFqNdtQ1rNjok0K18b7Lw0yI50rDV
Sx5Tq+t6TX7QAL7JgPjTM9VH0Eox/KRXcFyCusIsD6VZBBFIiEuPLF5Oxu2bZYDB
a7C2BDKbnt3+uurUDiHFblJiqouX50X+DQiySa/xKE6w/9kY4iaiKY+WI0SaGMxK
I9/Rt2p9jvgaxws+ak5k3HwKW6jpGpjCIaSGuyysV4M5YGNwFrltVqK+E0pwO13Z
zUuO7qZ//Waw2+eWgSb+zbrFu38DtgSHWSduoCpEVguzDK0oZ5v05zKvJwCoVl2b
4CnZzPBwoDXYzRFGkutLd/hPNDPT7VefiYdiJJX1MBndljEW/n2Bvhv0le7m3c63
+edp12v7Foxtk6VoxFUSWOLZ25nZniwIUnw1f8uoT9Kg6vEUg3qrjfw98B913T9l
dDhO2SBEeBpBeCiITRokYV+zLeBKonXGBY/hvE4/tgg=
`protect END_PROTECTED
