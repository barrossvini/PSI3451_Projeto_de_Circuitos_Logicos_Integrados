`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yEQ7P1Iq+IT5p87gPwNz5Qxs80gtUYiyTUVlkNZNPjwKMCqj6uiGv62HMQPYOnGO
58lE/zSCQ0eOzcPB3gTxJRMn8UBPza/KKo23HqM0dGZP6anVglcjmxB8c21M9uOJ
UDT/gF//ACBKlMlUOJ7f54hNd2xp/x8CqSmWHhW/ti9uZL1vnVZNaErrlr2gaeto
4jjX6VyCNWZlP0Pn88Av0o5W1URZblH1+rshoKxJM+yqYGqwPNhqV3YPipZB5IG3
6FFIgPGNOiMDk24BJ6rO1FWUtNS8Ij06GMO80h8K8ZvRxk1SLFmZ3CzlgUV5x26s
YrLaCSahCFgqpodZ93E0Zm9OaLYSuQw0qYG6MPPSpOfVPIm8w6baUMoskLLrjHE3
5tQ2Eqscup+6NDYTKOHJsDfr87vOmAoXbdc8cUgqRIs76gcq9P3VZ9PNqh3lNMEK
BxEHJ3/k6+CjHEoGCOIAknh+EiJMsHu0PVZF3MoYU0y7uK3UAEGbflVjAjLA0R8a
Ttqgd4ruUUB3A4VKKFpme3HHHBWNv95se3hue/eEu5UbpTPkVSqaDcCJmkQ2lEtz
HWyr7IGv/jhM53qDpEJrpb+/fKa7nrl5muwFJsDMlyVsQTsHdtY6z5zFTIA/Nq2H
6m3pL4mJf1Q+KxddNyHkEVaSiCzhtpZDom9QzhOFWVoFtvPOsv/j0EAf21ctyrKq
oN2Gk0QNhhgy4ml1YXimBJP4ynAcclB+QD12my7w141L/OS0p3zxM7gzUsF+fEO5
HEgFIjzrXdFLoGvzytnRiDL9T7SdfQ5Qyn8egKoek0h3ZEeLsXmGoXoODt6LSyMW
NovJMWgbQwZok9SjoMeL3lHrRLbvxQM8O2WG/1wpePhrNA3aObggtK9WsORyEN2s
`protect END_PROTECTED
