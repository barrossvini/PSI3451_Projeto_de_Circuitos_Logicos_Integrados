`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ThcqgHhWaNnnvMMoXedIArQDAjcE918AQIc8bTOImBRf44qYfH/OMJNtEpZi46Hr
EKPvW29zNBfjbrkskXNKCNYeuBe8Dv3Slph+4r322NjnPY21hFew1cRSBSPWsJ9h
8BsEHwQpGRb7nKgFo8ZGkvXCVIh1nmDuTYYuksRIBIP6AB6Ypx/YB4YyiObBTlx6
KMrHwX6NqY/JPMhVaYpPFaJkZ3a1ZgZkKnt/pTL5JJWk6BNJ8sRjqM4PLdndzE7h
peIv5uOpjZ0+HNJCJVltcCia/tk0LUsa6UUrDyHgnSPMX9UVNUrN9OZIaIQR3vJG
UL6f9itYqIo4upvObMvaUEnNcTkF8qqT2sqwliRAjzE5GnMKjpBWpaWG7NbawYlY
zFTiDHliiaDxU+seelJ1ShnSEX+CcsxSmW8/b7mcNduZRVVkuLbuAV2F5RhK32Bb
050/8hrZaDlLQtMVJLUhyNZ3ePFwWgRGUN5m53N19CuAFpdaM5bQpXuHp/EEpYfy
dga4ih7SVl8yeDJsJRNwyOJWFbHQWSRgnkhkhZ3fnekn1gaizylwdAKEfZkfTBvx
e3OPwDkK1P2A8J8759JIiX/tDGGeFcY73yY7OpYPdXV74nM1jIzobrS8MuJglIP7
/NNGxMIyqULYodEgwnfiI0WIdJCz0pLnlFhL7E64A6zGxcO0cbwVpAN4/CQ8+u8F
nYmKSJAZp4cbkeaXOsyeAnqnD/F8maJajzUj80fq5bkgScpHuHMBGXJfCcUuQJzr
bjtOJHJQ8wdSBMPTWzI9w5docxcNv+HU17qbZfLSsRgC1Mf4Exq3zo4qR0CH0rxW
ujXjbZgFWZm2Zy5u/izqv5fW7GOmkvK2VFx6y+rKK7wJuEvU8SHpyJa8Pxm6lSct
naJTm8ByyW849g97G09mmuQ3JlDxzyWXFaSBhI/XhMkNj+0VsuMnjjx+sIkv08Ky
fnaFN4Q3kr4UVHVGqRiT8lBB77pueuQHhPiAoKKR7DhrByFuyVr5tcZMbEGUOglo
jWYQ3cexLtCCj/j7d5IvW5zIjzvBzDMK3ioNX8YiCK9eD08PcJ/5uLKUuBm7r7sJ
cKuqg0o0yh7jaXX7C26ZqZ3VIaTZBlXXZg1u/yJDOEFvzkxA2tIopsW3swse3rEJ
PgjItlObRoiJlcv80e+SBtK1TcB9O2KjU9VMsZJ3s18Bf0WklOeLF/sgwCHDJSpk
O6eDfLK5MDpSIyyPZJa3ojRr19ZiPBipsWDWjICtQiLmRTDNwBAz+Z7Wucy3fJlP
`protect END_PROTECTED
