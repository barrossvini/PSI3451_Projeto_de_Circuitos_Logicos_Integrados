`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wHm6d3NyNtA9Y9RijrIFGXG20goO6omI0c0y9LzhxT/tqolEDpGFjQ3N9m2cU3tl
X9n5BSDcNg06GScX4FfWXe7N9xP5NEpLFlGm/PUOfAx0JUHdNnUC142IRo3Q6+s3
ArcRqmsRO5mBervw1B+RblCx5GI1UCwXKH7h2VBWoOwE9WGAhM5v9rtu/01aulDj
2D80VOf6aanvW2ftJdOZgc5eZgPLaaDpZniApZuaVXQ2tzL3oKp5GPLMAqJ4A+EX
Dr1+suCxDXVkOlc7pHUo+UTeHwUxvrnbuiNVK+/WMD22I1NP5H8FEnhFc/ak1VqR
wSmIxD0MNKE/i8CIZE8aT6sOj7A955DHMNYHDKGN607ouC0CrqrIJ0ZDqVPdUo2M
AZMm6coMNypeqw7DQ5iS/5zWWA6Xb4PfN9RJyKvdlPeqjXXJw7Qxb/FZVZMhXRk6
6u4NWOS773Q6o+rSy7VrRHhExNSPpU8MLfz78Ep6DbEbVtPbz50Pzv9f8NzibFUD
wmCNZ25+yJMNSeQjCKgcsi4n7/6hbc6UFIk0vhRBYGBvllwWagnyklxdN1HM6OtN
An4wvjsu4i2WPMx40t0C2zPrkNZG0jD1RvBSFeqHltEb8bHILMvemsrA7yozKFzH
T+7RU8kZHD/3avx0zYXQLWTw0K70mK5VEffmdQ8DO8NlqyjSMgeCgWGQHAqXuuuj
cwm8gzeHkFX7Kl1YewitlQjgbUK2+29KnwRtpOf+1f5y0+lMCyj5Nk3fZDTGAsG1
Kh0zAODCLhXym2xoI8Gm0C7wEriO+LUVvxLlnQRzUTP4RScEB3OFKL2vtVDDk/n9
61EfmhclxEFbPU0uW8ZYHHSpMXTBoz0Y9Xlm98dz/hBP7JdiFjnKKtwK6VGHmulT
eipItj0kGVejWyYbUcSDMiblwhNF+FfJbPgAgEWDk9PsgHzMnuc9p7G/+PoBo04G
4x/yLZdFMclo5R7fsaKkOiYTgyoUP+PMajzWcRbfqUyVXo9EFwv4THsN6O7m0w5l
V1BJEG5kSj7kQibR0V5orsfQrL6b8BhGrPMiTR5I4kxOVy7Jx/2JxrGa/OSo3Ffm
oQ3vMusFkguK6p9OtiQzbu9CVBDZRUWjgEHcKqLp0Bh9/acOf9fKTvx5r6C/w2j9
1LRZXHyoEFBqPWF4qLB9pVCDyUPtqSc/JEyNln335z66pybw8jxYxuXsgqxENFZ4
+Rg645JuFgMcUSfd2UlWfdsfEK16oYk1zOluQxfzNdA3X6WCX6c+g7Sd4GDcF9lg
2G6x1lSSMEFUKbzoDj3ry6Tcsy/gy8uKX0h8oKUV06bBZ/FGk3P2FGgJwUtZWBt7
KX3WChbzxysZiEPU81ph+5VHd4DopGvMHy92mH2EZ0njNI/DtUjdH6B7zRnqY317
M/fnS9KUF2BnwugcqvPp44DlMMeJHDdl7r6LCMIt5fEOPb1NBQ/qfxTWap+PCsUw
5sKHcInzIC4UarM1yIQUSnsBWdsqZMTzyzqpdeJuSZBCfeJmpo0eurwLGmAgumfq
ANbznMTRSEH6tbDOk6dGUev1571/c9tNqLch7/qnwysLrD83SVVkHgdRkbc5KU02
DztWi9FqCcYfVVtXAoDocecGtriMCKvEZ3jXm/cMEu0zEug9kI2ENDyvAipDsBpV
PkEy/VbcnfKqpoxiTV0Lhw==
`protect END_PROTECTED
