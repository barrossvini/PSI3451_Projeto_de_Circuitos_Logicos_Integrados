`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uw/9P8dZpONjQLsuPbyxpqSzgQXuqzekxmgBLobt+Xikm1NFei52oPLes3V+CClK
ZxYn+v51OWZC6MxOncx93uQ5dSPGulY5vQfoy0eXlOcSTcyK8ZFoBw/uD3z4aQrX
tPpXf+Kwz6lk5LK8MBsCDhsQMOXqrBALBRHfd0cPAJrGSLP4L7q3GObsCbp4CLGA
Sc9AbywyA9Lbka3H1Yqc3e6i+eLjkJ/+vvaghg66LylGdwI6MU8yTBWxe328AbKg
xpxYTt6y7+902EfDpbUGyKNYDmcaByG4elfcgR9ZUGq0eFHbsInkTf+2L7KafnlW
3rtRKlal/zDMLym1kGebI0gE4w8vMa+8XJHgtWa3hGJrNhVNr6Tp7ElhZFoyyYw4
WSFRpUW9KCmqLEIBQsn8RYDY2lqQLUbkYxzpUnUm5hMCx4AohBFk3UTXdFbzSkgW
CuinDS1Dq58HcdwXbLYR3xJgkMxRFAYDoV0zhZ6kHwWoftzkYjvVt7c+KEVdFQUf
GCrBguonFUPZn7j2Dbc5BHN6Pzij3yW/cLbG8UTKfr+2XbZmjEfbSM1kmUg/uXKD
UEPhDDZIkLUKi6dC8yM1YrwvlcMx6f0YQ4aiHdA6JQ5hZa1u8i4Cb790nl2fmELS
Ww5yRUWD7clQAPEhqR3xxjX2qh5qhxd4H0r3ps9VNQgd/i7YbheDJ5xJs/9iiXbK
x0SviLcqGtJOWv0+lQlxzer+KiWNwg9vDUtlkG9S4DpuY3kovZmwYFWuUeABJpxz
v8nwo9nFg7I+7es3s4ST2K1huyXraBe8cS0t1jUSwPgD/nte99nJP+XfZWPwrMA5
4j/tef3cxT9RgvTfwVEb7aW+LyY9AjQ3bkS1CXZU3iXzE8fA2bAK9S1vg3GtzbR2
xbSmbetn1jM9aSN265J+GAKw7+9gO443a0V0rTmV35m923yJMZIegtmkuLprVmM3
yJW7miMTOd3/A9K9MaaDOCQw9uYgOzS/0PvBiYm0UnPeWO/KaiotZOUPdmkPGHAP
NQ/vqFo+7Nk+7P0S0vQ4Lcn/+XfH3PgpaABJtqWF9eMr5ZxQjQUASzOu61tWjepU
3j9hx24RA5gOeEUhN5Wi+Y2JyfaNCXkXvzttxcz5iyHGZ4DZltyB8r6Uhhe03tFf
cHWKq6jn4324R42Tm0ryISoyQT8oOk63H+yEhI0ZimaqBR7DpkxycP49pTi23FWX
bLddag4VbjPMmXvelju/hSy/HKSHxn2lvV/94MAwRobpRBnSSojlxmZDXCubJh2E
`protect END_PROTECTED
