`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0HTPlvwKY0ik6Z5t4ujqDnc2hVsqum23t9o19RSW8i8b3jK/BdIarn2nfwP0VhmP
yYGqNfp0C69ntxTDYuHJ2kfD7AHbsJtGBw9n6g5zhPxxJ+gEdOdx9k+Q7Zv7NWOS
xg0PbzoOJEekThcRsCSNZqyJNlzEnDEPDcnmvS5YWhMf5bqEH3tF9awwz/jmF6PS
l1PrZWdHNrg/oroousW+QlE9H8oArZZFAm7ShYoN2hUfRQQzQh6NPeqrLd/B8pA7
IeDljxTxRakkTCvWiKPK3QuYTUUc2c3LWGZIakjBKE4i7qjRkGu2WXc74gnHR7D9
m5bN1ULHjc4M+TuNkvloQQfQM3JysB5UbxBrakEAmb41J7gHeSALbcEWqO6PS3MW
VdSzFFRgjalJImREN+n0vzsPqjrrQyRF7arHShOwvXLoX9DHXjno9Kml4xKl1Bo0
KZkeAPXdsnhVpio9KG/kLK/JP+FuigHxmoQP7r+b3eO1Zfur2BtMFbWK/jkLRg0U
lNsvceBJ3e0mFYtpW8jVVCh54V5ZXiro/ugP4LuH0swnkjVz1Xg45gHO6JOWk4EU
fbA2cAHNN+MuiGH1mFRCmqmHBWj/4y4BL4/6xit2wgMvYFE/2vXJeMgA1P0Ow9+9
NcESuzTmY4pd+1qzDpKUwz3Syjiu8L9iSd6suLaHCO04ICW9rCXnsrYz1mr3edkF
s/nZxWFW+ZY+0F9Q+92v0WgcUL27DSqv74iq5A12oKlBblAGpI+Tonpb5pxaWO3V
palgffqLvEHaUKAF+P/MeNJO7aOXPcteU2iziy7kY8P9WfbHA3G0zXmg4Mad1grZ
+jud3I+wkXezFLlRUtecleeOGugJGC2/eSrLdJYlJKv4EVfPf7w1NrrQ8ICsbLlK
/nGtWpiavL4MpHpXnAJE5JJn1Nl3B3Gb+x45GCPZr11w4N5qegFsKM/A2oxFfiM/
r/stlZoXPU35xUinhRbZJxzaHTUGNGO9gcWbqwpGVr3kEgcPVq3guhB0Jhy/B/ur
M3x/T2R7zVirNX14g9jk48nEd5aTzHFtEI+6tVsRRUh8jv64vvuY6kH1488+BESn
TCohFbvxybQGkYZyquzd5qMdkgoJQ4v47nbAD+9++cxnk3AyBQF3PDfD78V/bWfK
2BpDjhi9+cAv1NctAr25sxzVb3ZKLIQn6BdH2O8eZfEkg2pTneO50iptKrih9dJM
t3Dz7ix8SwDhbX7BXJWIS5MrtvchYUJlStRIqsz7tHiPSPXai9wMnQAU8/DP+UAO
aX6vBlCV2yVXEPkgJS+sEoE3JO+STLUP5UbaEfjgUkz4anNZ1xu5QwCkBAAgWsOY
CULX75aI9jKj6GDeqcl5M5tlxafMlBZ7irEPBpZzm4sQP5uJuCHIWHvwNDR/bv/b
95pUFEuzn5Uj08zeM8tcFfYTCD2XQ+NKaGdGDuWDOmuowO8tBY2K0Njtczlt+SAF
VAyEyA00ZYqDCIW3VymR9T/kRUH5a95P+6fNknNJqWTKRaDA4fqygW5elVV/uoR0
st3T+BJsNWZRZenkVhkxjiOsAdJy9CvV6Pao36irx16ehjX3vurUa3shCig9W0/d
KV/CF293qe3mLye42ozSI+WyMsl4E+vDbisCvjTW6xuf47brcL5xyUW4xASIrGVL
pstzV5JplAZsViOW0mYdo/BKJbGbfn5fhNlJQ3/g0mU=
`protect END_PROTECTED
