`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e41v5vRYPDIXeCPHThC80wbQsPTnXONzEj1aL/5vAKC+mRokmgPK5eg+Ug6rf9oB
cBzUuuigMCLJ3WkTefgXQQgiQFGpSQ8RPEdXabOD+wXkr79H3QS8sogJltsRqPXH
96zrokR23/FlH+KxZ/OX72KO1/rRZpIwLbpLMNePcVyo9G8bXVfbX8GLSuXRVoK8
S0slTUcjVmM38Y7CbA8ryp1xyctZKS0dzbDmh97B/3vCwtVGKSMybN7NZAwWFw6A
/J9Fbfdf7pZ1GO3voy095Z4GSGUYPCfOgLMvE4KHSuphE4F3P/0h/dMsKR+Dend5
uhn2w5EcZfpJ7tiANs8QnU5ZPi0FkqwDEFNw9Rfkg+CBJGgG8FndcTiw1GEdQpM8
1NuplgLqKR99DAa3+PhrGg/FIvHkeOjykM2y6lXAijLIehOUpechQKrKvYJO56st
9EX1CnTB4XRZkkyI5rQtiDXV8vBVNBa+ZRDOImjjwAM7R8HintcgObcrn0bV8ASf
5OBnU8/y1Fx/eY92VpHddiLdQStBiUMDvhank4LTl2NhXlIutdX+yJSYtzknpO7X
SP+lxprq5zI06AyQPewf8AV4c40QL7nBAwbwL8UVSmXQ3iVCL7VbB1+c3A4lhj05
mtzhFkI/763TgS/HikOhF6x1yGZcmcddX1JMyVRS5Gr6b5mf8twDHRG5cWDPctr2
4luGsl8sq28le/YcfavOrH1Ap38J8k3faqq4UVOvUH0jGtBBvRTJCqWECrX0F5DS
7uw1HPRwJZNu25PUO8qyC4/pyKeSQdLOpm1Fi/74fiS27ZrKxhcCT0qoazzqIyYA
VOBHndDsdvNWU6YiQYBxvTle6M5bl0oHtqjDVjgPsWvaiuVkEjFHz8H1i8A6FPFi
dgCEEfKKzORK2+DBq0hMxmysn6XSIGgjMG8GDxDSi1xR7ms91AnsffKySkswbYZZ
tuOnlxL3uuOsvhcf7ADfprPxccpSA1DppAIE0mbLeoA6tCDnJ8LCXc1pgOx5uP9u
2QZPc7CeYdRclzRfc+F2PnPqX31EwaD06nn87WxL6imtXhquNwy9Jdj12hVSuJ/O
BZjAeHDMEP2UdyZfk5Z/CNvKzvYi06kjF06AI8jBf4m0R/vQNoHVuEVYm3WiisyM
QbLkKXycbsqOOLxZJg0lnU96dUvfF87FAEKiQD+ptBMvDfgtSL0wwjJUoeDho9AU
zGSZ3CbiXkAgVhofR7NOOxT0FEcTOcWjwvmIDRENJmM9oCLJ0kbBq+F92VN4B33a
Y5El27o007HCRbKF5AZOAbpNCi2C2PTKSGSnQ9if+UZZlQUOBEmZMZ/i+/THvQ8L
1VcYAhxJvg89wvKfIRfQR5RSlnODLkaP9dhGSOLvH6WvJGEw/LxpXSjb2aTzsMj1
6MQkKziX2Uzrzf0oIBvQ4UWJEDs0jsZyd4SNf8kE0lLHADN5aI3oQMbl9DyF0rYf
cUEQDD214Z8dyDdOBxPMVUzFUGZCU0yVgqwMiSLtSymJfM2axBWg85lCimYPr7j6
P0vdrikELr03ECb/bWm6U0EFj8NNiTxhfxu9Y6m7eX4KZ4rxBaDvSLqlzrqtadQ/
vmzTTquP2N/3mAwIjgOt5xkP+db9dj/+GCQ0BIrs6/8VP/jtjbDSa5KSYgt95j4d
eaqioqBDE/26PjQNRdP3fBmARtGg7ps8GPgLVEhR1ro+zm3lAz+AZzmy58J7NZ70
uqV7lw0s9JdkKkBSmD4RXKUGMwK6Q16N1mKhom6tNANd0VSmW0W6+s6L3tA4i3Ib
vxy/DVqJjwU4vy9tVeS0dO1A+7ZnmElAxjym+fXnuc3fT+SHCxpeuLX8nSPTFu4R
Ylm6oXGKVrhV2LoU01c4qohfizN9xm4ZKmMG/9Ejvw/9m5wT8EwyuQygEsXBVAX1
7bpw3GfzAYv+xoHi3dSI5Bzc8XPOwPvnMWPdhYmNJ9C0bmvVL0LtaYLalA/Kzc6T
YXSSPLulh9cCSmDBnmxvvQI6DjyOPS4fZA38tfq7ePwsrIrNIp3Z+nder+JKA654
JCNTAAQ+iqQTqNn7RxwRN852czFBseoqCVZR0ySmPx2J+9tzrtJcgJzpB7N67jiC
UUkHWn8oyissd7C9OIY0r+X70rFqOVoHpEkXX3j/H5UAWnpdlBYyh52lZCfiVigo
/0Hwb6B4YM64/XkNWfwv+NYsOmyiEFcyNlIL+IeNlpfIA90mLNw2zZnbfvjRnkhx
7L5fr5Nk0ERp+Ium/IXN+cLcIMbhwFD4UJ31DHJ565uEfi4F4ijW9A5GK6XMKEnP
JYqFDdqWHsDZSv3lqqpO7h0yX+/C6jvILcNeuR3N5qX/vsSP9iiT46C+Fe4nlHUz
`protect END_PROTECTED
