`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XaAt1uP6lcxFtA5BXKPx+nDKyMD8HwbtNgGxBqE/MPclH1oBSFiKlCtUToPl+LkE
00VIPtpEv4/YPOb9zpASGI1Q7A3BGiq4qU0i57tr81OqaSKhlGMTSsd8KmppDb5Y
SoKFBlZqBzPHjjKxw/kF8BnBwQwUhJLi0Ocw+g4DGUppiHnpGWIWaOo8jxas/g2A
26tVW8dsszgniclHIsoA13w8grnR1EZJhg91KwbRN1kRN4wDp1yKYaAfHwfxEd0X
P0rOl4uONNPd8HkdPGoKn8jhwTu/Wt64jknCumEPOv1YWb1AZixKSxEfmCO6CUOO
sqoVVzUdHUph2NZ0uGO9WQ8V76PMEHlgHHwI/LMYzIQc4zfA1pEzroNLaSZdAWjQ
HwY9hXWRh5cMSpwEbPJv9mViBUCtd5WB45MPBmtjGVr0pAtoUIj2bWhZpHL2G9lX
EHBgahBqS4E7hOwlXBA4LhjdyaReMBZzCo7sihMlE7qTT73HyR80Iu10CDpfJcn5
92dxJcHMclvGhd8b8DmXJx4q1g7mFKo7jZmuzjM22vik3M4WbBJ3xMxUUiyTgruK
zHPzlHHpChLinqmCYn8g7lHtNzEPBvbxcjjr7n312Soze8hPm/BUzOrGrl4+l9jr
HdUzDxbD2oxwiLm5jE9puVnpSvY/Or6ZAa4sFW8rFtGZOAVAxQm1ZVGEuVAIfYvo
9zBVVlW77iDPi1NaFjyr5jgXdiO7eXNWJF3vLaXU6uDjdVNsWD1OUsECcp1HKCDY
7+Ecar/AcnflaO7Ydl8mfDTcD0XDXxsqrOskhD7cQUwM2D4q/9GHmaksWKnpAnL1
H9mfVTRl6K93BeBnsVX+gNeG/Kmz73iWPU87Kn3bI8nH0Nx4kU0pd823xx5xqYsf
horY9SRBatQWLgsbomCUn65Yqld76lL9eJzIvupAvNboB+Inpn1YzqBZ6zcc+dwM
It2VSBe70iBv7g+Gv59VbZiXE4sw1+U89kVdlcw9aq5Zew5fc6SRy9sdce3Gp1sE
2Yalf7RmwPVuazQWQIBBZQgxthm8tD79wnYplMwcGokfmAhGAWVt9RIenjj1n0qG
FUrSHqzPeKrCfHv93UkkyD/CUO1Dt512JDXUNX8Hum8FXDwu3mNsJpKGylFrFCei
ktAI0i9ENyXUkRQzg1txr4gM/gq6dYhwFATrJyZ8adYDKVcMRF37cdETeA2L9Boe
eOtoF6LaSRCLcoV64XgNzxMJ7cojJS/V3YbSRlb3LaQ8lPuv2tYsXxVeeLX35q2q
klxNF8m0WaAfAhYDdffZOIoLcHNSVndM+K1qWPGAO5OVneEfan7SxlV96WgpmnNN
v37/kq+wreKu66CXn+k20U7AdEXTPkRSBT3on21tUZFN0cGGBh/R/krqZ8bf9Z9q
DDyE64uy8nbpz+yp3GgK1rkGzCPtoqqz5gmBSPEJcIubva3f/KN0/lNYRS3Pi7o4
aM7ceFS60jRYLWPbR75pZ7c7LBGPi+OgFRIAItQqAl6IPi4t8z3KakVxbEPIEOY6
+UYP4TZlZPHwS9tw5r+lGbQJbU5rrDDTncH/gQR4JOPKH/RqMqqmf+vQa7rV4EXo
dKod5lZBanaA+AvCFbNHEP/G+YeEGl+ZEyTtIVy4Q3sftdw2aYKDdwS3StIZHYAQ
oUSqHcLHHZCU3IoGZE18UuTmocM+ijdE0n22AF7QSTpCQsPrytGqp2MsNOOvHd9u
O+g/4rQZPNQ4jGYjIKJ0aE5Dg9JPsajb4PGZM9g0HJ89nXbSEIRfuWecYcEe9smU
JurgtGeP4O9AZx0kacndGeGusBkGNKT2hwR3UCBJRiDIg5WBMx8rpq3sTXHbpfPz
4q05lLsH5i+pUKmsBSsc2uEd0eolk/hcqBmCESALMcl0/CjANRFqJD2x2uyYyaT0
2cm+U0Zsg1ZPSpU238VWLj8fUw5o+iVGfSlC790HKmR0TsdcEFOl+rbSYK3//4lP
/cN5cfYtS2SWPeNm0h0m6ZUxqHMdtdTObuKa1qawB8tjKspnupAQc1zTTIRSYHQ4
A9gZtW9MzA9nd8EnTt88l0Ua8gFH0r9EarZ8OuemfD24zcS9f4ByuLsj+SV2xJvL
bGi7CCFqf0f1sG35Ssfw9COOpkSUrs9kMWmqqsHpUK5Bb3II2CSM10iWBr1HqlQ7
a7zpHqeOOITRpQu2lAHRac9C6zRcCC1eElN3ZA2NGAHd1RjH1LN2UjnnkL5yhaNt
9vLxd9+jKL7CQ/XAdvO9L0utgrniGI7aMlJEoBt8Nl2F6LYg6OaHkZiEDv5X4tHV
JwAQp7Kl10m/LhAvQUglYMVDp7stKAQQO4yFi0jsqM/mBmJu/l1ZDbmM75RE9zoy
Hb7ZwevXpJh3O8sPqZrZYOvImUh23HWN5nnamHzltCJdckbBMCdtrkklT5JkCiV0
CpHFd1eWfSluHx1hUiAYPuLDKvZL75RZ2TTz4zvrk6KdH5ZCS0zAj+oV2fZ6jAKa
TU1N9wxgNYsJxSjiyYZkF1W/dPqoAgICh8V7C7IKfIndDqAEOQshkt91Hes0LCZx
kx3Nv8QmABxmLMWpHAS5L+Dvsj2aG4RgYJPoYl/+7BGpYJg/4UHAa+tKtmAtm+xI
TD0oxtKfyJfHZV7JWUt3Xqeq7tjk//xP/c693FbjKomLOw2DBeh5iiGCgLF3B83G
Hz8ObYbd2V06Iq8yBf0avBIJ4ko4gMRnRPTs2EKzpzA9RTjH9OU0S/q/MD3QtxXx
WTnrIE+P/XJ6AI/kmH9X+fprB9N7BD/cR2z8EENpa+4xcykNsXdKXO9LY25soiur
Zk7jKzj6qOPR9sFQAlPxNenx7dT2GmNsLYXFiI0dYvIY+UL90YGgljO5PMVCYtDe
XqveBNZ+LMkh/gvfg5IEnoE0qRVrFSUGz/WbZE6UHCHcEIjeq5L7hMdSAJOTD1GB
VJcBK25Vm3umTXcPxUg0WuYkfaHw4hjPEqIhhEhLwTP2jBC5d864b494IYMjQrn2
gKNXNOG2PVmX0/BwryTrsQ/eWYDK07A6TdsImuEj83GVOuUgMvqk9NJT4anE+a5u
qOa2u9vbC3amk6u16mnqKPSAArQlym//eiP0Yx+e0ypKwO0BsVJ01Syf7Eed87TD
tJsQ5UhQzeDB+s0hL2SYtKBvXqhO19/p2sIgh1JT8qSFyEdOhoqQ1Kix2srE6vRa
MoA9kF3UfxhHkz2ZBXuYkidSd3n81iXqfeQOuFToEZHZCAZhB7QcJLXl6fMKbDIJ
Z29Nxqrnfawbf6qta6NgOaUklUCG3TzVsEitGXKShmgtXkfYLyhT3i87vkCF2rPp
k/5BMOr/Ga1XAr1KlF7MeLLH0hOUgJqNyiim2MRK3Cr2Rt0LIsbfVdQg1oAcj+vZ
lPNQD9ka29hqVHoq33iL4ylkw5SpCt3IEcSsHM5XwKZgGY/Z4ljx0zOrUK9ZVONB
85aiE4R5oOnUmi7TbpnsjxyaVIQwpeM0NRXm+sBZ1khCa/NF2E7gZpf1E8Q9mDB6
u8VfmcRqQcT2um7uTSmt5E1ReLmNabdjoP8fnc5XAnMcKfLso6X98aCC/pxxj6cX
c8HBD9p9zCWm6MgEjZJfrRHkFvKe9sstPGhmw8W72t2DKhMBEzTTHMKCyy7QHDrm
`protect END_PROTECTED
