`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tq5sY+SIGY49SNCQqG1yinoPFcujac/Wj/hnpcKyDWkmb7qS1twBQKRW4q6a4YxP
hW2lLRZp0BOIv2k99nEyd+mVCqYg5ozF2uZYmjmKq5RY86hzYjae/H4jgPc8gn07
XEO+tekmS5I9Q5qghcSqGMa1NJka7pQEeUaf9HMInHLKaOOwQR5DZJRSupkZTBe3
BM3X0yMCFcMRr0uYMhHX098BfOxVaiCoB3XxPSoo6BsEX/H881b0i+n9EEv4WMJV
YUL0foO4hRQ5ifxbfBEdELUAJWsITVMJasvp5bwfVE0hf9Nh4eu5U/oQkbjPFEtB
uLoD9YL3OKUkO2eY+Q7Tuj8Wb4juJwI1fhF92bsD1EvhmQbiOhjv6bZPlyernoJa
vup75WoOInsuqYg6gL+Tlq81437kw7zFqKEO0PEftASNzngkzX0pN3gJyg3YWKzu
AcY4zLwwQcYC9Pi6pEegYj60gxaS+gZRZH4LOjiUmsbKnMmv0E+fYE9Np7ChbX/5
nXA3wk2JvPNCUKS8aaixIxrfintlefkDQ5XuwPQzvfC8YcWkJf+5XeoQjiPTtEEP
7c8WwMpl4+rVqREJb5Zthe4BwXc8rPZPjidEjH4nujv68gXCf4y2ly/DwtUQDHGb
3YVv11zRMmVEMCFLXA1VMqkx0SG1Leq6shf9F50VE6nx8ty4OPf94ZAGvchG5GiJ
e5HBfHVpPk5x8AHuEA33sFTQy4yyQ5xQWNmXyCEyS0Zk+LF5EtrQ7Unb7OhmkjTF
DSQAxZu+KUpUBw5TkeNUPFr2NnNYfEbXj2NMaTZ3B6Qi2dk10m8mdnfHmGN9/AJ6
sD9t9hF3GoUMhhEgdhXZP9AB3LqbB8kcaTKzXZPAPXxO5Ipk1bFF64mIzFuM+UiO
Z/KLs4ZlsVlYLVksfLNC+xXj0c2LLEZ6YGg8qzfqlrHHackD8ybnfEVrAWaF30l5
0dlDjnyTS+MKZxOz1GhqUftWGRDIPscUIMQyNZSEJidUlYX2tJHU51iLTrAK7tXO
82v9rQ8asgro1bw2kyV9r0q9lx9+AqT9xRKFAOPK+DJMs42lg1e+qafkdl/L1Fhx
F2+RClbuMXTYOx4SmpvhjAFqaJY5iLOIgoA02NpnDgc2/dpeW6ABJdPFHTmxBcFb
Q3qyOt5EAmbGOmgj+W8KAGGpFDX9BLVXom8KHK+OpfTLYxp6RGTXuR3brIbrUCDE
7meQNPIBefUJBL5UhuQK5dBSGFhieOOks0xYJj3PMVdRjWKwgP+WkinCgA6PHFIM
ymb4z9jl1BpyB9QLTIIOpernR1VYq/IZFIuHAF5jypOlzg/Inn2TOIeQlL5ZnYyI
uUSxWPJkjZhu0Djrd9yyusEKjGdXB5ff/9Gl81O/Vr/KSA0zOmbrYjQG9t5kx/4W
WLwdX64Xfg3Q3Iqwe2C+S08/LVe3ykQDerhXyEDEbv+OIGZQGVTDDt3atF4KbPDa
OYdrUMQ0f8mvu0e9wFokmD+E4+h53UOkYxZpGQIlbMGNox3FQAmfnEkpzQIt2llV
hnZgmUgOTTQXS4XzFv72cJe96VXhJj7jTFwAt+a9yc2hPRxxQt13DNwyuJpaT9Rw
SjC6vHtAVWXF9IbHR/MVudWeWtV566vqkIWQkI1db7FLEFGTnJlP+VP1HcI5d9d/
hTno+kU3x39fqtC75OZVwgu9Vpcy/6+JzsYCzfeD0fWNGUiepMZ4Z/ndh1SLZ301
OTlx6b4Zws+jEmGpPOJtV5trIFyDYDJQ05sqYdKYzgBksmTuUXkl7anlOtvvFvgS
zRTiZ7q9v3t76CDq8DYmy9cooVLK7Mkrs1nMrnqVkEBUXJoH2Wdm0IPOfj+U2fQL
UyOnXT3FlwcMpyP5l/NCOAzlW9QtrxAgMzLFqInw5rr0xS5MQGM4SLN28MZD1QAk
xr1IDeBahuPplcy4qLAUmpyRMEs44lUnRsxGFzQocpyiTg/NaVU7JwZJeWDnoX8d
6m/OT2F76y4dUCJxg60ZrKQ6avPLB4itZYiIFpsHzBncfP96/K10pv4LwqOscWVT
nnq+au8WHuV/RaXRlnVE960hcMZBxMwtBfUvc8ugz8MFK2dQTOkxTDgbdoamzSY3
m1waNWq+T3bUK0/bPhgOdpyyp/Ei+FxR9S9NkQ5J2bmMrqEcJZK8u7O91VSV+CpV
Ig9TY8EyZ5uu4xXjQyvcYkbdi5WYEtLcwToaBhjTav+Qalh7dRs6YhLf9MnEDELU
XgzSuOjf5Qgax/XKp10yQliQHeTMxwK//nUcaqMniIQppbT/wDNdZu5Jn5oLcGyR
up0WopdMK9/yr88UmAX1ZkG8cMvCLkmkV11fENUwEb6uIAmVgVZSZdUST6xw0+1H
J/ISmJ/vKOUJ5PhSJCP+gXolgQIbEv/lK1/Tevi2wVICCcbj1nG5By58dIi6wlsJ
C6TtpUJouTwyiGc7CAKimfZ8MmgtgTneOAPAF115DTLfDMGgZ+IwGWwIuDIdQzo5
Tr+7q5DqXBPlXyexsy7iRrqVpTC6N89COM4bwLWs6A0Oaz6eY+ohOD+ng52Um6m+
BkF9clcPa9vAAmow3R8jcimSoF5P3WZHxidFxq+ev7TqhziZD3a0GbmrQ1coB8IT
IMm945ofB/wPxm7jjNi3oqqUowh9oRyPgXhlq7eNkJ50GXzBy2xrIAmxmdTC3OXR
ZXdlZ7Hle9/821LMim5JQW0DRccoEvPGHkL+9jwK93uX0dMjzR5fRtqoFuN4r1Ro
AUYCDXoMr3ZHcY2ZNNQwbgUg6euUUbSGscEpuDjUGKfCHvqOPbf+Me/TcrLV4ekx
IUfTSp3NFEAewuj7CPfG43stEZ9a2igOYAeQgj+akz/6vNeEIAedJrLfDeZrUnj9
7fmsQS0Hw/RbtfZeaD7aXCDdGhMuk5C8qlLX6CMO0SFkf7AdfpCmlrN7IDnzVNMZ
fQBO6TFsiaPX298BTC0NDguA9EXY7l8Hk9makfH/dFQKcNuXKfdHt2aycuCKi52K
FRHHyiNO2hb67UCyiWaLF1Oilu5D+hV2jJOznIjBqMZ8ArGu3DyypHYZGeoJuAis
gCxAMPqW4vlQVgmndkl5EwBuS08IzvQatHO/p0lL8y6FxjhY7D2bKTs33YQV0p1f
trcTKD+CYkoJ5cDHrZL+/920EE/kVNX8uNLvlQQsnjh/99BItl8Iv+ATBAhWvlSJ
omaabHqlFHTUm8Mwx5yE3LVtQlRH4U7oMkEfncLr4zABTsLJDPMs0gzG2i7S+taR
lKlQtu23TmlORUawVfB8L0oqrmI5MmhLUM0mdFBpZfyjTfIpXLPoqe9UQN15ii+n
Ez4bYNPP+pYKpOZpUX7G9jul4IKfndW4bxgNDgfg6GgyaChU9x67z6XYdhJ9RKuM
3g6JXHByUCkvXQsAjZ4jVFUNf4EdlPwvxldwsBnAbWMPVmQZUzRLwlc16bw2p/y9
0gKRj9EmJNKsU05VALuxSgCqWraZhaMp9i1RiFPhqvXzVQFZCoktZdV8WycHcira
fIZLusmOjB3WVdDBCIDxNrL5oyfwRUDpi6uPR1YWQZk98HEzSXYCIHo4RSoQUnGu
a9bvz+NNUX6zeDmZwGOge9wN2EIUObASR5kSn3SPwomifFekxRpv5vq04juJYyk0
eir8rpl5qxBKmN0/43kztN2ZvBrZSilWjT8ItMGG+l37OTC8NnTpiZEiWn660GSm
jY+v5LUhSTQBNCKbFb8QgaoWmuDxTIgvWxzd3Y7ft9w3x3aoKkYf0BBGX2Mjqsyf
QF1BG1D2uXR8RApNQFl0VjkyRfxEM/3yzSy0lyyG9EZ1kdT52nuSCkgG+eODufam
BaBQrbjtYDwuXN7BrO740gkPMYMaaiq+80co5ePPxscKxPEHaKuJoa30e45Q6TKn
9wIGee2jV804mpQBIBtsRbTP+zoVvsSEkk73TqL1ZHwXAOxDz6Kx38nbvtCk9IWi
rslWJkI0I8CCLLOPiNBigK+dICdr/XZVTGgRGc3mgUMU6fZpLBE2Shb9kqeynAn1
ZFL3AIRv6ebpmc/OShN1GydoPxK0qercPXl3WOhHvZFJfJy/H/UasfjIbWOqwnCc
/coRgwTqvnGA1eEwC/u/YPpeMrsVmTbMeRDONXyu5IuL7IliKOJ0CX6IVqT3iZ12
vveWMOzZoi1LHwQwjM9HibVn5B3EkJ7+0YLThTlhmSGhWnEggIKGGpQN20EasYhY
PCkf6rtV6hJrylXpSJAdWchO4EEfYt+XHqgB9dBbLaZTPmXfyD/efWz4F+EnVceK
ryFBQWC5K5LiPx4wWvFUe8U2cN+IeCOFUPQS764ceEnMffbDEjVqfxpnuKcaUmgf
A70SpViMLATWiaxugcr+uQtHp75fknTGEz29qncKR50pdgQoDQXQN7/xmgCpxFpR
/Xl12dxSaFdK4d+bH0C4NFGyFxsrhobh44e60pAp3s0lRS4fIjNadnBU42T429E2
cM0HDnGM+e+tG6OoSBV/EcXzgbR8Ydn4M5a16YG+BgDQh8f5nlguSeddidjyzdW8
y0pr581jVBxgpE2WW/9PNEEIWi0oaLvCUMwoButWqyO5mmvCm7tG6logkI2tsYnR
QrQZFq0j5Zmh/AvoHjBiCWs1mcNHQ3MuanmJmHvMZwC0szOVU9whVspsKBSyevm+
ZhluwJr9N1i3UnEY5S1kv8SYT/erQe/T0qh5nGM8Sf2vFM6aRuSXl/7QvGHtkQyf
TNALdZ9/VVwqXt/BkJm2VaFuyIDCSHN5DoKuuBd0lAA5mohUmWWyXcdurAbz89OW
t1gxV0mbgZX5juHDkp1rHOfql2uv8RgEb8o3pTRQrtHs1SzLs1eL6WrbLztdob6K
WC0572aeWHcyDgf7lwSuvjoSO6APUm1oPY2uWsqChdTvv5T0uE4d0DwQa2vD5r8e
6P7ag+xUrngQVOdhStLY3MjmjSH8xeWrHzJchDA91Fx3J4d0VV4euUQRpF8EM58K
ySQtQVw6PyLgdgUENtKRWWCynvM7c0YkE4WFUC7q92XjM+7O4I1qt2uhCYh+K0nz
D7c9/QGxdlpZq9gG/B0DsGKq6TrvJ5RcNG2veWlk1MIoGqhUD14jYrsSJ08Frhfj
+Rk1wrYYcIJql9qODavfO+5N5/Jt/jzMnyWG74or73lTooa33dBcd+YeaJ6WYFy3
kcS48Bc/jwrqyEY8ob/yD0Q1FGvpn9uZQ1lmCQyBnv6YsMWbjN8JU4sKFC/EO8gx
OO+fPkm6V49r+4KLiM+Af1pR7PePm191qk4446FO2QorJynbHoe84O0vjSk2QgYi
3fAzH0ToGydxjt37iwIxIZRyMW0CIrWw1yL2HO2FGOvaHMuzVDTOMugNFimTT/5l
hPaF62SkHTMf6f/zn1bOQabTfuhLur/V4g8RW1kXny63swkSSmKtEK7rldJ8W4tS
iSYGtOp4cE+rIUgdFarJEojcwUUvESqui4kNiz4U4N99CN3lm63RmYqT6q4zAHPC
hOJIRiA6zsgh+J5qMt/ioI2QEaK1yLxRWA9piqmfYFwuvGwzE0huw6sWS+k15gp2
PApdeuiD/FhvS7xxRISx1OEXCj6eLKNt1W/9sF7C46+k0pfVH00BW4G+KxBE8GsY
WG5orLocw4AEZ5lMy6BFimXdz1s+sYDItA+mj/NkKKwYCNKLz2RbPskMxavMwPhz
29XH4fP0+PrLv1OYU/U+2U+82nGbsSovaWP891XeGNqlphI5Vc+zUp3yQbAtogRO
pvpdBOK8zXo5UGr5zaddqcRso/yQgCzg4e1u2Hn3MdUUaiLW3h8ujZU2OeHYvTua
nC+jVPnXNPY7ftF6I5c8N1wnnHon3zL5KzUKSuevhcgpAQqf9qVymOIenbRkCB+4
n3pjfoyT9afaSqbRTHk9NGuWBH1DR0mftC5XNAuSEuQ07S6HugZB+YTLaZC9yLmT
XMoWsz6IAktxe+HeDREFfoRrCGs9yfxtGNh34TT11jHlHgO8h5FrxP0PD2/WSQj8
j9gW43hrk7SoRZKYdAxgIz3GGK7TbXBO3QXxLMQOojJcpU8oVAZLlvg6CcFRkpa9
ZH63LdhwBo4Dt6OzMDypIAocWjOdLFIfH+R/2Y9fddyIzeoW5CI7yjq72A5Avjbf
A8+k59wHqlUG3a3TzhcbBO+/XVP3J5b761ASysQdBZ0bmjvcREDAIkw/yCxFBFHk
BXtbdnrhWsFv1VLa/5r5WA0d0dMzwJbd2gRpjRiuchyzArNdrMNVrB6rt6rvddx9
IkZNCYHX5W8YWIcXRvtFqsixXhvzajchWMQ7wob2wnILNT2XjZ3tdxvkVsQMdQbe
RUsEMXakVZmk7elQEpJw7CuSv7Z8WXvPGklPzBfFFloHszBdWd9C4/yUc8Fj/zli
uuUB2Zi4RzR12ifPZngmEZOQQpCeA96kZ2kaqrsIlEmaxvr8R9yt6M8xxzFUwT5i
v3HSTQX8TlZqwNEbmQ+njmGfxcy/0kdBJYgLyYBepmZZr3Kc5lOs4NbVvORjBcba
oRK8fa6ZTE5Nk+HnnTIsjQnSzD8SfuPa4zOmi9ZTUlhXzEipPleyKyrbI2w4NnFu
9FLMg+b9P/ETreNdz5Hqq39NEOaCehJfCMBRnwsnvVSLYXLMJiCThM9DsrZBPk1h
sZDmMyyKtubp5vASUJ+Gd6xUArYJXDa/QE/yQra3EqkNEqczmTROouCV0bQ84t5R
AChWOBynkobUu8y2ZYZFioeBOjf2WUmygm3WZ4T29eQRsX8T7OhglWnCEBvUPruF
MqYV1Z1SmRiRtdZ94l3vwu8VHcP6gMzxL3kg8xzzqxRTkyoxDIXgTUL/DYXPFpgE
Hv9+xJj1YbT0w0gHAIbf8W3zRVDlRSG53+uj4iTuqn7fez2Gj+mg2WLXAfPqzfeA
ueIBQeu9i4qRPDf1bTYZRRJv+7z6DsjZIYTVBPKRT2rjMkq0fzLZ/pZABd4l5z67
P4x028aIaa2ggbMFKPc1ncmDoIAqMivPX131qQBnQt2h374K6XMJAbM6YJopAtdr
TEFFU+l+tkI/uR9+XTfDMUIamrisKWDGbog+t6VORO0AAZNCPaZZJMCzgG3D/01z
eun8kghxiMKxQntskByTyO76Y7g/GlXgOGrqRVTaHbWB/8KDqz6ddwyT0MHEoRf3
HKgJeXI7o2CVWVBBBqvL7mlrTalT/Lf6i7B+E5kQiXqGgj6FDWWyYNL05WkiHSI1
x8Uxsz9fQrcV0A+auZWBTyvqaEaLmal7rBTE7ahyXiHnye4HyyVzDR46ymFxuAsB
rP3lHEB9zG7Y8eXqT5y/CoCKWB1HLKBR+/970rsHtOyI2a/QYV+TxvuhweNb7tDP
DVFRzDAz5YspyHUx8kL+UxDZBFS9dhuRAxGcnHLHtZUPruWPOIQ6O+W9RIUCDoRh
zqzxpheM2X6YhA8jOM5PfNh6BPDduUBuJ9Y1sQ4+urRfKSyfbTGXzVslo5gCahS8
sUmaGiMo9JIc6ybtXK3z0nfGv4fBPsoQTLycsmSC8CkXN/LVqtqp5oGS8yS5wCAs
HJOc5Etn33iS5Q/RHi0WYpNQurieLoh4a3jA406D+j7zqYke17OE+gfh9FgRJDaG
6R+RstkNq4QtcSyn2+j78EZeUQiqO2HNjbhcThi1zZ6CCokZHohjoYOr0dy6bFU8
+zLoxVR963ANPcZEQXfifU9WBYT473K8V4+l5Z4QPFY9XjDqDT3BkDAaHGGHkvLx
g2UJrag4ysOiEk0fVCkDQxTaX8HCg48oeJZKqtj3tY9COCFu7YeUBATGxwlfW09q
pvytWXg38aDC7uLowbcuP+c+7CiB8YMJzvp4onftCnGMcnUEQKZTy5a1bCCgq+Od
pwH3qZuOIP6pwqhOSikWC6pcntnCWuk21c4lp8l/3w7leXdQq52r2ioGemZLZDFK
QJj8VDtAgprkV1dHnx8J8KWaOYSlL7IGycsSsgQqQW52RC6R2layXQeSg4zVDl93
`protect END_PROTECTED
